// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ntz3LA27GlIb1h8I/4QzK+lnwhCKqrEfeOruTT7u5nXwXPNhE0oMYkfrZEcE
UtYxtbUIjcPsbddqvjziofyrE2mVSDmsYhxmrt/Wxz7+gOBKMAN+qmaRX73z
UwsmJAKIhoZCecvY+1Pn9i2inSH9lZ07DT/+Jpd2EO9xQIsfgmG+E7Loy9l4
of/heWXB92NzEw2SAcVTLPBrAOe9tWTX9p8KjZZvmDymHbnq2GOtTGaOhJr4
5rkiHrNA2r8BYAzvHlSpW4wlK3VWtgv6JWJqNeOi0nXGsXcjDIAIF2OSDv7X
viKyz9TM3F+EqxrLCggz/8btStvoH0MtNJJyCYPAgQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AbNa8cUCMeqNm5ZFCdF9R2vD75Un92cZ6K3L94UrG6KPMmOgwewjHv+3GUC+
aM18ffk/6EkSuCv+d3Z8YWV46XUugmizcDAPo4sMbQWxzNgnLuSFKWsdnmlD
of6dgpiy/XZ0Z9ZnKuqTKhnzgPDZs70oRmDr3bNSkLBMG4iZJbEcvAcvCM68
TqJz3zWEKA7D1O6rQVoweH1kQxLBcdxQKIG/W1wdLy0OlZemPDYorI3dHDNY
CEqXnW/xQNypZFAkUzrjWgBFzT/hzWljFp3oFqL8FUopLsTHtQss/URTDWBl
hekAvvj24ZFOe+/9H34fs4JEcFofuwM/rFYmCI9uiQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JqWU0nmYcJpS+hIjzA4JnxWys2gAbgD6yqwEQisjYaSh23nakoi8DK7O9drB
+Rttidd4Y1NKlifv2Aqxp3mqrfh2fDZrz5V6CjpiOS/0hFReSq2NnMsgRw1h
1poP9oCsShY9C+nJTykjJfWRYTykBrrgjq5MpJkjA3COemIJXIEddvYscqBx
mdwx0aBSM/WXJVa6I/ARniGDwqVsW9B+ejPxF5JR2bMD8zLAvbgZP+kDPBL+
OviAs6TRvFYRkl1RiOl0pEqkznbBlme4+31j93PTD+zskv+PpdO6UZKVCsZN
PtyR3C5FbmGDZqZ+RAXh/wq7v5qaO66HmcqYndTrhA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Nhg/A/5UTYyn8fa3kk02lQNhgTK1OptZwtsuffph3ulBqY9m4lCrGxIl2SgQ
R1pKbuqo5ddd1GSvFcPMl8PmIeU1spwoliMaiBRoXOGFVK6ijfjwUxYbqCNK
DZzgG55lWoGDn30anoStsKov4DnKdWQzMwYJpmSDe3DghyM5HGk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XBv/apvDCUaydCzxqpXi2wMOZCBlrXMec3585kX5BSlosyMPngCfuF8T+ziJ
JpLJpal8tJTpNqP9cbea1CRPV/DIAUyQ45M+NsRepA19mCNkOS4ar+cqr1iA
lGPyY1TMG54zMSRN2Yzk9rTfXIwlMjvE9B3M+nkKMcUNVUOkVFHCUmDgjmM7
RxC6K8tyiMphl+SMp7mGYRkOYqp20F8HtHjlEHC0som3Us1tgL9kyG07U3mD
MTjH45/Lnh6DWqLhGXuERSaGwzZolmWatPAZ7YNyVcTFdal79rCHOunwCmYh
JQIBkXRZTNSLEtEgrcyZ/GJDMZMrkZbRiaHaRXQtSbwYCiGIoVpAa6cqw43s
11OcQFUsj51KOCM5CU2uRnLZhbjv/GkPadVEI55Qbq0JXVe3AyVE/P7VeouN
7iZ04nTmMOF+8degeIZZ8UZTFLzpawVUpxJ6ld4SUXSCbwJUA/e6ACHzaFpg
56DoI31i3euwaNsi/ewXlSDtpgFWeNgN


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e7eeb2kZ9ts7kHOvCTtSZ63voHICqWs+iU7Pe8ur9iKdPJXfX1DRU4rmVP1D
yoeDMKboKBuIBhWT5E++YAPQq/JNGI5hR3AjzAvVt/Z3SbhA2AeXZTeLj9VF
gKKvmTMBOvavTnsHoIabLhumMLTTCBKSwGZ3giMpYx8JSlONze8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XXscrPPLQEW122j9BZc8DJrMN78geXqOpzaZ9QMBPHlD0sFPR4RMRp5zr8/e
U+qxFnitp+Zc8694yNR7dhdZdRtuRk+mHqXCRjnXcf7swRjH9jhBo1mV5L2T
MYSjkt7Ek/XUUQpAxRzmOMNsYYjlSVK7dR9uwaknczra+LuGhoA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 94720)
`pragma protect data_block
ot7Dc4D6jcrHcwIufFsiZOCctjQgnM6UPvZFJkSQpdAwSX4pWhD+jbs4smji
GGyY6JBo/ZrsKJwhopsLfvF04B8ktUoHFN4oM9agm/4cdTN42SYqLZJLsJic
To3dBC1E8bYDE+OvgpSiN+zofGuOt1xHMZaICpwnpWoIT+1oTDAeJ1CRqIFB
WcyLCFjDKzP+BCO71nYvjWosaclXobZIQ5OSU1RWJJsTX5oooCsUqc8ZxBB6
qdRWITeu5xCzPoLDqZ59UYeXcYa1SsZsFBFqebGm4N+pjcsgkZSTyGHEkGEK
peJ/hkRUpTPFSF1rciIljBQVdaOOHlABl92APKLVPlMn86BKCqA4jjfhFm0K
bc3/vUem+YAKIfCNCl0g76kNiwrASU4ewaorJd+SaeJ6/KFwXZsf2srWWbpB
IAkl29kHg2Pf3valoWcshb79Fk/9bmPDLdsn2UykJq/WfysXURsCUI25bBcL
/Cc9QOhwbiHpkFhcYOriEoxXp3Wyv2SEEpOlvtXDiLB1eOwjecmIMzTYRKz8
P69fYxSa/g55WuL5KQe78DNHbqB21eXDnimEClYVqfbUu2WaTLJTIQIrx89E
wu9tY8TJ3bk3EHR0kn1L65kaKvqayve+oOvtzl3LlDY7pU6W9M7G5M+kp5AA
EvuFcaYH/HzW1MvFz+Iqk5TECXCNT/loE/e/2JJar5lfgeGL55ShyF5Cv3r/
jKLUPqF1aE0nU48yCsxKK8z2xAWEhQtHNVwsEgH/fqvlqwzx0LzNajpcN1g9
Vnq0PiQJjiHT+UvqDEGpprV+6jYCEIR+bv3vik/DGIRscRJX0cim3hyOVCXT
Q6noQLx5zPqkexHBHzuMIsp5iuA4NIrj75SZvt6FbZ6YsIbXoHBw5GgBt+x8
BEI2KBluh8J0QNSFb5QZ9xDjePd9f+pAfv45PAiVBp945CLS/+t/S7uJFP+j
f+MQswdAHU22Y8D6fsPg7ezpt8aevlojoRH/Lcwf4pzujnYFA6Vgzvt4syFU
FOkV21CLHIctkKPPdWQ5lkHDmObR3/JR63f3EKcfwps2g6D8XjckG5z5yPQT
JEPFvY7qoc7rdzR3CRQZv3WrDOItdL3ZrzzmQMEUuiiLRZualwwOsL3x5ckD
6iPUC3/WabcP8CuzCgTyKYdz9VXimQpyO4Dcq6fZqnMAbqsVQxrAVnUMNF9W
Z/N8QJfLA3LFRZdZ/cxS5IgH2yyUm9Y7K1/WdYfGui28f92AJFMn+R631HsV
5xv6ZbCTlequDBCycWOuUFFL6ihmvAyZ3P0KaG8bOO19xc1qsUvulF7q2ViL
iUUFnVTE8BOFqgDvQE8vNEMTxRebTLVLjNFHdf5+O79sgGA5IdkLrInMWE6j
OY6/MAMrnNs6y/aPqC74uO++5OP//1PPMqG4dLsvqXq0OQh9Ohr9AQTU1okO
TY2k73TPZC2YTf+04z7Qpie8UOZCfGBgpVzD+fA0KXDpIg4Ia+27dWto5RqM
am9ac/RVslZQQmg+a0qj+eWC7EeZOKsYWHzc23G/allu/+7ZFlksuLQo/Yt1
1QDvKMCsewdoK1h/uMG+89RM14rJKmjhroTUb9cWYt0Lt9o/w62h1fE/2U+h
y8nJcqL07jwOujBAIRZHspDrpV4kigPJtbM4W8dt/RVlc3TuiV3PNUf26FSi
mrdut6IB7i5SM7gztUKpYDISKGDW2amJt2VK7y175kyuBrzQaAI3qv4715qK
AQRPXErX2nn4u/VWPEdzVJluZdUDaPJ+gd/d0cY62O+Gu93H+gNGmD5Oca0E
PBo6KxWNAwq6tOTem8G3tq6U3EDiG33OPcjdaDgpyhag6nM60mOSam8ATJ8P
OedB+o5cQK4UAJD9p4E82ojt3A+RYPP4Lck3V/rotkZR1Bm0NmMpG0v6BlSs
dksvdxWZail2sfI+Wfl2lTjohc53nYAQQqHoUx9rW7FoKDZifxQmm5PBoDvA
a1cz06SV0DKFL+k9wX7M+9GJOhbzoferdkqRkzG3vmIXQaSLwzbNiosMIkSX
13jxiTOYh5F8pVAtBx9ttkrroBruDOK14xH7zEBKlFG4ZJiar1sh1Hv5rvBE
6ZsO3c6OvVm2kQtAwu7JjEbIZt1Cm4LOaXWUXqsXWGhGHkzFLCryOt3YyOKB
qarkGq06Ip9nwI+M1YBJ1UhgdKjDA2ph6soxCZv15amFY9UKuGCTJ5Ifn83p
JCcJzvSo1srR/7n0wmEs027q5a/D3wDi0O6NqxP03QzP5OvR4imlIE4cvkft
eNxw7tTloZ5R/jY6BM8+pKX7kKxAdahuEOEXwiK2fU5uoa2IqGoJgRDXTw2m
unJN78pNzNXHiMg/rTOOEh3Ep6wPIbtd6LOzjRJYGBGa/sO4raYH3orRtBmX
RNT3fwwmux6bpo7b52MVlnUR2yrQxUG8AklCZakqi9h2hoIcmaZjJX3j0bI3
HCwwxdb3WFjc4aVlpCEYqLBkiz4HBsNYyLGQw0G63Crc1+a51LdpkMa39YH9
sCjfHcxtqcU+k3PlWzA3rOSo6Qf44hATO2c1l7RBk6UMtp23wC76K9B2vuIM
+MeG7tcrjYhIRRf7wfzkGKFO1k6AbQQlDLRI3mDnpQlGupeHtfViRYoiw7jY
TpW7rtm5O5Ls8TETcdAZInhtEhyHpNpVo4Iguve0Ub3Q4fL/WzVL4iDiwFMi
rbEj3o4mDJOyAuk0P0hbSdAak7qJt2wI4h0iWiRTDrstIxBkgqs5VQ5N3hZr
nRLCdyC4eUOJM4WljRwS8rSG3V1W/X+5W1rv6fkDXSlkT12g1tsLscwZfbrg
GB5dcPuFCMMZRh9v8odPx/J52nQev8RqDLrJgyRoKO0wjt9GnZFpslPJz0cm
m0YfMElrw2x+yRPSSA1Em9/rwkC51b01npw0ZcSnwJHVflrdJVvXKCWtb1Es
xhKs6kcangvKZyDeaTkmzsTGSQPkMKNONqDg49ZxBg8qLgQbMGK9HdV2Xh8j
mwM8LbrAY682lwgdghvBA18Owt9lay+ctUwL7VBtrcgZHlR2VAh221Jwn5QU
b55QbyyMll1iWorYG8eAYcI1mGTjhYdkOe0X8pmL4jS76k75jFgFJC+NDw9V
6pfNeysdMR6OA3zTLTFnELddz+vd4DKALhs62X5j5i2s4FaLMFwF88cWcdkl
4NAIJfXVU12t9FM1m6rBcSktSVL2Q0EmlSuv1Fvp9DuPhJ72iqxGeExOgeqv
a4MfG9SQ+wDSNnz+yNA4tcKH9U8Vll2jf4AgBo5PNkpkMg5KXjnqwens76vL
+CbgLgU352Y0FvHV+xlG6Oa/U3JkieYHFzwL+ZVtRUjMSmBZ1AKwwjRKr3A/
Dv/99j5qlWnRPHW6ePS52IUbUMmFrp/57dZhdHS6Q+vO6N9Bl6gJKOS1ZCHF
ynSCLfkhqTfWXZU5OfybsmBrSpZyPjnN1Qhia+iVX29Cp5R0Rw1Khc4B6IEt
7Mg+ZqM1lePkplCWsBykFHGFMqMBsN63Vob3AOAzuje/hK2BJdGa764vS74C
O/ILRtiJdFIvvNRGnZyHND/k0pcrnK+VJtFNbHC1aPyXgsinDGoI+hdzGBcv
VAS8hJ39cPpuPK46MEzcw4Cfo3+UoP+X4QQkAdaIicrvEZokbB7pNQYv437I
Cs329YF0T4K+RqpYasVpZjaytzQEEZPCMZH60wWNqCXchTE13pxBBFcWGjL1
J+KymUg+R6VC5h93jr6kKoiQHTlg1euyahYdS9CI6Cd4z/O3YUOO9aDpK0Xf
FhvHi9usOpo079bCfkcHp5711eDF6DjYBpawa5iUs1oQNhLekJoB7aF+DGuy
L1EDxhyUYctZ+ThmPrJWQu4p7ws752HSewyJMZm5eUt6KuqGNSaxDKIITADY
T/Md6YjQWCBnpQGlWDbEtwA6hBMD7WwGjGYyAJSdmRw9AAZHUN35dmN0FCfU
hbDFPSfpgidp59Y0KbKYfHAp2XpGLw1IHQD18BvF6wSZVbJLrpZIv1LkkXcJ
vgcS1JQd8Sis45UTWW3biX7APvdSFxlAIGCTiPXK9QwP3izb6pwH2g+y8xWD
VzvDo1vX7fln7p4w/9etcztq1tBQP1YKX2lcogYuyksRIRYZd4mCQ4Rk0e88
wYQ6xJig2kfxug2w0Kd0UaZoCW31Bwt2xvg9KDPZOhByoi7dFRtWZ+ehtfxH
hPPrtXEubkZdeditNsmPNsHurqdkh5od2R1zBf3AObHXuTr7lIoMekjaiyr2
o+aKeSelVUlPMy5iP5z69Rij6r7Jx8Ib2REl/3ok2zVkuaWOgxSnEhkuD3Rn
xWMvlBVDbVy1e4V7/+yjtuo+Y6lB/NFxT25K/+p9r5264XuSpB9qVJEALE4N
fVYsCE4A99M/OjRIwHxwz52f/u7oCW3tgtoHOgx3Hn9QROj+QvKLW9mVeWAJ
DxD7HFM7cRxdYawATmMl+Eb3nVk4pFEyHOkbHmm2Qa28ed+JuweOSgPiU2j/
2rJHruoVbA5TG599pWFxyl80lfQeEuMyGEhzkWe1y2BHL0hF3Usn6dUmMU7F
kfbtNnjRD1EFcu3+aKwzwVv48w6e+Kk0/HnfVKk40tMfpOABUPm5s4y0fvc1
u4dLNhT/JsGzVo48hOC6OvCaCV/VYRC3NGabBk0E9KIK8V7mPg1mPNKNO2WF
SlBrVgIDAzlOGzhZb3GayHHnaezo3B0PZL+drzgSzd4AC5Xo9znzhwMjYBpI
SnyE89KK6zij2ahhqj5AeXaRLZuPz/OjE+5wY6K0aaIF7DCMtnTmiFV39u+7
NrJAhjy6kN6LuxYAhmUJn4geA16tU5GUt6C68UVLujC6ZGZsDo9LwsoG8cNV
hMkqelpIjfMcJ8l5Un6OGm7LTafznnD2cCMwkSSe2Z9MDijxJulaWPIRtYlp
HECZUXLTgbI+BFfQdtoZJnzcwKNxXhXcuN2kWFrJz2wYY4xPSgqdAaRbxjvr
IXf7x3spAJzerR10/NHWFAdZs1aC2mpBaPOCGrN9R7Xb1ELq5NMc+wQdGV2Z
lwctaTbUAQJvx+KPrVAR/cc/k69k/fc/pq+3ILLesWm3frcpnM/KNW+3vHw5
S9jWyDiTlQjZ9Lf/FklxutytNRH4T+2syDAcOX4svL94Ch07C9x4zdw5fvIT
pONSwZnJtvVzEKgwJQAr44MdmXxNjM9SmRudtQddvxz2t1N7RSQYWFXImAIf
xTKJFmq5JHQUdGifhiAwMafbFXYBf4AbQtuBGoddFYcM3AUEwMYrzlEA25sp
wLJpHW3oswlukLXXhl3GzuI9byS/p37ma2u0sdchuh+4iIaBSjIBaBeDW0s7
NVrCk8kG9bWiQ4uuqLO3f9EmT9Qeg4HSK5J+O6ruPb0xIYmUDk1b3naWxOq3
2sFljOWHUbK8v9hNHyYrSbtJQ/eT1X2s1ZJ5XVlLMzR2m1Hjo1Tcw6p/464K
LBBKLoCALyiDhyc5vXWzMxFeUyNTqLcHqQ7Xj/RlB68Fghx6203TpoC2xqcw
FD9IU88lqtQ39vyPp4sws8s0PnJPJBxh5VHIQ5GboPzBdbz+ad3sIQ1Ohqi4
U64MkI/4rqNoEbMpu8gLtXdOSeBwST7AL8pgGfVaNk/pC7oPKJJ/Pyh/jRXW
+L6s5a4cPPZc3DtvuUmhQO4QZ3JsTgJmJ1zE4DwH0bD43udjvDZXJKWbJYNH
ypEytEMCZsS/xB84AZlgQ/qR7r6y/ofVeVeffxETXPUp4WlKoTpCZVm2SUKz
TdO40HMAfPkQXpOE/fZ0EkIfyePz+sU7WiTJv7XMqiLQpJ/DSozIvUlmR00+
GoIpd8YzusbbWIxJ6bHh/BxpWvGwmbUGOd4abXBWL/XPCPbto2IL5Eepf8wC
jTdReJMobAiQghP8tPiL8cioaWWK1rUaf6FRv66zZHBCOa4sDRd9r+hGHls2
gg+J8DfuJDuqjbG7McTNIcjfzcB9kK05U58J9N1ceqxL/yF7aHliYzyqND1Z
Ax6+gHtPF4QBXkw300SoM+XXMOqwjw1OIl8gtzAjgMESjnlSzotPQndHkJAB
T/iClGi+Z5FKnG9Vj9I0oEA19jtmxE+H09Wl/GI0I08gQbwHg82y44DQAUaW
/tBgGoJTS6rW4Tf164S2V4qATqhye4vlXyGvZhzDGBxIVP9/Xaacls/9HFje
fI6/hUzIHjhP++BdPVs9yGKFagq5Wocgp7fMCUU/Ys3kSQY4NbSbomumV6d+
tufvtY1526GPDv5R6MeXe+L5uKH+4MhU/Tp4b74YqUcyIze9dpEN9nSKkH8U
CJ+bnSp8cJJZLY2/ojBkPO3uidZiu7SLQCQ6FyNS9E3wfqTuCekXU6hRT02A
UatpQWKy0Om8AHi9uHN1xUl/zgJCKKNqBuke1Y0bdiBqgmbE/TEj1mMf6AzA
X6qEXrDb/qR7NzHbq2y+wLfOF6Lv5K2C31zFENOy2axIiDRcnhkY1EdB1lQs
YTlC0srJj0W7YA9aytqlz50t5snTtVlmFfJ/eZePPCUIBPIVtdbJ5TF57bnn
KUk6pypoTgum9rT736pFWcOpyD2hNb5HotVFwCBPl50Ff5jhaiPRwLv4inCu
QeYciIK69Pj481uw8snoogtYiK1cUb6nAfUT/ZNTanN9ac4tqv83X6OgyP6a
670nTN0G82VJT/NQEXQxMLQ7EqPRnrf9VOimMTmMPOTn5ALpTd3DnefsG58l
kZmlflzozJ0fcOMbUACkxz69Ct/eFplKm+bFNiEjCeAl/MM/Y7c6I3U4fv5u
/2QYUgBKgGtIhoynR3DYKfcgvBiqBb4U7BJ8euQYCaMKF2XJ4taq/6rVz696
pZ+80QwRsDGkelPD+wzmOn3EJM+ef4wdl03L8jUrOAHWHKe4Ix8uDVXEOLJk
N2hoCGMQzYhWIvVY1CpVWL2RGx+RRv4TPPX1ZDGn0u0U+FbzmMbuM2jdC0nd
/VaGHNIaer6P03HuXYcFR05Z+fPwPNhcQhGU7SiqHlYIAxgpMjQxp6SE3HkM
IsA+Jg4bSvlokdtlwcv0yQbDxawMEMb0pQ0t+FIst5hROCRelSwCfiXj9PMd
UVdUVtSnnDkPrrLLLXTmDVn6vKljNxhkHLGxaWY8e97wls+mgL2jtf1RHod/
uvlYWxKm+UdarExy/lQ4mPZLU/Mg+5fTuhnpiwI5jL4JG8kAkTk0y0AYjeKm
ABkMnERmGqkb9SHj5AERCI7SSTnWReoENhqjWAsocUMmWpWVUmxlvsS4UZhu
ViEttf3SoeezrxIRhU9+lYd6MHOC6xzom2BXTMC6UK1rmSGog5r1jpx0rTuf
WdEhc5APuv2idpXuWpQ/UuPio+bXedQM4M9tRHi6Ut7QIHyWIURUvbwEwcLd
Wa7v01viqzL3+ynmo9eNa8a/f8/3FSCTXFLl4fW/cigIYa9fwB4gbwzU+Ngk
r6eS/NEKo7C5w21oOGEBrf4h/ZJPI79FlLjI+oCEz63RKn5MXDWfUn5O0uhD
0Cs76owHw1cV30ig5X7RhI2A2TTh9qROH2vUWwo4rksf2jJlDqkIMyfG2OjC
eLGt38F1UHJ1amZ1ZvJto7MNDZk7q1K23z3rCr6Pmc6gyaq8F7Fdn64wSZoi
8AQ51AEqH6LFcDeCcdFY8WUwGpAz6Mm2em2J9x0c7SPoaoeAv1PQ81yglEd7
rz25+B/llQOImqo0haWCbg0dbJyhOj/K6qqxR25YHje0etirOVmpMZn1ypW1
mYpGqDRMwwlBRUtOyNN45/bq6eBOCuz9FXs+ru4K8A0sHJhiMAh0s7fPYsZy
VcW/NSB3rYBluxnRwiRrHLHqs/xGkKKWKLzJqXVPgXmQwrRRJLl1xApi+6Bp
I0gWnJsehQJLd40DSY7eiXtlw2nszCqeie2vqi5RaQzAf9DY9aFcZGTLcIMK
Vv/xxWVFpYQPVSba2OuRlrEFvPGM03t58WOor2L+ZlC4pzhCXorcvuLWd21k
3MPe6hF7PsZuIQTRLC+91MxTRVJzrhSiQP1oXkDhdherxkk3QnyUD8Jswu+1
0cZFe/FNR2jqgFFNeVppu59p+QKS3t4mK+mF/IwuDD4Txbjyk3ZpHmlI6dqK
xzQuhUJZZUH1QCGaThs7V9rrCduX6qDW4tYufgK1kq+Y3DuGFc/NZaZ4shMt
syS6i3MgXxHCdZ+V1Cb8YFkQgIWnWjbQ7XjqebGpbIRwb5w1a4jhBCVwhqKf
oOFkpqO5o9lHptzlGLi2fftMtftQ225bkFspale9uGj4+EMiCcfYxdTjQ+8t
1WoJKwLSxA4FZKrcvtUFiUu2wjmqVVsOPn/6EzJ7TU7Ntg8gY9S0NTgIEciN
P4odEOC6XUb0Zi7QACympiM4WjqJ+Q169epvd3MZLoyxyfB9xZveUdqQr6vP
etu464LH4+Tq8X25phCYMyoaJ37+Xl/IuR+hKijOy43xx4IZOomeG9Prchty
TU6v1QymPRi9fXxt6vtlVqbt7SSlQE4ynNkrBSFTRCzT4b9gPbr80Yoi/ety
Hex6dV7rSawAIGy8ne4zju0n4YVBeXG1BWNbaI5Ta0XtEr6YLLdTZ1S2SDGS
Y1N/q1wZW+liaJMb2ycZEZO/j4/BYGpDzYO/Bskrak0dLAWVo+j0tDsAEjJS
zyLMPEmGDLlnaCi7iED45HhbEPoWbpSJw7nQ1ayWnOPOSpP5HiuDo6qn3E2R
wbixJSVu9isf0+KXqmB2mK8FLf+S+WkBq0xMb/RC4RtoQ5pOyAFsY5rHCpWz
nu2ik5LFcJB7OjRaIUeEtYQh+oaVca1QIE7XSpbsiv1NwLn09Chb9+wea+y+
Vsw5qz8fjQBqIjBIZFO1N5XcVYoMx9X1C5W2ijtPgvl7c6fUdcMj283vE837
UUPuwJ5dAmq5TUltqZedXVmqrfOSWw1R2OYC3WXN9HwdowbGYeDHSTMpi6ed
6vo06u2bDewUTfVB1Z7j8/aKASx5+9dosyd7/0anrHvzAIxZ+dM1BVVALZ9s
AEo0fAL5SVB/22lzqWZf/KJdsVvlkcHTPaaWNL265E7U0Nn+HBmKOfpBTOYY
20sm4HafBwjTARK1SdvOLcT8CYm7HSR37mtEoKq1Ve9D0Z77AyIKUqSdzVnh
lc8OBd8Q64DQfX+mCeG1cFm+s26Dxx6WQc7InpClIa9pimtR0ncRVNEREwX9
i4P094Au918R90DKb4H3GrIa6oK4DQYysexjnwShLEFZG3+j+2LNQWfAujQS
kvBf0utNcLRI9/3XpBnWEgjfKPZ6ryrUcJrdx7o1bgwulvQfp/m98H5KjiIE
1bI2bizV0FZczTUe0QlX/t15H6SlnNMTSXVDczgrX6Cur/6GUNycWQba6/x9
YXYTakmTPPNti86kIcwSpkc5Zlzr8UpZw6Wr0U9YtoS/CNIXjjHlzONc5g+k
tcZ5ztr/heEQF8wfhsF6QkmY6hr7ZzXIX0kYcrSxNWs1t2TJotm5Q3fzBy7o
0k1LeXSUka9xKcL/SKEC/gK/sfIhoHbvWGVfBqJdkkdPXSq1tQ4bPfCQDo/U
ighDxf1QSYCU1628Tpr+p9VoyJ9feZEAQ8WnKyiEWLgMHyDjIeYEcxfxz8v6
4cmUzPNkQor3Tp+NTFtPEJVg8BWL2yklmLNYGup01qcxqw2S/GzwHJe22wa+
e4kzivnnaKN/hpFnU3DlcUrxRtSWqOh6OM3au0WKxr6HxHKZlikvQMNuvt9N
nw1BzAg8F+zRyYv57eDQMX3OpdsXI+F+6MH1EdzW6I/pAUu4Wg2y5bhHxAL2
8szkRyeInZxf7GAb6jUT7a+HcCdgE7bPHNA74uxplPuSd9xcpkt236ri1PPn
qFrXiCdR3oxq9jTUFaiycn9fAHuAkRc+2+plrQngWib/LfrWYutBcxpwxaVu
ms1Vhtn5d5WiAbAbHZZy+2pgyje4k9s5OnvAnoX6IWxMQpqSK/xsSapZfEc6
4NDj/laGUf/x/dTis1mR2E4MyUqYP1XcjwNbFU8uLUfqyRALlcmuwpiDUQU7
r3FpAac4UJgjbeXsQJ7jEIuyyjqhR+UjaAVUymkNnEFQzOL+A3+jGfEiT66a
x+eVCjmORTspgepkpoTvQDoftOoHVV1hthufOlPchlihzt6F9eowXtNBopTL
BBxafDYXgQ/BSyp0p1AVckEZVBm1vkwc1cCHv1XpzlWaXpggZJgylhhItkYK
+OLf8PC8pO8IGRFqAcCuotuKyTdo1ZRjQrCPjQ3tzo55fpvonHxu/do61MtO
b9KpeMva/q43iiIykW1xiA1be5MqRFwSEJGQEQIgMDLAAuN2WJCOIGuzulDQ
t756aeQPMQR2e2cdM5ZfLDaFzwaaPozCDjs9OYP8SNSN4UGTPj0IjRg+i5UZ
dXVypnEobFSd3xlGTYwrBSG0aB53l7nKDJnwRR6IY4TVEarQdx/+IkmvTgTt
lTPPeVq6v04rdT0aStOLdcHfuHhfRJN7fp8qHUyA0RkMAKI2EfgcSalHPEgg
z3N8pzPaYCLDuFqk7yZUIUZpLb/l+J+q/RdBI3O4sJupL9NWQw7wGqkJFpB5
LtdiASsyaQrGxN7FV8Iqitgy5GxNGqHs+sMvPdrhDQ/o2SsxNRrCV33uOg/S
RGnV+kktkdJgcF4NXITSHn1pL/iFa+m42rZFuryDbnO63QaCWRsWHaW9pBMk
kndpu4/K33zDAEvNkUqADKfuj0jDBiYFtW3a6FZf44bQNtAjuqJ72XimH1p7
io7oArcLFWVd3R4XszkUghVCzf4Zn1HhXwUHv6Tatw3LR6hVJisTyjSL+VDl
gWRO9oJwWobWWnXEPUxcc6eeeRdqweb51x3PwD+/y4eZ803qif4XRnmvLANQ
S1GRFDJ9jl8nsyycBayEyOsdZjLRZfywQ3RLAC6mQP6lpBUbwmyWQ4qYi06Y
j/DXTEI0Q+sgJZbJhWhXdF5Ns1m3n1Wf/nOXzbXWa7Icp0vyd6eiq1/9xrtM
814gzPlIlGuHTvzhWzfLfyHNXY6FT6zjWR8sySdoFqIRrVJxLpnp9ynegc3P
XYIssq+tPg238hHLJQJpgWDA+qmrxxGlq/P6+VLZtp5uNN1NKMnc34zkcPy+
5xwValFn7CB5C/LwPsD49jeRn5F6j3VP4GoDrfl/3SGleANEIGcp+idJ/boY
Dk1YhlxDtgUsBHUN093VFvDtH6mJrpotCPhLDXnGc9e0kef9jskilplXly3S
tsX/eCNxp+9wWW0Dy6b+lOYk9YPNOWLnD9DsqcwZvU8pbLzVvp4nmDFqFa+R
1o1Px9bMeYC5nOdiLD1j551M9Efmuq2Mx9DyoaDXaIzb4b1C/aqdZNtVdn/j
47lTtX6Waz7LUEr6NJqqLkKJu4yh7F8/u8DWM9nAg3UgVbI6+xVFrOMUgsH5
RFRw/yMGLzM48dBAlrZx4KMsxmbBsTfyovIzJebSjTZQpELfo/adQYEegp7j
NyMJITBPeVcFjAPUJbpZ8vN/JD5Yvoi9GYDHsyVYwV6oamaWG5AnUWy/pt8I
2hKsPfJEFMwTFo2QYkfcxYN+1dZ0bVDSR0NrBK77Twsbc5jryE47kAVCcSOJ
hcSRCu+uYkM51gzYrbMQRI8b8KrT1dp/h7ovm0ONSMSvi1rv6UelEENXC/n8
L2R7En4hLhAU2ASH0kjCKvHE6SyjfyoHGcdZO6c0nekFT0v9h0jqro4qcqv/
g+dF09WSUD2JGEQbqjph/Ts1aC25alpH2ByQQaVIwomn7VpeaQd1Mca8ffOx
xg0RnSOCmngjMyVEr91X041whi5qo/HEGS8JYGY5GSq2w8VbX7SgJ4hplhg/
oj5noUR/SLCzLF3HBLwroSFt0CVFQf0jgC1b24S3SSuuuD4gnY0qfEVeDU41
+xx3xtoFeYscp2IBXB27scoatHAimV5VimlVl/4FK3ofklWCIs4+b7h3FmB7
IR/CFkFi6kIrLRnMoTMgtA6jTuXKZThY8AOexqx6f+c0wNeP3PwWbVtWGpKv
leJkOvmoCl5jlzAMRJpgqhPHUQG4xmnDmdBuAcCz0xIoyxhET2VJrX8y1os7
ODPhOUliwFblu8mONfPP+TGXhPSCzAYo4bAt0hBCHFtrpL9GSL30VPjGof+1
+ueGQ9uXfM7wel0dC2Jz8NVKiY9dLEte/UW2hfqOt18daB/gct+w4JwEc8R/
xOAzL2isIeTEP3WLS3vsZaZslbHNGaThWHUFAAwB9fCEGscu2twRZaKRwuPf
dYfiOBjUi0HVbtcEFisDgN74TEnr9H2ndci5Yu1qSBnUxHoAfXj0lPGjHGZi
ypa5B1jLmLz0Bv2pR1gazIxAJcJgf2LjJ4ItxRCSNx4nEEDTy2Fk+Vcmu5+r
DG4KnkpNe0Gnwu+txhWmEf5qN6tX3A7f6p+XILdnFnGskOSGjiIPMY0xvEDX
0Ke5BlNe1xUtk8NDR/2LSN2V2d7608ZSl4Qac86fa8ttdY+/o1wWusFp4h72
RgLFgRO891rljy+iG28bEp2LQn+tI0lWcrCV2SQroFFM0+3S89BeN/sCVzHC
68OzXgtPD27qaqw3wJJpQ7Sn9YwY9igBnXjbJcqa3yD0viTctw7M9O8NtwBG
jMxtR8EN+hFa1dhj/xmWK9LdLKtBX0TH2lsldO7nBC9VABKUuAWX5JaJQ7Q/
E4ZEKIDQuqOoLTRRrI+gOPRFSfpotrNvbMuQ+e0XXkyDn2SYONOS1shweAAF
SWptAKBycgD6n7+DD/Vg7E91d/0IPY8vhplp5qgsPm9oRGIBCEQzbaqP1qtw
qNtKOC7Z9rkaCSpUVWi6dlYRbqQwxgyEPX7yE9bbn/dq58JKzJrN1++GHwRn
httxZnFRxUIxcjeLtF60/pdYhrLfra14zygGCfRIAkpzdpHxZXffJRtz2HcM
6zJ8XMy4bofztXwVnBBYGFHgIpwFtzBux0/rZT0rawUg+rZHmjFIU5XdE/jM
MnMH9n9riKgMoxn7ZE1XS9La8kyM5Qo8M/WxxV2QeBuzgZqKaHYIWoVrFeL5
5MhZ2NUD0sLQDwLRX5EsVElvivF09AXRKhFGXOL5LvoPwITVuIF5KvJ333Hr
eJbLwi/DfzplEFRypcRzq9O6pnNzzrG/tDnhD5hdmPItYJQuNEbdXak0YyKY
712Z5dyx0+M7EcfQP6IMp1QzBMQ3v9YuaUvw+RsNR6lXB/HRwybuQ7fNmm4z
PJheWdMVPde/V0gPgPFQVRD9Ser5jsyOOL5zadewld2Uoqxyy/Zfza0hvp3P
9cqTxDIsegLz3wufA5ikTPCeuTO2H+OGjY5TEmef9cjAw0imAi0KjK6IkgDo
VMzJcnW6/PyhJkvXFrJgyGu5Y6C9/s5XjA1GedQE4nWlBbkfArDqvq96O/Cx
wzVIdPw2moIJBxma6G0poEz6vsDDYXhtdw+2M981uRjZEvQy3feemnGSXY/t
ADaJMvs58OrAjuH93m3oCs9xnmGdBWvaKKPZVqqR0tESXcdmDdHnLwnpxirP
GUKwmi2e3ZIv7FEHaD/YSB7vEs/qVwOIlZ4mod2qm0nwXcOXKpGq5cADrRZ6
+8K8xn5GyMzSk2BsamnC79JzJ5qd4lM0yo3Zq27/xBlzoO2DSWDCoRsO1EnW
9N+rcvDS2A5C3ufBNEcfUmfgfnkSye1gfw19zUkdrZ00a2gJ39NUVedp4jyz
8YqF89FOViejfR+i/CQZO7PNbes2el/q9Mn7y2i40ml7m9X+O7PPsHjckcWa
6YBOJk9Hr6pbrRgtUrIB7V/NZPuHqsJYE5ykIevWu65KTsBBhyisWzuwQ3IB
EY3Nc7TmeZKQSRNPMnSTz09/AB+6eu/5gSePYw3KvcW3xbFLZTt/r8oMzSH0
mw3MBiOxDBDT/s4fQVXMD8OPPFvRCWJ+aB3bQT/qFmbXd49ri/i/CcAXtuH2
5ZVo/xNbp/E9ILQgERFo5ebjPSGPtS0fr1oCd1TAXYnxREaEqow4Gp2aicjb
gqBmL59QIPsyYgCnJhZm+cubqSQXUmNkZunHBtGE5vob6MwCIkY0Iogb8SRf
WJYhyJVwBSgiB+0Jr8LhfVyu52IKWSsXOX2gxYBzF2EKgFzHH9LZQge/cvam
lnu+YQLk8Z8FZ4NI6/U8WAs90lfNdL3cuDiHbyubBXHZk0YdmaXMN8hKyVrz
9Glx+CaMQHb2Me2w4rVI/r/mnKdFUhZiWO+bM0lHsGDPu035hWpN0r4mS2XA
uNDCUDxW6ysszYjKie+SJip+MQeuBYYdzY5svzqA+tYLNLSUQHFe6D0s6LEQ
PBfl9rkTcRzg0dGuJdqCTrGAjLs+gFVI0rCBH+H5d+KpZniuyk+ZhJI8BqUS
/B9Mi4PHqEOcnavxB4ffEE8hSXBWJD9afnNx+kSWV+Dg96YyWzBO4wI6MLzK
F/FD0XhNGqYXqNm6oDdNHl558vLhkGdNkmMTP7QXUuHx4whp0L6ecVsj0Ih2
GqJtooX33UfJ2EN8eeXeqjF49psVvklGTrJFyejVxKll0aOm7qUeTTZBqIu+
lLFTlRA5qfohpXytmXz9cJcBNG2L39ymEzphNrJy+kn2WXVLD9xb0oy/Xjqg
o3rjrAMwmwAm4kQL42sNvAHnG8ftRVNZ2HxM7jwOIGk/zxmEv4KgSuiGngA6
3E0J7LskdrfRg6XZLqR4ET6sNBNdW4Vph3tsWS/Ds1cmVo/rS7IlvhcQK/dn
7qsOCx3GHMHvCzz60+0ItP54ivcH/4Q1kkCdy7Txb8NMo0CPm5BB3nPpdwGL
vXjlTSYw8L7CV4XIG9TUDc5rm5ZF+PKn0ryv1eKkj8WgYxtfmBqMhBR042jm
4HEZhBHzWMGWFtkPwz5KjLrPyQekUuZLAQ6AYUd9U69HBdEfsvxSDfAl6QqS
SA4MbMJ3rNnbew6LzoNQ2AhnDy3BmCTXy6nLoGl0bIJnNzSj/VjCi5chi8kG
gt2sr2cdOW7kITOv/v6SH/vZLId1EmTjd4NHJm9KHPaglYIOCFAJvMslRLp1
pMKnHQ+tWcvioh9nslyuDZ418gX97rRGDq6+NlgmGRD+RES6PcO7iK+cNKnW
KkuM7FfnnMi4Ae5tg8FWd79JxzbwG5POsjbsVWO2uxSUNV49ZP2dVStbYH3W
94pmtkQKyvq9YgP7vJM+ZZxWl3tls08qnPVgNd7mJJXHEs7+hoe1O46mHstD
MQGYtEQacYAXvnsjckrW8cvKeEfhZ2aeVL2G/anTcfA6hkowvLbUEY8AdN3x
Xa7BRCggbj9yKPErHBgpDjgPlDbFfU4n+KEqOWSPaxoSMnIMyWDMsFYZadsp
bAIurJ4Wu0jeyfycwdWFte7Bf+/OonPXbES7Rsi8ibQzeeX6vFIKKc8iK3yP
zKZOKCTbQM9Vv0arviCNBT+2xQt87dzr2KfbZTm0QxULc0FeyLiGYR3bpW9y
ZnD+uhJW82ltBZ/kiu00gzhRqlN08pO/Eq6jSI1h/SZKvP3ey7ZPDUA+ezIG
XzF4IJBZLJSpZfq5Zr4ltK4R7EEk6XK4/6OXnVFnGQGkJN09mtWz08/xga+9
rPK1pauWq0tMuQqUSoY46vjX58xZuuZ+kfDOB+NdM3kmtxAA20zTWOfFFOTR
hOEpE2Ub4oFhcDnRgWkQUC6HqbhrG2TrTlBCuBrfxlLV4n/8KRdBD2llsuJP
8KY4/4WCDzNUe63dHEU0OTSTh9noR7a+FloVSKPP8PzWy9n7LPIR4IZGeSfr
X09oXQjU93J5QsggPRPS+87w9/B3N342daoNIU3Wof4oDSrQ279wFIhWF8OJ
iMRdGcU+3xRuzt2sm5KVnmfrOB0xfMEidaDqNhR0LwJzJuAsughP57/SqQvY
KyVRPtoARR9WIZugi3WpfWkEEvm/PbKgdkozZs9tC8jrhBbrJJxfe3Xn0Qcr
XbXoRwXJKlH0PxNnqcAPepWjgsTH6obvluLUgF/5QPzWle6+plLq8Dv9jSSB
fMxN0z6fi45Rou4tM4w10+QmPewCJVsFpTs/T9Um9Du8AfOSLTt8Qthwof4L
Z65RDHhXhCPP9cZY1Yb3+83/z29YN/5BC6nCON/oIeL5lY1t+C57Tct5jgpj
Ful5jL7FgRAFub9qCzQRp7Ib4lny8USW/Yltq3er07TInRo0v/w57KSkFply
sJaUrnCvtnKihHIS9nTF+Y3Jxrn568p7vcpA+7ZWYCq+Hk7E+7RqE6v5YU6/
bHRSscCrqv7qloRtOnwb03Gv8AkJNVmXy767Y1ydGTSzrabC9mMlZIFTL+vn
s9KMbMMhcXPUxUlldXKMUsVmJ/vPs0kKCz5yYb5Gnk9NkntxpIduK+8VcS5r
gr6WvDp8QLnoyaHzAkxKtg1i9KfhNULAizMCIdlMHmXeHK1yvAW+fknKqq4y
BnFZsIOMZhGHp/xzQi9DBxliI4Lv2SEt9rU0MTswpoMr77LfvFXXlECTJDEp
fJv5WIOV6Uk+6w1yUZD5vBiAKjD0NhjlPlR9Xgtjt1SqIStwRGed//tU5UFC
g8pM1BN5fVkLBsC9N/lkod5Ij3tUeRur+k8AoEDVxgpYsftWuUpMXX5sO7+w
NX6haM6Z5EwFEWnEHElswM+Db/fg7gM1wx1nmxwC759kJNif592Gh82m5EPi
fqSVVy4LLVrt/XlZ1S7O0T1HAPYmanwniWrlvMm3uqHbxWyxzr/iDo3zRntD
BWOabvFWHcIPhW7QZuqOQb3eyHN5zuRc5gCcr+0Fy2m52KUHl0SwlXbXY0pc
PReqiWTyUrn57yWX7vDk8bUE4vDJQZ1pBl7y8aLnI9M0ai5B0CZT9x0omeOe
aVUBFvzWW/KNrzOjubFk7E2SqBuzOjyiuJqWlh4O4b5Kv4KZp7LfHhfpnUFV
GPbIe85XbWOwLyqUZmPtRcMQfiRWo9IWY6sbMBkQYEg/BCSb9Wmd6kLDVTtj
wZ6dVkszQqpYbH2U+R7HrLxh9aJqYvJyDwsjm4bcI/ZlefNcG4EnpZudwUpT
EYFv6xySDSV3Lm8zGikFacqp5+Dc7N7fRoEloXXkYHIpoG0d8NAqTwkt+u3k
4VO2iBE/w5nUJxaSMGoEP/gIXxWpae2nvgdzz9YkZDGhzzlArsGpmCcMtgVx
3SckoVvBu9pqaPsY4vDWJuY8X472jJKuYnUW3ITI9Jzt50BJ65dHUtjC1yyc
rlmIC8+VPVF2Rhg9CuqJxDeBIWHYgeAmiD6xm2UBYpUSUf7+iLHsWwwqk4a6
4QgPiBJotdlLMyp0uor7vv+R+ewY3vkcOspH1Ew4cbFLZ19guvYm/sm260eI
F6/P/TZOybxoQLfa9fL3jFurQgZdGeWwfkbzqL6o0S3RnQ2cdiWACkX1BozE
mcuY6smGUAKH8A9O/lFVc5jf3pGkm2+0fHM3ebjmTwRmg2/L/JifxsR1vIIw
pB4etKtkbRmPpznPkVXcJgn/G3AF1k+os+Giscwrw9lqo/xpBzT/Surdguu5
YyW6rmrpFWJghYOHgDBDVCgohau9h1p5Utbq3wUgcuEwDamtqSWDhhAz/+Hq
66QHv6eyUxWssEac1haFvZplU9kFw6qgn1OBNseoF+Xe5+StBD0GSZP9A2Fz
0cht3mLdcC1Yg7UHiuO7GI8kN9O1C8quw7uB6sjS4gDorCdbSI1prvSNFIMe
r4iZT9yPcVtyBH+k6xBPeHwEH8Rghldpjkjkj5N4jHSBLypfrBI2+QE3VrkL
4sE+wNJvSNhHNEF4/j7Cgm94N5CvXEvkOINlLAbnym+AAoaCAGgAl/bbk0Cu
CWN0VUFkG1yzKmLAm7YJ56Og9GZPdBQdu/+m7o8NPX7TSutJfpAoCZT8tke9
EXT9AK0wiw6zE14hL4J7d5XQqN9EL+7rs33iquiwTIXNYBcPehhD8Tul7Wai
EB1YIaK8zVL/a26LVG8MQzEuj44vKgx9Eg42VzMRZ6HBoa9hzeQFIVW4Pnnn
xJiyV8azGkyJtAtfgQSy50/mACdvILD/0uK28Pi58rOJLsBkl1uSkcMSB/MG
0SyE6+3KbTEo9fI4QTMWkWF7i6+w1IpzDVale6mFsO+pwBIqkMNaS3uxqlYU
6z03mdNslWagq3MrC7eS5q2853I9OHAfTEHvazKkMSy62kPSB3IVaQQ3eIgz
KDBErCru60bX+sgNsUMSO705kinji3eb0mMzlO08FvTF8quB90988q9siYpF
XScxUElzNT7A26lYRYjPsktYA46EKipZwxqTgetM/2mmd3Wc9lvdkz4QSsF+
N0p6NQH7hmIY9RNtdoeHff20AAiR4pff2vJAEezLKxT6UvpUvPEf/aJMLmxI
AqXej14EDwtppbEA4s3NYOiux5JbWrpis6w7egVbIhFEw9mHP9fxylsZ6SqB
eWh6dfw3wbCsA0rz59Q3+2GK5UK1qmkPl0hZFToDqo6MLnTWhEoACpY3pvw5
WRpoXTO2qV8IwNWTQAt9wW6EmI0OBB1BwrORmiPp4MRF/Ji4F1Fax6vdlxPT
h2cfijt4w4PN2cG1/WoKVSXM26aoIj3oYG+93DmGijVeya/VAeg/FBJV/uEh
mgmJ7PQf4KiOdkl0wNNsFLclh0QCjUgNltdocKpbw2B0gRnSxW6Pt7k4v7HW
/HBV6buwnsU5ZkLpwBQtEdzHbd+obxeGYTjgw7rdPUvETdTAU7X/FhBtQM5L
3UwjqOwxWLiwd2L7EqwK5CtfJ3RdatRF5BkwmztNfTDYhZpkPK2l2b0EZoaf
tETroZM9bxJsSX7wIQd4P938Xz4u2VHm3CEOLwfWDVk2rBXm2/Kw0redVGL+
fiDCw4VjvlWTtcMgKwkRNWpIBBItZ57ivAexH3kitHHJyxDD96VJ8vJaJJF7
p2X0fK8KtYHXijPcnIatdyfTMj2tQeklU6FPgzv66aO+Q2YjJdYR0/bJyT0m
mFZqEqd6GCTgKfv8GIgB+sfYA9u+yHkAdbLzzRk7DZwMCJIyQu8l5rLwJUYL
3yc7Di6829dqclML/+VKLC+4hUzNoAUtToAL3R1uK/WW+i3Y9mXO1VxZFdby
5/u//dJzGULbN23lXzgwT4u5UgQwhtRMKnCzdLyhj+se1yw4gDinDUxOV8oB
2iHVcx4FebM83g//h7V0jgDlwHhX7gpJ6Ug73G/HpD5xNNN68ekKp3UbTS06
Kjp3JsXcskbqDjyZFxf4l+l1gutXPXLfNp8i3q2AvJO+1vn0LhZc0hr2BfQS
RNrLrsKOpoEg5rCD5i0KZCzrH0YyboUPwP3dsapdAhkMwCDESERMbv01Zrzk
M6ir7ow/ir7Wl+Tbn483zqYpQvBFQFtX2gb/9UPIIfj/tHtdO3D0FSoYniHK
mL16ViMY5QKIHQrB4vy0sUH2lvBSFgsC+5MQOPQpcht3Kgpg3Vq27z9l4cXZ
FIT8CB7oACE46yiNYTosVz6PUa2uuBb1LWUJpqyGcxJJec7IS+dc+FRMZpUf
DChxvfQ2cxAelwk4Gb1z/ItFXw+ubuZQOiy18MWZ+Tl+AHIF7TYxDpwQBIw2
4zoLMsmKCuXCY/ADGneayf5UJXxIH3E6wjwFTWFvnK55JqERuV/hnm148/jo
95F7iLXMfVPCAhPETqRWOEPB1lYkBTfrlW6lSDPAvNlWDOJDXD1uC/+Zjukf
Q68M3tvJ5X6LL9vo9rFWmVKJN9XWm7s2vpHzCHcfFVq/NPouXP7kshpSLTtG
dk+xcaMFxQKrU6VJecLfPvzVJ41nTRNVV6uofhpJ+oTA9IW4OzAja5HWodBT
QyOqN/UKKZTKemYOl8KO7XaasxAyXfzIXikbw51yTiiUjayZpO/Z/eA6ceRL
IWBuKLKHNVsBILCJ//8B+h39YgMaSxLKiZE0zkL+ihTJhWMOpHAB69gtFQJK
lAHYa3TYQDuscWMCUQVqPnrnYGln+y1IlC+d3yFX0nCKY2ZFy1OIvFZ6Gl4o
MOZyswklOzrl+f3Kd8wtUp3G86HiQIP2JzHC3SCEqrseFT4rZ6SOoqBOPIQH
XfIDVcCwWSMtTA6YF26KZrDHr1Cz94hXxDnUgs4S4eslaUyflzfHlOfp3QTF
983DMQXSZnzYkb8KMekwsYqY22PaUqCI5i+W8uR5GNJCvrp74ucj6C+4EoVv
Icji7k9Gjx2+KVP1ssfZ5n9NZKEpQFZM44TYAoMrqlwgonvmgFp2vEYZW8Zd
iAswSJTMZmVAS5pw9hH4HfUDm3lYcQ7+R/eTqMn5xA5nmRHz9RtHXExD190m
3fSppB1kX4ef8q4BMy2DzrrM1UNeGKisjKK2KKsrbRFJXSrnn30jVdnUe9e7
g19MZbELtSoGG34PZ3Uvyx2XekRinarAlYTeXaR26zQ4V1MDCHHhRPyHWGGt
CttGVdKA3+PpxOtjS4vX5NYJGslKavx0zPdP8PYsL7I+eVD6sc7sROFNvVRW
BIzhRYW21SDYetU/wDncW/0Ebebc6exhwEiZ6aVz9yxUxrwq5Z6XtwmfnyLU
fCMGwVaWH7aMZz7HqZcEPg6RDyuBMwWvPL0LXjrl7orb62o0a6kD1t94cnUr
lp9CwIBQ/h1WppD2O16WlhsnvC7WTZ7IyuzttebYuIDIpRANSwqKoJcLRGbh
WKO3wspNItnFZrYrrW9bl+TQDFrdM69FjSIlcsAP7o0bdPQmmuAlETvu50vO
gV2uYpii4iIsBWWZY40otHvzF6/Y1B0XCOuT0CH7n4b/rZqEGmec2YMkppFl
jHpq1n5Ey4LfnDp1t3VTG+dBJ+iu8H3SUhFBe0k1xZ1i92KcslnUVUOGgB8f
sWCYB6BrqG6y06HkbP3OrSQQYnBVQaXK0/cX5l4lglYTMZHCGJ8sCyqqIO99
owr9pdecRxCpXQo2OKva7ZkapjjNZYY+TgAorDL+Gl8NF/4SCFsFm7iapiW4
HyQ1L24vX3CDvaVXGPtBKWo6iGaPhbSSjnRDb02xA4Uhg1a89dECDyl7mQVr
7e1vQBztZJxfDOUoq8XupozAzZ6yrYkH3X57u7LEbHQhuywcXl1b7lDs7dt6
eEXtfYUM126asAUBXbP1K4UXBONUTtk7I56pDW0LJ3GttcwwvpX2ur6w06Ta
ZN38aQuu0C+vvpmrFSbGJSHQUG0xCnPXgCuVXxOA448KtKFflSvRZBJ51NdX
abdKgxUc3dgGaX2kfJNxsQFRpvprTg7t1sLzdZjayk2mrplctaIBTwkWSbqz
nEM2RCmWZo79yfnoPCGExtBteEHEdrwiB6+zSjQ+kJQpsTyZdFNJfZufCzFS
dXwlPr3Rt6diwxtAlMRbnyx8lLhMSRnIbDC0Hn5BL3LdfyeLyx/9HbTmbDYs
2SIoHewjp4OJcQsXO0xtwFroaTYKJx6EU/4/gJG5UyuZoDupfdtdKFjGfLkD
acHpbnVOBjmPg0UTB1yqo5ZW6YxEqRxYppWlZd9mgtKdck1RELlRsHryvS//
0dqiZOAQuDWl5tLpcCW6tqCoem7AVMD6ZivBU2O3zN0i0Ayi3QKsdx2++Vu9
lTWX0Q60eoWQLEo4SIXLHTHG0b2XMU1qZrLSzySEpUEtLFpkFawadc2yXDGp
FRm2W0IZN/PzjFNzPKUd3dM9ciwlpvCHKsUJha5wweQ8fCtpMM6nDapxnjOe
7eXEwIH3sVv/p1OXAP7o+PRFK4tjul7s1UhBTBMcOx/TJzwSCDgYLn9NN4Ec
tD18Gxjuin6BwwlaLcSwf2K4+qGV8vvKzwMBTOPopTzPtkbBryR/GyJrhUQh
Ynm4Td0XhMUuRtJw7LxkQFPOTrqlIMa+4PrphP63FeGi73mnkW22AdeME5nO
EjGFNpC33YIgI+udQBzHDZULnig73Ge+1DbXr0rzfZ2h+W67f7sXuAhAjR2P
LHTvC8NhJTSHJTIclAZQ8bzrSJRzsIE4hHnnZqNUvGSnpJ7kFvcVKjRTgUSt
KhcxkG0PhMrlYmQMQTnwBjcPGGsNv5a9kE7s9YhEZtpu9hX0HjEG+ehdI1eR
o8T/TIvI7iGVOdkhPWnlWgxfI3+sOZ+ysgLXhN6eWspCbvn6Jd0gEIYc4TBe
tCNI7/BcOl8udulWmjhUNC2u90gw7+bKRknR8fQNRWXsCVOMzLQT4XG658jn
7+b1r5kNZGHsWYboStLxYWIe2/VolwjjMKuOnaEOvnOnfUCi1VmOHYq37dNQ
AuMXD+6YshzxxANyHF+pWHXOJ+OGHevz64SQ3XA7ghESLgF7e+prSVKDPPku
fNAz5OKscaiTdP9Melidrg6BEILJyUvAs28gqQErq+bGYNprmNZtnbQRKcsl
8Zjb9OZ7IDOmS5KXiDzPZnzGjKgt9yFTt5hK9im1Gnegc8xapzYnu5uv0sGp
a0Eo7JX8x43H1iUjyBYEBNJ4AiW8H1XT38hP2BG8mmcEfBh+WjxAKzZ0gh0H
24HFkEInNf4rnH43/pXUaHyVvX5jxAb+Nmh0A0+jjDtgXLRv0ySG3WTxgEHA
FG1o/VjlAczPeIj66pbXWjrPeKhAovkxZT2ZRdcXUVU7jsxQHQMDVedV8uPX
JXvbd0OsjWuq8IctYr3Qhb2NGxhzcNT1lFsxq7boFUojMSnyNZYufsLhSgze
1MdRNRH3LLQkC5/ok0GVzTlucFWbpkD+LlEPLB3FCOaX2bVFNxnwObThhFWq
VXxi6ZZKa7M2BqsTwqMa6c91IEBsne2n7hWENtBRnbAwDN+L2obIfk3JxX7u
9i6elGSxLVMV8XMv1a4oxy5Wpf4L7MqwBKtfiii4QEenFPh5DueJnxmn7s4A
gCAstiyonWihiVJEIn0nZ6Vi7xqOF65UBCArokozRsyp47VvdOrgF9i1PtX8
JlDp05CJSuwdypfEjJFJHFj92JvVT8awZ7a95iks7xlkrbMtwFDoAS3XVUGv
awdijbPdQydZvBz+diEfCmnO8mHY+l0976/QINHHbuLJ1D+lIQwA1ajhWZmi
VRPA4vVuQiA5/Db5gXuDZ12DG/CgEkdeD6pkuGTZnTqNyuThb/IVHpHCDCmh
7mNPRQlXJ8omSWn9+7CFN267OSGuOTNKBzFX7OBvVaYKRCL2ey5/uDH0wtP4
jAGgczC3ie249noX9F49JumAjcDJKo/InM+44X6u/qd5MoCUwYqsfP6bPpDY
s4rCNb8E7xUdZaMfleNK4/0JJ16DG/xYYnSDmZbiHPjtmLS/rl+7yiskMuT2
Q0KWpKzBG6oJ/bw5VYbRWDab2bAqHKa/lGif4a9WhfbIOVPisBb2iQIJ4eqy
tYoWG82tGUB9RGJvbZkEXkec+NGTEbL4j+n63XZ9zFpLwTQ7OZTf2gw6bg/T
SQqaoxSWIYmWDT1yCxLEr2AbFVyklmr9ZkOWdEt0mZQc2g4RfqKXh2nSjyQM
pFYC9+4uyxaLeYLvbRfL2DoVkQDecueWP5nu1zlwVbCed765gyURZcBPoRbF
38WYfvmsaW0aIZmffr4aj5My7PGpPaeMd/7QMRSA2XPZdX0HwST7VpndSuTY
m/h8dQuaKLH4f+onBxgRJ/Qy14qORDf1gWg+G4FoVN5mmqx2tctE80g/1SZ3
vF5oecIuWQf7LXk09p8S6ce7j5Qa9SpmEvizMKST8McTLp/34l9U8+Gl4TCI
NPzwB6UrXeGUmj1hLLYvm/9uJu6+lKs8sappfjMv/nbM23EgJqXUUDWsgDOo
KkUPaiFG8YIqiVN23NwJmZZjod5jbUCUech57u+B0JTuUG9OCxep2VrnUUsg
zw5dYsfArAO31sV5z4LvVRTkYTeOkBy5PStkWEVKKG2miDTCEIytWdG7Ubg6
D7gJCc8OT+/+nWXu7HDu5GzwcUuqMW85unsVQQVjChSl7iPoXrjwyw1CEhl2
CKz56S3tEYdYPhPzeSAuu3KJQ3t1cpqhlVsTGpNmscPekY/tGAj327Kyi7jW
wjIO5BzxG/vilF6C/mF0ntS6BoyWtv2l2Dy1I1o/DODM84Sx8pILM0VIRBHx
mDsK+rKlgsfzwv9yKafex42pG9ukeknW04ip9MXJzM46hM1rnlhAQNRSxunP
0VexYpaZVcW7gQmstrZx6areaDxEj0sypqie3SvwysfEUdIxfKaPHGzPXRWE
XyzIi8y2e+TPP8DY7a6Q+zs9O6suoVFhs1JH+24ufg+ndBcxtBudD99pcUyx
ntrnbxGxXWI432zROQNC9mkdKhJrar0WczJW3V+9TsrJ1c7wh7VNDKAzgCaa
/K2PYouH3QNhZRI9j6y10Uox0atEOQ+5q3pyXHIilJ9Vh5eZBolAUiev6qw5
pGFFxt/W1GlBiJHxLnH8c+O+2QARvh9EeCB7jolOoSmgY43Sp4zFIcZ2KxNP
x7f8zyQeR1t/IHii6LqYTNaOQcKfUTScWA/HEPghqqE4x6IPIO25x/9Q0jnh
nDjj51Ifk5X20lBxJZ3sbqSl8ZRDLM7DdlS5CAc0uXExqB2OwXIpo104l8Lx
c0eie2iST+lQNCC4+X3p/r5KiUo7ZLVn4D5cLwjywrk1lTblirCok7GSJziB
SkigvWDouB7Jkje24Ac3oMwS8TAWbDjPhCl2zeMvTMc7mn1GinC39KnZHQyM
43uwqxJ37zRCTeB9MypjiE7Wl0e3IUFh4+gxjj9PHeyO0Zo//DpoCinHlnqq
EHfKexrSqUg982hlhVYL5EEhUwUiSkPWmxQt2qOOvFEReYQjrnjnYiICsvXM
JGzY0GYBBd030Q33KvScJJ2wBLpyQ9PKA9jQt/NQ58GEueehPUiBoq5ijzlQ
Gk3lLz86tQuyJwJrl6ws2/tckRa15zsVsaQpFLyz9dDjyoVyCws7PVDw/lt1
HhnAHe+hJAeF+U4jsN+zoniNNqKPYfVYDBG0hq/XG+GXpCLh/yDUg5TNoIsM
2ywNuwKKOi/w43MIY9lEU5m/I+35nq7cU7/9CBecVWHlHNZageWvzuCJnepm
S+tMrkd+JdMVs0ngBIJpCQN69tC1W54WlDP0r7YgWzyovTNARvkPCDoF7ZA8
sg6lgAafSQSo1COTCDQiuLPkRBGdjYRdfe5KXXTtuyG1/u/D8w0JwvJsebsd
okl6hjlXAY0gzljicdLCfY3fEmmOQVSiHinUcKsni+chTIjTaqXXpbSoJrk4
yK3W2+42NznK6/uCijBUcpNbTocmEd4KedEoPMf887i4toHKbKXrQdy0H+G8
sTx2u+9W1yPw5oazDfPKLrC680HF6YIvUA3Z0Sa1/a74A445EqTKufmndS7d
pPaTDlQHAW/6Xr5mq708MqfU6LXJYNZuEWbnvcTUde3GBuhjr+eOdoz5ipGZ
cH896AE2hsO8UvV35d5fy95IW2HGNifsVX85rBGLKo49FKwOJsxTSqr8mqK0
krFzq4LLvi4ZwyBDgGseAe7OgAnp0eDHb91GDg82Lj0HaRTojMDfLnjnyEFQ
xZYK8UBzGIh4Z+iQmmHT9NCNVmX6JtHdOoC7Ao+ya51YbXW4rG4zI3XPqPm4
qEurcQgFkfUIr4cuksCxR0jfnZr0pIKgFOq4C0+/cVL6Z3Qf3jHudpIKE1mI
vIlzApQh6BQRUy6G+RjojacWJukDMXyacocW7p/7c4XVgZXUtniTs3ufGO0o
fb26eKTYGA0NETjm71qVnsKMJ5rcwbSJEr0aL16thRp0m4YV8zajt/m2pjbm
hifOEiLERaRrDLai4/X8UlmVA5CgVmwgMutUrbeoTcEwKQgVVGXKtesb+Nga
rolnBWNgbGxBLRnDNZu5IY64MFKrgnw5o/IuXNK8qQYHPafpeW0HVi33Vq4u
lPrElmMe1lPv2FVLewn9GZpeK0CnHNbgcOxWwcz9uQA9ef2sE/F07p4G9blz
lLMibJAXc/nmJXvTFmJwOXREVzHqw1BMXaCwaYqipGFZHuHohay1OymP4SjP
w4tc1nL23mYk7E0elIf1Y9nWYd0hzLNXWt0MYy442djlf9y7BA/9MwngJGTU
kR6xJ9Kv9Hyf0dwUZSkK8Q3/nAqLnOm5Z99fpI+vAqbthi6/XmdqNqX0SM7f
DS77bbUpqe2WPTCVJftMEwsq6EhJiA38P+ypAIc5oLZcV/4TeZlD89MvKbgy
nCmov8mSTZgyoLE30KTxliCKOvQZdnuX6U92tO3D5kjRrbQegTKAErxPfepC
z8tu/vIf1RMM+IckYi7OZpB+XGRxlTv+ITvL5ICcJr033aYKhWiFOyIhZl5d
8Z92Y0lquaaCwwFebArgBnYunEJmtkRDd8QeCVcENOpQEL/L9xNf/SRTtstf
KYSAwx288uHNN1g6vCVecd4a8zUCPkd/Nd6ychtkIVfJ72GK0f9PYumdBGi0
RWBWuotXOMPct4lci510uKgjtW2QdnqGDvlAg2ZCMe0/IhPNWigPpPnx/rsI
MQVddriXO0FvnzL2da1fFfW4cm2rdq2G4NtJ7a8oHw+Bxn+Em2/IMZS6OVA8
vWySh2bXwxF1pUS7zJ3liPPBgrVcHx/3E6tWGxESPh0TgO8Al51jXFSbb4W+
QGWwKWVWJJnqYg516b7My5x6biYGLjeI4klEqtA2Fjfczx36yczbCeXz3F0T
xa/C7FLlPLb+RmhMgkMCXDrtxMhEq+eAqvvWez/ohVAPzhduGZwcRSBRUcYm
Zn8n4SYc9HiYMb5bm/Lst2sTRDiKiyiXqntz/6h1R9GNrcJ0CzbArIBss4ZX
OQXyWybIvPwi2UO9R2SRTT1bgPSJxomkR/Fehpa1FI596O5x/2pYoxdSBh6A
/C4xhvY4qaAbAoZOUouhwE2M0OAtt9aXhCKb7e3CPTV/WrfR13smZ8uMD2+r
rXBVVh+8Q35un8e1lMkDCBiChP0F25LwjikdNReonnQea51JYCqWitTZdlI3
iESs+t6TfrmTADLaXwYy9bU+79D9uh7iPojCX89LkZp/Pi+Qwkyk4CbyOd7z
b87pieicmH2UU1TpaimA/XtiC6Va5z839NZ/6NngPt09S2dKjULn1vZdMBsH
aeTLJv5F+Vwc5lmRGEURgosw++sjzLPQOIBqDdbpm0J8VJPvDIBoGvMKCoZl
Tc6fy07ydHHSd7Sm9Hqh3Za+W/hlVaJ8AZhNZFtATph/NFBTz5gae8nOxVO3
vQURIY57eli1o/1L3AAHIMJ6lrgid0caxo5L4l0RWwhPvwQBhS3bxeYNdV14
rvU1mTWs72TK/vO6SK0TwPDsL+tlAKxKApddRKf7WQPYKcfSd4GdDMTcGKnL
BubR1LeY5WJAUypNZsXtF3rM6ogA4KMYT/mzZVgup/U4EqDv7KLEEX1zUPGa
MdNabBsu0Y6C9g+rSlNlXYgfFGYhSgZMeCDLlO0p1t3SHh5cRc7uIRA+fnws
8VU4Vvahf6bd24PWAfvIY20AwYsXmUGS6FABdtpWK5PKRmjwKLb6K9Z2bSX+
rSIbGPrbSFKH6j6pDZ2+mYSrh+Hqc3eLG0y9RB0WTdqxh7gR9ufB5e8id9Lv
AjaXVrZjKCvBgsRf7zAjbBbba3F0gVCbuP47cQlV9ixuGnVFPnAd82RRB2Qu
FZG2uBazgkGS4+ExUzuxRHuvIh0kuIZZUndFa6cVjerusb9eieqULu1AVv4K
V0D+P2a+T+E08m+bPhWlXPaVS7ro0+/a4DQrSQMqocQ7QgRiMR54BB9XbCem
QqkF0QzQKS9Y4tRPmtWk1EeSKJYeyIz/w4Gmk1ndvnwm9ST+BDlNoLi9m8uL
XRl6o2dLfgbP15TPdMXGV4kWs/y80z+rUc0cVsX0mf715BmAMQcmego+r7BZ
ntkGgjb5zaNWzX9uHycj9hqaOAs4nsFUSSeomNxzuImVDkExrUVaE3SL+Sil
0XHimFiIIiMEf5EV4yKd885yJQxQbBDILCgqb8p5FbVisQc+NGsxlSFo7Spw
ZxpgEKg+P3NMReGnHg6NH1sEMfSv1uzOYq452E8ZyiAFEsjcFJfiHSpVXYWb
b30Iw6RR74BFbT4uSVbtG++PfHPrWq/UhLYXh53qwb4o51ZnOnzvF+W+a2pv
CRFvRhC6fNJMgIspY2TUs1/xl3QO2ifjksSr/fGcuC/9GvqwceK0y4NSCuAb
me6R880R1RmX7Gk294FDYtHM4q9paV3eWjywcCt8NOptBzHn9UuG3Dnzzl+K
Wsx6Q5qyHOnOn4d90hTGgevWqToSYTi6HSszjM/rfXJ2la0SnW7wVglMFh+Z
cC4GLfN4fi852MyjNb6SUn5RLdjadV4pO2C6xXrMq1zMGgBHq7AN0wOK++Ln
pfjKKE/rZT7IBuyExopCye2ZtnO1DeEQPoghwydNByahz7+VvwlMcqARIL6v
miOYqMvRV6c0xugNkl2q/Yt2aP3ZeEQLLHeJfPUgMG+3rJh+vWYMV8gimOWF
yHVX3KVsl5NelX9CXtpjURLkDZ4phsnLubCDH16D1ohC4tzlb6YTpeWjaQsK
FTqF7+Vw3i1NSGs4MLQOOEq1UxfeSHZUS1iP7d3dpRZpzGC+w8v0dQor9k61
YwvmgG54prCo4e1eecYeoBxDxiQqPm7yC84vT/76w+RxOfkJGjmKHuDwFgse
d1KF9XehAzPLchFTy0jtiNhqD6sAW6pSZ0g5N5P9ML1exL12TEhM3hx1fO4B
lfYvq1Z0EH7dmBwuLs0OIy9mwH7l0FihgtX/dJxA2x9sV3dW/Ks9cdM1mYrt
pAB5lMXMiqJxYBo0x0Gdr1IxRfvR2GPjjZ3JuMobVUo8gvwDx6n5cRAa545K
TwZRcFVv722MQqhkYOaguzddrRYNEYId8spBFwrvmbZOCHssUj5nC2ugZHK+
nxQrj02I4nS7jpg8WCq6C2k1sdo1D132G1goGM2tGEsO3ZHV4ir6SRj2/yEW
f68ve3fajLGTleVIOR7m8S9M2iXBGyZthBK0uo6fuckBPYymUCPFTs0qAgX2
zFAH7AXoaaa6mbYLwazQ0MlAnsmuAgCqT91MbqglmB1bLazc/FafBNBYi2oK
r2gONL/WM8m/xPUyuuNo+pACex29JemCe57dyoVdEnuM/8TNRgFTUPAyjdxW
UR+rTZpPzyfB+oCMOOFbHGAtTd8V7Q0CT3LgamVtOJhvE0/gNGvhKbv3MpZk
Fj78xau/RIpuNn67xbf4Y39dZGrlW4txsw0Z8Y7r4IBbMYpr5qgv7QV+krbX
g8y3obfA0afZmn3Hg+ynN8kOaLGAzpW0tSBau+w3KYTy3FSqTZbDxenYfRAD
lFqkoeL4ZRZaTWw9U5GyrxI2dwk8tweuiJNj1kARymFGi0PykXi0NXt3dm1B
Xa8Kki+1o1PkXtSbPeZEBuGfpNyXQymKmWXOpLBpvH1LNLnmSW398L9DEoM1
wndI9D/CsCWrWODaLBlubMIlGS3OzGbtak54hxqBECo1D76TpSPWFBecVnsx
2tvplI93YVLOEtfAqIZuS3u98vfT5ikCinyTWGnw4FsBoMOpduF0BkgPS6yw
977GABfU9Y+eH4Fzf3N1KWnGhTXe9xYGd8UPS3LmVTDeILZGPgRVQ0xk6i81
40hnbo01i7BPEnLXxC6UVbOFUWyKN9lzWeElamiPZzUI06sg0ZYFzvvTuHhz
hPNmzNHWTTg0TIDjqbl1xwGMqtwKcfdimBB+UUjwCe0D+h+T3i9UIEHrrpYi
X9uC/QUnkJ5t3D5F5OFPZW119DKOf2MY4ZawnKj0TFGO/bae3MOR1wheRC3J
kIih1xcAznb5pu3Ngxkx5vuegzaxPSsoYktr1rUgE2MZ1+iFm5KQfoQA7wn4
igO8dPnR31vCVWig2jfhtapA2eUX5hnHHnuH/kj9j7t0+e066S1gfX0Xs64X
vU9gURGbpyzrkwmW5RuvFzrJHiei1bTpyI+1zaWBXGUykPHRwUuZ+oBWJ8wE
ZsjgqJ7O6UbDzsL+4eSdn62dAVRtr/j6U+RRBOKPfQq9WtIFpDef+xCUub2m
RVn/ip47GceWWemTT/hyg7oDNcLHwMZOMhcKgJXpM6jk0m81SWaZPNuxqZNE
21wR7gpWI7ry4V99yMnmZmLLzCVLHnvkwJwDyTDf7Xfxpd/2M6KrwDQJdQI+
yaiieMBq2IohC5SNudOeuuUnbVDSx0bYqTnHn1VMt4D5sHj7ZbKRs3EuSBDh
JWxvQM3/MkE+8jdZbpf8QQe9xo8+AaTbjdQ3q8gdu76LM++XlOpOujmaBE28
KTq3ofjJOSZrGq3MhVpLfkQkuHfOiaYswid/yHRZgZIV3lcabaAyGYgCuYpO
c6PV+rNNAITqwxZoWJ7Gg6zHMSDtXUh97FxHUdxM8RPvWpuqdxRxtBfl2FvA
mmaw6BStHw8oVRxssS/Tu0vQhLaW5SdhN3ptKOHzYWBe6gIjL9SyFQNNGQW0
SVAfvQ3fntBOto/aCD9jm+qnsd92PmUSMz1FxTKSd9Ni6KVWMD5RA+f99BnB
fHVRh92QIhUsuGzqf7WAhdClBaYSjEESBJ8grMjlR1YtEMxOp0OlmrkY+441
IrXHCv9yb8s+yMG+XQ1qkY8jnAKxWe/CpnjpG2A0o1wgWSkE/J2J1ekskcW+
jW1t2SrtWbMgb1p6gpCMl5hTYBmQMe/ax0ZVZGKJD+wj4CjU6TP7M67Iz2ZV
v9KYicPnNJ2yzCvDL8c8KcNHU00Loft4+qB18jiM3164WpurWxjEkiC1R33H
Ppw3BEOPd8Mbgnw7v/HLZMtzpswuv8lBPZN/7JH5ErJFAVe0wcArerKyRhLw
9l7CCTd78hVmdgrl42vOea4pjrzUepb2D3aIAEfOENJZbIUsIgUWwI8R3cKo
8yHP5Ar5WiHWOaByOgY59ltykKANEGz4QM8YAk49zwLVBAplVmsFU5YZk2Yb
lpkanBQ/irUXvrd19XEL5hhPofMDJFymfY373laLvcQ3K5RXdb9/o3VzHBVE
R8oS+1msOzwoktimhAaZIuyVZbZIZRfOzmVMdqn4tFmGsh0XR0e7yGy2a7H9
sbDkJt2+fkk10MvERNrI4LjMXFgvVKI/ozJxzEEvmBgwYQlapLmsnJssWh9m
TrPhnLdIQCpxybML7SMqWPqEqV+Nde6GtKvKijvwp7Kbo//OrM7Bus2uO+hM
PPVE+pB6ZVenEDZyLVc32I46tXB9mjDfYoQxHL5MRgfab9v7PVA6DithMs+2
hyQARzNw9K2lQsstOGN0PJEiqEiBnUzgOnF6dpQuNGcFcy2pLjbcbIT8kapi
zGZwR0vP2RpS/ZYCmtmLgiZpNbYFggOVZvPc1ygybdS3iI7vQ3SyksbBAYYV
aT1TcKjKLzA/ZK1yl53rpgi4B1GNcZew+6rfBwikQyY6bt3gTGbXY2nM0X6W
1GPyGm6+vV0gunp6THYsBj5u0XpiibhQFXIULLs5tW3VRhY3jN9uULjl2/iS
qS/QoRGznarQFP0X5Ft7UZetzmnW2J0lEJV7HId0x20xuDtZvjynH2NkcnQE
LeekPI4SYXYtcpL8lIVDUjqNZy+nUz6H/G7MZR2ZtsRHrZeAPBG3UhD23tjO
wcvHvgbSh4GLDQzls+OkYaOEys+loceKTe28D82B+J2X20aeru85YA7K9d2D
+c8ohZcX56jRhPRHCTKpxGTQ0UMSXKoDZlW6SnJZD2/z3vf8CsbGRHodEF0d
8lQ9ctNtHFiSYAjdualxUk0wc8+o/9ybEA0Veobk0mkJD1nDPIfe+Pnv5IgV
OpzFKpeHmZsOdSt3p7tByz7C7oUtCJfatvW8mLPZC+1xwE7Gggzdqj77A+d3
wJ5hK+Q8CGgNdDHYOE/nCpD1tAB1fbMPi2AzZmp6VKpLJ1SCJl2+SkupafPJ
zTRDvdblVeT065N+XgRIavnh1FJCW0Kylex832nRPJGprjjV5eTmhT0/kliw
9TtsUJ545DbCueZan6wJvEvDC/9Q8clCHc3HsUFmBLd6toCV1KvAr2F9Jy1U
PBysBLuEfWJVHZMLke+ZbR1lu2Eo3mL9cQS8MY2w/YsbH9XuIxxK8Fq4Pafh
yYcHB3Fy94YMk7cM20/O/o+EeAOy7fI2QKSQw1Pyzlq/oVQqAcwAXoPRqCr0
PqfAFMMLNmplvq4krHAyxbx1wRi1xRtBq/oUyFHk1jSDTHrV9LtJ/hAtHFuq
TkBZS9SWC3rvJBZLGUapQ6PCrDjUReSdcPuZ7GiwvpT0DAkBW4QgTrpGgGVR
5DvxsKOQG1frW9tyRu3TqCIKu+RlijEXVr8TB13Gxyj3bWe4ISlt/rX7PKBm
Vcegnjs2YVWCQlOUDSK3t1Nktux8TNbzZpBDBxyskXabgKXxFvxZU/vmB0gH
rQa3Deoe25gxFikQZZ9stue8cMs/zqLfMcN+8N10csGG4QGCb4tZI8rcKJQ9
BuJ8MXsi2Lxc+g6WZuX+nusQqqguzUrgjltBVexJ0Fe1HHqlrF0D+A8WOB/B
EtUw90b4CdG3s7T2rj+IdJXGscWzRJXzWokaW+KF6xmVRjrgoG9BLVuFG5LR
gx2ZdF2XuGKyhsCN+hhVKisLusMUPttIC0aUo04Q4OQAazhqB+GK41zxAE64
I15CiA0HAt2g1CjKMyvyVbTyGMY40cKAdUMTbAMA122rBKUxWDWmkGsajQhx
LDMT1z9l/bAKARZBkc05+v0zmp7XHONjkW0LF9zo+RJVFhoLrYtHBF1Voiws
xH26AiyxbjuGEd8iv4JUqd8SjHgwtGS5/Ypnr89UuwfEtOEfpMsXIYPV7CP2
yJ3XWUbW5PHBpB7Wb8vBEOz+/wN8SnX3yoOz4EnHht5GxeVxuMlxsQWp2COc
1/ovcAu3KiR9B4AzcPLz7Wf03fhGkM6GfGkPpuTNxk2tq/eJQGE9igPzlqp9
Z9dPiCgotI/q2Erfu6Y0A0vU8WGmGoEO+jXAAhJsYLESb/iIYa2X1K046VjJ
ncY3jNtlaQGvkz3WDqHZjahrym2mvbYxBXJYSUYah28Ao1MN7KtbMUt7l6po
lbg7m5jX8IOgeH5f4qLsskZaeB0vOkN54f3kdM17pRq9mynyEkUvmBKK1mjD
kHvfGVXAmxVDsEQ3KoMAuR1xsPdV155csKi2he4DUme7hQd1YqKalHw+JsvT
5yVb+ig0KZlezqn4aziF/3luhZn9jWxvW1u7igIp4xQwT+FJ4YA50fd5/hgg
getr/n5pDsA+pfxrxhT+73IMLOQyCj2OkDRwvIM6XovqLiLjywS8kjhMT3Ht
Se35TIRohfBfnRos6w+E0q+0CehditX/DJmP2C2jSxAhJ6cEurNoEAM8EV3a
0GhcXhIEfPeUzT9AYocR57ei4ZebNb+xxRGuHittIDo8jTolhqkGbjBU3Cmb
4SJwv02w+W+ZtVH1U0ll/68SROMxTGd5S33E2wX+uzadkPjO2+vYd1Kzw8gn
2qwNjBhbNhkebIRlSn4IfsV0ugZC9BIGGHuCXi+sHSwm4A00y5QMPpovoPNW
FYxcM5WDm6OqXGX1OnsaidRVGYtDGUoNv54OVg7AmfmxfAm7SEwwwx+/xTrQ
BNHS+q/cMPE4ZBcBKQWCV6pM8X1ZqLLY/01mC4XlFG0NYC40kFaqbAeVT4lC
OJBvrbCnETaE3+qY0dqyNRaIPWcAqtA01Pf+lbGskX8OUdZgeNYVxN+3szzj
VuJGn+QEYcHDWCgzoFw7yK1lDDGztXxvmAT9kMWcBRKDI8HzJNescEoyIz5p
+e/myOAehg+elQtaIVNHoXZfsx6v6oHlmJxt9To2mNXze4K5HQYujloz+Dv4
g0TxD/cTU11k5Dst4oOq8x2SI7NEk/sCO4RaYcCcCyMckDJr+4Wmr9eA5sO8
gnjdnx2qVcRqCVzmwGY1rfCH0q4l+NfuuRe4UNl51lLOrNAh0o3qAi4HxuWY
oIs5NBGrs2CJCnC/dXmKrTJf98EQW0LKxdb4I1K7e4RWBBNrfdHb419v7jQR
wtC39WR60mA8BDe1wbmvNW8+ftY5f7cuZ0iVEfDspxvW2q79fZ04SX5VduJg
8+xioz1/G/ic1CnrZLPKpPin9gSxc2zl/U4xARYXZkHEQIRreNQSjfsgLDY9
+AIOy7JBORz4dzhUCnHLKY3O18bewhEmOEZiLuLUxW7KotOONinuIN95BrCj
ngYpiTMSG1S2D6rhYXdq4uLBvVS7aU0wCxecBmmPYp+zmT+CX7UiuMHEIwV4
TlgWvOgU0nS9SuAiPBZgTc78ctSXg0NiUTJbHRQxkmICPdwOQ9x92IAhG8cL
U6HS0yLdULYt/LaQPh1dybDJkymCrDCfFCJy/UD79iZZIX526R2GMrHenYCg
CWbSr6Fo25CTyG7/z5MAAJOYCrfNqiR+tzE6JYYzSxlbzOntE62lmvER6S12
FhwuUsrW8xGdcjAn49KEdQSG48CmhVMgGQMgdOZEZ2gFrg9cYybz/BFNKJpo
EU3qnlTuNbUwzFeZHfX8IGNTfxIqLb1ehpxxL68KEHuPRq36bK7f5gfkJKVI
675pvaQFD2/y1P296QK0C6FbDcsrW6ZVG8pf8NCkoeBWIS12ewOTvQgV1e5k
pAnjKtnRNEHRyy4Sws3J+wK/E3QfdIuBOvwjP/u/B1Kv2i0PHEONc0VrHGlU
r0yLgPUlwk29UOUEgxt+7TdBBesBdmt/knit0fBgc5vUbZg0sCc762YzjW2r
a9VoJ0qU0YiiLFOS7loqH2NUY0hODnxkLJcRjDbil5iRhr0jHmRpGziau0hU
gL8sdDeYyr9gT5nRHfIsFPJ+rq6Qmw4xDJLdJCyuulsJHlH+8ROdEm+CSYXg
iAB7wvFsE0Oj9OI2/53vl34WJ2TH/NjjbEjnOlKnYEDI2BJ71u8TIgPJBD9P
0fVVvUj5jnJWQU1d99j1oYzpEW/AmkB0mTaO7wg09m8uoOZlOFEHAjsAlarm
NPutae4QHWY9BD/jp8CnjNhR9WhNvbVRde99ruK5KCb7olNvj9CdmUbWDBUZ
pym/jG63Mipv8MwUKOV9Jb7QJpT1/FkIBJ8+cwGVCHJbdxX0evmtsyWlH+9j
8MbdFsRBrJEB5p1xIM6/vF7JDLHF2o7ThUWaMLLI/bDeq23I855yIP8ItJz4
2+Ji11Q3yopLCUNvK9Y03nRChV8gpOpjQL5fIvESV3mU5plA7ifhfKHfEUKZ
p6qbP4K44UxIaMFPakp5lRvljk3wRJpZ5RMx1qCEdV9TIXvagZSa4MFIauL0
iuanD8FcR5TifLLVw1TJpFLrvWfsosmqpQuyi9/87Y8QEhv/O5jJ+gyCPxI9
oheFrf8CsDSSsdxoKZOz6VpN8s6eMblFR8zt4eVfNhmMIzaZWFaL/D89iFdo
HfOJgrcBAyrp29buMWnQCn9x97d+oqClqrVCE1TVuZRCr3ebDvXFraHQYdGY
6Fj5I7ZMyZJy6cOMZaCO6subcMpLTrJf3Vgb9S2OkXNqK0L9UYdnCkhwCAxy
BYSSMmj/Ez+38LXSAajkJrWqvhp39AqO+1egC/Y5BKzfAIPSczd4cj28dJec
SZEdEPBCtFD0SwTanYDDti/p8wcYCg+ixtMe4L8pvIJ+1uo1juR+QFi7rkFz
5+P0jQ6mtpm1kJ/fFaYb7UrGWCnEgv+uXzIIyEHnPxazmruAqgMNmFML/nn6
aYlCNxrcUX08OjuZ0towHSN5xUGuxD45a8tQM9SPBX6tcv9suozi2gdja15Q
pPRuXwxq5PxFCNPJK/eH0fTsu+ENvVr60BjxBuE1kK9ChFN8q1/FI8lL8DWv
ZPWPGdDuofHJYAyxHwn14ISf0IN1v0IkqrEzkXEfYlrVIcMSCf+PAM0j7DdM
WqlM3XsC9bXavMs9JzXd2HG4wsxuexviUbawcPTUNrpK+ahEUlTVDUanGMl/
Ape+wGe2PQMQa0/ccQduT7j0EyXCdk7CJf8CI4Uol4/fUpTncK+Up8Fr91yM
B+AoTyJdU+bBiEndhCurNpN1qGDJxXj3t6M2DsEgLoCCSGKdVXS5VTZ+wOC2
z3PPuGuB8i7YdXiKKwR5UapTTGF/tG4hxB8Uo4PvFFU8zxmpg6HJd6Ph1zSJ
RkLxDAH2s7OGlhUKL3IXMSc7iImGHnKbLRHnYvBtiTT8dzv3NhhgcOHPpUAC
qrIOJobnm30dJt4tS0DYakrzX1emPQY92KB1JicsSnDmBo4ZDAaOLw+1J2x7
iHPMEjDaQpuYqqd/4zLT0OPTXdJon5Gdf5F6LLlVP9DKtfFZClPeuD1gNgmd
vL/k8FOGrSNeu9Ow42l1NKQI81u2y0T+ETATwCzYhmwUNLuVzDOTTlHRsybA
D+KnM4MrMCacqRptBLGQclIl/CRdOTtlG/Rs8iLDm+RStbCWBUmWPSEnwFHH
0WkMqlH0zxHWZiuG0Tb0jLHqn8kAYgB+OfPzMJLnox/7a4hL0EW9ATNDEy/4
DcptOU1VNnn+hgv+f7xjPbx3vKeWKBZEt0xVyoK5ZNI/gwXfySc43vIEwrTi
krnzql1pmiGLUDr7nbRwCVLzZNHruirmYyfKbiu5g0wfiZR6DJ4EHvw7U7GA
0+xBk7XGtN3qrKUMI9BLGlf9f9bpaF3I05foXEmyPJH+t09XtEjVAT6b3Vla
OzTuusLkr1V+UPicsChwTwSnsdtdbhAQ28P0PYbWlF3QY/XzPHtGp5JKimjl
HOkcf1gs3EYaV1MwSkcRmDbydstsZidBU/NkJ6cx0DWVqoQZnxFuQtA+Xpzk
w1EQds/kqO/yp4Hi+N9ftzb7ADWPNwP4WrYrRWjxjOpbMACnpBqNlo0ZbPSG
QztIBec+4D/46kfQFQyAC9csFXyy7TNPH1l+0SselZeQCv60w3hqGl5S1SHn
Be73PXRWK2P8PNsjJRVx150tVOC6816Fjq9sb0B015GNTz0gBOw9rQJqOaxg
yf0aLi/UdBMKiVwaHLh2M6X3w++siVPqrEDg0YuKA0FzeL/hWWWDDJvOMwXX
8/vYodOyh2vNh9lt7NfwduDrEDMZ9bfrt5/A0rGHtJ2iSX/X3UVqBaOwZoDu
rF2zWW2IWSbQgcKwJkjBH99/srShAxJXLhH9q8lpbalanq5gKgtcE1VAIzEA
V0ogw00o7dz0zSWwV/rgr/s0cL7ELhfK9t2z9Mv1xHg7VJEfYjwVOahc6GXP
ctiHnqefc/yFRo9Gvi1XgARJoOJ9YfcsvBiLrLCZTlW0eKBssjfa6LmN9Lpp
0Sbs356vxiNp4UUGbavna2wdnbij2SRt8kUk3W6VAPep1qv8Qy2+ZxR+4GdT
LTa7kNCac3FLwnqgkMJHiMxafQxf+L0AUp4Gzj4obWJXFNW0EU4Sk9o/csmd
3C0syen/GBmgfJBh1ZIU/D9UHnAaP31rNA1TUbO/O/1R/x2HumkI5d6kEWSF
YMHvHhuYVGck27ai2D9Y0VtEp5Q/DL9XHVv5ZpVuEGLFUjCYuv52U767dM7m
E8F0NZ5J4ojP3hpynG+VSCGX9VHPwNW3Bt1jVQoIIfUOOZFhVAvgReRMKggD
A9LdTVk6zIKk4dRiYl7g/ZvV/L70K0lb+LnQqElJ4jP0GpXsVWwbAETmnd/r
mLFoZrZinHIj38UNV+8vAUa1iXibv2qipkt6FHAxFqdvjCqyKSdW/dBRhmKf
28yLfjC9Hd34u15ZJoDMIqF3Nxgw9lA4HhLZeWSoR1Ey2ZPjc1U1GjREwiJC
ioJkM5Jgnd8WX2Vh09jGtltVASD0oCzcW+xhk/Axhw8qvuZlsl0cYA9y9T8j
L+/UDOwXQy9A8BF2JfWLumeYu2rbgpMTmi3W9W+uxLXpHr08JEMja4j2jjWN
LwXD3ClQKUASGjTZqk1+0pZQ+AnaoaRV/9OPHOi89qyInbPoQ5g7IQnvWYnB
rhawxzc+DPcAtblYKdtmWM4ALnV4+4f8G2vpYeUF9UiKBJRdB4ctGQXU7Vug
f747DnMRfjRA3lEv3UjzikzMOqCIHdhvUl14XC1PvMjrqHrzRIc0SqlP+Ut1
rxi0x3GPlstSpyqW+1ULCj4PiNlZJpwGsn9llWeenCZQa55YKYYFJqjI3q+j
FSbFLW1GbpFTJWiBaZcHbR0iCL6BN02kdI+LG5Mt9yLregS+2I7msEjh77Zm
n/gEUiZyUGKSVQO+KYSZatcU9dKpELW/8zV1cEUocCa7BW93UTfZLNlU4GCK
n2rT38+oQO09Q60F/zOavd20Mue9k0vhzFo4C6CZeV/jcMDHJrPVpY3L7G5M
XvNV9ob+iRKFacNv+r9cpSO5TP3PnWYCpvbgvigo4yE1kNd22PQBRUCMP96p
zGHxkKcTfpzMRdqXJtnSeGqwNf15dPgrb7C13WggNdzjQH41NwIG5zlHSSi8
ves9866zKxZS1I/wJOVqyb9SfIpvkGgzYIKqhb4BRSJlMBijtUWvIUK+89rt
v7fsuSKmcxoWUsI1h0ryztzsMIJhqMT8li3uEpQN17VrZOaH5Am2xerA6JvS
gENAXaY4pt0RP2eEAfYcr56eP5IYhOFqzlctDrlTuxYBh8bnISqgGw7VYMa2
nwcaR4jS+p1OdJZWngbJLegy374NZWlJdf3hJ0r8SR3Rx6t42aZGcsBDmU5Z
k/IeU4wtXigpaZfXOVX9mfgosU5OI2sD+ISlGClDJOLER1HE7VArHYXXNJ6a
pR2JVlEHWjFbMbn7QxfX5t856HNFMI/xoJEJrTfFHnwf2LYiQ180Jsf2kvl9
zlBJu97QrsASaHvS8TEFiMAjiXwAB/T0SlalmMdBxJ7gmbpBpffwF8QiyHY7
4Puvt8wKkyOTvbkj+K2YhyvE4+sLRn12sfSyl2HtLVkC4eDnszutC5Pit2ja
JJWSbhskUKvgCE7DUnHFndjhKyTgvNLh9pkrS4nNQTWDE5FvN89Yj0R4UBS2
rQgQpxHr9AqeltHqytbM2j4A9Xicz/+6mjHCwkOxm9cbxH5SVtutzl8ZK5xw
xcgFY3LhlfvAL0xl5tjhTR/82bXodGhVkqnycsF3Y69G6DNQM0dvZnepeSn7
bwNqWOMVdjk1p3bq+iT520qTPxSMf6Nm0VzGgDFz9m8h+xiV+R15gOMiSsJw
nrPZ4ESoS3lP+cxMF6++Znsy9EIgz0HvqNlhXXfWhNgiGo4JJ03wsTHK0ooY
wChaCm3P9w8vSJMrqb4sejso9pkuSkw+clxHgh779jDPPEq0fmx30cQXMQ0k
uATKHSnizhoN56kd3iT68VUQjzdMOMUmIyqGXw90Qn4zd8AAchNzpM9lGtEM
iONrk+UaCWzxelsetxFQmD4jVuXuiLe3tDDNQj7nOjPC9MUp3s2unR/NHBwg
1IBQRHtgngapzO6N5+Z9ruYi/ZPPDeomiOrut9MY56etqreue0f30OQo+A2S
ILHaQyW2iGgIqhMvSDWfMY0ePjpLiWB6oO1su90OA0BLKGcM0giA1d80XUf+
Xv+nn44GjKHSUzXvZWkLpX5Xry5ZksOqyLb4WbHdzSRFoMVYXsvu/rHLWhna
/+OaMeeQ6wVFXWNtSzUDZrPgxCllTLkiKyU2YgJ2cLMsFM57e4fHRkI6k539
QGleDlaAswl9WTqDRjSm7Glu2KlGhqflOe0Mfy64fOw3JWjgHNMMFKZ5Yk4f
gFkO0gDgKygFSh05wFI4X1cR/2BeUi/9kPwCcc1k03s7O1xpneO2hKmxP2k1
dpitBNtaAmTkroMc/zwXjpJEd3+u4U3UrlSr9dqASPt0Dw0wtJhmG1sPCyR0
aQd9PC9beKuRrwgDWmaXtVDujfxXtWYF6heZEC7V1jCVTIDs+0pA92r7tnp4
wpGhc2HkDIljWCfTWiUEtK+sN+9VR+C++E1GqKP0PpqloVtAbFdtV9s1iZFM
Iyr8MLfIlwBMM9/yjAVr5kL4CpD23BMkv2xAa4iUlbAsE9K2mq73aVsscUA2
7TwngWR3khSiah3j0Yh/QXXzGdD6oplYxoYPyTbvlVOi2dEW40Vz69V2gD0w
20ndA3MccTANQUPGAULHbPDKdQ2Yn39NAKhWCi0Vlmct8ZkCBOztLq8bJ5Ux
jicemw7bVKzc4JKoEsdkpSeauf+FS4elxuGmwoxdFulTksZVl1IiHZnB4Ym6
lIROA06DBzkCnvs1YTvtUptS1alXgr+zSiIEc5ADZ40b92O6dyMcU4Di6uei
+3yK935zNlfTG9z2/XFE/hpFcfdTMU0c93HE8EfL+sdbfHxUiFsYup39wEwj
9lpGfrv/hlgUqLvHTYXpnXSaa/JAPPwo0XOKRhL5ebL/UrrgWRLtfqxA0eoX
xkb1lI2D239z6cxF+zUX4t+/dbWWUq/nmwLQ2opCJZquG8xMrAz54lmqMj8n
dxisBw7AayUZp/0yD+RB9CzbWg19auwpONyG78wdBMXAQXhDADPruP2JdWTG
Jld9K9PB5B/9+HEg5i6lA1yRGXUqaOem0BWlEyty9qsEJOoGjXx7VLLPFbui
EPmdpUWVY1+kTpln0thfSmSlbSaFizGXwXw9mTG+jo26L02XLUAafqmMvlOB
tPYgfNQtgfE6y7DnUqPrZprC9yI7oG6dm683aqom2tbvkcyEKeYM8T7gjtUi
R3JKIML4D20gp/5oEjEwAKohyxMocihgZkwfdkO9a2TX4f6fQnR5rzWdi2sJ
JIo8v29U1BUh4Lyo2t15CwaJsiIPqGwNCnx3VmauV3GcVoQ4DKaPumtfpIXO
BXmXsXACXw5K/YRn582F9w20Ma079GwJi59LxU4XgtZvZjTQfPGeMD8JkJ45
GVtgecD5iDUCoCPojmHjDEBebck6quLQyDBxYwyEBSSLgjGw4dnQL0J7Ls7s
hHM2YGpbvYl3zBzcMxoY31Xw98gSYNYY+kkRBYHZfDbv5dI4+ip8QdhMneZQ
3t3kzRoU8wl/SDwdgalP6m3PWOWh8HhL8aseM5lFQtL1Pxbb+nrL8zjsD35Z
glFy3oAG5kY4+hAxWVQ+aDvFz/0RXMcZbB99luAR8mjG5wwEC0EcD7tmGzc/
vyoYzN+FLBmr3mKw/a+O+2Oew8Vqzmv8HZpXynryQkBPvDyjjWsL3N6F/c1N
fvIZv6lvXxb4z48MoJgmVwwPvCqrYnr4L6AiJPnba62b6k2VHQeoXFdf64Rp
AyreA7NPTuh+jhhm3cMbuxZD/YlqIVPZs2AGLJkRwZr7G1FNwwjIG0iqX/SL
psvfbS1nO9OS2bjNDdinr/ugww1lHB5h8h5PlwsFQw70V222NwS0/c0Hb1EP
kJy2ZIOsegXbp0HuHrdoQyM8bF0xe5NYbmkKunsAp3+IWAJqg4bf8zjCMagb
+4nH2oZzqRCJXrPZHA8vK6hqK2EwGqDYE6ujRC01IXqn5A79/ghy7zygyu/L
T0i4A/SCvla+a3F8on++cpLyxzI5sSdqod7yQjvXIlZ/wNcIVz+BbYQeNVuf
EMq0Mh5EAkQvx+eNYHcMBLCkOPyWKr/B58jQG2NZwc+Gpil7d3ROa7k32kIJ
eExsNJB3eABatCBSQQuBc2XqHG19zAJsEDF8c9YFEtoGXFzJhR8Efl7QChhB
7yTNU8LKxjWExNalnJU+fStr6quNTG/vFY3qAe0pc6CSPpojIwpXOCromOM1
xA2/eS0HHStLVn98dVxuvRl/z8e+O3dnUQHfJUbn++scYsjbR5BWvRY3lFmj
scZ+eONLXgIqGpbv4Si+aaoBOhTRykA9uLiyOaFcNrd1h7b5x4NwRV7Nb/qa
U2emSDogX2W/VJZ6tyA54cvgMiNSebr7LOjUE0jMdYvDqU27T154wgniTlpg
4F1FgUav0vU5NCYOcUBY/9A5I4YXr+MnIaD2cPe3eGRiiTWC2Ce6xTilhtWt
7Xyf64WpStG9sJYc8CfxtjxhyQivsD7FvmfjkZ9ktrBEcpSeeEdiz3bmLViG
92PX62OgM/3MMrLl1E/INxla8ppMurvmd5YEFQYo6u8VvLjL0BqqVpkwKhUz
+LecHgvA+sVgq0xez0c7IqV8ydbHq7Z1vQ1OmaECFVbWNX3b5RSIgCEPHLw3
pcp12QUzzlQ09qHpPDKHxsq/f6116w8ZxW0pU3zF+RiWph8Mm6e2O6YSC4WC
xrIpD7WVTisWG2TeBmJ7aANoLH8kor505pmwhhuY0IKdRTPwZrAgE5XfUvuk
0xLcooVkh3LVjYzkThR844gCPhOoHyZP9Eu3wKm/9aRLdpTf7YMN/A5K1hZF
r6eh8LtiDcTLzfAmEYnZctnLlD3Iyi7vMhBnwc3HXvf34g3OAvK0k+w+o66G
8/5cI5OBfj7K4UmhbY6QeAqfVolteFfeRGy1DcvY4CKYUzdSfNG0k+Hrs5Zl
18zUL8C+BsR/P9D5hsoylDA+/Li67hi64dxGkhlOMK5M0YoomU2cHu3rgvNO
aUGuS/x/Wq457FdE3k/A9JLfefjovmk2LGdQ+5uqrDccyBnf5RiQNpYT3jD3
WHpoxpN8+Ux6iP3khiRvZljNYkosWrHeZ/GYHT6Kv0xM9cL6FtUkJ9ugBi/n
3go+52PRAWDuUHPYDUlnR9Y2qHimsrPErDXotYtyNYZ8BUT5e1r7pqFPMUaw
Tc28yjC/8jjMC6GKTwc7vNluPrJwymPd6caFMBS0k090xmd1a33z+k8wXrYK
mpor7iIvAqB8vJODLA1RlMi4QCZlaKzjmAmPCCQdH7v560tjXWNuB+UyU/Y0
P5jT96JNai3dDRnSRqtWVuxaMXuKVLoDVMDpcoG0j9znBRFUEqiehJ7sSSkH
BDfnRhLlfpp+FkR+HBVbK5xKR7biyGXretEAwpmXd0VwMJgwekP7J0p2eJ9L
P6pXNCwWpDQGVxWt8SNaOk4eIhr1ndXhHiXx6V+HBrtSFZn4CitZ6hweO81A
o5VznE6+kIMxf5DFOxNknH/UEOijLZyNfEP42aJuM+mHgTatSkPw8i+kLJ7g
SVeFE1oVRSnOJ588T9S1SzV9x05V6OqqtHFZwJn9zEefKudbc7iQyD28w0rz
gL7j3v43v2D5HPRMOzFUzDrUMt85cIB42Wa1wy5iFme6YSIWsg4p+0t9AeVb
53dvFS2R2PpdXGMW5dSJiDD0inHnfmMyvshR+gppWRbQlF0aFJA+YxhUcH76
E70/zqeqUoin5G0hdHEZNSh65g0HpWkp35gTR0UWVDjONiyCT8Z9woyYG6oY
CZIb3NliUxt3CCIPP/43Zlx1KKCVYBRp8coA52iM6Rn4WfSspk+GNrY3tphX
wAq3zGhFu12BcZJxk+r+rrA63TjXinRwTDfW9Y7vAkplIAtoBpRkL4ulmHEQ
XDQin5p8wP1Vp4aFoFKDCWHsdjP/baMvmhKuo3zpPudaFI8VnsaE+JqH93fG
W61hlkz71wcZCq19X2OmMcifH6Ps/AZUblWj5SuBkE/CIalG9xM93/TOXMcI
Pby7XhGw3NHI/pSzOGY/gzFmNkUwnVRoJ5Nq8oR2l80vOnglEubD79v3nCI+
AqytQNbKSbpA0IR1Nhbg/y7i6SN+uSFqkilyx87mtsS4mYPdmNvQH+J85zPl
grl5i9i6jDHyVrCFTOe700Y/Z3W/vOQccoQ8toD1MHU3WSALo028fLrfYCV5
PFI0sP8744Tof9ro01aQNHyEnMMb7dwAyfzi4WC0Ca+luytjTYUcuG2q77Mt
qDcoNObXQP2TnpYncweXP+UTyXiZD2F1+ujUT2mqxMAhJnyBDHgz21HWodye
4UbO3WVmlo93Pd4fgU9oBk8WpsbRiyPqqkYxHdUSbSc52W22rA+vr83FLuIC
ZtV9WwKDXIzUGiLXbQLe3N+vS+CN04jLwtRvaKkK5FEKbSAxzH5G36DO+4Ma
Le8nR771luk5/h1onjZsKC5qV2It/qn8iXW3iT9SmuEr2txRcecc55/rx8I+
muqRXtCx6eKcxKx2VKKEva1zm6TWj3CkK61fDl9OtzD/Ry+LsKPnqNpipDvb
LLau+YCxGNwPrQ2odRAdDfMSl7MeAFxF3mG/tITpmV94FTCGg3r+gjws5L7O
HwwlkuWJAi5XEB+Zd1Wj9q/qfr8i06kulNGXAaI/HoWJtTyDbKFH/WR8Hpy3
dQEViN8Ysz1RnMEIGzIZwbo9AUDxrJ2P6VVvNwBeuj7GpFrkCqqqUUWaBTeM
d+BhEM/GBOV6G1MlBkEfbexpI0w424HsZWnjwNjrGy2G7+px8az+H/G/dpOX
PCxMv0ffGNl1z7FT2E3oYU4lGwQwsJC2CVDQKF9izOQ9MHs4wZrRZ64yvzCq
YN1ILcRNm6LYqESqGJZPrsqy+GrM3PtyxjvFZXQK85eUQkI0IFbC1+g9DE9E
PlZ+OhYO/j7PXyYujqrCGuAnCdMfRrHbCqyqhYHoZwFg/kwwewylQ2qe8fBH
vcAUrj54WP2Yq/HpTE/pLpGRGNXVH76YtxleS0GdwmDinF8BejG9GzzVxQIA
0mMyGfc3xcfIKVLtAmO2h8tmXHPbPoEthGah8Z8/Zjd8Vf61ggFiw4pIXowa
5UIVZig1wdCGrgPVgmho/MUTuGf3rNVWeX4RR7yaUXGXC2XoBRJKmWczG9hB
Qpr9JLxOXUYB5Sxlypy6i2t4TN8hns5OwRgihHecqqI0ouU8X5l9W5XmUbmG
QEoB1UCks2p744GT3U/ig2kYG4HfqJCojurvQwAUNyZ68vsa1LZIlXF/DLYR
PGaGBDc0TsPGVhMS5s1hmXXwkSfuWLorXehWWmBjQBS/O9io1shENUIhIplQ
7AUm7fx2LI9Nqb1cG+eXXHEg1vYcr5QNxz9uWmwsSz5fv3J6NsknCcYa4Hwt
lfAbU2SkoxrywyNylGtRi35dhuJxvF33Bj2hxrNIskhaYOzoWlc6g9EDz638
l19NmhGGDirs0cnBKPNBwotDijdkz9bovwJ1ctb8N95+b6VtVb4Iq1IYluGa
LhLW3szyRSO72fJDEipoaAja3m8iPWnUNQX043Uy40YdKWGcPCetHXk3a+w5
dkSfVk76mzD2zkZoHcMJpIgN+dRVHunQYASzvGpZgVTSTHoMVw2eWndjMaww
UP8IaUC9trglCttEt7OENOhuLDk53wXaTBCcngJrzB46Swa4bI6cRy5YdvtX
NfuF6ehSVabKNFFS1IZY/4YKMujqtaJ9pVbHYjBX5F5FluuVs1i+GdIgV2dP
qiw/4ZWH2fF/+CnQpvp/c8PScHnLq9bJHjVjnlOkLEls2aWzC01DC3Wrh2xD
+OD23m0zYg4tVNqZoYqqqEBRWbF3Nxp4UJ9h83sEOsZ34gLo05G5c3bRRTNR
mdJZ9uZg9k+QAzYdVwTa4FyaHzgTJCbWxnn3U6+BDHP7oBO06F+5NHgmi3Xx
gbiglCXD/bhpPvjKIl5JZKGm7OAABqbRjsswQDnSWefGJOOYHWRwXJjOUV3L
/zYu8fGdjmgK6nPkGCGRDSz5RXCbpRDyGN22p/LDKcXpmpswfVZhbvLamfbw
cmHBdb5kM9vjX+yaDSDCheTgGFpYMbfwv7F9SnB18IpvXL8vS90mWB2Hs6lv
tuSjSXDbf8s0JVHpXlLPI0SRw/pG9+LzsZMUqKAM1rAagrcdqMlwovq/usiy
lLlOrNLWyaC7w62MXOpKnrs5OM1BnXAwW2Px3deQbBED9jPLr7f1qLKhjmCX
uKvkk+uJtoTmFE2IfxmvCPwNC2+pnWKtBn7ieybsyMmIe26sTGFzOujl5sMx
MhOLaXhZr4W5Ikxk/K/st2ZZBNCdyqtIEdURKeyG/CIxHn3iAkEAMv3ujufL
PPFXQPxFQ8MfgkVnXeVOzeAl4OO09/3DMZizDAy4ptTjcJmXhzj3RcTfhbZ5
BsFy0Ym5OyaDq8EpHTaJmffdSNYJv5HWKltNefvKrNwIAO4KiqY8dRcisWe9
Q+agK7gBFcmABCRFplLVzDlyurxpbcxyfFT+VeBMFX39LD29K8FtL4+a1G2d
CIq1ieyxkVPihAd9HGRlGcRZxZCk1kMfRgvpguvP+I6Cfwofyps3OutrT+zP
aKD46/Vuh1pVaM1wdmJ4zwCP2LxbCviUhKrB42HfS1UjSDoPSTNUbWhgX0eP
SguPgy99HlNr4BerGEiO+rEpo/8sXN3/2xmlikaHObTjjS/pE/P1ye9B+HfF
kU1Gm+ImJP4oq+YRt5AFZB0C0rfcoUrzIWi412PhLaOCDQNxzdJxDSoiC0HC
QeZqnIv1IbJUGRrE2SS2NcFrJvaCe1ejEWCm1VVo+osljzvlSEohScXxbf6c
A22vFxteK4iYY3BDB7RSNW1NTt2/5ZhKJVzi2RQP0ZjUahzbtnrqmPEfkKrf
IhH6r8X4yKoBXeOXklaZXILF0nx/an6pbKtSIGq+nsVsDcAlvq95EG24aINF
pDp13at4y8ezJFSpCluWb1Q4m5tfWUEgYwsryD+YCPghFmDQwrEFIGVV54HI
tq11pyLkdNq7Vm04rmYbXFMasZExwgTYnniImfoSAztxdCPLhuuMgbD9kj7k
N0nrSY2drWQJD5j0Ro7k6JwM+F/0Fzy0DurRis2R8I8vpz7t8a7aBVmQCKSl
KJbpPPgdCIGZTS5Toeq2tjNFR1ahQAZm8qk+Cr9l+OkpxwI/2/CPlo6dl4p6
tOtDbNAXvkq40QQIBr9cKx8wY7mNUwx7LiyDxdcE+K1yFywvbQ7BUCih9jr3
KAGsJXJp4s5bcBGlbm0fIDAiAoDYoHTKlB7TjLtL1ShirnmnRZ7+XSX/c2gN
zNB++g6PxcqfUtrzJaE/MnEhsEtb6Oi1vrFaxBqXjPjbrvic18WZTGpoG1H8
tkzObwIxearq9tUp1zzmhCgefLz+EbChNooyg6PbrLpLzrpCmC5wsTZsec6j
NdhaOJg8TTnmvkpyNpcpM6SArZoMY1NYbOyz/6VBCT98ggkHnJAHJxZUDysh
89SrEjuMT5+FIrzxukl0ZU9hyfn/M1ndDKVBLlFyqBFaX71bPYIRM2SsPMxA
jXiA2amtH643YkslXN8cYxzVCccBZfFuxTRQ2gv5gnRaXVPNmqalcTi1fJYa
WA+RM8c4V/JlzTGV+1QhDnwt5zZjF9Hh2dM02Pg7enM6yOiMXVKYQTb9g+PD
r8gn7mRjqJmbiF9x/hDwa8ksrBsPerDf5ACMRDrQUyWvbvVCN7itGQCTjCaC
LZNiNPt33aLyXNfcPoPAQaX3aHID0cDIay1N4Gw3XKS+Unx9LiJDwO1ULWCA
N9iHdBOBeUAK9bHJM7QF9kZb4mJ+VOQvzGca7v/dUd9+sn6zrW+/BNP8behN
KIw9MQhel80/SRSHmAwiuZqtvYL6ot0IM/YaaHmKxwPgNLjlFKljARY056ca
YLZizG/atbjLxavBKq+kF41LdP/NaMUPW6E+m1pWe9ucy5oPyzv6rFeJ2r2g
OhePm65mV4w+hRyI+XZqXnqlGVOselYM8VK4cv85orSzA0AeJMVuyvyr0Nla
h4IG8xI98vhkKlwbdswnUiR6CHuoI3J9Z5w45zDOP162svOgYXhSuyn9Ozoa
4kV+S9r/NCy+MvTJC2CqXUNn71Q2aZLsBhTooEDYctOVS9W9H3Vcq5UtYt3x
xn4Tnluvvoj2lzOsvZvbAuPqNBLLdLPK1k9HMRBKDlUS+xgYiuYM7C8nQ/e5
hMPPe3LGbbz/MFbbTIxMSDCx5/wbKsXP6WZqAQ4W/+cSqwDSHlx0EFw3enG5
Ihd6DtlNL4RJdkH//wFE3F1WhRfT5WRQLTOKNYxKyjOSBNcK7L7uGRUN1CGl
U5u7XiKJPxnO0bAkmlUo6Uj9DZe1hE1/dbXZFDKDhZ6rpQVFQt4wKolT7gAI
Dgo558yM721CRiB1maAGByJB+rTzse4ot2vN8JxXi6XmchzTM5jv2khPyNe8
oKCxxTEppXFNlJy2ehzzJCUoM88pCe3ABXVI0jz7vMgQSSDXex64WWVjIoDa
SL7dB0wb+aIoZqZ4XuL19TIa8ghRbxEHyIAVXPCpHqPBkGFHENo8heG6qGQP
Ve5TNuq2qcRFW96YDhbcXtvu0k7fJA66YeddPVe59kT99pfotZ3C4QDsVpkt
pRQQI1K/EMCh7FjdkzXDVEDglWqaWfDyf+zntUasZe/f+v1leUIkBSwwKx4w
7ZebBOL8064Gl1fTX9fZi9/58Fz7oN9tDGy3vVsDmawvevD+Sb8JTDUPhh9E
G9a/cDHS+dpiPBQ/9xRXfpuPDSZcKP/Fgw/6DniXRO4LpiwIkG3la9qZALMm
2QpOV0pyWxnsgthsi8taz0ovJPnW130NQbFTbxC0jqJETBesqqHQGaXubWC7
rDabgYNs+oV9EYTcpsOEspI+sR3WzX27cGWaDbAJin/R9lgDAy/bNDYFTZl4
X44s8qtP9cXhcmElVUkMmpSK/1cCtPOAOb5yXk1ikaTGuzxk+V5twRmjhaFb
G4LFySXa2cg6xTkpYWrDb22Ou+NIPhjs1sWsSPKZiwHRb35+CYe6l1IUarW5
LcUEYt27UcmcXpYqwSiTzUSSICu5NhXSZH+BKxf+W4kSAhwlGajL8ENkrQ/r
awDTwhrRhnfz8aBHgHeY5goPlLcFCCJFB3oQSTMMH/9IeFTOdbV7aDWrVw9F
blvvrpCrym9PI8MZGIoVU8MAeclqEM2GedIQvoKuTQY75rJhUS3UGfko6ZaB
9LVp650VGuBggc5gKmSQGmPDTs0BGG3WW1SiViNJ35DnunpO7sSeo+of/teT
4KEgYSeFxi5/cD9U8L7u0x8d4qn8ent+f/BEONlOGcpyBPWBbdwr3UJkGOgr
PzcZdv6zAqrJ4YPLwD0Wym9kRC986lP/WZCmdR1AheFXmQOzY/mCRIjyh8SX
S4LYnAawQiXNoJhv79Gf2/1+Lu0d1BR7X2LjIvELtsXKHuhV0/lExbFUWK13
2ICXooeXpadjQAhYwPkr1sZq4MhkZc9h75C/aeGTwhsZmNXl56Rv+gEG3iqI
t660V4tbipzyARD4E29GIyBdQ0rkgxotqHP49vS/DYFcGk/8O+Z2eeX4Jj8A
n0hmAB5FffoMclXvKWJnTz+PkSOoi9Uqqqplt9+f5mZuMw+hUnfTSPUgoZfx
zTOknUnH20GUPUUHxVOHaEMiLeFy0+Us3JnB3LSXALV1RzjMZdeNvMxwYfrL
Z+ZkpDEiZX3jQhVSScBVLIptvgTpcLwO+JOsYjcm1oKIGP3aydHl0t/5fqJ0
gFhq6tP3Dh6IKORwwuU7MmF9ItTmQFkd2DI4zbsQfzn6NqCjfPDveWGUUmhC
FQTBUPcsUFfOzq0lY7pD3YFlucxACHQC7/QYkTq9/FJI+UU9wHv+b8XrROmG
ECyMPkaEw6xC5Nn2hahdhZYmz4utr0e2ZzUYVI0kQlHji0CHaTX3+90kOGmp
ZT3TAJ/XAB+LZmPUyv7Zno4X+FImxYWU4LxfjJZLI4oQf39EF8P86WKm7XV4
yjeqTjzHPKZRn/c4zXSX0bH1yVSQ3tlHBhDvF34P71nXTdwuRrkRLB22Q1fN
yWthAmeDhi6C8rNeqVMCo6YkBHGK4eopoj3vl2Jj3L2hP/GuMItPz51oErOt
g/2kXn5y1/ty7sEAQ1Bd4ZB9qIE9OfM+ylMbBZ0JqMHzVA/51UStw1f752DT
jCdRTAOZE3Ar1Ai+K0i+cQ6yb7BdT8QzIf7AsOgI9H1F/3GXlbpmHgAvPeG7
8c8wPg1S+dy4CdlMgXvL9H/yBeeh2JhhOv4ylr3GVLftAL/eHXQGli6u2Hdu
1vclQfvdOUjWxQZp0jwQyI0ksLwjJH3HzsHYvmoZ/9WjtX1fsnGbDNqR8SP9
MVlZnfFj5dxhyONQF0uNSPM4MFKIduUsM5VdXQoifcjkq1hGBkKxu/0PfgOU
L50L1Ea1aO1jVgSR3FZ9hb/oDSyZY45VJ6oHB6HZPcXqHEvBBbZcsPNuAb3r
S9c3u8wPy7511tebr0fJx/qMP6S6LEnLd1f/1vN/os2r+WtvPo/Dz2F29mgW
7dqm8QveWk3VohWqJH7qqHfwm+X3q70wPNFDhRHXTW9vISSGArE16THuHLtO
xZ2+jNmbwd99yu5myMzSISM7icqLfTHoWYE2zxN0WKySnsYI+nKx/M4GcAJ1
IRO2btyD/7WihK0sfPdIPGiZs29tErIlbHlNeoSYMQED1ncf87QSMMbfWEk1
oUd25EirQ04VxzXkiCs7/f5OwfL2zT47M1DXuPjC9s5uHUWgyGTVUjhM0EeP
j12wL7qkUcvT3dXgb+DxwVOHEonNQ9F+CJpsnKjAACwpPo/eNbCqxtF/ZNfI
pvsN8o2RZd7agKL34sC+UdAakXsHd2B+vrJjqUeQJjyf8BrN/FdpSCVKarZz
g9uKT6Doe2ILIsDObPIGbehBq9udfyxFsPAJ4lhUhFr/GD2rLOWvJZFC9VVr
B78Z63jCBwSa7QPeGqvqLgcl8Mn3y2OnxooWbsDQh2vZfP5qi1XAXEx8j5K0
rgVJFhWZinxCa65uvujYl8fLs+FTFOZ4pOWnlevhv7BPU5Brhs2gf9muT8iI
Kp7lsJOP3MJw1SygWhDP5DaTO5SE2hFXbzYoU/IMzEYj1tNY4q5jUvj8RFRw
rtullIzsLjDYbjMDkss4Ou9ZYfyHKNBFC5pJ8IqP3a+z/lZQnXkBxlVPKaV3
uAoguJG0sREUv4UtfTtlNdzAdUPnaUOTOlHSxidAtRvRY4TPaty0ykR2wdqn
RUGqfZ56foj/JDJ6+PLF5aZAv2Dl7ySF7lD13FCisl6JlXpj+ae5X7r9gzWL
06iFP1CEyIqX1qFiShvdxppxijn0n/h8kGnWHtCeHupG9oSdUBgHfqD0xxL6
E6dbjWFW5a9BPLWmnEzhpNFxBP6cptZJALTH82ucJxx65xcViBFQrryGcvdu
xpCUWrbeqyCH3f4OzZzKixAswyguGEdDDxew8CrjGpejMCbbXb7ZHGW301QW
MVWlmFzCML5Z17rs8//5f3gJPWDrh3fRDvpXCpulhA/isMQx1HjgrrhhD8J9
Ci6KSlfSFnai+ALSKKahe/SRIq4Ea7sqGu5XFHO+2fsTDAwa4gYcbfFrd00X
T5Msfq++FRNPJ5JLbH+mFNLy7iYU9htsIC4+dvqxX38KpmRKdtKnF3IMo0T3
aLL3JMj6ro8LMv4e+TPThRJGrcUw0u2oLKv+CkJvf0JineTlUA6VIqmC6L4t
CCf8NqSDjzqKC8Ix6vh19upgQGGXumcjv/H2suPzKGhIs/bS22yO3j/92iRv
fff8bbiawBiqa4Z1WTx7WEhJcxtOFKUv+1E8QujJj9gn7eRKInsLESVtxnl9
dVQ8F+FcrPO7JEpoeDH6zcHKbMT/5qO3uiAdI/jUKkHbIXn5ZP7xM/qodXmd
ZJ+O3rszzrXgjz3y9EX2m/Dl1/n3z8YQQR4UllrKhZslOZNMlb7TdhVF2e7f
Nirvs//s2lY6Ds0+5XJhj+RNvmsRzK098lKeb6TQuNjmaSM0KJLBSASBw8MV
CbIq9kUQD+4qxWCI5gbaPG3LmRGe+RseEG1EIDoZftWzhtceCzlWR5nlAlVF
8KtKI2xMxgnW+PhPs2FMZqGg3G8iQ+Ri073YWmWDn34hA+39l2LNKCkWfA4x
K9RSKa9+MQtbrN0F3sE4o/+88PTcP34IbxKmqtqcyxGPEvf9GnQXOSeGHaIG
R9ec1clnNpz5X8XSBj5NpCvLb3YOnDq2zXPrND6HlXCAk+8BX1ITZzya9Eup
cP5CmgjwUEeSgoeG6t+kvtxen3Y4ErEDMho7+oe8n2NopyzW22LvjgzRJkbr
rwUVUjaKCWg2b35oezzEBtwMPSaFi/9IbpMtefBXsUWXdWzwgRyvhAwzwf02
VbeGgN10ZhjBdYWw2gJjC8GnwLRSJvQr8dwBSH94tUwXcaDHuz4JMMxvUoBP
G9YqON+qetEhWZ3OdGjtVHI6MWqjxm94Kk53N/yAN2uSc7cvnUHd+1Ba+OXn
G9zbGgPw3x/zsgUHxlbnQgvXoY40wMqyy/nUhbRWEJfqiF2Yk6ZSKpaWhzbU
IAkpllhRcD1e3mstgxJLkItGjBsjYHurQBZmCV4NFzsqrDIfMA65X2LqFFky
LBstQwesWwZjQTi8BUX0ss1b7y3EWCtgCcXuQ6YGlJquqAUDUC3dYRpIAkqx
7+UUHRTlqqpPCfyajH+71dmBdBzbk+PsV7k4GR+AfL1euAu3V7dvVppNMWl7
bdbtpCYEZ43hUP5pXTuVF/694415YnMF2DzJq6EsSdrd4hmv2BEgOFnFwtAB
wYg+qaQpzo7guagV035wnY0CHMudsbyhYb0djLtut337Uu2QiH/sR6lWBA4t
b1SDtsxUKDxLEGL7N2xNjYYMQuSo8eOiI6Skx03Lz7gR4pUGI1yIxcvMd+Lk
NSwjenUlGG63kq5M+sddOADeMyRzWPerMZ5LQmAurPIBleYy7xreW6olTZqp
B+GrHcJ9W/IhLO2SkKdFrdK66oNooIyHEvhmlc85jqa1qDGXqcZn8Jf7e7RE
lTZeklBuKxgR1nFA9gBafOrgmur4Q3WuXiI2srRZmyTxrC2rDKkO7qApfgkK
QTqs57/OzglToKyg20lmb9KaLvyzPnC0A7k9OtUo50fOfzFtSxiVTEMlHDDg
rlYrwf7oa87fbO4GYWTjCNm1SZXoiPk5Mh5Lf0otOVLKGU6Ya919qx3V9x4Z
gRgiJ3aYGZPQzPn+MUzQIhIy/VaUEX1fOPapYsdh5tQVKTU0J118qK8Ffb7+
k/itTvkKj4DtM7OqSkwJ4kK6e6/pHNblKGkZru/YeQrihClDPcY9s8lunsbs
jiJqCdNESGijU647eC6X5Cu03TqYPawn4Kt7UuKlZOec4F7NIHFCfz4E/X4s
Ix2CkTl7sU47rhWIBBsPUtf/DQwpFDZlvtLpT1ii/71MORW4bPFacQ+Re7xO
/EzGCvWeKJEVewDtXzGS75Dv99lxKo9FS/CKdYUkjgLdjGpissakDkgpIqi7
dC/Th/oPBnbUd+Rz3swUoby0UgBdw0bx6gcoQHNHaFYlZE/1h6YYImLLj3X4
KuxzuYdic3HtwMWGzwY1GSjlyj0piPzeY1iNFwZ+bu40XgcPV4hBfNveHi2H
Slbx0xnfr3GXZkV+XJgBYLO/gpPLQa7K5NxOd1RneAF0l4j5LRolY4xclWDT
vwBHEuCqCXBHS6UlFrULr7LVi6HjmUuH4TbYfy9xA5mQlBb1KKgWKxxL1ZU5
9WVJTp/UMslgKHojbSaZI/gqIG5gozInU3jvAixzllnK1iJsNrZ24GqkanUm
7p1+ANP6xS9MEgsp6yXI5XYPBAu8VnkZTr5kAcq/2GmEMrgrv7IniHo5LIqH
xW3rMeGmuk0ygn8NXccXLidHft1Fw5zDSwV8o5TKsVULk6K34GXxkoTORnDB
SBIU8sdLsCdq/zCSFQgJGnbKI+5dh9OGD3GQEAIN8s/DkeU1Gh+I51LIUPmQ
WPG2VwVlwvH6JdfV0oRGyC7ZUxM9KM71wfqtI/F/d9BztzDzjBqHiL1POuAd
SZEVRRjy38c1+k6cSrSkn0ix57QUf1Jg9Um6fFfbtrlUXOJYvy6uKbjjl1lP
0GoOM4gyPf4deWR28VRpwISGMEw43GL6soBjsV6gYXmHW2k7We9mNHp4pFsQ
7ZG6rnuie65AJf5ahIn0Ylqw3SaQL2kR6zpBf4IySqsHVe0bV2zSWO4aVWIP
gDCEx+v7K7D/etPkh5D8obIjRa8A/bV420JegXNzvkqkhl3tAeUXfvP6mTp2
qp5zwKXYxaqLTalbBjA6zag8nkM1Yp93DW+riopm4mZeg2ppzV4m9u/OyWHE
F0rCC+C83vnssVLW7Bx4IPyW7KCTG0uvCJJkchrkdk+q7RWd6gUgDP7shiGR
yUJK5wiYEbmCI1ZVenR0XLa7qQYo8PE/UdpEo2RrQUDEDvQEdASWUOxGMWc1
85RpVwmc5rEXk45vYNSFPZ85saSZoL9zEb6IOvCRzJ7ojAEc0eLDDiLKt6gG
4SSy5FSwk4ySS8i0TI5L7YOrJR9LjtnOGwZqaCZgS7n8ivuezt2g50hOtFKA
Jtgk2fb8EkBG8XwCjU766QOQ8wV0Ue691guGdrdfO5+2VkuuU0ME5EEqmgxl
485WxUTnw+lRU5A8QGLqFkbXJoQaGGczb2MnsvVXexp4YZ+m9AgVoxcK/M8F
/MEErzFF3am5946Z0Ye1dBBwcZ1IEKXhum9aHcJt4XsiyEBZRm0TUPk1n2kb
NOpbBQrN3wDWuH4JmXzfuHMsT9AaJRMr6nHg5a1dRU7iqrvGIHexeGpvCWNM
YPDh6E2MY3nsVw8Hd3X4owgSQ68kS597PKsjrHNjVmWQsBXLSyDoTDT+Ud25
icndpsH83XxIy7Kc//V4RtzuroMHHqez6CGpaxv7WzROA6j51785vZCVFGzS
AxdaBJlLnh+BZO7MxDaIFFtIrM0rMF3NM4lL9K8I/Z6FJ11TYVS3qOl+OKEt
0w3Qfcke8iMP4iFt+rQDLBixpPwp6UHeVae7giZqcKIU8dokzSsATVZMyzEd
SV3D0PmZrsvljYGCWdO5zQyvLCGegKQyWmit+7AzdgxZYn3UeKVtAFG0SQuY
x1x9lYgTfnCDO5SLsJv7j2xOBszIrSRgBsa+RgNHx26WyO4Sgu9mmFMBfSIj
qvEho7X3/GnndR9uPLjmUb5uYbNQCFEA3romm875aCquzrpOkyUbWm+oH5uF
ArsqJZJBNI+kLkJ3dSVVIeKS0377PBA8rf3d8hO/j3lSCZTpgcDlJnM28ZSS
Vr/V9fC/dAZ/1SSS/HMaRbUMxIfo0UOP/aFjOkvk3Eo6kx0q8hFqrP3l5O8i
q8flIL7ouJbYqu1QA6oeltOkt9DscVsVNMzjCSDOEKoruF7YYNvcHEgp5Euh
DO/C2OiGnIJhwltdTG81LLvvVTxgP1acszA3eu5u98umCN096ZsbCngcV5HE
cDA12vBhLZZ+2Kx0I2V6BFWUerlrQqMjOGpcqeewiKQzNM66R6/WoVQYX+29
8eLmSkOQ4LdWkDtNlKLPrSEVCd1gVqiMKFN32wC8Siyx+X7rDkLOyQI0rmbc
86X66dQuzrhhRM9PEdxsAb49jB8mvazLNbRMZvNHyf30HqeY+b3anYFVREX7
07Fgh7cA8vfAJaHM+Li4aui1i6u2IlxfwJ8QJ3waetRq9UA71/JGr+YkVXxZ
uFYPPXh53k9k9YIr7aas3n/3MOGifJmUn10Ujo8r2xY3nUMbo3puzGvY6hjq
+4qb6a35uZ9Bx8NYfHKwz2oe8XPvi5X8QIEtE69320FizxOWAGsa8KTtzCGx
1P4e8mtHYN+ANna7fozn/HJB8RjymJSFneYf5F2IUK0Lx7sqiS40J154AY+2
AX48PmykhHd6cDIRV7BtODlMislFhi8zxUHR7mtPwoOi4eJWFyNJS97D3ZZ2
+FP2JylarrtZ3mbvGtmw4yZcoXCwsLD1TTD41Ljpi1HfO1mVO/EOT25tbSC/
fw2p5+68rMc8HT2PPgkYmz+sdQ+l/nP2Gcnla4Kx4DFbLnpKIxRI7BpFAMLe
H+STdE6v1TladsVDHr9NLoss5sHq+yMRTNgYjZ6IuHHiFjWSAxs8uj1LQzuc
JiGg6vJ4KnAl//zPSHK8TJvlWwaECmRLbApcGhJWOlP+O45x5EBnAXmAAsJh
eEivETCEM4f5Mj2vx9+li718UfihgA2WfVSBdLEKVMPL2YBwBRbMXk+kuK+q
dIGOMgmDvP1wsSyE2UfYPv9Kt7ZvdMS6WhI3LjbER+ccqUlGwv43rzpbAgqk
cOzoz1/77L4oZ/eifRfFR2/8nvsi4ClcEi1AzaS94Ue7hwXcfeejbG7ZYPI3
cM9uHLabBLTuYyR0juEe5MhLpJWRgxeYjCwrdJOLCcq3msVQAwHZlQhFsuV6
6A3xqUXq4dMmljYPlmVwgsCKr1by6RGC8LJ1Cxjphrq5WHZp2w87Zc9kBByC
xiR/zGWu2eMllV3ch87ynY7ot192SFobbkiWas0tAUwUrv7Ch6vSZWah1Dnp
mu+2y5trTPDUkFIBn9kUjaSsV2h2UQ39RL24H5BvgumS96dcm9+mg9UVu9Xb
glMTb8H/m8Jr/68EIzYdE5wm4dAhn61aQ18EtWjSZg4UkuGYgFhubAjATgrY
HbQWxbrP8NGT+lD4eDP1gUbJBM3LHJGes193fZvxH9TB+36IUL5wVpgh+rCy
VQIR2RRbpUOfkOmgOZaubOTZN6AR7Lg3DKPT5mlPcT/G5VW9uuWIDSRoepuu
F+gErYZYDulNI82NESCfg5CaNozg4vRPnRljVi/RQ1a7N1MnCtNcygb90S/V
mA+ov/X+jB/l5r7sqjpCS1QeKG1IsFQcXVmOV0p0DdaDeOka61Ex4cz2zG5x
kLZM1WCEWkChIdHi5znb7a+yMYa4EbvMGsVyr8gH6xTUBPqHsYtJe2QGwBSp
tHCBM+CmjYb2QqqIfjMk86CHFlaM8fi0khujZ51BPcbDuG5ohK6ExSjZ11+h
SsK6oEFV1wehXwOk+0dOI41PzXqAaxB6K3ZlEv02JIfzT7i6Wpy9v/SFzces
Ry2GICit3yorUBVfuG4eLMVFrvs8aJ8GcmaboVYegX2Frob0xirLvWrYNgBd
O4knjFJnlrPw9pH/wyPC+RMzVh0gl8y29n9edEOY0XW414WmkjsD5HtpQ453
+yNYncivNThOopFprYPYrNsLAjhgKJrZP5wXTrUog1LKk34glEZn/iwJR4nl
qOBBwaJ4XZs6Y46bMelBT5sPVNuCfPamdxJTUb6MRXxkr4p5lGR9cIryVD23
+IhWShlJ3qJjVQl8Old4/dqvOiyLJnlzGU9+28aGLLxp94CY2vgJ0LjcMtlH
3dB2h51SEsqrsvX9hRw46NgnHaxSxH+8orz+mKlDAiEHReBQsFMssOWSxUHi
hq2AX2uv1LLZuwnnCZc6OTGm90ch6EZPUci3SLNKnZprFjxTL0xftroxjd4y
2Ge+pHEMpE7hqoYZsYSzaIooBW/snI23xJxBSfQoYadr9StFzdNYk1NPLxEj
Ro4UEjQ+Neks7v2QYW0Uu61+0Rl3c8Mlsgba9higyu7dwEpnNRgogWo7j+EY
ujukmURMRY0HxJ0AMCFuxrJzlSbsAeGLzeNqFVVPSaHodW5dHfPl8BbaS5u7
c7OemneWCZY6peF94HLemHiiM8z3ovF8z0FtUBIs+Qi22F9i4U3im6wlp4AF
gr9M6sHu6EcyBLQ6Mm6l25cynHqi8QoVb/WcYH0GrTqOhbpjAptUGi9z3IiW
Qe9Rjq6X0d89pMHkM8wLN2dmSXTcZWRHxyjHJI5Yl9Okk2QSGdOoKfXz5BTE
AgRwjYTS5lxrMEU824vr46i5Thpr/drUSuUbwiEM90JmNRpmwtvRBd2cxrdQ
JOHJDszJzMDIohjIFI9vSqy8VyqRs4FMCK5y2sAGHY3Ltj19l1JVGhnHk01M
YK1f3qbqZtg5+9LT98owBfBPZ+o5azg8Px+7t6XmRsMpWLf/MJadQAd1p6CX
ejDzpXcV7+b2B75pXLW8m7MEZ1VOQSm+EHSm3w7RWGbOvG4XwJRQesJql9Ej
UVVejQ+MlwckgO/AyKyATagO3FK+DkXcgN68JyumYzCVV3mm5Dhl3j5X9Val
GJA1zGeTztPoutTznIMPGmAB+B6GrF2AvLTAkLSKrFRPWxTlbZ2SLLyBrqbo
8+/zPw8PILcyYT4jmPm0vKwJWItnD1FbAcTN0OCDs0/QjO1eA5aq7y52jeCv
5cjP11UjDa1tw6ZxdwuIWwHCa2/Letyj1drQFntYORIUZt0uUOnMYTlOvkmN
XUe4IbBvvYURaz+TENe9hBCA+XDWny5baMOWDwPfNRYYjtkBBZ055/i0pQdR
SDQVHCtWgxom9QREm+tF4DHg0gk0uEebpWnIjpk9DGvjzx6+GyghSyJCU1Cd
WSthz+UltHonu3g8BDY7RlgH92DeV0ZzsZ6ZoqlZ4i9XIbPOyWYJ2WM/WNaT
m61nU/j1iXkgL8qIJuImiToIM8L4ynEphwk9MgzAcq810KC4t0qWayhejF6E
HYbXuQHyTzMfYHF+zvKREANpTIFuh9rYk7yweD98J15mmVQTk2YBsKjo+SGD
NRC1g1Cvax1wVFO96NRORQfWq5ZMwphtH4byKv+vwr3ioNw+WT+bDBwfDz80
+KPrpBeei4RLS4VszuAnfaG1JeP0Mk2TgmNFaniqTLN0Xs+eLRe6FvDYltcf
7wUuQeEuXznjPRt3BV0Bq5hbDF5pYiNPpcpsdtdxZwAjfiwyTLlHxLSP0DWH
u1eqgO+Nar1pozSvdTd7PFA/3KJRPxWdNg8NEP5rjET8sJLsgWP29bD7Ff0G
NDh4WxlLxpr42Y4wwDz53sp5Kckhlml10XuC2f80LoB2doexjhHKypQCptCb
kE1oMuCEuGVLhDVlE/WPwN3hGxLiPFQohTcJxuYoD3AOSxtaZEmDjH2MHqkF
sqhYIy6Zv3O5KRnur9zq59gsWyoamPT4xpdbn9/xwcSln2BhwA6m22XYSNk7
h4nnifT8AFGuOwnbm/1mEShmhIGsmsXGy/slpDUKQ+fJJMYJr5Vru/4eU33h
Aju+D56iizIfr2SzPaFMZ7m2eF7RHFEek1Lf5weuw5kEQGOym6U5Pc1PMZjJ
J2svdG/4CXBZvLDrRpykNKixnTpPbdyPfHAry4lM8nMqSupMTkCR51x41X3H
BQktukf0/LGYQwLqmBVsj2+Fe0nZqYvJMGPZPkJkpMiebtkI3tmi34YsXa9e
dnBdAHyTpOppvR+FEhdwhRCf6tbbLCSLBNuz4GJMMoZ0tPeczsPMlmtJxlzK
HUVHmQc+q9slIUJ/HBLdo8kC7WCI/d1s4vpPl0Mef4r2b7EJk7DQyJiZJy33
MGmPft1cvbqER5M2uLea9XbWLjlvz4n3OanHIWJiuGbfSpcCGzWowC0RV1ty
YHTYSDzzliE00oN0f47lnhr8/tKI/FfTwvvG7epH+yWWWM8DhSWWVHs7uo4O
45zseQbZYSNVMoDHuMq+SNk11aJr4rmBxG3sSoxZsAe8J6MKQ5boTnenH1lJ
BrWuwPsyGQKQN+myX5XFmKX3z+mkkjjih78UWsrMEcJ/wpStZO0TePYnZF1q
pu9VyECusv0VTzSzsx4J5OqWV2fRBPzPmrruGDPbh3hMpvd+DV2v7vaN05Ms
boL4jS6qepE4i29nq2p+BGcvwOtQJNe8e+xNnr80uluo687sdpC+QGKq41VQ
X5Tf4p3GOvXrD/6RpClCsxSWuMAC4ULIqvwMrC3Z0K69DV4aUeFJu8vrKBjZ
uvlVjhuwQe0P8ZTgYGQTw1/f0qDl8qpXD+wWH6v4Zv+UvPt/rXnyRvvJ3kHs
nM03hCmyIn229xX0NcJwrNJafJJQDrNavrh8L+zway66JymD4eTxWbIuZ5KP
LmIC3YX0CDvNyicUxodudl2vstDV757KlDjhXeV8PUd05JgZXEvYwH3Ch8AJ
oVrQ3HMi8V8vW/g4a0TzcM9XABlYbdZja4ThH2UnUtyl3VKgUIfBoTtTqRBm
di1BK+J6EZ60xruq3i3eHEIqMhyme81tJ9LDZKVCJZ2wD4sVyir0LO+WK+2W
OB3AvEWOdIguIy55up5ui9rljtIrMoibzUfOBqT70AFWmnShL5bK1xeWqkDZ
qz3TuG1CmZivCGYXTDYIeVZB77uuEZprjUjgyxLL5Lq+2XwPMnA/V1nr2VYB
h8Z6zExZBb2RrrY9YLKerM5l5n+GsyiKtLbmR5DpxkFD/hhIavw9Sv8EbROc
WexBXH1Qt3yy2AkIvLciPUS9vVyGdlV6ZnSdv1APZkai16tUPhpOoTur49HC
SNKipuq39criYkS8YX8zf68SJfWbFteuzjdXoLwmlNqXLm9KcINYLZGb/WWn
XrAHIp7mX0Z3K0+lnzqUvwjsAvp+SwV1FKGyNngNQAqdO48EQuZjlb5JSnCy
YPw52a6J80ubkzgjkq5n4xKAVid6fljuJVO68CSJM5m3P55jrIG+ul6/D26U
yvbPXghA2AebfziQ8U5ySz903oTX8cAzGMxPAB6W5MrHye/yd31R3XQPwvIb
UT+WaKFxB1o3rR5/YM7QLS7SOyvY5MYa4r6WJKaCfPNEL2MCJos9+ApO7YXu
eaPtrntSZrz3PuV8KJQTDUKplU1kspKy932AngVAJuaPLd9Xep/VoLwIwgKJ
O0FkEpftjrpAjnDraWeAh51bvA0toi9uNC2pPsr0Azrvd+v6IrXcmrf7X1JQ
Ymb1nIGGkp2H9KyRMe7dGbHsv2TRXTNsLWppeTCNWCnPQnogAN7GWY0UvLCC
gcTSEV0HFSuCinwEXrZurNgRB4g3Qnhwg97WHW57joB4eppdt+2NW0Uxiaql
nFbVbaVia/sbBgbo49mj+vDWGmKXaRLjT5Fkt2XjEJf3hp0qSDZr31lxvYil
Al9v3gpSe6pVw+7byfOe2j0FOLFQj3Y4qfc+fTeZ1GNW8cIh1HqgaYL+8G9N
NlDAWdakNJEbHU9GpnnqBTX/7y28TZ6PhmTSkWo+4dhitkR4psxu3cx0gG9j
+6G2sE2TJ1FB4QXth0fbKARSKj0ybOPNKUJy4CyN9RjTbQl6n48MXbiK8hKK
bgC61Is3SeCFWL+L2vY7v6yOOrIWQhAYiz8IRf5NxnNqvhgimaRzLBLkpuOX
tU21Iv4TbNx0ot0YAO5KKxVmpts9Vhk7WgQkfq1Ee2PQXHpEgBVIWYi4RHbV
JFX/jc44M7/9IAtRLy5LtXaObfw/gBg/eTVDZ0lFMeKJSoNkVg0AXNfptjLv
nZTMTOZ7huqsK4e1OElNcU5M2BkmYdB6F00+CmWmo1Jik5W/bJEvKezFVwL1
2wYfr48Nz+6fwzeIDUei7K/J69Y4Zc1EUozryr0qBTAwYcMUNPdrY4iASZv/
xRCXT4UjhG7QpK454dWU7oFdz45cf1lPrmt2A/m4EGCM4/plLg7oJMa7dhi3
r5vHaCdO7gYRo7pvn6M6Ivi+aXHoOAFPnk7U9xbTS9t8B1aq70LsXMjMT9AD
8Y2lMnndTLKVNeaAFC2iUaSVGKWt47mW2TUgzoqA4joc455Gg1PrnE05Unlp
RnDokNW4lMhfelDkrLAz2+wS5wt2zB3b03wvspXhU8u5EqI5v7TIzNFoumy7
7/WYnNs3e0nds8LVT789uu1pYGouYTjfeW4KMNFSPDbPmc0Fp4r5RcaWJr8n
trd4USew/UNXwSIwqTv6CjqLGNcCX1Pglp6929Nn68p6agWHditOjKth9rvY
3xTvAoGDoRd17GKJsXyXMsoFVBFOOhLNVeu/6EM0peSNT6QVytj7SCu3prMt
gyr2MGL8D6WsFAK3dGfBJSHYuwi8WZmqOpcXT9bQBCtndWgiBkQM7OQHYn8T
DmIceTbPlghwESyKA5pYEkM1WMunmEiKkaC7cBL8lsQOeGjB+wu3HHmP3mv/
mQgwSSJC+Kb/u384wU/MmC0CgisEQxGefkbWTsrWqL3bbIIm/vqYhHQvhvzK
aI2rS96ExbLriSVu0jRQpGE3zMXudxwnBh1RenDj90J3UhDfwnk0yVVn8r0L
uh0eeHs1E2LzkuNkyGtqKUSKfQ1JcnCAiF0cZBpsvWMD8luguk6iYoekMrOn
KCyTjouNZbxi6BbjrGf6QLTNT7NA3TQJ5NnYKdYHAvPizE1g2nlVi+UuiDSu
3sGvxwCKSW9xiGAUp5SKjjXHZMoTqFerSqhz+Fin37l7YMp/jmsteaQ7QVmE
s126AoKnBR+1MGQKbO+HVNYrrIxvbf1KR1saEcilccdaptgC1WwQzqWotavv
4BzB4kQp687Pvh3aJQ9TAK6OQKS/CXnYuRSwZfyTWWacFShccdY/cbREqpir
at7homGSArykqKkU9LlTlzLk7fvM0IYbYUix2qS+yg1aw/tkiJXDch2SSK+y
nIcR/jyk3oiI2mbkRcfeICnR2SP9icZ4+KibRCLL/JG3cGWeEiNQ3/5em1Ay
/9NhBCiYz8ozb3NguYZ17xZ2cLFkOUCL+EqjeltBsSFmCX43WWwfPIY1Q4jn
uYL/NYPEv+1hkBxKDd4r/tOEpyzUIJD37hI+UKAWHwgreqbTQJVQPZmz25mh
AhE2bKn7AzEHO4/8ImtpuH7hI0o6Ghlt1WpoOUbpvoA6vy0l9AUmAGWWPrB8
Qb5XC+N9d02iK7tr4p08WhlcjybLn+/XQhOs4Z1YTZbQV0gU2kJprl69kMbz
8HaEkoFzlxnEpvelzaHhZs3CMYbvSkMkFg7mgYmioNBk4ocWZ4TGmj1dMsuD
2ow4mPgWliU0HrhYmVqF/QE8xW0XFfwgEfP/Luns9Phl8ms+Av4m+OGdaKcX
/+MoWxxXzvNJQdZx+IDOKUwpigpavbPDjcTVdahJg1YAbc8ibeLHpp0cz393
HjvMPLHQH//eg98+bmrb/jgfBmPkEtQ3KAuQ4WfB3Jt28k0ddBi3k+O6rVkq
n0w9mpxEP/T+q5A8Yig8DP0Dh/FZfhdLfkFGJQbZJN9O297bqafdgyDQvrvY
MDr1apbctZdRSiEenml88B0h+bzwBihZUtDm/nY1Lh77Cn6o8W/fzAKtuN2M
+iVmRN9IE9EWuxcNLmCKXDQdTf/g+rlFWI7d8EmoPwYhDtinogqnhSq+KADb
yCfG7kE+hM2K/PHIoXN/exwReldOiO+QxgK7RrEDThLtUTytsQPDrku+LBjg
MDqL9EABmVYdIYWhif13e3z70T7qY0jEFPVyaTQ+DMyjxM7G1oXJSd67EweP
Hvkh2vxT401LdfpX0PRXHeBEanLxltV1FzoUh9Qma1QY6hC7GqHuNfJ7koi9
fObswmcuP6IaAzAr4DpQqKpdxltt2t4/ZCbVaLIT0GxXh+XH4RWYzy8TpQdG
xYAKlBhXLT8aPsyrCu1tfTxMawN6a1Xq483OFYU+fUH3LY7Br/MLZZfkOM4C
DKNlLTvZ/ZNBDLZX7u581Rki3jhjs6AMeDBVcAukgOXA4P6JoUOCM71Vzfed
jZczGpcDgPk0AOBzG68F/TRNq5MmrRC6pyPfuvyfu0D8lnO1JCeoqlI0G/Bq
oPj64WgnYGUuu33ej5V6ZjIYy8aGie1SRItQS3Jh3VztV+losBLBPPX6np9/
Zxf86CYyd1LaehrHAWH0o30vQwULJoZiW7DUNh1gjHtltbVUUla/pc3DAsDa
QEVF0LBaMkiw/Gre6MvG1MbnBncQD5AsjZZUNEctQz7tiL0ayQrwH/yMtPMZ
7U1n1NrZsJtT29fTa8YSlSuw+BdRlB7rW47tyVo62NeK4AMUan3lqnUltl55
WJoV57EAJG5YQhQI2FQBrvHuQhrZOxiGGhmdesOcbEMANMVwuEyA4rO364LT
ONoD7pOZN2u1Y3v3f8Wa+0KtryHtkbc99Cp9Y9mOCEl2sTSOlNnIF1354jqb
9QHfmS4v5mozb9kIYe4wISXeRM4D0Ehqa/GB/Xr8fmAU63Rryoyh94hhbshW
RdffJHrothEZIavhtQKwSfHjlvgRF7LJYXrdU0tfnggpbXgkpVos41LmtYyv
sj/o4JZJY1Ld+xXdGycvri+4BkxiwosV7niVbtx3LRH+ThWSk7Neunq7W+by
arpe4v1xsVZ7iqZz9Nn7gTNvZ5LHjEyjEb6a9QJnl6xrFfOX9UIN72DGfdm0
/lHY+uzTEw22YQWmqsktrM+5rmJ6TlRRgxWHkC0LZTGaXKETWs+yH8v0Pzo7
mMuNG6vE45htGrOP/YXYQClWmPwcujTBd1RszD3uc1RHUj9QRRTR2d2Nt72d
sfr2aYKQ0mTsY6CxN1wwjJrRdcb2dMcU72g+D2Go+8R7mnAU2s+TMyMJoMIF
0dyk+Ex07uL4bY2ERxQxyfU2GaKmrtwCKkhpjdE9NXVrB8j4gSOHUw1NiKTI
/uok0vLPMkXaKGAyvB9EtOJ/OttHEG1c76qaONHKruqxAZGSItV0Hs7J9s3m
ReaUtzq/TEIZ/4NLnFbKZl0mywzwgsMwmeJYMrFkB4S9T1MFsjKHxjoc5LGo
oi4Sp0PJnVkVhaWefIUZY1RyRUKvUqulo5v9Dpek6ZcFE1EybSQ1zhbPl31Y
W500MG+shQCvPUOmrnwgqmjbjqXB99hr0N+TrteSXGxPmtgUJwmxokRD9T+P
+E9C9EYgRMVdc5rVjI3RgYCipEeCfyj4xW7TZS8TiCeANPHTq2gBDc8itoIN
nKZqkqaO+VGkF3lIuq2Vctcu+r2Ngz3coF8d0zi2RTLHk8WitjUIzvF1x5C2
QIO/2GPjEnraCeF+q2I3WHXen0RQdCjsFYjnwQsMThXX5TdWfG/dAerUJzhH
pXthoWpcbPnGNoVeT3KKuLSiFFPORXGg3PJ3nlQNipQQx8BH8bPDTozLqTFC
s/a4nxrGsMTzw8+h5FOjr9hVSLUU+A3wSvESjiXS4ypNWkGavyPfo2/IMoVC
dYf+P9ItZXIrySqkmmSGT1x/bTqcnHLX77+Q7r77b0oo4pd+VLFo4DWIccie
Xle/K/p4i4wkMjT7DS4yk+eUEoNmT9QsPgNL33mAZtjEHcFd2/ljlfUUQ+k4
cWjOey6K0sWr5zH4wqIkuTTheNX0udTFCP+jCk3QmOB932ilzsg4a0+H/P4f
bvkqOpcbFNzJ2qCqaLlaXtCYynyg7uIE2749nCPzKEbtZWFLbGEkeAOFu9Gl
dqn5Mw+D8mcfY0jC9+rr6ZMQ8tFWTbzQbX1Kvwtoq69Xjg0NJSlfR/P0HF25
z58NtEhTamKwc0G/ug2DmUwSs1k1imRpOEmBHTCb2Yavdq+tJMUOqTCwISlH
l2OgNo7GcWoEAn84Kwn3nF4jLrhtl5B/iUFWvdwd0W5rx61SrmmSGXQjia37
dh+zoMA/4x4Qqyj2y+9iVUbgB/6HPW6xlBBbanLwvvHQPB70zLS+W2iycpaA
0EgbZYeAXNxdo3g9oOp/y9PpjrGicRhEuapqKqrvBGfDx3OPfvxGmfS7CCZo
sPA5CHCDSlLt2raVO2bbejPmlW2c59b9k/XxMAFZZfcdcw9j7L2QRH1z5EOG
t/t0CJDduB07UBB7oDEe8IO/Bj4TUiFqU+vAGPAixJE1EkF+V7KjJOIAGTYF
uhrxCtxuGdFdtTh77XSRGVmwycUWwduInFW6o2Tu9Vw+lmqZ5ohnebj6KH38
yTm5avQZjdBO9eKA8v5kxxUZgSqq63cnslr4dRQBh0fPTd9IETQiW+Mhw3mt
MtGb6iYwR41uXkf6iAwmIRxtgfMqQwjICRoMAmR6fI9wBULCCy9qu0A3Mgw1
huF1GITGKUsDFmOoloQuzPaL/lgIjV1CMZW/Y1M+48SX/mMrYnNJq/xLCpJi
whw/r5dMlgKrpy9sqlatmAHURMR00uBNduf3ItBIciOr8kYGEur7zUkF8UeM
j9ml1x95CZ4nWI3QcSB1ATEnfNlFXrxyh4dsEtbahTOQVSBgEO5c/sb0VglB
KfcruUe7/C67Fn+RWiOM2TPRcr3f4PBiM6VIda0W9Zs/l8WQhfT/OkP3bcxw
cHa8FtA3LSbvW+yqptTChlMgD1j7m57at2+wBDPYoYdy74iXtEF1qqqJFuA3
tp8X0fW6eFB4SxIbcCJouu5fBQ1nh9rPJgMhr4uMfdLrlk+9dY/OByMHefGH
baTu8INQEQx4weCOYu7wuilLL+nZh39YFLCoKuBreJ1UmnWvdZqjJnzlW+A9
OqmprsGOy4fIOfZaB2SGOdzhUFQ99p0U1NfF+A3uQrpxrA/3lLAWio2Hk3hn
0zZTmyKMzicl9U3XNQ1A9In/IK6stP2VhgcBs7iNW1ZhbKSR9qA6NWDTO97s
IfCLwIlA14xstW4cEUFAZNbvzGtFOOMsOlU6T4kKudk7J8qw5WgBwVks+eMW
V1IyHxeDzFXtX1mcR4f3DdCA71xZtP2rDuYftDj/+z3fnalkgRfFVAauhfAl
t71AcT+xS7UEqCCAzJFuozYaBbQULd0PpA/+KTTQYghP+ANoP4G7pblbChJv
ATpT/pgBguiopj8S7uUUt+rxHHpebV2kWQ3nufsTGhRslYEDaGOh8oSoIRDZ
XOhv/D3rstptNpc2DU7z4YH2ri6swVVu9o/OBD0K/Va/WarJDMK1s+X5iTFX
epUr7blolW0CBd42ssHBrOrHpwdsy+Z2AGaxaBIHICCp8qR9qYy3jSy5aowM
b4elOonAvp9BMycUVbHCP0r4l3f+pnUMv+b3wVFZyLjiRRnWMEoInkXZRGwq
S5TgCzA6DhCEHAX/qIE8JDOmuwCwaxF00Nza9FNA6Y+D3Am2s4JnZtQ/XFUe
HYBNoMVX5AMa1XQbwfZxoKmcAcL78EJbDic9Gj7BYsICxUDwNpDMQp+BkxVW
gUWly22Kc79oGN95ey6erL4+ysWRjS+oJSPFDM7vXZ/5W7xiI4WJCP+mvCaz
UQ37TyT/9FPITKN85vh6f+nAMRBak/4fjR8k2Y+0+KWJymPP0hQzwXuwepBr
Q3R1Yv+y3eWv0+tSBYTeXBsGdhZQuYqF5TuFB+q/bSNMj9Z2K6rdBNJIeWCw
VNCfEAvaeCQ/hiBg66pBP7q1/vmnJya7n8S554eLh6TKTMTVzn+DHCDk8rTv
Ct6vHSjrZNEkZNlrhOzUPpsb3iy3x6InECMOjnqGxj3dUKCac86Qc4YMjyuZ
HGOF6k5SFEgPBxPluXB/RrwSDRWPcQAmtyJZD7ri8PgWy94EB2S7Bk1FpKVI
v5e+uWUsR5VtUSiu95/rjIDC3WAQVJ1Cccb7JBy2ERphG8TsWs2aXpL8LQuh
udgQpe0RD/zAOYVw98Zpi7cIbMWTbh2JAsxU/tjZSY0vosnFi8mti7zvurGy
F9ZLU1Dm1dCwXbe9CbKiPEea2K54g74FIwsWA37HX3cwWUd69Pn5rhGdtjA9
FXgVMTLzdWUkcDvo2fGdr8kgdmyGM1ZpoK1xF9c9NWuMIDZpE0PgBj6Aq72J
pul/3uSGrUWLA9lmj5VitSqJio1gKBetcGnZHhoQIeb259jAs+Mo+vmy3tI8
DAbJd4CMDtojGofIh75MF8kMqt4wbuvPLK35COsfckrnxLrXDbF9YNfaZu8E
K7cGBet6WY4hl1Fv7cfux+PAIdlhRbo1h6uHqZZELzaja1lIwBMlCtJFSkbH
cKDkhcuYSVtzpgKAb77yC49kolgT62GNBAOjjF5b4IZymQw+ezD8tst3yA9v
WOtR/XYgMDqbvOzqi2k1JGo20kH4/2msOXs65tNVKtJstVPsAT9Chc3WeFlL
uv0bcAVKzmfZAVDAHiR5xMP6sWHWGmNGf0dZ3Jfx4adJfNGJLSEr5pXhiedI
lqUKdDCVDYsc+yIAnJJUmv/92XxpQ8br392DYkO8nBYAoIZXc6Fce99ecn32
xy+jSVRcoWVPPsdrvj3bFCyQfm5lp2rFWmFt5CMSEeSrmuRGSTHdmqA0/c9w
zaHrHG4AAK3eQ5iGqpFeX+NwOoe8hiCvCz7aBfVKJ4E+bGKClGEacTZoVh1Q
HGJtwDoh+A9kNloa4cX5dJPq4WWv3eLY1+re5eQBdZ3nqaJ01H7DjSMT6K/A
fpkFJSA1mVIC9whGQiA2VaJttAd45DkdqGJNQjSuByO9L2mvjeCh31X/r1EO
kI7rv025sDCe6hOJV5SSO+JkX1/Ef8oT7OmfKxw0WAt8XieOQU9h5+ZGFm6D
zpwW4kMOPuhcTNVGNrMr6mpo8rXrryy557WPw95DPPhG8M7ZGUjFZMMTYMdj
J21Q+M5cLtyAOO+29/zeL2cEBbGZ61JkezxC53IGQki2DBRNKadXVrc/f2F4
uLI1xvpuO7qTxr9EfO+6tHdHGS/WXHQZx1HJ0Ts1Nuh+1+5Inh2ES1szAMGW
MoC6di5hRPoUlCu6HgOekhzEJ1J/6MTh8gXck911Um4vOvRI9iH5HFBhc+1M
SbPmH5DHQarRSC+eV/TvdAVtbqSJk/S1lu5rGLmWL1jE2itC+aPdSGnywb8i
M3IylQfClBjnqhbM2/y1EHNSs/NZqrbJVqGJiakDGCztO472vcSQsn+K0uu/
8GGFh1524Qj+xuPBUHgc14RhC2Cmnr4V49xzePU/onlJOxI7er2QjTJ9f/3G
HcCC/2WZxTU9Gg1Cn+6N5oI+kC4hhFpw3wQvyUj2k+teriUaay53Pu42nMsg
I/X42tlBDGHmiT7cRSv1+rCtRu4xRPR5XNpepOSPYIr92H6RBJdtnZeb2Z7m
OTflethpHRf9IGMmVSSEe5DOiy+wL6rA4qG2BGgGPt2Z1yAFoLellAp4pCv5
mUQ4pLMLaeBlBzU704JxKp0+4pJvthunoGgd6WUUefdV9JRD91yCTLOc4Cl4
zySnctaEz133LP4fFJmQ/58+WE4sR8MkQcoB3N22bjH0Flt8XNhJd+Kj+uqb
ELZvFVNHtVMdsUcgwpTXdI7E0+JgLWSSoYtiITwIdofX1LkkPcNqv14MsXLR
cymY3T1TmFIS5ztm2ERRgkSiOIFFHVtJH3Nf1YSrcsC5T5+mSIG+AQTej6x0
f9waGZloG+pCD8vptXa4TMILQa7F9+FGeGozQrnpe1RUhjZ8Uv11Dii+TlCo
1U4Qufu2H8UihVPxC7KzN1+PhDQ0F3QmsXMxEGLg57ucyxauyIBNxS0GRJck
NthoHC9Kuj+Upwx6dZJbTe7PYkjuhOqCCJCWDYL1upcxO7A54ACkonPdLoHC
pSAnX3brNPRRTq/Fl/0opBXplc65FVKhvshJkvOIRLGVdk5Pi9UD2RfOh7qO
48QFI7NQlZZEwsd7Z4dX8V+d5otvC8sCu/g1pDoF3TqGEfpyf/DMBcu6PapR
K54+YJ7rIt66hRxCVVhjfgyM0wZfR1wP2R1pK2XMX9WzLj0RYxec9LKhnRfo
tU9GInjXSKfUWQiinkFUbSRtNgnp6kqHfe7sY+kdP8Si8IhN3ZFNNEDOZjrm
/DI48lc0Im+Kopv2gqEFPuVThAL8MKSBB39395SsLeN+K59aOSbr+SK4D1D7
3Ciyj1go8l7fXErBeZLR+zrImOo+3wzY7uS4+Cbx7MuRma9xzn3s8isYJrBG
wAoGEkn1I6d+5ed7AQ66Hxm7YpAfPiIc2MFR4aW9+4eS2vqQK2oi32E57wvd
639bEg8Pihe5mI2lJXY4Taj1jjB1eXAeg01dtBE+G7/dIHN3K1V8CCy5yd8B
L50BZqqzvttGfxJPS2x4M+3Jo/bJSOQDJ6orZl81ACfl9hpG8enLPAARwbfd
MVp3HuoLgODGaQrLKNNSASY77IGDu07ElM5bieBWjfOpCOci8sjqa8rX7WXH
XHuHVPgR3dKUJxLxOAaRCgz8lkwzY2bstNike//fM1E79iITtTFitIlwMQsi
pGCrs6UlSNRKIcsHVdNX/B26LXMTxTsHr4GJHrN/CfxoEAqtnkl6V+ICeME5
0RZ2pA/IrOfIBsjAHgVXBTbvCIUkkpGOcK8MUInmPG5NEIVj+4hP/u1nsIOl
i7a4owuK2q359arCPIALFLYs+JUYlg9oug6Sey2Pm/0H3Vpy68ycp2UqkQms
YSnrjrfmVxZMF5n1yOC2JNeQDrDlxIm4qz7cVQ7T2PX14Sv7MwG6i9WBfON+
tggQPhnLZjFV6wWrX8+2Jr0n2BYlncB5RlB8nlKPdwsf2d8qyY5GIkcgZmfd
B7wuYjULErtfdjJPqTAknHUAsX90kUWLUPkrfXVoO22JDmYYFeFWnh63adf2
/eVVSWpcZ89WSI2cZaVF4sTah8Tc+8am/Cd3ppgC8UpinlAhMQsOo0tZwvQv
2ZbNOAb60y9X5UNvr5ZCp/wc0pPwobJl5Gn6tQe4VuofKmBDLsFJbnqcmCVc
TUCXkmUsQiD2z4s2OfH5+yMR8PKXhOX2UPT485E+Lo1tuNf67bXDwl+F7UeJ
GeiStsmMojgswhvJ0TlJkuAIqQs5r3sWPVqR5hOeVEOgL8gGzPXprozinZ6P
vCLbI8b8CIrdvMrBBZbAkV07LiVKDju6/Qj+Aec5Vb0pGjMb4gK/+yc4vD5k
u6NMg6WXzu0OJ1cWzqTvwuvbCjY3CffiHZ4AL+syi2ly1FylICbcDrdEbPz/
siQ+HiDbVE9fx9AXJYUWyDMiAvxVeHiMnRIzkN4gM6AaL0nBh3Y+J3qXzAzK
PNPPZ06SblMrqgoY8OTzjIRIKUcSvIjUjEa2YsThrDcB/29b0oebynUU8l4o
j9TBcr3/yWkhbImrJv4bk3ebtiVQ8OteLlWQm5jb2y7c2TSMuGhGYb+3Gmku
zxxZz4ZJvPRCY+Lzz92XGejsEKOrHykgVTGsrdykjsX2fUz/Wk+JB97507PT
Dwds2Hm2mLuLZNGY6cHDAvoIKO0HGqAQNAWLq/GRS9r2BhBohmU8h7nK2Mth
R3sqFcohmsPKOvU7ud8rbEp6NJ0rs/TwuUfHGyf0OUJKcznCiWYfpjF5QxGe
Veg9rKh6tNh4p1x/+O+RA/nP2abOtScoxy9/dipTQoaOsZHOwUDKrTj4R5Uw
+b8p3VEXsxFwFf5xbFJ+A9iWHvpY//dG54LuJnudZgDJ00pGFNH9SeKGX0FH
yugdcLz4TCmTSHaD42m7lm4q76OhS51eBLVwCTIVgcmdjrdGmYSmJ6R5BEyc
iz/CYSZpFAIi42ISZ6LKdpXyiotzV6dQlarCLkGn2ueBbFOA/uUMju/RYOMz
nOa6DRGCkW4Au6iKLzyFyRFaao6mMEzIvbNRXCgqbVaT7aBdxippPRL5Gi/s
8jhMonfMp7xf+ros1mDOPFTEQR1mnE6FLqOZ30eo0I/fgkxAeF3vmMbIljxI
ak1AzQwrkPtWMoc6r7jpxVDnI7uwNnjVMOFtU99ykca5UCcO0I8zh4G/seKY
ikjCb6K1nxH6dir8WLQOdaU0uVbIA9RwVB4iOpxEJ2z2l4AwKOHVvnQL5Q3P
GAhgNxBWFx5nZ7vsHw/WVGHn0/b6//BcDB/sJATjzM35LCvNrjSFu5M/Bopi
wEZB21GLMKlDlqGD28V6Cpw3vPXPOopQgYbwCvHAc2wKOBqFX40X9xwcOw44
6RSPEL6FdsgR1wzQ7WHEP+aFvjA2MRpCm4WsGNheldZp4900pfVcdWnksIxd
QTIAORRKfVTRBXHTVvOWqC6/oDWP5+Rtk9fpsBLLXjQ4hIGg/hUuYjWEz1nW
OXCS5cwetWlgDZDvtW2w/hS5c62fPRCnnjOo77ucTeLLN7iUJD9NUGmBbi92
0JlwzKJSVmnA4+z2sR3mVGDzIczJFjzWRRXInSiyFsoe2kxtQ+Fc0u9sSp8Q
oRS9oHMbpJdc/ZO0j+BjZ0bLSJ8iE5CyGr7xXDhmimYeTee3jWBkxN1vE6Zk
ekYZjkxrj5T6EiAIMB8R7cnwehqraYRVY1oX5UU+f3YgotbKC6wpFeQ2I0QR
x46UJK9/b2r222yyxdi+cYSR9ljd/Vx3vUBsh/f6kRsor9eQramiIxLW5WXt
F0A9Ze/Pr0cZZQSMw0Hai+/S4iaEl9S8qVj+Xz9R4HA7f0pUoCpxDU7LojX5
nmfqrzN6iFvFU1fe7O60qkx78HtIz7xbySzRwfqjlqhJutrtHLOxq9GNCcPK
8bVUAywbPAExUMuL9iCHnw2d0Q2sE4lACW9Vc3vbn9B8G2C8ain1h3hNCLu/
BY4EEkgIiDunm4NlUyVRyWF4FogOyrztObotFccFtzVF8mr1e1SxQcJDJ7Qo
amdXpX0uddHsAG+jiTbxMUEy1xD0t4xKueWWb233dn3V2CnCU72K3ah+XPCV
kpcLxXJnDh/i7nyOqPmPUZWQWJTMVM1mT0h+DJBshZCYNfU1EBhd1lYeIQHW
gwrAokggUgmBwrjtyHsmojFWZuz8Az+aru9SU9p0Bm1Zw4hbek9P4UGSROfa
vH+UO1nRKv/AesS6+0PoWLoAlP6l6/bsMPiyDpm5uGezsSezl4WwxyynzhVC
VnQ9c003vzrmZLe3yElAzi0WMeqlpEGX4prsWZk+9EMMF1/fgmZsdBXFWALZ
MVFA3i9mYDKwTUWRHpTF7LfeRs+ihAxPsOFHFGK4x7dOPtWhCLUVcqXxe9k7
WbbdZb48VvvNIffU4wZgeuQa5s09LlEz3xAJ/Q+sJ7aTDNKaP1Dd9YuRE1ki
527s1tEddVUT0I9tGLTicTPn/y0WoFwPqU+jq9GAgd52HMhxwsCeC8Qzn4WC
w9KS0kmwdbunYd9JnPnoBoZnU4DFxIJQb/5VjXscCZFo6tOIIWVaBgyFrzaN
t0U3W01p+wGP72hB4bhyaiXHnucVwPKmJNOnYheYjpaWopVbS3fo9ebKKe36
sExbjzPqQTV2np+NXvOPk2nCw3NvN4kqsMHdXf9Wf+gWg5vwpI3dtGenew3J
F1aEu4j+zl6T8E4rpIWNghzsVa3eCv/F53GN2mE6IfZiZvd15GQ8jywb3hna
ULLk3op+ol/W8sonreuL6U7xrMIJn6Ve+tvDaqaZj5lFLTH6cL2dZmKbK66T
ypOjkqX6M8O4p/fA+3q/iXYnsNUcz/UxoTLz3bsKwobXpVXtJAMPR/b4p3yZ
m1dGKAWGFF8APk0cIL5ymeKq6C6ERBg1btwsNKJ9936i2PIcCEOESX/KwDaT
iyrpQqcbfPYdwdlGCjr/hGDoWl7gDkVK+MBNA14qq2Cl7xg1Ba1KqcHVROG3
KuvcHz0j6fXl1cfibd3H4uodCyO9pz3f4D6xaNg54mmVbDGMrEPxFx7UubdP
xhiYkeguNRZqUj+A5ZQxGx0RkrSteRs5WpWbWDJszEJYRoZqwRjbTKs4Ax8B
FovDp6q8FV8C0FagGtQ6ypXAVuE3ibuW4mJCryeLsqnCEvFsU+uje1Sz1B+f
04DUGmbP5NPtIIy8+D0AESNQbMtRlNfyKJzLnQ8WSJa96jJDj07fqmuBvNQM
GNIbbORFCupAm2lCl1WbhzM6TiMIhRrfzIFo6R20mmCGukV0tL7onHnfO5iz
32x5Ks12+UjByR1xe4JxSlLqspn0oEINY2AgLW7lrDNMZ3VZobcXqnWaAkxV
JEzCS+ZH13TTn4A7NA2/y8kXRN/wTm95pb18QTNrF3XGZnGV3omTxMYFHvim
nj/yqz/zdEyot8DzKBVyFkWVkkhevEo40c/YsRSuzmHPLm1ZirogSYdjufk/
m5044XurQGDwf8GrxLg979Wk2vbbQcPwSUpXjrb+2Ned8qHHchFLxJOmdO0R
p/81oPkJtVJzq8HDQtf8oR+SjZ8DvVjEEGfFvx7poZ7opoqd3FXrRjawV2gi
R317GUUjoiUApSKrVRebmMHqAh9Mk+GGo0YtsvJUjmTwu2kYGtdvc0A5qZLS
T/XptiXdc/NiHz7AdX5rAOolws6mCIy3MFpe3Q0D2bLKul8Bk9dd83L2lPwG
2R/VX4ttCEpSSkBXQEuiiNQycWlR4+cLuedkgHyT9G/94BIpueAJaXjgis8/
6YRIuCfjzYyjJplNCe4G1HMNciNz6Wps5Rwi4oy3Wr1V+41cLKT52f0pfvC6
T5DkJgDhcXbbJs6cn2KKyCtxv5x8K+TUxcLW3QjhJRmyql+VpAqIqeBcYmlQ
SB3iG06OKppDBw4AFd8MhImRxoOCd04EUMv70+EEW/t7A+3Sxxo/g8yARL16
NkGUGV+VncsunUjP8bX53z8S5Z4ungkO5IcCbcqeyOGtvYHk05kXPbEq8ok3
LTttfi8l2TaMMabpaUJ7/DcpTkKmsTAwQqvH8mI3x7C1/g1/0MlO+d6t4Vjr
A3vNyp1Bi307HdWPf2ZdqWaqenegyVSFnmllj8aQCUIwSDdDkD9aN9ibtZZE
N7GMqA73CUFecWxQcVLszP+J1D3GzYncFQ8Rcj3UHLm+saQMG7IzlGUCDoRa
WacT4CK0nmvo2lfTuvrmZn6E2A4wwssu6Zc0NXpAW9xR06LpGGhtovJhPXlr
gWjmosSaMWEgo873+DuZJ2NonC9XkFJ1uKPLvvnY9tT77DdAsJ6AaLyaOgDU
SlFVlV+TZUtEPKKzvso7GwdoK41Y4DX5PGxHAKCyiFQl71R7PWh58tgbZpDt
Q7szCXH9FUVZAJ+pCuVHNYXm0NsATJOTQiU+tH4fihvxcFXbmd0r+XpkpKRz
K6MlI3tO0Si+0fe3IJZf3X4WUFO9sOvgjnveDI2ETf9Mzua5wibQFfVZXJUs
2UJTR4gmv77m26Px9MckL+orIA71wjHlH1ClkiKnUYrDP6FNIa893dQ6kEHn
Y0EE4CbHGx9KwXdS4u7IMUFkS+w8ho+YZdhCNHN0NYX9Id8rXu2NQQdSkwhd
A3WF5ex0V6P9E9YvqtMj/6GsQLrZsSdnkdldYYcYXi4xygEKkfSApBt60WCJ
EDt9WVQqvDKcpFnbxv2beDg4rnmtgpDJtWfTlKOsQ6iCOIoHjoW6gS0C6Sfd
buTES5smartfdy0oF1MVVkR8e+tl+y04dcpGV81WUYGMsKMIdMaj9th9tgak
z05x/DrMGfHlfSPLSf+Hr8/ouQNQbn9v2b8GGBc6gWeaS3OgK+P+RiFcReU2
rzqEw7hr+beKJphb748hwR0D8DS2zgaLhhla3h9wlnwRzmua1hcU7sQULiCO
zXgJZ8EvvrYG/5NueWpgVtlJSFXkx2pLCEvMn4K/jzzUOyCDWp2ew7L54fqQ
57dIIf9iXqP6YGm+MTGPf1W4B/GJeOQ/4ygh0iUUsdI7LK635hfqWtahPNPL
lloEEfj9anBo7fsiOz546kyiESZmr8arM0SPQ5jWM32yYeRF2K4TgCY3hzH0
6Pboh/3PZJX1HpzBJgdQDaRfx1ljew7Gsavf8vRhiqtrjheVcLNMRvta9zbI
mSrKewvPDTGjymNSuE2pmgO2QCu+C/n24cRYUywdIwOM+WK7z5wb0vAA2abT
K5KbFC84DyidWg/Y21bRqkpwS8jVTWCX9TgyPCh2fR5FjVmEMFTHzV4VUOU7
DtQIy7KGyVmFdPUA9KGIsB0khHi8VQPH2fQCaZqOA7biCvZlfYnguim9gSca
zTQWp9IeC1776jzohyjBa2hbB66aFwonP8qdfNXBnpfMQN4pVeQ3L4mAWheM
Th36lMd29rY57THKCGdkq8lsyOT1+ZOXhUqeawwOwO+dexRv3FidHWTAzC6B
GqngV0uUEV14q0obRsSPf2S/dQsNzAmvU13OSjSRroKUylxxFA7urgiWGo8C
4kRzIFjkyOuXYQlpTE+kbDEwTw22U7dO/JPkmGqY+UQgPUuKm2Dnq7Fe6+ws
BRpzpMEsNZJ6NqVusiUuHR6zxKJxZgQxBLRU/t9BNIAPzE+aF89I/t1Y0Sm3
DlMGXT2kfFBsLQj4cRETskOKDLeLh4/D6kAj4RytD7LPHod9M0H986LYJiYg
vCvMtslYz9oQVykzWw9KpofeWkb54lzjbJ96RiwgTlE0FReHmriF+2cy52uU
2gdmNxKRw0Tnb1FqTfEcmH7DsgzUM3gLutYk2oUNEIfSrjwQxeJGyN1787GB
bN7x5v6pmUkOQejlai4ctyMO0ftfCypJKwl6M6RpYrlsDJdYr5h5QMg+9ZIN
aw+k+5OmPgP5AQozWySMevGUIicYxYKuGdnMSz6fx7Gx8RtP2/PADV22CNEG
uqJedvlozlp2Yes8Ok33RYKgkFxC5o81nKG0PdO5VwN8qA2djq0skqTvUmFl
8SW8A898PLv7nUYgPTuRGUmIfAk9v9iCJoY0Ef2bXq3xlHDuBwMZwORKQVcy
4lbesjQb5P8T62SP4ThrvF5PQQU8oWKRTQCAkBPt19Fckk507uREUDjysdQy
D7hwFPEkJDqNLu/7Fjq9Z7Fkx7w13VCnBZrd1AuHxPftT4M9enXpl+Ie/ykq
xnpiMDf9+CCnfFApvGVLkmVfYyEuU3qrcf4uYeKQV7/FvL7VYbqO+UM7rQ/A
CSFlr0oxt0z27QNvXp2JWkQHIKPhldMaf5fx+h4LDacMZtTdI1kYb+APVxt0
Q4Anb1QOkGO0Cl5nqsXWIYniNllei8KqLo2+VCsYXL3ZRwA6I8rnAT/dWyb1
wcHGXKBNZhnnqp4DW/m1UHmYcW8P2hPWxe0Cc0zKWr898LTcXk7Af14g3YIE
MMiimS6fcx+rUpwaqMRnldhcuWQlhiiNqWaFYYjwBcfJuOenE5vuf8c4PliP
gV5jgTEXx78zn+/s/X4XC8KM7AC75f+WoJWg1NtFeXFh4eruGt8aqEmC2MLy
oTLsv7FE3DZyWxkdrZsc08UR7afMViWMMLUH2pxV09Ne9zlBhdit9P2Ta1Yf
INaDTtdGb2s8eJg83CYaqlMN040TnT9ETIFDSmWBnqWDJgjPZgFgknnh091Q
wJDNiW8BULOG+hEuKouH0GUHW0Xm21fMxAIvE9pniBP7bCqvg8a8LQGC//un
3eHPcxxdqoRqQta36MeCb0OuZgRmP+B/ASmQT0Mdcki5T4o5hOax3iWjBgrb
l80VzPkHig36j2IF0sR6uNc/1ynPrPyP75khwZMc7yVS56SyNeNWkLY1qa1c
Bc8p2/xHCiTkIKmwzupoU1LoREX6HQNBaSWzMcadeZ+NFz0tuaKtUJaCJCVX
ub0CCif/JIPYs7RSS3QKcVKZCpNgUYNuoBsRk7yQeLCMUtZOoeuQ2dtxtEA7
pQQXRlyIZS9ZSToC3Jkv4zBIcuW3+BZqtYblzyLoGhBgukhalWI7xnbSOQVm
QpaUSvfU3n6dUhX8w8WMTFOmInFh9Erm+fIgovTQjDNyVsAed0AN/tWfWYyU
KNylfsjrosUPiVPqPlv63Q9IEkj/GC/hXaSG7UGsJ3i55zD0W+nz1ycwCjCb
fr4GDxdR6bXq359M2IxC3YO5wOL9BDUkzB6kZl9KMGnLztjmi4iPc/UiogKA
5lJbJRruy5BFbjcruiVW/1w0NRVhfL76HOTY+pJ06XhrJW2x47BlSxeV2AcL
G7rEdTbz+GzIlD8U6Fo17I8DKjsmQJ7+KQd7C7O6SoO7RVs1x31lWF3iHdkj
37vZGTYxKg1UMoCxS7iW1pM8lTNOYo79JTUpESlhBQBQzkO8348c/jg7Gvpg
GNJmSwdMxDJ1qMi/x1K7eyuXaaPwf7pMiY33MTQplA7wm71mXCy+5A99lsej
OLO3iZsjtcaT5mp26sHFKj5e9tfiUKXnAssyxiJG38j9Y7B5Fn/FQzyfFLV+
+G4/lRrYh1v4HYa7Da8EZEWOsQ1unidhTTuRUTGCZSKTPE6GaT7y8YdxPVKH
zKusCza0n9MeewkHBMj6vU4jKrOXt7keuNsMWZFvJdR92NM0DzyAb89UDx4Q
H72qHUYfvmqI0BZquwROB5zXVednR340HpYam+hbBIIm7nPeyJ1qXOlt6MQp
0b3g9KwwSm8tKTo5wPCa/W2LzlYNtMiqxAbU6eGzWrsmR1JPO2Rui8BsbtEG
fnxejRpGQ/AZkB9YHWX6Rv+X39My7KLRF95sx666s+TXIX3RUhsYnRD//pL7
ywsYFJu88RQvY4lcym0CxURQQeVhV06gvOuyfR5SxSjBWdff1kbUNlg3sLyY
w8OYeGvh9q0s3/ooGhj+N4AMZN/qHxzPmCQKCfKpmiioA5hfnYimv0wbgwUg
08EtsyzZMiqLHkIIwXib+dWc1eEx3rJgRNsbR902ThnblFeWRRNC8fmJ7+YX
PmELyT2qj7lQFzLg90tj/k57iPzKHNCbxu/Oe0eoMVD35SySP47KRPZDLFwH
ZPE5xqWk8OBmBvalQDLQKPx+qdE2BrcxtjtxCldrDXSxaA6KRW1aY9vWBaOO
qS0BbIA0DY2QZUTW3cPf4bAwhmzBXVoW/w1pNozZ7sbn6oJDimXHgclqt9jc
gfLIo4Nei+NtTnw3EB/SKgwyRqLeEU+/PTjHKOISXa64lwNozb6qDGsZtA61
ilZThQTSZj6myomCvJwYda6GqTdoxJrcrtKz/mXj3cCgbzTK1H1n4ASiCeeV
TJ7hKIf7031R7jbc+ZuhoAOkZyR5fX8VkXtLBiQTXZFl7PrQeKPK7RDXe7Kn
e8TZvfbTltYwkC73p3RN8JUG2eTJjrVnmbfoE1/CBTSKfPf2/Y1Tpa7i3ZHg
8MS2ag2iBk643aKGNlDz8UjcpVadanL5AIEwRUBVsn9AMypCM9xOqJohrIX1
+KwnqXXy9gziqG8SM8tt4hXVejAevDFZoH7lshQEAsE90q2xjBz6BqoyWUlz
JrtpVx8CeqcHCNDZM43AFfDPecrVOd6U9Fdh1GTFqIcyldLhAvGuNgVvRi2b
XTICbgON3+bCG/5pbFa62XNJQ4X8fb7MdeZxQpKONfgGw980VnZ/lweCFJyx
qEbbDsSkVKt4xLY/UPnkAwDsMyXGwDnrTaoJtk2xan1fDZEDCBAzI1vpJxmw
mL7Bbn16j/dEuiwt07GOexfLvthPvzqpRzTjy1gXLGGz1vCjCyfL17TASQu3
Ovtd50NQ0UuApyhrpHZpjVfomDpG1I+pBoPG2vUSXz6R5RDjP73Ta4VDzkVO
nNEJTqxnXwRJDTp/LDg5ybiVpOIK62/y9eGWFyD/fAPifULm+qmeY4EDauUv
zImSQ8UDTN+kRN9GgsAmBckcwgTrySTLHmkzk/n/74EaICB+Ejm3e25Uc66M
Z24yljIEQao/ENKCWLeTXLp3Fyao1dTht0mw0JTk64MyckxrCJMoqNQHl2Dw
2UDE7Zh7Jje6Mu/O3YTxUY0x3DVJX/iNvrO9S+P/Ak/5I1BtziG1wC/iwvFz
rKJp4NaQjblxiPE88D7jX+PVZXMMLeCfqB9o/lUlf3J5HtcMOBWu4p9Rrkeq
loFbrevfeTio+gYao5wRAifre+uW7MHoO1D8tDVxU+eVMGpTLk9fpng56J2J
SrVsfafwdWjN6RlPlkY2bSmXW9BDJcpyGHAIU7fKY+K3ZeQT3WiPSrtiAFyi
M5wPazd6e+Gd/Ro2mYOPnSv+sGJkFvoT/Cp/D73IR2JltbAZ8npd4g2K+4/L
MNmoVxDt3L3DrjXIE4GndDtMIfOYa8L1Z8THECu8bqUko7dWx7YMUWRq/EDc
1oNrV0NvD9hGaFWsnnbCr4qbBwaoKZyMX4J0YzG7qrba40AqkSfCk+tmUrUA
75XGQwhp4ujdjbuEf3Sc2RLYHG+lWz4iDj9+6tbb0VpNvHF9mWaVYy8hdq9K
hlJOjCSOkC8kx+WF9HOu30/aC/tval4QG0nLlC043ubFcTA3BLORVyAXTTtj
aAH/pvYkXuVv/rxzIlMHROTyJ7OZNDiH8sIN9LMKA6kQQdgSxFogi+JVd8lQ
c5nfnU/F0EfvrsmvXbMsc+VKdzThrBqF5TJR4QeUP6ZBcYKB3XILD+HRtbwq
+5FKsQWMe8+DT72A8IYovC9K8flMeg44tg3FCvRzg7WmzcrIH54VuD349cY4
DbhsC/WC2N+nD4BGdzBLgjYAnE7g6cZdN/mqxMjBpLl+wMp+aGpSasz3k0Y3
EM2Bq+IybnfYtc02ei7qy27D8RVkJDEPiocpW+16RkihvrpHUMnnWKmk6zO9
+M+LyvZaF4HPX700OAbXCHIG9bJzhl1Yrm2w0BREm2DqGaQC7yNID6a7BSOB
UIzUFnrcd8E+ygUBHdOej/+nfzRiD0uCjPuNzaLQ8WdkfJ4ScV1rBFll1ASs
6B1NGQZxu2zeEyavBvH+679wa9D/DxoQGhZgxcrmlXv1I69/0rrGLuGMoGNm
U8ZGef58qF4v23DX+zGSXRYk1g3y6oyzrFWT5FuEUIVGi/VTjKCMBUPlq9A8
oeuMtwH1mI7gBAdtD04QqxLuHBRsw0LEArbZWwBiDwq8EMYkmRfah9dWm6ZO
35ysBym/TwbaLhTzrkFVH/IPi2CVEvC4CNIvfv/dg1gBuSZQ3plojEGr3b2u
BpSYcJZ5bUDIwrB8wJUakjY/IrbJFMUiyXXXfB1ywz7A0i1xZL1YhkSa7ciE
Uy7xZzcMmUqYQsTOGeu+xUmZSPUtnCufaV8UR571LvCxk7EjrwNgOtwtHVbJ
o6V0YlV5l7xk0DlYui5pKXw5qRuOlFHbRP57V8e5j4Azi0c/GN/lg+9JJMpP
4iIyCDk8HkYCuwjOi0y+efMi90/hhM5kqAIRXev7pzVbdRPtZ57Swd8wBkag
abvWY6s70uiubaKqfLXldvb2cRx4A3YDYIxjXcV3N8z0dGLZrjT3HiqEcBhM
d2PQUKWzjBT0ImFDLCi1LyOvfdJsS+TP/xsnzu1lMSUtQcIRNiLiOFfiLEO6
KdQw9zst1PhmL04gUyIkyIadxkKhppASvR8KDlyBy+mMj1V01QdgyfTgTmK9
EMkvf8fzGZ5DJuv2BgjaCEHOvxxSEoCHALUOaaPLeZvkoI6hnzW5Uw2N0M6A
nBJ5Qd5VqdWIjFsMmfLU4Qph1x7At4RUK0Txk7SW9QOS5hgseIKsoHau+854
uSfoTx1O5WimvAWouTDV/c+sjB75yjR1z8cl0Z4u65MxiI+LaWo+RQXOGlzt
0+EpGe70ENnlpYQcvx1F1ACwJYd5X5SOS6NGuj4XEboPJrhbr6vY2Xa2y0rp
+kQQMN5T0kcfTMPO380BZ5qJeLXDJhRc7wL/hWLJ8PXujKadwuC9DNphx5ZV
HwL95jwSa1Z9QBxxlTSTmvm40iQTbipNEW+vL0PoBRSbr+P7WkZBh60mNjM+
lwxggldy/SKjN+fWI7sVYDyuN8UBpm160FtVVvZUT+E/hKcmf9x716A3+C7g
ntBFYAUfKiJpnkWKDk6UYPiDV5UmuBlPB81IJjNlw1T/xayJ5Wy7Xwilca11
ht6KZ+9Fm+wT+Td44htfhiaCE6NOLeHJ+Wb+MT4DPZWqfQA+oDCAgp9WAu5X
3udR0AzJKZAfEFcdpaOxxaIgoNC2lLkVelg3xrbW1WBhzDExKZAF7ylRTsE+
6fqz5z2Z0assiKRR52ko2CyafbX+dnMF38RPElXx9gfxyVhyPiijT2g+evPB
LaYq3lQNO/pEIFg8KAdov7fsFLu7ySSJbKGkJjSntxq6PZy2j+1FtNEmnDvm
qRhKOYHdkrOBnIQQDZgkRzTovrZ6YwYjiBuNntwa+3a5a8H5y1E2SnCk5Lpj
W3UmZXECsEyZvdDWC4pc1DxUnQQsffurEqPJB50HwcEc6FmXFtq2Ldey0xAu
Lt6q5R7byKyuYStIC7yP+jxcLskpYffHlcq99Ga6BkFzhqpfXuCuWqVgMvYc
kqZlRyTiwPAVAjS06bsZDm69MZ7q7tro0EUgRJbPUo5vWnuZeC8ej7cNwAiQ
d7vOicUWQbvBvoWdZ8FACZ/NNOyofLeEDIPEyjs1xagaoRZU8tyo+xjEWkvS
TLT4u4fRGjj7fwHzzS1Kcp1871yvZzFXSJNZrSoFSZzZo87FX3U0lqQPYJ8A
JPKDSqCSUi9Kl0Y1jVo6curZNis62hpEZaiuTjX6bJFunSTHSM4wjxJ0od2W
nl0zBZ6OpTE4MCEohLbKH7R+qsLdyAshWLJsz/ZHqQIOCPr7+h+C45KzpYZR
/MQPpoE+J8kYa7mAT5gKJqyAbfUJel/nn1dKirQeaDVdP+bZP96y7rt/Xuxa
0aTmR/AhYVOn1rg276GgBJjE02NcGJQykcEM1W0PiTOqHBiAUZseRcYZxJho
M9nutc4vJylx3M/X7xQOyahFL8dEcNYGjjfLUieQGSIKfFcD9gMlspLcNgnd
ggvmfV+9aXtXKMLfPAfhdCkg2ucZGOkJIy6BTja2XMbq+O9YexoBpzHXpWWj
ZNPVPRP1/4h8qVdoqUXKDCfvI63Kn2WzLQfCIcNO1G2wNxLeDOfY0uOOlfwc
LOMmwl6phTLFmFJrdvvGa/KpcEjttNvKqSeSXiehS0XtJW26U3VR2TKPq4/K
Ylx4UkDWw8uOMAusYXaN9CNTYfCr3rDqX7CF9f8Mr80YRuVVuubz1yigkmsK
Je936yWcA8U29dD/5kxSg5W4ivJMt4Z71OA2hRz0PC6q5oD7Yi8hOiKDj65C
s1DiLJvXQWfSjF5aSnMs269uZC/vCFp6wOjtFdwNDZ1+jn5NIbR3nFypo3+X
euUpaO+SbqUJ/lW0czPNaTi4zPrJkC1mbwxwIPGWis20B2HupZ5Co38SDtUL
mtYGNxWEknBS0FY8TGDNvRwnWEA0R7DoYTWzhYhP8GllkPzwfsyYLBQJWnxF
xQxMdPUocUJQ8QbpDvDlBaqITWtSPavRSC9GV2MZ+gC2wQ9Y1uXd8V7DRSEp
Wzd9PiWGzx2qpS4qheItENyN+/feZhQGg1JGAHM1HMNrVwpEByoFPxhV2wAp
Q1jcM0ECKhHzr/H+YmNekeKbLJUUcysm1x1uhYG1jjVvIlU/B1n3fCswdyAp
OwLYgqNa6PaX1fuHlRdjYjXn5dbcHS5rNp6Z+zpWd8WtJQI640Hb28fAhJea
he2BnocddQqieFs3JmmPkfLMdD7NiV4woNVHUVKXExp16Em4BKqXzo9gfYRQ
Na89EV7/3LEWG4b60ShcXweDh46yWDF3pHxLPfSFovpvAzI90wdH9KTkPB74
0USbXUfAZGyqvXzYsLImHJineSVm5aEnQYj6BYcl4J9hZUD1rSK7iAe2MVM5
Q1t3b6fFmG3USAMrkYgnyIaJQh6DqhLVm4lSR3AvT/Ny3TdPFM+s1Es29112
l0N3vnZaop8gc+p26ZEQCm6RJ/3+mW1v1FwgY0Ep5BaqsxaDVOj+TR7rVM+E
eQXn6W5lvAHCPlSpRY/trJT1TBVBX1B4TF/ZJnlRIzufWulZ/JUTrZZbx211
As7jigbaNxJ0+DwXcFknQMfgQvRyMhU7/6QB9uHsVZCltiu4p9v/n59PZfId
ErV+tEF2vzSm3Ocl8Gj5amXCiK6bifa7OXZy+quzDOo/hxTEHxlErPiBM8fb
PFgSUuX4LNxxJ7GxQjvXJLLzKtl8C3uCTfP3hwPkonGO5U9NkFRb5twU0MD6
C0iNXgEpqP6/umbAiIkMfiGdJq6of2VfXCXL2ud/BFEJuV3RmloLDJz0FT/m
d6hkkKyhwA/9CAwhGdwifFoyNqGbmzxn7pa/jKo5CHDdVd/DReRBQZlR1fQJ
MeIrLYoGZ/Bsv9TI9xZVhYlLJjUh51Y8epZO2qHGuSBkaiCC365tXzUy+/Un
CpDCM1iINPYDiTf09fD2wFlAMUZMQGpxRaqHiqV0vwYWK1pGjjiBb1rzkP4d
jA+bDkccu6emMzeg3msKOcGD46xu+XnpHyLNCGgP8g7jlK6eIaxwC329tLVS
Dzl04u+sXcCGYVp4qb36pou1ARZvfbF4fnpO41jbE3lR99pEW6rR5lsFYWa2
0SPZfgPZdLyhmBZi+GQiVkmBmeM7gR4kC3ee5s2IpVd9kGSIHZrFnMTbbqTp
PpJf0a0MaADWTfMQEjpcaB+6vnfaTigSUdPYF/fhJbco546MBw1ZXXN6rKxZ
3frv1YkU8AWlTQCLIJj1Tt5uCBzA7sWigjGG576+/R7xF8WCiyEdFnXgXIcH
zXJNDc31h9wom+ca+rbGbo4BjmMD+KMxCB4sEecr2jm7nqkP6+/iET0BF/Na
iVChJQZXmvyAhoEmpXjaKHFdgW1VS7HayJYVe837m73E1MUxMapAPnEA84P1
ra0SehoHVG1j0PaAFAF6rDjloCDx10EEvjtHDfFxpkJNOjmuhMKuEcclM4Xu
oHQJbYI7r7F7zRTcqignf7F3jGtPBdk/9qYBlttwVOhsIdh1lj0rxBUrsPPP
XPLRNzPMgbXu9gBxgHzzqUGqL0/cP/Fg5ADf4GVIbyeYX72AbtM5QQxrzdmj
vyhmRbvAvd7t7QnWQp3goM2cfh3AMCICRTzvCzO7C89Aju5YX9v1B8woB8ne
czBlehEOQN/xKoKsrw+FxqNnkJYxFUfuPLR2Iro0Pd7Sa62sLet8cxlogCWB
gAijj0FCsM5lkH1vda+JzWfJo/JgQHlpkaDuK1TWWA7nUAQyV9shjtWtA0aD
nXmYoDUVGRtTzFugRa0ILIOCo+bPlS1YPYFKcSAbk2XfPXVmaFqZ6yCbNTQI
IMuKKELR/2iuHEYozhAJzNo/IGDIWid7HBuuqSfDzwtNQFmUQPumYI+Uo6Vy
zEjiz0kyqPPmhihkANckboAgrv5Bx9Zk0Ass33GOoKxxO134xFqqe/SWEcoK
WzMWWxwgToV+5aondd+vs3bwJvfG/UZ8QTs7E3dn9Q6YYSTIwFQWl1CcDPIc
+l7wTI0i7ZgFlAp8/80wl7frcCa9X3UpkpFeNkC0rwNpLmCjnBP5/utR1oJj
VIMoZC5aOmaDlwqC885/O/3A/lnOh7j5sI9tyk2wK5qafpDdk75DjDV4W6Sh
j1kbWEITdfzAHD9POqMcp0wiivMoIVq9dL1kEnKQl+6k+WPPhE1fCBX6M3Ms
TlqGw0lh5JEQckRIh631lUzK3m0ycqgl8oG4ZclvXdjTO3Kgw5goDamEWyV2
XZJMh4tG6OkTaNw52M7YA0FEA1NoPAYNrquzhCgU5YksU+l48jNWqCsStKOU
zuBk5tLMP035IaDY/QCqtSqC/IgYmBQBt3NJiaXlP+ODDr0XONAnmI6YkreN
93WJdPBt0IMFlh/UVZDNWyhbH9GPmxXNXDOpHml7CNErsvbF48r0A2BdXep9
UJJp50kWC0auBa7LNtckx/c6PbebY+jo0injFfG7gCTlRweMNiiqTGn5b/Rk
9CMd24f1zPnjTym5+dt80vvgAHaVAMgUshZ1Qs6V4NtjMypeprP463UQGiiY
Zidi07m+JNV6/zgaeNCvoiWwaddHnv3ErXsA32CYe2lOYhzwpDSPKTOJD1Lk
bGEusbFNi+DTfOlpnR/hvt/lqlw1WEk0F75m3xmlj17r3wyHA9WoS0RD++aa
uQxOIuLZGwV6YWpdt3ORTvfWcFFdPxV9omv0MAYvC6KBEhe0K904Gk4p+tYO
s+iu0Hn9hGphM2A6WCxJq7PHdFt+OIX77LlmMrPQhuA2oMKH5Bpbk35/sUw0
17gUG7onlG+KujgsoaE0qxJoYBkNvyl8pwzD8E1V8DmQfG8FC8t+GJuH1KZq
vY2ZGR2qyNLNgB7CSdImEyvCa+ZGw896prcAS0RSUAz64YwgWC5UEZGjJCkB
qYZUByAB+q4Ofn5ZRDgl5PdGcuvn2Ikd1EyaEAhlu3oFTpdp1ZInbXKjZ0Z/
TJb7lXvK0FBuu9cQ5yss/wyPcFaLprbMhCTTHukC6o6WdtCbjPHP1lY0YTM9
Y//kelXwW37yxpPtpR5Id7pSB0MCLEAunEkaBrxfxp0UA46X7elhVTFRBMXe
vWWrH8HtvHeDg/nACy5E5v0YIG8Oaa3cozy62fGDTOV1Mp1UGCECtyc69S9s
PkI6lgTC9RSHK8+f0/Q8mUe9KDyenfwLcqBkyEDY8veaPSw+KeSXbVquK1Ph
eeRRw1qL8SOwLqx6nuhQOMzhmyZ7dcIGMr37fhpLyellbGQLNVDAKevwKon+
4QPt9HbV9NWhEErWVmZA+3GmYuDsQILr00XURigeFWtQURITpe7XOQ8C7hFE
yqvkjS5FTpMQ1vAvWqVuP4UxpmElUSXHhnA8tdHuJkKA5Gq917JrytfxXt3X
lpiy4bMHOYWQAZmdi9D6kRM9aBS+2yuqPNGRmh9iBkS52jC2fRTSz8VXkwx6
C9UXm95G67TTVfBXeaa27AYrvgiP+Hhni5DN3New2G8Vpl/UlAf8XpX0VOoH
AtPsLekl6Si9mKC4HCjl14ZUUCSU7KNxSb2rbN6nXhoqlUVHlHzUXiS2+f5N
1SgMmT7aa1hOMo8LxwG6ddX3kCH3I722btuwAOrggJ6YY/gT/ZfWuc7/9jtR
rc3NdFv6UOOdK/HN3j/FDxPS+Js4S/LgO3yvh6ZMr6J2JkXaa4/tP9eD4Nrv
zWZCnCSMitDM82lNgQJq7D7gHxpkPMnBfMa3dZhHCQwWqy2opHleOFBZzi9+
t3TQ2V5M27XON4aO6KrM0D8QbrAZW/0btQ6vQkjfMhtQX50G31c7zMhP940s
Y74jQT3TBmYNPrzCeQXznVrZteWGgmoNKZR/CmL1BbMOC/z24paIO9iILFFn
n8DAfiwhZOKllJHIm/tzl9caLmBlnL9aDe3Q+KvF/BE4Bh6CkdIYhRxlIOsB
N15N4I63q+mdy4Aa65WlpV4IxfjJ9GEv8WXz0+/QyWt5CHDMHFCq6yI0xdZx
0f2YSt+STH2Az3ZNhGwFBhFSFACAMBIVO2dqduaQeFQYQkV1UatWTqWi3jpk
4ER0uoReZywhEInsTnbMbdEAuKvvG6BxSI1FO2Mpt01lPSzP2Co1CCo5JqIh
vvk581Mulsqf5KXQbNUghFuO7fKDzXsAo0FweXShZg2NBP4QD4u6Lhd4HoIv
9ORKFTcg2q5LZiDpKgjPJtDj1zS34MRv8xSe/u8Qx2TB0m0kx1I3KNoc6vv4
YQ3uOtZjVCoqPfj8sC2PSWDVxPM77faySEHTSjQJVfiD1RsxIxTu2Cfjxut/
arKkGTi6gFwRlguk8sbi9fmd1aDZZksDudxl7LJ4bX6jvf54oR74Gare2Nep
Q1fzHKDeuAns1XLYSm5LYu7LQMrXzd15V7W9MjM4kHw0PTkfGglQV4tzth69
8LfUV3tPVXvvy0xJaJ5KDx5bIKD7aBE260rbxrpDv0n+uDScwWmjlF3DMvk5
kh/7gQeKP5SHRXNar8ABwxLteGXKzkCSrbwyJjGwP7Ot0xQbkuPOFQO4djeX
re8daQFZ+lbzarvJozvZc4HmLOyDZof79bnZACytT2dsxe2mvVs1fqXSYuDt
nEdJJ7IB0F+o4Nca/95YN9f8+HbNTNFuWEe/9qEOCxoHt8tqxV7pUkLPjvtS
jNbx/dmEjfHR2AGPK4+lNZ38wslnyEhrQDzMRxzPAEziYoI9FrXRfHSlATka
60npfbzMaO8hy0dyFwOOwwDIBLm3u7sn0diqXwSNr3TH9z68/CskB5Jr95pT
VZyNzgdrz8cTJm3ucqUOtWEy4mjHBAPPDxij+JjX+MYNz/maR5opfCW0iHuU
S3MSouNiP5+Gc/QO9g2TTIdqW8auEjYfG+6rUAXZ9pezBxomaBeYVg8V0hZW
rinizshqTv1R0r7sQea4WD+o9uYj2AZMBo1QlvQJCGU7mHtzkgBTdzrpGos8
5E0V3J7v8v4KxBehIpmGfBJIkqeSXq77WwS+Lu05FibZ3/Ym7qZvVlrWClVu
wz+uVthUPYcrElxDdwYPt69zYZOg9OEUXSG3unPLa35bLB79LdURbsn+oOSU
6lnPxdCeaSPuV0m2M/9aTTYXOp19ELa3uP3DTes9kTkxrJzFk7WDrKF9UdIp
RE3tHo5RLvTE8Ye4TgwHqNyh+kah2Ru0hL3hv0RmZ0T1tr4kqe9lQRQ++Ynq
fj6220pWfRSExh/cwXvkiLn60PaSLlaqgRycgkPDehRPeupQ5NRGPcpmyGah
1j50DKRZtsuXmQLN9FUDodG/bup2B7TSVxwCFEgQdz3f3hGZkqIFfr7lFma0
j65Bjb0urRa8XYXjBRLjxMJywdvPVMOu7mzRJJgVpz/qW+J+vpq/5urK8oL7
oqJMea4i8T6ex24/8JFBW2xAPQPI7AZHODA57EPIxQdEuO86zLq3JYN6WY5c
nod8WIuURTaFmnaC+a4KEFx52QAfZF3SHYLz4yfDVJlwngtl0ZB8sROYHCK/
M7vofmQVeHnwVRB2rSCAyDvsrIbw1e0QRmue6YlclDMjkBCBNowl/vRcP5s/
z2gEm5VKzP/f0kk6IWCm7iZAitdCn+lMfhKLg+RQoW5mssXHGOaLYhg8qqJa
hN5Zj8+WNg2zVGilzCsay11K3EW9vZZQ1VPBSLnEqgD3npCN9Pi/jnEFvAvV
lmf+Heyhh+Ics7UlriLXpIN9V+ByfPF6F9VJIGWHyCTuxci8IQUiV5YNuwvD
mKk0KNnRLslH86q3iEdTc9fVrIzoWfwoopfGP2YcbCI4ghecvkT/+pHyMl+/
88B9jYWwaQZ1avaabMO16bJLpUHSUyA6SZiQFxArnMngBgsnIH3tkj23TclU
o2+dzxOyHS4hFIf/X+eV3DR5To/kn26DN1OC41ZcgUH2kJcocArN9A8EY+56
pDIKwssr6iqoKIsaQxXjO8ArmARntp5D512yVUf4fK/v+++PflWm7EDWgFvu
VdHpK/4lMRg8zq3C/TRnOYeOZDzvLbVZVTmD1507+Dwzk+QilEYzsOx6LS/H
aEsEwmAjdgeoqCTZ5x4V1Jf0OtmSvaHmP0VN5U3r5dy+gDubAy8osn0ZPM49
fTbYL12en2JcYZPk3AYsxtY4wmXpY5b/ubMntTLUcHF2IWbJt+3srNu8ftXU
4O3dFDaaeWJCvNnEMuitfXX2+TaBVzNOOn5bu1fMX903rIYPny0r1bI6A02s
38LMo3GnX75Uvt+MfDy6UiNT8FyejoOSjhyMJILo8ju8hXvutu0Ez93rQqOX
/GM9hPzxotu6iHtrm+ULjJ85Otj9O3R7gOzU8x+jwCwuj0hOOD1+nJMxzxzZ
Jg6aA8L7xwoSTvpYYthoHMDzIuBP8V3CHNq1n7hQROHdNtcw2umnN1lxDuuR
iFtzh739IqUHgeZTBkZ6AQmU2wbexeDuecE7blq8oT5Q6SY8e+oR0RfguOBU
I2g8g6HVs/7atsmLMRPBzNYhGiwAgzshnB4U5nnB4nIWr1zh/LB4zZu2vB2D
vgbjxw0QDR/beScvwHnCPvz4kuGeFmgamHHvS+lTyVg3kYHqF0xpIUwQks99
b4ogTetfDwUocGEBZZwxMSJwrh07gtT3xAp+p7EBC2Jp/r/S9cCO6Wt4p5C9
Dr+roSUC0LyR/XoNJLHauC50/SCCfVr58es/vh6zTLoLKrUavYfc95Iu5MOO
vspvQH5iUMHu6FaaUdX6gOlmTFyHXrZL3F2l+K1eVjak8HowO5Di692k7xGA
teiJOlBSRUC6KBdjkcwyWF07tdNsp/2tuvI1zKvzffCGPQ2yJYt+mD99Jwj/
k5hnL2YdaGtkEw2/y57a67Sw+3s1ZINEcbkjeq24qhHVpmAAZAHg2gP0hXpD
iEHKY438xFzd021OC8pomVtjfQoAj5KJgaTNs+jso/LmNL4zEe3sxf2QHU7J
xIR/o/wZdQvoT66aKpMdZJ9LLZrGctd1dJ9Uu3RFTdP6S3CFDrmmsrqNukIC
nBllLvVtfkmdSzvaKIRayQKFgykMO6SOzYEE+ZvEdPMSSBeZoLEguw56UF8x
mZchXzjkay7c0TtguigrAXjreArRHt1QpiPT9ZfZKqLmog9BoLkpGOn/5Hkj
HYkLt/Li9CuBLyPbkBqGYIuSbrgnoRCFarIAUHDsAd0hoWM8opRXaQi8qxS6
XcNJscvXo6TYy40JiO3PWnjfoWrpKQONOBMdkMJMTD9mNSxh79QkHgSZnFfB
dTiWhteMxHPpIAbohPXc0oHMM7krWFi3zMOFwkSiW6Iya0JJS+JGfLVnmaMD
X84HEfzzjSCA9gpbYXfbhUDNnluYE/bHC6iabt2H7AcaqdzTB0TPSNQJUNbS
WEEBnzmE5ZEZIb+1r17sM3lh5vFbhabSnSPn54QhR9ZYLQYxLlUICC05p6me
lhNq1ch1bY9YKd/2+yOp9Y/WM5JFiWGvdxh2HusYDtyRHn2t2jr73tls0tlm
2w8c11tzbHkX/24Tt+nsYUc9N/BppHwHilyDjzRB+W19/1cuPY+8OHdpAjJY
5emvEWSZ1IUD5NitknNefBB2wAx8b0GksUrTOSOMGJLpexkpdDU6PCg8zMxr
6D5TJmEXnjIFI6MK3+z1NZIUjg04+bHJ2ZylkMcak54yI9n/4/ChCcdjD4Pb
hqm5j3z/g7BoNo6+toET2lHo/agJpzf/FcL5GpXwXby1yJitoCe+cVdWxO8h
wpcy79yS3m5TUOVb4CnTRUtXJyOtq1fXrnNWGbROOzKLe8G1itczf1DR7a0T
0O1S2WwQhgjEBg7L1jYEVmaHsqkYiZBp7vmA5Z/MXbEewY8djCSyEOS7X8Dy
34uC4DyjxTWaWnO0wjAXSHEuN+ajmPU4ZAtdT6rWf/UJy8d2qTCx/8UUvswp
cPeib+TV5x5GWixllr3LRLkrarj1np085o/bT89zOEE8x8ZDS5H5MZZIQK6q
C8WY1RTwxZObDeuz8EL3q7I7WWjvGo8iFZ9Zh3NEQuax8e5K44mgBzElRqjs
zKjWxJnqSORr8EMburLLMryO3qtqGbHBvHRLC6pVFr4vcmwo/KlX1c4lspsv
EvQjUHndHxbUiNnVTu5V56Tu6Lk864V+W/zHQt49zoQP/kqvLdSgIm9tksuK
Xc41Wt9JXQRu98zuZdb20OqSrDwX82ItS7u/iFHeWHtHgB77ollVJM+rnBgk
OhtriS3xDI5Ief0cz8dVlsFHD/kfVQwd1P3hb6jo85cpj3Z/r1M7I4RRemdP
rferzaP7C0unzlC3QgBBuUXlaF+aoju45r8l+6VKLuk/Aifi6K2TI6IZ8Ocu
hLzj6ySIqwUYE4DIa64AbIvGKEZ4Dc0LHgq1Xv8HbGk7t0/y+X2eIc9cTVBp
Mi2Q6E3r7MIm97tyr0gsqSlGFPUt0giJo7ig6sPL8bcxMiyABtXCidoxupeZ
5+dNdURWuihgBb4pnRd5hqgP98YEkPo3ozuWgQRXK8XnwIpjceGaoI2u+fK5
bzWpy35bAWmPK0Ai1JfbCVPzzbiWE5KxxMz2LjQo3Ti/Khda95fAyb5zilIf
3Lr+EDV7ow2JR52xS0vgbnoBBwfXHKGo13gZhy8e/VKr9N1r8N/l6B7Mwl7h
bxkKBY4orQcJOPOQjksfFlP1m+G19a8VPcwVLu9hq7ZPRFYSLuQum3NSsYMg
thV+tP9yPVAWZsBSWbcAq8ST+K7ASE8gHA4wu3qg1I85bDjhptEUpSuBiQGX
nHsjmexhaPlvzSdCkwLwtzPiLVgqUedAjSNB8ejWGOQP9xilCqtE9ja7h4QP
QLEgEtrTY7ofDHt4dy4lFEQwX+YcVkfDes83a3P7iqJkvQHQbUTYMcuwHzux
791HxLBxVrOsVpWiUmcUqBncuUY8Z/M9agEJiT9yUgXQEYTXhAbTom/sI3rE
IXlLTAYam8WCIhKrtIpTh7YcbaPgFwnXJgw2rYrp9/hWm8SdESnqew8cQ1t1
2IKZA7roDGekHcjn1M3OsV6lruqvBQxYoQ5QAsBtKfU3GauSu8vJxsGcN489
LDnEthQU+ulJXUZQQNPuZ0dlB2ndCmcxvmI1rmSlfvK178VMaqCo4cm/nB4J
zHzuTOtcRM9QvVwxUepNu5MLrFToLJT5lHmXtqlmO75c67XH2XUbzGWTZe/6
VbSBNc7zJqUlDJ2zsLwp1ynJN+0Md320b3UqBCnrvZbOQ1d1/eR23qBZtNlF
Vg1nuyfG6tcGR+A1JiVPQw4KMK/SDGCUkeleQGebVmyBiSZ2QlNgjn683mTu
gMHmD5MIzW/slfrSyxyy2OftFbdFnKVvkyB9ysm+7cGxwieDa6XgjOwSeVbR
fV8PUnTMD8I75a0GLyNpAmxd/3AatMC7vLQr7oZqME9jbwkT4JAlUUjIfjJf
I1zqbqMM4Xf+oIL+I2qMsCRZJdcxpzJE1gmdZ757RPl9T8KhlOT3Q4gA8VE/
uveqfO6Xr9s468XKfvk3T56XUpYYjcROj1IU9gdpceFXuJA6apdNZsDiKjUE
TTus9QoWqaoST/zNiQGMiFM1WH6wfypXH8WNC80eK886We+TBRVjpbbowK/G
Tdk6XoHEHtikGirCSOgBmZfWS1xKpQguBWv07qJ9IJwvpy8hOJJ4yk9VkDNM
58Q6ThmjrmRNhqhmO2XC5rscYpFXeZMUN0Yj6PCXcHFvUlm0/KwnmPpm+o92
iERWPprhUfjnwuq90X5NeXu/kcWpwtMxtpReOAN1/GxnHYDu7cY/Mbjwu0WE
1QilC5XnYVm/lFA/IUkhzLX6E8tLBfcDokhXm2GiTCJv4n7dM6uNAp2CnMqC
WXHj126nEplE6jDLvZeu2ny7fV+B6Y3C6NBuVUW0a3kzK++YKjbeqQHVIKO+
bQtwHOiLtNQJm2E7VQzqBilOtYAPjUfDgo7HtiXpse/w2DFuUVt9CIl1JO5Q
x9KRw1gBYkVUKtIev4xS0Cnxm7Pf1cpg7M3R0PJxSD+qabWbQQeS7qitd3FK
yC4S9j3BzD/TVYQnA6jQo1nZV4X5yt+efzoB3ptE8wGfVHOwcsPIX6EXhh3R
DtCxvRPA0pNqQcX2+TBSYd563rIiUgIHMGNgg65u22mud4Vdq315AukG3CMU
G9jLhDI66fDY3Cz0IGE1VhuG6Nv612zYxqw9/y+P3LTsubiw1kdktjqrHRnv
uWjZ1zj//W85vCXiDFgfGAXXO5sPMCpttZMfYvIXj+Szkr5F9f7/Wz8HTqKU
xoKUICH/i53ILtltT9k6NVw3fvPFauUYgMOlQISWs1xKLfTMdqD+jmldWIdq
Dqg9AVsvuOXnGa0G29AK403yp+MAmm8nKeQLwRFVNtocS48EEVYunynOk4Up
njCEopcKElau6DxHLrdLRl8tiuzm2oKw35ru38TG6ZunU1rt9Vfpetxcb+Qh
DQ/TrnsEiR/wyu82T6QpB/rDQYp8uf2ayjrnR9nC89O/VQ8JtlPXGRNYX8mv
pKVY3qnyqSBEL5KwnAb4rMRurlcCdoAqNGQQ1JqhL6+Sop7Ag6mZ0TJrPSpM
xVFNrfA85FMyjfZJ1NXPIrR2vamJGwOZa07AYiEpdZ1YRY/KMP/ZnlPVSvYB
PC1aIphRjA1tD8JtuEYYINhiczDHe9gzC9TR7zeO1DVyT9yD05L2MWS4+vAW
NxQ4rKFPAlCe4XelLtCZA380t/o50F/FQq1a463oMk+NEpSAnbp7E0OrS+fn
rUYUOK0Xt9PzclrtEwjzAAjxpAIWF2qbaEO16McIT+UWNN5gEgjuRgobl8sB
ljN+LBygEq0BLXIa8P4c5j39u+GQWOuKYQYThCkgvwXLldnccpB/dQrwV0wB
NtE/l2tsYly0xqBEbpVwgdZEW3336h9F8jW8MJaqaYn3I8k0AFI+ozJ71F4K
OazntbExw/GMsRrvDnpgj6hIlQoGWxHr+2RhATLWyhzxUTot3mcD9yEapq5F
40cPNT/JZLieGRyTCIX8g13X13v9u3YiqCF6DAgPX683w8+NQp//g4yVgWTB
6SnaWHba7niWHrVNKYrgZN871CKw2GTCkkXLxMjrgmXFKS+lrKkmZ9sHiZMg
Hnw9XkfKRp/Vl1kTZRaO/fL3qON25FZjB1JUIvwUK3lUIGdZqNG7o6PWOGjW
GQDkR31YuIF0kOrAshBdfa61IB4iWzH3sc8ts6h0CbZzksk5gwDb2j3r+Ily
Y7qNCmCNQjqHi7W1Z0OKbjt6t9JSpeVPx/DHjiAeNIKuBl8VhkmGl9Hz3h85
rtYyqdYk4Oa/BmDKwmEGgoVzMo6tk0FQuTBqHHWb+rhkfIWv149G+Rxcyo7P
DkcOO0PP9cn1Kdpxbx4VX8FCVIlUJ8Zdo4lIuKBZr8x8KJKTIvRU8SO5Sn0a
ttbNYCcHNTfvSYluGnumdFN4WUD0uWdfICBu8HfcLIGUu1n3nrJ/5ZFt0FCB
fin5OzM6PY7sOyHfLEnZJ8N7NhiBnZUl8AD4ShL4AXUTSZaqODnDFD3kMTcz
bozemFyHmdPGBpmdDvqb5TFX9Gpox2O4sc97js7kz3RJIQ/nM/fALa8hQOgk
FyO1xBKJHDKnBLjaL6IWmD/nDbvELuq83IKwAWHkkEkish2tXxnEyC3yJ8wt
Mha+SuU9oAkcJOy7y3xySFOU7KRF5/ekIKIcqW+HyzoNYL8/pbeNqcBx+iyZ
jOkyi9ZMo+46DgFF2bgjMyr63lvrDRrJChE5NjpLC2Z0ysFM8bJYVQ3HKmZq
6avVOUnKoqRgbe8vHdtVIMgWx9sWBIMOokgJLvmYwr5LVF1YXJfDqoVxuWAu
ZZOIjlnLD6wQ0/r3wIQvgrcvj+ECt3HM8I/S1XC9EJRQ8OBw4HeuGbUoB9dA
m7IOi9+RniR7wE0djf0vsb/7C+4/NxrYVQe1gKXU1JeArE+Wmn+vV5+PI329
k9qmlKK4CjplPzEE6MqAq8UeVrdwBzfOJAiiXwhMEmJofEsVO8lJhG0y23gl
blQS6Yollkw+l7h+zcL7NLtGDmdp28jJpnLKiHGOLgxC24EYdnHI22pk1vxB
Ynj7mC8TOIdMD6pQGMVjUKprh2rg6WG9I3TrUv4LknUDCAhIhY6XAtPiXmkj
TCI0SUMBXKdO0uZKX6hhpWQ609TK+Vgcr5k/Iwy6z2siu+jzyYOHl5VAAKCG
vOxF7XD954XeW/gdXfgMG504rBn89wBeYEvjWvxmMrJeIyNvfvN+vS5eqmT0
xs6wUseUzYXLHuutDFNk/KFKsIZ8I7jPqpR0fg77wLlcz3PXLK/IA53P/gIc
NTcLjD3odwoZBcGKHLsD50TFkWJ6VVAijifMB1dINS9yd2IPJ5h/WiTXdlzk
LMUikGEdtFakDgUQ0D8AbI04cQOtyC10rQag0MhsFrwfn7cnqwVQKHtmOTte
DRhRKayR+EZciN9vVv8zh7ywtQu/gvNpp5uClVSLUIJZ73eGjv7hhKxztoAy
MoDTZ8eov2tHLI93vJEvFk3RyVi63yTS+5Nn39ud166uenSj+OEI1EjsErve
lYpOCB7gxh0f3U9Axz6kNEyOreiNy/zSqBWA9ru0vO/dEWbmWokw278GDpJq
f0Ago19Fpq8LJLC1D0CJ6qwuv2XT2RWyuFxCrMAjr+2lmqX1XdofGQVSt5n9
Wb6vQQ+8r9+dAPpNz3QTOCeb8hx/o/34ZB9H9cPn14UuY75wPJ1mUhMXwdGx
ZY+rmEPuRf8iA5h3ZuwqBlQeQ97z+AXuv6yDQdSpot8FnZYDUWSCFUvmIeq9
sCvvV7Vb3tGrheOpF1QWX+Eas57FtWlffBPw0v9QosS82OUjNbZbRJnzMjbo
ak3AdqAXq5SeKMVNSWvR7S7kz2IZVMtrvzTA+hiCSne+kk3TUWP3FRFxcH6m
0JuBav8759XXeE7j7mRo0kwUpGGDtL7VDXUlZliEkvgf9qrVM7FJgZbnD4vI
vD9Ttl5x53ZvQV2tVI40IJfQmPlY8EXdsf31fj5NgqX8t7qUXIL0bDJxSXro
irTNn0V5KPeam6SaHVRuu9XRpmtm4qZDFXngyEyvdTfJjPb7h8xTkAXWm5yr
sxCIIJIMmeZWrSKuKXpmP4E/iSUeyLLrc/6BCO+2sATnkR0nAVz0G4iLm09R
FkKdERPDTi6epEvIafJnHQVF242/0/R2OwvB3axa8L9bu5y4Hr8mK15tshUh
3xtyUSMa6VdT7kHMTbfCt6SGphrpXUOLKcV9rT3FxZNGd83bpTCchGMeAol5
o8/kMryy0yYa4TKT1YLvwwMwM0ZQFso+idaxpzzjXn1njto5QVcvjLc6jArW
XU1ULpTendyZRs+0dkdtvq/lCr1J0+mmKuTCCjS7YL0L1+URmPDYeKmOLoae
9yx909Gi/Iy2nbTGgodQjiNZQY07fawAe/1mwdrD5C0zMAHMw2u8H/3QcYOC
gSpoeOP/XQ03VoICHqLM2V/QtBUVaeFqcd9HXg0FM9Xt61Rl0UYlvVwxIR9F
2uMuFafM/kXN07JRCk8FU1TJBv5Ot2s9YKhVulWn2cJ/tXCd+4WHvYh7CPFr
re8em5YsMBuNBqRJ/wbDDg1uVGB1Wvek5t3b1im1Ac+i2zPQ1g5FLVHpRjUR
y+KcAIVqME6m6O1gdTX+eAGjcd1hRhM4+6phXEM5P2vQrzIH8Nqvl11g2q/m
n4pvwdvRJbbFQo8qWI8j/lbs26A4UULa6Ci+A+PgHu/D7ks2DRDjAzIU2vz8
UN+C1FxSnasNI595z7aijNngkwvJrELaPiNO7E2c+7+UdKtQAZzAPl0Omkds
zowz2Ux3bZ/Eb8blxyo/DvOAyM7UqGPHJ5dJO1P8tgm08RM+SLEWz3/qRVDA
NktI2jtTYIwJvdVZu3iFpraalu/suQuLDKjVmOrQBM+g9XgaeQkrSbUSp4i2
a8yWqgubcojdCKcWEYMvrfexXD+PK4a2V+z2DDnMwrR9BDGzfGY8rCyYZYb5
Q8bZRFNSP76MVUmv0dNJb9KtglDXm7NI0vDhqZ9EQxa4x+xWariKr70M01yN
zvVsGTIECWJ5gkTNN6Vn0pDTfq9L8wIxV2yS6KZ9ojxdsZIZVo5dVOE1GcQX
msLJKI74RTsttuJoneOv4qNZePBanf+27ofNmRi6ath5VkUeNG2va32BlXTK
o0GOFDH3ztfmTNUs6nxv7L+hZ2NIVG9E+c0O96f++z9wX7tTWMT26qFnMF4n
zLeHAihl8odmziG7r4UcT0VoDMfjtnx7W5Ne7ZWyisuc5nXS1qUjZvBdSMJY
22seYKVXJRw7qq6Dt7pl96W93wP4Id5A1/wLLOuNeRToo4eG+s1zucbPtjWz
o6qqMhrhAQBP4zNQ4TcL9Jrr+ToM8ILJfJ1DmB73UMsgs79J9l8RwUbDM7l3
N3cnCaP4D9FUZZi6EQsq0/vjW6XaLhqYcy9DLuRNABBYiSTEmm3ofE1vRKWW
JI8uYFYfVxzJJmdxk88ImxN41XCGbzIXPtiBst8NDswz4AzYhW7Ip+pAWswU
NaLjGH8Tl/+rs2uNhAOz0JR/WlTxxWp/WZ3gTSoDrt2EbU2zyb2foQHBthQo
C8Dl11H+UWBMDmbykOgBmtX2v5pDSOU4xuTdUJMqoHjK+BMRnYLYy5vMtWiy
dOx0L5gzytM+c1+xLFKWobXSOLsBn/LSKInWNGZ9iunyYn9/mhk3SE4sdeUF
Jy3DOIa/6+3nJVARloO6vzIAGPofFebwa9pOE5mkRgJ9fBCAShbc0fjuoUKo
NtZ3T6CRDiCp1iOKvlAm5AHcVD+iPoA/t9oSaj8g/SvQT7t3FIytT4RPfRna
F+av7BjgJiai+kJtHkGJAqm6l2mDPvV5uF4Nlc1nzNu+e0L56zOg1nwj6qgI
/6oOCShiHXDRJALTpdnjYRdEY3qMo04aaUu166uvj06/RlwfidpJ+2GYfPEd
SmaPYVFDDf8TSyQXvpgh6mCxz0ZGYx6ZcWKRPE9FA51vphse22LPnEQfpe4q
Pp2l7aPsyCK8EAilTOkqHqJYP3BdzdWeEBAHmzi4nJPczT7hfgrjYyc/+YY/
wlAvwNxie8dRkA+nDfsYQE2Cdly4/DPB2GIs0N6vWsky0NEjOKBf7qw+DHvE
6zeuS6ibr5HOOoY2uaHzJVlT1f+uEWrc4nTCGcB9gkwleg6gPknquBfjnlFE
YcGpd824tLO4RDOcIyf8pQntJfSkvcR1x8tZKVfXVW44c8rxuc1c11XMSOwm
jlB67qqcMHLPs1miyRlUpYt0vlyplhNtlY++MhcXiA7dHMWX9OH47TSHm/4e
hmIUnliGjCjMEDJxop8Sdt9gwygDWysm7bqmkrgVonKx6WzEA/0bfWbEPs3H
zLkSIUKXu6VEOYjXRFQKCXrZ7AGzsazlX9HwY+y2fDxrOahLmKo93EYyEuNK
bBXTBqM0xvl3oNfGUJUJ+U1iHq1GR7wIJJLnTHJlfbNrifll0XXkYVCblT/T
1k4sNp8y1PrH9iG4B29fYnKeI3QMHtHmEXCT+AOoPJRTC6Uj6/PIF8Y3cZsW
66+B+oVtj5hZZRRAPI8PwlSqgUXyXNIKSHES2FQZ103zdDKFwTK/ftJkMwrP
MfKeL4Bll6WnVbsbfHbWFtLMc9k/BPXL7reLmwGbIy09GAOkzChElhkQ+DpW
KZq87jnbUItbu9JtlzpzFZ0zrGHQ2mgJE8qtIRGaN7mGDNZH6ZGPZl5cbjL0
ZRJuIWfmdRXDx+LtaPacDXm7/1bAx2ILezTzzmR5N5fNW/TZKzZlcSRVmJLL
e2ATWVSJvsKQ4CYt24L2fS6ilfdM4CUCbM+d5VoCjfkp2x0LTSRlqfAJhoUD
z4ft5F/OosmajJg5Qx5Mq3YMt4tc4+3N23V8y6G7y1fEg0eubO007s4ukdNt
bjrhanvp5SpLjGA5KbXlENjh77h11dEEX+Mi4T0hGzBQhsUOcAxjEy+CYb+F
gGluTdT+My5Q29uo7vJkf/ctKk6Aag9/IziZcc+beu68fEVF5Yz+On+f5r03
v4G3oaobD/5OUIqleiTsLZemKB0yzcgvF5tfFKVqxbN7k10KIQC/nToAF1iT
7zKUjecrbY7Yw6ZBtL1+M7y4M9PGnz+ZM2XR4nY6iVxoHlNNbg5NQ9O7k6IS
1KRNhtLB5gYEXtYE1yLi7NmTSa3teQ9bxn7tTpSWk72F4pA0l5EnoDqnVmbs
K3L8ITJXgpp0LUha2uyKeUI0mjEa6scV2A5bxR/D4Zuy9dnHfSF4RaelLIEW
y8N+DcZw35unrt85UwJacHXDxgy3PPC5lY+y5kVIr1fqrSrsfwW3s32C6H4w
FV02LQhjUS+vzW3kwYZAB+wD1ETn5Qlvgnh3V1kZxv9niiEGZsPYZ5FnRKRH
zfH1tDpxwehaGqz8cHNL8aAv0VccYM9h7T2lhqlaHSn1hRYqOJkDZ3Ip8SHU
c3dG7vsXH/9ZLara3o8/o06lxwjg2Mi69nva9MSFU/ug5pRP2oJgeN9MaYLB
yhpMCrqgv6MAFWEgoA1BvWbeb0KOrayj3/JRIOAmbSdvuGHsudQrMKMoY3x1
HB6NuQGH406bfwUL4xbHISTNAN7165F5xYYUYt1Ic0Tm1xz9erPuE2nXWixi
r9HmIWDpAiF7/nXkD6aXkeG7JHswsRRxOm1YkBPoUIqmltDZaRIdaEBV/aiS
tiLOL26759g9WpA+mq6Rnt+CzE5eZAwlczKAuxv0zXBoCTeU8JBVdyU0yWfX
WG6QnsAX1qfMZ20T+1xZ3GIPoduK9nuVE9GLo9A17D2X8IVrbqKuiKhI4D2k
jHNn2p1YFqbaBiSRxy42hjK77qoh4iO1c+OJolXZZzwq+oEQc/HMLzpicDuH
VoSmY2Y9QYzFkmaWwmZLjlKxRGYfe8KLwGQQkg9Mtkk5/uQEu8qYIh2Zb3Hz
I3zRRKwDm/d/doE4zVxBPH+hTb9A4y3GiMS2l9NPIojSXlKJIAwcrLS5tKpm
y5ZICB3QV5ZhcLDmhO4trRoAwzitfsY7lcK4/ESmpdqTuoloD4t5sk6Q3Ocq
u2qE0JSUv3ykMGxM7OWv0dWMQEdZA28pAiP0Z14wiD/SXVVY9Et6beAqXXyT
D9AvOryv3S4A+a4q5ePR6E4FjsnyjSMJ/6KMLVu3uKUOFf8m7grNCZFVjb/s
l39IAgCe//+p95FKMUQczXGf9EExQSDuWF4bc40vtAaSofBv//tlbaCS2Bd2
ocgoeUuGOTM+FWbea90dZFiZCx6oMs56VhfOS/DrW+sOFH8vPJceKDL33VJi
KJCTrfVJwL5JWURQ5NPzSb4GDIjQIfZDfEB0fZEEoxIzG3DRWR8PWlbOvLYP
wqwHggg76/VvQlKHntP0cfHwfWHH6xtu1EwBKSFzpDyhxDwYvT09EXMI0TuN
WDbdLT0I1oLkEQvYnt+9/c9BsjfkexqJpFJ074VJaf7GJX1BSqTIbRy3zOEC
1gDeEJkksGSFOxF65TksGpGBzXj4iO4XMM9JUUxD19CfyPttRQBQ4hShPJ3U
U5Z78D7JlZ1rNKhc9sbrsZ9RsbfZvoRaYOAFQHsuqWMevHyVquUv7K4J1w2W
DVTXWmZGnmJ5sAqdWI2EhvdTgHJOIrU+BQwgjOV8pa9r+jB1LmEzX7OCjS4t
/lAhpDaTz1yxcJXtfq1wW9gaJLClElMNsPwfqSl28yCLNaD1HchEs7D6nCtK
al1BR6HFw0JsOwgMMlnjafThMnLgRe97zcCx99VmOKbywpaou5MYj2SnxxvY
b1X8bPBbQaL+FePcaOJQcyzZo8hs7Z2sMcE6DwCoUuYZbSrkPqs7tim3ZWQo
N7kTXytNJWEn8O8lEuYaPiG32aQjqgQi7kP+PeuzVTM7i//oXPDFtS6xRDj+
yrdjbI/xJGClm1ac+OZ3bqTkzpnb15j7gnPy6qKM7OEvbZ7uVzPV2DJqxVP8
FRysBMRUW1KKcxn5HoZiC0kCYrR15snKsrNZaQOqqrnfn0K/bi+/I1QQSGgh
0ARosOqaL3L6XKQpiAuOo39Sh7ogsv5d62qM/1Zd33WTwXu3YwvDGOtj8UhY
BXN1H8RuFqru/X4nPd64NhrAy3p0eQnK0HcQY0uk2sdW1MAMECIh3UmsT0Ex
lqANVZp0XlW+DcmBm/LX5388jl5qzuTnKgz9ekuns2t+BcdF1r3fxuHHzyDv
pndahpBsD8spEL9zU1oFCjG7/Tv2+n4ypRxqxk827IaWpbUqZxxCbw8IguXm
P/wiBhwbjVlxjEGeNGEfDgXYb5QQpab2RwNWIJSl2XhilKNuT7bE8K0ySKD2
ncAtfn4Re0CzsfWES7E6VN5t7zLD7kWg2hYk50WBnilmkqjTmRdcuCYM9/MB
YC3/qOVjMEyKzNb5huqmG4IBLvEOcjoUMlN7M8KXO7/7BrDHgky4djh07Pan
fCUqhW3OzKW6sSqnud8n2yeeC0PcgyuyeN88uKLPTeoTwK5d3xH6UOo/L1gi
lvE0PWHe0FggLqo2g6tvG4eP6xIYwWnt3oL2iDJV7pldpWlUf0BfWaKvxS6w
vLCladmYdaBm0oJvIgF0gNp6ruxRry8bee7xYRSHAdjNcenVsA/FqK91G7vL
hsDAEcxi65A5Pl4CvPVAItRjvqMNDjfkO8gL5E57bD7COm5bafmppXPiN+EN
U75F54UuNjfdnBi1x601MbhAQwDfczmk4MoiVkbfO7fwrRldzRj5nBYuZ6fj
xKqHvJ/0SzcKv50B8LUfR94SU4elLJM8Encfm1aFi2KkMXK0FAxXga9o47uO
qYOH9BCepm16dAiNci1/7YFVaV4Z+O9rI8cKoccsIOy4MlVe90TyxWj+X0tQ
0sKpPFvWXKyFJtBrqPwPPm0y0K5BTmjoLxg9vMkQeshpxeKzyRv8Sf9FaMGc
md6HZ66y7D7Fe2QDcDhCdOmNGlUXQaJ/9x+8DI2nQAfxv3CYAQyn4S13V3AQ
Dz7WwOkMjt7eu2GhEeH9Wuz0Nz4DXNnwKgS9/EwX5srtYiY3omL+7sSwjrDT
v6fQfBDOLUhtSwfUaUJWp3xX71P3Ktf1//a0zN6uSAH6fTzpiCJ2S5mhBe4+
dwwK6TNm299OyF5g04F1YO7rU7pM/jlGappHbt1d8GYs/Lh1b7HbO0dtv4gc
ZB1mLw2uh9BhZsWYBFOTyxqjJNigLLV51X3/V5WvRgzYlCYrHPbs6L1sN+Qn
hOGkWYNZXuEL8HSpp1iu86WbtNjNZpBh2bPlub51Bq0ufoOuENh87aJer0NI
970L5kBcUaJEOorya1/C7XRpZl212haaYqyrBHgdkLaqrwoWOloZinuVvGry
37xrnH2X+aQfM4wDKjETsYU5vbpnqOZJ2v0I/lI3aD19I0F0EUeMiMk7IJ07
F/Ol4wY0egJ7tmXtlQtAxf+LNovK/jttsqCAclnRYTGWxnRchkG/KaAjbIu9
j+jnGlIxG/nUsAxzj5qVC7olranVyMSfSzIVqU38tAJz5IyauGn/K+/u08gf
nVa5R51unhdwFhD4/yZE23gWmZQnfWlcCWe+MTVssHybto9FNj2UgJxzfH1f
ky/JZTF/uuFBJ1Vjh3vRoEoycfmbJD2y0d7Z1tYnHrZ49AEROiTb4l32kQ1B
vd+5ckzW2S1a8m7MCPl1+C2MB38M6LsybYxbjceoiUnaRIjVLW8izBnK/VKJ
zh4iPNSl8gN/fsgIA20g0TsHQGUkqItkFLMJEo1QPF6mj0Twd/JEpBSWGwCg
lEJWVcqDlbJvR93ZqNStPMy4bYvVN+j8ziMpJXZm8pEIm4+LUbDGpLaRyiEc
GITN8Vy+guk28wtAkOyQI0nf1UPTD0jL7b11eOVp0Tz60EDSFTKrvBfOyfk9
i2ECspExntg1EIeDjan/msIbm4cbdWGchR1cYqfalpgvzOp2fA++PkuAqIsB
x83/z+RIJ0+oZ5YLmSyHxeFrglAiaN5HMN87Jrf0IB+4+MCu+ldQJem/Q35l
rT0w/zXS2U1QaBmsCqyfNwH50rOz3PvjPS5nAybhHp/Z+KqJFWRuDTDGlQsl
YFUrjjNRAS47T6zd0QdXJUO7oqxwtIhwIsPoJIFWZzSDDletrfX10osKerXs
kfYAvLrafdIjKMf1GNnQa238EsI9lO3poXH1WQcHzqoNXYvFbeTC/hwm/FO6
6nuepc1MPnfCEO1Gd2/2+b0q4nqVH1xT4C/C/TGj8l/JXBx6BSb63SwvupJ3
mGVbEtM6SLobPvw/M/nO2SKdPqvbtLe6r1QH8QQt/bNOvTpqwuin4keYT38G
voEqSGaUEhLnYutLe6fJEq1f9+SS9ryJzzbsCzij0nh6ziTrJ0BGsfnoamNl
NFJarlf7ejOn+h268Zn7CdiRIKgmIlhXvKplZxm/93LlGSRugwJ5UaHExQDH
LuYhjB7o7XFzqvJSrMbKIrxG7scbhssBfZi7spFfKRj9+sWbC1BFVwM/Q80k
Ep+fukQIby4PbdsmCZ/A5MzLQmYywG/zdwdM1At31CtBvRtVzVaweHX/Ov9s
/xSZUptmFAHRs5Y2nSqFvLXAxwlOOXtSYkzNNL6eJciHwgZifpukeRcbSRxC
4HoJ3Nsnm6p7aErZXXtR3VljBxdJ0ES37VUSrT5RWvX8awtc3aS41+xs4P7E
mabMdBp5zfmyTiZe/NLVa3ga2SgnOVeQuwWCA4EAIXqVIYmcMqrYY/uIF7Tt
CUa/yipjyI7w+PT7Uk7dkkcQrK4FZ7pysLmB8k7XeuuKSoWzVg2jpVUoijb4
H42dPkWOYiRwjwVBYabksUtBifVpURGegG1pf2qQCZaw5nr05FgmvXuMkv9Y
pnrt2ydBdkr9nhklfEIp2ccrcTxPidJ15fdfnv0/xBnuMmd56+z25ag6aAyP
EdOTf7Xm9hBIxVEoGEx+MtcWSAoLo6C+P0d9OY/tBlKTkijivEEw8GxWrk0m
XaQgM4Fi/99JqXRiGKbSPmBE3oAdhvBUH1RMHBBRdsK61qExgv9ufM1ZOgt7
CPPRF836tcVQrU39JIIk159wy5Qom2R8couk94ZkbRIqoxj9PkG1H3OEjwAT
JhybG7xHnNZtzycDyWrz5FVhJ39/JuLmAeo7oN8wAg3t1rUDViLHoCSvzFL+
6q13wwmH5jkH6pTjtnyMcClQ625KMbCyUI+0DmXmaBoqWWYOXFXFoB9/Z1of
bZLGAigebECa86owHI0UbausZbYMebNHAH6OCF2P1HLTu7CQiMEIVy9GPueu
5kc6bzc6ugWllxXgw4EhM/fdLNSpqBgSz6yRaOBgWXV0jm0Mzm5oHZNdrH56
2K2jN9SDpIq95FNBjOi7H6CeQtreXgxppBz4R+qocuzjiJjNgC/hl+i29gzB
jiRNP2WaOqSV+qRdPxFTGOpfHkyfpuBHJrtK/K9ysth1kTqvxqqdZPt/78QK
gtyUjnwFFGdEY4qHn3KdkkXL5q6UXaGPRmwRCUgZElkp8bhTEvv45qRuFVfc
uarD7KWaARYqkG6R1xwtCmvRXphT8E+JNlUeEpvm1QlFc+yBwOGrOt+wfHkZ
eopqwq/6Qyq/r8WljRQrNQ5oQGy9NIlFASJYpSiCVidaHLO6Wo5tGy87bCun
HD2oW90m+2MF5m/cExB436hKcb9w3wnTKf9+oScvhcuVdncJoAx1n7EJvWe8
a8UpfXf7oZheLlLeYttgZM4QJGtBgEt4jTlOE3Zp7+qW1Zo43ZyjMbnaBb4B
TGw+8BHKxvhiqWcPjXrA5cjkldn1D5lADs5Rg1HMbUZfbMCYacBVFK1GLF9D
uRLa3RBeqmYqMVjO3wFxYWYKUG47sW7aAgUOijnD68dQN1ziIs1B+EQRUQiH
XEv+fMcyLafI1jl8Hpu970P2HQ1EIPCgojzdYSEevxKv/woxAogJpkXo0xf2
bNEp/lE1Bbm8P+KN0Y/SuC+OJOAhqz3yYNSj3xK7+lWAzVO5S8jMJ/GOykY1
JtlXkY0rphqcMx+TqxShIigO4Qx7eZEMgGWYfXyoPrL/CEmY8dOAC5/WmTeX
6HdvOpOonF2rZgVhUKLEx1a0FfkbcqrnUJNJrwUEGkqC7JEwGU6lkMGh+N96
bbCUIPhb4v2WkAPfTBjssmLRcOpsM5M+6kJ66xYY2gXT1LzdydVJjKXEg9LE
y9jjY7X7Nd673b9CFzRJ+Oc7wyCQIGfZxHH7GB9n+6yz7Xk0Um0f8/htEPBN
D8dqfkycrDAzci4HW2OmQrUjLJBqfT0Cp61MkEiBdjxqEdMDEcunSItdJnH2
+XVAFZ6AGOuhhQn24Go+U1hmaTQBoCtIUU/Ua/Zn+W0zKyTvsfHw1ZZrFy3j
phiNjf+gaDkLEzWqzpWp84E11ajnSp+wN86yCMRO4NttmvjjUgMu+1L588Ue
e3USc/aGYtpRc02OFgTKvNwhzeG2btSRi3i8zJurPk29xjUHRM6SXcXAAw+r
LGgaSSIBWYr55uoYot/CcQ+cJyFXOMllqdm+TbV0PZXFX4Ykdj3hsZT/4M5h
tDLrbBO796Q2iewjG4H+M4m5ZlL6M0MkUxi1E+1ElwClnun9sbAvtsbbqY8D
H6KbA/P7DRlUQ6IG5qkRnIxCGdBqiKDICqnNuoyhjh3N+pUYq8AtzPgVK4Xi
m2ZbijrusvYkWet5JNtJMC6jLfbNk3JXgFy8I56CDnIIwbdE9EhKSevN1UTy
CmMT0K9bKqLc1BndJ/EldpuePOTAXUvaCI5dXKIl18hZo0o0BqGEgbeRPcIu
czK0EKccEyV3U3qC+53NmRqdN7uEpWvdjYVUFG4rbDU0fZ/X4JZ4OmbrHuVr
znEMzMDHVTk92AOv4+Sa2N232onTKSNDPC9UCqtKgIZjJkz00rdbgFN2Hr+K
5/duLmTDArc54uPRt94a9I0AR/Xq0DdvUEwk5MpvJ8IlMnZQEvFE0cK7i+xj
HzbGF/agntZXPX9NsGJJigJmXsQTZ/MKs1PScSZelLpM6+oEnsIeY1Nbin8I
y1zBqDqrzUVkB0IF4UoCcqjc407afoS8NqWbKmWiRSwgmxTjk5iWkT30Z3sG
avnZaiGWsRmoXbaPZHDYsVuFGQpArVtctMfzcVqxIfdCsIcE2ye8v3G77HVo
NcIPHtKgMw4QIHYncCvyNLAzYX+vhVLsx5IDxCENDSFjvfUJZKrEHbCfO8KC
DgewQXl3XgjHAFKnOu1I18Gvwc200zuOIoEB6wyjdkSneEJgiq4V3d4hH7mh
2ktA3woBW4gDvIlAsIQHcaAdre0ds1IXjVE02nRyVdx0v3dVCrl37p4/JWQi
ZcYH9OaRzs9n59F9DJpuiYLUZAsAaPl1q5W5svJJWS5uQbzoS0l13HmgbGE8
UDhA+CW1kRGV7qhrxNsQEmFafHrNti8fWxJ4/IJO3RNijmYQW2Z2khXldSeA
cb6K9+d/8vNHDel9+E/+Y8kj2fkbYLu6DlSW7LVo5vRgtF7KYopE5jNPHoYy
hMEGUDzibN4qwmpVC1XnYBTjB0tgsU1+RwxwfQSeW676GSs/Ppc69JFR2qeE
2PpFHI+Sb3MfR4V/enk1gmqnYv5pkwyvbU8reFNhfD51TeGqhCF3fpJnfMEe
pJavcZgqXewb/2TqG72eXenWJ6h04nMHzg5nZ+16JUjuEp5NfbZT4VUhfO3f
cbkcXDgodOkzCv1+5/inbH16i7zYUxVoXT+9P6XrHU18LWRZVyim7uEugjV6
sW7iqjw03EBqW/YajDE1KJNrGZS4ZV+BGqkgZuaH3+p/QCLVtRpzGbLVO5x9
szcQTdqpIf870F+3DmKfe17X3fqA9ssrtGswe02h/tjj6ALSGw+brqy6gZK0
t9p/JLhUtu4ZBA7SBi3aIeFrn8Q5+ms3+Jh+4kBuzRKjrnv7MorOpCbkHHK4
c+bC5x2x16sFGIZ9iiLNtkP7ckjx8Er9iByKE0E/BPj/RCqT+eoaZ3CgO1IR
gDaM/kwocu7DMlGIsndba+cZyfJcP84PnagdO+VXeXvGVKF/N6MTLWU8daLw
4TC87lXYuZ+20hSz7ofsFK8fykMzUkBSzpEPqUK9ZKghMfFGqUN8bygDSchm
x+CqFHyLGZOgojD+f7QPy/Y/1vb6drJm1MxNyTpyaUZdutS9mhMSDCk3PXUk
b4UwbqGxW+eRgqk5RW0OjmkNBvWPIWJ6RqIK0KPXwfseMFbzvgexwHFHzHrh
5Nqqqb+VkA1E6IhZvhhSvf72lBKY1SSYyEJkGZJl70bAJs9sD3qkPd670FbA
zv/EX/WBFEhbeMK9Ur/1vm1Aa7miaqRwfLDMHPBtv6ztOGaAPfjUiyHdt9pJ
JDM659c/2HI/Ix6FDDj99oTcVfaBw7cOX8xsYEcdmK6jljpxMfB687oErooP
Tx+Xk7ALuTkZ1CbTOSjaS0WU+TeznReFVpOEXIuq6nkkwfEPQQde2+woqne+
8gD7igEYR5vDtjChb58iPGyFlgmyjF+e81Kdt7pnFnGmrh2RpX+5SEMDTsZe
+Kjbl1OkhS5vYJbgrDJtXZqzYeEHdHJO1iOqMccRdEO4rC1QlsJSRxAlCtYa
NPT+QQM6mlETCfN4ImbtKCIxbbVE7bV3NolS02hWnoswQZj1uEZvwTiJ9Ulg
eQUiG+Fg9FqM4Zx2SRV2kN0yv3R6edVBR7biHY2gvd+6lCHeLZQn7QZx8ka0
+GxGI0UTicGTj/kzs9fL+97kSI2EpDHt+pdDO+At3lhJsWepzo6vFwdtX2bz
v9I2AviZOG0HUBGJKfX5UXhkr8hXwlFg099uW66y6uRC5QCwKKppiNdAmuse
V1o/RsKkUADxOAsc86caRWWG0D0LJl7j1RFWf32rT2p/Mo4jDxdkOLf650I0
3nb42t1hRGgBXUG2A7XbcKa7oQ1p/qV7+mkYNTIZE+mPZJqzid95mKqEP2bn
ra8mk5Zi0sIzKjU0Hghq2S2BKZvShafIf4GKzJsYKWM3AMDCb8f2A4OfNyJp
HwVFTzByRNXjGQkID6ZTZqM3Hq2uYKuf3jrz2Tv8vtCYsiH1urbraYSZ5z74
ivPoLzuEFhg7CieSZcjUgtOL5hEDYiq9t2f0lq4BDbgaB99VI7R4DdsUx4tI
B6b6YKkjVuxmRjVc+qeJZhpcpRb2PAIStXFnisb3ldMxdWpP4ftxAY/M0C+m
8xPbJ39XvOHlnkReXKcIoRvzD8cy8e4vVXTB6wFZeMpXTLx8sqOnZ/KPf1a3
xJ1AXYE/wNyRvBT0YkatpwLSruTYpLkgqMIlx0/5fiYfGzDykhgkdgg89KXH
NEUwRi5nz9CG3MNZfNxahgS+xE/YrudGj/T9UX7XJ6KcYKyw8J4WWqdPpKHx
0AAyKYeDRY1E1I6F4Ew7uJNfAYTteRcnKLdxmTjYLfMvq+pMwDaf3Myw/0XU
CwTXncAL5gzVJLtsglCM0a59s90dW1CRcydd+tprkctk2a2MZeWDV8nwKxoh
36ltufnkLQTVbI/b7u4tfXe0fBfnmyvNG97NLbkHK3FTnZbDGGgszITrT4a0
y/XLyNKXWyKEjz3NYiti0rmVnPFdJkiLVnorf0Qzgz/QfBupzlc9Z7/2bRN3
PhKOBxqbKPjtR2K0ryp91vTGa9tpkUwaR6EoIFXtDxucsfve1gwPgzi1Z7Gm
YtgCSO4A5Hw3yLzNNaLU+NeGJASatU1HRlduByy/9tpDWoTQVJa+Dm2jzMd/
+h6fW27D6MR4R+Q5angswg2oB8fqHH1Pc4bLlji0JwoJRwWFuy7uCVIO5yNr
KWUgrmiHfBCbC+glbbc4UZ4QH6YtFS/YJNt1ET5blIAMdv+0TK6RXDTTG3Zj
BI+ytAy+O7OfnR5NhL71bYkoFP+f3/KtM7eumZeyVI/ngFVhyve159dQhl7u
1ytkpe6OAVm8jolFgBPffOMU+KfXYN6yZ3lXhtQy6vdf+1m5h9i2IN6bZqvt
+T25O+GBDb/+ulslG+gWuIOYWDC2d2Ul9V9yFAj2UQCoiUKFD6e9qF7CEZAZ
68XLSebOhUDt3UlS9KLfkusCLN670uNdELZwsB9pMhhdP9aHHqGcegFLV+03
IB570A+c1rYeiCZj/8+Z/sdHT5UMJGuELvlGw2mmiwfDuBSNw5lGkSGBsfgt
AJxB7NBVQp8av3Cj7Ya+lY5yHUth9p5zYCpFyVMRZCjpthEAufDcdK7jBtqV
GyNmKi45x2oCHN3ClapqdBdsZSK9fpwB5bH2fttXIQV3ETbc0BV1A41zPnpx
H7t3OAQL78zuroMZ3EZQPMQsYmZeiz3T7rf+9+vceu4bRRU1YP14GLy8xwJy
IinqeyNSt6vATi0lEdONyxGvj96DfqwbJp5rd6mhw/lcJka3febkLNB2PGSR
6ve3zGmyR7ZtUouUCSKMF+5ghnzey7sqajnOv+1kfv6F8KlbfFvCFshDHo3B
i5OI8pL4QcLZHhz6vEkm/D4ZG4FlO+Q/I31k/l3YyfMPe5Kg0egdUFTf7Fs7
S+mL0RvrdRmmJpDNyIkCq/uViwM56cmOyxokbYYppSx4u2jGYZzvWFHQLrjd
QW0eDQb+lKrJgoWJqs2za2XtJMiT/XEEjPfIYe7TjnNZWnCtBcB1+m/oGMOD
hTFH912zfyDikv/68MufaWTy2SIECmUv85cmTYd0s6JJiR76ZQBUvh9wkP/f
jeSwPnSV8w6YhNWNpcJh5Fe2ZkQ9AYtXXf7LXhl5Gb+kQQYg8cAaTbBPIHuB
IKVRC1qRYRJIRFUuTmvpNtHF0eYPbuOHGz4MrlgSeanJmdwzFoZ2sGFFxgL/
JDEBS/gl8BUDE9S7EYLdyA3GM6IEv2Et5mmnHVppm5EAur3WE6rurY9UX6sK
WF3QEa8ywjTOB4onCw0gUhr/6qjX6AZvDHZRm4xeUfez4wLcoLvupevb/lw1
Yu/CtXLVT/mhFha4vsu/Nzfqosr4wj661LV4XPuO6qmeDR9cCwxw3mrgq+w0
bo+EF7Udj3a1Uxgnp2hOZMiFuCTy2s2wPbY90e+vLCJ4TKQKfhRFsp31ASac
5TXmvbsA/lfKfom2KRPwMO1gYQJsoQTQNbiCiGEH/rEjPAxlMaiqX+ULiwbl
0tz/R8AX3Mq5xyXwIxz+HfpJoUuzdRceMvb2JAiCYXPD1ojvXjXtZhEe+r5a
LssiP22ag0yo9ZwJGumfHPgJEJ0IkWTXTluo26PCHxoDhtZVS6DhHiGj4Ba7
5wQ+n1S9Dn/SQvGiZO6uSvxgMigQtD1XMF3pyWRnkr8zUcceRXwq4IkcAftx
MbE+Omj6CwgdAvO27d1+MowlQ2FiLeWwYF/IjbkA3thw2/YdW1ETwYl44d8D
BbOYkSNx5Zd373MRlbfw1DBTCkz1SUBgKv8gubLdOZ7nYO81BR9QF/Gvc3KB
1WGgZxl79ZyPrqvf9VUI+5w1g2Ij6RSKf9bxmlDWv/kuvrC+yxaM+ELcqh63
JgZ3L7HyoFQemaHF/r6CfKVDnknzItB11kjWnSpjnbdINV8Jq5qYEoVSjvSo
l6APeriShwYq0nwdKaJY09KDLgvfK2/2oZReGKEXO7N6nLQFFDFhWE6wJxOu
y1U7CS8z1k0ysRdGhnbK/+9RJyjv8hONxG5Eb6nu36eJP8LYqnUmmH0FVmKO
mh1gCXhZ9dG9LWuodHyUHK4MvZMk7oSlueCXHBuELqq+U4CXiq1DOjpVDcB1
+PbwL6bZdofWpl0hdLX0FKLJy3TwFlC5rNetpugnoj0H+c1ZPycq3FdVY08h
fA/UZbHF5RcO55zSfqNlo1aXIHOcmq0HUz+kGLT/mIlfUtEUsBJD+OFemAA7
vfqyADNeCC7Oad1qtxtf/up3S4GTLIodzfvTKUCewp309yvX3rO25xpAYXFo
cNGdLLAJ2Awv3KSUz7QC8QZsi32xjc/O++G8CLRfkBxBxSxOPqNyrEtTL/RO
IoBqZxVP9wdwLasFeE0mhW1l/LN1jM9Wza/hN9cqh6/R2//6JfDj/5+7Y+BO
QAFnOrAGAQMMu+yMyqnyG4LFoxDej0JLpKSCZv03xWFHuc1bFwCt0U8PQUrg
Cl01JcqdmoJrL1TZVB5vR8S0NxkMu/WZefY0zRyMielO0gxqKZEJALSa0idx
auikBlmiKlNFLDbIREoz+mXmqBBzD7pJA7KoUTTi3wXLxjzLchuAPbfbXOSM
jBz0/SMCIZpals4s5asq7Ri63d+TWOr/aK8lCf/E4iVOeDVtT+SqkT2xCZCx
iFrB0b4isw5Sr11ojDOnsPUBxKpNyUt/sTedU+RCzJbq6IdcHsVq/rLEWA02
vBCUH8YTCfrJPXa4+cg72+1KTHr8GUIVoPh/pftvRbFhq5YihbQVvM5alS9a
UCU5lkR/hWTfAbn0aXp2yd9VrOXF6K8462XalJr6Hu/1Yyyfg0dTmKpqhJAl
8AjMU8tL2wHp4xL3ByDgatF035H74Ql11aKvi+CfhlTZPncTHEDGYIAvF54d
puVJdn8uhHWme+kJqUJ/9TDINiz3idO1tqYPIW2jbXGsgkZ9/ZweIcXCyhHk
RNPVHLmhF/4dKwYzrEhPbAmsuueD5Eiob4sZsgEr0jF715is9hZAYiOqK4s/
yIKQQgeZon2S8gRO9MJp1cnmMgZdoX+0TRCn72p1wYsCMxZZza8RwNlPIiwj
HCxO1UrVEcOkylVR1iKoWOrHhIdq5iYWOMionBDwe/5IaCPqIqaoiyvV5g2a
wOkyXjQ9MMGHRFgBhLoRjGTu8oOH2AP/79hp/g2qr0c4pyI+BBtyRmYFMgbb
K10qarJn5IRcleS7b6ZNGLfimAyxehENtaVgwhzXQgTpk68K2BX+OH9OcrXG
jL7HoHEtG77bGdT+3W0IU74+1XaZXdb8jrnPdBnUV/VbZi8cmbqUFDSwX/ZI
mOc0q32hWdvp2gQHlLUE50WDaQHA81DiKHkybVwgiHNI1JqnfXb/fqWvvEnb
drW3SS7jOmB2hd8WlfgQy64nblYYVe3+3AHr0mY/wQHyDOQSWCGii5m6XeFX
IowZRQNfYpY3AA56Sgp9fzjSlOQRiIW+0rnCkiASTzPXA51YFkcuFAknWZDy
smL5jy+cTRKTQmF8NfsZ1XG9NieqWJYs8hHkPYGtkDCPnaBtrIDP8uMyzlND
0ARcMacxA1lT6KnMCq4kJyi4qbfVHlYbWdOn0vtKkJ4c3NoqMe7MrQvNbcuG
jMzeu3Z0rkEXi4TGK/wipVwDTBUuiia8G7znbLZDM6eQCnAmhQJLWwndvSyO
9aWZQHbl3AB87O6P81WbrDO46E+94ly6tk15/Aow/GPbVEYoP0EZp/EcNy+D
5zTdN2AxhGpd6Xyn6gl8sEhXcgnGDuI6pW1rDZYgvuK+NtOSsgnNDQ84gee7
ifaHbwaKGN5dkopg0eriTMKx6RtmDAITQTvIsoIqBYigD3ez7hmNmWgb+x40
V0YZ7W9zJpDyFnQseAXvaAbc2rq9dtSMOEO46mR4yQA+syUo+auICIwlbO1E
nd47ajuI9UIH8Yrtgf8U7bvfGO4B7UJ/xkiTnbNUipXNvfqM7cndXGo8crL/
5/rItWokYSllhjGqhCEfYUAzC69AEW3Dsq/6Lpysjfh6dbankMLUmd4KTzKF
zxT0U3Ju15amvXt97CWHxR1opLOVVZlYHlpoC/gK79Y5LCBWDWTgl32KJVnQ
PVpahv4L9N5oYQtk2ZDpQ3EP8ouN9MVYqhIJeghqfu1c/0X+3Ad14Q9cMYST
I+RYSXncvcc+R62lREB1fmakU8BO4l1DoE6F1qFEwDfEjlFxskR2VZDlq55J
/aV9ep1N4jZs7ozoJwj1UyxWlLTgg88lv6N/aRugC4WSTIzROdPWc7h6zilG
oNL1Qn6bJmMpppB+06HNtYWezGhtXOrCS7e8EE7/Oz1P4SyP4iQ8Is5w39B1
+olLRQky4u3gN1QdxYTyB6g9SPQdDua2AkVC0+vAQ/gy70aSpGxvH538g6Ei
M33puVQY9sJLNmPJxmUZ3QatL5yiTnKXMZUAiOguO6XjwdfS7yPn+6SUfbTB
wKkxtEjvH5hGm6Gas6Sn0HkZrXuRpPcjFkg+OcuZVpn3CsOM7LY8KfFmQUT9
ICl5HvxtiqpMSEBOvR+uA+w8JRzmdtVWGrYpzdT6BaOv4U94v2n82jbX7g4+
x+HoT8A7qLGkE7qZHX6odBib+fLNH3iHca+B1KgGFlB2hwateWjJqB3FaN+y
+tscqotrjZ0OjoHPZxrsagPoFXsexS2Jkd1JVdR/IPitA0U9uCAZb8LeyPvx
bpVNIRAc6H2oSD5for+Y5PoG1jgbWRwq0tP9JfI65LCr4pTqEjiANK0qyCeZ
ioDMDCoXoQspO+QZFRuu89Ckgwq+oLgr10IVbGkv/uCl3dO5vE0go4IntFQG
SiehWrRjOGK3gss9eEo/Kykj1s1Doyfn+jRp9O+fI5oXNn2Kg5KFLkX/9I1g
3nUWLd4Z52Nz9tJ9GGusPSyZdBHimnLG25pWZ2WblDKDN3Vx3hIrr8gdRdL8
NCd0HC9tpdV6p+Fo9DuP8uKQH5gdCwGy0IDqeQ4449C5TetV4zk9HqXboFO/
S1vwm1jJDJLWNroVxpgKq/yKSRsScVMawPwicIv2P3rDq3W1tH60Eoy26PT6
By+CnExeWaz9r2SdqwNyptkQ1z7DdLEU656v1KfdWOAqO58Itoa4M5Uzl/p2
ZK/6R0gfsDUvfo+nYzswwAd89vUgv/2LzB/S4r4CJDYlrPN+Pwa3zSI2y3nY
cubiLw5PuQ1F5W5hOL3LB5YTG8ixtKkdCcndYtPPRpggcFoIud8B94/0uDhp
RKJ0SyDh1IjE1J7EYbKiaJ077oENwqdkCTtKrNwGCaBNU9+RvxB3N1LejFME
CeYOUHlXqGuT5J/u2DR+7AyjHsxX9kWP2sXaucwy/zXhbQMseZIKeOa4gU0b
CTkXNpYaeTMKcwwSn8N5oraiZDQmmrN3fqY2FO9tnYbQpO7nh3qeiSHJ2sud
HGnn7rXY4S9WwpoIjGI6vfImXK544i5CSjjMmsaETGsxo1xkghcwB6ZRCR/Y
ziwNze6JLQKXoGiL6LKRC45ldhLv7mzjCUT9jGWERYt18ppXZz7XfO3I5yPZ
kQzkWRBbr43e05QkbC5ouRN2HCSdR1CQppCYHqqEF6IvP18jAdShzdQxfOUH
zL2AismckzxfgWUNpfV4oBBL/qebvs3khhCd0XG6Rwmofbwb1VwAI7cbrvFk
5JZ5B3khgMmJLafRVmKukgNugXmKmNoL5HZv44wgUEuN60p77APQ2OO+yEia
GmbGCNIXE74x019RaWws9Dxt89tEobRTi1KPQmjd2SXLlGnNmNrMtcAKVaiw
8fIHmUCj/R+y6UVjEi9nE8e9St2EHYVnQ7RJoup4vWv5Mxs4V+jqwve2KzDt
+3iPB0SH+1qYSCX3DIR9QmyZWcpbKtwpTDObyyI8HVjcMwUR99cRiTCiBhPX
+QHoL41zmRpaCggKRX2DHt83iwC4rc0mu3JUxihLVDB7BzcgHV4bqp8fs6+W
qTJOWRUFnJV4G8H5wWrvZbWdPuthb8vCz2FKnPOLH/BuFOBrkLH9Kn6UQtei
2nHVJbg/cd11SOV8vdODycPhVL5z5XvHRaQQt7XueJcOLYcrypEFtznXEG3F
dDXSyDZovNI0LoITAgVZtKSGQ6xnv5fdXFEN1tfSIl3wL2+qtJgEalKFeiNx
VY4/F5JwXHKl4Z3OW0vRO9CuTJi2a4/pZpHZC5S946cD6Sg1ICNZPoZGWva0
LSyBcNIf71oQ/W6n1VbSUlNQEcLkNR7fVykbfv9+eW0ewiYoRIosOK2YUsC2
VKcXZ3w0wDZr2HSB30+CP/ueiLowcP6HzgvkTXqrez+imHUuvAxd/dOBQN1y
lVDz5m4h57oT3cg/+F4nVLZ+D/LYZwgfD7DpF647yETvkRIpUeBYfFE2cqOJ
5pK8thCeiLSXyn/3jrZ8wwqWt9ZBzG+3WQw1AiWc3GJVrkn4haTWk8QtbGsf
t9VfwX6isWf9/BlxCPdQOeRiXuzLdBP1ITGrCnKvIgd3RSik9C3SZd2i/IoT
hn55/ps7xOrYqZ25TMXghFHP6nbk+EjfPVvw8q0LKDbE7x3ORvpcsyaiDEm5
Kj70SeistdUfRXn0wgedwIEXv+OKzCLDgXHT9SRg5Fb+CuDQznYjKMNGPk/y
lIQCxmZJHBMGTQCn1tvYTSEeKAPOobLKfPbSK2RYhxjDE+dCzFypzvh4LPis
PYNBNTcp+fZx0kX3J2vrwvNjTmTdRaY5iPGtgtln1VovHhdQq4yjWEY7/lpW
SuwIR21RyqusRwT5XlmwPiWtxoiJxcKTsPS1f2YvWV/x/aSadX01DZoLlg6M
N9nYeLSAw4m5aCq4HZdQ6dKDOyVZQmabI8Xy97OQpfyuRAvQGsgKkhlPuPXG
f5M11KTWJkaMmBQ4yV9v3afx1hm+FOAT8VSx0gQFeg8Ythy39HpWRO1AiRkt
tAaccTfNqtTOd9mLeHMcwnNWa8z35j2qLLwj06JePnl26ng7qpG2IBTJTZ5q
LYHrEFKPxyk/OtO5WN41/jVb0E6pxF3Z1wkM8FZEAyYrESQOouJpVX/EwwEa
meGzXL1eKpYbx3acfnfQ+1w++DkED6vAsyrVK+21wJ/Z9HPIE88XlU6PEmXs
LzfNl+hQtjeoS3SK9mRUV1yHlkcTm9lYUsLn+d9QvS285hkJmxfmR25tDfJe
zBIQYn94wJAPwEvQlPBJbrmlgfFSZvxyICxHKR6CkAXmqaKbumAb+JU9beUP
x3dNZQuoRgeQ9FpMqfAP1Mfr5Y7i59FacpoSJPMhocnwKhBStF6DmpPznQox
4HBKG849jBBFJwock8OUJjR+aBKRAd8J+kD4qyHEqtpWaB3DVcIGF6/yTPsI
BhPizJJ/JnIaxbbNBw6RILExWfyac1G6s4Iurrm01/ZxOEijGPbc+QFUnbWe
7LEq0XMNXHEtEIgdTgng/SACtHEv0L/aQNvTmvweKh4lnvitXuP0Ev/+Qlwu
fuOEh5YWJPat2JxPlSs3G2fTbb4mQX7jU0i6JyAoqmvAoXmnfCI6GvPhpk/1
0WLxKQbU4MeP0YUAwrk3uPUfbm2ZKlLpiuveeDjBc4YlqJSjtvcb+qpz3pFH
Yun2729Dti8VyTU870Uu8uGT4cBoglVBr22BBFFwqm80pU2jwdpTr1I4o+Fq
tX9+J4lPpkqy6UbqwWcqJcn8x3lCZPH0GfGEVxpFx9gItm0ajHniIUBtCOUL
Gfn43mPuxlZ22+pEJJNQOfWHwY9eUi0Bu4jQKPHH9DHfFa5FnWsTvvDjO8cg
h63xx/fZKMkERRYJ995FPNnDnhKaqyo0AguwgqE8DvQj/UFygmvu29KMpHyH
2z3ZzaeRZE40k+VaLGwhmE0ok5fVT+X7y+EFtLyisSRrOsQ/tJ02NxjxWugc
LWVHjSd+bb9kxoCkmHzd295Pv4xAFB3AHuGEn7+7/S1bC4wMZuoMr9ZS1KfZ
t5CsjqIts6r2xPGbfdP/CnRmYeH7Fnm+XWDXLYYAGJnppd4LyskXyYwqAFoW
MCr/0M5UbJMyB0xO4ww4MTRzKfnZ0HK2ybGCnAXaVpFNomUKyK8oKw0KIgm2
PVmxqfHuLTcr72ftbNWenF9Etyp7QeieeAA6d9+mDVEuA5SA1x464rU3ABx2
GX0O8ReKdFchL9Di+OsvUschNGFSAT85iWI5MZk/obHdDU+ZdVqcnLauME3e
1AFZG1zBfBpicjmVeOyzy9lKSz8UILaWBUFBKJE1tu3dy6rtIv5QTpQ4nyTT
vtiMG+blAaps5aU0wyBctwCa8qMakbuoiXe02rRLkA231T66GplZRJk9fRwT
Tm8tVnlgjXFBss1NqZdiXDF6XOZ+id5ZWESdvVrdnm4W/f7wQKB2UObrC9SP
cNlMdTt8BF+dPsKo6o0TZCXPrgA8RwnEjOChqQt4HjYbxRFM1/ILrvaWfxAc
I2HhnAac4aRSyKMLdyQBkvYfEZZCd1Mp159tWamB4jweGUHgMJqhapMR8s6K
t+BqdKsJsE7qoCQFf7Nk0lrAq4TvnG4YtuQPY6TgN+zdAcJcVByDlRvj9FL0
NdjlNaqfoKtLuivlIH8Z5XwQP9+GuRuSft6YjY/0mXMqVVEj6E6HtmUNbICc
GOXiLJ7vRGE9CWyE2JG9s5dxrgZ6leRgyrYsYTBl5JkgGvHstY5sEr3qKFTf
xAsvUMoIDwtFjsy/ovhxaORBxGpvE+hf2pFBP8mguLkr1pmKFAlxMH5wJ9dA
KfKh9xkSsQ0S15moJMrCS0DGXUowvlrrEX4GT21i7KvqzFN9xmgFRTZE+xn4
D060IcpCM0VvIxqzTjHHkXrn/Z7K0T4xCLa72h4YMDL+44XbfCsfXGkjj6M7
Q981PxsYmiBpoXFMQctbo4rlf/LrTpyVt2LI4hpJxt3mPaAz8N89h6PCCZbt
KPv24T0zS/feiD2Jvj+y9BGgLwjnWCYMMl+yFW9mxm/shqOvp/LL4les3jLU
5xZn+EVKkctyPWL0vpVJ5A/uDYnMNG7r9SX9fzG1EW2W8XOnTEjYAtxZ98hO
YUsKNDgxhF/gk9DuuowbcgQo/XMuJT5YSvLLDOqfCRc+P1xU81fLsdN/ZVtc
8tW/3cEcqTrZ2pdkXPIy2cFgE180Flc7yiPtcIFycUVzZjhSp4j2QZGv0j7t
TbMldpl3Eh/vchu3IeNL6QmFc4zaUCPk8awrIFv9D19sFsAZ4PO1ia+gSkYU
GatP7mw2kDGUgQ0VZ9emj0S73pILWaAcdl6cASFqFrzN1c3YM2TTtxKrqXm3
n700vSJYOuNxBrj0HT20kZC8Z9WYxPRq9o3Z7EtOhqXSsbBi8UTbshuoTfF2
93mOrqSvmSIkqH+isYk2cBq7Ba+81mPAl16i6W9sPA67g0Oc3yYZus/qIOmS
sZstkbfdq3r6KK5p9gro9V62H1o+rvxdluRIsJX098uOKfnGEnxjBtaps7y2
689sj8ZRQHjBBW3gicDeP9cHlH4gQ28xK3yBHN4t/6YphkQ9X6e6h7Ke1c3X
eFUm2ofaTPhttN3CiUMNBSN5vNGFWL0dZBkOlqZxuhyXBCpzGCB9AfyGO6yR
/XMooi102jJSFp+gHLA98mDz+Q4esOgac1gF4yzAWfFydM+PhlXBXX6qZ73m
UGKLYq9Ki4Gl74rzNkqwOtkpiMca+L/DT8SxwfDJNGK/YGqlLi9XD0uJ38Tb
b0xgSd4Kxzl2ZSJkklTcPWxwKQB6MXVbgfZ1A2UxkC2zMzOrbBMUMAkdrHgU
w0JO8KJV97OuO1ENlUR4HCX+Dqa5/TDSrRo1Ixz8oAWpAXuiBhoGRcIPPIhZ
9voFVCP7+1S745PVF05oXqJruoz/vcPcZGzAJApUwLHmhkeS84BrOrg4lJNe
cWy73QX3hR/ezPeROhYGtHav0xmTzz1om0yfFz1lAwf6+TNhmtPJQFk+I/LB
kBrsFvAAZMXG4axP7rKm2f8F47ZkwuHCj8ZdYrF1m0fEiYF38pwITwqFcqjD
MRZJ4/95sBjXhPAb5m7b/J1DDPd4L4e8F8W8y2swUHlEtUbLomHnM0p0wM4K
9t4c92X2jSaJSbse3l9weOn+ueS8r4oHNZ7CUP2DGC2DtRm1SFaRjnUcmwdC
WePP3X6p74PiXHyEuctS6fglnsY18vsYmuRqR0ideXrD9nrurOMYkfzbW+ag
4jjtK5/sfdxDItm2LYIe/lDbTtwGVf+hBSEwBv3eA2rDudHfKFcC/MgljhFv
S+9uEO3eB6VRSiAKsDWj6vALKBHzpfkh/RP+lTJPEyEo8EsFuyUi7DhDmOjk
OFgCnAGdeUTd8wNNQAcPYDV5yvWaqSf6NkdLRPb6yTyu0TA1XuPSp8ZIzpmj
FAoPZgQ7VfajyeZYKlYaqW4Bm8P3QD1wTvq6WGY1+tUdlP9OqHD8fHcNJNLJ
dRLMDcexARjBY/B7YqJn8eXKkWq3TicrWsv4qfMKAj13LbDNFKGJ6PgFceS6
j6BZ1GcPA978d2LujJ/Wejsi5DqeKZ2al225T+6YK6ca6g7Wg4I5BxUYQmRU
+UXKbulXHylITOFdwL0PMm8my7lhdeeHLoiGeQREhetQEHXukb/VTn6XvFuE
flfttHJlOHd443c9d0FCPqkQRgk+40nv+b1rJ9/Vy4zX01ducQF/ZzrEeCoD
CXY4WQOw4Fmu0ebOD29z5wOAz6/kIc/1fgcWJ6VV979LoJTXMoj97opiNdhu
VnLEWkJ3ifuKDb8e5UUz0Oe4FhuCGW/Gr8j335UZrGAWJ7qeyosahkRy3qmV
CI9/iZackKDy6oek1JQsxUt7PEzIeccblQtW1h6dT3TvGQTiD3PJSoFxEQYP
VfQ+TD9ZUd1LyD4r5lLl+6tHIuA0bffmWSB6KT2Es3tFue6imrdefzEwfB2+
s6FxmcaZo7nqaq2fspcWTsNPHNaoTjVbWzhVrk3p5g2vFHcuiL9BDZXpex4y
UuDztluV2Z5jQX7Weou1gp7XunoiXcybxxm5jePmL5CbG9ZN8Kcb7UIjw074
W09n9WkWpZsesxDeXlpe0Uz4r28xwpsAEkVvE1E81nuo6YuAiFCi/oK5kNyl
77Fu6NNqFqD3H95mWei6tmYY+5cF/rDbvBpbGbSbuBrbUKLuB+gR9NCKmezc
ifGpBrgtIuRtz9oW84OloQ/5QVndn+fL2Ik/KbbrjwFjb+VAKFLZ4PLvCTMV
u8gjtVE4Hg1/r6vUHB36ynALyon+xAmv8fF63wcJYdPVlKUud3BjrgPqHdD8
yAOEcP02Ae9UWDjmDclP9DGfiTct/QhSnuVD5JErK/SttGZYwWQgO3WbIy9s
GECPDmROEfrwX+BeatgShe1whnbogI2SHE9ZjOkm00YlgGDwftzGKguAyioi
+vwfaLUG6B2g0khACKdlfi0os081iGAPSp3ZvXZB83rCxy71fwqEEwLGCngF
24G6dDT0oOpHD8BEiu0DGiOvIMNEREDumnafJdyWLiy8OzJhaAVmRFVgckFq
eVVNsCe9xEV+QxFki07i9knu1hqXlHBPvudbav3Z1Y+cwzriZS0tX/bvbIJC
3GwWYYl2baZcCOvKnTueX21NrVKimrzD6NxEVPTNgxuO23BlWpkYsf6VYw9M
miivsl6rLT3FMMUkpIJQOAqSMOMVUuAEal+3UQbMfpuwFHBQ2o4tnwJnosRy
bWvpgeijA40nFnZze49LS8+NG/b2COrr+7ekW+V7blweGpsp8KSRCSwNyJk5
thr1RiragAAxfgCeYAYv0RGOFDETMd3Hjf5mVt0F6rK1UPsR58i3d7Mkkhqf
sUC2PQIFNlIYKd2QDkj/buHgMA8Gqgxlt33ESMOYjO0iAwJu6v1ZbYoDJv5A
oF1MR/3dt2LYzGuGmMFC914ecW0FVYuR9/QnpV8TYi9u+a/LXd1gDRoVvmwp
UMNaoqIF/2gEPBGBqlZtUzRN58wo7t+z363AZ7qs9/k7+pnVLGBjEPnVWk3x
rm4W1B6Vi7NAg0x3vMWdwm1vuxHncDMenftbgbEJzJgElSB70JbwuPKREQAj
hzjW/w7AOzKOqt+8WAiiq62pwGfh/jU+owLxnYsvVCVkcI2yhCfNzY8tYnIs
0j8zTxVSNA4q3xBReJBCl5BMsCUuHWVh439icj9OWHADzAY7elaTLUweFv29
QTj5qd1h0sKWbg8KmtuP+TdXBfmeT4xDNXGmDgV0BuA8LFKcjTF7rhuvlDt5
ehSe9VL3JxBKc27gZEIsQUREHXdOQvYAlPoeL7HvErirGU4hhYSR7fl/v5OO
JbJJLMq63RIclIMEtkE+j6FW/p0ZoucHmutw/7U7kLvJkqGvxS2jzMiwvNaP
sEckpgE3L5r6MZJ8aOLxV7dsLkhF44KTaQgi/8N/TFrVHIgwwCLlnUs2Rs+B
F1jVVZyPSzGuIWMb0F+fFY4unZCcFjekaCveQb7DLeeZQ7KLltLC5pLqMGHE
r8b6PIkhLCLaqAQm+0IrXCI8fy5Qv7DdRkh69zd6Dg2l7luAyI+zUKeGfl5Q
MycTetjsKo6Z2T122EzDeXEvl42uDmnaLTeS2AbBtyyiDNnFntEYWf4W3jNS
35AFTu29n/t4DI4SbrDECSc4eBKnpH/nPwTpHqVH4PIeiFrO1EPmiFgpge1F
Apbq1qFkz3UETkVVfIlJiHLfDbXZcxxWoDGeV5XqP4icUyA2XRSD7+1H6L1k
1evHEi8XjVhuC0jfDf69dNvt/anTFVlvVXerQzD+lwm6YyWPctpFQlQkwd4m
UARrERYQA04NB+tyY6EGJBlmS9sAA58ybb5H9P2L6QW5H1KqZsjLCI96LG3a
umQw8CbZw5aUTb4fuyoR+2uMsouJRcGfnUA0vJs4+W62bvjf/nKGIJru/1+N
DBIDgAFfUsaC4OnMwhq6RENjuHfFtusHdOpmPTRUxXcabMj/yhAb625Zk4m3
rvQTZ2O9yls2kRNJ2BesyjgtjWScmSG9LBIvKHZjRgC1Y14RD9kU9WQHeaP+
bJVTGzg+FBAc0hj9Q+Ray0AdPR8BDsM2JcqSE860U74skHVNIVknJ0OfhTki
WGQmWiknRgNy/cXDYRhnt40/vunTpgL8iiz346DQpvASuU8Ll6L6w7mmhjb3
Ay5j0PkBi3Jpfs9XvLLhVbBhgwixVEiegNAXlDDTJ+eQTZHhHCIpoHZ5NVho
zfcU7KZlcvqgTmKRrisRO+AhZ8jQJTzA8GqWb76kETHGAKKJXrm0KifD8k3Z
DR6AWiG5M5NRc8HXUtk+v0VaC4loJsZfS4trDxwbDWswfRt2qdOMR/XW+3gs
QeQHySmmAR1zkkX1oMn1ZrTu0+/6c7KL9sys5HakCLhdzm5bAPuV8lnG0gNE
WjMsQ60IFNlU3RNigxqCff5HczlyRvCDJmflFe/I4TiwXROZP+FgG1ocVkxe
1XiV94wes1VRN28ZAF+54gJrVWs0NJbDBRI2RJNFvAGXjESyag73Lpfrjh5E
zfiz1vHiLaegRKUDbo7/XEcMrQV+ggNSD8+xof9Wn+asRYohjAJPizQEa4+4
GOdIveoTK1APYN5NHdVRNtoRtWuVc00IjAcnGzbIjYzLcWYTHT8OADiFsGl5
0X+CNAJhBaVJVPDPkE3+B3U2lsCKnfsRdXTVefApQ/Sn6A+qHBJUdCPD5YwI
yRbMsMQs9dpADUarnUawBlwdRu2iYS2o5bmHTXDj8ackdq/yv86aTUuuUKI7
xBDzZlU3QrCDqh3mrJ8rJYjb6Ai6LTKXQgx9T2fp6a39HBJn+ImLE9VsHv3e
b1FcNJG2mjmrt/d3nUtX/eObVUubtPrFVsIWq6BG12S4fGu1xSjA/DnInVGk
XBTrH6KMTR0SODBVzG76D/UxDGWgmi6OvzfXuWdqv8C8mzi3jsxV+WlAoquO
5SqQ3eIUSmbo0zgpHw/yOBqnGBokmPsVQHn5HYpfvf/nJrzqaT2WOY+0EwZ1
D24/DyJPx3AtXGf3/209+yK/VcxqGovfQHCG68ttcAL/6kJZKaSUIK5AZDHu
w08AKXKW25zdVbatSXrMjYsR783qADxNx5tqYAWrCxHSyHP0HhaSejgYM/gc
nv9QrYhhaaMvClqFnpNSjvgQG/XVRfyI6yjrsBMzU3NIbAFKr+cSbmoS3cH/
JgCzajJkGJmZfD+Mud2VG7OpeFSL/lHU+4wkmuVeFAplDmKuoyvMTIevRvrb
z0kbzemIKei/gKhmNqAklr8ZydMqOL7l/9jZVTnx+uWtkPG1VGDnV+jtsoT0
J9NLrH1QILeIKmvi0BVYTSqEGh4sn+bD1xUVq/HixZlL7yXM+puZO/2mf++9
aczqfyo6caAXL6T0vTpqeWMPi2JqSxRLrlRA1fF1/O5QsgSCsnCR0StAu5Zu
s7+hRq8ucSSjREzDdtAcZAG2QIUXP4fajvddMBhKYdwK28shn19bJ4D6g7Up
c2novpdlz2YI0JUPVeqw3atbgyjXG4wPccDtdk1ZBNvdKhAtARllj4/lR1sS
STqEifW3zbQFX6vJU6pzPKlw07k0/ZT3dP4GHnrqO8pf/nyWx7ulImURo/RR
agGLKnjbXMZMNsKe/sIA9b+3Gm8hMMH9nSIr+xdvd8UPw4odotUOnQ5Fdru2
UdP4etuwNvSAu5L8tT+Kh9dDtHGAcjCag1tj2XVO+dg9tE0YYwQqZp7DS3G7
0Cv+SVLsVFS3iL51TDciW7M2dctSNzSWVlGrxj81dHY42nrtQQyLNTpZ64k8
GOf+sK5hyUVr8itCrPq3bxtOZOh1HVX5W4t3hc8bUcZzPlnPp8pBjisOSUsZ
9ORkENcvr7zHFNfX8chdaPxJt9u0KPI8fIpgF7VTPHeObdD6ypDdczU7AutD
ntrul64aZdSAJNzdUMYLUDvXGOPbU1q3sIcQYr4vinliH9NikHZ5W0Jmu4/K
jbcEhusfyylCoGJeprWe1xltzn/Uo+XFG6l5hmImTrpWRf2Rb3IjqJWkZGvs
h4mQrtrW5OzvPX09RuSmUv6n2BzN8Ylrb+hOZ7hZHNTY/R85kq3oOtqUBsIH
kLNg1Uo70U/IYlEvJhmajwhAzsud+NTASbUt2mlRZL1OvE9LFHgXm/o11NPu
rUH068kpgUG7YSAcepZWtcFTdBeK1kuH1h8hdDhML1Ju2Dk15KAx7qvVQpdC
jxLUB6styfpi5j3tJ0s/lDh3P6wxEU0t3wHxnCpH+YJ3ONnL5KtOioPRJouX
2C6eOWrSPIPci2tihVt+Lt0in35V21d9dVP/LxU+jUUfBtn/XxKzLORAesiM
1Hq5TXO/t/a+K7lThaAM/TZfCXNsfisIdrBHquRLPHv2bOLpI2xIn6KS4coe
ctj01YxvKvc7ugVQFI6cTkT5jCUkBQAqhZzpD5MY7LC3PwTyipz6wVM2HmPg
nAdPaOCpAahgPAemHElrH92dnm+yowBu+22P6uus3FhCiEec75qwBghAKpdA
krGo4odQPyrhjW5dl06JZyUgsjWF+4s1ljLWHaeorU/j9QXTqXMw7BA6CMA4
0S/xSuH4CIJ2V8lVHsgxqRtKGaiUCiwXk1CeKlIIekQLGBtGu9OxUFvFVwcB
2WdBMf3qoi3C5tF3Vw8sCjXBcqn+uqxtjmwVyPRHSBmjv7nhW5ozjVSVLj4f
FEQql7YiQwXctkE97TRDS9+M4Wc/mpPtLFFN/JYN2KHOZQ+O7dO32koy/48j
/JbqjpvN0LPbb2B8GTiX+DHI1/oHZf0giJs72K/OAchb/WmlTuM3LqYZ1wBM
iirvImWQ6yijOdofpb39jIJxT2VVwgWzZ6hltZTmh03/8WWIUhlpVReQtgJx
7b7yRhRxvL0FW0nbFYYsFxo/E4+2mA6UUtcgr9nRx9PdwpxsY03qaYmIDeLY
NwosZaPQujoJ8FDgpKq/MkZbFjqAHo/vWSSyycCYRnkc48ECyUaPH0G00Ep8
0i9fPJUxNSE1sFzUDt87ltpkqOpZxhYFxXs5BLM8cJtLJt/74AS47gDSPs6p
oBxHEp7LxtBDXA0Re9zCg/2qlRkfHEPCSR75Db5QdXr8HNfvo6/2nS3vxI96
e3aphDw+G3dKDa7Ba5hOsW260Wj4vqOZxzSYLSNfc29V7QuWcSRSBxWePZzD
HWGi5mWrp26BM6i3Q3eiQ8SpnxlctTkK5iwzoUCiBcUm3QQdjUcpUuXwTMKE
SwrZQnxbVGmKosb0MzVOyaHrZtLDsZVuhJKBkRr9XpyJARSapi83dfoBgOUx
YFSGLZDFniU5UxkwwKQtEeu0xV0cgz1aCFiq9/gt/8ET+3xzI+P9kYev3xoV
8wbuna+9YwMZ/xLGF1KBBawy9lDWBv1tPwBJGX2KjmIH+asF+YwvsiVEpz2j
eKcr6S8waKw1Bn9yfUAJKHp0YuZQHeApEXeMi7AryQbNhHdTUt1eF0ypWsf1
VahBYzK4E6Ed2muPlFnXQ67LIqRnwKtubVHBNgejmsTPqzusK6jaVzQdHlFZ
uldiYJTTIgyFHa2MYVNq4ro/dV0Mrs+ZTfoYm5PvuJuBfv25+9HFft7wf7uh
tsTGsZpj4DMD3tcJojZqliUSs+0X1cyMGO91RhD0Z8o5pTMRWirEAVcFXTxC
W7NNItPzkA4iG2CUwDlGeGMfkB0tkbDEcc+WU2V/r9zuweStfo8BPvvJ8m2W
VwHWyPBzZ0qUXKhpVjX86amTntczEzAAc45W5QWsYD7rLJw0DQn5yfyp7Vhe
zioKQ0kbjPqKBXN3223EvpvvRZYQwLSHVyfRCz63r51ybpPekoKpb821fQ3X
hMDQdPhgu87n33Jwd0l8m66co2TlLUST2Nx3qMwZ5AqyFCGiFm3mn8HjHvyF
+Bz+69RhozRp8xc2Hcz8edYWo3/k/dqVA/0qdUEMEThOitXCQgxiL+ewO26m
jeDf8CItcASdZ3LVXyHQkZTrdw0eC2dzBv3x0ya8Y+MTVnzSka5TyjWHNfHd
0YYNCIlLiDGcrDt2LsAWPcB6j2GTNWz5LwpPDb6O18FE8xg67gImwIeXTdWT
PO+epibeOVVpQCjWvUyDn8mxN1qLp9lNs90CoGNPpHPj60pa2fUq1khHF98J
70fnwILAw+QS1KvlCI5sxo5A8duUccYqwvalRabid/sKzhG6AkMC3RX6b6C+
kYz7WHwABTZSB3G5kQGmY7gtrOt6lI19GAUhKfnlKBVQ48P86BRmCXbFGYgu
msGl8PWHdPj85/FxA6WHo8TWTOIHVBMHiuR+30lyOk/6jAKorIrsW6KORFhu
FjUED6ETUhUHZRgIxKUfIBJD8RNsdTmZCZEp9M6yWFqtsOTxWB8SLK8ZvKM8
eORGXN2ofFlZwUOdGcy2SQeloWltMdt4SpOr1qJ46z3SuomlRLyiWCkmS4ES
Wx9XOkM3OA+7LJ/2qsA5D9iv6wPIPWysZGuNJfIYGBm1eo6rxRox4LB6XhSW
DR5vy9sAmznaqUTC4W5apu2Syo2jo4YipGH7wzZtBLybg2+ekMtkxVObnNdo
EsN0SS5nngfTzeCBLVfEf/gjE0z28MeOcu9TW2l485CFa199Zd9ZtB9hfsUP
N0Ii0OQ47i38R+iWjEHIIKiCt8dT/Ek3+Ke5epv/wYtIfNDCbceqVuoh2RS4
O2fUGk8tmHQKObm6SrJBCxBbsgGyTcKH0LjwSYmJ8PbFfYdSXHAXTIIVuYyt
arXFoYmUDqJOyXtkcQ0WRRiT1o+r6N1QlnA03OcvigRGbNUSkUc98Kl1KwAR
3l9gmZWquC54uBq86ofmFHMwEfABBcSH7CGtXG47juSTkNg6oTp2B699srBV
YJBvUDVwp4O/wpfwkxF+NDu9s69N5Q1GniblZS7Yrsr5pBpD7KMfGSPwAWip
dXuhaLdeMkFjaecz2wcoRWuJQjCOKWnUK+bKv3wXX3CM2gGxxwDJusR/P5iB
xSVfg5uOejh0G1k9EGvPr7h5WSbAYbn9iLZs8jwZX+GqE6JqTaF7WpfdLiY8
Re76l1o9knHty8EX7fXDjr4eXOqZInE6B0zjAh5PwhyPKbGwdMcIW5/RAMyH
FgzAX4kmrkor63CXUMgtwIWafqp3B9zIyw9dO1ozxt48hvEZRTXG1VZSCE8M
a72D8CIzyoaxJSZarfPTb+IdcRHWBp/OTka7SVfuLMTzy6L1NQFR2SazZB8J
SAWBKJXcsHXatzL4pUExrAMpdH6OkbLJJvZWNfwYRDx4sNhsfr3xjiSYZW31
ox7C1hBrZEKKyRqR33lT0idpG3u5ncM/WAus94AsxzUz+IsOyBuVU2Ov27QN
jDNc19pH1sCk04jBfKAGKFEpbBftM+KRM95DMfBYA81AhsFq13DLLUuOnBxm
/CUQ3NAd068njvmixzTRSE93du5PBLKfQtOUzhMtyxAFs8EVSfjycwHbzyJ+
eUmLK/W3YMk1TJ26HNWpyncTncx9lrf0ANy46C3AA41VuxahcvAMVHgrpp6S
GFldN7srmsW7GQvpQiL9VKEp0Dx0lK700pwEBYs07h35K9cPtj67p6W9OF6Y
JFIMgCGofaQc75FvYdYakfrePxokH3j1uSn1xU8r59w/W9QgCptVnOlN+MmW
JSTNvkLWkAKNoJzrfD+zU8ONAMyHWWUHbWXSwssyOO/6LqZ3s9Gg8xfPAawn
cJHV3iAUxXRdWYlHceDuZsjA94UIdIsbzXAS4AYmCm2+Y06qwSd898T+T/l2
a9t+3ctgD5RiWCC7IbsowC8Fx+nSLBemZQBAyp3NhOlLTflFmpARSg==

`pragma protect end_protected
