`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
OSwhp/A8Y6Bx+Bt224YUWdmVZGNLoVydvyi6NaETpqhIKgiSrb1bORhs1SJgmGML
IZMMrx/eGj8LAp4XMBIB+ClSQfaYARzh0qdaSxNifSK6DOg1A2lizTTKIUq3pYra
qOM58A8K4z520wFktolF8XYepjdG8F6jH+Kf+Ha9suk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 26576), data_block
fpPEDf2iRJgDhVz+js7HJlJUtVVgIdG4uvPomasbD3i+DATJzH/nxs0I7mQI1N3c
rXSfHFB4UHHTIlluJ15rtNf2vO3IQtAPOqC669fVOxTHfbyJKSstFuKe+PLLjmM8
gR+9bk0z4XNUZags4/EogEdDZL2+TJBUdX2zcgjfj2BoiN3flSRi6fmJOJ3OwuR9
MSqwUs8//NMXz7qloapV+LWiLZOp3pLFBMK+yIfVzQ6DlrRtd1kZWNh51JO86afo
E+8xf4PeKOHGlu44ZWVYXtW3GiXCco+n9Tm+rDIpqu15bes8eqiERVhNsdp4kizh
OiZpK1ujIHIqh36QV8Kz4KD7X1iI+i6onvzD/ln6hmTVna1crozCRMbe3bQtQxh/
u+tzkUySkICvSDUE/zeB5MKS2jIZCaM4KBucOB8FNMS7IwWDPvrH5SVZCiXbUXsb
EIZDeNmDuYzucQWJGDlKXNXF+SjgsjQyKHDyPJgt0HKCU6qEGAi2HhAzR9D7vPAT
wN2k1iwktg6rZs7n5DPDWLT4H/llQ+Z5GObKK7n1YuQG/mC0mgrdEEkMejyOET+I
xTmrB/rUvs0ZyKoKfJsSSLslV47qEWYPu81TgtO1M5u87dXLHg1bjBZ0yuGsVMq1
geh4mPpHzrxn2qncYY8lz/87mjfr5rBRhf7z1Pvzmay8KLCac6UIoja0PDY2E6ZB
LzXwsko3LZ7AEHqTCMGUOUoYW8bRybrrz3Kv9fFv2wGqT/TXDYHRL1cT8pm5VLIr
ATd0EGhSspfvXn2pEVhH/DTSvPUVu5vGYgJrzSXQO4rlkMC81wrkDraXXxp6OKSA
IAIygcC2x5S2CI/IkpRu/I8Oh3SnDt2DebJL6lcyxs9LRkuW8/lH1/ah+Fiyn8Vd
cGOPRUgGVLB0CfbQhWcysNMVUc+imtimQ0c6Tp2X3H6dvYHciBla3XuOweio0zDY
OxfzkzT+oYBJ0KeoJ9o0LJCd/AuCbHeq5J1aJuiDEtBQEdLxzvNikTYMyjcmY5Xs
BEgWmoiF6/eN7h7UPaZsG9kizW7M28u61YiwWxIEkMfXlkUpgDx27o1hatSq2TUK
GSKIwfkW0K/xnGabforQ8pbqXvznFs2Sa6bfR5BpanmL6sRINGN1KsUdMZoZkpTE
8tHukskkv4t6JbfH6wmFTOsnAQZP36DVOwLG1MnHgwPot2FHOHiWUekn7JlZ0c2W
RuvtCGVTu8AA0D6l7x0/pcnnkzKrCF6fMB8UQhY16PTnTNGeNaLf7Dl0i1qXQpji
OW84DfV4strj8EDX8qdz4a+QLQ37CLnT2mxn+5PzimGK7Sh2UAtUx1e599zzUtaH
xvZ3vfQIn1x61EDMlis5OmhSbTpPPFDV2TC6FZ+WZOpBBlH/E5Tbmy1Lnz/Gpurf
c+Ysked8UQVEhEaix/ba/ib7xQpu+NJAf59WS5x/tMknwMVisDVDqqsey+A65ac0
0wt81Rb+PBif+zNLab7q71tQ+yvLyWiu4zPEgcr8MOnhlzpCzeatq7L49BhgVp2R
grVkwQS97TZpmr9hUoM04eVj4h9KlH4wgwv1vLDpowQFVKwq7RgGs1XBNwx/7ffs
jY3lczejmRsWZesA0YOgLuH+2jYBSenZPcEAcpweG2kQhHauZQcarpREjP+uFrVj
GrUnl++kBGS1d7ueVE0VWa0d7lE59SYb8JjIugWHT6kjkzuN9SSpS9VuttU6w9k0
+QYlEukgdRgnSubb1kZEysITWi33INmjDZnj0N8fOom8W/oCSRRJum+RAxqzQKYa
O22GnUueJpawCeFul6z8nPefedk/CU+pQoWrZUYebst6rBSYd16kaSF63fCsAC3s
zxVYeEG3qyWK5XHRCmdq6nSQchQyX1/+ggjAN4k8XYI+a5sgT6B8IKcczYseBc59
HvpyidrMGiHaBC5E2tS+OpeB0tqFQQO2VdvSRUh1OFlymSNFtlnI0wB6SAWYM8o9
TAq6Y6zgoyR8m3nGLOldc/HtXYXwJw4rdpEcrwzJFnk/IUBf+1iw/7yqvmOOu8Eh
+IUe1BsWKpA27w3eER48V+lwH78v/yeJoGZ+LfDjSTKgmXIqu17bpkAXVyLnWOCb
yQd9l1JHFerjxbZgLTQGBjrAyfXtjNIdl/flMWq8Sv9m+ozWMyxfoJeT1sU41pJC
4yNGLqdklm+p2VLDblvpcegJ1EFX+27Db7pNsa3fMCrfI1hyqDEVyedpqwIvjQ2u
0zagkTU0GCw0AMKR+A55xYkFL0xs+/XV9c8kB36+IGjWVrRWV0WW/ZdF0Nb+WH3D
ObXySXY2ojCYabTarh4w5DTFOIc7Ji7UkWeO9bVwqCco8YlpzbEw9ps0vNaGqTkR
JxdBg/GnHF6W2+RvTOO8ZmYvbJvZNr6gsDlBDQdxiNTu7QffNj/o+wwUFdea9YnF
QFfhWYsaPqvWT+ux/R/V4YLaPJtnNQCdooIJeaEoXqCiO+DdDkKNQnwCr8Cy9Pnc
F8LeRN5BVLioMRdPGSRw3cbeWH7HZKCCaKP4MTJOZgOicZTy7R44qllJ6hlP6/lL
qnQuZ+KmzppED7/QbfFuitUb900D8PdcE1NbmIGMxw+LBpvsQ+cK7gqD4FX5NyRf
PjFwO6ru7JSR+r6RIA3Ug3AB2g/kMguo5DnOECmPcqqT/tXFaiPk+nSvKfWqfUMe
aC1kB5PD/QkLqXNZUYg2c1PNpUQ9mb9xyHY76ZxrqrsL83h4yzeI66Hr+F/jchlz
cDjEw6fhmVq0+Ik07uTdrsudB+Mp4eccc0AHF831yV9BsnXZ9eyI283V/SYZPiAp
0nuTVcAuMABImHVlWWqdAT9cjpo5wAI2D1Q8RmbDiBWyEWFno1dMo76fGrZ5pqUf
+G5XdAXgQuWYdvyChWWDxejPTg3rU4NG635lDy6qr8M2NKbDVU02EWEry9M1qaKT
iBFUbG+DvRAQBXQ5c7DyKlit3mSiUFHztHkRKEgZp0LBF9SA0dEy+BUVOmZ8ozW2
seo+FxmwH7XxhTuN95+SYTLXKiEyIMNegO9dzJ1eQyFo9Gni0RHBi3My3OjFC3eT
DZgLCgj5kIfebdflMTctlGYICUiyU9bzIJbR9Er4nwfnJTZsCR0v8x6QVNo4/80Y
n6Sm5VUqlUNu0DjRRNknmaK4bzx835yAWCbRnOdZD32VjKIppSEfZdqKPnGVx3st
b2l3oTY/Zsn61VzPpGmxUsctl81T6ljWBG1sGm78lJMFUOnUSpSHJ180vJefo0C6
NlN1nRcP0AYXPuFdBqQBpEA0rrIzlWjzNLmm9Q0QWfzYbdZ/wSpQDbNJuoU69jhr
zjH/Ndnij+pDMlP4W5ly4LWg3ZLsn57Y9VqYaq63qgR6+1jPCOq19gfacRjSluJm
NCApZS8BzD6VL+eQTRW9paSo+5S3mke3IKu/8pN+Ln58XX+cmthpTT/SX3GClJqj
Ygh8R+h76mghafkyR42Hy/XGhByse0bfZuEDSKNuAbYp5dTC1Mdri7Af2rz2MBdh
084U83Oo56X38WldiJgY04VNhXjEMZemRb4R17xiXcmMYIVIR27qjUyhJIvlVZNT
BJ0qdomQy6FP1yh5RVGpWYpbIf7/hRat/6W4OftN6WMrp6FDca8UYeaRyCPWB+jD
g0Fwfh4MsXBj+YSfrWzuRlO2RagxJYkgttwi1AV2viddqpo+QrNJijQ1NMzUIxaH
k1jmCeH5Mz7xxuu6VwzWR0i44zW6J3k/FYpSwvJFWHwpIuP6xu6dCC3VWgSUhtls
IBMGiV9NrJyw0oppaUV/kBUJP4ohatebMl/jF/3XozaK41GQ/Tu7HYx5nXbaider
Afm/BEfHEJiuNxUExn0yzhOHkayVGqqcbNdZo9J3LQgrYcA8YAYAHtp6LGt1XRet
cRP7SZS6jyd+80aVWYzALRBVqaUSUECDnOjmjLA8WUfYWR+W9hbpagdBs9C00ZLd
SesNLhAiptIz73wCyH8fVc5MlaVmfOkcoSGhwsGHRL+pSoVxBU+0HHpswo2xeCAi
8lRELafFZlKqUbZq7My6E64AOP9Tw/IPGsm0DDv/kPSKn+LLrnOp4+woOB5QPKlZ
ZbNsKiO7dI88sM7zgrHLK/1QnzdIT/XfVZfetGKl8z/CqyRcCQOjghJODUksCJWV
If0LEfAoDcZ/b9Sapg7I6kXLtQq1HaR7sptVX4E/+uGE1xzfncNGGgI/vbxVpxdF
PyZXwxbCZ6Xxhqnj983CleXQB1T9ALndyThIZBx/gFajmWtse2hfiPk6gULvnCdU
5/c1PnordWJ56OI5kuqzCTNILP49FT2OJM0zcDZ0f+ewnFnwjJ9lC0A9uZFAVrmr
sCf8NQRzrGsZaTgRIxfnOc9+rdtXfjs4t8MRVZvT1xJALoeV5C4B+lqAMxj8wD9W
bwOUuK5NtQRHNF1hkaD2aK2h/Hp0TNVaJAd0d+/WWn0cLgM+8F1ftdhUX9VbGf7/
WXoQ90x+c6qNvL4hKigHxkBa5rAvb+2DDmV5da/ANGk/2jn64/QuCVBsXes3nYeX
x7JC0wHLqJVImC8ThLm5ED3jIIj+lm2Y+Gn4bK11HOUL6h+Imb1bIP91JOMIcRoz
rZewXFYukT/MTWDlVXcvJWQ2O93iDL86cpRUY6EHTqNxB3o0pfMe2sqZqNH1cZz8
LMQkJc74VKnkwAtcadHIDlqoPeuAWWJW+maDprnjdp9vaX9Hxb2AfgFX9pfL5INW
nvEnrvhcbatvta0bR5X0kMcH34d9sGbSoVCkyOpXj/NVSUU6wam7xxXX6WegD2nU
jguU6tpNGSADLKwQFWsunOw3cKerzeMyMV8C3/z4RGz3m+65KujsZnPKV1A5XfX2
r/UvlVqESHK6CLX+5It8gsXHzbb5hZ6MudalMDFMyuhgxdsiHD5K96Rj6s1QHTYs
wyh6eUp6vwjKY3WUQnbHb7nFCVS1WudRRk2AXvt4t0z0OQMQZhi0jE0h9wMQguty
KjMwfd+m4875b7P4CtkFYSttznfpNxoG8Wv572kLw1LqyFhQyefYfODK6e03FZGY
gT0Cb4/4tKvYw5nd7QJldr6FqZ61NI4PfETWX8Srge7UkWkZGZSAU7xEBWbkb2rH
Qf9LUNC5B1p+ZEg4Ho1D42fF1aIGiaCPCJmy5o1yoPzArMCFHOtlM0B9YmRhLXD6
41O5v0AeOpZYgZOfYZJPq4fXqJ3N5PQjloy8pIxbyMjnQ3zUmNz05wimB2n8mEec
Ppo6OUyGB/wFX4SU3LZekCtG4Tpu66D/TBUrmUU+ym/2BiGkcKedlT6t8xtvJmIt
UUTAXNHqpME3QwDflwRF17VTXf3FT8gmasTZ73FqmJK1NT/eJTA7wErHbOjzOqH8
DHKNCTsSg2Pq0mEQBiMH1AZ8wxomBZxoViOXNxeuyx1rI0xduKx98W66+E7nev2e
x0oNoEbFjnBZ5qEvEiTCe5qmb+mMmcW4U0RTdKGYKOqEifjnSjr5g4Oa1ubUMX4T
beEayJu4rfEoDY1vql7m2viijR7PMC81vrIzCf8q9dHHUW5W5oq/hMlJpA4iXPbR
GI3DTbu/tmpC2ubiI6kxKrD2jalEum7NDIj/9tGigB8rddyh/6xlYcLK3wZedGew
cBiLO4c87C+T1mVr0/qgW/6q0fZUL+6fT4I5P2kJ6hHv7+g87EvKpvNGILoagQMJ
XHu8+HGI6LZ4oQTSbm9ki6CRyuDaW7aSer7X/ylFK69HDQO1MBZ1gqfUS4D/Iaor
sW5VFJxhWznM/qFUld6FN6OPoxG1o1jlhMxXQVu+wY5RmfNcIcoqN1FdRSG2qoEH
B91qOB3LD5sW7VXR0CS6fRHRs6rkOtZ0zpILnJqCA6mAtY8Z/K+d4u8VmKVNqrND
lMvR8Ax+8yOfvLjCtjUxzh2z1FGWp5+iInk+T6mnkrinXU4b1s5WUHzrERNVg91s
1eDY0OFvNIa07D4xPraL/0RKaGIEbFME/AILVmXOzAPZ7J1+3GuI4NBQNoEGWcOx
Klg2/ckkiVt+rzimxQAVHUyXEdTZ1tvkoYhQFh/0doJC1rekjh8zdAbUPE6YbTzD
D9k3cV2MWWeJle1Z3sD2YHWsCTa+2+gfbN8Rl6C5MTHyXIiQXNQOy0UuepkP19F/
VGCqv9SxYnDWg4FCy3Nm+h/MQd9RmIaF8fKBFJV0HHojP/zV9Ux7zRdwT3USje5R
s00BEewNkdKQojeyRe16OlyGSTxVaxipW+sL8p5bN2z71GXN67NNFS1xWNPyRZ9e
Ssnl+5Z6On1CNu3Vcr7V/1q0uh5VYV12p3Ia7NNyPAfKPC2Yhp+DjiHQUQx1rIPr
QYbAdNzV3+qCKyRg6X2lPwJfb6QMStL5q+HLvEbrZt6d7/EuNspCafpP1PBFQ44A
wyXXIZ4pe8Z4l4+dQT17AWmN/LTMTKO8c+SqdWVm4KTIPUbKHy4/fBzGQLh/sep9
XHsok7bEQgOXlC25qx0jt658rap8ts/ztc9nloDcAMTAOLVxu8rSmd/WBaBJTcmh
d4+IYD6aPs58U82Wkj1Ms8h9s9xxj8mFH09jVVbl98wS/X3kHbDyp8hx3flAcf8J
xFzZpntCUX2XBmgBfHJrdFNAlzhTZkJpcNhOMgM1b95GA+OBNLr1b69UijuQQi3m
31TxOamtC+54VaM5KnB89DV+PyjSmoIPJzhBzZ+fZIiAjBr6FcIVxW+yxDYThJA2
CrdfMfzukEWQrjGaOf+F5eH3kB3na2V6V7/Mm2h5MbY3yz9AZsLvfIG1Vo8LaNyc
Zn8u1hVGOBvqgMNSnpzDXs2yLb7lprd4Eq1/p3WbkzZIKJrEjo71+4NYrKuXFF4H
zxShLX2y0K9pOufWRz1oCm70rZpw4QXkUGgwcJ1uXUeUDYdMLFF0ZbtXyNS8UiAE
k58S37GxfsiizWSxbTE08eCeFBz1TcR8rt/Qgo3z1vUpWhr9nKyBPsk2bm9B3jtv
q0hLPIu1ATcs8rMXYA6A5/iale8JzY0x5EvN7YsTjw6xh0hP29oElFTmLDEujhCc
RuxF8QoXKWLIoiom9d31eNmq9M3lEFu9Ury2oFwZ39gcqkz9HN/5uebyADCaZojL
3H3e3tCOlHKdgjUu1VCHnynS1MoOfE4ihXpIswmPbox6snnIKDQqZne5Q/vlOBzm
FYJdWoINVae4WFFPYG7lAEsBkyHxydOHI16/9OxD/mLaIWgUCFDprqCzj67rC1VG
8+1bRjtyKE9KnDrgnihoFCyyYDp65phlgOdzVP2FKjtDCMWyPIjPhFNqCNC2EqZE
huMmKI3XymintDklSPkGrOuX/G7baa71o49L236fLmvsfe/ac+N6o+SQlc5Lkrrs
w4U9GQzyYGEWyj+xbQKRomXmvDq91+3oNI+GAX3hY/cQOGljqPNF7wYN2VFOcmcb
8f5PTTL5Z2pRD3TZHLzMKhwjglAwMxpVtrisVST9XyevZ+e4aUqtYitcOhoy7J13
XURu7H1BG6Swp4xswCR3lssrxTV8P7OFTpnfaiI4nnVf3fuA9rg48OQ/q5xdnqrC
PncNTNZsHCsWSZGxFR40j0MOzLNMHRAtOqRP+vJ5WjGZ64/WsJWpRgcyhscSSPQd
EZOqaaI5d9tfBrKBMJ66fBQajL2hXECCzm/adxTNj89yGHS6fyy4Agp0bpeJ14xw
INAbBWJIH3KUl7soo2tqFoiuXIlnTOckuCwqUDmgm94QWl9WHcO81IGw5j160Rc1
6t9sc32SWZ1EjilMip5g5AYIKXUjbI9J9774enF1JPhUEbL0Gt41l9356vFg8N9u
6RvEMsX2wzwE2NJP+MnlFZrx6Zxmxu2zo/y9oXYdhvTo+VJteFpYkyunDJx6UKnH
sos2tnNOMEsepT9Cz9B/9MPS5cSdfaBn80CQ0nHxjAx4PG37o7k/rT0u3b4ec2gI
73sFpUzTpXL5ceGz1ij1d1Q4qf0/lj3wDXs6mkxNlsy8AsECorI65Y5TvbJY0YPp
RibcuGLZTlsUZl0//iHna/qNYqGrLrS0cAPVC6NFLgll2eMoDDLeklda2TVFeTte
o+yXmPfcfGUBjykOrFSNnX2kZdglKM+UnOEse/8NzOQfENPQ4Q5SFFgFcvYXLBdk
T56M22fBLzVmh38SHtVNUXL3GOkWF8oxavs2YmgeWvCq3SyS6vAazJIubdbmHp77
9NzFl4GTYEUTWZZLXi8mKV5Vn+c+82vHpAUq1AFp6zE15STwrmnWYogrF4YwyVuk
vFwEucq2uKc9w684O4D3yu693gceVzuSQ1zTSUDc3jPNZ9lZQRNXXDNeo1ZOnsQs
HDWT0dlGoYWR01JkXhx3wI2ZRG8sxke0UBSsc9OlvrOabmBQ8L+tLLDukXCBhhua
DBYeLl9Ty17UPNZex4P3WK6WXQ/iXM6KiUSXhPE8f1aWoglM0Eq5qCL2mwsjeLJh
AP9cWP2P3kRq7jlnFrYmAvaZiq13bOH4xLR2zR+gGHrSxlUjGNQ9JSHsMZtcu1Ts
/5G6otRqMZtZ8BSTvhswnPcNudM4FEbGkBMQnVzhtmtVPfraHWpEzE9mnWOxt7MF
6BZhDgCLtSM3aag9cqaZ6vAPcuRVlxHM2waGOiBbAO82dJ8XQu1QdPXYcGstWE8l
6apnUW9BRdRNlWaZvOEDufiAqrlk66UabpegD0/rSASz29C20JNHBIJtJvg75EOH
fdTpox6gTQ+rFKp/hIF9dCrRTvsxGWnAcUdSMTqcr3WPBImcNfIZaXzWgpGw4fbc
Y0JEDsWFBcCfph56HqHqKm9Zb90aLQu530DLK8CUGgOxY47gHoG8KC8fajAlB6Zg
MclNNji3pVO+kFc87LRvIWOK7vDdn3JF4+WLQ3/Lvay3uH08MhcIaTwZw0bMzXjd
Ci2dctZui0deq2jn42ZhgS7CpyGheMm/EvBiD+HHKw3Gphum6KTgIujgdxFw63EM
e7gtB7xdv60Kilnr/dfo+sNPjHQxEpugLpNMDFnJCISJqHelbBFyQEki1Ddy88BE
ij1QEUhadWiGVTdmaTp8a1Gy7JfAPbAXEqKIeRG0KBYosUJyYCbaF81bgHkenvNB
XFpBaZQ0nj9Pz/jIJ/OgkPpcnRTU4xgweKkTxtPjcyaiKZdVqmL9fPhMv/jBJBV6
fjFtCOsI1PK64yQZouORufeneifXeGqOQSU/pBwPt9Nc5X6h9b+iHbFq2aXhhtkj
CPffvDHuYUFNbST6hIQipR5sH2yIx7kVoZOkyTEdyUuSkiT140dTE1lIi7i2P5KI
FK6WKeejOxlSwasNOMB8y4a8cxYKHSQ3Pvxmm//9OLZySX1jyR7oirF29TstwbiN
FAnS23QVbjuvg+o/+WQHzCZvd9zriUvNFK4bkIXk1XNCX77T1Z1ITG/wzm/GdGZB
qo7t1BAlScDlL5Q49ljkosysjEaNfG9nkQBp4BDTJXqYpZz3samgOXI8xg7O8Grk
2fZZRpWIsL239y9ajf21bbxj0N+XIuePj98OD5Fs9QJHytI2ABzROEP2GGet3Xrx
R77xeU8cZD/Jbv4kAPZbiMg4byNg9fTqrK4l9lCtbKjsZcq0gJQR5Lc57DPcgIfB
IrYAEQFEsLWV+Zx6fygZ1vRD2BPbQ274zTUO5tV5ENklGyU4xsnsVS401Y7UFQ9W
KuZ770wHUNyqM9Qi5ReedhksAbJTdBlyIsG+2bSiSwHWsvWfd1gTYK00V2QU6BdJ
ZbBNkvVZSFDca+qG1XGrwj2JDrRzpPzFQX1TLL+yKCKPsVPIGOQULOlFoJebAkLk
HYPyNDQ3KKaG1zlrFMdLxrOXFu4h+1K3TmSbC+o6XyIg+9uUVi4cKKVtUeoOxdUZ
5vVnIGaZ9qRuxOwdznfx8Zlo47XOccsToPn8wef2nWKIBB/3otv7T9vM95I6gU4U
X2mT2+iNoZA28SM7irn+dCYPQSiAMxGbr7BUqQU8ufIehztdTlguDqLbXQVgHHOu
LsYqsCIwDBwEekFsrbkGd4SbSkxYWbBeJnotvcurwdtAl+pMtBLoTNL2748DNZpE
ShFBbTUcBA1tYConDXdEuhoYkmuvmfaLnJtvq3KbBWo4/upKA1LwqgRMkbOwc8du
sigKC6W7G4YKbACHU+++sTXPZ3RCEaT6GxC6oJIfP0YrUmbebHx0EmrC1yzCVQs8
Ju/wIUmTT821cmwGQvi3HGvcPpJ3t6pGxZPsK9KnTGFzF2whdlg7q1xa0OWqQq6o
EKAye2u6ZV5dCN9FWKlLZGhLgq1iBiwnPbjIpRuDJ62SNZF9ZEtwVQlXQlKp7tQ4
J+GkSW4DCa1+cBceSxmdrGzdG5uwoMU8g7bMszbxu3du69l9JE5x3is/co/lB038
PmTPcHxuF3bpoMBJ6RW1PWJBTxShEiy+dW3ObIe2AhL2M+9uPvLjZuJe3LinscWG
IzCNx0q7xe7FkgyAI774rCdJFPdPTOm3ZcwxuMM5PGGd52/RVqbA5w1/y+C8CpJt
waYaJGz1xvLZTpfWxP0XqNBjB8wjy+ZEKuF68iiLKhbYs4D1WpmudMCZveaevPVY
Bdq3fjydP5Fh+Sb+4qtu3gXhKyR0yZrBADZGJU5dxcjC7tqIGlBnHliqYzue6a1r
YOAPMcksxOhVrcsBI0/fltDqpfiNmDLoWLXwOSkNWrUzYh9kIt//KPtF8yoZFfun
AUBAwt9qC21+Jvzs1mi0HNN3UJ8AKmlSDJ9Pb91qAwa8y+2JSwSj9o3kxQQWLM+t
yuyeh6ghn0dUGB1LfTsP7Ffhxhf1/wp7szCHM3Z6+Ch516PPRQ604zhZK6VxR7fX
QISjfJ1AtvtAf5mVYjM4UlA3niQNXn03jzWXLbO+PvHX81yf71kzMwI0gS7MxYmu
sti4wYn6m638oFJw8hgg+IMjDxZKpnjSbR0ViOI+apLCwxqsYLKzLMnkogQerf3x
TI2kDY+fInKuRl+Ho1LEX6qyj0dJ71Gj5KgRYaya6VSTbhRQw9m0GdizFA+cA99y
V1GYI+zNZgnay8IBuDJ8/2qwl+Dw5n6ZiJM2VKsIcL0MuzOdXi5ywkqmor+BhIf+
rYL/6/VnHY3BxmWUTsfOX5OKsQ6Y3tuFEkN6K5Hgjnn4u/wbnZzOm5UTeBEnyRQv
1cMgpGFqC2qxqDfiYXxNAEj2dPae5+PyyCd+YTteKn2eexwA9m7I7CjdhvqKEm13
w7vrsD4hLt9g+HGHBVJs3N09QUL7MOHtzTow1EOEoDFcRn0AqbBITSPXhNlITbdH
Bwkj3iiV4zx3zReo0LaZ6aU2bILStoNaYPXRyX71rkOO4ai9KKGjBVX890GX0IAC
sGb1fOKoXoRPs9auBhByaBfQEzhaGheueJD6j3fJwTMCl7R3yvvDCPooBQ3rcO69
SrjnlYm+qxWp0ddQaBBr4OeMNHUuc5l01Yg4Y0xw2RFf+iSR4pgMtPc2nfvzl8xS
DYOnY1/Eq/GRBI6qYQji8X0RYJmh8PkIPoarmrLUY7OLqzCShKtyYakaQLYNeYKO
mBChluK7O1r5ELYL+WZyYfvY9vJV4ARysWQu0H3YXvvcUL//jYxa1EmUHOz1Yubi
SqNPABCE396oON6AnjbZV38YbD1hSeVYSbxC8jtswSsIJWAhUSKUde9Rejxe5/+G
b3PluKAbWAxvEUsPy7rsudDC8MxB2r+aiSPqoMVY2qfkHFTy9g75jgEVnlWnFQ7i
crWx/S5Qz1iprJFsrOofqJR9hUG6FrKKeSNc0nbCjzjysj2uwZ4whRD/O/s0OjJI
imLcgTVwDkkTx+9rvjjjDDn4Ht810DU1PVnFZHZuczTmuSC1axh+aX1i+rgEom0k
0qiqmePKYN2KWwWVnR/p/tHDp7AblYkQ3YnXAcvdG71OArZuCdPi+4jgVAr7Ezen
sun6mAtNGLFj/qWpTsa787Ar4nsZD2+bxFKc0/06WyDqV0P+iM37udEbjD2NrEPl
gw2Co3lUVX+aL63MO59ucOVUn6/AfspES7A8LC8t8pGA/2aR8ZYrS4BR98tscms6
JKss2iSDAGfZeEy38e9zy3SHUd0i0yPnGmo34cmKwOxWXlA+LTDlWIgk3ro3EtRO
tgK2BzFt3ZyeTwNN0hcv/5UA6d0wXH5KRIfUryt6JFNxRRiCj8GSCeF5BwBUX2/j
ljpuvbbyg3MkmjwvEuhDctBc8WAJqigr8KdSpiQdnVJtJTFaX0UehQ6paY3uw8bj
kZOolMtAy4Cyjshwy7bCrl4/cCqeKB/0PWbm2XttmhI5hjRMSNYWX2FE9s7mpsGM
qSa9mCKaI/NZkoiL9PXDUDcYJ+i8Wy3dhSaKgV1Y+pWiIstETU4HnFGgXAa9lrQm
RfhX8OCaysI0K8jDU0JIGLyOkmO/6fYUVesruS/ez3jiMEnMRjWhd37k2/EX4/vQ
UsJhhwbt6iRkF/GX8NVI6dvqlx48tm8iwYtHPEzESI60TKhbw/6F0PMPCup4gtyM
afjrQK1QMB12cYtc3VprzsdLP203Tj9/EPBuLlVHLuP8c+veoOtOUy/jUScOUllx
eo9UCL7e3qhxTdmSObnAraumWAX6LXeVyFM6EEcR4N8S+49zTI+h7Bcm8joNld9O
GzDKuFkpvrrzVnbg5dojDJciljsfDDfB7c53WoAnm8CpoFs7Ju0LjpbN1RQeeba1
2jeoNhox1pf2l0Re1djs3Z39goaNwkKsj+q2sMkmzN2hJ0U5kG8s361df4sEwYO4
EaXO2FyhPNtPCWkhSA1m5u6XzVMPOJwFss/Gi2XKAhEIasfR/J6dItFoyriWnYPs
DSxjuByeXerpJeaWMi3B+MkjeRcV/smOxcN9pla2x5ySaN4B2nposl/FD8ypbplJ
oJfvPJ+nqyh9OK1fMoL7Yw95iTB/rtdijKub1OhiYHpbpP1CM9tIt8QoU1HE7yDu
EPbQz3t3EhGUhSUAsclT11EPwx8DB/COfa2fRMu9BaYJ8jGWvvykr/QE236A3bCV
ZI1dN1ul10u9sOy7yDYNsdGxcLoRJJa8ouomlulTXO2JKzwtBZAR9FwAPwuor44o
2IX0qR0ygg/e2MvcNuCk5DS4qPKMGP18q/hkYpIAxG8TYlffd8b5krZX0Hi8/rDr
uydLu7FF+HnaYPKwtEFZIrbsjJUGAbYQCjTqwjEJsO9/h7ldjvPPsEnUpiIaz1a6
N84/vnYy3ohUlZ4Et6RjT86MxznrcvCqT4Is8EnpfB3K+/EFtovxAlcGPmUlAEMP
O4aU2XzGeIXZlfcW+m2ayHUFimQsWrTzJAka7AisQpEk+ifClFzW6GCD68TGLXxm
u9yKLsP3WuUzTdzR+NR2T9fOSKNMQorH0hyfjMmhxHl23x554Bbd3VUPfOhyFVVK
NY3Twv2fBPhJXVP9e5R9jf6ERc16O0WM5jQ5WG2r+CC0Z5IN1d6Glu/29HF9paoI
zi68OHV7lQ0if7jIJjdiZ0nkGl2HGUd/ZPWvabgwCzGunJNv00sOvzcvSluO2Mfm
wJdoitvqbQg4wr/Uli3JAdGc4fH5QmRxMlWrMsrV8eTILLEu+I0eiPflo3upsTKm
LViOYijvHvu42TXTaV4b6PKtaYKYUCKjS2ilRn7FfRCqxUv2eFwdp9Y7sz4NwGZ8
2C7ZwCvBVdRl6S4hJOqdHUlRRovpgZt24FWDKt3+OWVEYv1dWi2kNNsIbF8/6H/S
sIsnqSNAb8vQ9qEDlSeB268C0sPrWj3QmiqypOO4nt/iHnUhFEC8Wj9gsh1OxPfg
cihpobCWccOo/vfvuOeFJ+dW6yCgUnyufkDY11VnBgrnxQohuOcSHLZW47lDh2h8
5BiH7YRChWf97gzHYFVM3flanQWkobqAF4L8z+rcafSDv91C8qxPwNR/hIx0uFPO
LC1Pzxn3bsOeRPRg2WnwMPpS3mkxHdso8wXp3vQ1eqO7TKb5aJU9lvAwCDat8KjA
vsHDnBuGwefntedW+QbgfdjriDbTvzQmJnxNpHLjA/R5mMHjRPjyYe5d0OqQB1Tb
4wCYj7nshRLk3zLoPycIAyz5jA+8GrxmR/tDOjAbL3fJCoW+OjnymRckJI6t5NNl
FAaBYq4aGCJhbvwUmd9uiCj/x4p+9e6wz0m3qaQP1zPfIO0PMbgpImNnjasmpcOf
9cvgiTT04R/qjgGq4KmJ8P8xim4sDEXTB4KQmBVdBCtEKDfLn/3A98C7FIcQHAt6
fEeHTkD2hAbx02CA9NsMypamCuQSVC0pl900KelaXrb8WKSVqRSjmRa3EbXwAj16
fkAGp/msRfv2ontlbInuDw2/HYU1uLgjx9OH525q1peyFLsOeLloT+pq++iPSd02
9+KOM7ndtFTgD2tQ3SYyYVD1x90/a6c0LHJeqXkjOJDwHbFXf1hJwSMwhC2dXdGP
uHKcOZ+FNBWzm0H8xfPHqI3zOCoD5f/AdggyIm+tR6DruHF64XcEqPNC8P5/wxGD
ilaLyXJFbD+E8mngx9D3Cu9vOixQ3hiJabrB/qUPbcaZhMesp+iQWGk32UJWiHTT
ACY3hJMb2h1mX7yA5/td5XfZnCJDGW0BxRgfuXwzTnHlGfCZHFKZwm6UxXZAjCgm
rJ5rLpcmoPXOaMo2S5A1ueu/2sOnuf5R4NCAqqCJVmaP0H34MEHz3nqr+c5QoKGi
mYT/izWrojVDDIdZI/tO+O6/0mWQCh+N8YxOmGqWS+WljoNs/wu0pe2ZhpGdDwf7
1Ws6H/OxZjPWgHWJc0Ct+G70LFg79u6vf0TMwRrhBZYnF+gZwFFn7Q66Kozcb98C
TfV0W6h2V2HsC+Evj0ygAkvRphUU+PdrREiJG2oJ5VQCTN/NKa1lcMSNYDKirWFY
UWhK7/M2439CFN4gYNBM7hlIQxwbE1tIOcwFBChCVFiJZhT5XXb/NU80+tu2kn0+
OQhS7X0WGXJCbNMGrhBRmoU/ymFV+tnl7Bm/X3yZDB7JgigZ4Vt31gJYJoEsxqIU
mjWe3Uf0ip7WTeseWP2nkcOg48iZleVXVMvYkl3rTav26ttV0atAE/kyXCxiWE/c
LRZ9JnrlTJ17yS2deE0qTAFA+YKjA1VYCAoAIOO/uG/u+XXcfp1LDYzM1AM1rCX4
jV/gTXOWuZBeqaWGlUGKR0xh44MaiWZRxUvYoZHr/HOoTYF98gP0xKLpxryod2mD
bKPUICdVE31QtKXDGN8bqwAAq4J1WKFlZ5w51Ojj7S/700W6wilt3TsJV0Awhjwd
tHlnZoUbX3EH6qDq4E65nuFWkwZ91RA4DUgJ4ymCv4+672EWzU++3oBYYZXERKu7
18A4+30XaesSD67NlJSqqimXkrfJYwd/RNuXmCdo3ia6FVOBlMqDZhSdTZDDyDqU
P46Ws/eVeifYIY/Yy6APOLUfE0vBEIpaSb8hemmsQvWAVTEV/mvS9MIQvtzmcrT8
+w4Yv7YoTgnDUkz8KXjbpwWqPmJssq3nqruotib4ijnss9eh9xc/htH0P/2eUED0
wYC+A46iFaQ4yxOr7VJ8XGpQ0bs29+f1zHyTVsbTR3P1abHIqH8vyENqN49CrRzX
YFF+vl4CfzKHJWyuwoojkL8PHMElASJMro9BJWROk4eebp1zrUWsYL2bNpDI49Np
PwvpM8wlNEaf1iZOeiZaFkXBUmaCR1pa2+y7Y8okOYvjURrOd29ByqIzRzismsGg
7Iq13LHxqLbpwnnCsaqtPrALgL52gkrJbLhuKAItlPPxUA3HIfn2QVuEzujEODrF
Z9L+9k6nVVzif9gZw1IwQnXUmQRitfLi4683NFQstzjMQMRKL3QnsUxGvjT24J6a
FTHA+UCWbPVVcIFjn+jN8lN4TJ0UVXWW+dsqMWAXhrFAXpwWAqYdaOPuRDvIPnuD
xuSISA/Mf8ZE0O4dAW05D18n/K24CNKUzu1krWAChnhWGBjVIpM7+W3BRjEe4X6a
FF53KIS5pGS2pKOsN2sSCdRGtXdlsQ+QV/QhSI1HyUk3av4dFGHJzRHHJYixPUZo
Joi2/XedJi4eOJzwQhSCeNl+f3w0fHX8iijIn5SCezowKtsDBb/24hO8doX21iC+
uMinMlQtU+5Wlk/YLWdDPEq8VYerlT+vZrZH8JclkBniKdRKte/loBfxqvxBTuZF
k46hxR0srl3HUdvdF7Hrc21wkbCQcae0Y+VrCvfRPkE5MU/euCfbBMiZGD33tDfx
0dQgsjFEWO2lu1Ecrn4XswqWS0IhrEMcCquwp/xa1SB8SUtwSwjnD5eHuLncclD5
OfJSomqyorFw7Y28GiVkXP8yU8vUCFiWehgSPr6O+Qk+8JKmB+JobfFyz+dAHMHm
ahfErIWEkkiyzKtsXQ9mB5iJCtvofnyuiKfRPtsWegwR9kHYTCvIgLgYaunIMcwk
w+hgdJzLNWZ1oZVsvzJt55qnrarFPh2KAP6zQkM4hVREtkCowuJuDjGKP2ifcQWU
emIKLYcHwi+o4PZaiIEju/QZm1hl5d0DJS2iO0rJLJgqPQOs5tMd6GLX/mT3pWuZ
+dIEzVhPH531mjDq9bzPBNCZNaEUw4OjIxTozww1zgy+Dxn4UXmoYcTEQI7oQeXX
zDMGQSzQ3aqp43Q9v5yswnksE6WQR/FQCaSN/WNx6GAp+mVTEoiNZCgW8YwYj0Em
72B1pBOi8CIj4M7fxQf4l5Ybf12TiJHJOnyEAfob+LL4tvIhip5UW0DczZkMZ9t+
hzTJcpredkSbihknEImbTBQjA7+tbcw1afxV9Xqnr8eQn96RAgSrxK0kbX7Pg3+U
01RSaVCwKvx4CgSk3jj8nxtCZB9J26UfLJ5PdgH1GCI585OAkgyMBgdLtXoauKww
rFm2nVTTAKnGUCEB5IpH+pjAZpgNGbhxxQRcw1ULsgj10lz1rtQxs3GSP7iW7mnr
vtKs7k7bM0InkPGXveKp0zBKZwjOLV53Za+3vcvzK/zQ4WFn0Uhg+T3qn8O1Cy54
qAnVoFQYl0iH/poUDt/SOYbDPZ5kQg2bRsAr/n/oH3GjBZv60BXG9VOpT1sTEwIb
f40h5Pml9j773NQcTBaCBH4c96BmyfZVNObU2PxmZQwgfjTYfOPCgU4jeQmlfEdq
wKC/RIQTFVlHqSW/VKptcBtvGOdagcjvX5GtecbMItD3vuBk1SikYA9/tcJvQuGa
/zoQ2B7gn72yUdm7JH60h8jymNnRppv81XIfM/GaAFxDvLZPI2VWySxX9ZYgXZza
93JtdZV5xcxJPen+ep0Wd+nmJR7Y/yhXH5E5tGfZCXwu+7jCGSpxISCWlBAndE/K
5866SL29bwGssPUUdyIzVNfxwoCmqkyMbLRNsX7c1MTzpuTFk6s9Cj1GsmhX2fMy
EYS+JuqIBiPKIJuH4/Vm7hHGvbzY1MTmtRXs2u655mQudNIzVZ+MYDdungARjG12
ln7EOUyVTA71Kcisdc5gHhrsAOGjpSMuyoj/jeDqoeu4/djtZcdpCFlvkZ1RhlqS
P6Z4B4Mt8MZ37TwDqOizI/MFwowY4JB7KpuqqEVSpamp5v65bMvMpslOx7JA4sJp
FQzVxmJBQnIS8OLE1l28b7lqzQitSWfhUDHKV/9lUrVahwQOzrX+LjSMC8G0VmHn
YxCc4o0Ph9vxkF2rlazgBF7NQN2WSXcwz80s/4gXY+Dj42dssiyCoQRit3IMvor9
p8Mu3rCIV+Dy5aQD/FaRXAh5ybPkxfbeOumfBPGWPLl6cKhKBH9cA1sFss6wL9HG
2NytjuyeBLw8jzJtTpgX5uYY7NiqIy2AsLO/PWNf53xANk4hgeVFhv/yRC6lHPf8
ptLd+R2rIxRXgy27KePUIEZEI4eUZSucFtU9lIxbSuxb+RoEL5wsbC0WJWhId01T
SAASjuXqt9i+OC+R/QDhWs9LG24evpJOsBPiaQcUP1h75SKV6iUlGpFOZxkxq4oD
Rm9Jjgs8yKM41UnMapTJBFxVfuaeHNjlQ8whg702WepwZhIfyfW0sgi64KTUve6c
dngf/AOeyts6YA2Y0oylQz+qjDMOqG8n03T2jEUZXOudz9mwR2bHqmHBatnb3Hid
c6MuoP7LIyrS/8bi4P1ZzsTPNmCIYz7e+iz3qzoIF89yE3h1IJZ3j5jEDA+A0aoX
lNYcWdY6JfXADFOE6jodfXCkmTtKIAclw5vJkdLjXpviDP53qrhaKRWHsyjrM9n0
EVTg4d990KRQ2+BPJp7dZNgEiHk4wuqeDV5iakNUe6CczrfRFuqoQk9IsJG0EW6A
nLUwQjCG+6JcVJE+rgOmQaKSrc9W3fQw2STza7JXndZ0PL4dIFFDPwxEtPMtpZNV
7X1c1JbKbw7QYbDa9lDJ31DsepHsOBp0NLScs4Ma9hzky2pz42PfUFctjEIm99Le
U9HexLgqv7/3x0H3p2xYzJfdZ2IxLzN/xxZUb3lmfABJOAoes0GWs++kgTH0YgiD
W82hBRNy5XHAvSSlT/7fZrrSg+lvIUnc6AVLK3v1szmt0+/gGDM4UHhWWKwPbFtB
t8WqALS6sMsUsfm48c5v4Z8XrV/FdkSt/i06UMTroeKPsLHHS3Q5M57jzK6ps84o
r4W7EZ2ldEHyiWcpTzUgycLrvTFntsVDxlzG8Xmbwf4Rj+S7G3RPWXWGWsck6Hbf
TWSEmkgSVzcQ3Z6S1vZw8LnCiHwca8AW5W63kspY4HblGCIE/SWwuwgyU1sXiQwB
e7MppObEizIbzD7mSbDFSZC5eh2kifGCJSy+sVqI21qhniT9SZihvpsRo+nVH3jl
DV7XDQAsZU3pS3jYCostiwlG1a3GPeHDoVA3xVLo47DOFXStWaidCCbREwLvoF7a
79u/1ltoqIPxyDio3vmIFQne3CLtqiB8GlrCvbxnGcGmYHztRRWaOB11f83is5ax
3SkhviLeZojP3turFHdoAl9AEu5P4qxmX11zfcWpcONiAF7TQ0fLa66KFtf60U5N
4pyQL76mbpEo3W5ATmv6Nz/IpIAP52Ki1p6SY9QVoYUZots7Nq6dI99QqPd//n2k
bEj8wsZqzipiOL54o9MHTpIe1zkzSaD/p47VtWtfSQLiKTRx+y4R9cOoWM8ENGIM
6l+1YPuuyR4yJNgcFN3UtkjB7aa1OKKw4WDU83rDXnP8QQOZzqShehkriDAliz2T
N9/ufhF0csJxLNU4bEmvNO3qEl6Hk4sLW2lJvcBE/vdHoTsWth4Gp4CEovZkjdWG
hPH7vyhHJpv6a0TQN6bOUvVROuA/EQOWeciNGoBeK1LeMIWOOXj5I7WOFTZG/UMh
VWxcNJvYlM1zURe5Mbl4lq6r6IC9lBkj8Z1JjxCdJlY8GlleMz+Pphp7a+JmuDuV
5cDFKf1RKpk5L3DKhxVK8H4eSaagsEGCQ3bmqs8hovJWhej4Unag2t0QmuiMc57E
usSJsgqfMUvyiS9uGrTwNhlcS0RGsscH/zt0f2AeaPuMzqj+mJ9//dGPkPEYRFqX
UkAzp7ANrtcnL98M1vunDrEKrMkSVp2cAqLdhpsQTSsiMmgZG82aSgZ8mHOd5NXV
X+v7QX9/u1IUrZaR8BLabN05EDIGgfSLiVCnSryvQ6ZyhWEkOWJeLh9sKvhEq342
dsecn1ENWMEupBrEIoFyq/xl739uN57vBwNnFgjbzu1tszk3B0S84zTvXT6TIW8z
c2VWGDWdeon5RWTcdgCYYdQZ95CZJmwefXgyYDHj8kol2EIx5h/KAa1Hveuq5a5x
RBFs/3l7tULkzCpW/dsM2ma1/qhtU/LdX4ni2UDC/EHNBYoDTJYiSeR5hyhBiUz1
H0IYGKvGxtMEc8RY9covwyDh9mYftilDbQBL0vGrbH4defrkFtgUK1qRQLT0vJ00
K1LbQ81IcryR8f8ljSIsZ+SGt7/ICTnbd83mgNLcZEWdcfA1Xa8qIix+EX2TOiU/
HjeaRQMVbMCOl3wTho/pUbzOHvv5k6q9Z/oZEydtYnFOt078DCsh9KtmGW6tiDLY
gjrWC6/QjdyGL0az3Jt8DoIxZ6KaRy1LTzv5bgTtBYRBfpiNlHDISnG+srWrdB6s
epPmorR8er0/ZGw7e50MV5gw0kxlAjwtj4RhqPqSXO0ZQW/ebrTklM6q3IUb8Cj6
ViWOiBQ8T5n9n9614gxWBAgJKjajdMPK2cRke70cTycjf/FPxySqHSuElDLKl4fu
UX9DurQRjQqA2nuqCcnJ6h+Qb7XqGGKm4GuQapx7ENiTUY+WVmn11LrDAqaFsQPl
4+nQg38zhTYqirYBJozSE5FP/2jg6pvRDWdORyl+cbR08p6yBEN3kPD8V704RZfX
6pJTlzd5SizZ3JP2MqPsihka4OORo2qRHQEEy6zzxVKyL0wkmGWj8P7mD1eFWVYC
Um0gD+hB8vlp2gpAsUlGUv/wkeUUAGZRThpuLnsZbNvV/nwdScJaTj9G0S1pmzCK
NVu4L7Oqjm3F9tgY4tIj20MaRVEoEYT04b4l5PfwU+9xwEr0bonJtoHE3SqZA+VG
JTcCrpKPHG6Q0TctfVi3JpkiMFuRqKB+yJ4c2gXpHmpZ2ig6XPxTelc59T2bqZxP
EUX2siA1VPw1oZMLQu72smasIM8aM03jUs85gTwHK79+jltEOcEgtYRTYdLInA4q
tbwn8d39942d1B4hlFxd8lcGMyx73OvbDv6dRFJDat+IZK29aDLcSmfZufjLRvZV
YqfVozbscvEvYomAGV7bP7S0RmNrOfHxEl4Ey+bCzvcEiGr7qR9RGoRCNQZp2//W
qZDpfq5mqldBaTaHdIpZ6Bs7bIAI00QNIGRj9TQDMPR9JoLF6hGo5gYUCSrva8dD
GkFQGlIki2Ru1R3HAbYy7NlcunqW6qa5uLheBT8/UUzvHHYWpGns09g/aqWHTCtS
/QiIiPNuDrQHeRmpnbN2EbDXvbPn+umCyqe9RjReAu14TqOaCUlpTftZe0AOzZey
3xPTqhKlRXAnLZpd4B0+B98PniFASKZOtyWjm2Oe99ATG7X73y7jnAvHxMLF1U+3
rb/kGJMoFRB0VpOIvnkNu4eswQNtUEtXNKPUCLKHscS3urC2Dm2KoE5jN4XYWzpu
Jt5oEWX9DgRs6uqtFksvmu840z98HyVzsXRzdfIDvSBH3Q67REZu2oYuha7pfE/S
A5teXWH21ACGqD0AORqFv13zK22Camx02IY0ZmuBoNyN8qqa/aFpSIdBLmlLqpjI
n+cR9lQAQdKWhuRglMLVs8M1l/NW2jPQNwGlsugARoXwQxBlnvNNSlMriQjXR1En
2jSQJS7deM2SmXhPfZXuH0wLQLketuFZha6oUQAbFsY5EIOFA0YU7ZMATN0J5pHe
Q9bb8Gta0woicPazaQvmzCCAdMlXpQxi/COjb6IgayjvRHoehCYW89fangA/FRrf
mtofJGiazC1vsevwkXprY1MWIXIMgH8lORqZnpydb2WLDQKJJKtUAuKO94It6M6R
OosvFPzNFBJ5zRNkK88YMeM9NuS7H+BxqbZQWVfdFJlo/PVbUg4k+Wro26907UVI
AcWU6AGk7MHNxAKOLHAIAgJbhVyvDWrWWiV1eAEKVt9wxXBvtfoUliHRE102wUjs
JCLLjL4a2l4O/S1V5u9Avd37ydSwnIlEkt7zX1qdywPvu/tZFM6hFIiuaNKL1dxp
CVaaePkcXY9+9zP4YDUm8RvPlE+9a0IlF7Qr2LaIuP/MnqP+KS2VPYRFf2HdFut0
bqAgD5UqBhwBQOwS/BkZ63WCedd9SjH9KrFm9wSOD99KMVG+wLgDq1CiF4FYz4Fg
IEUGalk5FcTv8pwL0kNzksEhtL9rYTdC5VK8z+75v7+95Q8zlLe6DKZzgPhhmgTf
WdN7Fj5eDVvzvQnbh8zzkGmY/aqMpmpIC5nJodFymCeL170efSbKZZrdBHF8dgxD
eFLuIKeTiMURgOY2Yhnk5ThTL+jx76f2i9gjemgTpJu2FeQyLuqYPJAhFnO8RRNF
aErd4JNtRXystRGZWKHYyLaUGNdOXqBwV07wWh15tUr7okheLkufVuNBSUs9Hkrp
/+rBlB7kn5q84YYrGfCjvtg6B1a+d4YPumE+1lJfUQn44TZY3VV3W/kOUUVMrSeV
6wIzqTVS7YlhAyVjDzKZLvmsToyld9U5gEO2ZolpECP/yxXKnDC10JzUBnvVPQML
Kv9XztZBLDIregXJVPXixyTYQUYj8x5TsfR5Aq7qvn8otIHTl8jWd5bsXLCXk+oX
SpDpbtmQcx3UxP2MOQr29Rm6uZnFkXdg4bRyem6tTSPiV5qdpHrsCb2Pl9dtGCQA
K/wYEGhIK4P4L/DY+lf7CWO/5SYRR8RevXM29WZVo+YTSgoaczbNaUmTMc50TR+I
DXKYwrliBLQdl2kstaUyJtsDrQ3w7640N9Ta3+6+alOwxGPUSvKRKSSRnjD9jCPL
0TSe6VfRw8H6YYs4eRLzyimnNFtYgMBq16IzOVBp6lbr9MtXk5vz6KXZUjnMHYEJ
3hITQl8BWRYouCrOgb6s9wNsw9MSqKQLwTi+9D830oRlgKEwt5foSAxWY8GFx4Cl
mZ5Tj33vds8fbl5q8LqiCbQClkXCQy9C5E9bA+Ss2yCGx15ANCpQSatQk8zFxX5g
IfJ7kGsRjycge8hKsYFOGyJfKMmktuxNNRknz8p9kLovycESgIHVNJtQfAxQxfxr
Q7jvUBN1mY8yHXxir34tJ7AcNg8L5CXnMFV1BgU266MW9Niqidu+VxcFnPpDr/rO
CXQ4jcXwlpFhAsQlpax7kAEfMDvfsA7l4dRh4d+w6iit9PZmnB1MauPC/faQ/sjg
qci6b+it0JKEd8Ouz9o1ug2LT/mxgyLTzDgGeYLlHmWIFoF2dwCh0Saiby7D8mQs
OnUgP9IYYM8iN26uAxpe9jg4lozKZ/LLuo8lnGrdrH64DCSYJMBlL+xOWtQLwJ2c
ks5WIvfO9JNANvkEFcmuTKVgCljObbERTi3GzgYw6exeHyo/rpt+qHfhRlZPeliv
X07fOKwxtSrZXqo5z2hLszjszgXewwz4d8tWDvi/7K6VpNKCqfbmodLZEwc2fkiS
S2qMi49jxffSvtQvKhkb+pUu1cuytCrwdE6g7Zlg0uHRsyX4IaqizB63Axz92ybB
xa41/BtIOLSHS6mD9ytImyrvS8OLJe/az9HTl2TNoZRrB/3+S7OPb4CJhL49oYiV
r9q39PpsExOHMPJsaRxlkVCEN3sSRaaxjwrBm2NwmG0avC43dCf5IC02rP0gZ1tI
eRJFochWfnUAHB2eMAHGVWJLCu0nHwoFxiRIk4J/lmuGfSPFd9p/zjWv4sLwPm6n
ZBQ4BXPAiHsNrD+se9gHJgTgOR29eiOe2CUqzsQu9EmQtJW5ZgOyqPXsncgwzlpp
ky7cgU17ofFS7kiXcubs7k15CGJnLwA1AhtmXpjGQwd1FKuMf6S010gNDIXIhQY5
eriHRXXjWfMQznOsoZQmHeLdoD/9oO/YaBNQB4HBWoCM0UY0IwpTLgTJrvDk1bs2
5xBtrMcnFTVnds9VtixLxYA8xtIAGxXjcwulY6gQcIVo8J+PYuVnTPn7KD4E5M/H
Kf/LgAdS771Z07lRaRWQ36+y727gqspquT4e9QV9IbBz0HIgyRSFXjbx9Kk2cCfK
08cUFCFIxFF6VgUbfw5ZEfl/QINjxkOgPXpcotdtOBG3q+HVgA0c1YzWUK7zejf/
KlmB39VBMlljYMcRG3mbXv1s4n4mNx/QZBCsYZOuDRsfPFguFA6u016h+/bXxmGA
3ArcsuMehnWAu7epytJ3U/lO2SRI0V6jzWuHPCijuc0kIHYxVrOYZvMMO65HDXAV
iLDMtCeMNG4deAfPEmJ9BNgJnumfz4oe+vRF5UYgRkxezjrhtZ/OF2ES9/8YuHn5
BOVFjIDj2UywhfMoKths+7OKV3m+TivPiu+EowgpQoAIGhJ2aWPBNeECb1x4xtoT
+gK2A7hJTg9bzt26ZF45Hilffj/I035bSY0/tm9YUP0lzCCebuUCrK4uo1K2yv8V
jp1NV7qRVObz6AaUn7D1d2qPexsJP4wT1c+UpvH0s9nPG8zcpW3R+/sux850Rg+s
nV+niVhNpCWxyKNI+fZbWZHb4k1qk7odgtOV2tVBdt6cY0LigZNn9QxJo//kqMvI
7ChVY1Q6gpqkMRoIC/ZqXfDu1v1nS8/E9cJtb+k7k6uQRLRTk4z6N31tpr231mgF
/bQsotuICcmLPcrN0IRLDAH2lvMVbKsdUbU5WOSEjEmMgPvknpMGyBI1BO9JAUlb
KzRAMJaXrUteMBZGRxVhqIXUba/iN+TrZPTjPgVof2AbcX6jBHCZF19kO9E2afPN
gcrFhCZFX65lTjFRCW3qgCZ+7gtmOCK1c1lLrSGItphdY3Krg6r58FZ6NeFM+0zi
mHXDecWOTBHYk74ipr8nSKHf3noF0oWYGKHM02ijGzNU5B9/9n6k99gbeMmFKaCP
buR6XM3NncT+4Fqkg6aes4WrQ3nFieP96fWq3T56RWOTt+vf0kU9XVY7dVx62lVv
stkmML8OM+JbEqJ2SHtfSKO85oBpBM3Y+evljTesbnKISGjcE/nhBC0cyBg/MM5c
HgXXkVfb59eO75HPaNZzjKI2adFIlA1n1cXF8ZCS4fh6fHD5UDZkq66UIThsG2k1
wOKhXEbhSHXxATS1UYEoU5xzWHqSL66aZKDUZLamrQ/Fxxs21ntl6UBtq9MQDkha
o3WY+aF2D/lrZX8WE5Nictwy0fPJlCioWU950OuYM8L+NRnsXfoVb382I2Xx19sV
5mT+dgeOMe7ahiRetxPFUEJtsJvW7uF63m9Hc34Q7lqY8xsR783lzgHwVhbwRN9t
S3wgB5btGumnxb+CFJRUNhs5vCadn3nM0R2OeQhNIhxS0CnUAWwFieYMa0XW5HnF
uIDAlP1s5E1VbkIbqS2nKvL4T7iPkiq+uCbcoky0ymH0i7Ere0L1n5mCVCgNef1U
iiQsTKYSboJa8S3jB1KlFiW6Vw2FmR/hF5m7aojBSJUf6PNPVQo5k5ulbiD+zu3y
KzlpvhezB8tiLFUPM48/WraxpjOvvMDwceY8CDfIJdL/oFdFdBdIYRQFtqXUrwE1
vIJn5CblG/xbnxFJaOgUtYM0DedOgIolkgwD7dSx0WGXrrr0u2SRew9qtqiJn5C9
sqhiT8iqwAeLZG2CAS1e6UVyMxgQ8wKjIsUMtulgL6e7zJtDQK3mAQ/XtJNYiFdS
l514GFGTqdanbaWDt//rBg9RApAkyS+XRD2b+nbcRAKFPAJe/goSt0HuTIeQeKlG
cvOheM5cy5Mxf3kfnqNFZ88r3dERxEilPX0fKECkkplCrnzXMpF6qhyuMGxOC8px
Ykeax5MzT7RlvROOHv7im0Q5AoOfx2jC8UMX0hTo8CKkYxgexlgwnHQOmB8PUbDj
3GoOzAO6Upo5e4GzxhgnsYNVjaz1unmDyZA4H/6Osm/KE05Le2i5/YXt0cEe9OXi
U/vEPaS/o+9za6xG2CJuu///Jlv8lsGlIPNv0YiBzBP4mUmw672XB30dbzCF7R/Q
x5MmMwRNTeETTpdASO+7kJx1nfX95IqZgg8Rq3+x3K5DrY/rl3JblKQM8pLHK1CJ
qRSyS0VhUeXCfDCMckLixZTnSj/WTIjuE6F8w56aNVnPlsrbRZEVgGD/LueLAIFx
jzESOKC6zgkQxtaafbY5nbAedbHr6r+xzxnkAUb4Np5qgRNH+XxjX/z7IQzHTgDl
/cBzZftmwyL45RKmKtWc3+9D4Rtq982ziyszdDCjfwdLDYPaFZF5Gjt6E2+UiCet
v1uUgPJhDt3MK9I5kYRoL1XSf4pWCpTa5I6jAYMVSxn7pcrdpK/joJ10AWSLqoAi
ifhAOMtOzO2EI0I3XmHJSIqKGE0duUdjxt72JpI6+V1sttkKrXrsxdPGfpZsRjYC
Vh+Tgkb/fgnpYs6egNaSUC0Kll1SIZ3jK81ezvkSdPmGTUrVKhCEBQevgqJvnpt/
dTfeIAxD6DlVoYbvg7efHC7Gp8sMzTzKXYFCZNMKvSYwwNxNbpqMXPfdhsyDZ2OG
+NOJ5cc9lAB8VuZcuuhBkD7T6GGGW7BVvJ2JZ02QFztvFE8LiqB5Pw0Xqq5jCRQf
7JQJWYUt9eatofiAUzbFLDHP0PU68qr6y/gAPXo+Fa0AXbzF+qy2ruVyYsiSHDWC
mgomLGoohxkiY2WaZPSsT/DRERUnV4w9bYLhRnqwKkyuNG2vKQRo4Vjur04Ut4Jx
VKI7fI9RyUcaqi+wwEW+j2fBwqqxXAw7fX2HBFJnJOgLSFfTIOnhYPfesYKo5SK4
UiGt951jkM44ynhDwS16yO2+z0LDkDKDKv24sNZmM/g3Kjt2GcvpVfnx9sM/q+pW
N29rPo5hMDWFbQY69k7eSaUHL/VqW7TxWjGts97DAtshYnBhntDyDqQbJTDV7hHV
i1B7xqm/cvyXnhiCv3LO3sLU+7Wh49TZMZhc1CaKB3Yq78Lj7p46oEloiiSTj2Lu
+uM3AI1O0+roMJogptKECdpodNYtPgVgoYrSfsXnRUoKLJxLbRhcnXwGEry5FdGq
BSvGv/R+Lp0ZVN1msm/Ips6I+wtBZkfSgXF00xdYRijkWJXY3/UNT4zH+aePK4SI
ilwoVXXgAX9bo0ijL0bNmr3yULUPJMbjcDQCsRyoxYl5j+4RTsdKhMbREojKLCrW
rLhsRzeuotgdewLysO4LiuawDutSN1Sh50lg2vjbiFXuuoQ5+V/1RcHihBRtdwZK
LygjU9N5sWrgHNssPS0XG5dBl0Gy3sHL2k4661RqczZpb8Ak8k3a6vQu70yECarJ
HfTLtq/PWskYYd416B95IE65gcN+uyt1VQCSWo+5vACa6Hdj71NZB6MHHv3yXg1i
67WcmC9I8qncDo2D7DfrBCZfWQk+rNWjgRYl4ppGOcja4/ZgE9SCLXGEJJTUntVS
QcHrrhDRNXN8Ru2fqQ2rdE57HMlPWWY0lzF+cefUZHWqLeO7Q8Wa6W6v0rBNhoKT
9pHKtHAZVUTK55zb7oyq0j79yACIXJLIWlhRuJ8/pBW9yjlpts2kcBl8poZmET2J
hTUMcHIVsyr/fc4ssHK0nrrri9iw/cM52LMdq6El1XRhBh24cqd2hkHwwLQ9QmA4
7+67DmrfdyUJQxce0rv1azHot262RwSnNcW1UZUPmCsahzyM7EXljLe+6aMhNZlu
adi96MLVA5j9RAqv4DjT8iOyi0ZdxZWw8IhhcB7gtj/i/Tz3zRSHucO5MhuviX9H
VCVnBRhtGcPaxAM8XAngLzQK0oBxlzdiGYCioVju84oye3W8BUkjvUMYr92hYlRh
aY4jU01S/TNvyU/N7sQMN+5TyvTNNi8AZ+gWRLUMXQoYTRjn38EjLqaTjhQUM60+
+Xj6vsSVyHrBFl5Vf4OAG6NjlQoAjCa/m69YMFHhVjG76Pwz566qvcJkigSCJ3aK
ZhcdtUPp9ML88N0C7/3YoqVNsJDQDZA2LIfcWfe5mETK3/pigntNlbOsrBywQhpH
VLOagFRpIED7D7aRRv/Rr8ce8lakIQcrYrqyZbmA1A25VdiIJTwX1OKGv4wfowcd
vTfdMW1enekMNPQaxVTtRfwSuFNIEfZqxL2ITxNdfso9W7usE1D43GDH3s+eKzKd
qKDpy/er++96ofB3KNTPQf0ROQh4iPeDMz7P4Vj+z9u9yD6LM+FL9AIfyiCEAsg5
vn7KUBoP8InMuByfVrjZc8UrdjK0necjjCvEVnTfHkRQXoskUQk5aaeGWaERlWc9
1CPI+NaQpu02Uj8uPf/H6jCPM6t5DQBaGvswWnQz0ghBX3I2bphLybvV80eApmO5
7Ncm59O4k1vq2rb2XF/Zvo5eHDsoEfHwqskSLwUrcqSV7Z/EyMYY16EB3OYSdwUm
94s0Nu02A9K3ea7b6o7R+my6vxomZFGiKa55GUxXEqSp/0P9vqCp5nmmzEaSSppO
AI2IvSUSJqCZJf2/NVy9MGys6d624EpUcfhfwkcQH03MBxVNHXH7gDgvh5FUd1E/
U4aY+Fi5FULshJFRPLqiHTAEyU495Uim71OPHmWBdqqLbBOA/jY0O5foFs82KmSO
lriizVvYIKh4NNKfMQ64ihuN8YDk2h0fSOAq3wkf1n011TPRdx5eS7XJiVZqwCTD
3nlzjRrIXac+7oW2dK9OKjteut+q6SCoSlrLjTj/6++uHFyQpWJKpU3dcdW0xt4g
OVPueE0+4Tb3/zmwEogZW7QDeV0yIUieKd1F/ZoyyUGKGRERYp/mvNhNRm8hzZLA
guuN33J+NwAIJCNLJSRQe+X6Wa8yCepRhnBbwXvWsZRp707XKm9lCpIBrKbH65ag
7SvDxVATrcqp+pBNQ+ANmR+4OUoT7fmmwOLv7wx6oRk51+b37/MK8ysD2BZ9Tt02
rUgomzelgpNA7NwWtj7lvkdowiO7HWG0ZjvbIQ/EEapkwLQJtO+ChRrF1IPnASoo
J+Jm2Wc6tl829jtSRowvNpiJQ+di97KI9/ZqbDQ5Hqqn77bmIX3JfOegStqTgVBZ
aSykCEmoQhNbMfnCyrVBuMz81NUAkMgqkuIkxA0Z7YiXtZWfEJmLSg+eHZy29U/2
fl9JP3JOW1T9eS2U0IYyX7u7rOMaWWhLGxsUn+IvQ+2+QxWp7xRYBg/19aSohLFU
VoTbx2G6yqVEp8vTGaWPm8s+5jS106TWacCkrvMizGYhvAv3s9C2pOlA2MiiMtI9
asJaopN+pOR28ZTErPLEuMOddNxO8yPgnRGoXQqBzbQKHmwpNLRl3HxR9PWwc3vC
yzAyOXhwf4kNaXix1t52HSQ9bjhn7Km72VlQ561PbxSxgLI1n0F8liMpdZ9Vxy3X
Bs1+tuD8MivZKhY8hmMGiZq9UewckAfQDPa1+ME0GkqM3ZJlS72lu5m/i0zFx2VJ
MKJh3Y1CwHVSCb+ZqcI80cktFzVam54oVtbCKSAYWEPlOzvo/mZp6FI2HPDiOVWq
X3ifgK2A1t2AZY4IVh9CpjxZpDkRtylujYb3rJ3ucuOAyA9qafHXdCbCfkKT5Kb+
YkEqkSEmxyDdCG7t31zCzEAVgg6zWoz6qM2Tkd/YrIi31ghs1opkJQWmvN++Zdt+
Q2CHRQqT6SB7werxPO1X+HGqwACCKbkemmF3/uyrIuRHiHFMuA6NfmueBieI/0q7
us6Mz6EsT2ecXqe6OGARuxpoKOxGZF4xf4VRsAwHrUpbAvxa7I8TCXXOG4dBbaKq
wsZrqqRKff10l0OLgykEw3/v7cc6q4j0km675AXmyTgnGgzGPaVY/YNjXn53vpF+
a5ZNKLpoggHMpcpYPKddHaAYzjhH0k9LhjY8t356L4Izz+YXAtZYgWHgQ2sUE8Cq
Kue1tTiNXs62tyNvIrdDIc6ofslDmY2VTOSd+Y2voAG1DuSurSzji7TQlPBquZi9
AhRLMQYdllgJmwBoYViktyPuRvMavIoOJqZHtI5MRGRRhydpp5lfjSD3PxseDEQE
VLQ8KWXFYonI9eUMSJllMryiUCbBeYRlwoa3ZxbnpOuHIG2MN0DJ/1iNUOMHVBi3
na4F6ZRf7y3rzAoHVPkJVsO3wDOP71eYvG2tvKpJF8Txw8Pav/wE93xCyG4aUQ/M
Bz8K2uWS05T9X6OkdqX6BOeML5GYfa7sbXqbfNJORg6eTvz+vT/2/EIilb41CAsq
yFsM4waS8kNRuejKsPV/kQZaF9QzRLQ2RuDLi4f52+c8ePxsA33/AYlLZK7eTEyn
PExtmqT1m+D/yKlYmK8+ZgKAgAc7gTj0CxIGk6d7VufUdlEkeGbVS/gy9YOjUHPd
Vk3Sn6N72eKlDrQ7FFGQPqMnn5IkN84JmYI8bLT0VY3zXJ72WAdYPqecX1mamPOz
qXM9AFn15aOcIChlkpd81nujnpO1FXXHTXK8WYj5tFDQYaWVWNL7UIg/nD5dDaY2
O8kzRiZC8iQDc+yoVX7n60Kg/Q7nrO8aBLhjJYZuuopR4d9jGj+aFKz5Kst8Fj0s
+flDrf0YHEzZrsi6t4jh9xempQvCuO3++Yt6l8vKfWFpEirb5FBHQLsPLEA6sBWL
DjAEEON4E1eig+Wzll9rNhe+OTaZYO/1YyfAKIpQmrt95RTquKh2tLS26OZO/heo
J3j6tKxHzZrgo72GJKCL8Lh/imK5Y1YZwjZHzu2xJWUdVr7kbyLZ/HAWv2L1bEWq
ujqjcyNZ3Z70inZo1lkYWej9DlQAOzWgfX2f790QMXMdoPhB/4psuksUmyrfDKV+
GsCe+UwJhU7QzkZlce/vFvRO2T3cSNtZYdl+0nfncM+zZ/nfeherpehnMCTDW0+G
FACqV78u2MSMCp87OjXjR1IWbIjzcMZe3fiYRiforaJcR4qPuoSSJFQbpXrWNbeX
utdAs47AJlL2VZwX/w1Boh6+/S/2dKWTjTySoimgKY8OVG1jWllUXXrFaucu1taX
axjBZawucBRniZvsZfRjUaC1wpbdvxQuKjk1sBHb5dmhw5PdCAZGDIclGXHafyXt
DcA7KBpJ6akq0qc4NoVNtl5I7kiYtNqt2TQpFA1r1gx4nYMukGvF7ZHYSJVBmaly
XKh/QRy5kHyQzIuOYYBNhDus+JFW2tiPDdyjkbxfPR1nQSutqxAldjakIPLURZPE
iOgKfGHnVeklaejczL6xMmuaYnkEyJ9If2qzVUdKNxfie1XvM3izqOJthJujB4Sf
bqSstqnK0b/voOdpUttybeigDumWi1fSiE85t0g8IWqY7k3kizuUKvU2WHvSK2ir
q2khC0YhwlvMLfb1exIQSO1GnuWugniSw187VvMsft3c16AjUulRFqiDGugL0xw7
/KUyKH+O6f2w3mTDcDYabm5ouQT0TZ0+33URJanogpt8eUYjrnMYJFi8bXPsyA6y
vCMfu0VEUAjbKmI69sqKXIfTL45Y9ilTf2YZM6oFNzRPKaqWgs82BoCkMf+/BQ8K
G0zkPwUNnvCqMz0x0v2GPBokkW2+wv2R5r5E3w4BqMwumQXnU2j8FdLEYVamJ+np
xy2GZ3KwvrA3a9s/3/rT1peTd15QciJIsUxUROBTtVsdPxm7QU6kyIyxqT2uJyo2
4ri1qQTKTdFdBZ1UVcWV5Sif72cQVItRLJVu0DB1nzOH1jBbOa+Pc5HHjKUjJPIO
LmzxoAS2YbKRvWteeEPbG8oLcBXQXWQ45h6s6mgMz4m3VUaRRGN/MQoCJSb/LK1j
XqjxrYmfVTl+ZJFTbF57npIyFWPKkcyLql2wqs1mCp4caX/ihiynFBXgNnmXV98d
pAOSjyfsvJI/XHjJtqwnTZdnJqwBajFVsJSTezCjHskEnbQKKw/h28cM/74pMsJa
OosilHmdGr5INsOkDtpmQuk6urvDW99a3xEmqgVO3qWnTQCMNaNMh83FgTbQXwgi
gqkPqaFOpme7tkULdHfVkAs8lknE+nH0de19vrVw1VxywBx6ll+vlzMkvWn4JCyB
U2VpETxYoaGAEQyL8kk38gWMTyECKFOLl0NhqqJTfWFl8k8Z7UQsAlz449jguZuz
xirxzTaoBDHqBAwLMPcYpMxbnTuYBCOEsUsOdwc7J4ahrl3dfF5XXPzqD0Wegr8B
UKfaQ8Pkhm2J8HEmeKU0TaRgic2fZN9N277erpI/VtPc8uGbwCulhYcxZMUPVDWP
TedmzsejqlelkfClVePrXHVtYwY9BKMoVbXtP1e8aLjCmBXgKaTJ7QEEtaUTEBkt
b0HZ1FpcC/flEqqW02S461aELwedF7UDOiKntivBgNywfsOxohhai+IqOUyH8XvI
EUiQezg4NkMQQIe+F5dx7hv26ef8HcWfqQBy3QIgwwz8dM2NEVciOAmb+rAzcCIS
BclqQmWxl74n0XGfsW9KxrlD5IbnNR8LaKABsD/JVMyMlX9DHw+xJwmu/AY66uhX
sYeIzp1wn9qkW5o6AcYY22HedEIvnkxzxsIsXpVPjbSB7TKNTkUhtu3XRas9ECoQ
JWVmEdwAKdCbAiqq7AEgrD7VA81xmkafhjB+YTv2nEFiso48rcw8dWbfyRRmDi8K
eJ0Oksvn+S6BRdkIO75wVFN6CxKiRyzM1mIqJhxoxQvoJjQP2ADJDQwt6X8fUzm8
63zys3jWaGEuQeUAL2fbFF8fSIiBToMDd3ZzBO+DIZgq7lZtxa5HXn4CLVU4P8Tb
x6jBhZdKTOuR5P28yFcu6x/tdI/altU0ji6RCqbLX3UYu2IuRPH66SU7MVndb+pm
Qa5U5RhZlg2rkc494xVh/ieaRZjdFsiLFTMg2Bhs2vzjdvrNTJbMS8DpUs6/vUGd
7w5PMFMLjg+CP3roHYrJemzs8Z/XrIwc1rBydC4X5hZkHM8EKM/Lyi0ENUpFEdXb
ltVzmVUpGKm5l0pN9ddRoLSBWFuDY9qFpTwVyXYc9urZPCpiknS5MItHqqgUNKeP
7io5G85R15S1neOQQFGZ0fNCQF4NsIlDOIG+81vTEjMJP2p9Eq3eVe56nmP+CO7o
YROnxr28tX6OBUC+AEp98xBU/7GEzG17/EI/McEmfKBA7GThvqytbEqWVlxc2Fo9
zBbxu0YlBXPNvsngxpzuLibt4D0ung5kCoV2U1JGrwDPyoKmrZ3ua3tl0fU+Dscu
4pGl1wwMdLS0lV6gzuBATqHSBoX2tcd/6Ifl1J+1tOX6M/AMGmq6PqJDZGokOrvG
9eqeSb9OoYKl8SsUA3FebRYhJhM86+EBrU4X4Xe7GkyBZRDtQ9vMMfMQ4TrihlLi
YzLobKWvb3WGd49a/LYF1abvkgYluCiUTvToETSJCu2AvGNbfnQgZHZ/7BD+Gy80
cS85GiF+CUYBGJxlfG0plS/Y75/lfDzCu8pucKqEtojwaySzddOguJOhRKlrRk63
gjNy0ZxG3p55vfK+fDVb9fDxH/bcqd4HDVbbxZFPpkOZ2g6QhvxuOI3a0jZGriDL
IvLDqXflAZxApCBKY14kACq9vRKzHPVDdJPS3E0Ihs2d6aSzprO2PW98OpSWzsNZ
BZMPgQatKhfNGl4oyx6lAauVWqUx7A4+fL12GfTdvXxwIgyJX5K8pG+fEhbQtgTl
LBgMKtV9PaXCaOJKYLzfkWTf29ExoVnQuaMipGDb10EVniT4ZBTqFW3vNy/BfVAs
PIkLCHXqwJaZiRS6UHcDPnwbKIyp3iPOE/xeWBjpBn957n7HLnZ7b6Ra5iENZoeU
GREWTYThuxv5RCESLSBUJmX81EysRk0B1ELCrFfFRID+5VSrTZ5fzIFKU65AuoUf
vz3YIrXGuZCExhWCknae7yLdwVLCFfkGD0pnF4qWoPjp1EjqafJf9HbnD8TndP5k
FvlGjEmMVUSyMk8vhxND4omC9fmNWcHOh8X1jcF0nWkGT1hAjnno3jC0PMyNvC7M
2OmusEHY2W3581O+KqY+8YUYYpSQ5MXYffWrM87PDYNEqGbywYC8TjB+a4F6q6Nl
2JuJh8MTILSKLp81QHXqA62H2NSafWdnG8M/7+tV6An8WHii9BOjxrUh24goalnn
4blxw80UbGFs0K9zIHj8FM1fzHNg3g2DODDQUEDQHOjo/k5jIsFYX7P1VEsyIKEh
bvsyplVRM6bSgLOMfrcl+yZTZgzMv/P+bdk8tzoERERirTd6HbX0wQaomR8uhBEh
x/ZSjxAczCWV/Ae/aVzzo4QxOvIDBZ9JeXWWyGEhszpSm819n5Qd4FBhPuN0euYL
bGp5Gw6CAo10J58Re5AJD+i5Casgw9zVF8LkUI4yW5p/ZtnvnZi/f/j+w5TCwE6o
49NXPaH8FgbmHERDqidII9Et8eMRabCkdpny15qQuyNCiW82cB6lvudxhcmR4UMN
kNKcfmqDvh/xkpEkU8n6dBnPxpbnA0+rpwwN8TewXwop7oOnY2mS7neUjFpG2SXV
9/eUyHeEjzKLa+jTWQYGF4IF6PdnYwgdTEo671Rate0BaVwQWziB8pcusiwjGrBN
uYSKcEL2xhd8tfXHc72FOsdDocOQAJISISYx5+SFoOee26Sc9wLbs1OU78t/QhCn
JoH05eG39Kk9T85+lYjzsIUys8e6dkwMPCmLT0SF0n6c0GI95ed98hXzyf54PFOY
LUOhbhytehIhPkoEMrrfESnNt+03/cpdTKAKlCutoj1zoduFEF/ilzYj0p2YP+Mv
cJ1TF41KfLz3QbtdJWGH7rtN94fc/Mcq7UYAV2ztw/D44tOOF2NztV7DgvZRD4tB
GtZWhTR0QEUvfkglf14UVE4M8XOWGaK2ppVXU3+l3aRqwKRQzCu6ikVrTNAUUIQB
MGNBav9RL36L/lanti+jlglwVyCPpdSRW2y4BFM2+5ax5vSTwT1r9lHV3CKlSpIg
LQXJHalEEKvxywEmhlpanXQYbHRtMP1slgWKaxf1oCbCDpUI0Cf+HfIrbVA8fHad
AtxuPHIzzW7/DSeg7+ArgehNaYS99JEppnU7u69ny4i8BbfO6+eEUxdyi67yZk/A
hQWK64/zZ+GuQKqG/Xl2ugosZT7XXrZ8GS5bkqta2KznCsjp3ODJ1b1wNPE2nczw
NSGliHZ1lcKLeO8TPsATwZpCEe9joC1cCju4554UuAQ5rHXAP9lch0iQoGR2PvIT
L+9fwWG4zX6clvWy4Blz/wirJ1Mj4mABoYTU+jYkiGHbTf2kvy+nC25W5XTi/SbC
R0Qh2QDZ0FRGFCIof2cJpmgFnAWUYceemaBI6iMm85QShr7k3B2JdXqGWV+GLwJI
WbKbdcaQq4jCVON3yakq+PUUDUi+ezabPN0LgMmY95Rd5tYLkCzthwSRdNgRPjZE
+rWjnolhhqxVBJFys01peBsLappDQ4cCiu/HEcPZdZePsEoJ3BgYb8tSoPU3WV6x
sWWc1j5WSUb23hNivKDuQqgfxWEuX4R7dqZq1sUz46ZTZdjRSJfh/IaqnL8nYpaw
cGbJB2JOzcgOtViTgebLy3wGhlrvMGMUJMyB9yyY16bdpjo4b8KDVnTTI+yHrRal
wnXMgYzw3JViHkDnKxZ89/i0jrouMiSYLdL6QK/Ugsbd3RdqXiAaVZeoSzakPpUS
ioYItAOmv55jNmjXE4y1OTG9xdGrauXHdPON6ubspnZTlfdScoLX6gAZgXop5W6z
dr8jaXzER7vXdSuqoaKF5S03SOeE0ywgq7tOW8A85qExbDpEGgzRGIv4GZ73b8Se
DEFkhBVqTFrq8cf9383DHkP0LWUXJUykMAIlYNWeQRZ7ESXjgrqXHAlHijQqNTA0
I2tur49PkvMnOwI97HLlImtAx6gsebUZz94PIk5hOxJ/EzfstdObxJx+atj1gAqD
hEjlYz6Ys8NjRDiVWfiY1QW2s0CrhWWatgROhcgC9oYNVKGiFarh+hlielB3IwoK
VnRs20UpzboW3g5SeqThDDNs057sKPRNKq0kFZmDOxU=
`pragma protect end_protected
