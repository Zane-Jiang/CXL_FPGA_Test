// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
wHE5Lu/FSmVeVd/Nz1eNKjIf3IFc4Wo9zK/jq/NTj1nEAjrVLjRBURdvUn0H3EvI
r0/XOAnDJPSYa6WQSfpcUC+ZRquEWRpn3cnGrO5SJNQzbul+r4IFJXtmDAgAvLiI
nZbimSu+EZyQ/zRxB4Bx0JL7SII9oQvX8qFkxwVZxJsPFZ7ZdwetxQ==
//pragma protect end_key_block
//pragma protect digest_block
amSwbhMFhUY9X0ViKNHiZdKSBr8=
//pragma protect end_digest_block
//pragma protect data_block
h3kSjrizRb9r0ZPQ2fFOAWMlAqVjS3GI4TvApvJ8LIjmu5Tij5roxalkS1kUFBKi
JQRXNFybb9GmLLjoAEbF8aYLA1lhxTDFapeEvrO1lZxt1UsUjDNcufT/1LXOshCK
uFgGMOd0VnFlSYLQn839IgDAqIZKMFRnsK5SQheIXo+awiyHkKty9cGn/U9XjolB
tru2zT9e+3LcugxIPXLFWEx7SrLxcvIREN7yGvP4sH7vs/6dZ2lF2V1AlB/TGB/a
g34OvEppDBl9IacZ878//4Ls8mVEtvhpW2aNW/znH26qWFmR3uLY3cOdNEIwWx3u
588IU4t439TruivoCY24x9ydUA5yUhvTZVbnMCv6Sqzjs41MboikcsyvYSPrnRKm
Ernk0NMbZbAmOwWK92MAlfmTbUNzQAY48JF3jNaSW2kqBxtMB8wWl4nPsT7Tfy9D
AnIuvuzpJM7wAgXIQjxExpEzv0hoJEAxtWOMFVFD0xR5aasN/ujaBzN8BAeF39bF
cYONr55HTT488L6XnjNI0YZrWJt+vW+lDD5l6K3dJD/Ft1/9eAACHFPkoDDvkJ9H
Ns2Aja9OgaYdt9bM2RBOG6R2gXDuoW5EcSvniuIapfId+NN4APdkCgnqNFIHOID6
oHp0zkyKvLlWiyqfZsolwvMhDAtoG0/H37wQXKZog8ncMX9OOTDV7cj8anWIxA9C
HkBB5iF2pc9TDExAoRKFMNbImXBH4+hzJasPzL4r00Ayha6FPWqfc9g37XEe8XjH
QkWXdrTGFnKUkaltzB5w5KZBcCIDVba4jSZQOx+NKOhJ5tHbBg/7lBZ70hJ/2R7f
n88PTl69mfmyh65We3dBQNDzVJP2f8uD548o9Y25UotIKGAgbgPVkyaKlaf5uNKm
I2XtxBMYCoQO6CF7AFmYvgL0o7DiNeb3teD2V3QwojKUAXJ6LENoeVtc9gD+9fik
XiPbPt5XHWFUGyTo5oJcQx2pWxBplzNVGJhqGNzgDS90ANMyi+b7P/ksq7RM/rBg
btPeayRvs4unSarJSqWu+JHRUEaGdQqV+YPch1FGndqamhP2/T/qpc26jrAA0gkh
C01vs05WLMrnirvxWsIR+SdQZod+qUAkClw7m6JM8Ugs3TpHsoX8aHdQlH4ZLSTI
slfUbxUFmxrWEQMu5HItIv5jkXQ3lYZXo0tvHAFFXLonHM3l3oHehkesHCxZs0Ya
syTzZhhJ6w1+JadqQ2MNQSdpwdFlA+gIJxTNtlTakc9CEd4F/cQTva3t/s0YObRg
2JRLlBG5ddGVOaKE4zbqZxktLxRA/hGGxHs/pMbdJLBnAxsrQrkBa78375K9DMpt
SPL2NkZpXwCCKXd+0mtfCFHwd+trbBkO6SEpY7wu5KdosvgTuxU70qfF8KT66HW+
uSpMMEpuiFF3Ng+cyB3d6luNuv/EIwgrChh97UX6+wqqddjzRvlfpgSbYPZpjwr5
Eft0ziSRwEKrHxCT4Mbu612wxcPKkk7+usqqTnM7GUHhwkOvXThqIKScF2tTikRy
4vrvZOwewYOAJwrQvDNTcnpjSLrBpKLyAcBbHgsZlY1w2Bdtwct1nUV8eGO0tBS+
/uPB1cHNq3p5VmyqiMjU8wbhrvJOOuS2xibzB3HD+1lt7FfFtontxXtRY4c+pzU7
yoy/MrauGvZLwRQzK/MVZSStRbbwiX9rcjlMe3Kio3sdvyCdCMfaexFJKf4eg1SR
7rzMwf6NnOgo+2nfzkRoO8oWn03VmLkaLDtjbTC538PrJ2MQjbng2FjVNkdcWq9e
FOxHMtU69KcE6X87PlsoQSRY1MaTQKP14haxOFaWaPDaUwxoq6G7vDB3msBI1cew
XWb5Mz+TUynMxpTYwDQDQu/GgZnK+VVXSQAnltmEZsxhnCJSAetGDNDspXJaI0ir
5p73j0pui1jrtfVRNegJi/+B9sIcZ4J8EvJo/0zIXNdMdjcwR/Imlq/MBkCnfTrg
t9ISKfcpMOyd5A4avscolzCxb4Iis3CXPPxyLYMoPSFS9FCETJlrntZpWoW7hYN+
MXuwCsXV3Hw+KImwHfZj26A8TwF592hNWIAp45pbI3uKZpBILCeTP+ycv4jNVSYw
0UyYGeVO+OMNm78xEduZkxECTydcG/IanwoJ8unSBED6wQWrl6jC1AqICRDXMS/3
pLBjXAySoz1SdgHebGTKhYJeXcN8WFbaRpKukva1EQ5e0Ow9ZMtEy78diOv5MI7E
k+eAHEH1+c+zF+fmrWEzNJPs6HKJuAsv+6aa5zmTUkhtAyfzxHr1qpqBWypQpBX4
YieQK81LSoDxcpngWHxAHDZM7YpbzlfgAsG4L1wu6bMnYqj6uK6LtYJuM+zPAj+J
hkM/M7TkD2uivuKQB3dugQdDCU7oyFfSOHcU48dalRTtywNTyIo6XbRaDy7udevI
PNploKC+9HAQ+uTMG9pdEAlKSvHezwoMmXiKYYtcBUvEpZHWBQZzR9eHq86136wS
uFB5ek74VWLnlO27IyNFsZH5e+aE8ZwvnX56SXUy5wnWx0EsZfFGigce8gDudsqh
5Az/6RAG+nCqB7eeVj+4DdM+kF+24z6HWPq+imvOSEuslPK5aRq2ohB4l8cSjFtX
ZYyONTFakKmwOdWzH4nP4xCch/n3op9aiZRZi2vXmFjgOyF3biTcsOW5z/FWqzP+
SswqHLn9EJQd+1OfneskSkSNtVWjGJRA4x01BNSLqrsYqFu+V+7WAcCn8HjTgSRP
Thwau1yddzNs/MsF9MIcpOXlnhdxZA7kDpL9mb3y5vGU6BEXRF706g9K6yyVuihT
TdgmmWKr2t2+9C2DRHDdRX6d4fyff2xOnbfxRX2Gv/cVKP/ePRwAW5Oeu4lh105d
uluGZ2+8oXdPB7jHE1oMNJOsh6SinLtTdMKwDH+IuYWHiH9geKnPpPida2MAxYjY
wBp5zA2Ewv8VvNi8twWXmkgQ6cj+WcGs8BOrwspU1suQo9KcSg5UmDtpJ8cFzyKG
pJYWgdDynAlRmn8w7fKA6d5M+GWw2tj9RjWKNtSKN3utQE9/wBb11kmtTHkZByno
DJkXPWKv3JPPbAzKXTpbCDp0WA08zpXp9n4VoLyzknlRCXaHSvrEelU6DZIfw9B0
a96kDfqdvnzUNZpPefwLPh+fOvF8rErzFNsC83UT/3heBZNMbWEBFjunOXoCnU1R
2rvc1/ZZhfODmh+UTKohl+hH5e3qwx4qS1WeNhuBBF6VbhHIXq7pOogw4OU0UDK0
4wJEMBhsOGIs1IwVb1whOoD9HTPUpzfDMXOON+xZmPJPsEnuPIQnXQHszl0lSEBV
wtJaJ/FJ4DMljF9n2DiT6TY1+PaOvw9labRn0KyiPoYYJmrNclTIH2J61bCTStoH
Z4+VeUuJeaGvcZJ7MEvVlkYKx49DFtnRdaJL/r/yzmsRHNeoPwvYxu8iww3UbLR5
6nB8Zk1sE7X3WS1+5Jy89PzqgtOTXE0zNDLUlkpGAbU8qBklxrp5jz2GAw/bjcDj
ZwDmvdPgJTWUcpbjungmp7BTU5BGxcb2LnvmJfsXcD/zXafbxCaAz3iFHrXsQmoJ
Hj5/K+pSjHaPD1q7vuDVaJW74S6u2W4tjp2i5E3aJUzR0Qb+bpCI13J0fw+RQsjQ
hIaA+GT0+9xoULwWCOziGtAzEE2pxCAWAWDEVdhCgumu7gRZqFNjE5ceV1uEwA9P
CefQKgEdMcOe78ytXyMcCaWcdsXau1n/yD62BolGJbI2UZnIeRal6agFGczF1s8I
AILVy3MGrIXtUxIEMsNuUV945gjF0DfV6Czs6WF1+rn6EVM1MI1924wqfaZtccC6
QNgoB0ngfo7+n9nhMc+vIMmX9WA2UAB8+SqkfATLWCg4idTZtZfY865CZvHnQNlP
cu0IeEE3jweKjds92/sy7nVBnkPxhy+NV8yj/8uypRSAJYKrJ/o9w+qdXlzuxDon
gtBVEI1Ar4b0kDT//2ZOVpr7c93UXf+afBIcZWMbO+zstDPlK8k1efpx3mLzb1Rj
9OlKLDmNd/ieJhcvLT9NHQ5BnUr6QO5qsTQRS56FqFp+jrZ0j4tx60z+x6gJ9Ig9
HlS194Gow4VDvJDRKw29XFl8e7ahdBohWmelccIg2jQkYiAyuzckQ0tkJRvnw+Ok
Jqmx03EIt2DKNxRhS9zmBjTvMlvfBsThJZArmdWiSmT0mspI7AQXiiIKLWLcxkc2
cZ6jWqn4o3WYBMWLrBgettFRP49HQ3yMBQMzkWSpUjJJhySFNkkIdqjZZcQlYhcC
rSMhw5Ikynzb4erbG4PKlRmUfnsLGBfyXUz1RK0sWNOa+8tCWzbO+9c3AMTbaTR2
5sKzgRc6LKiBwz5Thb4/17/PEdOpbi4mldak+XoY69CzTUqjbaqSnYQLW3gVm83S
T3HEdhhJSYjljVYwOeL1SfNnZRHUb/CaOmLDvB2mf8zv9Rg40tmAjf7ch5UCuxrC
H52NcLGHcpWeH+y2UHvrMM2onpFrtgNT0dLCewiDBZs13VQlt8Xa+xVTwpBReGx6
BEoCQ9Wm+p//n4J2dp/n6aRGIkz/XXA8oeoaV5L0Og7V/Mrib+ZrUfEAuwiydLqE
Muk3kMKagHqXPI43X8ZMCc4GPMHl/1orJudlfDjrhsplk8I6yybW3ILIZO+/OhtW
BbksDIy1xQ9a3FRXEnTW0asiiftu+6rgqe/vUbRE3umUpdStojwCyegi2KnK5Xbq
SAW56bWB/aMq+CHRaoxBy5OeDr4HgEwq76JFG6ucXaK61UN8o2G6qTjm2K4kzLUN
/j5Yuf5TlLNXCE9xpP1AYcunyu7SvtckwdD4+TydlIorDHtN/5ci/xR/rCOzWRnd
rGEGHFSpm1OLl5o0oM7Y97tk6dQRJjEtn7t3vrupoGfl8QiADtsxAVrC0o6aplA6
D1s95URwqzWc+B9dzsfYmBluwvJLsrBHhveFXuoPIBKmzZZOpF9esg7gzi2bAcmc
EIoWAU3AgGbbtgINFrW9YYpQslQVl5vCVG/q1MpbdC6N82G5o400UMkeQxBXeqVK
5+lrT7jGzVDF/mJU2GWzvBGZKS0RoxVsS2uMqx9STcMeclN1AB3ExTZeauLP3xCN
O6VCQN6ipxoKPAOsue1EiIqxh6knFSe3NyXzR9fgaE3nvQepNSWvSgD/+68QsJht
4yw55kksfHe/9Ik+/ZeAGZzUhEQPfCPpD+CITcLETTmcv5nI9bnGXeKKfG6r0KOH
Jhaci0RV4PJGmWZLOPW/WGvahy4EtZ6kriP88sLzocTH7PZ2GoFOXQB1tDf6/3CN
i66ibfyFzObwgIcqP5ZGJNfccF/fbrZLOBUYgoRnHg3bCnjWSX2fOv5ZgZhwZn5v
uVVIyIdX+PPDyVwFqi2ijfYiOszsW+Py5+rIikI2rCUupUp14y0Of+mCQRnlvto/
U1A/frhCqP3AAnUVgaF2g4trwH3dzRADRLL70eVtUpOXJS+KiKwJxRlT9ahmjFvW
0Snvy/ODv5xs10eCafpdAVMuaOC1qq8PaYizFPsb6rXpA3NGql4RbV0O2KKOdpHL
JFPBiCVqTcit96UIcWGCXtXKWWtVPtiVLK1Y3RGVCXblwmtq2ZLsqPwAGSQ9IEg1
igz0P9Yhg+t8EwXN3JtU4m0dYYC7CPpO3f3+mLXVtT1utj4teT+avMnUxBFOCwEB
C2nw+UPic3wvsZVaQKwjYvy2M1q2necvOkH7wojMlrGhgG4Zxvi0PG8CpSnnhhpc
On4IsLSjj7z7IwehFZaTb+WugL8/fB6T0/zI3MWM71eEcbzpaplU9Uq9f4DULjoS
XXVFtUyqaogT+aX98ndUWD2L6hKG1xEkgMaf/q8smEmH3jpFeTnh3uCGHCsecVfX
HBpGL2eV2bmTLupbVJR9e8KcDBWOPdz8nlqn5GZcxkYRq1gSMq3xhedDvkqHl8d2
e+V+rSw5P+sawKlfY5F5v2omnKgy4G5z/4WCkAke7Ni7Vl2K0lPln9XPihIbzwaG
IxKjAx5s2SW0kFpUmeMbY7bZp5ls2f7kqWmXrt/+sitW4sbqmeFLycNNKEvaRToK
EcRzsmfkf4jSJyApUlocMwUSHzdoJKNktx0H22BIVAlVpZw5ChYRyL66HmpsoMmO
vS2TNr/5cH0OHve74uPeY2cyorep+O1AWP45ffXNfTiAJDvF1iGUncZDnK6rybmS
6Br3iCLLTAJICt+9BcKRNLB38wtVS+2wJYGURZBrY/HUB+7/Jw5nae9mNGTsVQ7L
iyn+bjjPyL4sVsYQShjNcZr9+tYbY1KXk/ib7ro1syfPSo9eQO9LQ9MGh3ExcdwD
PazsrHXjhcEfIrKpw875y2WCIhVTwvi0xckGAMRI+zp8J/c2KEytKA6mi5odKg9B
z6/AAzEteWGZWFsramM+1mlfqIPAk8Dvc8G8L8bh7e5Ao4GvXNrP6KyJQYUgnEoP
8a2csE4oxW3YFimiuLS1s36UXLfEkNob8DDnY1BQFGXbIy7Bl6ReXkCbkN9Zm+AY
fqQqEAu3eGunxUk0r6A0DFnROHTY7X2fYqVLo4jcjp40OrBeVeb5Iw0YVK8h3PK7
Mvut9pKc2uWGV3y9OsvFsaIX4hC8wOVZluVxnjNW06qJr/YE/x0AQAFAtId9N5KM
7YVfZ9/FC/xFqzeAzRfXV8ihhFvs/uip2nILO/cmHU0y3Cw7jfSuEaW3RgR5XwMg
Z4QAYtGxvu9KytrXIXwcPjUGEtiRQrmBllCNEQ4ywnYYT4OCIZ27/NLesikn/zZ3
FW47vey9HDKTLzRtL0vX40qekXNP7cKqavOBwkWduRW2StF2oLEbT0GIw3vBOGwL
V4vuNcdXtWqCI06LsxDjHULeq0luYgfngszg1+Kv/ZDy/Cy5M8XdqkYf7OdGR/Xz
w68YIHa+IdWNKlg8iZyQRCoEzrf7owCo0ZoDO2Ph6+TaLTDmDvFWGeOSa4Wpad+p
gtBCn/zc+pzj1Urpk96xUB8NcMLSAzeHYiv8r84xKDB5ifYRX10+vhAeDDVxR4TJ
BHBZpReIzBJuge84gqQUi+Y5jp3VCRRlQcDmis6ICjBtTMOIKdP8r90Va3VUckGs
XuDCd43mr416l/JB533IwVQ/POPCQ9YEPt4hB+FCjbSuz02xlX7Af+dmDPHkOhdw
xuNr4qWOjNRsGo1DfDslLAdFySUN4U4RQF3hjwTmIT6EIW7/AnGYunBolW6tOPtz
xe9YD7O55x0Wlp1Zbp3AIKIg25S4bI9m3mNkaDKuDYXhFYi3WlwTxgL92FyZNQe6
xvPT6LbP04RV6wmBHY052B2mYsAJz9OsvVfsqdGdSMngaeYHXucly1DbYPpS0E0g
iWrCUOBQW+2f5JPdwnb0WR1VVwwNm7xTzb3Eh6XXdfdDGThJtjaazGG5LZqhC9hi
BSQXENJp/kAB7Vobm/dhL7tfPIKu2cHGDDJiOtCmShL/VRJ/nGVntRtBXhVNpKwV
ZR9pQkS4tf5qQc4eBsLJyvkPRUXkOEhdPaDyLqcnYJ7U5plC1kuTUUN2OyyNV7/J
jhXMel8seYAprPaq8syTMtgLVUw8lzms0AUt+dhmosRLo2egv3YK6kes1NG+nNpH
JKUxFmy1Orm8UGtJ/H7/7UW7S7era2Z3jtzPG+ciBvk9s/enfsz11f3W6a8pkN5u
+7U9uYB+uTwCIs8/a3EB/YYGFD9pCCGN9QAtCcXxYAcvEhoy6a4VqTUDba+bRJUR
rCq4iZiv7eQjMpSWe4SJqZjqcjl6iZZ4F2jPihfuk6UnGhu3lzqMQyiivs7UlTZt
WpFZ1PwjyCbhFYkm7Y+YhmyT+eLlW0C36nYugFwBw+tK1HxVj5ekGxE6JqRHK2jx
pJg6ap6p3P6NMEgp6Az5FmlGCU27jmxuZBqFX9BL/tRoSUPXqgjzxQc5coIL6EyM
4ja89bQeQG0KdHFvOWCsUlHz+IGToCDApL7EeX7KjWx15xy744/pOg1N9/6sJy6F
v0LGoyxDK8gqv8Kt/J4rHsKSLC/xcibsC7cWGNvcnOFJ3xHVSKn7j+06J7jbKUdk
2eeOnx5t+ZKrPOo3cnCyr64wDR1QZd1U5s404bjV7fiZS2mU9R5iUsqRLU+xRBzK
LdUJnbzj8LWVBAlXS3hMoh6NNlb7yuhKZQNfSwzA8ykc2giw2qfGGikn8BbWvmXo
TrVomQgmuUulEJ13uoR0wgh1ganu1OkuxL4X/OFf6e2jDuALEBoPvpbGhB0oc02h
+WagtVdL4RpbvPfNTaxwmmojswsaJMqG5EDChmFfn26oKsKkmMSUEXFsw+ey3Bqi
Pwy9mjfA1l5baIEM/dWQrKupNdcTJ8TDLCjJScK3bTzGXbZNNVnZm9TtfTU3D0o0
u9CHGAWz6pDfUSMt7vLZ7JwPOP93zaJ+8O2DuI6uL0xmgeO9Gp7Tcm36AyTOs+lI
yx0kV0o0r5Yx+yDSpJuNWu8AQNelO4iy3PzDcivqduGTXSD02+LY78Cmf4F62L+v
fR9UX9uXxFK3BPF/FtQm3VHHYnTVYswC9LszZdRQqGSulrag8ARdC4LYEpY6NJ8u
kUYyAhKNr4MyWZ4ukNcFX7CFnRfOdEl3pB0/U8xFJNDnjUCukVBI5cM2emW5PrbL
Zkk5Z6Oe1G5tMBpnCzQrHPZmsMQ23o3RyiGSfz3BQUoLgR0JNtwGDH9h/SUsp2KV
0citHWkFi1TK+Yf9VRL8d4ob0ZxS8g0pLBpnhPWk6NmYfStR+Y873IwGFYPSnlOI
qbJZNugwBkDga1B+5pMUmDNurIormIVbCvYW1WkG3VYIKSO0Q2nWGrTf0rfox/Gi
ELRaEz0UUF03uZDSZTJHHKI7J0J+CgHrfcpuUSF4K2flqTOJ5OfrBiOLtc8VSp5w
3qPGUzALOFyz0nmvXOPs/aYGzOR4eb4lXks2PYQ7/kkOUzFF/wEUosQrLEQgryAj
tFlRlqXUlWecRJvPVSfUWXFBdwVRf+XmIy8Adr/LB8IBTzsA6+FW5y3kRPvYpJ4s
H6YdkZ7JUHd6hkghBc8h0EoeOHxzl5enRi/KeQWu5Dm8Kr/4wmVNmynaLSpQMrZH
Bjw6EvZ735T2YdWITe45rjLqXNK2sfATvaqbbp+vrj+mLnF0qsxpXhqnYnQA5yKS
tbFogCINVh3qEu0uzti4T9wp7KwZQZRqQ1LwRpdqgyl25CLeEqVUqaNBC42Q3DWw
bCia3oKVDt4tibIn1j/xLDzJb11fNaZMQcVfdH7AMwe7D/R85KgZDZLX9g8iAU4M
5YeNLZKGR5Z5bsHyM6gQUuCrQWBSaNp3MZn4UDRSEy4LaDDd9/cHTG3fC504Lqfi
R/92cHcVeCIIufJAa07bfRrfZIwZC9kWQZpQCVVp/e3YUUwi8l6yLB7B+UGFOGcY
IGYUZxCrB1Pyf2ckjVo88Bc4COJB+SzVg+HT8p661RY0TOhxt0a7PGWZxs8LCw+0
wxqu8E/k3gXp3LA7y/WDBmLX+148a8LDJ83gUOGCibW+Mvnpyj74i8DEw4ocJMWE
p2OixaM3rWnDmG7a4A5VEE9bcQDdFXyKIAxHUTc0ISuWAjvsR+k0CxdEZ19Vkfjl
G/NpxDihsh7xldHN05uSH4N0j//pGpfjFnRqiV2I7lub9xeiU4W81r2z0skWJ0kX
T0g/PoI0n9a7CWcZyvCcxhJUrFjsl66qCNSWJnKhrrxdqF9llx+0Rsc/WqCKyfxb
0Y/a4fYzmRkD7buIoSQRYxAP4M7aCpjNPh9s4duur2VDcF5dPgxLaifLQAbA31GQ
2Ou0hVpWG/xxnfthKhIjQy9HqzXZN4/aLVd5q62AsMHQPWYEwBI7mn4OrZcSM4o0
uWBvXRJi/ydstGoYfOaxfNaECVYkk4i9wJ5/Ezq7iiUttVOJzH6GZvIO7S6PjGmF
d15QRhbDQxGUWjYn+K808VEtC4RxDPaAbTsT12cLSKRMBe9LXfY6hTGT/NW8VAqw
BnlK3+Xr9vxZUg9zkMvF7MEwPyNuGsP8RSKROEsprl9mgxtVqrX0XdD3HNZWuKpf
qdgFxqf336J1eBTRDvMAoTY3qIce9cUfLit15uolZw3c+lWYF+dhfMymmnnsAz/z
iNaHoJtMDGXBFXc1OazMQ0CAnbw7SY1fIBNCJUfjEP+oGFe/QyP27OYe6rasbOOf
3keS8Q33K1+NNM54lGqBD8kgb5ZcD9nIff4t/19oYozt1tkRXwxN3rtqfkSllB4G
tkY2Rd+WYF4Mfl+fG343WGM7yP2m1tAnydUzZKJC8pl+nVUXtiOB2ZyoCFqJs3Od
fQe1wdf8CJByLhk99gMtvrCmhGYJ4CoctF8VeuDFvfxGaw8sMxNoDVZH4jPToC5J
LlXIy0jV6GQR5spQWItEQwJ/P+i7k2OcFpjzEmYSwZ/4Yk4OYDtq7f4akX+LV1yu
zWfUPTJ79KD1Mwrzq74MNDxbs5FIXWpby7CrTtRMfAMdyBo1itzyFc43C80RiAl0
2R9mMkPkQvhvvXiASXdqymMqp9s6QKwH0nRlHVI45VT3cJPJODMzJ8PVveMVku85
x4498WyrggGR9BWdewyd01cAv6HNcT6i2vglNWNJs8Xw07SIgzkZl3VPSVA7g5UP
LgrjIE4YsuTAwBu808pyjWFuPlXm2GByettHFwMEqkDV8y7cAvr+L6clHaiorUiI
Bie7MjKUgRUUSPfVahlDk/gcuQkdPVrDqyR2/IoFYjRKzBGNzv1qM5h9MTFhRqAa
4CpVddQQk+wJl3uCNd35XXTeP2XRT/bHu/HUA/FB5xLTJutlKSgRV67W5EFMi4MU
ng+c7AChXDaCWQj8XPYNl3SgqEA/1N+Od8YlB/Qe6XVuIUerMpWHhPqvfPZIbdtO
vSKt8ty/nM9JKoISK+zfLykcp2vv0vyAHjW4sUWTbVTyh08Tuhr2icjKlzTWNcMb
6s/cmZktHOJ4/4iDrDWvizSu+orrgNG2BzhgJ+8pbKoHE2JZsZd0ENRD47EhqjGV
gjis4MeHbE0JVjKv+0fD6L05wnG7Ghets2V1QR8R/x9svkEfDu0oC+x9B89zlYej
DjeTwUx5/XUlezWGhY5WEkojC5LYneGV0p4+ulr8AE2kfMaVDTdWDzLz7xPUHGhS
yEf9HYjOP35yOe535drmYasy1RMWXjhTxPgAK/gOFDEIP28w3XFZdwCLqqyRnRqF
Di+lL4U32ybJQges1ZW+iBa39g+lYtwH8htHFGjMX92jVaXWCT+82ajQzCXycTnc
Ba5UHhL28K+G5cUggfA2CToDeqgMZ7izhhdblQRTGpS7ze5dL6OluPOzunjES7g+
5TvJEfX7hpNjXamVvvtWVS2SkJEQarIhWvQc2JjMkLy99CTYKE5g7fiCriv34EBV
trcO3CwDGC72JFtUOKToejuGPkOInzP2YHEa6V8mLSAmMdjocW2w27WTn1/MTchx
V56QX7qAFpxUKEZkmCjZirSLmEMZRtlTqjnnBjjQ70IboO7VFhkqX1zp2mL4L/7T
6QjXB9didl6/GS3RiAk/tmzH+WY/hO5hVWhTROBrU4y0gdCyDo7JnjCwUWzSq4va
tdOacJe92t+BzEsjWB2Y821fSG4GZiUGIelFKdk/y9/fp1iDrNybs1QUYCOXbC8o
yct6bFlHLh3oSYo+9/2dUn13fUy8U38D1K2MYbfgNKMd/y8VBh4RUFrakT2Sc55o
nqhAWt5Gb0vhD/zUz/06E7jAyd3NyKH7+oRZrrOWPqjcDFH7RJHO4Tty2JZSBSCP
mEVtspZoiOQIXSMX+UOO50wvxUfoRL01PcO1WR4nehY4Jush6PEeSvhaJK0AZ7kF
aAFZmzxZdxYDDesrDPIsIPcOM90ne1U6W7ToyZVVru/a4uTJXn24CP19i6qZLwVC
w1BUoYU4GEk0q6xuIw5UeIN8rxwpc7GJK/uaHkv0mEEib5WT1xxaZDDAI3YB4FF9
aiuVW7OuX/jZz6lIdH+0nRMau2JEerxmgklo2L+91Urbg2mwe5+klGUCZIOhZJ2Y
16grP+qdB/YWGUFoxZ5KbDdvXTJJdLGtS/w9usHZBPHAtD8L+YHhSQjyWsE/7kXz
O90WIvRT/hJR/qYJQvTDBS6cezZGH+v1t6WHTxfEIRDOul1yajDpvVF83mucnwb+
VbVJHF9Iaxnixhj/MEBi20Cvn3MNDjV6MubIAul3sCK/OoZcISkvAL2hiFTCXFt+
WMoP4Nt8U+r5qhss6cq75djgssnLfF4s+7RyEQVfz7Ix0QVFvenuZCQq9OOL7hoQ
p6ryb1on8OxHImulzAErzllrGtxWwlfzalhh11AYfZ0ld0eys97iIt9jX9pjD3jm
HGctVy+9/k4LhLE9scGqNWucW5cFi32d4C1ElaF0tzyybzgV/VaUisEFescOzhN6
ovG6/PQPjnRtMSXn1EACs5/lOw+FV1Ba6KJSM3O5vyaNAo8AN5Khjv7BAMUK9zls
DL0hBMB39zU71q0wKw4B/v6gO8dOMDV9OjycSMDcslxbTKVj88wuKzi+8LCeHI82
HZjuYctWGMSkSh+6JHnFRvBqcSjt7MoJlWk981goMG0dkVmGGOZpdnxiYltJfniI
H61sgUy0fqFBQz43t+Zlw3LLgjGMKIE1rsi/0YXwpTZ9xGCoOXOlY7FCz8X6SaKk
iAe/Q9jllAFvwbX+lOpiteNb1pxzfvfEFvdN+PigIEi7nhChQYJy+ZDAS/+Lr3VZ
HC5Blp/l44bOO+gUzJ24UERAgJ+u5pxSvwIcDpHtyDzyJ7G80v8IB1EfcfXpyVrk
mRvvXlQuB0eawsjd4V4SSH8CcZ+w27WFJkC44kilMiklOtozn80zo7AVXO3DZOoS
UBnwvTKPPM5UGaXho839cXcxcOGIsZ0Q2lIq9CWcAmKepjG8nWc8bjppMDNdsTY/
uBOfnWxtcI5uSW4xUOf+h/iaI8yLVOCoxbtTOOIp2fXC4WohIeeQj0JoW+776KlB
L+KN+aoda8mTj91ppTN+xEJ1+mKUXNu3hxasJGsvUWTa1tHdAj4unF1d5XOG/p9m
O+FQtM/JxUQzNqNPa5Staju2s6+/YwkGTtWbBOzJ0Ib/gSqIexusT33ofiYzaWDI
5u11RY33Yo1pVbb2imt0uHQ90m0XelR1oQca9u61mZKlyKx8l66EEn/+iGYbwY1p
DCQdAOEX6PE+1ldF70owpSxmHt43WFPnRLtRD4HmWXqKMB8nYry4uzG1AiA9ju2e
JEkbidQgdp2INaLdUztVq0nDiEFnsIB1N0haB5Ebxu1UjwqfNjeSgP1m7klbTUkm
92JUBrV04qoWQGeEOvi6KnEVlI/9LkXhKBRMQXYx7upJdf17VkMaq/uAkwm7HECZ
DODrKkaSGj0lyuKfA77g9j3JtFr83oBos4hmMA0HOWOF2fg/ZUTGp/Jbi1U94v4Z
xTtGUDvfK/O5GvOZPHNn/tCQMdLcGtY7rnIHxsf406MF2qlzpnyMRNs5srhsH04P
hic/T8S5a8aDNMqUdGNtOiSJlIq0dQI8Dqrm6zWsi2Db2ZWKj84+rf2e7606ET0P
0imoV9HAxTXoCb3d6LB3cQmb8LUl+5NosG7gRCvF95kT4SmaUVAFoZv9Sy/bwDg3
J7pSJLVsHIoqCKRPcq+NumkPY2TRigRpdjBJG8OLFJ9yuBP9JMk0D5L1lUsbuP/P
/mjTeoJnb9XV6YMk2YJovXX8yUfauw86Ltzj04QIvCdOrlMjScfERDnrq8tdZ93E
WIpNBdEKiCt2+g3EF0zWvGqHAw99nVIDTLRcCcxK78Zj2J0G7UK+VeBwyZL6c5cA
ELqDE6QnbhYydMiHKBqosUlmd1LGf3ptg/IP6vyowO2OZxyX9LSAmP23cI5kfErM
USZ0IJOpoJna4T1+MlrP1tqJ2I19zKkzphdBkgMhzlt9FdEeHIXZxL2FbHR7R6Rt
wlly3UDjqTM+MR83vXKwj6A78ae9MF//H7LIu38Fj6nlouwd4BEIkHrZhNtQyYDQ
NXkOHCDWAIC81KFC28rcC556hI97e0Hda6Ud6w1EVEUtxtLh7uFFZxfE6ruvPEPf
AUsHDA4UWNhjzUPZ+ezUc5BM/YfvxWIDSlLEYU569mNp/O5klwCyX+LfqDeC8kAq
1ySksCD5bNFVD/Cfk1a+uTp77Q57bsmT64dpAqMbD39k/weS0ReK9knzZUGRNyaG
DY9vamlNIpDoFCxWTOmXcBrMCQsLP+XaYOdZKgww9Tx6FF/pbw7dcuZzL6oBs1ZE
VuAZ+XbpiF/ViHlmMoDmD4+Wl2r0Py45yb0kKBKwmQSRwtKcp3BSIJY4wHu8btOR
otRXng72Gkctorf03nJdtmlmTJNgfAVA2oPCiYlXVLKYJA4xLG64wA7T4ZuTImzb
L7XxkdYalFh+VeWDKsfmUxCydtIYuFox2ykViH70JoAG4nAfSKIIUEXlC8H8A1Ky
M6t364Q2rQt/Sgot365enFShW+ZkqPkCLygDLYtkcAZRyXAU1xg69DcZhnZsz+Lj
0dj+z5EJvqnB1ttYBVIwyqeiu3ltPK6MQKDI60p5IVc3PnvjNS0xVVNmI7ot/EKc
ewS160ZCtJqoz9OwPoDix+OMPrgfqldRWdOA3NSK6ufnL5ZnlvX2KiFIvabA/dnR
DDuKsWPw2ZhiUc3lh35zvKRwu+8mdGvurMr+SKY/rbE7VVUdEa6c+sZ5IyYhzgJC
nIrEVy2E/dVSl2Fq7Acgo005J/7UB/BjrPaPidxrsPGZ4jSilAzAGI77X8wBoSQS
1Ogl+eTOE5NDoG2GSWKuVeNVxYd1zGP8cBcVhzL2lBmodh3d3v66MJ74SBPJ73al
bSSvOxH07YVvXbMlPLdaEUBmP5F8C0VzF7K685Xux3MRUPBD2XzsDTIdLdlxoSsA
VMcSmy52733VCdNwbYPM6o4Wtxx1H34ROtrLjuNbCEfyF5qr9S9P44KRAZBT5QhK
sfmeGK7yCEP/24GHB1iwwWtd9JAMsReByHtf4AgP6T2e+3d+ipKUAV1AwOKkGI5m
uUcu/Oom+ua4Kw3jooDWpI0iidjGaE5pEv+7jTYRJTvS5wOUrbKeQ3dBd2svtmim
fG8o6Fa1wpkP+PpDIt+Mg+nsenDYjpNWNwvsQg+IIPk/ll3uBtUTA0ik0/RggK/Q
Q20GK1q6LYws/ZcpsrJ8sVhYmlrex/Xb6XP2HJ1flG8p3xqUxqB/B2/l/pgXrLG+
/S57Nso28STlP0rAnxf1lRAso+/mJMNahuOehfcdkVdGMw1Uc67uLj9FYziNvHbO
ybNgOZbRWsuFumALDFC3aorMpvB0MngCHtpqZrN+CX6LtTKqFFVniM8WCAh3XqST
6EUYSrLu5kZjfYC0JtXLkGnzPoHM9i6O5lg+hCoy4IplhNcIukegfun1vuzvuS3s
xW9Z2X9RO5ZtnAFi7OnLUUubZ9R4Ii6cVWO3eI+8D0Cm/V7qWPDJSV7Citl41xdb
Hhj64FePHdWpuNEO47AnbFiLybu1xoT3bdUBwpCnuybnjFqxoPj1TMiEBWxhf0SN
k2ZkYCqw7qSWmVKpDx6nPnzIkWIQ8SCxcL29NEhS0rxhu7rQROekbCqJy54n8kbH
nYNDgiDKgPRo3qZUpJ8a+g4+p9HHFWDTFJfAhZ9B/PV/5rp7bCDDgSY+MhYLTf1b
PABW98WWzokwyMU4OV9wR2PEnVAf9tBlO+2mpr6ubG0IYoxGMAVAxJ1lYQuR6+8C
YQAbnv3f3wpbKuXv+n/2t7J30trOHwkRk6YX/uu6ie8AVCaOqIiS0zp611pzjxY/
sHbR8gv9cSXlhkc4PZzVWXT0zeATIu4hOgfQfh8dAfU3tYK55+Oz0yv/+a9ax0B0
/2QOjZ4cKnObRP6KMRX1yGT1i1ya3iXOiQYLHF2ST3kv6i+ef4t79VXRwb0PdWbK
uuAlFps7fmVzqZAMIIzVd+KJ8gVQXtBHQQqN2B+e7EMVbeCPajQus70g2m4vpScG
Gs4ZRNNlz4gosDO0S6kJ5CnYkUa4qIX9bB2G92T3jRAqKBEnO2SUAQuzHF1/2rEV
QmtGbVf/cn16THB2D9rrVDNeT+P7TXn35/fQGQEof+sekSN1T1Dudek95xA9EzKq
37rgWBdPav47KZ19uXeP9mMBzL9Q2uyDgQpKSURBfEhmS3G6PDY6Ak7KxX7zV18d
9CL0mqhU7jKPXyhj9Nre8ciXdlpIpAX+HT50fX0ZBEm7n9ocG5AKKML7TkAPLxn0
VtnMs0q+Rb0oVF45Q2MywWwXhxKFPrea546r6KLaKHe0rOLeHR42/abhxvTFk16k
btArBBO5ocgklXkXMyskrwGYlyHzFn5orL19XpoujOIziwY6dd6WuLRrq3rWxrNf
Vr5RDWjSdk2xCih0+ioqtobH6UXV7VPBiXPDid+kZs9rjIa1yyEhc5Pk59CSIT57
1RKMOHM7M0laJyGusbUn2mk7XglTT5GgBuwKwyctRUPKkLwXVBkKxVPQs0Sf7059
EGgHqbHSZlrtIAsriYOA4sEUt1OSLZQ5BfEa04mfrT3TeGJJ7AwajWkoxSU85Ffg
+lau2cS8lelM2JuYP8T0FV5tyu8ubjDyactlY+2wWUQXC53n449HxlkwqM/hGMmc
/8nuge0Np9FOuww/F+uylGcef7wb+VLqHj1qWyES27HnNE4WFphOaGflroCqpZjB
z6nMD/uoShH+yslpr7ezTMFKFs3St3qdJM6aumaHcmClTGNYEWxOPRKMVYtb+YLB
r9QlWnIQ3IOF2wNmiryvj7Lw/J0T0ZUmo33PVkT9e45qe+Bw2DH21HCkMzzsNQTx
ybmzF1kMAX5r8zIhDEl72kYXLJSjstNw6xw633O08RFFs9QNOxHRCPG6JIQ5QjRv
YFsgXLlw/kiL7PSmz1LoZdQM3fR8AfHm7zfXqB63Z8r+thPgMiM54Y3tGmtxTrww
vUSZ+d+pDkX92eBql83XC3QRMWAxOZSqu6zsG1ZoofKzI1hw8Mm7iXJitnYKOM/e
2gc0qNeEfvFOBM67PfRVydb1KKWhWx5SWjrStn5tOktlGxALyuwpPB76WKgJ6XBX
lSdv/YccbEmmI67NxNijtsIRYp15X7EAoEiOus1pkLmqCRshe2Gj/nx9Ob70Kpfb
voSmcDjHndiDtrEkXaNu9WXy6bdzHfKHQH+VwN7WVgmSOrSLbXyx9w8RoO13nyD4
m+U84DPEPhpWayxwAXWae0x4ELzLSqBYtgRrmLcXuo2xo7+/ps9DxsWru1moQuJQ
+g2rCLz35k8FX7Nk5rPuPAFHwUovmUYHVIMvRnyx2ah618Np1MGXZkJDu9X9s7ji
EGSdlK+Y3o+9be8vJq9IerABM8YZXEm2xA3c/b/KMeipMQosGol9YlCe0vs0C/go
Y2NqD7OTSGgnzs4VcXNA6nZrbnViaDv6EHB+vUpgYO2E4Jkwf1NEFjIAArU/Uunn
QAyvFq6XoNqG9i555BU6UmCaf1MIfoVh2EnMvxw/ZU+6wMZ8NmhYVhZWETuxjeH/
DRRaeXTOYHtl9Np+PPl6I0kMepCYHJyOdi/xlxPjbLOSh5UUb1UB1+vYUK8BiOqA
FlxRvTdIqv3WlRzGnhIBYbVtfhrgqHS/3ololAvi89y4q1tAJJaVH5ShkOefRPr7
mu9wr8ugsguYYaYkoL4CFNVG2nLeFOzEOgB71uUxqxHbzLgot/jlxcmUCWjm+IU+
/e7CmTNUD6ZS+Hv2PQ8zHwbn1zE+40CrnaMNKyvjpZCU24qR3+N3eSU8bYYNdQpQ
MseD1/Vsfgk97ZWD7wARBJu6BADSUpNJQDglDPQrgWaVzU0VBw5il5rEzU6GrzNQ
d/S7hylSDdQhuWu+19QqdMZSvUXvdKwl9tPyoKHAIgoAqCEYWoN97NmZ9kc2k34s
BaND/2o3KAg0mB20VzJhDXQzJQUsxpuAJbgOFHiZczFQ/Wum64ojfSXvVQUAcToZ
rblRTh/KzI0H3MaRIYd5WwmcJdwoN+Nj918vbrcQtjrGFClsfe/pR7nyzHEgQ8rT
o5nQ6dUxRaF0AEp6T0lUfWATYlTmEh4ueMcvHd2vUchPkblJKP1+G/Tm0MpwsbD1
7zjQ4rQwpOjR58qBdemz81tGpkrXULaNOHXXwF78URzsmkbFsixlx0VLz2aC6X38
KKyIde93qA0W0Emt+B48NZBRGjHY08UpvfZ3ixX9bEtJMYmesemHKPQijbpYX6NW
w1TBi0pwjF1dCAx21OEjFnm1XKsCjAWrwlgCooYPsxu16tZjqrs0k0NihiwQIzrj
AayPv3hdXDOaZEv2QuRD713/SrC0lQRCzvd+/PeCE0+ToZnvYPTUURnkSD6Kru3R
EgN9HydBD0xa7aW2mZSFBngoSiSFXVUiDISx/mIs5jebPjGYHBLJR8REjxTrhqMQ
J4O7He/TCvQJ4qlCqrgIGlOIlkp7zyYYYDz+6O6Z8sPPsHGM/916shZ4KSnne93O
MyY+GyDW3u0IYtYQ9pP+gygI2KLHIUnj04e0JW4urY0eVgz+1LiYgvNfqzjWKmSu
AXaYyrQ4Q9NHrrt4BbDom28V8rp51z5deCseAWQVZPHXxcwexxvrDlvvvToIElpn
hkJkGuan67UnyRkdnOXatVH6lf+v18G4oOmgw8Nj9GyGEZbNvbeEs5bLXuk5Kkqg
ilF0aH+FesBbwwI5CJN50FJxselipuNdMZRu+Kn+J04OyvsZmhJZ12ZBDyA0G27Y
qEj0oT05M3aa0h1bB4rkF83p6sT3QseQ3LyS3ea4kpYYvkc+vOGkfu/IadqSLuLX
5rc7G2+HKGm0E/kyf8UbNqdYjCWVjvcw79siIDO9LdtOxzk6JnSfovL1s3MmNjtQ
KWuk7WzVN1oVzOEjEKoQmFnI5DHQBzvxYsjVj2aEZsYxVcek/UIEtjxIzAOhGeq9
5YpCXAL1Vo73zcWMpbKLs8gvudlXFhg/35QSJUlGSVe6A7yFpfs82Odc7/7QABZ2
/fnrlQqUWbGdDOYo9+q1tL+MyPZyDLqiPJ2XtsvSdC4I/QjXJPbcHup7DDrSKhNM
roUmPJZYsGmcO95ooPCigiy6h/2oc+loPZuGjggL75CGdSdg5pKKeJfmbXt/csac
nAR8ykeYEz2UVQ7Nv4jpClrS7Cv01JYlP9h9xR1aUVTxs/54xhNtl3cO70BR0jM2
D4yT3aWofy8UGDHTjQwfoWeBaMo0HsjU8ehSnnQZMIQgLANMmfg6wvYtTsnjMWb6
dETmmblKckHb9+nCLB/THuWoI9vnelg1O1xH3xis8DPsKDQk8OYJiNR7osfsTbCq
/MUwZTaVAF4oMPRikHE1RWK1jsihxtWntlWqpu1aDhLU57kJTuF97ur6OM6FIVEP
kreuqg0bSUJNujpqQ9eLT52kwCAAoGLuccFUYCAlh3qVWmP4RcTNjscIba2JbNzA
pSA/N/2EEN9byCBAicEkgyOzkg7+7o+zu9hbApjEsSJFjkNrVIghPXFvSRo4c5qd
iDJrAWoMlewmvEgqXK3M3WVPj6/H76oBjh9SF4SKzC+8A96JwYLs2yrxRW0L7fco
Wb2SIIprZuuf4EKU5Mv8X87HtUailGi4wjSccQlO7+mpUC+w3vEW8wX7XqH/KBZp
IBTNLmyCGikdI/engYngJsPOlA/wyTVmwrDvQgDDJfOiXzjl0DLIk2lwlsrV4cnX
BKEX4G2916cjZHaEmZugnWbjFG+1a0D1tMNfGErfoLYRrDqbGlHGMAwYz/Fa/Dy0
0fmYnsEEyiQGkaxhdx0O8/VTML4a09r/LsZXJQLa2BVaS87+J6c/8F+0cO6qTdlq
P4LuJpRygMnegkTQW/D0BdmHyw1CGIL04PheOeFqX1nkxaM5vxahutnMq1G7atYX
kFDvnpF+yewKk2iD+ZrgI8iN4WMY9ecyYvn/PQf2AEBVr9wteioOlGNL25zzEjOv
qB5L9UYN0PoDtG6x0YhpDNyUyNxltmO54APnts/ZAIGKUSKqzZiNp0do9VUHE/7h
0llE07EvcDETz4tVP+Uhc6DjPKcH4NB6MhbRAX/2tfNSJqCcI7lJy/fVT7EXM9Dr
dDUvk2FFc8L/SOKFwZm8hSiguBUlNWKz65L/Y32OZvlW/V3siWeC+oUPGsb6GhwX
UjgyAfmL9SkbaygcmnS62CrPp/JrQTT9CRAUPtrV5w7Xe4fAKCSbLIKy/JOdQrwp
n18mDUGWULip+Uye0eXStBrvt//B+Azoa6R109cUxM8I8NAqovrF2eyh1E+ugc8Q
0yeesxs4z+IDkTz2KFVsoMHytTBpCDQp5JbwZ6K3bW6Y5xqJply40al/+R2E+YKh
LSpSLAKt1Ybc1m0AGm9JlxQYq04Lu2C5aLUbZ6eVfpRDcAVs6AeJ16SpZGbbRiPw
11ZCC3p/O0K9jK23wJB6Hq6HERg64s6XvMRIz8Uw4YzjCM+6MG03uLsqbUA8dMQ6
rGw+qsPvuEWyBb9vTueKpPde86MZwXYKF2/CvdM/3y7J71RcXSVlPbWll1Sm7Z3W
8ek+exnfjc46S2wbYxI/aG/OXf9JA6+iuiPZ7Jk+ZxFxzjhajFlQt+plc6RRu+LV
fwvxdBXmHS7Am0yZnUWuyrDspTtX5Mz6uPTjngKCPM6YHZHLGSFF1XIotSIr4D+y
u1PlJwMECYE0CBdzKkN9qVT3sFWF3JyEWglxZ9c/UxScHjjrsno2CQ3zcDmiGPpC
SDDt1gBnW7s0hQNgbACoLA6A/Ik742F6EcfH5GV3nM36Psolu0c6l5WegeWlJmhD
t44+LsuCLkTQaJdshT6z+UvtLpKrDJ2SpB0a9S2riADSa6+OOyuidttoHfvnm0mm
iywsUDvkibZt5Y54H5sr0uyJfZhBFRPFhx7FkvUt42vkxhmLXvCvTsnPbHFXpkcK
fOq7D9WUTdYFhQzZdV5hp/TmE3hAA0ObZkuqeMoGah+Wtpdnbib5ANQft6xq8ve9
uxGUJL+6RodwG7E5EE67I+ZfYZUm+URTvU/rkTTCno5ZksLFnPkCbPLhmLx8WQBv
dpOIHKg/K+bUWfelP24aQLCa4akND3nGa/Nrg1g15xx6z31TOHgGA1tTHCw+VMlT
NE2+j4l/p0yVYxYjCkHHKfKiEXt3+Kjp9vTIO8W2CT42Ree4cnjsKNUcZsMQXiqm
Y3B9mddIrViKc75wnPSPm5P5JUpQviSO7IzHCYarnV/RU4DOlYZKx7kGx36dQdAi
I4RTCpfzyQToNEIBLTI6xzfz5z+lznWQUnXhOGIxvgz4NRAa4d8vF51JNrDHLPtZ
C6N5Gkzjpqm+8r5hPKPFXcjqpHnfmpPsTq2uE5QHSG4TwS6f4Hwxadm5RybwzQy5
8b6nM4ho2enzbYv2lTzf4jnIoE6UnnFqE1mqmKooyqTgGxyogrsgny4ObFc1q2ss
IM40sjYlvddaAk3IAlhhP2DXlkJ0oFlN8+r+8A0YNU+X9bVH2hv0Or9ItyUR2xSa
z7gJ1HFBA2Nb8tZRuX/W8mUTCNTiIUKQzEb/CDnstipnw3++uskbG3xkBIZEYBkL
A5YT2NWw8ygGseHUXFYFhrie90Mw94lbMRohH1u/CKxLCNIoWqZAexRl1AeX316X
+C6k3jtAP8B7LqY5Oo3Rd2F3P+AE2HKRR7FYKLEnsRGVW8TFPlx9NSzsg7Ssj663
Yb83GEgwpA/5DjXCL/AI5zztV+7lFIKCX81bIvLmlDZMOkCQ/7pxkmVadJRz0fH/
fwbif24zxAVOvH1R/FqmBrmYa+wSR0jUqE3UAieNBvtG0/AeZM0mTRvmyw7o3xin
wlmboG57I2udgnQIx2CT8h1U+QVjxqpmFWtQCwBTj9F6OVRn5RDFNUMa/Q5bb5u3
7dQA9GggO3PzFJpsBkT669c4aYGGiFPmMVJ5IhXqt+HM77RcINypVbjkwzYc9DYC
C2nEEWJ8xtRPh5BSTJa1Lpj2J+U2oJrAJwuGBykiOcOj3mW35I9IcjKE4EIt1qCA
Q60MW/Jd4RoQCpM/9dCbQtqWdAahEVvCipRQjVXR8qkgz5yGVWddLY+p6/n3DQoj
alhX4oloeIW8hBBtiz45vk80jjUYnkloF4QrACFyXFELedMDx6M9Kxy5deuzfElL
j7BatmHt8tHwgnA7K/SZiscimQoQuoOBJtUTqRUl6KYP/Apse3jTU63JOBP4Tdbo
ntX9o9Q+7HM6pyBTZdTIpa7IbafuylvTrtn3/eOnYVAnKen2m8skZP5uPds1tfDi
HZngV+2UWtd4fgt3ygEoDVvLejUHtjuas3wPwnKC+388sJUlI0x4A58FaZ77Sbi5
heiuVmeRnnUA7FekUi2onG/sKdg0V6gfUInGXqbSrcWOL6ypAiya9K7sIzU2/95m
aVsYZVYEwghXe5M7PO4tUN/uQs4j62GjaC7oESUP+Y/s5qbI3ltU1VTylmHrLaH+
YGJV1D4SFqxPLuUuAtaLtHvVt5RYMkm5+0oZr+U5jyre8nIy1T8JEuttG5smmWHj
/WIxRL2gw/vYifoT+rF38Q9KkEMjUzF8aU/GbgNwaUZ5aDRYObwF6kwnZSV29MDd
9zVn2z0BAoYO7jVo8JlQLyPulX72OF154wghby9IPTxCf3D2SbHzljx7MYnIMRVk
hKpTqRMw4/FGoW/AUyvHUyEIEQnQGmowQpn7hGH4ZHVbN+jqBqHV06KyFC5lL16y
O8lLjvD0oeoxtVzhrl06Ut4MnQO0P9PScEQ+Z17gXthTRXmJAUZ6eC2CWgW7XQih
2BrhMxSMk7Gfljkb/EJV1UXFBHdgt/gwxcHJjsmw3FYHCRQgytTKKNHhMu4qaazC
IdZRhpXJ71jtmwTSwjCQPy/T5kpBPp3Kz7Rk1EphB510q3iPwHHRv31InDmjdi8K
U3SQFvNCsHW55Kw2UPukwr3Ji4eFefsPtGkigR47TS9RQXnSVivNjS3FHFypHvBp
8hXWPanyKyvi2qlaqhWslmSo08gJMHH0rJ8/+BDPM5TGMLnF1wriNJzZv92jE5ME
FGt9pYIPsbdMm7gBPGHbF+1YuoRqZhl18cxFw1HeEH91Y0OrJXYVr92FBKdDzyx0
yTbm8HE3RswvTLjv33XbLqTmtTZr08IzwuWyOxd/D+wNyvJ5pGStOc+fpvEHgleY
RZeIUuGjYV5b22/RAIuXr+WGmAkaDGPbCEFb5shT99I4VgDW+r2ui9BiCrEwofiX
v3GCh27ARy1PN45NvWpZjVPF3hEVxTQwAG10p97Afsud0Hye4NMdERMx77/8AerX
kLFUiJTiX/NLkJO281by2fg/qB7NSgIXgwlnSnJe9L1LiNXSDR1aUMyXR7NbZiKW
CuQf3cwejxzm7euJHJAAPzfZ/7oN8WO6wMBbDRbPDW2bxP4x1uq3eAUOPSw2bphS
JZM2ww/lHYPvEUBBNyJMIQ9NeSJWnHXun5/BuMFfOB0A3MljMh/wtNazV9IQHzB+
23y4IQ90xfr6PwT+JuTDiljg+KMMas3AthUIQs++nK8JHHL7Dypy+zmD9ECDPGJo
GcMG8RluXRUtbqCKY6cUdM3txeuzfollddQadEO8pipImXZGywpAQTwU0Oow64NY
Id8hWWImdGzPTetoapnOHtjjt0TNyv48SdXiCC5xsMio9P1upmABCGeiO4MWK7ZU
zmnvBmKiy7cFN4U1U8+gAQEieLKbwcDF6XX4bGKAgVhNq/FQLBOtZ6W5y8zgxhws
zM+st/cK8EFiT74HqWa8jGZiWcxwDH4KBO5HbBltNhP8Z9FDgGEL1vzd9nd71mMi
uJ861BKqhlAlMq1g17osBdPXJ0MyWsEmjc08P3h2pR5i2WiK7IUe3q1qW95i0Vbd
z6W50KxY47mCqhX5XmaHP+R60NuQrtwPs+zdXACkBkN/yYVEEiT2DG3i4SNJGfnY
XWQj7++lA6ZXr2KQ7wGVvaBMxtNB0LSiDrdzjIiOKlauLasFHZ5hAip/onN09vjA
94n98qj4bGi7xHeeGUU3OoJhC6mIaiuEFt3bPTNaPcFI/3fPTm4huH7gBHQlHVxZ
DpqEmiKu+fuU6N97ynSmvtGwAXNNWPkjVIcbQssX0LLlsK8m4GnIHIL6NXsdf+Ik
twsY3x5tM8MmroY8trrB53wBnYcTx/6OJPeCoGi/WrWU8RAsnOLgXNf17SpEzYNN
LNBhhRQ0RIFdqDTf4kxbgn+C+rEtnvkS3+IuvpKa5OuBV3Zgn2cmfghdQyLZ+YJc
vmS4LcgAkkcAjlktmzQajgaB+buctLfCf3SLOpck1YD9zCxEPkk2qWJXA8OSx5k9
qlcifjRIkGFo/nnvXsYEwwKmHnyzqRsT2DjZlG4zKtsb9yZHptQ42x2ZcL9HbuS5
Pn/GTtPPf+gpznEqH0+zwiPcRDTzF+UYkypJTJzav5Uby+OJ+qjzC7o7OP/dBK8Y
G2LRNMGzpHcd7mIUrHgaV73GCCS+SeNDg+Aj+zhGFb0AXytNo7dlAMDMSWWQGrN5
dkeJsEWRIgu5p2mSAnDKfrAZj4WwlQbKACzRH9Goco41bSo6o0ZqlTsC+E5tG+lf
BZiXHzGNEjWLVvDnb2J/RDkXlfBd2I7kkBr554dZUrDQZYAA7/ff4gqhvMSGc9jD
VtMEpPhEJCCBybEcuFN/ODAiVdUsD/JOXOmaLySlqyI/ZKJFfZGgNrxcuivsBFEz
+j0tCCI1oI5NDOumtgZgtlvzqs3I7BEQgg/WbtN3utXBZ4pXWGqirt45Ck4TYPLx
CjI/krBWQv/FblwrmKTOrVuoICwlzFSb8rXwVW57WL0/k1gMWoV8zoyi+j3E551l
dU5yqcml3RTrSDCljgOoe0NAWiywCf+cpPHXWYmCVK6wxabPywA2eaXA9Kc1EV/Q
Yh2JsIBLv54mFN46L+ysHJRBj3yU9hFw8W1R/+HHviBj1WkDskvqkCGNZX+/ra1q
HJFPVmTdfHqphFKcxEpHA1nnWMmr8Qd0fB51iVhCo3CQzo1z3/YlUjQszSIWhh4Y
IDAaEIc4PY2A02iTwZLuC+VtjOXz3o48zzwjRehKX8lkY9db7RT0ti2cMYiHKSKr
A9rprxAGau07tcpH1v/uKGGez7NoMgKrBFt29nwLlVQvV14bOBzn3nimXTVS7GCD
9NTmeAYlBM6HxEeh9PNS2eX7vOey/+EoRfV5LqlJNJtUzT62r/M97pCqCfwOdpk2
c+JqNxeVHRyxzX3XCMdg9pJsXhxya+Irr92RVwawSb9m3T5mpTmrevU/2ZpLAdWN
rLePFThjMOUvkV2/rGV1guqpUfO2IkU0wyqccGAQpnL0NlsWbat5c/lqWJWl14lF
GqpH2BYmFf3VgLHJfGKx97CaalqAqEKb8w/Km2X+zK46ofu1j2EU/5Lzdd0y7b43
Zzhy+5TtwNWHoe76Pm//kxEaagPXPq9ixmQVyjjeKAulJZuKKbl3iWDNyfSA0Cht
L82I4JhMSEok4tDeWKcw0fuwPSr911qauO0auLFw3HOF7JUQ843jDzHu0x2WeadA
PCW+jHCn472bT3PmLoXVtvEa4HWSqNqga/dBtIBHX+4U8tcvABAd5Ird+3vtNBfn
Xo/gslMW2XAEEizO7SBnq+JyQmNUM768NJx5tWd846EmVPytX8Dobs2GjAdAKh9g
cnIr/erVotMFuV62bSjmve7nmDMH+3wHgkxIVJOYvgaZv9DaVuJKEFPr58/bTcPN
DCZHH5lJy42pnB6GAnNBD6Jyp/o3MlEG2IPXB3yn9PjvqDp0YyZVLljdYaGsXbav
mMAJtvEs9UiqYka37S0DkKUxqsg5bXv0WmlZCsgG7yBa4TeatW4iph9kJjbaja1Q
/b6jbDBeyUm4zeT+UPsaPsYIZ45FXo8TbUIeXhGzAVojEbQfpr68GGS8xDcTQg3D
83M1EQC23joD6tKCA63R3STrK5ZflpRoYxk+PDC8Sjhf2mTtfemF6VM9XZOsMAa7
y/GpFbQDKriM1Ppz4osDvB4FryGTs0m5grcocegBsUSWuYLP3oZjnfiOCSWn9pkO
OjgUfPEoTKSILWYusjDhPWcUGtb83660swfmS1XyGbc3mqs8U4RegV9K3QcAYWV1
S/uNjc2jQYmDKZ1vdqPMP9wdCVoyYwXudA6xRnfP5fHpJBr09xemNgWRv+8y0e5O
foC7Gk9ubWFb8cygPBF8RtL/Ah4zztrG8mmpK8q4gUT3cSTYBWIDrMaT3zjPeeir
B3BYuMzHtJhmnK09JKUUO1OOhgeXETENmu93HsIsyvmXZMdvAev6Adna+bQ4z5q2
w9mu+Eo0itY12CWQYWoUv7YAVNmxxzejxIg9+Kbk+bVXW0l999OioqawFMUn11Rf
SDdcsazW8pWvNq0SOTAyyfJHaOvUeycnnLXI4MUrCkuMEOaozcLgSi2GORpa4q6+
FWU1TTCG8H6eqnYsLLkgTg3kED5N4D4nGA3PmK8Q/+y/jZwbKDatDDuxtpdnSkPR
vbZK1nlo830zELePBKg9sTpwV/HFHLGfJtNTy6gAHVcc8lH1KK5p5jk8tSRBhETe
CS7ckNkuQyKSkJKSJKOqmoYHG2pYlOcOyPLo3D29rJlAQPrnmd33/1LG4SoA1yC/
CgiNvpMUSZYUh9sMqMdZnuQDuVGpdkqAznMA0/qg8HCO35cUvk8IJm3XdrVk23wH
kUAx0305B6hYc9+IQPLQL5lqYJED0W312AsSbFM0xNz1HHI4QaWKLjVMnsWjYHFQ
IYIpOIeMbiwjloUVLztOlEXyra7w4Z1zUVMPjbpE1MDAp1Cti146SPT2MdXr88WN
j2BmvuIGAj9rx06qixeyoV1Fq7527Qz/gTEJLuW7pML4Shxo6QIJ44cULmg/5iqs
btXlRU4/5VqMryZG+Asb5JVMSjF/nchG7tt8mzYDBdBn81yv+QvhRxArsLXyoJyO
Ab2GOjWIARLybQtGn+xUwdIub0pakZlNJ9jH0S7L7UMm8pSdYW5ERJVI7o8+6WRY
01CRXlbodufi+0advswb4EoTFBi/vXeMGvxn0D6AkGcI0SDw/JvWILlWX6EZIx94
i8brCxH7Dp3ivaKTQ9mLilh1dMppRBuqahLF2pa4idNdDMAk73FbyeTUy05gWiXd
KuqiCT0sBxCHgVOf74in/toky/unWcT+Jhdhefn7Ohf9VWOfF96/7WSVZysnJqrp
gaSWCRe4b1xVbflN/vH8cu7olHu063LqlY0kv2HVKunsHMwjBuLn+SvnQduEWGZz
Fn31YfcX5eXxGuDlGnE/BA2JkQgLr584qVCm6BoVLHGoub3L7pMNL5mXAhJssz6x
iltjcg1Eeye+CxcFPMeJyWwEdxO+D48kBLP+psYBhzI3g58ilM2nrHyKX1KXcI20
Pe6Fy71Nmy4IPgM865PweTH762qMGMukmqOsdIMgNJo3ShC8ObaQn8CsF+21pkFm
L2NMceWC/0ROpCOFKumrS/bfKX8tMByHthR41POD0JDW3v+eT8bb6yu2w3VqQXAa
Uu41vT/Aun4fE2M5wwCMdwkW9bAc0xsTPppEiFM28HZv0QkrEI+0BEPWrxKEpsNW
DD33tldZMUCRSL83dWaMxp7QgG71K599rTEo9xTd1Lp3WmwZgqNZto58JQ7+3XP/
ngxfLR9a/bddTdK0qldYYXgG4QcieoAVTcTitIF7ytJmtb67LpOL3PLJJWYFraxB
I9SvtnsUV5NY052QGaqX8HXAijGb5nyp4kTYE2FQNDoseA3aM4yJYuGgxNYp20R4
J5z6b/4M6Jncg272w7nBm6Bajlca/a+kbqUfQ3SGXyL99jUNmEGGgDq1DYSoP4jF
sGiN8qnYNebyRWSPRxx9POiwCAmmKN/1ObPbGqWi9t66IkYx7JRcceBzeqNtsllJ
i5DAZ+pVsPM6vbVGrzCTPvLFfCeob93OBXji5EFWvyLFRv2k3KaYSDnDYaBxY890
mgjbfpgSzxFwtayxNsNA9rY1MwiZ+PuG1HI7+1l104HMubjB9FMr/wkgUgQRyNPQ
3MyI2nGV+tVIq1GHjqqUyHS6Au740a6d5L9Jh/cEJsAluZjCR5IDu2WSX59hzBf8
yeheEbOYisTCXqLPXy1YWwjp35LclNr6xbryTTEjNdIuzkqhtHOFHYlJahTyGlKZ
/FjSqtwWDvCoMnrUhqEvXQwq2N1UHTWcDMGHrwD99p7KpScPVCTBVrpkF8NYjl84
HW3AermaDM0iQH9DvWt6wV9v4LcgyKhgv/cH+SenAJPYsDoRp2Hyx/Slw5FnUN3K
bcWGQKSCnao3gV3Y6GdV6mHu3sTpCOZMBrbiD+p8MyFUio8vyd1Xa8nI3cBRU1sp
Oc2gzO+yA6JgM2lS450PwgglwcHnuX+7VeuaHUeODcyf8L2FdgIiRX8JzZk7uW0w
lpwcOM+hjuZnQA1CxsxILvq54WAAwAHtmqnO3CN1m92RuG3m7nx28sHVAPMxBTTk
kPhTXbLFXINEvSYsfIeCJfp/8zwLwaVsjr9HqpUMsZIUMcjU0j4Fu7NYR/d4NRNC
aX50e9gTAiUPet7FcEcoZmUCSawwcPUMrWsbm+u0bf9xomg12pCorXfmyiWN6cVL
MYsbaQLpK4vmA77nWwdnyiV6BZo2jxNkl2JKL/4UjFdW6Phj7w01aVNZ731vWQCh
ZRVNe3xCmuBUJUE+B4w+WjaRiyqBR07EZ0diAlxNFhQ0BaGBJbAIWu+3bsVJeONb
iGeTsyV/SU75oCBcam20WoWHlK3s7pkywmxQpViHS1k8XsIAflMi/gK/WI6+VPKT
Soj7MNzaJQOyW+4I1Pe4En1lQPaOYgWCBlkvbf1ZOebFgwd65wibs8ynXyYAa0rc
Kr0YsEboPKdho8aa+fsUgy5O19bULDaOlXcXKLa3Ce78q5Ov+J4S8SKsmy3Nz5tu
g9rv9BwAySwjwoTs99se3w2pUl55avj11SvBd7mMWK/GqHmu2o3iSc6K3Toa97wT
inzKME5BTQoQGLRyKuLqleoPYKpJiwYxxNJ3bQVGXvoss37Gh3vcsgb43vEoBi1k
kemsHsLM2nhcGXQkPlps9HMTRh0672E656g6ojAU4K5dmdWwOh75517RPuIv7HoQ
R2//7t3TAyQch3mGnCmzg0pB3V67SGyVRlnF8m4KHAeE45Ov6NXwDe/fh13S7b3z
AQflxg+FqjmE/kWeV6vkkVJ/dVzv2N3MWZ1XGV4sjOzyDKnihid7tFxmT76FOOwj
JYo2yYiYce7ZHWLWcSLCde5iuUf34SsXMaMrmYIjQdpC7nWzefZKJc5yxa+QC4tL
WEXtbmOs5E0qljBgawJbj/BMucsPpq3GllKIRoG+NRJef/T45/bn4bwRMey2vORn
RR7PwvUjY2dIe3/dE97KtAfRFWqEWY4m36NGCdY0HzOnzIeAZuUzYEZRLiV1mUJx
tdwEu1vor0+eTOMnbAh5UXYjyUg9OjrMY/m2LvOHSf52JYcTxb9m5AthG5U9PGDx
7Sl7lwxHobuYYj1EhrFQUe6CTnpfJLMpO86Fn5t0VE82PIj6TGzcQ4TYlVF6T+LH
gpbkA0cHiptawLJ5f4S3VrqyVhNvepnRAvnRrYixCJBOZSl7aiO6X78o7o7zeOo3
z3nNXrtisv9z/kNEuAqHuUm2xmBq+gQnqTwEJeMYRb0GpLUxl4wyBeWeH3fjnSEo
dT85tBHnLpWE11JxN3Me0nDDKybkfavhpaWSVxjA6bffBS++yvBh2zSHdxQMlHRi
SUdteVwCntO1jmuDSqs7t7Myrm7xvyATEuF1NJC2Iu/FRmkYkZCNWf3sFf7qoGfe
80NEYx2YSIvkVnfzg3eFSKf1xaX2wOJMlD9CM1dFQRJkksp2P4EIA+VsUtyyF6yx
166CxXQms/krApEaUr9kCuGHEl++I1+x/friUpMx/S16PARcf80w53DToZZFB8a7
J6a0swC0dfUkbyyG5gyF6J3j5ePdG4re/Rcz4XBH0S4Ea86JwoW3SEi3u3xZYSkz
iK2mxsjn5BPLybJf7W1g86GvGx1GU+qXDxqnTbrOpWlWBgtfTkU/n5LNXOQuZZm+
dkrCsSYkLwVfpgWpaAxPqRNUuPSCNd8WzBuAy76z1J6WL+/q3WNoBmhuY3NT2+8g
DtIgl1mo9sYmgULH1uNvhCDkVT0Pn5V8hQxi97i/t1SQKMmBQWoPIknDN+QsRLBY
a3c0h267y7if8JlXCZOw4oiCpiwzYzU6r39vapHaIF63/bVhdpGsAIsxR/1d6g/k
QyaMarmdjktBg94MEtssZU+HmMYYXZgnuZ514jM0wHQULbS3mr5oMVBrXMRhUjPE
ON6Wcs8renY3uS9HCinKvRVXypmd34TcuzRyYIz2kaVwFqUeqQj2ZO85NHY4OH6y
L7Ny0b5DAxcW9lfgNuAHfXjFqx1pOqkyUSk3zTUWdwdugKafbHKPhlej09CVs/4V
oA73Vva8kB706wrgiuNry9dCQWMmuCTgAZrCzmfe/W0DTLNcBr4HEY05VQTLs/9a
4DH/4Ll3oJAfPVbDibJUrtNf2LfgOESALvrJ2jGqvPZluFe5OH1gWkp1qTgmPM1b
P5+hFn1Fp4E8OyInzFp2p4s2CEdkLS+63iQvUpCx+VH6ZVb674IcGuxbygpzhRC8
CbCZOD/2Wz9JYyy79yGCIM8duSaMzGSODZ9alhEQ6Mk2bbGSHZC/An2QRjUIXyA9
iJdi5oljMBlGFE1yHax/gz2CooNxJLq43Q/MHb5GsXy4CCksIcWXuaoAGdSV0o+f
At9Q/tJH2h3/Kl6xDK4ZtdE26csN/knGO9dZH4qeJELnmLbK6ULCpmOui/tEpYGd
xc9K5omZ4cHVPba2SAzEjL4+5Zgcp3KWmWi+WGUh61eHFIgi58BAY+PXKN3+8PD6
FmaduKJtoXL0DRaSqsWX0+wcmwIm4u3vi+Lmn2mweaEfpXobjcILkKEwdBlRw56N
QaAKUa9FuWch0JhKp8j9shpVDpCWmZ8ZWFrdn7K6rrdQ50E9aaba5PjKDNA05X7A
Q3Am3bwPrMPLF4v9d8fvSWCOLBXuCei7LSnA4LFgf4hCIXFlAPF52O7F0tvlpetz
PVIjRqxzAnEGr8WMBnsEpUjU87l9e5SxMHchS1iFlRdsziyJcA8JeLrC8uT/N3MN
ydpYKV2APalY0zCXVIbUmfRK62Nkq1vz06qVkv0amTqOoCE5AfXU3WRtUXQGxw1D
G58/W2LAE33AQotziPdJ8FYmT8y1NgGZYWuppK4z4wNGWBuS41Blkjey7nMFiSwt
w5qBlTOnd/jpwbmPliRS+wo5nsI+9A0g8Ttm1ssuWlqEnOlhicYdFW+H2wKrCErO
NsVXcICbL+MxJUuqnHQVV4aLUhgbQteldxNmy7U+TMG40duDMiydbEk0ANczqA4P
uNR+vH/NdLSzEb5DXzHAYJSgnBFn9oaKPPyJt1zEimn7z1Ku+lh2+r5xBhD/spFT
zy54h1BUJ4RWeppszcEpnvgLzAt5WbwyNfSdo9JDIHBCD6B1+ukB/b3PQo+oyZp4
bk7qSFzLN6ncbIkvriO8ulRHpjw81E7yvFB2KgPVmRFvfB8T8A67u3j0gvyyoB7x
yfKANqLQwjqBJsSkZ4CblriwvukMmjG0WqMXazh1yqyGNTR0fC8WOzW2c2THu3uI
gVRVO978zaHpigeL95iJaVrwHqkNN9XtmQxxUMV1++8wBqkjW1TUbRz9PAJ10JTw
NJhBymimL0Ce18BK0XA/DxZsm5I94jDZjLG3ALYNmAE/zociXXL+yFofxB2YxLz7
O+8OilspiLJcCh9+CZBBgmkMjp0SlEftaMHv9opD8Adgne2fO0WCefMIGQXrxI3t
jhHoSQUkI0KsyL+WQdOAPmLfBmFJ4F9PSMwwD7eYdf8+U/GZI7pOBuJ5A53E5X6C
UYxwKlvZENsIAVw3CJtiGkfsoTcGoTYcf/3lVw8aJdcgMPfLmtp/lZPM1CY9HBmi
xRQW8GnWZN8hAcxKsNHE3u790zsQIJ6XVLj3UYA47JPi4wFael41V1sBKPi5qC8G
HxFeAVvDcxfbD2eTilEYCeyrYOeblE23Rc/UPMY1HqADXJF7P+E1Uh2ylEL0GymU
ftIJ5atEdehAdo3JixoV34xcZZ6t+EthhPqEVI18jIngQRq/3ZSv+SqcsNMutpHZ
EZ0f792CFdg22StLqnKXhj/BCrHG9wFWI522mceNSmZecWtwHTy95puu+HQxKuJy
G6wPrj96VCOftk1Tx17MEawlvbzgF8BGTt17zs8SKFlAsoJkwpM3jDnWkkscGNUe
7M1BOKBCtAQjR6UQMX+8NMayrRtawZ0u2Re9gEn9LCa3mNeeVkL5TGpp3sPufMGC
7GGR+N90diLifyvp1EplWbjV4minqNMURvPjuo5qvYcgPySrlTyyY/fJMnJHZYrO
pfiVyh629STq8vyhDJwMZxRabzkbcCNzU6D225PNDu1LRsoBVJjahS9nqPT+nFDg
QH2fhgScexwEr3J+J19zrljTDhyIy99iBtr1dckwvZtzK9GEt8wNEBlbNJWaSC4n
2jIGuCpgux1R0o+7q4q2KX5MEDqgb2a7JVUSpiqDdKN5F0eyACNgVDbKnEOH6aEU
vRVrC+OnRdc9022N+VrQdeQosHUHHs7PHcBSExtcDxgaASQww0b7fM048GldJvZX
NKv4RvkQbXMS7c81qGJTIJMpEc25w5BX5T3mH3OjxfDJSs6U5bDkqByerZR591UB
WKbXZyatzaGAysK4/dn074W5NrsJnDVv5qzIVW2YogIFhWoroWFnY3uxi8cREkNa
10OpSYy6iitp3qwjmCpxu6S7oqGjf8tVgTAhdDsEpCE/7n+rSpKdRVTX0b2FsMF4
3z7Tsv/a6rrFZUifiTHnMtFwaa+54Y2dy/mZAU6n4TQVRkpOaXiLzfcqtPYWl5xp
Q0bZrG4FrG6by6g9AwoOXLZdV0gXJsj/u9VZsFGK3BcfhdeNCGyUVsIYwYMGRk/l
qilIsj+XlgVV0d1B7BCqsehUCpt9XhHDQwMko5K2702ADKqeuKe9k3WZd16wMzPF
SXvMiIGzyUr9O/N7ZamCl3w9eQ64vHCdsU6+iDAA7O1ziO12WYizRHucdLxAW1E1
UL3oPRqT2YzGj74ZVbE3xyVfT4pLbZRkwtcfqKGR6E2mQygcWWPyQncq3m6HYV8N
HceoUk1tlKtKN8OniVNzd9T+OWkp+FrHNI+weJHlnT4q8tNjoYc+1OwpIcT4jczV
JFMIOhErzSiWKBiWNfyspTSCXhpeiWLWxfEe7KZdMqkV2h9/sOzjsLZVKRZgzJYP
GYur7klOJVecbp2e1OyQ0bj0L3JF1kA72Jo16abFL5bWLTld89P+DBe70N3pVDBN
fZLNBpY777w++6rS6aClns9pgh5DpWPQ6u09fmHRiXKZn6mLfBSMIjKKUJC9L/Pl
orMGBD6S5DnjZzYs3iL4gz2MJJVdvNk2zh/1sRj6CQdlQIuYG0NGRFC7rqoOs2jl
H1xCtsxNLbEcPBOez8UCiG/H3BShnwbcvpjFxwD0hGr5ZYaIr04k3UZMHJn2/8PI
0MI6gwgFaRoKkGxewDEXQMGwA6qfk6YGfNJbIsiKaAsaL9wur2iMXa31O+4Sfls6
q9qVHb5vM+BZ+Wopzkx2bGsEgwV5frTgBCqzPxSvtQCIw8O9bhFrBzKAgHUngcxd
NJK+uzjLGxwXPKhRap6zi/MAEp3fcbFuff7O9VsCET6aIQFine7plsHO4XaX0sIF
4uxcQ8mAf1175Scm0WhkWA2q9orLITkZOXFaUrSi1SYwdLiK4tP+Hmzue8nb8l4W
KiwNccw+nXq0AsP7L2qBsATFlOXfE0ndhMluC4xHYqxl4j/cLeHauSQsx9fUFLQp
Ew71ZQS2esUREC9gsdQaxn5k8HOxVD3Tv+HAoR6oZ5iFTp5pYAOkUm8rP/BuQO9S
vI3ovw1e3zp4MoxDrJ1upwc1hjCNgckl+7895C5lcKIeT0CVhucMigmiyrZc4c8M
jNGFp3hKN9W4+osJl58Czfv6PnKPy9RMQng9tqFXCnyzIKinNPquknkrqm9DBUo3
pl0sOiG2xftVHkkPBjmYtN7pkZqOiaE9AUI5QS/SMolgH641uA7sbEAR6mtBY42s
1kozphAk9wXXouHaycM/jRYCweMH3DnHRN9s5KKezk8mKIG4elpBcfZeUPEGtPnQ
hzLI7va+k6+fxaZUk5iuSH6kNLqvkk2jit9zyoFJ0EbF1m7x0tWxH/qsu7wDGyGt
2Gu9C1uhK82WxrDbTKc9BoFkUE31bGgWy2LcN/Exau72ZTyXW/tN6mwdjXQ+03VX
j0MtMS8eix+CZi0yIHtZ0RY5chOadhvgCJrkG1owEXPLlvf1w+N7uxhPwNVxdtPU
7cRjdQIV+Bdi04rWlG+b+hQH2s/qBslgZFtm/5KCh+dBp4G2atrCqfiFCTHypDkw
9r4tJ9QXIDs/G7s8Hg/gMRebZan5dOmGj/lZxGhEVWW/xbvFh9k9UG7ew/f5+bZC
6HSAXyVDyJQEAk4i6rLH658sp06HGVS0c4wfonqgmLaoTw9x13TjmHcEZspTtph1
qPrwLyl5Lz+EUqJCF5uPvCRIryHrYGKx7vTV3rt0bTSvZUqScqj9rdfhTz+1XGLL
tNxExrVecopzbk/PxH/auxO5IZSWa05awN2+jg9p8U3KDR/fymg3RI5yRGcRmdsx
kzjXTuAXGmmPBh28AB3WgazES0U1fFz8JSRCZ7CuuFh5ENukGnZcWEfU7SL7wYVh
KLDZ4TZDU26veymjAf2h3qlDFYp4ZbpwMwwlSJaVC43MTKNy8/P7jcq3KGYLqsIB
kMKk4oucdxMCTZ2BGDZZlkhD3pYPmKM5G2Ltrv28MY6zJHLhH36gMbysy6m7iS8u
HVSaQxliZlC9dFK9VqF7PWAILE/G4A8MQUMVyKnbxWLU5LOqj20dfKlLTXSia3xR
cKFVgC2pEd16LSkhuuuaIFdqR1Of8NRm9dlHMK4Qk+NyTDGmr8jPBfigozXVY6SP
+LE21fM7zht/T5sFxWYaoUfbi4T672sFHF1logvTWg6KIZtqJHLG7Fgi7Xunovio
6ikzoiEz/ApAiRECE0bXalYCt049BfonCD3atZnXWxh/+/DUfyDCUeFuxK9+ItB4
2xJ8GM43IFcjuvoFIk/N0UsQ7kPTlMiEomx/KDKV5+TfsccYrl8F92ChFRIVZR20
4HRfzL2Mc2XvH/ynq/4/fecAciMGXTQPiXIwbBa1VDjhV2LqE0wMDuRTr1TrjgyI
KI0PbAJ/ebPGh0zGJHJFns9O3KohxhA6cn/zuTJu/pceqdY3Uc0mhEQeUR4Wr9xp
zI0C78ykGqDWQKEr1Ss78WCOZunPxmAMavgj13ObxcMBpOfsqCvkiQTX71wUOmqH
lxNJqtsxRYhpbyDYByFMx12PmPgNDwChbNFDnSF36mFPiqfov2A+don6fhKnK0Td
Wiggik9JlPPA/I/QBIlg/xO4yiA9io12S4LsBWbOJbjWlpMgdb4q7cIdodxqJd52
pRqs4VhP22PIrdcLhTcFma06OzN9FBUDNLg7aTCrni7fXr3iM/27YXmhHr4CuRfX
bRb6P4RF+lVdDgJvPW7GwhsHnoH1M7Mvv79jGetlncJInduOBEcsUod7fu/D83Xc
F72Wm6BUExwxGrE7Asy/AKxuneaIJxIckI9S/brPed/iHP1YzODdfybLIv165b1D
Brr0IsFqP8n6s+h7v/x2h31SVDdYBCO3dyELo80tPXGj8tTiaNm3uhjcBU1zUNhT
6ntu3n3erCi/48wUxosDgDwwZVBN2BA94hwXrYQuS0Z2Q/CGL2a401jRMVXr5qQf
MKIi4/YsT/ueQlpTUPONGg/682BZD3Br7/Q3eb6vGmlDjWocwf4mOPL1Adz41Lpm
ya1HI9amvL4D1Ag3Yr2KTCtSEcjCNHKDt8Pq1oZwii0pHce7M/tCxQhUMAtyHg2S
SSrS9uuubneYqe0wnU90w845GJni9QeK0fGD5MhxtltpnWJrwin5BMm+U5wJeDgM
YFf8dtjzE4z2DNz0qVN9G16GCtS7XVhXwMebC2c5rLfo6YQCaGINXT+/3ymoAbiH
DJ73HTTwjSYg1wVzTocKCcErTmoj2Q2brNQbSFcLy8sa3bGR6j84H0ko/fsHHFZq
2BSudMKHZQVRiSKKMGrNIx7SQMpdIJVwjkuaWZZXXX3UgqBuZIJ+/kVVXntvXdq7
RGCWFO1DFd8uWkJkOK1A12wvT8dxXedPa1WyyAFG9L+TriD0Jd00AgdUZ2IjXuYC
PvTPI+11p+rNTt4FBklxT+FcLT7QoukQT/oGE8epM4iF9VWdr8hTtlvQ1PCRLOYm
aE8VwGv3FJ0S+MPgm25b0QI+h7tVyxpPfjomeNL0+WonroljKsihdpW1LkmzYNFC
9FwfMT7Cftqrqs3BrOw5FL2cXX1kEzwkuOqqRFO3x0vPhnTYnRguFkvUKRryISF1
l0Uj2ej05RnWnf8OEOnJU+xQKa+EGrdT81fXvJbmnMjtUQ5zioiBS6YjPvPH/M13
uHOQfkt7iPpS4t8RM5Kpj2HtSTQ40tA1RtqvvutEWCxtyqyurW1zyfyNqjkYaQmw
57NiLAcNnht7OnUbLbABPSTx0MXVSPwgVwj6CDhSiDJlw2bZ5dJXs1iogKMkqLoR
btnO/2CIJs1Xlloxnd/QGIP2zAWGlQI6oBw/76yFTGj3MzhcEbP4pu+LkxmVq/zK
l7rYKNrzbZh2V/sRCNbwgXdLsz0pzSr+VjkGMoWsQ+fywnrM6tULFWHfL9zvrzfu
foMk8kkS+UOhes8iQakJ60EGjwEga3k7lrW7horR59hAGJCNu0ILsZ/ZFlaluIPM
J+GhlCStTZhps+N5sWTtt13D42t+HCrQxbqShRkE2LL35Wy4X95fLIg+kSqi8Q82
7O1cmI/hAlGhUuAV6oQH6SrNe0AsEPpdXxM3sfstG1dV5938dfvgbCvkza0+mNR4
4zBlusA0I5AJ4sv+atbYt2+GkbewjonhCF34aprdKeqQ0opebBhXcrxi1FxFl3l3
xphaliI2/YDjDrBVje48OVJhTwCWNipRwqIeXSBC0VNUGy96NDAiZgiGUHLLtozX
HPBqvynwrLEWTpjwYmo2GaRy+Tv1wh4MazhGZ/y7V3szuvaDgrP/NZAc00e2DCQz
jBwFZ6A0w5KlTdwtgNraJxO+oXbna/AWHKW1dwN9n87uYLeas/nLD+c+RS2e2T5p
QtnCi13rI9BTzRnlVrF+tzOzLo5FGPu2M1+SkbvCQisyo2zKAf9RXJhvos1tfxez
8zVOEQ+9olrigtf96k4XGuaUx1IRZ7HSiU1n+tfoLuq7TEpNz6CnHvF1Dmq7nsyX
pkqTTb93c0JkIq/nrCfLawzTA8eL76aHBETPM2GG/x6pIypqGC3Eb7VFOSVPA35P
KY7KUhUp1cPlhBs0xyGCmktSzQWLPaevJ1MaSanH2EI1aL/11lfqbDFt+JW9nLG4
ZGwy86y8uxqM0a4hWTQ0v5fMQdKQi3liIn8akhxA4jNPF8fBO7HXI7E/5Xr+HBox
GTCXO6QiWiEdCAw0do9i9OcRTUhOlI03BJsi38ECPBWVY6m/9GoIi+j1cPMN0olb
PvqKeQwWvqsVgAIc1B2K0r3GggIQ9p4WOeYHGvP/Ef0Go7z0u8hlU4mUjuvXOFxf
98LyB8a8IzYfg4l0NnBIApN9luVgcYxW6Xalaox8aJxKgrzB6KP1aRD8FxxvsanO
Ly5s3Cr8NjXadSwXBzRvDiMlT0QRLlGmp9+uMJWJVJabzOEiQ7mhLmghRXro9ct7
CBYWXP67mR6brBqu5P85DYfyqTDzchyUx96LrYnexzk0K/V6/NI5npCmsHcYZpfo
soS1q5UH3fSpFP1M+Cc5DcFJSfW8tHoQAE1O2iR33gq5zhdIQzq+a4qsPWlkcFWn
zqK5Qn7dK89yRBdQ2RljbCgeGp0gQljlmTG2FOdpI3IMhdVhytujvZbJbnmX5Slo
7uIXLucNHDQLMBkkPxKYucpF3fRrCKddpInhv14+eFtNXmcSMhmZqMjBy3XI6rGh
oUSQjXlOc2NPZLRyl1bx15zik4br3tUeNC/V8NzNxWwtP0OTneW/2wdhBUUDnsTa
8V9kZKBY4UXpuKnr7J8f+VRGk3V8Golr2hSEdyN+IC6VZnyIJgA2LzLi9nXJ78qB
INw1uqQhqRsWtT5Pxy+LD/p14E5dAdNhbjE2+It8rguIDHwg9yBGUJ/0ltZsFOAd
csbTbxPCAYKC6u/sEk2vTlHaDBfgFd2FgS0rDPKf54eUAoFODYN/MuJV4CFG230Q
297LT7Wq3/ze7BDsbR8wJXYmF5vnrE6GpdnRW0sbwh7okNFAPImTSdRhbQSdtEuk
QHj1DCIo8ACCTv8QbAkfV3IT/uNy1ln1d/HwfwVhI/vPqu208/7RK7kUNlYkey/K
lLi1t8SE9aWbLpn1oU/G8Admuwe1PX8BPkt8lQ5uhQ9f68v0WF157MdYwGzOBuDR
UxqziWXE75QEFNXYBczmZwqpjHfg12LXi5gxJDXyJL4HKDJISeqlpNqK05NvSfiQ
k6wbKcnEeKHJzIR+NYNVmh2k4jYAySx+jOLbtEJqJv32GV2xJ0MgtXt4Kj8ocjNx
+5nNgUibhDQRMzS/f3BSngLb/KgU2gR4x7FLEMBBJpX40dL/VU5eNdRxPj5Ms03n
8238O1Sake6FsnlsLBt+cUL3/8WHjmVlw8teLg2VTV2S1NE4QEPi6jfavIA5MhiI
LzhMzTSqA/Re9YMoIzIC4ggfrdaafruPav3luPQPuUhk3v5whsAFmBts8vEM0Mgr
WffKFdk7WRif7qh19shYfDrchwHjXz4gJ5bvPVkdwICUjBz7uaFvrEv49ZLYgm/g
kMwtUNjeEn+hI6JmaW8J5SkRL5EckDEApQyswRl5ZiEy8uumjMYCPmaXNdjzgI4L
dvV8IIuZYWyIkkf+VGWcqcpExZQrnLXIsa3Am9DU4r+8WHmnvGESZVbuN69aKgRb
7XHQwgyWyZtJeOLaHmthtQBPj6LUuzK2ztd4WLlCHupHUtdkCz9p+Bu+/XBJQ6ZS
b3LmVXyd8bba8QS34wLXd4Jv0NdY9H7AgTVo/YVmtXFU0vDkFK65OMK7yRvdnBHS
mieiMQ6HWuF5JVYmD1N8JZeQY5RWGup24Ohjfo8UVgYSraJPlWm0m4CrY2LhQU2B
/iCnZkdLYg1Pkw6pPsS6Z0ZEkpnbazHXBWz/xHdGF9rbBLnhQBuIZUS268ZDhfit
tGTKt+bcFfmZk3RlEkaETtR0HsoA+oWJL11ABLQwgRqavlbG9R/uTpot/ISDWPvA
HFGUopluDYx4Dc0SJrYYa+KszdXXMkAcb+ZO+XEqfjkTK3CajJ7NiXbZCePTnmfs
Omtm01HNGaykE4fsqbFnDRiUa/iujFqBUy1i6XXOPo+ugyjuI/3sbdh33VEutUDZ
4z9qbTSLpJG3R40JUyJwL8n3DTkZDWTn6m8Bv/uIbFwQPXkMppmkjeg0g3r6D2YL
+q2+qSIOX5S2gBJVuZNrYf08OixznGftJ7Av8yi9cLMkIVhTMrHGCfrF7qCzF4za
NLOjtXDs98CyfIaL76baXdMU+EI6Otd5FZw8yDPSTGCgJnmBuUZDMip4P6tcIoBL
X+qoDx2vpATaKciMkTD7ITZ8FpJWRpOpDR7iivqArLAsC8tIP0v/9brMQOscWIhu
MbO+qfAQhojgJORv8tM3/QzfHOUMcvLn6l0kWAekGMDvznHRaWVgPNw5zIGNYhOg
brgp7LUqoFN7ipoW3XIv3izslTpL39Ar1B7GD76CnNUOPPgsCD17SbBbcEtilNHw
/6sO1VLMqYVmA5gFOtKcdX4zxnDlg1dS//wGlhfbfDC+5FdAjUgeFE7AtnvH/g1L
RZJrKPpCbV6nq3kldIj/LHQYa23CiyJiKKrrZI+uKT/qq639XbUaODSxHGMJtPF4
8QP/vppLKh32lyqGYk84DofxP1d38qQs/9hTD/KBUXk+8G1fRVieBbrSMLAw02tA
dVoGenzcPl6Kj8MuJf71iaLYXttir8pq3DxKTbcA9gL1eRtqlVkPnzTJuPiG+na2
wBsGgK2XJfsfF54VxjVFaYcTkyJJvFrGe0tnTlzOUvZCiSVCkZdrp5UKuxeNG1Oa
zdZEeMfDNWeNgSHukUc8GOOaQWxBbbKxwsX3+nl97FL6FL5ZiGYUiOhfo7hpdb1G
YEoXafi2T0S2k7VIP/GaR0lJr0HN8mHuPOXWu4+F7cM+Hq75jbWkU+4obwsAN/Pr
1+8G1ln+6gxv0XK2bpCQiAfovRfjeeLexQZArWRSHk1b9n8aPT7Z/dg9o/2wzHMJ
9/ZIqxTXLB0JCby4tGBWq9KfEXCQzRCpPP3iEbxuumn1Cpa3xjSyj+EgvDtAJdMD
F89/ncypkpCFX6jQgXsa1J29gv3nDSRF6wpAcS8jKFWpUuC14Zd4GGpFN6yzmAzS
boJf5lUIDx/lHweoXRT71QTW04AMHZsSrQEjF1TdZHHZkonR5HOdXGatWg4rYiPP
CHjJ2RjZAlLycLNSsMaXeLTw0SxU8/YjKBnk3aqLxwZkwXSNeAfZ1IwUhwmS2Dyk
71lGrEqzgryfg6DQDReGwqoWbwKuROcAdF65axMbb5cArWW2ory4KeLeFYcavOlk
BLSrk4xT62BPgknYGgkkFyksbxhZWnhxEO5JCyx5bpb2tyujKOoTV9/E/fSngPFY
+c3m/Ko+3qjbl9yH2CAXcpEE0VYofpJJXWK67UhItbWDXrPL3Ee2nmG6EEyCb8CT
52s9su1KAHUhJaU1KFmyyloxWf5fk/BP5rl2iVihpl6GRRn24DwjVQjAaP9+pL2T
2YD2l3CsD/vOlLDu9Rk8HU1e3EbgagBZ9hJasmDZ2j2ihf7J79sthE41syhHjJsW
y6DEkrwqGQaJwSMKAYpNwgVZpWOuoSaVqzOZ3AjK8ONcmfyMa0CPp2N+Van+dEci
RfK7ncackbV2oNPDI5sir7GEqqncJ06/j6Idva24m5K1UjuLu/aeKsi1FuC80mFp
CmmN/WXK4ILJUTOqDZipsa5n6nMw6RlYuijyHnyUOTPov4D5BvGg+UvcYkTnrAHu
7Ra9zj/+or5bbzc9mSWWM3oIJD5CzvbL5wxDKPqw3a7TxKqWyEsGmn/PKB3IRpDx
WgFpVmH7k/RRwjs4D3LZ2YL5DNCtoWx2ayqMj1PguKzU/4awWsDJsm4kU45msqPU
S5vpkIn+zrFd1BpRhC4t8agwa+xQNI16qc+0U1M9wptKurb9ORHcTA1oIHt36MKr
AZ+M+RGKU8D5Ph88qj8FoWUi6Qkpkym1VCVPV1/zRkT+jJLU4br+prQGwWoffnWt
Wkz6w3tlfPLFeJ10dkY0PKXALlUh5C+H8VL90lJqo6RCbmxwlJPCRa4BCtu4HT6A
G3abQY5sY8Mcw19brx9s+1WYC6V8cYfRf0RhxOzRaQc4kXoBx4nxE85iB5X+I7vB
mO9C/1VSWdxsqqucl9W15z/qt/2KxzHsMH21dJvzhbkWbSqocezHHan6ELhQmtlC
8slcGJPVdageKiHO/9LsR5Yt+WMt3gWVGyqfQEVfCbAFP/ECjz4PKoV3lrbBpt7e
WFcSQjIDcw8ZsNAnk1+Ys7zRDWvpL0FmNUk54KViIDiYIGTyYBxjoTtEfrK1S1lY
mhjb+ILM6Ljs+9mp96OXkc01QIjFDF6B0LHGuZ4SZ0ZmpBZDJEUyd90l81l0CTwv
477lVU8QQCO38eL0jkWcMRZKWMsLLXt4a17kqTG0Bu6JTeFYFCxUJdyZvWYPYLwg
pPzpUR3tvmHu85oSJXe9qH+yEUuFGrpqF6JJn3R8tYdoI9NdNLh9FOkN/BReeNmG
6dvtvuonbu2E2hC6qL8pX6f1ZnwSjpEAo5io7z6mGGnv/JPnGDUDW28hNSWB258K
AT0ldlHPPbi7B3NtuSSnFjaxfhMqCY+j8du686y9FqZCEh51ZErynewM8WSSn2Kb
2FWYMYGJKw/6nAQsiVKSZ6DJ22EJATXyeKFAD9j3FjCL0s8U2jJG75ijsDM50K9i
MdzVTmbREQjpvMfvmpC9X5RdEIYWYXNJR9DpS3GN/O5BPSyN344pUco/WH2D2uJT
q1t+c9mFLNqT3lidOIrqqt2HLzIHImZUwuf568+gYqJHKG3xTv7LM15nxiGjnZMj
asCVByJsZST2ZwuLGi7uPNfu8uWfNsdhUlh7ufA/UEm87qWNPknvgcDOdMtfmN4o
q7ueTc97Qla2h3ocKVS3RvE+fQmSbljBuiH+1r8ctDSolFANwB9KWm94BLzkRFm9
oiwwyXA6/tC2esslAlj8uUN6PScRSNReol9aUh4+7HpSgL36bxpzzI0/iA1tevg5
84NeWP1ScHgJ9iDShA0cnvRmXBF1zuYDj7Q3bGNDdSbKN8A4vSpFcL4L6cVFUe4X
8h0/1B02zFgCzMuCWnm21rHiuyddVjNsjwirVNlw2We+7KT3ynAl5XWIuksImN2b
ztPreCboykN8OFs+gV3834GTp/mdjr5Za+KrRMYqMRuqnLeZkYePMsYEHcfj+bJN
FJTwi9rNPz608F1Crm4pToZ2QkXUfqlQIobvzesMYAbeqwlUZDCmqVctSG3CoTqb
eJkAiMmoYxG38XMvQ+iFlL67croIk7lNdS1h/KRjV9l6jfSQcFaVA4/65Nc6UaGP
NyPrxltpDkG1RnZxaKNptfiH4CHbweYYTendHe0G9GxCSkWifHENZbHI9ILostpH
I6HJwJB3bE7tSrA6RKBWw8VMDHWmIUet6iQCnEcjcq6YAYVHLE/y1nzDVhoMY6Jc
//n+aH/N+sWVrKfGFhuNRO/Rm67blPxWi6PLt3Rcc/wUJxYaR5ogjbX/o3iM2RX+
u6FTYeHD4uG4ImfBusEH5wouTe4hi7zwUI64qhqeZOIcsL3Xla/cp8Z4WlvXpN9e
DdJdhHOAe57j3rzJuPQwBfcv9LutC7uRPZ6I+Tz0d7Z14PYdqef1MMaEKXJdeM+N
6fRoyeNfam0CULYe8IyRsrHkpbDvLBD2Od8Kh2bowvF8Lr4sO9P5BDiShsBd/ycp
kiPWeNZySUZERNGZyWHcyU0j2jM4a/yFng+oVsLL1aHbdmytWtqMfP6fWGLgFUkl
ttB+I/T4Yp4ker0ju44BYaYbuXgjcNXSRqYi37aGHBvJbWgXDahFNlSaI6Hv4pXe
N+S0lHRVgDMa2fXirXuXY/3+uScfdMkOCXt5dEUqbxalcGkOxuV1zrmzxjFwA9o3
AYq0jy4sFjPQB19Ja9yipV1tdfQ+/eFit/acMLqQRoAQaEFaHze8JRE5aUJhnV1j
s31igY6UOT1VLKruaWw7dEKUm3C4AO+i8F0KG5LXQm9pWHnv52NaYnTDMsXvlB3D
JwaG3YyC75L6YRE6OEhTVRC15K2QuO35ubZaHTq4PrgxB/yaU9xa5J9N9gc50px9
H3m2gBmrX1bqeMp7RztrgWFhdRyYJIjj8x19QbXUsEE0a+bOmcbfHRZE760gjAbu
JiSazsRTRsywH6vhFBR0Y2JHGyDu/cq8zRYUd3usmyqgJaDEfCV3yIWHvSzdGc6e
Q7E2SdbBUL9vIvmUouxrParlle3Ni+GtD74MXXvtELqWgW4Pxh3hdAe5VeEsv/H8
pbHkj/1EV092H3Aj5Ay34lbeh5c3KZjd6UIn1ZF93Lg2wmi4LPiP5olJmhKEavqr
9lde3A8DhbDr2eWtzkv9vgAfJWaec1CE5173TFIubGKnWANs5ec6VwsYP7N+QPbw
8qQNJjwrdj7MLYndEH4db0KSga/yDIhJeC8AvjRLEZV+wsFGqKxgVTl41XF/eicz
meQ23g2hUHCAlQqAi7LQHdzbeLX40MpYnIfiOn35VACkIhzEVam7Dscr39SVORpM
HiLPrmDOsRiUNszxcvH8EJS1ozG14Pk7ZHO46OteiIq4ePPYhIMOihb2FgSFHRXz
f+puJYD38htclegmL61yt36jJL5pKSxMy98wO2t/KDSgdOnF6MlNc/KDrxryyzqv
btqBCOXiKFuxXsPYQajlFDK9ID3Sz9W4x328/p0Clr02Hv9EzcLUT35l3+97y4kb
w/+8prtUEdXG0EW6tqXejrrPjouezo2HmYQreH0a8w16wPysyTqKxIhHGKysnOtj
O2MvqZLw49FULEb46ax536gDIoVCteVIcVJuH+OFaN37L3tuxKqdls3U4tHoebks
KzPwAbHViPMYONr6Y9aKozh2fHsAc7I9WbPd7dkTZ3/Z54qjq+18PqBFT8y6Iy1a
6W7rSY2XJMuG/F6RjKyxnpE3Xza8PsAnUwGG5hEnrqySeT0EOEvTMsBHnIj6R7aO
5yLB/8es0VmdBs/bl7D45dBACq3Xzd6wOPVYFWZLKFlTe1rmDIdcs7EDoZgqYxFq
xh8ijM3Qh0kIyPNiMOW/wKtbSko3HTJnHMDhsseKLJcaCjvVccY5++mTtW192UpV
OZ6efaDjrPsJiMcFx94HwKCBRkuqOM8ZvbOLlYbTvjTRAR6ViWOz0Om1QHx/rgbS
mvnXRiIdbxVeyMoYVHVaIHz5F3LvTPbj4Nz7qVvQc9o8QQJhoWhghftkTaQC5xBf
OIdEOh73wL06ux/0A7S8IXi3V33WMiwR9raZgxqkxxFyQFFbTEEjiT55Bdaoh4K8
rfkV7IcU9GdKGcb6KmP/c5V8HlHB2mTYZuMpHcMCtnv9unxVNFxkOUCGxEjSnam6
LsIO2UywpvNamKhtEIptorQCbI4UQZb7eWdmLQR8i31gBNyPj90YXGdrNuDBmk/l
9b+cjnx5sCvQ0XKdl8VYlC7rp2nkzdvrYwTn7oWESfDHlgK6kElo+EJQyl10zYZq
ovciMXGH5qeFd177VXCRrTUhNpX9J2Nq7NnVY9ByKSLz2y2yZy0b9XgEv0YJS8jU
Tb8edCozoggxvZspba9CMRc0+Fk5lcQl9f9c2xtRQsp7sCXr+rlIr7IWZsDa87K3
WnCuaiOTJ1jbINAsuMggpTH2IMBEwQi6DSeIf5eoql6Vc/3n2W/JfTBaxf/69YF4
M6xzsWkXr1vMX7B0Zck6OLzO4RJ7UW8lYxX0HJdz0up/1FBhnZY41Ucn9FjIn3dM
0SMViKBLJtg5XQO+yYp8GeK5bjrIkjvOZR4PPRZZ4na2OnqY96HogQusEf4KJ7xG
HDlfmIvk6icxsUWUUYJg/Op3HUhBshbxOssWHBsv/mxM2K7TlvVYgm6pTpimCcjR
W95GAoSpJtlmi0UBAejXU5gD7kWaITWqhP1w9nY04dFpP5pm5SY5VVlRStvWeryc
SZCctNOVLjNnO/gZPF0r0PRASYQP2+Ha+/LHDsZzNUyJT0m26hx064pViau3RqnO
aO/HrRwo4TFl+CzcEouE8izI1AaLfYK3xQVtgjNzewok0XhcG4c+AG+CF7ZA8lSv
Or8Cqh4lYjrGG6Uc7G4EoU71OsBE5qpmQMyBLPjCUryA4snSBXET6shRVc7A+YJB
0EvvoI0a1lDle+mA25I359jURv3lgQinnBQ7tARMizYm14j0NLwiF1O+wrXghQBZ
oFx74HRs65673dNt8k5iGBhL6EiAMVtHSji+hWrt+xjjijoq7Eqb9jsXofndeWK5
lkd4rvtN8VGXrLH69DEUzRrr//6tOGPkX0kasBztHNQS0bzb5MAKRcoTz+6aWYKs
tddde93U9FdC8LkVQN4dM7OBJiowibtqarhdDfWS8q+k+DOyTaizH1JoAsc5jVcq
YVl6Rpg+ZxcI01GbuDLiSRmN7nBeZ7kZZoblRLu5rbm+SmyqYRG4XGxoQuynZ1Ij
FTrPwEkeIkcrja2MQokQ70fHRmOBeks8k0bQRQ2WGS61mrs6DFJQmODy5UIssoIA
a1p5ee8nwRqEMCVQsA2/CkowfOnPJEB8d8agGniQrOT8WeK7osV4w8BaKsn0Bn2P
uREzKNhO4LBGRRJEBBUdolyEJ/fALluRAFHHGI2uoN5UkFlUSidtTwXINgaRtn/T
RNO4iZdl/0AmSGaCBCgWtFXrd4UXAm/r68VLnkFbc4zbd6nJzqwCG/PI7R71C7J0
hNS1BDAEsT/4jRVZJINZ6baUHGjqb+zGQSAebwNAqC7ka02Mawxt/7/ZmJ4xYdWB
00qPRB+91knMkslw13X/7PlVxtACB8gSMuB5d/xH7LmEo/xpYvL9wClrRSVOuaSN
whOAL8Scof2uwxQho/s6RXfl+fUPxCcUj8Y1aMnIiKxPDg6lB5L01KsRCRCNUfyg
Z5BxxRJCw8BiA6YIKut3M/HkFe7OLi/af53LSwAk3JYXxSkgfx49fgN7QC7117Mu
NTaNRZvZzg17eZxb3t0SdR3lT4lqD7XOZ0OP8MlXaay0DtcyVbMrE/qKx4IAhcth
2ggtOCdJ1gbnIsPaIxHujfQUZCIv34euRPV/wb4dgiEiaW5pu5Sh+LKtps6opgcF
Z7Ph8npKa7ulQUck4eROFmM2ErKq+wW98Hdm8swHXqVbd+rshFD/slXKdWe3ZYmN
WlzhVcI7Xd3x/XqfizhilJ0n97vMIR2AfDtX0uaLYE8wHw1iFLjXYOJzqslMthFD
MXkM4m+xKmPZ9fTrCw6LzQhmotEE6ncIu5p9aF/L+4bItusEleO+iAugAc2EvG5O
Ki7Q5RbW7rD267MowafZ0+hLevCJGFPHelyC53MaeDRK6ETRX1eAg9/gs+g5GoA8
IW1ObtQYOD4t9MRCxlpGgPt+n5fOwd3WiUuHQfBisEPrcoxkpayblGiSJNi7f6KZ
aFQb0iWo9ETqUs2aUDiJDFBwxVZ8aDSKaGLT6C75jua+Kg8W7mN87Sd3OU3iiePg
vBswmQ9pw79T3y+kc24BP7x/jTabmQ7VWZX81wnlw5M6U4A215B4wc3hEhoLxPbk
c09oWCnaZx+2KJkMLAMMBeWtfu0EgtjTiOPYd+nLihX2c5x6xcKuEIPL2zzYZt2Q
QX9HDQnqGGutExAJzb3+399lyfke3Wy0iLCrdE+ge0zLLcLXjptm7Lg+hARXt4cv
hCxyiYecDX+ccc3yO6ZzCq2SQt4tVWFpBSC+PgycRKUe3lz86FNYqcJwAWn5mmJq
r6N+Q2Bu7GZOURVdl+u5X1sgmeU/tUVlf0+2JOXIq2zyUuqlKGjXXjN7ZH8+oceJ
gC5CroXRb+NMhCn/NRFauRwYfwXl+Tbt/0nqrL5JQpoSi7bmh5iB2nSJD22iRVoD
eT5fEkoHAax5IxKPTjzlsPvs9uJgVlRahZcr8H1lm/oV1othHMEj+PWHSqfULIrH
YQrKHQBxZPWWfT5liwbufSm5grGSuM0dA4Y+MsX04wQvXkolnfZ3RI+I5oEGHDGP
TvnHTyMAyZOU4Z+HMWuhOLvptfjRndndgbZdQEcMD3ABt8CJHx1hzGSZDTRo/Fgj
w7NEpD6i7EozWgLJsomec4Ug6ya6qVZ+FqjvaM+Rktfo3cAZ4tkoet39D4hGo4wY
+hIoqbbQP6lIWzhV2yObxl9nn2WN0Pe3O4zZddfRtx2m4N9bDxQfmgVoxdPsQ2D6
6iM4qXU76Cw21Z+JW5uNaeHbeR/MNRHq9McwH+hoVM3qeeH6+x2UUVEQLfmf0tU0
WiQU1OSF77YhoPi7vp6KAnDGfwbHn/uvXkMkf7LUDW/j6leu57T62Je8/7F+QdpX
phBvlGMj6nhZvsJT7PUWGVVAz7jVM5CHDNRBQdTAh68qQ9Bk+oKd0rxpAVk+tANY
fThb72Kh1/rxdrr+e1OFY6zHGgMllPdLzF+F42iUhHku67BzcXHXh2gnEIBlDkAX
wtPuO200F9R+rkSTWioHIbAF0Mcvjve16s64WrW8kK87b/ZmX0AwA5xB85UUrrDd
L5HcI1LPKkz8hwxw+JR5ELhegULu3KNbM6Hgj+mq80vh28q6t/CKrrna6Guc4XHP
m+PrUU+iw16p3H0AfY3iM73fNgZ77D0lAwo+Lm/kzc6pwaJLLgfOeMewojdjd/tE
DEsxCCfpncmHAav3oEAKVWyGk1R9Qmwk3b5voQJ6yFpbKs9N18GTA//vForbHbqU
oT2JkdcpBLm1uAMmXXfBom4HzSPzOX+KawCmWfxOQN6Dwcr+BbXzgD3sDtxTX6SH
4hbdysrKXxOZEt5AuMkLdgxkuflmdHX+FEodPx+DkwEMCniOnSjJ7jYaiIkd2tu9
b64EUqCjZC5ms1uLLYihYO9/sCApWrpeSWNa/RmAPkEdB8NCMEsBz/5mg80mHGZ7
uWwpwJNOo5OY0vJ47jH0I27mwmBTt1foAMtU5AQzxuyON/2J2VTl05HJKtHeXX/x
SEHnqRk46PK/sjjfCOW1lKnoxfwZwGB18JOZWdlh+6PFY2NA9WzJyXf/J2SsNUCS
/mapbwbKzbTBQOG3mlm/On1AdxSVk+QinEte8Z5lfTjjf56dNYTgpvXXsEYPRN+D
6NWp7cKoqbCZSB+7BT6qJBpY0h8HxQHFI4PvTfwVwhvHG8U/rqaX/LVFMCCmKStz
rLfVE/Uc3qQJKe8iAv5ByYI4buSK6RCr2kW+SWX+LYV5NK23kNBvOUYlnr3f7s2I
l8bbCUna33WeTUSZn/+95HMnNkOg64Wz3GCkl+ULqDyRzkz5mE69JKAQhqCHGHIY
xjqygiIANfHuzi3KH9z1Qie7yI6CtP+453glyOGImpXPhGfVrQx31OHNf6fmKkqt
1+Jt0tfQKmp8F+U8CgLpeb+mp+RRZQgwTdndqD4Dv76obfVPgDod856ViONpxALK
O5maCJNMYBrtlRWNsWrq2sMCb0Ql4E1wHtBbCL9h0T9OXrMTC4YPEhScey44cnx8
Dv7/iTiCnSjNDdE3kWkRBilfMh2Fw5hTJgMpdDor4dVh099HvNu57F2jWBC9R6Mf
DP4u+Y9X8YiDTZQ6zyNA4qmSvizs0D6E6VWCqG5fDGHZ9UN7reNLmQP2bMNz7Fvj
bcYp/IptwA7LPiIx/cr6p8LYg0eIONXsDoXmaiZ7kxBt+phKVQ0jmQJ23rQIB3rn
f5MwHl8JFts2qoBnFRsN1lVDI4gng0CHriFEzU1TORUlPrKDHpT0U8v/Rpuz/9qB
jgsxeNP6GSQXE9t3RUUE8JUQMWFgqQIEriUumBz7FT1ceMZ1mMrMFejcFqQtoSk5
fmDroAGv4DIpZE4mtLtYy9eX7010sK046kh4k4Y4VAEiBAj6y+qiw/T6gHkbG+Vf
I5wHA//cThbzzKh1KC6/nNbnI0uzkwDCMSimC4xQ+SNmwYryRxFPgKobAO9+0CnD
lK4cKG6wgtckRXEmKLvMApzux15DKtlxYHNARZO0hDoV143yW/V9Ltz4q68FoKzy
08X3p3r+zCofPWos0kJafgNhbQ8s1S4BW8Imrmi10wObSt7Uq0WwR+9XS1cok+11
do+FLtUMrmj3FG6uaNWczlL+NWNn4ksQbiLuFtn0xsybsoCPJmPPmpiNAvu34v37
nw5qj3BdiMyoTDKHrSx6vOIx04xk7DN7eNQpcPUCZ+mJ/dKWC6Nxn1/ZKUe8cO6t
m8FtB0cl2oEJsqwXqWMdBoDNl3QyyC2Brrah98UgZ5CW62M4eGcFhtGEB9AgjQ2P
txfO3C45a7zYjT6V5xmOZMtH/YNtRhTZPPvPjUTvoK/8HY7EfdBV5pqCrrCRpHfp
XLiAdsW6OEZrf2SkDwYVXmnBsyYsCshbhdNmy1W6R9rSwb5DpzC+v+EvFAiZ1fdS
EfLEBlV5STodfCDEI6GXllmxh/h0q0wyNQAul0hTjc9E0kDwjyu6iAPQk8lOm9sJ
X2PAxd8lArNdiWZKm8I3CWZZksAHjk0kh8+W1VE5PeqlzFKHr1SlYQEuG8wu8vjG
EArUYw0fHcujLAZkz+Te3O8kBryPJWpleXpOK+/zHvCL1Do+VXOKLzWVJyGYCPLv
mzcAX92SWgWyyV9s9EbiLQkjqjvsqJPGts0PqFg0TulSmGuwaR7oTYuQjFb0Z/oi
JJbQJnHN5czA9gEQ+KCUUsARofEcShQ+045OeJf+YUAvQoK0rtD0raPl5PvjAyQu
GvT7b2FqC8ACaeJfNUjL790jl//ZV4CsNs8CYUQp4SwnjMAv0nqv2pBUzQSWqHTC
8NVqLFqCAOgHAMq5mmVtHDXqK3pfDplDWXC/JRyuTdN2/ude6Nx4juriAsldQF6e
RSaegzM5CwE+17SoETfa9UMcV0tiIUTe/+0zg59Uav1StvsfbKaCosDsLrxrJBx7
DcE7//TLSOcQ0CVGPK+Z3NY0Jfn096GpQva3RPIo6mwjY6J1G4rzzMwQ4JYe2+mE
PeeNX/P75tdm4sGVeBe5QHbCdaYdfSOgnW8zwIwC5r71ps96AU5pPWHwPbnpl4al
QHD5SSgnSxqF7mr3rwmLfG1z6Ueofr2H7bmeiTaFxRZr+4Br472Z10T/fl9YsYB0
K8QXsAb+OrhkJiNobB3vTjZQLNI3/9RXbuTGYbGldJqoX9Os3OO+moIfDDuUZvq8
jOfCVdhsAhdu5zmLDvQcGe+7W8plmxplXKQ9/mdo2ANM93XIgdhy2lm7U9668vqS
BE/mrDTQjhm3tIaUuQwiN6RDxm6e3Nl+y1FdLnr5fBap6ShhO2WfDLYPuGZ4lK9Y
HsZIhl2ocyjbrcfv4fd+ee9vGxrIujNXZt6gpRFPP/u3+0ypb1N2syKQn4Jqx0xo
YN454AwoS+oHLkKbxUuMz6HfXLdHaXEU9jzt/dBAPB4eVpBZK+JoXCxmDflf2QaE
I4o6ogdyTWZ9gZpviAlmT+xaErFDy7Sl+6YsQj8ERTVboWyl936xj1fSlckBlo1i
aWPlxLjvasLjnkTvVlHCsF4FW7FQUcZg1XphWwXL+5W01SB2Ya9nK9iQPt6oed3I
/VXkJuuEbBJ1gtggPrjq8iE68pemVzaALzgq2WhR06fB3ydtU29/L7s3SruWRJ7s
MCVSmzC3b5xf3QovlpdM0QsKXOdLdnVQDgK7bp78+pnNLw/j7tvNVEf8liVFdgzz
7WlG/ChSaA4BihdBpQo/W30Z0ypS4jnG4EHcOrNTdRgKG4cBj+QQc68oGRrB5IRI
Ba1jq1k9m/H8JMGqczM2hb1/uz7dPaFZIXWLIqR1Om1wLaBQI97NSqE2MS/D2Uw5
A8MmIzjdUtcVluAmADnOEFRH6Lp75MwRWnkl3svTvnWGR6/sXqEBUJVi6Vw1anfQ
vvD+/zr7doc6cVN5+H6iyF2prlrF7+vEQgfydyWmajEIuqOB9eU3ljcKxbrt7ugO
9BdLHZEAQuGXz5TDiJwZapy8zXBQJ9P0HihVv2MGI2dYyXgJG1Qeiwk33Xc9sHpC
LSlmGWkTpx5es3zzVcXzTWogT+rgW9durT47MZzFy7mV9U/0LJWKtGAZug6XXFib
5qVrFJ5tQIbylPAl3nDsmHy7B4sFnpZ3EdwUWbIZBBHUqvZClSPPrt762xGKIFFs
B1x0cHXrLtYIDfTDHJcChLfYy7a42IVWc1yQ8i6bztlKDJizpKoCCiyhcYtyfXdG
VnP010a9xWxMkYwGdgjhDLeRhb7vSHj+pBVRphNuA4nR8fEcAgO6mJghv5+B/1xN
a0IeHL78A7zscvy0fp+AiZ93545NN5Vq7nEg0zb/f9zuXqeR9y74bTFwUk5u4+Vz
dMSbfMnYgCXJbomZIA6JMHzM9MXkHxTSAMAs/WBakLZlTarbpZwfOiI3eQbR2cGb
ZBfGp9QRcSajoaf4zMxOS4oYl7C6DqnbB7KoCLaO1qdlxL0E1nHM09nqvQpoJ+gh
quK3QKFCrV2lIw2VSLQ3+BpkiZMAAxs5B1cfeM3QRTjqNwsjJj2r/fEIT5pcJZ5r
BKFqzVJgy1+syuXCgyfLve2FWoyVBJRfx7J3F2kI6o2Q2/0D0DfSxIwUQ2Tfvw4Z
3B/0nzzd6d3e35a5QSYsYUDLxIFNJyLFcX79yPPjVPhSnQwdyTfy5dvbUSxxs+J0
h6SU9QzRuPeLlwWdimtC3voIUZEyjyiBa8Z6z+zw0d7wHFrZAOmpunUElGePAbo2
uO4ssmk699IQadiBFvgymF+519AXBbv4qZ9SXSaAd8cn8HdK/z4ZQLGd6baFFo7U
C1LhaQdQnL4SaOoXUBG7r7Q/fcREQhtkIkVA9T0zKugydERoBp9nmJCJPSSQLcHd
hmd/TsumEc10uN9FXkK7IfjYvSH8OEkU/QfBeRYpTzVFmNDzw9+CbTK4rc7WuYgP
6wvE9JElzMNbXA1nIzQp9McTOkJCxVcJmvQsTDLO1aFu4HQzMRO2fmIDHKuk4wVK
rMqy9J7Al7o9Qauzo8na3RDaXlUE0UeOy+cQ6e1Y6FrimzME89PK/rJHuhsSsxhl
TLKYqWFleIKVIk0F7meF5xiQSco60HxzWvahWrSpn63NxQwXNf6VdZ4LgeevmNeC
j3WSWIP+AkIj2lpvIveyQhWBpVpixAfI3BSyBXJKXa3v5/+Ofy/r/UW9BzZ9U36m
w/rwmFDO/JyZSGdDccx7BH0sPUWai5aakqyydneAz8LRgLhnXuL34zobSDQ23FTX
izJuc6Wds6lhedB4upej8igZIb8upJjhnN+iWJ9JgVIuFkKSf/gn0hLXZOqCNHim
vsPJRGFumkGtvsRGpgKbP5ypCpwQvTxKiGL8XeJjBJuC/cyTAfUxqhGCRtKb3jYC
9Jcg4EUzeddsStCc9XCCEAHR8eGf/Fbg96vC7ch6QAN34fvVkYan6oRaR2ZTwpSe
EEqroEDEBOGFJHXAAq4jYRtPsGIrnWFPnz0PuC79vDF1SVrnmcWyIoJK1M7WjMjd
InogB5NfB3wHY9B3WEzHvavHk2PGM+KNC1vbQW6rq1sE3/tZrdaoIN2EYpPJvZig
mPJpVXyZqvAOOroT8f3BARXGuk2ZBFprFjjf51TboaEbAi2DhiXL0wWeeprkkMwe
QahL728/XWPsEWJzyLwYUwqkwX8zfPu/q6BasovvdR8qziamKc5VFcye4yerhzcH
DcPC1U8NBtUQ8osP6xEwq9a1adiWcW3Ke3b4oKnbYKS6n8l8lUGAD0PXLGw+OvFZ
xkXram4t6QWhfV0/tKX5y5DGhCTKzlTKY/rro9KjGsqd+3cq+BJcHwaqtzT56nKp
FY85Mjt2I0nt53ShsM6qb99AknvqiS+Hb/3/t6W2rZ9kM6nORHjgM74xfdhoFvYK
9BO2Iizy0yzg5SlC5Ukz+/uzZzdxYDguIbZoY1Gm9Np7sNKiQHfYWYLdxIL035re
CVoy2fJ0bV79T7KK6jrck9AWpEKBIe1bFKufBihhJsteEWuLrWMM3sKUjkZ7igVM
YJ/s4hRDqhuhxCdvNgT7FZgzX8Rw3k/DwxJp/LQLwpe+H4qcnHsjhA3ipByHyqx6
f+85KbZ4+T93q+BRsMT8FOuj4If/JqHdiLBEaoBXvm1lz8c8HlH27nSs6AQImFB0
PE+0OBOe71QnrtwFlH9gvlhNryfGJH8Kwf1Au6ZcycAoyK5tT1qzV/7fRTcZ1dZP
aSmAlXyFGbm+Vu+0vVDVGzZtXCukGP3kUgRMl3IB6u40xdMdeJtKHY9GkTVm+X9M
rc3urJpT8pDt+VsFeWZvHIBN6dgC1LSp4tv6U+y0VJa8PJULUa3jR8a+rZlDmytZ
IVS1uWQjwLgdvXZT/CaitFQkDBlSKpUtCxbTfIqmEAsKFj6EqTn39yh5cT4JEv9r
Nh8N4a25iUeHBZhNgnjai39nSGCs9esTcczTtJeYlsxNKfrVjn4iq/UXkepRw8xj
Ovk7UgFaoO5I40473jC1TXQbcdrPH3hAB2ercq+EmZQpbU2RpXMKTEx/wNnJhrIM
S9VIm5iS2vwOOOAxW0x4mnVBPdz01/+yZYISpCKwa+lQTOaw195eBDYC9WWJszBx
rtMqApAGfjP4Y2I+1vSwvZrMLiry+yavhEb/9YuXV7mDBWKFywz2+qhtzDi4jwwd
cJvAvzyI0xy+EKAhuMfhaX9IBQIIwmZBvhOfsKuEt1UaeWtny/oRpX3FDV8FhhLe
smj3S7kXcuDdztJBRk3tDH40aoUwGdHDg1vFzRjDZCwPCjDMJI3f+wApyFg0K31d
2vNjjGFY1ZRkjuB+0Q9L6BwdxvQg1p1ikRFiA2GaDNwjSVEgRNOFc5aXUqUm7TDv
gXTXecxF7d1QO5Rl+rSdoO1Lnv3frzscyl6g3V07o/0LbGSOtDU/1mAgldf8JcRv
faGOK6FGf+N1QhQfwQopvdfVjp3FRIgRL927AuhPehioMBpc7kglzI/E3DCj+lKu
W4WRsSyVhazPp4JmMaGSNMA8CazmLVo24V+y3th7r9i7X1mfWbAxzvqg+td9+Ykw
LGbqBNOzNv3f1T06OoC4etMA94m/HGjK2STyEifd+O9S/h00ZTIxbSlqDV8QabeT
x1Kzq50v3NHwUYkUoD8TlxA9JxU3EidOQ4cFzxmfVom2r9Vd4cQMV3DH+Mawsbc7
/eTxw1omPDKl4w+GEG2AaWfTnUIkeeuIvng3imOmK7yC8VsxIwfcMvxgnebS+lBY
Li+sCvDfpb/HCSiAL8FCx93zqYIDmJsHhvcocpNkSkK4iDiDmTvkdrSn32AduSB+
ftVFNKxvETbKBLQ60P7MitT1ShTaa5zKzLb7E/aIelrY3hyCpJBZkQGAVleS7hMj
knQGPCGDlh30bd3CmnXJKt8Fqu9EsjgmJu9ESc0NL/Au+qU+YBYQBjU+g/M59wNU
syE0eG2bAKYqfgNy97zSP3An2hlqOMeQPxHbMpMygmGhvBbOcoqAwDJj4+1XBFk9
GwMNO6vRbKWhxlB5IsopuSfv5LsZaGb0KAl7FxDauVL+IEnOvlJ7cUicRrtaK9vE
aWrzWRr/uPx09sRluhbr2fSGHtkAU+IstwA92DCR7FoTAjJk2jXB7a30WIR0Oaap
se0U5J+m5t1f1qW8KPEyTLbvu7Pf8ni0FA6RpyvBb6u0+nRN7EfoifbVI+UjcG9F
b16Z+hkIJ2SZpAhpxoqSOYWtdEgfm9HM7pkus7dglweRykO4Ftvv7XWDLdIPAgTN
VcwM009dorY3iGm/99/MWB8uvJYuNwlAOCpt2dW4jgUaK3CwLU1qxKoSsVslyAKb
VvGoVGwfFdLI4v98FhPX8+6m0tLww5505Acdoblmid1YB2I6y4LgGVkVlBySBnO3
jfjqXJH0tymEbEHOM7hQNAuUUUw4wd5fY0EZINS1X2SsqmphFfpqqoYBsIjpgdLR
wMiz9r0HeYWiAW/f65+b++WxaI/5brVdcRALxs1+ady0c1g4XyepcRntPrEeQU1d
ZR8D6BXWJavV1l+ePY7KJA+jfD5wzh8c+q9jmWVkc0P2GHz/QZtWdFYKS+aY9etG
9tSgQfwt8r96HpBP37TliG0+GeU1ZZeoqlh62gDibYnFAep5Bgzw+K7bxiSTEq75
6dlUeURuVjYlFzukth3Lr+tiYjFVvgBtrkkf1qU6asrATtIOfXtUQT8e3m0aKmZ2
Cdj+iQZVE5AXDX7GZQterDAP1fiyVgaV4KDX0vV7Fb0h7ZQnMvnqkr3GDpY5GcKP
2SXSjdTsCmcoLDoAs4Y1s7tarh6AYoge8myXIgcAyXN0lsqDttutNpWmPcA/RB2/
pabPL/yKU8GjXffHxjI6IT+0nhK6kaL1ENgNDgK9lffq3vwq6j1fHG62igqheBA+
3Lb2fWb+ikOkzKXlEU4xJI6oz8UfM4bEeH+nUKnnZcWNvAvj3Ss+SCRnVgTLnEtm
/Il1b2IpOw1CYQuF8IVV19yUKoSUdwM4/SXjzRXbMDlyU1t7NR9Q9pls1tUf31ZA
dl+TQCizVZ6FpgE6m7ecjxpjSFvcXWuSvrLRUKmn3GQd5MtJA/hiQ0rtiRWZmRsI
AO+MazS+LrPePa/nNP8aicz4dtpPnN2IZk7DJuZu00Ahr5+ItwYjyena8VzGVAxE
R3zpc7uUzkNkRtx+FzSreXHqX8SEVbLPaeMOTjGDXCE3p7/CaKVTmJjnPvVO3rJA
Tp/FS6WCPFhLHRTkHgRqoK8NBRzxUpp0KHTnoTMaF5+Jcq2LotuXoRB8739QF06Q
E6M3CqDaMk96RiRCDAhVcRiiFhg3eWoCIu8zIH+aJRt6pvmjEQzL3crYbTmNHBjM
LMSN8Vnz4xEhF1Zf2RdBXKaZGNZSKvbI+Qj0BeYCaRWUx93gL7hZ9ASdyrRune1D
QdWwl1i/8U+7iJA3PTwWzEngjlgI09KJ5tr70R3B30dedQi6pFg7LKPBxR7xywMp
d2nRaoaHxAAYUHK6jzsPcEEAmgLp4pW8zIuB8tNICvbJgAu/nhqZy02zu0S7ffeC
xlDbokiLSeR7on9YlL5NK+VRxtRMCSBqvZA2sTz7akRpKcxJMDx7/ERxmA1BX9Pa
XyOcWANy9H/gWpgb9s48l1fSAgNGwjZzrKLbUGiUKSt6883mm9y+HwH0CAvLG6Y+
XMxkJRiz0g7rIZN6nH82UsPxe5uuHmwnwXzIPjw6Qr/BnGpUm9Al2cHa+bTdb2xK
Rch2bZCcheuxV6qAFGarO78D/i/n0rbNVn5xm070D8ppAu4jdeji29Lf0V9ObGUQ
D0UyFsHmch07pOS4imfLuyYeLZJCrBZ0idUZBXz8bqb+SNOsIkVy1es2+SYklnww
POJnMEA8oXoS+6zpAqBr9Jt71PG5p0GS6nr8t5W+pzsKovptoj1VwsufIjjdDfSm
haQO7e5MxueK/PgSt2wrGkri8rCAPfbZ6SCKI4FfLKv3bLK344V02dYSgdbD3h5q
bW/aWIVDvSER7iKPvLD/sGq2gMw/c/3PJZ8nYkwMzmy1HNde2VuorQhwc8WHaB3L
Q6WZh/1xBZYcMmIKlFG1Q0gaD8BshngkvaUg7SVYCVFs6fxn/LhTCPTrzZEFjB7H
feivWcL5LvxYpWya0NytmYRXmf5/1o/4NU0i6WDqx3srNMtTAa/eiZRnVkx4Wo5I
02r8uxi4k2YJSxvcolKJKERiL0MrBwn7D4+FKZlN0Pn9dSAwpOGKPlcugj26jg/e
gq7L/XzjzpW3h9X256mTwIgbM+CIfN63SIOAffDjoNjAx7DKPvmolgRgyGsmeNIO
FE7CkHKe6TYRprGEI6xi+bJc2q304+ylC7AnF+TrW+gJM3k4RdoESjMWKVuCO25d
kl9NUFELXeOFm4xXlyEfiOsIDudnuG4sdpOSzDUsWCatBCHDweakzwZ/IpIRkUcZ
CBXwNFWymGGfWOL/r0vIorbYY0KeEIlyAZkI0ML3DPfgQjJsVHwPLFwg9Rbg2kgb
KasY0G4wNCgcGB3Cqp7mDLTSWPbcjEgvC9Skeix8k1yoNTOV33Ies26Bzu2wkpDs
lzxqy78TfWCOchvMHQB7dQTYsch7SYmbudx2SGD5cMMUVm1nR3yXwz4iZuNGmjuz
xLotIzOHSUUSOGQMioQyCXKLj/N/eSzfVlK/9PnrXTjdUPMX94gJjyfbJoQIi6H7
OG2jfabFbXP55YLAi7RPdEOBZZstgBrH1GxJQzLHs9Nj2umLo6BsW9b/mFIRN7iK
uy5LLoHko2tO4SpV11KMrQMQeUnmsNlIhscz+ewOqnSPLvKt0kUypD6ASF46M4mZ
vbwR0aucSlXr1BflFnt5F9nuKWeB3PE8Gq1Ysg+aXeYEcsPD4ncu/L1sut5SZDCs
eMJ4JtDfHqhbCaF+mvX0JVd/r33tbL4yU5lfi7Zwl4FQRF4Oqdym6wpciU2GyhYq
Ow/vXkI/BL4ps6eQFesdBxhuFNyO1okc79m1Cdv9afN+rg1KBtGRehMQOAyNPLuo
dufGfmd1ZFH/gl1fahkLyEJtKVfoJdmAiutDNLu7IEPX9EeYHdh7EdHpWG+EjegX
0DYbilLiaOwTEDU1M2Eekw0AdrWFGpcn+UMQN85S+fCM1JOofTcE6OgQ/FCG5dwn
RMOy8xFVnYcnC9bNfPNuVevBUoiVOJwiCYJVSpS8B3Xrni+9lAEMYSUZevD8du3d
2KnSlUsDLTNWP25ylNr3MXMKRZECOIVwupfuMqgZpzjLjR+7rCcpTvkhjIbcQ7uy
yPQLFHQdZdRix0LfNNzeiyYZE7khOS2940dLaJxfcjTFb6ZqgGMeY9Mhd7uT3rkh
DCz6pvKSyMwG03fwrqR7vKr/XaSuWLlGMKa6D0aoO346AaK++AXr3ZhqNvd6F1e5
CQKtTLrEEPpZcGS4O+HQKPls5DhlB39Y5rvEaAs7gf20KPm46D/OY+fElI4COoO2
lgpPitHmrIfnM8mP2rQOVi+x50UqWzvfV+8qW7OiZ5JcozE16znb26pCzthglOmE
nRuzgi8b2XOjjNfjwVbm7mZaZzc3ItAlaL+xqSoICjcgCkg5IhvEHVmPavNioLtQ
bp4bgRPTxc9WZIX2sXciiKEfQC12Fs2g9HqH4S0wE9oUEu+mcPiAQ60Y6hHn/66Q
UC153DPmfX4Tlg52vDBox8dL2QUA/JaWaQUWRnbeV5SycpW4x+vXJg1lqLVvTYNl
I/1kLqK0hxKEi47rS36a1C4cpihS8dWk4Y0x2eEmGSDn9ahKppHstMDrYglwn+9s
B1ko6XnwQgWPpygQcUCmcaHwLQNKAzQ6dPf004kCftzAw+9QY7Q27IOT+s6WKWd7
06qhFvF2X7mc9x3aVo1qchB7XpiYCXAeV0n///OAarLo32yvktwiaGc3E5CoDqBw
LMPjpHo2+ejm4G3BObsmuIyBzavv0t2XM2NbpnVWn94UtVquZkkiQjayb+wc+CBc
tLKfgI3hu0khi3WfnnXwU0TVxFcXAgKSDfAmnfZQ3gOlJlkZJYhYeKxJu3zghjEm
p0W6M0GVN+YXi8bDAR3ZkEcHiM1cVJiegfIXbWrkP9LUUNzauDuB0VDZ4FvBUTmr
J/T9k8+rH9KarqZRW5+5KynOQGzdp3VqQobD7PPoImp/OnWvscdK4Pjr8RCNOfnG
TeD3XeQ/DiO3FTNCf/bTCsyQoifPOJwfJTGjdvnDaLXlBZZHVPKN1q7OCTUWgxbK
4KtWBpyFAbJOIyMkNqtDpJpyKArIuoNJ6xI6ZZeJzWiUoNFzVvhslA1CnMk08lPY
Qu0rLD4h3TtkfpwEpYlqiOwb5YJP+BOXQS9alZhbBHu6VcqohWq8DAYsIMFR/1e9
WTvljSGsSnN73kr3Zqx8aBsN1A8MuXeaOQiw0TtxCUPNr0msdb4ISHeHgJUbnNU6
bkkBDGNyoyrCwLbl7M5uZVZRlH259gOgPDr9pjCz43rZ5UkXUsMkChtvnkWkzKgh
qs6j+nkNYA8HFwG94V+PYg7F3YUI5sf63U5mWqvcgXu9yXn5XdkU+FI2M/I9/0sl
iqyAfcJgI2iw7zwurlDKSDu5OBoFjpSBcn6J2ppq1WUSWVf/tWU1qIvxLwexJWRJ
iem+vDhhwwmWYfsk1qSYKfof8GnsjVTwKSSoaU1yXWKt+hI3VyxgOChn6cH6gdcl
Wjvpf/Z4MVFTZWypKlExSWO2gaa1w5XGqAoO28dc4wyeeKdUiuoWoFFOzN+MTd2T
IHnKM9TtNQ/4dhF7eUuRs+a8r+pyxtwPyDhVCA4kyYDPU29gScQXKgKwV6gACB/S
XjA2RthvemeJlVGq0dC4onVCkVRKLR3m+1FzTXHC+62P7ZBbWsQNyZo65eSFC0Q4
zIRimpSi3aYv4Jg57QL1WccV9K2FfbfnUgcLGColR1eBCYx917peq5zU1MAlIFKY
vC09XG6UX6VFXDVSVsN55jc/JuB0AGEHQ7Gyu3h2Z1NNHSSg7NCgWcsND+SGDwYJ
i8uTWk2aGNmQXkUFQWFQjcwWtOVQe/tg2gif4m73U2ucK3O6cQ0Fnf7Gwxck1ZeE
SXyHMwsNwuPBAhRuacAXVZhyfCGhvjv3zuP83Abhz4FZuLU5QNWnUUm2/XUDMFpH
o7hUZ/xqH6PrJWmfB0eWBo+jCUcBgfIimEYunH0lCYxplvk8AvtUPFc/CVll8jA4
afwod67Np+CYhGO0pzhcgCzFrSPdVG9H3BsZczZLJpnqbDSH7DCXLO7o2fFwoURv
gTraFIUcQmzyJySHZtqABkMcNaKhPS10P1RacXOqBilegw3vhC654n82u7k/2V3a
e7rlV1fPvnyKXlcA0TpMvpvxi0mSOEBXyD56pXxKuwcU+vBvdXWLpmMihr+gqECS
ipdPQ0IIxjn01OP1EHG3eS7MDYHkOe26o5AKEunoUkAD3udljJa1mLbEt1ir1pn8
z/VGZH1sj7mLX4UvDmlTyffeNfy9E+GGLDcElwcNuKTtNjE+6A74zxE3+o4Xurla
2sb9zykafDTmTCAaE4IiNxgnoheb2yyIU8+sTW+81/O8LTswPwaqsENNHHyu1idr
2t2AvP/QhqQ+iTpBaiRIFXSxCRH7II4d4SHNJo/p3oTqg41dm1IR7gyitk+VcvSw
detfGZ2O18hQ6LmdWlehEe3P35eMVMVOnyzh78/UltFfrR2m9pd6q1+swYH39N3I
ksXSdxnqqK7tZ+7/qF2m4IMx6WBrJABmX0FJ6akSOcbqDn1CgJr0m3UurAjoudqj
aZwq3UWRWzoIsexgaQmViLXlVa1NWqti6wetY/pqdh/SDk8cmWUC2de3EMHcBXPA
Vpk/Lj0QAEDyBUG/JsP7lZJaugAtA7tPJ/uDONhWUYT5fXuM9lQW0Wb/VMm+HmuK
9eSDbVzG9yCxhyCEtI98KOcadR9RUnWBILGC4/Wmwz4tQcJTgmb1o5cbLEK/PRz1
Fm5AiTQ67tlA74U8jjOt2qVmBS/r1Svyy7RAZMsEgf2w4kpCI3VY465ZU0EUGQer
rJcCPtx1kD3snyWAp/K3x6Ov1ys2xORKpFinDxbivV2kxaBHwkeGk8Ce3ZuDiQoB
svEa3pq6gExc+Ejjum3ClqP19Lcul7l2beRUSFR7wzv/q1s891cG1y4O3tD1tm7u
bsJuCPEQnkH1o6soUvfcqyF2j+F+UPzuV026lSPeo6Nn4n4pT1RDZXct1vYi4im6
IU4HvzQAytZINgUkObcIXqst//6T+gAYvbKH/ipQq5mh7ECNd6yZQDYHBH1CGt44
pksR9+jZ5wev4a7wsfPgVVNrH6U5bHI1HfDRqQtV9IDHlGwu4uRbtck+9Q3VOHCZ
HPCZmdmOV65sZZTFGQt04FnNHARTb/FtYWtdTc7lnF3jthPmcDv6SW8Izi7QDguS
p5oEZKe9tLT3z0uPkOOyjuu0pCYYiFjhEmFA1Za8MqCeeQevF+IMQvMDpWa7Bb04
j3qqY+xXBFyDfEJeyLG03wVk0UJq9Q5yapr94qEziFDbZdDj6pKkK4Itx099pwAn
qL7T6ur3fBOk7gyHzIBIAolWCCwzNYN0mwQiL+gcS3M4npWgcZ2ul8K5RjjBWh8p
x9XE2kN+eeHVb5uN7OV/ZhIv27txmBkro+wYw5nq2jQQZZyRTkx18mrrzM67BPTG
Ahi3O2dOvmVkjhFCHe2r/CWgVG4qAferMMLCUdAC4pxjsMenuUZ/b2Rvj1PIle2F
Kxb8T8TO0+FBsjNeytBfz7vbpNzqrGi82QWCdg6NjpBePxIPsL5geLT4zS/6Feti
MbxCkUCgKnGQTp2Yw6IOKX/62id+u+2MCvvvPJ6A/9BW6Hn/OkI3JnoI2J9CXtl8
QkQSBGpVT4m3Qa3pG/ICVAN+zgP1JpUx1HZmGv8a2j6KV2uTvavrGwyjbZiS9j+g
gWh6aER+luZ4yYorLQuj7aMP4IsV7VYPgVPT4iMwIN0N5S+fIRGG52zRo+Rwmh7b
pd41SfZsClBJTaa4Who1k8d/Fqo9DvLT4gfqYAqHNs6llZaV1vrTxhscGb2ZEpI3
+YXYYf1hsRYcWfn/xGYqqtlcB3uNlz5YF2Ns6oaNDxvyQrhJX+wSGzawMvo+TiPv
yl06C0KgJF77Nom75ok/wV9Ne6UJpnHxQTGr1A8LGpU3xgUrxlIcl66m/OpgyhIM
s6i1Z2GE94YP7RwevxMBbqL/hfodwRCQQj/pm56Gt89sbTh4fm9SyYWGBN859zRT
AwnjMX5Ds2yBYop+UFfe6djf22CJ5/8aFR/SZw3POGK1sdzgOxL1TzCgqO1UFc7f
YM49cLrnkAe4frWdEyAT+uLXVw+hvpe5L34/2q5iCgNAG2nCOhYfgbZgOpx12hA9
WFinLKoRorjz87vTbOaKXqD44M3Fsw4+ZEhHB80pij7rde6bMvI3tHMHwAg8Gfxa
RR8vw7zI0OMFA9ophaCWNiL1S2/HluGFc3PnHmstSyQyMSekUdM4VlbOVesDCCly
Rk6PBlZfqk8eXjFZVlzzSlk6ALBb+fGWLEU7xgG/02MYY0HCuqhERrokOueLZGsI
2kYRbZYyKpuvQgyyeYZF1a6+gC173lBP7pruI4D2HdrZAnbf8WLXcEiUk1/vcR4S
EsIDgzZEVZZU3sUQCSjoweC+IDf7ZN/IyYscxFL0dKkxBk/gYlSIeKz6AbH/q9kE
/nWMzpx5R/Bl9+F2eBBxswDAvOfoOxlG/l9LN4XGMv1IZWFC+s3JWfDh4FYVbzhT
JB4fBufY/WBp2DUT40+GTzTgpxqj3xNiJNaAMwzC1LOhbZH1T5D6+Bm8kQ77pmx+
M3Aw/xmjnqYFVhlkBuobz5YCgQit/eYV5SGWm80k8synaKqG7uvHTdz3t/WrCeof
Vp79WqPzz9lrT4xqL0v+9UVyfxyY9NzaYKX2vzG2L2ISWRv8vvlvrCHE/DNQl+Qd
tifKG2fxo36xckeZ4L/bgMQuFsgrOcEq01x79bhXK0IA0sXz1EjbdYNFvuKDUtdm
tBTlvSQJ0DQBvhYu1RyU+oV1cQVZCze381YgGJgSlMYl0TGTJ2/G8E67FrJOFPUD
9aQqIvtGy3a51PA3MLcpYXy/yV+Buto8MlUAdoTmLPMTzDmbS9B2v6CnGxt8LgH2
fte5/O+WJR60e7d652VFPFcw0U+wa5GXxRlmkGFIHClYcKbjGIc1cxeXrpV7/whV
jdH/HQ00/2K1Lvok6lO3nnioen3a0QeAPIDiy4Ob0Zno1v2zpLfAq5JoZWplK744
uDMcuMaQt23ldqln5LdEg8JXVZwOQcGeuGFXYvrg3ptOyWK53u6qcZGb9FsTpoxb
ULAi7u/N/OwZgdzKqscmAqGH59nLTXR2qhh9XUJA+r+qELAc9ApkfmdYPDKwq+wC
OTksD7aSkvESjTSwb2gA7cRvq9S6hnCNckiw5Hp7noBJW9qnVmJ4OYDDG7//Yxp9
NtNfAegLZQx68lprg2SWCyK6DT8EPpAK8jK2It3hLODX9lP+XD1ioFNobESVtSog
b2SXtZKoU+Wsid1LUfQ3KhZI9wHwWJhiJ+V8c6tumw0gpJvYFFwIHKIDvObBTzlm
8V8J84b8xXFqB8CVz+V2Bzic3gO1pms27kHE22I/v/45n7lnO6N6lt93DLculur7
aC2s36aW+SD19LBA+VNb+6kz2dA0i65ilol1YlzylsrGPwJhmLEf9fnUQ6qJDBDt
HAPxWcxjBFLCmE7JPk7DzW0i577jR77TAX6Lrj0Mw6vA66nBTf1jOkz+kGs4usqY
HHJK/Xg3P6nlWmtskcoe4l4M3PqxMW1OTlTwL187gagutEs+lMxedEXtSihBQDIp
Erxw3inl8YdTNUPq1XVPh9Egg84z7qjgeE0qALsfOe1JU18lrKFe0wsft16iSBKw
diaewEuY7cgO38HzA1JdXC2MnFgFdQkxoZCScvHqCCWyQasz9MlxQjtHg+qtjqXa
IX9jgAnzalBzh10bMtyehCVsHQqIZtQh3y4oyN2WiG9uZs0H48tZ+h1ie1MWu/79
E010jTfdqDu7cdVl6g/ja/rpysgVXSbitBqy+TVMYK28+BBrEwY+m8TWWRmFxhoK
nJsu7ajNUNLGqPmzZQ3xSK7+bgioypYfjuCMS3ITUJ7N0hsLDlas9Dn0wM3tTr8Z
fm8zMv47Y/OYGSdI4v0TtZabbE6wvs9anfIR+wMvOTR+P2XgWri2Znv4Zb05iOnz
pgLYWGJXOBk2FhmtmPJASOSq7qfRNrPHQxcW8NS9PUOzJZGNmW9Av9wz8Ayegt2w
2/aIlCENQ7h1MXX5zSgNKwo+oD2vbIrX0fsNBx3qb9kbLRhLgRFIDzRvdj0FpQP5
xRzR+lxD5X8iZkuQ4W+EC9rFucFejIwxMqj6YdSJkxp4S9oGi8/FkxHOOql/7Hj4
4u97ar6WFm24CKdGiLyK0I5bRvQk7CjYYHWHIyUtyMgbbPI6FGJro359WmJ13EgI
0WgRLMINkF7YtLxdsaEjDHEjKGSjIxzplbVIGOH8KPkOpDhGmpY1uQV//3w67Fic
sMI81i78FYwP1OempPx/zfxt8RidWB6KlPLYCjUp/DEwswXxCYz0yWFoYL56Cknq
dNeuKhYSL7FHBwBcTzCpKjuHoYEJu2zb3Fwp1QM2bJG+KRTNK1oVjUAv+q7x9KN2
+/qFN8mTTGMpFel5JUJEU430aRIRDV9AcL6MMFLXeSkz+tjiTgdVw4QxGbsbIh1S
eTisOUfc3rtXPGZvcxsie5k8wUwwkjPVuvMtxsq6zlP/PD7ceZRE3kbNf1YMfyV/
2QL0k4GQTSQiSDO+7KB6nXg0rWSmEKAEnYsM+o2b3lKB7bpADct3o0/YHxVx+geJ
pP938IlH2xvHnPVJdRSG+W3oK3Yx2XOxqGifkGYk7lJO4M8UL2A8lHoRenQR0PVC
aQs/JJjI51exPKOHmRBjBHeO3veXWopqFKYssvbeuufPlbxTLkXvDmf1VIBo6UpL
rDlEDgP6OQ2c0VBzQp7MOpZ0eE5QWcVuEzQeyS8N/KG1NQAtyhDz8SBx1hTIm6fq
oi4x5xnOJcl7njaQG144Gt6s7N6c3JP78IKDqJ0D0HNk0qPA6kgiJ9qjCvWIrOIl
ydkjeun9+dOJYTB2ym/eHmzNthI3qMSRTBNH/QjRkxpRKWr6K9G2W02GfBOzkInO
qo9jX3bLAH+7OT+N+jGbwBe5F7Xl9+Co9Iqo2F2vBl6opUk1UtTS6qyhygX0qKkA
pDfIcp1DtysZnFYr8a24LObSqvDE3/Zs8mfLZJ0XIdoXh0OT6UuPjRuP176QaJLj
XMw0fvGyUyQ6sCo1/+gMM4W8pkHMPS4rBrFku6TPAFB6wg89FB0oeC9VVVZSGvkV
LkUHh+49LC7pR236A4XYPqWgyYN1WCADkeiJHlI+yd4vzWvJy1zQ/9nxBZkjVttI
pvd2nUpjQ9xSc2WcSFBEa7wOoPGUl8Y4LWc0w6P86vu7cbLYgCNPvOwEQrFEbruE
0R35GpzE5L0bj535+RKTnuTwU4CpzwEOOkhhmLs3TGtPd/Ox6L+6ghdDqTkIIssq
yh6RWAZGIYdLlrCjmZvFhE7t+51ZbZSC1F995/LnH/2LqLgU5irZ5jusKdu0sUlk
ob8usP4FsrgKR6aLG2W2s983RYN+9NKKcnKxW0aCvK4pikm9KIWVnFJjBHH5dMOI
FgkBm86VjSzAspcJ6tFr+2AwxZOAb0SK+97KIMrZKwygpCU/myYG5u+zdVYqFlo3
KS4xK/2JLRqs18PTljGLrzQkyEX+1N3XWLJJkKAGEvfPK7ShP6zyQWB6+lCGJiWK
7n4zI1TTcd7qXgo2NT9MmLOf3XRXYyuolX7z46a8K+K5uPCO52u7j7sRhui3/7tx
p5kgBV45cQkMDVhVLUvGbvzk/RSsiCN8FgupRMLL6WloP0LJmg8BWdG8bQ7lTagj
tIharVHGGZNujTWftOWPcS542dkMoV3HyJeADC2PCO+rSO12TVN8PX4jDh7AXFzf
0h9GTzdQagl13jk9GT4t3O3y2Srs0IZ3tT4HGoRSUkYhXow1NSFeVhv/jXyGojKw
ltnaeP8jsAR7xnyp5MpMGRUyWWclDyVGsc0dro6GrwFQO0gaC/+3WCigcZkIiWOK
kOKX71txKFVcDq/1AaI8PS7WG92Z2oYCZjl/p6x9GbdGUIZdFKM23PSOzsx19b6c
RDaN+sZM13qR9DdKRKxqKKk4ucXLsBK2v8JJw0esyoNmXcPXu9VC4Ur3JYRFBzX3
bAPbYtvSZWeGCIQitYH4AK6BSCopdf20mfIL9r6F8RKIDErmnNar1pflXbAxEyE7
NnTZG3PXCiFN+zTyy8z5Q6NdUrpHcutTAMN4qtbUx3z27YVdYY/VzMR+3TSC9XEY
LTGdbkeDnYgr/l49paUXxNHL0wBEceRsmrizQ2wdJ+JveByn4vCGATDVTuKjsmmF
5x/BkSDegiuvGk0bNJSccBDJiwez6fFyJn7+N9FpbvzSwuZ/+0pUV1hSsA/92DeP
1Mif3TchRyKb8NZZth996abv/76iBJ/WgCu1+YSa11lL9/lyW0AGuuLt/I8VHVsk
DxBaXPBxxxyFE33XBy+keh+AdXG8jwuzCokKjZN4PUx79JxYjL0f1Vfr4VZ9WDRP
WTD9mkzuwUPEDxq2Stphq58YN3dm+gPtq2IpcwF3xzY9lCIih0FnEZYh8Zlbn4ab
Kb4GdXeuUlOgplkwP+s6z524g6fBccE1pvWtul7y+4kixGM4uH49KI7r9ysR9Ief
3NqoIyUKNsFCzEId4ZdUnjosCTRBHzKOcTcvf5AJKCTyY3L2ERlOU5Hv4Tx9JH3b
OCRp4u8ypnq6KTMTkQ1E02gbn2/yqelfq/GM9ia+coYYH38IMf9MWmhBdA6QQleB
JkWdgJ8WL+44wzq0Q+zmwWdvA0uvQdOAXZlYTNaNFI9TxRD30r1yxu+DUDcLDSOf
pGhH3qMMfyFPYGNTO3urq1jHjFVtCintBthF8ENG46lt0spK0TqfjpPbezTdnNUd
uPd/ARt9UQMINBgBAhVrBKeyX+Zj9lqNSOr/mrc5O0F34PK7ukaQ0jQTox4uWl/0
wpneYfWgz5ki+ggrdvEi7ziJibxx/AaMcpZbM367MjfgDWgZWLdbNgNDR/LkAs0y
S+TbfSrJbzNtOo1n4AOMyuid+/GducqOMeCcNNYFzvA8BdLq2TggKeduipqChhWd
SHIJ5XbMwF5ZO4Q1lWEwDhbd2vahjIla7I9QYkpEaXcpnLgPqBiOKlDeIt3cpD76
X/WDDh7vCaqjqu/N/fXytQcu4x7QImfrIWt6sGBUxrZXUct3np2EiskLESY4/LkH
/xxMl79+YdDl+BnuhxHOb3VkQWQCX4j7ANBbqqZtPz47uNVU19hSZOb9mWfYEB1x
0j3oHagYn9fl1OAYTshAVGYewy2NJP/zzsYPFDqx0OJbAGrGwRsDlvpTG7phZScH
sP6odmmCftSsk1vyxhUT7d15Qk17+k6F/Kmpdkc6OcVSvcmLSfZDwmNyVy/mU52N
iHUmK9pyvViBHQyZFbCN/cW7Rggsw5Ix8vm/79CEazFboTvK6djWawBB0Nc2EDF7
8ey19lQF6VeS08zvKFk3WyZbas6Z9ENhu06tfXtwRY4thGUBTb5fy+IUCREYeMiW
94zWJvSptjnUkEigPocNXSw39HRI+IBgMII0Rexrb+wkRxwyFyKGEQkMectYFsWQ
/MWE04gnqDP+G6Uj1o//v2/Q5axQnfHM22RDFtXAbt43OKMVFxgU/wIbyLiepYJe
oXQghaO0rdo6xvjP8C7NoT35G4ZDoYFxapyEwu7Io/qO9XmaAtH4l4k6bmiHTEba
3bTZdIysW2lF9CpWj7bNL2kV/hqN3UbS8TXU/ZpA5vuaVTZG3LfwYW8ngoaGbA3i
NBDOHIFZ7Yzwsref9P6T1ArT54aTj9Tqu7vE6uCzxm5u4ry6Xg+hR1h9J1wpnLmy
mR+dQGTQwMWrHHMMibK2tfB5wMYwVNtIWFCZl6rcT5mLgftUVLufCo0Q10v9fyU6
2U6P20GBAwxp6M4njLg2sYH1AMnUlAxXncgp2m+zuYyU/JHPDao+EcdRwNl3TdcG
MmiDc8pE9FT4By4evGLG+GtFx4VJs0/+n001xRa8GsF7busN2O++utdj3WQyTbBb
7k39SBy/RpD5hpRonK0LDISmZE2EBxcEHOuQIK9DnapAdWTe4jTSQu38yjs9verO
wvoLAuH8N8EIjxcbEfgyKD0Af/yNg9GOJzX3fH6TYQ75YkJP4kuQFggdgmJYBUL6
599lUJ1ufnzk9QaWalbIrQqhcjsi8qP1vE5BzUNdAQLGVbY9RHuwKUrPyNF26Xg3
X6U6SBm6U0SffBJ3pVOERcMAAU3UtWFIcy2bLOLrY84iVaAGuLQVZ6BqdlW6S6eW
zsyfI98jENlGf+5Ppoj+aaA6AVW82ieBOUrOTEMPWSR5utEpix0AbYxdD1aPwl4I
bumH/o8qUw3E7TfMYFTgmzWwEWYjyRvXcwLCZnmMLr7TUi0qZ/GL7+ALfGeZc+Tn
+WY1VXdfdf7F0yUeGHP2NxFhoT/V46bYxqOSwJzWpYdCLPhxlpPmr5cncmSTuhQ1
bl7uwuExiVA2ljM2KQo0j3/8Cwq5auQgRi2HWYc8lLV6G2C7/Eo/JS5VtVGDOcOK
A3tKwkDg4pg6+pKXjGauZbCKT3YQdOHbaeCoSeRIOygkuyskWXQhVvsSV39W9emq
9/iPC9S57L+C0bJZlwQbMFbEp1uNyg1xOGWTR+ol44wuBzQsP2k8ZV8+JLxGEBc7
e3aB1V/WhzLhpz6LBZ/6imix0fwbQfCS8U6gqSq7DkY7v5mwf3uNtY6RVBjspmzv
zv3i2dUFjjl50Yumacx7No+qWBxdK+fpqCznPq4mQO18UCeVLAn2fteKZF3hYDhi
+s6NTDmGgTIYPDEPBZF2zcCmrYrJRVKb6gxWuwi3eA76QnKp2xDjmI+D6oOR7E4B
QOuUHxno4WJQs2EZqZuK1hURpp3fxBpNSPoebcAxmKHTRGbivF3hwuGI5u2LNvYh
sLUGzbFhN3qZVU87BqODdHXhw7cEZ6GCeBWtJK+lH13wfdKZeYRFPH55I2D8r0yW
2Vldb2CeL0KUKwWrk8C7+3orkSv7WSOiqNiKF8hZeR+3ERRrWWl7luGta5ZsdlBY
YiHPccbwCR/wkKvOciTq0FN1W5AXs8YJlN8/xwphzrrImoB4i4jsdXpFL1puJDGf
INFssJce1DtO1J7Sa9Sq+YN1yL14kHCmQy7SXGKcyPjsvyo6uIjTA4wcwhCKl0wC
aGseAVgPwTfDTUfTZtZw5YmgFQ6gwD/jbJnE/GyrizBF3ljTdkEcVvHwEvQiiZan
LHLmm/Yu4zjch6cnf35OtTDApGSXttLKcgET3eb3GgifYWtwTkjRRePFRHA6Nle5
DBYhNNZUB9sppJHVpO+eErk4igdM7qmeV8b3ceJIvFq8UnOvTlPAOKXVdc8laLtS
UmhTcLaXOwLJGSu3bzTRwbXMSyVqlZT0KNr4Yx9yt0j2F1pU9feQ6Vm4k20va5Ce
vvVNVx7DXnQvufCzHwF++y7rUOZlICBiQfCIZIMA4uEjtq3sQY3Tv7DoGN3grLSo
h+4DYP9oGo7Bm1oPzJJRBflZKHzrokEq97c5woz4TXkWOsar4pit5wGTerbpKKyY
KL0bEOq+AN35L/9KP9FvPSggmjlR8q+2/bQzbhd+p6MEpFBQ0H4ZttljJOVqXz7y
63nu2GzwlYdTMy472pmzbdE9JogK6JyvtLEDK2bhXdDAySVOgiq1xSJvSOjhVN1n
KF72mbs73+dNyHViLzED95iddR3bVdsswoCFvJD9BD3j9aHHYgilih/ixdlC963X
X4ZtSXgxOzIb+NMSJnV1aaMYogVvrVsRtG43L6FpZYaKzDc6ek4dymXR2NS62L2j
826OZ88g6tIBnR3zY5h2g9kpZ0HdkpqPXOiXN70NhLTMIkMe02JjCEzUZYas9rJZ
TTukzrXFeL3lzPAWBdy8ABSadNkHFCVnxo2t5eP0/ov2TPEF2JivQr2gP9FT/0T6
VKaZO2cQ4sPHhMre6bjGgHPKt5l+3oogfD1kNV/mBfLcOZQhWo8bwU+hobRFFICd
qfLq9Wvc4yXJR+H4S4RLcPxlBdJNmZxd11cD1PesIlqXn6y+Mi2XCEz5/TwzIi4m
62kdTRCU0pHpkSPT1VOn0Cph0/9nMvnFo4nV+Duka/dmH+wiTsJvBMVGXXaUbCgV
n5yaYb+eZq1ysimYYdP+VJz03DwEf5v08Y6qXxD/2kX+bWP2ZLm4zwA7wkVti+u+
6h8jjqFmNBepezL7aFyas6jn5lDAaoDBD7nGaaHhjAExTjA3wOF7zRyySuRwhwk2
cznIcQ7paIDZQQMa5K+PjhsRwN8sCjHrIw0r8gWepUntowVa/BpsgOQwuHR7EpP8
iMN8QPMFRlBsr0wJVhaPuQ0iBW0/Hqhx4eSL+/v78grvLXSurz+C/3/7ENS3PZvC
XyC6DK/mP8jdAwFuFBoXziDiU+gHW5rUthcxOm+VE6e6tBv2A3rPR7ZrcayFxOva
OugptwQObge8cGPCm8afM8cxGSTAiyoNqc2ApkCwFmCjR+759XdHkripLIX6pNiu
YtOZZ4X8dwjhE1s/c4z0T7LI+nZvNGaim23SN/atpa2b/vPm9NWQfFJCG99i943m
aSOCNF0R4iP+0MticrFAWmtqXwNLNNMI4kbjN814cW80wSaRe4IeRBLxLCvw/j6X
7yF6UX3DMbTrAJyjFj0z/qEloPrfMMkqVwTKvlsfs8gWi8p/rzkTbTsUzUP7pz2Y
CFYN/0Gefpeynw3JhKTYL8xj7VBQeF/qI7p+7OFB5eopn4gI/tkvk15uYnsIUfOX
VEYZ5Pc/AZMoFdpBzqlaSoajB3MiCOt0m8uZMW8Bw+oIVTrlnWhGolhQsqeoI3d7
PJhlo+hAu1TfH5xs/coIHHg5DmAo5eyuwbsq3QMfe2xIBbEDed3ptjJseujdtBAo
DblXLAiQBQGtKh8C8I1NSmcDMBJy5OfSWxd8WjBIHWElyTVltA7T+ttMPkbbBUqa
fBKf8K14ZDMe8sOG2dM6iB6YrbaV5E75caA75m/E0FIaFvP1K66bQo8tIMjYtDI9
Rwscw4wpUgbdr80Ik57e8x0qWod0vtbkluKEIUGbJpRlfn7/jyYX66JnrHvKfhYf
aAd7xmNr06V/tp9nfhi3mcEIJTogBs0qPLMUiJv1m4jKcP22xMdJwkz8+D5pcnfw
dL8PTTjL3IJc6ouz7cQU63m12MAzakTO7lRjHlur7gbvNWoTrz1wsiJS9m/T1l2j
2uUhFHtwowxCXb1O8beKiPaGGFCT9aZPU6XOFGstSXfaS32I0f8bYlGu2PTKmXWj
apsTJ5iwnARwzD4jlac08rD4KhIDgxpessPb7wbywRcy2gZtxakSUguhY6VB7T4W
idie76GzRdJPJmBS1kLtWDKx7vQ9XpApcKOdS4mcdUEyU9XXUwpoZASTLvxWclD8
soVcbZdHPACYHc5wVMXaAS15bS3bWOn7RMN8n5HxEFE3W0OtPq+oMDdcS83aJjSF
yvzkzc4FAnUYTPvIW5L5IEECT5fzTWYjq2bRRQWxzmmUkW+nwWHtTmReO6FoQXhf
p7HYSXbLFljEEkUCef0y/tDSzbrdSEK1HyW0n2i12rFcMAB46swdw25az0lbKFx6
GL6Qc5T6sSs6FHRP0i6WB3VUakoRmzUZx449JyYyehd0FgugW5qa6hhN91yfQymX
BltWKKalu5WPKqNNjXAzLKgoV9X3a6W4kJ3iCqvHY6QAYk9ZHbNR19v4JGlYrFZ4
RwZ3i3uToweXUJyw8N686wPfYr5Sj8DqiRXs2mPG2HHoazRDGy32d2UkYhMvrgQN
lDM9PiboJlKxZMpKeo9TZzlnBKMGcmMa0cR4ClZ5gEGOJgBIKLDKoJWzsb92ywMC
GQdXvgCdN7svxkGY56q8udruxBCgzc6x+5IR++7oBhOrRc0Qya08ODxuiGF81BbC
5a29D5osFsInAxpbVSTtuL/02luR4PU7NlrXe7VkP82qEGI6sj//BIWk6XgxCbfC
Qave4T7YJQr2JJdqTgpCFGaf6qFDFm6RfovyvILusdHv/I12e1A0d+CmCFzxE9uu
rNCcSkLSKLZMon7Rjd0PzPUstyJWWfSsysRBPOoSUcaVTRJ4s0n3/zjDV0aTiSsE
n3YUxQ5R8BbU9fjR6H8XutdsEFL2QzodEXrHoEr9oRyZ+xieGOxUQBtM+a23gFkg
BZCgyMKKoQST4+4rZb5F5+vfd4z880KKg4Gp3B/kejahgncxg+3aQRnzNmbZ6v2d
zNQCxrTSbMjNWyqv/+EZkXAIsIovCYGvvOf3iwpcgGVH5i1EQfIOwhg5zWcvChUC
SHUZOz1xhUi93xFBnpsKmmBZRFIMcWevl0pplqewGUxeOq5Z4RRri0FBaPG32wCa
Z0gXMw0AsoQuUS1ODnVpcSThkNWorBb4d6KFEBXyKhEjHrot1sz7GxYkqsDxluVN
wzrT2VkdjMaeUl4EWyfi1j/APDppfPSVqJBOhEf8Zv0mOR/Ln7tOnZLEGPz2Trce
A05LF9VbLvEE6jJKgS3gevKeQWYhhG1sidTh/+jB7ZoplvyDJM7Q7ZKZjaAgYGZV
kIG8tUY0JPO9CIIgtAD6/SvQCY/EMwxEZrgCVsMJIVVnis8ReyHIiZ1RZut3hJcN
n+FwSItwxaRh/UPdDUgRptmTnZ9WVybpVlpBk2ygBLPMSaNmG+D/68YT0VyVsry5
j+1NGjuCz4A6MZpRKO41kwUjsVCPg5OY+MeAzPOseR06bRXyCOU0krgr0NONF8aO
ABjqSAfbcTuhlt64Nnj1X4FJs3SsPSBiwC3wVlMEh9ZgV0kM2udtbHM/qJ1MAPlX
oTs8gUvckZVd6CNURgHjTAwQqSCWQqAR259VnUsOI80tVX/Qe2E2uwmQCuCmoXPy
juXpzcV0A/0Oj9AIiX6DuO1xzlPS3TTXLF+VwWrUStEEkFtpU9OeyS9vNtHxYuqP
tZvSs3IBv8KZrCSPb65Ina3DDQXrAuKoV+v8ux9u7RoMYckDqi6S/fmc8RoW1RPx
5EVu+B/i8i33LntoG/BQt2rykWj+0Ub9g+IXv/p3R2tZgZjLkNk4l4B937hlqJvi
jtkuQyP1yHV3ojPVPOLGx8VWq8VKsTk3vZWRhunxSxAlJ1nml/HBitGIUQ0d7DWu
jIu4SgYzA+2fUvr+8awrYUNhJbKpmScCil5zwqM3b/WwrqQLk955n1y9PX0nwTsq
IYp2IdR2Jge3yrELuBp3i1VbMNv7qFFzrNKuxyIkKAZDG12Q6UR7Iy2yRMD6XklA
Ri5I+CTtacbBhntzKKKYRgtuAXq9yIP44PvDHaouFlNYspxttvSX3AxDpZppp8jH
f1hj3v2KHjJjdwtyWwwM4GLV1TUu+K8UbOdRjAVTiZP/rXJvsnc2PZ3XmBCalonO
8H0a1wcrBVE7cZNEwJKjRIIRhdBzlPdC3eEiFNoxjv6vfOdJaR7UgfVxIC4FO90a
a+ub7vWTAVs4JVhP3kGdZHH8WA0A/TrdqvkpzSerqK5uY0xrBVRNB/Od3Fiq7kVr
IZ0aRFoEn+t7MzvX09r0QN9lhSflhJvNQ01FHeaBfKDPq5NT1GPaDLlb0g5DPt3P
t2hfRJmftjZeJk5gKozSNlntc37QZdMzKKpzYjYr2wIZA8eDZ6vczN5lIC7my5+X
qMUs4UFzPfePzu93F6vW6qE2RpGKunGL85ipSfjeYLx81giH60A9IQpxei6UkoKM
nTk5zykCOL8vGyqsIBZAdfe+Pf/OgwpF6763Mhwu6dygCOpJFLkoXExTrSqUUJEs
0MeHsXj+TwZC52ZJbxPoLkFrHqmqqY0MXUV4ZTPUlKOuachoR8YVvA5dLAFam3hC
cs24bztGrt5V7zpi3UYMhCammRFFVjUCvwdmfUsyKa80A3KdC/IV+tqsuC/QlCax
dy46eR48nJBE7/5u+4ApPWmHZ9o0XApXIWL2T3hNQqQH0B96RxSGRlDrzUbqvtH5
T+kFYIJq30kV32xkJ2SBTXAozQNYVWmfqGPE4vkdPNLHsFoqZxJWD79zm+OsQQbr
r2vViIk6r/eR7zesO0iH4cNxYz0y0oiemm6R60LmMpWLoV3Q3a3Q3bI9PzYUDnn0
SuQQhlKqoWo8o64T/LHxgLuNk8cUSTc1IiB9gG3W9C0EyTdZKD5jENGXyFoDjy2c
YIYQHandHBRbMRth4acyUJboa8u57AcSePBZOEq7H1JmGW06fDPOoC9xJs2wo3Go
KxjCmQdZ1sDDjUFT0VHAdLLrZzem+Y8UpN7fU/feSA+mnFIqnb3PNc4Vwr3u0kEm
xagAgxkXcQOpgbncVUCFoh3MuVvWmqUwSgduIMGW6cy/sYnDyrMou1FjN4u3pe/H
3yWbq4JXyG/BhCtVujpmu5QktGPNpPdIr2dCQZ5pXY0wIG8Cy3R41PwQU0oglDHd
Imf1PZo+y6HlW+FKWESMKm3WRAT399gL0fdtnzbgwaCNQruwtsYCWVR7h7J/+xZO
Xvlx25mxj5jjXBytHdsBWPHgd7xjYLw/TT4r2+i/gzncpL3YS8B2AHuHFUKGqZrT
bY5O0w1YZB0476NMdROdBymhZuI6C1pxtBMNdPuXZqdu4qTn/dJhjW5HUDU+UFEU
YNlY5fks/Lu8+D+Ul6W4mg8lzI01qRng0h2hHJAmK8Mp2GlCIittWxXQS03AwK54
5kTsr0WtLfgoLCfW911c6Jn6rDUbIgIVKnl2t6fHvGFqnPbhjmuYYXvlc7DUuSnD
Wdf0VNBHCoxETnkUS6ZAJDWbmlPjuS8cMV3dY1GF957+9ewwX/JKS7iZn9cQ3Fih
YYI1pufwCvk5TCp61vq+x9FxjGqgWbmfDwiGigtocR4D7pRRklGK35GN979tNdz6
PJNaxnhP4MSXzzynyYzy46g2kSY9k38oWKP8QhSIf1xR6DjzrLKQnF0pVcEG/0SF
MN90H5hfCBijToYqSSjcu9nRs9a6NrtIYGHD3/y7LPtCZgtAf9lvCL95hKb7WpyC
ejPsXZbrmejkryhQpclTEtxPwh7Crp7hrlVHdmeNBoYVR7CNAIsaK16v537p2eXr
VGh5iXPw5glKMHiECyhGMc1/Hd82qEWA5WO9TJguVglcD733AGpmcRn0rvQ4E7eT
eTFMw+onui4XEzcTlueNvHHpSOfmCbI/nUzB9zmSCPOikgqxEr+2ped6UIiCk/KY
CJehkvcDq6VmzxoBq0t/LOXS/ndkJs4xqeyBtQijOpqvszoc7rWeFbd4RdstplV5
vdmBoeEILhpBli7SfPZhzcRtcVN0X8imWazSU7dMvZ4gnYmnNEc13R1V6r6x57b4
ZdxMSUre20eTUWp0d5EyyqNg34KJjGn2O1Vu33GMtsZUmVm8urHRyIFietydy/3A
jbkttsmdYDSJX95JVqt6aQjYvgvnH/xz0+Z8nVfOYL7BS9KkuBsVLgvNxdYWUMLd
UNR2P0bOL6BFUu2mkZyvi/xF66KNMMfrYydIMPhQQYK1kPgys0Ye3/vrk4056Hdd
YmNOoGu3ksfJo+U/phnUrAyCO8rPThKpCSkz43X/dloh9NKdtzTo3B9fuzip5Fiw
LPNkI4uxe34AL+cd5RctCqd6cWpwTpqiygQcrodOPlVWyxRMqdK3EoM+FLTgmYhp
+aDWD7werZ9XMbdnIIbwD+NJGco7+12vT5C2Jm+H3ShGNO9TIgfzll4bDJcMis2L
Oc6fiOmhifpa2gCU/bpssNPfitr6AHJ7ph7mJRGBKk+wTFQBVsJikeFVO6e81tPn
aGMhriWQ7dkFhVSDv9kNkVIrAegC4ESIvuw5pw1jLVUHJ19lPLh5thSzX3ncmQZB
eSP3EyyAkLyc3maWf1gayeH6r6kqJDn4D652rM1C9L9IFsLUgmEvxgUeZNZ7Db3Q
kqibtVuIM+aXwIPTMjozf+3cbINMNZ2+yTOScnwvg8CCZKprX0x23TpqSaMY692G
jyBMOnbRY9PN70/8dmiUJFntd7d3cHgEaAtwtjng/JhxDaNkftRbD+IVnnqWFxix
w6FCQqLFLG4xYi0x/Y3f7xqGOS2NWi7r1lcS6hGra0QENStpWA0wkmg4dtoLJpyA
luGordiixFMiBBSZ9pXMo3AN25PkvSwizN4pyXdNsxAJsOi4WjKTzHndKmr6mOea
AxFM4FBQKTzz04W/+dH0GaKtl/XtP3deSqcnxsy45Or+/A0P0590nGtHX53peeO2
8JWKZBdPDlbDeCKtEtP1XeJr6QqwEnTeFMbKTBgH44tpD7hnZS5iHJDBRHCt9bfE
VI7utRJ7GZaNhttRFAT7qPI32oVxE9MKsH1MXYVjDQMNkNGoRrPpI2gwyVIU7A50
I0sC9QMUKfs3qwj9Zop7R4IyHCP9DFDQSbxypfPTSlIMhdfnEQJgDrXBLCJtjdxc
Tef+MA1vA+2bZglx2D/0r/NwP61royS+QnLyM1PUvXyvo3CqY2UG9mGwNEyhFuXD
ZfYW7FksfOf3GcDJo/c+6b90XCwAEpsjF0MFXDNd9NeYGVU5KWn1aD1r4PsAwjDF
q2o2/+bl/PMiWqW+m1oLAfPexGGCXjMR0bw298RMxfptz9lMqsrM7Rrhr/bmZX6V
+g+QJdOGKLayu3V6DmXCYvZUw7JoN8b04TosGnLTPq9TYKJWjs1RJjAaGCGyuFQa
/W3OqXllYOuUmSgScfrubmdT9ZqvTh0Cmi/oibeym8C5UukxMHT+E3g/q9ZU1yzJ
IR1FfR7TbeTBmxb6CQ4UJi4xwro258HDQOg9STwOHfDQOq4AWY09+L72s1vD48CO
wcnfC1DvXlSODStvOEmSh6317vhqc+JucG1hnVsOE0AeioWyvvH8ICkiW/eE90eG
F8Nlp1lm3dSZ+gPtKKMyXz4pueVXPy9Nb1hceepLww5La55xFJmewamoaExnOs9e
IdNVOYLJUkecfxWgCfLpzlw2PZWa0NmBXd8tItjaaWW98x5ZtcI+m384L8Y73ciQ
BluIGFE90b9bYsZH+bNDC04/OKgdfLI5uxQkuuOeCJkjozkGT5p2jtOICxuj0B0/
WDLd801Ht7OwtYi/UUdnp8KpbMpi8mIWiqiKb7EkYbUpuPoYmTJJCxKVkYtdw28r
KzjreBLWVmLQRTdCUR0pp1l8L4gxHBWOIOiBZ49jxwvsW9Ldk+I5TrrwElscv3pF
qODMMbc4KWRoUjzcxTfnt4YQPjkv4CtPyR8CG/mWvSx+nXzHNip2KzMfQiSHBqyI
cSUXXULnixxM4iUOxRFM2hlrNj7V7bZlB1UARhfn8pA/+1Gkg1YVxsJ2JqhudLcS
P6axGbKv2mt4fbeCVX/oB6xV7Z6h0FElrGVJ2aiFOKxd8rbCniev2L+jTSg7wBNP
mFQ2VyzKT38ssvO+JNXSN1fAK+ZydtlLZRg/4g4sDpTE4FqUYMeqI7Ih1KxHUBCp
rF1/x+li9R1jXoJDJ3LAH2atpEofC0HV4kAEedUQ3PYF6PvDg5LL2dJFUFWK73Kr
rgHW9Zk9of7A/OcYzvwpIkyq8Y9/xGVZTuMeXM9mKtTlfxWXrSfT01UxyEDaw8KF
9+Io24cVpCmnrwG8RWW3dWvUCJ8Yw5zdqUFqdw7yQDWJjIedyeIMJTPfJjRSlcfp
Pgm9apLOdML3DVqlq6u+K3KceSgEWQQBSa+sL2UfCJQOBZv+KPcuTOq/1N2ksHni
vJPhNluwzMW57o4Uv2P0h03KZ8F3VoSaBJYCwmoeiihn0O4MRt9mDoomdZk+Oa58
uxh5ab6tMHDaM9QNv2QCmhsf1KTe7ZbyZJajnU1akvB0UjaYNw1Mh2b/bAjCcX4r
gNyDP5u4NIU7ZRataGxzF+6N4NEEBbAq7LbCNGiDF4BbOaQH46mU2YragUCtleIY
0UQ/fOgYHNXaUrGAYGmrWxvb8w1G27uXNtxVV7RSqPXk8oAPTbsXQyS6LvAo2Iou
dg0jsHhf9EBT5OP3sreVhmVCULBuPi+zDPeEWA4/mctBcRNrmKAQR/xel+op8dDE
FjHGb02B7TU2gfePQ+gpqTh0TOu6a3xeJKBmSDNC1Uq/K1JNP9jQj4HiR8ayqtdf
Vtp+amFl9GjxhIoXjBCSDZGz/4zrrqYwyrKSa0LbOtpqdPi+hrEV2meXNNXnuDJ0
cceMeC47witRIcNvnmEwr8v9wLim1nAE+ZvO3fNMQMSUW6I7fybpDJh59TAINa/T
c6L21uxPBxj8usML3qKSxnyt+7tKyhoLK0N8ATnYjhncR7Fho3Z1nS3D+PjvJxOj
LiUJg4jmQxUaE0AIbEvp05qGGKOT4HKFrjM+dFJF9hRIS/whf72zKKpYxSXOlMIC
2tQEU/MtITkz3s7aZdmp1pk5nSC8c842dNwjfJC5fF9oxqgdl2NprnIwBJpTbcfa
9Y53oVIJxO5qbgl1zgo1XvxLaOBp3ltcsX7KENk8CuFW3Y6SV6ffKeFla8eM0Ar8
liR0lgtZLHWY9Kl8TUdVuLjdBw2iRSR/NVW85omMDXY2w7xkBvFQUVtsvWnlPo0P
HCRaKRFGkRVqqQB0KlrfJ0q2LUDb6KldbS0rGwajpE3Jd0HV7AlnjItzVA/hSt8f
ChBjqyltyZHZ9gw9hM+lhFITrmMZC+a4uQui/PIulXBH3MIp0d5bWqtAzYjbNXt6
uahxO+clgyegOJSX9SDQDf+n6vDlWJAtNu0++7M8134UwlkWLwU66yorvqZhkmEp
0tRyIJm2CztSyOoo1pOyc7V9gTpGNN6c54vESGNX1vX9kt8PU5IDjUnoxxoFQ6Pe
YiDNyQxXfSqI+luyDqFl855J0ncZh9zw2nv1Q3aJJfrFas3R7n7WHEkACGsQoDXQ
/qB9WZScQiT+g9aoamF1aMONi1fM9QuSQZNvlJbhXd3VWKNqd7mfKqQXuZ0osHoy
WHih0cdHQBYnceBfppM0QDTU7yxoKu3rUdmsPWofe8RidwraUDWZpeL1iToMnD58
t7JU8TapnH7KJpVsDDOsifjaCTZ2+y6zKtwQqtiPtGgoQ86F8BwrwXh8yTzwsCBj
LrZ+GVFEo78LoMqOTxE9NmvSJGf8gH1Dca9V2wn++Nc7JYsgpT8FA+pz4EXFK/gU
fO39V+/Df4G485p9YhP9REtQBJk/udUr/fMLvNPPnKpGzq/Lf5/59lZp20z+W5G4
vFZXnpfnv7PSSGk4YvNJnPi+zY4vxBxLBZVWEyCkXYDk8H4dbMtmqPHIvwjpVF76
+MG2t5QwKNebEm2MRRX+MEpEAi6m2CSbJ0lhFthg+eVeOrInYk8myTEreDw7uWCW
mmbT83PLrg1HFdH+leSPStckvgixfwtmgNw+FDDPlEJj92ALKxC0zWjZkeW1dSy5
lirxm8Mo+f7UpL6rFCxDjPhPe0D9Uz2oeCJS81g3oXvr1SZlQfOpcRepw5lgJbn3
q3of4vjTi79z7M1m8udf0XBFBs8KKikvXS008i4MGYq+4Y0wmHY3k/PUz7TaxFdO
DNwSglSL5SPT5HQ9C8iSuNrt9AdPJWOa0PELten4LVG2Qgfjm3biX8lG/whT2vgD
Don1quGzEBsqKNwn07XZI9Yxl7p7IdQjwLGo0lNIOtXsS3trR/a4SNCX2ulU/nEm
vaGT2FwKMcPEXcaeXjzJ2i4WZ/lVvwgTEPh97FMhW4E24GhdzRbTKYI2+hKHUxmu
yUWV53CkZ3oOMoFFXnzaLzFNrAZbPLTeHZa4lB0+3ebhh9EfX21hDn4EVkwHdZQV
teDY79ge8xv73cabLDARw2QGZLkzQHj1gyaV6VaXu5A2KZze/+Ha9ReZ219xx0M7
8aZA5kziXURfPFRPfZL8B0CA+Eg6DUckMCCon8Z20P46TRjMlZE2KTsKaBDWLJ+d
rH1TAfZaAkr6Xou/P/bvusPEJZSq3Mra2egGqEE32RGaexQd/o8flEHk1YphTJqk
11mHiKcoTkAuZJjDkWLNEkYlA3BfZoTQQs1bS+w3Fd5fhiIFOqyJmFL5YT+F/P8Y
0PiLQ5Vi8ljRWNFJ4HB0dkgZ3CaPdumXn20O8G74I+ges91iuwBmX3G7cG7kxUIy
0yOI1SfTaGIvrOX5xoLJadD9yAzSf1f/yIycVKVqHxtFYqVvuCovNm/y2TMiRVn6
AYz7kZQcoFEYBe+66FNryY2Ae//xs/NzjVYo5jLfDDG+z9RRkVxKKKsaw3IXryVU
DdsLJCHINWC1mKYQjSxMfR0q4W+ZUwUHlqMd864D/MuUAfCPYvV5Ta8S4gQoiotV
MLe4FmNFwpKLv248gtlcxlNjwvgxnI+szz7XzsxfQwkO0oT9oQvAALJ5tMnbfoUY
QTjwASjA3r3dqaZORYhWGSFhRmFi6sMQpvUctxSasM7ZZkiCh5IxD5YiN0k8dNmD
xFmhFerZNdzJki+stNYV+/IcrakWL6H7cnGE3yqXWxHHag3NsifvIKyuNRo068Ga
EsKZYBZhelbkY3FxRDxbiPAazPli/XsEY+Z2B7rPiJ9SmJ0PPrO0HETdwuCLrkFI
dB+PpRbFOMEC3fRfQgBK/VBEfB1hxn2d6noFuWsJuY4iEq6sajRMvIDS46hvVHlj
oEPewBSUvEkQPJW0i8MTDAtE+f0LrBJ/Spu8hnRSeHbyGgxhk+NSDx/oWe8EC6Ou
mEOZCsDR7aS2UQP+VFINX/9rd1bHUg/PGwCgq4yQiXzj9OuteoEvHTDJ7wv+NZKy
mRCBjfeNIVCErlVtX9XYmnOvXIrHZNkTLTJ4nEYTm9wtseqmWblWDEaEmPI1oDHt
5CQm7KX2+gZlIXslgbRd2xoy+6/559w7mc3TcBD23qLyZaS0KzzAsNwzxqgqySXN
gOfLyZlwDOmKL533k0yyIWDX6MPBmDqMJAVmel1RdgzFiKESlDeJkEwEKPbwi16W
NLYGIGCthGYTb5piFI3KxCW2O7grS4nxFA3JhRFL0lfGITmjPaYw1EyaVgjwqVuR
XEvPkde8aY9aDjmY01jv7U3uYct8cPOQhtBlO87RkOz5MVn3a6bIFR0FF0DU60g1
8u0oS2AdMMv1DwNwJ2We9r/u4N67yzwix8k628TN0METGsPIJA0X94aEetOnEt7e
lXKbB50YI0kHpGBbJgLuquA77hdrd8hBuN3Db+FXwTBeETj1iFjJbEOHHm43Wphc
vIzWdFzOZD/OzXc9tZ9NuJHRG3+Qdq/VXo0yDS8oQ4WOaW/RSKLXFPcWJezL/krg
AgFhioyaadevV8tVs7fJGGoQ35aD1ikHdXncHdNMgHlkTdXpDo8jPKbAT4BAQOBc
j3qe6r+1u8VMPz/DwvyA9HnBC0wvFtO+VxLOedSedF9VH64btF340wzEbSVnauWf
AVnsuugiXdWAEszmarqXUi/G99bbn9QmDrylWQeIiO5wt5Hiyobeouas/+V+xi36
FDQoNlbczfHHvAlRMjJXmfLVla0xVojUYZjlA1oj1Vf813alU+HhyrTU5mTeo19Z
kROA+IqHYe5+biGLhqtaacnEb3mDjXWwT+YOn8Unnhy3lCampUGGooqq2GjeHNpC
5AT0K8AQW1UhgifyPAfm43V2H6G0zKXgznPD+wbpANd+K8AeIaY7XIF08uxfFJPI
rnvGnAEBsvekRwE7LgbAWa62ToNgNr58al2yQ/d/ie9FH10X+daYFDMh+PD55syk
3xgAI188fGIw0/PXTkBLSh5yp2NAqsj/ee1tBqIxmJLU1tzdAyYYEToxGxueJyHQ
RqL563WqRD1oKq0bNy4prFxGdHYllsGvgCqSn3izsRXuhRKcQE1L0ggWOqJiAWNX
SL8p1xNofj2568+eVFbV0C22MrH7Le6dREnV6Rn1OxyCuRjQD0ki9eni5z/YGAnk
AaE12d4J+ktSGG7oZkww04GrrMlAw2hPV7luUVQG9TBvtbelVgKoqS+xI7OgeyQt
tlWyRsAltrkDlRM40hdcyfIQk4kZLC6NATFc4bLKa5tuGYxNnhI7Q3Wi2bYTif2s
fy+7yZF6xVct4k86ddvWEYHOrScPlUb/ycn9BIegbjtUFnfw+i+5gj/u0/pGBiIB
1GHHcjbMn7TVGFA5p4Ir+V1AWTz2hZdyocOZjZ/48P61d+Vsz0rZxCeolIhyNIjA
ojZeJgBw1AYrDAtP6mk9M/VHbq5Qte6nS3tXl5HqUaEbptba7wJ8mfwAXpL6VQrc
IRZMw2sfVYXUrEqA7Nj7dxMtkRqiUztMgDK5RzleKrMxqt/M0YvT3fZqZ6x5dCLX
asDcBSmhVOzpbivGOis+ZEEkTIWnfZzK0ovx0sRX1eTbcSqUExt184YiNoLmmcJb
tIBvIo4xVXZsoQZAKCsQnoLVM891b+agEAosiOzQ++YJYQigW9EVVkveXhQ/39lI
S/+w6hRPA2zFxUBOqsz30Lonuf9mhEtF98JbUEDThNGGY1YloNuym5cNrh/ihmHT
xmenDcEeaLOqv0t+urBWBF/uKThWluXYDlZPKHJSp1wSf9f7fO6Uj+LPxHOmnt+8
qxzbJMIxrQfjb2dBEN/8SkLHOyF2Bx0zmi+ahfvOkrKC3xxryB5QN15fRfs430r3
/filEu14FT5x5NbndqutWbywbFej0C6zSNOwU2VBXWn0Qm6VHBzqcIjLBJyjlSjz
QkExtc5yTQ8KgTafvDqAQigJ0+nK9tkbZOqvFwKCFRvE45VodTyyQ+g2xyxG7Foq
hnskH6MVDmfa0vmU7GBy9fTfYygOVgnqraSS8OvsNvQhvzVIpe3/BapuADnrV5nY
Ahiux/MicZHPYQGY1aSIi2r9YAPOw80FlhdQ/8aI1feK4nNoBV/4ZF2D9ykDtW2l
HQ73ZnDGFo7n2EJckiXEF06f3VIz2iJtNUAGEjS+aDQYYSTbo1zFBGtVHR2rns5h
XYnkklYenbE/yi98pGnS2fD0MFZV9QF1xUQ2iTi1sETrcjgeCqRjRCQU/z8ItAE+
WnRSfm84wfUNEvJC79DwoT09bCgWFoZhEd4EDpoo0I6Gm+ndrKnE4hXYAIEtzFu7
Vka23zR7sjRDPrGuJTHd06qENvsZp1kZqobD78oY5XD5xqnbRbej9D2p7592cRmL
etMxtYSoVD6cM/lpb34tvxI00TG3HFcrResPyTr1F7Phspm6ucMAuqI6WoF73T9c
rw6ZF+l9WliL0lG5vORroBzHJvvXpPszdHeODgLniM7A0j4JwBo0MlaE42tL0hQu
z5+CCpOif+HoFQeXG3coJ8b827TWrZ2/+uWf77Ur0oRxZ0UzjB6dYeFvVUIOIWh+
kZ4p9SgwrLvj/LYbYgOl8jdgWPwaJZf1ykFgy3exleppq2Eg1oAvQJGwphsUtW8d
7mv5s7iHheDFCa/ftjfSGFmFx6XYfC7RIsDztuHfn3/xr7KbAnbuPZ/Wu7SCpDR8
DiE7jPVeFBaM7xLxDo4bUNV0iuqAnvb408mgw0U/aEteU3Mxyn41x8Dt3SLDiB5i
GOFbPKHA7QOcu/OKtGqs1YrJw1dvuCWC5oDKPHUzqjeCunZoM1gHDsHedS1SQdik
LGHWmoHxNZLtvwToTl00FtKM6gJ/C8aJiQNU81bPdWpgolvheuSpcenO+ADoUaAh
okt4s40KuL+GZNCCMIWp9I/HNrPFzkcejgXST4KJ5hPrM7IWPn/U5ZX2SbwOWiy/
NgV/+hyJ7Ik1RSHWEQB/7Y0sGxous5b0xi8ki0BMneSelx8FZQ7zQ8mXyAyboV3z
1gY11z1Gbqj/f/CMlMU5AxCWgOMtOn7qrRpCBxyX4LadjOwlALGQh5owyA0EbWLs
wrRnHOL57UYPDu+IIINZVBTEybciOWF/nIoowKT0Oxo1A1wrGMhASdbDRxmDPtpB
gMjgHhnPOxyniCcmjJ6rgp/gCnu0yg37Pt5sdLYNQTUCqnXbdEAxR6B6Pb+tw+oE
T7HEraM1BaFNA0uAcoTssRnrB/qtgpEk8oXe5kvuVoDvJIwprs9neyHlfFI2Zmlk
ridEuqoVU5d6zplvvenaZEJ7MS9CwVkzywkNzWb8h2HoZiVN9PUzP89VMemY7lbn
2ybyoSAO+0XQo4I4qU4LU7miK/TwDCFSGUna8WiA0IxVI5I3tQuBQ0ZbD7lnUnI+
1zfatfogdArPaGl5erzAo51Wfiv1cdLwFs2qHVo/QH+xbPTSqboB9BpXI4gfJ03E
CCXCOFMQRGbrr22Y6fy8Di3auXE4YGKuNIXbG5Ba5LBo5HiFJEkj6EnykUUJoBX8
BdJ3s4fnQFXZZBpmqfJk6feJMxc4KpElRUcuwaAL+El1EHUz63dEF8Z+iR0DSLY5
fsboJRPT0WGjWdrZzFd0t4T0VFeKBOrKmGFn8l5nAXzyceWzxKRD24Ts6lgQBsGP
8KNSgqn109WX5TzFBioCcthACHWaMDbEimyv5B4VZWdgek5SaB5P3sMf2mWEsGdt
fIY65n24UAUcpLXtybUARTJ/LGVXiXGaroCcbr0IIJcKxvqxZtaJCSCQNBxPep6r
N1tVtYXkeYwS5SCrAIQk892yKpo+UTecQ6nLbyLiVGHM48etyECvUUA1ZNvXF3xH
obczFty4QZftbIEf3IcOtKO6c8YPo6Fs4xaTliHi2vtwpkC11+FHmm8njIjnWTem
Q36ivhP3iBiWGQSeIWQit4Zcwtkd84kt4ianUUcR6nF5L0Itq/tZ3S+LPSamJz64
Pibae8phC3BXK7SFEZ3opy1tFGFpCShU2u5wssZCangIb+zpV9F7vGq/J8633MxX
Ev/JTsXiNkXZx4r7YUrTS3BZLeDcfYCJIGJYFSab8yhNdjXTPy+ZJbBV/Y9D+o/b
kuK6q/I4bEjtWhk26TuSh/qFzrC7aGZaKNc+4T+o43bWFrzVldf9E08gRR6Rg08G
4M0kS2jceZI7VscPkZdof8kvbncHRgtCKAwuy/PklGRFx/exzScQKk61MtdX1GX9
Bx03zKpdyCnuI0zij6CKqmt8lL1KLIsWBzVvXRCsbVZPGJF1E89L1W8R+YZ4frFE
HvrHMPlMKjGxDQwGGxc22X2jEAG6zRLx6enI+x20FY8Br5oXX5TKHOUehiY5X28h
1SPSDJD6hBVxJBD8ylC1icdpuI6hZ6QFIsOkH18V3LcLrSLcUia1zCu5jfzQfDYa
LmMQgzI3dlk+zpEnz1OQm6kGcJ1ilhsROjsrGM1TF5fK8+1OFfBD1DOH2ExZYYec
1XQh+XIWEvULSbAxEGkgYFPrSWs3vxS9llOBFURaT1IBrlpKGt/KjwIJls8ttdYN
8jTKgKzqr0bUlDSOlvHZVgiAY0hl1xQVYgMUY4ui+qcS429HM2vulvDb7wa2BD2Z
aZOFMF7Fuq2TOjYcVMmpfEzT72swbFdmIbGv7Sd0ieIAs8nwmnPBrP3Wq2Fn2S10
TU7YS/E+/jBqygAGS+UIPnFRwUU6DFPlxXbGlFMk+2wdYd+K+/672Z6rkLkV311e
jmY90npDNIv66tLtxpbOgQujsMDvREtG0eHM2f115GPiEGAA1rBrwmgRz4VdQShl
37Az1KeA0RGC/7IebKde3kf0Q+Kl3cb1QlaLLzITLVagfS9gt9qJDTJL+yepWmKO
vcW6W7tWKxy1wJz1+VYa5r2nnuLpkH7w6dI74S2yUJ1+0sJK4ceIkpZa3BkqHzBK
cDnUe1eg0DNQMMQbgZ6vjsCQNy6K0W+5e4aUO2qJRM4Ra2hOk5MNYfL7lfzC6DJI
6iA1q3I1nZ2sG7jgWJ1a/T9lci3ceLrXn/V4cSfhCZGfOE+mKLFnEckKOr3QEBby
PUBTPjkXudDbIdbvhaE4a2Ttjm8ZGrNexUSGQlEsQ8+O50Hkm6C68W6TYwflMBGr
weiCYj+9qJcV2nupHv0N6tUwlAtbd7GBkheRS07ueqXL1m8bljDm3cXiRZlrAd4h
Bh0AoLuQufm7qnp+FkNP/DG90nFHuOnjKx0T7i+NrZn9y6Z03xCyklmhyX6mF/Tl
I+cTlgRHuYTyn3Bg4gK+y+7vStrhdmXcJN/T/rpjK023tuJUK0OHfdB7QYyoh1rT
TtHEagNvw6YLYLjbdO/J//7GDDhxGRfY2TUFNmdY56NZIJs2YITKbzzYDFFDTSU2
BlkhcJWBZeNcTzN2VOhW922toOiMlMCYEld8w8fOMJk20CGtGssh+PERvzbdtrNe
4LAKFy69Og6qKdksDfkcmR/VqbVfXE9itBvAHdWGEnietO/B8ZDU6Bjlz8Hi+rsU
FgW2Bd4tuMw9Y77tMvVMIZNMumdqaR8PGgeoDuohsfRrnnurIi/YGNt+5Lp6Ucm/
TUz/KXk5TjGOf5ZNgqvGXshaB99E5fTUWNE2BiMMB1RzWycFHndwTPygczECoeNa
C6P33u4jF7pT6zmTdmYIwGgEwhbrdHI9VKjNVETK4scxLnmFI3h0MwpxnASzHuMN
7+11o2WHR6RimaKzVo9synxdWOPxju4WVDV9jEPdaltL5TYpZM+cr1MsKYCk1FfR
FBptEcMvLybieu5/tpQoygK1BzOGHClRvZ7Pz6mve8dDOJjL2FF56900rUtfw+5R
ohQyGScjMgg9Z/nrg757dhbX/mSYZ2vXtvml03rGgi9OKstF2XAhPUqHg12HQ6ZH
n1GYGg2LrMwHo49eItHjDo8xYXGk4CyCxt2t2VvGXX/e3hgbyBwiI1D2Q0wefzDq
4rVODQw+JVwR1YI50XKdxDt6U/YA2uxpfzPZwyuVxisd4MMh0dkwERcpw3yQjabY
MMvIA8wbJkhI5KHDsd8WEf5gdSrmKavrUkrLRKNT16zn+jZiuC6E6bZvBqda0URr
F3aoF1ryems2kPXdAIBLbdlYe4m7uuWz8cVsh8bGAKItnN/2cIR8J/H5VI/vl6lv
XHpHWeGW4DyoJqDfeJUFbg/z2ULQ8IWjNKKD7lnOUC0sYtlOT07ItivjI4p7r8Gk
ZZ+F1at6ac/ms/NplxvgcBKu4hBQOKn6FOkMZ8sOMdX4A+vdIw3DjolIWRsYynUg
Ehz/oX2alqGdvrzhEXEDKrlGwpkIDBHS9G2qgIZIKNz6k6GKTCdBw/O6XJk+4W9U
pUU86hxa/09AXEp10ogu32aQOXrJMqGf3sR/cMgJLVOfZViC35oom2yZB1QZAUST
Vs4Fq9Qp9MNmbCYXdvSjdTzvP7bf/WDizVPrWX6vorAsEGNOIpac9G+8eKbLGv5x
V0lPXPFB8RpyleWG7ugoroRDMQOkHQ5QuNM/t7MmST9OD+pEh41fZQ4DuNriALi6
qi96VLIjtF77zkIMew65z3sEtrP5r/DcOGQ8brs7/t/DZ0YtlAmszgUfq0NvCwng
Pfov264/jN/F9mHwCVEI2lMNK5+K40dnxXzv5W+T9QwHP4s0dwgCIRjx3fqfZVux
auJenYcxOt1123jOsPXBi6UwPEOsIjUROa4d/9SUDrIxGbBacikUFbknz6PI8p6F
0GDyjv21b2aJs8BRmqzOKNdlkr7xSSpeVJFEbkusBM9Hh63r/jFAzy60w5kbQj5z
wpGY5HCYDYJ95HPm4dmCN7YmM8X/X+cvrbB92ScXp8J94acY1tYctrT9Oz1tgxEz
UUPtFyBIwFAZPVrPFwmHTEaozqoFIlM6r7ecXKrBX8R9cNr+juZ7a9774rDEcZ6N
Hr02n9wsOkN1ROv2mPA/4jv8WKiHWm0TK9KPhLQiH4cbPVWIFyPzDwMEqIP/PPoT
MNyUwjtLYn2LYKiiNMLaqPOiSGLZA3z7kJc2CuiX/qFualhd5Oo2NBoqUsHjHHOM
KdVChLClOV8Ofl2hvsdPTRAFG/nssMORDbMJ3tV7VJIdAq5sin0/FQfLnsgL12Br
4p/yQfVZspz3VsuYwn/TQZRAJlsmv1v1dQCDjhS6gB/J+UTJpFvJhc6O+6kEsw7w
EejBnm5j1OXsV8FEhLeY+sXpySlH2UK34KLhSGflief++3HpOo4LcrcxpMHKUpiw
X9L7h5aUadZjIVF0TobaRZBC4St8yj9jSyW7GQeYHaagA+f09L/twfSZl4sZF6bR
TBUsg/BwEGV543W3Uf9x1USTiUB+c8i5kkEz8IrAfhRVq2xcvAI0eaxCKOX6uCu1
PatpdPhmEsFXsGcCJEy9UmGJsRs25eoUcA1WmD7wDKy8PBTz5Z6NLi5a4GuBShlI
fhzXic3hrFPHJB8iqa9d6nFcsK0+qYyrQyWeOjByt9jR+WtnfSQwxQHST1qPHYLC
FiIn7ya9uEB6TXc+zYb27czlWTHIOND6QH8/RjvT4UK1bn6bWEBSrHSdbDk9EEcE
KSxcab4S/qmCNtcqzFGwWmTA8S9RXE77WO642kyWEst3l78jwyLuVS0POm09Wh+C
W4XPx64rH/V9mJbnjrLZbFZtNz+yEH4EbMn1pXQHIkmZGlTBf1zszcwYmfFy5mAV
ipiFhV3+ObGh1PnaYj9u5FfelMhYSKRx7BtoLUgoHb/ig8exsVFAP4Fe4/O4QDPb
RCAp38k6Oa3giwIjWSIjRN0zUVCiVVFXQuRB1HTwIeA37tiao5UaRIm1tdY7xYsE
Xx7TjApqsEKnYiqRvbAwdxJILpDJdxUvoStKFOb0FhOXKaiwbekbSdEniEBIZ76B
YRjQrglvPM/GsXnwOlv/nWhT1VOl00bYhFNoHIZULBjOZ8RwmnF+ml8hB6vnlm5F
Gtvs1WnWWBsDe4qagfGQpCspMETCG15o58d37O/yBmSPd+30fAQfbyfpbg1gUaAq
9iEP7nJPnsX3p/xpBb7jEqX4tsXUY+JN5JSrRNNbZGKaHZ6ggJA3MR8rL+nREHnX
YmyQxaDo4r3KdAsSG8c5096rXLepJs1ZBse+f53n8HhlZofifsuMT7zV+Isg3ZBc
BfAbGNcw/B7ubN+FTQAwdFrKdReXbVNErTNHOwLfHeQyYQeaXxIixT1jT+uGjqnY
BpDzAnhg1oYOK7sFyeuYfYjDs0h4PZRALkdWUyyuMjbhS1JerPEaozjgBOVZabX9
iiS0TEK5kPAMTML77jixFCm+Y3BRitpGp1kRC6+GMl4XtQCCy1q1S/z4z0hpX/Js
LHsaqnOX3P8RmaIYhvQ21SaA7lj/9MRPGzXyCvEzBPfVM/7awubqomaywB+c32XP
s5ijtw77DHBs60NGlYTnBSQU0DNgwD4ynsNLYusNXCOBAKZk38YvMbB0KozxrJlk
ql7NeHqkAlUVOp5YqAbE7qvQXjy6mu0PezuT2zzvAyR/XVOMbcRSWNGnv8mpDAGF
j3k6TnVCTay7zzsAn5GrfV4nn5lxGC+0f8L1kd0lcDhoYTJyJZJf+xtf46fatTFE
n4MfKO8ZDWWGDVowBDFrCjRPCgWoctrkYMirKd3fbhFzfRZcHRbp9VnvMST2j8eM
lL6PLYVa3TbOjI7S0hK+yWTrGJLwaQM+WVlMg6IwaZXRCVUWx4NoVxD1iBwweO9R
IWhjgFjB36Qs01RcPKmld46ewQIKHE/HVeARArHjctfg7FxJpf5vyu/+lZOrsdsQ
10JtAWF7ddvfoqaReuvjxNDmf3+ahNeF+9Tt+YztVYRfbR8hXD6Bvps6SKU+SoH4
vtFa38VoRqFA6tS5Vtai5rzzDeXr2qzfiMlltGx9JCftW5OhyA/eVxqeYot300Ls
iyRiqj33TH62mVHRpJzWyPYc3DcKQFW48AORBg56WCwPE2elL+4IBPLyM0LX28+B
/w7aPEnREEu/eD4CZuNhh03klAgItTNTZVef9BwPTp9Qv+FFGCTOE+V3qqrukeO9
uRg3Jreif65oyrYbZiLuQs1bApJvAArPXuc+Q7dRw52NXLnQkpDH3swAHSrMmCSs
LagSvymJ5qhMfT33ohEniBPjk8qJ1rTh4eMONVI/QA+L+3vyycqMqHj49fWPgJDc
L971kYJJvTIrjY6BdSZ5e1WFFnMdsiX4IroxM7i3dPJrlXSpA+Ix7LLTByMhdyYm
fM0IkJcaEZSkUQ6kEIBkeGnAS6SeABHA5XIjh1uUc+asQl5Yr9JbHaBUMpdEheRK
QE0YwB/9QTKXej1/qeOWPyhOEQAoT2dhDQefdQkYIRTPlSnxfvcokoVXwHpnUfgh
RyIOPKz0usZVoFWtMtIVy1TY/SmjuS5z0lisFPBq1ZPN8RLc1bGQXmpysNhhpGTS
4To2U5Kc6xSrj7SQLLGcMzWhrABjdIDGTiz1NCAa9dwBQnoBYON8W2grBGiWRE5h
d18V2B2lREopMpj8/I27xycEpOq9OlsypYr+rcp4zKJuns0HnQgtZ/ehQ2v3y76W
F4/M4yyKb+3WGyHQ8VGPIvY+LlsIYG9VhFOQCHXtXwARnQlShgC0ySueQQo12cM5
CUsP9WyFz+Di10rc0r99z84AQZyqzxuU/2ZLwCVl79hy2xdq6efPrzeQyLujrOK4
so5XGEoj9u/ZTbcCKFxBVdj0h0jwZiBszKKXMs42Xt3oa2mEpj19YIsYTrv8rBri
QKXxjTjDuMmpL4f/fivFI1558/4+65uVihBexMv7iNWn1twt7BqJpmpcS8v84cby
a8pvScQ5WIXDKMiF3wnr2ugc0CmMoGeY+D2NDroUH3rFaJS5xOVmxNVY/aYjA7U4
kPzZvRx1uk0ZSueJp+zrqo8IUdgC+0hM3HL7P+BO4929NR3sliPASxJmYm6t8zqu
LjARyHPf8fOgu2uxSeyyOpjbMO1Lsc/K+I4mnj3S0h5tNd+1bQBE4/4CAOmNDYRn
k+PVMEFe/Iizyu1k1E5yqqgDug2Tb/2s36Scj7zVWHfzceRPRGd6Nab0l7xi9x7T
TztmFhn4v7s8DdUm/Hafpyj3g9JwD7rmV0Bp+NZ4Q9U9aPuzKFISkYvYh79JkmE6
bs7suuwR0GTEZj05eIr71LN7Rl8xLz5oimqEaPW6L9XCikZ1uK4FxVXU4VM1Os6N
/GzmoDlqiJQHyzgND2Tz0IjSYdsz/Z//gf1+5jSYNcSVI9ni2J77YXSLBZj97iAs
rI2X+OXXCnyI+rAzWUIYygWd3BIvwWIk0z88vz0DqMse5D/X0nTdatAVGr10AYAw
f2GAr9HKZuzA/zN+Qr688dxYZc00hAagCRPdrm7tH9O5PhF69Ji7QSW+pORV6/t3
Sl3megpxFmfbTRJLKW0mwE8YMPSiwAFPJR0+j/Xhbj1OVNF62lHpiibSiPOs6oTY
w1fhcxSuvHSCVTKgRvr3sKnjT6SBu49R8RE6/mZt9hY33IEMTx2Q/uYfLQUk6iTp
/NVjeo9y3AMrFQv2N4wfKVfewDN/ncOiWZob4K1bsVgfxgx1ST70Qd6F+eVmk45A
ou4qKzwoNn7LOyFogL5B3C30W0wbWaNTTDFDmQsQeZclOYIKioCDAIS+wO6KCdqV
g9heXz7moThDD30yYoUSzZKkBUGZ3uw6douv68MzrbKbD9eQTw1py04awdRhI2lC
Oze2XKVxMYD6kmPLrZj65cSlBrBsbPpQ/zev2DQAT2F7BE3IeY3v8Uga8jFDPmEc
YzSErzp/upMoazmyLuHzukst8Yx+FrpVrkZkVMt6iYoQTszFimuAmQnFgftM3b/a
GGZ/sF0CPDNM7pivZBsoJhgy/9Bv1a2gHoMe2kEjpwLxW1CksODrk99PW3n0scEa
HtNqiIDxCvA3FPgT2RrzqTD23Cxmc2Yc3xqC4u+tYD0LSnNogCNOk+ZTwY4xTvmy
ZPwVF8LNOtNVjLNDXaKFnYtn5fFqP+f7XKBuDLatcnh2SDnSwnkP+/FcIIXxOopO
RcC9Eva5Dped+t8dps1lP4bq8x1JuTpp+y1JCq4Gn9crw/8+ObsR5tISA48W3OXi
+lpKnJxrYUwy3Vb/iqf/fHjRe7gOPW6QjU7cIwMMKwBPzLXd5cbXNL+d0VHHeDfZ
o+R1lNYQqwOG3Cre6i2OPuT5HdIYiXqsr9PWI9SBTX75eNyag8raYP7qhymVEm3E
MPlw8QklHL8xOnEj9I6nU79u+HSVi2h4BgwOhQo1QRVQtKVturfZuk/dvxYIXHhC
rEM2ipnGbTfZP+1gaXoO/3Z2eVxrKqc9LOk54qkanSJ/MQTf9YmPYvE88nf4LbQH
SYpL84QXAclY+offB6mU9o6OA7MM4A7bJMvloo3kZtxdcStfDVfvuShlj6fBGW3V
VpyTh9QgPW5yKSIewVaO8Mze4h6cvfzwNGIPpRQ22qOqDXGFLiE3ZgrRaOmBoaOv
rDtw2OjMET22W+/v+yXY2cA5yOx+h6XC06PL8/cn6i9naB2unrj23VMVIsx/9enB
RyJedHSImE9Md2QHVgRaSaQe8FOuxX9Wng3lxIhT1JLpg22962towA3uYrOkj9yF
j6BzOVsdkBtHWt2WGQBE+ql1OuvRdV0E1GOBAN1BRVEmEv0p0dpo94CboY5toZ5V
U1WIum0cmSv1VafiE35Oo9s31NaZzb29OpyHld9X+PByCgMdVRBEQhtGHZeknoCB
HawyRPl4/Vp3Ne0zhMA85+OV+194Kl9sWaApOPYsnR/vYCGmzKJpbviJtJJwU3EF
nSRJAUUJ+2lrm70VKcIK1+E4YQIuva7Wd4tKs3RrBx0YcHLT/rRvE7wW8BseM6jX
/sMEvGVmvCviY0g3hXUSmXTz36kC4gMo/M7QJkWS16O6lku1uVNbhZblNciss4Kk
zpTKMHAIvqUHq6qgBQGEdEFFszDw3Ft4J+M96PBmIOW3z98eZRytAUPi7MiKiDE2
GZ073nn3Cblydqqj+Tn/R7kNVjFK4bxla5Ims2oC8Ji3kQBpmf3mqx876wo8HpLa
uX0VnAfRlChA4EKC8KnV75nyEUu3gxofOYbh/XOpyJ3/+Uop4Jpz+wVmbUvuAAtt
pDyny52RgevSbatdijoabKEl1DBh+5G5OXX19fyBTlqGVprrFQSchsMHIXtVA6QD
mQa2Rag0WObEB+eiwy5hOapxbi8cKUFuAzv/OIeGy8DXX6cjPR4g6DNK2I+bbWzm
Be8DO5BIfKcoxA77HRe526sDmFNNmwa3KkTq50I18e1wnu2WcJ26c8pvQexBLsdw
wUvMf01+4iwmB7MgZ/1/t41xQ9Rm5XttCiUCWeBc7mImxOZYpcgkYpIoDxoIGiYr
reAwpjs5FFNnlc3rH4SNNK52EJhrJbkTPWgDGG42VQutGBF9/Xq7SATCUVol8YDg
ltIVEnYYWWLqplOtDoDr6RmYzJ8duvsFU46ddSpSVc6J9NXm8plcwttwNiLUvkin
/NWG1fi5UhnWKkjSN+AS7s+1aacaDbdWgmk6HFdyZEJPJ2oPksgwh7R1zdWQtacH
UG062uasyTzWaDr/f2hdI/HC1JDVJAPcDv7+lrVQvfSXQk6Us+1EtWU8n0d+di8n
2pUoIr/Aj+KjzSIJzg4JtW+v+frLmjDpe6DDhk9W3S0k36fwGk7xcUMk9GfZU+1g
wslSHYqp29UGgrrfgiX9FvrP6mO4kEJ+rHkk4bSWxM4K0bQfWpZ8KAStuepKxrgB
8785TNwYoYK3jp54Hn7doMFylOGwoyLAsOnNOPP9nNBFR/MU2FdLvHskUDGcbp0z
ABd+AJ0h1i2OFm/uUTCIIGg2M6YjE7ch+zgt9g2hO+axftXe+owF/ry3U9sHFsSG
wgvzcEtfAs19iuX0oJALDkiJp+dZmdBrtadjZjTKIZYoVfSmp2mEtj9erRY2JEgq
I6+am06h0wZML0DS5YBAxxyTpgayFUOjSqU/559ArFeovFur/9Qr43IdQ0fVMlnB
Z6S8FkJCWLXvTIBlp7Atlc5aVfUk7wrZnkMsnQ5TWTrql/BVtcFyEtIsbkmbRlwa
GFFkVw57CMEkB5+n4GG2pe6rrExihmF8217cGbh/wyYPEPaDBWkMe1Z4Xp7sRbtN
jD9mZmp+/paBSpJuofbI6thL6eW37oWElbc229Yei/VFUmV+OM66Xz5YPKNn3Fd1
tjdgSCPFfOV4/MIL+D/XNODcXxQVwPCV5CTNFGsuNsHyz3M8Lg/xBWoX+QjcckhE
YRNVpiccRRPwHTT7TEbhhdUYiID8QRRZ1lVP/Hmrhhg02cXQ1i3onQsbDb0zRrpr
/fw/P53uGUQ0T1aSLj9CNnqR/ZfF9Qw+IzGBMDMrv+M/0+MPVJOoY5MJdfJDj1/9
jZK5tfo2j1CxkqIxdBjXPWwKso5rpQwQOxPc7HNXFVSGI03nxCaaKF7bDWR7Haw0
DbAqwU36FMnuAwnW5z1VZPK3ZRFOIkSzRZtsA3QKKRX/Pv6f/0wzuOZHLQpBc5zC
U6Re9tUxi7UIi4+AiQ39vqZIdLmCpK7xYWvdN9zz0Guxq4nkwZSCDERC/N98vpj3
kMgSInXw4Em5ub+p66cZwrUSOAWMtTW6mWR5X14ZJKMbURdwJkbiPBcdgtkgmxO7
/lMYKOjXGgZaZTDWsRbFWcxsROF1RTwFAD/gAkKren9hUYebpDWrmrS+eZolRFzr
prG/JMMG2CMYRIUmZJMaF5uA86mUodaDBe5p9O9qhnNxj0TA9QOQ2lZnqh64mZr6
hyFj0dDmPXJIoHPcRo/kWK9uOtR0W0OnLBx+zpTbdfxN8YOlIcQfbK02X1LnY6ll
ZUvWzhNN8fdVaPsYmnaQIE9aIh6+9heWNUoPGSAJ0n6UoU4sDrV4sSOCr0F4uVJm
3G4FLpq3ZnN48Jbl42P/ljSRIhHC+tXqfEY22l6dcMZnCoZbO+IFY7RcDbruSSiw
xrPm0IDHoJFPH+UZHOGaaEwWBWWZUjj28ufQsWhvfC0ihUgLpVdcu1CW0I23yoYU
qPRM7wzwOejdED1H3lo9FNaBB5WeX5Te2mOlyD1zUmDXenRm/DOvwgCJEjSa1wuC
zG8gZSLXq5m7qJJ2bR++J053uJxZgLpDBmve7vs3OEb95eO7qpICVgXvn36kLQ0K
gRw4UgcPQSWQpGRvLGqvQKpL2K7dSxs5zwUmHdG72Ubkzx+DabPWPk6Pp08koZOp
P4iDnDYsYkvTazv9vQpSjRN/NFkTrdXaqfTxME17/FpOR8nVouBFMNP+V03W+l1L
KYunwTzVWM+bojUCwnQ5p95EDM3ZiT8k6z/SFjiTrNmeWQiTx+aS2z9x9UdeI6+O
QSPpoRdRWjdx5ojJQExNwGLvI2h1bB4yTHplHY2iNxOssxv3SSqm7iMBNhWcZ4/T
UADGhP126+rDAh+h6nsmhWmCU/OROBrHS8wu4YqRKqwQ6v35muy7W0oexaD2yIlu
KxRPMUMDRD8LkIdMCT94QNy7/rDCjEJlcAqMfoxJNQrRkltT5EWfUrUCbpFg6opv
52dFIymTDg1roBkQ/UtUxGCJieNXvF0+aJWNDyvU89qaZHHeKf4UlsPwSfitneVa
p2x18aKuJ0YDO7FwM1vyM7JaBXdM6JnqPiiOkg+qG/AjbUDSmtthCJEYg4qyca6n
hMDCp7UTqp/Wro62RiMnGGUMsouXEbYIe9UZEw9qBMZEjH234z5fhjcMxeOhKoy+
RWJEGq28HJEq+sZDQP1fSaZLsEk5YyfbwJxiXI2H4jbvJbu/Yl4spMmyAaG0CstZ
WFInqtSH7bao2pXmESHvwHpRw7hNxBEjnOJrNjsCtgC+bEczBQ0N2jlUoSDgxiZq
kikbdbvIIgZfj1aRxMeStnfk7aeFc4yuEi3P9PSIdlgQFuvmPl/ez1Z2VhZmf7ZG
5liQNPFL9aaC3lnj53l8hf4exBnyn1DkOzBCLve37HmNoCFRvleSmt87IqI+zNOY
x3xMHlRTgUWbRsnqn9QcycMf8oaGMUcRZ/BJECcACMAhy1KnLRcizfwUDPsfl/Fj
RkLJOsajamhdxrLlXqloIfMGf5omCtEyLBD8ZHyvAIvwbFO9U8WKQV9eCufGYS3+
5DQlfrVlD+5Rra65EReNjgLh7JmvnjU4r0T0sUovrq+pkuHpGEDcytcwgZ7Cp5Iv
XxgtzsyLhOBtKXjPZzTEMbQfSl3dLFPfBKC2tOmSA/6pjRDoyOuoaZ90pjdU/Lqi
ETxBKraaPEcRubwGx2nZJO3dz12lzOjFx1/TbxiGdCnI5FNr2mVlpndC3lfhoLML
9FiIGTpH7L95AskwGdJCVYlcfnMEdm5jZ2pfIsgwJ+xc0B8Rgd+UpUo/wBdXaR+u
OzYZ2ZlAiE6DOompYTkSEzeOi9kfofhiL8tQYXDLzwKcd5JNsvXSVPSi84+AzfYo
kr6uSnvG3fl845EFOE0yx+VsWqpLeJNEuLb7hoXcMUlWLLZ8RMjmL8Y5l5+NhwJK
n+/npCqIGhp0I+0cWTX+YYTGooExghtv1zv92ubFwV0BF5I8Z3Fen2ybQxUTXSsp
ODeIPuXM+hK354O03yGeUJqn8tYz6BzfxXUbpFI63ysaDJlv2R1wtP6lcaJSb+UB
RUpYRKgbXEdEau/4xC/PdB62uEwKebxsYqh5MkhppTormKv9cQm6sZ6VhiJXdf8t
bAPtmQlLeTANM1yJtoXcPd494afxpnjxpx8zX4N4wYZZPXuZYTNVS3I7N386rTup
kUO/BF+k1mhZHO8xBfIW5B7mt6WXeZLhuKbIkAt0WLIk+Q3s7cxFR6YhpMOyymnt
HFIOe5oJbmRFC4ZMvuqwkiwL7MvZqFB+l9+t24njsdRZVGBM++D2T/gJJmI8jEL2
nTy91HAcq5Z+wBki/ujeu2Go5be5jqw/tYDYTUM2Jd4LkB9yl//gUQwUuq9jNTVe
1FfigUsm6gFaJcATBxwtP1UUzMh7YBOWXThmAS+dp08njlNnjOWyvcd0y/1vg1lt
FxjSBLpy2efIw6E5UtnJ9NdkRCJv/RBxOjHBJ/EsErC7uGZWgZDad9JFiQpC97Sn
iOJ5PIyiS+d/CRv4Ns8Ng5cBy2EosdZR1Ljmn1wGSdORDJmPzlqAgHQTfJ4W0oOa
0kBlBanDVBH7zzEYSEH0JdIsH3JtgoBtazdyCgGB9ISNtnHfzK1Wn4FqIpPx44xI
vE5pdyAe2GmElgcApr/7xO0mxVPhKzudCCDPg0B64YBAVW0hz5XjDmmAYpWvIVdS
J0nNN6YKZ2Qw1eOpizHovodwLTy1xifS+CJ448aCKa0s+UNGWdLMiY2heV+TVk8x
c7XdvZw9Qjym5Dyro//gw5MNY/riIfL010NuBd+6onrS2nuhgfm+halCYymBmFFN
dgJ6hDkPphLV8ECMflfd6LK+U4cUREDTWFdc/zVdyibs5vFtnywf6GTqJhA4mSPc
osjP9SYNbGZzOd0Zl2YM3Ctj0jR+Fe5Czmfg7fv5Lovht7FQGR1pZxyrXwZFui0/
BsNgRnGoOpio3FkmtY3K5DRM8kpUrkh95Nofy53jfIZsT1lG6LmSMBr75H14ocVR
x3iPDMyhnjun98OcHPfj7Azir+CncZ0lxqgO1FToFvL5IwhM7xI357H1nN5ipHjO
Nt83x7q2PfLVrr8ASuj7D3AKNZPRAXC2oGxWdATsbvFXCKy5DNFt0mDtfD8eFHcs
NGXG0WqTJfskcOmHof4xwLmadd06Pu9hYysvUtuJ0LfVnMlkQDDNvGvFgWkWYxBk
w6PEBVlALOW2yd8ByoKCiQIk4QJ0NMFQk9tzbcwVdMYBtg8OZ7dxGQFs21EZsb1J
t+wiPmkFVeq2ql64xBmbMlCXfJxBuDkNfO5f1im4mRHfmQkGsJMhfvgssLUKDnop
2XFCfcqgCt8gVilAZwinVNA/BC270FRS6cvduzIloyWDJpGe+9hAHUdiohAovkye
seDS7mgyBX5ksoEtdztiNapxLmHkQ3r7n81aYrUIUYp8iXdPme+tsU42D3L+jj32
luoiKbrq0NvBEQnX/0HCRlg8VmniWlD97xQc02etQIuwEiR1OwZhdY0gkmvUcImL
z1/J8yHI09GYu/CoOxXgDnXD83nm5XCR9bnx66roOOH/HH5UpBl6wftMLcBpWhAC
nkQsCDRscXcoWi/bqK5R03Nl70FR5zmek53SmFgZqh0av2k+AzO5sSxYP71gru0q
c/PhI3cU1/3IxRkTZ3LQal+im4F6jiFFJH2EWNszrGSbz9YYWu/OmSHWTDC1PQR6
Mg4wziV1V+zZix9TKGkMmv/3VclynLi+E1OsUK9BkPaHzunK+oXkPz9SbsYSgHO+
UVVUKJAiLtf0qSCn6rknRXt96fka5PayjbZR7zLWvz9RWcY3FBrZERaQrl4677qd
BTDpGBw9r8b+Sjx/3se4631zh3ZEWSbEvxvcjhSzZMu4ARUd6iwQFOWguDmkpD3T
Lh3W1hAQHOi2cu4hpkM8YC82wbdHK0bV4MYQSF7NgYkrkPLukIx//JCyD0z0/g7G
XtelNkjgD2Y8nVwHlPyiWqwldOfAlMjOi3HNAvmRPRLBFsmqSPXm5LnfG6ucdCPq
3dsAu0lENwL1pE6dhwJRJjyjT0Sgv28QslhiyAfnPS5Pbihe4ItdnXW4cfFXpFZO
Qt/YfwCF3WUPUdv60KiZPXy2Xv2GkOZ6MZum/O0trmRZDP2OJ0ekbKtI747moiJM
9wb1v+5NjGp36PhUw8wtJfRccBKdufPcGXl6r5Tbc+Lnz9RYUbTNwyRLkVjbz5cP
a6sThGRwXoQkJPF6Ma0X5fO6FtA6+7ym1ufYgq7B54/jdSvN3Cnzj2CZPFJw8r5N
EUkdO+b0I4+0z8PXYGX68XjfzbQg8qotjycYv9vtHXyy/WoAgy2Hj+zNKf3n75Ac
HibVyYTIaOtll1XfLFVdYGeMuUfHqtjtDFC13ZHiMyi+5unC8rc3ZlEraY+5B2eT
yQg3/eTMa7K/FHworx5M9MIZKu6H+QJ3JXfk6cGMizGdiFUcR984tx9ox/xqrVru
xfEsTGpJTwBYcqU2ZBa5SQQCYwFCjaLeb+SgToR4RsLwPqreffKeRnxZ5xuRrSIl
LWyVZc8U43kNsZBFvl+/L/iaMsLgKKY5Q6mG8AGuKREgBhE2aExY+vxnzJq7xXq9
EtnXGju9wFr+LzFTs0z2tBS1SKUFBtQENsewZsCdHPN7qy0Blmbb3lILTD2CxcsP
fbFmhUGB+H72jMwMKxOvnEgDV+HKPVWubSVZmg7ySmHfPsxQHZztUoFFmqp6lV6N
Ci84zVjPOCd04avnLYUl1nUjzjbKKXldBgiEamDAbrQ6uw2yPWAqAYNn36UJRFeC
A5+e+rUgvZ7WP7rKkzsvOq7mbKVPk9QF8MPG3HxnIdh7Q6Mz8jYcgLEJ2rWWJj/W
MtnNYGtumIz4GIiYm0Lv0oMcedBUdKaf2A0/ruHcfF1wLJBwoG2zLCKPzU6ocrx0
kfpdiMdppKFYKLEtCiChgq/bYEl3C1XNY6VvizPpHiXUxMfA5m7EwRK8Z/Qdifl7
mHWpNBU/ieRcZOlZuovjIsLO3u/nr6XYfTxFc3XLhtB46YxXiBs9iqmvU3rgkir7
H0+k9ty7Wbh+4lr/4ZRysKa3F0gJHWZcEAn86ptNGDv7lZHit2rCXrr0SNs1n+T+
e/5oidL52RkIrhQmqAFAox6GqruUTh0zfe2+fmOSGdKNTpft23wCLrsvVaPPV/Ql
6P2OF/RDG7ZsYO06IGDVzk2sCemRqKn57669ny+UkOcv3MQTiRQ2sUz2edQm8B5G
qf43cOg1mNHAer3K82i89AYBkw7sm8woKBnW3AACaLp4mccTt+39K7H4fg555MLj
AodyXNVF7/sFhff2yzkyiPd9no7pzORgCHtYyHPjewaIp51TmzoUfERmOPY2c/gB
BitVKNNPzC3e+zagRlMvs1xi9k2unJX7qWdLDU1cpNFAp7kQCBGVRmQTMDZcG9NO
4P4lADobS++UaqsEp+xg2dgRnZ34JAdl/B3w0ZIRspOCbgO1YKsN9qb3ArPNjSxn
gOye8qzvSoYLNTXgQgRs1z8D2u/mbjD1mViZfx5ylUE/Nk9/n2ND1dL4rC46fdQ2
4uwj2LLkH8OwPiiKLSbFbCTRjCiEwsZ0Yv2BUpAAFrWengbZM8ivAKDY+Jg77gFK
HZ4n57smlE72PrtBkmhDPXE8tW5d9CAHp1t/lbj1FxOwXA4iy10qI7Ek+PjskqNK
XnhicjAQYJFHYnBHsUdIi/FUdR64+J2RNw7CoIrOPrweczXuq0cr7NGcijj+l9vj
YyrMOJ9Rd1v1ZvqYGTAa4fAJkO6OE6q/KHMxtLBtY45oyB7/vakx4e5Ge2uesQBf
KjoLaGN+VUAnDIY0q3WgGEXgkKEK74tZLGwpvdysJ9ItIuOn2cw8ned25YUTV8+w
gctCS9ykrIZjTD+tPOHopwQMzbTX2SPZ1me9SWVbtlYxGRRUMLHomvWsrMaifhnm
ojeX9ihfp15GO63k+DxMkyCt4nZy5taI2MgyaxggSVFWawsjZr4zmAucVDRBrfrJ
Tq1K5gQP9KU8g4Vrvgci9CkCLYGYPEGTsrvIFblaOV3Vs6Vll/l2YFQBh0Pw1io4
Nk40hN9w8wcg80HKFZmruWbhwEmF8iP99G7gSMBwSreeQEX/mgGK+JrPb6i2hWsm
8hIEF303dQGHJTG0qfpzpk9jGYu0IkgH+ovHuXgoYiF1rUXuHRWDaCfmlwljxGlz
NQsHSapy7KhgHb3DLloXyRYS7AnCY5ewojcFk+akuuSXDsFrVs1VwhJe82G5m5gO
qgJy3q9sx0r3XNwlpP6VUT8b90bkY+ocSKvtlGM5ydKlx4mixzgGYZ3krW23clhI
62rHZaEQUvgfLkdSYdkkNt2iNqSoJpbA3uCI/N2OkzCEnQqgH+Ya+gZrWB1P7/Qe
ER1fTAQGy0J8QDANEp/2mvZoDoPcaWq6rnAW6F4VqsNdHvYpjwbgXfGcLudXEvtL
XatWLfGofvP8AeH148jtzWW+xQiRyfKO4wzJRjmay3Q1ErN+kZiMmCG/Ar1P58RO
4U7jYvaWP/aDdS2Of+cZvliP2OzbSDMeZlUu44oOPBN2oNhxkekX6Fs4EBKrVEr+
xTtzpr8Lki4TWzuH89e0Hi9/Ue2VjzXrnQu83wV89pjMzEJLo4ByR2H5R//kzLJO
M0x6ZCl3HdIMt1V+BjPx1ycJASb6CoYvsXqeazzj5+EWZUxtdVClEjJtMEcj2EDH
I74BpDshTqlYrXvwuoYje0oG6MItnnWY3KiQ5+lhfgfEwSdkN8pnPvFUdlev8CeK
j0QzcpziP8JPP+j2KFkVuP8o3iEsTGQwq0vN5kPE8AVzjKYaueZJwWGwvk+n5pBS
vr0c+BU0udAwNZFijwwP0kISDYJuKZCAbkIq5AMcdekXiqoFHnJQv1xgZfqcOSgp
94wx1L6JSLu9LOg6jVZggEnPqmq3wxsy7c6Zzshb2xPGC4YNBFbEHU9sbAkeudtM
SgDL4IYcR2VWOF2qUkpKS2kkxsx6b1CVEm4NPm4kNZj7QISvD7sbZxYik0qfGDw+
lfQWNwMvF4UR72gpdk2uEiuo0TI2ius0JMb8X0RXV42DzBzVZEb4kqd8VWSqOCj7
3hu7Mzh6PoE1lXDssSRiEAfuB9BGSE0hILPjarJCW/J8F9TPHxhtDfkzFcPf8o15
hMkEjyLlE/Wje2ztHcMQOlrfSP6GW8F8xruCa0FSDsz8JDQGwjBSSdHRceBghtSR
I8t9TAGOxw82K6gVJxNxWQECDCVDVMVqbHUSjDxz+bg5rnzRC2buUEGQLhXaeQcH
UvdsJRO7rAa7+LeFcXnxrGkOdWdZALlW4MtskaOOucEp40zcEJJKrrO3r+suCSGV
AgJFPw9u2L3KHc6k1ZTcJIkwb/R1Y6WpF1kCN7hEXkoA8dpbKxnHrgcwaMKXdzTf
KKHal5VDLVkPexfpaWU/pmgJzpOJebKP07U3hR88Qj2gSVK6iuW3ng8rBtBy75zs
INVRyjo9BXZIto5i7hNXlSX8spqayyKZxgODUa0uZzxsw27zsdUX+TLS8OV5mI0l
OmGOT3pBnY9b7+AujLOSKrVThOhcaNE+Qqzk73TTqKV+2VUSEO8jHYhDJd1GnbWU
W4o6Ew0OYclMLvf0dfOqIbFb3io4YZcI6O2eF2eF2fD9X3UEzbkMi4MYsXgSmqUK
kLiS2QrttWfUg7aqW8mGibK3C4FOR+ND4029p3A1lYY/0eqhY6MS2DVgBBrk19Ed
LooI7d5qWAdR6TmwY4s1l7F9Wa4alZPVAdqDx8ZXXwthAfVzxgOZyJGowGEgJ1Bf
+y4p9kxrjr6Qg9POPdFArLIxwCXFjhnTllBnkgXfCGWFkTQgUCgtNxurBVBjPVGA
geKISF7bz9UcoB/pH0fwqPbIdjB89q7JNLvuNurw0HA9YxiaZ3qM8PX8FeJ8te/L
gc/d6jbTHqOXvF8tmXG+wBUtVfsKxN5dYm1CNhA+jo3UMUtv8VBU8js0WAKqAiu2
4W6MFe0C8xXxNPj7X2O6cKLnhD5vGtp7huppatH/+hjWXBAAkhpXzJwwptRse7to
+su0rRKWv8MoVNptxxcpNwyAANPRclSmP4bMvWON2iUfBh0hKrP43mDnKgUOUvPd
WNgpLVwhqCO2jkC2JN/3cnh9wm85KihhSZaHXVlsk8LE5QhtIv1/W1X+dpYo3IpE
EeodfYDpBp0HcGsKQHyCSCf0ZauB+8o41sQrcn8lK2lLQJB26ROAiAHQnq/9BTpP
un8c9taKjvMDJWDhV1PP7fQbMlMd96HIqiWDg699biliK4oe+vdbrMxc774xrZvB
Wp9zNnlnhSIVAy3T3uZzSdzXu49jqpH3ppEUXhJUQWPmWJ/nk5JlAasueJaPI/Qd
T6LLnLkOFEGVVQ5gEiFjc3YRh9DTh5zDzkPCJNUn3t4wWQgQkEveM/jETPPx+H1k
wnquRGWt+DJNP3g9jVOlytSxlJHWukmpC97yFT8T1e2tbh1pXoYNFTpIdNJAdzqc
7jAQ4LK0nBEXPkPnbsYaIw2sa2GOMVfFfzrwuFP9lKek1DTDyl/yZQFl5caTma5l
4X4ozAlr5n5BN6CbupoB1w7un+3UStfD+0xkn8pieVvUb7yEGFxzvZjCh96Gfs9/
RnfcUuKF81GXB71uWFUi1blvmILaFwEWj8hW4Um2/X3PKfofmfW92JnPDObDa6KN
RJm9XfG+xS/G4F8dtK5KC8Bf50p6gFlH5oCpwdwGXqZEd1IkC+AfcVCN7vhZMl8s
29/P54uAcQCaS3LrY/cP3DDgsHWXuN5tXQ8lcuQEsMPBKWFwcGVpVTB0v/sKVWYL
tpQr/dudGhmWnkhlG99oz1wUHtgs0hPEQPf2NMOJ2fEka8fU3eTmewsHlFZ0t21g
mRI5j8chWY+dqZrqgjFwcw6EzOSG6SbaqxcTunpgReZTRSiCaXM6nFv+MxXGzRE/
4QsEvQ+ovQHiDoLwfIj7ab5/V+vUtktvzvMNUgp3yV6vAAd+AW5xkd1ZXuRZ1Lf7
F2Cy9fWAub4esOm4EJjGicR9iS/WyjT8Tw/iT4MI7Q0ie1kpTpQ/mHLIvftJ0mO+
Bx7QKd0SSOkmjHKfZaFGF2TwCXKfk1uevm2zadYNi0mXf6ba/d83hwtYP2b5oAVq
bEeClHqJfejFPn4/iHxkjhIeEZuHBV4DbSKsaByvXt0hMUe8QWf6nYEMuU9Wb3xN
+ocEgRlbBWTh/8RpirQReHXYwxJQkqlQEED8B94GawXjcvvznIeAJO23iYPN5QMx
PxqrnR59alFP8wcU6DCP2Hz9c7FJLo1Irn0/h9EVN4m83o5N1VtXL3uGRusk//Iq
81LrWs9w8YgFWnxMmT9XU6qAIJfCKkETllDHWKQ6oK7vw1KmdX/gaf4odHH44aVx
MTHbt5ZsdxckvOlS7y2Nfva9CVvAb3zAx9hDo3E89cPMdtb0RoPRNsW0V++LJGwh
sJwINhecDOwa4TiAWzpMBEEjuUEK1W2l4hjhgJr09LqH0PqJ1W10cqfTqXPd6xDr
yJVMxmVqjqB4bv6WU0S+zIVfgQuXDq24cbecojK6TbRgiR5cVK0MQfyYiBhG4Ne3
B2R6Ueo4fYpGQAatbUF98awuzaGCD+tbZBwdbTYd1T75KRDdpBxHOEaGFjtlv7Xe
dt6fCh9wjjJQI4j/tNkQKgW2H4cl7TnpykrQSckhGeKT2Km+k4lNiH/v/sDdvlgq
jU0mxfqE5YYgLvd/1KzJZa7Mk+sLOWS02yQpOCzZ+UOVbujr1OxFbo4MExVFZzJk
rpbFLKew1h+XKuSuILC2ZkEg16tcao9EA0gFAUAPrDzjk+6cQRHMHwrAk9iQDRrk
j4Q07rvTyi/18c3bA1B/mDHryQRNYEe27jtcH+5Ww464/kqJLp9MQy62oGQnlOiZ
QxsYeI81gtj5IwdFTs0wU1iLLPmq303RGZxDYRj8oLWce3w3eQYbie6ZpAITy7Eu
ZCkSqjj+PNbhYtuaiMBPZEkK5Sq/D7jiLGCQAHS1lQOGfW/VKYT6V5IOeSUNW/RA
7n65F/jDE9qF/Q7A8BruH6qt9ks84fzHBZJIGd6aZ6bWrzBm110oZsP+OgeWNR5b
rLSTSo0ksqvvvLYls6WKNsF1lblxf2Hu/B/iLZDQ43K1JsZklas6ksnCuMT/UG5F
wthUeiTnsQIgkRRt+XEvOQ4TxAvRIkJTqEHDsk40WOM18x/Wos+jXjCX5NvdT8N/
JwfyADRtUzkbsZOT6jU56HQRYvNivMPjmySdhDTZVJ6Wk89rFPMDa2lQbiwI3Prx
RTykxrlfKJAc7NyEs0cqFx61wc1cZte4ZHYSvYtQhkktwdPbDZYkd0rU4CwrDXdL
6Dtb0LbjC/pTA4z1U6QWvwFE4JEc0A6oTtK9UufKm4N5Jo0LbvxENaIKEeQt+SvD
d9Rofyga7UAgWXOtY289UwRAC0U1tQS38RGMvA2PPbMbXfWBbzMoET+kleMV82ad
l081CDHRGCu0d/Nkes/svTm69nBJmapxp+b+RmORH7HSa+LvJdbxIybXiaTAglCs
qfeK8Fizal0CfxvL9TM1ulgrZ8+GAGhUKgCLpJUAYWbrfJ7kPagzesONo8ZanzL0
HcXDY2CtMpsZM3KxVVJizcoDeX9kCkS6Mkd+ZdL8zZkHAOxP7d1G08nVisbVwY6N
umqYKrBSJxOsmwEpO8pmvT/SzSMBSTJNDxVMdwCZWwhkiBx2BPqyFb3eRaTyyE0s
zIBCPcUIytUcm5F0+WeFy5U4mlJ9yLtJtGb9xLfPJunUuHN2JAByooqQ8WJGpIkh
Y558PoRvj6IOkH6I1Th4RV4Wy8LtMA4ORYWLzCdK/4wRQpWeNz9M8gDNK1AaSLZY
kXgpagkUbudz6T/fj37++O8JI2gQOl818tbBaaxfS6ZAANBiHf+08yk8ZFpIpZqb
ZWjwUnAekCkI5j5f5XP7370NYmbLetJwHFayyqxY/Kf96z7rfShx/UdeFaRZgQ4b
r4q3vfW1gXhJaIjP7Axz+Tr+iEr/5np+R6vpJR8+CCl0PoYCDzKVRxb2XJiQg6r1
5yLSjH4umdsmGP0fGcF2EifSrROoA2QjZSBRZ8LnKO1CDMjhMTbnBPy9EDwUKNMD
nNbUFkGvRanGL7a9sjpDKv60f2bB0um3d2A9JTUqMEBGaRdmB0LZRCvT0Mj/ZHEQ
p6ldN2yO03fBoCWDvewXPQNGfeS8oTBrqkB1NCeOtJBtIK6tXwM0q/pqBFFIUOFD
TINWCb4XnZxfQ1SglNftoYrRLg1Lv/a38wxl7i8ZiTBFvGiFbMwD3H+herl9Afgk
MDnbyIrG0UwCf0PHXEtgnUx6TPI9HFUBJ7YVg7/dFYJeXFPnzsk/pAsRkdr12hsn
iWVX7n3GZTC9jtiIEXt959g7XDJc9Po5lET90i7Z+2j73EYWzMD6ESUKq0cFNPNE
v4UQQ5we5WnnoCNJ67DgT5iua47QWX7NbsKCVbAA5kyotAomp8FagDu9fTlMrELx
iAkk+3VETf86CmclppusE6ZctL/6BFTUCtts2UV3+DsGvaYu3J6lzyLFpI4GcNFY
e7mFSMaAAdeDqH8tu3unshe2oCjGdxJMUYHafBnViSe6Fpg4D83JEnLXfPUZxsFE
gRjLLDX+RQy/hwLeFHznFP/SlK6LXl09b7Ky0VaBiy/Q9skhJuM8DI+dnJSuO/da
W4zIeMlQq7oowC3D0H1b+Z76bQ6zmIKamVKxv25CuToCZB/HCHEfp6Z+7WhpvIS+
bTgBh3QVpm9QqE5YetEo/27Zz3ESlGT2qCFJoOQww4H4h0d73pqQ8/7tWpyqen0Y
E+IPZStw16NbrLaKLxYR0wdexe+RrE4ovC+57PE5UcQSBLTGbcudXWauOqa3vZ3O
ozaW6hQ9cpP/dP61DolV/CvAV2lohSO3ndEYNkaxUU4zmB3d1Q+20/MVARY49fUD
X3Etfy6qIHzyxzTZ3lBUAgBzgZoxLgc3r8+DLWuWnQEF9OOmzDj4io0909UR/Ex4
dFoFfVpQTRIdcPB+z0wNVYSqGk21Ve5tSV+YskTmYlym+ZLJCOAvqnSC8i4FHfO1
zXw1vcsORXQkZifZrptzK4ynncXZSR+88FKnHCZLkodBALzKJ+OWgFVyFdAnuGLk
YEwBOkyjnQycuJnG/7l/9CeMsF93otewB9tn2z56gPk7tzIL5/urL+RfHfvO0E8t
lNJx5mHyLEpi9uJu6bz2zPGrE+4gO7EvBxrOPr0ncwrTE8xT/a76iqU4lk/ttuzG
mduKnN3uf5zCoLpBohAFdVALBtOzdqvpcWYWAc3X4oxb1WjOfrHuKk4NVsXht0dp
AagAumHOC4Lrn1+PEEOeXwWvoPpdMDA0u70riqrOtsRocjjs69jmZwD1CJil6gF+
ayqsoOY2ltlmpuTgmE9FICMKIerOakdcvUU9vupUKOy4N3pDzV11ItklW/AwnEej
wnQgjDIz8Xj8NPrJ3UelYyY/PxijxF7tGllpMbTkFEnvWkd3zjZA2THoDD1BsdqK
Ls4RwS3ZTBNd0YQwUOOFqiludTYWLeJ0FgZPzHo6OQKN8Ggi2bYvC1zWYYFLyit1
41HEV/iAC52i12w45C/nf5ECnJii2aaBfbpHXTXyhkp0lBS6U4/M8IcfjircVzZs
UisCK3dLcI+aM5/G6MmlDUahT0tqVX+6UMANWCLolXAlKQvMvTJpbUIiN0ybcUVR
I+V73vyDftAjP74z8lNPxQbICSozY6EDS3CKKHPsLgpvEIFJfuEFpd4vS2ezSup7
Rw65kFOeybqQ/Dfufpui9H7HRhYQf0NhA0cprFOwYxp/OPSSceZqxz9O+Q8FjJdD
EA6Dtq2RtzGcknQkcLAHLerAaq69UgSs/bf5I9gfqh7g6EHLOWMQ+1rDzAdZ4A05
8WbhABbYhhJfDi6jf+nnGiMtr4kh3SA9KrP1YxjMdLt07z9FzPvZOo3lbSmHYiMt
Sgam5F2mIoz5jdFl/MyoJbdpqQhT/jis7fWbF6E6i7JjEMBJ5Tbap1Q/Ahi1nHPh
7ew2gY2yexKSPF+N6gWoS1fbywXZduvOgME+jTnzL/TTgQOsuHn8oVJuuTk64t+u
6I8Hvi/ib1VYaF21rqgTS1wHvMIei0fNJ+60fjNRs1G7Kb/9tiuCQwmkkRJQlqYo
bT7A0+PRkKPNHAzEp5o8IwTQmAxNwlLVnBsEVG3Ajy+c2pGp0pkMFgzytyz8UmqD
R/WzEbxMRlG5/VgeDg+GyKVOevNKrL6CRgtsF6mJM5sLS0um8tcF85aUmXUyNdck
wBwyGOzLJ4piMEPse9GFRFn/q5JA7vYNPQlhNSJR9hc/U/DjTGdWwfp4ChpIdIro
bTU0Rb9Wra6lOc4dstorU+U8v2YQp2I8OZOtMbnYO7ej5q4yUpY6mTRV6Dmlvshq
Lxw76rkhhH+ZqDZqCyJdEu1dcGnIWUmcXdZRbpqpBgUO1oo10p+AAKdxBoQNPlJv
hH4IZhUGtCBrDnqfT2+sX/3OagKC1epo+Kmw94z+tChJ/Q3BLTKU729pFyh92xiQ
oEjH0/1D9tBtr+RzSt+lJu234gzXkC0xOVlUI/s1cZkzG1D7qs9K4oe8UsBk0h9C
TNAMhidZDDjBbIJl49sP6g8Tz7j75zmLi2jHEdYc0qK1cRtfqpFR/erhQZVy7kil
2GmDZV12Agk+LuB+5xlhTV8YGFnazE9A8c+OrcOqzMgNQkU5qm0W8y85VG3yhuRa
ewBk9cQn39ndcjjiA2CVuy+j5MmIBNh0LS3ZEoyegRStikX3SjxmbfISp7dq8mcp
4veqzTxCQ6m16dGTc20P8TKAjGNvXX+4+/1S4lfLglc+HBMVNY2sizpriwGaIU1+
AN6inW0VFujxjDYbMpPKdMepOmKSTnYsafS37fBQ9GA962bAITwpaavvu+Q7Y5Z/
H/TP1dXeUzMp8ApQNJsbqKEFu1KRlq7CaNFHpWp7/EDdHXp6Jy8kdqRoxxBhz1Jq
hmYZMqFZoN3f/vQT058+92Uob74P2Pc7TLYg2xCE5xi+8kxip17a457wSx0HtrD9
0lA/uSPFmmS5vBZSa4wHR8HdC2GEyGoROhd048Bwv9pvNKCld2JL/vvVqClAquLX
rCpwyHVAojmwpivIxPdYdVglsDB1E/YGIEVuKwJb0EU1FwiZnozyFsObStIgSnT1
1JWpU1vqAeRJVtbJAl2jctycwUAOgZ8Dc1E1GHOWFtK/B4L5vQ5BuGQer3h02GTA
x8H0wuAERxAOjqpp6/jUZSw7REf8JLSg6tRHtovlGhASiRWHOk0LEEnqB1qB3Fo2
Ens+WNF2+N00ffoDggkyfM9zA9ZcDyGn6KLPD3UqVzG+ZKIPsIK6vKgn8kfDbnLB
MSMtZwyvZ72HdjQpSG6UJooaXnde8znMHwmf6CK51nZLT9mt3wk9TzUA4vyWSJRW
Em0YIFQ6ZQZgQy5o2o71RRrzs5Bf/ByQA88kwnQJyxFN0+F5HbXYkNhUx95Dgjfo
dvwIqw+o7OQuDKeFbclJoMMzkrOKxzGwByO/h5njH1YGCbaEbylZb570/2/R+k1m
MB6C3rgEmaW6MpFaXJrCdXg8CIJUMMh/NIqtg7lTxitNFeDPF/yunK836R0VggFh
KRERuAgF1ouTh5u6pKh4coSM4Qs/wO2HKSPs5owtXAgnwL1s0XETQys79Nd1vbQx
clgEWtUW7N5yqlgS9AthrZliY0UAWCm47M7pn201Bjz1BV7uBq3mYFOu79uKz1/H
Kl1EDSn2GNGeIbiMkzH54ltV+SsaQi925gGAHL+gbdyLERQxuxXpNE6xuQ8yTDDW
4TOFrCHK/7z3m+azyKRig9vvjf7y9ndhgntX6FADt1hnuiWNTjxVsvUdyveN0bL4
a/f7iVLmHpAEqu0x04LgVmGJITGDyTxaFpOmpalTHDPw2tYLFp0hEsp58ndtxUL3
t94KeQ+KOt2U2PE5EYHYcMRiBtmIp/7gTjGpJUGDm8hjakr/ClNJtnJj8JTz3eJ/
KCcJ/L5uroXoU4EnjVZp9xfVBxh6NFxhvGD/fvdhoyffnnyFx3fl1TrFRTvbRsUS
oOGI/utFIqBBEzAE3vgb+qAb38a9CQXRbLcW7uLgVL5/6R7CJiQHJYmpz7WmMQAJ
BTzkKc7sUwuaSC0f9wCExi+ZEe7p6YlYQ8oEzYPoE1T0WZ1zhSMlad+493LyIczA
HikVlQpKl1YI+94dsZn5jZ4NhEwS3GIiEL66S/3ZA/q91Wom7xZ7q6K9lNFCskne
m23cvODOi4t3b3wNnS5OanQNmdR/8TNizlsivBK+fNWE7jtG0s9metuDKz+nm1YK
550pj6uYBkSPkZp6QYWQ+QsBw8zTrtihJYbEx/Jv9bzOmpY7yovEu8Xxz3YeWV0e
4CosCzPDqisGTSP3nRu82oxEmFtrpb576Ij+BYAjBVH3XNCM/0GVFfQSyGutq4Fq
heopdFrnCeKz07/fs/C1gUxyBGSEWN6S/gHoINvl2Lb+Wx1PsI7JLLDUsLzVFwkz
P2BRZA9FeBdy5VHfvVqIfLwWf5zNvXgQt9S8kXMkl8Vtd2ntRze7ATyST9d7ZlLn
INH8HsWBY3nrSk/R6g6zBK192BQtG9iEvH4TG0jt7y6NBuZZpfUpI7ca5vVJXUKv
HE4fkj0tPFED2KBtTEL/Wb8g/ypYgCExwGVgF1eALJAvL1agOrE96XCxyNy6JFq0
ekQdqGkbQbocq37R0Nsttkt4ARPNL9oA3ruCcx3MJcGdiJgYdYjAxjLe6MqB8EUs
UNTE3YDABfkUM5iQNGskJxpdd1c84C0DW8bFYGFBypXkAaaW/J6s2qXncIDdod0+
cfq0tLKj9smyW8E/kv5PBb4s6h2l4PI75D45UD8Kk8beGf+IwJJA3ROD09v6qOIL
kY7IDpWLBGCyraoOS4L63EOc3MInG1g9DYMBjA4qRU4uxzAWfSfI9g7ia1vCpZg3
fCDjDSfPYCyZBd71JwQRdqj86SioOHoRdQqy9dGMI7dtM/SmGcLTLSu+Hpb0dCUc
CXIEGOpUXDH+5Tzu4zSfPlhHr7OYbeva+KD3ux+pB+JzUv8cgGsjnPQ6aq2cccN3
BGrrw64CaYkrWIhfazIoDeox/g9pueqQkyDXZhYEzdtvLe4lJeCLzKVx2xnDxMfc
o+TTqAnfONLCYBhMoYy8d/GykebqUPyAks7cM+lukh67DEYv59vqhH66t2bw+4PS
H3WsTlLEpfbsrYOp81bBvsClnwXaV5LgSqxqNZYNPlo/hLUucbaOkoHOmJbjyZpP
92kCNnfC+4yUJzq0MyXtkmgVj1OzWSb7nRNY0OIFYmHxJFLUTunnMa+skmF6dBt0
mzZGc7Y9uGjnovJqz8Wm8/dL7tCXeZPWX+EMtxs85peUWJRyYFCHiSLy3qfnSfPK
9RcUC2t7E43xCPUeZSjqdmRK5eQUd9tNAFSrrBWPOsbx/Rfn/OrARKTTrtXBZqIh
eRhrtPeebIZfKPVPuTXXu1ukp3FjVrJM8+1zs0YcMnXFC3kyvg0GsugCo5f565V3
hxmRx7lOZGid+SaVKbJDWC5FuJz4I5iiMV3c3VRLlmaaTWcIHMhhy3eIo/WYE4Mo
oE11oZoDmiAWLDF/MJPWxquXZRPRRuddBmuwpQeXJuAd7plqUog7fL29Dqqt1q9A
v9GhwDwT5nfI6kCTzuAN9zr3s/WV3tewvGfIljkRfC+C8r09qGFRlJXQHBpFQAHA
2DDEVMONa/TIj7jbnW186F2EtOChdvaOLUbAdixFOHsUCxqoehZiJBWihu9YUOhc
OqSOlkpOfk4InLXpjblhpb+qUtD4Tjf1Ye3EFCOaxZxDFnJAgUUJA7qiCSMlCtv9
U+95XDjWIyqnJqMGFzVE08i97YH9Rau2KzrZwSuzJWftBf7fYdNCKv36z6GrGMbs
uL5nXEHXBK7ZjSuLap8rxm1joZPIReytb+ZUOx32Bj/MUFiuY7n+QdR6o1YOrD+A
zeeTWoeaOFZrf+wxqEzayE5dG25SNwfSF5cSUuCb4jGSgkYVJTzEOD5MYO83yS06
hNTLN/zia9ZLv+GJQ6+AKop6evwMKSryPu7vO9a/eQXO0joLilnzSYAnrGp4Olpu
XEE7kAgCnSRu6G1BBmrCdwBISzCNr0xpfbCzQeNtIop5KFvuBIu6dqQPxv9ziYMU
7CA6EU141cPx1k+Vd3s5gWv9gYCw+DjAirI/HHCB0Ic0VDa2TK+kBQhCjQIBx+R4
UkPcB46JWU8x8oGX/jrVH+fG+x3PMjVNETsjW0PyEVH+ZXqV0YEpZCkZroORrFfo
IJe0u0fC+7jfPjx6vy3h8ijjhNBXzL+wmdLyCJIGzy3D9GcyyQWiUUpEb4IG+moL
ZyGQKZAyxJmh+R9+MoI5bYBf54LmvTug86uX5iKJnkh3XJo59wMZn6jfvqo7s9fG
ZI+kakhX7WyRWvSxhzUEeEpB9E9cPcPqtFhE/0OkAxpv9VeHYZJBBO2VbL88Ibs5
oxVERzyltVZp57DjuY4ccwA3jIbZ66oWKsgrwUbD4gHYwHsNyHgG9Qky5/9pjlAd
tYSIarRtqi4QKExfjO4I4AKoW2MJOxvQeJ/5zBjfqQY32bTjFRoJ2Z/cDK12IOW6
LrhlKjh0L4FPmhZ5YBlYK0BQKoq5AMBngBLfMRhVH1nvqlHg7xVza1UW1neRW78U
1n2Cdt+/9NpJxq7FRTSBukVvTDhhL+YmMGp/ZUS1Bi6xdvEuJ6fkSiqS0yO6j6li
En/+yDZLc+y7lFruZptJb7Ori/yifeQ9QpSOhi4jEM/bLyAAvMbIqhIcMMeB5CXB
RWD1WIpnPSf18pju0wAuSgb9tzXIgm2P1evbKTawfYfkbuf1dhHFSvGaHZNode3g
rVoAI0RMa+cj+cgQQXn9m4q/0ijLjcfjbrSBxWrw9t34M23EVVGOSPDH5xVtpSUd
ZMl2MKu9UqfKPnU9U9IKcz2qqtUhB8pskKEVBETGQ4lowJ+qPfbo+S+Rjv+whfUy
MBRb4UdL9S955SsCisRJ6ttXA+isTTqB811bOsPd9mfvWS22tI17IVSiTNQsWkww
Bz7/vM0GGBUhDIUpwKLT0eqCMLdp5BsaxlRWuTgzQ+vpTTB549kS1QgEM+2vOQEb
GsvHrjkW6+eT4b+ZBiZomZvDNaTZQ7MRpn6ixTMBTi1pFzYmKlIp509MgGc+i5JE
aogcP+KWz4eA/GxyT5U96/ObxD1OMU32XuKgKZiXUljbTIiLJiBUqndKKA3Rzptf
S5U9QYoP/loFwEXlX90Nd8E99/TKzXTzwZYq/vnFeK+qQT+9jV33RAyBplwgHWAo
9eeKqbF0W/jhuidhCIhsx5M6qfHKNxgK80iOEueBpb1AjAO4f9j/s/pUexft/z0n
/haBbfsJObLhAu07/EEZWDHh5wOcCVSnnGJbGqXYbfGI+IqihArjZsHVYB/gbbUI
iTtCbdoXjKr5dU26v2lgcqK34Ay/YLfoNyIuDaa6VNrVtK71pnugTapvdzerYt1l
zh1WGdJV985oZR/3AnQC4dKjXvDLZAR/vmMIB5wdog5Y+L2biqVdI0gUNbWHuG4M
+Q+Cr4YTU7efrR9e3a3j59U6jBJEwJpHSC5VP1y1BmUSaiaIv/9S2eOoweNk0Alp
kenwZEBESxa4oa6LyVHqpch1p9dBU8SYJUgD+0awCgMWvmYzKO/ALVSK/WaWNtI3
Av3lTJ7sigYppOjVUPdfy0jdzVx5SWFCrZRyoNb3a3HwNHTpyTfk19oXoP+E8EMk
SFMryXRhzaZlvwMYnqZIrkExkZnxrX4Xv3pcQunDvMAyrWxTpwaQU8oI0rMjMWm5
vZSZrTgKsAfjjDXemPnjR3eKLUboHEGCduXjgrxmw1PVLzSIDJZqIjoWwvD50s0Y
lFl+l3AwMI6ubowtqlKxYH5xTt8elK9Novh4ZdbnESYwyRcBjFjALr1pWF07g3al
upFPObL2dLKuMmejRG11b3QviXE8D4gkKOkr/AaoLWon7Z+XBNeYg2DgtyyFtY5R
7vtnCrJgqyFfG7ULiqtyQsBOXHyI/wQTDau+NRUVCQ3umm0g5wuVe5jqXbLcRNyo
1wkqBVB1rwLC/qHSdv1sIRqVAGPx79K1WAfUDw6ywWt0yTWOewosvUeReytRv1Ud
WPHYxNJ8o5xbxJOwrHmruI9RMi/GUJ1ktnqp29/iuVb9QiG9sA+OBWM6XYl29hP+
hWF16NDBebhnCanTUgom+tWGzHbBSezgX6vKw5p91fwLROj8gvqLRWuN1AP3vLKs
Ruk8JAbAy00VsgQadH6AGIzHF/plRJ2J1YhJctD73aE5YPLo+sPvC5GuFXBah7hX
wqSzRSzSQzueo6GdQhckP3JyEqxH90R+SPLXDKuecQvExdH4IlsB3IKxpvR4fX3q
ueZeZsgihmix0kHZ6pnvH3PCqFP6kG4rwUGpCVsB0aQlq4dvSJK7ejB8pxNAj3Tp
4/9ZruqUh1GeNNeXrRpQDfwGBcZnsL37IDzkOmWQzyNySieU6H2RZFVaWHVHFvf3
TxXN1SGlILIlo4IVoHEHvUo9SpJoiFAnkM1i05G0YNhVYkG1Kek2yY72qGmNapcw
o2m8lafXmw6ydWAiYopuniKr7WvKFrR8fFrTNkdVcldEJX5T6dat6kZRYKfZXi5r
GAFgbr9Kmawd01Jd9UyAjj+IzJCYsFYAKP+eBMm2ityI3kW3+dOmTY4vA3qN1+u9
SLk+qvVGjnkSlQwzMkJNLHOMUtPPLCaYp+Md4XLnLxEuL4KIXmdlUrjeL5K3wgi5
BUtrXGJ1PGF4HXJnEgXcFTOUktTGBF+m5j9d6IKEbJWDo6E4i1ad8PmC2yiddDav
V905/4AqIMJ39YblBmHpDCSMZsC3fQguqVEjp3TtahpgRjVwR0HPNw/SdJT2gyCd
nSdma87jJNE8Pt9zOM9nuEPfsOVzWrd+eYcuGhI1BAGbtPpxgJsaL0T1rh6VmbIj
X6VbMsaxPNOvctj7Qzrjg4RpG/WBzpU1CHTQUbZqwfUlCdr/Aa4B8VGHYHB8DXee
rqBF5YQKIzN71tJ/XHnasmrSFU/KW3syJhkF3xZS/t6sUnj4ZC8FwnsBokuvePbL
OpJ43idcsXoNoQLu7KLVDqE1klLVuymWpR5Tlcqb/U0NXELtvS8fra+AQHqfLlxV
LEGZiPyJryAMsu7+EXslyvD+UjVRiBm+v4s26y0Bu0WsO2wsszXDKnNsDGpckjZl
UpkCoAn1r4R+qPHrs8srI62/NPoAoZ1vCCwrnhEClaPIKMTksKkZ9+wnVNLy3M6K
Ul1SUksHxenVDMUwXICPooD/fVWX44wNylkNHMEgCiHQwTft01dQivlyRMIuTPy9
pcADOMVr8Z7i0gzsozc9oatkSRhNld3Esemm6DZYqFyNH3llemREILepezOqwSSP
fGhOxgBw8YwhcRmTgoPYQiVHEQ1J9M6+jbCbCCHRS/RrvWw26UJDlVJYM7b1aGem
yFWaAn7/LSuP4Fte3O4oJ2A5NtfVp1AWPlGwRN+hadOVglEuf3PWwLWqs6v4bEbI
0hqlHD5PcGiNkJe5nKSzQ+4kGlNAhr7lS4QANrp1zcWGrfkjEJwwkWiAQWXT1aL5
/B9byrTKXn8IvXn5n3Wd7F1ia8Spb/iUzBxAFt9gp3XqbJjiGQTM3WsGo4nYB2Ot
61TcRmtxSbgflwoqUWUO19uj12igMG7VkZTrOeGT9CyEFqz+fFGfbkgsg3JAUU/I
jm5J69EktAhVkTClI/bbwFOt7H1/cf8nYeYOT3A+JLwH7iU4Mc47C4h5Inmf3ErV
ywaH1eHXfH4B0HG6cxmcXz+Ru4ngPfcDhQFVxPVBAK6ipwvH4xX/u8PXYpox1cQV
7S/1abRAP8XW72TL/OCTAl4+O0wWTFP9D0RS0KDTmuP+aVpdWk7DcM4VvGLopDl6
/Ez5jD5uNStWAMUeKSjdZL5yOou00oVz85mK1Vrg5/1Bxg3uUnd13g/nbOBAk8ok
uFnrh/7hCmOkuSI4yHXZ0ET1ununLsP01yJnGWW+vv4rGjQqal2siUM0OqWASJLA
jqjRY4p1DeGKH0aqrAWoCTGzg4afqEnYzUTKK+BWijX2aYYcoJ8ukomQkomUXBdL
xBqAK4OdyZJ/j+O1rDTYbo65WmwuiNIJwEWL4+CTi7f+krwhB59UU5kLK4/BxISN
OR8a+oTYjz+jPrnLOvWbyXsNgAEOeVfR+FtkdSZY82lNNdpJ5RMC5XGDUDqPmWO8
+R9fEE99Ywt3IfA9GD0abO+nYOU8Fjq/++uIh90ir0m6/BgEW3InVBn7NsUNxi6k
X/pARaO6DMt9OpevJx7oL4NFjnmjjDabeJa7/sajuztpWWFCnJxHxCYSJoE0e0Pa
tNk2rxXH8AK2xhZtWPA4larS3Jl2c0sUHFgHcRrPnWim4RNvnYysyMB670QzHhBh
3NbHALBh0E9ZtBee6UjoqNg96twAdZBvikb70JW3GdUz1HuVUnn8qh2yzol9PiWg
3ZWRB/442Hpgi1K6mgDZzAra1qs4V5vRdbx28POLDLFZkwZUbXbmWzDbjG2gpDiD
mjXvs5O+V5vKGX9BsqeHfryWuWjgeg2M0tWRlx6o/jmhkpNxG96u3Q3/TXk3pMtT
Ibj1o7WwP068ZTP4T1aVGPnK3XpH715DQkklFrPb+GSZ+GVxaRgOfCfgR+ZjpOSz
WOOClYAqHtF+HhREV1ThdY0ugEdJ5GDgyeoYxIionekEZ4yug+8vsa6ZeeCKlyPz
lcQbAc9HfpEBgQUSG4rc8lHtqfl57WjrOZZY1A3sehruJh5E6jbcd3SaeF1sp6hC
ZnQruD/KOIggn2glruLnWlb7VHgOPp/uGm9bCoAAENJtfem3DkxS33mTEq1DvwUc
3z+YeeUnShVZGVXWevi5uzOcAyEjQsv1aYJ7r+WNz54+Y8v8p/ep2ni+5zgWDt2t
dKCtPqHsAwypox2PfcDVIz3jaXnRmF5IPZkQItMOMVzC/vhP2hAUwRB3zxMMpHgU
pMilpbpOAMsJpWLZExLm9mAW/xksumFvq5nFhRwiuMGU+DbVH8CJfGub9D+aye8/
U3JXWj2yHq/U5OaWAZCpKNPROTCG6y4zM44SZELz/diUmkmZk9yd5gPxuT4UFPIx
RgoaPg+h2Q1q33Z3G23hRcxVuLaXqsvObomHZng957g31OQS9Fl9XbmzD4hnwfqm
zluH2oxzIq+MShGdCvcsyssMLbONt1b/Fg6YSJYJFV578R1oVgX+tUkLRqcgMsi3
Pkn1cR6ObRzjr5RkxEKbYz+qyYMks+l8A6nQK1CBZoSzUqgS7w6O5nYhq1qPiHl9
vWh9UbHaUj6t3K5PjmbgMjy0SVah7g2YYzRqbd1LdaqykMZCQTq9qv5wk/HjxjcE
dmHJITHEs3nl650ekJZU0wDWC7YHuDN7VgeJ7mlrXmY631Wq5y4l0tUNRD6GCQLH
B/Fa9Au1Vvo6UX1wkrFE/9lh0O2CWTICQ/Ag+o7HWQqB3vS3TfLGF8fEcGyynbJW
VuZS7VMtL1kuTwUSO8baLZ3yQb0ODVTgfHL8aoaz4P4OOSH8kgzEO+EdWSYZQ36X
JrisKTTBvvQn9tcJGeA2J4PkuBCMucS6fK2i9wMrDHQWSmThYmj+bpID4v1a+PaR
CfDPt5OaTRh1z/8UAmN/TuX7yCaQ9AvEAi3GoEG+Tp4NkeQumlZ9ka6tAZwGIWqz
yGBmMok19zHxEOlSiu2YrN3pzztMHwAdIMKVU+4h/+byjQbjUxB9mFh2D+DLXuM0
Y4afZtv1j0a6A6jVprCr+01bD89NJo1HBu1cTWxde/+8KmUo3Iqdk8KEIQxywFcc
2XAgI8yVbl8ORac7ngMezcAlV5WS2npaXj4oiNDg8CjishCrjwR0T5yPJYkDo42o
3sorCbKLWsM6P4lVSU1wK170E3qC0STotXCVKUX6Ix9hTHlkjkzWCCyqtjlwtxjO
QpyCMwfRLOStDKx2TzVSIiWxUJTCNeT5xbD0uo556xCJWPdkEnvA0gEDk7IgMwya
9itQoFonTt749WPCVU8pc1fNLOmvdzGOU76UnEfXmUEkHQam4HfbenCjfzXd3zmh
tYjNOlYnQbTCmBnRhOYPoaNAE6E7wDmnlRX/2dPn7ZxvNVzZ8GOLKpAvNEVnvSYn
JuwfHKoxRCwxtMMm7kpdwW76V6GRI9Bvat4C3Ec098Qbz39DOMxoq6cz1IRRUSsK
I+15v6ZTZ5oTSVXAPUlUWhNFaFOxMSAi3SU6Pl+4fBMhyMK9hZSazbm/yq4I3S0B
m2Z8tQuVbU4zZCjWZxT1Ess89SR6iD1OOEZLL4cfG3scdAkBFEDw0pAOh8JgSp+Z
wjsUK/uaLkJRnPXfC3orfbFeVAPnhVMYJB86ayDtTHkFFkHk3kPZUx4I0AmJzzQ+
9dmwzG14G38ooxReRcUp9Ofu2MM4S1EyQge3Z5YOqQA9QY4VoEdcWleUFehUv3QK
JVNRiOHv4bAYOEFhnTtoqx0PlTSdk5nU7nvjc+IcTGIv3avTpBx4SwoKp+QGMYDA
Ksukiqd+v7ZtkzRSDfb33Nfk5kxQ2rPjs1PSItl00/Uvm2aeHWgWnZofGgjg8M38
H6/kxXetIJgXO2E78N6Yov5lVh9XMuIW8zKxsTBync+EGkqHymgnYsBqqBqbO2KS
mh4DkT9LltcckC4K3DT6jwvSa2vlMxDRAWSDXtaT/TTrBtxKHwCqGZ3iAqj0jzWE
V1sl4bfddF4jwsmX9nBaWA8BdB1TbWSXoTUhRsv60dexef5+QGfbTt6VMMppz8pR
RSWKTup9DH5qLEgGYOGp8q+g0AooGbslfFhWq5oWWMDKNEFOFDWehLH+BpibwVjz
pO/FvboYYF4N8yr+2RtOD3FTnXCi0we46/1/cDZ5TA2bWKVNGhbz8T82uUZEttb3
gZLSKf1hqcJPGc6yMvvAmpNb1xqIPOUOCnB3ilfUh0kghp1wXvo6G2f8Ftp7zKG+
V/sXLFiFZoD6tyzKJN43G51N9mYxLibpizTRa0Qcd2SJVyGrP+H7N2V2uNi3Rwk+
V4o7TBJDQJvJnRysuKfGR3rMNDsf9vKS2Wi7q2sYn/+zwXz55dwLLchcQ3a6pVYI
lr89QYMIWC3PxndXBHbzVGNdutObftXGqLuAjnwGI6E9fMc8KeSMmOqM+GqJre2k
20R/d+AXfRFZnl1BtdK/jlsAeNgUAq5QTG4zbRsgpwRUdBO/8srk3SpymmSzka/V
XB34uDInkSMbXTOeKpSP3qGC3hRK4XaYilVXEv7peozbukuTO+1jHs97rfMQm2Lf
lLZYD/Xq8SE82ra6fnQnVyqEfbLA3aTFHzGYFhAOGNV+6tYcinzORmJh7mlbFnyb
qzFt+3Krfn+Lj2QHJgtxBb6RfwHdCm8NJFr3VKGKAOp2D2gTdxR5Li38JQltbSy9
SOGhX4kXEhSKunx6WhHIIDwSClh44w2rRPfKNMapRtTH1qTeMbUv7XEW9xgwiVZp
9Wjk05wEkFDojEHq5NsudXR1ZCgBQmy04/i7uZPzwtfVw+jP6Y1S1dJWESl6yud6
WZ/En6ftG3GFYGkIHN8AmsDbOkv+ZBpXFTuUu+F2OLACZgWUIMWVwfg5SAD3Nla4
hgzFCUz8mUI8owq+tGBsDnmeAP/Fl/xTfLK7VZTUxz8ruRffIVCPEswLawAsVDG7
U2CaNaiPYockmP2jyDWcnW118eWipd8rDsKeJcz4mYaXEOT2xydq7+/I9RYdBVow
FZ0WNSjNjXha+H0//SCu0i7XyCzGSl2l9hqW/CFiWLxULFv0Posv/GRwAqVLlgge
JZ8i3KHo8qqW79fgLVuatHnYmnX0rOoXCqCY8tsURoiC1PHkHtgFdk+KQzzy5Gmf
xSBJ3YFpoJvM0faKQh5bNglQbUDcJqlD3SorSpu27zQdA+Biwyh/ZbO9uXE0a8An
wDmBpvnnv7MKBPpOXC4W8P/cyBfr3hFEZV++gzC1sXiBXy/9vgOmAHz9u92iZ1Rw
yMGBTnkJV6T6kmaWp4k90DiG5mqGTP/9ANyY7sla8LzgjeICsbjVxAIYoUc1zlV+
Vu8BXYr/Qvr/Iq/zVTkEOsUpeot6WZ7/6jG4XuWEBLZDIzuV/9Z6Y3OJht65dnYw
FPjvgkjYd3VkhJxPifIf2F3pz3hsbUZpjEWZNT8zMnsKWJ1RT30Gt9754Pi0EaHP
QhbCccKkRlGDgLQT99cYz3qoHqdxJg76wq0Df6KV/MiIm5d2SpyEIR7xa4yLfDhV
6GdjGTbLPy0hs35FtnPJmNK0A6TLkBXu0iT2ETYXR1U7k+kpToyZaMFI5F7M12En
b0rGKebzA4uUwQAWu+Mr9rQmEq9JmLGv8WuYhUd5t9ORGyQLIk4w8xrlT0degWgV
3BSh6pQBV+88OmCbtAu8PqkHsUSQeDVBFs94DsrwXyeRW7h5DhufY/MsWwtkXvtA
UbZP17Qqg8BgDvmpHw0fuDcRJxvztzGV/w27+qoEKrMv+feQG0OsUqHPGvxocoeY
9guT/RcKz3N1w2VyWO4JOVmgSaazGwIcXYJjqkMb+v6rFt3l59RV6Co56vHgA0nC
WDcCcM5xi/bWtB+20pQPFVgICgRfbCdywk9Qn6Aqg+8BnM+4cwAc9CzP+/bTXa5c
ouKsnRBjWcBSlPpuIBu72hc5bxZ4UMfxCQKzjd4Daiz9sW+GVmzhnpB3OFQnk21o
XHsYONp9Uk9bcJ6/+GW9jMTw8DQ25WuPBdnXR+lhGobtcHxzIwlR8AxRGZ803sp5
4fvERvTV8a1be10L4k3hxvA1G6tp9uLkn53FlU+nGbfP+uoBbL1FM/S6WUsZuEFk
7RP26GzNACBsdy52mUAbHJzAZLeUQW8OIUqD9/7yoDvccZijtVTuT7qc87bMkH+N
nAK7KK9CQApGbI00mqa5kVLOLdedUQEwhYlKoLReVP+KzaKXsSTXn2kWg/lfB/Mm
sbEXiweDYKwzKbWK6w5AikTQWk4nV02jtKqrPW6bhRGLXpGXyr6eOEhQ8M3ez0Wx
ewbVZxRs+nDZM5Ms5vZDJCmLLuAMk7VxKbyk6Y0+8PDForVJI7RMpNZXfFe6c4d0
3ZbXH8DU8m9VjMqDrw+gO3Gy/JBspRHeSHRsGmL0aMVtkeC5r4DUj6Y8lhJSZiCT
Dgrj+4dWYA2Ju3DNAJzi8N1GUcMTrN2PtksDrSBFw3QTCxQYqQr0fuYWBXZ8NJtf
922DOCdmcYgKZetvas9RO6zlSVenBO4WwBSwNRLod4YmWkzx9rcTEhPX0pEDPTR8
ZELb3BQFzMhV7G46qRPsUENZHiMgRNJrGwT0F+AHqzh5dis+CLfs6U1XswBLl1hm
RCgLfCk2EgYghZrCupG+mmDNyYgiSMB9HvRAcXMoIkLxCd5KO33bRZaKBCZrSXmD
dLckO5BQ3IqEBEiQJeCnd5Jf7fJOciIoypbfiebCce9z8fKkt08G2OgR4AsYRgNd
E1wN5ObohIituoGP7xlLOq/tCxNuZFXl3iZ9RI/jhKtB9tc1sYsoDiAr82pvK+e+
txmf3u0BPvnrqPJr+hS784DZ9XidRvqHSuMula3S2cKIBBKM774C5JhMiSER7Y5E
SAk2DCOYbN9hicPDMqsmMhXYdUmY8/rOWuWlTRSEd6YlzHU3EI7KNUe7eX/DovAL
IjyhKpSR3MM1FPcf7xQGtYXFXU5bkTzgvKEctqRKwiCd62LRqhn8f4l0LZJhSCs4
JcCvSZubXLXdvaajAoLYUfaapN6xc7Gi5Yl721peoPJazz2NED37VG3yTAIm34gU
g2iiyCKNErRWb76z4T04c/0fKTWTRBdUSpWzror0W7AFxTZt/Ca5NTpGVvz8/u5Q
t8fHykiRWNB1wKaXPlXlfNNI2ae5RpWBy7FX/8++nv36cNBYkEuBZkclJDj50F8u
+oGGfBTYn+v4uxIBg/zucGGRElAHqQCnFIQsKW3DqsX/jYIB/PYvDlEFJxM5caZ5
w7gzlhgcjP4YCtJc4Z2/ZqJEZ+k2BwHi/5P2mxxIEyoJ4g4/UWMkoVjffWQ6xgot
QT9lVcp6nlAmXB9s3kSTKsBg/+wau+UwctCcPEDrayaD7v8br/gek12hlDLXUqp0
GqyHnJc3XdlPsCB182suy3jENrRfJcxY4MHa8sAzrV5gUjK40eduAFDJBEj3be92
eWBdY33c+Y+seQrSoMdlnSZcm2fHuUGwAG3CrK2Bgp5O1sRtVpn6SEnJCqjK4B4R
+9ZChLGGNteAprdm9tEdMe09Vz6x/r+82CwQbCNn15uZQHfeBAPtStAACcU3fpsF
aEAhzzJKoMzxHP0kD87qfw==
//pragma protect end_data_block
//pragma protect digest_block
hs++EX1k6GFAqVEJV3I3GNq7Lkc=
//pragma protect end_digest_block
//pragma protect end_protected
