// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KsK85jblFpdrLF3EYfsHkds4cTwx4CsrPTcDcF+4SSa5JfQk/DvF38yCpPZT
P0rL+f4YoXevm69nCjOODvjZIZbTA1lcbiMCXaMPS4XoKFkSfM9qWA1JKvRj
n0V9fcyBCj1LJnC6ad5IMG6L+Gny0tVGVSYtU+GTJBpoAD10NxC56emLZwVe
FAaKIJFJJTYtgwLkCuhnH4ML5JYg3wKe1NAGtOoEKPuz1szXncqyABd9khWn
RyAv8Si7MvF9lLdVyTrfPIjzphvxN2rNXoo/oLqEBXkShZiV//ESdSA+8Aew
NCI/b89hjyK4Rkwev1/eIXKL4KW+/uAMbEOC1/mIGg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FTu2v+Yh28Frx8QV3C2p1Pqfn4mfAAGxHYUCXuOaYwlOdAxvB9CaH/O5tyh8
VbCrgByTD1kNjKfIBlbNaeC9mA97CxtZMxm4GcoGE2Ir+qwgngfLHM+DD9yR
orM6GqewOdpy7BY5Bh6Oh+IFlOBMJNECz3XSL7uZj5E4lXTJRUaQDuUGDlXw
qAX0roL09s/MXNR1nbNAbpLU/LRGgZzEKyaudKGiqLoW6dauLgmS+wTLFax9
Va+/bdtK/rpr+kgBwYXwBmr+cD7u+2Y4cFPfaD1peiwi5EOz7LA6mX9gZ7es
aLRlNzJeuCnG4jkRAbwNJv3s9VKUmJcWD2u3GJ4kew==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WC5ihi5oAK8U8Mkx4eL6lC9LbrIY4GmWTfaxAM0UOZnuOPdzZ5znyJ/+6Qng
+qWwXg6FdX1BX3gJCriTfVlKJ6BI2chm+ONbBdL4c93N1pm7qVXSEh/uJ0jI
2Dg7Qfj/qNAJBd65/gJug5/VrK6zlZsMJiRvtlCYvAFonXdRAmCfD9nvlJVA
YQ1MspMEzOofI89NCLfUETHgWltGUTOSBisdX5lGUi0ZHxc8vsu2dbKLhu0Q
mn/lmbyfh8tgM7+4KeqrVBOvkCR0BpuzyhHh/gn84Lw/vKPrm7ZbnSxQtNLa
O5ZRaB86wlTLibqqNTC79l2sWe8x2V78dbQGgtb8vw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iCXX+NpmsD8XdptlnxabkMjZdRG6DWWIT57oagzIP8aMGW6VjcUCA47QzpFY
AKUuQ7T5ZTJaMG+wWsPOzqM9eQV7BFzNTxCHwzBzdftPCPmjHqgE9u8lGoZ7
jAWqSIQqGb2XZyWnUk4GvlXxmNdaimDzQPIX/JlRnGmcSVQLfck=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GP77nOqayDC7bfG7h3oXsXhYjCHIE7pgGuVhOOhWKUkMOPM15KSpB0tO6K6h
o3gpbkSuyhE4YArH18ycqezR9sueYbEUsT+ySLd2+Lt+7K3myf+NyLZB9mu8
80Rz/vHWannzXJCa5b0QQ5e2eqfLK+hbHrepB9mmlLjY/2O9UF3Ll1QUq7B1
Lozibk5vvgkfHFwzh6IMVemkBYxvjVKXl308lqAYLXVSvZ1hoksWra3RMCzz
HQljheuOxHN5y3Pq3sn683YyhIv5h0EYjWTAyDrIYueMHcLKmGedBC2iOLDX
Cjn6VrZR5ZcRH3rUXCYVIx1CCmsdNcb7BnmUubbGjpb1DrpCQAWZSZpgs8/P
FkSM/vxXVZKPT3zXERx6j5VtsHjgdLt6XKQsIvT61p+849yTgN0Xj2oe66X3
hKJvc5LRwnV7l70j0znvrX6kZMoDkWf3nYKeT58is7kwFSsdSAb3kVSjiBPy
t2hha5Chi78RUPLsCtNvcwe62s5J0K5S


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QAax7EW4zEMonsOGlesUy3zlzhxE/vC2UUiP9dhf62UER0Vm0GZp+wemr+qL
R5UPAScOin/+OUMV8QnItPzO7sI/sc76KmouBwX3Wnx379YuCKFTS1GHJcEw
3Pr2xLvmrfAsOBx0NjHSmF6k4YHS3e+6JHzA5QmXwchd61WJv7o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pUZv9cQOrT5EzV4oxcYfD/VSURAnYTvSPt+thvZh/c3iBtB5r0v/8WOad1ik
IDmJRGPuesIAiQhAQgHmmFI2xfTw+YxYkJAqZW3cyTKWOvilU/rSW3uhK4D3
W7J1FnSiXVud4UxTkPVJguY9xcq1ZTCeAiiSTXKb5R/Bl/QulFw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13184)
`pragma protect data_block
TAPUiFOKOV2PLq5OfOaDH/Noo+NmFBTyuDmdf9cbi1NbFSeFFpwnqVRI/AzD
H58VBN3j6k4XsRTpP0HoiehSgD50pLrQWLcsH6HV6PykXkkv/VOHRSoPwfqP
ohGz7ZqYEZwuetFr5sQmD3VM7qaw6cZlW1ZfX4Xo/vcBJdINdPolrNwkZgmZ
uG/lQ1YbwhJIxES5UQmsJxGl49ARPgBPEUCO7575uzIeMByFSzoToi18KYCr
13MRgSL0SiJpyJwlboQX5VzBQniDYywOIvWUxgTo7fJv0kxTsc25E9N9ImRP
uvbM507K/sGrxAze/z4/e2n7bPgs0e1AVUX8FWfi4u+hhmWEKx2IaBUs9/8n
p14PVzVM0b6zxJ8ef8JCyGrKXzsKFAqTFAKoADc7HiBi/BolQCsQNp7BHMgY
tnRcxiRPP8uc1ws/PfC5V9KXg5oK6fgVIVtRTb92lSFTRrbXkGf38vopuVMa
TFBF8QpNnQiu0hwHmkf6HH1kP4xx7ICeNgXQtUVLxOeBxxRo4R0sYOG0Tvaa
nTY0x4QFFok/HkJ9Z2NMzSrGEQCJPQFTBpt+kM6sKpLH3cPaXmcoDMv4Qr1W
se1QEo23BTE73AotYmxExTmhbCQS+LsjQlTtxELDa+J2F6BECX2VYYvJ+eZ0
B/DEL/uhfSoKDjyydoqzMbPtPcgQtZDbwfzTIjp2iVnM4xyVKZUkTOIGV2zl
jBDXTVHfXRNRVjXa2AKn6xecSzQlf4FQPkrTralU9CD0cidwR9NNpGmU/Wf8
nNKXyqPpiJ0ydQmcjNgwXTb143KhPJfuXZnZC2PhPOWH/w1V/DGjn++eF5Nc
DFaiYjOeo2ePYcXjq0EXtlc68NGv+/UIrMHmOF4gTOurrfYQQeWlRYCSjnUd
fY+MFVJ8NUm8TijOhKtjUaN4DjdWhMrJRT2wD4Xrd3pnK6IWAguYWc1RxkZs
xzac52GfaZ8mfv6te+hW1ji0vD3jk3klEb9N9cK3H49QNSUYJcZ65KQr8QhP
Ue4vK+/xWGvVQswZDctbZTJys/QHUs+oXrWA+zmfNpCFEnABHoFVdN8qF57N
pauWXNLoeX9K4dsHVGKzMh5/xHW6fnhXEuS2F3Qsc363kA5Jx6Qf1Kc04N52
md0VmnuRNI0KfLgmMDdCLtpFlv1qZRTj/BbDDDlWXq9tLbSYIqrPhl2mb+pl
Pm8afPcNioBw/UhD5FNB6ALVc9qACBc6Gm4zBPNrYv+9KyTXuDv6VR0+whC1
uGKPWIKGtThZ8GVsV5XQd+aRVocYIFnjYklAWRBUkp5dTEuBvISx33Ybz+cq
o9eaE6haLemv4iHDVVKk/lDUW1ti1YBTe08MY6SGecQ/Dvf+Iaon1RXphkQi
uYhpBkBK+L4zqyqCMF6ysHy8xntF+0cZ+3i+Osafe0585HjZQ8fnSVzuAbtT
LtRvEu+/SVhpHbzVSVbbxEaOGQB5cVD5YCIgtCsLm2hTnmuLJkK/Sc/+XWdi
h0D3gx+TFZNyKeoIKLGFZxxXjj35QVd3K8amvxSpD4S4h40qknjJLE5QYxpo
ny0DS6kXTQKf6W4uccehOG+l0ZTrFsX9wB7YABdqczhj6sOXnEI2Yr1ZHwXQ
TQLsdrY3u8NeK5pSJN8BrUt7PKz+7Q6uQSvw3XkoAvplmMlIHaRGzN81GX1X
NCe3dqt30/6whD+YOhiRi/f06Eh0Ibi/2ufnCASagzqjQcME4+IUnMN2reob
545WgLXt/aiVlIuGtlmfdkGi3dTjjiWu4LE8D9y93VtWU+Ryn4TwOLoKk0TO
jSzaJpYWLbDcyJr3+5/FnpDtjr7vLCkVH2njjjQFw0iHkifP5VQdSBWZQrQW
6me+xdiK7xQaIFJOgR5XpqqAxpfrQm9kbqdfhs+T5GDZSw5wXGu8TMgleGfm
KgqrFpY74p0yC8MVbrMf5tfWkm4JzLhJxfTLtFENnHHJkZKp8ixHy7cSjc5J
SsFEXRKNMzZE14/h4hRbO5/ErjVNrDIqVgHgFdu/ycDnB5nAIvRprfqiJEqK
6K1/rJTTM08aOAoNrgFDd8/yfGztYLm7cZuHMTrvOU3nzxTAhG55nQrSIcC0
yEvzVBtaXVwqVx4/Fku6C7gHEXYzkkvwcKve9prUHTkC0IMujLlBJZQ13d42
51AHmP59r8PH/dK9kYKw9xs3t7nyinu4dvE3Idq9BcNMk0z0oqyZ+6fPr49T
MsE0lbLo7Qt0l3WFjSBDYPvh4bBu3xf3I37tpys08BE8VJmUblSqvL/HcJ1G
c0ONdJLZ7+iDQMpztX7qMYtfg3eiEcYd5K2I2giJDZbnb0Nk9sLILEwCL3si
e93cibPBfytQGt07Ym5PTo7V47D1rMQRT8FbQY204r4rXKDYoVpzzRxWvw3m
JtqwqCwYma+z+RcSPyhnKwPVwcWL5aFVmK5t2MjJ5efsy3uplHY7o6roiFJ/
Sisr7CaQFBsUt6EtNdQisuczmSL8Yfs3eCvIhgTkjV80ja52A7OOoBnnPKV1
Gs3aGKHC6LN46XAVuT4DHCQuqoWVJSaE5zO0By8oypfhqLEOhbPO9V6LpSwH
uRdg1QXxemlYH/NngH8vDs0X5JbP8O0pnFdcjckn4CCiOoRKbjJFKCDTR0SK
U7RXN+2TSKH7JxOLn/o3Lj2ez0OdauscyXXZzL+j2T2bYsJ0bWNnsMh9Wn02
8X/uc/JAn+KQhQcoWbAtVTSjNtaODOjHW+UBq6GxFR9uGzQLCouAKwiZKX2H
kXgx366zaIpZSYhabMZhQeAE2LHHzidxhAZlBgHOdt0PZ2WV+c72BCaTwRi1
ddgh2iBQOBDjosn4pHWIkDcQfn4Bb2uaWdzPJZXfImC8a4E8iJlvHRA5l0r5
omoAxhnsfy1egqMp3Nj+dWAQ/xboQTKY8kl+52Gzg3/itmhBaNAcIjJtx/jf
CTQnsSOy3aM3GvxwU3BaArl7DYlRQs8JpdkyYg0hoHKJiX2j6DTOEzo1NvPy
Q8Bo6I7q18q6yf20sacfN4p3dOZABNJv3VbiyXozAcMcVImm6rAcwvkPf6Q8
xCck5eEM5CSx/6y5ZKIKBb7SamWYF0+g4w2h7OY1Tn6zb+XWBVXmGtdXETfq
KHz/NiEs9GhRtuw6NELwP+D2hq/XLOzkYfRXRUU5CcAR5vhWlo6MCFaNc4la
O766xww2PpLFUtloexCAmwwYRzul/KVa1fz4bAHj7VfVtKSy5nQGHZAAq2ST
/u2PjlNe1Vo4oYEi+HZ8lxf2qgOx+WRPEQqgNH5qHZRMMog8IK2VmLesxixG
7Wzuf9aLkMHSvCJYk8931B85sZDBEGgLyrAhmj04pSuamq4E7hPpyqDn8rS7
f/K14yofKaP1o9U9elMFcW0JHp/Qgj01SFb0lBiKdO1tEhI0EHtBK5M20nPZ
RkmhYYt5E9UU/OvbliQo3pJYViR0Bazv0aObYaJdUz5rbfuFTfTuxzXOY2vU
T4ZAMXMTtkSEm/JIQoRRcCf8bMVZSKD7A7tCufZEyr+wfm45ptFXpx6PUQGU
SMTWnVlgMM3RXMB9umEpwk9O8RVjto50+sTXniZ/zbMjtJGVZ5JT0AKtj1un
p6yWK5UaEDWX843Voh+1slwq7+HOHM/V5F83kE4tIr+Kbg5AF17SVBZeZFZx
JnSWmrvqv95jkcSXXdgi4ntaV9BVq058FCwloxI0AkYs0d2ZTnq32jcqAXEY
Vf5ZSJnkO/CUP8m37W3rvNIoMPt3jifCjfOSp6zb2784S2uPO2l/kNR0LKoH
zhZJSYC/FQnRu8Rmeoq0MK6nMNMSEEGBMQjSmDoWFB0NpZJ1mIxVWt9+owCr
U5bmVs+JJ29or2NOR+fIAtF5lPlIIiyw8fI5eHKeVaA9zQj02iIhVQc5fmn1
pRuphZ6VvvvEAt43sxVcf9sf5UTVSKaGuefwwHbeTQtv5PrbnGn6pqSG8Jf4
6RRp3qQcXFiUKBJh63UNhxs51981TnNN1MiOn3EUuv9+YcX/K5vrosPF7OFd
hHzC3rRE499pWUe87niCkQHRNFAN7rImfRe9dEoiXYZWRxrCUAPWLY5Y3DW7
GJbAo9oT/h1DjjRwRmpMPEWV+XR2CoVkvI3ub9PqL0khdJ0vRUXC2XEB2pI7
dQpiECLccqXQ4lx2OLNgsm01B9EM0rCXj0nX1ByCPPkRHJEfj2mR2K3f8S91
BHZocg9/nTsiEzpXYxOGHLFCyeWyeu8Ia8rJfFWfFFArDFN3jYgPlsI4dE/g
wjRf0KHVUgw1Y2CiHVROpEB2JdCuu9W0SIhrl2FzTJH3WS/sM+JKBFir7HBx
onWxGHcRwE5Lg7qhX+sqF41Y2tYc+S6TdiNFq3UtmXD9Oc1iae/pSJ4vhfvT
yHQ/AbChZOR6+hlcXRIm129T0ZFUa9cIgLT8sWf0Ux/YPbLwJcc2UdPaMTuF
L+pK2jFBw3eVtPw+j7se1dwsxi/XyxJQM9m+KUGiXQ0HGvMSDF6JNHC+5wkq
5ATtwirIZazN8MSLwvivgiylqC+oKioVvHbsTV39ZPobMeFFmxQTNwOV/70l
Fa4LnnRutM8eSF4ulbUKfQSJnNQxDtza0O0u21HtlT9HRx62SFajtqkljOXt
QKpqVm9BA4xBi3ZOTLoHHyeadaesROdCYqIjcFxashRwmaDS+1/X9si7+ReW
DMSx5wRkr82qTNQjQHimKTW8tvIwI10YmmF1nQdx7oVXAzEq7G9NpTPMdEsr
5NkTrObpfs+Q+Pkbxo7m48iFpj6LLWrdE4Xuhd47RM7Iu4Yx3s/MV/yiS3lW
KBFS0/FUAAckWhRzsBGP2RnXdREf93z/4SMTHAl96eKa+OUMfwDyBZcALjrA
2aT3U9Rc8yHnKnAOz5bzVBZNB6P0lR+E9NNEtinved4pAmlafRjW9CV1dHhY
hse7g6XjbxjFSKd5SIoUZ4wL8G0SC/kE56966B4VEzCdqRJPmBV22U6vrGsi
fJAtwgqn1girzWJvvyRiCLoQ1ws734w5TX9TmyVOpW4oI41VcX+qEZV3pLu/
Dxr1PPu+fN5eJ5rb39vq8sr6o6e2Pdd3YJYrtTDMsQe5XfcdRPb7D9sFAsKP
r7EMIMMLzKMNPukaz7IUWS62dLHh92R43NYJVOysJNg0PoPsNXxsSt3uh1Ww
Av3qKIqU+rGGZfM9c1p1JYcmdS9Msx7eQMrp24Ew42zuXumt9UKYUePge71G
svwmD/6hAS3Ra7Hqbkv9my7rMVSpFcwz788FmhnjezXdbDjP9BlDY4rd+d4l
KCX8J38thVVTxRcYWC9UjxBrOh6lDEMA/p8OM1HwOhE9Z9kaAwbM3t9T/bu8
80XXOOJgMM0Ocd3TsA3lB3PvazwR1DyEgR+iHqT5uOwbGyaOYdXTdTVQhl3h
L5CBc+B+3rgubPmnp4OAOeCmasMZtCQ062pz7DetOhlL5K8lowQ0837wBlg5
Vvk6PdIvSKwNgZ7Hym5njysFUz+k78YkGoZ3pnEWohlrIO4msB+q3ZjwluWD
Im2HTPJdByAp5rZbeAXWy0oDcymye51JRv2XWsqUlkGjZQOImG2qAxbOGvjf
5G74qBMp09q2gxmIb/WECh7MbWtHho3N5FFgAlgvrlIu3ZR2kYPh4c/ZyGK9
CvPQgD9cPES3Iakvc5himi03kfsOiqTihr41o6ACFb64HVf44VFC/L6yiEX0
eTQoIeVzysLaAVQQTq6hvldirNxrtVWVgsjDYEElCOvG48d+yPbgm5ZaTEYz
Ys7neBQzAOwYnUPTGaHlcbaGCpPNaTNE3UShkSnqmStsXEyfX7h9/i5AgHMJ
ulPwjrlzLUVkJyczm9FbKj8v301YCFisCppG/jAY/3tP3HUoCTXz1C9l/RKV
ZGsA1QMORlNbrN4GVXdG8VUR0ZKzmwzMeQx0/EybG+WcoGhxntnpIAnYAmLE
Y73nMlVbeUJ0MGmYxv5OoKO48m/PZJYH1MIjFYel26HEzoUdtxsKihOHp3Xy
tBhWS0IbtFuQxJ4HJffFfzXZGeYgULXs3tqjWLOs0c7BrU3dV07MpUBQd32z
aI4dtFOLQjwrqsUUi8xgdAiNct3DxDcq/xWMylQ8+RI4x9P1pyJUV+sr/hE2
aMFvxpnVeaqgRixZ+H9NH1pYwGhJlAyDf27wp04YPuf2x3SJqaEKfCMhJ45F
xd2lzq9njcA1F2BxY5cvF9KDZgnL7To35tpxRO1ECIsBrXpwkCFQBnCP1NZ5
yA+2F53cADzDLAetlnR3ispkDijlziNk8yTF5c8iozqXZYjX0uQQwgzxpGij
u0P9p5B2N5TQYv/t1g6ksiNfQWCKBr6laBj8XP7i2h3xolzX32/bGFbVWwIi
h4sLyGXVnF3aZVE7prx5SHWbTtCCy/hKwia0De5a2IQeIA6aWGzrZvZvlnWx
7DVuvkS83Qwpq5yxvPWM25Ag4l00+qhiYemJSQVINibfr0gcSfEBCwtNqyxT
x/KIrNfCglXt4DuPROxN9sc18qdFYi5IHair6+FgeDonu8TsFaVkBIprDEbZ
sBmtDRtwQfDtVUid8phPPjhhC5T8ivdpezjufS/qO4rq1o0Ca0YxYgvBkmKl
ifUvpUks2A1jC/4EbEmBFEWSWi+m9KWlCKjZ+s6Ob8xfEA40YEalABG0FHXV
cVXj0cOE2EE0Occ3vMUGU/RloKxd0QjKWIvAjQY9ytu/KRXf8HGe4UB+VpS6
cSxZ2IwUYyB/XbgCWc8BMqhAHiPxKCITEardWJx4DVWy36NzcgSD2iB0jX+4
ggISYdoCSproc2Gr1bOiVsfI1eqmS73CzxvqZYeHScLcknDXXNixZrPUNdrc
do8PYTA/YqkEaEIkfys3aKrCueEo8dIzLqOYwdOWKBLLoMHka+XoHrzYmTiQ
UjlM8Ya/kQYMKgWYytNGbietdMHbgTxSyNhAAGFc4wsEmD02622ndtQkNR54
moFr+epoPmFTyOMdrIyHBeNTyH9ygMwZuaydkFqCCljjSitPWURmvVEyPeZr
vFb/jQJ2tGHmADtwTFkdz1ZvO/KELn9YDZnnyUP+iC5zRkPyxJtZobBRgOE3
PxSuGXv0tuZNPufvGBN+Jz7vkG4ih/33fNR95imyajkJbt6u4mXteFxac/7E
NAmzlWGfVWfCORVKxANxBmc+qCcOyUefjxOKpFBsVu5ZiKlM1roeF0BWLQhK
zvdZVd2NpUSUEDAiHe6jHClLV6jMpodDAcAAP61Y4NRjdawYWosL0Q6bIsTA
8K93rzJ5/lRHEyxGX1aJSVeCni/CyoKEqX/n/jjiqYIetzJTs3qLC/aUDgsM
h5pvRWTVsox9fzJTwhE8vvs/eL6/RMjUADbZLjFt14Z7UGTPI7Nc4ZEP7D5E
4kSl3ZKu2dmk/vo/fGFwzXr9Au4XumuKVZfVbkjy4Pc9nCGpzR+AhaATEo0j
8aVQNm71PZTnlZSQ+9fepqEClZlbfz2fHQh+zVvHVYwWF3hbOG4l7k4Vmi+r
CD+vApbA2MNdTjIBCnXiQ/jEY5I6y9A3QiaoeRPrTrUUpd9S1gcnVaCfIcFp
xnHksXGS+ZwlEQhQ/6XFK4o8AmV2LvakkVAzexrVfRYhuGSE9T9HN3Ls/gEx
BJHV3OC7hx3jf4IDrmmYq4l26Yt9OetmkTzBsSKEmgpzTFs9Rog/eurYvR2d
VrtYfyy/GqLZiFWNxMBsk/TTNAd/16nnvB118b8/BspaWhidQSs5+BNcBAot
TAkmxVCxsRTjA64H71YV0+ChQXcHp7AnYbzQSP//sd6RV3e8zG0QHXXevWCO
VmS3z7Gu0jWNWBIq7y1qsLU1QUZScqYT04VYwTK78ABqPtcnGI9fFOKWz5Wo
ZBdDRCwGcABJd2FGo4xIP3yJpqcTq4B3M85Ply3VIbl+/zOzCJBIlZzSft3i
FoKEP5JcpW3XM4UPC/OPYjvCdWelf5Qc/9qKySAFVhqotZhK7ICPOtQtUZFX
jbaDEJzeRDkf406olBksiN26MUsIKSOCH9Uf3XnpHEBaxaYmVzDK00tbqfHM
8ixJ19YlVUFDd/i+EikxJNU6k92CPOwlhaOE8JId2VpmYvC5oAhZdTHio1GE
K0dMlpDmz08WO38qM6QW9DZr1oI6R6pxRiyvDlKnQMse1pYcpacZo+RG+atZ
ybj3CNybq1fQ+fpCraiCCmjFfNp5uNJMdmsH2XdbikzzN6F4HB4/+nOVI8sA
EQcWbF1AH7uIIHTVjQi2CvbZS/rf1XUjDzMY/YYaXRpsiQvkD+vYgHdHHf3I
84St6Q17ryDgJgQvU4qq/ZTkAXKdxYGVrZi3MqYDSWYWu/cWq/nVFKIGHrR8
d6GBbJJQ/tZdjMendNg1c/m4e4yHivFG2mloMs9DKO4dh3XwB5tasIxsQ6MQ
Ox4b7NB0h/sGy9tkcBnTNtUrHl/NKgKN4ISz/uDz2fg2oWv7U7FRyQwfy+PH
jVpAVaRNH63R75HVfatcB7IwvD9EkrKcxC568dT5RYpGIW1l85UM0tcDQ9+c
Fxir5zpsE2cO5+zx6720VZmcWD2hAII+xx0c++N/8RUMoXhC0+1aLWP7WPv2
bsScVo7feFUbOdmWpU4aDYvO4MxW19LT7vQ+VezjOHfia0MkUFN9s9wukx+g
jNBuB9VMnrnB55zTUMQRYz2JgtQWyoWd9oRXGeyepIkl9WGLAcD3oak4YukH
ubXXVsL7v/HYx8KPCYghVZr/GtlZQM+2I/OV7b495zNcPuJtMwmOEwnGMVBe
h7pourUfhZ4z069FGvnMZevsPzAx1nnpDbQ8fxgpWnBUvtdPREelgfxF/mJL
sJ2ZA19z8GmLgD8xxo9184l5TsjrqTpwK7ECGHMZAgv8ugJN8H9tNlSZdVL8
cf9zg9JRoYgQYAL+RJvDwnSZdLV0+YNWhzvkCR44RMzsduxjuRYCDXv30rfh
xG0/+RloDOVNtE+fChXmp+Mayjl8mOLEd3V5gupLgR7XmgNeRiH9ztPHCz/X
plp4tS67bpmI3ehUfB3gML4kc/l1YGkoqVybV4lvKeqlEdEseW1x2cjG72fI
ODIg51a5lzJ+rrXscW2TZFJdDYPulPbwMWfOvMS9rrTeOFsloS+9uerAjFJS
y8NMRnhqlxuck2DJ2CkJqDbL7VxQhSy5JO+WRN2zss/ExJV1JyvJ4CxD6Sp1
h1XCwEvDBV5Q2yvZG3+Y8a2KhlbgZMmr8zbdpz77mcX8jnFsktDMp/7St/14
Vv4gVBlczDhTfQ5qG47xO3yfrDn2ekpPsk9p03+LUaTbDHPGe/M3FPrP3xns
3PiVMugfE7n1Db7OZmgDk6laii7chSL/4LOLDXabfRNkEE6o02UnB6XzPlZo
BxNZ36X3AUPpnpykFali30oqpjedyiHpV+TMgHXwA8mJYyqkvH/Z5u/aU4nr
0Txo8ucr3wpK7vyLE41vFo5W8Yp7tEiNYQoj3eByyau8B3szzr9okrZ3kgiK
2/Zco/wMN5krwNILOVkj8aBFLYvzyXyO9jozWR4khSR1olBHrHsPh0IpHrTj
ANX9+tFjax8wX75gDDtdXS95GsOYEqPAQaE3AL4zhAZVCx72VMd+X1r8YBB1
gLkOxEn5WNEEL/0SGTkaIUBCHZb687RDEK/q7bdMsg7MyXNkqQIGYqbkz5Jn
VR13RDMs8+iEqyypHbdBNN4vxtcEzKvFd5f/XBTeQw1bZFGG82CKFT3RrtiL
IYQfDMNOP35jNTSEFwBxq6DkEZR2Wz83YnjXM4GgP+Bu31BAWWE0eojGuxh/
zOu5JWN4snQRl2GYGg8isqq85S6gjtZhGl9eDYGBHoXh3kHIeGdVJRzfLLq1
FmCUngbf1DsNZhjpLvXfftBZCPps4w0Acj3LdzCjmSevLgQxkqGeYSvJGW6q
TX3dGDudaS5M+mY7Jpz9dwhXlYkaToSb8d+UxxqjLe5eBJu2tHAAEpEnSJ4y
dsnhCD7IOYSfOmtutVUpbJMQzjruvCtIJe/U/aQVSNWTl5dfmGB9djGDr9k3
GPkBFlP6Xn/BeJ3CpQO5T3W0xplutSD0JQZE4iL4IQQ9YXxaoGqwOEBxgEC7
/uVNpYtc5qu44o50IkgfJfeFMluyP7Zq4CxS6huXo9iX7d1QaYA9jX0PKwr8
1Ko9R+bcrr1wtsmd+q4/33JmI0kDFI64Yt60cCamc2NoKJD/19hRzpadyXoC
pD4iRzScebHfmw/lkUAelwgMwmXTK/GeG9McHcqgUo0MFiuB5d8kK62s/IO2
HtEXhu9jyptZFB7hWdb1S+onincL4YGsDKet9n+TtcBU5xZYfrx6PNbyvBv9
sqaYyFxaQVpxwxGUKbyXAA7o3YauV8ptS6bYPV7onaWYOCubXIjs0HDSVw13
u7oWJyNzd4xsRreoLwhj7tusdVculwmSGasYtvLCGeaEezj09YKREir+Z9GW
hKpdGPWUwu7uOSI9j1VuRbjvug5WRFieWDPDgxwrYTLa/vLyJBsxS7u/iJlA
5FepKkBvWfnX3Mv7ILUNEFL2iYm3VVt81t5rQpGyRuwW+NhpJPfC6/I/2nUQ
0H3GaBAQ5YBaCUNVdGZmIudX11ecW2m85eW5YQMk0q7yKIudmONgWJldvnO/
u/DObG4+cMYQVGIaWEishbytAjuexl4hPM14DM4YtaQVDrlPdQEReZJXcdLs
zpBEU5kfaO+0vUsmUta7+Q4uqnsyBTnuPrB+JibqQoUuHMtlivn1jjyD7NbP
OQfsgOOkGx6dswlnaMOAsW1vx0oxSuDNVqkfLmpHBiJ7H7h9gBhWtYX2c9hU
OpypKfnRFbVsN2jLS5B0W+CmmUQSSEKfwhhCmSPmdkFCaRF40hOg3wN7a2GF
MUDjdzKYWrmmptUVtpLOFxD5gb8FxmVgDfQSJIUE4R20rxtXfSL0FBaKY3le
OcQ/rdieJzdaytTku785jAU5FJ5OjEDX2cusYNK5IceGAH8D/YRxt3xCa8zd
gphD/4tEHMJortkFq5KgqeVo9+KPLnml/no6acjeOFdrm0klMrSEPOxQKzR0
8Mm8GznFqEGGzFtoL/8WovswC6KnEGRBDR7lMfkmJOJgjvgTLx7ImY7SjHqP
Sp7zWGYMPJKGUE0B0Cmvnt0nYW49sodk6d2QK8H5Xe6mC+7pLRO1t2LYQvtM
HqsfMcTbx1AC2J0hm7FVhbG3hNfE+Z151WbFTUbCn4cAWUROOzMOB2pkIYR4
bQLGGAUp3PVPlB69alEISl4Zg2lZQOvJrlcSa577ksPBki+2sQrwdfoltQbG
UbE69zEh3hd/FA5v62gVrHrq+Xj8dMFdEpajsRLGJBUTvsyNSx9DnJxZaWIT
TnbAfiar2nXbSm2F10vPbYEZRYhtchhlZHVEOMGf1FRNjAfKK5ACIfhtpi12
iXKsTMv8NFLbEWCu/R/C2Jf2Ycqhn48mo+BpIEeyYget5e5Sa1BjBQ3Ty2z3
oLfVw0aoMnh3PfBouAk9Kw9RSXtg52Gdiyy3/799xd9aT4G5E/ORJiSjld32
seAllbZmGuUcdu33YtIZYZr6yvTSoBIfx1pAcM3Hhq4S9m8tXB2rlsk0XY0a
3FO+GZdW/Gk/oUqh6fPH86Zll7xJwO3P+hgFJPf18nCdNEbS+QxkUeUwmenH
2DiTuacYitkNs0jlCaPT9PCnt9+Hc3f4gg5Pg+K5pQ7bg3gNpb8Xi3xjptzI
tcMjPUeQwN6V8mQj03AvvXtLMgclENYu405wMM3+xLHNu9kAXw1h4O6AhAkd
mqL/19IBo4P0aCzFCMXeX4hZLjD6TXupvmBsCfzZAAnw1vQyUspLtKjrh7Bp
uM9StqNp4n+/0BFZzOjatIl0rs8+cYM9pJ05whkpi2I30I4nod2g5kBSsRpa
lcLGW2wnFUxAs83DKoZyCXArIJo4q06KYHKBrTiLSCITWsZUQNhH/LAQ3nFP
HXAd0oV2YP4jJObrNl58OmfOkfWswttKFc7lvzHs8CAELTUG4Xqvui8fTfG4
hc6SyAEnz++itNxH+M8gLWrTfitUiywphuJ4Ncas7GvVvxhXGHTrUuh53/Gw
YsuS1ne9jhjPdisqlNcZpuTclsIa9Vy3Ra5oUZyq+pgShmfOh6wMk+g8VDbc
ZFWYlz8BL/3FpkbDD8ex+G5o3tKxz8IaSGsqInYLviBGyyPO6aq9dfUuicPe
ZyXg8RQtnbspx1FeF5BqtQHzKNw3piia8twHyekNzpZwqasF61HpWoOcrXdu
ACCO11RzHU7EEsG/1Wm1yT/XzoevQHUgBsudsbFNSnnDiyeeW6b1Q5SU0ow/
O7/f4GPsxGL4FHORK9gEinrin+Ak6tJN1dcN4hgEcJW/le3fLnTCP01QEy6x
Xln3zNKQMBVlYSqc0NKVvIFq6i4MztV8OxiOkmfJypeVIVWg4DuI/0E2FVew
+bepRbi+HrBkRcI4zcMdWblT0CA1J1p9eqDCWZOug3kVPu7mSIq9Q3ZaeJgU
d9HBAijhh7tKxsilLoz1BFB0B4MOvqfhwx11A6DZyhP3fG1n29LUk9DkxJ+5
U+AuHuMijQ8Ge8MnjYhBSdkNjV4Uwk59t6HawQrU7bNeWhNjuF26ND+yp4Mu
CH2gFF8+Xz7CUB4HyrMKCacCU621kJ5pduPtU7zM/Z1UqMIGfM/eoc4zzP0U
lJIyKfW5lJMfExv3GYW+GPCpLcv4qGAcijCi/c5plZ6422jerzsJxdj/wkzD
56tuLy+EL1YxIWy00074bMZaILTk3C9bcAVPghy1lmxXCqfGbnZpNWsWyZvH
ll5p1OJ+n2W71j4FczYy9V1duH1wCX7pFBR/ZHSEJ2zUF/pKEy0VfF4cAGBe
2Dlmm0tUnm/eVIgFaTqyqLpxmw0wLzrRYyFj8AIUz4QQgf2sRstB4UCOjBgz
cKHgzye8cP5gmg+JlxXGT2lk4UsnWcjp8SH+b3j8x7gShuEXRQ08x7oBxTQH
k4qFyLUZ80TAP9avlOo2MhB7ZWXRUu/wCSRAS9BJdk3DkRzJHEHvetYB/Fl7
nZ4G6UpgjytDxw1TI8b9prtlOGeX9Uaz1aO07ZPzh1CnWjQENxFY6MGGTTns
bxbvCvBSmb9Vwa7PNjmWCRPMP01mCpklAbZqY6qT5zpNINhUcSqdEsfeyVkP
cRyspRKinF2y0jKeXbmt1UvY/3A7W7RW88mJp/F1KAr7wEQMFMUE/xFUOJ8y
Xs7P+Wr3v1LBG6qv3cIAa2vnZK1DR2HBZADE28WPd/jLh7mzlqQ9Wjwlj02Q
MptPKUGQDvODM5gY5lbKUTkCODHOYqlgvJHljbSKcY9W2egMo3MiWEGmkBNJ
DQFUce9AXqG4dRKfmVS3l2gPB/HhXPUcTqCAw0Of5ZoleboPDZN8N4jQWxnW
FPKnCnJvQ4Zy6qMq7FwzyH1QPXh4UEdiCStxxjC4VO+XT020Fzw3IGhTie/2
pGxOEdT8D69qvQ7kdNsZbIMUo47VO0xKwp7NyiBGTWqwdVfoXUCtCExmcaqT
Rjec1a5xFJc86yPNB/rav0aIgmv3cZ0HB11Zo5A/TGsly0da2x9K97ct5Ib4
f8Ihdc0EXqCThxRTXGIJGrUgU5qHNjpOuFxpV74aym37ck1e/BCHv6QFrWsb
02qKGN72hfcD8TVxpvhlXliDOZjx+D6UQBvpKqW4vAXh8lkPVqVtxLgQxH4M
z9XpKfR0CNUDG1Wr/kOuMVDo9bVphDzWZCkmuM+vwpyf3UVI/Bn9/H561mGF
jzzf/XYYQPSHjgaVPfcYakfxSK4JGRGMcxzjqsgrqBz8tkG0YU7AD0tQx7ha
jV3D0K4eNXGIVvgZFWBKD1Y2+iVisi/zYo02gxo1rQ4zVt6R1XCSbfdAJ7C7
dzShoYiDgzLsLDHQSv4e0PVT7kABb2By0EmImy+bEXgOiyW8v6U632sBD+Rn
GQfyZ+89Hm8wzw0igHSABq9yRMp0tGibkgPdcEx6W4bEMKoEssc6d9+zoWGY
Btzcd5/K+p5atrnr+AyQq26c+wE5mcwYmn4NdEhwe/v0yAt6t70ToiJTPwLv
D3+XXu6Aw09Ci0KYGyWomr1V4FvEcZkWHD/91VnsnHRGfNo4mP46usyQjx/J
ufL/zxEgVHhShpTjCffYs1gsWeriTz1UI7ciWS1uZODhSPM4uCR5El96uaeA
pxZBwlrNosokkfpQ/QcbqQI7731+hyNv7ChRgsEyjxQXjV/ptfHk5FiXw/rS
2ezL5KnBhhZgcxLEXOHcBdZ0E1QWkI5fAYMLhtYy6e/VO2NVkOwY4XGlr9Ff
ml/hqfpp97Kgcu9/WZFhrFr0IRPVzMqYLjr7Go92x+8u4iKbrhgsTgS2zHVW
HqDQaewOTtV3EjBjSVh97f1ir6f1D2SdH/t2Slzej7r10y7XbS3HsdcrAFcr
ep+Ndc/7U66kmnBAUk+3b732jIzNjUnbYwHWctI0aLn1JTwLmqRRT3TdRSN7
Nr1Utb2e/QAfdSu7wRkbUQT+OdXv2P+zlPsXk83mUohkfr/zMkbZUHiIq84h
vb586KtO6tDVJzCqncoS9TonEYfasPnomhBsSXOUvd3O42xIlhNJEIvaa2d4
FBt/fYjTo+oD4UkNqH5pBt2kuR1/GV1ZBuYjowcdANXuBIpJFRJs5sZljhFa
AaRkECzL9dl/m1NefUUKR4OIJo/tHFoFVTwokUCEjUg9KfFB8RcryZaIzlBN
Aa6EAcxUCfBQiTc0oFyb7RsZXzVXRSsRZHTuP2SGKTZ+Zn63AS48fdyoLwL1
XdkNwEThCNerCN/M+R2vXXwSwWjTUGcnb/Cmk+jzafhRnlnzkwaSpqSsC/Md
iKFHAPreny7Fj8BwEjcKETIKL2bbqInagbcnu6R1WplWhJjxP8WCyWrpWCJ7
Aa3ii5bo1ZQ7xm0B/RmTDAHbcu6+6g/0gVsfmSfo1G0iSreb7NwtA7AXGMr4
jf49NJXCJkC/SpqnxafMc7WJbNTFecSzBD815/YiwGvFhf+gDsRwxJsEooRo
J2W4ewmSQtuc81N+Af8yGLeuBcyfdHQYPldPYY2OFDpXTvet/gYFbUhr3IKL
Xp9+R9Gl6BpDGT33UHL45rf4h8LCE1DVYLc9gq7CXgAzYZcvo99Dj5e6LJd0
2gsnpc1H3O+mTfNdLt+HBVPpyOLbyrcwZviK6fpLfeObHF67udHg17dMOvlD
ElmOS3b9sJWz1LMgH5FqAz9UJRdH+U5/MrT/EfA4Gag5CsNP7lEPFU1MEId7
6mZZddliKXuW6FSMMq1Cag+diQCnQp+831tdYGGSpicY5UQAflS8FWEXacMF
MVLh10VtKHMuiHx/CKXuf5sUsu1jxHVA8mtV3w09Vn91FUNOFcHvskp8MjCn
RSIuHWaEnhoeygMLMO0d7lTLQBi763IPpT6MJag9xorOltJtw+XDTnkoeasN
NNRCV59w+2EeGXAOXMWhnPsC8Fost8f1yPPfBmtKQp497e1ZLj/LH0d6s8Nm
AoySpE+Y1zEibZq76kEsCioLy4YSdZStg8knKcM/4JZrEM8gK7H4+ra/FDKk
1T8jep35tsX3E1mVq8ij+xBeHWek71in/9TOXqWr918ehZDBp4VCP7r/tdLC
VxlrQUPNBlHOWrs/jAirvEjD5tMUPe2aR9gxGiNKt7zO7VEKaO8N3jCZeb+Q
pHWYP8M+ywTfZZycrGRgJ6+jIqGi/ZP914CCG0OSeCixpUZ6fkY+alluGr6k
teClQouw9T0bx07ih1xPxEdNq1go7dULBIYQExlmkV5Zjc4RpPIMUJyezUUv
tirc44/ruR+YK1OyRRwgciojpAbV6MM8VoJHZ/J3CQPhUl0DwX0QCGvGxfsP
aDSiHtoKXJnTbJSONqT3b09Q7TLa970CV0LlZJhVsvCDtzMh6zwD5cSXBrSR
h9KT3IN+3CKDon7FOl2d/NuBdYxJX6JUJvJ6XrX+1HnBGWg9r101VrwfOfOn
hQZPkft0yuBL9nsi6J/cMStJPaux98+q6kRiUs0RYWYfOK4QzDG56+dhZkMS
NnelCdaA58DoHX2JMqrlvc5/AnrPKY3jclHXM8l1Bf1KZN8SWbHsU410KVSR
v2EnfpuzhnZFwqHZstwaW4ijoT2ROTLu7th7mGhQ1uUyegGVDR6IPa2n0UMM
yCtF8CMrbDP5gdkjjQbLFKGca8h/dfFNxWv15wV+XzfwjO1FfQ+Eyov1uuZN
kE98jqxKx9BtIx2N/P5EZ3CApSY2I4XZSKs7WIFWVeq6Y7TB22WtiAV3ClGK
6QNQpdF4ayQNWjHNsaa/KEqgkkqexkFpmi+keDQqqvtOgKz/n+ffEt0bNfr4
vVLZANMRSaygTkopHcphmJmOGKs911y2HX27kYZfPopIroSm5jxVtASzvQuK
Im8TKk1tZ96kq5RrY/GJYbHGHVGaj3+Amb/rRf9io+e0+xa8J3zs46sPFAzj
IBJHz+nGVk2MEf73R4Zs2ZkN3hKD2kbb8SpZz0sma0NOQYaqDuuPGbzEWgPZ
OQkedwSIMQQ3IkJteW3x7QmI6wUGrP+dlai+/OvB+Be3jTpA2exXTLY5qwM6
o1Sz8rREIZyXVeMmjV+ZqK/P1dPCJ3405cmWl4jyFv/GTmnakxhfbwy/WoId
i2ehvL90ur8Fh9XrZlPBFTxzdM76BzRHvMu7oQ5qrsWQQS3JgJa/fi5SKgF0
iZcYx/kg7kOHYf1gh1K0cm/LEJVD9ohjWRBU22qdvr+rub/2EgufGbkn5KoP
nAUm+IfiDyQ3KsfL891OlvB+1WyD+P3avC60EsldTXW2gb1x606c04EnJVNn
p+n6QZX7KXhRtfVbCfyb8GcDeq0E9P9/FSNGMZ7Qn8qFsGMlc4bwwyrf7N77
1eHiUTZllWeK3B8R6Fh9I549XJKRCEl0Sz9Rbh96c9aDZsbd8EaHTgpCAprx
W7OwYn4SqroSujc4nHfVsfybyQWHU10r+yDseYYAorAl9jqmPTDYbuHM2Lj8
sAPl4el4lu1iR8s04lqQXZtO2wFf8DQawLE+ezgnIUWxwcUGwG3c7kH0V3/Y
rs0N1Fvu/KUY0T25S6fsNvhnJL7bgaADoPtUBbgGNvUeBpwHYwbo6N/oZiWV
Mwpfma2EXqDR/p4yn/QySjHTZIOGcDYD6EN0ltQ9yXxrx1V0/Zjc7MXhHgnR
koHnvjRl2Z8EUnWFgfw24X9TKeyGAqFlsqlDnLELAv+2ZoQuHWhyRVwChfjL
JXgo4LCBqexxa09GPK3ANm7fedsWFR3cCI5aVrbvvqOC1lRiKeZ3xry9Zd+h
ZoPqYz5xOr3Q62peWbKvmHkKNy/35nw5yU7sqt3MAclAlOCKFC7oZ6aSunm/
P9Y4W6szQKIK/OYIJscrXm6o5n3tOxELOaW95yCya07MUxWtrlAHOnQ/wr83
VNARRbXLYg5hKyW/4k5xQAU3qrnD7IG8wbNKNLShQ3blctJAXktN5PaWHQw8
KJ2kwdhGwDccoPXt7doebcIkEVIfjJnghYT1r2UkxhsQD2nCBDGJSEuXwuDe
bwRpgV680U+BZ1VXe+17F9DkkRgYlQZnmKg2riTbLKJkRN7Mo8diHGIgolw=

`pragma protect end_protected
