`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
t4SdC8rj84Y0iw88Ex1dsbsa4Iqjn6SuEqCHIG8HiZyHJmnhBs1XOHUTNdMbT3d7
KWU35mhC066HCsldUjhdbB+vFtxopvsBlLZ8sVsII1s5hZnCswoQZPs9VUHVhDqG
Yp1LDc+ZFuDBL2OSfA/8KYPh3J559SVityZB8OUMXtU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 31488), data_block
a66wYJAp8cgm5loUn2m0pgw4wP0B33ZwmxyUlw5nlRNVnFiiC54EVyt6jcaHPAHJ
oyoyp8+IVBUMobs1Ox5IrNdxkk27e/wcVxa7BoyVgB0fm62mWgNw4M1aqGcXpeGO
a3jofD3fECKx9k0KNBCuAB2JSF2V2iXtxaNJjYxQVMeGcuuF1MxLmQw54niehl4S
OPfSbn6Wg1qxYnNkK/yY9PvqYVuxxMc1WoGyXiGNsxRNDrpmd/1CgotsbwQ9xbMp
OIvGwCH8CelGh5e+Wdd73wO9z26KglPgzy5Itje5ApXB8DK8R408fp3+VxQK4BWO
acki2fq+OS8BB8FsdLogF7E0nDOW+slI+zEKxTaxGjjraAZBtMCJknO/08dfG1r7
2iQ3qd0TQ9Yr9oX9L/p3b3UWPGJLF6Jjm3/oCRGUR0cnpNCWxlfJmw0hz2VGheYP
5leanxKYcnlFcbMA3ZyeHhODMbql0gp5/GniW2g9iI/5h+2mgg1yo7N1RkoDqTZp
SaprETWDPV+Cjs4lirUKKdf/7Jwa/6crEHNBd1vLeAeqPVPaB5so8eKnBd99MlBt
Vjj+RN+1NbL7HvQuFwpEglL3QeRPrEx24bJH16JcRRqkOcleGd88scpZqF4tIgbj
n202wqGjQ13yLHOOprvwYeceFCBXrRjz8neNKBaeYxoR/ReWYdUmqviHbIfZXn3+
ptw/kvJ3n8mNcNGjCfMnO3Kb+9wg3bBg0fjQ/sbRkn3wjMl9y1m8ioFvTctXV4Dq
Nl3954qdMFCUTsRhOFXQWHmKTrOQBJEeMysqbEuXfRXKAuBgOUAPA28pb/5/59Xi
YaPQlQcYsM/Y+ucgSgvSTvuKZGNRGzWlOEIIuJE0M/pSe0ytjryqBL1Hg8wxA8Sm
+VZmKYK7wFuhBTeia3sBDW15jbXHH61UNLsLZNCSAe37UYVzP0TSuX1+u6WNuYPC
1Zn/3afkjkzGGL9w1Rr8AIVnIYzBMqYzBjQhbB5HAgVCrgO8eCMuiKWNexHj27eP
hBzqKfIkq+0htq6fONvQDcH67IEeYEBv1q6+eiDnsUXUv0nDQDK1Re4yTTg11xWw
9dUpMpjK/Ly+M+XK/f+PeniDUQlG+o4AG28gVasn+zN5kQOreB6Bhz71rIqiVlKs
+XE4bHcCjluo3A0w8EJqDt6SyVc2zZ9yvmVKWHCUGzjFGoWtucnEOBZMUCxNUuFv
2PGwt6BWF+CQNftOcZlbBEZ5C+t5TTcoUvmiVRP/Kb4wDajM2E0OQ9MS4ZFFUTrp
GpqiAL0YTgXuL57opmgkWg+qxkD9YzFF58G1WtI9i9qzwCDu2BJ/6vDDWmqJGQ4P
VtnNSyhZjXytOE7r2gnF6kwb+d4gfPFnaxZlsc9tpi5qyRQoUGhgSVF3qYdLTTfk
Srt/Uh61nwzcxc6ovWwZJ4frRfYbH5QPE6mPLbMxBINXCsAKMiLStNiU+ZFWnZ5Y
zU/l0qQ20a08h6caQZ4+l2zWFbo0g5lsdjHEXgEZeUqOBqlJeQ639uDcYCFl9O3j
kHuCb2j6+kvxwYYwuW6Y02E92uYpB3ZNbu1MP/Xtiats6II9b2qA3e2ILLYRcLRp
mOI7HnaYWuDX3XK5cQWRANWo4mUQR6EI2Uu/iHmQl9LIFOWlPwDA0zjUmhu7TuCh
2oeRBy5Z6BGfFUM5AypLvMTda62RlsbTZaWTkKsj1adjISi2k1PJRI0TkCmOM9+b
iQ0dl6sm5qVoFxtm0J/I+sNmRB65GJl+Hm1CA8+0MkkG7Wb6GYmjswCY71QSIxhh
OKOklAJ7OG6oyk8VLB8W6tVlVNc8HoQJ2INX9Ka1MXC4Qm7R9vqrVhlczRzD0zZA
OSnTGuAZyyS/lTpm6uhFWmf4dvh9uuE+i21r3/Trv8IQLfOZw2DfZw6//aQkhASn
BV+8U1DgHph9Bc/7aEeeR5wx14uxpSHxXu3weIqjuUT8XtCIipj3Yhr5s+1pyjD0
71Wo0Nxcw5bPfWW4YDPg5e7XbIdMh8iHfWd/d26KeAq2qWFU8OyuWHnldTgSX7o6
UUxU+Yl3+bDH0yagPIfwVXpDuhE4rUSi3uboM0SEcQHOANxgrQG1DlIlKBWk0zKN
DMmItN6f+rC7sSssX+GphaXdIRC5IvpDr+w8EWQoIabLrtxQ81CbDQaeQNRVB8l8
x7eknTqwMygbe3TpRmrfUhSbE71ZKasxFXFpyUUlIHOOmoiejbT8CW8diuojBdrq
bd/nXLaKpTpyZgDk0XptSbP2GPtSOi5MHvPJ8x2Aia3dUaE3GTGPNEPlTtVAbS71
TEAX3aMolVcLt58uUBEr9gGfQ/gtHbPxZNKF+EcKL+OTFzjCgrkm514Sfxfy0uK8
AMBnwZbsrfBPYXWFV6g5LZX3Gv2yhAmOVpCXwOacuEMyz40hdZ9k0A9rC1A9WNIm
fHL73hKloQ4d0+TpoEQgMs6bUfKzenh9x4BTm7quyKsOsa0gXeaNIYvotHD0aEAu
SDpq69euPNPzsY+j+wNP8wS/8acRIj4J2m0SYuw71JinJB4sDYF8j9HP3G98wstV
kHMgOA2BRckYIyS8cDOfJFuwISJxqfucAEqIC+w4J/6Xexwnc/SVxoNxX3tQiCmx
4PnwQfnJrULZ4yQuPHIfXLZS91hZeo5lKzPSoreHdPDg723mEchW2WUSQH/EVmkI
9pOV6iOaDO0R698J+P8IKb/MQXV0iIOQScf68frDCRh4eyn9YeAUerw0Ss/FHhqJ
NmajBEr6cAFHKPjhR3h3tRoWwwuybyCVNtCzhEzXFuAh6EvwvnatyZxLO+uqdor/
mZyJvDDA1IEv/NGiSa8pcYzG6c+ncXAgrUVgm204leX27sHWNYKTcKVTyhWYlWTw
+q6zpfd0TPeDNVY1M7xAxl1E5w7NxO76IicYv1TKAyiSXeDlsD8TjXCH3yhNYSFK
hu5ytQhXoYqn2ccPpsTtjrBfaXO7Umv0fXIHw2AGe8KI+UqHCSk50Y3JTuNYh8M3
mOJiBDd+JyjnVL7havOwjTP8Vh+wb8ZEWHM9pOcArsQ+zHhx5NuFgtMoyVrtNCFy
qndsunQnmb+oqRiguxp167SrTo9xLMEmM4dkbD0UPNygMYH7iuW0iodWKVGvErz6
pllJrDIhFPF5PknkPziF8n3bIZmKMdrrXAKCAXELiOVpZJFwbvbFTkL2H2QfJ+ui
lB2Bc22FukM7XK0Myhp1C/cGS2gU3DGjcCrsGdJenvWMW/U97ObW+5grc7yjs79B
b0h7zq+9ksgOO9J5ODmfoo6hSvwP/oPwwUzwg82akY2nUmANJHKJ1uDT4ggBBIYi
w0mESlGgocovx8liliuX/7aNcW7HCf8+abswyGVx+y7BolihsB79zt9Vs9SyXvef
VBts8JRCZ77S3f05393/x3Htmk5WyJmrK9uH+5YjvrCfBnGbTsUeakkDoA2LS/lN
VB/k2Cv7EEKh8nkKUOOMCkHZDU4BtsgGEUdUWE5B1fQK+Ty+2q1F9M3m6zhNmIxD
L7vmJOeUVGZnQaV2u2SK5fCPT5508jcrX8/TtxgR/dXrK9fKnwG8npA4dSFzmYH8
TRQs5eUO+ktBEXdlzWI7KOBTAmbeNg+tuffcITWJE7fTnktm4jA0wj1nvyxMG+aZ
BNgpQRBQ35GrrZSg1/YQLQyYeGFiEwzD17u9Kb7sLfAgtk8X1bPiNfutkQcU3mNG
GuiIFlgNNL4V1qXgxMqPrAp8KgaaIaOP6WAES0w32999jTbq1WfJMNuVgqDyJEXU
EYCJwq8MX/zWENj/+Y0SBtqY5NZOFBBI3hVHKo2yYeSeGEFF7rJavZ14KT0CFerm
aCttspKBt/LkBX3oK4/b9QFwA+EbDP5VXuzbIWOIMCT+fmrozOj+LvhKbI2GhSXy
AhBctD+19Fj6l3vuBf6mJ2KlRz0sDQhhLE4BTDnAx/sOJbhAie8/baRUaldHSR5Z
QBHOaupkfGx+VFDUdPJAHRmY574wTCzovaZZ+a1f66lznu/6mvkIbvYA0HTNDG6q
sE8/gr/YvEg2brpG6QerugyuZddg3km4S0jTCSVcwFhiEFRMdCmJKassfn5PV3Sm
R6dgbzwiPu80+81xScQ/WKHb68L2lq4SdajmIfxBqSnc0XLlLCwsm2MVeIwhIq+G
64S1vWfnT4Ur6qtATe/uRKypnVZiAr3WMmUCIGhYGg4xljJBZZ3xGMF14jVOKOmh
PlZeajwt7B3rItNRORVk/pVinJjmLTfz3k253n3DWKteQBGwbb8Lvb3sO6t1MdZi
YSFmEpgvK50MLtmnLZzTiQRlwsWPLgZOe7Mu9Z5LKmZCya2n8TdRRRcLl307G1qB
/hUiSgrc7jrGrZjKoJCeKmWZNtdpus3YP7K20BHHSruCZdKAjkZ1yLdfrHIyVox8
o+pXlGMnCjgStud1Xh6k04jn1URcdD2hmSZX7jnxuCIoHVXN2znkF0uMZoQO6l+Z
xkpUoaGOgEAxcVyhwp4uLczxNJiE92LSjWdPpAsz513PJEaQs0QSA98e1rxCLFTP
Jdmn+rBl+4KUX2Ot5IJJa7LklRSpC0/LQxOjJSklfC7Sk5j7OCimQdOIxEXUpyKR
+5B12xKg7lc4g8EnK5kQu4ikMpbCPhjHqg3xdXLW8TgU5J30qS2ydzFaT9f3Eumv
eRe3h/z5u5UKiUC/uqiYYqmopqg/AC5+kvWPtNCoTA9ykT/WS2t/7nGNjvO+CPlR
xr3G0hTOv10ds6CUoeeyTJ1LX/oGo4d8fZXwcqJmfcHQqB3eGl3Y0bnouNlUth6a
tKiwUuslzAOhmidXpG1reZdvmv1o36eMm0rzluR8CSroZbmf2oFhDLJaPk8/5j7w
17cyOB/mR1nRuvnDoKmzuRZvaPWHTZsSjYcXcH8S1LPaWls36Lv5pkijh+hRmxh8
Yu/wVLQEYD7N5tlpyG0iaPJb5oQd/7DBQqiXOFACqUUrTd5bM3qnSlZVLPMVRFf1
YkMSRVtrdH5A90iThaRtF6mTj3OiS630QBTJ5S36kEQYIEAQWtdCuWi/EiFZLON1
nW43WRtAZyvCpdBGQ4x02vJO2fJJZ+6NwF1y9lvMgjrrzS4mFxBMiKPNSJ1CB7W4
EGhyWCTH2esr7VcPakkNqxI2xOmudtVPemFWkUbOZpV0oOtjs4hAqdwy0o0KuTU/
pnryWw9ut+NYalKtWcQQSNif/3rqEhDuh6mQGsOMEgV4o1IQkFKCZwwoBJjWepEZ
lHBlUcX6q4u/g1fHwjH2TYHBDIVuInyzOx1dZOkSfYHv6Mtp+mR4S36ncCO0cnPa
NWbBB3rvqRrzUBvwmVzqaOVdTtfdrlXlgx6uWpQNPj559VTX8YFzQIK+SgxsNMNf
g4k4/6Nd/vWHU0cKlKY0DsPZhGfwx37z7uW5HqU7GHsHSgsLQDJ7KPjGzupIX61f
Du4jInJo3nOXMRxCyEGvYmAs1JdGEZSEiVcxOUmkZBkgj6FoputfHn4mYNV/t8kO
CYhhM94jHVwenPSBa8m2rNtSUn8f+aGH7BaV22uINpMQh6pIPP5SQ37Nqg+qRyt6
jXQBlg/JwD5qSBvJBu8JjllY+vLq84mYJIQSH3NJnoVZo+tevXrGXwptnLWLEi05
6lXJGgZkGa0VTHSeL3Rle/r7czf8Vk8YTFpncAcGg4eqe+93ed+IPTlKzH3h+8VI
77VchQvVTBgrvgT6yWT/xjK3bJsTgLOXaj+uRD3TcP74AP2gPiz4qOKyWmQEWv3p
0+IZz0zQN9Em0h7BvFzOjGHeY/xTktAdL95MTeUui8YHX8m0l3Vi0ye4UBUZ+9k1
PAX3x3WpI8deAM8VLNEP96u7dx8HejtlBzgOHabVI1cMM0AMJjP+Xt3KoQlFI1v6
KTxjRc4Jz2ZJXMm6mAjwlwDsNLikDl7FD8tukL8+1eKIcuBC9JJNo4hdph80ATsg
zf53FWt4OzmRhOkAyf0mVrPId+hOljAO8+izk+WX+ngp7slzT5VWR82yGhZdW8sv
RjQOIBKh+NUhg/VNRTqt96dR4HomNWM7Tzdu+D/0y867258DxCq5z+CvsbTSFsLm
yRN7dphg60IBkOeKYzEa2VRYR7NrLPbg1eblCq4U5ZWQrpdKQFKlR6Kzg5cdZEAo
W9XmbEr5nZtX8hWPTzWCOyLf0UzlhgtWKwyhTsDaFq6zFJCq8q3rgkAizULYqdDe
GtyEST8jRzVLHHi9MvXGzE407yrVvrOGyQ5NhHcM364MsZeGW4xMowZJ61X4DuI8
DfxxwaZifHg53WfghXMoPEHqGGH9AUn6HJp38X/Ox0jieQ5c30RAM4Q3wI5rziiq
FlYZuAnCnuK0r8WX1s7p0QOLm5ojZSKAtWQJrLXRcihCHz+heClQHoOJmfBKRVpI
Bk0xLg+ZgjhuljsOjdkK+4U9BnQ+Qng0M0UbtUocIcXeBXIK0CptYxj/dFCT40Id
6s0J7lKxLoEJma03Ackd4NVQiEr6NwlHBAVvWEwPY+5juSGybY2MWBTaPE5KX/YL
MA0V6PQUlLI1214TqWLwJ32Dz/k2N0ELpXJAzpBc27c/pBHg78vKRr+qGUVHDRf2
mWQ/C3mgTx+s2Fvd2/qFHsU5ZUTJhfkeW9h+boLA0uFyTf+ci9SMkLpRowO1YeOZ
n/9SHPaBFKtDO3A9kTbVBrN4NvAIw407V178aQDB9mVVdexNPx49s8HTiCaP2ihx
SJ4vG+RXzUXkcX/UyIsmNXl9UcXWcIPhtQNbxBK0IpL28Y2yQDmbi94whRQMCisC
tIYoQQ9sT73XW5m0Ws7dEs0k3Oj0Q2HNlp8rMvv4QLZAWcN/hPtV3UUAz2Iq2sfo
4ymMHhU6fwNpm6lCbfIpQgcjTMNsRdUKEMvKTdgUngSrLQFj5YKWxVNB1jmWB8MN
k+0EEoaYNV37rqfHX+47tqlXTzPXHhW7tmxQJ9eK/bYvAnHnpPEONbCcDUD62nkX
CpgACkP04+jYxc8U5szZ5gc2qbaM1SCuBY1zyXsuY1neqRVmzcFEwQ9n8Qbx2Wbj
H2y4g6C26ZUJEEEZr3tyhUhpWb+/7rjxx57IzDMeIh33hy/HmJqh3g9EIYts88U+
GeX2Ax1Zuq7hMpjqduuX1rnNyimPpiaUGs2uEjuJgl+3LePQ+RCij8xFgQezrmOY
jFu0IYaSkfj2bNiXgs4hxVBUssPT7WE9IAcIoCg6fGMopJ3XFD7A/1yW/uF8MT0F
rs6AVGt9cJSBFQRvVBctX3y4ROJuCGBAAmg4GYnbR5XeVyIYXyHVEDavAwYd1m8I
HVzXzpScIgKN+Goypr+WfLwIKfnNz0pkIcj7zH7KplFC2VGQiHBXjQYfQeMp0gWG
F3KEqOga3t0zf36hBrhhrxeFO5jt4eBKj3XWex35RcaEJknLwaPK4UKxdfdqopnB
2cBXUYxVI6G35szZNFHblK4fyFGReBriVXBzgLnmzKFL6zmSCQbzqcACr5OYiLoe
TTi9M2MU6VDls33xG6g6gPrsiVgXuBVQ/den17LnqssolXjsiEAdHgsv2LNQr+Hp
vD+maszunm777QQnbExDk3xEfKk9LfxThPvxuLRdlD52YnwoyKhMyBCFzMQDGqmN
xNVeyx4/BaA5Sd8NeK8kwQyTOdzGFTxPAx6vp1HYV0IlbTr+KGgR0YsgGQbnCzLc
06u0ZbmwXEEK6onJ5f6D55QxCIx8Of8wpR1vjR3eczRPWbMgAT78nqQTnHDfPCqf
H2+7GBt4I5GN/lrRbTlJP8r20IjtURPgFY1TvW5zU/h8Gt+Zcn2KD/lwY3RlzDy9
1OFaBdptXV7t94rJ26aX5zGP+tUbHlRxwudOTokexu7oK/WP7TrH+IJ8A4S3QxGQ
/UsmiaypEhG+W+4BI65hTNn21mMSViTzrPuqBlAPNw5KcyTjqOBuw3kcu/yBhUkk
KVrS2J5ZMKdPSma4ne9YaLF+fhGQl0cTGyPbkJfraZpLLNb3bDgnH6K751FRRUmF
uDA3XVpenLi1bJZg4dV6ydX6E14uZ13RzIc0e/mWUvpRbkiCMPyAS02g1WnKqRdv
o87D7eERTAFR9H+4tSvV4/homHhnl0t1ovvFo0mMoBibk+jzDTYkk18f2CxgjdQa
3EFTbOjit1eIOYr7PgU7WDGW635CYH37uHj5Qf9CYywUo9JbnQ7yZOlT8R2ss3/z
VqcdTTpm4VXWY4UyZoL6lyajB1TKaSvTLK16Zyc3cBr4UASfMq5i8UXc0HU7nAMN
qUP/t1qmvjJDuzyAPVNUYGy99+lQiDKaWwE4oHFCEAkGKounoE57smf7mjveGmmO
03GW/nhv1286jLQX316zrwN7U57k9chr00jSPFu3my44kyrtYstaDMfdJQhnoXpI
9CI78y3ZPXxMWr2HkhlYxvWwaEX8deQlwKC58NP9XPrdTTMTOrpcWr/gfarBmwzf
3BvGRcAP2O/EghWZxSgcKEx4zqWfP9Kg4OYwwW9Z64bwrje7CuzRO2a1D+KaKWTa
iBd8TfzTthi2AinUUSrFp3Y9wqMWuScDf3U8grSnXuxB0mnuQSVwJ0nvWYAKO4bz
uEfX7MYIwU5uJX6hIQ2KHItOWiIi3YpZa7DF8Aq0HRE6G0qv9gc5aTik/Q5D5oYt
c5IU2G5smPciGdFhJvgNnLDC7D3nybEb6xqKF8ckZgMsKFlBL35hKbdRiM0AwQV+
D0JdTDbWd5HyqrPYFCgRvxxL3pwRRkZDIISfu9uw6qT7MnQqIc8zBqGyhZD+Aqpc
AXqul9RtUmAPs4n83f/Tku2zlJWGqWsUHUEGF/SPiFa1s7nUp2DKqK62tux1wcJd
gBR6Ehf5Px9r49d36QfjU9Xy8mQ5Bkv7sWYKJPq+5wNSF2ahLX8sM40U4MWMqUJ+
gdAh7pgJGy+0gBCr3LmgSiGVa5F3nD+9WXD1wOyW6/raHHz71tzNMl+Zac1pEWbs
b2A0BHkXiuRzFq+9O+JVSBfBcm0odBCCoErJOfUrHfBBpP0jqOiGM6xa7P5Xm/jg
gFk81CRhWJPWz20KWieHWacGwZEBaFcaO3O1RmRTcoO2uyXd7h1543x+uBGAXCv2
WSd8BiDcYmNNWQ1eQ6ZZll2Q4FAYiDHBdKGNJpm16BPXkubYlFksXRKFZSJArqpY
kz9BNaHSE8NsrhnwTCSiCQ2kNzhyWd8AVOWubFrPQOMF2uWVLuuSmqOYTy/Ofn2p
rtskoHCeyFsIATCs8tc/DLCUy8xOshP0BivlBXad1XAAI8j8BBIjs62YAa9kRDbe
7GyG1lSdyyzyEG4KXkwdZw036lLnYj6zVxXBVFwxnpYD5NqvusOo+gKzsj+NgWYH
7z79+O0ZhC39wxLooQKpLGWE4apyTbJfWZGW+PW/ZlEEIcFPr59cn6nW5JKlmxqa
tlEvfq68iI9YpsMAyLq+/Opo6bRWxDSiEiYE6zNjCy3/hMkFQtAZGTvznc4DoZqH
72t1Hg2COD3mfsl2GE92CL47ig9ehjTOhgCH2Fmg7pTJXv4TSAIsvU/r1vGC2gbF
+YNd/i3lnNLm7EWGowON2GfbR6zc4xb7Pw2M1IFDZeWdPjvCs6BzTDl3XVMZwe5w
JftPjoqPgUjAXuUcgJeoSi5HU15OAOsiYDmQTSBUt38jPeLDf8lj4vkhq2IgEXeb
S2nlq3z9T1IksCXXDqIn8X6d1Ypld+VuTtTYl/5zhlwtCAI95ZbYfWJhmPNeZb4J
1GMLEDNRplmd0s71KQpxyFbpjWtPwX2WIGbJD/De0vyc+d1T3livLMXb9Xy5+mdh
JZ7C6Rk/tZmiX3aBEoaZ2e15Q8FsYMaFQIinFsolbwCepjSLlXVb4mtWz21H3mh3
ZLaZreEg7g1OHxfkscGN7wcXj/2xMI7PTirfSiaTa5d/FMOOvmESAljGVP8pHZXb
e31JPI9iaCLobGOx+m18XSCfUSSJ8hf6K+x6xVT4Kf62xHNnIurxgrVjrsrBuUsY
oE5fUV8pJpMgGu2G65hworpFNfbKM+f/0OvtFklwkBb9pIhuubrZQsnNpaSMR0ak
lcMFHQQ+pc9NzSWEOz1JJDglBucozFWomUqUOzoZ7T2pFILDN4hprg1Uz1D1SivX
bNKjMQ2MMXam1+5FklBqNM2B/GDoEGf/+zG+8r2CTdPgorc5PwdRG/QxRg+eWQg/
eMOcWWiwn7NuLsJKFyQIe+nyhIG8JCj1qajfYuAEXU3mc+x8yCELPMXmTj7X68Ck
9OnCFMoWo939BgZKM9T52eve9Rwt7++nFxnkjiid1YouJXURt1Vbcz0YHBdVeBba
3TJiij8LHH8qbVr/3CBl2THy5Ecr4KFUv2oeFhknW0r3iyZoNfX8mIoYcfx9fuQ0
j9zAnK60/CZxQTeUZbqP8QwDSjJruKeCO5AmSRF0SKQ1fo4c3WfYA+3jeZcYSCym
DwS9GhryjP59SdglcgjitxT5bXgLoa9n5am8BjtZNxN2hKIqicm5X9zi+fpu6TKK
2JX456fydmksMp3LaVvQRix6cHe0zSfcfYXqDhtEO/1aEHWBVDtq7xkiiGdCz1Mc
R5dZmO7ybfIAU9cKKnMnMhoeIew1QUkRtwvgrXEUw9+V86CmxN81ZrzcRiM75ADn
d0bJk7WzRCtEvsC352Ua57XWsmcf8FupsFvZNtVPO2IBKFwi1FqhPrOzVsFEtNL8
TGZAAL5atZdI9n5gOgjP/aM6UKzW7vaMpa76wdyqN4kLBWf5hsk29k1C3lOz7u5Z
FeFuaBqwesAU4SEGfZFJWF8Yhat4SLZlhApcH0VwWXsLlAQDZEdu40mYBo95KxG2
K7p0SjD+YVIXY9goYChCisXagQ4J1mCEtgODW4H9RKMb8CFcI1OSf+lfKjw+ouzZ
W/f1wg1dwndJNI5Qyki/yHHhmbLtIEs+j3bsidBtf6zycf0ddTsxvtpmYEQ8iV0f
ScRshqHWd5IXSvFcVLSZ2KVjMvYimIaHJ3DHHU3TnW1RzQfvkV1Fx+GUrk3/7Ze3
xqCBR78vM5y56z8LAsdeOvy5YeLJGCMSNAEgBii17pjqyDSzpRMoh9lMqanvy0Tw
gbgJSZrYbTL+wtg2vcjvB9LtMvoaOGY1WKOXfv0H2R+XVOTinIlPZMllcVTieBCJ
prxdGXo/YP+UdnheUNNcftuNRaTFT1eReIbBQB1o3KUEmR3Ds3nw4CVwAgX6Th0R
rpkns4ioyyGv2awyActEjlOrBhZviw4ZwujeEG6K+d5mMibcRZHFfGsqv4stlpyF
GpunjshxpgYfqoUstDqoV+HPZIKoFvBBCry9u1qT0SKtvtDHjSwRt+wOlg8bbOOW
RF9TKaMOeUjS+RHmXXJ3OwTRB1VDT53uczWpjON2gVVwp/5VXUa+ASaszg2UUont
HyOZAavwnH9nL3YiQLUmJupl9+B+PMMoOHhApJbQhleuVrTgSs8fdGBYWt+xxOdD
d5BLL5D2qDB0070xCycm69wzUVC0P6+K3KoGS5mOm/IrqMD9957PSDq7Bvixgy7v
J+b1Vx4Z9jtxD14LIaoLZliBz7sycxex68J7gUJTT2z9xJRyL2u21zCfzgXvdQzr
GheT2aIg/7pv/YYcVFnEW1fqi5F9UP5V43rEWz28Ay92MxsiDT2ZiZOiHwNqwWJs
j49koUOIiZmY383vsgMMYD23o96GsXYzgHQWfmSI6ztdSYH8hV02UzjYRBaFB7vE
9uwTLRFh0cx3/cmj8DAEilGRUuLMYzNsN/dMpRKmCs/g7ICkhsMhQO/1CEMTV6jC
KCzDqE4WgsFnYDsEvBPnxO8PZ0L3O8hUvP64xv4Ct4VtLo4upSXsDklgllCsicQ3
HqCYu0i/vyUAdhWYoPHADwXYVfXXK+rFw4iNP6KW6RKoE3LXmWQi2ycqeHO6Cw4/
WFYX1aVOG2No5NM3R3UAE85H1TA0vQQ4O6LPN1zcRqLPNyWuQ3vaxwiJoCiF6Pew
FatU/y7HlDOerLk4d7sRSvk4ElGj/gK0O+FKWJQ0B+lE/mwbFHlZdteDD/28bh+N
bzmod+Z7VxGBIDnllIxHKEbRZjbELx8tJKQgGOFDV3FlgFIiR70EqKDYxU7FgL4E
MHOxukoNGuhv5+l8rhBVG/kLJCU3lsEyLCe2ad6WOKRc5Q/L18WT2i2t6CCiHQH3
LpGViTp3IS8ToRs27gX5CGOydBrDcyhk6MFsLI9F5p/9/jweYcZzacwoPx1CK3iY
4WMg70gE9ngDaenU2EaQKsir1IshkFEzKHJb0mV9WEoRYCnRx9xGovmby8BG21/O
LcPxigtCRrNFlDkeRmLUR2H412wyu+TmP6tpb3DxYuEDnK1ONLfaSt2ewkDgiKbf
f8a41UpeyErMq555I/05ucjlux3RS7xoGNXyf4y4tFzONVgk0R+8ShSdh5b7GCN4
fF0fhLFiUUCzcwxYM3DZyxmjsAyON/rhXeOljhh/xUlN9sCHms7pflsTAngUsy9I
9m1ss3ltNct2kp12ll2mOvVVIVLsVNFKgQ7NhORQXkrfsGfU50bwTPYgz7kVJmmW
RhrYnq7vuBDBr2YDJquVl3viu/Qr1TpaclT2LtoiGjzXU/hyf7afsAlMAmydWZnj
lgeaNY0DSOwKIEpvxx+CPBB9SUZkCVvG683bMJj7tgM1skxJYOUTL2CojayrOLf4
AfivTuOHV/O4hgHB8IOSHS8c0NR6D7pDI9e0d4UNev54MRDWmzmjik1b3Hy3m9wF
JesvzMKfwZklE34/ccBqaZkI8HfmDbt4/BfYypBkzkkq2rAY+xjY9Zz7aONjl2OH
Iq6eFQv443lYz2Kqg7OZEzog0llqgG/A96dSpGKfvQxBHa6xaEBEbhygXKG4jnWy
0VZrQ2StwyzPWdZdKq2UtmXz8s+SUKtMgA0V8CisliOGk/cOj8IXBl/SwFhTo4Q6
a6vIveXDXVDoJ9cYjpRTFTkil64+z5fs4aGAXyEioUYwtzFB0pnuXKrtd/pYRayu
hJaDxbK3m7tLtUeA7hH6nLpvx58B2H8yzimBfP+F+nQESC4IapwM1ljPslKrFqLe
2nhDPTB11RgNilAue0cBeZT6Mvk1KGo/kRfhZKEi0H86a0yHKiLetbw+VYSWo8+G
2dayZOkzYP6XuERBqBCii4cHXKKAXzUKwngWU4L1Hh96W1cBFC/QuobX9eIwNFcy
dN/xEh5j5vmgxXsnvOJouhbKgyecXehbIxzRxSUc0wog0nyy+eE0uJIiVIzytlHp
Tr7bsbLLaQZSa9qRgYu8Mqw4PGyt7XjGqvkBbtE/1y7bCeAR6JpUI2Pwt/RSglZU
wEuJDb1MIAU6lXutv8WH9gNjp0SFRYinY41dAObB/n75/tJrf20ve4NHpzFMFxAX
JKEOrGA+AT+izWOKdrRo9Y7fi7iv/6WvE+Apq/AMWFlApEgWuACejVDNSrkvI4dy
02vqpfS8T5E3+cc3bkz+25iK1pq+KmiEyXmkSt55gPJDDNc3rUceLvjVhSR3tiJx
I/svtTYe9EeSq3bSYus7LYRRMYUWxLv41kfrfc+GNj4ZigZenjXaHx8yMMHpfRhW
dCvnFSqLBQpUWUZmYCrWrfNXipJoHN3ZjmIqsfeaGNF16iiGu9rjyteD7OZ6lQbr
gDUYXiqamxkkhsNJt9AdH+DkMu4BozrUPlYszfjBa4EhLBGKlRQOP+t4BlHhrzr4
OmH+BHHIjizwZNUeTsV/UpvRUUoYTTMD+qdLhdatpQS8tWafF8dQ6DqidxCnr9X1
QbZ02eDTmmOs4Lfi6xAkGrp7NPEWDzyaGVTkWiJLTx4cocJV672LQ3u8iBNYgrVx
TdLngc3YsIBi3vcQJKtHqaakTmSGMryfby7W+5lrpecBr7vS6X3SOiWQZ8QjVgb6
pBkylz2ujkw9say8KsKrMxDtVRyCf5McZGvbcUoS3O/AtJqILdBKCTKhpx2w3diE
x0gQn9Re19ATxPO9Ff9hMxWyxevjfUUPEBwIAe+xPZ5k75eT9umSMagbz0hhUMLJ
zA2Mw6xbbY6IGvTloumloz6HWdcT2RI5+7xvEjSYtsb6qXyGkv/xKTPAasKWOxzl
aYYciIwqHrfl0dbhFph7fBViHndiGd8i3Y5dKxueJ6Mh536PgcGpacTnN4isZhYD
T7HENDEdmgw6+q6X3oMO+FmVEQfctaagMGjMidhaJmpFMGGjtgxBX7DUfvuwhv0O
N1Bf5UryM3eU/PK33KvHN8+l9G6YE+goa2jQNM3G92s45l2vExZTbwdUlseGIVSh
GQeA33AZse9Rz38eDuZk4hm+YB5WVfmufZBaLfkHUsrvmjeAcUJi3HcqPkiZooW+
CIlNdIzKcOB/O4hPA7XYbBbKQ3jXsa6a4fukvnz9ud4cJzBkeX7X77jTn/2T0emf
jAFOmopy1mtEED7vj8L5elr1GRGZIbGc6cc+Ilbg4sSwqp09mRYalIMCCYI/sqcM
WV9IZxEndvI8D8E2huhqkWaLP1TVDt5kS+4xt8sGix/OelPwnMGZmugRIzSmCbrH
93HkFtK5RxUc3sD3o8HoarQru4U3AGDxMi9HWJoh5OaxIR7hmrJKIJa/sZ3c9+Ko
R+qv21khaD/awxNWhO/tbZJKSc8cPyEcTUufZWNuypezYcrtDZ4BfMY5CLFRdgyg
N0epmgNZ89sD8NdTWQ9hAtE/MyMA9EK3M1izR9Z5Tno9qOTPAtbkPDWxCJkK9Zk2
PdD5q0oraa8212H1DUOakhC+Nuc4FDMugoYiepiEt+v8kmP1FdAGBdTLB8qQdtRq
g2pQ8lOYZvEClkgOEmdMNnzpJuNWD+RwA8N4S7CW7Hp0sb7RkxEw1/JqKzxjBn/T
gn5oDtGgqPHcEi+Gd21hW/70pzoBPSVarpO/eWc7l4HKguTscwxnHJpAdt2Fxx8Y
v+2bIudyO00u9kdKxqvKmHaB6+MIT7yY3ZAbmQd+f2e2isofKmUNLgqjjdCl52tK
XbJO1eteK9zvWuhqprN5Xo5AFTDuLMsIvF0S5NF0zfgjbJWn9JRIVDR0bZNCY8tT
0Okrm0ZpdH4Sg400Nn15mNJ7HUSUUg3GLjuvUYHxpBr/hwMXw6wF9YHdRcA7JvMs
CjuSyAusMM1sxKZalQ45SiA1gh5e6WRqlUPYYWdKNb9pf2kO617D4hevqw4u9Opo
wHZpTYD1U6Uldn7kfV7oQhKwBOIESP/PnVdICC7w9G1HSumcKIqe5Wa8WKHRGDjJ
e9U9RHUjpw6LNvY9qhjiFd+eVt2FePIeh0YrSXM/5ZDco7pVcCanElpcvGTIKo9/
AFvJetIYOkxNsc9MoNnlU0PBP98yj9o+DJ4mtVO1/Ay9bB2QXyazu/EKtdJfKtY7
Bq/Crdu6uuwjz5Co+l9im4CBOsCxi1Lxt4cQinDQm8N6q5kF12uFJyHDNnJF39zA
wm8z0CwzVFC5gQzwe4JDx/sFFHdmpkA5K5McaRiNlg1kBPrN99ilq3ebtFvSQtcV
Mn6hHhfZob+vB6rKNf7jzB+rk2RNe9XXiLE8XFwVJduY4H1QV3PZ0r0+GvOwp3HS
0m4ZTK5DrC7eQKGGQiEgXB2Lrq9uGtFDUORDcF7TxbTMbOPYVvrYesct15RXHwiP
3UGLgp06WYYocL0jOmTY2PcIqkMDHbJcRtsJm2HS7bzhoCgkQiS0lt0QOCotqKzj
Wz1BXxDWD8Ssu6Lxg8fSedKKD7EDUHsIT2LoLOYHyqyPgJAQFKPDuUsZw449oNhc
TZ2P8/zPPMgBzu79JlLqiY25yAFB0jA3Nck0ApGzwp5jJU+ulAla1EiHUCkmXVdl
E+bm1hHn2DSol1ncWDJEQ9NgWy+maXAwDVcNTJ9PYBH5Dcg1UxPLSM1jOfak1Ghu
ERsM/2xG3JrW2fDM0+SAQwB73YWiJ9O5dff8FYHMuB0QfDgvqwEZQ2blj5HAR3N+
NLJW7NCvlupOb+S8R6zHMZ6cmgxAECDcPQoS2dBTHVR6duZMcbGQvajCGH1r4C4h
A2CFsT6jy3cjmSdTuG9ur/IooCTxV/lDPDUZkynAITBhRyYJZXUQKZ81RHheqjyF
I88JK3Z5y7aqehAjR1biz0OnfisI6W1y625Kaq6AM/lNiI9uutDLj51Q/pJ6gvxa
lgBL95OjxDvwBqWguV+rJ/xhiuij+h1NUZhPu/WK+q4xebNgT77qiI5vFkWebC1v
ha3WRgtb6cY2WqDE06klfDnx1ifRySjV8Ref7oPVZSUK/jGt5Q5tkSwIlwyt+Sa8
2bdGXFUfED6QFjIfwvNIgCZ+Rvn6mpezBesrjsIuxXQG3dG/PnIf8NQAUPXZTvbf
8s/lEawG+uXlHjoxbeNtizw6wxU8LOLCoa2vbGzNTF3Jk8DdZ8P6ky7FsqhXsHp5
bTQNv4wyDNbhZkhvRMPDZaG44US0rYfkvkIbG77Rnc+KGJuHHgEeipfGacfH2Xwb
drNj4RV4BxB4xtnapGkBMBATGRRUViWcXvXCoWthYLTygOGER7t3Fmwo5R5T0iHY
USRir02eci898j4SwasYEe5CnlCFrPvx0h0DtASW2Fjxc/+W97h1Bzd6qzHDVy/d
rWYHdHyYdyQvuupiacNlUy67aiO16LH8igzki1mLj+/wEW4wyZ0Qwbvtxc8ZTLBe
onKjxftKezKUZXR9HFBS0m86kU5LqqKHW6PDdlNH1bUrKlszWqPlAmG7oA3ob862
bC1ATj4BjSEs+PZq8wRQMouEAJsKaHBabF7iUWtBx4xAEi83WP/QN+BU2a7P2H1t
CLDQb4G1pU9QLyiH4ZhSHpGZC4CF9KmWWGObRr6vdSWa9x14HBdoK/1rkkW8MEpB
vv4iMHnq3gdgVZEqg/KLdbWcJBZRBak7Cve5avNLcUDdSc74wKoRriTGG2DDHeSx
Y+mCbbNojzfFVV1noS9ujruhe/Q9YMTvSfu2uBz9clDrRRQFDTXNeQ716WwHsETd
mtwqn9hCDnWDMupUPAHBd5fkTMoMJAp1jHoyKP9XzzfjXvtz+rfN3n5xMoXWjCuk
iJvYuGmYajUWVsvS9sDwIt3+z3WQEy3dcpeORBvkdKKqaSC2UMiETggB71AZ3XMK
HU75gcDc6qFB3hJRs3Sp9/7dOcTu91D1nBSc7Jw9za85WaX/Uqv6p3PViLG0PhNo
ydAh6uMlyW+eyKboDp7rSvXSdeyYj1gEBHaUiM5woTMTvGE6o9x48EdIWm6eCKml
d2pZy26zMrFQcpgIb6iHnaEs5s/zvI4nJxCjS0Y4BwGaOXc6jqeeTHiFxHjLQba6
ZFLKK0JhDVnuVFn1fGsZqHDKakTKC/2tUZv39sCu9/6n1WIYvXZD9FTDGze1SG8u
HUeFPHVl0BdELan4RETDSlj8cJ48n19cyQd5By5hSS9gT+tNo2BlP5cqiT0DdzJ3
+MWD+5xC5bIHmzDBOfCOPVZtdUpMAvQC2mXXdt54OQoMMtRFHUiNpZD7uZjRgFVj
bSYX0/+SOSamtP7rC+h/UXNLyZVu3bmlnRTIRhUN26s58NLy9cgwi6fPGNA9FH5K
DFKYv1YEneY6RiQC2tAjekclciuNFiBve3+FoqJyxMzxS/vnvvkCYwkny0nLk9Dw
EHlMQBgmdi+3fMMXb+Pdgb6fX69m41R6HvQhJJbuTfkbiJPGSgVfq21nuqkWu4bZ
pnIUcRDqt3VxpPbTPCi/ysQqQuzMhnaFWuQhIuHcpZ4F4qi5PVybY05EQRvDHBLF
5dsNOoLDYmY2WbBpnaL9f2ochAtfOPBWgg7ssZy0A59PlSZiU8/ezUwZ/LkUp1hR
PGYoDamMgWgOwdmstGSK2Mwdq0lIFgLCU6wJV7hPLT6bVrwgt39KajZf82jKpQ+T
dZKHuKrJJwU6iZDEPmsdCBzqlJt+WsxFybMfzMddYXM4UG35LatK71m9TMc93WyD
fNCCdXywZL42LktnjJWByHhdpR6ynML//l0tQxPIPvtdJnLADByLRD1M8ciqQaaD
TLy/r66MElYozPNzm+45aZ14QSNImKEauLAzeyOVP6emNHqe6GqojLuxPeYdJLCs
2UkzNE+bRSczjV+YPmEQmCj12/OTYo+x4d0aRcyxEFVzfaeDujGZzoy0t17Qwp2N
/5XBIuUBp3L6rZzGMH+zXLZj/ZLu6+bfucD6MCei05pEHvKpVDiZZqbNLlnpzfEe
/WhoJbInoA9GJlP2b8qHOf7ddhVubzk7IF1FwexO+eoNDmwrTfH6iXeWj1Ps/hEw
cH38EbcSRkRA2kAq7N6iZb3WHPh1wV42Nfl1f8rg8/ChXjL7r6WpotoakbzMaujr
Y6bfQaOJ1Qj2UuRU3D2e4mWY3MWdwsw6Tpd1qtaqNbd4Gb5bdG8PnOd+TJnSrj5D
qyv4wCOjRy/OlmgclY4YxXAfyDdezTlanBsbjWFoFF0NcXsRF2t4B4NcvV/CED/9
nisEn9M+KWl1EGAnoxA3VOLZH5W6Awg/Joz9fO0/xx7jYpUYw1uruMA5sp3QDKPk
+pww8spakxsdAMwgz0jspY6AaL45gYcsNuRDyk/IgGsKGlD9bqLQY3MDOdl87iG1
4MQCP1+u5BUPQmzE55hNsduev5j/xp4SjL5mjT1si/xC91ZpcW9n8vptwONyfGI5
vu18sd4AwAPrkF8m5CvaZkWuwR1LgfbWJsmwbbLwpm81V7PVKTSRfzCiaUS+6VRH
VPnRgxCq13I02FJtjZwnjyfULljUpL4KMKHrbvHMKtH9h1RZGaRCkAaBPidJImIB
Z19fPHMdxPwjDfrX6E3B5RIQvbbGU6Vv1Js4RU3toYsUFcRlH4KTbjU6U0zEz+jB
uvagIqL5PgxCbOHsCRVcqui4n3RLngEXdF18QkDeln/+8aUWvb5g/Xd/lWbEEnTK
aEXkCF5a0WKmeXGBEH8TGnNmlylAZeM3qvLQTHlUrwG55y7XbKCzg7pBEEx4wyQf
gXwLYvet7yGlnS68YYqB863ntS3cwUCS1orrjJdKnV+cfhaiJz7tnBHcr8gB5ke2
NRdss8Q8wza2pd7UYXCVV1l+gP7H2uDKabGsfsnvhI8FRejwC+LSRlmfe3ggJxRG
TegwLJ7XSwnkJt7Yj/CeV/FiUGCwq1+qLNOcS7ixpbeGTNzSDKYLeiZm7+jMHWvu
l8+CNp7H/f7I4BV/pQoft861GVDkIkIAgc7vJXJgcQpMhNoo7fwc8dOw3CZHdmBq
Ro7IGbJerfG13q0JuXkeC8hbDI56KaGaD+fTzc9QmgnB/z0ZO4z5BoEis1Gb77DA
tylbXwEg97YM0OgD0MJ1e81hCi95hA+zJV1Gr1ICbpw/KU7mLkCenkySvhTHnEMO
k+G+eXW/WTcYg3qMT3UtDSj4ljkpxDElGwgvkwFltoDQDGSaUtDOJsE5A4j+QswR
okhi7pBurUMmLj8lpQqzPAdXIINh459gkkVyTPKa4K2OKRLlsmk0bnP0mkbE2Iut
fKMs7jGhw/ZLoV13tVu3mNjQZ0+JKjNxSxfQjRxYqrwHEjhoaOzfpw4IJFuqB8m9
RRa2l1my+e0r9w+NiBqBkG1GjnkSmu7B4yKRFFRaeB4ndqzzQiVssdEjf0d4XPxJ
manOpq+CvLKuaqDglZGZlrOnDiPGm01U5N6VwyGyZwnxD2Zm0X3Z8A1L7IVqS8FE
QqOxrZKN+XDeiQjPwkcid9mXpqJL8gUNxMiDq0FzmSVRtV6ux35vnfpU4owpW6u1
Q5C6a0OJS7s7Y8/927dUHgBJsZsygUwHYQCxoJdF3lYc2RoIGe0yt53WW8UCuXiu
yImQHHqY0VNx2c6nsmHPZ/h4YhgTnGAn6TJE19s1XW37u017xFn77EPCu6v4OeSV
ABLhY3WtkPRG1QDYboLj4x04mt0RH9lV4M2uL0YLH3SlJt1j+NlKWfYSqQmCRovt
QMSQKSz7OD9f64dtuFaePrubj6fo58MjMO72L3CAjCITMubc18SaSp22C936H1iX
I/+aapaNZZoRPRoHWqsaLaihkfHLp1mIoQllGCULFkAHFYLUHsyg0BGVNk2xzeOF
xIDOPvmRq61xz6BDHYZgyY0gs0pjOQUN/Zn+Ge3dBL8/5a5usil3/0hmKw+ltUjc
VUDtwlN/Oq4jC1Gmjro3YkOAZ4x2jDyEZHkraKRe5eekLRda5nLvQdJAwlT0Ho3Z
JCzprq5fbB2ABXJNhgWJ4g+lg+viVwFosHUtB7Jlp57JYK//iJOaNk3zRA6YspM7
t/qX+pEPLOhSej3wk0b4+iKUEeje2+o21R5r/XiJRzUYDW8IS4bRPmjTUBwvn2R5
S+52K30xolZzEHOKIIeftAqpcH4FSN7jCdSLr3/34e5WBzlqWsqWMsmGz9/2giIM
ORHAEb/eeZ/JznoLWc/S345aZIMT11icmYa5lFl5r+wdIGOovgTG7HfPL7c2xXpd
OCopAIkLvkfdRgBLlEIk1hO8rNPv/JdcDKnDFSKUEmLhKDN9Ptv75XGtnl4H0J3q
Urfbaysxt3oJUQSuM3VkOgDt9pz8QRFvvwmTncVh5iHDTe21Z8cWELAha7vGw7NY
NVjk5/mcpbBegVrNrbMHI6A+vf8R6efekS/GBXihuQg8+e2NUEEbnWkIu5v7HDY4
/3hHkVZD0zM4jngSBgz92TKzZHBA2blQ577pGbK9Pm6zMcDT+S3A6q0wVDxg64Bu
kMp1q1LmLq+kqOk7uQZvQSa9w1vvV9QwGKBjXcSy6c203/dol1isTdtWj/Efo1Iw
2GGB0zsbFJLAmmaws4dfcN0POz/QELD2wQTjn7Ku/CJek0U1z0H/fIitYiBq5P5a
uMbe//Z6Jrwgwop7Xe9MDWXYPTTgFr2E+v8CHJ3c3+VlTOS7crwRjZJyBhgtoNfu
S7BRlsPTnLULos6xfQjJ53QxtqrVLKwX7U8BTcadAyaDqFYzEqfPFfqpp6eWxsVE
ZEu/TcsWb/elMHCCB87gFQUbpwS1xelB04sRG+PjeM0np1z+EPvjz9Lop8dB1Z7x
0Bv2K44BJymIy5iHajSuxgmutx6zN6WrGMNuRLNY3BVST3SOGVVb7ivWEGsOkle+
AiC6KCa3RAFGud8KtRiV7Q8Z6JjwG29KP4YvrjMdDQVZjlXxs+P7y2Qtkj7DuEDM
vJGuVenSTWKAsVCdfUn5UHRXLmonbJeuInsdiuPVu8xMdRxnXyJUi+wfy1IiLbNx
z0TnY11vC67jC9FanjBPJnL4VZpeZl/MuTEXuXjs5HgmC5ajIEhvEbd6CD5n25Aw
vxgxO98W90JFHH1iBrKusMbzn5NOncnoEYbtbKPuzGWoGUoTC/E7TU/iU6K7kBS9
zXHOvLg8IJpQfjrS4CNMIoCOwnG9LP85O818n62Dd3ahrHPkJUT5BzkCrhr/4kRU
ZHj1lFIF5Im9NpR1hkzVbE85NwPkt74n4h5077P5g6qTHfT84G6x8do1lCQNhY4b
AeKUs04jVOTPKoIw+Lfm7WruiOxP92AgtKJ1DKY/I36hERXI8Dmy3khENkGChmhs
LvrGe1HuDKdjKMU7lIAybNxeXzP6bT8nw+DB1WJAYg71aJNPYhDEAfh+JLHxyBrD
Bxih6k4iQVgLVMrT8EpqncIaT6GShIZwZSaJZOuTFtuXsiSfvizBZ3eyw4SMwYbS
H5OcUCoR/2vy4EitjWLC/EE/gkte/Qle9xMaJmNhkG3zTztfNklCGsKzuEmPdjZB
f7/L1ZyV/GWlzd8NTSJFIeB0ReSCNHkN48TUSND8V7+L0Fr9Eyj78DdaVnDp/+yd
GCTjVHluDg3z/FHo6XK+WfTPSe6qGUaJR1QVlX2FdX70jNmF5dT0QeM3+R9KgSOt
T2M7E+sCn8ON+S3JemwGLPy2n7S8QoQh/cjrTdJb0mKqg4WU6aNW9XeGUp419f4a
wLd7u++Ys4/eZ3z3095asFvfXdycSRmSLSUtKgam3mpx22Ak+uBQWEwQUExb4wdE
p/L5aOBzTqab+F8Om7IcUNir9Inh3oFOYir0UWPMuKHj9lodqJGjho/S6R4mjPQl
7m3WWrKMBEUqdPvgQ8RXe3+7gKsDTTGTV7U5C7w464YpyX5rGCx27rV8ihIaQaqO
VcX6ShPiDuxtxOa+fPfp/9HRZzD+j9N3KEgtujzy5RMLL+JHmHgpV6zymnnA8oOU
wCB7xpLiOSn0X5JnQ1JqPf4k+FLqTmjf3Mv+WMdIKahfiJYX4AzIYw8ju0wBzRCF
iCPx1zSvTtQV1jCtbZKR3Kfq7HeZCynfEXIQ7/1louQKQwTaipsIbJmWktF+vZr6
axRAm4YYVGLcnpj2wIhnWyvXhIFaKBWTltB+W7+Rw1JincdMWG5Xo+oTvLdRvXor
gSNTyCx78My5u7A/0NtWZTZyWkx1R52j1vpkBPd3kUCOOHW9liSV/+RKQtbCZuuK
UDVN8WR/6zxhg0U2E7uhHjhaovXj35xuM7eHR1ECXC3Cydb+rq80l4K5iqw94wDJ
mclWqMSqXgHQpL4krQwZu4lsQZl+ccgJ+VRNIuI/WW8QOnkxZeITr5EwBTkQz4G4
WEuM78H5w9fJ0FuxmGeXe3i3D7LizgcO10vQLzU7oeIrnKdR88eVZ5J1n8rAeDOz
j2l4u8k5aR3U12j//NuyxBIQiCvmtilp1OIO0gNKLKTyI4GotVqv5UXPSuttOmdA
7Qz4g7Pn2SF3h7BS2pWBlv4PoMtQXsqfWC21L+BY/3gHDLTR39+xIIE7kR9t86vV
uv1Q6upHHpWy0sZhFlGswDIpb77XyKYQcQR/OfZ8fg2ODen6J2Lw2u1fnhhNuwkh
lWImIB2BWIGPgsVl5nMnfJT8dHt624E7EZ2ueKU1JVoGkLogKycQZCbsmORz7YFA
S7uGmB8MrWGlzlEhjLKubds9locllaExATw5WLbohEw5hdNBqH3oFk0UT8OBTlZF
sl3v6xRzNorMr/oxFoTaQRRPo+8EPMaWYEEVVgjVUSmpWc+CZBc2PRD9dwYfDT7m
f1R9DkYW4d4QImOXX+Qi9/cJfRKVscmNHDFgLYmBRU1r4ZuY2SNyFQKcNLyAbqFd
CJB6rg0wqFQMvO7hIdO+OHVM9RfnOrMMTncyAxA+ZUZmFUQPrs0q0tIFoq2E2L4+
u0C8qjz7hKtCt8AL0cHk3FwqWRxWbCbvsu2rxuudXsYU5gId/YQOo7DPmnmPerwn
Lp9gIkpUJ11sE4N2yAgina+KO+4HyLMHJy9nPTaQ1/NyItskHo09nV2bHAUNJAD3
qb+TbZn0szqg3pPorhvaHl3K5pdvv2CgHFZoF75JKZdrXlOXnwggsajoPV+04cd4
OKEMwPWH59ztGtU27VpiQ3tWQpog9xN6wEY4dDSCz4okAj9JELUKLQVV2CSfPe6x
hGCUOlL61efMnx4+C0AgustIWdLPU3EtKvVROp/zy0lIe9TEc/RzUMBd8Gayq0oq
L/tWUyVMb+ZnWPJjt9GesjdZVdvLcL9OO7UXU5XbgzL/jEdiX8Hg3VQE1ozKF9PT
gP3q55CS+6+z17C+8bVqWWonDvkb/H2AbjKSREAUaAs1PTmmeY7+CzSzo8vZU5dQ
iYsqRTxZA62yisTdvkyyIEvj1QKzS65hfeC1Pu+KzJLmx2zStB/eaZtk5Oq2nwzJ
tKXUl3GsI+VN3oFydrYT+kv78OiquiiutzS+E3LIx7Zpe1asqrvaRgP6ZR0F4PV9
mdMiefan+L5qBOkAMPoB5ofv8DLM0q+V/RNYVMIT/KXJhlBF9W2HxUIhmu1IywFv
gTh3RVdv20xc7/TM3ySgIOMYZHEOStC411VfCIFLDEiTeMtiSe7MBEt1+1VHemBd
y1RFPvceFtHQmYkG+rA+1/p6unwWpoikHeHP+S8rIWbrvNGC4vrDTiIh8wMAwK/A
N4gKG5uQ0w+D5Xph8MBiwhWAd74idqX9PntNdl0MYoiZDXc+u3Iyy5Dhp18Sl3RI
QtRxAzWAC+hubjhGe1PX7TrT9597gkFPqISuZyGdpVfOHTUaa0s6IgDTjSL2G1MH
GrucOGd+40HjXGTo7heV8YxANjC0kf5oE0Zz5B7iUgsfdweUhkPUSsbd/EvbxX7V
rUw34Zqe29cDS/HgKYA5Y/VQ398c4dzanDuyPmxCA4oewsUQd1RSHtzVr/WED8t/
EaCckpOiIK6kVEOTaYs80iLtIhzfzehfS/Xknpig3erEWwrEkGlEwqfclUl42ey6
+whf98qfj52aCJehi5N//zevkJjus5GMhy/dDmk2ugvnXohhd+vFuYQSlNJum5dg
4x2QZ6ORLnkPfY6upTlMMqZPgGOhCHPZ9evcbBtSCmgSRrZRSHABWYciOV3RJzx3
LlYeyp5Nlw5k691eRvonlXBcKWdFS/6kT6eUuSZTeK5v5jE7JEqD+u4HJfi/LXQl
KHvPT2+Ps6mHUYc1M+84smDdilID5qi09Y/JeAELAhaJYr7ZcVm8lB95J/JQQCci
j+QZB0m4Hk7oFCJT5t2JNd7WMK55zOcVbuFgOsshOXU+gqbE41qDF5MJ8VMwSwUX
77aCPa29HCJNsR89hUHsvEwoRO6tSMNGa6Vjk3Cn25vLhL4oq8ghzcqVSnlZ2Jy4
k2RKGGLXFnnhyxxBAcf8Di+VXYAANpXIvPWkHFq81APx/4sRRRs4uUQYBL3j5Cre
LuorNbR/0/chcWol7+84rL4OQuIozB1bKo10J7yzoZmE5HTkRyjZlqvcKpYRm72o
ODgaCAAtqcjJ5t+4O8OSJPid8hL6dE7oWP0IYizSnNcyLoiVJIcOPnVQ3Ga0UtSo
dBqFZdW1LB6HF1Q5vXudFwmNPIl3c1C7oboxPLfsTzFNWcdvY91+B/9eXKBVUs5G
8zqa9CBYh4kNpW1AfZrfgel7fRzFNTXv5i78LUig9EJdDls0X9MTAwAElvIjqEj5
vCzB/fjARJBRhU3GqvrRfwwfqoy2I/ezjL8Bk3v6Np3x0X5jgyCiG/8O9FmXSK9j
3/oCTQVtU3EhZ8IuNz99QU1N+vea+xXKGv3y7Q6T7n4KQ+q3cQYXcNdKV/PqjBV0
eonW45MWoOAd6KaPcRWB4OOy35w3+MFCOv1YJyq1RvSwjRFKr6UyQNHj501G9LhK
1BAPUBOTp/zsPmc9+3ImAKMaMPLGmdWTzZ1uwRDPDhlt/f+Og1Xy/DdzAYmwsmaI
dbVAJwhE2AuVbBXu0i+pTflu6K+xYwoK8QMKNvAdF5tYwk+BCcQGUTdHILBYdeaZ
a0IFddakBAlv7QDhcgluq5v8f31fwz7nqkHNDpuEy00mDvVrpDpdJgJCyRpS5P/7
kFgdP4NTGAH8KI/PGnGHQbjnkEyl9oKDC5wBCBA/fqIwKT2UW+7mM4FEfxgPw3id
cDmSlbASQrAUuVBNbOhvVkumRvl6PVM4swZAj1+eD9N1qa5++24v5S1gydoLClTB
+310iqSZfyDDG8qtTtngXWYtEbytMmvveDDIlj6zEYKgrcVW99e/afWSJfh59dng
MroqBmq1UmwdljwnQM9PL91hssmK7E5CFLmCOlWgEW+KjFnqXadwGgOWflhxEA/j
G49W8k5KS8adPvQ6VSrNxRvcqd804Zl16ae4LSAX/nAzTV/IHlxWpR3Av6Jm95cH
DiIxLg4/n1HfgVg2N2CUUWdTTggt/w8fflKGBNTiOeddyLAbVLY7IhJZBovC4voL
G/ywKWiHBLBmfEQmQHjGt7jldVrut3fNBrpy2QlQypmtaeYXQ0DlZgO9JCemUMCT
Ixx2s/Cp5LfmUUfPTShsk7tZpHUa2UXu9Szx4tX8XjPAhKtNxPaoDKPnwvOP2hD/
U/PM2EHN/Li+OMyELsD8P11o00NgvlQndrJaeWYhZ81WA3GIvMhitGo2uNU9uKTD
4nYk5Iop11ZHUbQuR7i/mDKdlDdzB2M/cO9kDyFQHPz/+OjctWkNLC2ELqgpre7+
borNqclsYRYFInG59Hz4skFJ9qJ+1Z81ZDOnA7u9mKea7PRrYdOdbmPOen6WVjeP
9GgsKv28VJXGGgVU6z3IZdaPWQVevywI9MZ3hnswJb+qY90x/lf6kzJvFkkE8b1I
Lnkrf4Q5YZyxrNwHDF5mriS3qdXQAal59aXImpbe09kZTgIS16ZSE7doz0OEH708
7TEgYvZP3YtSTK58BuCkrWxUEAMggtKbHXl6HD/WY1PXVGFOyvqaVgHHFVwyLU9L
4S8hmOPpkR6dqpqPZN+YMxPtSK0E6CSp8ikB0wul11xQjzBStbyvFROD5zJ2Tens
EdUzYzI4SdJZgXf0Z+j0AaZPUZb8FsR4N7GBYaBE3mtQqi33egAMRDwmdJyXb79g
03cu2SYvuSggcU13fAX8iW90FH751jBYqynczeqz9BXE8tDkVctsl3AspeuvZzOQ
931gU93unDTpMQ/j9CR6XaaLRtmvVGXaettqWbr8UIxbFWCRqT73xcLUcV74/vLF
FigAsUoyrfMd662BNwsQislXYwrBhAXE7FwNR2b1mCMtPfYxTL4BNL5zEjZd/kTI
Bh2LAlQiDqWdw9TOLqNsM9w/4ME8GCc00a5P1rBgQP1ksDo5vq4T/rSQ4sZSAoGF
DKCYV8F9ovRZ5TZzY/SdMemajhw66Zch8fiCRjbHyJgDGyIBGdFUfAbnirG139a+
6QZR1Lgq0jribQpzngTZRDStDK4m2TbBaQra1jhrdVdpBr2n5WdqNgxoL6uoepfh
Gb0XQuCczAISMgqeKDVoZiCBIxDqwcolgtpTlJi//vro1eyfUMLJi+qu8beCLEL4
17iWiMfWfPjAcctP33kwXq9jQ8gNPBgRYjCOOsH5zkfPI0E4vx9K8ktTZzg9dHdE
PJKx99rLxH3IgWMRr5zdp1BosUwQ3Mupg2LXA2jH3UK8hHiq9J5zh8zFFl+A+6+t
zpaENp1fouw5oWoYmLvEV7484h8epntZJ9QY9hfZaToIRowYhlMBWoF+HyeBciVI
UsPO8WEiEXQNvlLWdxWJN7N5TBrMVJWlLL/a/1LWvnhkAxW7DqvzG7J4z+L6zMSZ
zugdB3KyHpUgMZSieqGQJxBZxRT0gbrETs6c8xyyimoMO3oDggtSDaC+NPC9R7k1
5mkKb1c2LzjpUDJiO2Ezkay++Cuh2xBQr4ccl5ZQJe4Syb8hSJiXFF7XIkhiONbY
aNF3RPN6sTo9d7QhvR4I+iLxWUrN6QAtyzXfwOyQ7N4xUopE+SLYpiHpTLzSGrkg
g7+47bmL3BWsENInqeJl6McAmRgMkCI3rfteILxnKaUYjuqfIMdpj+TOV6/5sN9i
qWSsiAc1Ng0QI70E8tBtcTKG7rGMNxWB+CbZfLc4vyHcsHITsS91f/e5cp5irFsZ
hj+9f659mLzbdoMC3w0yNFI2kCh2Y5YbAJWDTQpclRH6XthEDc2XIC6RGjlVkgVQ
wwPhNCeEIl9xj/cxF/vDZTWiojTK67LeY9MT4PrTZlCrF7jmsZFDOwz4Vjq7bhDJ
ilQZYOScrk6mdeFH0xaO8YfWTRohVWNXTBAyOxIjWr4ZgV+hQwv5exaMJRmjjVte
BIbqSVKkXjg1vdAbQFBJwcMkyd+ThtBQrwTf7xUp5ZrIMUJQfr1Q3ovxN0Z/tGnu
pl1nMOQ+AEIdk5WihxqhM6Xu+bpNrWiWrm3AwL4N0WIKEJZmv3XppEVfAfwK/C0A
YvJcK/Ie/eiT8yrD36WeSqqdOK1ibLmSxt5MhMSGyPD3qzUAMw9by9lBo1rrkHQv
Pwx22/h3nMSCCRCXv1nm3kCVNc3Qtch51FsQGDwSfAhHl0ZIcsJN806ue+zGyD53
OGouQqq3juLPANuYM24131wyU6OdSK69UKJEdHh4vN0y/Ik2Pe/Ze1lO+lBjnJ2t
OUnIJ54oKeGSRThW1QkkPXRZwWl9Keht7bgB/L0Qc3REKBZfUE1ErTKyNZ5+k8yA
HFZCWYQEhstfnuZNqtoD+Iw35i9mhlxIKqrbhjSuAgB/8twOmID2u4MdsdZex/Wb
b8VO7ObhoStaa3aZx0KlS5Zhnd1GIYH1QkeqaUmJ8uy+V4KgykoWhBTzYMhJzZJD
Dw1NbzYScblWKgTqfFfAOKdDz4hwjGe9K1IFYHrbAFNTdpSPrqXogFQhI2gcU0hk
+Kfxmet+ChjWsIcRhS+rhCdf43nbBOLKcg72xRHnZ53fbTJ1Bc6G1RMNtF1COpq3
+2Ph4ZKh+j3/P46V3tHIsKg40OUUce8re56tkkVZAsBLOr94iY2uKqv1SePNB959
EGA4wMlcvxYoggePwXkz12aFrkeyCj7jYsfwPGXVeDlWpVX9GA9HfU4PrD9s6psM
sigQsafEkZReJ7oJlvqmUSHauGVhMT2DCrmwyJ9pk8sZ5bm/yi/qL4arKk/KyCOY
B6i1nFtwkeu6qUYAhRFoevVB8ai7KZy9txBMwo5xCKwZb10pifzkKQccoVEXQ2yI
c6UHMcSg1oFXWBPb4qR1/YL8Xi96MmLOrzdtKyh51HI10HTIY+1KopL3mCFnTHrS
WHqw6PBi2oo3lCDAAEJvb6XofLJcC9UTHvQPoFoILsNeR7Lm4LKiZm+LSt650Va/
4cxiQzgICrUzmYq0aA9aschygFsVnu2lZb6gvcmNJNCynxdZhp0Ka0A1RHJb42WJ
WDt4rO69SDKaIZYocBfgu+xXJ0FZUYMLFyg2HOGTb1TZIo/xQ4uZu6cx+VRViXBT
tOLTrJNHY0feRlJd+e9LzRDfDvUAOnydCoJ7g996eniwQ0RhfWTABqTZL8fvKTjM
UMVp6iWPbKh/IFX/6IiU33VLI5H2RiF/8tkka2BYlcndZeSRCThFnCq1H7rQgJdE
qr63w1UgYa/YRCOjCmuVM7v1qMhSwWzigx0rddkMqw9137qSPZRFf7e7T3hrCphR
Hr7dIv63okgojGFOECCtrGlxOk7tU0H6JWl6ZNN+Ozys350EGh85QMRWPCiqa1iP
D03qa6vFQ/vPS930zr5IoCYSiy2vXSXE8HGZHQo4GcUfptvpc7zmTRHSf5pr7+OS
pancYcSuyeKAJh8eGr+DDCWm3gzYl2FZsVYmZaI3xwxPBe3ZvjgN7G0FkUy1PGTH
h3wCt6wYp5zqk/JZ3hfcMram3EkQl6jiQEydlvvRuGlRsEhYBsyKLG7cqIqfmiFF
kMz29zz7MDXM3DxuJWGrSrS+NvXRDGkCeDoe6OxVdaUvjQ9eoC1k7GlkoF9T6ie4
gAnRHqluHV2rIfXs05nOJI3D7oL7zHID/Or/v6kHBFX70SdN/YHP2xCG9Nr32gSb
AgrPRjbgS9KHv5UE4HX1CQMWM5oeZNIq4wvLjuvNP49ArQVVFre1LF2Q1scc53HV
aAyhNktYYbB++cYGq79zaTnuVeEEPOeX1IPNZSYtMa3Qgo/nZ5v//kzsRntd9ltv
+rJSGc0iedr4VRRwHNFYP3rJQqlUhIKNk3+jflFtZW3N6eTiM5KOkVP4RC7AEuTt
8+WDDami6rtG1JL7MFo7+n2nHFF0o+u6koFq1FVI3SmZt1wf2AjH8HAjrWR1Sa66
wlY2wqqeLygAHGpGjGx6s3NzuZzReqqUpDrZ4iMvd95qS1MY8Tt+H2SHKVDliDoq
PU7I/tXyE16PcVU6kBjps+AJMSeViniaWFLvLqk3P3xrdg7HHOF5KgrVWJ9ZvQMG
09BEDoFBkAM2dutm9PY5xpWM38tS9gUjZn9Q1fAEo2PZsbuQPcNR/u7rNNcL/Bly
dzpLvjnZ5vMU+pRN8FOb+XMdtGsWqE39SwhyZ0hZrVtsoJeb4Kb00Lg857edcWAd
BbAnKBkLpnmvgJU6MV1BsgNXiEaZkjrfSqpwo1hjQ9iZ7D6iWrIY7k/ud1Lz2KBv
RtZSecTbJ8XP+aYsAGa57Lm4DTg6m024TKPHghv32QYPntMmjtSbSSyqx8fkclVp
00ciURILgmuNVeUB+WoXXMM8xRP+ZlsBbEmccFmv++2ZKDqzgvGi5T+AK8yChxeq
R3B1TLeOz3/U6tIQJrIfjlzklgYGPvFqMt62w/sx6mYMJw67yhYhZAfimWBEvwac
6xEQ3biQEjubFMNlVve25EvA0kYZNkIWl9OLMTukkmW67QG9MUPf3luhRBDVbuAI
Q26s2ZxGr2lrPnje9wokiDlEeZZbPr62ucG9P5ISCz4GZw2SgCx6mV2dnLu8U4k0
OYtZlK9T6EDsUNTmJH0JHvZ+6rlQwgFZPN3SIsNotIUqh1N9ESbGoWk7HLf5tYH6
aLkr702TmczaT5rqyzbdJEW1T6GMWo7lJU4TK8e6F89R0e0e4wn/OgG+VhHEdGxF
1qtxjRhgwT8xHWTbl5aPrje3N5DX/3un9vGIa1FFRVbMClr7Iflcti6/4tuAU+nn
BEkSMzvQEF07wYqaiNSUJMpCjt1d67STkqFMUxFnhYC0AafX+CtUtQ0dvfTiXrQ+
gxHwJL2y6UiyybtEFgn57fZBKPlRCBdYzC7c7K5PtpqyPKR5EIDpDNEJxWz/U6Yk
KTuXXzoAkexZ76t7txX719/VapNIYF37c88J4gDjg9reTlvEWxb/RMVunogZ+Cuo
I6igFilBlpF2aiektfSWLb6RnwSI4PBBy5PNVqd1JpavNkyZkXoyOR+x0khyub+w
TO1Ggh/sHEZ97VLDw5yPiEZxwsTYYVWUvgMpBvaY4TxdSFMkAOOhKu10bJ25euc2
x4hu5zdQtoWLucfWn99tp8b0qRCLJkevMq/FVGNzdbZUqzVGa6gOxt6f+qWZLtVw
lrnQMoGWqnwEZ3b7PqnQs8maxJN33vz7YQxrWA2EEInsm+ahmSWMv6bPYkR2MMsZ
D9aJOc0+tHmCK/6V2mDJp9HJtrvZFW7r8BGko3UBms1S7gZNQipsWbf0WAZRftYg
s5Qah9eEwnoiIsx9kXJSN3S8ubIgUEDCi8Dv/84oWE4I8aAk8mHgwHSdCV59HQE4
KcWhrFe+alSc/xiyr203FUEl5KLOitjt14WicYs5ABLGi1eOt8qh/V9JeDwcEqwv
UerwHIXEH1brwyOmTEbj7k2c5CPTnatcpKziOW2t4W9NRCU95dP6/8KbA9FwCIHT
/4jWkGJFkfO1Boqw1hUEcFAjrxsiagbk5GuQD08uBByRuAvVkL+rsr+6oU+6eTRK
q5m3R152xtGC0M1yYCYaapNhdXJfSyttSgDFX/6R0zqXIi2PUovQdlzseiGdoKIB
jp+C37Y7paG//QRcaRvJY3+Bq5RvHlN6c1fLdFyTt8r3wI0GEzolEyApVVlJyk6d
i9pYbY7ys6bwCFlfE8nd+MF4xr1Y0A5VmqeopyQGjDssViUAA5c6z9Jm2Ro6XjOI
1Ph1iBOqszVQbBQ5BFRSpbZvhmVI8x3EeJfLyT+35gGqzcBa1qg03XJ+qB38LSyK
GLZamAdYZ9ukNZZ/3zfTNkbTe+cud1EGDofFVivtdDpDqS+9Hq5hFnFDnFsEUZYW
YS134qNA56MmkzCTTeue0Y/RQsaqyGl+kIUsEpmJqbj7z4ImN7bYs9Oa/yYUjzwS
1qeORLslxd+fFkKylYeA9mDV7u9ZDrE0GOWF2qhCus8EhGhZD1I9MH6EfNTBBy+5
BY4GwWlnBSJDPieu6noPlkQMyxibbkiUC+NotjAOuQ8F7VdllJaB9gez+h5ZSfyy
5Sz5vKslzkmOqlRYEtBdWZ/xR/sqhhhbPL5CE/CSGKJMpFG7FIs81KIRW/XwevOk
P92i6sST54v+3+3dwJ3WZjynRkaA9bm1MgQvkOFrgRtReONjXm/DLx6C/zsATDGa
LXdljMTy/uuXNd/4XyXN4hh/ttkgLIFYEO7ER/QM0s8XSpj8mTSMlb9rJdjUDZmg
P7rGl6ncLFjHE6Uxqw4ZQcqx7iKOg2LDDKxhXgDnYYSxcFWTuE+y0WzUqWqsabgm
pInKozd24HZvA/RTq+f26yl9FSkeqm1+UIWv4SIqII+vx0iJJ7zi5ZX7uVNIs9ns
QWMCLlPwrnotmjscq4olA4lDl+Ke58dI1ZkWlkE0zIU1MIm4o3AJm2XRAXk/NJQ7
T7PIG5vLN4RppcpNlxoceaFU2TMLxHvMXAVr4Ie78rrkYpJX17PO/OllpYZKwoqv
eOT5fEw/O3NI7+p45xQllHnqDFivehHUteMjuNZTEcTz+pYCXIC8QX+A/qX4P4qy
lYR8qMJCYmJTBcqaaJZLrwNIHO/KBRA8jl0Q/4GKvdmwMwoP1fzyFnv9YXpna9c+
/JWzk3Oh8gTApk5giVP5nQbKhXDR8vbCEMw797Q8l5K8H61baISnSJg6eUT+t+vR
maSmmsmJO+nDkGdSnuwEig866scpDGdxnwboMFw4oLyvgotg+3sVeWOM4m6Yg8hh
8M0aSZCpaSdOhG81rwoltDYlSbbGwjIMf29vWta5QACnq76Wb0AkvvH8VPAgGESV
xk1fm9B2hrhJ8TKLTdZdWWaEigfny174BvOMkZdJPMTXOYuPAmn0hopiIOilUmQe
JdAvGkLdLXLVwGe4nKn6x8Pe//Nb5DQmBXbhpA1/dwfbbBAWfWxXQ0if8niglnRU
XwdkzjfKZAxg6mDKA15W+sUZSwIo72277+UnJ0EBJh6UrJZPUBofybwBoPPE8uRP
47pyL8QKdTxvC4+STzBc5F+uooHRz7F8rWzXZC4L3ucFP0PNSGiidosd/mOJBGUz
X8p+u/x3EmD5tGpSEoQ7RU4ZLv3eub0aTGTbsFk6879JZO6tcPbblxmAea16dO/r
NR8IVgeHuQ1DEhufdZdlN2fXxDliMI/YRh0AHmf/IzIDOYHVwTe6Z3mXpHAmawBD
dNiyyp3Gr3JKrJCgvlrQAJ+QWJE9QWMyLQ40GE8wQum+WRsJLkmn21IcquG/2stD
fTGRYmarcI8c49igUgCG97BetEu0ZAj9+rRADyaW5BCstWJ05itkijnFdOdIOT42
htvf4C/KHpHPtRazbAqN48R90idcjCtXnk55SIRl41Q0S20C7nnDFxve04aMvadZ
lppMu5eVP0FovGyah8tjOOm4QXaCUb7gX5gSV6EzG2Ac6pcPt/5oqQNfms0Vj+MG
NNDt9wq+tD3T23GCE1Hq/bmOwtn40wNYBF8vaf86ARZoX4cSuyAV+5/aEV7tYvoj
xJhdU3h2f7NvsffJtxS7m8HMHXBZ7PO3xsdUZ7PzXSCn1w9sHrOFdcXIi9OAheTQ
dHH/CAEViTXCb/lWp+oZO1OePmoqHc6PP5Lws1xICkqRT+tzEX+ak9MwTqg6/oLq
q0yynGo+7ssO9mbKRah+oUVRH7yS51idHCvmfommZQu9LsWSxuMAPYAyOEeSINKX
0YUYETgObvBlbbZvzkrWxaKWKgxrTn4zukxf9oLWYISVPdSSpXITs6mFgGaFSXcO
9Bm9h44Dqim8QztdqdIfxSN99lAQRMeWUTAdJh4rkJIDZslLvcseg8/nmbhAspEw
fT14fiwOo/tGh4j7RsqtZCWshg/ROUQbgxhPULOlFbbRQ5BfDR2JiR86Uc8J7UU4
RwLNWzc9Ccy4P413f7O1OJ05RTP0dLPVuShsSTV3gt37h91CNxc6J4qbGdG3S4Hp
+MGTX9LPJ7DvqrH7qHnj2GnG6eJLQIKOWmWhXUjOYLK4HbOdHjcNQxGva6R1PNHl
6nL7M/c36sZqjsvcEmwTwP5QrgQZ3fqvIk/v0NExIxDVci1BtmgL17k09Ku5xv6l
tp21fA6/3fsz1VtW+RNb2UvCnEuAfJiync5AYBRm6ahVjO2KAaTv5cTtDg3FxAK6
/kBX+xsj+KqG6hsAPDb7o1h9vQcrbWRz/iBOzUTm2wXjDt7ga/OabGYcsThJf+kP
Ka+kYSlAFvQQbF7DzEJN7Hjwh39w1Kd4vkasudp4evk7GJH/3hJ2AEpAYzTfE9Dz
aeyD6iU9yID8dYWAmt+yVedIC1WFIqYQD6xz3MJ4mq+D4dATUcE6m351OyesGoeo
lRWQEHKIe7gRDz9hCR6hQw6Ie7BuW/jPnqf0j8BFCHF/zxMZo662bN4lIMXwgi7y
bz+sl597ztoYiv0cwelkQ0R60GNCpbfKEcMzjky5Gg76vDr2Q2D7kUoFbO2u0zqp
0jQEVcrMBdIchwGMBdY2B9nSUt8K4jZawgUZ+xrPCELwMPTUQB9pxnJxSjTX5Ii8
KI4AmVMbC2eJDZQZbtoRJBGkMpqkFUFbYwhM8L3TtH5ga+qa6IOHjreUOQ7ABo9z
arFTYMYikweCMzcOcP5GKOuQQ3txkpoweikIvqXKwgcpcBzaLsUtuyK/6/cI4kiI
iAcKwF6sbJhLkBIT4AbCsGiz0Stnu/MKzRej1yY/+MmqSV2T0Dmc1Zy8tGuZ3ael
UbCWfFYcaJk4woSgeWLFCOBppNPykd0m+/SQfXx4EIy5U5STAtPVCUGTZePwJqom
CHJUdjJaQgofiXnPUyJvuHvA4v/+sbUs0YGii9wbRXQAkDqBgXo3ASSCaygZBour
BQqUS92pLJVH5OXsUa/Zp3GH9ROkGaV3YDekCZhx0dWyh07fmBVjXJGmW3U9HzVC
JHfnYZHo7P/hw92x0uDQNmxCTXUMG898JFuWG9pnH7HXDtIN4Qi0WeLyr+zSJuSN
9d5JJODIio+h7LtLmX71v3ugWomhGND4HM+NY90cmmUaaV2T0gwMZdGpDxyguFY3
MjTddHMkquKL2GJy1mMAxBjrC3kHgF/ty80hKrzA+5CL0lgMZH3b+hILDyjCAKcB
vWALPo0PM0Gm6VrEImcZo6/qqqDmJg1hSqe+cs+Zc04HYsbjKAK7H7VWVyYAyCwa
RKPQ8fCrWlb0cqoCKH4+DUopuxnZJiORuFlDQht5fMyokdOcKkFEc6Y5cXUEQBWc
SxP64hKVxiFa6UWA626Ly1jY76hoo4x9QmPlDsI44NJKHYhrsyrsWQdlKWtdHn9t
mniktCV6XZZu2tnXn2K9DmXpSCkOCo5RE157a5OpCgb7iYcEviElVp+j0/UrDBaj
qygUTAvr2vwBPIu/Ns4h15ke5J69iW2GtDsR4jbDgOiCApJFnScsa2AwbcItBhJ5
XaIQamFOrnonZ3uUKq/vHAbIGVRUsgaJFnx0fzrClVVGyRD/138wj7d9nNaNYqbu
PkvEArHjrPZLlIqEO7mkIRrsSWaOXA5RSXIEqdr3u2QUrnbu6bsC76YoSBj9ozKP
5kC0n/WhcktbIPB1eG/ZNyH67gsIOGmsGX56Ekh97Kk75+x3VxiSSytIyJEogAOD
vNbJuhdKdo2oamEPyV0WrTHW9+G68meRICF1n3faNqYiKLfLqfjAi2IBes+JJTDQ
nN6ciaQnNlHyBv5JdQVjeWxL8Leln3TKe7XWgvHPN7mSFRc5fhS/eACbQfzHHNZB
JayuSdhwBJO8tZk7RsQw0zfPx3XuNwvZzOkUITDTW+oFE7TqBOW3TIRHW0IwmJbl
lq324MrpJy0lYS4VXrfJUM/GMKFzIrtIevaLrLnPqn+35RnuGIxYrJvoX95mA9/P
rwOTN83OFzF25ZyQcz2Yq2mZu5ZfJxY7v168sGpWV99ji6zyDjWxrFWbBdv6qhfo
JIDvxtpgQ6HfPuUApg5nNg6sWokMghFh14/nurTPG4JEPFDfol8Snrn3QpEORzg8
KIynSF14j8xVu+V4Up8mygMPzRUUkGZruv8/COSKQnoXHuTADBABUgu6RMOOnR9K
pXZUGUKHzRle24fOS732Kl++hH6ag5O/08ScF4kmnxDH/LnkfzzIOiR53rlYGJNw
s/iL5NYyKkKAHA2Y7sqlyRo+ctARoc/uvSW2Je9uRe76ELJU7+hPxGGUvUGGCAHT
/hxzbu3+CnlSkOtxuk3JsKJeyn/woRJNWQlEMRy/B+eiBmsCgdnkVAmfyTpmqMMY
bLz0Wf/JUifPG2pj8dSxK656Pwm58g+5IjN5NDganNKtVOOWa4fMlcaqNAhY5/Fd
bRrNBO/zeArlnYi/nslonQycIIYA0Gh9tEyyvmNL3+KY7q3OQs+O70D4yyLJkuZ1
sblZQpG1utZvzF+P0iZSu1JSuivU5Bdhk5u97OMmwsEBjUDEAEueVfxFM7f1mM8n
DCQZP0gBM13I6+Em2vNGGqFFfJd2+NGfOAkVEBFKXG22Zab3mekF0AIjvKseR1De
/d+VYXLEpOBbgvPhFLeU1wm9aQ/peW4HZDyE1QEZZLW3VrE6Ck2KFzI8NhLNGcLS
5aUoVQbqluo1pbSYEXWxU8fHIhZWGyPip5CBSY5xj48vpPzC7FPQxHAP/2gsiLG+
RGBfpTIklQVKSItWDOwU+2V899+ZQoZHkKqTcXwHFX2KCfDr5jX8t5o+73T1xXBv
3xbSlW5bCFKu8Dz/PdbK9Y8dgT5urXTUD0mbTbpNP4XD+3QZ94fzmVhrBtRBSUqr
7s1zjlDy0Wi7RfPi29NEydrvlJn7DFROen1CNXPCJ2+O9okhCANOyeU3B2D6ZeDR
rmTf5yRX1PO9UvUabRLDHev7yNQe/D1wS5UtTphAz2cgAy6jw83NuhxlgG89tEiB
HGyX4xoFwRme8WBIv0I9Vxuhd2VOYmSMOZKLNkt8yZN6248LdFsySy26JaL9AxF6
wSQR3rY1gOwKDt6fMcZBWjAoDAQneXuWeH6Bd/SHzoLTlIVGRcJx/YRKpK3QFu7K
wzdM3xB3yIeZQ9ni5gTD0grvD+ZGpjx/gGEkY+su/dKvzJSOcCobOB4XU9UJCwHm
pyqN1hNcy1S+1ixfb+g6UeCBDcXxn3BKPArksGtn3gf4tT0pEfBiLaAIt0yt05QS
hL+J4WbgdOfkZNEf4rkvGWjJVi+SxfKkSc1lK/EBgv2LShiHwuUfvJJ629PfLvzU
pF0wTUqxOOfCXbn13EIRC2EBDyuxBvnCWHrDIYPGtxeja/FnbTYwYelvT1gUzEQ7
c3pwxslJH8y27x0DAHMHWgR9LAPdGpHt+D061mcjgE+Mie4eSCdY2/06TIhwyRpl
DmvA9xJPZBGoQ5DMGE7L8jGJp5s7eW54ubByC1Jhb6bjfGYz9HjAwj3m+nVpcUdw
eQhZEKGJOt6Cby4QwJwDlG/mC8OfFHvxHXTINAT80Oypm0z0vihbAmmH55PmgTiJ
8RP/siG68uk6JLyTre2zTPWeeoYutI8jFCxeMqWe+Upr0Tc3r5ygq8Qih2fxysW8
aehWKtVNXmRLzk4wxa/kBUwId6zXqvbfl02oUTBDwm9twKindmHqX0aN7wuRY/MA
Kv9CWMHx8k8//7oVyDNvL+bNRXGVOGt18e/Bv0TTDb6S3ID/lX5OBERlZyupGOku
ciVj8dcM/lleTJG67wRSS95GmrtlT6LN9PZC6ErgvITw+ntEQW6RliF5/WOHbsWE
czt8+vgj7jh9JStCGNzgn+oC6gdIOAaFbLubj24qhLwm4mPOj9IkB6xJCLICWg9z
zHJGag5Mug7gVXR2Y4q9Xukfi+qFVTyqfEPkMCQnUMMXAt9QNjnkdNIEEx3VJIS1
DBWOAHf378KbJQicSHWYrXEpP8ASV3AxtCMrs+l1EH/ceVzLS2IIRfitdKCqFCsN
F1xMvpf3pXOy8eJxczfXMppJfs8jtDU2u4Q4xv58ctTKkjegbQkFbN4y4MzYffqd
m6es+wOX4W08fr2nDC6BjilftbEe8F5Aq9JLpYKBSrRKXclB/cgdjOiWEYmdZQox
UkdBOLw0aRRwMzpl3Ir47asZIFQNVyb2oHoSmWHtwYYWbvUN9bG/BH84xxlvgAeT
CtaBN6dzmTRWPqyuaQvm+yPRo/dlw1rKejBAZNlZ6qeGzHlXbQzSi970HUxMN6+C
bQ/Y8gKvVq1l1YewhcTebymjJXZZURCSzeLxoqUU+zP3XJlr2x5KWYBxt2a/yXzK
DF9M/TRNdsL3Qicvhgd84gFqeqYj7QUStwH+O/U1H/ZVzVrdEldViY4dveQjE373
n+vvOELBw8DKD5Zkti8JKjvamIMZC5JcXt6dHM6E0nXhKsJ1mAufQeAH9tNZ6JNA
i1pxRaHX8Q3UqesPbSq2GdBP5sfeVXVzgkF6XtOg6AoOG0l49K2GNxzjRz6UIcSX
6Eq6TcXCC6oE/CYAyrVwLLEYGTuwvo3yfoy8fKO4zHUIAaIRzx/r3G8B6Gj0ZMfG
B0PZ05BABSx3CvF+qO3vE84XoPCMeXsk8hISXEex5ZdYno2utDCqSu3Jt84IS8MD
5csL/oAiVkkNZoJ1NS+ODVhu4Dum/0UEXZWpfjhhzWSTTRRvHo9AxtG8jMEuOoaT
Y3LrcPee0paGLR9imxH+D4aVbT5yJmvPltst3SyvgV0gwkTtJPFQShQRMzev9fSS
jnt5aa1kWpvQRKjXQ4sKMN9sOh5kQPCK95fbLLYzAw6qUjmDhfw1x49jAKuJFACy
dDhz3Dj6Hfv9FXN2ku0GXcKd4+R5FG16yUGBXvzXuGh/SZ3Xklyof6S9eJb5ERtN
f1vs3/Z4zjJP+TpiPII9x6X5uKrCWfZNtgHpPG0fhwUseiRKCdYQ9t6TaKh9iCVC
hjBKutvrHGC9KJiZZdwmq7k0CWICUmIiVJoSWu9xuGi8iMtwqP+tnLyAr0pV1QHQ
BZdXhaoldVPVQCu+N33VdePMzg1KsOzjmPJbvwu7p4eWMPlqBvKCzCCceqov084V
bpAMRAJ8r1OayVVBKdk3pQeswPiK6HxhwDNhXJoJUv5Hl82mMNq44Qao52TItr80
JnAEfHpki2qkRxMzFFzi8bR7Cpg3f+XKpzWa88QI729W9OiCWtGOTB1XEaizIC/a
llPuG+JSEgXOTCarVNqpvli5E4StcsfO8xkSjC1m5IfMFHv7eYm2APDhM/JDxRmN
XkhAwCG8UygzrMMYHmO4Zidqz+QOgD34ymnisSRYi5qSCbfJKht+/I8VoPsWZTrq
MPIF1lM4ueNOOoOWm2Zpqug5DqdKVQZ5vSJSCHsV6ozfYRF1jECLkMgnWPBI7kZ1
e4R6K5lT/YZ8uO6pf2DgI/3D8ssYroyY4iV1izZNMc3oLTJgqFuke0I6LBwy6Y01
ckbde4H6cYjEvh6eHzWqkCdFBYY9McJpvQwIpIs2FGaqbB8qFKBwmxQQRnOXUzOx
v74/mEUqT/QZIMfSL4EhnOhML7/YrU/E+K0hGt+axjdbvc7Fz9JfDbrJ0NG0aL2h
G2PRU29hPk5PEgkizGxcPM1No0JK0Jsd5aIk1D8Fg0eInjGvD1VtTCQW+cUr5EF3
hBVRIX9pT8xuK725z6nKH+Su05My9Con2Q2cCqJPXqTazGh1eW+cK6ttzOy3tr4F
2USrMPTpGJrN0TI+8Gwf9+bSKI9WKu4Gq0Tu9JfqXSBkumLUzwAO74QN33XkLrxS
CYHZFlzlRhjfpUFBkhZdTra42G7SeTjsrcMNx05mBVNXlmsofCimA/uGD+mJ53k3
5yYC9OF5Pdp5pk/g3hEZNc1h1M49aNPb7XA7vrf0HDYaS7bngWkj/rraMkunMTQO
WFXfy65e+ufI4X1TD5u3FvxBar91neyAOiOFKVWse0Glf8TvT4sQkMnToMDMR7CR
87mohNP45+vL1MLlKgHbJOpYytDk31aBjGKBPwfp1jA4Yp6uOl3MXaDwEaRn1D1v
vuUrwQBRHTYnmJuMRFf76cf5dIpigCNwYXFdM3+REVjzFzEULQ43GF8BCmCeuD61
ICIXpJft/UIimoXDlg2hxneFggIx+yDuabk3L6+aoUaFVZSbn5MdMR+dPK43n2ou
GqYKY5WZz44msMigPsFKJLTK93KhQEQ2Mmu3o5jM3aKiCCfqZwKWcxLLycneG0rF
Rg84/qhGmnR4pbAm8SFSveLpFPKMLnF+CUfs2VUJU02k4YAZAGAFPI9U74c+12fs
xk54QrCuFkBywoqNBDvA2bxyVXKCk0YAEwqjZtzJrFVq5Ft/CXlQVc53kC8blRYA
rQPMtPEnr2++pWIPKjKmpLm0tUgppiwEA9p3qgR3pHgaJd7CjTGyIDdDphH6wzDs
5upLwLOBdb0SqQUUN18EcWadS5UwF3q8LEYWoYtXbnpbQlD2vfUeaEKQgr9MKaX2
yV2TEcBdnNwZaRq7DPKcNoEc9OVRnKhzhbYrc808jjI+ZhRSJ7on3tHFChXJ/akH
0YiEIRw3qZkVPRO+UCXEireNibir1vYkfuYv+0xWS3G6vVA6kdOfxCNGWj1sgFwe
9TTmTt/kBTjHnE8edksQrJNxSeBmWrVEkN1/pdJDnwqL83Mi9nje0iwA8u9gsK9y
r1l9LnMERdQopgaT46b607/W9owrezo4fKpY7+y3X9toXw2eQE+CqxPTfnlxQ7/d
Hz4NefqGq5pGa0Oj+7/PKbnHkvoYr6pOI+1N0+QuXU5x0SH/Ol0eBn2O0P8S8RAP
UggxbAR5hfeVpGyG6tKa8bSEWnfYqzG6G6iYxNhmQZU1AcwMmxKTZ7vCPEHwikt2
fhVogiEA1ut7Cd53ZHuFhoLUO1osEvwF12S/ifwFfs2VKFLMC0WfSt/H7ep3OcR2
TmwpJcEHvCaCNyXxBjkJTa/e0abZDNsSSAh1m7YaXL1zJXUINE1GEcgm/W3LCIxa
d0+p0FnPiTIXbg7QW9fKmhfwiFBFdBLND0T3ktQTdI0EhuVJ3Zwcqk54AJolikwG
Uc1hlSKWNeWSn/P/0i6mmeur6DEh045TAY93q/IqbHk8l/eAuwOeRQzGWIs4EnEA
UQ6t6UJE8dhZk7Bx+NdhAFLOQfERjaqfuMpLqamP1NFEIEUektVGkoeZ4tZRXcN+
tWn2Id4g/j0uCWwU/OeaGdJCbSyjzMJDuOzC9zKQG054SkizZaOdoB8lQJu+9qIm
W8qhVHH72vVzVA+O/7S1rVi+AhXFLzRKwJNsRyLfWdbPtbH31AAGB8ojTR6CuJvO
tLUI6X33J6OM3feQoN96lp1w3ZnqH9YxY8Cg1GQrXaEbzRTzuE4AyRhLB+aGTTm/
bEMZyNzGynyQEdn99pmpptbEqk8eYBsGqTHWLRT/jOI1hANRtAOEnes7WPNHN3Uk
pG7CDFL8D88yq6oLoVrc8g8BR1+loDlzSnHyhAI2Y4uAUvlimVDNe+W442zi2QH1
YlF4LOJG4H00HilDSmu8ifI8Mu6ZpbRnvAmsUxEdKIRdpRGcUC/ad+Xawae7TWDK
X/msHglTcWy5CjUkHk7Mf94RHuS+cMzpC1wyty8cXFAbRByBfCxeWkw1ajFV0Cr7
B6eElnemF8guU5LF0QJGRhTYHy4RZMYJFN5ORMhA4mhmcHXwRxBsjdGvyVE5VwQm
FGH35oyvj7iUwhMiuyYlyXiv0Nxjc8c+wGvLkdFc08umrdYkGjdNdB+zNtskMOwd
W96TFIAEgt8v+/twkYs+DLPRch9s3iUDEqVDsEry1DVWI0w2xe/DCtly8uH23IMJ
NSJcvDuypyovbLFsT7qk21nXFeJlVHimzZRf6tuXgkCifkFnSSXpZgpXgpMjdm1z
9sZ4jXX0iRQxqAXbawq7NzHU0q4c81J4L4lsnYz52FmolClVB9q8AjPHPG/Py8JW
mxjTfn8X3aU93eIEplZ4fPm1MFxdK/KkWmTo7FWCt3hGSKwHZDcSVnaQf4YtUcTT
JMlb2FvGnb0zCzFNrX2T3WB01Ehp+zlKGS5MmfqdXAE6ZHGJEIHWgbetUPS8y0HV
vZ052VDnwL93l7OhkXnvod1R//ViFX4RXE1lVDHwYnqpQ4Wit6UPvyUkpquTfsfC
gNv3Fahfjk7ub2zLSQeMTHbBGUbX63zRCJQa5Hq/YGogNb4GrsMYvzFSmSBtf2yV
sZ1RY3npDOyZZMIkK7SDENEpqKT6G4qviiW642Zx+QTroqThpGVPshXb12Uky88k
E/Vr9TvkREyQ+OIPKo6euRryjIu2Ebfz8L4owSDFaqPrwx0gQRG8VLrOBvMQrkhG
6D/BQ2modspaFlzk5gjIrTQGtji3VgobOLQOhrOO3Jn3ZR5J11W/F9EsoK7jY/+B
Skr/BkU5Mp8lvA0/17VU///3dI0iguOmIHMVHwlUSP+3nErQ8t21pog0mfp6QhfV
`pragma protect end_protected
