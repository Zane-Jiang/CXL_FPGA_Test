// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
JI2Q+KFiE712/MeWZI2zn20+5A2LFAGZpzkfffXeAXKOraqieR7Q2SEqmuFBHHev
xDAy/wJ9oVbgIizg2r4UIRm9veLG5q1/itq3MXAU6PAQRiNKtWpttt1HC+7DKjNM
x/OhzU3Ua/M11zVrKTgZ1xi5oiJAvkPg3XQRaZkMr6M=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 11120 )
`pragma protect data_block
7u0DENoyged+gzNlpD7KhB165c9vbhQmWm7z9x1//VbtefRpPrVfsZVsuPpDnuC9
fOzJFYDCs2G/BQ53NpFzScsD4wLNBFq7f25HDqhuwmoUfVrcO4CsTsL9tBUYt6uX
aIOikabNFlR7d/6erUKQ/VkvsEThH29nDUplhZ6HIcXmMheZAxeCcGH1rmPB8uTo
vjzvYGBrnoTsVSDGj1xZqsMMhm5yrNAWP0cjas/J2Bh0iR7EDpXq/XLnR0kHUNzI
sgueutkKnjeQaLUISIM3xRBbrmXKCDxSZF05APAzTAAtxbAYjm0Zsv3+45K2XaWw
WBJ/Pp/RlH0VEIjiLRGTXDndcYusAXmhwwraSV+S5tKar+eKwQPwdFWAEOqpUaRH
rx3XAfenKeuO8aWueWD2fGlKt2tyI324vKv+ArgnZ8oBrhZVwfcGO8gMXahTxpuH
cdyKTbEH3nvx0ulXV1xulHihVKy60OodnAmZMQczD9qeB5vTTnhjEYLfUs56ttmp
YjPX5+X1Q0JZi/ctfO9499nXi6nxKwNGrurAph0lVfmB6NWzg05zH5gxg4BS3oyj
dn9MiWDqQpBTsKGvTvSqZDnEbHb2YiKCrIA6TKpN3eg4XrUEUcEoJhfTsNc+m59s
C3ttfknEv1O2OnFM1jELhuFiB4pfllIcVE2tk+zS8mxR9jBcIcKaVTipHtUPFjUN
rTpUILglO/sVEBUDetSlxUIEAVrZOCxtQRqi5RGFZr7mPqfmpji0xcN8ihITYehS
3nII+2VBTt6ho/kA6Zhp71Ieres2ueifvw/WFRJqYS955fkhKUpy/oFtUaNlC0uo
hdr5iEsKAk6/wZPBadWOvr4o/B5DMKzv1DMLf1mGmwZg7JHVeHeJYnSAPbNkck22
2VqzYT9psV9l3TFe+Qfkrd0F7+bga5OQ53+X4TwFqnUofGiItItGN6vzpxDu1vmh
MY41d+EaPuA9URXW7O6dU0hpC2ifiM/fh/ocGUgfZd0oWDEBUbdQtTHKqF3zLz7B
DM5x6TRNdqdu2er/oHl/FC+MJLnElQxg2ByoBPMrD7zl8+R5z6KRw5znNp+95ZPb
+kxx29iXB7LFAg0yADnHK+d3+/r6fo0ErJCpY9TtvX0VxmZbcYhlNJ/KvMBhcqPZ
2PsTXEkaBfp/OuywnhWNEiyiJ6CzQesSR/hOT//1hdGhok0u8epcoicwEkaVXCgx
17Ckp8FDsvq2HOdTdBiWupP20hCOEnO5zNL1InVWnHZM6TgbLr4Ni9yc2HwX9FE8
gsvQvaL5Yg4Tg2jYE/b3Gqi/ctnMXtvELQN+YBz6ZgJOeLBHu5XztEdPbNlVaoCO
RuCloQm+2Ah6/L3w3RGWmVpWEsZigxcycMcVsqTChC1COgdhvl5Vg9TAhjOOOlEp
v13ad2ymRD03Fpa3PUbCKYaEfc15WYWbAC92F8dAzy53yKHqsmJyt6MIVjcvjyzy
iRipxGMgvFLTCDkROYv9SAmQxE+BfFJKISn5eli91p8np7tmTVrAH3hM050D62n8
E9b20yj9uH4W4tTC6l+0sSMTj5NEpfc5wT9E/cghp4SFcvhNITtk6QH+E5coPOiw
Mgpa2y3xAIOyzSAcM55YQpTfOTgERQMX+BfjZVPpHeNJj5SgB0ovyfu8xJul6q4z
fhrDxH5kDDWcniIClQHUsziifKQQRC22j6xdP1HbC0iLxYF7FP2sEABKJfVkJC3V
dAJh+vqKfMb/7y404+0z4r0pO0A+Rhh33ZHdmZFrpEqh3oinBuMIZR9AV6iXFOCa
3YIdz6avKtysmqJI/3uDSafACPQClsMtOHGMr3i2FaejlXbaK29JA2vcWnzU2TYO
YvGb9/9eHEnqfEvSkdaYmHc0cDDEngJJNmXBCrpB2H1Op5Uwy8g9kl/uz+lHDRvk
5A8Ij+UuhsRKLPZRb+9QZZ44IKOvgEmtVK74AP6cwQ7oUQDlQk4U9v9e5tPNyvHa
PQOpvg8xWG5gROW21DsJ0Dw15Qkdh7LdbrB/nAqBNR0TIBs5JQyGBVNYhxTdu9Ga
IIrCiUx2MscRLJuoFivCqNERbC/TnW6yMtUNuR6dz7H5CsWRhapBwYNocDPG6lNO
ojB5S8PQNsOaB3J6pNALn+QOZJMaxdjm7IE4uHKHOl8FIUR8Jyg63V4EWHvCvTXZ
oR1DkAF1lUmV7nnmCGVr5+ivoe0xVj+6eqXCh7IdNMabO7PFe/18o+ldsBhH+cae
Idkke46aSIs0Tmmf8Ngtc5m2NEZgcTtRNzGkLRL6VHZs/1VxdnvTAzAuNn891RRa
Lvzh1TgPEh1Qm+Gw/m7pNF3ncEWcuEJp9JSAnPBgQTmxTKpTCB2DDLOlaeSr8pAo
O4t6//f9aHfNeiBvWR5T8d98zszCizhE7OWISWJcMwSOeIEVsTx7JIvU5olYwwy7
bF3OvCZ2HF8rjHrO9Dn525PXjawv0+SChk/WMBaZOqGF5cMngVaAjDJbpHJ9M+Np
an+PJQqKGND0WarJ0nh1+SliAw98SY8LrWuag68N6jFAXwfCsa0zV9eBVz6Gz92o
KdcDnw4hlPyAY5+Vd1zu9CaMSSWflnNCJptg+TSpRvx/WFI2WRtMD32gdvhfLJrh
ZOtpg2Vm+mXAduOgVuFtPdtF6NG4TcEAYR9V81cTIfe01Is67PGuaS0aTVGXtt/p
8ZPX/phyc7qGfgZ2/RgrtE07SJ5IWorEuw5mwNQ9qR/GIaWAG0/VrqG+EZstPnT0
78airRL9urI/EArpm534XukEyu4Dhk7RA2voCSvupUg1XktEhksttxXkiTgIC88l
bK12FFTs35twQg0pEdRFKMXgpnEx0/bc1T0HNYcI3kN7QmgnVx3KqOJ5z+pO0Kgu
qx8uqG1tIt1QWENS5dPK4EsGHP0B1vOy9cpuabdSUUMoYrkU22+z4hAdjkBCGjRs
l2jK22JLP3ouF2Gy8XTCm4prhzNIL+y3KSlDAmGa7UsZVJcKXSLtRvpZeB5YFwxD
7NC/5j3oXBVkeUV0dx6Fd0wJsV0uy7AxrQZAnKvUOrbr3nRDqtZlry49YG4NslAQ
NxXWxOCUj5/aJPiFcTQjJ930otcaPwilpVyptRK1M0ncD0NXZk97GCaLrl/5ag3y
HClrvflwpCL1d8/ykoyMoTnKjUYdWqdm9XjyyrNw/JLikeot8YKziKzJftdVwOet
+JnY624O6b8M399Rp8322BLUDRGlHpdOvYjborja8Gphj75DjcbcE3rJEtdg1JiJ
MxWB5JAxV/Zs/nw9jMd+XDbr7MS/8rfMfG84dEmSwwk6wMNadoZtjeHbbnNMfhUK
f+oHjfzSgJiy8oknNG5VJubVEMuAtRuDzH51XDgK6ly5gpp5i30BApxv1042J5R5
ajesGkftRcHtl5teUxqxbCTJkT0prSL3ZnSX9f07HqI1KocgbGiY3qrnn8mkHCeT
nGkncxAYiIBNBHfJsD2VxZeUsR7mMrmmZ6vK+ySqvAI8vC+mVhOCOg71hXv1OYS8
B83oyJHqR5lL8H4weI77289gxIRK0pglpa6z5DWm80lCAu3SpRw0Ar3Wuv5AN3u9
YwKSU3d5IswEytSpe4dFkOcw7e5tzu5wPLLxu+u5uVJRF0XpiB1/8WMUxQw7CNo8
kotZ0abHCVZMPqwhBcoy5q6T6ZfPWEThgLAI4kRJKL2o9NEO2yXb1kAcdX73l/KQ
W+cBS1kfM7g3n8+/CyaFwhdj01pOqGCZcttGMpO7An1Rh+JK3fh282G252SfFxo5
dPkZqczWtth5v5VCiloZBsjSbCDDf/FebqKwUHZraYwiSGtp97piFylkLpsbESlK
u4iOIfZLxzS5u8WThfzrnmY5S1HC/uBFVEV+XpBiMh4IBHFDFjd1TQsraZS7XGnJ
HFZRY7ocicEOl5FxLoVhfPU1wcAeQxqdm36tqazSJeoedC+iriemVPTnR0+u0iWU
hK2uv002r5XkM9kj/rc10TyT/Wso4QHMD8axJjRNDxkXma9+NmgDoRBbp2ApUiAZ
CtN/e08LlcR35EY77DuICKpI5geFFVNLoWrXOd/M5/r/rZN33e6wBL1dSoRBCZKE
tRiXmg/r+JMdLOsPizWSR4ab0DJR9WK/aosYeeWkzEh/PYAmXceDCS0S5aQv1wj5
xHB3fakPlsEPq19KI3VW/41/saCnkxulCjN3aYiPXf2hGJ3EXLBUcGuUyEjURnrj
NKiQS3u+OBXCo3R7QfFX53g1FHCTRi/AdyHJArCwqnB+HMKD6AukSJaecBKvFlkd
IygsrSWD7wm4eLA0nda+JBP5E2UGD6rrXwa2E7AA/x3jkqnQg5lb8R/8pZzJmTTi
WRLuY49XE8uDtf408+H12hDp4Kkc8ThG/a5Uv4SUCSuotnFS9jHCXwoR06EZF4lM
e0Q9/hOsk3s53WvAJcZumW6WnvoqpEfBSWR5NGMFo8NUykIZTMuarVhp+kFOZe/k
SofCIdDo1Hrpvv7ZMaVOrgaiL9i02pyLwPy20/+ZXXLT0vYggz/GJX3H/HK/A7Dp
RqAObV2BoHyUhjQPVX2v2/B08crAWN3SqmHGj9Vj3jlz8e3tTZW8J4tf7OoOhs79
i4QATfi7Aq03DnKRXFuwRLRYm3rNCtCu+wjfi5gYP3+hqHHEctEIMz7FXh/lHc5q
SbimI1/1oJDVXsK0qmUirb8RJkg/I23PIjHPwtHt0g64CSJs7bUIEqMAKE/2W5ZZ
q2X1aG0nM0X0il4WEj9jaBClfR2XijZXVhJT3SDSW/q6AO999D/igLoWmGzd6L2t
7ABW8UAodxF4THSAWbCLclaSCJI0co0pvjMG3OX9xg60hx8xosxZS5cOQzSfHvUv
6QoYTFGakcXcRVZlOH4JMvp0c9ANPqNDe858HWr6mfTaiJl9ij/QYD5AUgnetwrT
lJnFSbxG2PGwVGXEQhbOvZNdkhVOcvLEyiDSL0qHHr0EAE3KsvjK02bhDy2Y62wF
6hnw2z5JRl4Iad5oQv31CkGyyibigFBu78jZps+wqFWYQpvNjzPynihMOBHVKnbr
sFPBtX5ZvMyYTy0kHr01Hlpotl6CvAxbo0V3oXS+hQnRbA9JjxhGRMtqJwMM3J0D
ePC2F5Nqjtxwspz4vjrSA6wAzSGi2+bVpPQfCKPFFmkjELyZ9Tlkd9E+JPvhVnab
3aIeLUeR6I9D4146WbxxgaS5wHnbsanTMz35SIEuN5uPx5IJ5iKGhNiEXVfubQ+/
4mPaedE+tYsPJ+ozK+UBZY/d0EkUgNlDZ2GxIh00VO12IHq1htIk3w+1zJrpTlGK
O5NUqRdsHfo2n8PmYgQRbX6ZCZDnRJLihqNQQ+SM9e3HSrdMdM74VLzOT8Uq2xRg
JuMtKGqkBsGztIPV6wNkjWCfAuCVs6RPPB+0FkiNKLfR87YNTZixzIZfdNu//xg0
kc8vTcqtdPyDCNKXU2HRziUMoTfxHuYRs6f3bxdbmlXYB+VHiyvwOuJl/r6mLy6B
9EGNJcqMqb0AwC63dqEOih1tdoGkoHv6IuD7n+qFpt7KLIEkv6YJr04uKkXwbXRE
r0fEv8OAITaYnb5f7W/+9effc5hR5Mh+56MtWaXgOLjboWHa9fw2rcbaSvdcFXGD
ycqgkHlhir+b+qiQK3xfRdN6y0tp3Y32tBwJuvz1d/8rcTBjwWOy9DQyYreRCmLM
iBYyIYbv/NptpHy9V3Ndi5o056NA/YTY8oXL5AGGfQ9dBEFSnjrnvxYIoKvOC9+6
T4KWCG5Y6aH5opabGONPDy1CQjf9U7jLH6kbZLxCm6p8HChZqC+i8h6chBh/m6em
ML0n8cdX0lepY/suKbV9gZxEfiNTqXptXxt3zEVTXSh7/hEZ6je63tTM25CHCaCy
W+2puNV3zvaRSULP0D89LNpvUSuMZ89/s7FCgADCvoWNyr92593rKfU9R3mx/xJO
gHkJUX91ImhNK1h6ywex4h5H1ApoRrduRITgJV+TLiSGmDMRGAsizaa/8fqVhrzU
JbaMl5C48G8VttJUvTopJDGiKQ/j7hn6duHFwIl6H1Jch/iUcaFW4EHVtsqOw//u
ds+4BtfEmcId7U+qpou3HYugJshf6vQop3El5avaXewz+fBX2SETB7aUf9ChaTTV
R7knXE0oYYD6kOjfbFeH6+rbyjR3cFPEA3cxxj7z8DtmUjRmTDtWS792Kkpv5HTv
bMFhqrjv6sY5YGadFoRPJm3Z7VN+W7cB1FsYA2xqcnBJANyNEa7YombatlraZDMG
7+/bPDbHoo4zjbE+tLiRVxonHA/j78ZTDcvfGn1rsR08a2HTG/RNdnEn7jzzibfz
TMQkLJnR3qkEgLGiQ+BUTtNpYFXepgZpv3XLYs15Bgst9UWv/9t9gFBe4xskcGw1
PMo7Y/2BmzglIlOainnOX/zcx2XhwUPj5a89hM60VrHVX3AsL6TtHSlLwPYAGxln
3Ejfsh8CRSi9eNLexry80FVc3LwV5Z4pqnDnkVbf7GlXzD2LTxM367yBsBpiQwXM
ovToNA+1bU9YWlpADAQDM04H/K0L/umK/chVQfvc4+uwhuY5HFGg/dXjIJaYO0Ae
2AC2PijkQCjEM0oCk3awCqI3sc/cFqpF0jJ3RwoKrHnjI21mJ23UiZT14j45rrxT
QhR5OyQKTGPhj2GYVS5uamsKV49yNTFtwN4QWCsPyuGoBdjr2+vIXp/BWXBMaLT1
kVFHIHlgnsQ7mkYQbmLagqHb4MATCaSMHQKjzE1mYwuIO/VbXrqyo4NYdftZq+8M
ZNDmk34pWPuNgArin/2kQinpBbsQUZ3lVK+VEG1c883jtDJpSBPt5Q6pvdhgU25b
V87ZqcxhSqkSLeVuHwwi3c/k21Z6I7qt3c3X2SH0cgGxUqKXGSGc4vVF05LeU5zH
4idN9KzdlzDLpJCcSbAD8cnwDVp5ut6fD3siHU8Z8OAgafYPJp8qRuRhRX4zy2Nq
H0ZGY5ituGUwCEvQPSKfpjCotpw2+0UO6gHf0IgJcTLz5Mpf2g1x7jypf9S/IKp2
pEdT4wMeCk5zWpUkrscHhERhKQOpAn8tzMn+8FEUBuEZCPiAkI41AYLruUkwHO2Y
UYS6HPTPnQqdwlrAwYAA2s8Wmp+ONFeTyZD3NQC07xgfYDS3V2eYJD2NTQyjg0WE
8pQrqNJsqsOJej7BgB2jG68qPOrX7Y1andZetDtSYvs3duOVkDs6MBsUeHwXQWoh
CI03wa/Cp7CVbXznp1ChwRtaUt8jQxnA9OobeGJelB25cpbJJrICZIeSppp9ERnx
ejKQ2V1tfXgLYQXG8fFlPLHtkgYGg41rA9ZtcH/w/OprnKissv5nlxdlp+al8ckz
JblCa12RILWZnsWqVFWHgF/h010GD30IK/yzO6/Zq0OFtwX20EQxlJvf4cgIjzcu
Z+EsrsO9sCoB/B9XiHDkrhdM/3CDa5Df4KyLaR2gqhfnr2AvhFSxFeo4+57urVrW
iGNANZCS60idS/7Ygp+xPVIFEcJzozxaqt5Ra2CheCrdSeiaEb+M4jvH0llvZcV1
+Z2aGS2f8Y1dKIaaf1YyjZe+HS1gKCZYuEcsurGV+t/o+YdE3MuQI8ifPI2PHv7m
wRCLThsOxuWdxmgKKx914cnmIRxQnFU5yV6CMh/l8Eg/xvWTJ7BE9AbOxZRH9fRb
nfk/7vWnxKm9pkN08WN5paEDN4WKuYsGA3X1hKsNsKmsyzHYwB81JZkPKo9CfzT0
wQiCuuaCLZWu7N+GgUFq0epgrYESKtqXLR3lpr86o+0KmA7mJRnxAHPrKCWWZSw2
BIT81mPbElWKhNcFawQ+JGu5+l3+xRslLf12fm4wLjVk8suC2jf9bJsR0djASTPt
bFBnpYbVMvmYO4aYs4vrnSHS14pq0H8+qzshkJgR/u1mMVfoUPvfCAK7npWYa6+f
QcpogliNpCxQZCGDx+xyfVDwZL0MJyI7GYvZdrGEv4Gqgq8LXiztUF9/adnXFdOo
X5Fxrr5Oja35T4WsPlU94Xs4IuUf5fBCj7eTeOtv59TR12HrPXDz4JnlgysSVU2N
POG+lM5HB2FzE4Zn8orCYpyfjSYgnWjz10JLH/LCvPCzWEyU14lGYk8jwDZsXspx
030bNsE7AU+VnGPc3MZDwVIF7rooIv9aIs0LNC8S9k44oGBQuBToP1XWrfzEO1dv
x9uVaAeuyITWbwFXlEblli3iokCuLclV8DFbrWJK/+/2mqi5O9ubziZE6L5XBKoP
Dh6bENHZ2qjfPdqMRsyb5Bv7d4s9vFtLB3mDuVYGDcYvPXF6rJjjuFLXostCz4hf
DHDLgiw9J4Yrln7AhhpwsjzvwsLs3pKa05ARz0orTdbDH/HbC3ekwkgSasXBs0xM
P0xC2DKIlz5c4hXCTpmIiPPzVBbatqgS1Xw66HnboaFoktc8pTKRfLzKLFJf83zh
IV2KsWwSFgv4PIw73ZdLZ/lyDBkhLFm6sz+qq81bAZ0guGrJ6+5fSFpSxNbgR3Jb
Vwu7uHTPot7WYVf/GQGKYESQ24dtHgI9P8TCuldto0dk/2/FzpF1Zd6ilQEDqVQd
fBpDl/NWkrIEuX4w9Y2D1m1WSYNimmbhRadin3KJk2A8GiRwPM/Cd07M28sZsIvN
n5JeV1SQa5wFlb55z8y5XE2YJWbQ3Cj/xLS7UJtz4U829UO9DSdaP180D0uV8DB6
MOir58/pv2wRWs8NCAcLyEcwCJT5Nef7c5HBzvBUcfCW9SiPt1yqxWG2qrgmCHSe
R2+6LHcIkHJHRec8Nw6vabGB91I5H/5r7LIZKnHIhQE+FwHQ/69KkVc9OQGtfxP/
nwpBZxGJYmTSPvD/GDTXuyY+JpgkhrhOPPqsb1TMOtDvabtQWmdhUbI5P8BcHBaf
glvLz8v7mS390H63HA9S1P4XHg0m0+NeN5WXhY+Jt/GcA5eUI8AEnsUWDxVkFP+L
jRNhHKuv9nPSGnMkKEIoFlKRlDy76RbM9cOl2T1PEVgExl61ys7xI/kteNIkeaN7
TjVo7hyZwUAdXo99jlZp3pw8YjU4UaebQndGEsVLejv8xdsa5brl4h9zt1SSRrIJ
4I2P0TQpnTFg/VRPW9w7y0pPPWoKNwQ9vAXvfCKoAFeAFbXoWnaUIjza4zkbIJDH
qeANeM/cWRJLPZZ8n0DOgrto9Zwec+pJEZTT16I0R52DC0IL6pdIqxCaO+iqQ9gq
NtAd8frn2eljpjuMJM5tGl3qedP7WNr6ET/NKeBDUNvvUo9MFB0P5DMYd9qwocGn
wYRyQdfkBhffQO87UdNiHYuOpu3btLI1NcLhZKImrr/CI9B+m/f6SL+eb6+fXKX6
k9NKB6Nqp25jt+u7VRpgZvjZaf5mWpAh+xjS/93qvlgmjz8uS2737USpVGL5sL+t
y6q0nEXqq8WWsMN0I1/au8/z/xiVLJZOUm9i7NIf0SKkSjS8UaCmrOoPnprfU4PY
449ZI/konwAbxGyZK1dK23Tmf0MfT/YLUPQu6hLJjTvaIfbRYM9KRl+oq59eDsPy
Qs0ywoH+mzqmolsIBTwl8ZqO6FDpqUqDDk1Rfj1fjWV12dPw6yllEjgDaL8s6EjV
rG4w8NutGRiomGUROJI3nMOFcKZNMR1Hss4CsFrDRqdBkE7zcBRgtRP+q7bZiinP
ik58TGGTtei8+kL38S6bKJjPTVtusGDTO1H8xmC7CfWGn/GK0qoaEkS3Cjdi3hLC
JxPOteN/wH4K7rnnnq0Vmr0/Hm+WnkuzYckM3HqaNgNVbGVVuKmzA27g9pOU+MBa
Mk8W9JX5/1pgG59x66aaNyBkzU5A4xyl6eySleYt9z9p3cvCcihjt2DSQCGuar+a
pOBVUu4SAfIjK7DY7IltCQUSN9FM9iAr9iBKNsvGMdFJqYfv5X33NqVpeLgmzuoW
mWfllER2Ag2Xkb/SCURufpuzTrVD5byxp3saudqccC7Vs8S2D/RuE/1NkzzHYoFS
sSA3Y0OZIyridrgs5ZlqzZNRudemyZDWql5YlF+atmVkxCfahD/APm+vFKtrxrfQ
ae/iwekdNXgJhY0jVEYz+tigVIOUDVg4gVWBskrOVJglmCL/wkg8pnKB9l5T308W
KZZasensG/3fd3lCsQNih/KowOcKJaci1cbvLP20ZKWpDPnP8zY8rgDle99j4Ibm
7IQOdZlD2er9SM1SpSC5Zi2thvGFFScDLvYow2D2gcwnQjRGux7LK57eKRVuXy1A
eq6YS6MjfrY4vLaMeUJopfApXNFPk2tyDIp0w7W1r1UtoLXT0UffhjZyBQoPjinE
0yRuk80F0wC95EIsb6D4E9YlkFuzDgBF3GtcLYA75rJtBLONkbdtTIVuzvL4fR7G
mCw17ss4TiEp5G9AajE7k2Dw6mgq0Tu30AiTJaAHg4KVNzvmsiMw6+CBh6ZPA7Pu
p9zrmplSXFlReVFosoAQsdM9q0sEkWdlknm/R/FDYVGmUzfxMcj22JBcQ6THd/H9
Z+KHeoCg+6gZEcTz8Sk+lwsWcnnss4OhwzHIo8tHHqfc6uEIJy440/MShuigzLcn
JD5T0Meo2P0EGiVr0YpA46taIwmyh96OPIZzQEotiNfT/rXpL6Hs1e5Bn86aVZrW
QvsiyzbXpuiZE3NxmGpnZNf5v62ZK3nw4vdlK61yHRRJAXrCpeEqRYDp2SpXUUSF
CrwqXQjn/VkvPiGQ2ogqd6Y+jUtZMC4wZ82BxE5S777Wfv93Bwr/DAXlZNNFUk9/
VqbCiG12HlhBJmS8uaeyf0zESdzJalaHoslP7SeY3AGVlzAmF47DQMQ1f1aibYHL
Zg0bf49/vM6u0OV9CU8tikAdqMZDBVgcGol3Z8AU7ZX/ktBkKwooOF7E8VL+55/1
LFKZ77vGPaeSfB3tqilZjH6WR0CI8o+YDcGn7lD0uPOzyqwJGQtbFsJtlxRx50oX
LpweGFr/nYLbMF0lu8JglUmH7/chLmuN9+dd/7Zis0z81mOQ0fRigNVCTqfToTWj
cOHZGVXHOzas56q9gIwyLGWGS3R9oAasYBF20syMvVp+j/5yJ/rIGUBkI8qi6fiM
Q/qxIjkLGLbf9vU50v8BbqZCdwUy1STaBb2kwoVlN9WPuVdyhfHhA8KEYVAzLiaZ
4nXTFziXYN3GIjfbhroE/6Ls1Msw65nYIh9rq6mcoGh45yRPqc7iwO348/ePcQnb
5arUd7xnsvi/5hIXSIDEP9BFYkWyG0FsFvK9AAeECOOLq+dMXcA/8CmxUHzfsySq
i0Dq9MCkkEv0TbMnIARz9roqrt0uHQjd2K6AgibU6oTbsYQtmiISWJRYnRxyuHUr
g2UpB+QSTWcV/SFix6qli6c8plMKv7RocgpF/zCLzmjxa/TCHN1xLeRzH1UaNBEk
vcGFrz/BFZ4I7En07jc7sHOOaB3HBS6JWk/l+G3aFHz5B9RhtjjrEn/W20NtFKEW
eAPCFYZo8D3M85FbRBVGWX/FpGZSh/dF/kQnQJ6C95UG8Omk78zHcoUi6ARn/2sG
xohxHXdrWRS/aMueKQbkUl43DtCY2rAhlHIiQSODLXqrbIsR3j+qPDR3HccQDzN+
72nCTHkBrIAChEjIeD4t6vJnOkJY2i+xy44/QhUw1Cf8P6Ur6JtDzM1hxzOSA74N
E4qkx2Im0ToNIfwfbPqZOC3k8IYFqqH3uB6gTUeXCx5iJtTRq0861+E9fv9BUqCq
5xSUSARM7Cmdl6Vt6ygmF6UPggwu8SffSC8QLxp74LpKyfPQ5SqVvXXV+Xp3cFOX
ypgS7OKdvA7GXNupL8CGjqB6vrGMURHH977d22gsfP9pjZz66jjdT5KLv6S4yIxZ
E2U09LTuH+DaVoAhNc0umxt2odxqlS3Lkyi8hplBU7uwzZ8251w9f5v1Zu9ynuuM
A/sKTSgQH4RnWTIQT+he1PQCVAeyrHWzKDNBGEePMmYsvE5VEXDD/WcnALS7mYTh
jDP9jnh6+17Bl1ySoRrGeImf1ENZmXXMKPvB1hyYu2FGF86ZCK046JrGGW8BzyPo
cBhZGQQi1dL+hPKW0tTUmnvKf2YvSY5+qolr5BFkWlPWUQuSyphwVjE/SBWYSBGM
6OHSv9Omzhr+FxVw7jObtHTZt6noNYurLBC9TxDdCQKJJ8lsrCs73n9O1ByCzNGA
ADvbWabHgSAyzrv5Hh93rY26ly9ffG3P5HouYPOQsnZWOKsGdDrQiUdU+sG3ge4O
IrGRZD3DEo1gljRLKWx1N6J3+RnysHXax5cGpPkiII+qSfmAnP6cVXm1FxmSNUSu
Fc70Sil+P1Rb1Hmvdaw91BcfwzUJmSSQHk2wW7YoOsV/LFqCOQVIDrq1KqX9RPHd
0rinwboEUpAw/8wfU9oVkVLnw/9B4dDYfK789IPUD20nvC8P+OHqlV4AH/v57Qug
af7gNFnOb/tvyogAobaWlu0V4TBSa7hsa23+vMDdgg1N9+MsAJIZteVDWdGIZ3H2
ixe6HB44HMO38rLUsdsUJ7LcDuHg2aixJkU3XmV3n7yvPLIETl1TmEfDYab2c5F4
1UE7DroUEt90x22KCShyvLvMmzx/nzxI/q68uAuY9q6cDM9lkDOUmtpKGHw0XROj
5kxj/vnkjsouQwReDzC0KKQreVJgqRQHKTJdmtadAKXiW4gM3yjCTgQKGtKjsI1+
IBUwtnvfhYabziZNB+8uF2xc9XhS7YbSlXKsaGBhh8OGOn7G1hKjREs5uekOnwR4
n5xg4C0dzvgPzXOizTfqMgb41KHwUCGkGQbcDuSGzuLlnAfVsXXuG1vJUTUl8wEr
v/fVduFhFXblPLj9zxdfOW9QegS7eNwxD5DJirbXIJNHNjSWfsiXNv2T53W51zS7
xbXtmXQG4yXszfZ621kNnWOdzpgzwb01pNCQPBWZm13mpV4x1W9nqhzdrfzQ5pf8
PgNn5C83nfeGNL/qVzdtHaEVImhmvsZaxTl57l1esgOYKbq2fwHgtkOHMwbSVaQ0
EIkz5WAXXON9gwCoEDM/9i7U0HyhEfK3WLwZ8ES7AQ8rLBSODkQHnDQ93VRwlnGh
StNevnq4DtaIhxxYxjeeJJVqTQI46CzGTcbGiIu7L/NOwNQyFy9weR6VQ4wFw5WT
1KA9zirxkAnwpDh8BDm1ZTcVjJdbkvQermDfJ5/pySHrrrvD5pLJ3GgtEvoFfZ4T
zozs09bKIyyQYv2z/Lj2cWwqORJhgLz3pF4XyHHIXdOXZH1IPRvJM2Au+HqD5jjk
oEOx/FAl3KudfuewhMneVTMbKEn8lmwtNO3FeVQ9wXXQafJBg0k5kq75jXCXgfwv
b+MY6eJ9cRQi6YUDU/LAKDd5RY2Egtk46+C1PDiSuUjxkxP3EhO6xeARtFgYzdfo
MAyGUke1vWnr8gORqnFH27C/Ro9mDKAEhhIVEovKP867FKc6R2nLQVfZV4eOMl1D
HnvtEBRlVc6zOKfb4ltXWlzoWS2TiyYr+XAKTd9FFOmCUsYnRGK7aUngmK0jIbck
AhcO5vE3UVXTfQ1oxgS8OoBkcZ1B3wLh1jOfb/gGnd+27qXudKc5bxRCfTpptsIC
mZMl10FR6n77rlQ5jJjZ+x2HoyblEBGFe7CPRcuybuXcUyC2unPw/P6/+47nx3iE
Uh9lShQkgQ8XGS8l5isTlHsDkML4QM5R93Ah5CEXulVbEyDwJkZ0CScsPGiqaYsy
uyIDKQWPKkgkQlNQdydKQ8SUu8oHJCuwwPl2qmsUR4BgtXld3Rvz+onmUoC23XJc
jTINaR3ZSZPBOBHeP3umHGwR0+npyROXu2rVh5K+sUJyaw7BaXZE5xsggZt72AlW
3lhq0ARWHNGWK/2zQitYM+cFd0Wmzp3pCeeagj1WJ4CC7wnjsGdkmx4WSGo7c0kB
imIhsrg4fZ9uh0dR/FuUlhIOu8VkwSvQ8SY5FMctKn+YxxuyfYc4DNdE5ktDA28I
h5QSCCkaFRY0Mwd7TahzhhemnFQw0OxuotH5Lon4V7Ze5WyJ67NjMV/O7RvTqEIZ
p3YNAnofpcyCHc9TEO+kuN8N7vW/Dkz2ES9bG9IvQcsj2TAiciNJ7MlFMdSpW515
v5DW3F8shcGmnjCLM7CIT4MTRYWfxhZ0MEKRylU8H5fcVIBVNo87HR5TjBMjAlls
PUMKAcXNbBziYo7F9cszeNcNZs7ZF5hBMso0CG7U6jt/xZTlNvKQOGtIzZnZmb+8
e8/NjJcscx2amSw9mHP0gZMBhfxBQMxRFyfYlQmFAC84ep7PUgIvHvGngU37M0jv
rDR5Vp99Thm2oJ+pCZIeR7bgkb+hFyn+LO/8/MQoCMHohJf0o0y1/0lfQMHmhZ3V
A1mAT0eKvQCZ1M+fTse9EVbhjD3AwuAnkp5czdAh/QUQhcRt71NMMutMBX9CkDAh
QVRGswof4NdgS9DpKeDVtaNRFrBs2A8sodJ97srs7LdlIg7uzUUy4bc5KkQoH8wE
XDsrHYVnjNNueyEBkOThd+xCgmJviAh1zLqBs3me/b52d4gV/fAmG5mUYiG4NvoU
K4NYcyJdWJctBKoOniiUvxz/02h8gLARC8N2PgRl9BOqL5UsLvpjD4rKn3TJFI7R
pkd08D/gOP8pHQBKRWl+nVn/CzmnomVQfgnm7sDyN6iam+PAH8UXaHIS68LNflZs
AQVET9bfSCmWgVZ+eJAy0y7u9zuUufWIFj3wQx+Ce1F7G0/6NUA0Dd24p4ph29+p
YlfyeZsXiTWV4Or6MF3LVKXGdoIJn2lM6YPVbVfmoUZ8/1mjVGrMgdHh1lFRhclq
3GQ9npzvRnVG0oLVDtziVN2s1RNjzgdNUPOeT3t12M4=

`pragma protect end_protected
