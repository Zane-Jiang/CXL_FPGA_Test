// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BIzs6GT0qjMqKGY9lhyjf2eZVNK2rcnLnVxssoidcuSagh0br2+u1V7Ltcig
woOsQvdhemtqoEvvDXn9sytgLI9Vxo/J60ACQ10Jm50vt6lZAcV5Ua/6YCMG
XSLM7ZCNsuQwkwiuCqHpZ9VUrG9VaIFajVESK9LcrhLNBj0xR/wYq0LABm9Q
tyWveQ6F7dCCEU3FiiXeP3SAkdbWhuPAzoB79qK2yJpCborfQ6fBqOG++Du3
LILeYC/dA0RswT3YT4fBt/HaRxoEhN6eKraL6upzG2NgfknxnQFN2VHbGIaL
j8eu+HI1Z2OxnY8EpjJnNAtNmsQ14rn6pngjrJH8uQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QgY2ORTHXAszwntu6Ps2O1rVH0ImKXC5cDJpDPEoE1MkOZqorlBXn8Xw+qd4
CvrabwSroOvt+G8oDxI/dHH9xYuzPc/cv0QNdEWjuTAPGocsYlOu8lOLS9qC
z1YtJqNeIGvvRjHTKsqpOyOcU35oDhWbIXVmm7u2xMiwz5Qdmwp0VXeATGjO
yYpCzQsplg7+O2sDpRqsPybGDYOAFb1/isEqPKhRUsh6Vl5Zs35yHp0UrgIN
sz/4SYdPlyobaJTMBcJ6o/ka2zMgcNkEwt3Qht6LtPuxYu1xtleb7C07No1R
SgRxeATQFGt1QpmI2XQPcfgvvvriVJ+GWFLRm0pFTQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MVvhzJQhkpnmaZPgvXU2SjekuXlHT1D8klmqRB/GwZrus7PzOfRSHG6QeHyb
kjpy7W4Zo0qdVjWdBz2NV/HKsfrEY9QdM0aqUotwG/ZxWz5xiMbae7s8K+ZH
39jgb9EZCacqSOBY1YkeFrytpd48DuLA3xnuaXHrfwsDkP2jVRITKGHSrgj9
OF0451MG9CmR4y3C0P/W39CyMeBQxWXaltfoNtfCtf2jxHmG8vQ0nFH/YSD3
eFo2ao5QQ/BCWKc/Jd47H3YV9RQAdQZz8fwmXD5cFhx1rs1K9aYhYMoQi7kM
GsiaBJEBOYrCI28fEaa1etiOUcwBhys/RCRQYyiJMA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hG10tcHSCRTU4T1gQInwURkPXEjKzFx+EtUe/AorNJ+L+fzJol6RrC+SdcKa
tSIqvlEVovDlOFeV7IK7tcO48g0BnFMtPf/G0VM41EY3kNyHGKT3d0q+I6f3
dzhPwka1YP7F1TfPefgwon7VfKazQ9xx95/Kokzb68Q3kH72tuM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GsHDc5aVe0hmVnymw53EvZxSX8u2uyjPUGOj68XxE9Mas7tJt8ucheWDtKcs
vXbhEN9DIu/rqi7WK555hb2Et0nOTWAAn6VIvkUI+JFGWsewfu0uVIb4HvRh
6bKiyD3bNAbhpDn8B2fJehAhro53071JsdIYFanEUwGK+SQVqfE0ol7IBQKS
C/zI90QTuSA+OELLvD/uzjF+m1JGOImF7xA4n+vi0epzagqi/il0m5UskRBq
Du8flGOHcK1ZBvX6f75z8Bpw8UPdzccrvlSQq++2d8G+oqyfRKhju1i2FWRY
ubA6KUc4GR0/eqMrJL2DRh4GSC1LWtyvxbLt3mAhyJM533slLhv4S5t5hfGT
3FvX5TKwC5DFFWiAkbgGEWgi8SzN769l1lPjG2Q1Iu4B+ghWUP4iYJXphwb9
Rx2k+L2Q1KdaJW2aeNdXFSYBtUz+LPcJjQT/E4t1gRS092rh06/sXjObTHA8
Wl++vDl0jkWSSVHUTL9o+XNmVu82FcSr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iBNKrlt7DGUeZclDQeFkqHHjRWLr1bK4qb61HeUjYyeRL1nNsXcZN/0RvPtg
UQFyZefkfNX10pWQ8q8sicSdEjOXZvsrLe4cv2Bc2sJanICdgTmMX7YRF7Zx
CbqW399+5iAZ3xN1iLPg5NgLJ5JC0pkSNSiYXX9//7ZU+TZBnew=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DmdyLOb5KIqdM5oO9ZGP50Tiha4kQJKGFGkkwiWmEzBjnJDHVFUiyD7A95At
KYAFGFi12IUfKKxir9itZi+3ubDq0w21y9IECoxwp5UkILtrypyhpHoK9pFA
F5mTotoXldxZwgD/YCGzSE+/lPJwLLzLMRD8XT2ZfKPm5aqH7ZA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12112)
`pragma protect data_block
dgS6KKzwu9sQfsP+aoJWLV0bI5vCMoqAB3/llUHUiDXyjF5OLWXwHIZiA8Iv
tTtGkERgBAo/ON7FQdMuZ3ZUqEh8orLhxiQnKftFDsgGu3eJUb2jW3mtzxLd
N4x4MvCfU9BibjbGTI1CxLoYqbxdvbiN3WwogY/1H6mkXBTWvuGh/DC6o/pi
f33WSG56PCfjrf/0LNxjemSJxJV4IofWZ2nlfhELPNokiQdr22wNhDJPoYnc
XTj5ZBeJav2PjqJsC3OZ6iMfWgcszbtJVpyG0LAPq6I99kBsRNJhNN36RrxK
428mKRCjZQXh+2wYDpDFNsAr0reYfRP8i3Uzt9EbdUIi4y3IlGTRLWKtqviE
KyhQHsRpbrTM1atGsesGW1moPAFVKgDdSUJImrSu5u0OEj6WO7UKbMHLnVp4
k0+UgvunzPErSiSlxJjKl9xAexL4zz0DWXo9Egfz3ymJltv3rLd8RcJfj7W6
kySFZ5Z3H3U2ePrK9S8NF0sVXuzayt64IK6t81DUJc0g/fYuNdE1ixVDcbzx
hqjDq24OI+c9C29xbLqqc2Trz4C24aZ1uWW0yGNBo56M+mIG6QXJGKhBrpKP
GEb0cqzo+FuyCkiQ0TAT0SmOK4Ql07BY3rVbSXEamzCnrAjEOsYXuEruMOI2
Qw5kmF9D41z+doB4LytQLJTvI1gWBzGZ1ieykA1JP99sMfOdj5keFQIKdqTd
Zyg5S1bvVq1+93FS80DlCzhPgCMZLYEzGbgv1aCl8Uz/trtskD+4rNXPnZqd
W6QxiHne5B2MCMen8m299P/d3CSkb5i4ahoVicmYtxgNNJ5lXUrSDEu5XWvu
QMqbO9NOfTVucYSy2WfanmES1WfIkXJJa0FV93BPjurzo8l2dgMMaVxGnEUX
UFzyfbK6VMS933wjGOTkJuz1kSa1v3r+HWI6pQJwOD4jIrg6oeEhjAjh8Lal
IZ4OjAalxovuUWufMV22PhTfCHoJGvjkCwOxX6uEmdkE6yxwPzuKn1jMZUgM
MkdFbXKpiikYKPwnQwFXp5ykYq/kSXJFkvNq2Fah+1tfAxtIq7rqSvZyCEPV
tXq6gMnhxk109heUtRJywo5LoxGUwRBfSRmt5rmnlSAQ7jvRAcsV1N3ykbHM
HdGAWxhPJcQh85MrqCu0PHtFmjABeTHMO7t7/T7Kdr6mXitDfqIsSyXnQd68
q1uiGJgCsE3fxEX7Z/4l2yh21Vbw8THxE6wFfkFxFq9JDMsb0Dl8bTRhnOMW
PSI7JctACfOVIAZD9CfADwKV3NWfGoPmZqAl3oPGsJc/zEwsvPk2ar8WsnWh
hQLL4hW3F6U0RzCEGtzI8TZJr6hRcU/HG6aaSoztx/pxRCHDS//Q+TA5/lIs
1lhGWepcjxoV3WXKKe7gv+sEJu4dxOKt9SqNsJtqj4V1ucQI0ljtl8iWFOfH
+dGcn5zE6i14uU/Wo52j1E4prqkKBOXYxaUs8pEyg/lkYM6cfj+0ImlBuK8H
YzLlD2zX3sEb4r4DiUkwEPToKNsb2yc6qCIHlTUshszmeVl6XHayBju20B5E
KfzADi1vB+GPh3SqNO29GAXm0+RCCkAAjm2AxXrO7rezEAOF9M9PdscR4qiA
7mIv3FiEjQ2+YNFtYNrdFubMKWGNElQn/mepCrKeRrr8BPWf8dGySJt22iZu
zKQudNJewaWO0Hzln1TdCDM5hvngjZQJIgePjft5MWDerTQS9nrfKD1QMtYk
7DlQe37EIbSXtKIrLL92UGL8zsbhYnEgweKsWu0HkvDWdeln7ZYbKrlCBX6I
gdwQP94m7Uub10p4X/r4zXsRFwNdNK8fxou+d8rbWLdkXf8hsx7MY/nMrC7f
0FbjJeH28g0JLKA1rXqRnHRpQ9u3qP/bKIsLLDl5BHMyePeh0rUD6TBNi/fy
gd07hveG5gz3nlSCRaZ6E9m7yMM4czBIwJIprEpjRYx0q6y0ag550KdQDGzo
0GOODB37ecdd7BJVQkjeq0ZJlaUPmYeneRqXJLlI6EfXr0gNJr4zPNxhlqlm
kfNJ+38dHHeobkWYg+RR/bColgtobL28CO2FJdKjfTMBx7JzvGQZ3CWx2aem
8UaZpBaEov4M0iAVPC+0mV3+zW2R1P/5LHc5fw7jESUEloCRFjFPVLbub9H5
jWtaKWBCpTbxA/osKBEeNP3VJDzGY2qcU+4whYrkiT83+Z3RBcCHJrNpHQHH
GkbWj3x+ItueYHCk+nFe8laG3pdF4h8TB2fD1lzUK5isl3FPjmbYbP0wGAeV
3SN5LkrsUogupzJEl4vxkhX3+4h0wlO7uBkTyPvMfE6lWjXXEiE9pkS7n3tK
DLM32bT5uZ8gqisMmyAXdVNwT6WUj261+B20ya7pUP57KqaTau9SyZ/XKjDH
ideTDIfX9VJ2AhsrafNcUhUeBGYjRW/VMdE6rm8NKXKvhPb1klwTh6aMFkHO
K7E1hg5hIdURLFWFADXhjj8UhRdRvk3TJNlrmP7DqLDZCl9sdSkXqAdd4spJ
X4cYjVr4jiIJGBT4ROU/8EafCmPNL+N6w2myFUhQ32NybVZgBrCEvsYIUZ3K
LXAO+1xYIPqvhXgpTmqn3L4StsdeM3wdzVGaCpEmmDLyZDfTKZASOBymwX4w
HXlznXzI9N4SuuzF9A1qezb16ko4iO48FYH5384lZtVbIft0PUGrHYsTo03c
wTYVo+IZRgKqit5yYgYtAqMjHgGpr9KXZs73w5JwwqVn1GnDO3vwvPRg0+cu
zigxbaX2+s62gzNzdUdxSKxpBtAhPorRZ5ur9BXa0tU3owAvYQqNFuSBj/hk
4qjHCqBYohIAfzXKzUhctVW7+vv+brwHqu2QyxlEgQCzka8ew0s67tW4U0iH
2Fpdn+UEBcAlj7id13fdG9IbBXkTDXb1avW1wWwEhDqzuE/oBIXtJF7a7dsm
BcCCVZ5AG85Ic5Bj7IomZg55J6P6+ahdjLnHUt+KTTcdgwvf2fqFl18AKhIk
b3irY7verlEgcOuQmlZ3OMwf+CBWoijE84JyCGBZq0n7bQNuST1h97OOX/Lt
7mOd+C5z9uEgiwOuOYYbXX2ELHULqUksIh8x7w6/Ouy1zkQ41efMdeCiYiU8
L6UjkQf4ffjqD3itUpqb8bOVfq5IovUAOz7kspCo5JX+QWTsY9cP+jZkls3A
NdLDBRJJQjAZQcIG4rq7shnxrKem/PT9z3l1X8oEwnYAbS2Yik0pBq+Mytmd
h9ZG6C7S1F6AEVa8Q9HXdOi8D1D98S5FIAmDnCIRIFGImJpTbxvO5mOLDzbT
Iq3l5OobiEJK5mCo2VCiU56qn2FbsJPrtWHYyfhtHFICYWaHrwr+iY6gk2L8
/AG0SjmlYDV0I00PGdSdlvwN9IpT3Q8e+T9zAHQr2aSi+lSGjEtZEEme21FE
LEAUgwzXeQsmG9xDLGpa4dPFcsIuJGABDfi0hgFoIRpvH39EXgknWYw2Ks0T
pO8hLuMN28NXy7epfDNUp9pF1pWQAs4Se8ECXwHVwn784kgZU6ZkOa2x3+K3
9VCQTHhP291HNzyE9y071geE3ewYiiO6DqlhWkSM9+edVB5EQ9ahmLL7TKtc
e9ZSlvRW504H0s4FS7w2uTD0ZDnGkT/tTp/tB7oESfzAXM63b2aHCW/oieDL
fx5jImxa7pmGCGpUtQBIln4517Yw+3GM5tfTQP8WBuyStXDtJtK6D4fKhHGc
BqUwwwpkpQ3gVHc76CrF3PLZHOa9QzJJoLiDqcfKSaJhcy+DGxY3eiSd1MQu
vu2xKgGQx0gUT5QtMam4eAamObgyKuYXee/fm8+NOUKpJMaMq7rSwO9kY7Hm
cGD/Awy3yLVEWvy4m2pdSVkSltbqq6Rw1Wi3tSfkZ6xEbbKvUYwD1xyS28Or
PW5LJzpm/0l7WqUqB8bYuo6pUYK+lxnXJy52HZ32qGT9jrqv/rwKV38CD6/5
RU7gZhutDfgs5rBsRyRUhMAefLPaSSrBmqfC2x7yqPlKJas0bDaLEzYlm1Xw
mymCGQsiTYIqRrTrbDsZfv8C7MoOJ4mW5ut5SL6H0WT2apfoyNlGAbdaNFuB
+Iw4TMYt70SNlRmzmKSlTxmJpXlY/yx5rBpHhWEyjp4Gxv8NjEZsMIwG2Jx4
M5XBzfwNYDh1v6ClgJEzXHKqDkJGiD07skOOJKwDdAJA3UvnIH96Zf20kBIF
9icFdNOXMG1jQDF4lxQhQGfHsi8sbptRiDxOsgwGeloWHjIZ6XWP10TvxEij
qXOhUdANT3OiuJB6SColjwAUe3cQpJ68h+X+g3Gk+nxPPni/cgXje65mMhmc
3E1vjHaG26W86484EtlvAu6xhJBubHougTvt3sN6ZyeUqEjEuyI0H34NHYWp
wt6EMX2kFrbuMIUpWEAWwOgq7ZxTP/RtE3EiZ87qh9S+e/mDaDEgQjdHIv2U
YjOHX8Okv/9foGQBESz1RCEl5AszEjzyjvEH+IpfjkRKaLmNGu+21MHZ7EIP
cAyzZrbY7C6y2ZSYT09EMKVIJXLd8jq2c0PzQmCsW/c2b/1rYXIUTz2Oe9M5
Fme3czRY4bHeBzlA6Tkdf6Ieb56zzKhmUc4pdbD2gY+9p8YHJHDmAfbP7bcX
DfEGBjhn+pTy4eNvnAZJsrnstPjWAsZLus/UROMIA6HBvP3jXceUYe47uKHM
rPHcdCjIRgiKhi2ApIVKefqZOysCA64aBVu+SbjqTKXu0uqxe62TlZI5gDkV
xh5wAX7D+XwumuMDkEptIfejfBLvp8CNAFR4dVoBYySnpREXyxMdyHtETo4W
Qq6kR8hhTnJ5oe6gUfYstgnQfOs3Gk8Gh9VHplq/0FS7ebwb9dttlWlUoYqz
qesTQ1m12TDNE/9plD2SrV/HUcXOjfNM52ZtEhR5x9el6OC4Yt5T7qIEfq+w
7CuETWSrSq4vcYagqJpofQuTohhY6sZAa4f3aWpKY0TglpMu9SwOR+GXWMpA
3aDE/0Qw3wZgAB+Q9Ja70BMIQUT8MAVStYJ8yG27UbVxL69rL/rss1jPi5qQ
qvnlN+KAAazxKabeJNH0VvaKR/eE2PcLBC2wT4/sUns3aLTKsZ0TasIUFmcA
sseStC6TmeIS83wLaI/UzczCRYIQDhYUasbDXOPjqvh9tVEpYVO4leVJublO
NUBT/vV1VaM9syJoxAQ1o2x8X//RBgdgwb1K58Mwp8sllO3J/yPPMEtVZh1+
+h797y2E1ZrFa0jMNqHTsFu7dkdzRSfdVlUG/UDNRCbaslTjZcTSWj23MqR6
SyM8W+78kYJ7EEFbjXs8+vXxT7GYJtT35F4axxBOW33eX9rT/s9kzerlbWXY
wU4Tre0hc6GtKbSQLrWXHqU7q6zI8IF7u4O/yhNJFUwwX3lhaBc573AiIlXO
c66y7Xm6wNxVrxi6hTZrleknY7z5cElIegFIQU5FWv18VpFjiTUhUIyURSiG
18K23MgJewHGv6+xp/d+W3IreAbTzLMmOZ2T/s1ogeUpGi62S1GfpZ5ISeSJ
r1uuLy5kERMpUzhk1icuthj3C8GAfQycZtQVBMcFtZrQSKPj3B0G/TxpcuF5
ukltCEh6DTdIFfpbfQKI0ds9FK9XHlT0iCWlx+VdrGzrzJcS8cTBShEkhNqR
tDRqvYYV4Ovwkp3/oHl9HdrxaY7KlF7FaLZIgRkX5Ebbg+wgIxp1Nb+CgPV7
5kcG0krhMJqhw7ODcW05qIlLCxyASDW7z+2HzIhrlVNRcr4i6SMu9mke/X+W
KQ94apRELAyO8CyX/2kqFI4mk9kHDW3f4qinbZhu5uq6WWRMhIgRceZXuur1
N4kFDvEkyXCnomc9bFVqdRhPqKK+cFWyssN1+5Q8krNboGwOaxaNGXcK6bf9
ZEC3hQjX6z5ZolprVhvcrG0ny72t6pl0A2QQ7IZVFEcH7CFrXBXzgag9G+BU
p9IwENArZ+4EjPTYGcPVBwglPO6wS7SQJwwGD3u4PFLJvv62DcVejT+JVozW
JGsFZV2WFyQooLh9BiGLsAMGDjHiaQc1b5oWIkUc21wF37n85E7xtJi76FA+
dBEN5osk8GH2FDMMhdEG9h6HccyPMualZf3TO2NADH6Eiz1NhhgGmxb1QqY/
gikfCUUKiznTNBf83/0LlftanbD+lQUTqidIrzukGumPN4sW62lXfaqeIYlr
nuddob8LhjSIKtMQ7olc4UzZHa/KYmCcOoyUDpW86PPTw4SZ/RrrEum5OR2B
/8MDPfMAlzC1brZZKRkAdbrnAUO9lXT16uv/qnBB0NdKTr6zD04NNtgmg88v
/DD+XlEN7DOG1WDVzZEBEs1DMyD2L21NAnU3H0XaxtbYga26K+Xbm2oQ8/pC
7YYsD0/IFG4ZWb5OovNXqR04sh3dERitn85w+LEAvS9qIT0gAyV0cCLBJasu
7FD+4h6O4XLuFNI/xQDJnLpDazRlTEAmdZcFyIjYI/szTU1dkVTes+PRbJs/
G8QAbVYnYaJmBLXi/4aIEgUnyfwE6kLOmz+5ZgCcu97J94k3f3+RW0BTU9ZP
j8mFhSsGVp07nNrMTBlLIouZJgLcvggYk0GoMhQuuNSV6NHGnvQpxU4xDodN
9cUv26N+PHdmxXs8jz5VWmquP+pXGgDkei2flDDMc0553NsDnqc0kOKgHYUN
mpO21U+pOhAZZqHEaQi7GHfVouEWzueaxuhq9nIEIGBsIvRDUosJ6MCQ/PHf
Qk9O6bCjzAETlzocfYZpQJ8TLbySZo3LtH6YqQo/NiCEHPl3jhiZXclCOAmU
w3n8eE3cQFKk+CGQa7WI4lLfMXYQoU7mg1ad9Cny9YM1m0MBYzxzw7hHXtzG
ssuM7CG6bm27YVWSIk8QgPX0PxEtXtguf0BK32E6de7u/lchrqHB/ufGwkj6
8uPnjki5eZIo+D0cBh2tUPml9hYGhW4rkYRWM9Y6bq3NHKyaj8CjZRSzsUv0
k5RiITyZE//ySdJy1F+2qTnpJFytj9zQ7aSagUhAxrDNlnYF0Wp8Qs28WgG4
7Ir0QHt8b46Vc4pihb3nAteL6pctK/CXpp65k3Vpjqh/jQFl2QGSAKhhPzRi
y0j6jwzceaU0lVYEYMPYljbAwPPnnDbJJsyK7ILDrXZB5OXORgCmh8p21rlm
M7owLViOcy9ZOaX/kzgUZ8H1W/7uMr6Vg9WObjkZHvOrpcP39fkxMg2ye2UO
FeSXYY73lTf6ILrzQdVblH8nFffmdtCmzo1/2W5clfHr/QzPK76asGpdsb6s
l1iByi8kBOYTbJkLq7RiIY1cWsCSXWQCtJQ82kqeTckhF4RbanvpdJoJvxi9
deM4xBOStUrnYQNpT4VP7tbHMU8pSedJCbN9Etvq1/73xug7K9hRuId6Jgvk
YWL9dsRS/J7dAM7WXxVT16lNkDwk600J1RpjdlOlj9DqwYgwz+23gDc64no3
p0H9PF+TBAAyfx6EgXPaRZjBTds+8/2S1YGA8aP7Kz/DyCU3jrMWgAkEYyJ8
aTO5gMBLqGSRv8HHCFlLhyC/afSfctLZb7G7MLFnOW1a+qrJyzvryGfmZYRX
8VSvVGGMfji/AnI1p7kRJMb5nRujzW609lmlXdL/pK7YfxHL83PfMVC+Xjf7
z4O3lkl+OGclDGlhkCYuvK8zlq/rEYvIO4zL2NiEMIGcGzeEALa7MjU8epoD
trMNiKJzyn0XpKh62NmgAZiL4Pkyc4MwMFe0v5pqhe2MYpoTmeWiWM4AmXHm
LnWg9KVFb+Jy4ti/40sK1409A0zmvrzqKsKEcsJtQDpqCze2sp0vX88CXMr5
gG1ZhYZYCDloFtW31tPVcycJogzsKnKoGGPXDo3NvBXesbGRascJpHqVdsAF
e+ah0jmskdP/+ZNlpB9T6x0sP43sR9+kVd7IU810rPTLTnUoXcnUdN8dVJc4
4hbx2/GTMuwSJ66kKIKzRjTXJfV+5zGxR2tZXXLMUjHhuYKE5CJCEBhWyWqS
+v0UhZ4dHYHX/Le3si2b/cPoudLAkIbGcX53v3YD3h72H2A1AbqOwtqnIh3M
gBlGbc4Hk1RCE8uRRMBsr7ZuiT7ot1qj9uVHOS7kpz6PvjXqWO/30KaRNL1+
GqNHX7M3h4jFp7Ga0pzul2bid6nNUSyX/xtJB7rxbEPZKSsmVFd3IX8FN2PB
Ul5iqielk15NN+aUtuY7Ntfh9FIAgi1BV4sorteEYLwnzjNGPhjNjFlaI9In
+DI9wdvrJBBmsBq1Je9wysAoDocw6f6d1KzFMGiROJy4v3PGQx0zsRwOcWQP
65YWksCVnpZIP939BT+zm8MwN5PnhtvV/9w99mRBBYpVxA4CVFwZn0r48OwI
nOxKyxDNxb2Jqi8qhTX33l3dZQLOZ5j9zdNpmaJpsQzjhNwYd5o1TPbufc+X
cSfeuwyEHY0MX2taNBJooy2zhim48hT7yVqAmX00HxpFnQFlGcxNtNiUv+Kz
SHXJyNM13ZYSPnlEfzYmmS2eb1kJ6MhJ7Ttik7yMNFdpMYf/PX58GCJyFAYh
DMBfA0D8slQLWwDWPrPS96l86Vsgrtek5svLx/0oKtgy1XjlF4uinaFu2OMd
xBqVs0i2+9ZH3l85HlJ5fx5oGJ3OWJCxGckbfNFfwi/kkp8XN1oP97BVppYR
EWzJKaQcMWab8ZH9Zt1xatebhegp6g2FwgjW+t7B1ViqK3Q0d5jzEJrKxQDj
hQGSTe6qTHQfJBtVGBSO5oL4EfTHLl+XE3TQ05cxNAoSlm/KDBRAU67zKf/3
YKUxi4Dd5DN0ZTvjNeqml8spBB+6nESBvK/hvjYSztZ+QWqtF7+Ck3NA0jdn
3B30KvjmyTEbVmJgu3cEa80DFemuiztB3JMviPJx8jTIKNtd01o5ncUMHoi4
V6Q20ifaUMYPaa7cBQHaaVRjorXfpfUlxSdZW2kVYX6GNCKToHiQOIuLSqb8
+CwKEfLgH6p+tI7L0JDgJtbJr2KcbkyUfEPYfeSdGdPkvI9G831Q7tgSH7qW
0yunVeGFG/UVhEDex4nNQwtORaatPrEM7gEWkRrfP5hQYECiSeR68OI6Htlo
K5o/hTkSDyTqCemoVOwcupNwgXYcKqpdTs3jNh/YHN8P1f8K+ZXutJ501UFc
OMgzkUn0aopquGXPgWTRiiEuR3yU9/S2qLdpXGvL7xI9QSGq4D6eGXHs4OlA
vVkpq4inT6gtr+4tklSPgOEK5Oyw2aIiWeQfaHh5RqFYY4qvXKr1oGYFAUxb
YEncDf27WwdOussXmzf+QEXylEHPPIEWBmI/7zFlByBupZDcrboONnOokMlq
weWmlldAXw13R00/+HbhzbMUvVtDevORDymtZEiSVgElKyeo3FhE6HLnxEMu
qgQP+GLy3ksQfNN4oT4n3H6msbpAQGH7HYJAmtTBeuXTIkqwOidYqFi5u8eF
Z0sWI3SFEm0ndstInhGjJ0rGtUoEMimwfuWyJ+2SEgoQlvgJJmfIKJmChUz9
/puOjqCSJuyC4y+nVnde1PXHF0UHNC1zT4dcThpGNn5HTytZrGoeCKCBgoMY
SVpt5s0bVyuTwv/jpEqMzNls3+pivOMQyomewt2CGHCYxkQ9RMFC9SiOK4TI
GXwE/YYiBNovc2VdQ1KSULXqdS2rbXJC6kyGAmMKofOelnWcI+1nPOleb9w9
ZLeTKv6kjVNCdYeT5SNJ3zR70LPxY+X0gNf5No3Lj1tXlZZ+j7c8tIhsYsl6
zJ++9Q+KmLnBAnpxu21bOpCNpva4giVfFnDiOyJ9sFP+dnNElVvn4cAVOSkB
/Qsswx6c5xBKHkKbjI4HkNWVYXCFGY6lHBbLt2zJyR8G+E9WyBNcpKIxGpwh
gc2quTXAMY/CyzBpZMvQzHnZcShNswltPK9YhCuAwUv7cTyibX+D2340uOKF
T+Ia6EgHndRrveE0jeXHQ8GqUU/S06NSmvdFR7pUGUD466REnCe4vuRHs4Rp
/NaLs6HIRK1tywlJeIdTWOXN5J7beJazvclf1oh9K3pTFc1+XxwTm7MX5Rt8
tHIqJuqN6jVFKgjx7CclHIgrFAwwQm0cvZLDBqjsaXxvwt93wSYfhN/2wW2s
kxVVFVmz3nmziL7OFF5qTYZe6ZlBOMVJNOYgCikwlN60sRhfJt91aXn3VdBm
LqxLvoViR6h5iaW2w8JvfxI10XMeamgcFOCKgTvH24KKPv9hjMQBaxCoIwaF
3rJ8nuywGQN1gvhGf+Hvg1vpgRAXgLqQZ65/QhR3dXqRAUhPL+HJtWtu6i95
IOAhmmaNFLVEE/cq776Vgt/130mC1caVAYG+iZGvlFEMcIMZLx9A1NP0VafA
68Bj1vHX4N0q7buiNR44Zi1JlpXMZ2b69EEZPFJV2xkKkLDlhZj5r/s9nQwN
qzmgIBwI0G1HeK6TMAOGF2d5NKYPOSpLWR7t+xqNn8lv1j4IU+D4qDKYhsb6
H7GWEBHDNKwkE7bJocbTPgbHB+yIV5GsmS/rpRLyci4HRhKLv2oFnbqfyMki
UtC9SQZ8HDli5975P40/QD+4fvn+kMs/U6V0Or+1Mp9TYHhPjkDOlxbQMiue
NIoEu9eVSlReORiJTS+hrkDwDRU6qSEtlj9Cx8dllrQS6ynQ1uZ63O1gblYc
j7rYTdpE9OsERvavc0kWz5HlZkya1rnFXeSaZ4Op+sBL4UIRuDLoh+UNLpz6
kzA6H1vyVIXCXOdTtMaWAm0JHzt48I4r3qsz4sNtEhnNrLqxG+xiya78vXVs
ZUEP+tbzql1rCWfETpYxVz/Rz/czg9Za400sE7yoID8ocNZfKegQ6JDcVYdr
1tvT6aH4ajat/PROV6tcKxi/6StgSH3kHefgIJaFkviyzgE6lLAeMt8rNwWZ
lzvcDV+rsX0OYgLCnG7dYxI5AF8okvpUzYh7TM2CALRuHTbldGBZeCs0YKLN
g2/vMezEZeRqDXqdLfo0GCv8B22/dqfUS0pOYic1kiGM4dWyDzRNBHHDw50B
RDNBHOCm5xywsPmfFZWvxFIB/gPA0egESNrzjXdpRiErCf7hMXwtENQRRgfh
zvyr2CAYxbsSrUDH/UM7KkB6OjCZ0+SChQrBfitKIRJJn/HLktOZqHAvU/uJ
5LKK4U0CPoWP5HWl/MpY3vT2RsBRGsRsBUxCoW3T3yV+Uiyr7OmlE/VHfBbW
YM0B+G+F17m+Wy0ZzyCO08I5GN4H61FLyB4Bx1cbwH81kNg9HEi1kSFTvdV9
5OsucrMJ4L3LLKzeI8+IrprdDY/ruE9QZVx2scM8pLTApG8z326S0RwVwxJa
7Toz1pIYr0tyAfuKbJ/MLvbOrF1nui//RyGvqJovI+vobdFijPxFLMO6JLpP
SAXggTEpexENde09MzmPTlYxYitwnAkuU8IS9QDVbBcB+4xOzMcdQOTeR3V9
Sas6oKXgomHQIKy2XBzGEJWiQIGF2uWsuvNv9GMtR+1uLfvERKuk/a/blrUK
XOHwqdMJBcA9yvRfgawbPR14YAqzWPXrSrEeYZaMBBuwP81Z2MfJhJ5jsOCP
pYFuzhseD24zWpZLCe0unbTLGMZv8Y1s6NnF8b911m7SlyTMU3lz+GqwOkny
VNnfi7R/5ZXgcCqHXKtj+UbmOQlsnHt5uRgfl+0axXg8+1mYSfFYA5LlgoDE
WssKiTXaUxUpjdJI6pruMQBr/5e8v/9QG+vSxFgGBhwUQxPrOZHJr7o/NR7G
hF2hxgDvBJrl3qBVq2Ks2rBxsGtiOTQiG4r5g+6emGAC8olKIRSl9gnkjzk6
ZzBE3xbCMsapplCa83dOdP9IjeVmCUomUOcloqrr97UnycV8r5GUZ6+djw/u
QhZU3zxt73GwbGFqF444fuoSdJGythBqwSg2104/h+ZOFlJfAfc0VnB4hcit
CUzA2wqXQKEWRqiSqI7+9S8M7rHKoKqssg6T1XpKxViVbyWv1LTx6t4Owadv
52Ci+Alt34/B5gJvohhrFXK9uhtDVyc0ny/G8WMcfGkugdOBfNgalYOWTgIx
ACMehB47pNYGVF8kcOpVW36eY+L0yNjNJnUik1w0bjk3mEHiJUQLDSwAs39G
QFcbvL5/EjxKt1nTb2e9URZADIBc82/KRSagr24L6twLjUH4nb6s/ieP67I3
xm4PMnP16jz8AMURyvCMFIdXTvCGlxD6H8f0+rMyqbEEW1+1D7CwW3icxDu6
o+PK4GK/W5/kxhfTfPtMtJfI+FijTxdxXhNIQeDNjf5d+61kEMk6HIZ9p9XY
vIP4keH1qsfgJc8/EpWpGVRQzH2LLJ4q9ascLmHVELNbk6ch4uZKBUqqgv4f
/Za1/fTNoTmCjNckwEQdP51QjSQAudn5RszehVr2Y1CvYQidEDurwkGVh+t5
OgQGjQgHPvG/Bed8Qh/s5rDVCLzlvcR/E6d7v6s1R2fekbNUW+FTXY7yM9ea
t7NFSveHRcXi5vw2UQ8nVvbwMRgXFFdIOmPKM8iPImElLSfgqGgwlPYTYsI8
eYF56x+Ax8wWHYDTgFs2Z+upUr+kSHPjGIEGNW/S/Xs7WROMQBrgvTtStWMB
KIOB0LfC7g1TfMrlraQSTjLzMHZxFgeZt4YaUu/9KjWfHB+dxzBJA/oipw7z
4xWp8JZmrB8cz7yzh8anvtux8qcmA1rVqLsaIdUvGcrP2SHfFcmpfobnfiKQ
2vkXoxcs2qbcQfam/AY1DXyWWnbiyRHzHJQqbXf1hp+aVSwdXwH9htDG3/Tu
0ysMHX+UP53U++UZrlHzItKA8Bt3ZuRTlrSHqXj6CiB6V0pr6O4vFWRkCRjp
v9AnSBcN6mqSeSEn7K2BNVUBSniWvnfhjB42faYNZkDFTI/rH6T5HnXO+Dyf
U04jB9++1GVrs8n/f55AVO9CdhYb2151nG8UKOT3VpYTqkbQV9rjQbl0vFnT
hOl0Sej8bkHV1CCxVhv6NJPWah0Kvc7WYjoUV2iS0uYm1R0gSdw5wUKjAs+m
vGOdcBfG7AQJPBz6Cl1GO5m1lpPyzXm1gyU25Ymv97ugo+OaAZWA4jBeRXVz
E48NgyombAJ22uR0v0nKrX/OqvTqqip0cwTCNg7tQPG367V1c+GNwuv30xGw
Ctz4c4YIuh8mydbaynjiO3UwK5T2kcX2DA116s0GM5BVFjd+FHIWoW9/1q4y
8eP/+Pja2vrYJuCNhc3JP8Ahnw2Wnz8r4c31WBp02TKmOLT+I6udGvivZNJG
RaYbDFWtuXfAAcxh+5FHlVhP19aLCtEPJH4UXJBwXbG0m26XZSqXD1lOJfWy
22b1UCmgeTnIdHCon8/0woV3g7jlcp+wmDFPh0OVFDuAJlp7jZSJMkf80GiD
F367fo2teKshpw9XtBmwWpoaVseQZ9od1J5gYTEgoemFSsmU9zgahurTOhkl
N9855TPQy27SMtQV3ifJewoSXefQVu3PQ/+ZJyS1KaJtE4UeMJGckPraX72W
sCs+SCE/I/EQDBieKDQ8+OHeoMMqB7k9CgX5f3HlrsrEVm9EiknJ05vyCfjF
bpMKgE3bX/1bQQZ60CCQH2rrYvTDTl/DtCD1PFAe+9s/1uxs5DTKMpcTlMSP
pHbUBmGi5OOYlAq9YutOTMMMBzZ3JE+bf4f3fAi+rqqYLZSP3SyTO8lKECN6
F1AHjqcVTmK7YKaCH+FoHoBKCc/J6zoDuqyv0+zteNrX+L17d0idOhZIoX5w
r3FFs2bZgLYXk/UsKQB4sIdYDHDOZ63/Uh70zfvda/0pTmfkPLdR1BQgioYn
mR0bQ0rZu98PB01GMlSYNrDAT8rS6z3AIWHBSJom46JmhtVtJ89BuTqX3waU
CkkqlfZc+ciaJk2xSaaN75dyT8008gL6G1mffJ7rSX1gGvvcfJeBrgUm/NkU
cXrlkHpP7aL6JllLCY9iAVpmSGAPb2SmNJ5T7DZ5I8l3ZlsrKNlUz/wpgMH0
YmX0MuCexpl4e/9gSZ2oqf3jXYnPpeAgH2XPmWz4/QBPoiZz0qEvuWfh547m
UHptB0K4+R3dnOOCQsDFe1dsgWxAyWTRpnjb5sNqE4ydn2DV60EcYdKFqNZG
J63c7j8/aXZBqCI1ioPlR17mRoQvLom6V7flm5vnulaNszqNPuKSW3DdQowm
+GCFJTR/r6vP90ngbjpLLImC64ZdcDUnHnFprTlTwnZGvt08sJo+ItgWqv02
mV3vHg8OHVKCAsp8Zc1G7PLjyygomUK512fQfCdtzbwWVzXitKMIvF/WRrAG
rUNm/TYyZ9OuTqjD2q4N59AMfqr9YQDHaAFTfvSZOkv3pb85vABwBqGDu1Xq
0mKXSWtceZtafdOJzDISc35l2SuptRuWKhuxFN7kP4vdnAqR6Y9uYPXFQRV9
eHW3kKISfYAKeSbjiOQv0TyYY6SDazlst5LToXZY3ypkHO43LOnQpY9aKw1S
gKLRI/daYh8sEMxXsJBb00TDawvW2Z9o/iVh3ExyWqC4NgHHuFi2XfAl4v+y
0Nw5g2OVxi7x55CgHRKLiuQ6Qvu0+FJqQv5Xlt3jeSQlJEF43l8/2hmEL+46
dn/k9puCj+GZLGjukJ1yWnA7xWdjhRjxZWzCk1OIiho12Mt16kreEY/2I4k4
4oOYGpP9aEzTehlxEeONYRPpXlZTVJyEOf3r9Z2Z9CGVB1g78U+u6zblqkvZ
1W/WcUQUVCZAQtMmYM3hsilUiGSBlf3ZDOt8xm6kJbG1nW0HiaBnhb4WzxEa
PBJVi3St+SzyHOSYLbtcCnHf1UECiQMuyPbdL8XpnQfE7OEXoGEkjU/0wCoF
0gEZQyeHfcSq2QDK5N9PCVpxXKDWgPwPEWgY/nUaSu6q1+rlxsYXSOH355l6
yBIFoPrWifF/9FHayNEVGkZVA1mxbrwayQfScIZ/cA4vQvgD8CpXOJc/6udY
lRjrn5+679y1i0hmPsbio5fSrLqG/oEaAxNz2FPNMT4RcHH82C4Pc0aUjDIe
2XIRp8pVHHqmvcoU4GrFllh0OK2kgztYagm+2gfUPc06hGpEwNpGXK3ALpOK
QgRHsyPtPUZkSUI61tSLOwgONe9jXgXsKhkv7V+RwZGG0rRs2WGTzuU/Aa4I
P9P5TiydlI3DKOIGUyTqYO34GattcOZeQ0siQRHoJLuLs4ocfwEyhTYPCtQK
oHV3Q5ZPt6Et+vaTDlS7ZFhTl0iaXXwd0iUZ/ITI7xJ2nFAZBsJmMZNcYZCG
5CDZcpe4Q2wvnP4mLUreJqgZyzZze0rYjAOZYYxyHHKgjRnVXKOVYZ2lLUht
IyREEm+VHat+sX9LCqeg0L+impWSWbVpD/8WlPGfnRa1TTv63216amzNmzUA
36FNkJ/VJqlp3YKzr3mG3mwbilXdPGTyXwh7Bn/mW3c/qRFdElG/vrpBj03a
9yv7u8/ElynE6DW8smCHNUiZ+iAO/b7J8rTRWsBjgYJxgi7BCn2e/IX0Ww7i
9s+ZRpMwji4SmbONo3RUwBPw+2FNftnbytNdEJg3Iy672EerYO05Q5WRFU3p
d5BeuuOncLRu/xAjlkEdJzvK6ugIYlcUbmA3XPFwSasSvjojQAjQU4xbzjNu
xlc+cC4BXBJURloSJErnEuN18PRO9Fb0GhEtipujndW239JYXoSkOKpzbuR9
ccq1/tzO9MGPthBfNNB/mv3VG2McrgPcbNtAlc3MRH/2mJ+WR2cQCMv/YVDf
wNv7MtpE1q5od6FHqujIehJlajkyz5YFIhb/hmoakdxYfydLRu8mXF2XIpAe
i3swDhbdSigl+oq0KyMroMXGziqKXOHS4mLgA5cDn8VKGcyEfePKd3JAPR62
IqUuIqKSZxkyeEjEIeuK256Kvf5T5msJL374A6Q14ofZTZQcoLHGrxsRkF92
QhMjSBVGjDVYlvBfBuYm5wZfHsYnK4bpygsRaYYRi+N/RXBOI/TRJ/UUqK+3
DMhO95ECPfQ9EAeJCwMVERUhgIHaKXGo9RHun2eNXINavJBKUWQVlOkP+pbj
tlXYaFA4D1b20h/3n9oSzKntmcNZWxJiMpSN7pATOz4ZvGdC1ZwFd4Awi8PR
jvdcua6b2CTqERRl2HE001H2+Qelbk2gJ4mMyaUe2d8tHkrntctB17pf7ukU
O46U6nTTfRBYhb7qfrKouqkLPR/hXu5FLAnl9eaRTrep9gDxdvJH7ufRnUYI
TaOvXQdR3Q==

`pragma protect end_protected
