// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Oamo4bEVjI9EbNgBxQG6V5f0FjcFgaUnXpn7ZE/2yt0SWCSFx1NWA6ZzcIXUSyzn
/afBjZDzIa+8s0WZN0bumL5m2a6fqX+ACQOhzDFAbk1D7I6VVoC3VNTpB0XMCJBK
OZsmJEC3br1rjD5kZrXTkhTBiCemmjPcou3OdA3H1Ufi8jV7/h524g==
//pragma protect end_key_block
//pragma protect digest_block
P/BIPZj0A5AMe/GC/2t5l6UW5sI=
//pragma protect end_digest_block
//pragma protect data_block
6rMy29hGDZnXMzbZ6FIXoLPC3k9GzdpeCqg8oTMfRmXZ9QSwcLKOIGqh4G4jyoED
4tUx5GiV17Szvgj3juwtKa2DPwbXtkiBZuhVdBs/+LvXWiItxGqzrb3NoWcZQH/U
Dvj4ykKU5Yfq8tz1XDfHcFv6LrFkXVpoWnwHRMZzJqoUvJVPL9mYCgHOC5r4Sj0z
V2n+GPdM5uhLUKyPXdL8/Jo+V9YtsIB/DisqeTiDEsYqBSQLr4mkkwdFiXOAGqQT
y356+ZyPCjoJXS6a100vy4cHKg+QVKl9IpaZPXIjbmmmfuCjSu5UxWJw2R2kK/g+
2QAuWME2so8KcxyzZJmTrKZ+OfznIOY5Njxa/f7JQyEodrL1WXBCaH081sSAkriA
3epqLoPMxHWHjDcmlYyLPQvgXxedtWJ+QFfNo2zoAhoNOYVktitwvDu/loN5PSqV
Sq9WkCeneOMRRrF0BsVNrduAPXvG7S1ITIjP36NA3iekYcaPkdNFLYPisEhJXpg2
Go6Hpk9+Tn69Rjvx1pIqPgC78olVGKwmGeuEaZvYIgY1PZbrHIJ0105jmpb2lDZ8
5tbi9oD3k/OdXeF1+9gWqVLpRDLFl2+OcLJJ7X4vCJx3BNgMhPCpK1ppPad7Yj6Y
I0MBPBkEQM4ZS430iBvJKylujGB4WEQqSMSBZDG2NXesasJ7kEtATLHa60e1UWqM
S4FAt7onU+fES2FKpc4OEUOMkg71hpPUQE0qZRMS0J4rX9CesXgHda+p1Sno0oiT
IuiHDE8+NuGgySWVz7ZMJgXg0Zih5oDexi5hAdyZrniJLy/cUzjyPfeCrUwuWs5b
vq/ZCz5p4QpG4KZJVzbrwo+DstCHmZIxcpJ2ZQ5mzVDQu5ctEh303mSUVOAsQnwM
UD+oYAtOTqBTOiPXqs/S5e2ysw28Nr3TaOp/vPxY1dW9GUE7hbQAEWOr1eKs+0D4
qIHInNAv80v9aAY+zYLoEWfd8xckYDLp1pqjPdag3WNrIpMwQNSme9Sn3++a6H3D
yInTVPnFNgeqTsccKPR0n0HVN2OG9PxVXAcafjpd9aW3CgvlZmSS8CGzu4YU5Rtm
ZS5unxK/grcP4K8jp1IuqXMJ2D3a0qsWEg5ER+TCuR6fLRO6u6g4B9Y5BelvCB/L
BehC6FQpZyImHdWPC8hYS6K31hJdRWauONBZ/Ubv4Yvmy3usBoPiBvXggN0VK9JI
SVa+z73UBzrMVtXtLhPtmMVYR8dFZTj34RbJTRDBRdO0XrTFX7hIxzZpLKwupo/W
LiP1HSJU/+bEp79QwY+BZhCHa2BETPbMK+hL61q2pn+/Nx+PONYKMryDChYFyP2X
go5qu8KWX+upiVPy9zdascbj0I45OGB3UX/lH6DJtX6AI12QXOgq+pkfuGeUdsYQ
1MHQK3raf2nOXSEx3NXVDBzmplhA3nmnjMsYSE/lks8EEGD9i6XJ8C03CFz4+2jn
RuEnIl/ZOCysdJfX8Q7NEdyfrpHCOEFh0MO28wv4VWNUZf/PhNP4fIqM25QsgM6C
RYBbM1xiH4yFgJp8nelDbVc2OvI3unzWnBtJ0wGGcUFIC8k5VPOW+ZY/C/9d73MO
XTtcI0u9EvG/h9uaiqQUOvTnCVxHrzt1KBsedcDpzVYJZTqYlpcFMfYWE+hVzyUL
Zctq0rsFF+1MLigJ7GYw/bUjx9byb4WMRdElk0zYlgOkk5O6MM6QkrtRnwaCKDDG
ltL9zFCuCE5SRUwxs7gRyE35OjSzK8L5sOjauQR5Wa7jt11KrPIsVVL5CoyzTbIW
MRa+ymNeug4HSyzuSP2Dhi6nbRf6AdPZ+8YrZ59fxU0P/+Ex5OFzbLhuqtTTaBG/
0BTxMsCItRFyXNLy7aPjeRCbXfX3tnmgFOzmHkLksgI5xlpoiL/e1I/cv7y8/Xu2
bMOUTc9pf3fW5lXbknALkVhV8lzp5+lE02IeRIcb3CAa7VzpeQCFL+oDJo1QqyuG
w9nYJZ2L0d2uPOkfxCaYJO2266Xu888/SgE7TA69tL5AvEGvqmwJbrLeNNEF8muA
LlL6opZDQTKcPbNf9aXGO/UVZQBir2jXyGj85SKMX12uHpStBDahl6w7qgJ+ed0R
8l9YevTTQraSnPXQ8nxu8U+gaWngh9Nhw/pWer67BAkGHrfQ0MsYNlPN0tFLAPBW
lGgJT88zLOljTqzxBhR6CGiizBAgjDyquOexAFJ8bJvNg6qlMfbe0hSw+HFKX4cJ
yYN+2h5BQk2JScwiCQgZZaYczA1oGNasmrIXEtdjc5RYMh6yOtxYYQ9qT0wnc4Mu
+y/L/HY4iiDPiBYy525B0nfzgPbAk7DFZlaC3dHiHRLEua0ebFjF0DVDpq+jg2CR
NkNhpb16GS+ZrDMPievsWen5EyIJ80Rt7pJ9QLMoZ/0g/5yCIPaNAhsHHsqxK78/
LnAaVhNYtbdHqdH1WT+SB6UYr7/I1Zw069Ikn9w/Cv9pJL9eb0QsXmh2PCM6Kk4T
4BBuy6/HWgP145LZKdSuyouamLgKVs5pe+S26GWpiwRsDobEhxxZct8NN0ELRCod
e6c3ENA9viXThZD6g6DzOf41CyYuB8/rxxw90ZkFCmdB0X1z3Mi4qZbTAl01TM2F
Bu8qc3dDZKRacJiEl91PkxOemDvwD+ch9NdMs2Wzs8Jer7bbCJgGZhIQqe/eNwaN
MeE9LVe1MCDmr7W9Uzg1nPKTuLL1+AuF09YuJUUkfNW3K8OTGgvjKsfV6HidJbnk
Qkp5hdPfPX2ZOLN7rYjPxv5eItBlXfwYxpBumjKFDJ2IV0RRHSbjWuWZNs0vkTXF
RbyOSGWIxgwEr/tdGOzveBF/mvHoBbxp9SWaGnIVzuh3lFKdPVoVL35ZuY+HtUc6
oMgtDnDwFDAU4OqLi5Hp+oVa3ntuo5NbtOYLcydfQKguMUONbX4DrpE6pf6eHkKh
ON+aPVIo0swbjIo8atOi6xQiHrz/ChEY0KiCa7NP3tni2fXlrlCM0kuZnuY1dwX/
XYy68iaQw0R8LQP3qQZC0TtKj9HnlBj2gUFM3GMDwK66e85htvws7/Nxwg7C7KsT
qYOLMeRj05kEpdk5EHHZqCd31momBEBeytDCsd4ZVGwQx5wRwF8FpBjxqFdK4ILG
xfs8aXJt8sp+hWkD18osNlnPs6w4iKCy8CO1UCqFdySzxKMtVboBmOMx6YmD6XI9
npF8FTX2t/+511eDhb7sHblxIN/jhvK0Vg5EcPOfRdldpSTHgtTdLic4j1jF92Nx
gD2CRTeTsdS8tRLmTRqfaIyWMtC5YRhJ1dXuKmH5CFijj/D16//ex8C/DjaqDEWt
x1HqPmxYnNwGUHAM23LhLdIvvEyBv3XUWYvnJnSVQDdcrRPwy5d68Tr75hmvMQNt
vJ+jIeGmKm7P4eBB08qBJXkmcM8kDcz+7samDdmBIjYXSIsAQZC+EdshdxurQfO/
NaDJnj0CpnzxjWA3vt+8EV8+BTTKeSQpe93yBzzQTWy02tNjGzuXe59n21rvyF9G
h728eFol5b2KT8/nCcPMcrD9gA/8QThtMswuIO4Ntjwf3tuxCH3gNyP5CAQlmazt
TpeJAVfEIdrM1thQZjP6MaBqAXgLzP23ywwhlCQyZqTxY+gsTQARxSQAGvktdcF+
YlS59TIZxiEAsIHaP7Du3ZcMfiJG2juWDGlFow+HMwQNpWNobFin2yeUExxR/fw3
hQ+Pla3nv9RC/E0uDvzG/UdMj5vxksCsA2No/QJwhGQ21cwBKlR+MNlAOy/kNECI
O5Kq/LthK2BdBUDfq4BMN1E4Vsg3novWFMFOUIVm+Z0Rk9YB0EvjVOVuGmFbzry8
WzFJ2QlsAUAqqRuFIOuAVcJflLPbNjYqrVJ6tTKAyAZ8lONPAtfRv0EJq6BzYNNZ
Zam3foMIrKmD9xOBXQWfl9Vt53sF+0QHx9jKV8wmDMYENsp4YV2WxRIvos6iN+9O
DQIBHmLv59mNAujcOygnfraPF32BfE/YlXHYe6sK1I1YrLmlm/2jDBKzr5x3OlHH
+2eqh2myVvTp4Su64v6Uw8mLaaIq1y6kmKmfVh6pn2z6UjwNQtDXEDiZM6XCA7JG
JrDuOwLRxZPej1+tHd2uytSKSpbjckKyR42OohfEFJEwguh0s0y9pe/n5STAiSH+
p6c9TtzfEAdCBWY7TWaReqGKoBLA0wIZt8ZLy1vl2fI/s4+7svDE99rodJ0CV2Ly
aaSLKgRU2NbcGV/35Zj4FS0MCgpX4Dk9hlM/F01nGsE8lVbB11+VQVn+Jb09V8Fb
aF1K2El7goF/KtRQrYo02ltovE5j6FuYIqFIeA64rGB8PN42dM75ImKmAO2zylGs
RUsYyHNgF4JvdH8M31fike841FHQX2Efsy9m0mPIawyyie1+JsAze3qjh5+IOpNQ
JnW2j8zqTzBg0kIxsfPHEfkurjFHf+lb+rLm3EK1trW725kPMTSJfoNJ2hdHZWXI
0sVaGeF3eKPWxeMgYOuVDVtTR48or9pLVqQfJKHBw63qXya9xhUlREMY5UBhD752
P07l6HeIDpt3U2CtZugx3QhdfUErHpWOBvJW5/+KNz/L1kuWeg+uAyIGN/64uvF9
f2sq+npRS/WL7ZDqnWf4oG5hvcKuDUZQektQr/PPcGKVBTIbn18f7nA2W/BVAoiE
uldNEkXok2CwyKRTkXsq/pGwvqArVvYdD2I+6kEFLb9q/a77FJjBd9MU0VKStOra
WLpt5j13Bor0Xc8HA3D0VR2WPqOFO0rGSa2iGsSsuIiLU4fxtXsUuD0Hl7NfS0kx
1o/MepkM+6c4hMBjeWUURCHYn+SAtyranCvwwFXjsXnneRD7sNEwilEYFwoqnaS5
ZCdNLlcqqg0FhROkYhM8lYFt3/NnsjA8Hl3Jg1tR2pIBcTiGZRNao3o8d493Yson
dK3i3Et4lhE/PEb/6DFleA0wZM07yHSX3qRrP0yCrbDghWargD0TkYzu8tcedxsM
9zCXkE71mpfDqqG8uozFhjZ4nnlU28ixus8nvNmNQCpsr4JNntR1D9nziSjuugzO
PpwfbIe/EZz7EUKvDcJq0AA/X56VhIG3+uY2clJTzfPbNOHfhctjfcZE0M92ZHYE
LMDT8tppTZY5wq3sUvjfeFiPxkHhm/8pATO56AoxB+5f9s4m7n/d2UaVE8zzE+rf
78Hj8oYIkj4WgWRFPKnhGmBM+jOaeYZziHWS7YrTRhnkCkUgJQ6y4xAKX0vPNRIs
zLA2MgSYDIJgQ9Im5ViIglgXkDtLHbXNRx9Nd1raew694Q1KGurkLedRQpGZdr7B
3S1S8gcn7/pXFz/L13iEO+X+MP4bY9DvGy9DmiJK8uIQhMGAMjBBPpG99vYGLBpd
8Jhfupr96nE6R5wAweTkDeeo0hV2MAtfHTLsZdWnOX5Jo5DdrqGyMixFn5C20hf9
Q2cweO+MGVJCiGKNHV5s/N0R7+rB8aY8oQerLVdHPr4SLDTnuQXlnQGoYQQaWzB3
RyaHHcYRbg2RoKeyrR9nO6tVkHn7hFpLe6y5VYRAYF9eKK73+pvLn3IeK6mAu0p2
a2adwqM/8w1Bf4c7HwN6LiXQyCQNdk9MD3moCuKmDcUreC7SSHdb88fr0a5aXY+/
O/7da9vqIKEUO7HRq50GAgXYLNReoyqti4Yh/fTIX8CjFGrGxVEnTJ+g+DW30m9a
GlgjjS1IdloNugwuHoRW38kKCVckCYDkWx6Cdxrc/VXBWdUMX9f6mj3aZsFyeTUh
4yF7IvORmZtX8XTj7o5M2lBepJgiZOuGtE0Ou/FftvLUagb90i3jVC3rc9Vs33nf
tRli+YESsm6DljUWH3aJ7+y1vvVTrWzMFFy4x5qPLxeizFcZkwRDcW5oduaYmJ50
vrN18owPFPCSmP1JEXeGmA/Pb5QB9gcYtfnkmMoX5oUFM6dylDvtXtPnNLVZ4llp
EllGTGTEfCwgMC3lGc+wvln8XhYKk5keToE+8KyRKQs0bsE5vQL/kSZaZ9sMMxep
VdhYqDOK4CVtrM6JkOGBQ5wwU4eC8YWonIMOApAJOgTo5BriZaZcumMTjH9hfFAz
FwIiozfYX0HliecZzkeCzCmf8+19WueWCup3MqpqT+826tB2q0a2bsQ6TyOx+PDq
lSsEr2CCWYnhpA9hr6Ugozua7dzb9UzWnufo6zAFDJuKPv98Rf0kea9HsOb02Tbb
XOjOZ5vonH6uePlwk5er8okfnTxV55dgswognRiYhhSUyqleZQaX/P5pbQvBTK5U
7zp7ihSbY9sCoozuWhVFcPPAg9rd51vEVK78me11yKk1M5r88+JglXm6NqVnn0JU
dL4xhLme5FL38o3bB44oWE8LiNVTDZmRv6IyduK/0LpTnlUxCXXJ7qwzsg0Gspt4
484Fh9cRZozmv2n+CbqR7TmSxk6s9JDjSTsxQL5s3IHdDQ4G8CDXlE6RLfja+lSz
tDd6r7cpAP+YaTjMKCPMR6KE4lshXZkgNrH0vctWTxf0yrpXtzynaaEjyiv6UR9a
764Sx64AKraVpC2cljljpldFDVtPaErAz0I5T7HB4wzPQrcwe3yxBOsEl30Tfx5G
buD5WlXooygl6USGigCUf4wAj9xC+u1j3gw3Bm9hGNfRRecbET4Jk4Hd5nwaNYZH
za3lBJHriV3ADJTpWMUsBzsjwwRIMZ+WM8McYTWKyG+mzV239xvATPhTu8oYI3vN
YJVhnPAEDqyWFE5UkMMsQDPwxJDB4gQYjC22AtQsgS+bH7EGlA3s+PjrbmXOsbdy
yGNssultvYWVZpw8b5WYLyFhVYvbVt7ZZeDrTCVNpBD+V/4ZpgbyHcRTRBodVyQn
Ej8OZREneNGkxLtiAgKETJfyEF0lWmE1X6H3LETN3vwqMwvXweLVcTEflssWOU2d
v0fwDkh6s7eyHd1OwU1lKy1QPpXBx6eN/zqWI3W9+fO8mgofQ88T9U7jimQQiP3/
YJwwz1xyvu3QCO5Gn9GrATrYjL/tff+xxQAa+u+YIGFdctbn4n4+c1a/Qt0rTp73
lk7Dj0SX2OwukA/A7SiRMa11/isRXd5wPcgVySt3n+uJE/mQcFlCLhw/DoaWUc2y
RPHvaQeowfteMua9Ovqv8/lQM+h+Zx8VcpYz38ZLPT3Vr0D6AepAHUk/gTgmiVMc
CeWLjX/n0jA48PZZJA64Ft0CXoDj2i0OvznDvyeDMNNdk/u9vwtQZmtgxj7oVF0p
g+RK14WOphOA4e75PJNPm9NoUrllHtskHK1x4BO20THyKLUkjy7h8vrSmk/8XALN
Os06IZpJCR6U+2by03uHQSTfl+S3o1MMF218hYh8ILB0+o9f+NGSJ+wAZiJSL3uz
Zj5zyXZw8qpUNhW9i9MhmQuwHuan+wEyuFYdRKyFDFwRzrNc1wa7wFRxzMGu3Ntr
cRGkY9m6fSToSey9kCNfT+oGIDqqJdXozssjAr4sHgypuGW0AEBkhP+bv+faBh6F
Nq5VyJDqZDMipFf9KiyJaid+VuIgwvBKPDnY22/fBI7MH2TjBIaDGAnzxua92cGu
3U3evY6OTksoToX8WhY+XWqQChRkud66NG9qcE9C7QAhqDUcZGXFKmHt7l7rg8gQ
U1zKSH/DyJC9/J/FEJHDeufd6Ttxr0fEGJz7Su7BDhcT4V+Bi9QCTsz3kLm+UoOB
jTh1c7wy1I5bavVr6j/uFHwdHxEn/WD2ofmM5avNpz2M/ViDRsKjwPpla6mVIvL2
32K3/VBa/4mZxmPm9I7wLLAvjIuVQQ9V9vftoappFSSNjqL3ctVZXI+yBZEahHAw
j+MystDV4DtX/FdL1mfJ+iYTC1ObBF//4O9Jv1FituM1MW6iYX90+tM9UHBozO0A
lE9c4H7nOxEfdxuSgC/pg285kIicR7/dFV906QHXHbpySIE4+Tj/DZJf4N0z5ZAI
Phfzl9mTy9hG/ETQwnsaSRIkkZ9WgMtZGCARJPy3wRHZ7ViFHEj2KoNnIC9xhV11
87HIepreyo5vFqXF/Lt4eJB1vrFARozerZDyITY+JD+Z2I9b+Ah275RbaCg6Ut9Q
TNpL/hOrnYm8RVgM6YVaptsapco0sXNIer23pBp35hhXFSkImHpe8jv18RG0j+9d
A+ncJ3n09ch7KeI8EU3hD9ZZFq5WEZpK5a1f+5/HSBfrWJ38G4GWzQzhFVJUHKtp
GG4xOVyxWBqrGGXN5esDxVGf7DVbNju7vLCA0TT5mDlDLcyC9AuDes6Z6qf7cXsL
ltWhpCGMZ41RZk/zi0vDnJFATFPcrnCXTIlafmP1e+9K9dtu0/pv5NPQ4hECjc/P
aZKlyaD9WCtXpcRVIRb8YYojjxdcvPtjCt/SkRnF6punldAG8ajiG5T4No1tLN+q
V80VtCFxi3DLldcpCHZ6A9hSx8CpzqA6MCKxtEegQAe7g6R8aiCa36dkDeIBUT5r
ZZfgLQJQvLFHlItO02bDyhJ8o5LWSzVGNUf4AJgcy5lvxGxs/4mUrPxQ7vMfX4d4
rtB8OVYcEPpObeazUANCCeMoNDbo8U6f5AnXM2fwjpapoSrsqqSjOwMnFYPTzSIA
IKM6+8+3eCyd/yoZYZ9WArFq/DXgFgHJypjK7rjn2cor56rTE6lTLFaa6U5lZiXI
aEVyecuT3ByceXbPQqgGMf3aSnJsW62z7TdHzsQoH3iB8fq95udoqHUvYIXOXFwI
I9sq2t6jeMBELkq81G4ZYmfH742F4aaDU9LrMjimo+D4XSUsuaVGVf2jxzFC0cvF
sHLc8cLAG90+aEPDBs3iDv4u/hG3kZHxe821xn76M18XJY2VQlcXEm3UmHECQfKP
fjA7u3aEWnOjO3x4wxIjKkvxQxi9+w/LpjALdUo33bU5Itge0go1jeWI82z35l3V
q9CBVfLArUQwB7ypGb1ESiBYHzMpymQ6H0y0ASjlas7BYTrqTRegLXSLM9koNFQx
SI3JHUFM+E0l37wDSePbruyoulINkyQsblOcMnkR6/0EJ3lzvKMUTrdwWu13xS4n
tY4T2Cr4u+kmSRD+THRD3DQ4IT2t7iHehu6bBSPIft5vkA6vu3Vzju9Z+mOobrxj
Fd5+BgimR5uk1jVoRtywCO32tHP3ckuo9wfFoRPVbjSttvExCCp0AOZTDQqsCwIu
b/6e/iJsB0XvqnydCM7eoOczcr8g3gUHcdiGw5y2cilZKdJSPz4jEpnRZSPLEtoZ
Fc3l38FS/JgANFF42KMXpknSCYsUzbRDT7OfMGMBp+VjdYZJO35dBg4uF7/k9wWg
lOXRbLvziu30BF0DNuTiuzeYseMXgw/bJZZyWF7jq/S7URi0exQAd3+c6ZPAMh4U
r98Gt4RTewKg2FpY2CNBbWaIdCrSqRpiAgGFe4/O58Xih4UAyenzVyC43N2fn239
0YX62Sn4gxCODbsAj5S6G2lBdIN36DQMh7Ss5+UxS323fR9PB2K7cjGlmA2mte6F
lTlcWzq1wlyGbgRjM/5WhhGZo4Y2W8Y4W3ilZCFW1ytyMXjoP4UA8/be/71iQcUM
a18JC/pbZPJBcry7MmphTpvXu2HId/15mTB4I/ZVoKeZUsdPCiZuo3nmGDxivuhI
CDW61POShggZpcVzBeceiKu55bq7ekACWWFizirgU1VtkqUpUPFgl7hRFwzza030
Tu23tMlz2yM/971hXWz4fXc3vUJwDagoZJ1xJXRw1uQj7yAp+2v8qeMCgESbIrYU
R8kY2z4k2Qt98Thb7Y+EGvYkiL73JrQWh2Fe3VjvMO8BjX+thi+N6YJ+UVhW/YfU
FNc54XZj0xjbSL7/lt3QrfywW3vI8rfNEAmzzuNGFB2l6qkBs5N6EzcP6MCm+BYa
FHM718CmVPZMdGa+gQZBBgUhDdrGrOAOZ0q7xwd7U7JZwmfAvwTihozOi8kcI7A/
/4sE7GM59T+soYzvEiSPIrBruVUuZi2NAm8gT5uEYujAjrF0wKjH+1DOwToSmkp1
0pnY1Kd2ZhMfd8MD+6Z2R4LlqwvZyi1wlO6hMr8Urx7p525TVAhl0V1GCPebF+P7
rzywFKodIUJyQXkNvWK79sTkJLFTVPakeoqAAh94dOvw4Pod8BMqwf7JeO3e44XJ
1sisIwAUwhKhgmBuyQFXoWLAymKgzrEJ+NRwWYvhYfjfEwwVskIuxlsJShSeA20r
fCVJlUrhpAwN/p4YefO4nqJ3/XNh511xo0uco5oARM9kjhVJvo3B5+kKKUhhLa6b
wo/afRqf8NgTKzackWMndljmJiS2IQ7/c9hyNDBtDPxZ4f+yZkdXH5irbVF/zE59
J+55chIBE4+2XImgspWApXi2oEKpFGRvbQt5BCecwwBd3dylMaILZ8rpFd7DXM3B
PNITX0NAhGhcECjpzsr7PQnpQQSaFKFEQKTlM1YFYWj24YxIg/u1b9qBt29WKyVn
bneBc1Xrv+OAjmOdkBLZnbDryxmLkPHt8bP1rWOrsalfNxWMepzRs8P9eTGolk9g
iY3XnCIxQpbTSIK5lz9FD0mw9r61X+ggCAYOdc3fYibK8n62Dr5CHCltb/sM2LFj
ndom4jRifDRajwD3obrrjbH1bWkXhC4n06G1yeE/sHaOLU0ckeM511+ZJej1IC1W
paJL/7RkLnTTxHu8DpDmoH1QMxVIKEQtQJUsUa/U4oWziw31GXzeP764NQrgWdBC
0Nx64J9Vhu6zURXX6Z5WOq9TLlBzotoTQyhZjopWE6w71UvHraJAPUf7POwGVkrl
PIVF4dcHtMqaKYP9kv2Nt34WpvPYwrvGmpJqCQ/WuI6ePBMr2nYju6U9kEELLI8R
4znGf3fhrD0mXS/idV03tOcFg8QraowlOIvy4al6IAymhldLzZxO/DhzpWWEswtH
+X8CuLy6l9R72kL1H3fhjKqEwmQW7nZQ/YcEMK94LunZ3DkUqPVR4Lc7MNYEHd5w
GaDPQLiytpTKo1+h1GQXkRddRThPW73t8cZVL3tuxnyMQnu9v0Y0HGuIM0375yWG
eeElphRbXb1yRJCBe7y7LPn9ALscVdhrRhD7eAT3Zlr6M5DEAn8IEjRUXKUDKXU7
QjwQFBqrjxAMKXmhSAyeLhUHUazreI8zWIRFYiER/oZbeaS9ES1e7wthBAlBP+ML
MCPa6nCync7kcqmAB8r3ptAmFabdGOXgKVm3yUgDhi6kk4s2Ha6cLrCbIep5iVb2
s44h3QI08KFVfwFMoC4YSkzBeEiXt4FEVdNyKCdRQEUsqR1iXOmGPRIXhgsC1JiY
8Vl5Bc6EgpZsgF3C2cprLhRsAQft1MUFeKfHq5n1x1nFaWno9bO22ZmC/xQieHH+
DrpsqsB27/wfKhZXH/dGqZDRigHeRq/zx2ty0koNg330KRzgrU4DZgMVvrS2HCub
MeExLIYaZoWc3mvHdyWJnRtVUZApT6lTsCdq9I3R6oXhBnTpJuxWLxiWh3On58ko
cv5kYMBJ0BrhLHu7Hd0rHv20RYg2vArsDtp/DFbwUOhQO0ozugs+gTxbwvuJcaUV
qGvY9S1t5SFqh8w8aE+AF7xlUVWZcZcK4UMdQ6+chpG9L+e22bUO19w+8N3Mae3y
WKM9Mvc38xnLnl5iDU/HD+yuYzGTMccISFNX6m5n2v1ZSDsyecYtJnrlPL+2jtkW
3SUu3YfAwDQ29CrGex9eqUeVLcRRDZgMa9DgFGat3bY+h0cR1So4XBbGxq0RempK
WH/h2JujMXoJzqGH2eY1mdCcqhHWZ4RfnPS3Zy1c3diUfys3xMUWQKc0zo2cYocR
1gFXBZ5RTvQT8tzx4tH7qr1bMvUhtjxlt8heLP+ynsGjWGTOyHy01+MYGN2xYQ1I
cx/EKqiAphMcke6zRlJkmuKZ7KD2sf4FZRZpRaRWGhrs2kdiY8gcYO+YuidcuFe7
/DI9yhEU34uQBy1oqvDnER32zqIZzNXKk8g3eUSsFh5AK8xVkBMHCu9vjy/72rDx
7fw+Fk/iw133HXSdXDeCosypL0Qsq7jD3rdlw6Y0lKN2FflWzACb/hjvnpo/Kr3N
HDZKXyWKjeAEB4HLq6kvIrKXmO0Psdm9H/d+wlir7sgdZplZ4nglSubszCCttxBw
JbyVYnULYM+bGxVKve7uHsCvvYbEwuX3+xEKaIwWMd2mPmT/mMfetKG1+TlhCHHB
nvNUcxOzZQBloz7tpO8lpKHhwVNMDwklt2+2oFfd4/8ktLHNBe4BJnmpbA1IrkcQ
mvh51vlu2zX5Zx3Ar4C8ALSvdXEQtgUxLDigl51J9EwaEjutGACsvwdvjea1fazP
j+YnR6YqqnHk25HDipKS736S0hDS+LwsNJ06/R6VDlyprK0obX+mVj+RAzbW8wHl
J6E+XCi5xqLD+5jM47msXbmt1Spw1d5Zf+fbzau6zQ1q+oAeYoYIq193Hdomw024
KjC/GlZtsyNaD6efCHxpl/3nvEzU08jGEQHdP5ke65G4jV0znqOig127LI3ZlDtu
MEcgtEvBVUiUZUHmSwa5N/k75rhmaX3+3s96CmjCGFkHVB0o9P0s7AuuIJQ5n679
iqsPKEzVn0ngNvv+5/2ELmo2eBWOLzZ8qGxS63hGxTsij8+scjBkYndCLQQ94lKW
rqHZ0ieyXP4UVX8aCYhoj0pGA4aoSr2VnMUC6lv0t6zrEb2Ns42jPQcQoCxo+PdN
ueyadraA14DJUMRnGn1ybVXeDFf5XX15dV8OTavebNPpI0yfrrdybTzCSgywqtC2
hHbaOkAp6z3Cyf0gxUlASI9lCyZTbPtSOuXhscMdK/UcUjzxaKdZv9MAkWksKcGS
UzHrg/RPZT4X3nnllMKz8B/lHRS3ObIuinaXG6qeQ1T0hrxnOE0knwWhjrU6FASK
j4Vr3eYloVQOTCXPN3SM2nZpAn0qVhk7vGycthsfw5ew2RIuJmoHbKoXeYViuqCj
Qv2WiqbdFwst+KGykzLQMPVyy/nkPGwq10jQGRM754SjjMvcek56ZnYwKi1fxZoT
p8sAuQVLjSlT+VwoPh7oVtTnfFeSAiql6hWTkjiZlpUTOOqwaGEIQFX03BXNQHgL
eETQbc7gUKlkHRWjfnntQOtxEjDXSAODtKCQpLuEccwiujNZyWhQfutiKKCLZume
LS2ZR5R2UrbfV3y6MTH8YyVINjfvJcibkLmgH+1XZISz5rmatWjUrS/ui/QC3wlw
2JkCnuD7K7X7lkCJw/JxcmJDd3d9kIV/pXH9ZWAcx9lbStlvXtz4L/Oi3LdvHUiU
A/OkAPJFVpvu31YM//1KaaY4UzAos63wLX1JG0IfoUQU6YHo3QeX8c2HwPFcnnht
azdWsIsqT3qs+GILJgjGS1I1kptyVGXkrJRRQ+AZNZS0Y80NhvbpbFvYLVpnfZNs
BoRi1dmXiUvfGREOXOiR26NAMDXb6peRpHVo7cSsEStV5TaRYDFdgxMDgSTPbwFL
SESPBJAYpBNazeX+mbgv1JJwKVqZKUInLwNeeC/N0lbPXbi+EhWYkUocnGGIkvZo
CrUoP9SOsA566nHuXWow2gX0sQOJIIq2hnwFvubB4GCBxNbmUGN198rqZ4SUC2Lm
vSNo8q+TXYVr9SAWVgWL4v93ZXye3A78tLvZwP+vVevGR+/oGwWwOSqhYqqnj42C
jskwk4g8IKRztjBD4xf8y1Dy10YmPKdIsdA80rgKyXlxv42vbMHVkDr1X7NPSpI/
cL6k+bp4DtT1ziNFMakS9D4iMGuV0DW5S879fpJRrcrl4pRFCxm5FjjWsHyjIvOl
xQmV3+GsYIPtk3WMq7e7XvSdJed3Qoad8Thi4U0Z9a78yLFexVJoz8YZmy1utjy8
OWFWwICR61YWmZC0RUQDz5u8VFmvOluLzAI347Oeu3ooL/baroTPPkiURBlq7eHA
0GykmB1yeqJORTmYX7ldQP7lLcHuyO3EtlGJkrioacx4vlB5I99i6WiIbxlUClMr
wCraGqhDEK4nHC4ymZ7Wx7hXSnDs7bSoAH2jRAoTqPAGS8uFIqfSHXz6MT8/gPAm
M5IwF3LpUyeLP1yGGSbS8r3wdmtOmYdw4mpa9sC7MFn53FwrznPzTCsZnHI+qGvl
v8WSpVbi0/iecTUlfCM3w24ZzjCGWtKnvBG2NDEv1iUaab7IXC076003TY6PvICW
nkarOjVF2fIkUSfirFj3+tnNn3xNAelbw2Bq/ZV+xU18sFTwtpaIz6AsPogIqzUT
cxBJAUQ4iVUSfyGO6s7OMdNruJrknAweJOSKXkrhfIKRhhwCQglxF+PBQcx/3V1W
LVNJzJ5tjjvxf+4xjFl4IqrOBYE9QLmnWHwoGP2l5+rTLDGpmPQb9TCr8S+pANoc
P0jyFOkcC24s0xn42eJSNA5uyE4tfU5kq5txIZa6feDptB7lJSGLRrREScew/Hsc
H5qyI+dnsMcdUfdPlz4UDCYW51suRKMd8GsOPkeaw/7k0fvuUUYZAmqYvwjGCubl
tu4ceiETdFDP6SjajhMG3VWTDMMR1K4nXAyYEfZuBoLysRPQgjD9zeSu4zDP65Cy
IZ+1MSBgRl79ChBokmszyldK0foGzZnWiclRw1eh5U2ZmFeoPLurRKZEXWVukvaZ
QB4G/7ErP9OkQyh9L4gi3yDct18eQutPQDBlh74cl/Ek9oFoRu1wVPW/ILvrU0qw
jEeGHMpVfO3d757kLIDcU2LVicexcv/k/92fhpkgwjNr11m9hoINrhzihytRv9Zp
OC4nMvzAMiMqnIDNVy+p0DRsn4ekzV4WyP+cp7Y2BHFP7Dhc2hWmv4U5paBMgMjg
h4pDmYxKwteX+rnlnAhsK5vlyDfe9oY+0e62GJYbOk90DQDq5gm5u+rw2Y73urIB
0DwsjsGFJE9C4f53red7NVWTBDyQWYi1heC3toHEMEwkqb8orVCkcFm+RP0u0zUD
MH6EGN4TlFYF8BqVxZigCVw6zhWN5c6RSF+dnnuifAlgyljbYfIhN0BlVd2PwZa7
F/6qN5PAgLe+/86Mc/E68ZDyjULzdu0Y1GJmqeTsHBGbb0okqgK2m3lltSOahYub
r0ShgtJcJ2HQYTGMB+ITpbVGYpuw2R7CGi5MYR+xj+L7dmeRFqqK3cYD2VH463RI
RFUK2EAa1fe/9T/QZosomTW7fnVyD9fK8i2f+lQsJTFj4LtHexCKACObO1HWcdSG
MGphEs1TCU8/IRwHcJU7Ke6d9v+n2EMDTvLFwCPd+f1ZGhhnJ1Kx5NxT/3WzW4fU
LGWvG7teXTANl5aj+8u1yC+pDDis1fOGI8z/BznEMCjxaynXqhCYpESNmwBe8Im8
w/ISzxIgPnc3s3WLeO2ja04kZwzYHQwI4g3IzSGEfHIYQPwRT9fYs9fpdkVIx3mT
7EhngdMMe3Efqaxm9SO67V8Q50mtle5sKWxW5h96apoKfmtK6bZAk0ZVcrlbKeXv
7jQT3YpXGesI8C1F0xP/mxztDJx1gQrwb4SXl5RZ7dm+Ja/DOdif2EIOqQ+ciOP0
1jYVTdr2B2un1Xytf3qJDI9+1i9COpOd6rtwe6eJIpTT+UtenLw7xoA0+D9xqu0c
5up/c7sLNYfsDNlzjZma7pF6o9ShHsC51CXcc+H3HM6eDY4ADsjjQKqd9tfwk3+S
1XyrWO0NtH3wd//gXG1vNn0Y3+GZ59J1eUCPEJL8yJTnEdOVw511V7S3MfkDVvU7
h6vnEeZT5Rvo64m9dMrs+YRwoxomt9QQENK2cK3UrQ2IZzWhnmeN6UVWkNFkpuWM
LOCzX2k0VeU5JF0apFCVi5I/M2vMWOpJwBrc3+wfRqws4+0UnyOyLuOKbzxuWSZn
/ZJExgJQ8dxXvQEz9BIka43HtNQDzyhvANAUCJFlrW7GuSYquz7Ee0N0cEUuMksS
pKxJc4dmBRmPtbNidsyPgULNjhLLcYJuM2MGOL2LAr9pSQ+/NSCh1D+SugJoYzxf
0qvOajL3GGpO0l0DKQoSlhBfCnvRgjItKaemBcYa8SyCRDfzpcLZ2RZg0T4xn3r4
ZrqB1q5MU+DpqM0vdKh1NNdOBoHlDINzSHZ5VTI8HOsJOm4vO60RliqJ7ms+87QX
xMdoEGxBv5x9X0f1dVbl4X9TFvJKSvh+7bDwqtYY14/3vo9Esx21atTpMaiRhHGz
Ni3GUTOWgabwCZhzTv2l2fhZS+CjqlMQeUSvsLZ9zAvnqUYwmpgyIlgL28C4et1B
yEAja8eIRtlctWTOG5kRU3tCf5opyIXlftgASoptHI0GKKgTbojjK85NIbpB5fe4
1+blwwJwXhY8k9vK6T/uv/rVeGJmaW91cqe+D+FaLs0u86hGj/spcfYfPUANa5Hl
YzJ2LFebEToQmUzpQAYixmhleuJ+2mJs/4gptBYTHye6TugPnrfoEKH0TsTteORW
XOQc1g7ka4nF+kCsE7y7YZif2XVtdzM5lACSq89ym96KVub22PHUUU2Zk1o84NNo
QZHq+cuFM8Qwh11lKByi/hTX0XU5/BNBRKtx3ktBybmEJ859aoJXay2sYZmlk10h
ajZAIVoU5jgKKvAJruwNGov32EBeN2RorXZMWjtR0Th7mpxSYducstPrytt6Y28m
lhcJy8ofA1zmgnsra2owsGXj7tiE6JfLL8uXyNjH6VtzQ13P7B1pw5mOluBDZstV
+DAUyS9uWZXamQ7F0aee7sNpIj+uIcWNOsSy69m9sEq12mXLAV5JUXNrdAL6nwEX
m2ExXYBzyL+op39bagKDJQXmbw80uxOBC/78TVTn7ZZlPaP6sQDTvq3XN2enus/g
VbW9vThEURbAINzbcsBoXtIHSMwpKltUPl8K6P4N02KNfMl6sAfaI+hWIx/Cdepo
puuMMcVUSfPJAu+CBARkgLHEPkyQou+KGWSt/FF0DCOMaMAPySrDn8I+Kd076T5U
5hhRPCHwQVa6WQ3yqje38GSGaJoAc4hVI33KSxXWmPxxBKNyvuXLMAEy2DuiYTWW
eQF3wBPCT4BvHBqHtJutQPft18fqiJn5BV5ZZwLNaKIYKIyRG5Cr38f+AMatyrUS
l3cXOV6IxsdtzY5ePbbDJS5abyYHFG9kspj3GCBJHlb23zJDMS/v4qrmDlKh33Xr
vlYFt5DBDb6h8Q+xHGqw+rDUZahzaFVtq39InnT9jsS0rm+1xffz5zYs7kaJQ+ky
S3VnopULLgKZHrMBufeadRGXB9QvSPkaGH0xO3WW8ktwUNlNb8HafrlDJGV8rdzp
m5BfWlYK/6FOJDvmkEtq5aHuECWHgUGAE4a36nnug5X91oaLBSVYMOSuU3qJEJbv
vBAOFFDVpmBjVwWMI9g2KyDZp3XlUbcAx6Si2XxDNiduhPMRDCWAjabSxI1jvzTZ
sLxyE/+sWLA9NRUbW+Ds8MuDV7THHcKp4+Mu0Lg9c6sgyq6tukPPXbs8cunRLtjp
q6uubt/ckcFU1TovI8RedSHQybNd+PveSuWedkH2LdH2KPi8uF+0O0N6wc7+CDFE
pMosFHw2Wpd6fNgXQPb+5TnVzJ5z/XRfL9SExEuKo1Hcig5EJyJVLOfQ8L/3rOgx
1thm7580tjTpxQIzN9odPrNJK7mnSmsY/1foLke5nIyMfVfdiP0qA6myFBBFnpGh
K5EeR51Vun4DpUeoTqQ7wqdMNauhfO/C4rByUHZt2dE/g+0e90/+9GQsGhqP7eZ6
3YGl1lwudBId/xC+oWwlpUekrt46ymhpIbAWKzPM7Op+f3zyI73SVbS0Jav2UaYw
ZLDmyAc5Ep10TyMUZODkhT4kl26azJrjk3mZR5+iHbKx4ePSiRrLJc7gcMHo0Ma8
A2jboksoe6xhwUdCN5G0+gpYZEwtgo+1C7H6dyXGaobjowoYp06xMKdHI/NxDInJ
n4wlWLDekcOG0R2Zfwo9sfbViLj0s6ItCzVFyEeYDe3ss3F5o3/aRUsjNA9nEAPq
1pNpwvM7VHnphGBVsNsEQYUkf0EfDYXcABjLoxXKkqs10iGca1PXcBWTc8yYlXaP
ONhbcpRKRRIJbNkLDoV7wJlGfzLFdPzPKi5YG5oZ8aADAhSbhahD4dh7De/ONFWY
PO46mt9JAINeTGFQS6AAqDtRqryX8RQ37RH5c+S+CNPTdK5QF7IYp/k9JED4g7pS
4UAeBsVz+H+EyA9OA0MTW2g5Xm1M7K5sZkBT5VJNRD7RUQJ7Q+SzPBj5OyG/M4Wh
G3dgupqSER1Nzlw4mObibT68yQ/tczq9HI5dNDyEC1UezrbgDPgRA5xkvYMpSQET
B/3T3LznaCoYjjd+VBSKaWeReWrW8YBGa8+bcPcJFfyP97wCWjKG9nOJRSOJeVU1
Mbkq30GrZ+jlXKj+Ef2j/KfBXZ+aIYYi8wVsdMCxn1Y6pFSGrQzlFh0jhShhacSk
rcbp9ycXP4TqTqX7AVzPkgZ6awZz3lpi8bGqEreCQGrv31Bamz89KW/FvF+AyBUI
7xEsmflReadId14SusiWeeSXFo3Q32haXpWSZwYDlDWkhDTsv4S7d654VH0mnv4p
f7GLyBYdQC0mQjip0SeJunt5YnZLSFeflan56ohlfPRyeLMQfs6bJjIcxJK2SVqm
d8DHpWOoao1NFRj9oWO6iha4wgv8OF+Bc0sg/rsuqoGdKR2U5PrVxsjMYCvu5o8r
i8TH0Fmw6rdUdRfdvyaiiNz9Jt3EiTRAskZzVxqXh836UIDAvvDuX6OQY2wltovG
aJF3eAoJFVnk02XK3stZLK3b+de7xEYyYvDUW9bnsSs9d7ydyh11/sEtp2IzLWl0
LZmR65zntRxx4TN6XYIkctZGKrlBzQNBR2sz8pWpDKpzwOZFrePHGYJnXTqWGINo
b7p2GNRUMTmvVS4r0K+KlZaR1WSzXM7GxH4FyIDJtDbdtUUy2d9hM6iwXKhxAbGe
HDLOWow7MjkLHfA7XNeuewtsVs1BAi2r15HEuJR647q1uvQmnsdNoxIwDIkCgyUJ
hpo6UE3I86yqbXGhHQXIGsuG1tB1pVbw/88kyz94xZ3zp9WFK5xnsGIGkbbSyxJG
dyDYNbDYTH60Sj2/GB4SZxr1L8gQL5DoVc4JFuu9HuuNVbq4byrkdYGlsYw7fbJA
uLReT4ATE19jWFjnBmSdumeoJr5BZz9JCjdbt3hyaxFsru9R7DsX9UYlUMpiyT1U
grP322k13jat5sWnBOoVhL8sSuGKvcNn5mO591+ueJ6vYv0RLmlkyWJ5P01ahN+p
ZNM/JkNW4qawMl7dX0eeAWirA2Jwo2yfLiK9bvbA7FUv87qu6pzshC8IFFUIefl6
cedkg+fLge2iPdd40pb8FyekTHq/EKdwXYBPA0VoGXcBytG0H+t8EdUHb1KSvmU0
2Qj9yx/pZ5JBzVfGnN1A44+mzsIEQXNdsSidMvoF+UBEY79Whkl+LYCucDY/wlx3
w7EVfXBgYF87dWcdE3pdJSxm6312tk0itJrm+zyXnruHBBTLXpST18AkGNJplje7
GL4Nzghnp44ik4bcyVwAazwlm10c0d8N3qUVkn5t85ZoFXf9CBSnuHRJ90ew1ULK
sv0SOai5bdArDL7hZmsnrgL3gyejBLD4gXpdlLjj6xNg5kU5tymiQYWb1e+Id7Xi
7Qwyg6sQzRsL0sdEjA+BELQAnVF7yilfjzTidy3EwaHkMgBKrWGxK2WIvSnFAImw
SKy4nPAgyrPSSiyF0xhyHsG5hOYOM75gcpMRl7+NiIdxCy9nHOsIAqaTaqLiKP8A
+dYg3oX4dhZRMVvrm5WWPyoxT2FX8dwLbQjf5hC/WPvE/9O6zMgDCmwtkEMBqy+S
rlnhsj7sBqtA5hHIzx98lPFLrv5ybZ5HpFWMJPTo3/24Dy2IWKnk14bJ/pqBkJZS
xV8D0jx4KvKNcOLyN2IoS/tHNRvYDSKBR1LVd7sgliPtDgG65lLrIcIO1qRtmGrx
AvyA7jLksgg8bmbm7jH/ACgwUXfCj0kgjcYBIpRBQJPD4zB4yEqNC1SFqsh8Sm4L
HV+6whQZku6VOmvHrFaRvURpPOp4SxNVTIFZe651qHPwvT1ewTkVvm2ZBMKeyjjP
zB6JTU3WgfWOTWQJZAwQYjN2fXS5Kxb3/GHottTgloUHynecMCQom7TvGRyyWMJd
MtiqxF5px2BCtH1uELihmedUoUU0qTL2kG+BH+tKV/xg7qjsyOQjf7s7VnKBeUOX
VLx2yQ/QA56r/1LDXXa9xK5iS4JAI84mL36kDqDl0EvwBXBkF7CKCbM2tIgVMvnE
K78kPt62p5GwDWHB/zzdQD1g8hxxpsTVZCIfBeqsul9UGjCkBOYJFbyEbbH8WUf3
UVHmAhRmDO62Zn18z0FgrJPFU3GkqOIKE84oUGusljbbTO5K0nBLcuPfkaIKip0+
86N2IJY8gzK+PL95eEYXsyGr4fhQXRm3/bXitzAwfQ/bpXp+bBgvK59xu3NPIeEg
q8YY0t0vOPefW5mnAIgwn8LhUXFNPG5YuHK3vH60wRZWIz4PfI9kRLozuk9/aLXg
4pEoYXqI5LGRgCPJEPKHc5uhDCdx2m3K/HNj0d+r1+Lt/4xcHWV2u9QH7eK0lRPO
q8joBy2p+pin34f56rFEMJb66T2+IV/Hbf6CtUsyWl2CTsFD0GWsLWXDzV40nDf2
Fpry5IXXXGSy2YW2Y5ui9qAedPMuXrhrBfH5sY7vXCRaHkjlvD6uHcsNgSwl6L31
1QC5S3mf3BptOJF+oUyE0YW0JZflDCH4SA1ITbhzUVuAaUQm6Gc5oZ7wCxAqIdb1
/HAFkL0QkSH+6sd3m3ViVEDjpnoAQrRQnYELP+K4o6pWdKGvijC20Hl17VcbjCzq
luo5gOzMDzcRGKtHZi1hhwv9VY9/Q6ghq6uyJmnfe96kXYyRX6H+AO0wr7+L8Z5c
TFM6yECAkW788dWKjp4dw1o6XoU/Y1/Sdksx+jfvpmtDJDu3as+xnb3aZf+uaXqN
CmknYOSCCBviRvQJBcZJo+uKAelAWa85+GQcvzD5OOrkl8JlE/wxdAKRpyx/pdyG
86MCIReG6aaiHI4LYlF4Qnf/xhpLSDSV1BCruTFhlwcMRscN7wkdV8q9qtWsvvZd
889+MS7JTy6ATgYZU4KzSwzEttAcDxMUZ8h4iEmgj7HFO93LoiAwey0R0qpy9F3u
+5SBDA542DEjiVwCiaVv4AyqgSJ3uW6miX38eAROCEu9Ozik2h3xbHCO2q75kO6f
lbq9HIhXtqe13EAc667aDsJB0U2eHCb7mKeBM94i5aaCOXEJjDRDsmWueTVP+7GB
CsYUxqBRswrTARHzoyqYRKv5b3ay4Ky1OsIlZqPttT4or7iigaq+A4L7DIJCM4fG
48aOubhzymeYZCquFuhK5YBIpt4icXHrzg8r6V0Wy9bA3yC/KuEdLUbxx/5DEMdE
YGXT/D5CPe9+6imJWyFn0SGTSN4SKVTwQqWmtPn4TcRl7N9hszL2UwROx/zR1ZiP
6cYBVy2EDHR1qLN28nnj1HhVqwz5saDK9qD7syA/gfXpFoew+QqSqpiR13DnTDLA
H8Un2Z3qn0S6yi9f8vE1moIwfWRncOS4dcSTIR1qK4ME3fGHbMn+QfS/SQN99TZL
gYk/HkzIJE6ac/LdTtVgo4uNPH5SSHEhbwqStCY1DeSfUbnY2dVZy6R6+Bth5njh
fxQu/SPmM3CLc5NIC77xQV/ICJYXOIIfr51EjIRtPa8EmU8MgUMS7ZnLblC94byP
J7Hlr7/EU8JMSlb+RprT+7CjBXz7z3vUJjFQ1yrDn5jRrIGtFdo3ZtWYsFDFpMJW
DN/B9isr6NHmt+pkgwq9EbL46l6DhrB6s1tHYPXqYRqxLq3wiTvDAw4E9eoBlhOX
NPCX1ipx14+aKNqI029O7Lh2s2QbGr9c9HeYGrT8/SYFHG6B0F7VqBAXqooM8odS
kYn4pc9Pk7urO5Ctp+JC6mo3ijQu8Qus9ki7S19ie1J8o1fLDA4cuqI89YOQQVJc
D8LMnschNximgi7L3fQ63FtG8qgSliYL39WCv3Thcb/CGTcddSrdysyNakx05CA0
LQscybhzxBHm+jdK6yNZLwP4bFFQ03DeyJCFR3eRVS7FSwk7tfPUsZ4bGOzHhDrU
UqsDTfboru4E7GYpDnHNUGBLso2ZCKzGDid92gP5QCiQSF/g1nIcnxb0+9JBYvj2
nQD2YYcuC37oHSLXoko+rRoB6VjWn5kBEg0NmekkUHqQTxzjhyP+kUFgoAGLNUtg
e802UE0U2NETSK5mg1dSL/XTeIp9XQsdA6yQsP1n5OBtCPlgaarw6HdMzDmwVBxx
+2ACLMBiFrkL1LBDjd9k4USBr6hLtrH86M65hXwJQ1YBFYma1AC35o/qoalRU+LN
Fgzfmw5jHqqzNmnoKZXrFweQF2G+BnwWGd2CuxWflgB2gGqrKr1VQZxSe/+SQjpf
vNQ1wzhTKWsto6ynMvzLOBGu7Zz4ERjqjgUVXAPSOEtTysDnUuGvYRifLPZTA9Js
qYzZ2S4AWpMeR3cjRGRuhK/LDf1ZXxZTAayOBhYQfDCDrbCNXK9IV7AdFnTlIGtZ
54K7/kNVQeewkP9EWgW717OSbEMoHZI0daGkekCNrE0TmJ0lMmHraYm9n2uPFgBx
OS3VSrLJhmDe2sTCcCVHJModLrFWshoI8S2YjCRjjJC6VCxsVtCko5+qxlr5vcRM
sduX2CMiMwacFA7v2ijiUTAS7JBL0XO8lyFrXYY1oOzL2yBZEefaJtyF7/NIYU7l
CctrDYyyOYq7tNpcWNW4g/DFgrWjzYDA/Pv75YDvBsMoV3/ZL8WCb+C1NhKMtQRM
wI7wAL3aJpZk/FDIFzmIpomh0bcAjS32MXZynJjh8DiSIMJblAtOZ2V66Q8JTGFZ
CYxAdJSYeW/+ivVjGbydZQ7jq0pEhshwn3T9khCTUZRgC53j7otTUMWhOcsGRyWW
rzjqDkWFj1P5hvgRlkjM52uLQztuIgunrDuW4jMTjCaiW0MuZHgCCfcHAH2brKtw
avMRle2aHOqzM/lkWl0OAht3IJ0MHWoSABUsD1Lu8hhXsN3IKsQmo06QQFs8YZ1q
6aqeUZHRpWCnG/iAcStVsAo99U1p5tBNLAITHonMlr2a6xZuXWmLOeybqk9r0V/T
Y/pP94TZ/vhv7ki8Kb7JSaRenpQeZE08wcXxA7mwvEbd7ZDnH1hhrbDH1uzuxM6u
9d3qOwjv2G+zbjpy2FplAm8XCEUi3PchNnYBbfd60MlxcTmz4JN2qLU2901LMWzF
FW8Z+o7Ool2sCHTgy3JhgPIxrY09/XRQ/n7+zrV+BBhbul6T3YE+S1SG9fdpCWhB
3mnfrxgQXPC3cJAb0JkBz8sVi3fSrV3z9YmajXHy5I+r6BXrxUgn/t7WpgSrmjPF
eXn99uf8oOqYl/mU+RjeE/EriNDd7gP5UvktJq/HegBPktxavBJldo9OzsI/v1+h
J0KKblEFh9SIyHluPt4wadlpeY9a64EZDm/mLIwiLujijCGAfsACjMntrGIsBUky
R+eBLmWi5pbATJeTvAEaXK+3w9O/6jfHNnpeODseNMwvmrqgBOmDgoIG8iAqvApd
R8tUUQ80lk2Cq+1NnQ/2tEJ08IqsZtR5+vknZmsX2HJEyuFNezEhXb1Lr38o/emg
hUBDru0z5Fh1WaAjsBd+JmkIk7agWPqt0pR3PffW59KyWJX37gD0yOTl5WVo74fb
23x+VrcLH9UmhCloxHEEem0CSXxCTlfX1dv+6GmonmS9HSnz3sCVeAOAZOgMKneZ
G42SgvFhMSXugIRwtaiomZ+rPAU+E4CKAHgUDKnyn1+Mru4R0KUL/lwIWHpPfVbR
RPdxVhn1Dsqg06sBXRxNcNKArc3MMLmf4OyLgfEgBZpdTolz5XUkU8UDc5Gw33cF
+DO14di6lDQMF2C1ZH9zyFbDzNTuEVKgpMI5FOuMg/dg5GUBxaREqxTuE1QXB16E
7x2ofoW7GkQe1qkY8nrsc71SMqMA3G48YDOBiU1JF4ATn9srekQ5u5bcZ3UV2bQK
siun5wK6v4bxdrdkBALBFMS7e8ZSwr3kz7lCnGs+bZIJRhXSy6ctAmpjw6Ke9QqZ
+p18OXtI7J5fKpV8UHvNvxro1STrMK3KNINv6RNe6xerC6rtwKLb2r9JU6nRo2kL
hUIkc2vc7F/nXyli25RpExG8qIK/qfmc2f9YSIR/plVL5b9TtcnBgEkK0s6FmOPM
hy4ebaHkoYZDJFK0FqJzQfFOjYGflbN6uW1bf/NdA6sIgssZaLFuGiHlDyueFXrz
BYBFmr+dNmSvMFNqorKByv4xWCkqWDtFl4iQdBs9zq7hv/RUUeo0cwBrqTrMbOiL
wkRdpHylw3Fe4yBRVP4vRhTAiHonCNa4u0pFyQmT+vQZdwGFZulnkIbl9B3dFKDv
scDXjyMwQtmf+sX/vYMZBFQAA8SlJ9LZYAyZba7I4in2FacDAXEvwDwTsDMdgPed
fFRDjnFR5vIm6T1C6TLPcmQ+vxj4yhCjJCzee7tCQS8jsd7F3Gh50R0AiUr8kwhB
WzXUsz8a2vO3GFOzHVKM0bdxE6fwbnxVO8qcZvqQ1KlCQKikvzqEMpeFwlMhtFPm
tQQYxTdj7LCk3H9J8ke1ZC/arbAntVuNhQZAug6Msmb7hXNtgInOjJjJcpOLH55P
jV3wENMdSxtnEWKU3gT7A0d0AlZ9UjeQwrWOkRIpjHf36STXiekDDRyY5af+kmK7
QzXaqSC5O48oInCaqah4RpP+DZB6USNcbjK4CGk7yoTzP5XVfD+EzYmUTJK6fKaJ
1o8ehS1AwpfpyWrazY578QjZdsQKh/56V5b07UBfVWByfdHq/hqqhsHHFhXYW1TY
bYx4qjRX277cTmRUde35AfyflaS50zrcXuFSA32td3xEKoHBRskGjuNvSQP1xS6L
XlS3W3qD4nw6mv+SG1TH/5jxbIPgQbmfaG/8M0WuuQQxWQQl3b6n7tSb2ozJoyXD
hlPcsrB2Y2hcaPUpbHMPEaHFg46KRjGmBIg9Br/df5QSjBdqTd3AQPHJ0P4aEZgj
mBzchvU0jdzFN/0rOXOVbPHOFKDBl1Z4oONuPc7gGR9cfdDMdk53oZiZhsrqDVil
UleS6v0zdY5xivY+SmIIzBJoiUuEW4bmaFGkTsdqIiePNP+W4rfaWRISy0zc0PSu
uVL0W1MgHBEuYJgJX9s2J4Eu+0LdY6+CnoLYeyNZMUxDnBJROMspqSZwcW2xxsA2
BrIbpdwMnYqyT88sOcQ9LHKF55Vr7TTwhkmFT+C6fHiwflwcMXAtz65abU7w2tLo
v5DLDFqJJyxsG40AJIy+Fox6jC2Xrz7VW8LSQh9kTX74kTVstGe24NhlxcfFGRZU
1bfvNhhr6qyH6nQeN5IG8ufRPMcXHMsS9hbsqgfUKvN1CCrZsjI5tkdBQeZAKUY/
pmsX46RlDjB+qd50SAFP86btTJLE6BCjH0OmUpKYzK8i258+1fzSsezxIePy+4HP
6WdgbnhRNIKpgSkhFPO9Z/SE1ZQr+bOlfXEezzM1lQY0h8L+zKc7L0mKVkkwe64F
at6KXKrp5SZ6WVtVCTl9G6r2JQLYwtHxojsvI6sZ3rtrIBCfSE/SL0dAM4u67tmr
K/58/XC103AiQMfDyPYxzdQPx33iLBrFWlGhRX+pyp09cQwi+TAWoMKm1KHlUHLu
2KHfn+7YujkaFrvWN1uJM3vxkpnFnNd9LqHDuukKwv4/6kwDCyRPnPIPJL3NKTri
noNTzRtuJU5BWVNRlkKcEvMEkNsr/DEO8Jp5eTO/pai7ZmX2zmjGkbfSR1nS7i2L
IUKKQJ6KANlHOBo51EpbYCEu2K0SAZRjslM9MgNQKA3XLTuuwi6GO8O9kpoWInI7
zXXi/B28wB8z+Pyuu56Ag5cHEWwRrwYe776M/hzf3ytJzEBMlZtDspB98uNs3SEN
ply1sJjOsyIj546agPaFwFKVFk2S016okUdYYd23RsjjuBlfVCnaiSSe9eu61ZgD
tTEJsVV6R0pWV5cdDZs8jnKGlWyblN+xXnJL26B99QV0ayR+D+N4Ztcw/xuAmanZ
F9wL4s6MQQs81s1FqXTCxFWo1RNNoUdaqamWH5IO+gmmd7N/HPjtyD4JTah3gk7s
s2iCB5YiFNe+B2oJC6Lh1R6tu1Hlt9SeKJUSoEHhBTHvj3SeE8AY3NakfH6OFY80
eCZdu0+Gq3pVQke6Z1XPubhJoPxVpQFqd1774PqBj2PxKchVhQ3Bb8wsCnZI7G9j
UqqlWaiUUAt8ocJl5aWATJnJCP5C0wNY3lbG9ApzxRN4NhRnNsTRIZtcK7k05Ks0
PRfZG7JSTyPUKDdVSf1luUSwlbnLo5oPu6+QAuahePysfCjN5jok6ndFJIheRTAF
ic0j6Z+KQajtjHo/HWy45AliIFbYVD39zOKyfebKs1zJ6UFsQiT4fIvjWUmZFOGD
Jsnn8Ao9U3LQElLYWpL5QsmZe5zirGDB2XIvBR2vPDFo3hN7u26lXsIFTaq8yNCF
edHHxjEDd8qLKgiSGHTbC08oo1iSxkEO8dsSHgEAoKhgCNr4oLnZcsPmGWeRd3v7
1ikbXkoKPQCBni6/cR+LKWBwolwB3SFEFo+t/5YNRNIHTqa4bfFKjodKaSRcIBtq
ZXEjX3PgHZwnibaUIDuvzEKF8YX26OTl82h8e3U29emQiZkYpUSF93T/XLdJmwaV
5qjWX2nqqUD/eDw0ot0AyfFJ2rn6MdBje9jebV18vcxho9bvB6/7xtwzJN1hRGph
9IdtPdQY4NMPDsH9NUi2QkCegNYM9YssXYqGSYU2yw8skkitHFzkBLKiv/dnT+87
nCY0vwtnraQ3zqL/x77pOCuvmz0dsLBsbLyGiM7/4yMFvU4w9D8e0EGmo9UoTgHv
/TnEueuMeJJgFrPclxL1TkRtyPeDuCFiskwx8aGY/7+rxZMjdGtLYJ9cxIE7LQnq
u3DI72/gnXJfafUT2gI7L9nQugJw29F8HqcDXeCiJW3APJ0sK/UvqB7/WMqUkXFA
l4IVxqJpw/YCSvbSaE/A8P59kEAo4IwUwBN7GIbXBzv1+4eO8J1XpIPNmPyGy7oB
9EkqHwNNjK3U0voQu3a5gMIadUxPJ80yXzA2AUzDvOVUkoSsMlKhpfvi7QYJP3nk
Qg5ip8D3oXv4lYtWEKeX4ddebPU6NAQcZsFD0sGzmoM4Byh0tXcfCJx5pVraL7d0
3rDESSQNS5EGuGhQxURg4d/wEW7evmtXsR/wwp39IUm1nWpfyXYv22h0GQxjdOrZ
GD9oCMXToamFrXdXmyqNU37DWTEdMiAfc88D0Ej47B4fyrAaFmoRYZx9NljExl7h
F5hQ/8lT9Wb9F/qM739Glqg2HbjIxhBQNMuZp96FZewBGaCF4eiD/d6x3gJFOZZz
zZ5oxYMXlipC4hGgBc8oxbUoPqLQmzu5ckcLBQ3Xvmy6S65Pk7It6ki7YvHHAX2n
N/PjYHYrRA4/9Bay9wJkD8ghbLht8FwiMvJ2UTb9/b9Bg0B4y6a97yKvFxip4imi
E0vjwkMl+cO+Vw8xTorUK7d8tLtAZoOK8HrgKVmEMKYAqggDk4vvlf8Fg+4ooGpR
E3SF0Y5AlHIMX/5NSqPavdRwjwkBSgMVLzXQXCCVx1AzXriaBI88EZhSgzX3paSM
bWoxBHnx6r/Sn2pFV6+omESaup9a7y8d7HE1djuteYUwmi+J3BIj8gRm9vM/tkg0
gAp8DVSSOWito7D6/ti+4G3wVbkzQda4VLiBmPIP2aGIL5ymbZthaHeklRAyNjxS
AXLQVeLFADrgmfb++b0MwaDWhz0eDctj20gTJ1zIAIIMOn+VoXJnccvR2Fma/+FK
gTQEbtiMvrRIklrfdQMWaF7kCJO7oZnX+Fiypg9ONUqXwlRmyUHJlVSFPpIobTUJ
VBLo9qhT3nfKnwx7iB3PT5Dvfy/IwvtkFnDyQarVQjw+Idmf1TJ+TUPtkuJ46oOM
JHKFeEbsisCQkMQfw1pHg701T+iBQDmTVGB8yARFCYMVEOV+DTc+Lxpz8GbPzbF0
L3H58IbCR7MIusXUaRTV84eFU2E2HwFdlwtDu0X6iQEzSUsV4ew33XJGc36IAHtE
1ilJw1lKDPIhGkksgv9/IRQi4zsashl4bHLLBh3WK6IE6qIfSc0KXF1McWyjlhSz
C+yxWU+IrMuRE4AdDwBHZQaJmgsQbBJ29kzZddGHUnXwGm3nZhUjvwjuDAJR7ZML
LZHpm+IBbp7e4oUYfJVR6I620KJvAGrm4yq0tYlJcOiYYtHLpVORwsfxhpdxR1Fs
/+rF3KsBm+s+9AFW+x5L7rz0ed7FYunLv1BFpXpkOzBm8vBODwvV2UypPP2f6HxY
47H8yJiFB1BjL79vc4NX/SRMSAQAmVD0PXx/ZBsrt+wlegd/9Ya9Hs5Sg7cjzfYX
JcPQdY5oTZiIQ1dBxDqetO10JO7m1XvaSgSgr8omUQUPiv3a8ZO8DbhZyOgRzdFE
6YOHPMVLwv5XUk7ZZB62Vask39UpjmxrQNBsV5L2Gj+oGqxMoB6pLp/wJGXDpjkq
S5j8RG/yZE6DsfQ4rC/l4oFwSYaz/uT2ESZGz2BceCojIZt4kMbMpgEixlPRX0Ou
7eTyCJdb9lu8UVFkSnGOzqhgx1z2mT/FP55p8FesJoueUIOtIAyn9+OONSJ4Dt/w
iAEacdw195cGio5fnKQ8gNch2yu20ECef/Rh/sN1a7U0re7a05hi1wI54NCcvdxg
RrQ7/KsoSpGM9ll4FOvwhKq+TrlGLMDTrD20qXFHuIy3yWZ/72gXObmM/riJOEAz
81ddqTjGZVnwJEFVQ6npZt1T3efijlJ0lQBifCkwLkWftRP9Xd/FtEkhBNo9o2mU
5zYxFi0+f/qzKMjV7y1i17DyUGgD8AYa9CNjMLrNi1YvmpmfD4jITl+KMx618NmY
OWAGgx6JuovGkq00u4Ueh8FzG62B6Xv17FcU9lWkTaSuvVq6khFlxpRJOSemD/ZW
GaIBk6R19pAoHIgPXt448Zu1riRZSf+xXD5ErJ5OHyClmvXKqgtj74rPpfRACYUP
XZB3WEZNj5t5fOhp+gBkFzHOY9SbOcoC7A4a4ClRFj0luJT1Yx6tOH2diYBRUruK
AZmsyCR1KEaX7WGBis7gU9C5xykd8vtpDiRGO0AgnSHocvKwZ4anD36nC1RUFbbU
31s28FvHbNEQrucSR1XqpmcV8a87ElfiDza2Ew0yQtNkYKD8BcsLuzhkE/8uQiXc
fRgB8Ru1QKGSjHD83F+Wc4LIFrVJPn7hiZOLmcPVutIx0StSvQL5NzKquA4GhVYu
JBXEja1B6k3fBc1j+ksfR0zC/IAYL6rSnc/eDeyHjl4SnC+mjIYEr3rIMly+yRSp
qLcB2DzDCJZOrie6tJF6FdedajUhFtnXjPVZcs2YHURUSsesCOpcVf4ohM0gIXP2
1knIpw9HaFTr7YF3ZQ+YCst21HZ8U7PyuE290jr3aMf9Uu9wkmMWJiJlUPgXRN9e
Iba+JeZV7B8m6/I/Tc8I2frHizKB81sU1G8hRBNfuR94IC5Ziiue5aT3czqGQsbZ
lniysROspWDH6RmX39t+miwZngclXSPRWlD//inEGleU+n+WkNfqzrxMRHJ2oXhP
v/Qj/9vv08lxrmXgk9MooXUr+ZNxtzynOEdsJHsawfpN+4pmPXEZF/18fWWfOH4R
wNFEB/wNXdmL32WBY2cxh7DKqN3WM2SLxKRsYH6WBMNfnyEq6mChVron8UngojXD
wkBaPqWqG5QyV83WL9k5gyQyGeOxl1zXRLLlmiPwr07sDLBmIbmY7mJIv/ti8UV2
cpRqQcZELvT3A9ofkCwJyZQ/XwMVPfHwEm4vsWF10MFwccrjrKS/kUjp15ynGOai
6sMqxtYB868oSLFsjHsXlN1IZV/Wt+ZvgVrNcw2uEN4wuzRvzCXsN7ssfRMaXp3N
dz+EnZzZgmB70y4c7Rf+GqIWi1Om/XkOBWA9JDhFZ79SCt5rbN1GVa24PZBmUZYt
/sJVwD85dSzNW9FwyaGpp75/i6t+hihDIz957SWZIO1H4nYLXiNRodKHP0AWJyeh
qU8VJqtzWdAw801pPXfqOwzw1lhDF7Dh/xXwvTKbpkTZAfBMqfXzERIl2X6KH8vy
A2zMndgenjfYqDIQSePo05IVAjt4gT1DzOMgiS58kSzGhZ5x2zSs78IrKxjduYh/
qPQRIu2I/K4uzPLh2cp4mseQm4G7I4huoTKrHOaQO4oU8ugDqM6Z/ARlvdWVagMZ
H9G+2AGAHDh6GAQlxVIZK7Yejf2IyjFzCGXHLZanyATVda7TBjr3qJ6UPD0Ok3RV
u4c99+uKpe0zZ1P6UO1DTKCWB5T1/pwdB/jErK872IDKOmECN71ciCzR8ATjt270
PmZxm5qtt1kk4gbXPl1iI1IsWAsu9g/u7olxRP6DqBE5ssFuYARy+IrZ7E2BKrCD
321OkJwTykI9XgYFVuT3enu6OM8Oi/dYn4sZiqYJ7MoSRYgYLMwudDVZhwvUOzS1
G4YQi1B5ukxNqlFNIB3NDLLMZGA2z/5PSr1O83Fc+Kq9usLbDgUyFdIwDZTmVCWQ
WXCzsx5ncvleYeLJjC0hy/SY2P74V1pOzPmG4HEh+GkRbnxRNjOFj6mHo1vAU3aK
mVcpet8Vpt07ExDEHybBM3tDDf0deTub/LnhqZfDf4EPbQbq719tP+rvvN7pyWUG
/Fr673J0TNOaynMpkrRrHCqf8mTfI3y1xiF+sWsZ6JMA46P2Baz5z6cHehiC+o2c
fGEFKCaiIh7bdLm5UzDrgYaKYOOUet6v6mJTUk46k9Q0kcvBB5KRmIQMq+lza73B
7LP7l3HwfyMxWMY4iC7FolsEwF7jtz3X1HBq6go3J1k9q2wozwVmZFJxkuk15gWJ
yL2u4Ny1ir4nIatmyymqWdqJ3rwk4EBE0o0O6aOFS5dzxcYtn/nnPkwEFnwpl1Wa
mZPruJkVvyJoKiFPSAajRiJSye8zDRuE1BHhB+iZvIUtPzQgp/0v2KMeNAFZMz9z
1/9Nj8CQBqCmgxc+jpoNAcdeZ5D0fU6LXDbCaT/c6Qc35j8asnFFE8r9gtyq7pyI
ugCkaedOnQZHqse/mmQPZaj2mGtoRwJ7cl/UtvH9i/7yQk7YFbzBoKfBPeUsG51E
HUFLF1NxB3JS1mViIbYStjXbsGArcf/ZCwoSL6nTlXVr6ACJtenCs5UdtDqdS5g7
4g0wOq2HQHpdeaIcb9GRaH7IGuEbyAM4O/+30bRgBWhwEgZ7JpdYyRJZm7dXA6ot
y8faIVjWPPH/q02VwZh5itTwz/D4wBgu+cVdyznYn4uR0HgJd1ZJSULjcXOpWrPt
BbO/65oDbyVlOLCkxdLoaBuXzdHSVJA0szxXrECQTxKTUxVOOA2HSI3Dl0bU5hKf
gVhxZCUJIp3n51wWI2gswChWXXYHfSF/ZJaOl2OAiK2EQ0aOvkx1fkfa/UUcXjog
w0+c+8tWhte0jzUKDetEIvR914mRfV1XQH6PpIGPfKMD0YvT3REu6NxkZH9kxQG+
IYlsoS1iRW2l5iyx8A4Oo8Q8D1pXS8WwAGjlAXQnymaJu9eEELGdHw6RJISqpXjz
IjHUsG/mYw/gcJqnQzaJLMdt7hleQVCtv9faGtZNbnnIvJfTS/0AOIjf4VP2wvnD
vZDavhCpgMSX8PaW37gU8ziXivnnN0eqYYgSf95Sei4buEtXEqLQPTOxcvqrM/f4
GZUtM2Ab6wu748vfiH68d85TI/EFoLihnp0lqofc3d5SMV/qASJvkvR+hILhH08+
DImyMPD+T/LZ1DYmtAf/E5AG3rUnasGl8I4bKQA8W7iOrn38K/zkovILycWDYCX+
73P2P204e19HigF7rxkmuzYhisM9MKivImUzYz/qZLDkSEXqB8tamwoGwVL42Pys
h4C0HH6i+V/ijrse0iBau+/p91h5XqNPPxtZZwmgEiub6CUwO5ZkmWajBPZNcgNp
1z0WD4pDk4FMMXEPpcuRSrkxPg7dkRLiGg3CGjYHoUXPeAAt6adiOOsu4ecL/Ox5
PdxWWXUgDk4JU1X8HC5P30z8mVQ5Wuc80FCqCEh/x2GLa30x8sAbfik+HSYjKWER
3qKyQF90EgCHv8StcunFgSKZlsXtR5IoKGqO+u0oWFel9J7+yB6XDGFjkUhVjzyv
4xkjyIh3LpT2B9ZAsIZePOEB5jbbppmk2QlmoOVD2RC/BwtihAaGc6P5MaIUrOyG
ILCkAjK4x1umt1jVySyGh7Nai4pmFGO0CQ6E0dPdlFkq2qmwdC13uScEeFB3ua8s
vHFFuUoPNd6gzLj3ictAPk/9i8mxGygP0z5oiq/VkGJi3AtOiSXaMMF/IfD1ChBO
+7/yTozM+6egOnGpzMFwJlTaxOV/jDft6si1s9vXBcpHUz9iXPXtQfx9SWd/wmFc
g9XhjfCPEcLEUY0MKZ/IM7QLpuUHLt9BPAjzuW9SRKR08GtlnkYt5y5qsGuzGKuu
kwizaT3UmZjewubpAKDbhZry96T4v9xCYkhP2ruAjy1sVDDdEZF60WkBElZJSNHq
2PxgZ0Z30wFcigpc6JuBXcYZ6AkdqsXy1ZgdnXkfr/30aRDkvdgalbEKYVbh0ohg
3V1LkYIspwrL9Gpn5cNupAzYgc3DZ1O/uyQKNS1EUzpffucRa3DFQYojxBoyiSey
pS0dr0GKUxiF3kemDJiYWBZOy857OtH3lzo2plE7zSe87gzw8RyWt+OgkyeEDSRs
9rKN8W01Pl2r2l/93ZBTIcSy7S43i0a4+GIMtLYuK5xtwjrNqrvKIr/ivC+44TYr
i3t/LKAsFbNLJ8Tmo5hq+axzQaH15HmZRK6sL/AEMm/4HM+Fk0XorEa0uG3Yg1mW
z34FOiGCOtBQ+4MesqlfI+T8qlUKSFEyANV+mvBoGSORUdgg+Pq6U9lDsD+XdQki
6KgKGjtc7dVfrWwzwO1A3UAR+3Lqe6GAKcXXsWOPujG1PCRRDNwp6oNwNsD/PDX4
hKXPAJhDscTLuXgpl5KSEeCtbdiljQPF8CXCzAImSRZA+ZTzLyEylPagFV9cIoFK
whv6xWY5JfEC5uAVjyT5TJwkdSJqSApdCXsJ41dcRSsKfeyeS2RYuHVSghR55Krx
kKvVDDbE5exblatjENRHRi21MN9H6rjJLAs08u7+nPVO66MM5nO3eFQcbmOVjdo4
dE0GDRpHMNpzr90KrNcww8j79bWC9BHBphZaekRr3iSw4q/LLKL2IuJRCZEgPEcm
n4MFhzTBm/s095RoC2kqSrewbnNdzHOMN8G2yAusbvy2sx3ZhCRnql4Qqo6xa5Ag
ZCKoS2Wetf+EvMyc9iRZYafmuO9XIdWbbk+TVfA0Kp42flRTfoo7kxipNTua1Rhy
tOiarOB2ITyvt/PEB/WSZHGVJZZkRj28MtITMDbJ7KVHv+u+VgqKaZRhhc9jy/v5
ZGFxxyyVgD5CzROLfdwu08d/g6Z0v573NxNFIHGAy8O/hcKW5m/8ETNSl9WRbpjp
7xCI8XgRYi7Yp4yaHG9kPqpUqxHoQNGBBWBvU65JTj+kO+z7jE5sH7o37YD17CGX
CJDwIvCpmdJ/7G7OQ74wdThf2LvmaAB47xs9N01pySe73LjdeP1KmgEmArcpHMlS
DQbQjkXNHGAe6AG4P2AwQJeGp3AXKY8I/WRJGCSdkueYY1tnfTXq2SzGdQMb3zZq
YxDqdc9HicAB5p44B21nkLJSrWrFFeRVwxn3QxF4uHDizYnIf1abUyXqkUhKaB56
R9BhgIo5muMWHAbKyvOqCAzbgs83PUfYimQzAiPwDV0W3zsZkk2cDmqhonJbcGR/
PnjjW6wxCDI9ZO4kc7/pfxU9R6xG0RaA/G0z+amnatqnpnp+wOmfn/o7xD+fjrg3
zECW6ohPsLbpXLOt87JhDFYiMy7zKHYeNjaDMRqi6J83GinxYhQZhxYMaH4Aveov
TYlo72cwAR6iw3+GR5N6lyie5dWdvTSDuOrttplVFxr+B+IDwyRGZvXaHTqo2PFK
lV/gABtceU817Q32gjcyRZ+Y53CXgERTHzmHSLbWE4CnRKne+LgGzyrR6HdpWw6u
jDo6L8mT+vvAnpt3o4efEcL0FIgefrzuuFMbfpn4MdTgbCfpsiqRpTA2JRZAXcVP
552jUZNS0A3kIcRmR5jVi6rYP8aBzCKM4NhdAlN7j2sG8q6uSo/lyeaLssIveval
ho5uRBDDsTQSDpnusmd3x1vx6i/gL0cYHfPBA+WGb9/W1tPy8Zb4unN6DDKZ1JPx
PUlKcvCgcfTnn3xVBwLfQcU5YPv+zdQLhZanqJ1BnxMGoLWjEBG7qB3ZiRxoE182
7OWRrXbSBsPAKNSySlVqto/IperiWrLO99mj8cnzeUkozmYPPf/N4xbRNhqw72LP
uvM3dfzOhd2y3LznMNI2hne7symKiNTRz1VtMbsqrqiQD3Qi/e3rTB2IC8hZTM8g
sTwBSD5aYlRr35ZJyhvZN8NJknzwPe7uSzLIpvGfCgDYoVcc/E8Wv935emwDh6d/
usLPhFFgaWPAytZsArYgYl0UODv/Uzf1LbMMv/pMb6USSpgWgNYeTV3POPmv+7DD
O+adqLga41JRLOJc/OdGRfJAWk+s5x4Uw6yi79VHsZEvsQTxU4WtcHIKdB62JDfY
IdV+4UZcoouNNNPCmhea3Mo8GO9LbNXtxphDQcfayVhIMXez+xgXWN52lp27JWXu
GW7BJVFNx+CG7dpJOb0atCxARjkwXpkchnRBW7+Az93tQ4YcUuThjtkmVnEEFv6u
qZrU9PMfhOKiKXDIiGeMTWQXyhnXqfzlC6Wot2i2YF36hwUDpCd/VI13IbIWtEEJ
SBSVnKDzOxwJ9mrfIoZj9+KKjWUD8T44jwccMtfZ8J4/NAgGHA4peQt1kPh/rHuV
2NRBgPRcGnGU15k07jbGUTBq818aIy7dkY/4C+qOuDfSKshPi0wdHRYuh0qJ1Sh1
vi1hJkSb5quR1bs+TOVGx9xyf4qlzESzPNJdQe454e98/KdqXDQBjdkLOauvZ4ez
0jvRB623TUIg+Jk1pqmBO3Rm8cVXFdkFeUvYOWWxw0ijIiz2k8QkXvwwEhO4KCzB
krUU4zuzXbjXE0kBxEaW2YLzgz+/+ongQSXnioLjWhWgtnuZqW9poiQgymOtZIWa
G9+6h5PDKuMtqeoi/77GuT/AYR35ylNmWRgdPrznUartq2Vhmrn2HDDBhv+IHXIS
Kb7L7lM2KdYIveRtuRpyzZS+US8o1T8LVn9JOvK79zw5yjdeQG2UxvsZlVTzPfQE
lpel+j0cqQs8wZNnN22nu74fi0csXKVQ2UVpRV2pmPoCO8s5nk1y0Navdk/gqKoD
4N4gSNDBpVqmlz9yB+kUqTugyBbekZWWNgmgqPjYEf4JUmYqF8IZ7RL5kUUKkN12
OzQ8r9mRJdo4orOF6Bm3aWUKW0TvJy94YquQZh8T/U/S1xQZF/Xyj+Yvo2V5YXZz
UJTAe+VKwCEz3Oh9ERnlDdCee8dKf1oHWc28WvCDgb3zN5+uoLidaHysi/FtBtbB
p1Mno1xkaSi/cN53/9MzOeFgRJaoPufq4m8vcSlCTiMepgvdMLraoYJZHmQYLNcg
CtK5myYjTGspWJIFNHXn95bRhA4HxaIJ68FUwS6oUIM3RCK9m+WXteSQE2rSHMA6
9HAXEyaaFin/Zeagpn8U07xUXvL4wxlSV1YW/manEL7IdXwRg0G77HsBVAXxZvQV
OF0m0hcUEq/MbNf018P7cxJmlcS9yJlhwotVBZ7YV4+9Kqzb+GAq771f00omg0VK
t/diE7svXuJV2Bt3X4QpHTlMUbERRykmn36LNsz+y3oQIPzt3PJO4kkkVLFO9V6A
oqjNHrGyKbq/JAXbcrYIoH0fZ0k4w2VpmRuwSpQninnHGBPWb5xkr4v7pK7pX1qC
sS1K5E7GdMUtQtyMJkCYWs6TvtXPgkW0lZJ5q2bwf2wMjIs18GCYBAR82dXKrQhX
HkN2DBXSrGerltus1lNZzA/f6Y65+Aaswse7IH30aUmgfdHVmDDj3++I2blqBZBw
p+yxoix9R+u/3QaFk7M7wVLabkht+FdXoCgE0TWB9XnJvk13eHyFs3yuTgMEEIeO
7V6BxwIe3i6FtFb8fUQx6EDU47eD0yzv2qwuCo80XKtHiJUxmhuOCBqfJXnhDTaj
5y21TRQC32Seg34xucza0hYUjkMMjZpln3NEr7lE1ogUjAyQWcQnzLgheOlWZS8B
XawjIRGC8e3J7pwmrq+C9ku+IE6vG8Gt0xSV4tE9nH536L1i35lzBFmP2zJE16s7
utFRgrxnmTZxohOHCiZuSvARy08hkily/0dPEvZOfCn34oFM7uqQ1pr/XKm9Vi1/
UWeS4NKJUbfPBZ6VLseFrViTQQxBUC6LgYQ9vSB+o3e0juAyd+vjETFQ9LUEfX93
s6DiSFDRanNiaj9/rK8/BCSDdpLl3tWSDZmq5ubLzxFHCQ1Tf3Ttq8Q8A6GU5cna
Rm84UzmvwglSPsELJBUZnuSscldwUIzTMypoQvU2Nm3iilVRzFIzK/4Cnn0MfCnI
CHvwFSARJtrKe1coMIeSRgdRAur9c9ArDH3QEgSDPMmDN3Q/a1m74eT6XQwlgQ7m
yU0GV27lV3JL38wzajdRVG9R06goQSJuFoLMsckshArgEFLxGGsqniz/XhKSV7gb
oWgRmpww/FESndXCK/iVVrfrZzJe1bVjV3osLSDb7DSvs2B4W/b2vB5in+DdHID7
1jFDQBDfjbTcAWgvaDEEE+/A+xDUFbaMTJS5g71IJZjnik24E75zZ+gmPkwcXQRR
FKw8LLjkytr1EaHlUcq1RJRBsGI0dokgd4yElHJKn4qg0mIAp+L7WOwVhW+0M8F/
vcdjGYypkbg4qpR2nb8ozvG9IpesE9OWxtpA6wA7/SMdj6l15yK49tyod3vL4SFO
7aDrwjAetx1ub3YRwkSv9H1NRx1tYCQ01i5HiWC8OYBBghdzCGP/Otx1+DRrCvIt
uvxZSs1BHB/qZBGhlYny045xHhYqRsRcTCNoXCiApopprPzNCFX/tZjB0cidCkEI
6icuNsYHQ/sW59nyeoI+JG53G4LxLjCF+PkT9riC7qmtS6K2nKaZ281hmZsFUXaO
pHaHGBEscUj8evt6H98nc/wygtMHO1aoa0zS/JwCvWO2UiQyygHI7PL9YbsrFGXt
G/LLRXEVARrR8sco8SXW+RXX+Uap3OtFVySub2DY0Ac73xSYCepc09ODWcRfu3c/
kmWHm+o81jiHnQaOgSeLzO2Fmv28qT2lXFJ1vKwaRBsrfqtB9qpCW8nwH/rYs1dE
bmHq9aN1UNxBBEsisVErpJaQSqJ6Hs7IwYcDI3haUk8ow0cxS6IKcLZl3FxzFDyA
K2MWmZa15IWgWDu6LSZZOGEemTjpAJ0vYXvvR8kKGfY632pqiJUphGPTifMCaA1p
YAZSymwBe+YMSRt4fb2dGiy/PMSoKJy3YyUGlM6fM1a+b5kzlY71QNxz/EWcHKJB
hVNQFvGklyAQ1FrEQcWFImozUgeEpYLmBhF/jbDFk9Z4we98Vox5HCp3alFy1sDd
e/242KR9SHlC3Dc9Vijele9Ap5kGHPKeFFL73nW9kA/o30PFpKZvVjcoEoV2d4QL
l61vHA0AcxDaKj9ljB6hcBngMEZLkB+vzhbo+GI874J9LR1hb20ei+kAPUSmMZbb
ElC0Ui9KKtTdLjhWVxtuPZ1yGz7gMqhmfURhWr3ffooc4CIHzIpNynqUoM7YsKWJ
RJEfrPjme949I+kUXI/ib3YqmNG/2V18T1vMJUIiXN+xiOOMyFqtS5MtacPc3DY7
FekqpLyiqLEP2g0pMICyh0yRdWetEL+ufGWUcUSCYVFUW5MIMME/xT1Fy88D0w5l
lf5vQDiLOLqXxz6eAnPwewqhnESQIERtfjARgcuM1EQypn9cBjGvIXHPF3FZTiOL
4RW6ZaV/iGDvhzF6dz3bOm28OoAvZvhSNPLL0ovi0Yog4Qtbd/BoBmYcHraJEnig
QMLqjn7iJYX6GdyMXGtaoniPfC8vUqfnp8owB3ROo6cBHrCT6zuHVBLyDzDMpu7y
k9BFI7lModVqL3NUvEOE7gvzdHui0DLGY5Tv/kAgE9kuXcn++S+3bdBNU5qBTYqM
cA0nvztEBWdLqqTY3A5vnBUMFodfY/lQ280zfF6sZkysD32VE4gpkhOkAFs33wvr
Q0Lyug6uqIdBwxr5TUBAGBYMI3/LF2IXrEo5k31HA+2LnBDkJnvi3q1qd5FiKJkm
Ou0bWPYnUePItSs1Pleq+Q8JjqssTOGFSl/gMEF11UZv3KdeCbfPzKpCGa9nZhEd
Wehf7iOzdQBCsYm9ANo94W5TBhL0aHv5Jhdg591Wyzzxp+N9C/ale+UvXPDnOElA
1sdilhOza5/Om6L0H20ecme75XFsEnTOTjwdR9c/OrEo5+EkPpgsb3td8KBp34ha
ksINVhOTyXtn/A+H1YD7hSzX3nza2RHhOmQNZIKgC/VXbG8TKjJJqRBLf0ziPutk
Hb+G9mSmVh9dVXHcGsZPjmEkSTSF0m6uaGEPqXLGqvpJ8ec8DAIybYhTmIZON5jo
9S3fsPl1+JWgGwXqT2tro2pY9seborUnvXcprhY0iA2KQC50vT03cR8biWKYwEe9
lfFlP5inxOExhV74HVyZJNjARk0/tFrAkZPxyyNcwi+eD+c32Nquv6BkgoUZcfaJ
JE3FzucsHpG1Jucor9259C/TRYMSZma3dX/dsrRERYRp7diOrw6JqHFyqS6EFpmd
WE8LsKbr6pxRniOt3JrtOyAz1B0Cxx8PM/IxJzNpAEcume/ufATDnj1/WRpq2HTR
rbGkw53kbt8I645jM5eNONCT7wVaDlY+luno45A9GqlKmaHGO7tH1nOyrRY03onx
ZHByfejtuoA88sjc3MUe1AN9WmAfLyHf9Gd1oUh8f65VAvR9qEPW/D3DflWpeoP6
RU7CPXMmgTqyUQfO+N6He3SGNoWpXjjpeFSDJ2fzpUoaIgdOszKEPyGzceteHYCi
jIsImnURcdFfJPhvBqtOHOehUhTKfxN2iGvcsDkGELgE5UnxBFE11fPC2UwX+yfD
4cvWPH17quS961ctap1N/WbtFhDCyvFlKWyONEifNkqdtyDIpbixGEnBI1XXQRlO
DzoYXlPYdoQYyi8SIhIDCcqM/fozga5I1JsNggBQOmgpZp1D4jlF5hAMgJosAi/i
NM4JQq8Ohx30eTrx+//kSyFIoxHTUjO/gCIwdSThY1b/MHmAV2NimXHJxjSr2QHc
IBQEOvNi3Bst5T+NY5a9QtvDL25/L1c8GFYfgvMyhQTPsSpSGA9ljJ06prZadshd
AgstF5/uEBq1nC99SErlThzN/1AEt7p3flrFXnC5/6Gw2b/gN0ihpB/RsjLf8jmK
XOJ9CVXWGGIpCvypUgEdlghd5QwgoD3VPyBQPydBjA8osK7rzFUFJYjafPQNZML4
XKHSGPZPLLICmE+6zBy8vFYKcY5Q99LbbWnxfb7315qbUITPFgDcJSaoYmEo6Pt6
8+yRaBKYQ6BProm0wN7U1prz3aGB8ieaMNxOTgZs65pfhCcsj3gYWCNduYnkIvlO
b1lUm4AldLnvNlNevTspIe0DDzjQ6+D8VSEzdrH+iL8Yk6KwhIxIubgdo2Y1AIhU
7Y1kwkKlDJA8lOK7OlMczP0aZrnbiiG45sFghCD9eNQ/PbZYPB7Z8HAw6Doly4Gs
y5h4DySI/M859z1DSXwM0JoptwKAzxwgzKRUMX+KDcZUfIHvBBJjT0rKXCE53dMs
g4sMJ4aWTDJEYDvC+rBjvnH2ir8BmZVHvEQy3yVrYdnaBxMPOyfYtYAbOG4gyQ+d
lq8nhxhGlRgL7uW92psI+VyQ3VGrKR+e7caQNAcwDnl8QXGTiZWiiR5BqE+5MBRq
+fuxKpVjrTB7iOrOfHwoAQcFgqinlic5P61umRF+vBh1AdK78LwiOZXfIOgiEEDG
C45KPgc5kqZSNZoqxBwJ/I174BmIeDuBdd9SiN20djyklaMyRteQJoSFvIHIVUVj
oWesleQAWomzpSvQnxcfkdU+DSwfqhy1raOG2F7GfvtpAO5+WrJJfK8p66aGnw0i
q5VGPpOeL2ekVTGyz8wodDHggyd5eYHHYNvFauky5qv5MzjH9cFuFe/cYNRSeMmp
0Ox9FXZdKR4R5cv/LidMsdd5OMsWesL9HWq0xQ422rZW8/A5O9od7n+xDDP7IBT4
PIrx+HsDksR0n/eO6lOvv7Lkx2V70Jmjr9rF1Sd4RmFvgSEuzFjm6CgfbbOoKWWt
grOgN5DzRvnSmqNmSkSomji6Xps9h44KIFB4nEn1D09AYrijkQr4g1l7r4U4TdhA
ZCilwe4nTYCSVYpMk0EsR+0zqCMFS+wUx9ZRk9YzClvpFseX5a2y3j94w4cCrwqp
6EDpTAZftHYpRFZiLCwk3ZEixsH25xB6igcNporCmFR5iI3SC6E2MN/Vw/1CzFum
OyZKKCM/D0x+wXjuaXkUUy86VbDgPjUr/F2EOQS+QHoPuGzlXZYlT0Cp7inBlW8a
eeytpAiLueRT4yrclRe7sVP03qBgl+ovm1zYemYRu5ClDSkGhz15Ze5QdYzdt2cT
sKiMD4wqyvPO2OUayJP1Du+2pLB+B2JSdarIsuSkkZpxtq1Mt9QWYUVZEZzUpNs+
UwWSdvGFFiV/AoX0+Jte6BF+U9jcG8K7k8IOqWH8Xf1aGQAZaDxabeVhad6yG/Wp
O9I6JJw0a38mJf2XeGxPXZ6GC4k7mq2fyQ5WqN1+3SD8TBWCFtQs2EFEFKYG6qOS
5OEeZfueS9D0hP/k9vqsX2UMHRZGFFlfQuOaCBCKWkgf4Ji0aVSXeYce1ZC3YXRB
c9nn279hxS+GqDU81ygCS05NB2jNuZysIQeQxtZY+M/IUZw10a7v7Sn8j8uDZChH
iNV/vJiBj6W3MDO0rJHh0OO3LuJs6vWH0e4r7mPvsi1Y0Ng5HrwSCR0u+3UUc08e
PpSMl/w2VTTbGfd5/KwZIhQVEJULQgt0CspeDw7cW63MhDStyGK6Pq/DD3ovfdSN
5D+55wPMeN8DQlw8Zx1aH7r54gFTjWXtjbFrssJHHm0mC+oSOr1BwN7gByDudSy6
hLLGoiWkZ/H80FUjnb66I765k5krydsbcXcn36C6P0IfooWYMJQaLmW9g/J4Ow3J
97hwHYmTIYDUHsTTHLdLjhx4SqFUmsKRPYrmYBdvbLrD3uquZNnr+HmXusvCEp5p
ICsBRnD+qtc3zE1OmXMXFES1X7i504QtvBJk3aqOuVP/5+6eY5Ikn+pKP0oZeXyD
/ipRvQFi6RY9F+4yBS/rhfCNR7GpUlxbuY+YcMAikUmNQYftOGXPQH16AmcZmgjv
GvYudbHIAlizw5ksfiLkznMI/4XsLXp2qoX48krqUMAlBkmurrpdLh861+3ylH54
I1WV6b5dsC14dSRgLgdMHnE9alD+gwTocAzYZM22LzFx1TadcQwRY3CKhtYJ4NAJ
IwDxOf9pc55m7PIjcd4PZ0YaXvEc1C2WCYeofrXndIx9RiSVxXk2k2D1AxAl4sRV
zTxPYj01zG7RlklcSQyOGlB98VovFAlw//bBenjn1TBhqkevL9wSwoo2QPhfOLm1
T23EqovKctkImzusxfikfCV7ERmLvnHEiQ0YfCp3V5IPvAPhduMVqrJu59ZG4Fu3
A0AzW6cn1M/1BNMOgABCFT7qkYNBpT/CXXPLeftZ+o7fLZOSZ9ETlQfWYo70OnHj
rjwmTeUGPJT8c3BDx/d68I9vJvi5TJiVbi5Kd57juzWvEZc7BW5gehYtM5puj5er
FhIB0iafvajR6k991CbDFcRVva/bnte+VQZPSgBgitTFzpt8cepSe0mdXlvxAjCr
Ep8wo+l+UcPKEaR8Mb3iKRM+ARjzKfMLPistSkAKTP7KEVbFDh+vDzV+reun0Jfj
eGc3k+h1kGKwH1/ToNWnP9Be3ehkKWmhUiG39kb6R2M2vHrXIuMDhd3DA8kq8Dhv
MDwtLdkEe/earWE3nCULCAoVr4GgliWQ4gKk+EzWF5K8iOXXG9ZU6vnudUHYW8e1
sk5FryXIFxYKAQuGkh12ja8h5plq2TNGTWdYC5a4RGt0AlngKYMFG34VTgPu/5N3
ig9JVOqcUMPAiUPQLpGtlAv5eN0L8J/kYcM9+vXVQJ/crdfAzw0tGxzAxEEE0cjh
XsHYLjWqeOLu03e8vsiz6NbtgAWB6EBNNaKMDoP8b+AY9cdNQbAhF5Bw3GBvSjIT
XYayTwctM5HPSKp9pWQi04b3k+oMFHawrvbDq8C5ReJWIib6Vi9ayOPoOWW4AyaA
FBQ86JAdTYLhshLfKj3OdKp0s3njinO1xXERQbneeDFOHWWhugb2hTJ+yMkbftn6
gxDI4E/ydzmFCGYEpoUO17yVQIorvUQPSmR3iStwtvH2C5PWWLi1wS43gs6bT7q4
l6pzWZqnFmWnEx2JGXoqBLfb1XOZYVQUT6Yd2xzDOSgYEttGPb5daLswuXxAQ8Hw
WF4Q9/mswuML2Bn5b/OW3OP3Xp+hGEIbx2PC/wtwX8tOwXO7MiwRooqPdIyixoOm
+/zHUyM4rmc2xxYCQTEpts+SMMaFAsjiR3eMVtSzfxp5q2qY5J2g+1LMFSI2Ppz4
mc1TGWscl7YVlU0JSnrWxapcU+LgHx0QatFKoKmdqO8K7fSSqHJNzFuAehkCWj9q
Ki5OAYF8U8zW1fW4eJbbBE2VlC9itXoBUlSF/pkNFbQU48UhPW/oedmh/3Xoc5u8
DpQ2O4v46Q9+Vpd2hzBYcG4k51ILAEiQ/cCTOQPpb/izaqOYZ75OBTQ+vXCqMG5O
cXoWz3hHu8OT7vFcCifQ4Ma14bvI2XVx1o1GPRPW1lUDndzuz2ZD+TKjBDDjtsoD
l3ubJ1ob31e7sCaWMcyKdPmzM2Iu8ft8QTWOOXUSvAGL1GiSk4c+o0BMQHA/az0+
ao2BZqaFVOvzreD44TrxSkrnNXbEOyLeRZ2tcOox/E/p2kwg2sLoNmsD4lsDfs8F
Bc89ToYK1ttM6s5meVxF6zOfr9ljCgjZn901zbxRSxN9hdGBR95DT2PP8jGnKKd8
5ZzOcSktZd72q4lOVWI04juebxCokCwBddvsjc1WQ6L4XAfass1+8sfBQXCcB72N
b2LKS5TO/uxquZHypIK7zZsDuGDFs/S20YTuPVvQwFdjY9a+juUzJE8Qd4R253O0
E8gu/DD3+XSSEYonz4BPGP3OATrD0kOZXgQO10ZqsAdWEEqaDrywFLaNTK3dLzmr
4WxmL+/2WGYa8FRTYY5wIzgDUwjS2l+/JkdYYzGJ7oGSkcXTMfxw2d5m3wVyj1S6
6hfhwRT82PusflUJGG151r5/oLpAR+4qkqtjT4brLQkXKLn2h7DEqfI1A91+Qinl
xdQ0kGBrUiDIZLzJd+8qYX493yWRfJAM/LLTM9p8ae/+3s3W+/+KEtfOO2q0QmTp
TSMCoIV2ZN/2dmfc0inMPi3nujrD1toZBX4XtQwNK4wM2kY7qUShyDcfMS/ZN3RA
jmScRjcHLYue3ypdRZ2vqbk8iPbyYrOfxy8/4jqPtQ8WL3TmMWQzTINGxa4NyhCx
uZ0hl9vclqFATzaZzfwSWU+r9xsbiRE8e4yCEXnE6tWLFd9u8d/2K0JXlTlmYIDn
nImdvaQcIGl03gcbTitb97+aUi+ye6nrY7fbIBmhXIIlHpAlDOfvrqqGYEx+nt6f
W4Tr+fEAbzotIFktXSTx9rnz0SCC3ST2RhZLNem6/MgkwqJzvoEGH2fXi1331iU9
5KmOQ/9li1jVVhKKWMmJBpmYxtyni2tfXRRQ0naZxw4z7JCdTqdLLDpzYn3bHpdf
yJCczFR9T42ibkaJvzuf0RWce5+l+WJHpJ9Ie3J+6Wz1WkAzAAP6SGvWKXEBB53v
PDRH09miGwDcTblV2AQsuQZ6DDJDyxTPE+ACyJcnbWkkZcoCQ/G/4sEmEMSNUK+P
Ht4AKmUk87ARx4h9khAUzkzjTdtBFl98aiXWGnwMuC3DlqPNmemRYJbbR8l0h1Uv
wVpcKKMOme5lKK1Oz658vnZOEgRffB5U/c2skbGoDf1IE+b8StN+05YW3rMb0X3b
RBAS2evHjgiAZpU5TmuYCujbO6Z9p+Wwl1wlDYnp7mmUCgRSYoqtz1iPw3hDO+j8
6KvVyXVMiLQrg/JdJ7K7cjpYlTPc1kGsdxESP9uM2GY84tAaU/1uK/coC5ogVnFa
y7qktSJChgI2EhoCW7QNnhfrxzMOdNozFTbbfFEj1JpgWGdZ14UHsqVvwt8xs/J0
MubeQwUhiRSOON3DDpGfQLldpm2pMXSRMwRs4lmxaKgP9RnI+X02nal3R8kDDyiz
AkFASlt4g7BQZZSFYMYafZCKLSnWmPv2NmfKaVnBRKpoAFA3Yz2+bxvZHZNSzTAm
/0p3aEpoTueUjf5oI488CEwGU7YepecuAPT6ZSTFvh1BLKloVT9EaxjmrYkKVfAd
sK5WU6/BGBmsTRT1FNTksEmV1h4Gk0tm4tnN7Zs3AaqJi0gGSZSBv8RYaeLTjqr5
6hAOkq4l76BWrU90EnfiXG6bdQLQ735IxwMTGgeg9+Fk7OrJEGf2Y9SjEsV+KJeb
KC0cpTEqE3ix9jg41Lc6gMdcJEm36UZujzzSU29ZAn/m0QO9MYbrvpj6HMQhn7OS
BEn3o5BBExclNoLmzOtt4LgqajMoCTWxZ6cz85CO78DygXUHx9+/xt4b1gq1i+Iv
vwhao1S0Zu6OKG3FefoV70BxjQ/vUMg8Q77C9j+sA0vnafSPuZViG0T2uL3PAGlm
2sqsd1a3ObNrAOCkskfPHXhzUPiRLMIA8SgnPwGkK2whkDbavDeWUwz5I40qZm6J
BPo7SZdsXr89nzKB4q1G46OEzixloW67lGYi7XLZq7qvgRGU3sE0bg/VqgTlVZ2o
yVnKyuJ5iBTvjVCY3jyuskZQ1+sljzYRKodB7PswgTe+PZUOPuJitcioI1UhCbGx
xdB4iQGlk4qJMI6Ue/6ax3JVwv2qY3DB9NVvbVhJXytpUL1a0Q/QKUEo3iW1MAD3
rUYjcsMNwkGUMnlF/cNoliSr7WuT3Gy5fE1scUVE7PdNw5nRyOnmswz79nkYdZfD
NJRYdlyVyjioAvVYnEgXeFfq5sYnd5uW3YnWoHE1YE83vvRDrSZvNNrMFjvz3iG2
MxZ/QBs6s78e8pRrpr7OppPR5L2bMrh1a/+iab3zO6bRMxxW3YxCqdmuxML9YVcr
MuBCpWyO7ru7bS+UQnNo4X4Wf3dtmuVunYm51uldYxBbeAmn+SUilZ53q6GqRMvU
fdJREdi+giO/rWMOxmNT2qLcMsAJlCMtV842sLgPIjxzUPg82EC/WytXyO1qVHbB
3aIqEXmOcdr3xwxHclPL9XhKDLq+vy4WQK8LJqV3jn7M103ieW7JfaBg2D2/3BHR
5g1yClif3ircwBTWgCuHTM88OmcAofcQN51Up/F2YvE9XY8B19rOWRPXT9xs6BL7
JigjT8xPox45MU9ih4WsRFG0B2n7wmKuNWF/a3s/614Xf7RLgJFeRvrJgL6jSEkF
ebdaNnjO8QUFbj01PL9/e8wceXaXVesoTUZlgKqjGcf5qHg/5aE9j3KENVRvrUPp
AYJDs/RrPZs39wRSDjgZGBIwkLdHx+UpyOf2xsBiD3RYUH7/3nH+GzgBHesoq6fH
9UNmQfoq2A4/OrL+JO0fDERcTwH4KNpmcNpNOIzPuGP50LnM9mzgcHCiRhUSMVBm
lM9lkxwsfxGtou9tIb8ybIWkBZr4Ud17ygJH1Q5qu+8WmHh7b2J0XtzFpvqcolOr
WrYpeThO9cQDUFTFtTJNS/UzV4AuE0teKPnQdtwuSWGNe6JUhJDhimm7R9K0YPtW
9SAVBO4HW67CO0fTp8qM8KdDcgTscbgNJrjYUmxVwHjQEhnzBnij2350pw1dK13r
wne5qxesUMXf+rO9WIHgtQOv+rgZo2XfiDCXJvGisvh5zGCN8U/WosWmfNo0MDCN
AW0nTuv7Xs+Mdw5Tkkgms0wdKy6vSPuS+Kt5kKAB1xKiImm3gSlewc2DrZhYBcg5
2GfGUn+69XDtPrjXXTbwIwriY/L2ffL9Ymz6IkpMuL+m1sINMnX7eE5ErZKpypqR
f7GfxDCe23AOvPIHpYwHgFjHM7DmL0XQg5gloBKRWmJ7C9yXNqQdqttTOZDLMN75
F4/kvS9fOmed1UoUmJ61ch2Uev/aZbfo0lbxloq4Zs7diwXwpofJW/9aCumykmjq
QVUrzVP13RjZJooTNT+TaPjybh4zACKjaVdBMOeQR5robYFp4wfGAiLIvNTQiNOB
Ja86oMfDmuo33RBcl6ORVYIiieiHz+WwCN4ZtdmWiPOmNPn4q367XkpCSF5NddEe
tQ1dT75X1m43GNdGwRHZXAKU7BJuP2j3zvwAUZ92SysOJoQyhqbsM/Qzj+FIpmoV
DI9CLtfnzfZXzyo7sMAq5NaPGHMdophYwIROSUr3OIBKuAl+btNNiw7Ie5P6yo6M
D09q/EJ84HEV5cXNLcLBt2YCsx/Zw0cZwJUcgmDsOj1skDOhfrbWMNSPRS01ALoj
SijZYvxR2E3j0tAL71FydwtqVPtcvXBtGRGrB1P8KpDTy6fqqKPeHrshhY8pTGrc
wrw6iycluQm7djvq7oB4PMPibyW62moKwgLheWCFt1MlhT88Rsk2jl9oVkge6fFA
5ZJYej6cPHpFC3i4T3hLO8x25ej6EJolSHdi8w8kKqaFCe8O1Ko/GKsCyCqllHHI
SkbRrj8mbcn0bfGazF6vX8SnQ5ZyFAMDS8bLmEYCgD2BKnzQ43jq9kGpJo7209KF
Aj/NEU4yrZli5WmEI07/FpqBAG7xImQW6K9FW6+UT+4w/Tqyu/7TVffWa9q1Y1jl
/xTrahDsFKyGJ06h3yPZHi++NRK6GeBd/RR+UBdmTWquambt1kKGwIC/6i1PxSBD
fU2Vkjga0HTDExkbGTc4510/G5oAV6rTrDpD84qUEJ3M3Qef9i1ndXHSBy9CdKQP
aPKYx0cVNshOYs8OoUwAQFom6+E6MrINjd8NbHJsGfN9M7E466hiKWEVjCxgKWme
QCBCk/fbFotkDHmYEfYlzv/XHHVborS0LZOJf2VmZPnvDnpZ8iaHUin4jPrzLSn9
FonmQPNuEFcodKDcwYf2UUPmpFX/pzGZ0Xl/k5fn2gnizX76YZ9DOc5GgfkLpSGN
z8b9SkTlukdtylH8+HJmN0T0eJnOdH0WCQSowdrbDxcMVCIu6t3awTfG3Al9cIRq
BRzFSdnIFUFWKg42H6hmcJmcvhu5b5ZWrGICVrgxICdFp5mDIVnMFeOaAdkbGxod
8LRUjX6Xfnz2d0eHCYKj7ilBO3QLbq/Z7Kw7+B+DGlE+djd2t0UmyabOKsUlmMt+
OewCxN7NHuypN+N+f8BtfRo8X5OYcgjXuskIcYaE2yTZ9tdKjFLvY1snmKyIPPzE
6Tw6ERLTvKm8ktrWCOXDC8YM8fO5AqIpm6HB2HxZMvINcBWjkZwQ3QOJQOfeVYqr
N1vNjRvuufyPpd55UV7wE+kBigVw8N/gyl2bGHKG67H3Pg0hyiKZMfKc5V9ZrruY
CwW+IA1XtHabcjvrLg32tnRKS1IdH5uym8oANrbH1k2Jdx5sDlmYkxbGfTm1+oqd
0af35XcNbDt4+Arq30y3owLLb3nULrWho9XjJLVOTr/uYnQONeRNSgJZF2aCZGEG
Q0+TQLivrv2LYdYi3HnOYBWK/BTcGq3Jq7R5ABX10mkwE1Q480z7k5U3Vqw8TdDN
Ip7QBsHV4rTs5mbIos+W4PRef3bkBOqAdO+JqcR9/pmI8q9EskISR6SYoTObxTJm
d1O7ICTyBQSJjQZsnsop8FZv1WeFVUZLh80z0rBvUKBsE2sRRNFUBETUELkLEqTQ
J3YIePIrHnDSfvf3V6j72uwGQkuVkryPSKof9h0/xM5Peym2mfL8eLGhMEYp/X4j
nrxldaz93yBwpkCmGgEgVcx+nwocIVSmRP1Rw9eRLbK1tcF/0pMgmIqzyiwauyjl
9GVKPP3xxRn3HOu1ZiWeH1gyM/Hbj1ExwFej5Fi3iemalkksTFwtifHTO+Utvj7Z
8x5pNbU08twqMKib9Wsa9QskIEiBh6cTbs2miZtVR0efoxizMRkEdpeOBqN/GVxM
6cNQ4Ix7AitJI4JyOprtT3H54R87KF/j09eGeBI3w9cPfp1bOyhWEcVI3Hhio7zW
FNdO21tSsRGUdDgJskZoPUTPEf97arv0TmnnrQlXN975/D8KFThyEmv7Wc25yq8W
mxNdhjWNKd2JNZxDWu87m2lwdjAFIL1ErywWoDK1U0QnCnIwPswyWBp2annTqqBA
aORBigK5y1glczHF67X1tiDs4W9ksps8+7jMC8R+63JQKf2VcisD2mhXUB2x2Pxq
pE974wN5EoSVvo0sKxbIepl5cHZioenjeehSEGG57kC15adDIsbOwrHWMOsQwPs1
sCAyYhPDq7xVXW6IJGqArbokJIjqrVpfK/5uSDXp8GiMyCg3c0TEfiEQJEl8VJVs
jbTimfsgxxbM7Z9wK1d5lQY1eiOiBNBFpIrY+HuhFXZrs57MRvTU0sGlIAG3uBC7
6izvJQEQYMyPTyj75Qzo9ZHBTozf7+eD4V4oET6tL0zJYA3UoHntFUnG4askOgDr
G1XxJ+jDB+cdpxyfN3lbHPb0B69K2E/nxituZ0U+hCAY8u4rAFzzEgEhCnE0vltG
1kJXw+RTcBxGe3q7tCMuQ6AOW4JTsgbA4bWzA3Sr2PSzMzW48oKGAQfjrLxx2wHF
p0slZI3QyaBILkZRZPPIiACklVSjTzBsGliJfpT9haRFHa6Sh9y/BQKDeWLcrXpg
8/zZ4SlDHZ9n5Yhz/lKLIijbOEFfYRsLagCztxD+Da3zu4r/aUzf4joNTObhaWc/
RbngQuiOuLJCS5ZcgOZxD5646V8ijp8K8oWKCg6/Ejw5VVmhUQ2BO213jaA7QML5
UHLXrzbejSsNfNnrvjmTXRbD/iTftte44htf0JGH0F3RuPwYKxN6ks2uU9Of5ZVx
e+t7PUsYE+Z8T9BueyWIfxRiVQqOLWTm+YE/ZZd1CEZXWNmghnWBEjHLkhLgFRBe
UxOnhYpcAnbjJLdI8AzeM811Y1EFyYPd4vONiPHAlRwVnSlCMwtyiDP1Kb3Xnn+a
wj57iPA+GA93FJsPGRBfl58yNVh9o3+rLTsiVNBfqxumZAqoLwnQZHsQwCZwZUuV
wiAlb2B0U5lhEYaAVdGpmOPaZsnqxMdK1EuJaHX6ScBVT6HeefHYPsarz1Rnsgg3
FxvGdwT7IErqBMgNE+ATchY3PR2Ole9ds94lBMgWB1raBUYVVw9TyzEWyvfYT1g9
/GvHEGYcZsn0LWalriGPwg5a3SDHFHa+tZoSfLNr8N68XjXDWoEzn8PDsQYV4ETk
gH+m4IeX0TP3ihVNT7UdfE+F4Pi7ii01lSDT7yWQMtgz2nMdEMgKmF1JK6X0p7Tq
2ICfXl8x2XB3AZP2nVoc1Y3wHZKnzUjQQWGCV3SFyvFlWvyGD1ovIHXofOgBoX51
xAWjFrBSeGz46zXksZAT0QGglmPbKteyMZBBgFtboTzO0lAp+88oyMFk/IoprGxr
hH4NMPGQ82dmFo/2NGYrCBzHHWzFbjtWpd9RETc1u2tt6RVKetT7ck3K4aWUaLJI
xxdX4KDkON+AFzgK+rmGHkGXCecf48cC4m4Ul7Z9L8mOG9nXLAO7LZ9tJqfAWe70
I4UllhEW14yjJS+jlAQPMyp4VThiy5ek5pvlyV4jdxYEuSFKzGYLQ2k2tHk0O+xK
ijW6uYs3MunxJnZE+F0T/8e0Oj/k9aRWGHAW6Ki5hY56QRL9Oeo21SIyMWcWy7Mw
5tecXcInNkOgRaJDEGxWqcZFgWxjjBO0qeIqzeLI38xgSSdyi41FV7Lrvc0CbGrl
1CouJLbvN+Q13s+dRaui2CK8dLiXzW1nML8/b0XiMELzjl5f1y39ASsci6BTYZIV
IkCRmvpSSQc8gwL89kKImHWwPTsO0ilsccIYQdiddLQBRrE+S5OTbbBfS7Mfa9wP
JMZacZkeJIaw+vofydazw/WSoDk+Yu686wj65rtAYZHFqRIMQAiyDQGErMWjniGu
jcG59hA4pq14cSVXduHcyq2cuLrARNHbSwYqFj/zOTxb06gSoIyaXejQ/TAfRxF7
WCfaqDEbTPbXHrn2tGfODxvZIlgwkT4uFtgR3teI41IKZ707VPUbzHqVxbBHKtye
Cx4VFzqMAJzbb/8Vm5Juov9knGbrQpa1zCAAXb/nG/lzksqKra0ssrDDxRX6A6d/
ohmIhNNRy0+JpZ5OnkkNbc+uMt0Wn63FhH15EhUrdaglxcRHK322E2S0LAmrxBF0
fhBhYiLIhH1CgsQThWC0DKPdeL583krA4wgOisnuNbjU4NgaV0z4SzP1qynO+NWe
zXrP6ynHTcbwlWdsDiF8oWKSitIu/OooixHtG/vFz+flkNXzC28wQk8nFXRln+z+
+KrKwTiXTvDZRgpYOKBHeWwnTijWLXEAbj4a1lMVg2fqBl3bQCPloBNmfdd4ttAc
SvecnxSrbyVWexDtCU2xBfzgfKzzQSfQOwlacJPxa00uNiTZw5IbjNqIOoJ7Hsiz
bsTe/7Zqc58bCr47tECdOdxvPsa8CJIidJw7F+5uc+R+ZNMkDuCZVz8crYHWRGIu
2YxXUdlzU7cTYyotV5CBmBqBC44Ff3r+7DBINHhZZvvbiTbIXaClxfv1mZ8I3mfr
BJp6PE9hPyIODUUyiGnClFvfdl7eZp86sVHbvt659ycHUI86D7DbXPvEdLgCXXW8
rY+dcvuGJUW+9aVmPb+MJDpxuHs23LqQd8nGC7PhYov8D5+sGmo4CKjWPbI7LBq6
D1rSweqk730YA1NPef0piXePt6cksft35Oprrs9ia7jVOyAMTzdilgoRmvURJQsv
V+S0RhqSA5gvvDy6NkI0rLMm9G8+skZoFySxIuAryajgSxJhkCrWOcaPLpCq1Dlp
uo2A79NaFHR1z6dCQcSWbUgQPu3/HmlOS7gPwLNodxQaZAeBBtK6L3jQt0nO3zrJ
TZfbBklDrIFoe0wLz/qjyrocJuoVr7n41/Us+lvhHc2fieoXoriBozUR4n3skWD8
6PDaTJTj6B70/OkHRHj5W1O8wb3WNf6kZ6eZ5qVlIL9Tbp31veQ8S2bnIatnhbSR
A6gZowYnxMRXq/yXLJd7JUHXZu+4dEJc07ALwD+vN4enyDEcKwy+1/FduXhYevvn
c5VB4pxCNYHpKaOV/asMkcplGEVrO109gHCLBp7Cu9fgJw0IPo+PeZrVqVokxXJE
SXs9a2cnHRcTJObWnhZW7HR61GvTbML29ZsIR642fnNWGnocujnb2PUAuQoj1IyV
nEx5MTdfTssLxpumSzDMtIdqr00g70jsKLw913VwwvV5CsV6jCcmcYIMeR4RHT1h
z1Q0ldrO6WrrJ/NkqDhqQTFxCKq+ZgaB3uNWadll/N+hj7CLzMqGvHh9Q2gIwW4+
pvkGnHyp2FefTDT6BxdoXiwVk+YGpUdR4wFqWXToI9i1J+AYU92HBTLbYN5fqFQq
bROJpYVggGzrdusN/NKessT6ejSdxV4svZUMb2OftWDyM/sn3y8Q4qyEw0iUkTrs
Q/4Yhy8cyCA/4URwq2CojmwGqCpmtV3cUV1XjF1Zc8XFSMcpQCU0BAOSfIr3kpyf
vvKzfy+xvHHCv408fmqeS1Thu8psv5R5g5FVLxyOwiqOCk37eFBv6Bdf0Hj7G/Pt
1qs52ZOZIMk0SRlcJ6qCfFul4uo/Re0YX/0gEnafLbtSK7tkflRIWLnPvtx+UlKs
878kaJ+gAIve7py/E/3Vecp9zJkYTYCpJt69EIr5a1SQb8GkWPl2o+NtCvpVnjuU
2s5MfBspb8jkVOia+AsS7C44eY1q3pIF/2MR4kOEeRsyUyOgX/MMxhdxEwtMOYA9
a5pcX54ZHWJtWwRsxbEdMVby7KEL9fSyKLSo6bzPCi8BWNwbGfFxHMaT2jfgsJ2A
1XRsZ9qchbj88GP9cMQk0cZijDmoeAj+E8wbwA/a44lgiKepU2w4ZsMUndAoau0s
+wmGBzE/Sf7toeGpJDdybbbSb4R/eWJvzqRX447DyHFdzJQuXqgRBE5POCi8L8fM
7k34vX2u8hboB/ZiKpFJVZwFXFsKTXgl3XlYo71oRJk0wewUgXlM8sIoT89qWfT2
qk9mN0p+Zs0U2TPpu8jxt3owWrv4gA9ZGCVRh2oy2luL85zZ0AW738K+/5b70RDW
pof/sROb0U3stZrQSFldKPG6gFj8MfHWHhpUdZGIJXG5gfwc0U+19UecA3AUzH7Q
CwYQuB87zikhKRssHOt4Hl3LWVhL8OcQmkF/czCH9eBbpc9jShSmPWneW+J4I8PS
IE96pJz1SbOt9WRz2xZLpN3gWmOVW+qSsWmkwrsXL/6WyLimYuJ/0xoQNqC4uOAf
RiHnMjGFGzplTdS+2N3q88QHHSzFNxqZd+1CE6LGC5vtHq3ul9h+V3jQhtx9ktN1
nRhnEJhevtiQFiRC68BdLKlbv1kIrizUQPf30FXa8gqNP+4MGFivt9MROdohw8TR
rTVsHVhTwSBwqq9DKel6uYH3+99OWth3a1TJkQziV0154OsnZIttWUx1w6Z8ueiF
fi8Pn7JlP7UjWCs3MXX8qf4o/pTHa8lZkJHFvwyI2XQfmtBXs0WEMYGN8Z4DC0Fh
1kmcOXk5b4ace3UBZXftaDnFohA2UaPZ0MqYiC5eVd1F0IH/Jj2+xNcAZnvMqoD8
qZfyYdKhmSb8C60aV4r5aZ3b0T8VS1D9bQabYnlY27axebqUlrVWAs8MU/byJL85
j2Jed4GRc36De8vapBg+s5KjYz5UVTvXvj/dlxQOeU6L3laL59B7Lgos+8FZWlL9
8xCOUWAv+ls+pF628N9uT+2FqqphSGS7d1EpEDAX5q9rnssnWomzEjipOc0DSRgK
T11Xs/VynnzB1NU3OcS2VjcO6wwZtXp6iI7wEHfuqg4p9hCr0IEydQVf/ceT7uQn
czLB2H4CJ/466Wu8I4l1cfOZ/mOM9DupRn5I3bgDx3oBVe/rnk8FjUg97UmSLIGl
ww9cLnCWfskBACbpS9/qIL0q9DnL7pUvINdu9KHV7NFm1CR6U98e1WtCbCeb7NgA
sKDUvfWXeg3p9WUKj3Lhkol4S9m8J/WABFY3HMhY0YMNwZ/59Sf8s3QUzVDwjwDu
/qp1b9rVve3I3IEnv4bdMZ7I1rU/L605+Vmtzh09AN3/Ha5KRfj6z2d7mVL5dbTk
tkSahxRqzUeq1X5tF2aoXoq+iJugTIGznyzcgLU6Jac61fw4fxKC9cUVGlzmPpZK
qgxSGBTuXu2DfXtLNUJZEehDar3UC00115xBFeb6tQCwXl+S/0JqNmJ8o6gm3/mp
1fDpbD8M1m5cbsKAzCs97uDIVoxtAi71/JkIbHlNbKRg6TvvlNgorOjxdazLCNv4
fD7P2pgWbfx7ry3D1b+4cEw1F0yEhweCqXHnhCNrQuVpAiNbgnq09az7LhpnSnJS
ffmiV70173UYCXaPz/BfBFFfvkSapNg+qQVQOxzok/ftbJNmLCet8o5glyyNPUfU
2uii1DWw1nshZ+GvmdpLDQvj+o53FUHE9J476TAs/T918jh2HiYqb31XCxcASAZj
DvBhyQEBJ0GI3l89EkZxMLaIgJLOinWTQDTG/Xy2YYYYNSwNb+OACxtyDZaO5qdb
vrvWaDxrEov7dBeRMqAVMb0ZEO+GXzVK1ArowuxTg+XHm+vNmRG/EBab8rauggoE
k0DEFW7V6Yu24vtK6qsQTpiUWZzzVWtBoot90rKxQxnQvaPsTeDdiY5ZPPadczZl
anRjblL9P0IspUPALGkOEDxRcTtQOZcMwyZvAGT9DKT3gPltIlvsMWWReGtqfnLd
dU0k3i5WHgvQoyvSaOz/4jEP4uWxpGeL90P6LdB7LHMzJ9336nGj8b3FYamqsr/Z
bWwQ9hEe7do6wzt77TI0P8aaEGjrWm7onvuGw4lp5ADEOBOREqU6gmoEspdBnowD
mesLpodoU3iKOo4gJerc+pa/FeX0yF7t9wau7cGt0ixjWtFfNvzJ4cWEQQhEMLKH
qz9vVXJ60NMWsRmu2FxVz8EAmP4obngJrG9th1JGFhZzPfDF/khaDE6GUAcr9FaW
M++sEl2gYn1xRQ+o2Q0wik4JUZsaBd8blo8LWtpr7gL/QtkUN6r3vMeKL2rxLypS
Wu/LrF65ktOMHv8QLQuK58hD6fpRxlDQ8gVcv6ROngNsbBXU5A4IdV9/yJibxAEG
mV2K5FapSO4v4XFO8MQeuNA1N06FDfVBzQjrX6x+DFGKttjyiSr//JdaMmgBuLh2
OtG4WiP54Ij9S2DemycD+SaDgTCwrel8+y1VZ+SISIn7x1Oy83Z5UTrHTbvacJsK
e08EfjsRMqYJvhLLj2+fToCe1eWPqC2pJEqvkbU7QeNCbE9PhP1q1er62fLZTZfm
5+cSfMazMOyQSsLejxMGHhf5S48F3c1KvX+LfudTY+S1Ja622HMfPDMpWcUNQSvC
cCuci5irepyRImNelpa2+2X+iObX0Iitdo92bEt6v0KivuKVnsijEl0QrTXJC33K
K9k9RImbbJemeQ4hRlR9sjYxBzzzfbQ8Yl/HVP6sbwAtvzYENzt6TAT83siQqqCq
4kPEd/sRbWaPb2rtuyHTnTrefr62PlccwTHKrHHEQeMM/jvV+4kSRjOo4OArY0lo
I5oCYCxKkio9uQhEbfG9A/7kcDy1FCjHWIe7wrsRsIGtOG7SvgLf7o2lRvFZkJnX
QRNlhlnIQoeESaQra1CkeYKygk7ukivzXQv3z6SnvShmkSBRBLMSItuT09L1Nw1I
uY89T4J3Gd6FhzzgY1f1PcGRz4zfJO7PMvGpTlZWlubWTzLbeXtl1727VeHRe9GH
OIJ5+pZiaV4rgiXm59M9vKiwZrw7D4iXiNRQnM1ezwC3q1eqDYu2CvpDaL358z9s
6ea1LYl7CRDQzcwcN5QZmJ7VgR67KMcSK6foqMvOILRdHMqY/cdcKoDSf0kV21Kl
Vinxdtefu6rH3zU/5SW2F1ci3katUHIrIzJW4el2HlR9+Nyj/3C1TijHElwdH4oC
WAbYK+VZY5ryIi7k8B5JCj9JNyhv9TJnsc3PgjMj0VDM2bVn+fe1zCY8g5H0vBP5
7a9T65ZiH/4ZPFtv8aP2bco7nr21JUKgA3hyoMEz1hU9paXSKwgtPQ7oBQQ9GtaI
BfdkK1OrpyeoiRDydEKFUuwaGprBeLPkKF6spIPacpB99xwKrecysfqRwLbaVy+P
El6Gl6iisEGjTlaFUauOLGdNdfQvMt9AKqyjsjrIcdGFZUBbyRYMbeOO5I0uSmEe
11fZT+Lx2qUOfbBNl+O1YZ4ZcXnT26cVvSrlds3HingbZYLAZFCNZwxJkJ/YW5T6
9Y1TOSjXj90SoRYMtIOH9oE/g5lSBcWwJvaXnoLxjhbUiRCz9bCDGeQMlJtULKgw
NQZcih1qFfJb59toQ6Rcyq/S2JhvrScgdtvPZ6yavEHv5QmAAZgL0Oob1jkeoNqX
SHL0SByYhxZyZKrV3GNp+ufMxAAzwaM9hIATaTrFiiPJDV9q5wBXdFgpTSgtn7VJ
B9IySVFyK05RyxwmrsOqEP6X12tjXc1+9YYt2Uu+tazNgXwDrxW8oUp1xj+sYiPq
YizfkouidhG0kNyX28WhcWVUYsg6PpuGqpWju2ZlCQYU+W3U2iRUdfrWRAPDHtz+
l6eLY9Gi/k0aJwEmT+eDsG4CMCvbb41R42lNqlVLmV7PqoShAHxBfHtmaaQP9tbT
Xdaucdcju74g1LsvzZOGVcqfZnw4IsdHnptCXBxqP0+H6I0M1N6+hro6qm4kUKGm
VhUNd8e7kEt5FI7pRsONnulTje99uKBUpjhTGUcbpB5/7X7o6OvDuafmQ86M+bde
Ugp00R7lZm9F7IVVIsjyK7Sx/yi3ywsltK+CoXMv/Ks7jDQB7HRYQkUDEuFgd6mb
kUyQSaQQQoJQGjERmHQqWdlV93+YSIJHXGl00zp7UmNhAxsN19/KFSp+pkpOwbQz
/rtTBk9YK8CxrwKbYnD7skndoFq0HRgXrOmHk/JF9rRRwPFLHm0iUkn8qsvNjT5u
DRRqzQoXbGVtQamwxeDmPNY/EF/7QPM00rqwmHiNqvovswRMEqJXXuBHA9ZUFcdf
wOvfvO5Xd0gCEh/odXM/UQOQVR36Ia7xJzgnQwSJlRepd9iSMxhpgxK9LdBkn0os
tijo0ESW3jzJ/Y4LWAxuuQ4+XRA62LkyLNdgSwVr1y47nkP0Es61m1TP3oT2dUgN
eJ3Tpdnc9SkDGDBRV7yST1yfi7dwbLQCMOjJtC3jYof4iFeUg2sDUeJygwew27Oz
HXVR/yZGjCJChR4mQJXrgrn1w0UeEfy+0GPCelnHBZf3ZuT59T2nmFmswhmApcmk
DLa7dvDUJV667YrzrtzpbBcHuqaFAd4HndLsWvaWnOgqP0EZ4g4w3RbPggvS8ixO
Q+ctGoPJI+6Q1RFOYACCqKR5TO8XlFMQpI2Hmt7GAF9fJixW9TFtLGgTTIxm06gs
Ns85OCV3N3Nik/YJnYSDYsGUqYOwJHORqr5VW3SARZC1If9575amT+cGmBnIHTBh
KfD5gYPcZA879XXA0YMd870s5SNtOoeLeh53NtDv91szGFZzGkUJTyWb7YNpLrnf
wOQ7AAy/aNSb44zLolLGURYDVCZjnmrNCi+1Lk+y86FNZ9pc8w/K64hZM4bn/aze
vLBaTdbaaycEb5V/auqzMhh7dY5gS7JbRl64tPOxL/OHPtXr8XxvAf8V9DEcXMlg
0qASGBIuZRbg0Xp8A/Y6Qrf8QmNC85mv1gFdWh/ZQgPj6p2epVv+MX5tKvWGuflH
MlWfpJ7Kv96V8fVbz61/yz/JwA37LdYFAElE9Y9CqeMPY/NQIoCOjt8Wtt0k9Tcn
Ugwc10gAO3ygcQ+wHsgtBXr2a3/pEScp9PtjWIvF4uUMRM4pSphsgksgKg/ThiZP
bSbN0nCrXQJXhPpzzW+udOY8Z/OYxOhKHRly7Gt0EJs4Tgieht+3zBUfwLYeoYtt
UfOFq/EhpZcj/xS3Jqbgo+zK1CIFMcYB+DNdcd/O0porYajbU20R2QInORhBTbPU
FKV/4gnqEhQu1LGjKi0FnD2zt6AITxFn7b8XGHxIe2BeeSjFi/c1YVzwqiHjTx2z
eaDGXKW5HS5B37ZPrGhJ7h2E7Yw1lpQvvrQPn8U8BdWExsgx0/Oamtiz7D21un0v
zdw96AakaTTjwnyLEilQ8zafSjGr70EXqCJ51U3woeDaVj9jDODy7jP/3PerhKUi
wB1U3+HVH2etnVggCR3vIuYLWQcImww/T8FWS4ByWlMB1SLC5A+SEDrmhKSICJr2
7YLCwn02NzetZXP8o2lOlI3L02j/LzjjQ33bYbUfgFjVh5tJIcr3wX6wrpjmY93c
1wL6eXmmmXSFo31Fhr/P0rHlaZScEvq25xvVkguuNbbQ0RTS65DKSFKvLBCLDMRE
CDDQcl4mPHbCbIO8gZBszfW3lSUMmFGjWnhxrsrdjzhJrqo2vbqQeCNDAUy9g8+p
AgCyRMDhSu8TgOtBYQ8cFYgarGFBFmCqKg2lBT2bfD0EGtf+rRczwRMT2iZLs6jx
kOSrj8jDHfE+CgVl65Nu6YxQsiJNF0gEpxzkJtAzcOM79hiiMEsYxK+8FiceSuZ5
FTQOLdXCzk5cOkLetnWuzqcKzjeZrI/kLl36tR1PQaAyhePrnKuWkwFB0U4d6XOb
qlVItQZpi253GTWvoMZ+o0DzASpBG9cHzRc2XJOKEQNqCaqOaRElHIVRLP+TxCVB
yndxskHio/Q5HXMEkMDQbg+gOnK28rAf0fYLSHAtt6cdQQDQQedxnltttSatpWWp
0l1ZG4kOb1znoQWmCdvCcwc0I1zPyNzdWIz8g93qhNOrYnVQGrwqISVkgL3RhCwY
Piz4pwUg1HEq2QogykstWWmXJRftur07dtVTOdcPppnssmXmqlLGLkfH9HXnjk8i
nbzxZn4GPgZzWbg1Jnpfw7VJJDERHlzRxzzsGmjrUsv1yWSDxX5BjSyDOW+vUFMZ
GxY3jnxZjiKfOvFbTKzw50LOOgoV5MwnrNKk+Wlbqs1Z6rQLnHdGfMUiGOVplpVf
OvK+uL2Rcl8+O5vCYy0DYR1r7kXtJM9861YUucxmZdVrFtfDVt5MQlJBQ78zrn9a
EniqbgKhfGB1QzQuLFevSVy7qwqiltJPHvv6LxHM22cg4UOx8835+MpazPjYJ5Wu
9dPNmd8ROmURxULZTrXxuI5YJGiLpCR6owe6/VwZS5Xwv7MOAfX+6WUBgqLrO/uV
KbepXojcqhGkC6VBSKVtMv353sU1tZ+zthVos12ajFzJnGy7BfHXiFIrWYZcpeUL
MdGMe9Ibs77WQsO73pPEnYUXMEtzQIYbh0/iQo5nT539HNfgxwnimL5PNuPPi253
I/7bCZng+BCjwfL85Q8erIRHfFNYfiJPzIMReyWeOSdaZSlE/bYeZumE7IBdrHIF
u8t349lw+gDlmR4h+NUNLh9sCJUU7sAjKZwG9gr8k2HhoPmIzjkHtFwGacr1CeuE
AW7syeaHxa42W7DuidBXcjwTxC6ReKXH/2oqvloCeEkjQ4oMXb6HV3uj7b20zGCk
ExSnF65cKJZ2u5KnhCPwU185j2zbsl6ePBDqghQVGC3sq+vucbApzFaZSeewLqof
fA/wABGD+Ner7rh5CafS1Vic9h7l8h0oxuSgD3GAZDRNSyIwNliwnS0uJceq9UoL
aPMEu3EpUKeEwCjQejPRqrJQYAYugcnERKuSR6iJ9Jxc+Ktgttcq1BbQT0U6eMCf
vzgbmJxqemOa31+5fm5f2kHCJ8JSGxA7DRB5AHv5gQkHymBQknzI8L/Duk+6yMYK
mAWKQ3VzHLrsM8kG/w9SXwypXRUh5zRp7jEXjVSmCnjm0Xf6AETEoTaKf2E2Tfsi
A+5kaaMw2b+Psysyr26lfYjXPgDnQMXl+3/hA1bwGZiie2neiNLuY7na51Bzfi2G
wQotHgvu6llNUxcMiPyBFGgWI3lMWTIJ9bwOelaiRcH9O597qV5ZajMNsaFi6ySs
lrFEI/K/J989TM9ewrzGh3AUmvatJCaYCqpBSIy0+xOhtSCjptjVdMHXAkQOUsBk
HmQDsgtaBotlkAAtdvwORIUb8eEJhU4MrNQLYh2L4PWmyG6DOmKhKQk7NQQ/bxYC
CP1EpgMfEguWjUqOeMkH8vDn48QCmgmwJorOdC0hrQpcT4tYbmHSb6z/RYqwUVRm
KoLmzeRlK+hHD2vdWXK6gORryvzChXfWc6bnJ0GLo/yTAXm9ukbH4piXfjvQNdtu
6ZXnXJJyENqDDmwJRfGzH4Zq9mKeKMzNDJKOAwNS3ZDxUkx5CF4rBswzd5oh4SBE
gHcFdloVzp8NMGtvu5ebIAVS1DSvyMiOrVdfPhJai/i7MEWD9W+EZFCZzy+5DGxZ
BmJXoXKE0OGSjP6Q/xxASgThLPrEKe/lAR84FAk9BGgstfRUqcp8EOGxnyuU3jzU
z1yjhs6S8ap7VXkZl7TeHEm1UQZXic1QIUjTC10u2XQoRFWRrFb6Qopa4mjhwRid
GYfcEoUa0PvSwQySYbwodoHb9JEhEgMVJLxhRDWfhtonkB9/e/+yZZzODTbJ5Q8I
DSwSPaFBiTbqTCK3gvxW041LSDBlzvPbygd9zroeKluu03jT+dHQvFqQb0+lmfYo
hw914mYvQStLiCdB1UANpJnyrqeJWm5Sv+uLR3ojjBCbEz2dj3LzS0l2aizuXvlk
Ftik6xrrilrwVv0iAChHsFOA6hlxhKwqezM5UrsEGDWpUouIyKpPDb2uy8+3UkRk
ZXFI+eZFm8TcYR6Fj/6F4yyeftM3b7/ITw4FC8FuK+HXg2KlXGtDuFwg/W2KCcGa
rRqqjwCYgDGx5bBFQS+u3euQgjlpuxvUsnzIge5mFr5C3Xc2+PoMW+GJFTkS0GgK
PGqXOra6L9i6ap0LeBO6Mu44gvONzy+I9ZUdVYIVbiHB4N3YClKDRz5c8X4h9uQh
ZhxpB6dQsPDPQP1MJnvhIKxi5c7kZ+DxBezFZ24BkJyvsIoWUUSdcvjaLI+aRdVK
PPQb5Xc+ga1fBLH6P2QM88kCfmFG2z3Ns/qFgbrYG0Z31TrHa1/Sjon4+Itr04xI
F5W3GeRJabIOP693kt/9J0Re7MwZ0ZAGXZYMjguvLII5K8dbzOVEbR6KJVQsGKsQ
vGLfI+EfxwXOi5xy29EWHZo9utvlbxNOBx+HUafsQt+C6WqL9jlKCxwH9Q2EjVsk
yd728EnsEwZqL8Cp/o4U9C41i3XtY0j8ye6H8/C84VhqWchcy0chcPoANeAi9Nhd
3X3An0z67MOdbx6bkkpiEtPUMuYY/LYjRrm1mA9ViBv+htHYeQXd1YSA3+eevj77
4aeT/K6/34buv9FrbCL44PEvaOyh8ytBuzPKiB8U/l542rj9u5BBakBBMLyCINCo
6JGNePkGrmAoWVIq8h3si0wak3Ypac57by+z8cIIYQiP9pTlJQyDEscQZnRaikag
aQPIgWBjIXlEXoZ33agWuj4eqXVDEb6gnl4D7qf5orZZarK1VcCkuBqDhbIvouBB
qaUqDWzX+/NA2XgLHxJFOT6tcB3RPG5D1xA+wNDq3BJMS9hViOcJkCSZHuB7P2FU
FEXmHufJU3v2VA9NUA4qeoDHgfv6MW3ghhN6x2FxhV3PpC+XJXN3GyUV+uhz3SGV
TxxAZR2jt/cJAQ80kiIp8CWEDbipJxxvG/6eB7/kCXUvreyoEzURsfFVnVhElbL8
n6TkwgQC6mOM+9Q0V0k2zU8YKzAbIRBge+6k8yjTT5TUq4AlmVJcqYoEpOGLvhXg
6fP2yQcEXAYEqgqYzyDgQgkJAhXSkfBGI5HHfcIq15qatb33XiANMqqIu1jQNgzQ
KI58CeMPHTS9UbvgE7AQ0se/QwIdzPuCQXKE1z/YeY+WqkznhyAIalLi4YEVrCCU
VdywtBip/WzkE6vAlpFQxEuLUiMyH0fnmBXrWz6Y0CVXkJEJpXdkBGzCNBjOd/Mz
SBr2s/6ZorWWjtfLqPGt7UoSIKGhPhzmjz99C6bM/pGOVw8/KU6EdQTX82IOjQQm
a9TesugXyO/zvCOmJs3YMmF26q3ilMgSGca1+U7YKevHJJAvzL2t6LtRhV9E5bEy
9LJu2BIe0t7VngUD8cRj41WOL6uM9/QMfWwObK7qzIKmdGkq4PRue7HgYD1anCEq
BBQ8EZvLJSsGhcbLIN4elieWPcSEpfPuIcxGUhYVNxbMJhe7K4nHwPC/YEckVsRl
XjuXotWnsVJSAJ9CIGO9Eyo7kyW/5611zR4kE8gSUwiuPskak8ilScyFdHO00xPT
9Pt3pB8SRUcxR7VTESTemaQTqEgDZU9RDV2JECK+1CxeCpIdRiNdU1xGlmtZZAkY
if5EwOe2AmpYOu8Oi377Ut/sm3GKGVpoZLQT9qsQj3KLejQ3R+LIVMwNsxf8XWeH
kW92E1uMJ+Bdq0HMX3elS6lTIuFFr4SNubROKfbtkGEHA6Gjj/WhYB0V7wo3OJx4
RVAH2DNu5lakFwQc3/fKozxYB1wXOec2BV/NqgtHx1UqldHww/rDNf7OM7zE7zzv
HG2sFHBH67kixbZO2iBT59BXOLzkgoxz0WU14Q5v+wLjZ55KCvW/f0IteZTLDJIG
sSA31mlOhthjCNMOlL76UVjoTSpDbz6Aju+/kQCmVykUZHnX3yJpa6ved1XysaAu
jfoPTDN1EsZbFrl5LFFh6moI+f8/DoLMy2d2g0pFMAgaH74ThUcYWWR26JWB3zs3
HIS9sOC9on7N1/WlLf3bOWA3hkYTD59oLkTbgLCGcNqbtEpITtVJ1jw6ySxV+yw/
8kobPC3fyh3CxDirELN/mtE22nlm2hs7iXMRiJ7MMTPmRwxMV7MXUjEWMo/wBWxJ
VoqYUcovUD9CuJ+NHgVfL649wtphuvHRRBq9J+TIWAQylFx7b/Glc8kN9oiU99Ax
8zFjTwz8DikP/aOJbmYYedqpbO7XLkd1TPmaQkZ+WZ/TAR4sS7UxXlnrGkpD3hUm
R2EsEoI4/mGx+Son9kBOkc4s8WLXtql7Ja4By27zBuDxgDDPY87q9W6ASbMBkscP
iFQk+TxHWNK5toQtlsYiLHggODmpK2g/SaAegRFcA9bXgN5upc2htSjqs935PyH5
qnNGJ+oVXViPH0bwhO0UgYDuTJBO5Vs/4bFbquxRUPw8xkUP5jCZjJnZPaxl9QfV
8wkesydb2Fagq941P8P44Uv6WTlO+uSGFtPbK+KRLs3aIKGPKzHf+34UZBrdxKji
6OzLvQIpy5ql8A2Pq4rF6EDi0dZIaQR7/shZ1lIsL8yZCO9nBBA8UowkRrtDSdyu
yCz+Go4mSNPOMefA3/WWC/h6/qtAyoTf3l/3faPi6isrkindP42st0BETawzZfhv
Q9FJBhX+43RZetpR4JmWm2nbfZ67SQbqI2pZHLXRG5kloJ0tuGuBl8g4W4l1p3ys
fiK8GlV8+DXjBVLxace64WZTNkHWSSku2GJMsDgxHssR7RKjTWJHPu8ZefQ+6yqJ
d71wyg0Go1RN4t9DuL1gvbTcdCdlu7Fjx/xKQutJK6RthQ1TVmM3oIpkH+r8FPzr
tUF4W/vyMdY+JoQdkKA2KaSpVsMbeFlJVVpxdsiNRfMNCVXMUBM0ERUcX2NtiJ1/
Axg9eQ/sNRhVb8MfqIld4+zauooG1SlDAr8KFJtzPolgCc4vYc8LwCn6jfkqDmP4
ujh7s9L0QY4MOA9e5fDrUFm+ETrSsvz9Ldkl11gvUgc0X2CRLwkcgeFLB6sZDVkM
eJ6PLMeHcXaPFW4hz6DM5R90PXhkX/GCLYxUEW7fRiDXs8hg2aQjOQWkm/v8woV5
bd41C7u3no4ZHBCNtarIgm2sc5D3BojPpFYBrwiKblE7V0XtCAC9cFzs1W6ACl+L
3aapwNBecsT3pv294FkkjVSNfnfAT/GhluSAL1CwicaulDF/9Yc78SEo3ZvYvo7t
9mrtVV6zzEHnyDDypJaeHNcJuK7QcgeYlmd1xdYyIO9ZbRKdek+xfoeVc6QQFBrO
+J1ycDdagojI8F6Wj0+WiOULqp7PZY7Cs4ZBH6oitQaKzcEOWzN7yfiiAylXlrKC
HAoiA/1xkI2uDORl6EPQUtRuuOfeAm+jt15jjl4Ey8TU+ETWBtfFNcvBdTBZrYSJ
9VIcQmx3L2SqjqaMxB1mge/Pr/Vh5Wm1gG/sNnQlt1WFHNIecpJ9fKFB4EysAsmT
RiqEFu9rh4FTdCldcfjKJjPmxZzWG3vgxRw8dGXNLGTGqg3ZjaBfALZhGGJxBTIV
7kYPcWqcrYEEwOGiVWgFTawRN1+dndpWAX6a7AZ7MMfG4Xo/I/HMRwPEFKpjzaa+
g3lVn9+Rrx9A9Izp7CtWvrrHx4JlEznT8yAL3gR4hPqTpzytJcx9jRmEIplnLkwI
CxZ9NQZrN5FN/Bf/jXNUyfWCOI0P/WBlWIIeOuk+zSao6uTJH3O/8H6DCRPQyG+u
tnTeHEyPCUezG+ugM0ekr5FcDM5i591d4x1qz7O5OY7vPJuh2zT+RmzpmUsSAZZY
IM50fb+lI1y7NMP3UA/kUwMgQA9hfB+WUA8zFDh099FTOsEvr+EDi6xDn0rtLTDr
y5sFB27QbU5s30QCQoyvA/uoBLz9Dm6sb2JFQwuzMHSZ9lsvsGOGUAB8lvlnCVyn
S7tposs4ayhl4EbVoVW6AlBY1zUAaet+C8WpWT7Sq2puxTLA6A5DdbDOwo/HTHHr
sI0d1hD4Jq2+OTHp3UADlp6gq6OSRx8+Ddij8e+dwegKkOnhWMByg7lg6k8jkXzN
ODq8GNU7UxZQ5n1WJQr1wlqY2fcuqLOdr9uP3aa5sGn8oDyR2976LyBpeblwN0s2
c5avHGMaLgIYl5NdibBzXywP1dvqGVzk0/nTHsZvcasAJRoiMhQWJppvXQaRxhl/
aW/AJdl2BgqykHIyHsFUjeBBwETenFYeMxL6+r5RP4z2ZmeeSfrdqYPDArfuZk7h
2yDfbKQtas72UFSHtivo89rmBTGZkSzkvHIHkE5CF1Q7CMz+07Y9AR4LbVgwTsEs
uV1DEn+MlFn2DhitFVKXuYTkgVPc01Qzgko0Z+oh58PHYVQKR3iPd0BMAade4m7z
NEabHaRj0bwKjS6jFv7qBGvG8vUWIahXRMrYbsHxtvpoxzoyGdi/Ty3rUBLRqwcB
JorvAr7NddmxNNIQX1y8rveXvZXkbOVe1J0mOK1720O1riHTM83ckzVjsLIs4h8M
lzG7A2FZ6vAlm+Y0ZPEuyzl35NvGEnumwArlWDi7VZuLmUc4DNrAUJBkDtD3ZntX
diPzZz3p6QU4cyWqjXsmcoJTeJ88SBNv6tq6KnQUe4SJUc5vjg9Uw0EhLp8snoCc
t9ukb+ch8ZzKBmumW49dvVSJEqkQWSt5FCPgNddrMW6WIUB1Nf2x02VkQ1VXwofT
WkgGSYUgbm5hmDprk6bjjP0JRK7ICq303q/MSSnqRLkKyIZ5Oc+3x8O42ddbEU/S
BxssdcfqSgDgBpKsYuYjAFgaIXpI5RPr7mrrYZ18tbHRPWOzt9gfimqKGikxsShd
7UcrDVsQyB7J325olwfu4tlw5zfzFNNtWWgdbmaZQ0rw4XmDiZ7PMmdwk+6KcZfa
wQeu+/4bW2kopoLSEZc2jw9Cip680EYFn4pUDw9DBimGQcrgJnfvgUyh/SHNIjRD
ZSsfn5xp7hx2R7kALBQcU1MMYD/jPwvyv1hKKO0rsm+aQ+q0naTLgmZZgVUAnU37
wLp8XZYOGFDtQreARlxdDKT1H2vG3hCAM0V46t5nxfD92MbURiygjQ7w0fV6AQsI
JgWBczol1Snb+0SKwoy89veeyPfyCtJBjvVEfu6X8siI/mwjnLjw5vh0F0K6+wlN
G9gqinuGp3o65cvasefPOBUStXlItPe3+tjWUJW81PShtzeerkwe2zRCpm1OAXks
j9R61u0sLXefB3sQjmR5dTZUEHN6Nkz8PAG+LKxSW/4a3HJxviB9ps+75CXMSrMQ
Y0If5oQ7IDyLzVFr60HaWM+tX9UHdhacAQ3doiuffbT41S2+BDqlOG1RGoWtpb5u
op8JpJmvMGd1xMzQjDsFjN3JIEwdTY4c6aWUrbroJv2zD+jfTLSo9iT47v2/imcZ
gX9EzAmQcQ+X4wDawVx2/NYubehoy7HjbKJOnpHGOffbYJNl6Nnw7o/5bs/RdcDY
5u3nm4OAzAhvk+wvi6lORwRnW86p5/ePaF16K4/+o2Fdq2maFPd41mUhDYxASsjl
jXngE98GKqC2QGSmWPsAJ8vcjluynLJeJcXC5Td9XLUDXC1jeePYNcjT3RJj/cwb
dpIr7LNKoAN1g80v9NrzG0ZgWhQ+uvOJnIA5eGd9ByNrTI88zj1TIofg6pfwqCBG
CAMH/zD374Skh/R5bCjjXKtuLdECNlNI0RkXP9Y/czA2Bf/w0HRCXpUiK5VsRpML
UnFlQXReLXLFHiLOpWJrGKWas6ZtHSpVLvvmZ5tEPzhewiB3XTZlziAegdMYeyDM
0s5s1jDrJWzrmH0KM2hnPLuqz/bOWiihFsUMCY3xBw/N3eJ2JZZ2hRBFmSpy3Vu0
uBLOtcdcXBma+NyzThjiPZdQsiRyvq3mDbtjAbunuYyqMBygij7GOSHz8e2dLqoG
6TUzLmmjEMyRTG39CWI01e8yculbrNiLPLiZDrsSLo4ByytpkdasuFLjiN8MIu1t
iiqEuooCeMEaEzImdgzec+dCv++BggFHZxQ++mtNlthbNmS/2HZei08UCPvy7O41
hYACJoYvdMEV1LvTP/p3PdCIZg8c0GViDUQkes3ctJEwdGUeGbdLiV/f2UO1hgvI
9V5x+C9a+nVpeKEJbtrSBdzZOzhE3vcJopcp/B2rTof/5/vkgw6brcWmOfXm4neN
avbcH9tjiqJanECLFaoV9MAiAxs48d/5/RcWJH8wK7GLJgl8x9Pse/K7kyEyn7FU
sx3nFJaVhAC7BHt3RZSQlAWNr7esohHt8IJOIH+lpgF2u4D9x6QFuCRfEbfoIGsk
VQ9FtM8x3i/rGV8Y/OEEndj5yTxqtDtXhyQDVlzNQCFMHbJjLUh32fYjWhnJi06C
lURq8m7jwrwhsaIiJuF1jjvx1WCJHfGqFOdXXrEEjVjQYWDhgFcjJ1xkvCMQgHwr
BeHy0YKFMEKvsu7Gi+CphC/kBfKGVe9fzWR1/pex4pt6NbOGw7L5/T19/R5uoXAN
Mj9XBZFVTvz+JUD58BtEgV0YIGrRi/TkTU1ru9KC715kvY+DyfPrdxyF8ix3lLEQ
QGVplX4PrZQHxpLVhYiMfi3UC2B2QLjDL5s0nc+Tbm3mUHvDlpWzX2aKpIqvqrcX
gLebbtip4DqaVJhDWyNGeg/rGpOZWwDcDbpbg4zIFBFfbQsyQTN/e1DM4cFKMjBL
rBdRh97mPuXfnrI6vGONVcbGBBcuhXB9smc32Rm0ZAKFOSK3LOT/CdRCLkT+4VKV
tok0g29ys9nO4qHieSU+ODp992V4jkvOit/yVne3KE3AlzKIORYQlcuqvti0lOFC
EwnGGyTdWKblxxw6kW7TxcgPUBUK3ErhxJCup3/oeYYAzVntL4/DOBR+30+zpgCi
jc2IGMuLf4TT12OudAOmIUp+VAXidndSWFtxMduGHJWDIEYVwUFv6MfRj4kiUwIo
K8zChLrW6Mwu2ECa+DXPE/23/Gt80y2za6rMFcQL03z/aBITXYdAK+LGs7CRrMEN
a23G2eATkK0oTVk2UCqX6G/LXahUn/EK820QVT/QNwQojlKVTEtIUTTirk/7XssK
UK0tGV/B7V5kP2C6aCCj8FvIS+Nsp3coAiKVX67XuirTvZywxHnE2T+8JKs4aaTj
NsfS3ELVgXMlSyJAHfpIyPtOwOfpMwEa1O4ZHgVbIdrVOEQpQ7bLlplHKCsX31mn
iceX9PNM+iuWYBuN/k/7YTfc07Y/dTB5b4fWcSxVzaKLyhwuDntr/CQsITZ0s9Ff
crQtpuX+BGCEMqEyhheW7DsQsuVvco5lQOlPA8sO81/qte//JZroeIwloOlK5Fm4
WEEoQCXJStHKFatokGZT+hj/5TEL6yELwBdplwlxf8YJlWDIDnJEhHO1JpsgoqHI
203KAUd+ZK3VQDo/Oqc5wkavuYJnA3MN9bWLNe0idzIWnly2kMytTI0vOQne691B
7WLMBGjQ3fQWV1tzziksfazN5i6cGNnouPGBtiA2Ni4LyY9sWQgepf/1vXNr1zML
SepWr2I5zRSMmp+iFfsQFDRf7advjEUflvsJ5xFdH28xgtZ5DC8mpurtxKQjDMAD
OYRr901bX62uQbX3sspt2OqMUJ+My+9n/oQHAPh9Q2kYpcO/6txhUvQbUgvaCUly
jrm1LVnhBNKro6+k47gRUjGOF1UNGuP5WO0r1xTSfIo9/Gtxh4pqqf6toL7OoobZ
xuuEejXrGd8h5H7xXX6FIaXvrvlv558R3aOfqmmL1NuZkwMtM+VGbUNo0hhjHZOP
jwhfsgRD/1ht/a8TKX8GcdbNECzo5t3CFmGb5IknKNKUG4myx/XPL+t520ql9kW3
Gd5b/4TY5rEJwpVRsSR8r5deLf8SiLkgYbyi28syuL4wla3qSyYskWvj93kwcqBC
j+hkBKv9Pgik9sFrIswYwQDVlSw6d7S3MZAA/zBxLbHkWh1NLWwE/ITxr1LX+H1K
gxz04TBqc0XxM5HjOEshB09BF09559IjloVQIEK0R1+livV7dPXrmisOP0oDdf/N
MVNYtZ/rX0XbjgeOAcXv2D1MoNhDx9EsvT5PW+dThFYjff4oTIiRYF/ORzx6YGsE
5SMfQihzXxEvG/L9suzj9sDf3UPdL4UAMVZUY3ihQulUWBOiKZb1kq06aMvg4MX7
6UqqudrLk1cXA4Xi0aCr+zTzvU5lByfxEn/BJZdjMN0qOdPCSihBlDnoISQhyTCc
UHea9Ub0dREAfaUYEBCQ5qLuolD2mwbHhQjpEIEKESrYczmpCbVqmMgCESExAasA
bRGXdSt3YvYoDlW6vO/+hEJeC5FeGCswLpdnem0fNjYvAyi42CP1gSoCu6/Nqekj
QfQnHC6Il8pBPPMWoQ1eH3NVeDWycFBr836VoRlGmfuxfqN/RqRYg1Iub69DugaK
FuoGG88La3MuWtd9RdkS9WMplmsmfL1b/HGvO+5j0LcpzSaLLYEhCvHKsnlaRsnS
slAU2XrJALfLJfundSlXVKms+w2VFNwRvHmE8Ewpu4n8GHjZx8YXLPj4oIF812wg
MDnA2IDj04sFXKZLcnA1BgLuLD4tKrKq8rZFQR/ZX8hO/45f8ogwooPpP8toDa2z
mJXjUeimZ1AnAim3U66tDJzWRxws7Gz7GHEM6ujp2A/75coWj8gGPJD96uqXk2Td
OC6cQTFrqdAkf4mxYbbt9XYjU4wKic/4Nc8rTmsVJIDiHxSSaMmmyQYA97xR0L/h
+bugMqKwgJXMKF07EhDPP0QePHbMzqC1DVkxsahF3SZd+29ZaSdDSGJxZa3eRCE6
h0j/0zZdGl0M8fQYA7GNPllo4Vfj8hsSI4MQ8xf24e4m9UT0wX7Uj+9nIttFroyl
ZSzkXU97L4ijF+Y+jMSq8H8hG9RCWI/WhbwfAv1kmJZ0r0aHDbU/7FyZA8O1LV5M
iFLPUlkho3fchJarRxoqR2O3aZbKi2N878WiQ6K1W/T9cS1CaCee1GuQn6qtCvZs
ks4gTf+Ei0saojKl1BMy8jl+BFdJ+01O2ZOi7lotQdB3z7HvCO19q1vkhGRqqEPh
cL0mF2ntdj/IW16kSu5Ll2VCjAq0HRlvqTZJrVbx7yFyXra17SnNkVxCjyGL02g7
8fYV2IsyKzyv1C4OgiD5ZxtAP2wRxeH7qPaL+EWTcSfTw+YTWd9Xsrp4V75yeUvD
pmWVJuecZvzFv5MBX+YFdtYEJ9zYQCTklVxTqCcgX34VuHlZOt0mJwBP5Npujqdp
bLsuPW97+xZF5OT40o/33r/5kR3EkbEQxDbUqREPtMP1fOWvNZ0NryrTc0GjNZmI
p+sW1n/O0pyfyfYIGkw6OaLrKZkTgMFVMEPitmsjAWh4uc/iJK8lmYVHiILhAnH0
wOjGWRK64NS/nOKjZZ0FaYWdS7OnV2qyNEIqGRJv8PJtGydDITsrQY5be3P8ljOb
OWy0TgK5UWKe2mk4yeT/vc0iMulUk+5gSCCi33T/q/DmzRTdIo2a4hoNajqZbuDs
dmbMQ6302smo7x2InQLRinhjabtG1yGubhMq5D9ciOa6CuusJeQsOMiNtluRHPN+
1Gar8Xa/wvk66LKCSvWKpw3aWkMi9KPOp64R5NAxwj/22HNNr3qvH1pvTHflvheR
dAT2UykNcqOwxwybPkCBvp2vXkeA2afmlbK2MYTSif1Gpm0EtVlyEFhLw1uvGpPp
6lM46pfSWXoLEnE6juXsf/NhuyNHttoOKyW59H/iIXXw5CybU0Ztw9OrPHDEcHiK
x1pf6CRm7FJtA9Y3DoIDfQh62s2gbEPvfPd0MyHaaNE0o/TwEhejWHuQJbdNWFlp
dG/8pNQQs64a4UPsp+Duj0ANH9oCd/NoLR8parRBtE3ACzWMVA9v7mSC/g0toERk
jl+u/F1Nb92/Le6ZqkCOFxnSt49IVRM+c05cio8uUgThhpmZFN6LFU4M3+v6o2If
Jpt1pgii6WiZTN6Rs2rwlM60HHsfOCeiv22aH8lPsNeDF1BHE8jrD9kuonRHRRt2
MRjI/lTQ18QUpd/JJu/iPTQ6f+IEw9QxrG9mS7JRle29cr/H4Y8ktiPTo646iy24
LxtvAnZMDiOV+DWKtU1JRQ4wxCQ5jem/b0E7zHoYwiBxKitErZLNz2CWbijiAZfU
MfiHBr9k760NXrC4ykTpTcWWm6Wc0eZ91BghkUQh0/Xzl7mKF2p7fyif+TDfyuS/
DZ1Ixxwad3VpYQyEnUd++6/ImoSzIqxxliY2/dQ5h0BBJWZlUGfMSIvUPsqIYaqa
j8ctQMrHdJm29450YhOnFHznCpxZyT7mjpPeOcORSS2lXYko+1ITWeg8fN3HsY4Z
s15qGmHWWhXHboZRJ2HN99pPCIoiMx6Jci+0DkA2dWU2wSflMOJuLCgpRHOJ0F5n
cp1yjfgChB7cL7gCXrnV9SrjEB1ghX4Oyelf5xraDrkS99R/GaYD7Q9536T7KNxN
xNpaduGYHROlzBVm/97ueqIBImTq55bFB1I6MvR51K+kvBUzPnJj5bTl8QNJzWtY
FudblQfG0KIhPXyT4nWIdOWLeTLUJ3oO4l4DouwOBGnlW9Rp9ruAlLq0/SAHhqSG
Be1R1p+AikEaItLebnUtuS9z1hOWWkeRuB8x2ZyjEz5w0YTlDggmVLYum7RyYwvR
+ZpTlS2CEie1fyGt4tWL6QINU0L3vy4E+9mYEent4kBZrH4//lxVzUPY2sKdKdsH
JsPmswfdWZdTkkDULPTNOwZEAIZpfCBbTEImPhKBrrH6knnqxOUviD1ra/+WpNFN
o2YFlFURAKgJy6oNgiwS3SJ1iZAOSVIJUSz+vAVteXc3Db+QOgoGFpnjzhLXur+k
nHlbV5kkjXIdlDaT5WOo5l+705fufCOIB4QXR4V9BSTpMWGJlPjw7o7Ynr2cG5qj
7JLFyPXPhMTkwClGeiQvMo6r2aUyvUoIxmBxSuEDXO1RoCvXQD0AeIV/4AyOrx4B
sqvazXr805IVMoiFd+JrWWS+Du2Mk1dTaTDlHZ0M6iU5VfECZhzHdPwkogDVH1aE
oHyUxT+uc+E6iCGuQrfa2zjti+8UIQDPaDE5ypzjJZMZ7eecArL/SU56hL4s1OWw
88QZE3u4LcrVZUqWIB4uGA3oKrYEoqiF0glzlgqA4KAme/myjLBr7/AXk4MU5rOd
kIB1lziAWKT+ASX1DuQDtyMTndEXL/9gWMwy2k2mI8Mu+AQEpUM05J6nLQNMLdnE
CYOxTU+b6flWcmXQlaMqz5Q9MZCqvHG+ObLwrAaeMUR8HxjCB++y/DxQkHkVEp9t
KA1VcniOnjl+piH3KSiUXUcBHlGhLQ2vUCzwyiu6s8d04W7YbUK5NP/AP6c657jA
a5e06qBVVb3NnNLOVfeHjYia736FsazwOwaHM7I4kAT4wPWrmTnVVDW9e66pidaW
Bp18kT3ZypjnS15xPB50iMccUCNWvtdmRcBq6LkZhmBW/IoRL56kOSYJDZf720MK
bmXRm41aAn1zejSNRaDfdrtEROV3qJh4dlAjgY5pYNrDbY0KUSoH/yA0P1b+foK+
RwLkGTCebfhMOxg235ac6m3a431A6LapAiTGO5y/89/JX5lf+k4lwpwZsqdQInjF
FcfJvgmKy4iXHFU3NMX/1RENI8SuH32YLBWCJmlqDA4jE2JPGrpUR9j02RjEGnTI
UxA8ybf1gk1Q+GgIC/KXP21ZENTcCUZPCf4oWzi80JcyM0zhXG5RGbZbdl27NQrr
PsrhjZbsKzy61gCrNMoaB5BjmLXffyMvmW00wxMyO7qg3QrU8YU/1Z6fU9attREa
GvZp+eJS3KvBAFGUbi0Fenm6madq8HWhcVYIIkNHjv3brKvadqLDxxfKhY4V7Jkc
Fh5n32wOjim6xTMC7BJt+EvxYUF6ipvJOmgfNKYpXTX9ujA1e07M+22uCCHIach6
bCC7LOYVXKWvWAyt5UFT0QnQM35GEA1QR0VdkCHW1qEUX4n+zRyeq17mh+P4TsE/
Y/jNQOcHaAHZHezC/x4fB1f+Y18wsbgZg20xEIizbVFHfhpveoJGHJhNSBl38um1
EmSh4QUdubOiQoLdFpkxQupyOwkwJGPyRQkYkoPHvdfXm8NNCBCajDeezGp4z3DT
W3rl0xBLum5BfVdjz2g0zR+USp0qnqlVbMjZc/1d87UiefvqqHYgHzDv2Vl/SntA
GPowhTc9AokC7rd+4Bvw/AK2qpCm2uIcBBUPazl6eI6z5smTA2G0SJ/Viwe4BLuV
x8NxzQ+dRrSZiKOUU4gVpt4JTQNwf4mEMraOGcsbcWnbd702nCxuoOr85jp8eK/K
c3//UTNaPqJJmELUJlF965VI6Tc3mz8Svyy5a0EzlV/pAeaIez5mdEJ9cFIfhde8
yqSShDQUck8sbhP9C+uWe+CuDOs7VBeOskUIHtOP5UDxyVlOnNcmNbNO0VJs9mh1
hCDrV9uPtKrk4kF5ouFO65h78JrE9/C6u7wgYU9/uwtk2kI4knk/T+62sE+cE3kc
upOI1lbi73sjXnNlrowijkt2JpbnDLYoM7xO0Fdos2RyzZOvCitZwUmz6KdZJxb9
WA/xe2VU7gqXp1fVHCh7tbANBJQV/LdOzxt18kBNWHkdFvZOwtgydtGCqOP7idrX
e/TS6H8oWdRPcR5rB1YGiPGemBUxi82UjSdxdx3XSzYtk4RRJs1ylv3ayEIpQ5aH
9yQX4AiPrXsMGQv0zk+KA+YnwwTNzu4f+rClnEECY0Z9egL7/PwTC9BHOXUcxyif
bD75URAFQQqW2cRHZrsd82MlJyIuxWW4Vw2NTHk9fVdMPSbzyO2May4wodR/vaYo
s0s3nfAdTKILD/JtC24tXADnnBTPx97emO6atbXIZ3HmCtPo1NTG4Vk0kqcx9cCh
svxZGJ01+kOms75DzZ6ltZTJ0+aBGK4cYyxI1hN7nGjSvbbNrProx+k9npJ29mwu
gldpFdeppAIB0YiZVhIttZ4Dz4/2+c3EMV3gjEZCyhXSkHWF5utB8K/d5jlx/qkh
N+XjPIm0NFj5rkzXIbDRMzH+uWRoi9S6rjGj+N2skq7JbbPTtsHU+aB/d4fCYN3E
ghvlQ8cawaKhSSgifrcm5zBap8OaQy9Mt7QafKF8Wv0SI2LdMc3P3UoWbcMr5y7o
2FrSqPpho45kX2kyU9j7lkrkDG+IwHN1xAzhzO84JTTQVqWzs1xBxENpcqXDdDbK
+P1BD5MVjF6Mi4noSIwSG3lcVfVlUqv0zXY77Hcl6iCbYp2NqoEeTSjTamCU8VuS
pYzniEuCqe0kNpp9/k765xqupq2xW0e2BpqRzjh8OLZWona2ZuFt4NBB4depytvP
ge8Hgaw/pdboIB51VRmYbx593bpoGg8BasMEyf+9Maip3U48b5pI28Ox08e/oXIS
V9on9U6h/vlR9clGg9skX9xK8Ffvulej5sAgJGF1dxKqbBHxhQGGCMsGmz/655pq
q4jbaKd9nww3HnyaZ6in33eSyNLbrE7LQTZ54FiXEEEGkYe39YVHhpf9buzdLLzu
pjQO0EIG90RZy9Q1HdV+P1mylSzQqmL9ebuEn3Js2qk+QElZIz+hnG4ijU/H8eK6
CJbLM/5Hfa1ehwgaDoOqN4Jb2sOEPo0O6DvybXIhd1ZZydVBLPriiddM7kb2AIFz
ntHLZbnuY/SfOlHK89uO5B8k9MuO3s47jl11BQsg5heaGmJGKPpKzL8XsQYFYXzm
gHZGgE408i/FbeRvFzH5xLyRdGwvSgoURYV39l/MzPdjoEovxVUh32YW6fCO49yB
6Qi/n0uW1z78TD5zif4nfruK2OR9D1s0owkkxUuE9YBkys3Yn2TKCNAtFsNZfYBR
E4j0hreZdHpJklRdVgFuvqEfzULkRvH1y4b4iZnSgWUMzQPuAmWQNWLtdTfQLjsu
ElToUlACr0vSFGhpMdlDiDscNT+aGGoiJ5lOMCbggQt5sQG49YzC2emcn9+hrzC5
5MzVCUQl87lIiRjQZwxo09ibz4bgW4mkqKgi5O5X2HbBduPwp+bzdn765BN4aJqt
zMxuIHZBKTqlo3RsI1mUVJpylOkzU60B4oGTxhQBXAjaCfiXUbUQ27bJKOtbYbiB
F/wsyiyktcCckg8NnrPSQwy0N90euF3u31ZlM8pbdcfbKE4UFiNirmoONaGj2oKQ
8hxoPAYl0N0k4Jm0iMjVYV/zLeK5nu6qWDuZX2WwbCbzjJOsNtnhxPP2mlhmedIM
AF+psa0xwcvoXh8a6/N1DfQBayR+doy8YMsJdrFsu7uU6+i7iIL4+SOUHtjkkxyv
PhrrcnJcoLeAY2tXI2yycuxB9i6oa1rRSw9GR2o79QTc/Z6K6iaqLF6kkv+tV45+
R4DA8/ltTZat32G0UV5blwYL0oF8lILlRfC+MoNx+Y9QvsqxIwZbhyS/nNUv/vLG
FBN9IBsDxI+av9d1pVv4WgxjTOoc9OHubb+v7zjV6PY7PKiWAtPhy3zKU+8X1ZEP
3rY6Ubw2P0l29j/NJBLorkq9zovnrjTRsG4tgIHmUUesj/bcuc6JII21tjQZ0BHg
5Y3sh+VQKJnbTzOFp4xAWvbwDFrJhrFJNf2Y/EMYp7KakPqNqu2gRISBwzCrfZpy
qJDNp11fkKya1FcuJqqQXWktlVm0ETxDhN/s4Bt7BxAFNnRTQwjm7w1Sf1CC6OhQ
+mD5vLL83nb4mri+bXn9hzs4DKjHWNDRrv3CaX6TJrPgKVRjnCPqPI8bot1OLkx1
tPz8xo8waoBsypjXJwtOArw9hWB470NUx6kV+WS5OLSz8qCbgif/P0YenAfKKAyD
HWklsTSYyeQc9qEeAgRL9dkE9qVp0qvSH6hVcGiJYV8QFZE32Bt2ojvT4Hz8mSV+
DhhOW88N5VhfGL8U/nw39T+R5K0ZevP+E+1LHwJqRby3Z9D6N+CbMurA1t4yd8eh
jrgBkCxRTMsf4GrYLsmby70CMqiuhwHXb/sxfKMaxC8L6NosGLmXFIdk1fOhOpsl
NtmO/omHflQFzuR6LcMObRg6OcUM4IyVLX+E/Otn9ovtjvTSs1z3VPuq8HmSUXy+
HoDqns0HRYBpPH5/bzgmi9YqLQr9c2mxx6zTTeA5V0o6Hi6yJyfkJtucxpLKAWcU
5t95FcdbGL74td5yKzKB5AJwOREhyXPJBQBKO6ZqlPy9uBbTlAasc+TgDoN4rptD
+gsO4qLbFBf8JRatktH0c4PFHwsPni0EiOfq9WpNjeYAwcarb6E1bgp0qjj0rHjO
+/Kl+dnZjfzr1j+sSb0YiSQYi9dwVMTYWqgQ9FUf0dmMX2Jvt7C9ezix9j5ROqEW
MqsUc6A6WWxzI3LrhIv/5rE/037iugNMujFpP8yxXyI9qLvTQuy7cp2VaPu4ce+t
6+VfVc5qqh6rj8t2uANHZQHyvEgT1Lq6s1uJ8qXPSIrhDhRgjNqiE8yn+3Xl9+iR
/izdKSPpvQ2kpAlL+HmdN03fNr22WJ1HQUUnyf4lfz6vxC8OdWREn8yGeLSapZzR
4vlsb2W14vcPnG0bVrp2MLMqaoYbK1Z9yqC1E1Zd2jjih+Y2GkNYQIMC+syGK8vC
ZXp7AAjERIZOCRM+DSaYai0d0oYoNtxnXCXrVnDqWNIS9oATtokwvt5tAQI5+1pf
CtwNOW5/v3XNkK1bxxmbIRMSLhJdU9Rv3Sv1ntFn4CgV6Hj+caxtV1ADsphqxU5w
OnLs/ni25mYNWuE2xpXb9SbUxC8Vh2Q7B3E+mLprJ0n1rvDBaR5h5RgEyI3K+uUa
2f8rcakDmawy9Ad/cJkm3fRbjhyBSjWtmUEvMIi+V++qN8DQW5Cx6+JfNE0KPx3F
xM5ajtZyX3Yi45gZIj2B/K4peEEGvFnS7oFTz1ZdJlFvfz562ZqVdyGRWRAozA5F
rRaeg26sXBRGtRwqmrhZcPiFAsOih3ZjLdmvcykoor6Tre3Pfy+d1XrM22OwRzoy
bWb9q+1JSvH6TGfrT0Z/3dp8YLA8cRW5GNNk82A1T0k4kupdbqPplpmxw2LWesYa
CCzy50mIvo8ggjBxSKOj69j+XmhstugkF7EXAnhjrVih+HHEKxjBzzInp/4Pld3+
U1XYctHfeTIKjSg91G1CmlCHDFI0N1qUWKQqoynfrXAmYa89DkFZ17hWh9kN3Xv0
OHLOXiNZ7nKSsbB8YsH7sQp2XpzK06i/1wuZZ2qa2z7WRKKC5cJMWvjt3XZFfpxo
1zRkayLk+Z8eW/iHRdSULGfrTlLar3FM7FIw1vzt7zwBtb+4WWWfV+jIMPpUCLR4
eyrMGSquXuBfhY66quRoRnnPPkAzhZlQDfhIocXlATLsdHLwM3T5jMnCweCrLNHN
nq2LAHrmWS33AfF4F519xQIAmh+xE2/Zon/p4OTmdiZE3+/uE5Gded9l6ClKqGyz
lKBufuF7MPwoNJcZBLB50X4pZvzDPTuxJi8/f+C6Y1Zx23zxvNPumLT5NPUCkeyk
Du9h6yX1pJwfvRqmWp5e3duTfxpw5hc86oldklC1G46qB7TOZ6BLJINgVThoKkzo
wJyCrdzg42rczti02wNhB1ELLxKL3DgyY5gIRtkR3xZ6TmF5Ko1HYAOM4GePIAqr
SrelDRy+nJioZstpjOp7MIp2w46DPqqloYZdolndqpPcMlJKe/J5inhok3HsQuha
cMzdK8J/I/ZzzankXuVzUunGkoSJJTPWe5NXUyPhJOkJBOANVH2ZfF5QCZTQj8xG
yZDxVLP2v8nA0k7QG6VUbBdr00BMFkSZ1ZT0DY2iVyoEhqh9VKcPIuSiJapiYgpn
RUQqhMIKnUggAguEIj83Mr6yrNJrVd3vfZD8eV3CeVErhaRYZ4e3WMRgZxpTi3yd
IH4NmosPL3bkhYLDTUp57LnrglClbjnHSAemdvWTVEq7CFAtcLgn/EbeIn2/YJLg
vA82BY9Wa69DBaAjdiPt9tcdDAQjUIq1ASD1IwP7dFT4cKGfroedsh75Vah4rpvO
5hyoTansGiNP7UnOS03l9VNWll71sdk18E/b8o2USPGwJ5uOGXgxFgtSbPv2gblv
6faD3n2TAbvdn82aQOp8q+KmHx0zvW96BGa5RTQxJqkoSC4DrJrUK7XrWp53JOyl
iD7NfoihIg+LA+XL93yzcNVsxm9kR9XTze2UW/rxqJuPI1bRe21zkgtX0I+F051R
rwh1lF06Gw7WYMtTMO34DS5uTZD2+jQY8uNoUui/J5m4CrSDoF2JqS/T3By2Vihh
5fVr21zZKaIiI9nXjaytiXxWhTyfLRidtC49uZLq6gAKfZCMmpTx08SAJwp28rJD
wzY9txvZw+qg7nv4858uJnZYxQ7u2q6q0LR47jbmu9qfNjFxZjBJmAB4CxLSNCyz
5IOcPzfFonEJzsKDV1w4y6CJhfyx9pHm/9SapTRe1mpDh3vS8mk3afo5Rqoi3Tmp
KFPStZxdNiJqL7WhNrJaImaSpSwYP2hkAj4hG2++5mEbwF7ubMXARmwVrRVDhgws
STG2NUWZRpIVlg4v1D9TgRB4iJ64j0Uk0Pga7jGYWunfYduFZS9iE1PV8ex6bf7a
dShr4zy59qZeKwRVKEZ95eppAMsv6YNMr+wJBRpeAD4TsqZT55CIiYOr3CbBdyih
OlrZkMxgii0omOpeDudqNLCPeobJJiUT0JWtILTQZUcM2aPPLHBKeT60DvrMf5d1
9z/kiPSPHYQPvMvqZgEX4fv9eno/WCsDw4ABk2phcssKQyXdetHJ1wynbRklIei7
34UNAFZwwIPK6ab9KyOz20rxi1ps6XlDDmbLLfStbaqpsQF6qekZXxe8mHETzJf9
2p3PyIAvLghgAN/ez6tdoj7fKXbTXb2xyb2eht8FeAYN3eb4q1PiAIaacQtPdY31
R6ZqWyVP/fs8rwLXDAV66BTRdnUVsKTvBKUxyTwAf2QrxST/WbLSmqilK2e45Uou
VpBPAfJ5VMyu+HTb/5/UAOtG3vPgDenGXJh53dbsouv7dOOFwJue3zFW8o8ZzUfe
ReqBM/5JFwlmCFfaQ2l7BN/YMN9dS7tgc5Gkux/WvRU8kgCcQFyb1AKkCbfxPwYt
D7YowWK/YmX5JGj1n+aiBQ2/IwmIDk58lmjC0Nmsh7FW6/B8sX3un/2Z6C0HDFuo
cbB0pEAWvcxB0X/jxTQgvbI4wMtgs5siyzFg4G7SQmTB6UpI01Ep6svHB2r/2jsb
+ZiOugk95L//bgSX83+bStqHLu3XXnuJBHqTnhUgeeSxZPcI9ZgGZSkJJA0F88gF
g6RUkVdBhP5OTsuRXY5OpEDTpiv0JobquuWTwz81c0aw79II3axNIf+fzL3smZHN
/Q7ki+LfNlPsq6gbe4s78GU+rDyjgzjJF0ekDW+cjRFhKeAeDr3J/uxK9q8GWYoN
qW5qSpWhwv/CQAQ+KesledEMIMAqmz7BK0EwWLwz1DitwHc7DFNIibNX1YO1zUuv
x86MULkoRcUHyK64o1Jj/YEmRJHyRadU2ojKsdFd5ROBiiBr1Nj91m48l2Qzb+zT
wR710kj/cCoPstRzKHH4mFv0nPtyNB5vCNS0QV9pRjYkT0X5Tma3CZbyPdJp+NKV
gm+8T+sERv2aMRN9syDtPMUbpTRaSPjEnoUSWsAtiosWbW/eoJORebMaqzMY58qY
bUrr/QGjCt8zre2cGDaBaBmL+b+LZtGJZUYSbInXBGtCcrTqXbT2Ar+0d9Y6CtSi
Bb7EVUuHgoFYdVFIbNkMdebNKc3B3VgK3LtOsXXmd2XKvPoZnsZ/CLTB/m87ptNx
A137UhLBf1xt4VBK+89GkHpov8Aj65f26T3ZQKtiFUIhjzUmnRLLViVvONursryI
VRhUgAjcwEtPIrP/dRNlImI3r0fVcY8gRi7FHDwlFAm2LTFEV8IV9hUCZiEXRIxQ
+q6d20GRFnbihByLBf0B5HCz4xn4hSgG62SNR8cm5NLuvy6JJ//G95ZCTG5xo4xZ
5HK3olPRiipeevOkALt61mEk72D0vuTaeHVCn2vYefd5kBP76SGIoS4DTy5gcKPw
Tlp4LJR0rdk8kdC15qz5os2wvQKRYH1M43+nSyv+zCci2sUt6sKwzAJYilIcIZHj
TDCMhpgU48XeT7Bie5XRqpD0MVJ5zwIAjdFzJoQlg3N5SHn9gAL+W/9fHK1Ygjwz
Z5oAHtWMlo0TsxJwOb1ESmW2SV084SGVnBpxLIyZTC4sw111vrBkgcfNDpHS70Fe
E44Slf/RwxSssadUTj5Mmf1twV9OivAoGTqoqInfnXHJNqNRMm98XbnXjwD5X43Y
Yp6dPHnEwJhRF4KVb+39SCMX5zC3ZDWz1aBKbWj9NvjZqCcArkYRn3eB8wSFfjtu
5Y5fzV0pUUODvFU/nve2vj0tQqC2Y+YWFo6pCntVbku6/9jHzeBWoGJmV7kBQ0Is
p1GlPn664E2GD4KzFMS0/ENGTdduhtOpFcp7JX0PFkf5ZKPLCrHzDkUO7ZovQ56P
rtu0aK2Eul7pZUzgF7p0kxK+N6Fg7TWYGYmX+XHOmCWuh8fyQujrFpA5yW2UUA8n
7Q1etN9YI99NgFMQ3zdXp6ROJto1cZ5Hn+OWxSfAGQWcb7VzwOtDBKN4NXqdmzaZ
i4kwcbVGl4Kj2WK4XmaKOUtg5PX8u7XhTQq3DW2hkYwYsj0WccwMu8EjIolerUPG
DxyB40IX/2iUJBLADejYrsjT7/lh73xXaxWppBUSLbRXaBr2xP2OuevxghLpE3KZ
P6WVB1jd89LmR5WfK70UHbQKMrzlNz0NurjJL7zi4WZVohBk9iouiPONiRMaQMRI
rbx9zHBjLTb6XL0zbD96waHLL0cM7wum3MVpTZQL8xB4A61bHcbo4tumda0XLuZN
XyIFHDAuSpTAOV8j6sE56Zad7K5EF7Q/e23QMka+WPS6rR+3TphrJtJ6Pn+lIrX9
j9JODeJ+dh8zlvOj9IuQ1e/zMM4oGYKr/OR1BnkZ6nXmoeVNrqlLHPhTeoL/BZM5
nPWN/MC96DzGP5NXaJt6kq74aD5UvvJL/fxLqAl7jq0d3b0MH5w7/S56DE+ekl7j
buAy46sKY+Avpsw+BG3I7fIX5GjWoot2wCjVVwJkX5wLW49v7QsBtZj8CUMCps2D
v+N99Nj8njfabV3Wx3KP9hlF3sAIg6vCuZ9hQUH/OmQzusgkUjo1l5du+gOHhBCD
+73nldmAU9IU9XKccw0gvlep0cWyEhIqxkbm62DVC/TCc7KAsRQK5RJLXf67zWRl
98KJUVNCHjh3EjKBra5X3lgCtZ0e957mnpWfGrET09IK5JnN6eT+4MBXJ7BAaYdM
zL2RHRzv+fxXjfxnuoQb8HLK5zY8nAbeS5p1xk0P0F+pJGobUp9yAU1tg7gA7y6N
PgaCLi3WaopxgQk+gsElfIdMPLbXhSfLKi5RTrPLqtBErGBGRxcQwMzFA4gzmE5q
rPoyXKZcGjYdpJ6OWKNws3VKtvdcie1L7JYOINpgE2c3X2igB3mN0TZpMb5sfZPn
pxNkFFWDVw0LqomPiT5VHFGw84VjyBLnSu7vyxUOvpqEpy9ljFpuaFlfJTsIBhJP
es8P2cKzupJu8FJG7YzK+rx9lIL2gVk7wpzXHJWscmrZTJljtrTUTjtKmXz+cUvz
ADwljpGIYwzxdl9egKWhDrFLedEzgPj0xSCsD2o8C9NdR8DpYZ5LRf38JgxFHH1W
cgMf5GCosBmvKnNPRcV1POmNpU96nLOgUHIJSgO5jV5KLr3iFOPR5y4MJeutRRAu
vOtg5P1piI9XYYZ4GUrZ5XYwAfUosjKlacuZo30SBCMsojFBab4UZ8CMVkeo1uei
B5qZKHcv8el0P5yn6obw6c9xlpZBfiRSzum02Kc0K1uTOiCBioecVDdb1m538ae/
4CG8DYdNm3TXKbbaTniqkngUXC8yeYviE5eB6XVB7S/zI2PhdCSJJAOU+0quxhVK
t0Uel5kVpb2g5fYWBRFFn/jTafcQ8zuQ4W5i0KbDDc4WbvrokrPubBFBOk23Z71I
fxAw3DLx8eYZ8vM3yyJ873SO9BscAE7A6AIg8ROpJre7S8sy1j12awLw3Xs9v+a4
MJv+MpfyZW3TLaab8thnejeiYPQ+UcHS7cUGzk1Yz7ySgYLeJ4zIDW5CSb2jF3bA
u++kxoWwjI/00KX4bWEupExL21LuAWkVPyuXTYoP9rPZMY0nOhO/gwaC5gHskHvW
ecQEcIBTN/cASrtK0YcU8Xh7hnkynDvTpe6pR3mEVM0OkIY1G3uPRkMQSmvfj2II
VVR5xEGoQjSPv3ih8tc/x6b80T2YPoDrc4XX2ab1DI79PqiaTE+GXv3vkLGEObGK
+StFpnfV6O4G+QBE/Q2WdLrCkxxvbm2epUMwPnt/cvxcaAe6h20EVYH0hI4Hek1o
HskR+B6sAhfFjEqRONIbIbU5Ff1EvyJrmkTBkjHmK8N9elKfd3yYzcBV8V7Gbn+o
JYU9gL86257t2bJtVDfLfunrz+MvfsRFJj72TErPj8R64RrxuhIR3iTAU+HpV7f/
wt9L/s7xfFZr9JLyTjy9f2wAfhZZrWouWq3ZVIWS+ZV5omyJWCA2WdjVc0RMUl3R
QBJKVMKE+SIsghMao+wRn7zfH8vosFm9BFqt4VRUjBf6AUNzm2ibkHHnzn7rrjsZ
s2LNDsoUsqJX6OVmdipiibq+FWQWW0enPVXMK2Tl+V93HKMk2unQOCeQwxk1gn5n
o45TnCe6WnWoeg+nFh/nw9FYnHXIPNNVIZYDsz1TqflSKygsyCtOIc79c8MsFE2a
mQkxLLzQmVX8Z3CXSr+v9W/u3HcVf+gnZ4dQT7qdYQ6Mxzm4Z8v5Sqi1CTd3YAN1
N/8imdxLUOIK1OGw/F6Jg6T97j8NlmpW2eU/iLn/VDaaEvTqcIIrFePPvlE2/hg5
TJkWRa7hyCSbGG0f2KMp/91dwNGFDPHufHfae1ybmQNPE7XrkVRMIdNpPa8lkP0a
yGC58g1FP+szNu0kgR30PnZoysqlFKf9IiXq4T/RMXcUXqFy1YzcDWT2UevI8GQn
IjE4vWhV8BENbK/wfMPjSKn5yEctjkQ6uJgJuCI4evVKgST/iapLxjzQI4/m72GF
cGkHgU8092CYrdWnC3zZEs2VXOnI+Tkd1a7wES5mv55jCK3gHeTa9N1m7i7McAdB
lbDGAfZxG8bCE3dbkBTC9Bf9Gjz7bKqARAp5ZzsFYZTrIwkQgdPY7IPer05Ixlcr
/u42v9LLJkNQlb5q53Z6oBzL4GXpEfG9XZiqKLyzwVMDUpk/nto4tv3seqLEjM3X
yBifnTwk6k3gcAZnDQg1rQcM7G203k0sgPep6jRVf7b6tGzkTC7d15XLbQG0kmlg
vZBroglJb5clb2D5Kn1Jcn/FQYS6sTCZ2H1bRFIQPB5K+eXliNawKCypey9cX0E3
vSCJ421yye+J3xTtPvdLHv12K9AqLnmZH+dnDgfbpDHUEoLWxZyM28wIyKyMNnv+
lYbBStMTZOYpgFfmvFV8UmufVzO089l/0Spc5CDaQEQf8GjZC4oEZpkFzPDpXVmA
qY3POtGO5AxTk+96var/DqVN3wsAbL2HZJuUMKgceMRyTH82BGNREUTHCgZTPtjD
I1IOlU32pVDXMggx4ld3/faX/vDv17UJ6L4sUwESBoAlnrnFwcmx1ZyjouD7lmX2
Gza5BNd5L/q5R5+X/48AYHVUC9rFTSvlAI711kbAzL4bLW3KG6OQkpr37yQjg9hl
/VUKUaTyivDGhn8uN88aUWuGe6luSOG1PiaC/Mi1LtLyJSVYMtirvcxvqN2f5ztE
VtrzcDoOrpNJoo3EbKT8z2dCu6kKXsmedQj3rGt+KlBofHCoi7p1hIrHUmztFfkw
5VYfOd622CyjgmQtA6v7dTwnyscqIZzi8t7ovZtmLJOe3XUHJarGRxPFPdU+OzpG
950sssMv4pyo/Ym/84rrH9iqpyin8xSkA2COhb/HkFpmRYqf2wDbRfhcCu3deDwk
WdYl5kUGr74f5YEYBljA1aQT79acXbWBVRGPlmE96zBE6FAmOPxmGlz6Em2UopY7
jHFPAzPLWe2XdMM9J9JAbJLGghn3yx1gT+2qw/W4aCwh8JknEzjQdEyWmDmrZ9Kx
bZ9GRi5I0Wmq3L2WxFIP6nYt4/imE1zQwIzeRRyqYMclsYJdlpbmuVNMPdMhYY25
7bpT8FlXg/vibt0zSuKsiRmKISOKmYie4z4armW8KeKLiiFTGf3UOMapccDC/FwQ
sj14xet2LrrMLzoIsoRhLXcBJWVg5p628K7X/ujNcLpXlre5eDjxopIF/DFm1gNv
6nHXKwLaeRQb5quEIBWheow2Ks03E6S1R3zs9CnYBZKVerSLwU0Daw7fOKDcQtTm
rAhmbMlPjlZby5Q493tQuggB8hGVA++n8MqUvk66cb5LVQtg2khGOkwySxoVxdOD
9CYMnEyVNayWGyfmkUrt9fieXAgIurLm+zv0Y8qbmYLQeoVRCNLxNNRmqXkJ5ruz
GN95Phho0HgVnczugRleX+hRNnjK5G4+Qm/a3N8X1rLLL1KjACdRcZBI9+XqMiK9
PDjy5gfgzYcjEPJ9uY4V8NwomZ+7xEvoABHeEVm/uBJ3JFQCpEtwC5kWkvaN9A80
4OrEUhX9MJyDbcGPNoyG/VUyfl1MxNzUXhU7yQE77/74YcWHCeQYLe8il/fbI735
9oZ5vVCEUAUHKQzKZ8w3NBya/9PyhSB3rDUpb1y/8E0EsOgGLSi5DRAmRKp4t48A
QshxtnvYI4iorLa3szjZCGMsNZTK6LcLHePxU3kAlE1Lm0weIdy4AjR1KI56RLUt
ChAShMvfaniq8601S8CmCBC5cSoNDLngyFI089eaxg31v0Q8lRKIXc6feOTcx10E
tTKZgh35qad1/q+AGGrkfJDIW4ng3baKTHfDpTRAnWy5VIZjpTK0BYpZBZNyLpCb
SIzfTG0POkzFsM8UppViQ8wWKYxF+4uausnK1Mt7ugonODJ28GPZs77pgKNHtbIL
pkBcHJo2hlD5R5G8Ikyo2wDBWghrYLWBU78sXXwUxKVlU83r0UtESbGyvlxZzD9y
AlY3pZz0c2THKMAfgUiPPl1GFuh91c4OlxZfaba/cT7bHSW/ZFQyGaiawyO/TvQH
jQf+GTl+Nom5YeTx9x8r5UnNEBhbosUNQUuEBDZvgB91VVaZVpxlCzVHc5E/foRh
FSTNSyuRt/wG90foGpHMIPAGCC/5NriH0K4ICzlcf9Jn+RIhpua7cyzH98P/YuX6
CzHJH62XpFPDadxjoFRc5TRB5SwaEFQ28mounQGLSHHSKaUoSp2DfB9rqA1+d+dm
lKGJ+1N90czl0+0WnYf3FjePQQWkz1ilJcDDHB+YhQdssWJc68Y3pkOEKz6OK3c1
ZQtDDPPe8HaVEFlaRAeZAdWIoH7SDUUCTriOOfWnCsvpFj/kfO4GW6RK50eYKVF+
RQcN9UvJDz7QYnAhalk+M3c1qmZh1aiJy1baAETXsmP6mCLONl+PW4+PETVkSmgu
CtwRyU5Ls5amBM3rHbOk9emQaf6YiACdxlLTvCuCowLPFHzr/KSwrfQspzmLbiLM
dbf5pYFg3cjgfIjDgvF1lGA3v3X2cFryJRV2PzcguKC08eQ9J+rpuxZ65Rc/Y+wT
A8bgMm2UG4saLywp23KhyC5XwgP1aenZPCtdIjdqy8JxJ+qtFPf5TYKzgguayWKt
ZaIFMU7OQwbmOznBUGvWr9VcTcFcSEOkUm5bVknisf4DXxbpX6nS/5OOUCUs9zng
YoayR/34pGGf5yFGiCSIljxCjbU3pd81xoV3ME3zKM7uNbBwZWjPMr51w7vLFZgS
sUMU184+COrT02FFVO9SfCY5t7jFZqvmHB1P6F1GszxY/Zx6jtYsPICg/9ZhhEq7
aoOFKEy6H86Y3Kpaq3ZpnZWNZzQ5u70lV9FwOOfUkNzAC1X80MHJJxloCsX0r1n0
VcSt+TLM9IHspvBwBA19oFjIou/FwRc6UydZQ3UPPrAePY9oTm04oTLr4jcr1CcN
/r6OScwRVuojPg9bnWtqEpfR4why/GAAFI3R9bgvz93hfahHrXfPEuwt6KIVP9vz
x34aBjTfIpaGftf4JRODZtzwkNxeKBDfFwjLWvjvJahtMfV+ICMdY0VR+/J6ekta
QAnYw3dOuxqe8E3MB/KnMyuA5cJN6CG/KvY2+ksZoHtzyPwrCzzvfhRiPcClsUw9
MfFVRY9IYcbsbVnQj6FCw9rcI+DqnQvq5hSlSLN8/Z6H5JXzdyL2WUBiQ2uTlczY
r+pO07Lu/ewu9YS52xJbaFtGyizWXGClkcmQOmVvnbyN2sFG6In75mpuAq+qqvqe
qISOPWAg4KIFSr4i7X8yDgZG/masPdM5JpzrjT2vkZXugW9zGjFHaxRs0CCX410y
spJh7Mdjf0vGHF21pQy5oTkIxuk6q+CIlB0udejA0RhM4TGOq7Fm8D+ynkVdTefp
Hx6kbEocs0r4nLKLWWT67J0lj2kcTPpod7NovjatKaZFMLNfatxdQWtcxKNJcnbF
s+sWddnjcd9ZSfqqlBL+b/oftWCIO/Tsana96YO7trJIYk3Kv/77NKlsng7oYoG0
OGw+DL0+Q3t9OEYpSAGxN8xHRkL10wkWIf1lHNrKsIwbu257o6ooWx8K1TekkadH
DbkCmZMQeQtN+FWNBo4pRpNLS/n0bzlyf6TpaJ5ymgn0jV8bsbsekHMdY/PKx34l
3+cXzKRzYhb5GpJAF2Zp+7RxIW+eRcBCytJmtzDqWW7647pyDi5JYtE4DYroENX3
FBAFBHgEiLuzF2VLZ6zNcxQABzEjGVSa7nbQ6IrLHx+WkWuqutfLRSUD04BK6FMq
AZOciWiwbqbdY0V3XqK9pzPfBLbIOooiCtPEGPzqUNWSqr+KpY6qN3QhkuFTJMkJ
Szg8+DJCIR20dE+QnqXhi2gLhUFVIGwQy//UeD6EurPnYSDlhnNCIMX0/b4p3Lpd
AKO5baznXpAJdprflUl31/CiZUjxkG5PJq7BBd9gv0VZlhUd6bUf4Moi3pe/kN7O
bklYe2zcpswGGokJUFisaZDrQxGvMTY5dVBOFJSKT66YaXWNk3Yz177SzhkTrqBC
7JULiPoRcG8dos86Np1NQOhYYH4wnODexPDaR0XRwe1yNCjQxXXlQJOyIC0UxoEg
jWk/3RpXemanas2DtnNxL7VsgbnHCqEyAcQhvDPwUDN9jnSD/Q9HIJY+F3E3QnDe
lOfGcVd2lA0lnPOji1a2H2/lN4OJzBDGBSBPFXULAdjUOuXhLlmYr2+hD/qsyWWU
56kLxMw4Fx+mS0lpCMPCLYIyFIsnX9iOTDW6aSQBo1bfCKXHDkMZpinKD8oVP7Ix
fAsf9dOxNAao/Us3wd19rWCJNN2uBn0m7K6TJKmrItpESGfJ3YWu/mFk7rZCMGJW
JdQvl89bCRc3gygZRsY9Rrt+tdyWCP09lQ85kyUmytGSF9LIfAynDXWSrOiNRYdw
juYDqFwqYV4IyvMSKvyOqV5aSA0gDj8X8GKtz5tdBVnteiUGFeRm5rwSTXkeoZV/
a6Hj1MDpWvG+5tOjmXeHz8Jy7pEqH5jicBGnxmnPuRpI8tunQvmsZw5etaCNaZhb
/Nqj5PNTLcCFgpItHTrbFYwODTpNKxd31KDRMsPlTVnX6F99lvVM0A7EXcgT6752
XIjY71/OZV5a178ie1921HGft6CB63xcUfipKJb0dluZVnhY3lmJDhB9qoLJZr0Z
UiSyHPeIe04SwCr/seSoWb8EODZXAenm2wWEHnOqiWmlOBrQdt3efXOz9Zh0OGmz
LzFNVMUJEozt2wNyIwJvwsf2xWSMuRab4vrrMZUkQMCcJI/gFcnxfdmmf8alZpcO
GM10ksm6/k+Ic9c5wTVK8qd0TWhjR0vA2W9UtMngKSwnC66CQy7XMYfyLb6d7EA6
V7UxBiDaYETVnizyQElYuZXfqLA/Zu8pGtjsJIccWVxXWq4B7hE3er64lhCSS9sh
636zwSzygm/dCH2DQ19qTj7q7fmj5q4dneA6ArKZ9J2FfjS7gxEogl5+S6Jg0CsF
7I/YKVUieBHo4qWpz5Hzsc1Fbv/IJ4RzjkeHwhNgnsyk12wTX7fi+w8D4lWZ1a+V
UkHe6qqjlg2CgnmTAVfII5vblMoFfGT2LczBL0uEvX6vwNRsaxOsW8VXosyqVM3X
qiGiHBN8K+ev/yqZZy/YoYtPy7Yz++GI4q+oopXuH7aF0AhkrIbxKXtPfrlwaLIJ
sGDS5hXMoIH6fEMGy0Wg57fWYNVRciXasHeOUlrhFeUVh751xy0vZFJpvIFG0HMF
JaQEkzRDeKEPwWDL1EiX2G8EiO5wVi7CPOlTEB5Qk8rot0IzMKNgy/2zdGV0P7j7
pfmjlUo1E9YUl/kJzB88dOgzILk9slhUo7vgrFCgJsyUpp9vSwwl/sqiqt4L7jb2
fFthDsdpegbxciFYPe/3ZDxifNt8588D8C16PEFPRGFlSea89q+9YrYr/a4SU/kD
sEGX6iIFsVQKpsxjJui5NGV3j/sJyq4S1T6w/N0gDbc42NrMrKdEc3tPGZU+cgNG
jNUiEfn6AbvaBXC8hmgX7BR35uvgn6rkVbIdZDXPTuXrLqAGb8pdTgoGDS2nbwgV
8c7RSQnZ+i8H6euPC++KZK4Aant0bxHEiC2F5/eJo05pPmde1usUZ6KeqNNMqN/e
FfPcrKXez2pyw+jcSPf4gmbdF0ybuP/s73ATEB77ra3JCqxIZl0wvbwtn5yS3UYd
GRf8OCcNY60mX88prYwqVrYpYVg4eshJDEDMjAeGJVCGqfOE5VMzhwLXLdoxrCmX
u07EdG1OxQZgcZ/M3Q8bSN4LMvOsxK5rtR0tBh32QrHHsh4VmNfac4p9UfNXh4wd
axJEfVswZ/+0ZLY5GF2OGIZxP6i6ZyTAj/GQUWUqQfGqB7AJY1nZHa5iGBUHOPV5
hAZMZo3FYjEnp96XF3yMzFJp4EncTpTv2wF09bBA7bUbfQ4Ikq7kQmJdLrxfmwKQ
PTmrY15FhSW+8DHOlWxDFgyh+avXa9rNdU11IUpVAmXmExVqA8tEKcd45fWRbJ5P
26emHJ7ouEHTwOuNXZjxR1fecv1w53KMATBsZmIUxcir8nZu40wWiT7/X1lgCHuR
A1awXTwDbYw2ZbC9rfmEL5HND0RZ4RVSzQeEEx8TR5IMs8MqnMGEYsEE3vAmrukt
7UCVAImmkIPyKPwhhzi6BhUCFjf6UFBEltYr/IzsFtKL55jCnkZz/4QfMDFwlCAF
gONXtglZiXwB2UyVYppkZo0O1yCbQ3fa7nYDf212TAZB3GEPpbtFOAVga0OGJUGV
IixWQts8U6BfBQmlA5HZZVChStq86kWrK1vtL6N6QhaPDTRjpyVDKAhBDoLspNfq
pL173GqQFmd+NVyEV3GTPSD5hCIm8agofe+fKHpZxkUPNoUa4g7jlIGbIMg/lfmy
uITD6eWMiBvx+bmd6AtJe/Av6T2nnzYvU34yTYuUesGMXu9FFNbPYnNm72qF9EqS
4zpfIXqHzZu0ud1pfXit0SjuvIgLlyON+M8L1hwwmbeNNsbbN65pllCCnAaT0mK2
epEq6c11Zi9Pip5XQe1iLy3qh2YEkkdJaCz2um7KndPf4PabviWHcBXPMbCGRfFo
rtxA+yOyPlx4Mqt1orQcseL5CuX7Ay3VNAPNIjHcykcghWuPAm1nv0rMXxA7QQLi
CnijpEbUZdDJ/wpUUYNFhb9iLaQAozdyiruC4En5ay8VxS7gYD4FA3N/CkgaOhoD
1Zuyykw0dO188XPO6MS2ICX8Fz/HLv8O7r8fldw4apHcSNnBHChy0wmp4ZMMft8f
78iVC51/odezyrTjqT/MVeSXO7Fjzl8cxGKYKprRGZOjwnD8jGMa5/kXo4jL1Kxp
GOA5oSf0mib2B+1LfIDBRLXZbnjVqNVJEWxjkjT/KKTV6t3kbH2EjRins7hKF6KT
lD+sXElTlkxugv8OMLryot9iPJ805cjljd9KBwsjfgesfr2pV6MbdvzjUHgm15Io
/uqSYEhQGcG1CojJa0v3feKo0Nhkj5PnbWJCTNBp7x4uxq0Qkmj0H1PWcMdzQ6Dw
ivxF86GcQZXUi+LnG1hG5diny24nHjr0FrNvohDxmFABh+NMuFiGjretmKLlmzLI
BYGgmyRz0/YbRA1dAo5YQcEUQ7z2lDyQ3bSiT7tf/C1WCDClhbpySrb5t9F/3l/F
S0VyaWN1Ymi66uK7QcnGCiBXc/xLnEyAkYjRIHPY6yY6Y3ovVHVU1k4Z/fenUel0
lpQLeGrPkfHiOYC7mFW91DgFg+rl6OoTZkcj8Dx78Jks64YQN1ZDwxoqmAO2+xjb
/Eq4yrKmCXZ2LSoyINV2hMSNn5KSQ4Yb54j6rG1bUCqLECu4XTzlMrgbMT4nvBZc
SqA4ld37WvoGdTxYyMgbZCnFheDqbj4EwUKHQvJGl2YQRQRRsGh1jpgCAEwbhxbw
JEritfOna+fZ2Y1XzAYg6o6hYUu0n1iKZ6MAovLf1kqSMJ+J/zPT8ze00vE/E+LF
mNHhPQGJiw04rbkh1md1c1c9bKmN06yIpJBxVaL3kRwOC6UZYglQVPNh9MSl66sJ
m9wbZdRmei4tRmRvafPwwwuBZxiBbtAsZaLr+5qR+7v8ygC9soF1VJgxjI8Y3xXf
Zo8FbvJMyB/wyMYjGPnuXN80m0KVpmXLp+diWxmi8MkiUVqp+TwtzEs7y3gfl3kn
x6NbDKsaOZwZ/QznrnLNYDueOil5v8Ch5xf5ObHC9m+YJSIJwdaOfV3MK67fJ6VI
T3IrNcG7eAPeYaT5wPfb1SEdHOWndBnC/ZgwRaLu7CN2EARkqPH5IIrCq0Dnu4Af
73JuE3zNB2Pp+ZGCLtF53AWnq9LebWzD0ydU1SrxzTJshACPhR/cgMOF9qGqDnR/
lYSTQIQu/3FbGxTrrtiGhl0xc7gRF65oU7N+wjaSf0A/jqlef09QjJ+m9yOZn9Mz
z6gmIzvMFCod2IWbxSLN01cTqT8Fp5RXsYIo14QtL1ZPvTGY0U3L/Ulx3ic/0iFv
AroPD0mM0nePG6BiHESVBkue9XRTowOCAlx3n1Tr3V9z0Jk++ViglvOnKR12Ujjm
WHJWZelyuAE389IVUtnajDmpvBT92uYO2OawQ+92/e35OKVuGKGiAgHbvlXRte58
5VXnA6vAYRFYBQHgxqfJXAX+6JKyWQiqifod0LFv7L+jV1kM3XgsxZTzNbtGkvI1
/W0Z0UelBkt+tNfL///3Z06sH5Yv+XAHxbVLg5MCn6mQ1sLk5VJEuHMn/TNVadMm
ogUfitGc4ZrvuteKby+oUeV3dPevN1+9BlRUZYFfA3DRsiJa+CgJ5WPNJIZJye2a
nXJ9xpcCdkQVsE7JLLZAa0Ysd+9wX0ElJ8g7Q5WDh4y+azfiNo03aiWpqOvv36DR
QRHC1uju/5tmWS1EwIN7AA0X51yf24bowOnO56+bY5ZJixmCF8wu5iHpThiHyp76
MNCO4EzUj1CJGbzTLpEpxoy6NCNINuzIB4xX02Rc4goc62C81oShf/l/N0yvnzlq
uZfL0XF8OJCKIdBz4kaQqmTXwSwKbAvb/qRukTvtt1hc15T/0x/Wh3RTkl0xRvc8
XF7B52WJeTTgZajQ7YqM+kMg66kArhPQA+JY8iVLIOjyJiAmpR1aoInu4uNL/egJ
TJHWWOONGykFcyDJ/5OFOtPu2KSM9quwYFstcQfKxYa5gGzjcP8/S61XJ/mvDkwu
ALz8AhfylOnF3/WFhOtMeZytSB6eBU9egVodyMFQQWLJxSMJIgSApWkUKN2CyThI
vud7EqjvsYFexBwztj9VLpeefQLdF7V4IBw9ceSXvUym4DXGjJ/HIUZwU5evBMNw
CFDylFq/dMYSmzRZKvNLy0ksGi0+IokxvlkZ/Ir+J0kYltPmqk8nYr+aW6P60tIe
I9KAPHWeex1m3+je8gSxW8Lf3mLNW6qL6IhOeIpMmw7+riXf2NMiq9NjhfLFJS+2
Ef48GIk2Mkj2crfh8C7Rx5b1Bewq5ut3sdIFYok92KcZg2BOIxeNr3wPtpIJIgQ2
q5VT+p5hUoIiLhPQc4d9BSgIcYuBDp9Xl8Ub/1Jc+jUDibxYlcuxG4hp+xKNeb59
GOGz1P2BdP+SzJfcmEFKOgPaUzcS6WMaBQopMjNWh5zTsNAz1OntxhQoBDqWzwjG
b+tAeJUw3w+oymqi2/frbyfLgZZcrjN1P07FARVYRZPIEaAzRI5uD+tn25hxEYqC
/koATGJL77/xcxo+XDchQe2wsJ2legCrynDt21GqpmKDjcv/i+k2ClS0dp9i95Dt
ZL3VsgJ9K/qVJAujLcRR4BhDzebyOc87tA8BmYF64KTdmFocmsiWpK0hLPT4AuoI
4VwTjOIsiy1cHx56F7hXs4MJfC/49egSnv/k6QaM6no5XWB19dZjVjcPn3fh+eoc
Ss5HdRnadkH1R2g6Dc2FA90j8BtInpDwSclN2drd8DCVSWRcE9L1tMtf+uliRjPy
rUotFmPuApNTkclX0K2uJ+QEav4HGmh1RaNiE/zkkPvmceh/8L1OOvPwJW2BNvsW
B4Tc0LS2WNoR4TcRoaYHcbvNnci8kqIhlCM2BNiGV5NeLgHKQEZqwZkSif3AiwR2
Xg8IIJ1KqUw8MJ3l0LGwpw+LtWP36R/QtfQWyXaYcGK6pUd6bModmHQBsiuYFqi6
bPDVyMPkwH7P2T9ofJbQKeSjo1a4oMbfS8nQGj94Zx/WaQOGhH/1FWLGyDUZzBMn
5npPK1e5drOJK2Yk9c8aCi2POxsoIrT/fPzbP+uiGGcjiOzMriuyKbiqjJQr3EmX
pB97tQ07+RYl6VTS1Cgz/b/a/+f1Ss3/sDD2j+4wMADynCs3JwFZpdL43yCmzvRc
lfhHD2NrLoVdRWKcwP4vtZgyc654WgsbJ9QPfNE3OG57/InsTM0sYQq/+Zwy5IUS
FyV8FFh0TVosjQDQr5plLBZwUt+3KR7vLmc/1C2EUZSRBhLFoshJhKrpSlXXwUrg
eld+SO0aB8ErC0KJHFbfi2Agym02dZh1P0TOMR8+5QJSvq3j3atTgbz9gvI8R4GN
x0XHpHMQhLwpCFMrqU0dtG6WnNlYdCXhUsnZn4CEZg6KUvKy9/ChM5JWh+W6Vkzy
vUyCMMrsfKpRiz5bV6wQq7s9yHI3+nYwwsCHPaVc+PFCOOMV6ej2REpwalhXcvqE
xKT2L0HodW0y5tpFOOLB1ww6D5ezB9D7nJDt0fBDf2cAYz+vXkWHW73QZvhVXE1q
J6UEnk63YimiE+ip9MBs8WJ1ZBTvvoeTqEhRaeGkoxWj2hbF8xJiCY+ymPyWfWPA
RWzD1iO3WtV4475uRkEGK4hLAX0HN3N2UUiQZ8+C3fjFMfCvFpjadksBaeoXKqhi
8PN+PA+swZyMN6d+i9cfACmNz3iWzk8CKeTGtEyNNjkV2hZFwW9hFGhSmVoXMPi9
121mUXqdayHS+8DkSBbmafOo2OPJEF5OvM6tWU1EOEKAqbRV7NgoKseYrgQb6/Lg
vfP+MdTpQV79xwpKUioZAsioM/k4Irh4Kbw/hjUVqavG9szRrFRIXuBunG8uI5tT
mHt7oUfJubudmntMDaWy/KWqXgar186nb8+YS2xmyx9JOQr0M21+Cs9nkAdFof5m
hGjIWMLdlB799PftqR6cuETrCxGG/vm0wgXxJTJA7XjThkdRSYFVzy/974vPl79z
suyolZvedFAuR47M7mynPPKNSFDEkpE7UO02zg1YFfUe4wmK3z97Ep5REyS5DKLQ
W9QVzRZwIi8jzasin1JJ9FSfJLtwQsbqX9hDr5OUaG5OEEu7JkGdafLw9nHqfmPB
r+jPO1PkEO5tqcVWrXblAlSDe9miEN0PbbiysJYedqIx8u1xVe9SGmmNEt8cAT/B
3mQ+0Onq/ChkfW0/TGjaSQDeghTe4TYIo/+HlltjNoHDR/uVPWKBFNPenGsAIpyA
Ab38zCN84czFaArWjnmcnUqwfhoI7Cvkvi8fZtiIuFi215okPfKq49Dd+ZcjK7sL
RW9w1Q+p6stEzseJz7C9MP4B6Le0ezLezs+GUOpg1h39y6m+1wQ7F/GkqFlY2g2h
aoEkxHQFCbUPQ3VT7AU+/WPvmKXWrrc48GY3dtluLYK9fHPOZZ22hM4p4wLkJ3T0
B5/ol6m0KH+V1XMiGgJDYn82HQzeKkDRZw/E4/IqS9SBlptkW1VQrCuN4vP585OW
GpnBLoJjI2uhohXQMzIJGJsOUyOZHSyv++a67EKhxHBxcw4dc/RIT1lCXXikrekZ
LYFmWBt7DWqEInGVFs2afu2STBTWK9O273caEyIyASxSe9uJNSfy3iGTjD+FLF7w
xch+ccNgcqVCEpiKmMczv+fd1Ejv5tCGz2ibCziJtrx99rISXHXqx7A90+YtLwgG
u73kvRSMOBvrwMJ0Ubp9q4e6xTwLUyeRItU7aCLWiR78NuOnxo7R0o25bl8Haq88
Q+664RJVoQVfFqMzROggTM+DKT8vYxGo6lVvrOZG3bPjnVDFMET0SX8U31+CnY90
bONHtTu9OgUiWrd7195td3hQ2nV1zrbz4DZsy/SOHMahjfegW1DSG6pzP8rmWxZN
8BruMb0uaaaGKQFJz5xyr8v0HRNjrIMARDCILJ4Bgy9z2u+A5koB6n7haHV2Ikbt
KC9+6cqpByiEsvbUWTwyxgq6EdXRkH6H0ykAeKLK9fFdD/lu2gN+SKfFfyeFKHCa
ZyTZK6ry+My+XYNUYklwAtqu4kdtzxNufg4IDwY41kz/4KX23K4lQfqG8PSmwPgV
98M7S9/yLAnkQRfqTgncpYAWC8VcEKUFHgToa8cNR66H2BCkjGZi+/2CfxE8Mj5S
sWQaNCzAg3XhAx8rwYC5S0opY2cNO1o3U6cTtOKEaDkK9T/Qq8qUbNkXdcG5NWJJ
84kt06yrG76cs34LvJmY3yeyrXzp33+lDZ7rh08kY/gy3kKRPuuie0h18m//6e7b
suAgSYPQJVtDECI+5+V8Uy8nyrLEE0tCH3xbJ61JEerHL7aS38u3xSF1z11pJEr/
3fQeTnVKyDdqrTFFyhpTfBOyVJIoPDOPJtSm2xVatZpj7brB/2vSjac98X0s/uAF
UswHADe+Zt2/R0ojq9QrCyip2nqoINsXupXd5jM3lribspUtsNCu6zabUjZSIpgL
WxITNu4e3YDaPbyTriBluWZCn3JmGE1wYeb4Aq+c3DziwqtI9TipFj82KyeCFwqT
nVYcDeyHbrVHVFtK8kE4pntTBrFteCVEokQO7Ji6yNUIV+i7rz87PFnacW58HP/l
HTxH3mWZ3kNW7nt60XUq2XP1ejwevKbTNpeVv97L7JbnVYWEtj6BtQC6v+Xlwlhi
GBhh6iwls5cqTGuhok6CuUgPWP+N1QWhOKuJGxlNGWf1bs0e9tEOoAjerRp2+sPD
PqLl19yPfckY1r30iLwBBWNwvHYsWO3FY1ZNchgtJt4TV4kNi+B8Q1ol1L+zwXZG
C/4MFXoIA+eb/W1xYUURE+NF78DZ/A/VGjRXpmcZI+IH5LzmyiUiKtcHB95fepNm
HPcfayyuTpf861oXVHp2NpiQuSizOQFEsRSksU+EAIzB+rtJRdASHOyJb6lO7oKF
HT7TF9fvEOwftP9YkdJ4Z01d0lRXon5L/6iSUexM2JX1yFKEPe6w2EnOGHtjcLs0
HUAcMUc4ppSqZR6dNvp/BtKpmFwoRpxsJAJVynQSOQdr2kOKN5Znw4QBtVyKXHxr
7zNlfQCHo1b6MRChJ/6dtLcwFzC0Bxlm3drpdETrTVaMUHltEHF/Y0ynxiZmSOIe
A+7wwg8pJtoPCSRGAx55rs6s42hUrEJKLzGqr1hsqfjnZ9SUCGXspWlbLVgm+Qn7
hUWydVlElnsY3bXtg8Us6eultvfju/bAV8JkMp+RKrPyW1OYo4hy+d/qgOq+uh77
uNMSg2Z/MUKfZJXxm55cfHjKUTwe0SsNRf6y20oEgJO5NW7gQ+JZYJoWY7vJGzF4
ZSAoCkBkPWyHJPvxDbmvF2Ke+8Bs3UpvEjrcU0TJmhL+qV2SPTXisWRewG/QXLqR
A2QD+f01SlhdhEa/W0ZA2V0Q48LzoqdjkYGiJv/MrNI4vRNiATe/vAPTX5pv3uED
eFEgJ0YGCBgr6vDvkyXoZVlItlX3w0BUiVBIYWc7aqSCXB54Cqj8CAfZR64GXdNy
WlAcouwaLswEYGVBT0P+69mOUwwDglD3TekbgWqYlewEFbBGJxyKK0GgGJAEevXI
dFAJcE7XFlM+Ncve6spoz60Jka9eml5Hx2Ey6gFlLD2GsZZQM9+cf4f+uNuVzuDK
PQOBhSQoCqePH5fFtHCWvBS9ajkSayTYHKboa6HCmTnGZL/h+BLNMzoiRXPIoCQS
+bbkiNqlzadsRFpgYx5EB1xV8WS+9LxLAVz72P8ZPC16KywLfhgnohLaVXT5XWjP
xwJxor6gRhpn0s1AuhXD3nichf0vd4iDotpKe64azlFwVgCPCl8GTjj8mu3fWVsa
58/vrIuhiwD7C8Z8gdk7VzklGcU7Regmrt96qklaoucLuBd/BEHgVTY9DGefsLJg
bpmCXxL3m60uaoIXM18f+rxXxp8nFF4sCJmGBmjDb7kz/UMg/qbFT1UGm9w5BE8x
0ah3vwAIIr7PvQT4sjM1WalkICQARiRaloPSCudQ0NBJRndWIeyEzIRdATx8T2/q
8BV/+ih4dIIQymnzb0MNRyLjeU9hvR+JZFTEDpETMYgQGtSdTATNfNUsEMcigaWb
8TcvAb4aH2EAzo3rldHL1zk0r8cJnG+uOuQoZzfFBI+nJ4gAwBxj2P1T+cnDzZK4
cw+kyxhJvMsfkTy1A+u2hAvWRa0qXxtxHca/4SD5rrbWSfiKRWLkJEZyihV4E3eN
r/ej4rV+RAvRQzmJav8IrPfS6ZhQ5nNnTyQQ7gSUX5ezqquqyzYkuDX8BAY3qIK5
EsSeNVg0Fokq6b8rbLCh49YwCEOCpil5RnAct8IpNUlfb2Fxnc8LOY6dEvbLnAw6
Bh4GLu/ur6rISEsMhqeRZF2WBAQ9YsWyv5qDjrBNAV1lYUdLo76YoKxS3GmyxGnc
ozXKSQuP2rWgE7Qe5SDebLvJIUe3o9jXks8S1v9T8zmXsx8QpqII5RTew4lGz1hA
sElRTAkF1XK7g+RpO6fC/A9a5kboY2diRh7bdv5yWegUomP4dZX5Pq1cMMZNmVeE
n8ZGX4Hh8u60DOp8s/AwmWhYrzl8Xnjz5muWKRodXqFSwycZ0LUO0QWjqZ3qR5RP
gdrlAtJpCHk1o0qHMPlkfg5hez1fiM1raLsRxyBgQ7rWJxgHC74w0AB2NvX1nym3
sZAnwtTHo6kkzxTHA7ypFu24SDw/DnK+Fh7xVSPApSiunHQMwDGqG3UgrmIdQZkP
9QvhkSpiE6UcM19KWEBWiIqYyR14M1/SkPKLIC2jeQ1cAGXz3calcAlQmzGJ4b6O
amG/Jvu/Omgbr4L/Ochfad9Sr5ySMemf3w/AhcFHia5REj95kevno3QR9F8/5Ukt
yN+EQphTHLZ/vdVASqcfu2D7TjyKV+RRnaWIa2/dwZsHyFPuFJM1FcED4einsmJh
yLJPUsy0yElzb9Ynh4lxC5ppE9M/eFMW9tbi2B8SrEnDddSCQZ26oGUAa0NotCqx
In7Q+wiePiBra/jIjbjUmwwVZW78U4HsSFKAG16DjVtct80sGj7uXOYdla/259hS
F/tmXFQK3iHtph4u2Cx2yJiC4cjH20xU+D88S3DJ7N3/RUglkMxH3B5vTMWSdI9Z
zTc+aYtU9h/U7oyt4RE54qgIAuvHctH/leau9kB8YytatNfSXYiLr6Gc9sjgz/Yj
uhirET9Q2BasU9zrBcv03p/ucgBenlpYz8l3llDX2zhfjnI5gFSnegu6ZZD+5UE7
ULoqSiu8rhk7FwwNcYBdYZ3nMPP6ZEv50xnfjpcryT4CHADPfnV5PNVekRWD9Epw
9PQN6o08/GopsWA0M8Xp+fQfy4ysfWLYlUHhynam940vnVv+PqMY5fOJ2A2aYQUk
8BZLEcgX2KRlFtG4eUYxw4kVq0IUYo22WEA4tfVcin5pVm1Td5g+LqgMqJVJgrHT
bH7gfxtmAdY4THPyYFAskrrlIF4rUJ36ls78ssYLebx2LZyqJPSzUSwcSJyNR/b+
ixjI38U5WvK0APcW9ZuqvAjqjgZHWr3LcgGp4OsqAZKkqDMTmGuAN18Ca2OZ2lVO
/b5yc4EdDggVop1iAscooxDFeDofvXxK5CWPEy4YMxOX5FbIGmydjqrcv9YdAovM
heHGMLA3kdqLuX8JF+Voy1ITL47T2rhroKYFy07GA63NxwZqPaTDevahSGx5+nDd
+yjPNTz94FmleWbIdcFbqQzxg7tInp8SlLOJVmoRFczxeC/Ox35DwmleFQ1vKh8+
hqhBQR81Or7X9bgp3UhzSZJnI0KfIUm8X5PgknByG7ZSpJWFHxcaE7e7cUIh4x4Z
ksBKo02x3SomLhNA04hCvCh9cKnbZZrmqF/Tj5CwHeHSvLXWg37d+jIrALV80lFW
KTtqPX3+yn7XJ82m2LbqHzR7YyyeB+nYToTTFKFjPg7nrG2wqPyDeJRMf7rUkTJ6
Z4kIfKKb/+bRExGs08J6zV8gJX3+oSsChcXiROKPn4Z6UbQ93ywK183fFAFOdIa0
b4LbNpid3eta5BSou9Jc3fWyZVNTCdNzmYFuTDXWlxLe5ahU4xEKCHFL40fBTZ7y
lmfYyCyS2e0KxoUwKpSectu3xJggOQJFUjVmUiokt9827dbU/mX7A+K6parWHQvX
0SgLj9NlcJRFaijIFytFeiGfz8hhKkEzyfkebztmzZBRv8MXhyNwKdmPHnYR9Tao
zbQZ7DXZlhI4snwCul03wrv4f7RAEPlKaBklHjWpg1n3b0O/pi2h2VNsv5NJS6Ku
iCUedY1ojUmxjqccMqoLePVsUUg2mSaIc2dyPHknvdunwcnPaySnHNc+6PxOleym
rYWJutYaG+AvDcRaUKMPiD05aq4mYpkqczHkJX6h49ST8NYyAVOdXq+ZJwIX5Ldz
Jwv0L3Y3RTT5/sNBl+2sFDHmbCexSgW4JdLr6V2JYXNBsbo6gaULNXgd1Xd5qM5H
IocVBDm5enoNL4k5wju6hpBk/gHAyu4xYwNhifpWfGpKW4e1mxqr5mcxrFk0xzYL
3E+QDhiBqjyMAzWrFQpf9D2q4hii+q+aKUEXGdXd7Zrt1ivkhMEN2JTTvOfC65/N
2+QTJie4+kcUyrQGDV4xnQU4SDK0NDxrFIF2rZgLtO0SQE1z28eIz3gSor7PcfKc
f2wd8ClL9UusBULfXH8TsGYlzMZiVZMIwY5naUg3jQ1TbxI8HXc5yGlnf2HZ1LD2
MHfTtz8SRxrdJEU33vEDE7KTcUrSA0tfUz/xiR8As62/dYMYIHnC2BCzPs0qmuVR
OMIxQ9Kz9yIUXzfdhhSn2Grq7rcWGovbKMQwKXUW/H6NE/CuxS97SlSp+wL4lI8N
fYoANdv7hqak5WbA7MJUjQQTJ4QkgEYJSr4a5CBNtBZ5O5P5ba0kJFD5LnyrjbUa
gXX2b0/hXQ88z/+wOxSOruxIVrwAx4j3rXHxx0OLgFeizsrbOjT113tyKbuQQj2k
yw96M7q+Y758qjU2CGvUrOu/fIPzXnUxUQrApSYOXDGY42VTJ+JHVI4p2lIVWE9f
RWaglEdyb2hNHoNsnK2WbO7XFOHE+vyjGDGA7hLtsEiRUgDbXmphsZuKV3eJYGPB
y2HLDVOkn9x/M76CUFzgQRGfhhbmJglGvNWykEaqtC/dzrnXsRnHzsw0fzwzAkxD
PKNUZAbakLjoheZNYf4hYqiKyIaTLvbv4Jrsm03KsVaQtaVdHImCBdmFP1YGAEcW
VMIML57Uwu80dAGPkyVFBWytEUQl6KiAr+R0fiYFSW++T3ehtUU5msD1ich98kQu
WR7fp12TCN6wcWs3wKWJKogSvtF6A+CG88/I1uyvazrJvG/OBEmcAk92bSQNSNur
5pxp1sMc9KbJciPO3VY2EBXCuomYMM8D8OzLzX4HCryXYpunb76eM2ovuUPrX7zS
3KFw8NV5JGM2vCiuUXxyr04f16JtNazoMiFo9tdS75wg4pyraQVCXfJr8ZR3TYUx
QjLATjvflpstTeM850ZhEzq0vgAgGDL54dDJDWNJkjw1/L8kvp+Ag+fwa5Qmekhy
9ZCqxZv+FUMd3zyx41kTxEh5sO2Jw4nHJtmWNBnU2q3l6bv3yRwf3VGLyI4Ra0wc
Srh/jLxOHT0yJWDsfCuNKXH1rsX0Pz9HKyr/QBZW7wIpm7VJ62hXcO7V0SPnYaHY
4dziJXpl2XidO2CcFtzvDFwFJ9YjboySlPPvy7qHt5JF4TxbdT/N/ycM1pWv3eCL
2763ZXmE4m+0fJeNFGUxU94i3nF+puVR+Bihfpi39pxc3Isqep13XqM6HiVshIXS
JsggiWowa0bUTNJ4IAB0DyuTQsaoa6X7SbpV6+uFxORTDoudxOo2+37mMbLh8QrV
OFTDVyAvUdkj+trg2x6OJVMMJyCQIMYhiGKB1q/6X6bZUdT98WZ1vJQA6iRUqLP7
y3bycNVjZrNEduOZflucd4c1fKCwil4XKSiOPM1vxI4wIgAsR12gHplXP/q5yXCq
uMv+UVNp2cD4Tuwc6+AphSasVJN4+HP7/JmWeHOVMJHNS6AvxAv1br8m4Fucegu6
zJdFcE7uQp99miUgPPgZKcI7LQZdimR+WUDPo6ac5HLi8svV/Q0DTb56TYjyF+pN
ljtGCn74d7jTJZUpKA3yxZevcUkw4N0FTj2CSiDfT6Lvn2zferxkilRlz2Ja4ra6
QG5ZyfbYhMJ84W5o49JmsyaU8oMr1vNmwIeHPdGBODycFdfrx1pC9utjtPs14FUd
wnqujzGHQS8Lv6spFtCrj/uAIAGh2rt3R9PbJpmKx8XvBTwcGo1oqGL9TJ4OYUXB
IIy/oOTtcya3csM+PAd/24nCF6IcVJQpi3BBO3bsO1IfYi3AD8CeYMSp8D1mSxcH
wW7p+NAnyJhcmuujGGBSi/pfeIDWirll8Q6vMR0wajJasrgpExIXsDjbEZbDQK4d
KWPvMs9kfC4egDsYSON27GhXBoORGkoYoFvALESeQFXP8oX65Gx+T+8ZsHds5/vN
LV1kaqCPo8M3iROqncbkmOiQXiN4lncl3i/j3IspeHVHTnbKBGD0qHFsxgzDOL2b
gSkJ501uTpHmMnGMlBq+WUl5K5v1zho6kDINVXHcD//zEKGolARoEE73mUTDzTWO
fn9ANXqC8l5B0iK+f2yoWapJ2NJfej5cCRb6LZvz5lhKz/WA08EU2MKTCeFA2Y7V
BvcMbFPbU0vFM+Al6CISdrRlfXrQsyeJPUnfhHfc5ROBYQaFeWWFYpOjwblpIE8P
pa1D/vbwXTL7qVf90TFk3nV/FrVrrHpt3YVQhewqFAgNA0PlV1JT0xRnKUK/CcSr
WdUoVY3gFhnv+zeQVqwbBWkbPelv85zC6aTpbRpUvCctJesIP9UIchQySqNsMOu2
QNAdBi3i+3BDG7wzUpNI18lAYo26NY68jQpvo/NUL3YJJF94HMdkgEEd6CzXQgTj
pYc0p9pwXmCFqgLTzDMHF4uYmcG5TM9m7zGQNAiiI6uClhhEhN7Tr3ZCmP0PTN9u
F76tuqVwi36jVt4d3F+WznRUjMBHmecsMyV6dVK7aibsAzy3etW6LiDZXVPy2VO4
9TVicGKfiM5b1UP4nfjjrA29bfk7F2wf2T7W6GM66jaJ4aAJeCA+aY/9PXp/rK5D
3eq3F7TPwFNQUPxV6uGfjBprfV6UloTFMl3UfQQ1nthVBNz5M3K4FwgVosDmm5kw
I5nt6gQKabnzUHG+I4ZEEmLEmJ0c6xT75dxjYXXBV6zUyZ8r16OAHTFFfIXgWzGD
/sHN5oyIMWMIpYDhqejtTqSw7ASYDdGEA1Dy89exr/K1v7R5iqqMo+4xZ7tagNzU
iTu3SGxrPXiOKpDHOe81dWTPfsDi3VZ057KzsoW0KPMSIuo9DBhjHmj08dZxgrah
b0gkUME0awl6oJFKscFfZRCepPiniciFwXMn9d61fCGp59dWL86LkPqkkIL77hd5
n7ZbfAQAO4D4e2l1dA33A/AcqgIZBDFfmyjqUofQO0+KzguqtVU/Lev4LTseyG21
mgdUr5gC9Va+LRHTwtdXi5z2ULSW19m/ezQlTrmrzshr1Gx82GEy/wGL5U7pkrRa
2CpzqX9nBVbSc/bEjfzTKrYQ0ad1pcBiPJaASj9GiRlCXgi4azF4LxaM/h1bvkK4
yV3AWTpIB9q1XWcS6ORbPjIh60pr1hbhFD4IrCx9LFP3zU3d/RbatmJtPWLpLW0e
zIochO5LgJd02IEuDWDCUMbEGpzsZPwfS4/SC7lvGWO5H/0ig8cIy2N1CyoSQ5Gm
YypDOx9jK5Qh/svJ2eTkvmKdPkUOA/19bTMTMvzHhQa96t1EJyqkJZxDi98GOmpE
3Tc1t0XYeWixzC6wVHD7j34sFIVlQYTlyoROJ4baiel1Pva7vlJjExcQqEuPxTpx
PKnTiERJPFqazcekmMFxcs97SmeBEBIvPALJ7f2luxW7a7kFa6p1CbgZ/8DYrDUc
MNGX291aL3DoWgel8bQHLxzfzVfxjLcgvuvA4BxQ00F+3FjOKmbEDRvuMxqLMwk1
NIrBVt4wBdYFXg8bqA0OvAi8VidJVcVpk9p1nqE7grVnjZZoCL1xkDPbA8DZQRC8
FnHJKMKe0ccfM2WyCNIlrpWcrMxWIeIuE7IKJaseTXOO3jsiKLiPaWRstxSpUFqQ
iYEuCPLrdH7JTkgxDv3/14WScqbwoHY0zXWGGheZgzYNrly8EwqKhnGDYov0KdFg
CF2j28Cut3Gi4vXNe6y1Ehrv3FBps0Y83egrewSH4IYLWKeRd9i4neD4pquNYShh
PYCmRG/cN4+B9VefLkq2aihrATNP6a44Oi8tYWEH1IVa17rNgcSXotUwTUKF6gey
sE19BTZtRGK8ls3P6MdSWyuv6/lRbqOWiq04rncpHjEJzqjB63BxVxWJ3Fv7xoUo
ygk+90YlHUoxg70zF+iyLBKTbIrDzftJkGpUKF+DzI/7BvYXVha3bgEWYmuDO36e
R0mbCgsclpTO73RALAdnCIC/l7+lBUueAz8a7qnjLWlu/cAdgN4XR8PpHcW7wWby
msR1Yp3PD0lZ40izm2fKRyiMlaum/05NCeJR/UhIxIy0CjnPZzVpLch9mrBWfzmw
iYrZD/R+Ij2WpMgJAQJn6cmpwtgS79TQdorNGgld9U6YbOtVZWxsNMcaxOaYpFTg
d1crhnpgFen+2JWs1SVGjLV1vCC6t7PbBmjNQBvPO4ZinTZHYl8544VxJzhXNtN5
drGJgRlZfYODSbWch0pbqmuhgQZZEmuxvSTKCYwPIpeBYKrXW5PkyQgJBb5YVybH
88Ml3vuiZWiCAu/m4zw7/vPTsAG/E/DW7K+YlITKoQABCUefLKgjOJA242/y3vUH
gQJJEwf+32xfhxcbAoDihnpz0csD1d0v+wldBI/lM/0=
//pragma protect end_data_block
//pragma protect digest_block
L5FM/kESpXQFi9GxVolpCakC7ic=
//pragma protect end_digest_block
//pragma protect end_protected
