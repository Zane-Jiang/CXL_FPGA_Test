// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uFpXnZPvlwxMeelMCR6vl6O/F1QiJm+nEAupuzYLJqObxNT7tzr2BLSU3kvS
1n30jDeVOoIY1CCx2lPF7R/DGrSui4QAenmDeVmtqmyXjeKNVHbniWBbsqmp
WP5UX9n2Y8U8CKx44G0WPFgHxGFjQcQPGfgJvntDngd9AAyHa6qisEzX5Zla
pnhp4aLlfEiP+YqlYDRyLMrMh+sKVEwPamWBghgcMn0g9c0fNfVLhiZFNPy6
hTYuZ6+EE4tiLsJskSuhCBHvbDFS9ZzMrFiVs0rEqKxFWXGZMVTUwqNhzI4L
c8teppYbYeHmSNuxUfhLX9I2BvnYi/p2sR/AOkOqNQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OwucRawYdKbhV8u8ITJfLSkcMggPDk0PYKSRFQmneFa3we9xQy0ErxvmNhPe
jfKIrbN3J+QyXZER7mKtLOPERNpC+0E542y6jDlp+WqBog6tnYB1MBQEmmFL
ypOOzD5hKF/o+LpNQUTFogjnvx0Mc/fVYrMycWM2UnUS4US+2V+LxJjKBJVq
ESIhyfz9GyZg5N/aozovNdBzgDoG5IqtfBtK9rCFO+3O3EKSgdf6tIZ9WQRz
jxTvuPIu8y94BqDxenA7npO5pgr7WHQq/D05IOHbtx6BiQjg40GlIPbvMn2k
3/xE5W1DaWSuwNrxzFkSsWsZiOF0V6ps1ASkhL1ejA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KYJxA5g6RzlpLQDx+Be5Xi0Aa3mJudCCMk7AURoeuJ2qEi4IMfhTjrmwNpSW
WWCGp3jB7xC2sMvYtbm4/5O1/HAjUbjZxfQQNUO1g3AUcBriJ8Q1U/KD7FsS
u1rKNTpnOhW10giubHz1dt3qVYN5U7LzWOR29it00FQDiFTlBiBNsVs87kOb
qAASU2PZdIE/E3UksvtvVQg37I6TW1QNZeYIj9dF139+ulJK8s65WnZ2Bs3H
4HSHXe+8h48rOnHgvF7ZytyceEsOK9fQl8r1i3n0MgZzPpQ6WefNmDkqtdCu
9yOwwsk/H34Q46cF8R96RsemNy2sP8apOJuppI+Vdg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ec1wEHvL1HXzcZZtzT+K7gf/D3dmKOigee4fDE8rfXLO5l6h1SRoUVjr8pix
HzG+cJNr4pmOjESgAm8tVRZRMeZd8Kw6yqgaI5FOYUove1bQeuk4mJaYU3yf
2gT+oLnwEO+NGVTGK97xCjO/jbCc0yTnQ5XHhCNE8gSFV03rEQk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xwODS/jNRQdutEFS2NpXgSeQtWGmO9CKJ37WdBpX9IUVarOExPfOTrzu94fu
xrdv/yO9PY/05y/GVFYQAWflD+L29qqrx6o1v9kWkupVkmDm3cv0cVFfkq+F
dFN26CM+irzWmz2QQ7fvWSraaOscGZcrS8JfPd+bjGIXusdnoYtcH+B++SID
t3l+PtwjJAGhIpGmFvqCtsura0sceVwpxtMuXtE6o8NkopxDR6sJiH2C7x4l
JoeO0NejHNoekOKVuuTSPgZRozwez+9OkI4nB9Oc1f3jqdRE+LsUyEf0Gfh7
qSfAAI3Lzd6Y0Mq/3u44pTo43rzJSVA+nW+4nO68Wp0BUYmPuEvSax7bs+7k
IyIUc4jrjgqksZQ4Vc+tfW+BLRiHXEZwYQeVC+LDcMHUl6ZkuwghD+02acnj
ovFOkt6cA80qzcWRAOnvhSatq44bsaAPFqSrdp/qZsJlxRWBt+HqtaPNPxjc
7Y0DkdEgv8AaBzL9Mc7f41tv4F9M5arr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KpafX/uERYcWTG8YUIQjlBXbchDRBduu3PXEcwizJM1L0VEVwerHZcWhfJFA
zPN22FMY34RHpPplbf5/aVQbUHpiU2g4jW3OkoXQXpyqg7mSADhht5Jups2G
9zSsVkehUt7FCjACEhbe/qkjqvgst8h6PzximA7xkxZzXuz8XOs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n6MScWKJog/Skh0Y+4BCKc2cxPLIM1tQgF4kGtelWJvcRZBHY/0iet4gD8Np
Fjcz5uJP9APpWl3poSECUck2Hs9Wfmp4Winc2r6wqld9DDZuIhkSI7u7qMEH
mMJGNGF6NyihgwsX+CWFnjdgY08E9XIalk16QM3aacq4Kee5p/k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1024)
`pragma protect data_block
rG+dLLv8HUUbVGkvFdEqhxdopZqtZIAWXU3rf4cl2uBLJkMoQkK4W50xk8M5
Txv18H+iO9761BDMtDuzP+/D9wZBtr74+15GwEy7pVJZLHRgYVKn/eaYNUE2
89DD8Fb4RtwWMmBjADrpeevDv+7qoPu3IEcsRzGCiSM5gAO+vikJCnJ/2rf9
vD7PtZl3z+It77W8pmUh2VSlnX+tu94oLauxsvy1xhY0yDaekppiPDfx1iqo
WGNsHU/Ud+25lsVlHPH77UygtyBL4M+VvEmeKvcrDjQAfsb9zxEsIaeVv9uM
Uxzn0yllv5kG4XXRZg5NIEXjEKAwW8ArEAuOxyAjkK+ZPQMFAXztE37l8Rmf
55Pcg9ZTAYY2+JfOG8DTVM283ujqClESsrhvgm6zUmpY4m+iDAAHhxZN2AHP
iXBYVI8j6GVftsSFu+FOnV6DKBJj19s3c+js7sSCPCkTV3ZoMIaaTfJ3cdY/
B78cpwDk1Q72lUvCWVJsCYbDvCtv4LFX95z2cKN+uUxHpneJcghs3vUGQWR6
adx4+NezSYbbCw5ExbL8LzSDpsAqZHjcd8LdjHTu3Kiyv3PRdUVMUsEPu3Jn
vR1chNu7RM+cqxWVNcnF0HOtjLR90Usy6FAfP7o0epTtzhNarXiFyDzsKi4B
97HTrBdWKeEH4CrAz23K01kZVt6jpOJbd8DFWMEQnr6c0th/dEsxGK3hBqu7
RcdxUoiL3lbyYSDs9cfkVxMMqQHWBjjPnPmfLrJ9MRRoOfSdsh1iBwvTK9YU
Otu4fZhIADUTNRcuHUCVgfqVjC/2DqQ+PxGJP3LzAXvt4RLgCfCZ/919IjWW
8RczUjtFtIkI+6QMjDMM1n5woMyqJSjo9+EcqfPh6KR4UBYTufTDMcwz91uF
R24ojkFusuOYUg5n8H9mo631+k3sBMD07XMhMXfMEWfkVvFYhoAlYY049eCZ
OqZ2yM0mKd3BMILqulUIlcmwDHj9p0gmpudh1Y0es6/rhPxbv95UvzHiSQap
/RGcMMqrDB59vrf1Hm7nV53oE3xcDiAN49gFgeaGbbEgi5EuNqmXh4MBAp1h
yFGUTSKVDWmWaHOCmPdIf93yM6HyZoKf5XXdzYPzT0cWOWzRQ6VJNBX/lGJF
FpQjSV8fK4P4y42BEPApDsOX61jTen6lRY9ioTQvOGpr/sWTvtE7jQnrREkq
F/B5JdACoChQoiQ/bfpZ6ddRXyxEK4tjQKrhxETlJcHH6NFviR+BPIgO6IvT
/9L1B6OtWObvnFyW82TOR/F+toPgf4aIsxYz9yqs1anWHDZhG+7DGKt29TMQ
djPe29yp9+mX0IMEIO7bdi1oz+agvHx8C2JXrhj9LWAY8A==

`pragma protect end_protected
