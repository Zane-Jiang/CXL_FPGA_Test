// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
UmNJbeziWp3C1TKSnBYomnMQmavPnOO8+xxtfqdpMOv8LvvxmpX+kwbf0Ak3XJC6
+Z5Pjvuexmrkrg7ZzwOBlCNNU4G6ibdX6UlAs1gc9DsPz4MmBbw1n0VAJyDsS6Df
CA41m7rOQ71fkdh5MNFrLi2zdXJp7rA22IbGqnbZbB8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2304 )
`pragma protect data_block
TZ28zhxh06Wz2J+bnyQiQPWP9ItEMDR38uGwhlr8ZqCLKT2vGayuokUdNw4NqOEv
dMTtDZ5v2q/2VATNjc2FnN55bjWwHhGWt9LP/j4v2B518+SZjAg85C2uxjY/OkDw
AUXzZ7BJGKJSk37tecD8JHPc/0A1hn3Tl1X9qBAW32bvyjzPElsDKpBJE7nAl+Pb
aKoso2zBuJ9NpNM/vsM92OqiZV6QUKAWlKcz8FJOe1fIB7aroSdvHSO4o9yJGFGs
PO30L8JTqrRK8HihnObK84d2N5zLvP0aWFv5JT9vUSdPUIG/O3foZmkJ7UXOcps+
vOYWmOQ1+tU5uBV2WYL/fRGo301IkxgSiqrnltgQ4Ki59/peDSYLIeHy2MHx6DBh
AKVJ4vC5zNv/wiGn0DmsoGv7mla5ugLqj0yPVx5r6f7CIr/ShWYcKKfCeK6fKpR/
0vvR9gJqMWAj9tHOTUqpHjfbY04PzdrG85/sVL0kIUaBdSYZu3+3ItIE7zzQELZM
hqvXz/Qql0BmmPTBBFrEqGroT/k0P5QzKDZmYhV2/tafHYY2fPLz/+WknSPxwTef
Py81DhpCX0z9VWoT91vL5ka6IWr978MTsEoxs9qtF5ZBVzPBl511Fux4GJB7Nk4+
+Ksonbe6pVDmFHwS8eP0AhaqyviSsH1RPACUFNfRO0k9fEyZiK5wOHZNozrAcLQJ
RPie2L5Fuq581x6dzn6VL1ChHbfj5JFDLD/XajNkQ4YkdowsV17NLClHRSt2REHx
mTmQ7u81zlm8xDlDjCvzg9pm1SNj/bI4K4xRjHoVUlYeC3eEjhscgJUJgLdDF5jN
88uq4CInnFmTX/vbIXL0BgYJt+9WoI4cNfa7RJWXi7bV/1jtoISLoAXyNIjUEaIs
dirPx/5WooNiIvM9f6Bf2xIVQa2ip/lNuYZK84LjuEGLM7dYktRkqrpIe7/m5p3Z
nTmVqnY+tdm5Pq6x7/JjiNSYAucribgda0Bhh91rtv2WM2bkUdvvN8uHuch3tlh2
De9YPOUI97y0Hwq6HroM5esk0S/I+bqWUiIu1keS0f81/TI0naJLOUyO54q29uv2
mhGWOOn1faH54S6G+qB1oR624yjKWhDcPeRS4hXehORJg8xm5HrGRCfMHTtd7g9v
q71Ckw+FZ66pGsKPgV0a6YS7QbszgLChDvMdYU92gD2tZjYfslGN7Io3cZH9UvEx
HxQ/a+KQYuM7p7B9YQryULL68CrHVpyCJP1WGPr62JRJ3s/v/4sVaL2qw0iAMK9p
M4RKNYc4jYN/5BpakxbBUomrWFqhnAHE5VLOdS6dqHBIB0TzpnTLex1Hv1rn/0Db
c5ps33iOghLPeEQHZabFQAgj0jlNfOdmYCc8s9euP8I9O8q9gwWj2vYeF8CoBj9o
JsiCg3qz/93yTdWQb30lif5w+SFhz4dClugse01xf8ASggH0CGPul1ExGRri4IEw
x3DLr6YIligjrQ6YjSG5/5n+chlh5OVjUGE9dwhZ9rmmVvkevH5MQ0hhQPmZaqTy
tKLOmdSzTNkbxKkY0IJJS6+k9Mi8dRCB97afKSjT65MLRCmpEs0ONJ2kBYN4VnIi
H0gfRdwzh+O+KMUhrP7Dbh2UYKG4AuniEeu9P9Vfo66U2W4HjOpKTZjX4ro6UgsT
O8XmBqSlGv6Vr/YI9Bm+eVI5GQPWk/LsBf9p1DUgGyqQwvLi/seOI64wnGqp8Pgl
zg9vqK67KkU77IBXL1v16MdFA+/aUsDhKXjlGCKDMbXLeealAmgUsYJ/VN7fdmbl
qI/+yrZgTyYXs55DWKkLdzI+sZDZgopr77lxoXL1dm59jwndgSo6zONIsrv/VKLl
jm9sgfrNjytY5ZxzdtuQadht5jX2Y64UXx2UF3HqD0FUviTnDZWLNeYALH309Q0N
dDbldh1u647ZAbiKjmuWQcuc9VLBIgfE+lOMUJzWQvAN8HM+rBRDdZC/wWeSIXVk
/jz72HcrLOtCMVddqzQs3/0zN3NpAVcEG/u53ZhvsIjgFIytsghbM/1D7Hu+mxHn
xhfkodNvB2HY9xdamkuDXiI5wLhRzb7KcPaOI8U6VIuzv98O5QsXMxmqAbMFFhZU
OCiRQCYMuriFv46EICgketz0NsIonI9f2dRZtJvCa8jT4hXRffy/2zzRigunWIBO
JqzEYEECoTqpIWaDeAHmruh4TfoGJF2SPk/J6u7g6YE7p8C/fM30Q5qULQFsrVy9
EKIM70maGZ2+4zSb1xblrSJAgfLRjqHytAy2/Kqwx5AtTw0uZB5bgGwK8fUXyWjQ
muTgb+fBQwxAQUQOX+iMDNHu2nj3ULZtvvgUoryyGk5CpwwaYUWTr7gGU7BkTuM9
GcOwQdPzEBFdY34JNELYWj0d9x9xjbcRKWq9gVSAuxqNPx4miAR3xFfP0oLpjSXP
0WxBatAFlY+szMJl6aB/GTau/jW+Pn/dxEDr0fwBuEAUw6byxIqqZlMmowlfjCtn
YNx9JKl60C3i3WvIoBkHuApEHhqzmWvC2hVmwqxftlYR4TpAib3G3JR/jSZ2tsh8
NpDVgWJ2NhKA7uFqcUaABpADMfRa+mALfSuwwkW8m/k9SvzqF172bczTn6BizgFn
y6GNusnFLyPwku6dgiIihRuwm3yJkznf0vICMke0m75C7JeYcWUa2T3KYv7ztvXH
Wqgct1AnpmVyMJ07T3EUWtS28olexHYRHwLxItmcsoR2UyuRFTxCfJDNVb0TYMSP
QhK6YWKeWlcyUKBGBWRiNDjmYMnRqC0e1GauSWlb31elNjX6EfnjwI/hFgcehPtf
lgPUV5JdIfEIDVkr3OVyqzYGZTaskJKydm7PzJDxNFXdv4VeyaaBarTxM5DLUBfc
IrYB2LXumuWM3WQw4zit63wdhQBkFYOuwHbzpU8zPtC4kopmFvtQhMj/jodUqrYM
NDIAT+vONCbaWDAATgzjXNjUzrTsseXES0ZncWnTBq2pC6Ce5PNe5ZIwhlf980+h
V6q7wXcCTYKHa2eX5Q/MlAsdELouyAYH9hidfvX9/quCBN/PZsLMaiLLjUXlGjpm

`pragma protect end_protected
