// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
V8bkC0MAHhew/6kdUcEgx7/Oeu6W2uxUy0+7pENIct2tXbr0d1J1eJxQa++iQOkk
W6te3gvdNPWhym5GimeCdsDHbhBvT56lOjNf3yqn9vC8t6FRdljW/8lUsgaYxb08
Y7x0U7Yhe9kfPrCL50ILJ5R1wz87+4R9YnbleFekhBJEh1X590KgVQ==
//pragma protect end_key_block
//pragma protect digest_block
dAdKjJHxjUXq6BRJoAJ+sKFeIQA=
//pragma protect end_digest_block
//pragma protect data_block
8aWeQJUUOXeDDRPJC7EBUVnYWoSQINkrbrUyal8nwoUNiYl98A6ZjhPbpe3pt2Q8
3CnYsv6uMSL3PLFWXxtj/NAusY+xq9YhnG4oiqXbfXWqURUN0OrqryUUKQVQ+jRB
kjvRYXOHvgojkAqRws1IA7CrQIfb+azt66QdBuxJAt5MxaPrWxdQSJDJAycC9huP
Wlsr+4B1M66r3f1ngB/XMs28P6Bs5Tz1LCcV9c07MkOhHZK5upIEAAbr9iEToxe6
LOJVTxqUKxc26loAtkMgOv+ohnnhlNF9yi7kgIexQ8enzDWocE8LuopMgwFCcPO6
ur5ODdcEFKeg3DzQILdJ9QFasovQe7iBZ2wkXv95vHjOrT/4iC0qoH5WJ+OFL5uf
NVE6kNJJSLqWBlYyKbYokKRZVO4LYMa0rlYL3M4x0ZgYdrw/9BgnR1WWQws7+PG4
0Yyei4LhxUYznGwIm8Tq2zBJAU3IatUY5Qt0nuK7GBwgg4frZf9Tnl2qpAVyT3AS
n0himEzs1FM3qypqk1y1u1LmBgFjUB1mRz9fQboAtleQo5LnlJC6ZQCwpW7SreBp
4uAZ6zPxhd/Bsg8my/f2KEvb6SWd7HgZZlY6xd8XCQHQwTdasYdVWirqqg/WMQLw
vFPt7x+xdctY8bj8L/z7RQKWRhTCqge87X4y1sXc6mMDtKVsrd4iYEY1OjK/P7p/
EWisc2XTfMczc/8DC7X/muSvkjd+Ng6jOpq+HBHPUWLN5ljnBrhMflZpYmwCHbkb
UWa+Gfp0g8KACNHdcMfyJ9UEKu+xQmAffQJ8mhm7lmQYexc5d7qis9781l3BqfGs
9s2m1u6Bf1TrYTNJEcgOhvXPI2HQo033riAKLqB50ivEo/e+uUo7dtkG6NBI576X
LNXw6iRZnUESq3acPAbN+1hHXp8BPoudwyzVX1Bx7cS8XRxglR75oVPeWqk9YWD+
gOx61EqcKYzIMhyMYdrEMr0KEd1eCQUVVJFn598xFHQE9hXedmBgmx8uk9dhusyT
mc/O1H/QXRwhHvfik3+TBjV6/fxjqu/4U01lFGrnK1uoLgJEA2PPyUN8joMX8siQ
Q+c9LAbdfH6jLyYCYL9vB1PVOX2aZY13ADRlW26JYEr/rMO9R4CUrLEEItJ1QRhy
CDvIob8p0uUquij9VQdKnFR7pehOMwRMGulSWlCABtJiaIQ2fEF139xbf55oM1ui
uD6DDHKzjCWq9U4tAK0zCRBR/AWQklddy8/geJf2tsWNfCTCW+I9s4KB0gU32tyP
2NUzwiiEhb+DsVOwDYJqjusoBnrhiEiLl230T65d7PGLuftMhLfQRuiSNi+93Y8v
lMfQKWKcMRymvZhLMtbfTN9iC5luNwZU8JMwxrhCEedK6xSW60XEyBgmdAPWmIIo
m9iq1PMjpvgus19ybOSK9HBYmJwwNNVpJoAGaYywWN18wxMrFJcp5+GM3p+dCmVs
kGxQeGpc+rfH+NUzjXIrVzd69hn8s0Ht8tL7u14xkWWyEPpLBeuIgm6Nba8HkQLo
knbtvWJqHpzrTRR6b/LT7sq9j7FnrJiGJ1xbM4yQcdfwpehwhi29xYYL/eyjdidY
t/CLdxbX9e9v26MVmXRY9mQei4NpXkvHn4ZLYWG7a7fCtIoXOM7ze2vHJHfT0LeY
sJG1OSvApx3LMeLuJOzh+V26oUAkSVeojNExO43A68ZPucBomFkPZmMNvMz2HSlE
aFCoPnXIb/ZlmYU2nLIXDEko7WTL0buBuJs7fyWwOdJ8rTNXnBxcdm3lBKmbHajw
olUBNKTHn2PHQhFPOQs9eNO7gW3fqUYa3pDvcegPAs1whtmedITHNmQyDcZLfIUO
6qUek6ArdE68UmIkzObRvS3MCbzWt+562los4gLlaO4VkM7tiP0Vi1viNL4Lo6Us
zELilzTDsJmEsNXjgqtFe74CprE6W2tRpa4lNllu8eP6BmK/3QXdUiK+pqzFRSxb
ikLi9zNVbj7nqX3fRKIJ0dvJgfq96eqsfElngMSsHzCk6yTB847D3xJb6mGKA9cM
F2Z1Z2YC4G5SbhQHWH5SVj3lfPBH1T0+ArXaEVKTIMCMeUL6ou8CvLR1HXJKoaDO
9H+s7TcvPumQ0scQ4WZyQFXyUnL3bXe8NHENKAHxZevlOdObm2TxEBECiG1VFDgg
Ov8bMyND5DMx1wjUBLNHjqbViFkxtGv0+X8CL7LKzaug3UZOeEUpri9CYP12VLKf
m0G9wiprdJGdlUvMNeqKY9niSH+Z27sO22QR9B9dnggX0QvpnGMuNA4O6gQr60lX
gVq98EzAL6mTHfq7t8Jt/7GJ7WJv3WnnkZzztXLRyjGNGgzKy2hWjMPA8RIxXcqd
+eWoilCWoeqX85wREhOxSc3MmMuwqjqkCVDL78selyF4xUEu2N0JyDjBYCxaMwzB
bMxim0B62kq9tTw1JKfb7JLBW1limMXfffu/QvpQnHL0jOTd/EdA3RDbftiMlKUT
qvcIRwgkepiG0nWtdgX0XQap2B1f7vndndpdT6vBc9RIyrZ7EQY07MOeINj531JE
hMfnYi/Ho0vSWEkoYlI+Cb0AdZxGI8+/yK+SW3dw0cID4MJk9nSuyi6fooRgmz1H
IMfIlc8DLIpvJaJvnFdtRS6o/fO4XtAEBcfWxyY7OriPZ7T/IAJ3zAyZw0MbS+bs
gx+4RMQpJkNDBTX1M+X/iXur4f2C7tAiggXwfzzUCAdu+gN8NuSUjdcxpElA2MOE
aRa8gpjjKahaw46tcjXyCcyNlNIR7W8TMP1IcCkwP4t7nh2ry0eth94igJI6vOzL
2eNAYCw0KgX5/vBe7tzuUp4gz4XtsLeGRRX5CGQhokkT7R7S7R7FrB0AQXekvlaH
PwyiKB0OPAKL9IIn7tFF0VbomKabcKyVtrl82fAyw9GisaXEHt5O2zC6MGQAid6T
cL/Gv6q8ktoWNDFFwtk+x94Yd4U3bsvXyhg7qlicDTKUwhIy8ED1ohcYPQH2xZyx
A+D8h0R1OgAmR8zQqf26fGxCS0726P41qPuq1zoaO6etAUMMbPO9cOR1hhh9ZL2K
koUckO5OGVtD8I8F2DMKrgjHwh8eD9w6a3EBhqCDA6WIjRLt18/ClQk7RJ5yb+I5
Kyl+LKNEN00s4tUYEodxJYX9Zg6Wlk7wbbrLacaoE7hpREgRqsAbc99+kINUD47Z
PToQ8RytgZ5qC/JanuJqORGvhDKd0WaaVXsAnBuCWBFl9Cx4rxBNq/NOGB+Ax1a+
kefZCds+17ZUEovm7+qmYH5HAT64pfMoMJ0FBnQofsIX3gmStG6a2ySU/hgG+93L
bpB3pe49XAoR3OktV8kf2FuJerG4te3gP+VencHNy+d9I33LX/4UUJb9QDSJBc03
Y4eV+wdwW9sHkQtj8QvvAuBrN1uxOIs48GsSWa+N8LEj0eP85l9j7sXEfm59tv1Q
TH3pBpgg9n9MEHmdvgaQkY1udc/6lJZ+JEa560bHp/SXnvdhVgiM3QKVRrlS06Ur
9IPzHV/u0bcep2Yx8BSiletQoBm7qOlj2uEjHW0PNoANOlIQ+1/VlQifnG9Ot/VS
K3IjHFpGEKOIP+YY2KsiImZT5Q8dG+PZY1/ohvcmWsx62gJJ/Mu/i1dvpQKK0EcS
YIW6kJjEgm6SX61DXdfBiEgD5m7igAwRMeogNPi3DN4ON9FRJpFIcL51aWLYHP/R
c+lN1QDLtwRon6NlxG49XzUpiujsTZ++Sf2sOeSGv2c0FGAZ37fuiiBmFKktRU6w
qvcSBcS+Nv7prmFiKHLbFt+gbg65MvLg7EwbLJwleSidLam6cnWQlj1/6Sg+Ce1+
elanQ7yCaB2x4jvPXG9gyts8JF2TS2sCVky9TSnqkBmys8kw4EDtqmp0DGk22FGf
1LgGJGbK8ntcVDi04zfgGQyvz7nP84Ra5A5iAYAnStin15MYMGdUmrYl0ZEiY4Hb
kEBPnd4hpI/El3wCX+6KuwyhjQqKs0STlw6KwibnryxFTi/Y5m0YJJJdiQ8dsrdS
g5aHwAzZQBrV8BEkw1VipFB/wWiB+D4V21wlvF3Gb9xMc7JmtsmzroFbrZGiqxAB
cOIfCUxQGTVE8u5ssg2tB/mBHrmWcQGIufNvGPI/CYLYbwO4ScOsWuK+gZ6Lo/Dp
lL0BsYYLHI+txqDNLC17O2ca1uw9uPjt99Ob4HHl9flgiVd6sGQJF4kQThHtGGqW
FKdjmHQiMRWO0KhecH1WqB8b+uwVf2gy+DYS0WzQZ3FJA8KsBLxxOp43KcGOuNz3
S0g5ASnICvbnTswiBXFVQlVvDZep5hjSXVr05dQVaTX2RG9nn6qyc3r6Exr7fi3X
hfkN8vVq0yU3U4VuDO+6nQjFefvWFlDHjtLC2IfYfFFLGLN7QcIPsK6HylpGGk2k
f6sdBTUgnT/tFjikZfpoQep2erw8PoC8Ef2T1ZCZuCocDF44lGhCkjo2VFZHAYYm
rCNdKKWZeTXtRwb4UOscbwP5+CtPe6+JDu7RU/sGjWHAEpXzl/m3COBkqRaihYzl
nSHQ3HTll9NIOdlZmVcIUVAn+moUJTnbU3ZflZhX0Y359kEYr4aq1jmh1FE+Hy1B
z0dGd/qc5fmQH1gXdpwy+1SG5F1xJf7p/zdCPChn9jUoIcLAY+O9K6RpUlepVY9X
TIeFBNUrEwuw4NZaD+I8W0T+C568D5HpDgnAyP2D5PWBXQDpRlP1kefGPed/tTMA
L1a5DrX0YkZivaButOvXh9sLTv3CeRZO7/wYLmppyT5R/yoaCr+nw5/eWPAZ2sQo
b4cfZ21F5uQ5oPFm+NnB+umtJFMu+ksRoxjzb30Xn3u998XECrqWCbmGZD8amHPs
Z+VrnVQrFpCCDeZLxhcCUVBgcdhg2fAc4SP4hGVxy3Eq1/4/FjPUZ5xI92jBeAH9
M6D4l0Znt5uFJIqMcHZ/v2bns9O/f1+DApJTHi5DYwjMQ8YhV0ZXohcQR5+KN6tq
NAFpicHyTD4PnDvr/QaNtsNHWzFmMXVQq4XZ+kfZX5dzPGiR4PCmsG/5DMMw5LNF
WNK/Q47arLJNVkeVhpKSP402fvMM2XV3mhs7oxx5FV0pNY5qXMjiLNAiW2fYw6d4
+qQHvZ2jqQk5U9D9uUfpMxhNUsropwaM2IZlshkFzqHNI1Oxaf8spvmu6HlDMMr/
IY8dXa6hrb/f2XavvrI4qEU0ZYTEcnLNgoubkR+QaYytai7zEgNSUifyQpDMtACP
Lr23vUthlPpIx6zKbbMKQwko8HHWMJsTy0tdw6PNl7atT2ryL9RsohAfIDOTSw/d
CgHuWj8vngIKlQTbLTjscXKzr+OVyKlT7RmzzjGasGP3xCStu4CuEXUidhXilcbo
weFQavqJgbsAk4Jnyo/fIbiDNjfCscq1lYdxak+6paqktJHZAv4FJWX6Ow3TZDsJ
uVuhzpsST0Uo1jXEepqTwSI/70qeuj8QzLEqps4J473hf97va7pYm2zVRmbYRJPR
PvGYx2+6ZXm5RHP0Xucr5uxyFYYWAAjpIPIYPeX0IKdR6Q2zppLmZ+ehoRBYNo2e
kxj2EjSWToS43h5/DgLNML25ONeCOHTQymcg5AQkMCNpO5cUEwdYjupBnUi1SzUs
fCyb9Tt4ZWzSxTQUsK/Yi5CkT50o7ZhNvQZ0FUSY/BoWJAVd0o1vXtglEl9NTOLs
Ih7xJ1lZeAIRWQmywk6cOPJ8muts6PC08V7nnqt1DUEID1KyZHgwSpzqSjKgwzLF
mTP6PvB1Ifv/nlviL5vExoteHMEdhAnj01qmYAlbYpBe1Lum6V+fuXOem57sPlNQ
NWovLeJUFLeF2VpX3/gff55rnGUD1XGPTzSp0o1m8FXGd4CcnkQapSuevcDT9JrN
YZBWR/v5DEhSlFjf5ltUWUN90kxRJcPRItnP0vEXssH2v3Gc5VSX8XDE2oNwrv2w
esO7TWbQ9vtZJ/7T8MkvhEwWI5yUenkHDCafE1X3KheAN0wAbJ/rBQ+ZIsHOEAaV
WAYgOPP4paQOQDMjELuyWbBLTeqkDGeZQeqyxO3x7gcSejN2DgteeczDE/drTM8w
ndZzPeYu1+A0fyHedTYBSr6dYllZaFd2vDIjAmdAWYBrlER6ZC0eeAE+ZvBKCf3M
p3DeXODx4R9iureQyWtbNCmPKn4c1XhVHIGFutbs/WAiIP7bR3kK9Hn03YadZ895
fDDsEUP1e5TpNCNlxjsQvDjME/Rlw5ecu94lRKpy5oS4041cJ5JkK1nB0TIINQHO
Vz88R7EpsFxDgiY7+Sox/KcYwhnDOSViMzAPHxD8c111+zArwybLNJSgBAwcMHl6
UwTXWQSu2sSuPXxqZK5pNxc5xX541TNXcLhN/oPDA4dZjQfW+hyxZuLO86HACym0
n/00g325Mnh8wiY9TRHWNGasaQJijgjMLTcD6APhlRSYTP6YWfF5Uwwgbex2C/6p
gILdqBd5tcclSt/Fb7xDu0iENyL5FQ3dFYuU1U0w8AFIWxfblNNYvwiWyVETw2ql
X2Prib0vjoZNNku9rcc7/S6qjzg+LsGxPTcNULCGs9TOgkfm03uqGdEH+yYme5xk
Dzv3Yzs45q8Tv9mQa6OYaZp4BKCBuMJBle5Uckycx1xoU82p06SdHBEd1BOfwLQC
uEbGcLt8epunx7/jv59cJPM6b0yLD43FFVyDAcdqqfnDx89AfqK3cB+9aLyd5qML
vzGS0BdPsGCbTgn1qS3puCtCMyWo9MoITtXtqCd/DhXhacadbztoNqOvrArNEOQB
vyv9QhiQ8JJWBHuVC3637KhYqHppb2rHhbKhaSVQUYrwJkjFzvyC+UhlXs6visxF
7MyT+jb0oo7q+82wfPtwvSiXcVOOVyIlBtWKAwsTkGLYM/jrZLzay4uQp7QSCyjp
NsnFSPEX6fbo8S97jnDmgbuupIdgtL+BoGOOo9yXlpw4VqTnKZGiPe9mtiQnNLmI
8mnlD24hqITpnbaVLTtKvYAdz/CbuZPFF48Oy/FAueS4lBR7Wjs05EQwFBRVXJO4
/FzD+Vb1sa/rkNJMA50TEtPN9+RmtBJmOozYGm9gxLB86EQfCzzK+yGVkPv37JSo
jS1heel/0wb6g3hATr/hXU2OVMH+XJsLZMzzJI+E4Aomg40gGNFslzE43yq711uX
bxTZNDWQt67BUIf6kbpz91n/oU5z3GW7oNytVBlL2IaVHER300T9kT1T31Es0Rqu
GB2z6mkvTeMc+Kl5VRvgeVE9WpsnyJfKslQMbUkJkZ5ijdSYP0u0hMC7hikKsT4r
c1lvE3eQmOm7gNv8KrGcvpV20p0W9NcS34GNI4OYuX8mLyMOnQe8JCvLRdkas/1s
WlrlPDj+LvITGKrMKsRtmUpnILl4ubbXt+ls8bN1Nbbt9vQKXcb7rN0OrDQ/1Pg9
gFXZ6vtRveDsbz4d8jhfDpLBLs+vBfT8+FPRCXfq5sAoy8UqTofHCiA/qGLoh54d
xefa7lCVpXDZw+EE+K1rixUD5m/bgU4VQW4877dZ0JR/EHbLtaGRWDYFjhfaUUFz
8kEuEhQqhw/izbrsDLohHtwFeuKbwis8EYg1Ja1pjRpTmmtVv9w3NDcZWk9E1WDO
TPIH+BElKX+8AXltzcXeARkAG12eTbva9Lqlk+0Osj3WAZJ2gkgVLj3HLGAv1q8w
lwGRN3EhYJtB/yc7ivRoyXjMIacMDcuMnQ3pGGtGpMUwqxmk/rENZjlhysF+1k75
N6h+/+Lz7ctHlbfqV2WMpAjp0Yv7M4xJaG4pUWLkiP9eIx2hPAqy2uXV9uizPzFh
flJUEaZflIfFRM309aYASlPohcDrSWnuNEh2Jno3Q4ycqSUZe3pmcxJ5udQ6RSVI
RWr0N3vPptqmMiKunzOXBhNTjE3IC3sMr9ISZldOqED7ghe5GeEM5bNfoVh5p02d
qNBwwbH57QZeHb0ceKL2JJkZc76aFWvFZfJ+feDz+nuiQiZwHiOhA+eH7mlTHuQZ
8pWWznLECjHSVzWJ09UmFDJEwILDscKSXjRP7n2meoz76XsgNcx1dqNd+V+g1U0N
3ru38Y1X9RtMzkEyOmVj5JiEsGr+YF5z0HfMav2jPKyAX0EnT51R5Ct1AWuI3sJa
SjRQPvwzRKcTsrUSSE6ITK8eYIK/3HLLwSjY3Xet9awM05w1Bm5+vD3JPur69Mtr
OCZS+CO4d8H/6lf6B5UrQaTD6NfozmDvJRPmCtkJf9M5/mePNgsgUug4/LZGI9w9
eqk5I9pu8Tume0bQAmdhLiz5hV0q9DZzJfOSJAgzuTDOX+BNn+LS5M2XkW+EjdQO
I3277QeVL6bTdbTovTIYrmXNtapSa4oj4StnTBNLkKnsFeqRO9SRI9c4+OTvWhcX
rH3q+v6lSU3XrpwQ3gXI5yY+0GaX5Mf55b3aaUT5TR1wgIA60ZaRhX0q2MUZNE5M
cPsAWkNrOmVMomWub/P2TEa9PS++M9aHliKvKKSiHby+MGCZZLnYlIJ3e/f0ysy+
wugdFKuU0AFvtF8BN02ALTykuTpRWND9RhW1KvVfTXLaMmA5AxWCIdWjIDaRnWJy
EsMYezLC+odTUN1FACGQgIcfOEv6C67+doBAKSqHXRK+bp/bEkwg3+YStVCerXMc
v9m2flhAqcn8xmUnE5zS6zpkMBFPpiqBATd0Cbsa1lPFu4hBG8jpxUiyY4vIfS19
BStBNE9SDgV9CokBNoI9CB0fFR3PPN/qagUoishzo2eCxiarsxvO3YAPi2+LtuLE
1kBSZ3jWpRrmE88F4s2bPORj/c9MxgoK5/PH4uxMxoqfgU/oYcU/INOdF/WP5pDA
dt0CNZpgLnyzw8eesUXGc7+aITyxRr1vnTaZA90Vp5savmFM7Fg4y4K/W0u+228U
jFpQsQOdRUvSzbGbIvMUawzCcGzEUuTAwuoEh5vvgGjQnXkjWjJEVr9D5ezqVstl
2kJ/pX/GgWwmkgrgA46lBbw48kev0I2lz1ZguEP/HCDFJYCtLF/4MxOWNAGiIit2
E4kUrparCD5spfGbHGhkvwfCAUasWD7ooN9rYal/q8BDT/PNnIhqBr/pYclrxMiI
n9hTvoezm5YqR2SCRwg+g9SptnpyO/49DJK2dJ7NKIGYl1FdqqFkG0PCI1Mnh1kg
YuvsG+ZVQi+Ni7nl95SQhoriK1AXIR7yUm177iFuvc1Q6Gj2lY7DH4z2y1dr6WAx
CV4wCZQhCauhsWu4kgjosyV2JLF6WiSIhnf3U8uJ391LcVhq/aqej8x9t5VwSZuK
Ek0VcPx4N4/yhfC78AdpL0Ue0eyrgKrXxd75WPVAmziuJLRjoO0reOTaWM2AyqZd
l0koerf8plBao3RHJ4LKYAaXwHkVOTp/NSrDvdFTim/HHpYrChOJeYiPPnaOSUNJ
FZe5GtBPdgcyoFkzcT69rKza5T3vzzriMNBNCYoEWNRa6NaFsDHTs7wPjrYlf24u
LxKBgzbNg98pEkCtbszYzJzLaFfPhCfsSiysC+Nybq8VmgdEls88ukuh61Jtwuva
1MA3+UlZCdVuTIh/hn8A52Pc9ijs2/vHduzAlHilZ0SMVuHIxVt/8qgi5wY9jWJW
4rA6YnpdJ1pAhdsazyCvyQYdTUFT7i7t7Lbsb6r5ancLH+ZuRs29rZPzN9ItLcVR
1b4C/0C1Ywgj7QHViAtG300PirKUz3kNQtwZ42RyC51JeqqBpvSvc2csaYuI3KOq
9/fzr2G5lRxjnAvUK7qrtxborvpgWyGkrVeUWInLiZbL1Y2pkymR1eUB0Hg6zqvH
T1crd5WFJtPtofZycx2ZKq0zbJY1g1QFbZx9jDmlezrkzejvybfi/Z91vhCxeYSM
72+DyrjeyB0RoxPJBowz0rfLuP9J6Lvmvri92iBpc2uw6n4vjEwrJexqbrdIPTPd
GIj/4vKNadaTak5BUb12mmxMcjrI52zjQOBGlCFfGD+nn3ZzWa3VDcONfkv+EkdC
pIG4V+MyLqeYc3cWl9zISuv8Q0YBUZrynz3qEZL7/S4oMicKJyKO2K5y6QPU8yZ5
3s90b7Cjj8kcWoZk0LbW++3Aitq7/yQmRnc3bEe7vAr0DtdNc2pQOuRMQpxmRe7n
YBNUTD3KcLjWUEzLsHSmD/C7yIXilvs88YvIW3rzGU2jo7gTB/35CS15lXRM8BeR
9N7Z9cSHybHKKp0w7l10SXeyjDM92LZwC66bK7wU+VMjgoZCsa3AYMt99LqUEYZl
Gfkg2c85/kyylNmR2AayOVdBjL+ZSmmZNuIo4K3ffKCTk9kpJz9XW2jdiOuBW5wk
EJooONyaEM7LIyFerALVicZVNXnhQyjZgm83KxhCcPkRPtCBGp4fwnU70btjqnbq
opoIviEehgsmPGOS++pOR/RRG4CKv9WRlg8QKYc8VJc0Vv7WpYOBgdKY+XaOfMBD
hMzmoCZ9PW1XJoQ0cZxi131kCKII8+cO+K9bnLckZMND+cvvOk2UIKbmWl9JZcoO
DUYAOQe9ymZrKbTDitnl3I8HaBuvQe5zkex5ET6x3VVMFuaPUjaL8kFtUD22sl9f
NCjnk/idwudEsi1sM0rSUlgbTcCvByMqy8VUsUWMVMfSc6CJAHTuUNJs0PU5LLYR
/iqBUx4ci8ZWAQ8tQx26WOq7WsxIL6KYEI80a84LkphNaPm16cu1/0mD4BMQbGfr
w/PvbOvojKJFBqgZ+ezvLJw/K1+Ocx5vN8fvmsGuUhCmGIWOgfn/b0QcbFzAemW+
edrGHhwT4UPfMDCE8wJ8XKdvjqJIp3kUJpd6NDssMDC27PZP4GlBZXfHDHjz4l+0
eKKMqKo9Jdt6Qrsi+rKnE1foZKy+ar+um16AYFIuqBlIEfolw4W6kB3BbCoLnq39
NpHAMJWB6XNjwYTVvH0oNuVV8jgHdrLlU+Ub4cRSQ3iz/ZnvShpb3XHM4GgfnDa9
hl17LupEv2ItBJIAXpz56pmOe1oMUBfYaB0TFqIHJsHAs8/uU7ujbDw/UVZldgpt
LhRNLfIqsYcP4Vu2aW+g+Qr4AyzhXkxEYzE8aM8/zBnlt1f+Cw+nTidZ100KnwYf
Ir4NGcB2b1cRbuOwH9HB593Z7WubZDTKfwg5GYfAhSS/JtECQQQIreApLZKd8cau
OlGdUelwhoj/ncIm/v9hPXcIy95wlyjSfoUqSKQNt/2a3fUBAqZqvOdfwzI0uzkN
MVJXisE9a2SV5OvvK7H3BGFDMfarYI7r3Uk3yPfhOGCDOQNbzj3NW13EHtdB+hj4
i0y3b7OWTOE4Q03GU4mdgUYIRnZltCaqiC50k8ebCyDhmSHpsig+ao3PkBOAJ7RD
umtzUN78NidNupI86Jkdi1xbx7ffDEozoWUjITGGO+3xzzARbEokHFM6UgbUpBhb
ypfVflWsFjWKrPUqiBsPgDGnDuwE7/oO3zlkBinrQTavTr48dsjkF9tF0GfhxJ5W
3Xe3scRf1P5CpK3PBpTeaolsUsBp1rm8LamrspXIdj1IRYd6Ov4q9QAuCwGk/e0c
yxKKW20p2QBvGkKvjYrdTLXGdNbV4aDCkDhBYAwuU4JPwMbA6AM0zH47QnqJKFfO
+vy93uL/vm2lABzY/nT3AEuetb6tGxdib5q37oUmPu15ezYObQDA9IcT+wRsFacQ

//pragma protect end_data_block
//pragma protect digest_block
YbH2m5O5EXsJprvyjIf+Igcas7A=
//pragma protect end_digest_block
//pragma protect end_protected
