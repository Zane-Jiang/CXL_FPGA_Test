// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
B2YKtwS4eyWnWuRXGQoCM/oIveVKGGCRMsbEg74S5LNQ4jJR18nr0jf5fN1Z
PFcNZ3d1eLVe2H9cze0IUAOlDTQckINDLE/SYIcWkKCveW1SzFlx4eDnk8X2
rS373PIzanzQfZgnwgbAxW3Zs3hA4E+jnQ5Upq9sq2coLR9I9HwmZgnoW5fX
eCVN4/VG4ksDNTerraPb6YSS+iGdV5MSV+E4YyoK3mZB65Dkr/Vj6IN01Emd
OxlhkUjc95fD/vVam28EDBfnaEg746bgsYorD1473XYpz0FS0ouJ+zYDwg3E
7lmRmFJfA8fsK/P62s+7FCX+P7ObWn1fkG0D6kojzA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YuX8TtrQuXyNgkjn1Dii8zg8SA5+xEYPuEiUeLXqkATsYy405g1La66jMWK6
4pQJqDPDSK0Frt9euzjuIOvOIHID90vqy0fTa4IzsXmDj3LlkUn5F86IW/0o
6WxJo5nChqDTg49NqsK2hFpvUWdqP4hV6KjLEVBSioNepPxoIXyGEzZJwJ6e
WURcxfZ3y+N2KALD2/UHtp9ujifFjHr+tMNLO+gX0xnJCTOgjUcgmjJgQ9jp
oJB2vX7IVKgYwsynkZZNvwnkIVciDeqhY9uTLa3RBlYkMN6mq0esgkWz4oCX
YyK9ZFi+BCKOgbJPWvqFcrDe8+JDiUP3rGZXKpl3Hw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CMbAaouQpcdeyd0bYwJpXmgvZnDhnhbNLH/kv43BZs5/0XYyhztgd3AZG0a2
d+KO8pNijFbV0Yqzc6NSx8aM/j2grp/NgVuVbjnR2aatffl3jSLsRK5AaSxw
BJ0/KSkrw2RfE08oMkN9qI+NfiTQ+tWvV3B7OUoZDMRlGYgt69AQM1D5CR77
Bi/OucAnmOaghr0BUsvh5dS+G9bXE6mocQUu+iaX3fyEZ2USRGum7iRYEGRn
xDZ/QOta6TRWzyBOfv2uYi3zhKoUlvUOs7TIJ+ram24zQxm+T1W7NnYMlaGF
dnzfySOBMvmUv6gG+CZzYkf39G2R/tU17mbZK4zbHw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J9HPuI541IOLWRxTF9iaToIve2SPOPIb1ypeMKeFZckm0hwRkLH1anVHdsdu
mv2rlPK6dH/mf1OkDWzXgztwrouDXGqu+CcoYNGQr8OFlmhPCp2qZJuVjzgL
eNnZBpGs0m+sgUXJ9im298Z8dytetBNn7NS6oqNXm+8FD9Pr2Cc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wiCS3IKboqw+GFRNLXs8a658SGo8Mgzcnyxj27M6N/N+r1QyC2uRioelVb9G
nfs1XRoIa2rQieKzB2FQFuLKGEcH8v4ADVTtkEo1/u9CeX69JjEcpGTkg8GO
Fn2dX4P74IwuO730Lj038Ym5jh36LYzGrEjlwN9JgTJwtaVzAWKOVtJPyPlQ
iMzV33qYmhsOspKSHYCF/2RQ15ZJCZXSt7Y9+pht+JAufzbh9PhdcKcsbImN
YncIagG7kvvGBNg7yNR6gF0jt5kN6FjzGPxITR041bYIHJksOoc4gGe7dr9/
dDdQG6Cf/Gsbnu4+LS8FF+pXYYSmxZPUEXxblM7HgNjTHPTAeZc9WJ3fwBuP
PooujOe/lW5+URlBu7ZsRuZXoJs89yFHSXvuYf+QSCfEpe+ufqk1iLNC+EHH
wVr4arxseCcSXBrAdXUmh52PoqeuxnK9EVXDufv1Tdb/QLIEao+Pqh1HR+H1
ehsIopEq79D2giKqVXg1g7alp9eutQR+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kF+xUlYMR0HTqpSP0z3CeGzHSDqrNglvNCeyEh5oOTtPPdLeSvKelzUj1btF
Li8NbmiDufaE34CAKVbbVkCEEWz2tEX6gSuGvCvgyP580d3VczOYORS8SH6W
AzOUsYIUYIqYmPbho8iulvK3zThkMb8sMoKuH/KoQqEN7AhguYM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rz4+CZKkcc6zwd4kORCrU/tiI8BWVE2BPJuyfGe3MtobM+ENozfWPJXYDTvp
pKfgoBP6nXtk0HcZFkBKr7o+hvLBPp8nDl7nxNCsoft1QwVZc8C1QArvnnK5
bxq8saJs5yL8iB+8xmNWjGK/i+3MIpV6btCndv218yW+Rl1o5Ac=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21792)
`pragma protect data_block
X1/TWvje/90UXXylli284kiEdZK7HWaVbhgHXKrsUgoGpIWAA2xWVC/x5IeY
kpuTAI1hphnwarOaPo+uOiOMjwzoJG8FoAm2S3G6Zd6V21aO1lCmbYcl3cNV
xoKzJhIQKps58208RGBf4Gbp6kKomQ+2usa2yXBrmlHlWfmIx5k/JeT1R0xA
hW4xcFnl531JaSlIHEskm2N4Fr3BF4/7BTY6NfEW4BIgEp0QnoIjm/TNWS8g
ocmkuICsi81f5xweWhsIoFJtZqvLL8LIwHu7wIa2puZ6Py+FS0+mT0WndXkC
C+7Shl218e0+B/VxyaF7qfI+ZRcEY4qO13RyAUXZrFXcrXYchjwubxwAFrCy
wVgwXqLVXh5ew0HMZ16zXnWIGM1mTVr+Jc6SDFaOMIMSFwmhqYsKJh/Pm83u
YwYiOccocW6A0WR4r5js2vImBdE028iXLekCOKzLzEHx1uMLwkepTB3EJrgv
cum2eBF3NtfcWBK8+70RD5UuAjLwB6gZIz9e6XARSFBTEy7BmK1dyAE/Spfs
Hlqmf1q3i2Y08f+k9n4Kj2SLFAI324nQRa6WMXfsmLqkDsEv+I6b7Oqhx4/v
/bRMgnR9bPKYNGw+XG5QNNKHGSRcTwgu619kLl3pIXXthGez5mGp/JOM4bbF
bSWvMygucII6Vcfo1UzjrOIE1NOakp93ZBheFs9pMNQZyF9JG1GTTH4bXiJ/
bclQMojles95VgAUDCUnXKWoke2x/KAeVL8Y5aWaVM8uI9ElJAuyR46pOiOW
8p+u9VRfLV5De19zHcoj7LdI77YQzOZ4bT3D7/Va220uFLDMZ7WVvpaM7AXZ
lHNinyOvwMlGP78J6UaIiYR20YiSet6kZ8dD+xQ9BhpCm9o9xFlHgG3TuUYw
eclFOxAZjVOoNsQZI5vKnzKibGaO3euEN8UfPslt5Z3srLZS77q843w1sF23
nXGmtPisCJzFVbDJR9bGDCBnKEdMFjiEHZDvRK36V+qiuv2r7C3iG8H/3ADM
dKURDVfM75MAPqN6n72Bd6WpZVkwZqKtKEEZDkLGafkO7a4+/Q5lQyaBB4k3
DN5XjyfDXp82BNr4TZo5I5jsxD8n+l6JtJcZpLQGDNNp9AJZv/7IYTiHXSNp
4ediHIwOJ54h7twJ44jZ/GctKxhRCSyawavvWrQtLXPK0P390pQDqi96sGKx
7cCJUMBMr3zOjRC/CVMWU4J8Y9jeYACHBniwRgKsv2W4fA5ylMXTmaQiqJjn
ywURYRkH6+wDSJojcevEavq1pqV17ho+R6uyXOHmGrtqsV7ENShsYgJ3btje
wFXPOHAvEHv3/nBowoEw4hKJcjvWvP+2OO3XDsfWFb6N5VHPSn/lNkp1Xwdn
ErgfoFPkJMLl/QZjd9zgv80pLLQ2ZN18s6AMC5KXOS8zSej5Cow3cA0seYPj
QTFFbAtJGbLRVBXrE8ycZo7ZTUQwHHh07SEKG1VZ8bFxFKreDNdltseg7G/S
69Ldvk9U/uheLs33/45plG6qppeB4k4/sEhuKealbEkpMozN1Nen6/0HfBld
zyh83+uW9qaGA2CMyjyBpZwgVxxHDVRnx2ffGRIt8akNWXxlF8y9/XbI/R66
1dFH5H4Qh6Xi94LxBIx+h6lPhGf+axXOTEJMfLvDD6586cCiPgfqKwE6gLfH
mUYzfOINicwbc49CMDyrKSbPez65iicvhCpvrL4RCAgw+si0GReqXluVOCzR
n2WkCN5cUxxeaHUTspUY7O4JVXf47X2IhqwAybKgvbbEn1Bk0aRJcN1c3nEy
rECA2k0bsEB33j/GrD3t7uK0+/zjPAUPNssu34Qr0CXGTUm62DChGSV1qwhh
NFujT/kSOA8wqC/aTBZcGWsUcEx05cysnUAS0Fsh3c4Ot4KlPC3mpM7JIEpW
74UmWlIhQCln/z0Ap70FjRbKI51W+IuyXuF5vYCREwROBk0fl3xdWUq4XM9p
x+52OQKpF10tt3vIIKjK65x3MODHNka1jyneWeD8r4Tt4SB1GxJct1oj7dk6
wy8Rj37+I2ay9dSoVoc1WmkwhkPmAylVMoi+vNv7ao91VrOP4W2PPFKA3cRp
UO01ANylGhwnDFgUPiNkA9DQBNwLND83DDrLsrISJUTEKW26OnLXRz9TrO6W
G/ulPUDtE1rsm/zG4wdocgkMCWlfpGYr53ZaSumqlnMGaXIGNyj7Zz1Trn3G
ygEPionm1zsmoXQKRUL8lLADk0IhHyNJRBAWV2oMf7Kyv1Ywo21Me3jyW5dW
KbOAGJYy90qBuNzaG5GtuJwbcl1O5Y4XGe9a3e+KrAItkZMCjzGhRlXCiIEC
CMprUT3EV9fuReAjmrzenk9Py3XqRtHP2oxHa9hx/HEjnM9Zyt5iCdCTKYSu
Uri2UbsKassFHvS9KjVEKziPjGYZa/JmT/SuwbcHWzCoCgtJ2anBzGAQLNKT
mgRITst38nmrtUlqG80kka9SQzI1J6QBXLX9qv5YKRRBKITgwwrGF43m6svk
2+3bWQO5hya7j67gBI6jSOxNvqf72/JIKcKxhIps2LKs66YvpUHNZDJezaTD
KeXqld9lYlU/V17/shHBzTue1muyRp1XCthRmr4BeNor60WPznyvz4jggTOH
0cfKH4Umt7hYOt7pt3sd7Pw2z2lS9kth6r8KgLC+9hrZ9FNuBglfrIR5MRqh
160iG9gMJ81O5O3RfQxG6QDpIAQ2AGnP7kx1UbcMAyudC4hK5dc0pkgGrGX1
/kMEuf0XM857jwBr4UxhVNvXVV68/hmD1AHADpRWFyDzcbOBwdANviziVuWp
zKVkaTQTiMXqbAw18wlofxqyZeEuYcomiQ3CsN7iSv5pia6yoIxyEVrpeY4N
h5OdTmZi7w0P5L4xyZUkEEcqRk1JOajrDCbnP2s8aZM/KOkWPTeGFX1k2p83
hRXCgaxbSGfyXYlsWiY0XJ8EZGMZAxYihBrI44E0bhdeXG4D0M64YZPxxzDZ
RedkzUTvmWDREPiVpsbtA+HAsEFOCODIIAqXVVdZc/AV68/dmhc83Bi2dQPL
1yVz1n9YkuENpx3v6m6vl6Z+5Kt4wcrpuKLGUqpTEcIpBIfYomXmAMh2vsr1
uJ6VSz5Wzj/oSB9yAcNF7Tyvg5rPtM34cO95ePFvmBGxVC1SlYQFS8xaBNtE
PlVrqKlpacNH+z4kiuZ9cmssgCCuOsWr8H3jQA8t7G9ZMKozhv9yKFmzmt6d
OBUsv56Bh3FZEd40nZjwo/GSqfWeyOUitHm1+b+Z4cfI0rX5kTFtHqKxIYgY
gZMDvxZklGNpd3Cf5GyNPbDFtfqmdL+F2G44c18O4Q8Xe11RihWLst15h48/
LN8FbXecEJROM524KmtaLXjAa3u7Aq6lnq6i8ZOfsQROC0b1j1RzazzuE5dM
F9JHsqf4pylHPtM68F7mYyeCFf6x3Dj5b85fTZVV6yQtIKjbJivhBO3BSMBn
oiYJJv1JB1CYT7LJ3GcU4JFcY3bWEgvpH8m/GvzaUNe33pYf5eKILNaWS9GY
YXnyfqVvbJhdA/Axp4sv58Ypr+cywDNO8tjK9W9vSk8uW0g3ofOdULUEROzv
gdRGmhVwjJvlUzUNJ8kULlNhoQft8ltX5VcdalOJTH2AijalNz95Sj8/Fq4s
ZVrCGIIOU6zFSF6eaw+i8/4nKpv6q7vFYUZsnO+bYJo4gpdXIoZMupOzeuuH
jFVBOw/0oaX1dwaE0C/d+54OjxMs7b0/qJ0gn89qJkZjuGOMdMInfQtpl/Os
wjtQ94fD/uPBJCGgPEwPDxAj5Jg1n1VfJBoyvz3BedAaAPP+7pk2Idetef4m
3PkJsB3sN8tyR/M1rArJqWX986zHd4oBSAMDuJsG1sSF3M8MiVCe1Oxku1fo
igMYGnhrEQ5oNZDqZ26k2kiUCqUBUhj4BdqS0O6jI6O4iz61o8oGngIMou6G
8xBeEDBNh/Aj5hjSAHVjUMQvXY68m0ENB09vjxRmgO7lLEXxGUkB0BmH2sKH
Tea4FKDgbEQyBtlxOHTYuss1DFXTtkqR3EDrHtl4tGO3LnxGfXMbugwaowhI
8uEBQUb5sij0mvuXvJcuXhI17PGrRLlztcrczv8j2xJuhkHdSDh/TtzMhENZ
MPflrzklpfqWzePWlltzSIhTE2vzxvFCBegSV7AYnndHqloo8q5g31mse0w2
t6faoXaVvd8QdOh/PNfc7qwaKF8i5T516j4YN75NDaR30OZU6pHlQniqjJOZ
vg5COwv9ecPve+AJQXl/3TjtLgCs61K+LV8L1I43fpIfBSkaaoyP0/s4yLzs
ON+/CZqH+m0yDt+UENDs5K0+1EReVhFfkhUNYl8Wk3LOla7VSsic/w1WsIlb
35mzK/jPTZEIx9vK194maxelxi4XHq3mv36UHTK7H14bZwukIITz+a+zRtQC
VSAy3ENC2vA8wYYt3FEetFj68w88xRKoSe3uDO2gpXNfdkr2O1+wwy4A7agI
6u7AgejkTiF6ijzbEUb5aV/siB57xrZzkZ3DRSbFI+lpbT3qdsOr7RyajFkn
dSIn/d7xtTkP17FVDHicr5heFS0xWOgvhthLxxD9I1XmQ6vUEEOAW3YKzxTh
o38Pi3xaci8+YhF4c60oeroHG93A6aNbAoKmjpudj6HL5StIuGHdrnb6jCgx
J+qJJVHHUl/iSfGn2rRBLyk6u7NZA/gb93pwBcaD4nI0uKIGpPvPsw0rrIbq
evxW4cuhtXLqqzrad1zhPZ8Smp1176x/lVeFdCXs6+VOL+MZewGnYiO4tmHz
vGJJV1juBvMXCRTct7y78uOLIa57Rl8Lbne0KlFMInvo0K+XDVz6/CHjnv0y
9AXmurGKzdUaCoU9vn6Qh5EnI/5BydpLd4PgZhS+ujmqcDdn43H+/eorjIm5
R77dbiiLeKZ253iBe7fPy0JZN4EwGWDWs+thHQQ4eo4Dw3gapDyfjDeapWL9
rww1P8CnyNcsjVm6YBXfNWWvNvo5eg7Rqg6KRi+0J0yORVN4pU0/1XhbWQ9V
bouRhS0LSuuORek0AYRveGaXHahm1I8pnTeiIYc9UxifyfoWDTchMtRImSAr
isKNKB0EMizy/ugy8OaD0BQ1vAAE12nbqpfZj5ry6C6y14kZyamzun5ctbWj
uXQzkS/PIHmx5UyZ3YoQKpYcwovlEVv2cnwoojxnvWx/fISowozOfUHml0cW
kNb3Yzl78NXhTl+tOzKsruLrAOSXu9T3Eozw7EnOuHHf33njptVhsIL2jQVy
YnZZzSP87smUaoRvgCpEPtndbsTvXyZ6gvB/d46dqt8zEYOU6CBY51O0gta/
Eb+FfG04NzUU4IOuWMSp3tozoYdh8HGA2pkjprI2OObA6JocMfgd+lSlikoU
YizAna4oAsj6BqB4G1XHuiFdABgdHdbVcic1J0DtUSRxeg01Plw+Y+zzal/u
Q1aSIo0QtrEt7+K4RSW3j7d1yWJzDKL+XPzffceVFZWkgNsuWZfdB17Vx0Y1
npoN3L8WOLYpMSwt/3ISOpHIdhgiU6VrGeWufz0e4JNPvOb4iTpTcdHFXCAd
0iPGGbhN72dRa2aKOSBEHwCY9kLdF1C1W6QwUwGow1V169W4H7goIQzq+0dK
/XayCADMi+9huNeqmeX64zwUHs7yGnvuXV8/vM5si/w9A9UPFXd0IYjJgG9P
K2BTrt+HQ/NQG+2t+ZvoZCESfNXe7wkHeZu8FS3E4Qe2GitWCzVuHCG/DeIk
qOf8D0qxT7D8cv5xtirNQzF2NL4ZUumylS1NeRqz2HUFACIuMTA0btJXr41K
BdnrXI7ITbJNNR5HMUg3OEAvoOocUFH934nQjeTSEOpa8nZXPrQZA2Tdwoj/
eXDulmpj9B4T1e5dmaQNPWGfrNwLFZL9uAroYYa5IWNps35VlM9q0ByW13I4
PpJTtr39rjs/VmHDLYBZlIdrj2RKLBD83AuYmlPYIyS5UEs4aHnUdkSqXu/l
LmSUfCYWw02nP0tRglBcL/8QM732XBpLJvtBfn7fLyFG8ceaaFwOgePMo4xO
HsMrDp3D/CeDa1SBln4h6VQXLLBuMRPMV0B75/i9Vb2IHJWYwEnfJtxH2pHN
pdp+byPSbxFglXdeknEpNlWgYn90uBXZ/FRsAeuE29Ur5B+x3oe4JFOTudVW
+9ahrQyCb36zNMvs/FwmxV+3zhL5EElW+ZXa8VGaxPX7O3ibGCY2BQQpWR+u
ojRJ1UPoBmv5oAocLb6WwAIsfW1SSf3+YapEY4jQJoDOuM0kjidWujM/uURj
vRsGFSq8r4v+YV4ap5s3j6n7DxTY914ZxCimkyzVasuO6VvCwZQFZ5Df8uoZ
wdPkFKvA9O5xYX72GPykN8U1fSJJ2leYLZbPw1Z7XTtJNcY5DOXBGAqZOIVv
SJETArBkB323cpmn4aJ5v7esDAXuDfZw6dsR2LJbJemhO3ABfPH+5EsAVZpr
cAHp0QEPxpDWJNM03HEzFjIE2/nnfdBWCzBJME62eeP1e5rOSJcQfakoTsI1
SMc847khijOWf2bQSP6fCHCiBiF0tnqW/lknhXAQcevGO4HccoB4J6+a3R+B
IFzrPZ3WemIOlYXIOG9YsTZhmSypVShUxFlOM2cb4t+xwsBKE7i9bDWVv8g+
Kvapn2OPpz7uJRSoyR1IHuNI3lCS4wxzVmy8Fad/2Vh8qrniMQHkT1byCs52
aJK/1gTZiX5x2FbIrtqJW6vZu2FAx1NcX3xxTEQwzcLiIooS8ANFOAaVrVTy
xkkK/FA4Aw8Anpw+KweUmkSn0PVJJSLjmEQS/1PXPaB1KEFyxdLCsKqkyRmw
w4WyEj+2W6uYDg23YzvH8/WyanJTmAOYmnVjag85mbHzYE0DjdNNZJIFipb4
K/WRDdfiEVjDJQGNylbV4rzYTpDaPvXpC1wm870SwiFOVCF+oEJhgi5FcYxz
q3UIUlCZToF0pDPAAD72QbKzmzaH813ypKOAQau7TClcFRt07J3Wt3C3kPtA
YL4REWnXpz8j/qJTv+ISyz+vHc8OY8F0yQd3T0+fhCKKREyLt+srYhM6ANRM
SyvXgW/9nGn+Jb4240kSJa5tDcz28zFu+S4JojhqRKV1LIzk8JLs4H6dfj9P
ES9p2vPGiASM45vdkwRyw2fDsZPgOFiDtvClEQn7k/8ouraqb2E+T84JHCMz
JaqsM3zJ6VwMom107uaGR342BbN5IvJrgFeRlicO+ZC3uxgsQ+oBq+ETfu3w
3lLMqwWdIpc5AcSjBIgkAGjSyobJXL1iYvgA3rV7WyHv1bG1Q7HCKlvTpFqx
9E5OLrJF0xbUaFhoI+IYRBeUPVcsMiZf8AwXCCszWzofRmAlJABMdWKqeRbM
zBC44zMKX9NQCF6E82Wurz1CoHP5xlz4QOrupS6GBKQDioZkogxZXzshhmPQ
uKn7WuzhJd96xGvfuisPs/g21CesI9UVe7EXVmc4ssKTYMOevPO9LjlreDS/
iyUqIjFq82+6YwlCRftC4mDXYmdvV3S85LnRl1xG3ePuJGTRwl7qdTG6WWG0
WugYfD0U2hkEDVcWgBvbDq60pmj4zV+I7LaX1UMLNLEg/OZieQabIS8zBDx/
MsM0YWvBugqVzahfQ7BJkCgay0ZZlTsIUu0jBPKdcD1VuavpelTrUdBURL4M
Szr445h4yAzQx3vhHIXT8k36irCOm5XT4Ia8ntESEewwVFo1NOCP5xrEhePe
oAI+dJWAaEP04pyKBoauZs+i/nMy7zbEyB9LmGfg0Ru9UfsmDPIAqZC/lbPm
BQxdsFA5nfiMn/8vsa2RImRupfLN2gPizUbVa05/k8FVENWWE4lPEYhtd8ME
ePgF+JYveeoX+XSosCNGUtym/18MIZ1K/I9cIEvvYImWwGtYuh5DPxjnQBEB
d+fQMGLymPTmZ7NDVN4PSZqw7uQMks8fbvJODFOJGk5Esx9C83/9Oo+nrPgn
OZLYmyCOe7Ebs4gWrkwuakhL9BQG0qXH8cKhw9zOd7sbM+n0/a6xketxn+99
0IFpzRGK4RNktKNXazhKxw4f3bYUeuBy5T72PNN4x4l4daJVvFZ7ZMTyBa4I
E5eUG3eUUPB/SV0W58tRGBiRwBqVA5hJ2ZiTWbVnhmX/kiV6AQpdCXhFWJzD
Jg2oOeUNAHBxvdw1b2HPK1dgmRMGsb6PqJWBbh0+Kr4rbEzABGuojSNa0ja3
jZxWi51d7WTKOYosSAIKZ42+asnl1OX4w1J6f5e/pUe1ITS6CUuhjbN+8Xjq
S+vxfzrhy6kEZZzrLWlAaPfLlxhKhHMd/hN9Rd5WrCEFzuBa+LpkPtAzUdkt
oXRw6+/MFElP3Pop2edcRUsEGmUMVFPjA3z2ZgsMHyYoAe9s4Y8qz7a5yhdZ
uhSq6tWl2BNTU9mF00MYbEg8keeOYa0cDJeOjnMlyBxhSfwiVgJiO5CKMIei
ylv6qaJcjKbU2FWI+rGHd1J8KdZzxLRSJJfp5d41rk+zxwZxsyIi42feNRVS
wk+XsE6sN7Xk5kAqKJSkEcM8zxBaA9vTIqDzJTPIL0QL/TD4YNibvenJdP5N
2bVn1H9SUUV2+MSKG3EPOQRR5IH3L3ugcjjnEcGuqrSCdF2ykHp4cMe91eOd
CR0ubrBew9e8Rc7zx0C4QIn8iiC11IcS3r9/VuBRDsuCAJyUIdIPcmnXjals
EfuvYvevUvfoa9XHhWDHQR5BR4PetSEruHVG6xGKe+xwebcK7p4G1r3TETEK
3F9M4Z2k0amzy3IczA61CWsxz9yMjFK+DMoxYw1yckzJb/1J9iiSqevxKHmU
/ucxPw7E7CGcfFSkeFcWicsGlO7d0AQ9mH8jC9LGF1IwhXr57eLXwXUhjPna
QqIypxiE+/kneNklSWHbtIHZE1lF7HBco+/sC2kraP+9dXbzAr4bEq3+Osu0
cR4W9sWQT+zdjLsl4zTIcYDNW22vdfaiAnnbT1xL45fgdWKewCJDzJVQHuWG
0QtGc7gbRQJv0jdstiAbjng3yj0YFEJHPaA2hR4EbgZJpc4ULlGSx7iRpEBc
Or2N02F8g/i8DqeOePMeJTgP4+KwBL8fIGq/yT1AZWxSbS1nEZbkH5d+kOUU
aCYEq2LNwj1LBM7+AnxHOsiiMWmRcVoDKaOZPSgbWpij/FMkmsfxhUGAR+HQ
onbXv7MHCW+JMRrQMv+njJFp5riESXeIxbqftYHp2tmX9emReK5oxzgm5FPA
KmNQDqtjr/K188CrQ/zq4el0LNetjg5VZ52Ijuk1yQPDNYuTTkFPjvYW9MNc
axkAZgRHxdyH4iRSqFTn7t9kDsHpmQWrqyu/3Cg6fysgCcUHfPbQIrqeD/JX
/KeTEI3BA1cB9pt/xyp8bzJ8VrCaIsUQ9ZwUuF4m+kBPjk2r/6AAkx7IWHjS
ClYlbNnNR33lMLPwcs5inMUDgh6EDppnZhtRfTg084u5CPLOXenXvTklKRxs
qBozCcP0pjEmVSLSFJUbZlzL3pfA1+jmWkDm1hEBlgQjotHrped4cGDoWyMs
OlM97THsIjhLsZV1wbwTdhy/znPmctBNEPaown9UPazv4uzgeel8DfuV26ad
HFJqNiQlq+DXEqKxvhEAzNzRiX+oV0d9tKE5oVZTiBEdReReDGWn9hBl8kFC
we+bYE5UwW6Gc0TZDTdEk+SE2DIZRmW/VC4+YkqulZg/5k5ks6TlmKJsaNR3
29z98r0xjk+9pwz+Vej8J7caf+Z2qtr8RgNhMMbK7tJYoGykT+nVssxffd/Y
O+fVOMdX0tDDFZZmAA+hmo958KI+qh2rhr8p/30oeheHsHkoR3wi3CWAnXTx
Axql1iSDT3OXe39saYxRBkX9rzBitU97cGqZg8V2JewkZ+DAr4BF1RKt59ee
FEdGp7/GlpvGNxMlYLUpSKUiRO96UzgZNCGY1pjJtNeRSAIZHGzD2RkZi585
kwZkG1kBeMHxgzcq3O6hcJtNMYj0zzxWO/bRgpDlAc8FV7Mb6mr4J4YrD8UE
gOaFRpYw8Nm+8qYorf/i2TXlzid2DSnM8pCSiDUFaS0x9ml2GwSzBSuNLpDn
07Sz64t/gMEKuwVINFZ44+lwvSsQnMTt/nBUSZYWcqvu78Fa9ftXKADi3ugs
9yxNQBcdvS9MGPvdmxk19OlaLJ5Gh/w4WiIGp/ylaYKhKt7oKzwTCZFb5/Wd
/g7Vs1F9flvEvcsYo9/hEugRfg/mfiWYWZs1GB5cR73CDjktXIi0UDhVRqIB
fLS5ew9OJF4pFjl0dbYuPUYWBgXH3LuNHLhF/dir3imd+ZM/7m60AdkbFxyv
8O6R9IN5tDCC6TuHBrFAGvSElsSWj81oOG7ScRYljPrzBqejly74MvuFYELB
dDEDTjo+wzYWa46iW5VTh82+6wlGuHlBBMTUm28P89KXZb47B8GwBn6gmg8P
btKZp9FMHTMamgkdIOzAv2gdCKR6fWwwAxBl/1HiqohBmb5ODkyM1Ko9p91g
7VNkOLV3gLATiTg8d1A2qxCu/wfTTLCW37AGjGPwpxXEvDtGN9VD3zrf1tv1
aZAXIox3VDAh6Tq8NidunLcax/sohMiw0vwsn6qwjgxKXNzzDKYfGvq87wi2
0rJzcZbTqyVIbDJ2owe1KtQJeeu6OLc//Z4qjx3rnViY/uzG/20U2PfoC0lA
eWMq+l9oFVC752+Rop3pStaPsa19tzybGa/e7Mrt2C0RovWeCu9MPDpH2Ahm
chU/kb3ZTf/aktktqDYYv07bhDD6Zn3TPvvH5CUHFItlC7kT9AItVfOkzmKg
du8lOZW4HqlX/0PzSKtqqy4PbWmpSTvHvm/bbCSKCj6Oa4mgkor9bl1AFec8
IExwq23A+0OHAoqvava5zTILoj7X6oGgJthDr0s52RwPvuoqHwtXc69GYNZ8
+shiVBVcZ34KUq0JWP9FXfUdFrqVyD4QmNU2jcyx0Bp3VGEzalZVi5T5M036
EWfNFQF+qXGv+HC1995QwclHnVbHDSARVv9HTaQB9npj5dR/cBeqUSaJulTD
jVhdy3zG9iN0oZwzSo8B9JpEKgrn8NHDGWZVl/W17ikcjF/q1kQ2mE2ZKUEU
BDmo9jmOlCdIh++/2zU3Cq/iEX3oiXIhXF0tFSWfOkrA3B5kGp9EmedIY7BM
GgGm7q70tkMkpU2XRt7dgp5a94t6CqhYLxVS04nBurlrb+zN0JbuaPSFO1hs
l+xaRevInMBhKibCTaN2kEM2dxLbSaRL+LuzvMBakFqxR2tDp7rCAgudu0kp
78Xd+F74TZ1Tq8jeOnmA6OkQeM2RiXqo7RslZzb8yU2Vjtqf8/3pEZsiF1u+
CsHxXNP5csGD5qILOu6pCgg+zoc+adtPtAOH/9cImc37gIbka6IVM43F99y4
Q2/mLp/xd5BJNfds54nllD76ax5GXG2hqGCqRrZ4UCUGAz9kVu5ZEHrrJx3b
BU48pLasRAobCrSpD3kAMMvMYtsE0lL/UtzPT2J1oFcRqXPXxYIQsBHD+zye
MWgtzM09Z1fiEwcLl/HH/govvO5SPJlDjS9xtO9HtESofWnI5+mYOfD7TflY
SLblW7cGXMIftByeoJ9fd5HzcLS7DLmEqKe5eUBGiJKQudNG03kPZiWscrQk
sVPlMiFDmGVWbBGzFeEouYh7CyF0IdsEIOOyvD23BGt7zwnrhX3WYiSqvBLL
bAAc5ORzd/mMTw73BKQKZrWVnOwhQXpEo8NPqz8n9o54fWinqJDGMo+BDvZ8
e3T8O1VIdPKfL8vAIpGo7DhirCWTOZEEk6Sb1RO8bFaye16PZQqVV7hfNzoP
OvkTFKoLK1CmXlAsTXV+jYI0VtzZYdo6i8uUS8AjxlGi7/BfvXL2CSxT1MN+
qLBR3Aw7BpVYgL6jP3iiF6FpOS6juXzqh/iOPqFe9b+WBK6bXIwqg7knSa5b
PDVE1L6hHsDgDDiHDJ+XsoXPglI2rFG+64Jq7HkL8Mg0V+Q6l6PtPKX4goFG
0dyi5BUPaZgRJc0pORbh285TqPVk7b1vuaBFEcEFPvVwR9Juxoies0o80wLq
VWgcL+rekRj7HYnnindOmD8dbEjdfL1jbwLdTAvZNEOsnBvszU1qcCKgFwxF
4npQMvYgklLKONy+hDWgwm5XosllW3RccgDhFSuRWNYQSA/8j1HoXdhwhp7Z
ikgow5GPSZI7hJszg5FIHUI1+wePhxKkbt8AV7LJ0+aWaFqRE4mfRS8+zDyN
GqEMebmESv/w96PMEKs7EEHlchVJmurBt4sm85pgyyEa/HrqEfUb25YVqnyL
7/WZFwWt6GVxtI+AsL+HSuMzpB0tB4C6OrTdcPZgRIJtlpHZsWgfut0lTxfy
wN1iw4GVmG5bsKK8mUjw3cY12diiquM5Zp5C1dhgTYCwYYpttgIBKX8SaEUo
CNbd6k0alneP01fxqNQEPFk0SM/52lXpRPBZDFM7uEaiwGoe8b9IfUBurj8O
V+a6lrEcvvN8YkocY6HD05kEVij2wy0KJ0Tq/zuACynHm7YOLuJwobRk/Dlf
f/8gXBZ/QiAVlhcFpOJ59TKSxKne9XHA0/HdhBkeEwYicHB7WX0ghFAJp9VD
ZaB9K6J3qj+gghVjsQ/etlOl6GFwi19lrAiJrTLPcSgVpkn/S9KUx4zhnV+p
CGpg8ojxNgIE4OgrlLw0LK6XNGIlrW/9XffHgiwodVIsw5+26jisJKDjxRgk
VqwethD0LJA/UKc8kBtagczi42SV5SJtlfOiUNBERpmLcbDe9j2eNI621rLk
Kz5v2Xy2k5a8FylZyqSeqK9j4fEgi2w2MufkjQ7z+J6tRwf+uQrWPYDs44mm
3oeDMcGuDSQ9Y8wfDW49lwjV8gNMqyw6CY8hL1C8yuhqRUKXLgm3YT2aWMlT
PH7qY/6IpvgS5Kb7QTGgXTi1Z8gVCgvR7H1wfvN+LIzmxhT2OzM6iZIOjZqb
OMq4XVtAVMi452Tt2xzF4gxI3V6LWOzJoOWw3NP39dxKy3mHRitSGoeJnrhv
Omwp7rPMZ303lspW9XJavx5LdaIAlk1Mz48XTZ/YW8IiNVrA9BzOJkH7CvB9
zqlN/ueWj2xWRDBcXh4UKqc8y89068A6CnOoO7jkDUaimu2bFFBZcpN5Ieka
FxAkgUc/ObkdOsq/JVuGjMuRx01NPTgHHrs/FTE8U0aAHeO2blktnhyWjdNV
XlZnMGgyPXGsCk/ZohBJesK8FA7zLyiDkhaprQo0yZB5HtYNIk+ow/4ShVJU
1uMAm53ihEIoyB4l2MPtNSWpzFwUlJuoM+HD1AXoA+bXPHxJxZ3I6kEd+4um
9TccibnlaMf7QrQAJsDWnswrZuNnDErosIT4Mk3GuzRS2h0slyuOdRmy85lT
4p/A/ZbKrH5wI6eIF1W4MEM5++U5cnufyvFlTe7qpX9fF/U30NVuaWbCfGQQ
1udvw/ryrpLBBO0n31bwT+qcDIDL7LKa6pzFhVDnvP/xCZrr2xNvfJSq3v9j
1qbWXqeu+DF3oXrtwsSRLq9MYfS3x2ybC4ViA+15dZwo9jUQRyc6b7ydNiBq
vFX/z+B1WyawYIOh9S7s9RjUk4E1PDDXb7sDIhyLKnqX+odXX7W5DN/qZykq
KEISYxzfVxjVyUujpfHHCJtyk5w8JMnH0KeYXQUjukDhgv9sUIbKwK24PziP
B3ShSbCIMCmZY2PexXquFNpngdmHuMF/kkeyM6ZPZ3z6p8Mb741wKH9shMme
3UHF8OXvTTkU9VGC/6Cm4OiXM2yfGQhiuw6VNJAX7CyUKnPbqtuXpGx52UEq
oC23A9OHFG0415XSsEt2KJEK4YowFN/HhkLCy63w2DgGLUGav6dQ98GbVcg4
OUvdPz6BZYTWObIM45GTRlz16rBC+NmmtrAC+LYr093T5yW35xmLyrGtfabW
I2+VHHFNkiWkd6g7M2Kyd3FYgopal/nyf8fh+ij0IMp7bqimCxFpD4kCc6lz
x/qIBCq4q6GNvvGYC4GKpqPUMpzktA0T1wCRE3yvB6Rf5a0iPru2ydpS6UC1
5OQzViUcVgz78xiMu6R38Za1jQWxU6qJIPOFgci59KokORnaVBoVw+uJJN5c
bqKMVTpYpkJmTKfNdgB8nQmIdpn1TWok+H/QEfAqMtdGntf2iKE0hnkwe5WV
O/A3telOPhFgOYhZxqXUfsrc3UT6hMF1YlxKDpQz7ZipnEJeIub25/DSVzD7
VyYGAliTCf0uMPHXgSLtd0QLHx3oCdkBh7IP/b1ZbJuVPXqSBsA+82TCeTQC
UGraBgKDcbOF2mzrhiaZhbf94EO9payGsc2/tqPJVzXYDKFgLhiCIUow07Qn
thzpZu0zVmanRPQbp1+gTHIOC/cp6xB00jEtoV4SUvaiIcSFwapAexJM0vnp
aYpZ/GqyRkgZSmGAMw+1KswaRbURkZAfPjcnY/A8yR3SZDXu567K+/yIqg65
qNt+x54luVDvesj2Ug3F6Yslo8iQL6i+UilJJ+XvowZ2rtvmoiwLD0igoc9z
AL55jBJLKupliUuml6HydRd3OxuFtVJrIpRxe0twqO67cKuKmVrgRshUxIJ+
ObCqOBgyUt3h0Z3z+0y+GyuE8HJsaguI1uGmUJkIPipDh/RI2cWyTgG3AV8l
CyxY0U8FUg7eSV0cKSPSgw2ZyqaRREEWkbhS1IZ5E0cxSPdq37Jy59HSP83a
ZYilHTFKy3DDyT1/3EtYuxMSyC6spNKWC4d7kEu+/lq8d5Eajgcae/kkxOUh
FdiGG6ASqCZ+vsHACKog3A6gu3M285ksqvS245bY00l9leDrBcOD/7uey2a/
wOde2pBW3lHPCPWB4ih1pA1nW3/sp6JOuRoTqCyT6j+dp7HPL7J138Q//RAW
2FZzDT09khrJBSsyPu5gSMi9R1FJpf8CyEWaR1VHRCHYebbjcoPj1AImDUEY
h6xjEd6Dkz5N9K+ovVTPhqWQlihLILoOtfPAqco3ubAuMk7dU1HpT594Lla2
moUW0X3wmbyY2yGVmcZiYtENPMNxer2dslAEthbyZ7grmv3bDGvybwgRNfIf
xp5SwjZkGjxSFcrlLSv+1/RWk26cndtR13CSOKkIz0/SS0UTpOPi6SHM6UFl
hzXIb82wYNdV1YeVRr6C8O4cBDP4DLhkhFnxJQ2RvHQxSXgp/aAaLctlSvaG
oDRvcanrO5wWbKzNDcwyUIdSBihTIhf36ywSmo8GbriGnJQzjtRj5HnmY08E
QwFhNA5Psa2KcmUQabxG8qlDpyue+eeGszRqbgXzAv3H91cuAJWgwMLoN+Bd
+9xjGxBL2+jLg8jrzCeUL++KJVLYc6XtBW1v2cMyN7YRmwuvm9R7G5LoH20e
w9ZJ3qR5AnqHPJFyCmEqqHtWY/EEqu5wU1u/7PHkY5RqLNBb+sWNLJtRhiU7
PETdJ2r6Jxw5JjT27ulOLB7NHbkCMhqAfuK4HuhmWthKW9vw3UMEbPIf4+pN
e4D+QtP+0Laj8BcZs0u4iOi6ePyUMecEDfwtfXgFmHp4MJH2TwHNa+V4U3PU
gt46n/MgXNLNCvHS9MUoNAhToyBj9f3qnkaubHel5uC9o+zjRI0Ot7AkdEOl
8Eis0867g3tTnOF7SJAZ8Xm92Ap27iKJgGmPpFwNIPT1GWjPo1ta3kK+IeKV
TWnzWwdXVp53eY2XDwKWguD907pw4SoR229lXYnog70cvuZZU2eU0kQ/BUFX
T+3WZ3qmfFaR3oLFLlfk04udrzvY+TiYjLHm8TYfgjx7SWAXsQxpvZl2ct2V
FOhOd/0HSShq6mt0ukQ2z4OwlW+5QmDdQuguBr24sJE/vj8JjNY9XKfLsnxj
H+eEu8ZTDj4wPO6lZk0fIoNSRapkbRyEgbhkTeEWLuLTjw+HyZnhX1pHD5es
zQYI44OsSKzl+UquSLW86b/VZQ1qtSBoALNA5Ty3n8DFgs04OFdSWS5ayJJV
ev2eAZmMygjJ9Jba9nQPle9FDupj6fYk8Q6zHQiOf8vTOEOCOlf1P78vmOsI
7iPxUfTfMd1gjD4TKaAXsDsVlQFsrw4OArm4Ya3waxYqbnFEjYdJ6jAcbT+n
dP6T8Rmb+gLdhdhANsUQevxR+EgDbXS+oQ/Dd1l333/ejU7npH9W7SCyF2B4
CKgMjeGbSNQoehSJtZ7vtrpn/X1u4mHI+8fYOq0lcm0GYQxA4U6gLyxYGOp1
zgD1CzvpQdxsIwS3SBNyrv/TlspC3eCNt5vvYPzj4bT9hYBPlcrE17/AjRBS
2fApBHud7Ad5pJWJD8IlAvuuam9qt1rS/J01nxel14halTELQyAhYp930hC4
5DMZSh1UhL3cmFg4do66GdLrDyOjrlG6AFCKUEFcq/0OHUxMgc7vURMSPS+n
vUaTS7aHoOZFux2RNxDbtbgdlLaDr8BanLtH4XK4ounmh6EiZX6MWY0czXrf
Sa6EH8UDcmhVhccl7j5tsBHI/IvQ9IkpAmkTy+V9vmM9vHSWCyf/umPvBSgF
NhWSk+mr7HrpbmL6kVrKH9hA9ho8LDST8tmbiFt68mgOBSHOgvrtujb0kkvy
HjQZLRZzYJZ5JfmGiQQXPGK/9tLPlTQydxq1fY+10frMzpSPF9of2LZo13Yw
PfaOKpXrcTB9eiRc2dT3cXs+5dEi+Jd/VmrbRxWfrWLaXYwPOicHoJa099LV
J6c4G4vlr5M2tU8I9F6t0mnLJyGNb7OxAK9wZjs9sCnUjTO3294hRALDV8s8
LiAANZTqVdJIYfvhZQXIh3WotgkggcDuqdYEoE7AAyAsWJtFF/Ann5qcPZN1
ireTjLZllpyoLsa+VbP/JLBr4h6sHLISZVcsaDbf/OU5o/8CcyqPe0V3LdXo
c1y5hw0KOaN39JHGjaMr3In67gTCaeBmDK4W5kKb3ycbnD9S50zbKnXG9FxO
VaQjcEZ13Jx/yxyj3h5VtmPlyRodQp2CSqUL7dom7Q1QgML4sVOyQCvVStKk
Ah+qNhFQeVBfXomomcrejTXeW497akPcKi6vO7vir2qHRgfa+i/MW/N9Ujzf
9t8zP7mHhD3r180jZgpwS6OIXWCSRoFlloFAQer7rVvvlYWzhmcC5yiHiHuN
IOYPYzcgyxQW8V12oraZPafeV1NhL3S6NY02CMIGFtYr7EORCYI+/DfcJgiA
Idh7Xa1/hK4IS2guDgYAUh+7uqh5WJgFEHXA2x7C+FJ3qdidEYuZrk+31XrK
QV6JIVpcj5P3pnolwSdDjl01gsdCiWFbu7Ws2B8khISQEz3STdt/VD8Jvp1J
miHfQCd8j3yDPgDmr4QqKEu4kGzo9a0OrNX/ROCR42q0dfU1c5CgTQbxUILG
MgBuriy9GDZ2QZbMNp4kmNIsKyuRqCh9q+AkzOsIaEhY9ie9/8uT0VrUqpFC
w1jqpRCxS5QSDycseobHtJxhqChSIr82mBFRGsPQMrUexrfwGqHDyY/mBvtv
Ax4H9UJu0WsWdKuzPpSpzbj9pjqC6dVKA9mVm58pbbSYRGbGRJTzpHyfE1q7
8pzC63e7mcVhxkTUjlOSiEBtFXYufhPUB6wvLE6cgvnHwlYY2LyXNhz2dghb
0b8g8PTYclXP+WdojeW0nERNlbDZpk04j2Ri409PAGnLpaDiujSbsWpI7zoc
hAWe6VjOymRkAXY1not3/VRCQYCWOJwp5QMVHcReVRIRrPhe72AfMJKismHW
l63yPcakON87ktQz+yOEPu/8sWJNxWvDSXtd3DQfm/bdgdkLBOegRxdssE91
EtaDDzl4dOw110rJJTUV1bhPtooA9GXUjPog1UI6RZ906YgkZqoOJyhoyDBV
Z01zi61MyIkW2nkv/hgFFfAqqWsXv5UGoPdqE852PIPlrcNYgXMF+Jx/W9e7
YxmAwGzxonMziydoj30qIwIXfMY/bR59nKe240EoAVC+9vAbxxjn7kPyqP0x
a8Pyhjnd9SYp17yj7lY7N2SbHpiqtZm8mALF5E0W6nITEQh2JG2rk0XNYhju
hIejiQOyBeLaulWpeex4oOCd0Qzxt9cfa+gMoXcE/wecqomPFIPRbhAizjsA
YwrO7QrrfW5HD9ChRB04yqVM29yqW4AA+9h3boqzcSGtHwboHEvz/sGMblgk
araYNpitRwgTeeBNFJ6bnuhu8LqTDo50bjC/t69zry+0Mu5Q90qeljYPKO6K
n+YGIxvF3s2hQnA61qxnlFE+u/BXHnIUdyP5W7v8wrFzXt2sxtgdxGmyylci
ZeRRHk3NmGQ5MyxejOKnlt4d4+clVHaF7BTG8rgQuD6+9cXT24sqAM1vGZdW
ZnQAfl4miPagzGh62rO18iNyIc9/6bzHPcly27NsP0glStItyLPJ3UAxNMZ4
4SeBsvRtBltAn2I/BwWQGNY/R9S5WPkNacRKV0fM2FoHVRbqYQLjSqboC75w
BEoWuwDv1VmPuiXg9r+BusITCJ1bm2/RW+la+KhyN4da3ggeYj7P7jbC25GR
qdb1bb3HBP00tA3i3Q2dQzQmhtIvv8JSzvxXfX9wKwC+QbYxH0DLb2Rbu4pO
os8PqB1Axu18xyYVBVdTd9k56AL6Beg7tDg39wmjGLsmhX+MqTBuSKDlHt01
BDWZr2ZQbdcNZslq9Lmwhx+2ZFYsHokpSbgf1LcLqMGbvS0ZrpMtCSEPvFIy
DU7npLvJrzGeG48EYaZRysHrZHX5VhKe0jfseiyTx2apR+SsfuhPbbXGniV7
zJkjchj+KRZs0YmvY40grsLO0Cd2iq0lRWhhb8d3MQFJOfF9zguB6voDjFa6
tNEqKYAoja9lieqT5OarK3FLYZmMAyDOn/vyyAzO0iUVgmyNgVdigYYyxJIg
s55W8ej3xciQjNNvlvoT9krzsB/6ZsNa0jgK614hi/mFGVTfb2F1IbZIANJ/
P1BtOoAEPSnHQK2sc6V7gM3kIQ6Rt6bPHcuuqkjjvthPuyoTWJ4x0GRzjB+e
2ZOPssje2rI49wgS0qkswNBIcCLwSv6mi/BvK7Wcj7isvq2rvMwwgW25N331
hEKrGAXoh3or+CBwrX1Fqi1g0/7/2Fu3uRy5LEKoIo5nodJ1BEJfHkTGlOr3
KEUVrknTv6z4Xvo6co6Jimr1FjkdJPdCQSbXS83kfSl91DQCWDoO4oI5kSSM
X5mMT7+bpYQx0AV6c5Y1RRt+r1GW61mG4EUSgVxDDLED+IcJ7NI9GL/lcaFb
iYUtXnJ6JCxJ+ovP9mQqK8LPhlEMdQPKAmuXQcgjvsd/pnyAUXTq0LgkFLz1
F4gR/fhxq6IzleMzoIr6elxuqBMIYDdAWIoFSigAiywEIjvm1YYjairwT+0v
9VYAzCcuEpxQe5SpMwXyJq9RU7k94BWOGrXiGuNIsqfUS9fiMDHxOCaNEv0E
/+IJx+4VVSQ9NA7clI2gFQopX6rhbamWoYrV7ecXbc/m0FlT0N9j2OMgXYMx
ApZVZESBoQibA2chz/HBQgzdrh6Jb+OOw+J5wzJfJl2ldOBdpZ6AZ/hVaDyy
lKpCAnHIWMdHTVTjnJe2EcqapifUfXZzB68/Mzt0mNY2o4efrGLKUE4KNTJL
SLuR9y2g79SUIGGyA+oZHhnUl3m4kJrCFppisB60OOn6aYbmN2ZyPzYjTVgp
+nUO83d4jzSDrH8s5OcUIiyA2LRvV9mn8E3VZnYjIHf4tvh8ykVHrQHSGiuN
s8mfOZ6xOIKMnKzoP9ZFnok7NiWn1mUgFlFXR8U3yt0PuedJDMslv/bXsPUn
YQDROswwnuNzeg+2ckmWJKJdewdDq44k1Ci+l4gthJ02IkT8z3p/kkes6JMr
uZ3F07mjvQot2b3c6/gpeEsVIc6BTHSVqbGeVAHF4sxyrOTCnfoxUYaNV3Ch
3YJPOktLvukOW8URHdwHy5YTfRMLxsLpVlJmJOjMlEf8p/BLcsAgpyuk490c
OXnu47PLY3YG+p9PX7mnU5nO1zsUBO6EZypzBJNjDT0Gw8gFztYJ+OjTkgFn
6WYiTXnQtC4UKAntllyk2Pt6OeAkyL1xgIXMdDRk9rxSLbwFSTrZm5/4Dxkj
WpCMY/pJrA7sqc70zVNjg7sEDSGvKfiAqgEZMX87slmDAY/QW9/EWYKelXxP
g3CuhJUV5miNdcwI4WtVvQWk1Z6LCvW7S98J/HSKvWF2F3sYwdpnM0+IfGm+
uEfY3rLp6LiUy6YdfzrsQFslzhr+ONlApu7rVyTZJP5GpVpMH1FY9wzUqT+a
bAYw4g22nzvVLLbAlYjdoyQYfyeW0bw8OVKOmtw6htgQGcMG28Wv9Yap+BLZ
dv/bkZ/Ttri4RiSmjklwRaYVHQT7HVy/oBo778geDNshLYPkYsAbl5AlHNnS
LFKBZTs6RRoGGzUY3kTzMTPEoWEwDCAonWfNNLnG4Ow9i1ZjEgeIPVfRq7OE
2ayM+ow/NhZ/93LR7rTLYrZlca0uy0TrV1zOk0/iJHUvv3EGyzSj8PbfzNhj
RtgOuck7vl6xQk9TaYGGA5sd/Ng3rYfYibVJ6eQpMXKnU8HVJ9Ok/JOMK928
OghFqnHJZ5HnEufovvhasfKhbT+d3Wd2OBVmep32uKxjCQYn7/9ORM6Re7kU
VeE1XgoUFk1t9DuPNQss6ClsFsPqgsOvDHZF9efNuKu+IJWjwn5sOMpUa6CM
rZver2WYTaSJtbEwspRztOSVF3O9iQ5PBEszoixCRVv7zKqlKQeuv9F7EQOy
CTLMhRbS+ahQUbb5sgW1kv40PuRZKl4VBeOPhoWPTLTwQfgRwhYrFvM2Ta7/
Y8VzezyRhWIEV3tz9FIR6j10Ew/g0L7UuLmcOf5t4U2kMR0QBJZuZVZCaskx
yVmkhq9wp9nWvB/tnwNZOmYmLJ+XWQt2RnDiTx3sDk0AaANTTP1grueGKz1w
EB2oRpdoRECDNFxIwbWdmfbSaOYaPnpmpaPWK1QyZD8As2y8YZD3wIUUU3wp
Ow/+E4Jf7g0UxdElpguHfFFmxpg0260C9nSjMklynIu0Kzy2iBYZfGMzxcat
+3eiR8FvwkJfh4rIO9Jg0Uhbf4YTpHTzYrBUPwJUonak73csKjptbfCq1D/7
bcoog+1UngoMXnHOXHCpp7++CQzKMRSKzWHd+d2K4OwXYw4+leqnnI+WXVkF
J1XAzD+uvsPWKAbEONg4BbTZRXY/Xg83nykS3jYjtIZKLuIYburUZ+YjVaZi
oosQIpSGrtlh2Up5rXLUx3AWs8OaFCjqWMBMGmmK5Wr+T4+Q/fvSZcZCkDym
1ZljlsozYdZV88C3LMqAEsH3+Z9Y/SPNCt/UDyq6eP70G+nYwGuNI2oTTcY/
skpaMM7iOHmPWgbsVAAljoFMT+SO7mKj0ws0D0Vud6/uM7D+dXaShgEg410N
t4i9jUZJgEDwnVblEcboCCxTtCoIZ0QPjkGYcPTz1KAwbg823XfULhS/Q8wk
1q8h0uoKpO+IR9Jd4duzIzrgNPOH8mrClsp70vOsuqfC05I69Xx/5T/x4p5F
il+9UVS2JM6P8J04gdMYKsK9DZC8RCheNPdhOOIR0rgOe5HdXaU12COYvFM3
5oVJJ0wrFh3puE711lc0+qhSyWo0okjpC1acecVaS0+mW1jEAxvfVhtoWPwT
arI0PHICyfNrSxgOilvXOUBDBmIIhhzh18LEKrEao/R9p9mERhmU+umEg0/e
/yBN/dScEZusFUzJiXE69JId+mNu9BLtGDsGlYwFARIalShS2wfo2GxmWuAq
kOowJdQqv8neeBjpW/y5QepaLWLVqU/W+CjAvHON/h8dePmNbDGj5nipWizd
bpqFa19klPmfhO21k1ykECNcE4oOB6zBp0k5Z2qIBcGltgr1MPR5GUnNgozr
CjBA+Cnkvvjr332YtNOsgiP9BwUPsaPDxL2diXNgIPyXx3jhntHbBExOTxVi
IasC6L5Wy0X9jxJXvTVIzH+b8ERcfC6zlA/5aq0IdDWuINY3C8sEq3QGL9wq
wTdrb0CSpIoxQy5PLoZ9JxJfPag2mX8u662No13eQA4p7D/zO6CS5GLhSp0Q
trZnGOUKiTp1lUcIztCGUJFxclKmRaNbonHVQ8ekJMviBuhF8aCe6GLl4wKA
OaPv6AoG3Whzj1Xg0bSruNp3zg1+ihDyj6r7nXLdCkn0FgPN4q19VQHBz3JO
KTki1F8cQsIurnetmEK4rE9USlryXNyxYRHrZb1gqm0dL3rCI/XflAqF3Set
1sTx9VzUXqA8B/ZsMigsUN5DHDgybiA8XWlOFDz8nfAD1aropd1EmJ3/Q9TZ
V1ik0jLhGeHgS5DpFlFn90/yCLGH86IPEaqer++Yet/Oe5b/H6GKu7pWRlI+
TFb1TTeDUrU7p0xpNkhe1VaOBrPIVPE8ubPKMp70AivzFjWvqq3ToNscaD9Z
l0H5kW1QRePQfVSyFiiJKAkqdszigK+uWBZ/PuC20P1BFhHuBzuio8Y5IN17
mzo1o5ScSTbBxIcPJCFyanmBu2wXXzMCIy4lazmbt54HQQMSGfHk2pNOln8F
RlNYZAINH6q/gbHoGy4GckAId/qTdymMW0pgGG1+8JpHVNaa3MNCsmG8ck7Q
9kj3yhYUC+ql7SasPVVftRvSkIrNFuZ1D6zmLCSUohQb/wX+R3aR7TDEW+6F
Sx3C/nCAqEBQTD+3KWeNtMnvu70YT8O2EosOSNvrM3BqgKy3HbD9/zof0si9
yZNYe0yYmzr1rJhLiA/N+mRTSiiZrsVc6PFZoXPtwHiMYotQVGEbsNJfNZsx
QCSTx+zPAYq5+djuRZfBSJ6v6vEC8SIb3St0L9usmARGQYQ1kgiV/AIEhYYG
M9+Mw65XIlxsu7v+riC1CNSu6mLM59rbD0HNZwsEKLkroi7UThrfe6uUBisc
aIFYOahPe+NzwJkm6pbTZue4xYUqGN7cSm+4icZPciWYBLgz12C2k3D0H44u
RCwROW4faSxUIZND7hLIWwn92upCDm2uZpoGEO51/oXJh+gE0Pc97j1pHjMa
CKZaRz4HkgX3cMCX6q4d7YlNqOfXhaohQ7UduAT7KAOcMRar2LyexIzsl2li
+1PlNcObomUhtACf7/9qUAvwcafptnb21YX6apL8cqOSkhXN7UbI9cNmmR8L
ZfumV5aV4kHUY1bREK+PJRD10vs1H/85u/RnyKla3ouof/7rH2Bhhf/aeenJ
r/6tycjzzFa+vGyP49qGht1v8B4axFYC1IVK4UqJr0zx69yo+VWZVHn/DKrI
SHyctAsBPCoQyWeFTzu5Xq8MsKo/ouiUbabKBe/X5uH9XHPQxGzt0Szdq62g
nOahpQxWifTCN2vhBtmMXVZROLjNXPnWyeNJvYvB1fOPQg0oTpiKj7BPTfyB
2KSfvEcqE9hDUd/bD2n0PQI2VFFDgcgJaaDDMa6PVZ05w3NhXnD6Fqlj+poq
PuCZm7kO42Wc6pjuCZbrJPjnlbWP280LRY5e8B693LUpiwIWoeMwdMbFcbgM
03Grp8MedYe/lMQeRVScWkpA2zneB98SFjneqZkbgZ2Tg50fIx+yFxDWFONY
cK3W3LIhAxIVRwVYsWZXGKn4jhVoowE0/mY+jUCmVpK7mro707ezkCJNAYMK
d3B6ZB98eeFqAy+9HiHwgYmIfLUW6Jy0hzlL4NMyZXZZrvAPqEmNlQMLi3Uk
Dr5FYkRqfJBnH48RRX8jHq067NnGJl/Jv8ozbfZGSO8d8G1825UxDAVzGsx4
QX887GZ4EVbHP/OFuxLCNcKaKtzpwW/vtT0VTq8ap3MXNmQvJxCGO40Y0TcR
JHoAnMoyTsAV89LKetNdz0Klv5btwPsKIE5RjIvLWJI5bjOYO4MBPKOJrix6
mgOG7KVp1QOqcmZQT4/SSme/uOUXzW7VMlFjWXhMo5Dk78tYiVm/vB8QsimL
6/xjExP4OF57UmJCdjWczVW16i6ByI5dJ50jq4op6GmlWUT3ZI4P9kcIuRyB
qM8TuqGHvfaA8ttXVwrRz9jExUycdHgQlodaOWqwrfqA8h6AQYxNEN3aZvX+
PWOJLJLVGkKhNp/fW+kk5dwDv4Hb5uo0h1WpBa8lfTUnitVATLzvo1f7h9e0
aZbWlCwinz5v075qr3wEcA0XA4Xb9SVmDowAIWUkoHz1QKpQeSp8RjjLmy0e
l9Og60FfOJfVrZZEuHjsNtRfDeb07FyJEK873PEyBtc237Sltxa4zrkqP1kF
SHu26/agLr5A0WHADXIlppCydVgWDUhIcTcMZvzvn7qQZ+MDupm1OYekE69R
Eact0JHGX5yq8PY7isUObxJ6pVzEmahbCcbyi/omoEKMExhbnYYwFtPdeKfC
51lUCxQOiJLSN00M75akqzRoN5ceGMleerTFueGLNwMw4wqvGnnIG/IuUN7Z
ovM74pxESoMB1uVX8rEuNSPjWVKg+4Q1+CkpebQxUZQJNBTCB4wbBVvI2tNi
S2oLWgxUtJGoC3VJ9B3FeMFTRjXu02STXngj0Q7CVPFdY/LK/QPM515Uuzy5
5f61S09sRzYWh43aqNcZ5lp/R8fKZyKGdouekZnRC5BNbREsL8GCJ1+k1tj5
zJGbmMbOkDWJZaoaEZOeyqTGJNEeNAEJpzHeRlKQnL9lxTqiyWnNzHFKtwVP
6xcUEEY9BYqKgo3zVEE3g56DIPpCYPDrQdEh/VMEfVS9fR5gE33odY+UNDUB
M4Fu93qoXNyOvgqscwF5kk2ReraDEmXY/yesTx1mZhOt+4tMSqHfJWftVAQ1
rJpANfZfQNV3kprPoYX5lUcJu2zyKXCNrtnuKDzgnlTa+xlsO+GQvNnTTXdP
NmtiKQdAGsp6DGRZ5fkFiwxrjZC8e0h+ILEc+bvistZVhsi32lx1vgAZFLMC
hifKOmlkL75g7uhW2SPWmekShnExerg5KGcG+5ICESI5b9Xnnj+aX8bQO0lV
PcPopQi5bl7IKR2uce31DFjg/Q92UCcGVPOwuZAU3ZKQ74WwvSEhZFUkEc/0
lHImsk+mijuQL+1Kz7jxqAxUr5GBhZ7VjKhFTn4UMT18y74RRPPQB6Ygilbm
0TdRc/T+/SAKm450Ji6S4oXvBb8+nagF4aFnOEflwKF/n3E/ol61OSbEInYG
uaBTm2cqELhkFbhExIn8Y6z45gW5IZII3EC+SL5wJFDTp6hiduCi3iIFCsAE
LE0f9U2hYXNsbcTnXBK4sijX+rEArJRCYSY9IGUNlM5gkOmQ9/aD1mdoh68F
3Dp2q6dsSUw1FKDcbbv2yT4eWl30CftqrsUU7wSadAPn8iKNVuxNMbgCc+Sm
hzJjR8q4Yog91I+IfsXOmcZmS+Ub1xS31Ep1xFEwMxDRi3wsEoRDYaslCAcz
7viSuHLoeWHjFmPdF9AoxjXIBO8eodwCyemS7mPKlEAX1aPHHseG8WAMMS/N
oMK08Zu5aA3q9h2vdrN0ZYV/X/G9bIedU0miTIpqrojZ7c9PX/mRuZWauv3/
kQDuWLylwD9+BrEQesv2fFVpEtBF1DJxdMd94ylxr3+NucGoAcA3WlrtcQZu
xMQB4yeDJ/GIip9LzaujTJlCCsr9wAd1T/ZFKzLt3+k2/92nYE7qGMxVTfG3
xzhGSi1zRNop+ldmQp2YrkHBOKlrwisgUhSgAxLBxUObCrmMoRv8A9nNZqOy
y4e7MifOYd636OwjiqFWbVYGNvfNBLG7vw4uecDNpiO7DwKdBezsYmZGMBKC
jZALZVdc4PRtCEXzkJmZ8zFUYpwncvBYQAr/frTTLwtIeeCciYG97y4ufnNN
C4hjLaht6BepVBlRmEW1Q780fe0mDcFvLiMjYgwLD5BGEluMGMjDxjnFAWjm
BWUXaawaZgQsfI6L3//8msZ3y2+e2m8O+q6sPQM7BYm3kvIGbnuPMxd1o3C0
Hit4YSUnH6s8qJk4tXOs1ygritjEHqvrx4zLwsFnUzS9v+ULxaNc+JPanB3E
1V5QJArkBx5vFqjMlzGMrpBQ3546oEsLxekuvWeqkc2kvpXHdvAuQToDLD/Z
krIP4eJHKGWejMETXRapIsi+E+zAXKrnzfNog55lm8sHnLSXSA7wP8PK8n8t
IS0jr+hEG89j+d1HlGHRYP69PyZQmoB7c5Ht2GbGN1nq9wGrMwCbP0kzRuQh
q6JZDIkvza22zYQl2Hy9Ur+VtZkUPDY9Vhj3MPsIeqOmBufyPvWg6z8QnXJW
Ttp3jVN4Wj6HZonBjypRS7HGry56xexO0NYN7q629ElHLJstWvRNt9ixGabX
RLFUrHe5JiHXAQ7BBgUQm/4PlUDv+AP001zyti8gNxem4wuqtdYx1zl3Gk09
TDsJmNPUD/Hqnw4lS8G+rQJh7d/wpHEim+DMVnwGoLj/KOBTLFn3EUfAovqS
4ivQiIsMvCTr2/n/6e06/giu+j8F2F0sTk+MK6o+g3PVUbx288NZQTeQY9CH
ZZAzY5RE2VAx9iE817hqWt7iWGNLAz+YnfvN/augq1uag0nYPrmR2ryTLguK
QKyGaOUeryp4tbYO1reR4ZoXGi7RAa4/j4jwkpvRIF8eeCnD+pVTEiG83aB2
LwbM1lRheSR8SUYeUufgMgl+WAwaspL1pcK2um/qAaxp6iUBwWNfLunhHW9N
T3ueKxEHXoNpwIklZwFC/HKruMTAcINTz3qMmBH0xNBGa1YQ9z4zX5nH9XGz
O9GKBG7aBOtAshOGZ4mHaprHOz3FyoVLIqipmSKPuguTlmNTxTiU1nMdcR7u
AU3u4Cf7Sc/46FcCTn2idKke3HH/l8zyPWSmUBw/3QzF1pEDNFTcYPgY45fr
R8PGuHO9EKCUx9IOqP5wHh9CPg1617NRIpFKVuX9+0ypyjhK/L6njlHCoEaQ
cg8oWd1r906AhLJvvU9Q5/c88PoOuXrtQ8VRZwLRz2s6+amai2zzyxBEBOnC
w5ZuvWxx/FbO18WXi52Q/G94O7DIoMvUaWMD7MfdSDwwaufRmdO5ggr6f8Wr
/SX8n/k9WXAt+AGrW3hLsLMcv8mnJHELdrYUxtCFrgR0qgoLQyQzHBMIfROu
bYbziYFhk9r1EAsS5VFMNahKKN2FRp63+4aViCB2v2SLzyvZEuQ+1h5b1lrS
MRlyaeI1uzt7CXvTOF/xkzH3M3Q3atjNeNdcdc5S/oQvKhEvorJAHwxpAkP5
E1sbYhfNydZuvk9LMGnikIJMXX3aW8d2EX8EeGMthP9xjuuTgUefxYsWWuQx
EQq3GKoNy1qwFg9phdfbAqsCYTRsxttI6xgHsfzL+tHtqKeqd4UOUGSfTOG7
wm/SddM7f6wNDarwJ+Y1SbSl/duSfwiHspit0WO2Pq2ab/qAeB07/5fvPG1j
mWxBvxp/JXMQgZK/mSAVCPHyHXdXUXB+CKpED3ao9GyGi1i+gGqh09jazc9/
lOi7CnUv0D9SUweD8HQLqU29gh75b4g8UFasp6xUTxnCL0m3XXB6zPEQr4gx
vhq2Co3qvFYe8NdSqLgH92ExUkINU5ZGj2ej+B4+ZfdJ/DTkZlMs/pHWtaXP
Q7NSpx0v7HUxYEwPoAxwA6wOMpIIaLo6D92rZoLXrTJYStsqwOFfVQBvEerK
J9To5ThmwO6NwhBptuvmbkvT1KgWppkdj1DZI0+O5BJrFALEOtb+ZKUZvjVs
GLVPoQuADH8rXXz8ZpiIycRh8o6FwZZtu7TTLh2/tVb7FiFHvh4MlqVolTy/
ohHURk8Ima3b3LBZw81G5kvhlPxa/XuwdD4K0cege+LV4aWcBghT7dbIMdf2
BiEyZ9zq1OCopFbbx9kWmlaADHXP1ApZ2SRf/5BPTzM6lHD4JrPFEqtIzM8s
V7U5pAV0a5gvBX47CxcJiUedCLEhFxKw+drnnytF/jLqvr+Sv2cBrMRcYgsw
PwPZ9vpaIx2Jy9Ud9o18AkqSdxKGtq2Vwxs0bJJM1KpzxH9KweOGpKJhELM4
AxY7z9RFq/xT7WOWvi43Y46B56n2LqFYznTUb9f4I08122Trlvh3NEU2E7JC
UBq4itabyzYnhSAXhsMR4lioG1LdmQ44IUf9g5jkrznGT2TXi2Ag5P6K7uHu
frewRDrxelBM3qFhBHRF3+R4OXKj9ugp6F4ONqLBjfH50GZUEKx6+/YpsT2m
AqRxrM59MUtkWoF6io7T4Od27PJ/93ld+yaPzCLC0X518x/iqJNxEfrsY4Mq
EGfqmul9iXJ3LdqTvHVMqV2ChcUDEfjmo1d/cZKOdOWpu7Bhdni/rCh2BSu9
BQRnv2bHoVZ4j74QGgfo5iF7FW61NFojOF4Jjsuhl/vRBG+LRoTA19sUu7ah
1g/bsv4CbwcRrI3JWcHZXUyP+8+UwXSqA5oz58Y/CrhrcN4e7gs0c7sg644X
+3IVmiohbQ7tUpO0hY7bXxsRcODgEfLExLG1x868O6XNdSXTrZ1zZEG72RAN
EO5qllGr+GkggTdcv4n+ZZ2Ny86AqTUgKw5iSSbbWhu6l2kRieT0Go3ou8fv
mBFSRIY3gC82+ceUHovDZrA5Su7/08sOFByRqVjeyGt0oz52UGfK9J/7KlfF
s8EEilnBlo0wggnxLMdT8LxkXesYs5nZLNmOFMaLfjAxVyRScWlU3RC9JgLC
ph5uJu0e7RCeuj2ra5umv4EnnRIbWu7vUPuQoQCnIkR6trn5xWs+5AhAXiUH
FHdaKQFuofEM9pO5m+HEHD3RfdXyWO3wm7bq0iHD72uxZBgx/ywwsoydFIZD
PYNFNQZvWgyPOAyi2Radclqq/PLfXfuASyfXAT9iLzQtPu6b5AwYcW3sQtOd
a/PpCI1tC91NYpDsuZK6R+F6xuI4+C6bPCfUiH8LTEQVHudFs2Ma0tLC2bI2
ydrmecKa64nVBzpWTDc7lujvauGIXSsVXwzoR5yZkros9ZioNhcGceJAyIsJ
a+IT8RD7Z8S2TrSriIskqh13p1qqjod4V2rJzZD86T9Gm7HdmS3Fz7tDF+GO
/qOZ6FLOLLv9YYBiD51heb9j8RdByybuyr3BspSYAFDne7CFqBK8SEQh9HVZ
R5k1qMYnFMjUTL6Vy6Xie/fGLbesj6dCO9LUFEep2g2ky1JpeNQdeVmrsDuK
+cQH9cAIAbqNmLEj

`pragma protect end_protected
