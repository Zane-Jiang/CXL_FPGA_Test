`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
TTPGx8D/FNN1wJCf+liMSgryd5UBSit8DnuJzPs4S1BpoVGRoWi+1UJjJRnntgI5
SufMs7HcpOS71RmiK4apiTgk7IpchWepuLB9rEwp8YPMfWmvAUYjzXidH4GxpoU+
RVdcsU0Xie68opcWyETcDarn41zFOR7uE+6WfVkTVuU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 37184), data_block
VNbwk+Vk3/iOJbTbkqBCMEfJ+re32KOv2XZ7mqoNIRz7U7AaKoD4BbdCSbm4q6K5
NoFN+j7jjg3bkQQgcP4neWYKmcjWg7gu94ZjkKvy2KuMiuZJYmkW2guqJoPyEbOR
qzdIDx1xL0kXM3wMi7CC6PjWGF3z9Ug3V+odX9JIRuZnq+pLvy2MVGz+d0M80g45
N6S5utxkONMPESAp5s3aBIWPtgumCrUe0G9u+HdoxByljVejI74LH43xiHFE71QE
qq6Jp1ACXAuMYhEjrjj9Xh2OrDyiqunYcvBzrDCB8FeXN3b4B8PSXGa0laGYqqfL
YclEoHmIlhNGAWbdsieYFS1Q5KHL3rUfsLe12I9tWwQrINDs3hwurIrZSh4NqdnN
kXB7PArw/B/5L9TJejJyatQp/oVYacyslq/jyFbVnCDzieKElGpLxb+DXeIUYEUu
W4Y1pD29C7ajy2OIRznkbR7kUcBLi4U30esqvGmKZi+Iqo7isYpz203wX2VGZi2L
4O9nezZwht0YMtgkIgXr+n4AixRYkbby1KtJok65UJet7K642IRtSWqP1XvbifHD
rCqnhtmRhT6zNxrvD+IcGYftO4ab/nJaKS3I7E9pYfcupUxXlg2/n2fXul5cqQmN
ECG2S8uGXVFw2jmlI56852otQf/iGdmXpRndo42FURqsmMEyF8FvJlt1zQlGQRKl
sp95LmyQ3mYHqTCJgBe2g4nQutgwqcspEINgxF3RduYkS+KBTErXxvwHCrbtzRk0
JKjwE4I2bPk11nbUP+aEnumc9JCMXUX7ldIJT/P+ppF2OOsX/uA4Tg3mk1eUmkN8
yd8rx8+CGZdbMygWr8SS10qZibNiIvCrN7LUXe7tPAwayQCEDc5cMp6MNIIGQeQp
OlwdUFvhZHGQ3Y1VO6C89fnqpTuYKxlVbUkCvzaxhWwcYNJp4b/OPcQdrcbvEl1d
PMTZG2Z4J//qrOS+R959IIbTKvApd2X0WVvU2GUhiT0ANA6AhRg2u0i9REZrS0LG
mPvZlO1vNRQqYuDJBamRQ7/HH3NSgmvFWsLUQnrBWKOWxO2eLe0vLsCzDDR7Fs61
uI+a17xe4tzvPhNGSWN6clkc4x9f92lQXGtkI75S83kOBBXRj+UNdjaj/AY38x2r
vBFNIbQLJrPVYEo7sPyggCH+WKdqaNcnQvM86dA/BqcWf5cRY7NHcj1aH7zXJ0TD
JIlM0pZK99Mn62SNiKR7FqtPXm8QHKRtKfBZNTstK8fdrgqTBpSClHoIAZd7cOS1
LE+yGESgwFPb1vWk2EvqogGxXg+VZKcgCvhUwvQb634GxLdH1UcoenLz5XIh0CK1
BTxOQo+seMLUhtbehhysmufggz9NFdQgxvv9YcopihqZyi90dRn2grf4kAFJ9AX/
zSfCmWAm1193WJ71wHgjrAqA3YBMas0LYK+hh1FBlWf4rTzv9sv5OmS7b7cS/C6M
cftCxWUoPAy7ecG6yaSIha8XYXmAf2ch4Jg5PDeu3qAQcs5ubUjTthjx9AgqJpH5
50sSt6YaOIEeCXW8TMkbPRzr8iEMpPKX8MlEBVm+RwXQQ/7lxLWRMYQBAmF+he1n
VgMQOZzqvjgstwtVKV3cGoy7C0QUkhBVVNRq4ONG9vAxCknRI2E+ZqDRpocu0xR+
V4fLlv8gGbXfonhjZLK1VoOXtdMMNvxs8rJhyp4rMagsaPtoz3u92r1ALZ2+UBLT
X4oJmBGhghvroKfyFS9VfoIga5vvQHL/HEO2934jCXMVQ4JKzWT7T6TymBLzU9tG
2WlxVCTy9hRSAAE9PcAwi9Gp2pc8y7Hb/hjWVGkGlkAtnxJ429ATv6HC5pk5Og/3
54rx7gqmQth6I7IbPzJbaiP8PZWhQtdAAyr8Z0OykySodtti7kVcB3v4S4ygEcxL
VWeMjwkj6feGoXoWqsl/6UhG9JODUQXks1QVBhi9gzcVrigCHf+ISEOyNjzIr02s
3GwooWGeMO9vbLp1KRptBvCxq9G/zW74R50k32qs2dHnDf+20ELH1S3Z8CpdvC7h
6KwqhK3weYQaCAGQSlyTDL56enzQXU6Sc0PGUX17v2ahxOtOOC9gpK5YZSJP1iEZ
i4rAyeVE5dXqGt3gKBSHx47xQ8FgcAJ4w2VBLtW7xW7hvaBliy4ZZF2cS48NRuuC
MgiNLbrrHQEtYNQSZqc5SRCjcryALa+D6ctXi8en104/gzKfi+PFqMESJmMbKOjR
z0VOA676APP/XNSU+MK7THAGfNdXYWEZl+yXrj4ZN2KeVGpG43Z47HPmsFArZTS9
GjqI6QfpzIVprR5B5yC0jl9IFbmimqNuqgwi0bogQZooytl6cZfAuOVDCVMwfjol
6HRr8p4QRi9iGgP8daf2eHCVT9ZXDkq8MfGmJX8acnav5eix8kxRRUb26c3R5kVk
Xqbu+BgmzPFBKLJNrGTD0nw2h6iXrPmiaL5gy+868RADgZ0rnJm6ikdrs03+/rQM
8sxlP4cfQVCLSGP1rc1Z5wG9zosonb+0xAs227sOCKkT9IoXmsJ7yin7j88pDK+K
te0BUppclGk2eMzxKu7X6upjVgVfh3I1u6QjMLjguqKMhG7bjwv9AD6QKTx+Y1Jp
0tYY1apZpYUwNsvEafJjW0YDSoaev5AwRNJi7mr0fKnuYF9fm5x6NIqRj9pUStsU
erhAGVpB8jAhkk9ito9OKr+lTdd/m8cEC73WEC1NICWCUHxSUMg2G9wZwkia7ayT
RjOQ9ISoovuUvS91l1k6FdXoD2dnzgj0uya5BFkB2HSocKeXL74aP6XH5B2KwON5
H7eZU+EPYW42wPyk1NuGFg8QCf81E/WkTWmjQF43wbix1u+8v1U7UtaOovbgXk9o
l3r+MMgTW33bBFEeGkRsI8iI+pYs1JgNrfnYJAn2i5G2SasN/n9lPMkDuTVnqazd
wEx8XHdrhrkuaaaKw0XPPSiLG1++kpleOp9q17wD7o4eIep/HXtl3ejw+RDeZ8oz
3EKwOw11PYyWZ4UjUqqL0dxYV3oUv5am0fJsq3c9GEjQgrGHOEqv7yls42jDlmkh
E7/rPA2gEG8H9bd/n2/GyuFZB8oyJ/ZmTU9E24fQaTUM7xnXTHOAiiEfRXJEG5+L
ue9yPLf3BvX3TengAMZxQWio+VH7GqAXiVBR7amGJK1CYRbDruz7g//1NETUcsP4
1ixvdT7AdPqKzoUhQUoSvN34dI63GuNy8RLGIcAsQZ+99XLWzfwKZZM6gHD0+DOj
HZ/cPFlFtsZadOAfknenoufB7HVARNePv+CDpU4ltQFIg0eAUg+4MgRY5DpDmEoN
v09vO7URCQ9zFWcwkjI+Y8pv+5K94f/FzbGbwbRdT9TVzblxTHsPKshdPWbtn1WS
Bm4Mec8dM8UbqVFrT/gwAygs2lfs+/7msogrd/gN/VBYxaqoxVOAEiDf3PrdvA78
iko03YGr2j7RA9BEvjhcoC+rXmDIYutMGUQLFJ+Yeza7upNypbPFDYXFxcYSa1l/
rS9pB6r6aD20oidua+FKzEQ2TX/RxSG4y5rf8zPBY0uQonG1pExoOFjnUo6fSfaV
sRO4p+HPhBsN42M+xRpeVlXg6oBQR5k8cMN4bdDLHaX/NPeLWgkY1HST7FPQU0c9
Di5IROiUaQWtbzNloBz/C3AUZPg8GkH9fyLZALudY0Zds80WicXKu1DFHB/JfdLl
AxHbhKlx9b7eXzH8Da9SzDp2HOdEv/kS6oQt47NS+LxglZcYaYy8I5Gb8bCtcefj
ujiGC+yjP6xzrGsXmqVvFhyIcNU15I6SD/CnXBV8lq9ALm9U0++s+wejapw2PEyU
Tnj099Gtv+xkP539ZHteTWZwbnc5A+8TMic6vzrHIEocfZiqUdpHrvUlh7203R/H
7SDONjiG0Dpv0Q2m5lvInwex1I5zgX9KVTzcf6p4XBlPzRdiccDpL5LCmT2S0zlp
dX5FLs5rLpeAEuklxd7kItkAir/KhIyPYa2chGXdVo3wCbwd/Wsew14deMXyrKNd
psjMudgY7GU9emXTbuK4JNraOG4NFqcqj79KN2SDKzs5mYIOs/gEtHBxcoCgYaRw
11RONc+jCkX2u4EUa6GMfOCuThoqxOBjl/oWwUCZVLDLR8zt+aAG3tBfZRaNuNuc
Zinelu/0KVmqdJFRqq4Vpt/7aVsXAJi5eqWn9NINjce8BwzozoTefUkAcNss7Je1
Lt6lj0NCvSHvdxmT0vHifKpzwA8xYgLVKI3VFMqwLSp6oVEWQaxhCM0mQlP2u7yz
cNQg832DxXrwkSEuoWmy09/DwodnXbAwgM5Tqqwz0/qvA6qaMetHHAm4G4gApMnQ
qaC0eyaFXS0SgNwbU81nEc7bFhIHK/nHjY1PsTmnQcJRKWHyYUb9cFMnywHWsZ31
yGt4uEMVuYxExBsF4cFv/+uB2WMKZk5+E6PQEA5M0L0lAvI0AoN2wX0pPQ0C34T+
uz0lu+mlacmiGlBH13BwRbeyZkGVBzPCdX0LJqhQKr/SViTiLt6pGtrCB+YgaMpz
Jig8yPAOtujVW78HphsvKDO4hIR2JuiFa2LSiA+uy0FOtY4jN+Vi1AtzdNXxBx4B
UpGW+N8jQbuvD4bt92GQajz+ZWBwxCPLnFntiNKYUigrTRhGYz1vwDdtb29hl+6V
yUvbO5MR97FKZf0KlIkJWdow4X/22JnFrNSKfuLpGT3aypngweOwazETLHEJxThM
X2352v6XJ95e+sDekx6ZlX5b4hxannZB6FBfGaRBwXNZFMz/COb6qiScmAWpgJeq
hQjkfO23r6Jv6ArjSmH5MMJSmgWhfFvqBDfuiybM6qvp9kqdIcFAFPI7khN/zgB7
HahGSUWliQkEnXimfEibGJ1wmRqKKei9zTx5yDzCVh2f3/S+Qu/N30JOAr/vDt/d
TJFdy6QDZ0QLtCJFUCogtamDqL+Gw0sJixRkZvQkufGi8GOj1qfNMhA6TV0cHXiT
Hy0nS67VQDoCpJNcAmmc4ZlKIlx/58BWt2LffAJx+w59piQwDsvTK+IsuZE3otny
lt32QTwNgaBmCj17Rz+DW7f65gR6uGlBxvjCjM5xqu1i/exGdoQwh9IjJq9xkndT
RcbfzAGfvevUKlkZiFH/MrBTJvUMkLSf3s7pfS7kx++OYjBVdP8pwLx6GJ4/25qK
ah9iF9STOyRxRU2CzIM0DpXFd4EzoQNA0aNHEzZwZDUdI3wpTwlffiRaADHxzE99
tGKePMYCjgrlosmbG5hIA6v9gdAm+PabX5SPN0tWKNqZcMNeZ5AlkPT0lhpx/Ni0
DNv1uwfci3NZZRzhaCEl3kLaPQDSVrwY5XV+DZr7Ao3UYCfvhzTJtIi/+DOiqXOH
V4SnTMXL5Y+Bfkw0ApL2GyhrJjWe9ouBk71DnjXbQS6aDnGmG9KYwMthwt1DsPDz
sBgj35oGRdZp95KRxNPtjXPRfFi3HbpwkD+yd3D2/SJRKP5s1Cl2Bz6VWcvairCk
LypFL3McMDXpj+sPdHlErsGCXzgHiu0kzPK/I9BKLywZFQROpaCbCiMLYlnY6USk
ysPhGe78XWZFAINqt7mioM653rGfZyYTyQOyto6m43fgJQVB2a8kuXU9u2jdJmHO
S4HVskHwn6bzdJolbsOWXXOosVOLpgPiOWM73iwTK6LH0DAz2Dm7Ha9iK3lGlIDL
DjXZTanXFTkEn+j7+scBkRAAH+E/qEZaTg6M4slfcEG/ghabSVD96zlXJpaMd+TS
eg94FrHxAK2u15qJAx2wqKVvJxE9OUNPgLl0hSzf/DqUZpQCzdyDJgUHKS/JxF6R
vJdqNdNhuIuvE47jAF4964zqo2BY9m5mdM3vamTqPOi9LZ1+MZJVow691PG4Sway
YnZIXEnBAJjAt3BycrBnmrrfr+afar5VR1HOZJUZ4Ak6OOdEfkELlHZ/3lpW9NmI
/i4W21wIn3O+bW1/0G/G0gsV3XkXu/YkToTiPfRHyvDSFYWCxZsz+9vbUCJarWyS
sOi0AIG9BD9H1bKYnHadTmIevph4gPbZUZayStjnYL0oZlFLv/rbv0afwJA1LVvI
f6aWxDHL2qxVckdr0s9O0gro/UjgtjjInwP2uHs0qNtJermRoezm0Ou5sD5QwI5v
nkvoWgUJY83Ipuk8IgzlQVy7wOfg6ptRADPOCjP+oJFMsauJ0BTjTZqkoPpk4iCL
6iWfHgdZ4mzZ97ZNavKqODdXim+tfuiCZOG1DWuRo2RXM3YD9ZgDz7pm5m3yKCW9
N2mQXxkmRPSIi1+nmDAmQyb1vgm1vs0uc4lcaym58714XYsUvUQQWDathPRnOYZL
PLQUQ+zMh6cnAuenO9ngSSDdFXetUG19ZAm5RSLm3m6U/dh/ZHz2D+Qtt/PpqVn9
0cykx1bNRW9LjQfy01Dfs1UI8266e6Iwm5ez37QUQTZoDCIBh0lhTlD8R87nt3/6
NVzGBbXCsvnOoyQ3aoa6BmU+rUKhXzrEbqiL0mWL63PKAEZ8vzrdgHElQuhdgURe
Uokt/7ThsV+HTEe9qSnKOVdlciBR2rnaGMIYv4DSdbFLQROcjApr4VXFc4Ldhxof
PvnSD4Z5Mn3sOm/lAMorpg6dem+kpR5rzeRKho5OoTFrfTrehaW3ICUESrvFx86m
xu02S6JE+j8DbxHgAzeJ/uDCXRFEaJ6bLlLnJ82Nqul7iEXJYcl8KoWjsDz+tHFO
LC4L/24BBh/9TttAGeZ5MYs7dcqP9VP65yvJGoUphYCaTf1GXBOEgOKTWwjpd9zN
HAyGQaHdvDtvkSpfGNYEFvViWZonCWcSvCcHV/IdVyLkSXuHCsGRWrrFVcJ5LFDq
TlOPcyRU3DUPpe8mMzSKRPL4KWiSlWaqbD8N1yjcv6887sJKXazwBo6iUf7ScqEI
iLliLYVyKtk2PKw/6SvA/Wb92e9kOSaclWl7TBgI1FKPwoJFjIgArPfbYdXE9hm2
jSh8u7V1LGS06x94c2Jd8ltABtFySfKC+piEqEQ41rzeBKb12mU2UxUzK/VxEZI4
3I5I0i3R0SW1wLMQ308LDxEV5oX30YX7z0iGIay4YYTu47BpjE1adrTvng7XFtY1
UoD36436Ht5HBzMQDS5gqI6cQaJYweGQNruNUgNUEb6o8+gwqVOoqWVdODxJD9O6
SzUubFMFEdkQWjvEjSfpdi1uTPVKlVLOmL5Q1RzSPL1j3QB8bI3l9VdKN+uCoRk2
U2o1UHlblytmPuZHmPf1WAeoop6aSpP6xI2yRVOOHm88ayybTcWSfNjZRSbjWNMz
uBY2hGABwaCdNwh0d0auGMEXnDSbZ5WpyElcVBKp7QfhY+PIOh3AID0HQ7ufw189
8IKrZ2D3FbGQNe029wDWiq8j232Wg7zhLEOrnW9PkzMdYgZqibne0l2IUb0bP1rV
OkWF47QMyNO92C+ZhElrv/7xtxsoxdqjuPiVRqUpZhw57Esn4/bgy5zkubOuMgVI
DSi9B5lYBUGn08aw5+Te/x8z3zZAW6b+swBL8DEjdT3+8kLaaP/NpKt4y6XPaf1x
bZJ/RPc5BwEd0+DbeXi8NeemXLJCc/lMFMIuuA8BL3ZK0iyvQ+KjYxaPUCpaXwZj
xhCR7OSon78AyGSYAiW6mYPRQHte8AOY2/vgR7vW8vvFFWDupbJI+vtEg8tTmxo+
OR16WEE2KCTCT2sQc6w4PZeePIGQ7dq1BgB9pkcrxH3quEEn4aZkJad1hdzLODSX
hxIGQZ1H/MsWboBrw8/OlbZ27OvPW1B3qn541OibVvmxApuWydnBL2wU3ppDbe/B
MPSLqDtt4dQvOqb4gUtRyUdrahIUrsN0G5X+mN5knZbQgM9A2tKlLAzGSss3mmdD
dGMWXSZdkBdM9T4EAGoKoD+S8xV0ahrQ/4igPgrqh9k3etXnXfOBjbdI4gDDCgPR
ESmmUrysfIiRgDUBhiDtJbHcdHReF8CdVZcjKz0u2hhfdxqqSByCsk1WvYdU8zgG
upqHPJ4nKt64N1O7R9Gxp1502XjQ7Teu7kX5/bjC4yQ/ER+4ba/FXD7a+qvSLqZj
WCL9rY9wDD7GE/fQ4Nhbvyb8f4mYHGQ4RgIEdWe/JagUHRsMmWT4rKUPRhI3Zsi0
wxe71//DjHXy0qQ7vNh8puWaXwYZtLXnKC+0ZbfkM8YLWrmUrLnw4c09Ljn10Fha
j16lL4u/hcjJj7j21L5y3bxNG3yu5RY/xIj7SQbieGIQful3jTQAfwtoNDve6Lyn
ipujvstjwUwDBVwOqsEzBTWwXU0eBr+tAFTelP2NmyWdmIMJOSZmY1vM7I8+K+cE
+uU+KFnLPRlf9Ynbt6200qQ2LqlCRhLPqb0WR6m3iNYUEk3JExtbbXp/lIDEaUfg
KAFK9rwSWWrleQX78FxFEivs5fMSI4E5icK3L7Jtfc/3Iaw03C7HQkzwnrVOlDhA
pNWhu+cXN5APtiOSI/JcvJ6Z23kdFAbGY7uBPDbTjFJzNYFE43KrQ+sfrmcbaGp7
7Q9e2/Z7v07mr04BeemUUwyPst/W40KoIqefEluP7gZPvy99AXTW5/PI5hOt+cLu
2FiiGGtMC0VyDERn61g7AwXl3Bj9an+ol8PHOZAK2NzDeI/P6AYuGWoIvRKRjLVi
SkwF8GBSc/7DIJmMtu8otw55D91vKfkZQvZllIxg7ajMY0f5WM3umSC20tIhrN+z
z0s6Ws1K1jTq/8jh9bPw0cYlox+8oOK4wiYJL52dcek8n4B7IV0GEPhEh0pq7PeC
Myho8HX4tet3p5+hKCDITCF5Hz29Dc2nKETZzqMI+o97nWeRcIlBKLe1ZewlhilE
spPSk+zRDtZ6JODToz8UqKbaKWPnoyieQ18evnEvyD1DcJqSI67UHobDjkhKBz1F
k51tu+G1tVcuTvIj5Rf7feQ/+FBghNsHN2+UFJ3arjkoETBos4+2eRb7wdNzCzqA
hivWm3EMOyIvEqSWvEFjcl1cCzPHnYX6XuGKbuThVq6w3+oneFMKFXkmvBgpC9RP
/OFHNdqKcQD4KaPBG6vDY32zwKm9i6KW+phYqUMFY+MmZNkpjXLHBedT9otN6awG
o8mMSjbBHqOA8zvwowPhDBmNS+ghxXHETHsiY0v3v9y105NGwmGa+SLB6SH6z9jN
ri2JLqaTTMIWxPt8K5wIDL7APNbwN+hhH93X3qrA+8wfnw3s3Sc3LNj9N89HGs0j
ldsuIyNPBfYV30NR+p5NB3tIUamTqpDmh+cw8awF4FbB8NoGDbveneGMkiyh6TNz
ZJOK2nLzotE+FO3uJ7uyN0Mkt9Tv4GAk+jA2dR86vL2mv6/VBmUCbx59DrxJUgn6
95D0ItngT75/gZhYSsZMsWnFlIlr1PIOF9Fkq3+keqm7yRJijCr+h5wmH3b8taCt
a9laMCtyJXwQgpsCEjdwXKB1/gnMVzZ3GjLgLMjPTCh3coj70I/+uDyBXGQ7DQo7
a4rz5ELrkix5e2k/fa2xHaf8HumzXQ618IkWO7C2OXZWKzZhsd/eaFjznXkeqIXO
lgq5IRwf+gp+XZv7n2QTLIu9C9eI8ADZFQI1+x1KUnyVQqSigIHKq2cm7C/udUsj
s8KuJv0aYFTPpU4IB2fFI3CsnSUfnwg4Rq1c5aAgNw2/QzYsnHNjfqcujnuXzR9j
l9bHteNITNU+1AeGac4lfQKMTR6ucfazp0kzrxZcbMU3oVB1gomCiVbhjw1O9Ga4
sl++XHLS7bJwSEZAZPU3ldE5vMd81sPzHQYKIJd9rKu66ZDjYiPKBVnYoFs6cAL5
9kYXJLzKYk8IEhEBM/NEO6bFRGlIYuv8chsy+yP5rTD9xo+uj7mzNuEU04E56zlS
pLdy5y7mlVALRx03M02/gApG9G3OnBVZTJC/eLBc92lRNxocX8YEZ4THU0Gg0Y4r
wgWIE+UQVpcQGKZEYoRDtk5/Qw3rQUtVCunQdDh6bs3Afjn9CuceIHGttb2zBlZj
hJJ3CH/3wraQKqqNBHnWyP0rDioOi+7sWn3MYa6gbg4I3BId+gUehLx3XttilwEu
9yp9yDZLebltZimQXeBlPMqBRYFC1R+gR7kuVjtrhIw4oOoR4s5aeUQFJR8Y9mel
ZfJ57QchGrHMNq/mcPkx9q6PzMYmzmxewCwXwooHfDWU7DWQE+NwlFK/wgOmUC3H
1wZTRody9vDAcaMclYUh1ZvjDgzywT2kd0PrmjfnmxLatEATYkPqkRBNBgOkv4pK
ABZMAWUOVTYB35mxblVP09uqVTjKaw4JO0il4KFTtOmy4VKk8C8AkO3n7DwxlOMx
Pc6WHbMOleorEAT4DM/w541jrK1RC8f57nKejmzYnw3nKKhV+SEfAbHUQfBOvG/E
j78JDM7ZEKFoI5sKpdKvqU4e+4YUljTd4O8pUF8SuVCs9aR9MnA4KYhgI8emBHUu
QivJ19suJhj8FRfmEwsgu0izUHqkaqW9UwSdnthdX6H/Zd7r9j3jjzmaUptxCFs1
gefN5tjBpBUeZoV+2kaACjB0cTYGcDm2J33zTeIKbLUYq4SEHkmjTBgbQHbS4YIk
gc4RXOSF3hqH8upS1JqNekL6zHIRg82n8u6TWb7jgx2bXTOjUMgkuoI1WO+f+E19
QS/wRvVOJaPDkljD5L+oqWVZk0CNNnaedr/8/VrLRNd/kZJEmGEClD7dKbCkWb9Z
757o8u6aXCNsg5bxL4INrJMgKPIxg2Ok2QWEbfidgGFN4fOSvqEl1lwxWbToj5L/
v5jcKXvHOSOM9NNJ7ljB68geScLEpljzo19JLJfjxqhNIzhe4OBBHvvczUN2S/4g
aCT0yPAeZqP30JC+kvZDAyPPgw/V59tem7QmrsSer7jCHnMhDfT86s6hxQfQ0WyP
PIqwyPdaSuXQTK8L6p5bNvXRVNuZpB5ir7+6AXFGond3PvYHrEWLOOshMbLWRfZB
bLD5f3FIen6gc6lUBU11k0UdtRcUGDwblIWTARXs6FDr0DlN2ZXOvC2wpYnWkVng
TL6dQ2agZ2Prqzx6n7iXdUW8qVqO1P8fj6sp7KtFM4fpIGQZ6KpSpvW6Ct5y6M/U
giP6sfokwpOR87hQe3TLILiK9WGGEAMJfzN0GpocmcArBKB2V47sVa76cGWzEb6v
kow27hM8nkgrSlEJFgWH1wl0lZljJb3OUIzPwZRF0fQmOkwlpoe7D6TIRp4IDtg1
hwF5zdVkOTc4lM2Iga2ovmIoRgt3GSNKkLN7Ur2G+ogTSLsn/y2e4tK+GTbo7AVq
xiMbU6U5mJf06udOOUkHJ5+BFGzWsyKdJMNgy6lrwV0SRfLBnjbNIBCAQv3zyRJy
gXUym8pcrlKjNXXscEjRNx6FGuvxOXMK9gEdvHWc8ybuO9kT3Gas+mKXz2SYhxCB
4VGc+sKPcQAit6HGJDWNqn42wJSPBaOoRUhtGUITqhFtEteyJrjULUxvb+Mv7CbI
hUXKPZYigxJgfJxakZOakvbipkvros+txSUFPJldJEl41xeGeNqTWu6m0dkj7D76
Zwysu+Yo/rIEfbSNJap8cI/hQrPSuuxEbCOQV+uM1DNIyn641OEhx2FoGecTOcED
72rqwiePUBoGiSqsoATQTgYXW8T65jGUicxDAL6RNkYY7WtuvScRISXu14gqu3Sc
FY37iSVatXO7vLG+xqRCMAFTJs7Mx93YYHTsnnOHvsFuBwmgcNPHlpyanY0jSu9e
06zLU/eB2W36KCVX2yRJtAoCxliVxhbSG9hpax3k9zLnIwoFGTFExW9kLURYDdxm
vRjbMvA44siZmtGjqG7uBMvJ2DVDF1U7L9pYrAabOQhx36Szk8h0DRqOmTBeDqxs
ADcq3piViZ1cxSsLDAeY+eRDF93UPyfk8MrN5z9CfHIw/NtZUXbs4Kq9WhKroO1/
kOXIxEFNQooMPQ+sh7CiCWr4pGYN/XfWVPxpaDS+QVPYvzzyVtAkSTOjrieCCwLc
eA5gi4xGEkovszSXzut3ftuLMF2NltfJMZ9YvhLu868Uj7aoUYDziXf6sRil4uUw
qJwUpyRu8nIlSmVbwFA50gfwavL85SKbzOJ9ygQRgNl0uR7uOjM8287X8F86bMlv
/4jDZ5rVdlqR57PAgZzf3aB1icjP+kR0m7DSvYktiy1OFNaQQqMQmJkZEJ5RwC9L
di5MO43sVdlXP83CWeWles0G2Z3LJXKtWKmu+88cdqqUQsZKhS/LTG2Bt7YEHBwd
X84O/AonmajL21yCbHl66JIRZ6OXtE3XtnsWwoht35hlm08v0aiAmp97wd8X1S2x
AD8iSAuW678E1/KwMbt3pjgcr/NjNsSH4sVZjqGRvxB+oneHEhzWXMuBQMwsU8sx
11FaWHDpqBFC+9+uPToN5ODwuA9KDA/0TYVgp5qFLJS1efjLkUvCBcuXLKJ95+rC
ys9shsT8UTLhn/LJ05cj45TuHI+2pwio2/6VBg8Lt7igBrtdg5nv2RKmnX6jagJb
M2vDel5qairse7yKsrR6ZymSXjCei3a+G2KolMlHx8mOUuFKD9GzN6A+oVyxCrgy
bmOo/X2EI2D1kVxNfwwqSigJKE89IMucgjZ/i2NJtYwn/ODWUNxrgte9DCflVxEI
VX4bbDMZeua9ASn5zZfQyg46RcZqOI8mvxBhfOzo3gThf0eF2/E1Whm+p4u2AHd7
iVTEjIr0Ar6km0Duc7P7xEcvZJjgnEGGJr6N06c4dMc1NtSm9q5HdJdsRblZCG71
Tr0+/DyIEzwZXAxOxfRpKWFUmXuYnUmlQyz/ULsZAc9iSot67WjnvpLyMPNLB2NE
mf3MaZtPD2Kypt1tqEDlINVSmsonTZWkwCXdfe6rLhvUVWvrxere65kZ3UJse73N
MZi2/Aa05DA/3Y6cCrqTaYoLhFIfg+WAPDgZl+GL9DurI+rpKR5OvSL3qWhhjUgo
XLttgQlnanrsMp8m6sqhdWe8rEDurz3xOp5AxyCe1tvm/gk6AHYbgAKiD5im071I
g69eW+7GlchzCl2Rjjd7tiTXUzGPtczVaJKQSn27q1JcJJxuGwRN77A5jDxwYkJ1
1EstDjGT7+6lMY/HkxGS5Ah3ipKDwx38wXZEMNE4bAnXOMNJ1/zKGHCcLiF4cyBS
Av9S1A15MPBuh5UP8YtLopFrAKOEkh70g4F5RhUEcS8Hw0qxHwd31YPGG2UnbfFl
SPLKH7EVr2F3Ii3HSyS0ImeAHzrxCsEQaWhZ39LbyIQXqGGRW9MFFTjue66wUxrn
3db3291jrjMYyMcftL6XMuNAQ0J7CR3bxKZDspEQwhs1BQg2DV0E8LY9ubyeTkoH
9Hkyw2ubMDiSARSnWjlofEy93IknxD4scoPlXymQKIPZ2qsbG4vSsY5ozQM18K2w
nYXghSqjMWiQl6/47+gI8fbgwh3nn5Ue9NTou5QBGg3JTNSg48EjvbQ6v4uOpnc6
fxrSlA3+4msQnWE8iBVlfSB5/whi5UYtc/5XP9mTt1popLg+YpIvfBIWaH9pk95K
VNzf57QHezEmlTr6Jars/U+T7WIrHN4Z+xJ2sHpyHf0AMq23KhKM5LxNyOUkC0oA
/d4Grgvt2W/d2m+sVtG/ayv/fTxEX/+S/GOX56fbrfL2o9yZMnCB9zy0kfKBDARh
rrM5gyx/OVfvlmJyOuD0nQjoX2Bmbvkrw8IWLtf1X5HbCTRHx7sK7hDBZHzwWugC
IerLBE/zUy9AR19lbW8uSOfl6ne4naXndD3IQREAJ4kZh/uuoZdotu7foHzpV8TU
q6Lpk6vNLWJOUfVtnNLPL9P6YG8XrTQAuXeE87UDToIKPeK7MFRHPJ4cqAbkAPRk
hBpYRLryufpNmK5Z/RQIjp2MKSf6VtWaHtU4OEjHdd5fdkJbxmsM6j7PgQ8pWphc
sw46sVJpXy1qBhfG4fVJLUPXD+sAUN9F41QpDv1fIZ6VTJ3Tx/5u+fuzCqDYiq5K
WCaBYtIHYVOJRMEHOn0uUaTck0hGj4c7r7m6+22Io8EMIQFnzmBMSUWPxdbkbWkX
1vKdUL1IsqmVgMJYIiFWTD7kWcc16Jm4j/ivGZUgG5D9zT2utkAYtVPTCFWL7RAz
Np1vfqcnsV9z17xb9p00oMyXC/0Jaw7Uzq8gkAuPl1z2vomvSm65P+A/l+tFINiY
W1aFBRduBtaXMliRuSapfWn3/BXqDsti5BL8YK87t/DaTgg6nlNm/bEPH5RcPb6I
W5rPwjdUgowmTuYuHShpPZxw7NFjCCOeO3+owisKl5Im3aDTxlijiCeGhRGluoQM
55C5PVKXcdXJl/+tS6rZQeKP6puc/h+HciyQEuDUHDCtEIN9+cFUl/Gm4fFAhn1V
IA9vALthp8VSYWZrzT/WMMLddIkYIPVgzcYvfQbDuqYNTfE4IEj/E3xLqUf3qQuo
lpqEyOA0nL2KZ4SHJyxvSsN5C7TV5ijYy8Ok/qKchd4Zd2lrzxQZlfbomyFlSVFm
msJsNssBJL3Q7hrJfQaSqJhjdbx+Z0drOXeht2CVvmkEAGwD4+Cc9p0esfkUFjVl
yqprUTF9W4f+Va8mJwfVDHcj62SWiCxG3Vm85tA8fuCIA4BZYyTZnjrPGSCDSZnH
o3uWZLVGWpYpA7ZEfGXEpXSgQmuYCaPhkwZUGoV3JqCCE8SrOOeCzTxlj7duRlfL
IYZrKttbZiw1C5RCSf6TnNr9OB0yD87Q1MpbHIaqoOthLveaLs/HdPtdXhixUC+G
Of1GWeprASxJUhK6b6YXggH856xilanw85oqZkrkHJG5FzTye+FgMfnkP6sxbhhg
10KhpYFWDd0EzYkOooKa6CHBhpcxd2KrRgtX6U/tQAkdNkfmKuIElXGIxkmjbzDi
1Ccu3aqlR+zMKguvUx2V5oZ4sjK9Ukku9JiogpC2tXJsL5+HF88Ao9GBF72tlsB/
kknXwk+YxfXgQqhlnnbG8LK+kGAJLcG2OBlO2UKMFFWXjUHx3gP7DkB1E0lkyG0F
WaxLqfDxrIsMlgNjc69bYdSr8UGovPKrTDIS5/Qp91sLlfd51f1NJWuLmQWdRVDL
FElNF+rgxoEg9ugvKQT6dR9pBOjYZC/Q4fmLKllqNKIIz8QOZ/CbnlY/mYB62Jbv
57oDR915ynG3X0OZCHb5Ye6YcFW+XRnQl655mWsd0LfpJeYP8bVmDPZTRLwgwn12
uoyMiFhUgfWVLOPhcuf8x5HiOXr9aU03RLdKow3wUbveaud9JcFZRIGYqNkUXPn+
oahbSe7LdTyzyf3Tvs5+zmh0UD3v/e6iVvvNLfVo25RzdjTDAMupqP/WZyaXb2kJ
pQxxPxqU+dU89mBZ9AR/W01S2BB8fkbGw8TgIE539xPRGBEao/XI0muvModqjD91
Lylj5YNgcAKjQmwO3uORmGAw8QoAS8uihkS9s6KgabhrXYBvJbd4Lk2vyWuDew/O
J1D6waTTZHi3tJzM4T69T5PZiF/kjEfpuxEnJVXw1ILKpUYdOY99x3J5qXLM3XEX
C5Plxxvtz1i0AVvRpgw/weo4VVQkRPU+vOstdrRCB/tTCXrTcvu5BKtOV99PzsN8
NkcbTnV1TlTMXZ+PgC/RvRBzIijpDAoLOS4iswCBIHppkkV/IZUyJKu5MrPuYlP4
Uz6DkNGUdbHvC8Bbo7np4iAMFnWcJZKOES2Iii08NBRDIqAbdHVgkNTOM8Xx37zB
RczvNCFE6S2QrbeQMHp6SCUHiiJpP4GcG71xGq1IsuQNNqVssqR6O9LOkXduuuby
rbyaXy14dPkNkPQ8BUbJb5CRt5iP85vuCAZRROW39OS/Te+H4wQDzqhfpijsa9nV
xNgqlB0iWm87DzHFh5cRMSfZY9gLPpBQ+BNJMhrwupE7VxdUAplzjGQjDsDdTSGL
T6QLsQXMAJFOyXbOkkUjB+eySm1Z35NHmFcTFw2VisEeBhEbGHZ6c3vm//9yYf1U
LlHSrHMwxAXfySpCcUTTq6FUCyYkHJWTchKJMWE+Hs37xo0nBPAJfCouZh8GtC3h
MDt5b5c6h+3k26TP+qUQfubE/5y2cFfgDPYUlPXgIuHeAVp57asXsf3pwJnP0z/n
NRS7UC7u1nDgUEI06shUuEUBZBYHw3SZPcvEvSoGuQj7qrW4SsQnXtMKS2oHff/D
fQ51Sx7b8lERNTgtxZfEZyZ9H2c8R6DB9SxKXbxnoNlDCmVWmNk4bItlxPwBwaJS
uyYoEdlHj1E6j2yWKt2g/N2C1E1nyiZqWUhErBD2KEjk9Hi/KxQFAjRaDPGDoKkF
XOSZx6jfaO9FlzQmUG2rWIPYxyeIq//iCYdtrxAmvf8a2kq/0V/6tEXZMxDKHHA2
U9OY6YqaM9avQCdQwMbyf22YGoQQX6ltmsRt5oTZpFmptOnVWxRHAJU69dX3LHW4
icejkmCcZtaOr5o8ExUJ9/xWRUvrYlbBvXOAl70SUCr0qfW+K7BAOzrF+jLvlcBy
GsVhZsbwOBadSvn6f1mNmJDqDepGgHWhceemA0tmY58R/9+HkdFCFisgcl8OKsBb
ZlLDnova5TtfMt6lbu9rtBIhIt019cHz2ZfSmQtnxtg10j+yYBxZRRI1dJBgCsPG
Mt3oC+8JurNaW7DPYbPfwQXxd03CdIxCdwSLN3U6xFC/L/eSl/Vm1RQuhwubO6mz
VGXMK305JuGPIwSFvRuygSRB3teDNY1CUzFsojUMXvAzHW2dWb6EHiqGcDcpTsoi
YrQpOF7DOuSvzQjpv8wdHHlxImevTRDrIDP9gEbjTLYmP579TpI9A9Tkwldn8Fx2
zzFkd2GUfL/wbD4cn4aucYAX+1YN+qj98m9PczCMlL6w+pBJ3/Tvd+E6eObFl9ab
cFafOKfOv62qZ/JQtfcyf3d/3UA/21LuqMuemyqZnXm4jSAckzjpCFDzN6GxzKXE
g9xwL9vv+YsETgaAG77MReJnYZv9K+OBtEtPCDuTX4AEfPms+/kNUeWjjg99ZvOS
k6DQ1FbFYdL4CdJkQCVIDO7CM3av3moBYNPCqVOVsZSrpYlC/gns0B/w3YB9axLT
o51ahi+yGRvDz6bUzcRaaf6c2vMhlTX3zo3+09AI5Obd3nSfQK8SgdCnvQWyLTO5
bWLbfVMUbIqyLpryDdeqM/sQxoajVGQ1mwndBMebgHIxnW4MPg6vbhBIcWb04E89
VJ/o37tXlAvak3EupeoAtSc8W6XKDGHEz+fTiAE9sskgqXrfdutEH8YKatqq3+eP
fotBo1RoMTeyNtbmKNVack7ZhzuF4BEuvA6QYo2hzmEMmu1O0HEAx1Sor47nGOlS
tX2UO52c8cywkSiMWTTqyflWQGxBbz/WK7szyvICTxufq3e0eqMT5nL98aW2n2iw
hdhG/w1vbT/055tg0ZrJ/IzDusPnJYAmaMfXxkl/EXUnp0whgYk7pgVgjoQcjCfL
ILMP/KMMBdqu4qXmRSi2bd3iuK7goQ2o7EP3hWX/hdizNPtPLUGVWv5QUzNQHBbF
wMxM3/5tAK2zVHX6EpODwYOi0xPVEaOzbV+gy7h7McV5RnmHSRHCavsXUnfPAApy
CrnxVd9PTaOckyprJHh9BJZe0g7sE59e70kBKz7IY/eUkvKC7kvxJnWfYWpA/j0w
O2kzxpk7gszui2yfyUhKhiW4o0gk3DgpgCNkS6nk9TIwJrkR2WXedu3jtZumGi43
80z/I2WywbvLwc+44Lds5dHNfX+LLwB1yr5o4zoVN00GQpR62qWxDjoAMxv9esBY
uFAFtodvAkCGC0QN3AbXMlQ0HrsryTxGIt/sOqlg30PYGzGa81leEtJUjDz80xRK
ZyJWshqlGtYL6BJ5PEs3d9HODwdwBFSfWts7jsK8x703cvrwKQV1Jc8DaVWGWIx4
/2SyBoTtH9hPtu0pAwsapTNlKTmY9lrvaYL/5qQDLIdz6TdzCiWOC+QQL1ELvNCR
FQSWyGiN4pQQbBhyQ5zNudA/4bowZepsD3SdmBMf7IuLDLi7BOWK9YuMds/u7FVD
nH3qqgXCR1nt6Yv7SNf5iIkwQ4Gz35hbU0b+37lbTi7u7TfRgOvg+S2El2Z2dqj5
SEUELQnzh7nWUKBtfmOPk82gToCXlQlPLdBcRXT2GwYa5MWpAweJNzoSvy4wTlum
1PMyxCQxI5To76D8UgOcRpsir+HXyr1vVWQvav4cihc2srtTCLQHSTOiQOMqUyEd
iSIdxiHkkHthi+cqTT8kyAAXQuz6mklJAYa3dZ30El1GUAFoMk58L0WwlEZptGBW
qxXu6vZlnO4OftyUOYQ+WJkPl9rbf2efsuh85vC0vv/sdWGTzzCrQP3QKhvbelxH
V07yIVXBpNQzl9ELtNN1uB6FCD5CcPcVoExn+bD5lb8ihZjCljTOX/LT2xC4c8BT
i+fGnJSKuG4qlhtqCaknBCAfxjojWoq0rzc0BbEcG4qsAlghpqNK13yuv6F+iPHM
2Zqo4CfNJA6qHH7CnDn4WyeUYZ5eiGGOEn0HyH+HXHu7yLS4kXrEQcHg8qGQyCxX
WysnN1nw83f2WDJN9sfwfhCwOtV3J3gSDcNg5dW7AW1AQzgpi/HsWcuX55ytrQBm
xjyLV2JsVz7FxtTBM7GGF3dTkbk6GWXKaXH7Hu2QDvehu/ksJDeg8IeQkZZLtxzD
LzMUgF2NpQ8eVXmcrZdOrkY18K9H077SRbmP5T4l+6a8wGbyQmZ2Hr5tyCEZyEvp
zkqRWIdPdg9IcS4j8CPbzxo7kb67NuJxTY2VFP2aveQJH7HKIqwkNp1ddveeB6Tp
kH4OavPsUsngt5y52khAPfsMKYmD5EnHVVMk+WMwaMdaQcQXxsZIfbe7l2zSDMjR
WQ5sFlgazQx6Sc593DXvlhDtY+MK/0tj7Ik4v2/RYGtdoterXMz1Duv6cAU1Kd5w
3CYL6INXGU+N8MTCRfwhK1ts9Kd6xysgHRdsTnH2XEoFxPk/1kbNk+DJTa6dH3OS
x+6Ixcfvr8axwGPTu64U0BoT4hdAj+JbS7OAf4g7UNCX2Iu4j6x0rIE8n7I4VU2o
tjw5f+TTfkh2zpM9LxlVwC7gU/zG43UE1mjosJZK/xQ5ONJ/obHfpzJjKlho9WY6
bUzrMc6N3X58Fj1RofMowduKpgJgVO388UgJ2L2auo7nI1yjVSuLToGT1ZhWlnyR
WxeRp5LtUubJxBLdY7yKYR5qHsDN7sGXMNt47SoVc1WFawO1hRZSrYWR62d6oc13
HX3g65ptBK3NmXHZKPlTWljF+lsIJvXc49NnDn+/NL1Lnk0tZQ7VgtujQoeEA6bp
CXOgPWBLFr1xBWD42FaGYt4BoPLFnFrN2B9o3MnhuF7flMJ7b1B3uIEp4kyeipdt
BoalxAR89hjOpbqnEh5MhcDS47nGIxp1czAasiZz/o68eX+O6UjBkk3pgcHxZC3M
osZU1mTSYhp7/WUVj9vJwQsJqmHNi4E9t2eIoMpG82tPTTRkJOC7U6uAVvCoXVqJ
UWbRePOiTlzd2/+Atk+7Kn7ZA17YqVz14hxnRxPcxTfZQ5oODlE0C2VdODLAYmQ0
oecdK2WwCCkwT2HssCey3V0XyPIu0jWW2GwdAflatoESIf3sisqq3IDsk/pz5iMV
pfWNPmwAblxEW/gvp3jI+xai8MxQepF20cCfJu1IOhnWFrW+oJ/MJbhv/KMDMh6m
ejG7ihVGp6VfoLcTqPV1Ihw9lkGxw8ujWOidn2DaYHsD1XyehbNC6XXOd6ZI7ICC
gtOPyPULNAQfPzJmJLPufSkGOc3gIW1A3J6Rx9sWK27P66qcf/s6ZEshDpbYsqN1
XBF3zPczThtiQOj49ui4gpzqSFR10dAYuOfmM0hbwTBYVL9P+cFQYx0vwnU5Ta+2
P+0qy55GRkHOkwADQnaPowCL5cgTD9BF5V7sfNJG4UItYnuVE4kdbisCtcA6+evZ
qszEyYwOyY53O+KhJPphJX2m+v01wmYOStrNPn//MkKJRboSTPLX/xobRd4W2PF7
N6NVpOmBUXDUr6kb3M0Jtkzb33MTTad9reiNYziHG/L8j3yrh6UhO0nOePmyXGAO
Shbr7dZproi1wrlipXHxmOyxji5nD4G55Qb3FrCKxX3uBf0QNEN6C24JqKdTah0l
ERuRdt7M2rFDvZSDRsbpyv/JxgkRg9xO2q2VRAcjlPWCYOGomCOyAMPP9xUlq2IW
m7tkKysDM2CMdWKaGnqg9vEXxC7jA96nDjXD3KSvrT8O+uooMI4THvUhF1+xTEQZ
SJCVFFAsrEqkrEupHtJVJGqWo41xzO1UQRVu32ilstprpv3KtxpoiHU8AvCFTEyZ
tvjfmu+pmLNgL0dX6UjJm2E1UTdzpWAItejMhWp/gN+vxwYcnteI8J6d8JxX56lC
fnTw72L4vb2W+WmfEJH4U2KjJYwAhN0KjPuBgrEiX9hQPy7pheL+V4KtwR272XBK
sKt4JUlXLwM2qzSxJ/PdAZsPFbWFLU/WJWejM4GJwVHLYd+483oc/FV1j2fyFK8F
+GVj+iCVIzxn9f26H24ed7iVgMAvMlJul4J81P790IqSD5X6H0inO807PXIFpbfW
eIAuq2+vpVyxOBkCerLpN9H8fNLBOp6hemKxori3krRsEOjM/W07zFCn3JFvTsZy
P4NlH3ceQ4NlN9jcAfWPH6IKL5HOGduUMLlmkaLEVwQm/jPby/gEZRVr3YtopTsG
Zb+vOTLgxT7B7pKSJSPwGSy7hXoD2qx0/dPztwiR2f4aLEafOMglHU24BEaK4a3x
2sYMx6nYHNFrIlBgoacD6gIPdxiZNmUVX9xh9qNrkMOY7t/J4k9Y9n4ol6GIKu0d
hzSGU0qNdCdz3P40l4m3jbjLH/ltlBNU4MvulvT2msEM8DdCzbNoTr6GC7WkpN0T
J8naRqEORiS6H2UxcQu+H505cab43psEKSPrI2U8W0varIgJknV0FTfIQu76tK6/
gfjJqbBUIJYTX8j0fKBndz2oDoG4vSGlMXax4fWyeJI2bVi59sotFkYW8qjICUzb
s8IztySxiKqToPY+zFYAaHHtWCqtQ2nHwAvLySLg8unRV23HBt1QqlMwldnD+X81
vkMz07BwOIf2bpkrZjZN+QgZJoxRZufqi4xFw8tda6/qxhwtO9ml5ywDNTl+SBCw
UNoX9a28W1x+L3Gn8FhV4kVUDxVUou7a+zC3aw5booGs0UhWsW+FozU1YSmnGIXP
uJw0sdJszzkzpdBj8Yhg07/BE2s6F0o4OudYrrtP0liBEKt0Km3Mg0LJl/c5Pr1z
SOX0Ae4mMBzWmwX0zZnW9byYUoQunGR7SFUC9G05M4RuhGkbbiJenSmBSBsZ5sdz
u+vOae531XQsyzr3Aj3BR6lGzPThnbOCVE3IkOVVHabY7GYsV0HqeXlL5TkRjkeM
+xjRxhRqQXcAIOWpXYrnXguCwgCnVuSnkmqMjFML++POV2EuQP5UivWPcaepoIar
SEwX/gOmtPQPrk5ni/NMQQI1QCISe0PUjkP2/xT7P8HvbywrDt/CmbNJ3jWsUfyW
MC5vMhuxt0g5YeZevp8YeR19xnNrtj3GD/eJgzwHZ49Jmax891qJ21mxVY7gwDKS
pW7YT4ZFqw3kZZLM18IKGZnd79Odg0Fyg57haWBE5/cqEhKaE8vNI05B1cpnrW7O
W7o3V3JpdCgyNEJto6flamZjYGVUC54yaesC0f6QKJfCDYH6UTxMdaiUJ2UQUwog
lMC4iDX9lkC9233JjdtMncHhYdU+laNQGRdAASGKwz8lsqHw5Hen9XQaJWCU05h8
7xzp0x3G6cJtytwzoI5bLKQ/czJSXRDvV8CElXxP6iKXm9jHUf6tf8ZBczWbxhOB
nGsA2iL3Nxpaq2jYal7tDgjiYHCjXuWFWNwP/CSDY6DSjbdeRWVw+WbAdVccufsZ
hTZjQuDqPXJ3j12QVCvSynY1NMvW31cr/Nu17IVBHtXPvZYAdznwE0TQnTDqp7L9
7h/nMx/PHRlhRcI7lbAF48C/LPhd76pWjRA2VPerjP140UcrsabXsxys2ADKL9PS
CKSL7RqWCR+NA6CHWbZltONysJ0ThCMpnN+kdf+eTSUzfMEmrk2GijN/cgE0gJNv
RJWjzlwBWHNA04IMW/dw02jTJLNTw7ytoFDhX1Q4ZIl6BpJcndcwMIo4QvFLMiG8
suN9wonoGhFf2g8/7Z9wu/O6lMGZ+WpY4oYJEcU6gts0ePqUChPHtG2bXSwa6ZHT
t/lyxXAsgDNfF0WaFHpmDK5LI4bl5EkT3kI6g2c+HFeYkOIC4ymTqpv9o0Jf4eEe
9kPml6g/W1mib1uVCDedu184S6PyREouGsbqENj/vbCIT/eJ2lOJfDNswcIMfB0I
W+grqFKdqxWyPzhIdkNVlq7cqPesZZCrKMF77qiVyX64PJMZynAKQgio0asl2S5l
m44wa1I1ETf6Dlo0JUuSq2TmNwPAC29J1alFfHFR8RsqzH3+fcdOF96WELa3dDyt
M706s1PvPLDoF78EylB0dMwr4Ct/Ml4Ku3lP1W6iRYcr041JPZDQ6l9UwqKhIT+s
WfuJKl2u2erRpI8iLCqLO2o1bAsxU6WF7rF6xB4joikyTkJNV9Ka8D7BbwoGC8Hi
bfve+Zyvz8iXf+abaQsDERxIU6ZsNjcyScwjQnOe+nSsJEmXGxkCdtBuI7PMfQDn
M+eMG81xoJknsHiVsxs0N22k5s11u3kOG9uLhI1p9lYC/9fvic4KQ5SKZc63rygc
YGyjtMgY33F91GHqp4oXb7JjbZhiiJFa0KGT8llkyf/J9pVAJxt4lZyrMjXHQnXg
qhUtRzL61T+YLo0vUx7mCDifcwJfUCMiYkJmf+3NDeryNtpoBtwARP52Pd7Yc6mw
MrBnQDthHIcTEBD5PrDiQ7OQ/1IIUQlMZNgXPAP1VIr0r4V4/PFfAi4XUAOgwu9R
YatbRGPRJAmB4Cuw0wDoU3A2Ex2lJD523APGd1WDgXuKrRLGagy7jnglUUyjbc4W
CHIkbad3/YUxJnpCvQ3IVtKV2x/ICE0u4Xw1okAy6Obp9vENPFLRAhdxIjIP6uNq
W17pBrSvhCg6NnvKBUKbSnyqRlLmDITZTjBjtD2RA/SPq98IOj4wqcioVGfXWd9x
ixGgugXDKKBdDySzC0fNwmLywtRa0jy97SmCEzzJgpiz7CeUkd83Qh0ro9FixFrZ
9vchj7r10R4H030FxkeMiym0GDMZG5X3WqUv5E92JjxV0PPECZ1/jf8Ib+N58rRe
eEmPCK9Cv5lRLbPusAs9jMup7fCV6r5FhAsoJc3hfIf+3xZgESL8CHXCNxtNSZ4m
hPWv3wcZcrYqbs35qK257X1HkAUZ7b/lQSS5O6KbiCDLUgkbxKeQf+StLayNtcDO
SWzc0ocOxocAk5HPzpemF3XBHXBlSoLDVAenlcon3bXiLbaA17J9q1hDXrCjctRL
OjSy2sB2oskjUQRPwasMFev6ZAwaRoUo2Lsab7ZGuoJD7JhHeoTDH3qp5RUa4rWE
H3MvM+ADqt/l02wQgQRhdJo4lLBZNFGKWfQRepv6YoY1QNqmfbZEbwr0FyxeKY83
DTP1KXu0fiTsAaYWMD7cq/DU2KpDVVTmESAM0FM3f1iy7xJT6GNnfkyx3YLNRI6A
DFwUhJKcx3Wrppd0Yf6yqMlgJH3KBbj4QwN2gYIOtgnTRQnRqlNjipZCEZ9ogg3t
YcX4nd+7vDUhqHyEqO5QECPtUJKoAMK3/qyKgSJU+JhzWwsKIm39CosRlELLpwBF
KbFpBLiOoijmd0yQr7AqUd3WebkgzgaoLX1EfCjyHqQra2qxhit6QK6U66tCeOW4
loIx85Wr2jyrg3G408I0Xtzuu71brcNyVe5s11SgIWysLp0S77/qfTf3/oqNYQmw
/1E9N52dL7iMSBP1UtNN5oCS5IESb+q3/9VxlmJLv7uLl+6bERtX7gDvuz037O/t
hbE9i1gEjCZTwSw+NIl40R64yJlLQ2jXWPDqGFzKoenR+NKgdbWu+JXHFAiIc/zk
DrqCD/yda2LN/IQEPpEK5me0X9gUp0dUJgh5DhBDxUAjpS3cqh7jkAPUmbqFjLTa
278cyRV5JlOJ4MBhiFQ6QXsFEm5gtjD/wOIdd6ZiSs5XFasx9oZ22w0kJr4yinwd
TivWnmcFsrPTsKLsCLtpWo3CzsjVlzos88EaMtWSQBN4HbUcVEIvz3ftNgl+a2H2
83IMNTOzJjiJWU7eBozESiAKe6b99w4iLMPf/TIU1+iAMdJfdMJCJGQmohOu2C4B
uoeKcvD6H84z6CLhowfh+Gccm4wTF/94imQsq35hwo0z0aGcwo78NO93R2b8bZVo
VTZSvX2yxQNqEZJruzoQ8phhXvCeP93QLU1v9CJ9Xb0JDStKChsZ10YQwh9B9de5
1h08zwxY1mnueJXd2DDUJZa/En64/0Ap9iohq6d1GTAULi17QRz+ZnVvBIZMvEf9
pKxsiy4LETReWFK4jlTZ3743gbmSgpmjSHuSBgxZmCT/DAj5Lu1B6wAeElFi9h4M
j+xkh/F2Vm/8KEmn73tkZ7vJp3+85Z6jMcBalkP0KSNO4uos8u3JCc1IVHxRvUW0
dbRZn/Z8kAyDz1M5gZntKNXZ5Kw6Q2psuiUOmAwOOQxK7iYoX1HzaXYn8Iw1bmxb
+NXKe16PDFi9RGhHxe9worHDNfDQhnk3tkMXtNbbf21ckuOySCWiDvbNGorrjamJ
fXyI9E1F3jVnte3kLDKCq4XWFwdXUi6xFAllf8fCc9Y2+2MUn6QFjSbtRqEhS8Fr
SyUv7SWVRpzvNN4YFsCEz7F/qqSjr0N45WHbmyfwWYFIOmIWkRbglIMlPEOZmafs
H/+/ZH1cqsShclwG4MRk6bWAHi7lhWmYWaklym+5zxwgMn1sZJN/zsZHM0dZxUJk
4tWcCAqIIDPrcqYTZZJoCJhILZIRrNzls4VerR0fi6KGCtdM/lUWppVoYi17rrwY
hp/LqBCykcvIsiYgQeDStVhxAFEIZnO0mqvPd7ebwhXIt0mKl3Tyqp0k0oqaoi5C
vHieHlCUU8Fdtbx8i4K7WQThZjTimjgKfNMks+nbulrvGH+V3iIRszI9F1/IOiEu
erWdoBnnQh49Fzm4nFeQnGa24jpTiJxuAERMNgzUbRxDnsleGvU29O+zgxhZYrDu
DZig6grutLoC15MlPgsV2BlmXMWvDqTuiGTcR5x92ZVcRo5Kz6CtdZWu49oVYH+M
FYGrLBMUz0RNyrIp82Rnzh38J84seS9AsxSfNdJsLbTxf5vKtTiEkFzfcjEswZXh
sYIkNi3O/++nFzX5KYh/vHwykyhGD5VlStL34wfQK3d3B7Z7QCJlS/E60B4GiB97
qlCk4tgsdg3XAKF3MrK80WjHKqvE1akrv7XjSdtF8Z5SNqi1yk0uqjEQVS473k0K
j0gyTM8mFRF1TJN53NG25RNTZsPju7MDJEZA5JvkXV0eQcaAK4CIh2dqT61ge3S3
JUS5D+hoMKJuGGb/hi8+btp4ecQ99BDqMGXgcYvcOZQDnOOEo9Ajq9ImjoeZwoE4
+JSar5s+AZP5YiRZH456tSElh8WCER+wdtNkV7Z3u0xHfjWM1d55/botfk8KMnIv
lPAZLCIA3hMPGTFAuD2nkGpD+dYL+HrJ3R+Mp6JtK9vdOa4f1vxpT86mqiECmD09
i47LsXu5s+7Z+a54q4k3We+EcxZ4cMBlVQ2eum8Eq+b/DQL5XrtG7bTTcDC8xmr0
/6Vu+iBqdWz7PCPV9Sqw7UFeOrKSyEoMOoX1D6fLFlkSJuosXt6xcBTNEP6+6bkp
uhUahGdcFf4QhWBiN4X5/Nycp6wuc7P/rmenO52umhtB5u8DTvNP+cFAxacxHRAk
iocqjTUGyvcpHxqvv8RX0z2AOenVRvSJtQgLzvVGjBoHPCJEpJppLpp5sNi6zNRH
xaDL3lPU+/FXZNFohpmNgd/wvT5o2ZKvm3iygCxV8w3UD5vKmazlFObvW6WqhyYM
/mbsZsYQpobK9YvcdME6dJZc122qCAg4gcGO+X/42mDOfxexxmzeo6kMTucSzVvM
xA8dYbFOQ5fQ6c+zy8hI3dxT4BRYW125s4Ycn1BF5Y5enT1lg9+GzBvdaKm4rxa6
UH6yH1DcaSd2HyPf9VizLJWfoO3gUpqKqRwZzkbuNunOp6DFnJQZ65Qj9g3gVbV7
RnvcQ8y7BXwMpcjK8RD6cKiG+lhYAQdSRgbbEcD4pnVjYWbT3300bDQ8KggVk9cq
J+3c1hZvOG53RHhSAqNYWRkzv1A+zKxTAYrPHg5w2k8XM2MZOQD7A5WSFIdUJhDU
fC5K8jiApk24fsSFDnF8UFYhr/tUdWTykQwPNdqVzTTBu+W1EDMSk416TZ1loQ0Y
5F1OZK/ToPp/J+LTdIBh0YyIrvnqk0MLqmD5yOJqyawE1mjoHmYQ5dXEupAaioox
DQy2AaNMWV8cYjXrUddpY0eo//609qgOhAsIYgqp+CakmD3Etv43wUSOB94eNqWq
loIjNtbojnoctv2ori2WODKopJzmNKWO81quN4g4mYyKskJiDQ/E9UkUTXLyE+Ot
XwNayMIo0Luv/7+LtixNbi3K6xAQNbI+s48ibI+YNRWstCcu/oDLNWAzNCwbFDK2
y45TZUucoXzKNOchX0WZKLEty5DEwyYQVk96FjLLppmLYuUROwkA055CeH8ayYU8
aTAUAgZohusak6LEc63XHnYWXLRhJ1eapqpu22iu88tsERuPYNEMT49FepZBURbE
99MeUo0wnltz2b7bft/+37uRIRJHdxF7U++RRGobQjRjfiDPxftyKMXnWPiMQ4+C
8Ph6R3bHQjlr5Xumynm2ktrjl2H1smRMcI3GiZJuOqLNI4cSBEjVdTTXsM1HKIak
7ic1uzmNO2Px1Sfhy0r6YlRSf8ZtkjzlbIVYY5HT73XgD/xS6685dsyk0cTLEzMP
/ZaY/aQkqKLiMIHMBXQRdh2Hrav6P67JDaKkKeE210f2TIo0NFp9P3YGIk63EKUL
9qs3Kt2X3v49XZ2QlatGWQYs/51wYlA7cTeTq1o+62SoqzJCd3+O2h5aFnJS331G
l61HJWIYq62R5HNnyGouJHx0spmD0eZkZsW+cjSR6fzjTzMDrRDQb2+zkHWJx1xz
S8H+tu/oiSmPngobw3+wa2twIOfnqNwqQmUHCLjt2OVHO+XRwCIvW43z4qoUcV4z
37m83LojOD9w7JmpeQvELeEoxlW3tX38aR0TlfpvlYq9pvvB56GFnZl/9Z5IC7Ok
b+gzQoHdQW3xfzRyIr/frahm6rKkqQjeeSycubGRGEUq4rzq1foMgDo0U8ZJfMaT
zcQJwmimk6kbCmXZ7WtETyx0m154C2vbGsyL+TNxaI5UhoekEXKulKYr5foCg+HQ
4jQmcd8PwWRd2mB8bPVBKKHtxRwdAOl/RzdpQ0eZWnjD6mD77ENcxdXB67p/Jmtb
aHcKAKU2/H8rkdf9ArRGUvvhYaesZmKxZLfkWwQciEcZzE3ndVyiC2dRzdy33FJG
XnbtS/lvtrFUcgKF72C3Kv48PYaoL5LkJPmiRIi86adWFaY3ZG24kqiy7ZaI1FO4
1kGlVoc6WkQ73V1qpFIwc2+brwfZZhvbeJN49Fu8rVyRarnrPuGZxKEZdFOvPBUB
D0Jp0XuT5WBHZ2tDY/LriuecN3J/3MWwfCPHpc3ndcQCSWQ8bTKOWNBrpFeYy8e0
BjfwTouhVnB9qhAbHexdpnY3f+JXyAx8kV403h205LGkMY5ug+FQH2KDFpoHKQEH
0dR4b+Rd9I++nW9J5iyNsd+xN8EE70NE6OVhPmVFGdCH8i4pqcMRupcHnBjpdvH4
UYWxPjZV5hzNFJpdJT1knc1SQQbayy4bIWtGwuQfoPjMfKRc2MNwtGCJlfQrRsw6
TAGnQeTy3YWOHUSW5hbqd97V/CALvOVKXl7COMA5jQzr8dssAmIuTtEgUpDI6EOz
nZPskEt4edrlmz6jyFl8TAnD9/JRPHgNAJK3acZeTGUCfPhDo0A3rekjoF+PIltj
g8fAVNnKY00KEIo5JHjESAY1clAWd4QCx+NFxRma7yRdLaOSDb9xGTONx2h4rysv
qeECsGAnrd2ciy94e6Ml/0Wh+/JAPVqMYyEeBRak1/bTNqoTPn+wZDL3uu722vXY
T8irnigm/YS0ktNF9LdiEm/Rzl570+rNT3LvW+5o8oSdJnE6qz/+HNO7Qyub0As2
kidgjBmeCP2+0ZxVuOzBmbYPWbJ5QD6GNDx+GUDiZ2FEwsU4fPFzx1t9Va+sp5Ly
+I8OTHf1x8+7ggk3y2abJtlZOLlld6R/LI5jbKyCEdWG/xBcqVMGEPqXhu7jgJ3/
SJcEgNKN87VeP6i5TXsqkeKJ9kchvaTf7SPLXOUv/dAac5q+i9PYjZSVNdN94Zk/
Go2Xmtzv+y2ZttaHuzU2ZOx4+PEouvVLuNReU/xV1ncINPyzNCAXXiu4YLEVUotK
RUpoYjsqBprJO3YYhwih9984rqmjkp3ZsRRbscNyDBawAfthqufHPeP6ljXIgHTE
cb5vUSV4L/MJtj3dpqzWRVrtdwD7FGBw0t3SNobthaOizJSeL0m6gJZBst7Ru0a0
bHJ7t6PEAUgM+1cn/PX8DWQKSur6DLavMgNDT3dZSykI5ttFm5Fv09douE31V83P
gYYtvnGYrrG3NialgO/rzkk7fTvduRBPzJEog6SgMQGALm5wULUIPGpfFvETouUp
efOBElPeuXUG2lO7EPuTa3CNZYoxx1zVSkBLf5plYlTwYtDpTZiFvwfjyGF52KZX
yiCwAxjdmB4DOwkL30y+TwF9R4Zu8WeoxLsKpvHX0hwwiIFuU4Z+4OhvAZs7zZp1
5QOW758EbEvNBig495gugp+rruKKV/2TJ8Qu92yv4rJ5nHJGQVoqP69EsbFgPYAk
LZDTsJuM2nW0QHz+F3XTvVlOA0HDYs3/DzL5H01UrMYDZWsZ6lFRrU/YmXSrgyCG
VwYxpElMd/jnjgy8gRTjPBP/49hImZhZ+Mdt3oP+82foAfXzW8dDbwWdx28tzSOc
thSfsaKN7E32efrrr/ZeJXYEt/9LaoDgD3luM7kMmLSa3sLMz4FDF09dTmM+KD9p
VmMehEUm9sD0nUwSOamVqjJkXPfTAZi9hJT2qz3J3b8A6oFxr7xsuww0psquYQPB
sp8dPnAgdH2zRU8ou2Rl5pApRmdGDfBQY4pfV+AKnExQAGoEbVIBloli3O7ueJTC
bwqzW/LhRi8opDwsoN1fgKdWumEM++jvP9/5WHMx3Z/coKtTD18F0lQ//bRxA2+h
/+qGU9/TEn48PWKJXI8mKGuYh/dwTk4wn3qQ4Ufv7fvLpuZ7Gj17m7sE5SuB+1Vb
6XCmmx95dDQ4NajH1RkyfIqJ1HuEiCCp2bs6RLP4Se+SuE2/7RAD2G52GcbVjSj0
ckCVaA54ti9zceLC4EKSTGehvkjPzvN4mQqBE5S7AfFtOSq9KwZ57oH7qXW0DK6x
TbXcYlQrQhOOEsVW0rpemFdY4b+X/zB5uFJceO5P9fVNGshhkCWqhSeLUGSZLwBR
0jz/D93y774qUX8Mpm5t4+LsuN6zXUK6vfWn7Tmmf3PkN0zTnaEj6szXSPfC+0jl
CIHgnXOQ6rQ0hgyS9djMSbif/xYOkQj//bxkXYz2Dw7wBpiXDur7Y/3Yi/pbXp2h
BTA8ilD6BM6TM4gOfVSzcep17Z756T3p5PqRxT+HIAsJjx72qIrXd+869rVJFFIr
0BaSwuOUV8fPE+1AGkurTi/r2YCYNVReayDhL+0jpyd3Zc6XL1RK7JymuStP+IQJ
3SrVEgER2RKy9VfRepYjCuwX5yMK2JUNeds2wjaU9bVr61r8za4uJ3i7ZMJbkQ1f
Z3qsqCVooHSR4jlynsmTnm+stEZZjyhlYLR2q3o/fsmHaxFGuwHKoF8gq/oVBAOM
b4UbeLpkm7KXhPpjdzjHa8z3e56N4TsH+N8xXK2PPyrZrFGbsuyPEYfG/WKmK7lE
E441I2dOmdss0E97CAGKjyM/WuMAnzoYNdVMFfFft8L1K56U50bNaMBh06wmXTY+
Vy8NwfBNXtkKa9qlBaGLpeRVC3XdTOxEmiZL6r73bJO3BdIXgHxryA0S15o6Cr/G
Sh5LYay6un88H72Te7IQJ4uy14BjUQUjCqObguOMn9tVHAh20+JPA0CWhnHjLfpR
6rR9lxgvkm8T5bL2HT+Zv4K3aqCBpmoxADMHJYRHdlYbIUgX7kQAFyPgAu1/PUZ2
VD/W45FMjLtK9agbEEhRU9vo3Gl08BWeERQrDBQRXx1VmgDar5I/6kuvBNJZ8cdK
dVFHJHmh0KtCiH4O6s2Rqoy88MiLG5HEYTNMzIRVp2/H9Ky7pBJV/m5vDxJ6A6Zw
tB4l/+Ly48KgZv0k6Z9bT5dQpF+/luicC8M1VnEPvkCd/Y3BoeBr/+c7HwGAPzVV
4fffhhfXaJesJU4PT5eKBCvrlrZcpN2G5xMjkkxltH00g/Ml01BP33pj0jZ1DrNc
PA/ri4a2SX3CfcP7HUJ6QQITqCPKJDP1v3kvTjT8ZtSphjdk5jpHzAJg/fpUQzW+
cBXNag/l8Hh2HB0dVvyLTFupjGrXzFstK1pU4KAbtmiYIgLELIUiAM6wLhSM5s61
hrfEKTN44M4QVj+r/EPb+oQ/GQj6x/2tnTMK7Rg+Rsq/iSy64AtfS6yn5iC32vER
OCl0GEzWqXGMYMtf1ci7Hqca9oC5R1jew09MocyiMdI0ddvkS7nyRFIvMX+s8bWE
H5e8I/WYW/KCfPrtbzxF5iinvzdwlnyEtrE1pa9/cpKzPZC1exP1Gsv2ARLBCvFh
0dNBUIcuTTQqLX0z9nYiQI9HlBA0vP30YvQT+HaLcZwh/qlYOZ1aKqgtg/rrHFT1
GfmLNOTli6uWyLVxc50tInewO2D6I7D5UBs45wE645x8VZc7/3E/ukKS5KdtC145
QOqz7RSgeV3uD6y3ns08XZzVRnb0yFEw6+AmZrkYoMl54d2MjCeXYushM30wXhCO
ZZnoIZdorIuF6ug5VPoDeBqm7r/kUqG2HxDBI7ZLFwI9D0GmtXXOtD+UhT1YMLKg
HbCMQFHXKsIprUrdFWCvVSCL1T2zBOODTn09B+vl4mOJEpVqKRtYuG2kwORd08Pn
Y0J4ycDFcRRdEU9n5o49YnIdMiZKa7vAoUfI+1mv1z+6dIsNg71TYo4pBZM3Djf3
fJ/7Ad4xVR61cHG8tOMPmMjR3qo4W2qCjCiFOln5yL3MOu7TtTvHlUVjxEjnU+ue
0g3tUJboMpIbnN4o7gXMVbI593oyTIkCTKrSViYUbh9ZXKWr9wzvwSq7UHqveiuC
wGOoA4Tw0wD1LuAtoZCyccGiVmSdCBUvTUGDI5DFrVNVWCrnZ6mtSnZAEwqisnVx
o6VECHh72vMTToDVeLX3qqjrlkuhsw3nb7i51mqj+4nkJibVZzhzZHDEwykD/MfJ
0YMxNrt6H8rfOq0neSbIj43CiAdKeIB4PsZOUSzlyablKD2Nvg0BKC3JPj4VQyqI
QkOxMq7vMIRfnEzkHqzRYm4miNTwv5mY+1Co2JIGr1rDHGfVbBOG14avQ94700F2
t6S0cj7s8QH4xEb6YKG/nRr3hQHaf7+2+j+p9p/XAjXpC/NZv/EoV4Ppu8DGRVQc
RcnvAmKvo+onqq8NVjq42NPPFlsshbW0OeCowifRja3ZB/I25XTzN9dY2Y5ZfwcI
8TfCSUZelPHX+mGix0LVESnSax69P5CmYTEuCTZqpjInOiD1vH8Q1wwI69arHHgu
dZXF3xPmB5B9adCe8VC7T6fTlCDpBga04VhHyK82tLP6zyC1EydCB31xZ06qae4R
peHBB65ltPTrgtsBi5KD1O86YpPhqEq9WQEGlhAiGuMKB4qLdQZOacU/z5JFsyI9
IiKxCLrV97Gle57DRUOqGPHipOewDPeqvMIkXaQzlaKe7wwS9EU7t73tawOd+k85
hFVePqnMP2QUQmbBs9MQoogsYLgiSROkyOBNwdHLwyyE7Kqd5rmcbRQx8QB5cQQi
VRizFO9zhgWREsLBZIhlK8+m5DO1BOZ+VFbJV3mp1Aio7SoYVfXylB3ipEIrgXxr
jz8N84DW3bJI2gOX9baLa81GI9vgpakHPedgY46XBUd+QLUG5kJb1Jp3wuxKMoI/
hIT3noYOCY8AYnDn3satY3WP/eZee5beB/AAUjjL5n9MI1qcFYmv9vbRGZRCkE/X
oBlvnEfR0Al4Hlzv1b0z4tDGTtb+9jrdoNZt0PmHZNq+omal+mkeAOtOthV3yE0r
VTORh1WvCGGaPDCUI9LwirjH7A/UsDpQT23JE/OnPiajAgv7tDGNrWmSAI/BFwW6
roprE4108nV8mwCm8V4uUdNCL4ZmhefvNL/BaTGC+CkA5ap8CHWoWxr+TNY88DuY
eFxWiJChGmA76isImWiAuzZauD2GNtuRgU9Ezm4TD2btYq3nfLxGaDxaGaSX2Ht6
shpobNAtdX9A/CuGiJqBnk6P4hNsKn9oJX0jrTUf4R0kFRorNnP1+YrCzZ/7/+ZV
JODls6eOtGumE4ZpJg93sFYt3j8DCz0g0eoTWzP32n2ddKly0WWtpIBOMf4QRomC
M61Y0V6QTw0Iv21ECJCWGclebEuCxiiPBOP9H3KqEsqnxo1n8AinXgdiL0YntuSE
W9G2c2hdKTpP+ET0P2LG/b5jR5JY+Am1VuZkvKeqD/DfvgDeSQ36kJSDHA0XQR73
23LL6+fIdMBFjBLLTfhjoWTD3hLINxaStDO+Mm2/LDjOWqI7fo0IkZF1m0OrDVGt
DyP78T26mzqh3K0/G4TDird+Diq6GAYCoSfFgfMaJ3n+Li+RRpcNyGSdpjuDHoka
qtqknM0Qllycol+CtV7xNCDdlWfcPPWp89WlkPRUsqAyb3/4Jg5kKSWoeY15nbJK
aaseA7rrMxhM0WNL6TGlQOCfJFJHCFj+asZmEeLIF+rakaDYvz8wCON38ZqLe1fc
pqNrkeiaM0zkQKgXkidAbFuLP1mWsKuM6ERohrj2RgE6SENtcQEe+EcuQveiQ65r
GsnQqcog9twkHMNTTY+QiEzz7V5l965O+reg717OcKBQ7K+lG07pS2gF+RiGHOEf
cC7Gp2H1zClrSYfhhECup52cZDBsRdmgvECxe/Aqh5lCqD+0TQ/4wkz33T6j5k76
dEU5KIpnJHLDshgLt9rzhTrjGkL/7n78IZ3vBX/fQdR5+QRQLZmMuhri6NHQcNK9
HDYf+0SS2vn2PcKIufgnIQ9J8nVYwqeIqR9+FhuMABj2WMNDXE11yltdd1Af2NRj
+efwuuvMz9snDCPLbjiuPGadGQBNrPuFj0A9E5re0ggQE7tLFZBPzJBA+0SGV+7i
9L0WkQA0S0qE7XvGgto4wfkQslmDmQJ3PW0lhu+RhiD4N2M3jd3xFlzf1ryUu5Ks
S7YXBMbSDbYw7wyG6Sg9y+opLt1rScO9ssZ07caXIxgcX8D1PF8rlVtujeCHIqm2
m5ijxvzyQpK2H7liGRAYs3JzogwV2zFe4zJnsolOCPpU4yzHC2tXqI2LrYfqYcFq
aWSCEIXoEheTapNd669pCUO8UEhBVoKzlL8tUXNkkv6wYFGZgJK8C0MP8W3msS/H
nItsj35z0HY7C2rhz12VZfm37WI1UbT5CzKghXh/nX12UCKfzhzkKkNTeqw2YX4s
WUeHuyFW5ShjTwVT1ypYTSPn0OPme9mpn1AFVFtpCVqRGnj1TWgwzY/j0pfeJBSB
wj8QV/85t+4n8UTey2OqT5ss3VlAj+nZAoVBdBGiJc2Ql5z3Jf5Oiqsg8ZS9AXz4
boC9EOweb5XnHqjOQbCVqcYubuO/dlY9Tfxd8QMBD3WNm2OxG1Fd5cFI8v4N0SLu
I18xhp4bscIzwn47b3gPYVTOKJCWOgmebYrfTlWk/KFoF5IGoYPXCIA9bWzBJM4Y
jyDC4JeQNl1pQ4bYqUyAINr5VGFdvr1lAX6dhKJg3mpxVw9LJMia4TpepjQUmjnm
j3w74Wyjlg/IJ+2ai3MQE/E0csFJ9EB2gHGknoTlgaL19Ob5iGUBissAtjxuT7uo
ZJOSYij7su6GlzbABbI52BjT24YiQnJIjbIRnhdY4ymp2fCEpokJQ3+OKatN7wzh
in754DgATncUTMKA5jZm8YthiMUHUpzud0U5RWnKvCyHRkIal/HHQlgkytMn5ps1
tztIwgID2LN6XEiU3mAJ7DULOV+9B4IOf1+uOtS0cJ2CTvbFU1wzxAJEdH6jvGiw
ieMRdaLLBgZO/rHQHeIdWvdRaT4Ujbv06n6Vy+wJEANqYTQR+3GDd8a1Wla+cGpq
ucj+0kodO88S2F7XAKY6dQPvKMduw9csuPGU2x18YZMB/M2ife0SI+LY+qh+WpYc
Di/SI59mp1wiZkTd8vTCD0a8HpE9O0CoZ8k+TI175c7gT4EAIexvFYG67R5fID4m
Jxjo9hIjDdiNCvNvj2K723munqxOlQGMqlR4RE86/j6K3Do0Wq4YIjZr9/wnKKYj
Vkwg8vpnwGKrAoP96cXp2I6inq7MZKg7NP45xOr9ounm4lGxWQ3HA+FYCxZf5kOO
X0ZMqGFc9wHhgP8WXAHHMFx4eSzI1D9JadGJi4u7B9XRyx4jHR6AtJTq7oWlEHAi
aOfXqy+8ENsuqscq5OqyJBQclMDo+VN0edF27m3IBOZ2cJPygwkfugJJ68nO4WJZ
GoQMxJJ5veaVSb9nfg4COdFsi55+sYAGRUdtAlrYMyysmkIQ19aTy9vvg7xtTT1i
4uTdvre0pLOxbsjt5+kpSWNdADnGBFpLa8OCITYJMKEz/NgOxIXcdOPOLML+YZXT
ctcxGWDm6f2zmZ/m4pnEZKMqCING/jcFKpAWKRgW9p3NOItmkBzdsqxVdWN9BPXj
FrSZpFineSxWsMi1e8OPkcQoSaxm0vVXxjypVIZnPppFwI+jnaItHQwhf83cn2Fb
sv/GGTydLs1fpUO3f8LSUbuNlWXq8V+FFN8AgMKqIH0H+J5CGGgY1zhCxWwMQvPh
n7ULHo5Vq5GYylwB87wCXOFz+yyh9XGAHQQ1fPQrzh37SVOYAzGMJPVtfR/L2SZ2
eACaZPs+dCCEPYZatuANcI0FCnMj8cKtrpVUgsEP3SbFa0FrX6HMS3et/1diBycH
haELejzZ7t83pJveyIaN4TWfDEL0auuGxjgUMkz9RyHGGVcPwm7YKrwlssQn1AIR
BIyVpG8uDZcGyRWto0TOTTJ62V6S/q5z+vEl0uANTgQtSq/dozCpWgouhiTENsNA
TFxGYXc/xAZnbuyXeC/r6RuWEwoA7mAUckt5SCM+somvUsnrtbDE2rEXnt3rf5lR
mX56v6hTRdo4tRvuPXUN3IExVXeyLE/Ab+swYYascDtrkKhqdp0iXeaILfswialL
+I27fFCZDIm3QDo4LbxPJUgz3qg6lQ7TNKhbVsHO4vU7+NMcjlcLE5Yek964woQ1
oGcLmZ1VHNYB3t+H9bItPBPZtdSFj1nwvm/OyvyANWg1O2QOdVSNsn82FZyx1ziB
5Sq3pI+wTfRP23KTeQq36brPj/FOleY03dOsokCYrBOfNXGClP4SsgFnCTwj2UMB
MeCqHzhv2bp5kXJR0a7B3uACpYgDP9m+gHR9pUH+xYZVlcUXvVYKENbNa87YL+11
m6+RojlfInWqrqp5Zw6J3OTWhAodf1OrgQKh/tbgh4gcgI4Nnj7zNfxf5IPCA+GJ
6Ok2LAN52WLwgFZOmmqU+QsEHjiR89AQoA7grOPbJdcBvbjUdDMflSdH7jjM6RGV
y0joArZ2LiZrUoTkd5Mbe/kkHZBmNo3ElFjlZNDZeOTH88Tc6y2E1wm8AWeolp/L
6dDPuy5rI16tNlGQM19roy3TxObpt4XwMuJQZ2rsbQHQ2UTko0AqrT77NIcKHoVh
CMHmzQ/DEPXqieS6BJU1PJOtqBLFi6HY8SmYsg642nSnIs9+Uw5m5jmabCUlEWGg
DbXn2K0lk632omvrLsiG12eEmf1Z+7Uo0aEec+5+J0AzLdl5cLGcwOfp+cVxm0SE
Nw0SbuQPsSmFp0vefx/xw1bjoMEsMsLfPpFKcuzu0MrQe9qPDvXwYYaxoEalBgQ2
hJyf+/DOYcpuy3qY11ycveUtboEPFK2kZubeIpnjTLc79aEgAAP6Ep4H71OgntcT
qGhqDzFWMdC/Ji+NP4yF5cBd16vISs5EJW4RRkEbsk3RdoMeFec8pyZQOvdSLDMl
hMI7UDFnbr7Drny6Uh8DtS+S4abCW01L53dHgfeFUqN9RofLS4hF7mdFRHfHG0H7
HgRV20lTvdP+vuBQlnWzPd5MwOJGB+klUwnTpGIvr2LiZn8bOQEvAG9F3sGABc4E
mHpQurqNghu/JrIdn6t4+lXuYNSyzLCV+FdnEB2gKKVjgeyXjYJI9IYfsBYfKTXR
ibiPsOg8UfY4ysTuD9Q/EXjdZ+dTom+VhMsmEJthj5sYD8WfL8twxnq4/cn2Grhp
G6guAosT2ZP8d/BLcBNbFbm2V62rnwxhdTgFxfaO3pVIZmKjfEOg+pkBadnPMJVX
UM+Udio3Q3opWaK0ZYwSthuIiUKq2OmX1iZ/WKoIE1OH89Pwgzt/LGSvvg4hAfm8
0AIkwl3ns9KHLByM/+jpHzepu9lkryIATP6GUce2DpetTgv4TDHEu2AcGNSWUccv
DxXq2fvetFdEHdKbjlZMPdFe2qCrIf8dU6xiZiwbjOaCD3okL06/u1BHWUuieBO/
eVkNvEkCV9CyV4HwmyIHnfPAIJRwvLFeDPfCw9H4e7mCidCDbMJyFlJP4yVOSClR
iDuEfT9a/ybkHkComYCX02z+hDG0cmFFwG5xnBvYS5lLJmZUSbKwuJXq5JCr+r1E
aRmhAjSFiFe4+CtwgW+e5DuNdzwZXLLawpInqA/R3QzwhaBNQIGu/QIG37/kPzJ4
zukrwWo5ur8DQvrckACg7ZdCTu3Ub5xX3JOTWIGnxRrUTDGbQU09eFH7Pd+rSyn0
MG0Vb+W9PMrWtvL3ZJMX1TIKuj+EfIH5pj/BwzifexkFONhp98xRwxQ26P5R2Y6i
/EbgkGSyHK4k9REzOTIqMyVyc2H15Sjc9IfU08phdxQfvq6DCpKHlZNJ9rVMIxw+
VZ68d4gxYEJr4n4dDq8fJe1jMIM0UmE4jWdadZsj6HNZWu27Qesr1KZ72wdWF2gb
SbjHu6Qn7DIc92dWuIE5Guc6vonleKrkew8X+CIdyaEkS/kDNiqPk6EU7OcRO1Cv
mNB3RoYXyMQ+BjNhXhNCgDSTNKdQcURVJn86U6Taj1NMNRw69GETRVq63GU3eRTm
46jH6ucJT2Blcyr4chDhseQzw6vtU5RDo+FWqpLC0VW009iRH7ggQObEu1cKKiv2
JzZKTw3xT57FzvDknGbQ+lUhy1zF6/FMNv891FN8IyzYoVGn0dp0Qs6+YdP0JbWP
Ny08FYg9R9jSWx7d4hAPOsX3rXEf5wTjMBDHGcDhl12SyqjLluE6hfIfIrOD9v/U
GcxvCHX5MElJmw/N5tmhREuzddnIJbvjMkAZ9j1OPDEimgANMtXC8asonwEjOSO7
Dgf23bY1dI+wIO4n4eSTpwc673qeWWrGXtrPKrm27r6rNY3FkbkR6rOlAbdaaVAW
B00y1+5dDL4WiFEBKcyQDNC/LF6R17bJ3WxRNnBOLDr8R+qe4LTbFygliUl1mlCy
QmfufZO8QaZYY/HrGDCbaYxgfJGFBmAc7s3Mcw5RwpwR6yIUj4QVpbmJidP0695d
SroHfHoDukX8+I3YdQgmHy7jvTx3/aCXHhyoEyS5fvCL/g9dhYmRS0sIeE/sE8Dp
NscPlzztlzpmoj9CgLuLlxMlcnnFvXmAN3aC6UDeLgiFIrC0rlw/z4a6cUZh3yjC
JPQQqmFM4sOvH6WsZtl7DhzCtD11kFg/Mg8+54X8ApiGVX7GjVsM3LuXwmycD2Mt
Q9vHMVB1Ihd7ulriKxsyl2u2nSuQ4/bhkGoGROBT88g6yVDxzc3KsOsY/97oDDUU
oCPZIGnw77YZikhA3P6zWIsegsc3cabbh8x3g5LfDUOW8C6zHCL6iaQLtK+EpIcg
g0jvca6YT9HBeawuqqQsrYND1o/ccW635JcSXFelLM/MaxV2B+9BJgyA12i4Ohqy
9mxq0JIHatGSAf8jds40qB0k28mzx/hH2Kf+7DflE+cPfBGc1oFNr8+YVtmXS5oC
4jhEECJ3kzdM54zkJRXkkrgsDmFDXgyTdLuOBperkL1BQGzicPm0bYMqV+uMDSnr
AK/gjWBJVM3kUr6RBAEE9HnC0yJ12/cutWEklA6EXtL5r+7X28lMuZPAGbP7OicL
KTal34D3C9k4rpBBKMGuwDHTi5owMMNQZVDEDo4jb+tJI9AN0clMYamaK3wjjUd/
7kLv6NWrqbOEN6NcgySRgHVvSP66vMnseeNvNf2aKS3pV4M1h1T8vTu926KRmpuP
YMeQvhPCLScTbcihw3nxWQHqHNRevi9lwM+xuW3lY5gJKWoBEVJGioyiO+PYwCrL
TrhzDEkxY59q+E8THUm6IrIr05SsqIMm4ojFvRc7HDcMntGu9l7BDg9yIz/HHTUb
GEa1VVZ4c6gypZKtwMSG0VDKF0WWHYlq65ymY+YWRDYa2nYdn/DWi1HMpdgzlIzg
oIe7SrXTzy6BEXLuwWx6J05XEk633tmer9Jck/u5kwTTgzxvU/kpRNx/BsPJaKhf
pEFvD6SGZIJdEJ6uCoXyaTsfGqm6SZh050mYXEioZjHBSdPLuIH1dUyonibfj+kl
V3BZuKghW+dOK1xS+U2SUm1f2fsLaUz+72VwdEgrXEv8wA2IjK71G/qZEZgLljYT
JXoRDBmWPdo3IoCcpPHFLfT2UVd56bjWTWYfW9qCdp8LB2p7AJPBOE6AP1+8GYtl
yP08kaZFWVIXbP5+tsbW7XIaVFjoY8a+sNLtsjX4uHkXvfb4+JKyP8KQ4D8MDL7O
vqYFqtDCucMxPKmY2lt2XFF4Zq+pd2Jf9lrfExkAi7AHPqoU9q73xi5p4W1bZNy1
rSUd20N7mr+Zz66KyG1QKKxLMikl3pwE1iRznWebiJegmsOW3yRuUsbt1Jjdn3SM
7G6eBvjmVm8oS6QbADYu4Z9xtK2sjYnReAkYv8eFOJZ9SgqL4SU/3TDRJfSsYZyM
Obj4hBag0o//U7iipSMOczo/P0G1iLbC7nTdGmE5UWT6+DEqV/tLlpAARqIV/iI1
D8alpte8XLKxvK7L39pxnHyHZ+NC/MjCKF/sc0mSICZMjAbeqsTWPoh+JG5kVtzC
WlC34fWEnTtnbw3hi0rVvDU8c+e9RZoPmdT5/e1AXrkmUhWZEhjid1S73k1RzBQd
P9GJQYlhvt+HZQe78rA6ctS5khn8Gg1cP6BGC1dsLOjDIlc8+HrCoNv6m/DthuGJ
74bZbKmC3tSxhZSkM8NPq7+M5tldMra9SAXqvOS1iIaCy+EIv5bCNuOPXejeWj3d
3a3Supc3s5tHD+xYi/9n9dA2ctYhm0d4/DMay43OXA8lY8l/i+hT9mVKP7A6AkiE
7Is+TY+hpECc41nNjX7kxMAhfU4RxIpc1FshwdU/aoDtANKlcmgo+4iqDPAyiSeF
mM8P1Uj0zwZ6RReLwbxu5Y4aEC7GimTeuD3eylmIhavx0vYMC37NtVV8DgDg6RVF
pTMJ2quCMAvkW+mXMjOcMiFhX+rHf+0/qMFNKTsZVEynQwySteC1yLAffr1/PNgG
/ev9i9u+SjeHiicxiEsHpG21Hyf0ULt2PcQEy3hswYsh1ec+AwBBWXGve0kSACYg
34REes2gCUlf7guLuGVC+K0xg9lKvVGheUrsAqnkSvSuhHsqKsxgHs/rnOTnhKSW
Nrq7zPi/MELJUWUKjDHL4ulfaImlEv8DtLpQxG0ZNYGCH0bCd5PfwAY9zLyJlhfd
iwOoWLSGg0T5UdD9kbV2FS0eA2sd3d5oVQmZ70BhcFKj8cT8IpVaqdw7ewu0W8fp
A1KNR66ONv3I+TujJ1ZhVShwuuGzjhzOJADxLPN4KDXybcuOJCl+j9p59GqWB2y1
NThUoYxQjYTHYZvTmSZiTgmK1lhwsqUJzCGs0DotGfVYZDzcIs1Sn/oJvMggPnFu
hhWSseb2uC7EraSfsMKPAyyifujSwhwDrUAaXdUzSUamcnzG7RR+HHy3eUtTzXtc
zGgoFQXAtKQUUlR1rzvm/J34rlkyQTN+YfZyMSwuQf/uRzdUTJuyrMm7vKK8pDJi
WPaPYampp3/yfiuFnc2uO9OkNJ6lAP3A+5UtDUiVAeJ74K6hRktGwqjs766VFGo0
xZ/W9dKHt5THMkG3Ga0lnsX6GOwCvEz1WVwqsYeMxeB1PffvnVQqdBepgImjTmrd
mtDDmwUqgQM14PPzUxY1wApph0DGYpFRV72FBrMD30NMQEvBr58t7mWJPNae9XST
hcpjilbMXAd+Hd/QzzUn4LyPFYXsNA/fAKyxyJjb9/6PPxRohTS2Gqh26IcY4l1O
brxsCWqKZYD1p9hk5cPWBeFmoosI/4tRzNXcaTqWxRqvtW0Rr9d2hYxQe71xBwNt
z+34z5O8WNiXtoxbsqILu/Fh9px6pE3nFVzEl23CBfFFI/4fl3jmQl4wmLY9m0hk
zXHuVuZefgpEAZZEpGh+lFgc9KesK4oZlhBFmNRUsTRzMRqTFOZQFWSTY2yMtPNa
Lco0ovIJzDSwZ3HncLzHmTnDl7eDaEOzb/jZTDT7Px9EhRpFPzuVEG0EiIjI0XCh
OY+n6R34P5sjpPF+0gDDfSaH3g2ZPFD0hpy1VY2eF0AnMMQ25W6pPaivQYUwY6Ky
kl2khf/g9Lf3Kk3rSsyouTJfIug30tAYb86Z57Fbu5U//wCgfJAf4sfl2gwSfbvJ
htverpxALg11z5aH+X0BEW9ks6NPkOuyVVqFqyVaPwtzlcg5ffux1LvZ+6tN3Jm0
451zP+kpzsAV5uipiWpR2QfyPmTZCUYmKVfgaMZFjiqXU0vCTMY68dvynQXUdVcl
e6+Fbm5mX2OZ/nLUHFCIx2XBiRtkxf6TDIkp3DeqlHxJUU2Yt6lMXpdAxmM9Ps21
hwJM6Dk6MPgw0b5XXeTvZ5Qw4Jo2KbpBA/aXY+lRTCP/E6NP0PU94KCFdKh4iJYI
ollALl40L7jMo2EoCzZE8HaGN8JlJmxSGexLhu398qED1JeaiKpkcJRWUsz7hRkr
G5f12ZPhDgjrAHCr5+A3qJOT9qr/IfKb/SIb2bGhUeMfZpz8qSNkLZt36Bmd/uqd
VkrzeLFUA2tI1ptuljdXiJLqrpxvCG/4fheCs7pirEjpD2poMD29VyfOlScKzfcW
mBkMPU/GmNX4816y73kuhfwlX1BvNIEi9FT+cq2jUgDOgnLapZ9gtUajxqDI8kBp
HEVm3AMjsSZxIUVlD05i+XxmfyvK42sqOay0NL+Dvq5kR1jOzxTMdPZdQWq+6nxp
PbaW2OfsnVKLOpsXUP7gpZGmootzmAxpiWNrZaIOY1xprAbMoYqahu8XcS0Bybwn
MM8lL5z/FHsG0H5QmuYnUJQ79MdW4G2f7aTBaQw9ZpLf9DEPL1TL77U1D4zf39xw
cNUSQcFDoOjGT75wM1i1K27gksZM0UhGh0MJGYIPXvo6OE2VmSRLWdXWPJteXSti
R+VViWnb6cmDDe8/PKGWmnTWaG90sDyoq40QjXjYbJUaQMmsNHwoUi0ZymuRuXBx
G4I7fyqdTIvWg7jh+JWPagF0tJx2z0R5dtorBu5hrU2QSw/QV3pNwKf0d/iCj1YE
jTw1DSRq99R3A3lD/DnWx5fg0idHqV5DfNYJvJW8N6DUX4qyFXwLQQPH2HgJmpkq
Odd86TeaWe37jz5J7SJWyLZk/6+gcIrXtvuQRdFOYp5ysLLwpFxc7cT9r3IHrzyz
W8DNrY5msjT3umBA6DPCpyQowY/o6QrbImW8gWehwHIDMzOEIInv3yNoPPWineEX
3VgL1ar1jneXsOPUsEyFNJpN7Gxqn4HwWAfb4OjmgqyVXnwv3KrlUc+I7DcM0Bch
wja2hlklADcgY7dANdTs7lLajmChS9U/bxhQvNd12JrtwFq6xsMjvjyA2Sz8bz0U
pVmw4hAW9t738IXnU1GqIBt3bcraNCUs3L1Xg3GnZe3mJEhwYILvfJY5dUJesP4i
ATpuiXoSD8bpU7BQmRlRtXQhN3eKKiUfU8eXk5ySfntgb/ZmdwkVmt5hgjeal7vM
CQ8D+R8e5/Li9JNoMEb94v+8v25cu7ySZkEnb/sox/lxDIL9x2u4796QXoqDupKB
aV02YscPTEnYUSKJvUoAkaPK0VHEmSImzWWf3cfVyIbQKAFPwxJwRxj93ldGYmAJ
oBS9l/7seCvvdyUct6CPHLd8il49mA1S0lovEEMOGmJ0RfSb613TXzrP49kh42er
Ycxuuew1zSUYFr7Kl9TnZlg4QPDnMEjWDlexvpD8ETq6f1sbNZRroiy2fisQeSd1
1ddVsFiWto66EGuq8YSNGvpIXdH4msSsBFqXThR5fGSscRsiK0YdKzEThZpGFIeO
OYR3qEjFQPVG44i4noNWNqbdcDh6XSwtD47ZGIf07G2lIX779KNbN5YM05LdWM+O
SS7Wcj3tA1LHZ1p8CYLYnhoGzxz/a176nC5CabYoGdwK/2GyLwrBUUmeFoRW7WmO
Yw2gUhMvLA+9qrAzu8AlhcEsyDPdA+AY+XwzW46SP6tN7wu+UxSI+vTPDUBI4Rz/
MpZvOYT19M8Kql42xf+WtrgxILD6stoL3+A7swbZPoGynJd8ZryjiITxn6YVPdId
BR+la4VGJx1mOa5qNRSftOiqqfi1A5st/IRdv69pZ8QRJtWtL6R9tJfyP1XIFZLx
ywfv8fNUTO0GdoPnDyj56SaMCxnYd5jXFp02gfKpES69wfJiJjPukvwkjErXkycy
BXWsQiAGbbuLI/GJGb/GJHxS7hUMgrCK2Z/2seZMKhH+/m//q871uhbG0IkKmFGh
7wjqSTgtQruDnbKoyhUj8CzaWgoX0qohvrQ9PbJxyml3+sLAmK4/QWOwP4OnN2Iv
AOVySfi1H60FCm2ZF6vpdyAtrvCL4Lu1egifqqaTbZSvjdwtzrIlyXRnDnSYiTl7
ZVZ51MIUBhOWi4WJJHqr873r5a/1esrYdreuZUMwklyoOou4+Wrs9eGiTrND16AB
+recjSmTiWtZbsSNDda81dpsafSpA5MSTmQ9EHgmpBJWTuBmb3+DymFPhnCT7hV9
/GQn95SnL5X8b82gcXz5LovodXe/ilA6NsAwmESnqnL2mUfLa/M+IpisJ6L1YTpW
HyJO6HRsrhtHxbAG7zNTFvCeAIIYtHmQVGpykHtai9Q+FsmWGHlTIkegUxBWDVVv
WQzKljOIcWS5CgqkciBSBD1RtMXcjya6OmsWXkVUfkBGjM+ceqgSQP9BkgAOZnrb
gfMSnuYQsgTbDXiafsis0dLdONiInzX2EhtuP7Ma4t/7IRzYbvusAJpBtFexBfC/
H/9HI20PzmPX1QPSSj3k5GGve0UeSlHlb5+tOyNddy6R2Po7slzc1VyFMjuEldMP
XIRVtomWkBe/xV8hUa0KmF8fQsEZA1VX7JERu5Rjg1cjT1n43qTwnB+Ulw53d/fh
EDD+YVroUMbzfLr+jhMbuFKB8hw6VTm/PVE4UROHT4XZeUbw/xBdy5vtGgiPD918
MQcYERkIOfcxT6AjqzsQHwzZn9DRKMOlSI/BHpx79ZdCD10O4NvuAU3JL2upWUqY
khMlwiKcdolKvL9zYrlZ+ALghHzyDCTDGvPedM0xcizRpwozMP1pWkI+jfy7O1iH
cUt3kgetnO2ALLeVhM+zYt/NB1SKqk3GaIPKsrnxByJpolpjjOdsDpmfS77Xq2QW
GXMn1WviuPvrFOqoWhMAzlxlJbTe1BkblSdYI3/N0Sf/GoM9C0rQL7D7w6Fsb2LZ
Q9Snld081hBfrB+eMLcIzj2H0Eam/eXaHbV18Zsp2hy+FhmRMsvKSSox0kRJb+Lr
uS2VXrQ28+mR5SUbZIPQwmN4t6CvlE1UsH6gvr3xYHPLxjZ0Lcx278XLwhGI5WBd
RhS9xKRpLQnt9T7Yr9qEFY4KSHJDXkjxVb5NoHCVg59Q5UJrA9taGCUv/eZHAq+q
e4KQeVJHW0ap2aocJC01d2JY7VqTaEyfCg0GAqBcmyHmCGvUaoYL3H9NL9RxZ3UP
Bfo6GSSRb1+7X2o4H8gLGpIiMWrOg4r8n62VW0twkX893F0pbF7EXF86Cj/Ryi6R
nxcTCdIAS0AvlCTS0cJTghO+DRH2myOb3CS7GL7+oKNmsIWKOvmGUS+cnzanFnDB
A3DiIeyqZGr29REpn0Ea9mnenik6Zy6+mV1dGfycePKtcwT7J8MIDm5bIjidpUA9
uMcZuF1+/nIUZaIRK/9ssgbNamITDAh9lIq2u4dCuX4ROf4Ui7TbO9ma8AYHit7P
tT/hbgoAhXCdCkx6fGtaflfCuqOT/SizTAzXF4rAbmvHalZb/FHI1kTHEOAgsz+2
CtSISmXDTmX/hvfvM1kgFwejuUGJQdCyvDMdW0Pb4ZPKAOPLbqJk42BklFyuFb4T
c4kM+58giTW+ORbKux8v8yYZC2pKzSmODsbIirrphWzoh4pXtg8VZgOR+hrWb9Dm
5YJg8OXHcwK5a2AmmmjO1zluYEyNuLo1auCKoslttzCcKadwcwMVIUrM+jqr1pHb
+F3chFvIaRj1zoJ/7jvDoLOXcpi7dO4n0Vmt0kNHJjQzNXXI6FAv+BRXK5elnxBz
3SjKydsHOwOTdv6w3A24ith2DF6yZ6MHq2wFQ/gTxOhk2Gs6ztWK+8z8IvAqrZck
FKOSqcTlN4O5JnEU9ZWNopaz9vEvtfgjTq81VDMeetIE92MfuU9quhVgLC0oEc79
5vQIcGRhgR3TZ/hETqN4K3zRkCH+qZ+AKbJjiacZd8d9PsE+ne/7exdWkhlTc10l
JkkxVAaIcTLUhspxIAC6HMKZnnSH8MDYb3WDRPSBK69pU6zt/um8gHAscztx7/ev
GzpnFLFh3XSgTpE1QrHCqZgSUiVw1LFKcHCieULn7VbTQDR6sAq0m3nwgOpWlLI4
mdleAAgdgTLqlnTSWGjk08uqwrIJdqlnVkPEvwKyAIZU19wSHhFBwguc2YVGr58n
uOS4Owzdz5zGjMZF/kzFSzgkWeNj7JW7/N/QoKrBfuua2fj4YUr5c3GKttTEhDCU
S67nz3dtMiBRwQZ6Ygczv+Xw8RlpGiCSX1OOEkYKknMHJTYyoGcco4Gy5clyKUOv
E7yGPAefT4cgwjRQjej2USc3jzx7LqHDSWKoLNmt4dE7DV4IS8MmPQ8yh/6TJGOY
NGLvRfg5KpAAdyGNyV6grd0emyw3JyZ0oRkRzT60DO1HgO8V4xJcUzMahIc9DiQp
0trCKrrhChPJdAN52+3RVEVKBmix6fS1ZJQWZEBGi3KJyAew8QqFMXzbQPedjj+V
vZQQs0+oBf7zFuDVSz8JVHWbA2hV8rjQhUt57ZCZGGGrPng5LlrgFtJXq2MFWBWn
8G1CAJqYiUyKqdIdZau+MS31f71lLcUBOMylScKvL6dcpE0h8p1o9bBXc8LhKBZ8
0lsU42HcGBVbycZpfMNZ80evp/qvdejvPQfy6uJqj9/wUKryW4Aclmheg3DUeQDA
FdKi4iSAceKnpLc/wJ1eq+r5/n19Jft8X8HEraPcbb+Fl8lOjGFTV3bj4c6yb8/c
SDb6T1noPyvMNNoYIczCmZo0cIbjYuksrSKIAtytUU2EBY9kVBfJ6+0yDcNig4Sw
SRQGHoFgmtzufRInMxOjn866zv/bKOnvpxTiVstMhFmkD8hMKDMAKMYJSIfoojP5
QXXjWaGnR3Uh9Yn5lLDWfjxvcSQAbxSCbSGSkGZcbG7FNtllxLcjqR3AW1j7sXfZ
yM9/zMU4TyFfTFXAv7F8UIVpCpLDLly7vY/aolTGhPfsyEA4KI+cJesZiVuJF9Wh
IS29iR7TlvlltBOBM+0og1wiA6zsFIXhOQh1Ab1oveNSq4h47pLG6Xk/pLyRULk+
tJJKAL/GqbY4n1PfN/Dpv6jrA3+YfaSd3Q8yjvMwW/cLJFlM8twJdWR8udGqitmu
HkLGX1A7kl6ZNXbwZh2cUWPNuP8kBTE3bAch+im699zI7ErykWoMOT5afdZiyVRd
Uw/UuAb3H1Xs+JomfYrF13blXFObsA8/tF4U4kjTLEMBg2Gqqo3RHY2E5qc7Kngw
Cj0pGuazT8NtkNZuKtG7cl6bjZHuMuzcyOteJ6HxIsULqwvEROsXCxK1cEfoPkuR
n3vL5hytO0+5t7Bn8JoClBeEWIjHk02UMLNLCZ9SIdTDJrLXjlkLgDyzl8gNZgOz
+TLeFaPAsXiesA1n5YqLx42CO4Zk5t+1YJZxYxxHbIik0WrwEAXtqZklzTz9riLw
/OkTdgUOMGJr2WNnHK7fZVHXOUn3pvgvltbF5Ovs/A40Qa8RVoLtxApHMroc/s9U
bOVPxVlGmVack12fBGeSrtvyBk1XnO4TuSziCwmqhoR1BQBCcPyS40zktm51WHZx
aGlOWC9dUSRPWKplmSFMFdZs7H1x/e9AHt72goyUHgxkc75+HBMEWqO07dJkVSc9
qdZSrCJVLSTkwHp3AWa0DgjqsAEJmT48uOw1UY9mdgn2gthev7FGh/cp0+Mk4Ul8
NA4HpxnfBpJUJjNCYOji09pmWhRgdnc4kxNE2vjF7AhMFUtBmTRKQn0CYBRDU14S
EXO+OytfRFGq6FhtNFk2/Mqd/OS4OLiDXJhQnJY4MLAujX1iWmbu9FoMC3APvi+3
vbTZCsZxPFmPIVkPL6nDE0wzXqxKPOn5+mP5aybAxTPX5NZfcmpzrfvvYy1/MHsS
czUm8AtHZCOddP/behWVLrFRxz7E7Sg0rn62SqyzYkVo6cVKxxXDScOtxyvnslDQ
g08SC4YppcuurgjRjOWIspU6/Vb5n1Cf4KqJ7A4/jw/P/0bqgv95bvPyVnM8UETJ
i19jt1fu5woLccynhwgiUnTugJFoQkOcbQ1NQLdLIAu7qoLZBJlBkImxtkw2peCw
1brIpRFJJ6yBMKfw/DwOJcDV4nd/aUCyep30AyHaz2pISStSXPTd6Lz1UrhIRddL
I7PRAw0SeaejEs4SsCGCP62fWhGn1Dup4MMhLCVYMb4+5wQbxdxuDABnh6TTdf8J
GMuOKL1PiA/d5JVRkq0mq5KcifeX56QJx5k6J1yf6T3I2k/VdQU+KKathss5ssVT
nTrAZ5HlKItQ6b7P/T9QmSLfPCte3FVkd4kHFD4ezPXNf3M5UHRQgPhnZIadgKTr
OastxOy2KYjTN3yy6/ZyIdjHTIU3gOd17R2ujH24r1ttgzL6IDcJ2NAJjanH09vw
O2l8TE2r7csWjv5or6IL/FSSG9aryQolju6yjVN6oVG8WdEte88MgF2468Njco0S
Jnk3XlWSimUGaBGQwGCK4J3z6zufB0v+UNfpPpq6wnh+0Cri4vbQmNNPt8f5VQ6O
FNe6tiswGsq+McC5X1UdtvOQgaGA4uIV+IAL74il1YOFQNpM/5x6xWTZhHbBWVy3
6/t/ilzfaea7lh0KOFrhmXyxtqmPPAQCFVOkvIET5NGF4w7gIFOByOL2QVQ+/POf
Hk66IQvOu72VHQiWE18Fg5TCXchrdQSjN9XTqIUdBvr7EuFC0VvPxb6U0tn9dWre
OmvHooE6vMLjRTnZwssqVY8xVY71IDA5dpLnUJl8iVVuYNtYDwvqZKZ/idGuBwVS
Q5JQJyv/+5faHWNkZ9g86mgyFX7feTmv9PBPST+X42FzQEmM4KXkEauKzNUwzcWq
7VD8K1NJM+ng6pLDHmlayQfQP740x6tK5gGEgCx/onTNgKBqwC7cCCGJ3JLWU8oi
H+dwOS7+cUMynho+ZyofboD5ZhmwpivTzHsE+/KMnzZmTn3gDdriVMPMguHED3NK
94q+Nq6UpDW/PQ1y2IGIAWhudLx2RcALA0GGcyBJsk+Zc/k/C6StYwBGnx4f/tWJ
/104mnionGrw0/Tgqmbzj69kBgvwnRM3+JbJQY363OQ2SxS0zrCQiQBdxKx0EveO
M33IIRYhpKA0qZoHLLdG1iASZbNnPOONVJlfsb4f+Aul9FnRRNIxbdI56AXBIOOo
fw4DekLcRJDOIHXnqhfhHTxWKER4Wj98TROo08xeP6Mo5zbVJ+beICiI4PE+Ro8K
OwjO9MX8RSBAEhcTIGvqGCfbBeFcEbcKq/QKugjrgNSItp2LbzSwuHPEuAgALvVr
NdJSjm7P4KqI1zk3wPMqBWP+0BVqcoh6wLoZmDt52xib1tPLrIgBHKcOV/3MBvXW
asfIeEL2PiOgvBtt6zuXB3C9LYv/Ho7tL0/OrH6PC5SxgChGHG3ZEyOCdVxlYPhZ
10ySfL9/Kc5OtvdUdF5iOUg3+jiIn29CSC/z86RbaAJHKTNnEF1GPNTK+8kFMfqC
ITMlFFWtX9UGEdCrilGnhYgs5EfieLE+0wjBbn8HwNYEK/xXQcA9Po5sweYbI0UG
NhAtLweb7d4JMq13iRa6SsIIhtculo6BicBg7MtQns5zWt8ggER0v+Kf6nqAX7rK
7lT1M6q+5p475HxYf4mgSfRtLdBU9JreKARDxedZOJHjXOiFw82PW7YzaCy0oyno
+4U5WAlAScNpSXWtUFthYATrZwXFuo0qYBjjmwAIrsknkGvNTQw4d/tcSB/gHGAv
dCJhKTxVBzVb1RZVZIjKQcA7AkNlv9nzDHILXMWAhgFtyXNM+JwKVgeVD44eJz4H
lB34GvAxiIrxpMPvWmVYDGtc6gFvkEYoRvT73pw5BoWuyPyV9TP8onnmw80ZHDeg
gyHt1L+HokcG+FzhIzLfOa+StGD2s9Xs702pDlzMG0pZW2yF95NV8O86NNiDP59v
hJTw6JKKY9yrhmX+/lNhjrMHDqqdSvI5c35p4kuI651EiBckf8Rq+nU7SulOoZbx
qJ6FjT12f4q7vPTcNeUTou7QPw0Yas/0YPzIC1g8HLvpWeFIiEfx6bh1ZkFiSg3S
MPgiC268YXFuh37jE9u3Pl+eq64OsYvNTP7pH/Nz8RFAqUd8Y2Iqc3rMapsHCZVh
l070GV05lec3fRLkvj9wh83Z3+Q60sJz8auKi197bUYncwyN193A5ZE/IoKe2OmX
LY9ZkdCQhtYRTErdX5L/kM001epeyYs6NCW+zOccknmT/35PLxxwl0eRClMTvyTb
LIbJDF1AyzSubAYLc7vCyPge3LWiHYiw5hJeAPLxjZkCvhnKnpA1cvnN8BEzVpm+
LOy/KOmor9Ppr+Gr7wutGV2D/k1QuiFNm9c9M5kFDoQ6z2deQA3qkYyeWcKtRe2R
em7GZj9zf4gIbV0UirOdidwauEBAl15Fw24L7Apftiv89dYLJS2jcBwSjvm3PO+F
hzPy5Oin7AHjCLRX31IXRVasmQdo2PXzmhds6a5Ks4Q=
`pragma protect end_protected
