// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qPSiqAVJl8SinXah4sjgUaO0LLENN+LX5PZ+WiaZaCGK6uRY+dgqNvUkCDP9
+cSUlSGRdVNCS9llIKxKSo20Gj7brNvwKzZ5L7v/T1i7rytIfTUPFbW1uVwr
TrUmvOG3jV/nmS/VcYELC8CC4sYYdmc7mjCSWX+NOsFxoZdr53ddrl9f3PF9
0Q1LQjjnIBRokEz+hQzh6C2AZHQp2IpCgVp5brD1Ti+K+rh+DNhnFpRnOzBm
FbhBqeSRXuJjFCvaMrtWXTNTix5gm5MltnGq9KaBURghsTYXacWagDrkXGis
ghaFujw/EN82gChkSmZq1NvQXdGDULsB2/poyCxrHw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MInk5Izh3TA9vvXwAqkAr2xONiQQoVCMQy6mp9PO759BHh7UarnK2a2D+GP1
JFoDGtmwwkFqipM1bsw+dG7k2yoFJv0Ka3KtMyVXQxVjvf0bNpC82fPM9JkB
YwwxKwi+0Uvr/pF6ZIfGEl+ktZjoTkrci6cgKpxjahXJJUKTvTNbkmMtJ8g2
ms5BbpoLSuFsqPMjAROXqiCBUahvxe2jdP17b+CGBhCm9P+gVDUFLtHSLij3
AqDaeO8Vz5CFxwQyYcGQnBmcU2BlDJxZC+wb47b6AFYeb20YPHXDD1K1t41S
RpcKhmO36JO/a1JyhV48h3cle3k9YodxEO06z5josg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ckwc+OCtEKoyJpNcJbQDIqLR6BcAcHGXR2BUpPdW7zAnfm9lE+qpJdCwv0fG
fUWqrqcXfVgZ1aum1XQAgwzMTA9Vscmq78gXebyhL3oqUN3Vo/pNd/dRK6zV
/uqAVVdzcciZP3MUXZw9EjLJxi/BskM8ftfGp99zJXgZjypfIn98BwIYJyWi
+YpO/VHmfN8NKiXdCO+o4DcR3XjxhRa3heRBisvspov6cyVYwTDyFOs6Gbbl
erbE5KltALIDPTxX43wkAJfETAii4lbEGoq7+aTXeRaq5sToO0UTwi7MXvGg
XNS0yQyMbH/IpefMmWl8lmRR13n7rJn3MUMl47+1mg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k5bDSK0PlWzoV8RJZaM5eJP9MMGo0ixNwgEd/ySYry7jcxPutl7EnEtUzl06
/AkQlHqO9ouDIDrTModscBkau+NVDgqMLlM4u0kaJeqv1ERXG8xVdZ+r8+TD
Tuv9jJfsNNPaZ7a0+RNvTEhJCengEpJ5msPGDjqXOz66OEWIza8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Tx/sbUlOWpz6racqKhA7mr91rHdQCVaSrQavQbdNuEsdHUAKE4UwKBRHigBX
Yxbrdntxzgrg6HQbi18LFgwR/LPGEUfcyXvZpW/2uEq6VmTimgZOl/DOg2Tc
GiR2Bn/nlFen+Qk53uxDUqKLXiR1hfaPwWd0xJEjTHR2BwxhR8LVxMWlwXq+
lxNbkc16TRZH3TqmiPJPE44+AgsYrLwVrrH2McD/jxakDTXN2gBWYOOwUhbJ
AwdFUCSdE5Dl9JZRUBJy2gtwbUXc25sd6u3NujtZVXGyqyx4/CNcmXildrr0
LnmVC7L39GKgAq+gfzJ/j0cUsF+8F6myIoEuQg2vpSvLGTG7GPnCN4joTlGq
8jdwhiLGA0mLPVrHsN7ZIu0rDCanx21QmgyYsBJ3/E5rcp+GlXTb2vlw0YeD
MgMKmcQL4rvP7lnwK12W7utMjIB8BEXsWdxmLghp+6gJksKMAto91peg213H
BUVlI2c8wz6zuQYpGlU5mj4mIayqhNqY


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A8HflW4zlOmpq83iOsLdmFQY4Gdw/kgRq55O2wIp97vY2Om/VeQ5wIfLanaZ
AQiii90oI6DDWvwr5mE2VKNQ1KdmHci3AWQGmAflBoDQTyIh1AXoJn1b4RmQ
B7XNQfw3q+twmpRATL+6CDdK0Nh2vuktUo3XnWBco63WZ4FP6D8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GSS0kSFTLNfpsRJlEzYEmfJ5tAfXTB28ri3CMvaqhV/fIIabfBdwDNl0GfbG
1d2BRI0335y6CUkq6+7x4ku9nAwrVeUHy7uSynXzPGoDp6zjOvHIGpks7Iqb
S1Yfrq7vRp/+ysbSNighOfBNGy9IDEH62R9sEOaOHtlu32zqH/0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10112)
`pragma protect data_block
Xl8E4ZqChW9m//WGWDH89rMnpwQcOHGi8Nk21F2BibNqQQ8P5QlepFqYIfZG
XeaT3rlyLlnw/J4O4BQ/XMXIZAXgCLfBtRV11Lp2BDyXWfZilTck7yCEuBWu
b9LhCTq0mXyv4lLzslc/j/z111Orsi+slEWHOjdJl9d7sBQpU0AKZgJFWT77
NwARrBhWRiaNnrFljDtuAQOkXrSpDXJieOWhF6YAUKt2Oi/PmCEmPmMruqVT
Re7FkNhPbiJWbBz9rb+peG6/h7SsBAFUSalrEQau/iuya5l+fl1fX6miTXfl
S0lbjoHUvAVUtpY+/kQzZZK2sOmb/ohrqrBd25zvqcDXe3tSLna5g7IkGMeA
elMgIKYAmKHjNcTQ9kHTrwph1+xwTWX7e2NLs30kOTjohG58a2bHYSINQjdl
Dj98dcKZ7LuD/9Ib/O/7RgzrzrK+2GhM3cOFNbSIbinFQs1NOVGzxCq9Unoz
/xO5wvj8Efr5dPVmC/Xt2q8LNgdOk4n1lU5Hb+EmrEeZ8nGO1k1xTiX1ifsf
zJST2iWJZ6hcJ9vElv/wPamComKH8sWEqNPmUtwUzRelqTHY6eBwvpzq/8m8
a/XB0rDopajl4k7bBuLiQZQR+mfvieSCDPXJ+f0qt9eYvfjSUWVB/xJp9D/t
w1H6ELtW/7gGVHkFzjTMRl3oe+Kjy05K8ihFLBPNmTaA75h3flplrWgb8nXg
zi8x4y1LyWAy5lzSjuG4TwnYNySglmIGbJ/Xwp6HVwpP6bV0qJAN5c4m2kb6
qqrDJSBHIKLwhHH+QsfRCzrMVKQ2Gg9+F/Aq7EspE1PDgSpymVdVGxdtimzE
yWKRUnc2nORGLyYY990Hm4kqO/dZ86NvlfP6M8CDhXdUPBKhQBUvHB/jmZdp
pQano0jYtxZoKJMxX65I8di6yho+ZsMuLqyldtf363Ps4biHComEZnGZzNJG
6Kzi7kqGrkDABCw34+qehrBdjeahZsCW51tToWiNcyIo84L1mv3PjTAu/WXw
V/I5CzQhd/lSBnC98XcDN1aYWil9Kr8chrKPPRHjCQPKXp7spWIafwdJJ+X2
oo8kdiaWTvhCY/Q19HgPe1jCTgzVZC3w5BApJ4lAJkIVpMVSLjg9MfJdFheB
fwOjlJY+n+AlzqpS282iwUcS9NIgOPlwRcQUx0DSqV5ubsVk43aX/dr908+n
NWgKBvsl6vpFhXu+bn0Ul0T7KhnfDpD75lxZkt/HZhg5P9sdQKqrQbVSvCly
h6RMaXnh+ibVYK9MkNXn/xwWUMOYwkKtWHnaGA706OMbKIju2h7OgBhSYVM6
UPjJO7S87DS+dWScQ0LbYU2LwciCKNvmwnCC/aHLvqOfDCuQrJZaG2BzMfro
TNMM3lsFbk/K2Jq/haD2IrIFa3EnHJznUNQOJFoSmDjib+YL9182BlrTbvLm
3eskOTlkji8/bCJK+k/swqlGawBf5/xXUIHXQ1HIk8Foo4yvLTNO/B694Is1
2HyEvBz+hpXTmmoRuswxAoOjf7nUX2X5pZmFuDTu1YPL+DRRxMT7XdytOkNW
pXHLl/331ttjVHQSluI9XBp7H/RPWNgyuVqPM9IrfPz2KKnAu+Gx0BNWJgEX
mUwVS+Xuf9dOM2tdNsBdukhyLSjakTx/cJNAMHaugnP1v88Qex9BWaw1fKTo
qc0cs5oi5zo//voMOoNNFqQFP+RM0Pl3EKdkvDhJhjWIDYk3mBbZceGkvBSz
dWFkw+GEtMny68ewZcZWlaYjQ0n5mLYR8GveYQu0169iPPwtgTBGukicqwFU
SsUc/gg5V7D50k3fOpor9TfAsuGESMZhPer2aGeLjGwuXwDPWkWK1jQA5mU8
7SmIm8ltyE2bA4T7yQEdQzNGjXoATgUNDK5tZZawlLY5iOhMWASYLOwXKc3A
m1wMGbCHPEFSRPZxuEUSAerQuSSLEEcYrVP9sFGk07SDYsj1sI0nbZNGT6D7
QCYO4TCI3qSa1E4WXAaedE3mASnSN1NVvrLo84MnH74UKBahroVd861xRWgl
/ctHLlnm8+M7VDc24YSmAJ5UNZW2u9E6FsBalP3T0OjqD5EODYHShQFu2B82
1yW8rcYQQoQKtYpqRhYGHevnpYxLp0PIJ8ic+CDTUApbyj5QFkPMrX/6ox8f
QM1obWQVA05eVqVAroTkNH0KXkD2GcfdqwwSI+NIfPX2PHl/xWVUPNYH0oNY
yXIhSDZiilrICao/1fdZU9joY13pT7FJ6P+bgH+2UY1CgPXJl59qEqsIFpPF
WkAWsnYJuSn/Je8Fz1uljV3OlbGtIQCc8E+8ey8Tc4w84LFCySNMlof3eWjS
2SmDvTjRvt5h/8hMZTPWY7G5UhkIMGJ6V+0C15g7vopocbKlUajksAERH3Vz
T0WpGX+Z06CqWA5CDmP1SRPXSEegKBarRmgCtguEHuu6j4eTzRE8dxcURaSB
w9HN5PpS1+U8Dwcg6Ewqf0h+D9UyfX3ceYR/XO5obkrM6+ukQ124mi32/e+z
Dfau5Izn1mrpsZNlgYI4Rv0eTIy+gNK8MQ+jPd10bmUAda2G9XKK3mvpRX8Q
h+AZGQwTiGJqSFVAGp7l2LB4eUI+I+Y+oLGhL/MEsn4OKeGCqWlkrOUCpGqZ
V3MnzRkg2h09k8Qg4MiDeNHcu1/bdKDgNukVvnY9K41S5zcbqQjnwek4aeuy
2GGx5zHCPhM8xMZ5BboyxssOBxA/7wjXPwAq3Apgdw/6yiYgYjLUlkzp1XWd
IbatiuTbe8W6ePkjfFNI7ZP5gAj5RARc8pz+8Cvm+YHictWbxw5SoXQpfepT
xqheogIEkZEW+4kHGezZQMbdZYjTvAmJnKEt++VPhXPwj4YoxImPpFORILhq
Aqbalw22jAQ7BQAZZ6Qdw4Ly2k75GBEw8+5NB7BaRMgwmwdVIRkfCBnujrp0
I8vwoxFwK6sjuShSpfA2UUILWvoHqOtomOjPBP3vCPd0wUf/JyJ6HD2xQE/Y
BKv6a41Z6I7boLDzP8Ts9rjESn/k2qOYVSdODpQmbO/D5lFs8BOidmkieCYW
HRnsRlrPRLamKqiIs17c921OJC8c5fb0QHB+3yfteu4aKzivgIbxdfyJ5zLU
htvaTKuLprI286LuR4oPFqEEXMZsX6Et+8C71F5StitsssEL8qlJ/ZQwFr/w
Cxf3ZHbc5eavStck0cFWQ8E2dzA+wwG70dKN4eoUM5aqSwOBdEwzmLCmIw+T
2hr9Ghax5OvtmYKdSu4X+xLXvlEfyEJ4E59xkTNfXHWN0wk6N/4EJ3clJeII
pT+Z7HZpfzzqrDTpYpbhomPmgITmycDD6ibKN1xASW26H8zOxKhZstwhVjp7
oOtEm34Xw3Abl2VzjH/9pz8HIB9YRnv/unnr/sAGuf2YSzmwJdKg4uSM+isy
l7M+V446vyhJ6I3pSgpCbynVc1wXB9FwdFg/lxuyOwtnsQJ9KQe0iiTZpomk
treEJj2z22C32U2/ZvMuzo7UYdNXvyALDxg60YX6589H+oN5TkyVVbV0wIZd
uR4LbETLWaabic4aOFHCwzN9xqm6pm4A1kQakZC7pPXXut/6/DrPzjAvJBdx
ooNTcB93lyvXChJG/rRFDhZTPQKHbEt36O6/Jn6IPk5/tNROZLBW/s/GXB8C
zv3+i2AHZRnEZXJKXLQ2H8U93ffeWXTaQ0RAuxwN2lKea2XbDP0FpyCVGx2t
6l3zMdaHPhhjdN/Yw0CMfMW3v44PXyygtCDTLBMruPghrM1uWld1hM42CVns
OBY0a+bxUdrCYwFWfqJjsPosusR5s5asiSIgAaJ0kcbxa+YNcVLJUzRXUz6E
6JwSkM06QfyyZCc4VAQMQ2gaF/pRHbGFlCpodzZPE69OBAQ+1o/8Af5dCYoV
c69sBw/34KMZOE1DjWDa0pkWl2Eisg/sHkLTgtqHYr0POD467UFq33lZ0Dm2
da6Ce29KMGzMPcu00spEIVYLmj2PIpzgafP7jwJU44Rl6LixiGNF3wP7EopF
/lbXUShz26WJd9fpQvHssQpH2bBkhrOm89Rbxy+64v6mqx5qvjjm8noeq/rl
zOET1CVj3AM4TyVZ+48tMU/m6AZXS5J+pn+CuDGTENfQGs0hLKEi1oniL0q7
/iQd9BKqsIgx+W8wlJ7vjplkQZGdLWgGY5SOzx0QWusdxMBjNwyUNgdVejVv
HvSygr7g89e2zc0blq/SbsNVpsXuPewPJaXTGQLkx3HILt2u421APiEqR+Fg
gmmIr1LZZ5uCx1nkX753RM5m4kFwFMT25BW4YgF8yfeLAxmB7Z1SzkLtXQg0
ebE9xsXBigI5FHZXnt4rpR3WZgyj8jVwHc1xkp6FwmyAhVaSq+FaBGlcEfsX
vx/Ee8hVmHVohG6P5Y8mprksiBuJNJyO0bSQ2peT4iz9fJ7dWmTeypMNcTSc
FfpOdEx2eowg/1DxtC6jjl1izxokJlFBvI+l2mUuPk8P9qNIYoSRTFUKyVjq
71+PkGSHYaYWN7OU+7Bq8EiVMBbUvjE5pORtARBeSuPE5FaXpNIUfealRNpa
M+2XFXmJ81Zmu7cheNiBy+lJREwnv6tsx6ihY4o9EdH8+oTZDWlCPUbIeFfU
pGUiRuR2OCcDoVVsmryy6LlzxZTdT5OfFqCml13tUB8oaUSPTSF5JO2/ZLqR
mFeBg1oafuR3Mrf6HnRJU9MDupddC6+2IOd/hVHsRrhXxMVRvvqIaUT3XdXg
KtHqgq7ahiDuGYdOBj9HJ1wEY9HhUSyhdfvFQ0swfQET3qRj3McdS+HmlNMu
eqgIAyoCczXNt3KgOAtovm+moWs+MlxqijXuSzRKAehQuVgNq1QegtSoC42X
OMWsZSgnvWJ3HaGtMAxd0cbnRNnBFXFERabS5I8MJNNKJNcgUM+wU9GhkqzV
lgKlXGVASrcvEgCvPa4lmkLN0ztjYNZHjLdvW1/xyAIeZI6bQLsnjXeMp2qK
znbpM333pEhDXA+qirsxyiWPCn/fBOAnYtWHOd38Xz5HYTB2knxDfcyXq6A3
PhoRst3pVx1HOz8kkOQo97uPEdcdTdkADe5MfOb+IP9ODFs95w9pw49zsQps
3yY+5ELaNoatnBlbaswlJ0e8IZsn8KkcbZqWkAU2MEUra+z+wlZsH/2xhZ1X
3DSVBqQeSIhCrZXwOs0gV8K8RmFREqnx/CxXx97hOjsPzlGQZ3/Pr7tA9OUz
odnxDK8jJtk+VKBFwDZyg/Jss65ZZw9BgpWMqSmozDRGR/1B0McEfmhMs+vc
XvsMUd+NwMGrNRMGJgqlKMxGL6FA07s2WFzgYRsCNdsXHV44zXfiCCW/qwgC
kiScqJASejfGQav8lxcVsonli9JecAKLVp/8TAqfWUS1DB1379cvxD+xl95i
OKSX9oqiNDTXjGORYW5kKSDJJ67prWH9C0s2Jc16Pc076Lx2JpBY9u8TjrCv
NltSlGizP3+372DKODNid258v0jtkSqJ0tURfpsQJuA3XlMN0YxCMAp/twkh
Lqqt4K2Ad606Ci+6cdq1CRThjpYsOqrwCpXY8lkyMSVxw004briecQEyf1jn
CCpSI2Nw/M3nyYZLRuSe0Eulgo72f0t9P7e/33FahyMhVrUufiJ3bxganAQq
nXNIzEhTJFPC8BDLmIVe3l/7u+H49r9uuQYKoushMFgoj0VQ57wyxOvH3mok
t28VyWD8Cfu0LHyER/EIisHiuL1vtcRXZKzoQ9lxOHOJwXj6eg2QGjWDlPQw
bD1ZQlZ4SB84q4keyOZfrHg9MFfbYfpUR2kpgVKhZgJPIeEGxbX2eMCpZZ3z
R0Bu0eLGAxtqV0zVmQEl9CFVMvkf0fggo2Dj/k96TOOXO/XW1rl00vpVoNYD
dOZzpS5N8q9OnVFEzPZwDBWBwI74pN1YdSgYJNAKJidtCU+lvVo7E1oH9j5A
YnQLV8AG0OLOMabip0HPsPGmZXhdwzniB7BWhwuUxkV9WPvCfLMc8XUXGtuC
slOc5X1CnwZw+1tkJpQyYMA9HnORcQAXr9J9dpIZocPIma8D830Y1pn5pl7U
ElgJiy8jMXfME9aLyO8RoFCWYtTmQMfgCH8lWt00HRNSQ10DXZ9tRX/y1o7j
n3/6NoAAK2SA5wBFCPyMERJEkkZmWvb8VoQUySwOB42MgKFfBjdEOxHScvhv
kdMUPlYV3c4ic3+DTOx6z0fwWbEppY7Vvq21Lq3Fy+Rv/uaz6M8lv3tOd4AG
Z616IIjAnKIQ2IywD+rgVfyU5nECQw4B1gH4ypJxRXCCMOxsaX2Bxbefihoa
cgMHQZ78n+z91t1NKQLO/GnMfXSU+TcX9EKVGllQGcYRRGNziGPGeiJlkJVA
rv/JG8Ao/l46c7TVi2z5LQA8dYKUtDN2u9oacBLudq/piCA3JdOYAKR3tpci
uMNGs1jSzQAGeMLRGAk8pTgdh6KncOntExVpdDs8onCtYDPv6OLHV9NLXnHD
E6iqcWlGAj05Z6MVwo0+4QShhUpv2zVHzlaRgdqoJUEAbKQLKdHI7mibbBbB
3FqttouQHKmoQHGT7v+ZWVGE+H8iEJ+qLQVg+LDavfBU12aZO0WpphbDLzlJ
4JBqIQGnPXcnG+JPMDRjQ0AHJr2lJxTO0NShgGX429zPbnlgieFdcPXuNCga
9RGR7iTpzku6MPPr9NQp3syON+JrQmCv9KBBM5WIxSCXfpjo+Etom3VjgKM4
qOsBFbwgSth/2brGn80HH5EKlsXURcIHJDZ4aXzzyCJL0AdHVYDGk2afEalX
w9OsQuIlPOnGec1FGkh2WGeWQ0MMF7N8G85ri5d1WGaU9DZM6kthg8bExV6i
YO4ZBCsPbjON5vr7J9+M5JfPBR0fJbYlpM4Z0mWWkSes34ReVYK8GhKIXh42
YlhoHs6f59Gkw+m5cfsZtvYXsfDfoZE4fxNv2rRC+4vJjTWTGwQ5xusfYt3c
4AL+YPIx/2PwURWhgxE8F+QZ6Tt130AbbpSq9QHR3Thq8N9lRxsBnS2lwZ2r
+EFDdZcwG7wqd3n0YWxDgSOoA9DYQ9aZdlUT4AFF/9sQvtgYZz+ahfYXxCuK
u27dUY86atkCc++3zR2f+K3sNapCO4Z4caUEscsVJ3PepG83JCVWBozvun9p
tujOT9gOoSn3eZqFTx6WoRRdIa/MDnu+a0wxy8a1gpOZoHDT70yYNajzsV1m
DGfb1xnyRUW0O9wE7a62X6alT1malnrsdPR9Q9S1E9j9skniMu0woaDY1FEa
K56Rp0q51nGEMGhtQL1YuE4XOcN+oSnfSVxFfi+sYzsELyRl/Cb4GUWVjxCL
BxeehXubTyKf5+BRVYMWizUT4MD7W1J15VW4Y7NI6rRK+u5K0RPlduNhZV/O
RDWfdQ9xpuycmKrtm0W82JDxx7jxXixjYx2E+JGChDSY6y2gArahZrzbcNJg
SKJiwf4jHHIUjnLUZf3UTWQ5Knp241tIndrQOjcbqGrr2SmpBTlqBTdlpUWP
ERhjHWgghy6wU6byrb7A+zgrv8Zskp/ObR5A0FsKK7CVAibMJhleHT1mcUyo
PSEAhlhNxcDWrOwL3ULhdtJLd0DA8nh6cvmRVYqsyQDI8GVVtuaMZGkcBjHP
YHE0KhVrzWP7EitNGIJMtFADX1z9rNbEYiueAPjBzLfE9VEX80YKknOVmOyW
rxKFDsQ9wMQbnGfjgpqNwQzpqJflXIqdiFaPe/FkYpOHqUAMdBcxmlE7Cy0/
nmNDbWHRycOvMhqBduWqjkYl6N1mhDz51USRfphr6KgUqWObapnv4DSEUcZA
XFe2fWGSGeT7pQTtWgMRmYGGK8h+1CK2qIV5UTYW8XQDeXSO7UhYGx3lBG91
qMTH+lYvpVMd6XZO0TNCv6eA2wv1VKE5PgAMAsMCiGrqq7n6Xi8wAcL+OtCt
7Xlt+ItmzxRZRyEJ234y20Nn3ZW0G+qEJMBkWeZfB5b5rVikZ3ASfJ/V9S0c
B4U5hxr7ziSOthTZvUDUY8RgAJlLNV5X+xNz3ygnmFoeJC0nAegnIqsON3vQ
W1mDhZCUVhUG0y/MUaMEfKoAx26KEPCjYqGuMPxNtZVk3pFHyLBOQsACRUK9
cqg49MEGtsOZaByFlUP2jSYfGyCD2ph2A3AIbSRbc6p/L+4qOg/RmOjyl+FP
QykF2oImXdn4b4fcUjOkYH6/DAcazQWyZ7QkfnD+G3uez1iSeTDTrLMIAX25
A+5IW8IBfkxxfOgF0Q6WJ2vj1aMjUpbLjVz5pS4fBVn3r0cX8IRAuGhIhZQV
ymiiRwaIHMl4r/kNfStdULgnjjDkVKJCT4gbMnwx5PhiyoBO06kbm5KhL+at
hAYPniW+XCNcMN+2w/vOIKDxO7bDmdXRjvgABgai710HVjoLio7EXVX1LBtf
TKO4f9VT4RujbUyWhPPksbMHHGJCU60j5fgqj3B+dGtmZkkhkmyq3rMtNgJK
yiVS+BxrFmFefe5o+SRrgku1VNQG7JVjNIDM2SlU9jWWp1IyPHv670i3NDys
jik1mEi7j9ztJqf0RruzxJE7EAxudTqyNPwvLFi1pXq2P/Ng8XduC45VMUpS
6oFVvUsPMFQ56/I69wqr1YvEuv7E+7dMau8XhUpmUeF9VEustCKvUKGGGBEc
ct1OEPV0zsAZMBXaxyGFv/06Jz87k50OuLypWoIHYA5Xmrj+zcrkeyZtybmL
SJGMgA2kG6jp9ZG3HytQCmf0JJ2WJHiXOxR+lwFmXVqFaSFFqO6NMk1arB3D
IUpaN+KgEHvqQZzFcWl5fB5alTAVCiqb8eDlJREvYW2ZVsJItWDheKgsoDSb
Nr9C7Cn8ZWAaJvROkDXkgabVz37FZSHHMbIXETCRZoOkshb+TVpoUxFyNMKo
ls7q0zlKYTgBes5/lIU6BXgpPP7CIGkFd3AqMKrr3i2W6gRkOvVCFabHcfbp
ppGwR8KLilNfnjzMENhAC8SPHtzNRqgTAP8IUBPZfOn6lpW3v3G3xtRc7iTX
VIJC7OLIBwbBwFzB6IxiGLS0vj9KxCJ06+ELqHzW8Lo2AIzHuy38kmLw5ud7
l8tKtVKG0xGj76kGE3u3pHi9mFaJf1E5oJe6XaAznzYuvDoHXUyMMTkDQTkJ
rFeWmx7ZjvQDQQbTdQhzHzgqIxNyf9mMAH1092SZemCXAtR2UNOzi3cOyIvC
15MPgDQ981lYkqhMyX9ifZrrdBaffCWWoSphAxLiZsIfTDCxEX2Q0jyPqyKL
rZ1GMNygxStbd4lPnkV9ewIRtS1XJAMiyzbRuAI0yOnVDyZG55+xZqjAHTyW
bQRpiQaIvjQg/pl6yRKYoblVVzcVNDHiZmadYbFiOEGodMbCawvFpl+klYxr
1XRdXjeulGb16665XHMtYAmsTIM6nOCu1SQRQ1RdZqwO5Xzx8hnTAiFLmzmz
7Av7LIx6EC4zJi8OHuxHtm1ssF4WQkwiUzZZV+esehH2wYbXhMW4qlGoBTSs
FqaQjoRWk7uhXbtwVY1gzPx2G6h40YtK2mylJoRnNj3bsuGbSCrRcuKhCFnC
buwsQQ67k9pL+D/kP4y57HvjhY4sgAQDuyHNRmEhs7IZcaewM5fvvZsdw2C0
L+KDlXUIpij2pJLs0+AWPhOhOwKZIrcxQpP/5axpTOyGXqeBYr7xS42iy7sD
ik61xV4GWsC4uVRPISyFUSReELAjWjReBefqP1Vuc2jk1wrK6Gi2QftKLfy1
I+GVgMoIZaZY/Vaq4FfXiTVE4sCjg8bFZGbRWCplF8FAUqiipHODWC/J4NRO
Is+YzWz8i0oPMhqVvkwlNnnZXmeMT+yOl+0nQ9AmU4/ZPJwG5Yp9+u2QkcHx
cq9VcXa5hc78gX0u6eOlf+CFvQE3qHqz+009twKN3Ws1ZgR6Ojksrz+/Lf0z
gNPOxHzh0o9SuSyrRRWnX85vjHUA1n73X+etex8artvv2pJ+SXitu+czmoRk
o9dPSKKJ0OWE2sev6F87AluZwlI0j7CPjB532o893qinZqszNkcEqO8SR41H
N/D1NCH0vmG293ONove0eofKysWRu7veofll/uHoayaYRIPTwh7nEjTWAVJw
RvSIk5wxhNSYr465EOrUamEMi8Jqi6g/8noLoEfzqWzJ+eknU/P8Mppo//6x
3oZrFXFVN1wZFdEG7EcViJmBN2GtGGhR5NgKg54mgsD5uwangOqdiRyo1kJf
4tfoeIT/jIyQ1Sw0IFKj92GKLVcP3mLTwWzlQg9gG8U1LUrkT/Aumt/cz5fs
7VwjcmYl6RN4Yfu5MIiBKvmUUuRObkIS16x3hFKZdQf9KFPgTGTRx8PMByqw
f67TtTumFPNa7HvOhYUyyGxlE1613AB6d5VguFyhUXLilxBif8UBARu4bYtz
BZxqq4d0bEhaaqvCxbtiiavaU/TQCNpW14arZhne6qJFx2wKJyPxtIB6MBXo
tYEn3LNNyuAQRlbC2K4FzhJMf4jJRAyCfWE9t3PCupaHC67JmJI3BRswAVLS
9/wyz09tA3whrKBjnMhABgz65Uemz74nKg3zgTymmCVMmN+DENQTU07MjiK+
YL2pqW1xEeIJWMoYSgZzzN/wGJ7SQGAey6P1IuLhyavc24wM4vPMP4Qt+0ds
7LdeRN4hhb+BwSHNM7J4Bum3GMwAuVSMKhAaosGW/Sr6pVw/er8aho+QeHNA
FC10EQqCpL2mRBYsLV0eRiXTCfx53cyhV/GidOvMro1BzZKLhk5g6VNb8g+W
IoFqjCSz8Bb/liYHOF5pL5SArK4sxaMM0ygjbu4sffBzsl/Y0jRzNmLzIRNO
beRUyg7ZO3EXhHUfifw9Baogkkr/eOLlUeY1JfyZVKAlFThxm0AzyKgJRX2/
WNddLzrmTeSyTlHmXGpR2a8IvYX2o0lL3gvMp7p3rSkONPlvhDf+y/6aHKV4
f8/lyFthrrYq9Gzy/v/BZcL4fFr5PR5aBLfC2ceJpoh94BdK9udLxpT3G0T+
Id7jkAiPREm1UPK5+sfpsKchPBpPjrQYycHCt04OSKKyIlWyJ4CVl7Fn/SnP
m8ZcEHTBP17+kXJ0wIs0bgG1e2RhT5u7WCyjeSItIwix7H3zdyrVuEkyyqYT
alh7T3j+MaDF0PgKU5499b8stjO7am0oxoKorIOE+Iyj7uKkQHF1W+MxtqNt
ATIeVrIqki/n40VX3EfB59q7eZfuuwV6uNHVsUMWvo3PxfrUlkxikPzw+tsR
QWfTrUa9d6FAmvj2hjWirJdhYzxDh2MCblu3lloKpu6n0zSdJ6L+asuGY4nh
JQJAgGTe4qxIXt00W2Hoj4U942gQERkbGNt2CmDizg4DFy7HXfwaUHFkI5Ns
nuO2MQyDeua0zNS+hbwveNOJxZrY4LKDJIVBESyMBxBbMUqGsufAgLdvayYO
wCKota34ghytLdRExEhsDQL8IZ2vZbEb2waw6PtVrUFnFld+H6ee46/BbhBO
P92gaALteMs3xbjF1EdeMyw49CJU/+7guvTgXbB6Rc2Akcv5Ot0zCNkIDPua
K/3BSonJdl/yP3gzrhfu7WFeJEUtMQr00uEq2Bg6aI9j8lJVJ8JnZjmfsM3l
W3jfSowa9MlAEpUAwoKolkfnwQ8/gB9lvUNgVTCY3WCtRjE8x3TZ7hq2r7QR
QG8EHFewhBDNrc8GghgkB4FmHYeoOdwsKG8aU7kp0HE8lFk4TyB2I+vmzhAD
99oL5+nptk1P1psAKXOC/+x/rhVt9/ICMozTMKKKEzGCgePsEiUOb2uqu6g8
n3rofVBnkjfAAmpXaKFOTPgg6/u9aPeR+s5qxgqAmtvObt2qe11U2eM7PGnt
PedbZe+lNHLE3vpnBRPnV83Opn7HizJYFh0pSUafEGiU1tBJd1tgkePcMddz
k/lCVQyaEIiRy+peMRPjKRQj92Nh5+jD5B105dGkVBosyTHCBwVLjbH205ee
uKaZD64OwZzxr9VGev1bJ+SBHPJVvvIIS92v4M89RNYzh1306VV9dDeFSUDW
sWmESRSVROe+faEehCKfwnAe5cZtZLIIsxZmBiN2iNC+HnDe46lD5SV5sGe6
3PbzpF8YmBcaO9DjYpJaLVlHTxaG6Cz41Oq8/R3b0sAdFGHTedxpKIdv7NMB
j0rx++VTv/SzGpYLZw+JHhW9gOvO8ZaRhiVAFSn+0cJFQ1EBEdEu6JiTK7nq
MaK++Gdh5382bQ/D6nqapm4nm/m03L5m00YpPBlk7RxD1gFCm6SLK+DJOBfJ
rpAeRvnongLeJUaoFQLf40v+gCMRyvX3IYvLAgAIrJOa68SxqXWarXdxgdls
rjpeMsmlEdehNuxO5mEw+0eDPg9VrajoIqyi2e1KEagx8n2tejfGQ1OY7J+E
L//R/vAD/QezP4KPJBYoJsKgqXrYGfSuF7yfxBHmUdQSmdRvCy0YZTo53af1
ONyAbAF/MCovkkhrlgGiM4K9UUzSSzNsCLvtt9G9xyllEKGOiysDi0kJp0sS
5ZcQXYhgiiqYyo8UoeV+gajPp1FZulVMZ8KyaeHS2imn/iEVX0zbaPBj2GVQ
yAAvkNYPYdX2W46srryuxBsj+Aq4QCUwdKHtjm48H6B3VfYJ3O0F7Nto/6gq
nZmMO1HS8qVb2rpCItCbm0540QhnTEuJFPZtwoEDEq6zINJ/b3KcDtojfBYp
WAStwYLSFeOlfnkEbcVvKg/HlSc7m4LKza8mNbDKShSAUe6JoY1zrGARQMw/
cCRCDPZze1Ryk79N5S6scMmcW9piu6irzFqOUnFE99scN02wHmC0e7iywPHR
lg4omRWLLtQIBYHk2AYiRpXR2LZaZY0URg/ZO+/PpOj8RoDu3kDSAyJlLvV8
8A0wHHPps7aOrgksCH4RUx+P4dPw0BMhk3/YJ1CUJxs3FQ8FQpr5fiaHAKbH
9dJVYcICG8L4KEkDbwnJtHg1iWsPN/mfAVWBEs0uncrmP/2s3CYc/DCCsJyO
1jN5e6hSy1SAHaZpWdFO898mSWVlg9iQLygL4VJ2zdlTtTXWf0M1Z6Y+OnZk
vrWF6ySosIKbvLf+bhr9CZyhzDEePElLLKcsBzjn7Y8f+ZGmkfNIfvG5NjIO
Qg3pxv88POmfpgxr9J1LXo+V0/XRtJXSazz/0nrNgW9RVYmwG5IBb5yAQXEG
odhIS4AvJAosNiChH+dAIqCFcB8AdSLOEqwP+0Sh4iRXLDuuUW3PHA+3HUEj
klhT42Ca+i8hUNETXR1KIhEZuCXuHgB6Y0Ayre0sV922PkE2rIKy5wayjD4s
UsHSPmkEqUtp5gyyzbWv4R30lxqARbPc16MVLt15hswQBYi4qoqm1DjSLq/E
GlZbq6+q8zUD9qJKIyaBvG6K3k5Eqj5ySYDgPZd62IbMKldjvmPpneSHEjeY
ZXwmAyENuUSi8nFvGDhXXEzv1mj10C7gcyLLBWto+OBLzRc7f8uOV3HxjT6h
4WViabu6x1SSFXoqrGK3OoQbQuFlUN2dteZt2QIBhN0=

`pragma protect end_protected
