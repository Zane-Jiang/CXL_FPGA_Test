// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
cxnZktVn7dwdo/fQQgUrQ2vlT3D/sDQJOjlI12RdgWZblxmT77W5L/qUiFcq9DA/
LcUGvo+FFF55XU7uZB32vksgakCmG3hZn14JvgYHg2EalimI5rTEMj7YnSoEVfp0
NgEOWyj4bh3NHpS1FOuhlnMGcIdq1xIgo4gIKArkmsU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 18624 )
`pragma protect data_block
swNkMG6ioazniQplGHTL6nXeWBSV+8HskVtaIcju2wbneu8JJPgkuB8yuLCcXBS/
tdH3mr1yNAlpA4syLdv/Qs9a2LJ144jsoVjjs3F6IWKE8egXmdVPFx6sm0naKLGc
+taFWiB9OTUqm7Nz3dvr405PpLdmP5O9hOHnpByMvTaLu1WvFuAw/zHwOETPCeUy
C09Jy96y8Yjj+iK2Nz7n9YypcPHjShnpBTItIfrVQAKoKfmjfNoEk2y9+D/C3Er5
So8Nav+6WGFrmwj577tXVMVcMuniirVq0rjbp35WhyElTydEnP595uY/eCeaEP3Q
ufGLFpooGi2tl8ixhsTb/hQimxXoxEMUk+vnMjoQptIXQgZVpk1pV3lCJNXyQdUr
PYqaxxhoUMjh/Xxh3SLPk97GUr7f7QqZD+PFA2KETvHYo6sVVcEiYfLnPCqJRTiB
dIqs9rc6tAI8hutH3WJpsi1qBgncvwIq08/1Ws7eduC0i85LTQwFjcOFHrhH3+LB
xxvUh+tFxN6nycxpoXDGCuyM28wNqDyQ2YHbAtlSe2wgInc4gWYAMRL5jYEZysSf
58eKCSJ3BG+bqT6zmROA4CVanhzS147KXxByO2QmVCB2pHooVfr0p/c0YZ0GrFx1
MmwZu8qLUOICPN9h1tugqZcPAjso3zzZurCj9clIbO9tUa4sZeYScOSFUxAyxlCT
gGv2RuvEDKQ4eT8VnB35mtvnn92MQgLWoLzK9yKEItKAiVy5d/0J1HZwVnLAu8La
xqP4E448UlM/WbTvoXvR+QBA42SryMXqeBW/ChavOmpwNdlsUilOHvkv8at3w94C
4iv9QkAVP6RIgCgE8V5FKGCXUhtQ0nAsjFDx1Y/TtOahPWTqbTBStScsOzYJH0Tc
UuDbjwR/AGXkMMe9eCcPfltDiwHU4WVxhzvdTIl3AYC5vZam4TUrsklis/Yj7Z3R
HRED8FmpoilB3p+Z80Tsap7beRlBHtenAwariFh/W3G2v93QD3yuz7pVqPlDebft
r96DxTcxB23zYCBNnqdidn2smNH2ftx77Y9e6a+tGLZr+LEa6e5anrlEf2xJNRvx
BIfVuE4CCRBDuy7Yi/neQ2Lyet3xfKsjSAGxxDCPENs/nbUPn8QrCU1CSWhvq5s2
MstdFpx2heJZ4WrrgyiF/5MWME2L84iCbQFnpDjjBUKftReK/dH1aAu5Tzw8mPq4
6XPCUMxjgUMtzVQTk8pk/FIW/NUYyz4Js8CkdzECHf6McsNq5XrPUWLSTG8MXwCk
/POYwVLPBOUPA3fBA+8/MY6SHl6VEAETGQMoWcfNPAtEftXAGCw8BHtfQfnsXonn
32mcL+QYpV/OKM95hWOUwTZmzyYoQuYrx4JdmzMY1rKEgNkr9MXZZH5sGsZ+19SL
NWkNCy31SQnVPfS/QB/SGYEtgLKD7CwTka3SgMpIqnnZfz6NXhtwd26WRkurUMuR
IF6L/fTx32JCfFioKCHRaitfwDi/VWeHZHNlywX1Wil08xSQjneliW1gmyZ7ZJkh
jZvGnexJzSqkJQKgR1b47QC0TVZr5sCweX23mzSXOhilyticv1Q0KX2j4OExB/ut
KINvPPrqfPkJvm9EY8Wug2mv7OwNruQH8vKYl62fjDhmmG5oXcimlC50OHDvx78O
5ftBGQdMA/yByZ6GrvvhlEOz27+wcySqSQBKVQNq4N64mU9nkKUlMm82AiVaDf9Q
sJum5l+02CUDOr0FnfV7SbNA7uAPBazEYtPdkuufN1cQODAA4G1qr1i/Dy8+NvQx
7N2P3wVuIli36ZN2BK+d574Jg32MgOaqYATX4p+dMNuTGI+652S+D3z4eJUZLdcT
x4EZezWsb440iLpIIYScWqmGmd2Td6xCrIx2Ixvj4ccBJPBqaxynPu8tyIi3vN2i
872C+RQWZZ5qjtoRU68hE5AtN9Dd0k/zpXXKao7iIeC3/TvRxhMWgwPCE2m1u/hX
LSM5K2J++p9iptjou3v2hf67ER9oPi1GuyB5E0wfhWpMtJcSRH35Y6V+Tg/itrCz
AqOdxB7G814qWAZsiEtW/nuH5kR/Mg8FXMakX5Wp+iGTNREUxVXxrVLdKSpvGF/U
N6EIxzDAf/H6/ilO8OdOfMA32ldGAIh6sd1O7rpqETlCYnPH13H3gymuj1eIAb7a
cR6qgdE2NJ8CbGaiFpoXtim6yq98Ir6YejaSRP9xmdtSjapd7QfQwl8XuoUPf4M5
m36Km2HvRGFmVvKWmJdyc73OxaYtXQ5x7qlC+XG7x3hOqvZfVfc6Kt9OBavNt3lg
ydAXgUtJC9ESveVoebnQV8qgcGITExp66Suw/gsyX9DGXSKTiM6g2hkKIU5/Yrs/
N12WZtkuOsIRNQb84SbOAicF2p0Gaawwa4iGPYoUB+SLV78YlrrIvl1HAucaszTX
59kDgspVLf2PyO7VUealuNfftVu9+G2EIBQ57Jl3EWBG+izuIspLboUHr5gDoLTR
wP3+rE85Y855dXDu7nDz4xTuq4VYRxT3N/5LKxvbFPOjHWvPM1ez+NZba9ShHKsA
gZaKrUj7IkCRsr6nL49PiFANRwInHOCkr0fouz3bjO5i+r3B/+8g9lCTNN7rjN2p
dgm77oU9NoVGtWyMSL1wzdajRR4j+ZlimcBbpq4r8J+MC5BJTDB9zqCb3fmEK1OU
h2fR93VTviZDNxd6svSQpyEbyoWHhR/I5Rmtmoj6+lJe8GXFEoejtV3zrmy4BVzD
57PSp794k9RiZbVYzzaVnjzkw6ZVLUugslEOsUNIT9+lN7e6OkWAxRKrWizKcl2+
4TaP0CwDVk9UrLdbG/mf/Mwpj61QX3of/gDX1HAO8uT39Hl2tho8kNeiKicJ9gD/
YGEHxcx5Q7wgwwS6X7PjDGMi5M5vztbREH+ACwuplE93AAmnyoMVr/G5+b6maXHr
rN61JI7zyMpKI6C0exDRORgGIwySouXKwPLPqxOb6iB2FIwKE74H3wgCZcAdJVjh
hWWBlgsHdH0vch5DbvQOfNpp/J/sWL6ocgbPVFA9iIb3Lt35enRu6lTIuXA7z+7q
rSqYB2Yr82i99E0NFnwgbqOtYWFzeBGeWbgYuWGnfmZbBX0yj3KN2gRzc7xTQYaI
qamUq19y2N0qmTuHS3q25HrrEOJhFEvOTIiJmnWg4IcqqJ/jkzkkNVTE0ytaSazL
5e5BxpSsNCSX1n3kJ73ltAFxB8NWFKqegxaInqYaZ87S0GsSzr2GV1LiYUAR6Goo
R1W5WdA3pIaSpMaIVr/NSDQuWncv2BIkJA/yGDqPpFDdtRfXk2mhj7yYJokfCSZp
+aYWIdcob/5G3uTR8vMnRd4hvx0ltSHGfcysVstpokFdEzVQfvsciNVLLOfjWPfk
XvmidaP0Tl6B9pKQrxaO+627GZ2tRuUm+BeDYMTyupSR/z2vWx18FB/QntlC/6Tr
RYbiZkqlHQ5Sl7xUs7jBIZXlmjUUkBRsaDW8hWCs2abOTYMjxMnjRp+AESc6A+x3
Qda8+x5NL1BpvVmJ7NUHqS9xwzlFSmXmCfZJS18C/BPS5oLdSiag1hnuq+s5P0Ud
3I72LSZ+VNY4LpHfT51SAjUxlJIsLsMs89s342fhsev9QlBa/go1FjDeLIZD3uSE
Lb+wGf6BgcS+qS0z9tuzscM21uaJyuD7Fk2ycHZ2zJbiXPeKbdS2JF7HsLtiAqpu
lSclW0Pq8wTZcF8AVE+FqHxWlugDv2samSyN8KW43KmVlPQ76hI8yXgQ0ELrM3sV
SBIhd7u/NQkN4uyfg/zg1kRaIr3k4o2B2FKibv+qo0TsftURZ+Dx5/H+rrSRtfH9
Yhfj7lg0yeion0LbmJ6yMDVDpthETgLa+jj5KhMiO6ADmnSwuC1d96l1AohxlJsU
oIX61gRNL4xgDgvroLr9HVbQlPYcX+HiC2axf0+5LEUXQsRUAHLh8ihJhVjTJkse
tNO6HJ2aQJZ8JZAbdIaL83N8sBrH7baupUSR2b+gwI5Dyw1Mq5ytVKyvJ2XInv3x
np3K8+Hv6Ck8lDBBdzL0eaRJis6QEEnIwFUdThkMtnrJrkvogptNCyMjC59ZydAm
q681w34TF4sQddFJAe/zMKcMXH9nxT+ytabCcgCzEtx8dFFs3dRCFaZMlc+eIVfp
R/Bm2WXbVK6RM9xuGJu9lBxBoGx3mz7dTOXgNoP0+J387T1raXo3o9yeWhjOvOGf
rw1y3AO14JpTtUd5C8ilaJk/SR4WVNmxk3ae1lPxDNNZCNx1a3S01xdVLS3K78rG
bDCnLuDqaAHckJcPVdt2XZFbR6HLKzk5TKIL8Urg6KlFA+1Lcg48Yiqzb5/+EB8X
ruI1bjqU3QXUeJzLn/K2Ox+L3BS6OU9pqWjVbzJLvqn1fv+h9gf5Tkvoz8w0xd9R
+BWmz1fF6ZTpO0c9ZKDwfY+hJliX8/YDjQeM+W000DXQaAUGGHqy7TYljspboAbe
fqyvp7DuznKfdvaebDOFYRa0r51DpHMWIR31LzXtaEDZJWa830f9F36J9WtD6Zvb
yZtEIL6hr97qi2C0J7C9xrrtCMsK4n+eym2OjlsZDO26t/rpxA7HLukho2Sm0i3T
7TrIS36HT5uCIFZl3gRZjTK3Iy12U9EJvCMpbTN2uTLfLv2Rd4kuzEXC3pU8Ue+P
C5aiM4IHAjbwPBGsVxhyLPhoT7769W7rU0Fpof084Qb0TVgW2QDeM6r4pEnUxFrY
SIfkJvVyXA8ziBytDnejpmLmAnWtNZjGfoHzEJM67xDrXFnn8s9lKp7YKyLZlhco
6s0qVrqtGhAPZ+M9WxjNHyQ1H9OGYdCTzp9DNCPjeo+Wp84hwl67zfglJF693CaF
IfinHQ1MalbKeSkZfFLK8CxgleDtC0K+1gOP4JjIPkc3lFN2elqAavTAJ5RyCzJK
iPWWTXDBP3Onv5HeaWq0hyxpwNfbXrHztQ8j/EFzmNKzGyJk2rK77l2m50F+SoGL
EiB0KkR+j9ubYacv/J/Of1lDNYVHpQHtXS9Rb2RpSrdPbimdamnq6Qz06VFHwYjU
7oM9zeopDju0VIhhsI/XEWGbl5Pd4rm4A+QhIwE+YVnJSLkNQezjVyFlS1cQtCmc
u73qYESy4aToUFnC+8jb9n7TF4cUPr+4bFf5rhU4j4DvLPtT0rtpMV3PlScVK1EU
NYiU/BvLsoMX3JYfIALFnYki8LdAR4QFS/C5hAjndq6The1v4FBj3S1AVJr4lul4
QG50Ofd5roW6FgVaAkPFKfAdEB8K6D+2671jXBCsW5YFpHcXrYlHuaLZarspUmkX
ScAu8siI9muH6FVnkycKxicWpvWfHDk0Mz5Rt+Aw4thgo9QZ8V1uS4gKiliAK9LQ
/N7L3jKdszDUAcmPjV1zs8mjORzq0VOBHfeQFW96wTyzGymLj7ABKVWH34KiXF+S
7aB6voyRCg/S74BYCtjfajgN6us0YbgL0mqg8+8wnqICYurnNKeTtT1TsuQ4qGDI
XakN10vY8ow85Cs2h1zOB8K5QX10kIsyRgZrUvHe/HILaxKr4MvGhwdtaM8uWHPP
2x0pSMR81QXgUfCC38+WFV7l2ky1JlCVynufqhOdbS1cpfA3PalE/wboUFXmS6tJ
jDK9kNQdO4g+HmT8JGbspV6EJjLiMp0+/cQC1cD0EgoOpzLmMsmQukAZu1mP44UG
OzdjzMWn+ygWafC6zD5vrcfmlO6etk2cCwSCx4+5Fuk0z1W1VkcoEdUZDfy3mZjD
yJgVOrlU7tYcZuX7nYGblr/7pPWG9W4T37PXfUD8iri4K8b45IZ/FU8In52y1W1s
UW51yhNbvn5K1nMTnjzfBFLDj3ndpuu/OMTUqtqG77RLYyIM/+7RJC+tRTynRkIF
m+ghBKuP+eVNmSOLL++O7gD2NWVJ0LTbpSYONTYfo+JuddcP3kjeGaxN0KnVM3E8
sHBS/V7hxf+czJ453Bpd4X9e8RXDQUB2oN7B28euMkTXuzc0sOFZTMNskmejTMFj
ctqMpwxSv962MhjTCTyjY/RSe+hBr9SUGGVSN4n2wB5VZQz5RzneD2WO4T0ttt5Y
adJQtg1fBvFJOVQ0c5+I0csznGbc24DbW3Bi+QnJ/lA8UA5YJIqnXYi49QH3Yh8t
vpgui0YPTOlfvdYWvAzoF1Ht3Rd14MyEsGG+YACO4v/tvkNBuh0Jn3Ks+UWqY9rf
qyaO1tl5J9fRFQRCz7VNrrT7BPkfomK/06W8rN0Ma2cjXS3OPVjxCApTGX9gojQY
C3NRcRxhhD6349HPd7oL+bHz+2F1yK81voi7YawSr9FLCxZw+VyobNCuVRoDWuMu
xDBm9llwgSWSRZEZ9mPsjTyW+94WKX02kDd8l1LVskDn7sT/cmmlM5D9jqueCBOB
0pG6n7fXP6uYnQfQw0h6EQd7PDIPgCJkBh87pKjpZS1t7LUCmOCNRAI3HVKa3Yjx
++G7oHDOfQh4bvbuibpoB0a7JT27IiKBKlahUSKBS++uDdjGl9aaSxliZ/QesZN6
XmE/DN+X99KveisW+VjWAH53FmKLVPbzWDnyciJr2t46NE/fwBwNn/MQu2uZXUaG
OwqLDlUZ82yJ/xkKho5UXcIpZPulD/9GVHEDT9wpWrva00vyHjLmxQ3ShT4QBb/+
16F3NM99nI1/ouFEB2JGQhkT6Tam5dPa5l1ar8p5dRdKEk8bjK1pMWJmIyZ6ymf/
X4lO2rhTtvFzpy/6CMULM7Fj8FZpUQ7hQfZWROtclzLlF9Len4wwQV6jwNOrLa7V
HvQ/xaz31Wgu9Ts9Genohc5Vk2qcK3umTzUTdTFdQed6QKAe4gu/i/fQlcLHznKi
EoJGioJqwLk0AJbU34eoPOaF+En4V3AyoEW/r10LXXeEDgYg4JgfAAjMpV4vkX9/
Vv8LJ7QHU/U1d4wGmaB7QL2Bc7EpbO8DeaZCr8rd+j2lBRYFxWBpl7YTH33S9rbD
U20PuHlH4fXhaKwFyk3f7PIYg7utPt1hEodTQrOSJnKUBGBS/t7wucfrZW/VIWlJ
yhI4nGiu82NbBFKuDXJWiVEw0K0YoiU4h0G78Jdr9+A1ZpbP8ZrSVLeXMW0uI1JL
MDtBDsSeHlp73wlFKqxBXpKkOO968oamHwvK0N4h1luF61cIkZUpKf0PkLyAwcH+
7l5kn7batXJTJj16u2Ve2rJuDc4nrHPqBa39LBM6rWb3Q6GeVA523lUARlZaWzSW
E9Y+//52/aT/pjC31TXjLRFOfzYCZPHDKlfxl6/QUukqB986Yyzsfy1rStyb7E8c
Xom2JiZSM/U2iUpFM1oLkPDPCKL3JZqdM5E2+CfJti3p+gHvpPDLVWuL6qwNNP2V
6IVeheMrbH0BMuz+m2jLZs/fQCoX3oalLF6NQ2Fkb1/7KMkd1HrGFMcvdB0zkYrz
XQsLXpQBjZJ66qyTF/iKq4IHtMlFrvkUAHbyIL1PeBxQpJql/oAZQiTonGacf7Co
tLj0eNpR8pUlix0jhkZnxYHc/jfCEz2yblPE9pR5w/ocEAYh1oV/vHZ/2beb78l6
h8hKDH/wR+M3yr0bdiBIV47rJGDgoSILKeLguBy5o2Kx5H4bUvex95OQREi3siqC
5mxlazXEf2AsV/AdB+jiwJJvU/BhCOAw8qs9pkk+RQh+9pzJ9PnwanicSD9RO9eM
7ummtQpVYA3IrkqqIYXy17m0H0GmV0B9VDWq1NYTFvokZebo+NToHAEbz6m9PCee
eUfPFldp11tXMejOJAky19TXV5ZQdA8jgQV9VkWzTIb3UuOkVjah3+KQkTAmr4A1
jUn1Wuy6KENyjGbTf9Xy/hcojIS7lSzNy/DrAev4qy8IENMnAX6/IFfYnwU+P9Tu
2rLOxxc9fuRzDhyGPt5eO11AYDTuA7UzqdLDeZ/z5Rs079dzZnhpsF1FFgT80Q4x
yd9EYNiYZWS0dfG/9w5GOzdiyWYdVvnLwm6BNjfz6w/RN4Sm1ywCyITnbGuH4/OO
ZoK5KoPqQwqpLUj7ta7j8SHgo+91Dt3RU5YjJvXjCYBsqlloLDyM3Mzf0GR8y5z8
UNBQt08aUz+neKjDaZhtP8pK4NPyz63vdyBQW/XGKOi95HS9tFErBHkX/gDFLvhX
8Qdnpntc3oUnuMOBs2DA32nBSHoVE4gzuaxDR55gaEyKoRYu58WEumiakiEpdkfL
CZ117712TOpm0LR7TsDtHbYBNZESsyXz41pKjkPPpV15n5bNiqhlDVvmScaU2DU3
iOIsaWtikrsZzbMLTWV9ZIjR+KdV3ThN3MFENzhiktoiWNq7RZTBnai3z4XVuR9G
bcPi0ffcQzUPwKm2JhMWgifl67IDvw/plhem5eU2wjf6rLz8Yz5RJQkMFp+o31FO
V6ixILQc/mjqQYYMhGkbK560OVGHdYPUe590eqoD+HCrTZlK0qPy+trJdBhKIk94
ErRRhGl3WgLop1Ig95sS78vLFyzjxaul9/aHdzlb1vicS2PB1NhGG4y1i6Y2mD3h
t44kkoMS8yhBdP8tAiTqSz1gdILdL1Je9mz45CP1ErHtBLDx9xVia6LE+6GXbrUf
9WdQQuWogdHwTOIADNwz4pzk0jflkIzPevFdoRp6ZGT3qJn9wim1eursDi+iso1G
1fEJyV5aPYvd+vKBbq6YC45V5OSc6qH55F1y8HOeSkMifpZQsp7bT5kpGLtbPP1b
u6B6I5AOUil8X5Qqen+gciM95CVZDSXbqA4JbJoLMIVBy5SXAE1Lwq5vzuzuMQC2
xTGX7sGNSux9weVH1ZEtpsIBKOME0nHmzbySbRiNoeFkvcGzjcFrFCPluhi0SD8f
ll8NLIQ2LkqCy0gvYXBBxAVRaj1u2KCdYQ5po5T2PFB2E6Ah6x1jHiHWlj0u9LRG
cT2OKgW2pWxQrUtBbQoOF4S/p/Hr/rtzc0RfiFwdUYXxvDhA4W9qqhPeD9uOVVa1
pIJo2rgYFxDjVP/sITP4WiZgJpixTrkCEtcsEqSHngjC9AN6fhPP7cSyPyWx2XgV
yaUwURxCgTC3XKp97DHMXZv0Ga4Je/Zii7lsCl3JQ4oIs+b6ZyLkNhqYHI1XxMRM
WVlOaL2QhjKReqPBJtphqOUvzJX7I5MUsXpOom9Sa6B0SQPARLF+rvctVWrHCqoO
aHyeFD7ud9QC+b5CThd0FKZCY6dRYuwZz306ZO6ZMeGKS/NIPRdwTifaGytsl25i
AwJ3DaJOb7vB1q01e7sds9jZ7ooYlTgW99jwWGd53tErCf6DCUDQIclRuMDECwea
X46skOL56p1/lg+KnKS6VNXthw8t9DGLHI7tdSUQUyrk6I+fDHtUiGZ7jcUHGc0K
aoNGZphphSdalIG6lJE122gmz5s1MYUzGxcls8FAhszbEshMV9+w73ZPamvCddBc
IB68bCMSVzDVT7nk22uiaWD34W0Gk/ouyxgWjHfc9RGaYopM39x+lfJE1++BJhZ4
taq+gyluWapdOesvnILDpr9oC+rDhAzYoKHQQ5S1IK6qeLlYe8i+dO/d7FsS7CcB
R8KNBEM8pYsbEduKE/eq9koqU8hRJYXJQz9fhCbQRpKMHotEOV3SiZcYx44qamjq
GBD1T0X2ZZmWEOP7cQQXaLxRzCcC2/0dt3sBj84BcakExu2++UarLRwshPxrTYGv
SAv6OiSCUIWld5bJhfxKc0xjN1f5MUUrslF2B8J4kPPkYdLBiwMLAwLCOwRmbHf3
HhUFEameV+2oSCxAA4avP75BxbEL0Hjnv8O2peAUPqmxzfapfKfqbaruXjFgHS3d
7FOiSIO2v0jDUdP1g2te4iqnW/jFhokIZxu0CJzXN5IkECJ5mK4dDhCJdpFFpp6b
QdygGPACjUHvgQevIp+/A2JT6W9xcKfR6j6OJ266xKNtVlCKf076mdQ/gQFvZSjS
WNj/JvniFFjHyc4GkJk+hkZsBTxl9j8hTh3ef+owmWrdoYcFkdo2MoW+h/kggBsa
jCaCaj7D3SLIvGTGPhYLOevpRtO8fnhSBbzZNsDctgU2KtSdBT8PnZ8aGuMAD/Z0
XTB8rAFcPxC1Rihiey2CmCQTi7kgCpJZ2l8G62NYkLFSxt9ZBvmqz+C1sIQocfNo
YegWmYfKqcbxtj0K4yZHq4c2kqCuo/W/JYwL014lVbR3sGFmj9AmGhIhUac+hLGa
Uyx6n2Yt0/DcY/8WkAf+Uw2/fdrAlQEfROeqm3S4PRuGP/1BvTYfH4YpAmRzCe/Y
LWNtqCojriG+kJgbyStsQGyCdQVf+hqO1DB4iQYTaAYSToFi4nT0ovXgyyeaFO1g
2ymQujAyd3+yXs2bp7V29rDhCbrYiTyoMifP7h0zxqzMnmqfqmjw98K3I55OFTWc
S0RXOPA5pyLeMlultFgK1Z73eqQoLDS8bWoesjb5g5Nwp/qQShTq8xyeBAkdRLxw
O+kPbGXqXTeb5dtFaLcLtuhRSXkghgz68mM8Mz9PvyYKaS//8NqUKnFZ/Fay9N3Y
LF2OMB6FHdoz+xkbvV5kbotKlvScv8ZMBbh9SyqpoRTptNdwYa4FTraVjvZ980EQ
gowpUfNwMLvwoK7Kve7D7vEdmAp7VpP3HOIVZRRWv394lpazneHxmCroVK95cewi
fKmQeo9RrO0iccLAQ36FoDkffBAdzz7/3sDW8UlSqy83FDQDIGBXHCrBObavplLb
bpwBHZrPG30zzNrWG4poRGTPzKZ3GnyJu6x0IsqrIHS/gVTAMVS1rAIO4YKP/h4h
R3UOgOE6+iEiXmYOvuOIW/xiteDBSTipy8Wdx7LKc6uDn3/tgaAPEthA6b82eH3y
tzEtN5Ff+kF0r1ZyOpjIYfP8j6TiUS7RY6nhNwICr4NOd5y322upeWeW2Iu0eV9y
YiC0gYv/ul3u6V+qj+qjMDHmiuK1piptdAO5CoJ1MqHX9RqwWqmdLs8zvfEdwlGX
9xYYj+MaTMi1gQmzzivzXWiI6WaRjIkcQ4L1+Z27GiyGsPGRxVMuRIdAipVTnYOu
I9vDIMaJ4qmv6V94k9P8fQRqzRZxu8aLAoECYiXa95koNRzUpe8X2fWi+l9TH74z
A7E1RjKjaNV8ZPCu+qY0/llUA2yvq6Hhed+8giAVXSPkznG5r+NvyGz+W1ivMwAW
fHVo6/9Oy/Soa24mwz9mOkrNkW1mR/FTOmokTgR6rkQK3Clspy3VTRQjOyl/Xv+8
Ahl185/pc4MNGiQUxq/UFe0XuCyZEkgY6DsaMPndoYFA18kXhYYuHEAa+Vh20gWz
V3U8hnek29rv+endAs1pVpST+o6m8Bropy81TbiL8J9oLktYD38xNHEcHjg1CO6M
wkiIVJSXf1zEg0eAPxNnK2o34iYslHdFj1QAiTDFbMjNEcdfOCq2+vk+XQ7RBzvi
x/KUfozfI4qxPUG2c811VmrXgn/0sTjxyhb5soF/izf7TRDfo+ofo2fN/4f1WoeG
/K8AhM84iNl7typ3p8cHiXjZGSCiHzPK3K237VIHbcG3Pp11k2WIaUeBxTp5me8c
r8X2muLyiter3oL/0OPvFwOdsUGYYoWOGTV6ZFD+974q0OKoUI3cHxL4Nn1SCcqb
NoF8GaM0abYJFOhPIymTcC+D5kDcdQPdyZUpaK04v0X6hOfo/yx+wpTjjCmGJQKd
Ax5g/2elAHfs/jx8iqW82VfcaWxgmnfGx8idZudjaG1DVxHOStLf88MTglKKTfv0
kLkSd+u2OJeVZZwsu+niz5I3B6k1CokmysJohQ+J00tGBw4qbeRUUtoDP9JAXcRb
YB2CccR1u9MXWN3TVZG27+o4zCDLanOpJDnQv5iYvLx1iOu0kt2CGVP6BOVeKMfX
Tb2x+l06YMasvPg+2ykTVyl9zoUL9DM525b91OFNB6C8dTfdht+C/RSd7xYCyfPy
3uPFbq+KipSc74kuvMc5+CEP1OMVEbKmvIEsKSBp+gvH1ZjuGtXzb2TLWmyFDwvw
KDJsudUTGJZFPFmGpdUtf9hZHGZB5+25gTVkvTesACxuK0gbemD9aLqPi60bzNzL
RnaZ/VRSoWjEWXLbczC5DOFhlKxztn6DIsvxHG3QhxAx2kNiy8Iz7vs57zq7iBXH
r0fONBcB/GkkeAAOnPgxBlYeTcK9uVdL/0QBExTpasDbERgGPPeKLuVshl+3jcWU
GsxZDzRhlQ1Crcz8MSFYLkJEnJlDUvVhjvVJhJLCaTTFMq+f/cM2TUGEjuCvycZ+
o+qopCMFh5DbVbbzXaXfxZnOWkOUb1yLgXcdWhbi1EBTRU8j6OXdiIiTeO3/GWho
K+IHeI2WK4KbeuJc/ij+fIpmnHjdpcuCYIP1QRBspBMpmU7OhML3Y3EUjb0I+HCi
y31rNNOSbK4GcCAa9y8+A0x2zYJ+RZTtTZg3dKQeWg0dV7acXHVVdOsspUQOYSoF
oIn6nhNMS8qL4EchfTeSXNoHNEdsaYJEyszZ1d7R5sgTU4RC0I/S0Rww5mPCTR5F
LcXXBUQ5aAT12EjFzmxcjgWw4y3i6NU+cPn11j889Tg9rrfJlxJ4M0lfr2GEI3OM
mtiW2UuGgMdrG0pVRO3B9Nz2sotbfET6pNhDRSE1PSDdfIQ8K3osOYbr1Epkxj03
Yg33ERP0WxWHlNQhTsOXyNIf6M1SX/JyRinrhjcdUc6WfsSK7nsWdJ0ufdqLFBYD
DHX/JV+yww5fkLl/cnRNIWaECz0VK49QrVF559J4cKhaji9DmzNBXhquOszaO45Z
w85betGxJQW64HI3dfoTGjwHEq3zjI6K2w3ihbh5KJ+2ijH0+7ZHK6qfB6ySbHIN
vAqAC2fo1SfFBA544haMqO7N9QSEiVqvLT+fmhlhgXFNjXmjFlUh09NlMDfioG51
Ic5SMhsdSaKLmtIJNvqNm/ch7HEDjmDK+sEDwP522DMe0NKhp04odFBTNoOK00DU
6MAV3F+sYegYMR0j42gHKlpoY64og9URgNkehKbV3okPnLXVcvcjmFlb0ufDMl1C
R33TuyrTgi3efoqdqBAxFess3HpPyEhvdd+2kQPUCVa5fyPaQsjGdViXEdOxjGhv
Y1/EzPgsSyVKPgfFjy2gJBw/rkW8Q/fXwNEDJ1BjdUqFQyMbxbIQgEypPbwIMssy
cfzM9R3Yrxf+nWpIHfHixYqfrr3JvNY4wvRriBblyk6I7rZmwApBPSm6JJVunErE
1hMYnwm6eDY7DGUATx1FpZ5mecmjP9JJ10+Dwq1eO6iIHMhXJ4sI5QDAR42FupJh
ygc3TRXArPOBRarXp56osRRLKfxpY0VhR7K9AZN84VzX7INtacAwjXdV8/rNQ76/
YPR3lyY0yjKCz8fK6+MB+i1IcOYxkYCw80EsFVNNeDFE2QbT7wexcetsBo0oqf6g
iitDtDYA5/jIuKvVclWk8l2tzcTusKGvd+vg4VWkuXG/qtwoLvm9nTZmamixvWw/
ihjHET9+kTDRCKoCnoYpAIMrlPZTv4eU0wFUPho9aU2xkZnLVPoKfWNED/P4Qr46
/4cu/5j3ljSvurRp0pJIxIfvZUtYV1ZcjD1E1tu4rv/+I0Ev0wPODjP32PAmzC5y
f/mAFuMG2wTDdA9eJzv8mhzjDmAOFgrdOXd1zQA2FieleTIWzqRxkGDAKIDrAWu9
deZzXwi6iRqiq3tRNH37YevQBhRGWgUFM208T5J01yAYmxzRrB4YtQXGdH7/icsX
8ZXJDS9XYlGXuhMuL2wlE7MivzN9o3yayIuVVUhMzlDKVydfhXsdruUhKSfXSN86
EHNKjF9K3WUoOmm0UUJwwarVa7EZsogDRc368TSXmtt8hjOJiLbCbRybvAC4JEN1
3rtvs1dNWWxhrbMV5DgQdP7hcar3C8c1qrmwHP2yOH91NaWcY73Su4DlByzhdqSN
UKJHDE8P8E3bvVH3N3W7bPAvALcUUI2p+kwlw/IQnzuLDBbQ6k6va/+gkgJqF4Ii
JF4ZXAj4GoyytYPHNsDEGNIPZQoxoj8ChFqVzz5b9/LMUcO1qWoh9a94+kmbeVmA
sjw7kb5Gx9fzwioE4IgPHAaxxQ6bPHfTWfIvH+Rj7XSMh+GsSDRMvMXHWU4b7HD5
LUKsJGYMZg8lJDkHPKOcn3XMpTwvUtzdVmoAN5oqf9QBDDniJbcuskQ56SRf2h5e
xmTrx0J8QNMqtED3eJQdMaCQHZFIt7AN+dOfwJzNJDGz+1abMryyo4aZAQAXDA9Q
ih9rMPiCtfl2P3b36qXy+qtNYQA6xQauDQLGhR65xyfdQM9OPD3QZjhBWhFKToVi
cn7AQv/F7uO9Tk+r4S88h5uXXiIRY8NplJVSXJLKzj/A9Bg3+CzeAqkS4dHfWuFh
TcCswDBJ+KG2QPinWlDmkDcwTZp1Pn7c/7PLRvL399umaR374ZZGI3zPAYTpyyxA
yg/sFPL7O01YjE9+1vTF2llcQ87P+rmI2t+k2E57y1K7DQDm3Ru+q4MpoYJzA6u0
5s1Hoylbv64yZRDKP5Bp041vuFibEVntg9Z9Cn/E7sT+PT3lFyRZUNFXrkqHwJu+
9Gzpo3ZHrZxaPIX/C8ldqEf5ljf/tx08GmQdgnjcDHNJT0nGvKB/uljJYa2PVAZy
2kXsPfwDToKY28oy0ziIRahq1bsd0o51T2Pep4MYJffjL9Epx7LwfeD0ooRZwOJY
2mG4oJFr9uo9uFqSgWAhP5VMra0AeiDg35dxD09hpH1Xv/4Zb+jb+WreMOwL9E3s
wHoxJrCwDwSdd3S2IvfWzFxKJSB5Qct1IJkelHsLt+CVWXFDn8ibhksJ4/LRI0cH
LRWfP2Bym261ITaAAWHXLvSpR+29qZrJ2iN4uZA1Cam2H+nu29zaT9au/YZvuKWL
MZg+0+FFX/oxmtPu8sh63azstaZvC2aGssUmYASvZIfuwxEOcFr6JwCwAipVfgPR
7PyZ7PzFWjHKyt3ELQVzUb5hkpRPQ9cBEt9n6iW9Os5ynUC0AXRrCdf0We2TcBzr
7SQ6FWGo99TY0YUc0Mu/GIWJ3YbOznFBJLzcgn7ywdvTqpXy8r3sRLouQlByRUs8
+kbp/1E2RFbiJCjafhdJpHvUfy86nTp6pzBEGyxOuFRM8cStfj4RZKdYKy2ARbln
izk1ud4RvkPq0THjh/slGBVcKol/0oyq9etK3KsgyRkCPUAAy7F7ltaVAEhUQJSs
BR8OXWTDHf4hkScSVfZOfLrb65IsPGoQUhIE1ctGo+OK3kR4B7Y/YeKD515MBaBX
88XYZFBTKz+99bxaxixZ4AXxCKbkUg32CnikycvyeQtBNWbTUJclYwrDoEZpPgJ9
hH6Ug31M2wkC7ZxAX36gLXRxexks8iQ2iBGo7YBwXU18FXi5hXorGcphjyHqRlkA
odceTpYeayDnfKUGvxojgJy7YCHNdnd82c323lOPtOCLQNnjT70vWHC1e7PNEf2c
jk6LNtmCNEuisHuFrIj4R2LDk26T1J3zlmdZjaiAmZtOIEofHOqMrBKTGBiA4Vi0
BVJDRIHF9T/gDX/BJ4XaK5dLtcyyAlIbp4VhxQRuiIKgQzyb+M22+f2tid3gJGe0
2z/IEWoG78PSewYR7ACEiHDiSw0z+plzYh3I78c7NTF3CMEG5DD6LTlEeLpegE/b
cjYH04eYGN4gbfP9throl+b+4e0BwM0BG6oN267TTXzSJvaUs74+SuqP26vVirj9
wDC6yYFIZZs9qtaiR/BfcIvWU9TR1PMieKA9JPSFFbjrhLOGwFklW4wl9iWs/vW8
x2JAAYnOivcQQpHTArSp2mYvB6gojXhAZmjVVOpoKUuis89j0dMKNTMd3y+XWiQb
jiVnChUsd8fo8ZqkrWlUbyh4EyLh6Yz0ouc22bIWVL0tgZSbgISNOrqO7rmKuV6G
z6G8Al9SUK/8Zu39houx4deBXIPD1fssteupiKvntaWKvV+Z04+xoG+sYCmJWxN5
O4rKMhmgA+wOaitqtkomgsX69NqbVLz0Xac4U5RDBWiZwu7IeSF7or+kjH9DWPeJ
BKvOtbrtcdQPy7aZtSTMo7IXXXmaK27t6fmhypwjRu8JLvVuDmZJ04SvGkE/brd1
+2g58skgcUT+q1e5XZydLskAjRe3b+qO7zUX6N7ECVt499fm4ZgO0nLXPVI+gpkf
dAgnKkO/WzMDydx2fbM6DorxsjHY32XeaX6kilD90vWUsjP18X8Eb8FbLBG5zDrq
pAl05pGXPcLnRIE8lzCXDl8+n5feYBnAi2zGJsqS+5ZGy+fJ8umrTFtYEVoJ5dZN
kW0z+kL0mxYYdTG3RuonNuJQbq69XPU12cQW1LkSdROUjtD097zPiK/gM+4PMjvb
rOpYfQ2VdbOgD1O8hf/a/xdn9r6HF5ZERenytDaOk/hMu4F209rydZiQWHAjfan9
cgcMgd5wnwaXvlaTbKMmBwjlsSGrnKDnHyQEYgJLuualJYL0ag8PwcvBt7oVmCC+
8IUs5bDteM/eJ5laafDOoN2YQ5QAWLwrt9cW+TMNZx9c7ESOZpT26HxLxFpurcER
kp494i/oFuziwOmfmkwjaWfAFZR+7fSevuOmhZlo3DNWC3Sh7h5ZWHU2TPnwQ+Uy
PnjzBYdHhsl/Ego3dXA/igrp9DK2KuBwpAgBWik6Fp8nf7d/PYXwgGDIoLXxQ6Yj
nwgy3+aXYCVdrF6aGmYPwr6Q0sH2Aj2e1DF7hpmAmTJ9ID4KaoBhi0vqLOtcHVnt
UuKGey5Bb01SSQfuaicqiutv2Ih/TSeF69uKWgX68369Lex9d0uTd4WtK/a18ix+
HFGsR4GtNCc9RYCz0VJVF+TEFf8hV3mTP1msVDizRKRpIRI7vHSW0QUusAPPD7s9
0J7ENsq2XGwIBL+68uxKA5hi5dIMsXXDxqcjAy69dDJT2reLzoESVwZRA9iOGCTC
gW35CTOYy9Er5p5bnHQN0PTje7s8gaIQdEIA0R36kST/WCj8pSddEjxVkDs6OrBo
pXCSb5/pN1KmCqQADBh7+vpZbKYT/L4gQdYdsHRugwsr1jDIzgaLR5cz7eh0PKMx
vyIp5TiVSaaWFZmRJUn3Ri7ipuc90eXPaL++huaGZY7Bohrftzk1hRqLKs6x2a5E
QNcNFPir7zb2P4WSAH/uV/pejzjC1WV66N6huC56jChzfdpMuwG4y6WRsLzzx5oq
d79x+9u4+/NtX+ZcFVwe/KvdVC5uvX16i5DV0lttWz6uVN+x9YjWGvqWpZJAfR0L
nUcmx5x/MH2QjnJtbkGwYXEM7lbd0SAyz7ucNxEnEq6e4P+rV8UcXOLCmvDWXgjD
UqiS8KcGchf7B3l2setUien3Vwa9YvTKNxw0Z4/N/wTW85oAqG8KBrNrrVCzodY0
+w+ahPG9AFs8/iRvXxrbhrMqNDCciVW2359bk+rerVel71zqbpmDwNhNtqd44+YU
oYcqiXl+9hk9HG4X1U6Ern86UK8FB/PhAcBY6yWb1wXYU1Dh2OlY6yfN1qYsGn74
7xWW0sSPQlwBtxEtwo2vOYIsiuDXGESVvPxXLcJGB4gyQvEHLNJGVIOWoBFCAubt
pfVJ9N9TKXsAtshpp8AnZyegOFsZKN1w1x02KRNQc71YMxxdbMCN3PjeJjUmLnIQ
V32mS+XG3SlSl7XItC3qPN4zCtSXz3HoEJdA+vI9g2Dr6CbeIxX5ucCA7IefgH2t
Ka69VFlwwrv65nim90Q1FCSjUcwmEi/KFUZOnU4MwSXgjyNFF3TIhRsdG2cCuawA
v9GqtBh1B/pahalMQOEqh8jbJi1OHdwmRQm2vfr48J57Y6L+2j56mpDIxJhshMry
z6cMijW+hIIBckQhsSC/hofyrfuTFAKCQudWEzBD1UEnFmSNRVkhD6ir1hkrpkFe
2dWjrSYqszD/gDt8HaNwE84qjRKw0paC78aCSWVslZ5g5TxA6k84reGrQUUI8ehU
1PN2DbOxXrqvFbqsrlFFkWETYslBSf+ERl1Td2me14Jt2PKhnHNB8/mCohcFt7Mc
WytgLf7gKwuSE7RJDGBn0tH6UxbfmmzfWFCp2khQOI5nvvMcrg6GSRjaVMRhXMVl
RoiNsDJGcUEfC8ZdgPQtDeKIZLw4LEyj24u9XZKfwk6MhBFuz1oUKEQ8h2UWSnB9
B6lH6GpQATHfmpOsQPqlIzjv3RQ2XeoflPqXrJ0OJb3QjCtjiUTlioxaqhGmesHL
QLnDjyYhtez6UDfHnimFth1dpf1T5SzLYFubArODYLGQIg7+al7sehbObHFjvdU0
FKnnJGw76LvZa2s4eKfk3pVMCZO//ITib50X5gGM8JrbQAW/FxuR3NK/1A/de4rp
WW8YucAuS5GcLNf/KpFnAwhTPyTXcVnZ5xUN9Xv1EORpmuFfjJDqle34T1ymsn4W
UI3edWEhWABw/9dVG+CZuOQfxGxYASvrQNKK6QSfVfJLhAyV8PntqG+1VaDzDbf7
E2yWPbSSrwUKr9yZOXikRQ09EI9L41PGSB/8itDMSwDNqhhHFTwVTSfU/mJ5amZ3
IesyjVJn6STckv9HYnf4aUB5Sp6XHtQMR5/xLVPOM+o8jz0As1++o1TgiaOuiGBz
oGVae/iw+EjWzWQ/ieDt5wVmMOv0lNPje+m0sdD2eh7GZrQhrkiqKT/dgE6nkyxX
ZgKqhMR73sWz9Z6pGO/auIKcQKzTG3g0B7sNwN45EyWm5qdJ9M5rfRgKvhA4A9pv
qgO/8hTNpXZz5HsM0wZlHMTHk4zknDtoGXdhz3eaYIg1i2tOY4JfD6VQmZpLTWEI
zBqern0Po0O5MMCXOw8tG+VJ09cx13IWE4EY0dsmTGHMqdz4naNL21Gw+RmxLVzO
J3twpdHIgFYn8SobIksOqUtVqzCYpUksiK7N0YUhr5hGMHKVcVburCvSZ4ktAKry
KxH9VAPU7hEZeF0BLR8gdgh2oNqaeotYC4/QgCd4sCeCJKm0ezYwoQih1i5L/nB6
sSMBDuS/GJUQfbhNSnEsm5fPLK0UPARuPxJXcPGquo8iX/23fP5dMaaP/TTCkPe6
8ntypHMxwLGk+wmYURVdQgYtFr274sfQsgi7qlFN95NOzuFakCizNWnxatyuvvvQ
bbvlmNVAFBjqCsGAoto8SB8DFdTptVAiHaQWov7lR/8Prf/HpA0SjufID6/S+S1E
qNUy1/x2IVp/30ECKq3xZONbfUT5iaT4TrIym6k51LMRUfI6/p3I+VAFhAjhxXBg
gN3e4gWmKkTQocYHSg5VQG4hs8SjG2mtHBUzNFYZJv7em9hnoUpKr9M7KrkTxmKR
L2Xv+C0MxNZtQZcJakv4N8JUs+sDHFqNsWt+0blwgiWX7SqNMd77sjwZD+zM6D5L
RWC6ZPNhvp0b8dNXG6qrBog5x6l6W5JmK1kDVX7YBWsZ9mGH3f8iCvPWgmCYBUaH
gw7HQnmnMcWhoc5km70xXk569aIEgWMQYiHTinnVGrZRYCkehrsxZsIn4MTw0w1u
tPZxqY0ZkOTm8XbiYHe3QZT9c2Ewb9uXh9wUT7yK7vHNLZeG8RkISFpata4MkLa6
FRn6C3zi6HB3TRGu8ZNDOcjXHX97uN9/LC2YZNSXdZvOsO1O8cFoBw5dYSzbqS/n
0Mr7H8mkPYlixYJht0EH60isaciAvtWpo+EVKceBjsiKAD/8lUhfsgLjacLV7CYd
XsjXHvoyNYT3mDfHJ22NhAWRvvU2n8gBRQqE0Q05lfw9TKZOX6k+rM5fTxIJkD7J
wel3dvVTdzyv3R6Ch3PY85mWkIEMTw1WnkPan2I/P16vDxmR2UP99NObft6ZaPwQ
8OhM0vPHTTrH8ikbY2zzOyWkIi9gYXGZUl0Osoi0fbRo//baQ03MvBfXLcCn8kD2
HO2J46kKGM4UoCSUVsI49VhkxVR7t3MMFV/fS9aR+m//jz6Kj97BcW0TTB3CVt6Y
Igu5o6jsQUZRTG49XFX67ScXN8Ji98/2WkRI/9sUfEmAk/VY2uKKGQfs7qNWHbWy
LsJHHYCQcr/ECWB2cuEp7YeJ6XfY1i/zsRdS7rOepKm/O9K+LrZf41z2E+6qG7of
YARx1VUkv0bdWTuiodjlGdQ9Qy6COltGCJxQp5rPlSQVQssI6kZpxjRimy/f4Kmw
3ESA5GMAt02vJSqJaRt7H9n6nm3ACTVREf03OuTCgnAvexfCTLq1BMmXR55zAeJn
Loxqpm8FwHK9salel0zDSHvp7Y/P1+KcpquthMXFqADhe52j314jdQFphAGlUJWk
wFb7SFU6qL+nNhBLIuyOM8ZiXCSUfLm3I4XwB5fGL8it3+hjcroOS/znoeJzOWvx
lLwNSIEC7HIxmAphpnesRyEnwNHmYHprsc3IXNeg3H8HUodHPGXmxUXCNr6gas+9
FkpIfqPvU35/91dOJqscMtCzFI9rH76a5OZsQ3nmUHIWHw/V/cFVtHDa5tD3vu1j
xvu6FPSvPhIptGw8MPnCg7hVIPQXuAL/rbhdVVCRXEv+N0dUgG8jddO11EcNV7oh
SrPvwhGlwoZDrt5yH78lv8NyZqmSTCIDAS97eftYBA7OMYOCj4geZUaFPuMlkcuG
yYlCZOb9BvIYDriAuBvoTudpDIjoF+EFXk9gxzSzcbIiw8QZh1TGwJI6jKo75001
WtF42s9N7czBf4LUniELlpggKL2obbamC0Rq88cJqelVzOtlaHienvGt5gfIRL/E
5oF9DjZu8/iHtohSI+Zo6E+MISPM0Ui5eQd6LUc8Ryuy0klO9lki9AzSrXK8O9ni
cmFXrVqlgS1SKBky6QJAFpgI0NW64raYLFPNk8qqSxa0MzGwczxBbZAPrpkqyGLb
5y8nb855/pZ+VMgpKE23N7vL4jYEXkPrtnC7LaQv4op+fNLluluMA36MsEDqeWpz
3Kx5ixDhQc5r911bnarrDQto3Ltqn6FG8ydhSqf80qJP0wQvfuJuY0I0RwyVYeha
8qHgCzKLiKgfmYe7mWxzKq3JDKZWtRC1DgleAFKOzyrst5HrOOUTTsjDrHrgxLra
acN/jSWeYepelJjXj6MAsLtNDZaJKhx0RZ2yX5LwKT3QYm6fYLCDvzWYXdsULTxR
AfjmG47PALy0GTIkUtzPxwENEDXOSL+UOwJDl5DQ8dAcW+/AHeAvcgkY7O16rP6c
S0PBJQiq9HTYZx4llEAJeQWBPtPYxd+0Z9hMMVm+vzbw064AgYXCvXwRTeTzRdR2
WpNGFjpeGt0QvaD32FK1RbY1Ci6eB56RwtdjR4GlvnpVKYnIFiUGPvtVppkSi4NQ
ss+4VCz9UfY+jz+vE9DReKZrRGotWtTeQp/PU9zxhwlPm6El4CKG6YXzBWN1P5JU
ubQSaEKbUetj1EQOES84Nb53pdp1VGTjEkmMoN4Ek2XmZHBj5BsLDYyV56Q/V7cW
if87WKKI5ONyTr7NWYxYGb8cGJBuMUOiutOojD5f0Vu035bTAs5OAQTEFlGzCxTc
hH6dIRkhEgtEc/MrJvZxp1dtkGN0btGWVUvBmwDjR+JHLyjoI+yCVogXJIen7xhX
6acMkXrJdBnbZ1VqsGdUKdwWtufWozmpnF20r3Ob+iU6fYDsOoOWVjtCr3pE2mMj
TLTws0dcj+lNiRoZ+Sm2YcA1hT7YjM3j1Y/z3KrHCP0ERHeViafP/RLSSML+vP3R
/sSK765fb9wzsviB8cD2D8C4zKzu4QEBi7jR33ZgSC/oOjbMG0ZIiWoCqM53+VuG
wk7gwIt4hYiplItbl1iMwyo0/awUrlKhzvz2MjYFJ23+IZi8waAMoBwu6e4jQjws
Nj4O16JXTyjcnKVM1dx1Q8XbHD5LuNtXlk/+8oEO54YOuidrRmrclZb+KiIRQRDn
eYU6MFdUZXnZi1liAVcv4X8wWIz142Gd26nqO+o9XlSkaTSL3Dshh0QmR4wi6kmH
xZDv7RYdM1YP9k1gDgUtOvKTnRBdEI6ERa7/DMvBjs7puzVKLT/t9Sk07koD9NLN
TSIPW4mlys1H5VRAQadOZ1bdG4ZMhqhiSeS5nOhy449ywG5ZeBp5F6e6vvwcWSKU
xzVBG+uUnIBWnDzLQP+HcAnq1z9PxWdTEPKMyw5OHgvwvVoWkQFLRHjvITWMpQG9
hmZR5PpWbGhPGtXLmn4Qp0HiDLrtrV5uF9mqXY16eBJK54XaJ57wXSHJM0LnB9zz
YyPTOxMKgnVavDdKa2GDp2lBWPBq+Qm7fvK++xvOUniowJ7ths3x2TyCOBVdC74N
AopenOGYjYoSXBcyU8lP1LlxpWlelsJVx+0al3bMzxV5x/YIektrWdt9C1wy0BAM
ySPpy6Flb6e5AdcK1+wrAfLKjP9+ekLV37AjkHh2kizhOn9MmGTMtcnYo6/uvYzn
MyC/bTSWxsxp2ChX4wJwNbl+NBsBKKuZzBw71rHvEMU25Pr2PP2bG5Z3uYvJII7P
ea0QmUXxWYWjWK1c1KnMO3dTSqc8iL6ilufsMqqnuL3Wx1eL65YZ9rSXy2GtM5OO
hEAnh7AzfExpU5I8n9YsfT5FxkMYbvs2qLHG+RDxUh0OHCFEXdwib6r7Tt5BYur4
I6flMfuUKgUJAPfYZ3Ul9TeEFUpDOM+0Yiqk1CDZaVMBtaF2zdub/AnTeZuDnt/B
2l7e9uTTU1A2wov6UusV0mVi67w6uduX/p6E6MErtbfIpDREYxC+h6ao+vRMxO0O
SeZNVhA0VaqvspLlP1clHWkj7+0Erc+sMCVTDVUfBWUthj3Y3QQ5zpWv09Ax60Ob
ubUbEmqxpF2z5Q4H/Gm9uxV0W/kXkBvsLiKNWcD22EALj3SAvP/gcnCsyq2UoWAz
4QpXJCpALh3GYEn1FuoEbyRVDCm6pK26U3aroLIY7J8KoGKGPssCggOt1GOBr1Bc
J1XDnCAvyUki8c+TiHDKkBFDDyHhr/LxDKbz9WFd9R0azxB/I2HYbwt3fjdyswoN
183PMgqGQLchHUreNiLC+Q0PdZONot3COYY3RTTTJlTPUdyLII2+n2LtNzDEUgHo
n1l6VGTvFoDOr8BdjTuTsu5gRtIvJ3/ki/uPpswIksUOq9KL+5IIs7VqoiMS58Bv
EIdJyPWSuH1gSCCldTYM5EvRK0qinkqkiOijcKSAyBmBk4+RJeAK3mz/LTtWs03Q
IdF0gwZ342t6Nu1K6Uy7y5Jun3Qw5L2uCUAGKmqrp1MoOOSQsGoflCwj8RM19HXT
KTQANjzoz6TiSq3d23+scjr8anpfQbnMmmZbjRe8ei+c4jtsGUPTEiBsZtRjhh5y
dBQJOK82orM1UBhQULWKosvzzz5XSakY7mgKx6mx1nRvtVQex3IP8n9ihAW1kenf
SfjnsZ5FbHnL/EU6ptFPb45C2lHAb79BWAGoGH2N7GR8v7Vv/QAUZ+gMeMj+nunR
E2ABm8dShdCeD28e7HqqDrrC7w1PnPdnUpF+7X83M/HEjhPBB+NrA6hIG68/8hkU
6c7jvKD2gR9LRCYW1+Tf/v8csAFUnMeJoq8Wwes37Bp8sTj7zdUCj/ZVEVHih3dC
to/FK5TeFvd2+zufi0d2a3yuIws7t55zEZhLvy5bXdIpsdQ85rNEGP2rbJxfoczK
i4mqr14W5m7M2CRbh1CqO6HC8yb5wqMOC+8kKFvNTw9gfvJfe/B8o6SvCwvLAgl/
xe+4OoqpofuUjH1bxjsjWMECIzHF4Qb8+YAWBrSRXWA1FMR43wNV1njBOVBdXD8A
ubp4vkeFqFZ83VhGa5a6bnYZmzuIjbALcd1RCYuRiJKIrcX3TbsN5Zpn33AkRilB
Ig0IC1ALEn/qxia6aZ4BXgR/42vdfrYlVGZIn/VAJ5nncD7DK3662HlTjOwgz7Pq
yNfNhjaowPxtqIdTqFO6Fk+xqPQAWTBzFugFNvYp7H1sAvMrYzQx53WwoFmmDORE
iT/M2tQl0qYygCJRkblcBwpPO+llbSLxhjbX2+zEbctporW0cRAC8LLL9/aSP5Rl
qaYBmQxOEMRTBeYFLIvmCi5Z5Qy7CJBuH10QIRbZ+0xg8mJNXH+Trv/nIpLZ4P3I
Xd+ZuT+P4yrD1g8XeaDBc47qeHMLtiOF5oqsFnSbsDPNiF8WWv7NmT983UIqWsE8
8BDIBcgcvGF2qTRQp6HGAw23lYYc+ioNeLbl7/BIWkwDtJn96qEZi5ZKnhEaHdvc
KzYoI0XSZ7Qvdko5oJRgtQTE8vWLIKZIhsK+2NnLW4diaXH4aUu+0oLEZF0vvSha
h9tSPsvwoqSmjuclCRJ9CR/K6LgCZf7Xa3rMeIi6aKD33wAWTLQ2YWRPqaT005O3
XPA1+UfGFTuEOY3BB50X41KD1/TVl/dN6+iYBwzdMS75TXyVOt1Y50FL9DSJm4iG
hd0KBZGBBjeCVIWhL5PzO06LXGC72UgkAWyGHPHVEhOLUJwJRUNIxMT9Sy1NSHmC
c5dvrdqyOiglbkcLa3gd8sfWzHhOzn9lOj+wqpt95Inm24nGofc2o4zTZJ61FzW8
p8twgDz9tCMf+07c1yZvkz94ScsPLUv2pcZFygbhi9P9byct98+Ifee2eRDgw7uR
TPRnawjgvuLdvPmr3BiTfp8Hyc4Sohz8lS1rBSfKvBbqGBX9EcduTK0WqmYGJSlI
QgtphNxuGgCFgp3rPc7GWR6H1BzEygJw9b3OpEDVdt6z6X2tFWD4JP8M7TKOAOMe
lCQOsctox67wkHT2y3AJcx0ifw8w65ADOwiJ+rRUOxyZi5Xpftikvp5Hr2EgqMwh
pX3PYTIt8pkumGaFvEl6Fbrrz+JFwMPhqq7yHd64/wREB0U4hfALk0W1/sBLNa77
/strpJ7Wj3XDWIfXiCuawiEMCKQdMgZdkx3Cq3bl2OT1DohVHZFMRGiLWt0xXisE

`pragma protect end_protected
