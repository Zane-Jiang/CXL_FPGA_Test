`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
cZ71EzpnkVdLzDugj8PuyEknHXXITXVCvcWWL4OlpKEjcCS4l6Ortwx0a9nWrDoo
fHcTSuTAjcPmtQ3KNs8WS1jC5KWfOixws0mydxUdbrIdyReGxD1OogToZORBarSO
b+6xA2hee1wdkTRNLlGhxDM4Hls6Msl/6GEv5HjJnJk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
uA9KxxLzIBV97owM40GZ4CBYZvtHWlJ2w3T9PYkDnZY3Cg/yIm/NvGddt+FCY9/2
1gu4gz7FaNQQ2hHyWNiqU46sAZRuSkmV1e2ggqZCchqdy91La/SntBeyO2HJeWls
hk/6c5vIGiAIpPUEWPdKAEtYPeoT0BVyNCvJAvEYdGkrbtI3EeCZH8jGF6p/Og+k
Q24ri44qDPRwf0I7anYgw0jLIZxA7mi+Cxs89nQvD5blVI14+nrScV3agGs5DL8Q
DH7QkhUMvjJZV4CZC4H5EtJCYrFFgypg4qbeikbWX7pXW5d2Iv7zwtwJlgb09Cy/
psJKNUtXtNcN+Gs4ydwyREY+7XVZ5ekI/JU/xz/aSok4IzO0QZDhKu7Mve4vRh60
8cru4qrKy2K11fMTWoMWlP3KO2BU4Br1XlmpEPJ2dIYS5c/7n2J+HIKIOeLKhtad
yk9YLitCD7twBBRSPbsXjLklvJ3Vo8hhubxE3iFxGYNPXgeXip2t+QWDwI/0lsY4
oR4/5+cTypaTf4NH1D4HJBwnBbDLJ4TP2zqUL8RrEXUdO4HhjEjrZx+M2MU5DaFR
B08+iV36e5bVMJhIexEKaguMQGPRpaHs2gjzmrKkeQfkwYfx3UoXP/Sd24uTynZJ
PZB6o/vD+4ytX2LoOVPMR989d6U5H17/BphANVt69//zVzO9qhYJtGHoxJUWb2xn
h4ay533VRBlCL9f6/RKq0Sy3OXTh65tANWsq0vN9ttb1LC6ODzKQWn6Wrou0zdwU
7SLM0pwOItMjK7imEXC9tzj53Jd1d0TiZJLzjhusdCJZ1y4weOJUTRviZbJh+yx6
0UI/RUgp2EeYouR4jAFiUJ5lNcb8/fi6P7B1dQdyn7F34ll1I3o8ECvYizxkeDK/
dBmh7/nI6bQsULoRADatQprumre99etUqz9AJXkKKCqGy2CyNRKulROeII4Gse/l
y+lJfh43kvfJ+P5kQq0m456KgmYPZ2bJxmVD/syfdxN9fnvMqmdU3Z6ZBxSM+94g
+QMgEuzJvsXT79jHDQqV4GY0/Wo0DtdvoZIRt3AybL/yGTyo3OJB5GBgR0fMUQpg
ACEoqmu1aghKhbBGsA1A6NiS2OB3Qx1Cs6HsZ6S4BmDb3Qz4LnJzKyyxpY4vffpw
EyFvYy1gPMA3ytYy1gdpQ5TsxStG0TVGSJ6Llte1BfGFTNMj61D69Ir66aMEIq89
vz+k/doJrHtnCdf5ZOacHgowOMHP+z1Wb9zcCC8JdXmxrln9qAxxpRrNE7YihPbB
oTsPQHQid8GE/HB/BwVCy4JyIdAFGbhMqa2Ld/lkZBLWut1iO19Tuq3nijaYaQZS
TqYtUizXcAm6y4oAeWsJNromIxOSkeHsTHxwuCWTCXeCF4dR+q5LokOkk/SDpnZc
aw2doL7kZ73LQ126/2TNTfr/cQcc2v5FzIZiWVoqvJPBGVoZhQY4g2tr4R4mD48w
1QZKbNl9A0XFitSqwjHi25XO99FsnoUWZGtrHQyUAXaGlsv8mOGmOq5xeEHht+KZ
4pKQI2cUD3OLAAorF8Mmp62nhqJPQqh7fw7Nq6/c1JdUPg3PKigQ7DQw22isoVxN
jPVxn5BELwm3Ztl9N0dd1ANdmp3KgXXoICv1ISvWD2NmhrjaMbYfAiZ5EOmhU0nU
MBVcT+C3mcz639ovMhm+XlzPdEB4ACwSblc82fhllqRgn7mga9+1nMewYMOVQ4UX
oq8SZQtlB6QOgaWlSV/Ebmu40ytiYfMTzZlSeFoYMk4Sjl+i9/kWEFJ9iyRBbjuo
D3osrx2D74a+Qto8qtxkiIeXgdX4WBI+v0tcVw/IbunpMqSEnFntgK6fPk1RFgiU
vZdmJlNdhhd05np+EeiNIqPrAAteHHyZjEWkTGdS8RNcXf9D76pfjoFarComL5cA
DNSatCNeNo2sEMHoZL6KZBq2Cocc/IFLo/Swt4Os5fNVMwO5GplzROGjqfhYSuYT
NQHvPZXT9l/HvE2KgpDoZL/QZz2jgi0wAi0HS1gBFV6YdrRvZlOx/ZgJhulAuMQq
IAyJR7rDUpZzi6BKzB1ACb25VNOIS9NO5h4Z8cWAx9DCGo99JV2GNIf+HOd446Eh
ftcQeBIT2UHXlerHvwtxK2Yg6J/1xMdSrzlxAK1mw4JUBXt9QoY1xnqoovHcBu14
zn9QgvcWdW+4tjEdKzd7DLv2PuM92hSsnwezQ2JOwXF7MXRwtkJSxKxInK9YMHxO
8Z6FL/Tpp9Das/2atlTcVapNpq4lcNmu8usXOTknJ66dvzcllFZ3r0alIJnbdFs5
8aa58oGs7ucdCjAyzCy8jLhBIRW9BPSCyZgIB9xDJhR9m/VXN2K7IOvK/pgrsA5m
JRfL+7XR/NrRLaZjE+MacwlxQuQZHtMVc50oQZDazWWxtQcks8X+EiU1DQpKJudZ
n8XES1WlN7nbfITowbmiQCFRW9ylAEeV3/Cp30+3i+0aPm+mSf2bn3m3MDtt4Yhb
w4XboZjfWk2F0Y21Rx+ObmPsIhd4mO/qF+BzMx9koCNdJW71garX3ijx49wjEEh/
glAXAGo/+q/YXkp3hmF/y6PfxvFRS0bXTIXAeUJmkIYz3x7z6RU5lly0YlwXuUa0
RPw0/boQaPEcwiPUWQDnagJqHCkGxwRW9TX7nM4zs6NWuU0tEPGfuZed/eWMTsfl
KShMLeUQiYKg/8uuJIdCjgVkpSBWI4AfGuaohw69XXZLLc4BjZpRocN7NvA71AWV
H0SbIYgDYkT2Lw1Z5M1mLxZG575/0UW5DVy7Y4F8G6ptxHhf09INmesCtnU34ATk
x7aU6fDHLxrehVyfV89rDNJGOVegI20V888XUSbrXtE6ZFRQfvVyMBUH4BF7UXuO
3WEWawxRYGCtXG/KYha3T1VgvJa8zmeQ+qTDsYnck5y6RsPHjvir8h6d+idxz7Ru
jdOstThK5Swn+ApenY2Rle6p+HUMR1xByHoNXWE9M1+V2X+JAuleSTqlZM1tRx48
O1Gal4qCHb3sdUbFXRh+lbwiM9YO+q9pm0cB8SFqoldBpLJiT75r7nSpdGk1bmGh
tSLBgfi5bziYTpJBwlMiGVP0tTN8FYJs+GGjPQP2nM75zyLjQLHknauMBcz753e1
aQZcM3drA56EYFg0wo/lTeI/Bs8ipbJ7tWHVtlpBnIBCWUheYLxL2DlIlgiP+Hyh
6JZ5zuJOLREmS82+tjiVDXmupcEM5AMS6ULfdYiSfjmXIe76b5uwNYhtcSS7/trL
uXd8SR5797HXXD/b+yrTSfeWMo5kfLy/BQtPuwwhSHbfGVjRrHw3m+rNIT/vpVy/
q9n/TDY7QHnkZkyCF93vj1+oyKf+D5pVy7rTqmIOmPonjtfy7ICO0WkbZF1WngLd
AOfZ7NElSzw4CeqQyHHiTuDgo2K8QdV8SxUmkDfxUEFR0JPHkYI9ecIf9t0Ze72W
xmEUsKI7zOCO+/tmvKVkO8LWj4CD0AuauMUwxpJMT33o7nKK1Ey88ijcF+xGGf6z
8P/+6pM3u7AAaNeTxslJ4aLOgL53f5oYOCXkIl61asoq1WSj6llc3L5kQKEv6MWK
YNXMOAA6rCao1UEvkakfwL5UcB3QGpoHuNE7pVQBRPeh2pz+cdoAHQcPajDT+3+1
rJmNkJ5Ubveo3vMsEkqTH2OCKqqIjJO8ACswp31Ug7ALB7FHrw11NnEPNyhBE5PE
VyjPjgsAUUcVHYpsaMxS3PesfXk1qFcLwoA7bF6mwmfQl4gSvFGMBFy+GcKEVNct
X+B2Rd/EVffUADV30IdUUvZEkadPUT91f3iYdMH04d3PUw/KCAO1J8Ut3E07Oy5v
pq0R8ldbSoY5M9iciXd9sJa7C36PMWjDlrUhQVps6zyiGZr/9jt3d/DyphgLCgbg
pcSeXuLnUD/bKCIcIv8PH45w2yzKdQRRJdgxRlmvOeaNAKvWZsi7PUVHb2n+czDx
U/g2fLv9dYzTJH92k12TaJbOejwxREtdYU4aOHL2VqXYVLuaby0DrDz9LD6DUkmB
NgXKUg5dUYqaQ9fKUDmQKrGwsQFMyMvlg4PzSB3oxm37Lu6cbNa5pZlsms+NhRPf
Q/2TL/j04CvDimcB9I3wxLSk0NcYUE06MBTKxFwxKJ52bfrqYhhMLoRczxmNq//+
4H7jr+mWmT6ih26trm3MaH0CdP6weIvru2bZagsP7E83xkzjHxTqs8WgHIcTcD/p
J7BFp0N18S7UrnjHWDGA7p8j5PUjcgJxlLF2PbbA6S+TkN9t8aqkdPNOWViWxbqU
fQRJ55D463z4iE63lXSTGvtodk3/MNd5GVwQQ7qRoeCuIbjV2n0Ns/vQO01shAp6
rh1q1o222zvv4VQIyen9RobBFtzpe0AJwxMTEjUxjIfy7k2QPsqoNIdNgFS13AQQ
IXM4cZ03yWqb8X0XwJTz1VGIiLNkbbSnuUtyS19gber/RmrckUZ5DAxDCOlGfI9B
W6PIl/voLR80qyBMvYs+DgrgNTBG0uohMSvisjS5rof7QTrQgsW9GOPvhYRSmFFo
Uyy2oaCzgx9OfnIEoVo8DJ1uNt/lQSkP6Cw2fF54VjNmmBOyBne/USCanP5tnokx
i1drGWMlppsWcjusnvoQQf0/TFmZCaxEm+JUmOSY7hsukk0xXPCr0HbOhzXRFsL3
Q36YCfCzb6RgpPKEng552iDtCd82XJksl2ABkLxgqClG3nvc5y66DKYKZ1RvIVlw
Cih/WaiipVMbpBPO3a0ytFUsxQiPm7p+4+jdBukGNlIACa17Ste3rxIPOich0RaU
L6FmrGmUOK/V+bF+RaFeIByU0+xzOHCn3XIDLrbsUu8Q1KI6F8rt3iRoSbmm2jXs
JiNQJNT8jSpY+5bdQXaW7l4BElsoNMOJ0wKW7XcTm97uKJdrO7LqtpGxydgHFL4/
oV7ifbMR3VmnY4Jpoofw4Y7pd0PRMMMFlbEqP0SeFhM4qfgtxtGlk6eq6GxzHpc0
hL909PwkMuZ1infKLWLsS/07Z2H/wG9hb4eZNkArWlkgeVMPWNXy3UtkydcNKhDD
BBrtZ8zlnYtD6H1AKvlctpL4uIZNV/fU0GaOcMfnov6azteSTKp68Ytmja8DfSED
ALMI8q5ySuzV04Ys2BDX4KwFIj4KtV8T570nbnjy4Xz9gaFEnTxQI2DvYiFFw/kF
SHCd3gDUN+Pk9eDSSnmahMJ4PzX1yVw6HkdnepH3tG9RwpIab9VR6n0yihgszvBK
u56PmGelkawSoxGBOQklAJtSeOdXqTXshjP0Om4+ZG9i7pzANDcNa33/Yf6GUaUu
M8HU72KNO1bYhlp/Yon2nLpqlewnfSy183jxxH8MX1ncyKI9+mh3pNHVpQ1Ssoj5
6eHWl38rCkYe4Ei/wmyqhpmbPBe33k9k1c8y2RUXfXLmNkgOasQibkKKSHIpoFBu
DEN/Uu4rPEj2MLTdX6COCjt4Pts0YxPeFA/0X9xSMdw01nmnoqFJKcjWwqN4wieq
lhneP8ga1+wHNhw17YOURQlLjMUQ74nOrh0qu5AHM7T8KVzSjocNWYA8olanVmvL
8fkIus6T771I215ItA8QpzjLIePnHfDswBf4m6JYRMqtfRF/xxZIwZnFuQxReTIs
DfaRhjy+N6s0FWucPIJEJiFtdik+OuwPi/iYtsvFi7w7MJYaCIQVvo+JQg6x7lwF
YEg5u21im2nik1xLWFmdcMKOwowTeari27SYmkVNiGYh72jQyiW6rjZawU/gO9di
3HHPPwe+akJ46S4KAvTv4fg0dI57wAmtcxAhAp6f/Vo3q4Cfu+S6fNtR3dYCakh8
5m55A90gGVkNfw0DtI9OPmcJCxJMKjptM/wMHmWHTzP7gFxJsdHottzW3C9hZDCb
dlMRzPD//hBqR9W72+mSQaA5LUeMFhf0pD6UVY3PK8zeWrwkpLXhLWBMATEfNt2J
yTj+kdzd5k7ygCTMa75r4b37Nx/gN/5FFZSvr5hShATjbYNJywLE6Qo22i2pmgja
avWYN08Skz++th5Bm8AAS09Rh6DEX632V/rIEhszV8q+hGYCdPYb2FQTcvYPXPY9
PhAULDY+bjnB0tAU3hs89tj/OLqGQltTwF5q9sQ1Yd8mzFURT3BqEAhVCnUbNtFO
9Rjfs2b3/keyBZOia+05YNk32okAIE6q0sDO/iBrd/qqneu2R2dWVfjWJ4b5/+og
e4WuDWgvmbrjDUfUgL2GYItO4PLZ2MDZqBAAxp94Fy7DZBeoVvFKqzq7hpDelLAu
JShkzNvFZpnl+ZNqtpVeXXTXIdQiUL3IntE0WxTjpW9ubyxQn+zMpgjJSOIgicWh
wNwh1nXpmzJ8uzRhb9tCBOSQnM9y2pqjTXLD7yFjg8L06lxWDK6XoRZgS94FQhrc
KnvwLKMm40mpkm8xpjDk7aL5LjAkAmMTNNawRaHq1WevwPpRhqXI0cF4TFC/bIfI
0L+73QTxnLh6cKscJnF53sanHSFJQS/1pDdp9u/LUi7c24G/lWb/0LeLNtKg9o36
Nfo1TQ4ShiAAeLr6nu5SezIwHf7pv65juvaL1OC20/Ojo7XcfbOU2cBnLDD8yQZJ
/Mk7lb2HN9TFbP5Amqn8aTMQLaUMgaHFE9/n7exr4sZaB1SBuf0Ji6Hj0TYUDmbl
Ys//J7AfS0oBsld6u7/TduLWfnGBwSjNajy9Fh/HkOItiGOagip0aj2KWjh0OaQZ
/ZCgDhFFQX2b26+kXl2ryPab+6sYsfPVBU/qpOLTc1ymHSZIpGyBhI3lqOdCISNF
IaAH9dwtyrzAtwlg2gXeaEmy4rg2bHaPOavwYqhCpWPelZ8D2G+gDq/eodNHRFr8
kqRYqwlyqXz8m9NkHt0F2HXyd3VLnDxMwn0pn1RTxPnlExskqm4+8YIhRCSTasna
VDvyoUMOeYOeTMw3VNYyLyUZr0OzNyGiuSXy8O0iM37z0E9czN2su5VEtYri9XTm
QvIKisMp7eknNl5YAn1nXss+x9YgRMAhbjP/Q8Kj49tVegxBqeqVLLC/Cwevaw+U
XW0XwCHwTV9vpkCxjCRBX0eBRBSblAXIg6UswbYf1Vz2Ce/NX2OweJyWACuhc13Q
9YYNG6O8dmMXjRH2LrD0NUqNEBgAuPHP0mSa1OcsdfQMBtbaf0A+QXeimz8m1HZj
er+dY80I52BwXgnO5XUv1azAuOrAmZqS4G/RmTfVH2isXKxuPGcFoXTV9uLMc5bM
Xv08rSmkZcB9Yb2OGG1FxwdXnQeeQujZxkX/QUTzbqBejHquHzRFWGinfopTlRh/
RZaPvdosfD1SWyTI6Nzp5aKdPGM9zvFbwKLW4q8Ewwl9U1wm6nvL99HItVSW7M0r
RU7EeSFf2xDgbRewRoTOt4dAPXsfsRapgRjzXaroXVOQdn2K9/OrHT3N76jrDfib
6/uleDMcopBvuP+pIvjyeAgPRhDu9beB/LykXQltKyHoh9OJfDufiKA5oUDsc5+c
W5BlPRJFxep2za2Z9rWCFDkjK+2MV6tTe1DKPx8wUa+5WcjOLdSU3NRH9HKQIWfo
7GEX6/FVgLGekn5iaSNS5glrGT7qDHm6v/1LDA2/9tyzyYlr6XL70WXLvTe4QKgI
xeNG8KH57fPCA2AnSVKohamNKN76FQyYADx5hbIHbSN1xx6TfQPlHhADxhXP50sX
96mrGiFXRmkAHzcWAmeKl1YsQdUL1ClJx9YnAu08ht88dknMZq7xqUJX26nf6fNO
PZROsDqYRJPn7JDsNKdX6qQSdxnwtKVPy2C2sxQsxYg2+jijUK2sRmwBa6Db1+vh
XBejlVCU2KpmJBFRTTlrcIYuGLUNXvxGvHMyrC/x2nUmuWwz8Ig89r4nmnva177a
D6/qx352dK5uUhd2gfdbn/VaBStr2/r3rPyjCO8MhPiTLmM8QQZuhiSrLy4MlM3v
/jRg8yCa51uOL7dDAfPr566ZF+YAkaY8xHAwbqipgG0/bVLyzDfd7Y2CtGPVm1q7
aS35Hd2GMo0a3YT0HqQrNlwdjjYdDAgI5amKGSACHckzto1j9CJwt7M/l1dbyZs7
UZn4fx45nNDWbwt6lPb6alrC7QPkxvIi6LwdYSrFwLDdRx0yoW50wP27+L1L8In6
i2WUOl00MzcixZzFqZVIxDGDSi1FXh2XoIt4sHwxayTA3EeMcl8wNIEvTXy9Clqb
du2CWdswiBoWFhiIaiWXFkpFZM69L3K7n5FL0wMcWbL6S00OOD2N5HOWMQJLl28B
v6iuNSzo8vfhETpCd2PCqSQ4UaLCLzb+Najjinh7DyK/BFVEpd9Up7fLcFokcwBt
UbhkYq43vgJ6VlhCvw3gm0Rw61GyhX0jbyqph1bsmRagAvT4pgsL+kJZn315R+Tk
9LgfRzF0D4puSn2nsL6EvkdxnsnZlYmTyHcWfmHFfAOCjDMbk3hRL02sk5LZZoDn
pTAyIXmx2ppSLpVnne/YbGsd7tOKY/V4J04xv0dK6Z37DqaUWHFo5s8tTluICqxv
PdBc0VGNHiZ088LN/dovum5yt6Sv3UMO55oLz02NAZNtzhkRngzalnIF7uprAv02
hQX/PO8LTn7l01CreIkh5bGyFadWsGOJInYADrWA+oxOKRPQUdTX5gk1UZAnuoW5
yYikLDWUPYOFURgM3Is0R74mPWLqOatbLz68NBlEc5hfv2Ji2aS1BXmQxv6q/dXP
ce8RAi0aWwHOd07c7wGy9EhoO+GSnB2XN6IwQ/LfcqZpuAc0H+jy+eMvPEweHJLr
OiOG8gd5oO7gI7fJd1fJHwOl8zKkIOD6Dwpd2k84E7fn7vR/N9Xbt0RQ5oOL5Ifh
RVOPtZ8EhbXGwhjdQMywAQgegPZj2BFUZ5gwcllZ0zAHN2gs6uRbsc5CtYMjWh9H
OUN+YTShrvBGAZK3Bm+91DZ3122de0CyWZHQC7EZ2SSKPfMHw0wjUGdqu2tHt+Hr
khadwzYx5lYc+I/11PouwjzqUaCN0dYBZJQp5V4KpSwY0a55SkHBsRvXcSCiRHBL
3PHr0gDl1fbURtY7Jk7Ds1Qes7bfHTj4iA6JBZtWgufR+Klxo/RJqRadZ5/Bg+gF
NIWbF+hdnTlLO6AlSLIMV8q/bmuBPqNHkAdSqHVTMJLfuYlFgqatesOY3f0mkv0m
e31/vgmZOHB75wD3ckkHf0wd2IrPSANzh5lBr1K0q6OQ8ksJgtQEF5JPW2iCkscG
M3/Ogyc0bulvjOirpGWwaco+HCg+vCuGceBTSGTp+eIg2ed8/ZPmU28Gdc/h79nc
ywNe/Zhplnjk4sYhcwe8RLWzk5FdaV7/kTqem+JRKSqNrRsE27dCQD59ioA7ESdg
5dDjHLBegbvktcZQ0cP6njK0gdXPdAgK5TQ3xFBekt1DSoqZfsdIcaXDuVSYMT6y
2Wk1eRDK/elVXA6bPyW6uGo7/qAgyAaI+rpoAK+aT97bGPJc5uOo+I3I+tvlwYPR
3QHHuzE+8sZxPtHTnC+K45Opq4lxlmPIS3YsTF/MS+PWbzj7A3Il1XUl988w+SB9
jG6H+EoAPG6gHEMrkInVUAsErFUOcJx0c64Ic4hHrDdlyzXLqTh9i4Sk4khGljww
84n/h2//+6N3uivSOcShVziERhNKA7SSzWrd7ym9hEkJ5Lhz2ZRJt2lEGX8l/IBg
+JRhuLTWCgX3VcfvqXuThK9Lp8K66P1+3Jfo5EtZArWbuH7lr6VQHDXTz006/x8C
NUwco6sdpFjPX9ABybhy+ciMDKN7j/+eeg36gWKfj+HuyPwiTbFltMaCf2yAeYBY
ynNal/9SlB6ukFc6kUW08KjuuPG9soFukgtKWC7ibFULnaHvEFXX64nferfSqw9q
XEpsmO6qS+gT7JFxcqKaACSFB7dX/FhkE37873GTB/KYmqOfkxX7q3pDyy4SG7Ht
4mPf/bzqEiw7xGRpfBRoU3etk0qz41l5b2918o38I4641BIqQa8oofey//na9js5
EQGa9iuKwHDbBMffxPXfEWCxW77PcRREVprIX85+cFxYX9Qx7Z2YM302g3iNQM71
oIJNHZ4EHFUvB+GnV5CU2BVfQeu87/tAHLvKnqDe9kuh12Z+pTABWpU+2OLgMkE/
6llmFaCc1w/vativdDhpjUpfXmHeLp3oy5ycpGi1zdHc+uQEYdqMOwYV534Ss6+v
k8v9tNAiSVVxD3O+JCQGk6zk6o7Ac2DstUyJpwqF3XFCgBFNLiqoEdhNeZMj3IzG
P5u5rZhB7T0K69F3opwgCRQZJDbb6I0sgINoXe7dWu9biMs4DaI44YsYojIpolbX
vBgctCFRCSZi9IlNUBnetgb8k3xo9lviRQDFbcWZYlSe+HqMEpN09tbNU0Smqa9/
GcMamBWZZPpSesMB/ykqp4M2oMYYIycm8KxoaH16CuOyd3aZqBPPQWG1SOef3stL
CVpacA0dUz6H4LodVYcsPi41fSlMRnKLnNHBR9h7N85xYheSfaQjJxo+2c6h0Q/k
4AtqOCxMxEcorkq122ndYWpv2uok9E2A2P4YwFstSznVBTFuzPCrM8AYT1LJQqEK
pHdtfg66rqwrPXXxfzRpgkxOAMgC8IJa6raryWgnUGIKF2QjAc2cPwTj7VoFRUgI
VLduijOCYr1HjlHojveauSlOhYT47gczJkqfxrE2+HoqAgKIVvONKcD4cXVIS33u
xqmRKug3olbv/PqNAZhqZ1cXuifJbEPI9siZ5Dc66l5/vQNvnngqR2jL1s5neyRE
ReZjVkrxz6piOW+0oWLT0nJXye04OBesSIA0T3N640ZtVWJK6z1B32P4S2cPvWvi
TDxTErn5YA7M+SYQPjC3wyVCZ4DLYAffOPpTvebcHHcmWFMV4/8yNdpDoOyWTVL+
2OsOmm/jOzqfSYh/6NSW6JkDp5tT1fZeFmQ3fc18AxRTyCgyJaIz5JP6+rG13gVw
ZYH/3pVGotBJ3YegaBqp6wo0//PZIQg+xKvkdaWNr338HPm5vAp1om6fr2dBqFwa
iCUiwVO/qO4cWe1U99HOP0R6x3e2C+cZ3brrwC5mp/jJSiAxoSu6ZH3gzjgCGrpV
zd8pqDYzEhhlT6zzM39h8yWRqtF9agVaipv+ath16D6AZkaY/6GJa/vZ6fWHnFz2
t7j12JpAzdzWQgLwYg0hg+fagkyDc2Q6f1Dhm8FwPwqcYdHJRRWDAUx2R2Wqh25C
3SRSZahTaDoAoMkfTD31KYzjzAarCPYXLdjg2ZthCG1yGlUt/lg2D4H6BtxW2L1m
iFk9wAsneWit0mB4XgBiAHmu/NxlzPp3tqz99GySs+JjFlQRG2AgU7APzdpCxdmb
h5ttHu8rqiGLH0JJauB3BXpqTPW8ZLGieLRbZKTG/NNF+WpaMmSfrVeoSNZ/guFv
dM2ihQ6Z4Und4LGnt28kNUH1tEPffMwIvjYnBJNAt5Y=
`pragma protect end_protected
