// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3d++bMdNlovIKUZoxQGtA5hF5Um/Thg/CXrypArp9ffwMUr1dDiVcTgxgIDNrn4F
MqBhqPL8FGqPhTUm+1x4IUWbXs+bKDOhEXHZvp8qsnbpoMEUF0FGsjLlW2le83Mp
35sBsrFYyU+nJnjDUKZdaJlNgEWoPG1hwPYIo8rfLX8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 23552 )
`pragma protect data_block
Gf9DNi7ww9NKf5Ng1pmAcXueRZNkTMHmubEa2q3ILrgYlbLG61DZ+t4X/xxzVyuh
BjTk4U1aRnerYSl+t9AXroLno8Uvb6TD0TanNnAuXsHyMEJu4nVI0DLveEEfq5/y
q6XPjSPvfYMGfTkZ+b9S+mQeggkxQHZOXVgqzq+yBqv0ll2FyrQg4xTdBVhQxzML
+l2pcbRNOlIm3XS4iknNz8CLX1aKh+djozdHz2ZdesYfNSWm0h1zOr5+zQHJRv/G
N+rv6ak7N5iiyJQPxNUquM3DWrtMUJ4K5CEYE84mR3vzNJoftJXF4bUo5rFjnoyZ
L1TtihlZrIyi2mYVQqFFEr2rXfPJHEKSlh9GMH8TYY7XoFJQAgbIt5iY5cXK9hSW
cI7/XVrta/EGYfvEXD0ER0Ltr72SF0FZQ0G6e4C8ZN+Y+aoi7N/mc1X3D6gFF3+P
nmi2o6Ogxct7d3nAse9lHDf0wZpKBviiyun9bezZMEOaP9jsK6lf/61gQTitgKqb
RQlf48w/DQ1+nIDp9siV9qzUX5+8V5bh6dZDxdz3gceDM1S77+QJe4qh++PGldkP
QT4yr2XPhyfEarJqMN5Vi8NoE1Fdra009U+gqjkhKzTeaodCjCZLHedr++dY8jHp
HFjJB24lYCDlo0NZ3xczmI1Ngh5gu2EIeMDPVmGxfYhFMGkISb37sTLSEbjr0r8Q
yBUBGvI2HpfWmmzZ/cWFxDtxRKmVH+aUjjdWlc+5Ttmem8QnLLnRG23yEJg20cok
ydqAdy2zoKmBqy2hBiww50roC3qOu6oJCVdKheBQKm4kBmnqTQpHACgr02gbhVCX
02RV3LmWBbSW5crAr8kvfXCgYwsFdo/qRfb1i5zYSp0n5QlI+SRJ5M6M+F94Nt44
987msamggmiwjrPR+2SPACnhusMDj13phm8WZySgpqDTjFH9/0R6yt3b2wS2l33c
ITeGVfxXION8bK1inRsOPeJuzWuQEUtB6m8Qympq40mg4/2qrOssqIB0CXAgq7fO
05x4qZz/pFwSi50/OCoD66BngHi8v1WQ0lURSAcGr6Vbm039CL6ON4N1NWg2iMLU
uIwfWJP3757f+d5u3U/UtuTbg+lbhEp5yuzlY9COEH0wKGC3YXwy6N2OqNCuELzf
lpC1xzpLOHYZPjcLWCCU8HR9FrJ555NZdX4yIKwl2gMCMFcNlUwjf5nkryTAxQ2q
YLxow81/wtYPCbUQGUa1dHXDQ95R8mODccfILSK6MqkLT+d6FGr5xD3cfJ93ItT3
Juk3Wc/tFi+gAqxp9OoIRS4qQMM9hqfWGJrAKvlnO9JX0Brg9bIdPI9671FURIW8
2OeCtdmr1Q3L0iRZxLkBZ/Qf+DsoP2ggdCDZ02/aOQ/yT69jWdX0Vfk0YtH+c4PG
rEo5pWjmXLO7arqL7nRn9ftiKFN/abDXkFyLh57XAWfmVZjUG0l7FSnkbEVcY/dZ
9U/x4tehBoVHyjK1+b0Armj8XrbmHkGMo0RkxvMJOwn8cptXk3N+V9lrgjLPUvK8
OYJkk8JqbzxZXyBLkVVU03w8ZKCON4r/JaeBPyD+Tw7aEOoEAJjUgOgc08pZm3Xm
UHrTXss6zsl4K9eUF6ZQvZnO+a9aWlW/DJNcPD/O92uStXRtBp9j9445RIdZZN9o
FMnF6L69Lj9FGJVkB5KTqrYKqxtKr6TWz4RFPL2vr3V1wQ0Rn5UqYq9vT0nlx909
r3XbMQ/qOwHc+yqW1GVbtWUF1DB0VmMEkXQA+E3eeMS78kvIcBkTuxxheEQ1TVXs
SX9fmINhYJ5NCemH5YRGsbW4Up7lfIV3RcKkf2rLN3QgdccPFvbLS2QsFB6mb/mP
+Zw3WYv/7PP6ArkR+ud3X+Tq0xA1VZ0eGzMN+3L+BTf8DkKHFATZbEr3GNp+jdLi
3ZTECaNJOGyiqnTlJ74GewlWB7ud9afJfoAKvIPfOGDW9fzb3nq8LzVx8QPVlOM6
jQS5mHTazkvyHI5QcpaAl557jevZlf1jN0COZS98lXU7g6I75xDBGytOT5YxbP8k
HbYlohcC1msPSLSQp3cMt7a0l0NfjpQg/69xL2sVwoG3S5PgSCqRHaQBdtY15+as
s6BhHOFZ1kQTxhptfrrIe6Rw8DqZo6+od3Q0eJeOhsTKtgXJ+kwOUPZCcHmupxyw
+uyRUXuee3tgg8zzv0Z7MGxef5oNHED7kI7Nk8hh8ozdWqEslvmRShW1TjtfBq9Y
1unxlCauH2q05iH/xmI/+l2V/rzDmCLVqMOUtpf/rvdBPfdUMJw76nCc33NrNjh+
FbMupgf5Q8zP7uNCPsG9KsgRm5xAGC5NCp5dYZJZEyhk+hY9HMf923xYZ6wX1PjJ
+gPquOedU2O3dOZmWTjXmvXmeBQMsSl0DC8/meB6pAZcbE0/04ZXUVn+CIsIZ0K6
kvZkT2NcnjTrapndTN5D2dtDUnEoufDJrjJgWJ0AmnXEe8xhHy3J6HuKWFioCCJZ
o3MmvitFJfY0/FP++CAykHvC2De1WAHQFzUvBe9zb8DNNsAF00yhg4UKPezKzzt+
MvChXpRazI4YrgUBRQhCbv8V7jaulwKcO+P+H2WgO+EYwo/R4HenpzxoycDrkOpQ
5fJssbTsH2a10964gJil1a/AnlrmV4LKCx1hvoQ0GOwDPHqohAswhB9x3jUPmciG
E732QhQnPv82ic/W+AWqHK/YNAiVD1jqmA6uZt6yNfPuVmULRoCHcSOyMAwleLgD
u+zXwCAu6546Zh/OvMLTa501h1y4SnoKC1UMzJ6bCkKAyu7MzgHnpWFakGUzNdZP
RvUo1nTET6F6iOxhUp3VrxDOXxrgZOgBmVu5zBe5WDf4Et9lkCx0Ti/zPxsFjFUp
FpB0gu7sHCdwbz4L7gAUt6kpA39PC1VoH8YxepMscPMZbOrQ3SgyWaifggHWXssN
zEwLhzD81jeYs363ycA9nBDm9uILrQpDA+7MtDWwCYeuXEBHyQBetwMAZsy0Jjb+
7IrHVbc3QoRpvIGEeezYmWwYVdAxfi612OZEMY7EnY5BiXVM9kz8BmIYZRsu2Uuk
HxZJOvPYpB13ESku50bUX965xEi4xvnqZPAofFm2XsuugU+BeR5NInnqQoucCj2R
XWoNTYssQhekLauAJ2Qz37D10FB1urd7CD1mpE5hgmQoVH4bAZbdTwh5Kv+gD8W+
16/DDJKpDbbmSdOovYJwdvFLf7Se8gbthCqCaFOOTWt0a5bsAFRmbP74UMFNj3CF
/IDBrxTfj/tR6Zev9ssXn5AjSmDgIHEWrQw4X3lA/RUk/XIxRLaVfo8g+XDQw+ZI
9iWXGN3OoVShPeP+6XkTUhS1jCbRVQBq0Sv/Ozsb7j1r9Ofx8RGfmMwy9jdcNuaI
P5ezJ4aLTZoc4Di0tDHlE+hVQn537M9W+V+lj0HVaVvXkIxe66x4Op+G5RG/Czxn
nCnVmNLN3HMqcP2M+HKMktAY1ekCCPk0VzudDHHdOSItZmn2Qx0Ed20SXHne4TcY
AoiwkohRU3pShkqM38pArjtSvH6Nybqns8Zd9n27hZBOC62TPBTvu3KFQ8pio1yy
qOL3o/M2AfDN0lgoqvJOWy8YUtNHv/gkWA+Fj9WDcGAIPecEuwX82f4p7lhg8xzJ
5skj/iHmJ5oJ58ue4uzyZ9hVcqyOeScKLj39YjuOUp1HiK8r6N3iIu0Slhu7sakA
T8M2GHd1x/Zs0rYJXSQxQj3Q/Ssn9AFS5E7yNmwnwlGiBEw8npEHnX00GDdBMq51
uiNZpDGnh6wyP3gWSJI5Q27kmuvh+1hB+ivWzgK19jdt5UKcknm6RSuZVi/F9s5I
X19GC4tRhRkuonXq/KH8LKJ6cWNXGbM6tY6I911xeAM0TJCHPdi+XPakJzqIvJHr
V294X0w08kXaqCjiHQZK4fPgiS+mBtVpxEx8KJalw0QABSVRIknUmEFeGLve1aYa
7Jjf9YwQiHgyGa12QE6JuhG34ueYmiFK9lLQNdtB/k7TlRZT02VxqXetPTwEZ1pp
fj5DyGx4ENjPEQMPbFXbjWvCCEb/FEEtOhxA36MsDXZyEIjYS+Xg5QrSMQL/yCY7
aljhsy2lsiHmSCji7xiKZdlu39FfKE6cR/iNeRqEgay58j3dU5q6bYoNacQJIIOd
aDjcN63vKEaOxMbv2xIE3CDwST+Qbe1WhzSkUOFHppgokww1NGVPU94lsFewy+i9
a2nWgjvvZbtZUao3aw4kShmGSrOpaDUfKaQz1F44LON2lSbV6wkUx/5nFkeYA34h
fdlPLhDMpQ7+FWiPvXPFyg9cNaMYoj3Hz6tkDkiabdIMjHs7Xk+lnFz8K9A73X6E
EmA34nd3hAVFj+0W89TNXdJ7MhJXHzjI8wNDbDc7ZRR1fwX5pPfwvHyLMuApkFyZ
4aVKeMzuBTliQ9pSBiC5eOEy5QiTedVuPZkpktsPcXoKaf5c8wrSN6o5LGL4UdVz
GpCiM/u6EbmICR113m1uFHuLv5UWpCrV0h4s3YE7LbdUtwD6liuQbzRF7xOKHT0Z
oDYBQb/dOwD4jjORMAruPQ96LT2ECDexKWPD9B0jpjM61erN+3lBKR0UXgP1IMvi
iUj5UgdhdDG4Nta8OEffVoaMJRENS6s9yMFHhBAFRcHaL8gkDxa4Id3UN3GcciHg
OLljOrdnQZTwFrgFnUmtv/tTdHyj8qKNFFzBVQAyklU+Yy6mgeyTk9KwfAN3338H
EWqPRiiy+VkU8gM5syHKWzlYc29Xz3NijidOjB44lKl9wCgHeQGdgc9jeC9k8gyR
5zzLEIYx1k5nd51kC7+2yPDw+ZVVh8XDMCQG3xvlZj9yT8APFau+mwMqq8HzvRn2
q8gBzcPQbwNaRsOU5kdbJ+/bMCsPU80ad2n+Qa/sqlCzEyw89PFzXT0D4twzQpVX
XKArnR0748I4oae8MCkuik/7NFBy//thsYHqWkG6x40x/lBB+e055+eZGR5qwf2L
Toa2Lny+U0u8f7jpnl1V0GMmWRap7ws/0k/2dO1HjJzKXSA7yjfDdm1VQa4I22GH
gjN9gU6Eh8ktn2KvewK7aThZ9y4ssEdCDNKgM+M+46sLwvl5hkN96t2PWfnUYaIk
06V3MzM1QyKpdm+KjlrB5Lu3QTLI6g7UHfM1z2y+N5B2pzvmdGi5lFFnp+xWAi5d
ntrrvV7u8WrTM225flmAspA+2o1FfH5uQ6N0GKU8zTsHiW6MDn1FQEYT2AKvuBLH
LlL8PYeYYaHrjvVRUtQ3CTgOLlU7qdLLP6WzMsB0ExF1AUznpDTVEElYjYvZH/ML
MD9Xg4MufDIxA9AEdv10ma85nW0riIe1F41B5ITyr/MgZu04jb+0OJzovbBur0Ao
Z5Vi7H4wc2TL2ydj6G47PcH3V/Znvg0ONWQLYkGKbSUjAwdE2lnhs9dQP/jBfpC3
hJ1QyWNjt+/Ns6c8ORDPtUCNAKxx6M5Gqdv6blBrw9dCD5FwILsJyoidcCDKOLoQ
/XXmCSbtzdukJRtpSwPG+7O+Jzz0FfMDEwlKfAlJApVU310f5hirSYiLfgpPm4Ba
r0SIkuytokoonyJFcxYiSr7MS+06GOVBB5WjeyAf2xktF0uHFkM/el7G9gurrVs0
ZDwA2AhgBo8WD/V+9cQLIQmAxdq3nJ0tK2D8s5HCqFh3/L5UKdSr4JWULEg3sVKd
/XWojSq26mzhywn58lme/AAbjJWszTNcNIDulMROiW6RPjm5TTkmPzrcVXglw6Pm
aQUVqq2JVv/+5B5J4BWPlJTMiGUCnmE7riE8ObcBkLMNRUcM6hFuPAbVanfOcD3m
oNGGQfqWJ0ESlpXbe4B7e2cWUO9K7eQdoC/HtzVMNKVzaju4Uhs9Yo/LR8E/7N/e
4JwJ0/0lNecIQgdH3FSbNBo0PtNE/8VVUqbbfgEvgmptcErm55tXvp/EqX02jlY9
5WxwLSp9WerYo1u2hUvv/SqV8DuCLHRJJUYPVrFG2BwR4Ato3FzTknB8JRLxWahQ
qEcZlWtEaJ+99TC3eaF98AspLYukQPFmtnJNpkTQpYZzIRMOfYF6rgKOBAiQupd/
d3qWYDYwqmgJNnopMY+wC53WenhNaa1fmNNnnG4yowWDmyxTmxFtNyfV99Ag/2iN
FBz2JaxOZI4GpB5Q0Ej/sa30wD8iaDm8rcA1BzEgGVV404Dzb10i7jaMwpWtUwwD
fT3fdMb0GTgindwjY2BZmNGt2sqOjIBaC3tAQuWT/Lxk3vSimwSi+v6NFq8nJ+ee
5W/bLKxNXkCuZka0S0MQdI85ORAYqi8Eghxe7cZj6pEzKGcIEi2I2xGYY2UMEgl0
ofOtNcq3ASCKcl+98EQeO6c5rXVDGv7M7OyRb3MZXGOafDjAkLUPQpoy+qT12/8l
Zasr1z8tRqdhtQSDf5k8eSdpYVDShw8d6aE8EELFRJwbQVMuTl9q+ndbHGT4TXPU
E1nuE2SH1dvZC8w0BfH5/GV+KZCRxx616Gd2HMIpSya84Itwykra23thFyftpafC
bdksHM/z9A8REFRCK6gse7hgmw88MbnegrwAoSJO7xvwGARejvfNijw1iHu64Beo
qbC7OBoFVqSHKfE0CP/ZCAR39UccsVLjf5Qwyf5vI1vtOtyfoQtEpeLLb02n0TP2
0QhAU/8/7GXe/p95TD+hxCXrBgn9WsGenx9HhMLKj1J+U0vjjR0chefn5sGsmLSe
dNXVhMXQijQQ/vtxukPnxaG8cuUMg66G8sqzK1AAeCRDuvXeCaE376Jy7hhhat0v
39bLoxHqBpUJtGnag6FD8V06A7VkdRIGCaMN5j6azha2hzFtrriwvfJfCgEmOnfr
ZUm3aCeMMC7Y2oPR0BIn0LOzxzR7NAYT13RAnov4lkPDYuOJlYbUxrjucjrcB6O6
X644G/K2bwLI8foi5V0xPRcbXEtyhucGCOUXy5FBff4bTRHpLpZgRit81WAGmobg
SHWIilpPGW7Qy6WP0FwHZaf1+y7rA/BnKfCWMDEF9TLYR5Hy77zDOIx7JKonCIBh
9MkxYE7PZ71UBzXLQi6AX/CXT8xUBKpxZMt7oSpvlteYcjrBq4+wa6L+BdSPUGka
XWVnHgmPhSgKXWTEtsJCsHfVdnCMG3CkKguEWVHMy32ReQuNMjv5vhkeOBQ6IlvG
aTolEq1PDO1K7lCRPP6Kucyr3AV4nzdFNjLAlAsZULxKd0mQfrWopQw1+kntcydm
PjwgnrerdIanruR7ssMhZq3AGLPWmX+ubKliyGsEvjBXtf85xRHRxOs3s3ta/zWY
riy2x1qG95+NwfWxUCisXSZIN1eQ92HMlHs8A8EkMYA3P9bXrM+xGjTJZ9x7YswJ
Hk9sW/FM2ZAV1rS9KvDcwgHeXVKnvHHc23yhvsNE9rmjolOGOZcAD202JbPnxYBU
HiegU7Gf05do4+42P5KEBygKRFBnmHJTBOFkotEKejdn+7/SVW4UfilDBiHH3Ixn
/2z7AVl1Vg+9Caeq83H59S0IaQk+a8Q+aI5C706Wqr4N8kTBYJ9Z/SeU4OvANh/M
HNU3TirfBGMAfbLGhCVgogedNRD/ggD2srispBNjZV+6GU28MsOUCsLfIPnutHR6
n71LCMiTllbellOjJ4Jb+MInDOB68GvIai3alARn8e4bfR8wX266MSkS3QbmLjRg
VZxdKAQueOh0dgqQ0Hq9Jr6qpBIHjHQpJY//ODv0FMNueYKeSufk2BBOtFPp6uwF
8qDta9RgaSxqRRZam2VGjc7vNntEmRxB/SgGTvMa4as1Q8GgNQXWIvJh//AnzZ3I
MlQZQzzTvvdr2WbLNyFgAdvdLoSRzv9cRLQ1mIaGkrZsRpptMQw6zA3+7ThOvl4t
umJmY4H9m4iWj4/+AIDRE+s724mCpa1k8L2sLijKpe0J9vCwjfUReNsVpeq+RyqV
7V/Kop5jpCYjH3/N4Cf7okA4v0+ijw6R1/4a/NYjadSGGe18nAHILn3JgOePnL+Y
HXXkYU+UYkzkS4ZMuL5F+PrUPtiNvjxEAGEXtO96oaStkzrYEfCaeZhKEomXMsOQ
obhu7Lfw8znn/hAb6pZ2INFT2ZhTWVJZyAydDs6qRkI2r+ez7E8o91tdcpCzqDaX
mIxOIwpuEiDWOI3N1/EmsVvJHZQhG6iq9oDIIK+vYk4BE0KIDlWhTVwv3O2iI80N
Mq376rLXcHg0Gu/wkMUtKZ712gQ0RDNTiHFLT41wISdUlWZxHdeyQuETuwFGaMGv
26u+6B94AqMGhW/fSav230L7RHeV73NDqsPG0u9pbAitQmVgF2ML68jEQjf8N8b7
AhEo+/J8DFq/GklLKC70TfoOSYScFhkEFnPflMRiNGf/AnsA25uIK9nR/sZlaFJC
+vzgUOzn0NCfiHk6JI4mYc9yaylr2fnNAEoyesTGNe1yT2KTKoazPQE1pm5s3R/c
Nj8Nwyf5W7XUvtp0HbGIprxwcw3RGPTsiEFxATVfJn/ms9vvODdv+3uzLh1g/cN4
6m42vGtlWN0tuiXI2K43J6lBVuvjgUwHYYqYOmXf+L0sh3GYU6ceImvusd9TbgjN
IV+1RJ5zmKPyopJ0l1ObFh8IKidRUnTxdcF/HFfzO5r/9kdxo3syym/k7Qlm6XV0
Z6ydQBxP+ZQ+ZsNvkUj2fUWrisWy2wCuVp3x0W4OmvFYWbN35wlgQTzy2bGyZrDX
ZVM39YJNtLToC2pG+GXvcxmPTd2WrcrSY3CRdTa/MnPweqanUaZ+K/WSZknp1ead
VLj9TVBPNJEGIfOI8eqasOp1zURBz5qvqJ+YpJ4v9kdGCeJHAa9svitx+qZe0uIt
HETU4sI/z6YUMBX7BS10hT3DGl8/JowfywZi1YozrNyfC5TsJD3jJWpJKtM/UUdX
y6AFUW4VKlR2A2pI8yKRdo18Deb3dCoQXtrvUb3QVg/IauaEy5s5YKi3FYJbQDon
ikPzGUkPoEYXEHviIgoG9IGPS2FIXowecBJBRIm8WgaC7I6xawpdxQt2Eg4VJIK9
7jIoVdF5ij8pdEdFA1au0gOrxCWho5SjJFblCpD9fiHrdY2/nv/4mMOk3cfQKcdH
h39egWkohywZn6jDTJ6mYd2JSwGPyGl7nlVeWh5/KqL8PGBCIDQofDVi4VwDunhm
M3rjC93saAwR3rPbGDYsSXFMJdJDtfXpf7hhmAudY6q6nWcK40V+VESr7FiT4zrY
YUO0DU3tezhYO9EHuMcPgkgG8ycWVLxwVIG1GEe5FuNf9h7/5ZVAIxCvqo4gHmvd
m2aw+N2zV7t1HW9ajYnzYWewZttZznlca663w2S6UbGlhTKEy1C5BFHQDfdc+FIr
2JInP/wzWegeGJEKrwquHZcV9ING8Zga9yd93APmPx4QYQFMcLnRNznZKTJV5ZwZ
OmnudOWeF1n3OyrkOZuCpaRElxDWZZqmP+dFqXKH8x5lXdw6Sk8pNW8VdmiCrqGp
sDy1J8Aql8fKEBvHQLM1PmXLv7Lvi+wK0Yj9lPfbW+ziU8slbORDXIRrOqRsgK3R
SwSRjo5mHk5Vu6Jw9P5vw0BSktfPuYJ+BrGAm+dQzBZXCV0K2Qq1MDRKCEVa2Azu
Kt0OVwm3gwiQr2Tuwl86arntyhs1+6eO7eWisJub/q/I2FVSqDq2PwPGKWd6i/i5
dA+RTJC2kWp+Nhp/kI3h2w15LVWDdoT6QX9HQ1upJxq3JtWfTfYKrxjYbENz9T/b
+0Yk8f3cSMRWcLOEbxt+NzXlkHzNuMpwSlecwFaQ6QsUvY4xL2laFWSsXMP/w4Nz
08/DHeCPMSfgX+ikohXfhVQqeSCkQq1Hpe5dVKvDB9M/+OnpkQU+OXuLV+MwFHFM
sosjS/cmaQ1cOE+NsK9wmVscTiVVMnLrtLs9Z0FYX1PvIbKBhjtqL6IKPVW4YdS1
vfsIexoTYhAR+byxcoDbk6LIA5X8z9O2K7j+BF6Pk17FV9ZhlvmKyjFYZo0stCsM
5axQXtzYreb+ZpboR1yu1Xe6zLkJEqN7ajfQx4JwRZ8n2X4F4QGO2Xhh25Bs4D7Z
A8aDqTCR50wW4GcqRgolMk6drcsATxO57pu6KA7hUvJG04Yw/fYEg47VATodMYo2
as3uZinpKmjuirCcOBpERlNGCRpBw2bMdupu6TiQEpIBqJl30BLXM/VuM75WA/Av
jsHsEB3NVP0TBo5l0DoxP12o0d2uSYoPBgruAtq1wZrYLwkb0Kn3jK1WJxjep5Nh
zLtBqN76W/UHvofkU8ojCyX5l+wYJWUX3GXgmXNtcpT1+kr3e+shKjKFfQMB/ara
3TUTJCvNCDNU4KaZpB60VhUJJp9/tr9wdhMu9H5WuPdCjbeiMquAWgfinO82LUwa
2pJvayv4FgOJoVKdD7/573+7LB1XNNVgIE9IV5PVH1AA4fgI53/diyRTDz1MX9ru
ZnCSaT3x8D4rKvQ1GtjqepOau5AUCi531vphLlgVqc0Q03esfYP04hYdf2YziI4T
bH2F5ZMik/1jZ+h+9O7If0dPIkdLCjGFXQfZ1ZZsgZdJvZqCa5sgFG0IoNCBMP/k
U/hfZ5SXrBhO4cOEFsn+IH8Udom/LCH0dYNobgPqlO0rdEhS5s9fKcG34q3pzOR1
9pK1Hnhz7cXf4rbDfq4EQ/nnyZS37IOhFbGTnwI0MqJ4pzstBGb7qB8QtC31xjsJ
HXg1pVioSSY1wOI1VAGKiBpd2gDeTzvTjVmYgctqSJ0Cy3XMQdq4/PGGRVLHcluU
JFOSYWouWG4dcP28tqcuDMx+34gio8TJcD45W1RzLWLnuhEjksxe23wCjKoa+uFm
7oyII6MLufDTYwUG7JR/1Shtf9gc08t+z89Evnaic+1QGMMSDkneWlR5M6TJS+WE
visFhPSsYQYlz8lTlQasd04yCk/IKA7WSt0+t3g753T/ruavWXVXeimNcI0o6VaY
HAoVXcJzVWXB50ekG++mUfHV1qgru7n7GFfuc9WzBOyv75LcBM/6LZmyucHdAYtQ
1rIpKqVk5YwBkLhs05ECEB+ynyHiGaWIxnM39oTULpVy5PAY+HbLw8UrqUDhd+ru
vT1yIqvl2VMkxEDiyARymI34AyTSIT9AY0vzbpAuwCILy/Q5mOdRhM76YrblWBnR
sc2Y5TWywfRMQfCjvJizfBs12NsebmcE3twEuSLnb4Ylx/vPqqKTJlutyv0mt+jy
r6AIV45qMaDkfQKwk15jl95qkXxl6ugvT/PkIWZkx2obv/z8Yz3AY9rQdM+/hALJ
Rf7lTB8/nEnCXOQ3/41xVofvD6urF2IxVT6hU6AlDmAV2PMTLNSpHVeb30E146AZ
pW6ii7deAup5fHs3FTJhPi42FpEuxKm2nez2/mVxBMeyAYo2JNeTFLi/L8w+Ka3s
a9ni35aAmcawl4AtrgD0Uc8Tbg9Vx3dJujMe5Dkj60sCGbPePnLAGicgUace+kPR
YlNMxTahvaRkFyp+KlMSjTVTYOkjCVznMWCLbsUKn4xDpRJBVyI2guiXBh7txRr1
gyZ4kEHX8zm1OBpE0yaTMQhRVRExgb56x7KSFU5xgukMA+fxZe+pH1PTtvLpWkXG
M68yB/BAEQ5+qqBGFumY5J3uJ+nTppuqsr5TBQ+Lmor/W01jjySw1rrq5C63Trlv
i1H0xR7QvEFJA1m176FDutyDM0HCXxRuxJM6trQ7yfItvx6UiW2eVE924opxcJvU
z79H+4ZzyY2le22L6Vhhq65jeSUqvWiYejab7kieNjRJbmsXdYRUEvqmGA9/3ybQ
8J1p3UmTyL4Neqq7TDblrdKYPDN5obDldrDJjl45/xPuwPgIzdEK9y1Lblt+qqmk
2CXtKtvVW6yvRjvO7um4RCWMVoinPuoNeVYmDpljpw82//3edSZKW+wWQfvUGPx7
WzYpKds68/pLE7cKWst1Jjr5MajpTbaJmtzIFJLOURvEwd5n6yo1xi0QA3E9jvEd
nipf26JXeEeqcqhCprpGJk4xxYZ6btP/KjPcF1SNPLH1JOz+j4xCr1MwI3HedWS/
ppGZzzAHG0vLXB95huyIgFSehdu3kPUx33aBYs1eOxwcs5xRkqzQs9j6A4j67nio
p7UGoOc285ipnHRMUgCTNCftxCvZqzZ3aC+eUkfJO7qH61CRQ/dgGRyGvsjwoeNB
CZB6TTiFR+khKqMw3yd8zzIddb7oYqOryAZzQer+Du7+9KVz+NUyquAr2MHuWC7f
eI2hSBfieND+TrvLAM/GcKB2UQfU8ep8UQvUXhPOaP5tc/MwZiqY3Ca6f/MrtoGX
PVZIiiIIeJBzs/5tbG/uH1xrUv+CKxuGlQdMNW3AGGc4uaWkt8GMdNZmAScKoLI1
jomzwiQtSgAQMECg2t9kv9/HvG2Py65nKJbl9Z6xQKbjABLGO/q1ERZPUV9HBaC+
Z2iQw3rpDlJnPGWRNRNzHPbeyhLXm1R9Es8WkQ4I9bddkTyeQWW4xpAkjPnLMUAv
buwy9JInEaEmo6ryEysYVsoachFty1VNQsMceW5WD16xPNRGC2srLs/UJZnVkfwc
vBPifWep0do9xTpomBT8ZRVGYXucQknKYxPJdu0Ss4krejtnlXJNw1O/z6ByuQEg
VolZyNt3bXipXm2D5rkvb5c7WyODc3wIxW5rvysGZGqcjKh1uHKB6hvwE9cCVoX4
Go3GWd3Nvp2Lzintu1y/+jN10DP/oISKl4xRqyy5Mse03mYbY7M+82039GbFi7mV
YJKGhoMc4MtBPKy9a6OggJb1HGm0sOgHwflxa28GnpqFFpd0A9pxkamgxLzbwLga
OyS8LssSBgX8VWFY7d5yQUVZFfMIdztn4L3ElT1f3yC8luSM5p56JhAtDu3vbE0l
ojwmJajynzhWspkRSZBdTcu10GhOkcQZD0+wtJ6sGZqQZ1JHJz4mNwR0PRI71SJ+
0q0j2Iubj0lWWvciLpG6oA8AERY2lX8+J7pXgBTghQNKnCoVtYz9lsf63EvhoANb
g2jc8ZrUmB3ZkZCWVWOWMkPWLJFcx1+NbY/hxW7SqIJ7gW+p2U24F2IvrsDLO/bF
T6TW620xfEAdjhHj2XTb7kM5/yrXyXUuypcmjpjy5pZRYw1tRiZ90c1mtsaRmj6e
wh7GFEJMjVUdmC95FWAfajhu/qn9VpNRdPrEvH4GoXburAwLtcWQistLvqlSNjG+
oP2vtYBodpwmZumAmaDe2Q4FfEGmftSXwUGRvy2yvMSwdsSCi/GugE5Y6iWTCVaO
Pt4zqltgQisk3Mxd1i+rGaTBDQwzc1jIk+CzGpepFcHQoEF3mDv2IMovzLMMUW4F
TEzy3u+87fqk+f/J1mS1n25ixA4tIlik15zrnATUkUJyZMQ4CnBi4B7o1siLOJgL
SUS7/qpvyeSdQvtbcz18uxhAS+w/HXKioJQ92jinGN3YaZrpA62aW9yp7MYYJJSF
rOmgPC7C5bEstnNB+LFiDyi4vQh7UKDS67tXAl9r6LrIWBIJ1FWaSXYqfgpVb4bH
RZlS03ZZ3bW9ZsyX1ZHSour2t50DM74i4W6afaJBk1BH7sevixAb71QSzDNVvXlN
WL2qV23XURI1e+3jhXqwn/m8wHvLM21X61mBaKrAyk1xSD6//mVCy2t2moaoTW8E
+5K6xfsdjvQQRZFQ8IdsnGsZR09mOJHWyLPxjL29ir0SrQAPE1v3RC7pu5OI023s
Ylt6FXalfnC4sUsZjCL39Ol6+0pUS0aZEYFJ0TPrk6LNLZLK9LJNhfTtfGhXCdv+
fk4/2aHSMB9m9MjE72+GzWYcYRzK7cJMpWd2NuKmnlhaFDP2PB3hqLo4DT63yaId
UP1HLNHfVfSB1gC3AFz+ITxDt85tyV55c4xN74Et+wKy7La88S/yKIko1aRclmtO
Xb6c01cBas/FBDP7OeE9l1ykdCJl/VvxI4rN494Jg8z8t51DwTVEoka8MDEn/lAd
CaVkMPJ/1MBlSmWIaGQiePfgtKZm2BkijdTBa+jeaPD5KsTz+1RJCJzsCv6kiKyi
l0PJEruM0H+R/ITRQrK2PchQgbZbLJEUq1NTzqrvfz4J3dKXWmr8Sy4FOsppVLoF
3blkiDM/5nwSO8SITfj2A9QdnYuRaUjtWbt6qbsRHi42TOOKg68LFbwzLhwekmFM
7s05sH1I3Ie0AGmDKpMxHG2QiHzw8Akw71ppR02PW3H1MOuNxsgkhFxTYaXNhGR6
ya4bdisDnfxKz8LXG/60dAyCd4naXRMHSng8/MOZ32J6p18nX2Mo0mG8UxNr8eni
7EXaiG02lZ24LVjxowxFHOJcs4GN/0XUQ9+mER3IVNA2F3RVSc6igQVQER1pwFfh
qnmk/F/q097N24ObSBdesppSXhDZ4nYbGeB7PPcraNhpf/pNCMIxh2QfJE3HiqBi
hrBxpGiMvdzfFWXPxbMlEnGuIi4A63B9YiR2Iwh5+xtSUE7Z+4EhZVQgy7DlYbq8
KxZTZ8o9kpgZN1VsS28cZw3X/ECntlMHJvODZGrr9PIJjHtP4g1Fzj1qL0Hho/mM
D3ujR//C8/ECKKzGatE5rRRB6Yys1EtniYjXHF4cbKrKaHcgavCMlJFrT8Y6OfrS
m0hp/gozKMchdRVSBZsNLFG6jbOmChgw3K+9744sEnfgtgfLFiIC6mYVVG1Casw/
bNfNgnG92uqIvnG1TQxC+DsFMmnK0pd6BcwtPkKhODz3G8LGsKeF2GMYnb3YHO2u
auFTZiDGmyDmfh9cT0oEqwYmE3Vcj/TCjFHDtBYoZ848DG2xDYYFOEoyq6s03/gm
QGR6tSiP65cLA6wblZ68Vnyf2xdqt9VJe0N9fOKg/FcBvG+4aJr7/UHtMjJebLuJ
pHD/6oxz5gIur/G7y2axzDI9Y307a8SgLxh8cZjphM5OZVtAgx41UsSBpSBaA5+1
XP80N38yRjZCd4b44oaoN6Un66XS7TK4g6mX8ynf6cZXpVqFZVCXK5ntXil74ni5
eV4Hug3ZKomk2CdivEDgQIj+7/a7alyvM8aUyDejEuwP+GTwxZ2mYb+CrFp0Fyh1
Zxh6sNvC1kUsBUdhk+hbUN/oCje2iYHDLXCRrEqqWeKDl0oepZp/yyNE1LLXbSzU
CmvMhQ6fgkX4TX8D9MDt+YW35YzTWSj7LW3z0YbekHIvJ0qYksOpG7GxCcIvlQdS
eRkg0Fw/LBx39R5zLuaScRlcP3x/NslzEmHcP00fhyY1uQCXAvkH3hzOsezpAgU4
dBXsygFqGY4ozjS8BOI3uDpEU+zA2FtbRl8Gn5Vl1ZBpI4mKwAo/cBSGHmp/cptR
CgrERwiyqPDy4p5RyJ7VLcKNgECWBii4x364UUTbbTYLsoc9UQLAcICt1SKCHwox
e6YU7Qmzc0ZZR3+lyTzYX9izxCu2dH+1RWgsCZL/wD0I+2sYiLkWj3DYy4dnMyVt
Tuejist50umeh3L+MNh/nqNtXQW103NkPc2WoSqPGlFFPzEV7LfBRbhX62qlwJ4H
7Tvu/FMEHbE3T/g8SHpFYSuJs/+efRvGFQJl+Nbh1LjVzYrJJLBK6V8W7hJ9M6eE
dj7ijs5tqAyhnZ2k6URmj6fO8RwK9YAndhsP7YA0olTLQlT7nouiHI33kYX05GmW
T+0UeHhNBtReZEHAvSWg7a1AEdURN4ZRleFUS/5EiJ/g3RTd5u2qQ90QMPHtkbPf
MXFSNLFVObs9zvlCjkmhchz1uUzxcHywuJWQ9fk0oWJuDrB3KAOY1B5RlFEhltdS
M7UQt9TKACdY7I5a8NnkUnjqCwMHsfaG7ZcbQyRT8GlP2DPwHD3bBFvvpcbu8YSw
vhv1aTcI+wI66PW2VWi644tKQGjdW3EWkm9ohbvwFr2/V7Dp7qMyAJiBgDRwINZG
8eMfh3ZCScKFpLm3eO+CCKJnRrqX3yUGu0+xJOaa28/uDNhMA+NaHpT9fcUcKGhA
RHjoAG/0DnaDytL7iDadQiMG96sR9qwlgFnkogT/aRJEfl6DoDF5y/Og0QON5sHi
AkcDcS9YELbhtn1a2Y+3bQr3q/HM8GHd9alZZ0KOMZbWVXFDqeEQWUQFN+CzeScq
OkySuKv60Ts/bZ/6V1qTh0IJX8gG5cYIvv1Vpei3Zb9t6jO/kTOb11BVBhZprUeX
e71wLPhxnc+y6UtRl+YembFS39FQ5I3uNUxgBAOZ1x4kGZcARdb1OVo14GoCr0rz
2D8lh1AkL6viLQBN1HZRN+mg16txDjK8FYzWaXFDYSaZ62ApGWmse2biYRfA8mS1
flxIPwke3o0d/u7nCRNXZ2vIQi4iVmDWeGxXZ8O9h1H1+wuvXYm6mly2PG8iEzcI
1z81skMTcpsaL7LrqVuS/p/bCWfO6XG+RqBZhstXFL4svXJpFmir/xJ7n8q4A4yn
Ksy59ATXKgXkGKXUOSpgl13S1uYFiPN+B0K0gkhnhfs2D/XrTHNrjZB4RFfpdX8k
wMhPMnPjs0BZ14jopSENfv2SLsf+wrj8xUDesmZQKZfhFhyQKxHTkKCEeyJKM6m+
lOzrsUfpLxyqZkXb4bysnoHus98Q7rGJfyKHAm54gXWE6WRebpjMe0eU8UakxHt2
6Ke9zqJw0oeA0dTbvnxmnMg9+1kuoqZlFXqX7JmcpNUgfAHoqch9jyFdG2PuXap5
vZEBIonc7lZOtL73n+H1KVIheTGe0aI6JT59Z0Akj/UAhT4uIPIjq0Rmb0DW4WZT
ElVLCxXRaREg8ngXn7rWQoaxnzIn4vE3V45QevuHSAf/j+nCQSvYBphYLY51tfNV
tsBouUuK5qpD1wt0llPqr1u8nmX1S8qB0BkJn7xYnfjiAAX1YFo2fqlf6JRaogXK
FnJ0xLEYxCBxE15HqHBJtb9Ie/Bl/GXZoGlgq2bZjk0aJGgVvjzil2I83KH6RjPu
9IRQhi78hCQ8k1Wlbnp9OI79r61FrWCjlzn2Az+0d62IWqhXTra5QmRh/x9vKpjh
QzjbRu8b3jB30VStUaFNCKuB8iqHWA04yjNDDsCQn3aoBufbg4UgSFDLmIHzfMOj
qZKx4RsV3ZtiHZx5E7o6dz2EZm85bxh5oUZiEIixJPe9+ix9nwqQJZ83csym7A/r
xQRTRafN4oXBBwWAPq6r3WushkusTvcDz5ZFctJq6nz6R6BO8lSQkqN1cACL3CbL
91Q/LwZoWMEkiPz10nAZ/PykG8l7goVc4mqF93VV6xl87IahpqEX/saoE34em7F+
lGMoI18h5f9WXfvIXio6I7mGNyV88gqzzMGY/SJdOIEGSHkX2eoOtswmc8DSmgZp
4SGiQrW5BBdp9qMRfompdwcVhJnsKZMPbf6/rGQjjEJ0Rog96LU/CkTxbHyIwpUa
Vr2hQTVV/qYh6fgs+BB9fW2lqqly2O4U1eRDIbc6e2U9L1UowB/K1RVYnUw+TTZy
SzPOGqd1aT+jcefgrW+hn4s9o+Th9TN/Dx1t7eSxdBhjhmUsgDqQPrUlpDulODhU
WiN/aNovKMk/RclUY1oAncTnSSrSyLPAI1eOhyMa2+FglZtI/8GUaFDhhJFqqYvm
P7VQeKgDggU8p2aNsJRFPbgCZx9RkEmJvCf+JWfBr7Efdjuqpxe5RL7hlozlPrp6
WHBjG3fTh+cOJVbC1GTKy9zvvfHOh1HoQEYQJJvQ67llQyfueZRwUrewBPgakkIB
N16dg2e5XIHSqrZHtlBK8q352SecGwa/R1JNhRmhyU7eESRg+LIbEmT8e4V4CmLi
+0QjgzFHSpJ50la6iSr2M8MPF/+0zlgC7g/sn4ng7bms+5AeWB3AL8mvCiCjVPXq
x93Gc8TkBlV+YtkgwPQ2sAJOSG+GWn59dylt0fkv3ejp1hKT77pmixIhrL72z0pQ
Rnsh+31qctzYWfGajwip7xrVJWUV61ZQxNH8w2qdWTA3X143yzrzaZEGa++qBAvK
Ec86YtnfKrMAE2i384h5cj4q36TK8TAxRAqgQRtWZijycL7pNTFpNJUV56iitet5
+eUXLQxAVbwe3DctkX8fj+1UsObwpUSQ0kXhC++AqIMq3OceOJfGYRDMP/qnf+eV
S4Q0U63qFUzHCDvyRSDRuqrgHW6XHHmiUKXBaRaCB3FzjBPa6BtEctFcGr9dsu61
huKNNjbl+/FPooLBTRC0UuiJY4Kgw65TTwTLysyMd3LZrBS6G17M4y3M6PXvuklt
oKYgQb3id1MdWoBmKL9//G3gr1bFpX5PmhcDptyX9aMPXFa34y3GzGoR/n5ZQRpa
oQa4krEg1lzCdBdOWR7moksWIcCJ2t6aRWAa9XnXtRuSlR+6ZHv5mtwpNUNU0f7h
KuzWXf7pqCuOBGmCof5ojJR9NK4yBhxupUBkrcfR9IkTUkWgQQVh29xcj48FtFXL
p8wrDDn9UPvBmsNLEjv/H18hd91twCHZGrsExEmyPTMnJqMI/fQAhPbg2R0BpOQq
C3Fe+wBGxsGgdvs9g699SXubUBun2BTZnna7sPZI2LtzGlx/lH33eMRVgN+u1g5C
5uWjK/qp48UfZfbMuySlwSiVdruubCZnPpHUrBRH66YlM0qXSvB8TrMdJHV5Kl6M
dpw+A/78JDIGXfyf3IE1WiL93iJDFy5gTuvJg9KKlvN5Aw1/U+7FDmTI/4gQmfnp
6npFtaYxLrwuAK1GsQv1FVkgWCAGNBZYUmKjwB5XMRZ1J7rPCs+3BijMQqFpFEzG
WfjDFOK+T725M5tYQgFKKRIYqAtEatsUarqH4fCD5TI00ztosLyeBveBX27RUmdb
ViqIMHjgHWlL/gmemL0a9Oxya0XckCwSd0ATi8WOJBTTkKfw2eZjyxxdLK5s3Om6
8+UoHu3/j6UkHOpBY/VMHCkj7vQef9pi09Bf7NIQhynys2qfAE55bjldKVfK8gI1
nle8JvHdIBAUnq4GRMnhe4caVMD24qUXD57cLQ743sg/iJ1NC4P18UwdC2MFgpqb
uHb7dFq7jTKWErD3Dr5peAcmMQQ/VcZiWEdToyQpt+kSKHkZptjO7rWPWSyzTrgf
QQj6gqKLZzDGmKcnDd5NXr6TvxCIWXdQrGF7z+b3qPI9ThY3TlNv29ysbupO98kM
pxAzlG0msjmcgs31V0PQI5mzHivx2l5G8+fwP8dXXYXcjkTPTKwHg4vShzVKg1UY
7NUjwnUgEIK7KUvDKdxkdq3hWVcf9ua02Tpattl4QuHuuDtwBZN5lRRnKGInCugC
wRQzIHqRkuFOKSRluT8j1Fih1XC8wt+4ZuWwwf3Rb28WF2BWJMN8+XyJ5o0v0Nr0
MjLZfRMQq/3ZOh87Cprs/kjmkq0iql9G1QOLJnJE8tpiL3tp63auxQRIFtcOZFTU
CJhf4Y7K0xJ0x3BP9ZA8GrW6286uBzUR3wDmr55es2O/0nQcpCZfGYuDcQuKXKbD
fcNWOzHExyZkObG2zPPDcwJMB4tUnhLcZ584AnVGu0wsoa5WUrFBVRxbdBKvT8/Y
1Qdrz8zR54v8Q/JNwa+pvi9pLP3gMOmlpvoQ+OLkaWtkeOfn52/bpbuQBr22zg+U
0HKQmbO4uYCuu3J9t4n8Gx9GiYpjq/wcTk0gxPW74H8c5ZdT7pYKnQKHERynlyCG
VpaqA2A76fbwj4isDTr8UwNmQBHda8ie6V5+jsgoxPMzqdBv8lGzPNRgzclDq5QI
pZUOPbNpbEt9kd1VJTOX1uJqiVjChg3szJXfYi10B64pmseTmdWKQkuPz1UoFYpy
Al9f2eKr3NxlCe5EDpWyUrc22YQ1bXqI1jdBBiaNykV/0HR2rp4E9+v+lZ0XDcMl
8hZfRl3exma+o9l1itKmY3aEbOLHpyAdXHwFA7La5kdqX+sC9CNibUXiEi9m9qma
M/c/GHocjuSciqQ6ihz4Ke1OcuUpFq/bF55goAKCHbPMGTsDc3dZ77mgFVr/b8Rg
sYNUyJsKaFz2RrCLb47k8o7w3glgn6CDlCUTEathQTXlcKrYGjwt/DIfdpIxfr3D
DXHZRJDfhzvQtmKDC3BYu2QOpCVoIL68+1jvqZ24FFc5s9a2VsxZNraHMSk3WOsA
Usol9WNsHyehLtflITmcGby51diGj+pXyY2vUIq9XHyQRQtlXdteqNFPxXjL8Pc8
Cm5C+t0lZJrGo+0N9pTJ9mRJ5fd4uPpTckdB7g0miNJmhMXqg9RtqkpTDtWJQB7H
3HsdqN3Szs4rv/x/xG+SB5A3S7vRa2cvlOmYxrw66OW3gOU/a0muvnQb2rkQ3ZBU
V+TaiYuhXynVVIyidUXcGs+6QhPSteyPjtPQb9URCcU9GdC1dj106v6DTAbo+JG8
djeDi/6T3xsK5dY0ct0sBK9dz6ym+x1a0n7U8J45HM1OKmES7b/ffgK9k3Wm2woq
Hp7thrmnlxQKVbpEqkKFMFunAfRTm8LpL5xAsMvcDIJ7/gwb3PK4gzTC/a3StXaE
eil9c9S5JHca0KzBV8EcpNLATutfrjmMzjFGfueuSxQqiOHeCUK2Zb1GZHIN14wk
vAfaT28gniiwUAPS9mKUWI156X1Lc0EBJIABe8XNVWrUkha0VI7s7D6k86RlQmMU
VIR7Qil4MMu5G6wJghxhamz3jDy+tFK1sNAn9dIYXxoGLE1Am3DMUuDTIAJgzWOA
Az1hfOtFSLjTRjQR2xxWYCZNrxLx5phiBWPalcTu4zkMu/oxRStgLxJtieePhH+C
z7NbFz8lIXYaaP7pHDAte+Fh777PjvHwBjKvarrV0AIZcY8zLgj7heLmByhhlyfg
GcPWsi2rUwwiGlBE/1xi5wHIyb1ZYeAa4MRfWfcFCDnJ0Yzn5AE7uciR4/rirbOR
XW2GyokO8Ja+VLjs95nuDFhTZdxVGYcsaRYP/eHVTVzmfeWCldTYaV4DzwK4UQxJ
vMTf0y9PAdpvtCQ6j301XBcZup25CzBNjp6C5hjuPqZ1QFRfIefenuLkz0J5bKV5
j53kTr9rYdV3be7vLR0Cb5L+yVQd+qHhNCcrzaNarFJtRhIe4SphGCwCpHLOWBni
sDNA/d6iasuFKupsw309VYxKHRY1A+jrSXzKm0kljq0T8Tvi2XEBcL/CFlPf5av2
dmTvufPop61DaCd4m9OsST8iM94UUj8rvev//mXTvGPZTZuaRN9JmdaoNPlJwLnP
S5X1GvP+Wkbre+S20LbGffwqSvoJeEOwGOq/yq10QxRklVFgqhkbPBSUFOxDyHdi
KM+Q6rSf9HxJsgeMubgz3nt3BxPu4BLNqo9zdBaDbMh7abI57RmSsW3UBF/Y5orn
6i0AGddPR1CKdHBSC+LC+okF6gMbZg5X8/iJN3L7RkZPAGj0Yg7zgLvfJT99jYeN
92lxpD2C5NP26CC4XXCxvkO5TCdQ4MX4G//Rqk6beKY2tX2+Qcj5ozutq0Qyyg5G
36z6NKVMQxEeuMFSiHFz/scZQZaNy9lJtUOxWfCZwfKSy7xurspj1Asg214nCBbf
Wa1tHZYBgRSozUMSUnURUxm6eOohPE4JStILM6zIcKSM65fGPrSz2tFx7weWRRv7
wn1b6+d83Zlg8MF1rKgw5hEzmuWTtGWMlUYe3LDb23F2/wuJssMr8hIuDANQVYku
R15aU1M4LWOwKMSwY7M5W9AQ8yEHrq1nLntIDzRZaL4WRBEwudQJ4uGgch3MpsJk
EaWyy8DtTe4sZlBLzR2UTTzvBS+6IgxzoHsxNpwDHVpPZyr7PZFWP1QLcVlTW8ZJ
9tmDrEdwQoUspJxl/BAnlOfTAtvI0nicp8BHOFnZR8gg8qWmBayr7KD5WQiYCjEt
frGEMb5/D3I3j515VcOisC8Vdc06Vy346o8ajNKCrqSm8HnDnqa2fXGJNUr8vDKD
6wy0aW0V1pyavvGYJeNoY+bLE7lieUyTuqwQX2d3XzBhnVmn8unO9HOKY4Y/7LgN
R9iREPV/QndoxMsm0aToRb6jc4WIoDWzZh7X4Xvka3kiD3gX0zLQAJtWwLnaWXmm
Ni5CDjZ/aoqroSjv507L6EnyPY8FmEuZyEZdis2qU4Rh0yhp/3L50+T7907LnJIW
MaBv+XaJpdJcGGz19P4KDJ+8EYxYOvBnYrzFXSkQ85Qv631JfPslarKI2/3fBf9+
Te/V5GeaH2PM76JJX68vMii+ORlRTGzUfhMw9WgK+q6vnZobttRa+qjw3rFKzbHO
Y+rhffhc7JOCw3Dv3w11IxkhnMSGKwXUNnq5e/smabsccX7axhiaf2DqtoOXF5C1
sRpZm5naMurbjKVjFfvP3NGBQ6oK+jg+R+o1ht7g+8H6BBWBGGJBF5iuaIv7eqK1
G0DA8mHs1SmPvld8TH6vLrM8BGW60q2lFaA2gTVv9zsDB1mAuK+x1I6VJgZS/A6y
wp+V34SfVkPRSf2flUoNzD2rrcsqg0FZkTJbkzqd4+gaBYvcx/0mdqMwdkQIWvpg
hQmHVQAUah2yBCxqQ7ePW/oWdv9wFI8NfgtVGPDkr92pwK35AMQT27hoqvgckZwA
IuDaDKOdv4N/pGEQjA7ipjYsV9mEnIQ98cBP4XpJlAymf1UCbgimYDZU2ljNOHvl
B23rZpO0Onlunc8w2Vwce28vX9hsrUdur/8cRst91LG8+oFLxd9V/nTyb0/+yPn7
Lp+gxkw71L8zWQ8H6zGK15dS4S6PdKK8fydsg4ypC5DlCoK1uHJyippBqIM8tPov
XjXuS3GrqMLGDlNHVkkBoAXHrMfTmYZx+x3qyCxf8VR5AVYt7p+kQUmlPSjNKMHy
GpEJ2OSua//c3JVFLBDzWOs6r/BtEk4KgIh4c1rlBrYMNSiEZiuSyHhK6Z9rpGpI
xZntuqTILsPYFA8ISBOzP5Eh9IBBb7NHg8XC4y84Z6wKgOBy9GQEDIXlI0ZGmk1U
a216kbi/cIKJzmPNjOwJcMWVzHy1qcNGQtWX/SJfJVUbNmEtgJyMD0813RMoA0//
e6a6jOK8FRz/T5fl+RnoVERkDWOUtQhbEtkkR3BYpQiehfg4oGwbzY+MvA2k7MlL
xCkdFi45DmkreE392SDfY5wbddFppSuhovBkBePOEafZrZuZ/UG/JF7JAIAqKRKn
GOxtB0hRQBUdY2bgB2HZBL54iKm7JGzoYLw/0zGDxuU3AY9IKyO/jA0L6cSj6Nzr
JcreZG6BHed9qYko8C/PNwYye/8+SGy1aOTAzDeR5/DFmCBR/yf/uuNqwCdb38QY
N+uraeWxeFEUfN6rWFsQy5KQvhicBJMfMrLO7jgzgal/chk1KGWCqLPDWrFlgcfx
RkHIeq6Y8Qv91v8kQOW20DOWfkq4+8lSgvLgoLBqHDzEIEM2SPLkURB/JqE9+2Uz
Q4BKEAJ9/JKtPKSZ1tAli+Pr9pZtory6kk421YPGrCG6YTJcFKmEhvFKCegtD3KA
QECr1Ix1HHYjJzue5ril9sbHpyoE/pO9cAmXu1lr3ibNlRDv9WUCsUaGMNx8eUu0
JLKrCx3TpBXFZRVbcDNzt8YNnPYljZ+92PXO8yQzDYNcq5vGa3SOZqKnqDF+RnwK
fMo/sNtrFqSnDRDPc8xcZVA4292fZ9Ll0sRa7/0ELUYsLUAvYzhUOMNY5fXR4QnA
uSK78xpA3SC4A2br+JU01LCD3J3G+iTk4eVdvoyBouw4yx8QqTFDX80NcOI+ChC2
p/1iAKB15MK3OZolPZtQZcLdjtTEKPmu6RE90Ut26f4HEELjYDtjH5Fr6RoRTlUk
R5hZ6dlqZNGErnN9gq8UZpkqt+MlAv/N89uxycxlRHSSG1swgzBkkuI1zQl3vYs6
PX+lSQGafZHQer218avLT6Yd2ZsNeBBykzUKrqg+KmYdR2rMP2ZR1QZXaM4OBFBg
MdBWSMId1WfWb9kqj3J0S+uNwnfi1qNOYxFSRwK8S4wxYFpedAd5uNlj/5g8kulE
H6zfqh7Y2kSawJsOxiowO8ZcC2CmWGjtDlZgkkrOAwW3idPFu8AauXre+mJwA28k
XT0gdK82AMQyBGKZqouCa4Jh5Dp86O2hUJT+QJoAjgAeyCWl2nFCh4GN2dU3bcqw
bz3g6e6zBqy2e2GsfsaTBdUBkvVjMFMMAgITsDo/CeXPf6E6iqhRVefCSef1txU8
oPZqsbnfFnOsVcviYnaVy4ceCBa2gqWWJFTPp4z1XfBIHMJQwC2kvSFmKjnbZWea
IYg8BwWLg7uusn0I2LaOXpQEvs+MIi2h42/PiuQaR8ZSVZjt+RsEdk8Gva1DYAOa
wtEJ6TJTQigW5sXpGSCjEEKOP9Aigo4R6VPZEfcKdyAb1bYV2W/AsGuM9opIFHX/
jV/VJ5rrkj+5LP7/+TcwaYRZ2p+qgPn2xAtBOqS0XPpVnketAa8iJaZEAmFWdIwO
Pg8+mdGftVRDSMbCQp/KKUZCyaqrzxxez6VhsyjMXNqpRwpve10/uL8WB6pHHF4/
/uuDdJS639n8RiCJIoYhv4HSdSFPVxJC6gzI+LwV0h6mSLVIq5vETbcEWolN/j+U
4p7ypcE8J6Agis4mYlJovS56FRRFWCCMahdJCkgUQ3ww0v7bj3sq1g7UzQBXJqvN
tQ1yTxwzFJU2+jtVc4/i13lnePDQw7E29w8EVW1AcuwhE9Je1SMLg5G+ZRG83GsH
PlziYDUCQ58vIl6s0mA3+LVMdK7oYxZ5+2ImB5s8hKu5m7QE1eOk7kuvrW5tJjkZ
G+rmHMWGVu21h3WXty2E6ZpQyaXZF8Jf7nRVsjp0F27Nr52wP9NLg9d5vE7R62qI
JpMwHdo1FB6vDJGF2thvXcbO6YspikdwLv2QoFiFrxar3M2hh756F3OxV1qTia+R
JLsGVrOOgDqnTgw7miCUIy54r+wWRJehjYIvRcanK2S7gjLwLOnL2onOXGAZ47Ev
HULPGFxhTBpGYbsuBXCoFP8r8b5o8GBCm6N51QpL1befn08Wan2gPR4uD67+KOpK
V/b7uwlO0QmsPRF0mrI7IeQi78WeB5tkqUidL0gOUG6viB5IZfa/Vsh6kpIO67O4
7O2Ruu+FjhdKtcm+9AIxBb9ZDAnM8JNamTGjxOgv2zj8iUiXvL3Qp0sqMWBxteiQ
bIUXEhc1ngmLOc0lzwvugz8HvI2yWN8PfAzKyp778RDUTpFAMqamuRPgeZspsbMp
bP6UaUBUnx9hC2v7v2tlinHJwfgYIwtl55g0JS/se5Vtk6MHp2TZbOtPkM43gtlH
+IQ1jGmKbXWM1ymR+J+VT4TMZuAdRBvwj/9XnXklL5Z1NIoiI6Ubjr6ix0w4f/+F
L1svX4JAEzO2IIk3adTTl2guzWjeMKwokzNoewFeu39bgV69Lk00gwQjcgnk6lrP
gf5qeheZGAvDWUa7huaY6Q62Rn7DOfIA88ud2cI51mhtripj6Ky7fzb4CZOR2CUC
Nz+4VT/LzfD1boyUODLhADnw+L1cKUMikYAOYKaUlKSWjJk1lQ5vX8de+pgUcZQ6
peayTrnlmlMBKYiYaWxthZ/kBQp7q2VCn8T+TEerKUUlf/qYHUOy7JzAbvt0z0qO
onRh/P2moMfMI/JNxFXAOawQrYK/tNeLP/afmarf5piauvvnkknsxOk1HEoiM8Z6
qIXld3rEkUFnUTjgt7W+fV+9ctJq1L7Xr/0vIsnOG7e7MHE2ZRMQrjq2CpHO+jqJ
yV1QpWsF6aQ7GfOAaZxvAjY3ChR3cUW1HfGAVvS3sBRvLtVNvWG2kKgGvGIuBb7o
jzTwSuLhsnlMgaE8wDq2Y/MZylzyOH0+m2AmrJMxuCX9pjEV166/pKgZrBxoGToo
bOjMDbUgN/UvNl1OTtvDwtZf05RnMyorCm/eMhVQxXHucyNtVysThnZoWkZBs51y
9UwtaxS7U3W0+mVUtq007hMJ8RNDKzpBLqG9yuSeLVCruh/JmVWIfXw2kzwh219h
WRop75ULFE13JvaHbyW66HTtMJ5Pv/GZ7ucb5B6fBfjP9FdowHO2Cc0LvhR3xuF+
rVyNNBfMisl52vW5clA19zeXkkQSpUi2mJUAfLgNyzm8LmZzEOu1xAhaJOmf7/Xk
gYTbEO7xVTZtwGLa/QmDxATXFG4wZzBwuPyrZ4ftJ9XCtG2HqfKhP1uY6lnHm9bl
9eIbcJ9uSoBxX+WeTOmT8hjesLO27HHHFBsnOZITMzitJNeWcOvJg9PWXyX+Q88N
GlCKWFDlkl1knPHQuzDRFqtd5FSXycJynzycJH+k//lZ5aYW+9WuV1YhBs1zHcuQ
KM6HD0Yz5m+wi2zYAbS/O3zgP8LX5RUFLrtuklhRRXnpcAuUy9cyeMHHhYWFa35z
iilzIdrsVUpnF2EecMlAKlr9WuQt9IuwIPwp9yihAB8WdNAN7XM9W1oaNUgg3Vr4
D7kf7nMvbdO4d8swHqxQCZ99pZ4+iKiO0KXxKtsliXVfYuC4HhtOpc1ltJ3ceya4
A1S2uCz15ICSsDOeJylDPcaDJPduAhIr53JrqzAVPXb//m4qclXD90buoFg9yyTV
TJ0qTh6TXUmmaP4QqBSZPbpTo2tn9xiMW6iZJFwAhq/R9+/m+5Xq/hnEaJHtkwGl
qEsa7PHBMB97N7chOkS+FdN+8Rp0v61NocowY6JChiuyXiJC8g00Jn5DZZ8uA8gz
/ynHzzEyk8WfwZunEUkplrEhRvOmgUEQx3jmImoof9ttcXloMl494OxVbOuKkgR7
h5aT+RhEw9nqsHsl4luk3ZUtOobGvfgr2tp85rVOZLY5NEPZMTrSvskIHo3AWCkQ
F6+1mHRqUeyt+VyE176UvYoaSn9joZEQoVmhmm6MEyqjms9WhOibntEFW6adDij1
MuhKAtzGyedW55VYS6p7wtLdJb0N5EIbxmlFgAOi/sFyeKcGVgFeOhxJ5Tp207cn
PrnkVTpIkdxcbyP5HXbc1T9dONFx61+EsM3DS321NfU20xeYK9d29NwRkenwbjnW
kGMvaR9LHgvt6ERRaZ0Gsn/9Xud0r/jPWT/sUEGJ4E70VHBnbvdRoGHa7wkIC2QC
QCKmZ339Og0au28CWQWhfSvZxLO9+h/ERh4Ofmcza6mN0Zl7ghuloAa5wLJxyezA
oFpTvjQwzKIAI+pv11XTXQMK5vaeo2VbBBtzer6/q7vgYZxX6nmfAxdm23iiPgu/
vqUKdXk/t6j/Aq89W0sNGLgxAkkYFjwECUu445pbpZtz5TVy91o5Lnw5TD7t08SU
CMMBV0+bO/ZKCBO0Ihfn8qsju4e/vOKXLTZvlvsuAiWph7ji60RNuFrI7HJ7BrVE
/xyzzj1UPmk84wzOQ9mNAAD8HfQNRowFd9e8As3Ms5dVIB7n0txIjPDzHsXwxobd
N4ssiZfftYKXswWOcsSXhuMGN1d9hho7ojrODRThc3Y8cX2MQlrwURABMDbE9JJQ
LmB5LEYXLE9exWSS7VyTO0zdozP6zKj5+/T0g5TUpr9yLWt9WKgW6PaLQVmuzzWm
ZWT9q0iHEkpthsF3K9i3JMs1XNtaxsblQojiTRSupQzichA0YAmkGu5EvrJz/a84
m9+Z0SbCnL/t9qpvhQIRttMH9FwFL89GhAYwISe2/tseV3/Z+aU6X5SICN7BEhCf
c7Bz+8JrkXaDXukluq81wfAcc1+vKIWQS9hZ74RukqfXdjwFhpfgwLkMmknB2JKD
XVSq396wYwx3CXcmIMUTJfYM1O/yYy9nzZv0SDnnTpENzktyl+HFJjH8zdCq9Zuu
nEXAUMs1frsjAVqDydImMuxedyYZAZLGoih8FJJsj9iIJM0YG6ti0b/Bp+XqF6c8
ghSAUXUv1684w5R7XGLGePnC+fLLahhHI8tBy9kG+svCM9zE5G0BY1mEioRRxLZs
YOehKWDOzzCSCWCNqkJxMDdQTFoQQDz+BW7PGPAqS4RWSG8a32zxBJaLvdIAgk6r
ZXTQfXNLfr6A7CxJ0jbkObYHDHUl8PmxRhOQGJZLROWUaAOOWopXYTb1K548y1kA
ZZfYQlEDk4IRHEvv5cpDVQcekjH3yPi0hTpI0WVfQOcH9AvazTfCNPssEfA7U6xi
djPsHhoJ1x0uiqSWylaWDkDwMeAtdboZIhLrI5cAB8I8qUeGKsA6gzPeg53SDc1h
hsI7TrW0DrWde3O8cPeR4Z21gSwXHslaalhNo/Wo77C9S88WK27EcUE1kv/dP7P0
Vk7bocL/PyWi+uE5egM/MNplI/oNEIrhgpxQ4zrUVx9HkimNGjemNXn5lgWyNLx3
CunPhCX3+oUZYIj2OTCY1CR9F5zWFr0dqpATJu2v6STfZ/2LZjzlVz5nwFITOt+p
J/xocNC08CRMiJBWtxTcGu/sli/C7nIQUCVbELTVfb7v2owt/FQOfbecTiPxW2oX
lvFZ2Kw3C1BY9oNyLAxLBjxiSv3zGCiNQcETYLCCYdFoA664BaDElbBywFIoNAHy
fAlCLQPWDus1Xaxz9IpF3OZE9Jbo6k0ts9VpCZ4AIWLiLjs3EHjlV5M1ek2tyP39
K3TH7wGVTBHsoM+OfVuZWZJgkFGokk3lg5w1O9wXLe/4MKEHbe1gunY18dvo7MNY
NeBc5/s2mZ/icQrkgjbtoXhWwOu9LvFTroltx2Wrymq5afX/owZTw7yyjci47YE4
4Jf3ZAO6doH9ZpQNzxC/YDzXd13U09VwXLG83m0GsGvXqkL0jipswnK0BDmni1rB
/u0AKmS+exWtaZUvUttencx++phOGTFdkK850dW/tEi+llC3O7FAC2k8jeE0D++M
L21rrXSUvW261rkvwUqCVwdPYkka3QoNqi8CSUpSW+I1KenwFNHFMeL2F3/gTjh4
I5GnQndRIaC9oiHg7MidUvHPfhta4VP0GZlFFUcKpcLse2l7kKutfk3X+ErL4+lH
tSkO8uWlxWak4RPcTHOrQBsOpW79GRWB6kJLjTKXXENlhAo1JOUVySbXhJTX+1uO
KBkG2FGyS1fEI1Q/8sA5nA7BvCXruNnVT21yAr09ku2DYmubieC+hAh2QdhKPGJL
6VGkep5I5ojqL1jH2QY8dhAA1yCA4C543LvYisI8FwY4AAjspiyrqBGaDqwehaWN
CpGKktXYlzLyIwBzueXvUwIQid+ZI+qQLPNcLUVqQVvHvZjRlx+y56TJ11g4/ueV
Qdac9cdUaj8ktoKxMCHGKFvApwQ8l3oe+BQjeuN3pdz5cjmgNSqG9zRXRmxKY/Yk
OKnCx0PWeUZ+SsR+z8dE+tAYc4lVqBMRFb3BwpTqG9XpO3l8UUbRHcPdX20o9Utu
8pLVqkrhM3ZK70ZJHahmWSwOMH0aADN7SSHeNQe7ywDtfI0DoSXluhNB58uPb2Ft
EdAiX0jMdz26TjLM4ibCQLIBGeS5GoLSZ31ZnySDEkqW3M0GXm6nLsaPQK7EzCfu
uCpwdq8fRB8jRMd6NJUnKmXb8E652DABV2xEtNC4Dh41APYE1YOWyhhX4qpScibp
86DZNKzgaOlJkMMNynk1EvTsX7RXDFRVW+QJgoJdYr91Rchf6fxhFcco6PBBD3Jz
wrrxEiE+Wuoj2N75XvyWOPw+WSdXH2i8iTKzoCdrO0Fdf/XBH2eKOfWmOoIyumSE
wZ41fwSuA4/MvLukuClYdQR2L55h4V/xsV61xAQSKE7jpX89SZn+OLWyza28m4wc
Qd5LnvgxssfDt/4kAmnSDLhaW15pbFC5geVVu/JQKXoippUFSd/dHe/viKQ2JzqG
g/KKW2s8G2cCKOrX2YwzUc0eCjMzknFskWceLQEutsRvdjkJR+PEU+AvJayf3g0L
P7nyfct++3cobFWsbzivbuySTi8/5AjMMZDppPqISOpvH1C9HjQ1QkPn8K0DtHZv
PkE4TDoaWe3qe3WSCkuGFxH+mtEdwNRlEbRRJl5/pk7IbOsnQdNXb39bIepyQF6G
4ut2C9OhUbnb4dMau3AC8ZuBxwdF8eD2M/RstcbC7GkwRYvDXh9lMb/dnp880MMF
ZOiD+Sv1R8A/Y3CXLauJIRL+B8wCGW5i22cSZVy8r6vkayxccibapxjJqfCkTdGJ
Rwybwb28D9Wv2EltjGuW0KPbKM57P1DCLxjgNwgVSlY5DbgcwI2L7vuV6nlpjf+P
jWULT0SiTxtTgFhkZXVQrmtf9K3l4mHVSpdpiTIf6eTlBwUftuiZ/CUqnJnAIOBt
g6Ui9OgjwI5WTdDlZ+F6B3Gyye/45DFLJGEWce0qa/yFX6Ezdw4s2OYgvgKxJCcN
Gb8YGJ4N67bQwYBrekFX9xN2OkYTBpeQ6bJfw6Kg8tDZFz+ImxXEtlZixCFRexBv
bgAzzlv6O5yPAjTOsM9SX7P1WU+As0P6ELl0ev1SsRw/Phds7RJ+xQJnsQF5FzK8
Q6xAk02+AN56kk/DaxxdAUt9JE9iMQefwh+Sw9EVrSiDFl1YiY9jyMi7O3ZkXBj6
RlCB0MKnxM+ACpUaIAZBFENVXUCgdCE+arJsnzbdxQB76CwmsqZplGLonHSkoEdL
HF5FYHhwmmHx9Y6GsqfmiYueB5hwZIVSM/oBZsXfUPX8fzuZbugaEErVps9b6XGx
26F13ByT2li1i1+4Vtrl1U80zKuBq5iTfwgycjFthbC7XWf1wcgl4S+vSxly9c0R
Ir/o4tqJ6GfmBVEKg/Q8zu7C5dmBuPseCP9DHoUfonBUzBq6yd5BSflNH+JTjwCw
qS4jhV9UY3ue3OhPEGEiP7PDDfjfqqsSfmqM0YOp65NsbE/4zddfmtODtWxeHURK
WuDGtcGjcL2NwyrSMvP1VaNlULqBtjK4/0GolcrBov1RbT26Bg7WGCaR/+U3Mc6A
nAyKt+GtaN0M9CZ0oaaGKz9cDdDAl8De1vSOCThFjMvl8WK8ws1f6Xwd03S8Y6tb
ejXPFtYzwZqkRjixTC3OCYa+LA0SpvKt8s7ZTFCM5DhxeqSgEkfPc5l+P9on1aoF
AyBiIuo33il1dwZTxzUf0IjWbBsouIVomJlMmd8skxYuFmp32RQrH+/NCve6D8y9
HhDRtC+Z1nDEaQXH3/SzxFyTWtw7YtySmM8rCKn18jlTglLvjMWSeVcMgcyZ+Lex
aM2HjRL5wL3g29CsMU/nLEx0Ktrk1/L/mxIx+YD1wDLtJhujF6Ng3J1o5Perx1pr
8Ju39NYGghEej6B/ugmUxEOtqe8cWIdJuTusxPlLhuvmaDwrLKEFcQaJ6nB1CgwO
bZE+EH4frV9chkJXBhC9SQ3hpr+fDcFJlEVAuQh7FFjKHDGse0gEJZWmiEOTDfS7
caOkXEWEMIMhVexkreOygQIJVr8vYJoitpbWhMI9/Lb/zUFpB3V6rRZZjdFJUlKq
QsCJc+Hs383BacoV5YN+3L6oGQZtZEznVFNMJ0N0QD/R3gBmp8FhCAQQfopkFY0D
eIbwVcFpOmhayHffc9424ES2PB6+gteKew7ktM1iTM/FrKQoUfI9AZnh59IJbGeT
CQ9xetTRG/6H91MIqs3UY0fL7a5UdjlNRHsr+Px5Q1Q=

`pragma protect end_protected
