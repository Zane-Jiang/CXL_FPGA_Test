// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QaJmgy5dFJEVxRvsJinqgxj+ehsRV2MPOCOABz+mxTN1IDhZRuKknjMXvqF6
M8AErdGmffHznGf1obNS2rbtq2lkmTUwySnTVx93i3Fme99iwE0gPoyAwV8h
xQN51HtnOgrcSy7lFVEGWY+ZEuf6HuSwAV8YQwngYgho/Kb3txmRReQLU01y
TXAOgs/ANWH/U/QH2Uk7362QIsAoOEOfYpbazuCAW2eAceao86gRTnfP5U20
FCK3OzA/eEhXtmVVpd/6pmNAsdr1xGj32cbtRyQnkkWFyeJ0K4EtcvBqes6X
/llR265/40FxygE5YUjUdNAXZrnYebcBChqX3C/pcg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
htCIa/KcYZFXAwg3ic4yMqcbv/7BtlelqxegkYGvXka56Ov9Po2Ik03fnXlD
rDLmnWktbtYF1KT1DUXYAqHshMYMIsLIwUw3cLP1rfDHQimLru952yG72cQ6
bK4lw/Un+4J8usbUxVpOx7Cw+lOsiqgpHYBb1Y5lPF6ahO63sa42BbROd1Cv
lIpI/vXxlsyDxePN2Vfsl5fXKT9RIV1Lc1iFN3TN3f8X51Wa5desHQwUxDHi
Ff06A1CzPtr62wJ7nb8+seDUSmHBMaJgz7SM7K8Ete7cRlrQ1TL9mNiBxFHI
nX5RIOCr4FBb74IraI/DuMc6njDC03f5YKZX4XhbbA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VaIiOOKZnbjL/YS6dNVWmru0UpKPbDpb03IAWO/FhN+B7dYxEcRJ/Cq2mfhW
efmum6seUy92ht9PWERbrhDv7pB3fhlaFoD3C2XFa43qb3g3xYHz4aCXXxRH
6MxtzQHQlFgEAZb4/vxoX14oPYogHDnpUNTZhL1SiCi3ziFwWg5xXhBqXL1I
ji/24J6Wc96aV8+3uAnDqIe+sd5+SMKY2y07sb3mIwV1h/8J9aO2JZebH2VW
kgd/vsE/GpBL9C9IOYt2QpjjvtFPFBJOB1vfF0hAV7qMAaOwgdF877XPMMTX
gzo05RIABz2ONsmUj4jbJB2cJs6Sxn31oQqNUpFCzQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JSuWxjUqy6+deeZlCHTHZ03CyDpw2Uyj0ySQ6nBVyUTrQgj2XUujGcSYAKAa
6v/hqJIFPfFfkp0L9zQdWZ0MjMHtRzlHgh4PSJJve4f8bsE6c5Y3r/nJ+yHc
SjXB03vVANx8u/R1lEnAiRbHtK8gtNR066csEGM+svBopS3j76A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
EhGOzqeFEAxkve6epwZNa3HoQqduwnF9asKyo5ncPKnrhxdNRVswI2Bv6ve2
xl3QS/wx9ReZdj3I/jZiBKTEmMqzFEqqo//TSk8nnWWpGB+/ecUHD9ugF+mI
5hMW7dfNdPya7n3ZXWTQM1lU9XarBzTnD9IKGBcO2/iMsgp3vfhTrbMAwHiH
YOLyhEYZdb5ffYkAChfuQt1Erq7gJmaaaa5zRf2EWt7w2V8+T+3BpTegXj+d
QnQTij6sPFO7jLVF/EvpM3HVCUHfbOc5+d7P3fOB3cq34+XnppDDRfrpa5JC
mJxtFphObag88Forrs6AV+XWfZdHZIovXW07Lz3XSStuvXoZ1MKgLcrh/4yc
RwZX+xaLDsV4yuny95kmXJ4/5Mn6ao7oquUF39mrgRDqhGffe8XC+v0TC3us
iK54Jz3+66Qk+yE+hLdihzMrEQDgwGlNzqZMt5JqEtTxd2AiPY9gzHrfjBoi
kJgci8v7frh/v+G7AsWtGebScnE8jaoP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SEBFqBEO5AmlZ4/z6CnqdJxEEkjC2sfP9pBr4wy3wJg+6rcgtHPKwaIbqrW7
p4vLH+Eu0UNxmDbiiysxvG5IstBT+iHfB3a3BZ1VPmkcjpaHgRZHFFiblkvN
XY/t+wS2MPFCLISe2AnimNG+YGrkhSf75Crn0aorUt8RhMfUUXM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KnMorat6uXAOzUZObFlggQGQEceLqyAo1rPCt0XwXvWoT9jnnndttVwe7ZOa
G+Gb31KS3nNXT1wVRp19WCLBHiSiHB69Tqn6oUyZ5z4ErYS+pW85ZZ6fstB/
7mADzUpAX+p+rTGicZ8fJwQG/+VY+N72VrSRxygz1/itgcn1nt8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 237088)
`pragma protect data_block
lhw2wSQBiTZYHbrFcy+h7zEVuvYpnNMd1r1y30HDbUdf7bTulA1/aCiUlzW9
HC/RKAh4msZpr1fhsHwEmy2i7kh+Z4JNy1VoLY7KfXAPed857rqCSH7BQo1T
/LwRBp1tA7wofji+iYnMgVdwEbYNDzxBFb/KuKfkvgiTHcbmTonCAOpTK2SV
DDW4ZByO7Naz50dC+7rZh2m2dXUPQg3xfQOKNpYHmHx7UL89w4aoxA3Rh6Ci
f5XxZT5jac07yZXKdoagaqdWGQq38zOd1qAJMG2ZZqNXoaOrh75Ab3Qn/FlR
92lOayalPSwZfaxiKFZ4mqC/1TCjyQqv440IiDGkVJ9ZbmOmt7p44WnQsemp
PUprj1F4msPMZXjaz5qoYx6/a15A5Cjd39OU8ZXn3P/+p4cfpAO1vgxmaws4
4svOSdFLgdlSxmwzh2EFs/a/yU4DisPictVdV5XMEvRsTwWfrownywI7TAoO
b83WWeuGtoanIpdLI+qebrxhNoablycXCMavtD9n2yrU1yzzhrBP1TFWmxTs
YqPDbr18F8dJbVqF49vQ8zuuSvNUp3R993qec0eWFK9Pe0RNYpqHDbv/0UEJ
ZpuS0OopmNpzIj1iQUq/EA6JxI/vJawWBj2NkuTCY/vaXDOl/GQHHSy/v147
TG1WSa06lqDTD66T8wH/TawkkXqWlRV+ilgAC7t1FN3TKBt/RIQHxo51mN97
aLoRdgjTi3DL1riYmbw7mvklDtZf6+7luiGf7L566TUsvGtjRCe8MSP7Tkxg
Ts4GedeKIPG7nx8ojV/M6WqNDs6r8SDQDLBhHbU01Rgaj/+FrkvkMqJsQ27c
LnQkW3pndrlDTc0KipC+Ix9jNdbdP+7/xZ0E35C4tkiRuBDO9UdLSqvTBznF
eAM+RhAUSPAmWF6d7U3/ChkFnor8n+PKaGBrZQxx7APVfLyoGFVGgUa5QxVN
BviFPbn4JjRLZ+JJWaAhoD0cpOlxYV1y9ybuODmrY9zUKpAgPeGk9xkFsxEE
Rbn5Ba2u8jxWYn6BA+kXccRcl59bJva7QJAVSm5J0zEAW3mx8T9q1SvM8yT2
N3nJ7vMFDisytHwR4NqJkCxHvGNKo4nAOrpjGZlyi2X0OfkqQIi9hMHrE8Bt
cege/J/xq9MTAjKKvqxFdMWTYEsGI5veOrlFmHSXyIYMYDb4C3q3+BedgXoY
WPzoW7r4+lxNmDgm2SRkx0Mg9j6FjzVY5BFwgn3z1A4VVSU4XJe5VfqTxKu7
KujqzaGvbp8AQA6ci2FSkiB3LSoTwXBfFsCk76s0mr0AiBHT5pjjm9qBxtwz
MTJsxso7l40dOleOEc/mKhmFaVLOYHw3mrkeowE+V/XyCOkoLjvzNNiqWoEs
vTMGlhQZQ+Rh4FyIhECt3SuRuk6nh0z8Fth7zeFxGV8MXOTJxXlpmSe8W1eC
9erFJ+xgCz706pVCj+8fFWOFh/vVgTB5ILj3veO96A4OI3+Icx0XrXpLVaxG
DyslE5W+xycKOX0qpaBUJxocjaM90Di+DMopyzU8HVWif4zOMH0ZOipAT8qI
3R0MY3bYfuMu0v//2nqgWRI+/3vzok2gAikhMldYyj3orbUFT/eMqkG9vsXo
G1et+QgMUS1Z0M/+Kxj2wIZU82UDfoltYAZn2tqn2D7n+GS5AsIij12lMrOF
sbIkHpCrmULW+v2s3OWY+X4qUjEufshnrO9i6ex52iBMd1Hk/eHBPTV4tnUR
i/FE0sNmPNNYoqCy+ezAVQl5VwiwYF5fhomN0pNSRmCF7ZLosa23xxsLw/cz
PKQfxvUkiotajri3XKjEFrRYKIBPSg1HNs9oPEfWowIdj5zzGa8PjVftav/M
LE1MMlgzz2e7TCsUHjfioqqaphWIQoNNBlxcKxJFg/2o6illOt4ycjkGGKHT
aLn6ataROm2czxBIr3GqPrq6ic/rGxGRXyFoBVEHzGqHZzbccrzzG8nD7HDG
5Lgp2TsgR2cfMlPJDx7amtzbOYkvYSIzcn1j39a3vK98owPC3BIdy7nHKvW1
AOYNrnzHoBytkp2S+Mpz1YBgF9VNWI5tSXItrNBwAUfFrPK1oi+WKITI6nmq
nxGpiRxOgg5eREXLk9Wi0WK51h0+kMWKfn8icStrO65XLmzBw+J3UoLX90cH
pHRMoGnNmwd5CWvIQhoWNauIN+9TQjpN1IqRjJDfT5gHP1Ml4Z9yjlrZuTMG
0Yx0t6ZOKB+JBV2QtkbVlTn1PjJF+IYECfLGxVBnu5XEU223+0svAh20oJXx
17fzxtX+h5XvhBGkOcJ3HxVG6t9IFZhwERbhTMVOlEtPi1hh87Z1Ef7E04vL
xJfjU6vFWRAMgSsJJKiB2i/QCx5pC0J/3VnDozfTEuoij++acJMA5d4FQa9P
ZchRQQbCpzcXPI/hyVY/ivzbv9g0ZIwdwwj6wnjUJdvozZAdkcItKIveKAYw
vDTVa2KnJrsFsVidRNIiGO/K1cpJt45YeCxXwEyaZD7qEc26MVb76YNtV4eE
hXObM+sbhjnPB4iXj/b0r/NlQWOmTIcxSWMBcoJVAEvzklh78W38vqc6fgKm
JZSJHfBo1xwXOhLT2YMYgqMqyvuFwEe25uvg/pk3CUQq5OXh+wPUxjZxEndp
s7LzctCkIRS/B7Idwf+0skII2nAZGFm4uNjUMhsQOaPaOZ0eOmj/LNeXUuP1
Am+WN4bS63i5xju9PKevwPTAy5yZyEQkmAKLTre6LwBt8L+JSaKwlng9Yia8
VzvLZ2PtYPXG/a2ShZdsxVuIp0fUhCwBf+8el48LVGtyCHZfN//bggSn0T/M
HJnJ/eI/GTnc51yqqOSL9DXoHQ4uIzUN2QwDd8g29qtDyU5DrP8N3QXSQIYK
1xJyROFV/1OIs/qJCPJ9cRXT/A8Vsr3f/JNW5ezJKfvAVIG3tPLudxJB8Jzb
KRI68XxXTOiNpOSu1QAu5DnqlAzDW4mva6lR0qfKkDq1NpPpaq/n/DxnxbwL
wSwOiflBaIuEkalSev/PreR/qVJcDJMUOiew41/VEFUrHsmdcKyYCeho5fXL
d4A6mpncDpd4f+m32cWYQCWBgEy8BBBR6UUmcvFK/MPXSp40izpDGcG5CxY2
Y6jl29u/GBQu0Ds5oV9FCy7hsx+fKZJhJfPcvoBviuxVYyMrLJzj8YbiXL8I
Ev8cv7YvoDK76rMsTdiefx9hIeDn+GOQLjEn6j8AP2GkVmSpIoLv82e19LCK
Ss2a+zJ7Oup5ERVQAFFUX9JmBRFp7O8dJzQ3JuPrC9RqDbWJ+2riwKRc4b8x
mVA4q/rbTn2UtFDo5TDuKg+ivpFLpgHaYch8L5OgcvJ/fPxTViARbzapZlz0
sCDByop57JbIt5FBHbABY8QyxVg2wCAQUgA82jqguQTLyx9zAz93wvqTZM1c
1SnkFmPyTdv/OaZ12yuv4LgQeISjnsKIpHSGNerUsM/GhjAZ/o7482uYFISn
+943irRpPIB43fpkw6/ACx/RzgsGoKXcoKi1Fs7iB7WQZp7g6q5d0MxQkGnC
uRPM4Z/o3rbCQi3NisRCSTZtxMoIazWwgUpi6jWVTLM+3K+G8TvRFJATjKyA
l7IwYMt0UoWPYuuY5FlwxJRyngnkHrqTR9eQYk2nR0YHF/JPE4JpDuOZRsHc
1q3VsH4rml0q6sHC722e0SSvpcVMUzWY4ZbMBnzjXXyrDo7dIweIFWKYlDfQ
W3xrGgwcgcGfOIKQvf2MgWxRxd6+MMSHPOxjqIHKs0z7uQMPu3P2DRLKTO8t
na47DdZvkLFpj4FkNwnqjmPOUSgJvPCtu1BuoxzjmmUBC1WWTEqiLOOxoXdJ
dXHH3h/pQ7EdYC+nrQnlOrW56e7M+w3haEHmVuWZbVfRfirr8aw6DLXzJ+oL
bU7nLeI7zCIhU73b00T9DtxI9pnIeEz+LWhe+hNUZImLQoM7389HiUiiN7IL
GsrF4INZGDARbStOWZ6fzXRCxl1KZi804A96z6ijHoYbhxh0AEwTsdth4bxE
0+EvCQb2ifgJP/DYYSatxyFSDk20aPfoJkWEoqlhpLddcDmp1T1XL8qO2Wsk
0A/4QFedxDrzi0mMB2Yd2uNO2X4curUe/ALRQugq3wlNoHZEgkW3Dj/p5eLM
kz2iFhuC6WvKH7K1wfV0OwHu3Xcd4JpXWoxGPE9Yic+P3X49JqQZuYSJjTmC
V+Bu0Lbi+NqtSOtAumF66VKi/XblVLhTKv6s3+5GR5gER7owLXlD3xqndnf+
QjF0IItgVKqGBIh9y4puFEsEr3JLsHJqspsYVMpycFgNAZE6zIUgyTAS5yPw
U7QIuTWQmz1xJ6fvHdyQsa4Ecbp72Si+CP4qFyFm4yCTBpGJxdxZ6ZFrH1Uj
TKVvcpXvpf5AZArHrqQpqq/v2eJziAwdiyU44DZVjr2DDNFFfaag1UXiNjbr
hScTRewA/I89s4Pq0cK++CMdhVtVQeb+WuDnl6jEQajyE7kKNvQEi1ItNIo0
Mi8K+RYsK7nu0wH9LN92/ZGCAAyLMqqLSBHroRfL2OY/8HCzPn1NT1DlLdVi
18gNMq7CRTQ+6YqHXW2Pt72okbIk8ah5wArCOAmk7HXLKQ97Z2qv4LCiTPhh
n1xl5d7UCSOcnv9plk+rhR1XUxD4OIBfMJFbCqwlI808etBN5IXDaSO1X3dW
Edkl1xZFjd3TndTbrhd+VBaa5NM4vcDOg1czN13iC6oW5O5HAawYzkIJG4U9
ESIZfK/qWKqZf8S3Wn8p2MLtj776X025WANugTr3T7X3THVz/VkH5d6Djwwu
9w2HBeph69TP6kZkIobHoFb4faHIs/5Mz7e5o87957oQgegZd6JAQn1c9hYs
KTLBNhQ6BZNSdWwHF9NLmGlCXDhS7P+N5UvlAfMkFXDfOwSOneaC3Rcf2D8p
43OrRI9M3b3AEJJyJeJrAMKctZRIIw/C+NJ3eNF3eo9DpbHXJCW7lb8it7uW
yIk7odGjc7vdNcdFQoMjsih3uPeCqeM+n6bHvZa79HJBCol7CtJSQBxFqy1y
3I7TGGIg+vVkvd8bBFqCrzLaQZoJTibXgXhwdILGfk202W2JgK+cp80hu8g0
7iNWeNLCX8yZbk1lSQYaEeHoWvtWna4gDhw/TU+4BSIdJ+kW9u+Jf/rjuuWl
kjgtFfjUaM2ZXNqjXrois/TEZWY52KWcFGJvr1XiF3d4V8KqXy2GE2pbP1Gr
c3cV6VF785fiGbGMDIlc95SL/Y1TOhcrkbUS7bXo1ofm25FekoVH3lKzovNY
2p+RaWfF2lii7TFdvnDYupxq4v1VFGsQGQ2OpFN/esm4ThlcVL+jgTUdcSds
G7TFnXtNWOYI+8Udz4gYt8FfSLTUxwxu4QCqSRiV1S/sJhk8ig3EtFm3ip31
tKOuq4cbJ5frB/nlTJTR9wIpjvevwqiKWvDpOtowNaDptxo5Jor5QKj+ErCl
gFc+fqBvxNJ1ClQQGiT1Z19lUBLXdcE0nT8gr6xc8Ssf8UPxh+RyYGaUJBas
Z2Q8U9X1Rz7ORPiwbeZePijYMVzg7kLRRg2HWWv7XFqkBaA0XE+s4C9dw2QD
1lq8FeFmms6MQOHeFpIwLUYjVGDmwOI8AyUjOxBamM0NEQhZm/uqyZtrW0RB
Yw6WbCZ+yoAJ9uxqtPWRgk+ba6qyytgG+D8pmnDHoPlXJz7Q47UI3i5BvqD1
0GAR/ApiR136oG0WdnfYDG8/OweIQyiVwlaoSHBNp6R98fdDMV2eAHjcpllD
o51BgTdo0JiTZIBp7Bqp1aBEaM6fZgdnmtPgxsCqbSeQlP0qmDBy4qHZVqaU
MXTm5r06VWPzuMlVp4TZ7y/2gXNaLjQH5mtpUpHTuSGxJ70ho9E4kchJbnK6
AzKWYy0LCzQ3Zch1Gqyed8HxL7CPFskZDHkDQkN6gdpuYkKs58H5UDREBx0o
H0SXZnfQaivxzfwIue6xuhL1zP5FfM/cKcDUAMcsZb7QU1MrvukXvp0b7PQl
r2APahTUJ0NqjC4+idkwZHCjoj7kiwGJKW/ojlo+Ylgx3Tf8FSovNxgOcavC
up7H/u2YusMemqKFWH7i0CSw+cRUn1YPJeV1zHovYnfrBgPPTwW7QHVSLg2b
lLc6t22yPOPT2thjd+ySEvQhcmtu6cY/oMntjCfaOnVwA2oMFN/UGqz2zQ9p
2RXATf+U1IJjD6LAss7m7Dh2g4dQVUoADCgOZho4EIQxwZ7eULCohj7xmPqN
Qvo0KfolUzZnZustwrqYueahVJxwFf74c5DaqzxNu0E2dzukAFfAObfA0twz
x1Pjhtr6r4o2TFPUtfM849KOZPVrY/ZRhvilfsSezDWYI8TeGQ9aumGTO0WB
fOu2s13TlYh2w0bZcaXGzSFa+i+yvF1C0o6ZiFCywTxi+fpCe5aJ5aEGrFLS
Ve/cv+qy5YPSEE9/DemVMyw41baycnUtQ9qPdexsr5BnuaBg7Rlu/1kFUlQP
SpJN3LK2+nRZ7XzI+zn3AKOXrZKEZYBfxl+FjLr2h5yGe+TmaiSjuuZ+5S20
dBTjJ1fgfyL5+ZAKq+6Xbhkt7s2TYitfPUfVdQwvk0qOU4KvVkEFqpI4kVvI
fDimR/cx5vsGz08PXEw7vBByw+cYAUN47LlLX+oMfxKrynxRnEEEv/pNyMQT
3yB5NaDTmtUccaU3UZW0vHfDqJ1f010JdI1S9/+V8XBH13H3hgzobT/zeUDl
sDMM7blE22LhP01z437cuHLvOHFQupiqit0ltPhigZRUxikpIE9CSzQRA7A3
EqY76LsHnWE9hnBO7SFVli3kQHLS/bjYgwNVv97pDxQOyxVAPPGXXvUKpiK7
jIgOGPTte6chW2RyRM9baH+yG87epmROB7yNgJF1OfnJeDbdeAtv/7fA7YTG
aeWFuvAxd90H5g9Ynyl1SgU0lM9m8ydzXUZykmDpGf8IlojXgj+AiclUOyic
3NxmE2pNgRnJGnYSJmQUpnmD3/8hTKH0FGk35xPgHNcIvksLctVZFdsaJ4Cv
0AkjiU+bKCjJAQwDt79Xgx/cU9cSF23z3ouKMGMKkTG4Mlq+XB7HlOFBZRsn
tk9KyHK6zBNs4czg09pCM7mX5Nj1il9bI686o3F+GrQiX4FWWi80FqVb31va
joXIfYEoUvPlGGU+9cvgR6N2dlvwjSrnFEpXi5Vs9zhUImKp+rpIbVVYN5de
jmESjYpEH2m39tjpQTAaIGFcmCSR8w8aDCb+aI9gFgLanSI9PLne3rEHc1Ex
vd5dMS4sBdGgOaugE9XD8J+ZhNYTDdg5Lne7Ry8wX8MkWvICUDHsmE5SME9R
1bvRO0KAOYcYEPZHf35UIhMP4B58pR6sMadeod/02lxGFE/XIHuC9KoSEpBq
L8pF2PmAejLSqSaoioX5Zi7jUUo9DNCCTthoylo6ww7PnqIn7uLyL3fYU3Hb
4ijUfBxPpPsYCXYA0pwyuvOFYQ2fsOCDqPySUxpzu5DjvRjnTdpwYBWGSHvc
0122W09h4z7NntcwH/fRSpE/1PXD4pxqpRqATVx8WTw1zxyVtWnF30nFRH65
YErdRqG5IpCoaibudmvjb33iywQ89SU1ok/htTih8/R/M16YEqhF1ldIbmqS
Pg+u72YNs9iA6mR0WAzd5o+I+hMV0E2C0DfJOSnXJfM5GjYEphEDlA7Qr+Wb
8QFo69SQ+l/6Bv4MFstv8oLeYA0a1IXHq+5YcA3VC4/GTVFONCE6vg4VofRs
KRj8PIjaPZDM3v/CWen358q43xYyU+RJD0hhH59l/3VPVSdW7xWSW2b4F+E2
PObENGm8qhwm1ZIh/OHWJdIj2DmNUaN/6ADrAFqEp8RwrF1aZzZTsq8Mo8nu
6fGHjlODprvOgWVzSNi0WAPkwv22HMqb47aKcA4SmYOKwl8KyR4ItXujEPYu
MF31mCOpkze4g4nbeGmc7ndS14BKuCB48WJ28u3SZj0qhRvTAcP6oc3dcoO4
lrcudcStvlr3GJPGaiPfyCOT5/12EvB/ZIXGQ74xnK45hL/DkuFVBXxXGa3j
Z1A5Upp8ymPagKJqkTl4g94+X8T72CQj4QJrUawzMFa894TMXNJoBfBgpAcL
uqZJr94YFmPnIsh7Mill87DaDZYQKTPIMedykInSp/Ucy3aZYQDQpSJhtEWF
regHptcTBvbA+XmfxENhRk2zLPjCqjSb66MU90UVmzTfs0slkEZ+KrsnnK0b
De4aO6W59jS0ao6CLi4NyAWTzyJzF0wlw4biYc8kaXjrDOZzNb2C/wnz1kN0
mYLLYa2CexfNymzMsFTtYZ3pogxtUTrSRfpuyJQ6N/2H6+tIRpngsBEVZ6j6
JyPanltNsNpKHybRdOOthgaGPrktQD/hBaN5xzvI9y8H4IC3lVgn0wZ/F3K8
k7qz8xoyAoQFyKWQfi7XVGOvndij7SsKX+x+bxNMOMM8skP2gzbn+HCJ3PxY
OE3f1Wp+ZelyfwE/5ER0bp0rWTWpJeYJRYUN5g0IS+loRotRIj+z51GdkEyu
x4N9zSJiJOVpo13lXMSZbA9YaaM0ChN/znjCrMmiXSeaLaXY+cX13x+giAO8
n64Fipy4OPXrIa0ZsGpBTO91MhzvCrpa2aNenGviNxxyUNMB1BERRCMMpDOG
kWELYNkjmCt79EBaylBTIoVbzgdkqhGn3RTdg9XfbOUCIYuBzQ2sIID5XqKE
nt64lML5UanBMttE//0Q/51JzCmIXq/3Y92OVXZQ6kjlJY0APcGkmWBAt7by
kQICprYilRXWTtJ+VahpRgBZX/Fe6sWXZcqNlvBPk37k3zsUZtLeT+jMKxLb
yHbxFGte3nwM7Z5Y3UJYMATJ1BkrKmpz3xv8DzAXG7CDwrjKKSFrlbnnAHDc
o2jgX8jZybBhKJ1UfkBbdqQS8JqI1VY0KT+YVVRmPD/tMfU7fPQdryVF16Di
S1V4wwnwygyqJ/XHbuSaeZuFsEma1sllrfCf9z4vnwBnqLTLZ7DwFrKce2am
V7uI9shu6t4hNz3pMGH3g5iakPb9epDWeQ9CCrb77fTm3bPiHt2TCTpmp7cx
avke0GO7IGW4quGRI7QYyQez6+OhlxC2UlWBKQ52fuBD+EAdMyDmiHlzUhvH
Y9jxegyHrjSGufl9dc8+QkEkm7bkfo518LxbT+4NGX+VT8G5ZfbdWiUagSAY
raDN3LxFVn0BsVGan7wdHYP35S5H1XpFmdF7i70ecdwyZqmiuIzGuxh11Dj5
t8W621jdaPioKkK2FgHYfMojYeS/zjc5vyKdNS3XPRy56L6KuZSQhKX4wyuO
tj3M3wDRXp7U9a6n/wQ9zMoezvgB3TnKYegwL9EYFWX+kyGDbPo/YjA60k4V
X9qS+rwx2irvsSJ4dmMUS1y5EAomzzUwm2V2slo+GZ+at7JY87lH4V+0zQqd
RfuMJRFdwdHPXLRajrGuCM/D+pwLGOHeamALxgQ963NMxTGc9nnvuiMja95q
6mPDsvhiesT5iaV6eGHrvN/SpjvPaUTGsQChY418TfltSCmwWkXEHnwUNJGL
lDRS9mN6/IRKSemNJFSnZJ/NLpX2Mn1KTzQVUqa/dGc/QeqDbLjidjyejA5/
XheVEzZUFiYBrWkTLu6J6VWq+Xh6uR1KolzSyLpdghsfrCtqS9kpDSjoYrT8
AgnFzyhkYm2ldpwHfPF/SPcSwsVw/+wolnnv3psO0yN6ASCz12yLl3exYqkt
/e2BJVC+QKtczQPGvyxxDp223NKDlXagGvfYpGk8jvR5nlryfJehD8ctxOUI
BJ9irgf0eXMlJ5hGe0skg+sFokPeJkgX8BOn4U3cvAIgS1eHMA8R/soZ1dY9
ssWb35qzyEDfFzfCKFZKlq9u2RFMVsh3wsZVIR1TfqdLMZWd/UY98B4MPNAb
7EkydH4MSjOdXuyCfYzWJkvcN+g4Jt7nZnhexK/sMs1/OwAMKNwR9I1pqm9k
BSGp1jWtDIfIaF0AkFKdiCOwEzujs6slL58bf7PliiDWO1GC4H9eKI4yQ1A7
hIeASymXSCTHjpPK0eoWU5i/yLpiIYNyGzBgGFWmvjCzDi+KPUtFkggRlAuk
ntARCkgk/vT0YFSAbVTIVi5vxdWTbdAWd+i/4r/2tgAS1bxpjmB9YDP01/w/
KifhlM+H9xleirQPBUCC9uDri7AlwNQyBeoTvF4lPy5Nw7lqjVxKrLnCrQuq
+q5oq/+rH1kRBWTPqTP+NeFhhGub/tuz1BA5nMuCo2iM1q9xENQxscYgZ0IV
Rq+UsRLyvHSDVDXTPhf8MgHGEhbzSql9CjGGJPQFMgrzsCY5aaLAvqK4Rq2x
IVhXjh3wxL5Kn9d9cUH03aEbqMsvTds+diAOfKochTGBs634naW+J+LyyNne
9BROELyjQaiPMC9GPuadiEbEl07RmpLMaj170Uk/YwXXt67mjz4hlMcIPrcz
+LRankLLad/N3i9/hzrt0ZNFC1XpQ1+d7iHt58M3ls7awY6FwdoryFdrns1R
PWr7+UbWgz0PAnc3IsF4E2wUbOTaUNi4kt7wzdBqsv9OPgqGjYEIi88B2qk3
51fo/3wnPKlylNprFeSIaW2h5r0S9NVGvCa3hCqjdlpKay3oH5s3/L688bgE
ajIA6oFYFZd1UxSsfL9WYiZvCBhgD3jDdMTbNfgKgLVEgbQxqtRlJsZLr55u
YtbYJ7aurCSTEjQuHIWgG14SbYO9Q0GsnDXf+8pjgnn/Wwv2nOFSFyvhMbi8
4AoSLoSYQCwGIFSsEQ68cXzYTu3hYXKE6D3tG+Z2xo4L8nLlj7dxxxHgHzhU
K9p7A/NxY/gCyqOEC1QWY7pBKD4El1pEjhNPAo0OZ/0w3FRmVqbRwyFLrShN
UrwB6LT/OtMz/iDM1xUtmcId/mo6IkZsms00Akt0B/FLM6kG77wqo69XLo7e
zv2bYZ7yYifFtPqmJ49W7YG5cLdc2HgyzMUEdGHs0zRVSJ7cNMzrKmc0iBRO
KiCoSfujdMmRpP1vimrTBjiMFMXcvJC0OoyRBUSIYFJ6rmOm0mvYsX7eOaXS
RGo8I4vQDsLCFkbr0eUytsjiVNSFIcoLcdM4Bkwif1HCDdubww9rNVlip3Wk
93HpTVFkW7AiOxBUuSJmpeMeCCxMBZ/KZ4M2vo4EHNFDj9nV5tRW6NZ9E0UQ
py0of12zwE+WM27rb1E8pb+kJcdtrhcxXix2i8yvwVStgcD5+b/9kr2yqBdx
2Q635Ar9BGIDWmzHJ+OXaborvgacvNVOxWLtRWjBSv1xsP/bWLwUvIx3HKvZ
MtfUQYDElA0LMhfL6/+vyt5CB8KE4S5nFJ9haJK1uQ4XBfsQSkJA0qiGeAvz
gS0TQn7y74HZ/yAsgigR+I+TtPLyzX+VUL3wHvS4wDcVmHaIvYTiMag6kD8W
5jOVm8FnQnzZu3goNcGbbWnPIYP6vQPPHeabYJ/Uf2w7zhfT3tCyK4vmUTWT
RHRN+ATyPFxbrI7AoYfTyhhezoM/n35AdUGLS2Ob1n5AxWwzLTbza4ZZZaZ2
7FauPuljhN4warHYLgPav7wzD8mNLp2EiVvb6Du4HfKLAPnZ3+9+t8Ff1GFg
Eh6hxS7Od4iIxjaXbc91+cipVvO+ULJx922O7btf1N5mm+rZjJ7yv4IQ8Cfy
dG4CCHDdiQqJQjwy7Y09vZvl+prs/cNXUSbTJ25uWLq4Ax2de/Ky65aFWZHz
5+ZYq5grZ7UQ6/4aEfCUz0FLH9a9WoBad0C/4VKoRBC4E0r8CQIiQaXt8+VT
719/ol8SgdQ3gLOcM5XVi/DI9O/dW79Ia2X/9twKjSRdRAif1uknwRB+zkLH
zJ/PNtrzDxTmCncwUwSgCvOAPVyGKwbfSCNmv8rwWsxutvCA/TuqEPuzScx/
/5EY+RDsgXAKz34VcCvFsuOQ+C68BxBr9B5RftO4deev1ocVV/XQdRWoR54m
QmNAIqRyRaAoZzMiRyut+o2auoJv/EFa6oWPndcRFJbAoQyrmZsT6DvJIA1/
d40CZfH5/6DqdLorDfpMfM32cxliXfwzdxPO+w7KsEH8NHskvDovSqpEz6+i
Tq/Vy9PCB63hhavokS8PAEcp7QzilA/gBiyswJu/5h92gr8miB+pg5f30hy0
PStVHgOxZKMeSTURqWkxmwq4U2RZfDT2CY8DxJTxXQOnGU6gedAUQQyekVWL
Y5M5AWzLXM2Z7ibdQ4nfE9Jyab/qrONlUMDf9oOTa25mEULrcvDyN2Jy95iV
c2FnrLAiHlVcM/bolfJjNDAT/yKrBhaDNglszwDpSSb3eWFVntMdb+kIsyNP
1FiQ7z1cJseBtCsbrUQwkNEkE4XfsfQXvLQozGhdZJZLxk4o7eRed33DrsTD
dX8uglEL3ZD5bLRUD68RmKXJ3aoH3S2Gg1XqbDSVq1b6IYB4zES1KO0M1rgM
PRpoCtIiCd64Qn2DOdKmmWasqAwEXBhJ12LNdcsb1q8m5t7TD9AIFd5N6n12
/SVH5zxIWf43QyJ7IeeJ7fp33WJBLKkJjOniYb7AXOHB0wDU79aqYaaz2X6c
Bl286PN5hfbz9ZHmnWEp6ejAZw/A7cKGYeBO2a7GsphtJXvsCWEHHkgPy5d2
LmfjAP5g+K9YQMxSRj8r4TTNokj/7GQ7MwTl9tbQ8sa2fKl2CfKwhqfnUpvG
4Qz6iiGeB/bhkFtwFqvZqB4yfodx3XLkPC4AD4elhv65fQoRN8+ZdBlqfgDg
RaNWZBJ1rkcspVIpNKdx7pWvZack6yJFSSGjkySnYwWbLANj1GnkflhcL/T7
e5EpuJthUds2/fnH0CzoE3wEWvJHzNGRKJhBoEwkjXhIG5G4IH4ePkVlQ2g9
hQh9ZJcT/dsVn+vm2ulMX/hHRct0YDw2DGU3wnOGVbdEpvBEK+5qZfU/Ba5T
spLnb3vpPySgeMrWI/vmiwB76N8FExQ039MaSQxI00Bzrb5JbzRdJwKq5Gkv
+5Xy3pql9MleEkX0+ADLuxr/GIqq66vi0xSTw/0GUZG2gk1iQos/j4TgysyS
Ho5azqTA+U7bvIItulPQYHhiq+3ZYaL7Q+Z56+WK1cQaTZCwkRKe4F70WPkp
/OnkGCqOb//YuzieL/eR89hla+gjq4mYdKCOBLpFfq+qowdnl2bxRdmGL2Yw
8b+H1Px8pE+QLQXFiuxfiVJUN0eoUkyCmMOlyeqMZ+ywkevgdtL/qd3rfakP
C1EZSOlXClDnTFbQepG2U3niRgO0iaF7Tqe+QdVgyv2U47FIsk/M/GKSwtsR
jKhdZF3SwjWRH+ggNrYFE7/GeCQxNCmH/os+oqDERLwYrGiArVdnzU+p9fpr
4qlVS4Yhjb+KiuiMzzFbfp0GWlTBJnVXOaqQgdHQ+GHVaW3Ai7e0azkkx8oC
vDG6j1cgBYnvmX8pnsZfUaqGu+jzfEwao2qgERsL7+6C0M2POg6G9smyyniD
e40Eord9d7cigGzCB6pxHQuEuAXDW6W4ASByMb9MgjsimBdtwbdVgcRHhZmf
Z9GqteJ2uUOoTnaPowu2uEgeee5ojpTuAkxzUDRvMXfjF6ZZqTy3EYMZWdff
kUAnMAqUeMvBLBUG/0u0eeJHaFGfRTOEzmo1jfiQoJmD1eOiKBrQbSC+QfFe
XVAMmJ1Gg4c7XapgCCPpLoFqxz45vDWlg6nAsqVdoEI3o4KDha5nkZ+Ivumv
5y+W1sr/MRlodgCUsXbxGFQ/SaUZVS4bnnIAbtjoZydI9sd7c2HNCTnTG+Ta
OoC2XHBkT2gbcIwwT32LdVduALnbFWRn6xHIfB1YK9LIe5r+gBHhF7+5F3ua
XomqrLhKOznjN8vEk8yG1tRO0CbxN4NPU0L9Y3yqMeBHnBYd2jH93QxAHyee
eovIY7lcFUOqYGo5GnzFhT6X8KxAOO/jEHfTUI3RY7flvOt3GOV9rK7ZEldf
MwMWoQOPgscvf2jWeB6ywwQKz7HufD9tcM2xSZh9ac9kWtOY0UwBx3zmkg17
IUMrraaCVyGN23RruaFjlTnu4Zm1Si51VQEnUxdxTGJaFJYlGkTVrUH5jj6l
J3Jcv9YMxnSSZeucErVbtgYnHy5lSWPQf0/+AmPdglX35YSpOQmB9qQ1HoiH
m3hDoDEFWFJKGJEGjbB7+ituYrURFhM+8WiBbcXwVBflnpalgXlCqzs7fktV
SlzyHB3lFVJG4109o5lrgTpwzWD91xw9h48kxg3FL60GtSkgYlsbtC/cI5I+
saWhM9caEAoEyKu30xLBmdOoWVo5tM3LhPTkEEbo+WUDckoHSBGuVTLHwKvp
P0B2ujuW9oUC4LJDYYXvKUq6aBihWZkRr+SuGYCocoA/Fw42EY/bYVstUTkv
vGSYmiuj5wYYg9DUNq194oQJrFD5yNPL92/Z/TIlFFjgUmViCD9+GLJTJoHF
9mbsPySOs71km9VKvd6ehjAvYpt65PWNZgoFQcf6G5epHIEMILKtYDoALlDa
NcT6Uz05FFD0dBW2AMegwobqXf47K6T1gFGPdmP65+XIeS2QOm7WU2SjCbQL
AxxBpeEek46gAJ+HSWUHOJM4iSqC6VDEzePViOVO3SgZxXMn8AfzWmiPQQv7
RHFlWIgR8Q3G6SdlbUVoCGhGt5Ort0G6OuvMTVAyFp3YuMFTK9G8Q5yf8DVm
MCBJli5VUXLnO0vz7orhkaTdnV3h0VEhmKFhhhdF544f0gMHjYe+QPRlQPpB
ESttcbVbpd87uD8X1qTPO/QmlEi8t10p/VoDJliGFDE2/FowlANCyMTqIIXg
3BZZCFZx4B/qkwpR5iueOgGCWnzFTB3azhDBxZj9L3VSS4s4PWaBrPiKKYya
KzwRapjAeIOjAQP1ZsUOrx6SXHegMasedUI3XxQD6OAQOrKuOKUz+OrdYdZm
sKlfdHiIB37W7zIb1saKYoQQiq7oDZItDJGvaPgPdTWLRKHqfeKVYknduCap
kxrcYD4+I/bj9+sCnedFZxcZ2e3uTEQtyjgzFKP/RsYJ2yUeDSVfXugnzeAA
SI0d7griI/9bQrwxO4oPsQ+1L4bU4gw2w884gMDu+24JnUPwEN7q70HVclTD
QYxMGnoDC98Kqi5WFNU8W6PWfVbX/BJ/Pz/fvao6rtASPie5VBJ9Cu3F6qOC
tM6c7AOcQmYr0k+Yo0RrM7tW1T/uC5x6ow1qyEBGHvB02m/D1MBYWMvICibs
ib0GbmDzFzWJ6Cw17dRG9wpgwv+8iqn9jNBSUYec8/1B49y+oQHNg020R0fE
I/nrs6CLUpTlh68HxQcP1Ptw52rzi8Ar5arZeNK7iuof7n+5Nz10e3/MLvTY
02w9if9LGd9xkwAwc9MoYdBCK6H5iFqgVnNSHbvfnaS3GHeraxdt4TyOGOvx
JdIrbVXhYT9YROfNnVi4oQN7hJTlmiU4ty37xmaoe4cbbxZnRdFLtOs8AMU/
LG762WUC/0AT8r5yyKk2A2eI7oOB1cmamuxJiY/TZphNYFgLMFZo8aC4WFOg
larlhVJ7OsW/GV7k1IQKXYbd9nHvFFLNh4BymWIl7ECGFnFKxi5o1Aveq3LA
dog7yCWSYZuMkETesRtmnajxH9F2PhnfJDOKVkHRQIl/wgWxOrnkP5scNvxf
EEcPh2OjafD/gGPTFqXI7oWpkB1vmaxGxAxFBExW6WNx3z1vX5XbUt+vnLmt
Ss1BimAbjyGhsdkvOZCllSm9TgFSoKMiEwXaTEgZpo7AjlFZOjdap1r0H+eR
Qek07nK6jiaY8tZcaPSMrXea/pSaBhB5GyMZ6z3OPfc4KDLxqS39FkUXerEX
6LhpEHyzvpZCR78alVQGDmgN6AIsKlcgF338Lr/ns6DdCcXIeY1hh7nugLDX
v2WB0HmdbZ6VdVAMKiEko+wqNdm3+mygAYVmLlZuZj+J85M6BaYBO69yjM2c
Wau9UOJqu4euyqJhg9Oa1rLMwgODLEnwr6lv+3kXaJutTKdqj8TtHYtNx9ua
LLvSjdf+SghBi0o5ebWGc7u6MGnxC/VxauLKetwrofP+5cbiJz/m8AtZKXp1
dSjDlE50QonR3g/TCXhHFamjeAGL5l8M4XzkplrkYy1rZSeQSaZqNX2DkjCv
beyh/u4g5IHf78nb17JjnqkKq6mSU473+Nf4YjNwMTfOVqq42aL9IgAMyU6F
5VntqYxtIl5V4cp4me6KtYRkedgCoomQ65tBMJj5m+HG/oo7ojFm1g1Ic/Qp
lBe9Y6TcC9HBj/aaJtOAwkIkZBowCkIgtwq/GdE7l3xGtHaThQk3dBdn0c+M
WVtx2DmTzm4yuJ2WT+/76yDODEl4aJPlorEZGnAP4GxQcGHsrEwMNUt41bxg
aVQRYM1NJv39/6t0dcEGoFlM9VkEoPMUHahvYxDd1P5fFJOUiYX3RxaJr4wY
tBxMZwOwFCJh/VLefe89crl6XgTvLVjAlIxN4b7I/UV0ebJ/j4nwSKuK7Bab
x93iKa43q/tNXPIkbc+CIHwM1qTPPkddbD9jC8kV4T+aS7viptb2ttbQejT/
G0883o8H0zrKiUNRq/9+RJfLMsLsDqiEy6maZLOzN8vdOi2R6xHX+DidG7BI
uZaMbXOES6YcTwfJ/aD12nxDeamoWmUb4Ixom9gOUdAhMkQTLXWPK+k8hpdW
EFU1t7WOd+zyNuT34A1XEix/bf8VyAcmT/ZsE3sjfsZenNeWqupgGpM3S31t
Vugq1brM2zFjgTWbOPvFUnZz1XGG+bPmpt6hYg9zY4oV5bH0qoepf3zI4bxK
IiLNumlktvy6lYYkoXnp0ka5bcgYFz3v0DlccI0lYSfv01mOLKUTzrbP3mDu
eDc6A/LnHq8488ob2P/wse+C+2DJde2wGI5zzL319+SRgCRlY8DG3pS/OGsS
XaL7i3j7Q5UdEyKWL39hvknjLW+psUrQAXe+xH4re457qXUN8N8AEveamOxt
Agg0YetYfKoGxSbHCxdzNSl9DR6IK1DQ3Bo5dqXOJVOhzQr3fed32lXPdCjl
Nw4DruSeVBr58oMkzeGQ2a1iMWJHuzSDiThM2OJYBxSX9wav8JOOigs3ywRJ
TxV6XIaMN9+bk+k72S0joAS7m2pjzWP4hUqwKluI8XaZoehTOM6V3gozidRw
9VICsAvqkAEygzk21eJV3JWyYKxWcBx1ewRO+64Gp9NtP9CPPQ0yPyqzW2mr
IKT5tppGHHYT1sruC7/1dsBzJ+2XZm9GxLdsKTZi3I9Ba3IMYki3Ie856QbF
ZPMdbqafKVxLJ1/DT6V3R9mR506NPOE+S0X9e+QtDYj+zEBdJDvCRiOfJCsV
sz+uMuZuxUvOi2wpnkfy1Ky6hyxRAeo5N/ZQ8V0RoFvdLhIN4xycYfV4Evoz
S8mG+0wb3sy8UmeVW+zz/q1i1mqXNM8HoEEkjLoBj9k+k7g5GDpM6/Wj5MUt
4i+F7MwbnZ36ASLrolHfzyU6602RYKDiFOwBHw7z81fvnQerP0NlqvKXZiwy
+FLzSidDruNhRnOlIsm7KKwWlGsFw/75A/w6wdnPB+4QUM/OXUilqZ5xFv/d
F64dhpd1HNfsKvq/Mx9VMciavPuBT8Bg+tGnMFgV6kIA7hnYuzXyRq/n/mCp
y0vhWKCuN4g6X42NVq/PUdPtlfpOe7liYXX8REJ1/1cBtDnfb+lhN69aJZVO
E6580tU+v3uhj/O/Xd//YKhNCFgAz3g6V2MWSutO2pymMbqqGNfkGMKl/8Kf
w/ndFpwh7I2Hcg2gWNNL2qd2FUtp3QerYozArt7xLTr0luHPnzO56q7hOT4D
A6QFOs1Gl252lVPgVSw8htWAt3DunK8UBLgyZ2hqBO5N+HP0l3/Df+aSnlW5
1z0b9qeI3rZtR5d96GPxXghL5CB+aJuj3oFCIUDCrBLbEdrZFvpH9RIgMqTm
lWpyESqazlsiJsAT5Eta80YqVDlhZAuc/KXSsj5DXTrXBDvPZG63zGsV4XY4
A7Azy9NtQroc+2jHBm5XtIzrJbalZrGSOF29eGwdJkp1HSyKOS5wG488unBG
To4oWlp/0oLsws18DLxPFagGVNhlgl1fNLzdl1bCQDep80QdzqzkgMUgrenl
f42b1MWgQCJmuS9F1U7P4fpqPmEv/8iKRTj1TeZ98/7Cel9Z2xVtLt9cXtwT
oRxktlYb5iwMlKTnNTKj6EicJF2J68IxijLihz5CN6bXWHp4F5d05bdXmS0O
y2abvUtOoA0QfuqT79uKp/psYJn3gkzTSEVxUmEUz0MbS/h14C5gVyuFwZDw
Ea5w0sI8yyR8JMOAXq5rrSPBK+D6HSMYArFnWvvpUp0JlEI3yJeATqHsCyNf
vsHju63LIzTUJngq3lJXQqxuzhXZS6SC4iGmkKDubHhNNgcuSm2lE9fL/uys
pT5Y9k2Cvb0VNcB6FjN6YjnUiWGsZvr97tOPto9BKDw4qEy24nGxnTxiYnys
2nOE1N46lu5rl94x9kutVkAVK3cJnanIEUJmz1hIaZRXuB2L3jftr2yR9XmI
l2fv+to6MPPGW6KBVT+LtOGS7/Tsh5oFmzV/KucsJofyP+aY0ayxtsAg7+oq
j8EIz4u3d/WFYDdNzdYxPyfH9aXidnvCcKrrZgRFVCzbmzu+vgIwNTEe/ovs
sk5xwvKvF9tQ5KzMA0twiNFlZ4yiyVZlA/08E6Hu/NRPy42e5YfAM8QleAMt
Z6HY5nJLvQZojFP+EaL+iNse9kjo1xzCoEKag2LuFIHYTnUm0FQlAJo3pqjv
ICopue4/ODFOiOFlW2VtKGKfyErsZZISVbE2IuY6KRrKwfJs4/sg+SDkyBfk
8Fg5vsZsG8dZA3H3wMpeWwUDJSJ28jF+xtJFIqrAGTm6lz7KlCQC9vIXwJPc
2Jc1Gl2V2IOwM51NxJpsLXalZSrInuSnlnfx2yo3s0T9Q/gHAqRrJzF9naJQ
P3gjUQO0VXcGUkBHxaWUOJA044wiJy4YcLwYT6MgDNErJy/bbK6mKI6djCk1
HwDCEJbxNTNlWifMkDrljrXEknscTeGgQR4NXd+/4bfss3Myx0gAKKWbpbf+
laudq7Ph9zGuczoVqXW2YTjGkP9+8r/b86xVZ4mC9THJ5uoJAcmZE2SwTDo6
n/jc0gf2CXlnDaQ4nukvJ2bR4zMmJZV1w6SSCrYQJC+IC4s0I77FB6KVacHh
BDifZY8vuSz3fmPRkQYOKGn6VlPms89TzgUfFLKMl0PTtJgt8YsBCZ1iUlV+
r2EwmqZzEPnVpb6f3uckqm5PYmoiVwuZmSmZ+YHbdyt3fVmuCdOUnO4OxHb6
NybGgJJaWq8IE43veQ2VzclaNOJtEZXT/yuuTd5ClBKDBpQeSBpJ8glBEr+i
6rurCUZUNEoiEg/HV0bvZ3gUSS/PX6QBL8fKoNiOb6nuDjdau8uUlm1mi5jS
o/dcUV8IipyBR31T9LktoUEWXS+yAmzEb6dQW/WuTnPF8EuD3DwDlYTuYxBE
zJ4jGs8wyqqZL1w72KUr7hAYA+S9G8eA/9eflBt7c4/biGmQ9gnsxV8glLQI
+56jBRqBDUqA8+P9xmD78USwmmc4JeOe4SjDadbLz/ovGrMIgqblmzYrHUt6
eYZNgQE76VKAFSVvHkyeH8cL86l/eJdfib19a09qINlYs6BRBkiIOMTbLaOS
B4JwYefL1iiVTE+G8bR03Z98CPBPWpN/NqBAvDnMObpTFr+hxOrR+XSKwvuz
rgfEEIqiwP2BD33SQywOkslW3Kw65cw+sPrpztMws+vAIQ2TU+GOzTYxKu/h
Fv4zl5sb/pWbtLhHgJA7VEStE0BrluHwvH2TRiy5Xq0cskcLOcyr0RQV5UWV
N78cKpObPntTr83F2lypvYsz7lEKYS4zKqlWy6ZOj2qUGibJNiYLkqFsfbaY
seLza3MoY7GAHKmyY9N+rWu55BZlrTxVO6MN0PJMX4XTowaaFVQTzksbbaaG
5hYagYfMUjWidLqfKB3l3JrxSxFh+mZcybfd1DyfrLoWIZs11nJpzkEdlzXQ
SEdgRo48auiKK4S/hZndYtKS7k2p46RTkPxw6fYv26GV80sph+PHkO6ORiD6
Xt04nPiybWX88Ad0asZXZznjZBCylGYCDppynu/2mWtqok2JFYo9qkRKVVeX
IZvmZoQIjqC+LqPdCKZqL5TVh28T0dz7bXEydezaOBDKjMrmldyOV+vxvPb9
id8AXJn1KqpaZx/qfR2fgh9UQYy0RFGIXF7oVi3AxnM234Wr35RkDRKB5Mj3
Jfk/8SGwytYfKZbB2TwzNqyS3ypGZdXFVoS5ETwWYHU1j9EZmyoxfeA2yDOR
KBZ1YHqXn8RAV5bGxQgc4VUhdEqZF/aLdPE0++mAfXCUlNzvGqY/M47GFNwd
NGdb13L2iLnUnkqUNUzXLzDqrr6ggkOXsQIfYnb5+yqKie6H+KxPtk982Z/4
ukLTi20hdTgzdtQRJH9lP1P9Xlqdrv+23tPUDXWYmsTacYpGahg2dhyz+Z78
0w2hgOG40ZaCr5rGjRzYs8G4HSHmqJuXJKf+TBerXesT/2JDr+uDlAE0dOqn
xiosOCIe/PGnlfxEOsFKt2WkGzvrgZ8lB6CDqf2ptACJZPhxwip381RZK6UX
wZh2Kykv1AgjQ3VghoL9dEvvpBgG2Qyt/fxi++zfStXYLZya7AHIt0s9G2XX
7ubMoFSYzL4blitpaXZKoJgfnFXPBO5i9lV/5R+km2UCkAH1WZEkDim4c1pq
E486kLcVoW+nv25uAVdLg9qGbrRwdUABhH3p2fx/2ePFDr87tPsS1+Oq7cFh
dAauyCEUHuYdEaz8w9fSHlXwd6ffCKLyVHUqFaMYz9b02Yc7Gk+MQk7Hlonr
rzVVoWa5FtAX2gJR0unfLL7O2L01toh9Ds+deCZ6izRfRlnCAeKkfWGqIUdx
z8U2usAMHsvLAqsKhOd3sgLloD+b2s506d63qhL+03XKVCZngE+HYEzSWOFt
DsQT6hrRzoZxyQql9Mcak6yYoaHi0vDvMvWthF0yMPvTgAHkHNzITI0BavCO
u1e2Wir+G470HRInu3pQyNxna94Knd2ZOjtehUOgXg+6g67OFKg7Bun6tzyX
dktNENCvw4sf6VCEZfJGTeOOmW72/8JZ6O8vyUU+kTHy66QQlGsShXs+061D
bMTnanRN2OQSxJDGV9DoktogMoAP0S7NC6TBZSwX7pOFBaz+YxgHQgK2IzUz
lCOL+Yi7zynZmXG024ewn9pQtZzPcxN7JSmd5qxTauIsu7tS/XscCCbuqdBa
I5MohjisXU4DMttoq8zs+Uy5+opr6rqLOmI+9cNO/evOVhZ+jDbfI9EFHQCi
RXV/zN4lECNhnA4Yy6ysUVado+QfnQTZJTiJtIv4fDQz+MkwQvvhIxM6mjMj
RO9LOtAtWv+b+FBDd32N6ZJ8tSFoA1MPl1Wsv5OlpKJRh/1jrM8IQaO7TxzM
t0mtlD/DOM51I5jHQEE9MSvPfahay2x39u8aWVGgTmh7wVhnyYxB5xBUONR/
hxCEC4a4IN6iyCwB506cB8N2+ud95CRtxJKRkylxkW2lDdI2tN8jgxKV3h6Y
5i8P5GoopFGOuP+0NjGIrzBAXWpqdcAqlc4+gHX0Uo5qFwl2/2Sbq+dJDUrP
nedCEr0+nQGLmeO0UrbHVwUTgmW8vWGzo1DFuQdMU2x8DMlHXX6QxuSepAF4
1yJX/8teR+/RxdeBtaC5eRBg+/FsdpYBN0RFqpUBnAJ7cNfkXS6OKtOnZal0
wDAKWjmLPSWW0mAmpls4zILBJs5l3buxhwfxGfVWgGbKoyr3hoXxpwLbOw+O
oy9JPgTY4YPLxiRJqQPaqujLoz1KFh7wuUgPiNPjGOVzHey7mbT7z+J4tR64
afzKjyLM9EUV36ztKzVhEx6eJ60G8yawRluP1MHujRYlRzs3g0kMc55xR5+u
klPkE3lwR6SX24MEcHXr1IL3pjArTQKvx8QgrPWYiTU5A7W+vsVVDCxX8vC3
4iO8qH9yYWlytuDMh3tWN/2vc5QcilfH3b/aT9Ed5kYQLTdu/QdTm/tawHNm
8qGTqKkyy3DSf6yo2efv3vjbyrcGIVJRSSVfLwKRrjdvHJxkFIsYBOQvA0Wa
T5eI+I0uW0qVla3KrRH6t7S6fGF3Yj0UUF49ac04ybLvg7k7uIf5VJYcUXhE
wyralsW1tz0NArtc/xGDdToShJsRhzTV/hF1onkpgl7VetOVln7Mk2A0Bp52
eh4BQ1Z29rS6sr5jNYR7HF+GQEUyzP2OLMQs4j76ONhI1e3MVJysrzZkdc5F
7IC/8NjDRNZqMeSutOxZJsoXH4Qzwwfev3m1JTjkZmrkVHd/Fwu6j6ruAQmZ
LzvD/LalmXuIEn96Qc14jPnuE9+badmXwWNi0ebaQxiuRm7kjJM2ryirAuEr
pJlZVSCHoMinABFPJq8tI1M6AdvmYXE+XTtmUTSj3knDSbOVwJMkS2O8aPQF
1siVbU78RxKYKBgphuKMQiyoRBXHO33ggO4iCcGtW2RUi65K1p7JNUIyogXK
Ydmu2v+lM6G+Wi4tsru3mNYmVhd8pnO/77tVJu2DZdn1tIICRt6twpW/ac1D
D5sTPcCb7VFfThBamLDocietSr9dsrD9yVmeeAmaVVQFFa/MD5wimLLLVSpM
roy6zFew/wb3LH3p7siJIp7zuc8D+cy8+raJ1I6x1u+2ozfglLbc4bLTMA8j
KBuSypM9b+3h63w/5nb/smbTgIeZfz1UqY7hLL8KCnar40USMaAboCiPoJjL
+/8oabLfrZyLOwrmBzddVrPPs+cOUarvTEkFIaPihI6To9QNPXZa+dsXLJvS
clOL/05uYkGBLKuPc/G9Z32MAO86EIRyw5xQbirfKjtz3Hz097fPTx70stDM
AyKh+ATS1fF7ILmb022Xl0FdROPpA+0yrX1Qzj03sHVAeUcTJWbesiDwjJ04
kBVWigQrEy9nLUeU0pHtDHndXewNI2C1uISX0G903DX4Qomw5ykENIIhhwO/
q3IIqXz9dqjSztG0KaJfBoDAZRSM8/U2QliRWTntSPSB2IOjWUVSujQ7A2p2
+2M+VWOVieiY4r5mK3YoTE4d2qUn67SqB9pUaFwfWbPgEgfhlsnO7vQZGT7n
ng244F++0Ws7WrsCZA9yzj/TYRTK9OC9VnL/EiP3va3gC8s5bsJtJVJ2YZDF
U2YAldjTywvYLdJWlkPllUdR5Kgd2tkyxnYXBmVNkTUByv/EYQE5qjs8sYqB
hwi/qQ7EJMoGobxc6g17VUHdcoNEXw2RsgcwJxl5Eph8TKHA6B9JFL4IBL33
rB9WM2inr/MAXX55EFz4HW3iyBu001coa1KCVu200BVqdDLUBrkHKDAr4xsX
nVODaLMqwn2rB186oxEg1SFX8YrUjw/y1KrR0vRfm1mg3ePeVgcz094VK2mh
Cbng7d68OzDp6m8cvwTowOEvLIIjICv22/DdUTxWmxhFMXzYwaLEQi0u9SDT
hev9oAl5XC5NES/KFDbGC8FLLKdckSCnbBfqHKmM+yh+L+CJTY+T499WYTcB
8AHPSOPAKy88oQhJIhPIhpQSCsK+e9Rf8TFusnY/CR6BATcDybpIic2xHPZq
RJdQYEcMescacX8Q13cQKuAc2DTw6SXpysez6rf1GAWzwQTMCyeUVRcgyhbG
aNCFObYfXPSJBOl/kkEeZWKhMER6eNAzWTuVVAKC6oHHaMiSazmdI2yHhJZM
2/+TKug8R/npAf71ftQtHb0La9JTnO39Hb0GZB4HQKTNM31+NlMD1wQTL17/
Av4M+Q8UqdTrm9b65XqUrtqIuTQX5PwXcxO1+cXo5EAQRiqOnL4mdj4C/LNA
KBZjjHdfxXXJOEmtRu2YpHhzj2zJJRKKmCc1qgHbAJE7AqmYZzbgfdq67zRw
BwDc0iTzjFrU6+usxUw5o9ct8qFk70VHc3yjv/9Zw53dmR9N7xGcqBhH4OS4
sF1jZo0LTuU+HSqIJJymBGXW/IvB+o/6NCvonq48znrjTZmzkPOwVLYzRzXW
mrYT9cYVRxLh0PIwWPqQf7aivS/IKRFJg6kEyv+veaxirus55tJWEIEPO5rB
La2ehOzxQ5/OTAiaUvqptvW7sRtenRARRSQAZwOfHiJS5CED+rbQcoWEb8cv
j1loKiQaRODoQDsIfewVU+chx7AIW28Av29yIL9tjQc6/0FR1+Pfj68/a1vx
6qX0RP/M8JtPIVXQ6C8Y+ukrTH3edQapvUX071z0Sm07nrPTnceRNG0q7Y74
BC7QWlw26kYQNpsb2exRiqd4WACKYpnVNQ82xfDdwXb+t3zciK6lOi1dBvc1
7sa4dXvNaRpXH8FO6Eu6Ql5TuNo96z8CclMSlCkhiB16liiW+uDWl1SVjuNu
tYTlfrYmU1JyZAmZp9yEVp2Rkn/9EVImo1+S4QDlCbYihLMxK0Vm4kV0xPQ3
BAOriptEV3hTscYAckUOSA/+89ZgIcStK0gnSdze9H1ZYGyE29XessA+SJyE
aEVGRgBlYgYYiYEHsY9axT3JPVXRUkWFfx3xArVQ2Yre5RAffzSRvYnZx36J
g6Rmg+G+IQeNN2XMOZM6iAJNM0K1b1N/94q6R0B0wORLk8Y42+kz3vWMbvUu
hwwai7stxQV1l7c2VzqeSGuajysZBT2lfftlIqy/+mXDxvguubU6liMpxSN2
AYG0cs1zpMf+psmwzDhDn4vAFfUoY1PeTid00mOhdDXsFYW1yw9/kbtMjidb
ttUxvTb3LOcLG5Jz7Ezh6UQRkccFsgdrY/wtv5baEvVL1Q96ajAPAMFr3iJu
zPmVa30IBXjlwNUSDfs059mhW1Hw826Bo7s17dTYeBydxr0S3CEgf/tjRrKt
jdWOqG8YLu3BbpfmbaREHFSgj4Fk0kBPzGoY91wuk/TGadjdFTXqOgtlK0Q7
d91vJOILLgHda17pV041puQA2EtJlZmSP/jbhNGU7C1HX4OvRs0fRIEywTD7
Lfd91USlXWoRXCZZ48Eu7mc0cKXwvzEKLHNuq2xs/Fzeia+VglFHUwzUap2G
y+LS+4g7uE4e5ohBg+8SHrzqv/GCOzo5tl1/J0TvZvSr8ugRM8wSnFCxYCs+
ieqMpDxiXQ75rH2CScBKkyb8jeIFXs+ilTUx+KnosbMckuIuGuMk+eLSwvuE
Qg5Ssok5VrBlYWS0mpM0yPQ21NpEnluoZYcHxzkQUyOBHM4Crh1B9y+VgZUu
GuBq0m4e9bY1xZqMeUOiqR37ZTZALLdpuB3MReoGsO3Cyc/TFnciK0MtQrsF
pvBQVuaPsj4ka6r/0f7LMVoMF+5JhkciugiGUo6nASKtpkDu4cXw9JBGdYNB
t9cnBvNlmywWgnO8jQooysfpf3VjL2svIsuyENXWcNiQBRVmn31VntPz6fa9
O8Pc0AFP/FauyiPsFHPFuTUveJjMbnG4Op/7lApYXRz2mODg7Sst8ldRxK6p
7V2+IYxt/c9wYDlPmFK1pWF6d8Ztudk/GxahyLfH8nz7V5TmbUIRS+EhTNhS
sxPj2P5xEORqKxMWfpEYjgnQgn+U4RCdVseAoB5L+LjB2wO0xxoqTlU2deJR
h3FSaAkt16ogLZOTU+vg9h6+u/dPGQnB//8qy4oM9purvhyuRZNlS25Y2jEv
N9Ur1Mx6Jy1xWuKz9Kz0nkfjBGr0lyX5npn+M+5ErgXfB+ZuyXFlD55JpsJ3
Mhwwe4Aklp9I94W4qsJnvkHfBPV2QpVvn1N8ZnasR5jT/hu0BjiRPMG0jEhp
MeY//DSxDyodj0DgZle/WPwwQOGwy9BCYlShIWSjl9HhgkM825ejKMXr6Cqa
rKsm6kAkyscPKA379WtYhurguf7C4NSA34Bj6DYj8LMO89d7/+76Y13+rocJ
hCGHKT1rEGg0O7wVJBJCHSCuAAEGf9gs4AGPgaYR9Tt8m69OwY0Qf3BoKaJP
uUnz/cavjXfw1t5h/xK0q0zhW/RZKBUmkLO4ZNKR9d4sQeVP3izPzOEvcwiS
Mao2NtuMCapQ8/w2TojeSBQh9hDtkQfEUeMvDyj7kaCnkcJOoudW04ebQdHJ
ONBLP5a/POrtOTV6AoI6sEyUcOHLpRXhQv5wglo73V4VLfjSg2lC4LIfWy2w
Ug+PVCB/LeCJzkxs73wVHyNFwdnYBbDnh1PAOpWXXfbzf+ltJ1IoQsTMIlBi
tLl8vQgP8N/5/kFz2OrShdsljRoTX36stfHqrYp/qGykOd+oYvETKB5sTiAN
4LFNcfB5+xoi1wdaEuka3p0RAFTIHi3+MbFSTrB9Jp3JR3gDOvOdlEXnew89
coSmOoVtTUI6dCvYD60DyHOHWaT0t5xTeDLhK0HgRBtsC/O7IjWzxYp0SdQE
ONkOJTdJvMHeIoARdXcVMpUiPUR6r6YesOSBp8agCy8+EZsL9uIGLF22SHu7
FKiXlVdjei7c8NV40v6N0lHGw7f9pP9GV15aCqDr63dpIlXzOcz6QfpkLf4V
HJccGVkPPHPhWIET0KcAHoJ5uRwEbhTk0FkonfdYpPTv8bLsR7riO2YXbF1j
eLiHBN2ETA0n/VrCKkh/BN/IU60TERyOpTNgbXXbF1OcfWKpFTc3EZIMwBor
3MQ7J6eRpUQpRkPKRrsEskrexCcmxfRFRk9lArpqWGHEzXXbl/6usBZu18EE
FLJpW3UK+YNeJc14MW5L6vFbIPUPw1yM+pnEpSlbOt/FqqCjyA2+ZpinFKFv
oXk4C5ngEcdUzKv2rsye4uUfPaOz/JXlGLH60jQg7LGgkiDMScH4AdAPHCRr
sH75b08oPkDxqxiqzIs52O5AMxbDAGJMtWbOcciDuZVUU+LH8JWl3Y3ADF28
tEPf0mWC/f8GJFjkLMWiQiCrUplAPsH+FKkyYFU3BAn/ickQXIk+79mfNRcH
harzszncJDdKU41+MXvoFGgt4aI5M0yHQ/UMrDGov6WJtSMBOU+ffuwG2uEs
ydokvKvzo4366oUEcuLCS6w+i2+w7yYdGfY+X2N/EjxX+Jvd58Jl1djCbttu
c1stifhUl3B5y406tuggbNzjdRYOTX7789Yr9zRSQ+tIGtAu/LVNjATIO8oZ
n4qCPH3Qvk5vXlOSzr4l7Lxrh/ZGWTVHD0yVDcnzSL0HC7KfqgZCNJ5FlnPr
SxkdYSJBsdYsLoe9AJ88rkZWNZcQeYBcFQ5Yi//58U5+DgsGkXDiwr2H4G3c
YQu/70rc8+xj7UL3nZ+jEPJy3CYJPpzPxq8ngPsoSSJj0uYkw4+WhaKgFSkZ
XpWqHYM/NzECsdt7DcHQI3F+fsBuLOwRqFeE9Eshb0LXnbrj1PujX65Tx6MI
SnJACfved0SaSbwMhZ1Z41P7pZBdtuKC0P40EYGK73llNKXotgJI5AtH0Fxa
xcjOW8Pd13WCYEt1MKkoIfIxxHPVufK9fxNRcJbpgC+8Yg5UJ2nSXts0HatQ
4yz/zO7MX4koO2wKCXCTLUS/eAunQ/8KTnRk41CEY7ThSsrnlKiFCNbC3R6H
KeQyH+QpNns1sP3UEErtVuq8vp6aYG4xb/B9hzKREPwlhF9m4DccW19lTByE
S3Fz4YRnC904FQON+0jKvx4SAP9TFmdkj5WX0FOAVTpTxrPgJkjoIFqg3tx9
qxHdANaxUu5RZvkW30VVbX5tVy+im2r0tdunjCxuebciTHvLlTu7WcvXIJbJ
v7fPaQfLh6jKGgTH5nDvsU3UJo/umj7xhejJgchbJAg5D8RGbn6WPOkIO4Xc
LJZydCWPVj5RmwubsMZ2EUGTCeUAy4rDN2kGE5dtXuSg/M/+JsRkkoeTznti
NAviEjOyVQDg+K3ZZ+UN0BXJhn0fI7osrkp6+WmxFQZ7RvF1xWMkoZCCqPQZ
5uXwowtXscBrGdQ9v98a4cbRggSDiaEK55aZSf9bHeyslUD5BgVzDGZ4h+/y
xo5euj4MEhZ63Y0tUeljQDxgIkFgUVjctPBu4v3kbvmYPFX1WfTNzPiRu8Pj
x0gf2EtLSz3gO0xgqmInH9RvB0d2C9ypHJNe/f7PuE3KMrh2skSLCq5+luRy
TufeX61egOoY8iZh2AyRv/rrprVv+qhXlhdzWSxdfzMP7MpEh1oegS5UuFpI
9TR5ybmAheXisWhXUyAJNf4/EU84Bw34V7rW/AlFeOK9OA5z9gaiqQo+rIT+
SXLut3/1+aioIyzTHjcRoUdXeJMEjq5hvqDRBzeXS9mOjD9/2h4qpAE1UNhw
z1Q/oD4RbAV9HMpdZaUowCnHwh3hpfAfprUonIE43X/NbvPwAHDLzQ010e65
Nn2ELGguhPvtqkUeQ11k3x1eOT+omFXONIcUQlqfJkB/kdPH9ZDfx4MnrgLh
R4EsTLXLdFQOKlfDy/jBbFtlwX5wn5OepkMkMxW3K/WC0LYVia2e2guw3LUx
fFxMsSCVcTqFVNnXN4fb5qXgtJGw7Tp9T4qIK8wHv+aBZLz8vXwbvFHZGBgw
NzV2n3X0CL9sbJckEGgxqtpaH0nCiXjhG21l5ijOwX2pqCOhWMl7qK0SFm8j
tckJOD4NElGkBerjG3biugJCJrIOwPaK1OggsJhyFoKgDmuT+ldXsfGmMLSr
Jy1mOVQgDmtJgJ3COxxhyvw1yxOwj22jvG+qzQtoEP3ZBSnBCQ77M1O+DlWu
HIsNPPK8Awl9nW7MiFl/sBcG2AsAD0RS6wobIOby51kIjdoNnTev8o5X2SOf
0dVz6INZ9AU6txWF87viQMvmxMTdm17qn634NbiRgVAv0DYCMmc3iA/MKAMd
wNe1O3kWTr7MoYbusLIdNG8jhhSck0hRMy8xYjcL1a/pE4Y/LaNE+o26J7UP
qXjIxU5hHYA7PxFAsKi6nyIx5qSuFdox3kDCxfHT3xXsJz4DklzIEze3Wdf7
2BSKCO95IjuUL/9hENVrlwq5qb/fsMNqgf1umu8Do5PAp1tocQW+MyY42q/0
v5g0RAzHFFu92TrudIlmQeaUmy7p/B/FpUkYEVwzpJybfVTQro3IuSlLaVtf
gIUugOpEF6Kot0T0yK2UJn9GHQJ/A7veGWx/JMuGe1SwD6DEsl/+w3ZXvD3Y
/Rsm1gbaxx4Wy59Kwg93KvJ+pYRwYQiDP5j7On+T633GoE2NGGm3xwBr7lws
mUCaIl/m1T08LH+nOMvNOOoyqZ0PUhJGNiX1OyQR5xrQuQlnha2+fbbX5ao0
lWlTZTa5pKOI9D+iV6Js2/+M7YUOH7wWKXkQPpSM/rEePrt2yvJJxFP022ap
sbXe22c+trkW5KAcJscIOCws1jLso/RnqVWXrHFhDT3KIifR2mnVD7EpPUT0
pRtvKQyYZrflbgAEZ0y8/qMpXg3vY/AIDvUS2sb2ipHd1/tCh5RSdNBqbtMd
eoy3lnDarn1nnTWZ5ELbSv8K9pMLEcoHev03qJp3fxV8TUM5z2G/bmNS2tBi
8p258vWjVwcFp1xBKFJdfyqUwnkthlWTZn2yVw7m5JlUuhdi6XURN0tQlPyn
ktTkqAOU0ies+7C/3ApsrJy/xg5Zc53RTX/gL4JaUxgQRUEJM+IFm55bFS4U
a1Khxn++6WAsQGsAyoEsYaCSPxt4u0qvKZE93CMiW+ar8R2iwyIhlyMRL//k
E632dnvXe/YN+HHIHV3E0nxfmO+cmgm7j0vbcJ+S7EhcscA+afmyGthi0Uqj
+ip1qw9utQTkVfxDvlv8mPi363Rz/rD2ZbN+loSTSN5oPaiqhuvrkAkZYuaX
gu/nIRclqDQEUL0pZtDZPpQnmXDf0V6s92sCMQM0xEF0NAUrluLQO9mWwSnL
8o11odhI/4+C+9KEgSonVBUK/aDYjoSBwWQ0k9oICnbyIrcEK3Nw02o/h1Dc
7ikTQW0ykPCOMaWdef2TyWpbUIEqVsBBycfAPJtSp8bIcBjoWJM0t9JU0Ufn
6H32zWx+QKhYKH3bkzJfGvIcSWu6oUUnmhJ+EVzG99jfQaxLcaG5xzsz3R99
x16bhttdgIq+rLHmczf2+eEjXYPOtnZQKpJOMwKdJP7f6axl62VGfjEiogng
mH9bhoBY3ePBXm0SF2niXbOwYKy+0UcdB4qm2FfL1Ao25KPGpT61SilHfHcz
UuJojGenXdgwHGIk1ULSHtRjcowKkPvG834WU/Ap2jUa52O4KON16PLG6ur1
WBqu0PPGdgVel0Qr4uR10quqJ72LMfFarze6gMXs6VH+nf01eFsflRYfnyoC
1ZvScNmSjENzgAX0EI6c1lC0Ber6ERetIm9Sj9qP3mQEsI8MI3qYNmlFOq/R
Nl/I6IHsCWOA2HHa7hTxqqQHvEluP6EqTVCe7kKBx9oShUFjMawXh/C+HhYS
S7kqF2lFCN+AMnxnenmP88VL9vN7iDUiNw8CfvntZbtvHrGyWE3lOMYWSLlr
qDwJamuSiZcgbLdOggVIYR3YSD3O3E8JeBdgpKSz2inT0fz3HqxIdhbK8SU5
xev8P9sBSiipXjex9jQUSbOJ95RCqv8QKAdPsVdoGwW6hQlsnZhD7OuCPLK2
hWz4t4m0jSMBmbsLbE0kLxguGcl86KZAEsYFJuVOx0/0j1pbaP3/peAPUZW4
vKuS+BJhou/ic52w8JRehsxEz/nohwxVMomDfa8KXq5HL4GB3zff6r/H44PX
F6EuYV0zLlSerVshwNXIND7trDT2IXjBF8EcZ01rWndRgJMhgZeKImWg6gVg
knUC5gG22U12zUQvywrIy8cCNLLt1+op5XvlNczIrjLARKyKk3ELrtDz4kk2
7+vS6eIH70hvvzvZQZMNjkurdq95/ySGCSlHtRt9nnUpIgrUiOJXEm+bWkCh
drniidwj0sqNMjlK+mc3jcW1Blhe/uIN9DNMcjhqrWZ3y5iEPDdlH1ROFnFD
JT8d120g2zDkPnzsf7VX1BlGSe06hGhStUix96lwR3q2YMfaxXTIwf0TyoA3
9WypMnknxP083X46H9JvAbZgaMzH9OcSJVsVPC+5CYotSn4tbTh5Rb3WVDit
j3l80WP1eJGTi7W25BKmv+dVQ4LqPPPlPe7vtx5W5OeSE0CTPIWNjPTkjffk
aBRU7jxbjVKDdLeXzZ3eLIkTaLdnJnL4T7GCSZgn5L0I4zuluB2xOo2b9IVs
GnLnJVDXrXTDN2VdVZOiwbYF0hpJUMJToYvTILuqddGJg1QSiD0zqUD8EGVc
m2Wam/QiDFIK2qPlHKGYm/kOEdF6FVm7sFSmQKkVNDRlZDUdkrgNudc+jiM/
L9cxrIE0LnArLZU2EgGwmI00C5f8t0Uf25KOTpfbSjBD0qaVPLFaifRP3RTl
/D+BS7rEaeQ0xJa+k9jd89JtRC0yrtH/MPMRuU7IkbKABVdpPmKIFJjH4n/n
ZE7CxB3FZ8FDvgeNAXUl6Mkev+eOsdjFyh3iaKsVlPGZqLM6f+GzGlxi+0BU
E20RKBOezQ7bf3Y1nA1Lar/B1uUA3GMB155V7gThM3ZLqfdGKFs7Dj+KVeUa
d28r/ifS9Cy5+30bBhn4fXUqIuWeMLISpQzjHq9BYet8BMuOQoYRWv3Rj361
2QhloJicZ2cq7j8pg6reAao2Lj2z+lbmn8oY17LIZdou4D0NIjvCpXOszVzl
DOVM77OfN0BSnQYDZBXDoOy6svJxmFqk6snvov1Jj8PvW89pS4/6KarJx4CO
hhbUrJzkQ5/2Jj+cD6ChLBVP+jpZKfbOxldj7KzUMlB9aZXk1XPfZwUpQmrS
wfaYZoP66FE5fVkrOAnazS83hnR1RgyNSLvA+JvZfWEiSYcM0jhm8GCNsgq2
SdpRDqPULtTwskCWF+G8NMHVImzmt7tY4zCDP3kyKGqTDolYp1xrkUCJeIUY
ob7TERNchZ/AC3OGXR27gHAdMWguDTFoVSrQ+NvcgIrWqxwIljWCD0tz3pWc
9avXKn7P3cqRcuhmuuTks1D1MicArkBmhCVtXpbYyRnDd03MIXgIKXHwsXWg
OLqqFZ13pnF0M4VaR+7noK4kyDmHjxqYPs5rE5mKtiqcjnbol0jVsomQrbnS
hSd13x7jiF5UukeqKBfXmBEO6NUaFKUvR0XLiuB0fPyiknMKN7acspYP9oiM
pGhBrzlnDaTuoGWfUr4ojWYWGgM8dQhTo5hq7EIDAL4BSi61/G//SiOAMgaP
ui+2TvmwFoyMojUAaBa0NAKpnrnia46xGDGOc7WcZ5cm1pVPn/OQtUYL58F7
X8fn7aVGoNcNmwfvOvvASDniz5aENC4ZpShpU7rAx/W5UPnKqUSaffY2U9RB
ZoCD78J3Y1pXfnd+ECHRi53cRYJjbizUDBeZJ316P2VB2aUQcvFg9J0fqNtm
NccILWUrozTfCN7yy+N741SbVkWuerICQcbQk/JOzFQ+oAzUo/BpPvbumP5I
NH3mgJ1efP3n/+W/r/GyorOkt1VZN65gJCe4+37M64ogYV0r/HkFCiWXSdmK
PyRGE0mPC0M4GpHdnt2THqtRkoSHeU07fzKD8suhoq9a7UlP+KybTTlBzENv
lXv7Y6Lc8SjcbPDZ7xWhx0tIHL+PiD7K/F7+/YevhjMofz4+2Lue4eutdzvj
IgQpGm69ltAmb5XNvIV7nwP/SgLY1uYMbrlK+VfVSuanDA0G9H8Jxjbahcc3
dbWeHDnnbalpFXj+3x8j4HbWMz7ApmZThPKMfGkyrkbSJArMrHriIHfI72eP
XKDH2hh2hGRJo7H5dnsk+ri8moG4ZxDyV8trjg0P8HLoVyMA3AABHxlJLFH1
5zkCbLgs3lTFMnigXRVXCl3mAbwKPTOz8/hPKaO0wwpHnl5JYD2rLtLNIOn9
ePyA5dSw2mj5EaDgSdTgRwz2BkKXsSPP/P/+YAZrd/pzwyWMzdviDvdaiOnz
m7wTFpBdrodh7ubZgawnfczncZ46OESyr7prhO8UbaKihREsN+o97IiNcrv4
1m8Xh8Jm/eBToNlmP0I+W4YLDQ/ntA1twjQJVK8WaRy2qZQOn+9TxfB3xl4V
H4ByTkEeAPqeBaId+M7TjymbQXBrnm7U4gcIb0ZT6PWm680S3Xv9Xf3kB/n4
8fbcpCzAY+kwEmbzTxIpsgX++wy40hxsGA06Nh6jh1F1nHJfE+DI3TSSWi01
3ryrQIBEiXFBK86MLswaqewGSxs6uKpslu35wUJ38iGkbsMhkaUHlBd8Slid
kDiVv4RvpGc7CdfbdvlRzJAsOphjbNg+Z9yT8BW8qu68VcdzMP7DyUUn52cy
QKibVNc0cxJsr2My6qjZdNPIM8p4GZ3A3DR2pfMvnJB8ZOpCaqNVwo8Dkjia
NG/vCK6tYS/FlIuZJ4Je6ZZF3XCkRXy4YMkqR+eR85sXD/xo7LEvc4EnktAA
DXn351ey9Wtfs/001zSlT7LBVN5v17ZDBUcDDwySnqiiFWTDnMmFlyCKFfCz
AEXB9hWDNCtCsiw4TowKCvQ6+YF9FWTST3/EznTgAo/l33Vs8zqs8F5S2P4D
BKtu1zb5A88qfABs+4s3bsERm8pR2oiFaFjhm4MFcywnq1wFvmABSTfZ7K/n
wdyk5cgJQ1P32fsgPDnkhyWusgOGzvLcpacWcjFLL41oFIsnZ7wCQMO1o8wZ
uWvKfjoUl7XL24AwKrApTtVhH9E0WM893V2IfLiJD6OUwN5lO2uWcYft7PRH
ga6NRiQywGqcfBbGL0VllRj3CvORZg3WVvnBLZ3M2304+PkiPtpv+BIFoM61
/oN1VlMrIm4r34jY73joB+9SoIr9ShPVhLSCn+Mb64RccwKpxBg5thQPuCj2
XfkIaON49oQyy64/hLOsIUXVe5pRoOtfm6lz+ODXjQ6kZbn63Q7lPMIWVPsO
tRv0RsDK2q4mlWGK7ItsiepOQbZ4SeRShONAfHswF6T6+mfjIprYHE+q2wbi
1rcfsQbCelzmQty0KARC8xGSJGGrN1b8Ux9nUEufbDcUSyL/FckKxvDfEyx0
ufp3Fm9QTPQyk36xr4A0DcTk9juHKu6eoVimLHfrjmFykCKwDbEmAG5MvIGa
hRcQWymSnLEml6xnBaQE7mKA+YQ+SHikuO3aWmFeBggBR5YIiXDeCZqQaTuu
e2U/+qcFRkVzmJyQfFOwbWZjrGSdcleeM8DvPgwcEehe0EVNCVvAdAQ1X9np
nSqTnDUW8r8Wh49YIZ4RtqR5PJvXWW99zFe8kDr4sQ5CMhnKt6ZuIPXWKPEN
u/WsekX6KXfcJLg0BukS9Q1LYghqIokXRI7DzohV7MsiGtMqUpcrwZ+UB6za
LFVMeXOFvjAZxJHB7cdmlWGIS/YyEIcJKhhpQGFo3DnEQ65rV6Ts8lZw2MZH
ZPi9Utmxhn4/dWEIhemqYxatVS8687VviEIpKfyddl+Jiz77ac6q+usYdsy/
em+PB2Rg5QsHpGh4mSxslH6O40SBS/K9RhKtysviUE1lATFiLv2DzHk1wXRn
P+csRDi5XVlZgE9RTp9/gau/DthzGemNH6wvTnx6t64A+1PNSejfvT3D8IaR
44LEzw5+w1dN+KCHaUCw3AwUbaG3yYNwxH3bM12kz9YePxuFIroJgGCmxdh9
0/+rvcAxqrStekBdAOIpZWzjNUK3E62LcumwS9x4uIfe7b/tFugkL92Us9CS
o6upRoutiPgIKUSLSIbyuFnPqzy3PbsDFZZST+1rDrbe50qf9d0nHskLO7s/
uVadTlN1C8zVR4xK8nRdANQRGJgZJdM0FdviST9quCw0BhV07BKCzxWE7Luq
OV9a45emXth9fAzy7F0OVLfnMazyTq7ncZ7ORX21BJr0YwXlFQUgfxsZcHRs
WLzGo1UGLUXeOigs+U358RbRrUaO5loSvr+1AEePuzPjnH3Ablus/Gx6xiIf
ju4h6O+MTFx5dOImOPIoUxCDVc8HRSUYlXmxuGV5tVSHbqRRpfTXaI0KgTjr
Ojl6io0UkyzpJ2ZJybI7zoS+4AgJ8Ae/o5kW7G/SgfMP/6bsEQShvpr4tJoj
9SaP7j2koRFrPkC6LxLc3O3iQ0lpSD4RcReYxYogzXtFnJQQZJRyrzbh24d2
Rah0j+99+yb/SjGFXeeQCeNN3pYIDTlJMlJgE6KqhNqJcZ6/Nrl6y+pQizj/
gG6miZ0O4JDgveER/ATGRQ/dSnLCMpVLzBvAyyQ4EOtymb294OZwW9tPCeYI
HOzbE//7eqDpGsMTBkYGL+yzZAz94jaiYDaeyCR+EROX5lAniKjUsxb+iW4p
kMAaudAvS2l0OLOrJZChFToapSuNtdQuoriqdLd+Z/GRJzHexOJAYuTvGy9p
m8rdGdYqKso2Ipia2wGodEuZ9IOU1gD+Rb+AtErPVHi1LoO0ec6eOyhxm18q
r5HJWOo9MKFMKuBIXfy97ZuzNTiem5GF8SYwT/6wms0xqbgRD6A8+9CKd2gI
bwghtm0zt7qwQC4DNywP00bp4ljl9RHwqse8O0ulcAHDMTRNpFwy1p6n4cI9
kaAddq/9hiKpG5VSDziOyPL/SzafQU0XKF+tSG8B+zqBuLRC+9ywx4UfyUSE
F8kfbJVJH2FTC5qMhvHh+CV9iCFKWoe1o3zMfRgRzbDnBe2s7vab3Fgb7TrE
AcPC08FSLIU/UktKd7fbnJPjX5vC0uExdsQ9jvyraXiLQeniJi1m5DKByc5j
a1W3U6VfcR7u10fKomBlleJMR6z4VgymaDKKRFz745v0lJx1dfoYvvVP5Pq1
SHfWZ2/DjmFSNIc3I2wLzqm8ovPD2FhWo1aaAoCa0WEQ4BPLd6iOF/WR9KZn
TEVNYDTnZHFDYbomgKrHlZZhlaWs0T2OUyKJfPDo2tXu4Iy1Kt7ET6XjNN7M
wcraJ7bj1fEm7Ha4r5w6sCXCK8eibQbdkAT182TGPCgRSJajz4zifJD4mEPb
QYTbJuuHw2Tx4iQy9E3pxpCL1Q9m3tuWVsvTcxfbDo0mmzFj1UifITwlgk5V
0p8VXYkqDl7lS95zt1cDK7/F7dueD2G1YVZmlDeLzEJIN7kdchqyv5BM4nVB
FtY0cpi+QifKZVbAUnooyu1ouDkIWKdk10oaCT8mHwhNct6uUG0fg4LJSdXB
Hq+BCTULXjTbPihdFERcJ5CAXhX1erUXALka0FnuCrG46FGoC698i4/uhooi
NHqvMdT/PHBghn/cKAq9dR9MaFBdIUYZBYGGPbUJDdjjy0eWw2t2o44YpiWH
VwuZt1tJOt/jLeCTLJJMPQ+Ifp42d65z0HiT60EA+fa33JQwH0R8a2mAANi5
RcE22tcmzEiZPMczrnor1Vd//ZMnrGg9o0aVR5wA54vrxPHMFHzQD4dZ4VyP
SGICwGzVCeH1c9/0gWS8kiGKF0Itvqb46ik6FQu/X93ozd8O3PgRIxJqmwtA
fTz9C/U/jc/dQom8pN6iXkqybuavohaYurzz4rlWn6DHK8lComM5cZ6/Y6D0
ZCUtV6c/AV018xvPnLJ3zOWH2FXKWece2s3s7OJ91xAgVL7pwYg4uKtfgiPQ
jALBCPmSUTKQdr6GhIsXSEZC4BQUzQJne1uCBi78OLowKnXv1B/CnP6jQw5k
ALIJ4WGutoU5S3AP6Ur5ELmySJT0QqdR5f5ZXcPMsJIQhq2Hi+DwiMS3sRd4
ut548p/IVLs0kXRWkbGXv/tIbIzbzzC5RjSUpCLrBnWUFHZKvIAfVqpgZsrC
vvCI2BnV/FJrHmNLhvZxk/0peo1SCI2xgNVqdOQhK0TFO0vlaBS1bNJD4XSR
YasO5OX4bt+IQtjH2DvGkTuHibyZRwxNBcVm0bgTzxyzagBJnVDzA/X0zDtL
DSn9jH54l2WNz8E8NfpNOAGBEiMPJB64ZXgV2BFrTq4PpkuMbkv9sTuOH/bK
lTNNjLq6V1CPWf9oUfgScTLIjbAzHSF6y1Hwg4wMAQ7R7J6lrI6fUU/yw7BS
fAIFdgYT/y0Jg0lNgCo+X4ZUwZUtibCHRsh9ZXXDkuMiligNNy9c6c5VqoqU
cypjypnAkzElK8uBEAJfVOQaCtQVLCpoX2ZRkb0YOgOPj790gZGOX7T/HqP1
Jmg4O7O8By/8DgfxNIvVgfq6pp/Zheg5/wqk3xJ/NYyn8xVqMa4IhWmqHyS4
rc2kzPc0PvReByfVt9bIEYrvCeW3vttdmSKEK/EchrTzBZ6Eg5jmLILBJpWq
w+mqLrGuP8d2tjPv/SepcUcK5Ub0CxPDQC84bXm3hObJHNJ3EFaidUS9ptG8
ZC1bta4SQmLA8Qd6dGzFpH2zqbmgnbeYX1AySWcBaFKsyRTYSg2zM2HPORY6
qvBWBo2jZdnhwFPaIKS34h4Px6L7N/z0MmAajl/J+Ve9eVpUiYrLAimuS2FN
rm1svymQs3pVpvgRfpR8cvR059IrXjkh63ZU5fYFcd7+ODshDCFjaSKAxp88
c/Fejfox5+sz6NECyzSXgOm+RLf8SyTNS+Xwt+noF/d8QuL5i4P6hGX26PmZ
rRSTd298Rw5XSt9MeA6a64CKEGyfLWqUn9oUg5y1Qvqs74E2APJ2hwJhJnXk
bWtAsB4NffHj4HUAsVLFwvnyKbVTy7Zq0GSNG60W4gRJY8ltqrZYfHGGsd27
rwy4cgi3YTJLwM+O25Mw2OqN59gLyCVOGgD4WoATvTbc5mYs6mJGHMy14K7U
9TYoikv3KPpZ9h8TIzQTXA58x8Fa4wKhSQ1aDUAwsi3xE0+jra87MG3k9nIC
QgfhaM6+V9TtoM3Uc/wB2My17zHQnl8KEeQnGAcdl4kTehjA//UI8FkL8Pfv
EEiINSHcp+/exyU1blavrRKAn0uvkdacWZ41KUG1US0gAkvDeULfbYVIEZiy
u2oFKnZVh5sV7wf/17NB2T5nzYSAHiXeg+6cTUKWLKIv4EbBriSPtAfY0Rhe
0Noh5pZiD9hKGyh0s/e1fBB+Jb0X0Hl1o6ForC4Is5LQcuMfMOd9xGmUnaCW
Z21mywpFDzBWwY7WlfJaVcdp48MTw9GfouSizG86oY79Wwm1VKGX1nVdbTQW
gPdKyRLF3yqtyBfYDaJ0jSf+krskeZZkw+DS6p98jjZMXPQguDZrYgsa5REn
TlIorRIMWVcVpbn/A43A6SYvAC8qQJj9m/1R6sJyErK2UwCUrHs71wAJKybN
Fu1cRf9mxm0FYbsW4gTRR7bo+KF3L4squFnzg4GqJQvryuASRM6hb/mNKssX
+qrDNO+DIzSev9G4glyOSgDr2IjGl+ne/m/i53boLeg7NmL4UMHcQ9r+HQWt
apZc+m2zBn22tpr9YrdKQSS/582WI0E/EE0l36fODo5vVKAYKRSwejk5F+cv
HhwvVT8O3t8OBc1EqUWNp4hWrQ6YqrkRJFsruX9E5PNIxG3sM5Sjns2+CkUo
MXdJpQWgIEY/e2D0wNBj8UVXPGVvzKvYQz750BB3C1cftNZIIN2SjfcgdBj3
INbSIP/teXddyGHjFRcOI86BzWrbt8aG5J1hHrLgu/v7G6xK8klInM4AjdtT
aWU+RBC5lXKWQO6Pl3r+YreHUmdFfl8cLh0JTYatxd2qlJN+CO+reulkEpU3
fUinDv9dign0YAcuE/h3+PY1k1n+4wDTlE9DUMS4ClMmYUyv0KZ6RVvWsX9C
bJHP4wB07r6E96m3sNrKAT5nsb0efVhtksIMcXTkirqujVbennErNZDT/DGB
2AdCwiRgNd2MCM1dOYEOrA+JSEpfPHK21hniyeHeqWLBz21rS8q6Ugi9V//U
RxmcyIJQ6nJeSwec9J6SRwaTA1EEmxKWEq6ndw3LeQaP1mjb9crtz9KUsC4r
Ht0CjEKXLNt+1i/LcSM1FMySfZVNz0S4CwUUD+ouoJNaX34JSL51EjNK+fJ8
UZmkdHqWaGEIn3FlpEuDik0f3kQAtnj8+3HP72K4rxioqcsk6CYOkgByXN10
1IqTYpLgEHSH77Up8pMaovuyK+NxNlwWY42Dmcc6ZGL6Ec8qC3ZsBRDi0Gel
zePE988XEL+ymBkzG+9jo1dYSSppisxWrNgPuHbQQewoDgwpmc5nGuus8ylV
X9CaXOcBrdCgRgKA9Y4SwVZH4Bk8GWaa9cFvgvK1P3cW+n7yu0+IThijYPxo
Ouzc3ozbtzhnz+n0Jp9HQ5wyCP23XVz3CpCLM4NhEE26/zyhuZH9aUX7Rtps
Oz2rkFvfimFKgi6iHADavbHi/acCMxPcnPx9mm7L8pqAP9wTVPiG/5rCJxn8
hevAib1XA0vq+PJ9w0AYug91tzxm0LodRNHBUU3JFDClKnrPoiXG83oD1fYJ
QrYGug8Gl0FxXUv6pZc89sNiqtm3jZ8vzeG40ythtMK0DhPBAcZwvt59xeHO
Vo3kkD7zodS7w+OZECRUnqvclhSmaw0zLio6j1b5gYiZAQEnJ7qWkoe+o3bj
/uBCrXZA1lPFoxFG0iNfjIQKwGgKzzgqfkqNiV3rccvFIvivmaTPlFM1NVyF
VacbtH8xuFx+GyjHNQS3zP9B4DACOwdrms7Xg9RA+T1+vDihEd/CAUS2LooJ
wZ5iPO+hfW/QnJJsz2Ep6QKn3vP8crteqpKxR7aamyYY4hcN7axSEkZiTS/+
wB14GaQYgCEVdX5gue4N1MjMIurDz6vxp7jqgrNSTyJZHJYXvPjPzcPZTEv4
cGfd23H7kbS5POt/ZTK1F6JkqtV+0MgIEAmh4Ly6Wifm3x/7nmGAcTx7mW7z
iXbyKZNrYRDpvKrxUzZnIduApaCfZ6uyHU0xfhMCoqbfC/QLEy83M0z4ovE2
plgYbjMgr9nDCYTrYvbmAQmphhzpNYM+cZUhJR2puPnR7IAxHvwoqMBoYRBS
HqZiEGdc3bTXJp9ktOxEzPhx/pL2Z8h12+6EUaFaThjtkhIbxmDZ2CGy0Jm9
WMcyhth/7ZeQrOX4nQkCshPXQrCHgng9FzcUJb01Znq239+fiYWsaEjhNZYy
YRT6XyzIBpl4VkoHRGS8YxpvX0qrBOWbb0iAaAuEwZN68bybBGHzuWN9d10e
/swPa7FxTF0px647dhNEea8NAroY+x3mWRafwZ9b6Dp3JLXnZKaOgypfZLVS
0MNud2MOortU264k1ZqpQ6SPrKuvjaPd4Iev6c0AqGp7B4D2rQCS0NsNbkbb
hVrJZOhtXVfwtCu/nqh76PzigqOuu2TBI90zwon21CnOV5N6gHQQ2zZIjJDt
pJczW4qRN+CjPgEX0jbXzbDTXCKNgEpMrPL8lkjEZZMehxD3R6IcFZY89y9r
/LjBcbAroSg9eaxYG2uo6qBWqfZovGjxbjhGj1kNHNeo+861ljlHoy4/uhhN
plliKlAB3KJDrbgmJZ/UDLEwxQEe1RCTpTxpJLxQz7vbm/bRot3/8q9Jn+UC
PVZ15TdUZbE/docwgkO9aMTtuXA4Kce2hN/TiWmDKB6IpGXu7DJkq+atn/ut
hnqTnz4sa45zO8B5LvUDaEnJvWI5kyde0xHuj8Ow6CWm4pMaSs+UkBwr4iOn
0z8XNyHAQeAaB4hnbufxrBdUGiZj7ixUZVnNvsys+YJD7rtMUX/D53RM7xIx
yy+oVyHE1nkP+zhdEk4fClSi06YS/qIIqlf/mJm6yArBihjYB32KMGKWkeNf
/KJ4wpIqVp/F2Q/A5RQvqnC2Q0bUt/4UAFN5TTzMjrrf0vknEEeKaDzK1SdB
0kVXrubGsZn2uzfqaGaMiA0xnDKygUojkJsOo70gjh4YhUGVRBNZEaQbWCYm
sBK34bzzqq8iLYMs3zrKK+6YVgyCyOtTLUfsZUje/YPeeFCf5fsbD63PobV8
w1sERPZV06VS76TMcYY45ydmo3Std6TkjSBSV0JGSXFufeb02l9FnkVm+Rfp
hYVZVNXevwc4I+JyGAmkWFn5tdsdymJ3QCaWFjxr8tBNGlldVVVBFiQlZ4ly
Fh8ezrp1DaGONbRuxNf2RWmy/Wim75UEztQohPoq/pK9OJk02vgj+ume4ioh
KM7x6/UdKYiidgSia/72jBWMdhlQvi62N3ygvSvF4Q8i/n187mWClQBaPdzr
NPoN0qSKog5i6GDbqGDpu7Lhs9y0vrYZc//+8Pk8vy2qQTaVNKDRYVUEyTpL
51gb1HJL6lhOzVK329jBSkxV0PTLhNsAkCDgntNErMwt1tyEBRcmt+am/bwk
RTjUX0yecC2shIcpWWNi20vEtAEPBI1WGtp00hzdZjtm+lgAX0qsM/jQs6QV
B9ajcXZA7BiQPHtIcbXsz0HV+F57tuSZUwroG/dArgB42aitI0QFi6+EdovS
4EkJG7OxySAyaYZF6i2QrG+YjmcYeDFD44RvWmypX/5BEZ4crjsV7bkkPGX3
ebvsjatYSYSvgqOmdBaqpq2glOs7Yy7dJHD17JFY0tJyaZMyJ/7jTEQF900X
cPYfSPGv3/DghXgER01tUOZA28Pt76boJBIm6FpMkmBVtaXhqSlXoxfFTe+M
UaSaTr80cd0qlvRY6h7EIB2EZ2zrzcno4qrVZSdu4FmpEq5r8QFj0YWIuWKv
vjkbQWkDaIS42DyhW4m/5yX6Q+wpC6PzcEXLW5Mx+0T38YHutZ2g77uyJZQj
Y+79g9+AkvqUZZrdryMX+Ix3rv1pt/vuPOBESflmkCqFMqMYBcZFQMtiLA4X
ZOGiVXzEvqbv2VYckiskxEvos6vadiAzWyVOFSyW/ZCLNZkpCPjg9oZLvNgx
2cM1RnBRptSY1eIlf7qRaJHGK3ed6yJWqFx3pSG7PEf8CjjxXrDI/k05i3Hx
Yq3M1LhEp99Tkl0N4kuanznvrk51uYNxt1idelNAPxCcnsVLlXcZToUsy5PO
WoQaNLmwP5r46ukve4XI6LyNqSTn4Qg1m/bPWHn2GOfdvFxE+gPaAr9NU4en
bSpQbZFl0Cn2oTgT/3l3tLBKt5SbMB3JnTXxTOnE8eJo4oyXXsbxOqDmlNuf
60QBM4uspB8Rkt0mAE/fWi6CNZotdaw+a3tCdSt1v0HUeV/LAz2+fa2giBd4
gNHi5a6RMm/ZrNkgaGacWxbBmKX6K2sxI8+SEX59z/yojAgJyt/3ZdHI169L
G2UelrhcgtJvEnVDR8uXWD4sjCxgPR5nGQCg/0ZUaUmCOQHcSKtWEtP4XwQW
hXkbA0BYE5PuqvUZWMG9LcvRTH0ctyAF6GKCqJTJ7JDfsFfW4PmN9gCh5Dgt
CzoNw72kmJyFOkvAsssLIrWCeUP+0pzduHYIwloxvgdACJThsIMWy9c34e5Q
uTXPHEXpCq5/TIukdDZzGK3VgE1kIsjcRM6ukljqu9KwoXeZ+T3fvg3fwL/Z
JjOh+QhGSBsz18/ZH73KbsxGsrAHEs1Ollju8eZ35f8o1iIqFXwhgNuv0fhz
6F5S1+juxRD4wPlJYHeTAO3YywhIUyPRgaa61OFYkwvHPdSCF/1XMAcLC386
dNiqZSC2IjeFEmGjwaWgxTefylGmeDgX+gN5NdiMg0+PeZ3zKpbkDIxOly8+
mC9zi17doPsHT5Gm0kG+/r3F6ecO28E1mocUkcc0wkdSUeSPOVXYVJqj+SPl
9qIMABBld9jB4LbusQogyjRmN4IvF+EBKEVPwSFTddZhxMluD6TVZkaMpxND
TwSb5UZeBg0XmJ7mFnfzVLIwhHODm2Vfdm+wl+sKVC3rkKoWDQDdpJGgT77D
WaIixBY6rxV3HcHXuxS7Q/ygqUef61N73htB8vG8IJ2Lat9lsxJ7edFsLN17
BH6UkOq+wPAmMd4+V9itbA5OP319D6CaJCqKUw/B15jJBACSO3KA3zcZLkaU
l+7LxYZL9ce+5X5wwrodOXcz1qvxIgWBFzqjizB/2hSzhu8Eofbn8DgDoHtP
S93YhZ1+AztdkilCPDHsAJ6/jmAK7IWqX3v25jjVb6YtDZjUmH7Y4lZ0xb/I
zB+V2BcFxatFJhyPFkObcna1euukafXCjEYPhbNt/ogebfH7YqwmrZaZfciC
BDzX+47/nv/ayNkD7Gz3JZnCI3Psr2RJbm7yf7gLhpyDCwjJwJEMbDs89zS/
F7AVTls+7GlRaeucCncvLpZHxNaVfudum3kkTvRK7tozOp2tgoCGYBFZTPkx
oaj5CoNQ0oPLsLYCstZjedR8WwIHp3nUvdNlAS0qZ9LafbX9GSzWZ+69KmTD
xn443IbQX8rDeftQmXI22aQbPzrHFZsKRbusOu23wFwqoGI6UMb9rLf9YBrD
aKEOf92/o+IzTId+VZA4LRN57hEZBcB7G92UJfX/WHw+twHgmrcobrBjsQgx
+HsJzkGGFyqG4bESnFUwuq0TZY1zPqJ6JR9/eyp8Ej719biF/ck5Tr1BpNW6
FwRZbPPEzTPk4R4VhLpF1+VWaU5KrxtPszMQQ0C5dZ7eIKtRdrE57ZalOnNh
J/05sCOavd1wLnIznxRudGiIel7t/wWdZJ6kp4BYpFueK8duJcqjizXhsN4T
fCazlRnFSKgaz2CQ4RoMv+FborpeXSoaEauy2cU/7WD7a98UaYPKmgMPACd7
3i/5OUysxAVVDGPKF9Z4LQes2Hqng6eCjWJ0q8mAnbc2Shbx6wQ7clobcSZH
ZkyOEjPigUhz8V+txZg2zq1lMEkNuTfHINsx2TMc7eDECRxVRQKvN5qj4/jn
hBK3aCrIaT7imSPPJUwH3X6WsQnj01WBBRKfOJrFTCgpvclh5omYdjZPw2Yj
Hlgm2A93P/Sj211xLPOOFnOjwQpSFCud61S8azHs3OC/k7EvtE9Vrj2wn+J6
S5gZVTuAUMq4wMhJXHzejJAu/PEzSIxkLPK6M+jIOFzhL1CbIyW0+yrt6vfy
RIqTiFSmMFf6xe899hZ7rKzvf6j4uGWpoi9/XhpgiL3kqe9PTNTZLoKRz4Vl
lh9Bt1d1QHWhDZ8s/VYF4bCXBk7pevKT5Qa4BbmnO0FYJYrT6BfamvccAWZV
6S5FvpPEMtdi5Wl2zO74V/GmWcr9+qlh32uLzYezA9P5SoVnba6gaQ5Np8FE
MCQ6PvGNrTTmdbBxZoOcN+WSfdeJvbReRkayQxYIAtz9bpa+HoqXkFmkq1Px
stMBQKQEpgo5EuV+KEeSW3Fxa8sdNaLZZbmtcXQF3M9mHGTiu0OJTN0qBkvY
L5Ye5779EaXRV60CZu3RSD69pjFi7W7w2sNS9TUH5PpCrwWQitNK9n6hmukL
K+jgHvHUAXCh7AvNU4rZPEtYqZJf1mhFZUsotXyrHQ/ha8ET42ynt60NM02C
2amzr38Y6DiFQSfRYSQxC53bAjkbYYE8OnMaQlkhByr5lNdzHyqv9LyChz2M
qTEK1N7bbfvGA+6b97XOlhfw00rENtOoOi/9JcumFjONszeUdjE4J3tNgZCo
groqrXmxm/bf9jLwj69DizQrfcaLA0FeiAv5X+D+GHKH7fgo6eN9MeGYkwxw
ItgXxOlJHoHWTPtTUjijJU3K7jq1WzIz2LFlg7VPGwjILrQsJzj2OGHU4LVr
gqAmxNCPX+lepA9y1HRpuI1NfZ3uUAtlfTFek7Vsv+kyLroxKlbInGYbE4Ot
HH29lmfCw9gSeMeKThBki7G9wDTwdO8whGg7WWc/OIdLSQr4FxH+lZKq/U8p
heqHzVfytx2W5Dir3mj1+w0kbI0C9auDXznz0oSjDBzbizCCO4d/fVYL2zCp
WEEh/Mel7xFUs3wsPRXeMsR2A2I7LUG+W3hTGovhPoKEHrSiEYLaWESVpNPL
HEkXX+i/9oHGK5aXhQQloipbSk8mqvNA2xDs6notG8hOYsarxpRwIP1M+jwt
ul7H8Oj0wjtvXYyK8MaFLZrtFwfnhtP2LNjTas9OnrCiaXq2GSr0WpIubNTd
SwzRJi/RL/nkf42Bagtgb+ijwFPEdMv6i1NsUiECJkqbrifkXJrMrjscUBi7
jVD5NSU/hD5bPWy3Zpw41jyNZv14OHtWGFwC473Ag+a0yvQaick3fElmsUC8
TNqSHiiaUrdDn70J6QAePCaDMaDwdCqOfhOjO89czUm9KJtMotOCd4/7vnvX
3mG7Pg+LhGI/CzF18LluEDO9PGEduJa6DQpNJWLoV2Pm2Vb1i8oyem9zE7jT
mmlvMZ0jqKHsnvJA2ku6t7UAuC1jh3YkdfqfrNl26e82XDjqzZPl6igf55Hm
JTgXQrG9+r0YuLGJko4svVY8Au+EPRCnfSyI6CJDWIdgHDgWl97aw6yHLTxk
qt7SCAlu7PYA9DOz5CAaUfznL/gDGTfyATBpMCjDCcB/kvcl6zI0/IYkjPXJ
ph7tmEXRyrvqiyL+s5dCGhzabkdWqQc3XayiRytKqGFtYzbc3iHFgaqoUpD+
0L4L0NwPCHQsp3DnN9n9NFBngcQGRaFfOQz6dge3SSL8UzV3452bD77r/0im
7ivdhXAgu+i4esC9kKZQyuAoR4Q21lwUy6lfmNsf2S0LyJwF5oB5HS78IaI3
QrN1s+5sigt0iuNYTDZficI7ui5avaolrvmlxCgdNv67RcfjxrDlepo9Vlll
JowFYmkhtgRZtajp74yw6E/StR4S+5G4WrlJexChM8BBCYj7OfxaWYGUIe0y
y+jJgWbkz7nx4mcQ8bO9N98F/l/ZVdw/lA55Zfv9PGOLPaJ2rIo+KtFQX81F
BwFGhZl0PJQptCGHE11YMO0aNA9aDriuPtnlWDHgVcN3AYMNjK2UeKQ4I6Zl
hTIJNcq/WVOV9tTtCuAK41h+h4VkhLKYxCDOqbKeAtconkUdOfo6aacptnM/
AtzDdx//2DWvgftOU66PFjPM5r3mHc0HpczmZae58MdK42Rlf9eL7welNUh0
XOS2XmEIqD5wI6n5JLD2SmcqUGcn4uatdivPTjeOya6TrzOd1Jejw+Lnf00m
QmeymfbhLAwo81Q1a0Jfb+5K+sMPbwpbTaqFCodqQwP3upGbl69M5rAcuX8G
prvEPmHSrM3gasHXgRVmHGj7Cc+LdQJMhaFa6BXCedN5+sgWpjgvvjFBypk7
sMNHw6zOYu69dYOEtqfpg8gwyhXRv4SsDNnrN/sAvcLZybZKKMoPDYrtP1c/
owCHxt28YYrku7V9BPF/k8+RLxSz8IqNdcwDo35CiCYiPwpZVU9b9hKQGbJ0
3O7Or08uotuBrYabCWm4UsRV56L5S+YUH3fRTIsYaXQpk2pqvSOvgpnMud0Z
j7nNkoiJkt3EPGpB8mOk3VgKIEY/keGE4cuRX1+SsIioBVKeNrM6ey3yfzpS
uNDTVeMvbojeqZS68VJ2yrvEMBEA8T8UKDykJC7fSccTo4j+FuwEs2Y+4bVO
NsRmh89UxZHAReIw21wTMdzhVGNyXrGdnPu5sJpnNTptmPkEiHAK4ge2kq+K
daxqlSMmCn5agtAUlbGjAdHJD+9GCgtHidOdC04Cu7BExE7Yh5ydqkUFR2KL
NR+jobgkXgGOaGTCG9P+lcRnqh10gcAOZrlKncPA6fuMfi7qAtuCQjsVMBeQ
yFWQJTvk5CT0hMinr6uouk3YjLOO2I3FT7Pqkz2ixEF6LthBJe6iTzm4gAI0
mO4jGpYua5lxUw1ECAxFYZGiDOBLQIxoBnmjlYhLLJZMRaQhhSiT8rdbRh4Q
NELWWiPhNsscJW1M66SnnhJ/xpXY7ZZPfsjZ4RUj23qFNk0Ap7b85FWh+tuE
dSvZlP6ipXKGIEMBNN2kzo8DVL+p1YalkWER3DlR3E+XdfmQM8o74HLkIwU9
84KQu+iKNDZKowYm6qKjpnZ6IaeANxs2w+ho4hp92VSxEtV+Sfk82VPvgD/i
YsTW+GR6PNjjP1Q0Bt1Hdl0fqQUHppbq0xPBbRrD2AwNS5mSfwnZm2KivJ3N
KD4H4ZveJNGNgky5X9wUaAeeLr69eHQH2t1g83eCRA+8AualAQWyPlhAUQt5
hpw0BHOaZg3lmuRYQG1v+plgVMsuk/8FoEmpWWA8f2JSQs7pOsQpNFJS//La
70mdm4UowMhL4sHTLlj6hS0JtklYD72rGPl4aJ2BbidssRbbcSjBZIAUZs1n
k6xqm2x5JOJuAbxBrdRQnJzL+HxBzHTI5PUHvHKfKoVreh8U1SgZjesAKnzz
AF9/iWlie+31Lmy3IokEaBgKas2JoLfa9b9uwRo3RTTIIZkXw/NXmAJuVsEP
CUwaRlrhBnPZu5EcU3zC02nHg1vmzFhRjG9pBZv4DrihmS/uUOgtkGYP4BlF
NsaBN6LnlXVMspyaZ5UAb1TBn3ZgaYpSeUe908KCRqz6L+8tsZmtzpeI/4CR
soi11RINVMycdTBuSmiYjjkKTRjg7ReuKJzZShDfK4aQWSnPsM8zWNfWvjjk
u2wjoe60DNPY6NPRTRTFvPdFKloj8ufYtNjZhaljwGpRdFHM3e6P5NuIDM3l
i+I3Yx8XINQiedBrYEJCI+GV5a1MEsw72oxBC1FBAtKSv21IW+C3X1XxvQKA
B12I6tZ+ZCWXu/MRVJRPTydK+80H94l4sPIK9fL2C1KIJnSjJ5kMsfqV/Gx8
uO6Ojrlzov1ryy4y/TtvPmenffSH8pPSWQHakjpMc/uKoxAT21gse5eX5R4g
+Mq3U4NfajKUnS/o002h+w8vqR9rPo/zkslUK630HoQO2YEbTAC1OkZmUqhA
1xIU5t4jUxYVH/zmfGR8e9gTr65E5cmv/lQHf9gvmG3jyrDE0bogLQ/q0fVP
SbprsuklQMM/IF//11VOxWZdqSwypcFEqS1zQAGBmfD6/VDZJ+3AmhNNiMMD
2RblgOPpWdXYPFcsLYaV2CaxG+FAG9UmUjXYowB3aKC3XUtiy9YkS8PM0pxJ
va7jPIRb9TGXV86gAdv7u+RF386B+YLcyeeocvv+KGVVmG2g/zujAEohfY12
jRtWTOmsR0zl3VLJYtfrarQj2xacrgUSCY/9Eowe2BNa1QbanKDjEHxpbQd0
zE/cc9V5E39Zkeu5a0zTJRW2aUgqWLV5wEaM1K8YrIzASImvpwDUBaPy5K3J
k1IWykUApzwmYmJ74MlK3xZgsodME/rj1aBwCevWk8Qk0bgdviBEuwa6DV2V
d5VEsy7nlbHzaQJ7H+2KiBl8yWS13W8ppu+YuGlwMeV5hxfekg/4ui5OfOd8
xfnoy75qKbl06xZArGVY3WVCW0acGoUQUbuV2tI8kxCEpijLylsf5cj/81dG
pDPWTa4njnIetGf7wa0heY07m5IM9UPPAnvszvSkDOjoyOVSCrPDwTN4MkJ6
602LdWURoS0kttsA8Q2XlYxMqS5fe00GtAJSF0YLX+AUtWlChIDGuWWHGkJE
WTxqF6gEUn66/zpVt/Znk+P0TbRmzJLoAZWyaUaH6+WECr+LoGFfW7OAydNa
t5iOiThPTFClzlWHNp6KEk9Um2KV1MPufRjF3Bjyf6poKPwXxUqNOfgL0IR0
JWmRX898fQOK+BcHOgWSwgBX3v6cdCyv5+jBjp/+km3nPIAadTbBDqs0iz0n
brpEknxMLKg9Gcef7K0G1BgDnOgeHBr/y/mHORklRKrpiezCn3JpQznMR9Yu
kNmHZIYITMrK4W0ZueWLGEZJXYeHzrI4yfoHBzruxoDKL40Bb3oC5JyaIlJh
bQ/3bz2sEbdZ/IzmUBO1hl/e2bNkfN3bHOI8agBokXrZDb4h42MAAJDaUYYD
SPM2LSLzeEe/+ElLTb39sqoRjKfVwkjIyd4uuBtQeg/k8DZw9Vnx5QiU0tio
3kJ5aAdzDnalB3pBFQCOb76DMvazf7H++EVRlABYabWFdQC2fkIRqrlDtiB2
ploDgRWuT7hnamxDY4J1Fq0gbHyy7QMeX9jLrM3PzIk5ZMAPiEsso7ytSBmF
V/qLgXTTkl7+Leqx088eKf5J+zaStMXp3HMS3zLyOnZwoRdK4VjVktAfkUEt
5AH8RDnRzTST4bDaOcMTSMAwXEDwD10hO2E78txk+RlUQ/PO2fkFSc6CSw+s
/jFDoPbRyxN6rbOVAR31yN1cV+484kGY+T/OY1Xin02XmMTwI6gRkujU9Hrx
QtskgY34nZIHqxX86tGTP6Xqe8QFVOtSrm26dc9X82ju/O5rDOBQbG3gdCve
qXTClSBndXrg59VNywMckSMsEvzc7Z1EAz/VriAZwk8n+NBSbHFS5zCfKe3s
J2nBuJ0Xsb43c7cW8mQ4+6u3mgTw6hkpZwCc6VPPUg/kv0lFWKBUe5/qKOth
EkMCXkx5oddV8EFcfmHIT0QQJmhMgRqICgtm7f34OqpFBCfLYuOaBjSRRCPI
EWP564CRHOh3aLjnrvUM1dDjtqyt4nc7JYv9UcxMwLLyi+BnZtfFLQkb3IA4
bb5xMxI4fojOY8s5tSEGKetAgkqmzF56U4v5lEp2/Aj1u0stoY2fwDgc29Vp
qupbi6qTtkhUEu0wHTW2czwS/TNM1EpIahq3xopNWvXOjARVurX0ErZ5BtRa
stgOMcuqT7iNxmw4hjbMrEEyOfXMMm0sanRvc3GaNFhlZXgB9YVqPFsELdDQ
JI+H/fIsXTEfo/66YbBBHmhe01gyLHtoPTayW2o3DY64wbd9z2N+Ph9xRRZW
vXtyISrRi/s9krZdvacN7MKvZ9HMIr5B0axETh4Ma3Uw6km0rfkG2/hvI4J7
d4tHxHjcLcV9OGK0SBZnIcogqNfeuQ7FzRhKxdQ2AlQV7eeDHIdPMEU/mnk3
eVWHKI+hixEGZKG6uBEnseRVEu0hVobJRCyzq150FNA48+uw9QqBv1kM1eoE
ClcAqKq5jSDWuwq2h/TScJu8ctoAY/k3oY9D6udkKnSN9bbZ5fcCtmPPhkAn
h7aTWZ8jOzlwzAkOL6AwzX0clCgPhw7D8v7eK/tpWitziX28uBhSx25RxzkY
m8SrkAXFKKSlZlPIFjE90OOHeVUZNR4CuTvVm42VqXST9dJSJV048LfUTAGd
b9SfunHyUE6z/X6k7U9XA8Bp3tZ6SrFnsdHCaNJz5PLL2hFJBKU3yTc3iyoL
U+SHJ3ErWvecKhEO/vyb3SX7xYnru2MapAC+27mCbx8LsmEZFGTashXgpMZ2
kO85Iu2aXk0Lo+/Hmbx+B1DoRH4QY1o2IfNNBmmknT8GCw/7dbYpm267Easr
09lNgZaSm9TKwYxmG6n0I3nqNn76LtpIcQ7VGOt4E1Y4wobRFgEjKHAopg2s
6UmJ7m1XVsc2yrUmSKt+33z7yj1KNLuqse0KkyI1/n/ajvyZqOFmDlhODGOa
2BiC6Z1v19+EhoNyjVcM3QYcUmeTB29BTN9Qq99ius0W6WSoDoTnZ+FO3+TG
esqAwT2pmjJT0HMRacHrMoznV+V91i3MZGyk8gcDKXSpq3EH3ZX+lWaWbsEF
TbxEik1yRTWgSxtyue6kgsW1TysUhETfyceA6tuUxLxrsbDj3jiPMlt6oGCt
rG3Nq9dZ/y+i1vsPTvoSCvLUu76ENCbrS5UsLGnVe6ON2ljOWU7hceUVObeF
GalGl4xnonhE5AWqzXHjyKgtNguKRcUVAVYaIR1gN/DgkUjnaFXVMXiYZlZU
xJ98DfxJB6gtmRSLbzTKlh6limjZ5QLYVSNGF94Z0b1qusTboQZSCks/BioY
y9qIqGEMfRrHHDQuUqBte0Moth74ywGDxDyKZjQKQ2PSGKRfcPkkzCEjGkcx
pyiL52GOkz0N7K9yKxorYugPAqnDiBxFK5oqbgaoom605QVmNgJnJ8/VrYW2
EKQ86+9ltYvt9XnCQq9N9RJxUDhwpw7m/4RVPBjBkYqgXH+DjQI4BC6aeZ1H
aAvJy8G0DrYV0tSzngQjM1N4JG1Rlpmua6cgDCrJSULcB7MAeWVXU2QIYd/k
xvkP4DGN49asxnpRmoMMpL6ET5qWaTcb2yao/ntheoo5x6/xXa/54Szb4QiY
Bwa16cmxTzXtVtmQs4Un02NGcwX4pOmIjIy6uxCOUCKnD0BAvz8teaS3U0kK
vnuzrpRLRWu0MkYAxsR9kMft+0gEg9uVQPI14PIeCibNrtKhUT80fM0yuEcx
XlbL2OzK/66FfX4pWd3a4E+tUzs1NCfHy2R0Tx0p2IKd6ij8isARFRBjHirV
cByrr932NqkSEA1dSrWC3pEKKi0Wo4bpbKhqS3pK61k6A1+0OJqPP5M6vpTB
4fFChtmivel8CHC5DwRTEDq4CHOBKUkwzS5AhbZiTxyPcZ/DDkeyjRQaNTw5
TN0GQvHCful1Wosp8TPP7/YqOIerAXRZe4U6cxDHtTlnB1/oEqq/zPs47I4b
HwVxadWMYtdQubWP6Bkhvf39oT04xRkWutAi530ryJiK4TMQ7WadKWciEA4/
xKNCIfvGh4N4q2Dl44nQMwIrGk/+b9nJ7UWZA3chp43ewn1bMibhRlU2M+JR
hkh7oTFM2FeEWoBJTe1LqUh971EVBCqWM+grU3v1XO1SLbtGSuNBakSPKeT0
NZKbcu1nzuFc5vXtJ1YjI3xv4qRD+I7cXNArKgv/QfrUoplk1rKX3lwmLqTt
SD6GuoQHc5ye1dxFkiIv4pdAIQGAbK0bAFMmbY/Bh2ic53yEI3H3l38jiG58
ymrZsSqgHjNk4/BCghbsaMU23hY1ciFN3BXWGLTaTlfVSV+C782rE95FJcoH
4Kgz0lufkoa3zPB2m4N8GCG2DAJtIWo1iOk3A4w+RJiwU3j5srosCiNmmDOM
9E43vAZNwQyywTxZJZ5IBnwZaj2sPOU3+twmIz5WLfHp35XTBVX9CMdXdIQU
1PVN5r4N5Ma4Lf9Wdz3NfAVeUwvpl7UsZ2x2m/mFxocvKrBG1bWfsx/yOMn3
uay1kQJ8XsFfv/5x9/FcdHpg7YrOOy3b1yOJsp0YtynDRt9QRjK1kcbAIKvY
o4p5xYVRl+34VJ4L91BJ52SumSKWWrz4XpnLzUnFjIyNZdGcSdn/wgzcpUrE
6Vu5m7gqk78nY6XRH41NE9g8eaZQXkB11HF4n1kSy51kBHYmR3SnyXptuq0n
QI7Dp88KkaL//IRX/XgDN+KQK2RlAyvF4RAo3ZTKmQDXFyhIwgVw1Y87QCO3
LG5kJnYy0b+k3QbH0p+7DRl2dXgCZHfMxQeagAs8y/fm5CJTTwJWdtS7YyWr
tEUfRBGiNjzywQw5yVAzC54i8ZTo/tztON+DLHH5MF5XKZCcW2zeparsEyXS
DqRoijuq6KNz5UbP6fqUqzxa1OuuxtF96zEPPnAhsbIqvmufJag0CSxhOHS6
XSPThXZnO40qX8NisEA6a2G8H3LRmH8m+EH9yZc6jCfTilT6V1ZDKYt6opJZ
zfMdb7+50LopPnLKJGmB6pOZFttYeOiK2lqFefP+cjPx4nWxQhMVlVODOLzE
GEJkhwDCfuT6hwxz92Mj4gd5vQTA787mhCNVxD1dTssF0NrE220eKvnmKW+W
iYrQIr+VJQdtwwbup+SSzUgwNkT2Oi6UjMY+BYySwAcuo16i8dJuMHTarsIe
IFQetgW1z06jVgi4D3FTu2Rjf5wFSTwPAad97YekHQiy8r49ARD/7czNJBVd
9SlTbT4UT3NdeYU+U4YPjcN5Bhr/Ll3dyheGjE9HgmUmZhjKLwXdnghbB4hR
d7oj3lVrxABiIwGr6oga5Mjp94TrfGozQOT/qB4LvtrjAQOGF87dqmgY/UHj
+mngXka8TraQLpuY/gKdOv2FnnbQWFE4VTbuUqdXTm7XhpF0xXmpM4YwDx+8
Q3Kd4GssUSPTphZJDdNlJwJKyceOAZMBvVeV/pkhr0XTOIDII6/kDQGbvDEU
vpJ4SNrOMp6Ri1fy9zolPezc0+8zYFSotEbXiqXAeGQYkMXFyMjYQd/bLuKi
fXEW56Y7Sol3/eLKImFu+ymed67kt7xAx5vUprJzbXlhV8THGo+tRjDM3NfG
I3ZywL1zrgsScJJWg3hpYoJwkmnauBy8vgDP849Pg9XsKxKuqUO2HJV0sHSy
NBl/5nrnh5hebfg8lFAuineTAphQpctj/tb4cqaq/dMNXmREF6fAZj4Aiuag
a45oiSWQ/ztLYlIoJt3uu+2gOx4BOW0iCpdc2aXEb/uy/p9CeJg8wYChtOFR
dXC/oGbFfP78VAzMk2XY4Va5Lu7WyMos0Vmq40rH7Wyz8m0swdSFme/8rZ3W
q/UkkNjfz2GMuiI4oiP5fooCBljLV1QTp0e06oa3/oAvlwMm2IUE7Vpux4jx
vnPbo4i3Tk/AAMg92WrSDHYsdNPg+2w9K9BvT6wCJF5o83/hNppwW9tmpgUh
kCxKTK183hFw7b8pQxAgvLDJrge7ELpFP5LEW5sxF/UPUQDbuD+3IwyVtaWx
sA0KdfOEfW5HEwSlp/ali66h+NYDHqGVbB3IEH/B+3W5/lYnLDnwAFf5Yjh1
pgcSOfj2lLtpRzZcy283BNRC2JivMtR0zRmDmhD2PODUi5tI02iKiqmkjE2M
ehWn0CmmObbAWLQKFthQ7ReGLQ5C0xZm9Y7/olSLLKSjVxNJhbOQ2m/RdFRK
jPh4nOtrZ9efObYqwNhNS9rmm3ZEINGNi2Kmsuf4OgoHqzgIfKTFVQ7cKfUF
svYT0wN4bJoDlCZbO1ZWkYUTsAQHo6LgZWe56iBr3+WJWikCkJjfeQ3WRlJ8
KI0bO/CwO6F/iGRBx9gjXovVsGphZY+HycCBD6eBi92uMWEMdUxHxfDJAm4+
iMvDAXfJqvD1ynd00D5bD1SId9OYQ0+TBm/Psjkh/g/vclVmf8gvgpYDDp9r
ihZTADuakdCXjcTupoEeiNBbx5SVT4XqlZb1MAx3P6+f0aCHm2/yKZfrITSc
KfjfpY3eg1VrC/nyMRLb8PdrynCN+dJs/8bFGemUXI3GSLDX5sGrtnle5StA
T/rq4QjkcZfmdpSfSNwXIqGChwO/CImr167t5HWm5yo1whqMi8O3FVLrqQD7
h3/KA/zxoSxtEco7gxbMYQltrIAFrzY+ao/PM/YN6jaGE8bJUBsM1BHffNR3
iueuR3bOqWmvLpE4h/PnNFegGHm/1ce1q7Nrc6jhKkKAXoajPJQPVKAkL7JG
m2v7phQZ9euiJZNwf0HLVqdk49kCZtDdvAn+T6FrkYbGrqJDh9HCysO3JJ2v
+o4GZGWrv0KoEZE7F+C6SaGihANyLewPEghC5OI3zy4+O2lNsfl+ROF1zFcn
fGox8+bFH/Bx7N4tKDuWrJQLIzc3lbHQ1tNNGocWrm4QC2k8FR5u9YHOULqZ
supL8bXShUGg4R/quZKm0o1Zv4UXoHB+TCaBaHf/9ZtUi5REMQQAn3NeOu+V
oxjKmsHS4PoCdY92tIEgjFbJrh22PDpkPVSCK1iGgY1RLcDtGQLBR/1Hq0AQ
YIOyBec8pme5KAie9jjglt7vfyLrdJl2V5Nydbgct7HauMl9vEQs7p2Gf8wP
irjwCmyKBexUKIjF9zbKkQdN2CuinP7UAyo68X7vAtmsrL7T8DEocfpD8cnT
+U4ik68pHU8sToMEQaGHhmUGbGe531HYXRn6c1nkLfEngV5Pf0leLEH65puK
NWIsKXhNnFA5XG67oiwHFZC+jjItbQRmqV3BCi9mo8tLW3oCYZH3dw/A7rbX
kv9Aq/S5P54QrIaZrs1j+Rtu70LPEmUjtv5Xl0oj1kakCuT573cWLImR4kxS
pjB1S2aUy4wQlPWM4+rBEjWvBVOkwXYICxCSyiYq2cWZli6z2rsVUCkXlNnF
8czMgNyiXmhTo7LIvmHI7ZPm+cI76c4+Nmtjk/vjH9G5I1WOD3EHrdSGXAKz
9yR+gTEAAsAORCkwWSLaci24d0OgueShi599FZWwTHuzjjjD4Cz6jnPe4lEY
MUuvFlyU3jgwMtvoeL3rA4NuzlvV5M/lKkNlB2wUdpD5k6MvwM2YDaQ8RM7X
wBFwhzL4MYSZIza/t7vQKPSpk5Pik7rhernVVrM2ZULMcgoeaEJBNDYcrMoL
SZ1MpwdnK9h58es+cl4d7y0285CK32xSYaQl/Q8lB/sjjrS+OYlbvUouixaC
ZVfuEYwvYipoie+o9+YS4sW1OakG+GJM6f21JlcCebC42hquE9qBkl38M4kA
EaENp5CR5+GIcegJ9gOpm3BEJP1nEPjCekTNv6JY2CtE6kGT3CVyZBwitVqU
MeuH/ZH0f/YrFBFTKwlcX8udHFIZ2+H5MqdZue9Mt10bdrvBPpUqTmj+QULj
xsD4pZzsQ/w18E1Vj9rp1mW5egLYMPElv8XBO5Ek9K6YYSu4kMBpqbO6tH4d
tW7J9YVUsudQfwvxpgc3rLcseLRS6gLfe6xMcb4EZ0B1OvPH1ICm6vnzfcqE
Zm2JCQP5BoHDNM3OJH/bbP8ieRI5Wcg4ZRcsn5m8wS96yfNoZ9jSqetzswFT
UTJ/0yXNGbSSzSIX/UomrHSxal/iH2jZEiqQOZHg9V13MD/5PoiIlfy5MiRP
QszgnJs6+qbWUT+D99lWkzyYXHtig6URXeguddBipRQazSJ+48uiefHQGand
ZNIKKd4nFvuohpzOSvCAetshEHyYUT8DGLDImWay3Q94M4AGVfKFNfgW2pQy
d1+e+poIBM2BEqRTO5LQu2OBK/UlOp9LDmGhp+2iV8EYuTk5qi1JPN1vDgTo
7t0GQNxIvrRYwMjxhbRRgA3g8g4YTD5ZHr597mY9qobwy/YQWqCF1aweGbN6
OTCiI0OFcS1F1P/i4hz11+GLtguGlVJVlkb9NV5pxynP+0lEEXuc4FxGb4Wb
C9GmS42yMP3QvJsS7+7Od/TjXb4amB9Nlr/Eo5/jb5hX6i0uk+BezAoX/UY+
jg/GjL9dpBB683Scl1eIDNpehUqkS55hpemiM5rs+CxTbak45WtNDFxOuVfT
iby9ixITyQmBWN/iQD+2QjCjimMsbe5Jbn9eTaK5BMnAzFGiadLVQM1wxRsP
BAP/0AGSkfko7KNT7ZpwklsUpyRK6jXtYpOofk939wyNc29Bs15PAQ0cYIpu
L68JsCNd5WgXrQDkeVhHFbhPi9H+qhzHyUa7TChTcSu6/qOQVSzPGmcA4p5W
vA3AQS4cYfdZTFeMBDxgzaBs3j4JcTWvkCK7rzaoJ8Q0SzPHv80Slg6sqPr9
YYnLjtrY1NZx9s91oAl7fNSiVTZzoUvtjwH45wWOkfAw15bkr/tcVO5PYOPL
ptPfsxmDoOhXmmeNZAyXlWEc6O2bafg6ReP6fwHsyolCkPossGcumbtxIuO2
58S8X0HxZYrJokxC/7Xf53/DepQsJ7h/MVTuzD7chMXYO4C06rVeOAR+nWJP
Q+R+cN4kQGzulaw/U/u4X+3k8e+IdxBb0TQtbD5KREEjwhUW656t05y/Bkjj
AyO8a4VYFm/b/MpcQzpqvqOug477tI/v5ryTkI10HxR2lN6ZufnjSkZFtbLl
ytcXFO1Ms6gyO7x+Mi0DsyvLb5NXZqps2fFEMwGfJjI9kVnXWJTyfDCOvBy8
ysE6U0Fu2CCL+nOgki6fsHuCSp/gNYw+VVfXoR0QTKjh3pzBFAURp98qAzzo
VbF7jxLMZC9i0gt/LMaOJVR7garFBLVBUKc/jnPCVg2qb7kfL3NqRmj+rQne
cW12gq6ZXuA4LEVR7BsUz3bA1gStjK1EIFH5azrwQdmBS9CUMjfpfkN6Fb0B
LIidgFfWYSmfpi1roZnkRcPtSPRrDLphKldx7OzV8B2c19C55g7ADtyvESsh
Racmv8Phayt1wi6hzdg3fZFb7iUMh+7rznqYQwybS+zbDFypY3mDG/uV19fk
W4LEYB7aQDugLCX+YxdPCE4lYBU4G9ynZX5uiIPjcqGr2WtFwzDq7cBReD1D
ZXQ1mvhIGxZg64d3qiExcOooVggXkMCHKMTkpoNCVwdgoqk0Crk28WXfqwYs
185LOYs5RzzX3MJRU+v2FR4btPAtljJE/FHYrEzbL7VWjVmQdR7XZMzMKl7s
zUGpyex/sxI1L9MGvd6QCQz95HEs/HxV4+1j4HKnuMotSj3gleAUGxh6vtmp
saCgCedDBzdUkyp8dt/52V8k4Jr/3C1mRLjYOs4D6nfHbmDYbSrTQQibMYLa
hatBwZwuM3IR/MJ2PTyM7XGKQAy02gtJWdHf68fgdmJFitgLnxyehjdAnZpj
4oQAgS7mt1Hf/bI4aHxk9gUK/tLKg8x2LmFvq21yMCWy6lRCbeRYnZf1dwie
6AIHF0yYqSWS0FHVYaw8ozuOwDZocatZN/UxAPU1VQSZCF9WcSFiUtdSLPRt
kuTU6LnZfhj/fgWsfhk5sshxZkoYPjWhOS0orPe2XPU4Xfx10ZEcg2Woc/sD
Aj+FpPeQjclWwaWGGLLycd0PSMRx5x2mtm7DvBV/QoBGcDtcwVEIy2TYHovg
j6Gc5sYUPj5sdVim0F97HZU5JQvonvLi6f+fYaWhCAPZJ4jwBvRGjr5VN7BW
sPtKy5DFyzwHI5ZLjfFm4+kJkYPi/WbY+nBGJ2am21yhr2sRkh1gk9Bt562e
/uMQI+fTJS5Dvpa7JCYPmKIL65b2xjWwa6lNUgaJKH4aXNj5tRs4nV1+0Z6i
A0AX3LBXyQXLRczsuxJwZSSX/zpV2XCRiXm9kHUSttaLtBNG3IfpV1shBc8X
ax+wK9kmrTftroeDIHQD0u7lNZnsx4EeeH/1v9YHnmS4Lru8o9TPzMPPlemY
Cv3iLUVDJqj1jshtYkjYBKHqxf/SNmRKLKtTHg66EhXzjLW+jcvwZL5OEb6f
jeHcU/WQlaPkgR/8xQ9xIEg5bWRz3XSLcfI2v+IuhP/0nZ2ReKjJpSrYY/EJ
d071i9Xitt35PFBhxV5kmzHxn6kLkaoimAHq9eja9yjCdlaanta2UdUa6Gsq
mJIXZbN/rYxVrpExsG445mMbiqf/EZ61T9oG0DzGhUeTEg0a6h9fP94Azavt
zR3sV6z7sCHHjKYDU+3y9GLaxQUNLNkBj0yewZNxiAdy4SwzXmFsXmhhlhpI
F/EeDIH0y29LBBIIGQ804dmIY0Dpmp2Ar2KDy41U84kknzNZntC2U3fGcuhk
rMdZ/UNUEDv/TlW491+U+noepMPE5X9PC6z+tDLl7B0Pe1hqf4PYOUkOtYwk
RQ/mZSC7O1SpbLhuUmKNVNdQM8wGvzSI0TgNTQ/S8KpMs51SLvV0tP0sjjv1
ASkhjOIzOplfScrhNYkYWeLKgyTisS6A5kc5k59PVFJ8TCB9A1EZKpZF4LZA
lAmUZCqfL1nvgrzdFAt/CV5ZuOn4fSX7KdSC0wfaB+WPGoLiIAM15Ap6mNw0
bXKg94Ov6B979on/iALEuWv6sKunJ65JGkeBD+/7d415NYdGvnlhlF4L2WRu
YqGl1hdhEGc7+DMAPvWL5zSLwQ9tooPw6uPJTZS9fht5+kR8S9993uIprJ2m
tZapGaM7+4qVHs6OxAWknNpymh4PwpNoQmnVW0S0A53EtI305cDjPR1cn/Xo
rEcqTVU57CuWqDk3SzXX6PqVXkTc8aV+RfgJLlD9UrDpY/wfB7wZa+wpGNlU
horQ1E/pKJ58eUzsRsMQSfEcKtlFuiZE/E6C8lc6LqOLbJAreQm5TLBys+rs
96uT3zdlVO4p2QOMD8aJE+gxntyrP8jnas5YbyP+nq+D7kpn6FGkRBQHn2wn
lk1NRGsyche75UoQL8Kel5eFzlq98F/y+W/p/BmDX23PXd596zcKh0vmVQMO
7iUsLufiFMY+sC4sFcXQBm8eZIyTdNPWHjamcDsBkrGdVU9953aeMSyFqnjE
jF40zVdCH7T4EW42lpv9zhn146SmLT3ZCuCtORFtD5Sy+TQg5GHl88up15N1
mmuJ3Q0MKyUBsCGzJ59d3yq4kpaOvfxm8DScabLkl9dFuTLVPOd46sb4P/mY
uB4OLEWc8boiKXJl7wBZjJ/tpC+yPebsaf/Qsq1yNomT9YQz7xJCulKXrWvY
elU4DOuDNfRInKocz5jlA3SJJr8EjqXVRGQmzkt9nHlVEQF0kTZXPUpP4aqi
8jcU0AFYfdBC3GOAX51TEHV/7xKWQJInDhpEmf9wqyglFB3HWTp8YNz+GrVR
WbJCWbffJQGfDDrgSosSHh4G1d1o9aLWHrAJxUZb/1jW4/0JIK3QNtFVg9vo
lhNWz9nU0wZTX0X4jU2//YTAMKnnjm3KNjCE8YnXVPanrtebPz5HQQCbvAP7
BPlLqJqQVKxLHn5dOCD+3COkrm7W+SjEPL7/fGUaV7IaPeSetr7w86X2p9xq
CvIWh3CvZZLVYOlibmJ8ppI/7xOLkAe0m+gl4Va7RB0e0+QLbyrqXFe5uBmf
NGlgsYUnO2Zge79THcuzdNAR+J1jCmVRtR1hJdnOYx3zoI6oVur+UGN/lJ+W
/BxHkhplRTgZlJjRp0uDoL1hwUDD0km1bPhEIkaSVXDmpG3nBlBqEDQor9pi
tNzNn2wDmPBNR2mxwTxAcfmtjULOqId82p3Gb3K0WIcsbBwZx8yoCoAY0VwI
v/IIeHPjYvpJjpHDwX37Q2xGaPcG63WmThHVv8yg96ZP6P1umNDr849ZLm5b
C1GQPIoUQMpo3grvuVrlQa/sOwGs9GtEQ9KjqO6WCeM1DfMy1UFbFHNDzDZv
Cl5RqwJjlRgjTR5ShXtKluGduEZXHkwNw6OoUe26bSAhRVtryT4M/Rf1kUnG
pHCLIkp22DiG449oUM9AcLfG8a9LaxkTuxr+XY+mKodoQus9Jlw0J//NVFq5
2TEyTJwmwSPVXbwcchFQclPG8IynOpcB3U7ra3wUfZNFINBrkJ1BJ6fbrMnt
EzCESSjGPRXUomp7o5brkt0ggdfZCmNNWZl2XHajndihVhDVX0GPiAeo+6nf
1saNf4Zp7BT/UTGJJ3cLI8vTHAwrouAOVcEvn99PFCjuOYADcE6YUfCwirbE
QuuXBU7ObETcKUbujbAW3OQPuk6IcJ+UG0WfdqtUwXcCiXTDqHRRVByEbu3/
fICDJS5wR5zDxl9paqPvApxsNcVbLEdSaCNc2/SEDuKvfVKkeTr2Jn+EHbSb
0svGWVdu48BTWmnpLvyDvzDFPTYGOStvJcN0uhDpg0TKj1+PnUmXuZ6t37sG
V7IL/aS9vaawxBfj+7ZvIfQuFRVLikeDy/StAmsv72z06hf2HXw7C/+gnujL
/m4dy34gPsg4Bt1IJN1ynOOiNZajY2lczZrlz7WU+NwI5+043Df8eeqbwZKW
U3t6q0GF7dPp/XM5xRtgxOliJ3X6H5KpkkNvG+GJXe/gDnAy+NnMpLJxksNR
om2x5IP3qgkLpfsy4kApISSlIdVYi9f2o3V6sM54VRlDojLDW7isn8P2hiU3
mLOmqEeSwTsIfN9nbvthZuFkspq1iHm60FC7pPSXUxhdoM9jlIua0DbnFwai
VIY6kqFP1zNzwSs+HzB7tZJVf5/BbmTt4UttqP6D9oj/t0ni115HkdyX4/XT
iUqjcX1ZDHcAxO0dTYoMedROBi4yvQJGzJjmj9BlDcUSxcyN9YmxTHJeggGO
wWPOEkT/tgN7c8O2mEUr52hq31kxvPU8DNPbbx3CvaZJhGy5GfB3VAnpAHr3
g09vFqi0RR83thdOeSGmxmkkxlCNCbfBK7H0WWCz+0TliZK4uL34zqtLOyB3
PqqOsyDFwH2BdAXa6/KNQ9xn97Pl6Z+CdSjVVxSNIJsO7XzLvTQlIu+XMYBH
dyu9TOm4BHcChRYW9rkOjJsdNsKF2X++/gLuYg8uqTMNmyR1OBkg0C6blZHZ
MwxwYSNHVgZfr00ImB234roVG/jG9OIPgZk2kajkir5tBIs7I3mpJ7dwrdy0
IonVQ3W8E3ZqjeQfHTaWLuR2NMFG00iPBUOeqcgBWtu2AgFHLYELntfvpPia
46j4lc/XYrLkX4QM0ZIrjpISSO//EIG8fD5fL1fqMGCsHs2xm69LZtujnxZN
OfNQvU41dynggEJ/O6k6kjcv8rPh+3YXFeVcrWmCDXPRjjjyWXph9O7dCZKC
PIjH2soM4AvikHqJ/E/Rx8jtDErpIeR8kCWKBsvafILTiDaegv2IuC4rRMxh
oq31V3AZ/FQ/dPiZ21vukztMYuB0citgLpUhpg2ZSn8hh4UFfV9Po68Ar08J
e2spRRgJLJM0CC+xOIBwKrj0Z0FStQcFr5qtS/LPXuIpmjyNb6SkvVpiNnLy
keXh6GiWg3Ez2jKLyN9+8VQFMcRR0P7Hl+ZzFgy2v9Dqur/+uz0reta0vrGS
NAFNDpp/sSXYtKdxH8CjTkFOguqBJY1S/Mxm4dMwt95gwJS6S15RKTFdBXYh
28MYCFvoctemrfMRQCc4IFKvQhHoo4aAB6W4YwttnRsKJCH4TGx5ZfCqDjl5
8fazlpbffQ0MKFR7ZA+GUrVkeLzgTBtISqIyFf5ITPGqjtGoV/WQMpH6mecJ
GWGLz9zzeXvsIQkFizws/NgGRSHWehM3O0VI0+I61GSq5Eer5+pmVuoN46it
W075hUhWO0J4zdQdLlzQAv8dsbR8SCnNe1sdmAeYZ/RzjY4fGUsZ4gHWwijM
tifMR889iEspViyWtMqySLPrZuZih3oWHWcB06WWmAILNokQG/gpHDHSeJSl
2hytAqdmC2B2BfyscFJaTOt8BtSInol0eV/ForEqANhUN6vMTS2txgJXuCuI
fTGU7cRevUu8KP7XUscdFBkVmczYP6zL1zs8VlhlXX5FVxTDuP/W+ICFR0KX
xFprOHyi7X1Mif5rG10vleaIpMji8UmcEbi9AoI0NzC1zVvAjAHQIevduvOc
+M3F3CTxBPZgiEQWes6x09D9gueyNuub9XRfopHMwFv7g2Y2lnZOTNvFd9is
1xf66rtcuGePsIs4SWNLQ7/so5w1t5V85ztXn/JJkXDle/DqITocYmTgjenv
Bx3VHz6ZuHNBXI3knsdJFfJve1vwi+mPbCadWC96wbRFB4zNGQXvw7dOWfUg
OW8dPpAcxXnHpGHxvtJwyrjB4WFdJuDUaDJ8OiSrw7sxM6ZAkc+EI0xBvPDR
3JvuNGKRy5URGF1Wlyv1ngBv+6L1KwsRSHk6D3KE7ocjed2KMXPRZdurSySq
RE/MOlDjJok3YgNmQsiSlmO2rH8nwnHvrqJztz7C7rgknX0fsnN1B9FIbi8C
Lf6H5J9eMmkwduRMIX5iqUvI3MHXtZuU45A6ZD8p5bQn5kaio+PZ2q04VPtt
ZwerlcY7Z11klIrDbRnvnSWLjDtau57r/OE46n4hU2fuqpdBmUDlYzZUFpqL
WaHTh3thtIwnlDsRjllQl2g6fX1zzBc5PKAN4l2p0IZlAjlfODn/kWjq1sRd
/B1JJXERL+HZiXvb12ma/T4tCVbFYg8VM6ftMeLcRB+lcnoDRvmN3sMgpCjW
XYAR2M3zgpcDqtL5jXu7InPkSobbWd0IyR2Vh1nXBoP9/fm2lECn6h2zHU0C
BZQmh7J1OStEPJmMCaHsSVyoUHG1TKBiWVE5zJzw4mTJ0JPF91UwOw0cFb7m
MVePct2OiW2XSDiPL8ThddBtHfZuwFBPjOgg62ic6sRvnnLjYz5gdPz+kz+C
jhI2r+hgsVau5NjQLP4bkuPihssrvskmg+vqJ6Z309sPZTZxlXFhmDWrFugM
M/SaVH2vkfE46EW2uo21fKLAZgYj/JFezek8y4IFxsWX8zXEZHLw7rcu2V+a
j0nr0oRBSlu/FJCZ5wcGptLL7SAcx3G86PhGqSpAiKwcnA+DYQ+GHochUSkb
rKU5aH3oxnJubNUg/R0mCJ67JQRsjRm58PSf5XLCiG3j9+5Clt+ezwAh+0wo
zCuLXlmIDPPs0WSTXMlKSgr2gU/UF4sLOHOWbTgRZXsKgHkMA604HSffFvp8
q7QShvUlU6MExbdyFU/280s4ivxxqEluKJAfJTCk2GEk6IBp1+F1WOhVQJsH
CXtS3Lg15SO0IsbPwkpvK2ONCrs8xsi/zksVrbDGcR/go2dy7LrewZyvU5/G
QT3FW2CLwChXP9Cjp7ppq6tmMf5Ex5jTfENAJV2oCcAo61SHa0oKRTNSRIZL
hV1PFejHAnfo3KkNlUyh1WoXdhJOyI6AOsmooAv4grnOpb5QFy9ssOtoa0Te
RUIahXdazpiN3VkgD1WWcpydQ+WvE9t7MCOFvQfQfh7qzunSalMxa9H8pj59
S3zHMygeP8qKx92MWHxWhomlMSWkoNKqm31oPMSHym4/lfuAh1H6S9RoLCbm
VsntuSjyyLhf9Be+A7ch/gJAEl9ddTHcr/sLcFW/cz6GOsRni7etW8A7izUv
j5joNdEDLrWfUoRZlUlKprfzCuvc5ufO2yCA4FOwoATF5Ioz3LYINjxR7Gvx
UC1FOM+f0T28BRvB6u/FvIOBaccHEF14B2yxT3ZTSgC060WGhFNl8Z+Tltya
W88Xq8uSweyGDhA8DfS8bilJl1lgUHkoiQykObDjrxdlUvPo5S96QX33lAWK
fu8SFnK8phjgRlOLnLBzsQnZdnbpYHtrJToT6DyfUDZ4DhlfUzZiSysXwpRZ
kM4cbzf/xxlyEdH6jdpToY1FTqcEVwEIfv8XujoOAgeUTY9s+YK6KK7Vt/NL
Fg/rQfBGtTpSkuxgSLQf67dKiAftmDs6uz2p6QyqwMahIlFvmhBXGZZZAGor
2DCQZ5QgBbCeVTieLWWvlZ2fKAIAfiRmTAk1zQbWXHBLQ3C9kIJ8fETeewg3
+pdZfJgf2L06/pFp+Qzc51PXqH7aCEqhc1+IZysRpuAcjIH2lipJW/jA/d2Z
6b5xJVuWsy9rAIVToSeh0+TieUy6ZpkPhNn2GNuwcY4SkNP0Ei78C1UADa0R
0CiLe6m2Is4ii1xJ5Kb2W1SuDJsbztIarK3KIc8rrUWRWBNdn4NGcvIbv8Jj
5jO1ajjVfXlrj2bLyWnjHnnCIaHmUmoCSezKvLEO5tyFtNGLHZ/R5mmLZhot
bYRcz3S7xsdQUKOexg9FKZlSohhTLMkY1m9rK0mnpKyfXLsv1jIsFNcxiQ2m
Uwxdq+gHFFcslSf6XdkHZQdo9/LJnWXe3/QHpxzwkYLWEGumoSCgYFT1bfrB
szEgDqRiz7G4HlQfY5VPrP7FGtmn4BVSOSjw1F7vDNXEL7KzCvVsgVkZk0tX
e2+/qNNgE+/d0D6S3cB0KiC703MYXzJE58hxuP5MEhd9kVMljUaqJ7sFx6E6
JAanBfsM1ISXfyGHWyBnwGaD4KY0Ugif+RPfy/Jr1TZq/roytKnMB0CUHHbE
yBfxp3ou4HrHIw1UlFRyAEayStM+9moZvxZg8UPyoZihPWL94rCZV9ct9NHK
OUurSv4g6SxT3CcGZidSA1ZNUZl5UgjlXmE7DK1WirccU33/lFwNRShBvM61
ZVjfRaDhNLWG8+CAUjtn+PaUzZNkLxpbWvBsjVCVNWQfILyypAiMXOnXL0QC
JWXUNfi8fzBlMXFjSsxWBTJZf4iab6U75M4q8OQeWqKb1t7DbAVDkaZ7T30k
uwtOEca5GdeJJeX2WxPz8CrKPjPp3bFKTv2MZHBdeXz7RFVqqzo+UeIeL5L0
SKeuD7CF1Mmi3AFQHlwVAKAJT1TqeagvmHGoF1F2fUoi8/jy+5d0ZbzTNcci
8ZwO3Q+6KT7DMi3DuPasVLtvOBjSlHd5xCGpNB2m3yOTq/Gn1Ly4N8vQH1ru
AjHzyFICOIT8arloUI2xohfipxQud9kIYeNUOK7bNTv83RalOP8sHmVvC2+f
FRsCVeb9QLuiDvRFy44+OYS2g56YLiIFL5keGoExz0dOJ82JGIfzOU8RKQG+
hN7h1Y4tr5GqipdAH8o5QMiYBqV+F6ATLGU3H3kFhLFI0WP3BPn24OilqlW8
Hahi0QTlGQu9MJMQCX8zX4X8p2Lweq/GLepV8vP0zeiDW1PgDrxn5hhqYmxp
25CioNaHcKkD7ZToT3ETKMP/v3KBCp2Nqd0TH2ftCLcMfRUNJpORl35bMIGw
IAFaYetqre6T+MqgpGvHz7vAeinhpPlo1yqnJLAkVN5s4vMFvHbvq4JylCyc
7tWRF8iVnlbkVD9D1a0PtZuwADbFdLKs3Nk10zQsEX35wQCsfoE9Elzujtfx
Yz8EavOlJ32YQzbIi4xkEIbG7UOD7tYhcUuh66xNJWYOJ3QffXxGbKN/WFUa
RXY7OEJwzDO/oCxjJEyE+4NLtWabhFNSNSF7hX9K4a9ze4SVI25pVlhD+AY3
qEh/7GBAzcO74nBCVsfY/CGgCNW2joIXpjd6HYtGRPfMLbsAfLiYm6lSeTNk
KGG35rRQkpscSBvs1U1a95TFUWOWZcTbT3jzz0Gvifvkz4ZN3+BY5lZrtN/M
5dvmxfsdSjB9tIYlizMwLOd/zq734KCgDzmkkiO9LrvkkFP34XWSoQB8q3E3
wGGzSChp/fYtR16CZkwdVZVx8tqrdgEKBvdHytzXj7sXmGEqANb4JJpMpFba
if5PbMGhj5Xz/dCOAZ8oLr5qF+LiKHV++gMEWL40sdBlZ2MImTWLtU1ZhJqp
oBMf3J71u4Hcbn8AQZIHPosMyhURqeTFduTNrlYVu8hF0YcWWTbdfS9ZIa4Z
H/6XDKcAiqJlfPtOkl1AAvlMFkanABDLLnu1WtJShzQv6Gc/3tTcReZzEde7
rUdcXy4UVTi42TG+eiKg3BNmwEN3DWIx+Jyc7CkB8sR5sVUH9hXxxNsXKqyd
2Yl+baT++Mzrp1PnOiYVbZV/KJ2owsF/Bu46hLaHc8cgGXmLAnczCuQ9jPiu
ay6VVJz+LtIKSohz2LX5F+IjvMcvaravRg60u1ZHxohENlepBAQ4ypNgTPSK
USo/DgnGn4FyA1ercRPUiQl+ljbozYQEXPWVMuQwKlsOT81qqHv+8WjDc/cX
eQssxXN97XvNxhWrWFuCGZwkk6sT2gMReAtNDxRJTU6+jOCBZWhXL5g6F4G1
PLOtUc6rt5igkmXpEL2zMpEZkZt3CjAB1T+GlXbQj3oNW1NvN+NuUv0RVjxW
+N8mDPHjMuaE9omWOtfZZXbjWSktOzdkcAh6rQv5WukP9tvjZyy5Xzm+MM69
Ht0OSOSC7++uExJsNgI3ttbf2dIYgMTvaGfVySQK/vsmetbrqZOphRfjNfLc
Y5XTd6v+kFoTnTQ17e9k9+ML76M0OoGtuOBQG/Hj2Zvm7FQmoYtB25eMgYJa
K4NZeXsk/Z16NIQEaTfx6UnswF+mxQWkYraoEZRWtHBFxr9shPVUv+8c6vLC
QhBunBe+tBR06FFLl/E6fI8fgSTevjZanVXupbBMVkszOGgRkimL4eneH1T1
z9XCDA278vYOggpf2yHs6cvF6tKLXGAsDGDTfGu9M1831r+eX0pzzteZSBJc
g/T9IjDetMfc2ywEghIn3zwf8ORX+IIJiJNdzClnmxgzrrK6F4bQQz4xsE++
9cAoUuuPRQcxubnbfL/oa/a0ywqjcOYaNVrcBiEb35O44zGp4hHmCOAmYHqj
5Ji5fgU4d2HL6jKFq88ud13MU5zncRl7WOl3fjeEIbiDhtp95KjTkQIA4CO6
VGEgsjmIyzBp3jZq41Qbbt0c86q65OogvWFiKZ02i5oeGeWtjscw3W/7A9DW
jHB+ZuVMDYZGZ2+pefKewGyCuSGnIJZJgKb9gCI+7CKviJMCG76S5nsjFmpH
SeZ0Jhr31U9puZGpwNsJfAPRBzpA9Xp/PQpGo7tuzxbA0IqOczJdQQNlajkf
zhb/sTxL9+3U6r+01WQRqcWosZkQ+ray+u03+2jf3VbsGAQM8omnTarjaH+3
xBIOR91E5WuvrhdETQp0J8ZlV+QjmlORWCtrl8C+q7KpLAsi50MDrNQom/M0
82Qb0ObcwRY5nBxOvqgm+UZO0eGW6WMJvjFD5rJsgifeDpSMG8QDxVXVNsSX
1aa8mIe/Y9dFsH2Il6vygMU6kwGl3aW4Rqta3+b0eRnSi/OvgIDzevBLH7v0
6aQzqqTKyV6Y/IhxuS0KSmLd8Ef1W5lQFjkO0RzXb7xduhEwLqPMCyK0MZFO
wbWEBeBGziyQ5MCc85IPHsouV5KaX+VYggX64QqErwIFmjPpFoqLebibpTDo
+Lu+u45dFHJHuwBtxzW9wAV11GdkodAwHOxgQRkpF7kkLoXnvrvkIffIukcq
0FYG5kARWnLRJ07esQOZ399K71zeTIzoaEnP7H5o3Yxyn5SyJnYpqCKq31zR
7lcGIO+4eqmQbvHwCd8MR32EI7bSmBcsgqQlR4DAnzn51bTGthfQT/lbMBl4
SN5Vj//wSFTMrs/fqlO1XZDuut/YYDtCCDylimhF8iErbH+05xFc+N6W3Xy9
7QAoE68x773I3oYGDySHkw8EveGdN5Sv8IAZ3Nucb5yhhgkqHvCIPSBDNNI5
QX51dsojir0uy9vMznAGWmec39UiWIJNUp0wgy3vUl4ryoEAVqnyetZSBs7T
zcr8zO4Otil/FPncqYkXEiP2jpBG9hslN6mt4vEPv5rcRpZrPiB7D01OMm+i
Ypm7rx/dnhuLvqZ8jHpdUJsYmqXtYaVAEqM/KPc3z/NGIxzLweOslt1XGcFZ
AKAF+eoERMdLMqK26dISSktDJf2plsH8fjlU276rQit3sa5PxZ/+MlYFP2X4
RVBkGvRm4Sr6Lip+FOnD5EwkfwuaXCJJqvprbZa/KON8V8HelXfNvLlDXRBh
AbJXE0wQ+hjtVQTqqQaqxRqb+U6tbJRt1N4ft7S2DKs4hrEu9H4yYajKNENO
JUFYR66tFVg8n/BaOtGghMwxsekeVQo5V3rO0SsY5EgzYk8dY3BHLDE5rz2M
Gahe+s37nfBAOA2p/TtX1FnmxTDE+vcyqQJmJFXLl2IE+QE3WiATLrD2/rDQ
abnUs0r25CTYKYtrVxhNTEsX3mJXPr3IcjSOtZMvXABSoqITHm5y7kRe6ttu
vkBKxWHJvQZ2hcjEUWrd8MmdC8DUoYGQYVHIliRBLYHclMVFwxh834+bPkkI
B8qYL5LfKMo+jawTNHtqelKMlkwP/bQjm8NuxlLZyegoIc20xicDyyBO6k2K
mEf7swtH6tgO3OFPhvadOa6SW0uGm3Q/1YXzq6uv8ocfjkP9dqeSNaVH2lE5
KC0z82X2f9FUcEQERL3agyLP1Qrl4C9Ig5iKkTbIAJxcmnTbJy6jEv5LA1QU
aT0JJvI8hOoSZQKhruABFf0PFRjqieI8no1D/uQRousZg2iS9ui+EfHtrmAZ
pbWTYpHOWSOVBlUPh8jA4gIrfKkbrqMl7aIAbjOK2+RTAtG5owV8BcIwUlGG
HuYLgkn6/fMx9HVzGnp9lKjOAMj5RZyQ7cdAPHfsTfgLxWn02BHWBrEGAtlO
QY47rVB34bGBuwyTPoAXjO0qppsTvhDW2Hg4PggX3y/ul8PnnCjQrNhXOdbu
FgHLh/3u6DkCJ9T1YxtVDTLQxHJzHbaDJlnOfB64vM7LfcQ3FxcvSK//NND7
3Tb95yENgqDPUQ3zW4bS0j2JNmh6UFF80yZMXla/55Twikb9OaViFlvVjPdy
8o7MHaxTjqjUX03SsKL3vmM2JEn5g69kpMGkaVsCKRv1+wawmo1y0Ymu9AY6
ug21NPN4KE71PS7vx0bmDu9SjB1uQZb+AYiRZYu1Bcoj6YAXVFDo/viNY9jk
v4szzcX1dqwlbUX2ce+Ve60ArbO3CFFs1Oub2N9hOtJSW9AZixpjCXaXBSjP
2a8NjS/CzHyTNI5hQD+SvHmwqsOv3sIhZ6s8nLQE66tN0dpnGnyShg21tqCa
gxLZGlx9aTkfNdiOLkD2B4vB25KVUW6sfFGvFgl/Fwki7hsvHy1LpQwnOdRw
iB2pZj0+ARGUyDCoLeRG20dArcB/vphdVwhv0FN6LgnqIQzihf9YpsOTw2y4
2GTH3uY9oZerT87wC/xUkly2aRGmGkkcXqFwyS2dDilFNop1zgyE1uejbEnx
N6p2QCkaVJjDojCEnVYJGWpIhEetzwJfaCRC90iHlrOaEH1ivIyqVCMp0Ivo
kFIPdQcWj2q5kBa27EhgRmEtDaLEaSsDNLfIAyIUzl/86Empd6BGsaiIN09S
0/E51nneUajpNngxUsDuM7G6MbBN6Zb5P3sT9goUcrryA2t+rlillhAeWbq8
BALoIdtVkuXk1/4MR3s60bW3IplgJQgMvAgihK4nAUiXi9J7hpCsFsUD8DmI
6pGwyDioR/Z3jCVhLXedaZDifSqWfPlEtMipp3Cp6DMkBkAN+XYJZhhPzT4c
aiKm84Mx2fdDgNsTn5APeIRVy5GILWNBOPw6buvMsrIQdmvyo9RxnWhuVqGf
LG7NRHZMPQHAZvmd5/bBiUtNCJ+tsVdRn4ObqW8U526JPf+jEpAY9KWxdlB9
kDRXkah1yMFQbdamtdWMZTXvSUQKM3C3JWxb4d1djdDVV14wm0fZWfk0CWuT
6FVbEAGLCDl+WmVZzvfSKZprNOFpOvP6X4MTV+LCHAM1Xq6b8urdTpj+jhPv
kIJFcp+fXL/D0ltLofC9v8PiUgWFMREQYY6lTxYdydQ16KLoTyOWAzh4wnSb
R0q/Js3g+Rz27Hap4wg2jlUtXnnWFj0uqAkbGX1H8DI4KEhpO2Muubnh8RXJ
ny5uI/S7SkLhIQePQZayjUar/2gbynNkatojf3+OKQbUyb6WOSbY4N6Gjbgo
/yBHxzAf5RdH76DF4UNu9YmbkCljbEFgVm3cHAKzgR9nY/1Dr+EOHLtiucXm
JCWsDqcASSMe9gljeD/dKhHYHFNYPwfNM3Zp319keKAW4htibeAy5oBgAcQB
CX9wAV2+WCpc1kaXIGvCb78cr5qcjKw/vZa2JsIMaO8l6e7wiWyRAAIh3ISZ
vyRzFvdXfNFAR9LtOh24Xwgx1oPyr48jV+0eNE3mMozwKuvwQKOArTkne+oO
reGgCJw3Nkjh+Yf9uw/yS3V4skH+1339P3R8A5a0naE2RMBy8JE9yHk6z2sd
OwyiwzPuX8cxZkDrCYuYCeZUzI4RjpU8FcWfld/VnMffsriOpUGSKuCYAP1b
5L7OAAPVrIK05AhekfBiTEdzeQq7yj0/zeNT4msOnv4e0W9S0VpWGmSEMIr0
sz8XG3hIeqV9Rny1J6zZClqPaFqwfTyeVCZvdacsuE5DySJtkYicwqAYmYGO
v7BHqqY1OtXxdGcT3Z5CntVNxGwCVY7Y6VREPet/AZyI1197MvahJyEGMeB0
dfF/8FjqZ3Dkxlmu7x/oXXX/J6M2hMyFojc1StSGBInYzL5lQy1UAmk4qftN
3kHt+WUOTNF0tTAoafFjsLAjfH5CRhonZluBu/lz4v+UtQo+8DxpR/e1bqsq
fjOLn5ghgcbIkRRqPPE4wXAxC1ceq1y7FXAlnTzCuaggoe/iNaOQAF01vUCG
E12A5cztOUUnqu7ATOIiPFpovoIIh22Gstzw0HjhIDOZh7lFpRqd9r8R3Gta
5kY3DcnA3+nyy2DZQgGf+1nI+IOuJzGNslOgA3O0WNa6kiaeHlEMmyL+HJer
Wacsb/O4Lz3+HFAjhr8qOGaSkB1Xb1XWyZWt//qFg3KjpyN4YWLc/urmk2Y4
0wSCHvN6iG4LsNGLLsnXQyvNo9ouvmYQX9ob5YBNF4YvzyTM0Qmub4NA6N49
+B5fskI7r6raKcTWnKXl9PRN8XvdFQXBYwENIa3VFBlOPpAC12WLsIXEbufm
r7gZfEPKDMwSJR70FrJnrpO0w42qPqL28Jhs9wuV2UzaW03Nyu+rbkI0JGhd
QTbpi5xxY6mfLLh0HI3NfxP5/cUs4sx0FyJzMvRAsbvR209xYcAx/GkOXKC2
BgfXj1Y4sRe4J7KcSts3KC15mS+Zt/3RkhBxXSjcLPQfjPjo050m94OQt0Dx
7qjCgZL6yEJKv1Xz38iDnqTE28eKCvxJ5mCAiLQB0YlhB8FBbdCFdW0L2/SV
mBNnTCI05C6JmMoCNr6ODK1rRmcuC/otvXO3QA/3EwxKKzaqyC0gYXnkl400
tkVLcF2++ZkibJQcyuPBpGCSHb+pFNkhhH84gDS1Ie4duUGoRbEGEdo/2V2j
/2yWtOYUgm5pRFM1JELE4K3l6dD1cH2H+SAs1eeLxFlAYeJQBPf5BOkBqwyc
rTuJXO4YqbSGRk2rcI9gdmV5DLffc39rM/QjS1liZlIvIRSpkmGne3yhNetJ
+Glzf6CnID+DmijlRHZWPMGi5oxHB9aSc9CZ/7Q2nFVWgee+dM60tuBQAW3C
Ru8NHGhyiKhLpnsOZG7mvb697sJKqtpiDKMG5SjrkKs+eIkO1rzV6C5GCPBX
LwPTOummjebE55tI+o3XQvICQIki5XSZvn4VJx36Xs6M9owBuiAFzC/sPhsZ
8tW003uyjyLz4P3c0InzOTEgP9uQAmOUoXJdr/4HnFiwsab4aJoN05UJUa+S
QNC0f1BXOWfHKR4JAJlPlXgK/TZRcE1VkqomKWNsGiIsyEVOM2Ydw2mi+1Bg
34WB8IOA21/mj2wRM6nnjY6nLKtGSh1gP/lUEYyCsOexxb0bKja5TK/O26LV
irXQd4pjzGYbh1tBoZxP8e53ZEz8ltPKmuRuOFvVsrbwk0kIkExO0N8kXX+u
hEFjZ7ae/VZk8ji/NYEz1oTrWQKzmSdyhM1lcCNAQubjahxXFCubEhmbS21h
Usu/PnAZlXg1Y4YFVIr/EZnZpUzX6mGxxFCuPGTPaMA3NApKvdxUJTc3ngCM
DmQSqK7V9D1ApGvb4wdd2Jsqpe1Om7k37AdAAarw2NWROo/CWteEDULGBxs0
6HM5GPqb91IYU4qXiGeges+nytwMXC5bar/5UH1cRjVYDIwc4L+1oC0dGSdb
RQGP2dMxQYOkKy16riUm4uaBednZvkK9N6IprmTz0NVbWK4cN0ElHImJcaox
W0FDNnLxsfa/jrX7k0iRfME625xvIiFaB4PPHToIJpGMLzvyJlIqn5kI6Hhv
Yeyo4ptv/RPTVZxMvZkU6/fhwvxIO2jopsgkVsXhQonLPlIUuPpfPg/YmHBS
zATPa4x/f1FlJGuXUADn42cbt6CYEFcmRJqmLWo7DVh6VJiVuwbm9tHKTLwx
Vh8xcGrY6VVbDEmTan2VBrmcR0d+4ToHrRmA2vNgLgKiYdo0Ox6El5UGRHze
NwnDtUeB+/zrl6ZvdjLoTTKUmJsozT5RL6NF9FXKY8uqsCWep2qsdYLX9Izw
AFJaJ01uzoOPMsCBE8kQmhze7nhQ6oHwOXrA+xFhOor/MhKPzdkAVbW4g6sn
Zw0H3zM2mIGW2KerQt0Y5cZGzwFhvZv9uhXB7UaQRk9vxLttA8h2Sdn9XB2A
LZY/9og9b+S1+IWNj4D0qEn3DGdwZdm7uqW1UMdZ85fnlKnonyYABrCF0Chu
baDWHXnRaQoJnqSH4auG6dp5vmG2QNFaQmMalsZKXxUIaqoSdeVYDs72L8Mt
pURkCcibu0WEWiQ6+35U8rT5P2V5mDB63G8+3+NgdhGiI2zx3segzkMUEmFO
rUBWD8Qk7V/CG+uoIi5MTHzDCQpjfhuWzGwzx7XOS33MAOxaW1/wihnZrQOX
nJyo6gnh48jP12/nAl0iAisE9/sYoVUakBDVInMUacpvpKxGt/tg1UhZkzxr
6WoAwLG7XGfKRNOXi0ZYzreLS1f4vUadtP3nMv3PWJyfkcNybLOHfo8eg6k2
2pJfncvJZqqtxNHDXDk3ULiwS9eC2WK8qkDp6Im2q2HzjMj1OKspqdQ6UE7y
qVEuyMxX85tThBvwZ25KaBSw5/3wkqgzgZh+wVTQurMGuQxdqi/IsOTUcPo6
34zzscbacjVDpJTk/O4FkLOxyK9WRPRDB4IBN7o4B2r5HicaeQU+PC3p+mU+
i3oplNTJAif/MAI1DUTBGkBxPz3L6kwUtx9oiKPcpFcp+cfthWtQXMHGKZVd
WUnIgKgVYUpvfX+ksRAr4pas/1x6AX0cWqx+qZDoCKJuxc1hFcTdAbIxuLXi
GZ6sDe3jnpulWvTZdJ9wW/tyAZ3K4LaI+c8HaCrbzTkArh68JBxQJTkq5Fis
N+P6jMxz10sn26pOS5+lAZ33zbBf6AcbFMC7B7dq/LZpLXBgn3MBNrAcSLo+
Rr/EAyYP11BM0amttBYHmfOefRJP47C5XcptjUNR2Snw29wZXRdQPvQxLUpB
psPT5+/0L0RBQACj3bldV9hyjzC3cF4R8Ja27F8CfpyRatSuB7jvZerCXFGb
PQhZ3Mm6rVYKhMVjtAkkDllREuxOuKtyhwbJx4i7T8S2vXht/wmMYuFXwTAa
DGeM1u9xZPlmCS9YPC9tlFamML9XkCHt20xWWYSROab5PcL05IXx4eKAaoPO
4U2uL5l4KxdItRj5V0gTIzkbSLYSoiG/iehlIIzlLc2WnoJrjdLpxdrgXtFJ
ZS5QjPLGzgPfPwcgXFk1EWcXjb8Ebdhldg0rzjwrxFob9eIMKEUBpAR3IwDM
RJ/AVjpUtfjsjTeDLWUsWHqBOtp+sL/x6TLa9KzQHyriGUDfPwUOH2HpZjAB
efOG71Sof2VQDhq2lZXzSi1RFOwpdu0GzOyLq1fuAAGE8rOZpzVO87lMhbUD
1veafq5TSVitI93RR14rMQAJQH2LPaX40+g9Cy/uGqvnly/Lvd9hMKC4RPP+
mteVTRpwh6NcUVZTxZ9wpmCGzbNWb8BwCh896J5VrrUZodWRnd6AyCwK97D2
aWJC5kUZTND6Sn0GnPpdg1PPE1yG26hlJnGN3A80u5wfmLhMlBhF+7fiWOWZ
rSNxc0lDggBHLBr6U+yorFc1xCfmT+KilFYRHVStIjJ8Ql3bXkMo8ljug4lh
F1uWWnDkU4bMP+EtUP82HlWM6/vIZwSknkzLz5oylJflfQZRAywUtdk8n+yA
foGIlt5eWrCG6gjqb/xfWTdT/x4GZfnYQRYPIby6Ot7TchxfzuoqMSmYyM6X
i+M6DixBE91Z6nPpDGBZCzUYwRSRRJ+kmL7b/KIZst/mlborrJSyjXG3jWUl
FphUBwdF2FljkBcPPfgDsxeEhLCGRPi/hEiB9xmWPsnZpm70PcFBQfli/6H0
vz/ZGmtwfXiq1L2WjEKm0WaiNhbq1ha17xCS5DhvYMZv2SA57CIwf/Cg553p
SnQ6eonbfjgsQEAtKIfjg1zjFrC5jsjBVd87q20Z3be3fxMD8ragMdo0iDcZ
69IYqOrXMpKCOEkrXQNiqFB6irtOTabK/VAr6kNJifOvDFVB8Hk9O67qwLSg
wFM6vXVy8gzuInk1j8iMYz2GQAqnHAvrju3lfdN5Nb4oHZ0NbcviubmZ4Vlg
wyJHKE1UL8+h8qr2CgsJaaz14GaMfzAY1NCwMqXsScAcFrwM3EzvxqwEupXE
6EmjyuGPUvn7R1cgsTN0YJ/lfdMQDM6eP6QtQ4jbndRXK5433d9XxRExIpED
62LD2m4YsbIvwIUk60LWYbs+NkOGtbt1we1jf9AoeMtVfMlZvuHFXelVAFuL
jRj3jo4tP7PU7kuWhWdJjjbGj07YFDMo71uWcG1erU3mDmP2qvj1zjQdukLG
ZtkbXmbRSJOPSrK1Ad+LRDp1g29v8WLIOfwjAve3NnZ4VReGiGCCcacJyTUY
IVIjqQS458pUT+U6zovJTlDXR7nJhvCPvDdwX2rZmv6RRmMuE2PRWxv8rSYw
gJnw5uKTLJ7pyf6Hr40XnBKtub1Lzft+ZBGMIvsRz4BdBLBxZWBVQYoViY0O
YuJsrPoM2sIQUcMoKtqmuAWiYzbbtSXtjeILUC2FaiAvQFEUwEsdQcgcDjmE
mfxhsfYoAcZa40aK69kkn3hack0EuVojUh6NwEqnlpSfTieB09Od9Nv7KIXj
nFfAliSdOeZ1yu95vqt86xqKQBIUlgtLJ/AtE0VZAFsF9t0LLm1eKG3ALL3t
1JW0HcvsyS0gngw0jKMHOYOlwpJFTcxIYMocuB7DoGkqUEFw/AVaCQbbXsCP
1RBihGDHNKMZ0AgR2Or28matqAL8tCa2ToPl87gDw2uJXI0O3foBK/KE1B05
4ET8xlE0NpORHob/F3F+oENEpGYpC7b4sx6FAtZBlgNMps+0v+kC5EU3TMfI
K5ppiY07rJVejFTAbP9MIXcnPpieTdaq39/OcCgl4mRhE/3ArJYNkZ4y74ho
6K57TEsxGnL2bDVh2ekEJMwG+NNBG1slgZpH1CRGx28EJyQXqmD3TC6vh+qC
jmoD4emGGtjwP/YQxqxZsMHm/Ru4YJI0F5uUjhTjzQzCvgcRBZHF/JqoKH2u
LIuwt5dA4PSPHpQ65KgRR+quk1nm5U7rtFWZBISRwxl0FAF5E4Dz9xEf4JoS
i5ABT8QmOcmgTsYRY9bEN2t4wsZVpen1czdKrbaJjU6c1U//YEVG3SOiumyC
mJpb2WYjnqHKZLCRFlzH5CpfdBQYk5niGW345IH9diicfrNuhCRuxmbyYkV8
jHTZnCmns9qSOm9Aozh3XZ+abc/wTlYyHzmE/JQ/Ex4hVFszbf6R2wwZoGB9
pJHsHu6Y6rTqbArWtJ+EXb5XVNbdj1iy+fP0pdPsN3HuwpDDyM9mcY9WmSob
nCrW6uE4DVeusx/JnMXsgbJTnH5J3+QY2L+ytrObsbGuJx09XqiuS+ikpcou
/tpFizX+TcCaQF1tfr99FMK6vA0SU3mlcCTMXYqozEvCRc97z6690qcWdrLe
GG4rV7hLvTbvkmQVcy8wCxrzp/g4ZBiyfLacYrsbpGcsFe2kouMQk504S5la
2YUa/l5+/zOACygwpGAzYydaZBpq2NanLpRA+YqKq4ojB4L/cv53B1A1t+QX
SoWM0vgp4Odxs8Jj6BS6twUrhuiSuYUG7dT3pvb4mAfKwRmiNH1Y58ckJud/
rcLN+NCtFBlxy0ImoWg10r5P1A8BZ4lDpFtdVAdoIS7w3fN3gPYhKt6lHSOo
YO+SkiKbVG44B8/LK7mfDQSDbkQyY0IjQBqterg3XgpEDpbjVFZkfDs7pNIQ
FIINHIzkaloakfkuTtJEgEfJrAeIeS0XakAB9mKPz7/RhmzWNoxnmZad+9L8
ZXwqYRiZYxYkYt++TEBJDWeXm7hpjtfkB6PvL9ErdTGWQx7oy8Cf7eFMg2eh
qXMdkj4Tj6Y0PRyn73vAIuIdedX38mngIU1DXKf9QUUK3BcaNA7dOku/sJ8L
rj3I50pKNQYRQjj9hlbhhtVyDYJ7z6vQ6qvAT6Tm1N7dF/ZTShmDl0SMlO4m
i9PhmuK9OJH+znoJOkhCNVpS47MvvNgrY5I/uxThl6cHugqoUoEfIt26hgcu
ZKslZ36kHZ/GSxnQeIknd8JgsNc9wh1HwWvs2snZvUlwtIjbCiddW5xBLCFE
x+g8YP/12v8m45euSv7PQdqdpv6xsjvFb08GgLAmtCKMwVJiiS6QwmUMx3T+
l8/RUk6pTJgfaSF306iUrPiUff+hAFjqiiiRLBHpnUWuihGkdogw2CqY/wI1
YZ30QiFrSus5IouIvUJzr6+2sN9OSRNN8B7qPqQxn5Y43glZDcRb4yao1Ysc
PAz55rIcaVNdJxeZknPIeh035e1Toys5WFgwa15p05tFoWaIKq4iiryRAKJ3
dsQkZVM5FOXgT3NGZQm/BJNYy2bg10uKRAl2aSZH+nplBVNrPH0q/BfzqXs6
lDCJdY7imhSEPWZxJt7224Aikf+XfCCMqO4+TnGs6LpFAWErkCjabT6cNn7m
VVUd0wEEquO1ZoHciw/xSEzrt1VpiaIyCVWvGFcjsy3jUkW2pKykbj8sMZ+p
uSIjIco96Hkux+U8o4q21RfSaPgemY4QaLFxTLyUpvIaTI7q4G02RLN6QmGt
/yANbnO3/nqXA0gJ/gOkHo9YpnxoDvhU+CrRU/PRxhFRpthc3g+345PbTd2W
jRQbHTsmlBp0H3HJnUp1w0Eoqy4ncV/neoC4jwdhZvD6i7NvmdgwRV875CC1
BJNhWUaKAJmqLRDNQasPB3Hlu7YvtRhDo4nv2dWRxkrdms+YRUtMkEyls3iV
K+vxfz1H0vkz+yfzoalh3Cl6aLwiwqImYLBvtn8SC2N888KZtt3Mm/izuaLc
af+ECzsLtCvGRqsIRakjaSxwt8MzQ1anKbNOfsPmclFQzMyBuxr3r74p5+Mu
k+t1VMqoemAHSaxonFfNS6KuZzVKMi9BxdNbv3CGi1U1RyhZUwu685Dit43g
/whqVzZ8AlcilrNDMGoQrrsyd2KoJB8G9Ft2iMIgY5bcLQt5CkQFMpUXPr/E
Dbiwu2FWQmd63/5HXVyJ+IACUG7uquP68DhrSWPViUk4c0hLtwdfifcu0vjF
cJTc+QUCqF/v1Sk8MoTUMwOajXUL4R4xtD/fqOdZQ7JMgewhKdyDlUo2PBlE
ZiU/RDU+SOT/E1qu6ciL1VC6ykzcgRMbMrxTaZAiSAR1PUOa6wnps7wNdsnf
FqDWrn8GBVbInD25p7hV2I8G555tAr9fCgrqdygT2stbYYNftIxQWj6PxvTA
MZstZcWAYWAcMK1VGboAAKUQ7rNNpVF9cutYSbLsvxvrJzLw50Q8ux6LEKLp
xdv+ex7WZ42aay/syV86AQ1LnQZeE7M8A3DIu03TVE3m1IdiERhI6UsEPn+4
6przcSEmttKfd9rOEACiNpZUPmeLwp2zEDbYvMeP9aVbi3AozHKU/2fAIth2
LToIL6jOtqo9bq8mpPDs6fu56LY122SDgnkKYlWzEPiWkBgQtag30frtvYGq
jJMbRu+85I+JRbrhlfa0wEEB/6GRkjpbIi1RHRsHgD6iVdTtS+AumR0rc74A
12ccFyT+Nvb5035D0ZE5Ye0RcgBBYlxOzrGyADH3TO3LFLFKUK+PApya3IvY
JEEE7dd7BwIMJueEOcBS5j4M2FHm3XmnMdw0j7uvmAZ9tz5uA6Aq9JKW8zeK
EffRi5it0EPEjnUJJGqAFFz3nuoqp2YZtBYa2RXkA4y7BMh7hZpqK00bKDV5
MKEb055BOi53RNSzYhoDjQWtTVybOESCRUmRoOkWanb+800tC/PWsWewM3To
cZqcQXW2Q5RzTfWqpHraASNeYNYxJYJCermrie9sEl4rsBCZ4vfMP1dQKilu
DGsBz63Zx1esuCKQuMZFztjSeaNAJZFmLxxRRWcvbrf7+3494Zpe8LkAv3p0
cFDzN74gkWFnXFdiW7y9sl3+IP710QiF1Dm9lsQ+k3qzIOK8P78Z6uBk/PFr
nN3/Lv9V975B5Q+goFFEEUFiMR5/nMXAaBwpgmnfbgt1aXokcnT2ve/ZJbFB
sLV5+VdLKwfnQr1wkHKPzVHJ+xHr0D3rPQwZ5UgZewAE1i8ryS6L7Za9gpbF
CzVXScaYiwKcMwEM7ud0Fq/Kc0BQ74rtktfeF5MNHVCyEsCsITDzdz6hGhOg
7UsvXwSuDKPXccBLTGKuQVD60xBh+3GeKqRIWcMwb7ruQjgr7EWj37k3qGdB
vFbgp97LVVmG5FxhVwzr8cooUeR53npC0sb2lsH+oRiRgB3aaBUZvTCgmzQq
IKocA32NgM8q3n96KFSHOurCIGxdwI9GSZFeISZXM92mcdynWVBjojIID4qB
tyGbT96xoYt1JW3FlGdwQ5gUEvbUsEAR25FD9xuS00iu7I0I5kv/zqOGatTr
RKJ+mi9PnBltJO6dEXfPt5fRNMYeaRngvzxoPFiFWqNjvbLRfiQjDhCnyshd
TPInszjcsPjfSaeSPTD2Dj39bJ67ZTRJCHnD5m8MsmJ9m7NZTqsUg5Ew9jUX
Nd0fdsNWyxnPX3P1uTSnr6lHNTvjjEH0IjeoHMhW9fHfJmKWnihSUQWQH29N
lk9l3xiQ2qY+rB3+35SJOIJ2g5kevR6idMb7XSbJQgRqe2CO0h/HOqUdoNQk
4Ld+Iy2IyNlaySc1y9vKwDegnzkxI6wmYalxOIh8mAHkNGp3RsjiZylywXfe
lQIaVnfXSuzJEvhy3RDU2JG7khlbeicOGFdiCtpblQ6HT7umo2ksyUkVPpYM
vo3oLEwhfaMhCs3ucVUYGVKNOUDHfAdAgP1hjQlPkX01Zzk0xhV5N2CP/vII
wyzijeQn/RsW2vB10TGim7rZxyhdFU2L7mZ3jJ555lWR1cSDgnlckR0FuQwb
q7XtQtNKd+jPOgGuZYqWsfWpTTTzjI441WTCouvYWB4q6iHWb7MAaJkdfkUd
KZHIL8krQ7PQJtFLlTckkXoyUAHl9qalgiOAA3Gcka29OjrLGzVANTj8c/4A
BVp6VzpxLliC+pp796FkxR5HvbOjxHB+uPQgN5nh1siSCrdm391ODFccUGNX
0EsBRHkLLCRxGxGowFrwYvknzMheW1yrMiVtV0woAv69r8lsShYy5dKCZ6UT
8i001eiJAXn2L62YlDax9E7wLz3BsBy42xK4OlnVfDbFcsHFm1Ov4Wgq6Cnz
r72FwFNMIcivvNPicj9Q0wTcMEA3fRiTJXgjzziN4w2YCnhLUTHk6MRVNwss
p8Eodt750nxOmh7CPBSIlymxEr6DVapogH3L9Cr7+gg5MYyWMiNrDCLzbr+Q
kl2RmJ3upnvSu4s+gJfRBVC2AIaF0oyDkqS8nzBPcELnkD3y772XJ8z62cI7
X8peFy6SveD1Z23F89V9zOkq8V7Rx3Rk0mYp9q1AuCOnov5a+q5G6QUXu9lm
iNhrwJcDbpI/ObG1XxgSBFDKKrvJjwv9zyOnaN90FoZ+CBQLqYyt3CdlA+rs
DsJLP/l2VXFO69E6picTC0CTGg5LYdOFsXk69UmcP3nTsEY8JwYo40dQoK5B
VZpi+lm1UW3bflsTeAJci6Ex6iO+T4q1MMNTQFl/MnO6omernbge8E58W7pw
WMW9OuaKwQck1uwxthZaM9/425KIyz7/cWdiM4uh3KF+XbYUlm1RuVg4mfDE
SD608SuEZPJxf5sxRwLxnalm3hpdQVCTyPWo4gXvvROSeKjWKo33LPs8ozNV
E3Vp08oWWz85Qqdjd1le/c3YZZt28hXXq8SNaSuRfBg/kUCBJTJMh0WzFmcW
Yqdur0S3EZFFiAtvus0ak34FwhWBUbsgiRKFpGvWn5qvuJlNc/JINOO9f1Q+
HcyMB4RaoRvP2iaET8SjXo+6bh8YDXaB079OwjWkHIR9u7VDBvEk4HcGCM4v
/4lsJkbKFy0mlYb2ZrmKydmc9uM+6BG223wFni1UZvR9ubPFO/L38dzGJlcA
3nm0ggMQtNG8t4yAAQBjDY3mkz7lx1JP6rdqeLn8E3BDrCDmQ67viJEUPh7X
FgIfpMd1kBn1pDY85Mf5tFTIuqnU3u6Z90z7RUDFKkG6xhbidisjpE/SQzo5
SuRTcsPMcsH7HcrrN1UZ3sPZkUyHSjzBKnZ88NszoRZvsk6I8YiHCqq6niDg
XmdAyvc2R28sSK8Fyv93m9O5X/ljwBRMStKQiNYMBzn+2sbpm3l4HadZ5Yye
3fn82vzJIve7oh7KsvgObwfIZpGTtOZYVZusP7V6fxEWZt3TaZLfTbf9DIrH
tSW9OzwRnpPLtVtVRVfE5mZF+XlzVTn4/XdqM6UGxsV0BbIGOIXkhob4aMCD
rTfrxLsayXbg5B4tc8vuTkNUrO30rn9nShjSAEIMVa6dvh9MTeU+gjF3rjsr
me/NitFu3BvHMTf1379FVtEPOM1PBhwuDwo5BjNagGm+U5v9W6BTZ7GiRTS9
egj0HbahNWeAol0/9nSlFoXWF51qP49Vhb9oBXbLYPOxjqwhM+3vF1HV81+X
dng3dGR5J3givYpZlzhQlbZiC1X/wk/1Lk939V3q66C0/yVlDTAWE/tg7JUb
4MdrQkt9PUeudIXpZmqQE4hzrscYDH5MrTmpXYy++Xle0xC9AKC/zuAhTI+X
mt2leDlNyAsDAGSeosPrJLsuFT2Glre6u5n3ZDoOZVnnXQlrk2nTTY5WGygY
Q+sIYDHrNCOvfbFS43T7ZRFp2huhHSPUzn16axM0O0qrH9L61J/0OP2kJfmy
jnuGKzZZI24DzFKpHxgD9VGHtp18GfwW5JjHilbtY7rs3ORi9d0cAQWkyY/e
8ijo0rnd4DZavmBz9kOBiCNiGbHFkrJEdPGUK5QJpzurKtM8tRzUt6P6fXEq
uGcMXfRjUTQKL7rVVN9PCY1GyTqpM7I83p8iRHjZ48u4RvxkJg9CxHWyaUss
dbS2kBVIWsP/McIsWwSqClWBUyplDG0HTCBhsWdiyTH1avGkpaBJjr4H72lZ
GyXYNGslsDUnA9PtuxFsTk9P1so+hmZfS78Cf8ryJ2IbIoB6xCNLOXYazJnC
ZkLjS7sT7ushOt5jONDjmG/BHgQIWEVYbe6yQZCk/BNHWfFWx1Mdh3BVhiwM
Q71zK2F0bsTxeMISkKqsq+6jID8IQvF1FxVUQCRIr/wtmwz/DJTSWoegNaCq
QMtsyhSOfTAFXn3npO3NtkdJtLK4cpuWoXkOWz1gHLjPspammQhXe0Vs/A8y
y9mdrnFTkpBMD5JmUTY3sjA/WXyYpdz8T7cH63wDEOKbMZa0kUPlTmjySbgl
57di9ejzEkGeaPk/dT4UTMGuNdghPCl2hPIk0vdS8R4pqM8QgjaQN6lDR/28
6SCO8Ds9GmL0UGu6yw/WfaXJotFJs9GIhC0D+yNRjQYmjj/epTwkW6MaAvvo
KlvbA4ygg7blQ3SkU91+v8Bv2wN8+lRtFSGbbACRjd9UQAgLgIjd2oeWrc2o
NccYBRd0jqVRWEBR0/qzxTHs9Aa5rIydCbhty/8EqLCYCwTPjdArlXYLgbS9
Um64PFdDbum2Odzrdbj6G/88Kuu6kdyzu7m19Dyy4E3twvMaCX9+URA4ZiS5
BnMrNl5+2sU5lKOvY4+eqwBsK1Iw9u0eHXecOvr6q4ILTEodXpoxVZjwwGtG
zaU0iGKiJ1V3JpBzmvVD03JY+LyHsiYTfR0Ui1pFVLu2MkuR+XirZ4gCcVxC
GY5v2Fm0q/VoDFeL+m7/inM4c2wCo6Kd/x2sC6+aE36V7JbmsVsK/v/rMf3P
abi8CLMWZYYUDR/wfxm95gwf/zN2ya1hV4Y+n4ZnHAhhM3kuUhbVwtmSeA0O
/BHAyFgb7CXQyfDOJqSpItvAIeJM5+d+YlsKIKPmZEiFeoTgza9nK3ElhIsG
uyz/gPFvbX/eKtZ268F+2itLSlXc+EVzWEb2OWYt+27/O1lzQFxVvoVuK+ur
jmgKj5PlRQYxJnrt1o6WVbxdkGY/L31d3em4QiLSwwrx/7FtLCjNryyfKDCh
GQ8zSAgj5/1anDDyOspAl0aAlJt30gfPBbFFWgaNsU/HsciBjkfBVKEW+VBp
MNd8kmurJMv346Itw4/LEsXkVH76d5+1iKk2ZonFZ9mImda3GJC63vWE9gfr
GEyT0N6VT+7RHHMHDUN/0S98tBiYTW1L1nM8TB7bSjsS3evKdyJ82nP89nla
Rhz3zHO9/8lsCXJOIqyNo5Xz/vsTFZ+8hrCTVRVlsnDqk1W2MGEsQSaIE0pY
lQFnCypiUgtvOs7v6lvz6qJso/ncqYfCCZ8RYX3A4BM+7/0hGVIpdsgN2woC
TwywnHRgOKWO3CnaV8tVuxxFuyKCGRhsOk8tNE4fBt3hqfBgbXDsWjrcuFal
CCAti4Yui0ZtQrQyrvebmeZ9qz1JcwBdyG0Nruf/wm8ivaGAQo0nAbWFdiVR
E2QtKZHcnh1Ct/xcGdGiRfsq3ULW24paM27HUQNnSp+BL7KF8mgZZs0WnnTa
TgRC4akbttd+KOrxr1AsDwnnq8gEtk8NQvrXWWxMNWjIZdRG9j/t6HtBCrkT
pGk8u+8OjKlKnWdJrUh5fE2V4QSbHdTKypJgWjsGt+2khpgAEPzjzjojmwxd
kQMeKQD7LyQep9YHLGAgV+Svw9MhYVNcO5kxdlHkUbd6SI6sRO71+SGMGvWn
rJOLV9Q6RtrK95bQoyN86W/67+pGo7iJ+4m0TPHmMY27N2b8URPoPN/rQm9m
wzL9TVMk948Cn8zc65O4j4CebQPv0aLY8xFXaEzCyCH0xQhCPlKuSm0fuSAA
fJDYx+Xq9SyvyM9i3dWPlFXOhE9z1Gcjg2Yk/CfwCTDm+rJtX723nVy1mJgI
SNo2FPf5WRDniCD2WVAtCTwLdkFxHiBpBdSF2VvN/3Y5f5OFvVbjrxisHwDp
1t51JFzbn2vjUPU7KcMvN+xtm0V0FsxzFSTUVczkueADVOcIIo4YHkg/M/pv
fC1ZdSMZAQRZRtJ3Ks20tgYjGNo6ig9QacchkHFLpAXPo9hHwuL20zZBmDC8
X3TfOVqRbGHrSfwWSZYAWgXFT7zq3/O5U+H0V9+ICK4jhQOZKD1UA6m9AEff
3i9QdkEOgq1biaTIBxEwaVx0n4tUjBGcaG6NU6iWMkCbQIXVO9LCvx33QqjG
4Fh2neZgowkHYoj35HmRVBaEaK18YsX+bd4ROrbt0bJtM/xGX0AifYi6xNat
6PnZk/7yhGcYIuwTlImIbht1JJi3vTSCh9afxvlrS6lXJn3XWR6Aq0yJq2dV
PkAyLpe1ujQOyErAPIhG6r2AyUyzlmJis6VGRdaQVrkl9V4Obd1DcymHx1OF
eLQBbo/uC68BGcqHs9erfaSUcEAHZUmAg5ss+VoCi16DmAptXrlengqVuKEK
7LEZPqFLxa8/v37HTygvO+2DIiCzfO3+eD3YORgkdx8+1v0et3dtKO1ZVght
Hth51DXl22T3QYQNTtrW/HmdecsBjRnnUdHMxUE1SSFSnpT1L+6BqvZlYjJz
n+psksiJh7Q1VMoWgDt6WbYWfD4Scv0/TaGUTZyXTZU/6wQmue6+ASgJ9ImK
XR76cgFqvYVQd6onCaXRmoyXt5aKfSsS80BPRGu5COrFFCl3yOCjvaCbRU+E
3IhHzcQGNWwjfpB9bARAn+2dozVGxZcY7JLG6xqosnAmoMtuAk+1byEoJgQ1
dhYrSgxfvvV62c3KTU1RP5/DRl/U6ayNmAqGG11oK/4g+cJTJ8Xyj97KTXaG
LsaPuxWNGvPc/fP/JLASAxwwbJoA+8o+dRm4v/74UXPoAHoyTz8iP2bVoNJK
MuL4bY3CmrjczmvlQbzc3HlpaH/JdhDBkJIxanlPf1eWrhT+LIqz4JHzZl2j
HVvQI0KrwKiIOCnEsiSBnzCzrAxDf2iJAXgjvwM42vp8Jaw+14S+rYydlvZJ
N/7bg6cdzwfYOpRcMPBg6cDnSEVcESum52+FHPJ+zWydisq9XKpg4WPOo1/0
xIw0HuiEgEBtvKhqafsv6xS7TCtcA2BqjMiY2FwNk1XywCXqVS8sHo4lvTaS
VxpffudrBwmFqhJajRzGwnSHkr5Q7Uwk64r7VMke91F7cGuSfyuOYVMSPxNQ
fEipJCdIwuqJr8kKipbzwueDDTnXa90dPGopw80JY4O5BPzHZtLvN37ihOu0
JeYQF/d7ka52K9ayLk9nq064nT5EU3v7rZ9zUtRaBsvqgKCoTq8RMDlf+wC3
v0N9Rzz0m4nQDl/KS886j9b4JszMLywekKnDwHzfcfmWa5yljK+vmsROeb03
sDQfklBSC4+ghN1ph6gDdhsqU78LTQa75RE1sErbb8GVU4Z6AkrK5ssa851q
T2KbJxEkgoRXyPdKpOfR5aIxcZ7jB6vr0Hj6DCYp3R2Mv4Z7nQ+JvP3YQtEN
ITbTroG80zSyPtzo0Hk41yJ8OhQp2+kohhhv5BsKJIBDNHObCv/tVR41jaDR
kSHjJq6jiKIUmfCZQ12MOdkpUMqsYH77S19KO8CrYY3Vcc8KgawB+S1iHasp
82IMu87VihQITMu5rRXPhCwG/IdZ0VnwhR3kmfFqdOEsFR6pWC2kcLEsj5Aq
XPhOOe7kAmYqIjlAcCHqL/swXmQJ0nutryxbrb0k9NvQLR234E2ZvtUb3Gt4
k0NU5Uwg3ABbMD1OLeIy5SqTdZdZOvy74jvm4FLvslvQyM85Hux3Sgkp6LG/
04WQcsV4RzjzLyAFypiIy8hwma7BaD/SmhgSQcOCRype9AfbyFP1yXZFRSG2
srmPndlaGupz/74bnsEdVVOqO71ax2hqD/UNjbJSDb5BfsAw88V4o2gO60bE
Jdgsmcw86wEwo2qzWmUTqQ3i+Y8ovHgyRV3ScjG9++jYjqcAuYiBFxwbdDtc
76vnN6mMvpodWzEAZpx0EHt1lt0WNIHq7AJyw6YzsBXkEJ18RHRwt3iMU8I6
f08rzT0XMRw/r6NIvxgZXi+4PLWcmNt9OTbEcaT34J4/PfOEUsa6yEM6v9cF
UZW7mSfNMGIbZ0Yr7KA6cQWj6dAlwcejLSITzO5TzDcXQPoWDBtYcAFOgoQz
ZYkQNAyC7XAxJFo8zsj6VU0xpc99IMqzDI2CetMbWOrAxaw/Pa+WefJLMwGw
2jn4RseRSlJf4MMEtPt+a1H9XJ2paqnQlnBJkOCnlNj0DRAdHntk8Udv1LHt
rVN6kXEkWMc1Y8Niz9vampnCBUWd5DksRRbe9JeldKyusl+Tr5yIJWKButT0
FtXd59brAZyXxDyl3hOuFBMXBRxnhWA5UUEAB6R0BwghHPdCQMAAKAIVJLic
N6jQvMK6islHvbDa6dLmwuz2PXyV34S/XJAAubhv6szCRK30y/dccL4BsPng
GN6jO5IHsYrm1TDVlxZo0ZuTdZBEiqSfzSg/d7dDP1Y/1ejtJj4d7xjvNk8v
SB8iHExADQ/WBgMQl4qxYlYVVwT4Agpz+0TlRHb3gu6/7bjWjE51yZIGYM2K
mz30g6LvxHS91covQ7f9KYnAMPbAx/UMuR5MOzIV9kn/WtWYR4C2MFJT+EpH
KlO3HqJ9rTyUhgb0uKP39pDvJFc4IVH2pnSpMtqZdzTTzHllXzjxO4nnR2zY
ba3yZ2dG3OnRRsL3qUs2kUi6gR4aHqyRPfXlrtk5NGTLR0ESjPl+SmxU22E4
qgmIM3mcoibETKk97SX7oOazR2oyNvqddh7UKmi7z5e2hjgSASdYylC6xIj4
Alv0ZsrNzvlBliOeq3hP38LCSrv9n//fdoFr4NLhvkMIfdLTk48iAZDNlUz3
NBHZcwfmfQbPPeufQ5sO1FHgkGmGoGXIU27/JuRBlOMfPqIVQ4mIOniwQ3Ei
XeBfXdFr24RxCYUiYRq55Bdx3Rww4kqztTiPRByZlN8mmMTA/ATzmYmD1yc2
gadEhSTTmEnL8NzFNZ/V8XA6/VGQnGW/46E1rW5GC4oAlc3XYAdW2zA4yGqL
A7885/CtVN8MArmR4ENbCeXpyKiZTcEO+BGQV/ZOffqWFpWo85QkyfD2csFs
Rx6E8/ygv9ipLQdUh0GBWot+Ny/bUTD+duVr9iA32SpKuPld9gt4IHob9Wri
sgV5XTbA5xNZ0iYlgIsqxg2frfK8w7vduL3PYTcfe1Ql2fQEDZI7RnypI2rf
P3JmfXy6bZYswh/Qj8W++LMvOZhrWDBDtlACdhCyXC2oBZPi4wiOxKnfvX4j
C3SQ+0ebk08g9v162iO8pY5yKO9MUnS/LMaK6y1cqBqHzkjIkYfz+PLfpatw
oCoFeNrkxnf89vWkComncMO/1x9j80ldMyC/7lNts10ldahEvAcsEkceyMgg
pKsV60skAgaoxm68w363qwUBNDRORj+NEYW5Y7yijzKovPTOS4QAKVZsV0R5
FEqHxkz7SM3+NfH5tH3v+2eUTploFB1PdJFtruoTYF8BlAWB89elYbpTM+NA
fJ+jA/AuZce87sXWWcqkaSR3dvmDQ0X4RmNEqtcme1Tcgj9DITWOtisy/Je8
15U37AEcs9GAcxE3jfHYj8JGYgiwJgv0umLwwE0SwH3wdq97uRf+N3lzj+bj
N0uGpwu5Qqp+I+B0iegMk4ZAN2pJ9tE5yBYenVXvLNgrMxsAFVBC638rSDva
+MEzeOFeB9nFguz0T6rL1PrizQ/cGyfcS6TWZ1nSn1ihPb9T9mGulI0+Q7KI
p1k+kv8HtRiY7sg9xL2vfHi8y3LhudyucSbiCf6sEmB/dboRReISGEkzhZhC
BBhQ3LfhopnYt0xc8EYyOpLJfZWCUUPxYanf2gp7txngNfxSAtffs21bRaOq
VqgNR8S2t9L2hkbWVlUFfCQ2d4zMQSWXoqZDNF6Qk8OQKhOqghRTrIdb+Av+
+Tv2y7zdMS6yBz/DjVaPBi6wa0bAtDZXUWvdTMxRWmabsBzOuBAeP0WZpazk
sL9K7gsrxFUWTvLHItBFSh93da1FlfzUCEakyPau6oIRThdShbnbpAei9/lC
nLHLdW85KVosUqF94qoZn280zGuvrKjAn9ToneaRG84EXdqQlPtXJaVBV2zf
m6u7LDj/f5iRDGaSxuSwonOpIdC8LnjuO3nG4jeWoeRRLWOquC9ez0WMCyqF
ARx+39W4OFvwatEFsQfdYOyYlmfN4iulikiuwXjkWA+E1yweJdjuAlXbPUCe
0jusZLaecj9r/SEeKSQ+90jIKEo/ALCO7cwotWhTMRRNekG6jFl1kvxTftcr
Rg/rmkrk2NlH793WLJgmOH90xSmpvVoaSy6Y+NDtdd+k3qkdtujq+zP12z9z
2EsLMWMLtmZZiBw28+uwlcCP2E1G8PnMq0U+Wo6/lF8tIaRKaXmN3Ddp+WaW
m1Oa/5X8DPx59IP9whnS6ZGrVVOTHzVvclkPXFJp4ejWE78FkaaHEeYrzb9B
9oufwGEupUnKiiYT6rm+c8VYYntjyRv3sNs3v57+zOWpvt2KKzsH1opYGCbl
PHe5qiq6SX7A4KMuLnaKprsAYB4c86bVGt2uD//2IKryIEy05rKSxvc7AyQF
xf1AUyAAv3DI/SHb9xhONYqz8J8lKA5YUHhu1JQGPq+OxxI/uGTEHic82iP+
LLxE//H1oXv8Ece0l+GbRq58E/grX1Xc5njhZIGZxjkju7+pGnsGoiocopyP
Y7ULi6QQGyxQA4NG1Ylo6vlxwJlTU8gkHgxMuswZ6RQBIX19e8de5hl4VAy7
WLRyhYivUuokRLmXm+gtkf/o6as5PG9j8k83RNEZvsFBL5uJM05ZHAb+1/a2
UmsfozdNB4zP1OlPSWRdgwVIhDpz8fhOSurH85bTxQGPyxChjsrE5BABL5Z3
oHsQj7mIl69HLxs8cbG5llU/IuLNlVlA6vwKyHQDodqwJhl2WWdf4KjQRUmI
CV1BZT+bM3Hwg55y9zt5ln8GjyLba5GRSde6dUjReIxCYKWCUcpw7DURjdDe
NE6VE7LmTZ91yzOKdZkJBfWjBzykW7w83NpLtH2Bv99xoOdvqIdD4tHgcXfu
0wmvq36a7O/fNa7ItQNizct7mRHtVVvB+6hVWP5MU8nX/WRKYLeyzgkxIwZv
vYNki/LEjiYwPxWVgKvBIBN67ja1vabngxZe+kZWgX7Y2fxbgcvTNsr24YJ2
0fn13TqNobPCMZ6+lkvXLYeE2HynlqHantdcIkLcovjX8ea+cAxns9zHA1A5
Egs7Z4vRzk3atFF+ZAWUfYxzbzJ6/RoSaIABhpS8oTWZrtnaqG3KI5eqEghV
+p961rdQDHHVQYTW+LAdLy/YSvlFR03o/0apK44uOs8Qas7DIwTvPBlWm8iB
PllHSp1Cdf4Y2amnaprpkxT25kjpZ9VxzByvXVgvu3Ql85QTq4sBrcscdHUD
vGXk6+zwyu4eHHjjqq5HZBOVvb5caNUTa2K1tazMSDaFlSM/xHgo0e7uDGTm
+/DX4GdTcb2LEm5juXozaqxxzxqVjBjDTzVZNYMWac8ONnAIBbX2LZFRw3sY
Qj+Rus0ZGfZyP6h2QypzvaAcG3Pfc0qyraVvnU0QAbSgNLsN93D6+SjIbA8l
8skBiBDUNWmM5tWa2VbH7rDmC3ildg7wnXEMMb6ElxAtd25AZOCzkAG2LZ7h
gIfQFmT9QlHIbVf+9pJC0Rb0TmaS2D5T8U7xUSKqpl2uaA+V4l1xUGEwkYoY
4FSHPzZx/ZeGXOlv8XJjYfZaeXYPv5eld1k4tZxdBYwE6SarEHAq5vksxIWq
qGRUQbEXIzBBKRxTSkZr0+Gi1cLIRE+Ua6jAUX/Fb5nTJ9F785E/hd8cNuPD
FnqFHJ/EO70B2R4FJwxhuz+nEHLsrbeX6yfB8XKDdgIVbIHk0Pt3ycPstgWt
4jTxHfSTpEG9ddVfV6IvFj4dKx3ssG4/kDGhz9zvWqS/7M1u0LTkJF1z9M1m
fd0ZfHPj+4o4AvJSAlMc9GvMx4psOiJ9M1n4vQC3Qy48c5emc9IVULw6bXu9
BR8rMCgP3VtMab6Jwqc/BpJzWrj/YpdBZAJ1ltHEbuznWn6TgaLvQ7kbql2B
3B3DmCS+Hr/UD/TQzs5u1Tz/RYkrQGsQ/x8k8TXsVJF8uydR6SAnI9nlE9sE
apj7sR8fVpkNmH8TIIVl/PdyvMWAnTqSyseJh5iIzpSzafxucG+JkDO4xs1t
X6fzTVEYBDV0IhRl8258iWdy4PaQ2VXf/L7jCAQxqzAQcFMTH94ogKqwYsQM
0LfR7fspC9gPHovHKBpTgdt5yM8YOfGBKCJRewgkPZynI54BXg4rvm/0JrlD
dp6w6Sv3PD/m0UpAjLBN8ys24OIc8nkSl/Uk/fyrwS+9pPTNUqVrO4Ayfpa0
JvXZwEDJ5+h6VhiN/CC2wlwprbl2SqhVguHiBiWu7w2BTsCIx8zw5FJbdOG8
Z3JCk6LeuPym9u1qW24GUlbxasuqmb78TTrRlCub/5GyOwNR4acKSOPm/3rU
P3Sul4eINP6gfKadkG5pOlNZOUzpivuuNQhQ7qBUU1jNaviECFNLqH4mZ3mL
H2uOc1khXV2mrAARcOPSDk1ahXRdJvJZKknTZbXruzsDAWmUahFz53WCcsN8
BZyoLM0c57tSAH0K6sIvY3dqplRKUcPRNAAGbsR1uaKY609WP2UVqrWO1ISf
/MV49b1HYQ8qLWGLhJZRaKj7tuAUQbQGb9KKOzddp2yaeS7QuAnhk5At2D8S
vqmo+1PIJ3dvp2uDPpS77ANV8t3CyHtQpfPxKJHlrlvXqFosTJq2Jzr2ojaY
jRKYJHm5PfQ64Bfh6EA3JAOfJ4dBGhm5GFcT4tO8HiSGA4r2/raxToRnW0Uj
caWkosQttZIapSmHr++Ev0loHygQm1jI+P9WEN6dp/PHmGS+955xTjsxG8Xy
zMSxD7KnIbG9PINvItTiqrjl/5NMGLoV2ajohaNVFMZQLR7kxSvYRE58dLFm
hhl6K9QXmNOyUaxIKt8pVaSEDaQRj6p/N34YI3RnLEvbopBs3bCHDhLazIW5
K01a+47yoJKNSUc2FlmFAxmzKgdH9nL97zvhs4/KbvtridP3LxdE4UL/rZ3R
vcDICDeR4fLE94Kj6QCSkV226rBZnHO6M84V3xT6uWLn+XZB3vZLzzwyTXSM
59YPXNwfYIB5yz5FbekWmY3kxh5DlvyHTe4rPeG/K1Aq825ZNVF57bnk0Rcy
a8RL22LkER1ZkvR/hs8KQLbDTZ0JdyOQW1BNZgMfgl/MhKHyAOOYYTiGU3Ik
LUpSQoDvZnE4CWnIoL+9GCZNZGXZkEKYeYS5o6O/9VE15lVl89JcMukqdCmS
+wELQGqtNKVkZJFkt1Cdzt+9+SXgX0kAoJQX2PoqEQbnXz4xK8l0QrXxVUX2
6bwpZxS4gFkbA0KZAwfyLzT4blrXsH0z+X4Yr9hBZg2NJ6ip9IagzsuBYC00
Jq7lFnXsfk2vlvXfAOYse6DwJtMaTOJMP9QKBzNoGjHb2DCtkIHYYhw0OC3R
Of1maHHi2D5I2/2FC4JJW1p2vT9bV66yujpEaQGtGVRV+g6zj/Vjh5iBUiCD
k21STelx7D92YLwZEhHVzSwoqVEasa6rkudLHpvygacF+gyOUZVO+qpeCLYW
VD9GSWp0FmE58ecP4oA98oHnwQGJk6DhgWU7tmKEkQQzc3M1zemcLWfbt3e2
Qx+lqPn5UYoOu19MRfveRnzjN9cV/Xh3gf1xONYEoNvVSsSWNqSclx6Mn0hz
fqhm/jAaVpyz4wwBRgQzjhQM4XF3QqGFI0MLsBD8SLuYh635J3amytgb3koQ
gPSh0PNCSd1GOv4m2pkLFmJbi+Ks67qvTNHZe7EB4XBPwK3CpkA9XVaIpt1G
qcGSYd2NMQ442CrjB0kzvhDy7WQzPjYXxk/3XW/0djymdsisYxvHzRB+dCAB
+tbalZxWrl1kFGBl3s0Hlrrg2MYHicYhBEWbo6WMGCfb8RtX0YMhiPwD/o+Y
dEwpdj1iWUaFI45tQkNUVTSWnaOHaPOP31i4tbAJDfIGoePn9Si1YbtbmVxp
QSVSg8FqAJrtNMI3n6waC+Ulw/oUEu8tVSH0lOUh2TR9f11sXKDQGARtizZN
J4C3ZgDCWCA2bDWafyHaB9sm4ANs3Z1LMmLLpMYZ+mxF7Uq8VoLAfSwdUoOr
taTtzyR4+V8Q4Xhy6F/4Hlru3kXoud12+9WS84b7rH5sXpyYsVGGyAOZnlZA
OjG0V/MQZmNjj6GQa773ZT0GFqdRoxmb7DWVpvQar0q09tek7cA8gg2p2bjv
duSU/CLMxz5/hisYk9L+kNIcMTFbQy54jbK1AbkLdScwhHqGlBJiXJUEawYh
g2kOCPFn3wVcXEPSHKO5sTrHnPirjKIDLAl7vjAQwuvoc03CDhGtWIrkddnH
lpEb42WKDFwXmxcrA6RrowYFI3JAWQa5vOThNjX2uomfbug86t0QI/nn3B5K
BW+6eJknUsPK+bdD3S4G1hyx0FqqBM+mpN8SmDEfQ49pToPOR4zBBn7S1kyH
cNFP3RkEm6as0+5JpLycxmKDSQc6QigNxhab3E+YXLiaNY4b+CJAhZC9ifXR
fFgu9QxwGjN8AKV1edLH7VRuzvM+YEp4XwVzGL2Ynqk3nFrFZvh9jJcMTn28
ByOqBmvtpnZKA4uN8REckowFdZDrLqWfR7vEe35pyBlwLTmCrwbkiuaP8IWf
mewQAp/gNIailq0fPYIP6Lq2GzXmNCfp609Tr0oHv78tb5Xvnnr/8pVjdc5m
SgkxjRg80Mu47YgMxMuWHlx8hv6nMLWVKHLhIvyqNVq6W9RU7GcY8bAeUTOZ
KCTu2JL5JA+KAGYIEpVNet8LhtAGAkaCG6JVNu1dJv2kqeixPtcbBr3mXEoQ
m+TK7hR+/U9T39Tos20ng9CH1zkG29figFl05ECqSRsgj4TmwyYrAJNjFbLA
3h3FoZYQeg0gf8nifZnEGErs9rIz/Mta6Esyeqp6gXZ+CDfxmEjTrx0qTNvd
5zIz1pXMhARuOM+ZkebuGItwI4P876VX11g1ncEvNTajYLqoh1Oa2dRgrPum
xjoiSQFeyw05Eke+l4Z4FFRYVyNVC0B5tCyZGJi+pJYDywL0a8/aRTYJbvc1
xDzj+qkUcn2uDsX1ZVMQrEsoE9J8Efyh7/6irsy1PqHwtqol7trBfFiMO69g
SRr3o3yQLshbm5WRowXwx7fPwboKexIQpRffmRwevYjN57DexYItIGbmugCT
sLHWgL7U2gBn6iVSEG5XkQBlmyCd5fwH08oGQWCnhsdUXPOtl73qYXWElnxO
JzdwTKuJwaWvisjfPEHYJGuEmq+Kbv2PcZpxssN3ABXsNu6Cv5lEX+cOMM87
6f8ByfMNGx4cvSQVEuJ0KeI3vaBfYEU6xoTz51VYwTp6L9gF7J37NWuFuuRS
H3UCufMS9JZn605SWDNiDGvbL9s9KUClIlSS7ZNU0VM+aU3Sa7/Yyi7KeS5j
oCVuaRy520MwmK9J3yFFB5jFzVmTSo9tlOFfvnoe2HCtUKHWX2T9hf+aPuYe
/MJZgFrvO0gEGeQrEk41ePlXZ0K7X+MprlAJg219c+Ja2EwSymwMCdrbwaww
ed1um3/4OiZBhYzFsO9zHyVU/5oRZWUunD0nlvySNDTTTjTKNlPZDKJOT7Gi
1NMR+j1IlFDyOMOw+zByal6d60N9m6XSnnCG0C80qlW/Be6LsaPToXZYDkPq
zu1pjTSGRgos3+iCON8nwEj+Gztc6suBCXo3OB9DaLNR9WcVhnEXOTRmLqnX
9hFWkkW3Y1pp9PBiknNMPofQRWmKphsT//9nMBRxoFtth+9lWTCwOUWvyr+Y
SjvqFD+fW5aiv4k0nE2DMRkxETUEz1/F+yeK4pGcdPxFBb73u/MFnpRhKTQ2
XhZR7Vl+qsuD8Y7pPkfUTgdWWCfLK4AAyw81SvjNqvVgk/K8EIomnQAw9V/N
+6Q4RZWfFBqeejxR+PC2TnGqyuSY3hKT7Fctnys56+1F25t6cjhOGRK49y0z
TL7aEfid0CyRmbpVR1EAaNrf109DhKCnRRpiYvECgZcmFu2K5qKae7LnvjWX
dvsUx0DsE9LkOfkL17KBK7lQ8pxHVtznN/oIldG3xdXjbLNlTTNhThBn7NGP
5r89HsBcy+zCNva84sJHRqUgAg9mfxJn2clwc3e7Ss57M8/UuZSn/dzH4+ql
8LZraaRSrb0IPfe3ASM9PQnMP7Cd3jlzs9MwwKhyl651JIyRJbzHRq2DHsTe
nmOG5XDac3n+sizlRjEGJPHgGUPVpgwuMSFHUEqUicT3FGrGOjgVhuLuPKFR
LyYbGsjVw4KbrKg3xWznaA6rWSfKm6pfD4TzrYDdV8F4OvmQrEj0jn3Hddmk
oRYeG0+YOm0cagtJDi5R8YGkOtjU750+h9hSMCjP6I7WNNOpcBXr2PFvICzd
sdYmD8JzgPi5PmRyBvEWAgjLnwzZWbB2NBdk6d1nv9YgxlHhQI64bRNoYPiF
5ohFqZ0RV8Gw0JWXHCNR9n1sj86+RxDdOUM7a86uCHSU3HlpZOec/D6KfsXk
N7C4B437DhCe8wr7qKM2SO3RVe1dS+XSCsS+lS130wKAcvxbSwdV9qAFiAVY
2vU1g+jc63wQaLO+qtZ7XAqvCzCDllO302JyKTwhbgVIlnMyf36mtZdWQURB
28bk19VQ18CJoExFnisArZD4pAFEMJ6bCnsp3yhBUl/dJfVFE0Kr3h1h1Gvs
a74tI8w75M+HFWxg2OHTMOxBvp0LIYNX76a17Ru7eH1LTYy8t9LCXIfBkWeA
lhBctRHKIa4DBriMZOM2aG4br1JTazMYBmn44Afx3t06ANhZIkeTsV/BcHzM
k6N3Vh0T+Nn8eVOJew5C5qauwfh+CbES3hHrzc93R/XRzW7mjjhXzST7C+94
qZBnS7dhOdArVWwlYTzNr6F8wZTc2HxLTssHJ/YFuWXDyBkn2VqsinhNYsvP
u4DqKed2tkQat+8IOavtRy11y0n5VKSuOwCyEhssyizOmecsMiUp+r3aVk17
rmeeZxE8TxbeDbCNMbltg8A4TV2HIO2UIPc8L8eRC+B5BJVJaqkLX0tvoFye
zytYD9qftms8Nlf/0UnpbMtjJwB69hu5xk6qfk1YthnLbFBtBV1ba7Lx2260
tbL6xLyZpFtdnAkcLkxze+8b44F9iZEpuILsQ9JUIynjY48E2BICKaRqeCBZ
UkGyuH5Q/z+cjNGCPKtTX0806hn/6oEYMucQTiR7sbMUNC80kXA7twnMK45R
L/oj6mfPMSBAiFEHVrNt+Xn0bCokMDZzHEkp9VOW+Cm8PCXEO16ywDtD3x/4
D7lVk9tfnWdxy6/lObJw7bxbly6uKc/K0D6n6BPs/DWxPcfOQ9h499zJg1CO
j1Q7A/MgItGCJf1KCIbLgUcyZF2pFl0HqSlb4/ELCQpU6rdoWfPmNk4gR0td
14g03Z9kr2uxBWLV3PgDhy04TTGM7xWYZ6BdHfKLfq8i6Vx+ZBQAeQUCN7EL
qnt9rG787I4aqPiExdt7M66at5VlGswzTDsW8VrOV8f07uoQgLb1vzgI1nyi
28/Cb+w0ysDD1FVVAdWJzLOrKaDqn4LlTA3HL2GuQHkTEMj5COK6fE8m2+NB
ueCMKP9zWsJKt2sptZ7n0jTdS/ZxAJ2KnXoC4xP81ZThSzip2OAnl4wWQDsM
pFHGFFFobKAgNW05ZTW9mp4PhiSGORfXZg+ox7SxeNYvisG7sUuOwNRjThlM
kL0eiFPrY5PHItkkwm3zKDxIcnojiHmGB9PuX0gRgKQiJvM1jR6Dn11Yvj1i
V99OIdP4+Evwb95zrIwXQA91watKdDaq2wpXCDKVTHvMU825QnM3qZaVnEKz
n/rUfD6ejWQXq4z91WgXf3qMOHVQ7At2Uedq72cO9JM3QLgufvm5XUBPv5iZ
Ip4PPioOkGAvdN1I87Nrxp1PO4xg933K6wFV0/Q5ISJYO+Muy9ZPBcfbiSYt
XNgZym7EAzcmMInZaJL4X1aWVzwMNO1hK0WDjfuC0whwWiP/Vtf+qaHPWDXV
PggQDcH027AJKvPuouFzgLSX1tI77DpTStEXt83VgwGOEpxCFkxIGLl7vHA8
b8Kih+nKx0GtBclyfJdMnDoWLs/L+yQgMXg1Z3MOryo2U07pbPG7BPTZsk6I
8ekTBWOBUcD/Qa6HSEmUAzKdnk/ddTIHkqzxmPLvHG2c/hflVZxh6uIwa/zX
35BwLRTT3mOwDxfMHFJTCMtXTHEm2m1jGmv5YYF/ZLeQRSqeMYX7LZyAZbfe
8HgwRGLUU2iYiodkOjsP2/oHGkZp9eNuJmagUcPcOwXE+ReJIwRHEHfUBhZ9
bFAIibvZypCz4hM2HrTqO0vCtElnZeBTc+4mSVMqJx/qXgLudcT5x7V2BfFu
UavnMtBFr+LLjymHaQyxQda7Xp4pNSWn8nmAVES8qmX0PAYRInqltFjtG/jI
mYU8Coz7/cPpEG4oDZlDwnjY6k89CbMhlxVTFK0puL8sycmbmwh95rAW0BKX
Frf3cCsLd8t6wqjwzkQIwJ7TVRESpAR1NxL2qOT5dcnW8ilJqCSINS0QNej8
EjKxL3+0I0+jrY1L0cqteRXZKs0SLPcBAAB0Bx24DJfnwwYA8QkCfhSbW5mY
u37u3b4Js4X2RX1UNpihNSQpDCydScM6SWfZRHLzhREK0X7jVugZCrrmhBYH
Vo6C9TfxOfKoFoCG8uPy4rGKr1WS7Q/ZdXE8CrnEVL4C6DYU177CCU/mH1lr
YR6GqiAFJa87azdRj4+LZm6JLy+lhRsMo8auULDheMxrVyDB2cS83CivXYE6
9VZnT/h7n07l//2BEIVj2uqw35xXSyZn59rYgEmKRrJSsPwVQe5MzIORgtLr
0wCZNGU50uCSGncuwhumKVqCcLkIOyvyMC+ustqPXDcpdnqRecx5eF6gu7xs
FGkHuU+ebbc1LuSzMqsBJMZLHR9C9jXFR4lPMYjIUrVV5vP+UdDBxvvpR+f4
U6YkcF2Rnb552eMPC0BEiA9eZwrPJNDEf4yhWz/ClR8nGMccGMud6p0cy2sI
AsBuGNuIHCwZkSMOkTrUYcsRG3QF9abuvDTytlI3NPB/0vIEBNFbHoWBErMY
smgv7SKUIhK3w7OcdT8/Na/WUidhYxcBgVPQ5yO7Ne6MS/WDCkphkyOdvlv7
/29egRqP950JDFr10zcoqM1gYHFwki2XBCp2nn+HFjBBE+zGnF7lbD3KtzrT
xDwI5qvQU/LkSX4tXG19DXrg52+pg/+EElWYxpuK3pnloqEvklfqMtMIN798
sHdllMLW1pMIATTICUxv/laMMRvkUCS87GTs4UcGnJosScHpxsRIQrfN7jS2
vw0yHtSethiDyJu+GNBrES7sJM8xDUkJNjbfiMEu7RMJYLLQ0m6O+5urqh75
BCAbW7gIxxJ6JUjNdQce2xdXy5sI/WBlaY5nGbYahR+m6PGt40QkO27CLm1b
z45oj4RPn/mbAQ3djDykuQv2pyBW+w6lA/6fANrbr8181jKRcPy5BZqe4Er3
6SoHMAn+A0rptAgDjH+KNmtqlkza1Xyk/+OcfXw/XyhTjvU0d7JCWyXwPEEB
l21xy5VRQA/Zu85Cjt8Aip4mhw0u14XF3C/1IJ8iHR3ZmLzFoozHMXoSBamP
xCzLCUkAOGBIFixbnswLt9oUvDsM6YCF+HstqIQRos682xQa/m6QE3+tKVVz
D+kZp8EZcRBlN8S1S1WSQlj4XvD+WiT/HM+2QPrVjGJy2HgEkLI6E0dSx9dt
EKIOwGrofhEL0PorOUmwfjG3Kj4X+exPJi7eFTeJ63hDQrjex7MTSJ/ciIHg
jFK7s5OuJkDRgCo5rnsC5LprsVh7WVulUTgTpHBG/3GglyjuRuVYDREeUbcL
0kzGEYiZhQUTOfBUOdgo1A+kL7qjg+vCwtrR659T4vX8cphbWH95BjSrL0Yn
f/eYQOVmoXyw9EvPajAjcheaagvaM8BNlRkksFrmj1Q4Tk972gGjleC7CN0d
aIWYqvubM5wJr5bB5iq/5ZWDoyVPVWfsW1siZhi5dXUPy5tIMG1SgJ3L2YeP
Ej1PidkaWo0WqCfD87rBgPnxEZ8YSnKpBehAQ2tI8wguoTH61wj0MTz/Hvt5
B5JPrXaJU6o+Ocqzx2feUg/Y2elfK62ml5oEgn/G4rkg2WUhAM1dnW4p27f6
js9p4gXPwoZqV6B95EoFJBWGB00m/zTlfDKRS9osTrFAaED8x4Y0qvt02xNl
lj91YFjJZOa16njiA9zAivin1/V3PyA9gy1+47mzrkKysp9Sc/jCaJ8OZuO2
sconWVUs3k1hTi94+BheU6SWTJLnodXThK7toEwb8aIP2uIrIFBc+H6SQldg
03sYwkyyIsrVbJ4t3vTCnXK2E8V2lftkNngYUUAWaGbFtMfQS28XsFpI/dvs
Sp8UeOkYNQJ0aIL++Bn0k+nNqEoqf66/CtjEDjJS68AplID7uBlR2gLfyF2b
MFhtgAnEW/6jeZtYYKxA6myY6Rj8G0TiTTEbbqKCeek2jFeb87RPvIKxcxly
gdHqGzUW+84tzoTzyCWrLirskjjQtFHh0h3RcakqR9JwXXFeNvJVMZSvmXcU
6VnZgvjREE+jcCyX9EQ0obprEIy39uiyBa7CPXgBWUpI38LCDHpYDFnLQAOA
grWGCtKWA7z1MhYK8VtuaNVqy/aS+L6E7Nd5Ez3UgJjDSDpKQBvUqcncroy7
+PJTvw7dK6ewd9rFwknQmFNXbyJuCKPfOwxE49OGR3+H5PmZGeoUeSxZ4950
s/QlkQlLNp9R2P896ASGIrToCJrI+WElk2s9Yuz0Ud26ygQP4o1Mu4OkTOiR
WxLap3RyTIFe9+JinoUOi/OsE7u2KjKLTAbLpVRhBpv5GWunSduf1nA2Rqls
8+ojuOBR+/lzDWs/zvylo+o+a/7Au/5vtkIowQsEzgVSw8AfHDzFE/3LwBIY
gmQDdnlK7uotAVk8cyqcPQ9B9YX+icGyINMJeurDKLPD1b/ciSNQb9crttsb
2Bt5LChA/x9BC6/g4abWDXYzNv5o/1F09QctvFuuUL6y/iSyQU7qDjQ5LY6o
RhG7PMtYIBbv4I6Mh4h1too/gbFIV5pLTVrI4LrzslK+e83TRdD88FNpmhEF
b3bOC87vCCZ+VW+yEb1TNwWeX4vy17bAmuSzq2Ev/vn+dHTcrA5NxB95uy2R
i1jO4W3RFgNbca4sFNQHZmL/cGDL8fCsimX0l8djEQukUfaND8xkLnFO0xiq
Rkb3wvDsU/HITJo85Weo+M96uqUiinAoCIUrqoXs35ATKssGvHOsJAqPHEjp
Av5FI0AucGw7qV0JhNWyPUh5iB0wZBDgNDxmzgkFtRkI8OX0GraLVvNOSMMF
efb6Dqf9czJo266XwRfYyx2fa5YwvQd61di2/RDEG3Pwr9nS9P6koCDwmwU1
6F+zj9zAp8OfqJ5r1hOHHqaepeWurU6itxWAMHVZIjddX/q523VKVGjgmqL4
I+xLqciI1b5YOAIeCZfAW1NXhMq5aaqFbBatwyHOoFv26RD1xhqwzRHLnSS0
mfLCdUkLdnFKSHdRYbCCQ9B1r/cm2qQ10w69BTLnWB0xNoZ7gs9Td4fKhzft
ugkei3VALv2MlDvNPA47ynhELnwVxI0Q+xnmuRwu7jRw/yCYvMbURkuGndpN
xa/302F+CBJqQmSeCEjhemXiplOTdsB8kWWUi69fWC7sVWV4zSjC5rTZ1XMs
ypEKzhPQNzW9iWG27oKdfBh+v9AbJ0duSVXdQtPA6MqDJYeNhwnywTDSeL0w
1f/eaHw89AC5g8zpqk8arxPQqnYe+wkWjdm4dkS7kca+GK2m2fCHl7dZ54S+
LoDlBV1hv49pKzAFxCjJ7ystticz1tnu/wzxIbNcX4mwloN+0u+2rupiiU0z
sPUEuQir6rilX0uDkHcx7etykpSLVwioWE0ewsqqllPu6uBbESzuWMScHyGK
f7oupJJYSM2l2EKh0AodlozhN3WZKAcXuRBxrcy+4tnNF20dohnLq6Yq2QOM
FEEvDqGTHXxob4lvxZXpCfHRmeUcdAByHQHRjpvj6lUJhgp+9tZ4D/i6IZn+
7Q/HgmcDhg5uLdAAiwc4OvVMNANqLrG+FBzFHSyfu6l8x1+SgzGnEK8rCn/S
gqY3v33laI5UGumBCYyWr7podaNfYyw9IfAWbuSP9S7e4hCOGCYafDYs/WeH
zpS0QGpkAq/MQIIXd7pIWihhob3YdbRxGBx1my2ubk4Gp+i4Oe7jbG4/c0lH
YsE1urwTtcYr0TJvIx/CmfBk+MLzm/WeeSLMZMvZtIQNPyz3IfBDUS2JB9ry
j9GvRjRgtZh+VzSccL5CYt0+WAqlOMDkNVnVEebORd4PYk944tArH+Ela/sa
EspV7MsCRWK/UsazKEhatLj+nh28JsEoMCHW38TyEpyQCCwz1zp7qNAIxQ6V
MK07rERsltdrBoPompJ7tmt5+AuG126eHwCl4VBeoW1c/VlNGC1mMmDA3Esf
+wHgCxu5egIGpiJ++XOx6fMbHX54NXsaXfmNWpJD1IR6GfPl1vlmkk7i9n0V
1NsxeN/4eG9KSDb9ay8V1FxMBVAxd3Pwo1gj6DoxHj9jzQuWKQK9LtQxHA9K
cCPBilPEg6bHtts/y4tXgpcckhDOhjkJyItbXQKGJvqgPDJe8thZYpWaavD2
OwwYLG9nzZpWYw8sYLHxtOXR3ZhGmoQ17QYdqGdCwKP/QKEgrn9uJu+/pHl8
DgHjNtGb2bzpigI+i9Lk96JIV33xO/MZ1oTorh1tNp3Cv1HZzCylzXdjQTmG
s6T6BeIicRNN1K+pFnDmIAktrZjnrLREGf9frTJI6QKxuqzG6HU4sCVS6ysp
XwRBVcXBCsa8/m5UOm9lxcOD6Vr0rMaIhxEHW1tj/sy9Z8Bac3/IFDVHjwqz
gBPkeTfJtCOaTzVUNDexxtPbGFZ61JNp7b+vxDJRqqEQ+SUyQXvum876FPbh
PshwM5QwBQZvzpOHQAErnzxDziAGwLTcQNn8kFlPLpCYzqta4q29K5gR04LF
4E/6YyJDn6uQEaV36wKN1uLTSnFfyUdguWJBnWXyGJN3tyY1efgacRhQiq4S
zxxZhM9sCUl/Q7xNMYJ7GytwXvIWSDMQRMCYr2ijN6pLoCnPe4YZ1PgROOPf
a3mMKzVp/wsiiqmk4RkdXb1mhkElONMkok0LFn72ERtvCjsGHp5r5ld7bQsz
u9f2mZxDSml7MQNdH0HpVPfX9CWKR3fbL4Q85KO8x2UiA7+re6lVggcSfjqd
xdZCbaQFSaDYMUimfm7ZncJWt8a7bMtTb/cA9bU/XWCU+QUy0cvDN0H4bLc/
4YC8/uWanPgVGwFOS6ja1T/K4isxQJ6yw1UW/qqKMG+w7K4PDnL0qy60Peab
cVkoSW6e60Fe/QeKJayvk/4nHbKbIpvk7b5VHLJpsCs3O/WMaYnyEPFqngMu
L02A4BMLEqflELq/TIAs5aZLbblCZ9Qlz8MXvRptNjgVJuYPxlCdXlzfFK8Z
k2xfr461vxFraVXG9yoKfEctYIf4S1BHKsv0fViuDI+Z0hgmF/4FAFwHqbvB
oJ6S7UmYTqdZJZ5IcMt1EcadTAxbzoykzIODfO6AyIwDbwSxj5ZaAgwRFkST
P8eTb7T55QMCZ3KX3YY4Z+Vc8TekeBBwg3X3njYwc07e9HDX7yn+eYW9yVDc
O//c5ZIu8vFYxcShhl5DhPcG7PalPevrMp1k967S3twz3uNFFm++LIJ+DbaX
gaIk9lUDsN6JguCYOeiF3TapQX3NxRBVEHgpjbty866CHRgtvvEfCUaax494
644hyLUYIwokZaus5vhs7V64EKPu1quImaoF6Ic1eIrDooXVEJ68qrmFvdRj
KaV6+CxR9qD4CagjMHaqK2Lt9WgBWutDYbJgEaj3lvfwsT3tbaUBKLM8mhDN
J9+KgYlaFqi6xg/2C8hBfcQ14a2qRirfVL3cfoTBK5f66blWBa0v8NFUXdas
FYguH979s/y/zfHPFnZ1XTifrEWfHFx8brVmxh53vwTPSZbd/NVC39PE8KgW
zN+ykryOZ4se11SFAAuWKTyEA/ICE3GX4CLf6oZ0jGow/YNFayeflOZaYmpu
wq6nQB9wue+v4/2XHpl0T4ewVNYf8TayfEG1h82Embz9cU81VVnRgRdLhkKP
tr60wSf9POkaJfy9dAhQHATJnizFvkLB4P/LvT+1dAiapFlVv4GffouZguQN
jfLYJvd6m8UDoCqGv7Z8IKD4mrpH0QiU4jlQPkZ2jrNsxrYOVYJReyrh63k9
kHitEklM9T4oWTcF4vG2+VzKqEDnfSNYZHXq46xQZt9OdZaE309M2drWjqVe
fKgqOZRE9UNE3bQ9DW8fgue87zg7bfkEFPlbqFUR1mOz3xmXgFJnyWJ7AWyx
6f/2N3RdY25aI/ESz/u5YvgomTF5wjFDAe3Kva4/Wn1f5Pm7ILGQZ+lv5Ehy
lISjSD+D7XviZz8gDvlWXJ8gZZ7XXolQOaXK2LWTq5zQo/gqYMeeKR3my0RM
nYOXn7cxq0Qu8TdgdVtbhqO0xzriHylLWrFdbV6UpHTHDINPLfUt79+Nrxdt
V8JKITW+V71/CM3XoJ5YKLW7XZWBGj7MR5kOVNxS9spEmZ97JWtggU1WE78m
ouZuy7g3pVjRtYJDOgOocZRoxJmoMghWxlzK2wUZo4nA+ysA2YTlD+6QVvJs
c3CLS3JBhe8pxoq/1DyVZc4cVCJGFcypaG+TGti+K0JOXn+wgd+YOlBrB0Oc
ussE+8GoEGPfCYjZ9HqgLj+3lspoBT8JENctsXyvVkeERbbJpkqFNlHjm43N
YmMkO7Yo9rUNYyyjQO5iIORdUfP6jrruXroscw8RZ/j+cVSi2F8qtaVFmWJ5
mQygJ/OP7y+vTYpc7zjSCQJpVmxIqralyaNho7CMwA3MC06MVGZP27qEUsPi
Pd3uGeB+NC09T42f6ZXS6tg0TTB+tcAg1ZPJc+9dbZCJrSZPEQx8FloYBn4+
8UyRLyC2HjJs6InifJnzg7wrcFw+DEMkZRi09K4kQe39Vo0AAJcK1ua/2HN1
lIm/ORnEGe+BU7oWdH8NyK32v9p9J5eoS1SPC60TvPKOfgShA50opqDCqUl/
nymC+dOleB9to7y8embK1a1I6s+EjAptrxC86VMhMd0HI/jxNy4KMnneLels
gxoJxd0YFP79gnuwh0LS8Yl8SkizsLXgN3Fs7LILGHxWO62Nr685I3jaKHIv
Dg+pxsHFBef1y900jkicTP6wvS3qOhnzzmXVPpvcg6vg+J2mznFQ//gpbt4J
CKOMPrqTIdIXoPkYFi0njAO6e3PtFCJLVaGbcPNdh1l7wsHIEbYdBenceIzS
zfaockX7px4t00dEAnVWcSPF5GT9gMVtXy7ea5RE6Ji3wRdIELQ3CvuaUxmW
L6GfYCx8pyX6+gtfFsZxKH91Ak/pUZrTBNA1aZjFZeLdKlVrfb3PY3+49v0L
o7eWYMfvTOwWBeQOEFrFGQwkHwrTe4cAdvTUXy5LU4EaL/BbPnVVhT5Li3WS
/+rNhHElhn4Tr8tsBuXMmJ5fnGl2RTb3ha4f1sSyk7qOe2+yZ456YtP2rCQ8
ckL60bJeCGqXvZhDfnqygxkZV5iaOpI52x0UVkTlW5EAr3VQG5z2V8NirQEy
tXSxC6rN1RQz9DiwSwPD8cNPLtm1ucetLqsvY8NdZZQ8Pl/Z9vDfkBWh22g1
uffs+sKVTr6/1QKUvVPfEoYY8YOR2zqz1b8U0d0wdm4I0poyldK3OmgdNvYE
1/tR9Th2eXEWdrXTltAt8+BBtjwSXU0vqZLMnjK8gaW1jZ76s5KADszXXVUk
J9Lri5qKjtJhy0dVzAgeGXhwTmYYTolihWgrnBRKuKeu0jbkExZ3gpB/TsWH
OaZUoKNM4C8gashpRFw5IsVqEqo6U+0Jez51SyozzNFVU2tVsOATgvZ9ecd+
C28GM3OyHZh3HfKoBVq6QRTROQrZprQiy0WGqLFc2kuM/HQI+mVpLzOAfCgL
fRYK+RZKakn7W2ERFf/oLbbBnlBUn/c3v5ZcGvoE+RVIVveRJaUJ9xcUu1Aa
teKdVuIbZQ9t/JW3ZsfWyxwknx0I7Osp7G50Oaqtv2YvMAUxv35cIgs1As/C
9L+psr2gBYh4dwea95cyomcGKFaxzO57gf5P1AR4hNgADLgVWeoFyk+izJIu
P8ZTcIIKYf6/0wCxzO1myCtpSU9noVMtKEjqeRhnzp82xlP4ya/a2dzc8iu/
p3Hly4dwWX/UQLvUN49wg6piHlOEV2Awsb0JuOLIcrGAtmQQBshtaYj+RGHD
nbwHjyjqJuslp7OGi0IulhLdErrAgJaqCilmkch4LY7zh5fHe+MK997kk0ve
sDxYOnvxUavERYunXA4DrIE0RobHFxksFOOpfKgnLac+FuTn3Qf3TUw7q47O
GqCm6T3QFOksb9U7y6IGxcdVbthoasJuWExv7TZA+6d0kORYCF1oy7ZPvzx7
H78FKyvXeM9GCCRIHXV1q61qWihdmSzTma5/wT+3jAmJbGvFQ645tXwkE/tH
MD2EhO8mDiIUMz4gNOdNDPD/w4b9Mq3JsYRhFFEWmr9XUZUznfLv8qbPYd20
HSpAhWZ8BecQVi19HEi6BLr68IWug0toIu5RM5icXUCpY1ANUD+VnCCyyivc
M/6DkOZ8cvDdZnu9DQ/U5q3noXDUQ+6ls1Y8Lxpt6nIctRJ5sXoWh85UJvz4
0gyHIA+W9hw/OUfb5JJ168ZLpIzI4GV6gk4qwDn2oIG/ySQaWniaMMNiFAHQ
zTm4+z+Qk+Z538ZmxwCqLaVf9cqyONZ6DqSCao77On90/RWjVUAcYyimlL7G
zGHR8ztSRKWDQi7WFJrhJCOxQuo0CIVdoEo2h5CfJN+vTOdng2AujpyegD/V
ql9t13dmhW5ErW9D8lr0e0LqbpU82Iym3aHgdGch5VISU11kwrWuieXUtcR/
iESMpPOJGNjfM7OkSxFRrEi0dgeRVe/n0iLph9Mrs70h6752C7oA3J6cBbTS
BXfBfZnmtclG2jH7hf6mkPKelNn0umxZLKphZ3I/D6mE/bkDEveUVMLXxk38
iFvgAJRQsisRzCiUEzyVxVgRLaOpMUAtTqtc+026WA/0n9t3fXUuxfFh2Je/
voqI6duv3iLzqXYWBhFNdSxLhmaUvyQYgBx87sSN1BrFFyThDVVQ49tvMWFF
bVQkhVvB/Kkjy5A5O6gV9jfT1+ZT/yPLYQd6Quf8fFuGbrerU4lyaO8AslqE
2Y68W97njQuonjQcLBrHzppGWgBTAEZtbU91O6PDrJDqupAmhQWKeUSjTHIF
LSHMnI63VERaw3TgnsAPottcgI4iKEUmF6yD93NwPexy//NAFdP6rWAU3Cbg
sIlwpS1R2pbq+cpmIY/y+5Gdh6LLdNM2y0fkx21Q8e3wN+mHbgQ9aeutOYAH
NaJOS8KpH2MaNOfsCKdBVPa6DZ9JbbF8kGZqKVK4TwwyCkcJfyzMkYcmAxDr
Rmp5OeSmmCdH37admwiU+yuCIJT6gFgWFsg5R0EjECMCZcEDUmBOsFRkRmAB
qhcDgpeRzgxJJYeNLFRd8+5NF5GGVosv47cfM78DyYNSOGguIhtSe+7PY127
UW6DFWIM1OA+L6fOfJF0vEt+E5ddkntc7OP6YJ7a+yTgWN5VSFBjenXTc9oZ
g6YLy7uvmpGCH7MluursbOzaGapA2lWx/86rHxUZIH9kh/2466a1RyzD4Etk
tFOEDi3s0GYfGylmUZGUBqfEWHOXDQvd/6Rmb3DMpaM1LG8PtcWJ45uAS0+x
XY8dSdsYbaK67bxdmUXvasxkggo7jqNWPXPKCKoQWEXXNcxbqYCbUhwtaw/V
w+HPGzOvOqFGS5Q9t+ct0enwprTTxMhUQchneYo7Xs6aUcGCIr2U+rjl+2LO
jTOHkRN/wapU2ag5I/HhBHoa0H43C9WHNqDY0gkhy5HacdUzdAavQtuUYOh6
ayHubOnXhdSGHghrFLLGVFbPaTYxkq7jsKwxiBm8+Ow8S3K7fhTKXNFvm/78
xkPi5LCHuRZqGBMJjqMf8TR2TAOJjqsfQ4fygE3e2nta2pUu/vdRra6uObk9
q7x0pFYKx3sImqdRwg3jm8ys37niisKpdAABuZOYFgCSduQboimCQytYss3K
tVmFHmCu+Dn+jL1v2vbQNuJQGmZvNJnsys1BQ09CTnl/38E4fFME7/PKPvsC
6vYwc/wG0REFTN8MQMfx0ftzvMf18G2SV6t4ZC87FCTvMiSnFHwFGI4U5H7Z
wrqZEY8b6VsqsQ0Sr0EaO4twtho1gvhGJDqEzXlg6gSun+3pcUpL648mS3UZ
YYkzNWQIRkgRvYdoRCabuoUhxjgMmmsiep210t/J9AXpDAANjixL2JRTgbnD
KNCw8fINeI4fXq01qNa8ZQApxZyWCA0FngWM1RBih5jVphwUMyNgzXR4z6Nu
P/l7FAJ6S1SXGo7kued5ZLgwGA+6RsiM4vjyjOluil7JrLiMajKa/xqUzv5e
JDKYa/3w/jm9B53D+X3uciUL1ryhWPoZzwIxQ5uaZeSwrmTCFquY2ub8uDKt
f0WHEa+z4Y5rvN50Re4GQw9IIE96aHUUDf3UtDt2c6lG/46F6NbDqU+EJwWQ
1VCXiHQG3ZxL602/TSMuXa9Q2XLSHfzgCa0yOLKZ9vd8Pi1aWuqDDcIDuPIL
D04aCa3FGIR6uPpTYucheOMFwbw8SM/nUbbANIEDNlhfJDOdaM1ckLrZ48Pb
zI++VFPBIoN8cXhO5I67vFWVGLOxeFmKeozCF23k7pyxClQ9qeheSObl9mnS
t+W0SNXbaeiosM2ZL4/O3HKnnjTPWBdX/Pt3y793P50Y2CBu0dLMyWuu3XWI
c5R0//Ff4IxJaZHqAXcQyE8UGCy2faJ8FoG3J+qSFrbIJzQWhYJS66Nc+G2h
LD+qSyxt7BFBte8/g11gw+FvFVwNpLVC84ev+F3a6jiOlPMrInw8JAg0vDLz
3o8GpgHcF9M6lTMz24Nm8m7L53oAe2BrBRgRse1mZFongzYYkf1GkOh16lS7
ArxI+paBma96iyGQl/5X8gUy/CuWB0sIN3WMqCRNS/Qz8QdFnDItrVR1VugW
+lJE9WIfPzRWwn9aCQhgR0B1tzDj8QnZM5zWIAngVSZJpVT4dkfzUOQs0+HZ
ghFMkJEgcRo/8Il7AtzVlFQhzHM3qI1YVlNRJCn79Ei/WDAJaDJ+TZU2axzE
8Pc01fc3B19rIvOkXwMzmvTs35x8Md1E/TMo/5L16oDAImX8PDFufEP0Ki4o
V9yEUP+D6leGI3dOtu24zWXA7SvFqIgMtu9Hlfp8lJl+gya9Q21JrrLY9zRQ
I/gxCZQXPpCkryLmYfop59GdB63OLpBJuqZRS6qlF31nmY6/D6SJ6zfxi7gc
pAMzJBlwKHdKx+rRe8Hohso5P0Gu1kGXZPoPkx6KI1c299tEhlZ08DWIuLpr
Vz4sSaiNHRdNsrd+owcSTNlCbQEaU2zLfF2/TjoYvNnChLODubWgg3JBr8Bn
L/SOGderJsHw7S46k81ec4umKYWIZyKd49HHd1O/78Bkih3T77IaYBmQESXy
MgNq5IW++bgMCdFu+lxJ83A7x5Nr0ia67VGuz/1I0eKr6Mp7/TrjX7TMLvCj
4njRB9zmN6qJWmVnIze54ExCaCix3qq+CQhlhtuLb8HuonxbebtfweqVmBtx
QJ/0hLjqHeoz/eZJrkmot3wv0hPLpJCaNQesyUH18F/JhKCM6J4L4e2C6Qw9
zYd1ugQ1hp+upuBDePKnmqypUnKRNxwn7A4pJYYOcX6RUy0gK7ZbzTt7FlE1
pzRYMcIjYWInpukr/EjVCzzZdIxLwknaThKWCkQOMSIizmASLcWnEdriXX3N
FG/yL+Qn/7oyA2eZ+bH+Slm562d9h9BD4aK57aiBkZt+/MX9+3I+iOYzv6ag
NZRVErSscIdMIz2VBGba2K02y7dlMQjxTXGRDdxjoUB0cybXpOZ6W1T9Pz8T
JxMwYfBkTVKrorvuVGg/pbo9dewktduoBekKVz9knCTaY8dre/jU3mUyw9HJ
qyu4aMI/NSBxrtBLT4qhqbjZ0a9bBxSW2khWOy/kvdGKDXEIicafKndXICNn
7avXZYZgyLeFyd7kbhFw6yiYF+vljomXKw51fGpjzPe+lR7wzJe0DdxRVKDx
DS1aiZBzXi0cKHx7+79qLjWpYFZxyfawnLlSiwIIp/nMMLtvXUE6ACRBC9Ee
9XKPZRI501TXVvTSYtkbcJ7mEhe9ln6/jML2ctYYmztCyR7LCjmch1olBaVN
2mXNHA5DbVY3pm+jeknIzs5iIVsMgv6b09H24W5vA/OJDnDDCJ54vwzdeOWC
SZJZAtbqaWQlVV6OXXl2ZCcZpAjcQ6WWT1OVSMbaahU1lpG52p+aBUWQfHEy
5s3DrDtq3AxXItnolJaPSd2UQE5KI0SuisDUbc098g7ee5NJOTLHPGow73UZ
rU+O2kqrWzYQpNH7FPD3fU1lQcOWbO/XIjeA2m5nvUx9LD+EASFdy1D5HqRb
RB7PB2eW2ESypLboXuLCwu0IohxZknIFyXj1+ntWhjlPn0NoF7gF6J08S3N3
SeFSazCYO9frwtneWgYQK044tUUlFzkozOmlLqOMEwRr3K3znNkT6CjNrVuH
EbnNjplFXQraquP+q3SIKc92YzkQpN2FOXtYj/FId8FLzdESzYVr8YNJByHh
aKYZPUWElKgR9m/MHE3UbJ9iCKNroIxXbSEvu/e/uWZSKNariGz/dJQib9Fm
a+DnsIBPQKa9U+1B1IVgs2zM54u8p1sDaKmQKhBNKeRxhl8odCCnkPLkhocs
KvmRNMzDx+i5+dcYvYDWGnC5CH0dYN1hixMr8W1gtZ1PgDfjSfFlHjDlALEP
JAqK4c98Y39Q4EIxnElH0IhRdTqcjsRCvNIJyk3s2wW6rTlKfx7GLU4HCNDZ
3vr6dPFuB5dctzh5f3SgUFJzls4/zSCYwJpY1AIceXKl1T6/8Igl3LfIgNZD
D9sOgaTY6T2DOYrAn45zACk0Vo30zyKykVULENs5+APaIBiwYcff39orCwQA
G8ymopzhbC/X7JPEBO25M2xFD7vY0ycznIt4ykxESXVQbijvZ9lWShBQ2J8u
i+AGfZyv2sICaa+7KFMUShrzHqV4MXFJBM2JPXk0rDDoiaieU7OdxInLdbs2
raDb8B5LTnj86sPujNGRDpsHkjAvv5wD2y8p5E2zWmY/nYjVv/dIouVdng9a
sDlXsbCq23CIjRsYcNvaofdlFpRvBTtzlOXHJv05ttTMEzsPnCeemDyzjT4U
o04wqWEZRITlbqxYAqcltNxiF8w+AVClsNGCjYOqJhNqH0JlqcqVpNvpx+kB
nDN5yFau+AN/0sywkyO0hHJbdHONx8pY5vMCgY0Q2jtRlp2UUJ/EWanDopr2
G6Z1UtocRzISAX98Hssd0TTuqFDKMjMywikja/4IQUIm83t6EjZidUWTNEQ6
0LOieglGja449yryGWlgLBxAtCpb596UZIgVqeFPxXmhH7rnCgxd1i1mtYrg
AFWgGnGevbfooJEg3OEqZLTeh/zBOyw+p1VepS0ruiGLmbfDXV9kwdFwd4OL
G9KNLrnCPvY65RVxCFhYqZTlnnPGZUYGOnvsReCg1FwKMI/2VwVIMn0h0yWQ
EbUoBG/AtwyrJO+cfkKtHucDhZWIZ9mo3j9z5Zkcs5bUu96PXAhP6xQuqgob
gesXI20Az2Z+Mk94oj2k+PS9lsOO9Vpih3V80483fcC0UsN20YbD+arKtDBo
5ilvEFNIF1KJG9Pj5eHOG3/pE1BHOJOPsU3r+WOoW2liAFiX3QL+Yjng+oKm
rdMPQP2DDgI/8GFwpH8s2zkja9kY9sgoGoQ/iWgSDvZja2Sjq1Ng7z2dYaPg
EO2WuARQhlFu4OcFaLaR0Z6Eg4z5fJLZznHQy8qhQDa3AMJWysGSd2bihAVx
xUrEpXw+GSkoxfhV1i2kl1H+CoIgCgnD3deTT5N1zvAyDUBBynP+O8zgcoYu
sfy9QKgS/U2tuxTdGpB85wNa5JAO5Si13V0usjFDOY/W46oubZ6dbn7Yg34d
7yCuFLaEDLYBIXzSFLyO3YkZm/o5fYZGvV4iANrvHKmupEVkFM+cWze7H453
NKdAR0aQo+DXozE8VqtBOkkQvn2/IYdR8pkBTo03vvToCKyR26+QzHyGwEqQ
ffp+Ayqtn4BynHV4XEzzSP+1+6rI9wUK9hzERG2xCOU+aEbxlXLLMsFGv8w8
q7/nMSx755sviWkWCvE88P+rMI2bbTHH33vqhuI45aqSJ71y5u8NcSpi8Z5y
JrB1rU5ebDZfu1u0by1RxGomFDxsOTQ7Vd5W5kbuIUPaouNIHpFEQxmcOLoM
94i3ibzKlcCM43wJLpR1scuedKn2rCBdej9DmHx0Xzaay5SzZHrlVhQXtZ4M
RmYLDhBr545zIt0AGWZryTcqEa1jiHizIYCUjMuS9c89qHHEbtYQi+YFQHhU
qycrVje5mBuRtOu6mP9nWLgRLmmOEyrcW8VENs8SSr3sA7/mYw4Qh1WNVQFh
b7bM/GJKLKLvgN/JpeJQ7gjy/EuNX4buxb4BjxZgNzA+zjtJ3fxvBWdRaF0r
5nzI83SjDhOGnZtBKQTRqhBr4sV3dT8H75jbGwJOou0jGElh4Yr0RSZuFL1v
yzQs7E09v67t0+hhBuhQTAaDZ1bf7F3LKMJFCcmyVanFd7IO6bxHpkOEu5vT
DoSPCDH86KNP/G9lSHj3j9Z02gqxh/NQlzLKNdfKPWr5VYg22wkw+fjP7FvY
4SkQDlZLriE1TXh2lNuz6Vv/cigy0ILt/hmHnbkMlpuiGXMTADnGPlVI7mJ6
11FXV/UufS+heo/jPcMee7uQbxFJQawwvW3OufDNRBBOChgkeBU2L5Qk4tzX
iGHIxbkGJBNfUabV0TYomfovzSOHjMYVvH4kkeWFg4kq1fTTaO2f4vc+YA/N
D3ACkRnkYS71ifIjH9hESdktXZkwj1KeCkMqac1Le3+Ed+R1VNewyQzurdea
3c1QbNdP1HZP3eHor0bwLQztEa0gYCN4T72CXDU44tUDXMAfrn2hBE9kWxqe
8iwqBrR22qu4RfKuBNK/j4xedzMA2V0HbPg4uGdF87R77c74rx7mWDv0slpi
iWDv83e7uOfGc38xdsP3/t5W3MrTP/HBw4u/x0eJVxsA81ioD0KqrwSyZOxz
uIKkTUtxDcLBFx2QqVqLnDd+PkYlE+VsAK+EstbTnFr2XK73reZh2bK7K6Au
o3L3b6/itPv+NS5QKnv1yNt/e8FZOGq1Gtcz1aFlomaOnIas0y7y4sn1atzu
dPqSVDcenPr0xrI1dlmcqQtc9yI0Akz0l5kIN5tvvAzjxPD20SLfEE/7JezX
hr4OBpYGP3Lhdqw+W59hVDC7f8LWEQsNEvWhiDFScdgSVX0gVzLj/K4PioGL
L6H+u1gwIKK2PxhNdAJXE5bjfs18NdR2wi+wnm8S/7msyerHpCWW+g9E6i2l
oRH+z2x5d2wXJ/J8fQgPQOE0ApE9lvL089hvteoRa55f38hEWXdZYbGDagVV
jaVgpfEXYdYOQay1tbh8dkp78BXOo+Gd+u3JUTX69YymnGng4Wwd6IWNShS1
pTMBCeWkvPuPCXtbfzvnGrVQ6e3JfAMFcO8qsM3WAV8E6yQVH4NvNeANrEPk
b8O8oB97fUHWGgnOK+OSOcolCinXBlXQZng4H9fgEf9bWQLnidB0veCzpumY
QvCkKNqby+i2C5ynu6LD1hEVmEv6x2BQpWqZe/p1Ns9czcYtNKnANMa3tD6V
6C1QKgCAeCPxGoMasiVf0OhxoEEdLttXOniCMWfrEf2ynMlPQ7uPFxMfiBzO
qD6pXxFc6FSlqeFINMO55xgEwJkIHIUEF9YN1iIWKEYj4tQUBBU/jUdFiqUW
mHlGxZ/3URFvZ9e1CKC5lj3JYHeip2I7fy9Q9Da9Nf/ZBgwcMNZ53nHGZtnV
dSLdyOtYM082iirDOA4xAm5NJIDRJcdTx5EKGgjoU2I+b6qfYk5rgG9SLHfB
9Y0VqGU754rTHDgxyBRp6JiKuGWkCSDSS1CAmi7ABIB4cmQvYNuCQtjTTCyF
Y9IxyL6kTM6Ovo45mYKWJebFN/epacTJIjYYuVNlpfK8Vcj8oRLPo7GxckJY
rGh2M/SpEsHCazKGpIWxd12iEvOu8kkwmnvuCtxX6RMfzDhOaamNI4uuPl5F
bhrF6LBVuznAPsxzRn9fMs+BrX+d7vcpKwUmPfyVciy7HCQtt5pxO7aZZ3Ck
KS2/V05hePl/VILoFrSj/3Mf/V9Rt8J9Ni7FlglbGYnL60imLPTNb5Ai93kh
qaxQSdlIsk9KFhaSrY3F0JQSE3ITmX6Fg2ee4FdURGOXw2jy/nXBENzkSH2p
k+ChYhuxDbQO512poKF6N8a1+gdj+K6N1Gra/Ly803wRSdifIYQPGv0WxNTy
ElxnlnHmLKh48IVhRyAe7XWtWnqRuEYoBUUWDhWKPOiah7kRvyRn/O0dgzU8
kRf6u9Ayxak1LGEZELnmOgSVKLbwtb9nnVrVuAStfR7mwhCRZKT+UNRULzhC
e+6IQ7jnOAAiCiDLB8kw4+Xt/7OOmhPg404jTN4xmGs2rwPs/gPNBBJNT4YH
8a/4GXPC/jex6EWsI2pob816eAA2ZKyMEY8d6rDTGoA84PHfQo/He5IJ0K2D
iOgIQoadofPCmo1ofOhY8cklVZplxH2fytU+2+hfZ+p5g52UDanT/uqieIrb
SfzmDzO4aKgTBH07qhnCAiOIunQCSIqsxOWWDrbkI+UG60xjHZoPj5y4sc63
1fEk0Q/GaW1WhTBtEjqgz/GUuAK6FTR9psU12/YakVlEsJd0yywjfCnF8aff
aII2jS6W6LKcxgri3bzX+rHuDd2v9zGL+az4YoMS5CwXVKvVP4Y7Nh1Z2fui
i//DiR8PBxwpRawHns6VmzIIY/4vN6wp1qMi+XEU5QgrJX+3j6UMNKYAA+mI
wovbTUKxBUmgDRNJ0su6mPYIqGLSHBFitzgzIHyqjpxPnOPNaHIhajrPHPdI
pd5W2lgLuP3w8sNuMsCZDGo2yISY0Gb/aPfH0gFM5+XVYXdsQMM3oMwwwwgh
evHWT4E5GGQhkUcD+AXMZjgOsYcEMxp2Wvs83sqjajC31FsM1ToBYlMkAXGQ
cSu7mYBsDclyWGrw4t48DvaV64vmEG3PuWQ9QfWa5ZguqWMFYNgUNzGmfhtc
gpibdf/17Tf/P9qpVbpBrt8xM21Z76x7RAXZb6Uf8F2XwGeTAsozZdGv40ZI
pwSpuxkMzb4947omGW+byMiXvxxJ4UbqsB2E2Lg8dM7UDsFdG2o3XV5t8LRY
aK0NG5wei6OPUa/Jy7mzfn/F7f+HY+QltrYtL1IIteuq47rulj2jK0ojOVoM
7uBLrrGOeKQqcGykrO0rBEfGeEfsE7STrcuZ5pLtv2ZPLtU3NirfOFmzN2or
9pVETRMQmBGB3Y7Rgy6RNQQYvzXE0fsauT5SEhzDZ+oXSs7nVd/+hUI7tuxW
mPrtXaHdxxV7trKtrikf41SmenKp0LJPVN0/L9XoZW3r04WsHC5O0uFnrLxE
OWGdhG3VdRGo/ifosdsb39DQ/A4FMYAKQ56Eyh8XdvRZX+o/lD3BkLRQra9S
XTjunDIsKlvhUj4wDcRy0UsKoGCtieBuA0F8SZi4IZh4rb6O3aQPNStiVZVS
JAjmnT84W0g8eJbbGHdAyhsvJGeh5/zrSi5p3YKIFhn2aP/u33uS9RRa7ZBk
OJLcb2byqBGi+GQ8Y2neaMI7jYsEbCFW5T6qLtS489t7Gb5KuUDjpAQgRVz0
zlmglCiUOTfpA+++VX/ITG/lGNGFj8w75dEmBmyN2P/DJOt5Hsd/hXsrIibc
xB7TMfAEM7iteuF8Ozitwa80ciPYkuCjV4nHR2w9Z+QMyZc+7zyZuiwbSfAX
IoBU/pat+022KEWzRzT0X3PneYmcGA3EIf3g1gB7ZHDelB/d+Ufc2LXQ1xe5
cktsM4Nf3oIyLfyiXCaXT3gDkZg+vxtueX68cDMEW+s9BYj7vFak2qu+izcY
qCsX5UA9Mftj49fb8iHR3MRN6NotDq1M43nLJ6PUA4BDESJAFfr+I70HtXt+
xVmylEFxPV/KIPF6i1gCsZAFGnhEj+k9NWynEFboOPaKAat0ecLWdsmkajCZ
cFQ32jXxLvplI93f4dyiXauThCukjH4ACvmBPJVK1lMdJuYuL9udWcYvD4vs
M6Tk3ud3G5MWcCLnwNmlO+RH2xKf9QcpJGUFqMlSVLrLRaN7hbFveQUWuZ0B
ROjRiChjdf8SsCWi6hqjonw0HLvyaedstvWhEQMDY1jbxTANYlMvlDj9JDMF
8AoXYguPxHjf1S0cwJGJjafA26n7bTf2IGcGF1KWnCnXWncbXx/MPZnFf3TK
AUEDKK3goPJPlPBy5L300P23hxO6wUmDbJ9FsAg/d7fABc2lJWvrVn+ZeOa6
W99FViqfGzJ99tLYYRQP5KpvWj9gP8tLyVoi+aNzp+BRx9ExNCgl9IEeBZ70
oJpHmZkHxN0k5oEau5In/5yXOhhSWJ5pFySnqEwyDkwtxq5E8SrEE07HZ0N9
fxdq5Z2mq0SyVCsCaJE99f3b3L6mQCQalefJmnoeIClfkf7o4M14NVyPwKuM
3hSll9Lhez5wgU0IZCgY8ktW4B782crkHtG7Mo9qKGtj7WRbnbpauYgKatEr
JZThWnE/AwOW0ZrOj2k4I66Aq5WIprVidZvjgWm97GUE1YmaNdc3GKsVy8wn
0LU3okfxI2XNhyU5jWQE2XPaZMLTmD2NjdvdGzCG0tDRrcbXKieLO+VziM4k
oShqprZH31R27BZlZnsik1diUtv9F0YasEMPx75MF5sdWKsre0/XI7Z9SRtL
IhgaPgJQorcHqhLQuv//+dw6nB217W+6AaWpIe55x6xkK84WfcRNz63oFv7L
NSwyktiUtbm2Zh4q8jCatH+wiWNDV9CINQsz5zr9frFOBZkKM558PD/h579z
zOhUA38VkCrjmS9POPCoBTOB1JwTThMa7tC3TiHaSmveKkkUqBKuaESdxj6T
ZVw8ri+V+9rVnp54LqDhwy1WGuvYWiKF7PK0Jpx62eiKHfh9d9HDTHEteXOK
hgAywt1Pr73xe/Gt+mbZDVqz+qFFcb5+wC1KD00fYjBkNd+7utztK1LXq4UQ
X7cpBtSljy/iOCZhp7sxqxSQTnUsrdSzzD4gOjHonuP4Y6hGqo/0o9OrzqN2
Kf30r8Fx423cjpMgBc21deKfBKSTqJMAAtkjtXNdZOFHyERH1RwvREYx/eiw
WD0Wdox1ZHf9mZdEUNibiGy9/N2Tht4Dzg4PHyUO7s8DCCpuReBPt98Qj9zn
VX7qYAsCN2+S/V3i7ko0XkuYus5ZWKyKpJagsGab/2L5LJWzv7FCcufoktkX
AMKNvilIuqAKd586iGKU8fg+o53bA7hGg/BJ/AnKul7PnaZ+v6hZ8nwyq9ph
1JOM20WWIC8zCZT63+LgHm5FdrX3RuQeTDWnvG8IZpyXhja7I7WX5w4CKR4t
045Q2j7y+3Abk5a+i+Wz3asJo0b2pM20XeRY6iY9zcXdcS+u0YnFyHQvjFQD
2yisaz8e+aS6DrnkGUzZmW9l/EFHkHKcDM/DljEuelvLh3bFSNsVKHTMSLhh
zK3m7eN24UJlAb5JW1VfVNtI1emCIXQ5EVmHUYFtwtMWumodOHQ+g33z/KBe
SsH0H03RiHwyUXw3Xy7ju+7dosUlMP4ud7go/o/DZgqzphOMhI9k97X1/Jlq
o0OSzRlKijhRMw8kA/Znf2HE5F8UVvmqnWe5CxPUOZv5d5Aczcu96iw05e4e
ujNlTlafihY7qGqvS9JWeFyCjUahVJJPcbWE69SwN4fjZkEPylnJM1ReZ2yv
vjKx67c6Q5Yk3QUXD16HBM232zKgQoA5gQwn0A2Hdy73LTrveBptBxwFM5YI
csFEcy8XRZYaskQILifzxLLzmDNIWOOM4BW6m6/YYozXElmppLugN3YqPNVg
D/6LwntGLSKBJF/+xHYzhUxu8R5iTkczS7x6hyl0whG0qYQiRc9PbdCeJOPw
NJ0jltKDUmyVLXGp2x6mdyYpxuLXkWuSpKTnrYTWtdjxQtAeLDBd6v1NaHP7
cbI4k5zOaEiLF+T/50Gb71JAH4MnkA40fzfREV+20UnXvU9iyUCIyCeMdC04
PqSoR2kkNVY62anFiOKFPGLYzTAHPVfBIwX3fs/LW0Q731zJrin+kFPNIiVF
hqBErE7bv+yoteY4ekDJIclIW72ZlRtNktmXz4f52FAQhvkYcqWAruUy06Ae
z7RlZZ/SER0TvJDvEv5FlglhcDXKMpNhK6eX2/C1vLypOKottJjjuTGv9CTr
EveDnR0rFCrEW59Pcd+FuIPiZ5QOzCkBz7f3IxwEKYh8gKW8cB0+JzPonfQV
frhwjcrJl+yPeEiLwQ8i/1HqPBpyl1xB98NAkxb6Jeps9OYB/DlEdFuwZ6W+
lC8IjTkjROu9/lK1Ut4bd9XeD9U7smve2g0/+CEIcA/vcNQzf1paIc7G70q6
S3Dk8MAcLc/nGxoLNtmTPO9AE4jGqiLN+FRZX0NcAuVxaTPrFBceR2xy23+5
qv2CVHaL2z/3j4YpTJgYX32eiPZEvO6sk0LcBGL999iiyl2s662/KtvL/717
8FqbW8olzjeIzz0xMX/jQqfJ4qxFzC9ntukMlglnE3q3klJF07bCM+YlBHy/
m+/WlqJjkr2dpPlg8frX/cTfKg4pDInisVXVlxvW2iBjgq7PCByr0s/WvcJj
FoieoRJ45V61fDpQzhe2uXwaAMPi2dLCjiLFmMeNShPLz0IXYB5l8Gs7MU9C
bWimygFtFphe1+wblOfiwPbfdoBYynxC+dxeW1Cih0ZKWxAjVcLuS/0f2cuF
tXkPl1G3Hu4AbBqMYuxa7edlHsbhHcCWQM4jC9ARV2IWOB2BvTAtEHvWPRsH
hAv2LSXl9z8ABabsn2HMw6gStEX1hxwxPdYUq7IJR6ufifi7lRAXg8zFc1ZQ
C2g9/TtGQlvjCNnQFBt30zK9kyLUZha1x1/+WsnjvB0nHRophM/N5e5w0ibj
5F2fPyPuHnYJJhZXkCNkt5mmgTemjpnGTp8uOecvU9AelbKb85LTb/8azMzj
/4Ef4eepfIuUwJCXNj2UgbApkDvlos2ocux0eJQZJV0254UXdWZvhUzAFLTp
jo0vfItRSHYaQgsWHMx/Zdip1VDgNqtW92cgX34Zj2Vy21FZBETBrVWT9Tlr
FR/SS45g8Jh7sneOO6mE9OuZkfojJP9mKFdrI8YiYvbZeykU0wMQOVJFlAB1
otO7fBHnbNEyb7bvKzla/+lTXT97Ylsr0TexZGc4HKP0aTjoKTyCIzyTr1YV
/C7En5aEi62NvSQ5TQdByafDS/2E6/swDo/wg36yqbQggdr2in+Bm5OOm4y9
N4N2jg/TrJQNzVA9IjdCz9+iN3KaCf7/hqseNM3EvXmtzdXIfw42Ss4WN9O4
A467lMfZA5D4ylzVeXPuB9jpGMGCvPRlodzB/rwd9MRL3C7QEqVH6FTHV3zn
FV8jRk7W02XXJY80Zv9Gv4Tycj02wnJTk1hM1zGLk8Ol9XVO71Stg7EdCMi8
CLqlvR3UwpQU0opK+qJ9cCeBmlXMAmRWh5Gsm7qVZisMsLTNUbycAqT+E53a
kyHusmtXlf5aWo7m+sAMAJu0PA9OnkOc83RHOPqOYppTt1mId3H5MffzEchk
rU9fxiFOnczy+OQpbPuqZ4nqbzRKV/Kq+6As6LR7Ifcs9z2TuqANAq4BVblz
sfolqU+bqlJEObMNjd0a4x+puhz/m2o6aapFMFNwshTm+drCx3bfpkeotT/4
N/aWMbm5zklhnziiXQ2pUat1Iaz1dQG+biTSW0KlviqSR48f7BG+s+TocesH
DDxsHRwhfDOXDLg5uyQm6eABOZ6giE/uXp9lvdKTLrSVp7fvj8iSVDWyZhra
UcCFBlqkYAxZUlvFfCcIKHZOp/6FFmMxF9xZv2/GvPkWnzF5seNusP+8fB2M
zZt2u1ROc3ut73Q6Uv/UAsQsSbd14CeKXbxSOUp8e6yXNg1fFxoPDRzlDyu3
JLZ8y9Px9zyIos5EqAVDLXkOdnwsLVF5JUybcbrfELPo42NkbmFzkN2LJlmN
4ICfze9wHChOBK4k2a69r9kNj01vueuBLvifDou5lV0rzwRXL+OQRroMdmZh
2wol1WWO7mn9c4isxa2sTQBq5jbmpR4UvOwmHHOnEmd1p4YKWWaVQCh5LbZT
qYi0LY+84788+VUndWSDuUlsRu3mMT8up42ZskiSnf+VbVNpnxUXZDaSeqL4
79nMeydBrmsE7l5s/00Er96tRkZ1n11QxuuNjJAhoIAKbM0w79nzTXAWYjac
VY1g0uhtLNxTwLgo1DKV6IFfXh85Yprc+XcBiZi1BUgY/DdwDJE5iHtNTeku
zLSRSKYLMlVZbseEKFFgo2l3O2tE/UuxvpgO8z2uwqWhH6FqpJz0e26lF5lh
kifNXixZ41dS/YD+wxZCYKqHrjjSOI9tM9By/zmofq5uNl7cyXfMgc4O99yr
h2d+XLqe3u1bIE1BVWziwkymAhvKIrb9rCpZbMwOBCoxqJQgAE0Ia+oWN1ng
39T2LG5f+gETeNny3X7vhGcIwHd0+zK3V7qgK2iZXijZU74PNDjb7D7ihg89
Qb3mrxuhIzszyzbvD+y0E2kEQrBqMES/YyMoYIz24L8lq0SCwY0H7B/orMKd
A5ypjyQWt//4QXvDq+8GY2ddH8zRuvu0zK/4mG87FWaSnWovbdZeQdaDl+6a
scOb/a6zis/TzjfFSCYhDuR/KEWg2aLyVbtdBSCKFtMd+L9irBlx1jm5i+VA
SZSTwSZbJmfVc+Gg2/SgLUZ2Wi+Vy4t1WQuVuEICvsEsT6q/bULeGELuxTzU
VdoB/KqJ6xusBg3nllOeNuBDpgZqfNziTpuO6ttXPiz+OCUSO4QnqN225+t5
omV/jiIBBaV+q7wRbH9b9cqHVcmJnwsC94pb1Ogy0r2bi0rQfMM3D5Sx2NxU
4wDQHdBJM9qDSepok6NRWO9JfVlq4nO6RTx/EGLqz3OalSSaxaWevRegnnbV
aJGoMDjE4WUg05PDKehHelD6nmNyjt72vE/Wl/Te22BQqwX8s3G0hwJqU8vy
LziOqfVqv7KziViL0GnNdhj0zOtqBr6uvjtXiyfTMTcGb0E4K+JFxV+8vjOn
HkAmMexRMnd5sJxJ5trJLplCSaO/ZzNGq8EJZLwGNBJiyEXBL3BiJLsoszDs
59CfD54yZIz/8JRfNKDCfj9yfDNog/yYWevZ7NoA7NELhg5mmwUS6mVWC2fy
XSt9IR/qCnHkpKYV0c/2CYK6iqAJ1/1gkkfKyQ9VgIv3HlZk4NKbOdmc2pSf
uxilOqsF661RSjJyDl8iA/FsN6IKuUyzbzgRNc3vQrAe5aasXGh6cv11/TbZ
jwAi1AQjIpSBQNOZedoRcVWUpIVeuKaZDE96nIDFGfOdW2PtExoR45io34TC
iSLdPZDMme+ftUkH64d018/5xNItaI7Sm9dh4bKJfO3rYUw6+ZjtlfruHTKs
pQsS42oUScxuE1IgZO/YKZOx6BUuo94F0rI+2gwIEuvz8T+9J3x8tPLGhW3+
pakAGNSwEGTCqnGb3/77DKR+v5fYPWwFWQ4uwTQSr8qUznG9tKJk/Ux3SJ77
0ENMZGz7OitcujeIat/IGwtl1NoMT53+TqrY3HH0FCWS4In3vCXSAB6iwG4y
vC3dvPBG+/DX40qEDnZtOvpwnTzrcxK75cnaw2Teymn6zX6znLtymKvy+bQy
h7vYLQfBXirvjyzQtTsaRfo4LrU3u99lCjbuW9Z6y+0YQoOY6P8xN8mxxFMp
E/xBvnXObaFc6WCchdO7MucsUEsJfjKu7tKDWAwKOpGHH0rxCZzO7FNKzJy8
5OQLCTwvPMxB7ZeJM6jCw3FTukEhJQ65pjQxea8CI8PATaTFAC3L72+ZcAp6
XUFLWc2dHjrfqRTrrT9rRWyn6Zpnn1DjACWZSsGC20OHNUOGH9yB8apLMycc
fiDPAdj71bRrX6q4Nv6TYyEIrukdwC2TxBHINNLIKcu/StRRphoBKbbvxhOo
lu9qzvgCZTwEA2qjSfkh+AN1inrKSzIKLFZANlTJ+LTsZqB1Vk19LnVOFLIu
iqa17d0hvD8qJueA2vy776JFChPwn966SmSG2oKS4cAJ8xPdJnNeWjkjZJlF
4tQqti/wfg2gfHiT7SCxaaRZeiNnOnh4nxdc7x34VkKG1MXbQIcVmW8Vg5JC
4PRI2EBjffT7zw2T/UEZVXg/6XsmhI3rZ35Vp6/6xT6uqmmHLO5BuZ98z00S
eYYwYc5FqrquXB3SBcqFfLyEjjYcvLX4ykXi5JbvXrNOAprl5qrz/meKJGv1
vbfgOPA+wjBgUZZY3UmCf0FC405/Iza77R60BMew3By/BII2b698ITsusIWX
tyctj97Tg/JGqMYzPUQSsjn1xFL30fFFaOEOICbYW92+BjnHv5RmI1C/CW6R
KEy8PqfP1wy4HzdpLF8UKabK3JoKldeAPUVa0bW3P0CXmvPLXc8250bu068m
Jf3XVkWB4a3mgFhI43FEq2OPeYar/bzOB2ERQa+shV6kXpJgGdLUttQPgnbv
+21tc+b00Igd8GQ94+pZX02rVLK0dge4K1BCu2kiMs5ycdIhRc6HY7hHjBwE
lMoYa5LnSmBEyCVMHyNnTxEt9fzNZwE5MRfgJBuBOC4CUyhUInwvIP1n5YGp
OylGTlSgTyIXyub/Oy9zNI5BZonaP/tfcEpAnRGXp/Z09fTYkqSoQgAXdIVb
ZW6iz3ywnI0N0mMEG9iVbfJ1Xe/5EF8EoNV1XFpJZiaJ4N/EfoyN2Nkzv/63
kwjddq+cgHwEuRKBWDlJ1uW1a6ZTdbEo30/WN2xESXcxSjruknF0WluLu6Ka
3hdocE1m1R8mZ7QULv6DxXplLXHav9TqrBDXSiiIIyW0rRCqidKcLemFJCY/
WnSPV01W9/I8OAI+ehj4082E0DDiMrZ4ykNkCQ7bO7CdnfgWnBOcn85uLmDz
vltc6Tq43mIJGiiKYgaolbO7M6vhNJOzPKX9L0nhqtHoT9BgiVZL4axRexI9
fKWBGx9U6aUYw6edkc9GKHv5tzYShGhUmgv5Ahf5RNWLg0edibdhtQEr+q56
4/RTY/O4OUzIbZzLlWef+qULSjZZFl2zjSa26FUByuIChIudfonks+z0R48Y
SgWfKBU/p46/R6Nch++G7HbaAiNhNZhaQ1yAugctxnvRegx7c2q/dpDRJeuM
2CpavsyrP2YCjoFFicDWsmCBjPeuplqMXTvl1eRj/4OCCgXQme7EjfJTrITZ
r2s7wGKnAlB9JgLJPxUo7Fyx5fFvScokGP4tiv/fWGKzhTaIHHwbNivcX0CW
ZVwxgB1zag0m5s1YXiYutA3db9WCsGGRl+eo1k9mzb8AIQcXqeq2N7kH1LXN
cLo1fY3ebTzMD7alrhQUQtL0VYNeev5/7BtWCspNuYWz1R9r0U8cNle9iOK2
iDwjyN9ClssirT8t0EIMdQfq8+tRZJ6bZV60gbUo8EBWYbEzkjaYH5SRCvfe
p+2D6ie00Vn8lNznM9/EJ2l6jD0N7MCc9Ib3wOs0qp3yculkpKTd1QsZud9v
ZPAWS+eZibTlwMOpqGLCygqOfrI2+RVON1UerN9/dlA7EZuW1DwR2PfODzxS
2f9G+d9SWKETNx7sQ/aeWZZLlZ/YbIyJcqgpNMsoByo1/jXIHZGzfVXZRFv4
KETUBiJhBLc5Y9pdHtG8qJAvtFNOeV204txJo4PxlXmtl0DUMnu8d45e9JaP
I8DhtFP3njtcXf58pc82oWJk1Z0FdLJ/roSz7eM64+W1LFt5aEMjcBdPWhWC
pzmeXoSFUiArnLKmwxSvpLfll6dOhsKVKAvHURCQ3rJ5I5ThZyB19HyICYva
Q6LaOP/kXvDHyzkNGcKkj8HIpxPlOLYR1niaZiFfjRmCEKUBQbhqYXVD1VcA
hsSiW/9mEuuaP0SFffu7EPsk20fAxlyqkzsjNnXKLUyf7LJ+WNYY8nqYXeAD
delj/6wciCWZt0Bc9ljhJWRt8OgKg1bhoSpMqiw6+alPNwWFELYschpgCuoO
3z/Rsj/QN1NJpvlELmgfZ+XUsMrdVybbOQsNtT+RWvVn96jOqjwyMZb0JBXz
G8yXA8jje/n0aSdZR/pMzzaBqzzy6H0gQ+5P613WUy9hxzPmgURvKu1XuhEe
2Sy1RuepYS1KkQ3EZMBHhB0KBUc8jb8YwbUh0SFPZqnrXCeixTl50iih/zT6
iA1syZu1wsXJNbVxdTu1RVrk7YIwmIbIIHAqJq54Cj1xtEIehEyN+BbWmkfC
HlekbU1ebgniqJ6481pfWh2LUZlCoaH7wkOSxugraPsjjJuUXt+Sfp27eP5U
afBnPRX/qMtDRAoViFcI5mIZyVXNIfhGQT7rGhRKTwlV8f2t2Hen827KlZNv
FFmO95PE20WLzcepItHUBE/NAX/ds3RA7UQywQxT6D+LrON1wOIkbCmB/z80
EHJSAxmT834sugkmuHQQChT9SQjrz24FnIITTtVXRBz5xYtYQ/TcZYrdioaE
yz4TQusz5QN+ZLvWEm04nN4k7oe3ZzJCY3Lf+oUAp7W6Cff1cE4TzouLjKmT
6q+U2ErPOE0nSRHz7nWYFN0p/Czvp7FaqAjskvn9zS6kQFDQwrqgBsFTqdoY
zSXF2jJpf2GybocGWgAs6QJt91Q0fUHhYZ2KR79MB0LqrlpSoaBxzsSBufVK
nF3yxHP+Q0NAUIB6SPDcfmo/CqBFw8niJR2rA+ApxBYV6qgCYWv5ut1HZjqH
M9GfFy027D0OE/t1fs/S0jlYqfMvp6QmxO4Sv5tWsUgVZcUMocXsTe8C7wf/
JippjHW6K5+gl6umrdL48U1dooozk3ACNxCGXTmNlFK4/RCzu/M1Ns60WA/h
P8LLDVmRSt9Xf7K8iwuX9eQfEPPx73q3PkPGlS39aNOQzWcfy1dX0wMk7Ynd
F/sWgjSgBeXpVA0k7hCDKRBG0iRcpozGSJcZ1zlElsXmNKDgm3Kvt25fOPvu
Da2NEBorhHfyjR5ZzH2s/+lWykGmSl69pNKQse4/9ljNWwmjDEilk1J/OvWs
Q9SuGcogVTZpdm4uXJwIJRwUxEQtJ+oCwnNLHQQA6bsyMQNZDhpz78AsWsf7
+/PbyUMNZnBlCMSsdZQkH5H0GgVnlkAh4gr8DJ4EOfArqOMkpfOW1BTneB0R
ZCpHhXUrsKif9JjEsCcuSqfi8s57OHw3MCugUgKmKnpFHolMWZXWuFXIB8OB
r5JHZKCkb+ji1BF9h2gRW+bpB4+o5G3vY6V6oebByS9vjDcrrl/iZ8TQTyaM
a9+9cGzaS57TZpH1lPO2cq4x5/qSrDw1K+dNuVStRdSHzniCaInqHp8HwapS
W/WnI0QXd23wf7JZOKfiHonfmgAACLA59fI20x0/fLLbjYR8NHA0h3K404tg
ipDuYU1BHgjXs8ATF5KP0eck+FzMzhGIgZ9KvwSufGeOMgvpgVeitVcqfBJB
fNEVpZA2GEWgyMNBYYVvnhGFPag5zNUzRG2iKUA+BD+fxEmLtfgYGpj98SHI
FPiQZUFE2Ym6Bs9n7oCj9Cr58FQA01YD5Mnv5IaSI1zxPYEg7WVsGH4MC5eS
3iiWMEgth0ooqGnUGhp8YSkK9EJrx1fBoProcT8p4nBDzArreepnN75r2H6i
URysbUlcoH2ZeWjVFEQPjwVIqZu9QmmEf66zNG5HRZkCzKqvi2AlSIvKP0k1
dagLJfMBGzJRn7MqDgf9IFHQLEoBG+yN0SHcPVuSh5/tORoFY0jaf2IFNbgF
8KI83d0nbFkgeWPFlwdGnHOE55kLg+kN3SvJeDhSnzID37xfZm5LD7E4g30o
q0I6AGoiAcZVGzWjFLHDbDhdd/JklBcYP1eYKNG1Qa1bUqqz1wz4qDPQ3ak9
Es9CRqJTDI+aoYJuQZQ6w+9zc6tXA+8WAamOCduoDdIifE3c8S78iNKcN13Z
QUJPnZzP38+iGiPz2e31tpG9N9p/9IyGHkQaUgWECqu3eLK4oRuUvxmjvJ60
Uw39NQMQdYQsKNwg8Z0zbx0jZ8caqbROhZMtheauy60GSx5nl4+4Cyegfvrb
H+gSzhMYVbJFgvhehspGsUDu8pETyZH4LE3gjQXkba26Jrht8yOaqxihQlhG
/omjH+GV5CrH6JTT7yuUxBPSasXALDHYPt1tZArRqcGED4CHb79Gz4VmtUvO
iKnyAVTvE637VJuhAcLAsyeAohOD+rUhp3kxDd6lyMRL+FsIUSJMFoaqA8qK
ukdaGRAPyJucPmDryvGjSvi/Ucw8sVLzw0hXes0ksd0aJJCTc0XQXx7+qTme
tSSMfla10RxZfExZ9HyJKOoeMZMYcVlm3fgEfApJPYFW0yQztwp1a50FeQGJ
h0tjr/BiAYijyETV99tZwKpB0M3OpgQIkRqZO4BVbCDAMd0RufuGmk6FHpd0
fkBbDfP9s6kHShYGbw3BTlsWqRI79s593lyflHyyirC2Ytc6JhlG9203kZ2n
046EfDgD/cXcN4lOUNoQRw+bBYkTBygqOiOzsQmFClHpkZW2Fdp59yV5K9J1
tGQW0E1JnOfJUWyHZ5KATICPsIPd56+1PoTaQulQ6wCPTDg9Xv6j+zTIxyLI
1GD6JXaiLQKspjjRrOs012sj8RscC7ZY4QquX20Qsq82oKez+oUZbQDNZksU
NDp5i2pGkKQSKgQtjhfC9PswiQCseoHpCMt6wlx+X2ivggiGCnWka74jR4D7
fYNN5f7AY3VfoewFlBRaC0R17Mu3i6aKU9EUUXDH/eFhnXRoJVS5P3AAlT5V
6Dg3pfw5nUSnnR+c4Iah7tCRbUBvH2EQee1oUb8jkA6lnQgFHvcCMzsnF9Tv
CdOEaNhgAhMF84UIBDOBqAMcW3UrGg1WSynBuLHiP9kC8BU0UbMduFrHhdIG
UODS0osmxcNM46ayR1MXk8gtzp1pDTrOQI5OEEn3YVg/K0ifnGzUKY+9Kah9
M7Z8bgw8Of7Y+ZhR2vNjMPBzFS/S7F9bTENeI/vAZbBGUn39QWGXwT5/OOYq
PMS3OU8Z2++092JneUSZFGfygeOKg2mjb4y27dzqVagK+HjjIq4uCm0STvG0
f3b2EBtZt39qeLJi17z+Z38KGBgVZRVD1NTK0fxI6naXGDGzRk/CFp9DbaGn
zJSyDCWXTnHKBIuGkHmw825tmY+1XMv5LnVJHZER/6J4xud5d66Kmpiu0Ptr
XeeUisLk6GdjuqfLXVmGy+0z8yhBPvWK4ZqJFowYQR/z/hfJaLN8NwR64Va0
wjox2KKxvbK7a2WmTWtEl/EWFSGhX71R4EnADeEfkUal3rqiFo6mI26xxjoi
gciCkzgFihjIMc0mhy8JKyxllgOJomrD+Gn3ab7v7p2QMUF8CMz5lzA7Hikv
JbQh/OCvQOLphkph4j34s1VOwtEpQG8yYDjKLOElywc6qHuahTbchGVOJVAw
cwOlm80jBtec1u9GsDoXxNE7Mkz6TXnriWBlWJV/zkAJYGP+QHNp8neWByqR
drmY1Tz2DPWfAzP9fGJwU3iKWqIs2btUztgNk9Zvry/Gma6S78Yja7tDolf8
uPnpIrat+XQy9U5OAUPcChiuR5NiaSUOv5y3TKLb7BwVVljedvMOPZLvoR2j
svE0Mu3ul/P8vyqfswWiMZll4IGP8YIh9LFXoYN+rNOgg3PEkCYsGX5fIBiB
UnGfOt0cHkec9Ue0V3T8LHvTkPvTlH0AQQAzFelsrUUKz3tkBkTBfGofQKQJ
XOZYnVRf/6esKebprMzR7F6I+emKiIN9JskA6DxfMvKAOhkXI+FJpnt00PyM
dmj3N/e36YSg7fVXezoPx9EkxdQ7lPfwh8HDQH211abS8UyuCkuSZ9lHegjA
sr3WyoNWTNr08pHfUWk0mz1y3miJA9vQfTn8xCeKhaHzVk87f/AVuOveBH5b
ynEU1PBBVblN5zVkSJs35+rzXL42vjIB1M/vY6amxmDqhnvZxmY1q3zeSmHw
dJ5IGrTK+9ICqL1ANF8MX+tu1X3+i/vGRlaBYSletYcSo5upn8zQlwkol9aT
eiBnJWQ1aHdzmJQk2qjVn0KkBIJpufpyHtaNHjevEFaRgnRDw1HRR9aeVwQW
drM4RTODaqIHdbY8am1Wp+8krOIEy69a8Q6SjVRdKWnGBqgVJbiz84SQNczf
WELLO83HgqScYIERsPZKEVQcPhiJ1JULL32wEOQe2aL4qpRA94VqG+2/0Fms
4blO2PrDjV5VuoyYptqhMm+fa32Ft4Njz5aMhYqwVgONOAsVL7l+AH7nujxa
JqaYF5pN6FX6OxorfbjAz6ZgOY5TczqtajrlG6E0ydDyP3qHh2VLWF+yTE2B
79OB/aJaqFjDHefLSiWX8/qdd+0KiR/+jGZdhuRk2QJO1MjiZu3LJRIkZWbA
fQaaNUYejCoG0nQQHoZ/P/5iox4W0m3LnzAjwhGj94uth3uZq11SJc06tAcB
VX0eJPOLeAJa4WfmTWNlTs8zjtGdxlwFm8Z+rS5+iCndfzYqwxBm7MKTkJ54
7jAdMbBDS2Z4lSddJbrS9mhi94nbTJK7gr7EU0YiHfbxspdwsk9iIPDThzKB
MnWm4R1cN0n2PRLjYYF612cKF+HnM5/MRk/qiyq1USfLdJ9cdGLHRT//Ewuu
2g84i40ByInqK/nDf+8yp+28FOM82+Uhj7OdVsut3n0f1modoA3V7zoUvtaU
Q4paqZS+d4FKo5UrWWCx18itjwiorlcWozLNSHoMaE+zLp0FqWUs3dRqRt/a
E6S2ZkEvCzTBgbVl1Ej5pBHf0FC58hQi21/3Z1kySflpZM1P3xCgnhzefjbY
facfif9DIcLsDqsYaJIjny8T8zCNIeozauTyefDWhgR7ervGR2Fi4nAJQFFA
qcOGdRDpDo/xE0uNoZzoUWrULC/PXIa24zbFZCeY3Z/mmvKVYrNSK6qDd049
dWRAcP6zsDyxX3prxv1lZDCxxAz7E+w59gsmyoorwFc8tS22zpY63GpCJomS
dBEFBO4IIGOZBc7TxZIpgnG48i6R39eJ8WSlDJhHOYvVjk1URsMvVjCjRgqL
irsHBtUNfgOTbQjGXsL5WC8PxxkK8VGE/DcelN4Zcg0jMs3m3f5tQqrnH6KS
X358uo79BY4wk4RwutLgqNA1AKX9xHIE3kJIdRMHxT8DeoZpi5Wf1m/apMvR
d/xs/WGZcyP/bArkGY8lCmfUM+UG34YWLsd6M3v3UlAeUsyqfJs5OrGJ6U80
TRr7Hz6pi2+/c11TrGa9ysHVc3NkIdixHtJdupV18SZWql6D4MKdGaO4q6i5
hruFmROmLAjCuqe6U5UmCk/3dzcD69qnAp22Y7qYlGkxVLutoWiwRbh7Bfgm
IHX4xXjGIg2/OPMyHaNfD03Io+6eisayDnOFVjhuYOu0yXOur3OeAuoR0XyE
ktEjMXk3DAzmzZleLZibrg8U2MWVvc6wZSIOBU4f1HqxRtcGJV0vn3iVznKX
OcmtVAlDZaiDZHl6fxNw7/ZDZoIXCx4Vp09bJ5KFl0ym8UxNRAoLWzP2WiQm
SlYjSe2zAts5E+6dIwz6pEYxeqqq73oIHCqXkJlpF6n+afM2pkYdviklLS0f
nHC5ygux8tEe0a9RwHzVjv4vZ6Of700JvkhD3hqYNTgBKC39LSsIMysgxGIT
eYyJR5lmXKwss8MYqwxxER1aZ8V3EO5CQ9+5GyYdAJUqcqKR6/X6QV5C9x8I
nZ/nutCWa1FXg3IuEt0d6+5qEmhj6Y21dKX3s1gImS4McKpSE5Iw1Oq4f2jD
TDlUBzLtjG/bUhNQrsOXV76DJaUsAYRbGB1oQBZwvhcLJijJR11t+46OB1Io
3cWSKojpN09WZAkxZBYVSWI4qo8Q4lZ/tDeJTkg0VSKTxGOB/b5DMz/PYROR
mAr6rhLpuXw/ApsEhtrZeCYbM0oVOl8uaBzz0yNHY2EcWyf87U9ZLE0x8Ifg
z+OQYlEM413UanK6cXLUMYt4f1Cuuv29bbIvongvQRLyGkq+6P0eYkB7val9
PYE21G9gbRZEcAfJRVkHqwl9LZ1bT9u9Kvmk0H6kTbTRnU9r4oqKL5DMs1vr
jKCJ+a9B8wcQgQl+MaV4g6fhwr7gnpqhMeQUGTlXin4RP31wvdk3cmdD2e0M
Us/6d5fXpow8KkeJ5a1RUIHeO2/8ZkRtAtH+G0iysJZFBO14s+NvdFCaRKRB
g8uxfLaiDYwRhyZgqr/U5kfi090VsZjv8EcAus9z2e/7h/giTx1+kg/5+qNu
rUXbcKH8yvKlBqjlsDt6MrAJttvlpkFB1VNr/R+Rm2Blwj/49v7FSxQEGiPw
S15NzHNIZXw/OeHGxQWpEuO/oZmXqtw85MgDRclQbEln8RAj0Glo4sLPOTFj
7Z5tKUz61v5qnMWB9vwoIRSuS9yvKBA+V/KxtcjvUSc+ostljPqJjQNAQzE4
99INbwbAuwwpR03xgcWSb6shl2CPbDnpY0PQJOgstEfybaIPM8Meiw2IBKa/
9DT332Uh7jqOe8I8sPxXeRxsfYzPStdDSbxXuJo51iCySNf1NwTAo26ekGAx
3lFS/Yo+nXJRZCLTYk9p/F6BjUnqfGcd8LbWXEbP2W0Gk1umuE4uq7P2h1vH
0LVrZS4I8qoZlTkpXRBzUaec63yP0HZErMAfYOkeNOlSknTlS7jjQowlhwz9
ozeeTwV0jI3xw9Br0XWSLy3YpZ2hNe+RUwrnyv4+wlHLmg0bVRR6j4AxmhcU
UcMNwhk415Zkx1hl8HZII5AZ2HyDeVtTVdvIcfKTaH229FoJtXt3oBTlP3tH
MQqE3MJJ3/fZi8TEayFK+fitGSGJi70hHqo50gjCzzDRVpMQrHMkpcT/XoWQ
yUOztNVtZ+8v/DwLzIydzYwvtUE7CFcmkGINVItGkmz0Xcar913caOj6kWez
5ZzBk/rVAWGca2bOL+iee8NnXL8wFmTBezhAjqWxrXyPqK3DqvJ8QlxzZTHE
LTYC9dm/ten5hN4er5bQ9L36pJxhBG4jp6sEh9DC/uTP2xlXsuBSfkQL5vfx
HXs07MjaumosDcr31sWuvqBAhg4fL//vCwoMgwZTqoHHpb3jwsKhyXl4Kc+w
MqkcndJzxTrID0s2/IAMD16fu/pp7c3TgKbIn9obFsrMjnnJFcLdTXBm7pA5
tKOCTRUvEQJfIhxQtNh4Hes5Ei0phk27CPfDcwxqdk/HttRAFEr66E7M2rdz
2aOGiDTMPGqLbCFWZLr320x0kITd3XtsAH7iC+HffTw0wbDbHpL91msroWw/
nTad0m4mpm8kXBebauxKhcIeKhbsiSWv98ohGdSVDUL476tWDK8oefms0uyk
+5Y1Ecnk+5lw8H7nkM32+Mk6zFrRhJb8qIPdW8lpmb3x29U73IEvDT1C2m6p
V5YdPTLS0rhYl2XOx6oXnw9vqo80eHa9goRVB2fSc4vuTLb3oaSrHGcJ69p5
mrqIZGuUYHuZjQsbHiKC1nQy6MfYe9JJdtMKKLY3q7J1xWtPAiscSguVNuv6
xdoWWKAhXjPpqbVJIHS+uKB0gHUHHEAgK045l4ymRqxEWVsXiQBG93NjZjXX
fm+J0l+fHxm9lK0nB7UlHbOoFVTsAHq22fIov1w4jJAT/514A0xUCRliosBp
w9rYsv1VXL17wsxBVP6+ujK1Z0v3aoLnAN/p4yMGpLFHxlWuuLwfVB/yijn1
Zbg/vxztV87h7HxJJ4/ngQQoTRNqiW/DM6rCbfPNricHVr0JYLlSrJ4AYg5z
6RyWj/AU6V3FLERiUaxhLn3V8VBVH+6ZWXa00hj1pxx0nPNHUUtQFm4hmzgk
06Zg45T1CJxu0QYwLqnIX5DBT/dZ9d45vS6xc6r9S+ljOUPcNT1sYCEgH7OY
EZVu661/7yUxBddLFEFSNWciWvc2YD1/fJ0gZuq6YgZ/jg5128T5doNihb5o
RR2x0tQPHblgKd1DnK89zboHVJ3cBXzwTRJc54k/ts9ndSASvirDSkHqwlZR
B74AdX+n/27cexBvGwG8GQlQetpKE1+FgIvAv9G/5osNcpfTovaZV7OCH1fH
DTMADNyXPb3fnYTPDa17at0DWcZOwqfxEi1pkoOz9sYxvChoJb50+6cmzZDH
mtAShoFncCJe/bthbG+HqJHS8uZ2eDOWDwavXOK2TQRYo6baFZOYFzMUEqe2
tsoN6njxpgEAVeAQWNZQuP8lu8ASTBZ5ay8gwiSIlzNJ91c9iKPAKAJogx9Y
h6NdYhkeHf2mK/XKycOTmIw/VrEiqVYaP1xHWCtqxa8TB2L6j8qFNz6mhTXo
SfUACvGJr5vfl7CSrPhZTLqqRmo1jCHxpns54QbdPWVJ+et12q5bns2xFPzj
a1zJ8iJyfiuZL9RfasCIW1lA6ICNg+X2HJRc96DFhieLd0d/TjcIT62sorqz
UicyuoccXpRNU/y44D4kBrk+WKBymEPGUhLJFK6J9DqXnCHYndL83I1PACaX
zE0Qs2O5neWb7A1kgmu3MCew/cuziPLsm0Pkn5Ku7fWrWFpfCfW12pFT5INa
SD66Zri7CYO2VN/4lFLAsP+zjcWHa1XqW6R4U8surlIYIsbOR0Qygu3Mp2aN
4t7+o8dq6ydZVElBxE0oMiToqwxm1M6cX/zIpYGle9Jehv8ta/ML6Svz44tV
dIzjIdXbRNHWEJlusrXP0Oj2GRfm59hFtvtQwI0floyY86eD0zsBfS4YMt86
H6NErQTWIUzyAOyRNcWirbnLBOBNvnsMJVa+BhxmRFxmWZZDj8+gb/as+lzd
ZHgIwa/HPib+dkjvBUNdUjWUS3E6Jq0rpGUOJDfPp0jXEePpzkTKkxKeiX0a
563Idqvzwchxw2e2pVgj/aDR5ESD/vynR0JI8LMqcfjHzPC6EY7S5R0wPfA6
KDM8Twb8E2I+/FELR+sWcMrufnlHrFmZlSRn1OPy3p1TrBT5Ri0aRAoM18oO
007bDoiV+yfw5ankGZLki6bqb/f4Y9kfSGt/lzMI+jvWhMyoIWSdwDL72XaM
C1sV7HZqormBjoEOVYxpStpFkRwD6TolSR9juKpdo7JavLOPRuiRx5ybJZIf
hy3pk3+iGWwK1GYZBneFpvz8BfFHiaVFKnA93ThQtEJVndY9XmTHCSwDoMuy
Yw/bNtHzaktfSvGc4LteyJ7qKO2Ywj0Jm+FwuvtVsV+HtDTJeTJebLoceu5B
ZDWu1SGfb6n9+3NBTdY9DMLl8DyRs9MBZPwt86WOTjSM1TiVrtC/ICfqtXL3
7B/4531Yr+xv8oKfj2cHqUQnErAf6gKzFBk3rUdqdU/yp7fPb8E7rf+o7Zw5
5uCNpwB6JIimmHR1GktXGtDlRa+8eZw2U672BPEh0o4/OcJ9g9OS5iBcg9Zj
hP8gdysInq3nMq1lt/x6YdWOTJsjmH6ZJfv3RzFFuTU0J98Va6zZJwdH60JH
dRCufFOXqQsjyOAc+VZ/tIKaznSOkmykASsvXRKMf9cCUEZvLVOxRWViO3W6
fCRhs94m3hd2bExaCnG8hb++GYWJMm07jlEFDlm9XvQsqDTCH/HRSvZxESPc
k7fqu5wRmxBtDioX8OHRyRf1bFREi2LjD7/rlLSG+k1AlfyHTfQe3FeIWRTL
z42lcAK5BMhXA1JnYS+47kS+6xiX05i7QpTidb82NPkm0oVBpqVPaujSn4L7
oVAZ/tkYC/hG1UwPWhXLSMbj+R3LU3R33Zsve6d1exnQ7W/7MxVtyNb6EcuX
YTpKaIfnGnFvwk09BHEZY2evbnYKNwZTGtlJW/PiZZfWw3wq4ZFY3jkUzABL
fIjg6il4o8NaCLz2RPRtdgngSP4wP4p1YruziYEjHvzAX/AnzewqSs9xmFif
RkUmMk+WjUhIfiKKye4lkoiZDgjeG9iPFyN6OFyprmS8cWzBMUKh478/6InN
4VVRY2dwCihxgwniKp0QYLgGP4x40r4E+IGyE1klFTO8di60TtH2PsCedmI8
aaaRVr8+9chp3w+1WwXp/dZ6Rw1kpAbKSKTnuoCF0EWEnakrgajQED0yVO2V
t+yVL6PVTtlbNnpf61o+yFaVuWDVznR0aCLJ98wqHZPz7GqOKqY2VUxn/ELQ
SazWKpQtdGm7w17opb6pp7e4/QfMn8jvpZy+4J63xeNyUT7MTLAW40faH7rY
ZeXH7EsRaoMehrGURPc8Xf9jG3ACEddY5XCAlhRoaZxpE1j+mSMKuDv93amQ
rWFBtFTx5vbkCUlN9pDZYw0oAwc0g9LilQab5GkgzvapWcrfneEQrJv1/ecv
py6v5rCgezz3FMZGjXN+I5cEFERdOUV3XXy9lqOFnDLvCFdl5gi4LoVJL2qv
qdjOj0vrX2OWQ7mctVeTge7kF5QIylbvbPNxEjLDILZCcAk628rXhV5b7cuz
050RUDqha2xixHxg1Pf4jJfZE2sIrtZbB+FttX9MV8tuCmhndNgWXhdUwo0z
gf5qgL6zXV8LFvSjWgJW/8X32RP7iViUJPTPwCYbgPbaFqc+PqVUXGV05/jQ
tS24sM+BGtJb0J6q0JXhypEH1lz6AfCHAFjLDcX11DRioAx0J0XWgD2/6dig
ULkORDUvPhDkk7ZRrPe9AOAjqfyQVVODN9cI9W1Vg0w/oY9oYjPaHWJ+oqLU
fdc9bccVAm0YsAj7JAYTnZTP/CmZ4SMWwsekWKpwlFoALKUgxKvTZh2XnRmv
IYmtQnQQkZ7tDU08GMrfpWg1fteEXvgvanLsjRz0EibolsoMnDw5dmso1ui9
gH3DwnkNNSADuEcfiMLlr8VipKoraTVkc5EdqNR0hKV+xLCWNR7WNQVvI1tq
FeUebUUkWauPNCstDrZy+L7napCxA4RsJTKo1VF5hJFg9If4IdJscs2EpLSk
J9izXyE0lgjDsPwKxS3gGg3VVBZwq/08PQfdjUFfel2OfLFx5aaocXW0BXR/
YJSsbs0rAp5bWCx9/fwHegka9cWhzImMwrLbxCQgDHanZbFzNV2ktWNOktc4
ndJsMFkz9J4MV9k2lJLjfe8Q7AsYm4if92hKMxns0nZ9Xbb8CtL8mZt60dAe
ZKyXY4Sq30e/YDEQ+mdKlO5b0eMmnj/NzJqwcWqmA6PfrB8pOVDhnQ/GBxe9
ohnafLcxWuoWaT7IQqbdm2l88uveNILAeY9EpRJvlRxW6oEMkcqGD+KmtwF0
UoILcAzYS2J7b3Qb0qACSJ7Z/iNgv+FCb8Bm9lWBGHc68fRSnrEp6+qRdeVV
I5eXN16O5JvxxuezPEXNVntlSI5GNem8gPF5NpUn6ul9qZSXpT31MVq+eDoD
eNlLYUaDgPftKhhELPeZ221sL/gCVSD5/pd7GUFKyY0F9rVaGkK37SAzIjWo
UOc/30PvQPNP5WmsuM9gk7nF28hcabQm9psu4RO+GPcx46mm5zLTQImcMP/a
Ah+Zc6hq9roBXwf+zundvx0w9mroG5bLXdMsAVu0ONpaC5HrndGcTx7oedox
ToLWJSibFXYiuOeKbYSWgpSj95drgvW8QSdXibKX/gj2br0Zs+jiIAR13Kb0
A7REz9OSRnqhQ8NWNv8VDQlfdWC2dCUuswulXwMCGKLdnxOz+5R41TKmH/D6
ZxNUPO2eIbUG6JUEgd1SNd9KzKZv7m2fMe0VzTwx7Xi4qrbKFFAH1LhjuiJO
J8QxrA60nv9NlldBqJFbCXo/W+0Frvxf8fL5WG0GpWZzhZ7vUsE0gMp2FCS0
Reat4OXCHaAswMJnhs7Prus40U/PGAQBw817mgfZA28edpBL0iBnIByRXcfQ
/X4Bvg6dr1sp1mm7vBQvw1+GaarxkaIu5VkpP9fGmi4UYO53Cwk09fX6TLh/
/ZF10Vh4yCOeiuQDnSeVnCeaf6g/f/rB5PqDE8xd9/Uyg4zC3m4cDY+FTp86
LhyROqqG2slq5ymDifF01q3uK74OD7OuKnB/n83bV6Dpzwez62+0GCec8Cqo
vtbmBWkkIPWkc5U2FqkN4vNfsJZlCZ3K/Ar8Du6l/hsmtyAWKhvvuHlOUECu
qiTVmB+4+yGWCMrgnce031BvZdDm2srOMrcMnzBef3svundNKY/zoLGVni1Q
2xrfcQQK9JgqIAkw5OfQTJEupUzL5QNi23YehfEiocT6/sMlbwzkTwxhqYxF
C5/9vK3dyIu4tsUZ1wSh3w0FiB4Asq2ysfP34G2pUQFunHidXNZ7ZDRRIZMV
kUDKIGGD4DuT5t+6NP5UWFuFW64HXzgYamX0iR0GP4jG4Q+xSZ1cB0SjdmQq
lwWHyI7Hb6BMdSjlXMu1wCz78Bx3rMpcKu+aAOe27ztczwilAepA2qsXg5cN
5mX+cUuwxGrbtpV9Y9KYdseO5qQUmFX6hRh+XjhXeEXaaubMW+9RhPaucHBH
UDMwnVmYt7Umaq3aF9nJ1T4+WF32XJDa5Z8mA55p+/2RqBxV+U3vbedO8c3T
1HfU1S0LAtfdxGjETh/ooAu+ZGaKhkw9OEO2GGt7oZXI5UEf686MgCuccV0t
g6Pg8rvWlE/vu/ZHbJxef5w3CYmOnbGfIvKQOKNRtPRz35+A0Y0Ttz1zosry
9E59ni+JG03kZf7JYbi/+ElCpDrLBGPJiuY16Bo3nYgp6Y0CktBcmQVYio4T
na2zk3NuSomz11+ghtbLuWgo99xE8vHYZ2aEeHq1YZOxPExG3OqklwwgK0YN
qWnsSUTbxrAY8THiLvpxlzqjpSN0RG48xCmIT74tbORAj2P9QWp9g4hwLd49
k4Iq4JVYr3QVTYn0k6AOccsvY5XvC8y+k+nUZxdc0SP3y/jioCPms4uUu4XT
KFMiuxUc+6nR+aC8WRBKLrBRF7hBy51F3TVZ3bcODtBbKQmth+a13TrTlB8o
7Tm2HXQssU8HUolYVAjpkzbisSoghRjCDyjSJ0IcQRPvgU1evUCetdON+o+y
N2y3ZueHJlGlWMsUm8HkBS7uvfjmlOdj4UX2WHP4RPgZVq+ggRPNuX41Y53x
9flRwCyy2EPrkA/iUN2GZh50J7Dd83Z7R34y3BSYzKyI7qsbrpYwlxTe1bc/
aSJcX+KkChxlpgBB9QxxWaHmy+1K1zUCgCUybc6KWCpcJSmCFLWR7bi3UkSx
DHqvj7ZVmnTls1b3fy4M/i7fjprui322VCP2IOzH4WLbwYCspnhQztWm/juj
1u/oWSQCXzY/WZq3uEKmfnKNZmHZ0MEJolwoltLK6Ww2v+bEAlQIbPowzO3e
vbrlyyirLBQ7jFeLTozm6ia828aWGuYHKY0vlzRHa8mnwSobietu4FHp3dTW
PE8GwswwRdkTygSPiFjkvV3gV8ptJaOfXgVj2q6LVyDAzmOmAS0kSpxCAM80
Wz4CPVBi1KiDT8MEMx3raOXEAqwinOFatKDXMiGqVqFhjYGOgVc8EJhU9P8V
ZHgN0yvJkQj5crnVoznWb1zhGMEVFMAeadV9w0Ikdj1/25gA4f/yuJ5UnCK9
+orFZEFHXdloOTgYnug+PgsM5ZPSadSC7+y9JB4xgNEiOXTaABEHmixGmazl
9MuHXY1v0jXEepc1CFBAWwzJCQ9aA6FLYa4SJeadO1rzUdL3+1jKORcJEomk
PEuS4ZpNS82ALlkBzuC8iQrXdkQWXQuO9CBiNP0qLEoIDm24m4n+UBF10xzk
SrgHHvHlKJjeSXdGbt5rmNiADQC1HXgn2fX4kw0vCyYzQnX90lyfhg23V/eP
N2HaKka0Mqsg+baViwCLGr67TrHR5p3MayObPrV+RVfbmeLjXDOeK6MdiibO
SpJvF8LvAYFtiNvcIjBquHnnoU//B8zioxvqPKTAMpl0LWi2k23ocmSPSVSB
ln1As/Uj2ufRyuWc7XFcUMqOslWwZoER1PEr5JPk3n78yXW9Hk3/izBaZc5/
KQbaqBsFj0FCeBiIcRus8w8UWRz4yj675ifqPbjU/BJtT1S/hhra3xRuHvGP
wUI89suhJiMorXsc3S7jhpdUo66Mudms7yxURcpF7LhJM2+gBHIWurp4zHio
rQQLT5NCbw0KGYUyulWzzsnkXNfkNiLZ5NdHMjXy6Ap/XvRrj/TaDBwuQMnz
SDQL5KFVq3nEJqhqmfQ7WM8KaN9f3aR4ticbpo4ezCJwfeLT2fknxBWE8QxC
Ei5fQDDnwUqcOGdZMGIjt6cP7Ij3O03hi1jkjqLXkcg/Jh2RURWZq96HM1s5
EhN+HUuF/Q6Se9thgJZJBZL2ByZoe6GCjVJIJ6LLdzaIjuid5Fuev0FMBzoJ
d4yXaRAlCJFvJMi1PtV79z23H4FrBDAXQEjs4AYB9ZNlm02RzEcYaCApzt0F
kb8xD22tOsvgyJs1DPaP+6bxJ3Rt7XYBOYHrkYPLBlgXfvWBBwMgIzmtI70N
OiWSfASXDmou34Ql17ImOwIGfLKOc+GplLyOB6Uyfq9gGXgek7VcFudsy1WC
MvnP6Hp1RHOzz77qOBGT4mWa6IbJAGkueAiOOUbAShgWlR+qsA8pyGZb4SYb
TBTKNeD4oKnc6BztryQq2h2/NPvRRV9+JGjr3WylDEBUpFf+zMz9MfBAq+PH
IK60inSZzOuZyTccc6pCudfEgJC8SoKWYT+vUpU6W9jgvTTQxAuUT3YneX1m
5IpqTOpvzFRZ0kJFMOSUbeou/sbFbz8XLgRCGp/Cr1uEf/+GQDdKoPDIwbp2
xowNIl90sAQ/hs/7P1ZXKE9hxaU9S1yT2BkI8f7Mgj5uBGE3Ru20rHV7b7jV
BHdbETJFJGu0mcAvKn+7Q0l/6OmPAVhUs1CEXWib/A7vTAR8o1KbZE51tqmX
YDivo3O6jDjPMqWH1ZiEhbQnevkn9yCr9T6wdg99+H8c8MlJ50VqYnLjXmG3
IGAiO7COIazW+uFMjNe36aBrKjAMocFIHXKSBtb/qYBR7lsxnbBA9bpuAPtf
VMiwgjzTWMe6FrmR5kPGLVDnksWUM7Uwuk9dVCgVZx4O6XXK5C89UlKNlvsZ
AC3T4GerqanUY8rYFGL4nuIJCygUCcrAf37NavUjPSwP/BpPc4VNQvvMEN+Q
Kc4JjAxQZIs/HpONSeBn3eBCJqE/gSNQ9fW5pb4/CkV/nazKqQ41O71VuvvB
6ZmXcaOEfD2b2jeZrh4r3Q2QRVCBsupVGiGELUKFsdjJROTa6mmStjEY2Zud
qYDtjjwTjW0wv5Na+BMd5wvctanhxv9aczBEkIWIHLZXWel1hAJPihy9yQS6
DdnMqlrqraTu/w7/q0F7il7tv1PUgDVYbcjJPxbQLytfF7gPGiaTdTM55XhV
fd9XIcFhJHfD3//pjn+RNw+b0NPB4K4oIXlwjGo2PD16bPYOsKdnXIZXqJhu
YxfhdQzTef14Yr/Ms8Krp20oh3mvqQ35p7OHkEy4WhHX4g6jWWS/7D7ahDbn
wNjoP/u26NucKXFMa2vYbySqmuPIO4YpP6EQcYYq6IHYwV4BI3/x89EfRy8r
N497KYGi10OHSze8Oj1rR/+TcQYOEQrXF+GbDDEiAVNQgStHSNuWTJxmV72D
RN+UPhQ0GECkvS1jQO+wEZ4tZUURvLZuuEFIfSZ5gLM4OjQ9X2cBzsNJwKGq
P9wP6IIE63K0Rg5wUiAxS2ZLDuVTH8TCzJqMkOS3XPKrC/PZUFfN2LIUoCjd
7PtRtdLh3bzjU6MflKDmWXsWw50UVETBlxn7at1VEBzY36sQ0bELlFaLYp9e
MAx1BTwWYEk6FTLUqEQ5YevGfbkyRVIm1kTQrgkwnw+1atbKVyLuJdpLYnST
Y8XGYRGZXLzy3vAOr/9xIVAEpJmhP57oFfwnkwV4Qv+MTF39qIC+oW1di13C
18Yl9P4wmd6yS51iOeo825sogJSY4XqENV38pkuMAL1C0BY1puA/I9dWcP9x
T5QEwxmEFomTZpEbj3lyPeVgmmWHAHVu2mjdmjHW59vCyaN2v/MHfBMQsORw
uhWYGho7PhTjly5qm+0kPy8RaJ42yCIi65s7bTearU2EweLyNLO2Qm3Op9D6
Qv4kPbwKOK7dCU9QgxccAwip1jLX/OARfhoP8jFMlOpMKlpIVIomlGs1ygO2
OydkRKJAUKEwGE/UUAqWLg2QIXbu9fUr/b7xFIpoOXhYOt4WIqtp0nLocFcM
M1x6eaBpa65frpdpmNdT+2tBJRWzeCy+cqd7w81o0Q4c3K8kEvxtJ1v1Wwt8
zV75VeDkD1bFilgxNGE+QBLp9PxwFSh2MH+o4XD5C43BZ3Oxh4PhcZAvJ/sO
xSq6Y7eyVnmyI3S74Cchr98fUmyUCk7ufGvGRyY9vB6FwI/Xdl3PmMY1nYPU
yB9CMqMtdmowHdeBLbEqaCZnpENdoRLgXepWvvUsFyRAMlRSfywpnHUfs+AD
AAapdMvETdOcrlqeRtythBoiwljpcl9X7ATM2CPw0AuUFhdxk5zzY5j7HXu/
ILzt3iLG6MHL6aXFZzultVuvPXa3ldzvH3CQFc7x6pmHbUDEkfeE4xLm5tCE
lv+PfXXP2MRZTs+3eWW7uTv5jPJCoKCMde2B0mBPOD6nYFoaFLhJCly3jvBq
cIu8XfcGQuSQV/8jyqlVCFlEFKESv74GWHP8SgPGhItCk+J60YckuHqpn795
JSqL+pU4tsX0+aTR5GiWsaD/ZvCEE8WESRPXbquZ4dYvOVgMzRDvTL53HScq
HNEqm1ZbWKXqKVG6o603xkhy/djoFoKfIhIcD1lxcDBNscifZG7gV0fRMUMv
nfLkmMbjikg4XUI+9llI9KbEOCeHYx/KaTwVrPhlhuGk5b6gmdkfceGnOVp2
YaaPufVXBqnqripnNNGStqps2uW1LJF/DsEMG3niCelNBXspwdKvOsKDL6Gg
JW4Q/xRZbplJq2OikxtmntcsciRO2sXioG9oMf3Hln2GG2HKR7u/cLWfq96R
mz1Y1b6YGOj/6jbv7LVHp4wvxKPznocAPqjcRxuJQ2HDWrQaKVNsBJjW0IvO
dvjmLDNv9xRZg9QTDcWtr0xKSJ2t+NDZYM0UYJXDB4UhL+V7BGm8l2WhCyWQ
RIzUyGL7ozWW4rbSf/ENPBPy7uJrvhGc9NEhhFTKvFPYk9O6S9XGxn4y98gn
aGSlX2D6Q7LGhLPywoufHOL/+IZXR5+B03txIHcUy1TvumENqyxYkpIb9Cv9
36hdT0EhM18h00C8JPD9OJKNbPU7x6tuO9pFt49t9PR2vnOxMV6QNf1XJoGE
jjbXC/pT49WdnTrBwE8XCugU3T1yAXQhqrrgZAxsResx1Tj1hNxfuEue2Xl+
QrKQft1nO61pqMvYFZtfcqSTfeYsxQcz6IR8wB4l6AN4y2zTiiXaUMrbJSgj
B+9mcb3CrXNO1nJ4tVaVpGMKySIV0G2S/bzQJROmKqVyPxuUAeNcYj5FqBnr
X4t3RHq+IqQJfT9PdSy2Uh2oLlNclQ47RnwALJ9HxTc0sSH4KYybsLBnIZSo
j2ZsXhj4irMqaht6PHItZ0y8tcfz7sc1MSerL+CmNmvNkbIXi/Gv26jvZE22
X8PeUcSkFas9H+65qa4iucV+iujciftTtOL1vtAllGvZv48QE9IHWLh7n585
TJGzls4BG0ncMGPD0CHWeiimnmvP385heFtaOxiIfnG8mVESBexsMhIZheos
gU/Ugo1aWTfZicKrkvoqObq8AKICQKQTzk+Pb3rWztJOhOMJPog1IOZoVb9g
/xfcp8zSOJHeoXAH6rkfmYLD5c+PDXQn/goMwX4dR0cc5bfdYz47ZT1MN28Y
ZVPjDfNK289LeRoMRNSNBci415t1ZRxb0ZgcX1usJio8C+14A5y+SXXer32q
KXSf3Rfa2I/UpHUpM/cZyzhN5im+K57/W8AZ1zY0xTPkuSdgXmSdQrGn+62W
HexxmBzn45bTq8U/4JiRe2hqcTLjETmOJV6PXsxzgLFJuasRwJwDWJjjW7xd
TTqp23DlW79f10coFOlcPqlKo9WZ2kVT7l/G0jL5QK+OmjS2gT8z/B3OON1Z
WJMuVP53UW5O0rb4ewFgaBuSxmI0BaVQjmadAxpbqOsYSTTkt462GOnNm9Hl
gJiAFJqDaIoM6VQuxasb6kVtHrHL4Bm0Upm085Ju7tKQikygMSlsMAM5QpfA
+BPCpgTCbe4pU+5Gp1MgTPM0mmlmbKnZxnFznqZ9tfWKnafGlt+Fh/SUOkA/
Zd2nqJk9bp9D6j48H1GY8x9hezmN6ALCyd53o+e+Hdnm4aVlKfvXmRC7M1d4
/DtgCYVfCI9TD3pDuZrdhKnjvLh14tfOqwCamIoQiERIQOoEyRE6tG7FlfvP
JZhiPSh2MLLj7EXdK6m6gjuzCGPCOB+wRxLesQLGNRjTrgjq2xmJkbEjqxNB
aS/PLS6htl8ZYFqaQdNkvLOWeMnP8idpIvbpXavziUaOMAZ8LTLQRYIOg2vH
g4ZtQi4K6a4vr1zerNTVidP+kOHJX/VIepREZZvdidc8+yvZdEgScheAqwXO
vmXMbrvgghaC3eeBllYB50X+ffiA1k1HS2H8MAbgUK5pu9XEB4k8NLdfyDDa
vw1VZ+IwEKCXiHiyq6KyUIyGtoeSWBD1HvtFPGgC1tRB/XalVlMAkhUeT4tf
+Skn90Xa6v87dVflIRJSDUFa/2LirpYrIFvxwk4CwwMUWqeeS9jSXJyBFHbJ
zHjdRbL7GBiLCGQ+fMtpNwbGGSI9nq8gvJRnNpmKZYwojbUx0g3aQybuzUd0
s3ZYgserF4po48BrQLMJgx9mKQBF2T/R2ZY1kbPC4/9I3WPNYoyye5aWsRFt
scFV+ukBZzrH7krZbXcLh1QUXrRT15fteJEhTPpyAGh03NZlxZCZOuwctVWu
obh/7hTHwsFW1FTqAW2Y9Cg9KWoX8Nhh+YEahLpFmuYOK2VbpCQzuk92GY3i
7H6DRASWUCCi1CsqaWsOh+5bKIeGzsEkakgB5h7zCdHzJJcxsDoj4KU16TNJ
CImW6dWCH1F1X6GkwHZsfsLiiRIvrg6C/HZ8VvbTbnuAOxKoVvfX1618oDkW
vY7b5EhY6K41tQ0tLbK1RHBVJ7i59sO8+YvvhrDHwmXwpIcv3m8or4Pf1efF
GB6cQ+ek/M9/1OO9BBadTI9sSgJIwIXGtydil4dvyiiu+d8MOwqHrUiRXusw
VXk7JWWZSsNShOqbg//R0xOs+0XgJVquGQW/V98I+EiO7slLq/7LyKCKaPUz
MMWi/0VOywNislLatpqwWVOlUvVbiyDtgDpsJE+CPGp760MkBrzRZmmRtAqj
rCqjRXTNgM1gC07Po/GzQ24S+59xx784xu4/vLV5uGGX4EQsYb5f/ip1iQ4h
4e1t8ByLYCQjTQWkSN6AL/crOjqqMSYtaAUlp/CrSY2mzakNbMGmJNVslDpR
MswlCEx34gEtBpQWv0p94LcJc5s8w3Or56xCmPtMxy9y3WXJQv2G7sVPszXg
rEGppzoQ2gEDMVaLKmfI7ayYXazijB+rMQkM4oEaiL2tuh6DLumJ/PwATFjO
T3/DiKUA0JhD5fkeIZD6eCb1fsTU8bDkVpm8o+BC3A1w2RX2Z9BU6QJ3nzpB
2qeHB7e4i4H0pALg+Y+qf/+TJSdcIod/WKgTtGgCat++zLlgwMoCBOJkvtu1
wNhB1aj3rrgPR1c/g/fLdnpMAQj2nQhCfJANkew1O14Tp2TG6KJ/pEebf8ov
iMDcHfzzCtMQq1dSF8IUOtmgQLC2m/voNFIw1LjW8KJw4viS2+7kyR9f0TSG
fEaVN0v0LoGzdesIoVPc/nXvwllOSPu6sv7ldibz8ii8zC1G1gsJpCivAC51
hBShrGM9qqPvB+WHoF4AsfpiF9bN+dW2ggS0jBhhLWHIsqytSZT3Laf0eIg0
7ir5AKh4Pw5o5shwFOtB/UqImLzBC6R3L/E2PRUcS7f5XIvcGc2aS4JusDdh
O1QpkiinHHS44YJh1sO41NCH2kRmjkBH0oRJNatgEAhnbkAn7p0cpPLrMNNZ
DiqsT2GT4JqBkdz12dYrxe9R2y0SXmm9MrGWJ/gNUMef1HLIIiYyjd8C7Han
FsMlcy4vB9FZisKqOzYSh1eTwmYXk0EbVQx7ThBHAcZbrfON6h4qDlt2UbLk
+E+wIKWTHGpAWw5k/7q1lNarnjQ8/qLckUa7E0rMzJ56ZxWtnfeY9Whu2NQu
acGE0oL/1B0UiZdI7SXRd1mjf+cECV7xrA+E0g4DEyWJ7o6PjOXMLQFIw/g+
x3mqnBwgEmsuo4oKRXcihvAsJqZ7FcoGxvwuyEHiBevnKq2mPnXGE28cCrA9
Ys7GU9G2t2Km4qrqufXyrnYxgjU2EwL3qees86c8+lFkCmidkC6aPSqZ0hmX
t5o5RHTPw4QjsyW0qn0EDOkDTrNCLMzLku4PTEhFqVKJj/ue47rdBZ4YhhXZ
redAseYgMWVKVqmIoC/Afc5DKAcnTvdUerLOgwGVfqTvSODpdzSRtnOtWPVE
79Wx0EyJF+0jCr5tJmfXdAnNaNAusw7fN53L9JAD5qHmVEzupF0b3vKOcBL3
eZATU8TMroR6Uijjh/aNKBp+82Zxia/nAfSU8ObylEImg1c80AWo0Bv6gGRy
QLC2AtXpL+Nr8C+Qk6sOeGUzfJ66uvb456yuhvGZe1gesqpL5zRjDZ1fsuky
aI2enW/2zpN7sdgWh3PBc0dbAQsIv/VxL6FgMZHvA9JjPGRQOEdtk/anTNd4
0lG3BScdkMOhF1fWJs7gRwNNoaAXwMQ4N8ZwLC5sGHZ2aDHW/4oDOmL4xLNk
hmvcTMM6R+Xy4oKp1cj0vZPziF2588efDW+b72F8rCtXqJIrpd6wsgxnlNeg
bpPyIpx6qK+C+cE79Z4WSjSWlNoJS+Wewg3S/JFbZmVBa7P39bxG+Sdd4Hf2
56JRIh4wQaEcMBeiR7bcUT8RwPHuCzg1kcksNJ05L4di08o/SBd4yhMkMoEf
3G8m4oWB4orCWzxYkBEjnXhzMlM1EXiKqfTxz8/9nOK7AgVYcW8sBt0Udyxb
9fySsN19GqbjDw0rHUmxwNsaoSQ4vwc7F8cw/XKzT8lVY7TiwpfE4s4A4GAe
0VRT6wvyh5B34csjunlK2hK+HeIHb0GfJY1ywTDTHxxxm3EH4LQcFEWrCLGU
9UCJEEwgACxly4QuCycNiHaTSnLcmDCcxAM+EudEtlz2DDW6bNg1kS0cAYMD
aUoTaTDq1DawnFTci+A4idwlaseQBCn/P5nyNQu/hfCL7nAC8teIjNvbH2LZ
yKH4tZVyc+9GOb0TrO1GKqL2lBn5oAhs1YBAOQSbi8w+yoJ0mbO9haJRsVBc
2WLeK+s7ikg/YmOQKHmBPRIOmqj12xOPobjZaZPjpu3lbPE0mle26BylaEJU
beqp+/2UZj1RP88OpFeyZtsAvSBLP1mefudQk1cntoaYroOXjU328WAUIL3q
V1/VvsuAr4TAZPLA82Nt0ryRzLKdFAuidHnPnNOejnUiuZMh9dpMYusdHmM7
xn8LbAa58KfnvURXNEZGIvtmLBGm5uKf1o6W2njEzhOW3X3j4V4bDJF7Hzdx
X8F2sn2VaPp9FL6/gnCwcWohGjEoFoR2aq+BizCB7/HmLet80WTevScU9Nik
+PiFNXOKYdg5mcyKvJA/SVxg/SyRKGa5mIczoH5V5ExpbXSHewTUcwb1pa3n
1zk7VdZh24swqyrvzmdqaBb8PQSiwIcjgSpPZEqItDSX+bMdjfYA1Y2HnMtT
KUtFuCNEXjM7sSBEtCS7f4In50nrcuCgm43f59Ooqs9WL8sf/KPtP6O3yeCY
K72/sur6+m+kqqpImxnlOCajAsOIxjlKuFQkNHW1AcE+71BPq/JnxhpxFG3P
xTgn30lr6qXyIbzjkO68LFF9qzTfQEOILfNy5waNEjNkrKTUbA8XOWD+XUuD
DKZqR1Az8fdA/KMYuK/QgmyirfZMaKRb1gSgdL4I5/1Upi6YIRr7Bt36iPS2
iRjSAqKktVLKRRK5MeMPasAQZYWJ0bUOiECfqp+isNsPWaf4DYEkcEbxmoQq
udutt6kGM/M4jJxwvAHN6G2ed2zVEu9E/ZJUmi2SZcg8BUoQh4BoGF594wk0
lK6+J06u7/0h+GSh/U4xUqL2B392470474UTw4egte0fYzijXabIlMis/ASn
u3jwiflLJd4S+Rc3YtTHmFxFCWklvHzjsEpXaletl6b6u7tOwhMLVH720039
+aEVYZp89ERcoiqnWiYFRR+/kynKN33zFNIzqlEZ21C3x004lgZf/N/Izz46
zVm/ArOfHEwlm981VhRBI7IReGc1mGks9fvBnXq2wwTJ+YNuzNAPEO0qg0Ex
97YYXk9mUF8AxSrGZhmrXqLcwb/gthLIk2qmiQzLr7XkYARxzWcCUHtfECiV
wRzW/t6gxFoOdqOIiN83ujmArmtB7D4XhDjjz8fXaKg26F7rbV+mcJE9XSuN
HVi4qJUnXED04tSWAHq9V+lHOeTvkUFg/8XVeRHay0P3/bxbamX8pnOibmkJ
xxHMcitkz00cCYYtgoA2Ci2WTojHqN/nKkPuzBYCmqUNjEAxXULAqGu+NrB6
a5l3E2XcmpMLrC9E1ZwaDBnKMhmFiRTf1TM2eRq6QhMNedwHj9oBpLlUnfXU
MR5AOl4C+rMtEVi1Gd92kUvTewcQSfMyexQr2Zd8vAZA+fM7jeEuTIkL4yCr
EnADeBsJRYSZw8rE6G32f5jBXvFvqWkHCF4V4Ek3tfB6SqeLNats3ACAl67I
dSxBIGYDqAtMgAiGY2f3zYpXHEIqqKHeCK3jKZE2SBFdWHj9hRbKhVRivofP
QSgkfdaTLKNMM5DdnHXc/tPYiAwYSXQ5XfJWqBbg/01Y5xPlxxYYTqTA374+
q5dR+7xnatw7BV9wgJw4x6AiIzd8tFbP1PBJ24P+SKr3u8P8SRP2HpwERcvo
n1GNT16pTLxRMaSVY5I6NYmrhXOE94GK/VIqiO1X+NAG119GVy7vgSx/9Lxq
trYGYyhw6+9bT2SSrIHaSEkhR97TflLg0n876F9iVQ2c6wKNYaZfEF1hrX8P
ecb1PuztZodglQiCh37LwEunBKBCeGduuX+RkvQB0ANgc0K1IXLlgiHdmZHf
hEYj5uTW960PYLs9/7GyfIBaVHqCHDgPaAV6qTzQKh5aPzEQ6ItqS3HLW7lp
o7kJFlM4EiuBX6gww+LlAGEwNqFBnxeC0fnSHnrdd8PlMUs2hRUQrxLV8tbR
9hnfb0niOUXekIDwO1vy0x5s7tRKGYE2lqqExX8RAcZFWS27XIafEyme+gPN
emju82sA6OYFnqLk4OVb7ihZLBz2I4udJod3HVd/oZ2519AqMqsKJSwzZ5Rf
gV51SgbQzRhlHiukfNDT+rCsIY2yaQ36hGQnf28GxDwbbwvR424sDPmsa89Y
IHApXRfIAeNNqucQYIOxiQkRjxpvMTGej3ecUiZKpko5xPTX0xwrLgdGhOI+
JDzUwLrkSyVnoVzP5vlXeOmzA1WroNo58V0iM1yoTDVap3L4BsmeWTWY3tz5
lt4GZDxpLrqFxtv4e3WilTv4YId2CvggR92AU2zzozluHqN/QPAIXfQAjk/6
J4mZ8iAmMO5pvObNGGtP5t6KZB5zJj+ao9q8qsgly5t367YXDoC8X2sliIes
u8MnbrKTSwou4JyKr9ej2U/JQwSxFnKlivuj4va/jniSqWUvd0WeCkIBY8Yl
AXaBq7XI6F6q8bhK1soij78gBXV/307qj1Nl2H1Usr3lMvF2DLEBc8cbHs84
WblgZD5v0VvTXL7H3Cgz2mrh5YwIkNnqyCYMu66jcM7H4uDnf2/s1cVw49jF
fxvO8TlMwWeC0gbg7KcO4R8GNpbUzmkErd02T5GRJyfKOb6iKwGMCEucWXVa
7nDyZwOJjtUVoEGPAoaGLtK+jW3xYyKqzA/3+u1UzCyHwEVzJBu9lDPNec42
AKXMzpRDbNjy92y31WWJ/sSM/pMwbS640meX/ref1u92lZMalDJYT+jAiiT3
8e8UA/DJLbk5KiW6XZzxiE5Ti20F5M7sIJULuDJ3ZrsBME1oUX86MDPAR7dq
UGcAalIqfDryI2P+MM0bxQst4OrCKqCL4+w0W6leojCr0/K1mykZDn76p1/2
rC28rFdetod6nE2n4WgLyMZlmUhOUQaddN0e9R+hdnIylh39rVHtoOmJIZ67
pDWwrn7PhMXBb42P4IhqO9Fct+a//IWCrLDCTO0SeQLlhO4h4ZyhZTOcLnSm
7wJV7B1hAPfhO3QMtKWaJlX6Kyc1XDEywytf+BXMXbvqP1lbnvEKa/EI+i8g
617i9EctmCpum9vnel8efC7Ms9m35jJgf8DYDmhp4WDYCXbmqoLeuIzrJt5J
rCL8SGsYvxXU7sAFvYEv2sEErF8ANJLaPO/lA9AgMH3nNuHYrch3+tj9deTE
nNAD32wg4DAiWI2IThc74JfJ4t9QDpjzm8KzQ0K8pgR3ktmc+739cgnbmqlR
1JbMsvpaDayL8/pNpvwJF/EqkfmnIfibNXcCjPXQQR3biQKFZDd9EIiiyUZu
4BR5vJ2Rv21nurWWSduXcXQVfNbZWX2bb67M5qxGAONqagwkfousXM/3qm2E
h81GiziGgqsR6n9WNu1FWDgeiK1Pe50pGsKdmzvpC4IOb/wiWSoSPpqmGN2f
X055m9q0KDNgsZkpsHPQeQvX2ZPwtJCtivSzfF3XN1wWJqSQCXWS8aKbQVSE
aYxtfXQEGpLw0sV4XADtVaLpPENaInYtB0PiFLoeMHkAQDVa4HanXzB0knfO
6sSvTSUaCAU1M9Vi4qJic47mVhaH7Kb9rJhMTu6RfUJGjrWPbUTNgApi44ih
5YEOW191FOfNXqFIjXinre9LNWyjQ3BbFtQaHTyTn1h2Iw5+oadWr26M5g1Y
JOmM5T7YO9+828xIPzJLAIpY0M+FRrv8ZkaYnjjpULRfMd9CqOg81g7l3Q07
vH0KIUHqM6XmJVfTeINtecu5oDpBQe/LegfJalOr6FNmsnEvt6JAiQA12sC+
ntvHRmZOuUPErx6BkdGnS6McSd4F+OoKot/S3cvPbaANnqnJJLvVTDl5RSgG
jV+6XFAaM10M+jefhjK+dffbInRXzJ2d5pqR4XeWPlDOs9b/UZAwFNBHsTKo
mzbrqGDmXNAoycK3GHlDPlUeAt67+MHoyyeh/jVil+XhLYCI9HtFqvKA2SQM
lMeYPaARFiuwugDw98/qc5UST+B2QR49aSVYhWXmPwCnQruiRecc2D+A36A3
tUqT+NR7DFSWoaCic5d+IozJqOtIgxcKhfmDwS4qQls83zsZ+NNUB+E5TnyJ
8O+C5HC9HL4H9OI5H0v1qwmdqqBA93mN0GT2fIlKk/Yzk8vzcSTIcew4Qje0
/qTTSsgkrt4kR9KSX87Ni0Oo3IL4CrGUfCkWelP2kviCVKNH/4pv2cYAWw3Q
m4IGfJDMoa6cpxWsDdLDubayzRTvdAYpqH8k+sfvR2MRAuLf9RjalXcPznJK
xcWYlIOWlKHWT1ZOhGELjlAIc7Yc7b+/v4Az6P4NSkajD99hMeLOz1lCXpy6
AGxfhH/e7ox5grCykgSw7OR8Ral6AeMLM8bVbhbRkeeQoEJPjLInBKz6LTL1
PBDqvFH81KViRdV2Gyetg3ABtUE+9DkFEy0Hrh/q6GWIgwaEn8rFhHxXKIU+
ryjJBZZUv+xwiEwxGz5B7jBRjAT04dGRif1Zm79TwQyP4yS1GYxAxM0UvO0j
oXIL5IiOksAduj5WrnoiZVy2kJcf+ddy8u2duxH5IXsrH0lqs4+XCREO3j23
DbSoZafGd6F1bN/ndUBLdr3O2Q+0ub9319Nn1g2kNY2NOgqkXuiSMdvvagh1
Qd8Vc6WRHTkzCfwwUgJIq4cXMtjyWpA+8w6nS0XgnmZz+DcdmTZab6zEPnYK
MVjq34t6hTJeIGry50JYYwUC5kKY8JsoVPKxreds3JicEzP6IBpWQGfx+v+X
GrpB/kQ2EcuXUsJQFZc8RluqInlg05DoxrIVkEJicRbwbsTpNeXIz8Agx9fY
ylwsSnhCghk5ra4FH/qteOnWlWS+BmPYX3CL/1+PUpZpWKa/KqvWn2nCqG55
cb7Yx7VWV8scn6wNuLQVNFBbMUN5JpD4fCEyGacHIlxSSdPyaps8tlpEq5Yz
Nyo2pivSG3Md18clScLJVhzF+YP57XxKXZ1wE5qZc9eLV5lzWE6u+N6ysUE8
wzUZ9Ha9mEXRWTVnua7USKtmjcSTy0e/L4ynmnLBRm9VFQlLNWnhHL44+uSp
P4dV3wnkOkRI6nIqcVd7kbuP25RXWb3KUD5UP0vdrqGiiUtC3fYInTV18h42
NIgXLIDrPW53/6wwe9JJDelSMBsM/g5DkUtI3dCSYUBPPZ4kQ5pFRY06lhk2
v4ISNnpnzqpTtFiE3P1+KFwRQzamk2oknyoiPsa3twa1zCL9Vdb4tja+RxQx
0Al8SM+h444PimsJcrZG6qZgxbLLDXYP2YH+P/h44oFWBsQC4f8tPFhY0Kp+
OgAgqorgX7hakKY49WQS3FVh06vIyI1lcwWPZO0PqaJ9EkXc0BcNJ7oLR1wb
+DrrH5x4mF+BXb9Ly7VPYbeLufqJRRYGbAnISYFFrRpEoj7HGiEbXjVHTUQ0
C9eLlVcayu3MtZ/jHuDtviluI+9Tfj6euvM9Sxcs+SelSEdpYPbUqmyBa42h
h2IyDHi2vCDi1dORNqyavH3ow/UB4F5iMZonX+XLKUsCOnHMsPoiSKepzSFF
ymr/W5K2et/MkHz9LiwbYiwpiOX1rF/YczJ9fefjZpSgkReQWeOgYA/2htM3
QCOI5+JenWuW/RLGo27ZgzUhu/L7+o5t6hAHaj7qjTl7tBHtj6n6Wr1iI6RX
iGyz4sIBk2z1qkbWl6QE01LzMoNIesfC7fh74zxncUkTuYPHWekjNYgMDVAC
8km1Fo0aDQSfcdyprNs0XvgtKrO0rHmFc+VR7jqlliYX83P7TWRvxHGuzWGB
Jm9ahmC6wgzIsIsrQg/160k5LMQiggQPILqwSIR5xFFFWH1MLeCAd6mI1lgF
wUc9H6ahVKs7QQgmfMQMyxA5EqXYrKnyyC8h5wj3Wn9mt1QIqch4EcXhfV3n
3z5K6YOBnnSAjnWdAXm49L4LxAjFYOVcGb8jrnERL8JzCDCQw0tIfIFbKAks
gpbiXt0H+H1VKFPtcR54YyyJkkvMVF2uzmIjD64bL0slskh58QLIo9qSrdWU
XuFN/EzZCjmQDM7s404rIFUOMxFj9cjW6+gLYuQoNlDzscp489bPYUtZdgXB
oVZKOgbqiwNrsXTHnFi+VwThAqeNMzArZl7IEJIJGPXEbL4O/9b4M+bm6E9F
glDzidcbsRNn0Mcn5P9ENQltW6Pu+BJVUWtKfyT073Z1dlhXI7QVWzSfWLS5
uriiH2cA5JNR70iCDEGQXwAX8doQcQw4DqMqT9NB3Wu0YBSqPc0863bBXsD5
vqqmWH/zYV3Y74EbiAeKhbEh0yUdT6t+AWDo3dbdH1AcGeWChbQOgrbW1fRc
Y0SxncE7lUVJUDROGIhwpAw2MMAzhYNw2G/0r89BjRAqkKn2dPCWvWa9+4vj
wctsj4IDwPIZAwbybPXigIvFw0lgXBIY9ytkUgrUuf5VGJE9YrBxmT+WqU0b
o+SY4qL3Bt+2D59ecrTcWzQ4bZDBaJxqp/hdX8epvtuF0cCajRZ7LqarJgwL
ZKVC6K7vExhbiJ6qQGldedAQBiwwIZYBCmBfk9SUUm3u7SxX6i8jbcXPuTwZ
CeJSxGEd0WVBSvQNao+EElTN4tTgTzKRr0KMead75LrC/O0A4gbrv4/Njgk7
1Q4CVTKeKJm6Xg+VB3pLve8/9gZafI+1rTtPHfYRGkBUPdqFezN9U2Wa3mnx
Uqo4lxUDwuM/hgc0k7EF1F4Jb+jKYhxxLJt7uiuTbowM85P7Bt9EDcdfQJAT
H+KUIkBnWQ0Xal86N8TECpt4D2D1cNP68G356QZAFWvmSMVWR1pJLT7KzKlT
wZF/adUqps2x88pYvRu63MSVXDyDtm8gpngZmNM3pSHTqQROfe4BG1uceCzG
CkaRPFgAoPhnQX/hoGcdc7nNxMOujTQJ9jn/fz2Cv9I6ioPl0icXPCAynzGx
2c5sT2NOhy1iCMUEqjEwfLX+78rWoUOKbm/QX/3C1ikyJZvtufmywSlCqChO
X8Z8xb5nCxiE/XK5bhCtlHTGX4hj/joiEzfg97v6dmXEaYtW0yRf25wUOCMG
jXxb019f2fbMyhZmylnnpKRTp6Lqi50ZUlph19CYnr24Z/t3aHQLXJcltCsV
El04h2OgV7m5lTX0u6g4HwhrKd8SFmdXZotWOdI82HS2jlTf2KYjJWlA3k/5
tmZfL1p6or4kmKUQLxmOA4j7oBmHTyZ1hX4Jb2GCkgyhW0Qx+b9bqz4rri/w
r6yFTjHp6Cm4Vf+iQoq432QyKHDV2gdElROOO5kjoktQUkIWwTMLY4q/F/jR
AU7oWdr1VTysYX3iWqGeQqc23VDR5M8eNGZ7SUQlVxe9IOGb0QyGALYGNeOB
xnNFtarsFMLVCamBjiAyrjm6GTrPSTDQz0Ha4a+OYBWZhDYmc7hCQy20/YEl
MgeYIEvw1zrll3xX3pSuRvG9aaKoYjFx7Yv/Ibokf/s1hj6MlgVdI4EkYCAM
vHzUVnnX/JlHam9uutYNJQ9lYQpst2M5r0QRDdCLUv57DzdZrsSxxyyaD0rJ
VzQr3EyX7HFJS82c6qr90kExCEeFSEf6x4TORqw0U7E0k5XFqiTYUTnNNcQH
rXW+V3X5sLcEKSQpkFd/+iF1Vfm5OCTQOGY2pXgdHd7tRGq5Zk4fZ/1EZ4Dn
eMRbCge5OaE9CpRKGivwpLewR5pIAMkHFWQLP5rk0WUmvgDr/V+3NzW3B0+A
JYk8mjaLNQPmoctkb5N44pZ0+/K91PQASKRWKlJcWJz0E4mskBvNKDDZ2LzZ
yKWQi76cohp/u710pHpk0v0joqkyoK2GoNtFNRjhy3Wm8HBIriVrCpqf3ldY
7QSYaaY+ud5QmMFhhh7iQNycPElajTC9WUqD7hIK6YzSR7t9PmBsNPaQ5GTG
cT7L2bH1JXMN7bRpwZHkpXom5ZEX7E9Tz0YO9sSx4PBYjWfKgABgJW+PP+iF
B/Yca3LUm8wZczw3A3Zmtq3MxT2PN0VVQTn5yv5cxllbvKsZQTA06lyOSAIn
dS9RHbvSYVwC+uFPxEgc0uQyLkaX33pVipO6uq+DLPhICBYWVZnMa82kes/9
Fx4hrNZXM5OuiEGm5jjVbNB+SpoFYivu1+vr/9j/4dvK0pjkIFgCI4la/j2+
haP7PZrDQ8Fj2bdDEX0Ru7jdFYDK9aCouPixS9ivXRE5+hoR/NI4p73s9HYW
SB7I/ggNVG43C7oYJ/gLkI30EnraNfsGwhTqg6gAsUcc7iUnXXrqmUqNXUVI
p884gm9g9pBNqI5DQPr4MJbJ36G5TSLwSnPzOMB2brElnc3xFqt9w4wLNpCl
1W8DXhio4HuaKCGz+r4Cmvvau8h1qdgC5t6Y2lSvNGw+g6HcHR6xnBEidn5b
zuaI/fmCahl4Fi2l70ruVHW4ukh1L0GZww7aBldnAX/QRKgP2Wy+je60vVYH
AcOG0Q2jJzkVETCqW7vFekkLs2m0PHpOUZ+m3tTZ78MN4OGhYE9m8bWBGNNu
thqnqttZf2vu3IzoNrAw8OFpShZebvdVR0TCdkr16qrVvdHmR7JjBzbB3zTD
YKFFaFMRxZkda+KgjPk5VHjfE4JTb15mIgrFHIlSn6Qizk4AA/qETAE/OdA8
3YWStsX9H3wUDTCmNW64FWvzyRiZ9tyLIhiHgNNdt/BrkrIIvfMqmM/MVgPR
rXfXysDU89oPjdNWwqfYo25PgXjeV6yv/ILeBt4h5bJLWuvOWWXrs/VY04jX
n+N53KHbv/AmPaxX3HiwlFI15f0WlN+vOGL1nU8RU2Tx+bP2T7P6/6RO95xL
uasYdKm2bdY8rzScb9lNZWNurEgr2hTSks3t2qnBi6VZ3rQ31JN/sjx1HwF9
EIpdMLPXiejwZ7yFSmp5zhZVf71VnJJ66vXYZ7ca0s1hFb5sKz6jVH7DZwU8
IVzjPjzeYjh0OtmJkBSWYfOEB4z5iry0Rn6dNEa3g4Ru+41u7u6lGmIRPrIq
T4kKGMkFECBc7VnO2zpGC5Z1bnhSy8Y0IJacdDdMsnlLc8IyH+MTNj6JusO9
461aRYLjuxdusPLWwFgY5FxCrzZBbZf2H++uqHn2zRxDVhbtcINdBS1AnZCS
+fshYD6LBTxcc2AT1/Tip98vwhsVMF/kz69fYpN9q/NvuMvM0OoSZgH2uwfa
Zg9MUau5ymXuI0wE9jsUZIbwCxVPlJqLdbUY3wlHkUYvmkxB2fI+0lz2nsAo
R+A4jl2syZsKdDpWrx/d+42b8OJj8Tsy9A6ZMStdveEnKJr1T/EKC4o85XQ0
sOCvmT3fRyPFda4U5Wf5E7NjtPb5iMvsD6vzbDBRf2MIj3719WdG0se8I0rw
xkPiHP/JCoAfnDOfts+JP+lDH7YK6FTIYud4YkPzaQi8xAlteaCnH1jyLZpb
Dpba1mEUZYln8O/9GEZRIGMGAl4MYr03PNnOAhNo4K78vjfOXrxO0YDOvWXY
CEQJbyHFDzAUGnM5SafX9rbsOS/BOVRQCICLDxDfeGw5aTSMGxVnS5UTuxfu
adjA7QDJw/VlsRDSnLRj8dzAQhnOhvyyNA6PsgazNu66LUPwIDda4z1MhaVd
ghAQI0JulAmISKPMfZAvURkaZyvUs5OxZGteijTViuVI/dPUkRdVH668EVJc
pVs+t4mTwgtaXhJqxuD00VQy2MUB5kzCUufE0uFyXa9MO+FdwaUXVXSsjXJ8
6ieFAdBjIJ2/hl2RCb7AuCg2GEq3LLgh6qg+7Dw4zmTjSrfTrBdRG7crECX1
7zMj59TSu8ifLxpAVfSYonc0UkyJRhteldTL9lU9bUfUf+B7b1q485vy4rAl
xwyZjm8GQ1dLRZWH+1SPlIk5Ky3uAvnUKU++7OjxsGMLvQ+AkK7driPYcpaa
cDs0NJGCmdq6hltupTGOCsJLzIRc1LmV7ZRU4udiH1k8u9J08TIgf96khgGY
YM36DOeHHA8szageKd9vakJqwOWyn7gj0ykgpDLXWV0g6bQ6aBgbPxfxSiuN
2ogbONQbab84SJ7SPV1Jakkwe5jEZjbHZ1rJX9Bzpr5823UJQaoOSLzBdicR
TmD1cuKQU28SRZ/n3ReSrxGJiw2M2lt9yAvnEZUvPxSvvqC3SbZc8hmerN6m
c1KUL2d/k8KLNYwXB6UIlcGX6jcw+bkt+BlUQf292DWmRvkXicQ2glccZhmH
0afClHOOcGyawnJfE3I67RXARimLuHOFCixbmrCFgUqjLfijuE6yTJoO0wkJ
seIhURE1YwKZckUaKWKWjq7d8p5CTODLLdRbI5kN0UVCdg75zSuzw1GOTJP1
ATW8xbjrpggsB39wtR7BGD0NScrnG99U0Q/hPFTHfFPW8hk8u0eV3D2MGtVP
PiSOT6ZMGDsp3BdJByPmEAzNPGs6bICeJexXAaPwnpHBzY0p5NB52xMEZF3N
jLrFbzadZQ8JhT++KN3As0/4AFRZEE+kV+43/0DmDoEr5IeMX0YT/LqH3yeT
6ZpDzcmeyC4S2G0S0KcS/uy7YGghPP36nMfUvDcB7jkkN642Ch2gmMZZWhi2
/kxUYyfcO48846xbIcTFQmU8cPStc4NM7wN9cQ35ZP3bOUhYoi7fqlF/VoNi
bTp6/gmoLrydgk7uj9ZC5J4B+amBbKQuX6IBf0cgw4vhrGMFVR3sbLGgK6mk
wXaf95Gh7OeWHS2fsMH2wo8/6VzzsIkkilosz40ExtYjIa8pSxFr0Yw27VwU
RPDJfIWXMnFZ6UYPpb7FsA5hzL9oNjv8DV9ObHAXkV/fLFDsvMpPdlLmi3He
s5twE9dlRyJR7yPvzdshMzOp/qjreropo37DV+lHcWRfKrrDmAgl8rHGY/d0
5NYjbnk7EKTBzSOz/0D2U0sjDZXPtUWVHeIyG3VoGBA/JTBDzwMtJbBYK1nV
vEf13cIG2JyrSFJeSsIoJnvUfs9iYIPxbVS6xtpV1oSOq2kkjRbTbYa80e1F
UV7xRRbqWygNY4SKkSLgm0Rq1KgUibrG26R4IcfCTBpwMaVj1LIpchyQzasJ
j7lv6IkuUQZNytp7MsSGwaeFerYCoW1y2TLsUNCkzs8PF5n7JrOnDs0YtwR5
kbANnzZFUeWOyVXm2b9KAN4WSBQRTeS9WD//6CIY7D0hOrWwSL8xnsluAgSg
L4I8jLYKedm0UnOQ1b2UbZDHa7mHUXWea+NBdYFRDHODQKNYpsDP0vutkvmr
H+bFeEXpY97ZCanJF54wsCb0gBhpfGB0oDt7ATTK5JO4hozAupTXm9wkUJFY
Ts7rXMSJMf+z8nXtZaREdhbBqeSuNo76oc3vtFSAj2ENRb/UhpyAo4+Q2k7c
kEf7I6vyxzb3wudo1WCn1u1MWY/gtNnzQ7VhVXtFCT0924d8kucVKtZIDzRx
GPH7cJpn9gSqRVx4iLv/3tiJC3NrnAACx3mQfXZU5pAl9tra2urBIn2pEjYF
QSquFdStpx1lMs7fw3C/wee6EKZu2oaIk/gFebxQP202bEOCGnNviR8Qmm4a
TdYEkjDIEjSBb5qo81IF9vbdjV47RSx88tijOHA28gaFX+Nfwfq8CXKpYWv9
457OQLK1BBLNMwcC9VmjK2/AmJtGdGIkCbhyNUN/rQWvcPic1Te0pIvQN7Xz
RJwNBRSl2TsYghPdvg8DNksz29DMcling+Z7MwRX3ZjUOedsvzn/ifXC6DZN
7MudggllEUyqK6p3V87D/QFRU/qVqCkH4GR/t+iFbIkSQXyBIurMVleGfoMr
zNXrRGF/zwgBuJyoX6Dwjbdz2NDWJiofgN2fjrBhhQB5M6yYmExwWGEHbNfm
3uEiBSPLYTanYJS5BlOL+BJ1IVZf1m39/+D+NGjulhvSmmcFvBVLIN2Nmh+B
e9IpSjgu2D3lpUamaJKSnsGv3fO6ZOPbUd2cxoy7vYE5gywleOz5O9UO5MCu
xMsiv0BgjPnGb4sIhfnN7OyOVL+rakHqgalnm/EDAmquo7bngxhlyzuaxdAi
cU6HNaWnm25MXpTz5JKMPSFt86tIQZXK7W6t2i4fDr7i0Upoo6kLbWfX73LK
Wpnupppv5WqHYX6eRxUrCi+CINDhU9L59RtnDAK3maGPjYzfwuGhz+2qxXbe
41TTm/3pX81Dpg/gT7aJxGgEMdrsQItSINrGZcoHEkmZcVNee1Wo6vHi8ku8
Ey68Lss1JaXRJG3+T5f0Ah6L5K+bu8Foo/2VUmU/au0m5p446C/QDNd3mtK4
czZx9gtz3v7MO9ZATfeGLNMwucm05GamYWhPiswd+wp3Lwp3vMamitrOMogX
++K9x1KuyfUzyO7IN8gbvapfv1wHwLjbR9qEBiLeNxFziuxffZx7uM3qPcvg
ihgMvgRa1R/PwfBD02T97Rj60ykQr720LMtlMrEnx/9SZ9KIXrBqNjxWXiop
iSVvkg0IG0ItSBubgyK53REEOT2DF138IlBZj6Lz2HKaZIFltRubC9cE8gIE
T6W7hYmGHccG51rh/16CM5QmXRh0UyUQX0CwaMd7UWcIeDY1XUqpS0/tcsch
yvZFGi9AbTqpzzWE1JSK55LkrEJn3C/+FQEmHp18QEGeJtJJfU4ueQ2SJyhi
3LzezQVk4tFRmAg82d0kJM3DDZFnh+ks4M5BXYtoAOhjONzZc/RqsaP9XgDT
n0+7AHykGmUwUjaj7VyFn0dYHSLoy5Wm4Og88Cf7lUrFnlGVYNf08+Y7RzKw
nYjvH7A9lPb57OUUOcBkPNn3KW/tUCx19mPzdLvM1jjzWM0rioIkv8YugAwI
dc9VuesnjOhpeFeUBM0FJWz54BGjRam45W4GGwcuM4jsK8dKk9roUT1VsM1d
FAiMjQ6G3wTgToAvQcSMvaBQOGSaxM8rO4bydfU3ngiQBd4HpRQYZ46i1UlG
wFFyYDTHm1GRoV0FbDSp0vCTn441W/kgc2sFaa1wjpOm1LKaZn6h0fpQ24SG
gW+5p2yssEtlfAxCsJqBWU+gqeT/cZrGY8RcQscg0tkC+qZ9WDNruT4UOKhw
pO/84uqXiOCqPv2sioHmjaE2QTfhb4pPPnHyGRSmgn7jV+kcXRN2E+4j/WOD
U7qGc7A/Gw7ONw0y9Ck5jneBkoWOGi0Wlz4nKmuVDfj/rbLqoTU/sDPMZf9/
yFYXVio4OOgJmuPpNiBdJbbikWlYjUVUGX9/1xf/vUJnG3pWB70FHS7dOQ0+
IvIdsTC2spQRDo6FTlB8fjqIczsnsUha3rZ1i9W3diwkUPELDTCjBbMwulrC
qIEe/uHDe6iQPj081ZZwfiaq+PStk2xAM557eEtdK3sgDx5m7V9Ow6DWdm+S
s+0ziKhRVuJWrjurOVXrml+J9VkSLoI/DkuIMKYn5fKqtqU+j2cbAtBZ71qM
q1wP5LDigSBjQUg8W1D8YN1XvN6OnI82atTG/wFg77BLkHGhHumnxKggj0m9
s100Wknbt5PDUDnbLOGJsfI5BOkbUaIDNu9zLsrLbANNh2xXEL2sEX2LCqUQ
nIt5UnRudgz+0P15UunA/hRoQDSHR06MuVc/Zf3Li52hj8uXPEYoeahV/OsA
3Y0xCTeHYLaqBJbnFU/l7pj93H5ZriZzHJZF22wA3hY9R36lLiMzFTmfpqzH
FXpfdEAfLdlgNY+5VnDqWyM6kE7XdAp6XquOd5g3n1g9D7pt9Rj3WGh8iXvh
213u90o5hR2pbRzlUnI9gohAqamo2WJuvY3+5vZugoCGUeabKkYRd/U84JyE
/xTM4T3h8rk5ztqcKAiiFxv1OyhpT/Z55eL17TTdOOFHEoKbkP50Tg/F8aOz
0fiGChTLIibW+6fSi5FbLexEkYqlrypDYv11JiSEYignA2BB/Kc98H2LuzgL
4ufDTlXUBOv0INs5hWrIknlMJlz6gNlHFtakSZ0JU8msYhuDoFjOr3nUldj5
TwEaNQsHb1GKEo/qlB+B3TknkNxTyz/XGmI7vfAIFyZOhep81x4Prc7bkoGT
/uBrT5ExA6Wnh2RCYp8h8TBsfYUowlz2sNWFL6yt9VAitnhX0QFhZru0juKh
I/qJfkSEZjpMhhIb6vmvvEnqt3IfTlpOouxLlrOPV35d0xQv0UZjsLB9yH02
uM1SwfBgeEOKWt/QIdtgqMoMZFw4BHJFI+sSlD1y9xjT0HyASsMnZGw92dOq
BggJBn6XX3EQYD3DpAw9gx6S1g7iGFIkBG1KpdCc5A/QZKYA/nhJ0JZklPR5
Hd0uQqktajD8LoZr3Q879H3PJ0vIn5SFLCcigb/28Px8bh+eyE/hnhbjOOEv
uuWlb08ytULbicEV0lwUtuvaPbBdjLaJkh2UpQHe8ZFwmkqKL9sLc0MIZOo9
KqQO5cwc2DKvSLi9V7CLJuy1Qfvb/IbMNUT1RgmbGuKwdbhtix905JcfqrGw
5CGAHtZq4lQj2FGA44gvYltZmZHvd2o0XCC4B00xkTJsROBUePc4OAE67Tbb
1Q/FWjrzBtEVFbXhCZUp6hpQMp8g/3w/jZL01jTDcmK/EQKlzjesMQt7F61k
un6M74rVMk/0sHUQzJhwn+Goy5i5W8Sx0l+paTp3u6e4Co7VmlS8+o8cPstW
cTkWFHIpxDedxjVcFeag3gGWkvSLzlA4PQWOMr9rXONG8vKuBiNsojPgXJ8L
bbvfAxPkPGXui9a7oOKh3jEH/Biiz9W0n5es5Vp2/vt7DVTG7Bv9l3XxxmbZ
XLLUXai+kASJ6SfdNKNLrKmejylLUjr7dg8vlANEmDwfknytweyGNY0wKbZ3
FSwsUt30QzzJacKA0lYyyvveDcfflSTuqhdEg2koL9smxwE5sOiEQc6+9Ksi
aD9zEAe2z9t9zEV+kCXa1MgMpg6dm53fi8i7hY3Yha8Tmqin3BCitbii5PM3
8RacU9aRZm8YXS8w+BiF9kKsJRLdvtq6+BSYqnzoZEt5go6XH4SJnW/sjXK/
yU8hDh/ior8t/j0g6eOI3lc+B8aNL38mH48C7Ot/xazczmbtGNiBgCZ57v1f
MiqUz9pXvmlgWeiS5cWnjXokyv7iQ9FE4SoQRfmVUg5YswhDsm1w/JiZyu0P
kcBC8F9fC15tHQmcrjbkJfz7X74IHUtEd4AfGUrSZ674HqnPi/amTYqDkZN8
04cIhMQ/ePaAavzyEgd55WU5Q2Hc2PugnU5bSmz+EVusYyNabDu6EB4GaPpA
hKyXGNkR/CaTbzWopp/2CmpAX0XiaVRjoDOo8nJSj+5AoN66VG5nrgqNelIL
heS1Ta/xQic9tsXDayhmIZvjSwMpXqAea/nD69H/PXrQhQhk8kq2Ns5f2LEP
allqjs2L4S1Y43vCeJl0CqEXYQSIUlV+YI7jkHL1+Uod/EqBElv81oL7wG1c
wFNi0myC5GuRCGsKZET+fNTiEZSinpCDP0k14+RP3f1185kn1Vq3Wi2M3gsH
CsMogJDqxC6FrXlBfh2Uu068Rt4KQ0qyA50q5AYGkNxVe+rfKKSZZLALRluZ
FtUobpvDV4lDIYwfXfBkrtIGGJ9b5I7qa/iAjSu2hK7Qk3XjmUCctcHCIRPG
eAeiAKh+4dNejO7hTym9I1ZZ0gKnTwuZUM7v1rv+Cp5x0M/w7Di8DomQRNl3
SZL+CiDgNajQcPkHIcg7CvHeG+ExC/psoIUzFeW9OMUhgu7BUH7EE+78JDT6
hKDKKGdS/MPoDf90gUpMwiEJ8XV3JN8vc97iMj/OFt5ZOE/yk6Uc/SDpN8KQ
x3Np2mbMfpyEzMepkKtArfPX62jmLzZliyakz8LV6HpCaroC6Qj7T10UHhUT
quJ9k2HHMU9rqxbfeafo8Ph8rVPrTaAV4CZtUmuJjrpjFrrKeFiy+cryBTKW
tZCLGszYzuPFPzYIw9KHrzhlOtAzSwFSkGXzOdG/WANXsJJkVQphtd0RnNUP
M+GYfqacIQ3dZ9SmS2zRGC6KUrN0WgWfrzka7pBiS9OtbjujrBA/DB6g71JM
cDwI3yfFL+6wX4ElCrNSa9vxjXNpIO64M0YUCE7UF788HO1ZVAdmJmcViNx2
gwpwEvelvziI73AbYFCpy6wuKWQRj76wGRtSKta0d1ueo9xrVXeieHZEKau/
KTa+qpJjZBhNsxpkkCP+UwadVFK6B+IGR/gpMByAbaynq9h/kWGcEng61yX5
Fo3z/3FaWgkiHjtvRgCWqmHWGUUxRPalaCLx5/NqFboJqCMo4lbG+WK5jh8H
ELkMJjB8lRBxrL6RuAhUsE0K/OC9dQp5b445mBimeXUzPp7k4P8NWm3QzgfH
OL/v4YA4QDsybhMJ285Sq93vSbUod0iI1lxoTygmOAGCqKq7T9CPI2LECXt+
JeCRo57k0tR6TnuC4gWKxW47ud1YWFPyqagg7gSgpXDrgbZR32AeE49+b2SA
w4qpHjPg1dWqdlEHMfp9n6FTkDfGs+7ROG9/Yfeyn8tT3tHJRnsn1aJczAsV
DaJFHhNxyhiLuKVe9gErS940MHuaG4jriMQV1c/UK5zKR/D/xevJKtptBerO
xEflEbmdV0JdKEjXMmRyhNvg0MQpsu2ToeAvTEt1RVyj8/ZzNlvDm2DdOiRE
ZyYAZvlKm9GessTtCK2YwNCkeQa07wlaxGoKEqev9iomTeoarz5ru4gBucQ9
SZqpSa7FakLSzuUecJU9K92H/Hb1R0TR7g3bR/Ii1BeRPsBKd0mYCLRPMSpY
M+RceBTT9OD+O4qGSq2uSrrCEV0iKHAKRsVYv0MmLUSpplzn4TARYoajmKkk
fxV8M69Kn6kcraIb82UAIfXp9tQBPvnMfZEuguxQlOBwfbAruDDpubIEi643
k/weDc0F+Eq8H796hj+W6jrW0EggT6Ip2OeyVG2FLMzGHobQAjPktQdWthsv
gdo1fx+aZIdcPF5MWVFuWQB9xeb/eGsTc1vAbegNhuJ6DzXvvS6b0tHYDPPr
IKsllUlreTFffSxRn1gFsR8exoCDHTV170+ULlAwLvNh9OW2VSvv6g41K9fZ
yncIXvbw3FPXpH5RlAgtT896BunUSHXx5SK9MMpOYbpVOcNDPeKQXoiSJSOu
BVyjWa1OreE77E8SINsT0Cn5Bt4KZU/f85ONrGT6IX+HADFZ+/cu1GacVds4
a4NjXB/uqBE/ac99w5+54aDu5TphWGJHzgCIq+zZwnSRDWhnveMR6EGZ2u3G
xwORYvL6h8LeKEnDB3fkTGwwFRm8HUqAWZ6IwqMqbFsE+O6AQT6EeSXsx2Cy
VMjBsQSLWDymrnM9TQMWL1Rv/yevyNK/NTqDUr/AfQ3NRfqbKW1wbyhnmeci
vpwMptu1mJZcKQ9830UAZmHs0aB/rEjxafqkjRaYGkUMp8LPYZZpotXdGEww
p5EkuwJ/VgCtNuQCbAEKjKXNCVej/pWreUq0q6JvoYnJNwy/fbI9+hrsrq89
MzABdIqOsz9GVuDBRMWEH0LQy5ACQzju2Z3utFAEDF50WUvifQwBd2SKcLJ5
7vn7EayOfFFOGt7Dqm9oa9EOQSS37yMl5A5NSWvDMZljT17ogF0VPgCDowyQ
aZP8pDsbkImqgKydu5wJ/h3/ZEvUaulcwT84xY6le/QHzV2piOg63XrftQ7u
g00kZyR6OxagmNrorCv3HkyKaVj3zryhkkpcObaHDB4Bbg7v4H9wPg1pcDPC
3e2qg+iWk5YoflbpYwe3VOZggknpV/o9asRY1KQ8A7/PB0BGVaRBBchcXWQL
6InTIvAh6FHI5M5RqlaanqXSg5LH5dypCXgsZScWOXuPaDPvR8ZExxcnfAaA
q0k4PYcSP6/fs8aEILWRSPrtcOIExIBwGprD54bL9u5Ihq2NjNa8BZHphlvg
YrFaEoSl9eifjhU/ugBYQFrrlMr8rvYsrqO8tHmfDs4qws4xqxq17mN7zuXv
8Mr34aNcsXzzdcVyN8EvP4toN1YYpuDVwMqOa+Re3WT22usJeFzrI3ZWwpps
BVFAgC7j/M92eiyRb96YOhobjGdSV3yvNy4yOGCeXrCF/FJ5ZUXBCPo/V1Tu
4+YZH33Rl536K4AfsyGGiynyLpBD68eAuLxXGJlgoF+EBw33QlSbWtpwZ9N3
f2eaMgVEycne6FWkDWQAOMOmfUwajCrHmJvmBYSP4g2pcyTxo948r6ODyg+T
ytdm1dxbfN3dP8rUV91nFTsP1B7ltXXivhc2ol+oNOx73CwNay8mP/DRdioR
Qg+dF8rrbnDV0BKHtT+6X8M7s2NJ6ItCtP0hj2qeAKHlDAca73muAOD/+GJz
k4OUUJOnRvvdlKECaSUsBdfXAumtgmA7n4MBpNkYBe+iDM+5JZbBG2HOn3dc
afdVTSDNw1sEugQbGZsYkE3P3XB/Xw3kuSd3Jiw3Q3vFKnsb3kBkM+9wJZQD
SHhCPgzQHPOOJmZImhXfntt/Lt0EEx+Mc0BOs3wDoRl8/85uWAh530tR8q2r
yqFKumh04/Ezp9RwaTz04Ff7AAqymtNdaS9sWduf+jEsLXTG0u4srN2UCwNr
w0Vc3QZq2IfBud4m9ho2tbm1w//fUdqszHfTl+Exq1dm5gNmnzggylv/9gpN
BGW+bglfS3Jb+XoZnPv/Ry6LrNOpBmlNwZaT7MWwZC+FMRA9414yB+c8NmB4
aVRHnbLGqQRzOuiNhmuS3utzaITWpbTDf+uZHWxh78rdKrS/lHeHSiT1eDm1
aH6oL6NDIw0rqO6/JOFOozklpkCaPtoXhhoN329cmDkx55Mmcg9fnOuIp0NO
CbaeNiRjKQAvJm14+jGbuBmTCkW3ctm9EQ4EfR6qQH/gB4tggFDKJF8Zi2qN
kIHRx+2kBVmAlkTO2+KYQfv5sQ+5UM31nzMpzceYUIRohhNOCiwQHlpR0zVT
bb6k3L/t2Djubgti7ekrzssSvna5QyaquMZduTbIF3WjGtP+lXfI4NbBYfCk
5qwbq4xc0K7+CFtnqznkeAKdww+fn0aYPKlFo9EjSRTfhi7hwiWAUpxfIhdF
d0lnnSZdXKrXgDjz0Ox05Zvr+bKlH4OIf1sshjA0tEs5oDuxv3Q2aPSWx5+8
GulbHk8vnzRpuVWNbU2hENvkLBAbx7u7Ru5IH8ryOQ5Lt8zE9MGVyeVCTKxR
uhupVSpmYP4fQviyfz4ytBfThhXXXq3ZOLBXJ5ptEzxJawV7tXbxIvyvjScb
O2jJXa+NGCSbH0oBMopXAZzdlCaQdArh7TpCfJ5p6HMbLU2XjjDFxlYh43o2
k5S7fRnWabEb1LCfeVs4k4Az3tpKQfMtRRGVuwjIklHVbrRyoJbixp4ymU/X
yAIPFR1afg+swrCHYk5Co2M9jDyuzUYRqQi65NgTBWQwnm/IO3vvaxj5S/Ax
Nuh0dzyBBmjNGK7pRqQwKDcoOmhcIe5ENNTCNgfcGszA564+sWe58+cABATf
gYsIqoF4JJfUcgpTvA1jgsaFRlOVPwG32zp6+gz/z3nMULCmhBCshuX6scbK
BJ4Vy6+m7YEQtSlk0UQySvvI8CzQV2ksnkCrF4bMqcPPqhaix/TOYDw3RVsN
Oyk3L986a/+NVD25QDC+jjzwvRg4fCZEhQVJQFE5C9ULQkj0sIK0eiqU7+pU
Bpkt5rozX81udvnjBEoLkIl3IDuKk4s6CuC4IlYsttZIWOtAbDWAydg/JwsY
yKw+UU1+X7l2MZ3VE5tmrxggxnWnzMrsid+LJQbiHdqS9k3FTpP0bvF7Vxag
Oxr8WmPa4GGQvxsDtFGLphTH4iV8Myh/VG1L6oJUr9gVeypLJdn9VZwkWKXH
rFgkFWMsbFSVq3e40XtpTGMedEZKEIWa6FkSY07b75ZRZDZWeXnV05fn38/x
ZKzuxgpERNfswmc4v3CP/aTyToP91nLHq42hObx7GC933k419X/GYj47qAu8
/8JnoMnXBpiVrQJnWhNIOzOhT156b+T7MCgG2indmLZnlQu/0a61t5k891k5
aXXUA6XDd06vhHK07KcOcwVbKbLu+dXLgSgf/BtZlK28ymOfbIOokmBXPAaP
H3pweqmUcZUJBc2Edfv5oP3Oh9zYB7MUf70QS/xHQcFvKImsEIOvvqrcZFCx
W8fC7EozFUgmeJ7XqVDpJy6evilTxJSaeKx42AwUvwRkIMJG/cVJBMdjYktw
eoBHjHlaJANXAl/msExZ/PkBGPJMhqdHnTdozQ85RMdi9uZOSvQzvWr1f+99
2xuoU10mVy4+GSMGRcy6AVWBEbLLKnjGVLviMt3QwCpPBfE38870TyHbNSYs
HCMLvs8sBqPi9Wezp+bB7BgtVetonHotlLTj9nAS64ueaV1hW1HXu4y9HnY/
bAnwxe0mUfikC2siZjxz2N2CUNYWUFDQAQGBV94w7DqMYk6qZXcQDixfWbb8
B/8dYRIxviw+b5rBG5AiFj3hNHPcLPzkSYFmFcCtjLk2Ykl3BFkWw73BVITc
1XPW47eh5OnY0670YuHPs/kQi+PfTr741gG15oBoFh0+ZBXv4heWBLKRWkGf
fXiKe/ZUeq6t2c2nHGNA1ETaF7AzHugvtZPxjCJ9mVzHGKlB2NK8vSdQnAoC
iA0Lub5Zhz7CfeDAlOh/NLYILFYXKne+8CsOYrHAE4HXBsIAlZaEpOJDbNA2
/ObHmHCKf+RavRo0YWRmvVPkGIWmnRXkL+kd3zR0TuYqNa7cF0C4jiRTPpeK
ETHiMDk/LIzI9df3q0U/beQnoQLwHIZ4D9ggESUj6QTavlG6sRQL/q5mBmcs
NtxU4XDnrT19qZdWwpViH4+mPbZvAS2RG9I1V7kZkY8nKr/ApWLTZHH6PK/P
rLsILrWPdL43v0V6Qyi5zcfhZ1my48C4WoQIR7OvDq/HubxKmmy/2K3Di8Ju
G1S/jhj3Hawvjod934WB3H8x+o59v5oc+K2Y7+bFaitrJ/eEUbQHwFp4ivey
Vc3Y1qhrOj4waDVopgcJlQOzBT/qNECeJgIpZlVVnhgnh+yJTaI2Kk6ACIDM
jGyOtUcj9KtSgfNzPjGwaMD+ohqXP0fS83Ng4q0uOmsahJtEsmXKMhgXcGpF
gd7wFBbEtOk2iEGnykr5zhG/rTcPuqtxdsVapTNVATdgMY9WSt82OmbvkYsm
Zd5kq6YUnq1KeNM+JXFxcXmKQ8lfUL4IPjQ4yrRZjyKeVd0odasJ2Fi9hec5
zIXbhvPD2bQ76qEbzdIWPpR6PYEClfIaCYNtJgkyaYWLtd+Yw/zFwp2zPduC
gmAmnvQHjDzIbZjWBCEgDoHIJPuMxVON4WcZjx/n8Es2ZwfaRH7PG9bjrV/c
fomWCx0RYeSxm+O/zMjhgCRw1Qb7PW+r7SjntcuUObhF/1lXcsnzcZu2I7BK
0qNjhBXpzhWzMfJK4Zo2eVt5mP2MYYWMNxtjLSubqCHKXys4PUFYXuBJZlPu
wUw3u3bGBfxiFelNtfF+RomqQ9lfGPgrfY7ryLW81yhzWgj/lXrNY+lGzh8b
wsrtMxYCbyIxv8hSnfZWAQWore7ZQ9QhJhp0RGsa1HWL2niVIjwoiQ7u0/hv
iAWRbrDJ6LRg7iirvrDtOMEczNoJZZZrkB2TEHomsEeJHsoBKyN7hXK80gmO
0W6qFC6p7xnOIVLTuubtKrR5AwQrrX/JpLwK7fNmoNibf8wtD0A9cRJ0WjN5
zHZOeT8oJV8aNxL8WHlxrlguTW93kKoJeScEGanavLlfIMQ4qxs+5ir2qP0J
4vguQRTllBoFA3vA7ZijUuGwBII72rYoSO8LbBLzYbzE5PrimyWfxrmil3K+
Dqp02A8kIdL6vZZ/2buSGEtgiHSkNeF1P6Oi1jyu6Ozug1ozZFSaHhKIWPj5
vnZ+6+f6QVW0/G+LBPL8Lg1isLMzfK/eeDWDHpcE1aJLg0/yWE3RPVYgCGsR
EHmOYtRCMblzcjZgtPXyT5USujQKTAOj1hoLwEboDMYysS7mv5jm3yS1cT4u
saRfY91SWW7mcXxKD+ACKu0rLNypcHoRutP2P74fOJKr0Dzl4O+tIXIUgXH8
lPWW/8uD1RM9QiyVoiYKkUwX77F5NgUSQBgUDFMwHrES+6pGR6wmOVEDxbpC
Z6eWYWZXH3Bmu7I3nCUYLJpPC7Q1di7LUpIHgBGuxeuLiOFcsB5eD+bHkvAM
+FTyfm0QXGsK3Kpz+TXQejnYpzTQ8O3N+uhfFtDszHgAda4hOKVYdUKLpcQV
5OhENl3nqR3kXfTqMKUIdw208af8NwNwl2uPJi15fIENEUVTLIKbLQiSvq8s
G8ClOg8tRQ6LNyExSc9MsIEFIZfRSNN/hahf3fi37UsM0OqtH5cw9vBDrnb4
CNV+8MFWHnEf3MhNLI3ngEHuqKfwoCFV6ZUlWdNJTpuiNKqZ9Kil3PZncABH
mjr/E/1zpa8+UITCL+W4rrm7o6Ep2/miT976jUbEoMaMN91mg5w1VgWPTJur
YXgffFcoTRWZQIBLoxMBC0i9UrrYb7NDAWNcye9PKXZEMasTj1z0irriYyAQ
xhroJklBPrAuzQG3UDfxIuw3ksM3eewPR4MbNx4Af+7A0+Jv2iehtfSZtjXB
wP0YNg4r90G8Mn/olfBEHK7F4yzixsnLA3Y/RE0Kq1QuiKe5e1PYmJjNXI6Z
sw59SgbQeKhcN31r4sgue42Kh2WhcrphyhjyKl+Gq4sGgckp2I9ikB6Wg9P1
JK6LI4qdyrVH8T+MAS6GVa2v9buv23Mbqv1cq0Ns7kIPzkfP5nz69HFBE1mR
T68WUwnLOo+U6KoYDLPriyR7OWUDNxybRvGDOhU8Q9Fq/1pkZ6txxIoTukQb
Pt2tyGXl4ZWz444gEPn93Ca69ZqCpH986JhT49RNmFcz0kYRJYh6yYagC+Y1
PquQIaqOJ/shaKj/bzywl7hVbRd2DMrDaEKvvmIpksxmb8dV+Uq4C1hqb/VP
pFWYar4ioB7FtbG+90U2TwcvnpJaHPDRPFS3vBgQ9aoGTetbvr2Yz4m+4oIC
rH3U1KCOe2atRnDawhZfN7tPPKKZrgxZ0EtuXDEjt8OaWVny4qpknravcwej
klU4BUdwwBZS60FghA895ZsiexluYOFbrfPFVaMclwHdPNZYy2F12magiD0E
C8eJuNA2okSEG04WGDt+Wna3MN8cO50nm63VeMGR+jod4bKYIgvNvmmC6Kr/
myDIrW9Kx5RiFIWzQx9IqFqAaOlt65a1KMEa29vqXvBqS5/rnQe0LUxfCTOe
5uyRwjt2DmrWon2r7sq/GdeChq0UFu84ZL1vlv7kXmSagv7J8qRfuDEcnrai
YlqkBHnJ9hGGxlXfWd8prwszpxpLaYYE4SeUZd/lKZdjnmGGtdrjVfsJuEdG
2dGkt5EKZJPzUpXvOrWl6Vu8gR5kosy5GODYZobQ/NQLp2igBEgTOEBt2LN3
sQXmFLA9PhEDWdQPvh00XAO89MI/55kvJb1rL6j3IbfJk8TeBDIa0U7elq1w
1aWHJO8hUj3Q4c9vH4mSjIZv2BFkvoeNnbUigW3yaIhrboN0R+jaX93vdtnu
1xZxJFuVC8N9sa1MkXQMSCEkNE0VRqiFCQJ8YCuKkDjefGf5aNNaPe7NQ4So
IfKNfskxPBqR/SHEwk56cxgFFHrCgsXM+CgcFicmJzBZe7BSTK2AJocyxZQl
BK/7ADN/bnlVO8meBGhFoJy9dczGliIJBygEZERIGZ+BYXYeGZGkIvpKcXdL
VydYuAdX6DveToqk7rQw24T0A0TOGW0c0tJjYVi0iJNjm2nw5cNVfJYHRsU6
7Gbfv1bUu4RCfKQ1tpMu5p0S+9k8ZW1Y/feWQZgiMJ3PCC6aOfKhys1+GDPA
ScYs/RTLSx8Xn7iOlXr8aYn6a5eeeP5CGrl2rNCZOXUP2iCUuSyT2W4SgxZj
3gzRFxyAHh8irAR9qJJA4QVMc8X12zuI3FzRqXE7CGoO8dRe0qnGCMo1zsFS
a7VMXTVTYFTF+TdiHI1jw595XXyJQnDrWeTME0IC2/Ji2zCxDW5xt2wepd/D
E9QYY38ANlVbj45A1w2gFTre8RSiGH0+gc0D/V1UTpKHJOp7dK/6YLDtvveQ
4+AkNX1fv+1OfVafrHv+ITbM/qDn6u58XI02tYgJIQcuj450OyvHRbuO3ur/
8ptLEypZvBBeQTytCryjZStN5sHZpFDUC2bbYk4qOrm6qiIwtdDB/5pgHA1K
eVe+N9RQkYe/hKW80/O1jrN/2e7ZGRRW2FNkKrzP9X9TxxGxyuK9Az0ybAot
I9PliPiGU0SrRj+ZKKAAlc/wil0GEeyxvQE7xvT5qX/VJxiH3VdA40eKfI3x
EYPafKPJID8ZQPw65WuIMPdjDJXowjpGwVAEXhfFugzLPhLzTYWOPdTPMdmN
wOftiWBEbaPMAfMp3q/utcepOYQ+aSnXMaN3we5J9CluiyJZtQjevkZW6U9N
5I47m5cQpuDk4lvTBw+oN0IKayC82VfxKIfIX9qlvZpoljrlZIhfTvk6rZSQ
lWWw16m/071weWf9MqkdwD/kwaWzw8WH4UPQyQF6T0zJmrOdUCr84A21DCdQ
JWH9LC10O8Zih3mJhEX4dvuGCM6dslzkg/bZ7PHrDMc0ELGyUrcGHfZSxaGI
fgFYLpKoCBDCAfEDzvwQPI2c4TIceoUVKySJOrQltBz607aDcgHm4lVAvL5P
9wDbFyn3aXVo+3zy+Q8dDYnWeFv6DXWKEMjnxt4CTT2gfGCEDUI2nVELh2TO
zHAnjRS59yZP8wqh6H2dmbELKQgA5WiIhbxwn9gNHSDK5ZQcCVbOo1KkrJHA
HBJszHVSzo2PeSL5mlI9nMizUD6Pji+P3+0HX0fc8BooVe2y6H7xeqfvRO1B
HDVHtLEuPfn6N6GDPkI3ubQIp+sedU+GNDL3HXxRzid4p82yviFJt9vyGOti
u8LV4xXVrL622/v795n/rqcX1GvkvIoF+jQhWK6yfCq/DQXF0ZVOSA3fj9K4
O57enLMj2Zav2ntIL4BC18UNATwTKlfv1feg+14W9gIq/N+oN+4stPIzNBDh
5lV+3rdtlwTkvmMcSJ/veO5SJpnOzn2cCrcD3dVzYsG2cIHUEV9Gk7otlSij
aEHohl5qn0Y8NKQb+lZ/EUNmFAPH8DDlnVnp8tHQW+iZrXLkVBmXIz3EMEwe
uYMVMIpkDku82c7OpH3KcwGGHaeYQURnsJzjhazrEzNXLBnECNSwiAisHaoX
6/zJBCnyRJfIC96zr+tuVLO8r8pB8m+gQHe7JgzBl3iK2WLAEj4nBjMJBtfv
ENjfHqdcpFkltsTmAiWYYrD/1XkExQ8MMvKhq09dhnfJEan1MKOB+PDYtnXY
63U5IubgkAw23nYLGHYmgVb88ahekwnln5wrvXvfaevNiDaz+XHAbRjz+jqt
j9ei1TWG+h8NDSpgj0Q/t4tl05TeNSoynPAw7LzlXn1ujSYZKNbsh2dVJE7A
pNbbyaffAsWJOOTOx8bI0UF2g5Wjk9Qb2ocP3VFrTl15IXxJ0OAi8fhgUSFa
oCE3xGvnMMcoBXaJ16Ppx0zxmvvIjsMSf1drsXVJZK55vN8ikCuiTDwkdhQt
abGyXA46PJ29W3Z24QzBzKQxKCKEm/4zVyVj91veRuxjoNwRsBigklE1IdSZ
QHuY2YA9CRhYTTinm29fuFKx7IoypgYhJHCPHAYRPVAf1xPomh6EsfyybeuB
wUL5HfGtzaVb6pYKp+q8Qconp27fL0GbJGVvZgxhWe4BPdoEm/OGWMebZR3l
Hg1E9ARDphZ3ambNgw0WgkoqKHgPBR6fsRS+1LvbbtXkp84+A6W2jnS5182K
SndXP/1kjdHw2tx/zBieUloVc03ha2g48CC3TXVumdmd6XZDQ44GK9IDfCr3
lnLGrEkJnEi21aZ1ml3cGa4UQX72oX8q7nYtkd29c67hl6YTXct174QamhgV
siLzGr3Z7Wry329rfBNR8jK5mrwrRTnVxpUbNfFyCRmu8+wep5DIx48fe+u8
ewIQ0dfTtbHFqgXgvveC11Nb2eEM20XYi2LcCQF65K5jCbpi5NjyEfjTcglR
loj+sPLxnwEpNJwMcDguMbZS9zzS+Hqt1YOImz63NDXqNtl9ZVa6PRAsR+R/
RTQuRM9IN4CIdAKB9zOaeOmEDKTOx/dfIshbyiKVUOhNklTG/nQGcttj44FQ
JkehKXFMDb9A6KQGZRPPhIq/IRzF552Fj0P9L41z86JLlhclCi0V+sVvB5OO
It3z14atR3rR8EMTvCQpaKEg3gaVEyocsWoh+6SC9WmAR85VDt3kI+QkC7Dt
dNQlP3chfjHx+BOULFF8JrhR6sKtAETzHcaX9O1sFy+syYA5fYxJ7e/CsMzD
UvMY64qxT6zClldbVmYfpdgtMC+z6hqJzdrjxdv5aB0iRyI7wCWel0Wgnjf4
Hs5ffY/yu3JeiQNBZ6cYSwkOhyrHK23C8xMJvxwSnWs3Q1I8tlrPRNjEzS+i
rFJ0CvrlXK1n1xhs602Rk0RztyOAxtFDpIaXOa0XPWChdnzRS+IouwDfdO8B
x4MjcUP05A/eMmgp3UNzW4gr3LWC5pCtcZC42zb3miP0ngdQHhbircj1T1V4
sVCunQ8chwfwU5RYnSlvv6ayoGFQkuwclBBCD5o+kpI1AhZj736OhduvC4p0
CkI5UBZFsM0lm1ce5VeEZd4kwCHyxOap3AfnzEQgoukqmLcL6CVIzo8Tb3/r
RSJi4oK7Sq9x4x8HOxAGSj6lPBth3RoS3nCyO3/Qe0oAYpStmvACBvJVzT0D
nMge8XueTzO4gLsKINj/8ztoxqMXYZ7TBT9ZihigNX/VnxjncpOqZ92SV02l
vULA1IyLKDOB0z6dxIhz/piZnAInbZipeQKs0z8Zc0il8VEOhiSlvoJ3JwgL
ahG/a9AoHMM/8KyjWGo1Rv8rrgoWWEL65ZdwHxpUCGbwniAvMkxiRG4sqrOg
fRCj75ocokbh9jfSo8R/wdnPcknPNoyde40yWQR8YOa9f9dk23G+TPeMqamG
dEG6AAFkU99U6qz1a2v7Ch0W6ttWq4XfLX0JlfwTWn10YtlJ8wUrEVrlDtkE
pS07T2sGiH2SbMKPmococ9Dr8MhOwSzDjnV1zjKvPPx1u9HX/SE2ecQdCvXC
Vl6aSIw7gvr2NsW42O+XoBZ124Z1e0n+LOloTYBXvTAMR5GvRDn3r8OLRLwn
e5MikTO1QYu0r1x0gZJ51YbEdAflhMNO/tsu7P/35okm7wjSV2uZ0qG2dybI
fdTJkBFq4zbMbAH+wtHeI/vCux7nSwXNXTFkT0DMcI3CfwRIABUSyU9pgDza
F2D2AUx0yToAsUFqRww/XrfDEhaoMv/p9ScNK/QkA8iwp7fgoHToErVtLqN5
e+FCMgC9WVFpbrIaVNwQNS9EmJV399cVGJwu+EqgRAkjWdzvVkt/gJJuzdlo
GreRXEP2YHJP+JkggFLVUgllCIewoHVTwebfVUQDc7hF4UniyqQZ7x0ZsyMA
cHTWd8uBWl0IJCqHXr6hFTikl7kitls4oWbUN7D+/g+9pt1s+Ct1rpIcHUSi
+l5WUZNQJZvAlUKuOCojUsEhROiIrVy70f1oz4wHGGlSwVEUTh6tpYA3pI+z
fXzaEVYVU8a5nJo8m/HZD+82mw/Z/HnLIF9cZSPmum0XBkvgTvB/Py392d2W
QZVWgva5EPXA5mDFUsFHMqrof6+kX5VTezKGEvxFuRdFiXhMX/YQpH02c3Qk
aMJh5pnWrqngZnHez5v+hu+mvosGaB69isblvQZmnhH3HlYGlZd26Tx3TW5z
/Ta7gKxCLHWywdK0jj5JTdaNVT/dD4d77YutW/KOyNeIYY/sALUTXZWvuLNg
ambQ+D9Ewvf9aFi9qqJFNaPYm/md99GXmBAoV4anGn9FOKW36Sf5TvdecszV
WSBkg4IZLl8NYH50ETXEmZgMjURQomHt460RHhpkZem16Na4XY6zyu5KpVOr
ap5bq9eBd3QSPHyQrAddOszSk47D1Dh0sgitZLKHzX5cT3OrV+4oLEIN8p4Q
J+fIR2pQBm1DQgUDdGNbxCe08sTqQjtn3UXG3huVgKzpuexKp2rkKt1U7Wz6
pQqDc5QLIMvvHmy6yXjmBzT8tunr+ASisMD5cUNsCXWkigtYsr5kgFgGi/gl
2kBU5zUp/sdihvvvcT6y3H1tWpz58TPy3VyRMwnlLT2nSh9Wpv7JWCwPMWf9
UlDhEjYOBBfpVdrOhOTRF74s+/gCvlo/9CpNxvm1K3mEMlGmQQ8v7sGCNxqS
WiU9wNdDWvYYfdLyu+YfM7/ePdlaAAejPLL2BeRuqpTZrskDWEa42JF35C4B
2+CJZCOAbF14v2SZLwNib7EuawSQwQPSUNe0cVwFj9fAZeJZH5evp/paSIYo
4QuzqyXyKsllWxV7XjoSJYzf+rj5B9V2m9h6ABaNXWfgj6MyXeX3dNq16C8b
12vU1cY3sT4B1gi9A0JCoW1nX2HmwxiA8EvzBILxU29qKwdeid7Yunagu3cl
Zcz26f/+Wo2QgfHtbkJLxmi5V3UPDHS8Y4Rn+die0zmtwtvue3TlWLpKSPj2
Ri7+AOdLFyWkSGkVOmms8uGAwJHESE786E+YZ/WLWsgahZXBrJrqjhle/Gd2
K8BZOQFBAMiEhKolmjgGp9x0dR1e98xovl/bm81/Zi4Qg23+hhjIzCvTngX6
WSzxJ08hqLvUs/XtgmtnHDKty3WWsB9nnZSAHjFGITbOHMVcT4frKGRFF+ZS
U5Fbe1eWhdGdXZpm+QGp4HBmiAT+b0dll35dcZ1yCRVWo6NGU10LyXEV9YXx
4kdHzreb/5rjtOJvyPy8i0cdfZjxWSCBoNnRTKmrsal0b4f4ZSrB2PmKJ0aq
izac/F44vGMhBQezdYcZwqMpjdX9tuxk2hBdZOLCTArlCW6ecvITKOW7P0Yo
SArn7Uw8lZU2Pa1aTLLBegS7rDK5lA4+M1w7BYYH0mouJgXZYEd+UK/FtN9x
F1pveQ4wncAqfmtt18MN3BHYSUzi1c8K/dX/jkqfOdI1RImVqEeSlZ1laznY
eu1GgyNWzMHMD0i+ONoV7GSHwD1W96tUho6TZhHp9XGYzxNXiCz+lplKaDIT
TAdZT5w3TdgHEq0DJB+iXBm53lYdNuq6NpoXZ0s/JBdafAmm6wTbZWbMncOP
lQhxBiGD80ORfgjYtMYXVwfCQwkSYykGQ+8l0+rub8v3n95Ikbe75HvT+/+P
aodqIFk3Kzrryx37ow9anuD+dHsTwfhxOqRKPneMyXH3jzCBTLRl1wuUB2hr
nUTZcxZDIEUesw7nDkC27tb1l+ZPQHVVIzAljyuZfBFXtDWtv8qPFJ667/rH
7F9Op/ln1qcocSidv0sMs9D94kVr6F4BxqH3/XnD5iAFhLvWLDyRVODcpTur
pnFxm61mkRdjyQSLUhBMikqmmdM6ECgtDBLDnb2NUYC51jahDnbs/Sr6UUJz
f9XpI3iN8lB1g+lg0GwWfrSyYscKtd5/++Xknt5G8RoRlaw/b9oMYIeBvdG5
x95z37qlMSxfLzCIszEDLuWZv1CBhIDEduNwdhwuhHAxOrQZMWr5NSDq7SK/
oTbsUFVmEdtuMvFdx3SDB5F1y9aYTD0pW3LFLceoSI8kglPnKWiOl1ZhsE6m
wJn2X6hxpKbz0RThBwD/OnEk1OJR91l5NCVqyo9lM6aITWUfI6+1BwZwzOCw
pf5WKi/KgggB7RXfy4Ni2bc9MeGFwSJHjsIyBVTkHKont8r81dnh9EY5b0dx
91y7w9HVM1wI+EtRpIsXkNBsqB/C/9di0LulMCBK+Xg5+mNBY0G52izA4wgN
YzqOejd4n0GYMF4tUlv8KMKzW0R7a1Jj1Mrw0huDyA7x1wAy3GlTthGKUFLH
E7UXpQOc2CzsLRQ8zxBmoEphDeUJMZ1Gfl/OxlM2MKxKhh8t7ldUnjIR9Xwr
+8hgFUC972bdR21xlJUKgGm60cbeJj3sRpDZGu65CTfA+w3q1J/jvOGBFZMw
1L+wMPqss8MUIY5HXiZMi6BmZ6KfvfYdkSQJD9MrKpSsUJn4zzoBYfgDNqBc
dL0v6cRKpobpOmBSakInmryL1S4JDbUjTqtffF/q+WqUxtp4SBRgunobwhdh
Pfyvn/Ydd+XVKvy5OXTh38Nn9LXEetVFtJPEx+L/iJSpUzUXjSkLFhtOEgP4
OD1/kZhtlBvJum0eNia6xnBvyT6an6zTk/MBQafccM4toPObPzT/BQJel0el
a4C4VMig4LZpyE2hFchCTK5GHBOxXhPI9hrPGK2ioXqmYyWdPHMkQikRUH/Z
d1m2qLLzfOOLshiHALvP62g44lGcwUa5eb+/8Mqaohh9MGsRTJBQmTT2PWpU
dtTABOvaxD4OIcM45vMYCK6lMv/8DVdm45uc1mOKWRHWd7NWQ71QBwlrY3Un
AXd6zjxAzbaSMixgCCuNV0sHIpIvISzxI58OD5Mmef+p4/mZb+nvFH/YSNGO
5VPvkNLEJhKcQwg0faj+2umGgbrGVrSD3GIhJ8Qep9TE8qsOSjAaqGp/TRJh
7MOwzX3tH62MM4DMd8nPDJxwI2IqCA6gjgJ9jaTkhIY5NzvAwI/hLImvqgMH
WBtZVkpdlPrvduQ6fKO5duf2SZmzQr/du6lGLcGX56Yn9Si/7yZ9MQG//IFO
ulc8muqB5nrfLlkGElh1ieg2g6azbEcvorR87h4uIO0pYfVMOEAaOxN5Vge9
4iLAA/jmfJe5ZU/ifsAZHKSa0+Dwp6Tt6nlPJIxJgag6gjWeBD8L/rY8ogzn
HgZEDeGpXYxbAAqv819oeaCSvq+gsDrStOzpXvhcIbKP8ejD+EV0R3HM3tjo
fozbOKI71REi0ImjdmBv8cOscqsdCcKK38oSYUuQUa6x1K0tVxcadNu/jm0c
p+m2n+ob9vG/9Fg+F5JGRACgpx2NO5ieTc6Vcx8P5Rx3M7HowepOgzCcv5fz
ty9zzVW2Xi/TzKAnoTyS7cxxTVtvkPOazYAsOojFban8imcPMjY46N2wpssO
/hgISqRONwN+gU9G6dGtg4GUmwCgfcYxBZxF3R01jtRQLquxITnMM/G+NnXC
1FLnp9sVsZLxoeKlKE4WdHZfNmqk5AUyFWrAfVV8ZybUOEuux9clOi85Ucv/
WsGlcpfkKCpxXEHpaVPRZqW+ZyN7sLj+Osd1CVtUg+hfOq9qzQEkXKnjbhkl
Mdcn7p3qoNklK1tpE/i6+x2ypbJb5v6w9k6PnKeK5oIBdzJxaUdXXSCqkeeh
wVHFlICuaJ+DrDUnyDbvW6N/90Iw3rrUfva7Kk9QwPDORsgj6fM+5mWiRlPU
NMqzFlRErSiLDXBVCUVLiVGiG44cpTBj5FAmBnDIsPfbK84IjZaSAlCPC0/l
3adMJBkTZCDJW+OUDxdOzW47fyjMiIVRFBFBakHpI1kL5B9/Zf70pJRycTd2
6Jl6Yrn7gDidtyrLLkndFew1dfoMKSsN0ACDx1gJoAwCU4bNdEtaXCxUuN++
HyKCeckCYdrG7nzzpfbv4L35IDWqc/cslUfu+SkVmIPyIhs5e8GWrxen/152
C9dbvipjqXL57MmVKz+U2wDxQzRw4eP90A95TNTr3f56/XKDQuymO6L8LGTL
Mz9/5pKxqGevV9xNfc/TWN1S/26c3IBHM3ON0mwQ7mRek2aEweQmyD270ept
woJhU93e9XIxRRRg9yRwFMSCKc61I/JiiYX1UqtZcTUflc4UX+LFzoxjsPd+
a8IJuozBlW0FQ8TgNmoH1F8OdCGuPQFaSB3xYWObjjd1d1mPS8Q9SFjGroN0
KkhlZ5j2iyjt0fV/0JTVW7KQntPFb7vuFZNPs/eECWGhK5r/EnZEj8mdQ57V
d1cmXDj+836QVqrP8h/ZZfgEztjZjlitTmRMjvUsNDAtutc3VYylKu9oEFbr
D6jiK/CB2uKb+kZW1FwG2SBS8yc28YkpZN+onrduECpb/m1B1H2M5eECWH88
abl02vssnKliK6kWoFK4zzUbL8KFtziFkwPQKQyLz3kpZ1VkDlAgEZZloBAF
usJrqDCtVgXYac/cOuz03ir90fqBdTq+iV7tLhk+/9i3VbqmJNF9wygq8uPS
clQKNU5D22Can1ntfPvtFZ5eKII2s0GzifcgNE/+oW5YLherKJvI2TP/femN
PyFIyVf/BDh6krivKF/MaUdMU+mB1CvX1A9Uoyeclrty67B/0f+88l8w+4x3
EzbUcMnlSH/nMdKURv88Lpll05oVM65nMNQfQ8aYJU81Qbw5zQtRy6faG59q
aaibNnlQuPSJEJVEYm/nuC4UwrocDTEpgZjGiY8+bN+lolNDR9B6dYK3nBSc
wimNBR8fXgP804O2O1q9EwhAR0r1iLx0T7nh0BmN2Vdxza0DK5EUbkFdSXDh
6Pe6YA6Y9YEVfBX8/NFWQCmVE3Xq8RiqZ3B1iDKF3tg0E+x0TmaRHxIIdxBk
ANt32I6pSVDIrURYUUN3G0DFdXgoZUj5FSqtcQFtAPmUSmU22dYh7GHfwb/B
JwrDpGP+aipRkufkQUl9AFdtlXa+O5PssUtxVG+S406+cl7Y8p3mfqe8fbwr
3AWPyfETUyjhdqZh3KvQ/41CGAfyDxrLDrjcXLGuaO+RzIu8Uuo2kNKxbl3t
5qpb+OwWVyotcaS3RRlXFwo2cw/2PidLt+HOQgK20euaFbBv81S7ouYGAfnK
Weqgn6O8vsmWNHFoZ7gAwBEGp+y8xb3/Sb/taFdn8raQHL5iPAFyY7O3TGSG
qdO91VXvWb1sHXwOgNbub/9eNQ+Bgg58PtIdIB37JhVj2Y7IfC7JZ7BXH4x9
IbuWzvKqUe6EQuMpYYB9r4RlG6ks+DHx7HYKlQGdhzfB+/eIZdIe2QBK0W+y
GnYe0oiR7athaU9HQYi3iO+XG7bb2+HoE7C8maf5pB4qw/NkmBJZBEeNA8mP
yuO8NjFeU/T/yrGnL9c1sbwymz3RMKlVlUjbsTK0pMHHgGFfJ3QpQbvtHCY4
VTE1nij5QpDoKPWvunREKqKoUQd711Px7Gr2nvxOAxQ+8N5WQXs23HJorOp0
hk6VJdzRRqCiyxMcXOQv3Y0l17RqZh8LqbcI4PgegkyVQOYgV1wK+3M6xg27
xZ7Xqcmb2rKZd5UyoJt4dDaJX9VdcSTZKyxt/mH5nbvYpmbDB73mM/WUyiHk
tvlHeEFh2DCWFjZB3nZU9K4CdqR29zThJejtUykJQ1Ell4Ly1j+u5ZjBj2AR
P5fwKZjMc4od2yKRk0A/jfBqvarojou/pea/aHZ2ozGiXjj/1DV81Wb0AJvO
1tDVhB17YF22EJoFyFZx5qPNf+zZ4ezr0htpwxtdOfA0Zg5zf35SD+TwuL8H
WgwkGUETj/WG2/zxz3aXwtd1SSSpc7q+iQNBXHliA7jCuw9mE8lO02pW8fF9
mxeOI2CD5HfYYciTpXwI3mJw1pa0N3LRjUukjNlDRmni+/xFOsmsGJCzVwuO
qq9czUiwDtDI//P/o6pOsur838Ba6T2blUR+s5ALFPXUkYtZ2nVo0L3gqopE
W6ORwDX73oTaLZUc55iivKSkvkNdkP6Qs6UThHfvPdo6jjNklZHTZB2tIKVX
AwOnFJsPwBz7zE+NjlmaYjQ4ZxGd1FBRVUYr3eI0KnBGzqPyrRIEwS/sceWf
5mGXZlhDCH5Hh2WVafyuOW1CWVC125/A+jqBwkxtWzI88gM2Mh2Ej7LNrvMO
Da5oMWxTLfdMiwQ9aRRRy0RUrBUShSGe6uTjmODsDdqMbaeE7KngtNBEzrZp
HOPTVc783x4X2miJwL49+tjXYn8L3rt2SdW9WSYFnR8SwU1BxQ58CPlJbsg7
5UHBX8EGSN1AqWKj3k32wGoNbFvru2BzQXXpKnxYo3IPriI3b2iP7/wC1S82
pFVnP7IB5A23uaq7DNc1mziOkq08WG+P2XCyHjwMDR3zaidlZsImSiP1+hu9
x1kgjuGFT2s8J7N1sFpfDngFxJf4fC/hnbLeEbl33DkXJ6r19gzJdqZJz9QJ
g0/5sE++pvjHBO0AyT9p1VZlsZBN3OYD2S4vtNc7FQjW9oPA2KW+qBEg9wpK
r+ULbgFEKbZ+0o/u7Sw8cmeYRcInaQ5IDDxlvQHbBh2JdvSfVEOfUaPvzduI
oCqb3UZycR0460Ofd8QSnglxBqMKMb3VzwhBprATPZCHibKyR4JgN4jrWUyp
LYxzmB3PwM9GmnByrlxvmrYolSiRrpC7Q3R/dafiEgUwcyE4Z5e7Po2OGaph
g18ItcG1sjcOGYx0vUmPJwmxESeGf3sOXmsS9vi71+9pIjJPrwTJpjoI3/3K
OvgyGewZ7CluUcQCt7HCdCPTuvyTKJ3r/X4ezYDHO639GJV+0kkIr+1r+wu1
sCMv7vtPCb3ohqrqOq+F730jtdbIU6vbLS71yf/Ff56jXfCXxbJgwDefGFo2
d+IP8gQ+7WTzotn2J7fuUQ53TatzN/9BV1fxwH0MgNK+SWhTyLUisEJkDVTI
lT5ZGgdPQxYuL6lbIprG6IslB94Zrl+sdwYMz5hciDi7VwOyBCMqN+yQkvH3
4OtbzNoSghjgqp/7Xrz8TMQcTy8Tzb/iSBWGEJOUB4rjLF3gJh8eNOryHnse
wNghGGYgbyEMf1E+IxRuaOKXqPqk1f5mF5Mjm5oA3t2YPogM7Iu7VKxq51Kl
hrVWJ0WC7Rmz9YXHKpBETboSpRsuqpIEP9Dnfmasy9s06M1MIHPwwDf1u1HX
vT//NjMvn+U164rT/sJJpxzcvPd1c5xaUiYNAsnnYQXOzREdFtuIcUh98R40
NMhl394qjZRBy4imVUKib9H43S7UQCQgHzbJPaeIDDbCCpteDhT/72SKfYu5
jxtW3oYHO7+KM7YnkNqC2ZUoq2o5qOU7gO2LMoSKi3QbQ0wltKy87H7Umyi7
JyCNlJzBjv/wzQKp4Y2Uj5ttRYWfhhzilG5F45mrvU9rbNjhKYS3rJwsqBQu
e8JrEkGy++jEkqtPLpRzeiM/WqZ/SIKN36uEbyWhe/A/twvfEtNBYU5pYUMs
GXr5Udn7Or8RwOSWHhUaQXDdWTSY32pwH0vwTyUW/pkn+52XJznIxENcw1/H
TGJPeEnobN0LtBHYFeD+POYS3PrvRl/hZ3TkPX7iUON6c6Cf7lNFuAQcC47x
VKO4fhy4Blb1gnwJixu5ge9LO/14/SylkIbJ+jjEeprTCoVfDvepR4vZriyJ
stw1QrbUY/HeYlD72WWPSnoGLJukA9lL8vnQY31EWPzbU08jirvnrxWhDtHV
jznvXUiZE+YUi6vQ+tk8fPyiaN5vt1lfxn+up+vhZTt0U591JD1KM94jPpOQ
Gav2XDg1YWJckCSBGpTBdulDqxIq1T2d8Yd7bv79hbyh+3SFHO7EUKy+Br1S
RWYro5WvZmLdaXig/DyZkkjX7ibBJcBvshypyllISWSWSN07zTLgtzrAq8Ks
qItuDLFYgIcGGJTkSs1siojdm8MqjELPrJPU6YPezm3bZGb70d+D9hctT6m9
MCdGZpg4Gg5eoxVy0Gft1kxg7ekW6jkETKcFGfjY5Ut1lcYYISJtTeYbtUcS
jo03A0vfqNu6z8qSpIBWaQvaZXOH5zf6CjiRsfdyyhklJuGwezAHORWPxX3/
ZxzxeyMR/aN6oDE/txkyppXwSmqcT2efOQukfFBwacXLKCKfa3DebjoFWXz3
W3nE45p9L5FtoyuACCXmz42QIEWmVzy3fag/PUyfRreCzfbEwPmRm0mKq4RG
aiPDoDkHfgiPAm8x9Err7LoXg/OxxGAW6S9FyNoHozPgWD+QV285rWp2QrEp
ZpOx7MC1qxAgF1yX8I+0Vfiot5t6jHoBMYkpXffXLeUWKthOQDO9qxC5Plfa
vitW1S3VIntbntFkUq5Os2JF/N9x0RsIe06sT3uuc9kGnm3Dp2HEVYvZP+Fw
OB0Ee1PUakbfpWSBHyOgIxhQUQm2D/eGZ7IbJpcUqP5D1D6n2RuLUy6xwFdX
4vtSqWBVmN1LOx9MNEDl03Go5w4uUlz+4z3SxnmBmkojII424DTtUoY3sVqC
BIN5LufMI+LIUjEdD/VRPwgULgXwjKq8gftTR6vy+FTtt1RgnaYc6n3BncC5
RhOVGqMCxE3gDOxSphlPy67Qa9ARZbowPoKRLfdJUBYUltmLZvo0VrdlqyiP
CMlySVm8TuSTVbCHKzr2OnA5wrrojnEpn6P/4b6jawL9dYw4OegD73NlzYCr
D0q1AiLLBCgc5ujDCac4HC/CS/W6/49IGfPc4b6NU8mmZrtPXUBBShsr8SqZ
DYP1HDyLX7miQyCAgds8Oke6Y8+g88da1Fujjqj18JuFUDPpIni5Mw6CshX7
VIJUtlZIVdN+Ra8v7wSk7Qc7uFBzjgptSuqX5M1BCxCgb8MPvPkNUzWpzniS
mu9tXnMa9DYhp5VNc/dwBah74JlXZhj+PpFbFJpffOOUrLQYiR+Q1otJkEO6
c6LLYbYcu6bK4BmAKWbbxdKaJXXcjSALXVRrf+0EkexjobFB7HO03c8Q1pFl
eJ4cQ+hhoBwxRFIRwwimQ8kpYZw5pPRWetLpXDbxO5iAOJQjCFWTkggR8wYa
H4/N74ECDf0vIss99ndp5NMvHo8PqPc/quqN+Dacvd9/4j1JLFz5JjkQFgGd
zE+lhSxL05T4kygX6DxVoICEgHyrLqImJLbT0IqKeodzW6eNCV2jsZcUg6uU
HWOUXDrQOTAmvvRVwOQm1GAsdgXJR//yYCuSwsLPDgA0xFmw7aRWOQooXXN9
5KXLdfYPOcyUHr3OVp5By38ImVKM/JIkuHX683AGfpfxiCDJGQzNcfhHKaX5
L363uf/U74IAMttjUZzj10FKdKYILRoozzyc1M77d0ytGC8TkVFHU7wYIZi6
CPKFi/jjyuMqlDb7nRTjeWb356oWMy+HV0LJ9uSUOcYzZFcmPDkAl4G2xCvZ
C1defHE5pC2UWM0oH1y/vR8k+JjR56DGe/+Wln+cFdUxadyfAaqFzsqU2RHZ
B3UNfSn8OxviHymtheMX+cbKPnTMdlkDUJqHMyXqQCgkpD1K4LHRdE2ZI4lW
u8ClYg2X0GeHT9JIT9ZVpVds32LkccXl4ChxggfwoU5TvIjhNz9dhFcM9ycx
tzAUV1HEQGj5oAO9BRoJLrCACBhRKh/6ZF8JuGEuffFC/FsMw0A1KRC2HZej
J9T+Hzx7AJOXxRh/zPyRJD5QCgqqVZnSRAZq0nwzItJ2v1IMg48iJhVxnV+e
BV2rHEdQZfEWiBEa671NhgtmtauW1Qi7bUnUQS2Tbgw3/tvS2P3UdiwYdFWS
fiQFTx+8vnoWmLMI8lPfKYYo41BQSHI+fj70TKpKeDdkqqVSqeDTAFF7lbWn
IYLv8WmyAzj//1tAsTRHdCn23dQqvC6R5sA52G44otdY1sEz9CFzvK7ZL2VJ
A7yG2xKgzEn5GMUXvMSS2fb+Zm86VWZpr1mw5kwGFnUhOjlaa0h0ONDCJNdK
jsbLTKtGWyZi8kd8KcekYlNGuPftZMko68tBm/sWoi6Mh0Pc5t7RWXY3ME7c
e1hghooHlj52f8SNkR3JOVhl7QeSenCBR26aqOaceFu/sCnPdwCvviPmxInq
x+a/ts2LUkt5ZgNgktVsl/c4krTgXBbh+HokRKzxLl6l8qzja7qguydy7aex
DgAjsk84gC0l3CWNDwnQYzCCL+cFlebSijM7pyWuQaMJ3nnjDtR698n7SVmn
f1qhesk4V0IJNTFIvWCzoSDz+Sv5mTDeC6B92p7wh8OlC63XaPBzH7qPm/BK
OTvDN+VU4ysrO/NxzG8o+b+C5L3oPvZB5kX8PRMSCQhgOucVYJ34NsdFU3v8
jA+sabU7ZwZBCH0FibEJf4QaNsbSvowK7qtHnYEyBwUStaUFsOouZBtsXz19
lK9zuv8+Ca4xYfyV7TUfdcfTUZpKb0O7EaGYnTnMP4wLMdBNAyp9AaEpZ2GZ
BqUBykrSevgc1xNqbt97fYsExJrQApHtISITy0zwhFk0Lvnco8VQ4HVz3+/U
SnI372B0Uw33Kl8zvLTwEQNueYWb5Dxqnq52jvjD14NhR/k+LhB9bxcty1vt
XRzGxMF+CQNOEq4eDXTc7ZhHwZFfFFeRjmOV8zfJhnKFbUzrCA7FuwTiu0Ew
6xtHey2beGKz4Tl/YvOBqBy84JLOYTWCqjqG3vrnV045LA+emEPTg2+AakXq
cx4/Vk1zOTtvm985IogePitxSpp6N4gcALsalt7cUsZNiR1EzSHxTJvqgvQj
4HQHTeT4wsdzeBPUPbT4EthhqJsnJozz5f1eDt4Dqd00VsDxBoAPf+21JPM3
fnvzauYRBTAaTvBhb4+dpE+zcxeq/GAb79Ydbw6+dwOs5aVzJ8rgIKLD3Ci3
0JWni28k4f5vl87JXdH17dZPU6ApK+N7LM0FX0m83qP4cbALSP+b4at7jXAP
Ro7e/ksbtpQqpVB7TdqcIalrI4+OgQXmLTOwGHse6xMpXFzyM0kaZRgdwE5c
q0c3NX6vbf1yN0GWzlziKJXQux/QU6BjBi1bnx1TmtJR82Qsx9/7+33V0NTd
a2Pd8EAlCPb2Uvm6KSwt6gVXiiTrlV+/C9yHOh7dCcx3oLSbQKergBUaF6N+
rqgoMhoBvgFx7KCkG+rOmG1+1kJdGxu0QzId1of1TZIGHWlrdODo6Fta5ewH
yGltFv1DqLo5PCW4AcxUrS9bPhR28rxzhJKvfomA1W5SdCv2dAVcZ0u7aUKm
oDtW/RyWoHv3C4W490Abx2By3BtF8bVtGTXji4/HfgkX3V9/4/Y6tzsWTx/E
ZhJdp3WgfDBf9ItE3WbH1om5jU7fiwvGry0HdbAs3nmepgITfsNitoID1dLc
xYu6Z171v55A32LRrzy9pLGsUnFw44HD6DKrIVnUB1P8GLbDLYw6N7oAQfG5
Y7bEOnXyoi9kDhKf6/nCgl2I1LJi7qsFkSRxC8svZ1+SJuEl/lFk1fRiTyE+
q7piVcTtVrZGpQ4bPoTfqXy55bx3a38MS36HWe8HSm6K6kfq1Tpj4A5D6PHz
RX9zuYYlLMmlbAyMbbma0PPol1axPtBpFf1luKvABwnH1EWP7K9Do8K4uLQB
jTXnFvlsvDY6iU4AI0x1yCkyTIxsaCnxdkhP9rhGWaOvM2/R8wAy7K3+x5tp
49BsQVgwkm46+QvORJW8ZvCGoRxqzE4hOiH9uf1xPJzpmBYU7eCyUXntdG4g
RrkgqQEb6UWnRt4j+cV4wdmMoWuER8UOQJd+cJV3vBB5c8ic4IPd/PRp/zJN
hbLgmkumE/IS/E4rE+mc+DKeA7+Yz/MNYQica7Ws6fv+9a+MI6Of6QMt9u0Q
w/f+qn1A66ds/RQ2YIARZt4Br05x3xPwz3SEahy9WFJ7kJBHE1+Ms99cp8wb
djbWMEzUZ5ClerJyGwoSUZmHlQvM/dtrzVoKnI1V9IuphVYhmkoA5kkYcVCL
QrPpTxpPCWLTltobuJ2/xNa1y0b+OE/C7epyZfBdYfC1v0eupOkOzgEEFDij
0VKyz1dTAkWGcy8t1TQIpopiqCBe7Gs+YPSTcN6goDrVMq3unRfzIbLxFN+R
9+90iKQETdJ/BERXvN5HTNIMrInN+LKr/Te6DMQnF+QHaPrEFab4OiWBi4zE
n9uvksjKa8FG8tDmQQHCRS6voj1IGWdc5wc/hOidPpd1IvvNDdp0mus0Q3Vo
kfqUKW6MkdYS4EVynvJQSXsu+2mTUdkhXUhDYTfyMgqIBg4ELO7jt+UNENx2
zLuUis+LjmgXSA/059AhOZAoxqi/3uRLnU4y29BVgcreLmwSyfjwaopInaC3
ErYSrqldVHKIf1rAkhyA9bWD1Hx1GtEXkgZzl9GH55Rt6eyKUXJjPJxW1okU
d5/K3dNFSrhDLt7oHuKdz8lWnehbeiAhO5Gp+UT/oMi8aNBdMQmv7joCXrZa
yJ34jgjBi/Vb2VVDSt9Fzr9X3gc5sozAPmAKDocX2MIAI2Q2T81jqkBUjmtL
DomCahV0yEejE55BWe6ZZ+3iGZuo11LfgRtZqteUp8hlABFGzonX5bO2n7+Q
zSHPMVc3QoPlcL0mWDKwv5nXpm3aGsoR8JcvAdqZkJKsheEUR0DmhRvZKhEu
AdMpt1YrhGBMc0W9p3DMX7kH9yno3brsVlmTnJfuny3BqX1dsK2t9mD8y2It
F3I5FDYTAS+C7T+4I5EGxe+ZLiADxKYX8BWFeff05XZort/7neggvl2HDua3
CUjGk1qY4VKsJsxRhl2qGhME/ZK7+uj4vM5mgrZvtMPQLjXEjlNAa2fRgQWR
xYBEDaIaB/aW5jG9SPDpeUthl1BiVCzqpPvamaULS2LAgTjDwsULxAS89WWo
HQccEyxLY+xBrOiTQgXKkUDM17WAYpdwGPoH54t95PJi/jisp5NGd4IUwoWS
F2qJ7JFjpd5R+1POQ5vYi4u5NOK91FszxMX4jWIUhBoCQNUBh3+nQMyrguz7
kmuL6FT2aFoeE86qvt195wUgD3AhXbFxmMiKg52Bu8mpkmA9LIdz7wwIP5b7
3OCD/1efi++FraEUusU1bTNdrs1ph0hwwc36OF0LJgx1rlge+qtQtdZnvGSM
/bV/KYD4XPeXvNWjAZZGU7gFRF+04FsTp3dw44dwjmGFqQ+a3w43qlfqlBA3
6mJwke1yygIc35QeXk7Bw4lSTjNASkhJMAqC8mPdLRteN17Dz5nL1JweRl1Q
Zk0ZdDYgv0mncnlzIOOiLbwvf1UY7x6Zip4lhNolZ1kodnOPxpAFUtDmSEmI
sevSLBODyAK+lFPfzZlSYgtjbYBhS5XlU0WTGW+Xs1qjIOxouwWPePmqij4o
1LemyhI4Rekiom3zT09xUBrH09bWrCM/QIqScOpW5lfVhkncvQ3IEBUORxSM
Xk39ME8ZiuJEe4NEWpZGpKjpvFuW/S801VFQCEnR/8hEjlvUbY6x2mIAG6cD
lNfK6uALOEK44ZN02Wo1ct5AkIMCZeP8ut3DU/EDTIEaPh4aeJMhYaLqvSbO
DD21AaamujujSs7sSnEHpEahLD5htJQfFy2PNMBMSx0xQvmOFWFmYFoNpVen
htsOMU3B9MJaBXFWak1OqkJ7kTipnQ4mQ9ishpwsOthJSSiBswJK7j0eLPVm
gbZ5HoH0rTHeTfy/5BwUBwRnTO0HrmrShbF/il7TYL7lmo3342Jlr/C+CvKv
dLgvZcKD+8oCVvFfxxr3qhe6XxwsKKuReX7e6jANVsamEJ/lq+AxChNXhi9e
xJfeZUODvCdWqxowQkaXxnLxAyJrRw2yuXZxn7xHpQg0bcqkaqzdWNeza51U
RbN08J9b2APuLwnnL1NgP6bDNeEEuM9mE/FJwKFtPLMPPnkvreQhXIMvbZZm
w9KYBZg09zecDMWMW2eeZOCljcu2vo5LRP9tVYOL7e6Vm+QDOYj2CWT9QG80
tNnMAd8TQY2fvGeur0lSxDBZaCtxVzAqQnhE2MxCfva2JW9NQo5bm8yPKCrM
sxHnRVOcpzpqlyW92o0eiekTwUTt1zgDFC6sltCvPlnXBGRn47aKKsC0g+Aa
DC4W3Eit6v1odAqOhOWumom4HL2+2OpGZcRSY+8/QlxrInP13opvhLpgYc38
3W5t2kweKwuICIOktR3HhIvM5lSUtYn5z11jEoaW3hPRYCDnFLoZuOxmN20K
JkG8kpyl7lC7OSbh3lVl5VF7SIyRoCj26zC73Cf1BrUxNLGDy76CVblPMpYX
D2UH/no1ZwGWrNCuqb2EOqzu1niH7gJ8MXlAua9Tvl5xgq8Q1wkPA+7R9IDi
cwAskw0DYOnes97b4RFg2Veiz4AnE/vC7hWmqxkxVm4gooVkoNRONmJt0QtQ
IvaOYGgZbRvioKnhQFXaG/kIH8J5khwF65NQ0ouZKOCLRu9Xw1i3H3YvddkL
7u0+4wOtAJNp+kSKePw11guFqAIoLUNB8mTKUH5s1QZvoTHOzAqnjuL2fdNN
0IRdmrBMc+Z+8Rdm8CPh3rLD1o/YhZX+jAhca9uC4zomyZy3jMnwnJAPY0eq
LLkj70nUAEHtznq4p6Eu8nR7CWC0sHSrUOEvSAHMf8zG7bS28Felkn0BLa4N
zq36+r7gq2+0AeCl1y9E8c96EXODqMTr7cBYKlR2G1su8GAEw2UpV3/+GfaP
vkDiwVg4440wa6vRuuZeCrQVQ7UqbsFSSv7rq7u7sEw9254UPGTqY1DFyZbY
Mz/berFz4kxyQCQb7iWR7JEjsqZUB/EEnIK/Jotjnm+wESWqZTuSw9vTwDf0
t55FXm6XGHMp6TFD4ihQpWqYRWY5DauOkxb8vrGLFC52SVCfnCLIuPgSsldq
edmae1XDdniSF3k1iYwEh6aNOdF/mMqOqS5mW5aYEwfwU4TP0LDE8/pbIZ7G
CoqR7C/lWtKP/9QHHEtNPKFJMjtV+xkoaTJxzndhtKII3Xqw4BXI8oE2w3eF
xV/nQX3LupXDXRU6TI0ViM8GQy82J+q4B9gwpFX/cM7Dkhl2AVOCZY79yMka
5t0MlpbPeNWcOQj89mVuNacmCJb7g8N1RPXiSrKTdF6JgMKmWIPJvfWhPUn0
Gsf/h3L9GotBWmHapD9ChZxscCBfEcE0PLQylFoBdvVXw7+Irr21/77SJiZ+
Pb+9VUR4c4rWNo1y9YdBsH9xGLcUYya7312hbiaR9dw6f3LLVZZMzbJgg5aw
a84y5IEeC3hDpelgWH7JwxsiiGY6ybHL4OTF99IbBw1FofwbFe86xCIdTvQY
Bf9gL2jxJaTJEbW0f8rSb1+ETsOV1CORKS2Mh2UAMm2Edm8gRLN80TeQop+z
CrfUfu4uAk6tLLzzZqOVhCMUSl/keN1F5bLpEDT0HmuaV6ZcMt9nlWQVSsNT
vvQhn0aGOH1oFSiq+3YSNgNi8xiioV+mwcZQuw5t3/xjaauMQrCxemFgRMKh
gFI8nlW+9RdWWmBeVTnPkWsrAGmqrgJmqx5axrsqVn1vSgYJgxk1MfMXAJp6
T1Uf6TxY88P7ZlX3tN4QTUsLpqWmyEQtMnROmDmFw3TpX24WmbIB76vOuMeH
pX3rjDN2UfVFwfe1gho0i8Gnj5hD0CSoIVQQGplx1JG6qJEmyQa5zMRzpI1W
YxaUcsfHMGa2ZiNCEwNml9GzzdC6wpySuK6zNc2wT2pIo511E4Ys3SkkBr9K
zszHm21WahQy2WpB/7JAR3yRTgfEFaoqzHYVIMt5zl6zA/J+ufN86SAqAnOG
b1RFcETpOdFEVz9n4yHSjclVkUvsyUaPFEHehZ728G+yU08V3SBt0otgn+qy
bSHU3UCUShvEjH2vNp/XdQvQDKWUUfIr1VoBQYrv8Ste0HvYGUfXfATvqs7f
dqS697RzyNAt25+EmsN67+6jUMhUYf1vQKuYvh3+51SdSIDHp9f6uyp8SYnj
fDHgfXgaKx9wDocDXTaUeS5PbnrMaWb0PJGIpsez9ol0Z/m6jtP9REaVAnOI
sIhQYcsKRzAGeCIdkBjYimws58YI9/dVUKpuS7DeyfNtAxwk3pbtQk2kVOo8
HMjvZnntTC7FnE5iHU6w3oSAfM07CMgPDohQBAPoalHiFp9KzyoEEDIV1bfk
uFPVYmDYMaRqk4LI7Byr9EtsqjErLTX4WJNBlfFnLsxLOZbAbvWeHEsCbmCb
Rg/Vqt/+Hcn+7r4/7wrOUfyoI2ESVI0/9SVyKFr1putytgkDNJsPFHSDZ4yr
VCbM1aDxB95LiLqtikbST+qrXUFDZWJSqkt1TkbFrvqzQKYZcCaZWwGUz6ZR
5lwOdpqTaETrV6WI3z2FTaCqpAerpk8pnOPI1JmNu6HE6uUvkPTM+ghqgfoq
NHmFJgy1bbGugKzsBNvF9psOmehT98VmQOXQD+VxmbMCKh+2vHb34lQP4zIX
xWgVBWCrz1DACbHY0pSwPYdJJGHyV8n2laEd+30m0HP5NKarlF8pFt1E6dEA
EtcIEYtUH7msI4zse0/iMdH7/98HMxKgNL1B4Hmzbt8uBsENyZYMkfk8KVON
JM8oF1kEHiyef4OMqRRwoRqR1VqpakKPnlzIE5Bcol9tD4LQyvIk8YPR3QE4
pUw/bw5XtCBOni3aOMBvk6MlUBBxt9LCA0JLTYs9mDivhj4HwFZHxaqWDGsx
nR/Bdk+31W4d5dNQrLr4Npu8KwDcoAeZwIWDN2nfpMy/h/pSTf9pvd5zyXa7
FCLzABQZ9xAcv6xar/EY79WjSnPuXI/rwmneAxJOOt+eKUEIYng7Uteam5UX
VOy3YQBqpJhgMOjprVSHoLXZuDfzKI75rxFJQg5q7p6+rJYGsgffLL464UaS
UfbE1q4oYWTd0GH5oovmShUbrocORX4ACk2rYFKuEf2EW11LnuQLK4tCsCGf
MTyCFiACBZ9QalFANWlPHbGEvfZIv8Uujnh0VoCiKIn10BC+bE9ygfmx2x08
ACje4ULqwsJzDOdK/p91gF/8aNJ7yU35vVwNX/jXlgM8mM4fMqmSwTt9Pcvy
ATdekdIOaUkknsECiG92SdsBZgKdzBnrPBhPU5N7gYliDQwaUzSBym6dpWc2
yNTEM+tzA9A8EgeW3KX7amc09G80ukrTNXy5LkHhmX6UBN/dsWp3Z5X5ebR6
R5/cT4+KbynLMMmo2I+vvMcswfaIaEzh8SPOTExLZZSzcJ+B8i0Y6D6hEBk9
kub9MxE8vXx/crJ0+xpOOKnR310h8i+epc0fjRG6yPHlraLzjcNR9IadCjaZ
1uGguV8oWji+KcDQXSMYnJthh00vJOUTylxFlwDyAIPN/jVJa4n2IJPOToxs
LB+iiBQhyEwRCN9GWpOF6soqDsdQ/9o4nYq5bD7LMAhVEX56PJQ1XANIJj3E
W+2+VDw8GUy6n0OZWRuFug6Fpii5UsmkmW5Zh/goPA1qxS6d5RRIrmU7Qat+
m061r/Gl0PIq1bR9xOsmppF/smj3DVbr3QVi8nIxhKdCtqeqolMUaeekVzru
nmdL9e5NubdWD1Rg3CO3tZJC+66bm/uuv5M0FyM7XduSkVNEG4p3T7BYiInR
vKCFihaFaviTjaLsrGR2d63CkqCiJy4AZKFaZwhbkAXZBfAPZno2NyEMjU7n
yZUYjktKkMz3qjEF4rFZ7W9pimYVfc9WPw9xgz4KbwjE0WCrlKNg2Q7CqKtf
yfXwqo3gWRq8+wmZTzPP+AfxkhNDMgzSRax2XNbOBrh1tVLVpM/WV3iE1ni9
CkCSb8H8Vcjo6PIa8r2+kigD7qSAp0gf/B8sr8RUeR/XN7mHYMg+Ftdhc7tg
mWRfdO08Cqn+GKBZuKqRwr4BgSxIQimvCUwsTdBPu7ExByoLZgCjTqxV5hKU
JeYLY8n03uTNpdLbXbsV98C/8W+a0dZBsn5DFwK4wDopG0aFYkGNiTg/V1xJ
bKZqvR8uGApuHjtT6oC0JfsnwMz/85kL8ex9qg1opZaSAv+tMowrNZKIHKvk
rBQ0dsmaRZs7Dy5KgfcoCqHb82qtQ1j5OKYQ3Ql3DBTF1fZHpP7pbtofEBX0
/pJzCd4spD+FU8FQWZVIBbLKXuFbtp8oQyuNMUrKjYkk1hKTsD0v9lBeqF7/
iEwlF23mjSUNbNfEfEG+szjufFK2cKNyK1FU4x0Uj+YnIYID1U0kKgDR56uQ
fIJVgEsYh/15T5DKhkDofcj4XRduWGP0vGV0ncAWuoMcbuZdSZ8+PNZvKNSf
7Ly+z/QYJmkJDZvb2vn49LMMKx1e6SVuvcUOQbIRJwqf70iWrrmgjIyuz4Ih
9rMfpgRg5Fs6sMkgZVI85qU/83GeKex/TphY5gtEDlGeqUwEgLKynvYBclTo
FnwSj34FwdqAbtuFdTvsUy1+FFUUBUtH0iudZmesSCvTF9M9ZLg8H1dx4fzH
cMO0MNHHJvadWqK8XaIDts3z/eZ5HDF2+ECJybh+T6heNZURK3cKrq2VaJLr
G0BjrpqsHW2sILf6P05s6BkTjud3U9Uzm3J/ckG/aMrSvGv+k/gl2Vucqa8E
Qa915j4t5qhsj4YCZp15pDi7tFvris24EUOxi7cUgmtV9bh6vWIakQyXCsS9
UHbWlSiZzSX3yHm35pfU2Pkik93xfwSBd0DkgakFPbEOUwWQaAt3ufTaESAT
tsNw9uxNQRYVirn9uDgipGOaHwpdEnGekjvZBX2PIZF6LzbiVHPbn8Ga5IeZ
/T7PsCrmMIhNwQ+59CLItVk2jb21UBSdCA1Ed7XTqjuk3p/zqtd2xPzAXmu4
ur2OJniazMNtqz6NHqVusjOC0B3QI5J+gfldJQGFk0+O0wbSTA2WZHqiVYBv
azUdwYar2UOUjrgNe079gC9oR82lOY3nuuR6qF/05NdK1ppHTVE1yfSQTYb5
BJe/5l9J8KVzCEioRl5z398LtqEf20jc/K0s/tkI7Z9+/3BVUMl+1+NoHMIV
3/SlpI5YhKDygyeFY3+kPcQLIsLyrhYGL84T6z5itCmNeX1FobUrG99Hk4yG
7LDjneJEg7snzvLwaup9bL/G37BSNX1YhIAfn9DSi1t4pu5THOEixmZcRX0N
qKg5d5U+7WqH5ikDghx71n/AEo9fW6cfQqi98Ax91aec2Jm1q9N37u+Gw+Xj
35yt09AoKWKbjx7wA6N5mvoIyz9Ges1M05Nyihi2suapC6E+rtzjl3sjySJM
bm1MpH4U1GA0mMHv3130U9HphugUsb452HYl6Q+Zkq3an+o8weudKom+LNtI
UfA3etbbfCu+FQc2wF8OCH+2+VfHVaN/h/kRYTXdYTVbVlkeYdNTNby9lrPh
FCr06TL/nP6vk+qAB2veXhtU8qcL8fxAlEmbzapGRbDIkafGjQvj763/2VFf
YHVeVmVM1AQ93xLDUxKTW9in2wSz+/bS45F4WEpCwLRphNVroXfe1nMhA/yX
yWsU/oIH/Y87ZTEDAXlcHCQHf5jNS5XmBKzixMPX24X5ygSYyQ6g1DOZVbsC
JHeUtfbQ7C5yXheEWgTvpEqkZRwcj8bgg5iIHwQ0nhN9gMPTsjxlmnNpg6j9
Dj2VPN0hyacUfPHm7zuLrnrlAt/X04DGyrWN4Bq1L1/qL0UD+ubcMErIBGyt
92F///43jhExvLcXRE65ArG0XcvYiX8zXVdLBGUpALnMKjuKVPxhU8o+Zy5t
NoYyLvXzNP2wKJgw3HwaJH0FsIg+Wpr1AZTPiGf03RY8Mugtk94bQihkpATq
YMBcb4KU2ZpcpC5MdC5k61MEShKwVORiSJtEmYSqJPsIE3+2cHnhSpDa6djy
o6NddC+EFiYQDpkLt66tUVuXNNKZoNreYbmQOYTjgG+aJ0kXTeCkEm4DxMn9
8sq62wt+8HDvMqMP9AnlLtcgMh/ZXi2Cl0gZ+/1J0qBJdtrOgK6+t5UdE2h+
s/WfTP+oQTTyA7E9Yp22ergArGUwx6hLanCIY10/gtRJqcirqEqZv+qW8fxX
FSkYIEKnbaNHAFqHd5Ve7eQw5oN7tieA0syeDyZubS6zQf20mW07NXbFXoW0
h+SnhMIP1jF0rroIuu2f1Hyay5kO9NZLjPtF6tBRNaFFUvH0VtDHH3YvA6jg
/WcoXAWX1N3GNyuTNH3CT+7xouOXk2qsJdcRst0nQ59DgiupXGIEziHW/EKS
tPsBe5ya4Q4tMq0M0wDrSej9Nw8rhb59zbdstrqmuc51Z1A7GLCl03CMg3AG
ehRGUMZY1Q3FG9ZuABVWlD8u3A6OS7t7St5M72pvb2BpIQdFcrSPoTGbVRSp
U3bJc6h4QlYkch9l7O7uWisFEp9OXi6mCGioBAUmvGITkiuObCegedwqQQk2
mESTbiTAeVqBs9t9Rf689wv86fNBNtEhnQfs95K3m8qifLIoY7hAoWeaH1UC
Q4CQoeYAw20Q3HohKs47OW0MMQMTmFFIP9C+VKdi+1sV+E+0kg0+QQjhFHaD
5kZ3c/+vmWgRab8p2ZttijIqdEJJpqfJk+NLPUzmExH6nP9YXIXGTZDU0Bp3
N3JUyWnUae/+IeUff/52YPvH5wTaRE3UEZaez+KUZ2cR4k9NsWEJnBzbhu59
nXFkL/MhO/52Nqv9AlzyerM/mbnM96wisMn6e1TJteqXx/5JWsNljMgiGr3W
oP6opaG9767UIRVMmArXtAmK4aFtxx2rBeHjMertvNV7rp/dhqmUt3MjXzV9
Q0CVzMY3NqEhaKqF2amXf+8/1uSsumpmS677GISX2WDYUyK715IADNeFC4ci
9HKyc3ijU5Q1vuX4spXywboNTNdRGkxH0xcwpETJ5EjqEOWEltOjLfuQaI7s
wkTvWf050+TVKu29noPVfWKbaFPqDd9GrecbIJKe8yS9OHJW5A0okaXqRHPo
jdLW18JXF3+wpyOrgp6H+zE4VUO0xB3e2c14c5euRrHua8JcBKR2NhmTxi31
nWVeLtZbAMJhkLlKLyUH4H8gvVbnJ6C46QPdNlkefr2iPURmudUaMwPS7U7u
swQf3wn+xktWVW9zo7y1Lk1tPxJHtwIHCtc4k0LccRTwGe67qD49QxTdFBlp
FN68uBKghEjiFSqT7aH1J46zVYpkaBdMBlqLEHFsmf3NzWVS7Mfb/hnP9aLu
AtE1WSztdVJtSVbcpSonMRn/IRS5qpjNvPUyD+T4INdOvH6p48KspiYItiEm
MrKatpsBI+w97C8FDIPefb9oW+eCYp9fxwRfxTVKDAVuwpj8UQmQoznScoMY
OvGnpL21f4jaHuVrVTeb6iUtJ0hdt3ta6238Paa/NQOgwSel5ksN3QwhOy1b
hZdQUqZl8DD+igBKS++m9cKt6xNXEliw5Or+YRAGujcVKEGOb7p+t80I/VQX
g1GkQBL//laXDhClcSlWL4wQOPpIRQA2uuJeizLHDi/bhQtsnDbXvzvOOm27
zULrFjCO/TKyc5hwlFBSxlzX3o4X1OY2BVGmQF9B0Fwit54XY8QiiWmZetNp
OwMcxnvLFbeAGciXIQ4ac20nbfArHMPuzxraGngd6y83lkaYY3D6tUwBuWMc
aFsCR9qbYO2rcKAa1v4MbEc2wgUpQ9aPcwILakMg4JRh4CC9Hy6bWAYqjtZt
Nfj6aGJbXBOeAZQdIwc2lQeDZmyEZ93CA8EkUOE4Ca0fFN3lbooSHZTKhnyq
jaXbX3sFZKNHXMWWYusqYG6xCoYsK1HU3E7cvvxWMi8qSnXlx6+4FOSHvyB9
3gtS8LgK6rYdqdf2vVPTFZ2nS+xTnBCVGQpa+O/joiINPnVzrLszTyVIXcjL
AAANMYchS0bJoqc+Q+a5rUfxdTVbADDJmA2n0VI+X27Wzq9NyeweN4sjtQ/D
uoqguZ5qU6oQ2SX4S5+cXVWF2VAJmPm6zK4sroTgqYEl+Y5QcEcjAzvCG0CR
/eai6BcnwUexzZ/JH5twwZgTrRA1KVwG1z3L5CSJPWt/CawruR5Mg2QYVeEC
sxpmtm44UY53RqtT1RknCaDn+GmBYJAxoNOHjXyCx6FNpgP6CtSMmKUZVqLQ
cUAuVjmow63vvljPbQI/pSXn8QP4IgOv/YMIkEMc8+tN9IZpk/cD4TzpoN09
q6442EvMsFG3UwPpspsb4NBd55s3OIAlvuiSRKLH4JqRtdfe6WGcE1nVl4x6
NlVDJlx14a3Dh6W36Mt7PhzmxFC+XRrcwuAAzHOZMwLKl4ogcB3qZHlEekMe
gGxmfFaVeUh2xVGKvdO1jDloFTXoPYSxidXxQMiKDHAsQX6nFortIMx7wwt0
84QjZXO3+AyD2moGWFULWbXfiE8r5xloIEbeAStYc/rvgSx26cmUolKnOIJ/
TSpbDadUsL14hOHkjr8DHo8fNCd6WAdc9ebNq3k6z64FJGrh4eRcFcw5NiEj
J/meh6r+rEBA6zuRsINhM/TrNU2r2UTmoNqCOxL0aFOUdoBuvU1cg3LwStq2
h0dw7RlGqnLeudftjotCEDS7JxkZ03ihFOy0Yk6VjyHAaKn4Enesa8lpOQaI
FJyHPpvVxipJmGEatJss/Y7GRql8b0V+iBdU6nipiGSbfRHEkxSNj0HD+IUG
IAZRL3t2PTXVbHZowTMfzUuSTx0KsrcfgITPTZ3+Cv1vEUpmKXZN8vg7RGe0
xHZog7CVmODdGPpGGKYVMn4DABQOzVU+DCyz0GSDI0PsP0P8gIDqVNqJv4wz
UdkJEGaPEHtpx9p0n0o/Er9126t34OwFArdFQ6kRtOJ/wygNwF6mbdCyTBtS
nHklJLkwFk78gum6t2GJ4iSCmaBNjjgJn5DUkCsyk7xBeCXHYvI8pRBZlMG2
qmuH4VNRieW1PhgD3E2fz37fW3Anc6PtGM7b/bF0dgf0wBF/nMtJT8fptnIa
DWVlP9j3vfHNI6O+RuG+ybaJKBvTnESFtyrg3fdUAFePQot/DlDYPXXxQhaJ
6W7WCHKE87JAjvKnu4/J0e2FP4zWRNyxPqELOnJqLF2Lgk74qA+2gXRwo7sU
XxgSZkd5LMfHNuJpZOkpnP2fAyZv0oVHFD5dIi0nqCB0p0oDl9vL5liCVcKT
DK4NGIgNLgR3IEkK0YDYsK6ksS4a1BBJG8Oe1qwJm6StIZwHFgjB+cRH/e6G
b79Qwn6o84MfLOFwePdewpxdtJsjqY7TgUrLmTx9AGT2JEQbXjmlCefck8/p
3+k5dTdqz3LylRrPg6GhCzdOqKTO8CrHQAw0bp74ZuoJq6TnbJSW4TYkRaDR
NyZRHqUemICDrKbHE3Mvo6jVrIWdJkL3Ar22xGH8b4pS/Md4elWCtK+NTFe4
hvD2xX6yZ8bXEqJBmn0ZsMsuqH104FNCrjf6eWJ73fCDYjbDECBa4HymUpBz
HQQ4bHoDRV+KINddEnMa+qnzmfy3chuvqTJcZGgWzwui22Wx4192btFG5jQ7
O/RXS20MLWEf/Roi/ov22JcsK2RBRv56gDnrbeYBloJ7ROgHXsNsDm7ct5Hx
qBZMczZ2iVaUUg/+cTNDuTQegDNXL3Mkhqba+fQrzLU5eozrgbjnsWzFLRAu
vn9vn5HeZ43SzUNifrMoF3x2Dywd8YDHTUOy47nGFS14gexwPBC1ACU36wNa
slsRmcfWFqauvnAzdK1ny0J48Gn3tUJesTGBLAQ2fFxVXxKmjplMzFqNlzXF
1qZD6TWt2yWXkA0Y1scSnm7ROO8X8N+tsL8BsWFbWnYf5domkHfc8yDIDjKn
zTwGcoMRHkj4ts+yG6tdebQPda0ACRYmoMZOte2LO7Ya4fSp1gW1WmDLmHzF
BGg8wLKSv7cN4T54/Y99iF0FRPZQxraEonn3DJQmsCQ1yJT14qIK81qlMK0x
b5nUO4J3S7muVyxLM7dbwLV8R5wI1FdEVH6TR2nU+0VeR2TxMX4XxpCGQnp+
8KVmxwOh7oVzsXpSESgcySS4fltNXSFmfJacDSG3c/wf8XG46Y6tAOacCGBu
ASFpJ6UuHaXQC59Cjt5qnIkJxWuGp1MKl9vEnH+uFpW5puIEzF2ltU2mvcE/
6IrFxz6/sLoRen176lGugZ2TK71LyZlBAZSjhUPmZU9fGHy09q/ubcOaGv9H
9DmFPJ4wDXcnzA9vrIvAJO9QwDixHA5OqwkJA0PKCbELR2GeFFnh02tulo/G
6Jz9dS3hLhhXmTri7t09xD+fQGaUeo7vp61Z+4pwsK1w/gIVbKVkq6cdvkxp
hsfDqMNXrG4ZC14CeKADk4AQzWqpB5sfXAFP1eRgMQ1mU/uZAugYgLLfdI4A
/wXw3Cu+yI5s2mHedkW15EBzPi9TDE6j3UD/FWT1TP//Qjzfuo/n2L0T07kR
78eVHtLY73Wg1WhmUPfbowb/4xux/1nwHBHsLMPoWBHygWNl4JE5B6oP0Fgr
SXRrTLpTfY+4zVDVa9zx86xu75fPSeXLI5lvSuWmSZ7oqxBz5GKlLxKoTr3s
yreJcIPd+uuwAT/GZpgr9K+CJWbn76TPjn9N2qMRzV/OTkY4KDym63dsjr5t
8VnjQ6YRkfqzRNjZKhgPH6fQK0hThRJ9XAQSNQvANmLGLPOzUFDzSd/q1ai3
siwsViVPD71lUOuSNix0MtkozDyJVIuwK9DBQQ1Q0hZTtPmNH9RYlf5WwqF2
9Apw6wel47vf5bzYNuRWqQOsEaGeb/9hIXCVEsW+Y7rdcur01Z00IulGqgdz
2wZx1zdYGjAPCyrplm62cdelnkEgfrA/KPLalfZ1alwyQOZkKIpirileWBLP
sy15O+fdV1A9hX3lPxLdkUELwqPXdYRoE54IVgnDTxWezRjdyOORfz1kOHKk
SRymgYVKzJqgxlxS6M84EMJEB36ooz3xXCuGEhKIyD7ZycmnFAPoORRKf5my
b3rk+9Fd//+xqauEOrDLBUg4j6tKcSZtJqVnU4uIu5h6nCYn/e94bwm8GPMK
8H9brkbepHJOF9tl9NqiuriiFo/nosZiVXhh44yhO7PexKEnzkCissU4JW3Q
uYxbblr2iEVRy8GQN2eYnkzrI5+JuDgTBxAvV2mo7P9kxBhMAhxeG8RbJf8J
nBZATH0dYPCPb4D+ERMTyxKe/o+dm3dnDwwAbWU49kRaEMvFMX4M9tN+d+3S
ZzFynJcyhhJ2WIsBPvIb7L2LWTUe7bul4MnkPKCRyRGulsiCqFa8NKYuKkde
P3HT4bF6VVXbS3qBJV60DHJSVzhQ37pYpaqBklsqimrQBcG8uQAkRAzmXmgI
dIEyVHXlbGmdUrMXI7U/0LbWmTfBAOCxE4R85IUTH+tTdwRk4ScTGO5TeVMm
S0m18ycoxwix4ARB+rhUBeyolI6VAa14xMT9jKty486cSFsPTb6MM2btLTXb
2mGFMzgVR7Etp5Nz/R/68KSs1gWomq32U93sHB7FGrsk2Y+j3C1x2UtWlela
E2kj1Ya9fIMvI/ZFyg4UrN+KhTgXSj+L5OdHcYtsFoEGHiDa7SsZ8gUgYqzf
C8zz4if+k3dDqVZRNBjil4t9mA++mW+O4ZK6bqpO1TM4NwNbJQ3H+EB969vU
l6VG85DZNj3riKO5oflo/f+5F6c4KnAt3xexy0gmDRjWloqt6t7YKCyHXJlI
WVEbqnQujW4+oQuP84CViyymW/Xu4W/jC0hv4Ze9Q9ZUKR1QvGYwZGwlteUV
pV3fBHofFo/2lu2BGlgP7D0NfrGV+k9XAjfvdWV/uULxYMbcun2YOcOASyXQ
rYT7Y7tvr72QEc5N8S4ZbMhn4A6B/BZV+9wxwsvxcNEsBjgSX9Vm2hTZGBRH
13EcJdBF5w3192CAToN/AHZWJNGfT0P1HYoPiEPVxcR4iK0acs3Uvvpx0wo6
w0YciH8X2f5EtQQVHRQI2tv1lkxTBRfS6tzFj27GweJ7MPr5QZ6mmx8ZCXSK
dp39digsNx3MZyarpIn1rgpbU2/VvmXpXZb6imf2l5fAAhM476S6q72cSYV5
elE0Q40m+CYumwxs2yR9pBVUpq/Oug+IOsoGx78DHWDSxwzmA+ciOPoCuEib
oyLwPzqCfT5aVTYcggdCESLMb/A1VX2sFwDxFy6VfJKEcaVRMxI02vU93fNg
KY2i4eblhkXrnlfnlmZ847hev5NiTpC0ZiQz/hI4dMTB/4DLltAEV05+HPMw
K9jriDO1n+pWqaEEtwow7sm1TFD5vNodzvf1wWjscedT+w9uljpGSDiGw2pw
zMgw99xfGW6wSpfXLvUfIFnkDImB9DFXmhoqkAsu3G/zzYpU4Vn8KC8cb0JM
IaE9viYwcNVGw4QN2i1zGY3Q4K4MZF+gqBJuXA/hf687rnfjAehQxMS2CajQ
5Ua9rwkkbG/5Oxp+hV0rYEe/qAiZJiv0zC6KZYcQS2G+inPHRo1s6/jPoUV6
ZMIE3uVryVy89bNURn31w1q3nICkqccA7B2DGnee8O201LQn1+Y4hChsOQPt
in8cOw/QPVHItveYQdEdjzs6oKl9i+3UBlizR/YJqU+B9e3WeGNAF+EnNjxl
7jd5V6+RSg93+7lASVClqGzU/7eg445/wei6JU78stxUPgoSXHnc0V4RQQo6
jTMwf5Y2x9uFBSVGnvmIN+5L/wVcxUWD+I1Xm6QFSAYmZ018Bq5Rkpe0xI6+
5ppXeSYcORk8xk2EMxdnKK7ADKlTRfBY9RUJIMEjIep+OZjzqo4lGTRWCeyL
cispTN9zeYMrCdaNxVuf2lO5Gzgbzh9w1kNvjk1nMuH+uCCxY1N3+uk3nBYs
YPDa2nHhgc0G6XoERMk6COF5mK9TFzfzr+L8A/TEAVmIcqM8bOkWB0HSUdKl
MQOFdainu1ntiz5nS479mwH4854KoKRWDycp5/gkoljl9/zLn+YFgKt1LMaR
smKoVTnRZ98sthh3kef0UfKqrBfdKKKVBHVjtaaSGOwTHVqsvMQtEBuiekXU
kPhCZ7qlzln4aktyaHx4GRJnvysiuJxirbHEQ1Wb8g2qTTzqG+tQ48Cjs6ar
QAiT1t17yQg04/tJ9Qru+9VnqsAVNIXEwVx6PrOs5/H58mTvR/Ko+ZjvdqIY
h8qO6QBWEooSYAkfwcVLJpv0awpjxUufjMmKckXgKK+5TyuTYRGpNwRhdlgi
WQtW76N4gAxMDqGYKV+8nxFFx66J1/st5ojlGBLKRIVBMyVPnyRJOsRGCEHp
XIl07shT/bh62q6j+8r0JLkCTaEK4fTXRiM9zT6klYpcSE7bFM45l/ZA3QRc
rgzoxSkeaa4y3K102DF33NYTubVkayQ3nyVcbPGm6iwVdl82RM/H6W4/c6RE
+QE+ku/g20J+sCV27cR4rOL2kyXZ/ffZCvvxbjrlLEnJQWqVN0RtThQv5kgy
7NSEIt5dUPHjU8pURLJw2L57WmujCITSe71UeIRD493lEAV4TG3HWr+eZw0Q
mR2T7pcYoU4kS9IHsMX/T5s8zRAv0Wugd/RSAeWASEL9CJgdZOKnJhw/ZYQQ
lZfWZUf23VHS/zvTtvNkGyFCoM5X62Md6apx/x5rFLAykLc/04qOEgGtGGot
yOnS/iMZaUXoptnGciK5TZJDc8NXgvxtnqNO2paPRmWdE3eskF9tllSMA6i7
DLNN6X9CVSbCkaX2Y7+h+77PKFgQOU5I13WRbCu+bt+kC+51DtHbk0k+YJPn
xtBknmf3rOVDxLYzaU45K5Ry+z3pZjI6RAj4MSaMnp6FsQnya8ons2MBVCU3
brYciEtfjr8ZzzMdl38bWJY/eBH8R5XpTQh9h+9cCcbd3j+AIrypTR9vNrpk
fx986zcEKISdc3kXLnfGiOsoCq98yih9WlARLnksFbUcOP2K4Qe+eUQxaQ8n
+7DfoYgd35Lksf1gZo/tiXzfTXP+hqdQKz7rzQFhlOFkhaDBhcj7Cp3yOgTi
MEcabmFeq21GQtPci4jBq3W7MU812r5tTFGTFJFDveIsTZtf/IYDA/R276qv
+NF10z0CXRtUiHT9UJm5r+2WoQuIs3b5Q4UO19JmTQVKWnLrH0GcRGRENQlM
1jPeMbOM2eYg2KEaDQtlwA9ZYh7x3I6RzgiS3wL9ILnB5cgjKKTAmCmW3VUE
ILfhBwGR5UMfvcMofJKvzGYVOW7yVvX1Iw5m3PTQHDJg17OGkFRAHL7J/CtD
L8C5DOGTJxM1cmRQiSSmqsVfSYg2Px0GBhgRrIQB0pjrP8ZmuQSk1Ln8QSi4
6vfXtbTausMoEhZplH03skSNDQuhVcFNYgefTLlRzjP1IINoP8FS/IaprNKi
vXmu6PPcCr8csk6ZzwA4zcc3yQwP7DCsyFy2yxu0UpB0vyN4KTuJH0YsEbBT
HpN3FjHi2t3UMN7CUzzCm+Y+aEg/UtkSRx9xoabavT6IY1DZwZ60WSrthmWf
f5P5IHQxvipsy54LsBgyA2KX3M8fVUnx/Z1aZf3tOwXvJZu+yyiViDsFclEL
tAOdapVB3D+FNJvOr/pbaxsQFBJn+zL6FsMQimfp2j7Ibw32WfGxt3murs/u
XCpWZFhflcb+4ivV/Kd4ijVDh0I+n6LuSczY0uVDB8cVIiaa8TRZzbnsB+jt
1okRVAp4LTegMKchpUNT01GwyEiWuPABZF+mzpC/kSxsr2d1u0QAuu0YI8YB
kfIOvFrAbek0ZlYWs9ufUAY0YRw9HvZOiyIS88s/weYDWj4E7L6LRa7oTFZV
+Wdzu4DheYad65lTXbPbNwfhW8dFKPqd/xHZezPZ3EdoZZtuc83ZOlgZ3ukq
MkDVdzItteO7gwIgKT9mZ2zVO8wiSO8C522wo8p5b1HKsIDdYYcHo/hwlF/E
xOPuw3uC+Tz6ibb7Kuow/hnNUZtEaSCUGxLywA7e82Xjl/DFNLkh5OHVtO9/
ppawDH92PaHCdEsnB+0m4MoEBXezV45FmQkopE1kgk2XtgL4wxpg3BHSpkNl
6LMRmiSSHPG/FAYCd3OfncecofTYxZ6pk105WWnidWe2OTwcqmYjjUzbBze7
uoTZFDIeR1TQZK9PFOqW80PqLRMuFRYQ0qML2cYEr2OoGIwTVvXYDzDnmCUH
jH/uAa3C9xgWngeAgmDeFUG8EIvcKuQH/yO0cC1ZC6IZFnH4OnY+bjEK+VCD
q1y7bokgd9V14K0x3IbldhHQY6/+E8UX6b3359Ervz1gjXDpHutYrjdxJPQ3
JxENz1BFW3FakMvYg3H5v1t6gqqK3LyhGe62GNa+0D88zkg6YczAKhZlUgGL
0Ea8PnsHIJ4Zb9y5B7fMg+1aFhZIVrBJT3nCnfTdG8MIkCzwHXWYk5oeXug5
lObvzP1f0k5OZo/mngOWoeyNNe2VDDfFtUPlJ5mP7qMhE3AZsJotVkOBWzdn
0Yk3VOR9lZK8tblFuW04igGx2rEuxcebtgtViq2oY4OB5ZL9NkGlu795aWS6
KfXKpIgu2E27m8tqPmH4+jJ+jDnEk9C2PQhmMRhCiru9l9qrIjUSg/4JP6sJ
Ekhvw7XHnRP6QCwCPVapF3AAOmbxNNxePZQLp/kHQJHgGSm1+kA06wql06kD
6WTLF3EpG166daNOPvEcPbTkUUIvil07NLxYlklAAYr6qvGwWD5GUobwhB9T
i56+Gv1efX4CbGAqpn8kVi83ZpgXetD7okRvrJtG4sQxYqjxt0sWaG7nXtw5
Y/wwhxYfVdskbsWBRNI/beiAtMTcIfsByFn48+5f7B7r9WtC2dGt+MwA5nm4
QYnOmpNg4u9hSqSG++zvfQ4+OzTOJGZxDnScW90D737d19R3wDPwCT94bdjP
BXO7QfFHIXmw0hIg5w0d9LYRT7NneI96PgNxQmo5xEFmruVhZFeJgRKF3P/p
BWVgnMeZZL/LInhJ18TkZxAwXqjoadtGijyMHGB4iHczxsFo7r3Byy9rfLwW
rnusGosPNsIjRYfqwRcdrD5EC1ElGVAjyv3E5Als8Cj+1jW030n+MnvqPSgR
+V7rV5DsFFiJpEzDChuIYKDsj/FeuK0CZ06E40T+9GGUAu3CKV3o0mI4AHOD
s2JPSHWloBNKA49g+Ch9yOFLnt2hEpDegSQ/n/mW1wXsgArrEzGZNmX9Sa2y
jO+RMOXe+aQ9Yys4T3RG9NnHKeF49B5SBOkl9r5TXph1IVAjuPC+4oE2Dpha
QHXAKoBLdDzCl2QIX+CbLaV8mN2xjuzxQBHciUH4eFrud8kNcksKZaXdDJJs
18ns9zWTBgja+ARZJvKkRuyucCmsL8GCZZyvCOD4eJJryjYFaqoUVjJOw/a+
YTsePAfcYz4swO7efDbygKdc52N60CG026ynXXLxTDr7kMSCR/b3MvbAFd4Q
/G4DmPJUFLlZyOynobYX1ae83c6w6HFdmr46YLt5C7AkuZKi7dZJhjvsX9Te
x++lbWPPY00gw43+cFsxg8QZMz5rsQjZQVioKKNtaKY9qMuXwOvXnaFBn/NZ
OwCM7cmPKZgJmRaRbWnIMzglemZre5CDYHBRY0+tQ+wb16EKPb1b6H2WG/o5
8jF5Hl7EG5ne4md+/093l6bq5LWuJ25pTo97WhSBrszAL04kvykHAz3qx+9u
ZEhgIc3ciUnOoZVMk/tTAE3PzPFCOjHXCPsSlFFwH0qf1v0bA+uDsJcEQEOx
LOHBqlzQFP5c0hMKNW+TfL78ImWSnlBTRQ1AZYI3ThBrSdx0s4Q7l46gNTf9
OZTbA0Illrh1+FxmQB87ZnT/Wp35q6ydj+D6bcVBuCzKnr2fvJsKcWgl94Yx
Y4V2ArM5SZ9PRaJB2ydDcAN7Pa7G5Z2LuNzhSpN+Kn3VTUjefcV1tarx+GW0
8RFRPShfDzVWpAcz7NSXXdtNurCUIbJgP61Zr12mtvN6PVPRNxXNEQYeF19c
AQ+iJKd2TJDTiizBAiahcM96gpT9FcWyxAYKgFgH01HiF/VJVl1EJIXbbeFw
xo6cCjPfCurvlot578qbUw020XEYPZhxAZXt0+OMnybYEjhJCVf3lJBQgqeB
UgLTDU1/N+XbsyjEqLb+WtagxCLt8Ga8/uMoQcLNMREt1XMRmxhlLV9D1tui
AjKvQ529zbayfGtyHIGx5+tYt/nfZ0hAzIJ1Yfl1Pdle4ba7he6UtHW+j6h2
83MwfQF2Dns64rEbGhHdDknm640E6rz+SMGtI6SDiQa6tlAbcd28ErC5crBL
03rNZRCwXifIa1EdpsggmlYxnckJa2CQNxU/vJJYcajPG+9kWFiGoZANSvfi
WXn7t/5+eF7zuLL1uBSufRZi3thwrIV1It/stjgFqNnt8mEj26mIDwvNY4/F
VM8kHpalaDOD58HHhbk1NDbQhNJoY95mbvZlArU42WUgEe2vObNVb+Sj2ksE
oBF5j070QOvtOOKY/1GGyU5zBNI5hf9GPnVCBc0FJYqqX4q9QZjLYe0G2gX8
etHDOl05VhE5PuX/ZJ3uyriijeu4sG/EjolAlmLsIJYC7cOtkdxwSdk6UDha
XtlEs/5n+XVqfw7d+/mjF7SFGoblBcAolR4gQAC20sLC5ZE3qBjCCMZnEvja
c+j3tgMuTB+Jc/7f0EKBV5OGNTkzXDFxOLK4ehNXH+qqGJ3axLK37XAgbQcD
WMIKpruJtOXNNGJRI44BjqSp9HL6T1yP9J2mT1p34+p4f7erAsKxb2e7m7Qt
JiaiBI8m0sn9FIL1fgVbFOLmwoeHPyrygwPlVaORmOQ15Jyu/IV5WOhuLjDK
TpAMQImD3p/ft9nOef5HqpI9kDSzNOVK6A0bI2xCVHhzwSz+cPYnBJ/TuyXk
IajdU9mZbSMC4dm4uAlpuGaxZUQ9aLjh1oFliEttS/0JKeN9hfcPj8T3SNjL
SgBM2FiYhint5Wbed7hD1A+79EZFlxovhaOp/mIulYgj4HakHwVOhvuxsmgm
/uQigKhgLErOwypgNxKvCTHCKub51XmlL5psjWw/qIVHa4A7nsxh1pTz67M+
lcLB1Iz88YW84AMNzvd+MZBtxzjpQana1hHtpFI5OnvOAqutyamhWtiw7P3G
8//XNYwxkyG6l9YUkRCKYN8IBf5IvHgxD1/R3fk2Kedj5WMv4VJ4a+7ZhI5t
0vVNjVm1mRjH8S9wiQuHzCsp+AgnS1A2znh+6Fmoz4LKNjBuF891XQEiX9ed
nvk/qj6HD03oPYMlmgkCol64qwZ/oVjwtn6FSAR7Z9f6i084KgOEfnOdKsnn
uGujhbVYDU5suXLt/PkbZNUXki90Hf81nGZ5Z51OyG9JbF0lUarIdwESu73D
BxKlVH/5hIm7FB18LdoeVQA2QGDqBYrRmRaAK8DJu1Wdi05oJcdbCt5Xo5RJ
AQQUcyChEEk74Qaty7fy99DRE26VEKgFc+ySmWv9OzCYntHQhtaOoSM4n2Xg
JwykYae2+Xhv8a+7JQU46I3qsET3jLoQ0EPLo42CuFRKzI4bnXKqyS+M89Js
G3r+1ydEvoBU1nux8ep6edF+CJcsgiWmLAH52PYfirOnR6xtF5cy1V8392L1
v9KzLmHL4BoCfy/e6+msMzTTF73enPq8wY3M+og0Owf07Citr4+ATQRLemIh
Cmi0BVvHHjHdImRgCvi6iW3VmAzFckhfuuD71Qok/QvCnv+tTsr04Dttx3yr
dJb3rru0v3vymJYK4aNnLfDSIA09zqkGVV3m15b0djEMJc/QN4RkdwWMGzOh
+5XiEnss9phJdYxUF2M+Q4UkSla+G9qHYjkVExPoDLrWeJUD1qD0a+BwG6d7
54tiqzxfKrgQnf2Q2ZdPVnEM2QHLsSncAxmPc087B86bODdvbEJ9/UlZOy57
AFSdtc0ZLhoOwWe57c5jkyVWf6SZs7H8vqqqvkCjJr1+ahO//GIjbKZ4ZadW
YJ9HaphIicoYV01fVliXKzxVeZof8FFzFRWyzUw/RNBEIGj5EPkBd90pA2ZI
oMa3+80aOzg34PxbMV0gRT3KSViu3OFg52n3XkEbprHM/svxF8BeWpUnpM2f
XkX/85fbtFyMN8spvpi6jiyBZ+tEA2u2Vi1RL7vaail9oCEczrxlM/ikxl5v
UIad43i8af892kI1ZVLEI+qMEObqP3rjX8a/sVKNYdq+wUfAAw1CPwIb0HjS
0lU0HTJK1NOkeYJPMGV6dGoAm1fOs1ykGFv7wemug14QSzsTxZa8k7mxfx3Q
k1oRiyH5De9LJaINcmS6yv8ebkYi+AuxiDtzCZI2/oIBUA10b52meaqKCYjt
vIyv9ihFed1DcNiri5C6ooOTyd5x8LvjU9lFD37OZZFzUJiKv47CmMeQ1v4O
7qLHWObHNTod7LerP8gRCHoz6ZR+favsmDT93WhvzwL/GRtd/RYsxE2rNztW
+81hZXBJDxuUlw1xJLwCl8bTNl7DjdtKDG9fjvTOpNfZUkl8B4C2hmu9Faay
wGPcq04YRDhUbN243UDO7Zo34MmZGFOdIm8sGDeC3NzPBAMI+og7Yfc7oqLr
wMRV67MmHMNynvY5+/TBAuReb8sh2cZqgqzuCgJyW9Or+ASVbUjl8hKVWgdH
Ak43apbmQWgMnUzwmDM1dAP+VFtDsvX3h0a0KsaM+2MFq/RAMvlfLQ7KoxWe
WxisVz68w9JK0nPU6U9Mwz89vXFUVeXMXvOYJ/ce5tza6FTGHEoSfSO7Bi7g
2EuCKRZiDKGihrB2v8JFjB84hSjvYys+/jUYkWA0ujAX55KDLL52SHvrJF+y
h1HSGPc7SDc02yMEBbvEgB5VqT+FphTrNN+xsF2LGU1C+E7ihWftJWZnWrmE
4JMXe3ZQpx4jvsmFxq6938eOahSMG7/ecTGNtjAjYfDTS5h0BDBhHy3rlzdU
HmZ9Hb6z2Non55wnUdLZpYll65qtQQleD4dNsUpbEwpK32038vG2SUsNnBJv
4GnP+XiKEjRh4SZdFtp8LSaM+jp2fP/M3Sd+34GXUVPVxLjTCjVfwbiNBrIp
7YOndRuqxuERriARnRjxu0JTnGvRx9sErdqQCcAye6ictlENJFwr5tJbYiGa
1JelvywD9ufEnwI52+IsSqUIGCLGsiIGh0GOJheJhaWziLqczsq3cmtm+ywD
viNMJTX0lCHcoQlnoLOt9KQ3136Ordq8neOLEIehUbzE3y3I1EaU0+lCnnga
1pyxLTqyK00XjZxxQJzqfAzeVvsLyslxTKFNCc8LhfdFb6nPYbNzcgaIxxId
LIS/PP6rxk/Ea0Rl4ZHY4bAF92+VJfORTaRgAgMz8iIzOeTCUK6pCQ0xbSZC
Mgrq6pgD6H3Amjb+bbCpm0Yw51qwrikY8rUF1zopyEu7gwC6zSC1NY69xKHS
oeCTIqbYP+SUP1IqYB4e0K71rVbnIVBXAW9t6kg0x5vS+mEgVqx1OBmo9Ni3
19Doo9hFWAjVKiwiEY/utJ1+6lSixZiBQtp32jetxHzI0XnDUQVCYDw2HkqP
uxc+5JPuT5kT+jnu5g/EfWbjIq9r64eyhqpMPRS3YA46p+uK8xMFepOSHiYD
eeW+QAC+Hf19R23aM4udaUfjIJLp7B4JDIOQoWCXk04DiZsFO06QhIanCVPV
Fu+TIBO50CH5rSuq6zOfZjPqW3zmVk7Vl+42s+5GZC76/3D98aIzO9yh48Eq
zNOHUMjjBD4UXWowILpyrIx/UyY2KR8LeFbwDr0Gtrd1wqD9YTCr/YLo3zDE
E6xDQpnuTtkoiw7VbRU7dEBTlfH2uzMfNY6U9ULsPQ+RvasXJYJIz26BVy9X
Rab2EWKQWiH3rdiLINb7oV+ECOnFWd7QPz+AxLkl14mczmjUxowYAz0Je+/T
IRBKWyG1AwqatDhP7gTjCZkKn/Xq5K9YsQNCzDlgakDamWMmvalTX18koY7L
OCf+EO8AbcCcH+4yii39RokSD26Q1CNAe/XIt0sZnRpmpJaORp9RRWkpzvtz
+b5aZOHvEnZXsCYZGLb0LGbDTSk/B6Xc4tV1jqnAIVYNX8BpmYTw+uL0tJU0
x4zvqDVziUIQHKtbKwoWb39XtZ838EOROofE+7hBQUOeczBDXI4q1IlruA+q
wr8tGFNtE+WpW8tk2gE0SOrhk7A7dYDUE3gHVriwyZmpAJRbAOeT5hyI3qz1
cTgKhrAryjjxm6P3rcHFCuPTd/sPFZLDTqsVdBMdGPFrct6qCZCX4VszP+Aj
heAHcYrULQdJL96XdU/ZhMFjJKyAg7JVd0sbGDo6Vg+SGMWsSC/JBHtDzU9O
liyiiiEgrfGIT18CpjRGshgDx02pwAldEr3CbbfZWgAUu6CvD+ItbMlBLvMs
EmGAmwTApGNdZTREA26qrEMZTkUODJDMKubNuWPVjfdhyjh2lNhHcNhUCIl3
8HtJJnKaAoZWRsL6a5iLlVoAsiEVjLK7aiGCXXDa4glcVFNmc+A2QqezKUPu
f+pfEwps4clEbIjtR/4M96D7V9ddJv2QDwp0iiJArmfrWrMKnimKwPD/eMHR
dQW9dA7aHNTw/1rSQ5HI+wHxO1YSe+E8N+m196k5K/flyuw2NbEs9qr9B7XF
JGbsuILNwOpo03K9pwSLB6FND/4TOonLnsf30/ULXQoVLyIEUqzcdSAiCtuX
HKbToS9CmRMdPzUddiPiO7fOgsv5aDsWjUZEgy9CxNcvzQ6X+C1LdCsAxHve
uGwrmu96kI5yGv3yIGja3xSeChnQDaKxdqmGYQcvgpQgzdcY1upuXIGwt7qP
mChkr/ZC3EJ+fGi5UIJ55w1wdeKuS9dDISPiNNoioreUFRk+ctgGFInXgiqV
DEEg/z45+vAf3KEIiPBe0JaRUYfZIMy+fcsLf/SehS7Ij6oI6YPWCQHCIkqp
/+B5kRvmp72jefMyRnhUk97gdoSQWrwut4MiWDwsg/ATqF7JskA4l9ildHa4
s2aNnt5b0AR7Mn26wJtMqchy62chrmWyqG2VFuaMRSSCWdAhnlbFeawGtULR
TQ3SbePlLtEXLm04LRZoiROlPSfMvsVseEHJfImY3+Xa/NTRE65oKMVH+wEH
4mlS6T5XuXHRc14p19MgsU3xpQW3BWqsadJ2ubq9fT2J1ktIEd21ELWUafFg
YZbgeeK2SHrBN6Q3kvy3/L+Hu3IwJs9Y3IzLMFdkeQAsDAtWEa1Lp7/Vki5t
+E7ZohE/C6Ld7W2TC82j1iI4GCCL+DwLbeCPlLztv73h829PP9mie4ct5FRZ
WbM7bJx5NVsE54as8Zt8HIJhssvpuK7ndwAsV0W95DKK2O8jIJQEUxvVFyPL
WHOM36bQZYi92FHBgGa/Hzz18qh8RY/TVHbO9ofVZTHPgonMeQQkb+73NReU
c4IwLWrN5958jYz5EAsYIV9kor9mu6Of2hNYUfvqXDt8o3WmSmhi2HyIwTSi
kh89QVpYAs7iBl61m2qnh9frPOnrQP6n799a8hCzFZ8leQQVzEMYivk8HLih
8IDN6YEALFkm+T3sRF1k+LYhZvoE/HNtJZaMwmUIC2ghLo72QMulP7301bpV
yKl6un0NnubG9KPehvagf7C0mG0eNt7oNRQTTbUD3GhmGHwXe1ekohWMIt1K
gpL3DJWXKy1n3yF5laaWokxdp++LuApywIKHd5AZM35E/MA50EwT034lUBf6
6zMsk8LHBDQSHqZXczHrWGp+IMBekJjRUBrgbdHsIqPCaDG8nsQ3YjkMvCsx
G7QCmnhptq1lxXFzxjLrndzqB1Yyjtms/JUo8Xb7ApZDQ5g+kfYBz6cdFGkx
WX50p4RrnWxpXwuYPxs2dJroYU4F7qvYtnfECTIe6zTp71zXLy+mRNvpY+Cn
gZ7E2vjoSXtWDCezI/zr779c/BmQs1ZA42fsrLday8FD4LG8EEklUk8OvQ4m
jZWmDjtrtQ4V+OwoYqMWQ1F6iAqgK9esLTxqjS4h4VAhL82bj4T9lFaL559X
frTvCtZX36IfFym8/QHt+CRlwDvJtScHD6WsHb6LD2VZkeo1nxG+TeIdxImn
txyluQJ3yzlJqUtBZHkb2z1c3Eeb/pzLdL/aF3PVKY4mv1FXPVcA37NQqqBO
+EZ959RqTRPnzQ4E8c2BO7Gt8pBeyDsPrFDXq2uI7nLUg1MWCObNzPjFrd/Y
4HjtX/xdmkMTz/sAbeVYia3gug1qL9pGK6UJCj5YsEmSewEGavKxroSeAlMS
NhDndPs5dE6jPnjXl0YBZgQYFMFkgA+yCgmZEm/oH04YibADYj59sFI7WAYE
Pzc4rj7EnluYggoKo750miwrRY+xhd6rXukldFc8OtdWHs9gVvWzSgXX9PCG
pPbl1pxeeElqz29pTixalLf98+UrHvA4dDBRU2fnovJO2bSyp+Np8ry4lFZ6
q8+nV9Ubp0xyXF2qErUpXE4mI9deMRp2qaohnv+1ZeSnpAjHlmNGkjiZ2zCx
FMxH4lagkRK88Ak4fqVhrdnfu3Ms35kuBYwHVLkuywwRNRoG1raQU0TsU2QJ
+isEPG1hCS2cvGUwmx2C8S1nyZeDpjtw+T6Cy90veI0rrbEU37TKimdqqgdA
dkHY1iFDBlhSRjPNp6a5HGFbT2hJm5DBb7zripKEL5Vx/womJEo3rTwgiBXw
BDcqqXO/GqpPyIZR5+wM9ucTg4c/S8nqxIQsML6F6bQriZHpf5VZUk8lkDiT
3gnydD3dYH5bvd7B5RuRAiF0dE56ASqqPMGQRwmfyW8dvDKKepFyxaIzqOFm
cCs4dEedPAnhAJnZiZHAmq3STvJVCZiMp2W10eAjSvtFjYnw+0GgIiuuSZc3
8sAHFKAc8NwLTIO5VLmKccR/bPp0ETSNSaDkyhFOIBdRMOBfmU88JfNL+CxI
NAbWAZLCMsgl5M6UcPNcNE14rgkuYMj7o+LUPjxRzu0NETh6LI9uuLGy136c
hhisLsa/UkO3BcU0b9smLZNJEwaIg+fPlB6ewN7I5I76sYgAqPQzTq+BwbHC
6IwebB/lnF4sfdPYPOv8Wu1EbCTZcRMZ7Y3GmcOW9uRMqa0+fap4429ttv51
y1fYJwdHt70qeUaoFnulJhRjnqPYHouxU66KHo5eSRk93yfVJ7DW06cpAdh1
oFCmc2XTDyIHestAQgWudZXtJwetStIpfTINd2enIcqO5F0nHsztH399eJS3
y1jUsQYwN3QflfQp0Sd2r4A/oYdtqtvAfqgkr27Cee5Q7ob8e+Ah7YLiQGvC
b55NRw4GCVW/pH0pOFu9nUBOyyi/Grtu3IV+q9+bh4KQ3tksgsVczF/UR3j9
jABX/7vJzroQVvVMd6KVq5dLja+2+vllLfwem5SozL4QbDOEVdV06vGcB1HM
gP0aPcCRbsUGa++txYYcn4tMuvrBkXTnp0uy2s32+cJGGxRq9aUVeZEUA89a
TzNPNMpfVZchiklpZsQgmxQ5apNBI6ILenqXGLJD/v/E52XsnnbM9CUKlaKh
8teopl3yzaGbK1vsf9XXkL0jq18G68ol1CH2lQ49c8/l7G+HG+Q5M20v5O5n
8RebZ9T2mj71x3keu82QC6Q6JSI6qkjVR3oioFcId4PIp5A5Mv9LeWXtLcgd
0kqHzFQ37MdAm07kHR4uKSzD/R70q6GD9tJ6U3iz8oVtvj8glTKGx3Vk+k0e
AvA97r+B1/6duCmHIr70A2cPf6uW3W6ML91bGKDPpq3EZx8DMv+7WfGBs4SG
jt7M3cWXtnz7l83gaHFRZ/8OvsAMeqfs45f++z8aL9nhHMaPcWnLHGMcfmSC
MK5roWJxe5tVghAy8Kej9TmYNzyUu+CCqfyAgemniEBJGLBLvkxFPw2aO3fc
SYLJZCFAecOJxY8U+GMwtoucdqYOB6uX2MTIrCUo+x8pHJY0nUyMohGKMQLx
/gt3+mpHMzh8SprPIrES7oGmaGNS78FVkjZ8rCJeCGxUcT3+gjeKEBwOLwNi
bRr04cAwnhHJOgg5dMnMPLZSSc9GYT8XNBh2IwuSpqNZ7SWoUiIxZKw5O6u/
GGi/NzVko0PKAbv/58GGhe9IAFDwa1dQo1jicTrLh0LDrgNqeVv/tg8uCH/a
6QssqtU1F7e/T/+jQhhJPGZOggxemgWaFrsx/B/qmiFgTUTYdQ0nm0K8C8pq
k2VJIsMF2WEcJ6HlwEcKF+Uq5ZryXHqNeDYtAakS7Bhzt9pfUx3kB65dnDvU
plCDc5B4BZnHb4hDBdaJi4j8jfzAV2jiyMdmwW0TIu8BAQd5Sop4bZkcd2VN
XR8xTmImIH/wqPA6uFpWAI9rJHTwTTo8WqJvE+dzHMG9nAA2J6BeK0U9APZt
D+rvz1ybPQfw/FLsFN1acxdu7hMIrvUWmPct4RsDifJQ9MtT5Zy2rvRgYiL2
bIKHGIJt+z/au/RF1ZF3bMc9zFRU7hIQjzPwTsvDAlavButbCZQBk698uy60
YuD8IdSXXYEyw55SgGoR1+t5VcipjXVkL8sJ445joUCsiqRKUhqOsHezt/Ik
vY0KuWtbY1XmvMnO+ztRyUvQOYuF/QLaQotTCaO4mvw0jfdzh3R1N+ohs2yh
yDJmoNPwzHgmxZ8wq3QdT8a0OO+Wd5PUrnyXfYgtsdTV63evHFaRwPyi69MU
ptIXLUmQzKmsceaoGswGB2MDTp8/qpGnT4FSl9vD3rok5uNT+fNqNZs0Y+DY
uQUtngTbOSs87IcyDogELCZDAR/3pM/NAcf+hQxrOIKApmwNFaSnr0UNBeiU
nDye1sLLTAL0fIwqfQq3U4zLUiMS7Yfn3XZ0GGtdQrvMs+wLusVW6Wuw//BO
Ayvmh0m5IceVEzasTkMwGAoBNbYEKaxD/lLkX1qGv1p9V+oOQJB6988lp01w
dzrhzo7XxW6z0CZJGteww5v+fJj30/JY8C1si7cYTf6yuBapKdN15D5yAE/2
041/Xs+BPpzLOhGYBpwG0E09sdJQxSLC95Kxv74WqPIiFhJidr5qVITGxoR8
eBu3zDXaG/Ecs25iJcH9rXmWYsyrLUZt1mnjIcx6SMn/shcapG8NElc72P1l
iFu3m4dwH5jjxEdvlyMfhHBasXOmEUP2Y1W+ETyX5s1Fxw2iPUFXtnWJx22u
KLyaMeck4V+Q1F0iHrUprdQclockQtUiHnG5gatpyG/6mMpYOphBeGr/2uzv
BCWEMqMl1YsBYdN0lXwUtoNav8rrKzH5nTIstw3T3p7664PzyA9LUmg6Xtud
IqlZHK3a+N6MSY36RcoGNM295s+6PgVTrPUwomImevxImRJymWGlq7Atfaxc
nLMMgSsgTKaAMYgFC6BysadDayh3eZZ8atsw95SggSPARgKsfkXWISpRM2iH
jDo8delo97PAofRfDAh4JIoxvQixYSuOCVR5xlqqPUXKfp3ckBp8bDfcPbay
dF0NKgukfuqKjtwapQH/TCpfhcb+hpWOlj1dr5aKZfm0Wh5B5D1alb+d/Bt4
N8O2d67ICKZzRBi4iIy8/CuPdBdXb2dYcGi9RidODZDW9qCUosFqfrK5euWd
yw9yDBuS9uk1MhoS+7JDgHhOzA/rL660QcsRRHa74+AvtSV1GvLiuga5R94p
36WjMs75Fd0gjaitV0ZMUkN1mGs8W15FBXY5Tm5HlSY78ze7f+DcHNZl6n1p
TXAODeBPsAJ0pEsL54KABGn43edEMQIA80zG5DrpJLSfsvjtUZk1cqCJkqiq
avUdI7F4xvYV2+4kGEKy0x0RG+SprzMJdbvDo9e2gbL3foGRqgJjoK6eM73r
R9z32SW608sYKGMZei8Y9hpCDeIzsEl2BM9DzSG72L5HtY6E9Lv47i6NiiWu
GUtBThc1kyThdXChlo8SSybIfV3o9iuRDTICQriMRsvwQ+HkOWF0B+DyRidp
LNA7VDDwhrKpd8oWGw5tIdisFxA9afMKfAEmfdIm60/XP+YGQhYiCtpT2W/w
6phXEVfQWhqYEswzGn4J6xpY6s6bgEFkkiIKMsbIvuOM4Ij0L7n2gpWWwRuU
LsD2hrvUvYjjhSRJjLDA1RjfU6yyf333ShApwPLKqJGj4+PpnoVVqx9EN3jj
3j8+Lf/PCR8ID7rgvTfWii9YNVgt+GSJ3CNhdMKdJhHTX4eyqSl4w1ZoT+G6
/ogdOpI+hCtO8gqK+EBfOVbY5s2yKxm9WqE2e+nuWWRipnmQZ/0BIh4jpbAG
MgcyAKkNSDg0vsgxfIWjd76vmH6fGAsD9u/exWhKYGqWjrJjMPalb4uymUv8
Wv81gs9ZufjsRTu4Q+hlzICzWjlzNjPGGANPPHZRc/Krz1ago0NXwvGsSvBL
q11Yv+YK4MGGmz1tvwoM/+gGrVbZC0uoozFWYk4aUlYfuPvMPxEKjoDibf0/
OAkgi6r95wuK0sefGthBKcYj88JhCND/e+LiD+gJnl/4VgimkSZj6WWEVj34
oYWtAAHzPPl4quzZVQW0WsPCdgZQscf7ph4bFjpyQsUkupWnlmLb0J9+At9/
PAnydd+yFXDKHaQyHJdiKWyxX/5Yf21beqVSj95usHYdSs28PthnCLaMZgOL
jg3NZysc4O4f7856lLFvcug7ub+MZJQVkBuC9p7Lq+YbJxQlgAu4PlKNYNyq
mFoyiUQNpcazfFJsn2mYF/eGpccfTh1JsLwsaClwT2gSj4Su+lraJJvzSGNK
0mD0qtuIaRXlOGPkfcWlmzYDQK0rwOY1aihJfhnUscQBMBESqDTiHl53mHLU
3mHpX35pzkV7Ib4KBO3ZCFyrr3fRPksRNKGhaZ8H7gjuqELF6fKxBTEqj8gb
Po//CSgdMztsbCJGvkI+s+amjvDAeBW8B+xfWJxinurDNZNDhpcm5b0iYHKI
3bY0qVX5DoIlC48eGoqV6FRd3FAck9wVaHsL8yeiQBzuKDWaQ0Lotzp9IdMG
vfTJTTd46zKfcFH0R6V1Ukib4ZNyWMSoUy8cuLhbUmwJ9G3L0ZZqJ7B1xNeU
agVSTuHldq3JE1B17p2npbOSWdaw5Yig9qu5U3ZVkVnW1Y/BzDw5pecsgkGG
1S5f2Up9bAE6t8TqxOUf2QJO8Fi/IIy+q2Dk/6D91yI81l4k3rMYajAeR95Q
+ablgi7kj1YALeMHdGZz4cCUQwk+T04K9/Zu1t1f+QFeousXR1o5pnzwBpkl
HO1e28C0HsIn5zImilWkpgR/9HwGDuKd5GQonsTtOFLexK4+b8fXAe4J/l2W
sUP2I1/7sHRMl9Y+jkkCDj5T05Oh1jUJVbAZUXNTKjRfMgMy9VZyHgIUhiLu
kkooqyokYf53hvcaIoFxdVlYXmG8XtdBcKt30Lp1UgC/WVueb0psAXHPcl18
FXQgjl8/WI1v29HwB6fUqZXw413Pi1DWJi5OudpZM8nGfHE9B4xfoKI/7jyV
KDOZBTQml5ZZYDdM5zSdb/bVeayhSZjHEG+5eQsISLO9DX4j2iptJd4xDBcJ
RyN5RrgMb/a9ZNYW/7Lh1SPz9IMJsoDs9rbsoN3meYr3jPRoDbTizd1mnn6p
/zNHTzx+/WjdokJ8Idwa/1Fj6sl+8MsBuvWRFT89s8D6NexCTP50wwEsBn90
8/GXt5N1kugB5EZP+4wz2xgQWSa9taVLHjTxpAK02ksyoMmBglBWQDZIp0Ql
3afcnIkzFEacY8Z8EnP8bHAbllpRAS4nlqMaDIn8yfHE7ffz4sqz0YKSSyTy
LnAMSgcoO/T1x/+7wZ8qaoQ55xnIJbVrC8I6Pn9JlhRwJ3CUznI7AAOcau9a
P/+mdJS0nsOIMz1s83ClQeAT4dYcEZudR5imzPwnk/3YG5uMuE5tjDxrE164
xlmr43gg2bCpJW8/NJtr4LejqSg5PpK/+MWq0pKKUYmdvyGaQZnP34a4uYvD
9/uIULDVtn01VDbfn5rhwnOipsHM/ZlfsNdnwRWbt7D6hJItPcJ0d/re4hz6
TIpH4mPnWIDuHrzRtVR5KHrYwhNE2AN0iP+oDYBqv4tm2fuhgI63ZPzqmMMs
hGnowY16wvUEDk5eQ4N7bqSFM7HYv1QUrWULBXSc117oSX/bANan0WI3QG4T
o89890A9XB67if5l7C6kQDgD5h/YCvplQMhjzmj1pLeYUF6s/9Zq0EQQAsW4
BKNeFBRL5hwLHBBFfYt5E+CAeduEOeUSImoXHjnUoSfEQ1Dlyd6k5QLo+c8g
p9ZClg9EVyM4Egt0SCxHzkwCif3o5Glhu7wA3yJULIBxJlTD/NLJXa46UbJH
hnAcRpp5t6OMgcPXUud+cbauDk8Wrzt4tLbYvZk/J+XdkEML4c6Mjzkx+k+K
EKLdAXO9e4rPBADI0ZXAucQc4HQdSx+FhbtQnKgpt8wRL4jm4iQcTrMf9kOx
3hGKzBQtWqJ6PlHwC/W7T26OvWJTYKZ6cMwY63M6x3QpA59KG9d+SPJhruEN
FgTJPjn5o/6x6Fsa1UsSo5T165gM15aR76CxEDCnzIO2L/rzwb7dicI04WPh
dYGY5VDL2CwihYjIIYNEGb5VoxiLjDnWI52nQhP/sFiJwmDFQOrWGa1JHb7B
95RrO/42XoKJp+hCZM6ckONYCJ4eb6uwlvqzrVwx6PxcS16XDMFBlm/nkCQT
z34NoAHhW3+oetBe1XXxIcZuHonJowInVqgSUjUf3AenQ+zqMuwlE80lRhfY
wMYYCK5YFbzca8ethFGtYiXmnAdrdN837E/xaU090cStIAbRQYwGq8bFPE1B
GUwG8oBPk8E4ADz6neYoRYOR1avBzS31UFJ53zizTbmCLXiw68lPseDRGLco
XRLbzgMSWEez/IaTbMVkoGN/cCK8Gen5D6Ms83SGqy75ZmW7TNP3Fi/biA2P
I3DjZxzNm/y4tE9F0O6KT0jSSzOAqwMN0kI6e55Wnzve0YKsdQggGtSGnWt2
jk7hGN0jYakhr5KY7FUAoWAcT559PXStpiYMFpa3JTCzg6LJjqwN+4+IRmbD
orYaFjAMob0Ssx+vNs+P01OnwllCJikdYP1qzfT/KG06FIag5F9ueGu/JY5U
MFPnfcwZiMnFz6AqtcF9vcco6WnKf2vYWb4VTLe+Cn5tm24tpiXSkGN3fxGv
1AcHKlHcMnEDKUrV/CqZqDRB2+lohFeN2Y3kGvqVBVo9vLDbr1ldS8aXl28Z
Hri5cmHZ9DUnBqvHBkqrhX7ZwolBVOHNGZjOoIKAEOfkGUlqPgTb51lk/jOM
QDzmkm+NL2LQH3y/QCA0lP/mFT30SSyYJZIMLsxUSxvas/hBJXkazaHrVYMz
VcBe+wXte4XU/DU6/MbAmh3xPCkomsbiFI9HgiTheeND+p47RkjDaovj/vCM
LPkYjMP53jzy3Qr7cIcwtmmkk7OwDp+eqjUt/oJTFyJlX1hjsBSUjpOOZZ4t
UPC9ql3gS2aCftlDGVITXMOtCLIm9Dx3hT//cZlaPA/SwHv6PocvLEDcwFUu
H4xpZubAo5n0Cbre+bZ9Ipomaiq/qwEZIIxResPI+yjKUaOD8adPBY2AYm8D
hZaOfF+zegCthEajBKrVAx7+ZgqQEsmgvXrUc/IJrSiyAzGvqzNYLGnU2F59
4asrEIHg6cE8FcakviXY+6FyM5bkaspQl8QViFe05gGa2m77APN7BA7mAL1O
hQ/cRGKc9U+frutDLsSEKAFi1rTwYavX2k/9+fM7Lu5R9mYASLcdTUdVD8vs
dQUuEM4XgSas9BLSGVYgQeaYhQJNswoV7xKsIAPVO2wnt3/ExQDAg3IpDJEZ
xd02GyJTqH1WSaz/pZ4msYV/Via4C6lcDGbjeWX857m7AqMwQe8FxXwZT33W
Xh1WYe3bNZRsGNnmmkPoRVKZYfENX9V7kbJ2FecWbaYs+vymYSV1WQANSD2J
PeLWuBbDh0mFfovm4cylYPLcz63HYd2pzv+5OWXETXHEjPPsIyqqjm5pc9xW
kT3l9OHMM1/+nlhDruhgixcxIxeT7DBZ9zWXuwUaLkKcikdUMGYmKDjG2b1b
IKTLLZ3XBQJ3jmq5NxBYWpsn8Ky1nJNwRI6tyFvSc1qhVToXghshBRoAblOJ
PtQEaTVTFz8t8h8f7MFKyHassNg5VwbE003iWKPdXd/Zw47+X/4KCIbGhuC9
AstIUnBA4//whsBjjOil/IlHVdInFQjaTE3VW1zpogwzpif6iF4XmqG7vFBt
WaMbJYZm1FAoW2CwUB3FIL0hPkCSomw98besvy6fRQ8AL0gzB9JiOfpPZShV
JohBkcmtdb5o515spME3/B6y23REnpCTu4BQMiFC0GKmUlTOrqOJgPKT+EzU
4FnSpLXkf6+84VO1NCuBv0MTzibudML3hCJBoZ7V5xQaPFQPaaz2664fjDII
tfCO5gdGpvUVYbjXtMhcbP1ZumbiD7mt2KRw6qg7r7DdXF3+IYJ+rVKbmmN6
8p70QIRfPsXx1/tqgAb8SCWOs+5hMHhfNlghkAH/gFLlmq4k8Y5/PDyuEf8r
CtnGeW0DeHtk63GVsUpp5ZjbddQcyUI5kXlPTusQ/qrhjroO9o0fEXgEEIhs
rTBTbp7uk1nniyyO6rmwgKvK8PY56vxm+J+M4oYlxghAEeMru19DPEretnYv
N1m/FbzrpkXzl2ckFXmAEF4cu/Qox3mClHKCsCb12TILtZ6PZcmeCoMgIBJO
/57bcA4C59MV6G+b2ibkVyU5lwOSVgSWHA8DnbnuTkpJLsBvdpzhS2Gg/bmN
Iant1ZBLtnzTMkPccbm/jALch9a0RSvESq8Vbm+UmVx3zxzbq0MHqEoY6CKZ
9Mq4pYOoLMnZ5F7rACnaLwN4BxylHM2fyi+40lsV3pv3w0d6aKtusSF/A+9C
1/e+1gf2+t+edhdvsghnqk8R4A8j2syukIpcJEqiGUQNHZA8Dbye/jixkSqs
IrvRapU29SSQ8amlAXUrSoz1JyKhhaKKCP79w+QmhhztLOlIqjPY0caLSY/1
FCFQRQodz1DwgcBwfbTpTzlcZfuRW6XoTfDzRICW5YMEzsbepj1cTXgqMk6K
lOOSjrMMosZuiR8/qN2loYhAd/S+aQGgunQKC6qLfM8x4JbFE2ihKnoP9vZL
3iquva3JneHutD871Vj7B2O2/JeyBDFYu1zUBWm3gSHKrWkyGkXumIqa3v3b
0rf5d3RBIUtMLIP92MilBNslfkZsmPPCtFmU0nAo+e58rdfQsU3xEbixc8aZ
e73bL62aivdL4GtcfJRCgZbPMGGu1E5pjZZHrt339Py6eLFG35bE8lFkcPeK
GD4SnVQLtexpaYJDpo3CnOoIqNBF5HrLjA583/R8Op6zpI5JmWIo5xlXMxBH
Fbgavc4PLUIYyVFcbst3rQ9ae+9O4sBB3SYiDEBBFDt2dX3CzAW99U6NMTqd
BJfBjjlmrgbWfCksy7qH2K4CmLdgBK8eH5pf+82h9YAxb7olFKJieepmtkng
p/oMdnktrXwbJ3620wlCR6VKx8EQzGCD4C18HgZuUGUiSSCke513syYmrLym
k24d/o6t9f7NfPYFLrVtUHQvkiWiCvW9Qn9jvmdFIfwbhGmE/MmQ1jPNEBRW
gEVP2BgapUVYgtr1gjwo2qIeH3V1L5q/6AFcaHYky4YsHXbuch9hW4Q9WjR3
lU9vZXdrSOvH0W8/Q4gUM5Zbx/zREn4uvY7afPG9LJ29e6/t/wocalslzITW
xXOkQk29POVMIQhh2KHpaWy9RdikSQwfqj2pYEbKlup9c/o19ZxF2r1pmpQT
qiWwaHUnjsgAXCDqDqyKDGBy28uM6H9/FW2x9kxDjt3soT0difcQqdZT3rZb
wDICLQzkHEg7cVXBj5rWoPDOgzHEYdSLFEHuF8YTkTos476YtdsXGdJRt/c8
vWqFdc03jKQaKkB47FTjl5OhqguUGL5/vFd1VjU+BUlP+P1XRHahNgN7zZmq
tNQIqxelzI0jG4XmVRUbMVkGGSnhDR2yixVlyuYq5dNAGY4ltI8mEBx1v1fb
ns3wWZRYLe92JICPA6/Pphrinx8k3HIarOko9paS0FW/zA5Gf/GkSOncQF/l
dbeinPX7xVNJPAlCupwYKRnt47K/PTKHdQU1SY98OiF0rD50uSuAbyggueuQ
MD4a+ykV++diM8O1v7X8XJsWyopv1KKVcwpHB47Tb0D8p8VhnVCnZRVa0O2F
Nko93NybJPe3teWneX2penakanGT2JsHFHAkMgxkyJ/czkeOfxlSCsfBa0Ph
9MSYOzlkUn1oQkxx+XIpF4bSXdNrIXb2iATijqnGb8RsV4vqPWhW8/pPep4G
t8FcREDMih7n27clQbRpDr6yZoD+LRHffVmMxlVLU5u+Xk1Gen0F/XOgFCwJ
oGTTES6Ou1UyMYg4sPVg9nS394TppKS/un6t9l9GLtCXqri7utRt3lNSGCB3
XRUI9SeKErApjIcjBY6W4yMeCaTvOJT2uXEpJNr0MpduVvg8lyWzJ0HQcLfF
9TwTWEV3KdEB/K+HjxQfl/fD70IXAMRychPKsTYKChc3LFIh/d6+UlIzndkU
z6S6QcPNWw3bWya6VwYGWlPyzMKFCBNTjFCFbWzuz6hrUWufH/T27CrrAUxR
FWmiZCBI9OTCioZdoOC08LzB2IIj041jKAX5H448SyknPzrgnOTjsNrmGJqu
CbntXaEehWdeeF/3obRs+1/JHnslpxIhQnQ2VWnh+GWwQsvFuBsa1zCN4DXS
Sx1FqzaSrG2rV28OXjLh3Nvtnd3/zv98mOyrRjCBU4nIbO3wbhihKbPw/8DX
m14eWlDMTqRk2xKCiJaerGmhzqrSho5hIB1asr1Q1eBH1BkfCQDJdqSzQmyJ
1sdmC5/o0fYbclqJJ7AzAK6oviGGVwhOwMzAGBXbQeeiV86tP3fqMIdxniKm
SfQOrWp0YBUxWzkg56rD/bnAVPy4GYvJNMW/cha8fBKOrDPGGv+7DL/u8ILq
cvK8L94XmFt4d3gB1MAuIKGkfwxye1hqjrk7AmaBA1zW+K3k64k/sQOBaujs
cD2sgGoXu3nf4CyCR38Q/2CWC1n/iCvZr8ShxmMJu1CAt6gJx1RyjE+Opnsv
Ge4MVbKuz5CJYQ/KXW2klRF6dOsqjIpF6fP1igsc8e0ddS9n26xSAcN7obNG
9ikjFVvQ42fOljbZlq+59zezZJQP85yj2jd21O/qM4rxbv1Q9+xNqUwJZ1YN
3tMhaBhYf3f2YJ0p9Mo4ZmSxRn+g/9SJD/Qphi7z59wWOS4G+q0eIaKnl/NF
aUCK1oerl8gcTh0wAk4GlZtToRYVe6FX/8ZzGJSSCE5bWlG3JrhARxwrQi6z
RExvd5dFzzLrjAMWj7EgkqWp91i1ltIVwivAnRu3z53xrONogf9jjdu1GY38
qNseZNyLYJ3wHCWFEfCVGcTzRbMoq+/FThx0fSYBvjRLUpEOR6lzwWiqSy53
Npx2CUCSv6h1ssOVLFTOtNpSB1dLWNCR577yR5+NqmpIc8xu0xgTEN2fLyNB
oXrecG5rXlHRRyj0ghcqsMIF/K/ITr9gd7w/c9ruXYQd3xofpaQ2OFKBlzbY
8oNbGmGVCImxUjQ7Wqlit6kenngMtxUzNsuQldBAQhMWm6BV379rZLz/j4vK
cFL0d0kUWHzXsIwVSb51aaN4RuhEkWl6/UdeZY6ddF/7mkAdjIo0XnAEkNq+
0bu0E9RTOKPJHeMD1vpAe+rPywXyQWowHFGTx35/shrowaHDVlaowjvpO4Vg
l5QygENNlg0T3wJRMJZwES7EACx4nbMkmIEurAAanrU9Y9BgnGiqnogQBddd
9dS5YihOKqd/mh4w3LC/YBb6go9qxjl8HH3EisjnxiiaCu6BLZ0LGu9Zpd9v
JmrUCEIu1Dl5z6+r5k0qmjGfqur/KOzEuhvCHlcRyd4Tc6BEYOQrzb/WL/GZ
cn2v1uaMbTxQJyWF6IzV2AE9UPfLLJniFu/QBOOWBQ0VRQnPCospHbmleKxj
SdoNnbQY/H7+0J8wj4TtwaKNEnsygp+XR0WtmxWwH2uhK6X6X7uYelz0UK/x
ey4GErpV7GXfHEkR4PWzHSE86i/0jGVF75+pp2XerJZgDIopmRc98Y/JEug9
1vghG22aXJZwnObDDCSxpo6gtC+xknVdyyig56aeFsAbcnHAYF51VNWebRww
jlzkhLxCXQDw/FXmWP0nYqqDGy3nWI8IQJ/S8N0HATGNvyaSKue0gFyQw38j
gB4UMsLWI04xiRIbPwOuYE8oQ1ZokpwEpByWslxnJdiXV+ZZbsW8w3vpV71X
M+ol5mjwjV8qFWWoLhdb169V0KzE1WUrvxekI4WEmi0zhObbfcbH+SVJ/xoe
Cfvnq8YgthTyY7c3jqIxYP8Jo/1OIZeA27xc0qoKg0G2+Uak6p07FEYXNfmq
x/4VvMXI5Kvf2XF6y/1iCx5uyYglFCz6QZWJo4YwCZoEhVWJciAL62BaBaM2
bGDGXqXJynPjLiXbw4Ty96OV54tK4PtmdK7jvrKVhoLPr5tNB2Ved+iwhi2t
eW0YlxkvYMQpl6vqOW3ArLVQkDEHygSxa0tOT/4RcY8N3r3hTF/Qpz2oo7IB
iTLk7T6roeRQvTlTJzCqqq/FcUKW69f/taMImOdyQ57ZZ1OhwuL899SkQgpz
ca3u1UGIE+Gu2BfOm68VkjoThy/PXzGPdDHi0hNxMkAQiQgXKUhDTXdDbme1
fqX5OpCrELjg7ACJoATpL7Ttr8GapIyW07Gq60JYEv/pjWOM6nUC1apOERYn
2NI3DHYq8mOHZ/d/czQ95VgNX3mk636A5zIB/fu20FY9ylChvsfTXh85CQPT
jsUlTg1/VxjoW2MjZs7dHaYxNs8Oy2ZxPfvrQ1+yocva4cbKym6FXyUU5lRj
CHvyx9zRRbJonwoslBDNBIrhF2nRLnRCx7bJ2cw7ovx7tKSAh0Jo8DH9xkHG
9lMQ8qwTXW5vl5fGy7lVZVg4vF6+FHqvVcL3GBGI3gVZnJKWc5O19wjqTi9z
jlXCDSo6ucYmmpC0+LPSV7zFW3VlbS43A5ffnPS7Z+qjCEjNF7Ni0YdvBC+8
e7Lscyx+/uzzN1ltMMDmlt6I1EgchSscUI+zMTRsN7ulP0keOP2GlPZc9uJZ
81bY6XFt0ksZvc0bDyIin6k8XCTwrSoGu3xNd/rhHbLOQgHpO7CCkOgECSPc
2ZSpQjpdnj6a0wp+XuMacpGNlFjP03vJBdpcRyoAgC9su9KaRAWHN7cIwLRK
zAu/EmQmlyMCZ6gTAG2OC9uGTHqwbKiYizQs28XSnShhj5X5kRFcTEmdBIm4
r+0OLbTnG1Y4F+qxIL9eNv6sRIQUYZqNX7r8z1WbG4ev/tMZkjSdLd7Rrhhy
eWJLDQMVyV4z090itBS9r1sfb0+2LUfYfd+OpT46cN/+FN+fv/z3VEKclmTA
pjgPy1+l5xpNuUQq+KKUTijIg7Ditey4oFO6mRMMkB9w10D0I3rClvfRzumI
8Q0IiSO5Qjzctq4juq3J8r2VeZlu73jKwYq2TsmYhIY9U79hwN9RP/43Spn+
tX5tAOTRnmODaSHNJfRkUeHcnOV6dsvozKYk8dX2bAxdUwkmia9+FpbR5qJe
KdKjNV478YwdU1mJFdCDOoejK/H5DlV64fjqfVK49WyaylelgmazzKKyimgt
63w4m6AasEhsiJoqf/RZGIp2kKk/c3v/D0ISQIO0j1FLUUDBHdQ+1rZTWnyp
6nj4dWfOPrlB43rtiNJEwjpK9w1Ii5X+NoC2txYfYJoUF/sOPCYHgnJeTzGN
UhsthCp1407pqn/sPHYI33qXIMVe/iMKbyNC2LmKFI1LGWlBRXz/8LLRux5r
KE8aOSUZJgeSHfZreAaWrT+6mFlz/qNehls3R0zQSJ/ytRRR9dLi18eecBR6
eqYLt66SHVvgO0tLvB1t5nA2kV8qVIn4KYNoxYpFPr3EJKXwFRUlcS0zkhLp
vE9ytWrvomnnphRL60pxK2bc2K54OFal5nHc37t4lQ0MVUE4FAkHj+8DEKXv
YvNwQaciBYssjFdFLBP1I8Y9L/D3Du+H2zqWaJyM9N7jVVw+1AI+CLLl998i
l0AYbE0XU9Xtcn1zi1qNSMUX8Z8v9lYX9adH3Enw/PtDgxQ3/S9eLl1LindD
DzxYix99RaS6CM/TOx4w42dp+KCKzL4IElQLm8ZnhuhxOB6R9Tw8ixZYoxbP
2JSTcZibpdgB7zVileq0dcB5o95W6r4Dv0+c8pFhMQGjYB0BiH/eLcxWpfj0
44lD//M193wQqfjQ+dI5gMkQVbPrBvdRcAyF8ytiLK8RIs6+AfGxARg3GI0E
ntsVOiOjLSzRPRTFlLiqqsWyCbp4od8qiO88T9fd943hNI8pd3w9OEjO7xCd
SfP62DqhD66soFuzUjku94MGZaIFATofysOnsQE5xqtA3sR3PFx3wvv15WhN
v2mC5UPTmShhHYuVhZq94OevqdTbOtUKty07L+0EcM/sHD/v9NjdzjAEZ+AH
bDrclnJwvgNLdoNLnlLI9uUo0UKIUgeE8d5NCBRbmx00hs3hMVT3xzH26f92
H4VmTjkvnzcwWjsjDNIrbjAXUI4aNTpTFxFW4NAlz1Qx0HbyZMwxIoGyb9WA
Vy9aG1q2cKyfYvZ+FZHIZ29ecELBz51zRO71LpZf5uXM76T8vaZape4NrFgZ
VYZTyhIEcSHouKRRDtad9uaj4Jg6cZN+oXTKZ/HBMKzADSXV2t5Ge+nZ7SnS
EvhSscYhhX6lC2Lp0fC60cH1MTW+P8wDgI/0JtIMD9veKOt9P82xYojRYG11
i2sPfeSTeO/LAve7vW+U9lfd7QJuN6aTdoyjqNvdPa/BRuUsr+jjvBZEk4+O
FEL2Lk7EjOleDORPZQOjgAQi1E/Ft3/sSc3VDI2jgr4dwRjgnINTWM9ecuiI
ExHb/NxomzU9y7Rn8vWWAtoUoc3QEGyz0YaXKbx1uc06gZKM/r1d2KEIT38J
Lk7OG1tb2kPZup/G39TL0XrYVNez2fMvbVPpuHbntGI+7ddjEp+NKm8G6bEU
nlr9jJhjKs0mjLf/oHW2j8xszFT7cS8JhRMRcGyAyIzzkiSelLht8LasO08q
EoRelBE6L+fH402j/M8xa49xXN43IqPtOraBV7+2/fJoRcxM+Yctww8xPXk8
KHgCZhFSTy4ywgaMHx9Coqu61wTFnjOhMkuuMXa87qXKAppYfW+o/sINck6W
N20bS4PqK34eFeJgy2yuks+e7xs6T6uv1Tiqg0PTR9VYzDuKUD68iwhGCR1C
O9l7oOW9Q940sA8gMM2ks5WzUNhMdqij/qvxgXcYvq/dkACVTwh6vWoaPRYb
RE8jBbpI9ReynbkP1WL6FLJOoc0nzjZyEHa2P95iS0Kvf2Y/46221eet8NIE
1B1x9/MW6Hy8v/A4U40x1hQMFQh25ruAL4nbcVjgqlVL0YOojcPDnJQEpaL+
Tn65gD5m5l1lHKjM/9CH20peaSM/bpTR0vnyKU6jho40qfrrUMYxfJ6yJkhw
wrUmw9NzSrQFwLpT+5SvEnfvaZufnhu8z4kp9Zuojp3bck6y4IjUAYjG3yzm
NvD99q7t7qDF2jCBde0OzYXE2QNNFEvKXijiI0ChoitZBNQ7id1r/kfQfZ3e
1laYg3MsgUKyU1MWWYABtBbGl1f/EnMtqDrztYQ9QxV7TedyV0DHRyR0aPZw
z1awOKujjA9Ud2sMMCy6+YjRmCSauDVaPnXG3AVm5izfDQlg5Pw2TBzSjZ5g
Zg9NNJzLVo+ge7VwJHtE8np/hpARljJWq4Ujv+l94zltWERr8Ub78C5nelCz
2I0M5BFvmN9LXhhmyo1ICjizs9UhfK090byOPZ595MNYz0lc7jrDaHaqQM8p
y2TZbq9jJBVSN32gjyEUXM+YD3bkA0d+/qRY7r0TvnYg4rWtUgMRrPSUOPSq
eMwix2Vaq4QeJUTLIHyBlupTS7uvQRb419JxlmAVUqLLXPO7MRGia65jRwM9
H+bKvkUnxjsZi9OjqvuVUKaorivqDp4d55fv6ChbA1W+lfgch/d9QQ1HqcrT
AU2UUhaPVJh07e1L6L9gipTOMln4HIeKBMwuyfkbRZDfZ+6WM4CTLPPqdYH0
Dntv3AwWjfpRIy1MVY/eoQAjYumViTwQYF97vUsO1UoEXpjw6LvVsrPHBzQM
Ir8Akvj51BKOMr4oU5C5wUSqg0NJ/U4BZ/BVbMro7V/ZXdeRgFD/IoVKJmPi
dQirk960bef/Y+/1Cv9m998bolAD1hrl3k+5FbbREifHqEJJ0ynjnn20Msuf
BseG02DKl6od/sCpYGPD20OFn3gmVchxnM1AK75aD9tC0dt7CPOHa0PaeqkM
p59sw7GbhGy9W7pBFAdJEb6I4bvXceyffP50NBhddPvHOVySbzG7r5LsFl/m
Lq3NEE0cPgetPmWzBxxEX7e9tKjNwb+msczSNCc8SKvftVDB+cL2POsuU4oK
vyzbVBs5KAYfm593MW+EAd7sZ+6/ndC18PZTpfoBCGa24m87TWxXjC+XGr/I
49VKIHDW2XpCR8EXsWKTAqYxpUiaLSw4y5CmGN+W4ytuIV9mfDFkWJHulhXE
yLzdOlOgjVw5D5L5WN7NwwrovVN5eouYNrCcEj3cZaxYKBA6nVlp4FaTjNu5
go+6yrMHtYSmdYJQlQdVOscp90JaViH8UAIxwsBpKLptrmwT6Vmrl98QtFFa
wNuTEZsM108vq6w6vYF5h9MGf92OLUelZYUnO1aom97TPgGKMPTrLphNoJNk
Pql9vGEqH/dJ2AS4hfuXGZcz5fOqqDGfNDrynUD/mymHg3qw5I3oamliYPJk
PdC8V/lEYcGR+OCKsS7eELzsiceHc0HhTylqt4RQOYH2moQEeEYrFvoH0qlC
c00l+vI1azOndELgrxag3tb3CezBDnBhw2M2ND740czVjBh9Ouz+hoXEBJHq
Tsi9uo1gPxwFkyhLUu1qOuTE2MawHEyJYJ/xvdctbJzXeVkXjjmhbv9bk7d7
QpWnamtaLOExmdyH1OvmxGVDE5R0/k1WUhrX36P2wijHC5sZeiHBZmhcAJmm
43zKxGWdaUoMoByq9OdEzoVBQI3mYeIR/uES9x+38pla78vHJeZHdcAxtT8Z
RnQucpJkBGcJDU/bHCgiUnSL33MO5NPdixvSPL4U7hGdVE/hhuMAifBJy71y
Z2BPNUOXEE/A4n2UGW4o2FmFNkcE2lvNU5o3v8H9U4KoE65C5DFZC12o4ffY
WoeKUngmYvBzdBp0GwuDJy5Je5PUQU/GH8DE9j/Ej0PGJ/QaDGs3QeONKLS9
2MPRga0v9UBQd6Icg5jBb+1aLfgGlPiWUQKGA5WT+gh+VD8bt6hbgl2o2Ay2
tll5bV1rPmi2FK/pkRj4J+G3yoLuyyEzfH8GS+D0P+hhI+Nqs6CIU/1yLHuR
MaO0RDuBtzTtBGRSii7HzAjK75oVrJcOJuvLoqK5AhhCUYC8oQYoQJqloFIn
wj8/+Hv9dnqVpp9RW8cWG8G2EYI1vP15IAH4JMRN7shOu0/51m45sC4mJK+x
snA9dKXB6PjNrlKnj1uYeSeSJh8Tkb0ICTx9fhT7cptt7c8l2E80wSxfPa3r
mW8/vjcJqY1AzlsA2LtiP32K2m/bG02ErraGeQd8YPG0VNBxabkpQWJ1lcbV
izgYtlnwDYy49lN5tUDdoDlHo5HKksCHJ5ByJvTGAZMoL5B3KW23PTyR9VNO
mScMy+1Xm9jtVwYLU2lujHKYWjQisBRf4bhePpvjqEkY1UU1u5ATk7Nk/udy
I0Fw0ZHnWDN9RV2g51IR4rdyYNu+OoiLZcQuyOU7qAd+nRL1XcA5nQXgr+SL
Khw+zE9oH9bQNfsSBTIFPI5RAhy7EVIVSZSMjdTfiVlI8BDdI5L31vNZ/JBw
NhpQ1COfDKS+EjYEBGOXNicK35+nDKze45V0O70KGmFU9++xn2shENAYjwUD
JC/RFcmRLxKkBDnPqO3JmS84EDWwqiXnUIby2h0eKzevQAZHfjhfyk5SU/Tx
6WiNTim1yChIT/ElG6II+4A746uw7jktzMPc+59mV9wrhwY0C1ynH5O3frsj
tsH0+HLatu4QFZaMjMw6mbU77MvYr3T3Q1cmbbmRybVJhqYY7d2/+NPgwQyd
uVwZSnS7nLcIwM0NST+xdJsj7nJj/4YdhB7/WBQj5JcM7bq7f9pnNRneQnnS
1wzmTw/JaCJtvnMglPwrkSlBIe2t/ZGkKksSiTN9/ZVlMyd5Y9/xmyC4yB2Y
cA0ECwDZ+Rw0RAT+aL5qbyYR0Bcko8gpZZXx9bC+3J5ATpkdhChnNxj6Z7XZ
EQpwBJjeM1R+EFQVV3O2/HijsWrzIR3vnftf6iYOfqtieY88Oh+y62tmywzy
Ql8K7He+Wui6o8uCCdBxGoaERFgPlvRpG4Esn1TwxoGvhdTsECLEqR3lW3Lt
BZDyVZc4tZJMfGzjF0ksuUbDxTncmnpbV/YhD51FVJToIdV9Vrf72b/lIfcQ
o91m00p/pt9HX1Ekv1GbTFWq1QaXWCp2l9qXA5R6UBX9gvC/+yzsknETt8Pq
bQJQObOnwmtkG+IGkia+eT/gxhcZIOZ3U9qt78X31uUyinmdFHjX2PRsaHMc
iccIIXbJdMYYgDPQtbBNGAxRBFluort2hfSZmnlkK7awEu/ryQS++ER6idDi
NnRsPnhT1wV8n9acqM87WAfcHF2gthDnoG4gbjvxE+990AaxYeDbielgHfdC
6rSL+odWXSqRB6K9KIVkEzDJ8zCM6boC9s+rKQNyNg3pukdcMGvxPUTq/Rz8
o5MUsuqncBFJVH3Bd+8C0rTbPu0PjMGl9CoF8r+X/ewfOgoA6lRdzFsBS5/4
C4n4e05FuuDh8VtwDATWIOlEg49KxSysVdjiypSYwvMJLzv8ruM+8+9QyGOZ
UtW74V8jJ0z39qAhNot3mfIslU9zqVOF7dL1rnGVAa2PjfxC5Iwd9bonfg95
lr5jXPDNm+AlPZzgnSpov5lCRYdXekG2kfQ+8CGn838L7S/0xdeBexjCD9mw
TZKvP0K6xBBUs2Q8A3VclboJyG1B7+EVXn+tZW0CMCoUen94lvMiexhIxj/2
GClPSyKGpDrl5eeEhrbnKnJMZs8jZnuf5FbrF+igUYPvSpRRPiYrNSMaqqHL
xeRJqwSkfH3huKl5mOZeg5peK2Cy6hCxBDa/JDuZRi81njEZEeiT75JCIVNq
tbZrTqa1K8uX+BEquHpvIEA92pjU6HAs3kF8KtysgnZZ6dZvmXRpvY+NY4Gr
hznZ4K3Ucmpj8Usf+WgmuWOOiOk8TfojtlksGJsVTq9S9OWRJUm5GLJg1jHB
o7qc3LcJXPZx7+xi43yhO3vxUFp5zc5kNLCxJuhROm0m/DAjKIqZqmJxRUVt
nX5q8QYBdkuRr5sY+iWuMvHV6XZdp9El2rWk2h0bjgPtfsLaiHtlVE3Av2Kf
GUgg/P8tdorHTfW0l2i9fWQA4WaumGigPquCQTH8t9ichDitVDsOvcFwPL68
5wuI5Hu0AQHEDYUkqoXGAD2iZ70MdRGrTXvRB/QCPu1GTSSsCKhTakR6jCAZ
VBhSSDHcD2pYWeavcTai6CzeF786TvBf48E4Tv00vnaVCij33X7QixveFmJS
XfY2go/Vu9MmX1sepXZ6yy3AHkUrULNdwA0RUJBy3ZFkSwLucnJJEAp0vCq7
d4UzZWHYrestqUQKefJTSgNkmAZTCO7uoWmkw76Eu0iUTUAUY2aZti12ZFZJ
RCTRNtETH2zF9QXssJPRxogO3rnVuUwg/8sNnMbwIhxa8vKisxavLr1x0mgA
CKqRRC6FKdqLWTtbsU/saHyn4rJfp2Y+/01ew+ybIeESShsjNW0umYE7kk72
PJfdILBj1m8dZuAyGlkIVL3beiMz0J2+xzq60mBimaSvd5UzcQ80SBkKojHC
cMhN5vLKTSLVXSxgfJpUMd5SfwMEhBVAppqcVk+Quja4gMEgHwT+JC7oQZE6
JRLdjEPNXunU2kVSVRVXfvksIIeqEJhqI4MT9O2UOvLsc2v5SxtRVv15DJtG
Jx8p5/M21+Ff+eh1RB7JCQ3NhcfN+K/OBy2mixCPLhQbxxovIP7cWQOmeDvz
uc/ByP02WPg5bVp4/NSuI7cyEt2annH1gdVgBd8xKIbNWn03dvi1hqYjipUc
qR/TvXVHO5VJLDwXr5+SBnrS9mrYMnPVxxU7QtpHPEiAUufiyXmC4mXMQ1V8
4NcVv2S6eGYJXJPudQy0R0tgmXti99fO/cCEkDto6y1aIkYhpHxwS6gUNwvC
+OInewKHs0zftkz2VgUAz02UEje4KHke59QZzAkzy8EEbR7cnfUsfmg5jf6I
nF5MMr1ioiId4l4lXw4l0m7OebNMYiFFgw+W0keslw3/c0wRjBEtRhHaaPKx
Wfhq8e54BU5I2WzRmJrQhqv+/Qw+JG/cYgPCMJGagt3HCW0veL2vALgqXf/F
/WCguI6cT48Deo63zS6oihnNzVEGi8L18ce4Z/wMXgO3PvzaGZL4AF8Jz+9+
ez/ocGeAkHo4JfqgPcxG1LMwCQce23WIx055u/jJ/WPch17LeKmEGbOsboJg
bZuNYNTllwklg5YpzjqFHEDseWSXNZDBIUaZsuN0bP8BpYVwka/xg+uK9Ywm
1yPKFQyHZMRkYCdENFnL/TKyKV7++qW5DXvn4b8cRkYAU317xj47vqhA6S1G
sTwLG3aeo7O2R0bHHtkWfpm8Wd878evmnk21oZmOSEroebkzzpdNn/5r/cB9
WlVV//YguMVCT60bFXS1urAxTeWmyqk7sVY1A9kdPaXMzVHsDPIdVEaRicSs
An1kUeTn8gnsJH3LGNZ84CKkjoCbrGqblqs+U58uU0CCDlZxUFMTlhFwOekQ
RmC5Y46lqfmOPH1A4e/WPqjtYBkPSQaF4k4Vd3dx6WdG7f4MJE/N3KZ3Rlz0
TjqQMoz1oyxk7U6zGDJ2kJ+GQfQjyfZ1COunWZRNds0Q9mG0CsEWv2bR0e4E
mnehGFN4a3+hf4a8SpfNCRGL0Nl1Ve50iqu8w5otZ9A8Y43Dbj9gt35rt0jF
vaQV2hR1frTKDAOhZFj4/pA7HlrNWpT3mqlkmUDfzpJuxjh2QB2LUyuGHsLc
Eta1DJruKcMb2NIZgnIiu+YGkPpgvrAudxa3JwfdqZqGy0WbjmdJbzL5zyGn
pTq8RkI95uoBSnL5zbh/ObaQfiZ69/rSh4uCiXo4GdDiazZhMyKpKgmuu2LI
mvYxc0612VCWq1/v66gOIk8oq6zSGkpuWpcU5kac/SZMih2NeJvirrcfOYb+
owo6blyaBorQT08VEZ9dQhy/VeoRJzMj5mbpsRHifguh4bhPgdtNfj9KZrvK
fE43K/ADWD5A7TU+uGPopHTNZYTCXBQO+kYM1hqHx67tso/IX8pDcRAEBgzK
K+mnQw3lBYt9QrFEt/1Jlt8BTpdBxXEEpieZRnOPUbfrIM2nPiSTxeIlAGLh
qWutWvQOg0GEeLgtMsCLJnmTFsm0xwcYB/sG2XNfQelXzAhwo702RkoEsujU
s9XSbS5mgYPM1liCCX1m7Ro37iThSwCgwaLbQcS9bDEa7Z4NzUzX12sG4Q/j
oyFCSzolh6sbwvyd6WsbWrv8rIKtG9i42JUxTvOzth8Q6imdKq6w/HqLxFyI
Dide08uj+JBb/LBGaDqGzpSq9zw5PpwTTXpinVIPBsG5hIzGGC3ZDHWEbYtz
6ZXJ+ydRWRFbnAInxTamNWpsI660ABhp/xuSUWpUPOUkTW20ce+PLXdR+w1g
JHdGmnC6Gh/jepDmYo9mrzszEl23UvGvNfuEiAvPpXLuVkAotpdACH0w0kHu
KnlMNQ3zMce16m16UD1E280LCPUBp7gfm2V6XaZvRjAU2nHp1tsCdd1/LdlA
F8ekdiSUjJZWEWPfK+Git3AbRjncY3psKjVexLXTRhO6auoSdONl/sz9lqZc
hHycfgv6Kn7gsj4FW7biOt0e4+3XyEx0qSQtAn6KRmsnzJblk+PYIYzNucd/
FuSD8a7XEBPdvMLU5ApXxB04wSeIOVhJFasx71o0KrN9Usp+Gj0JOxOGjcQK
codJqKfzeGGxRjukvWNqd51X+B0eIfN7e8WfPix/mCUXQ2BNxMl6ftk9pqx9
dwZjDnKFrxxmPEcTAKYV0V1xkm8kyV4iCMs83gT2SyOECkC+MkAtacxekxqV
bhmtK851BUgiUypRkSvvrZK1zuQAQw7b/uPiIEPBEj7n8LZJO8xZpMFiuzqZ
msuOemJnpE9Hcqyu2l+awnzCqjvN/bIN1DN/iO4+7rTLAES9bdFS1hlaRlZx
VFTqEcfRggnmU1/0DNhK6TeuoK8MAzpXz2TweZiYA2/IGiwZH0KodgT4CcQC
2O6BJHdCOCkRN9eX7Y5ybdc7pQOdjGocwNVig1XCwfeLNXt2RGIxlWproopZ
jNdNDJVthtLckDzJkOnvhWJ/x6gB/9FRhXPTHrUOFq9nji8C4Mwo9qexD0xg
zZ55q/X5C3f6YyGAAZTAeGTJ6Ql7kSu1iiLM3zviOQVwafekZhX74ye3IZI6
OVm3T93kiUXi3rBbyHaogz/H+JLWtoF4ErDi1ipWsPb/E87yg0wMZvlF44kB
/Uhodk73qiR39b5KrbebBe829QsxE29SOb4ffJRHqNM5aI7biCN1YJ6iyzmy
aycJftvfyuZFPd5qRRVsf93zYWmFw/Hx2J75q1PUXRgrS7lHQIYjxLmzrGdw
K2HwXwn4EEvOoi5rTGvgqqj9hK7KZOI2DZqaST2tFzgdRFNB+YHdLkgR0u1N
7LBuqMYaZfyZJI5MB7WGOmBkrcdrhmDedpUgg53kzG2UWAXAG3TKR2D6EbSb
dW/H5o6WgYCVIdm+GV8b2TcRQ/eRV4/jvtezBAJiRynVH75Q6q/FFs3vCMC9
yeGY/yXzyfGg8GYWsgppd71/Oh/vpn/CK58DyidLxW+5mgDdW7Ue4k3nr6N0
Lbqm69igL1ax49Arg3tUIkYk8PG/cHg1l6QP1b+MtQYtnFsQV94QFEL1temk
KAphes+pGOI1flzsCZ/jUfp8kDncRYFGYuLoyuqEKLh207nms7TigJoeBDQQ
XMfs3hnGP96ThqUix5AFxqzwpRizSQ0A/5cBYnWWNDeIbMNYK6jtIvDRMejU
dZtTdHIDkYFJxHYCGakwz/5DluqgdKARjd/TRk7gOL+fQs/jzUTplcd32D2H
yhOd+GNv5BhTGW2KOtJd2TPD8T2IsaGQdzbokCTQ7/ngvajHxic6XAlUkZJQ
L/KTpzlbViwbZZQCReYc7KT3UKkjdXQK6ixhwnoKy24iiNrZ0OxItDvZ3eok
S5m/cWEMvCfUUzpHKdp7CFS4vidD2TDuYPKI6Ab7s3ZS8dYRph41jcnoo2Ea
rOKNVtGHovLodcxE0DKJzuZT79d/qd4iedD72NQGNiPtTzOtCeg6f+8WrrWu
BES0DpGSmmAd7pdveBCIHCAcgGxClVb1yLh7UAuEJv7GJVAvhxniqfBoxqon
oeZdYtrSIiSzoKMM+VtpvEUzcAiN8JJHdgXbWkJtx3cKUWgF9e+qHIoBf2nA
yevy/fPbwq/uW16IgsGD4VbdrwRV54OHKw4QEJpfIzW9cA9WwQ1cHQHVL28N
2xS/MeO06gasjlrjj12SeC7BYM8VIjBIcfylr0qwJCw4cXsfJ0Gyl1OjEKab
GAMGXCUz3d2Hgic2cP3w3oTxoka0WdBjAvkb+QOS+tIaR9vXkaaEHzVQVN3H
Q8XsL9R6VX8gbaU1oyJ9oEItYpISIsA3TPRAfxZDOxWUlSC+SPjsNmVBRZWB
raJNxgS8Wai6kqw4RcykXhcatdUk9mhKVY5d043QnnP2uIjj/wd4moMkdYML
YzBdaHfFXxN/5XXy0cm3QTlNzXftYLsE8WwetmWD0OULq34hloV0lEmgLABx
rDy3QC/Fy22e6CInpra5Jq1lqaFQ6mWoOAuQK/UkzlV7pZjSGliZIjizzORL
2uGa0ayo9Cz/uwaB1T2/MEPHijw4fJvY6GnPQqgHzGo6c0+77Sy5d9WnbqCD
MjNQ6YqQCojEtm9YHmxM+2y02Pdob7b2aJf1Jg8D2Zy7aZgBSPoYfHNMHmgG
kcfx0Cc9hBr8jBCl3x+a3GVEFFMbEMLzAedUH1m5oAgOYpwCRhXfzOoQVehq
FghkOCnEwp8dG5FOGyZBhW5ViG6M6pnhYolwmClXQuMvDTBbQq8LclkoUSj8
0VdcGaZIP05tLXwYQ21ccG0l2UMo1GfamMcajCYZzuUsYDM21hTf0fp0W3oz
ufCw04EmOAnfzwE51LNp1kaurZq5wkk0Znm4CIkmz8T1wKVTET83zvLgN/9n
8VbfnZxp0SuG3S7Xx/cVoOOuD+jRptmrtls8vP0PHcU9is4oSzGorgOmO2/h
GGsDenYI6Cdwf+dBJOTs+pVbapoFsC4ewhd3qeRGHgq+hRklx4xcT38TGw4+
u5pje+YdFqtzixBReeCNGKVwnunJodWfbp2oSbgeNCKPl98PHN/uAjauBqin
AWzb4pruhTyD9l0wgCUoOAEfge0Gi+28ikR1IowOLxCh3gSrX+1LnQHnU+KQ
th7c/ldZaqdOJNsseJzjasVqjD1Qoi1Ajk6LXBesnaUWDzM/5wWeNT/djw8V
XlOZaTNf8gQiOhfaEx0lXw04aBJvCUMp/FTjh9PUfVQd1SPz8U+XcSzYV/RS
ZchBXr/LCMnA/5Op/p527U/AqMi5qdxv778h/ElAUtZZqFKTlNqKPQdTDFd6
qj9I5z5ze/GBSDrOUdnfBQRyOwyHkcs5LshP3UDDlFC8kM7sfxX6vxyl4vR6
8WPjfcc9czprTJFe4palQUhMLfNRh7xFIc/lUiT5unnglxfM4ZlR5oniRXjg
Qfn9FFw7EIvG3+RmWp1C1/G0oqo96J0w1lTVOE8sMxMELLBCJnKpmMJjx2M8
1ax86jN9Ox4oKFHtFdCwV/0WvOKM+dN55lPgd6hDKh5M3SwlTKKQoylMM7He
y6Xv9zlZ/SMsi52sZo9bMhPwJNJ4bqS/bvN5h9BoWFhyPz57nNbKAXMxEYeo
Has90/ey31crAsazHZ/aLopUcd/qkhPywpLQsy0LF8DA6OobeUCYu7UTCo9U
T2u0jhIn4x1hCLHcK/cKkLgQNlX/bMuxcTrwP5ufSC1Ihl989uSpYY1dGuSF
4aA7wOrIJX2ZE5AmX0gdkMi2riRCnqoGD7qfNzeoK5RGZQSN5NxHN5AQmIhv
Of0YQ96qlCLELnnXfVFt2WkNh8q5w+OGrq2wjxlIwf1HWfBwAGrw4Imq3sQt
LXUfo2kZmDC2VKXo5BDMKWgViQDsB6on7qpOtiwzcu62XxXXHCMnMfFUSR6y
9jTPTBV8OTiHLHTOBol6wkOnydq0ORaMU+aS1hc5CzgsjL6q3haOkf3AXgp/
bDWx3Mdu9UNkBOFQzKUJi1uF+L1lz3bRJ8rhtKKqVv4P/gchPw5oJtBT9sUW
cHF3xIya3sBtCx402Hv123KjD8/YY0wPE2lzdC5dXcm9sTcPKKeohNtDgNQ6
xynQeB1tWi6zSSbzFk96WPGM+rSyDYEJgpshtQmUq1x2j2vreMoC/DSop8vs
ddw1fD5vD2kC5qq140qqR6FuMm41518rZcJ+lNByAqs17PfVAvaZVUhQD0Co
uU6FWoqKwNQLLnM3PahMd0QT6S3Tjw/yOTNRpGzdXjaa8L+qiYo8M5DNmtq7
tOcvREKZHnI2qNKTsDPg+HJgTU5+VwU9xuWMHwEiO1Os95oLG0/JOoZDuvo9
xhqT2HMwDV4s6ALlGAuuRixCs3idoVsNB2J0kZ3wyjqUqmrbi9XsXiMol0f8
uYfPZ/XpFwZ61sMYkc7sJr6J55A0kTsHC60j2rd6wafXUo04Hepgv3sFF1OZ
sLPfGv/RI5UopO7ps97NSbvwrp3hch02BVSs8LslENXiwT9BlxomSDtILDFf
hX1CMGJTRXi0lobzaOf1RYbYJLGErDJ/zaxOCOKx+ANygWGA3esnCzrLvaEV
cqHDPn8vLLPVb/EYFFnp49BlRNFjDlrUmF32+68FF41Pu12+4fhjTT2QLFVV
u5dvkgRYdct28cv7c/ey0M4F3Zgmx6Rz/Sn8ouvPYEMMHmlMU/sK8m6nzkA+
bkm0M4XijZlYms8F3i7gzLfGlWk+ctqIfS55x2F5lhyeVBcTNWHjZGyj5eiv
vKdDlWBdKwI9l897xzRcFAH5OwkRfSbJLbgixL2dqBipcYkFaiZxpYM1BHyQ
wQFBqGWMnNNP5KO+qRcGKacQuSBPycWe00Plaz8RxTkv0uXtL0aTiK4ST2Y9
3v0C436ZogWFd6o9emfbqYTALXOsAyaJukB22XBrQnK2p4WVZUa0FXBiG+JI
pSDaU0RcA7tlSN+FFEfy8uYuLUnBb4Zh5o8utYV+UefjyDzfZU3s1dc+cCaT
s9M9EKtVKCORatEmJtFxIQDwD5XYv4LNLRhEm7wdOwajnDntBhRkK0zDeIcQ
zb8g+Wu+pSavB4NWgHVRep6RYBVI0ZbGJ13t8nNVZYfaNpqP9eduvjV9gj7n
69sgsnKB7gR2nvqlnRyVO/UCrxOdXNsym89CQ/CIx8XT55hEmU1phmUvKO3q
hVpR3ntRAxXZ3nr55NdD3/StuGYrfZc3t/RM8KwLlvl4+6JX7jG3N0yT0TEN
Xk/oCJYjitr/+qj+Q4tfkJY5Bde3WzT9bGe0CX2Y17oAsUDV6ZW+bA+Nbw3H
usH/mURLHMVUmyGAcJjgedkDQgc95u057WfpaZIIVaYcTrXipjKmHZEyuzOe
svDDoPNMiW8Y6aGmGOaC9kNulNPZmyO6UocunaZmUSFf9K4vx1Kd9kLjg0Ei
II5O/KUgLK/m/BdJrTGhkeEyBKyoxk4+ZBsEeY4W5ztoliikTEqO/dS90O0o
3P7qNuE1raPbke43ctlGqxAgBaUt9boEkmKX++vD55Fc3EeKi+di/EAYuOr9
8UbOvBZAkXub5U+Eqe9BXMi0ZChncusLBhfo0DOjpRNt+ZJ2tKwDff7L6wBz
hmUd0F0Y3FNhHuGsdsLjh1NdHWhdJpKQWF3Z2jWpyrdPJT5TWnkP0YBm5aZT
y0jSvfdmA2AVdZ6GvRnQbIN6z8TiWFHc+YoDJQi8MTSVlWummQMTjm2+T185
fQunJot8z0VPJAUQC30cuR3HLT/2Acl3irdBcV3cg8HrK2ssihXCKjEOhwVm
FSEwkmgi3mpU0oOFlQO3GLXyatXJYIGOW4XpAPVfErBhLkQy9LknAYpPPWc0
q8jl3kqMzjv+NZ4df+lNUVV0vljUiqOpiFNMJwtemOv7EsVa8FCdWRyYGVLe
8e9AjhmVrUx6noRp6/vmFAuFmyBwfq/FHxsOACpu/WXiTIJE/K7dEfzCrMVc
seDHdIFMamva11MCmgew84xYLKzn041hNhaqkdZDL1bAkImqQ8kh95ZIw7fl
AFZkFdp3oFTKpurQRgQahyg1aCtAFcyIwwrnHjEqd197yMpgx/ji4bgwZrX0
CWsgWjR1YdG32atbdpp0sHPdXxivqeao9JDE7HUWTnKlNBn00yp+mtbLtGRe
lAqjfeMCGQx9boAXPQJTxQegXxo6Je1gdfxctexb8wo3e1rTlkne0yN3hUnR
roBs8bAcar9YHZVF6uhWYiLyOepE7OTWyU0zreOTD6KWlJ99HXQnUToLP+mM
MHG/yWudVhbX2jp4Z/qQVIsRIyuPltojicnwrOSCuqBtEZLpF/eJCQqfPhgC
4N5eRb5KMSKb1E2jeGBtAfmg+slLyrm0scbOcf7SBJ5D6v7au6SsSaB0tV0e
5XckrZWp+zrmbMX+drVvgbXWQlyLYyDbE1fY09xM9KWIv9tsMsRSTagDfxBO
y40bxGqMXj6YZbNGx2//A04U+absXODRfGATQQCqJTnvYjmIZ5fbVNLTIU2g
nYDYOv+NQPie71+QoWqsRLGGrExOGhM1m3Rloj9WEbmusmkyKdHF5jIpSNpb
QEgvIFK88TiApklHwrYOR2xMAzXv2i8180/j6UpAfeftxty/fKsYm143FHyi
5X5NzCkUPjCbVOUtgmeFoEPQG/8tC/tJAbvtty1rQV/JO765Gv3nTf1dV3nO
bfMDSAjgFi0K8rZoEd4G2bweo3FjfcP51YhxblNz0pzPSuhe3QOCpOriFXtd
OnA1XQkBb2c9Ft0T0JA58N2Nay4/blbcToT5/iBNj3nZEpzTxg0BvnaanV7f
0eZB3B2Cd0yhSLnP9mtV+V2jY72cYDMJzmL4jaotEb6DpHBECKh4srGzskG3
TzrhWQDaQsuTgQI+SkAzdrPXTZrNgmClilDTYyMBh/DqVdr/Mt2AzsN1WBa9
7QVW5Fu+ZWZvXPKmcxqo/WHm8xliV0LIbMvof4gIi4SyUu88eFyew+L1z0A8
KOb1XR4TlJoLmEdU4wTmJnE7KXPrIYk173eI2YLDCVb1D9lOUcTx5V7N5TdD
44LLkqTtQlr6AxTaQ1DTzcm66Wff9RsiwH6LO/pBJDJF4xz+UypVHv0ZQlXA
InzlvwUDsHNIZh3gofKQ/vW3Jpz9sfDgsRd374p3Mvx5xIPTau+ubVThlUZo
65HzeKFBP1jo8TrBZU4C4+5wNPlhSt7nU8U9y6Oe6CUn1rAoJq8BtfWd+I19
w+s92rasS4ueMoIFwOy0iR75T/kakBXyB1yvo9w2ktAuO4uJpah5p8gF7nl2
TPoONs1TmOq2H8HjZUFr6uqJJtTAgYCBjjIRho7vpomsLRz/eENXOsMOLAMs
wrS5E2SzMMsm1hSR78m+oJ+Vgjsw8lIejH/xo2c9VhpBQbYyduGooWRspYxs
Oudf3q3e68SyVtg9ShEhJR+yE53MMeZNk9V57e/eirEgYe0ALzs+u4vwcy4g
+8snHAc29ks9cVoQfkaThWv9s7uhuYKaEIfpelS+RHIbnAuURdj4ANSyJsUa
WP6SeAeKB6qqyg6mUFiEnemQsR+7vra3x/99tEgaU7xb/1VseqbbXkuagBsI
XKjmGI01PgmvdHcpiXaj3IPTfdFSFe7OqXfXdrKYgApbVcKdmLjgdOQWdn8W
sI21GKlTZUio93e6MX6EjTxKiYId6tWR4ObZSWTfF9nQNGFsJzk0VOlujwQG
5xdKfdzlqgXdURYMS3cGLIA8ryaoY6EJsnwRgT4z1os8j+iKrQ22UL2FLTdc
Gwm676bRvpEupyriLNhEo1bn3WF/t54jy5oDFdl6MzZnIHUyeuc2CngK9lqv
wVTPTfLyjf0KDlmh3+5SVCry+BojigNQIr5qQ3fAt5xcK05X20OoMA7G4KT5
jFGXLVVzeAX5CMuKmaj8ZwV+AHJqmoxmaPf9EFuJJVCaB7gfLH5egdeTOKBE
tC5W9RrF2mhQhmZkoxMR2YcJKWrN+zXo9xhiB+Xqje8NSVabKX5R4RWmMJGX
/ITK+foIUokEC6eCDdVdY2ANwpyjuaYT0Tf+nN3Wneu2Y7FBioW1wihewAXO
2Pp6ofXUNbfqupKrX8JV47jjLUWMbrTJdOvtXj9psNZPKCxfvUR3E5l6AQwW
oF8aaWH5o33psyC+PS4HBMkXkeH917NNLmdcnykAwIX1XRzEXr+U/0FcMgqA
7DNjgPXDb/44Mz+izOruu5TV7LLZBMZc25lAXtky/7nsITiGpOruZtmVm1FY
eU5zJTzlyr06NeFH6Fq1ATSVSTF98ZwMaSwacIKhBuW+o6j7ytm/wzQ8j7Qz
k3BrNhcytryi6N/0Fu+4gAw9r0APzlOvQbw8ykLJNOzAxcAI9P9YoC7ym2Nx
UOukiyN2BE0i03cgrC9P5BkJ7YQI4AuQWPvyBFu7QTgsoYWcWH/xzLXXsr4g
Uk/kiUc+keuic1iaLRPkE5lMzehArPrTJ1Vrs/nQwGuACY50sfufX+3GIiCw
7YJG9USbjgDBJ4NIt8ZOPVaeGNthynfp2GRYD0R9RdrpP4dUxISN963WB+A8
CE12F+7PjTvqMQIXTVORCJUPHLFFrOBgr0BcApHePoG1EUQQgPsFittxKTiF
UkLQX4d6H+q++tD+/75Li6CYLzmnoP4EguZ04rSnl42uTUvojJLowh+1TdBZ
m181pLSpEAah2Xh2gu+weREpek1Z56OeOxRYvP4m3R1m4sycAPC7ccl/qqyq
GstQYTSl8FsUzizDx6HlBqSob8sQ20Xn1dBztSgLJf9N6o1wVnoRx1fLM+h9
4Ri4pzdKJ8g3kor+36Rju+nvGxX+Pug2hXH9CwyVIbmEDziM0bxZEhocybCb
wbEV7/7/KNyvaSFCXg664UKP1nqBcrDPtbqau7LXMduUMKffZZOJ3p/WuHdN
/J53eUxRHJBWDww3Caf4s3x7ZxhCGp3vODPrciewGPCPv+ma+SVJSFR2GZiv
EJyKp7t8UyiFBxK6iYvsw/F2KXbwlEoSm7dKszdmbblnybySGWOhbYBMoZoo
Uz118xqkQoCcb2PJaUwSQFPMRQXEa3ZuWR4DM2KGa6TTxIa4Ggkey07uxTTX
YGgw2YgP9m7Yyfa+0TluPY7rWo75xCPOJi2zODpLQjBU5a4H8t8YCF6Do8ue
eqdv0zGfW+UE19wXj1WIU+xv8JCcTfs49/2P9cFIcgjSe53LDVfgGu0VOfIR
rEZ/0Swq+uWC9LaIxr6cUZ/WttjUfOU5C3JmNCjcfiYu9g8abZ9zOfbYSWHE
uvssH1Rn8Cm/UACfvn7v/7jPy1fDhHRBhmb1otvRZeN+YHXo4k7m0/dQno3L
94e5NErwzwxA3Q02TSteaVw1IYZpa7+WKYXngl4Cv7mI8alinLpRKEbT14Y0
JninRfzpzIZ8T0NNNSv1tBMEBjKECJDeJhiuzfYHuXcJh5QsgVIKpdw4Vfc3
ZONf7oK1oODMaPa6/6ToeOpBiRRtBq44Mg7EN3Ykfw3DE3ou/b/puQOZCwAF
0S93TgemCwcTZ7PYi+I/t1cKJ+t29q64WIpy2Kl1BNJdEoudYbujtvQxLTQU
auGLaiYBVayyQezcc7iyXp82bGhAJcrXty8VI9u+1nyE9Xj1Ct/VCs7sfIM8
p6ZcXnRncnaLGPkYix898dtPdqAlMZ/0GBFoLmgqXRLwIOT4dSpvNog7eAmC
17mVxnFwEK8+KG8e6hfxxQaPEV+R8CypA324Uepsq9YlV8jNvUOFswFJ2TfA
Iee0OiaIm+O85uVl4Qs6euBHlStujhvMNO7+4z3L/UQRoMXX5gp48Clzm3x9
zDew+b3l2fuCNg26BjAIh/ZvdFtCj0L9NV67Anh2hgprWJmDKwSzLkZeo74n
74Tqa5fpGf6NQGRMy8n4HEx7tvmtnq0c1FHwdV6a6jI/0Bj8ShPM7dX6VZlj
LFWqyrQgEfL2bQ005LzNvWp6y289jNu3iI3iqjM1LbX1q+X50qcLIrHZCN9K
BoPbRId2QEM6GIcoCLSwwbdZR6HO5rCLAhHq5NLsiOJRXTPsr8UtGAAcwl7U
QKZN+4ITkKHbHTiclHvlulY4iJDDypj3dTd+tdR3bNEL4kmk9rQKpYVHYbUY
NqmdO/ylickbJ3nDrNI+zXkX2hQIbsk902sSin0KiYf9LsEL5+TMfydmchlv
Sk41Q8sFBtx4yXP9e8V5w1t8v512vR/ylUZ7c0uh3Ia8xdEXElPqghlkk6ts
JZt43998NpKCj1k2U6JmY/8bGckTPP/3W/u5KZHJ6cLxzQ1ILrd4IboPj8Yp
Y1RxkhCc0H1LTFfzGaOifU3v+F9gkku0pLAOdc2tdwFg0kxEkNJQ2ORMjIGs
l/RbLDmqsjm8/q8Bu7sbJKd/ulcsv9MZrP0BhBP7oWA1aNPRku5Vha0ustpI
HBGCYXsFh0pTQM3O6yoTKXbxNFJm4EY+z4aiWBaTZ4EY/WUuo/ubGUpJryZ8
PXuhQtHigqRVrCu+kJc9m3lp8msqthz/RhcJXO4TzhqZ2kptXIyBC7ltG+oK
MA1EHpGVeIC4s2l+iF5tdPOY6h+wHGKKVAPcEHFhXb09uUtAAlcNVrIgBW+M
cs0MTs1N+/E2R1Du9GAPBzQ2BQYEoEvNZFwaQVTGB73EFvAVwovOKMF90AQH
v8Wp5aE7MrBJFuQjOSN8esjtAoS7d0j1FgzkqFx+HKm5YJW8dYCip1FEsC5r
WjCOkV80Tor+pdWYZZKaPGI/EmcqV0/qel5/0KRRBP6I+5y25G/yoSW6CzBO
VcaaIlXwRxZR+Qyr2J0/zikiBeSyvv0dMPJlfUJQ0MXll+XcukvQLj+9fjQS
IkeLBdO41eFjrS4niWt3a2Vri3dEiWwvsrgFsa+gVmcUhWjeBXan58G0moPw
AEf7i3QLgu9g9l/lqfe0YsouFiIJ/p66nP8qnpFGrID9YxiXV7KsYGHBuhTQ
NeO0JTk0oFWEcDl1WfzlOeZ3cs3l0CfpSmh4LG5blmy9Yty13w/m0JkMExmM
mGMQ5yVbCR3tpneW8URihBIs0LG7gwpH9KopUpvEzE75M7U0JxPFcQH5V7Sb
O4EL7BAgrdWWu/c/N5YJ1USxtfks/Jqrh+OdH2SFNoz4UovNfaV+aIGGprcH
rXbW4ceTeXC2PdeL1JF4uYf+vR2aClNZHaghS8xuYmQraUnzEAOCPzDMSe3g
uJmYOpMgmyAcqr6SlMD8jeB5vxWc/vZQ86FFNc2OfsLXvFam7JmOYGKialRN
7p/F8hdALYWHN5DeaGBTlEIpNJLkCd/HBWWTh5BaE+5/5K6Y1wyHdeZ+qemm
h1LaSL11iYNksLRhGFD6wcd+LCLH7ypLoHV2vo21G6EPlWM2EvMOPGemqJ0J
De/587x9CImKLlVI0gCVidanvcPhEWHmAl/vP/egSxMjomzVVSZMXd5rDZsw
ToCI/A7caQUcnXdrZhssCu4bQCdgYhhuukqruu7TTz2tKujOpww7VutfMmqV
h0EP1P48w+cUB/8CsWSo0eD4xPnJ11fWqn/tndXXBFF8AxESLwSgs8ziDyzC
IuBJmK1Qxf7LY4UixG7Loqg5DxfiTNRGfeOw9tzgq8aObG5HmzI56uuFUoXM
eqBc7YIWg6VvKIQIBV1NFCxaL9FCOmKDU15Hom4tPbXpgLZ2dSNmv1LEWjTS
6m0/wqvD4een21gmFc+Wmnfc32CJFxqzNkrdcLPjC8y26EHTygMC2bAHMIVX
YEUCEYTB/YQc1GSN38aQ/8JhjiRx3yJoe00nWguTs4jwW7TxwmXJjnwKXpkS
f8jyc9uI/4gr7e00rj5YfdwbWJ6cPcgZtVTxGrAXskcAduQuSnYTEIyuiQXH
c+MEDtKwcfADh69eAdYkg7rHm0RrBwZa31ompOrEI+P/WhOkJt8vmUnSFGim
/yqx2x3bdEVsYjOcTDzyqNz90rfzimdH3zX2296v5aonBoo+sCPnvhJNc8sN
BhKGd3bEhJPEjMZNGCbDspXoZVZANshHIKaK+4GGss/6dzqFfaekF7dxhUZV
lQ9Qclgkv29b+f2m32VsIMn8yotKcrUKtZIg36dQJTyuDz4hQ6PwaN9nHXRQ
wdMadCZ2xoXn8kln8dAlLeqxV91Q5x/l95HD3sspu+TrVf62qif7EpnDaLo+
G+Puz/tFYsScsi1HIVrFcwXYIRWbFxztAwAR2lCUWc2wpedmaRjNMeIzF0Oa
2Ij7JDQWrlmnnvmWPPvwNRbegiX7LrB7+cpU1kirD1ZWB0sTga1Pp8r/MeVl
NF1gGXB4gEuJWZkn3A/p/ahjjQQhGIpvpYCAn2UwlRADTQRIhp1Zd07bKTv9
SC7x6oI1cYmjyUlurr7VKVBlJz/SrUc3nM4rSPt/F5UgRP/GMFnzwjryi+Ea
F5hGca60ieK0AaR2z4Vf8JO22Y27rh67SndnExLgPNx48xWnnbqLVMEYa8AY
QwAj2u9CEwKelXsDfTLklbmZr1PMhapqHqncXIaGCo5wmUupr1Lv/R6fK/z7
r8wz1cqzeiJTxy1v24ghWQPACWdnnLB7DKAM278tfHWTWp9E+1ktXIvo76qd
fEdzdSh9GDR8DpLm2JqGzKyRVne2FOgtUJadPJxXFwoSwGVpfhZtRfBTZUMT
Ih+mplfr1nRQduReL488KhhZXeE4r3mfXe2gakbwjojkjgup7C1ZbNMwQRwg
XxXFR5cagY3zKipXoDOBbSCpIiNodwGJVWtNzEe0V669qiq7gZVqzj+kyfuh
8wd/SsrNGWgZJoPkjhRugp9XzStgCSV5Lhtidtx4Wbq3Wgzd3XTsa+iwVhOM
YNMm47bFdEJRflTSDVv8RH38JAg7Qbf1GSurZmPnTS41s9su6M3G6d9nfD++
KDuwslGw3EmsZdS9jJJMgH9ANzSdeTxdFcEzPCT/2L0P7PaUkRL7VXx8WqBO
7pHOOnKBndIabYiOafnnydww4piuN8djIMoutRfDItC/RqCBOyi98N6qCrE5
57p9BR33WipJ3dsjL66lpB97OxcP4/wBs7w8MN1NQAYubQp9mIGS45xtcJf4
9Jtf8uBctG1JRUepEHP94M6ADFJhTOCJ7MBgICxEkrwpOsgTFQrbw1FsNBc3
eTY+m+CZ0SGJ143JxNIC/6NY3eAcoFPVYvI4StLDAkLj6C5K3Ji7lvx4Zt0M
Suv/3JGCt0t111oSwT/NCNs8q602FMbrpnQyVoHiiZQJcZUILEjd+4SmGlLc
HYJnfPcgBQuI+XXZui92reXxlas+ccN5suTJHVncL5TSRvMKgVwlgwUkxoDp
VtlELBBwCxwrOT04HAs/QNZq3ZyoCgOcu1okEGh49OfsyJ/9AVobMb4rS5wI
4Q4qpoqJ5Dk7Lpk/daxsChrxIgkKjoDRhon8I7OyukmOO9jH5MvVjJKgBQr5
ZfyLJE8r6rCmmRJMsa/FgD7Lvz5emaqT1/6mRDlM+bL6cCr08FiZbeJRy1JI
DvwWgTk4eIY0xwtcsnIu4ZNfCFNprT1uOEciy6vhmbxXqkCvcUVffHEhFcMK
WxueR+nc6Xz1lwfvTh8PXJGE0uFAgot49PVNMO2nZDwDjaZyEIFHz6Ffb3Xq
NJXLMBTTYv23vJJRWff15uxvXWZFgVyG3XCqU7eHYteEGdie8FJZC43bkdVa
sJcm8JhjwrhEgFwNVYZsJQXl20raxxMOJQha0K0QZ2oKRoPF3lZHvNW/P846
77SLbVBM2aSzMJtvxHn2oKdtUeeDifrqKNtYfvuEg1f9OtXs6FKtOd+mZJQv
nOjPJHphtlFt7lVsniEzuTmnM14i8QwCS6/4NnBJA1LPUYSXjSYYVec+NH/F
K+3j/l62Wyda93MzqbmZoVg2xJ9ISMa28CnGtjIQp7pJOSNe6zybnWWfgA9m
nZm0wfY4wtMSUgsqq330DthiL5+Q/9aPJDT7f3bjh3CZ6Ggm8R7l9pYHh+UF
RRyO/Vx+XX3yH89zt/aNbSf+LVc8EIywnCLclDHe+zHpmNLoJQWVQIuszZxA
WwulklTtPvTj5J4NlM7yRVEOe0lgvbitPlLCHiOTUomHLmATPB2/iLHn5Xdb
oxBlNTnz0x/Ul5yNHREbhBb9+qYcxyv0P6TtqDVSLlMuUfc2Q/2WOtTBJMYb
okpdk0gvvEjCmJOllFzxn9NSA7+qRbwIhH7z4qgoFnyS3sPxTAfu4qfwYmoG
fCApAV75N7omW6kf/W2avGDC2M4f+yhxG6r/DliWh1Qa1q9+PKudYDUmZ/MR
M/B/tTdBJ2eYSnxaumSMJOffYo8t4D17w5cAoEbyTkATk6iLQvyId69htT3b
1RvOH08U3GptE2I0TS1zO8pcTgr9FjgrEu6gsxM5AJjjVCngC+fIcZ7GEGY8
+gjbqGfdVj7vOsV67pv7eRKDMbZ6UK2viJ35+l95MRIjZ+zRUjiUugPVYzos
Cgq0Qk2kYfzrXoidVpSIMw2lt9emgRrgQh9K5e9cWKD1llqGSDBXikSjG4ab
M/UBXPCipovYzVdUzGTrfC5qNmReh2IvHJemgC2pFGe4mD9EAo1tyEnUxK4s
nljGhQMJPJlJhauiW6lzdkfPGudSYV2qWLonpKsZk/aHqj5FEmZHyMkL70A9
kBpL1tu69n2FE/nDqFOPuKoXrpDyOmtRQxfecaoAroyQ9vWzRQJR16raElcD
K8WD/5YiPuZRVkUNbK4bOnvBDK75EZDxhmgP6rqwXGiTPPuMz0smRvoLIXbO
6w/y8rvd/RFSUQVoZbIFwNUz7didm5RN4iIo1FZjTEW7HHXRWkJnMlhbhuob
R3b+dHizYlrzNccdcTFqXDmMUpiR1kmDeDdLbKjywXbmCxhzTGiwmSxo2M3u
uW6X1IO+bv9TH8Z6cSp26PbV5vgIgrYA0NTWlruvHF3tVojtfXoSCuWru1Q2
jyD5346qCw7F35+FzofHIhkqCg2/la80ZN96hkX/gE/6vO1X9n70siAzEyGS
/NDbrggITYoMVZMDbNWNGe7zbXFvPYOxIwjxDUGDaWPGI70qLbvKEm0FDYyR
H+1pqfY65kvdcCaNaTFnNjI8k84Qq24OfQ4o4ucPjxhChgjmqFBRZUCZIQEm
c/qyX5R9yfnstEmHLARFI2DN25edcYTYMaCn6zGpvQQBZlZhwCjiKsz5W1wu
P7SBpW8uL2SfeCYAWzdChSBbnBkZ8wIZElyACPqXVDJ74qI+hBq+Qm/kmBP6
s+HswaV1d/6WH/B6q6NvXNG89WRAzhzo/sV9Myw6nPfbnJ+hwiw+vhhhr3OA
g/5WEoGxi50gQda0RSzGfq9vBmBx/fxpyjXJccJSGU+vEx7t9YITe7378vgb
P/m6CGOHkj7sOYf46DcU3qgvja3deYgKCsHVKDr8XNw0M1BgmWYga6EQHEt0
7TKooXREk3VIbV6W273vv/G1WAdt8o5+voqOPTwFh+YmDegcL61LMHbshFtH
Oq3Xn+z4HtgJqBURc2WUnvar14Thrllm3guO6NdTaWUazlo2ecgAfwrj7MQX
1W3z4LjWSm1iJfXVoiiBYxQaZM5eQTqyywK8qgl6nMFv4Erd8Q3irkwNlc2/
jVL2QRUuw+3OmBMtW+MPO9zwOGBmfMtk9PRtw18Kpfq2cE5GyvsTRsvgiT/v
/3v3eCTpNIJc3TRS40TqW6VASHOq2O3ivo1EkescjItZf6w4Pf5VAfjhhLB6
GfdGHmZB7GHmzzhqs3DLd9yNu2MMeYReLDxYTfrcgTsQ5JNrK4eGwlmo6YGG
M37owWIB/W/aJxYhNYcFjN9YZm2ca+y/obg3b9nctNVv6TX2PcHQxE9yXyG2
0FwQaHpeIhDoqibdxGnLYIOgeZrY6D0Gbya/N06/t7l/mjZHSFwsPFnaQ5zQ
fY/mRp6g6KNUmIy/eMxeqHifYcSNQ3lP9OpbRpjci2vtZn/cU1xG0PGiF6WX
7GV4uMH/mxfuyFevvGn/qigX8kJADu6NfqDPjvzPEr2LrNzkWYY8VdHM51AE
P0Dc+WWUoJk1TVAAdFi+tSbiJpEDuKaWaozoKV4zXRTY9Rkv2FAs4tYQUnIn
1B/PKd68oVLgKjsNhhV/n2NXYignazFDWiHCyugeIydaERmOdI731iIpS8BZ
0IXC0WyAeP/c7HZ+VzxuEbq4CuP+vFBL51Ppd+2qfh3oUe30WoYVEJIVhnUx
ZaVIIRJ3D6QJ9v1PjC94M8zs42KDFZmAmGsYKxsN2x0uFtI/4McgztaOAmjc
NkgTl13qBU6hm8owweKPwAIMI6SGvWR3BUTiLWBRWE+9ucQQTN9dztBBqI8G
gxvge26dqfB2Iu7IFwWmGYe8rFBfxRYemMgLrwRNB4q2GFXTfMdG13E/fOwn
f/100JoeapPMtKgtuVngklh1wU6uP+6HYtUSRVezvzW4sJoLQc4iDEPEjSUZ
7wI7zvcpVPGpwtWHYuZtUfIkbTEibpc8wEvfCHH5lhj/Z3s7WVEEDWl3XZ4J
RIDqb/oR4FBe4BUGy4SSYjo9YiwaNMKepw4N48WtrFQROuoULBpyMoaTXq1Z
PLP7As4s6PVLzGbCJlpa9H7cD1x+LcZ+QZdHSw9KgbGobiK93cnf4yf4GWn9
n9Ux3GHT4AdsLi4ocpO9HYXj5g0pEoC7scu3gjBWzpeTY5fXOcADSf5BAv7I
61Iw9lsGeJrhUNqh57zaJagM/Fwfe9Djgx7AWR6TgvPcXTQyczwyUfgdiVO5
ZqO++9CoJJFLbAUS1j4RfeWQnCnyqxauHOeAM/olxuL5nH4tjbHvW7OsWVjw
RDMyk72Mc5dTNue8ulvFBgsUH1dX4RKbmvDFe3/Cw1A2RUNaRiMcWkA/QGtD
3zey/3H60Igl9yT0w9rQxN7V7hXlX+7AEyGFc9j9JKC8DQ9pwGitkx0rJYYz
ws4aJSC9m4YFQvWzJHnut8B85M3O9chHN00iYoYdRlXwNJ8Piy8fmdwvNRZx
jcmbUr5n4dSd+pNoGZU4bm4oj7S4JjyEqV32gha7NhasoDZCP/7vFkVxfrLL
JuEXmaKO1HfBnin1sUphM3Xmk9MjNgTZoYHRbxdQ+LpT9huLmSAuG/2WXgPL
IRnOMzUm7u2vpILTfAgLSQBVgggy0gJcY9aa8AY6bGrp45I7Mjkc+p9kfwzz
n0eTlpLPozqAuX3mZAGdxtS3wBerM4mBxuwoZI7PLOBlAeiZ/ZB6c0fBeL8z
z2H7oIJd3Rsa42eZL1A2YwEfRrv6ISkc7xKoqZK8cRd7bARv1D33fxUEbc5W
iJOtFmYaejurem8prMIzTsk81WFCtOB1pBgHMQRUNeBPgTd7/9BXKFoHE+Eu
1PohsSu9kRMlIldcuD9GqeNaeQYfBmVspenCV4kEOv0183VP7M/ldnSk6ZTP
9VWizxEhZTdYdeAJmhWfWRWKxrzme+Yh8jaImkq9XD5g8fXlFCuLVHuv8XOx
36pvTt793ZE+SVZTkB8ph+oJ9J5f6XeLxvm7egXpTWS6tZOubkUgzNGsJVDu
ZqfAzdGQG2uxCzPRWbEZU6NqgIc99JecdpVw89i69CHFmy8gYADLSqC5EWbr
MsawNpeX0EYcg94gteAMgJL8rLTGzkvkxXEWe3BGPIcogeQeEA3Yt4bzk4uY
XjII9YOiyjmpqUILz8YkFx0kv3Njgq9lpZjKxOb73QURHKNrroduDH4zGcBr
NxPDpR03XIr2rj+NjCUt3VSbRyXbPpNgJQbXtFG7Bi/gOvFC3P+RiJcDewaY
Pd0lNukJDFvp4N9bsZQ/q0tRRh0PY8fEWmLbrLSltGQsl5tc5bU4Xz+1Lxy/
VxcBB1LZZHbgrPxMsB2Cin7HP7EiA0IX/jlzm+dARueUvpAxBDS1JlO3XEIu
pb9+ztW2nzaQ7O67bqmibA1OdPTbugYP9M25jlmjPbmMyjtkHDfrgCdnqfy/
7cLspG5C0dXxFpr7d2NY+2T0wtCxCEbDVBXz4foqbjObNZxDA5eQ0NTjgtSw
ZiG/LBriAYjzW4ugiQVWh47DAwzyhomvNOgTsyjuEeC1N5WYZjOnju8HwL0S
Tk1VGb5waCCmPVyIssgdh7VJtJVWNUsYVfnFna4xo5qMQhvdk2VUxliYp3bD
MQR6eLyAHuIW8nXjlhAbgBbZ17Q1LXl4m4CRkMRQ4nv50Bk8SuAqGLyWrIyN
znMp+AhxauULs3d9v8YijTteU3v3rzZKwMHSixEn+jYI0dYPiTHDNWqDzYQE
kv0eYl+oqxTg0EVP3kjWz/Og7rmwd9gL8abJ2fxxyd3wZKy8HMa4oasXoCQG
8rw7Lt1JBn5N8sUaLEJGytjK11VFsVyJIEURRMkkQZlJn42WPYgHsGgEbE+z
Za5co9N+kWesQTDyrVYHUl91+w1cNJpnun0CAyInvDKZ9h96Ubd69xtDct3T
j6XBeWbzKxNXZGW7T0nV4uDp+ywDpfwatoe+uqt5v5Qjxbr777dn2JBYG2BF
QuGjlizBC8QKxFbnM4fJHcbTLys/4PWe2m+C1X2/arXZLSI8MiNwKkckeFGl
0lhKjH7Q97WVdHr5mLq3ZElN64JrGdArI+BXJQHofRCzqKz2Sj6irL4Nmbm+
EoefhATtcxnyktTnsyE2U/pNPoWrXNvhzh1596m1aK/ICK8CcgW/gwUihs1A
p7WvI6wFs3kYd9rq08iqrowlhIv9E37icqDOLUYqiBrINTsJ3RiPciGqEv73
tAxTIIt4s/ckMf236n58vwMDLPMHjuIRLu3+zs9glOtVfa1C5kpeV8ATU6OR
eWmHn9sCCnZ17pXKk2Vx/v/FC/uzh+6PaIRxIeU3iJ2MKsNwCGtIvpm/ZZoZ
jhYGFvUnL/Fg6Nn079WeKHRUfG2yLAGQJWdpminndCfVYBRo9Pkdyk8YrGll
nJgN+UqzC4W37ClUBEfutTyOH1GnRpVAjEIVrhI4GXK1lS3jgVNomcZDJcOw
XCnGUR/vEm/foVBrJfVmhbbhHegeUBRX/Rn+ntfz4ladOwI/XtnfJZD2/tlo
ogS310PZ4ovSz1R2u11WvH9gkrwF1sqth5FR1FEOELPPVufx6Ma0AFyNfS4i
2WQLKSwxqGE7Lx7H/9go9hw9jZ3YvqVfYDwkG21sIU3kINEHwleiqMpkrXqf
+nxrtPWxnqZoFgYnPfI3oLe3y3A+Hvv0VfO6HmB6+19S+K777yVyIYJr4J7m
4y0dYgCr+6r2RJ6IN9Hu1nZr+2mypkR0oYTIpw8RVjerVi0Ahf/mbBbB0ilV
c39huy9u38H4lKfjDScZP9Dyl0gAThqp/2bsKfDuqTUwCQ8av2p7e1REm0EO
a8NQczvrXWr6B5OEMy8FOq0FbpUaPrpDF3WunW5ChJjq4K9sF7PJl+gQ8cEP
WWiY1E7y49ipat2okNi7vcSIAN/+SvKjFMzkYd3wM3Lq1o0uWiVK6THso14d
73thna5VtdTMTBfsHUn3O6hwtDwvxHJOIaOuXuSPjv/OmofHBLV49Yw39nIz
UrmTktvhCQGzMYmHSukt2tr6+UQa02S0YuMvTqTd5xdYGB30X6mBlof7SlXb
yu85m7538N1B8JhZ8GdsRNIH5GJp1QrIAEI0llVzfaHtErVIit+N0NDPMhAa
mJhJC3GH4YUmpQsvjPRAulYDVAv7aJCcsv5VF/+HzOFRJHvav9sZUXpxbOUp
spTRbY8ukGRHfGUcDrVggXeM98WxjSauEx5KPSAtkGdLwnAQ7U5PTO/AS6EA
NZhCsYOeeXVguxX0wCtx5goZREna4I7jWHN1gz1qVOUQsbtQpgW/LjGAndGg
DJsHwQ9Kkzy2nbqiIskrktSQV3gNAoSUmRh+j5VD8jU4ELpBo0fUtOzFDHSZ
3DI0L/wl+LYsG9Jb5GR8ycCm2FPLROGxA2NMAfRfvuNKAdMCn70UGz9Eoy7f
q3ULVz2R2ju3/3npIasy2cKoR8932CGNQ3VUBj2WeL0BHWc8UtAzjLEVHg8B
y54E9yYn72J2dTyIOyuD1cRTPfmsKMqhDHmldGPzNn5IlJ/4TORN1rKSJrVa
q81HTICitd12XcGugKto7Hc6q9pZ0AbLgR4qKgUBjD6F/+/UqxsRhCPTHNyQ
AOqGrq1ix47noMxGneLLWCLGstraYfnkqRGipHdF6GA5mvuYuI8QMuZlp29H
qo9SEo6rDgLLYqIyAdm9ZmJUgCzxP1F7sN6Nqzg6YZNLezd2l/2t1f8nlDBb
VQ82eCkzxRUTq5m3BWrdvj80893RSPEPt5BNxHW2XgFFrcpDGS4igmYHbaJX
SJz5eAu1V+C/ZR6H/iUz1khXCdwhXsu+uOATGYWs1MLErFPsn5yEsTngPIYz
DetMDdM4N0ZGLKaVi5wNJEt/1Om0dVR3PB6403lGioQwlvkjqs83/WiDwxEV
NlkTJiCkJm09LCScW7Eq6bi1DEESodv4+P2Ua+QFZSyB1DScaobBCpotIdhX
ApSldFIykC2mmUR5uMwZTGUoF2fj+LZvUH3PF3x7L94A0H3AC/B7cN+/qiAz
KucPjKt0Ai/9HSMlAD0RTqsJeQmfU5KPt1bNhFVOiswoqYfRcv5ThAUMaaeT
o/aOBVXvF3sPSHXoBBhcnCIGbDDdHtvN/+8sLjHihwQhChbTM0Bt3IFUJDgO
15Tji1yn1AqOabUR4X9qkL3yCTifr7i7G0aIYUa29d6wA+XtE1LMrdW1s6Wu
ChAQZeg4k2alW9Y9IJRyd1S/1jrstksAu6iwNsMpSrB4PYZxghM3hx7jfg1K
1xckVtpATsAKb8UkXl/2f6nQerOqHaC9nbq+0G82vqsfZ8P8V8F1tEjzzi7l
QBafhl+Z6INg2w65jlWyMM4a5/DnYRJjjxjIUt/H6d1bS23W7WjaLXV7/AP8
Bp8eR0/QVUZdfTplF6A7DerYtLgZuNbnX9zeNl7u1bIlx4NcrWUE9HWTmSjf
JD7noQXDove+oP6uX4VLqjysFx7oztgUGAVIgr4junf1we+NN4NJnQwWq36E
clh6A7vbs89FbPvBI3MPwjz12y5v09cxwTtab1ltaArooRSUBG9+DtFHHxDq
b1tWGBMBrWlgxid2Obpj6IaCgvwuVf+6H+UEmu3WOQ1k9u+SvaryqFrc4KBH
WgQQ8FWZ1nN3PWam94BsPQqK2zUay422+oagQUzU86sMGaukQfcwP07e4UPV
wXRXruYdP500IurJL0r47lYzEA+PaL4APe6eIE0HfRthoNc8RkpmzT9nCDyU
OnYCwqcIylI7PyhMxO0ajzgP1uB+yuagcIIhmRwyT1tTHPGfN0UKevRBma+T
DXKOZ4Rbc3nZwydmF3Y1IA2sXsIXTjNXnVdAokUm3NM1tz/W/eCZkBwfSWck
nLYMDEFzbu6J++JZrqyrHGoyBQyOPyi82ARWWvhxcMGAGzOgvcn/A701e2jI
zil488B39hY6jBZ4cKUn4RRxR1A1h7IBhheLTbSrjeXhPGMXDDe231btDqDZ
9wyexwIq0LDQrxwZWWK+QDQGUpUk6x7UFpCZ6zJtVObBgOh7ya/gv0XWMo46
FWq97xTF7tU5JhZBaTe8++UJR//aHqnE0FvJbrIQScZHKHVCA1/BsXmRLkif
jhbahrczcjMYagXQC2t9EdbQ89PKq3l4hgzcVbrSek1TWDrU3tWjYOzvElyk
6wiVNVn1J75BnFtHiHQyqYfW84RxrnrMhXQcYJy7f1FGmgHMqyQTJfE9++FB
Oi/Oeerl7hq29RuCE8vSnK6bSEGhcglAAkjs0szgNTd2eSk+wEQ21d9wl4+s
C3ej6HRoejfTr0T7GBJzvToX6pSd6XyCMhgG/WGjwtC0m8i1EXdnDCvVZK1z
NF3eOvDRVKOtiKydy5SfgLLaJyerTZI8btD00InNbmvqYfgBfu7e2ztBEq7d
Ky4c2DN26hr829r+IqcoGjwhfxrUGSZhGWjih0vAIqlQVO9Z4u52LRWi2iwi
W7oQiw5mIgkb1eC/rroyjGh2AKxkrVh6ODjdGsJLbVpcE6n3K4q+t8E3wwcr
7fr6W/Kd3rhak9jr4uHXDRklHqzi8cqBYtjrtYy03ygb42QRS2QHDSkgcqQ3
7SGb2oeKTpH6+kle9z4R7OWCRWK4uW3LCbAglZjoUeBV9wf6djcGNPr97qba
OhLXX+VMEZjALIeFxp4srHDv24hYXQov/PxWX+El01r05MYcUfOiw5NSh1Nk
U6hNBrBFD08c/H7raTMx9GnfEF9c/IkxCfVEfiWclEPMwkclQPTJvGoPHcnO
s5AeON/Rrajy53qqy9Ar//kIMTvnD51yHGpsVUJcWHD982VgpKogmtlcvTEQ
2fNG2Nj5VhQjgTMaEY9539IJEL3etpNMSEumqqpX6LGCT2HoMraY9m1BLfhz
zV9mjzIcGVam1I78ZRQZXEPh5Q2NdYh/ylEjB9pI+uEJBpJ6mdA6YHY3hK8n
PG0ozZTviqTzOFfWfvQle+40Ac3aYrRqsTpjJNotu9JlWqUENLGTLHPIxuxJ
flQpLp+oF7NqEJoT/LjyYapATEVYrBBPRImpMW5930QoBCSDxu1oR7wxk4Kr
2f+ajFR9Hja9aUnE/dR27s3emPlQcAIdm7D2WICDwk/pAlpcHKATf4PG0SrD
UV/pkO5HvxRKHjBKjKaNOyUhCHxIEl0Ns3tKd0ew2xBxWgozlc9kT32E1Rca
IOQFMTehcBHMxSrCE3MLQMSRK+R6ujYSz5Vg3l+h2nf0Z5oKsPnoKIxZlP5r
aYwe3s9rmSuImetwOC7Qo3Q9HhYxr8I2eizI6Zb/Y27o/VhJ4Oz91Rvn5Bvn
jn/CprxS8AjdEyMDKDmz2KcFiINZo0XMsk1UTRLpQEcNciyXMMXQTJiyR9Ym
tVifuHu4WedURMVoD8Xy5Px+rcXJ6wFakBXfrLisK+6qHC3uMpu9VGtlLZk5
Jd7IvG0c2GQohk1gtyHVRb0m6rrroNXv9+LJzeBRFITd2E9/n53HKAOIxYyd
0yTG6VUNZsfQdC60Mr5RG09dLwY5ora9FD3RzlurcPdG3bzD8HMIBTkl4+Gg
1Iqhvqr5RSUtmIdLa1GlOyWQPdA1Si0CsaHsULal9hIRve1uKmtagZxqnmmo
Q2C7jmqgf1DAKFUwtkWT4b+GUPyDpD3YHhLbOXVBdVdJF5G2rZVzJsDvQOPu
FXs5CjZKCtdhFH7ZITPV48Og/8UNFT0dco2wDUHrulwTTBXylfr4OQHaO7Dn
C8U6+BP1/BF0QQCSR9E93MS37UFVXHcekcLhRZsC0CJvV6WOGg+M4ELdQfye
00Z3SoB3Srp66NLbpkvlUtxCrAbr+K6IBAXZgbwtZwz3hvWNxtuAuZDJNnMr
ciNfHT0pcgrEMopkmurjaxm2oG9qrVDVnHe8ZWfZLqWuXwpWvf/E0R4+zB3k
U41KUTxwahO9Qru6tww30ZkCfSPIBSdJ9QRzBaP1f95hnsRsSPZl7CaSm7lJ
dPQkMUMHXrvE+WWApCFVxEZ/2QvhwHfW7V86yq4tHmp44wiIgitQ7rF4oo4T
e9KlWoCt17PNwpuIJJDz0LX7wOyj5itZQg7XErytvhxzGf79iPVRPzOEr6XA
rpyNm61YyIxZE4ej5el6ALFDU2Ywj6iMfVki8Kt76g1SNuBa1jrVjIaYkbIf
P3Gub92QM7EESIe84ntrg2EfiW02bItokTWXQ9AenA6qMN46oXCzN/o0YLlJ
HfPTaKc8WZF34S1xMutDYfOOCqNWV4suC+gJ0kHoL2P3W/yfgxOcV4+J41GT
6vJ+eXUsSDIWjxAhK0OtYIGB+JqlG4XGk1/sSs7QEsdOL2c6KhhnNP5mvkg2
JLeXghsI/oAxtRX9EaZdipqJYRi/uMknRPojzvDMh8vv4YX8tmTJ4FhsbASe
YrcVSh5aRHHhv0cahKLofM4RuW5gdka/8h9aC46JMlS9cvKi+oLp2kO3ymWV
fVjYZY7zEdBWgd7e9+66Ltbhl4ZRn6NoRNMttiyO9hY+nzVOFlqUKCTcOGxp
OKR4vHzpUVGhuL8GvDbc7RGisTnvNRfIGNq+zafgdlHBszZI3Y8/RLHQvQzq
NCbUndwHxFl+Tl2yV0dqjYDQSHnErGwYrekyPf5meYESEAG2bBVeumw0TTSG
2Vt1edmWjTasMBlrbzdR51SIOBI1dD1dSECC/P4GCqq7Wl0SzTV6vvngrVXu
LaaMaU86I6kVXxL/98OjMgN+P9yA4iTx3DSzQYC0DPBQMrmD8hpGAe5QC0y2
w0rnxium4YLPmE/NodfoCUyS77nMaZhHm7wH5L6Yp1x2GGLEPn9/2MvAZDn9
HQ+MchnwxYyp60OYZDNNh76CiEaPiJRUDjke+r+QXT32+HFh+Lmpl7ighV9U
mw/hgLyJMzySXeTLRcyvLK3n8gKNnlsBznXhlFjm2bQwm2wuljcEJQ4xTf6E
EGV8C+hhkdyRWI5JbKAQoyps9YfQ3dM+nlueeAa4bt6LczvCJdDvHmsOghzj
TMmEvb+zHqnO88C2ryFSXABWLK1YQERT+/SI3a8aXlA/SuLEGIsKeIF9x+uH
E2TsD//XS7Yf3tjW2KKTB6xpQjMd/cPXg7IPGVg/oCezOWfriCwNEGd7kKRq
U0rHRG2aFePCcFULVGAuUhHOg9cmDic3r97Po1EHdIZf8DUk/sj5R6jwAAp/
Jn1HsH8EhBgBMupgng7r+pRyqDxxKKTcPc46mPkQb3NbA7BqCu3YG9ma3kx0
7vcGHecgrGPQ640apw14F2OPYESHVnNuUR54V6P5/isfRcIpHN0XJZSvrRen
vUx29KLwuxfuUz2SOQpVcpo4EWVRxZ7Uf5tHWx0tu/ojaB3LwWAx6bhZG7CP
WgP5In4UeBO/dq6hAp2Bjye01KE8xrtCYoGUYnpCqGuuFuehcNhmXTt/Wddz
9FAN78xBERUQAOefCHPK3612gSjgymkNzwz4rqNg9xPD4k6/Vy+t67JoByHb
a6Xd17U3umuHWbnFdvnVXYQZxgBySqprnbNsKcdF16mIZ9vyJ8vfEq8vYUVX
4i9ZLbbE/rb3U49vG9n2lVJaTOqHJwfb/y4tLBS+1kP6NxynZmfEGeAhvKQH
4Dnjnr0vdSwbyEOiDrGdD3jgX/eFyYF7pSSX9EHpJGG3iuKl/1gpBdOdXGq4
tm3rT6w/5jnQFi39Anbo6snjpoxOmTolbqG6iYttK3qKOJs7bmH84zpBmelL
mrLiiPDWWlkADgrdI9a4MEZfC23TONUsQmvUP717OvUcug1yJ243geR1qnob
8M3C/kRqdoFN3VbSvsf2LdsVf5peFKkgq52GrJND8MnbBE35NXvqrIQHS5YH
mlHM2esbxL0CCVYQnYwpTcMYLI9Uc4hB+HLBv8nMIObBLZNs2SlTePGczJ2V
u9V+rmUiEVyNAjVgdgRE278D0XQVnQHf2w+cxREhNPUDzdCcLfbhMmzo06Qa
lLPSGrWTahxhpCYkkrK17aJYyW44FqO0B0ib1WirKcIPDszJRf3kQRQPT1Bg
B6RIAk5hHIn8ahA6/HwmY7/Csj48sqFOOUPqSX+AW33JwSiO1ATVyhWrRb+0
eVtLOrcNNuvkjYwzMlrposKpZEd/S0SeJmgl3fFDvs/anvgnBSVHUXdIV7GC
+eRsdU/9bZF2dwJR5LgWOHDpOdl4C7CBCC/YSOYPPAgCPcQfNGjz0VcyqwX9
3BvoCTTNp2JwYKOtaiDF+jTOBOx4HpCsHWTsiI7eSp5rTSTC1hnQTk7c/WU2
RgyMicwnfyN5+kWiLx178fzlpxMs8kNq2VZ7SvF1kO0VQOJ/NT3h/IyP7+VS
aqcun/SNd/l4dsmvCn0aDBETMnB586atsK4PAITueGVrsyQVtw7NUb3hh4WA
VWBwGqVsT1nd4kLpGYUaey69CgyxDciNBoDVnsWJ0/R+3Qgm0GW2MGW/g1Q+
1dpNf6FmnDQT1KzkZiCmRhh3tb7j+JvcXa9Jgd8JCmW5MqOxyAjWZTpLAUN/
66yuf8Fj4i7ffOD/AOv1xDByBIbpBKCOV0IRI7pIXadp8WDEcPF2UtTKXblw
1gchUMjZW0Nvf3Mw9fEkusPXrPud6X1FBXflYZ3spEkIsoPFbcFIbf8dQMkY
dXgyClaZBj9TrvdW4dD3t2WwIaeiCCLgSx99EeUxRXQ3MXt+ZReIzFklF03R
oc+gE3ua1UAoTcrDljynaT57x9i/oBdMuTSlP59yklLj1rVXOxrX3q7CTN2U
FVD7td51faALH0RbJJj5SI3vjV4NRnMNU2a2Xk3jes4FQe4cnKLnQrmgWyrg
pU3f17Hg6YDmtJpKWr1Okjocwm6Bkt4tEsCS+yw1OOoLuFStD4XuRHvroCGt
h5eqoiR3A2yyEVWZEiNTC2oe2MvVUKgPckEKoakYfPHmoAj1rMwCKvG6h5GV
DJBHe8eeHZni9CrW/mSco+xnIO6rHHBADxf9Wnx7rcmRp6aSbOpFTr431xGP
9x5GD1YRPmzNZLkJs9jRWo4lLMRKb4GwYw6K1IctzVJCVKXx32gtj97wqcYG
dhf0DvBqByQ8yvo4ygDJWmjJaGTMGZIQXwJE/IyAlOnX0xPGO/2gfvanRRa0
zfNtgBzrEGuVny/nGGIVoUaBcG2yokYnefmUY0Lrpwm4Zh0AT9UB5+vgFo2y
sjEAdz1ErmGobEgMkb4xmfpg9bjiq1J0EJTQiYoyLVPjt8a4mX4eq68NAFcj
XxhvZboXXZ+XpQptbzZTIlK3ISQIP1ilg2apDmV671wsu8XXW+qWRsxtJ7UC
art4L1W2grXoZd9n45h8ePrnwL4Cl56YFO8r7MDyN3PSxQKdJm9gOxcxBIir
ewPNx2zat6AweqQkToTObsFy4ySKMrPOf/yGJxFUj9l9ZGIsBwDe1mAATtPZ
DFa8fDbicyAKbXBr+85g7/cYJ/rQe2TH8NcWZn43cR0gwrHJ1xpgVqiGLeZ8
s8JZ2yJiQnY/VcTUgnVHZfKksfj5SoUSRVeOng5YRbFE+8wPeR5iyvGoKyPp
dYA79hF6fusFjWLDeOMckooddBomjI2vgOxwuXP7IqsS2fvlgbHD5mKy5ZnJ
xwx1c9VzUKj9uDXMz3+Rg54UngkuQe/9WtdUQMsNaka+UcX4ozdGY5r3zxmb
SZG03i2li5kbjkWtJW5xJyOsdGAjnvwU/FkJatXwBqj6ULIQrdm6Z5iLnz8V
i/Dlxk5H6kZnbkgPwONwUl2WhUsizODDdRpDo+H5HVfqoysYD7RwJp32DH9c
NOrExBhNpHj083ZABAEuNzjUo8xJUI1mTKCg0Ma5r4vmUYHwWTKKO2dadEi0
vCTtEI3UXXT+xYv3oqyvJPqRLLbbUaow+uWJGk9LOij/025LED6j71EQrQON
JukLvBmFAp3vPOaBLpE9z1GrYcF2VQ6eiMZOg0W3fkQk6m3PrHWzKjXIdiNQ
ipQdqPPNaw0OOJVYJNo3od585AgC1o33RC+OPrDWO93WmKg2j7O2DVV6BPZS
U357s0FNsLLojuUj4s8IrcdTv/zS+UiT3yt+rbOXTan/ntjXy1aZ8/VnV/lo
11gKC788i0FOWydknfegsPMFFIfAFbflGZGq8PVUBKlRlAKzItI5WhFUj4bf
Kc4Q13TyB5gN0OLDFwSy0Qt0rhQHMIyc4ZzmXpuw1bmqqbDJKe42SR0CU9ej
zUyuHRpzEus0zAmUNH3xiYPL9bjRizU6JEgMyn07GD2v8ttmngBlPSdG/ehP
ZdCiYQT9F4Kh8shAh+ijAeeNPP/PtsIqSoLvWD+LMvA+A8CHZjnECePXEKip
UZV10XRKTD3kAF3ARUIVivwUzolqa7nwEeE+zhW3iRCKOA+lFlqVvrCsU7R4
LZfAEl35JxfgeQ9OV8gKl7v2cU2P7telbeeHbx8V8k+2UWbnbdy0CVWG5Rqt
Md9XQzoyljSq5eVVf4i0CVeXl5MXiLKvYaIW8sSx4NQzkhAeefU5h8oIhQMO
to5AiqOxvkQHHjOb3BGTvkYcp9xQo4/t3y5ZvESJmNAZGVN78BI/RQlq8hnp
nOXslCxQnTcSeRJT3Higf16IX4AET9t8Owa2p6dzjS8AZvZeQOyHMT6TYQOW
b4VxlnurQCwUAfFt27yYlqhIrI1E2EkVfJC6Ylp5YfzCjO1e2AHb/jGCyXVz
HOz2PUZu+g4b+4M08YuxhxJY8maot31yAcIBEqrik3Ht9z68Nys5oZpXBkNZ
6T+TVPEV9oMx8UePDunOI2i71N1vSMISxfRfZUG5uTZLzIuHR7DuPkMMiWFG
tR+t0kOvOCBPt8Jnqf/6Cpfb2PYv+zzmRSigxJbLuXBkp3aOajo7ceLOFxfW
I6Dl+wBoSLZqSnB0JIJHZIFTZjZ+WZRhFZfFgBQX5AyYkm0hgzZW9SWAj4We
OT0AC20XtfTX9e0q4o9drw+2Mza8SoUbaY7a29zK/8kkcwnBdUBwOoHPss3Y
g77ArsZ5WGn960Sce5bKVh1nyCK9s4qdgUdRXCWcdZs9qNcUxdQI4sCvjCyQ
brvCWfNfJnr932BdH3hg1p27krs7zOK3KzsHwBpOS7DUpCOajBVBQM10IX8i
SzNd5wEzliTscvumAWo07+d43rW0UHfazapjENAMYU7Jy4EFrbvo3EG2r1aS
pQxg4/WzdEkYoy79VPf3GD6mjuVTyb6MlOJpmo2bUK0Q/VqT4YOEzYcgc3Us
HkYZj3nJXUwyRIG0QRJB/2ilYdeTVMkF0iWQY6hNAPJy/2Bomgf9CsVMauUI
TDsRgYYyYLci7NamivYEYkToA8THarnTFcjz5lHROlt06mgEKSfBfY/zpVGj
Id0JvbRzP8PS/uPSaXDfYQ1gMsSkKivsZ7NW3M7h9s+3/XO9KelzlnrXhIEH
1TzDXYiTkBKQUFdtw9Nxei2GjSwHmHXDR+rWhj8ZW8rBz+e9c9xBx9m3l/6e
ryxU/o7UDQOJ8roLMUuQgnR97YwplG7y9vQdLI344BXSGpDdhDjOgO8TqjS+
IvAqOOQW/sTyM/A4NkEAQLdQ3z1wu+pTDUyHnEP/L+fqS59Q7T+4YLiZX/Vy
JHMzGNFWZ07gvjClSgOJtNijVZ5vZOWm5YFr5QIFRM9GT0GMdmQ1On+I7jnV
0H/X+dpneD4vLhDp9CBNT+3j7BFfVY7ndXGasj1UrxiYjFOro1VIC08aALVf
mP2XSjc5TLi2nV0quHWfskgwlAgNDjrPod6/v8yjfHqAfIy51zoDZikRh0Yy
hLjiYMpIkTOjnuSHCAjVWmeiPMT5/gGl1G4fP4RTHVfCT0YlGjy+XD95jbT7
9Jt1QacolKCt5tj3zIJAiz6WqvNbG6T68rmn5RiIaht/3agGs62DQxObpc8U
0fnqBy62jXbMH6EmFAdFPHA1d/ISaaxZS9ZRdc8341ae4QDSNKPKlUdhjaSw
TDzl1MhZgH7tQZdJw8oah+iMx3eYXbAxRrY1tJQD/4oBio2VyqslAgOmca6G
1ryD+BtbXfsQv0dT/PGTiSHP/rQjQ0hsbpMwEcgTcv5k2TYPI3FghIBuiEcn
q+GBri9IMABWKIscrwBl61RMJey8fi1oy9ueaONO9o6IpAANqEG6rNwP5F/Q
GZSiSjBT1UIeLHBN7WNKGA/LsSBNlttYfKkOETayss6svtrrN1Pw5jkG+Fb8
5VC0hOfPN+RtH4cxKYIoU9r28T0aSGMtGfMxcCizWOIVD8ecWsWhXa7d3mCi
Vb5x0Jg7C/9Us85pn01ZoioISS87Omn69ho5wDfYIqI9tAWSrtAQ48slPE+i
g2zXy9TUxtm7KlVMZGjZ2mKuIIu56+lEarpVRnCR6JGI5bwzwexIkErHzUoz
Yx33jZkkMpKVmah2IEOKdYRzysdNDP2Gqd45bX2tLYP6xUbqvEFu3sUMtgpW
AJGhhWNjfjbw1giawscjz5cnbaBVbHXNSTkKIZssDAer/SRGejYJjTgmCMBL
xwCfw66sCjPS9hEDR3tWnWUY5Qu3HrFq1rw9RKcbfimnfsdh8VylkZr5tqPB
qAtM2ZAZiQ5JsQdABNwY3zXUwmatB9H7UcCq6yK6+uIdF4RnUq7JELk0GCJe
aEuZAVBKQyHs+EiJSP3XDLBINSr32kErznIGgOk1Iq0Z4UIXezLTendd1c+Q
2nhBc1WJVdR1JzRaVB2FtLTjvXYUn7i5zs7otipzFwCJLQ20KVbJ5wbSoT9x
2ANy6Zvp5uuvmm++Gr73n2gSZ/LQA55964+t/+95pHKHT6KQSPYnR3S34X9+
6+ecOnrpKHHX5z24m/DSFzWAkmD/ywym0S/3nFr3TPUrziUwQV85t0p1ZzWC
7ow1Rqq/cTq37bHauvrTnfuTAi4z5q/X++J7pqJjMStioNGQ5B1Jnif3b7ek
NCaX0ZTFm+N8Ukzz+O7hxbEkNSVK2rGNVlBfroEzynyNXsfp8gResNU9kQPp
DxrpfUwYe7wxSe+B02gc16B54aA28Yz0k98o4GQKEFaBLN3/2+CcImUpznMH
DoAXKcNBlTGsi1iKtaRoJVldOPP+TWTnI0wrC4GD5Q8g5PLQ2Ywr3xYwn1XU
omUiK3B43qcSsh+NVwxnIltfzvNFjuLKCYbRtRkhPG5dpymdIvuRdazsCzAY
Hf7JP2nWjww5vg0KOOV6uS8oCsYqbWac8IzLUygwErea76CUG+Y/2jaxvO+P
OOuUMTPwAP39+baj0p3nq41NakU1Fw5ax9qmejPeD1zrrXisRHogqehWgPc6
3XCjnLbmkiUwrPqg1Ouj/oIwe0WPyDg7XYd2+TY+YU0wS1av5M28fDukOLs1
64RkPO3KxvHzeaBxFZSDuOKkabeGU9hY5oa4mPWFomSWj36o++fDPd1/aclM
m9H2Yvlh54p7pFmS5tRRS5J6EiZ3THssxW8WscJ60fDzsenTLNfGI68Lr6FT
rB4B74xJu9O4yAgBAOrUEBRVjRtQ5xIXN8q0q17G1OUMM2o/8oqAuI2i5xE2
K7c305u4GLd0j3r3SR4Me4GzylHm0RR4ql3OVbOQa8XQZK3wSO0fVGptTYdC
7Vu4TPRE5BJPizQU+ocJ+/cMYoWPcOSawppJoaLZFXJqQ1S9pEn4QyFUdMtJ
XQDM30vmiXr7yzodytXDWgy/Fjmd2MSs+ubcD/imwVMmHdmlqRquYBmjiHDZ
XdDI5IPXA6XDGiQD5NdJC8SWvZwUxKsTTBdGz8B9vTAaxpy3rRrNlDOOiyqq
sToCvT55+SoPaLFXiNU8gw2tGnWcIXLHVgGwUMh5Y4ldvod1SutF2mRBBgdL
2gANliRKbJUHInmjc4SQ/pahLEsaVmv2HaJiK7jfyv94cNbHvVdgE0gjArS2
e24k9+Vk4nM58jJHARBR1p8b1FyTD3DAnGqNNGzF/VTnKnrOsZHpe0vNuNQR
L8KYcCdBO8VvJLlyMCIFr+huy82QtCSa3Kv4nw5SglObYJLQIt3flbd/9XDN
EbgSEw8B0DnsOhf10svoYnCKxc1HS7Yg0PCipODgaf+cVgYKxYbLbXu3YRKq
PYy43jqBXOeleD640m2lEx0Y8A9UTzlqEeKQD850Ta6j0d1RHS9C1/9nCRRo
ry+Hp9i8JY20LutRlVxU39Zp4hGBu+2/kmqb4SQ0+zrosExkyiwqiyqLoaHd
h3WH52LdyKvAf1sRsT+JdSr9C4f9eMMkVv+K9S5wkmED44xDGc9XJrDjZqJd
TkEI3aLNkqOuFE3tHnLkvjXpmQXfFbcUlvj+NHTnYfWR2ntIcwMfs4o6VhxD
XKZKSjQ1uFkXA0OC7dI/S8+kBhQaeuoH5IveVJ4slnpwD7muIeLDVAvvUDAM
LQyeP3i8zvqpGFYw7RMOVr4hQQXoY+jxsYARPcAj2FcQFu7VvYkuerP8XAMq
jjJii/MYJNN4spFecMOcW1yarm9W+xbUD6R+Cp98tPg2na/qiWGAvQlPHvpp
ETOfzK6E0AolyBWOYtZAYMnOUHvOh98r4etcSlq01RQh6JHX7XdKeeTmS1mI
7GOBqqS6kV9GoXVbrOyHWnEJ7BMINYg6T+hG9+t3kaFLTs11CO4egUYCRgnH
pVgvOXhLNGK5CIpmiDCDECiNYVDoDKUk2u68NHDlBCZSh7KOGuHRMcCYeW1+
L/Kqv3HR8CZBjraD6KgA5Vqz29gKUvszobW4jY0QbSck3jtpQbSM1T/Do8A+
w34Bm/5IGodJkoiXWIJvaAz6qpHB4QYxJlFQsDDYaVPIkEc7R7aYJTI4eLFZ
ZjCVj6vXCGvfyqS9JIn09PRV4R/fHuvBK1Od0Z6ek/xhN2AMWdnchg5+8xFw
409BEj2ahiGXHCw3lsvhHu5HK6z33m5bccDdvy7YSgN3CUN3ynWu/io/1v55
c3aXtL2+b6oiNp0scrqWdMU7jfS27+nonVTFfBpI/xcV5h962hvmAb1t0GEP
UOXVRolM4TvhFB0Ypaeto2cGxOa2uL1RyOFZM04sqMe3xkAKWADoOKQG+z12
NgId63f0FsW9VbE4pfvcLqCLygyq3RDM5veUxPHxEk4Z7kbfnZP7fIZEnGyV
ESjLzQFL5FHteoKz41no8yjW7seLtSxK5VZwnHNKhlcROEaeM7MoaQouEBy4
6jrPjM1s30nnVcMccXDVZE/CRdRqK3SxuAtXfrx1oPfOI+NgHgYPohac3hMd
+GMuw+VeY8aroM/LuVjOH0MUAZg5W76sSjgQUSVl8FkF6pFyOMElCTGMXpYf
5O5OFdWCLRqGCVfPt2S4BMdbML8o8rqdLFENOfwQ11W/RNp/H5CYsp/5xdgA
juNMPHawvk9hNiWIO2m30Hg/Bjyr/EuBqtxIh7k81HKl64maBgAFcJ2iV+YS
K5E06R5NW+62nwbYXNh9Jgg5buMX+bqa0K8y6E4JtF2W6BI6kOQ4Hesnd0BH
TlCZujRpz+dQnG5FTAKP2BC3FfT93I4u/VjDLrAJRweyz2Gj6L5RLUbK4q3M
EmviGQu2PeSxVoZg+T+enYQ7jDP4W5KjDa1Iyl9ev5NlVdgYPOJGszFtP4X/
EsBzZ8+BlZkT+6LKrsrH7Obfwk7QotJsAQ5nj9c0XPprLHuMaisx21MgB1qd
93pyHQwuTQkvyPkSnXBz8mSONRP9StgO9fkOiZoHeFFiBwgXDsY1/xP1poTf
2mSO6PFZ+PG6I6uUsPhgtGkvne8kchYJE9e5VQLxDdgfqlrf8uMaUeu21+Iw
kfJYTPn/sTZ3sEuZtzOF+5NzKCVBTu3lcsZ1GozOgnbexxOrSyJ2PMvPHXfB
7z98XUDokqAtnSIFBfpfKlkhROm6qF9451SP6e2CoVKl1upbyqwDuRSr16PW
rG5/ooQ1ONc8QXOAqOLbBPVc2yYzypRury71PyopGeDErD4G5il7O6v6JEZa
RE8RePKpCJv7SmeVjaVy5spL54YrvaXOsQBIpj6y2iWBsjiWsVOq4GQPZKPH
Xcdyhn85JQXNkxpTJg8LN90qpr55cuwyZiaL/qZHN1OAChBunjtD6NcqF6J9
fPqmN5wNLrEPli6XgFwdaF60WUOoBWCl56igwmjgGMYQv/TLEsRl1nL2++9K
Z0o8npifvc2Mr/lkohpZgOup1cGV75tGd+mvPr7WsFxdDm5TTWG+e/ceIuFI
azo+tDVQDPuxUgXc4QyT4Lf7xKiqIWbOeUE2RyZ9TKU8oSR/wjbuF0YyhYV2
ldTH3q9vzwyeKuLr4iRyqJwfRaCyDswSSy4rxEozt0jnOQcgAdM3ccQYoIFB
68htM8OgIUboizUCMR6gei3ij7iTTedT0HY8IiQkhjlHFYU9YnhgQJBNZNkY
00tx3HyscX0ojnQSLq/acdrGUlmjepnfhBDKTJisSgOE77STaHYiTCJn5cSj
axu1PWZFNOpjEQHpODIydRI5AB0z+gHKvqt6IYqP8imWm4UBsOmM0DzaouB0
Kyj8RBhqC1AB4DiViBG5uYwxv6ogh6u8jQMkts5Q36TFvzuzXeTnussAXcj3
aULMDINvBmCAMJKIposEddm5eVYDyxc9hI0Gf/nJdKdTu6UrC3g6sH+GUSK3
YwOvHnVYPW7Ec0Luf5+HoEm6MiHqmOPrOdGpZLdwmkUsZEK1MH/p5P83KaUZ
Ux/N1cyGbKGBz1jo8q7dTL1q5ROft+OCErZskQAC2gIOkZDGd+EN8xYaoAQ+
UfUDNHYmF7qt5Sw0SkDURCv4oPbcWcLCS9MNjk/OM4TJBUF7e4M620vaMv6Y
RS3JKHQ0pwwhn25pTbipyx9xwW9aCoaYg4R0VsGaCNQwDJclDdl+3JL1r9uR
XET/oOkxj7lt2BRrYpWRnPcTfFkVRsq5SKmjrFN6iGXKO0DjWlOs5YbqPVIf
/oFR14JvEgpqeRScCre59Eds/LLs9Mc07NgEIzRuToh1D49rRIXvmb3cDG7Y
n7bWTRydKpzUctQe/fcw9jZobsiHjFDtGPSVtmo6H+BZEg8GueEFdoGXmTML
RwrRICYEqr44CfskZIWrFwHJqOnwXCQZZ9dNyMtxn4JvJKM9TwqDd/Bm5X+T
4LAbuwfNe3opway9VRXVY1ucGEfwKehmBjzN4UlcXB0O2yQjqVZIqzHpvLQ6
nUW32Zh54m5+Vkx4BTIpkHVFgR0IO5r8MhIojgFxdvsBfZqgwNpoOP6YhMHD
tFAHMxtJN7r1Vq0mboDE5aJF+5HspChcsN+pjnVBjV+kzZcSGWc12al2+MR/
lU9QrjT3BnKaJLAULDb+t0zPGXiWX1ABYXIllcrwAhSb0SzqSTTU1TAPbVUc
S6FdRVFQ1MzMcQ61donE6sjDgEWA2/2UkLkXD4U4ExT3pa8ZJe2j+cLCMS+d
QWRvqKh0r2CvPiHMDQgw4HzV9usMmQifqkrGWrhigW1Qv6FWofOb/y0cRgwt
6tE2zVhoKJATR+UoA41y7md4gpFRlQy7bqdnfqHC3sILOremm6ZFOhZOFiKD
JBGaKVR7xxHEjGc7uD1wUQ2qpiZzOAOX3bwrCUqsVhgoDf0K+rf90vO7Xb7j
SK7cW+LITvDyJ2tna8Z9z4HV9OABhFZECEFlQLdQaexwnBOqWC2EuKh1AbKb
Ii28D2zmYmjYz/COHXk9Mndjx0PevJbqY+sT4ABEihY3w/Nit/9tSQUqelK0
35ylqr4I/ZyyyDDomSs4ePIs4CT6i5H3JQ0Glzt+14ix3/IJXZkAbvLJNIUm
5CxTFxaNnpSFwyRJJLcZYFN8nzZ41uskGzV3puAtknm7yfvT+4ZbXNIi+KHC
hMAaBQbELtgcpfNQQ7UH6dEFtmvpNDegUbOpMmeGVIiNjcan4zuQasUkI+sd
ZGF8+WFBSE1+a04ptFQxrW+GHSMWMF/7yCO1M9vJ2ow16cX86E6jXV8RmTUP
5Vv+/qgROrdwNzgMTLu5nniyMMMk3+KSOgo7rsaEsjjWSGsSO8S+obi0lDMH
9cldY3DeF5huhQYRttTTEq44RO4Xb5CXhymxHLoKPbL8G83E2Pqtxw4zcAZJ
qoO7NdFiwmoyU/Dvv406t+db6nfM5sw08BNKiUvZDMoNIbh/WaMYenpLlR5t
ZbffmoAUqPJYbfLg0heyhXEa8ygNSp9xJSmjj7mbDkkFk/Q6J1tjobHE0kcw
Mzpy+3qycg7TuyZ5Hu25Ap4xkknwNiWLX8LPP4Ax2HjoA1fnCMrJGPwCvMW4
UxSsSE8AO2uTSvUvHEb6sqdkFK9YE60gUPODl6UWf78wTsHKuA/5s2bQyMiy
cvPuV9sZQsj+L3CiNLUZ2K4/vYbLeMQsbl9IeKoqtIsSNbUjkUhtqApzfILR
ARrOyusN2qoCa8p6XFB0kY23Bpja+1bjsd/JpX6rvgd/IIE5loKYBCmREdNL
9IPgCvtGsPW2YGvphmh8evTT79rwFEvEShdus1PXVCNSBae8rTQZusDfghNR
IX+dakc4QKWiR2ObpJwBLBSwimph69necRaPY6HmFakJ38Lc5Njb1vV61evu
gCAvrq8LHYw7YT/H+1JetGMfDXyCMekTp7qXftY/aqI52hM3Lb+Dm5P2xTXa
nyMY6QVJBUiNulcouksO4grM7dbEaiSh0ldNgmZJRXweD3m0A3U3WdEIu4Np
Cnm+CQGIW2C4dq7SLHEgMYLdVpVhpEA7a3LlQmJkEerX4bChuoX5B7mPR5VU
oeWMjrlkpRcDawvyDkt782NtYGoQreGid85L3ZumGi6PvCIAHDjblExESo28
U0w0L9j3Kf9uTbNkHBeszvDXfXukBzwH1dksa3W5jNUnxpMFIlj4TZdGES85
YHXs/FpYgPHH+QJUqoOidTE3E0+i39X+riRJbmepFTLL/m+qacJwIWnTGHtv
9VxPNhqMudX5gFENf3ikg6BZJHq/yfaKOT12kOdnJ7wZoTl6CCB74jI/ELps
N8tE65yMzSGBfOIYIkW7h2eVhcjIXpFF76lLiSTxtJ25kTbwLicl5723iLCW
Ut49BJlCMwb/jrveFHuTfN+IDGXAIqP+OzaJqchnR7ZYiBSszq3ltHOmS8RP
u68V8M2R75xzTQ+T4Ge9ex4X6bCVzucKDK8Beg1ZXRV7JVrEWMp/8UZspW7A
zxTl0Smv2fsHxEAqsPyD6DuykzzF1+RVKspIAqvlbSGIl5xMQUVO8cMUU7iQ
Jw1Jj+4J0c1Ym2nSLaNSXXou/myhuh2UzEBntKPfnZUfA8lJWxCpIAKvcn3Z
7KN8x6hB29UsYvRi5G+s0tcEDaF0JPi5Nn7d5G4QeYtBB5ncbT1nJ8P6E9Qn
EUejisfXQB/sC0Cuqg3Wxf139vyuiPcXefuVQNchJp+0p3RYgkI2D+N4vXoq
hr5buJW1zN69vmsfg1mkRhQSmcgPdFVYEoW03vpKeS5FxelF/lXeVsbuUSV/
ZIXdj0NBR9/eSQMTvptvBBWKt18/9Ue9x4Ma1UU5uQ8BJN16LEwtOXcWL+lf
mAWbiNmOFLy3DkrZwHDsjoHpLsPamy/lEW+XU6+o2haVKy1Vpu7EWvLt27jZ
oNUYqxHNYl8UGqDSrO1Q/uYDMamixbaz9PpKSdJ3s7G9c6VnzJAq91jyXnJf
P/DlWbtXFAWn6v0gPEcgNdHzyR1Xb3HTDZv8Cp1cQp+aTKqAHV62U0UvyaeS
ZR+QMO5QuvMxgVYpoFKFfCSElOrsKgRhtYPnnvymHCLm+6jBcKEh6Bb3UMG8
kqdFQIl2k9igRt/guynhBBRJBCcJWtn9AGMNK87vJylzsjVDAbZm3XSzYate
0FT2LU3NPClkOq6OJYPfnQ18YjKyr9FVAJPB7igv6V988sCY9ti+NJMeLtYx
7hOn6aUPtfvttAafUz1Qw08VAcf7SupLQxGiQ8PI7M9k4z/AQN+5toEyCu9G
MJEKUssGoQgRLROyG2t1ss0Y8tSiTR4+e7iBtHkmo7Aaoqa98fJYR1xTg62f
oBO87QokvfTQVsCmgO6W/PzyibL0o9LcqKNWE8xHF/VAL31qfJfgnUanoE1d
a5vI/aoBftb5x9U9jyj7xhBQlxiMRD/R7KjGP9yT0FayXVYHoT8SgrBLPLzf
5WfBjQE2ZbXdp/Lxe8E0urZECuHwVatjJtPVU6q4NJnVQNPbP4HKBboIELLo
tCQRp1Z+eQ7N2ngi8DB31voMwhxgIPEpQSET5Cx42w6aEgUszh/alUA2cXoZ
bGli47hge40cwaUwQ2vb5ZIElGorAd/SdCQOtk92U8QtMffv/LB/tJthUNs1
cRHZfuTMWeYbVH1OlVbw/XPqZ+LBLmPMgU7yKVfmpF2VJZNSrSFGGiF72/wZ
l6NXH7xbOWrDvKPJx1Sn5TJC+1hJLVljDCQOPjBwhldJvCYSrqT57mzwWkFl
D+fKP1Igsdjfz8uyRB4dIztpDviMQSP/MW0ZNLOXuhXBaSKCJWlXa6UhJycb
TJM9EUAXlPt6956uH9Zws3ffK2qyTRBAx+TkKLGFFMqqtTuzIIIImuiYDh7q
Rismj2gF2mJ82NxqElrVpkDj7we8wi8DO8P9oBGlIl6l8w8L0/pSoKBohy7P
f18QkDH8psSjBbTQyPLya6Y36pEW7YDxQWFblObGqbdapHEH1jql+TsRPBA2
HXCZoWAYWuYI5r/7UGI284mAHAkDBb9a/4Z7mGpMlM3wyXxtCYGMEK8XjhFw
3ED6DAGSOWPsgYq0UyqEmZFg3PSHccNeX2qEv9TG5RbDlQdHNwh4z8Pdy3S1
pKLissLSTq+T2SojgR0a+nJtPJDwnLXt5cHHhGO4rLU1hYqJHHuL+QPTGi57
Tl4ajnknFOga5DBGRnc9VbyJ/p++3ylpLzXJM6nRjWsTI6TtnfTmta/omFl+
zV0G3U03cGC41bq3abK9gzhjBH7G1LprbMQ2RhZQfqgSeCGDAX0uh1iGsWcJ
kNR1rcinZaDkKGj5nUwCvcImDE4ECVnLkxvgDxYULR71+ACotQRtJTx61Zi6
F7Ixj0+8/kl7oLBJsmE9bcCLwX4P16n0lTCOYPA1JQqRoMS8vaiiB7+jmEVP
HEoq8hZuvg9zUBN0Gjio1ryWSJ9+uiBEaBgTe8m9pcj1bgEK4I0LfIWkEwfr
4XIeTsoSNhWWkbHPN9O6B1O9dlLJZETnGKmx56C+eC0ABk0OwTKlhHPZfmIj
G/DhszP+xw/eTbJQ3e670W3E3TQBHG/3m0Vq5vIShy1Z9ESza3KM9HIJ2xo+
AmDbY8bqsUofqk6CsXuIgg2+M8cb7VqCPofgr/2IlWi2axJCZst+RP91ZUWe
Dw2M4MtRM1gFacH8HAhoweTpG7uKljAoL910zZDQQQ4juePzNf9aV/7VL2I8
/QK92QWujjggjouaOE6DJF0ON60SRwClcKfq6y3z8OhQwtCleD3mtYAw+TKy
bs2GonUncpcI2QMgPagXvdvTaunVAKISa3qhWtlXcybe91O2ujRdRwLkJJ8A
Q8ZYoH1BI8zh0+KctcCa7xKuZa7xZZduen3t2/R7v1rJXnLwkSgMBUWNSQcF
ldtiqHNRZzv06X48z+syG/uK3IrGsVKEsDwkWXXPcBcTDuSNdiIWxqAwaUN/
3qt3/Ym7Nbd8Q82Y8fl5NLM0WzmL+iXaO8/yQJpHI4vYYqukNGzGtX4xKZRj
KPHMvZ+9fWKnW1AmQ+KxTbDDOF7aem+fPXPMbs/kXeWiA292f3ELD9nvnD6U
jg1cAuQ3ko00qvJI2mmUGJ1qU/dT7d8DTBGAddpe+oQZjg285CJDYjpLV856
oXKEfHqGOSCqn+POBwk67K8kP7tytEDTZ7zitoncBucdHAczkVNif/mD0Vrg
3STQJq63fn3JEjgQa42SS028kLKAQ8w6g3SvnqkeJLxnXl8geWLee+pqrEZX
T8w2mvVSaH74d5GQKCbblRCdkHLQLrNGwcq8HNObZaQ4ithEgFHsY9A94c76
8p4sgyDTVDw0a5QSmV0UP+wWbV3AegfbES+JArcsDfAEdwnVk0CK7ljtKJnW
bhTGddR5eORDsbuGWMSiO9sSO+t4nnZKYV/28IqbqDEZSh6uJ/1WaMtESHng
ao5u387XFRlHcCR2l/X+KaRKtjSi47bWwRHv793nn/XkbaG2Agb138RsXoxF
zSmra08By5TdrSTKuRXGurXnQPoKfxd/mUgsoFTqG6ckb7hibndOTHloXiap
LA87hC+YopJ4Xew2AJ4w+y+fA9+QlbZ/o3xKjTRX/PMPlvJzPwPl5MsTm4NY
dCNiAbry5A85kOtXByfHqQTmze+eQGVMJZAayiujYWMFJf3ZrDn7AP2YUqmu
NySkXr2v/fErKMX9U/RI7QGwlIxSYH38DTsPdkVhNA5rPAcUORpEp81iSAWJ
8MBtDDP7jFm2CfdagM0yrMST0n3mZ4ruDaj8aO897ZiADL+WKWF4Atyw9yzK
jUNj1oCWlcrOZ+0bTPwqhimMNooUOpClJ5UyFGaqJJzgstRiPyePH6NdgAOn
vnqK/DXp9QR0SntHlpZ78obb0FwYkNs/B02xvuyM1GXxsil5MQV68C9dYK/u
74Imzwpb8RiH5xJpcCiPWTtXNOAYRbCTl0PSrMoLKSv6gn2SzwLJzZdaRg2I
ZZgbIOIRLEuBFP/u+nzuZGtFsnJ9SXGBC7lyGhxzoZ9FM5BQI+F3bCp0O2U2
97dnKL50dK8293iUJuNrzaW6A/dLEbrbQwfWUNV1Kb2X2gv5SZbT8ZDAkkT5
SFWXJsJjPEKOJV2N9e7WH5eKf4CfiKalkS0Wj24MgLTSU8HNmz+Mz+hlWlHW
kYw4cdAIHTayEEY/Ud2kXB40VnlXtD9mPKbf+XD6rnE95ZOb55OIdg63vtMI
SaBF1hKrToaCum1uhcO4IIQrlRT2gqRNEHwexJz7EqmE9vGHqVyd0x/610Jn
lzSYB9D1Dk/Pd1ydHEBV9gjP9kjAeVmHo2z7ZI7qaGxesXXWe5kCJLCnaun6
tawPgjxVgzsKcQtvzD66u4CDTHpry5fQihjoDFeURce2vWk+VFn1/4qUJTDw
aD1D709Rlq1N/Q7NJUXxEx9ty28/gD7OJSLgFHUvxSgHWMvw2N0b4bemkYDt
c+tIegfa8RxN1reGt1Dnso3UIDyHz4JJA2k3HE0o6Rt2m0JpqlhzUTh91leb
cEv3phO8+MKK676h1M4CpEVWZLrQ5LkhL2glh+r8/b0cT6uK++87OB4ap1SQ
rCzqKWK5WNstQBJ6zh2hOUueMaWRZJSlKPH0z5yys2adXScN6YtojR2JwS4v
6XPEGVPwMUm7ICCQnRxrBW2Cpe6c0ljxSpoE6b8nMqyw/RXj+/kDyXUITM+q
eACr2sG+gOO9dNx8rti69aiTL6AbGfwk9aV/7AdGf7ks7Ooob4iDIgU7b6GW
oRiB6cDaCSIQOzcGXqhXV2sobQ5ug8sg/EGd99sp/fv/9lHh3qI6Wtok/rgP
NjVsTBlCRBct1QRfSReQJuvymO0xCg88WLkosu9uM5UQrVCJGTj1b2OjM17e
1jGYIA895Kpyf3qte9r06PPjGxaWXYpc3GEF3i2c+pkwtNW7a0p0ddxUL3rt
VBfMrODIjoi44aDzP7Zz1VEVFT68/po4qMcWb7g8SZF0SZbWLn8u7vcJnz4e
5dlvmDNsSDXOC24/Dkt+8H5C9c5Cz3r6Q6bX68xcdGRCLONiqb0XhKFO/6Ga
RzepWEdTOBmweDHCpwmJpSBmcXFwAgkcwWL8t2VLzSr9lv2PTN15Urk5dA+B
zENBXkFAZZwqJausZovS89An/SqYASO6lJBNYbFJ6sFjV158GLRqcF0Yy582
oElCrKK1i2yps6J9AU4Rg+FUVSdv0tCoXGmDm5avt/H+IwWjPu5qbRUbtYXx
HRmizuUCYM8Awh4vVde/cx0KWdUMuykh0iKb3LMMEmfyF3HVpZTD0xh+7Dep
zUZ+LGXi+lF5lrg83sML/7A7QaFg88TwbCA+//L2OvSV12RVChHC2wlat9rM
HucGZnBlTeyBhoFlqwR+OKxs7n4QMWK5wbGo5KPgq9XLSW4UAv1IM6o67ika
36Z90QGyLl9icOKGtyXl9aYkYDRZQQxvfM3RE50lLfY+IY74i1L3W7/yKDJY
tpscP6vbU+yJzunDSGrwVZIBAX/oUw5SzPzgVu40Y9JEfNXeANfkR18hhcf4
qlzaqlKJuW1oajFPB029xU3oSwpmGmyxZYIM9rSx9DdlZwXkkjt4WPyeW/D2
kKkKEvemFO6q+7aUzPWn5ESpIYuFteX6hLgXbLlEyp/gfqzmnaYBQT42KSoF
y1o5B2mYgbF0x7wEnUoyoygB/NX9cvdpEmoNceoSUBVZuF3x7r708Ad2CZ7I
yi3HEkaoScRVN1Og8AAakfBjiZ8hQ2sEVd0KybOXITm4HH/3QXdZYO6ucZ2T
3AOaacbaa8KZ/hAC4qQcKQiiRZ9JZQ4la9NHKeg56ikcEdWIo+7v3/fM6MBR
icY2zrcap4SZ6qr5F+VvzHDq6oz7Th4jy8QpfHCfLB/tCoxXP0zy2q6t0iVW
Qt8I5u0g6AKQ09P71iJpEenRXyA9ecdlcInxc8VgNyl16NiypNHDM/8jll/P
3HycmKeUd0cwxz5/Hb3p4trqVSqjlIB5+VRwxTiGjWZBNv3za7RzPuG5N1Yq
6u5E2ocLwuJlDxw8KCUdmnz0oBGe2juk0UD1MkiREZ5cDh4Y8SGupmjR+svt
DA1MIuU9YO54Z9T5laqKor9nXv+HqGmJh/62sAe41YoOQuXOpJLPJNfCoznc
meDIQFrSVCeIRFkAaW+TCknT1aqYxrBh4Hn2rDPbef5MQ5rrdiel+ymiQlKA
wl3O/Z6xjmu/r+3LWruBZrf2vksGvfS0wd+P3n3oLUccYDe+pZEbKVzpuff/
POYfs5WdJeBI5WW/1FkXNRyVDynisEcCC3XNdKWQVx5kiEC7eyQpPFJyJ84b
tS9VuUgcT3tsimS2WLJXLOpoPryodU46KxJdtfqZOlbNN3Hl+Ey6sPFs/9LH
J9dKMt58rkeTUqeOzTv6d888t6zEnCe30PguGyLhLbHIZD7hw7Joc3nPGE7n
MMK+2LXxtj3UNbCuPOmEsSOuMxj83OTgAyc05lPqf1781UfbDu6TjhjBr/6D
/jfu1wTz8xb1GaAJpLqgFUjdQH1fTSYzeDX8gbb6TOzONqoMcocISBb/Rgtt
hGboEV156EGc4BMSuekYvrIFW8bfWckTE4XFm34aL8haEas6E1zMSHEA3k3+
j8N5cKDIZ4e5eTHTMVFOffqV5wfGhUuvdoq+v+vxFS84GGOeuQrKg0rEXU87
UbJ7cXzGL24Wd74YxRxxt6IFbx0zvMyJ5PBqcMnKx2Tv8DasU8rjRdm1/TJC
e3Vk+MGguZemJ0WeTsEmxH3w93499REi/Aa267V5cbQ56JvmJ83KQjieJrJG
+CGX+X/vQyWZx68UJ+LPiS/4YVNhwE4juUAhEVYfRTPtHOEg2vezNMMZxPnC
e0z80xiJD4BUZaPR62NNdmMlihv5jSYX8gbQBmNzBS1LfoPf6tLU+cPCFe9a
a729l8bq1UHEQppiyaWwXrXHczFIwfV7609A9nB+GfoCvx9I17LhYmeg7L/2
SP6dXkc8+DhyVZIm6X6CbeuY0bs6KTrpBxcCeHwrz40fSJReXhP+z66WJKSw
FzErQ3hLJuQ2IQFQwNX6lvirkAEOYokACKLXAGWeONlg9uKgU6T9w06DDNhT
lB91enWqibxy1YNxIehdllguNJwtZLpi3IjCWCKTtFZU+f2DjxpquC+1kogw
p588JCiLpK45jySKmSdylfeX9TxBJgeVnwJPMlPuQIL1Oq8CIUARLiYiUjMp
BxSQcF6tnjx5XIVQW/L19rm6cQT0FvNMQGl5eIeoM6cjdzyEP45KK+41ErrQ
exh8AKTlB1uTNjbLVBEK6+tremV+FrfVtpzwqYP911ZDUs5CTyrLkEpjI3gS
H+5a0CdCxiQu7+0iKJh9XyitwOPfz29CS4w4LVRRgdNe92HOtsyQy2TyHVpU
u/J8oMGrhrUKko8lLMQHXffsOQZ4TmSC1u04+46HrNzYUNhcHso7oGPbQ6kq
5DvJPJCk+fUgJtKU9CL+ADeGXTt4ekBVkmxFyuPtvKDcynASRp9ptRUPOkmQ
bb+JdbJ6SnAlTOovhtHR8SnE/w52mg7Nb3h3FQEnfkFsL7gnjGWl+5WLlsGk
Cprdr0KxW7BoYgAF+7qVJl+u1Q/fez8NRwxf1ED6ISO9r8cAN/Ih+xPub8Wf
AXDQn2eqzczSJDc3Zol1FVP+z9mmvE30u0FNC22HUBl3JYpUGoWrP5j7oqwm
yK5sbGIu1UyXQCZBtEYK7ULXzOo4f9YCcC9WYqnYaDjCTV3YkgxvlD9AC6f8
7frYDuCL1+0e9Nmc4nbgPfPJubXr3qk9L6AOXf2mBKvbGIbVd6a8etLGKO4n
PxsUVV6JQjsVLsOTm9Nov40G3+dOKLGepAkWmJL8OmsgpEktuT+j8tdajSd3
Sa3KYBnoZ9TUcGa6/amSD1JWB3Ll1ScDIGpDdT2Rgceeap73AbAm9YbMrUPf
/PWZAO1BB9nDAfMSMe4bOx3+F10UWF9MZcbnLQPIq75rFbQpvFEKyP8GU5NJ
dhcOk/f0wnZacO2OCbOGQd7DA69TXvqp9lvyoW+HUcH8Nk7SgqiODrzdBbq7
ZnpJIqMI5Mb6U+1Q11z5+wEkyiORdDWlx6QdX9djlgkyQ1GsszJPU6lM6HpD
6iIoFF94Ibxnjofr2VkTTFh72Gf8spwRb2wnXgUejy9yhiOsBz//TJmlXPBR
mbHazMq4LNE1tItaNMXJ/Hm2Fd/wLn/A/N219bFwXlY20tOM5TSvclWs1OKh
TcYNVeVdJQyHKs+HD1DqgLq+BIHHyl7kgVUyQcD2+VUlo0eAMQ7i5izonQ8R
p9qjEe1OVA3V9zkIL/ZeyvM9UpV95DkV/UyQy2bBUgDjO6rgh7/6PKgaeUXr
an+dJ9MJgj7huwmOWj5/JWZg6eZbP0zEsmpeAKw0L8C8d3T1e64MjyAyrhlh
tORUsEqkQGDTYz4kkTtuubFE/yi8zSQ+cmGkQB32s1uzp/0KvwlYYaJR3Bqe
kATINIRHuf3oQX1f3IF5o6GUnjTPZFyF3bX7esuhQv3QGw1f/WsNrhfW9Fev
JHhN4MXqpSeRB0xgv2QFjXCXemkHyUDMYO8x4ybw3EtB2KaWBEoGXrXWVEgu
aHHAbYgf1BBB6UTXmuuNXRcbDjrsnbTLL6yIbN4NoK8f4WjNJGEWI1Tj5TQA
vcrF8g1obkxNnWkkueXXb2FLCpXCkDFTOctExye/ozzUOvmj2aPuSFNos5yK
f817vB1AMkEknw1oa5ihvlb+7jyisnatkxqed87wF35HEIKBYh/3a+VVi1kt
FWtWoKecXVUsxCoO5v+g7WrHRfKNOJkKEOgFUYXC2PR3uIXEgXu2ORXTKLuO
Winj5ajakH2dQwR/HjxvZChfm3fADCJRPog9iAlCJn3DUujkIhWwS7O7KjYW
WXefkmZL1xHGm2P63Zn42+4M70THSgait0KdFonWw7rPmjCUJyt1LUh1jcxt
XFyqWjJVZnSiPKje6Gn2lNlJSdS+9hxUVHZNwRIewcxlM/El1IuUG3cU5xtv
3rhMwTxGOIq3VUjkZ0mWZkfZgt2M8MmDLUsii2ELjuo0XvvvJOOOoE6+VexH
9sNyShv/Lvc60fOkdjUAs8P+fglQUkbCdTmEd8ECtn3GN4UyWMooGNluaKTJ
OIjoEURtZvNB228IfMcRgIBUzv7d/0gC3B6Bj/Gk2THMcLMjtF/ygqFpvnyB
WqHFnvqOwh7m561LLMPTgjBrcf7M9CwExpqtYs6DHYp+xjALklI9i4J5TZsu
Kl6j2HeAUlfO3kv/whg6NtqxH5/yCJ2OtjYtAwa4Y5HXmeSCfLZky2B36siF
frCp7iFDAnFEZzWmNQUdVXhJzci/BAY9t1pf1LQj3HJoBNKRW2W1LI6+baLc
y574HLJOYSdGfgEKlXNVplUJUmgvJHuqEv2QU+gwz0a9Mp01bjApZI8o+TNG
KUFoheBJHB0NunA3U3tDqHa1EdaoM053x24775wG8JlGRXp/+2WS7Tz44/RR
ZwtpWxG/IRYvqlgUpMGh57jd5S4vPMPIpaCiKF4r8jC2E6pr0kUOy06Gk+lh
DFM+pN/PJBPqf0CKewJqvq47VEhZXVCxKVDw6mkEoN+YWz9tyCXpWohMNpUf
eAd717nQXfcGo/X8X1kJZ5M+wNoUygDc210b/9wIn34f1oWpYPvdlJFLN21E
MVNAgSHDQ55iwfqsZQKBZcTCaaBm6zC2sZWxXlSR8hPQgfjTB112+C7TvwHo
lAWsN9yMWLzlfpTHYnWuD02sP/YRDmdmWc0dVtwW1nKw9vc5ILUwnlysIpEw
DRYEjnVqB68PP4PWdVRPknz17wQr3d0v9lOZ8jJtCJSCgsKP1xoCsziY9FdJ
pWgwGb7JEEpITtxnbVtQJ/xp0vkEa9VBn8okLggcdmIudF/5xI0G6tQ4bYTp
zRI7u0KfUYNGajOF+AzyXrWxE99zWVrNt252npZLheoPYn5eF4SdshQC0r7Z
T3Vzk2FOiS9h8K6kObT3pxEGgdZxNq5wRRZN/NDANQgZPTUmwhe/+qpSqC2/
yczt5UDK2A3aFHY3Wqz4HpWzUsUa1Dhcq9LukDYVGRTLP3mJKl5iRKEBvFP9
kuA4Pcg9CjHfH91Xb2dneqZvNS3XP4VRMYdulR0CmHFy387WKWU95a1LrSgm
pCJwVcd9cD4WwbOqtwc1GwhPO06ZIJYqTLSQPWx0hRp3ARBaWjEFusSNwq56
TdoXfg9dtFjXum1Mq56IaGU3XwI/ZDvyq6nfOQgwq6+65JLkiu/WciwZIAZg
Yz5PKGsN2J9kEr4UCccrc/+zihcds5uQN9TXssf1qhM9cCGh1ftwHt0nwNyC
KLpFyhGiPmjaWeUNJ/nMwwFxNHW9nf/m5BnLOe7QSS2d20QKrZ9W1VLzgrcq
FS6dJUS/QhUXVfH04cJGA8wBlcvAlMBmVZiBmqUp0q8FvUWKPv+FFTsSFs/C
FjkXECIU8jECdfifQYUayKryD89F/EqaM3TFMpq0MTV+Wf+z+ffhOtYK8ces
f5Vd/P6HAGm7BnY182WkdsL9um7Jqd9KVgRwhXgyLl3VDBsTnMm9z0X+CkX6
QWT2ozQwcSDGk7slA8PtM2tv87v81Ng6zTPk5K74sAOWdQzZjGI/HsNY55DC
FzATFSWrc9vSFFxCNgeZU+9DIgF9hWgrZte+em54Oq1ZO/9SZRkRBji+JXTX
MOLEZJA2ewfDniGccDn7KJ3EgXKOKAquwJT+mi9xzoOCSx2nv5WuVjJm15Ws
/vXALM7gzdA0RC1ih9JB4hUc5A1PXrEa7fGz0MYPGkDbju8K3k0AVbOKJBeT
Jk8SI+mcYFOGVBwmWBoRW1C8MX/eorTfn9XGt4sHB+lrkovx7UClYoP35w0L
Wlszpl7Dpzu8K+kkEL9Oz0Lj/O8QgKVt0nuaWslc5gzQRgv731dtJJWNZAhn
vaRYyJHFZnFhKramGUZ7Y+wfv1PV3Abht5kpsRMxd+IcPQbKVRI2zH6m5MwV
AdMsJM9ps5cfdirfOdIX56e1Ckvbbqi0jdpqbQWp/bqyD6qU0jtttLmUktgo
hLhRFJdAcF5f8b/gG+EhMr8CxqzFXXuULE46v0gUrkzArjw8lgwFYELkoQn+
1xyvAvS8mr4xoQRE1nHrbpXlED1hADOgOZUqjemmlspudzKBY0u5YnBHeFiK
xDNQ9gcqqA3unEudoeQ2VCiXZkwfqC5ibTrtPe+TSmcV3ClrRpNH50pID8j0
yUN7u9i9/UDS2iT4lau/FQV8m86fmNCDoAxWfBmwVflSHta1LowtfTTF/72/
L7iud9ccbo7zX6Jnn09deue5xbFCX1lDAH1guEsGNbmGCh3M5FVrgEoXNI96
lOVrx0RyA3PFbRVq2sOv7v4+gJanUTmTqWkIfN6vjuFimorGHjkjS/d4hffd
hav97EpeDsRMKLW7s/OGy+ZP3/7oQQN3xS8JSJdaqUw2xphT73GhlVEI+Lgi
16XksSgOMyzt+ASvJjGy8zfwV57THC93t9WElGUJXLiEzeIEsZJbJa1Yyd7A
Qk/DTevRSH1fqY1W1e91Q4P0GyBsF3yEpVJJwE7Gu5zDf/T9ivfxvi2wtpPm
LOy0wAFqXXv0oQswEkqtDzt5iAzPK8hWZbAWSOS1QD4cIl6taZ/Y6vJ0BxyD
6LnhbxDor1gWZM2C1zJgAXaUGJCFPaBYsRJbRqPeLSRqTpHamNq5GTiJ+qOB
6vX7zR4bUxDajaT4Lb672yD/Shzc0f2H2XmLD+bI1pkInqrLnbKtwWezpLlm
1QzPjgJOjuIIDWS+b97fPrp9H2brDVshTHjdEB2etw2Pnh2E1M0GvmX30z96
39Oq/LeDDvRpmXhw8JtVx40mvtYW7idJ+bkLR7XVupfW5B/PhEsutpitN2vZ
8JumsysrR4H53CWm/PygBhaFKTYgZNIpW/E08NkjTOJZ2VYNxuAPYbi8W/Vf
YhcfWUFe1H8hd5qLhLNJyLJBjEcx37oifcgVO3ChmESi6UFxLW/FPHYAYxPx
uLw3iSDBpHizgJHxwY5oAgfcdAkwgg7tREym12WWGeYwWFiU1NmTjwGiohcr
SaUUJpD1+d2ehvFeM+mgHtqQqzVk848xivLgtbahRm54gUIokmvD5XWsFrYD
3/E8goIugV5RzBHb4dMTy/QObk8UurLc6EmbWDRqEOu5QoEXZAatJhATVYkx
DMZdzLDKek53Ttrtgad3KY3YcUTHrqmQL8Y3m6cqrLonJV87dephMgd1oSsI
FYBD5aFVteDAHXiozcPPh11qzUv7P3m65YZb7B83vI/wSdeDYFYjnua9+2dz
XeNpXqGZsjDTRCXODMGtw3gydg6eTGVh+tfWZBEQAHmCffzImG8YiiU1elnU
jrMrM8yYcVI7gQkJ6tpRXPgricKcVAZPoTZfFvE28AnCudKl5ZX2jAchZHGg
iXFGakxFOLAzndWyeDCnWIHcsTouPTHESQqg3ocitG7LVe9rWfPYCX4DIHuf
a5Gq9g/bgXeq1MK8nOdYg1/yfPP6JMGD36sJ9zg7G05yplQ8scETF7SFYnUb
QF9n6fPVAGku/vZLzYvVeVXSQJJEMwNBLcodtUNC6YE5IRlpjAQeYfMJfXGv
B4jhpeoQ6vveQFS29zb7zUUHQMO4oi5NtlXxX7c3SVP3G3B0ro/bedt+Onas
Zkf5DzQxst3YdQxq7N9WvTwy/Qf+qSFzKEUoGcB6E1LYzs/KrFS+WoQ74+7x
i3RMsTvrbBl/Q0rsRt/iLzxpHWWI8CwOjywGV4vt6dKgsg1a2CgYdFj9UB3n
31Bs83NVg5YxchofPrzNtIaOsq+WGnvHFm2UoejgiP8ECzOPKiy6xb1U1E3m
vKb8sVe2zv5fP0/6X51Od2W1DoA82TV3FyN+WmexaX+4ESU/GCAr9gWjPcSj
TDnnTLVxYuFP6JDf9kE4eFLgbF6Ugtz+1Xqg4J8ApL66cznKhxtaRbrFu7Yn
t3pMk3CWAaMuDf59k2W/RjnQkxnKty+XC5kj4m5/qrSpay7m28R0Fwf7WFMJ
W/3ttxhVU61ZL2volUzA/ACxlGZo2aJqOIqc2WAz5jM9d7u2CMNfYaEp09TP
UosTK+s0mksbkyh28hfWuE9xzlZQlxxVVXGtojbjYJVYjIOXnNBc0S1j3LlK
b0j1ueA71R4YzeMVVJq5hjTTyrqN1fYdNVEeIRMPixEygeLeS7kBBweDaMkK
hHvvUCDDehYltAGbpLIU2RxWmBWzZzEpMmGPe7p7YlJ9gXfZGq7x8FEKWk8i
4ZttN6LEj4c9/ZI6dyPMM1RlFKN4wolaAYbWquSZhpTArNsNn3O/oLdXEvPs
NXW017wHiIAM+PBV6Fl1ay6xG7nXP7Ka1MJJT4RfQz/K9HmBAe7QG1yPJnla
DExuYwBRLPHu7N05NJ2ip/57osVjdlSX2NsdsRNAUz0mv3jT9VE2rRDc7p49
T3Cloi4v4aw/LI/WaocLekIyZv4Z5up8i1B2kgFWgQzJpnHVQZuFISvn2L0r
s704xLLFPQzVfktkKB1xrlbSYz06qeu6SwR6oZfzp8700y2rhjfbvXHw2JUs
Lp7DcW5BT8vsnNbSRIhkfvaIsyLU5p0R6aFscIdIb2nvB7bT/Sly0pZtSWZk
KJnBO6YdoVgbMRVBUk+DT8crvmamHCTmqY9WhkXrJssVMgAkEJ0Gd3srmfaG
89/npXgIASD6WPRL7G9z42XWnMrAuspYJa87Yq7tWPQpmzRu9hKZW3hWXn6V
qJxWCo4DUF+1JpSb+1cqS2e2n3xSu5omkkdC2AfXcBCAKMDxmlrgFfzEHjGl
x9QUo1Mtec+5Rmv1/4vxe+LPpU25zYlpYqPZnL1feTa68WE34VA75Tz7w4dg
iPpu2AaT0Ce73AcvS7AvbshAo2xvBVoUR3OQhUKd4UJfrQaeJCAsJCLxV+Oz
tNxqS3kRaGdRB8EyLgCOcKMR/jUhDno1PU6C35XadRwLss+bCXHotbj7Ut2g
bKA0IWhO5TQGnA0G3xOlbbR+teRHJaTz8HSn36gk6D5ig/arXfABDdoIJU15
GurKtJr4ZsJ7WVceyBCLIhW6WY9dLGaeWB7hEfGMYCQ3HCJ6C1vDampE/Ki5
qRnmEJrHjQ6KZDU7We2zrJHZNRsOtg6oI/bryrWLIpiWrGSkR1icOtbicwlO
kPg4tKO1gf2VUl2nDZZgND++yd70aehCqftuFw/IZYcR89rvnuyF/W+/4Dc3
a2C7TrMv/7Kw1GQ0YB7W61LDTZXzwX95swUVKD8xoPoJSOaTdpfVWB/6kyEe
uVSabH8k/QwlhZYKlNPvpYSEu2xSEYwQ1qRglLl9lX9XMCV61AT/wCDEWhgP
Tc49NdBhu/4YdHy8l4b+VR8q5QsRipqD/vQAE1SLe/q9h0zT94lVkKooh0aX
jRyI+5+kDS73uL9hRT+0QrscY65h1C4houvyXLZ8W7XMeNkcVOkAVIAcNFKI
Hno3He4ftcO8URSrUEKXKRU7ArE7/dLm4Ni8mSUkRKw9r0iVjbzJF+mFt8fa
+CO3HkTRokM7NcMKcqGt9tk7m0O4ejV1IvkNJut8jK2eSksZKVkwjh83yBBE
vwxr7MCpAq8rAO9RgmejBFOkDpegr05l3JSWjJ34NXnR15eUhtKU1iN3kbRD
pYijUy1LTMFidgP8kF752sjMyMNRI5cIXwTUxFXia/wk29ZBinrlGXc9sIQ5
5JKlhI9rpcGfX8JxyDur3uZKMjFFOU+v0PSgXWOgPrt4UYWo9GhhYd7NQ4QU
9iBKOvslDNXNXF17Ay3aMJ5uITGlLEp4BZZCAmB4/OlvP+ndjHwrRekzHEPc
1T8CJv/WdBWsZbe+rS0n8bdlTxAX3H2YM3da+aTnK4cqrnZg2w0LjemKp+4l
C2EpsodKaKko0NYmwLkUmQ0BHs4N6XHq32mfgcAPbh8YbATCg6ZKgzYPqVMt
XOxa6741TeeaT5nuuEqIDEP7j2yNabVEgRyv8m4qWfsAG9ubok7mRiIUrv1O
pxIW+JMTBCyIYZJVS8O5zQ0ohkw/2vODCLg3GCfXYykJpfSDQY7LOKLyVXsZ
oMH+eQDZuEebtin9WNXB3rvPbmAre+9BuOLemeYJWGV4OVs5W61o12FxN3u1
Hb/4MqcKVlGIrW5LpT3wDkIIIYv714s34lFe7L9ZQflx9HujHdduk7bV1MwZ
P9YsCAlPksJ3EmDj5w60eTnrmzBnp9DAWcE9QuVDYQuTkJgWdI8PrQE3clGR
7gZyChd/+y/GAjX/o3wO6Wd4yGoycz480dYTso9icw09mK/Z0Of8NLw8uBKg
Iw3iPCjPw2/xcp5z9PdFjzERh+G9Lu8hfwJmxYJKbILJice93nfLVWY18QEI
XNVauyzlJ9XjdpqJy1L1BktAYGwyxGdjcL7ie6ednvOeRJOt6gBPyumjlFbJ
jl/8vRPsqu3xwE9AAf+YaABCPP3zNMiqUmF9aW0vuA1g0UsIa2vYI78a6JuE
fAQzPZKTse1mcwWDGyYpqE4qnz7REL3R8ig59mcQ7rnxClHt0DfUB3dyZcvk
lZJ/+foduUrV5nGNSnCAn2Odlmw2oL3XhBHvwIJ9/LO8q7sWMsv8ylS+aaXu
5Em7D9wpdC4DGp/pXeE+2wboVcnmzhafh1ELcjkxAVEoi8ld3sf155446gWr
V4iDIVw45EGPLMpCaipJLlN3viMrEHh10fgAm3+9E4iCRNKuE27L2/4zFjYv
sxyvnikZ/kIlP/FwewTWhFBShTpFguMTbO2sbGXHi5cee+rR3vw9S96AoO0C
rhe54gTfkm2ydTc6otgSEJpQNA1bHryZa0QEkHLwV7Lh5UbAA27q8rLb6KZv
clFL4KKhjRDd8WDGsZ3OVwbLREd6cEzKycYz7HVTNUB+qKfqGb27UQhqjt1p
z6SX0nFTl5cg00E2ew6/Y9sUgL537igg1FEBVxR2ITMbZm3h4QfPSHduWo3f
YKMdqtZzs+tAAet0GnIGlruGmH9WHDBOJUqmOW/Nv7uQFZi+6j+KcybF2SON
VgJxcwYl4/asY8amcH/ZhH+RFoo2NCelvtuZu6+TkBAf+qEJ0Nxh2OF2aZhx
W6nyKFBo9EgKYRB8U2BHTxXjhUAcegQz2hQyVwwOSe9BTwvq2QQGQlix/z6N
mv6C++YPDtvy/9x/VJ+Q8p6dWUQvQSfRhIOHpoCv1tL1LJ+ZOPN1ISNNolVF
zw+dbMhRaCzHI9Q9P5IDzPi4BHf2OnVQ2sbpcm1Tvc1KKTvKbTLa2P2bfXtL
vBkusJz/Zvch4HD1rQFSCFdab6QAcJNkWTxsE09QALg8In5QgSnQy/istRl+
3PeYBVEpBZWaf9DfCmhiNOuaVWaIoyx5wyo5Y5X5KADvc6aRFaSSfmbs/rK6
fMHtAWVH00WaDFcrpZmWbvErIOlEr964Lx+G/ac5aCjvW9fT/l6xAAmWJvyt
XCVYU3FzNv1zp5TTJ3l4hx9bqMaLdcJJPaK7vHrDHEDPdF8DHXDJjU6Eqd1I
Jgsus2/PVHNPJi20wozvG6uCRuAm1baExnkT0GptIbOBJRLjkU3SBsvxgdVK
NjyyDtLa6Euy+l8c8MYpXuK/A3tVi7px7TQ0BVdtqjE8/v0agYqHMvsDjAy5
0/tKVyrecWC9V9yJ/ryRemQf2UbJVXQsGtukbT7dcRemm5V3zGuN0LcAxAKg
qHBxhiNEUtXMFTbitWy+h+EipXCsyp9cvN1E+kclbW+fEn8VxDjwi7hVJV+m
VgIZhVLdc2jGkfLUCeIC3jVcvvGTuJj/FnlVuobqSRzmx8EnrDL4xYyDd4ZC
9jq4bWB+6pT+dBq2m1orpLC1MOHskFaN8y3NgtgceFsUnP53F1Uknv6moaDi
PWNBiG8JkKO7osLH/a3O9l7nppkLSAC0I7toHkU2XH9v/aCA8WN96xvH/9l3
MRBI2uCAP//pius/Wh/cOL2Nn/TeROJ75H3IEbJsDBkNo6rbdj33tyfRFubr
fwEJZwYBRGftHHAu19kSf2L7gi+2DAEnjjTtTwjJK5HZSiB+c++3BA3DrXoO
xKNtwDsQMg3jNJD2qLV2JoOLi7ikwHfwKTKNr1mc0j0/yIFdUjYC9m+s2Yys
NkOUf4G1k5wEK5rhxAFKKtst7iL59mCDz70iVwYlL6wsHDQrZJ802ykp3H2P
vs4Xt+4C0bDb9VLcZx7mtrCtfx7VikVhLrKUw/QcaZQk6+qc4/Vd05BA+iAN
YKAMxCcr/wx/A4w49b+LoZKwC50y86s2p1AsRL2R0d3A1SZpCNEAGBYgmWg0
4ZVy1P6GeixLzG7ckI8XmlXy7XV1TGBDGzr4kl8SY3M1xSqmK8XNe11/CxIr
z5wCSrZ8baJof5GQGWBnojQ0HLJr6cLkVxghNm1jRlhTRITGI30wTbWggVXf
MIYzqvlB3dphVDTT7r34rbfPgjqoObpD7O7rOmOoeeABAG6U6mWkECYxrXmH
w0qHNLLRDIJ8SV+UlCjITy8h+unS3W8tq1hGgvx554BwcZUQXVgNxDNevD6j
C9P6yzAoH6flBK2M+3dFsd2R8HBWh4+Xz5zGUXFStBOuL6DeuZo1qv6OepdJ
iooQlQzXlgMXJQAMP8axttp6C1M2ePwiZlDBP662f+w0l8nBpVNjNPd1VYe4
tP2q32RZ0Edv+VzKx1AC0521pX8b0Cj7mVNAcBPKsFZerH33re0VBJAEKegh
l/7GrJwFXJYtqoKAsOzm6mz47hZaeyRX0OAD2OyHGtK+OmFpndFAepqFxPqv
AFSHpKQHDpW3TYqYEUMTaOxqEtHDBBqmY931Xa6hGNKRkJRT7jNWT8t6RuF5
/ZVwnPjN6xiDvfs4KaZypbtQDWXpPp/INClMHARTLki91FVVsuyDBpLk3/Cb
vpFK5OIzR2206KVvwxab20ewEj5FsKCYcQVxQkR5E4eGsM7NKoq0cmLn6cds
H71lkJ8WAuG49D7bLD/CNU/zArTrll+nObcOui0L605BxeYbnjQxAwmSdVlf
/j+7K7OZQ6lGaT/r9Sk40OlkTPR0k3s5Oi2DNE3yJhuYcSQRPbprQnhBgCzh
L1wkVWIMwm2qoLaympsJVo71n/H6CjpSTYOHtaReV8F6RKt8lzyXOSpVvIYA
5bpu8Tm8hc73abx2ulpD51qC78RDgOQqUKoaqqyQNaJFiq1F4O0emhWA8SfE
ybR14Pv+Rq9yXrJcVT7/cQ+Pp3+c/uvSB0GJdvS25jDj7nqBXtTqaGJCFOdC
swV8ocOVB+foRW2Krl04ghAjiyCbhJmxifmVSqGmxh/tuHxVsRCfUBQlxnIt
qHZqI+kUgzJKfffLHcRcvQUFpgX/2kHUHdMSP1yKzUea9ZB8fU7QsdzpXa9Q
rNu8Dt4OGuEl2dO+lDnwd7XZOVZjoBwfucB16+w637BbO4QHHBnXkRZhifgy
CkCcoI+EswCsg5bsP4EtUVAE0CkyCvQyxPQxYt5u/5wq1iGidC/aUusoGwUR
KBUcNMDpEvrc1B2MCzICosuyntAaNBJWDgdAM5N/skYagr2w4TgP0foFLmH1
RvAZzpqHBuy6wb9a4i2kog7KeUpZi7rtaWWtuXghmTATlIrPR/W7ZhFuDYHg
RJFzkSN9N6itcetg4RH72J796QIXxuoIjhCGPho7I5uckFTHbdDe5glFacmN
zlN0+3xHwLTOe2gjvyTAXCmPq+Ex9leigE3CiBfiiTpWMc/Dxx2tCoz5lObh
98Rb9FhwNQlYF8tFxH/S604Ks58bCaLuGvZLH/OBSML0ZNUqXiTKg0eIeKRX
F/fIzcRGgXEMmoH6Q30eqiTh+3Kq50y95NqoTyAGPog8Jkr6PKlvvXfcYztx
2GSI6M0OSIaJTRLjNy1o9fSw+4O/Z/2+tTfUTA9QtuiFUUyP1TDiGzNJIuQI
NvWgpXVQpSSmWKFMVDwxW5/3thyobEDZGDWm/9oc7kdO4pfAdjQ5UavOA/MU
IdNsidpDQlvJ3OTZe3/LHjXIp5+wIbCUUS7e0+GKSHsL3JvBZSULFKeDICvl
7SdFcMl5Bn60Jn0a6+jEzUWnJ8YbTEgw8Eu1yMye5sLEg7/QdGOhUUd/q867
Na32z2AxKqI+sSx8JpTVJx4e2aUFt0Bk3T05mFFWOqRlhl0FLRaZsRkVsi5G
7Ec73PENfVHLGd3C1EWvF039kOhXEbb/BLCKCOxONsFUeWyEG0jL0qSg1XbI
cPemqizqxVB0UhXcWIu4WCakXC4oax3pY4c1Pzcs2VsxBrxLjX+BAQdfCXfU
Aivc6sgS7eE8HuGzcGWXzDeRzGR6kFCYjgoJORMv9GdwCtOiMzoC4Iz4DvA3
DDLXwy3D7K/bUIqCLifDPaVaO+ECU4hQJQ4Qs8qI3TDD+HxpGbEbfLsHL98r
h+Gy81Ll8B2tP0QMjh3/KOolI6oStvoNxnq4NRtwzO+crHQB+LQJjd/HG/vN
z57Qyi2ZSGBgaT6hdPheqYOnfT8J31cQUiYAIJWZm6Gl46cOfkKgu1rimyZJ
2EKJFb68Xmck1vn9cCmwjQHoHimaaVX4YERq8DpXSj36ZblCBypR9uaB4XuY
KJOfvFDOiZfkcvKsMt/56K+HIc/5DvEcNNePZde0ml8R7wFi3O7/HS3qPeU9
GC5iVL52GhTh+QQQvEyXMJigTsdvT01DzRosz1rR1ipr0ldLn2L5we8a/BMy
ww8eNznyhYMjzBYwDGOPIItkziMze68PhvwhzAJ015yRzdKK9TL/tn9CvrxJ
5x/NKxgwiCYlsUSHb3jfXpTtpgUSa0P6mp4451reg8V9+rjgRTxvyYswEXv9
kOnBOxLXW8yu348aYWUHZ1iC2qtwKaxaiAgFjW7Y/YSi2OkkoAeMb7xwuY9j
Jm2pD/sUS33GWA6S0iA1o3nhXAl4Uyt2RCLyrEiXE+M8FLvJ5SqeWGcYJUf1
yk4+wPlyRIjkSEZJQcnx6KcFaaPhy5CJe33VFrttEluFlLcCApFUCD1ZSOS9
L6ZLUEo1A9mMRkW8+fQEIPlzT+Y6c6he9St1GJC4OiH35SSkmS/0seersa4n
KJxGfC+797pbo4VDVn8EMD7rw+Bluj7PRPt2RRHpkYWfp9ZfLaU2ct0MeSPd
8rD+BELlhZg6ixGMZKsCeMgHhwYwWDbegOG6RTlhJ1S4gV4aLhspsBDlLCBI
p9mI+/9PJESXTEK7TudQNOpC1lUwTQ9/jHm1Aazn1m2wk7m3Drk2Zvm6I1xg
5ntRXCPhcNPksZgRA7Ajwt9sMji+3Uz+2DstCWwrGNo3X/zSwJuJzV4Z2afG
Jr0GWIbgiyHx4Snkgl4Ouhs8XvhLizegjH6n2nGh2cBqbLtMBNLSw1jgpl7p
qVYCapQGuQUysFllb0N6dFDDagNIjAUHprSBP+c43ue1Y1tq2hEkIAl+E6Zp
nTLfG0UlnBF2K/h+xtMkio0sAZ+DOIk6wOP6z4T7BeRYoPOLxPrll1BPj8yr
1/GmX0mKd++kaMVTFPRscjydaBXcqlBYAerCeBVv5DcEM4j/enBAfwYYBfOK
Ty7+WTzTEcjftR3/zqiefoNUVm6sM5GK6pZFw/7q9XerZeWhm1WOvSrXeXgN
LZ5697D/F5wn7hlEffL4AJlBxdBSpZpBjiAM9hpmyOVHuVqKifEwd+0wBbfN
7fSObQIdXgmByu3RJMADYUwQ0JHL+lcqI2fCfRMrqoNo9NwC3kgfBTeup18g
JTzMDhYjo9yF2/OXp8MKyXfIITYhy56TNHGnFgqTzH6ORiU7eUYADzBBTH8h
oncAzlM0TngL9TsW6stlyZwIHnuyytg8FJSZXms1zExJNWAAejUoFOhKR1II
dTkVL/E1nLOfWnA9IOsejhB7esfITvAXFIJVw9hcbg/nYCl+xmBb2qfUW/nh
O8DyHPpp9HGNSOjCmhprF6LV8PEL9TOyc9/i5aKs4tmhe4muXV+zkoymTiuQ
BFeoXu0i7wfqv+LfJ04OGBxJOXIdyDpT2xmSuTt72qB7vgTpz72OoslXW/Uk
+kCFdpaxa0CG865Wne2C//Pn+iYYLmHQlrH+JRRIAjgbDc87R8G+yXjiMV2u
EVOQDPRAmlMI6hpwNs0J0PcJXj0sYIcC1738TUPYAaUIFhpXfPrLJEkS5kxq
57gxF30yMn2pXBIJLblPx/zIOFEiMqnBH8TIeSJBHCgRy82du4wfaO02gVlG
KSMUcT2E8PK3meod/LQfi8WgoRGNO6LrKELTKrENi4R7ve+8XQjNTt77zg5I
pEZDf3hBJwJRANNsIlyUSLZAt5kU1Ek5/KG/oaQPvOIOCDFXMbCHoxcI5zXp
aJzG5D1Bt3p6t2/WQJR0LbCgD3ZBrPUKWqJlVHhV5c+oD9OWliFQ5/ZGDsLr
YjG42MyWjOsdAWNRFKgzPSoFU8wGethQYQFSzglRCoNY7vgJVTvlrqfz96cu
3zo49DoG9kezumzN/OS5RC8n3XuhgSNR9bAbSSQkbVzj0A6130eFZ9THhLAn
9EqsNfxjH+KXJJpzxI1HrJ6o8jDPkljXJfbMZqlMXG+uwiK1tYlZ11hfgBry
VfI/l67JkY5jF4WiXRZlcqPz//2BMbq/dIFzoC20zAX/ZHHx7W7P5qemijVq
nel/Y4M++5CZ86wcrPqV5XYdXoXUamTNz6Rx8ZjMV86yWqgolo4upLT9T4YH
5Hl4KqpXFaiVB3+kUN1fBNltEpfrcLReG3E/80ZZDaD0hf27xQhlE6rV+YOL
023EApKtVm6RFcNVwyHE8Z/92Ol257FsUJpu+m/auvbo8ExexfvLuRGhnTGg
UoUaC8nyOIuA41Djy7oI38/N8mBJI8BfqcLt6KYVjBJtndSVn/Y/kZqRBI3J
1tS2qLNJiy3o3XCFzuQhZNlStefVx/h9i8L7qeKoWLnS8naL1EZr8PGolt+L
4q18N24pjaPMwrskdmWhMn8BBfqBA8/+7YAurkCaBCzgm5D6bdq5ymzvUm8h
xvjmjRpWQgre26hs+PX5S93TYC3NlGLOXtjU/KkHz28TT8iHY9basKDbeR1n
+bNKXzGAeE14ApxSoxvwmBYsedmaOyFFwHP0yTrBby392QGB94/mgRgvE4uT
gKzGrAO+bSfdTi1Re2ZZ4aEQJ1UvVLFuJdGTVAekDoWO8h8RLVOqv3+yy6+J
5/kyNLYzEriIBd2Az1jQx/7c9WMf9nB8oP4YlKop62F3ApqYd4D0vASQC3BG
zbxoR70ndx/q+Q3llaEJ58k73Wp0FWeVgZwIQut5ol3BSksgxl01nfMamXbe
0M/z/NwEObwH8qqljQgd7pjpx7GwD0ZV4u/9VdlZhERudDQn6WbPkHmPPPPr
7FqVSFMWNkhSjXOpzQpsA3pxpuNRu571XrY4GcPdsiuIHgLKzHJCq7vGSAUq
CDmss6UcLFxtwFXVvlkdTypP1SGUI/WbUV9pC/zaVaOTP/oOLvOKc+f5XtST
13DUYJLvUkHD+XTYclVEH9pORreyY+JryKggpC7JT+YynlrHaqAR6tDsDR3g
TF3iNURUk6y7tinXJjEOrQvhk0q2XjaeXAAG0rI6RChv85KetequRDYAkrAZ
0pkedWEC9y17pjuHKRiWbx+myaYY1jt1qxF5VuVaCq0yiLfntDwaYVSIiq1T
EsBP9f/l7EJmo5M9NvOSIHIxQe+16SIH4O5vYqfA/TmleUNGKUAOssAqcp3j
CG34wIeTaoHHJop14uB3fd0e4LZHj1SasYq4F5uJTomvZY6F9MVf6kPds1rU
xHZPEhNdNLmJ4mLkJ8rbmh1Qh9Owf0HLI8Y5hpiRfH9V2doGzSWivlIbG+Ip
1NXfslsFN5/NAhsy+wAguu9CgDi9Hl2zIzGkl17lt64WTtFkzeyx0Wv4WWa/
7cGNFUDWOZrobBVgFF7yIc2fJb8iS80cNtGrHcpRn9kkUY6+ioJWWXyJlg65
0RXC9/xRP/A3QanW9du95qrJi/NVKLmLm4cqkHbOtFot72gTi1hgjjaYpb1h
azwXqVwqH7sHfwDcWodd1JgguGPEtF8Kp431d6xgstrurIaH32GKkUiPmdNQ
hVQXLku7UWRZXXrzf9RAy2jbpL7OreOlLyJgNas5eDJj+YHZALMhW4d7Yb/M
aL73mgsyiHciZsFAWbvJsOjpfxv0rq5BUQu3Snrjyw7WMzbWrct9Ew/TmPW/
Jm++oXP7/hZLGMEXUxtWEUQTHQQBYLvrDp+sTo5cCNaNgxcKWOheNbJIN5MN
RFkCfaxkN+B6Gsgx6qhlc2JjrND/xZiIZfzW68lAVewThY/Lqqqae54Ejw75
vZyb7GpvSo+q8IxiuR9swgfc4UVm+ANpiScIDjKzxWnLB1KVClisUqRgmnHI
rE7lP0HGMmOpnlda76nEowR6KYH1vB/Lu2/cPolmX+1YxZudLAGwkVwsF2cR
+A81BS6YCWIRlykJnmQXZtYo8E+FNKWVPQQKdKz7zOdQr4yfdOX1UpoEwUvI
E/KICcdUMA6AGw9ArCwvqsgzoj6gGowYbqEPPEcp7/or9SGGIKCfyCsfognH
hyaonns56Kg1O5bCBq7mOS0uQtTt44z1jeTjKp8f060fdagVztHhkgy+nd2V
/fkhd1s6FRD/HJE/4V9F1xurKrRMOhiqQGV+YjpJ2fkOckcaJOakqtPeoV0u
LTLCeSSYBFdKnfW4/pEcH+IZknMkZbJ5r2JxKR50UwR6TwW1yBFf9syqHeCd
jylaN2Pm4FQgjg5cjJGf2OsfbtLsz1TGBkRiyYQ4wmHJGY6L56CgXO7bPfmP
A2dvRHzzgLqaqMofxaTXYIeuu6FDYZkUvlJiDqBQwcsAKbfKxLpEhsuEj15V
pVZTZMZ2KPk188QS4l/Di+DyM+kQ2yM5utySWrj47HsQnJ03cjZspQE7W8M8
DiNLDcSliulMA3EFL9/iFI3sBZF5ZPzMErxjfol7VDzDmrPhHlnj/hB+sYLq
POLLPK6no8bFR86V8s/n0GzZGKKPKDC7zXXjRuUgLo/SgfRWJYaauAZygmlE
v+hD9E8RmNDqIN6ZAw8LZAJMvrnLPygXzE6i0s3KA6/OgU7+FubDzL2t6eAX
nM6t+2GhhRnHSKJA1IMoj5tSxkxOYAu7jnrJYU2tQa7yqSr0J4cwo6mybdDJ
xa2DW90UB9MQNs7NS0me+lEwsWjlM2dDJSbIHZXkkn4Q8rYsRuyvEzB6Qazv
q52z5bNmfvebJb2Qxqs6OATctM0mGtcj74MwX2WF9x5VdTEDmlY6zkrVuilA
5h79kAesQhrwMj9MFhEnlO+DpfVX5nuszu05Dhqd9oICDx9TAGm0kC5nFn0J
XB0t7nmperCiYYN2z1n8YCq4OPSG3licPEW952kgMAs9yqqeWhAhd/MMZj/F
R8dMolOPaOp/pZhWCjHjskkLM9Uu8jqcvXJc8XvDSRfTqh+CpbNqE8jhY7WP
fsA7dw2ObtwzCr4ZXpG4BODux3ZyaSlFd0O8GWdXd+y+jel52uUsI8XbDS/2
8UohPDS1An9MyVZj/6KsUmftjFFt5Cki7HhlbNxb4tOKM+EusttPkLJp1ZXE
isF4aJKximtn1Rpydf8dJdpZy8jzTjfMgblyhyqNPUO4cJO0EWQ3eeKQI1Xk
QOphBrvk8+sWHIiGoe+rdhsMD3twTi8BXS3iYkWsYpU9quEyYQJ6UrzD0gEp
v/km6z59LS7AQ+C6T3peowpK8eTDXmW2IxTqFKn1rUy/PlMjLS7NS9q84HRv
/Y5dWHGKVbYcS+p8YyTPcThv4gi6x8b++4asgGYQ82dn+N7s+5yZvhIKcxel
hrtBmhYKnOHzhUsIl4AMtMQtSDeJZ2nKtlnUVEcQ1EGp+9QLer3srckr9BOf
a/jBWi8JLUiEyoeA/Z/Kp1FWKVSydAzgQ+tSWIoI33EymGe+KfAY/CPbtx6B
0zdXP4xk7uG4uoASZ6FaVCO6zlctADmK2bxn9DyCkc77bpoocS6jJRxHtOyy
bJqdZBxUaYcBG+ng8JdiNCSBPfDh0mPoXnwuGxGYcRFFigh0XKcyAUxBYIqR
ieJcwhDUjsZICHT8geGNVzqOgnHMvF62jw1njP33bxd85bhYkcTruaoAijPK
2Z49Soa6VqrpR+znTbI6RMb/mOZwxkCJwEWKFhXUVUKu0G7KCvdCJ8ccD8nb
Lo5ndkAFaBE5wejlkz5D4Ia4gQupteCmav/FG6UI/u4WnQens5cta6ymqPT2
W3ZDh1qmSNnF92t4/JIH8cjwE7y6SADDRW7Pu7XDBRWLLBR7TibprLWixxnF
vqca/2aHHLAvjIJn2jJkDR+wDV21p2zLkth6yt/f1XiKMx3uQEE9QTLRaESW
s+IFpu9EPssMqPMsCzaOUSU7vX7Obt2sdY9eHeDHfWNeKJ6XwAu8Iml0LHEG
UhTbfvH6yb/p+XNQHFD7oCF6FpRbh7rpnPDs3HZZjP/8UronNjQrER0gmcua
9VERQZ7cNxBV4JyE3PmM+nOTJ8yLMZf8Ph623Qwg+Qa+G+eyjy7hidKWSlZ0
YUMdKDChTCIqJkY+Fx1EV6NaH+enEWgcujUxTBpY4hoO+PDgWop68gWUUHjs
jPi5LMT2mvvS7DvV+GjlI48NGcRECElzxOxrqu4JJmFnTNoSqYRspVXwHLWn
i1P1+I7Vf1lAAvzbw20FZb8ZdAQLQIfYOR5EY+JCbZCPBYfp4tNIsmeWEkHD
lKw7PToGPAZcJKEAxUjVw0za9fJbda4P4Aox6xVWLaiZ+PLdwfJ4j6Te5CXQ
ujTGBmlHtWBzc4wH0P5mapv6fdyvhp+4EzS+Zz5wWmkSaqOXWiWf639+gTxK
NIgF+GtM7s02VVoTap6ZEug16M0C/GUVeOX4V+bU0iZui0jKi7RR/7oEI00W
ieJNElFHR8aIRxEPpWvaUpS28wny+Kwi51IfdDjQJZEQdTodN1CVpfmPsW1Q
DoTq6Uwg93ZFfUsePg3lPsu90two253TBLYOKmC1PZdXz6oC52u7/BCargjH
BogQb0KGb+IKkC/wJVu9gout0OPyMaIlWIYrB4AymS1KbjEpkM4HzSLhgnoJ
T58+wulpWLWDSCni005fRIxQwRxpRTYeHbcp6d/h8DvwQOKyOvvU+2600rk6
fxUKs6o3e2Pgurlx6Jfex335RNbqM780lp6djVhs2D3p4oCfKL7BReJg0NOy
pEEjNHRpjs6hZ5X6sUFebtoUMwzHl677NxR775AOeuUISO058oSZlTs9zFSj
xW0nLOG3AS7iXVP3VHyCjGnDYYl6uAwQ2DX5aRHPHf99FBP8un69cTmcj0B2
CXNdE/5qKAQBmz2Eb8DUPtgSV9m4uuhttJW6ceKi2zxGCGMgt/uxDxlzZTAj
KxZN4dTPNMMxvv6mZWaRhoI1PW9Y4h9n9r0/Pm7xIWjcd8a4T3lCdx5RhyzN
ATf4zUd7Zmnef5dIFsH2Y2XTyYI/fXh7KiwLDA7CJA73u/jDE4V3aMyA7xS8
pbjkBnk1NqxhCfemYqs5IgXQmKT2etEapeeCqo7mkIXoG+fzLM4ZX0Y+EQTn
N6LjTkKuWcwE2Lr0C77Voqov5I27pJorWIv9iPvkcpV7hPkAMtPDD1fnmEH2
sHsafZDp02it8c41/WWp6mla9b0txyPXh2hvct4mBjwDqoRsviOctOinO8jI
jQY87cyWkEzcle6wsy4ohCG9QYgVtsnxEkYc1rkvnlgpQs9f7lc2TOr1mHZl
pDWeozmK5gYdYsLVB61C7+gHr67wVck8u3ttZkPrvbBKduxBru1adssi8Gc6
XNEF3wv9eV/rfJ0wE5c6TcqUJk651wM5kXGaSgJGzC955f4SixzxTVqvqv46
r6cef6j2MsIBxpbBP2GHmDBIs5fX0+h5M29tW7iFMdrg6JK0ZCYoC1B6yxHQ
qQolLSEXim1TSXDtvgCCJmzPr68UTs50bYm27wDXKGyjXOjtophZlkEfsN/z
olsAjezgnceYVdZAMmExjUjymlJwBAsvEo6rWg2E9mVzGtV9RDbJS2aB1mRt
SfQJVnrA9mbiBwxgkPdIfD80jn81w+OAc4SqG5N5MEamLubY63cQNLG06y4d
cY3c4Tuu5dUQfx4tRRCXIB7Qh16fZV99CX/EFQV1TRovTZr/E8OfNsjz6/Rf
8sVRbFR4t8jswuPqkStiEYy8el0O/BYPh36J3+oIfx2pO7rX3smHok6HD6jF
PNBLtvu+mWYWEoG/fXKxC40L1FLPSu9LzBHQe/gDcRmw1cvY8XCLBB500Muw
Tuo1LrssdCJg33/B2GhgUcf7qN4yKI9Z/2hOOYuwVrMe9gorMemk7k1IUFAg
+Dem27NjhqEBsNzLNeaSS+QwuggKyOzfXrFc6e90DG7P8uKD+MCpneCD2SIN
S929+jdCXlWzxRChkZj9Xgqx8u5OJXZM6ClDipnzHnLoGoWi1NGHaioRro48
bITa/MLpxQMb/K4YsmodcXwZaP/q9nBXs3JoWERpmvh+mo/hG7kr9kCWDW+F
X9baMCYPtA1L6kpaTK0EiI6uVDOApkoN5nbYKLslcW5VqO4W+6MER09WkXBk
wG6onp06FzQ/av0YzjXPiBfTTfl/Y2NCHrWnKWOKqRL9+pvPWCTr5j0fIfSY
f/FXqq+o6ztF0ZDmp2ojoo6UgbdBmBjhZicjWlbQ45VV8EIj/VMu3fdjEWTF
IyjoIG6WI41ABVMrVDKLNRjaKbUNB4dzmyh5ZFOtKWzlQdv7ElEs6Pjm7Qbk
J2T7sUtcYejjsUiiLxgMCpV0z3elp62nr7wTyTwnP/Zsa993q0GRhKc3+fYV
sVHGhQHaPpmaXGWtsCufUCVqQsK5xpxA92FqtUAYRKGAvJXGvaDMbeyO3rKP
HHFXbyGsvoB7qI9a06MJ+JYopgLCFHEve8/Tj3lrdG4aivSzcUHui2XHYuci
Z2PzD5Wq6posL3nzyziSbWWSK8o+Z2gbh99EcrW8sGW6JUZ5BW1uT6rbUlmY
W3W9tKnqhHJcNT9zTO8cASLBB35QGqGbUGwb351grGBRLFkoylAb7ov20kzu
jY4s+/Dz2/DFgiPZXTl88Dx5WO88Iro0n+pZQuymYueNYnZI9b5C3CV7C3+b
D40VuKlC3lXAEH1llrz1Wq+aZ7SyuWoxbsQF6Mdb7MEi6Uj11DPGVvaPOZpN
G1M/Foc88oVfuEg6aTl/Z6VCXl7VHKt1Ya9Wt/H5DcMIoFCYksqunl/5K59S
pOQmY6eKXmYNjaBg0XTEgv+o9FsGTQn7tYIrW3Y7TE/YL/NHzufl2SmSubCT
0d9n2bb6cWLSjyIDvK1SBHZeOIT5OQrrFTlVLUw6zC8zSqDtBarHLULl6+5j
Y60hzwKjtvsbV6RN/zXbTnV9jflYwVlhKhLU9RvUNXZn/coIphKt0mvXS9lw
8D66k2zqXbErt9Q3HdbgG6TY/Go7DZ9DT9ClB8U9ixruwLs19+bkVh9MMEAR
QY0UOJBN3t6bqvKSHFAQZ0gwGsUAzdcgRh319HpfJ9fsNt5O1BzlWjtxT9Sh
2/KdN6z2LghqiWKd/iKQ0m9ktReTI/sTWD93SsQ/koxpsRkAgG4sagjhzGsi
PhiYYfhN++xbjCSopUJtUCMCRxuYO7jXREmFZOn8iCF660Nx3rf1+pjFkABz
ezw2HmEmkZu+KCnSpY5N31aXiqSLtMIgyoLRD9i9QcjJhDK9Pljetk61sx6L
lEydFAa0XCwqWkVgtHvjOBIq3V3NtBL3IgRYppASrABLkNuv4+4bsNFxdW8k
mC0voc9F9zqx020h7YSWTmGPLhFzW6fzZz5cqBEuz2G9h7Yze140iMOCQ8En
vzoQDGzIdOBAdeITW9A3K/PSAUWrbBB6+vlVrFh8+qpQgtzpRstbi2++1rw+
MbQ5cgObR0sh2UGxXuT/iA/pZLRJuX4eX68nMSL5QWh9tdbKmR2ZCoHG3WS1
/DaBZmiha9sD9Q9i51kZ6LbpylgKzVgqiQJlk15+n6jbRI13Dqrgthaf7AD8
40JR6cLbK5Sq3qHnMDt6NbhIbeAYnTGeUyfbjWxeAEeT2jhWR52/10z7/wKQ
G0iNhceoPZrB9wno2vVLnS4jv/HhoVhOj0enIldSyv1LqXK2+n/qPXGM37ZQ
UNpEGTosc3Hq6WrJiqS8lKGZLk+R+3sPHXYmgLkTqa+G/DzRt3/PRhBbsxkk
Svvu5Yalnr8o6c9nT3RtfZi1LWE/0bi+UL68jV0+J0VcP0stqg9jDugHYPt3
hVk5+ZaQLOBEfzsmJ5akQrt5uyPC9tUEO02RZKQMkLpBqrjuKl0z229FjAZ2
lYPsMTr9ZgjzMe04ZqQRB2Kk1FfObxaptw1soeOQmoz+PRrC8cPC8HHrzw4x
aMNYZfsw9elU6zCdTDl5X00R49vqcHG9PkU1NFw3DT6HxO0pIspaZuD8+8Ju
rwr8rTdg4/UcPjpJyg+igl5paK3mAsNgrYeYMlxAiVZ/7B3BDMxLgCBLAb3N
mTApYMni6vL9t2esPNQCAl1JXwdg/jPLw9fv1fJOxCc77s3PXD+z290W+wDb
dMzB6F/cDw/OnfAmwaAszk/pY5IrlIyVmojZRN/bSXfuK0+HLV0RRqO9Fd7r
d+Eh5XuF9HMSmJokrdxPoeSwl46hFThq8rbAM7oohgzHvbxN7pEVd7aD3aUv
deT4zL7dCOCDQjKq3fps2Z6Lh6RCkCB0L4wwNaHIo+yixsNW4sqgW8o6yRA6
HphX9KKae+CdhE+P1MW9k1SwQqpcdA0boaybvE6Yi40delqJuK9ZKCTajVTu
cNAOh98LEzGVYqKgycHq5atw1t7ha9kFuo54ExIZ4rKWCpgR4RvlXZtemCSe
aH22f720QU5I2WEPfv77DdU0S7aXrYcFucW2NR4D5TrsyU6vJN/bTOLs8Qer
+UJ8JRdIS7cuJ6PDbxu/Xo0Y/QIjn4oP6ATUkdQYSI+f1e/AMmnxOoUyzTWc
ubrd6DkHmtuac2R+/AF89DEOt8EWR9gvyFhuQ/5wfVXvcl0jmVtlVURvLUma
u+GNhXrKm+uJgKRL2sLB35JfQMlR5fz+xiF/gJa2usiwrnE8tvTdOQDEd2t6
I8EwPpzJ+7XQNAEbaVLKcBJGnAZqx1By81cEbkutkrjO6PQQXHcF3sVi50vm
z7I1uhPL72DyTRKD4xSd9Gx9tknPo0wPd38Zc/aXSEdM2JdQokjnV+EMfdTh
1dDhheF2XptE+hKpUOpzWDZ2lZIMVeMGtjUekWUnRRZrJqCU0kTuaoy2mU/v
kI102dgQEKP19RD04WmeLgtKdtT+2jF5X5vJTtnY7pKmr8wHVKVV7hC3xbxV
6eUI7V0TZZuWC8p5K46lt5z0QSdMitONHOt0rGoXfVmDhDoWH4Pz3TvKc/ou
KaDYj37Eh73fgOF5s48meIU9gSjI0m5gj+JbHapddjNkT7SYjKIKwmDcAEHd
5hxKZ6+0wVKbNYdtD6Wp/aIQj7iCcDnysQdGHy9eNIawqGzmQ4ybZNCJ7cN1
+5pHqFY9+PXRFahXmq7HfZKGG8bEDPcrmBB08UY8HLclq2Dti9iYr+ENK+gZ
oX84Jyx1aKQQNlsDNjp/JlutYnWO+mW9dBFKRUc4emHnu3Uu6UxAm3plIsVi
5ZsLsVRnYFpB/Jowb96Tq5ir3NG+W3ep+Kl9k6DC3sqa0JL2a2d9l5ZxRqPx
X5HfKgq75IhToAU6DnePDoSmubKCIR1hepciJsa/XX6xUcvBWDTaDqeJrNSr
ihaReKhJRxyi6sprlHnRTcwrz2TWlScHVvr6JdvCDTXRuZmRTwdrC1iQWqGL
stUF5vl3YEWA6nn/I8T3Pk1IwKt9aolOaiLYqYZSHySIRH2bLLjcUZM9LCJ3
IeeNav/ZmQlvIM+y1B0PVxNqYO5iyjFByzbhSjECOnks/fGIcSA9voD7gbP3
d+CQuAAfW36SjKrEqfMsTPIXKXkOybFLOCbvS8odlKEIk88ogKknr09u6IMq
6Lg7Taw5l5I1BrJoOF7r9nVKa9AsSC4MG+c49nIWXaFtNyLDvOEs1XNXgzyf
vKNpzG54QZD9RyllCfaIn9A8HFyG7K7vWzwCWsx9+FaMVLuh0yur6u2clckH
DXHLPyZowvI4YRjo+gpPGEFGwbmH9UIaxp5mYnfHKcwLkvCixgF7GI9hjDWW
cJrR8DCq/sucwCRw77Q/sDtunLXJzGOkxLI5VEzxt/UGFor3TjEHuE/BDRuM
OdRNsYMByVfTzpWsjEBvAs3omcssxZSlD+Ag4FgAizMlsq7kA/qTrSTTW4M4
+jOl3STgKoGe5YaOdGbm6XCUUtCZ0iZ3V2UKX8CrgQ8U2Gu9DHkTgFQN9iHj
khBIpeqZmVWomvo7PkBYkMHZbL432CZMr9D+Utxd/qUHuKGZdZB3aS0coBJT
AhtEw0x6rVWkkJYI1vjqVx12jir8UubMrVjU2zW5KuxnCU9DGtYlho5frjlN
ge8Sf8+aaynF5nlIlEX+hpzvfdPZhllgIJlxB4s9jNx4qs6yfdLb/cjQ8llW
egFmD4Zxz1gT9BuOZXAbKnaRfuOf1chGG+WRvM3wvQJBbuBtJ3TwAG+WCX6U
wZ0bdVLLuhm38lO1dj33MlsjjEpudbjgyWrOYkxatyKlwVHdhvMbbrqKmrrp
2W4KF581Voz2WB54clF8SsI2G6GbiOtuuy6dUt+uo+eFn/mphDkYkgoyU5ni
BI8X2LKxQJZs4DLfe2rccURFwSAdPseGN2VcS/tIIptJPMC7SA3o+w62Mpsq
IjIxr6SikwP+NGQWvOgjPXwEP+JS4S/91ngH70uzCBdGSv4/rkkQBINzt/XZ
pnzKZh9ZM5BWCXxVFSuvDd5WrYuA263APNI6SVxUxVpKjuKvvY/irDxyk898
jYgsuyIg+Gs7Nouuuim1qzxwQTtMAMAqz3sVDCn6MLgVjNVhlx+95lRH9gCk
vXRCuXMpOA0Oq7umcDcv4E/gXePDKBmxg0NbRacjg96tBEiNzEtMtCx89qVC
6GV1pBiIm+xiBpeQcf9alOjXN8DNIsa/jVhuS4hq5WJtC/GnULYFb3BDn0ML
7hGdLd8U3KrvoERcJ7h2O/yNQ5ZZIMYWJJOo5m4e7ubH9yn+kGWjnGb03/BM
fdw8rQydz3xE6QIpW/omgNesYQdMWdx8BKkwHsQculhhi4vxvOp7Z884nuXg
aBeN4WzYuMV+eRIVu8SuchMJh0tqdpY28YazUZ0XoNBiqxLAA9YrtzcQaJgV
KU0Zfk2JjSl+XMgOr/Z0/J5Wg6O9aCyYfmwbZWWmTEw4DTyp9TefPjQAeDl/
pnH/uF5yX0OUERkLIX8HB52em2nOHqTEN48hLM3dswio8Pq0Rt28B4cNr8El
RjkDSr5A8e7mKOH5txWvT6Q5Tgisf3hO6gEQAQyhuuKf8C+bW/L2Av3s17G+
CiWbNjfT1/TooakPQq3prgAioA/BCx4MB55Ios01/83QJZHTN0R4IgbSHH9T
z3JvSIlI/dKTj6MHSsvSXDPGhPGxCXd/xpmLTLh98HadfglQNms6ypyMhkBD
Bbzj9+ihM/jBMsB/MVyCCkimVQNTg/F2B42cS95A0T0Hz83KxKbocuSCsb65
zl3Tt0diM08NAPMJOJf7mW4CLysLRXImtiYLkjS0EhxSX9u5OETMNV9qnLmi
abt/vCaUEEk9GjMC4jtObawzM3erndGArh0rwEJtoaXqNX7uZe1009/wcSBU
udcqsj8sdY8TU4/C5YPb+67OTIZbFfdyCKHk0lI7JSV/8so65eNxLctrpVpd
Bc2XAGOiKySjNY9QPdCnp+lJMM9vLHVFpEeTAhyNRppvKFCVq5phTcJ08aF2
9keEYyV9Nj0RdA+SAUO47hiZMK88tR6V+Y1hgs5rcI2xFAUviDRAck4QBoqd
SBaVGa63OGE/awvTJP8OXpd+J2igdKzC1AsBmcpt66l4VHrgOjC3ED0ejjud
IuhypNIbx5r2JpGKvvZh6HKMhuBgCOSgzsl9vTvW8PX2YVfZxoCUqOsVpAe9
LVDhztubKF3IAHzhgLB3z3dg51fBv/9u7Almm5PhBuLywqzJ8+uldi/sbdoN
3zkdMrZpKh29moEuwKCLaXqs2IuIztfFi6Rf/qwVGS75co/UJz9/eX6FfVMv
zS+Kky+6rm6vBDokHe4nVf7Pr2IApc7qwOtbb9GKGXtpGpLRkUDEqPl6Lv4M
3L1VBrGFuBy/gBCBAuUcqviOFdmHsWvM7rddSsHdR/jLvppcK7HjthJbbYSu
5RbvJQ6suKwmtpF4lnzK9lvOWISQeAjMkSsv4RgBAxb/L7sK2CRjm4QVTVFV
EWqXnRu/aTGuGt7uJBeml8Kr51gMxiFdgB05VwVCC4i/Dnmo+qgnx5bQAP8U
UKS8OC/l10VdznTDUjrajtTX++yz0bVl9D6BxQLm4HLVkD6syZqNwi7zT1+/
CtUHMOyKDN0GJ3ncLpu5bv51JYgBa278vbCpT/fAsahgr9hF+EhQYu5aK5xL
zhvX7qLhCj0ETNvC3T2ZM1vVm/4DJAUS5mDCkGmjlJ4O0TaajEXjnGcebjXZ
OmfRN3Tp/BxRXEbNBi/+Gk+bC5aWdDTfYpAkoI0LPs3SDY2JZFqp/C3BedN0
AB5/itrfQQmr+IqXF3Y7pExmEg6mF7yXQNIVb3/5IhR9CwMScCwpiVI8NxVx
FwEdyNiug+CFSpAyMjVS8PvJ3+K6EC6h9euEFVO/L8cAZzE/M8RRhp0oEW8R
P3cqnNWHh0yeQiPM6t2cJsPSLSdiEYK8LTrsrIPsu153P3yasj3rXrPX1ULM
p0LyTcBbz+wnGTA3N/6Meon902X1MbAR56kBGlRr+F37IbOmcFld8V5ws6GR
duv4FPmEWjZCQgLt0zEXQWwKuJmc6Lf5xPNQMsClcSYc1KClVXuasDWX/iTY
Onxc9kC0jmXVfA//Alrx2P56gloH1ftQbP4f8vRKt/sYT5dJ+DLhNZGSnYxH
FLG5zJvUvFo2hcq5VHTz2yc+pdvFGVhVTOLTVpUGh3QJe0q+ylqrlVoBOS1F
LqD+5k02hrrFZc4ckYqzj8bNsVQsqG/rgQEAstl62dlpbZAAuCE87M6Rn1Ci
n34uujOfZMRF6wHSi0B4LaUoF6VgYFMHyfE5SknXqOskZs1430V5oTnLn3dR
jKp9rh/pDPhvMaIolmJuyXInScmdpWwwr7OQ7R1x5lLKEze/EO/D37JAUxlO
QkC+ywIenqbUe34Oi6Jub6Dt9rsvBUpLUweEFiDRKLIXRHOqaBiOKsa6vFgC
ULyqLiXIEZmKbL/+dGtUTU0xwyKLX6pq8eHrA/bH0AldrUTOngzKMmcXQxfL
FwM19T6DYZ8wqq98vxDPPintpzi9ptRWi5bQv7zH2FvsFEwgIPNKbVD4r92a
Y6AOG6iavrqLuo2ZgZxF8L5gX4My8fFHS0xfVJwmGf2JcMqQa1wZi1HPVDwF
hZG1/0yIzcFCfIwuEcReWWV6Bq32HF13OCDE56Z5ogYVlCrER1Ve6aBqavsG
cd+jtIm7RtQKpop2IF/MqgHa4zI57n0UCcQrOiXHT+k+hhZC6gBwZqA1qJPM
kD4ukN4etJJIPTVhno6BgkRHMbTFlC7DetLTPGrPHztM27+MZFPQjEtZhhMp
QoSkO5/nk3qUosAVOHdW8uhQTCDzZSIq5+ayddadch90u4aisuEn7v4nxCb0
HtNIBDHhEzg3rAkGIg6OvbRqKkFhRZQCS95QPBXm4Di82kRrPUyoc9Qkz+/x
yJVcGbyfIpPtUKGnCZNfIyZnSPyepqjEkbNYlLY6T886/hlbx3tSPSPBphyn
cgn68iKBq0vWvHQUnFWuoQ6+itJvXsEWxpjagw5NpX97K7VDeMzOixlFgjfS
Z4q5EqUO4eQ/aV2sjQH6pn7lLA5ECoHzT0c+B/rAju1du/Oc0UiROfpRs9zG
hg5a42j5pNZp08o9h+4OXuIqbRJOkOi5m33018HHksWkBLczsgVURGRqtrO9
t1RZp3eAnM6VORO9j21UInIfA/xADfzXNVR57KnaaSxhpdV3AMvZ5Ole0zz6
tt4tGqVWa8hGoqLbOFjiS+ZoY0A4oMtXRwQjrV4lDyWy9RzRHeuZJxjuGcoO
bVoyTAAFvM1fJls9130/5MF3HGhQNb9AM+velZY4AKypCsR3JzsbDb2IVKBL
BGphNgej24sT/09lXTdNtrGRTOemuNSoFRnBEuAUYTgFEuLca+qg1u4xilAb
kOQDKsXlndL2sk4/qYqUVmo+XxgxTe4ZP6MAUrbFahApsW8rKyXNkXCxNmYx
OsQWricWohmocgpEw8mIvbJ0LY6Ei0gKj9EdEAVjogO6lcKdzxdpe+J8x2b8
KL80wQTMZPGJWC4S0ruUrWU8PcmPgHIClLkA7a878m6/e3aWYbmyc1+ouo2t
B/zHUjTAJdRdTwQjZyF96yKxbJxHxjBICVUmhkaENuSx0yKE0vBDIWq+0/uI
YdQ8FhgU7UroWjlnlkF0EBpKzMhygnoiFcbPmFoBGFSjuklm3/I24m2DCinx
8M0p3OkXIMaD2S5PqTAEmy/PjzRGkwscMpOJVLfybhF4amMUBlQ1nwfz1JwC
GyPW3eHbrM2Rfh0DH0TsyZNVyUXVxNingdd5ShWdRBF4IUhUrI+uJNCt4wRE
dP0SBWvy2/zAWEMuL0trz/VlBKyBcmWy63bReEPjqb6xuo3+6VJIqw5927sC
z8feJ0GUkqb6vZe7nfISBggGeQj2sNoemGp1Sx0izVAOAk6BVdY3H+DReciq
ES19Ax6jjqwQn88eikOhF0FOUEuD6lLh2OX0sGskEcG7EK7+ESMjc9/smyYc
YikQVoKvHEpUnaEMXQ7vaaN8JRhHwPwWTDRHi9CpCD2Ktv8YMf55fDOaupNZ
P6dePJyakdyb3i2mXG9NxK8edvz1NegkX+78INXalO1dlDqClQzV8V2iUyO8
Xd/qdOA6t0gFA4ZMzXv+gd6Mu3J5uDpk1WG+RMCHXGQc9557tH6eFf2DssdX
3aRGvY0J1CEtrnuCSK1H/pHAMmaof7/h2Hu9VtlXlK3O+oFxmVMnEm+gyuWz
+yZKgr0O7NaqJj3SnbdfbXaFbkxspyrU49NjPNcgJNS44hyiShA+pxPFCbDn
DmWpkcHGUCjxvT/TPvIEOiE7SLM/mipXVql1aMVCTXPaD8k9h8oNAZFkrxhr
cl9tLnNqiNBqmFmK0CbHzZyLFW6GeF5xtde+f/ubEMHB8pXnw5OVucF2kHyj
epIO3o3kTXEOd+PWEd1pm2YAAuXoAnXPrjDOuHcpErOdLo7ZdLiil/3iucqA
LrBECkGhJle97S37WCWHM94iY0Qsqy5bs6D1EHjeVzW5ux+vfunKSqij6tZG
lnmp/ks3het+M8LZwAEYjdt3SyNmRW5F6aYsVb/2mrvf+xi6FoSWikU/EcoN
qXSsiYwmBRxUS8ZfsjXcpvRBXbPTpttvxXjgOl8zBHpWbM5NVuZIpdsNfykW
LFbsJg/L4Ync5N5djr5/Y+rgpxUAz+yvPcmgaZAl0vEbd91m0S4SOWXzcacL
fDcNczhDAqE6GdeqCn4zYLBe3cKtgeJs5YTksGmVDJ9ZShHAWEgSW9vyMJpG
TToavrXbUSCidkEfJCl8S4utaTd26dSs7LwBQhtIVKhoFixSEgif99Jrrs/n
dh3htpGp3wPrvZjqRNn80GeXdkyaSc1Np83r0DVcc05pvRBGgNdKQo7Dxe2z
FWxFPIYHIDrdRkeTaTmydWZYToDu5ahvh5YqDjtTefwfvCggyT+t8RGXAZcC
aEisGSALtGYBFZj/0zSTQml9lUwcbp0AaqSbCwp2Obu9NvuNQGfL0SFIKax2
fGTbyCxCJufKANx7BIktRIeJDc5IzHWt9pDQiYfDjHodcKczUy3rYPEFdrPD
NrrNrtINKlWzhaLbXhONCFWoDtXTw3Lghp1Fv+nDf7AH2mZvUdqZOqoerbdE
5fUd4A/17ZwLPp6z1rddFEy6qiVmDhpzac+ms9d46WuqbVMVh2poIl9yJQ11
/KOk7xTo87gPHVaobXxYzraqvJDuQ+56zCAi4IL9KKMMLcoMD2vo89uxTUEL
J7AlF3SbaXnHky9DChx39sS+eKbUFqphUSqw2E5ov2rQ8ipLXTmKiQqEhoSR
/lO6yEBVdDJxEPKKfoEGveRiciqKsgH//UcUmXIYKbLFNyyagCBAEG0lWSNn
rCZuwtJCpExtDSX0Mr96g0IkvKkHyrzmWu1Wxqi5Vxm2zZzzvo0hJbsG8wge
euv2l3Z4BfWs6+jT512GLVUhIMnr32pgEk1sOTevEEImD5f89i9+01A58tvk
lLzLjfHW9P7he9ZtD3m8hUzBVFSemUu8hkGeDQkiD7sydClmclR+Fq90S5fS
ZPFFz7LO/AXiVLmk/mAbHLMfXbV8VJqte2yJWZF8YNH8dEU5qzmdj9sVqePG
HeSCaPp3tyiyp2GAEFiBb0zt8oHvIMY3DN/S7zfZ9It9H4GdvwPvXDX3VysJ
WfNQR9UCvgOFenBH33XtLsFlHMMmQg1SiOGIxnkf9v0tDur2R3WV3FqiA3Zj
RJwcMlxB6Rp4G8h0vg3dhqEr87aeVVNCh7tPqqBkEDZF18WKmSa9KvXOeYh4
WcisAnP9PPVl7f3OY1cDFaDqL2iTwlH8+/rgajjGIjvjjV++x2pny4vUmT7D
dWVM5X1C153qwfpKMp4jlzvjujQn1I2nB0Ent0/HULJ6vM+sNoKc7qlrWZMT
zEjShyqL4F1q678santviIYCQtO+0oc4b0q4v6wqf+6eEiSeKy14q5sw2XRT
aCMFlaEILqRN8JzXLBxuWnyM0K0IR7U21SPk/7Mb4960SUNEqrE1eRToOASx
hOJQ+3eDJMGW0nX8C9e6iKy0ofVW3tT084sXhzPVE3EHhznQpRYJEGTRRKem
OIaV18zU/AFLGQKtEZiyOGIU+ipMWK2VqwBtgj3E/aXMLZHty0knvd/BZC/r
w6pKVgXuFLxY+bb49KcPE71Po1a+noUFpe43bivZhRik9n/ppo1zMJ0OPYS8
rrW+Sbzitc4MExpnkAmp4vTp840idIPo6CjSgMhj9YiX/BsWW0gB9/ez2KXl
OcM4d/03YkXAyIbnfaokbbPv3ZUejZCodsBqT51LT2RAtdaoChI/yE2rCdaS
X7lhNgQ5qQOTO7JCGMvDSinC/JvEC6v4ADBQO2TIb0RdpoqPuD/vaUTdKosu
jtLZaFcRJ7udRc/gaL9lEIJZzCeP/Pv4bd+BytdH7URyv5g5lPgKlOhtCpIU
jhlU3te2J0LbpX04+yqf8MpSg08tmZddyWcq0GaMCVn03vtJ9HFriPwcLyTT
4sPXPPLP859m/Nq1R8tgXgYBaE1fHStB6VQyv0g3r1T4U0t7RPBge8w+qZTF
6KE90q+eaXq7YvWtZcWMU3PqHGQWvVTdoVL4MJrjtUXs0/dxU0KtqkpDTVGx
VdGjAey+GXCcvqVbRnlweeLmfnCst82vru3PCZlnY3ZiZ8eMZQSqLWgCxngp
q+Hyt9iOaxsNJUIBYXyd6U2hv0o7q0JHI+t6ghbhHdZfhpumx7iKP2dgHupg
RBwzOug8NFtYe6Np+cGmImltoP0mFODedwuspj296Cegm2SCMK80VP56JtgH
2NvlJoDuzdsHuE3ig1PnQ3P7Zyzj0mYT4lJ0Sj8Oj6612ylpBFWIikHuvXI6
Oln0LKNz4kWH4YBvBDnUSAaLt5bLT8t4ZM71AYEkkvJfPTJPN7PXpr1wNXd8
mp6XQNMurJJ9JIu0gOLRTidOuqauJsdGxmeMvQQowRJI1PrNOPg0/qwT/dMN
pIX9uaA5sCUL27vxnKVmzJKjWhuoBT84Y1TMOF9mI6g5XOQUtfqLkTsmU37y
5ZNF9i0KVrfeM25mA1odMlfuAJWOnr3TqI5818FmNmg5t2K0ervFbklJdU5v
JA5KzIJCGPkVi2HUTC5tV0OS4UwH8wZNNRJpZ19Yx3gilDaChGxfl05WtfwG
zlehC9qL1exDvVdNOYJkuOr/g4rbIxe9S/2SG/b5pBS605wm+jaGyVHGL4mi
WWTVjquACnPQ394LMkGFhLtTNI2xEV42Gck3icL75bZdcolXeg9iMX4BS/U7
D8oInObogY8Zli73oc2MMWaVKO1ZEadiumEWuvMku68RCga6IexaEtYs0Auy
3wIHwPWyzJu1Myyx4h2W/QCHmxHi7fuY6W202haaUTXhdDSx0ggTTX3gK9Bl
MKTAQkSjzoosCKeNcI2N5plu51ACoRhvQVCAEUmk003RgBqZZa+b3/FHovht
9lq5VOigrrargL22Cze78kZ4+lY3Jjj9pP4ufXhBtdhMoUIhiXqGHU10yHTR
404AqXNW71vD4rUKkkBb5vwlXaTjR57nC7IELlhtnQtqlWZ1tajYUcJQwNSh
nGL/aG5oJVtSebLSbn5qwaEkCh93F66HEU1jsWf/QO9SLD3WSkOQlQW/1QLN
WxONqcot+lTHP+4wnq5GYq4wem0Jm5fI9cSM+l91TyufhDN9e3KWx2AijKpw
l45WoG5dhq13gSASMpQVI/6o0ZgmvoxngoTDZU525hOz2R9so3l7RWOqTcp0
ZJ6RkKVFeulGAu894TcoS+UioBVapaAYANtDr9oHLr2GEWB6MuLzckKnZ+RB
MyfYf3Sa18ZwEScDjYd6510izuB3jpln/shxXASJpobmVyBWSNKOAa7yNYqO
sjr8wCTuCmyZghbNph4qyQNqVNPdTNV1RDfM2pqhfr5zRQgMelM3w+Vl1ri/
HGvT/mZlmGO0LQs+XVdFYBfrXxE7OXbPuL30UMTTaL7Du3tMcI1ash9FLXGB
HkDBcC3zLaK7JtJRl081TEN32G0Gh1x3mRODNW5W2LzPtCLTf6UKRPJo4YYR
WmFAaNdo7zhDxtqi+Mvef1hL090umMEWLOy1N57NUQza6/V2qDRxI9SnYL7X
7D7eUQaIDpN9Ckh0Cae/ZWiM25+En7t81TkJp53DbxbyPiTQZZYAnjJAVEaz
E+deeS2LL8czWi+RhHN/sLRKF1nN66j57JwnBM/a8831ecylXire5E30x6pQ
/5oPQpn9tEJVxs3K25i1Fsw3OdlKd2L3lWyQZnSicmsV+mv9Kqb8D447nRN6
zRW/Rhbkf/p9IselQkoyNieBVqPvbZQ/sIFGRK1YMevTaCORVydaKEv3QkT2
QpW3CE8l/2jt8hSoLZ7tBQnZ7ITN1ynwsOninyhSilnzJ1qF/0mrftq3YVqM
MOm7VzRWdjHvK4Z8p2OeDjZDwVP572lwvbP5XR1qNSJ7q8eZAcbj6T9U3QNE
fchEXwZJWG1k9eAsP8Ru9xSj6p4oFemZjr8hiw+3YMmsn/ANY8xxhIA7qBTf
dvv/37gj1xbEyscRJ5rH1zt2SXQ4mBdyMmYykLoLwyW6Y5srrLRvRTbHBgeO
qi3/S4KwDcEA1OF2wZB7ne8eILsSwyVp3Jmc8+dr2Qf6B6+qPga3415yfp39
OyKociv30WZZJbRNh7Xg1xml7U9llrXelEVUSx1ilV52W8TQFdovN86s9VY1
FslEkV0SD7mq57vFPT/v1KPG0dnts93e82quW9oUC6iZakS1C0MrmLwWBpxI
+Ta+F8u6MuF45TKUJpCpUI/HfCce/bh0Y0nHNjsefxIFXhwO++DP43tkQS66
Zt0PcRBjfv5AuiLHzkSbhx97f+xod/rlIYdlY49j84RVhQFdq0UDGUwlemHs
Umn1f2mwCIxnCL3hkd5dn3cRS767sbI8mMXA7Ktb97HvHxfgCK9UHXnn+fcC
PhgyMiilr3JdJDkAgFz6MudAZDiUY/JstzEsOUsPxw/9Bb4edQW0B+02PVPf
57XVLZ2UaR9j/d2Qf54sz2CHBXsr/OIeZ7wmomNCxW77BD1caCagDaFxxMSb
FbGChxUmFpLf97S4JfTQM86YffDcFquvz8oH5EIywl+8y6Am7h5WWpQuV0Qd
gnna1GGWLpF7wXPDIvtNXbstkYqK9NPu++5OBbjvtyREleek1KW1PvdGwiYZ
lFIx4yiNRB+4fjEOXjbqQ9iVvTFAr1EG7oYdLvNMuVbuauzQXpphlwmrX5Cr
7juo91uh9tH/DkDq2CMDzQlPow+o9zd2MwzAKYXmPnUMmJ3EqqqKkAn3K+yX
Yp0N2+xGkHmuvB2Gh/JZS/0LSQW7vMdMy++vHbA4VFnGIuhtvsJX861zGTB8
tDUg2xsi3EhSlxLGl4UVFCVnfjVk+k8bBXF7HyEqeTDMisHbF1IiGcno1SHP
lii0qifnJwOyZ+M+UlcbX/4l5AD/fnoPlX0e5imX9FJFzWQYp3FQ05y7QHxm
BMckJggcKciT7FGQJ6xyodM4Gb3UWfKB89yRMimZ8k7/JDTHwNzhMFpP6xQu
g5857lLhi5YKHNxdDAVkpapWfUUgiEktIPYZ897Mn8uAjcbv5SwxJ2dO2dhG
B+ChgLnaNUiCT8FkpQ9XisxqTwhLEs1TpMqfe0M6B0dD9LOu3pmvr43JebR/
sqhMiUR1T4S4D8VRyWrs0iqYRu3G+h+3AIspHm7QyU4l8y3CL+622J3g1pov
Sg86UU5OhBdsq617IUIy2xr2pl70arYXIYVA3iSi+oYscsxu6k1tCpUp6ctW
z+nz8rUfITO8/Cuece88VeBurCCr9uYpJ5Yw9/qYeH/C3zlk8PxgMGP62sYO
AN8BY3GM1nlhYmKpgmnL/s4w/v/l79E8TeaxzXiii5OFvDFdQ4OReLU1rxFs
Dewz2fzOfrsLNn5eY156XI0klxq9Wqh7WRjbbGBVrcflmz4NFg4wA12VVoT2
AyjHEwgvD6TSjd02/SYoqbDfEj6m9+f95ozBz4vu3XpQMsIkHlUmlkPLD6kJ
le3Gp+lEeoGFBtPbTZChZ/BoFW8I7IZI7CEizkPR7D9Gq0Qd0No/A7wdZNAQ
QtHX1I42BWe7Xo3/zVJmaf34n2Xp2006iQM+RODjis7s4+obXGtpjuon1HFN
n4B5Yn+4hRlee6vF9ZpwmQmprMmfxjlLMQkFu3zHUvr0gAkFUd6aK6ybYzmi
nyb1d2sbYWmTefWZ58jyBaWOLpXasx5JaLlZlRmK/S3ZVkBWM6GNHaFQ5/IJ
xwHPkKyI5mGgn0TZLJSyrQsABbLIEMzV+EJ9SN1LHthf6nwb2dBmnphxeoG0
QbjKmDSRZPgqf14TbP90RZrZSNFdcIi8WJmr8bQ4H1TvsL/a8GPDIpRpUoHZ
xfiRC/aUa/S0oemISm25quYJ+nsuZjPwSZ8wbcdL+UQpcxz4+YyhASQmU5VZ
a1MdX+40Bnfx5zZTJs6BROhq9aA90dDVfSZtwn68y8DCWxLuzjjgn5W2KwWJ
h8OM7ClBuE7MSMuqQ8I3C0eJqcIofSq6YnQLaRZIU4Q7i7eOOELJMas1eMMt
An7NjZq6l8gJLr/7XYCubj1ORVlnr6DWCuO7i14Rb5Pb82mubZ2aG3icDbqz
Lt+f1NHyn0udbPlE/MqIETN4waoAovqPykZt+NRWrVgFj3qT4hMvbtXQPRto
FRTjONori0WlNSCgG91jrcsU5MA8KS7pLuvSQ7psBNodco1quoioY4dbxlLH
i/+Oh6V+rnbTXvrD7BRZQZEOski5ufcv0x4fqOqwyn1W51ZC4z++ofi7SN79
0VnbHRc1mrl2G86157Zn4SKKgO375Uj0Fv49OZhmekNkkDhGz2E2qFn6bQsF
4O6kOxyfRsX8QRF+CMJnlEKeb7K5IihUhc+BklyiMLa46Pwgl3gas8Tv04N7
R/79iXtyWo6uWW/LOsaXJ+KH9iJBb/NlH0oe+6a7IWn1cOqR+yg1nzVLy6R1
yvsHkgJbWCwUhE/R5y+V0GDnHT8PRLMYxUo2pY4MzrTOYIJwsTg88MzU9zNp
e9HOyhFjnJRmNt8aSnkTPar6i/eZD4DN17RHW5pyF0s+TGwAReUswJ34/wUj
lisVNoCFpgP7fgIwNnEIRhJccBXhcngdWeVrCLB5UAvRT1P2/wyk7k+r1TSO
dzKNuRmK6Hffs0WS6qMRSIRQIwV2MpftuQx1Ok9920YwG2snzDROQbu9ARPX
pc4aR+x+rT+6WagJVCsVu9gPw1bY6i6c+X49bb//xRIdvULxoPxoAFC4en/t
dp7waBBurn64bUgk5GXcgadDbRM5GyIwbjRpfqdhX7I5MecF2GTEIbz/LSwT
tUJHYZlSYMEs7fjpzCHltXxKCPXlOomppXkSeYWK5hk3dCBSINy6vs9LKz0+
wcek1mOfCXN1E7JDWiGPcwO2ztLK/Wpaj07aD3+g4c2mcCwUktmwRUJxpFyz
9kVdSGF6k3513TeoNfliRmqOZfNFjpSc9Xua4AArgw+Lawziv4Vk4yo0TdU7
0shadd7tiHy+jr4wBPqafCQwZJDsXxvfAr8yWnIBi6RyE0kGOpXCHQPeCRzx
28NgRxwctQgVWG6iPNRC3pQXpk/6veuJqkn+m8BXJfnVOloO7+vA6WWbKqwW
IHs4NrlW4+I20THnIHjQigJ/w8M1drd78u6bxhB4DndX/sr9i/tJOo6z7F8w
v5sCXI364POYLvSus3pJv1NaNh9J0B1FE3PZ7aW/h3Ij/Gw0y2DIciXY9egr
7+bDxMH1hsPiKiCWaj3/ZU53XpUVh5oWxHMxXtA2+0/XCNqpxB/bbyf2kdRA
KSNzZ25Rf3/XdH+RkLds0XKjWuHyv0D75j/t+1zPNWvii0mHXs3HpyH6hCeQ
pQhkU1TnCuIOWfKyAKmBYCjycbbh/8rzqLGB6TQEmGnunPTm6HwClFZeqUp1
pmqPIG3ldRzHG45R/ViqIVsbrulgD36VgxBBmWtEH9wzIXtc0fdP8lofAVm6
VTiECfnqYBhG3ePeYRWGVHp64WWfjTTb+kVZotcbuarheaQ57HBPQ8ijWjGV
qd5IsWSp36ZfNfL+ovx5wK/LJKXj4lJ4uBo3FW3JnKcPQ0wBYI7ZjCIkggY6
ZaDGCpbyDLsV5rymT2gCS1gTzIjQmc90qMDaU4Pp5bO2p+lOvlPAaOJLdYKW
N6AYbXxlyZ3FdgiK9rcGC0j+3jeQpr9RmxTIxV7hS2LwNcJKAh/TsOkRQyfD
3qdZkMn+a/ETpyIKDCWlHwyfL40HLKf2530TkpkLLfXXRtxT0OYzMAQv12nG
D6aUrbgFQu7WnA2v3wKDwoP/XI69FZIMgFXXXzqaUAbWX6DTkGPyNRh+vDGu
uNpkO20i6AWZ6E/lWISszeQ+bqMziTgf5FjfwiZk3ZH/l3huRZRf+y8oU7yN
6zANDMI8fgjrDkgnoVOoMjccz677Z5D/yC1iRRJAj+UlLJAhgwYo7wOM9l7Z
XitKjFeDRbFAuWVpuIsEPhpKZx0ltVSZHK1c0yOX9zPlaq9byDhRjd+hHlYP
a+hZVj6pp9HriFALqmeOQzbhOH4hpgQMU+VjY9KCEenAHxUM1mKH5+R4f/Bs
Kbqc14PThTDctoAHVdjFOoRz8yNLz8hjjdyD8bPv2NOZ8Rr7ScqZZ0A+kQ93
9Qq6tqJ/VFf39ICbwrZF4a9co4E2AgpBqbyURkPsl+x0+cWaVfTMdEqkKYO4
2Sph+BXpuDs3YadDHHcRTQjJpRjTC87sXsrLNoBjHWaaGWSABJjQ6pN5FFuy
3E7k1D+W+XFdka54h6fMYwquFqnJJX1j8xHiOZMQnQkiD7vJbqRR8cwSanex
gFbaCW7vb+bVNQOxocGp1/2sPIUoe9jPqzXxRfhNS7eDvZkw4I+XUyjXSSxy
MZsw4OXpR2gr9cnOOA9vpkOSaTjzII3vN21ed/eQ+q5W73UgvcraCe1BQUdi
AHOLMB8gqX3Uw0MNj3EoFmWm9TNolyQBEfDi6Ky5uGnuYKMkD3RN7dllgtPA
Fy6/GQ7VuL8LzRAZHjz1ne4d1QyQ5Xvc5W6JH7osZ5JhjStnMT43kP3j74Vo
8EnEufWRuIgJ0JuaFrdoW5+wb1O6obE/Vc2gbSZbpWv9vZUJQcWVxwXspFqg
GYXrQf9n/zSEc9IZPOMTgbI50yrT/sCy3V99GyhTReOUt3rH5flkuDjZVGlK
4c7zjoE83U2GjUIZsgg0kSc8la5W80P1vmgIFM3gDGbZkC6emqr7TBB44vmt
37MlIVtMkVypwO+3/H93ql9k5uhfMmblIM9Z0xe4rh17uKEXoWTBKfexC+FG
RuwHg/yb+iOy7IxZ+zEIywzl4ew0cnMAIYn1f8Nd/go4MRIAOtSPO/Hvj5Y+
9z6l/Jfhp6/drkqg17vd8pOYT4pndSSXFq6lDZOOzksbNdYJxPOUsOS9gHCT
sfQXP7EvaiDsq4CSmfXd/AWFX0J7SbaMev/q3/U+ls9fi4UDaKkexqtY8iYz
3j0zuIP3NjA4gCrCw8tqB5lQlUsJc2GPRKFYB6PU6IkVcP68KdTaeUG+DT7O
yolFjmsd6es/Spe6lRAEpBQQBjgpJAsh2plM3r0WzNcb1+8zEdW1kSVzvLbr
4Wfrx/sf8W0D4RK1chevNv9D9eyMex4BHsvv85zrLmw7NUxwMfd2kCaNJJCF
cFbCeqvOmdRnhgr55Elc5QGR2Th56GQagob+/d2FwNjQigJyDBSjFFr6Mha/
/lAp3JSTC2OwRvCZ1FXUkBDE5/56zUklwZW65qhE0HoHVdSn+AEAhc4u7Km3
RBU1EeVPqpgenkT6gqGE/FyQRDsx/ECmV0XdngHUz/QEEt4PnC/d94Xx6LNx
aDq0udTv5J+SN8vVlLI2ouRhznZ1laV3yb+PpvU2xIhZyCIejGsUe6IOsFsk
cNngEwDWKTt5ZT5cLFmpVOyG+ni0PATgG0AfKH/9dcxtVJaXgnkO3dfIIHAA
gYK9rkmmDrjYM/i6zevGHFs/BuX0lQJF1ggizqF+QsopxKESdMpuw3z5idx0
M+fu+ET50kEnrQAinbsr4PjPEYCPz23HhJFVPFiU/Cr+pnDKE6HUs+SMWhe6
wcAg+nYosqMbWahNbdW9k65wjkfuFhNHnB1fc4yAOb9TzBST3Up7AcC5mzQN
pw8wGyKrrSIYze0F4WxTRzUT0WK/tPoaovrc2ei84169Ne5dY/gEzOw0UZ49
vs2PmwvGRDTTvbZYEpYb/TOJy4dcFDzZBqKWqapEGRV8bfOyicL8s+h1yQ4h
qVIpq1RD4r7di9HH59x3fGG3sNrI+YDhyddazdbi3VR5vvvFQxSgAJ801dHi
PRAuutmL0LZhHWz3V6sefDI+dNlwsTep5bvLp3n4hi8FraW9PesgEtPxhZlj
mpi7DHuBiL3NXBCIBUGynJ1e6ZR/auhhd6sl5f2S/AhvM9KFEIn6ZNAYBXYW
rOeasZo+QDL9Z82RHCUceUxdYOqvIHhT3clP8Kzk1G7Pa6I2zcbnqNJeSzFd
owiVHJyPdyK3Lm38bgryqwtb7eLzVOqTn2JkY0lr5rnP/ykDkyIpWn74Z+IV
s4QG/dWcJOCcrULIF2+OBuWC5WhBHm9O1/pK647UOYfMyB9KkSox5k4iixLo
n5vDVmfGncEj0u4lvCg9Z+5VYjRYoj7UvQKD64tkzlkjVdNkPEK+pvrcivvn
EDC05X4rtSDOnf6drk+SBHUWB3cNYKTg59wnm48+0RkqNgkcpRxTMf9+yBMp
ov982v5YEQXVW1yBT1fGy6qW5blI8Fj84lck28bGLiNSykcrNdKocKHjhnpp
eDkeKw96o9uGkGq/8mwgr3rKE72JIwo0MtJcXLEOwR00pVXD/i1GJMdyNTr5
OobGtW+tFSTLPvCiNxUXwFozv/E0KuE3R1ziUnzLL8p8ammicyihMEm+LOW6
DQHoQhvc3Ew9XAYqRumrXLNgKzRexQXZU/wyGckRAuK0lidw3R+l3OVA44Hg
HlDxil3PyNYgzXH5CFDOpoPvKX0U+9La9S0hUN+W2Qmy5X6+UNiZP2eWUzzs
5z4awLfqDyTqeC63L2T+/NjN0rbu5AOXWbhU9QqXy9oT0hVvz/i1IR/29uZe
qtz3iKS6oHsNAy3Vf3ef5mwGxcr2xNgQ3rijP/PI9YqqUwZneAgKVKI6xrL/
sCN3W5BE841LRZ+rmyKrqthvs6N5MqAO+T4rugi6WSYok0MzBgnyIvnDX/03
i/MsmtUt6YMqpd4P+2eZAjV+Qy89HYP59+Uixz9t/cateIwmaETDkf2rP/AT
No2RhOCm3v2Tfa9zYCKwMw8rlBPIuvKA6cD+1YEbF1+aTd/ib3ypwsrNe+f+
XHH9n3JOug4E6/YAy5Mz/2B1l0YtCgNJogHEt7GmY8eexwNR6/XClB/lToVu
tANNER3swAaV+SgyUhAUcSC0MmqrVYvc6piwtC4aGp3lUJrMxZLcpJz3dltq
z485hRV08bTaC3/jM/UjNhkxqd+F8fVC+MLtz26hwV1tCq9duS5DSTFPIE2f
sOBodoFnfI+K08QZcalmnohqYuQ88t4046wj9Z7+kI7SUmkIHxXRhe0OrdH5
OBjL237rSWakg3KHSCBHG5ondhkwKb2+RM5M7H7vVvWgEv2HvlZ+aB9bHnf9
WPTQwcw49/+RKb6vVmKlWXPGRZk3q7ZsZkveD+QII62MREA7TGWzi2Y3BnXb
GtllrZyj2UiSqieTWl/EK4tkzhNROYW8YeO6KzDOuWleEQhz1dw5vhecxmS0
bXs6K5dOAodJEQYcaEKPikZQwZTV8Mg9/PYih1TqwM7lrVGBk389kdV+oPSb
ir1O887a4M2QhVC6WlzKJX/vu6JpNv3W0hmLHwESEl9Qo6Ox/IYaY3g1Maa1
z/rDlcoTjPRUueiGyFF7J0bw/7mLaeEtSChbsLzO/FQ4PzoxoO8Gd9Wnvk5g
LjSgkaxOXZnF/SEwIeNzC42APojV78+5u8LYy9sRtcCYDydN97Fe/EO8ffFf
kLyVN+imIcXS/X/7IBCkfmeTKU+FJuwgjg9kLLbEKAg3ZF8NUKINO7/XrZ3X
VcNZqRESql8kvmNKFn6YFwXzQT6Wwupj3MyIB3EtMhOh/Ad0SONtKohrPlmg
8KZWAL0/yGpZ9o+kG99mpvc081fgUPf4vDhwre1RozaL9KPdzyWUFeo8nS9l
09jF//2Y6xqVwrpcYcgtGt4Nlm8t1qSjWCLN2GA9KD7TF1qow9tlPukS0U2n
eQVxohk4sg5iAPOS0rn38PPrSJsbK0rrK8QUuFviwoGilx9HdQLK5nrY/YIU
coWcJR3e9Dvi0/IBStK4VHpfvJFXuZoxlMX+plqaT86pNoGiQeh4lagLTvlk
7CrkWi9L7Z74X2QIMyAYWFn13lVwq1Db7XMKT/ogUfD+17LJLS8jPc9q71/z
Sbyhy0AOEx0V81ux8wDmpt0Q6dwV0f9Qxqy+nvqS/XTPsyLzXzfF9/VP9bvF
VreTUecnN91F9PIV6k0MsCnuMd5dvKppLA/tLUyfRBl8z4bWNGaz7jRqB5Go
eCvbaJrnk8UQKfNTpYrYl0xU9jMVJJUhK/oHtZKxTiIUIkXGvBFekL7+lrrS
NXU5oUHu5io0nleQQHBioXFzfljyGtuoYHn9xK/q+ScNrMjNPumAhsIsmnAR
EuhkHtU2hBHEnofQSISdGygh6SbcYKih0bzVbWCCkFkJmewydGBhFdYzjz2K
98ScyQgG75kZONe0vy4pieJynw5km39YLjuqmyG85RYhi+8hXSRF6vwhOhDl
Zj4OEWD7f2QhSCVXt8rgU76Wlby+Z1urNN9m+qvrDBtrR1vlTmya7RxM2uhO
6bG+prR6Sq5lfaE15X6VcGnp+V6UMPvGOpVxq6xXcKwUyHQQPk32ucn7A/nl
jg3Y6MdxPXVszDb8P7ST/MhIy3n639i5kOjtgu4XwK1q6YX6M2aiT+AfSD19
mhzHkN+/YOX2aVwC/S2lUg5C0EeFrOVI2aRWuI8paj8P2btZVtAaFdvOkIPf
pyl2AMGMgq2slrMhHeTaf7SvE+mSVtDrqd2D4BSRAn2OOTtWRqgLzs5CXfFZ
kOZOViaQfKi8enDaCxrPPdVjP6brHJVHEzTtZAwoGFfJAxgdzYSSkhptrWCq
L5bLzcJ5efQ80CkTDwQrOAbTUBYmmlCEPpHZ/p0MVKl4G1LpPHIs+rckpxB+
9c90oyMTlJc7NSCzFLrcRZjGBpjzVuhAJZXv4vq7yN1C67PUkN0APlPIElyp
CdpYqm7JodP4+pgvyGr8d2QcspfeZOLZcCvXEKSk2j8gKeynx6LI9aLpqiKO
k0GptHv9f78zSkhKaprEE7X1d0sp2kRPxX6DQe29bj0rNDjPz/Z2cFRfOygU
708qaVqd6VmWxy13DgzQOYmxf54SL3QXHabSNk4DhYTQxf4Z4D77EmC1X54a
KjsocYV6ig/nT/PUW/wWy1ZmueyVq/V8D+eiDiGIJUm3FNY3JH+eAdNWzKRv
9hLdxdgmFYVTLb6rjT6LblwoxPeo3pm8OP+bXAhMkyM9A++ALOjHnSUY2jEY
8xCpCtqgqaCKvZN95G/qVFB50U64S4ZMf8LmtN+hRj4T7jZLL1PLOEjDti/B
2GfX9NHCru2R6CRjWcqaapO1wgH16wilyfrPEVFIR0gVas6aWqu7cSlW2H4p
/WK57L9OdcDi3R1edS/8pVooIfH9f6Rpk2KtCG99vt8uzRGpiulCoT1Q6+rj
B9L3M8qiB3pJqx6FzlkWzWP2dKCnuHZVuOZwafApx+JFfyI2UvBQCnlG9OG+
4Eltn2FHWURFhq778EHQYzlUEIl5/y4JvQ+JdMSYpda1WNsN9zPdEZB2UoEW
5jPC5YmDtwqJ6a3KgOjJeoOSKY2+7FZR3Mc4++nF3rMwKJ04w1Aovu8e9wwo
0ZuwdbatEEPW3WSv1/zeZHNw4WMFYxCxo1f/uTIRYfTLVa5QnEyn4UAvsH9O
IxC2LoSfGx96cwNsEPTKnVIJdVYyrlwDiW40HQou1nla+Gie1mhL4CASQpxw
0uSg1cs+RqDIUCPEcOswqmugsvWNpRHWXhut5ICr6XRBKCW4pZo7TKw9EZhw
DsHqLGnxx4mx0VM8ckm/Comi0vGCAikDaYZ73GuqeglkNBYiq3vKioKLNh+V
ddQnh/2Np19tvgY4gtLmwsp+3iwsXFeB63/SOZFfzEiGPBekuPb5ykIGnPsE
unS9u+flfBckoODLeDQ6QTTJC1TqpDBsEKztUyHdJrBKek1ou5yZuplJfOHG
BYHHEeel++8yvDAXZk8WkR4KghB0Kk9FREc8GZKCxFQelBpy++y4bu4K/Sxg
eVbq16YCgM8QU7hg6H944CjrEUv64xneivdzh4SMbKIUfrApp+/755bH4an0
ViSX6iA06aA8R7/MnKCcuimLYHljMKWFASsYk4mYgh23u2ozTJN6d7PO+fos
p+utkGkTznSfMM1gxDFMlDt35fwLsaVIHktO+Bt82GE+JHyRSFhYMNPPVhGy
dFHXvKH8Ae5pbYJ6QvGq327JiQyZuFVgJyyUdkJZNWldqjSbPruii1fx/bOY
5rVugzIw4nSaDhYRQyfTpUeFRz793WZT0ZiQPTcfN8lC5Vyz7KiysCU7Tjxf
5hoPcSTjk7QjyUWYqImIuqZsYHq53sXuKcO3hdn1MynloLI3I1++guHM9P5N
RlfCvok5kM0AgvOHrOAoTvSWWOeGq8HF89kTr7CjLzyctvAGLsq9c1kI4+Wn
XZfSH60z3MAPcDY1hpQrUlyW6HqPD4k3f8pUvlLqeKDfiSMpwqg2moDxaK/G
rKNEj1DVFVzBk8nc18Ga4OnyDDB/UQ/j4UrfXlhH/evaagp4wmuqCmTNPfhd
meT6I8musin0RlLU14kMvTjtm7ydSYvgcGjc5grmjAyjfCTFMRKmoANrTBTi
vdwxFz+p+mzxdLAHeDdMXX43//WwnaXNgGTnWf0LX4PvCqL7OPk5t55rufjV
oN2iJe1r8qYyEPPaAs52CJGldaFMCTiVnAZYkbDn6vHIkax2cMFNqbL6CtQd
/6qtmit0Rw3bsDGOxbmUYYmQmMIYwRndjxCZ28kcJqZNZWhbDKd6c4u9nP4c
eyudI74po1tmysCigSPaYvT63LsvCKOYFx4kjD35xUWJLGOmSfeROalfarWR
ejEn9F/PPnaZBgMsCa4p1Scx6oN54oaXG9WG/PJWik92o3UmIZBs5liM8Q3G
OLbJw6gE99pDjex27RDb2JtkK3jBSgOf80Ue/qktEn/Y6xQEkA8VRW2np3aN
/5cxgCAkPJvxZebWJNzQueMEXPghWHPXKv0SlWl0jGpcbBiBIr3SNaP4utW9
8MwI/Mods0Eqr8JCeQ44iJaXyanS8PKSFd4GI5pXEwsPW5kJl8GHaQTfP4tq
6ERW8UtCtOSfAdfQ8mnKT2ZjuhQesIFFxtK063s++PYRD00BrFXJjP3PKLkz
Zzq7FlqjUTcnDf/J/4jZ6l/x0S8I70ALATl0JQ7qoPL/UTg1Sby6ady/dpu7
2ULzoT99sfTmuGjFiswequ7m5zFeymaBhtBHxmN6qZLyEf24iGUPPD5eV7bV
mheGuCR83839WrZj8voxaV7qLpOb9A795vMVizHpR9HL6hQOBKP7IF6j0egm
jvM5QWML5Bw+xfYDLCARWB6gNpfU9BffB1NQqcgob3lQ4E5WJwA+4K69u2Qs
L/m8Shde7L0eWkb9FtDU9nra5Bag7VbeemT8NAe82vIf03T/v7sxVTG7cPb+
x1sl1xJ//h6ZdYCrcjAHn+ddR9AYWtDje520W0Uy7SGdmvXHEaGS/yFqRHw8
GAIpllEdpHkBsEcU3ybjF0QSsJL1JeYVa7EC0Lfj44EZczk0lkZY9fj5CfM9
2CW2/cNy2WF0IS3idOlGARjSxsxR2t+b6znuV3Sw8/nf1lhCdP5Ud7WdUEbE
ucSQ1u5nrxFRkCZDPn4ZoCh6BgKuA59FZHLdzCzbbccSWcf7IZFYwzf+hw/2
FUVYh3oYekkZaAnxiadoiWjse8Y/q5kGinG7cwoFjtUGcmUUYX6XVcpFP6bn
mouXZvEIGr8DUVQOe68GnAiYDecSlRp51IdMv6CGsft+u19BYKJFznBz62aP
btpzrDOksejf8BgPRLA0pwMOCHdri7bS1+PNRw==

`pragma protect end_protected
