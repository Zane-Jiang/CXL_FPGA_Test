// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rt8zcBtNGB0DvtUE/oxFYN+HjwvPKm0u3L1BXMk/nKqmcyRxFmJPuWvBLnRB
n266kuJh2iShgiSCQZH2kUfztRGaNUsW9lsA3JfmuRYLUOS+ugFsnJuSjv+n
xWzk9bed7w20psY5KL3fa03pldVxMSMayHRIw3N9KZg86GB+UDNG6gtolIH2
9bjw+lsjUGrOw6iawLJGKvt3AEDjHcwJUBpW3UC3b+0e+VBx4OL+1+5c8k4m
isxw8SqH+3juWAavzOg1pcrU+J9odppyToLA/SurlH3wkTCSdm1U9yJCO4dt
HtQ8j0FV1VULwhTL71i1Wi1z2MO7Xs6B577bX3eXog==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ChhcCYBsD/58HsmCfRGFyedsIHX5Prng5rA7fDG7i7+NsuMp5xbWFS2vDFU5
e9gPmsgLSgsHl+Tdzbuk0sBUlfutjUZ0m9T/eObFI+BbAtjLk4UJ49GPJo4n
HOuIgTH2KI9EeCKkvyfh3LcDiC+WrHYTrrDRhYGCmndDonkJ9R4dU3eZo5F1
qTqfS//plV3ulodrDBV4/bfkNwnwejEDB7SZaIJemc4JOQaTgK89o5iaCIAx
HiT24hv3w1FxNcuF2jJVZyuJLzQdAPgCXHbxIKFmP3clwSFvSf3kgEPBzCd1
Duba+gi9RWu6BlAFKSSn7aT7nMLJsQPuShA9M1q0Gw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O5DEpxFCbnabgZbOxlgO3Gs4SqE3BQkVZ8rwQx/3uXzShdXl2hHkMCvcQz0d
sNEm0rbbi9wYoKtqWrit1ChumrWUNWmg48tHbXDiAPALwqliq9ppIEi//5QC
1aQsMJVcX3EBUXLR9q6JCW5HTcO2cLPDa7haLlxbxK3E0CCVDtlGL3+Z4u8h
t+HJE5FmHXwzC6fbDwlV8XGM2NT8YGLqxzd6Bj/ExhktiA7wc5V+YzeLykqU
++qEh6CuLns765c65Qm2Fr5vOpUzFWplL2wByykc85JgEKTBNevxr0igx+tM
6rVyXm/FmH2YmM2EeiWtvD7cSroaHYf4x167fsintg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RyP/5sluOHGWTzaj6vL4pdEYmi0IY+AKRTd5d89P1kA59bVmOp/NU9GYfKEV
A8VoLXdjgCyM+vTj7VF4bsDFayZA7a493tTzzhiNpxBb4xI+WTJP5QAjIXJO
BpOtZ+aip42pu74rq0aCfU87kAORGa0HhFtJtSo+5A/G6XVXhZo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ppX26cdAL2d8Ae2zSCWS5Ge4fDZnG6R7o222kYwzo04snLTIF3KQ25f62WCo
30nnGzaVFUWH5MuN2vBkRUXVIz5k6TI1Cr6fcTBKWKX5HSLkAtTuKJjjMPGO
jA8Gb6jBpu8h8RVytu1Q2FhfrbZItlgL8AUm0fh/2ejMhZjZJ4EYU48g4IcP
35LWSgexwe67G8TPWNHiowvQjJ25gejESrHAtEk6JGd9MxOodUoVT0MFHxhE
VqjF/Ywp4UI7YcTOXPIJ+bwcYtjGraMHiS7qdOQpI1D/8V3LxQmNEjnLDXxd
LTFTM9toVv6JHAwVOOADTtYtRRsduWiZGyLu0kPRE1MaEr+UwrU8FSq6riJf
AMnobX/Ome5tIogw3dS4oQi0vY4hJI+oFgLyxop++TOtLJQWv7FSNDmF0rU7
aibQiHn5RPN38Tkqm7OIc0Y0sCIxe3F/eKcbKmo87+36hRUO+W+ALotL+H06
npULQyEbUZjd0O48aX80GG6OSS7gt3Ed


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oJbB0J1XAwGS16ZlAifj++rFlpreqzkPQW3RuyxDQ7Pkc0kpvPj1K4vW+O2l
+6zDjS/TczKFNlypHiCBG2B229eEjM2JzIFrpEuYNcQvaDph71RwSv10m+EJ
/MNBkxbv9EoJkSJuVOI8dvCgJ0IPueYdw/qaA5x7FBJwNiCx2BI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A89tX/JB2LmA6D7nTUtqLOf+mFIyl7SDmBvv2vxd9A/JAtiP237gODpHuDN8
s6AjGTIK25G6srrlxgStBG582VC6lzZeVYipqeVQiMiEc98HGF1qrhrjxZVl
dj4OlWX1RpCKy/fE8s1VXnMpxH6XOVXw4+kNv6cGC6xXid2MNGI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3296)
`pragma protect data_block
XUWW2VR6U3pKLw7OhYgucbSeK0dc1+ImRHpuzN4UXRmiuMpATpRwInPZKvPY
k0HpwR2paBSP3b3NSDsGToWLT/3R7uM9rWl3sueJqkYGJpFXe78/JNnNA0SN
0zsnHD3sP94QK7fVM5mVpzyy74a6Hg074UpVAGM9+jIl2xbMC/GgZUxc/eBl
2O1p7v/2PsIlDMfv8IACFKgjQ0zUO91TlMdO+0NjpH+AVxdnVl/ugtyuVOBr
VhAqC2VP21NeNTM7E/75JsICN/8Z+60HPQVfgtmfdV0cWtfjEAZ2YftId8AG
hvPCylQqBVrphvZr3KYwYszMApoiMhaqkvBtYxRHDMWVpoRJCO8XD3kiorPv
4Rf2sQw5AJpMLyN7Eg0vwuNyix7vzo95rNmDXwn9CpvYZWHU7dGpGIpsrryT
7aoxLsdsaO185baK9XLN/aX02HFP+pG85NGgftDk2KquVGl4xLUs5NaWLoN9
vcAIBVIqJRljCg4O9i19bKLFC4xSBrYKyUGZqh/n6GVzq10UJ0KnQzNTmaEO
e4qQ3rjqJBCPDJ14oKTaOxgaReVmdPtLdR9wGGCxslFRmfbTHfu2NWpfS+fe
WglafjNtQC88VnCkunGK6eSf7VhX1zzbzfKEP1SSad1m2zZnXYagFlBwn+Ns
0eBUB86IMAQ2K4Q/vKqMD9a/zVlvhZjYgsN7e/+hKoWKgcJyV7i4S0U6wf0B
zyrMtF0NAgyWj9a2XLt7u7JMXeVlYav9j9DpxmwbIf0tZGsl6tqlvq5PhkQL
jrHFIwh+ANJSil0n1e8VsFRW/MSmUapQ8jYIz5wsM+US3KE6z4j+QaFhmcZO
vDZOYRfruP8F1iTDW6WYRI3sEMfTKq7Mz8qv2dBL0DRCPLjTWbZfnMw0Nel6
cGtUnwTAIqiy5+nnLcYFXx+GaQkziSpdB/rxpxxE7Lj5hoqPTOYia1zUYg0l
SZEGMYFKTiDC25NjwI8bb3ZaCMQUxagYwLzzQo6087nIe1A7FAur7zAxd00/
tA8dIiG+9olE5UxGLeucdPbH5YyuwQhh+65yTOEGVF6OPdE+Tzjh/mcgiqGz
oKaSMXQ6zsM/50OcuPcxmTQh4MVIKHUI1xHVnaxqDCendviE5NI5gfYJnlCt
BBKTfWRMxkDM4wY3Gckq/xKMHoSBINuyeK06bEBffiFpF6bevBS4JJ3SYScj
4tbh0skeTS6vXRdL7RFZOKo1jKGe9Yf42UvSdFIKCGOfBkzoWF4L0xvwd6Rt
QC1cp9Il4AG/xn626VFjGbQ23TtqN6VqPMrIChZJ4hGvr+tTUF16fxqzEAO2
/XUnFjL107S7O9JBkmPXnXYWqGVgHKUgTOWzQq1AOfuSwiGdNl77E2+faBiQ
HwYUXEGJybwpMtxkU7385t4kASHlc6/smFy3CXfCUvXLOClp3lLs7VJvnULN
EjPxJ59/o43YparTudRpFWPk0vrlyI98jljZgd55YPO0XeHcm4BW+fkQBWW/
yTGTLaK9J5DusqT8ybSb3Of0Xurh/KQyORoKCsBxAAaCdhlAKMqdp4Fz36lT
2s9bSmlaI+NXtDy+c0SPG08octjHqNeCnqvGKMoTVqnDnTZw57eK3IelpIMD
4EPQmTLBlPU/Z+iiPSV2q4oAdI7ywHDC0iW50Gogn00cx6MwK2FeaZ6p8gI7
ZnDYmvBPlhIktD1GU0KuUWoX4ColcF7iOn6SWDn2+RLv24JjR3viLHtfuH+s
UQ3SkeMOKAFyzXduOnVhjyqQjsI3Fw5qWNu9Iz+2Ro6z/replfDsidTbe6SH
I0XPqw011OAIhKCLRcZqo8E6mT0O2yb3iH+go6gf2jCeejVFRRNuvq2duQC5
jhP10o8sof2yzyEAmdsd/Jz/cto0J8ynUCLbsorRTrS44qkXOmjycKY/i+Sl
Agnpd9WohoZdrEizfz/EEbsZoK/MNvzMp232B6dB+AX5Sg2VD3uZRB6/TCEu
LqjOyuFlajytehjZkSCuf5nA96o9n9W6qxNCWZOpRgfM+gCvGiF78qeBoEJi
Ok3FjJh+nWlnTTPTfpp1M2WdzQq7wvfUEVWQcG2GW2YbmYIjkRF9bteb1vDF
D+RZCw/0XBGRdeFrD0LMO/pIfG5WTW6Q5grdTeHi3cjbzdp8isKf/BBoPHAr
3QqZ8lau1onAbkPWEEcDcLcDJ4qqVDo8XcSm4OadZ0tT1K+dz2HWGTMZaTw6
wjtDD+S0F9pKrRuNCEM13YI3UnTvUwrVn9Uig7YZtlZ+5h2mnQ3W5nfhTu5S
LcwkW90aC88vIOSHgf8Fw+31yhM3UgYhwyS4nQsUQmYJ4j1q3ILgG1sd2fN+
kplbXEijrjpnHkJUhTyeshkJnuNTbUdqxEbWo7epc4F2Uw9blx22zv+u6BXL
sT8AFKOZv93eLpWeqyTJqkVfzirT3JU0CRhY0UXdtf9V4LBRpg+3dhQXqn3B
8Bcynexb3TlIQRgKdDJwy4mn0tWo4lmXiGHQzLtRumZxjytkqpt1p9mEPV+X
R7s8MQV+WQWf3c4lmbFmMsxGYFu94hmDw/hdjGHUqXc430uJSarvp5FQ9LqY
mIofRbli4OFYSNWFdk6n7yvIkpb9cTnJSGrS04jO145EdCekWueSdtcJjvRx
UjelLzInIotL9IjxWIZjg5JzcA+/SBube0C5vQwh5NVN8F/EVJwhNq8VsjAC
Pi0+5O5K9GdaIdR/+47G7IkB/0x4xy4V00sK4GjZePsbBGgCRXD+jt99ELx8
fIWkM+n5kWNVkdgXN5DtWPo41TZpnIiqes1FgYzHMo0Hb/R7TmtB4U2WdOhE
sgVjksIjOfRI3rCFWYi4BKxYi6R49peAi9Ns/xu+J+gvTtTKyqVkjBHfi1zx
2iL4ZVsRqr6brmAhWefAorFO3hUOEh722tqTrjIUW08eHEhiVewdqlRvoyga
QYAL5sl+pVNHtYqxxYgLFuK3/3LbwVuojLkdxNDKQdhYthtAgq1zPTqKE5m/
q3UeFy9QcPEh8slxJBB0c0rriAyw6qFIrsuucvOkBV7+mdsS482zHWkYC9cV
G+Zc91VZp2O2Df5rQezGcVu64VIeiDhyvu0/2gz2xouO+8nrOGJ45UHdFLxQ
zMPPsI9FNiNWlv2TfN6KUSDPYTNjBUdNrCM1PpmztWrzzIKEXmnQnHYyv4c5
u411HRQoJDyHf+3D3/IUpYbJfCam8+FLlbDSsV4pasfNEtfXZfQuqaVGDtbZ
l2roLD/xLFDCm/EAxDuz5MHPjMw0QPJVCeEv2D9dD41d+uCpQVl67KYgKBgr
tDZIbJRISu0JOzzG1t1/mdy/IxdzsKsHePcVAD7hyF6LmyVXLC7kYFCZT8yH
ijv6UxWF6dm1c3lKtaa4f20EjLcxr5qiZ4MqJPkwA6wRzbmFdBpkY7LVOI2+
+YaLu3SQki9UGWr96VGeuvHJf135U+Py6+Vh36vIrHhm+0P7wpgeM/Ny9lXG
XVjGelPdfcJ6OpsYPgYmOWJ8h4pRC0X0dhc90ZJdQXyBfjTfthLWr+54NgVy
BflLl5RTTFugcY3SMKhE/Uka6JxaB9dh8M1SXk5HTEatIid+6Cc2tg0AD6LA
0XpghMOOpTmsiOzpVk7V2rAkG6c4gfAE/gqByaC/pjI9BV4PsAEHnL6AVtNo
lvrBp2+0jdyhWqpR3CQDxfkdhWgNyUBcSARzdx1M/CgLtUSaYkEhDsDgTD7U
30MUHB6DgN5Slae+rDaUpNHeRKtiANrGyYmhtpRFZhG75ojXqCNbYdVFxkPp
8ppjb87MLKqQTwnhB7CElwyPrZa0Lzq/d71s8yTpEf/RCm1kaptTFsSyALPf
2ZCE8tt3T+S1CjSK2XgysvnHa/urZ8oDIXO6rsUNrR/MlrXLCqOVmcMhn65T
Q9scmD90cQucmj4v3aoYfLfxFDUKm9tfglEpcla4G6klBRplLFSXwM1DVjW0
y3VYWCuhRuPQy9VvwMGTmfU4BxoYWCcPCgcaIcrNjH1x7gkYEc9AiiVwEszi
T329WKIdKe5RrqE1GMg9Lf9FNoU+iM/sNuQUew3dWUaQcd8Z22FzSOOE/sxO
dJ7P6ktLybX2Sy5Jg6F0RiEUd5+Mx1YDghQZCxa9KkM76yKiiIy6q4TyqC4m
2qimM/Zz6yZbi7JR/mQxadBa//FLIc+mrwn92U93ucxZHGwO2GGihcWwsFrI
usVa+wcVY5m30zKOK6McfNTbAJqskW0gpITRWx+L81RWB6Zb7YaYZ0bI7tgl
zdO0DOBr/5rVQNL4ZcVl7EOMKua7EAgM8jAlu1CDGhgxZufPUpT/DoNz6kKX
eCQbj0fvkZlFEpsOOhqhIC7MU9/4JXE5cXyASSM5UZBDVeS8CcEz8z+2gfJI
J3+Y+7vKNf+prf4=

`pragma protect end_protected
