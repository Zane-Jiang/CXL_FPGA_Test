// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BE7R9WGBiIyzGbt9iNLn4kl2mENEaqTqsDtwGHEAzDHQVNLyLCSnhDGpdWCJ
OpcVsyae5ODfWoMw6SPUt2Q2UXv9zg+22ZSd5h1PQuq2RfF9EEC3iHMGo0fT
LOZyvC5fMY4knjFAeBp0NPmj5s0SdYQd+stChZd72Keq6UpI7QPgoFg1Xpwj
JHjpH+DWV14uHPIkf8M0F+hAySH1F8hvxitnacUkJyFuzBgmSCca8cRrUqjN
dPWutxp/kqDW75L9Djsgw+DUi/3qnc33SJpGdGcbbUS85SlrO8TnrB07N2hc
uitI6XM2xldmZX3pz9JCZQiKWFLF7k5T4qMAbgZvlw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jMJWo4Tte9KN+pwMd5ZxM9IfaQZiLT94CVOHP2ycnb5uRQKM/Et7Stth7jmM
IPigRXi9WfeMGg8t+CJ7kh/eEH0a3nWaTOq3OfLHxK3vTBWqOe3PVKZbcx8L
FNeBImMe84c1V5s5s+QeikFye6uP35Glp8ctpr6sCO2v85KHhi0dlaVIkfz5
B+GMfTxEgTSdulhyOzSvv9PQbhUy2bMg4/B1dmScDOZ6A73kRLNRwEa1D4Mf
fOJ/gzAbT0mb/wZt85uWCntJXFYc1g7jBAf5e9dMkL/UdvxjcCYT3jP0eFos
kIJlEgXipBa1LoL57RTy51PQD/QVLFpoiC8Xuo0DAg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y+Ev1UzexCikF6aRX3A08WheOna/bS8WknG3pTlQu31ryfnXbFzxS+k1tnfS
V1ci62shXFXQIkK3mNY+s8yDMLk0t1RzMunthgcxiF1FMD9dcTDAjJCDbFdd
GdjyF5Pq4bzsphK46Fct0ycW9lptgJQKDwNGsWsyQQJ9JizQmA128/cjvK56
TaE0IJoDRYDodcD/TM2xEzlxyF9STyHupW663Yi5q65Uo7cvueoq3nKQQbzm
ORJDa8sj68/eWp3NFNZwRQa+GE44CwZz9I0YLODAMoekFN6tU+r7LOXC9kTG
4DNt9l3mQEPdCIC4UodVesDNUDDGvF1kzkh8qnBk4g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YusVgGp2XP4aUKcwvjKWCIegR2pMm82c2U/mLOXc9wDpfjY5LAlVsFi6a4km
ZDrobAWzbU7tiinbZcS9z8xq2/zWoKUgoCIA8YblfqwY3M2IcFKUa6tnEJTZ
1xT9TIt61QpiCLH4aqIGaIz+OxDAXy4Xk2BpfeuGRUB4TwngTDo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wMgZtbtOl1KdF94Qtzzz9XaTvwnvKiL1W0P7zKfpOvJIjPGUYmIjZnzh8QV/
Pv6VHQXNGCr98HhFQEcFtT/hyCYOpFV6THPk/6T0aK3M/vOtbqFRcQVi7g6c
qh1fRioFw793NTF3XxSRR/jTkW3Mbt5vhvOJoCkgty5B2nzeRQ5o6UK9yqiL
0seqM6u3Rj6ylgm3RVcPZXKPhqJTv65dsGZinNWed0eoY6qrCbHq8xY2H0tk
jsYig2L81l5wdF5YhfYU+cbTBueSoKBIngMZLnoj2jvrKI10ruaNZVlqYZZY
jQ+9QPuCcmEhDrmQdASeHBTL1mA+bbnyKZ980+jBv/cNq/jo+8u3ASJNmFyY
y+guhotDoJcXfEP8AgrbHzA9N9MB6S0ss8M8s6DYpmlyErqenwGNZxqlGfL4
L0FOYUeW9oovJ7w0U9tU9yEGglQlBiOcf8U8Au/u4Ulm4n04q0ib0PN2f+nL
pgNsPvbVr4bsOKMYlrUDVF8F+kB26D71


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h7R+pcIdNvMsFXKUw6TaTPToM+jr4t+pMpvO2e4cauLOEXIsh8Cj2oiewUpH
sR4o9wO/Ilhy59UVI2NJxwgawR5i7sJH3E1ExuQZ4Hh/n7/TIpMkoP6hAvC5
OEU3Vb1cMMepZHjkPqPQj0EUcnTyyHPF3eEfcJcTsK2sZMlCKtc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IQVbu5iYz9hipYLv9qylzkBwGA00IIzNBJP5Ev1gtptaXNE8aG46Zco9iusC
VDe7I12BbBJv6A9Qt+UoeoICGr0NCKWRPKbjFd8be2/CKYRWYR5W9qdWDuWO
EKU711YjUSUFce5HNCEzEleYuHIoFbqeQwd0cgIrcSvoGTaOl2U=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
bG1zF3kEqLx7QlXafiYpRBqJNwCKxOJGdPR+qWmMmLN9yMXVzc2Ac7Ah7vrg
MLvUNo6DmjHOFbGlF2lq+y9kxSEgQy5UNeAXyV1kW6TbLwR+YDP+ukTBeFcI
sT1YvlBxJY4ygdQqhzxoFglA2+tlGx3P3S+EO1aEatj0YMZ2xhYbGyO8wQuj
hRo2dWRKUCyub9RJxr+ciU9UbJnuvG6mW2FgkHLncByGLcb1ADZVIeW2QofE
crc219AjyvjT3SpvBaLUmlF4ZzDnL5IpSwsojhgZp0hl9zPtjfkxGe4+4xn/
BZyVuGAfueoD55LwroWLzcukz2opIrhnTwvnT9900fTh2+NY2Wa2WVCQCifb
TAaji2A00XxCh9ercyaHOjOFVV9PRh8ac+ra7X5GEJmhQTozr+1JS62nzl0Z
fzqvWa6gYrLP004N/DWWBOXxjqf1NMkEbbSJlLBq6l1xGMc3DlJst9VsdnLz
Xv1zlsy6Z62RPOfl3U8gwkc6DPwBIBr/hZ46dtXOgAVuIyetAFj+jEOIy3F4
iohrLrWd3xsC8Ggb00RoA1Jpg0yDkpNd1/EOJ1zsN+qlRSa0nv6fMFGKyqiJ
cx4JQF17RHpM9WrL9uj+ufq9wt0dPn4V4oeLf4XYo9vBjJ3z01HIwut0s4s5
H85egtcot1Sg7i59IPEBTYb2h7H8j7S8h3yVSz/32SgjTRchwdyOyblmaXMK
OorPMnFpTb+lNzZMYFubg1Dv6HYA0BBq9jYgYh2HerQUjiT7/4ahj+aOPHSN
lfkSNsqRfsMQq7WaiZVjf6hEcQ+ZqOxi2B2ISJijAXFZsPM4JiGu7Zl9vTMX
4ktE4phCDA5ybcfeGTA5muw+MKq74A8fDbPaR5N5Zjc0l785D4skd3pwpBLv
hTByc1zficnR/OJ43QKiUUvoBDN4BxOs/3FdP0zTVNHWo9vny9RpY3o6MF71
2FS6w4rzN9vwvb874AGgrLZVCh/K7zV5QLd/I3Xe1Jz0+jjBsbwhSb8Udq23
2xwa9SiKsgKo65EbR2OOdkYyNKq8R2iPLpO/jDsfiAyWRa+yQ/t03zYeF0oW
Mt99oze+LuHISjU0DgXSuFTOEV3uMJW+n/ae7P6lJtRDi8gPnXHZ+GhQZSw8
hPs4muGVi0AHKiY8Tst1XuEaULhKLGMxMlxv3GN6staxn291wbGpIDf9RjHD
JHbXskGAN4HGJnAlpV2aoNsTBjJwaelDqTmJ16JT8c27YTSXrIGD8vY8rD7c
ACEQ/AkYv0sfVYnz2Mu+z+Z3CYAoNSJUthekbal0iNI4aEWwyhRRvKqK7sWr
DXcCpW8hMY5YgEt0yDOvxwtnCnouGHpspQq1fTY3bdsfUxU5G9gPxV3tDbg5
AwvEa8M=

`pragma protect end_protected
