// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
xxL2M0wjh1/CDj7kiywr1DYHQXtaNofK3FBr3DOTSBnyjLnSnYQIAtyDJvwfYRt3
0S+YYP+B0scm2PRjyOEejk6NQysPIXzR3KWDHka5xVF9SmyF5QnEetYIcOoLB7QQ
fdO4yuq5AsZMHMVodyYFEWhxSwQy58iXsHFhz4XtwhQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
Vt4SThAfxLq/Nj/VJzcudtdxtRItM0pGqIrNrWV9MX8EZV3+THz4CyQiNDyQ6nss
dEU2ASqMIHZWdLE1X5d1FDMWisFDDjlVZ3t8eT+8Sb5+LtAAbyo14TBSUdJBW+gT
PvLlP0aaQTWKPBWIkssHB3VtRmLXWdHlMcXk6CePCpwZ+uikV2up9uAtzkHRsjMU
lCPpm5akXcmstKXKWdZA6Fg/3ulqVlGFPUEnz3Kc00QXEJ8AqttT77wZS2aqa95T
1/p7MbOPJQ54EPPwuP1YTLygfw7ReHB+GRkV3JF+PV3d6RoRNTS52i52gZ/6pwOW
wLiGLs4eOIfNYo5iWR96AuhFWMxbhgnutoYCx3Wjpf/AAOBCfDCfLkKlObmOzMRl
hYJ6Mat+FjFLDIktyCh4hIpARYfbnD2eLuXJqr4Enyx5NHZmBfZcYpas7Q3qJNaz
GKAs9z/q/uxyP9V3PCmc+Sn9U2Udmq5DLhearToCV/qNX5aLCp4bNeZcmxWd9A0N
dFdpIFEVplLb7L6C+OYUKJE4PWMibvAivZSSae6O10qFG3TrZr1Bc9EelpTjCvLi
zHi2CN7NdRags04dYiBvACZeQcGpdRiVeRpTGCtT7wnGmiExPATRNPAyxk27mAtY
v35iYNO1xXkt8WJcEYP0km4T+WnqgiqqXAW3ud39sgwkh20fBCy/DqDfnguRGhGU
SxqFm6F4ttgfBYnLCu2xJIAR44MU+FePmJ734D52B1sq3/YeOXSssQ4x6l+PIfsq
8qanbDJuXh+ujYnzuXDusPmmKsmj/WPppNDAofVMOfA6+YCPnODhppy6ojDqND3Z
YtsTqV7CRZxMoGbEqtz8y5JWGhafgJ2V8dOG/ge0sA9rFUej1ypumgTfKSwj0V19
gxm7r1bybrKN3GlKxW6DQZrSZchrVacUzYbtTcy83HVNd6nJ9B6klBE0QnZPahy/
hIMpoO/2fR3j1w/+1Bff0ce47INzEtin1DiMiPgvyD23p7XxutEHWTZ4NxOcQO2X
lT5OWufNooqO8tgCXWLzrGjtMQyaUh/r3BNZHQ0cF1mG8i87+qXW3GvjiWzAs1yT
BOZuGbIjKBInnQCFUCjXyjrHL0OkCpbkPfhGxl99iGCwZkxn9SQLm6uwAxTPEk/G
TV1AQaZGiSasoUcsuYOYpTOlCF4h7UjSQo+mq9a1wdBNenkElMflFBuDONI4otqs
TjcIy3qx+eLUVOzE/+7Ypy+lfA/i4fFeqBxQ+Ug9aGRDfc0ae4sckJX1DYW0p397
XwZ3uZ05ivKcCQ4CuWXlSYPkWSfm7b4on0uyjjHSpl/wm6Iz1rcG3J/UBMygRuZr
SzfG6HteIr1ygL3ZeTrQz0yyYVT2z1chACnsfhEFVlGkpjVlzVpcOLzX8cx0xBag
HXehOYFswJ6akdGyMtOLaH57S+AVPphDOmWqBFMoDTNZSYKtVHAyIkk+z2PZB/8f
9dD682uPYHo6T6nXbddO1Hbh9wJ4CF3GecaWvyw20PQMV1xzMA32EmvC9okpqVN0
Kr2tOUMErsVuw8ohJvdUHDA+oElNvtokJtt0c8kHKbCIuXjqxNx51UCobEMzOmm1
wcln052wAu8T/dkBmYoXQyEMSiksIyiOa7uSZQMiJHweOjS6su2+a/Nh0ya4YaJf
JD1MFOdDDcByODor+/vAsJn5W33O9Gig83bTqbJc0tl9wE8bCaCXyc2vR1jz8qN0
+FkcaPrEn1+UDElLr9qHhC0xl0H73Z6+9AP8vHfO66zH/tEX8pzB7fZTSiwRSP2N
oLKw0Pb5Peeai9UKzrgOxcK35+3f9rGJCesscB3/HiGJ7VzIeHOmMRnzEWwm3I7P
0HuNDoqir4MOh/Rf9Zky/HySZfUTqRAaernEVhp4vnNL2oyOmz3NzwXJddM4pXw8
LtHwQOHk8c/iXKeimg0WW9t5NrKiFfGGP8uZbnAJPbg9rl+OmFJlby/4YEg1NOof
L3DzKH2B+DLCd11kHdECkXUfuGtrB6f6JfmRF2q3NNJmLNxNv7LvAGNERGwd4BvH
P+g7AHcy/ezWDZ3Ei9TztOZkbUmQbfdi08v/ypWaTDYJjLB76uuJ29WTi4VYAOf9
+HBLh3atkiIHXRtYCZQfmnwLmyllbzj5kYh+iYFUzfZx4kar5gYYJY3axdX5xMIX
XAWAuhdoO0AmveHCHm/SxLWYBqXSh9ChrgUh7jzHsDDeZRAgzzT020Xk2yhRLXmG
WdQG+b3kKNOmVyNyAooFV1q6rZffvwcxEAumcLexWqy4oYGq6FIZU/cMDbOu+jyJ
+aSREn/62YcGsPIhU/7r1e6Y7oAwv+ltLp6g2/RRHRHrEPVtHYbd0nggwZG2anez
6k5LFIFqMf8/a+fSbzTDrkO2iJtJYV63ZW9X6fBdTNjiguQhPonAK6BhyZT+/djk
Z7lpafC8LS0IiuqDxNxifZDf9gWmlZ1KAoYXzvvthbdcujoh+poew7CgItYdvDaB
RU9iWqoetWE2u/0rqmhTdyVvPQ/V36rHJ4bhv1q+5cP+Wuut37CgBqrMcyfni+WW
SkTiMG89HkNotdM25Gz/1R6YH7MxqVqJ7a8XL6pQ5yAFYdMGkgQWP/E6O960OACx
QtbyWwFsDjtpKmgwu1OpProf8SmWDJxbPzs8Ow7g/sEhvc3eY1W9lryFGunG1eBj
bro6IbFroD6NiJuCwwOcp6BR0dxAcoq1p9zkV9IMxxoGhmc5XPhcKsZ11v87K6J3
3CiryS1N1yRKEmfBsV/pmVXubxzWSRtZOW2vQ/OElphrZjUAx48Gy0p/VUFpAU8b
HoA84wVxEtp+9oFbBu/GCGhj5Zz+wNoqOkv4Pmi7ML2oapuyEvm4CPqSdA0rG0UV
bceK5EpTB4m7D8Alc8gXHcsUE2XuNdAXJl8NCouBMLXdDd/8ThotRYxqcTztEpeC
zuSD8/ig4EhBGzA5mMCTUvab5kzP2pFyiPSzgHNdwcLIEZKkqKm2pb+jxkHOO4sB
iOeKX3BnmpZjaPOWA5hzQB2glffYVcCmWwnP9HROOVxP88PtMlSQi73KF9bO2WCT
MN9QlIIsBAUMDGf+/CbdQtcvSTl83DT6aexg4/OhmIhGG+2k83eYy7uZdSbhWQ5w
mdcLZesoA0RI4Osu5exadfNCbYPDHGsFjB2lH8uHp3AAm4p1KUP2PKlNeHxLZVlu
SL87OMMfn1C0mIEPC5/yUQmNepLP2bCMkVd6K90YGjjCIgkE8DA74sTejAiJMmG4
TcCDk7pipZgeY6eD3wo2SfdXta/T/5Z+YQtBmSRm9qsiQb82HKkXOO9L/5nIGEKm
7PJBSZyTmgol21whxssOKCBYnmOqQE5lePG9O/pNtQVg8aCpOur0L0G4ETQe8Sje
shIuHG3ytw8rdV1VHbfYGu80x1S3BRwOQuF+ypivPslT/P3fpFVKaXnTnQ2V89gb
zRGLH+IV/TntQ/kxuI3UH7YVT91uReMem0muw+woFlcG1oN5Jo3JlU0wDbJME7fR
NdTPGILgvbUlBDcwDc73rOESnLs8Yrv4dJASGOLzfvlzA5vEZZns2Wn6vljngL6W
kvTb+fg96NUBvCkZ5tLJHjOCxT2nB/Y4Fu7zN7a/IaFSPjcZzDl5chH3SCIhVVS2
LDvrNPqslabqgoav0NnWdDyLXl/vaqgVvxrc998USAKI3m7sxV4a56WoChvacHJI
fevBpBbpm9PTO1nENXykQrQ/r0Gt0rojNWNm/ha4DSwjZtpBlzKiO4oPIFcniLXN
Aupol/JFReegRKu6NmvXJBICwdvtD7n7tb9Q03wo/rdDbzfl6F/JDn/nOOFyfhwg
ZswVSXJ1o91bUqvLU1bxTanPNxjgNse/DoJBJvySmQW2AOc8vKUEGqNMT/9zezCk
FT2OPNPog6FEX0vcJACPpTuCCMpvAgMUWTXi+xYI1Ek7SHd7TJatPO3Cx7EPj2Ue
7hN5W3KkWLAefu2JBkuENRDYbUvnjvf4BbQps4PbjjwRLhabFKwq/EtJRUVMiNWh
oQetuuqzqAiI5g+7Az6CIm2fszZA/jrrDMgxdDO1scIomShT4Suo2dNqn331hUUV
iNfR9h6jaaXPovs+YJ0gYJD8zdwl2TT7xE2HismeBfR/PNHk0fhTjWPbOyEZfZ0h
+yIE0BYqUE+o5pdFX8VbrjQhafJ/NosqYxLlly8myWysvfiVdyA8Wp4V2pFT0z2w
VeKJ7xPEd0+26hiHfs8Ze8FCoTJvUH/MokkuSkBwvO0ujgOyXX4JgLXJMpg+tnOA
QNzyBu9Rw4pAiMK0movo7PHw+TbOqiWsXV2CbIp92BYNSC9I3eKsVMaVx1gxh7y6
nsCWg+Nr3Lav81qO/YfnlkmALjf9ypnNKeiPg0UyDJ3grshnNU3gq1oz4c1g8w6D
wF/f0XCNUQTe9O8s4w8Vttq9W4Uj4hLVgFCFYffovsmpA9qp94Hp7sY14aWyI7hX
GSxP08OyxV+Ya2sXvB/UAyZ2WVqi9MFDlCaiTW88vPALMZ5RgL8bToGYJ+LRL33B
gPlNRkAFtl7kemJnEB7cFdhg6hrkb82qZVv9/GCvVcViQMW4rLCzyBqTKuWASdDs
RbwAs+gnR8evk1QjJgS/AY4aPhX7IJZHy97X7QHINJfugDfyI/fmA2tXOTjG+5g/
/UsmB2Tr1DKrENbesQyyzVx+xntgKKr7uqBchGL+45oZzzJx1+SDPclsgWYhaBVG
IEpCBrI4qbiAkubNK4Om/W0+TrcXFccFdrxSzQiA7ojYu+Nl+OOpMPaabJqCVNei
lFr/tiSD94iHKiosRozt49K8oIAwHddVmsyVTvTE/m8QqoPQzjSY/AMISsjLUe1/
8elDcuUkrQRpDhHBWl3JPxQXzg0tyjxN5XOs5/PcKKxrmaOhaYGSP39VPHk33lJy
yvDp149i2ty3WNNzgNA6lnyD9hMWsso5E9ozkoLLtUdB6sxhGC0ghrJSEn2oFZQD
v5k30Io9x8jI3VSSkCh255mEyAdOIF66/n4gUrViqNsLeNnFnlMs2kdRsaTd1fOu
aKmwVgLICVrOYDrJMrYP5X1ogWgHTNEelh7nz5jOIrhdafAsFfckdmTPsSFtejeC
mNLgx5PPE8ZlI0QJzd51FqLsdpc3CnM7DwDYeSoqlgr96IkorRFuMhA932r5G1H+
3DcInoBv69tcU4L6XbvBuMF+JJFlcRQQDebaujubKLatkKQLkSzSPp067QvVgzDq
baK7VYtx2lN5dfUVfTEDypAJF2uS6oct1TlRXfQWqbkQTXX8ovNAGARSMWy6dN/W
tiWLraHVqgclF+iyJllXqjbi1NHzgSFivwCEGKJ8Ak0tCyPkNgcezO/rKO67yO0c
EqSqR2QLGxGWSZVLi8TdW+LxRpbzX6I3ZqUXpiwMXhYkQFVwWDMrJGvWBN5hzPJq
C1HSufh0SRk5zpRDnBqWm4t900Q14iqKlqcAGn5nKjnUl3CwGc4YzirXu5oVSChs
MWPVzw51F6V/jx2sCD1+6NJQjySMCv3GaPbwXhMvv6s5dOQEkNfoqCKxw2AK4JmZ
MWwZRd25x2zJATd7ZERUzIHhh8WALoepWHVOngme3/gss0QX2MZMV+aYJKDxl94+
kazSTnSfTGvIqc7bVV7yNCPzREtts7c6xT4wGom1m7Wtckfktks3fL4ttln02NjU
C/8i2AXk5p9lxvoOIvfZd0SeTzaNDIzhsZ26t5MQeF4kxy+hhN+/iNWlCZqLo+n9
HWWBOQd2ExnCc3/0T8ebAhMcoK9sbWxWI5qcbCAPgjELvrHRC3wiP5eGqmBM0aAw
Gz5qo9mKJxRZRk9FK3rRTb/FxeZU7dUDCZV9FtyEc837V/6UG8u4jG5SO2o0Oi5y
eCH+WLGpS46Qb2lwqObhK9hqL60U/PRlHW5NZHz9FRAkJbMKZvvw+fbZryFu4tGM
16hmkBBpuA/BMMUWWrb3jLulmEgsqpHeSUzK4KPnHErpTcfal5YYVQgkrFyaPijz
W/lpkrDhkaiOXUe5+v2cLreWP/H0nTC/SlzFs1Z1338Lrew8ss4joW9qhWoEdSMb
OejKWGR5/bSKnrAcTR4xLr+xAa/z3ds8jFqH0mA5Fx66ga2Yg9j4BA9KFntG5vxc
syep1QizJGalIiFA2vf2PtJ6hS3EchJx1lXDeu7gcED6EIdMR+wztQRSjOt45TN9
H1vGYNPoaZO+pTzT+W+TjeEsxDddgASnw8ZJLMKgFhTcpJ+Sv1YE3pttJzdI3UKT
QvIOKATqFV3X6fQwl13oYpyuSn/MzA/nNa2j+Zd0MRZGLGsDbthT24Q0NEUtbyOi
Tbo3Q3TC/GBt7umaSaUUwia+P0a4xBITJZ/Z1PSLRMCgHAi4mWItPt060zTParOw
jEljuB36WpCBRmPXthiwCJCKYuf5gelup9h2TMkkmTOSJsSvqr+lqwB0zjF7RNQD
WQhr+W8lKoibua1qfSsMw9HWrvLYXo0Qlb/WyjFQDltbiyA3RBif275DZTYL/JGJ
dmotfNmBBfuPCss3Xun+ZySowvMIq+vDm+SdG8QG069A+KcQGD6XPiU/++UapZRd
wYKnxLqp8qiEjAOrz7bhhMZS7TtpNUTz1gh+uA2xAXglDfdOB7gG4iCsWmTkPK6n
P+YYTBuXIoWyN4/mE+J76SRcIpk0W6UAUbCHGm6zOl8bdxdUK04PA0OgXrM+L510
LKNK7ekE7anBAEtmFy8qUVugQpqpM5ZU5ft5HEBS0NQk7lpinT+MxIwQxfjx+7V8
Jy/RJf4rXupF63k4ubFVyucjCxV7O5XxAXTQz9EA4Qr/lEFmDR+BEJYdL5jUSHBr
H0IUkDhbzphL0EFANWqUDJFRzc8jqDOV195S2T/1uKNbYHt7BtF07dYhg3KfVrRY
xQatxUS/f454AeS5r7p5y/p4DSTPdJIoIeqEGkmSuqNWB2Hji9WfetUslG4ZY/Hq
EEvRuZPedPcJHIn1QoV/nYHyXetflfuBRw2l3uHB9bD9oXf4Mw36JE6707FfhRO9
KPYsnCec2MuQuE3KbZnFZANAUt7MZHWyRMOUgJ9VnL+wmSYstwGFxvXiJIksn41K
lVzBlGCcuMkt7oWRL3gyqq8r7YxS/uAzH3QY1Y+QrHYpzWx8zOaoRcU0EPSTz5pZ
V5DamJ/PUB8ro8SSBM+1bLjdx4G0GEvT/MNDIkdUYItNzleXqNuIR7psx2MJLhWo
Uhr14G9qT04nZPewWAc95VRk3+tXJY0NAF4CkWtQaGr1LF5EHmsrrILqAU/p2fZ7
MgUcCBnQ6MPX8MFuBnLzcjzkgjpRpPbh2sBeXAhqPyL5YHsHANzQXmuA0rV1ixOs
uy17bj+qF/xd1jb0DH9byZT1Infok7aUIfNDlJprS07J0XgVxPt/eR1PvgNRJ1rK
xaw1v1UEE7MURsKnvdACWVYRvVK2jeOf00bUBZeNoVn4rG7Jkp+dc0Si3UVq9AJf
jNqQBkYRrxrKnUCM4r0/0YuHDKoHaR/LbRzVzWuNi2KhGWJkHmvRdebmjhTiwde3
gnh/jCSgxp1B0VQEt6j0Gv3i2426bSFmIjFemvBN+stw1UHk5rn6R0Q61Het+OtW
aShAIgr0vgjeinFEZPQebyDmvUia0xExwCge/ha+RNLGix8DDEK4t+k6mfN4vpNs
yWNciKJDzSBJkm/ONXisoFlmCyrJtS8QrVJ3MD9UNR/YLuvADlVITMjF1As4QkPl
c4/HGTQ801Id1kH8Hwuv27Yo61MXwdT/2M++RIKO1YpaAmtZhX2FmminNVMtLowZ
nebPqmn51zMm2mp0Bk1efywdiA4UkYd8+l3WIf8xq6GVrLywn2ywamLD/wWn+o7b
097G4eu06flF6sfgjxqB+piaC35J5aKfYgT6vM6q3voRBmUk0+ag04uw3XeE0eyz
JFgzcWOAqifSJacoihRDRDwlKTsmhSXPie4DjBb4rY0KJfAaxMrHdP/P/kI1JJit
QTQNh1x8BYYnP+fFf2atpmQ1VX65PZOuZoiLSbqNeaa2exCLPojSsZqnxBQtQk5B
m5AsH2PVwBXXk5QRdZKYveTbDHbWSLF827DbiZBZV6HMBYI0aQvqrj2e5cqTI/ll
az37hb8bj3vO4622PguGAvWUoOmmqb/bHv8z87UJnXavvZzeM2NsFKlTw2cnS+Rp
tffSsOdhdist/W3ztAE+65+EIFVVYI2Jc/nWnJxN7WlabiNgLvpEAuml6tfhrLPY
k5NqCqoIVCAhGW4gWTOLnFxtWHGjz1w8MH6jW/bloOqbkZdRnX3JsInMqhMjSOxH
Eraqb75oOMjnOnlVaH+67MT/UgNjsIIRL6vQCvC8bdzQYjYJWYfEoqLfy4NwvYBj
PQnECTd1sh+RluhpC64yHBrDYxDLnv9LumD35Z3s04R/bXhAC7fNkbFs4EXQ9fpQ
dAOoTWm//u5Hum41ozVqZEoEem7aEfzE2ub5Y+3b0CHYwes+aBrfc6gFlCLeJ5dv
NvlPcjAfZlwlxglkZmNHVSf6xHYWzCUa77HTSeF6I5XCfFwIaRkYZ7fBbqF4h9pr
yvzOw50VySIxq1hKjmqOzxy1mIgfkVn9RNOY1T0kKCxltfGG2ovAsx2YgG6VcgWd
ShwvNj7hpzHdtB3t0WQMcWyPsgHryZEInXeaLyZ6CGNEEveqfgIxzpm4UJ8X4DKM
jH4e3jrZFou51YQwEWxt/VypaTY0fEWN5GDAtmVEaVARhmt1/aeTLx9nBnpYTKzM
ksF15jKw3Os/lCbs9p1yIi4T5AackpU1pQAWSGXxfxyVqDbDFZhT9+em3B4pD2VW
BgLfOc4z91Cir6W4Ip2hhDOCAK1XC7t/DEaRhMSlrKgqXVjS0Wf6sqZUpZHwyMBh
iIxB6wPYyNGtPVF6NgzHUntugnvOqXaa9zZxmqgF7kvFyoCOg/i4tA7yBi0KcSCe
WmY5og2Vp6tjL2x1Q6vsLbp8Mkwvzz/PRBDBZbd9VnmKMKa56fOE6FQMI7SQotjV
SAayMvqUZF8rUVU1YwNcHnbNjCDFXW6U9VJsVE9H7CY9nLMJ9bYLBHXBVFe+o5VF
CCWjogrgyO4QnCgJl+fBISC9+/guG/rC/dj3+ODnv6JtK+WilcxUSpDRgECJma42
qMw62IQI+bFDHnudhZtEgIKszX3ruLasm+hP6ClrVBtc+XUaC5YUAI6Z9B8Cnhrx
kRIEcnhyhMEUnmat0ghneyV/Wj10Ym0PbeVF3uuU9frr/wP6SzDmkBT9ozVpWL/d
yIQSdjmENsAzTkW+y0OViloiGS/rlaFg2AzeQT/NlbNPszPIYmOwDglWeaJYE1Zp
ewcdI6nQxCRUmEqFBZpGwyjvWbYOP5lTdMjj4jbd3Q3NmnZeM2OnNUXEYGbUbXd0
dkZ1oryufoS391ntbnCrTn8T2ja10oUH20LdwU37uv5kFsesK0pBFu+ge7PisV1B
XKLoWD5uhTYMZ2ehJqYVMtZ+9j7vVy6xjEIbykteG3ZlGc+kcwNm+4BexZiD9qAB
/0P4yHR+QyyhF3D6avLgv3/CWVa+/rIBx0g3ztuT6QNq/SPPGO42aU0aNJXFBWye
gA7f7bIS35KOZJEhEO2Xkq8/NnxUuLoj0qpintdTEGRcZVS6mEQA5q9gLxujuDDt
Rntm3OYg9S/Z+3jvuqLAhZ1GcD1G5CU6uMBSjfAyyujXNbOwzxK/VTJijCFZksGJ
zclox9LEUKTHJU4HHUgyRPuEIFVHdswvk+S7aspDwV4L/oOHfYjPtw4wHMe7A5BM
64cQqjgvmQk0jAFsTvKFcZiRiJuJW29rmUSxiOo8CSi7T0g20Ynbdjh2YuMrMRrr
HB4RL5mMmRtqc8pvnPKWOz6kkxaBqrmZcS6HwBGAOnSSXMIZKdSrWPDt7onbPlnX
+QGyhT8u6a5JIgDQznZJES9Tz7iqViatKF7SFQ9tKm/Jp8+KRAs2v5gU66F9mzc8
5wRkdRO07hg1LfAGs9mGI1T7Q/17li4RIu5kLcLrTfWXt68oXlAODLN3yYULnoku
+1bBzttehDS02YQYf1nnehrX+VY6ZdO44SS1XK84HUWSeBkqXsxuQrJUbctY/PEN
X5FXmjX2PwT8bngIObq0/x2u8hWE5RB+XGHIkTqPO+CmsnskhGuYOb80KT320R3T
zETCIqwmdq4Waq7A91Q4EWcIuvaTOzI8tGsaW7+yR9GRW5qC/MlMoidb2HNW1mnN
uXkPERr1NapqxNiIRBH9XaTfEmhDDL7/V5LgFIR4+uAmvKSRzswzzmPCQZaCSzri
B8S2mOviL/B1Bha8IIJWzeyfbTnHDKSrG46PtmHC8Jn+je29G/emBKjRR6MCVrDT
93HykdxGKo/WK7iCRRFcjxvtjiQHlKI3YqNhkXTfzSiq/b2in7r7s1P/dF0xxZZb
Z8TOAKz4fbUvlvP15PCvI/t61mfvGKORuEN+DBd7ApdT1d6V0zphPcozU49P1KWy
Bo3xtNKX5LJjzJSvwd/+Zr8fshSejs762FeYCBVfI1LgVqBPsTgcrOn3CBgDMdMC
+0MvWkucW9yesC7yYqZK7flsyrcTjviULF/xWknQHMbqeXtA28aal2l7fZufl10o
iKFmSzGrXyBO58D5w0786pqouZG7Q5WUdrPsbYcRFVlPQTB6QC/6BQEnB+LH+LWS
b9wKXtwPvniM1XhFnnH8dgQSrBqfEN0rC4kZWgJivdldmaBp5KmqPB8PsQnJ5D2b
tS5mNBprcEQRULiPDCcpIPmbiBFhbXF1klKgh+NPuYwvh5xZqPC0gn7HOJgHdWuG
6o73816OUnuj1aVBOwckANhFly5tw8bnvykCXfn3kdC+1K2tTkV4c1u3epGTUCq+
GUjHjUzYw9xVOgIrrfGXbcMS7tAEziuGu976mrIe+oBXUy5t1IotsJv3xq3a8jqX
aKSMV/PlYzGz9S1VQMBjCs+Gw96tgqYUXOZSbZ9CAkV+X+IeHQE1fbG51hQ2kCM2
oAzT5yv+aurOSEImqHeHI3gOlcYLE2MzzxBe2P+BKxWQtcgV07r8OR+UHEs3Ylgt
dcXUlJaiLtjJN5VIrpWjv++p6jdNTVrPZKmU0xlAh3aNlJL7pmeyNnvK0GM0yr+j
li6cHmXr85mcpWNaeSD+SfEMoSxL3mFJrIPeY7INq4/PiM3+XCFPVf3exaJiANjw
68NL/yZ/exM7qAeoSPib/fZ24SENTUgyOAYCt2JrgXrIn+mLbepfKO8d+troq5Gi
T487tCUa0+IELKpGanRdpHvX8h/i8guYnFk+9QhYDWwNQXNETKNaAww+YVCJWH2d

`pragma protect end_protected
