// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dWjBQ6GoMDzCKLUsa5ATyqt+tVT4OkWJhDdYb0sT9/b1wbrlRA5EWGQqqAXo
vMwj/Y1XTqc4xcTZxJySktCZA7tEkSNxe+A/8iJWhA26IpFvNUSToO2JYgqn
+wXHGfd5k0y/nYhU2QrjUwCRWFHvY1JrObvBObd0JJtlXMYgenXWyudNG7Rb
sK5b2vgWJ9w+7aPqFa1dK9LScRe0nryr59Z1O8faejPCn2/BkLfILbcMy7fN
n6Vimo3mgVQ3xmMVY/B08l2lN+RFOG2Lh+6snSwheQOIpytJeZpXqIyLCl2B
7Dr/djSC9zAhQmy4iagGCNdB69JwuinylloYSOAAXg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kWSu/XHIdn152/2uui5sbCaq3lV7G9OKeA6dCi1Zp0SdVWWXwxcYhQ8M+ARx
+hr9W0RZwvsEtMvBsWua8fLmdGubRJFGhY7Mp77nDSI+A442RK3bf3GtI7Hj
ZO6I3qB3QSZacmYTU/LHJIn4nh692xvohnh+7tpf9ljduSHlxxRB6VqLD8EK
LFoikhokrHSdeSL3a99Ddh8GdfZEjLC5U8Yp+p+yzTqYlViqrq/9dhkc3LVW
6uKu4ThavIRAjkIjGwDoxNq/R21UwQtZ9WXSKM+uGQUEF/KfQJiKUnfQB6Bl
2oEubdh48biuD/zyp2wItmnQICmWPblqb7d6d4N/PQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bkk1K5cpMVeGuF6tED0fmpDZz2hYX3ids3LoIK/f0ZzuYfiBfS1vLEGRsa25
3qSb285EBTW0HF7TVF8NRfZdovJM+MtysQMQKxHjezOnWLl7+Fuj99oH7xwq
b8uOlS01VIMcw3O24KTBmIqZwmIDuc8OfmJSvfR+y7Qt5yotMz1cTTquvi2/
G/E/TdmZmKyxLzRd6NzNADWSN7sHuApNMKmLkvrAr+S1h4yfuDTVhWX5Afld
jCVclyKuzl2/KZoSn8IngEtwdEkVnQUBSUPbwapl/TyiJo8fnrFkyP2Kq0mc
HhoqVVDZgQKX7Uv8N8swPYKKDSPKszFOAJ+RdRwiKw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
haacZj4cpeVsZj4FiE70YvAY2bLii07Q5H+yijGsSl/YqXzWeMbMmd9eagqu
S7Sybm27ZPfJ2V/rrmOjHmhIxHqAosHimb7Io7ZLfdzCLQPJ1ufmLLC84ZgG
AyjjpvFzMqfXcIL+CHnTAYxyQKyG0e2l+ky3Yo+vLo/kVfouENs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bRUPDWxxBgSsfsuym5t8y9ca3haaBWzIeXdocxGGPFMQ7nrwzmmPXHWnbRTu
iC9IovBuh2ILlJOxAtx/fimuF1kw5oUmeArQO/Z6y2PEfADXb/Q9aayvWssl
Vy5iPEMqUw3xDCg4YOJi2R1H/twDXfuP8zcMtcEINVHwPoIr8FIhCK7Bj1RV
i/BAab7eSL8TpjnYzOU6HT9LmVsj+IudjSj5iBGTnCTo2imE/i/jIlMFM+Gb
3YvoDfyMLCi84/f30P4Sfn6iXergRPEchOWx4OJdEUAzumBpzlpvNeOUCbmn
z77tmKGQyRi47w8bXj2l3wCn7bFXxsVp40QfZz/4/EjcyZ6eyJULwrxv8ycS
NX3TLAHnsAanHyGWsCP2fuPW+dnZv3s+xFvfGhbmGPMbgD255/4Brnr7316n
32ibncoos7SMj6s/EfIfVY0xsW9/tDFsKnjFeUXr9eO/5Tttq4DXkZ14PfM9
YK6sMz3kD3/tZ0D+aqbBiTmyy0gYZFYk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G4gnqv9u08eLNbXTx+D5vwJvhXWAegfcwcfgdVGBVra0jf3lQstaj/5peh+g
21l+JeE2xH6adPKiJiihQ8z5/j3QapV9hFgHjzsjqoltBvnFOzhpKnJuOBYg
a5DUj9LEqT2gnUPNkSffoEj/G09G9IVzGO9g2/HM12AQp3ivSLA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tlkaloZEZsoht5QXAXPdxKPNe1h5ixwrDQJUPkBgH19f3hLAQ8At1SZxkhZU
boI/XkMqtXWG3vcgyAmR8RMwKEsSlz8TRmAVir+RruBnI41ifJutpOaNmGvK
Fuw3wtx27yBBY7Nb120qq0a8J58Cy7gkRVggttg5dgQhfp9FOWM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
G6uPzuVpMe7fZUCVMklyRl1+/ADRCqvkuJ4a0sMyXAlP7xHJOexpvDHADPNm
w1ySnbzx+inpkU+4V4qcxFOsTzeMBP2FyaKs5Wq0Uuth9GeKL7WMo2XMZuWo
3nT/DKUgX5/GF9YiW6A3eoQnGbnyX8lSlQO6q/wPiwQlmazAom3B2KFpXOAH
j5bZb7s4ipun+pUDO6haCZyWiLOyYxMhCIjIXft/QyTlqC4B+6pJmy1GsgNj
SRnHPoR9hWBIAOW6zAAJp2fpJZ5UGRM8d+qbbLL1V1m4XhDDmU+W2RfMD7uv
arajTAcf2BDmrIQLFOM3uEqLY+pek67P1zsfbml7nann24lkrtq+Z5xLXa0R
WoOXrpcP0jNiH1keTclmqZBigsT0v69sj2YpCjmjsuszmyqZZ+ax0hjBdnQ+
oAxHwk4jo7uUbqG3OugeUlaGmFqfqDVoVdYzEYucLhIDajaiQBNo6T3oP4e4
67C8I+pNxjbpjdrgo2GJ/b9oddh15ZbOU1+Z9hkz76CW4Sr2KpfqCJVTb5tG
fBSW1wgaKVzJ5KbNouegTeBHx3sBIKXCvRob2UubYFv7Of5YSi9rL5HkM0Db
bEwGakS6y8ZxFAqOtTARelpvq1FgHWIpmCNWlp1w0qe2mJfdtay5HgBrfcYd
pwsSjXRMQemehJ4kS7SrTOc1LJeljkDhnOStphsPXd7YYMCEZxQtUxEpDse0
rOiPtrbWWqKi7tGIusBtx/LBhR9GsEjSgYN5UQf3BKhW/onvjMENHFwRPKqF
uOFJTGJPYrq7eNdy2IIwcVWSh8BrOmsaAqvs2k50EpVskaRhRkhOR6XyKaR9
14s63CqvRDR2JMGEPOLH4BhyQseFn0kufuD/Hr4MgTAmaHimBiRkGVyy/MN8
+xngo7eu2AnTJalOEoedroRE58fUWbDfZqt9UMVo7IezSbwqOnFjjyzg0Sfi
OccUVTSAFpa8Rr4GRHZ2ds/jQ1virPyziDDzrqDPxZndphNuvFz7JI/OWi3T
a3QOV4UcRPSDOPQoIOXIQ9s3VauF9hdT7D3mAA3z0Te3kj8IX5b1d7KxhDUh
LgQysFiFaOcp7atlg0Xw02iOeeErjdqaUk9q3BxUsdc0U9OgqbE7tGsXHcgD
a+vSJGGKfzz3ES+82dwbmInS3W8a4xKua6lYTW5xUrLixiwHwEyu/IzaLg/0
MEj9+YnbdLiPmMQJmKD26E2m8tNjmelbiCNPcolh9WTa6hJpuWLQ+sY+3Mug
ChAjfDcZ8fCA06/naBh0wwfPJtmUA0hEqLlmlAemQfnrx3mjYvPipFRoiMpX
wpWJGdb5WhatgDZ0uiCm+zpbH3sID1v0MVfZiVt9bS2bk98YUZB6jJP5Iw4y
afKLwoU4tfZ4vewttrzGcoLqljl8AII6uRHXsW1VQFfDwx4BgJ44R8PjBMa2
/8Yo/3K2TOpW8asx6N3mwmEmgEas4HtkP/8mhviEbdfLOwK7t68/uZ0f4WW+
A/lfQmBApbMPUWy5jFF0lcC6e7+GVx7FAYDAT0mETpv1N86L6T8tI6hCoQc9
Vy4DuJupksBQtYe1/hjQSfYKFbS3bVpRTqqKhKtyzDs/GwxxU6fv2yvHfHex
sOmy1u+ZoEv6osDrk1s6ysFGL0IxTAUmk4ETid0pgh1ZiLlCKQWS8CGdLYbu
M+Ev0Ff+KqSSm4DYPsVnwkHZ1TVuU1QuJXvTlHYbTX+8GFjqRTpMk+IALAj6
iLp/A1Qa5Q==

`pragma protect end_protected
