// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dkh45VyUsByGHi07keTRPWAz44PYdooHsUBsBDt3GF4magQ+hDQh2N+CqIlN
hUrz1F9JxACijTshrmI91lJE0Esbh96z3SWXh7minmxQwCUFvAMcmBdhmhg7
TaeVju4A/zIuaIIc7YpjBw5B+l1RvJMSOgDfB9MpnETnyLoTrt/FxTlr8zI0
3wU78EUhmmS9I1diTBPDpEh7JFPpgaIwEbZhOw9KDZqGUQMvyKhr2nRKTwe3
P2gtOtBC1vl4DMiBb/o2EsJEL9AHbtyhW7nuz4I2rxOGUKSvFBfxsHgzw2Zh
qMiy2IiSKdUu1eJHUPdQRI5pD2eGmGCkKs1Cj/e2hQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gT3DAqUg4FI81FRXgyYGowacrH510rRsJyvQPBEUq95lH19hItWFMBuHmHPk
XfhJeMK7GIZYcBts5ZwRjg2gBmcjY69W7x3nSxmHP2Jq/Mzcf/tKfVIeam7x
MIltaZIR1nk4DFurw5QkcdaN/bBwNv3y6hFpuf/3XFVvkFjVilWZM7+NTOmh
BWTv7ok/BuXYE5fhqdgYrKH0lDQK97sN+cTfoMBfSM8h7U3+2NKdn+M43ybj
GPULZtaMI5SOYOw7qz7xoaLFGRqm0K4gIb4aFxnHbcu5+4lq19DwqAVdFYYO
CbJdjVSw1cKEzBoas+xyvmB5RWm73KTqCtX0C5IWvA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UshpWtK6PIPDDFBfKiXL/Z63Zam4B+pfd7rDvJXilq4MNNMvjcNVNtD4ueQC
M38nphRyiIcilszygOucToJYOd0pbCrx9YiskNTep/TEm21+wfxrhdixzUi9
uhrMSN4ArhQuGeUr2w5uYGi6+wDm1l+2l74QXQw6/SLwsaWxsQStcJnN+CfN
RHUVYJ0HXDk1WQID8oVgVod1dEQn9yclDldG+kux8j2mfKtgsMnG1jyXMvXj
BjMY9piycEZiIlQ58ia7NMFAUPG7jXERMBtBldCas2vcUgUDar1Ow5HNQBF+
agJ/bfXcF5wiuJPjN07SXH2gXbMH5tXP1ZC6aeKxHw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m4mHNM3fYqvFlbcvT5C7etrCblGjJ7WYS9p688lBDvf51E2LAmmNBcnc4M96
WoA2Q1uvR+x/45dFIDJZ3HbqvAHJ+YH5RnFGdUkf2EnpW5Ukq3T+ss/aTPt2
qX4AGdfKyRTs0odIcGmj1FKXfAOMS0vWBhetyGlFoqF8UgYdRVA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lzN6C6CZrgTnLqxg/kKxaiPSxmaGMCWhVff4NbE3tNCAcw1cPcBN/5oCPSGO
pr2sHVezDkRFMwjh8EIOua4A522C0631qStUwUg9urcRutqvtgfRzGlI4vp2
oWlFKoIEei/zxXPuTa6P1kCo/zDhl+WXZliVEZeegH3bWoRjkldeNYAgoibM
mypPHlhSK4VxA4Ge1u3QwAJU92b6wmMIbpo0u/V91dVAvPRgzXzI/kmy0PYH
QD4WwogFXUgm8yKcsZp2bkjuo8gHsQj/hJwNUTjGIhmZD4mDSx5ZJdyx1cxw
mckktCLNDwfAHRvzV/A+9KS24UOiJX9LSk6Vt9WZ6UldiRFHxVUL76MhANFX
UN+l7pz3mrOZ7tPpPkkmu7bTs0N/3qfX2W8xjAvODz/D23toeIAPb8vlCzfE
KoHLwWM1IXvKNbTpawngkmB8PAG2IQDYk7OBDzTT1lOk/x0oU5Jbm1wYNUkO
QAYyDBvkrj12mo+xb1aRZm2wkMyUJVMh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nFlRhmB6IkzTEnpNgjSY8iNxjznAV6tIvgse1tfeMdmu17o3kV1wbZ7fmdCc
vkNbR7faTcPnEzpoD6aTv5DZRutkVDmFxgpxAg9nnY8r2o5sOrFGbETa+w2x
jzRX2X/gPt+GSNv/E3551wmVk046teXJnjkEbAlUzMqcANdtQZY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YujyjBGkqZFMlmF5h0rOjtRR5bdclIhEoaHX0FOEXXW/RILDFXQueGInCuqE
VF7GukaUjnC5BxEL8v4Mo+wdG+RA+/AK0rxSDO1CVdSr4WCQWExGO3WBkUFk
aKDQGFsZWZLeLySRNDgIjkUBXFqzJiNXcuAnO35vHz0NMq3LKQM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7584)
`pragma protect data_block
2aKXHS5iL0VHgi8oAifEJ0mMJibznJFDGeY/SoOLrwUorW6CsomuwEgeYsTc
JqOD2W0RVrJq87+M/TtsILI3luOVcfKDpOC24tb+JvdNo/Kwz7Q1QR4tSEs5
rkJ9GFU1l+3e8WqsY2dMHOQIEsqOY5BgVNXrWhisgf5rx+Etr+MJRiZBiB4F
jrpSvgp/pWziJ77rIQmIfTR+Jscw4LoXxHcwqzEzTvO5c6cvJ3qHxquqHkGK
cZBneiDx8b8M5mC+7syAivIPvlg0SzkwReSUjtUR2JhuhgnuypiRBt4aQw7s
aTpr4C61wAZMPiyJ/YNXxvBLd0ULBIVKMnk5LEuiQ7b1mu1nA7UjyEG82AdI
ppUS2OZ7XpzD+GBbZutChZjmMnsjVugN4uHMiM2IMbHuuSKCEo9XwCCjOalX
DheyKDaLFS/4fPDVXDB6F2YO1AYmX/SJz4znyupe0RQNmuQlwZJKxEra3OyH
//CtZSstQriS9gZvHIkodFSQRK3ZeidTonD2Q3WVXBIoACv1U50fj6XlEoFd
oVx+ZH5mDRK+TuqEY15Oo7HD8vqhVh14Ls1akolW+NY7zEj040OZTj1X9kVJ
HiBeM+3PE7i2brTBa6AuUm2WwfeSzxgg7LK7RuVC5dDBqVD7p3GWIcRgzHyo
mAAmCMumzfm2Jk/Fnze62t4OSj8eRXYFdXL/3iRmDJhXk6A99GdWz4Cxlvau
IHkTsmTEKbjgExGihl3fZQCBY1FgMMCp2Ns5pj0+odjJIkm2G9lXBgS1vj1n
SyZBu4LVIPVX0QMAmxnKZUHKXISaLiO5XSgs1RTXsn1ZrGj03vXVYCcSdR8F
5jY7xkEfR6VaBFx1nhxSCgvBvdXsFA4JwDiSFcCgnA8jDTVVWTMJowljMiCU
DjrqTE6QSi34c3hk6nlb6PB9jU8L2tLKYdqFpZNEmDt1qSd4qbVn3B8Zf7tM
1w/5KWLampjVJMkrArNlRwPir6tqSPqXY8d8CLxt7iPshz5jPyghLZMVJEvh
n7opDdtf+lVi2fAj6ZUMFb4c1eH+9YQ4XpS41DkJTNpR8RiacQ77z+N6yAGm
MrQMt7Q4qqKbDreJ3yOsOBu3Ucc/8PGaoPoVM2dYTzVIyQJqizAk2vxCSwyP
Ye7BaaNeJys4Ok/64Kkdsb55h4Ys6LUgwYt/ge6cF6Cf4MCOhhyJKdr38P6B
Y5t7rFA6HAvtoM4mR8ciec7uawweEGhtSwUFD3kZ/Ote1EKWxURMorJIU2ag
CaPv1aK4mrpGmUzOINzpbIqsot+L5y0NuGhV5KEF21kQKe3jPAxCGU906raL
CX9hviJ6/kAfgZ+RG5BN9NSHHSdlauh7Lw9nx+kbnQ5seigMcgAIQ4Uz4v2c
r04nWo9CmCuVwC2Uva1iF+j7tc4hwZm3NXdl8g/2sztcObxPN2gp08rnVbaY
b8cND6nBoMp1BgPG6zkDBEz+5qYQfGmDzGlpJqPt8/8g0CnBebD2fjdaNfIp
lZyVahd1x9znkKGzY2q3un7axh7zXUrE65RSNbC4GcikvS/KQ5NThTy6g1Uc
9XPY0nWqa8o3pN/uyiIyE9xzmqxFeDbq2ujYbf5WZSoYAGcYZ+6fZd1RUw+t
YvUto/5URRVjfrNMTK30jgI8zQzhGBjh2mKNRDHTSTQbllTPPxymj4d4BC3U
JaKXk+0RSrRvxgeYLEDTm99v/r2TNkxoixddVbv7I/ps8V3abwQKkSVIK7BQ
CCU1gdrWs4YeY5RuSvetNbvJEhh38jLMDlJx8xhv4oq7bzhf28JJYIYZwf8J
8U4/rTIIbh/9nDS2pStIYcnfGnzjwFUL4wUzYVoK8TEqOjnuKPt7bkfJIWFY
1MFwQxp4Ayink6OKbP+/tHUufIwn82HEXAi/FNupGPFS7Q6duGueBP978ZRK
hx5W8frUYu9mrSJ3zI5ihPkv0nCiVgElfPMgP8z2/thACRdmtLo7XiLmaMFg
wLGi0FvYPMdiNXcp062T9aRS/qdqpmxU5CeVSgKuZPAOvB/Fkbhv0a6mIEAF
/1mFc3zVq+igRYBtkEEczPXJO4sILX3GlshAzOy9crqSCdF0bHLIxnQ5Mc3Q
MWl9eOXJptf9xMHLYjAykkYNjLJopyMfwaJwqExMO2Mj1VOUGej4P5Y8HTVh
bk2ORrw6HZSOMdoFe8x28fFGR8IkMGh3Za9wqx4RT+flVBeeM5ag7+24Hng/
vJIqElLwyFFv+LHf9ZOdIwTiF8Bg2bfFqFLH0SoZ8y7aGUAhKy9T7hdx+vG/
ghCxGFBnXf1TjNdXR1P3YWIC6+Qbgmx0sJmJnXQGjHfjdlCEqHNiwieDoqAN
RBbAolgOHIzCqqJpVb4+n0ZJ95mCn+ooRMUiOyePN3Cpt0hitqIfhJmCP2TR
Tt/l3bSO+1KHJWfFMJjX2lyd6FRaRvcOXn2+FY+HAqfGb42FVYzOBl3KUjTM
SFnWCAd9vliGGxvPDJh+EAj8YVjZAW/tR+kbXmXJlXXunpVHxMJhmwhfR0f1
O9C0ac18Qa2Ilhvrzqj4Euv60/A6bcVAi3dZLMCv0gtto3PTeP0ioqxqLhBH
endiEMrBoNZXDzV36T1rFFfUBRITTUWjACQd5htsYoMsC8F/im1wgN6oTl59
MS6bbF+zIW62Gl5oFuah9EAZAsYv/iKzdopXi0DCw6aFRlWChCMtlbEXC8Yr
yOZMQUTWchtfBoWKD+cqzgkh7XNw1fnchX4l+LBI+nj/J5NfZCeBKDxYB2ci
iqolKSt7Zpx3yR2Kz165i3IqMGsPwht/AQNnzjsUsaGurJggkLjPADMP9JSD
MHHkfVE4SRbXZz2SFEU+5Xx3rbAbuTFSy1+IxGmuXpeZJkFMlVVDNE/3AOMG
1F+7c89be5npQQ/81BNpBnv33cq5uCK7EqSgrRbTIDsn4YU/LKKI8qcaiUOz
K3kDxLBwmL2xSIW1v+VO3ZWv4kvUxamGbFgTKeCkXAfzhGWdFzP18ftHq5V+
E+E38wbcXcggR2TQwoqevQTdF/FSH+CEZ0qPJ/gsjXLRm+OZoZcB+pX1TeNW
36ZMMabRwGsl9lRGo5SJyzUkdX/pobFy7I5QL8G1ljChvXQwlT93u3VKwnTC
aCWj+mnVKoRj1A0D29pnnHIZfX3wlpAZSAetxpP32jW8iJG8eqfeaqtVdCJs
6d7hfeuJ1nW5SdQkLNZjgmZBNQy0wnxPn060mSB5mW2Q6E4XE2w2nRSj7V57
UWjhFXIBOW8H8ChGlObF3sDJJTRO9ajSsVgPuDem66KZdUub5qe8ah8beVxI
YQfZTGOMXj/HonealLakiERzzVPp2ZmPTPWH9kl6w//NEGs2p2F6/KWA7gP+
17YOn0q/wnbD0+/NOEqQRxlGk6Y/l1cwnEDejLxkfOcrL6Go9LgrdoJyuOuV
HZPS7cgiUZMdSjAyWLIwFOFDajnMTw+m/FBGUQKz5ucC0EvipYfULuUVpX5r
hGjfCAPufkacI0QgY1I3xwRQIlygOiCvldGHXk5siC7Vm1gTOMNGBxx6TBGZ
JodSatqwNT2/FjTzapn7g9YLQ5t4MGRQ7DrnI4i6R4S0YrZL73rCQku0qnI2
DvS4pThKwYonioQ/nAgsnK4uVW5k+7l/2+pgrcUlpxjMFtlyrfyqBkv9uxsA
8hEslJJol4iKRGRuurRXPPJf3UiDb5G91+7R6742+NjssnFOUfMZATT3OUsA
R8FzAkRUn+qVNGZiKbgAPiTH9nkG7faAK57edJ3MB/5sd9999gd68ueXI1fZ
GbzIC76h6aoAUtjqtjNclhO9KXybMKpCajIjDF5dlFA/CAcmIxMpMU1KAs5d
Vmq0PAKFNZ2xYO52456+RmW7wquYy6CWSPVEuglZZlj3MpyuGGPWU5xyqfWH
DcSnD+5fmr1ywCKfqUQL53hPigfsOaS+SYHta9vCFbEult2OTX7M49lR9fts
iY8kkNQP37eSJ2i6Dip8ddNXQKBR2Z3Kt7wXix72FHSXd0wLyd/DP2rvavkW
5JUfuYTVidFxYZuWvZscAWjc9NpmTQjLdU6taWFxOZe8R9w872WwbRWOPko0
muUM+AnnXMGpMXnbXZLQmmR8XqjSCV7RumLXoIIWzVTEpIkBVniL/l+0afCY
AhhqDWjOCogR2rKwpmHKFHT8R4tUaQxhw+KS5TmK9bTw+cAhHlm5H/BuXRye
zXZUQoDmqpIus99kHZZXTHzAvhSOQCRTA985ezanH/0r8sOLYrinCLLSE8hA
vN6UsGFirlpRIGDwrt5cGk6nMn4koSxygw56B83ilQD+AsK28jPlawUePAqL
NRJLj0ZquUABqMZSgxK4kWeu/GymASLivNjoJ5KWF2EgmyBMbFjpL0wRUBKW
v+sNP1WJlfi/3BXjboZQ9RPB6UA4zl5Ba/pJMeie6btK7lsOefMTtgvSeBUg
9VlNEOAmMqL8+XeuXGK0UFx+0QMUAXaYr420DHaKrLupo7xQJwHCM4q+skOZ
PZw/f/8ACGiGFXJ3jG7PI35SHzsptNYsR+S46v7AcmgYmXa7kfuEzZgP0PEo
j+om/Vr90C0KpwD2555/3U2Kd8GTPX62M65PY2azkg9jdgeB4TOYKjcYV8DU
J2oO64NbHNCa0BZAVRx2DAvA4UNqTUai+RHwJuVQfRikLpfoiGskr9vq+A0a
NjdyaVOH0qFcBDrtwuxnolUucd4S+izH+NgUF1RbgpZsn4v6YLhl8/GsRFSh
AN9VXCyycfR0pB+z5dwRegori73BXolHiCKeH3hAXLWzLcI+9Fc7oP7cVNZC
iz4yywcX9wQxJhDYN2SDdb9hBMqL9gwwXuEyeB9iACvcyPC6ep+OvASOKjrY
mfDUDwvStAe5KgoMSCiHFvqEXtIPJJb7E294i3L0zFGNwpu8GFd3SFfGSAbz
4z9ONGCr1sAw231cpleCuHcRGQ5CUYvGZADbatIZXEiEMMj/bqeRDNj7wX9w
Q1pxul1RKwmaBRbAtgxx7F62LgD6ILni1v+tONiQBk2AT2T+BQK1bNgiCOp/
tWPpfDhtjLZYg+RY1IRjxCXsIaM26odf6P0+MRgUE+aLo4iOvWpMA3TrOIA2
+DhnYSiewFNa70yH0ZrRzVG2cSnnn00hW558K8qnwYF5Bnx0Sjrwi0Hiqr3L
Q6lkIOQfsot7Gp9FUHKckLZIApdc9Lw5zL9S4ucnU7i8yyeg26WrLwNeIZ1h
ZIR3kCbfrhHulmFtzE/lgAQrMa+dgdTGEsB1KlFLtC1zDdn+mR2eZ/g5ry2i
zJ0UAc1E9a+zERPEBK/yaf6eZWTRaZXua7QUZ/UnOQ853JLyn/NNM0UYxdz5
3h5437vrkdXVlVD6gBD1ErjBLEfNkKkVsSaYXdbjLuuNE4Wd54FgnxodAq0G
x5rYElC8sJcM2n1miVAbHbxu1VmEsHpk7GAAQkFnm7wNClAdGXCI+rrCOf7X
lGHW10aBdElvRWIXPSiG7Pp0cGoA9cU2mFTIX0/eA9pyI3GzsTb+zZ2mw85R
3rZOp0pkuK6KNoOvUmJP+q698NQcFciSKEFAWjudAIsJamQ1ie1b7hxUpOak
SG8JjjZeKMzU6GHCSVBO0kc6MrzJnmetD+IeoXNabPJLWdyOET6GPgWn50iz
W7H8xyQCcx0LryhqVYAKz75jFqMle4RCU/PSz+DYCu5KbjxnPfqQLt1scmox
Tm6k7v3zNjQ404xhBOOMNzEIOyNig2aow02ElLfqC3X3+zzbxwmEBuG5SXAy
y75zGKRo09C3/gq0OOpz0f4TdaUyNMRMGWyTEpUp2YSBmopcVMA5ZgLKjG0H
zIXPl4io/++VAAb54y+ZFIvUJCpz/E3l1BvKotM8d+lnjsUjV+1f/J7MpUiQ
MMPWNkJyPBNtOzxM3sGCT4ZuaPx4pZXq0FH2jx5WAAKKrPSnfHG/wIG81gE3
Xw6RSZR05RajolbB/c4RfvAwOhDtpEeySkD9nmf3k1PTOY9xNuweKtVVSYnZ
4PRhaPL4AjtP8oxa9iq0Y4NFTvdJp2mDj99vGe6qab3JKMVbMF/gAthrhwhM
6+BFAPqYLuUZeZDT1DivzTJXc0dtkQLW7SlY4ay8wl6GscNbdCAXxsFyj4F3
w2BTc9NIjmsQ+S0iTmqgKEn0u1GkaDwhVVCH4LBmzpGtWUbZnNmWQ62coX2U
0liCWR1/N6kN08dV66gfMfpD3XrpS0c7pS1bgg0Pl9oG5y1xE5R2VCC4Sr/l
Fo+IZP5g9slbRjhxxcYTiL0USYZrfzGeFW0pqrJZ97/iV1kvkU0/7O9nqzPX
VpvQaR/3jorLHMdcJKkViRwLIPbO/yvmGKKQlZ03QjpK3aFle4vVNEBIFACl
13aD7vBnC0LYJdfe2neLhJgYlMQQhrfuGVu5yPmTXtGmauuNzVY9eIEoAIxE
eGYpyZST49bUrGa280PSdAWx4db7KQJDZ7D7woMhxKBacBzRD+RQvNQ0Hn1v
o6xXq5T9JeIH5Wzv+mzFUKeCUrdWai/hDbLyEQCv96QTbHAxbOj07LCVf01k
WlDXczmj6rhnIXsZKK12OXgb8LwTEDwIFVUCk1vKXMQuVtJdO1fERHLcC/m2
ZXrTUg1nA98cth+z6TbVEBepx+FNm+Kz+eerR76iBAsEhEcnRGgoG51wSaRc
jjv9JsSZa592EDiUKK/c5+ipDfw9xOM4XHC9h9w6Ft3+PsBI6my3kRftaqpQ
iFrD7j9uaijIMfLiDDjc3jvIbfhDqPfRQqVl+m1abSZbnvMJsT9lQgB+h5+Q
nkRekB6OpSmqomrvRu4UlRVFw8/WRpwNAQsbXLrLmoftl1W/cRULLx1vum6y
QL4441YBSv0QyLAjgsolK019PXdknyo06yAH/IRlkfP9ODv1CZ2NQz3XVYe7
A458e3ZSLTMXcDg5gJs1u4mDFmVCxuBV5Z3859jP97bGwF6qIofaVf+PDPzg
N3+jm4aQ4iFElsEWG4GLTgYSnKCXwnsN54wHZV3vE3m7utHLO12w2eWpQX5d
rVbx7q8hmmvS6ww5m2LPo/dj5LMD7B94cCwDyxMUjo1iRZkt2t1a8VpTIRi7
FfJQ5ojdIuUj4u55KP10Db42i+jCNnVD96SeilwvL+1OQTU2tudfOXMxXZJ1
FqAi6RPGp7UqRpwGqz3ibochlVIIsR45f96OS/y9/nJNEzwDA9Pz3BqOgAIg
qx1OiX1idhSej/0VhU7o8iImAi+XjinV9v1Zeywt4awcIpYyqp2Am4pmZhep
ok8YOxnmdQm7n+Fh804ZF8AX5Y/F4GNxBmD6HPw5FGPhJDGjjnpOZoFdRmtz
epd94631vFxY7mRf8dOrCAvvyx9FONaw11sa0uSGvxqQXHsKCHiFmYQ1/3e8
bnJbp2SL+3/epYwlEBNLGxhVjrgme1VVXREb9Gsfn3WpP4kJ9CTFK1c5x4Bs
/CNEw4DTPT4C73ERNlfNbUpIW2eLqN5ghosPuaBAexkRUEgQuKzv2a3oG4sS
wkVqchPfKTqRd1+Mv1262Pi38B9gRkCkfFgw8KEh3fYECZJ+cvmQaaPPEY2d
q/B6Bd0NnQaqbmzg0m3mb5f0iyjZ2SaUky8QkTihEBefr44y+0DXVMda5Y5Y
mAQxLM6fkAAuYfz8pwGRD+NfdXtbSwLL3Fdr2C5l83P9Ra/ygObE+6Ja1jah
Q9sojckXXySuXkAkx5UvX+D76tlu+ZRRiGSjG7VtAb+tSu0VDSTuRhz8axBK
g9kg4CRqbdT1RIbSPAxrv8/zDv54+ktqnQXOHdfdi4ww4vUpHEr5Ab1v61L4
nLWVpO2sUf7Xsb2uTsYmtRrIWfRBA9i0xHulTyokRUET4HmugWzV+I/wphA9
9+PDtn51MKCrCm1ryOz9+/2/69pbRDQSB0mXcGKjf4HANB4cDs8o9c5SbnW3
guDyRuHS+zdd4R9wGMJo+zIKY8jZR/z1/csZRaXQbdbTUkOOTOo6ShiOHsrN
zlF+xMo4MZwpom0Cucsopab1hDwdO3quVBKjEa4zABJIua1I4h1ikPEXUU0H
bM3Q7DslpRRDHTOnBHLmJn2cS89xXMW9M2qkEu9Iq71IbM+Yq7IZxhw5BE9z
vKLichBmsAqpx/uZNRrhtkUeW+J2abtBCnsWZNgB7GsXSlZIMmZkCTVqTbAQ
lAGGI9tZ6r/cU/xB5yIsSjRwFNEhNMsovgREZ7ta0x/jbLuMsC5SXMY0qP2V
e+11oJdMot1C9rLyzyleSoEtIO74R4LjWCZT+D5ZhcKyCtVpmBjypxc8+JT8
4+maljuch9khKRAYwvq8am2BughM9V6gQfaiLtdr0aYw5Eqfw9sgOMRhy8sJ
Q0hz08X5g1YSYXQh8vx9V44HBYYc+VZFiYVH9WWR6epggO43ByNJOScdE5P9
8ZjeC9eJWW4dVyNeMDOOlFi8UdIc50GTjmD4TUHggXkPb+fItgaC7/nSfsjJ
XofceDGc66uWTDtX+LRWL4QzAlg62kcSHhPJ8oXxFuiJ9AtzODGaAAaQtuOH
07dFk3wsqyiRsfGh4a135bEgt4QgJck3TO2jGRttsgR6h9P555mGkL65uJ2r
t5RVrkJeT5WsWtIZRLoH36r6GcOSNNy37dXNlFNgPb1jiYo4M4G/EKU8Up/S
CD8/QSUiFNoOPvVNjp+tKpcz9rx2tjmgE8TC3ecnfbdKNFp5b0c8XSk9QbgO
B6FyDdlFC6ySpFj03wWeLb+QyvT5D1d5klFEtZhs7bPG1QY9/UvGNqJFU6oJ
Tzl26XsLyQTG7BbqEaerkm+TjCCLQRtgAC9YElnsi7Jb4qLuWv+AT1CFK4th
3eYKYLeykXcCKT+knPaOSjRTb6QSS+Cmv9UDADSzSLMDMbQ11tHne6hPTw66
eF8AyEnPaXNwO3vR90tEjJAC741r4V3Vx570HEdORpegzM682SsJt6wmhdOq
EaCjkKupXuEpQs9ekeFkPLcgrhHVY6KvmNmS9owSq/sqzwLHEGdFaIk91MiV
VkKEoUjL2aLx2JeyBubfLJ+IZV1wqev5p02wRwL8w30+65PwQaNsL2czbhS0
/nqiONamMGH5f10SsmLWjD5NFORcMq9aOgQoEvjPQ3IOP1g5S0pXoafqE1LF
L3zzzFENwPXJPsCe7deJDe2Yy/ngedJ3j8ZDjDzQakElKgAA3aOzKZZsqR+i
7oRSzzkaMDwr+P3I41undvLpM4GdKEoFrpNiDwHkcuOYI8FRTy5J7qvXsnEa
7Q7YA73aDx7pzEWqv/FYvVZSLSL8AGOnsRNMPJxlYwSIxV80ILap8ixrN/VN
Sw3J+PWdR6ONqc7bC+lqi5ZKpT7sAzEYqudt9wKNv9qxHP0KoGSNVGhkjVBI
KpbNEyYsajmq4B4lRJ0hfV/EXWNnQM2Zq/XUvXcL2ZFqY1StrNcqUKE5yF53
4pXL748V+/VYaNEQdL5vLYiBUbmdlrmn30HagqXqjbiudprlnyxKy/Ic2JiI
oDJ+MeWqxxO4Vyc9YiMmhic1yeRwMpQMVZ5opOLZSAwPa2lAXs55Po666iJI
TTu4bBTYpSdRuppGj8jGYqQ8FnuMxGH502q/QKU+ZlnwyQf8SKLYvpQvpp/V
IvSn/Kk6hUzs+231GWtN2vaPzGGTqDUNSYqFx1WOqyjBZSIIPPvhCmo5TU/g
O6TmRmuWRQcRIOSptdkjxBtE6rtOj5Ivp9XLkK8qbnuc+7OFHwA+T6WWF6sI
czvhPvVGMrVBsUJAYSQmOT0LxZpJTEkqqZwmo6Zfe3zGOqx6Ycct8zmLE/2o
Fw9p3cJbOIIsZuowv8iNFfMBOEySHAE9FNmm9WwbXqo6hcvJbWSUx9RKgSEC
fCDomIoXjHfU1Cfvmd5Ksa38pWoV3W3A4m71D/7rHZ3rudZ/1wm44IJWmiuM
YVDZu3WbJJB2wLNmxHmmwIs82yLP7Z3H+W3UlGCwCUXViw51sFEMcKNToUyP
xqbRMMzdSZdukLBujJBl9JXokBVsycF8Xbek9P9tlrmg6mxpiWiuvjf/H32/
Tfe0D3VK8Nu1lUYA186yoTwY+Bi26ODkz1S37G4M8Ri7fIuqlJnNuh9xq8QF
Bi/m3kY6XrEuAMF+tkLq5gV7P7bJ7wxS

`pragma protect end_protected
