// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OI2i8m8vJPVXbHCJ/NYAx029mJRwtm1ICsJoBq0lMqLarrLcdvq1uZLaFNY1
IYGIRtMUdAkEXIeOld8NkrE9YKIKnx3UW21LIGeGfLG5JwpF4PEp8dnoBloE
AqcIe2U2qVdFj5Y3gQ4miKA1jtp26EW7zJY3kX4VciIsixzgiBuPVIC5Qyy3
XQHOLi6UWY5HpaxXD0erm1DU6OujDpHVH5OuAYKnEaqi9mhaIpkmLH9ISi9A
/akbHCSbLT1Y+DejXcqrKaNMp6JGCACohsjbk11+97WgaYAwoPenEVtzjdYQ
/6tLdft07DTMSTxdVpNVJZWKj9J9RRiQcu+OFgVb4w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BIcw55Y5Ie6BWAUqO4TveE05I+I9pRVfgvsEJtwJnGl/vW/Vc/7N4dTSPATW
iTBBEtw0hIYJpc2eaoLDu0HDc02PCUJEz0pE1mYYTHbkrCREFG8avVCV+O63
36CQxpCJbzFIoeIK41/YRWIKUKmt5NoX8oUj5ZVwuXPlUqmT4BZpKHrpXYG/
bsMG6W5EQYqGABZLs4MW7mQ8vUZwxU8BiYVQyaRbjUR2m0WexNruGYI0lfea
MlPtce9XdYa6JboR8juHxnBmSlR9iMzkm4UcPXjNdwnooDY6Bc6IMXMXbh/G
s69nE6gn9w4MAxGk1xpWcCbNcLhQ2tMVewzFuzrrfg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C8GYTcVF7/0oFmliOtdkr4VDIpokWXJHAu7trCQ/Awr7C7xbzm7sQ8nIOoE/
Zp5ja2JzQBwi4pVp+ujOpnH9cogkE1TrkuMyNzVoMztfmB9FPFwYXpPPdKsT
UXgf83NfwkVu6A4e8yL+utuKtwN1nTTpaS+DuxLJU6XSTr5d9jOKkYKwyS54
s5SbMJYD4R+Uyvl9idcBzFEZF5vtwD4JPEveTd7EVg1li64z+NQoPx7b9dUw
bcTlQHlCA5ZuHkrpoRbzo3nTMF8yarmfb1Fonavj6aZzMFM31SqNl5GSiohD
m7vjIArPN+GeHnb4R1BTuUdccfQT3X0FfIszrmb42w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
asIPK0k96/CWZ8/TWq62d2hzfzEn8Y8IGlpPyHFONcIJ82n2gt7xbsM1AVax
XNPNfphzBavyntGmn8w59SNqnBVpEWxRIZu7dAQFOQPxp9BBGJEF786DudIa
FgjhX6BY4mF6yzX/RME2M1ZSRdNPS2P4fY5p9sfNHHouPyPNVhE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
has1Hm26pMNB/LwGiXn3zooaYgsQIdxi9BOvTNez2xy1WdSOqcR6TqZavBA/
02d1aBwgwBGbpC0kXX9nSM3eXcQI32qIAEeoL4rRLwsis1I2j5IMtwXzlKCL
g0fnAhkqIy3zmuhjTPOhadSDAptsDWVVTslLqwrNAkvAPFaJxwhho1WB5/or
p5T/SWZHuvc63FcG6VVtyt84FYaj/btUAlbBOF1cLK8LvxoVpbRBROOOamlz
bmgnzwLjg/GYZhPv4RFtyhxVp1YbC03HnOVgPMv1KRDjTEnzzpZN4T/fF8GR
M1XMgQYH+WIDbpkDg0kiDhpSv6Ebw9rEui3QpVXGvos2NTALUF8AmP5zA0x6
xQzlepWjINk1vJHVfu7n2MMoaP2XLLMp64AvDzOpfb2Yqs+fEjQ/eNX3ogWF
JoiE60S48WoCBuwsDdbuvLlwXk183Tkxg8SYtUBUUHoGNmd77GvKyhTJYb7M
6tqxCbBJsytblkmhbuUl8JjOU98ItIQ4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ms3u1R1dBqYCilUuum6CStZOj1Ga61hXybA3dCjoZiEZytv1EOMeuzlKo6bA
zoiLAoHwXS5Eum4AZZyryJFNX03ArumCD1LWFSUknbfgEztj/Pl8Lftuev1J
JNFigVCKaNusjI1g/IbG/3jqzoi0PhE6L2CSfPI3ABcZL+rhIqo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IJZ5jtCrAo3H1aJTkvx3iVy+XsAmSOzwMoiY7bS992M2jHTTYiaLhznw8t6/
QqizbquCHQRxUvmgBHyl/JNFyBzdDE3QYOppllEeTzawJNSZ+9FE9L1t8J2o
PFJB47qvDWkQGzGrhxtXXPaoZM9vKfTS2qMg4FGYNtXllOXrkrE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15904)
`pragma protect data_block
CdEDYuo3z2wyF+i9D9Q5o/zIPvGf1H+XNqxgMyDBiDqd8evy6e/VhlGBTHz3
HpZepcpRpHPgE3Ocp0p2fF8UBdg1qrsFgEO6VRBpHHLXevH8OK0Leb8KHR2K
GKYsIWMj/BTCphoaCmkfhfIZa6hwLVb8LQiFbkHlAus8RHzR15PXTeMm8Yh2
WZaHfuKjd/ThygAD9n0aPQdvOGxZ4l6ygIgH5aCcxThKPY3PuQXZ2qIV0Pzb
Iicyc0tiUG517io3u5p24v9k5QAH/nlUAqmWfieg/UD6OjBtCcW7VxeQfJkQ
aKM1dahR8x6wOOchGdLo2yV6NT7kKwm9W1Cfgujlv7RhafaPQ2NqHKGOgfz1
3DH+ez4dwboTATqb/0xSCf9AVg4zmjO52XCYmpvGYBLrO4NI1IiNVBz33Bpn
VBAvgxw97UaalSoO1qfWJ5ojBO/LotmjZUaXpfARBTFNJ9y4F9kTbQOJiN+K
ATusnXFc8m9/pdoaOHZAItDPv6SARbqngvu1U5ZfLiErFmdlpAB1b/8RoXPo
H8LLhyM1kBeZPJRRGzLagZDaqbAy0+98lRnEoCrab6GP42DWQgemiAIYAhJ7
ytcGm7dnj2CdYPIyx2U/XuYDHvIcd8MwrZuAoWawYP6Q7TcYPsuhS2l1mnCL
oemZiv5zAaM8bgi0HFNT3jBQTfaAKLUNi38NwZsDUJh9YgOmExzHKcyytVfl
sFVS9VAXa6okJUN26pJZZLUbOSgbWfw2MDVn2mX7GwgjCIBnzflWjGvza98c
rASwBVAaRI9+mzLfrpTrj+HysLl1SIj3UTD+ZZjhIRo+QQ0f7Trs/GtdL0Qz
VhOv86a1j9BCnmCJe8f0GQrm3s7SdoO6TqTm+kPKjxlaf5sXtIo031Pi2uNk
7RDwshrOaZsxoMzQa6N1ZZ6SHDDvIXnqcp7GvZXVE7VhPgE782g/glpcaTfk
BskMHqAmGhBTpIvGu9l3ahb/HOxDXT3CGmsMZUwXkJonZh2Dss/XeGe2SYR3
UTRksmdOrCc+zTOoY5KAJPyDjF6PC4v96wLxYkivil4+n3DtmtmTcYGHOPcx
tGbPXhupJUo5lLNa7Q4+A5QoQGylHVawAneRzJU1AHbvOXe+Z03acPBXg1jt
qje2oyYNe+b3DC3kk2m27NX6S1NBw9EdV/kDhiZFay2PzRkQjUKaQdz3SNp7
kc03wFswOCnZYXz2xfMxTiaMdwuum6pO4Exm91SP31TUchodXcHdjDtQ2I7a
2c+1Wic9gf6TIWZqP9ZL2JX5W+SlEDgk3VZIgyKpNbxkpJycF7e5Agxs1OfZ
n5lG5/W6ArQredhXy2IWOvTZgt7nCj74DsKfCZ3OO9I/uB9LfBuGdaGVJ8Mt
f08F2hkSHMbI61AKsmDZcwrTCM9NJcXoO8/d9eGm91Nlug6OHQ052fRFX9uB
AKweS3NQmWCDBlxrQHqCeNgm/s0wNn9zptIvECbp95UZzXZD+tmvLgu5lLZK
YtSxvCOnTdo+h62m5pS+C54O0Y8CMXou7uAOwE1LNOmDj36qub8fmddGHqsI
cFewiWB8XBdngxJlBht83RQMGxfEHT57MEZfVMflWCaOl/OVtwQ9oEI/PbWc
tcWLaVk8AWcrtOCMgI1H3Di8CgzMVw0SLvifRyrsqCRZtzEA4Vkso35Rb/e0
ajwEdGp3EzKk1jLfuS5+7MY6QDgSMVb03mUVcILtbc3nEZjIxzZD7SSu/yCo
dPPqameG+toF/bu+ONQOYaBVWu+DR73n3ScjQse/8fCGiLFXuxBaDvvLQV0Z
LvgHTnxqBlH3Xi5JDIkyiC7iXMo3teY0vfhQ5aSNNpJRdIngzFUvCk5h1AUI
nVq9LOmGK8wTxQ+I7GrnKldKFIWUtIC6nEom+i22GuQoaPCmBR9oM0jpAA+I
K/m/Cw9kDBF8rpxlRDdogk6Q7jZwUrkOVxCO821583y2azum83tffiWn/tj3
omk0vCdbFtNVRKb5+yVcDkYCmWoRaVhGgC89CGbwW8YsPLLauEpY3/55jsg0
e+ZKvw58p8HLr2xJTid41AssOUlD3/LpC9JKtHh/pmvzESADtvMsTrWv8qMB
Mh9CAiFsyZ2CaXMStZU+R4Z2EWizmeH0YMMI15DOrsLY5y2ljWKASR9HvNKp
K2GaJ5TvcK8brSJjCt0jYqXCq8Ce616AgPdDoKueHYJfFLPWbtqSGCZqoEm3
AsrI0BtmwVHJTvhjd4OAG2SGyDeWcEMGPkJhcuiUa0AkYmClSY58e1lmd7BA
U+48iUTE6b7DpNOXK7BoHtvqLm9RKlZ6G/TaDJY8QxfDtCUgz8nrxXEIwyI2
nFw7KR93Ntv2AbgCNYfgSpT3Obq0RO1ZYuLZHY6yCaBxFE2g/f0CLrsG7FTI
TN5PGAfrZCoxrPfck0HntvXoCvEVTgtO2YzY4BgPB0QjF5AtkDL0qJ3LoAiP
Tmt7H1Hxri9yrCeuZEP+MbhTQfTWHjzpBPseuKYfjPy0kOs0MU5I7u7jU4Zz
SHmoNp/L9RmAQ+PckSfw4pw0uqOJPHTtjb60Eqbd4mogcR544u7SGGgF2tPO
WxiT80IqRXb09hN9sLoBuNa+fMSeYSPjUPIbrXWVb3+8UKzIx2RC1CU25fdm
w0xzNTJ06q1vDVPF/yGzis9c6vmBpEHjlvEf9E4lB7xR+PlNOPjsaobrMCtY
7Egs6ET7H+7+g09aRP7SESeqrwdEtHYnWwWP9KVPATq/dEEA9kphTsPqtPyi
V5CynCt5ljyfIPwnBgNwY1UVOgliu/54/9w4aa6NO8Z5NaHTipiE/Zqmxxbs
geE9vd3xFf2Zo0gSK3WDhzTDB/JyWuygbTwlFA+D6mV0sJGMUkgDJkhfhXLl
fcIwnmGd/C49Ue0wiUHkzYEuNRJA+BqArjFE8Kj79PSWuycW201pG0TFfggR
cu6KECQhtnwIRmNuF5zVpJ0wjfnIhNCRIsDRtTYVBuaAq4oiBwg7OBsVWeMz
tCbpPLa9HvKr9W/ivhPLblQu0KhXGxf3FUmP/GCh6/8ppvY32HCIGK20+IBC
pmHjpVBag4x75S031pA73mrzYbCfz31Oi91dJzsdmEgrDee1trJRcLbQzzpP
YFF4llf7iKvoJc8aB7NkEZXXkHaKBa1GO762PY9XNCZgHaCLh9VSH++VAEeI
Z4YJVFpFmF0uvdugmCGuszWGJKC/ziu3XG6yzawuPoaBKN/3hldyW+oYbwK9
P2qWcOm0Vequz4KpdMYsAhpM8M/bLhQH4Da+s1eAWcpBbXCXqCLoTLkXAFId
O5wCIgJfVXykjskI3GcTAOy7AKiCFrQoPraGoA//vs1jMSh/g3NnWwoQDwyo
uBJeGrW6JXPG68tZc9RflkQATt6M2o360yCLBiLklsSIE2+l4AK2kKTE2kx4
+J3TqGxg2P8S4R0o4njMl0LQZw8R0qMmv7OuLdEx0kIP+ncEh0VxZBjSkhIP
SwznQr1U+m7nfSzeUOER8PLZa3WHLKrl7/efx9dcSUM2hKs+yzgyKx0UiJXU
LJC9M0lPbIHsfKei6TkdfeY6SUy4UNO0mw5vC/Jaf8zOKiQJHrG4k1dUwROk
ebFSeVGhoYTlgcvfVd1NdJHGyj3DKl9drxggEMqDe1wvEI20KrCIhMREZjZT
gyit33ModKeA92o+z0g8fuIhfzMQ6KMj6fagj3H12aCJUD+HcdG+57WtPu2d
vNWzDYJgW8ztzAXKdm5VZOeLaXY97MVawUmLM53UrVYeuK8OVzdiM1Ipq8cd
kjhkI5kbuKFbd2ya6vYfqzXnwsdixELSW2hlFmnJsUpA6N1NVyP1O1KpdIXv
o5MdJVQRG6CjkAqT7+XgMj0g6ZA+0O22WANl/qlvSgFmtX+oh+VeC0cceKkh
FxSAFcfo1U/suHB7R4J1lh5pOE28+PzlHThcAsjd0t8bvtnnJR8Wdyw6Lhu7
iA9MzTaecziTBzsx47Je0XvK4EWgXcSzfECqclLRNZ/dVVzKtySlqk5s0Tb0
rn3P8pE5OPvtbdxfCX91hJcMxy7/j3gJtQhXUAbENQBaBMUgF1hjBk6gNk89
f56AqJ4dHeYYmJl4jkikImppE3DlJxJ8opQNAkwKsrR41IrKRZkT2NUPwMWX
7ayI0R0Rkjdlo5jjgSOezHxbVTRIUESdtPaQ2e7YC66ozcbdcvLGBwxka4Qh
0aB6UK7X+yGuW49PQlBp8ZI9d44eyxhZWYQK6kRdQBNnd3c7c9ukdbObG7j/
cQq1C790OqPPWcOxDSwEmAsjh804sZ2zqk4QjumU8YWfjSJhCY3uRlgaEBS1
HDHaGRHV+jPmbu65LNey+h8Xw2xI+KUI9gdfimkQcwbSSN1ov5+b0ubxqgXo
HuOXCC0nuCS/37EpPs6hXUOfP2155+0AC8q5q33jHeA3LQ/9xwwLSp14M5gH
hhBaacaygUUsPpGeGxVHlIEWGOc7m3lnzKC5NtZf+3Zsg8+MPdBS1EYrdVNy
grxvtL5UKtCNxhYjCMFS1UK0IX6YhJ9KzGEybc0u/EW6aBr5ROPevtY/9lu2
Zbo/Chc/IuCTrl4D2dz8Agf3b/Y3iffUmVQnZ2l74V0LlzTbABX5CEZ1itrp
m20GWZKbFI0xaqQmLgGeywDFDfNkPmqINFN2+5vjplK4A/KZ5mJ1mVyPUorh
4eiJU0Y5lj+gJZlwLbr8Ica4EGUr0DJTXoDV0ZAi3kszaBONw+E0Tm1X5R14
QMbU08/fSvK/QMXb0cOrxmW72F/eqSPRPpELVfG3545IAruaNHJs7vbMhJrN
QJ02W9gr4jeywTnzdDnNeobzjeB7BaPcmFHi50oaXjw8SDEaVYG3s+rE+1g5
YfFmLffX2KS0z1zt0mYHgj40ObTGVN9VwElfnG1holut5ThNhtM5M4vAhfvZ
Q5RMsOxumsDZ0kuQnMdf1I05aFl4VnXm2ddBWJhSdo+AcKN5nN0xev4fVoTd
QSRTEKJK01MTq85QaPYSKtW9dWdesuy74AjxGVVbbSIRBXXfqFCN70oWrYKb
pkPWQoMacRemUFsTgmLD+/T26Vd+hFSisVErwDLEMud4OVMrKMDApMGWm+yy
yJMLizdur1vPwQsTE9lQMflSxM0NaOCXu9vqfTlvPIJAzAHJGgd4ji5TLTfX
F9FUMAWDEtlsiN9/v7KIpAOtYM3rMXkri3LHOY5aOEpXR2L35T7838uWR2aF
ddbjxHbTBYcX1/cjakr1jZEu8BkptAx5/aPoOa6Y4WLg92NyoFh8Vljd6NWB
we+GwwWjL6LMfOEvAaQYGO9EGP2a9M6L03RMLsPx6UhgeV++IHCljEk9hkOB
Z5kKAgjKQYzwwx/QsRC8c+sBitSY5WAkUzFxm1f30+OvWZANrkoUSBd/UMXJ
Z8XZY/d984pFh/AsO2R5GbnIRGB0A4+YbP74OMCXxh6vNX5Yn1GT2PCsJme3
ZlUKsUCeuJevH4dSKzS1CC/smg264gLkJ0vX68IIdtn0GIu4LsbslUyrlR/h
rdiiHw75vjTijziKNCqmdkLWwOL4flREr2xvkoVRDMOA+FhM0BS17q+aQ/4c
i7AYyBfMP1AsbTVt52VsBDRlw+3t6yfEY8CnnKmqE+0Di1rykWZI208/hdEN
k3m3SCsz0hL5qYVjN97HAWxaPhTreItbaPrXNZW390Z7hzwFDZ1kasGACNej
xpnxWaLhTrn/VZZYM5Nll8hd1yyLT0jPGYtq7H7yB4+NL2ZbkSW9AnSJlxq/
liEdCQh2zCOUzlpNdCd/YOC8bAMhS8xONhPssF1Fd3LNBc7oei1my//ZTdf1
luSVb7zfjSri5gb3U+iSzEIIGHn/cjG+xHx+dHZaTPLI8tXlF6GKErTQ/M/h
v6UEt6DSACcdhfOl3sUbEyv7cVtX1oKvSLP9pKVLe44pDGCrsk7Den0SVDBF
F8KJwYoff7kmBDJcUvTMYNGMk9EIwDXCq5fabpEbIA+wnuDxSW52jFPV0hLX
hByupQaDa/g0ISRiZdywAcMP0lQLZ0D0e0lr+LPKTyfQJi8wBnzVqcHUkOXR
s24HB2MmHT7XHYEIdd9O57WHdbqKPp9eNnpWYe9qt6fN5EFf0FIJcI6JcYf1
+N1+X9+r+7ddjyxC/vaqxvVltx8OVXeFIWTSs2vmLzGp5LGmoEbaqy80AOok
1iQXlh06FfEZR5/4lVy2ix+1HFAri0uzG3qUn/dKRWqJGVGrTNqKiid9RFhX
FwUMaV11nxcD6+BzbS1AOury0OLmWHVDfAr40J1oF7RzF2WFy7DeTtq0p9HX
/8PdJNqxHkAubXJEgLMbFk6fo7/txnqazkfF2YD07Hgbc6IUNoTDtwE+yiGR
mFDJCuAIIr1g6acc9pObLZJM6AGE06C4ErKRBk+WS9g1imlCysgtkxIV5vha
hvOjGJGMWWcjyqr9uJcCv4/lx0o3gYRET9ajUhF0eJ+1aA7uD3LCqkFsat5j
IYOmHLLE+8I5xNJx/+HOKMG2yntQ3a82xVW4kDfVPPAF8cKE0Lr4iB/tR066
mHBMG9gVJwI0mBjs7SXESsqd8JoSpW6lmnGRWmgxJ4iwWXa7a6aPiwVZdATj
5Nfb63KTN52ZQZrD3ayRiX5qm9yMPhbVr8LGmP1ZlLG+IrClg4l4HTTdcy6x
LDx8HhBzroSVuB3HMzjhnDx34nXhCBxlD3BLoAbXEdyh3mUJfZ5qNsG6J3DC
/8NgnLehY7mdUh7n9a5WtJvkimlBXgVOraSUZbsgJivVuChX56dSJXY0wZPp
FXvfGGbpml+IsE3nmG25mu5qGCkEix2mbdjTCmS7cVr2AcQOwlxLtwZkd62L
QrmDHnDJSVlDs2zZ6XXAtUt5yUuJzrzEhotK/RLjsQEB0bDA8MzcjmE7sT8V
U2Q02qnDRI0/v7Fo5V3ZpxTrez+1odTgSc77ie3xmaaVTyXkO5RG0N1Oufmp
18m8HCCfbou0ZuITeijBipHuzIozr5lAGLuhamlg/fhlDUPdu8FM/qZTkGaN
ohs2ndUYN/39fR10/f8ys+guK0Ejd2FWJdZp5wChO92bPKgn+vLHNQu2rQiq
qKooDrztuLp60/EjdSlbK2zYJePzLVW0byMSqNT0i6m6MQZomPD8j3fmBAPu
Edp+i5VLrsxqS5WJhiV4GvQASav7aTVWK7n00/mIza46t9FuDgYQpHc4eJ0p
vwhusWG7nYWc/wUNThZNQL+9fU/YrmbRNwVliAtObqyhAzwAVU+wOWLtLLuP
OEDueprwopLLR3sm+qV4gC2jf0p1+3Spdillq8yUGeWBIcB2FUBy74qUQ4h1
evlwcT2zETb3JJMEw85Y4fmtU/uIpVn1CZYDXI3trHaMYirGgOgbGG5WjeOM
sOxbctJyhKlQ8zizJWETu5xYdbnsvxf3PVTaT5aTucQgWFfNoYPXJiux0P5f
5DxKRDHbp4byxdWB6eOGPmPia4cthQRRwoG6rqVKK3+vCQ9Bb1cIEZyzw8a/
md1B0mG0ctU1WmciXwQSWAkPo+SfLz3YbhR7fTNs0B6r8WTbKijS54NlaeQh
UnCQMnf3kqRLy9n200EELlrpM3X20Jop/el1DaddccX27fqr9cGN/J9NsVYq
/n73SQsWreshjnmKU/qWcrdTagCHga3X/4OTWzUs2F6fJWvbdtY722l596eX
AgEU1DYKDx2ndUKAETjcULiuOjYCCTJ45CM47wbOUFdNg7ZQ8Zl7IiGwUOyN
oppYXg0sQs4EEIV5MNquB/WOPbUNFJ/ktAZhjFRS+ATO0IXdN2ZNegQ9b4Wm
I0fsSyidxBQhWaOecZj1dXUFwx0wOT7OVpmqprbSBmzM8JSBSuBkKeQhbRng
PsH0RjvX15WnhAZHhV7NEpqJhbCQVtXcvKLNOyJ+xrnDq/T8F4ZXeBagaW+C
ve17Jl7qR68HPBJcWFnN1R0Y4a5j65FrfKHON9J+S9+S3b7FN5RrsTFpe77v
tLikTipjRfYH4iqpmU9/3C2r80Sx640cq/0gRWAqWSaJ8xVlVke1JOwdxIci
DlHoVkZ9hHluMJmYqjGmCY6qHCxVmDaRSi3umnWybvz0VjOn+oIgXFv4srhx
DzQg0Zi7pLzG1AsaR5V5hnwHILioJSGE01uI5lsaRCaunTZ9i3Pe3pXBXWcN
dA+JOQ4+6kpptP0dz1UJ7HPbTalz1Yi7BGj7AhNZhg6HNwVfoXJFUz4EMs9o
prd7lddY0Leq8VYegDgAg4Cbfy7//nnTr4QlXUd8DwBkjxddguCMqObBNL0V
YSxfbKQJLdl+6b+gJYn2CqeS7nU1V6b/KzMlknDXyWL+V46cv+wwDN61AI3z
XRCEhzPSXi34M/MDk7qxRdoSwBdUIhHifUddN/Ulq/Ft9h7ueE3NoSVLoZRt
9oIoObtIbtKsQT2jFgG+Z7x1T+Ua2vpfblTygN93I0a/rmqrD1O7d3qDwimS
myWNiDtk+bOtuJUUWKRm0WGyoGpycMeMojPONuVnIAo1OdWW5iVg31C7LZWt
HuKnpr/n8hwmJzlmMfoEdSLrPbNI5FuRPlsZsENZe/of5ullvp/c0Yoy3ubA
9bkHl7JmZxnO9/effQKxhJKDDN4GhecAG4X9WOLvWY47kXlDo6WzOWgBVXlh
EOHjKsZS/k7akIJ/tbjO7eZDz053PnsIcgnHMZpSw0G57XxpvOAzYNcVsdD0
n2/MZTa+mlvu1DOWV34jOgNJe/+m8fwy70FyGdutgRRRlW1feen8etqVcGt1
jqCkxHc22bnlZGLvfoMaIrc7nKEsdKd7Z29yc8N7y1sAHB90s7xE/IcPTS/I
23VSjHHEl07a88bJHaxjHatcPQRXuop4sd0dmDCjueNLI7/fBq7Kqx1MFGdV
4W+hQIshWteCvn+L+wTg49zxoSoTCHAfgzkQ9LjyNjZeDtr7ZGJ0yb3lCUJ3
48I+4FYTgKej6w59S3kyGdx/tK2SRS2iC1kjNochWFMs0y+sb7E5hRynMgTy
AqYmYhTPzB+iJQINt+VXALSXQImlmelJ9oaYd317eE+7Hb10GV56dQsE9PdH
4L7dPHx7cDsopA8YEIb3EqmfdrfskGg9TXFtgORAOREMQbC5ODMt8SxQ8ThK
R1fUuU42Q7+L2r1eR+ydHeB/orNy0fLo9E0IvzHYU+hQSot7pbKY6fa9gblo
tayWG/a1UUFGFjx18/yQt6rOAK+Qfb8aHN1Sjy5SKYdTpLRUQXPbiPgJU2ml
o7E74VjfVNGIBSpegno9mSUusRH8bA1S5l4K12ayK5lT8C2HTK8BXMQZFaXu
cGyBT8QVppSl1Kda7BC6uUCGeluQg//6VbNAmj+EbIj2FRJAzXHi8nduMdTL
1IOaUjGdswY/gLRBpuUW8a2h9RUYuQtxEYoIFLUQ+qQXIAneR2p43TkAeL1B
jobQ7MLbNfx/4yt3cgO+0LUxhD5fp+wRGdZxLQ/IqknVCjZvFHs6RvI1w3cx
EN42JjPIHvZQxKfSVKMt1JriUzDaQrZ1Z2IIq+9dfX9n6/2B79/1szpoWz9w
bQyqt3r/0r7+v8vRLSSditnW1Z2ytpuWfO1zytosqpohsvsvRGy5gccNjVZC
IvnoW7kFAtAdY6IRNKSBqaqrU1fh1F9z1VD58WOZHm+Qrg1AJfG18v7z4b3x
Dhh72WYja7bMqqVuRC5dIIUNfVe3vxLeqxWUvSzsdKga7C0+GBgQnrpRp8g3
4j+IFOnGtHBlk+M/J2ymWfPfhuHOka/yiEqmVrjm9Icj44rghQmw6bKtrbWK
x47MXmFmHOlSQYSH7bmqE0MrCfQJVJJMXF/dqeyFZk2YfD5ZQFfB6wLTTLct
B+dm7iGRrqX58LWwHaT9hW6BzHgWM5pADbCa9VcgWfoWRsnZJ5Mapf8tbYYN
0XZGoNsEqO2hUzyhA0u/RtnxjjFqZ6DcwPrN5nT4mYsW2i8s0Sp2H8yMPBHe
qnbv6HIHk86uG6xbolWIoh2aVZYwy67+20ZRVCBSL5RJ9LcylVCADSx4M1h7
IwqupL59YHs1lXIU40u36vTItoe1GToBvqxSH9VLiJRucsnOk30q8lxvPLYR
6ZdEqIhX8bcJ6OpFj/YyAwIzzsFZxbpf8CfXWDQXJ5SHXBKjf/pG6qH/D1yA
XB7bxo9qf1CuDiP6CGl2YcunEdydiNR2rerjsvwp8j5BUWaAEzghzBl0+ycr
7WAyuRtL3zzo/oHixXlJcvBur/HJZbo3hJ12pVFKcpmlqUGj4oRPLxRqUE0I
IxIktHXI6d9CX9/CAjMR351yL3UPLjyrCmgrCv5rATHGrJqjLv3x3eUstiKV
uhLwWZUdrzMX0PMAU1p2nEXs7B9beTK/rssD71Sa5GhpdGAGMhGaINxJVR6k
4MVXgT/YP3W5MZJVq5c+zN/e4PCADEM2Hg9AViLL6gg1zzZsRaynj2Zdcg23
ZDdDhuQPwMEbrlYAm/ZDnzEgg06Vst38gUBI1E1QTAvaKICpnWLpdr5P8VyP
aRXk5kbxWSoyo1F/9vrnGaW/OO6qrlkv7fr8MRbWgLaJ3CQIvPUMufhHLQbz
kk07+u1H6lpBy0cVsPrtZEzqN4u1oM8eG+w25dPVqIOsqu2nSmpyCdiBsiOm
QodajK1Yza5bbnI4aG2djgMxbuNyNKUdBr7LSDv4uYZfeMnkhsoH9sItafnm
MnUSA8AJHCxzxZKMnViWtIEwtpd2tc+HaNsKlqh3SD/iWZGvRQs1fV7jrqFX
xDCQ6BgyNQ1SeQaus7p+sgRbLsLnjZ7Qe4guLCwjFsSX9x000lsuvJZxSzb5
fwuI/FwLP+yFCV7Q2HnebsbpKsWl5qmYFAJZNLLlIXoPdUUVCJEBoNMS3J64
l4eA1YtKQfT0IVDLX39K1+aoy0E44/tCUB478o2ibzSlGvlHHwpjJjHI6fRB
uiZyB/a80cKDqaDZ836sHi7Xd4IujpSjP1xjLRwHm0fX2if/B5k3OqU1dlGJ
2bOOdz4ti+8R5zTUw9RI9Zd5jp6NFNI2XjDmT6vv9HMLZ8P9xFNWNMNzD1XE
/GPt+0MVZxqPQhHxkVaFgcRii2IyDxh7Nf46APRmOmvO3PWZEMeIse5V5D7B
Tx5Yt8hgir63poE9X6aoBI2dNFY29Vb+wL3qNGf123Hb1oy238EgnESGjgcX
dPcJoxuKCbhZaLOJkcIi8ViTGPtXGE3u/lNwlJMcSB7nTOZ1+Jkeyox1Joln
qR9dqJsitRCr2l0PUx6QcNVUQ5ecb2mYUHBHmJsU6wGczTvv4ktTnT7idPpf
68f4ZwO0xWrrMq5R8Te73GTAtgamEZBq7PHVhmRm89YVrwjyRvCqBNf9wFlx
iRDPrNFLj9vIiknKpo3V8xwsUfQBSg4t8uXdTLfJfHWYqpyFNOabY44kH4x6
zX94Tkn4iKn+xrw1E/VAKOijvKxgQV+ACQueKbBwrMEAdNN7+N18mcK7rgUt
MY0YauSeL9EEKGAo9ETNiHGpguTFRjnXSAzLMzD4jd4+PcpRzeCUdhNpTHRl
10diLq6c1kY2MXkUwh79N99GGCeMYtY6rAeMfub5xhnHciwSQ8a3L4HPbobK
zG0PvglBGP2oh2n9MVyM+meU4Q64uTY3hTtIW+OeA86Je/9dEAbXv5+lHDb3
UDDecrEA39BDaWqYY0kX01tFSPoUnlIKUW9UFyLK0o2U2z33RqVaSSykaXyp
wxUkPRRHWL0oQr7oOcz33wo8uwTzoohIGjkBa3g6Tw1/NRJQiYIG3GihqTTE
Vv9bzBq1WN2gxlpSl0ZLxiOY5OSgadg2f0MwJpKDnXXhRDLbMpoIrm2WSy+y
uWY9PW+RQty53k8Jf8tKVXIK0Qs+Ep4BbBXgHUpc86Z5oCgHioUcvb8usw6s
DA00MGFFrQWY4Euq3FWOjs6nj5ntpxSYJDLf+f+zcuGZEUW/py1ZGibV7TbC
YHZQPz75sFybfBgl4LxqWp/KfpaYFNFEKT2Fkub/x8iEC7lKl2Ni8EgkgJl7
aUwXWcnD/wU5WojblfJO7XmfvH6uRQKaHQaek+hNLfK22Cd9CLGKT6ux4+vp
4tnVS2eRRRHgCS8OKOLNaJQ0/eo4aBVUqMJLRiB33+RS6PN8xBqCt60uqYxr
yirnpUrRT1FPbv6/MdtBX5yMTwK+OqrMCbjQcye+zLGvqSVokyzevcmnv6bB
t5ABMJYITX5lGrJXAzXor1IJFa7A55qqpA53FFeCzfbomF/+NsKWH6fvvRWR
d95tbyz9jmFegsBXNqzyMK1LdhsxwdNbLUhKlLFVf5+90/red/s/hFcfNMh+
g3UI+gSw7wFdw0yYQFI8RMSAGff4oYfaJDC2zeVlr+nR6aUNPUnW9MY06Hje
3Tl70WloO0yTXI2ldR2j7rIb7D0AjxshWCQmlvwbtftZjDD0ehNs++7ftckM
XxPwBprnB7am85xC5ShBM6nfS90RuCQR60NJWe82SVUdKs2Ncz38aXjlLf6Z
BnE7iG2woNIq2VUzDXCnjVZEPOWfFY3+AU4IyCy38dm8lJv9+DPgQhDznBu9
LIi0Om+MhOcMSHPIBF2gfMSqtAQgpc5SnZtXMRkRwMqKCnqcM/FWGPCV2KaN
Jos8N2RGD+2zFDN+0tnLpKG5dEnmmLkp9SEq1kKDNHH6f80vWoXn4tVU8x8c
lkp1NViQIHAuHIbHF/7XWGnn7EMme/HAVDq9/NftSFchLnpy6g2W8Gs2D/X7
esZSrCjQwv6i1rUhwwN9Ox7DzUrijulPT+gbrQuH09y8J5u4wZ08gc1EUtow
Pxq99vjXP/JcRAbYw3miT1RAtX+LhXphi0mDEDs6CiSzHiKZbb+I6BTihgy4
CNgcvZx+HGRlAzNeh6j2MvrmXulSiI+DRMnMPgolO3QGxWpl5wEFMcPsVNYb
WCC7jehepUpxhKzQpHMp/eFsTbcepHRtMGk6KKBAksKr+V09xsTyZ2qxN8hv
/8JIN7xs9vfp57zJqRSU+m97u/KY6jD028t3+ZF0P196x2Syi1oCwAplGTp+
PDaE6+D9OGXdauOxpwDzvzxOOIsV4MVfvUlOcHG9ce8COpPymNzq19uZ8Sti
G1lghsvbpWRAI0qEKq8QL6/Pxajvp5M2UfBoBpnEF0L7DRkrQ4q6atWhdDlE
Uy5fqs9CtD8G8Kk9/ebGRhvce8ZlxZJbFhJiCL4reIVFM2U1zbjSHfSHSV2c
29ikVxgZhzrEmgDCpvRvo/Zin1RTutTuwLKmN947yf44QDysSp+TJweqlGtK
DjGWtJZJALfM/tblC5X1mb+x40C1UMOONi7EABnpTgHok/lcSPm6VX4nq3/S
kV3lZx2iYnajLGFyg8FWx+08UeyBS7AByqZBp6mqbMgaC33ADXAhUhUJgFK+
paXYRbmeW5nt6etwZmybS4fNn1i5e1vbUAoB2BiTctnXQDZ6KyR4mdUJUbdo
AUnf2Vfq0pmSOf6/Z8CH33bkW0bUFODVHEg7WmKQj0eNzUAyVQgbWktEyGzD
gmG7Iio/1vGIElaJidYoSJHMOtOHEcDr+qXWqLA8IQYt7D+uiH0R/XNhajdo
+Ip2K72uQ5AjPf3VfRfUkOU8pHuttH/gMXbKSMj3VWomLKJT1ZoBNvRWMawS
qLPeOashqeo0ltLuDhiESODY6sVD2LNAVQxeU4fpV1jg3G2i9A3bUS5DIrmX
PVL9wzXs4IzFphN+QTcnfGooBWEbU7r52zxIr6dziX/NhjbufKdbhd9RBM1S
s3QgbgTAu6kgiesozPAhINUALzJekD/cdiSEu06591mOEsbrRXDNvb4C2c4N
Y8n3VUNWZot5hzkWwKijF5GCUz6dil+Dv3csNkz1ihGIVVTr7dDyjegL0Ngi
HdtVZp9ZCGAP2ogczAVnjqpMDXRHENuaStMwWfY5ZOLw81Hl4AjbBhdrDs2J
VAZkaa+ECujWY45EgujosRRmxXZEVz6/+8IYJpFAOzHjFDO8Xbo4MoO/YUF6
qMZgyTtrhEM9oYld9VH6jGvnrY+RJ+551TSMdXdMe79g+rGpTENq6gfpleZP
3Cl3+hPinO8RSoM8t7czM3xXu4Uf27R5higU9U89ifgK3ZA+7LZ6fOhW2CxO
kunIdmAQLD3BZzkAhswc7grHz5K5tpC0bQyLJbJeDLwX2tttizoUjrL9+Q9N
Lvqe3lCjeJBRctJIOkR/wClaNKepfzrpcrpwuuT5ELkbyDKlMmdEZ616lQ7D
xkffBKKnlnfCxjnaIXpdXuTO+4H312+zlVYV/yruPgmj6cKCHSjOq7KXo/A4
R0e0rDYXQnysaDXzAfXOko3BKZEjz6sU6NUKcXI2TWD1xEUe4mrTdPZWWjWc
bsLpSSo4kmis62kA4ZOI05NV634WSd+Ir0IWmnRLt8jHIwOEGoArb90arIA7
zsLqlHeJxHEIPp7q6y24hAJ6XqukyUSKORE/4lqF/U8GfZn+/BSmHDiW473r
Mi5jecjL642odlkJtZfJnvowLhVZJyTcQmGN34zEUKSiSWT2h5ccwWcaXwqC
tc9y0aqZTFV9BQJoJ8HnyQmj3cMsVgBCEPoWKZ1a8YiMMF4UChTtwXj04jXE
leopaZyfS/UDV60qTH0jMCOD3S/LnUcPGfmkGMFsZzz5LrG2BdV0UU2oGD99
X24pdb6BRCVgtuNgAxWHsWnkmwM4gjdzX2kYY1F9XFQKuAJRJDrGavEsRY4H
mnEI8vk7kQL74f/9V1VNHshIKcx0UaVyZBA6ClPyVGSBLsPqvUv5hL96YOmS
dEXvngCaEOzU6RAeGGL8M/4zJ/R1qRNIR2HXMb37GpASHbtNQNWbblwPg2b5
wdtyKaWVO7ZGqgKqkGYtvDg/nJZ7qwpgpdDJduceFCiX7Nhkh9Nl2ng4Hv9a
39XfkI0fkfJ4LgIb08OPK60FEMR8Y9iZdJjACeb2UMpBjvMNBbgYwa3Iryc2
8UB8W9NPBL0KzKf1TQskOqwEHDWcBkNfqO9/qXI7KIKnn0hUs3I1mVbyE10t
wuMg3RYBCAOQtROfJN7xozdPZKJoKTe1+pDtOa4T0jv4U30QqmVCr8FmHoc0
t97mQR9dDiSCFYjGvxd9Ky+vss059sETKVFPLw44eBLyGjIXI3ZVL3IXr2+C
QHxl8paoSCBS9zqTFFL/9l8g+PdBTynnbYeNbAIkoxRBLm1yIcs0wrhCshGK
Y0sRmv6NOYfUEV3oP7wsbK5a6nkDsdbloYoWVZBndDOP0YGwAmaeczP3fl3E
Krg2HCm4ymbwZkz30fKJWoykOS/2dVkaTk5i7q0gPDPzIxkBYKQ5v08joAJh
HJJ5A/Tui/XO3pnCgFExWOap49sDBeckgQUoCTawTfYo4kgE8Z3YavMXrvQD
MYXq9sg5LPvzszaB+SHs5XAngxlwwDgf7dHdU3CRnuCMOvmSMA7/LQpa0uim
8W/9+jNkMHYrOTeDrPp5wH5cm5TJ8jO+xRLpdyNMZPsw52Lx097xlBmZ4Phw
Mc+ZwbBFfJkOhWMD9oBXfkFg1J4nLT2u9ISL3Wd9p3hktvRMTVvvFN7clHU3
fSLkIVqO+u3OsjDMe0tVwk+ztx3jlOcRBTJ8B3107HLJMH8hlZKRht4r/bn0
2dXmIyWwfd0Tt5nxxiyjVldOszAkDHpiN+9HGxfycjtx++c41bQ+sLchIK6p
IX5M3/JN7P/yrsUFqVswgJgVWH0USUvaPsG1+KameoztJku3PrQ0qu2+/xuh
ra8mNbJBL1XAHX1glwYiO1dSxXysDtoYqZ+Xw7LBZBOLEs1VOcYwGALAVusi
7TCttUbZW6L2+wgvIVdk8RFt5V1LmyxjtPTpjdHns59PWcXM7BCykCsNx0OQ
vc7LWYPgoIJyFajkw4Q7MuAENPkvVcl1gHbdvzZawc5WKijZGYf6Zoa9Rd9l
arzmmK6ukeZCsADOSkoqrD8KdNzSZVOTBU4u2DHQgv9kaagmMCjd50Co4EdL
w52913JHsNV1Zd2szkEgZuOh/C2JCuMq56x/ZkERpiDeOxKRzF4M5Dp822fT
A5Kc68tJUD4O57L+3hVv44aOcLASetVtEuKujd7WGFMEYMd6wo88lkJUgfYv
8tt60aUi5XH6e1JcUs6WRQVgL99tmQy58bh886iFkcicpu9lxnH0NfJr5mWH
BBPLm2q4YEDyMcDc+3iNvlqNmdU5kbdUdQPi+wtKo/jjzaucU9l5fCvOP501
/oRmaeRTq5fpMfLc3LWBg1S/AZ+FH0vdZHoSzDyjSp410soz/woAw/t819Js
G0wrGGd5moAGdYjdXDzIePUYD97qg5XeuS2q3jo4lazo0ZAgw3PMQyYXa5ir
oK87RXwXFQC/PrHbPxJRUyqdl0Uk9dycO1HjzHEpMTm4kRzSMv24Q7eCmie+
vJj8scV5OIdKLo+HgpCXulWoye9KbxvPegoUVicSl3U5w5Y1xA/ZyMnlXKNK
goXpZ9p4xe9IBDmTjnbSrAm8o7P/7mMaLtkLuW1p+8hoQllBJqtnJPJI2Xha
uwFySubnrnnJQz4MLKXqR5sL1blKzPC0kzHkNlGu/0q5ad+/qwuM0+vQ67vZ
l35k/TddmW/fclDkUUPkzc5fb2NPmpE00qhTupWJOwKJPUN6wL9lWZFlvpQh
cKjhzqwYk0aek2YX9GH096+6sE1g3ZKn1AZOwhZVaBoVygaboIzMrpsAgaTo
Hz63Em8h4mYHcyNYVlZ68hQkN0JvHsBnow/G2RFxx1p0sNP/eCQAtYwK1tvz
kRqyB7IK5PTChkoep5tMZvXEgNZZTjyf4f4+mSHy9iEs45Fwtxt+sbS3dCTD
WNsqAftAuHdqdyznqar4spQ9zqMstxEHrBPYsLucT2F6gHGilpFtPiUJvqYh
VA0JQwNq4l6168MbkumY5ghthDGbjHfM3R2HyyKkvb3kG4x03WxeTpRi7oM4
fImGApd4kzaYnmHNqKxHrvJ2kRyTICnFF84fN74ZrBtkXxDQY8vXSZjqh4aR
m7Bmqjv44z68hEKU87xbCy0vhWy2tbkIZX3ZLxc4D6cXsn+9tKNt1Og5/Q+A
1jFiWF2XKvf4MSOz3wX29KBqEqNW/vjbUumsE85BICJUaDHE0sBDDoL+doNM
52sFHwNKC3CcWyt9iGONj8Wjv2dbs7GwfPk7qt699cmYKTMi6rYI/nMUy6ln
hIPUHZNwpRkVLnFB+Gek4eZt7P/dhnisJxtsEfEoHtA7HcnaGPqN4W+PdBMc
HSTVIg9ZGKNnq6FGBQvAziHgfaVA1Dn7dy5Blo/CrE31VvnFOUBpuA+V0p1G
tAZZ3vic12AYazomMPZraXFHQfSMUfGcrIHDnu4HZHDoSAg9iaEHSdNST6lt
SWDtOrXFClm7yF6zv06N31gE5xahMN1lRUtt6EuUYXl2v2ArSYwMY/FzbDT0
Z0jN08VpNzX9CSwtPNbwEjE2qmYEwbDHKMKYNaMuqLAoGDw8inDxiNm9BymV
n+UbJm+OPIH8RA1tXYVgiCpA3SQGJqmJ7SPuiXifakUi2rMHdLYteVQ5lKJ3
Di0uS927DkUAAM78rsuSgfyv3VvwLAHmTo8kJ8O2dp20YclGYe9Ke1vyZLJa
aEQSKmDlIaRgvaLKvgx8ZJJ5ATol+X47ZAFJyeSzKKvbXsFip30vT7+7vGW5
MXyP3WNHf3Yd78CmVQuY1kNf58PYo2DzoZhIHnTzyPcqjOrVhfvwYUWrBVk/
jVha1ZZckc8BTCj5qKShh6Lf6/Bz019ERZUibmm5go/i+TB9hH/VkLZst6da
6WH8RHT42ApM1T9RxSqHWhjCU59ulcTnmSfiKuPRs1V1dOPoGtALZmrgWWnt
JydAJoVZens2bTTiwHjyI/NNG2p5Ruc4NxAv5BKpYHl/DwDtpVyevzD7r+LP
dRplH0ICYaWcbYOY1bFO13jVQxkvjfG9cIkNZTqWDahSbo6uLHc3nvuEPLHP
LGqEvba8dTEPJdOfguh1J+F6wloZe8XQT5Xg7BifevWmN2Iuzp4r8HkEtinq
+uOFPoPrmZe8qIajKJJ+wvDYR9R44gEmg/eGDqxPhY9OoCZeIg5NjhUjM2oy
COmoxMGkHp8J7fLo9zg418aP5paoPCKqUmjVGUjKk+Cw4qLDLn0cm2AwxTgw
EGwheav7SZ28mtpe/PZWCaxJWdCyE/YSeS/zZQOebWBXQ253VEnnyIZU4K4X
FzZH7aWSLojzdcOm5emV7/5nR3gO80StYr5lQXJUQHUoPze+XF5p+xUg0+v6
xMAaPq3wTrtCAJxpJCHSVgFq7Mbp1wzTeFHy5H6ILpckI4KYYGH6lh66tkQH
+4kn2U7XIsMWnrLv5+pPcVEq8NTyrmAhuLEjFeXvMQY0jg31JG4cMz1u5MGE
57+Fj73eG/hOmeGX14cjHXHTwAc3PPfFCpaOQ3wK1KloAKLHKvO4gk2xvDYH
Y9nivRkVuNLNZ+lNfz+2pzfg6lg3xe5Jgm9XSLiebRGZ5swfXL4q7QB9R5eu
fjfNNRWXF71kptOLrcrG1YyDFGFtEXxnV/EiHZ+BH9D/x8E2CGGlhNNq946q
o0RI+GxDVLuhSGsDyz6me2Zzvs7VVV6tbFbs5ynzPqiV5OijYN3UiWzxvF5h
OGftMUfrIdMOTZiNbGsFN775MG3DZoBoY9YHqKRLmPBdt2GMeCXnTz0Zh0Dj
EV8TdU7D2I0QA3lWeoeIDUYJpWwfDReNB8+LDwS4UFaiZxV1Af1FTD6rQaMN
qIkPpFIwDkcOufl7PdzcpHxLTPjVg8D67Xwp/eHnSsHX2e1VUukWnUgQjyW6
67+7040aFHqqHvKinRrBRN4iSC1TXgz9bj4+Tf74Cqs0at1CWrGt7AeUNGu4
74N4E1ZemoI7/X2K2EDW2OW9ojEGb/WJarNXFID6ig0wRzRtdLmKzP/6ldFg
hRh1snaXdQF48xhELnZz5B9PpYN/F/wdBvqeR3yGEyQQV8xl9eTIntCnZq4n
iZzY7KVYzho0rucyUbbzZLH2FSMV1VWaa9plHNhWQobug2EU3/4Weidoe+zW
yCijXNrIqJ14kl9lZLa7EbR67nhjHHUOlhIen0N5fdqFMdoWTK+gzab0qdUx
LrACXuYMN1Hk6UYXkCINvDTYDEAxb8OYJ29S0bYp/ZuU/ZEifULW8qY9AYwZ
BKJXCzSQyrUJxtfTDjjKnM0oMSxuNFfWE9LvHhGtX2wT7T04gaI7ZKMSSa79
lYgwzYuMVovIAAcKsd1COFwCvoiFMq8R9ky4t55N5//ik36aSfN6flf1Q6sL
nwM6rbS91GXcVxfrIQvBgBTJuQ3XxzfYd/SFY0yRNfj9X1RfV2JKeDmQ8Qmr
EltyqHNV1JZkGlC/bpdRmzNv2LvAMjoGyCmIynBBn8EEoxkdvPB/gfDOWCyL
nKM6gkruK9WqhjmKpG5SmE/TdjyoCMm2dQ1DnnZ5VL2t6d6PhuasedctTsLs
hmAHqOA/HFXrg4omaYtUFzJAxz1FMJZGmf/GCc/kMi1ulmCPwjMQCH6jn0cv
7orxca315OQVTICwshaLQI28rNpj7qaiELRM1OZ9LNEZyMDhJawFbk+LwwoP
HJdvHSSgFcG472qKIoyG0JE6i0KmpPGaPRWgpCl9TdabE+8+v2/ODDfD8UEG
T+zSgVFRSWBeDuN2XEEY+P06BJvgobx+P09X+yiKDgzTCleewZGFKq+tqXsI
DFXfMoeheqYebBTPq3XmGaw7rz3UARspEfokQhR8UUgelWTQ3XAR6XjODg/e
IoFrDvySUyt4YtUDG3AkCWjtbQhTv/B3cBEekbXErZKHXfEfWKZ2522+RK3b
ePkdjrfpyZWX7wlmZaEc7FLM+Nr0Kd+q3DtLQhum9AEVOftvBRzg3joW3+QP
AtWcxpaoFyCszXh1WktDhKp8p97y/9yQfuFjVWV7/3U0xHBrnGC27+C5biWO
lpMRP8Z14xUR+0ZniU3mOZsTiKpzdZxh9Kx2vDci3PlYTLGyuPrhKR3kK+ej
Cs0wUOqg+tHQ15F45ADfar3CEqTjvvOjQTfELxkLxkljYKietB7zIa/DuFRv
rCkHUJkJZgUvC7FGzJgfQMSVW9F1kwHwmOkVmfT0pfQiCy9pIzh2C1G3CUPt
96Hk9sVEywm/tMztcsdHo0RtRSrRYpocLmu1lAZ9zvD5jX5BLQMVwxtGtQF4
X/2Oev+hEdBbUNF4RBeXQueUsAhgg6K9OW/SollBuZm3sna0xeMVLz4NmQG8
WB+OR5CILQimwpD7eIhZs7FSB7Jb7iH/mDM1e2cmVXa1/RO38v6qRInthQoX
c4nmQm7/0nrOltPtEbo5ytroMs8BXCUf9oX6gNV23O9zqpSLPCFal1kNkB1r
97rJKnsXO3vrSn9N1VpJZls2TwNTFnWG0OXZw5ZCE4Z+vR3H8ztr2lI7ypkA
Zi8okPS1G2EV3Q1kUt9DiT8zvXsOESNJ0gkPXxwbtQn0kdBAFjDhHy7uwQim
x7tk73yxWFXrWAXzQywbiZE3AbEorX/3SCbqiYrQcoOrCHo0lToznH+xgUXM
ncYPaBHLUX8Osn93klCoWF4o+vCa66uJmEixHnh6eym/U0AK1y9haqZ+cbew
iUR1tgpIKxycYjMMIfdUt4/wEbz2cXejNbhNUJAKqoWdZV6rUege0A4A1NAS
DdTCDzzyrkos1swvuQBQnzrhtjw/VKITLzfm0cQxzS9DOH7cw/FzcVwmEtd8
YMcfh5m1lxvaq/mFantuJx5UPgs3tnWPCWsh9i+tA9+Nx75FxgLY++X3UaBQ
acwLr8LpdA2RCGf1fs9xAunBNYIPc6Cw73g0s/zWiMYMaN8JHa1Kh1qbYArM
vd8TyTkxLueyhhVGS7Rr7KP8ncnXMshXUwWBtl2SSYxLDi6GXeGTLLyQXaL1
i2kmWg4yOAsimSSy17afufLqYR56NOh6qbFfsYfCrfiuV5J7uHRJ9M/FTnVB
q54YleWbP+RQCx2KezR7pSACxsGj/xh6k14unausb7uGD+c3kdxDWZ+bCO2j
zJwiEweVp6DVOWyhE6VZrkK+DxRjndHwUsXXloCvptzPszXLUmJs3dktnhol
b2Fyy/in9FCEISfgRnwtxtFQcgMH+lOsrpO7I2GqiHPNkBih41ZxoNnJv9RD
MTIcqbQ4nMruGx0UBgr1/v8XhmsCilq9bUZjzfyerwlacxkKqHlVjdiDzn4d
wqTha6nZbUcPcZq/Tb9VJrexpg==

`pragma protect end_protected
