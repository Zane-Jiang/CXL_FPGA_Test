// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LK09ruivl8UEmeBtCcSeMSX/KFUy/LnVyiWl9T4z3gDP4Dmkyq8GqkeYavtJ
z/ARMBwbwDoq0WpwuTuYzFurxtfn/r0X/9No3m2Ms/bPsxLOSd1aqExVA2mO
ELbCD9YIPkbymzfZounT7bRItjGVqtiYCJ0e+OgGfdGhvP95RyXCGBP0/SB2
MUJ+QUmtwPv6mFukCPIUaV1VV0wt+0CjOaD/i6TqSx2SRH2xXYjubgo/3R6x
VIkQs+TKa5ng4nJ5o78TmNsAtlcLPgMrJycgAmQmBHNSOui+Q/kALiehRzMr
mp88ngn7/wzb1zNIh0bO+kLSwWWv3zZntlJrvsTplg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
F2wgYXpUAcTQWQsSYkU6LMUDyd6g1H0JryE2GG4M+pCVOx3isTvzYrOa2TEk
EYkdPEbfYpMn9TbwAwZ9XuLzbd391YzxsYyYjvv4R+Sh9inxSopm2LZrD9PK
BA+Ni2kmHjWnk/Ohg7IKkId9XnLTSP3qMHSHUvUxwqbfGQc28FMpro4ggTt+
lbz84C4yZ7bmGafzBna5uiRTQajFq8AHCqczClKlxKhXsWj0PlieifPHn0zf
3FI/g67/dkD32+RqGoVRAyGCzjFH2iOsoSk0N6kGo40AJzIGVZpP49BkHmil
lEWhmHvKb6rIPMdwdI8TWxxvKtIljlS/yt2ZPVLxUQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pCPUhXI9+WO79aVBLOHvopw5YYzP6sNtUy5iIR5Uwh+Be/laNF8QHUUc+ciI
Ma95LFy9AJNoscXlmduKbvYW0jLqNFV6Zg+l3IwL5WIvhGcJ6OyBLghz75i/
BQkEGl8DVrjXuabu7SNWaS4Gkll8Hrc+sKoiT3nqxM7B3467ERIck3UM/MpZ
tdJl3oYgJUerAxcHjdKkxAf4rWtFkajSd1asi30tKPP+1v4txwRP5MLsDljR
+Jo3fh3CmmflLn3pVeJaOzkTpTVP6FdOW2MHTyRTksBNp8zG4OtjkRZb1SWh
xdO1U/SHK8BjNBtJ0VJO2bXpDLEgL/1ow6zKt+cZ3Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a9/7XrNZc2lBM2PXYWFodWRCSELDUch8fuQav45XUyxMmQws9kKSI0MR4kRC
BTInxgJK3b3yNvtDc9VWA1ETjCmoqLhH82jET5KXmGimGWMqSIdDM2ALTwLs
BuWvE8sj1hA0eYk5R7g4VELLHgsL2uqZoCni5e734iR+EkUuvUw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
v/4QTITb746y4qj1AyZ4mA9HOiCygBWpSIWG5ogwEoG8AD0tF6j+G++AAILi
0HMdtm+Qm6s+Wntxtz3UgUmKwXgDY97hdzOGFlzrSag5GrOSNI6XfckHDiGv
W51gMGY+91Ya00KwYQJNN1nYNIIn81fFRiexiQ7hGqre7Jb8qUzYxBVedvny
RSxtedIrl6HLxjkhCWiB15BCQRgBDMe0nmghoiNnBdKaRRncduGEQF3NVe60
KSWThAJqzJt5Oyz9OOOZ4R1P1nY4czfd5N2nnA6ZIHo/mu9EI4QJ8oL+qXDR
RMvoAwKJGk2/VyAHtd2Dowk51jK07zcQQBKTKVzJ1OpjYdwPaxY2aw80w9NO
Iuzx2Ni+132hjJ8F93/owD8FdnYOqn5hVs6xJQinSyu2HvprKry+ye+PeTIk
HKwKbx7fgRapUnhS/mjfsIW3Jwf9P1Ubt5hbku85CxLadEtjwCaHSmitUBSv
VHUI/L1dKJPOJWuuAjHNKOeOymtnhfuV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qgMOAUEyAlDGHKfYmPxzWJHFZkgvUArq5fnpivUPPYE2QCAV8oG0xM8sJ54s
gpFc/uC6l6mLcDQOsT69I1uXlh6gMGiR7SeQnI4xz9rrY3U1osth4YMlVbAX
pnRBwjIvAEVeNz3OYh0hoGFCBMV6fWwiCGlcasLW4mWVFv4/w2o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
o8N9BvP1BHt4K5TMn39priiYbucI4awED7HffbTZwEdRA+xwoxZM1fekGinH
muskFYeetFJLmYv4sUcj3mF4GguMZbe4PoQ7YsgaijRyry2JCEKFmMhucD+9
+ofeXSGg3Srjkka7aL5Ke+PME9d4NrUGC/TiACwL9ISSobY3oOo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3648)
`pragma protect data_block
nKq2EXzHTp5/Sw72Pyz8+gLUJeZ+hnQNpeRpbRrQyjiwrSSb2W8Mz3nQYFlL
tBNK6xYh9SUCAn/KCD4qzirHYwIjwKCa2zgyJFENVwkpNRyjFrnW2eaa0oHo
ccbllvUhI0ObEoBonyWvPMOzmFL+Ay1hZ7HxAGBvYq+ONJWdN6vltXphuJ+8
s6j8cn0bYV7u2UXuqC8sitqOxEQ+Bf0G2aRNG94G8I9PJDZ7kqbOCBYVb5pu
XMFcYpzUKxA/WAIyu+VIuiaQL/puZmOFm+0gyFye7RFb/++r1EnCGP26qMzf
s+Xb9cLFXuFtoF5PqHDZhpxpPekYnDPj7Fi9SHKnv3YqeM6K3/VxFtakqhdW
njf9Zyu3VaPE+Yl1jsvn41r3Z+SuY1vlTIJTOx6+3+dzf9LJFVOrrO7HWOMz
VkJSEDb/CgjS7yV3CoNXyY4LARqVMzFHK6ZRbJasz+7uY+LGDRcnj1+x0Um0
2LmkZf9r+b1WGOFu1SVEPymwTjzKLTukmFr09+hbdNMn/zDgaGigwMDjOMY/
Mo+OChABdQIfOCshWqjDnSwYZmlfWHqTSyIyju0tIxaVxZUvY0/wytSAno+Y
Cct3ItRFoJ7CroFAsLYAs3DmFWDTe59Mh5LUcSVteDc0SHqp7rvbgqTNiy+5
dTQapMV+Xs2e7jLMwgXuvJqeA2C1I+54lT1ZoiR5HZOdP7Nz0OF+b0TPoNla
IWdWtDF/7GExqNlHpuyGHV0G9wdwRTobDpzP0LyOiQELo0bZ4njIusr/a+VZ
dgr5903pc9qXBH+omUC/U0iSb0kzj2LFVY2skKSJNY+SQNsqO/h+7OqdUXFR
zHgoXUj9s6Xo24xAv+xinyK7FyxiBaZczi+oUlbtYTdciBG6V+k8WBfaaort
1UcBeO5oSZ3cQ22TmEDvwagKO+Hf9/EmumQLyyLHst593uJFSXGqawHBVsr8
PIt7PGhi8vKvl6awphZMDRP2FlrQ0Nltm1i2JoiP88fWRC1M9PG57isb7J7o
FRTQ5K/jxwI5rpWF8RQaeonmdmUHtdFFpcj9Xk/SgvuuTNCdF/A5sxkhqePX
EfNdRTNCB49fukeQDpGsGN1PBYpvhHrOjAjsgb9Js9kOX4hc82umysgyCdUX
Kv4hoU4QuZ52BBNNQaE3oRRo1uyrxskS6p3TKi80F5gEL6/iuHnSSoTjtAJM
jn6slrLN2lcRpRU9m2fN27KUWWdqtE73VJTzrtU2OauxaXz+eknl6epkY7Qy
U8oRFOoFRAqllhvVumQJBVVTomKfWsixBv4GJR4ThFLyyoFt+6nfktXLjQAb
YIx7RMWGbKj38Z3wecT80lfuKOJLAMiccVM0lphqE+Uti8vpTLz8MzY7GzUD
3jmk1GySRKk75KL9WqYtRyrkf3m6KCs7cdMR3xWwN+W5UeAnXCd6JaAWQe/p
GHkgpkeRSaeGRHFhXfSjuaLwvqQZSJfSQsu3UjvIck4/4julqOAkoO255H04
GYkK/XtA3KEH1awhHR1EnwcDPvjA8uXWYREKUuiAzc1m8NNv5Yt2mmIOhhwg
GNXUxQdYe2TaQAga46GsoBTjTajaxPkyYBmRWQkVoKnbsaJ6dVrHErNXEZcL
Bqu6lPsQYU4aZozZPz+cy8bJXlMdouxYgsD4I86A+tZFQHvRGvQ7WvuPva62
VcMxLXnUm7V9qKqP81vB9oWg+svqbXgb5jhnXEekWODzwDDO8HTauG/Ktr/G
EidVdJBBHnR34F0vZADmiGThGJ6/fzcNKgrpRni+y8xS0Xn9yQbDKOiydUrT
glsBJDCaNOJ8zJIDr/cncw4uQqtRvA04ECX9HMHQWeTGIuoDSJphuHIy1jU+
Rs04zDzc5Gv5vVPI2/eml+q84G43dGQtotDUE5MXmlXi/Jrx+36Svcglkrkk
MZciByNwlM1mFEU16wvnnyWIILqfs/eY7AlITCVzGQwMLacUSGC7lbiwxV8Z
rIttbUIt46XXILEL/FyNCIqS3zVNMZodl37A7HXzg+Dsl42iIclZv656BG1+
LjXHJNHpaHyOyAwXfqjyuWsCCUZZq1XGHpq4IKt9khm2P2rnOkBj6wKPtrVf
qx2rl74y8EXm31RW0cMpG3TjaAZYhl2JxU2oryp1suxydWS4Ft6Fhaq6HOiN
phqXdVcNGkBOA8gezszqETaM7Ofw+wLtiU6kYi0hPLfyk/u44H0/6ozHdAto
8zZQwdGy/HDuG084Ufx0NJyxMMqOHHVM6lyd5oXxkJQJTsPhtZI3Yev5uZPk
0mMhZ8/lAKYDqkULLA7nxuRptfsXS1HHTWaSuGIP39oplfx/jEEVjU8kbGeu
Uja+jkyLzUSgKBozk3AZZqkOB/5SZ1BSTy4hSZ8/jE5yd0/11q4L7OEGLQd9
IKuTm2XledVwAFtoGY4+gIOB5HS2TARxuhfObCNe+/BhuyvdVIq/lt1cjpsh
Sz0Dil9Ia7jA9SgtUcjZqphd2j4F7Nnd0pAFgnO5iy/cet56xuUEelTJCRQC
KNcQyspBaT3FyAgk5faD2x618YsDUelAreT1kkRye0Awj1mFa6Pv6P343J++
KslHKpeQIGqpEfCSe4xfDlw0MwNNIl7uRoTluMzsXceiRyRmR8SIeIhhyIZt
6HrpCmPHBf9ZHE+3eW901tKtjWDXMWPYQEmYcC2/NT/IwdRPgDnakzUMnB78
5Wm6xNU0/TQfg3XIsHazwTLbhR6geh+7Ri156cm3OCRUESRmh5sV4slk/Vd4
8Uei1YTqKu2ke8rQggdhIn8VzF/u3nzVipKyFpmfm55eTrOIvOUAch76PEvI
cR3YZ0csZses7S+aK31ZrhiQ7kByncvgJBrQrx6G1YHkg7Nuxrq2FqsHYPWq
A8F//FxEHcq+NcqIpx5JabJ0qi29WpAhilN+okpTALw0FE99SBvZA9TguIrS
Eo9tnWDvgM6W73g86IzObI4iqHsnhRiCeMZN4OYy9MuB19crUCGbSLJ9Upg1
arns/JEedZEwd7uN1YahqzPBb7/ZT39dvSFKrL+OkgGvmHoNniePQJAxMmbg
zRaCD4+sPW+u4Nxq8y7sV3gOJc9NA1PWlclXF45W/9nhknOHlRK1fSBGOPRX
IaQ1nlKjN5CtrEecoa4McCDXl1G/7IX65/MdgjqpVDHKEpIM0tKTrcMuy3zn
uzibRTz34zDJxb1JSnX/Rg7sXvmSoSq52y0/BmCGKSFVmMpBGApKFSo1uoAm
2c+dbE2CpGoK+2XtIA3qTySAJ2mndNxtdRnNdtDuQWuOBGmNK2CGJP1dBdtl
QiEZDkv+Ztfy7fRQnk51o5IfYGIRVeleTutOmok3Lt1j3be+njfA3LP99gv0
MZ+oYDzhrpLqE90+lqOm3ddm6Ont4k46BBRkB3+Op/1vHYAn1DMTUwpdlwNE
M9s81j+u2wlA94tVNILe1d4R0UJ1HKjmypXL6mI0TKBAakw8ba0v4jSlEEhB
5PaCza4lmiv9jUkb18Vu+eDrPm43VzJFT4FtPzc5iTT08OcIZ5x8vR3pgzOv
HESxFga897Ag2w1stHtX8N3v2yqGig8sFfCQqFcda3SqRVZGSMv1c9Ve2NHH
3o3BiqZYw22r1WNkBaci5SO3KxdfXhwdgfFVQkaQhw193pLyxMAqz7YahFTs
46G2PZ5ZU8m9pUlfdFF73Km+IEHjICtY3AQ22ksFigYQlOnpktjUlnIckeDG
FcW0n+LjMUek5lmobaks7DTaaJSoMaAr7SVQZAJ5UEYzxweE/ZJrsTX2TIQy
A1FDydhzq1Gl3S988doigBZBeIc1yMqmTn6e7wa0IfUNXzy/vUbHUsIACRMZ
2gxFolBoKTiyqAWkdopclyoPhGA+y0xO02nsFGA0qsrRu7sd9Tq/VP7eLjmJ
a9rEzuI+KpG9c8MEwW+3I1dGv3GYL1MpnVY8h54Ha4VlGkdJOAMPeoVEwQpj
sSuZWiDo26EvV+5NRmnS/e/CKCzWJCSpOXD1f6jzHaW/olQoRztam5bFAMSr
PGZwFI5Oy9X3HBoUyoopLtbNK6k12xP1xDOXbZmRg2J/7Dwu6H1KXNOZQrza
NM3QYJoBTaFKP+TlyMtVuYQBxDutjNG9qWgZ741F4+fFwf97xUzU+OprEXeZ
L7OLHtvT4xn7z5vPWcvAGJLRTZXM1mRV6kbxWGiyP4ij8efgA0eEf5cN0qT1
9lqPoA+Yp3AIIREJFRM95pOgd65ZZ92NvHVq9lHy78yaHw+8zZkUFtCd0B00
xxKOMnSULqVzZaMaJV5UI3T8H0n5XfWgYTZoGFt9itstE1fsnVxR6FsQL+p6
k6vDGLIRSAiKwX/1etqZP8UW2G8uV7qRisPgt0nISUQ9uw2+7jHpHgnsfb6n
aXhWRH1EmFXBMeazdNymBVf5A/hNrSTNP949b2FnK+sNQtI+e3s9vRwWMME2
Dec4rcFaV3baC4NxPhXpdILNUFPYJBk8qYhphl3CsfqCSYhr4rmXdFQpWCnn
VTnn3DxLo29jwLogFyF7fs2iK4UQz2Snj+gW8kNyr3Ip+QGDy8Q1Tr9YCPT7
upkNQFCf6xNGlhpcEmR5PKLyWJc2zfemt+rgeKFAXWxgpn8yGxjrN7tNCZcv
+LBugDM/tBJLV4up8+xTFDzjSc65SBEcJqvLM+islUZBCZdqZWm78RSHjpvD
ZBR9i5fzngMUlQmC6O3s6+I5xRN0azrtXY/SLIYtS3kRyTjubirYoMQBgskh
tzir2Tob7nccbyiAU1IQMzboARw1OpXrpiDTetrgK5PTmVAnraTkQi/XwZ+j
gzvSaMxlIPRyy67e9DYxevXGVfbl39HTDbknd7Rw41V/Hu+E8oU05nr7hOTc
jFTs

`pragma protect end_protected
