// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Bz4UPMbS+BboD9VQcBsdFuwbsu/q2ZKYLWZJ4nLUxkQalWGZIn2wYLfKsgXbj7Up
F0YrpoIq85jRWBKF+VeFWHarsnr6lHLW3EeKquAGj4qTPpyBTcJrGkZrlviLh2t1
ibHA8/QoIvSyB6JlKk42zQqHEF90Mpxx2lb6ZUJBhDzex5DBCswU7Q==
//pragma protect end_key_block
//pragma protect digest_block
X4OmIG61Ki7QpPUSSUdFn9hTuxw=
//pragma protect end_digest_block
//pragma protect data_block
MriscUhOKMOeAiLQ4NTjMEbhI5PCt/tNoQGZUnOsf4FYXm3YoZHDTVtSv3wvRhke
r4ApDK4l2FHZKkZkUfcVSfOLiYHZ3VlyTGlVI/e8QhqJnG3pOjrE4hjzUPVn/Ld1
d+Y7xxUeBUhjh382Rw9u8ukZlFuzVeg27673NKwHRQf7/z+3Vl4z54fp251/+cps
vZorPKMbcNtsMEJrgu7NWgITnoeiw9Zohk73VrV1kIRjjjaa2QOYyFhr1Glmmz+e
2AJZD0zpVKHjf+eCsTK5gOeQAPJEK8mM0RfFQnhO/b5tkzHwF5iT9cOB1Fdr8B3x
PZFC+xGxyjQ9KxrU+BkFJiD3cFU42kWWi47ZX84ZUKIZ3TMj2tIHtjmeuUTDqSEv
/qnr4ucdgkdwWLMRVyPyEGPIS1DBchYatHz+tBDfS0eH6KS8H+i4dDqLj6fmZ1g/
1vCoD25JEzE4vUBHDj0464Zw5QU5bemc/zTLR+vsGowCLsuUr4MTxEx1TGaIf8wb
lwfD3PexMqXYtGwUFblJWEzHuEyX4rReyvubRg0txDw1n7KdbObY5ZfmVB2QdjQH
euYTFfxbBenHgtBzIc874UdFfrgHy3w8cxqGPV+/1oCaw9n+iYsZc8Gx2rjA/jHW
io3/zYhuVf9FKaDys35aRT/KycBIGMRvkPsQIFHUSpDi38uCINc/4YCD/n/SZ8WW
FJ/fDwi62hRNcSWtfmzDQAF/nK/9WJ9zWmmjYM9FPiRuGGZWyD1Fo2kmQu3TklYm
jfHDpv0Zv4NfGnrQkWXV/EzoGECd4bHgjcL2A3qgry/EyD1ZFQ/cn35Ngxd9CSqu
+bf0U16lMsiU9KizKfBSLTjL+Ayb/Dq2V2ZwTmkMBvu2Pqwc48L5WUARh9fvUs8f
rkp9jLPjGTi7meAUQlfaRb69pnZR18vpdRWJX+1smPqRv0gysDsrjwzYEmYYV5cZ
fRrhxZVTHcH5v8HcDswGPScWFeDZElIWAIwio0lgeTLwYUCYwENtoJRf04wFS6IX
pz1dySzHvVW208W/6dC9HDslJCO/NIEQol+EV0A6EdhChdO9DeIWcufyqN32WkSn
PSdLaZ0755yunjD+hk2yCOU0fj5Dqm+06otiobKD5KcOud54mspJqD2bzSlGQaoQ
m/zfs+H3u6jidb8OkVKpm/JIyZTjfv8XppvTz3RwEdWCcIg/hsfKC1++qyNs2Qq8
YzYho8vjDzZuAkyowMlKkXAn0RHZb/eiLlBs+aSCNFMpfRUCjqV0dNJAB+Wu8jdh
APNPIDgCKBjutKLxPjI8Lo6Tbxaj2gD7JVoGB4m/ODAVBLpJprfZiB+W0DMEa/aQ
tZ34CN1U3TykSSqPd2uBWFfEGHejYNZb14/dHveXp8NOC9/XEyPXbeRrrMnCHxfE
XHN7rPbVdIHi3LY+ZSZ3yGBUPGXmAtJKrmc4p6UBD12yBmqDrW36DNw7vlvEtOsJ
/cHAvmi/BaM2PFd+xPf0nQD/wC+1/hjzeAbEMZ6aM5KqU4OKuxpwL85HFCvQGnrg
AmHG6R4QchpSrRQTOLMv3BpPOJgec6VByDMS2G0EYat9/OMQZBaTraTHqgJkkYf5
IB8/Nb2sqnWz4euE7rrIzf4HQKdScES11Xg/H/BOPaFCI2ll7l36o8NXOHXg5c0V
hSvwXSew0kJExvNVeGkXe1GojipIS/yWbUabxmYjgWsDWDUVCCDKLdQsJkwtWeU9
G47a+LeXGzo5pZ4/aaC6BU0ZPtqYhVkejRuPdiJDys8OoaJUZSpY7AbjTexbAaI4
qOzGtE8k7p47ykuVAnVAPJed9wYxJGGlNmrq9kVEmQL9rz54c98L8qvl9e1lPuIE
4nlPcDhW6Ogn/0/hpNJrcKXl0ETbJs9uG9YsRgZDUDU/iFLXJuyhgdsJ59vU0ihc
OnfQg+bUekUOjvw/7smzBXxiL3t5ZyCyOB4LWODZT+Nt7NqroOcUKoUpk4eR9qJ6
HHCGdCYhdsqbHOQuhQH8iifjFCIudh2kkv/U9Iebt3BHf1trUkll2sB4uAW6DphE
WM2VK4EREIGVZjKuQmg8ATSBgZaD5MxpDOBEV0Y/2AcT3zrxvSmi+3AH6zfM50gU
wXUUFfaXa/n6H5zdCH31eKWacvLxGK7pSvSrc77nU94cR0HhJOSVlGbnXR5cajWw
dWfvRq55isj+WolMqZQ2hQPIm8pujjjueEt9dD+bTZsWoYqgze7boM8j67lyrXX5
t8r8L59UagcykSka/qb5PaSQMbucnFwXi2bO0kIA+SdaLVSdY8eC7VpNOWsHck6m
b/TplKhBs0X/V7FF7L081H2J5EAFegSoOtA8z5Ge2o3ArU23vxpd5MIshrmkTukX
scYWBiNgGflIBLgt0w7feGp2F2ITwZvrEK4l2Q5fKsmerphiF8aAIoqEjhtTj+Pe
w8PzkbmwAmuEJDksyUeaY4qZhZKG2+Iax1YIxmOV8EX76gR12UJzZqY3JSC6TFMb
HmGjllTU6SgE1S8fHGwNTx1XBukngoCTMvGUFL1F+mqjNfan6WvUOzPkKGF4xX0c
kEmpDP7IqGMOLFuMhFBojua2vLOW5XIsH85lur8pMDl/cL2odwF07kiaXlfggnNB
SSXxNEdMG8iq1ehHFuzSKl0apgpwwxcf2wsPu25y+DzDh1atUtXo9EKfi5dYVdGk
U/OnjvQHG+BxLPiWPt9U/0Vir1Y6itra/onFsLL5F+PxTQJTx6Lf4avzoMd3/4av
MKlhnWZtpk9/MGrF/ASQtGCFeAa5N7gvAk6arNY7XLmuuJBudq+WoNCAqMLgRv4o
TVaajqMDm1qGopuvUVl5Q5/EF8HoWHQwDYpFVL3lpk2FUo8LfGRAKgPot0sqJoeI
yK34lx++KWL2hwbDSISnRItDCazU6YxtbgwhXAmwUhzY96DYa1vuwRyfiqZCAJnG
8gV2V25hxxYToXG2PK1AmyAsHXPsgOHsZytz6xrd8Lps6cviyGX7K3EuG+Zqr7bR
QkOTsI89QYEmE9IHXwszFlhsTCWzvnLAG/1v5jXEcI2dyUokWb9iZISnWXnTPRVb
/B+4NSl8tHe9I0ISfQH3CDx0nlogRJBEq+AdKXLVC2NXT1aGsN0JFiHc3yMDxJqD
pbLXItVxTR28fffT3EtzhNuckgIoU6EleyfiIL/KhPqipwFQiVtzN6dNY/QhcHFG
8czbb2pqqwYAzu4uSEJskIgW30qYwuebjWEkj4hzrfY9+8O47iWczIwLxX+oK7TS
pDkNxqqH3dbrjBbgFq9EBO2v57a/efq4x5/m1p9drWydNRz17dyBgnmm+ChCH7my
nW/wWuhzrt3XnH1PryLSvYNJB8tKN1B7ABnyVGpVndVmnwdesgiIUuL0oWTs2fsj
bQjV/U3RoY7s4aCzWH5IQwfuHjXogijKfE2P9S+3bxsSjf1KZNolyRjPMnwc0SSV
tQ+XujAsSe1IbFV6Pe8WwWyWtJsz7bAhJqlVJdggzNlUMPOikppmrvWh+/bIOcPC
JGI119p0pwts2lW3SJoesEh7Bs6XB4fOPueaklEApyKxsORBfHGOUZ1Dux1owe5U
d1z3tcJC2eLCteRts7Dc4zz+aT7c6ZhSOaTK9g6/aVNnzSFjJ2qB7n7cDse1FtJT
iKDPNzKlk6pQCXcSmNZ6w+LWrayjrsXHZucyFaChFdjh9dp8E+7FZCHd8928V9OG
kbmEK+sRpbut/FCV9qqDeiaFc+7+kd7QhSsP6vKF3dXtAWCh9ybl+uTS7o8s70s+
A/TQxhXOrYcgkXm74/WJLTotRammcR+tS7DVAx5+4Ui4wivSa7Tt4hDitLKrlIH1
td+qvDx52RFOzCqHReEwZ2tVpnVO1X2DvPIHo24k8mG9GAu2P7F/uXsO4iCKFDAd
9H7r22PIA4JkZHyQQri4J5C4Ll0515e/PjGq3fvkT7wG7DgLwYQvxw3WHZgKDS8B
A3av9BeL9qSj9bJz7d3PGytKJz6vf/0VKm2Ms/zadHc+GkSRGaeCaynItRibaxh9
XV0tCUd/NT4Cwm8g1Ul/SjGWDGfjtI9/A1aRe/Xu0NCv7IjDTsx64zCZScN6smW+
+DpD2VPFVy7StmC6BeZYZlknzj2Di/cO0sej5k0lp/kQPjbBErk09oBXcfMQ+Wac
0pGffq8XAuRoq7TNaj3+OX2pLSBvR4gzuixZyEU4CO3NEuPSLt+TnreE5rZ0uZ7z
NUHGdeVenIIzNZntWGGSk80SOb7gZHLt/OwtFcEP3hV3lpocBq7YLXwnoLjDmxau
5FPzGN+pbtJqBC+nEPc1ipntA2ZPlPVZgyZuSU4Zs6JTi2By7fUjnAPwPL9YxuuR
qzv4tdw41Iy5bmuFy5F4s06GFdoXjRfXs1RDfRHeY9AsQtG1QMJn8FAw74zViceW
OMPyAVYT+bfGjrYLKnZCOCy/smHJkGTtGmtXlWX3mVBZizws7E6i2Bg0QfDh/eUX
iNFgEsyEtxolsT/iLK7EWOgTp2OauKnj15gd5aajQcreiwnpkIy3DKBUZkSKXYG0
RZ4U2tKCsrz2eaLhYy2x6M84kIH6c/8Rx599Xb6DM7NegdDZqy5n4dpbKTHALR0g
itLHFou/IzGTm3NX1uqXdMhi6XaGe8awtY8iK1thlLz5zxcLn1ew3gQFyQBjY/9x
eG/E3JmTHMvAbG/6JSJJjtiQfBmsnc6gaH6jGINLiUzC/NiltIAktLlrOwn7ygZo
nOWl6Ah/53MYxdUQx/j7aXeVoQ0h4gy2Z9bjUpbzjqfG1VewBEIkC/KDz8hXEPm8
RImNkhyBBCNe5hS5jFpK6SzaWoznMh0+DxEIuTYtu1SH8b3R+51nM86xNScMQGBf
lKg8/t4BTqhSQvEE1Qt44pZsmZorW9yZL9XeMl4x3dR/H7X3eadLF+ckzAcM/4Gn
/EOPAl02I5ieX90LzrlG7yJPmdQxdb8IkmaIQj7Px2OlFYAPuvAqv8cusGDkSnyr
uPRrzhzeoXBiDDv/3CtjTsc2JSA9F5z/e/ps0bXBijLOYnu4w5vWEtLsUCUqC/1x
khuuySR/W9ZACfwFvz6M3udRkAdJjtDGX5ZZhL1kYE32uMzfjLdfJPRngSZC+NSq
CzS8CCjTy/SrnfHNIrLcqjsPVsn1v11h0fd3sclvd0N1Mu5HlWXURpZjO3k1bvNI
cm+PqxW8u2SfHPDRl5EqsRrju03PpzEfxVnB/REr++FSicBzeSUp5H9m4ldpxAYx
FkLitgxKxB+e7T7U1wmhk3c9NvmiMaH9WNiqQ+MVa1dW9i5xZ3oEKjFFGIUpxDy/
seoJrqaZa2+vV6VVBc6sB5yr2U4005QOP0moyphF6tzi4qGEomIYy8TT05/0qORh
tERGYtK4S5bDg4zvM0e0zLq1X+XLAZM/SG8hRWdihtancQoQ0aRygVDFUC2FVGL1
qTuMLHhcwCVn+HN48xIzuq5VPrZnJLDtWFFmQwD7FkTbQjUcdnCj2FJsxqeekOVB
QMbfFFCOLCIFFmVPZ0s21f3+9HWoqe/tppC4cuNTp+L6rJyhiVehLlTzI1fGqxQo
LH61aJn/2x33HQgZJWHmJJh7nxeroO4dgDjhyVipTfk/ka24u/lMEawxVkaOW3es
IuNE+KFCi962KGuuM3Y2HgxRxJ6eIrlW9xDbWx32n+P+LX6pu1wTJA93ZSdgnb1O
LvtTV2YlOJmFqvVD2QyA0mcgar93wRnWHfgxamqOPQHEk7SuPqMptBsvOzY5XYXR
a0zg5m57LKauiapw9cSmuGqFHZ3huvp+pMgbxoLDSOTd1CmtYPdUqij06oFcu1Jt
LFFnPRzoFCP59m6oHOsWSBT0gQCc07v4bDnJNlxu/KRpO5v5T+pjqTURgFLMjj8K
AzJkEC42uJ14LohilQj7TxscZTGzqs/MCFC1F16+hXya7tP/Wd/yFnLSeZUR5k57
+a7zu8OxNFqFO4BbVXn/Lgiim7DKGfkujUGabxu/U8BDZ5aphVaSoL1+oKSnPsIJ
8+GHBQ0VvVlyGvpTMjiK9E/njg1VrXeSEIbfO8fnTt02mO1VvE9174DzwUN3xvRe
Oh2ROCw8AOAzFROd/hGzetjSwdfFcreqBHxFWQ14FiaMw5vbVp/UED/K3oe9YtH2
a4G9MNmipr/h7JViREl0ungrG6EOAp6rmQFGyR5/eNwP14hO0Tk27M4tgiH5GwWU
alTERm63Ud8NE5DEywhTKseyAYzCpGwncxbEMdxZbgqNUzwQhICIqHcEbsmC+74i
Qg+mReKBgEAfQd2Lpr4wcxlFXrEYGy8EvWjDefoAV+TGeKXslkhpLbNPRSVJQ02r
61ODi/mLd5FmFUJGGyZj7hwulKCgot4E+viuigTBj03B52gv6t+OcYqnLIxhdqHa
RQIRITHuWSzPqeMLH1Ta8wjIBjP0gFDVOmqZ+kXvOaHE/0vEjTDj60zet3vfXM++
QmQG9rbVCb5qW+H1l/huD+tNP5OmYitoJBFJI4qbAVA0k7TpwBuCvPt5pE90LTJF
cQXT950Q+sNxm8lFfHS3kNa4n/RQqSjgjXxMqkDRcxiB7ii6ZWrpZeJ5QIfHU6o4
X+x5Rm8cDymepGgZemLNqJvUUrVAtWXglPpBXIXnMD5xxlOYEwQLB6DO8wRidtzN
Ge12V/F3SmP03hVL+ydYmbPfRiD8i282l3TNSzw2OkQTNGxkEb1D4OFkxUbCTUji
I2IlpxY1rtd27t19y80z2qFgjwtGYCOcUizYjJtoLCnTFJuFjq8gkgv4LLe3heNW
GHiXIzUOcWIhacqDaz9vDzS3KRAX+XWXfwDKQlJWlgYh/8mt9gjC696KzxbpUHIK
4Y5AtLppaEsg72c7Ih8TdDbC6TdUbSsCzw5/3RgoSY7oyfhCW4wuGw8oCzom8RfS
wJYezMGOCH0TQdgK9ALh/TkGNjIcWux5IeprjLG/xuPOIyRRJnIUOkBCqiGqJ723
XhEqqaIHcYhud/ywlQpynxa18i9011O55WsyCRNrvU/6p2FjryAqHBV4NibzgoYR
I/wYmt8+zo0Uh38nzzVHceSV5V3TKbl5b1SaCZjOfzcZXUjU2ESBz1SmJKBL8oml
800aTt2e47kRDm84eCdhFpPg0Da5rZxTlx8Ticw+DHzTnrN+vBUx29JW9i3KiUqH
k8fqGtkDUXh+LFhNT6xTLP0mrE4Cfx+6Hjb+16gJz1xf7XN43McSK2NHmmtO9bAW
8DDDMmnxn7h7cSfCbPssdrTUdKbGb5uomOBCJhmG7QjVWQx90BruvWvgrOnwtkfj
1vouiAFa68D/QvYHrovLvUinTT0TJ76iDpWvTfNnLI6DypYpwGS4LzoLE88Vj7tc
qQVWsnAvrDzUC3rFskcb1sXWBt1Ml4K7JMOulfu8JdnBqcvlOqcrwu8NiDnLzDFo
kj57WJ9zgcqLF9U8BQBnOFWI5ysqJFnsinGNt+DmT92zbBioqb2NtXbZT43mRX7O
PlJBu39khHn/PiWdyCO+9wtQiRkJQBukmPHenH1+ZKUmkgEBd52EarE21hHqET9U
jyxDbFkhgiNCEcgdoW5Pe5nePLlrKl7vcbZPRbYsEwOOqKzMsY2p8W7+MrSkN9cM
w6N3AM5oYY0K1+pbufMaA5XlGx/wChQ+lAL/oVwqyb9OgPvENu0bEsscRol7pVYe
2ZGrS9nyikZkVyPo8XPcY8JLJBd1sS+9IF+umwYFTWcdgWBzK+Xrv0uJmHWC6L7a
AGUCaqUqOR3hBMO4ymdA7GewB4n4ITP87VVda60pSsDb2kQN5URgthEHwOku16oq
7EYbOhDCCM1EPOtl8f9n7JX1fuIZVgAkQWJoWekuTUW4rjdkcuthhDZ1uZZ9cND0
PYnRJh7+9rdGrwLfbSdqLTH9OawSJsHeYI2Be4ZleDCnabJVyeZ8eUDPemIqAq+I
xxKIXFrOhip/UdxLIlmZKkvJFbK/otgUv4VAbPa4hANyQULqDHvakOTv3/9IQ8FB
6cZ8UbZVSFJPgCGG/dncuftIk07+5wW+duXrLLXeAfw12noKsqiizpaxJds9NUtu
a79POb01YKdJXvKzb69LuDLHLEZHBxqPyTEu9tKeKeN3C3nRG0ffKM8XxwzLWKfh
8S36Fj0g1PYInclC5MGqZf9/oDukNeopU7/PDSX1mav1jd7ICwRKY/E/X/YIwa2M
R6N+uY0Rhz8oE2WaVIIAFBj5XDePZFX3Zxc3DAmOPQOGjhQDKpm8oqArk9Se8kp6
jwIPhqHBzsoqKRsNhtSL2FJkw+Vz4yrGKPfmNX0knjMuy7bT4I3PZGWg0Mv6gD7Q
1gFtVS3lOw5p4ODEW3LpMcmrtIWHZ0L2ex6vA1KeMBDoe57QlaNTJ+Z4TIK48zx7
mKNkFFx4vA8BUl4qFSH8ratK6CwTCMiNP0JrhvjmaBX6kMIqRKVTurIytSAch8QT
bAoNPjrIfqOE/GmlseN8VD6nfJmj6WIMPC42JVEvtJwnznp7lFCCp1sSIoDq2kGU
1HHOpVlzlwAixyoZ0RSqZo5Lgvram9P6gwCKB5S1Q9498Fea8eurmtOTw8LVh0vS
PdBSTUsx2sVOGKW85xDYtRU4dpIOtCwNFxYIzRM61Fsm3D7oQqbCmB21Px+tZmLz
YxoMWcBeDL6aK8rjtMc3L4TmHa/a9eQigLhET0HJF2jeRumDzqfYdMItFOburaxf
nKdrM/f8LkOLqH4fJq7m1FggzfjA/s0ygqyJjhRfb0kvZa0O3XGp1S0BL0J+QKTL
SDQmcoOFeECnjNtBB6FMx87sdz4keo36WcXohmSLs87cS3Xr73Y3Lt680DVlK1l1
WMunoXmktBjJcsvpdbgjCvj0RHyFsLC8BQ2qxQGtoTnD0qfUdqNfLdCUYrT+fvMe
EAgETHHDBqoOYbtWNaEJbeMhFUgi3jI2kJsFEMc0jAqw0GDTFH/LBFM4W4hMvMD5
IkH2pYklHZEn/8A48aG4nexzAGGHTDADaxDZ8xZ/VerAuND8zStVsjs/qfxGLEmf
vn4DClAyKdP7ht2Pbm1PMEYLqDusHeptHWQTNMr451ELsXS1YZ8rCZdjUnE1u5hk
0R/WW8V3cLj+mUwZC6nCeUg5cKs6czL3OpNPwBdMGQPYD/A+YRybaunq/2ciNbaR
f+XgF68jg+V55yXl5ocIb0KRKJGNMj63st8Y0iORQ1Y5lgRxqPLIyh2Qzm9FNQq2
2SyQkqxkH1+FPbXXX6d/W6DvhXmdWcwFsPf3azbIGPkO5mmtL64pEhY4R92qA5vp
/VU0PpCdAYthL2Ap5qerzzttNGirWqcNqYvgcEg81YzkILFLSJUSUVPxkL9wyMVt
lKvXy9TbA8viom1ozpIPc2PAbqn6iwwe8vcblchdVBbrA79jTL7ra0Enm3g4fj3m
9ZuZxdVxPHfw26EHSpA53iyzLjsjwQoH8ZRao2Ald9bAlW7JJaxJcwuSp4CF8bz5
dWiqcmca1u0MbjK2DfLyw7B2ynqfu73U8WLYWv6m8W/UBmUR4e2uAMEXxLFghdVp
W4i1nbhxNEUnstRaKGdsr6LeGdKrnLFnEmx0k3HgyHLCs2K/KW0bPjC/mZyyQaDL
C3l8bV3/FFCcLkytKIIANoHuToKxM3xifXc2ppgNOW4YfVHxFShV4i5MO0XwuvKC
oXXQi5llnEGJ/241m/f8jnehca7YS7uKiA9sryF0Oj+yekowKtmSSlKeBlLKsXw7
c8+5d2NCnopW21w3j9EBPb6Uj84ZZ7xNtEjIS49QVawP66KILmwTsRrcRWNg2WnL
VVYygqiq5S+WuwjlErinISfvfMrJBEBDLEgyiXgO20chKXhzJjjP4ps7tgBV3vMd
2382dugCAnDLTnP+TYWoM8JkE5Z0cwd1uRHi0rL1S4TJkcIqdn8Edhoqv+bZEXui
jzIxeBTtkiGKRtFW+LjVykX//oUkrn4JAiVPgRLYS8lyZZCIoJWVQavesVkmsHTQ
WOvfcWk42gMTyM1U9dm9dqBsZxlw4c4koIeDCtz74OdVMNRXpPLsyHp4CKUVe1hv
n0PFplNMA63+iVXKTGx2FcLVUySn1qERqJxHUkwkGq8MCQRkCAwRoHSOSjpLb4Dy
Gy3+IEZLn5OpVqw10j/MlRAJAg0GfCdkJYUoMhe3ECEe3ZLseaVEzmmjPwoVTqjy
EhGmyE3PCWKgGt4VnYnwC6Wlr4Zx/sxHN5TR3PScY0BJS/3UsAqz02ZrSGKCc8Xd
nXexRatmxf9Q7PrSCej6yteUOyOdNduwYcjPl9/L2Y67L2Nbeb/ksN8l/ElwuyLa
oaTg+k0EDBYw32ntR12wLdrNY8CSnnRNZu6zm768/CkILNQq13UmQFtgRDbPoqtD
agC9ZaKRIOfiBWN3VG1W/Pbbo+0cIN7bnD7zWB/2Snv+ZaMQNogCwZb/ij5Tvrwa
bsYicCfBOXySx9H7hp6pGe4Lv3z0P+Ec3006XyE8DmKelMWp7z2k3N1DdVp1Y/rr
S+ILaBVQl4hjLWgV6lZM/fC572RIEhig4lbWLDHr012mPRsBwxxw5DnyGiV8GmmV
Ss0t6PxHt6v42kZWodlIBx6wJCM1IKIdVaK79gztTd7xG6E/W/45lLS0PkAphFMa
bLmUyMD+35HPyVPRwxy4u9ZreoUPfL1BqTpQa0vdUGjS0mBE5X37qjMYXriMjiex
JK/OwIIkYhJHuLgH7gObfa3BbuzX68YrudX9mcmnj/mGUChMolIiERebuNs37t8I
gyRPA/SA/Nyqo0OZsH6Qj6uDB03vivCsA7jkF+OkkpVcpP1vrbzaKLZ8ksTU3hl3
dtK9I7a5E2NPmYIt0T9HXJDcVj7MpDBqgULl/nAK6DWxNi5ZPy8DOea499IcM5VM
D1zXHNDXWaxO/WJrRfBwItm+obIXXSNlqBudMTUVSEvhaRNU497FACerBDqW/czm
5ED5DmAPudMOhOWqf/xxTxwgOxUmIyecL1jxxsZay/EBhaKi+Dc/L6FKo58SNhyK
akUegQhNFFK/M/9jh9sTCagDCPMLgRvr2AUiMgfy+8a6QSL76nA32OPKWSF7SCQx
+JyXhiAtnxPaWnFU3ph25KfoS4sF18ZwBmficI1hl8CjWTECYn2ERkA1MoU+M7Gd
McL3xVHFGvkTmtc14YTSw96arn/KdTq6uQnWo+tPTdGsDuF8sklsX2qYcOlUh1of
HEUXhwJlQIJuOdMjQifQmE5jsxYrbTb+BF/Gvx8equHqOOx48CY/KD5htjsBhSHk
hwae6zMJUh5lN88qvzAzSDPwOtDFZD60z9fXZvMLgd443f4aZJcCmgsOuChT7DxF
0YNjQDKolfvMNeelHnK91F2aR5NRtbxcww5aZvhWRsmFDVZULJsPzes+EomNhjvo
wsxiPVY0tvTUQucldpm2p60lRPDVHv8jb54UlXgmii3YbbMVswlOVArTNZt43r1d
WdHxsUcNIjHGNFVgYj4+/qwyhyVZCCdzchWzQ0tvWRkpyXFhcHLcKfqwO3+1RhBV
/UA8ePuQ99dz3ic47hVq5iXUdM3nGHxbNLuLA7+op1QFM3wAbTYJ9lefKIqXBNJ7
JhvW7HRil52TenzXekTkcne4v27IhuCE9HLoI7bvyHTKedOrsblctRuqmjywzLz+
ilCJJfVXNWrL1oCW8bCzMBK5tnn4tQ5n6EOc2Y9hS+/70YxO4X0Ieju2l8TaCP2E
wz/yGzpKsyXczR3aSaIG59gwb3KeQCC8a8iniclwFnuJkM/7ph77L5vOvosM2JEh
KsGsoXDr4Us+pPxLLHbutg6ZNjjRZZbEVWORXMC4JzxvLmjlS22NIVFgmIoo1mvB
flVtdZNTih/AZ4hkTZJzPyF+cwzdVVPpfKDjOm3voSGwzhKqd4VD2XXeeUdkQXKV
T+z+++mgsfOFCLjo6V24+CzSek26NBHwlj5BqZPREqQGSvd9Vkt0oy+lk9e2oCIS
ClIBFC5UoZE+NaZqeMuFewT/wPZ9d4l7ConuONV/bjH41DIiElKDE/XPmO5Tsq62
gYCsK7tNhxCRwlkZVjr5tU7Dj3O3nVANtVZmfgWQ4GFjq1szOiKG6QCeICoxuOuB
CNIGIoVC46fj3MsXgbWDEcsvyqwFjJgRRMwFAicF0U1eNF6DRQU2BOFNQQXGy7RO
J4lsgm+IILzfyoDkIHOLv6kVCTuACoxVUkNgu0kDLoYJ5UeTt9KWH1GXjOGFy6Fo
HD3DEVGsVLl3w4oUqAKjMZfDho2V99Hrncsa6CWmPQC1B1bnxiJH8/fLez/CjM7W
ZpO+cN3qfV/Qlzke4Lj8yxjnfYjIP0lGpdwkRCsAfdn48aaG+XnsoUtfJdT04yCG
E90CTcApyp63HjWaHOXfOdKyz2ypZ0mgiooQ8Od9S8BurrnL9dgQBhljx1Axsh6B
6rydSxauyTLYHrfnN+qBT+GBHLQyQaTqrH/RWmE4W9inKA/zwAX9xrByfww1OS7F
KYlZT1VxAw3TEgZtHmFGYN4aCrBK6DXfZGcspCom8DsnEZEcCJfJOfDLxMl/xqSB
xXzA/pdI2ut9iU5rSQN8+bZbYlyhViCRuIM6kZjT8T6zWuHtAg5+ubTpe7Rb7pEp
tN7ZWg9Q8Ez6OGdSeZpxFORGvZSsjFoNodeFNcyp3ewjYfwvoavX/Kp7uKYS9MUe
eA0OhJkDRrS4B6M/RTyQcPJybMKq+ubTo1I3ru73KM6RqsnZc3ai3lHitwIfozlw
8DY3TnIoXpZmdnKiUUc/e69wawZlhvvZnAQ4KUHzWmvqsgl3HqYbLWuWR996pqUi
cYlBZ5gAkGYQJjRWqSW9FLeMkVG7HpXx8vImQ4uF+BASJ23qxqqVjjLNMgYHKm9m
xbXTP6KGdZEnEDa5kOHRmm2NP3FR94KZN6LuSbgoioQxe+jOLm/5FDRnfCE0HMRI
vqfTQFLVFUAFaUET/3mgVNL73Y8xA65heJiXrvLZkv0WgNv2IelGrv7tVCkzMWYe
Vzg13kYzXhloGzwt3RYKADcAb+7BC65e2u641GP0Gb7XV2vm7t+QAfhSdej8AT++
+3Wo0a0BbWMTNwsXpsiOp2r2LfXNrV++FlY/aJy0oh2QcC3e9eguww4iFpxm+eZT
bXJctcCnF+D0D6MCUc1sbfW0ZxjjUMcY0qwmnojkUj76ekhfKufqPnTOy3WqPWyk
p2Fv4WShieT2Xz1EwV8mkzVFrY6SHURyleb2HVMfsXUQBEy0UuRrZD/T/3u7dzo5
tDTLVeI2yaj6qMadMB/BYFmbZpXs1byVrMFqX6AOlNB2uNYef+LhXvMMcKUG75JW
PXWhl19ZzjKv9vsZ0erG6tqu7ySI1m9QLBftMLwuEss4DSWRqXA1i+s3OFAKx6cb
MNMRBoq1S4VcWaU6SXyIQjYcdOTetWi+BzpaZboP/G133L+iA6749pQmD+waB8Gc
W5x83Fn66Juy2oTE5SAdiGG3JH82QqerRetfsmh7CIAKgpJ/0YzQCcpPmCaiseRx
6Bqfqo4M8QeLp0FLNaIOZhq87WuYi9d/ZDB0Bgg1OO6csm0NqoRcIBqzFJBBovle
gl35SvaLvoY3ExE8w6dAEH9yBpFpXgQ7aZ0eu61tmgTwuY03ipBsgnIIcs8I2RAx
L62HwWIQwD9A/hUNQOI3K2+TK/eokSOTXjPSP1VD6jG9DWG7twfFoJybLYRVWEyG
n4jTpVcJA6qd8jXkbsGR/UVuu8amDzMsKe9JlQVW8zwc2SP/Qb8artdxREGEu9kI
Tsz45IWcIPrl5DWKdgULQ8FJf8ZK16hmoL1A01KXcCD+r6uAwsalxqtqd5syCQW7
Y/RPL49x7cUReH/GktRSYRyCB7Wsy0CiYRufHMjDp6J/qxzw7etcP6FzWm6/W9s3
PK3CBJ1EnS+dz9OhVpDkLTajik3+2VFtj8gW7PngOlDNHXNIgIrKiSSKkctrN1TZ
fMptsdzr6ne1/wHNCcX1lLU5w8/k6NaO2KBkDHYHZG6KmIAuGvfOB2GJy299rJp+
AF7YRRXA0JS3PfayzrtXFXayCG1k9dSgRYYFfj5DYXtZQ3qLHNl2l4i7bB//F/RK
IOCuoBGMFD4ZOvLHEzwseEH2X5s2eXLAZMK+tLY1uH/rUbLcSHMh7U+LOaLbyx5P
q0AXDgm8pkZmTVoblHtZP1pJEfz0nFat+OpEPKj338+ckGivJXQL34h6R14iC4F2
BAsxh4xy20DjuY0F48PgvdRTFP4m/i4mwtJEb6+E74o23PQ8vhB4rL8XFfdzpj7l
HBOgz5hgsjh5qZK9oIJuiNb2NkdvnMHt1kYyhAX0rwHLGLWDw8cNIhY/QjjlrLZh
9xfevsDMvAXa6QC3jrb8qSAD8pvCiYxZJw52FErXxPqHqT2/wH8JUcaBvBD9Aqus
s+7MbGPus1NdM/O+b5TjBUTYyZmKjKRgu1R++pp6AwlQ+JexU3P89rkCmx0uM9Rf
9VtN2ZhL7y85Ukb/L7ALvWDNm+Msnt0e//uElKCzzIPH75d/NWz5iq9/YgU8iLrw
cOnrFbfam/jtpITnooQHdJp0UB7upVtDTIyDVfvf7DhJuJ31YQUWWM8MNGheTYeu
92s9+EC+vNzANBm2jvxljLzfpRbqlUEZC8J9ZZGUdHy4veSFvSOrFdpnwy7NscO3
aiRx7KfrMvs+ZASZzbsR46nEA6f41K2YX8dUYP0Jsq7/ntv+RqkzUP+fNsGlEYBM
tXVh+6HPHhvWnv/ul2BcL4H7GZVZ87ogGJq5mUv2WUFjNt7wjvLJuxHzrQd1ngOM
G4U45/VqZCZOjkxfDP0xuHCQ9spjXEizsyb/UwWzeAcO0fDtNqg4kvgRZOJ+8Sha
HLhmRi9IkEnkXeYErOyFaJCRvl+lIr/5yqiFjOpPDt+tduqFRnb6zjvdIVv+/7E0
sn/zT/aU82irCeg4gegUXEN/+IFRLRgFx293bpglqPRsFdRvM3G0qo3ZLDNl2KwP
EdKbSJdyG43kmMU9D0J5O8pfOkS1h/7hxBv0xTqBhn3o8dpN3bHsNvRx0buWkl5D
etSJteUi/bvDMGxBHL+GIOYRUGchTR/7D28mDhbmM1HNqVS3N0pLlpM0wYV62zzL
4ytnkfOmTI+73B73/42SPBrJXpSe3eBeFCsM6wDm6jNx7+CEJqFZa6DxEUkz5eI8
zFxOK3vuqW08cPyRDS4vJdlifPXLIXlhwNRJWIT06QG0slPGjuoU11QFcaDWg8zA
bF3zFoE8Gn0yeAvAFi3mO+GobSItQgnC1SP1AiKXgympCW063ebVLKcRA3RvCArA
NVzBA5/enJ5TkTQNiZIUDcJ41gnK2Ux2ahD6HNe1iP5VDkdNupTACIO8rWI0A9yq
vbJltSbhnRfUjL3coW5y+ElvdJYsdKQ8BOXP4gGcZFo3hRLa7TXDTePFDB7Iugca
VpKlmWSjXOcq5Wq2i6MpGYLqzx/1snmZDOs4eZflfauT54Cf5GEQyW7hjf8K8Y8L
CxmrAoH8d6OPQRzXSmwOZsD0PGNQDmhB/gUUHcKjlW8u8+K0ulfvKDCGKPuwLnO0
WhpPIOLcQriSzJqE2gsHaPSz3yH0W7pCi9EUA7jZYqZL4DBdEh8/O/px7wyzKwwk
rht9HQmAf7/np+7k5D04v38O3iw0CCnR0AwJMkWUAKKjbY1Q1GxdID9qWcu8DKke
w4LdBX6n7IcF2dlJD6KYDHyChfY5jsFVrgLRb36w88fvHQqy1ANF1UNE2JHNkn/Q
E8TNIGjzIS2NT50Wb2ceI9vKRoc5r5baklo4Unu1O4irlqN2kATDiI9Sk10501f8
/oKmLRpZXQ5SPPSa2gGFQf08Joxl/JEm152l1VhHNYzPlq3r+2PSEa1vTusYHWCv
5mPLTYr3MsRCEK8OblelLKKLFhqZ57J0eAoFWDFeZ+R95cfHVVwdZZ7GvMQeO+Xy
ofvkoD3X8SOYUfnyqE9LEJshsuXK4uN7dkjQnqB0DfOntqQUjtvJ33hNS2rEkY/T
oB7FZfJsMrbVHyfdq8bmeBWKG4Zy0VC6YV68ZM2kIn4GgcBUd9ZuwO67cbpF7yQ1
TW93qXIfN1t4rowtfci/+HzdtS4pwMlgjEUa923um6mAxfSyE6xzaSIfP3oMdw67
Ce+F2Qa2WDWENxoyhP/6V8raMIkz5WAnjq6YCygTePDOaEu4pQgK1c7Km8bG2CGv
XAALlmKdH3x9YRuda9JK776xUlkNfOkz3S+p6A35Y/7F3G8OdbHj4vJEwEaNWjwG
P4tUMZsnBT1QUt6QMA0iKjQbUiEKsSNWv+SN6bECdhOLhMsZb/i91HL5xFr9V8Jf
t/4zaksBIPTaihd0jrCIcUmjyb37TCcEiX3OmP4uYDEbUTnCjl7/S2okVCTj+1Su
bFY7EFcfu3tbRWGlyaZJaQJiCNvwPL704bDjj2NkWe0d4vUWZT/xTwx491tIMGh/
Yd0XAyO4yIRiqeVaINH6Ptmqb2IW49Uilvmxk05U5Z8A2cKdMGGJAxabvX1ncPyD
Gc5WFAleO2dPpQrn7DnsutCn1RM3yn4VrX9wJ+nqraqbprN2U6bDSRKLnCqWVaSn
U8zljircF9Rt9Injz6rIv78fqEmNUrrKHQEp6NFEeLqtLJXUp1OMQ4PBqjq2aEzM
1hQMao8VykDcHd+N19N4eZjMpWld5iAibBm3Edjn6VvohSEhjNK9KOQKgnPZRdlc
zV4E+0mPSuESpDVVXw7llNu7GceVQhbR2RpH9yi7VViO8rpz7LijfSXD6RmgN5fB
fnt3XNqFv4mZEnAKMcJ7B5GKmwsaCOFfJDEtnA27q+MXbBJ4/aOAzJ5ELREmugCH
PMLA+s6aYUoia/n94L9nb79yFEbNQFsT3Z/G7dCbu5DK62ScCb6gQK3EIFdNVw7m
p4tx2Pbz/qYPLgf9nx42hdm6jd6sVNc3TyQFSA3v2Il1vj8WWGdGkfp7kVKNFt3Q
4iOxhUE81oPiK4WIbetvPfXQFQsaZfVbM5ylG9L0LEthlBEBYNWm+q/MWikPjHWW
IOJNB/XS72KTWeSyRpNoF7LUb387JzJ2LWHfw08SnEYRK9BQBm1SNmdSq2A8oKb0
SNDkNUw9WCRooy8n9Dg8DQG/ihPJbGLh8hr/IgbZBBkR3MU+KpoW152H76/NoCaz
VMfBUpnCUi+fbAE9btqlhXMcJjNuNDBLcoteHvCynuPBiHRDdX/SPPkhcfcxucdi
Voyl75cpKavSKxcw5sRlqDZFtPKWHFTwZ2mmdipic9+Sp0MgRZSsnn2lKD4gAnpS
8E8/w2hv7ZjvvAE9dcXxU17U9QW2AxwouLmCiaJSg0wiMZMC3f9h/7BaT38mGxwS
W0VzS+POA7I4cYvPqJHIq0Uh+onT6VrEWJ5pRBerTGKk6qnaDQAUsT1PW2uQagQy
/cXAoYuAiH8a8bTQYaiv/2gM51+/wf8zILAskfFOGNjuI7Ro11qZouJcpPGfSYK8
7/J6yDRgwjWHxlCzdYO0dJ6n8i8/T+xn/ZhCzfJH+31WFNgHx/26eCu9ViEaV4Fv
juBIqBhEPbbo52Zf7hJF4CIgfaItaxDYuQqdPaN9ulil6+Luj9bem3o12NZrtTXO
xP7W/xmegD/Sk+foIRUcJrXFFTNTbBXtg8iZjEQsGHIxd8myhNJnct/J2TUJmIAU
eQdElgutgrUa7nO73paQvlUVOTfq+1PnfYQ510bYk2vo/jsZrpeC2Y7PAh5Dpi63
XfIbMCXBLrSseNyo0oYnVTjX/AGlAUH1sKx67qMiRvNwutH4e7Q5YgbQrGLKbS8T
nQNggsUUXjr62MOcXXsajCB19u/QEq2kerfTV1jbHu/bImzol47xDHNfAXsRo5XU
7khLQOzc3VvCFo4NJsrv8fWGyiNYDCIoxLyHGfD07xG63pkDP3OyN75LR3Iuql5t
FnGsOemZgjEBqG5cMOxh7TOZDNHsNA4i1Rx49508arXZnFFUTlbAciGmpIJD4m0Z
v2/Rn7z+19Zcx1YHwvPm/gFJMoq7Uw/HfN3UwTdZr9jQE2js2kXinHXT8cppp4Dt
bDIVPQNGZrRlkTYyhCiXpNmHD/VBQuFolNSVNTcemTbCYTfRtUYCbFGbG9eg1JPs
1/5eM5F2xpWSt41wdPIJt88Bo/Pu/hR7sim6jSEKvijddNIBRx0O5q1xv1u4HPsq
WMwBnG78O8nama54QU3stMVflpZXp6VVorwlFC91ZB/qOEeALKdqXCtVMyrcH5Pr
ell9SVoXDH+8BwGSZxi1sJT/mNpA36fcqDcztvjZYOeKsN0cw6h7W2lVMZUqcIBK
hRhfLoPXYxNPhK1MZfMeZ4ZK/J70g0Odu82EICDrWogUSfdb1aP8Bt2qlRRcgsjg
QuEaFNqDyriQF+Mhyc47v3ZcZPjFPSJKYyNMOImMYgzLlmXapNyw1gRqVsJ25nLZ
QRdcoXSZpw+UenEkz3diwZ4odZl0TMS3GYXMz+ywV6XMQBKU12etV3/2mazHIC+A
/shckLr/B8mUFaVDmitXcwrj2SYCRNcvbMzGxtYU0fjdEFaQ0n71xHOLdkocBMkY
+7sjT/A3dsKaL+I/Pp3DkZeGgFhf67L7/erHwkQOczGnE8cLqrKV/wEmO6zk5dSz
OCZOuPeB2VrB6YedtterNW708JzZxp19VoBllrxDXcKo9WqkPkqOpc16JBWongUc
PylQj03Ykwjj+Gy17jDFq8qh+w+aWdWXb2fRtMQhZCD6NvpcO9qasWvNKGfra+if
JQRgxVZHX4Th6IN8WLdOAOTr0aufTpJ7dCEP2bsIs1bGDrnV5HhXBL/QccrQBco8
W+EuT1xaZfeFLKBMOrgpB13DjRrCF+1fZoay8AYV8f2Wsgl8i+nsUfqZSA4/Yfew
6ubBwg6iwPo3ULq4yww9MvHuLR5rQDSVym4SnwkTQPZE9V+zPRyNIvSkaZMwInqw
F44vhSw4u8/8UV+pOQk4JUX5lLqvbXjgiLaF120jlKSuW6vc5x2Ile6BVHj4xaox
yct4wHO+LJIPQQ4wyGBPFfIGvquC6wyLykbJYmEfu5Dy69CPJCwXGQWehIBppMiK
UNk5fUwXwh0w0JAUtNe1Ln0kdmAB6UKfeUx9skr1hfWvL+d8yF58AaR0dMpScF9r
HBHwtXiY0Kb3wy4Tp69/BOuG7bEWGEz3z4QvP7+jg+txEaSbGm6SHtJZKruSr/Mp
tJn9p/hDUIesEv6fUmvTf6nJrThMaDN9s9VGQsukHN0qrJHtn36f4w2xJsG7hr2j
kHJNPhsysI4XicylASGeeXLBCIobDkF8UHX8t7gDcwaBaJzQPFfpbDy5Wu6HLxkv
jEFOI3+T48ofKKR2f7xswkX5I14Kd23YiX6EjgNTAMHte9RMSmxMVINNc/JSj4Lj
eToZ5JVoWr44YfjU66NQXtZJrUzcHQFc+5xMmwvypKv/441kNBYKXRz5xDdKv8a0
8Mu85m5KCuDd2VgNk++iIe2BM97eC3BtqDdJtCN2UGUPKtV169jAueFvDKTeWjBK
2QZ5GpcUJMLFFZ9rtXpOHIzQ2yCMe01Z9+CYvtIinGLk/J/2qKzQUYuqTJoZSlOI
SDvp8h/+DA6sNsPs+wBfPjESMxLpQdpwb7qjOIlNGVMG7AIB0qEuJ/UtBHjVgc4a
BdQQTX1CEe0CNzosKhbD9hx3JB88ymJAz2RukYUW1yJSdHQrUjKdN/IWkVAQuryI
vylCUevV7D+uXwPE5cnJJOfo/Josz3I4P0pqjkrtPhpgGFnD3HR9/DvAIHQSx0v7
u7Rl/vjw/voP1IBGi3zIifo21KRMDEnx/4929STu5TYZC7Y1jfZo4lQT/jUEiOX1
cpDL5UKyi8cjbRbjWbUF8Udi461Eu/0qbMOaz97dh5gZFMa7SiuLK5+iyPmGYiI1
1ElKJAW6dJ0vKhPBMnhZcS4YXjNceIlTSzxkE9ferbAem9rqn0ar8BKAazvRZiXr
uGP6W/202wZgoNMTJcSDElLzE5ZkjPc4L/HxOJnd9O92Vgi2fSrWkBayWrR9pDQ0
TnahQZWPXkBxC5BgOJRGvtJgMCytQwvGaCptIXR6FXcC8lCKT/daCDRkwAm0mVSW
SI5tq6b7Hkdv3kbn2Ps8vgtSF48h3wu5J5iv4cwcflbQ/bdXKf9hyN4CQLSeqGI/
Oa2xepvz6FtTE6VD+NxaWaMBOJ9XTV6c9tShrYxwn8XX+4z49MesyBhBK2U8umYu
zij7S+9UpLGweTAVIF/p5cxLa59fDR/q/SwwZHyanL5YGXsSljX8mJB6WhtAbLpI
wX+idpXC0EUGI2o526Kp4bilxi0+2ynycuo12IcCYS40YDG4rJ2h/30XPEgNJdmR
lPN54lrRLqa7v5GouD0E0MUoxr4HY2CK9DtNFlFbpWpUTQvC0LZSww9ACVLMgXpu
PoA9AAHoQKWYBq8xymvqHl95nEA/0e2/4CHnmO244SoNxPKeb/jOtabnYAiNtmJ3
GcLtuf1NsfPq1Ht9ShPzHe2GU9uRsRKit8uj9yPHj0c4VwGAQ+Pp6ZTh+j22Q8gN
pvcODpXOw3EghEPKnZ8ab+O2K7DPMq8ckznkJ+TBz6h/3fmAPUttTHOHRGVGjy3+
mc0fpR0TyKGEEWV9Lo1l3obO3LKkzorshvwUcMQ/RnW2+XmJk/r+0RgZH5OyEo5w
Cdb+haXJ+5DdWd3IwWvKwP8raXKG45he4+11p0CwOpUdg+663Q1DewrNFTtVepEJ
hNi1rRsa14JphYbxsCZIK0o3IfpOlQcC+8DF1XbBO3w98FvVsBT9rf6urVYTUU66
+SRvah9/XEA29AiZ0VLMCxro6eCF2iij2xfBkfePEu5HoJ1q1Sbc/3Ifc+MI9ylx
mYGzfFqj0SNZiWFr72npAcC0OrEgq0PTppA7sHphUJHCMeCXz6ZYZMq2bvtNDFHX
MsGlhFjd5V5qF36CdW+kzw==
//pragma protect end_data_block
//pragma protect digest_block
cH4JzyNbSnjeT8kSBgpYO1mt5FY=
//pragma protect end_digest_block
//pragma protect end_protected
