// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
gIbYSDohFkEHayPa6cOzi7iceEJBk4XyyNdmfoXtxK0mcdKL4XPZbGX90kJKKHty8MR5vei+RvxV
PcKje/Rspm3VUV/uZh7KhKYDHQ8FxjaE5DoDJvdAVO6GI7VU36MmJ1ma8X4pNywS8o4Gye5qbV+H
Ly/NktzshSq0rGfs4suYURHgT19V8T6YfO8Ie6Vq2HfxILMTinx6kXt5pFBpWKCQxTnMpGpMZGxB
Xjot9ShU8/iq1o/KUI3f3lCwOWPrsIXLXZpMql8IaXuhWa8TWlZMIFuOAq6Mbm+KjQ6QQDZLgh/Q
5PURncxGScwGmtlj8tgu/QJV/BryOehgWsVtYQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 81456)
+kQ15sOu72/UpNUgHBq73vXNRm8Lm3i3+/Un3wHEZgcYgjZp01XGpDD2bzqBEqpsO4ExnQRpxjAJ
U8Q1YgTvcktfIwUskysES4RhF85Badhlu37A/PsBC2b3uKjb29r4Q1FD2MVr1Xsnyt7KBf2jmGIJ
jYIwZ3rXlFoVc2SU151gcTs0bwrIxc0ArTO4RKuaoKNujAuiPwotfsmL3BEdKcUrpsblaq9XUfj+
j9XETZ1Qtj1M3mvgfrydn1qGswiFJZD/bGEnCKpr04v3JytwhTqQWN2/qp9K6MTXjMf4NSLXPyfr
JgRX1ZKsWiiNPSNceWNFr7hmOv8jeRQ3yExpNf9redm9V2troh55/Tme7UYywhyLE3Lwd5T0+o2h
OgcQDbqQtXWBibNWcT7EsUihl+ZDDFgGk2Qzc3WcELfZentVcNnSmK3npz9UlpIAxVMRfIdIUis3
xXHF4lG0T1llXzx0YaueDvxSoUGsWHmy+GJS68YSWwWwMzlwG9iyYsmiWOWb68jmgl+CrGynadgQ
UvJnsaBhlfp9xkDYlQ2GzqueruMKM0cI26eduH1VHfxBMZ84D/n8BuEkmrr1h2kVti0kNSc9DDT5
6s0LZfYoUWyoflnRLE3gjaOxdOuw2CJy1mxwUKKc9fQvaZmAYgtp6FEZJhkkBCXbXUpArxRr29vZ
ZgAMCuOd962zduW0EmLn2iNov9XnxY32SIlEFSHmht5VobaCwCFcD5LiPN5oZ8WZ5yuZctEWQrCU
wikwtl8HqKziShISD9CZnQTNbe7kuRjMsnFvfBDe+V9cwb37ZyYmK7H2MX+DTFE+eXof+7PDJtSt
6r+PZutQDWkUE1UKJNKOLBXPya05g55W1UYi3X2eD3t9oVsaLAFwD1Od0kjVNvrw1Zh/vRI1l432
XrzLWyHwx8nGynxR9cVu6sul9vP4Rf8G0pGe859Z8ruLG+dLxCA+2WUo/sC4G3rfbP+pnBzpoZlO
IG2PaoT6EGEid4YpbKHRQdr7anny6B8T1q33FeGoR45uQcXtwdlbs+XPC+NgaNtgOOmeA3XAWJmZ
+TgBW3FeE73V55jZB2SXyLzGKsmtN3MkZwuQhMfTwV3K69xdZEjs3pszJkFqk+EKRMj63fwvcGcx
NowvKvE3Brpw22cdDFjOLKrgTGE03AUlfDDJFdI5EBJh7WD4AcWsLmAtQwxwMvePtgSuK5UCcAaL
YtWIqYzvnSj/RGa6zSQvyLphcqX4qx44bpSjS+sOXRw1zeYLS7H9FdVWw+bdSSTehwVRLJUYyeIa
C5Bc3if7K6yJ1RoRr3DKRpW8NBjJHaTrCgZA/4bE+JusY7T0rjWj+93a0dvL6VcLQ5FCQ2Wvrn+f
tN/FP109StIBbYrUbnVrHSIB8vAD+4INgpXRow9/CQnmdKbg7XBVdf2XJNQu9FU764oXq6f/60XM
Pao4cv1KJZb40hWF8JWuFXl08843g4Fv9fSKjECfhwNN8BlCtB2YTKdFQuYM4HSKL2NEbf0kk40c
2QFqwfPQ3OJgBLu8wcYXaT8kf1D3bSf3dqxx8Be15/xIzpsSNd3DRGZ/yi1tHvfZ5DOzblkAPW+i
Luu/MDOYXhAJLnwGxfuKf/2WapEzJz4zs34tEOw2CCJKBwKYg3oUbzgCD0A6e/T64/0WsJYs0l65
9Qm0IwCOTE+cvPSsTgXekAn7VS3f/+ZuEy/rC8dlfhyN9nDGCE/zdo7JDvACp5feyyfClTlP4OPi
jzXrPpCJ9csRloPUgRf18WBSpOX8xh+9ic19e6eCN42pjyfG4eEAu4L2BnQQwpySbPzgOaDl6Lt4
b3rTDoAj5lpUF6hBS+T4S3b29nar35sbx2i9S9jhL+koZjAQW2pbls6lO3EN1wVGCKE6W1dwNjSr
VgE70JaPBj6zcM7xB0JQ+XxfwwbAFTZFatuBmbF8Jyi19ZYILCpZImqAHUj23jiLhc8ctf0VwhEY
VqgTkCelePzxnFt6M8+rLFyQxvIaHh1JY0t/+5yUPjhDZn3QAA5vJfVSexQOkOsvYllSMmqTeaYS
Kzuy+zNUt3x57n4hSPI9BKrDcwyGcjyNspi9RS2YzPLwUXg64KifKpFZ+oPq1jlyTWmLylTN8QMn
Q0Xp0tl7FD/FTjJ3C4kuuAuROagaFfS5Y4dDcrB/+f1bSyz1jKnn1TvxIkURdKFS8aeF2c242yvm
wDY3Q2WJXZyTHpy7+lDnXYWEiMbRlLGO/EJ6UejNzWVsjHZIhk39RyUrBKJSCZ4REsEy6s08QLLB
69R61QvO6wzTDb9azJwMYUgG7BEus0sMMiTP5ncw6R6GwanQJvGvqc5b7750q+gSY933//KmBMlN
2evV1NYpbMRYVWbRKEMDiVoqOkPqEHDKa5s2lFFdyzB1ejAqIpZfpVFGBrXqbI13bZyPD6D5Z1Vf
JsyMF7ABNcnmI4TwITBHlsc3db58hLNaIiq0s+RMuxAUiUk3SN8RPmKm2gXe1UR5kgGq/DtmDUWQ
93bZh0o44LOGDTnxNBv3x9uD5Dj/+OAZ65WQn6d9LFUSSjBcOz3dB3JKmcGcubBU1JY0+ZgSqo2R
+qhCT3xsQvs2ae+FLO40qyUQ8OzpBATVmvQN1F9wUe/lFLBsiV/EgqMI/g9tWNlrz44Iq4RvL/kk
VmA1hhK8btUCQRzKqrAh1qdPG/kjM5/9jG+fqV1Vfug46pAGM2wt2h74PyA5PQbW1zabj4qaLCjH
BUEt2P2epzkAoMrUs6RWc6j/Ue1jNRQQDMsX+xJFvRrD+YXCYl7jEf2rSJFZm2ZZFmveV8OHy+5f
3de/QC6dJEjEiYfI2pzdAhaUORh3W8iSX0nlZEN+lx2L67Gkhg3U0PV9tAJckNwQkreTEJN7ZPiT
S38quScuKBh3ZRhiJsvI7fk9v5cDWRlwwEtD0lJZXRu3xwGTo5aO7XsGLP4smRl6vWYVBQXHuDtD
8Vpc0a6nKAHfPaZYo1DSjFxm70n7VI5Ah0FJ8HWzchwoNXCQAfbweMcZVC/jNbvbTXUE48Y6qJ3F
AOeLzId0G3ptp3soikpo2fJ94pCPLyGJtI2CaAlbwdy0MWlTnBRv33MX74xdxWDQ+DEfOkaJjRrn
4q36/LM0C1dg+kC+t8zYioinfenL1z1O8l2KsdjH3cAIzLkEcLHoHNr5IHoWkhCbg3xYRwgUTZa6
VnaWbUF1mhJF6aYZUIih8ZfYXbJLMBhoMpxlo08IYKEM66fW8Og1bXj/6+j7cMi08zQAw+wLDzN9
fm9Z+PDOr79tr81BppdXseu/rSUaY3RZ9h2v+4MWP9SMEUTlKtGJ/eLCXwQPS0oCXRcSbCT3xJwg
2SE2HwtET5//yoqvCYOSISj1jzMXmeYiDIUNoQbZU8+IbcK72Ny8kA4eAjv8DfytumI7bWig0Z3N
78l862/ZGxKIG3dKjVnw1SKur9DuKSWlMYl4iwCAoMeS1GGxyVG9GtzccJOuSV5A5NhCblnmJP1u
ioc2s55d6tg6ZfpTYiZumdwjNnsIEITt6e0Gl7f1shlOKd/CLqpUVv3L7wPUpQHjKxDrJ1G9Gd6f
ckXeFQhtUoYrT0+ELxRyZpZDKT2jhboCRrkhCaliy5YAYAArvGwjIB8mMu7xV1UXSoanvVawdLHB
AxcDfqM5cffT40uiWjXolsDIr19AMS9oegnHi16viSw9/pcmd4UFPChmg/47gJTFqXl7hrgw7ERf
RAmUeYXwTpcaqcbLgIzu3PTgM7JZxPLBGhfHHegnldcETHb4wpL9UC8Um/l2GlPx+389Cf/YOHqk
A+u/wajhYDVTyxYbct0+5ogEY03FSaWuTv5x0PXbBumpxvJuB3qAwBmlhrZBBmxBVjT0cdViyBsP
D2WVfnFfFVpR96WfcuNhThZixdYfK0uf7RIMBIBI3uN3LDUijJ8M60RY2vp2f0pK/EdaXGGjGTyl
/vW3DpJzzRy8vP95cSKNujmSBcKy9P4tB7407jbg0PSna0nGLSsef1vjnCMwrDtYkc3QVIJV/nAv
3hjOJIGUNwKtIIh2Gcr2DdtjJ05mkiL8DShbHyHn1u9VAm7K2yeZ4VN6plrbQEDfFyBd4QSSXvLg
w+QRCbT487xKHv3AuJ+1S/uH/P6DwMtEUYNHyXWTbpFu72XSNGpGrrEJSNYmP9GJ+B+HSMmmIBRL
v5cOOtkmUyGkkd+nsePFQypAFgy1LCvlhOAgHIvngWMQ5I/8apyCeq78ibNxBASoGVIxG9yNTh6y
v076Wrqk7BOsO7rTKv/tGqXy5lkGHAIEOnSfDOd+wqM5rb3GjKmPK14MqsKU7ZvzAJg0WZfR7VRh
wFq+dZTzT+ICZ52Qwxba3XBEVUfEw/ZULVjq+/4zLom5mfJpkK4sSdqBe/DzTZ3itOfCa6WPbw+h
vp9r5xFamLM2opZjtgX4KmDe5lWnBXLmsTyUd9Oqy8QLc4zC+DJ/bUIUgv+BSj+0a4QXO7KTeFJi
ln+NinpMSq/qidAWK33XoCeEv46+SNKOJXPv/aL6LswlrVx6QmBROVmM7T+z6EgJHRL/t5VBZ6ag
6ZWbtVIi8n9NReTUvySKV2E8ntlUi48QAhnMvLimP7t3IMKHfniJYQN3vfV7Oh47A0Cs01QNZ0p0
W1yH/piMM3Ar8ER7v6j6hfS2jchsmqNRwAcc1p9NWoYRXBaYMOlCvmO9nwYENFnPy7Z9Z02EyDOC
drhe5UOuutiE+MT0LSPjq8Y+e4Z47W0SItcRkuPLqjPmjNUsAD0bbmysrS8foUwXRB/Z+ERBmzvm
5dwPmiQWcGnVbFcmkiuiFCwhkN2DwNd6/OJcBYTKZDQT6ARhid4dWqxb9JCogBylTgUImrGLnbxf
rmz7hCFLxpml4qkYK9B6ELJv6BhfrCYfHocz82MkCUCazPr21PFQjBXCBlVv4/AqWpHGgp9teQzL
3fIo+28Qp6jnv3w8cRYg74w0rjAbCaztBB+Oqf5h9qxzYvGarNwYCf0EERvTjbFdVTHU47CSDkS9
chJg6F+YNOoEYFhVhZasGpStq4cjqIAWoKxhJWsWi90rsWzk5IKo2Er23K1RQTu3cHFDWAyTX99j
KurRkWtRJ4A5Um3ox8rzweo7qk+fYcgQPh4z3tLyP6oDSZHBY/vbET83wCIAbVB6x2BVhXt/KgJ+
bmR5PynzaWTf2TILaCDbEEwgbVh2UaiLwS60R0cjrZhfaY/4vFq1WtV21iNjtMqNE9kxvlM0d2JE
/uu4TJ2gNiyBlWRsF1fKxdmcXmYMyvL4Av6ujT1kh3uSzRiA1zaxFNsVnHGMNx1D26+KVGTtC9W8
XOZUBHb9ZxCIgsTC7SQ/6tFLJ9lZbuqzY87rR5WcN5LaKL8iBlRS6M9FAAgNhd8KFQNyjaITLeBw
Z+ld1CNIZBJmG80RQQty/3U3U7eZwFqB+/nL0p0jfSyk+WrMOhgw1+YkgrQ0SsCJpofuTI624dD0
abj6XVZbrXOXZAHgERJxGzZRUM9GTuyNuNXrZT03wmkjC2nZmOdN+kV0eT1O3btlNyFuDIMvJNvy
LeCHPx7hiqcL8ry3U/e22Lc7You8h5tkFzhBogEtTTRH41sThrPUPkDvh3d/yIdW3cBQDxF2sKF0
+YVMp42W4wRMODoajBfIsNpTwjeLboKMDxDwIXYqlZisDncEUc2Pu/ocor7Z+N1WZ384NboqE5Rb
bNMXvLxNRf4N6zJbXuTJExsiI5ee0PZqJsLeF2IHoFDZ6KzZXW5vdDn2GjOuEyhtYQjOg37CzBzl
ly+DQ2riZ0VrcwTrp6MmHeXaDcWCJLnpwirNHbfohXpbmAH3PpR+90JqQCX6XRBC0jezE6+nll/W
RESVg4kB2HLa2o90qlHXRXR+kWc0bY2M8kYvelEiX0KSRj4SPxlEj6vnC87a+fk3lpcgVIB9Up12
xnLb/HLn/qSBfkIk1AiD8UN8peqmdw7wgrLGxKt4HwiSYC2BWqRWZoZ7Oj3KFMK+1AHXZC0BXCHH
pADRS8sN6BGBmVsdWpaVkF9A58nLu/xZO3WX0ABnonMH6OhQDBMD+GrEH57/V0pH014KccxnqOw9
6YFBdP+rH4h4kIRuhVs3f39O/ODot+rwgL28U8ug7d4i0E9Fkpxjj+KMu+JZGBrnfO+4+mUG3CIj
tBt99LU4bBB2DPSQaq5Nu9lcJItOxKjbfCXX+jZwI1ydAA0R4VDvgWWNq7FX/y+dsLDr6nm9Nooq
YqMQTrVHCrQIDV9+28Mo2i/h8gwX/MB2TgL8HzWO4j6rDDS/ToiLZkOqA3Qxn1LT27/LRGTlzzIq
hCUc34RBeNtHkAdAmIVA4fmcoEPqnUkXtRHTlAWXo5GsjRF3yQ2eRj6zTozQlMX1CmXArX+1ma/X
NN18vQi4bHiVF/j70e/IsdP8auYBLywaCV1jWmSmzV/WzNQyNUPwEbDiX6GtilU5XPhZkApCcnYl
26QfZTEab01Q1N92w+VSWwRX4pHRhyh0QXY4ZP0HbSiPqFlPTeN1Jfrdz5V7PPblgqdBK+dr+9Hc
3Hi0lIRq1JvhCo4WC9v2BG6Z1y6dxMSH2zW9mblsd1kNvMFQy7OVdVWhy/NSb/Y2ojbPo0hGGNdl
kj9lkJBglIqFYoH/Pr+G9TXCpnKccV2Lq15KohYGsctBewW1QCe0XLGJzZu0/FMe3aIlNkBOu2k3
SPUBSbMYaRnRuYoGanpgppF58LsbLb0zC8Im0+3pHuzwPjWg/ALZuWzHO497T5sChcI+Kzl9DMB/
jIg6wfAyJ35L7ZFvhQV1qJxG8/ApAWzWkzE7uuwtcGUkAaG4mo4n8pvBSTrtWxxLNAFDax804Jjg
V31pGO3U4/YC5GRhbAyjwpMeKMgud9tt+rkF+avDlFRXPvjKsl/0yWB5mgeWzJFtjJCOglGRZdAT
IalBYhhIO5uBOlnIt5rSz/VMuRnKFHnyr9OGD8rX/NSUyfXgZBZ84CODq50V6wUhblCoDoVb/nQS
ibv18sFlB3S2aPG+0jBdgBmGfnfHp4jhyHzkKGQED7n8U/7jDJmQCcxm2XhGuagC5yDy+PNj9aIA
+69CkAPtAadYSQwEvz9n5Omr6B8d9Wq+PazpRYQ9Vpf+v7ucO8yDwgG71TW6nxSovAit7Wque88O
7rtq046PiDZ6+psHkKaxMcUlOQjzxC2mRVhG0tyhiRYIuiN+Ic/BZePURwYWJr4/13YDtvtF0uhy
7kPiEU3vOqmm4wj7keiIP0jx4rVnj6GlD7ThVx7/7lvAcC8GXnr4dH5wTlNiNKIHHzm8H6H+sQDp
G3+8wjvW4Lm7ukGnS49bJaoD3OkWZdMt3c/S+YLI53jNUAMX44QUfJrpf9p8RYhkiVI5/KAb18qP
KjORX22dtAjlB7Xa4eq+BdiacqwSkP6sEtnEnSVb23MmZZIWnXXoy2+ZVavLp893my1a/VlkraIv
ItHfe/+YmMYOXZsWoE/Fm+9cwgPwDbJ8Cwv4vSGErTcRL0S3PpTGKP4zrekbOpO5zDlJ2dyRvPb8
wp+zKTPi7MZojsHfDskdgcQcS9/h1zPqdGL2D4r0Dxe4hcxWfoiOVESr4xYDmKWj4XAOidO/RxhZ
m++76/6vySUb6c12uEYjI6h8nuQt/0yq2cUBzrRYbqChy2oVSuenwf3lM4LS1uQWs2iBqSSezuB5
q1dbpNnR9+gch9GFaccT/3Y1tZdkTS9IjDjHvtFMvvmPE5vmzY/7c+1GzlFfZNSXe6ZhoLTJXx7d
okXQEugfPRkxtPUcw3LPWdu6LqR1voEfK+lYlYRMu3LwZM5v8drV1RXxEnLv58I2MCEwYbQRLwax
kK/XwOuYJw1PqLcVnt92LjdTDrAUUgGznmGfXFqmpnppezH3f64uph2WHxofDshiEWQRfHxKzWW7
iBouk8+uSPoyXfUG0drUphvTAFHRl4UfvrJrwf/lV3Z1cj2Fjzi5G5CcN8KWvoHiauAtdVSj2ukY
JGPlavd58aHUTAQl9ZocVoTtpomC+qsVTQloxESMD/mh3QA/Pet1dIpOQF7WL2hLNIe/xttMgB9t
neVUG5gb9MqNQJN5U0nm1BCvZskgTAkGvSsbOPxszL2JpFH2+GfojI9rWfM/dPlUF/poPGCz+w0B
KF6LrNniQMwDpTYjJvx8RI7mdQ7CTgV58vImniYK6pRfUNJ47avHPUIF07AF+gcplSVGB0KUwXHQ
gX3YEoPLm9nf2Nj6bo5jM8FVcmm1g8xQ2sR92bVi+tebZlnNvUKYnUMKTIvbpIigzntsSIcUQve/
9Ohl/9LYzqrUW4BRWwXSN3Kq9WNZR1yxVntuUzxOY7oxAViHslCoTxSiaCE2v5FGXxBulRIWgoZ3
s+rkAK7MKyeSm/nXRJetDUphIQW2/OcL553Hk+hxkaHpLlve029s5JLmRYPXIiMWBVcW7v1S3cmQ
eb41CJXQn3vLwSDXRmZlX+Sm21kW0PI+QpQ9XJIhkw7AruTAYY8Tx0oVhpZqnmM6ijlE+WftWDok
sC127E7eNaG2zXo9gLcKDjMouKX9EFiXjoMl0pkJR1D7b56gk7+fIDiFyCFLiK5wNtg2RJMgCqBx
mcTb2dGm5kSuq8eEVRtnC7vEI74h4e/FT4qF7sQn5Ase6l5yQYizl8FA8pK6ZD3BoD1EhYPX4GLk
MB1/P4YaaZcFsBCnO4qad9Z8sSIKW+0OzZeuK7HsBk8wR8wyetjCp0Ri6SdbsPbZOdl1FdzKWnQq
SPR1+tsKLA9cDagCwAGWvD1Pm8yvPgyNcj1oOwXLtvrmIPtgUBllmoFhezKeY0PhdhilE4xFguE4
0hMct0IOqY/m0rvcffW8P7nLd9RwTS0zzYDxc+dNjlqbRGx9hAcNWCFE1ymfgG6zYzB6FBEhq4XU
S/bgwD365zLCdvq3TiPIRiY9g2zve90/wDmkiIfAfRu9X3YgVShCG0UsM2h+jcp3SS76pgzlMCxv
4APXFaQA88dXwbGGu1hR/7ztLplzgDQQVCJXvW0n0SOfu5miP+fRR3Qmw76Ttk4gL3QAkLW0Wh7x
pFHV7e4b1AZtJ4ImdMHFoMgavHgD+1cKCHsZeSruMtXaQVYEcMQBvg+vs+duo5RvuFerZTlaX6HY
AeoPhJkXPeFNbKxXvb6849Tye/Sn86OjGZ1a1VNATAUXyaKsmbTdTiOZJbZ/jceOuiJY6Ke6qiB7
unVc88DimAaltqB8FTX6gA1nyYKrh73lrvEVpN3656jPQxMdN0dXjtDaxE8ngjWDNm5c2zCMsMRG
7+65BG/xKUcKv07CYvN908oTTnLvWzi83LBtVqsTuEbSP5FcipQG0pUWHfARKP1T0yCumQSQptgg
u08LG2NecWVL1Ruoh+VKkrmWS/9tD43zdaHYE7VWcjx3HMhzg9k69THjyQeV7grMqxLV57ZOtLCe
bDZ0N70i50UAobmvmKPBHgQdMmUemajMPw36F1SNehI2Cp75zDX1N6msnNaMvyB3QyHf3jN/c92Q
7MfV1wVf5yViOXb2/fhVeiA6kogXX0Tub4hRG7SUYJdc3fDmIgh3rXA3hLeXSMKymYPk9oqw9j6g
7N3YZaL1H7Fmuw/kqQ6CSSVw53ZfXhLu1De4HTGaGiz9i27kxg8RYshgeNhgqBsRqm3h6jSQW9n+
/nLgGQxyddEs3bEem7F8iYaZ4FemHPaadPW7AjmBfGSdxcDABuAnUUeIUkauYnOMEk6KUIdYx2x9
+DsVJKaRJdTEQX3KtGYYrLmdTk6AuD8iALSr2PsUC7mA4+QzpK5ulTiEVMDYeAoYE/ZJBg1hYyM2
tvu2Nesobc3hj3khbd4L4OW5BNeiy2+NDwAzO5aEAfM6CsMyyD2bPvSzanAg6V8cMKSjxYgAEtkw
8LRLn2tEdldIA9DBa0rGoCRF9EtwpBsMFUtJeYO3GFw66fKH0j7KrYMgDv/weICWxpSKL3UCf4U+
elx2g0W4s/JEIo4yLgKkeYo9kEGbyhOPDxDy71pyrS2P+wEE1P/IzeTc8QK3S4x+aUePZ/t9cytc
a+5q5LTE0MrzDcVoVJ3HBu7cO/Be8/MKvnC7ApDFeKt0YRwABr/jA/UucQ4N8EBC6pWqWqfj+Tuh
CufdEz7OiGQIByAgH2u5eETwFIZdeeFW3NnvXUeNCAzJ719YzuKJ8ePItbHpEHY7wDow0+p+HNfW
rBJYOl2TuRDLii/CQf7kCtmkgUj06hrKJbCcvgZM42GtKLSUy6GrX6DfoAlUszcQHSQlNGUPdA2M
+avXyft5c8EjcVtITrVElJmvE3ArrDzWSl1idx8Z4tyf30GX/Mv+pEO2SUcb2w/WWUtKWf0+sJ04
PRiYqW4wa3H+C4HR0fIQD7EcBOCTXzWEhQXykH6Bs+fR0y/S20U3/pmrOWNw6sDdJxRQ2KJakKNP
3i5/ajokJR3R58Tsk9hphU1fZ2xOpKvGs2XZ2V80XBOgM0MSST2M2mQs3qkLEVW0rmNmMtfZ3yxr
ZDMTjCV4DgRcZggbT1Skp3uXC7JlaUgV3Xx6K3OitmkuWF9omcXfV9Px7f75EseFfd2uosoq5A/v
NounPaJK9NnstUu4UtyhTxlCkMGIArvW67+aUp0dwM5RHvnWxJK2zu0xcMiqQA4qlEpAKWuK5jrE
adruN3WIFxB7RegkyQxhx6MZIXNGcgmtle1boSKZb3K/2jMVeGZC8IpraTy1azYZMDvca9ta9VgK
RMoBjr0/fWTfwV4G1uFy7FsUeEqrhnykKDBBD0A7ib5RpaomgIU4zNyFemJccXuyacGB+bBrGDzV
vOKmszHRtPpSLtqaDmaa4D2PAEJQUvL9GJOX6Z++MSKpq/cGVtN0nE3twdkFLHNhjQ0rnSjKnkEU
moI/Sw9USLVFv2ou8HCQ54FquSKsHgyUGefomh7GomZ4a69KtH0ZOG5sB/6aqLhphdzSfnhV/x0X
zm+ZyhGE4K99cWq3sQs7JD94iVLLU8zsxzLe8AKIsMWZhRrFyEFNgjGt65B/ks1EuG2K/LGzxK64
ONmsM5LLGzagV5fB+l4oCBzLbmfn5JIKIm2HRr396kFrromO07Q3wambwxwL8qOSYhzhRE+0ZzSF
BrQpgbCzrD5Ac50Ds8cZG3fXRSMSMJH9AOiyEHHlciO0yqb20FYimtLuc1QdyIC08qOvWDmCCS5r
mT84VsfrQ7qNY7LaRRE3JM8zL0c+0JP6cwzjuaM3Fo8/VSNqn2oNADtJK5HvYnMDymnK8OQ2N9VK
ALuTTNOIe2rqzKdnR+zuHA0h1IsIhKsh7UDqtgLB9VBE9oQGOf1sd+bt1RXLIGTQ2OhxuUR7vQ5b
qgKhvhTCW+ETUogbDJatU08MMkKPO43q2F7rH+gG4lsuFig95xt+UewehIjVsLjWASqbPLy7JvaX
wJgp7qHbAWQyEjs3jqoHS7RYhki4MEcwHt+uQ106l7h8wGVLTe5U/exxiaaKf67zbtsxHWunIKoZ
yrqA0cXb6uhJcZxhWT5El9Z8lLGPrVdSEKAE8us1T0xsjVkBaXZKlBf8tpLaEFjIy9Zv+eWp3V3Q
/2uMI+bhDenZBVoPalqHnKs5sqn2KOdooJMFUrlOQvMcVRkt0xzkAxEz/ki+ir1I7BLaUzkzT8pB
f+O63PSLihnKU+xJUk5/S5Cot5MDr9nOaCv8/mWQ5kDbXrCJRnvh5X4d7vO/wKg+os/Vhvlqh7CB
HMD2p9e229oMKG9dj6RKjjfDKai4v9/h9Lv94QyrAbLzkmDoPVVdIvmtzpEvcxYFXc+1yLXzMY4O
QfDDISTKwm4JBEDAdTG9SHFXPEW74FX593nN6e2Dr9WiF9cfTmvpcRH0azZhkW/YCaiiDY29l/He
UZKkHh/XdyiQcgBRCBZc97yQNt5asJLtg9jZugQI/puNb1atoUc34YbjEVHbIEDsOnuwPHdxVRTV
uTb+rd/Ywh2W8lsnY4yCopaXZd8EliUo8gVYfe3NbUaxet2MLrVh7Hsn/FpBGBEEnZzwxPk3cCW5
2W7JzPkMhoUQvCBRHfAxnBp8Ybt2rxF3wMMLiaRgkWf4N4y8SLTBefRVFFAmBemLFC7NzRv9PQyH
d0QdF/qMdb9HrNeAUM4FntufHSi/hB9sfCvH3fDBi8PUFnKmOGxY1Z9YZ2v4CpkTQo7Zc11TfvKF
q17nWfkZDIQHyuL7UqwyHuhrxTD2tE9iHMVnwz0qVeV667huzZyYQaf6dog79qm2N92KMaPblZ12
bEwBgmPjWMXBg8UxqXJiuCRBO1f3n7RFfgSSlWgHVupk+2DS66SI1qaxUsxywpW9vr+x14xLtnuZ
zFc1gQFLMB49VkeRnIo7SwhrBm75Gg8kYc+IzfidzI3wukvtSnnzNcHIz7N+8z+a0w9EtjaVsoH1
tsP6bRZQJeO2K6nCYmG4frK3jj6D60RFKIJl8pyv0QclAjD17gH23WYVuawpOJwtvdIiYXaNOmTR
4HFTjZpCO6ZHTZijuQR1Am+CgSqeHX+h0T6HUBUUAQtqaRs7muS4Lat6reqg/AtqE+i9/JPZlj9O
D7uq6ih4QQOcrtyNdTzM8Grdo+CWBdM3FJxypcDh3IIFF3wfZYuYpWyJGAeqN/MtD1Nugq0UGJ8v
eusIzxgkv0FZMkuUlcnDR2pPOzy+gtnphWr+IbCHv14HnNGz2UAD/MWBPf9yx1wzLs49aoPPC6Ut
agGonnvCPchP8bEwl76ULRtm7FLRT1cn3/D4ujqnAmRbWd2O5U1zw15LNKSbmPgpKw6inkXKqYhH
3tKhrijVpbrzmgo6ASjlYr+TQ9dailATUCO74dXKxHaC6wfzi1uf/Xn1SfrbGFctMxZdzPhI8Tah
JyeKG3KHrT4qxUK8ozcjOXGTxNASjJEYjdS4UwYtm79YQctrj7jz7yLYm55PFrbE2ISX4xTWLGWg
sjSJVlrMkncDdP5DObiXBiimrdc/kjh15siGrbqGjLf7gmduJFEJT10Zo+PnUxoRQB4MVhdOB9Ew
alE0SF0bNF/4RlpVhjgN1cqDl/Az7C7r6+OoNNS/xyNdpVjkpNV4ZDkYwVgyhSnZcKHpsxd++JZB
8MgodiT7hwesm/GH8MejgYzEo2o157K71vQD0vPGTpTVZTDW9FqtUB6BdRYpRxb2rCszkxQoAULU
02QH3uUS29h6OwK4jm1isHNSueC9rIV3bMQPyL4t2DZCR0I1L+htosAyjaFMeMFkNWgluU6hu4Pc
KQ92PdqaTU++8pkmifPn6SBnsTgvfjcsJjway/x+n2JXo+bn2FKMqwq3Yst9sGEsBMqXB9hLptiR
x8YYU+n/ZLLjAM1RyNfocHATCiJfRNRH3WC8F55IzGokoJtdRmN0gfqnzLcrLQNrWjMK4bFrqRRD
yPyyIJXTV0WXQUJckGhUiZI1VTfytf9chY1k5JfGCqPRA8DhTcJC5cR8w23+lrScP4BeTHpOIZH0
F4+o9mszyxB9RPx/Pq9zuIZ7P6Z7vZoLcPN3Dt//pCqdZsiqq2jfarjugLmS3IUjj6FP6AX+z5G4
lESO1RksngPh44mux0cJOjnxpEv3QzZIs5N6iJL2YSA+bkx/YXmCs8O/opum8MBIpee4ibOgQR5B
DPKyqsGi2xIjAc+wYVLvK/xxCdC/ZndE5/+xmpoD4fnlMFB7byMKW2fH4Ay4BV93qxTEJUEN4oZR
qIAxsmcmIziIuStiv+FeLVsXsTop9jbHK5BOj2RVkBKcKZoWQPP0o9rRd9PareHpeP6x/fSmCLvO
YPpmGJcSS5SRUvktNj6Kge/H+1wrx9YYwRUps1guPwXKP60QCZhRkyoFOf0Y0wKp1cFYcY6WI+0g
4oR4DKAhEhNKcjDKP2+Hiij7/ZxjHAXBIEx9PT/ggTkIx3EE0yvOdrBo6lzoLBqot+aVdtUVRmf1
Wba+UmGAP7+C2RLiEpxbfnZSb/zy2c/YfPq+AC2kHQAXhzSz9FaL7AvXTZMG9lBp+j6lTbu4mNY0
9M6DGMrC9SrFwKacEmrYNmTNSrhI/N3DkA5Us2sTGVMTDiHk+Z0KmaxE+Sr5HM29D7Z7OhmSrCm2
gZ6bTR+3DQGrdsrX3D9h51mR+duT1vA+rnHCoGUMPHtdoohMHH4Adi8adg/j1jx45zDkZ/MPuKkV
qxnPY0gWGhufvlCis4Q3Bj8lI9op2VrPUwDHvIZHA1SMyx7qezK/ZnXAH44FnJPnd8dpDr/Fedb1
Eqk3sb8hV+1OooAqWDN9OHsU9bBCLINeNZphaKiHisnz31arIYvQasGFVg38sSLS3XiTNuA7wxMh
X6EWUMX3zylBX1P0/lN3JQTCv2q4lwRaPC3WYrKg2h/qt0FwtLgg40W4zQYE34a7nyibal1AKor/
2ukMFfZuM7yTgyQq3zOzuJlwkYnRtzBD3I2fgvdpWcoIfbZc7Vp4aY6fFMZLZ8pmFmT/C2uRdrWw
uuZgy9bxL/j9kAQJ8942r88pNCCt0LLylfTlcQUuykr4jzURVmQtWajp4StdxzhkTXy6C5oy57gz
vzztVjyznImgOWNIG71BW0YMVVtiCthywhbhyiM3wLWwMlMvhTb6N5TQ20Pe/Tke6nhVEnRTzlAz
Vy8fdPdISV9MCrHtD+4em70ode0el4Lqe398f9iDt6F6BxefMpXPr9pBWd35QHiIQb9LA/hUBBCb
bGgoJso1XozDQbWmL67J1LWY3kvzKlSpEt9sD6kzGHsbJMA1vJ2zpVYXseoFcnFIO+Vkyk0T7Sey
fJH1gw0if3U9n4WVqCCjs2Uh4NdWUp3OsYM+1BuRQq5zGhr9pWLx3uS05iVwu0PB6hgwLs129Urz
hBhC+hHYAb9Xl1palomAWTorjs+oXsc8KTPujrOJ0/2cdwfaKJ3cnUNi1mfPdZsQOt6c42vuKl/V
sBzQzxvoxxBhg0AaN+3qnH8OX4uTQiPmtIb5wtJijznbfDsrWL7ZVfNgkL1UMjOU5V4w6+wNH+rr
NiRgmRZyX2JFN47EWHhaapOTu6zHdtnD+Uv7LTRm9kqGZe0+YB5Hmv3x/FHAHg4ctO57DJ6WV32q
bXOcf8DQDioNeVNS5IJ3KOBAuGRFw2vsRpNOF/FoM8Iu0nuU9IvAkfQfYl9cz9VFGN9QPPmtHLMT
bvYLofxe6oGVdA75fLC7yXFKbYGslqZdk72X92z8QPSMIInr+bH4pNbpDGWO1pzySVlxNecAExN9
Nhdc8qRppvtqhnXrHsoWqD1MT1yzVxvHRaKpLQTz6HCaOQRIzkqTc41aG4IBElO3zfGrmXu/SMw8
FVc6qNxP1bFR+l/erSqt4Pbci/IJDJovzE+4guk7QJNghSmQ/282pUXAx26sJMkEasYPYaj83Cez
IZSTz2viLkR0G3hPrx1uUS4EnKQw0dJLzIT/oj14F6+zPNHHLSZPv3MeH3lHtr2vHzunyZpDOdDZ
zMKMt9GG+7fEFQrQuivpjvfF5EqnbFk0WCdf56GcI7hBpXD6KhkhKmNN8FnX5ZhAiTMd2BWYMfiA
qrku8caNcuG1fVzSTy3kwUFIvooDKbmorO5YcB3T/vcO269Ls2nJds4fgHe8Gwg+Tps1I8TB+m6N
LbsIQ/hpxnjRc63cZDU6MgRqN84SQQYUcibot02VQiwiTDLX8IuZtFOR4CSq7Fa2zkEBWOkXPJCG
6mwFU5nY9yJp3M1kbxuSfng8K1Y/cNZagAy256n0ymM89UpdqUXsyD7HVKmwpJTg965ou3z69f1G
KZaPkCNWISj4AvqBRJwz2cdSVl8ZNDLDylATAjp7ws2CJMMiXigPHn52FcOXJXW2uwanm1Mr88+0
uUi1hlItFGETewnefuqxhDF1oMn9vQ26mGU68fX2STgFs5zhRH7el8J7l646TKggGNQR3F/RzJbI
AJPNUOtoccTqgK7vqox674eu1+5plPDUqQ+jjI1V/1s1+9oddDhMALSqTf/v7yI4FrBeZvxf/uC0
T7w4xbAZXRCtzQPLqi/tEmdERq2tjIQHgj6ZVbXBpXb9xMQHnR7xXpFb9QfDx3M6slOMP8/pBpMi
JS7jC+k7s5NrcAFUAFAuptKioxKIJrcU+UTg/hX7Bb33V2VM+zBPQV1F3hwRjJ9IG6ySgHWcaHAT
PKgu12Kpx5L5Mt2I0wC4Lmu8NpCJcdGel+Hjjlt6UKt7H/wP/AknSAfgcB+K0a4Y6zW/kxqQxxyC
bNpddGhmrigPCUctNewt++bXkZ5FmRotAhsHM3FW2jZeKXc/tB8kXrfzXG79EgAJfMuPRqVZ49A0
WOx1apXNcZQbe7TD7SzvTU35CPKA9wJdxGeRO+UdLWau2fYMRb55n/wCnL8rEDJEBYLOtqCekteW
r/ytR7F/5PscxaMDR2bF+sxaH9QVn7x0oQJ9zP4hEtFk5Fqr63BEHG5jD/6FVUWY8J+zoXFcnNae
QY6APjS2M0we4DwRwlegLTi9uf8ubv2KE4u/yqHyZ5B1VHhE0YZt6ueQbRDB+KU+vqlqYFaSe9GJ
nkSvo/J+19FwoEf/Bb0sgLkrLuX7T/6p+ogADjVd5ydnctYd3AGdResTsH2DxWbzPSseiAq3ZJs2
pXl2MqXA4hlF5VQgsLQV9yzgg10RJW/iVT9Sbi57Ug6TxuXlwoOZWpkxCNyIHDU5tUW7voT8nG4w
z8sdqzY3XP4jpUPptOyxBDMEQZ7xGTEbHEED+lg9r/BN+G/KZF2RXnQgykRlLr3BuEUSf2+px8OJ
LR+M+tyaVzkW4rcMxdfBO05ZgNWiNrGSYfkze+5w+uURFO7K74B0zN/wN17pz52qQh/lxFO2hV0a
2hya4iBE1tV8cpaom4ZWDEunHSy+a7fgyX5nL7o2nwcvJk1xefIY8ogx/wyOaN7TPuoal3Qn/6Bq
+W15YON3Bvl5Sxka7GpBn4U6jKN6NUb/sWwQKVgJ9TQFV2/P5bB/3U+f9V47aJAJP4ivYgyx/0mg
Uv2s26fvf10ic2Sw8s5az3ZtLhjkWchP/lbXNLDoG6ds1/xIy8ytKt/J6mlBsYNHU+lfJLdWGSUj
o+fQIv77ED58ElMz80GrgpaaRNTaSNs5wqnQEL6TkrWQE3UInQ6wQSeHf2CvF1ycg6wppTx0f5uu
eV8R9/vRHj8P13pE90iu2v3EJGlJCDT8Jkdp4Vv2SJxDKagkWLLTYrKzZaoJ1l+Hc4jgFLz5Bvo/
xGIDVCNra4Yhfh/6EvFS1UGqG5F7Wz1s33+Ws7jDgVzNi+WRWnsx0AxlZTdCLYigWNf9/1/j2XXL
dGowTpspTsic1F82bUeTh8FwHiOg9UjcJpdD/p9V90HRqEcmRkCOGZM95LXnVpPxmDzauNnNgDTc
9Sjv6+JKGF3fZmN/4nvCJwgohipwnzWRW+y1JDpJr0X7Ftk0wxTgPiXwNG3oaBKtl3iCLm/pd6AL
skxIU23zh8hM16QVXPtJ3qE2KpvqIijxovv4hojd290MW+0RSbZ3ilb4Fbxw7XN25pSyzyE8Erhz
HkNWBK0UA7nROhsMUbCQjQLCu0f72Q/HVqwz1qbVmdQzWQK79XgJMsXP2IioAqixCuNg3lRDlUXi
2s4uPBZXwzDkVlu7h4qrwe3nEgErieCdB0Ctb7TY9c+6ebZplbQQqGpydBaK3iQjn86pBN7+Q8sj
7uii5bsMqHawu9KSVHF9bomcUxWn0oeaWQQYbFnylhcKeNkbGZrn7fyk2RfU72/RA+z5ynWIGJBK
99EAU8HbUd4WCzpGvr3G04Aq1Uf4KRAvGDcqNR7H4xNEIsIu2cgXOBpsxQIte8ywmgkcqDU/Nxnb
UUC1Vm5yq/PbWkcikHJkeT4IBBUHM7qMQ8dG8DIRHhX1LkEzyJHQhG0VrXkuVWKcMcXnlackmSwV
dGJ6kM3KZKdOyoScgPePHUeeqkzqOa3oLJgpQ0gbU0vrSPpyPuJPVLu84EKifS4PDFN3ol3Ihj8h
/KGc/n52LgNJWbOphhJxDrU5Hu6N+hCqsObl0eCTHLH7VtevzAOaVFT4nEL9QIp4Jg8JmSDYPrCr
EjC3zTlokkbDRnefe5KgfFF0Lot4aKszOQDDgxLXCK5LlSlGXdduyZI8urqIco8ROWMnOko4Q6ki
MREb2dTYWtYtyKKG5LUFeq0ciUKwqBflP479uh6YZHpYVfSztTT9ogdRUF6DUTcITQziB4anZ4YI
ATxANfn9l4SFvNu2yt5pA3dmnOmw5bJ/oDmCX9ae1yjXGBbW9UlGjpAvMj2JnmtZeBqMb8g+nj/0
O/Q+mGOajXnITm4naVLYtgPPqV5ovqZL4pYaLYla6OTstUuBoLZJEaE8qEzazljvSYQtqP0Dj3fW
81OvGLPNzMmAear+6pYP38wq8gbmRgfQPx6k9iT6EbZWLjBlufmfp2JGjJ+mxFUYR/lXayxWzBiG
mBLlM8mMGVxSV3qjmYJ9BMoKCO7Ibh4YanxTk5vrhuTgI+rKUmzQFamkRBSSG0YHCzCmk3Ep6kTu
hPugGeS9fOxukMJkk23M5kS6ZeyH65FwHBnVmFW4lZF+4sDEsrogaYtUWJaSCeo9ecCC90hEcreI
Lf0P5dX2xN+3TvoYhAYkanPLoz6HwSJLVKwEiPyY/A3rEGh4dYMMvSJ9crWKuhwKpDVI/nphDgyw
fZWbew5rovqPKtJXtLIKdH7cOIf05poB0io59XrPvURwpDkKjY+LJ/JBW8C0FASYO+Jr/J+BItaB
l8EwAnoMGfskSUPkzfQoH8He589HXzvJxR4LN/MpEWFJJ3MXg2f2tdtFoah19/1GuoBXUoTdBBcp
cw1j283ckBKoR7t3o0T2WvKY7aPKNoQUCjZgBoTAtnYHq47Bzksuc2XxxY16Iyp3zkOJFR+ugbI9
Uyd4X6PhgP2ZqaXDXqjal4N7Y8bNz0F0or6TMQB15z1Gb2L4Xraa8k4zQMHNDsWm9pCbqP05r0KE
A4RdCNFpsYJHwSwpQ/g9M2qE9PpYpLRi9tdZUtFfN6jvwT2HbDoLbS62cdNGs9IfYY+E5YYD3g7q
V1nM5i9cJnZ6ZpGn2Eqb1Mgbz9xzJGd8y9dEWUKrO87cVIt36rD/TTxJkrGtjGH3vtslwWAvs+64
xLwHD932UIBAv53ChpYc63qNOHJNWr8pNPejeQ7PDSkYnHIdZR4gJX8mGJBrfRamQetJy8tIN2WK
f49hhIlyOSxfik8YtuNvvHeFZdLiDBlWm8Q3BW5jTSN6/OM5seA0ouNW/dzanjSlx57sPFg0rEwd
QUr2t+M3fFHvygSZHtAJYLl0cSrqnKRPhn0l8QaBHnEBDsk40B61KkWjPx0T+FcZRFkOm/Dga+iq
WLnLFpw8tFJxHsmB6Job4szSxKjfUe8ISk7FaEZuWhf912ryp+8MdVcEmjP7QkDvE/j4ciNofNqT
90px+T36sEqmiyVntbgITF0dV6fZWFgkoW5dy50m1ou9PJr1l5ZLe0tlN6Cxqpi7fcxyywnWnET6
ef/LVEIRy0SJTPw1yQfnPZjQbTxLci3PlJDGVSHH/h13RdL1jgLCL7znz+BmDrEYy4qq7cWMmslv
YKmGFrW3dAI3rsPJ2F90XT8DVYsJh/M1AWlVjd19Ck7fIkTYoYYkRnG35bHccvkcOPmKtAqybmE4
LAVA0kccyPC6OohuIYnCWDf8WIcwJFbLhW0oLsRbOwRVPKK5HdgdV/6wwbXjGGcg6bnuqXWok2KY
QhucQ+hDSPd37JN9B1KBKqdYYi7GFqSMpyl5ghOzifjlt3kp7VRl1ezPTBQnWZoC6yj+zx9Ri/7E
dwFAzsvUcjQmHiuyPB5RPPDarjVEMbggmmk4x5gVR83Pu6gdvenM77k5fx4pFv8QERUVgFSaTJWt
feRl1GA9aVUnJbK+LTzeXzEw6/8YFME0SLXySctKEThgz1pWy4Hwuj5Xq7P34OXaWiKYqiJyeoj+
OTQvK5m5xVbcI13Xfs3wR1N9YEZeCY1OFu865gyjf20NpEHRbE0TQ2MauRPvU7xzixkvsmtEZJZZ
nplzK6K1kcoSF+4rQyO46tAEQqlfaTB2iYjx1SzlneJC/XvfDfKaxtk7dvVCoYWcMEIznwA6DTKU
s1aFkydtHZHRr+uBgfYl2Cok9z+RydWOUfa0DKTw023bqd1WkTZsDlZSD9Hh0plaeer1nlSU8eZT
XJm5PKliyaS1FpP/YkHQU0mExVNV1VCZ/Sdd9+wLmF9zZyqTR0JeJzc+fd/Azfy/Wwb+ktvRCi8b
EbBm3nf7RW+fpVNIPxARjF3dL46llbui3f7LANhs6ZTaQmPlAUF4ii5fpNBg9Nm4rhCG31VZv50O
FKQeOPcD8BasMpMOgwDYNDcErxwszz0rDhZkF2xqaBJNqu6zJRJHqPN9D0OYEUEDX7EgIdrvuh+3
rzJpYE6NQ7d0m2eqSsOn9/YqXhfsZSvoi9Km2tFkhte3oOA5IjM/IVvZmRCVC6Kol9NsTAvZ3Ros
We0aqrGLr+5TaqMiEIIeDVQOx2XnxPPoTmNXb4geOhdu4P045/iM/NvRlQnQpK7cETRLhJZfOVOo
ZhNIFsx5WLuEaspPtZM1JnYq7hLOApo6RHEhiKkzzWcylFfqLVlPduosKlf37aafPDBGqCyJJ0Ug
HLuwrgPHXWrMA9SgMRUsGj8RR7vJQHuPhRH2u8KjC52Znn/hTnb7pCfLPBLkekVPObmZG1TZoGOj
qyyjGySH85BbeBocdark5Z7SiEeB0dJfkL5QTeVMhRgPOmtRzLFg2LOAeCBZ58srTITXZTR21SeL
IErP9Z86cRnYlGWvL2aj9X3lidW5zUG0nMXgL7ukONzEIaSvEhBrITJtpR8AgE1m0QNtdlDJU9Sz
WfBw+3hY4SHWr5PL//HoTd2n7cLXT7WSAmvbXFlcMVvjmEJ5aeLJfVewykMfEkigpDhW0Ge2TIGd
y4+9KMS5+2wpZ+lKYFgYS7PFAs7YcTwlQI0m+hS6G1YN3W92hH07thr8gWd+oHKVRFo9GenUuurI
0Ra90PCZHQfj8JEA7kUwtBwDcNT/SciTk1qX8xz/zmtTvlymRsxJzbEYAs8HxLVBNSTMfavNDoms
cW9a3ntOFukO/zOI1bthJUktH0SWsNTPP0JTV6jr8F+6o7Vuf0mhjIMDzq0AbV6AjorlMitWKoO0
A+lxayMc7VTEjz8cu20ygul5glUgY62C8Lbr+lzqy/m80qvKBy5/k3r8xNt4G5JctbvyYZnx6KE/
PUmB/iYQNQwjMWiOqHc2QOl9A1gMR0FT2BZcQcc179Be7BkWt4bH77iO5jcY+9wvFWcPpi6h2nu5
WNDmWvEwN3xixpu1eLwXFw4o4pSsr3GUzTBdBuNAbrgSvZ+8EloHgqqI+jZ0/ZbVZxDRR+6oSO8q
IirXdM7i9ARScUG5P8GvAJoZx/15dF0H/DkqbLvZc54j/wobi1XHxzLkz9S6KBuQvh0NM4QmoTsi
Zjk+3G2Emjk544N9SFTMaiNygMHSN44E6Qyy6Cim0TzW/ZvWB64roEYR5eReMJ/MV9j/MXPSmB5F
B1b/bHmnGWI4KVTuyWiEVrLob7ksXRzNS6C9GIclx/6JZ3yCOfT16NnknJp/z2REd4CvL7L+PKt4
Pox1eca3Po7qdGm0FpLlnV7L1BAk8w9gN/rwaCAEWL7TancgoDDE4Dxx4RCCb5dOfhe6V9SU4Lqr
AiT6nMMpMsQF3GFHrya+T1mCfYAv4VGCxc3ma5/CYWdICHcCNTREndHPV6ahOGS2bqKGKsIj+GGw
T/pPNI63DO+UyEu1SaIC6umqq9oSPZZgTJYq2YC1XwD6kPotjW7KMkom0QchuPuKdrbBeoiv0gmN
oSqF7Ghq7n3vPhaRwrmQqeyIVCRm3ZzmMqK5jwBEbOSUPpMlJRj/KrHLDb1mwTad8u4Rei+TShl0
QwAamjclNY+5vNdZixn8bdgtS2iUaZ426rCjcMa9fhm76mBxJBLResXXDttxV8JB8tUjZBPfMFPr
cK6vjLvmsZrAe+lV0uWvbbpoY5GTvhuOtt3I1DO2o9x2Q4fYBeAAL0BlCKJ+Zy3DegV1f2v4OKwM
iYO5VUisebOvNPH79CkEzuwVg5FZ6UAih61ZkCn+X582v/9Eo+KOHVJn6mFr380qcYkH64sYOggf
lATISKUvxPmDQMlwC/nJ6J2VJYQcnWSS8nCCswNPvLn97kP+Nlqw3iM+tPZjGdT7mcDVmwTI1Npi
EdcSUQHQLQKa7HqNMCFrgAD6+KnAvNng5zi5MzIizAHMEA3y+zhEyabB/7FbVHk5Ii4l3wXfHTzc
M0LY282tBr3MybvMyuOKKz5mu0FYLtDHBtb60bEZPz5SIEOdpy8arYCIYhRRBiKKUjpoBfTGYUFg
TBgvc0TrSpYhIN0iN6BkZNpV1j6MBqRJ6fAnVjVYrNB6mMLP0u53CVI8JFZzkT0GmVWgAm4IyTx4
3Bld8W7YXgT56DJLDyhq3vUP3VvAriBdTwQFDCOlcDnKQm/Wuetr/CFELWrwi9tItW8IYUcidyAc
U0Z3A5Wek8g+7zm2zWXWsoC6zEtEi3vUufjHKcARAJifFZ0z/jow6JprCkOh1gpgtk5p0DVjKDnr
jjzvMp14/Ck8/Vkp9FRZ7CV3gJ8xuLWqPz1JzCPSYNFzwj7wwVHeA+k4B4bA5XRdl/qjsCSrrL+s
0FMRDsB/OXHPeFcYYi02IbeTuNrwnnLxk+IfFHIQuDre+2nUf9vwv7zEpNtDxNQE8EQYUqhAu4TT
4QsQSrfp0D28S9iibdhRExrV/V0coqkOEbzbV85lyZ8DhREZLpJUpO2Nmtwn4wVsgDQ2f+uWB5ad
3IFtVRYJK+LD4NfZIfOF8PfJ2fR9Jq7CFpVxxKJI3d/VIpCHQBagC7BvMDYdDpBAa9J5Myq5ojQM
+OAmtfeah5bSOe9jchBKlvPujVNLwQqVS0Wyokv3pCbHfscs9soXIhOJZcIwGaLnXZt+LWcJJXl/
iF3wtYXHUI6dwR0tMBIZ+G3BYJ7i/BsYUbvstUVDcYwhW92xd9S7icR97qEPImBzIrTDAFpUHCQO
3q7NubOQTXc0Tzc9uf/9tGRt5FFc3EbEkVcHrbCIT3fKVeQph1XuN/wAaYLpdYa+6jBTuXGjqxTU
OVlW8r4nHZ2Kw6pM4NTH/fVBg05rmsRGqVrzvXd34oeQ/wiWhRzYCSa1QhNKv+pStt7uorE9B6R1
5l8jThFNO3jmo3E8Yw69X0uded9xbGR2IH2e6o+kUhzTX0q7UWzwT2YxEaBdEJ1Y87F65WqHyq5L
KWiHPkrGBwKxR3s5QKqizO4HN1eE+pgELgKHp2TYVisOfX6HSkrN126uNwPy4LY42krltZLFGvbK
vjTzPVo+ZJxq7WQzgr0CkeLwoIfeL/inMUmGthgoq0mWxpzfZePk4kZaEuAM2N5vcyOar7ArlfX8
/JrSQkQb/PzQYLBYhP4VWiSh4dpWsyLTjFwuY8f0fvltNJ1QgQkdoZJRo/zIN05fXnELa0V7cy/d
ummtI6rQ0lPfu0qkqhlr3QaSe8Yxx2cHdHEYXg3jmSPYASo3A7t7XFMRkcH9XIgIrJ2UOyoIZWKb
tyGudAzse95GUOeM0QjUG9mmyD5iWP5wWnYk8XNmGCEhVm1KQ6bTDNKAR4hDvO9pYHxKUR2rUczc
vw1ETOpWNMDKEOyES2NDKMA2m5u+/+tVDvug88ncy9Dwobrp+ovvXUZmXB3zp+Fbl36OUoHonBOA
wpz+9AKx0L/9WbZ2r+pA4XCu8LsHsPD+2GK+3J/Vqb7+8W9Y3K0qTTvi9sOYbQQddUNAih5Cfl3V
tPHZAMNYn3eLcpuqw7cpgx492hlT3rWbW4mPZYXKd4iaHuQvTP/DoDagH7SYBDdRNMDZEJ0wjg6y
e6t1YYd+gUP3vSv5cVQ2uHM0jxP5UYiv47AGNKyg5/x2VufIp1o5UMuTrpBWgjqHKMWhQmNAODf5
RjsWW5No5QqNeaYmNAodybGOU9pzoTlWpfMYtvjXlpaIDBE37EW4RqPUfkJSy9QexQQeH8NZcX/b
G16ti3OQkypOUhNyASAKk4SYn8sWmZlIRAJuUIzFWM5FiipPC0JqWWjpQOd8R8VvQheOTOyne8UL
Q+1x8LO0KMogWLiWsZBjkE1M3YLRdkn+RN96+shhklxVPL7towGrJVKoTPFywh/Xb67cl1xFCV0T
g/nA74D9GZspnt06sW4d5oSc0mI2kNUr2BXZ+75N+JdAVxB1YPepT4setbeLd9ANHVEqCWwj2rAe
3s2yUbtA9NAyGAjq6SKwxMBJ9JUiQk1VP7q8gpWC/LBd2oYOOBKvovrBjn7jk/iFZPQO8oPU/Ftn
D+Q4ceOz1Y+gRezq5/DAtMZmB9VU1NtD075HfdBvejSitbH8hubOaEUwfFinqNuPWKE3FH5T/gZR
vaJeX/YIQxq8jyHCVMInKBqVwg9h1+7gcXejBGaWYqIsmVvcQSaEcwgiBoT4YduoRjG7qR4P6cd5
d47CK8yA4K6FdIzAhBZOTQFcDCt8yd3GotvtlUZJRaSwo/sinYVEG0vAiSt2OdtaN5kxi4QOIXzs
IX6jcAYmcbVQ+Z/WuWT1BK0PZKNHXp28NFXLD3rUXeQfQDtNnGp+kPxwjQdaeXH7VrZEAQZv0aCj
hzFOOl3MLTJpBJVSbvCRjpQ9EwgaSsZECoY5ZuNUsAyQtVhu3kdcMy5b3ULvZhXBx6uS6x1DvPkZ
caumbEit+7tZxxTN0a+AyDY75WJ2zZXU7jX13EzCHnZ/ZJEJYjibIOU8Bap0hgLq1B4qHYpQgzMI
M8Ei2J9AgO2bZ4YR6lw2ppNp3QqfZNmu537ZMhejxk/+loxZgZ4Fe+GA3tZL1h4taIWwsCwfLDpW
Y2zOgwF74eWDWtbRkJTV3YCUPgHoHb9eMhpujO/4hlYVuYrbyxgq+VplZUzvKIRDOkbxtX7ACpH4
1jO3lWsatiET80HmBTE/33exLymzVizTud+Hr3lbN0H0T5ykt/Icet8qgDEp91WaTKrDYu+Uge3I
jl2ZLo8mlWY6AUv4cq7jhQEmCKusuMkro9Ba1V6F/VSuPHE0gqFv4EsZdPBR0baawO7nMVarsvfV
BVT+F0bLJo9HKAiHfabDtwkRUDTHYIwt/WORss4jpTv9ucH2QDokk8n5M+3gaPFuVltejqzsWLwK
pzv/dSaAmURlydgFT0G/lcnkA/fJWu8/e33F9PGIGBFYtQ4pQ0AOLBul15SzIZo7C01GS/idIbiY
MvaqI5ypl5DH3qdjGQCzHj/BpCHzd/4fXDXabtGsDDczlhviDZy87C+MUm4JqXto3pJ4DnpZMMz1
6lg0d8IKE6jy+p8gFUtqPtNtdSFAD3BY6FTua46hfzit/mYin5NCFfB7lU3BbADKvh/gXTS+f1SM
l6WxzXItnOuAmv/xUh4Q6+xKHzQGOVvJEh8l4+rvJaw+1v3Su4Him1//ST/t75V3CXumquBySwAV
jgz878yGsKMy96gClvlOiItWUeVwuZR/2Uoakm5qzRi9xcwap6Xy5GTrmeUf+3aqru5OUauTSvQu
Vu9sFhJzpVc9QlclC9kooX/oNLUsiZsioSFHeOnfDJNF10eKr50a0+PTmFQCF3ExTKdF7auAkff9
1HwatLMS6WCd/6XkwrnB8L7XTunLf50UYQukhmKzuAG6aLsmYgPM6hhl2pkYCvNpubSCiOfSDY4S
rW4OnTjivuUuapRAATQt0Mg///jh9PF7LGT7/DBK7tz7ngGskxyQNCMC5UKhKxQ3OSkSSDqwypk5
vuwN+N8hIdBu72bnQkPh3ou1wSbJoED4T5/urYHClEmyNe6i/MlPf0enBoLx9sySDEVYNYun52q7
6Itzu5jQ5ouZ4ysCRjEEmLp1oEGMCoTa6xbmmCYKxp5x6shPZvIwaTWk/XjPrxeVkzQNu1VtXrGA
lditGvE5LfkFuXSXXVTndnymrP3FzIpvbBKqSCeIqg+0dT3t6SRfed3cgOXD+NSU/3sgSU2ZWSWS
16gqhV1dTvqeINw1Ws3Xg/xIxppaDzglA7QuRjZHuUWXJqD9JLUxjHw7wdhT2AkYo7VvhenJEEXI
LoV3at3G8Ovjw7BaneHazzs0G40/hQF5d5lmbQIMEEyga5/MIi8Hf9ZNlq0NwfZgCYwqPnPf/dD1
HWp/d1E2y1OS+1xfygdqSmuhnkcBJrqLBUZCo1YeBTIrJnepu4g4PPWh5LFYReM+eLMi2GDqm7Rs
Arb4tw6v1/27avHJguDFOf9fh9TrHfkYBsJPzIu4x/NRl0orQIPuOBcmN4ElQDQrrnxFmcF5yjha
ALbfbVrXoKYsB0cjJ+Y4wZ4+1+jPddtcdpAjbIkRfSdz5EyeFCIv0mC/bfPUmPA/4j7ejW/6+dI2
+sEx/TNiN/g8oY2wqDDdubB7NNf19XLGR9ctx3LOrslawIS3tM4iab8W4Wh/ZI9xQgzIw4buezEA
1uF+Hn94RCCyFOIIwnYz5T/sw50UKBN/+eFxIUIll4KXB34nDSdSLE2up8Qnz1NcapVYFUnuffit
OHEwzscxuD6feeCHebQ4MpR0saJvXnWN+hjL6+YeKiDKVB4qSKDJGajlL0Mx2/GVRa4vt9LAorY+
o+QuYx3ntXlsnVk+jNsu0cOkvTV7zS9aI6R+TPiaf92wVJpHWOT/y/clXsTnZ5nhrA+EHxko/6vw
K4vz/FO8+0LHcKvaS79G2AUSUL10WYDTQEk2X1rcWSCJHQQquLnlzkuS/m+t81hC/IKmnva+HjRi
PHoHeO1yWjtqCWLG8k4NUIadMWQKNmg9NOCnfEu2cVMB5HLF882HugGQmAqBqqQiuJUOCU60laKa
5InrZkBEHCPphkR3t6X3oagxiovdcOvsWI7J95JwOs8o9sER190O+N9vrK8tS0H5uhx9LG2f8+Lt
/DqAQ6f6/Z/Kzb7y+I7YvGMOvF0Z3BRO8m1LMxYpx+soM8eWxUq+buJKhuOJjAkIXvHi6yZTf8Uj
Lrs+C0ysMb0Dfnjvvr3zF1RH0esAkSG5NyZ96UlPcNquRKAuCmdQa9oYkyKlzCyVoBmLh2wzkFMc
kV4aW3f28VSs7VzXSeoMVdcuJIkaz9bWWXu5yeVvVBzHQg29RUg9pQlI1rE5vPltBvoWOs5VAIk1
seoqT3TTRPczxmNtaIWJPPZ04I9YuHuq1/3v4+dkKH2il3ZDV6CRz5+FA7ua8EWIziSUuKn0uIBw
Eo5ckJu+ZFW3a2NakXxbBG5feOCRbDfeaKbuIYRM+8QgDIZh0ccCSmIgtwtKt9TSRwQlsRyaPB3/
DgOo7W24J4Oy+N4y4MoAYRc5eSpgvH1OcmuE6K0oVCl9Ir1LeuvSXhj1R8rdYcdNsS47dAVrCHkN
fQPg4fxBAxxGWyBR+Kq5kcoOvZ8k12zT9L7JxQhYj6dUtRryClZAaX3sRp7Kxb9cpt/RdtL2wEUJ
R3zR1xd+7Q6+1t1qyNc+svZ3HV4/leGlg6xmZE3Z5H7UxOcWuUt7UZdV65STgGsPdT0bbJzojliA
tzEiY1QQZkiUzIH26icNwFlC69PCDEVQrTbExR8PBbBnH7aGLowHbkYHCVPVhrusaBNVq3xfm+rn
Rjx1SRNgQcz/WrDKhenGclnIkPreH6aEaBR7zIUQKCqLaWyu6wWCnmVmiqjoq77J22lUL/WETYdy
L93JfCNlmQU5QeCQtH4sLKenurGxFMiRJARtbEHnX3gxa2w0VT5iDSJQSltCnUcEQAxEOf8KoilZ
Cb1b+WIHpZ45MHJacmXjtx2TUuWpuRxj/aPwfXfytgLykJZ8qO+OygCwQLS1EKm9oncWsUo16Q5x
Gs1qtDxG+TtZYIYqenzKEZ7RqxAah2lRdZMr/p9hYyv4Ymq4TZF3EkNlBMmNLA3q/WuoXFKHBmhA
R/S9L3Itz2rbjzbBtwVN10lTpwBeKvT2RK0h25tcvzpJpg4s5xUQYWeqq3jV0Ys99iHzlPsaBgu5
eCANn/CNXmbxsIbz2bAvLVBzgPQO8WCt6tNElQxs50epv4Z+yxEQ/NgZNrLtZtmOamSuPDBIB/vD
NuJWKNSnOfIDv6Vsdhqe1L8NSL4Lk1SkVuwfAjbLjpq44l3BGpfKSwDoE4/ZXPbdTw6+ajeZ2AFE
tpLF+a6xxOeuOzz71N09GHHKlKFdkPM0RXWPorvB9UARLH57Ko5ORIGCzsqyQrpMuDU/6zGuu+1U
GOGB76G8hPCAty1Chq93DwcWXxRe1CClZ3rQLbITv+UvorJ7rh6nzQzutDlSLAdH4H6QVODMPGoo
1H547FIYDOB4xlJNOiTnnmtEHiJ8Nqr0rE68AdaMTLiA7iOM3ifD9MGEaWGozaSnk8Uu4loGgPYk
xUfZMH1bChKUmcaBg3aCIePyBb36jLJivdkUWFzYGucIO/kirb1+sy0fdE/Sf1EwyfhlKHNQibo/
fSKWopmMXTkH9Sr0fvwUOf7H+v4fPJQ81xjy3XLIYbvkmf/C1Ab8kL8bHOyj5rIfwtptS+pGwM72
YswKQDxDMY31mkHu5DFTfiN2eUeLBaItrSlMXwgWVn6c8lMATQeguWB+CydPvLsRSEyMXjT1kd+2
GdmkLRQUa0Ajt9X6r1f8hoE0FCN6EgK0mqcb//lHfSTpBi9VQkmm3uy+MVQLkjJuxkFh9MJGM/br
gIN+7kSoop0oN/sPVPYE1KRbAPHsfQOhB/3+vgrcHbtBb1/+yKKmvOv8szwOfuB+QkIsEO+wUQy7
7V13GrMI74FqiKP/XfXBAXlZmjtLEj5LP459kpmykYJ2U2/sNM9748lRWcHOBkCweGSG7CXYUkbQ
VxGUUIvSKhtZm8SFwrSafFcEZpMZWs78/MbG6UKpEOu8MXB9BUUyPXWtRsBzxgdj8gb8BVOzeoKy
KtXlxffsybwpMaNmbrMfBrf2onpm/RxPorstDmjv8c+m7dy7ApCweESGQEP6MEPrWKvNCFsHdXQF
F12PguY69MKn2E5qwVDtD3Rq6kTxLJMr/RmIG450y0NmD0te6lPD3uquA821aD70rtqwxdxYOdjC
cHZA91ARleldiKd+07xBNE+6n5ubB0bpd+eRce2F0ZS7ZhlPJFnsHRVWv9zMm5TxanTScZnsR+2A
9l7i3PU3p1o98OozgASc+hhSHVbAVmjY/qNcTc/gG2U82gHnwmyaAweDZ+12X5n8HPNc4LGi6R+3
3Pv71QPz/17IXOCKNz60RLSCexdi6LpyGsWymTKQ7j4336sLrdNDhmCU2GRqpD9ishdRu73siMPJ
RVaHN8cOoApgwtPWpb5TkRa4zlTpjt59QUSkTGl6uU4f76KSt0cCPmFYVB0ZUglOCklPPwwqZVq8
mkOKkjYVmBw8/DeTaB+8bRFqpgZwCT5bDNmZJwiNoe3MYHrEteHJO3oQat+PVyWWAWpgIqs3nX+j
dwR/zl/SS0Kfb6O3PXeZO3CihpS2Q+0Mx785CEsruf2eSmuEMfxVNvMufVn+7DrLsh249fvGFXq9
71nBxMBWpAVhhfWPZDBbdErmtLAjlmTqh9bqPnAZBJtjZNMG3N0Twu3U0ZuJYBQuu0cA89+rVkrO
yNVirgcG45pVNBd/udZVtmp+/RogZhISub2ybdd6DFcCG3ntXR3YQ0tmIHy3dy3ajZT1fJrFTVrI
82/0fLh2oE5g3RuRFq5qeXtgupP8v3K9uliaiEy3M2s8NHcnY37cfmwsmz4GBVnG0ubpSeOWf405
+o/dr9ueeVYeorec6X8daaGg2svwUthDMWkjP5STs8+nDYGd7D/WpFLM0frNOMNaMnPdn5HVTutu
9xumB0LVA8w1cUFyrn0PYcOF4K+dZr3rxECrJQGi6trQXC3BOtJZe0YiRVff2zZZYMprTUpY39si
dO8iEsXoHCCMdQmKuAgJQqWLq+FkJXQw7tiYYVPVt800EkPYnbp61cDu6FCIJhCvys970vEs4Bk8
FsG3A6ZsW7TdjQCidI+igMWskCEfIdO3A5LXThym7BwTm7nRYyTQV0mAIzfKjsSgRB20cjuYyDai
yAhMlbakHGduOF9Ia+DHBBQ4duKXlN6q2pVDAOo0Exg/HwQ0DFptGPTm1DwBRgTbjSpYe5T/U0Uj
jp6XaKKgLVdnxVNV6MbZtNv81IDceVmuRdw1xqapl8O20euECOZAlmyA6HIU0qxOZuja0tYzRbMD
CQyYGRtmX2VSbMX0R5QBjtBEPcXYq6ZqGeTCdPcQMSoSY0yo4VjD12vWfAFvr0o0r2k0typVykE8
SpggiM9n5y2YRWLU+SThi9sMndkfNQPT4cRwdqxRmV0W33J6JpCDpeyO38lgYY8+0ZtHxI7hafYN
PReD8d/4O+JMvsq8OjOa8j0lv1lsm1s+nJafnWG56BHSljhi3FH4xzy+bsrvVN2Wye/GJk1CIgff
55IBS3hIeUFF7B4MaK24wGBvS0J1FgBjL/NivXkLFvde9RYX3mouVkqOBzp4Rxpzoby7QgitdnLr
UxgadoWRkL3NLywM1/EXsH2smI/5+kFiqPUDBoTNMJnWjNBvgeGjLpHuAFaKqPtycAQl4hAycr8k
iIqe2DJZ5+tkNosTCN5M/6t4gAoQHJfSAjQXV8uK6EN+um6GhtFCQdb2XGAIwMnoBFrubYXxh367
hNt9KCCUKS6AGTnlOB7EFF2ZD16jdE6jgeCdhUsU2/cGYQIddiWIijijArRZtBx9qlB1NrfH5Mx2
prnEH8OHWLwPh7NR0yDt04TmbHil8CQfbz8YPlgrHxZdwc2F7RZpegajY/sqjOsPNN9+AWgEKsvT
FeU/Wf9E1I2EpTKRkfdk9dgUmO2QDOd8JQ2vSHsJiMwqBDLBuqBJYarglPIVr/zJQarR2BkoAz7u
KVw0lXyzC+9Yo5WMAcjlYG8JhThXKW4P0u54KTvqXyxV9ccxZUYiTlQJiYYyedwNkIcnfDspHMSr
Ne95geRgt+s/40qMMrCSGuHPjYtnq60IOKYWIDx+8Jqb0kwHlP5iFIN63OQbHdqr4cjiF/+AJ198
7A7m4ugMwBQGEWiqQLvQeeiaMQWNtCuUHUE7uSRkE9Yrlbw9MoSl443HuC/8AH/2/6D6vn02HgD5
wQw7CaBcaO81pw+c39T3qU039/knsVidW36CNvQW99vE5hXzVbThiK9Rq8sltChmvjREX0jgn69j
UhZaa7S/2gXUipIf+MGaTTqN6/NNUPwpPvjA62XuvHTLAsaim3ikqGB4z1pFd1Fp47EkCrjqdKLh
ITN/IEBC/2P3KBm18AQUz960aMW6LG4Ep/kMYXLqG0xYd4+Puk7/u4Gu/qUV+MB/0DTOFdtggG38
n5EYLQDPFYwNKmHphU7/Np5Yu8hJxDDvnVFRLGFFkS5uESRgKuS661HhoWavx/s1epJtNqf487ae
KGXQB4qTaWzrY3TbtB80cluWVIHxhy3EpIkAtbFI89nMOXz+0WHVDeaoWdyLCmLPZ3TNWcZJq+nY
rsk3r1K61LLVWuVdWUtyEg51YMpO7dVjl42TKXFN4MmQpAPPlkM1ypz1Z2sf3cWmp98sU0JJzWjU
KKS71BNQ8ofUI301gvp7wfWGwkHqGyc+b+M9TA7Ez90ct2HBrv0MS7TKolxjaQJkCXbHnLYF+Wxm
Qi2PnyYqTtzwu1Qiuj1QYpm6lOed+bh1pUVypO+NBAdzABHetVB+LjESvc3wrbWpTPtXjYkBFZAi
CkvgOPLtkPRjoXcRbt0QUlUFNxwA0rvy3fyr1OIAnvKtwvywCCyh/9JhJGIqFneZs92yP0OYqwPz
EI1ijYkCyxtijJnMSHL7cjFqQ4uL+evxojlX6fKeWS+W1+qryxvbKukzl2SBSFQuuK9xISLnFnQ/
Lm0Tmt8h97FlgaLnGRxUfnA9MMpMsSJAHQ7zBRzjh6bpaYF3UTdL7HMPc0u9Z0UQgfgTkc6ucCKF
ywbbPdqNQGKDcSoLECFT0QrJ6jnbXo7Sd0uAC4vVWv4s7NBPj4eTakKXffewzYMZ/1XrJzsjqmK0
YQUqd6mIeIyywBs732CRFZupNgiOZx81t/3wq1l2O5Qi23tJTgtspiG0b1uHGGSVQHL/W7d/UdJk
Thb1c310VwnPzAbZbpfgjL1lcWYbsZRYyxvZ0ti6GzaNtcrkijBsgacTbLP9KxapVvQ8mm5Nhps3
LybWNyh0VHqM+nzmdEx4dR/XQtUeW2zZYyeQbQxAenML8r+DR3MzBvuJrl2yWxOqYGh8I3iTICiU
89ovNd7So9fXKSaayKDAZ2ZjdR6ztFzEshRdBC3ptOA/u47cPHXz0rCwsDzDBZ9ar8qTJ/Dzv1FE
MrggHaKZLaGW2OEtvhqlSgYnHNp6cukf57TxRffjSsq8sTZl6jRtvnIFZ8KP9p1WvBUhG3soYTS5
q+Yus8uVKCMw2QN8E75TvYsgL+OZeRdDtf0ILmlAs0iJkZh8o2Buw9SwYIo7A8sa49Q5gQ2WIVtU
5lCNLz+vJFBfLNGnjfD/TB6gUu8dkb9IG2BKQqAqojL7VxSmls/+f1sMjCCFxKCRuMutDSEs1VEd
Uv65hX7dGyH+O5OnI0R61acIvRBem1x9DIp6cuZoipaQbZ7Eh7rbIu6CDKoQsDpYcNzXg0m9OgEU
Jhv1kb9P/Mdbo1O32nGGS3Nobew6mP7QNO20Vbu/LBT0Sbv0QbUzIRszf1/PB3wwiffRUq4TkixB
f7nin8jQScdHtReH9E4IpP3b4+cp5AIGO+mmZC2Ic8pvYlL8BMHVLB25+hhRJBj/OdL/HFQICRrC
tU0Q+GndbrWRprDXR02isaUeT8bkEOZd7qCnduMNK60stJ6rlTjP5ptXQmRZT61P0nIPPfiV4r1i
Np7j2lKF35SCGrP11Msz+zO7GPHS4IMvpRIpf6fcPVUHfCsmKSDVqThVdT7Y/2AL5ObUn1frK32z
mvsYISDW0BB+RpB+D8r1UjmHlMu+lT7H7/SA2x32J5uMUbvqYFeEl20xKJ0CND239NFOwz9uEcdf
57bJrThpP/MBLIa5JFZmWTtNhkLLsODnSDkKTbVduqd1RmN3HPUsSfBoDTxPsPxz4r1pJGgfxvPx
JcFIqHip7n8fUYR/W8OKTRGawEHr2qr4mXWpqEsm3AN1oXlKq1FswyAVT0bllOI5seP0z8OukVlf
e0R0S7mnepQwNRfMQFnlUku32XY8+OdQAzSldIq1hG2SjxiIgUadEz9uX7Rg/U0nioMpscN5MtJ6
foA9E3hhdBeUVtmev/rXoERwllhEhn7wxhzfUzFZn/lF2OztiZ3hWFR4Ak1TuD0XnnP5BXIa381D
BXrv3NqU6hAuGVgQ07OCJgjJbMR9jPJlR144BJagFCWFnRANUAmnZPi7JSSxpUuidF87HJulpdXm
z0D+029feQvY//HnnNk2HpIOeWfpXTlaUTUyvUk6sFjMZ9DUpSOxvffitG2LPJtckjz9qI3Bw5Bf
SBJGMcsNMxmPamDj4GLT6nzluGPY5u/cFaM/aanJj+LnylRLPlT8dBFBao2dh/IgxkK6hRakupJ5
SoyNMWLYUHGpbPWH89PdSpFH48LhCqwrAwoi9tvbl7Kaz1FyLnWz2VyZ2/mju7HRDRxLU5/qi8PT
FMYNmZUg9MHdaYYYvVq4ZoNYSd063TNYuwAIyRuA2CoP0qxy2Gyna62/4rsn0HT+XwBq+bqwueTi
COY8RPr4RqsxVDEuCwbm267mzauMaQ2d7M144Wf1NjO0YsaOPiQRXmCK3q/7XcBIrTHur4HutOTm
UMdyC9FVQJOzQXQlmr+fh6muA1VP0TGnZZhGeBW4KLq888JdYJLVg3zjJYCQRH0SwlREB4Eem0t0
YycSRSibxf9ayR3W74Ac2izRoUmlL44htFa/PSbNYx89/j7VJvNFg9qbkCR4DGrtOMmXC2CZOhxM
EXzeoPHNVOvfLOmKP0tN6V2HnFXpaBoq45B2b9RkTKsNud71dAey954CUoC8K5ITP1afoWYZZ5aU
zbaZdcm6vrle3TT1uAoKRJMn1cI6NaDxw/FvpTJ0ZoFxeS2NIpTFaXNNnd7eEx0tmsOrKbV1PjC2
d5i5E796dElTMFLngpbJsOPn/S7rSet829ssTj/JBBx7ZUAjDKFG7+Y3aevh6/rohUGNfxgaL4P1
U0px9VuVU/p74W9QOLk3uptVR+eK2igEYe8n4laby73OePESCJt5oRhMG38eepEY/ZuXuS+0sDWs
eCGktY6Teh5R660J3WKxRw8UwLPOmQtPC/O+6EcQnqNxgcFNKpFfe5Hjz/OMqJ7YkmKC762fVfPG
UrV64VVrUWLQT2lTOLSwpUk6qIB7wsOoIy/sUmFZVkoZTUFw3akclPb8gzzG+URD8uIU8KJwBZgi
oJQWGz172u1ziK2dh2l2wAPTd8jy9mFfJUArgcX1VoMbQtmfnRL6mHOS3BuLfJnwlMVLgh7gJ0q8
w3Id1xFrCbNq14Ytti6X1sAffGOm3UE8vkJ7JCJKMatZ4qGAn53h9eGU8Suey438yPiNFop9pLV/
+mweRgjFVec/xQftrRiqYwDB0T99dItQBxtX4AtRXRavAjpAEYZOQqEQOZ23PfAi2ToVBG+yu0Qa
8nKKZNewt1DSHO91+KdB2cxpbK54WeqRhk0BWMUnztYkjpY51cykHmuge6Le7qOE4Wnunxo/eMww
C4Q3S6VSucFipBt29O6wpgpcYI5B315dbvZRGwtW2bJEb3D58OZgZBG8mlqpSuh4Jcf9/qjxf5iA
M7lGwURSqpJdgXH/fHRw+T97nqTm7l7GELEdUg+iNgULC9fVlJZcmvPTMd2Sf8ZbHq2OlX2hF5b9
z5ym1UhWt14YGK+pBF6Q7+1a4urNcS1fYy1xy6I2I5Twhvo944Uv0zbe8ahNuHslMOenHZ6GPRTi
Z2KNthO1WfMryWqkCr9WCeSI6Miqn4HFu6lAhJwEpQ56wap9FrkAN/pnvKToWw3QKZAllnHarUg2
3Gaf9bsfttaB8zhIBF9TW8cy+cpLWrqAU4b4ip+5XJRFVk6rEFqWATBP3peWUwNJYVa7tLIIKQ+R
OCXjBiNmKC67aKsnH0FxRFwUNzuWh1RoNbSzkc2NHgQec0NSRnIEGAmnosjoNiPdIxgjbqrhLgoY
WswHEhI+IjwzVQ7yKj1l+OgW9dKJ9M/BIDNlhmbtuWHMK7uKucKRnj75xMmtJO8rkY1gOtx/qWV1
wQf6B1P13cO7XnqWcvEVANjD+W/v4njfSSy5pqs9PD/G0B6O3wF4F4tjHGph/uXaz0vtAMYriGf8
qBJ0wk7zcuopHQfRXrXo/sEizu5zMDy0O1OfMZCS+K3QLDikTJE6jacJLJHEbt2ZKyGsmOdZx/4S
oCt9+wb2xLJP/j1ye5VmHXe/sZi7E9rQiUdk3uJgAzH4ekeX5TpWKe5vaa9K42ru2+mPvtY5Asy6
yjKEpo+QV97ChUyZjBlnt8QRJO6Jp1i+f6lIP2tVCUFDMf0f82J/GASlizSs6uMTn5L297puQyQV
SjVvA2sSqow3Dv7Y4CkopYI8HfNtN/xHSY46rNtWD7547q4FdyTJfD/5L7rjS/8Ciu9dEq8kauYL
Tys/n6AF1/XpWtZg9YWeB25n2eMO880m9M9IfdoRu+h8qvPpovx3sgilGFenrDehDK8tou1wuEMX
pQMehaVFz1l+s2F/JhJY8K2iZNjXJlAiZeY24Ic4FlPWLUgGR0gTpPzRymsbVFnBTceYfgOObnT9
eXBzQ30U24ZevNu81Ua1xbDBxBedxMcgg+UypbXPWNmkXZnjsF0dfWN2BMr6cgZoxyRILxYlJTZP
meH9IwkazQV5HJIVKQEMeGv9g7C4kC7hdI8H20VYep4MOTGIK3c8yVdt63SSO3MCi+cPGKGNVDes
p063llkFwcvwn3J0aM/+AgUT4/QZK8jMly8v8lJUcKjV6Ax2UMdKI3r+vzeaeQEHM89P7gsljdp3
foiUTn78z5H+OtolDsY+NzZ9MGly+yciesjzF1zUKZ5Wn84E/gJkzpmzSeCcxY7/509Vc/Al86AM
bKAN8e8oqHfCGWDLsSoRdKOheL4TX0QY+4tdqlyUAZr8oBzCEs4x0admkCmJ6lgosa3jTNw2UNbs
Ep0qQeBDMQF1WLYZKvhdAO3bH9+dqDZQZXsDEKK/LlDBA4pk4v2+LanrGfd75gceWVSQRsHQpFqo
K5QCJuiGgVKyoSKRn8UUNvcBtdCddPVbGkbXVNwd+g7QC5nVDMeM9eEHpbfYshAHWK8tEuVWgMlZ
5AN9cR2dVacDF7Yd8oj2LzhGxgCZEmV81JLIVWXso7BqAnjThOlMXiDBUtaCv9Fpe7f6282vhB4R
u4HMG99EnPbW9XrCYAcWGAdlGEiV9WIG4R8DKZ6mK4hvtYht7HLlcTWBgkHyw/bomUwXtWIFjqhT
38nTsPjmPQqDpVTsIDLV/ZEGAq+3fuyMOVPtGf/lTcmQwmXksoandNizuM9PdcScdP37Ks3bCRTC
bI1YsN9G1UpmWsfcIxwT72jIrexOQNLf3qHEKztR8kxJxig6eJdDT4AoyplZKfbQIMV/iMzj5iA8
2jJoq3cjyNTvj80EcRZXwFVRSijk33DsJrKlq0t1THgC2EVgMpMrGW5XLcmb+/rgRqX0N3xbdiGu
WIUFQCC46BqQP1HqzulWOm0e1BFnZ+RzZM3Jxj66whdNUTtWpvYGHguZxqq2SUzXrxPn5Vz4jUCn
uLTNGOt3TFrD+/B3UArILw8AtOd3KtlgOUKkq/tZuhmdkKinqx2rVOP7eowBw/hV2ukZtrjuV/78
soul/Dj1Ha2WYFhoATXwRjOIxhScjHszHHrWeZrWhA6s267v0jla3PQLvq12MSHbu37kUbvkAtXn
DeJEOvHeM0gJI0gMKaZHdc60uoU1l8lL8JiAuskd69Ui0aHqUf/1Ji/hKPP7eydL96QgSJrLEzNm
KdBbH3ucoj7NQTxx+0IHlILK/wZK4L9pVt3cP/mwyk+3MD1Ij3gzr8nVGICD38PtpTNU2O7Z4H15
UxFRUwhU0HDPd6TR1fcq4gduLsA+kHUDOi4URNZwmYffd+Lir9f8yf7WnLJPEFHJLdMSBnp4hSEN
94ohWnssrnIIZiRoYh3SWBJJCCz9wD7mTnCNtuD/eT2G8KgBywyFKjnqnQvTNfz3m68LiEwLWpeP
qcjkcw/3UzfHl7D5n4t47U5MPlvSmzDpuAVI1HwLDFMLTOoQrBwjdk2Wk41uhjE8u16azzpDbwD4
f62t7qiWNca6X1W5y5/DX7FpDfUc6DsO7AizJeDtou5FM4qsRmnsImTN1XWSUl78JtrzkDbURp2Z
1kvpcDeuLvhLPAdPJ9XadTKrSiKoigYObAjCrSmXoLbkGINrB48u14hRYzHq4IMf2baRyhqPcJfT
5alcCsQyeNgZ5vFpWpuMWRYEf9rnEbnBNB494o598yv2n5H67wd7LaVgOpMhF7B18BPES9MWXs1h
mBkyKfGNiRDBc/4ZIBwG4BQZKaEB6KccobeSXMYdeXjfleTG9ctxhqk5ZDO99Qn+BmzOqS7w+lAt
HkeVOYkaO7Cf8FUDEb9nn122XFZvj81W4jvObwUZ+VjUfhVK+r/pyFcPs1SGg58IMx2+9eBeQnEh
FtPUIb05GOo6+uYMuMdCoYL3kGWXck/f2CxNn8tUHrzOfGGpx3fJe5XXZcYPJQjxQioKugbsz+H5
f3MB4ji6YIkpcYYJlGORfWz0utla3OfGppGDoHWshLAdcT7EYjJuHjrJJcADaxW8nVuu/1t1f2oW
sy6QrwIrLSCwNAizyDLU5WzmEC4x7y+HROBJmpnX0cJ9BR1OSBIWEbpDj8cnWqiEUHKl7J7mHcUb
l/EsTdnI2u/f0StH+9mUgGcS5y+krNYgK+DTxvrmdWUXAdo9wPA4Nq2F/aeHgut65mjfoOhiJNuU
dDEJhv1s40kiWpQRT8+sa9JDJXIqGOjh405OWcNNq22Yt2AdSoOCVIX42OpCcbBbpTZqnqa40+rJ
u6WhR+EnVUvoO118+rkFii1V/FcJfPz4TZ/PZtG5wOj9ZTojZaQ+phENK26M0JLrHPANOSczubPs
zt8/4gTtCvjkRvZwLUTMvoYHFjOa6C4SbdePlzu05rmOIibJ8qGSW74BuBbKotGe8dCxZexcZ8bS
GxAHhOKJ8gpY+BpDT0gSMiql0Ghw/DPmMtstfZuvkKMM4nZDdOCvjCMuzwqC0gN2P98Icn7ZWzUe
HIvIV6I6Su9HDLOJQo8ITJBqEmldER9orLMUnsA51Ao7vo820WvNX4P3UWN4j4QhjBX6U0J17p9G
0Pp2IXRQHqm5CYG/5WxEcT3BXpxjRLHhYXunhF1gsstlrB6gLYQSnE+d/rXxXcfqOXeau/lF8AB3
H6fi3hWhB3FsKDPfwCfYq+0gN2dgyX1U/RcjdXLwVdbXUf/Ewk/UwjcQLq4Lkl2eZvpCYrmilyLV
CbUKp+00cOIl0G30z/BmAQDOhaSZ2CXyAVnCioazhaSOgM+sJ+WSgU74Zs3IM9vrUFFMJ3g7HmVh
bcZnjfriuA/qycg8z9KiY21sNOvhgKnVGr/2FEjvATuAehFmKnvSphFZs2yI/SV6Xs1NaS5dLDT6
CKqEVKQETMtyJihnpGltgQaAwR35fwz9wPnKIJlxu0q1sOMlFN7NvGSWB3tL2pwCZjWJrJHTU7GA
0jt2wMgoWfHCRZ5WuR4TuGUGgqj6iiRfwWxzNy+DunTI/5kWkoeGvOXRotnDy0ZyLuvmfT14XCNf
tAp/sUIqT9SgyByyBVNelceMqTneHG6s8ZL9v6hIcpha2fS0pf34wgz7YKSRJaUbHhLmI2e0yGo6
A2BBOYy3gFplUGW4BZvEPPjeqBbYtzQd9Id1vheb8oghpiVN/3lDndTZWKvOXIM8rCYrw6y8fPsL
RdTRTWRZNFjQgyoP8rSC6aID9X+uJD0NyViLVGcbffV0NExE9t86UCsfb7KLwRZMz+JsURBUuRa3
qpw/+bO7jD4nH+58dfWj5QYsVEiE9jdZU/2U2cslfZf4MpUGVzAFR0pZ5UY5qekm0V9xRzf+XvLy
009O9rbUJ5nDeFouOKDJ+ZwmnF9pp29F55Ic5ne9eqSpTcZd+yciUVCZsjGrxaMWSC+emBYWkUvb
0sUF2llYnb0WfOdOJSh9QoiED750yInjHAnSZBT0cXHn+gs8WuqnuPf9VWz6uiRFi2GO3T4GTGLg
rQDRs/r+4aji6r1iwi3zdzqqCQPF9Fu8j4ylAMHvzaWsYtmJMjZQsXaEv5cU6Cpr8S3w5WEPg7oY
EK/w3jh9yLVV+xaEhLMCJeaiiAy7kCt7jTG6ECz8JNBKvB5hxMYEJnELVzJWgAmlMYOXi873h4+j
lMkCPBAQAGlA0JbqTzcFa+CkCGqRjfi+bvqaDFT1PW4IgRoDjboclteVz0oH/vKdHGJVyGm/kGLJ
YTcGF2zLurpdf2tGgc9IRCoCoCqQ1zt9odSyJcmppG8p/XyCTqfUdyXfKdYQRtUItKJEt/LEREI9
z+6Ui+UeQePs/JVG1d8mPJHQbX/CXRmL8nuwI0sWqpzi1rOvjSCiL5Ka5mIXlE1EXHIWxVanOGyx
9XCYDI5fHLyvM76fIDk55/T8LkApQA8bda9eeC4LwpZGJpEmvNs0VfeDC6bzA0wc3+iX2iArrzFa
1a0F5rmPp2iraCfQ33avfMFHhy0so5BrQ/lX0ZcIzgep5+ObSjSEIaDaHFCMl7H25uf1Nh8WLUDD
SAbHEwVffh5ja21loHA70V0fXW1/SwFUfd47y3YS0LjT+fTqiVFVPN80Bnv3pnRgDaJVCX+Hdi5E
qY61YiOX0EeI1XEoOnwmoulbLys3J7vMfO7/3cTpd285OBucY3e6k17v+2EWHNk86nMjo8hGAe6M
hxbb1mnC4Uoq6l0lpAD/RfWV/8bAf0j/QZc72zYAaypuilcYOIVeuFjVZ5GB7JqW/1aIAqVBYFVE
L8SummFNcGia8gCKykQojpEU4+d/zp1HOG8timSbBAnQc7y/YAWe0XdE4zRzEnRenKSyBlENXDa5
80SIsRD7RTaMYhj2PkJp8CB4wmFklMgL/wNDjHNI8JVepg1sHcaLC/HG+ejf2IK0c4BFBau0XMpB
k21si9erlZJRcVnE420yqTbbu5A/ryLocBJnB97pShfnF+VMMb3U5ouxa5Av9MmTbZTwHzTreuan
c4v5hQQSABBQAyhKcRE0OMnEsQxHiS995xDpilJLGTOMYajYv1ADgDi50sUDkxi6JZOYdvw1rUGh
YAQqBhdOaKWv/pyF/j4MfPY7r0q8qlkJlm/a+dzdlDd50IGt0ay+1bRVzKLLb1mFmQ/57xa/Nh/6
yiLdzst4dDunbOqjRxza50Jc+iZTuVF6A0pvv8X3ZVEY+y8z7jDHAyTlTkit0Ygr/69JzNycbwlZ
D2OwIwvfYapZSps6r2L8h40nBHr6W+gXsmCFqyB3ZqfoHMUJk0W96BcIOIyvSbxBo9zQkO3DjPo0
Sc0AoB0+WxZXFx0yua7nMvUAu1lNpOUbW5FZeaUXaSLKsV2EdPX6VP1jDLnHHcYBLS9Sjf+N6OB9
DF5Z7BtEyF8kVkapfGte5aLNPU/heTg38OvM604EG6Bmx17u3fmB60UJeHix/t9u3v2gRPfg5lsn
ch0smBo6Lxb328Vcs3tfEfwdOqMfLjOu8XuPr6JxGE1e6KCoFi+URcZaOI+mNxhb7M2VKMbA121A
eU7kDMucjIoEsF2pQEkhIAmeT/8PXttEeTpZnlG5fUO9SLcC3fDicsDlEj24TKF1PwedBbs8CX07
xZjy8+thH6MYJGPKChUW+4CJv8EWzp87J1G/Wy6YJ/tuEmqdauo7Dz/yK+bnCYahNnq8W2acKAUi
ZdZ35KFw/chtSRL4ZVp5SHvuBixy54ponvS3d2Stlcg0CQjDmjfAldjJ0FtaK+YSa7pN0W5042+T
s/JGJSNdhwOF3+TsTul/mfLVTkk7Gu1oL/lB0bbOoTuhqrcGvirEnJp4yg4XGX5YeDiGGdbMc9ML
5f7Z9YBTPrGA26C3Fildat0wfQ4E0HePi4tZMbcDAOylnAoB7ILzfWAi2PbEUp5PGl8NrZJ6LmGJ
tn+e0U3yx0VUU4vWrAX5eF0R0JV5D0PJnP8Q5sP9FZ8r6VtFYhCR98FWHwMzbJo8G7y1w+MzrE3f
fGtMf3YE2Pl57MfD9M/sIqZxFirFnmUMJUtwQU1aLGUIZYxsccuLZM1J2D9sJ8+l/j4NC8W7OLKm
dVppZE0IGZCx/k6zdjG0ogJm7/5hIbTwWUe8koCkdRD38yE8dTtFSBmMiPFau5kqNpXzADE8TX5O
rgmCZ+yzkdBkt18EmY+TzCs5nv05OTDR7N1aCZQNC5HA6aHEbbLI7BMIzahXfckH/l64W20OHKzH
TnalbBPMsV481O3rmw0eoxywYqQpCveBkYRAfZCNmXZC5kKTo3KueW13bD3l70VUd2Js56IF/iZs
gsAThC8+tGH/B5+8J6WbH9IhUb7SZLTVibIp8NwnFoBE8o/zY8ZsipROEDpWLvNEy8cs5IoqS50X
F0l6xTMoyGV+4ZGCiCU9d8N7lGp7gD7O+bNrKGPuTDq9TpX9c/6VfqKAyifKBOk3I9B7XmidUE1X
w3qsN+XCRIscIFb6Sa49lrBkpw2V2PDd+zBvbhq+Rvh+0Ylu27OaT0rf4O80sUmAfB70SVNfgQna
oa0/A9LnN3XZxaGj5p6DMuQBhmWKN9QsKt6AdYYB90LMUYwRDsKnZ1n2mt522utG+Yny5yXs0TlP
uwC/mxzkcEHlngRT0L4M5oWdcYegUC/Zh87fVjvm+WgeRXcqWEmRFm1EfL/CNsUqy/DfcD/azc2N
WaV5fKwlBxajOxICL2QPvQ+xkQISMFFs6gdF4MDVTcSq5jUGYpwkoaKlQj7f03n2bN2FlwY7+YUh
ppPjDc5O6o5zTX6eVWrF2CxnTLfh9BYhT0OEYwvnP4i/ATM+ftcuVam1E+hyOHSgPTz7CbdY7ojr
MZGNAt5ibDA/EXPqmzxvgV6FMgt095W7X5fQymIaiVJ0wvIzDqJr+Tjwn7TvztTKxcvhz30LUEfY
Zsc8Tv4Z95mn2bjy2j8CQufnPOeWgZwWJfIqHVCngtAHTgOO2OEQB6eSSUVaHIHx+EUm6qu67S+Y
iwxkfEl8Goj2JljxGIDcMnhxxKRdKXMRsoLlEFRyAOdkTYTsMHZnRbdIrkjRWThLZfIHtYrSKwaV
1pqv698ClVrVue+t/roMQM/Z4lN7KFzh/O2KPgU+XPJsZTeyrKboM6VreBLLT84uroyzyFTTU0oR
B7J5fD4xeG4bs5Oi+bcNb914gfvI/ft04e/fEEqC/s72UyhhEDIFpYKJswR+RWfbMW2unyGMC8aB
BpjeQsMy2jk7iGlZ4bpwpeQhOV9zKvAAq4grMk8Cu0IjBe5V+NjslJ08FSQLg7O6OgQ2xD5CC72T
VhMdlBVDkYwvsXLZg44Pk75+yYTfDi8MX8z6UrlyrpXD/mMgMoxVfV2juYscZ5bucLs/oJYU1E3v
tHrns16/IsAvMnMnNHhbV9Hudgl3LnfRSxt+KNTN/FkzJT+DlRCwDwaN36+CAetT0ZYxHjKp4lOS
ySCybX+bpK4DD0InwclLDfpoAFtCP4/BjAROWbWRwpDHrzh2wkqVJmwpCU1iAJogB0iwgKzT8CKD
tU5YfPDlhLmehP64bhA38mxP1uVs07AlBa6trOCq6qSaSHYGseqkIpI/vsLQe8xiO3OUF6WBZ685
5Drbpr7zd5IpLwSXKRyQ/8dw5EUzD+8lTtZcBl9GdYvVDdn68JWKazrjFHlm3cDPfbyGL4QnM6iZ
50XpK4jRLoZKCKjncyBRnhe3ZuFaBtBAzOetxuxe+1odk+sSXLtMA4liwmGJ9JDllww2DvGFf4y9
LYwQXkhvHRwEpQ/hUClgowm1guI9+74D8cJC2ooNAQO/nUQTjzJe2GkZtLvmJVq8P+ognTUh6pW+
jQDtIAREyjFsAPmT7aODwRjZVDl6+wYcJM857tHEqClQH/DLiGHe3AqQREpY/OGFpWojPPbIA6lr
reJ/FmiiFK0lwQr+aejumcs4P/pynUAakzEFtoMso22czLUCM2jqKllZv6S+gFgcNI9eyECqiZgY
/6KBeET0rmTNy+dn0huvh7Ky3GDFN9fd+U0hIs1s/m3WuhNeqBISQqm2iK65bcpuPE3xCyNSFQgw
57s6UF3lZJcF2yiTT11k8sPpr/9HJYGrsU17oFg24+LTKiNFWSHN83HWTggATL1jbb7ctsv93ZEw
BuloVZyb62YWYRpIJKcBiKsAsQRKYLYtZw/+WgSoUZQRmMOPnTPLYLT9I0vg9csNHNocHzOJ28gs
HIjSdpgBm+RthsXR2SRmOaKYxRLw1mdvZUDffmEEQzUYlAe3fvHo33aG0Fwv6ZElQCuxXidrpXPG
AtRB5FKMauNsWmE8oMhB1dERbqLXlh2mzI0uUc1J6ynrWHibS1sLDPZ2ZvY1oHBwbFAKdcrQ6Ow8
mbog6WOfCyKf7diN3kjuR5cVYX5lxY4mG8Oe/P62MRMKrvQnd5SSOtJlGxCAOl0x/oMnwv1CrfEF
EgWJPdcx1ArUXYEWs0pNz1HwQigzF/I7kbK4toKs9gJk1T2vEnbv43aKLI4n7H6u3J8WrduuoIhV
EvugqHZEgSygmPrPj/os3tnySCEAZB4a1Y+T05+qhOEmh5PiLz5i2bML/H9K2dgd4QGKAIr6R5Ts
GgIMP3nRqvCwQWjt5JCg6cx8d1ct5sFn8oJZ+AbTak/9SruylpIUXwU9kpQhCjuUL9N5QuFI6I2d
+uugaaw0pJXFVJ4O04wwNOWqJxcv66KFJF0ASxvxEgz/c8pVFqojsWXWGatSjgIn0hSFSslhilNT
QuYUlT3grr+WLuszJZ5KifePMb+h6I4jwZFbVwQTbvOQVZkE7sdQhNqfFAfxNHcTQIWeQeCRKJHZ
w85jXZ1AxF1LtDFMw36iZ99jWEjIuzsYpPlxFOVjLxofRy6u0F54WFBr7ejXHFr6KQXiVydXBF47
yIBX/nVXINN2luxT5UNvvKjy/cggX5nxRvFx4dIgjY/UzSptJu+dqbfOYmHdf18z7mymAHVgJU9w
mSRDjVMIseCzJqTDUx5g8AMf/+CwpV/VhGlCFqWuh2o+pIB/yaShDQTcd2oYjGQHd6uWQI+k4E84
mavbpOsAoGswtw3FobitFbMrbRgjV6jyxAZIrtLUSLr6KyhzabTztBTopFp+Py01NE3zLYcRVjXA
TYrVd+16PF5Ts5YA6PbWr/ZfjjFtGKIds3LeN/tnZlo+1nd2S7NVsd/pjBcvJ/pVffreWPTUAWiz
xTnZB7aKnG9Bf3l7ZuBbxG36uSY7nmeL356gaFFFORPI/90gsX2smDvAsC4b6LOb+88u5VC/av42
G9E2Vci7tuL130M52hM2Vm9gGnc+IrrVg1kE0hFg1w+fvWpmloYhn0z1FaREG5BfpyzCoiIYlJYq
6ZcVNCdwzc4zCCxSaUbnW4HCMIeESiSISPALsoJNn3MlgKktIDvdYBYWhk/dgeCwqmNdGrxcY9MG
2tsmVCgwEhhSDdQ1RmWDY0nQlcthKxsb/g8Qu5C55GusgiE6x7CULW+15eC0kdVP/f+dp+eX9o1M
ejbVR12FTe5g4V7JKw4W/jsoC2ubQFy7fVbT2ThpJDecgEDBHek1G7O5sG7l+rYMKEicq/U5nNdW
V4pfeOzSqrLkn7PGhj6/fKeXHUKE0FsxG8zeVqC7fX+8SuWTN8AT8VKvxOEZxQAS/3zJCPPG4RzK
lD10ujoJyrSo+ajl+cLMejaBi3bwpxgxNLmE4PeQHQK6JuH4UzHLFCJlBFsfOsBrG1OK1ylI6Der
8YZ3bq5cc45uFDotl78boXHIWMVgocJIqdVSsKskptZVq7YwBShaN8lmpnoBo1PhNh3EQ28deZhJ
H9XK2J2k8gZkIVOSV22LryBiLA1H57IX5sjCQIkaiiZHGzmMekqkpjJRYszvaIf+9RwJwmIaArZ5
DzOHOXFEx5Er+mcyaXGxr35/DOp0Th5pHMogpTL8XszWlJoMr5HB32gnE0Vila8GNcj5U76tUKp2
DXcShURHFrnwNjkVYHSvsI5EKifoFU7NN+9Qsox+QYuj0TT1km5cBwzgJUF092GEcakVrTFhm2H5
vkd6UAfgHS+zGsKJpblYHvdjLRbIhnm3lDCl5LBgkhLo0hz0lkGJs1uCAcIPpo3nRtU6apkvPt5G
A8w185od2OtCla5YCCqOysu7c8W0zmaZzYFM+veHkjpkeI7yKaUplMJiQWbhOlpydp7OFVPsAMp0
95P5aOhqjDt83w+VlDDg4hsFbX6yn0T9idij9VAM/s37i6MbGA9VR7tSxvrI36M8wS+jYo7oGoTd
/syIZz7sctK7wmU/+B+he/9DSHw+2N+0rIkRnKdzZTy1cZBtNlZsgnSAq2hTTbqA/0CUj6jDL1J+
Ok/oPVVpBHnpdGsgLj52u1aT21/4V6DcwqsA5oimNEj564UtYQkbCl+7CTY/Uml6w/hHhZumFuQj
Hvr9zt2zJcAskktNKjbuNnTlLTU6A057gGyr8vr7xT3+ZQMmM5pVDPmKYl95JiwhZ6jqbSdsnIQV
Vwd0w93pmWCW73rOpxo1E6v/+LboxP45itGtDtlFjscCf+JLgFfYxTnmMVzdoIS85uLnwrqx+9Dw
X4rIG/LE2k+V8AI8VhTZj0cfverjzjzXqZwrO1FwxaQo9TNIu9fufmJdZk3YLnAJb4vWsA33EFsk
JP39yi5rzdsxpjFrIlF5ck4WhmiMnnigEsfd+EfMV2eFsUgxoYtIcHRek6CmdCDFTy27+QUYZhUs
A7jl4hnlK+553q/QOuDmgdBs5ash/wpHHZDny/EqLnk+uVGe8Nb3BgOsq4FTx6u1UDkZEmYeHHyU
RInmc3R4kGKnNfGScVWgNZbp2Qca4bIyjcbq96eblzCwjl61z+joEfNFE7rFUnc5h1tVmZxS2KnX
zSMjtlkbDs4qNbErP60BFseFsoPWE+U630en5fLy49jMN9chzTs5RRr/j+A+h1dQPzdHZTo3q9/f
2nyxX1zrLKx6bnpeDhikyCH/1TrT2CXk1yjK3zau78DraJfuiTb34zGJVQ8OLsd8B4IJzw8o3RTj
1AbxRBBVC0gh64YX+8arXtnKNP5cW0xaweuDgkq8PZS3xrvxxs0vLn8Q8o04yiNYdEDHqjJypght
q2NOzi7tV3AHcMTB2bafi/g6GxM2qZmF8JUBYl1zoTT7Cd0x5jjyafbepDh69X+2Pe87r2DQzEgD
At3Z8f6SlYV1M2QWnUhNMOMQy66WlwQ4iWxJYh9pYpB4nlCvdT/ukNY4o788WLY7T7xkUr7smzll
i6+Z8E/5lG2cNRGkP4WucXVImzs4I/MetM3hW4RlBaxlRamx/WtRMgBsh4U23K+PSJHI5BRWfawA
tK32Uzx2g9XSUG4bAW9dOBjWwLCyUvqMqHET0dUIWbbYMfjkEreWcN5irnEBLeI4b/a+HM1Rddnd
+Xnix9CNF5bfgEOUswm9r6rRKJ8VjJoFBuR3geM82njAKQUqNINojbAIIGtbZ0eSfqPena4UXvau
KZiYMxxRB0Vuz+TgQEvKiZyICOXCbRCtFgWW3U35SPCrmta16N+46q4JFJwyQjJjg5q8Enc++aJM
P6UPPwliKbZKxDJz2W5O9FzPMkuKUV/eO2MBl/U3qiu9XWBorexdLCeclLLP4mLP4IlP5dkeePjj
XncpFH3UMbQJ5uqTMQO/JETSowXWHWMTKrnb2b/irXOW09efGpoCCUYwQqOX8S32xwf1mHL0jYpk
+LDh/pUu3ml9z026cX5XE5KGCuHQu7a7vJ0tTLxeX3n9r++QR+T26g4DCZsMBMCkYxgjuVFU6b+Y
giRnKsv5Ugp7RMFHjtRZzseIaFjt78YYhsubpBcO9rQtFiUCSpZZzvMOT7ifIBrST+HZ+KaLfi/4
7p3r5mxtTKa6plhRT7qLZvZ8XJDPnp/U0wZ7rmSfOl5Gh9iir9ye+9diUYbyHuUQDGSj82V24oTE
KWaACsJTmKCy8FGDusei6cJfmcdkVbDdl/lpXkfQi+nxNAPMea6re9TzdNPE4+ahRJVTdBSI4VaK
+5FRHSD2NHFbYROPXOKerW7HkI49eefXJ8xRG8lnA4JhD2l/MeerWdbo9l+ePLGtgjIhCtNk9hyh
ER4Ef0MgxzbWhbDZVz+z5C28h2Va/PvgdTS8jmIe6QqxNwr2Sj+xHFeM8qjMMVKVoQ63KuXotJMd
zbKHetstEnT5yFOlLnKMAsgE6vR1M8v6F23RVONU4o0B5cImGAcECplhXoEZMcmQA7MEWoYlAHBD
Zp2sTcFULvVP2pZDzXakedZ5oWB0aYh91vmy9NWZEi9yLHoKbYMYilik6rO3tZQzi8sXZR54oKx6
sfkY1AP5VUDMcFDhnmyxpALWBw/PWNjhX010INQSPsCvBYKUSdKOLmZEH9tspiSYmiM4qtudlwCx
iR8jhd8jHMc3MROGy5e8Bo0Mtle7Xxd552DElZ8+3wqSFtqUEZqByKX12Py956/wbDHMoh6bWvzt
uLWK8r2/yofvl0f1ipu4WljjNF6d7XvwTVSRPPicf4VIx6Z/bJcdmE1E1hybkDLf7J8U2XPsxt3m
yVHjpFdOiyq3KDx46o1dPG5j1GRS+IS5dPcLTXt6VHiQ/X/5CXuB+43cR5mr6xdnptzC6vo2SdcB
RzR7S2FFpSocvUQsayMG32Rst3UzANudrQhoQYvaQVobRo3UrN1HbVOsAMTzqCRr3+XH5AoKUlfU
H957STQ/beaAErCEWhtmYDa8scILCu5kjBi5IfDPVfJW4pDb+rz1yTRNMCTXSctbkVSwAWrTDChb
+G95Luaan1gSPlCCrrd60/nSSI4bxxhtV8UEew46bO8f+OQscwJny9vNjzmFrXakXBu/q5DYbqXT
sRkE2BDoLTCdHJJjgUigDvM+4OKcWQSzgf1xD/xrEPPd3ZF4dcj//+1nZVZBIa/xzKiIBkdC72Ui
sZ1tOZID7Zp3avDX8ExCXRzUIBM5N8wJWi7dmbUQqHkJX5L7uBFZ7IxOfnwKlSuOvMYNduVceQww
7v/LSsgsNm4ZKI9HG9pzVv65lts/3tkfqyDEwgZ6BjmjcRg7s4J8G26KiIh7g5WHQpfuRoHgnLgM
cde47rMqua84thQx5QCa7k6GBm9BTVEhAjXW3hvIruGdy5vOTMhSJ1ib+J0okksjqDqeJcYN/YZp
4NOo7gR0yOkt/tciOvuGsY6AyLmU84y3uy4AvLdu5/2eYGk5Dz7pRddls1Rqq/X5fQ5imGa9EVWR
mVTLMIZQ0fFZAe45Zjhc6sSbUPi3P8P9XvqjqfH9fg67F8Il++ElvK7pVbQCxkmlIT6MATl5cyjw
fSDC1GkKrCBHcOyI5a5o+4C6mdszOKCMlsyNe2f9r0Z1I77y1CQtyupSo2bvKAHbLFPTnG89ITvM
MOTr9ImSxAp1+dhMciANqTQUgEgcnKSLQVC+T+1XmwSQFn5HEN5TObH04mhoqhN4ujCJwfVdTtEV
QNaUVLPO9WMVz394GeGf2zMbq/3EU2FzZc5SF5DffA0m1pF40JgfKfQaiaqv41H6WraO/zvk+HFs
d5kRvdo5tolS1CaAj3FlXPYQML/j2dXGBnIHa6C7r0JxkuJCFM6LW17asYp1J1hZGWHRhR2vdD+D
bV3dRS4XTtZvhb+0qKx6im5JqJ9PUIBs3fqij/X5dJDzZ0tYgE2k9PR4Y4SZ2BtxEpxPY1rnQxUB
yaqwHr9XUJYkDCGPgwZXSczzINBuePkqeS6ijgk5WKefswjm9fHvDAKjgoTRfDf92PLRXOjEgO3A
bpQTwNfp2QoP2pa+NEAAWdNfT+KdbcmdJGXa0oaNJ854SIlk0lt44i+5cJOQl2sfml4thRBtL5MV
6QUxnddOGqQdyStKssRPcn/Bx6gaGyyRSD5wNHDB5XRjDbXweltjrZ+5mmzchi4hCEAJ6zj0r59j
rq7/95q0GOaOCZp2u/UsLDIX2slHd+ZSthXMgwDDzPHoZqh32w1Mjz78ut8gLJzJgKsJJYgB7e7x
L4WNoy1WfUCyb12hkT+Fq6Vt195OOSnlp4CmB73QyENh+tcZrPaAB0Pfmf2/7BVZTFTQc7lanJTs
15pbguEiuYc+EHIyw0W0AkqMUS3Zj2ed26rRMf0nHj6spNVn2vcL9v5V5wb7JAek/kaUMHN+JA65
rDkLmFlGgOiP1lFfM3/HDTKyYVN5ZcSTXhljJ0aPM4cS0jeyLo5II4Ily1a4gODCUUjk2L5YESzX
c/zgDLqtBZY/iMO0Sd8UNwWAi7Y6z2Y2azDuuFVgB+lLPfnB7YHk3dKa1dqRx3N+2NyU5XCV0R/2
oqo/FwIMkJ7s0tMhdz8QJVBj/dh2dGYAJ36nYd2yPSPtoD7rKJVcb0n6i4yqjW1UoGSM/akXBpTV
lR4bmlB4x6IfGm2HCW7yEK4PAHIQOmqrKj2bnltoDNllzNoCinsKPALa8KGil+A/29BOEiHJjBnn
AosIE28NLA5U8Ez3mz6qe9L4lA9AJGbZHjmtfl8QteiMkj0fe3CRe4gwzix/AgHTCuGqIhT7TPAk
E9dt/S5j00mHH/zh1F1bzKdyCKUFUPQl1tqfGADCuU7DZP4lyzDeKlMSNkEeNqvDxx/88ZMxsmYd
bM3ZrQKob+/JUgVJQ/o/CFzEyTqxl6agMIgTdHtpIROEYo8HUr9zz4WKeBVGdzTUoQk0uhK5xCwC
AsQWrO7F54u1Y+n2goHceIyiRsfV9hu4ZST525TdkcGA14RjaMuoSNOu7LyPsJfOd2iAtrjpXbHz
JBmQieGFaaBM+IwZy2IOAVzMH6OnHND/8aevTKLtvPe8M6VaCPOEBo0pSbm39C6paGW+/vVldWzs
WiC78t3/fC2bk10ffvnf8LQ50Qu3/ecTgOkDklHJ4NzO6t3F8VXtMHq6n5X7SC3NabHUFw3yo95l
L8bw9XF7kAq0p4XWkf7b7HlQDa73jXYGl8nWbnetwr+HfeaVxxabmSVAl7z4vyGEUBMzyMTexrxt
J1k5PBlhQ49krMSwrze6DtCyN5rqMIF6b9kEde/qdw0YKUmSGZkAMPtGo1xLDAgVPkCNwuRrHOIN
U4NQCt2RrHzdGkAdW/nYeumuX1fDQcs2UXX0weVJ1dgaRqlWLBIYhGNJp88+2+EmfWXURVimIEUx
7cPB6WvuASCyioZ5bbTWA+foTTeGM0KGwlTOmc3gKM0HJC+uqRW+1fhst/rGzgynLWNx5A+igXdd
pn/UXnI/LfHVAdytOBDpAUet7SSlacOIQlxnJ7qt1Q9n4gYAyV1sR50zduFluRy36ezgv6j0nO9y
SqqZMO6M9Pl7bDAC6kEAap2WCV95MBkSM0ap6WFFcpovKZN7ovvVMPi9s6KT0eD3zK1sxUGFV59A
KGUgDnzZWM3VdQw+cCDpjj6livny3g4k3FSvHZvNTp+1pFegdujzWjPGiqxZcqBgqMC3LsWGPtX4
QqEa4kOk8bvZvRonzITW/oeRRiV3giwyYdZyyuX66xXNvaqw8NwpRiZ72QQCD0kh57zpkN/Djg+C
9RnC4GHAlye9HPFSjJTovG5m1iRG86RjalvP1DTaollgnuN/V20Cad+NRgOn+yWro88QewDPNwcX
jalHSyonuRuA6nN47+LgtDnnvfsWU5fjskG0YNiZRGkZE268CnD3t+Wia/eVCwqz98bUtgha1WTl
bIpQFAe8CoIVngqe3paECmRZMKjKK0svnZ7h0v1u6yGcKLOhJS0QfzoFHuwNW8RicQxaoTGtKlBP
W8D38NgKbGMLBoO73eH36cvgsD3K0I64YV6ki4w7Kx0g23Euann2ovVfyUMeXmAezU8RV4xH+rAr
CEzEXlPZN+3kxZpPwPePO81+wHnGYP2d71PmeuQ60kuCxGwdIahRTyWlg+c3GMJ7yDjzGyotb+4y
uXrH18zrNUL0tvVvwSTnavw+qtL6tPX7xxoyZh2/uSgIAChihCSdlLyE2tgMEy+Ivde/7+E3PvBa
b5CMit1D6ZhlLdBbVbaMRCDqFUA5lFXoF2o0q1ApPmIM3DijGHLJ9ksYU/DcnbdfX8p+1jkuLSiz
M+ITfGChZSjX0z48pWGDGPwzTdd3otkFhG1qETjS4JJxCNLXOYNPE7I27m07cHcsF6dnKUImkVFR
I9cmTFubk5TmYeac7htrMa6+I2RlBWENhGhcf3WnEEBiuGksCo34E+3KNFMtykltNTSwMj5AIwZd
+K+ClwcPo336gmZoTaRnfslWd/8RTw/bbj7DQwmEeU0TG9UsZSS72eA7wdLeDardaLioHrzEesjc
fkorQkiBaSbbsLQDLEcbxwe+F1fSo+oz9Moq7s0imU4pQ72eAyP5GA9TBrunxuo7YKtHFhm/IKJ4
OJWZR2QKhcg2GlLAhNQRUAMuJ2b92eGDQuwNTbCbFYF2TVxGX0Ic4OhLiY+dp29x5T9cKu5LDCH6
EFlvH3MUeTKcNuSQH7tIDT+RT83yPS8MDDOpj8AeElStUKdRmT2LEjJnWUkB3HShDSKphUBcxtda
UhGKMacR9c6wx3QiToFG/JnXeRcM19hcZpzSJr36shwQcESeKrBi1JRTqfj6D/rYwOw25ObjEIDS
57QnXcbnEirea+ICfgWYU5OTvYaFomlMHMzxs8Nlc+K+kT4aGwoyZScZYJLWDk1Fr16zGwH+KfFA
y7Dxl2yjiarxlllhIclum5WiEa8aV29DPeP15YfH3r9tuOpMuCl/xozYa88jcwTLsunmXXq3BU2q
6R63pcdP3bmHsg1T5d5QVlzuEW/4acr351rUO/4MkQLA5EOnnQ+rMoz1KOlNZbcB4mG0GDe5Awns
tx5zTvMJp+goOPC+l/SvgCjYYmY6lpOlL8aN3BGaSpKFPYDimTuJnn1Amj6tM+kx4i+DylfBxuAV
VA6VxvOyZ/QcQHW3JB04Q9xXtGFX84X4P2fgN1QjmRC8y9tDHWCFoVLd/Q/FNCd3GRHJaapg/U6H
SZg/NjlUTrfb+15tVlPTcQFifscZmfPu1z0nW+8Fege8g52xvIjlzDqE4xn/NBMHcLpg/1AKBKKH
luCSAAuVratuYJJeXKU5FraIAz5UD9dJeAxmhyvHEYB/5TtJnPMI+Jjd9JZzbndKZ6fjjrmZ0zOQ
j/bGRkuS0ABgv7ewwnfAvGgcLPKQ27aFBth8w6NhQVrHDmEJDI/XM+TzsYCmtyMBZM9xzFZtTm7R
ZaDP0SMEpb0rOjGd+5HuS19Ll0BkUtDcexTzScbHwASFjcNS2CxHhAWjCzwY5y0vDcl/GxHYCc4i
qV1y+Ot661gaUluDif+oWIkCk6sJVC+aMjClKAfSy01wPoVSzunTG5/DOYaFJt6a1Y4Yc3e/GxiO
ph+dsRxaO/102TbvjXGoA1+gsvjhUVHsfEyFAvKtq4VAyL7jYvYKCrSH5yhUzfMPmjFE9yP1MRNc
76PBWmo/i1bATmmAGzCm8hJ2DB3rvxeLeyBIBgOopmPhVIKk7ppATJsNgf4t4cgd92XU1K+PPin6
wTwJeWUMrLaBUFp2e7OlT8Ukf6l0Q0gZTXlsG+03QIS0UquS2N7EmPvDy6Dk0RkuS2R5K7VNAapk
qs9cAnAiBFWQqaHAYvEC8lEXsqcGpdm6dLpq4VqslMAF9AuU7iFWPaOurUnBZRP8f6ODC4TPNzkl
6A2yA3w8zs5L8sH3iPG9BGaFVO8gEHE3y55P/UrXxyqtkTqG+SdP+M4hSdA4ea92TJuQp9ynuYBW
GhlfdMSwRSSWCagFIUzaqo8yx+yE1uEOO+YC4a8g62XRiIH2uz9yrV3mRrfvahkwJ+esnZ/EqJSK
vNDzbSN0YotQfpaxGkQyVtIt8fQUgQ14GbZSvwjw+91grSUcLDCqfppnHLCQzSa6/WaoRM8ii3XF
ML3Fg5xNn4D1PoH/QlGVcjUY+wneMBlzrp1uUHL3mYNI03gkwKzn6YNkxaWZq0uSalSdRmzTf2yA
+g1qx879LJg5MxbxQF41MfcQpJaYGwU1fN0iDb6QO9VEXT3c2KvRDtFnkdi7/PUKWraPnTWWEMag
+A2hEjlwIxhHYRrvZzhwT9x2l/hijPH/4JZxIhPz+SpHE7ixLy0ymA5Uci3xsKU+DLBIa/Gw+D5d
Cps34ZwvX5Xz0vBQUocTo+v9ZvjY03+qdIjfMtUE4yrdFOKhlXys/usn9WO91bbS9wUvKPQl9Tm5
uvOdP5w8NO9j87Ev8EPHDRYg5nD3hIUvKG3bGuatROvYI6zJzxCn4fxbJ+acAOo3GG4/DQZprlPH
dTFHI5hpcenRtyJuq1yDKjnlT9xzuvnG4GwYu9djQbNw9LeCWPlEX8g9nXKZ781ponPSwkxHP3Gu
5zbN4tfNXiFJ6KYoaOwPnd99paNjnc8vYzdCCopc9/oWqG0VxynTV71H1PKtJr+XJ12CC3LaCAfa
yIELyD7Yz0c3i2GaJG5hFT7yE2yANWM+NlbeTLpOnwrmqcjvVzPlgttoXBJROKb2lkjKnvGa0vhX
+zDVVrhC1l/o1RLVsV7umE6lt4g4c08BaNSzrMnTorzWTECwLIFc0WRVE2n42z9Ka0wtzVWjJUgP
vxasfBSLH7fnHgxs6BG3tSfdA/XVwc4Wr0lf7SoBEXpfpR8ajrjFM2NZEoVRvJ2HwWq8t3MBbYRn
4QlK7eN41Ta9sHzeS2MHkaH/osTHz7gy8lLmTYlLHo03sr8K9qQ8w7xRP+G4x4YXVFwZnhUXaE71
o2h9c/3ZDoBy5KFJb7moPmPrK8H7F1x6ZwNGAFho47i9X0gSyOGvNtwt7+SvT7QSDCAxjoiT/sM1
rwu+W1GCVTasU1x2oMYnPqQQBR428rlcSS40bWIJhMX71iS26/4H1SOuRdXMXzJwUOJxSrX8L8q2
mcSd9sNah+DpPCdHx4G+P4r8vorhCqHARcC5f2Dq2M0RT7fKAdutbx3T/uhlP8R1Q8xBujJaiVr7
MxG0QW877BGzhpX7tlllfm7aiJi3RR/QG40ww39PuAzHXF6VMGhuUEnhUlSHFB3h7X4XpzxL4D39
SjJCyE8YVtxdyRXV/+tX6qdCWSb/JMTKBXsl3+MLt/Sf5HyqJwlktvVKeqTtmAkhhcBfDRCQMZAq
cw++BUrZaz/KACxHohxxgcDEVn1V30wriof+b+9l1sNQryW8CPiqFDHBRY7YyewoCW15FzHbRqIc
HhoBlJtmv66h7cLeHHjByw8Rw5K7c1JUGvwQicOb5JXqgZZ0lgDgznyep5Zs7pfslIVVDQFDGTWy
8sD6RxTFlPCC1ESFgUYTGcKdqnSZe8RLEr65/GI190ebIKvFVVvqxNBFjwAq43UO8NVAMXo697Xi
/SEpZ1Bo8+RLjb9dsXcC9j3ugNUJZZoYZm7Y/aV46Pbhls8rLVbmIUa25k1aIUclXj+Du5dE6KOx
uek12223elMRUJA9HmPBUp7YUlKD8OR2geYIxYAoC3dMkztUkGz3oGSqVkKCwg93KOE9Y7c/1/5O
HRedGGhiuclt+0s/4JbTKUK9QXTPKGV5f4ccO6dl1jg4O9PkSur2xAqOBySn00fzGdtC5Vps4Gv6
ISYo8htw3ncRdu9FDvrqYB9cPJ0806d5AKwXgw/OPGRhFaUbDM72/OLcxpValpPldApPe5dqlOAa
t2jIT0XdujWrkTSP8d2e7W7ySQxtpJx1uEheisOeAmsxK7ACPh0erTwJ3VBD8DWVM1lTK/uXuoGy
jEqewqvLqbGKTs0kGgcO/9v++wJIyVN83XBzKvmU7uBecgvA42IuG9HefLKRI7a1A1xwuvuaVLPL
bBjEovDMZHEcXkNn+ddU5BBsFb4msK8Tk1Fa6y78/r13WVkniY5QlA1S3s2+tNit7gYQm9pnz20y
Utk7Hl2MIVqf1nLV6On3TRR9HgqWcqnEMNL2mHXZs4+H94CkscAGBGvi9Mh8qoPIybgGXZm8UoW0
BKc80xecQ5xNsd1w0AVN3zgIcax3TwLPHhvSnhRfguC+DT/zgl1bnhTqis0Zasj3qVbXUP9+dBH+
ELAlqSgnBHrtyFiNBswHuehqWUqndIMW5cdQDZQ/MOPR6pZD2y2+uzC07ZJ28gfSzHGQUMamGhz4
nVsTC9E6EvUehmR1VcfMHW0BqNkNDLRYe+Im8IvtCGy5bYAZgSw+MkmutdFWYnIpx1G13pUxeaGr
1u3ngVbJ/HzEYoadebQqaXxmLaXi3Q+DNorsKFg+GD0Wloc9HYhP8cSUzWRCz/fVkC1R/RKmcLiI
Fj/VF+pDFZk1Wzh8LVTqtFFNRXrzp06tFpigSz+MqPt71Jdgi5SqdCdBjHKg8XJc1T0pAOcaHUeu
J0iweodupp/8zZdB2elOrsxpk5i4blncU1EIH5Ig5+vHODKNdWrIY8ZSMhrhJwyt1mGxmDldlCUQ
vZViNQIbYE33AXnLdrYyQ22tEsdQmOTK1vLTFD/FAWPYek6dNmexe03xhO1UDyia0S6KmIneAZNF
8QXspI9M8t5qEUd9OuA7NP7CM3ehXfgMCB2rk61t0AnfDZtjctPqVufIe1vH71PGZ8kPUs5OLcHR
gzn5PIDw8Sy14Btmf6mCnwMZGdvauxvz8HClwKT96VelyAhk88lAjW8aVuQ9Pvwk2Ji80QxZxqQX
nqBQn86UF0A6GBGW57WP2iDMutDyCj0hMuOIdEN5JA4LS1L8gBT5d07Vx+IE0ZuQzCz8l0TycfUb
ThlMwmEVgqA1JzsMHbImq2RC1URTq3GF5OxjE8jF3XrYTj/hV0NA+QqeOof1xV+fiM/6NSd93shc
dI+JXEzDH5kIKDXovPMfLG5gcAHrbzlPrIxsC7Mch5IatVbERQRnnQpNHDG2x2lXwdUNXaOEdiAq
h99v0JnGl3mlijJtOD/VxGyxac3OZlmfUIaihtGwjbjgf+FJAlXgERyLdaYEw7EPHn9uOjozBdLk
3kQHZZdOmRaXHRbMv7Y7Q68tn1LT3WFzdTtesnx15nVcvPO6SpB6nc2VHQC6KutGhzhoTiUqKURI
Y639lC2tf4EbNnx+SIz8qINKncv5dJ4znl4hpSyLor8T3plVLlN+HXk5fj69G7zDdDtdHRrkUgMg
AYihasfnHIQhrkYovLMYi4y2cxYsceUl4aGSLGMhayaamsQfQ3WA+0xImLZKlfIkopn4rimtHB9z
Sb6x4D0VDB83UP2wpjhHkLY8EhJ/onzzsmTAt1ITxM62X62xgeBgd6FSR0NagTv9dMUB9exQFDVY
6IRHXc3tRaJlSyjz8Liaq+dprfgXb/I2dm6gAorLcJV1EyCwhHdWl+1ej1ux7mYvK1QSqQitiNuf
0OJfBmRdTA34DoworJfzr9Os6noFrxwvlOSkHr/dMN8nDnUrRXKc6QHruN3OdDPYSiAirTkt3GaS
X0Q15E9caenvmBnW0YyAFxCLHaMlVMzjSMeqlc/ViG9xnl2u6UId9dysYPQg5KAsQq3kZppZlbME
ZFSrxZxfgUk43tCBJb7f6JrzxoHx1IzH06QAOMePr218GrpSgg7CklkwZo8YcZ1DnT6eAv3hUcrD
4kE54aFBSd4aefpkq26fQdjS+vwHT+eeSvPTUfQKwR025SoJlEeI0tpuz5ZbipVWZn3CWWoZhDwj
QwigTMkFy+kqI5TY15uKWUtFRu/ilEiTxA0+vYkFwv4kIWsTIfGq6/vcVi/Iasq7bNr+KNqUdfg4
kpX+PiLUPd08UV4inJM2N3/o322A7BkY4pef12Zs8XG1mwT6feyAFOfGKLebfeM7kjsIqR2vXvuk
oO95gKCP4y3IGrhoVuGAdfSfDuISdRn78X0DLT41pGNxF6CmgY17aLoIG8l+SCJf37X7mdngQDpz
jCRg5rfZmeUt8m1Dx+zNUSN/IxMw1XUths90SBawW90G1+fdfNbPb4iBa93GdolBvJ94GacGZOio
G7cwWufFdpl88eCz7+8zFdZOjRdwf7jbSw8KisnJmJP4pbKYi0n3/04l8PlH4j2rxDRBQKBEuzuN
bsp51ipsjbQHLXUQ/XOTWeNssi50oAX40AeuEZw9H5qlG1AmWa1Hd7XSeaB1Ivf9c2t9RIlhc9G0
9npus4gkFNnfdgd7QlABPZiZp5RxXvqZNn4qCftWjsLO5M4aR3y1xqBVNpcQ0/fCZLN1X2C7+ypw
HcVVKyq2g+gNHCzYihzbttVbfjnHOdYedk1UVOGIaaHa20k+GCPjEJwZ2VBMGzZjEERYLF6utzwA
kSn9XRkcNiBd9ZRBlQIiI7YRP2EYOsn9lF2qeN+oZ/thu2BslE8txPZ120911JxOcpUUvVnIENTE
7sSyNscX3NLLPARLQvDNNs1gQybMd9m1SPja1XUwBlB234CqvcoDrFBnrQWG6DI5Epki3zcd/ntN
1cIxh8CN80TWYMEYHcb7JQWyxToHCr8RNo0JBKPIhgkTS7e0GXfAUDesXCMZ+SBu8AQDLv38kyG8
jP2/SQQv1g44kTa7+zN+JUEZBbmxzVYNRtS6cxymInDXLBoUC4lunsExiQvQCVtgFwyYac4w1ZKu
9otXfbsgMbnXFdrMsE4ECBvu9yXxLUFcdjL5TAPgg4VwzVe6RCuU3KXIvswCXBeLdNEbh91/K+ZJ
ut/p4wUKDrA/3T6FITsGhQdvp3zghM5gGFLB1JaKIEx3fYozJMI3R3aMuomzCha0pKJmOovILTVx
vKvkOu5ViYtKt78+2peyPE7QlmnT9mmdu3826x7KsJy0tX/V74S+S9gygwJOqFRbiqQQ4Vl4skM2
9NHd1IC9npO3MWIRYIuT4olrSJDoIwIvYML2mKsEvoEP0IWsO6xFf6Lcd7tj1V7qftguef3U/Smt
gXAMzP2NFu1rURK9uro+6MYbrtKSEa7IccW6v/sCAXvca6gOI8TxoCau+nKgVKOELQtn6oHO+uyb
zveospZfBSD+uGT5jo1KksFyIRa0+2im10x060q01PkNfltxrK36QYF1sgikZYFv5g6fPNAldUGT
5ciCKeqUEyGjFuAu9RIaD/wgykbPwkjEYw2wnYqVXtW4CkdaBM7MErMIwJKDz1MI621HPGQeiIQA
HSXGZxhBkXQ4m9vlAk0vJTtLox/WMtPVTJ2R9WQ9yAiPOOChzaBQKI/yZYjWkjOV0Fd82LtpUeT4
tygiMDAZIMdxGwQsgpV3zSrgjsRpugF1lAcFzkFynMvYZquTTCXfPtHZwYFl7CBpR7XhMYaihmT0
FkvVdwizLCtfPSSryD3aq6XoppXVGGpprJhSVf+bscebUvMziYimIUqCPHfrqIcd0Ybfbdx5DYMv
+jOVU28DOWt3GvD84mfHF9jG3YyR9R3g+d67DHVWlhlFbTaeMTyWTWOZ5l5qIAgpigNx4ua3zIdV
TpFIzM6O9Hl0uES2nNRgd8c8N8tbHK0rD3PW08VE6W5esLmoJ73Q3TSasAq5Q8yO0PH9pV8b3+/w
+Vpewmb8yuAb3M15b4uGRg9/oTATDACiHDuzn7vmlFGL2XVvzw6oPo+exESKhpUQ8Jk/cNEwggg1
s790Z6+oZRBMj5t2gZQefKrEhc09iELdXVWG3igfrTTaeyiEGRjV189yRfpHvkkFgxD2Nd27rz16
f8UhKWQQO9hHguRm8TgTjV28a5XMlJp+trD7wlsXdgrm93DXLUhdisT6BPOoFIpODQoIWjzI71UA
Yy/rWNuknkfi6WmZkbN2vfA/je9MYEMngT/iQuKGoN+UzPE0o0jz7x31hyVWwV8c394S3Ux8fNu7
iiHqfGIXyiir73WW2ytSAY15cpF4LcguI2CVD2eISDqTfyWM/5lg2xdF1vpJkzEIqIXVWTAuVSwX
xgGl1ZnMPDBIi5o5XQPgLRONTVnTFYjrrzbftKyyycbbiRSJ4ra8JKSOxCmEWNh05QxJ0OFcuctl
aZU3fBbyGRT1ZS2mBlCZLd64l2NmZAgL2N4YadiqcTU06ZXjAOeX0QPH2uYEB57JHOn9yGI2m6Ed
UevmuDM/YQ+mYzDDqEYF2hrXeQZkFvo2oY0WD2GtHheykRzfOIACVY5Pq5/njT66eOMZaS/x2oYU
c5pFNTIEeoCpLeU+o34FcsSP5Fv3TfwLXwyMF5S7EKU++G8cQosI3X5FBDOJUEf7ijqTojp88LGY
2lXClbd3G5I1+88UjAPN65C5ihCQHwUy1fwofGoLJoq1WAWPYvYnGNdVlcCDMTNQdrYGtk9R/u1l
oct48m3q6G/7VGI9raTfzd9dzQG5b011mqiWslhVpf7kpP2NgCQ28AhMlU6Z46jUpOt/AUlPsPQg
1pN2prUXZZ/Rg54IPe70OSI+qzWIxsOF/Mczlkfpn3tD/b1+MJXPr8JnBfZLVkRahVmTSj4EQiof
iaj/A6e8axgHddJUVFFJ+71LOHspeKko9PMHNI+tEtPW1Foj6cbmu0bBwfq5Ce6F5LzjKSSDXcuh
EG7T/GkhXTra3eu1snkx6yO7Qws3VYInD9cWXSTHWR+1JUNeiDEhHNKk6EhUALsK0hxB9vttRfsC
6r2pGiS8GhLEEOT3zaMjH1z2/30hlbI8uVHQ0YnkCASWhZPh8jOB5f9cSPSw9Fe5FUJGcHy2jh4W
428H4Gz+6Cjo5noMGwgtCYdEdLJohQ63H8xzrAi+mD91gogEKnikAuKsgpggStq8DxyRFI/IYTmc
cchc5DPTaynufmCRNNSoxQ63F58AnlGrY7ngtlAbwjnjHHYSafUm9sfQy9L8CoZ9h4q4UcRlWOm8
jIOlEQjigcagah0AjwbCoMlrTbt5/ziHKzrHDioTGlo82W3Ul19Etj5dTI6q+9166wLBBuCI5Axt
7L+Lnft/Cc1NXoTBg8ih9aH7biwJ0l5d9uXsRhxJ+q+Hw2qqUI10eBRz60AoUjXX3BdMkjbCDBsg
yBPIVyJfbwPr1EgeQ+aPAUllq/+oIM/SJ7jScSjLwlVTzo6gyoJgKJ8vCrGujFdGVLlrv89Hj695
VeU+/hqjr9D83/e5kUq5Uot/vLVmlRLNiDBNtFQXWuMa9/i8KW4pAjmUEo2Be5tMT4VnqPC1V7p3
MHy6uy/j7iEahsZmP1BTBfXe5b9kqyLD4WXbnxA1FqUSUtc+rpNSQAj2AwJN9CCko4+/82C9aogj
bYU/2ieHlA6j+WupAGsDVDWC4JsCtO/YiWkXqLxij51EOfkliw8vNAC3brMp+BjQIR3KMurOILST
SJ2iDgHOjjE/74xm7Cf2dncP8T3PfP7y7adnBQz45IpryERicUdFMdqGxZjqZkLnF0vVnkjNdQUG
qDnupXhp/zkTopIRM4y4pETVfWn4GKC9QFZV6p34eyxehcE7ZjJjdVImW7RswX5ZgU0PyJK51Rqx
rSp1ajL34pzztFdcbIg2AbXiqfA94p040GDnIhbpj1uHHSnYFZJDuFvtpIGbvhk1PFPmRPpZJED7
+nVL9Xy6AT7w3FtEgocwzVth2Ag84NlPrKKtjXICSCs1IXcxsQ2NqPQWa+ovgc7Ob4ntddAqmB43
vzVFxyltxPBymZSdzfXp81W5QIePLC1ouw8h4PcQey6M/y86mFQXH3Z8/u0Qv4sI0srJVtP+NjqZ
qUaLetNFMmKK4q4vp7CuSk2hdlA/TVl4e/LjS02xR0/nJEFR4vz0xvIljBXVsg4BluAn9RrNA67l
Vlwmin495nYXLiG3XxwDxowYNLi+pYAX8YE8zAQkwBoeKoVreG6SDm5HI+Ho71hMg0IFE8RyaiCl
7M294hB1Fjr3JFMNhTiIPFDR43VKQOMKqFsMsVzz7m4Ev9/6IltsPZuv7sGShfqvWT51MdgKgOC4
9FISihNwL7C492DlCVyi6Rq1jLuCzapCK3x9HAbWQdCs97xWw8O+H1BNrDFa5nHfu1wYFplR9vBc
cnUgoAOOM3jrCBbiXJYG0yKsD7OgJlPBFZdme65TaNxl0ldsHf0jDhnUKJJO/mgoQ8RnAZZCj8yA
YvWUJ/WfMDoQWB0s91z68hZTjP7l4RcvfnTIf0PajMbPXuN00hbiFMP7k7V7M+DU4N31ZcDwZGG4
RUMTKJ2L8dpVYfjXYgwdUxkzirETnzefmyQQF1IPX3oRc+joJSpJ7xZ/hYziurlLTWZkWx2b1WXO
8hfTBwuX1DNXAhB+fX4eglzuGKF1A6EdhAElwyJXzBeRZi9Y3pHBJFcMx9TTI1nVTHyj77L3Qay3
bX/2cWnH3rQVRrwSKOHXzTjU7dC13ubfJI897kyPb2jYATpkI//d5mYspcCuPG76XfCjke92niob
ebT8gg7G4UxfYs39jJhK0B92+QTTp8x1JAAN3nOw6h+xiZ1i4FToLc+2MWqURm734xGWre8XFRnF
hbY80CSfJL/kNlIHoj7GrjbP7RBThD7KFrnqF1VKqNisDPdShR3ZmJ1lX+8H74itJItI1ip9UKKr
mUxa5x/FnXL1hXV+C0El/HVuwUCwLLY5otp5bX43IhDpYQQv3IrfLr7ZuwN0PcXzQWHhoux3n58A
kVGFxC7CYKESW6GvDrmOJ+8diQX/iqqz8bzTzVyioQv8auLv7eakImGEOjW8TSY/CjlR5dqiI2RL
4bS0tWzV/iPa6O/SBUESG3lp4ROICEFoHCHXY5YsNcnmSHTWIrYq+qYcmU4NQMfBYvLOJ1J6n2sr
ZRm7Ujr/+It/31M1CbuLjBME2JqGrRj8y2eRE6NvEM+mN+dGYU+Ibkzk2+tMr5DOs7unIxE+XW9x
X5e/eN+QriJj9HlyPDKvhuzH54v3OVZ1R8BxLvivXMYeIj/pAtLP6zlBNpcu6z5Bw6o2/f0zaz1/
EMuFXdISMNv5eSodXQMDhGJj3gImBBOXUX18DizzOvr+lGxkqtCh+xtVJ3Ws5QhrVmV6Kz/RUsX6
Inp61Ebu7H2vcY2h+X7IofjCAalm2aa2Rqr591iWKT5xALzN87yRd+xQq16ZK/2X24sHrNUMAFAN
PvQYjDoWCJZ5gxqAkP8Ub7gkQXhyaNImK9UB0VxPF0jSx1a3LF9oM/dDNroz2gyqSHU/toIq5PD+
qzvJayNkSzw6vPqtADKS4IFFM5KYq4tKFSCwyCHL73aI9RHBXgQTuFZN2W2IK4s0MTFfuC1wABK6
WoyaIYkTCchnykF72rr8uxbNAh2OGv9DQaOZXe03EuUalajLtA9wBShcmCputa7Xz+32DmfDgvu9
yGgvBeX7d8ooxF/E1eS7pUrL8R5FFsBpywLj/u2HgRgCSeRK8COnuuu5sCvXIG0IDcYpJ7C7S98v
MXwPXLl8LDhCdCx6ASxDoKPxSgM20YJRBajL5UkXK2AZmmuTzn8eFJi7t/heHvz28nfYL3PxTewi
zwIFVKb9WleEh34KU54sjLSN9ZL8yW8boMf7EjSxxJKOsxCzqN8Fqpom7kwUZ3efI8l6ZWQrQBMI
xy+tpAfG4kzjsiw4IISFRiMzu9n8J5VO44jPh+eA88pFLF0dopmXF0VRxYMV6MITv/G7qg707TdY
YkGXO/qe0UALf9D7pjmUiFiWb9k5AlzO41oDhYEVDwdF85kxCVDoT0ThxPV9mjs/YHkF9SLyDU4y
SMMtmipm0EhN7wBGohaN35epkAR7PVTFG13YpElNu/szp+uA30tlBW57fytZoGIOvL8f3Ne0iSOh
Z8edYb1hFarNM0cEt7rdeQR5Sbv2hkpfGlRX136CiGqSdBYOE+nhEQTqyI5CZnQC2W+K8lIyQOlu
F7oSuawg5MUqzLYCSfTvHWPgwS+CMxhUCAjILVBXtJ1UD5lsEdyapXcnanQOLaUMoPX3a4UWqPnS
E03f+JP9aMlUXPuCAvU322wqLuRhzTOeyCXDyxRC+8+1QQCf2KMfxuOCyJerJNCLkxANDUuumV1w
fjchwIap32G+l1VwsD/UKH6EK6zipt6/VlzoFM0IlzUEYvJKxv8MiHeZJuDrHRPSu701Z+GhBZHJ
BiIAQCyQ8GonUN07OtoS3PrSPiIptqaqJ839HFACC90sT328wtM84gzFa17jgLNbUuomPFXRUjcO
JLMimG7u0pyenZvIU50oVrgKEY3ruCvoL3PN4ImBKjsZltni9wnafsXCoDXQdbz3Nw8kmvllvFMC
0DdIXr0ORqnxInhLzGF/ed/dU/whvl5ApWpyGPO9RmdOHF+P6DaqH3NsE/06GR+ZEuGcO8Uz4i9d
KVCb8iqFblOA0VBYg0g067eTTToBtVVnAHnHQqM1J3HTIuZi8vqpGosi6nltw8x3EonkBmnafyd+
P3tudJn2T1jrdCsto65QkgZbMqwB4wlRWQINmrShnWicIn7sNZOdhYJ4k62353WqEWN5Qci7Fn0E
KZxgjK4tacqzjpQul2HB+v/wChATS6hZttHnHzuMCIjQ7P6/+0izwpWxdX3iL1m/FkmG62nYhcRn
bd9m1sLi0MCCkqiB83FXOpt51B5Z7Z2AhJb7v9n0BZiIzZeQd7mxdf6mGXDNjHTY+ggyOp3s8SBP
Ooe8t81jh4kgnJwekwHxTN9nfTK7pgkHdzz9Ager9Rjm5EOieWKkQKGqqluReD8iOeer0Mbgf2r6
cvdcxZhFtOBTV1ENIMcFzVJyXuLSw0E/HTj40dl7ucVYPXEeLoVdEUMiTD+6Va/HevDul5m7dHab
u25s/dyHYL5q9dooCtTar6e1pF6WpHVucR57Tg+ifmol3ajfD74AssY19yrqXNaxe3pzMSvNJnq6
Tvn1qvNMsikby5vKJZmTwRngBLAV3/Sud1unPch70YDV09i9OU4fTTRbuv+ztm0Ljb62WUy5nFQq
sWS77ZWszwz7Dmwnw50PRMDcPlRVhOWp1i8EO6IzmF2OKclnzsJoyQakFlZLj4ybBxevYqTVqNNp
cbD79UpF6iHI74VCC7LZI5gp+WsQXi+6me0bVO5qmdKRfH2E7QdCQPKI9mTr6nd/j7k9G5v753TL
O9tI3enaMO/DWVrRquCz236xFe5dCn/+OX33Nt+0tyH2XhveaOQqxQVkHxk0svt2poJ+S767kw7Z
ngf3ErcNtpxvcGqtm/DGU8e9SceJe2KYVw1NdaNGXrWhpE4+KTIE696S5TAdrmLfJdVNxeIGA8DG
/TUd5j8vM/u4JTEVpZ3bDmQAco/8SqCOZ76FkvQgDhJ5Og5kYUiVdGfxegK1chucrYdurLXAKnMT
kcBIdlH/UkyxGQidIHT9gt6EZhUcR21KsgzWEFC4rdXRbwtjcVR/OHhTNGBBMXYoWQjxrGBbZVGQ
ZVfbjJpSi/beie8n8WhhYbn0SXdOQRH23JNgqGs6PAENvY3NMGB4FayITnUZoJuK48sPWEKINmdd
vu123AXJoBX2eRGZINRO92xh49Qg6kY8q5Sgw2gbbZAjYY+VqQbeNib6/+zc65Qe/YSSZjK+SL1P
V5GeILiPhZtpIalw3V4kSk1v0/TMKixBhcR3P2mlxJaSOcoPfHu4tXAnZPJBBGi0m5lfFUaFNn93
LV+yx+H9oObpUjrMgW8rf/N2f2AWsujkc0TSC6kjRUzOek41OhlQ6QksaVp+UNfLM4FlfqXOa8EK
SAOavhZXQT5eu6w03lE+GZk+1wwImXtRVDRydmvz7pxYMhKkRKyqIIx8GeLvrzn5KREc/rqTg8FC
8z0zLvMAEtf714mNvXHlzOMHblp01QdeqJFtgo6Bnt479pwAZbg+BEQRha6ofRY34cVbQtjhbW1j
jkl8Xz1HAWaNjHuQXMv6i73XKJIbvRapbqHsh782ig4FAcPafaW0LW8Pt/QwBp42DVwffrJldy4Z
Gf7jbNjq+049tR0EB40pvX5qiRlpAPY9bZqJwK/5cbLGRZ0ZYD/kEHU4dxGfOlrc1bZ4+l/bzuSu
uphjFsfWDOkT1AjPPL69Cz7Cjud3VW9vHrQPIGG4fBBUo+Cj3Q915XvnHCvMKFt38m0mE4tNzMwQ
wSnbtOvCXgkF4u7o+yhwFd2RgoJStFiHKstliEshbfRfKw7flvTjh7OzsStHdAoKjzry+70wBMx0
M7lz1WS//1cJ+jMkxEj/55kwhTexUT4JixO1ucgnI3JxzV8QANZpL4NfypoX7vB807xbcxydxOZy
2jH/PHRrwhoY7k842bjbj06eMBc+W6ujOHF0ka1GPjgi6eUGGBmlg+St0x7R+FqW6eDJkZppvyRC
xQG3n6yWNVZdFgqbsb6kAYVd4FV1a4ZmsaJ+xRd6ATTYOjL7XTjZdvD7fSP8djN4qqqspWLarCo2
rgS5GpnVwwJ3mufa9X9gUUTOwVBHSdd8NppVy1uA2cEbD6ewTEAQt0V345JrelitGvj0DFonZeMI
Ksrv2gvU9Q2nh874DFCkPAwURMsf0OMSk9cqLAyRs1zxwqREz6d0kmwG68U/00epyheZgXA1CQbk
dOBloCetl7gnCdPBdv6I1xNgQNqHiGLL1LQJyz/pAjcw2obOFWGtRyTaWGxn3IwM7i74LOZyrLKo
gHtYH5epm5OHLPEX+1QNGbg3ewkcFt+BkV57hIQ/ski4vuax5d2M1AVuyPQ8+aYW6BNnvNRRzIi7
nZmY1dmUkKMRCglaP9Y60NO1JLNIsgGfTxkhzyE7BqQEjelUe6lKWvTua35d3KC5rqsp2iosfiiI
t+hSENvhWDgGW3GLOz5N79z9YnHB8xrcN54eXHLdAhIatq7jt7wEXEhRQ6rNpfyxqAlGmeEu9ya7
2+ze0NwM0C4lG9p2NAbSrSlolynb2tTESB68mFgqF8vdmE0ERB8+dC3WxbaZM07aj9qwr2qBGEku
fJ8uWxzJyCZKzdMVI/FJZTzv+Br3NmuhNWsUhRaStWD2AMhd4rb+V+3Cxbke+6+qAPm4K/81SchQ
DtVGSd5dHT06lE2tbFltHYynJNMk7pWO05XiGkGAqh7O9Vj2DgsODIC5oWmhWpInl1VglfKs/jit
M4ZZwlAODCaeeEHXQQKaI5CmhPpJDmrHuqEJOTQNxkF6xjhIEuEqoH+HS/IEvGymkjLG2jAxbs9r
DZX0uJHefWl+QKYE9D26RI00icZ32MoWmfMJDVfYWlJpAfuQ00DgGSGuRaHtMP5yZBiD8J1ylWU0
tbjz9NkFA42yS+s9f6TibtERyQVoeijolZEEL5BX0cO/9+3YbgW1s0IFv8dQG4cSPJBBCDxbSEhP
gpOwM3u4CQ+6SSGHoD4XJN7MvNJ03s/QyGs9og4V02SdPf3mjc9o+je+U/wCMDKq1+VcsVnIAkwX
60RjTQ8HbpdXKOb5WBYpdnSjAN3tTHR5RKRlJ20TuJQQTbtFL6sQj0Pv3mhliqtJwUwZc0DbGFfZ
knJZvAc9HRiVZF25IweBskJe63BbUSBojGvsa9w+rAJFjqQ2KsQi8K6vHhHKY/ShHIiUOn3CUfeI
cEUJpLYh6KHX6cUlZZ+T7THf8wIf+XKWCOuNzhJzBq68lyGRij32kJiDRExGiGYRChWQh4uPmSug
ilNxUO4MeDse5VJpRnE4EvLoAzOHzuK7ScJGeQiItAzUsSFyoc2x4+4egIjYQpgFS46o902FfU09
6YfU3ZXaR7mb59xeQsgurFCCxAJ9CLLjVzbUQOoNhAqbHN9ieU1eYYBqzJIW73VUQP4+6CuYRj7j
Rv24jr46o+rrL6+/fFWYMZEvveL0oB/jEe3Rzr7vbWQ305RbI+PJTxBxN5zNFoij7lUNR+KAQ/qD
eokFKrGRmFnKhZNNn2IHtLAFI85zK7B8Rdl5UbgJ1o05SpcLQerHXYkUX8l6MZS9deHSzP1+AUBW
zAfiTMaaoF/1K8NeZm8QeeGobqGOP72jzFEBlwp2q1j5L5efgflOkODuolyxpRJp7FkWDSkh1dDG
QsStfr/ILnqwQw+huHqG18btfbQA+i7Vx3DhYv1SuPvrcy2rcA9l83hFnisKBCbB+HRRheuV0ccc
6AirRXTdRWUh6WFpjiXGf7y8toNrY+WOaXm2TFdyPkDizJyKMSC4Yf7za1rhDGHp73MjimuX1IeH
3+k3dKx/eKpCkZDkZFBL4pnhsR2uAHbAbFVTfBqF7o+Q7mq1Ns8ry+ipSvL8Ybaw5vcq4pujlGNM
GgsfxzzRNG5+JdOFt13MCC5kPinSmdJrKL50FzEN/su8wcUY/91k9297go4xrZs/hM6UqSvjJ5Rk
DxJMUi7bThGnUQ4UfqGEm4yYRZwRlxAtj/ZDnUfRUP5gAqhEgS3z2HuAdSB+HRwv4GbCqL2o8iX/
xOahfd2LHPzuUxkVV0HU3vudpUZHQ0x1RlLD8SFU5m0/Y5M412zeGm+r890cHQhjjp/pdifygh+4
F1ix2a/M/6y+/ETeF5DtjxL3lm68gw2Z89eIOXa5NA7irmWMPLMyWay8p88RWboD72APkOSrgHn7
bTHCJJX+UfB3zRjfI0+OqzAdKlxpQ1DG+2rw3xc4oIx6oLt//vmuUVJU+O6HAFaUe3REmAKGtOdH
j9x2GiydzawwQsV7SFm/wsZa+aPIxsbIw3F7Z+TJ4FZcfp6xkD67rkcoRHpebWXx41hiUKuCdcxG
saO6qlsPnLVtcF4Xkp1dTL33riCsECUqNUESA6nJoKbLOkzs4BQpPFrDObV055LnRiEdzBgM8tIw
s8E0m10ECK88H1BKPPBiZdb175FzAXBCyoa7WA2pVuS8pLTQ+RggfIL8lkcye7zb3YpG++WWveVB
ytmqVY9E86wCgvheVxMMliZz3nj3OLXgyIK2Dgh+OxXtjy5oBw1icEcpeOfZuE5HOxDkm2hC4eTm
yqbJ699F90Szh9MhShsaAKBmGwahRnwskgEbsTzl+zq/bH2cMIZfUUgPxRIy/22eINjJ0XyMuzit
xhYo3+Cjl/PC4cDdyBkHm6WdnzIaLcLM0tIPl0gCl8T8u1/yrm0SVfyGT65mQVIalgZPxi7Ptlm1
NxB7OiD6Dznc9DuMSAL2QzqTIOK/eXyJ5sRUMrIl1pB96BAExITdhqQ3XK6j7lVhiW6YRgx2Tbnz
osBfjXOmRO5W3eEWYEMkE0BfO/RgJvecU25hiy3aehHLfxnqmTWy0cjuOroax/zZTBZuVFybHBLZ
fgpzIaEhw3JCBIUB4wEHCUCoXnix3tRnoPEiSwAfKwWwTwrQYW3/Ix9s4EWLA3tYx+FzypaaPT4s
8Jlq3CqcP5L+8saGe1p3TyTkAECtxMzCDHslpJGdbpzR55fqFy7D8e3WK6zh1an+jAbuw0rdpVBD
ZpuSH26XXjYHAK9iMMFSum2xVlxVtVcZlQik9cYr76EX2eyzIkHwQy5WI9lHx21Clyj//jgB55jP
4L8DI8lGDHf3+7BCvM2Myl7iX3PSv9hyrOVjrLQyC2tQ37P+6NH0kyFVFIUSVVfsIHuYz6+nXRnb
aFIV+kvGrS+JC46YcYaghJZ2xRiIihKLBkIRXdzZXRyJeRKKxzllJXT88KTQCCYFAzdlD9SlRPrM
NJRFQ6I3pF5HG+z7pLOJztK3Qcr9jcTHAf+YFxnqtQ7WAQizB2A5DVCIZAKf2Mdl9vrT/xyhAXEZ
V/q9NslCFrgXlKbdTcTEZQa6gQnJVP3qG63eiMHXzByRoZBKRBrlic0gdyFlS4InbIFiDSU9lrIP
NDclVc+PZyIEKolxmtNCI8IMtF4rKXYP5bBZATyEWXV3mARxbmhWTIAMxcrttocw0vedb/P3w1dw
SQXJZ8c0Llhg77bLUPqzHfaQxkv88rgZxUunfnqO0tVaE3wzTpyLDrbkI7/3yvICUbSZC/04lbG4
KTnFgzSK0tgM4RZrDUe3VNki5QeUEO0XmQFUBbubeS+24cxZ+MuzTXlvwUHegZrepPXrFuDJkeQE
BPqINhfXfXfoSUBYgipfaTulyzBqXlTVHz6WTC+Vagcll5Us9zbrJ6lN+rsU7Ko+AhjKo/UTf/yh
YtVhiGjAWt6m6EusKVfO0WmcquKp64CxMtK9zG1Za9bUvcM+PpSdbPlrYuBRGIYvRqhxB92/Qxnj
LFTBFIZC0WnQtDyXuXRz8mSyWkywBi3GNgVXsbo/8GmjjDzfFQrgeDQErG48QrjM4kqNaYHEbLVc
lOb0jERcszviuGZNPHsm430UhDXgvd6xiLy1Yx58hCmCjcmPhA7UQddWbHxYTUEBcdwJdQKDoTih
Lp8ybDi3Mwr0Jx3/MsCkVMu7/YM8ZiBw8151UY7UwT2LByuPlslau7EoAp26g4dZFHzYSLoqaWCp
9eEhxW0erFAv8kDmHr60P32f68B/jcvFTEp98ld9+sygxmn1/xXrUfPS9iZo9rLxxiYijsmKZnqJ
IXVwypAkwHjemTOpPEz4CZwo5eUrPrvLtkvgn8tmGqDtm4YwkZYV8KpFQhW7yEw7TXiL3RFNV+CS
5kBWe6lOQmEh3mBU2QOlo5G11AC1ItPjymkO4OrUeRZBdkbhkEyJKdDVsQYpkRPwE+d9wCE14CVl
7WvnSdpHsVvHu4a5Y3KXLTPJglCgwicVcV86mZlSyqNvz1Y6RYMYRXe4jNytRtNRqSmMvc/qzVZe
uWGLGX2v5SjRCPxYFDj2mY0HSVoRPGb65etE5a0Gim7xkKLzfuEKsvDQQEAemfSQTSOjpri1rZmx
hSSKCRQwX+OnSRXyAAqyLNSUDBHeIo4QMll/J65yDZcSrXfGiRUewt12l8l72ROWSjkFh5TOXf39
fQwhQBXJfr1gUmUc+183hM60Ony10K3l7113OzaoTmwJBk6ObhvINEF2xwf6ug+Mp2En61zHuBns
/zF7ae833a6iULTCJUnTq9xGsh4Ua+nWroVE+A82PZOBd0ln2G21loblup6SJROWZMbE7hkbHfIW
1g6TeNOkx/cXf+MNaeAcg9RGQBKh7yheflhH91Uk7t4fSQyZkbDg8NnSu+DgQkRdW/gA5OEek+l1
iAOSBVenkF5JVXGeXbe05H1eTDym1wfS0VT/XgQZNtSN3978QXgMvf7C/4V7IRJGeCvsy3C6ZT/R
sCBkxw6ejlnUHuxTmRg99pKwcMJ3blpxgB4e0/0BSyJL40HjrUWW7+c4fhkWYu0MKH/oNdb/wNnA
G9AEbcCJ55B6077+pe8Dn5IVeXOXdxL9rUU+MmHXtVN75HKJXzLeFflsJCkA97YWibaaDX0Z2cRj
vD5sHeDGj3M8dncg4ZkRV9zyMBnYpAiV/k6uUG/ZSTbqE1f2qDHXKRd89hZYXUZC2vcNGhnUIW5z
N9ICzYA9vzezMlhByVG51kvgkPOCD5PQrMmpeV7CCmVVpE4b5crK7QPPQgp/4crRi0uCD232fxfQ
GVSU1k0dJ9Wfq6Pd9xB0Gom1vHiDAMo8n2HLMnkZVrVrlngv5APzy50pYVG3SS0oO5mvO1CWQoRS
PN27qW7Fg82pFpDqZhuoC65jiNWRf+oZb+R5vFXqqdnMt8+1aeUgg1WVgnn6o7gJaHF+l6S9pMPo
RGBqJkHX3cSAtf7WsNKBZhURLdBEidZ035icIVO5UuV8BTJXBpAYxFIsmNwxJyp4QhYLEaqOCHyz
8hjoY62IxDSbukLBmzg/POFeik6CsFLshXQtwdTw/s3fqbLjeiwBAQdAmRv528gzRlOOKtVTyG50
GtyGIWmqB0dqNcZAI6YjGD5e/kZTQ8JXQLB1/owqQqmoeYjSECIuVMBnsyd4FWQ9JqVgJ8c7+tMu
uRGCq8X4FmPP1xR4CPJRrHxviQTBb+YmPKt5xXB3Z1F2ZpB8ERPI3u55OZP/dHrMEn7lVHzrLI8d
bAFyfSj35ljc51U9coKTI01UXDnI/lj7ppzuSvEbIm8TgkYg+DvUr8xmwOt88vzGVoLwLvRr/JnV
eTiZTg0BowzgmEcmQ9EeHQ2eXdn7DzTrgMhG+nghdace+Wq23USNa+sjVTcyiUE6seD9HeMragY+
a2n+WElT2mjrzFCCsKOzuNCLwvtO72zDbUtd1vX1f/KC0TwcrkhuEUKae6RfXgz16ONYEc2b302v
qx0trUwl9B4UGSZeBlWkck9zLI1hfFp1Dz72xBARyxaK4need5APbiLag6U9Ss15mAOAAtGqua5I
asZ4DRCoJuj3Co0W3fd61EpjUA1uvMrdGz4ER9I1bxaM3BfRUYIxmNVSaTbBgzOzOIcE0zFWZEj/
+J/4NbkYRxZAFX0ayXl+oPHt3IUrXJR4uKz5GYmHjASCuL3nUgAmci9XE0hXIKXmzefdnG67h/Oq
R6JQ7Dy3r59c4FhLaqt7KzT6X9aFAaDyg8WDE9thciF8D03IcZosNlpZmATmc5TAqeN/Q4cH5KE8
konV6vDZ5szc44eltgqC34L5nsnlztyWnldr6drTazkx6AYrcl4vskGdQHvC+uMi9r0ctVIMi2sb
QehiICjTycylwUru4FqvQujrN4bIwdU2Hh7L1JruOQa332W62eo9c8t2Ku9FuBpc+5JPtAfT8cEM
6MN3oGaoNClXrDK7HJsMjUoiu7BxxoKU2xAfPLPehdPpBb6G4cTmVkL7MWAd4aeBNShDAlVSAwyv
pqMBGAJkBiJKBWaFFgIniyIPRkec/EA/Kmm1AShR0SuVGqAwmllWfYVEERvkU68kNrxdNvtfBJnt
88q+JErhRgHaDVBGbXK/pPmrvcChzbfCJgpqFv0UautWrT9Mtk0oY91auhjhgflIPxuPRloOZy7G
XcuubjtUie5XXohGWsIdf2TwzGfdydiZM9x6lWB88YF5vSltsugD/cxFA4gN2zVxDLIXJRo1QIo0
Z+t1Z5fWt4GSsFmr6uziF/L7lU5bHHX0BszGVTo6wOnbvJ6GoUhnFYUEqjfHmAb7GYi1HRvqMKXu
sGwyaAAad+2UMGn4920D0BD6mOyPF4i+zhZO4heggP4CslxHq6s/KbbAynePJfPIR2kF9WPDxaRe
kEhClg/2c4+5wXA/i+AiHn/Kkfd3Td+cM1W3nKgLCntsy4HqtpyxThzI+YZJ0tEwUguZq978f2Bn
BKhU2kF12cvZZUJkoT9sp7tMwYRXwVdcSftaUvAgsx5AC+1zH/+zXIy3p8p8xgp1ux86Z0z5cbTT
18/4zDwxnRyaQihPo3sfiBYGtQc1MF2LrMdmj01vNLLV1EfvzDQDcFJQgpZvhecn1GbjZwCnxPhd
j8D8HFNGmdEUHRktAdf8Uob1oi386In5Bo3VkvISzuvChOpUA0eknlkFLFm4MzM3DC/TbzUzCwiA
bcyfUwmcx8IBCl9GwvGvZqG16RFSnBQe06RaF97bxgbyxMqay+KYz6ANYf1huWFaSDg2eVdNuywh
0c4zjEfdJd6kiIHQ2teVn6bnm82vPGYToY7AlC7spMjktBDYdihXkRVTX99nqYioEvu2bF7YqWaZ
LdwCrMRzLSnJ2SxbDzPb/EOV6lIKlqrbyX7NgDgqDOEwfp/GrHAL28Z3FUwyU21Bqwf6tXhSuvLX
uzqPMT9sIjVABBBgiHMEzOBRh61SxoH6JQH7L77P0RYmALRIn6kTkaBQP/8EtTLa+6DtftRKJ9YY
iX39lDAZLl6zUG42Us9kFNAihnHjSdtNX9cj7UFfzgYDuaI56EW5yN/tGTEdqOz/75iOM1JM7v4Z
DWWgjtKKdpqiaa6ZUU9CHKrH+fCHwsvIqDaUtWoFaNvfeybKo9PoZSYf0jQMGXcPKmdzrphskGIZ
3s4Iw/5NtpRa9oTln3EyZFn+zeJGwfMdtlFC5cloSs6SZboeEqywMaH3AdaaOP0IyJBL3qJDW7je
68jlpcNL5xOIc5aPLwp9Rv0NU3YfAPSaVBO6MQuBwgDeOlFLGO48q1NbJDZXDRd3WDokXUpAI+Ev
DWzhtFYalKsIn+dgP9m5eKuPyhwWwuSGQWwUPjmbQneI8l9JzrtKb6zOYt1r5g8PBQPAlm/G48sl
LSi/OH3+LBKVaxH5Sa20i0es037KcNMsL8/Xu0unSs15q4jfgd7Zxg6NNCsiBTjs7L0pQ2VFKgx1
Z7VvJtyCIUeQTMzktyMCdA7B0HquoKkoP8/oLUbldN0W4hf0KX3K6ZCTYInINWw6m0LcvDUv18gh
EeC42fcAPfAbcGqWccmIn90ExKnMxg/kGOSW8c8FQku3ISUpjOm8GCpc69EgGjFjSpfbRTQZZWHj
FJP9MasVuZnI2cbxv3+JIcrwMXe5PPvW8OgOdewBIxmlsx2slATTJ0LoNvHG/3/weAkO8EZu5pGp
38UjgzU4o9YKSBuZr0G7TwIKE5MiILcyXbr3MF/i8XHVthyepQIhjL2L74NiYIPrSgC5xUGw/PHi
ruu8kiBeQ4YHg1T3P+PviTs6LufP/6QaM5wBJB/SageWriKx85kS4ifNnFivr5RD143poAfS5EHU
vc3muIt+Qmzd6yvbVOShGxEF/BqpNWYoIa0y2AZj6vxscsm3h1OCMuIvAovhH2WXVoPd6h7pZiT7
SsdK6CpCqB+CUOk40Vzq6CLpclxU06pV06E3mwvpAKwkCj4UDL7q8TIZ+wSdsse5/N9FMXj75zC9
x3/R0na2ao9mcY0ilJw61RjDEAqz+tDW5epDrgY5BSpPTJdcGsGSV4mYqew5KMOqr79K4EUHVOdV
Rz0gXQqqNWjPWpj16iw/ln5DnKCrkuGGqQk76lbzf1LeW6PdoC4lTc9CCGxKuWzJkzq3niUGO7+l
a3ZAwZfUeppAlCdN+nQqu9otVkNGSXHa143qjTup6LmcC6ofALf+EmcHPvBUxvjriIj5lnk5hFx8
6cqiHUsRLI6WbO5iLEfeX3lfKzYRXroVImJ0nk2tnK75mbnYj/JWk98ANClwbg+ugnHkXTLBPxYV
M4uv7q1LLfdiaWBwizZuNoXxS6Xho4pfrokO7ITGTEgUoL0KVj9qSLpc4ZVAPtqVJVDs4g04XYwy
ZrYsdAcj5z/HbKOR0EM/0irIxr8wHWEcGkVel8BAGyOgXb41F7nPegPvvgysAc/5bu/pxIyN8bTg
L1+rS3Njq5AIUbgDO1RrTBLfFN337dkDy8fsrQAKIB/nhLAmnaDhZ+x+uA1lWy0F/DKADSAc0ezj
mC7u8fNgczPBIT0ALhTyFL07LFC4U8Ak4ibvjpKAPIUMZpv0pYZBZ0T2uGcByjkbgd9X5jY9pAm5
6TF/aD0GHyNujWDViF7vE0A0FEDFT3FCRgDwPunePRKBVS2xxyuzT8lpXf1qjiZIltM4KTCGIX4P
A6Od2CVFgjibqK3krq2t210E4ATAZeuadkEsqptQMkgBOwXCag09GeErZti9t/+ED6p99sGFHzwr
80hZGGhrFGu38/x2CyN7Rdz5VE7Ted8Q6Xn7WeaISBE1kPRRVWDfFhvBJBPJU2ZfoYD4qpLgvB0g
jPC6HdZHbQM7Xl2dgFO1KQoVi3qpzVD7LRwLqxUx7fohqhLrt2c3S/+nU8EbAf1BMSBizJQ4uDj3
JD8RwLoGZIal/oLddy59se5fjo/cyYkh3Yi/gY1M952EgKxFaThVOIJV8DCPvRg1FBewPp5clYl9
EYh1afS/+CPxkknE41IB4fv1jMYurTI8TiiJRRTCzVGKmFtb0PxJCnZAxNHs0Eqt6CCUp8PUymCI
y8FsPGQICU6fsLcAjzJNvXB1mFuD/5VHQ7ipJVPytKWMCUOY247pKNLyCt+tbNUZqYvbBg3/Ya9Z
vjCHOARD8RTYrkvO5ia+2/4i3d8bY7a74tNNTnXXT3CXypYFIQiT+mKm6308AWjWGWQ0vF3L1kER
1kvGypTfETwZL9IaLiclYqdxqk3gOmrPhhaEUV4LjEO67InCaActIMyMBJlmLbv6PBFI9/Tvtoc7
EGSOcDG6DF9BxAgsXkcoQOoC4xwYNgDIgkkZ0gKAYDBmhTJ3LagxdUtcNnJJl7VfOecrUWjr+TVh
P9q1lEsI216mlIyygUd5xVV04l9AB0iCuFExtV6AVd65GOO6Fnv6lpqmtFgNMXGKHcFvxUAPMYqw
M+EZk+XXGLkLSQT0hUhtvAAxlNEVnjGZ0Ur99jZUcQNW6vBz9Ib0arrlGkaKp12yWHEsCzJHi7QA
LcavhZ9+355Hc+LOfV+rFEYw1/wYBHzp9ejVE2sB0zT6uT3bViEsKUFxTYKR+9CLXm2DgOmua2s2
oMfFs+hrZwWvyK9Auw77RflUcCKPLEoa4cw5HpqmnQ+N1ZDpgqhqsjPqmOsbacO3R5LoBrMwZBNj
XrMHA3+oY3lo8W230I22Mhek0UdWMM1ptkCL+dAS9EdwMXMa1/Vyq/qyXszVDxltQO9FmRq1JGNs
GoWdr+48u7Xkv7pR3tIvHlDNjJSs27NbLVhqIXP3iLCEQOyLGnaIsCg5dxBnmGnpJ7CiJFCeEyi3
noTRzpBxEIyLwDKQULakQyH32PN1OJbGu8Xn2KtVwk+zKlOkBK46hXAtJneXhxFXchu2g63hlEcb
PXAhWTRTgT6Oxx1HNw+xqdUXSor+p6ysNNdmKJdwpVhbw1ek00zKvv24HTBUVFXqg777ILeixWmI
MTjJEo0jruTwMGAvX9BoHOZuiw6gy9RALGG4mKX7dCHnvqPtVlFOg66pxU1JYXopYXa8eCAvC9Rv
KwZvTe9lGP3YmRmoBmnFr8YJGiH8IGCxdSBHcmTyBOCLSBjFnFYPEuukb24IbKjd9OKAHQX/zcJR
5cwBwlCiJHWgkhmCu8B+HugnW2reP3wh4vEF58cVCaSKRcnOQVYMQndL0bpBDYpWpGEyRLsfePny
7gVcC9+DKLC/IYfmXUcqs+xc3ReTBUVj4F+vu/3gYTvWkeCqkjz5A0qIyjKGQCure/zq730Nx8bF
OaoTBgNw5fMPYJpwoBA9NYeVwESpTGczaGwXD0rtqj0tWnlJE4DveI8WENw5LhZ1359EkSgqrPzx
+bjUwKGjGp74Q1eNpyPCQzt7pK/FptRgBDF2BwKDxovCjZ7F924YD8U8Bd7uTAogzdrNIxGYhHCH
WNRvvTLRMcwdTp821nArXi40HwGvJ7qy9Q5AGXvb9UlZ0OWhdkLwxL1MGrHG2Z29gauve3SqYnb6
iLRAtMqrButNz2KkUECnYneF77DMFFuWcqkCG+Lvze/Ijh2FToWiLDP0nGogv3BAMxpch0tU1U++
Q2sif12tKq6eKc5g+m0AfQBYLczk3uw7UHI3oecLH32z9dqLZBq9JohQGpXkGOjZkaKpOUxc7vEo
IV7kC5lBKzPb92XwPfdulHZPWhqjqDRcYBiCHzqh7aaHNFIrExTONe8a7UQR2hn6d9HQNT3SWPAS
gFQwZ70WlIH+3DQHksDQZD/jMpwu0Yimx0gyYu3fo5bVXpiHTv1hSRJGaPU48F6hHzu0aZNaTiD4
tdnEcH4fmxrDExqJ5wbEA90BxBldCTJU5VaOw1eeTZGvF6NwVDq4PG4raia7T88A4Zi/VP0Cfkkx
pVOXQnelBjjiFyAn1r/wbVfAHaaDTOLMBnK/a9O2a88KVzUAOwaXFMlxwu+w1z5I5/uTOLUAKsDx
RHcdArapppBgN+4iLJ9rPSQP8pVsuAyiSle0zKppX6I8/52rAlj2Cc0SgHjNfBLz3cIvNRvnbQwG
HkiH2qRV/AdRXdGPxpRMqvrsjCK0yF+HAfK71FMzDc/ymkTFhkmyy+IcpILCcCDp2KhkXCabF7pV
dO6owPowLaG3vmxQRpbGsilf1ZxhWRxDmS8fgu9JCOpcpV11L4xhIyzeepsKaslxlb4QvubQgqgf
3OgICSwUnTvfDpxHk1T4PC7w8maJ8ag+8cTSYkU6WwXnGTvaRhIK6JrWmrNUn0H61CZy3pxppxft
iMlGwy2u6PPpzE76G6OX2H8n6QYcTCOrmoqt60LVMLlsgw8BPwR4miP5+Pm7txWUuLd8klHV78fv
ijai7g78en+9mP5gJxxkiBX7S1or5GE6KMmU61lFsbbEZDTvgYsVi27XVTsV95Jk1ll1Zpt58JOS
SK+KFUAyzwR569h+EEFPrmD5qt5L3bGYZV5e2IDHGU2CnK1PCKkIfjzzrKACj/b1FIBr3EwMzufh
r2uFIRguma2ux9Ryek3q3jA6Ec+YONIiI8OXGDPKSGVOPn/+4l8vT3SfsBd24riTMz1AqRDjoo9/
XUPMxG5cWl/DdVbSZz9hBoRoWYF18GPlC2hWFO0bAgMWACcDBOHnrjDEusImAT4IZE4UT5Oojihb
DDWonT4i7PHoCoQHolBx44gK0MdQkibT6rGOGV86I0szlAZzieclPHgz2Ono2VTdfFOMo+OhMFOH
MG/Lh9LXRa2ypQrh3XTDaabC27vHYFvIfD+LI/PCaCkzighLxezBc5MDpjFTTJnMamtdyBkQOt0/
hlr0VPUBTcml+iKPUuU6c9tqd/tW57z2gkUi/EvXthog+v6kNY/oDL9t/G8rMiZVE0/zs0zX8nD3
jPBFpB52PFY7wow+uSp5SVq1eBQySbD4Sl3ODG97+B1jkYwa+NNRlUi0VSbJYkPvf/2wzz6tnMl8
VpZTgDuYXQZSVkJ4vlD8S3I0qc58dzbTQgyKBd9TbhD2CvRzYhAm7XRcK5NRjA8YTeLXLWRo5WN5
oyWduoIJCjSssBijOLwX8oM86GIMtrwWp4bO7uAzdHQFlk53ahMoirvXVLnRq1URogvAuTpbT1Rl
28q1NWhsJ1zueuIylEM1ixQfDg14e/CVwFquU7TUl6Gzy00mWQ8A6poK4w9rF4DAi9gBmF0Es6uc
NVUf6xPt8UtzuG8UVI1neHTv9vb7C9nCYN8pHXMd0NvOe+jdKqLE27HFDW6usJKOwB70PDbB7WQL
0hnPoImI58pF0E53IjewyQQ2g8oP22IcMNWEixUFOcxQzs/8jOAs+d/SqZL0dydzbNuDEKVc67i1
xObh5ZjgLA4uB2N/hXy3PjPINUGBHz2EAXhvo12LZmuFc3Gv6xpqIdxVHoja6VNV7vmcOSFCM86B
YHoW88VZyMN/zmaNIki8As4xu4h8TU+cgWfwLOhWxIioTUNWnsIcQOLKIAW2aOj8PduGYkfNDZb9
CW2WlxJi2f2YSnqTBHtwuf5BpJqxKseM/lqxal2P3L7xhmX9ChqpdOrJcJyRJRpwa8xUPajdQcSt
dwYly7NXDeEE+ajJgfpHyGg0Ad9IG2kkxXANSh8bZR5ScSCRUc/jUiu3p0lEH0If5WkkdFMFYPyO
a4t0swCcVItfFCnChrWC6hwuEgsesBjpjWd8/AFvopxmVFva4EbsLNch/BiRmnhuV6HfjR9nYpTR
qSuXggBBV+lWcpiHNrT14luysjaVc5euH5KkKxW3jyJObY0CDFgA3oPerWih6JNatw3iKw2O8kiK
d5EAehEptzMnf0JXw/0mr94ujc27W3qq4chdODtFzHNF0ephO4/cjAW+Iq57JomVOy62GZFRGBmY
hnWilNSd+Ji13NzHt9Q+HYvbQ4Mh2E0zvVXm4ECGfouDXwcIV4uCyK0jb2sEXw7NWgs+FZ/yRZ/E
BpwRiq8Rh0x+eroIa5S9jNOrhhnwVLaNJ1mE6d3NQvtanEkQwfKawH6WhV//7VpcBw/4KXfEGjmz
yHPagMpqfvwbzG8KncdAWX+6/6l0PavFGF8OnJcq52fEl2Gu30BWz21KHbyTYPDxZNAiQdKiBt6X
myIpPAPYRDjzEoDQdpVBtulr7TouxKL+FvM+p39GPXhuiyFenkh0uNqiCdT9K2bHDiTZ5kzmteZV
aBHDnARrBwB/wbulIZM+7iiJww3CTwyA/rtUyLRsnirrNHbLQ25kxoynKt0et8Om+cwpgC6E/MCB
LMwQO3Yiv66y28VG6iW6TLZc1DYBt/EUPrU6m9akymB7UckGVC3jys1U9yRTFCKX4BGq2LKIDYpG
fesQQQ7KANN+JAzM2StdEDje+U1TmlP2OvyVDcxNkqpUjc1aYNFVwwhFX2I7ny91xxnim+UToTMw
VPVqqmd9bhwm3mSyKC4Kivz82meqaebvyhbqUjWPTf99LNGTIQ4VP9wmpsEC10f5q3esCeZEeloQ
3Cqhb3NWvYn0tlCm08a8JKJQkxpm9m7q/F/yu3lllzq5ptrt6gaEfTjfAZfjiKNLvM4mRIoen0lZ
hZM0ZStOcvsAgabozEKWEvzx+0jEiP0RoAs4sWA2UQ2xm5sZB1OmZ2TPD/M/SlGaVPKik0F6FVeU
WJF0dI/FPQXBHDTq/5FgW9ginCMGYx/1FHUUFqGCgEa2o0LU55uRpx5XFykLS1wn/IVydaDhXPcY
rngVCJFtCxNlm+p/+SR09TCnGAXrzTZdXoK2RGCGAPgC77IVxVfxuF+kL0WI26D/xjl03PByEIKr
exgbV7bHhd+NNj4iv9v7lKOtRbbNtriFZR9nOR1iWekOAMfcs3aBjbzZgTher7WARFifkjm22tNr
AEw2+wsE0Hmp82X9laXnQt4LkZ52+0toWM2uN+zNjPh/bMErHEmrloZLh22a8+3McayTnqDbynMN
kwxqWojBdya2BhOmoEaLQ16u2CfYf5qlgVQ8r41J+bpPAcc8N1UIr/FSSyDD/EsbMab6+PlsLDA8
UO/Nry5zDwLT51XlE3LEyeh7PNFwrXGy45Nl0pY4WHYtE30lSUwNSrQ+ExOsSt0ynspxyu8A/1FU
4Mi3waF1TJqs6q3OziLaHh5GyxkJaT7Dld+56kCHdX89AGIty9Oc2n6Ow6Mqg8SIBw1J5Gy8mT19
H3wzcJxOtNdkkKfgFQ+9yF5f9esCNhiCp7UyfVbDeUpe4SCCQSiLxKct/Yj3ZQQrBPkJQbKMWkuJ
3KFy5byHj8ZrNZ6pC7mNZrnLOT3cOpMcodTk3Wyqndnt7JadcLDPtNYjfk7eBaZ9td5ulCSCz1R0
iWggzzn6c/caExTyzB93nXMRmqqaAsp4uaOEdrnSFmsjgR8ik4J5IZDXR46WULYyuZFId7puKHfo
dfsnhZyawbZgOuAt3+iGJawwbnRrDTh01Cz7DXeAaQGoPGYnvyRN0y9mbOMlamBer1TKP//OlNVy
PElGRvrRdhgH7SwlIzA3Ja/7IROdI0nHv8Wk3dwYOBArArbHjJTr+jluAw0huYAflUk4gVGEyHKT
v8Jhr0cbrbS5EUoSMdV49/P9wKiUsQ7+BJ/K+n0azaBuT7PxoxMdbEYjvbG3T80MDRd7Cy+v5fL0
XYYdaF9s/Av9MQvd8mOw4iT9XoprGstErX4aSeacbs3DBKX/g9P/ntNQKF2nIQdefoG4Ul/wkeLU
0f8WUzqxnK9prKSnBqC7sy8dmzMQEB92wPdF2H2w96yjNX2+P0QSaJfpEOt6xxRhkO5KO+Xw2Bq4
XhRH7PIZZvMxyBP8rhwa5/nXKZtdhYC+ETofhl68QHsdsFzw9H7ctvT+siAiYlTwGUnRHWB72/7m
/pV3REARn1ES7lEjhmFRzGLWsm5fZZYNMAUAeuQlxzouH2R2CbJbb/6D3jzU4nIdVxe9jAV8H46f
vowcvPuUvxgvvdIg6J0spTS7DB1YM5uKBRn9e++ylGapw2p5Bruwtlq/Pa7tCKAFKKk5ARSZbYhP
b1hgDk/IWZzwnLUXjM1z5DJ4Cio7tlMITCowxVsypGpFaphd+EcioPfFwVH9MwrcymF+Qiuaww9z
t8UKuHeRLsoWWPFRpTIW6fwN92ESDh7pwi8VUAhj+ba06NT6ttvjqs1JMm7/kbCJdvJhzzn4h4Na
1YgTw/Q98k+EDM7L88EigNFloJ5eIH5VrHfb6K0XXSHHuu9tbwOQEpzVC9SsVeEKKg2TVyivpMzD
MMxm/7w9eTNVcUZ/cGNPal5As6lrLH1MvNNlpEMN3/nUnVPXaU225khdkaxJM0yawWEqeM0x7jLN
/9SellyoLf6Z2eUrb231I6yPQ7dO38HkPwDa3dEy2nc76dwzBu3CApiEqONctr0qjWJJn7dYvz3R
NZxRuAvNk/EbOtUPQQPwwONRPA56i6IxBKldZw/03c0QcCFPIoJUhqQLBnrJoBKmsiukBqnFIzwe
VrHKndxO7fp8a3P18hwcOwu63H2LIiHjsZJNTdW9GyshLFrOhXFfBY4YVrGlbE9uafjuneVkGrVZ
dmlL3nAIOnGuJTPxrm0PTpBw0eZDfB4ui0p0rk0tsWXsM3z0jLsDH6xgS+CDDZBr/4628hP8Vmdk
jUWaNFbOddtZhKVqUVgeHtNJcp1g/rgCbuNYUQ0i8Ue18OFdzEBngjmoEtLAxPMrB9SKI6/AjhPw
DabqkjP6hEHq8yFmRXhuU6Akae2VJ3+fgh6hnggMivqbpoLNCKGp9Q8lspDUWK0p17Oy7nT6cOBq
e2qtv0ByovAhg9aujCGeC3N6kLDsYBV4SMYJgvDUX5uTZcBjADfFXXQR99wqhdbiG3xGvs4JttQ5
Ixb5BVyTcPdNjyyfaq5TcaZ23AcjXrtlyCznvrWOplP+1nLt/WRUXTg6IiCA/vgYDhgOYc+UtDGc
dwE1i1pF4mGIPO6ipHGVM7RfHtNXYNyY+NyvhWekpG7S0S49Ysnw8grI6s8F93zjnuWlEJp4if3v
xenhX28E1n9iOCHZNEFPpk9Q7n5d9zygSjlQw9BHGzrjulswiq8bD5rD8w+ExD++A4YlkP9H/6Vy
oBYqm7QyyYr+HoRLaJE9+5ySQSMd+DHrxngUqEsuupSNZnc3eHvZOSLB0GpJSZ5dFRB2zXghcnxZ
ayiL08E9fEI9jI6yatEwqgPlYi28hnuKuplYDo/eioeRFXlI4VNFsNkK9aT7ior1tVx4dpgOY977
nu7/38psudaIgvNXwzP4fTxz+1J51ZL+rDpH+1gh/nwueeRFelBTSRixNZogPgBK7BaX5OzmHSUb
Rz5ygj37wgf+dVRGr98J0wQ18/cgFJ3aVMTppfdZnaBWMuzFXCcJ5Tqj9snA7WmBMcuZuTzJStXl
5myrjjKXwnkAReMVWQc9JEs4mg9nKuPlzwOhODSxNjsFn/ik3xwr4xvFwQbZkTbT0wVfHtrJgdRU
R3DNjTW6KXP98rKm6egSksnmB1ot//B5uiclIyB42gR/wf/BhRHp8lxLH60iBQjyoPiNX9wj3igF
Z4VYVV6JjGQD05uc63b+sGFM4UShZQOKP1KVH4cAM9WVmhEy4Kj1RePw2xnYGCKqrgWFud4rPN4Q
ygm9DXp3pIjXuQ62rQy5p8ZJcbSE/Ua6UP9pI1QoncYIn9b5orOOCbLkPFHWIHzAWx8FlNkxzq0m
4QDpDOSTwCVEsNO3mS5k1qWhR+NIF11074GGtpSpRyIlX6BZr+zqi+lPj+VZmwBVCE2+aD2PCAfo
0l+isWB/t0fbi9plUoP5iNUvKc1CgcJntP6y3lMIyEEX6H8NLQx9aPyHRkGjHAc7d2/+fiBq7bB+
PjZHwviPQyPjtNLjUtp6bFuhcKavK6Jf/o2K6hPlz8yc9X5etd1MCnlMXHhpK1mvXvg7DD9Jbzsn
dB9JxkCKJLMQAd2wLC3dwe8w//n13yer7gRgNJinHVDZElZJH/TSQ7zgxswH27j5CWvxW3UFfka4
ZRulnRqWc9uRvGaNxfNktz3T4sSTqREtHD1euaReMQ45y4FsUfwc0WgjRDfHPh/9zNht5uKXykOf
KfRWQuIlJZvUrXTBWn5nCvuYfRxW+YIgKmxeuww9LWFHCn72/r4SNRjXLFOgAhKaW1EW7dqgsKpi
h3AjUB7XOjGmKm7CrBeHDhJpfkyHevvUDCwKPUGFZJ/cAy/AmoPXq8nCL8pOB41IgL4uYcB7Cs6x
hkW2leQNjWjbGQ2Cs8MLwF5ivfOC7wPCAeYTrbnjtrwysTjBmOCvTMBkT6RB9nVo4We/SdUgNUPS
73DPBMcWjx58Ps1D5MTn2HB/5H3SSgrTWeqYcvO6AEvVypnZ5XP8+UJo0iqbFXEaDdJma9s9Trje
gH4eCrk7AmSutjlJAhO9PYeP6hY4N2p+lEmTxGNXXgmWZVEJH9gWVP8lscEP7Nx+vZ1OWZnbcpyx
h+zMaXQG9U5opaeHmLNZPGxLU6SrgEaWYZ8GA2GJoDiDqdyVL9Dp/El4WqSD5+dE8nRgFzepXNqN
L82StCY+OmQ9fJlnJphAj9g0yCM/QLTJiSInz2Mpq5NCRWWwCo5OCwEP8rTISM/NWrKVcdnKhwae
nAMU9jMBTiXTQauaoce+ROk89BRw5PQyeeWS3XENBmJq+fzaPxg9qak6ZlCmsyjJQsmHQpZ7m7yU
rpXRI7JxAqv6w4CFt2NvwHRtLBZlzsK+Ae2pF1vytwkD4cZVyl2h7rsYM+mEpPHLDP1ZHTCnqKev
QNvMKEoN2YfVgskokptPj9VvMpogZj+2H8NkH6NzxwHKSaVEdtZeIUj9syqTWit6mnirZ3ZZSlkd
HihjE9vah3BaehqCR8n56hJ0ZyH3Ln3KWeCvviBMeaEi6hzTeD99B2TXajRNqf8OhOKR67Uqkrit
4Cx2TFOjGc97erWp0NAMCFCG8EvGSRMxC1tI7wuKpp9z5fWM1sQol/ku/9kSgsuSut1/9cNGk372
WKU4TJaVsjTnx3eUNP6V/rjDp8XNzO3SGO0wIfeiOfv7/nZtvU8N5FVRW13syUdydHqDkk1BLrGL
5ypShRXG8bmqQRjyr2++VwCDaZLorRebSpr5WFlgDLnxCAO63Ha8CIBdmpWo2KH+BYVPhOdLy/v1
qPoorw9ZTMtpTLFCR7rw/UEkYMW2eUhH3JpeWqnW3jm+d0II2eYSeD8SHcK3++UQkiPu4iGrRgIM
/BbGi7HxlqIRnktE93akK7TBNZDMMVsFKqR87d/n4l9aKBx0jSHF3aT8DWq/CsoyAfanK3+jc1ep
SgaSJWwpm7y4jFGGAjiuoSbGS8oBF3xTGmMY9mH4u633xsc7zQqPZfusIvWsSbPFrJBr0M3TfSW8
HfP/DHHil2ROPOhpex5/RasB3tUK/gaOQ1pSipGyYJjxTKcqJPDPCdYmDPs9VPMvt0GKwzPTr85u
09JzyhOhDM+LoGUV0EbGiSmetKfeH3DW64w3JxeNUhDzGa05xN1WLNiVFI6b6/eSMAq5WQy2TY9L
thOQBlOf+pbIwkVHC7sfp/C+5H/SiQG4OMsWaBRYKRFwvFyzBeVWzhqLDAVSakBaFFx9OnzWpqjU
7070pjs3LTaxEaGMkifrmHxCrzubyyjB7s/ksBg/wwOraxPmsMZ5HlbDb2gAvamFtxqFPoqRWprp
A3qRc+2wtRmR9G5jE8d8hSF07ebBYxNAQ2YBBDpuXmJQgmNSwjsaGGvAsS5AoHY8N9e1tHyrV/au
VlXelNpl+ZJUX/0P+vYp0Ski6mWsQuL2VaTB/DvWVHIMmUR7rvrNj104XkUOWgP8AoYa/XbUxvWw
FaAfhv1+nmcu8zlAW9GBTwhabkqrohwLrPkTmU1Tp0byUptzyLIZZFSj3TY7b+i3XPaS3S/rnCwO
OfklOvhXBkEWiTaYKPhuL75sK3mn059C5O5vNicbtXQyZjUN3ZVBvH1/0j0H6JcqMTBfscZdPIic
ZLj1RqGUKZhjduy/bfOkp2bQf9IBCracDlEEqI3BC/RthKbZPSzwh0O9GjB1Px8eZbx+Zh1htzJp
TKNTgHlST39vYlXN3UYk/f6++Xm+/oRTi1xScgsGCkPoem+aVI8cpfHj2Y4HLi7KBGaXHws46uLo
Nu9N0i9ijHn5fI1pwpCb2p7hyqnEXNiryVHO5Y9FVLG5yA9YIpHZ7h38cFVHDEn3c9gVCqLkt65P
041Jz/k9ebg9njIDmNvMsD6LZUxvXBtgb0YRmlaOx25r7iEErd96pyieTbJfiX6UOdqHzVY2uffo
LBT9BPC8tmk6Qu0td7649evdUlmTaQHSMkp4k/1e4ozcWYqq78zuE9nYbjlige9vbIHc3eG21dLD
tWiAlbx6qs6nRjqsZ77ZJQB7xdtVg1bXX/LHWVxO30ETqcAqfkTSYLik5am0yN+JAj61zUxoys+m
d4vhTxqvXJnF8Ws1vEKgV5QzuJszS6EfReMa8gnCazO83KBFqvdMjepGInr8xP+cy5pbRy0N0YRD
XUYrPfeflRc7VJ3k2wvqrZDUsCyeMxgltzpL21ySZ/pa8E87iw2rZKz79qAM9xMEILnJgibb4dgP
KZpJ6xPdz60yaZwrtHcozpKcy/6nrv3X7rpxKgY1MbV2GftGqVwrwnE7xEaaI0RCZ+MIGaYCl5y/
e+TJ1CWSkmcLuEsi/qXHgysUa1Mx9i7hDXHcxLGDqUFU8OXNT0UkM+luqA2qbslo1eFTX/Qv3MLI
GoB351L0Nec4za1hnMm0owmqz0+9AMOZMop0wsRu/9HsNYzv1DJYpfIKiN4BjeHH1j5iNt9zNQ4i
MQhArq89JPzbc1Jc1HmNaAj4fe9aBBd2HoXoGFpS+g6C+Knuqi5g2DKdD7TrX3lkGKQ/Q0+T9A4V
SKLI5k5lRDQbO9a2xY/qsMVuy8LDw8WGzgERSJqouRuyWjh55vzxwkgqd58k2KCljSd/kYcWQALE
HnABEmFRQL7Mm+9ELXqmSHnWJvYXVAGunyjMexe0etYAe0QtdiLf2J0rWfMmZXFE5zrwn2vnyNe6
r9jezViumlTZuIzhBjy2atvAhk790D7hWXEtXszhFEQX91q+JB7uPCX8tUGHwPC6xqRrfwxuuMG0
mpwpn8V4pAuq/iE6axTt6oZzhf8ph2kp+4MN2i1gtntTFj9sazY/0Nt6/re2fqNJH3uKa7OJLWfx
Wm277THfQAwe/GhJx0WGFSH50eC8yyL1XCeLLBULmymRhbPv+tKaQofawlDdzJTJmWo8jxExCW0H
9JLXc43RrGW1wLzh9bW9nx3s/qoDlCoYhoHgT8JvBx+szgSfRtnRaIuF1rsTpvEZ8yVvtP3EGm37
0Y0V+x28b3gTNpr3xmrK2PDbHOsg1+5x1ivO6MIZaw1/a/xW2zDYSuX0FEoYqz+ySAA5olszHxPd
eN+RygrzQzxPvFSvH9x2XV8wMA+Er9LvwXWsH/OkFp8jhdxavwA8S8Ii9sDnuR+hg6s1SMn5BbM3
UuETrdDPCBVGojX+jghKDwfLqpZxLU7G3IkzHflLtR87OU4NbuSJOu2Og5E9dRneK3FAU8hlUeqT
QYS06g3CMrSzD0p5zmZf2QiBa6xA42qaO+NYgLonb8l5QfkKc2NVGcNuM7hv62E0XrwnVrI+Ilbr
XpSN3gt4LG+kLAK+1ntebesGkYEG6vG+75e9FCJRuxgi5ftYx4Qqrd7WE5KzsJ9nrvSDWsNU4Uh2
bBvkguOavRnuaDSXh79emQ0QUlgUcjN0xTxhrKaN4aVfGruAQsEYmHEMOwYHGWyz9I/kR18ukmbG
sYS/VaY3Jy4BdsW8Tatezz+RuRHnoWNsNvMtZAYMF/2Vtln1DTjcuzeFbgLOQmpX1HNFCflPNFzn
yV6oNrBJsFKCItvKZ/wOshvUlFNTSO2eBa21RuTMuKufM/6ri+rlYoRqoyV6Jv0BFj+l5Z/ZYNI5
KIe83jnmj/w2yPrcnanr4oVHjeFXQV02wLQDXLKY689WikCvcHyWuVfIkUlvuKLSFJhBNDQ2GSPH
CEIznF1tX6kRrq/M3Zvbm6mLN9LIiCI68ZZHbx2XIMPBmwPVpkatfBvY2inHQgs2qcVxtO6b0b+9
hOuFnsGLbHGmbBcUfwK6rUVizhAr93cB5XB1WluYqoI939qdhUz27QeJ7T/9S9EZz3grkWU7NZeA
NV00s7ZIgxzBav+O1i5ivx1CgVYKKTl+UxFHSTUIRFQMLOQh5qUzUd7qt+hHwE15n9wlzJGE5KCx
QIf4SWjUETtOC+gW2ItBqmqmfRKoJwa1jR/Z6PibRd731iiQp9kd56NaMMe/Qzwx6p6c82DzKsvD
mOPisTvPXUsFu6Dck3OYwWmQ+lcVa0+ajN0OHKnmCw+0RKbKD0NXK0GJ2ZTYfVddjKODF+hJJtvc
1XC1HmpC/6/qWTjf0feIYbhj0ybmvPZf8Kv/axzwls6MVkuaF88KmwuklxtY8ABL7wprNZpF13Ea
P7QaDsYQTi3mGpuoqBzmWkXNEehG+LlG1INtGyDINx5G6hfukJNRDXmHeOl2bI7s6LshL9E3UuC3
w0+Joa49ils6WB61AOOf/10gkRqM/sfSD8LL6Lqsb0+s5O9iDHVegmNziiULRkWysc2uH7jB5w+y
bBejxbCg4Z1hOD9WMzr6JV0tp81jD17uNYND5ZbbetaQ7iR4F9Hkly78736X5ru5eQieKKDjQTf9
0I8Jm6p23D0gEXdm27X7vvz/Z99dmcffcbvvbKV8Vw7lPAF0199wO7UIfZfA4xw2YChBIe9pw7oS
veWhvig9N20+iXEVF6djjUpqAFMPoz2CnM5CeE+ZZJpBoFiGrHtx/0p5aDT8GF1R/ReYE7GyMG2n
o61XOVsh/0mew1TZKaGvjv4A+OwpPgG8HBqzTlNVuMl8gWlHdBUp162PNVDhvQMBS4M7CLdwBX5V
QaY9OMP+z4QIboAZdqtvr58cwGuW4MLpVHI86j1YJ1l/1e1OycljkA+7FS+DbmzHLh0QguPBRjqM
T1oWSaH9fr4M9gcOHz8tfNkh6hxSuoNdhxxflDNeghZtMCJsEWLMnKv66JbG7U+qf+d2exHbiJBG
J1+K+jGNSGXx9QsRQ/Pbhao4Vv+H+XnqD2uDUTf83OEiZkyMsksoS/Yu8N591znnGRfHKVGvWFvu
i2MizU1/aqpd5+qu4RjJK0CmywIhsU4mL2nmOIaU3/5oSoSg4w7YNYDoRnCIjIVAeIpcC5UAvSEI
14GKK3Su2Rs5C3vYH49x7c4AZF6bv7VokMSoeDicBm8rtWe1BpcsvuTu7bB4lxIMGfdrn0A3xwE7
clbD04qP2WH8V+tCZImlT48jDnFOce3JHIP5P1qJH3A0uXZMK4zfyy3xxm+QAdSVWgNAJZOJ9+/i
CZlDG7MhbEjLvpWwO1DmFv4IwdAAo+8gOIz1dHK2UHo2YKCZcO7RIUpAH4wqSVxZHJSw9VPFR3Q0
3cpOkGHs/81VymGcjTn1nrWqPNi8FQQzHmxnX4Ns2p5abZ0HnzJqiJZ1HgPS/RA/acWkJUYn0xQF
QiRrQgQ4y2GIsPTAeCPC30PqCH7PrPwNYYAXfPnGgKEtdkTppsmDmFF5i+wwBjaeerQhp31sHetI
+Q2D4ZRHehNzpYmJKUvFguiJDsKxfyPFY0FijLWETsDiQ5fAsKAhAc4TFb9WSPq0X3Gc5l0nxWyp
9Nj/PT3oU4FW/RfoI5oONHqNceodMfG5QtsyQFHbw8YemsTOZO0gNPxUf4GbIpjdQx0niaxnhzcM
BLO1fNItz5MRyFuAc4TyRq1e3NWi9xYnrKQZ2lDdOM+ixVF9aSWdYsapr0IQ+fU1K1mWuGZYbs7G
OPulJFdBvERm859TTtxZIRSTWM5rNWYxCtWw06mFdFV4zhtdFqOrf89+1UR/Pqbwf0xoOi750NYF
aKeKymr6S8z6kpsYO67Is7pudGMvPpQbpauFcmxFXsekJDnCistqm9VieubVCPbWT6SDW04dmtjy
5F+Conoz28C8YcaIEEw2d99btntgOulK2rCBLpnhw6m8bvQE1vyD19Zy93xB1trG/YMAEuTKTSB5
gB4f5s/1kV1fUpQVMKNbE8sqx9lNhvXtOkPm6qBAtwQFmCp6Gt/MHyBXDbLyG/Wp2O79Tivtt8ff
O5lODtffofzF6CX4RjcOMmTawjeUlWL9HCDsrUD+3273Fog4MalvzAr2xdHM/avwZ6I+zVNU2Lin
Y/xjx2O5F7JAob1yQmiHpVKPOIkRJpN4LGIrpcfiJrVXlXnRCjumLwBxUA+hCL+CL72sUJKIjZ7X
L2qENO2/1n02H8TLDor+D+7D59GAHTBTc6zxNDO4XfIgPuJruHyZ/R4PRXqZMNvxfa5A6ufmhfU8
v+Vmd8Fw0w9y9Rymrp/T+Rn+JVYRQ0Wpk3liVMdWQExOiviLc7yy2r0+sarSTNLTKLBeJ6DWtowV
WTEeASZpgyfKOpcy7bFl806bvCYU8Dix/wDErP9EEFm8nNDqdVL9fJ01+oZBHkUgyJI82Y10GAWO
E7B7Ge0buIQjkzq+fP9D5bwr09FYoZm5oZOb0SqG7oMrNcwwhcO73PDF+kh/O0eRWZuKYHh3WkvO
Hd9HuhqnotHdalYrXkpjMoFUNfbNrs3jsPu696QQcsQDVpS0O+Bn1Az+jBWmlHmxb9WxLCPd/q8+
0WXrKUAJZ2wEWJahepLBAto8j4/eP4KNMqC+SAsug7UQrUxtvKiyonRepdWMwSA1M28sI3+9OnqB
YyQAFv9bNiRCBZXa19qr0otisBG76Acxgp297M0iS1oH65JbzJPXPiR0QUYYaWUzOEu2TJprKrni
PpYoBWk78xXEyeQAy2Mj3yQid254Oz6naujBTpaSkwQnpZ7TdBtOPnAjZwdh8yqY0W47CGCjf5Ij
HFi1CDJ1ERUZeqtoIrE7kwIArTrywchec7flFAWEOEIq4ny1qVuY6A4s/LLtUhxN0rap/hpUAlgk
x+XD08Pr9vKOH2gjND0ejXy6Bme8iuTdtHP2l0DviVPTQkZU9tIkUeY3x8Og8PKltmYui67CPaML
OmAkGrrbcaSmWqsGUNBYVB5N2v/vA0OqyiL9QA+1mBP+tTlzapMwYtgmSsawZfIfFlbq++d3unXi
HLcNUD6kiWtCtzm3LzyfEUpIa1NNe3kr4mvdKVNq1sMYSaq8ILI1jfYuJhp/WjMdV+48xZ4fQ6hY
hhE+S8ffMDiysv8JoQSyQf+oF9AAprkrhWo+e9stkWQmNAD4bZOKZpYO5IhWmRUZe0fcJoDOp4lU
EeVNtIW8HinxQ+LlKTCnNJ75Gp1Py+9k5atI64RwN8xF0+RR0GUcVdQaRba8/TJGuLrFhBK9pBrY
ZOS7Jt1WlsTPZXL4F6LmXWACUSxaQ+9kgXjDHdC1sbGwXAwPrg/ctL0bTMtfBj5DY7p8trt4qES0
K1P9Ya1aFp4GHNpWFIaTF5efxuZVMr1D8ayFKc3/24z3MPc9fiO9tWo4PTL6F1++9k7Gpo0BSJ8t
MA+8ASS9mW3HUOe/lHtnNXp9KU9aVk3kYxf63oiOCMvqYsHTZAGwsA6H4hLCx9Jlx4KVkcVpo5cN
C79DXKBR0A+n86o/gAL4HS1rAOfvO+p0A7LzKWDu6y7UJx9VsGUnO/dLfTZeDWYZeJzoXGq7VsQk
TExH8SQysHJ5YVBENfkqO9sN5GFYgPdjdQHp9zyzWEHDraOr62kJPJcwSY2otFkDzUUhv0hRgQ1V
v4SdNK9CX6WzenLchm4XRklEiz2li3KwT5z5IOwtEvBnhMEz1JdsaYgJ4FzQQaiG79SL6vD0HdDu
HVp/I6ApY/dDEPk6VcFqcli7eQmNJk7K3XRKdHxXfJthNwSqJxAYsVMpE8MJkoB9AEjbUdDNbGk/
HhAE18vITZLpT9egA8wsE7ZqRNberg1ShxHSF1UBiFctiY3BEQNP6inRgb1pbDh5O9IQ0M+5hw3u
GqJZhEhC1QaRqsVTlpkouvxrAouAThr0T/Dbt2YRAor1g/a+QCwAxVxv+dAoUCyNscelIvo97Bnh
WnuJ5vX3Ejk2EdEcSpdjIfrZGAhhWqbQQV8vXhsGh/elO6vMbXCN4FCQGbK35/LrGTtXWIDBUJYS
uI+OaCzacTzqkU8ZnCZleiT/Vf1+XJYc80ysiwuYbK4rg7B4kao4eF7rDnqkH/YVez2XiF1M9YLi
MRqlgZntWiqtlV0fMRJb7eHFKP9DMPtaNNKJQMRkcsqr1L4rBFMVccOxpQK19CyLiye7n16wtLSg
N7lAC27o1QCyi/eI8iDCNc/aZsZrBxyB1YN2Zx/E+uO1i5O/Jvq6KpdSYxKBfSE6GQ22Tul9y+cl
7SVZsur6Zos1pZ1yiHkJ3FgW8iK1GazOEOTwPKnpQGkYpnP46qmT2H2psGYljgoBFPPpBc1RKxJ5
dQvHvoIiDCY3o8n43Oog/pl7EjofWP/+ZZB8KMNnKrFGaumtpgV9s6FI5XAKUeR76Wi6UDDFmVjH
G+030MaGJyt60OvlYcdewQrsNddMacrclz+WK/UejlUscuwCjImy1dCx9ar2AnoemRd07wn+5Zsm
xJfHB245998JIPwwi7tVZR2J2UDtWdx9mURGNS3lfWRaWj7QedqudjjNdRX7PiFletBBLWYXuv6Q
8LgZxEjCG89+VMnlS3IDrgFcLlE/btCprfMh0xu+jqHu6FtywNz+YrfkXWe/EyaCgLwVkPTBCHfY
QBB0kblvY5dfbCFMXgZJbi74UD00cpA0FT6RH4gxyzaPercB36HeAr7emji81+1SzI7A+Ee+wUkt
Qy84zydPLptvxwUXujuNc4DM28H66iJRUSLc9mvw6h3Y0AwMfypWDM3f2P6qR69fu48ofrTuSgud
24+a/5m5Y36HwT6cryxmawlxV1B1/bI0MWYmKxqRz7wc9ZuLPq/b4QUS/BaNTZO0vRpE5gw/BKOC
ZJsK5eGw7ARE1T1PnX3b0/u7cUHhrowqXPtSAwOkBnyZcLJY4/JdZ8IbRK4/S8kgvVrajCult+v5
3z9c3KO28OSNamFjuN2MnrcRnr6QVNqX0x1alVKc7zcM9glMB1VWKBvgmhVp7/pz2xz2wXYu0Gz2
baGLGIiwHek0zSZWfdfAKUVCQHFBGnUmHp0VmDgZpHSm51w8yeFttLNVwoz2agveWieiOPVlrxgN
vm4cf4qKOugwixtAVA5HcWdCcdqV6GaLElXEX06V6vHwOyAr7HDjKpOKLNO7pQq6G1L2bfC7KoyI
B4H1H3bDh8nqJbeyWJETCC1eQpWAdBprSONvWimEPhlW9zMOsBjllfJkG6BWM1OsOgUpytQ7cMlf
pxR3y/P6kB4ZKs6uFvfVa8QlFERyBXm7sBpVj9f2ddMhLcVgKp01IFRVpqWlpxqWan3Cg+dw6jNG
xePHuRkvilYndrNhuP2B5I03BN4GYJBqhPYCj8KTG6/goHjgtGktOXn00DDvQaFYfwbtzOqLM7oi
NL2qPz5QuRrhauUMTHYCb83gFyI5+Mb2+Y3bDgp3t+rtWLGVDSvaTBCLR1Jvfv3lOR3UNI3ogo+z
vAajVGzCerkedti7740YfDhAu+zMlxnTe8u7YWuG4EIKi0vot2113HuHtrVYy7Zjd0ySDbJgUOoF
VaRIh0nLe7r5XBQv9T0cYK/7lI8yuEEMFQwJdBO+ug/EIcY6Zsv8uhnS/c3kOf1+d3ouvK8v63Lt
P1h0/1ncsB8UIeBGsEDQjzN9BID3/8zX1MXONl8uGqNPCn/jG1Vt907RrMC3D/jL6YEgwvsfmnHS
+FCpxhotVSs4lfBDpe3YFRbYdbndie3KsQzGBL7APn5Bj1VGyBcY9lymTLXxwthRlUMVjpzbGp3M
Y4OjjiFRze6Snl6ZQ9ExvqVEvKeXiLO+ctJu0HYFqwlO8qSKQ7j0L79RHkd6qwa2iGN3BJegb5gy
lDbZSQGzMnLPEreZoAuTz6xngbrbLFYWt27GTOtweJbSWB/ZMONdH/dXnhj6BGvSwNi0gMKr0Zjy
YyzoEVWFQSoZN3EPeSFXiCuXqw/W4aTVhgemLvvWjJjAKUL5DAz+xq3HvLuNwxCMzFWufWyGH4W0
X/IrUHvRZcVHsgtvPQeMI81r2wqQsraxm34eOz+ebnyYc0au+fGYIK8NlGGg4fBGwcuYqMBrUkPj
i7p9cf1u5biDg50pZ1sUxI6MLfkPv5pgoPhnE9yF7khKUZQRXiCuwSUEhAUDE+Res4XHjhynhMrt
DV2Mv5s4yamgUrtriyP9tcOhdK63AkVw48D2fdeGr9I0O2VSmc5ZUq3v2PnBxXM3a/NRlh35oWeO
3MSeei4JGa8O/Ry0dmukrbh1sx8Mur2B6OMxRBxg4p4g1yzvFqJ7YYDLwk+qSrgbbV5NT0uBH94y
hDD+YuOmRYX3H1aAUGF7k9P1bx2kPkTG7AocPpILhVNNcGU6s2vO0uNyu8K5NYD9/x6hkYpJT2ll
hX8AUgTGCfwrOVT0/HaoJ6+H14Tg8dXIFvy7NiHDGDfTfsgZnC4jySU6n+Yq9oCPrioljLs5u/c+
TwMSKwG39NIg+HxULLDJIxyBIACAxHrN34cOOQWEY6ZGkQc9mMzTh/g5tyuNiT3f3kbHo5spcx8K
Qd9eHLu4hLvxtDhYRA7KNmFauZuyN34V3uoUY4C+ff5Q3Jw1lt8WMHUC4sJqzGIrwsr3RyO6GI5F
q3WthT4m7+wvAxI05nJROTZs4QpITmycNf6I0B4+z3rYnnIUj5MUCTBsnQwfLwUJ7Fe6JfXFkhdO
T3Yy4UARh9gIF93HivmGCR+mCyKnjJfmyMATAIDIa93fiEXNxDGPQk1hTNE5NjhpKGK4pdZn6zvx
NU6KolDSoD+Pqqv6inSaxkFvuZSceiB24Lfavv/mJwS97qjigpBtHuQrxqUHRZUctofY48yYC3hU
yBifcr56zjl8Z7cd+Nxk4hkAHMrd+UgCTjFKZ6mitHnFhOKnW0tK1Po+AIwIEVCZVtUROjKwhPy9
sZbb4tR67lfZ/kMJ7rOIuF76fyr7IO7i65b5latPyBLTUdZz8eTsp4trCxWblIK0b4CmCKtCkr44
QcdVEi13hefHC1kLJxm+BRqX6sgPl9BkP5UvYJ8sKxdsW/VvyUqcMxeTQO9ekL2s4IsiHrclRuHD
cDsyzKXQ9VkxloChjzVNovVT5q3FJrACmVod/FCK7GsyRIfEmNRoTObuh+6TUziP0VOnsSLzLOPr
pYXYGj5YO0L91PRw2H1Whd+f68C94UiVeVsV4CbCoW35q6g4LIgQBLYVwEGXHOsDNFsLIzaQhrME
R4RpU1TB+JKxLyutvNJsSH5yKK0Zf7FHCRMJFthmIi/d9z6jj61h9nnpxrg32oKJuBP6QCzezZ2y
kYCgS6zpbSt2D1R1EygXWaTYka+chWeFe4suBA5btdsWb9qF0lYJMpjwLii5SZbVjgwBCa/NxlhF
dh40h4xgiOTgwmEkOLUMWeTz1dFcMtYkxMJDoOuriugH6Z3zot9cB1Dod813P45JcI2QkI3mC7HB
7XtcGVMtNdp53LmrgsvFfPA3I5DBpYR36J6I49wYQ3kBA9dcmcXBg9iwqseuhsL+bSML7Ndc7h/O
5O1UiIpeTPmWemtkhOGtai2Z/vfPGJI1S4pH3BDb2McqhRHMYOIxJ/fGM74Frl3RxWOY61O88K5m
g3s1KrmkGKOkHVDOzmau8cyrWw7RYcCkDKdi1GsP4d4ChMQbiKEZ40sTQ0c8s90g5GJFEbuI1vkp
nbLnVb/9s6TFQ6qd5/9x98zi2W9jV4DJ6Zd9XX/G0EgxTCqHjt0L2iu7Xu7HefAsi5AEjPVPl+ak
5KJEKKloI89EuxU7EXcHTbQHJuNF+GOaFROTbEwE74TZ1RLRqINxMonO5fPq6xeNt2hBSJP5TOdB
qsOSMS5SMAjcMxF7HZDCUdV5YxeN25WwY2pZYU+dWssP0zbfqt+NDYOvJ2Rraqg6UH5KCFQkB3sh
FrOYz4D521k80jMwE7dARFmZa4Xv9fsQrPfqql8ULtqFVsJdJimT4PkgeFY1aNtbrxWXYgJSeawT
ZY3ZLuA+YZ/N27ecBI500LIOs2ajyah/tbIQBzCbGmcc5CcqZhNI9H08eo9A7d29QQxE9AZIaZ6X
xyRlYA1wYpJaB6UuiOU8Dz3qoPKaQO1XmxNn2N2iMX8XEh4ZCWePBBywDbcVkcApAWLIBL27TD4A
XhC6E5Lt/HYYrjxXYW9HEflw8usRJd5WeKF2/1mkWJmsB/AQDU4lNLYC4hkTRWABV+/SsdcIy9ig
wtW8YtxOeqhvab7YQSb6aokzX/ubWFlYq8CYLuk4kDoG28H22HQExfdzSmatdSEp3kVznS2OuCSW
zsPLd8uXX9f3Z8nD3WWxHmq5I6eHNf6GSqQpZsrCvmtbMMMOm6yRYILTFzPXx8xZn0X4SKh/fgSa
ZG8j3zmUB2Q+01v8LvOESh+c12X/Lg4IlJJiO928LaxQWMK77egUPqHEEhaHWKv7tix/DdI3f/t3
9lLHPisADu+xj3e5ZJ3/uO5AMMnyC8XUHSeOFb5e3uDRYyZgEbYLl5UtmfxGP91kML3FY3JsUUkD
5fTAi7bw6SRDZPjaZBjRTTlZt+yFSsetPRyiw4HWxyutF7qAoVj6+YYwyjZeOpukvwDLCJN+95kP
7v2zkobOo46MhbSOzoXlTA7YVXqlfle3jKrgw06MD4ubIxp67cqm1MygiwxiMW/RhpVf+YPaSS/7
bw6CfMXttTdK0X7cWdCIM4njVotii8V3RVUWbz1a++LkqKv2bfZGO0dXEpiNjnkH7k4SZMw7JcsC
XGdy2dJRuiLsxVANLBKcbbdsy9cEehAiWcUAhw9ePelSSKP6yDRLs+lGys9DU6rgqPyt+fEdKM5Y
vTgCXTZHjBH17Cyh6H0pMDJc9KEG0/WXeARqV8g8YGqD7fZfPQqeLvFHsw93LwOfISN6njvfaN+9
33KH4JrrNdkSKuJbKl0Nh0PDB74rmaKFZ1qix139FtUGp6dRzgAGh8IDvciBHny0Jgsmz60OJf2+
dIjfYZo4f+xhFo77z9ghKDxNedK1XGGRXbVuGtEBNtLFwIZuJ6X8LrtoyAwWEuiNMIEP95z1EH8o
NeGWAB5Wxm5Mzn4oiMI9IKeltWNXrBl/mpt+EuTWBPdfeHQenmYUNy4U4TRD2ofG4uClyBhdpCaJ
6QijLoIHiCUA1cjuIjMNQBEjOdd/K2oUxVd/Hg3JTxk/HUKG+4E5a/IdzjawruQZL66zbwI/rQAE
KeBAXQkE2lR9mw0o8r3EB9I40zBtr0EZEDqHI6RbQLMr1C32VML/xGyxd6dtV7CtHLPCFNz9PmlJ
Q1ZxyiRk36r34eU9KgD61xhCCSm0XpcHZzXRSbl5BX15r/Tg7FB7siM1D0+vnyddQcK8y8f4xzsB
jYFtPTT4tqUpl+be5h2I2vzPrrTm7I0sYGAsURz8OegC06LEUvty5IuH9f8zSzhMUGy7PPSTlOZ7
KE3qLdzRj5f3PEmJZ30W32YwTdjHxiaREyVRUtQhrEjsRoQKBTkLucmx+TiHcQYgoNCXBHWsvXgB
neQtuivE02u07BLff9LFpKFR3BzjE2TCL//FQXFUZ+ILi0LQsvZTAWsLHg8YmV699KYyssxNNkyS
9TrGi67RrAuH0y7Ut7aZWD5QQsI85ue9lEF2VA6GBDgYjX1Gs2iFweithV75NSxkW9StZlpmA6+I
4I3LNCM6T/Lkoa2olULXkZIEvS8iNhROphap1nhRJRKaBmhEtvarK3mXEddm6eQZ/LAsRPhQQs/G
aqmb5Sob2jNaBnCXeJj5tA1Am5+lhce44mnjLCdI42/QTxSQyLRlCA4o1GB6D9jfwTjBEhUarT+z
+OhVV3Au9wcX8YjzjrKDlbGEclchgNeIiounOaMLWMVCDLmJ5FXsyM94P6qYso7rnEX2CJcRcL4J
iLiOvnso973CbL9fsi32kxWi6Laa2zaHd5OK2rftrGYtObeeay/i0bis3Abavng/bevBDDeWoCko
+oBiOWUtQHbCqxptnofheQukxwBlb76Z0fk5UfbSo3ZA2gWXBClUPKiKSsiYFF6QJq3kUTmcbOv8
nk4OwM3vjJYlXolqVE/c3UQXVKHhC/MRpn3rgn33RAEQHxDdJx3SB+loZzBqTWs1Vm/qRFFSaZ5C
zddD1DYoqAdEVyKTTLVyjinwJepGNAeUowywps9oqo3S1Lg642F71pQUA5X43fBGAfFLmsuT2/P2
PSNJWKdPV/BVd1vNj7QyoR4bT1+CDDh9W0SljZUu7SuHHwwktlhH1GHmHbEd3iGshMsC2wO+C6zl
mD3BaPcUQoPtqyi69h2PklVSwxjXn5j48RBD2jlGi0f29Kw+9CrDr2NfIjq0V3a4jMsDf/ag/wsQ
pnRnDJ16h6w71aqz27tOXq4NEiQ6TLbKhm33xXOA4kavqz8MoIQXGWd6pESGkd5P8bUQCasxe2xz
Ks50cw1Ma0mH07jYo9rDcscPC8wZ9dWHRnnryyLyWkzzr8GULGcYEtt6LlDs7DmufHUZdf6zxnRF
AuMql/FYODIAhBfnwh8xoonWyKw4b5FHCbJINmSkgpjDlHc5kAbfCwlbgsGVKomiXfwokugly9uZ
c+ETWZCKJEvnnQQS4I5EzYIo6Y3R9S70cyP7SShXDrNQNNo6EEkzW1RTdR5N9SRuRP4P14CL9qro
bdh45yWFBZN6AxNTptuF7g1FDDQv3azh+veVP2p69N2uGzN3blJ+QzlCAtDDaBqH+IpnzpInISI2
5bmzKaP5lb4/JEQ9kCw/Be0i+OMbGCbtFvVTBDzsmeBt9iZX/v1hw28cbwkVSVNmZcjtiUxppnyG
SPpQN+APpzEQ0TME+fFMijAnEv7mROk+5WWri+pO3d73PI0N9KcmmjysrRetkQVx0eC8tY773Se6
2txa1+q4Ws8JjEUl5qi2TkGzNJYjJSxJygfoNnQx82GbFsTWhpw/nOo0hx2T2QcNnnyjV2BIqhJE
D0AHkkG1/87pOVvAEkoR6rEkteE4nlf7/aZp/PKhArWKXMw/AK+ywXB3WfJT2xufZhVNLtsR3aSF
TRLzrCHEM57BqlgqOdxxABJXdJ/VnVshlkB4F5Zzw4BnWf1FRvJdmeUvCEfzrYMVZYHjzCrf/53k
fFMHfbx0oc+gYDb6uFhEzjHJy/XQHdjfTxeztaCa4QIPFr7mBcvvY6YXSSj4irZRQaFvSE/uIITn
pYFteZwRxywZHioMoSRROw4B6nSKrhROOVliZwqMMPV2Fj19AyYpmRS39yhjt5QoxEz4YxqI4en+
3p8ArUVZx030Xu/VxTW0J/CQtAnXJEgp2JHBzm/V85EuDObT/J7eKlvB3HLZC1jcCYRKq6aAGKa1
xx7giN7BXEIzfIxbkXCay83n6m/xWWn+sk45EIKPIU94Hm3kz9IVtEFQ4xBvKDIhGObI+lI+WIUa
2K6wn8UqtKK7DB5D3K8KxSkMCkTY+/+Adp82TtBoucgEC4se5UXMsI5/l3ElT4wREJCPeODU2PXs
pardFwBsMixN/oeTTvHFiulzBatmQmCeSVKEPdWedWjdk8IIATu+1k82elNaWqf+spqL2KR8FfBf
EUqFqOWQ1Mt7sFB/HgUFqu5EigPHDyxAN5zhjn4TDDS5Bd8MOdCaMTEx5gJEpWJdU+fZdre79r8i
3GXSSMGItRqch5wHMMS85qDmr7Mwt+SYFosye/KRKQTVuoH0l/XpsvvcU4sVP5rKdOTdmuHP0Of5
DvlzAm80BVO+Axv5hHcZdk4jBWPmCkCMy5zn8I5dGPlV0y/Wwjj3QuMsVEoNMT/T1XAQFAvB89cQ
RRBrwMnDiO3IDuMD7OILxmA+ffZFT/T0MPZ3pj5ZmiUybt3BHOWh283gGuokZJOiZyGwXX1g+WJJ
ZLfpnLelQHbhrjregDabl5L80P7r2Ik7dSNZoJrXUrDTj32arrISFSrCjnK4IsrZlKfnIuez1u68
LZ4CJvlXQZ4UyQuVKdBbUYfPOsWOo+HelLYjho1f9GIM+Rb+ndOLN3RYx7BBYPn1z8UHf2esE/yR
YRP2UedhrAbSL6h6+RghWwUrJabZ9dn2l6YbP6u1Wjap1XXueUZ4NMsaAv5tMkjX8CWhGWcGmj31
+JSqB8H/9lGbD9hB2GeWh/1aPd3y1fy1OWbRjoHo2/3VaNsU72Xmbu4mtwSt6/nvELrjHgundfbP
aaKNQI+M0HPCVOTc7OP/v+Z+9I6m7cmt5Z9TyUTMYgzpPTdPRTTC6AGsoLYoViAK+PXntVMy5mEX
SMIB8evYUutiCgwWMFJ0YPGUdayprr8GMrMN/uOlH/7cxSeu3Ff4JwGLog/vIpO2NQUsPehmkYzD
l67thRLLRaAh78j5F3LJMFaIjnmIMN7z+w6fGKWSkKrK9fdHAlX2ClzwxrP3RezZrSkS5NSlNuLI
ynS6J/e9+QJq1y0K395n2Ba/VgoUSk0pM56sHqVnEjCCzpI8W7BtSfmQN8hmoWPqCubmq6mw6MBj
eCd2DRBrVw5Z0LbawKbz7cLOJBhjqBori+X1x9NBOsqpR4/D3mNjROcxt21Nb6lnsKbo4FdGT6Sb
IH2Tnc7ObwsM21wgRs2tGitFl8E94kX+2kGLl8Xegkxz+vg+Ud4fGiEjWfhEYxTUVCa1+Vcrw/Vq
+xg5ihph1RrQUoIYKu53HEJcAmdaQxQCI5ZyGtJdbAvjpf6HfHbzFIYF46J3LA/95Fx0vtZBZqju
sqmweHCxtjBrGIFZ5TQWTUBQwGuV8O81DPSBUp4UVCsaHu9paS5QQFPS8xsvOTHqN8PRDufOMesG
mHD9KSTwZ7DgTSrbTrhUdBWv5PaoGdkF2nxLUoNmWpmDrVk19QjHZOAPWo8etiaI4hzOJ3msbXpN
zqN68fRVOtl92yezfuNsmQgpjFCfC44XgWWSZSDP3kNKJX0nY60G1kS8npyPODpYDAyTTlJilx5v
wfjp7l3+LJM8n5qDCV3xmGQ+T+6rskuyHOY0y3NqVZ0rHBTNeLSIOQyoTGE8BPPr8uLJd0HrFRu2
DOmhgN3Rf3AUxjtHowW/H8PC1+CSC7sqFA8UMDH3kHWNow2k2DkpL5Ka1qPPF6ejX7JTtAmatXcB
vAuU41ZBysObHY23xBRhpHVLsRyXD7HL60WesB3NDH5deUjhmBZ7Qjn3Yr4MBqlDgU0IzNGyLToW
e0I/en7plsgjDFq/O5QGqy2f+tBftq84HS/O1U8gMtQJ//R8AjMRZ2ZccgLO/CG5SPPe9zocNbvv
h9SAM64gaqA6T9uCfrM7uwmahDDcdB4RlWc+31iYvtcgfasZ8I+on67Nq7mSgL375t8+DX2R34jc
fcRWU2Lwhx4cL8RHlfM1nqlpfo4/1W+Gs8qcFeZsNdMSqjm9VfDobUFYIhbtEFAXN5uIILiS+Np2
uDxO5Onp3lJcFkV/PkuLvG8v48/zJxj7Ktbwq6fsAJJP+fwBRmXMGNNPONtdDU/11aoZpcNhrqCp
o2qp/FaRGPfIilDU2Fij6udfSIThgv+65dTI93IfmUwrjirKxQnXZ2qGdwHRpqkO3ooRwPpkC/LK
gGim1UPKh130YSt+6fej39rVJPLclzG0XXRhupeuMUnuzoRq7p9Ij0QsVz8drZch8k3dZE+3U5vL
f2tWv3glMpxnHd/kAaLESDxWYhn4CmN7Hp1E2KYmYxcqFMvsM0Lw0FoRmWuf702nT7Oj0/Cj9tHn
kQ7UhsfBRl9GxcQ4I2rYGSVcJdhAeFPtM1C+7AXYqxlYzWHcS9J+JdjZ6Ln9NvkgtROeh6wprFFu
m8mw25becQm9uMhH6NidDC8BIUIOfYcK7jbAe1zui8r+wVPsDOpH4nnZ2EqfotzDCHQ3UXWsy+HW
M+5kdvL4x4m3ft2uadU2+T/tes+LQozOeojCCzG3oRNrabI7iGaD/8Gxp7+jm9sTXfkNJ4HFHG0r
vuERhY8gY+Ks7rjjdRUzfM1NXtLhGTvtoC7R9BC9mcXtjworAgWltM8C6uBgnD0Ppdrx6PuKKVK4
AjI9cTzAr/6Blz4IGHaXevTYeT+KI/Cbjtlau5MjPORLBFjrsAQKA2j7SkFO7yCe0iP7eMUjCrYs
LDwv+A70aNAC6WYw/V5sE7OS+mv8o0px41vUWbyowb1HrfH2DM4w43QU6g9qIG5c+xRo/9IIwQg+
LEeHtRA2H+dSX/U5gNeaO/UvO1zSq9Ws+XmmTgm5qELer2OhXZu/LMcsCQUYNoQ1Sb863sueC1Sq
BCv6raKyT5jxUQoyMbAs9yJh+LHRZULmN69kDsOtqAY5Ucp3KANzGW1+TXAojEJM+Cjs7LnrkKwJ
2mhqF07ddwQLDMDG7dZi8c85MGjqLUBQZqz/pLoDRM7t8vYTsOCCNoBWvnrCwzioZR64enYpPeNM
RfyYeyMw+oFsQPaOq0qN12v0d7kwQuRBvT0zIZMIiu4LxJ7JIQrE8RN1sAEjllWtJrNAspXjtHtF
rpY30831U4YkJcRdPCkCEPVlPzWLRPx8j4PAyeT9cNtueFf5JhUZiNAeDg/k6i5R6ysGxCKh412z
7j5tTJoQM5SCOpwJBMF8MT+GhAFKfkB0YT48KOQBFOLeVTnPPAJijE1idtEU8aPxXf7CzofeOnBT
YgMpdBkCVWTGnRexBzO8L0rpSJk13MuVmhv4T1q8rrR72s9dXt1jt/nXRGKeE7j8CdhwdirXUbNu
6Yrk9JzyIk6WYXgVH3kBu0svXaLIyg3bPQHUh0gQrbMgIKTdevtYWKceza9ohRxtUa9qLz6iG9he
lHz05MS8Ugu+mwtV2/uLLO9AgaN9EmP2LUKmfVB223BqmFRtW4jDEB14rpF2+U4u7hzjH5/JchX3
xM+sqOmoGtHArsB8nfuMNvSW2/MiEGDiNWEJt8fOvOqyzR62MYcL9TAWSKw84vlDj6csHhnRziyd
hSAHYA3BVdCSkBymmeo5Sr+v1BxTxIY2KWW3nRPiYSIYdHDssr3oJ8kpX66VweKIdRknKFqr+5dn
QH6OydlHZ/UMHIUQEC79DLx5jrFPnzDMaY2zBPWtXAADKFKBMK+9s9djT2x7XNPxgcOqDMVXBP5U
+QVP54MOU2R5JOmDEnDdgLTblwgk4XDRh4bYT3CDQ2xC6CUk+Dyow40nJ3+iWWtqqEvHeAG6m2VK
8YUKd2yPjBZJ2wC9+TG1YXZxUB8g1YaPdkCg9BkCIisIL7UbxehvEg/nFJPrK4++c5PBz9dwPh4e
cAeFXIvQL++wKpshDYRn6PFWEH93Hcm4EPwGrlNdWT9el6Nld1UQCsArS5g2J/I0TqxY3Zk7zw6L
ZVsRUGcIrrwEbChfKAkaTlfKERPcz/jrvmCiv8RDvR4NX3QppwRgRjLm3P4lPqVWZnLRhAd2mlPQ
lW1Y8EzVcePYdkT6/S6wCUsJedPI7PRHgWMigUTxnypOOnGVX9X7PaNPL918ObudXbxptlrCq0+L
2VqPM1EenoS1vxV3aVF0RCI1FtzIYDEoYnMievKi5lhK25CQEaZ1r6wBFExdgGtck1zEiaf+/KkS
XuqwbC9HBKVkybWN6aVVkjxJ/LBYelGZq38dqRYPycV0UGJB32mZJ4JqO+cFCUQExhHHyPvi9hvl
jOanmRPiNI42mTEuACs5AHMzljQtWiNAD3IAqDFWZE5OazW/k7w6E8/sbNsimTSnyGzMoqJXYyrq
SzRs7JW1JhTfCVtpbReGvnxrgP+VNAvyj9bqKAAT53XCNPEsJKfLVtSSrwsv86dTDjwnjPLXxIir
VH0V0ygDsdD0LS03ztBIyjw/yOyF9lteLxC4ynAYLEuDZlHza92lWh1kr0gbuN+5OJDIFJ2HB/VJ
D4aY/k5VRDUVvwONsBx+uVwt/xg9did9A+AkyI6nBI3YfEkOl1wQJ4pSTHWyk7jdlED7rkBu7sbW
2PomsMSVUx4xG+kloLAot+JhJdR5XK1/f076XBD9yeDiJA4JDHzc4Bp89Xu1k2IYSU6ArDQhzjks
RRyAxkAT85FfRVdAJcsyW4Lf38P5ak4BLGONmMO/PSkb3LRmgvo3uhyrzNUCMnwOqjRWKNZ0xOjg
67kY/sx10e/URE7D7D/fUSkB/wSBeEVQOziBHo0wXAB5/Uatm5xOLK6N4UU7AlEVJknadm9GSvby
p1SqLmRWoUxKHI6xtSFIYCU9vpSCjPJVYowQmbh1QJYT7YdFh37OmJVvijyGhgOulqHszajGY1oA
MrL+UitET2k2cJpknIUwBwT7fh2jwdlZaLblVraFU4UgUhtYBsOLLpTSWUhjuJjn8VhDDFCqsIL0
g3wb4JvJR1lAou5cmhEOL1pSM3i6hAU2vFPmcuLeQPcqbjgW+gGvIRGChq+oNZI8uIyCyO0+DGFU
Mx0Cfn/lQfja7Cm0wsbxv0Iz0RkVc+gzbRrmkpJ3v8LasFTHOB9Rwez1C+rWTmFcllGeu7KUQ4NZ
/MyClYUdjBX7zTNberj1rfAKzGS0uE2yg86L1qph9uP2qW5voCnHxZMDdr4Rif8s1u4VMcjIMA0F
BBz9OvNqwC1qBocGnmo+gAhA8Kc2C9wWo64+Hm9TAEHXKuegQkbz07gwsrPrBZcOH62kyQbNPKCo
TSaqaK9d1xMuXsWlvmqLQsWRASuNLQfRHult+D7BfropHT/y0ZY9+GukfQK91+hRPn0Xh+D5xZkA
/rWwr0qyEjcAiUdtaZte7/JLLY9uDyc0fdARSuZjtDniRcHHsJR+TX1pKZyYeRHwCgoBBB+Y+Ric
FK/UDw83G+05dsbgFk+gbHPH+e+3FZQJt41jO/E+salna2LzoY2SJ/WmYEM6N/dOw9EES303s0n+
Quufwn+X8Hv2Lh9Yszm7WPgW67xcIrLl/NoA2sk8EgoGzgmTcHM+J4tIJpzTlmoe1iaSFFF4lDsJ
Q14DmJ9T+4jAS4eOf2Ro2c2a2O4dPuq88nLCulWGH+V7ykipGEpUpIgRRcXb71Xjv5wh+erpA+bb
hjlixNfn5l9E6kyQCNnHLuXRXL4FFtDtB+AmezAvCNst7y6wkeknRyB4FDgbqyCOJ7bHLhIIHMlt
dPvOou2BSSGbRZmuo9X/uRL2Sw10eKaK+dnjUL+j5ie2ia68wSq3/wrWMBSh9esPiMVOOw3Fok2r
ifRiTWiHeMgVy436JWoWwKL6PDEzjEIpMQtXpF0SqexMBRhSfjrUrHZoWovcTUBtfIFu6EdjKHy+
iHk7jc1dm7xB+Gfyi/7Beq5J9E4151wSv9wdpcLaOA8KPf39VkLzD/w/pSMnmW28QyLxelNF0jLR
msJ8YM8QfdjJ8YLf2Oq1F7aHQgKV/Gw6a1s9WZEp1aRidlPsoOt1aghbI3M8zBF8XigmQWwLMsrF
gmsBX+Xb5y384GPhe/ifZvHl3TCoIOlQytV6tUoNeKAs/xKImnuygwMPdhREe179LIrnL4PFTsVJ
kYofDqXl3jjK5Pnu6PJtBQJcR7vaRJSsZJfscitwQifrNCzKWY8UTc7LeJ1I5yGWI+u4NyMnaBuH
hNhX6xhSH4Zss2j2n5QuLXM8r87JXkF65SF2KxN7avvnIUziwQBTF6j3GL8Nrfc3gIC9NTWo8z4v
uVWk5DuxsLMPTploMT8YF+kIW2J2WvBQJZrlevIpdqgiX4SkKV8fx0D+uDW1W3wFmpyk12Ee5JKE
IuvpTHxl7vQY8lY0eUQ03vmsaEqhOII4PZsjdWKdzTy9nxWPZU7hsrQF6Ds3VAGXwegoS1Fh3C4Y
AJitD7bLnHSi7//6Z+kaAaxv3FPGJDjNlbbATi3OTvwUZbisx0HIiBrdE1kPjNMDF3RL9pj62wR7
LFgbzq6m3P/Ekketkzc1+iaz8AFQy0QcwxY5Oy4XoHz7gxvlIu6WRk73Kex9sD7meN7+aEbR9Ar3
fBTnZS2pUzTTQS/Lvym+x1TQJZzp7zGp97xTFohzSKiFyBbaMntLnVEnCnmfPUqgryUr+GvXMBEK
U6gyeCpBdIZzapg2Wj8dxHE16pYA9gf3Zlv+vEwYG71ONUbRHOT5Z+UHwIoD/7CJVijVNC2QRpBP
ENPd5bSvFfFaYSoRIlWGK1ZkOj+5kzkf9LaDVrX6wBHCDunBRpXljrzAhl172iZY5EAWz5OZuSB7
zZ77XbINixXw95Gf6QDOFNunqWnqn/G30aXT6trm6fQdg9DQ7EolhQOEhploxP0YJeIvx9wUx/5O
bdZ9f6qpyLVcT3qF71RGySQowMtt9UPWzTeEWbRx8e1ZpmWmpMpeUsSxlcH9f1gR8lxv7OMwem+Y
IL9Y3+1rYZJbKzZIPlNgO9eFgWfHmoTyeASkdDX9hVbFcx+icsrgieLitjXj70ljjoESr49xOm2r
Dt8Q0f7iQcuC9yjjkRceQf5urbtDltYp+1zBkPAOTYzbtbUeqO7xphaLjKnNmQg8GslmeYVvNsiD
vH7w8GcITo7STXGVlhGrwGApWOh8TblmwRGxvS0Xfw9MjcSILmMcuxCk+AcqkUQn1xFDvePgVU9U
ExQF/KXS3Dl9l8ekmQlsika1Odcu8Y0daozzF4H0cZzR+N5JRuBNjLmK59O5oCiTqByaLPos/R0Q
XSgJNMcvYTjLSzR/wu8Ci4najVFYSHubkkfO0SQ0T2TkEKgIjcYsuwENXM+lcT3qNQ8CYP5I84oL
PTyn1bJiK3FGRBk133R8HijytHZsQqm5lCBlA+SwzztuvXsFSVsdvpjH3CvnAX6VhsRYBDk7fk5a
GEt5zEiTabKjllRZVZ1Jsll0NjpqC3TY88qYfL0lHq4V9PJbUvaXgtImTwuazf64f9J3YGsM6wbX
2Of6pw1I0u6kVCYewuhKv+APLVCyDSlzgtCQL1s9P+AlkhMxGg9OY0emX0Ow98hFy9NaUVbrS7G6
3+mosd5zMwNXJsKup+QHMUW0cJ8l2d+HeKJlQ6sXl2+yIaq60k9hU0eIG9QKAIMK8DOSly6QPMCl
Dv46wwUtbNQJZq4SbyIDf/eYF4oblpX7eF1w/Y6zphpfAoh7JhpTVt3oVMpzo/9IbLadV53bL8e3
uwSCeefZ5mPC1NDmmURTGjd5a138cu0V8+ZoaGPODu13KFF03VJIxs3UVCkqJgmrdEanoAgveFmd
DzCzSYJ1n5ngqEgreXFmD1zSwg04p95ajLUZ2zQPiVgdLLiLjZmnY0DuJU3CTYPwGr3bzWij56F/
SOEeE3ZWVKB9Tw+aiJK42RK2+BNmHOL88NqtKBbnA4kgU1qcemDCEMVfOqQe0cZ5iRbJCaiz/Soy
sYbvGVDUcEbwxhV6Zd58Rgj+wHtOOp5iCeRD9KwswXY89p58AU0dX6R6LTobJoErEPyXYh6jJfHx
iuA+nyDZfd2UFhl82w5KM8NO/FVyovknMnAPk2fiIN73thoYKL3R2YUGl/XrytdeDel/fzUdI9nk
2M3mlEWrnbmrvJi1Ekz060TmXJD8LR9twoO1GHuYADEx4Lm0vKyaohq2dCmiQSzv7CFSLKiT+y8N
IRnswX2OOgXEN3IG6GcdT5SHqdoH9q9PGuDXbHfnqiqqWxklQwtbin5zWGeQg0K7uOroswe/JCzD
QXlWPWVPij67jKEXaI9OZWKpWUhoP29IQF+I2cAGkkar/JbYuwhH3ns6VCIbwPYH7+uSQTlF53Wd
E+zvR/ZuIdQHOsAy+GAgh/YHF3xf6W6S+fwfUrdzBMGTE4ksBsougy7ovrZxKBQWXq6iqiNCiJqL
gVH5eu+VB0BDBkdyLAztKVLWelXPyTW0jEfU6YjQpypr1XLe+QtE7nPNgEdiWQtBViEKzQgHOKMe
GA23EuvPyys3D+M//nE5gPKHGlL1OUKjPTcNqBoofc838taKQMEKKyIyddoQjuSbiVKIRdBHfatc
SGaIZ708qs04lyFUkQFbF9Jjh4PYRYU/7WCRyObToMrkoxbVCNhQhp7DOfrS4GwIJfYbfHo+e+z6
L8F1y3zTT2SLf9i88isPDCkDIIvp4nDUQNeC9iogSCwclnd63JepLsA/MjaYQU6O+oZN9tWXGEjP
vdHRQzSHI6R6jAd6J4/VTlYJKXUzGKf4W8igtA44joLiAfjmC8p2REP8vHJeEOOyynqvgLI32m3L
G5Hco73cTs0Qf/iU35qUrDu034+d3554jRdANi4E1smPsB5coEAoTCEsKm+X/aUWEI99xdzk2vgZ
PUYHT71cOC3+uwIEbyHCMqVPVeo76VOVmSTkQZgZmMcpd+EpRFVvVuCqfmBuvkgukP+w/hfZ/5nq
l1ua3fqihhtgvPf+6CQHsSc7EsS0C743fne51BUu5ErGwqg6FcChJo/aOLwK9wI/Y/sp3alqPCVK
j84VfKzWoIjkB6NdBQwZNWn6/aCouIggGK+pR0FFji5d0fq447MBdN5x9oWHZ6Ong4OjyYIoJAK/
TA6Kg3xSSlx336Y9YD1s/1WNFI05CBvvq7PKrO1lNGySNnbbEdUr4u1VdoIzqU5xVXjgvUv+V0Cr
W5k0mC0LmDI6EVE7wXb2iRGaFlmXSe9+q2mVYTvC4v0IfClEFgjsCp8zMgaBXuTL0bw93zGqRTdk
RWqWJdEhymPj9GySd8D9zW5+kjT4WYPmdi/LlWMx8+Fk9j+RVLkTWVq1r29oEj84vSnlN51GE3d6
1OOAQFnAI3dytq/A4QpA0WDSlVs8VfM4JzUOKNufvbwl9vb2+/lrva9VskbMVyKQ+78RModkaOPI
lwc0VF3ork0OrjYnAxm2w5WDAWfqHkC52w1yOMjrh7qUo4+5+UVRrIzk3/jxsxewwh0mQTlMSIgp
+SJ3+rIFpRbuIPifAIDo0RI9SkbS4LnkCDvWqas74xeqbBrvbFL+mcQhUGS0c7L7zAFskTBs+pg+
6wexf78bIAj5e/WmWG9vqxj/iR6+V+2eYyBIhqKJ2gEmNA5Ouf6SZzouJTQ+M2kEl2ZhtQbin7mo
73JMY9I6kgwPDt4SxbxkO1wd+4ku1btAjn6X9XRIBwV7B395hHw/rul5bffhwa7AptZM0FFiKmU9
DoFQJSk6KGKgs6d/DhGs6fZGR33Yma/WFnv0gTJ8/XzUU72OIU1TDu7QWymqcN1YAWIL3ohCOsyC
f/LxAT4K/5B63fG92WHYKkWC2WrHBwTx+zA3pYRvvZwB9evZN/AmF4CImt/OH05KISOCdRgo8H/+
KPBU0d5/U3EYrA00gl1DDtGOvEZKAqfI5A6zkpvvUSqLcWAlHMzVvZQrQMUXgwMhYdy9CKnsBd2s
1/pJnbQblrfjGh5N2fXJlvzPufq6/rUTRJ1Kb1dNN246iGJ37bTLJLmaakqVwtgURRqiHWDjN592
e9eXUyhMzk1p/Tl+/hIGsV/EfR+0bm960MQO63r0wq/nSrZ8iDew3VZF0c1iVLO4Wz60tWdeNgoZ
RC2OXEjRsnDL2MvYaln4ZGNx+nxVYK0NYVfkeLRbqx/NK/ntifBS0T3uiRCTu7U1Fea9J1+KfjId
uEBQDXfDs5RS6D3QC5SqEfBx0UM+Y4jzWweXFBNdFludRJPvC+CLxBCKKmyY4XRiieJ/lFVZDfSF
iMniec9pwM7K2SCmg5JRqfb8au4qnaQsPn5zt7V6vSrPiU+QEc6+V2yWHQ314OUNk/+Ks/P/WuDA
zL9f/6G313seohZdDrlxkdP0msZ1oHFhEuNfZnrjCOdtlesXm0fXG/rUvXFqrLLhzMCW8yn4IK2s
XwQuvNki7WonYGAip8uz9luIgqRCdBhgNXDH9VvfS7VAWEK6mqVmimw4BfBkmZtk9XiSSLkhkeyw
kZu+F4SiNUlBqcJHNXSWxeOrvBx0bqgcygT5bTFUApWIIAux6JN5Fb0C/3JlC5QDcYN+jMNIiwEW
32gJT2b0PwD46FivE7cLi9gDLttNA/MlN2Ck6od9fHlKqeS2/SWRv5NGgzDp9EhJ3F56CPPfSeBc
tVzY0Ae3r2L8tGXsuP6/Vceit+Z2jtg0BX2sPb+Xmei1eoTrGRBklmeIJnfIXVB+RVmWlIdJwH2v
XRkc
`pragma protect end_protected
