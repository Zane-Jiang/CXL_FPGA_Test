// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
thfGkL9O+Li/EfeN4E4FxY3pDWgK2KyLJNSB25GuwS+0UFQPx5ITpFsg21ko
fdj8gABjs5cUqFS2zNOV65fVktO44gb6w73zARg3OBFkbBNxAeZ68Ewf60rD
jMkqsRlobqutgxi7ytNUewPpvQffncRClva8FMTUqCf2YBrbjI6Q4qf49Irn
BXUanuZ/KilRwbXC+RkwIdLfYUZjZB887W89SMneomHLjDlQY89cG79H02Ol
3D0It4qa2hhn5jLDbByztwTH2cMFdOQigw0E04cu7Xyjjiu7s+wYPFl5ei6m
+fUsbhsY80X/RaxNMEZViMoXR4limFwVfgzx0WEEow==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SnQPL/Usg79WaPRARc9tDEan6TjVzo9Zy7URr4tvJ6dcKLZKDrhx7nwAqBG8
qNFCNfK/sAwLaPxTljphwrfP44XAuWVbPZi31PRRj/UZ+KzLcbD7aLTvHJqJ
2vcKGNeHaq32i/1cHk+bmaVBkxB1kLxDN4Czgu4LqdNCdokf74sNlRtm1Gu/
AeDPGoUoVmpqojhtwcNl5NHV6XobopHH+Z8CVMLzVttWiUFMx1rDKrbRCvU5
BiJtY2scszEqXv5SCfvnnvlRTKWCtUE2FxSBoYj959XalpA40KF0ekzpaa/S
RUdiVesE+d5tM+CBTUgKohHPPe8F9gQTbDEeIAIVgg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WUwYsOI2+uirH7WKaKuCQtadZBZroiow+Aj0hFLJCEKExWBVqibq5e0ejAm2
ODN3Tu7ER0ZbqJxefSJcI63ru/0mPhGd5Q9TXTJppBqppVPedn1+fRphMAJA
Cb4ThRWzXUqUVs3I3MVvsXcE9EgFzok+VwWAJi4EgQCZRLe4CD8ALD3QbkoR
DzhtlyOJW2mwsoBfPe8fGotvzKa7zShjv6EL9Lr39ZPBKKVKtS/Y38mzUa7d
m6HCBiTVS9GY8X1aEL7Miy+6yBsquFLrusTXCk/gxPfP6YXEi/rZYB5O1kSI
P+/XAkFxNGMLdVsHfFFtAqOA7GU2Lcsa7NrfydtBkw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PiivWy8M7TOUJ0c4o9dhc9UJinoNWXl1XB2yFNnZiHB0ZuinG1Aw3gYbKF57
3IQkVhaLujx35QTmCpSJl2pFR2JTXDmrsW+TAWpxVEChiUxBEIuHpOwKsD+F
sthHT18nR+HeInyzEQU996hN3BHxuNRzOCIFDkgXZdX0CezpFcs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gDztD0KybLMJ6U+5qbYMQarrOoT10Iq46nm4PVveU8fmd7lsc9cViiKRxSgA
0RLZH68PgD1JmzZ/SamX4gAQcvhJP+bFmBHGChPqy3nmGgAhCQm4ocL4+aJN
HcxhDDthdN2sEJDpzEhHxXm7QkzPknAwIMCY2oogy+CNz4Y1yY7MfuzYZyqO
JOSVoW/dXSIT7yANr/ydrj5uELPJ4OcsIHyLm/cLBOmCSaP7OUimj14Eot7o
Og1hhGs7uX64Nibc09sY+FxoGmAlNAMTlqx4jd3M2X+aD0dS/VNUQkyKlaVy
hOIXA3xJHpCoVXGzYL0riaUdHd91sxnxfn6k3sGWs4iYIJOotSSisAMG70W7
tvAfBzGAcGvQ6ChHsUMMKWo/0h1tC0iAvkJgrZAtAE/oG1JEjmaWZ4WbCWuK
BIS065aVhuud/8FCGvSTJTNETxGSe/sKEkzTZdj66aDNpA0cYjRWUW9IBjaf
q42NR+6Cblb1Ze+cr6QippM8iIie16lB


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iYWkJZNIBv6Q5CHagDkfZOGaVoOFK+z6A3YJfRXwDxtwed3Rwo4fCg291jHY
7alBfnKuLfaNPZsd3CrAeNoAo4L1Vev7R8YeQ1SUR4yhygceOzPUnnuY/jyl
5MJAyEtltsL3w2urkU6tIMnQ8jdrdQHrlx9F3o2sh4UKdzE7BIM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j/Fps81/L/OaxODBSAF8bKfx+e0GLXrsXo300obXXMY7wWwL1j5iK40NEeTp
L/jSeYTC3KsJ5YxfNzxhcsW6PeDoj/8mA8yn/BTKtHjQzdJnrk9X+NTyofys
KkMiq0o2SVWJNm6u4W33fje0PYu8XTPLu9pfU9iGzf2XhM8oOpg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1360)
`pragma protect data_block
AKUibchSV5Ff/WPKKSrhgL7RgihrnnUUqnkKrzT2gmmm6Zt9oGV+u1fPVBEx
FSzzCRMXNzZ51fsdlcl35k72n/ycBh2AxQQWrP2+ohxNHMDzTEUdW7azimnY
6YYnlraz4VS8VSKxprFaCm8zskwE6r8g761OHP2wUoeQuwBQRll47TxHDBUq
jRAfyl3NIQ48N/Mr28zdF1CkWjJGpFP9ImYces6RK4BSIqGew/NMBccJzeuM
WLKKkawoRQ5nqkHg4goszI5FmnbOy5454ZwBGV/QrrHzjqSrU2aA7Bf4LbnR
qVgUQeEaQgjIddfVvbDtwO31rq9WxAMqs5lFovZtwgHpjWNUP+XcmQZ8CbmN
l4fZBK7pk831qgoTbFgm4LLoPdero0gUkwo9Ghfd3XoDwI9s5e0spPr/7nD5
nrpWYwrPGpSL92v3lM0NLn7BVpV/X70ppOFii6JohWz6yEVxEKGJrZAyKuCa
9W2RuDAXz9CSYFibsZhzd1ckJD9xxmC2Hizxlg57jxhcUXwZt4JihdU24gGY
G2trzuCV0OTsyAsaumKVV/cF0xLYZJwfgSejTF092K8anGmgfWfcVZYN7Xvd
15N/V76dQGqpbj4nAWwDvZb+IjaJbi+iSzm4wMQKFupzIbO7lkNjOfaK8OSG
nU0hmH8OlYfGqEBH2ZPO/edgIMg+FlyIzLR1DGiVcX/J4wnsmpQXo4c8awjC
rtxjK1Z7S4e9HGDHmRE4NEpV4QpW5GOfN+o8+rJpSaA6W29uiIhL6h0mUMS4
iDDH5unndNYyfAWjMCvWzBi2YrGU4CfAAI/wQP7b7Wq6jvVnE0tXfTHt8CKM
YaEUmP+tGztkd6M17koDRm0W/R+sZO+BxDrTkpFA5eF7npJ+9wqWoZRdzIPq
pXsKBaKjwcTwDrS2DboGZmucYDmyhetu6+ibqX43o+h8AemcwTftWdKbSKCQ
yNOe1xzloqR4VqmwakzaKBu9KnbAIjxIA0lSiqdDNPXpqfj9wfki8E5bjQh2
HNUjqAClopVAByaq/JsaCUmxcI8onn0CmCmRd31gGQzMzC8KlCmXCQcwGqgN
u3S3F9QT6bkFZhc0TVzldv/qKD87rgEByZtZ4edY9tLtHINZZJFJJXKYWZH+
QJaIMbuxfDluUWEbcXzgMEIsxhZenW5r69g/4qa1/fURb0Pyuclwfy7hiyOt
d+n2NCjfulQdEqJzKewKdqem3Gw7Vl/nQbuvMxWr0mH+kcqVaouDLl4GVIgY
ZBsU/QAkJ3G82Ja99nLF4ua6UaAyVQy+gsMdljVgTRE05pJUBbM/OyQu2k8t
Ep1tnbAZOEPPLFWlsof5BkrJ46qLjIO42mNbzq5XgkhHD3KTkgedEu+ifNkQ
43xIin72Lay+r83CMnrcOzw0pja4HTpkV3hvlztdotcUVQa6dHbbJbubSyij
Fy3tBFO3dj3y3yV+4M7Nl2M1+RvCdzZs+bryUsiTXQ2XCB0b+Kt3BxB4jhB7
UjierM9p9rNEBf3E246CaJceOmydwtR46uTxwl5P/ALbZu3zl4nMZGB/MvkV
QSSCWz57ULjC0aqnlyhcYa6kOdgg0+azLi6JFapyCcMNKR2FVtm9fXb1lyGE
6NO+8sToeRxUf4U7755L4+0j7RJ/WCP6M3r7/4ulKe9r6a5a08+H/OFWIxAW
5nTScECnqvOH0hMsOmaCtIZfPTPAoljGwInbxFv9+7ewNbW2Pl93EbABpBnu
6UFbWJ8HdwHaOdrbDsn/OPOLAMA5PgPz0ulPax2R5hvBikvGojbxky0WfpvA
QVlZpNbBUn7Xww==

`pragma protect end_protected
