// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2QowO6ZfQumYa++FHGiD7wVEjqGbHrEZrFsbtV+FYRI9Do0KqZ4KXlt8Rn4k4QY0
eleIuLhOFBcoMkQE7utS1gD9NhTdxm0fHYj+782++b9qah5yKSi0v+oyGr2l0ly7
J/9B1glnF2RXHL0jYS9SpKOjr5EdK9/8+WeHHps5mRIsCiKiFtGfcQ==
//pragma protect end_key_block
//pragma protect digest_block
Df1lIzXg6bd/Zjpflrt7P30aGUQ=
//pragma protect end_digest_block
//pragma protect data_block
MGY3tQP1ix8hEIrx5+pyv7j7p1/aqrejhjo1W7RAratlE/GKTwiRFWGfvYhEKh/x
5rODp4LsrqEgSnAYmdRJ8EPq4EwF0TRA8aVCxYdIC/hKrg2kMlnIMhbcfYrqFJeK
tcv+1muwBaduXM8/BMpJKzToMSGkMFyGgtNDJ0FgNzgAtUH3N+H43qJgQGpym2AN
r4NLHXTKr6LycG8a/8gP1zndbo/sgMxWwkkh/mUW9SXSVUTkWv1ryuTEC4VvtdLu
1C6wCiB/GO8SAE0Csp6OjDpfBcuxEc6Q3vtE5MW+p8yb6fZmsV6DlGWHL+kH0Di3
SiuTaKboaTShJdl8bRkNvcl/blgDrvxOj2i72UdUqb46bME4UxBI4t7DB8lYulhx
EK3I6Lna/+rAYk1mIundUAzJ8tY4z7WheN37uOdRYWwgYM9N/Y+2ZN5xXmFnYIV8
qcMeZ12pJ2hL3CofAsMObsLBIB/3VpkazGP+arTCMEVnSrsUC7bLeU1/nBFZX4XC
LZRgAy9IRgGT4IfG6bDp/VqexFDMyIBvgAuWy2aCiyydGNvvhRXHHcgxp4sNEqku
ylGUlG79WLpvJ+M1n+tJyxOO0hPB+/G/ZkHeDaiLfrHv4ylJtTWvoXFlMFHmiLwB
Qj180jFncW/X1wfqjR/JWZR3dDQEB/TZGALbpxJV0rPI/xthNN3z/m5WDZMEf/x3
PAjPFuNb1LnCMgrpnU33OeeNTan722PDsLtkVzS5ddkJbLFdhjrXHS9z/ucsFxZG
n6UcNrYMoo9znfSBm7yJpL3Vc2f9DRPAPJyR3JEN3bOZo840lsIyS6W8zrXaYVOy
7f3NZbkdUiJuSTSBB98gvmXC0eAoqCci1QAw6GZpXtdtjdTgtryEgBFu3A76o1uy
F5DJL1iI97hN2QMPsRhBpyR228oyrrtHXBT3I6NOdFaHdx6AOWrOxIrNojxojiK8
g4uvMZEowZABWyYDLF+HGc+aL4+fSzlf3OyiiA4/57Lv7jO3FfYxVnBR738gvLZq
fwzpPs7Wx7KsU7S4OscPWbDGn2moL1dMKMLGiQkRHmm9vgCMFV0kO4uJkb6euvla
F2a57zq4b85zaeb1Wayjo3eZITqeJ6pxxPmIWpdGw3LKSbXi5sTwWxopr5dIGKCY
OmFBP/PE2F7EH80DLq6U2Pem9Cbz3WWuE/w71owpvwPWPA+CzEh5cxnqqwn1hQjc
NVzYyup4D0OjThWltNR0K/kXed3sIB0xv3i2MnsLmIodVmu7sEJAy9+XgHnoDYm8
PBOhfwOTLdfUFsgmUEZE6j6MSgRhIp+HNTeh4swUJt07R+9fO/vabnijaD5iWwm4
Y44Sqbd46kKlmS+3AILgu+PpT/d6V89X7VP7Ow8rUCdVfFB33otTwn+bSyaJ4fEv
7USAcOMu/ypejC+JjeY0EJvzs/4N6/2x63sdH17FeX3oNHT2XWt0STY+QpBazDVy
2/a4fiqCasH2azI0973iylcBwbTsDa/NNBDTPhgYzBd2KKHYccHeIojxqULtJx0Z
xu9E8ebKUJfyqtrCRnnozX3XNw3F6VIV5Lu7WTxqdMmaJ5YizMcZceznSddvlRIe
Rb9zPT6uHYvwgUP1wSd1zGD6DqmJtu8bKMjgA12FQkPdUHTKztZFO1sonxUwXJHn
6SwZ0jCkcI7rPf8N6Y8mA5ER2cuYV01+oPyPbcFMDBJH986JFax3XB5plpqkTEUl
mu4eL8W5FihwWj3Zm3SZItXWeZBZ86O9NacwUteaB6ocuvEO2fY1n4RxaaAMYXH+
RBkWKG/1UdJwSl8/s6g2clkOGt8DjTCqAALvovuK9PK/AWlqdXbTE/6kozl34O6Q
Qn38OAnjPCGGasEPsZMjrBV7M9nat/ea4z8fx3jmVk6lBml2fuac8ygEAIoyaXpP
+lg1dqX/+a+1feyubkcCeTXEc6X6qPhzbA3EP2bLR+nAfouVKW48UVmIoa+vOFn9
ZGquEc+be3Vc5KWGw74/vjEdEwpLnAGsbxqAj4fkmS/I1MwvlY7tPdzoLoKF3O24
6Cofi2JcoaxN1byH1LWTrajgEW+L/H9/sCLXz9hPcFdfgYLNPytWtAs9TQVdL29d
vVX34qDeD5TS7RJdO5BQWp7FItfVmeb/31SJ3AnSYeG9Iu7oRhURQqyIh1tQcLnY
zFSUw3p+maQxES52ZLqOkfrBq+TjpOxP6XPEzIKjoBlGnjuRcX/792ZJQydOvwvG
RMzcB+j0fYKmxZqMZlCL1dEdCVK+vpfVpb0/5v8J0ZLiToudHEPTeIH11t06Slpv
oYZgMjlMWZEgUetxeWjIfJ++r3qbeOv6CxpLUi6dSsGcS2RK3pe3Dkm9ikqGK79S
tJT0cMLk6JowMnQD09j2TWb9gelkYvfxu/CMcN5eHNcu1wNQcVx+AGdDoyuM+laC
4Ty1UApQqVJUzXbogMSzSiwH22ESaLgJ1hjE8tioRzdWmnOdIqFW5l0Ru9Gnzd4k
LA+W7EGnsax5tXaLuIILXyuycxeIpWxIPIj32F9cHlY7wSm2CfzZcDEJERadhy8v
i0wsPUXCEjCxP5tzqRw/xSsArExJQZD5EJPO9VapnA+S2WsGnwwL93hX5CdAX62H
NivGYi8UeNjpAshp0Uc079Q9zfgOmM6jvrnYWbB8BmmGC9XkeyNYwOH8WB95E0xF
1Ra4zp5C5GsYDDpHQjpOcJJ8pX6KO3C4mTrnMThOnQkzPTC+fRwkq5Hc4jtfP8Rt
EaOO8e4RMqBucHeZx/h5UP31X6ClWMDhyeNsiRuYg33msqarudKxxPXdAS9o0upV
SmegSgqJdGHX11Y42h7zYtrrqTCeqUItCIzpUYVG4iozUTpwUtPeP5LIjDZcTEuI
eHr5aNLwoyQzPZACr4XrOo1CXW8iFrGsyrR5CBmwFFSuKb5ecFt3vVD9rXjKeDul
Bzyb8wuPv1CxXSCYnbUnBEwm8Gwr2lbkQBPO1GKtogADL3hsX87q/H9C5qVHr+Ja
FAmJtp8cFjxmn+7ZN932kS472G/q5U4V86fUwYZmdECMeTRG5SiJdPztIdAjZ0KO
UKsRdpVtqk7RngvNnlzSAbZhfBWcYEI7+31gbtJtMlh+aRrGkYdiFelEsR7MaeGX
yrlUVsDTzEiLfAAhZCu9Uk7f2+bB6Ll4ZAgcA2oEAlxUCmA2pk125jQQNoxBMiqe
YwjX5+eNRMJxai8ADyGi+498XhlBhW1QCJ0x2mkrk1CtR7F5S3sQYu8a7Y/n/WuC
zSEhiMqGeP4VmURfaoNuANA3WUxVLeOHeQ3/ZY/cDD9Of5Q17vZNhHeUoS7yPnky
75BNFpVRKa4WnSRvH1z6PIyvhyAG2GPawta8Q32Xeo2q0CnytVVUl+JuWswVKtYT
KVsE13KUNf7BonbdxWFAEVLEritdrO9CmST4Qr0qx3V8KYk+qbrVH6An6buQbI/O
rrIp85/s25v+NHV7dqIXw8+yRp5SeBQQ71hosA1WyGUm3jcBkyLL0iUVuPlPuxnP
7di+wXOEiElEjyV26/Q6qqtVQK0Mf3iPaxugzqhosc7HiJ782WKeaZDMp/Nvbfza
8cySUGzzjTDS+qULpSLKMZZujtm+MyOdXmF9kskbgvtAa2VBeH91smxyISqCfe0B
G/z92CLYnY+zcuspBSuixQX11eaO7H7iPh2gwS6tv2Rv8/WwmyTeZGl8DZA8uZFK
2K0/xk3q2QXFvSAkspsnYv9z5oZeLwZy3MbFysoxrbwLJGR8wafXQPXt1QeXTYJZ
tCDWaYrl8ENG0CGoBZvYu+uRhQB1JnODl6dKBvYWXliskPiBgOTffyxJkd8rEGnR
uQAvY1dkaxsp+R49wUM4Xhg58gMfBx86zitNuXnLbjYnOW8BcrlxCd56Tq69nc/r
VAw0VIPqFZRsitRqJguvZH7RslvroMfqY3/dk7rDnFLU+9gy8ngwjuzhri7hUOAg
2lBi9BSrQIQrR/8pOwGvtdfleduBAVvt16kZFTgKQtEW0CSqflfqNCa9yyLhlxnl
E7x5N8Vt1oibi8DHuEF0mqSvcTaZvEuNZ3A45ZDRFdEV+lZWBrPI2dmroI/a1H3I
8mRHnOBAdU/AlFVod4RJs2+dXwwFbmUsTLZrFZLxVnyUAKwyYQlQbeqb17ZINIP5
YvKQIMLKE3d8z6ExsznbOJ8+GGzeyr0+Dl8DkkSwXsaTaWwCI0O3GcARpGLg94+r
gI/p+2TN8rjw6rUFXLPC+HwvZHC3T9jzZGt28aZyDCCpnIaE6td07sjp9Y3NsX5U
lg0Uub0W7A4mtqWQBWYL1uU9MYgevKU9J56brGsnEhGJ1engg2LNmedNRot3xU3p
tivkMFnMUOFfgLDjkOwgvHSzcQXipxH4YYKNKiWVO7qYexs7ltjGTAYjEjNaNiSW
tYLhoRQjhq5Qak45uJBmHsXA+LPu17onwTv6SwdMy+ZapWcVrJJ3Wacp9jar/EeB
kpXs5AiwurhS6XXQfOpXTp+FwIk9q/2Pv+snvl4TAuEZtqB3l8UopAUoDcdcrqSW
hCMWc3MVqIG/NOsia+JOtHBIwp3/129AcfLQksUBYqnJa7zL9PPPLh1Sddv2IBLY
3MgxgTDRR7tyoBjDEiWaKzGAmRzdeasCCXUvdNef4gdkR3GnKy7eb6/c//lJiHIT
Bo0pqYBrriIyFHtGsFR4fT+L73vH+v1eFO/76siZR321JTS03ENrhios2/+56IlV
YDcgltpby/m1R91slBzkz9DcILDtajn7EE7me0rCezQWqSXFAlHLbFjMgCyf6fvV
5XT+rDhZ/ttk/dq99vHdOwP2jOjmLQB0dWm+XM3fuwMQrSZBuaVqqcQS8eCsRtiV
ZztXA0MHoon9Y9aoqvjQAZMDTXZ9n4pz0MS/2EwS0/NVtEjKsEgX47cKxwezsAtr
+fwYqa3Km2EH1I39w8rdEhr/44UAXbrIq9aG6e1bLz8vnHBU8x9e9z3Imv64zTjm
SKqdVUi/Ve0Ii7XAn6icxRq4UjjPdMQiy7Z5trqZ1aB0B2wSKEhM1d9koFzXk0xF
QBooxo0e2pG9s8PKcJq5Xy812tbj4fqeNYyON19n8pWm13WPV39I5T8BSt1bgi7T
MV3gMF5QbaszjocZe+hNIwXbKTa8OjusZ2bgsQE2twn0bmVKyTsciP4SsxgMoIvF
a2AC4T/TunrNpcpQ9wCRpzA7F9BPbLQPxSOX49sX0TyIYsO0ADgcLFtgQijSJFBz
VkXssSR81QojBoSkmblPO7yGl+Sj66HYExIe8FfzceLoGkdcEys9qndzh9S+qKV5
ru5gYhJABI0OpNfBE7MgwbO2alP83cObHswni9tJqOFWR1Vmg5TtHAf8PF1SflU9
iYkeECyVpBpWAPmKCvW00m1aSKy0m1JAfiymSruopXrw3DAdPj9eo0g1Bq5zbe4W
g85ISA+sW5/J2E5VduMMZEglCBJzHDzMxajMPJk8myXbG6YZx+rHgWoxUOxNlttY
5xk5vFyUUkWvWOnBNjtWGCJ+yITd9bevp1Nxftlb/ytuVbh2qhAd4Alh6Y4o3RtA
ly+K75O8D3dAaF92ySfRSih2RlpFHFMOGklAROoRIb0eedp5mgehouub/Chg1Du+
gBTfTbYayk71r2GIDx1clg14NDCgZz+UxE2k56BwYFZkLk0tJ6+4ZTAvyDpKGPcC
vS8XwB/mUAmthjztl6bg1drJDsv60Gma8+iFvUFAlrc=
//pragma protect end_data_block
//pragma protect digest_block
YOuhCOe+bhRqLK0zghITO1WwaIs=
//pragma protect end_digest_block
//pragma protect end_protected
