// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
pBs5ZtSWwbsRrBH3JKmaSQMV5GWTZbeWaFgvv5W2e8iY/HF0g3TqecDXEYzlg1iA
WJmj456FRZa0B4N8giFm/NYiwtdnpeLG3xIDVTYOUz8OtyzMjm822giE9u6Saex/
xZf/7Q7FZuu3xLpzcye6GRXZ3VnChmujw16PeQilSLU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 15472 )
`pragma protect data_block
qesk9dp+wz0fm+8Qw8HFLnMODhQbWvOaqa6kYD4+OcK00I1LA6dty8TkGUcZ7buh
YDxGT91ledsXZeJsPYVO2UFJRjEsrhBTgFVTb5UK/P7NBycvpiYX0Ddlqc4KkkNz
PP+Jh9F+UfBHrVimQCMPS9YK2zTnflNL2tUYf7RzoP8QqNjKq7lxs5KPaUjp2kAy
DmFF6qMwCegDCy5tCWW1TF6YOm6swbpLgw3o+Bbto5VyhG5tNt4OfEYjqJYN8ETG
5+t+XavDeqUIQoyDFlR0FHqxH4UnIPnF63onCpy99Gx3myFZRmqfqHKMiBruUv0S
GjXapVe7HaTmeLNKEmO26GSIyL2qhmrL0pmn19KpTffbny6A/CKdPggkczbZijsW
JreMrwGlO6gy11/fjMxqXDL3ChLOSasM9TTi0/LTv3zl9oJbmq3azhzZ1TaSVvaW
Gmm9vI9YxhkLUR9VSGM5PE3y5IvLWeWCBHVE4WMbE5pdJqEUHEagOOX4LXVjE0vA
mOehW1JfydfqpZisTB75UP89xQdSc6Wo4SIrKIzMI7T4R8W8vL1WmfksVTwGOGgm
hrgOoeTXf0kn5/WAYKn3kmZPgBwE9+AQD2SWtnLn7Zy1VepDud3zt/RYh7WeKPNw
IWSbYOf/SQ5sjpOOdqD3rrDVvJfior6sckd5H9V7T53eccSkvyEnot0ZrH7KpHmK
C+s+QP5XbkJhzeqzk3OwssGkOmi2iNlmLKskDkNOogoHM3V4FRE1ra8IArBIV75h
aTmnUZhXeVumvHcu4Qp/JC8UHIjkhZ6ZMsJjZnrSRfq4P6Q7icVB8VSxgXwnCOKQ
3+d3PeK84DXHTFjwmyr4Xi2jA0NatL63dU8WS1NHNUDVRMs6Z2wvcHtqUS4JpZ+g
+OWWElCk5wNXfXVWUH9OuwtMB1W5q0SPD1JdyEgjbkDttEucsmIlhoLZ5ZF11ovD
b1vWJ7iPRu2J6W9GhwaYBMeBEu2BvSGfPQYQlsupnkXf0e6DhAFt9av4ch5yAP2C
jCxf4mRyf0AAfsBbeBCVZqQ9vBQ1yC4ZzItUdHD6d4+RcaYudAuOeg9DVBcmVInh
hkaQx+EmxPpnB/v759p6YximhXkWsv9VRpDJawRaneGD0UWt2dx9qPHa/7Rth5F7
vb4ut36qPPX9YhrQ9OkWpQMTX1x123Ra+WAWcd9+ljSSKDASUlD3c7ww8E8Rx67t
nrcpTCeFpUa6hEJdvXEwT4qMnk90VpEa61SYjBwbsD49mP5cyvDfskhHM88eNkmQ
nSsJOg5MkDif1nUZ6D20oVEL+f5VzEG/V1917Dy792Z1zP7H3Jgd2tdcFLcUpwLN
iRJeIVRIG+BpuY3P+MADlZ7lucLhwaO0f9ofvExmu+4g9U8L+4qhHANdBAGSlOOn
kbFcrV4EtKU16RiO0ZOLfRBl5qmSPDPF6IIDnp+AYhaa8rN26hx9yBzxYf+AwpnQ
sn2FWb+PXEx/8Ow09xsX4t+2SITmL3C1Y9/Q9rBGs8eSJ2JEkpACMtU06vZPQy4y
x37H0ioH4717gk3jBJrXjSXms86JlxEel9TT0jQgdQSKjHURNSaErHy+XGKFni1B
CBGX1zTK1s1g+cj8Brs6A2pQlm9BaNynjlnPZLSr/bNscLjO+zJ6pCb7KOqjGUfg
c0RfHGCvyetxBnKFcDjkO1ikvhCyFbfu/fC9A8BO1DjQx5N4WXf5XdtE5nl4sVNW
LsrN0S3hOjO1s0+NB9+oqvcAZjuZf1N6Ie73Lgf6DrARXMb+z8UQhelZLFnEKrpE
H2E1VATHH68lG9AFyQXhdAoZGoPmiLyL6YldtUktQ90uWvKum5oo36AL7750mnkP
gGJoPG41s0EV0YMzWEeDU2FJdGjSo5oqYDoRC4MkjNaDJxyBExmIj6nTzzGF64sg
o6nBnkN/CGgaNtCJFfUQv2k/SQFlggMc4qmstW3IC5qgC3rDvfQ4psgpuW/bSIVn
CxS84iUJ3zcfMl1WZ+xasG8yLDj/BqwBgD61zKXQsnfQH0XZMWquhWKnBqDqkAVc
UmxtLWMq5W8g3/f79ZjtQRl5VXF+cWpZrEC/Ko8LhNZyd1qCubsYPuOl9OBRfhZt
5NPjTZyhYxTx8G5JvIOV45/2GEHs7Shl8Au1EnU9EG3P6jr+Az2Kq2W0jsHbscIX
0gnz5sQti7eSlQ2N1WxyzYQ/I6063wY0EnFjoTfNwwDqa2Gq11b0GaA0t8gWMzLU
zDJOSip9QSUyNq4ujaOvLIaO1ilX4Ljh+vaLzxmd0m95yyBwsRYyGotcfQD28G0Q
cuhWsip90x3q0oUtYuM6DOW3zF20FNSpdtCeKv52RCO8XDLSINuyDESem9uTj5eg
pex59knlG7Merhrg1rMFKvLZFFRghDZZysD4HZ/uxSGOAHUEByufa3okbabM35Wf
ngUFtfRThqftUtGYFlFu5G7LfJimZQINpEe5p2znxRF3Z0DiBwFEC552kHHDw0rG
Ad3+c03f5Jb2rzn8gJU8TYyq7kX4ynuOr4lBJDxoG3r06eN54vxFdaZ+rJ5YbjHr
gBlo5o9MisU18mKZxt6ETS8JZDJ8OSUy+4gM8bVI8NJDAOuNnSqM+hX/yCO+OD0W
UtFl126boB5Sn5DehfBUyZ1vJ8yRPEQ+bpnwmRvLyB5TO8nuUu+MKfARbwyShs+Y
xFWBpMHxBVWmfKXbieUse77X+I9STDprVxASHacsnxV4YfXbVr8+OsNwnxxJlN0c
udR1IR1VmiwR2E7gcVIrNLOkvHAr/sBplg4gE+Vq5zOYhMnajWSRz8fKmiM9TCwn
WNDP/frDqO8nsLgwKRwsZlbiVTQsViMPJITc979ii10qUC8CYAgNXEapFG5YHrQ9
BW/QKOGYoSe75jSizrFTHO3xciAugs6CQNLnzbQXrTGrrgTvtswthDLXftvN1ag8
XHybVLvk0Dr7Ws32hljxtVbs5EMUGRusUwAls/cKA6w3b1FrCQG5vvpVH2Deikyg
G05LnTQHS08KlXnDhTLXNqUPhT2M/8EKBhUHARtwETJlfPPb/aq/hqn4ULtLSm+5
LmaNlnSqf5/po/zJsYbRo40y1YnVIxjvPgO2RvOBqgkX6wdZvTKmZ++lY1898U50
rYXrddkQAYRJX4ZhKxYuhom2EfTdLXVGN3he4ACo5qHKUohuLG9YGshLYfSho0gz
nYMrJhVdS7ZxzdPo5ysy9HCtDK+MrJgnmJI2RhxvYqGF8cfcMu3YzsM1yN8CWM5Y
ySfhzDeORA3nbmK0gv3ddHnmEMIfKQNn5uFH5vqwiLhrTyv0kSNaiW5VIs9HVqJT
RAywQvQxzo/NBlAi5VGaUJg6hPv9xI191CFUQgLUNSCzwud9DKUu0eQpAgyJ1eWU
+/ZShXR727ztoswjzkO4iiduJ4KMrHK6R7cq87o3gThMp+KaVl2nOLsrh0j5YeSB
XSVO2MGXp2yXv0Px5Y2PxEjPQmj0Xz/zG23YfnnIQFd9KkTJaAcVfc2G8uRE47X+
NiEytmaC4riPLZBDN3/Qg39NQ0u7D46BxzIsSnCZPAKQCCP2Zsbn64tvYW042AQs
cIA6k5Y+7P+T9nOKyivQ+v4PCQezLVnyscELKeQoBIZi6A5Dksi0bPUih/xYMRIu
detwY9pdI6lxBJyB2ooNKnF7NXxTdX1f0gB8ejCzkmuyB396MVBFg1IGeujGDAgo
lyz2HxcFgjFWm6wgZ8YxDrwmIMSgyFLXe16q5ryGl++WKfhlCv5Fdda9IicnksjO
63FwEhDQ9B1+nBbMAKFPxOidGrg9CpUHvOk0hR0/RpiPNbpAI4haWaLv+r6qps0j
QUiunXA/47hIDuyJyOFg6G9hyrfSUDY347tFspgotY9bm7IbQis9mtHU2UGVs/mg
SkMA3BZBeUn6dRLS/DO4jvXx8T0V4wUDJHoWJR+ihfrmzeGCoyjYxUgJqq8D79Y9
lhzNRKn7aHuyn4xIV5plDPyptDqCM+gCeLttL3B2IbaHtDWY0cyrZnKvJKPpCNRe
X7uvnIb2bjwVbTZqeJOCtgiRsgEnFplXHqY7YpkI9HCnyM1aKeWikkDlP3hES8oZ
iq759Sr2FtduRDPI/PxFNb0gETHpfQEVN96i7lJzXJOIpFH36T03mshfKM1KsXZa
RuJRvg2GiRdyghH1qR/520YUxIFYZvcQla3qioiKdaNC4MZ5wKflmA65preWqiDW
bYUMjZxzc1p7lPOwaqzBtxFxdUvmRbDa5H2RZpyPkMFGVEo0Zml3gegJTn9utXmu
2EAKmalcjAy9wSoLxBFwTluBft6eW7zdBteUnxZNb/0zOKXFwtfNim0QAH9oAsoD
W3smaqhBI4R8vWfB2DpHAjEeE7JxTqKKv1X3VroDbC9jFOkyLrW2ykQWeqOKzh9h
DNbN3+bYT4n70YhOPDQBYmoqkQ5ek+qMp8uZ+MKbcZXQJcufrMKy2hFnGDRangRM
DyfK5AzalL3PribCYP5+QkNr6u3rjPlunO9Z/tJkZ3ow+bK8PQe3NfvRSEz29n3Z
0oFIwZeU2Q3iqAu2blAfAlQ/7OLterUQx+FCBfzszb/zrAyJ9to4YhjoFGvBn6L2
OJntApgpuFvHfh4l9ChM55zB+s/0pwF/HwmNbud7sC1HW2ukl1hPrutFylsD+OvV
K/Wzatqjp2A6hRtebX8a21N36im6Q46pQBWGIlUryMcvCJmAm4MfItrqFF8yWgL7
hTrcXtIhN0f0uyYe8/+t0Nx5dyMzOP0icHVtLwmLW/iGAt8TfF2PynSdCIoTIpfB
u8qIuyyck+GIy8U5UAMNhJ34W9QuhvpGpHiHTswr8y/LBNNVuCG5jouT4JuT69Av
CUOr7DuS1cOg+rEIzjfkxzB2h7L0XY5iA0RqlUFhmHEz1H+meekLH1VrO7HIdlWK
iFtrrEWz3R5NvtgKNUptqo89b6wCwjimQ+YiCLHVceiDSjJ5M5Q6Mh3+E8YYVZNU
rmnZ/I8gIcKOlpqAxoMxyCS+eMfHQq+XjQ90koPi2lNYsmgRr6bgN1lfnGtd/FwE
O3d3PHIOdlBqgX93v3hYqZ2IDm13pNpNgxiCtS9v40dQQHeuH0BPKb8g8DBW8OQy
rGJFHqErUhx8vg4Qkmstq1s7mefScolwXj+fH8B5THDErRdWxwHwWYKAyOqHYx+S
oB+lWj8OmfuCSsz4YED0AUvNfr4hk5LfBvSTF2dhtmp15OUxWwCvr7gp0TgOolhd
c1h63HQ+hU2/EOMeKEA/AFm6LeV6+TI19GLUkqmjE25ap8YnqreUuWwEK0T5+075
7eURmHn6J0Tyvobmr8izTi57qRgzvMC9EA0XqGaABfHt46dAuZjBbcoVPTVDkfo3
eiqFL+k6e+XLaluMFZSWvXusel03m2H460wjkDlDT0vofyg7rgXecGWd92CxdY3W
e2eqtCcUHBf9cKxThysz4xc5kR+LXxt7w6NdGiYpLJ0L/CnhbZuaiijTbfzQcnFg
u/rat58C19gNFkxdcvjahW79k+NPAMpUth0a8L3FRL3NEPyZw4Y/GDk9C9oLbUU6
OXJbxxz9146W/iSgK45Yn9xdwj9prZcFIgwUc8cUjHJC4ZjGA9kSecDCqGYQ4PQv
Mqogr8gqMU7KH6F6wi0wu4uVA198CofUtDCNVsRcPRfpOOmhrMPtdc4iM9R2I1L+
mBg2hXNsKYGJ/sU8jA0L7HF/lWr7qo20sIiViejaE7/fmraZM1ImVpPQgGAMxCa+
PGIsWE/6Kzlp/VdsgtvvNebqPoXizlDidH6lCR4mlWjdQpOc8Fj6jTirRR9S2kp1
rwgf02FIKzwmO9meYuI3Fq6czpEDtDs6DpMA05G/z4S86e6mF6Xy9dlEViOi8J4q
tB7EcDsrJyK8NYzAm8SRFO4OgKCJlxtR6LsM6wHIKpPp+whl3pYRjxpEtgPF9/n7
agNdy3hBYkhNKNRQA1CiAE17brjHp/yf0Hwy1WkczkutSUuoxtQl/M1n15ZrY31o
FrQ/+DBSAYLaZGtEDHeZ4bZwX4BfbOEznLIJPeSqZKdACaRET7zukMJvA+Np+stM
oeFXTvA+zVVuAwKxR5wzE7Ob3eckYB7cx4NMSrPTtRhf+LngenJRqLh0Aj+k52nj
n1xILqhbZW3nPyEQ7l4hKft+zJ/dbz5N0OuU12ew485ZA0LfsIwOX5mTmeYQUXO6
KTeGhMQrRL0Jlwkb2bgHwVBKLXK8ipcdXNeiaGCg0mg/MRICnYYVEleSiHY8f52i
9fvjij810vqp1+oDLnjWW4qFG9srGYvwAGpZ+mQc9yQRxd/whse8cxbVv8v3r22y
E0fjmFoMoD0MlEzF+DR/Gy+psOV4T7QkYxY2o7upBP2kMJ0XNsg2Z+OrTQpExo3B
O5SyyUGqUPBwGx7SUuc23O5MdGv3V9LzLHJ0+J6QTHwY6dr6BrvU3fuJraGwjWIJ
H3jqXqX33YJIEWI+mtlmB0dZ2bmKrF8WHDM5HEw3Rks0MGWrGHAU9+aLPQ8ErtJf
CFXdshlBB+0GywKY/ET9Dg9XHSkFR57kIVaMDYCiAqxLqvLEwMyOs9FmgnobVA0g
vSn2/UMi1NnWXl8AgYc8x8HOB8jZn8EM3psk5nDTaO9DckBd7yuGqzqgw9hRn7Ut
UuhtOwyKZjEZDEVDK31BrCoLmIJuUN6wDga4rDKrG1XZ7+ciBrMUVyuZMAJQBaGL
+V0N+zMQVOj0bKfx/exIWYZQhdkvq1vPRLhm018dkSMbiptak9xMmzfRcC4wgam6
XlALmWnsLy4yvPmNM3VxGRhhs9GSBftR3n/xiNPNEk5Ac/WJWK2AzN5uomXF6XZ+
21GVH0ix0/1VmZ4hyxLKUowqyxWyQ0typDxiyIQodiUjnMF9qqbVG/VcljOtmOEo
5SRu+Tbxw33AZ5TTyrJrKDPEknDvCM5hchudCckMn269Bbge8lBzwCESBvlVEH3Y
eSDk6dFIZ4WR1DQT2RGjQCdE8F34hH4cyXh45FoDUo6wE38DNnU1XIMCvRCiHUGi
I1f8RClP8HRO4AZZBEzjJEe3ipZG2XP22UvVc559LUaE0MPQLJ31b22ogr6UvtbK
kV8kHN4oVuR853c8jxTMloNMbmy/JkVVYZY22Cc4Ti+x9kzqLzT9vUPvhOxxs0xr
Dk56BJJMfxDeBadN9hPmOZidbGSvl4lGK/DlYT4o+izVvwb9T4u5f8GXwSAGEVn7
MQmnvMwxG62ijl54rRmQrzUJ6Feka8zkVIqqkKr1mqEGjCtgul55/ejQ/R5mYcxG
7Gjlk0yXnYI1i+NYp28UG3k/ZbeFBB/EJ2E4dly3tqn+/wVhOkMUgYEDoFLVnNcB
0u3536NfhhaybXsvHqRfmES5w9VfZCpL1yJo8xShVjejT1CqO3PiEdo9ZNc394PB
n5xKz0urtbPnMi15zR26q4EnW110xxrnuNgtoCRFHyhGkC/8rk2a6q4i5YbldUOe
rd41Bqt7/4Lwlghf4gsZHsf7g54SU6qSpxBx4zMHrbsSvVcfGMxfl4+whi3no3mM
H1SSemuPb98tPYoF9lDTypi0CU+qaa2wXM2xnJbZ99zVtfPhgrnbs2zIXKPlljqf
buV8duK6lP075p0bZWLHL4zMgiiS+NM0BaGpWHIQd8J7DRxOZKf1sefjYSu7/loW
h96sdDhpzOSbdVteDg9/xESIVUXeRcdxxELgCPqRurKUuf0rUauBxq7wckh/aZOx
vIHs05o8ai1csgjKt6ZYxLHCnJNBcWnqz8JIozRVCBL7llywbr+2ZOLR8XPjR3QM
TqXtYsUbZZUlFRo/dde+WhdmDyvlEFTnCdGn0ii5t2jxRYdhcP/w0xd4SyCkJrEU
/8DRKVU+xnz+0Hsxt3qYlsImkG4cYLJ0Xn9NprcfCLcisQBph9b5/HVBPVnfB6NE
6TXQAWIWgOwFBYB5yG4ZVAyiVfksINZdudqxyTFFFwELfanGQX8JrI8h9qp1yl5Q
JOcUFgT26NtTb58JfUNmVj7SzNJmZm9wymwxDDZdHshM3mFzBLq0JNARIzFvFSgc
Ya7LH8u3sRAIsv9dvgZsduVbunynDjhH5/4WP28v2r0H3pK5tWt3rt9rvgKL32A2
J9ZxCOU3QZMnm61DB9j2aYtEIicqDpJMPMAtaS+yrHwkLdVyvSMy+PXTKO9i+eKg
3a+HRZVMS/IX7z8tPfUnaCTf0+kyh5rGnZBeMwilC0OBj1Sk4Ow5bK2gLXCX+lma
SJy7T/wGWFl7vQRRd1bwmbsGLrYgdZFrOxC7SsV6pmZlwVOa9s0hkkyM6JEoxWtp
81eaHRziOLxOTmwZE0CYfJFxFHep2A0MyO9I15OyC6gNY+hm7WWwo65HLIwn3O3D
ba+MNBVfbzJm5NbLAfl1PYB14ToaW5cPqsfPtVYJA9OQMrjolDaWtqTWTkCnKB6C
5WfiA1aBiOM9mHKhGpfoaAHDIUiyNumL71k6FytsZV/eJRGU6IrBrQCHdDaaCfOW
E4k7gle7+pWemZ1swrKpQubiOOK5XeknQXdxZ6/5IBRmoJh5OF/VIjbw/JNsObB/
AxP17nfpNA1ecbXJa4nMbiOWFruSx6ewuPviyPAt/RRRO4Ni5K5PhnO6XjGxfmMz
9j3Pe/g+zfNKVue+qVa7SrMle5Z6zqMeamYIktnOV432aQFm59IN6MdQW3rQ/QJe
IEYsEbzl69fqc3xbZgurnuQIjiWZXZcbiRvAQzabc+F9ZKnET3pPohj30pj0zmyp
M/qb7xNgTbSXQveA+iSIfUplPRgVEqLEttgUmCgdoMOy/JEXS7ypUakfbcHoPl1g
QfH5hvTkmrqY79UxmnHLJDWzJeHMNoq3D78QidhPTw3SINnRqThnr+y//MFhlkON
WRTdjKTNwJywAX7AF+wrIxCGc5vPki8Jlhb3LwjMjqeMv8MMPk6uBIlXuKgSscE8
GIfcwEsHbxOv4BdA38mBq7w10JVyjjYxK1fLWoFkv9HGOIGc5n1VrsmUr19qWM+z
RcZrN27ArQy4LxjG6MToTHZzJsuErQOzpxqqg2jB/eldztskfhbogRoAEliEqQ0w
YlDQC1KAj77ss3yTZ6dgnHyuwT/AfwltAFgSbvh+e2jifgWd9uJiCYJJoF/hATNq
wQlJXSwTcaGCD261mRmLfbjncaPTqEdXkp6Qw3t9qeetYjDqFQCu0IhPrauz2mR2
aXTNfXXp8+OMmWcoPrD4TxnE1g4X3fxWUmUpZV/B18+zmQIUEqR9+s74AzifWlR6
rUFBbn49JOHHRpgbgLeSRpiEzGuqaCrdXl1QAlFYEhuQpztkZPR6ZTgUQT52gDaI
KnZKi1yRPxniHYLdOyYpw2Eo/aHnktGH/QB49mzz4zvF9gk+6hI1oSEVdgcHhb75
QXZPFF0ydbs240fVc5u0L5haX2ln5D/iRQGIVaPzv7egf+w4DuqbWcxHN5kojHfX
+wLDJY/t4Sqk+/W+veBzvb1fySP60tYwimdE9ihzGqyH//gCnV0WfPVOQ4ELz8hF
KIR351MBYMXATmV3wgaI1BM+VI+tEK2tZibbp4fxtQzt1GV0/m4VA3OkWQ3X+m4U
CqPj0PEBbRZQiyPgvXl9FMHKEIjIe3aU/pR/gngc3ZGMBKV0EBWP7MjLxvTb8WSF
/AEODGH/DePW/g+iI4BHIV5FLz+K0QC4w8vKUMnj7w8UMLdWZSiXLvQcdcW+Ch8h
1zL7/X3w+ggMVGp8Dst1c+du6ZnlQYGsTqz542p7rQhw92x3mpqZlGBc6vTDWGgj
ZIUlQaqz4NHbVC/K0z0D4Ct4JJkS1uEMKQXNcBrQduDi2hpg7oIzKdza77D0V4Nb
L6jSv5hYmscK/JFDaOKzXlLO+1rfw2gxgJnFLXBTsLZbscv7q47JlvRlkhZal8ZY
h78YPVb46Hgod6Zfmuqglmuh1PZf8fN+mILbpFC8dLnvG45GsvEzwcXFsY4tjjjg
sEDt/7oWeT/AAbG5E0QlrZKhZwuWcGZnMnyf3cWf7YvwejNpZKpmDoouTQwyn8Ur
ETdH2zuAvMJYXNEhuCeCDpyVOpWXBWKuXrllNzIkJwbBuMt3dd9c1LiwxSUmliZH
WDodTOtGxkGgm0dKlpLaibXJ2CirDjWprUYDO2ApS9Z3dE/G+BcMQVZSZEyTRWJv
rOVfw5gGKskThI6ji0tuOrdrnhU6J5bjKK1pgxonggI89talS4PcZ6tNGNS1VEBR
Thy1/ySH47ggDZ+IRpasrVrZlkBQopmaZzKczgcEX10tu5ew0JI9Jrw62WXUW0G6
7YUvYXxnEVcTtYmfRrA8SV2am9/TIpszk6Ypb+VliwzGEB/H9tjciDmSoM5VI4Ej
VLPJAfeYwQC0Hwgb449knPAoOEXU7n8Qgy9EI+HZpRtbl7veUhCvnHLA24qUNVzF
XkF6Lh9m3+mflgq2OsIjqvhVwLAhYNlOvpTlResceiSTN+R05UEeZR53P4XDaZf2
I1Q0EmIgYJ+KYXjE+txd4lij1fhiLWJauwiPOHMXEVYLnrkOcqYX6mUiKPzgM382
d2ADfu55/rckOu6qbFEYL9q7AlL2nfEFmp9t4JN0KN8qnKTidAGXvAahizFCAtYo
XwF3qEDvK6j6gtjrl0xGJrjn8aCRjIQVdRu5oc50Wnu+gtjqPtnuhbDvQ/gW0GAB
taVCWy6ntsWY8P3MjdRMT8PnQ6IzBe62xO3fiUQpCHJcCmGWdj4JQVxxI76fJrnf
4MopiZFJcrxsi8RWkEjlIMn8oX18fKzPKuH/yrwd+WZpJsS0XcjaaY16hRxV8IeE
4tI6wIvh7k+IgpRHce5PuBKrlhWzksSmj+QyN7rJQjxVHJDNBnZjb8eQbCOmIzXn
LJmviKxTBC9U5gLgXBwgiFWxIirsqSPoIT5VtLgnJuxe+sv/EPAkXmdYriHi9lcV
38c/Hlr0jQ63qwnP+/yxXEbuQAeJhLiWdnWqJZ2USyW9HsrSxKfGau0BB0g0wa00
UeUh1P+x1LSWcUg43LxxOM/KmmAB745+oyTz9E8mTw51fsR/p92dsDFOAsAmoL4V
RiNs8qR2+L8v0V9ZOrVitO/HJ8GcWO9sRXErCWFYqZBgIQ8vyPfGECUNEMh0x7/m
rbnlW5rUcXrVn9+KcpneosehEguTbgHwbeuacC4oYWsBXWg+wvOjkVVU2dWlg4Ry
cjeIAbVFzDjs6yb6ddphZr5UGyAb+zFtGrEOJh+PzFgMNrNEQoo1jTke6T/UIIuV
GZPKmeRZHHBZrdDaEq6wuIqwAgNC404cu4JGLb4KjLLy6OgaxiaUjDd4PIzv2r3o
OWv90xzBt/GSdAk4m1HkCWZf+eARa4i2EAo9GHVMSB+ajQdhNB7CScFvzIKPKuPi
fxSqwKUkHOFVrfQ3zAzxl4m/2wT3PQXth4wszaebjzz52Bl/GwdyXk+aaanpy+X2
6F6YvgT91at8dxoFXgbg0SCGoGmpyllRjpyrJLKt5qMYV/SDPLYcjRNMEs8Ewt+H
T6iwbJuksvkWRBm7qFDY72Haqa6nsOs3J6Td4x4Q1RRukrkpbsjchrse3gESBaFV
S10XgIH60N5eeCSJqV14yeRUmDPQeyzKoaik4k28xjkqoNtIrHIGHZ3DzKmXVTFC
MlYqEk8bmAJrWNAbyfnrQ28Unya883ir8HjES5h8whzkwGL2wpelsdglhovRPnye
dUnZDe2fykLRuw5+99J3vIljUdDpRnc3IW36n13wbD4zuVpoP5hiaKig+yYQSlZY
EwhSau2dzGW5vgzDcHwZuDWvmZOtkpZLLdydx/NoYXKHbzVlL3mVOeik4daSNKuh
Oxv7MznovviNTPCe7+M/GOArMqr1NqWhXBioaZ7zmryBjxSrxQV3V3JnV9MvYuL+
RJIhBJKMD8+xanS9VXNlqa9KgdlyGQYML1Jp6jeJLwa8yeSqqJZyEvoefHVzWMrG
nFU4vBXXkfPu1ilF/wGWE5q/QQQ9pIY4f0FWB03V4EaPets7ifSuzFwg6Y8nvf7c
Gx706SRh12ZxlUGqmyQANlgT1jGbHWD7VF3k/I4ZTmfhlIaGIOVLgh1wyfs/609F
9w7txpyQBVDPOhtzcdwE0oaMycn9vNQBBqjtYzks7IeO7VE13Rkx7ezSgpr6B+JE
+YnctBmQf2FsD1khrw9IuPRebWf7H0WVs5YTaMKeeG++3/dLQDmL2wsnbFhNQwXh
fOiiOmnCv4sg+uq/Ag9adscjcjbEIswnQlgsBmNCmbSTL4er3EPINq+9+oiVWjgD
1n2oKXiYFT5isMc/2MYvr9z1dhE3XmVNpGQzu5t1AqUo9u0u4Uhki+sTbKEYNDJl
qucY+lPnUMpwhiJc2p43y8nT6Q5Y3VIuyxy6DK+7l+a9FyJS0K9Ung5EFoXc3piI
fv2QRZggf96Y6kN3kJNJ4/KWuZPNpGdKsUUQlYNW5BoFaY/UwBRgHTI+YQR3RJzU
11HWuKnDQXkobFEw+mevyhzkbBpnshN1r9OnOnZ/2M60PlaF4osCI7QCWGapI9BF
AczBOeQB9WPDwp1h+s0un81XlUeTEncG+OFnVN9pMtc5cWMuV1hKNPjlS1tCSblw
56fY9d0yb+smzwqLM8rdp2VACbrMQ+0CTcIfRRbQUkLManOdYWRvFqpsNq29iB+Q
fNn2FPI6m4grEmN4e6l+5o+UkjoBd8RnH/WHTlaci5vVRv2kG6238zSlaGA+QjLP
xZ60OfzHe9UZtw6jmM7DrdsUm+km50hVeNT0toQCy7UWiMSco+EWnYtegN78Ty2I
dQkZlsmpkRIAKqyEQCyyY/0ILjy81TjwNa6JL5TqOqzInNnxXQfHSvwsdmxU6YgP
6IxTfduQ0FMLKBnXGyEnVHu9H/CO4EgMIaCcv9yofTZHWIUpKSghVYIt6rWY1Kxo
m5mURL8mqrc6lrHAKmTEhJIrkQuGHe2xawXP9l4WiAj0wE91H0FTvJbHnW377LhP
MGhe12J7rIOih5flkifynEaJWJ8/Hk7w/dT8OpKJNqowq6aUkIJlaXx2BZNQat9P
2cTQB2vF4YAzEQINwy7ZutMkwUxfv6zzzOz9HH2EUmRYbY2Q6EmBqLXj5qGF4obn
YOO/P75D3Tld9jyir3YeEjtN4ftBUErsPu5hZwMQl0Az8/+fbN16T/ehyfVIOlba
cKPU8c19aD6c0a4JNIyZq4xlf4fYO1Vx1cI9f7wfqDGp9cSxdn+uFCzEMoGxrxdu
Nz3Y4+4Q3yWICHRl1/NItaoiYEolq1TYadkrKGC9ml4sEEDb6mWRLb1G6/8seBjC
jwxbvlt6MyGORK8OwN8cLNn/sLUM8Zz+C2TcOq4XjRWL/GwV9Ag0OiAkz7GF9JNe
NHHwiq8oqQh+6aMeX4H3ddIjRZcWW/jZzLWtsyTGh6fSHeWXw68811J4dFP1wnRy
icvIazAMEVAQait+kxWiHklhCmo7vDX4N7bA196TJTs75gq0+6+94Twgxw45u/hT
7SG4sj0AevNhRcHtgTKzPkVHhE0+D3jsIbIQPRsg+PYI0FLDB78jT4JhMKguhmLA
w4Cf4R4KvdCL2Fs2QAtiF+7kqM+podV3SSebF641b2YhBeEYDG919WDh1IWHTQOH
swI5j8cV8vh4PKWVKlVWvQnig3phPRceSPFyEpl66JfU8fHJv1Rdwt4rzpJBrAK7
J3BWM5Ixx1nrTnDboXsh4hfJAUNKlnVrHf1OsWm6DyDXJm4HWDMkIe1wZLeNeZxf
GFg6PAjhm+gY59Vli7TLNrJzBG4zTk2O/ceb45tTa1bXxmdnzmMNIQtO9q4KR/dq
Xo00KSnCCuByKGdL4/64oa+U747BF8GouxWdEBVfX/V48iX9aQq8zt4YnQBRigpC
bLOSWUVurVSAd1FHLnYUE2hONVWtkVaFpyhhNU87a+Gx9PnVCLPTqEHnacVOJE8z
HQz8a/cQ6ZkHmt3XWh4nhzIVz1LJN2zafvPVX6JZilWaVoYIg/qGjUiOB/SghQHf
r0g3z+IXjRSBF3dSG02wOMfhPOEu94XSrGP2S8WulToT28PXWZe8BCYwnCBrwOdU
hCukqCRsOmJRlnPPieaSfO75a3seuEtxasWulAHV+Tp1CqdP5KIb1c0f7w9E/gh9
ur/2/FfPzRZ0Ny3o1lDiZ2+5+u7eRnibAsuW0qbU4jVaiad2XCPyn9Z0le2xhtw9
D+7J1mQJXdVhgQs+X+nsxf+hZyq7HAFduWOz0syjG4UBDN8v5yNx8t1AvEOMPWLS
SypmsZHGvVM3amp+7ATy7nmh8CLB/VCtrI6YZzcA9fcwfacoDbTOlw5lb3wJUV9t
CLJe4piC8Ml+SRLcdxqZdv+IxFY5Nfo1+ZjopJZYjOhr9AmkJPXGxYsOishmU3an
CyyPtJAIFQkHma6QWOI8DaeQDsAngdc6CXopkoWY+ZwzL5UnPOGhhnvgk/aphuAp
uxxIVhWMDlcMlocYWKT2F82YZQdfo1verYhtghCnJRFdnr3vV4RE1ujDvagcD5OS
tlIwiZYE7jldyWaZU6zB/w7I1/I38Y1do4FNnLpWojN3lsPIsn5n6h5vn3OyXLVx
41u7nG9btNWxeDuEFEsezf3BHj7hQqQ1f/n2eEyYXTJRBoNaJT0vuI5tHCIuXHxm
aX3JeUl3K3lqVaKRBfXtI9f828CFyAQGs5jDVak7vWv3cloAseLQF/SfF63jdyVx
M9mZhR8trjkj6yWWr8tBsqx+UjT0RSVD1yL6mFvRLpD8FDHHTPCZPStFoaQS8dbA
nDTpbkrK3ZkrlV8H60vuvzsMmxKWY/a29pTthZ/D3BcJUy+w4mdZvKG/Eozn8IXw
l2Mb2G/IMwncDCP37Jvn3ndJR1Hz37JkOKe7oymvHOllZNgtJhLTLaOhxIw/93d/
Bde89SE/QUyLhB2xyoMaIB8W3cbTemvAwz8n5BPXidrHKZs1OaFT6BKIFEkTSCxS
RhpXkppZKunj/5Rm5nMi0+WzlR2FbwTzjIcG1C6tezm5jIfGuLu/hJeWM2othjc1
FIPbxvKV8Ta/Wopb3sWt5z6f9BUKePHab02Q+yFG6zlmAkhwgloPuwWWBDMFX91i
Vxk2V1CI4W5cARWR8YVMRO7zugvmZ2p4T2Nc1RwQ5DLmzAAp+8wUq/W5pqVfiabR
ZeElk3yNjcR5wLGkrqIQE/BCxyD0JkX2yrrM6FjCbvU9B55OKmdH6+SK05IDM7Ei
KFwm9FdLzI9BPPjhEPH7KUoPYzLICUippiwaa87eE/e7g5YC4F3VhALeNugB7e1D
lYws7npwuccNSsV5zuhqsBpyEkftYvkwO++UxUjviXA1c4VRIuPn7mYZcsNv7dsF
ceZaZT/nhhFMe+itsYHq3DzEkF2gy1wiuBe8+rG9Ga2rg4IkPFYcOPqZiVoKxPbo
zWvaDCCjGZRUxKSDZLj6rvyJdCcnFlsSt0VVvjp894Eek3K4j0SlBQX5zKSgZLG2
N5eXPlZA2qWqlPDkouDZbDuSpWA0JbZEHObRQ6eedWWTB/MZGm2+/15kOjsw/xlL
dR7BcAyCaUYsr7s4uLAMl4Icm1mnISy+k2UdElGVeAXFUjz9ZQK5zZlwRm3PTkGt
Orn0EctnZqfhM3IxKoKJPGRDGgWeSM0H77+c/jHOdo5vNSxLg4lH8U9A+OJJFM01
UI8g0IInu4tkad2dPLcydy64swVsHpkyvqzLFSATPrIe5kgrhL6Yl+xOUMGyvjTP
jl9fYA8Ov5FH8RdM+RR+Nm8sd+UeGnJvYBQbYO/fIoKnM9D2RW983DctngA0k2j4
d6/lyvSGYeVu4htokpB55Swe9bD3bKGfFeHK38sE14KZRTBsPoCV28PgyPFOdmaC
sYmK86WDQcS7ym0h32vmx2Qf81HCQpyl2dse7frRTGA254RTIuIr2gOkb3Dkok/D
DB/YAMawsSAZjXzq1RVV/sGXUULtFZjDpseIMwDNuJoirH2Fp13AHTFa64Y4biXb
A6UyncitHfgRKrJbg0MAOZr0VtY3rcOv7RdtPpr4n9WB2vpNfHCA8QIczOULEEuW
PPjr4lECxz1GHCik1hLfb0deSvsZvYaU7orEnFKjAMzkzwkCsuzEbxwv+wyc0vfg
7WvCDza0HKj7cK1jy3H+mrsyRHX2HmRQrXzDQuIhLloS5wtqPHeF1M/OtCdspoJ/
em7Dtcd1oR8001SaglWNosxiFjWOa4bagiMFn8ybJ4Gc/A9cwIcTEoeOtbuck2ox
onvQppKQ+xdHNKWIJyG/FHaJfNsjkWiNe7/jFPy+CS2e+w8XK/bZ+nw36ffVxFPC
zMrKt7aMl60HmgFvqw0yFUruTgtsvOQ0PciAtl4IpwsObcNWFK/mzJ1sm2vWZnGc
BfM3FIdMGwtzXE1xcDPFB7yhpU90qnnvxzuBRcm8hHsm83rAhSsvd+b/eXW+3ubv
vs5VIZGiQyeE1rdFqfTQTxNYjUAfXJQVukvdFtuUUHB5QqlNRM+c72eFKoi+sDFC
pNWPqDCCmJqsBxQfrGKOjnl4BrAoKda6y2XH9JOWovJ8i++Qp/Usf3bEUp9OiSxc
rb9ML+4XqcaWFy9n1rq8mcGaWXcMKJMLa66/vuoZ8J/fkMyWShBW4DwQHC6/ij6l
gBofA8gnsKi1WqZ7/fi9bnG4sIQ2TyIUdkLglZC16+b4AkwnmoSkDviiZ8npUEDL
LMV5zr9yAgLMe94Aj5iaQu60dsEfPOR9xnu7lxlcbm/b9onyiYfURp3OXbchb6m4
HkF/mLtAsdnojSb1is/e91dxCBUmqYaLUZpY9FaMMXqEIe66Cpqsu6hyGxALMJPn
JzI8STKYvwuDdaFX3M3qhJ/5kFPlnBV6P9rcO5Jd4mE2SpsDeaby7X4aRD0IQdje
on+gcRWZJFDRtuhLaTwTBF2zWliKO4rC1amdFMhyqOvYBpYSZ05p2zZu6lo/urFB
lwtuizXd4G04rhTCPOdJmvWhgvGSSAPfh4zXdCATlgT0IPwxbE0tfcVjqcgdpXP+
V3pIR6G7REdJySlCTzDpBXIed6bYmUpkDDNnxPPbfzLIJQbiQifXJ6eZ3HkATFaI
4UTaqOGu3CFWiA3ob5p3MQEemyPsRXtNJJzg+GERkzQ1bRt+CWfrRbnOtdKfLv9f
bR/MO8Z2vK/W4u4QAmchT01MxvibiyrNc8oWaSoEC0ZTDOmnb1mEm5f+PwAX0FPa
HFoHyTWHBNueSWh5nAJqGQn3tn3P1FUAk6b/rZUlU1XDQcAf0qauBGjFGOuJafap
Oh139KhBM+CFxJ+kdnX3iGqN4kcHMmn3NjurUPuDxaikq8Jt0P1xzjYeEsKo+nJW
HWqm4T5hVf4mUCjJa+QB4gPGOKjEVV9vK+nzzoW+YwRL7n3+mbYc3kRAS+WZQlqS
Jpl3wWKntmFQk7GWxSnXNfnw9fzz2NYwIlHXw9iKD6Mt2tq10v9vf2KNGjJKWzGb
/SNk6JV0NwssymKOLm/T/XNh3Ryaf6K7x1eWtqC8C0INQbVd/sfy0P94iEfO5KGc
kGfgZfYmJF8+4VxG2+Y21c8Od1JAhEotX9qEZZKwunfVDRkKvgK6bh6YLTZFXcR7
cxxwK2oO9cZRUi7EgzPznRFAwt2hVFq6eVLFbbslTv9685UjeYLNIWUgUU7X+Gxe
UaWMrTLpQzLEkSjvOdV7OU7uCGKxJqtIvKle8x27TdOnl/Q3riEgbypuWsjElu7L
V36Aq1n8tZYqeP1MBV49py/ums4IJRC49usWI6H9STDNpxkhL6g4jaHinX1VPKQk
CJid1onhm1rXury/vGixmWlmFb+lb9pZUaAAimfwbHRQ9zIN80YNqYp+AzgMY9e8
YFEIAR0+mPAiVJLOgKlf5CGmlJuO+BsirhHLdQwo23pS0Dvj5/GoCl98iSuTlE6Q
Oy0eCeOzHUDfNFgl2yP7+pF5DaQK4ALXlsfgBW0Heq/xKXgCMYJiNxWRdNZw4waf
UXOn9m0QHdnYEd8dxZ5lUZqJqycUgsGg76UDRJMKVEnq5qxCmm8OwdoI1twJGjEU
VqNe9rMue+X88fLqc/IkLju9IHh5nAgGP/E2h2MW2w6E2RCbhD5732XA66EAkhFR
w50zXMwgLCUPYjrP7Iga1takhNPlx+Qnr25cmaNhVAl23YlVAcFZhnvgqcDPcTJK
BSGZ1AuemzAHrQQDYRp6rxBHRamLQQiIISXems7ABSLO0c1QSZbQ7BriyvUJOlA3
lAHngNbhQeHDwU00D8gDGASucDAheNz9DaBLKRjONWqLyYZ7PtGppBn7PYaPeu4J
U88zJw01I+YuzjhR65+S/BHZOrFt/Xeu/MeEJfS6CSdTLeRRRDo41IamdG19Ofhs
VxxxA5Vd8dZG6VMfuCQ/KuaioThE1A9f3WGRQIr7ZbY84nRejOvPbkZv2LbNfMEV
2iV2aGvSqjEYYea7utW+Osn8xhJD3dt8gEE5xz2VfQFavbN57cUF2Z8jnMDcgngC
kSj8luWYRlk4PE8fv8R8bJnFd06OF4NMEvmg9BHFJGR0HZ/UIwhuw0DHviv2UDWk
4HPmVj//0SAdIb10nxySn4UyXnWufhMhbOGsuYonDS5taHXyZdJnPfqm7I+7gNAD
3oX69yEc9mIKMiqWo/oyZ/PSJy7amfOyANBiEkm51uiBVWkJVwXMW0w85eqNGPIy
YTr6tCFGrprho21rtRByXRwqZUGI0SVYrIB1tz6IeSa/juHcggenuZn11EU69bMI
I0EJ2j9BN5tbyfLxwIR35R3ZAicSttHM9ShWJjGKt8urpaExqPEUEgo7VfYqavXE
6+IGeGRpAPKSf4H6OefIxaawpAT19mqgDdDIyghWyF4FKa68gKgVeBqDnh55lBjG
owlgAJGqtZNw65+9UXGIupdNTk87pkC7naGPIna1mTAjDRKIg0h5lLsciHnIBYuh
+xokYRbJE1wGF2jlY5OaPSLNIJs0/W8e2PS8elPuu18cHyr7Xvjf74YbLtCKLCa4
UgPedOkVkXLZfqtK89TdE04cAGIUdHrpUuyEScQoHbEKTr88CD5fCDeDlkcBIZQ+
75kzduzVhmAmVPCz5YZJFfs4VDtmaTv16VpxufFckxXlTk012sCO15x7rxY5K7DS
O1PPWEPJQtF5ArnpfbCjNshpbZys5+lgWzkdGtXm/tcv1m/LP7dNwMGhcja1j7vm
6DDnUh1x8A9rO9SD/YDcfPiwt61X57f+OpI4OfwYryv1/pnwgtlv4xgwh6bb62vH
29ZiOqTKNbaZZr58PN9GUZPtEzwZm3XJGU+bNq7+312af1kvvYfuVZHDYvOojxyO
EphLK+L8awv68JkQf28ZT9ZWhgDfTmyk+fsa+NltC7ehiaTj0qblnqLkCIs/fAnl
luveYjqZCUG3MElJ+D6EN1NFUJ13jNG6vqVQxcfjuLnwKCK/SrM5KxaO4BcxnYc4
7f+G5IWZ+idNcKRXF//o2dQI0y105X45qtlEbc7hiHJtilxJy/HBbfaTwPWx8CLw
yQexuFZLavhqg48mhunQiZgiYjo8sAypkTkx07N7Ou1j5cmULnNCyoYrzkN2uQeP
4wlPe7fsFCVmwfco46yHkTZD+PNMpTkRQHkBGVJ1QfNh4PtuNXLeyQdi5X7OrAgB
paaDm+6TDMV0xWACs0f4BoWwDKL5qi9nE49MBEEO8oMSo0I32oO8cxSjm2Lr7AQt
5jzA5p3HKuHy8hIorcg83cDQFSQ/TddqiYK+f91sM28R70cmtPW2VXYr+CT4dESz
k4kHYkPHLxK1IyIcy8c/lUEm9zlxyU0Mfrc3lJ0tM9iPWb0U5m5SWfeIo/akR5iW
o8rQOW1gXTBRqX60tVChoe3XN+t8OixLRmTFx4wBNfYFJDODzp0fO2D68z9SCg5J
7y52FkjeDxYnVn+91uUpHjWEOfITH/1BkxH0qEKzypbJ7moMj8LznzuCFO/j9v2h
M3eUx3FesFANb1bBIoD78wJOu0hhp9OaLQ3zNqpjDDcc+XKEY25H8it2p6bth++8
OX+3TfOZvj2a8Xg4EtXTfWwSpvzSRQ93frnri831RbBlFvLJgfnRf7pAEQp1iK18
4vSBFddnvGn08vPIirsqNF9fjirqWhmF4odJwVDx9itmqw6++3YnwxY6gm5k/KrW
hrN8LfPgi2WS/aJG47hPdqz5bf3jROFOPy8EeTP9Fon8QGGLCkU5LsqfJ/6DM7EC
W74OM6dz2gUx1yMzn6zgpwIZI2OnCakYSYzGkUXXyJy5xStu1fvaxrLOtZ7PUnUe
fXT77fUaqmzfubnQqoul/PMkWGwkrERmfXqJd3wvCnroWn7Hadht//kS69JqqyKx
tkMm229B+QjJN2BQ3qGOkRdUGaOcZ8CFnIUP9PxM4868BcLNJDwRJ3EGQ8POn18d
S2nQd4oQzNQ2R+zuemTZRKuiQGBwajWDf33YRSsQ8qU1tXPU95vIJC2d2mic+FjH
NWSLw/fC5Syp2CNJ+kXVXlr+2SZ3ctyyU8JZzQtIYRTQmYKL4ncTEjdO5LSuciNw
GG0RSkIXNm+QbMIjDJx11gVJ2AlZawyEwjbqHSOYOXq9toLQMq5tp/46RyCy7MgC
6GDJpibP93phwkC+F9ZR4w==

`pragma protect end_protected
