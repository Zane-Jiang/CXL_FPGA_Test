// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
vkUvWTMEAApf3UT+61F3fj92nvTCPybGpxLGtPacrXXklZs16xoorM4FKWbwqrj7
pLONynHU1sVkG3QvsLaiXFFLwvZ82CySfChysmeW8RuGLmns5kG1AQMppTSfH+qN
OX0ZUJ21LDyTX0cG5jrCD2RVzJQGa4wrmY7429urpKc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1344 )
`pragma protect data_block
gcf6O6LSf6bwbtBqsf9bf86dCnUmsCvW0MQ7/SfgTH6LhQZPILomLuTZGIDaWKGU
k+j3MTmZ554G7HXOTkPXc4GvgiWuQFzlmuxFnTtGnucggZE1qAV6m8mO6sQxsgQZ
/8t4X/BQQqJbY47YUoxeJhLS6+QdMfwaAnbEy8uMREJZd0viIgrxcpgSrrdZ1KfO
eFisoxgYszH0x9iyKh/DAan7uaUYHBaKdYwaH8WZ5VFFjdATd/D/UA2PkXc0jhgb
C0BmqN9ly52/2fAMWtBIqljghrBGqUcu5KXmjR5o+G9CBRo3e4u94VbIfBxFyFu5
HRfzLTimqNxXr5UiSmM9ZcqYxf4eLRTaJ3fjo/iA3H4zWDEFAVE1gJVgW6IgOG7D
cLVkqCYBdje3DUFoSSN5iBgmAsCfMKbd7w+IXUl9u8bHOaCAbbl2sphLbLD6rt3O
iAAEZ1owXS1jzmfAz699p84Mdo67M9dueHZ43km8XpbB87JRYkV+lPzZLFLFcZmO
RzSSn2QzEURMQyojPqdjSmEkjvPKhMIVa3xkXIdecJhyDkzABKvtxgQD+V+FY2nz
AN0x0Ni6YAgpphhig6U8LY6nt9hsZ3t0P+otqtrvhq6n8c5wSw7I1Zdgeb19mWPg
BjaPhXiqYkkKfqUxU5MQkAc5/6SUjS83FubzvAPTN4QhUfyBqNvseCzFyd0FIjVn
KyRDrTHmuaLeZR2VpcKllHeussLTiy77ropLVR9ckCL0IX1kRK6WyJ5NwVZN8H2P
BOCJNtKtfkXTfZuCObsmrGWRe5cLknJSwoiJFciMmDyCUH4ha9AHHw0+tpDc+zfM
K2crcPhW0tzqLNjbCRaIy+qjt/MSdGIQPbd6y9ZuPpmdX6745s/6kLts/c/BVmLd
KxA3xikucUPRUohLwdeiyL+5wnDljfiVvmwwbyNpnRMNdvrLnsnY1iBHX/WiEvBV
hzvB1EwEMWE6JAI3M0Hv5yDonTMkLxzwwge6M1qClXlCUKN06QgUs4nCPXJ9CIfW
vhosm8zAJHwPMVUIE/Mq/z+cdkEOLBAl+lHBe/TnLcPvedxbFuC16lUxCTO+VF9M
++pYfC6qQo6TFu2bn2kloOmpywYXnzK5TmVzEvfuBQoQhEPda8rC0iYKP3s2GkTW
IL19lClePMvIk+6fqnZt6PAiS8swi5fb8A3gIQRdXzo3S9QHz/8voDk732IrB/4g
S/HSZhrp4TOq/uwImyLihhgZshQ2FBR1qLjQ3z0qD9u6K5ioBA7hbhH4C1CX0eN3
PISIjh/nKIz62jhILzubEB0+t86R49dH89Crdj4wErnpiSS8GK0hF2stU6clEvBU
AgejvXp6Pwvxg2HI+ysJGKbH9VO4qlmdb4V+n05eSK2ZwD/GFxF+Cwb47rzNs+Q3
sv0cv0VCQDUv7nU814/7GafW4v1wywo2ZsYIXKB/k6ZIolbNCY/is99G0Xbx1fEE
wrrEDdfWvi5XSwiDMrEcaPVqE51NqGpbQVmTr+MLvQi5X+1QCwtMsrex7KO5qmQd
CrtszAG4YMzRsEhYr6siGWL3ePkNNYuvPMOFMIo6StSdd0zHGWE5ooUEcFYgmxq0
/VayHg+8nUgeWgVj06aMyByImLqId1y3WcAK4HSINTG3iMqf95HPyBn8sr8Pd/5F
o65xxht7OjpWpQ9LA6Tl2KvtOsujjFAV/hLWIAcvMrrmlzzVz41bKFFewOVcgNYl
XiH16hEAX3hkHa3jAR+Bdm4D8YzoUeDtv0kFMOunnCN/1jpNr0NMk2RrgGjRlo2d

`pragma protect end_protected
