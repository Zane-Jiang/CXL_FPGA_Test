// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
osa4F1T3nByXLR6MHtVplsCZQpO7leloK153YaMdiP0XVqql5HOTmUYvzTQE
bvfd7j9F8YY/l98m2EQSYqjN5lkGpCeG4zG3NMleTdgRSA1G7oKLaIRtph7Z
QCt+1WPfEKjxhF2bZkinlltPdMlQE9Awy2SVc3gRRTlAag2JYdp6WEK3mWb3
CBa18T9pW9AL/a52RYX+kj92QtvGUR3MIygX8Rp/JYSkwHwcrQLBigaIt8H1
OnY6jROk1IavB+kYVW826c2cUBmNMVEOXxVPLkdN3Hk/kSMLIHI9cFE2SMW4
YqxLS4cJwzHdGU2Dh44Ln9pC5lUQbWjt/BrGXq38FA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H0f2wCO6c3tUvOBhuXC117GW3lS0GGZJQE6Z+Jxz4TW1Gb1FPTomHGLomnty
9vuacZBH4nrVz1oB40RDhBih7yC5Px7NMSmBgHz6C1tWwjmQHX7i+4BWstE1
ehKtfUGqGIDjyzbzD9/KWQMzUphk9FjvqwKR1kBulnu/YBHMrwn/W8e2CKF7
Je8MbKa0HT0KLw89JQT8MyqaQEmL9Z3emx5QIi+DSsOzs73vECmbjixOYOcV
FmXrJTheBBHd5R1Fe7ElubxHMKspn1mQmCo746ozHaMlIbopXfFSgVzA8EZ8
WNswZaEKBdvcFiLipwfU/MMM1SExgO0PCUq4phtoTw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d4yUfjybmmhScTSBu1PKDAO5amUfpS1Tj5V03dHj7IfwkQtoZhWtYNUSA39S
kBkOKKhvblBKhj1dZDUNr9aGPwul/lPSLW7ZfaBH7CjYwEPWlwIhMFmi63Im
28oUMQGcNphRgC93PIy9Wl/o2yxfTuwPkO/A1NzQA/HHXlqgfdnXTiWH2aew
hhSNqBceYloIr+jDesbOIxOuFbzDa+T8KtX2+kGk8gpFW4pcXhQyg1tJCbp+
h+fq12bYfLOWmtCMOCmp32+N2VVdT1hkvBRkq8VyJ3dE8OjXzdOPe+QaEV/G
EF5s+CuneeqaCDqNGiA5fs8mUv8NPI5pmWduEIn+Hw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aarZIJaoKsqJVTXo6MxzA7m0TFXJE7m1dnBoRQITA1/kG1VbX9nrfA34TyTt
0qaGuoSOLjFUV1bYk3sAW7IS1rVdTHgKm0Lr7HeaDeaSfhe6j8AT+xGZa0tj
E5uqVlKNpVKsWMpwyTc+Wof7vGAU/3EpO7CcurQi7+0apW8ZTNs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
f62veXKFM0Ze4LXIAddgPwEmxDRFidF3Cj5KbmWHUeaFt7V0ZlYIP1mCw5qq
yGtvz+x0ONrhZ5xpu7KZYgi0LyHxOGv+BV+hK0+2gpIAUkT9q1vlJipzu1hX
GZ1hfQB3ZNNaURk0LHewI8tNaTFV/BvTxBSPPdgGevFjdOwi/teSjUN26fXs
P2WmF8qTs6wpOGlTN+mC+ahUQGZW7A8zPzKrvbh6wy4ZuQVhZBtRKh0/hQHi
I6OqjVF6aEZIhHxowH8RW8eX4rAF1D9isVah8Xw+FobbXOnSHody9o73Js6D
YHo/j5qbExLmZkr4MdzQxmNW33yv1FQoDsOhHHVzCI3WpYgaydsjBlSB1cWa
1VaG+kxJ6sXmkjREvxSBdn0QhoykoPOi/mVmZBRcX1NZEsmIOLvwOQVQfmWv
wqk2geEhW24kCuTrrALQkwOAj/of9L7WpyUW6TqiNu1BPj8l3ZDtmHd4uEqd
5t06p0iAZAlpibsKv3ZnBI3gy0baIFxv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HHybj79V4QE9jrjT+HTFybiZdLf6kSDllgSQe0yJG7Mcb9xiuUmH9Ru/6hz1
z4HCPZZtJn2QHmr6Dyavs9oW9hR6MNHmS7PSAmqNRhp9CFQDnlo0TIyogVCZ
npiqUdMsAtrVoUg+yZ460vb0OFtBHV+wlmRqbkCGgX/DdsJJ64k=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AgoQYd04tOxx7N0PxjOiBCIWaU3H9ONv6s4LbIxWUEC1cd8FrpCagYyWffQg
iFFbOiQMOPE1jlRQmbyBr1BHU6eIrPoHVuyaRO0TXkN9vgyo3L6nqs3pl2Ut
UcBLBziffXfr7mLgIA4XHmm5H1VPg0Amar6Mo2Hdt5pMArGfypo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1120)
`pragma protect data_block
7LEeQL83LcL+H17fzyK1AnGFfxHo42+ROJznYbLaQc4wI4ubqZOhCoVrDshG
Z3y2jSfTUlhRMTh0RxpzKT1jVnGXzHHGaVj1I0IJoFYf/o0vu9xR5Bd+gvFI
Q54dwf+Oba5ROZAKWnRx+87ww0FTFXfR3FNldKDTtB+k58zLD8/h/ofI9Kad
drf4brsStxcdtWhtAkeskFfGkn7+PSaZ4QbtLXV6F0H5/Ba0DtPx+G7dLDBO
nF0vVCQyMFiwNNGYWyjKskHG46idb8zvUHV6GGovc8tn3Tbbe9P41QEjKdrO
Hz7Bs/Td9ZbUkdVqUnufaTIIql3sqZ6ekULt/MUPOkRxN419dc/YBiEZcSKb
35kRmU+1g22n1EgjF/K7nTFQ1PtTL9+nuqFB+dc+CpbApVADcjeIVde29NnG
uTSFIwfU5tK5MQ+FV5Kt/pJDUOYbYL3diwHjsXf58gRw2raWhZQ9U5JC+cyX
Q5HNX+0sTqHK05JPIb+kRKQFxIU18TSUiv5LDvVfva77/wfjSoFdGY8vpNvN
+uI/wTjrpW8fEAu0vdklPIJdtdxvt7F7ZRT75qhvS+TW297ZwUKAF/CAfhkZ
mfUijr53YrWxYMQhegLaA19fu4LoRRslv7CBJTPwdOK7aK0NQoN/uV5kJx5X
L2NsVuCtlECe8di5kBk+wR3fqG4hwXIIa41R41/IjhkmYfZwwGqp3QhShXpD
A1mPPLLCVrPK2RS/6A4RbZCmpw28svzFVrS2hXK8UPdCWqtZt5QiqGCYYUQd
p4SI40uDWxvX11NDVW4Xr/9yEDTHZOiFKmaeeJ8DtfbGba3n9cWHE3DWZ+BS
AGeBMvrRTy8FsvgVwQUPeV/afJQ4YvLuTz7Pk0iRCpf91mIt13wjt4o+jbjT
0BImgOOB1FNzUHHkHZ4+kuPRTQ0ejUh2NFTd1wdM7sFpFQdpPEnEh4rGd54m
lv5wqg9oxBKD5nYvyj/NEJUMxsYyiD4ikstREQefRwLyRXF2MEKOurMbCfYI
R1NmBR7Cx17/eun11LXpEiPFQsBcwX2Pn5TsyXtEyesJvIzoK4Un3zVfVCXf
XDlAABnlHDjR9EQNo3co8+nrbSgLO6nXDELs+sDn9mJuV6nLX1CZtZV+d8T6
HVVstn9wS/+ABzk3Ml8uAVPN7gkdeZxZcsToF6A06K/4XnpH/MMi9IoY5B+w
2qaInjPqjEa21GUyWhnxB4jQl3TDs1/AujBz2kb2wzi3qY1SLv9btPQFHtjO
MmcfJWQHczysi96CZEpzPWXz0PbTQ+NTyaKtgFjgM3BArLot0mbrkg/tH0T9
WNpUHWM22TgXDPV00w9qLKMbdXWPxeINSEGYMLq2wajVzs6FM33jHLoQI7RX
YfNVKNywcqNP5Ad21IBXLeenEUpHqVUVerOPK8eOFIepdXwFTzUH3fy4Xwbm
nezOcjoqmsmoW3cpM9qZ5pLFUQuAG8qCewZmC2n5BevaMQ9UVxU8Kg==

`pragma protect end_protected
