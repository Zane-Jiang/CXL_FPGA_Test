// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YpvftbObIASRt4+H7q2eoXCvsYrOzqTRGdJq7qFCU4d+BatVvRiqztxxQh6l
DF/lT+RAcvLG3y+YRtWJ46LYR0UHLeZxb4xRcBidP+7G+4skwbdntcLeFcXf
zHlnCFQjxY4SEWTVUS7DuayokdnK1RXY92fiRFygVKj7+EtdU420YQ5WP1qW
6QHjh7f2QmJ4Q37VschkQiz+MbkK0Ic5sTWAtilOV+ZMFow2Xw9iV9n2UNOZ
/AlcqrOa7w4cmi4mKiLrWpssyX4f96v+5hortQifn0rEdK5dt+RwbAXsZcsK
KCtWOht9lduUAtqbbjKewNmQWSz6Taclu3y9/tJl+w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PqV70GmgRAP6mx75asYfCay0ftH0QlgG928ejaY6IqEUc74SuSxKagmd8pKy
TlFoB7MpJRhGZBv/OMYG+y9TG2Cv+y0xFdNwhoNkSR7wkUEEpmHafuj6uhl0
wzlcG1dd9L9jcTuBrc9xGEXBMeljqAtavja4eUfvEwbHLAl3TB6ewsvjMdGe
i5X7Ruqxi7gS5h/RXu7mnCLD/YcB/DiqecInoTmCq/gRo48oDJ2UeuvAjF73
B+cd5+qKjKIMfqpG6hACxcf7SGJ56i4YKeVzMixdtOrr/FYhrjofeO0JY6g7
dfUqavUjX4qk2orl+wbytjp6kpdOcpVnGGueFVc5VQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kAgtNAfwAqC1ztveA7kLtpGYyRVQlUlhEecIYGPWa/KiPGdmFtaTD4aMhcGr
Ibq4xm4+F31aWO3d55kmHoSFYHPqF5MmGqcXzY9dSHrchuR3B/UDS3552vKy
QFRHs3XB6pmHfNa4EvQf6FLwiMy/8fz57OkINreZou5SswIOC6+6hmu/i2db
tVwnFPLuer8PczdR/BFTUYov0ABOwynoJj6ziznsUn51T5gj582PbbK1zgzS
n4n96elD7I079m3LVaLiJ49i9oxcbVTtLp/P3e4m/JrvMN0LfC3rVjb4uBMW
7OKmkEaRi8GosUWlh8dmL5tdeOigq+1eHjVAlUprog==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
raLi7RlIORK9qminnb5P/OpirKHezBfUjQGgVQ4uytmp8TvSHpUcgJ3irt47
19s1az9UnHrWCl059exmh4UyMtKN1xbjMKrgIfVEMMNOe8zTQB4ihiD3GIP9
v+gnDgf7u2khdLA0x4D7itLKD0mKDKpML3Pjls9XYXzyE5gyljg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VqgzG/xhOrT4xxsNnVhuUzyckc2Q+uw12Be9UbPkQbgZ0lCWmMdAKf3rIMTH
cnnjibqlSnKWmp9RCGohBxzv2vdoc9LUzUDl+cHqBxuMpueKvkhP6T5oJbBw
D1FEKWoON5vmjudnNVttvyBiCcN+rGlAYq4116PAFqAsu32TLWN7WEEECwZ2
nUrO3diAwGDv55+SdFtdQlfcoiTkWDcD62U6sNXUctPnnig0gffnlO95RQdp
IBeFB7NJGNG6vdI00FClRYNYx3rvQMdy90KxpYBE4M1jCRlTG0uYsMnYVBfu
wpVX0xicmIljRAM1y8PvdQw7GEw8+eW8Qyt/025BIUUvuXx21GqGuxCrM12u
WMXkP2Voq9GoCCNt1RLbFTKNisAm9dsFRZiM51PyD8zRNjPcplm7FZ/FDtcf
fyj9Omp/awsC0FxeDH8CRE+lrCwZ13JoTkaJBY7x3tTKgco6O6H7E4n0HW0x
bNuaWwUJS1b3AwlnwyXihCWoJa3RNhu7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
khl31+382N0IcKGxzE+kC5ZGMYuoo/rHKQM3uXM0gtpQnqr6Mas3P2GEWYDY
ce627hmj9CKwY1WPh/f3EBjDPK6S+puwvlroQvJ8HUvX0vSbk4AnhyRDZwsj
fuABS370kac7CaO+xqWi8kJ4pdzMe/55TlFdBUELqNvwgIKk8ng=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qa5FwCypXzxgkdT5Y6Bb67kTzvmTMHRibtPigyq5C7xC+oPiRlwBzYe8WsP6
Fy6LKIBN1pUqIaBDdS2sIzvI4yYqLN679e07U3we55zQYa1do3X/PZwJ5gtc
KXYQ3EhiH6qVGtzxySvxTrbVw5UjZhtZapnJLOJQMF84nnQulo4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 688976)
`pragma protect data_block
I6j5c8tBUOsbIs1vt8p4wP0l7Utj0M4U5MVVz3ntJdTUcSCeqPTgiLeP7O1u
Xh8c20Z6tAtnx4/j9Sp/Edw0ZZuOGFep6cBXCLyYBrkIXpBSZLv+S2+S5AqZ
SOwLoXpk3UTF9CwxlWKyF/YRMXtgBbXSbfFCTn+BqUwTXyFgUHjp577Z8tFv
Q/G8VrXctLFnhn2j+eLzpF5E1epQFTtoA3SceygZzlqmoz0ulAj2IlIlOFlP
7nXjmuWK2noTz3+YNn7seUYeXIdfnjgHEM5JgIjaciM3Cl9F9/fPl2ai9XgS
QLDsMFxsIuNA/mqpKls/3ySlbdjc7nZCIzlouMes8yj/J9Fsfi/m5qMpAt4g
gRkbixP3LMq/RqcmooKvxYGQ0Hmuq5GRw0d7Xm8fOvYDG1RmMmJ7f4CISLTi
k+o+J71c5LOgk2sA2a64KWKGFKe9y98YmBRqtx14R2gAx95H3rzdk33WDWE4
oOz5pQxxSzkSiYMZPV038T+LmFBaIoZs3eTJXPijhc2j/7vfrcmKsy3oqvFZ
0wv4U6EQTP1hehHr2ppqJCYosHCRIL/Z177XbKmyI7EGw21ywfauzspJ/P9r
v3OHGp4l0jLLq3A3WauZIoh1qQ2jGTnDpR+MkUHN8iVoC+0z2uo0YFSfQ4r4
sgwwymzvzEWoRnijoNj3YmTbE0G/QGXFnflyDf1w0BJYmSqgvGz40Nai9k8L
I2LJBPr4lzWF4IvmL9FMhKOoR5Kii0I6SJw1gYtgVaiezHefeNKdsMoSQImf
Al7zZwNm6bg2T2ZOLDyW6uodQPAk+WQG/Aqs4dBD9YJiQ41dN+uaZDm1aQnJ
CcG6Tqt1D5rp7fvIkvMbdGWBnm9y6ljNwNx1E7UouGwyc4H6416sVYBADtx4
gWT3v9ElVUMAOhcD84a6nHyfl5lLY6i7iTxgl3CJTPmr1Vr6NF5B/kyxaMKu
kGNWjFYtvenvssf0et/RorBJ6db9gq+syxp1yo5V7JDtxyKjT2gXsvEJ4ST5
beuZzYDtSMG12QPmQSpiTBdfLBOSc33Pfk0ATYBlvB2NSJ/ZuG9O735jP7xo
aG3vwLNL57k5AKNDJo9fzHEuauGvYjOEzX18Y9nF5yQlr0OTBF0k5SNb8IeC
rs9/MRS+bcDH8VUNWp//rGAJ5ttjVayJ21oom3SvD0t+12rOo5TOCcOGw5SP
Df4cm6QsYKd/QLejEepPQEZu+kjifI+fz5lAjmxkrhuEwH6i2x0qRJxEls0k
gsOIVtOYBENCImiulDxuhMX5rgJPa8YxpU6Ycmb4iD21KKH/eWtn5Aq9nBP2
pdC1J0WgiJGkRykT9KurSM/V06b3VjB/lzUu/YPea42UEF3N3w0hQLOVSqX4
K4hy1whGDPZdeG3OVpR69e+Au2OUij9e7sZuevnU+FOIH7petja5UEtfeVUL
2IDTXZqLSl7EcGXTHfeCW03iMFP/f8NeOvRP8UT+lFx5WBNMeAfS9mbmrgWx
m+r82iQPtegbKtWUv1C8LlzxfozSrUIzg6AFhxrj7KG+FR9MzufCYnYvsBvs
tQGr5oxmJYJwE0GA6tYJL9Cxev/LT9WmFkLD1wN1Ff+Bva8kdp5mb5F53y7J
N2YNoHz4v8fso5t9OqPZnb7epq64xqOHBu0pAnIPSqf/PjsdM+aEi7EPTUTW
dXL3G+esRz4OQ9O/6HkkZ8tPrYUv6+EVFssElN+BCZ88qc2j1zBGLn40ZmQO
BPvWjlTCVgSEh4Pbetigp0ujGcpGrXC/kLeTDo3p0cbJ6f3SHQas1LMA6hiX
PWHg5bDxH20BDA941mOFFvjyz6NoSwjPCdMJXXX18VWtKv6Mv3W/e494W4vJ
8yGGaHUNxQfR3NcrOehbrJ3rpE/icC68xXhrFZSmrE2ll7idyWu9MkTMNQi5
37ip4z0EcSI2pNx5IJC0i8w2nr0I5aNfVTVEH/pEZP+etICydWb9ThOatG0q
OEGAdmVklQ7YpYYGtKdXURHrUxFG5xsL1uuPRxLi0AAvsa+Bd//2B9zNwcZ2
e6DsIPHNDUumA++EE7nfZ7NzpdvovPmhdLYQ725AM+AwtRtCTC2OVVUgZXa+
N7NW/JodwbOpUSGDLHEny+Oc6juPYRZPKBm2D9oI/WQp2ABiKoXgauoLiGe8
YQ5jV4lkvPu2H8NKXsyFT8k1uqsXnWcGBi9+OsiqWxgZEhBwe46MmnetUNay
8oXG7hL2J8s1vwMfrxFLkAo4F21RHFPS6i4FCRqH7I4U7uecENiZxwBAqEQu
McOmBseyaPUxN0/KZ9P+nSsCVtAKMIfvk6GQtAMXn1ytncKRWxjLqUmWaawR
PmypEJtzFHb0Sz/Czpdahw1oFPMzHBvYB6Eyb317Y3FGRBMYzSL4mzZVOOno
zsPebI8JeHVS0M0bO8uFKpUYsYXDdPTm2flZauW2x/DEQiTKxqRSG+jw/0O2
kPEo+uDSHyahU9+y1q3acz1l7iODKpxGdW0fpmNymbxoz7xAt/lDX1LU5sXG
8l0D1CZ5BR/TKopH56L8KD1kpO2pcChPnW0bXt2RsJyx6KQq+lrq/l2hMohY
EtxxvtomSCLG7oDN+CC4p6guw1+hSBNzDdG9upGWwkbf3DbYRrlhFKqA2h3R
lNEb0LnbylLyk7ZS1agPPDdEVFnKpGe4VY7X+HFIiUnldlEd3bl9ZSpNsVe8
+n2ICSQiR8HVvrtxjllL573XdEn4clV6GcPMGI9EN/7tDvO9vAF2Rc73BXHZ
aSQnHusu0s4SLSIMT47kCvlxB9Tyr1wzOvrgTB0EPwEJPW3f6+Uvv4rseSSy
uGbBSLvVy8zOt270QFxGQIzZSkgbT7nDAJhhfJWg3geV9GfVKqSSfllFnex9
BmNcyOjUfWec32Pe3PmC/cdgq9qnPk7CBXlYk+Pw6crafu1PxO79DerxryuS
/H+2SY4x3ZEV4Dgp3LGMerw7UEckkVNBHDuAG5QdbYXIMzQ3D4J8BHb/AGtt
kolhBnpHgpn/Er65TQksj+W7cs6/78Ey6fS5ZCIUauCiqjM3cXin5CMZBmug
bFu2IyhKZ7pVVsh+4Y/3J9tuAEypFtR0FHZ9MC2Gb8uzreLn9P4V27TRVh3D
Ga6Rfy4JLBPYITKaSQjk5jx5oowYzum5GhnYyiEER5+820g76HAsm1F9zlf5
xnL+dkCbQjapKUUV99huVSfQHPOM/GlwmI4csWV7ZxNngWFmbHz2MKwolCyb
sgNe+hnZ1NB60YUUrPSLUhZ6763JKq8CIHz7Uyec08jmxF664bsNAzPgCGPA
xlynviZirQE1dxdB8qoKolr4NajFrwlT8lE1g1LYbBB604V6seThdkSAJvKv
C5djZDDQcsf3w+GB+6c7cL+63sDMjG9GFJs4h7R0rbUY5Hdd3mQrj5fvQxsF
I3x8kajhJkp7cqQ1AloIk78gQUgx6hx8dvoeX9OABZwiCFvEuMyeuq0UqW5e
z6cAeGxWaPb3veUXD8BZFdwmYrlwtB/mEpCcVasmb9nPPU4z8Mv223l4/a1y
8rBDwjCl2vGIw1XxLRN6D8oII7S9C7Gn4iAmXTPftUkxMlC6ts4RkwbHn7H9
5azk8lHimaX8FSH/nACFdtUPqGmQQ+DZGdvsKoaF6no7OYPPM7lTfJZfa7dT
9M18YxivZVyGR5NAOq7d+rCZKZDZ7qQI5YAXS81iiG3b/w5YbqdJR1spgUqX
Qwb5LbfyDkly08Cj6llnC3rBkdDVWyJtcfnzEqzQFPuNv7XxfYCcrEr4+WYg
G+xSUaZ2gnUEXaZo9/Whkmlo41upcnKp1syKsKQ/MM7onXjpU5jOlen+P+dK
lNavc9dbPobzPvmzhjs93qKOFXdfWDf0aEITNqGkQrQHzIUhHGb4yEZH897i
hUkXJIffVh72EEsra+mA5u6KBPE/eCDJRjg4ZXez7kCIB75zMa03VU2yxJH6
2yAHojyTU+uEnDyMskLJiRPgUjL1Gh4Qowm3O+R5Zh05hd4MhnCyV3NOaNvc
SKlw5DeM7ck3Kep+R910vCD5d8IZ/GCZUXfYX09tPaGcigZueU2ObE2BhJGu
dtKsWDzazYhP+bmISoTZn613HavIWUAdlsuj5X3XPcW09DsCGjfHSxYP0mfI
BW6pUCnSwb/iVvTUfyGrqVKYB34c5AJnSuqRSLZitdN0q6+GUe1qAQmk4Fa5
KvY485d4YSXYiQy0dCzOkNRgLBSwC9ZbvAjBqGTmpgVg3r5O3u7p0vnNEfi1
6HFdR6GsFMtZ+7KEbGg1Spn3wO4psIPYErL9XA72KI+6hKuhjZ4avc3OpmPo
6gGsDGWSfd/ZRKXuj8kgRTOaqRglLgy2eZIqifxe0N1t1l57JvYfSepy/a31
T6cyOKmkqs9b4MvJGYABn5SEUvAWp/FB0yWrPeGqbMeLGk2UR9VEzi/umZ8b
sLcocL3yYZE21yVCzstmN+u/NTWvd7kSW26smxuQouqAVhnvj7f016ZR+Hwj
yTLcrfVQ2/RueJvzmaIgXmotU4YrUIOGCiMEDlldHQTvNVkPLUsq8zz468OG
glU8yHJ/k4fswWy/iZaBUxB6ZWjeTvEEhjCL+XTVfTuO17vEEFwb/fjtVTse
53NFppzLnVP1HcExF8cXmuMRGtrE4J88y4yQb9inVDtC4wA7AlmlVXwjJvjX
V0o6pVPkBybIZQiF6bLtu4W2YdRb53ssHGS6H9tplMXGkeO2dqeWlL9OHMTN
DsMFxxQnegPvP/uqifNgqYBEMGLutkfS+KK25PhZK7Wd56Dl7NGf+uAni1Tw
OSG2AEcVqJ63NOIdjgnjrWz3p43ep0dzkVN4mQVEL6WYkNhwDdq1ydKxblNY
bfwyBJiMTBCdMaV7dhtNDggmlUkTEFVwxYkOi9vhrR0JsX4Tz9mveWsWHqRa
wg4o5bL79uMO4y0Q/RsCpv3k4sxfkzcuB5/rHRaQye0s26oDCM591udVMirp
wFLxT22cIlmjWR99FKzSxEBg48U8q3+9mU4idQb2MpSbi4a5ZHpHjOI8FLmD
rQ0mLt3SCBrOC0lbunfNXh+E/dacDwCcsYPJD1AMY3b+LXcbw3d2Wkm4OKN2
YOuxCPDObYfB5MSCpKMtDfYjbZjKv7JxLL1RtuIgJvhDYMhkwfTOAk4PxqBG
HnFeavQUma5TKruTHYq0WUakyRyWYrkYzc5sjuIj7qIYotYyTZtQr7FtpNQq
xy336UYnvLnOScx+WsI9cR7mDoki7Eoe3XocU8ISyxpdoymzlgCbzYvO1jiA
TMEe8D/MNOWnToFq51wx7yasE48bFTORMa0fC3NtuBSKPJuRY5D9X4YQozBq
Sk/OunG6y4RpdU9A/HyUTHXnxdKOS6qSI0aISQiUqtSERqxcy1FoJq5B0i0Y
Dcc+2Bh3lwNzvBJ24NTRXGNl3DV9VGXPhmfjRRhzLg4wn6diLdqQ83Cnjrhw
MrufkmL2eLT/QkAvzxPCmBo4ZnE5oI8YB3QY+LvSNjscI7hICsVGFTJ5/gzb
MNFDYDlBUFKSSh8n+mt0vFuZGQbDoHrVhMO+3CAA0evMfg6uSnBAINkRC11R
cUgkIEIYXvg334jF9XS1ozn9JXKwM6J9l5gh/+b6sS8yk1ehXzYtKifT518D
PcZLbY6+D12kkritVwzTeh9kkvQGLdHpqZrzQ5QBFv5AOmrrQpPuH3cR6W6P
s2TJVZFf1Q+cgkG1kvS8XFXF7g1vd1BBrvPnzrlU9c1ARkVxXoBSG4MaaKPZ
j5iyvIp1e7TjipwGwuxl/plMIofR08NIyhIyi4EX8Z77/noyeUQgT5PDk+Pu
v75QmLs20+jn3S5ZZ9rR+IkqJoEMLl1cFgLVexp3fz/xZUb61AE1PtCp5Zfa
Jb69DTch+nPvzFz6G+tblgUbi0vZhKL1RCkmMmJDj8dpG1gMbofHjk0xmnI2
/IH5nbNyfL0cbXsmF/geLJgdMxpDnsCoxeMuHG4nuhse7QRdI+hYHg7g2kt7
byzf3a7pTLsvmxoMW7rLJiDMX6UZxET9NIikonqtJAGu7cP6tiP7OO4G7Dan
NLQydCjgLB47Ml9HQMGmRoesgrPE1mgG8Zlxs6WHQBm3ZNbX+xsVuv5ESCi8
d/nbKCfFHIR1eTA3lFdsKSiAjApAzhjl4RqFfAja6FymAQdjjRY0rN0bcGLt
zvPXCLxt1h92Yp1UtSSIquoZgwXrAo0kNQrFgNBqo3l1QehQMjar72R87Jdn
0FABDycr+wPypzi5PW1uYVhJY7/5xRC9higWVLYpRVfLCROxPHxA5fw9ucKM
TRqJ9ECNTTvKl2FPP2f4y2aHtRPj5bX43tlOt5iQb8Iq3ranTB40HiUStQMa
RYt/m9PQREU0UfsutEb73BQMOpCmRnTQTxvDdkGheb25CPduxOxLeofKdjv2
Fk7cR3xFKLqd24JSNuiqbhJISV7m88EKVaZEwRC5M9+sPiI9ZPfD6Wf+1TEn
bfCkbVkvLxkS+u93vuk9RXszK5ePxj8EcGvhcfwsr6vTMU6/xQ0q/dq9RsNy
XO1kYBQUmBX7qs0qMfU5HlhEiF/Cg1xieI2CSku/dnD31LgzpdNazd1n7k5i
o9VI1aIliXGtrpjSOP5qLZSS3/uixAgJLCultk8K7K1iMWJOxzmLfEtfgCUU
TZozXCLfEZXbHfzzEg3kscDhVn2b9MbU5190f6IcPwJ7dXX+/LrujJE1o+fk
Ko/PLpvvHpOB8STU3dAqTFN5zgn9S+luCULtCeL7MYvdRgscVZGhTYPbVi1i
fm/Z3BaQatjKGXe2eUj/kp67z6999ZeqjOnQU6+pJ3uQD6S7avzmuuVs775d
+ZjGEzRF+JpTPpCXE456hGmVbu4uD08v6wLUGxXMes3zKI4Q0BsKQ+ansS7j
/bDVBnRRoQT116I6lUrsEGHQRloP6BOBbghCDBGOZs7yirIlxAu6qrrr0CpW
CMA6GkzMCctFerpckH2RHDrsIz57KwUldjuyTdrupEtF7APZ4srTi5ii7o6E
BzQJ4rjDwSIZa+kN52J6c5hxLbXUuiPLrKvzImHdfGYj75EJG6gjmg2NSDba
XtkhuJpLLlfyHcZ+9spv6NsxuArpXctf4KVpoAMQ4Hnc9785bGHjKzZRwknA
x1op0xj9bFgdPN3KUrqZxVqIg65qv2gdjNvXO3kFU5paZbgbA4ngvi7IUjTe
7lOvSn2/LNdqIJ5eiZZUFVGuCftZet4c3OAJwMAmFImQGFX/FIyzPI3PKzHF
bWIN2QAkBqGwgyyBL0GaUZMSayVzKizjUcMmgfmQ881pjbQ4HYYRY2hvs3EA
jDRuY4zDI5IMDP7csRoLeLkb2VdY/xUenIXBZ9X7DM1xpqt2Pcr8KT5GOZ60
xWrRY80P8UNBwsUXEiRyq+aVRX1C5k9TWDNoJgxcFUS2dHO7RQzjTAvvYWuJ
IhLpeX3bAd82F1wF3kbaVxln4m/Nk41oxGqikpQlDIT4TxDaY0B1qu407lRS
zIEkl1jYb7xO0N+UZ0NMwg9K4aDs3R43//KtbL1UM8p1qcPqPIKOOGxsyMRI
QegbTwu33k6RIPDLf41Wd418ZgshvveWyDvOjl5pqCC2kjj1ZirXuUWFyB7B
y9CknMRysgCH/WPPzRtsDXyHXq+hbnPOjgpc9Be1sNYLbF/p9tv//SYX20V9
8ErNWU5kJAHXxQF3DCHNWK0F4qdeIlLCE5dRb9y0UOD55Ib1FfY4cwHwKWAv
mlhbwIHR36pl1O3hJfUDupl57CH2ShzYoqGbsa5plDB+1gMT9MyVspgeH1a1
BqmTDDGBeF1WOwUNDhRpiyYKINDMEz2UQf4tDAMMbDqsxzr/w/2zLivkDJhx
2pLvzrEhXEweLe7l4wh3u2fBXJGWS1qVq1GglkVBrckV7GKB7t19J5O4lkbw
HanxK1s4QBIYfMJDQH7Dj0e7/ywPtiNfiFvsBx/vtvhgVQGc2vLP0hewjWGB
86gNFxbNDNkRdTtAvh3fRCiaQzaxbH3oY7S42+dRZatNGRssS93B15IfEE5N
oRESscm4UcJaYf2Y75ik/AWX+pxMN5YdLU3L18cgVaGt5Ixd2CFm6CI9vXKd
u8pBN4UQq/EGpS+fR1MfwoJpYSayNBDSYxaIWiy6kt3VNCa+cdMjaJdSNYH9
JcHAUA5+sa0p2JQkltlpGP6Oo2DgzefqfkpFjf4so72aa9Cq50NMpRRT0Azh
iuKulqD8p2nsMTYRlyZ3dXq3ol2paCSNTzk79MbsbDyow6sf5kf6LScaoPo5
lHyIFpnintGYnk8DHQO895r9uS6HE00uRGEeezjya9q3RY2T9rcYLzxjlSIz
ajBDA4U2BWgL70c/R0KoRjiN2SghjhypcPK82y5BBjNtO+OUbrot1q60qVK1
QzmJfh9TO1buRo4Mx9o9bDiE+P7QCUY78iZ29tGGekr7ATQcPAwztd85tVO+
EI3tzDc441kdSrBbK2XkEPUVoQXyUJtWL1DojWnLVfgvDWCndLsi5e4gYsad
tkzFXwRc3nlbHwpiGBNnU7Y8ze9AntcRAMHKhoTNR9IDrh8CV3AXW1i/5aNy
V5bn2xt00gIOtGYWIJC8yVhEaCLzyXSr2/XRZ1Bt+ylCSlDfH25W7mkxIRKX
6+YeoZ3GWwjvsp2MR97eNlKhB8WtiUsqfRS+J/8fD7VCYzAvNfOHPTHRS6pJ
YH1AcHc20eCxVnBLYiYC5JG2bKpR1PXjExgAOhGfH+QHBV477RD6vqUuw00e
vsxeJOBNshLyNgIopiVOiHjcaqaBl69g1vbFcpjfVldYRBjEDBWUIUPEhwao
PyV9DZ6AiVRt9zDL0eXs5WlJ+vHeZtpmwMYLZAVJSxB9WPHkIPUgZE6iY2uE
nTn7Y9ULzq+C1ioVIXU8l2NIH/y5U4od4FWSLqSvaiEj79Otc1zJ+mQ/h68R
A+BUsAbIz3Qr03uZj33lO+pFTH7vc5Vkx/qCReprN5lIf91UhcwJIoE797TF
AE3ohXMsajvPg3An53Q46FgWBBDhmTViQNBohNTtv5XHyJTJKu3En4MvmXiE
ece0TuoA8PGhZDyBgJpjIoUgJid477Vpv5BVgsp5WJDdQG/M19pBKFI93rkg
wGa19U55KbecOtQlLOkHONERf1Bktlfqag3aD4rEhAVJQ2busWD6MKtZSUUo
NidkE4EG1izXSunCejbmo1yFWSmjsb6s5zzgWR49IlS66V7EKDtZJvrOjuox
3VA+TqEhdnZYbf0+a+6/wDqoUT12Yl7lXe7JisGeEj2CWPhsdOphdv4j0HYO
MLD/WARVXq/31o6gZAXHhoUd67x4cr/x8jLAt89C1f7SOvZyr2CR/bioXgKv
1DqzfSFiYBj6FHLMWR+TSs5jluFUUrP8tIemwp2JPbrj+tow75UBdSYBxCFK
xS/biRhlpvPbl0CoVVZjLfcENKAx8mC73GzNMs83Fnk7/37TRg761qR5AXEY
dcTf/dk37x0EXZd5zvKwR1y1OLdZnZnVg0cm2qOcNk1D4LEBlo+fM4NOxh69
fqNymes/IrN7/y2Mo4DuWI3BdEnxHiQ5xVoLhDgjX7uWxXy8RBNonTXyFeFQ
W7w1MQNGDy2uZm/T6avikz74HBVjbjy846QW32XkgRAjbzSlDQ8gIFOK2hXI
P+Y417wQgpJybKqc8/hJ/z0/e4WfD3YYq+7WhFNu8uWNyMefYzEB9MmszwnV
Q/V2/whTpDd9qUtJ6QgYYV60VoIm4szso3+7licFMQRecAulsRjFbL3QfNVV
a8y0ovchJ0BNaSH3+v4b2028uAZLE147qfdsfh3a0vVGTpCqp0rJSSj1i+sU
3iWL3PqPkU58Ex5Rq0+S5hdEjJY4cIOSMKcfmWTmIEkXMYXG0ZlCFgy3vzjl
lUye2w4cz2Lqxs0jYmn1NhHET5KaAonOqi9HfSUzMRDkMnTdZ89RDWapqVeq
yNaG1g1eeXTj6A4KUuuU1aLye2BVah0851E7bnVQE04JsNbtlRoCWSHuj/Wb
YsSEufTnyunOptQA/9fYdFY5Sx0kzVZq/y338BuuwbD+ge7nIDXq1R/9Wf1/
WY7sHIHN5Qcoq+vy+LPQ2SXNyjKrfJvRkaZlQjjSGJtxG/VHU/C8/hUeRWb3
oriN+1u0VnfUQca7VJMbBImW7Sim/yyIj35mF2nquu/IOd1azM6f5/0t/jW9
Q+Dkb09v4EbJAgn2nY4RzYlxleydkgbFsvI648cYjFWIlEsrujiF2HbWuQLJ
gD8C8WGZ29JAmVmcN29RTzV7TT5+RALUCjQBjCbka4lnzU+N5UsRNPLNXDpQ
gBn9NDfD955b07cPOgzOrjs7wWJR7ObAqQPevwiNh50OOUrlnkk0xVRQTpJB
/3GCvq8OjCa/MjfWW2PZgj+d0xk6gZCjU+yYI+bNODFqOfu3YxtE8IYsiT/p
4U21yGVkWIh2R6JtMPlTzKUXTtU9zI8K1ndlidpIKqta8OzEkUr4Nyt45Lu1
wPyOBaMsXDr7f/Vszo9/H1ZWORn4MyWXZ2lYUEVIH+y5dC4ZFzkhEar9L4xU
Dv8PEYafnV6H1sVH9Ep4wEbkhqUm3ykjjDlDa18kxHCc0i5ZkSMR7q5GGzFW
txO2wTHRR628JNHCB65u6S9oT0iny3vPKQxww/kYjRL0SiKYoWtf+LDES+qz
ku2D40ACIhi/hGumy8dBJk4slngv/TbmBQzBPMSuq21AT/jdAly/mvesc61L
Qfsom1EStY8kkwbOVnPt6EBL2zKfoo8s2UNRqDXLQWe1TKJvlidm8k5ROZIz
jG9sVE493pTOsTsURC8I21lelF3+KNUc4XmiTUuz4IbBi0UKg02e6oV+sx6D
ro/N02kOEkHKpuLAZ99kOpCVYDnKcB6XlaJlfIeNEk29vdk4JrShfO6YtNpr
hC9Q8PKV3KJBhIPJTwJ6KvqHiHhh/+lGJSpiG//o7CqUqs47GvWOT/DWVz38
0nZc7lGdhrOJ08vs+mR4k503MhgRlCOJO+nqpSPC1sbomuNBP9Qn0YHnbpKg
jie9P/2iW09lO+rw91ipF9Xxjd/ClJYyrvYpsSp6nsoPzAmGC0LI0JglaMii
+nh5qzPQl1slllsDpI1zbrWZ61kN6qQ9KrwC+HJh1mgs0jDlRajef58AO8WW
fHm95mOjaTVJaExbW8/+nr13i2ZisghxPWrj4fmLVNLvj2g1kdiNbO8sl0LC
X+e0LJMQzLo0gYavdRadlHPo8D9Eysvf+zSXdbtQm+rF9VUZyNkHooKsCaNX
Lo4/2lU4HqKtJzRsBFOdVYXfqH45pGP2txqUBQGQtjK6g2JVk+eP7QUMMxZw
Hh38ktCi4Zs7f087X7t0EmlX7dTKlQlCIY8kkPf1HDwcFsEIF1+c9moc27qy
lX/WOuJTDeEuYobRjc03Q9Zj3/NRbPRjTGOFx6zNHuCdQ72sIwF1u761d0Rz
l2SodzibgJEdTgDgMTCvCQms1iuYbQ9D31NldjTLH83zaK2B5ryPPzfoN47l
5BuJvFO66+ImftPByDUiCny9tJT6corbU12gDsbDhxNHVzy3Mek8kGsVudW3
tACu2457/8HSvz0CVMfZZeA+TcV6RYVWnZKWic0lpYQAaa9H/BFzSZq53Szy
6Cb7S3sbR8kBE1Vfkl8VqXMPNGML6sTpgEhTwgOwRwGwP8LeCxQeMlGz13hp
uaHyPyGxAFqo1ETD93kNb8xYnvNRiCTwFKtlkZi9HFGmrI+S8qLABD0Cplss
1w2P+AJalmKB7ZgSJpsVshvpazUbLMwrHJr4zDwM0jc4/Q2yNub73PE76MGq
4OAHFJAgzvtkupdiz4quevoVFZ/fA1FkNrsrzpeRWciYP4COTOtKVIHY7dsU
6CZPW8WuaSkByNbge0wyjpE33xbY6HxyDDdQzeKYRbIqceJseChLVZuhtMgM
vOBlIaHyFrAcvTghkoLCJ41SHgKPzoV9BFcCH5eHMJlj7L34DLChXeIV1SvK
6cLMasxfA6qzv6ERvmtREQseA/+GNx/TCD8Iezvsi4FZ988p0g95IjpLBZIa
gwBVIQH2jig8zgct49bncEq54UkpDor8Zv8jsObJPSgsIszgysC6GxyCqFQg
BCIYxCKjrgYKHsOwK2/fPayTY3c+5a09MAWAsR1wfhXD2i4HEAYAjmsSN05y
+bxv9lORZs8ngCyb45OFXciOikN3E2E/uVadg/y1hPwHFS22hQ013CEhLqIH
DwbvEbftq/bmXuQy8EJZ0jYsQVFRpa7HqBUSzpBX5r2S84nMJ2S0kMoViHBG
j30ccNO/3/ocOnnhEwBqR1KQwvZ9LBDkptKR8AU/9wZ09bmU8DyDnjsJGnD6
3ZtPVRQxxRW+nv9qw+xma8BfCkJ6LGZpFLwkXQ0Ymgqj5/4elYx2S1rWi5OW
36pFzcixy5Uekh6PLGqh293ZTXL0Mrn/RMzgejOZMeN/cBs1eVZoQltH/R+i
5SimuOsfAJOLPsC2rOHFy1ZNc9u0uZgak+CtcrqQYN+jJw0ru/mUFFG8yEC+
GnBFNiSMaevPWMV/f4Dn8m2CmOe5Mb6d3mVVxgIAIO8DATQ1oWtLkbuH+eet
J7knEf+cf9ezPUNTmN+H1Hk5PIWwHZgjHjCA5UlCfKwwzjXvcuOP6P3NmDn/
A7bMvANh729G2chpws8srf/B4vFOvq0fQ8pC1jIuPpq/mPuwCrXB7vLC+LFw
5qJ2p3ph8bOR/J8Zl7T7ASnSjQmy4MmpFyAc3A1O1fEcAbG8YArc4BEE23Ga
RLgMxxUQP8MqHZtAaXTNIie753rSzUc7L7Cw0Aiq5H4WhBzQHbZjUd+SXmaT
TJvzLI9pnhfIpTJPAPgJLVpeyqIXKjD3DOcP7bCn1bk2RwjhFPJ/Hq682y+i
6z4RBXV2wHRPrJ4S+yNjv72v+6ANv3nHgJpl8/pyJIaQVFib/e49zPhfV3wp
6njUJq9b/IeqWtT8mQUzsaQXSBfPaLGzZdbQ+A3MqRMTfZ9uL+PVj+fVud4l
cF6gIx/zwaMVYdVFYTJQwFW7EN8Tym6NstZEwlbSsYA0Www3Qfnuhu+UA242
AWy2I2LaezwF9TWa53ig0gxryoogSO1YIV8EASxzGE7jR7wxhpISAVMzsXLt
dO4pdipSkpzAx833Kt0Szy4pX5WInAQbQNWbe43FQLdCcxOmzMNx4+vfi+q9
9bB5vdLDHjfJ9dP/FBeBLHTHKeIBGZbMeddI2YbgnE2y5h8MUHtPJqceTVlm
eM3A87jBi7UozeGc93MaxGtwUo2KT0g3/6tCbFwdsRKDrV5h4FWTdrLzihgK
cyPP842CU57O7qeP7ody9W4uqJx36wBae2gg81+ummnYNPDFmnX5dXZOWsYN
0C9MXJ7wyFPc6+t3DS7grsO0aB2c4FjOy/p/yXczVNGbrx4V4N7M5jX5yaMH
0Ueh0YnG8iqVoNhJdfii5somhVMPqLbjXuOdcrX0bhV0CuAJKEikHOiiw691
GtOVo6Nmr1731UJ1f8YxiRmqlWaSYFejILS9rfcDk3PTncvxVGWst1RPXESc
jXeqFSFOE6xdN6Rdka7zxOBOl9pgfn17HaWlZbOjCsArhAfBrcWuuVnKg7t1
1wU2mCErcqPr+yWf2/S25MFrgzIh1Vxp7FWwhcuo3ORiSKZzynmSEbaOMQXk
vip9gzS4mTGDa6qMVTVgxgJWwkMvxt+SO2nLjB90PFfAm0vv4fGyyFon/nzw
wDGeD2+HyQlnJPewCphizcdoc+b6SdE0LvSpGyl810rCp4/vZb44IhWGwVch
7s9NaEnLH4+UeCQo0WF7IkIAgKBc7qJBvFLrijA3tK4eif4CpwGrsQ+M0KOG
L2xr1D7y5kN3ZgLWpT+d2t5NAwHpBSVXBFcS9qBEI9ahOm4UC9KzfMeskszc
oV5lie8bZmBKOBwe6OZx8M+3k/FkVWwvfydk8wyfHpQA4YuYezMYEYITGkeQ
oAByYFOOlzOoDPoqINcOGnQ+bt2/GJzFkXifqwMm3y5GM6UTVvqjo/HN3WRw
Q01IsB9WSaIQxayM57eZwxatGgvynSzJOulTF8juBD7uzbn7qpcbdnxfynID
akrfFOUImVqmrjtbdoYKK8k8Zw+15I4FiPwlWX4gBphTrLQEO1EcMIlOyCje
j8h/qoNclh4u4dU/M81SC/dUDTMlncCg0A2jRV2u3ClJ2vrxBGGp0axM1y4u
tb+vvFAEDETwog2KI+mEOl6r6T2UeEIgZmzOWENaaX26kAetQZwAeBGdOA3L
yaI+zUgGSE0bpnMX3HvyFk+woYE2K9zEtWyrNZOmChlOAxqT80JW8StYxHEG
AWbSsWb7l3ZQYlBh6+i+6tN/7zGhRdjI73gvBBuN/EbxYhxROdHVmQseesR4
ln8ety+VbvMutbknhe+uM74Mkm8OUEihinl9sO7w950u9cggBjYtIeZwPnXK
4I4COKBZ/+JoqdSzdmNUXdh2SG9z6YFd1yPD0xWLTos8OfUxFfoKFY54hs0J
B1RMdLzTf04JXfGjrJXwSaiyC7qzJ6hWe8pi0YZWeTTeQ3x12tdpyzEbzDJc
IvFMk5sYctTMvP/xTxJ/k7aGshi+YUIfIN0g3sB604oVUIWlhVkn+L3dF4pa
JitR6WKnb/6xhnhlUzCvbZIf7LJXHDJdmGdG6BDzp8oqO6io3CSyKb80/s8e
oHMn3/judF0dZoPcIMWTCteKRE3ihX4zfmfsiv+DeI8yppf/XZ0KB2JAKFyy
2BobP8Vn1xS88ms3H4lw0IPVWiVcuJwWBhLYeF+mKjNGPqi4FcslRlkVEgAE
mqwbdX294BWAOefS70aGs0hHILgNbHu8PL90PrE4mF6PvgCbAcW+3cesimpz
Hbg9n4KMluaThodP2T1lBuHgLo5nUQlCWsl7wLhVCVClqq4HB/dYFZKJSdk6
EE7/vrvPFmgHhKFUhZZPP9nDqnkOLXnlzR54eKqBPO8xLHYjuHGdX5s/y04Q
C5ALBTwNhdQIJk6f6p40mQFKs0yEWS/WrrksF4w4e28CMGqZuS19AWnR+O6X
fYemTFuicpPKVsRXwMUzyM6eFfq1f8cYWdNtjall008TvbRNxCFVzVIWNjFT
LFdb8iskzf1BBm9wdxA7vxY+L5vHLlHDSGmP6/aCA9nxw+cFsMkNf4VKjESS
Va1axT2i6ZKH2XQe6h5atyhr08TxnlahDSZRfNii1wluT1oOcn0igSa75Y7g
Oas7l2iDKG4rpBo+6T0BLnINaOS45CKsXZIT3d9qXJZJMTEr8O1sMuFtqMHD
biECYsg/4ITRYMFhgT07CgK4HqDzvk/Rpo88Fx/vW2cS2WFH1tte22IjNGIj
NBVN3iirpk8/Kp1C6MGJ9sCQHtr/woqD5HHBwVSsdD1txjPxlQMcBl9139MJ
VDsQPI5PzO0ftv2vtJVONHZPiF6p2ZKX1vOcexHZPMkWd5aO7XXR/WHbCuxa
DdfmTBxUxOQ19g7ja7ctlloJAOm61jpImpGh/4hhBbjENe9uugBi0pOD8LB7
O0LSML+qSPZ0ckyxMzsvasrv4R7jEjEih0kBc3biilNsqZ4/jGn/2A3NwlxW
rTFSW8E/LUVoNwZi3x2TJN45Ec50BOpHOZVZL5md0+qXcdS3viyndR00IfzD
lxCX0vGq9MyCSXG8RVKZ8kGAU8LsUI30f4mxeFdp0S7/1e1xQmSxyfI97PCW
jfXRu8saYIxdkz4nVjSmAXLlP9qNAUayRkGYn6Y6SDKN1DR40ce9fd1GKMhq
pFGsN/kLXPN374TApfG7Uff5/zR/OMNU5G9gXHg1M+2afVsQdU1DCS6/zf8y
reGk4iFRZNuyl9zaSh62X5x3fiZ/DXZzfWDjqFsVV/CY5VHGVoGj4NSSvds4
bG3JP2RX7OKMaW03TVGWk5kQhJV1qhkOnw82s1x+aIPPWQZnRiC0Q0sH4Bws
Cdal8r2mXUVQNfDhuLtbUlEF4jEPAVRSEh4br5nLlFTC2Ui7eiUJ2C4g6XRf
/mhkNRN4/IylhpVzXWGElJcvv6qEkFw2qpn86M2Il1bZW0js2I+O05lwDSyO
wiH8NRcywg6SaUOSNETxCZ88gIoVjyuyiA8G6QEQAwfRLNNs3TKNq0jLkwLI
j9haRVWO9lza6jiKL8EpuruWfbElDuHX0pug4GlpXxRd05lD+tV29Obwn4vy
nr4yHvV8UXgXgwMDdJ7QIy2e2ntEHYEKWgZP+G9A/VdWJg8ogFeLEk0XpEfQ
2/YJSLAdmLtEdlloBHgDCtgFJWMnPFrdN52vbnpcmmI42KvBrDvfLxMiNpUa
sym/ZpDSkzf4oHzcIWhs94Sn02eSaXL6cMyaK9hdH+zTI7sTxhU5xm0k1xeM
U1dQzcX0UGXXwK7EEo/YfiCDoIxNCzw+/W9JmhZEzwYgyW/B/0pOES3ukoD7
MXjiN3amY1ClOJ27u8F/blzp/L8/h/6PuOSb9KYgOGVWFz0f2vMEEGYrIzIT
njdC5p+xqfXvaTwb3WB7u1STC0tJKtIVOYS80pnBLPK2SzL/kVe4M0UXfwP9
ypqa/5kLPBuWtrGsIp6ki9+NA57PRb3sca69f+OFFpH/7OMEgFz+ZAWxz3F3
LALxYw+z+jaDN/mcYjgAzWNu+LfSgsfVODNwY/ZhSP7adFJ/LQRex3fGZqYc
IIs1fkffOlhh+5tm69MURqHETSNKROb9MaLXe3s5oM3FX/oeKL58izt4Lh45
XejCigyUcBe4JxRUK1kwQ7I8uH6SQ5fA7138u22B7QAjDqDZMnCxwX9PHqLt
G8ur+OL5hXE2fJxEoTa0uH10J6+Rian8ZaH/ZMbaWOeeSGIjDtnt/VI9H1GF
zvcEIIoBU0TjObbYCbdFogdToe8KrztK0o6RtnPOHnM6qQm9ll4oj82E90VB
yu5IHlzd87CBcjRixkV6JHS2VVqz4tQ6a3C2mj+Pj2pPssRRzpIYVwVbyo8c
18Gpre9dxbj1/0S7vR6TswwyLOa4dFlWU6DNwLH9VLHbwwP3MWottSYGbhYd
HOi/ycn+x1ml/m9uXj9VLVxhvjWzQGvRZX3Ml2L/kzYKtbGUxbqLCvY21NFb
WjTxKfDfqE2mUXtgylkQkEbv2bKvmJX24yqlnhGj1Y4AN/tTDj9rR1Kcl52l
TR11XRiRcHxrwB4gEl15MaXFz57t3f/jZMqPBVC1/CII45s81Xd1dSV6NvKM
nfJLoAr/9yp0YyKQbHmY+pq3KFl8hKRL4KjIlptOHDdxwAbCfEPLet2TY+YJ
ShI8E70XbKZQ7RK7XUpiW2b781Lr0rHz1Uszna0K/R89i5O6hhhb9Lp1VGuQ
V5wXSYH/DLXx6FwVXTsLsC8LiUhwZvHz0cttpx5MDBSRiBxfJiijqsR3CiWP
nzC33M6Wlo4JUK7g057+gZUKd4LcheB1T7tDh+YV/OTggR21LSSdAqmgO5Ju
VzYuMHxSXaVfMIFatnwfNUucRO4XZzlQoD7K5g8D1HDuhUZlwzHt+vvq8oSL
Yy0fA7oKTlDy6o0uXRNNxG8HtY7UdaLBr0+SkQWsC5Kpurfe2QIhX69JEjhG
PFbqlSebQteFhkxsEkbnQ8uf9yHXYuMCoDM0/KrHLZrc7vl+Ljz2fTBz0P0H
UeVxVej2SFnlDOVN9ZM9u0HOro1mNcInn9uIz5/JMNzHQ9GVQsnTJIdjJppo
rEDbP6g2UXz3VXa4ALHEioDuKMkWTlWWCmCcVjthWVYDN6dFbFXqhSPJ1ghP
LnTKk+e1ilcrxXqG7mdDsEWSshl4HCGp5ZIxS+RlBZw91Qoga2m0qLBfsYZR
Yw0a/d7s3QmD6o9mRElPQ4/zKB1u/2QFCNrvSx40koiKGQpZgEnDZszkqH7N
0q0CzGz+StDwyFAyLdngBP3xcOXcNCosZFvtbv70/s3WYObq3TNSvHbxsq8F
nZa25fhtJXv3iY/BLFCSjDafgKMsHH5OKW7R0qt78zeO0BoY1Z/vrGE84+D/
jV2snSWPRuuVjnCF04XlPu8fyH7GOca5P0XsRmT90XbNsI/ZKsotQiTRMF7h
+5yWcU3y1Mqy7781ry5GlQBtRf23LKHFc51eKooXSysv4m7WcPS66T+IN7rz
zdzjeM6Q4WrpJ0wYIgIWzyh9PEZJIDg6nmfhSMoNwPNqt3o3U3WX7SN0lzAd
e3Y9dJucRNqFJR2qvFOpKbK9fYG2ccHhmKf1eYW1aj42Me0cPnVRiLXEhidy
rRI2oME0OYYvCrYCC4Dx1ueQ1o/Hg1Ay63X6T4VAsDn69Ut1jiWzrNqBEInD
9bApfAR+4p5lnDU5wGG2yYeSIbv0bSQxVy52ZGZWAajmMe9rgDRYaLRPjUqq
6OI90+np6rUUrwkpkDXCwod9X9F6fvoglYJgepKeoBqxgeQBxew5bZ2LUCyp
vGv+efC4x/ozXxoQnQqhYZkZsAP7lri/14/MZg3tVn1jPJvyZ217xUTISIBR
Tn+zz/jEBFinL67dFNdT4ze+pqcbTbYm0zlAWPC41zMmW0N4zTwLC8303ZML
BulAHSb1uPVt/Mg4Y//0yAu1B5UCtb7sNiAX10hBlT9XCB0bfbZeNMUu4vvA
Q170tfdJjZVDp5NWZVS/gGQ39Ogk3v2jjNmYfgGutUq+qjlkYE0672xdnEPn
scCJ/qfJdOadJt+y3FnUnr7qvlgq9RkSb+9XUNudkUtntV3/AnvzFg7Gcf3I
Pl/kRoR5Ies9pOA9rQ+xcaZf0mucsduB7atiy2szqmBS9JvZ46jyl23hGse/
buGsl15DThSK6NQPANRQ56p6f6jsQenoI3sER0NuyXX6V8D4UB5zThhtpy96
CTA3dJ4ewAcuZQhTpmb8dwXwRg0gyc6p0k9XcG5VYy6Mw0YuXFLaGybnG7fC
H6T5cZgWHjhAHrZ5O4vN4kuAg0d5BvI0C0Vl3HAywMG/JFuTUKwF+k2ayuEY
I65/Nbw8yIvHqpoyFLFHCycpvx3OLQaPapw++zGrMAVL0VkQ6tVSOT54mU4n
eKOvn0vZbDpSLwhdA/K8XB83YLHgBisdpPAUW5yiCGIo0GE6rAirQBJzTLKA
+YxqZSU/j1qVc4O5hxYhmnFqpnKt38nANBNPUzEHXORMlEX+hsbVBgQxLPY8
ewieamYuSrIU7eAk1Lk6F7H3lw7X02vRhyAN7YNMLbJnaE7FaI9ARKyhW0at
lijlNC1A+CJlmptINDJihJf9+2XYDNZAAvJ08gNQf2owU1j8Pfr8t+eVQG7K
fMELVt8umjVF3CG5ZinRbtEKvr+fOUeFdKZILkRLQjH4YpDxJiT6stW65j9i
J1oTVlHkpyClXU6O4MmQV+C4SEYYGv8rNm0dIIdDowRM1+I3MGsyaK23tUyR
l7Q/FIQMZRBQaqvSNJufcijnkBfdvTQcXXt/AZJoj7yWwN7XBCRiixd0w8K/
b6ES4SXwQIb2j237uxR22Rj5XeKbkTb0DclboRCuW2Iqxb6igV2q5fgTKT0j
i+f59e/gvq7mWOjnwLUMdi4nTOyccxLG5qMVPoeZd18e10Gc0BmIIpTUWbad
ed8ijis0Swjgatb4jVL/Jz/Gk6VWKIj/Rcd1tBq06YE4CDPh1m2yrwZfmawF
B3J87I9K6aN3naL0PS4GpejLrrL55tEATZAVVaDVzXtRvWcDFzk4mbObrtkb
UPOxPKbJbAOBcIu+Wew/sB7aplkymLqJmR4Tzjkj1Qf/r8O9IjA9cUNTFg7h
p9yJ9LvuagqkdD7nUy00W0m0I2pCP9FvdqoPUh/YxG/PKaLPre71mGmT4rhh
OMjZanXF0wRajwC804CaONvxnaEMcoJZqlnfIzzEvzxKdmdyiR5jFP7o0QUy
s+L+WdxWsF/YmAANtTsMU3gBUElsP8EFsOzfR0HjsF9ENf81mKxNsFbrAIIk
ytJAzly9681OW0r7J7H+tWbOAclk0G7GEDT5A8oQImZbJMgFbqzggJqPkXM3
aOGJKytB4obpUWcFEaCHNwT7Led/l2NoysQpqoNjF9JMPd3fCeFz54i8FzGs
QaC+7JYvONSzRILnxlx12QAkl7zPVbvnTzMmFjDTa3KEZlvuHAiNmWqtWQkl
MOU/udPOY+DGQ9/Ijr7Zt1YKbol6KdPWAPvuZc4znFi7Zx27LsLJNOeKb1GZ
BwVgBH4uQkzQDqkjesoTMmR1apoF3AABFwNhGryLQAwprSdJ3dOYyL2qOGN7
B26Se/pM1pMEl0YSlBMeaVkhcnIMPuBCKJJFmQlvOqJOOICK7KxNOqGtpGs9
Ee1Hocd0y3KBx7NpH1keT1UxIaJYVzoTl0TTsxjpo5m7ATirB/JZas4X6ghd
bfGvO9C5qFRmv17Mafj1jQ32e26zuiRh2XatJWusoPEZpef7cxm65FCKFLkx
o8ZNdthhq2pE71x1pWbQhSWm6VUxVSQgbGZrMzCL/wLy6ukJC84Wx92tYGuj
4wVKhA8aciK4kaM8ETKoB4m4a4hMacycvNxcZmnZQsrKzh7S12Z4blcgvwAq
cdTDISmxAVF1MbIaj1M4wimF3T4AZCx0RFdIaYXN1UWj0RdSjIITk6dI3RnQ
xfz9vJ5MqoU7pqg86pE3+pi3HVJH3V1U9UxxVv9BMXCka5iWDnGph4zGnE0/
o8ihz09qSpyb6lPwv+4M6FmcdjOtyv6fK2hvgn+6vpKArYL0s7Jmx7mJtf9U
NiBgeXBt2GnEJT+F/JCNcJGNZ/bs+GWaDyNw8VGBNXPcoMYvry1VVLQ4NvaF
5teVqsCRe3t7IxTIG90DmXczkdpuiV+AHNrGf1ijNbi23a7fi30gnXJS3S9l
2pKjQTKFkmvtACuyUFKzLuKy4nl2jX7dtmzZWhNIPx2e1jHkI206bFHhZzpm
7+zisHljxECbz96O8//aA+icAFRcPCIHrkNFKAxBUgcUF1tg7KChDU21mQ69
uk18TtkOKNizc8zphB0jX3XvtH02G/v5dCrkWvALBEKPNXAnHykvOcaVWk14
vXxcyXvZ3fAzMwJMLJ4qj1YofaTRQhCyiV1rAZL/ahrT3fg4Dt4zr/n83J2k
7177FIKeRBX0eO8X4O9eE0eOvX2zTsA56JWtQbLo782i8/d3+GaToqmAT0+2
N0yFmqio5Da/4vBLo8tu2ANvy453vbbPflHQo5s4RiU2nlEUoZvoINZtqLsB
RpeaQDdPiDJWpo+qSvzBCWQBUTUOoOJiNZmwGW5u6A1aYPybneVOujKbfvVH
Bm5Jnh6YR+Fci8ul0yeCJKJ68B+aLhuvV/5DAU0zTitdxB6kUuEWBJdUj3eI
P8ZXq43fimJDOwY1qE5NKppYie7nocNTyGfxiB8w/DwBEO+wfIA3wmTTmM/v
fjvYYMVlldoUPzjcWJojfabGRzXBEftCxMscTXXYX5ShMzs3g0CCggH8OQfj
BDLAiSLI1LqbU3j840DK3JNpKpKBr7/hu6JjP0L59q+cSuBYot8IqMrqzLk6
iM/rAZvDxbOkm/zpfn0Y+NyIxCjh0ddZHSPRMnCPcUpmccE65iCJ0Los2Uiz
KAa17AsIUH3VzhwFKZy1RzLIjwY9yZbCwrnL9tZiqV/IRkg98HA7FDHprqRk
bInzGwSOdUUu8nU8+0Ol1ernPzE64xvG+DCU7gfoxFOMnn1z90qZWLoVqy0G
HDU5JNdJzndEbkkUtjrlGL7rbGcWiJ1gKghjt/IzgLJ+1ZJgoO3h6TRqasqw
xA07e8tJDCV6bE2Eh+4IWKLcp41XLPLSIGm41Kh88du8kXIHJe+i1+yaSpQ3
e7wq8z5TaSHIK1UV756jWfbkuBOlNHO5AESITe+XMZVJSKMjfd651upiSeMR
LGGSfFcnrvJMU9I9bxSStayn3m5GwBh16U76yvg3bwkwXV0XbDJeuWD+S9kf
NBlrlPiwzeR9xKqmJcvuQ6g0ZmSwvD/52DJ2KqSP8B0yy812pTW30r9HQnQd
bhvzT3KXLxMDbclhQRthknuM1DtJB2z3MqDBLV1tJ3ozkEIqNEO2+Xj+Zt8b
82tQC+pzT+ucj8TR5O/zCKfCwD3fXVRo9hDW5AChrsWMhHMZm/d1yN6KsWHU
TRA0DJUgKF9cv9U84byC1WcEvZWMoJgBlKlgtTnRs/RzB+cKj44aj8DO2uKX
YhxDO3hde9HuE3wlUase+uJf5I5iVDEWJP20ksMz600r5UW+Asr3JS19EXGv
PokOMurJX8kdprWK+9h4mAOeB1C8vHvZdxbdU963qHTT+n6+E4/QAUdy6Max
hNVLdV+IgT2d5KCsZE5yxRQbBsqtzf4nEXzvXH2hIkh8o7E9no7YLqp2pSVl
wlvfoyvC6yUnRsydBqcsjmzZrcLWVkBIOo4eY7Jp0gYq6rNXUHF21RRDUDTe
H+koeCEzNKH4qTjTzfmyYw/Mk6GXCxwb3j1sb/EkBmIZdxEFcjf0TRmDiwdU
L4P3ZkCokb28nDeMTPA8Ulr6Rv4TwEg/ABagF9PjlA3Ks45o/KfZuytLsWoi
4GoIxDAiiG8Gm/aSC0x5SFgy3zgo6vfdfij96jHHVPwviOEgVuv6TlYdFepl
sLyyANWhB3A16fW6aLsQrSipUZD01p5Wfw99o86Ltd/kpStvowGfAuJBB1l/
nsc/7/B5FxcOUsrQAXI3R9E9l4MdO35Uqde0mspa88Ndf/u3zZJ0wGIHkDdb
AysAUqX9sksoDKTS+74NnJP09iC6xHkSq9+1BnOX/bQed9S06sH1ojFZVoJ6
jMew34MfcgEY8sfKE389rKqSHYWLYAvvLSqUrloyDp6z68iXnzOtxVFcxdND
5QFfVvFI/BRebBnKe+bj7siHZMBK7ESaxJlyfmPNf/9GoLoHwaOoLaXPfTF7
QDTnfewRU39kU5NciKTk1MtIWRmvTiN9+YnsY80RBXbbBYE4fDmABqOqwSL2
XGGL2De7CjHTqJdjoTjhU7ORb+ZYC0KH7v6FFQKRJI6HjdKgJXkI+k4HH+dg
ixSKVAR8Xf8vRb7ksnszmZb7zuv3KCaV2B+fyaHhprvznyg6/id0S6rwjo/j
QHFz2dS/v+/d8glEbByoI3OLr4x+eLbxIUYCOVmdG0nIOGgNjBwANy3z9iTG
Phq+DHVw0Ok+f+WF+/Ac6CPt9SwOfvAEg+uNSD3YosgiqZEaX/1z+jiajuL6
W/17YWOlkMbrCPihcq6FBQs3/ZmzTp6yY2WzbKP2KbuaGlQEmRFqrrXowgMw
z7m9odrICUNupdiEsrgoPpPMc9BkLjpNqoMDPIlR3T9GqEbwEWbwDUi4we4V
0iDvSirHCf3EqpyNP7wDHLsJJUPZHxy6QCscnq4WUyUveLNbPz4Aof5rUr56
XN1NtWcy/0fM6+CXZCruPN6v29yjL1PmFEse+/VZW3klpz3XsY7I8hXetwgv
PoR9BeLq0/tdcQJhIhudxfK/H+MW0LzsxOw6SpySxlpMG8PT1D6e8G88Q9s6
JmcRFtd3w7GcrDzAMXZQV5mcltP+L4fEQIc1HQ6c3eDGpIUEhlDF4cUBuf5T
o/1IgGZ0HE2JFPn/E/yHTeE1xwOwIXuXye5+0b2I3nX3ag1mZ2PiuvZjiWUB
H46oyB0i3ktbsyaq6ImgqkPZb5iyhslXkzaRpTNcS6y8d5//ZBDgS8ZVNYeo
A/jXzL6+uJeesWq+4DE7lg/wC+CFPB9I1i9IoUtX0pYc71nYnnrdCH2uaVM8
3o3JZGLZsLscdIC5l84US0AGSYqygoqzoDtvMyy2+E2DrnZKNqv2NDV09lbA
3X6wNYUXYIG8r2hXGZLpVWpwcKjGDb7VTaL1DGuw5wtrRIw0IS++2qaBvXIf
WU3Yu1ZNDfdQcDC1nmhvPakAGFU0mOKB1W9WSPDdzBxlO6ZdvuS0rd1d3lhW
TF+1iWUn50TxjptjjUbPBHzBxPDlc8bEY2MUrZJfeA5zZE5pQT/HHEMDc8/a
6/ZGYG6p2iZ9HLCtUMjJebvCgqH2oNWorC3bUL8icgZ6gyMOhOaxqCqNeJ3S
qDGQ2sDvRYF5pOGqX5gRHExoQohnIf06z7/TmYaF3zLFHtEJlFwUQNlKX63k
Xp7p2S+x5YQOwxPd67VicH3C7gfgBiXt1mFbOaUan3FVXisWpEVc/x7KEgtJ
xma2xFlZ3m/tZOIQX6lh6O9CuKA+qKF6Y92rkbzTJ6PkkS4DsirX85fENBoc
PlABx9x50gKoX+Txhm+PkFobiPR96X31tx9+EszYA9r5+d+JYuyfpQP47XXo
ALqr19Ehg1bPgOg97oA+MoBf+G7nyIZD4xJkZT6crF09B6Z+BSsd6HsOWern
EpzBc/tJkkW4pCbTXyPZJkDIAn5F0MVidH4hUd6x4EqFeXqcJmAl7/jbKibz
TWxBXokWZpXqaFVu2y0QIsgH6a/z1/a3QSoFlMn/wdJ77UPCyyE1bhviH6nP
mqrvQD8NNN0bho30fgM2atrH/HRpzKmW42/lEx9BkQy61mueGrILabw1/Vwm
UHlF0m7MJbzhMz0dpQq/hpwwhWkr6TZuIs1PS9bkyk+TQclw/1H93QAmKRQ9
A89psLfQiJ+ulN7SOhoOVKsjoX9sm6vVa5kJLBRFwnRuDxp5LhGxUvcaGagV
Klpo1ZSYoPzJ1iRKkbA3clB2y2FPeBumcUOM+mE85vA8sHOPwxdNlpxa4fSi
X/Rj/M1YwYh7iXmAImGFMIlf5tQvg7YEY4emodSc0F3R98sX77pKs+DQWzQ0
DOnmXGhTGpl9PEhevycA0GD2Z9lu6pH8AxlIZTwBasH3wQFQVjFysO56ne+a
sb8NyvxKqq/Q7OWveRCvRykLpClMseMzDNHVtJIG5UE//DOQl9R9AVWxeVM4
TXbyo24CH6AuSPkSaE8cfFzBwiT7XzkKhjwmuDiN/SOgvLl+Mzco+8ABSf2Y
aPGHjkLnzR9L3ukh1uxvp+OywPMQmWZJMtL58qhe4xNWPBemXV2qYlG/tPgU
7AR3UO3JJB/9UA+SdVA7/u2oZanFJUAOntkg4i9Y+6S8PpbqISvXRb0Xrl1R
sWFVZX1E3geaxoIMr7+lfhh0vb8xU4eySEGzYkK3zkHzz0W9bLQImeTheN9L
ElxhsYsLzue4jrq/r9gnQMj0h3NZG69iDHMvyaTo4UarsHb8PGE7BUingGCh
r5aysn5GxD+DBLuzCg+hWj8Tfyy5HLmQRQDRpuiFVuMZAjzma0xM9qvq/QqE
Z0HDD7hcbIAeIOCRfqalZJ53iyXqtu8WfPntxox9gq/u/KEoq1Qh7ux09lPQ
dCMf16pt9HF6vrwx6iXe3pPXCDB3v/0V2I90vXTzyHlsnG6vrQ8ICXssvasn
YrxfO5jjS8Zi5OtqAoKQ+n8LWJPCVs9Njc3+pAy+58Rn6hv9DzK/E8aB18rt
d7SwKvpfIR56tai1AWOkt020yuENvtJZ2f0BevF8ya3x5zzgdZVW+ZBL6JU/
qt6Kf6uJ0NdzB5+XLmaPVd/WVaIX5axajyzxwnm0ogHC8kLPBGvsdy3uFBJV
t5qeqnidOT2Et/rvI6ZBufyWRA+RXduMezra0ucxZg4STlTR13lXNDYw4hin
ijwFjTQUVasTRg1lsfykWSP9cHd6D0IkH5IjyXRL38SyiPfq77nZ1MqTbN9b
ELOfL/M9DGXgyos4OisRpiUn3La7vD8DytyA+1q47g+tvo2kWgYonYjJ3BD6
ftqtGvYXScAGlDqTcw2lncuRFCfJ4Deeu4A+faCyV3/IcH3pL3NSbV5GWuby
9zWsRTB3BhFoOKIPUanbmS0QkGXlexP0GxVWSioi01XmfG0+KzFT3mSQgDUJ
hDeqkZhlpfYoD0wmxADzBLQmTf+HGq0uuR4u2miJzHb0XXwIehzn/ED+M9B1
xZUA96t+3UYOCWrXxX2VUz+qvTDwXaUHQCDc/ffdtvFW2UI9FF5OWfHDkEY0
MwQTNcNnoZpyiFF9lwrqqyMXT76zUWVQdoDJIcwcql/vmvfNcvrkcTF25JAr
A/e2RJN4MO5KhEMhOK5Y7skRR76wT+G0gggBVcRM7d4OG6pJ7MLAL8te2oa7
q1ftH8RRe26Rodl09i694P+YeVPWE1v4IinWm2HKTQ2M7y3f5UsPRu9n1u3k
9g+CNF5mFd91NGt8JSsz+1lunfY7IixdvUm5vXLBNBO7gKlhzvuVNJkyeQNS
2E7n9e5HfRYUTXPSN9ZOimvfMMppB31KbLIEAenpYrWsYiW1VEOdBxkdNjjr
fWo5vYvo+f5F0K+Qc2Kx3rAyhuSBlAc8AGqeN6stoNjwZuN5TFc0Ak5+LqRV
QGYrDSottEj9rjfusQdIE6Gb4fG0FxE1LtI+CkNQ0hrGaLA0Tosx6QOcjzZa
ulbZeyMcEz9Mr+1ZGRJihH+uhFIDQgLvCmXmJX9MFtJAfB1uvZYEPPwfEiKb
YortO/glgrPcnAXg5UCSKaH5iL9yjTpAQTKeNqcIsn6dIRDybzVwFlIGkIeG
pxIh8Pw8UtAwHsrLoXkoxK2Zw+ZbNkZPe6gcFXcn7R+jEM96uU3zejtJtMOs
22G8FVSqFH1AkNOHv/T9IB01P5eymJu/vMSfMei+Ae8dMjDN5MriUnxHi3WA
Bje731C/bELamwWoRmhOVBs9qZXxhTzDM+nkKgVjImRmqdX7S4qJBdUQn5Oo
VlQMCqQDKM0H1qnuYHdHC4I2PcjN3m4g6oGBKRV7vCMcKB9U/Lwn5TrDHs+J
x/5NnKhzWh3DF+70tI0RYyQvApvcNdwMv1mdqSOBpqNFDCY8z38EOnWF/bMu
swEuTm3jqCWwe2g75r+tmTLmOsANr3NPxRNAkv82dCKTs1X/1GbpYnB1WcTo
wvXP3zOjVz4S05wpbHl49xL4kTKZ3zil4qSt8r8pCyIBfpekOrmzblwN7nJi
Kk5juV1ltg21e9w3uT2d6YpiLvqU6Q6Fyby752Yb5gMrIqqaToI8U4xRiW0C
xzdTs0AlKlywZLtjqxKjB9pV/9YolGBP1d4Y/4w+qsOv89dk3dvvYH3ONSoR
oBa1iAMW6Wk6POxGFBZItz48/jQzrR869cJxRLATYkGqdh8Xy2rzxZQ38MI1
80tGPnU5jTUTm2Jf4pZMkvVKZU2MGx8eBN58qxtcKG8hjRp8rEbRzVW5YL3r
SSUmOJ524gs4LRp8a51wEyCt0FsHJfCALIfMX6siY04m893pC9mh7Vnddk46
PlGUzy0DXyuLsWzJETq/5Tkr6xyEMoH6M4CSG5B7Nceq/ZjX9QIkzTP5zVJx
ZEfVuh1SLtQ/l+lUlFRnt67xQ2IQtLRUuDh2tTYB+lJF4qWqxtaPaXW1kgT2
TKVgv2X7xsUOv1lDRQGu9qvNqnTt27vGPvYf2AoH2C+1WTjH45DtS4YSL7xk
lVlxLbCEVhXR/FaL/6FnPPIOGhO1oslFxzEJdsbuqopx0TxOB3kYnKJA58+V
cR3bkkzNTrFo1Nq7O2OO1avfTVa8eiYfUKadRmRMu4v5bMHY3osnsdUtUF+l
TKdxbhtErKubkFqXtHNmIvobZ8OZUc6pokuVMp2P87dKKZ/JO2WUg7XGCMZH
2SqWcq8814onWqlU1Ks7NqdW/SNy726eGsBEfUYpV8X4PoUNlK51nWHehQOX
78oAJ/YP2KxTCcLBLPmMhDjTUnC8ME6EnLbEKySlwla3Ccmfj/rtkGNQLHrT
OGggNZ3Chz7CiD3o5rfQ+dBYDjJ3uSM/Y46XFGONMWn6tEWMIAdWY0K3KqX0
lpOqfE8aGvR5+SwgjkyjOzIWaoZRinewneo2wG/0/PKatMlzlxvPONtA0vF6
xizti6KS65IvDZbpD+zEzVLgiHrGLNBnpPKEjiI2ZQyFzoy2HXwGq43qLl1E
YuBw1zWW+kLeqPHCNKP9J8u5R/7YKGDBD4670u4St4mm5oUikhoZ173aJygt
cyVQ2tvnG8AaggOFqG9o3CsGW/GNlmynRRW07wpF79vE1SV92uM2xTpdhY7D
KnVRoOPwP38d+9LRLSPXkRRP0rfnfADwoxAlx/9X6BqHnMVixbOjfz6xlwC5
ifZCO63llykjtuiiV7BHXVpBJh5zxwrK3/sinaz0tltB49IXbqR2AWeBHM9H
Yx8sc86VBEa8TQP76Cd5kFZbAj2odnmUQCwZ7DkU7cb1WzMjug0YpwPIuWNV
t8x1/reek2sTJTx0Akec+HD80hENNTFKM8pBLimpgjXxrEal4Q7sQv8I3zbi
LifuTasunOu8sikC1qRAmDDqCCriN7nsy3YrVsLs4hlPGC0WhgHB/8wuqEjL
2M0j4X2ET5CiO348OXGy0NJK083k44wdGznLCgd99PJ+gtKysZ8WpG5D+A+P
4xjGuMfiVA00vd8c6Itm+TpcwCbU2G0Ag7Y4rEyFZ4Dm8TbV6iNzllv+Vsqm
65CMk5nGTT1yfY/YZSSlATevZSbzuoZX8c8lyN8XjmlAFZXuPa5lzUpmJ0oJ
DShq9gtEjalsgJt1J7N2JooUZwqdJmmLIhd8CimT1GtUvTYusbzuIuGtYgda
lCc8Z+mOzFjAAPmrhVC0TfZnDMnsbPfWUxskOE5MnnxzepYt0uUh3cx6cdrV
yYTKbNVBMVijsUVA63md6tIxv2YmPAgfBqYQrUAldNLF74r/cc9oT0Smw/BB
IUb0yK6C+/u75+7WHod7O9HbaYCCaecDsagihOeDbEnIP5zgVLnvkTWyvWfP
lwprEEqOE6FGxms80H+1ejs+Bwm2NpW0n2o3CBzECz0ibca6sNAgDf86+w67
EZUkJEK0WBNA7r7JdyVzAaVhHnDj1nYv0UnR6hXr7jp3RS/zPuS6L+z4qfZB
mxTRWtPdjHkEzwKaru2qaloubrp9j8SNxhfj8WWpq2LpdbS3e2rJkxzavg4Z
ZS5XQlgmt3t63b5TVHc+/5Y1Khqz320u6bv0pdiWcggPeVplc5lZIZrLe2bZ
x39d7AiyKGunPItxK15IIrOnmq9DMlX81TKFjVX4KEy++cONKliFAo/JhSMj
/VcLr13w9puaHwYpWn6Hgia49wq7YXknDYLpABKpnbhWSHvhubgFV0BJKYMd
OlkLPO/WW3e86A7OsTSuzanILnjj8mgM+wfzJiFU6GUu2+dPNx0RYHGzFTdw
MJKjKE0BilzC0Cz+vra+aDvKtMVFmqEk9zlgMLCc4Y8SbJMilNzDYId4rgxr
Be5UbSinV8ryaXWWPjbAcmJzluWOgbzATxiv4xtBMFeKCO/TDschSRgKlV9U
DFSp5K/h+aCDzP+rw26RP61auLivCVHZXt68kE/D/EeZ9kGiwvFY/E7NmRnV
sisBvRdMCG1zb47CUHNAFrFOnw4Vp+ol8BdQD7ixZoTAP0lK3/S5yxMie7og
aW+gYe7To8oTZsH9s8s7wd70Fv9K3kJuf0yR4YLiMGYTiW+gFPhUryvaDRQW
Se2AGKbOxVWkF3JEilawucTJguZNPk9rcLpA6XCEzl03Zxym/j8fh1FfOHuO
MRpgBmdJ7SnKFYryPqLps48FCARGMM9gRTypihgFaBQUia+U3imYvZHD8ubL
ZajsYpZdVBuGp4aeDbN0Jm0Sxb8fpmoBqgWwCtZtF36CHxa8+TOxoCATzAgy
rYIiENk8JYYAWPMy4kiVzJ1ITTaxRvl1M07EAb9NMLP52nQ4t6mjIg/a0OdY
ub8WBlknY54hyvLhhwnbRH40+ImgVcIZbMrjbrOytmXSSn49VRgLI03pIOh/
MOdHhm+CZP1unwsWCPcr4wGKzN3vwup15m5NZDZuKU1TR8ng5ETxqWWTY6Rm
m3gwco0etDbL14IM2xr7C352YTCLUCgVJUW1DPq1/EKaIMTkG4KiYv0vfN8B
29+QFl69tqKKZ7VSlmDoP2TzcQ1mpDu3/f9BAVN/ZAlS8im9fk/ODG/43Iqk
NbdEZMcprtLMfsAxf7glteZohV10WIMxR7CLNpraBpb1PDgJMlqYigSd6HvX
IIl0FNEVV9lSAgYzCsUD6iD0E0T6SH4NAmhT3+GDRkHLvFEDBvcy+6UJXkIk
ogn95T98FMducw/kQcuoJVv8k+jRSZnEdiFFCLzwYzbcnhwDrs2GYx0+5/Iv
wLuOtOsS9rRHZQFMJh9cT01EsIMcAXOD0qXMrU2h4RmR8p0lzFHiicTckA+N
Giktqe0ZihfitUq0UIYGr9k+dKXk0NpbAcu82VDUx245iBI/dfc/M3DRpax6
r8VGw+5aFWaITQ7NokHaNimhJXizDe/vbRROrUA4gQcXPERU/5ybvxQdBRwb
O5dhghsrsImRk/pFwbu7oz9Xn997qslvcLqDGDO6YZeqafTeg35qyyESBIqh
1qmebwNRW7AtG9DL30w76GjxtcpXGCLU1RyqP/cl/T4UU/IRaZYskodetE+9
DA4oNC6/fg7QXVv5MptWNFZpquGxTYfwkiy0WoF6Bht7oH3vp/vzdU5JTqCr
9uDwZtSnXbxiTTewQuVfRoqNqgJeGDjG9Zpv/2mU4rvIgGU8dZBB8IK6t7rx
QBXuUqP2pEaXVZ8SgV5E4sAP+Ta43xvF2Co6/ea2C15QYjagOo0aafxhwaxq
7qFsfpu2daaRQm/loSpFNSWKAOO4ab6+xHp5WONxQFfJvlFYSiByUCzVZ+qc
OjUzzRPO5TehNNKt8N4eSW+FvgeMmX8BFPBzEteXac4dtDNoX5Zu0YABJtFa
ebMl8UX9pUa/FnijqtlZRH6r25IW4j9aEuG3AWUNo8k+o2MuZCXHI45klBqS
p55mCZRyR+vgTCjAh8EYdBVrSUe9ChnTmeH3Ptn0Ij5oGzT/peZc3L50NEIK
2R5bJGtRxp33fSdof54+h7ecLHs8JK7JopbPDZO/4nVcOw9EAXLIW5qI0xIn
NEGR9l2IaK5hVRX4U1NiethBCprwNq80DOSHwGD61FC7gPCtf2M4FLE7VWcE
EOvnbp5YkLrFPn83kORkQ4VWh5mQYHQztqQzWhSnaiXi56QYSWafw1AKGcy+
84WBBM5zydY0Zs3siXUWeKoifGpRhJJDNmm+ow+BPnI5H64cB2uW2o41idau
1lcVxUM749qsDGo+1wsvEx8wYF/bAIQjRO0tdrh31m/0hNdNZc34IZWpwazH
VzSudlG1rC/Jp2Hk7RgQoh/BORw6A71GxIGbmE55BQCFKiIcxF95yvAl6085
B78nE9rbo3nVy7qzzm8SeYTaaPDGbsRy22Xn1Gc9eFvx/IlymySWDfZA7hOq
DnIwX3Y1RFr9wdp8olw7cv/bCy/6TC/0V7ZkUluubCeAwZW3Ayyp/2wUBKIm
8wthyurJLvuy+Xe5JBj+1FQcIJggSyxUYn8Wn4F9W+w4iqVqvJ3vkIyEwqXy
F3lY1wH7dwdOZQbDEBbACsOaENrct7kZPWIRKQ8/DZ7y4IiP4oM5GrbT4CM7
t7xqSNRzP8fittFSZAcECD1Y4oRmBI5G2zNzM57HR3zoyqVgqnig3FU0JOT3
JkwXC8ZG2MZe/M9A+M4IGYfsQpYLIvCVn2U5BmD8nyElmvCgJcME/QSf0tnV
UAchfFN7hXi9IeEtKn7J6YFNxvjA0wg+3jKm21mEPQE4A3aUSfx6XxWc6/jf
w8GrZEpVOOehePjfTX0scZ3g071WWEZBYsDgbe5LWSZ1gRUEMDaNMbtVxkJv
yPKOrhw2aXkfS14G54c1qetv+ctlf8Ah0gq0PnytPL42lCjum/58Z2SYokGI
iceH+UkvGYGplMf/t6Dh1vZJpz+1rjwMB/4wxzo/nUI7LolkmN94C2+yA6HW
OaRVSv29E6wfZjbdO3bIym8iWHy2wLgYuBiEwC+wSjagJY6FHYUuF/PNQMBg
fGsdvIsN3bgj2Q/C4p0b7mSTZQ5oxux8xnmhT3xONqVzNLvfMb7JX9X+tR6h
/dyQMypPYSOvX2eG8EBX+mMupAA+OyK5D8QLqqpbZ+xNqWnFR+m0O2th12ED
MrhvW/RNcVBFR2p2blwiFxK44LHeYtuuKikJS1Vts8kBE/BdtvGDJW9UaLg3
jwgGfvxfQa4dN7ge0908sOrNgS2cn4FR+iWQFu5v3Lxn6rNmim9oTiBCWafY
fs7tCePuYzkpfKi0cer62DlGBL+WLcqdMf31/IfmuwAuqajRfTjI485UhiQ3
03X4KXrP5FCq5l6/u0OLewcCH6RQLZ9wLsash1GJKAbzRsk2SFMneU28xTJk
3ev16itX0JoXsXshvFV0EzjlHavOMqToEj4/tHY9lPjLPxol500Jmok69Drf
FLwJXjFcMUmI2fBQ0ZZFS0CXyawjEG9WnwhG0/XJGgVzNxvuFkNWmpRQ+OtP
1/Xlfge0mja5/GMIlErCP6fN2E/2lpApdwBf4U6uEIJz3OBSyPePVjCmunKk
9y+Sn7RDt7nMVDUWTYahvaAy2I5g3sAesQ+RBSncMwptwKKGM+CEbwuCyb2g
wWrAuNxSo2ZE2XZ6mX99OZM/Z6DwmmTL1xWeLBRJ6JDpS5863pVaLayggm48
EaJWglVa28vkgdKYQ/QLLM6xfHX7JGf3A3eGVlPn2RbNNX+Wp/tCAUCMbywk
nKqolD8bYqarUUEwcsV1s9BRvmDdJ9BBfd1ygTfrefoMIq8Guj0iLIZkRlNG
X8+S1uwsFfknwwIG2OoDgdjTJwVr+Onk2vM/57sY1pDT8reir7mmguH6YSwZ
XhGNvYd7CRP6ScSGeBedkMAp1HK26TfqRUYMLxFMulXqpfiQiq5Eyhkk30xG
hr5yQuUQnJxQ9hoOGlF0ei7VJgRRdXex1kF3/wcKCXM/GHh1we89GbjeymXq
aygPpbEwbj2IUu6Xd9Peh9Ihj9TbdT0y5VOdHVnpyynWwUXOXY1gbhWTPKU0
Bd6zH9O1eOdYCB7vQhXkhmVV3+SWlkLjVzGdpCEK1yWOWdAu5hHCLAf7Zi/3
lKDsCbWrJ2rtJad/O+zQggg50HTVwW5uVCzecw2Im3UJNlQdtRwxu9U9delU
P7IoV54/ekiFf049aSe/zDXPqj6EfKmplQAFeiEBeiAKCdwaSnooFlRFcZpj
TD1uUTbtG3dxxG2GFW2K/i299MfF0rRhTx4iFN9YWfQCZ04+TjcgzOyFvjeC
mPg8YpEEDtjKC5CFJWj9AgDN3bD/8l7+fk1GX/91KfD7K27ObvAwRGLfTzX1
uLCS7KhFL0Jwq+FgwxIakjkN7YavwTwx8sikSdXPdljMOLuqBw/kawrR1ogE
gfMYV4lU18UuFMT3ANURcXtHNYcPFCMiyCEz6d6/PCho79cWcCfNizRM7DuD
Kcts8nod4keNEMVWY33Q0HU/pm2LYMUr3wBV3RP/I7zlGLUgb0bEojOIGEN4
rpZOV/Zet+YTdiTrbx0UxDAbNO8rCYeUWURGHEHCVqqQKDkEsTcr6KtbfxHS
e34Nv+Bd4TI0GEmSUwgrKGMforeQAPZ/3Pdj+vJcTPfEMaIeIqDd8I4dzfpo
WWta0TkdZZuZh+oxlstysd8fuZRniVunwMvJInEW3dfcF2J8vpW/r8hMv8hn
p4Zs6NmHUDh7sMvsQcKrSjCv/9X6AxehkrxH3IELjZPd6+V3liW+XYdI3sK3
Gb7ZXYBJpuIEfmdPFrmjjsRP+poT4VPPs+L68t7AI/inqhYcnFu3plzhri9x
8Qi9AWTpUiSr2eD9yzRdbPXKKvhetCWyT9zHvVMTZD0I12H5vZ8NSO3ppoeb
a1JyXbSZIyNrMQRyeMPVGwfwSOhpDMjgnHsZotERgU6b3qex3V8sd/Gm7/9M
FEHQPaHvzL4c0EeKeUp11Cvn7yID2MaQVO7eCXYYk0jHGxBiLSq0svYBPDG9
OIX+4MvzqmocfgTCeK+NVXVbO+BGPT7dGkC7XIJvQf9kJAt+UuH2jpLgaYjC
7DngdqZn7eLRGNFLEsEC8tNkuUebR7imJvDEkpYq9FNDLn6tBhmVgFcrY0Oj
qSA/lEnG1aQTUDKBemqpj0Oq6gE4ouXMP35e4V7YCAqwsgCebCVAY4fdJEAR
L7ZWO1TBJ9bx/7XHzrc7/eCTJgAovqw0k1r2oCt9VTWSQkSMb7ZXePvHhM9E
hA2YmRS0FWpJn48F0/yM8Ff4xafsrmjV+NTDBfLkDpdlhvpI7SaLXYvBMiMX
WcQyF9qzBPJSUsWb3UiClio8Ey9XaCYWPivsLSnYwnatcsYh4LaKEObhGopS
IH9vtu+Jg/Meu2fOCkmDrCzqXP0kTOgrE9BRozhNkYI8qDdKCqKaGWSRg51d
7IZ2bVkVpffoVfgcs+EYuZL1e2WfjYCZ15UaZAd4aG/aPakLT5z8vzCXUWRh
VMDZ3qiDSiXSwg5616yE+wcsK/1vaSRSlj4dUZzRUMTSzJZQQ5kS81fwiGYN
L1MoVl5eTaw0PSvin+YaLzkIu3jrL5w/txXeRI79Jw8Veq2igyuOjjAWPKwo
ytxO7eBOJnBxMbBTZBvNm7dwy+AheQfVIkNNcOfZjcYwHMD8dgpj4uGcnEJz
WYxErGwc9qIz+tO+uQsxkYHZlI29cAYZXS7tr1jGdyqKz55xatkfQgYQzDlX
xIPheYoGnZKLDWzL20X+09CoIFftDovgHZwLGOjUxL/eB0SYTn+779kcqI6j
dPtbvNXMCFfPItNujHUDy0twAEbe1XtYJf4XMgVU7L8jfJqoFwJ9ASKIynkx
y2gvWIF2m3VNRF6RVjKXvJQHd5cPuBMfUqjzvi31QJ4FmUAiSeg02GfxzP/M
Ia3vEz3VUmhWqNGzCuZ2TbbBAaoHhYHoFJKf+oU+7Aos/KS+EnfW5zaQyn7e
LbLGJlc/PXItGJkKRGjEyAF9US+dWRQhVanJs9TlTa2J+FKSTZmrfnglbXfQ
dDbkdazEH62kYwcjn6Fl8qeCKbgQzcA4Hk3OadRGxSmL8QzqZJwycCeW0BcL
W6RMPj2xx9tufFtipIjD3g1LFrAZl8aMqtAToCZlRNU8cOzx7N3B3HB41wb4
ING+CI4gjIaowY8zSTNmU+7rFE6kukKwtu9NufwpvpMf6kxP8A9uu1dWhtQ2
r0un7HN3IX2qyR8TuV36ydWZw1E/bLnSonuFKQBr5t5EHh7443V7mPkp5N9Y
7F44AO+2jel+eb3ojef7y/LGALzABzw4xU02nOn8nlnBgJMO+dNDKRxAGzpm
DKX+V8dpPDtxnXb0pp0lazlsARsgmRO597w2NOgbdx0N24Uzt7q261qDrkXu
1FzzIa3OrzmRdbG4/4xntWJGWCDMkBRj6GLTs00qXuvtkxIQz408roJ+rbQL
hDsQ17unczCpe0lfzF3KxTRQu8F7clycjILrvI0oqbo2pWB+T2h4lsxOJgR+
jhm0spr/g0BQsTJUP25l/DCmr7VQi5lBx7xfFDilIU/YmUDCwrKREFHPNarX
yJf+Qx23qB+zu91j3PCkw8yNb7Izp/z25IUum4ObF3YuYCSlLXmPcKwNSRxF
O4ozPkExHRyD6c/+jrjb3lF6ZETMhLJpupKQRM+BvGE964mDaF58npeMQrvC
9gfED6cTmJozvgaEZ2DFTiInx1L3mlpqmvtG0BTk9Ai4lqE5vEs7hq4RA78R
oaVmP9WjKzUOC0e1PVTnZWZVmwFhHmvtML+PCriOjYAW5/jRLqzDFKHxyu56
vb3X3ao1bWNvilDlsq+oqSjIjMxFCUf9h0e2ZpdiybvYCqe83gD00c47ZQ9i
8Qi8rlQx1eGlf/xU6jySvQk6Iof+SsOjZwX0nRP2rXSKI8fJN+CH1WAHqwHe
NzSW2u4b1Z8BY9QxaKrxgFNFyg+FF3O8KJzt9Ok5lgSUtqqLwJDDXJLSGUyE
EpT+Gf91DG4R4Pc5n3NQ8PN7fJI37uBN7uSWlMqieEqV9VxSy67uYsGn2Ml1
kaFQZ/UUlLXGZ3k4NJpL95ycECrkkgn2Io/TlCCvyw2ga3SOnQsHUABhopNo
n1z2eiOyXTxdUhLbmZQxwGi6QLfzJucM1Bkki+W7ZKWJ+C0fC/uGtmskzwav
QUYqBDC7+/Wb5W2IZLKQ5PSlLx2yfiIMRaWBthz3ufL9mfe+yyTpGK9T7OGz
CorHtRF59cV+vaUSemIBtLrvlxAZUa2y4qBq90Ym+VMzOYtA3svPhd8pcYXk
YyBMr1u1VWp5c1GguCvG5k00P4urqxfLb80F04mWTLeXk6HZuff+IZhSFPhi
12XRXGLJo2vFtUPOcIC7VqUN0z61G/dMDS1h14RoHnDIOdBjG1v7MVTFR1fS
NhSL8FINPc1p3ebarRsEA585MHxxVfgT6w+SzNHcxUUzYhds7WtpPMYenB5C
sbkLP0KHOHOsmr8EbJtTg39QGfshNr5noRP0kiTtC5nKN4ZOYlI5GexnVC2y
tZXIcau3W/2TmGxPaCEyADoNsV9JHtC1vYDvEWMlM2HT9CfHL9QLY2oe4cj9
IhbTAoI9aGCLEY9L4ZJbQq1a4jem59uQu5gzMcmYzyAJrLauweN9Qzu5CQfm
x9S4mc0P1ZnpT0oSmGb+rhfbhLIPRM9kTx5NsZSPlX0Eybah+FLcxXu/xPmA
mLSXyUZUCgQwSg0bWjeldv9LoHri2NRnxzIfbaehdxpNlgw/uuxrdnwKNsX+
9WG1apbBNTERCuvej7oAAlnWcJDkEYT7v48Ym8xvBN6ZqfwhTtvdEHD2zjIA
FMqD7wzLXPiaOKqExR8dSnf89xrOJuTK6Dd9xDethOCA8MiufceHa6mNJfr5
zAvU37ckr+o4tqxmdGWCZEVQ7XAIWktmgZZGgzcxKLBooXEdlty+Gqb//dQZ
NCPKs54dZ/FyYwlACrP/KMsmF9x8dqbl4nmq5qzqlGvfk1c28BHWAomd0qNg
6daVirpUJmp5BP3fnJlgLesBIjjWmTwGRJeUZdEuqKHkSkxtL3pxWUgMCaj+
pHy2AHnxFQwq/vuVJd/s6B3dUogbLfiEYjxayAQvhrW1fn+Sw96NC1sZcfYH
SKMBblHuWRX2HPGMcufzzqbqRBzA50BTcb/1jRDolyjiHkIaHxWK77TvPB3V
a9XE5XOyWOdCqiclV4nzIUdfoISb0WLW86ezawuvJ+mX4i3YxZYdLnjfqHkT
UWhMJGTxPnGyqOP6Ubydtkhrd/8M/bLa6lPCjAC/vKEhebZl0nPli/OxkdSx
hLwJ29SQquk8XIEZ1hZG5m1lHhUJOmYX1zniU8AQ6qPmAuL58LQr35Jda04k
x+lVmH5cDrt0JSp6okPYmBCicYwzm5h+iwdqCokTwisEsJ7mq3omxwgTm8XD
S7MkwZhgN5Z2a+E6z6LhK8ifMZYaIOiaTgd59jfkd/hqZXbcUI6Fjyg0QQoz
YnMi/G5qM5FVFbR8UKc2PD2x7n0tedTxNzY5WV1vVvukQI5+TnWkRVnympr4
HZCpRlOODwPe01exKrAdiWQvyiySzDUtw0XtQ+7vOb61pLBdYion/8hbVWVv
JD4NdRPoyp0/5NI5sYC1LtNH2fPFsczLWEpJJg8UKQ9piYjpXHsQdTO0ySys
I32whcRLvabEn2RvRfp1ev23FChNn2Kh95xelm1N7EWwxqYbnvY8CBHY4+IV
U3ywZxvehebeU0QZcXjmNya68DO+z4XKUZZ/iMqOda4n0dycre6Pg8AAkE6O
f0M3h7WV++6XrquMoFlvFHH58tH5LbJXqgM9U1JdHymt4OcQ9oifCNWYhnda
pHbgLmXDBZfFVtQaD1yW+yZ9oeIl8HBF5gUWhXzHTWQvQwgVB5g6VZfPahXX
ClKozYiw6ow99v5E8pcB4oukFrO7OyDir6yUO4EmnXmxIkjH00XT0KeXQq5Q
V4wOSlLpW9dEtVnkU1eaLJnHFpkaTSYB3NWfcvFItTMYwt/nmXDk3ETIHT+f
NYbU0aEa4OF/lbwKWw/IwuyrloEluNUKmLtRoCrbq1f57TJdRc9kyWvHDwH5
OwImCVvK0cSBXrosU4WsgOp6sxZ233k6JM93xz0glHfd8PW9aLKF2rvN2L1a
JboQJ2s9DbotT9kuPdjzVRKONIXjNtUAmLXVdrLgwP/IPWWo+0+FIJ5dQ8qd
/Tn7CsFEahgk8MwjSglpS2K0pHSMhJiJXa8yVSxLyjaIkCCw38P+Ky9FrqQa
QTU7jrig7CZ2ci1ldX2+BZj4Pr0GWYl9qqsQz2SdUhCe7E/qt7CVh2sZZVmo
332mgNg5lcTq5IucOYiDB0+iHDd4wBVE5hHuPWoG1XOgucPnpNii4zPxlMuW
aSSDdp1oY6jzFdKNbUpJevRzmLYs+lnCGSeBVde/bFx+n6vfjfPC8IswQDYf
xtMCl4XQh4Jsp3M6CdKxMjpq/Wy4xl3hwSlliyiAY16mVelnJtGQvkiNa45e
4LkDw1roBKIOc8Z58MBCbfUw7LUtwUEtwXf/4X2eAtIEmen7Rdosprh1Qms4
wvxItiTuBY/XNR1uetmIMaZowCEE/GHL1jeozquFROGKpfZyAItOL5sChaut
mc1AvjTPmw/DTaYR/RKb+yP24RH+t4HDBRHRKzPvkINR+iwCJ0CqFXWwoB0z
Xb3NorwtYOx74Xy/s3zaNLR2tdRGKqE5cbVhpaRQ5sfmHu9jDjGcjk1rmght
jEAxQk0JBfIUWvjxy0sSdIr8JlXxGKzPM/+W+bBLVxHv6V+nRHrgzCWe3WPz
UckILKcSImEvhoumvDhH3UTlb36MTj21h2hC68fi6ov5hTba7ArEuCDEpkYT
iNw2WD5IBOfPZmBU1GVc4fPyknDafYIhc6jT+PoSOpsTwJJ0WTQEz+VobKeZ
S4jOaaT2DJb2ubgjIuxviXBElURUDGZ6NDDEtfoWaSmejhurTqA86hqC50QQ
RXZubKJTf5SDN+Tp5l262x+AWoLKnzSyP+1hV3AWQBnwOZcqOsaHMMI2eLYz
kZT/eKjIiC4GYiyqUYTE06BugU9RyKuuhBUgPqUuCBK0CU0foYnDtPi4QgnP
0R0ZwV5BfHWD6p8BofG1R3OqrDAHTaF30Vt+si0IslOR9sXWZsET11aWutuq
NzzP8+Acii7FSzW04NM7Ius1S0rBTpjxkMT6/m4zjAc1etRslP81IE/g+jGz
XswVA0Let6ZaS4UVsEZVQTF4WG6z/Oj3toLicZO8vaQ4+OUYECE0VKn7R544
XhqCgmpWi9Zwluw38xVhi2aSh35gRQPuSbDPC+PYeIXBdtgUkGxysVMdk6OD
fYRTQ0Yw6mtUFj/IiS58+Dgq6R27yZM5i0XEWIS0Wiu+sPKb9YgbJk0jST8f
GrQKN68o1/cPHDQhUWzA4IWzxsUW3bqdq80j6KSIIAJgTf+pFp9KbOBWLvpG
jVuR4KjKGPO+dFwPpAlLNNktMbMdecKej4qe7hGXMinMaDhlCVN6G9SLw50E
s1eH9GmsoOfw9O3Y/TcPgDqH/J3eJrMsW/qJVNEt5SO5JGzL2fq1okVSo69s
TZs89IDWgDNGAvkq8XlFiienG5+Nq7K4aMCH8C7/ZO60b3+AxgQb/QRcnSJw
FAdeX4SookPUU9wUimz6iqtLh3qcFLM9LIhAwA7TF+o6EvRqzrRkXSkx45tx
nsPzTV71KZj4BmUlm2QIwCu4GmThWegdpQVMa8U5mppDELDfLZ6KWCukTkW1
qFGbsHG/hBFzhpikbSeFk3KVuBC5grR+2Mkq4MPHypd4sRjh56DdwiNkKcwF
WBV3OQvgUglAGS2NsigS39PkiNzF8R+5Pzj5CEGIl/q+542f45iy2I/RNAUR
yv6yP/giQSfiBRBD9zIQKtp60XscI6bOjcxQu/o87nGtLw/e1QUI1JPOAkpK
prWqTOoqdRC4rvIrOqe9beemdXNwKNQtFT5PFRpnGb12FNMg8DOG87xe8DuN
scEnoa7tjr/KZoed2F6H+SQ6L6NK4WVOllgBe0iWiwMCXFsJSXrEdK9+n9gR
WRT0TcLyOrZY6oLcr0UIWKkgrr7QS/LEbc6VEkdvkp3io3T2HOYLkShkkv37
L15g/QxVI1WoUQSvFWwWJ55HWGx8n8X6Y02S+RXwN5pUQAqG5h7nXQymiua8
0I4vcPilBJJ3pYaXuQYKXw+nB2lMYvTmYjZClwP5VNkgZrDWsIO76Ihgp+PW
Fy+nempZHiuzvF6bQ1YBZQ1uMhExosLjL9bEf/LNOfQHLkI8vtoOUJbEvdM4
AjCfU5Y+JdITKE9/5e9504xtZvWIWA0OLtyIPlkkZ9LZFF6C0YnHpFN3BWXm
wvaIi1HmFmGkRWNTgFCeWERx6TnLML8V6F8Fmd/DKaGTlYaTz9op5ZgYfFFp
E+Bg1RuKnMRHWbqrQ6c3r5eL46Or4oB5YnDk8n4IbVwVABkQ2alwyT652WeG
9grFbw4XA1r1T7FXBwZRiFLf4kdVyKzF3EcMM9z4rCecI9NP4FQspHK7Gwxc
dEiqRyO4K0lFlXxf8pVg4LVRTKHAFczHKb+rljyV32p2vYIvch+NSUYWfP3q
StqOF0QLnOkORDKuICzJOu648WC5vKKQMzMIf0h8vBlZEp7rR1qO3vXiWqcG
hdyGZjps2p8OkQYWZogfepACtQ+tVx24SbxnF+/ZZBiTvMbnDUcKgKSwpfsw
rmXM/S6wLksJ33GN+fyJtWtASlQIaFwYkoPOfvdjJprTZbnGmLhP2xuF5Cjv
e7mxhUHTXht9sjW/EEDbmzNyuZq1Eeybl/7sOtJ7ek3fsJSC80/VCTOgeY0i
0lZTWFSIIFiVw6M/eP6zaVoxIewm69iiFqzlt1FXfLsbA0f2lvXfYqwIXslc
tUA25O4pcBq7KJsr7Ec+PSCP8/dOlrJm39+EM60oQr/v+2z8mmYwjWdJmUi/
QX4QcNp04FjE6KpWhQhuQUTXIbnmHNJ9ZOnd4s1yXsdnGVGDMgliQFJmrq6Y
iKngeoDKeeyk+cegsO/qk3+7OG5Ck5TBC5B0EZgMaR8R5tp2dy4m5rlmBbWc
ZoSgoqqZux+GYLhs5R6IACPQPfi36kV5bJ5e64gU2GR/11vON8MenlRebe+o
voc+rXEctuSj7gceKiujYb/vj8Fy263/HP+rbNw5eOQ7weAOd6dowR/WTtjP
+DEj/fr9wadN9razewP2xUwgLD8SKkA3hZsyatnnl+68wfy39AHLWa4en7VC
2YdMGTcXAicW0kmNtRe0hrsXcIa3q1fkR6Bg9UP4+ludfQHK7Ne0LLau9N/N
A86lbV3Utora/k0Nc//Fd/srj2GHNS8/2v6FicdMda9NELSw8Tlp9jVRf+Pw
aDiC/GjmuYSW/Z2sZiW6GXQDQxqD6dPik4n2kxPweD9m8i3n8lqM/DA1dDgH
+4uKI+PFTOhx12M8n0LUoWlUPOF6KEF88g646qPso3wOc3BtUAPrlJq1ZuAe
8V2cOlEe9jlYhveqqf6PfhHJNtyaVGFAnDS+BGoxhoA13q3qmiq3Zs1EcUq5
t4Hd/sGnNkJ27ExzLebJSRFKao4cpIKnS3IHBTC2fqtsubkDk6GkdmM+wcJi
A24AgJmF20fmsi1H2/FxKxrtJPrlfz7YZLmpYx0bsko0GQSyoxMXujmp47wk
PE5z89HvJ/JbHAVv+YGHLtIOcjTmRXUxHEARFEdrIOhsoYmn4Mio1eGb1S3d
RXck2q5/YbI257eJYhvBHUnnPrOCv2X3rWkrubnJZ11n2QoZ05H3XsgMPZFI
pE+aINuMFtrh40VasU8hlkqdQrnWVXhz7CLQcCZVfZHB/WWNDmSc2rRT1Fgh
hRIQ3wpJii2jPMZJ3AHezgKt9njV1efai0zXXLq3ds91QT92b1+ioQ5zziIV
1uVRJS70WALe6aEe0uvWnOfdjwQzv487St1Iyb2JRqXXhLsZmn4Iz/iKwntS
m3lc5Emogj7obJbg38GOpcdcfhXK1ygfc8A+p40WjrR/qQuIiRdf6NhEqPx3
GIis3r5K/LnLM2C54PvvgJhDMZkNMKPvPLFzOQALK3/yElrB2r9NXUQGi5JD
BWZMco7Z7pz1JfJwcwvSYfrIpocZ1O8+KLAY6CRnkWsPB9TZjc30Ye8m8dAb
4XCBlnXjHSwvnRzZaN67w2EkRbDhkpi6Js4GgEyxwU5RVMZT+BdspHH4KzZ7
gO7wLxRQyBSZpYjIvVJlFE1To8TTFBfhTloMcSB1ma4BjA65BfAhcey37zvH
ODN8+IPozgeQpZ0f9CFeuDVDfTIkI2F6kOvpFhHdxpSswf5TeMWjN1bybUkP
bcpIgzUTVAlgoTInNJLOJcKIbFJ0kF6WclrlEOVshcUy8rGe4+/5ip9bzPOe
oaOBcCM6PpvKTuRMVdKcRGpThCOpN1jl0EvXpavDzXEw05s5MFaVv7puefMl
wWYXXsRrP9TTlyXxNjpHfsUd78wrdOeVAMcaAMGiRwysmTj5jo6ywZZ4P6Yc
ct+fTfHBM4qG4lY6Q/W04Ic3mdms1Q+ctjd5Ke+FdouMAN8l6kAwRPbP0Prp
jsyQnbTQCvjV2fJb3nTEBW4g7qxyYWTz26NEXZDNuqY+y0Kijt6Q/wTIEb+V
Z/WgO7BxWiQGTOWIIBtM4LXtq12XoHPqZi5P79qDSMRxN5xkHcw+QrJlFaSB
VixoImLKtt6ivRpnTkOwYZPUWAxmrn2KoMTBpgHQ4NXnLdMg9yjG1U93hcte
f4hHEA3BnRZVmAqZcPnbWp/3z/y1sWqJVWFNX1ATKNwnfrqnY+Y6ZwVPZMNb
tIJ/5IWepaQvDcZXmgRP5KSKaQPGiF14nxh3FFLrwEj8OvdOrXHIQsmvtxO8
ii6t5zB8Al4mLjIBuTI7YkY2ykOfK1ScXl6B+87QR9IMgXslHaD5hQAGI2y8
Av+2jlFIjkcsuwf0gywifiEF03W46KB/LsY7SVfa2l46KLpR2IliR0qIDTqt
JFCRvOaN3kQ4i8RuBuyaHAknoJovIrDJpJ8hOjUnBJ3HVErJ3AJhzU1QQGH6
vnOsmaVKHOyQYeSx5HB3E7RIbjE7L8lc/6STqujmrPaE6Tg9iVZY0FBf9ap4
4OHc4JTT3oCvpXQNCC76oqxh6WCjavbpPFyzrdDhcU8wQRqsf2k8h8FMaPTl
qg1aL69cMZ7ypaMYZMg7EP+Rs8+wx41Wa5xOa4vehKivVa8lsIIAksL3HXk7
hmDcfUVtK6gzjYj/2m/BBFH8cKw4zucBpCvJqoKyjNE2dpkmw8Sle2t3QdRX
sfBbwtUFyRtUCr018JrR5yEBtMC9x3QEQmfhzlVRBRcCCsn8FviUMbAjrd0g
tj4k3RbtigSc87rOaIsoJZQ5cxPe7tE55Z0thz1SvHOld3flluOG0JCVPNRR
M3rNCsIqWqpanOZ4cfwdJpIPyO07ghjzIZbj3mLCd45cPDj7xiPC2Hnylfr3
gYV+CgJ4F4diiG4KXr5uyUwAMk03V9J1qrpb1fl1sFzmiEUb+uQlWacAOLAy
qxwOe0aKw1zIEFQBkFm83vCMwAz5omYkdxlbOmKeglZbBpU6nr0SLTMF5cAw
ATS+NC6mBHIz+PbmmLug5TYXei8Mxyhnj496rOoUSKPj4CcH9H8QttCYXqXB
s26Yz++MZbEU7+YIFUN0vYZCLxzBdKaChoJYXFrjMyqK8aPVa6ZWK7ubpi3+
mixgpcd+HNfihSwej27/rfdBgibj8EAIRMtH43Y13ajecUUc2BUPSmvlmGzq
ucCNPyI9qlTPz5T0O9LIYPld/ysnkMs0zMbfmCKZl2U+0aFH+JBCndGvxHwY
mwBZmGsG2jsk3p5vVRjKCFu6R9BOQsSIl8yubmMqs+9m4VZKxk5KqoquYlf3
bx70MI2Mrit4AvaRmischXL6B9PavIZgmObN0AKLjcJZzcNbwlhwiBJmwBVe
ak0ZdyI6JqvENNwNRXqe5YrmDOsnGnaj+l3NRr2sT+zuOyN9CJknrrCxZaaf
5z1jEUDr+VejvwHczllqlH5Lo1mNYqwxHQTk2h9z2R+fSts7ibkyMQgDGtTe
9gGAKjf1oV0zIOAcImg0MRUJfQi53sSD3hcZAhWs+wTshHNsVsvQb6JCczQl
qqFKf8jeOe2tuOKlWY10h4TFfU+p9xXUxpCTxa+dxhVscGiBz/wXmR6ecvoA
rMe3wbgj1ICZ+ViFvhpkqIEtfjakW8gHmIlNfjzMYG5fkFni/tB5pR0yG0ds
PfDA8cKRF9Dtjg3SEZUVBeNJoC/H5mQN2C2AyoCo5A08QUn7i8XX2qKG+DZK
BJ85s7hK19NBQ+4mmKs2OgzzDghDVX1qh1HY3VXhFGf1a/pCjhgaleG/OtV4
xbCRBefc/yrYXI8N/6AeoyH6M2vt6d7yVhN++xGd019HdSET3H54h+7QmlGP
Is/wUnn6Ez0peVoA8LGmw120txTuMJ79XnUlX3j+JcnqUMK+WYXKhb25Cojx
nOi6lot/HDhZIm9WwbagMNpZdlkVP4fjvIhng2wd4h/MMDgYG2KpS41zGS9v
EW+nZUr6cBRi1jyNf00EFHj60guokUe3Bb1uek67U4OZwF09qwdGa/b+KcYO
REdXAzyeSxySw3CsVOMstM165u2L7DzinOY5pnjjuiM9uKnosu1KN5vtoB+d
j27RBiHwINkSMiMbcolfsuuBCMEkF/kIWI3p/3zDNFKaWW+zZmt+gCVCTgfy
A/UgWjGLa+BFI1+qS87xcevElyGmRYqyx7i3NXIxUZya10eakfS8IZfLGjTp
K+hfBL11yewwJvCUSgk3nF9BFXi04pGCFLRBNtUHzlRDurnL+lnBjsGjPICu
IZfuLvvvcwB+zpgGHdklk+iXEFWKNW13P3HxTWFyjacH1tqh6bbRsy5A2dxz
3RX10sn4Dw06Y0RslEnUPqA+t0aOinWJI2ouNABtw+qZni/yICSTjGSfGZIW
/EBaLgZ6WG3mjacp3uZq33D4Z79YeSv8z2CBTCxtvqtZG7v9J2G1veBJwXcp
yhJwDrS/DMiihUlmRUR2BSsyhGrn4/VaTePoILnUSoOxLMXkQ0xfRW4ONqLK
uQxp9r3jhBKI6RH3tUNjg7lGqH05BgpdV2Sz90B9Yr4A4OOMuMi+juIKZ34U
Zs42/kv1qHylBvzug43X/fmul0R/2A6H14RGWwnCI3v6MRYXco71JvlbNS2n
8hj8cE4XB983KiH1yvSpiDpk361oHlr6PwxliwrHE1Z12loyrPTM+tXt/dCK
v+ckFb5m0Tumu7ZaiwTSs0eeWv17FKz92FdLqsasE0h88lJOZ4+yTffky0BX
i4u6/Z4JimS7qjODUTGEQCvdwzjCF6LGJI79WFr7hYnc7R2pvD9S76XHokq5
19xXX4VZU08Qf790FwbtcqZw8e6rehUEvVQDajlGITztF8MxlMuw4idLChU6
AF8d7v+f5ptQdgn5J/lN5YZAmre63y2S3TPiQOPZaS6C3vjwVltT0RCVNhhC
AqpPnzD/55knbaM2Zglx/Jy/vDyPCI3Am1N0WDouVMo8XYBPxvjRohotChKn
pdZQ8GBNTrJSnjVctB19oqSWPvKGjrKTLtFrpoGipvXvUZay/amdztwkAVqJ
LZTmAttCaBH9FywFrgUpnVmP45zb3bF4+wijUp/qbDYsYp85za+WN5s37CS0
z2D3my0x0OJO1XcrhjxpA9eCAWfkkY/d9dp/Xu79sJgt78nHtcgHnLdmibzh
7/wMSLJOXIiQy46ZeekNohfnkf9rRDMaudfFgoh95MRD6cuVmQo675sI2Jbo
EjnDo3GBM3931pPp+j9GJi32+mlkBf1zP5qU2s41/bjJ2cZA3ioLE+Gi8dT+
cK6ghSn8wuxZCoYFKii/IgCVvf2dlFIeBm5BsIj3FY+C357BaMYDjnhO0D6o
UtsjxUWlPEV2C6XnBtcqpIbLrVjY8YFpXBtUNzp1wvfHTmnM9N6n+/whsf/y
SFWNw7PWq5YlR1TfACdBuN5kPpAiUizPbdkDSaF5i5tO3uO0cWqr8ySltl8i
4UOBYk0Ta/y+yCDclW3tq2Vp+Yjr3XH4BvcgP0d1gn20fo3ipzLiwyFv80m0
Xzp+OT0+LvgxkEAbxXhSrPab3tHi4H8q8E5S0epXXPuQjvJU26AUCwCqw5CD
ZdGbnr6MRVULrsoI+jDtHus42Em8IT6aBIPEuxl/1vLmNdmub14Uwi/M1D90
lzbz7Ixd4zjR9FH4uC3zuALFbfJYH2PajbKeGAoEeH7Cx1j1/8xBVchZz0dN
/jRJgtIvKrjr2gLMz9wVWGnLriTSKQaxptMGSwumPPz6qNeIaTmu+1kRaPxs
xPMKlKvvGCZC5r0NVuhlN/i/rjLLSLAqz8RVvbPMOz3rj143tfPDmsEcz1bu
HGht3HwvJgyKwm9FqpxPAOCzjh7d3HaUo8SFLtCV8CsV4JD1tY6AT8Z+vxgf
BXfexf1M7DT385DqzZwZIhiS5stwMjZAkFPpT1leDzSpHWyoIvX4o4br/vtb
rEjEYFkS4I0/0bXsS/zos0DYzrOjRlEFX4cLw+9nBXCxCytJ3ztM+D2gIxYT
eBHa5KUk1qLLtg6L683rxvVATp0n9C3rPR+kHweQP5Vm7GbiiC8PnkTthFon
FSJzm3IFyeq8NgP5cZ8n+7rW8sBLClsoS3VehtwUFI2Sv7XjmveIEof9sseG
pSG5X0LkJKC6DWFLDIf7a3ArGDijTRynd8rRer6+iwewR3h3WeMzdofsSrCE
FBvWh2hqEqJBpKMOD0pKu3RjEUa2BJiR7QQ9VAz2NmAYON2O8p4THf++uhvM
vok4kx+dIWctQcQUsRExnvcIlodXf7auEW8Buj6WeKUaNvPR26LZ1TWjsNoJ
NIniDJY0E9BInDrRgSK674D+HuKjelYTKYvNTUNBo0j3fuJ5X3+iQKGmb576
80454/mQJn0er1OZx3Du0OOgT0KMG2/xGdBwrHckjvLqTgtRvPpquJwQ51gg
m3t15f+dw2PwLQTylbatgNB/W8L2ATTv+l+04sL9VtPe2l2DhhVBgS4DzbaH
MmXhCCXuTW/H9enHXeXs9+P/lnMWZaZ0mmk69QPadT61GgFSX6u1YPte0Yyz
LIsHNoHYCcIBwjnS5tMD/mIcu4F6CfhH9DZFjaK/xB3+tpi+5IlwrCcs2SD0
0xIuv+kEh+ZKp79DmWPKECJvXj2iJL19prB+P+LEzIbYVLqHDxFVwLjdBQjG
hC+ELC62eYlEyuOTo3cUk4exQXfP7P26FCy7x9i79qODntynqtkZcUkxuncu
KiTHkrau2vg+0p/c3zaiVHYUvAwZcTbkO/H37f4hna1SSdZK3I6mU0bNF/Bx
c5agMey3nR81yyhLmov48pMaXZQ3Tyto9zyMD77zANUoEW55OYx4O/8na+Gt
eWf95HXMG9EnPBMyzuBsh78v1gyw1eWUROy0UjKoQL9X8lFA74vaFtdBS9HZ
EL5Ndv0IBh0+gfan1SrbFESLwT9DDZi5LiGSCs+90+bgM8hiHTMLYSii8tD5
co//Lp5/3cJjwbHswEMQFGGYDFrMpfd9NKPBrZD/5i/INZry+Ox3O97mYkRn
mqHJtRPu6Mcm4isuP3tvm/ZCMmHNjC8p6GQPjlm4OU69Zf1A0xoSlEmrQZ8n
a7HpQEvRQxUCyvhaNbJ8k7obSQNRvDCDy9AJhnqAP+IuekrYvZ+akxhQNd5b
y/Fh98ibKPqts0GMQwnTh14O33UwlkcTdQdvC9VdfVySE4DMuJ/k18gURyYm
pD3Za/tdCOq48/leza+9rW37DxObmZaNMb8jgRQ/1w+gbswZZoSQiXuIPxvc
MjF+gh039gjVOULgIVzMcaQWS/8z2PJf7Aviqrpx52jc9P1h69ykgwTOUqP0
iBEEvhl/T0ze30rbFtSUMcQfOZ/bVLdBBoXMnPBlK9ExvUi8ak5VEKIgG7cL
yYFO4ckwuWAlyHiLOrBhxLjhwTw1I4UGXtA13FIbTBkfNNsCV1WjBztjfvY7
+NKILZO9/zHG3J6hDuTHKnYTPGou6uQHmWurYgofi0WXDqCTIOjaA+7lWla+
UtYzDZ39IjQinywRNhT95aZiIWmtimTBm8z1b7ul3Down0GVE8R3nGnP4ky3
2hQDuAXv+LWJThtIacB+ER9EP/w0lI1r8Y43TnBOWuiwKCWT9FGC2ExT5kix
veL3QPR4j43MFs/K9jgBaKnAAhuQxRcCHaUzzX8bNwGcMFh7Y936iiRIpSBy
ceWN6DVPGK+67+dUU8EUzzC+fGn88IyX8aVT4QjCWJyH28SgI7UWxwN3Y+sx
ug59cllcXL9x83CTIiowfXefa+j8HgPuBN2CgOxIMLhqR+yhHodlk9GnNcrq
6dE2BcIeKUWZsGunvhJKZ3aoO+REE6zZXnQZkhC0DpRi5IAJQEtxcxumrHz7
olDNyiQdBVwo32kM7D3/EZJXe4cJ+8MenqNYT1DCZi18Tb/ynM75Oft25+W9
/iRUZcPV09OZiBPwHXuCpdlti7GnRaszdfkplYfZ+YHmKxndrP5F4c3EV6xR
Yg03GWsTCczKLEUlXyKNYPWxrUTogH0HsxnG5k0BwaB6FX0KNTDawamIcx32
Y6LHylHi6oyNgPXeVIa3efn3KihjgYF0pk8fqA1iZB0ztDhOZngdKmpLsTiD
FwisekSqDLyFEadHBI6Hw1qHBQbCeZwDMnmHDAfJ6A8f6M41cOUmhnFO8naI
oxKI9gnL+i9/9jj+pn1YYYSMf01Q7lLF5nGfb2pTJYTmte1z6uTkGaWL3igz
1Jvmo3MSNj1GzWumEXIl9F6cDBGcXvkV6cDgVmhJ2U/sgzAsjFO5DZBJwECz
hJe3I5+JNrn7UztwGhQO2hk41CG/GfkCsNxVzd5pcNTY4ocrrGnfry8ejF3E
z0UO5xFMxz/JdRgZUrJbLfSAIXMrBzSZXL8kvgd4TBgnQInFQho8NdGYc2zS
fqk1IfPGHT6WIXccUj+CCtguAUbcQ24ICm1K2In0uGosLBmdQiQD9yzl/p8D
+SPB9bvLijpitykv0J+NtyoAASPqsAH+bPxpCgD0IsbHPibwUFDpyUxcTvd2
OIEOATbmNFrs/LLx1R4qCt83OLLa40oY6/hjWOxPqKI3zHD2Js12j91B6TBc
j3YW11m7cLBCXebkK5keGLEs29xbgjheiSZjwqseyJ4SWS3dpL0pwcTtFM+K
edUeuCJE5b/oyBbvHmAqlJtOQI6D5paVi04IvgVmkQAH3g1vatsfPC1Vqwft
gecS2At7o1Lxf5NAANgNGePnWqGKlbBjRUq00gQI2CdeJme3eGWvHlXgXSHf
o+9UmhqRwexTyZfhjbto8Nh1F3Crz5g+Ejw9o/EhbqDzznbYXmokgiC30Kps
nl5+BMM5OeFf234Dj0d70HMZH0ZPZ02ZkUtNGdOd1S8D33Qslc9d/toxDeBp
TGjVtRXyQSq5k0so9L2HuR9WvFnQH5fyOnXHCHKnSfg6P1abNRRzAbNukuGJ
IMDajLrzsnTRcqS6EvRYMsBhTPjswP3izVh4On964a+dFAUM8nPJN1aGW8Wv
zkzOnqXel18Vr+qmWfHivErX+IIeVsZT1WbCHwljAZATrX/FOnNb5o0ZRjbx
IKPvYtB4oHdXayArgis8agfV9JPwxKIS/0/AhYdpPKcHi6+aJvu1gcwPTSDj
HMTH6KmxMBEAf0AW+XFk9rXLTbjqMEzMoQx2NfeKI4iCQYB2y+ifjPSB2EHW
j0NJcXtln+S+cKE/9QLDeyfCgzoDkilqkpgHMAgNI9HiKzqT4JThvbcqmgxA
MX0+POibP2IV50+7XGk8ycBf9rziRnzNQ29X/sA8ElmBZ/uLyS3DRfnGqSme
Ghu61gdq2tEsVELaPQ75QK3MIixQ3mFy6Wo6aFVHhVhV36SHbBGpuWs5F3Kz
PXevMgZ8IwCqvkPJQ25oDusw2/4bh2XvwVAajsA7bHlzR8ikp07g3VtGWjqd
iP+Euu2kkx8GJ87z7g5UJFPlClwoa/u5wBS/BT1Dbo05jpHW8OKn0iJ0GBlc
HZT2EWJLg5nath2mQHQCOa1U3CfqB3pv7wtZwBhJ6tND2CTQEURpL1ONU8Sd
1PWRJvVvItBMWMOnTldopoEin/vJieSYs8IvMwU3+5mZmsyHJsYcYQyChNGY
wwCg5TrzprPIn/vas3czh/arpP22eQ7aqfibS1cQk4D0v/c1hts8En2dsMhR
JKKf38w7dizKTAyqXaKuX/H8/3w3DAyM08N7SxPZ/4xKc/XJA+vnYqypyC5z
xWjSyi7tTDoDS6FcbmyEciOFU///cM4TczrjZBM1af/mLql4X/vCun+sEEDp
uuUt3flDnlmCo5qQgYNvdpBYQe9cUTJu2BXQlgweVh5piZ1B0RQRBdvBgOU0
yzB5gdLPExz1iA+XvHpaQRLKVGJY0ApSPFhn8WiNRLyXUH7Y03rlLa/azfKs
H83XV5bOls/XHPCmi+r31ltPaONpNaVNEhk17dANlr5kb7Ebqj9uDWOFnkhV
X44gVFqpIn747oXzuhGBX1heulUF4uKCYOME5bEsMrlx0MUEmM4cOiyd5xDA
6/vqg9lf5z+UuZ2ZUjuHzmWhOHzd7ZjnvIs9+ITz7kDSy5K+nnPtrZe8MAxs
CA45xoEqvtwDrcdaJeMCxOVA/RXCyU2jLOswzpn3C5WpDhSjX2w5tL/0fMwR
ZrEH5k3x+KRU2z1pNiT9AJhW8vIMxlaNt94lSU35GfA7wn+E5/CdAKQh2yuL
kwDH2JmUorCDhC0K12JVGENHSvof7LU6Wa1hYk4Ig3pQUQrcGEiWqntefNtI
CLEQPqmJkE7nXiGXY3p5PQzOXZnyLROzWo48zHtW5YJ5IyFeHndtzdFdwtlp
uaY8s+6kg+pPRWWYuH1I+lNqCs1bX+UY/GUCFt5QK+IMgZ14B41EPnT4hnEY
E74GM7cUOJnk/+R0TtT0nILyEHM4/I5BpDX7vmHNjqZ3AtRHl07shjAQoUpx
76JxuPvq4lp8lotSLFXrE5lkrCR9/H9HjhZjbJoBE1FivxspIs6yRUTXBqiT
xU8uZzHgaN8mpWi2l3ynBEf5CPcWEOIw3nlTQImDporgqWJLnZTj9kldEkFG
6F0rlD+GvNT7WfcAXBehu6vdNo+WQllF1BS4BIbaY6RX89xyRJev4tn+Cpv6
ECyIswFAtnao7xm6IEWKV0mm2zyjh/50ZoJZ5YxKzQjG5WNo+sbNMuhOWnG8
YAVWaHgLc5qHgUqQ67zco/KELhXUVeSvkCYEPHMzSiig81oA5s9OqTWNFtdS
z0ZaYeAWRF6O9qH7TyrHofwKT0oPld2PX5PY6nLHnqLEE5ffnyeqh3TEYoo/
3GR3pcxbW2dNCW2u80FCLEJKKseJp8kXwNBZ2HTM6clIUt1F/8nPMOVc4TqQ
wwajkxmb5h5DUOYNfiw8zCoCgynjufwZ2k4yxjLR/eN8prijRDTsfeIJOkPH
J/W9LoWj+r4AmjeutQdcY9DjSlTq4xMomgMzxR8/OkYuNi8/WqKXmt6HfE4r
91kcNW4NeI3YBH2AIhFFLXiAY66jPPI6MWB10R/BUtJ0gtCOxpLSP1qbmhbC
ulCM0RHNNxvVU7388y+a1LyisBP1ASRRa7a7LQK0KN+vXAgeC+28ptCR0CMq
PzBurKoQ7c/Ika1futitoeXefbKge7aix8zNLBHeN1biIpUiDPzomcenLC8a
pZ8TSj2YXqbFkG8f0qMm7qbA93T1gUOfaMWTPa0igxkWB/JiZOpomZNEYDS+
6J2FKm2B4+JqbvST7AST7jcm+LMAH6QX3Z8EvoSHo4EUy1wIWfWpydpNRjat
VBJsXXif6p8JwW0K7J6wtSIpRguIj9daP9rsIRqhgBozv71u8H+u1FVmtzq2
TTUv8sPaiyjUBaCB8PxvKZYnkwTtGo6IQvA8SGAgL8suAOyAPqS5IDFArEWc
gVALL4P9m2q3/lX33iGJFHHaATMp9+hd5PqfJkKXca5hLgQeaMFND+7e/Wcv
fpEXzqcQYGWZl+vIzf+3MLTE566JOVLtbD0okDE+K9ic2yLIk77feqwKKnBV
Eyq0LTDTYP+KCmkPgvsLWRA88RHqgklWQujrQyiu94ukD1ucD4Nis66UkRKA
OQDriW0pliRCLDcoRFFY3SMbQEqQ1iiOoHorHAf67APhBAnW4A9fs0FnqUj4
iJTdN133CRJHUcT5Xgi6rDUygHxxifWCSDtsnm+KdGiJ8p+uaXltzxYFtXOi
CzQbAakYzdTzsUaQMybryxFYBnpKs54R+KoWXysOSHCN1JqItveZLo3hpbqG
7Em6l0BzHxER4IICdm7Mba5H9IVgaqw2B/f6ozR8iZcTliFnXZXqZN9J4xWl
PC7PPAbJPpOerjZRZ2CXgfZe7vfqfSvCSxHQrimqcOR5TT4IksGmQWjCUGGH
/9BynRvdFmemxl3yDlk6OTM2lc6hyI89bzD/QMbF24f6yF+VemjXT2Zp7503
thsOPZQgPuFCpc3gyNxyGSzO3ZjLMXrtQ0L8i0oK7n3Qv8G/NU8Jv2NAjJaE
DSYwzgVvkVWoenDud0Gm0TGzme3Ovz27of8xoqoKPIEU96SiizbWjHd0d48K
1AqBmOysZyLLdtCn3sDBp2n6uIfMKoH5gtNiHCRvOR/mTYq4R0h7hjczWM1X
oefWda28S6LWI/egjjLUd4VAl9kYZ3fFh6KmzQQ/FNbE4Ir3ErLpby8lh+Fz
PV975Wf73wr7chfq+5xCfWe6Br0e+4rX1yXhPGx7V37jHClhtlIUyP1av2yk
P2x0A99oRd+smDjXxXMbmqrtfCcXc/Jp/UBOCyh/FWtM1cqNccv5q3QNo8sv
8bf3W69/qIz6UbVVUz4osHc+p40jLMw33PsWNUcCUiLGKLxFitPJU3bjXcqk
JmVWWdk5ugeJXpMogb7yi7T3H8AjFL+NVNCNog8//0TitCdl408i2YBo4CHP
atIPNwAB5XF42GRH4jVjoe2JESljrNn5MK1+oIrogfFn+plK46UHL3pO0Qkh
GlQ3f2AM76UkMGKc6GNVJVVrB886h4NXcn5ugcOiOWlbn5nGiNagWR5eTcdo
aY1NaoZ4izZkD1FOuuvUsyjaEF6LmIjoryfuoEdvkBVqWASXlUGTrWXbmcr5
ch3x0kPrIgX1AkJsVD2COQbaS3q2yEkhnD55mfmbqTCB9QXKHJY05mHoTDaz
WlBRiMJ2X89vC5Md5NoTQ3m38dZ01kz+cAX8b6aU2lvCHhNVfHEgMUg9+ctW
HuOri2ccnBPh0LVtylCVFFzhi1eEY79nk08tohwU9DD5ltdgrUUGOAQBlagx
Q/TVraB2/Vx9U5NItAnZWHZJ5LspAWuoM3pLhy/JQ6Bec5zKvTwM0UbmvuF6
MGXMY7N4x7OkGEpj8yYuys3Pu/+0ON85TIb7Zvd1Bj1UgPn/LN+ez7/95BrB
MSsa1VQgw1iNWHUDPe6p7W8jBlobCNynnoiUX1qPjbUzf4AOBIO1wzyPrzrh
esNJ5lC8J5OWZunf2cCeojsJR053tH8+7IpvZAQfjtNOF0fPPQw6IZoU4upT
Ddh3cOFfcFTQhSkL52VsQTdXq9j7Ty3qcYrFMnTS8HpmML7Lqdk6ITjCDNIE
ng+kut5jzYsXTMd6v0vUuihVQthi+uq0K4jQkhkJG8vFc9di3V7QDh/9iV0I
DKHZIwDi8FdzpHXTaxxdvaKLa8KO4bogajvue35Bm42F9ePAfjt+YJVwoCqp
OiJmPbvXyfdMb9kS6HRvUvOrW1vl1uGdyZJopqpV526eWvmvIoDOPQRZ4rG+
8+nWZnnuCYfD6vuwI9mbLgmDTt9hduQ0Wu3h0s+4pduxAouc+zBbdftDXBD9
+GDLs0mCdtOCDEpVtAfQsS6YFgjEKTVvIMs0+WeWitCPc494RWQuRrXwdv7O
XNEsitXtiR/axcjeiyBWAiNx1UhY4sFLgQxxALYyWtzCDs1pFMfGWOTkeDBj
z9xJ0X7GKn3Po2D7A2mEYZo2z7WLFHtKMXjLVERq/eQaUCjnSHg/c9kHyG0c
GqvNbV0Lxy+4t/APG7pLng92J5az+QddZbMZ+dEdatbjOT5KxokGwMEmGoFj
v40uiFfvF/w54sWVt27uHs9JKimLYdbuxr1RfP/e0XYYD7Dn58iDh14khNf2
+ImQ0/zvXOwccQh8xhCJrMfbWd0IAHWGOI3d/jdvFyfU7upGdcBefquoruCj
GbGvLj8bkxoJsM0tBY+hdd7pZlIdK8xdLuho7uQl5izy0cUWPjRLQOATcuOh
IBUL6ahyTdGDB0KM4GopeOBWhPxtyFbz4C4Lus5S8x4PVg0APg8ZtFXXtLhd
a4j+d35Bkm+4one1W/yoRV7PmV++gxTj7B7wkIaHvwjuI27a8jiz0+ZsIzgh
c052gGkIDc9fOFzWAhE17RtlhcgRCZZ32gd9SBDND55ZnWjuG2ULiYX4JTWY
MvRRv2XoOEYmF+b9onGP7odaBHVgJgw/BQnz8aIQjZmIPMZwMv8R4I6VNBnG
lBWanOMM8kRJnL04WIUrLYCGR9fIIUGc2I0j63ufqL2CzWcpIyPtogp1pxvI
+xrvImzDS72Hcu6Kg7TNNUdjsRO1rtJfGhpIkHxhZ1gTIjy9fW6dYzG4lQFB
frslveGqndHrknqqa3UXCNjPelJf1tJ9dzrW9Tcz6IeVnSisA/FLHw0a8S9P
/XcQoNp1Ff2z+PopUlcfXSVi+3QsWMBEL+e6prX5yIM/Qnhb+evrhAXgv1YD
7C0a/GaZXIxrWg6N2xX/Ilwm2AJTv+EVU4kr+R8kJMjPnn5OgLwQ+8CkPxQA
jkPgle+7BxZ0a8DdTp/aciYPTYLE8RxwQ7cDq2LvfvluI++J2epgEUvWKF/E
Rra10d5VS7/QxnJIku2pWHQRk4ILmAxNz+0r8qRtAIGVkKwR6bMk0kS8U1Nm
oeZg12a0ZT6b5/kNWz11rXfS+nwm1tKJAlpK7/EJhJppsyW4N/qv/vX2OnLh
8MREzYOCgEIt9iEPwgbrkkS84Q4qrKJ0NXOVCOmyrrF4FU3+GaBxd0FOeCZw
pcLUjWV8f2JuB/qZ16MQUDgCqwwsD91kEol41r0rcY6L5PRkAq45zE5Q2PPa
AmicjIV2AY8IcyZc+2ML+GO/jWZSjCWFRHCCp4kMVL/fvDV4ZMB1v9v/lNAc
mfGAeuFmINgBscUgXnq7ikFbM1UnvB8Y96FrygzeuWoY/PhQ7mHRrElA8+mK
qHTnxQ3pVjRd0hEM5feU9KBvuWqGru24VAD1XH/kw2E4DAx+Uw00UWqfSX6U
uFH5clOVHftd9TEHL+7eGv6lIEtFwq+7hHRWYoCm3hh9e4OVRk0PeEk4QNQq
7xAEKEvEgCQEbaQr5J0yOciFRXm+oe+QR57EDYI98fv+PSJwmfb1ksjz1hwA
/NPRXKhkS8WlpVK2j4xhBec8Ov0Y50hlOHSMSpSh3prB4n06QRsj2AZP9w9j
51Z70TdpRpAu8zDBQaiuJZCq4tGHtGbl9VSvY5PqrbLHxRDaCQvhqCkqIDGw
18J4RWkjYFC7n++WwhGK7WQhgWGf8kMoHqxuOv7j2udojQ+WwET6nmM1HZAG
4Blc0jzjXL9LgKuvHuGnsgVJBkE9/3NJxSPdRYn+x0HuQJNSrbC69ASUGbRN
o9KM9+8xqvQAKnmKUFA51ybzyw0+GAE7iZ/iMHlSYSy9Co6PfycWLczHqK4k
fr+SafCjZjkJGTssW1bx9Iwn++zoFg5tCK5ZbruIWk4ExuKAhtqDiTDwx4k4
uXGBCfcZmLwuY9FMdoZeb/Y0GOVLei90Cpo4Jzo4bboL7CxswJAieQDfd9HR
00fKpamSoyRdy5s8P47ltfEH5/da/V7bnM19H3mNeTmrqrGxyfkGTGS+s09W
fMZ6I6/HSPuGuxF3deuLFTt18sssn47+ied2fkUzo5T0fLjBfnSIz9QWnaLe
hl0FfDJCUJ2Hgsbt1yw7Z7BON0YdczVGhEHQK07jHGEbuq6UdmejbQmCB8fg
A4Z/xM4l1Taxv5j+8B+BR536fxN0akwNZWkDX8isqp9cIuAisqo6PU2uc55N
doesVD1Anv/nRFwsQEtOGasZcJS5hzeezsXJbavDD/hXbO9scL0bc4b7asT1
d1dfBS3iI1OSRp+4k4GwOhRpLhvGWHQuAl7CWBToI0MxZIAUSHOqyLZ5rFkL
D8EklrYtLtC6OMvVu7dVsK/vncxIu7yuS8S35RQ7MGHaR8pc+Y2v3GMde4tR
5yPjgSUt0JPsDODFtQ2BP3o+wcGun80J8fjwLWiZQryo3DJEv+X+1Vl09n7B
Loa0F+EoZ8A1SzWmGEme3o7G2uZ7cOJoiphnspGJdOmrfwKvA/P8a7Ys9Z+f
LoYtwmdu6O+HIg3+Dg7oJMAY4E2zthUhfXS6M0Tzv5gcHKgfPjdboMELOVxE
WV1MyVwRC4CvBBZv4Ern7/ZCrw4Fv0gDD3zgigCytmbaH0mBOu0vtJk+aQzY
L+pnXLz3IhnEkyHEW1yJIV+z8Ij9Qx2Dcuw1gvsahp3xwdbtLRebybwMogiS
O9QGGvK+itgmkCKgsTNL7Twrhh5CkXUzkhTVShT5sZWuT/F3uwk5WddqOIrj
31a5sS5h6PdvM6sGKAYgMotGAGXKowAYN1hnHnfznZcZVEonNlaLxnBjHV40
x7fYrvg1YwzQezvtQxpYWS+izNBlhwrFaQPWS8ICmLH29XCthL22x9pG8j7U
X6G0/70ck1G3E7ryc6ASgXg1gSfiyNRqKPA4cg64ivcTWuZIPeN+XMyj+HNe
Gz56i0ztwgAEOt2WmJqtlp3zb+96+D+2+Ce+tGkIcaqrM51q7YAGYIatKsab
seNY7bQ7zuH909VaV9/aRnQBulyfqhgDBNkz5awHG7Bj50VSF8jRapQzvdee
s6SzzYi/jobFSGNkNA5JHnTtLJaYtdKq2eyBeqxbE/yNtKNlKFRnFMOd2Hod
JQs9AC9nQ8ZiGLwwW7tkkdNI6qwyIPWA1+2ro7g2n+hK1lG5fk3PgFinkn8A
zQWsRiqafQ0a2mHKPg7QuokiUNg09KbrZv4Ciz3v59wVX4dCbrFWo9XPGMNA
E7sgxm1jAbOAqL1LecF2TUw5wnzKPkgnkYv7Zmprt9lJRS6D8/N3X2hLMzZp
cT88INfnkvdwPbh29yn8rIVf9RfPoN5Rn5ran3f7AVbF8U2Cl3AvZPrCte2n
5UgeM9t3HZ2hCE3JTSW2K/Oe5rbhH22TVzNeS7C9DY+LU4rZt+FzyKpaqu3V
fUek+kNgdcw/BGlvepjmPKlNCq0Mxevs3zVVC2leX2dhjvlVMqHO7e4X3gl+
NY0GH9k71xX2Gh4IgAxR7s8TwLZCGztShW6tYLTcW+vXPrcQs2ujlqIvXPiG
feUFyyQs1KnLIAEEj3SoznX+8AvepG5qDI3bEaJ4LpWAY+NkLtPU2vEM1lQH
llH/f3Zk7TxXhcWMJf/pX34SJ4X4XjGNobMLn4byXYckgFWnKaeR2V/b0rkO
y9PRgwyrMcO3fuTo6v/XdtD3rjk4ZdIaMu7otX8b9NosRnwldPcekotlwAEb
pN0tdO9wdTextywQNQvQbAupErgBwRWM3otheSo0jf6rsviiU0X2xlReCz4x
FafTgOAF3fpXrblctoEy+/AigOaa43BysOqGepK9Z+0VG5RZZjjGtZvtrJOc
GrxQBEq+wPhZzScASehh94KroI+d6XLDzu/0QPC6Vg5OU4uhs8yTEZQHjZo8
SMAQKDiAllgfWx99cGlWPoYHvAbhHb8dsOaj8l8OtvMJfKfj/Xf0EddFb58t
gdz/6Eekm3kn7YZREZlrKmgfYc1yJ0RcfVgsDI8VoD0IFcAzpjuxsFZq0E+G
OlC/An/R+5aMioe1iw6hdYetnxHE5aNX+bT7SN7A2N2qVfYY6nbj4IfK2nUv
m2Onif4Yw7vU0IZ5UD7FOo9HWnVUiks9fsixn6Yyg1XoNUY0h4wIsZdWqngi
kzXKh2gijlrqbKNZT/346+yBAeAerJX+F61BnUe6RcyzID+S+p+5IxWIx6pP
hFqBNBPBLssNeePTzP63zBPaG3IHeTP8MLzFutG+YdJT2dEs5GxQ+8gntBcR
EtdwMhRRkolEY6PzjnkWc+rDAKXO9J+o2wEmmG8ESQ/SdORDRHC2s4z4dJAL
kC5vNmaPA0Bxl+QwqVumdHE+9dUQDl7aRgdczf7D/00GT5WdoVurXWj3GDsR
nQis1lVc6xL02Ty9lVVpN3JxRablDmLgKoajlgHbqhoCHxlHiW62fgW6fGfv
4EKW/RrcDVQupR3JWtzZutYHtyY1XNCn1LuU9BZSxVr1jO0Fuu/S8Jw6q8No
4HF0gNmtW/kDChsh/NvE02JKLm17yzkPIKsPcqkPKJv/X1qm9OGzuCE/zpLR
6df2BbMljDG6Op9F9EONVr8kPHh37tDxSD/s4x2ysh02fQaEH64qIB3/cEgF
kAATrWDGwCjkERflUmsEHgj2Lr/GRcKTKT5T7GTTtaaXw66efalDLkusxV1v
awIVDzRI3Gvnv+FT2YZr04OOQHAaL4B6NMaKdXQ5iFhmmDGGTksXwfxc6oBW
+hKAtu+rAXS6iEp468QK+4glPjv4GvDPnMAIxk2QHsCPV9/3ti1+4vCpE75Q
I5v0J4AdyuriXNn8cKj+Mi2+twBgQy5ynP8s6fiHAqHFc0q3DJ+QwHVjcgCE
2tg3rCKvTgspoh5bEp5WCpbLcYZ+lQNT7S+Qz2oYuzD4OwG/B221M4UBo7Jv
CqlcGhTiuJ3m0KbT0IEgU+imj956wiNocVHnBKzEkUlykTR7Jzb0aVZRFtau
nc1r/NwbdgX5/OpVkXWrxlCJ2ajNZLX5BKYXHhB5MFBG8VTn0jpzkDDluWJd
YuYl6egu07nlimwOEIzNNDIoHJyWDRWkAZYuQBgdGhoKNZXahM09MDiOSco0
4sDjvWo1GZ1qoPeKR7j23llEUnsbe5gb+BE+7+SQifrfy2ZMGD42LSeMRS2P
3ZJ6MVpD37OIdk4bBpt7IV/GVF9UXf/8s67eDTV+3j5UBZbetjVKwoY6ulQC
0ShGAEqvGjNal7MYfFGbKbgqAnLbjaAJHFmMu9DdYArPdrcwzMtrRIUPYvKl
4jD+wjcp8YfsutmqQER6Rbd6vfjaPLfm9zi3F+4PAjNgesSLRoHZIe1OOOlO
knJhH2trHkY05R+yfHNyJVVcFkO3Rdw80BqvnmJQ8yEXD3atkId+kHUYNT2H
+vgEFCDmkkS0ufytqNNcKDZsVBbveV22luX+bqg/DUjOVw2zynwYTxAwUa1T
N7Xz38JqHFH0amcK9dHPHcuRqVUPxGp+ZPCmbq36lzbkBK/QAFaJnWZEyfiU
3mqGCMalx7XQLvmUll6Zz9q705SwHqA5mx05iTaou1UK0sJxVyi2myA0ZVOJ
I4uKWhvGxIQRXWxVGB8rvBN823gGSKbH9aEQ40KqED5OrrFFs4Ky0oyVZsbU
ZQXTCUDwhHw408WJ2eYHtgOGr35VSTrb5XTRXkOyt+iRTA50yz2UjAffauFg
pMY0nc4of8lfQL+fP8uBmuoPK0qjkdzu5k9qxQINKpPUWuMRM/SUajf78wfY
ccEaWMVgelwQtQPE9mlr8UHIPPE8aQyQWtQXQlE4Vn9lcMeA+ntFivQtEZpk
LSe8/qBiTCF20UKguFrzH9xT3IUQkDrRC4XXIQ6xv30oDeRBLXU0yjZAr1a2
FEhu6ehDGF558PEq8gYUkj/wU1kcpiMxKpcwXUlVpX9C+GNC5/o88XWw4jy9
bcsARnv/0tRpQ3r9SB+au6QvVOd9K9G8x9gn7o6eVyuTHX8GEwwXbWidcwZ7
VwwYLeX+n2waelVwJ6q476qiPhEk6NN3loYa5ESRQMdo1Fff09LYzZQOMN1R
7HuFozmHqCuCb2fK8BpYENo8GVgiMeJt3owfNGHeeKj37xoVdwjOyN2DAX+C
Ht8Nf/d5eAaS+AxdbBqhFnpDP2+t2gQkjBbirHh4b/HMo8MF3Xw6D7mpvK8I
E7ERoD9e1b8iRDQwcHIAcSgOf9aXPJIu19tKyVCPvMmRnMS2RHM+qKRjC3AD
qLlrvVzkNhANRowRm3dXPx4x2ArJMMrO0dlXoaZ8uzV4BPsXuU4Mpao1qP0a
AfLkIYG3UlO/4YcO5+cvPvr5BHsEBWU5VZs5VGILrWP025fnRdp7evvaTwPN
RnN9nEmAamgo2hcdP68GhzrKIVhzH0+GrPANgznUdbKpaD8En962wUSweJxq
1ynvoRPa4Kh3x4JbiL7knXfqIc2w0JtkvMkIX9QGzPWvR7cNcue81c7/q6lu
C4/K2Axz/Y0Gymx0sGg7QWpiNRw4qIGWzbZaOgdO3KHLilfAEWEXt6uIxIgG
Acb/2hzsxASB3ZgmVR1tlT7y/Cl7eZfgQqDfw3lF/iOVVpcGDhiJVKIaSuXO
yYbMHeCMc3agtTbKpzf8E38ByUAAgwV1nfPPaqLgY3UrI+fGIulvXRMSHPRd
D97XeGMUsJSh9kYEyjbRPuw0ol1yzaE85cq0+jaE39KTwUQKxsl12Z7T6Kgv
dEn8WLwO+QNvr2SuSO4mM0LDHPEVHv1TRFf6/G15tC5vXU1ycfBKEqCbXLFX
2y6ipebWx5fyr9T4PitKfmhYRdVrkgnIKx+8AlSwNH3aMIDo+GSzBgRItNYH
VrbNZwQd99+F52rJ+QTma+Xr0v43+FF5VRukQUfqBVo9tC8BFIaDBzfa7V6A
AwBxXJ7dwi4jf5wMa9AhXpR0fjTFx5tyP4zE5oJA1vuQ9YZebbKI/nMNAi6v
7+XgSq/qt2OIOGLgAVb75tTcV1SnyGGDmvpTxba9lxJTNGgCJwJzPSO7fM4g
bdPdmi0mP8pCwfX4k2fkbTrcIsFU3u35xpwFqI5edsTckn9hHfowX6B9Zvgf
Fhwb5A+jnlNiQpBCwJZgPme8rsMwEsWok5LS4WpeybqjSerJQtXhXulbs87o
zPpVbTGtrjq1coMcDktpfDsU+7nMvIbnHR363JpLHjmIzsG/Cm9w2rFCsfVE
OkSQrxDmL8r4dq5le5mQ7U6LpnGAgG6dFtK6Khj7EO+DHswy3/3tUEP7hUEO
SMuzwXL5ftwlhbU0HjfX4AnCE60rC2nsw7RbcNQcH596t7XPdpWsBXg87SOh
SR0XwPBFCNrM95IAbo9YSoBHLTRQU2qtQB9e+FDP+miZPT/nzh4+ZV43R5+W
3fw1lK4lO4lxbi2Exyd7rRnM8sIQlWM6o4p7kGjSu0ZcZZ5aw+rbJwPY4BKs
yYWRWi0qFXAstsQomLcJhyC7UtxRmjzGIZUhFyEw1CR1mI6LnEf+FODTcy/S
xymZ2rm5OG2F5SrRu+chEN/nUBmiMU9wF0iQLh9kgP0o07W6mczm/iAyX1wz
cVLka0Ludcq4BeMV9Lhd+c3Vx5u3lJclWTHGs6yKIiFWLggkQvlh3rdMLM1i
1lLuBL03Zkt5vgy6+sw1mDAAYRm5rqClSuLKZWpOQlmnphum93ZzEA8w6xAm
SP5G9oXpYcXnbzJhbgxerluwhOU+iZarRH7jU+LZADWa+ufsdtfA9nFh5aky
gHPi7RVzco0+iAYoVa4iuVS/gLgaIEJvDk+0kul5cL6BJZ/5D7jFHvXuFcT7
NKOW18gYJHJXLCl5ylRxethKX7smVy92iV8hRUMFAJSZvoRiEuz6ruM63LcY
BYW/Rhyekb7xQ3qaUsBpWlXFxhMI1SoFWNxvwhOchu86mxEgoY6jNx60AWnb
scd7qKpbcH6hSslJEBNEiWgfnIh1kT96HspPmsvmAYYbJf4ljkQgOtcTnyP0
t1uCcBeDSseW0bhFFGAlIfsGGetrSwkBDvo1byJJwpqdx1FvwZbYMzhmafYr
as2Q/A3MYtl37P+ijq/ie+83rg033eVkM1s02S2w5pDsyzRO4/TabZoGR6mc
xBA5KHRsw+7xW3774axqio0NdZnedBmC1Ss7d1CejdGZVwgj69/8ruSLI+EB
HBt+2KgNIdP81XoKRgPQCaO/bZ0zkOGyWhjw3SqwWubEhucw5uNLbVSlehZD
m8X9E7j7ejYeWn/4JHFrR/nXPOiF+rayGKIcbKbQoEgvbZ7O90ezoM8M58h8
AK1DJ6dndbw8zeGvkl3HNKbkcUpz8SR2VNAdMZUthlRj9JD2tr8HC+k4h3bK
TWPTkWf5KTyj0PHZshPwwsopn9rduo5h6DRJcmDZaCC+L3DvUyHXUOKE73kH
K9C4qg1NfLRfFL9b0BBSD3IjtZNA/PetC7GjE2g8R9gtZY+xeOfXDC2YbrHa
GgPXhJGxjD+kZPfWHxy9+884gjaMfG5EKKTIbSPNizqcHpIrig+inSNGq4Ql
ISKOD2X0Y86n3XeKtOxurEYOC1Icw0qzQi9rnfIhGu48EjCVscl+4+S/nGfc
lRGslgr1uaUNFku7fwJeTek0D6PsokR3Hvf8e9v83W0LDAEFqeQj7MenEN28
PlBaDnyCRIoBFjkjw3KzOTH81seUMrIuU6s819sEz7rSNaQo8ZwewLzqSGXq
s+q3043lKOzWX8Kg+v/h3dv6zJPB0zsKJLKgiklqZoShq5YGf76oc+gGKnue
gcQQysebuq4uTT+4F6Jg0EdKgcwDN0JbqWinKjy0dg/BPJaxGY0r3aALm/ei
gZQsSN4BxKzhZgq8z/Nb8oypJSLhxilofjhfnpLZbP/591UmPo0qM2qPF2FC
o3XKzHmRuX2aqHyKvZidi/WosfQ229bg17XWQWwK63XAift9mtG6nPtyhHx8
3mS25GxU8gafytpQgNxPKWUXe+iez1f8+VeC8sjzAjEoCg44/HBQIYtK3T8v
OyET9PRzuAr+VHoy2jf1pQ1EjHfn78BmUe/OS6CyVbFQ+tcbzh/S3EEObsX8
WIXOKIIp6xhaKoaNOTchCiXBdmAArUURohJyZL4OZOJgG0wea6+JK6/y499X
VdPxpCkReqHscOj1bMP7fcvUnrFumTeDx7vI83LIf3BBtRe5GTNmJU48w/q3
ucH+Xuy5Y6GiE8lQYjKUONjUscuDLm6Dmax2y0jIipMosd7a8fESwe707D0l
HvV8jzGhGutGjyOhwJEX2vkW4icXXCsN3x375rG1jNPaDBHuNNvQvijt15F5
3uVicEfQZ/yCYsv1DZddXoewHhJaU/qRZPlKksUhq/gLg91aMTmY8UjeHT8y
V2MJHciEpIM+AsJNlfDiSCkuUJpWHqCjsfEB4oap461fx5EY/tsBc/sk+9MQ
doTSttd7eJt5CwN7hTu3VfkLwW2EXEMJ1SkGkTNQvtnLiEDvehhAdpUbyZVT
OBKlZ7WuZSM2P8802ANHx70zxisOy8J194D2/ijy/7P+nzbXJA16UQVjbup4
ROR/+5T0kjxiySGqYACYwd5ixOOX6ZEZMp++54ObAyywIGb63WnOBI4poVst
rypTlAq6gVwbGZ02IQ351Y8f+ixujFPHO/gvsAJCXzVx//HVIpriOl4P1Ogn
f3I/gL9reir8syshpUMqh2O647nS17Q+5tc8IgF3iug9kJk2NqUkPHnX1Yzu
0mHRtgfgj/XmN1J41S9LJBIB1xCa/O7GEKyhTZVyQ1YEfgAIHBDYi1NPj9br
K3t1B6lXaHKb8IyIlGzqwIyU29+QOPd/9JwA9Wu6cLaaHjwAItkm85wF1rfU
cNtqsfjKlaC8hF0YR/qM7anEmIO8xBDtHncdSWwI9+Ns25920WEDKMYLYxQz
th/S2zJYCcmN2XX3aKiLs5TNHGjI9xLqQRStvYgTKkVw9UYfQ51cVdwMsLsA
nO140MqosAz8ViuoeVOapBIxtN4aueHzXwozxswa62+X2PNUlQJwzin8wQuv
aoyeCYP2RG6jzGjKYS9fZ/FADqlQWA0+t4wz6ZzlglT7oCjd9Q/p2QbIGL2Y
onwu7hlUKgslYDsl7QbaTWfdViRljA+pp/S/C3VzeyCjtkBHFbEANYcoOXCf
o5l7NvZM8aj2Iw00DOZGa0rua2O1L46GD+tmyOLybnGWjNAE8i0CKfR5OizE
9pHmrbFlS3VJ29TzIPBfFBsIFBHrrVB7eGBUc/5PXWYyPL7A+lwos8oKHL5e
Kod/I0XWXruX3PXp2KEneoh854fzVHM1U+EasmxQKKn3JFV/6MJO2fV/bniS
3byTqWZ1SVOju6xplLO8T+7diY35u81nKo2RAIodDrAtuhrOpuzVEFzhZae0
6641B+O9Pj1cHKtRdlw+EDYKTh24gubBvNcVvzaXdrkTAHKMGSyiLyBNsXGH
XC7o7uLdPAQtc9Zaz70VhzJunvpSL95xNqISkzLDXKwr0KfmJPMjDb+g16ri
PrB2BxUOWLBnGkymiOByOrH2hxv9GuLaXK57+eb1VCBcNVb6d9wmrbAiwPIu
FM5ui5MdbvLSuNjW5/1mhZiaJaZmOhsd+3IFP2tTchsTTf6LK7KIXdD17zHU
9zceMbUutyLeQ/GAhkpMgc2y5FmojhWFRiOI2qHqYE6WowFGrzuRcSLsIx/p
oMMOeaoofCPlEahpDjVGiejuQ8JNVHihowto2mEJPcsC9lrEEa9otD2gogxp
+bKdrNdjEsFbjCqUCT+a/l4jaUBhXxBJGmf0yvNNSLgcDuxxHnm1rhjFvadi
tHZJ3bD9ZZc0GxQ8aTYzdE0urJSaAGlqvxG+GY3kS1756AdAJmKJoei8ivy0
geg1J8r8DnLzJ1VeHhXOSpXsM/bVnRVDtUFstzcPGX0NFpjhn51HgyRcg0EV
kTnRoICxtlzqQ0ZkctQGpOSaEjW0Z3jhfLri1LnNc86rB+4uRyjlQYixbEp3
jY3CPxK01a2vB3qaQvs4nOFV2R6zucKwMcUj1sFeCZOez2qEz6Am9tC7fUZX
objN2s07BvsJ+alW2091olbpswRo704+8qA4KfnWA2CmY0GTzFHkkRBBZP5w
XqxDgJFDgW0Z8GfgyXPaPbkJ0qFGX7IB0teYlShcf1uS3Gch5s0W9fEBiDfI
N6HdDLRScmQN8sX/SmwGA6wIcya3jh5aS+EvRbBa7s1ntMp8iLKksBuPVZVc
VxvzRbbzMzdAU4pPrRr1bGS7v6gN+4Y0MqUH8/KKDVjVzaNFoWTv/yXqkf6+
uuZgWV00ZO2EATa5zAVdyzJoGPS33xm5+gZKaUDDGA2kFYXrwVf5carsZGxQ
qnUI6sI3v8Ai/rmnhr47zFHiOir03ZIbLZbagQIbw1TUJOtK+zAhzRyi/huU
I/JMmIbY71zLzAG9eI0JBe1hAp6XYVJsy85bJ2yicdzTDhL1at5qZ/mvxLjn
QezFZGSsDAZevYJ57+cECXlDCe1huwpVTDp9wYbYywS8euuvUmJ5FOam6Vxo
pIwQhHQuKP/xrxRTDFVH29FqmfhATP8K+WLpGnl+zvVmtfxgX+X20cCwKMzB
udqlF4o7TRNHWW+Rikx4qZNz07BEDSZuLjTFC5IuZarCv3PekjfXiKHMkqWa
e22dT1ibsSL1RkQ/LGRltKSaqSWtwpDYbNbitsC/i8DDvrL5wpPjqVUYZHJD
/TUMyWPIBydgNrc11pOnWRFuiUHI7VRGh3hW4FAe2LqUn6l8PXc1J/+d0Mxs
8dIgBypMN0QqiTgPylP00gyVsXOicELYg7kt4flvjTCUBhcN8HWeLJoOJ0lK
81YhRwc61JOD99p7oo+v5sN5UU+PL3BbvD5MsOrO1cF/C7m6mPteLmbyp4Q8
WtZrj1JQ8uFQf8O+l+HxrHIiW/LWw7jiSNi4mjfn3SoK+xf1UXFbIpmbYtuq
2bFYOGovV82DePVtYFJYBSqPK2gs2SFEeJesxPW+K5Z89ta/vl33RNCuPELI
rRo6mRB7WOp7UYeFkGk3W4IeHtxq6yL0WW1mF7KQ0nCB1H90jWxr0LWWp6B2
Xb62YdxW5IANzF2HrCHY+N56GjPtRFlnEhxoXKpvU26oJSEUHoNaSiHfyp35
WEoE32URENbXIXIPUNYGWQ5q0HZxIkuZtug9qF9sKZ1vcHJMArrjMzhojYOc
/U2cCslue1EzkYbkN1O4haPyrdNQ/RaQVOxtg9kjCKgPH1XKDlJvs9s8PXGF
Rc2fEGortGidQt67vjnyUneYuSoNvzmEczRsPIZrzk3jt/2pFLjfEuiV9tfV
nQU1PTHgG+e6rnhcC1zmhA2+mLv8/gK+haMDCcZSY6lgbZIfcjwQCGIBGa53
Crr6bXJCT0aUVCqeEm8syiC76El+DMRSGSw0oWxCtI8eZsJiZl/0z9C62AoQ
zbQt15ibJyOS8hih+uzEVVCf69ZCk8XoIen3vKhUk5AMpRPa8T8t3kppXpwx
0jQ/JxGlBWPULt0t4w6BTNhxuMtVOewBpepQGdLGoL74xq2c6HVRxMjPCRJ4
mCGoCXghpjiPYhiB19jVhjRjtlAOKHfZwUEgxciccGFQXVhb96UfjyQBZD6H
kRA2/9NvekHv01gt84isxNszvWN3qPWbIAX+B/+q53A2MHSVI9VOpVFLzkA5
BRwdFJs/T+/vGnAm67+LQLgYwlp9u2u5rz6xJAiuvjEWxhZ5dB/e4/OXs0BB
aa4IxQr5NnTHFCnDr+D9HSzbvllbPZPwkPtLUyz0HDsWQYn7k6U+fglEDKhA
OZEam8tiCqCrIltVYX5bfgXR5Xjl0fEuoC2ero36LQqwgUfEiLsUrfntqoIa
YV7xKdUcfakIW3H359rfebRjPdfIERSL/IVnppeGTFXeMLr+6Nq2IBf0pwhi
K3fkBjIfoM7RKkLtgFHhd7qrl0NzHgnldzXtxL3r3IiIKBV8/gBq+4nC9JEq
QtrZioT+SAxcho/Wb/Wjy5w7mJC3HdU2ZAUKzfhG6QuJ2pV376Y4jl3DsLwD
mMfSxjs4szcGDD+vk8T8yxNfPLaYwuXakxb7xS2IDQGvlUYE/7AJhDTTWfxM
0S3pUaAFq7Ac/RdyuspIdHGoB5FZAahvJHzOh/tR+f8aBk2+hNnrXhFObskN
EecSCBEl/aTr5JmpdQ9WGK/xU97ARJkB1NtddAMQGDYbg3ifVizDemLhwyym
xdrX5a/RPcD1k//K0zS8xZwqtjebrxveS1wligmgfSCGJh03+1mhMK9vUIiq
YEkT5xnAYGJA/q89G/o5bKnUG9kvvtiVOyoa++EQ6KFP9k49EE8zjxbnUH9y
6/lEq1G1On8Ov2WwP6vXSeeRS+05WR4aBwIIsLjcZDalhM/lq9hN5sdCH4iC
dlOkgZcgp/zvsCJg5px+Jrna/UfP/myCRQLz13Bc6QCXYfXIFWUdrEOsDOdl
MpC32Fd+FOkRyOj/cJtwzB6GwWckJreXMMLRkvLvrRR32pzTdBxjTPR8mOix
Ngxq7929D/i5wnSbjgWehpFJRpC6A50YR/I3t/lkdOfd6DHQyKwtkyY+NG+V
wC+PtYrfgmywoCqJpLSmTN5UVmhtZ0ollZT9PCxSFivX0F/2cKTqGCvElGHx
gfvo0AUyB6AMih96nEl1Lcak48x4TkfugaYhHA7avKBwKr2KBrkVFqNVolMn
JCusYsGyvCsgzCJCiFk98t6LTdjxHJdSmDL9yEbgHi1FZ2XvgPn0YIYGmaR1
Z9a2k997O5uRH4mea0+06yImi2Vrs9mMT/K34TtUre6Xi7MjIYlT0MdKvD76
MHll/4t8nLS9H4iQ1HvgCsBEJtRAndzuMTx+fUWS8R26FUhNbX0/lIc2kqH3
0KBQ8exaCmsHl+uYnmfL0cWUcF25JTWvvrMRINoe/PLXhOs94hiO10i35WhV
LUYvcjPEGd3eD9tx/C9dGPlHeyeBBBPdNLWZ8pw1rBwC6cr3ApwCiyA7vDV2
iJGk6tFI6CYYRPtvTssNW3gmXm3sYICF1ieprO6GSbuAwB28HmTibI9GhywI
wu3M9TF5z/yEn8+z1/agMRqNpBSjLhhIwnIoPOB8qtZjZv0ySEZ+yv6qbx/w
PGUqT/nuFeEt9f/UKzgwxmxHwVXBdcqgd0rFBLnOwcypTvRnKG3Eeq1xhmjK
3ZtNLx59JByyD3KppXJLkBgZPBpN8jKpkrgrGn4wvpsPolUtYDD8jSE2MgYl
h0BBQZu8D8bzlTJ7GmY/sI4wUhrw9JQq7mcnCeee+WaFsGoq7vd8RO5YrjaS
8UzRNSiloHs70UwY/808bt5+HUOVyj05GaLJOs7HErojAp5YtYT/VC5U7iDs
JslzyfMZgh+4NEcd7iBA5BiL2sjkxJYxLOrt1kSrvcCHNttsb6J6ej/diz4Q
RhCKTts5dD5JEz6KFJfCk6eEDabQwSytN55C4iQhmNxD2QxiC3Vxk+UYlJz5
cKaTWAjgS/7uuSYcoE4BMmNIzu2ajc+MgAaChGqayQsWr5uK+pWkhX6hE+V9
2y4CPn0SIGkFmd1BpS+gbKcFvVhccQyihioBvS5mqhHcEmxxF3upq60J3u2Q
kmYG+RXVSPHrwOG8RpgEUs9ZTa9zr13+Xa72yZFh8wMf4ETFv7seQpUwxcMA
TifXe90jyk51uJXhr0xf6AenLvE6S8nnlarUZEIKhzgJY7NAY9cPHlBV4mbJ
4rRbordgxwMwvKXPkZzGej0FmOGHjvhdDa3HBDsI0Yag0E6I06WTZx1H88Aw
tYx4SJAfOx8HTN+K/1tiFNtNK0U9+vR1F1jEkC+EZMRt7uat7IPdG/w6Bo4b
tWmbYACIC1CXegkNsGiFPS3xGw/T6P9sKmKCGwKhRw/qYJ5b4k/oWDnwUkMb
xgUMqcBTBlHwkWAjS6NAoMEtAVfvD0OyeG0TH6Ya+Dw1wX6h7zl37UBKc0Pu
yLm7ue8j7/wM990OdyITZcEKTsYJy1doIr0ZpNZaCG8/B/91Llvt+WTIDK6C
iWPsja1koTvEZUR/FZhJ6DFqw8fhsEhsUs4LmWCFp9Oi1eIJDWfQjTXPXp5P
OpWHQ4343Vq3ci8+Q4kcn8BeP7sdxFzA8D8Cj4XXbthL4dHPFsx2/X+EeFtU
x0t4Wc3xUUOMInS3UVg80bjkyPccq5deUK6frRfB2Ls1EfSatpWOAYHzqw9o
Q00thaSTIui96B7eFR0eUMqZeE97D5mi1QUPHWJGbvHu/8mMttsoZDZ3sdae
tt8gGLAnv0sRtAXVRIzwXrzYJSEZviXXVD8tMtfbaG7GmzXXv1grg1r6l0VO
6pwWx+RQXFuHAdAuoo+ENM9JzNAuFIJzvDiUAYp8u+xdTJqPsE8OadLbmVvh
laHDP4D2l6L2nbQRgJO02jyNY6yO87/jpE37vucvFKimsZ5LK+bdd0jMkRLV
7H08wg2txEtepXTklSySGx0TJHvhJF6vkO3WSVXd1tNnDHVG1pjOfmxnHuhF
YwKZWeBfwN59SmhMdbY8jzIUuDceb1KvHWnFJGkZoXITF+iTbaA6raeP6F69
yksHHy0TKvJxiDJZqGH4qHy4cynYl5nZpcPuI+quWCUwShTwaQKTKfjwjCCR
/ekyaIH8U0S01yICllGDuWg2wq3Fgu4MnOJb2YXJvbyhQokgB4D8VFTh9JT6
C/UR+hOOpe44YNwNEAqDbT5/k3j5N8M9dvrj33E6gMCoC2pUg5xT0hlT7vQd
sVIqYOFo5hytYDKDkWYeiYMALJK7ATYvhKwpDakaeTj25paWzDjWfIdCBugV
roKHg5naDsA8f+NflQwD4wNz2rHSnIoqWAf5fNg0wYCOUx8NeAKYGIh5lRj9
/KXuQ7MLkt5V0lrzWWudaRXxEhrLjC4NrDVRWAGLZ7R/cUNyy/hKlN1GVGnA
Mn5MrTIB9V/MmLNJ/nKorNlCwrvsBpdc1IUb1VQzALI5t2IQpKYxu5bP6+ox
lk/ZoOcI/rZITcYd6qbsWWwugH337yJ5IWdHDujK2Z7emgqlSoNQRdZhDPuJ
38Jfta+UuG3/5dHxXVsO/J+YanUfdRDhJbcyJLoDx7i8q3ZP7+H4HmY7b7wF
s0yu7uSaNUgL8oBnMw2VIrhkBoaWKvk/PgxC/8J9xl/a9xk5vPDA5GOPE4aI
sMfei8Kq5zDMngP4a4JG7QZjo4yrD8fZwWlLbRBNRyEVd9sqw9h/MAx4DCIN
r/V/XeCwG+kDus+EVqkyamCLMInYLyIV5xNbuQ7/1yohQAG4w1/NIMb39JHz
qiNTcl1F3guncNfWc994+DH45YkkwSwv6KvwX7uxZ+1qf4qbXdBs3SYF9nUL
weUes+DK/eKKsc01y4wnMyQyDUkYZDlAkFS2aL0fFTTFAlNvpw9kqZZVBbQb
99NMBhoGcYgrRxcu4nQx9ApD4hlqmsmz6MEEarkxALYtSTKvaRzQDwQ5hsle
N9lhah94PdMdKcCQS5rMqsfav/SCOw6sMUt8byhEP1rnVeqLqMb4PUK+npXO
iJeP+d7QedZPaiXan0TFu9DZd99zAL895OxdS9t9SYH0HiLncBtQSeFNLA+U
fsMBgqwCgaVAfz0rlqZ430eFCrcirk3CScb7gP+nxrsiLYJbGNDIz7EYe5Bk
xD6YKaDuU+jwVRBk2vAGzPUS0tT5i1GeMVBkSvX38y/qX2CyC/S3W2Yp9NuA
nuL4H68zeHY2SFjH08oHx87LGz1xpRxGwi5HACv7DkA94JVN2kzQgyXEayG0
ti3DaJq6H2Rpr1kT5vYzRFWQ5ePCBc1hMIdUhwva2PDtFPQAd1l92hr+0sDP
FfAs3hqu2Os0LVVLATDVE/dIf7lW26wwEl9PIzJwSFebM3J+pzoMIogQ5vAt
H1x5F4euEdKj/2cOC3UrVnmT7j1vIvWgvyde3ZWadIBLBYyDJWaxKpv6gGbt
Lmc9a2Mcosoeq3LbP/JDXv1ZFpINGTlTUCBq0L++2+Mnnp67GARNLzBW6LTA
sfmmJps8vdosEk6K0Ot33+wX0BI4YvJcSrw+q7yArpoRsb3LJrTvMPPx0p1D
oiax8Bz+gAyyVyjhHL+WVEdyWHtPBn2484uwEPpLzr9ZT28N789BhaJJ57L1
DP5V2Uffq3b7n22cv01yfSPaHpQjzAx9JaqCRwYKrcSzOcunj0YBHMMLp0G/
mURnVU8UQa14K0eVL9eg+YFn+3l2Q7DfKega4JaM74mZKxSeS5oJMnXr4Wn4
9oV03er3QkS8Pvue+KmNVGfh2YTm5TI9VYuIwVYd04FhwNICylYBpLIKiaeZ
QVn87YgxzSbQi4rBmcL4ikinCr/8EJRsXMJMixaWIboovwMWiU+XLO8WoRM2
N4H5fcq7v1eD3KqqbWhTE350utFKukxWlf9uuFt8Z0BSSRkMfGSm151POdAL
2Ma5EQHwuanfTPX9JPSbAUhoW9uLLrJwCOg8nkfer9FN3DGNKNQrdp17fKdx
7m3Kmq1Xfs3zSE9gXqg5HuqZL4tLAEqOfOfyQnp1dwi9nrqh3fKyAcR/nswv
+Wjw8LXgA9AdnpfO/gs+4Q/s+JdBKVuJY8ZejoxcxOw79Ez4oYx27HcoydFc
TFa0KgS9fNYw/f/BUWcRl5hGyplg1XzRiv/tzIOBC06HIvoJLKzQSGH80iLO
OGWB0iqigFC9jtKtG8yMUOIRR46gABK5EPW3w/22BWeWTbMQUppFi8SgJce9
ve8Ko7nUAGqJpgtCsxmh7z83Ixr9YWZEVpY3lgo26W4bjDiTsjmbOqwn5HGc
tJ5vKdRrPp39gPml/pMwYXQPhQer/O0JnB0zSldNaKjoLDc9xb7vOrqBscgf
y3scgMDbGSXl4LuQpG19kx69Hz7XDFnIuyii8BoV894KNp9Cp5yx9jzrqOM3
yvet980+9px+Yosm5WWOyiLMx3MJv1dmW6uj4WNyY5DK87ZqoAaVJGGU0IY7
q3+09JIZqi+9XwcaOorHCqIQpK7187fXtJYk+aCK4I9FUE3lMtvNHRs+/dc+
1RLruTM76qd5IYljNRaNm6JWNWBE9rpNzn9omdZ0MtGbYc2yY73ffu9tixgD
KypcrMNwy4f38LtB2PR5ph1i3Fpx9AkX93xHR8JekqLXLUKSiwPG41MX94NZ
aYIwh7dj242ZKUF/K82sE/6GjeQCnE1/lQqhBKVR3XmPYgFx4rWKkhUSToYC
5fHeepGrIvP3ztytNIcjN+C2Nj0+vwzxCcwW6JMTlGDu+6JaAbUVomU8MSAI
CqpJyzi61TdP4dVqUPMg0KGSrX2Xh86vpTl28RqmhsnVY2l9w5TNquAEgXsL
SpEnUUSlcIVvfwR0CmdjdX23SaEirejiWcuCtFYKdfjwbDbnAkaH1LSb7azK
9m5VWXb2YceMeAfToNt5n/z5kCuxKEu6CVVhxQqh4AyFTNyfX1bxTt975RH8
0T7sdhYgf5DZhjrsZmmAFTdPpRPBZQ0edN0vp8pa1GsoC/MBt7tQdDenXYgb
PjufJui1wuMMjHJGb3crfVW5Zt7ydd8Qbc+zAPexptHeMH3Lf0dveKTAtB1S
QI5r0PPYN57kAxjXK4+55FiXfG6lNND2unDMu07LOFJD650Zj1rjsF/InNoz
ZuiZDfuAlSQTFDTCHQBIGZcY7vgeaQYI4yQ/tXUFwETz/TcZf0ALXDwzm1cD
grd6wMQP8kWA6Xrd8ApYGRfS/KoVvmtFMNJL3x+jLTb/uGjvN5105N5MjTCJ
j1UmIT40dBY65bRuZ3BCQyYh1ej4bc0UBz1g+lQ528p6PU/vxNHzN23sEUGU
mf3N6RTwxhfqblscXEdTVgGq/IGDcn2lVIdkp/Wig1NJleePBHKv8TU73ILo
w7+KnPfnW13McXJn7aOHw+Npp0vr8iKPaUs74blqW5Kh6QNWs928tzu2k0QL
rVZhNh6+5gx/S4v2KD/BzcfxN/ftMOHWex/WJZYoPCDicKH3eXb/F0z+/cxM
5Im5dRNaYoMVn83qd5uUu5BOzF+x7bfU6cmTlel6vuQa+4iZcIr6T86b+M3e
qmV/SZbSrMDeuwP6ArGRo9OMk3TEXfKZaaeup4ep//IEALrVhrjoVahH6ta6
hwLglNY/lDRChAirU5QU5+TyuIzLu4yBzcveaXoNX7poj7QUFuh3ZajTwVsq
6kJ2oo4k+PFKRq3rtc0FPCAh/6V7pAMTsFq8t61vRqq432EFETfukYIAAHfi
kBpAu8nuKFfo7UORN4rBmj9ELnb8v90lzI+08/zxPYiH30NsXarVIb4MOV79
lp1B6PKd/i477QI8vW27P7c5Y8LTNtk6C5TcT05jgXneCJnihgM53gmggpl4
dHoPRGhMyFAS1pSJdimgg7mzwavGR7SBi0lQINtfXcJD8rDdd0arjqZT322/
E8dL6eHVRF69Ys6ktQIlMiI4iQoIpYm+EJOfLj0YPksYxESkswsIJok4Qsgi
bCaydi9/AuPmfoPu9DsB0xwX0TBX5Bv1JlVjTimtYSRRwcJcH5rJh9qp872L
BY9UxQK6GMq3tblatNlFvyVFs0Zm5OYsvxGSL8ZTew7Z/HEzl6LywAIGSetk
rkiD+VA0EqpTOxl1PSWdkxttxZbXli+LspukZrtmEWDgoZ+oFUpI3Qo+4uh5
g0JSadaqeuLo4nEuSSH52mxHkZRU+yS+vBtCkStioezb3BP/f1wriDBcA4es
Lyt2t0a4IKxkdm8Ytdr6gh66SdaqxqypjU+amE7+QRx0dxyoZ0rfwDT1ZbO/
PZJ4Xqq5H+thUvXikF5SEQPWWpeEnPs+5X0Hb4iVnt39oSHl8BqU4w2CA//p
JaxDQpeCPGsS5Nz1H2JBCQK4bqAivgpGEvPoMrb+zIcYsNSWK/WjLG1FX5Mq
rlXOBlU7PYe5Wj2QJXIQAiLKXlTr9iK58bttibQuzIX4zi7p5QTE3hVz14UR
SAgmY3MhtpSZBHJJk3V3Qm7OgGVjNGpqagIB/2UPV7Q/j1sLqCdE+SedSXlg
hQD/oV5GRBvCU+sd3vjeuiy9tcE/4e/IIJJ6Q2ynJnBQ5UeVrgB4IGPPWoYA
XnZsTgh8pQw9Zn4peTVc35CMz2ReP9/B+/fx5FhTiYStv0QsPqyK2wzPScJK
BezqVsYGdxvksrt1xBaPodo3ednOyhp1ayRyklp7vlPwB50NqIJU/Eu559fL
1jT7A2JBuVIOJSAvSIt4IYG11X2GfV4Cj4r6njhHldaa1AY81fQKNfwbVylK
pBEDXbw6Lvv/ekgrNT+RGrwY+NGNw0ZZUjpuSLpLJOx3XC+VvBSZBEtcVvP8
vEX4eEI39OgnEPvVet4FkEcaDlcUNf9jzF24zNqi5bvA460OkjT1gzWg95n3
g+RbzvHvEm51AWp2O5I/8gW6qik/+zwM0vDdIEqclGrM06HOYSP+p52oPIvL
WKo6hMvL+UcmmGqcPGJIwJyfxmKC18ucFWFRgLVc4xPADHENsCVCjq263rP+
rhjEcpMz9kLn9mR9bUuoU2TO+w8d63d3Onc8kBATMCsiDog5H17yPkNHLsCk
GoWDTBmMpztPkz27yYTCflcMblhs0dHZPjKh1DfecjKMt9m8feQYYwgwiCuS
mE+x+Nnheixvr4VXTrg7mViHeb2ghzZFaeiTpedatD2wcUdSBB+qRY1yj023
9koAeqD1MTpjfYVZ6H5Rk3w0ioP0w9FwCvgaS/yQzvo5KboYVx0pJWP932Br
sw3WAFTZAnlpJ2U8/X7/UoDUQZzrm32MimyRJ+weKjTsJeTWoRVCoOUTsBgm
y7ha2uVs5fA5l82v72NIKRvoXD/mCFGPiHjSCJzAqHXGCVqiSA7N+TKiHtAH
b4ArtnZ8XjU2+7hZ44j+/+9yLhOKwNNc9N+AjhxLEykqZQ1esyIdnhF7U/fh
QvMMPOxEeQKv0QzvBt5hKhK8FIbqH0heefG2uBFQpDLGwTd+h49gJWBnx5oA
uNjb6Jp491PUbr9+0hfyos80ShNB6Jy0G1xdsI8Kn5iJ0j684LXQXLI/nsPp
7GYwc1k5yZLgZu4Xq1Iy2PLs1vubUu/uhmqOYdG+9cqjc2wt5pCyPCx39Syu
AtUTCS7cNYQV4TrKDm315OZkgPgaxHujKevp9QwSp/P2UGnGFXZ1Td5nf/n2
UpC7F1YgJFW/Di66f7DUFueQNzQT+ioa3lZnGRNQkU1aDzxDcebPY/BmXpSe
E7pfQ0a7K9Wpef+BP2foW3MIFwn83MrcNeAoXwS5gJ3TwQLLotAcFKH6bCs1
X5aGU2IRXhcUwoJUKcNMLhQARB8eiLKF+HQ2D9F/vMCZxEDS2p2a6VlrPdCF
BS1ShF2aVxh7eAdrBY5B9eHU4pRiAz4XuMfnXfFnp7nlObHzfZKoVSn0c32e
Xi8MjwrztKkZatvBU0nBDEghvAee3zIbKXPpp3A6Jf/O9YK3Rmz3HzFjQMYr
y7VjY7ExwM80KiRh53L7q6Hjd0lxQ7TARIi7jukorKUnoi9Zf3T/0mEgUbWH
65+aSLlaJLJw06tQ7PCWHT9hTnLVlk/PxA0reH0VdnoN+tbvNpDkOJaPH37V
svyHQIDtQ6s4Imz/PjcA/XiZHZwhKIvRMnF4iOEF5bIgcKux5qGnVFvkKFKf
bRft0A8R9JGSYd4Wotz4q/hs7hfeyxA6oRCt0d0hC/gyGUbJ/pDz/+QO5Ee+
347Yp5pR7nTuF3tlCg41dlE/owxPXWJz5Kg7SbJlO1kWDew+3EB/k5rJ9Hnb
+D5zwIuV3NZ1jXcl98VuX6KyWn5WfvcUSvLKpJ+C0STAo9w/DOCh+nE361GG
oY5vTsjQT+IvtNH9QBWu6dNo6pMl9HefL14aE0NK4Dww+DnKltjNoaW6hsz9
xP0WaA4T423it7h5M7YiT3i8SJdMJ28KcoyWtcSe8FNHlA8wIGGxqLSvlMcs
YXUtIlXXi6W27SK5qQW70DxGietfkxw2U6L3uzXDXBNIqaxc1hUijCuqmR/L
0HMqhV4Nel3g9iPIx8rjiMwzTs/yeR3U4QQuJnn6EpPuZLhUbXZoHzVWHrNQ
T+JqeedDSwH7sV2uSI2FecKX/q2fEjsNpYmApO1mf3w6Ss01JMcV4dVZPcOq
WvzNHbPWeara1rNwiRjiAYP3l5QZwxq3XJ1EextiEhLm8b4dUqDUZTurP7NS
8mzJb7/cLAaXh+/H5ZmdDrt4lNbKTkwo6yDW7EeCHJ3MNYN/8YnWG5QSdO+3
PcxsOa579QoxgTds7jRkIDg73z93FAFQhq1q4+gqEp+8P5TQLjU0ipsQM3L/
XkW2XB8SK7jYre5Q3ARBUyDmntB14FtqltjYmMwtfhhN3bccR2+zpk0/UquV
84AT/o2CEj8DqrxGscE9N5XTO8yzl55Dnc4DDkMf8Ar6IqjzOGoxtJk9Edbk
mYrTEN7dJYr/OmJWqRJy4Fx+MWbc31BSfqBGTv8QM4ahs638bM8uReF4veyl
7KGy91JIMRhSn4ETwYoizrllkoOsosIdwnXE0hgQMHnbCE3FNdxr9MYWIYlc
BEh9OyWWdjfBza3Gb3D4GEafSf2XEwei05ZJTyj7YGz5xewvfZw2KBVmtVgv
EdSzBhwkQLDl7AVmQeHIbhHNQZJrpLj5G2okvQii/eYDSiz6GXAVCi5+upoa
4HWHF9jNI5qIybTR/JqkUGwOFbpQ9timeSvXXGCqUr3tVYHVJXE8zk+xTctL
PNFwb0tl4EmAn5PMoIhZQo/sRgJoRZuo5RmDItgAdbJtKzzMSqLXggVMk+id
nXi+/k9SGuZyvwh5CZr1gRo5NbgQqDyWXk/GlVeGClJHtwyKlZNgIfQqo1/Y
67FVpUEApCBOzMUhdrdG6gb9LDy19UDqAtmWraVzaIR2EBFVhQr1I9yPCyXM
SqWUXWrLpWRSTu79dt5w1MXD7pvgvSCaYlgwlqRSyj22A90oS+7F2dqrCN5u
JJx3XjGZWPEQs4lAjUX9wS2G4z86dq+ndDITzBRv+iJN1d0lwPGaHZq5jNLF
Ei+E4WEMibkTqLTmSivgE/NOfFpJ9PmtAk3uG4NIBcQbzgZ8B4TIX+SErGxn
65/jEWE/ssXqe5CePccQHgpbxUZ1jdOTdO5QffefMBCBWkgtzABcUgcL2ONj
OrP0Ld4jB17cjXXa7TsoHdpi28BI7K25eGieO9kHgIbng4YNmNrXURw+NiVF
bi11VTy9Qdux6mIdIXOoNpmeVxi5rFR3EF3agrzqhC+UQs4yJLD/pooCiEwn
MSyfZYjilv6w7Oc+2bT2uhYQ2PX6FmqC6W70xkCKe3scnUjMn4LwENCHGech
H5QWulgwtkyYDTA4KdjwlL1iDZUXdbp9m1LK86waTf5NXmM+J4FzZtKKAnFj
uIK4ugbOUKGKe78FR56q3rkLZOkn/YEplZ8TbIvDOUWDLLxNqxX1JeWHGBY5
Vii3S7kj0SnC9cLC5iuDPxWAqUDNmCgb7+bnl9hdb+oGO1kpypmrg78HZv5t
hZgB/yyBVf2yoPHemzir1T7pHkkvWPdklYVMZEa664+Zo+33AiIaMvdzrEiL
/CVPilYQMw0Ztj16qAlj34kOc81vz2V7DlqTG1zMogXJfPREua80qqHKq4KZ
2U4bvkd97EyngAJ4C7OqzdA8YuvTWHX6N8oJ0e18TAOzVIUxp0lrkzJV/YC1
eXoqX1HzpdZXH8cjojQfaDigLwonafsu8+LdYoW/ZatsUABGpFKOxpy+B4/H
pBQ0sZzSw4ebQhDxfgUy81BFwVpEF8ODhYKLkSCYncsIDO7OeWPsKVVnJGsG
Wv2LdetKO5aNV5E62hoKmLPZEIi+mVvjNbqNOerVgXJzLuX1iXmn1Q+uEQYM
iFSgn5WQEhg9G5xyAt3U8ILzldx5wGNygG4VS6YLGPT4xtUvu73h5ewKyfvx
r6I9l6Q6JgxAx9nECMwCQTlciFqX75TcdbgQc6yR3crbC8E6nrXD11ahXwvC
HRlRqTUlfAEBYdtKlUNzRormWMk3MI7Zhm04ijyZeT1eFO2PpzisY0uW12bT
sw9G3dGQ7zfex6/5SaRHkhdzrUtK7Vnq75/8Fb3RrtwRH2OpXubqFCdE65DX
bHTnf5s4gQmo6brE0BP7/TbyllH2CIicHb2OBYgQNcGa3T/uvybyYK7Ila4m
UxPtabp3fgzgeuuiyvuIPSJ0mBgTpKN15PbchG447Nk/PB3I10QHIDj0V7Vw
l6v9/nGyTfiyBYvS0WfvGMz4vjpZn+UJuEgfggosnf+ishBhaCNp1XOytrsz
gDcerQATdKFJER+6l8+PSF+FZ1a6n0/0CIH88EwPnwpovtqYwoTCM9LN13qU
/j+/Ys3JI7wtVhTTVVh3OZN8hkbZRHSxCDGLb3gJnD1Ul2B7eaHBi6gXNpMB
AYQUh5Lr26jTzrR9JW4sYeDvGtzuvhMr6kIF5vgOB3tu+5JRLiVheFGTagRk
kM63MYhF1zEN89piI/OWEBnM/dmmXgqtwKS9VuvdFxBXRr95owVrQnezxfSP
JZo2UA/Q8CXP4pHbFGSX0C4/rx8Lrf6F/tUhKSmjIZFvCwKkwEmjssbCfPHn
qqeY1wgWsMKiGdOSW3pLLKvS/4HKbyEyTZusM4T/S1pcjTpJ14lP5iscVr49
eo3YaI6HLRLLEB3L9Q1RQmyzTwBWQeiJ3DXT6VLfuv6X1IMvWtpoiYGF3eRD
Ap4cE6xtbZ3gJ5jHemFZiY0i6LiJCERRw9VySpS9wCF+MIFyvlaVsbx3sgUH
va1YMbXGBOZbxwrHns2VJUTO7mCbuBwcB7AZsfvC/K270lxr7Ez4ZU7HyNA/
PWWPxA1KKbFlDHFsx/3kdz+uIOLFqv3nOUoatd+zfwYSJUndWaH5kRDojE82
5Cx0ZnTWCBVijsMrpRKaS9zMD2R0vZ3nM9rE77P31qW8BV3nagXl25MRiuGi
ABHhvL8XuDV+awcgUbYEZQOxazwtcz+wDO/SY+Z44h0tAauGFV6hdBBUigR4
YtARmylS9HxsVhFl8sWdK2+XO4NrWh8LWs3cGAfnzI7rINAWaf2mTRE6DgKb
7ZX1vOuRiQVXWAxvmozMiNcdUcR3BChZwhTVPvmrQ34IHL8bdciuzHNyMj6T
YxYpoDpjU7TRbJzNCPDRwDy9UPTYzQzrbulY5/5haW+XrYfC2Rke21vXYiq+
vLSmusVyNI8mTpEeXoBJRs36U2j7dhK9pZApgIIBHLRseFB8A4qZ0DT2DH0f
AxcHOx7tI2/RXozo5ZUtjfUEEpR7mWUJGTRqLz5ZluLvv4IqmXVyBWLkGf7T
LuZ9w5IEDAi3Q+eefi2rBTgLs9gsFd7WIs959M0xfxioNlTkKwn4tmlx3PAK
WX+DnavzdGZXXoltBWjnERsBe62eyExz4yuCgMgj7iArwoe/ZRrj4d3L7nPc
WKuFzOB/YJB0EvldVcTXkJxeeKglziB7oiHBvAjJsl5076sRWO6yqlmE3mvO
sEF2X5YxFk/XA+9b+o99HO/sy/R6tAyFqkOMflUn+4onJtBzxybciajFbr+Y
bztx92eYk0tlzOuEeHitQjKbel1ZdxL4yCiJJHDD+pGBmF96AmLgbsNHGId6
kFb6jVgCB6YcGsH575VxVmNNVz+jYGZb/TelUD/Nn8IL1pkWKWxsyi7GZwvG
0XVozQevvdspfTtfh0Cr+OuEvwvqk2ibgKVqrynxQb9SKYuyYdUJWUThvv2C
1HQWq29vf4Fsqs2gAahguDQUbQ7SaB1ajQgDX5NDWtRagCOacsgXJro/bfoB
uLqCrZGnrVcnUe8ejBxi7+enx0q8GiuyNzKSVMRFXClq0QBGbZ++Bx/7rJV4
jcLheIWSsXI2TxQkcimatb3x0Cm4peqcLykP/hzlk9Oh46bqTjY7CsnAhln0
7U+yVRB9IEp4GkXpz/vEuyclmUr6JSsMBGkQoOdLqj1vL4RADIqet0Ei1n05
upoTEKtiJ+lnV9t3A42KJt2nGarRgkvhGlw3aoIn0jFsc9tb1q2l9IPPUNof
D9NJhcbnJkOOcbpiAbobUlOk91jQlA6Mst7HV87WARtXFfP31QXb6m1iSevQ
IufvDc5fPkLm4E93fDFwrJfxCuQnSICszlD6RNXYlWvjJcnHzrZG0Ogh687G
Lf1B+xZoPHXQKaqQYMB130gj6aqANBQnpmNX8qpXzmYPyEJdpGl7ELPUqGLR
Wkx0UMGtZ0tJOLywD2phwAfDBBRIJ9N1Q20WupIAcOl97wS2kEvpnqFb4iaF
gJq0vZP4Tyjrbt01HeXbTJ/xLTNb4cQfXyp+LFfZ/RmQ0vxLHi/ZFcATOQkX
9ipjcWenoxi6rBP0FMORjC+l9L+9q+AeDYN9q/Q1i1fXNJqbkon42pCz8b3c
dFYKU9w/BcOg/z38ROYcATZt945mfEA1pkjNuTm+zhmRz5dMOSiKIosjRE6H
OB7sVuOVpLJiEdQAcstRGG3fCi/RUhHMKh3XMxRMrTMH6tYRuKZ7+aqPKcz5
drzX/3ZE2IKCgLWf93KYjL3cGohufV8+73LDpzv82VvJiJyg3o4q0decvnly
H4FtpDKDlpmBS9toji6akXbFc5vYtbr86wG7NNHfClGOBz2a4/yFXiQCumNg
HwDzK1fbikB8Fj/M1Ae4+L+j16V6alRuRTQagGPumtapuGqRQrn0ly4lGBe7
IyKMUzJPAyOaMtaKclDS39ggXoOvicVlVOnosJGI+gvD2JmJ1dSGRT68gGpV
GHhWnlrn+i/T03PGTYT0b2OYInA7cPMIE7HGB2cKtGtLfwNONoRev1Yk6sLI
s3q6FKpP4zneusoY6o3lOWmjKd3G9vjpAWULy9zyjKoENV689/zvfrK0gkQA
UQJq5jpUNh9P6i1HQlYNpjRMQ97czzhC+S8LBsQnLHucC2kFulPoMt/YYOTj
XOo6iuV/2eWkeM20u63DEoeXrjvnaTsVhglpzLsZV/YlLhD27qY/4Ty1zMb1
9+u+SNouL1pPH1O4cRlvcAdFjn4aqI84mHwSIoyBbZCx/vPavWVCDQ3a81m1
5wctFLuyEnYSzQ+1jg1WN1DeiBTmgdn8uyykw//noMcIxJHyzu4Qv2Az59h9
cqmksvVzWmm76jDy4ma6qx4cMHY6oJiPymFIS6RYkooZ37/jd2srpxs85GDt
zuyHsd6RJs/oDHcablxWEaNOBoOS9DUcsaZxK16sfhXiaVAbfBnmOSS0WxMB
KLNIoLGrBJZ4VMb2pu4gIO5RH+DWgiHjxnR0Fqmr/OXJkDibQkyLmoAf2LKj
GB0lZnPNP16+r7xUBw5G/2QTDHZFoLcAku0FbNweiWAr7Qv4V6KdZNZHYsFj
KnYQjJJSr4XhMBV86BgDFVAJD1UqB/H0ZEvcN2tTl+g/m7wUhoVuafx1hoRu
7mu0PzOCz6sCz5nYfyx8tVLHjTchCK/Gh3UXjlgenvPoFuz1WOfsPWI/IxgD
YZ31KXzorh+tq6HBCflD4W5SvUUnwfLqH88ZC46zmA7M7MtCM2FrODEGqbms
iJf7mfSThJGqQldt/EfCIWJFUtot0bOZaMXFe4yoFFrK077PyAfE9mb601Ju
FX9iBZFQaoPC6lKr2YUUO9FzIOQf0TnFEWUs1KYsmvhu3s1mKBuRj+dm4WP5
o+WGdnM9g7E/BQbrrcYmUdggkI4MaeoZNPCiYNcWDobBWc+ma80VO6yIhuPe
tJM71bGkE3ey5Vv/3z/M45ycSXEesQ52ng/4sVm6irQffaIMQUeoDtZsQcAC
Ko/9WV2ItSeXiE4WOgr7Io+UncRHhGQhpLlrYVzGLbXlLR1ba0ZfDmkVJRyR
pV+vIFjm3mkSNXn7rRlBGkLM/eWnGFqt6O9kxiaLl+GtWRZU1KHUWQMR0Zd1
XIglL0uGVTeCPtvcTidsroMSJFj58rP93JOFboaaSnW+RwW2CsZIQB7SQQfu
w+FpD0s+RWNuFEhyXNhROiAJVY3SYqvRS4lHrrjpVmQiVx3VIFBVR5pQfTwp
p4UQjDD77U8X4H4LE26LfkAp06xIHdasrstvEiGLnPspveVVwY99rWWb2TEj
TEBgu1f9+38gtHbcnh5lL36T40YjmQH6BTC+1kZgUb7HHPz439Mro1PR4UBW
tga2224Kk3AHtbLGFjcSnUwK2HMUkP1lAvFcIN64MOvzKcdONhjpYTIH8mmY
Fyz4og+H+LHHF0TokzD2PcrngNiFlKmCe4SqdUOPwAlsrHCbjgFKqyYpsk3n
OmBJn8ZcWGrPWFQkXg4xRqw/BMl4FVT6E65JVp8zxJwHs9G+bJiZqqWFCuC1
zaUHPF0LrXQsgoikWj+kowT7fokCtTKAmoqrwO2uN3EeCNiTv+SRvjSnNfs/
5Stit5fYu+i/EGrqdAfeRg+3BY6FnQCeRSZOknjdJyvRTei76xdedVkWT27P
cKnFr58DTJIb/qwcgKwFKLv0WkcKYixs+AuLIt85kEbdQF/lyFRWutlBFsgC
Z1prrlf8I567U/oz4UIGD1/7N9/BFP8jDmVFSR9zy24Q2Wt5vcXi0dnqDEmn
tuDX+3LaG3X9Nltm52C/Plv4iNfS7itLS2kWajIKtpbDODNcLMU8XvfPbYU+
Gi3ZuzHcGCWM8EGo/Zng0WXKdxaLjNoIbpxflTHgbepF2/s7tp5EvY+ETIr7
AUvU2qq9Mdg1KfEYIg7CjWPedWnwVsftygKt5EOboZEy/9WiRNB+rcZr4ZAh
oKpY2sLrwZ6D+R1fUctzW21adOgkOko+3EJpV9IlYCMwTAxOiauv361FEQnz
F+Dmemz+km4r2JrYlUx9rnEF55QgkxLeRC24sa9o6VVMc6RHv5rtVdXU1vyF
aBEShEYM8qc7YHgHVPKTNP6LGlxeRaZVEketgJ2k556SbWiDYCBn1JNZ75LM
qcr1UFfB2YsxzOS30R8pbrNp4NIgHSUUSCQoppB4K9/E0IX192O5k+Nz8n1g
UNV/fx97G1LoDHLjK/oGH2Qr8kGIubE8WKHPhy/0trYmrVrCXQhoRDsH7l2W
8su0Z2+TLpkgvU7QibXKRlxBbxnj0J8J/UUIryuv6uwGWm7SE379F9h8TTI/
/6Oxd/q83rN1LHFG2C+nEbb5NEEr91TFG87MsNcAoSk5bwaUt5J35BCDMJn2
neR0TA0vWE1nl2P/hNC+TEUqy4NvK+tKBFHmBAZZxOSzfYgQYteJpBSBtkgW
Tf3hi0s9vho/g9iHSl6DoxChDPkPNMgswOeuiVXr5ZgG/SUmEXxpevSAsRWi
UWjx85Hd8664tcp8WwQbHM3Pz4ECVziDm27pw2+kDWUdV/awHG7Pb2CJzUqR
Z6sPWF5Fc6dWEI62P4bXHW1GZZxCe1GVEjjEFBD1ow7As+yuN/kAdSgyB1B+
r12UCludRFe7v+oQTOGDHtuepfH92iMZCWggi447XXCIOatcd/8B7d/Hwv3P
slq0bc14HDEpWeBKwhc0egt5PdCEaspXyHG/iGfBblcRx61qlDfHGew0GkgU
nSgklWcTt0yvwPqLA4qROBVObAHlpPuDhVOmtd+ZOlt9KzL2vuv41pZvKTlt
idiWXUdiYQVtdeN8mo/cLRj6w38zywmRbctWkN0e3huIG5gt9ENwRMOyJxJe
aCVF+HtlYMd3NdSLettBjU/Y3T1YCBSBWPxi4E+P/NAYn/Ivz0ftPGfh51OL
G8aSN3JGLP9obcyv1XKp+mWeDNUjjBbqp98ZebJFs37w/P561dcV8tz4wgu4
41aexDs2fNNZTSg75NYnFwTjivSGniwh2D5+1VcNQbLjZnT/shnunW0dJ/e1
9bLoIaF4VMjlnpEE/wLqblye1ZpigVTOHhfHgUtkZ0c6LKuS8vlrmk8FMtT7
HBsVEt47mX3TL4/gjtfFTQwMQ3HaErj/aXWHB85wjZc977T0pEpczxdXktF+
fX6GWwfVnGi2+/8QppWcCa87gUzHcOI1PhP2PkZdc0uycuo8JtRQ451BzPo/
4d9zX1xCi8ysCLUEyFhBoQzes4KG9L4Dx1QvTEKYM4q/99jyxygxmNGpr6mp
8YN+IoeeoSBkfUqwtpijyuMUuHsTGzKx+t/j8kZhLje75ahPd65FZZKo1zh/
ylwCK6Xaju2SnV/FkURIoWvNy5SJZzWX3i2fUla4cn1ViPioynBEq7jovuRC
a9ikSXttmdxhlaxYUCtXgVYGM81m0tX9Ls7Nml2rj+3nkFPtimGbdOBpUhKC
FHEFyqIpYso0Qv/8/I+fJIE12DIdmkpWu3lxMDFpddlVnlCCEXF16fq+gQCz
Od4MD29pzMtrYbOFVQx4jGKliCjCIdJfrOqbTt/BAjPJlp0mamFMtdUAyebe
yHVokz8tH8ugB+xtFtMHGXgo11mny4pQilRPGkgYhNx6djJees5jDWbipW1v
VQUIg3q0iqlpBEaEbV+/Tlwf3w9ALPsDStdLX2hYlbhzy9Dhp3tYssExCAY8
7doXthyl1nQ2DDjGaRJ8nw23HFRBKzsDX+gjBaYxim94SJjmVS/P6YiNoZsG
ezjmBmed2WK8BWUtdzuM19ByMbr66TXJ+vewDlAtEZ/Ps5etddNE1ck17quM
UfsEvGTfAugJ84pPsAfTFeDlWK86awOXJiflY7BfzzTeEJf3MwMec1cPkrsT
SMXOdmLyKpFyWA0gU3rjAKA/6SiZZHJo4y9cWPeIjtps7qW6Qh1gpuYvyYDf
pP1z31l6x58X130OjEVb6UP7gYPJwlFfpFhzwnL5gEmpxNSxljVPsQkaVMEl
x2EwlslP66/RyKnA/i/kI8MksViSo1voFYgWG4xlFmDOv5Hwvora5Ue7n9XH
aNwv0XEs4edUa7YGFXAGAfLZQ6//lqV54ywjvtDmPhqkkMP53RJiaEoNODYm
xzUCbgNSiP1HDCRKnZXL7qi8HEqJPtyO7w5DPN4sYfJl3AXCsF4v0ZPGd/ra
PBNv++kVLNRJt73ApSAvyRQ95R95qUZDzlJVLJ1C4ID+QkvtDXrEQGu2wJj0
Ui97C29gYJDVPb1IF6d8udaCZWHgFYzZEYbChRKvZJeZedaiGdaOZG2q7ZOR
mloMW3goNwP+Y9R1SMZ1skxkrv0W7SNTDd7D+NZgN8DJcxVKt5cj+D5CXaw7
Z9Wimf3TaJ5iQ57Ed9g9AYi5brSEn1zJ7JOn0XRZ7VFeUVKegrv1cNvRPzIJ
iEbsoe42PuVJZOUJ0gBe3OYfy5a2DhY841R/nCVqqR2gLiMF432pHu14/BG4
4ESPDLKld68jv+41O4mKu9Vw5X19FZNktDwLuZ9B9QLAS8yBl1Z85cC5vEWV
O8hfTZSm6yKiYMbqcc9JArn01sM0d3Jo2D+t2sVdJXeE+AVpBMQf1W3EM0DR
PdxTLCbuiAttzXBuyOFdQFXoItpve4z4lPgLDfvROuX+5G3zX/v7iZp28Q3W
HEAD771nUrgq4PQP/ZbCP/6iOZKYmArE4Jzph4rIuqAOQiIyUOBLA6ETVj3W
CEH/lvb1/+tuXr38jCTmSI0zbZA+ALuSaMKFpsaEXhM33SUCGD/iybmVMnq1
xSGkl6PfV8m7ylCLYylYJngF5y2sa5uhi4zFGOdEjDoRk/3R+reDIXip7rpR
tuBQ379gjx/QarbSpfIu4u6gWlpMpAM2sBwmyeYuyzneN/qaoqcuX3V1tLH+
9FeYG7VjdlTs3llaUdvmMULKA05M+MvG3e7AqNF1jLxi+31oGqkjPeaPHKCq
Uc3HEcd4WlfCKqP5d35DAnGKzD8dgk0eoy+mj0KnRrKvl0qJdjd6AOrWbGMW
xEEw2nLzmJX/QMPrmC7obhiVmwJyqsvXIKE69i9Wl22Fla4amBgsO2AkufLe
kA4Rrjpj1K3u2/YAa9g0Kr0bDjLvSbVMwNgrHl+tFm5roTiT6C2+VcgyaYe3
bzSgdTa5vsF4Tle1Ff5jrE+VaDVp6YhgFA67MoKj+63FkcxooY9PSZv1joUe
nOVk1/z6YQP8PfK9/gZoyfmQTI1OXHFYnV/XGJOhc1GKZ+eDEg/9Mw9EWGDY
3EK4NU/Is3S/sGPgIuPF3TVYOwDUDg5mpsebojg0coKofqUZeCMcFMBitceY
uSDIe7LlO6/UKFYv3rRSWSx85SmvFJl3S+fKBTeDUD1tP4Q3jeqk2v0tOdUB
qq6LwO0XRBeK29hK0E6PIWHwRDVZQXohof1la77UeVPmnhJ/DdOkkieqyIjg
qS974aR7irES1jJOgMSIr6B/ozPjt0bFZJlZfg/Oivy2+cppA/rs+Denf07v
eslHgLlnHJPEQDxMkg7y/D3E5bOMCf2VP/jLFICZWIU5wt+BGhzLWLNy0Swh
5YkilzwXQoP5844WvuUY8c28+pHszQ2bvCaxTeOecUXuBVLg4T8TykozK4mf
h8udfThrhl9dCsmDf+CziQa4ACI/Sad4XHYm9RlUfMoBm6MR80NaUkBgOJ5Q
gEvf0lzO1JDrQseuKyko1y7buORfWVx+hZNTsYPJEOZhMCa3ryOB0kkO/doY
QdhKXb3min1Hoo93DnesY2LPpcPZv8O1H8nCUXp7mVQr1V9pT0IfCo+aREGd
6CyVWsQCK4vKRbYTqjO5XT51gu7QUQ/QL1jYesWS5DV1YYeF7A34ws73NgaQ
LKAfA4yLepTuWS/OQkHCEUozCGPsEVXb0VHw9YpsMnwj0MWQ+yvysZMMP+rt
WJ4fCFkLPeAzTK4YqRGSsBsLH4nzxlKtelGrLSGR2JvpK54n8CpPOVGReFz9
G+nTpyjE2anT0lxfybQFjIby0+uILQrQvg0io2jQMxjtTGG2+8xyNWG3llmx
LJHlLyatV8WhQiFDeqzZFDXbKsZLpmXyCuY8CIjRPXIqqKdsg5C3xhvJWPw+
mYMgpmWz7u/TaYFNR+XOtNLScerMJ9u2V8kgkcuQWPF8pazQwzSvk6AOD6DE
Nyfj4t6+Zb6W34zaO4NWtJ6h7hAtovI1tok+heKKlQI3wDD2DX6IXz47ee0u
a7XJducIDTLNGEqDTsh0WUbF2NgJRhmRgfECZhsqewO6h9X1ykjKWdA6ECYk
UImBZa1HixgpmZQpDT3C+eTNQNbbAQl09Nu4vZ7RAq5vtxXueLf0UMdW1/JZ
xtdS64ohfTePhyd5u7D97sIt3txrpqA/gmBLuuSmr4gdHlnsZf2DH6ydQWOE
6v7tqCynG7HWeW2boPuu44gns/qEL64KVdG9RspG6s+hlogHtE+PzMtZUI5c
Mz3n/1BDe3ixd9a41B/zHZtcxEueEswCWbyXtddJWpPNbb/PiOcSfF2TVzpt
ChJtKByt1KsCSREiZK04PKc2xscTI0SteQcKOGaANeDZeJgg56ySxB+xuHn6
pcv58ohlHOCrFjUB2JtqqFyAeU2koS92kyIUIM2KKxUa7Vjkljtqc6SLnOG2
I5WFZfBBFtDyNk5vlhZQHQ7a1J4Rt0TBUkOmZ7b1bQuoGPEl4Bv5g07c0IAU
H9QW75762OSMyRcStppeua1O51M3FCl3yT1LPoiuSZAVRz2+NKy4aczWHnyS
zPZBRM4u77K73gTcWyb5PFXtChG8SAgeUiNhwj/81QPgoZ3z8EsXioX+LOe6
xnsWLKl0zlEJRK/tDWeiUqMc5jxToCw01ErSLcOACCMQh/vBD4ORq1/L+jg5
OLostr6y1wXtzOJ3kgYHeQF2GEthlPx5DxpAjnnuExYgaKMDnHvoC1QDUKV4
/BzfOiRN0NM6eiEmlY+4FQbcax0zyPC9hmcCd87um+8bKSzDYtxks5PLxFCK
AUqJutFaEItD3yMdSU3Zy3HFhg4hnbTbxBSur5X7kFYL6UePZ9YUjotcEwPN
APovmeHohRn0JFgoagCSI7l9goCMSBnvMcwpaSKht5/iBcNlBFUSKCTdXC1x
0KT0+UCk3KXBppTvD7VjSFZ80YDeITYAZLUK01kHfRLzFwQtYK3il0rGc+ov
m1dkBNUWLN+NK4j3tbmgAe6kPPH7sKljuP73e8zuk3OjTxjbI6GQfboP3qAY
gVTpAFuOag/6+WYsA+Y1G4utZMsAzw7uDqwkJZSbor8JLUsd652GxkWjBtJz
qFAJKZqGrLA3u0gKrKxJhKroM8uqHBxFD4rzd+IK43i8seVTuBG+IYeEaazj
OcpbRqqVXV+5b3RMBq11JcMbOosD9v84cx5kVxUnZZidKIKmCldJzAeVCM3L
mJExGwrddvagicXI/qsIcP+M8PUuiOT7mlC+vyrdSU7e3KwTtgQ57VRNholp
t3ujvz+2/2QaP4yV872KVTr8cJhH8D7y4Q+j4/Pj5gU9nliGAZSbMN9rUSu4
7r8dJD8Zb67xjmpec+lFczDd/mSMIZqOL0WrXLTaNsyHVJ3Q3fY69NKm9JlG
da9gi4e8+WGMpkvcCz93Pb0sUQIltnQBjpla3r70DUGU+EYaVryoyXtVz53Q
Amr0WKythh4N+HT9UsM00Jr0Er1H0ngITNqWMOQwRqCzf0wj+TJ1Y9m2yD5u
Kj6yXlb4h23KLbr7aEOuH+VGXWv8V7encX1nurZf/4/NIxfcTWmZGNCxwvX/
qCyL68Nbgfq79DT/ijiW4E0vHPiFiD7Ixg1VMk9coiEbgVVl6V0+Ei4z7xwU
z6b8/TWwrUiasXkphwUfOralnKfnjoSfsohougfnwqfqL8FeO2xSAN0BbY/c
bNERYo8YJ2r4Y5dHEBLiL9+zLlTGwnwNb4yNv+BbRXp9NIugZHH9SVozArRa
v8WMPcPjLSjZmjXjUCGt+/1QfAqe1oNZ0ZnWKieSUcFHGGhZ37dyZfNWyk3q
4dvf0isy7uNbdtN1HO3wXxisGRuV86n/udP583KNNr8KHc910RdD9rAv3rIG
CTNdRn4/qRSyt6hqx4KBXLL8TNo62KXJbEux0y23cqAI7aBSCtD3XweE25hV
VbPpS0RlDhr2r2OQViXr8zOnCZZWdP7OT5/QAEJxII/bkWYrjtl+53D0IoqE
78B3h1LEOFjbT9VhfeacB5cLgP68K3eDdzZFE8CzbfLwvHY7qbPnUS3cCVoo
qNwj3HX19KB3awfUvNKkBdkbYFPB5hD4ktrQ6qHuPvXqcGHyNBSfnqRgm53d
SPnPXVZH3rcD+oa6N36TzyKFeeup4yFZkIk/mx9UwDJkZ3r5e1JbKX968Pcw
Oo7JXvWLFmg6cx4wkJoV5+3hfCjYxToMhxYWDTknA1nTgRQc2vKU5543jgmB
AZ5p5YNey10zsHyYy0X9k0sO6ooqvZ866dKLvHihCTEsQo0cwmbyBcUy2Syy
zKPa+iS4BPTIFLFbKAYoJkt3e1KdFmhX4thdcKXz7OtHVa9euAdmeKIlqARD
YtBAmedGCx7DRO3pBSp/jfqH2h7ALdqEYYBgm+WuNw+lvh2wp6c+UmTw2/7g
el59PKHCNN4uzAHLd7c1tSlFeKHTvkhwfjw+LARMBCqlV8M55BM1428kOIXE
yGw/3jbgMmAvRHCFCcqQngYyo7dXEpp/AmcOJZgHG37UHwscG2hOoYIDO3bk
XL2I+Hl8I1GgOTIL09ve+MiySRgeElLitWABTSac0LnYsy3R8H0COCk1HEfg
YW4zpFTQI0o9CBAcl+y/1F07yHl5pQbhaQxzoR3gX4MjtBzvpvnoPj6uHg5b
n8BdRxr6PIa4kwmT4wnmhYuExN78qItY/Lf8DKBvkqQjRupm1qBLJBr0nxRY
KTvK1eBLbWJiQYlV0Vqflz23BoAFXEQAWF+g5u6QoQU4O9sf/gFpVGhPzaj0
dsiF9Gh6NFMpbFkj+u84kiY7jQbmgmfEiiJiGFkO126P9eKBKjBl32sCla9s
DPbnWrCTC+7lxpHv3fqQshOmomC9DXquXRYW6yvu/bYpfpgIqEVnpr1ipAOg
McUVsC4koj4yQpD18G+zEF+FnYDzqTLl41iFPAW1jlWUQX/zCgP4zig+NQQA
AFhKlqyhOuf1FieC4XIw6CfT/knv++MnVSdosDHUIMyOTbm282U+TPwUb/qe
TyG3nt3KdmUZ4jOYaloorKz1WAXlUf2V57222jDOLJyIzw8awedARAz8ayaR
6oStiI7+wJ97PQFajlet8im2k6ScvBp1qo8F201buvCio5wHrvBNhCvWT2vB
iak9B3hLl74lJOJ7qNPDKIi3yaFiwYnGIxDWo89vfQv+8tp0DKvR0Woz/fqp
0OiyYrkz1Hadi0TZWo78A+q7NpyNlwqS0++5TN2UOR5DLXd1+Eu+t7gEIpUT
kX5qcSBtq6B5v8nU7SjlvMo6qOpPAZ4aZ+1mdkhQNyVqEVIyJO/NXgL+776E
/Gntv0ToBvNCwo8gJE2PzMLpA7XZwyWVUxFXkR2+2SGFubDyhLa5KCGcV6ph
8p2PVLYx3qkx6aINVqHiE7xh8nlVF4epEgqGDsvjGvDeeZSboMRc7hSclN/B
6QOU89amiHTLmrN+mfoS0oCyZC5KJeZCf23r9mDlft+1IQYDOnEJkjNjY+4W
1o3zqfgabxIgv90uTywqCKk69o5Es17NdqJmk+TRAcFUoUSWAd4/k3195tqh
7v4/CUn9B1242ub0XmXt8qteRfDT23+z1mGWWehD1l6xHiowsEGt2lwvpwHJ
cNj6UyO6bTdsTBiAG3DD6FYg36BnnNHi8mQUW8D6KlNXHcLkwxoncioDDkvJ
RjdmREjVvqsqqoljQ9QYwkCoHM0gBOis7XaFkIKFI2dtMrk8iT8SaWlADvIR
OpoKtKk4EKwm/9PrDDFEJAP+tSJ8nr/NnvqZ/0oVWF4itHisGf1LJPzQAwAF
uUX2LvgVvaNeyw6CWyMsZ9HAVlJ2o0593usialuk7B3Nf9ppN/YvcvV3VS6C
xUrxBQ7+1EMVx7a6BL1DGDbsPjXbcyHLwbSGDjKDcooKiScn46lVjC6i321O
xf6nkEUwXDt9pGk+bj9Gx8abEOeSW+5BcN1/iH5B8wgabjxnFuwL2HP6nLEE
mJC37iwDiwt3iCcgnn2SKmgAVGDiqwbZydlqOh8qhbhToi4Povkvfz0fi1/E
njKq72k98Ds6agbYF9sqP4dKYx3T8UyguQZ9mrbQ72GS7g6uBPsfm4vnxgX0
hvrD8SeW28zkPlzSfwrKgj7/cDiefpej5wwSM6dOGWXqvLw9euNoivZjeO09
X18ySwbmzNrdPgpCuwwmgG8TM4V9yx8Nzuxyf3ctxdrAsME51NCm7rvg14MH
vydl19b5D2c5Ee3oqoMSgcJmTep+zlUnG2kxrM4WWYgAqmGOkbrTYtUgByPe
l61alrplUy4m/j+tZTw6tJf9phk3/yWmDdaIgCMXgC+UCk0QGo9ZxsuXyR+K
6V00MfHGBIoOrVEDjxGLKlftjfx17nmZi4mXTZy+22ObpMTKgsRqskxB1u3V
C7FbSUrQhDntPJW7eMlmz/Z8VIn1csMI//NQYAS4zgMcrAMJVV8eAGZFwvUe
/JbPDX/sMmP54nYWs4BGooYPR6abJVHDx20KBn+05ztNUnb54l42vrgecyjh
OhJnNXrvWKfH/4pQoYykJLy4670OYsjJaKYqbpP6/A3nyFi7llgLsFkaVQO+
K2J2q6u0Gb340olXugx5ItvbeqmymF3zhlif1FXrnuVLLh3BblpP4tK4F1v6
Vo+ifmFd95EwiNB2xGWhjcotupj6D7MDObQ1mfFfNpj0LmxgPuVRXEhgPs7t
jZxbIdbwFqDvCTI0Ev43L8Zx28hw0uXAdkjRi652Zy9/KCxU9zNPQo1+NbcR
8lhTIA7UkRy/zdfvqytVj8SISQkTYd+/N73pNPJq4VpqNcqAG3iHwawjL+0u
YsWNrpUk+nRMABaBhX6SdRvzJMMLoe+TLLy3eCd+LYqde87Ix5o5WWCa/cmX
SrXEcMVJw2JDWsS6243ZUC5DkjvvBqhc7wawkEuo5mhGfn3UidICE7r+dbQ6
aKEp9bMPifsyA7ssI5A/Ao8N7dHwOduuqJTV5S5w8ot37QJPSIOLP+NRv5H+
BtWw2Y4tXixSnRsRZpnODBqzzFEiYE/el5ZLZTbUE3ngwCNPOKhD2lwjgLdZ
iA/nLEhyxcvUrTjWqVSkl9scrteniVeALtckLhS0b6GWBCzkv5ifV41j4zip
ffRz2QpL/6esR+h7aJkyXfjzRkdCc9ccUzabV8bwnIQ6pPPsRsDirKUbxXw7
V/xAOwwkJDnirdHveY2aoy/I9gZM5KUhtFi8xXS7EmLB67sZdaiDl7iIphEQ
/TvVQJvb3t/ZBA4JLDGDSXicjaIM+glc8pPCM3wiAZS/lShBCFlWr/XWbvyn
eHk128Kf38B0P8ABcLnF8sqPcLGBOS4VjN52qRFONEqoTR58PsqE+07+O61l
03CcI8MiiPCF8iCb3/1uSGKW+M77uvg2y9m3FMrlmCqzinKFBlK9KAJmGs2q
eFYobOBi0sUK6nOVdvybnPnoWuD0sGptQZv9V1foV96Q8+xJ/QtwweIJlkrd
w2KjIzcmrbDFZ/CE+I1+3SsyAsqJtVYCygB9Hx7UhwxUv04Zku2zSO49qMsc
N8+sCX/KSAJaKXZ+tddCnqpAUS8y+4Xp+rO/Fqi/sjA/kK6xETf7MQYG2gko
ME4dPvppwaFoXoZMR1Qqxi4xxS0h0ubaryV0YIiamc8ZB4kUfnczEnnJPVzC
yRpqBEb4J65Ut+LMjdXgR5r3EuWKAqlhppA6ymr8T241p87MBdHPxwhsCl3s
gocNC0g1JVdQhgki2DCcDD5+Xuz6aW5mwHLtJqoGXJZj4fk5j/WMtlQud+ba
5CzUDOJ16soRbiChFV2vuvrSwnel6ywYBfsXq+HPkOHDUyFa0ae7WPnKa3L6
cYCEAlUDldQMa4ky51Tc2e/Akf3nvluK12cdyCv40M9cymuLwMwVj3USmFfd
lTJ4obyN18RrvpOukpnhVPrE05KcayW0cvfi0JAb2Ea1LEY2tiE/Uucw0zqP
aHoGNUYWqF0cQMhhSBhf1Jp0abov+ea/eZg6uewdE6EC2SK2QeRzxLYDkFMn
X0MIlw4lWuVtclzYfvs0B1k5SUsp2SwHXEQn8qVTCTNr5UQNwi8qabL9TNDq
5T5ABcbR8sPkGr7uLMv41NHfTVSwnQQEdZfnfR8EcQdvfBQuV7l8mWwfEUeb
ruyxSPVqzZlDh8AvbxrBPMh/++SwD0CvUoE8+EVY2Fn3Ov0f6SMD0AyV1nM7
H+j1ZY1pkkXZXRYhBBjpI73o4/yrwgF23eqJkKTQoKbsBepHXKjRYUkz3wRs
/cUm4hh5Ijgh3zxS3ba5BBqFC9nW5gPfFZphVvPkkLkSWzrInfwTPOjgnNWG
LGXfvipYQaf0WSW32D2C75eKEyuleueKTY83Il5UvGaZHntvqzOFoU8xGJx+
e/1becEZ3/lBuZvdD68lvKehTXAav/3o16k6QSyg90XwA6AjiEFCWGwSfwzT
N6XNYaxpkQjXQmFeNCIPtcP4YG2r9SxAsMvFkIrigBxQodobM23OHCLYRx/w
Yf5UeImzFrFrWY8XhKntHNGYbsgoRTlqieyN0VjTLCZFpjyv6pPgVhLn4/jt
1afsw9a8Efvl3hyoSe+wC16s/npWV0tWqvRMyEoZ5ka0v/upkuhMHzJR63Ur
b0hyV2s9wjnfi6zPro5+v+kkwH/qdMhaoBoxd4DPUC3x6+VA4svoMScUIN8s
IXuYdwUTNyjxMH0YPqCnAOhMLjGkNyiVqDEfBPCUTbmctHbkA3+YJUNBK58I
icDaRRemht5nH6YDI9MYS8IWko5S3XhxaBQYujkS1Wo0mcqgzAu+UWzDRp+3
wOESEkq1WMY9TgE7uiJiq0DqKSMsD0rIQVKYuP0HuacWIhW7A6H5LtrDXA0n
ol9tGA+lrv6nhRk8bdkJgX2zkn4wy2AriDlvq2vVXDwaUmVCMfNcIYJ3UJro
URTjQmjHSTefNs4544Kga1zZRq6YySXtqvs8fCprkUeSXtZgEnMyeeb95ONx
VJ7NaZuoWXssZLt8HkecLtetPZlVf4MFVDZm1MKi7xKwl2DYCoNg+Yqy7qQA
CpESNgsV2XheHhwdjp0q37HvIQgLiSQsfAslFGDUiaS23KFLozczCl/JVPj/
ayJhCXuKM0c/akOguqehmHesUSK+KzUfPSQ7N6BnBWZH+x6GmyPWQvl3W6D6
oN6/EBq+u9hj+043N3eMkarjjENZXlhhqz8gB/uLcFIj8OrR94KiLGg6g4YC
5j4pFt1Z/fwCjRQfuRE1X2kvmFXZy4yglWWov932sXhbCDornbbMhKcu0DXO
BRcWdEBlK28iJdmBKCYJVj6j9tXvB/EjdRKCc/AxrfBrqIR6xQ695W3/uZJl
1EDEEqbPrzfYmI9k1lcUCjybdfm9Z14TQSKKiDVyORhBpRd7xYYitls5aiGH
4VPO+NSw2/Qs8XO53pxjN919Gnpns1HG9mMItmAjRqygmiIHYKc5anX7QOkc
HUQvnjhamqYLkPFATRNOJDjuk6Ia6OLKlhyoEcUVyPw1p2nbOzD/pu4KSCdv
couv2z6rCcgN+uWf0oyW8cG21kfKCOOPPff0XMBWPnC2OsFPnCoEkOSEBJYD
Nlfu9Y56u4rEOkn1xb+4kB3HfiYGT1PxU19RSdmzxHpEfxeHf5UDbY+riuq+
Mhgz97IRqZ3eUdCY+SZp2yk6bsBnGC4gyi9RO/RoK/IpgVEf0Xls2jU+ktTx
xDxGv5x9PSZPjxn/NNMlKG/y+00+OLP7YA+2ZzFjF3Dms73sGmwlfV72Mo1I
O7aHK2n9kZkHhIvHVyqpHQiqts8MZYIdL9n5qpIk98rQuxlTyGgYXf4T1Olb
0RcHN2Cw1cqEj1G9aaW/b7eoHnq+lfdFo3pijNfVaMALxv4Y2e1y6V8A54Au
kcbPaKfIspYTZAG/m78tjHZHIuO48SU5mkEwtKZP+WGEYTFNTy475Zx2fGxo
atqiO/8rx8fvSCeHUco0k1g6Uk1Rw2sDFpetUwRfa8oXu9pclYiiKGKObf92
b1+gDYwxaiGNoCHsqR8ZYOcLkl3mgcsW2JC6HnrRlQOgMcf6zLy3BSie7a8k
Q9TIRybhX3pWub6uxFFk/66Jf5qG2rom+7aIG8kiiLA8grgRsyGblrrCeFuV
tqVanwY1mRQUCI8oGBPuPqtzlX03bZFvhirovL0jRefxGmqKqFLOWBsU2fcy
BzSxKYTYAm+4PYbIyzXbI5QCRIiYvJHpZiwjuGgZDNw0iiSLmIoV4qEMdzg8
DA/0kMU+4D0FWdfYPsEr/PyQ2j9TCel3Di072n6UcfCuLyb3QPT8VWpWp1R5
ZPcdhzREw3KQrsGe119jmqO+sOtZvXUi2K4Gu0o3D4QNpnTMAFBSlhHUiFxW
hYfcOVFGhyE8tetzcb5Se7XBIBOd2on5mpNMOy8+WfUuAflpGcgHeMvMzbda
62eMAKxypDGqKvTEtkeSe6QlJGo7DDKw5s9QCkFmBvj5KY+an/gbo06eGTZY
eHy+73P9FwUQDDO8ZvXV3E0CAJdqAAMBEPApf1Qltg7Cbhk9JwEBerQ+Vo8H
rVGA6GG/Z3wVUqnFBguhzvVkGzHO1a9EAxyo1ihOaYPCxzP2EJBbilkH6Piv
NBCvICAm9oeOrqscAWWGyKgjTjpVfiYua6Vs1yu0M4THfi+kV4xMaYeShWFn
lavRv0NbaAl2f6/quELtoOKZw2+1DSeClTA7Ogf9GuRx1bgBbms5es/e70ST
9BbkKjZBUwydvIYGmFPmyZBPh3TM7DIhI+nD3YHMiNDLDywXkPt5wk1eGPcR
JzdikxKSF10k4jPKBaHS02uNrgIlNhGI0HXDYrN9IqZb5CHiZFN0ryhXouGD
MIz8TWnoBq6QD3kb5EKnpkTMeXItmIOv5K7+Ug8q+sC2pHdhEM2Q6ifFcC4P
FR8kkI/cdbnyBgDrXAeFzdApXRDAy5V1KRASdDTMCJrqpjTQjHQJTEkyutyv
gDuIBBtJeDVST1Uba3AIkntmhk0y02mcgUfoSkgnZxiNFsVcjgLeyZxzCKtW
4gWGAj38GMCjohCIXr7orGoBizin+ZWuVxnnbezmgX47niSd8DVDZyw4WO6D
enLykXkin2GdE4cFTzJRRMXkT5YOIMtltLOZ67fZo3jvR3qJVc80d7NTnmUv
+sAm3CHO+HB8Y6NCSXFxIsfBH/hrzI3PCoRl9CSlal8w83BrzU2d6mCLnhKc
3PhAEsMM6GjP6/9K30jDqEumttZvGlhRfoBmWx1+GAZypW3oyk8UzRNv05HZ
gKs5UCIktDLkxo8QAOaGgqW6qbFNwcGDQaukf6KGsSRMpdEvzdqbXerFSKqM
i7a24Qkn19X3hjCGXfstn3p5KhbtzQ4N8ClFMJa3T2sNQbEmDQDMRM96tqMv
jkpWcdaBTZQVxYYzQVVXb4HFZuoNJAQOwRtX9JmD1pKBD2k+LPl3tqve2V53
LLp8jidR7tgWHdU5a4SsjjQKFO/UWge40ygMugt0NUDrgPMpmv+PfupShRn0
50BWzZ8PoiL+1a12d99tPi/FfZty4rkB1rTPvr+M01mJqvb18VwAdzLkXRgt
gE9JZx+WWAPOVDKjcmLI2HJzg59QXHCyvseYbY6KY78Vu41wiPsbxtFLywZY
rMfNrqD0FSNMr+cGjtFue47f1XggsccJiT+U3gUI4Nf1vbkhzOh4BCK4g5d6
Gob+EXm/4js2NpP71omIaimxAIdZt8nwFUpKXEkQ/LZEdjvWRKzTGlT4bO9w
zHlqUHP5YdQ6iW2woqGfzqJ2l9Oyq44TV0fxYDgRUnlH3kjLT+6kFlQptF9s
0ZQBByDSkThhAwCe3cWCXEEqTl4QJonIBPFmlcdBYV4ZNPRG+UEvmesrwtoC
Ee0Ko+epAOUvUge3qB7C+XiNzNLJZZg8OElctZF/85tELV6CdmhitCCfRkru
11dhryGT7zZOSXaXjXzdYyrVAYRWhXWnq90hp31eRNHkW3b3fUyUwTtZ3pFw
ySW6TNbyEsCLR4hqp6bNVLH2WSSnE+r2eSt+wajheh1rB4ki0fRs9C0zXDWt
11m46KnJ8n7l6zi5USWH2DHoGOKIVeXXaCBPqfzQNJMYyv8hOliQG/OIN7Oz
P9Dc92BdRHg2knLf6KwzjGJJ+/bAWI/Fb2qR0dZIw/p2EMMqAEyYAKKbGXmJ
BguRfkOmg7k6m9H5EGQb1XpV2t5xCr1OLdWqblBtDO5h8DYAZhqq+29cYnWX
SrTKe8/3uk9TTDgTd0eWGYHD82od8abji86qQYXCAOIwD633xKMUbrPYQxRv
6WBDsAIyqULEtUrJbtJOpkFeEKzKxky8rVSKKrot5NIpHTqqRddBnV2iU4Fo
SBV3ctDoAyzgaOt9psH9S4ac8jvuj53UaMqeHkHUAS9FjiatSRHDPviUubfD
0mf9W+swBeNT0Y5EkG2bIk/opr5HFOAl3OgwJQ6HfTwtTKzo4fW95t/F77PU
rgUU1ce0ATG5EmCCw3guzLzmuDUXzKlVy96zIhItciaVf/rCno7r8ZthoUqV
fkkUxcktCl73R7GzIgQwE3WkqYoo/TgEtFuTlUQTJcvbYigppCVY/pCpfqJB
5wkPAVqSH5xg3STeSdPoMF0I8myHt5RZIzkIl5oUlf2D4XUFv2rLsIO1QlUK
cVacX6nFXuiLZBKq3S68pT+/MVv8bMeUefPhzdO6Qe5Mi/HtK0gmZRPtuyTD
yEzQHcS3Ef/mYDVzfQQhWmaFGAfA+mLhZeIfZopIE9JL7TSZ1BxBsCzEd1XB
WBfpz2qSs3ieyX8LKzEjW4X2m1NqmPkWiH4iljnY+DEiD8m8m+9sfHD6HCUS
80zT5MtBXcmSVZUkrqJGbclm+8hRlbrj/Sr1gbn9oLPVbZ+0Oo986y0+drkx
tA5qdxlTH+TIKpUv/YqDo5mGuxlEeUanx+AexdzJda8jX/yjTI5goSdU+53t
8LT9xWmZ76R274ZpbObBtYE17stqLhUQTfNPC8ZglTxMaMkG4dsSg+wlpiIE
5ZUr0xD8CxGRTcuWC2mYubZhkYMvyo6Lnrq61KrrqR4W3ioT9ciFa0Vh9sK1
+ncPjMxHro8QvAx9QTHi+pQBYqVMpiA48YlIevSVZw0fEjuSme9Dt9hFonyy
09ot8I6OxVW7iDQ6QXrAEuWgAzWke/j0f0znCH7C64dGMRXC+iIHQIMQAVrg
BNxw/Idt8oMo4FLNtB4be0yNpUZY5gM3VGhQR24gwVlCjsvWZWEETkrHcT6u
dypbLVXplpErH8GbWrMRKYk5pyppepg6PJLRM9KkadSzzkKbOcdAlIwXLWlM
ltlXSSIwJjy29pBK+oMWlcWRzjgtD9CfxPAdB+zSmP8nu6NPjcUnVXg0ByC0
+9JxJSTXzQ0gRodYy5v+JJszVPypgYH2FAOIFEGCFRK7hgBpIp2x/CBBKCJN
q7zhudMIzBdckfo4ooYGzMFWJCsFQCKv764nULDRBII+mwKYSbJ2txGpYj/I
rUxQSG09adimTBmSck+kSIwcQm6OtRc9W2cOY9bDPUf0Z585Y84hVznJ4+Px
5+Clj5NEFdPNSptReUliqpuIELAogTMvnWb9OYOtvUC5ArxOMZXt/kNcEfpE
AYnhuUeP55vE65b4rFcg4n1V1Vrr/o5VspBa9LV/4zz4dyNLj6ODsJOJvaZ3
kJB4m4X3exCrM5BUcvur7G/cvsb2wBsZhLAfuFFnN6rnkL9zqbkzK2aWYxNd
sgbv59yw86uitwXTmZlgy21fwhwTkQ7Mfefq6QlEhL4lDg9pIQ7uBFs3Eswa
WBVFTASLHF8vmUD8jd/Up6IOzDqUUlTT5f6oRIFqU8xAYmRIgru7lEPl9nCL
CjmUjYPGZKbBDyB5c/XOdsF3SF9L05NrR/s933m4pKtZAtbCIXBtkq7+OLkq
ocNJg1HaOIOYKR9eVGZB4UCtW88I5Kp/WLsg1IburhXZPVnIkpY22Vyv7D5Y
ekFTsotLkEkBTMc93t7gpUcG8X3ZE9FoVXa2dGOMzM+bNP82U8VSJJngstDY
TqMal8CyOU3/k0EwVnNZcp3DWZpCVB2zud98GZWQQQhXFlATGsjZnsvnysHs
eOsblDNlS6u292H52RnAIOyHgjbhEegIJWXz53vQwDKqR+ayB4Iid01K4psG
HD1ljz1s+WkjiWU8KEhTy7D3J4X3aXxV3/SnFnleRJghdt1Yatsx5OKoj1YI
vxWXC3gKktiTxRkhlMBpczvb6ZSi6mj62DwwwDgBgD/Eevknl+qhk6vj5LaO
JugycfNsMscd5NC199JbqU0v5l0FmDQ20jZJT85XYw//sN4kH+usFzLub/AS
kzn4YY6WCMKI0qS64NAHyG/sAgsQfH6XfhIxTl8Ei/buoERuk1T8EwJGgNhr
mx9diKeZvPMUI95h8KdwB8JnM+J4Ii78tO1K/aUOw2y4X9pWhlB0XeP4SrKs
1VpBKSQ3nJF+IZvHG58MPWouF+fKY8/JcCggZyAOS+Q4/nSgo7P6oiH/ER0h
BKwoPxKs6Ea2EsKmSGxY1UY3ROWZVhwueQgG1OVuck4V6e5R+xM8T0QM8+b3
YdTcxu4FwQYsCRgen4mEYKU6/3++TcnPv9RK8Nt1hCqLuzU7eJOQQhg1INsp
BE5zS2l9MJOPd4npD0mufjA9jJn8M8YCKMx7/AdnP8QMvGwa5BqMyd4e0U/4
oyym5w+DXTZisu1/WhApaI4/Tx9j3MmMEYcBNsXh/cfUbP6kMc7jj2C24h9S
hXUPnsit1JKRjqLub9l0N+wXIx8QGq+TiskcntgSCb9GCHA80nGpdHXFooI5
FypYoP/a+btmNetITOYFqK0omCAd0ZU09BfFBQM6NPBqKj9ajdU5k7nFNg6o
yKEm/tfbXOvps57KII2lpamFoL2pgGh/LCbn8+uVxLEamSYalqR3WFDac8jt
5Yjile9y01twVhMsuB4HFPm+8gbad2cXJX+c7aM5rLIoC4T0lwKo6aK2xeRs
PqzNttiu1qvbOdE4yLYr8ooss1jsygQ0Df55zHHBdEBhg3jIfVqrdWPi18Xx
ilSkFjNlZ+De/aRaMKW0AqU6unSveR0ED09ZValztcVuVYxaViOhQPtqdQUF
pW35srqXRWalazO7gQmqVJZH/M5Ke3+fLWvfgbeqe4BO02IVXV2N7F5UtkaQ
H+BqALV6YS3jNUGjACi3rRzd0qtPB56z2pM1St5jSmXEAXm3xKP+/Zeq2XmK
hKgYbG7Nxj8d5elv8Y0IjQvpPoVXguaVjsjGMnbE6zUYPtYHhgn5MO8R3uAY
XsEW12Im6h4yKCZhXTY6EmeBEBW7W8pH6L2AtRwSEPwj9s8UKPIwlhRA61xB
Bg+r08y2jhB/uh5oi/j1yePzd78HrUmTzhrLMGkpRjP/3hPlTNcmDpUA9Mpg
1t+DL1gCKF8lnBLHQWNADmramOuSsBLQi+fWvPGVLD7A/xOygx9NBTAAaEyN
s1uuuYzyzq0fD2ydc8mDfpsRMZeMNDa2T9sVsFD6v+8vgIKP/ZZIN7DnjM97
PbtYvWeTbJeaCnieKWPFjN3bWVeh1gpuznOgPTO5z8sGaTTYNzQXEYKjdfWb
3luwWuNAYlbEkswtiQfX+3j0cICAh4krdlCGnpNb7Cbzrgql9TxLdAopoOQr
rft8+2iq5NqKbsqnQaqf8GRYM3YEyo8oOqK8tMrcMM532bXZtdfks7mCm4K0
85lWsJD1Hyyzu0V5a7nXueDRxblzwEcbwECDPjJclTxcexHTB/BT9rDIYd7O
8juUfBjpYqorPa3InWZzSIFEvx4wpkyx6ZmS7j0B8k1mQvVqh66Ur5HeYxyA
n3u+MwF2a8/8efLCvht6oMDFwXZBX6wpCF+tOEQ0bclGBMqCs2g9a038qieE
GZYZ1sKPYwuJVyo2hIFiX77G8CkI2ZU5O7QTctS62hqm6C5VVKyCBuj0rxdm
ERDJ34HtkzuGYK9qh1p5XZyTg39k82eMX+4STATFU7VTqXH6mNrx2bOKs3tH
e34WLuWn8bK69Ts+Y9VbxM2xGFBz27z2b/eJKFSuHevkD5JLmaaurlaBik6h
Uff9/8JNaxU94IWLAgHFbAifDYfPwkQqhExfswK0pfzoDjAxBN0pueirQclB
NlEOJC+DFqfZagAZJymWBJc5LwcvWjDzSou/xddsAiE0BGRWVm46ZjYwjh5u
dQOQmeBHWYrdMRiIp7NRLe8Jj9QstqZEaqqanfn2jhdb7U8v6GKx7xmbObd3
Sq+dXsjsWi0BdmEd0pjWGNu8psjX04PoyNuFqKwWKxlKgOJ3z+z5YniRBgMH
0NXuC0noMFHJhtV1geujxGC86VvR0euzInd62TdWj5Ayb2DzLnAmXSrozqsw
V66KhMo47LdkkoOq5ODbyys2pS3lup+xS4i20/sbugmsPQJfdjzJ7Pf6l/G+
PShPZfziIAYiEmzL14VAz+Wk6RuUX/FZW8GtHzROEomOlyTC3mqakq9Pqgd4
N9xCG96gf7eMGT2zqZtiHWO2KWCG7TcktdcEkckrrzAlZhP+ICsbMTkF2gzv
KUan5PhQC6OJcwGwoEBuRdbjkkfe9zFUbsgWptgiHrNeprxwj45BJzb4/q5T
Ow2npn6iXEPiyhBmsBW/AW1gLhKkGLZCFzrGdspGtd/WvlLyDfg1J6Qytj7/
6PvtGyS3+kXieasqaL2pRWv5T2AOpIxXZIADs7uNho46X+dVE2SVfoEvhCG/
eSAYh4x7/LWgHQZRJfroOMFgpTVnNzW4qyRq6h21IK3sMlrdDuUSILGB4j+S
xyyOSh4LQfCTTmAQs2yy5TBMVuGdP+C3HHK9Ztpl4FejLF8cbcsDabVgAb17
rbCEwojMCArUbHYb+CWTBdOgLuPcJFrrNeqnWui5nqDCX1gSsqiZbUra+SmU
HuIGfQ6YMJzhIosxSxjayXr9YzpGvu842htb8dgmYb7qOwf9OnAArVWKnnhf
JDFx9VoKNN7yWwwYVyHqGKyK1VN3ynBwwEPn+QaEkFPwQSCjUrgz6IKiQdDN
6/9FMG7grMgUcBAqSgsPil4NCsZrStwFx2C/kNnttx4QzeUfoSiadNEULeQW
GiWPkRpcMfosSlVBLsY17HjEkxsJ3rsllysE4Qeo6lvZA2MjEw2ki4twGmNJ
IYEg/2NdeSxOFZXdgDd7Sk1AW/W0yQp9sBcnuQBkZ1f0a20qYQ8/5cEfAPrh
9DwxvUpKJdzvWqPo18w0vYgnX/ovWkciTDk1jUzCOpajzaEd+gyo9WZC4Q+9
6zNQYhc5o/A1NfnzskyrWMnZxijaZGOfyyuMszzteRvaq6dTBoobYZ+h/piq
mMkHfyN7RZFbsi9dIp7hXsJHuDqEOrNYa/45oVkdBV1KqiyEsxKwbih0ZDuA
sfHZHSd9YNJMfnA0iDQU68rbwJ073s6TkfoSLkhbdhBbDC203+ZVMbKQ/vOM
ljXLlblAMBOx0dDZLhdZTItCepQci+Y/wdfeipjCLuS9TjR89CUJCBLGOKNT
SNr0XDFnL++ptUlL10MRmR63DCc1A0IEkRU/eWhD886qY360TOptDtCv5mdL
J8mW/vyN51UFyXXLEnEFupVH9qhxJNk35u1x/mEwtrruPPaVmpLK7DbtCImA
wii9Z1kvAftNAMot20vfVhJ3xyDfMP2s8JE2FhtjUix2uwpTPj9x61ucg5t4
evVjaXHF8Rdi7pfhsYKQnj9R1r3RyDfXO5Fekn1re/c9J9ncXCZ9dCiwlJZx
eczSP+NcIGUyYFmbA2CtD3krNfWLQ1JUhxsgdlPgQzmSKcyrPELyYeKrxLb8
FCDxySS+2F4Fs/8QAriMpbLxV3hdzhRV4CCkc2Q0hv9ocTeO6J7pwp/VD2I/
AjRyQamqSiy9NOtX2kGweu84ExWpl/zMoRXnU4x484XHucAQFsE5IQ7cR3Pf
/9evdJJzcr3ony40qsNdSMf6cehP1U1hquRXqspDk1EeIfwtWb9NcjiwHrOm
SR3MdJRgni4zvi9pJacaIIkYzdYag/VUI+IQ2hygmU1yPoc9+qIUEh8t02XG
LnR2SEEwdDh3nz4FM+BvksqWyxeMPRbQYfg+Z6jFsr82i4WPLCxJ0qXt0RcJ
T+Eo6Jg3c3D1wir+DfvbSnJgekHnxGK115JwjjrYs/nuTHQfX/LcXrX0s2lR
WKrFETz4lnqQO8tSU5SU7WUfuw7Lo3mvEOKT8pcpnanNUD6QlKFhR305axuQ
aNMoGGaNlRG52qdJFsSPe37kRgr8qe0JThuo1J+nBvz4xkzeBdSyzp9/MZdX
8xKwfy4NK65vPUaIBPYuzjpPrkRkElcQ3ssUwdTR6tw41PD+bBQcuAMaWU6U
TSIcxiDFRJasEmKWzndumJLnyFiRt/eN3BfONl5hRk8TV759SxQfXisXw3Og
ByiKxGCPIWnA3T/Q/VeJV7yuqTJtkEmLvGFF8wyYFCulrIdMWSSxD4ZAMMBo
PD4+Z5bC7vo17YvX5UkQW74xvd1LoQ1CIzGu4w1sRJf1Iv9bqaN8WeQjN5fl
3aF9Hv9BJPIk5yU1m5K5MQRo5EIxWxTIvSY5nicbjbnYFnppzvQPdMFkYxWL
kGElWPlxUIbWDaMpUlQ0ohcUkyT+YuCR7DEzQsoeHxZ6wuU4SoYU3wlGesut
pOAYPherqRcFZmiRP1EOQa2HuSZCfL3r+GZnep+LBgXKKhVBuhMGyysHum5a
WVA6ySg/OAf1/ujiy01t15FVyGzQ9vFaCwhk8BkjCKnpeqO51REHF4aKVTCS
U8NZTk830bCFOTP+YkmtCkQQ0pb5aSX0dpO5qacDZpuKoTgT4xOSQ6T4wIVB
rUdcC61K+4QZrOQ/w862gzK/x7yAljRHPy/tX4WoMaOzTUYFNgCUZrSRiXkH
RJA3QEchebTRSVXSsaXgxm4IFV9bnuuIMEMWQUxGF5F32qr20TEL0hFQZMPB
Ay1uYHmpu5EEtN7fhYD6nMdabyEHIY8SJKkxDd2nwMS0k215PBcBydepgxzL
Qlpwxha9lDQxwacHXfVVciQgn9SlJxoSj6wHNNg0IqjqAX9tj5ScqPzWMciQ
dq5hRgGHHD5a2zQHW/Nqrvq8X+gvZhvOOaCymKQrHyNY1V2ydTaS1AEkhDus
gJh0Ox/vldnTtmuiq3BAXTI5KxV0aeh7H1Vp+b1j1P29+iwAynlTWo3FbSOc
uMt3RB5Ht3yzPS+3lEfdNlJUQeM3kXv4BWnR6VMx+ZtGD9RX7tI7LvXGsz05
+QMUxvW3z0bPcfFjZPdSzb7bZf8NL7Hf/sf7pH1vFM2etKz50k/H+6Qp5V5p
Htm0M/GhAv/oeQqTe51TouMgUz0mmfKLxAq2pZ3XWVJJtpFKdQtIvSD4L25F
X8w6ClJIXsjX+wbR/Mu4t/5IcJ4UHi8yOz7GwUc3QGUZS18vw7m6tPLzAg9T
a7bOqGHJ6pepI6yZ1bgZ9LQQEqc2Kq2m60Qf8l2ZqfU8WKk/nkXqH/OGfvOw
ASx/NCl9AlAaBs13O6NPayD1LqYz7KcuB7GBEwB//j7AEypMN1RGajtjN6Hn
aYIcROX8I7QN0rCernvWsSkHqD6t41MIjLmIrdK0p48NhPaCzNprtewBJq/k
ZQmJMe9qz9ZMvL7ZUmiJnOULE00GWVrdVWah5XEwmj5AxXP5iXs2tiO/ZO8V
VInPO90CwzKpbDEzXaSyHefw18+/biu4uVFbMFyBP/EX6WqL4I1Sm2qecKZF
DpRWjIXQYt/yZHEju6nxbbSTCfJK02D/F1Se4Mlr0XSWHcJWGj/n3xTm28KU
S17Pccb+rGo9DOWVzBBUFUfQK0gtD6ymlq/R31x1LdoSjXGSia9sfweer4bL
b1q+mdCfSkqFzi/blay0w/38XIJcFjHCX7ssLgSbrVuFRoO+b6/0H2ei4DjJ
Vc+nAvK8KwdqFccldYoFZ082i4WiiFQCp6q2yA5KmOzaJnF1Jp3+PhDwCLec
RI7TrECAVy85/GY/fqbC/ks3WVwkI5Dcs7gsYn3rXAHRkS+OTvBLXmr8Z9vk
S4ZBfcKPf2fnR+Moco/sbn68ANSOkhcYAV/HWFyk7hlMKHmLghQ/CbTlR9zs
AGZ1REUWBIH+OWFPRGIgcyKfhwrjghcK8jKOkk8m8mZ45ah50SvAh4v9GoiZ
MUqKgGB221IGDAACXedBH3ApDBABAflH8QtkpuIrm6Yy7JKh9cfAumyDXwYG
E3HPu38PCX/0jWdnZKiAd5XHKqpi5sdsbjSLCaZF12jlMn+OlXDj61qvbf9P
V4igYK86bw6r8D1KHtVJJsQA1uzLfeKEpcHLOwJj9GpMhC8J+13jC+9rFgTj
nFZh3gHFxJxcklgkM68kxWpCJJM2xNNmKT4kHhjU9vqIPVqdunRNkyweRj+h
ZSQfMiKhliu4DF09YFd/9acoC3zbxvyPquDGsBwy353biMqnc0TFU8aNL6CO
oJYI79mNVEwUtkhj8cdxIJ1yVF/yVDQ6xDq+lwAKQ+/LwreNjDNunqaxc4pE
tKgDrtQPVbhpf8Zj0k4Wl/TjPuNBOpRj9wpOZEu8q934oknZJVxLupDCoz22
twiopZrJhOTGUNk7+J4/xiwvFAfy6J4xN701Oy4eqFYpgoN76ssIQe7NRc6e
7fuVjDMayyaue3iCVgrSrFE9qZXntI4RQWN2T5f6qZBJWBiogKly55RiuhqK
nDfWuLbIgtaxCDQkAZNYRkvcgj7k9+hACcw4z4EEYRGMX4KufKOFdMbsw7wx
IJ5kMLJ9hQeyiDnqd1YOpL3KUJrYfZtfUPqvTWWMkz6R6arsegGaK67Ak40j
agvnToaBHdxmeuwb6+ST3tXOmyFd5KhdxQR4YDH/h796HgolAjiaSDH9MSpz
deWoLsxeiToic3lLA+MsV3i7A7SSk2NZVplTMhZEE2b83C2C/N5oFsrRMiUN
C6kJJgos38Henaapb9NFiuEdX7Q93mA1k/av90zxZZJuRofdma2tCaPmkDq6
isOoj4sA5x4l1wGXdb2Bnt1drZaP9Ys9kce3QoT8OkcbuGuHDqYcXeHJLrPA
+ScYhH4RolK/y11tBYnZdUriaYGvNodHtS/Dcljq5dbpSwduIh+KkxbPZYEe
bquBXHastNM2jLCW9a4qxqWdLh6vY66x2aLXqp7vYdutAZBa0VMU7fb0Aueb
xFIgVJUEPYwOSXj/dj71zk9aIfJW3tVmaefMTl1eq+C9rEeSoFl3hIFNwqLt
F0QrqO3tmDfNDYAc2v+9aT2p2CaLDAr4eobnGGz5nnkOHFIksmQURMp0+2y+
nazxL6ANk7TIGZHllBon778rFe0+9w4LpkjMSkJNpY18Tib+TOxQdGKsgpYu
rLgVIkBoJ1uMejYX+RZpYydA1e/qJT8yQw0w36vy6lAPQnsLLphd7X3odIPx
f0mMJik5fE5Z3XWy2h7F5+crb3cX/uZTLD80wu3bRDi71TQrmLDpaygQwc3a
ptSJ+mdkgOOZug2Pt/4Mc2rJXOpm8RefETThqCSZZY+/wbDkQ6iXWYG/r2jw
NBbQsqDn9kvGswQCGJJM65ptpOow2qF710mU4ojFrsTAqPMsuW0RBcjIcdFx
OM8A599xAUZZg24W+G3tZqidvXmVZyB5+O8Gmw0c3dQL6NAVqG8jU5YWsYXR
9CDvW90UA/qnSIdYmJKYqVqRVEQ2JuLfbs6sXqFoxMvF1AkFDrhm+oA4AmUz
2khGufGfkZfeLAhefmuOme6lHlGbgkf2QLVVM3uKyW2bH7ZwDSlNUj2CZrj3
2yQJdKSZD2aZb0ap1BzOUdXpxK+ViKdYs5nLCd19dNF5TSrQO469AmU+saZt
LDCh4wX+4TGSeho4CD/VINptRUrPWKcZ+x/f4LRXeq01g5/YLbfu5s5Jyibq
xDdhhTOrNChBiERRixJHtl8KuovgWG4NiR3Dmjj9fxLacfzyMg2uajuqH9I0
S4uSNoySDpcaQLvndjP/AlJgeZh3BFYHg2mpG4egotpgdq/UWJrdUoseG1Ox
fOa274a2SX1vzUd1HiqcZvDH5JdDui6AES7Z/wxAp4wajhkxVbkT97DOL6Mw
YKzkYfP89c/F75QywjXBFZmB7JrMut2YTMQWHAz7G7Eo0OX4qjWAYAmGUuTG
0SgC+XWjNsyg9kOd4oOuiVLQ0p1faCLn8XmQkFI0beCeNNs2hOTloXK/GX9I
p4Z1UnR6I8sOrQLDA2UmXdEtmeJDh8g6PFq57Mk+7nl3khxvlj1h5vBNs9IG
W+hAadgJlp3Phic3boavJ3UgtUK/gxI2KXWcN1PgwzRZDmWH8j3nFK3KqNrU
jAbrbsV8f2MpCTCPJHPxBuVnX0NF+2ai4xqJsaTU2BgoBxNrzxPlpykMBlZU
SUekBjiztAx3R5op127QysZA5EJ9BlPhxDJcx4RaUFu0lJldheHIl7+7H8sv
IEtACWcLE+DMgrP6tOucpMV7ck5mUKAogODMKbD1kKieJ2G3c77gMVeEm5IC
LXynamKFYopJ2TAmPhZe/7oE02vj3G47f98dUgrd7lh0YaRAIu2Ytt9LKoAa
vS0l8NqW0ifFUzmZ3XmAgTYalOw6wuUbWfCP5oQ2zg4er3kKIVPSdMqLfyMG
q/WiqFI1AsCYiR2TZwTOoK/CqRTOD+q/WSCuA6DEcIU3Bav1GiZ1bfRyf1Gy
lXBcRfGCGm/4ftyqiQILIRE6xmqHiUX84mR6kRver+1FaPJxqtZMz+cPx8o0
17YxTP3RqMb2dPDiO7pYGDRsFUBSh9XOs9KaLC7NEZjya75tiSzIxLg8XvM1
y2go9B/j59YiHioBpPByFDr+reTEaVK1rY5Oz2ijdtaOp+dHc8EW4xiElDku
EryBrL6+nwcCOSZCroLzdlDsB9hQJi2VzjZVcpZ1T41ZKmu9nUUZA1lgFvQ1
mI9iJxO3mDzvH30DqSzCpcJWK7B9no1lo7V0IcjtwWfKfAvzmEC1RwMHQq4e
PXPdgKTNDiwYkC6PcakzLaKHJdELv61QdNspf2pyAIjHWwyNsw3HG1/zS+bU
vCK8f/kPkPMqJUxZ+2sWGZGBmq4dkG5YtIfeIqxrxiWbrNevrTYjbYszBaZ1
P3XYAHRFU+XcGrLJzl49OUa6SC7rC/e+fP4sdIgmFn50HyDOfjEqHT8/biS3
vYD4IDz2Z+Bq0n70yrQkE9fkIShTtf5FEEl7La36B5AbwXk5BZFcn3FNZxZ4
m+H7zkfsc6W9ulyflonehP/IIVHuVwNibuRZC/is4nO7DNt9DvZ4W2DLP25B
n2cvy3AkYUlbe4x6KCUoyAem3Kog2hcL7xn1KIqYtradntcWUvdX5eJvJ/kV
RJpHhfvXJVOhBksB55KPGObY2DrZy19DTkCbEiqXZtQJ5GADLAMCBRmSGiTE
iC3CeOVMCPE0G5bFG8qXd4dH67o7bzNL93FehLXWXcUK3ZIO9QGj2BERCm33
Y1TcrLffmYm/1Hn3ZgTMZZUO2XgtZZpYZ+fiSWi0v99B/kSMJGf0U6yZDjf+
XSOgmLF+F9pRxFEFECJzkEKI4FTo9qyIJ8imBehddzD6Bu9SpzBZ6jQ2FqQM
evZTiLKZuLWFNJkLryfo+zEHO1Qib7vWCCwqH5Y3hwlWU9nfg9jQkIHEFgEk
jq+RTqDHSZZez5Cbx6Mn528hlyKDkqNGwHQOnDYO0OlBOPwApfWoO4VKPoE/
u77uOFgol8TlEXS6DvrtSANO5fG3qICFEYW1SOtAIfGcyCTCZkjnOlpBkiF4
a66AjBKJci/bbzLQlCGlqDWeztGBeU0gy+bVAcZhsL1VDMr2ERA7UlfQsGDf
SIMWRbgvWbxRaFGXhzS+hiXErm5Rn9IJek8mhpXxASDnNJLo4HFSaptK5Wn1
jqZX3cDsozLDsde50Nx4mf/J3mZHcZ2j1B4pNlUDInDMm8GhBeIkxnxBTq2/
4/DEm5SBxBupin8jj9zlCACCyOt6PYoioRjTGyZ/WKwJsFM2amCBHGPKNmar
rA8VS1um4fKGZyuh+V1KcdM8DiKp7GeTH5xGl1B75PmtsINqMc5cdavhHLar
4hGik+Nr0Unp1XHzEMDa4jlvorFwNHpHvuWSdSSjAByIaS2MJtlbPfXh1kEr
nllsH6AcbBktQ3AmFnWtHTrPbsnHL67Voe81ztj1cA3vjAf/YZWRNGrEy/8u
Q9mRarapVBV2dkJ4FUi8pDny0dVlcuHce0m3C9ZbrAjOlZfpVdriuGQGP1Vg
vkt1D625f1fOc0M/uv8/FupaD6UoPqDQr3VTmS+FljqoeU2yK+Zismi3i/Ho
SzyEfbuKf8WlgGXK7KQ+qrNbTiYcLmZ7i+51HacYekv50ljR8eZCtPumo5Lh
jSgIiLDv384QGXjD6ucf1CjZKBEoGQHzJrRCZE2UAQ7GF0APSYdruHXWB8Mh
CNV0Gl7ChTFpR30yK+vV4M6zufGz3X7ixHCh52GK3+KmL/YsQW2HWUIB+7L0
AI6T7ybIfL6S2914pYedUo6LFZP6ih2k72RIJ03vfefAAg2cDvETv7KMZGkh
Zq2srgyce8eicb51P1bSOe0peXMhGHzj2Cy8JmUyCPT5fJmxJg31M0hN+m/Y
fRdcYcZHTwsXhKgY/qdbGUQ3B9e6QsxUfmfLOBUv+zh8jGsajpSYk3QSw4qy
QmVZoqvxrhPvyqtkH3BSSq/ZThOs0OSPYEX5atcKZPGYa1uNT4eSzJ8SFkhw
MgOf61iKq8kwO4DCE5MA/YpWSj5p8BKukfkJyLtKkpfkIuufyXYEEl6Tmr8R
y7wS3VuuFtBc5vhJe9X37a95rWJ9VMDmI8VFn0oudBerLGQ1KfI8QgLHhuIi
xt8BUBh6vzVWVvCiFg2paY8LSfau1vK5Pu0IcuzdaPLRjD2hgKeZqkLo9BfS
dfTON62+N5hVx1+uepQuj1NkKOu0uR8mq/vSS+PZtdldHw8N1GzpB6brvvZ1
WmBJqv8RDwMjRGBsh5XQ/1etWESAUYFuHDxmycWF3nfGyn2gnU9RwQ2r7HSK
0uHJ/esY3a6z0R4IUTUcryzRWpGXXNZzK4hNhzj4i3m6IGJdWByABcqVBffm
ROA45K5NTIWBM9YDvLapdPkoa+DYYwHOid+ZffnW4ECXlBSbgFyVvhPY8s1f
9sZh7U71u5yrwL1szCnpxl7yukLRAPqel0IeMjZKJbzKauR58dwnDUP25TZX
/ezGAIx77PbHF+fxCCl2fNgRHtKIq1g77PrE9EfP32FzJR8l729CWnNaTX79
rfGPG7RvCF12yoMIOUtIhUmqPdy9Av2WEvjiUr9uA4bOn0Rkl1BUon9FcVHN
i+QeAtI5qLE6/376YLEs6JXVyOCscWd0w7vZMmRApd/D45XnEOWgoQiTIUFi
7J1iGOmtWlKcPcnq1cZEgQr4v0Yp6qEU2Fv1+CUSDO+aQbXdesdk4fbWrdll
15ypX43qZ9feew9wMzCsu6uAWyahtFAszz7MogtLs3UhIRbQpExo4YAMYVX1
qL+Hn/A7Dc2I+lPko4s1MEKYtAMOrra03BzynXjPnGhuKTd2vccitq+5vt83
drDSduCWmCcADf92bnq4QhuurmxlwRl60ngg9u7pOX0rImbBjVrhEPKdFw2J
4F+/r3YH7RJALobq8NaiMZTWDjsxYOsN5dywFgmp83hWDuWbW6jiORhaiVSJ
qV+bPszGJysfAJxOaMcxrMHjDVPfC1Cejm8qOLE9gHKaGhX2uTPcftfE8lGa
l0ZbstHYeZD+0MeKBW5e83zQxqGJumG/SlaAJrVnf3xr6YWNvnBkeoHSn3ZV
UCaZxycA9FOKgj2ykHn6oflyqgpuz8kA552Rtsy0hSRKyqyp/6WwLxj23ocJ
0Tp3Tks0TQ8cU11c7HtTrr/g3Sz9q9kMqmVLc4gej5AHr0vCu8Wf4mCut7Yx
J970Bb8RrBRMJicYeKEyUuWz4zp+vXTx8vShirFuxEOZ007w/+fOuKdFqUjd
6IDKQImlO9zWShV4oy/51lvKH184XIAWMcDhyjeH3YHqewmgWkS/33law/D/
PSj51kS3pGeXy5HttmGFIDrn7FLgTUusTQ75NgHskJOeWwVUVm21/FWG4Joz
vwkzSPje/rurlNo2Dr+T49PntrbDcRxRdmli8qAJ83RdKgY0cI43B5DOew8c
gvDE3OseCJwZHbBA5RyHLBGJ1RxenWnNyn2+K1Ig7+5plNPj2bAOpar8Bk4z
n17Hg5EK20mGwWxFuCj9et2SMzoJMzPhhKYfazkBJ75eXRKlO5rsZXaqiRww
4riLwGqubUr73qRCKe2ztn8WtXA/wzMA+yvvm6qFlfrJpoKUH2Kw7AchSvuf
DHFrJwE+EVjzbLGvDnxiPN0kYDFl7lbwNUW3MiB2qrZxHU1vR8ON2ahQ7uGs
h3p4/19iS0tz6NeEO+yb3oom51qQ8lnbg+mZFmSrTGNM75XjQj8I3+/s6wXF
4t8722ZXcT5yw5wPv4+0322Tvpwg6qZ/4rEKOB69XKVYntIZIBZkiTV/jEkG
3LGkGbopi1y47jwIbktqQO8FcISwbI3MvDqgMPML3yWHIOSFht4XglzQ7M5P
o4oTOSH5JL2dPnSO47LqvwALdDF1F0h3GOvs8t+UcVpJdYRY65+fR34Hjryt
AZdMvasjO3Tzu0kos2fXJ9gP66n5bFy6h3jzO7fWTTo9YlHrWz3pAw3lwzf/
45SBcYjzNYx4EgcdgNnKSakHyF+av8QsskSLMJxNCwfh43TikbpsXDsKTYaB
ZM6Ufuc5IHVMHlaTirk84q59yyRr/MsBOPvKV/dxNTiND397YuD+jmfv70r0
5Umh5Zj2mEUvKc5OaOvftBxW1DRyjEXOMH8Dd/bW/WLeazyYIa85ELj+WTTW
NZXICj79zp/3uVIGb1Z2LnkKJafz6814g6YD21wUMQEZc3QM5qFd5MmOTijm
8F5FcWEbS0Ig7b3u4k1R5ZjsyMLlfXXml3hf6lGnUgxVUn3jzhaODu45PTaA
L/g2ii3RAAs+jWWyLZOsIBiooZ2oWlmIxaIuJO2fnsp5x48c+gMo3VTkXUTQ
XqkDkZryS7bNQzqp4mH8BA8mEIBzWA0sVtoLhm/1h/LCjNOUVI3s/nXn6iFv
A7UGWfkBHlqB5QsAKr8ZmMyZhvFTmjwcztZNGUxC7LVulvxJHki11XvKG3Sv
xEcZ7zq6zycPIyi1vH9PIRRJIiw/1+NwC3sCB80WOdpA3/G8Y6mW2HadF/0S
W5Z0PKQNw+bd0I5e/pxHrZFwV/TzCI1CebCbgVoH84DOK3aJL/REb1kdb1Q8
CZfhR8tEPDvJ5my4xuI1Bh6rPN0be9YcRJZmgfBwivrbpPfyyce2sXfKpsyu
WVWs0NwbSu/y9SLeRQvGg6GG2D4YMyxViwsF+GMaQyjCagZIva0EubPm9itA
4rzvFjaz53HTf/CA0LsY7kneHVLHpzBKpCjSrOpoCOP2avOamJhL7gPQIKA3
Laeb9W1QLN486J71mU4u5pkIhxjOxiT21p14jGzRKsylpc4Qgu26xTpMOIsa
BOx8JuWbCWvB8xGFPH0QIF7mcP91MbZrH2tLXaIiYBOcmJEy83fqlWWPGoo+
8iBDYTKUzPWrLCGquMijsnKyW/Ww1gMTWY480xJtI0/MB+L2XJVdP6uOL7DG
RP0LAnMNkhYOi6mms0fVuh6m3Ec22miCXpK4GHLIGyaeBKGiQ8debQ82Asnw
cBTDq0Vg6wGIBFqXcTIF/syNFGzTO5NQkZaPftvBsFirJlKGX1J6Iflw0j7e
Gq8xBCLpFovnKpG1hXhBhteOwk/iOqbUH3NOGPOHPomHhEXuGIJYtgvq3ziL
3rixv0/xrQ1ZJrObQozhCGkXliRaEq89SBXTAmAMCOVo5XcpqcfveiUyOjdq
bcEdjPl9xYP82b4D3iXW3lA4RkuLMIQAxbi11UL4qHnfE2rAw/YDvi3ycFfu
rxrXGpwa28mwfnW5lX1Vazi85Xq+DFSZhTKohwECY3/3LrPLUlin4keGnY0a
FD7LjUar5U9dYGc5IIHe2ZljuqJNu4LQ0wgDHIUm3n8Ncc9E5I0YWuCOCNPU
Fef+//CSisia1Igm590VBNKEwnDq+I4cDHacJIvt0+BZJEf6Ooix0LNNb0Rj
AZikFUcLLDhHDiP2+PWBFD0tc5eawoZ0pMJ2LRawWuv9cea2AaxZjWG20BTy
RlN2pMnSZ72CmbZXiqLXPtOdpLrswztJFKvFomClyTjAQeHMz6W8VEIKkq8K
FjVNfhF3Iml20krBiZQ3fB1CKq2L23u+EZ4+XGM7ps9Zejw5hsMP0cH3GPDz
aK/2DIeP8yhtT4KOO+fkXY2FS4PrpBsSDiWuWY+3ryrxmpQmu71XQVDCZZTK
NMDQJGK0aNbEd9mSdbyfiUY7rxoiwBqB6eQMta40+U31so+izHiReREy+PJP
bNunNwuGb6PvpXco+jJZimbDaHlHXSybjiaI97J62DK+Owp3fM+Rtktlp/fM
BfBur+32RO8xBoyWF/BvEoZRUj4qiekvL0gMuNLVx/TjVrKJT/cFkpzqgzSv
yflm6HiReQiQi8lfYWl2e4DVGguMv7JkJX+ligvb9IciRsu1JsONouUM56Sd
iMuFUXtLlC/Lk5xVI9HPCAYgblhO0d+DVEUNA4l2XixTla6/pmY5NhPo/H26
3M8ItswoDzXNnMVGhT+UWSUJC28ZSpkvPrEhquwn5QMVOWQaHvBJsp/Dvyg5
RLd0/bpyKJ1RxD+OlMYoM1pCLeQcZCvmvxKJ5PBf0e18y+Lm+9finndLDhqI
GLmsoXgj446HU57VmlQxlhScOYLjAuM81wBNCCadRa1OynCruFGY8Qsz3Kos
La0tfhVpivVIErFgROivlOrmd2X8cZDs3hiJYSVlIabc++ZrDZqKHUzxzCdn
3DfxfFemvnQ//X1VQYEDsqQ/mS3GIQLUAKCKXQHNWmmJum4VWYUIaXqbIYcr
pmmj9Gdv3oKl5R1FQqQfMkV+0QV5McqRil+7QOLwuBceoE6c02DUjoJXzOVE
NAny5SrLhe3jutd6pMh4zJ/7zV/VJCI+WcATQmHvMgK2cLJ6GxGvNbm59rTW
BJ5eFu5ewh2x0ydxKs3kTWF84rvjkeode+ZzDzQmjbA8YUuQPQOZJghA9Fd6
KhA4ZTR+QlIId49o0348W6XWu63BqQ2sluqJOSNqRm7W7lrVn0Rh+fuSp085
MFrB54ldoT2S5bey4itTZXkzeESlHRS+gDJ98cOPsqJ0PGPImToYKB7MguRW
uw/bqDQ/zmQSyA1jicHH7M+r44ScJmr50VaCtO36WCpVMJEq1eE/LaeuFTwB
FZaXU+WOceCe7EmOMQQyKMlpNZYjpt6D4CJawk4Wj5tW0+8mgPXmVjvtKsCN
AHbSFlkdF2jYm6GDW/CIkg8AepvF3L0C3u0u6/5MllMcEcBZcygZcRjLtLsp
XqrWXyxaOBWxWn3aRldBiZMsiwXJoLc2bAdGt+hEVcSu1lk8vpmJdmuCINew
lSFvm5N7yY8qpai8PEccqA5p9IMJIEO42v9Vu4GT4gAvLYge7HyHGixKGgOn
IjJUUvn4i3qxR4SnC36hppG2+wMivVnc453ehh+eITsWjvSiBk8Uus8akYZc
qwKvk8BZHUvAWL+nrvUxZzIftrHNHTSkaeDUhU+eZWy3gZGvGOLZoOwdRTX/
vrDyOq1YVR4eSxKirhn4GKk53PKj7+MMgngw/GYtbHRc6r9tiBtCDc+myXvc
tcv9Ny4jYPngZdnS893pqIVS2OSBgzfdyRflIg5ZLnOqv+eZfKmcpcc1Crb7
pH1ny5tnMhkLKKylttB0/MnZMw4/9J7VoYtWuoPocXOxwgIx/V6SpRWffPPm
dWi/2qcbU2syUbIBjfmLWbDIDvghV7USSSf9Yi5IXgAzE50pXajKXRHtunNq
6XBwbEQgGj5fwqTzUyOQdBDJvOl0K46fjxNNzUXbbzCKbotim6bbNBdmGhM0
Ad+B0T8FfXmBYGQn8FAo7SgsUOuoJsuXArfrPlsYP3q6ZucMDJ7MVHo7szsm
U4kKf+FQzJ/50Xgq2bsCuPArtBCWGjfjXcgJr6xuwc4xulS1U8rNWEJ2mRFU
zvfRIMr8UaRQJi4r5A5LKRsAUPKY8iRPsL532ETOPDaWZEU058dh/Gk6PZTx
tLACQ6t1S5Tgocnf1SPJM3Rr0iTsa3czeIoPKG4leeck82Jo98LeeSd/gWEC
qcN+dyJEGxH46AlXKz9PnBPq42mlHc70KZLjT+E7xQ/yyiLKOuSItyim5lcq
p21BYmYYiHaRcPk3XKZ6/aYuz2Zsg69pGXWqMfkvV1wIvZi4VBYOVLWGRBOA
ah5I+6/WrDjRHDPq9lJWYtY4sRlt31Hl4m2xRkLS0m4MhQqNt+ddd2VGGufm
B7oLUmqYOsQEqcEqY8OiRLG+pTIni7dDy4/2m3lIJGqRJMKIgH7k926KTtOV
TDzBGuK3bPjZZEFMIWcKqsROXeZAYL94aDb6DP8IB7AXiEWkO1FaBiJfMLyc
oo/k5jGt0QshoE8u17yPqeGrNxkVHBJ/zRcp2xgaGRGyEjOCtGTVOwzjt6g5
Si9CfXDYKyVUxQOavfHoGwe4IdKCeNTUvCPsUihS9HfY0uwPgJtmjoqE9tPA
cmJ+4EbmDNyhmt7gEjGMLnsOcMkWEfjciVgNDn77MOYdJbiZwB6XmkvNun+G
vk789LnX/zYNzKjAa8UIvfduwS38vj9sB7lMvaHvs7H4qHAUlO4SHstaZfwC
IbnOwn8JkaWWFCqOhPx0REc2iE1T2ShRq1O1PjqUBJR66sE04Fnrd/YVkZzE
Goa7tUBwhUTv+Rffn9qI+s8+X9pY/gst3yDnlLbBAxhD2kDAQK78o8j9xEt5
de2hsdw0InODm7hgAGdE8WWHYgoTzWCLyEPMFOrTy3u5MSBom8lbYnmXb/cy
zx1CujNIMSnQiKy5RxANAqZsVDUsBhvZqpxBw1kocTV29hf6uAovmA1xl37L
0xAQCf9mMPK8lf/hqz28sh7EMKfmnOeZfOXPeSPAI938OlYvT4qQjOc7Z9sL
gC9lwigikVnXjWSmpJTkG9ubYo5GTzm58Xy/1ZizTTiYbIVALAIwLikeS6bQ
IxIG2JuJaHl2npW3DP9HjWP1ymf8Pr7y5OokibTTjKyH5FDSGHNrhZQQnIdK
m+IQ23CkGVhPxRVMr00vR/5U8fvM38zPY/uF3P6vN+0agnoncYcbQswsJ0jB
UNGfRd69I3nZGA0eBl392wkKP4ozVdtHBr6VMSA2fbBtFwUPio2NpZq8ziyU
4DoVbLijDq/PrBTy1giq4+zCnZPSBjr+NDyMeiXAOoBm7U4NGoHCHDb4lEOW
fHWqsjkNYI7txvu73O4EHVcUoIoTNQDmRYdq2MTeOAE5hw1YobmLz1PNNWHJ
lLQGSfctQxMiwSGaXL9iwibdjgk2iWU9LB3xWyQSRtiXtze6QZhyYPKw8m5g
op5ncb0W8/V4AGl+dL1FXWHvI7XtDab4EXj1b891bKxHJ4oNpTTnxd8OiQi3
8EYTIH4jGkXlMT/t9scYOmIeQq1OaxvtlRxaI5WDPvh3i7NmePRoWmODZ56f
7BpE7nnzWKl43+nPcv8KGYMKIR0tecftnjSExwPwYs7AGagZXOXAXREtotdy
Hh7X0lR5tBuoULSt/l61QFaQsMWhfc+GOSe0+Lb1SYzXV8PTD969MsXj42uV
Z6uernOAeGMG4GBbd+ucLneBMP2CsJtXRbKLY25YAwD6r57fXXDuShtQZ9v1
4QbZI2twgJ6gsTY/v+BtUDjm2hePJozHsSFzS/bhEFw+0ev1QCwsvzE60Sn7
ntCvlOhjOW8sljALhSMOEvyEoCVJZGwrU4fOFo4SZx5xI4yp1IfArSaNA4Ef
Wb2jGlMOI5wQ0ZEEWeq4Sf3EbccuyDej/JITVVP+wu84tC9NdFOLohmK19oz
o2gqHB2LxtxqR9TDbNLg2spn6rN20hgcI//OQ3oznJ3NFAKQ4Qoi81WHsHBL
zvlrbX//Fq3yRqU64FgG1XAF39MToLd/g1tGhGiX4T0osoYGfx5kNJGOWTDU
etjmZpZtb2PD7iL2JiLaMFSTH2Z8ZLmOj6hbQFZ9ypneAotm57WJdsfNaK1X
wAvIb/yFezJp9B/PzpH6OyPUXjgWQ4eOpPtfQpXyPhMdS+auK31Jszx0EZ4D
6xcakfDSpAQhaTYiBK9D5kbIbMWumpCbK+aWMVx9Zw29eG66JCGnc5x/41fU
n4i+zaezhR3oCmzCgX67SRO2VMyrTi9XfXa47hCeLTxH0uzAN9umVHhEqJ2z
/ktZRZrqQny3DaEFL3Wdd2OLa2tyX2i8p5xDR9CgB9+OVHU5Qy9dHu/sN3b5
9uRV6dVqUVoa/pVKvtfyJkZiRWxz+n0DckRqG2ozEAiDOTSro00liHs/Jtuh
D9ut+kU+Tto4oacVibpbDOtWWOTVBQj2ebyWnuJKvvJP3ptuZEEAaJJMkjrF
Pmvx2bUbugYyXPG7pgXfIQADrMVjdD3XcQgEmXMos0AeiD342BoH+qQ35+QZ
U1l25N3DmWWCOg0LrrxrRCtYDTBR6Ke+6UxO2VkmYE8GJ61IkQZTVS2lU12B
jEz1eWoQA5tkYSa/99u/zXn5SI2u67z4xTNhL4O6EUvFfeQBNV3Hokgd061p
TcWA72dOKxbI8+kV9ky2S/VfPJ8VI1M53oqacnFU567FeFqB7WbItX1iKurJ
cTrRkeQcRJo8ujg8106bkCZW8No44g5swTOvAVD2dX7ZsCIbwEa0XQdTQw6x
dHp0uXkWgiZBa440vCd7KzolMQb+rhhy60k4mW5vLki8UHkqDIC81ossZ0Dl
HciRD+5DC2M6SGBI4tHsXzDxmYc/H+34eQigEJFhwPo08+zt6VsbTyPnYZA9
RAudu3HaMoouEdjYmpoK95/GfVICsT5amT9QIZDZT5XsMRc+KZpnymccDdMd
Mt2UW5xJ3NO6p0Za3qV3DTGqdoq46hTzHSNVzV7+OZ1f5qJrXNB9gePAuK4a
1SHNFEz7/6Zpw1guh696xweM1RJkTnnOVVQCpZbx+QmPxeNZjrxh6xzH9+uq
BAqGH50WJ/On7/olKXq2rHv1yp9W0mcZO2CZal0p+uvBV+0wBJD9ifOyCaeM
YRV+6xI5G/LUGR3u08+jPNS0cpwb5p8Sg3FcWW6oF3wSAKNpzFVj/1x+oK2s
ZRBE5KPni+LEI2ebt/grLHCpwOjSs756xbmCbys4YmKQhG6Ayp+D7oOSKyKB
RcWh29Pf2bMnRucrypQ2CxevVqIb/b1FJlRVQGDZohI2WEbJC8wKMVdR+B+D
KPyrIffPtBGGgtOm8bbAIBHjAoNYtpOVo8AsTcezRB++o6pPonZMgkJ9JZlm
BJHpjDAGhS/23bvAJ2/a/vqHGC+s3pUpIXDo9WePVwomKjwjGjc+Iuug9pJY
Ub74RFf2EhbcoC/ZONGdMkizPMRAVj05YJC2amqzfN2ll5hMCjFIYRBhpVwa
AYxoMlgOjdWS/19ULrDLDG66nZ3Auo94s29p0mB7DkTfI26Xm1Bn5a+ZGB5y
sb/3AD3Dzhl/K8V+7xKjVYZZIo3StU2OIYtqcotoU0kuryurlP/P+GO+S4gg
5HBsNlmXwHWHriKh6CPyjgp2dhdEbI5/NCHbhnLB3ijE2O1J/rO2OHTW4C8A
p4WGR0bxzEZl9+kwesd5DRN5CRG/iQDrqJQcZeQ1NWoClAhckTRdikw7vKo7
+WYcZMbPMZRE6umNRPJRmAOoo1cNkbgNSMkQsG7URlJfz32IrHZ8lN/Efr7I
QugcjEI7eaKyGcyWSPSBlsrYs4D42cLrtFYkcDSzLuv7wMzMNKn/dDqwgHLR
dURs5+azhcVISX0b1uwEilhvulPi4s1tKhQsu82nMJ11t/cMFw1OY1qpHiMb
hxGwJj92lm3dPFkPbS45LCCp5gdvE8ENF4eE8JPlVQhqWPyhWTiiAUxQOb/Z
Z71NsPfxdoL4u467j8fGVDLmddd7jJQaU4kwqWl3WccLnA/AIQckJ+OmRmtO
blIZZ/pbPxP8Uv5UngUDJp4DDVPgwiUqfu8yGjawCM0BCxUbGej0oaZCbtyA
5EnTk/KvGzyGwdvUhCli2xR9Ojj1diD33PKTKQfjcodIwgafnFXCK8h4GH8K
/PoOeQIITnYye8IZTMs0KMndWX0JbLpVjbiTsFLkvxKzp0CH+/Y8cszv3zkI
+AbArhKIXqrmnVcS66MG0P/nJB2jpgSyHGGJnXZHCRwqNO5nki4bNrgnskVX
OTYAjGxF8mfqYsjGq72zGis5EOJEwOeP1OjwJ8KEyo3ANtVYo0K3I8tXk8dv
Cb0/e/NsQZ3GgjB4h7mz9hJmx4TwQqYslDBwN3UHE4hTmSw0H9R+ZvLzyYlT
hVPT61MViuCjOhzlrrzdD42pM5Aq6DyANo8Ex1PDseG6PbePfWJKhCaYvobv
l9I95oMj8L5IOqcP5OIKaKTAN6x5MqxkHRua7xr0pmnTbnSiHueUjZWXEYO4
wf6FrWrId9skObo5mvs+BbX81Guwq/TmqGRoX0o1agN3/Pc58IHnlIZirWDJ
Ff2fb5z9zgOQ1neZEqdfUsZr9zkOrV4al68oH39xyKQ2lpKyNcO0EXHS/utz
VQIyt4bzLvQAKai6DORmZFNidjsTCY1ZozqRm8kQf3ESvTAWoQJFpm0y1PlG
Q0+Up3tGXA8UZqRjh2dsyMA66x/jqB0KeO+EtIjWbEKaRnNP5+moLHV5+i5L
K+g2O41dIYHPkvcMf90OdZA1lZUDj2JGtocsgQFpcn6gWOomzrL/b74RMnyI
TElkRDlHNvofnEWABoz33K3UEz5D+050uurlZ9mwMCLX+9BnAUMU2qSmksm8
NfKsTYNlEDm+l+i4zuuP1eb31sOruiFSTIkSaM0WBxjR+zDyrw/SIj1qccBB
cseXCgpzo3Q/SHCe7W1a2qicLiBzF9+TwkVnuQR8xxEBL3bhytU79DDjuU3b
nyGEQbp0xecXjtzG7A0+76zZDgoGky4wQQ1coL2XL6Y12tcsvwcr/49LVFh0
dM3ELJnJysNl1pvQoNHkl0+/3PdmFsN3b32C6NpTDClKppqItbsGORZlCI6h
Qa35SzCrzhiLhfO3j3k2rNH5v9pNMyUntWteGsxwGutpFdYpQpjMNeUncXP2
eoM4V2maXO8IBGAEATWCf8kJTbRnL8nPOlU0z10a0p2MBCPZBhF+r2YGtrAb
0CKd7bbOJF2g/hT3RRL5wqN/rzEBE4wlCTSeb+dfeLUtWVa7i85oA3RN+wKO
D2SZXQ2HAemFJbLs7iyTYmM1qVjB8NFDsq/vKM10rEByCgMJwUBwhIbERcDP
Z6cNDlXktVwxjhR+Be8OqlXK/YcV32wSCp5aWX4vfAsvDjkAfQ4TqpH5C/lX
qV5kMUQ8etjsLOzFHkYtCMbRlu05JalB00Ol6rrNFyjQpWBhmfwppAVpi2Wo
/xZVZByfHoR7UJZTleOb2ZMLsZqjLx0uvigFKtYbM+dKj1OPb0AdGzICQu9t
eP6ATyRxgfj4RLvZVKuc6CYn0bQG+LMMsSi5QGMyseWGWS9/VLZsMSxxSWz5
XfxQquRfL9ELmT6ys+Nk9Cku11NUWWNIqetjUlt23W9NFtZSGo/S8ufX3Kjs
Wj9sSe2EmllLi+jX72wHZmZB+6632S8uay81dFegzp0Np6XSo6JQUh0Ci7Ek
vCHaRlWj7CeqnMfZ2tnkywNyChWLHCIlt7p2zHwc9xsbqBvCZgAGl/tstBiz
BcEytU6VZB90faHN2LsOAoT1EOOSH8jMggfwuQaOHmOtEWfCsLGKmUJ+XmA5
9dG72FnLW5zTXF4tiMyWgkv1pIdyNF6DwvN2Gfp7Hnf2wj5MgHGV+/1WFO6T
/QLCiSTkg4dvjPn2/uMrG10UTojjGS6IgL0bqy6CPWZSeMvF3Z6wMoiJhL2L
RSRcDqbqt5UDSC1Xb6+nuHcvBbWOUxEs0pzpcZbQRd0IBSYzMh4jCzoIfgP7
zeWmurpHn/xhtpF/jBiGU966IfrNNCQGU3vTZ9F3E5zKymw4Misc7SP5m4AR
vt75npHqg5AUJPRIO18rABMtmpFUSTNTdK/KByQbahVYzgiu8AJBLsnRLa2k
UMZI2Qn7/LDZjRRTihD5+xdGsxkcsVUr123CUM5fb9UkGmwDAIlgNmGI7keb
3pf0lrcK92tzAcay/O7zIRRVt2SotIwwXg+jHxNW/ffDGSDMFid8z/0iQeCR
1GxZpVcvcQZlN0R38ra8y/03dmUmmN2Ki/glf7FcP3qscg/9qbwQmI5Me8cV
yVkjlYIcBBNWz0eAk6fPfdsNOe2Lh8OtV1CXXwG6gSyd4RAtSnQ26h8C4IKO
BM9DveoI6okEmAGpsfwPYhOqz5/EJd+j+vBiI4cGuG/wZelmRlDjCsdPD9uk
GtN4OzWWg5ZTUirfUvM8R4Yy9dnBRzd/jECptU256zrpTgrdo5w0Fds1cPuT
2hIdbTAmZfzpBeAJXszYOX4AI5sNfeo0XFF/fnbUybKLqm/ia5FMMqB59JdO
5dziJ+9WNridLke6iOW+CLsCy3E8tt3gWIy1FVtkpYeF8v1UANMtMv1ARAMt
iBlQl5XRRUaMl+qsGM5lzZA12X+q/fAd5pB1/ttsLcctgc0yeIbfwx0URT1l
vgBctDNRxsJq6VgRz82KMwwQQgicQiB9BHBIzrYYJ9kC2la0DySWUZiyhSUa
O6t1l212F9mboOi8pXIkoVhO1kNtCCJQIP3lHziScObAu8uCS6GIba8r+rX1
zeH/esLjyKC7wAiliUL5+teNSD43y10ESWl82ZlYAvZ5wzTdvaMTdHCZGQQ5
B43FXNJ3tjPjo1cM39O5kwu0pdwQqSK0hxOJS/Dig/ZyGftPZ32fxgrRWVxz
ksD8lB3htKWXeA9euGptpGgTmUflJsPFOp2nhwhFmygHOmt3hnF3VhEngXyr
PMc3Am6h+QzAETlLwOaVjRrmcotePwgAbUhyveVougEuRLHaSHljXvSM80rA
TQPynA4TeHjc2ll4IxvHQ069mv40GxmscEGKsccoxDiRXwkIHDUUky8oJJtB
l8blTsSi/vJNVu6Qf8qKu3Njkh4V/7L64z5xDgj7ywHwxpzTfAsmXGqQHO1J
QVIAK8tzBmCj49j45zlaQbetg536FLKGKNZJM3dEkOsSE1xjX9ghKjh6spAV
LhGldn2nh14sIbYr79jsnjuLO1EI79QkSvV1XvfJ3UcaagzxQv1vlEfT1xHE
nMCE3co7x5bXxEV2E9br7NLW8ugEIYcMV1hOvs+yfcbZeZ0cIC4HpRl3jdmM
fKoMnuRb2DwHJwHtO8Px/qv9cB8etd+VLCyt2BmZsGRTEssETIHG7TP0SLJR
XdpbiH55tmJz0mNm8jbxmHdvi7PMw2r6ZZH2tZydNi6F6jHQ4IrAGAcq5SEE
blejjtG05HgD56NCojDBzrjNnSGeEMgRXsDyhxyWndVCR6YXY/tpp1t2Xrof
OOOawqkH30h6bLB97/LRmykKx/YQwqD6bv3/sKZTUpPfToA+X0D9HInaMKAM
Vae/FwUpyg/jNjsHcKfvVGcLAhU5vIkS8PJIc7nKmnOjRbOXoB1E1bm6zwqC
+QBORVzkizOXD/7o1bmv1vNjV2oj8yGsP+754OtRLgmO8ExXCZLIxJ5h2NVi
ddy3Tz8bY0/2nx4CGe3M26tEaO4sXhHZyk68UVwVd5HQa1UvUie3jEQrtWYg
GMBVJ/85xpW9BoKlD9pGmaVL6/L86wm+Yms6gR/9sKQyP7B9jO5wWdTN9LwS
1+PkZXD7P3wTowPHCyzu11leetBSngbDy9lLBbCc3/KrLAHFn2Ow/qYD+f71
oXYbODIzbRUg3A0co90XqR1RYN3Nyx9Xg3IOuKKuethxM7qFprt9RLO0DpHB
CWwOVxhvQFTGlb3pqzEmCwX8JEYjNShqhxB2LbXE49xTeGMRtn9ka63asXu4
p8Y4aPE0s/pn0m9wPWmkpKwGXzfcYaaXjX4W4P+wixxROGudodiFe92ae+Em
zt5H1P65GBv7X9SmSMhdpaaPHZpK6SvCDBzESMO6+/bYWhuw+bazqvN9nhu4
LaiKQQresfIQpsiCauhmpUUd7AecoGY/00/vkLWTBSBkhP+KL3h5J2/L+MP9
QXAykEV2uh5j/Ui9YjFNSbkVUFqiKtrwqNwFOl50ZG0qWp5lCsbHizDTzyNr
heqUxU7vQiiizUQfDOviYCZH7lFgZn64opjQxABiJPWA2nsXpumavmt4F5kL
912Hp25iD+BMjugHV3RhFAMqI1BXSvFsJ3/S9JuTNDc2JdXi77ZeiXUme1t1
mdmYVVkOgLsrqLWPBgiYdx/uMgcof1sZov90cZTr1v6rcZARwG9mdGZWmqly
mWK3XNu2K6ZJTWlfdMgcoA/5lDODi7bYJpXLi5U41bPcPEOu77CaFUt6Buiw
gfK/74v8jVijppEJLAZ7ddHzJnR9SuLGn5Sg3NfY62oo0fOw2opciwr5YWj0
Bp6qAuOnDei0UZyCNNhTKuvQcig3Otg8WnbuDqIQArsWxIhdGFH99AiY04rz
zD7eVi4nNDRNGyn0aHG/XrVSCqXT3k9gaMezVjp9A9wgA+aAep+O7OhbaEGF
uDLKao+UNJHZUAwQLeg4VPsV2yLrZCVbgFe/5mWorN07d3TLYuSPlOhvCW1N
h10o05lWMgK5GCl+NDlUPHxarnqH3tR/tM7joib+sZ0HX/lJ4ZIWbVAnMChp
a+RF0Tuqs//LLkhqGcb29piy8hppQkbqWrDPvJYWCPBVzjchKBO3QDYSie3i
0YcH0Fo65ux8cOc0u96Iqy9DmqCkGhtbQjYUer6VquLEEx0+tRJq+tAryzfB
7Di3peeWF3dRCtkYbYtmrKHUnTSe4pwhsCuirlY+BrgTYkdHXnbjtI4P4trc
+B39YsfLRp2iJn1pK1WYWwMHy2p3K4WiOI1izHWw8Nz8AnvQvtD4+s7jOp5s
9BKs9RTPkilFBVdCILfMC8uELq+hNjkkwiNBmbw1y81C9iUR410hPoFYo7te
o8CRo5VsmzhSYOIXm5bFMrVNpKRVdttWZdSlwR1E4wOqkFZjORhOrWOdgBSA
xyiLDBj86l1DJJann+LgeVrjpxPhUb0JVgglHbGylKghQrYuKl7snn5f8Jho
BAQrJA21I4yx6jD49lFizZ7m/nwjyI60hbAwQVNhGMfp+8GJLmUANUuuzwvh
HI2TjzbcWDVDGBKtMMaNWufJv1bWW0qglL1Dfu6fLkfR7oPEnVNDNsWaz3tw
8vu4Y6fFk0SsSTKIlPIPbhI0+jCVDbE15DUy2+Jv+BXxNn6tDigZyrq0X0Kn
b81geGp4oG8KIohFpI3+jx/1zkAzgfnnVa0n0sz5HGFd8ztglgNphoho4KJV
IAIkCAS+b+wBTZdkmZa19QsRSF7Oj2xCsrHn46nepVsWl8QHSYh7dSYT0mrb
FMSClbrvkfEJywqeeBnM3/TWWctbNEUxOYPPhbHDJULJ9tJyG7g0s49WzpKg
5x9aECwPLg1Zn2Q1SMNPZbxexiZrZQfChGJrh1JfBUU/ue8xG8fCKijDoJNn
IyEQ29zbEV8wK2vWFV6bsVOBp1KQ6PRt68puzEt0pjj+kRmCimwLL5HOhrl7
N2qDHyxJrDM9EDIVvc9gw2VJ860tbXdYZQbZAwEU9Hcgv0h+JbLcoZBtfPtd
1B7EwKt4OU3VX34+TpH6DxcIHUojle+P4bBv2839q7ZbgWsmreJgDaqNiqWA
SFIEIqELN7ptA/V9agzmIMbT/EkVJrZwMvo5kkfVaeXfhMNUI6tjPolRS8o5
NIdJihiqMPSqFHc8Hkm7/9XkZdegRvwNKRigBLcUYdnS3/1wG3+YuPs5ieGs
8VgDxgbZf8liyT8+c26BZYHfk1Mx5cuJ88npiecpMPdN3whsaUDowjBqNcBd
GkVUQQZVnWVGkNUeVSSIP9BcW81x8TWYHz8Sfy2H/weZnxUJ+qXGwlHIPdgH
ss2+jt3CkkiGL/tciaUTdThrZgDnZdYtZqLHW9cx+1PJ72PaGgLIuqpDneF+
Vxr60gGJvePOvlMO0/mTowjZjqe4awB912RkpZg8Fx2ZdLLoO5Nbn5m90Kyt
RAWd38pUn65LiBX7l90puJe64EHQky2NrX6LgLOr0M4h/thq/+M0007Fk0jq
wkVYT0ohnkicUuBihXunBq72rX0mgvCJR7n6RzNPb2J+pADcr+zN78JWO/qI
Hfk6q655oeTu6FetXCHpGBN5+Gx0MueZ/1AuFqZpYPi6dNvZ3vQGirD8VMuS
zgsIeD52vGXyRfBia4CbPFC9TJH0vW62vLT0bmdRvoFm8Ixs4JgpB+GNmwhP
TvJWOHMdnRAV+tlEZMJioabS1jtwFBwiPE1NZhw27LI4fCTVSRBMW8SbmyJJ
FZFOIivxg2Kvb8AbK/6xQA565LHYZSapmnGsFBnO2zg8Bo7FLm+H7LS3JAgn
4G388qSfeNaqyobtUhcKG1HSRV8B7/T4UDISQguwTB6DpzdL6J71yejFEc/a
3RdfC35v9ypTzT8Y7pIm93MnHVcahpHUPNiJoh517DhnUPbrc5DVGxCQfBTs
aXoDNKdEcvxTvjtxcO2bVVpW+PehfR4otXjO0I32cdUJ86eq5vtFlGJofTKU
mDtqsbSSsH/23yUrV7GpPW6vC+LP3bp1NVNXrgxoOxG8Er1kTclRY8UZmici
ZB4pKnfAQfcllRKJEKZ0lEl5Q2gWpWbkAwKskrjA18lVTwCWAVxB9ESn/IoB
VIhyespeGYtPeTMPLfZ++RG85DGn4Or1K6mub58fZIQEO9CjX7JIqfru7kXb
qV8vj4duRUOMZc3lU6qXApvs9Xkz4+8K6wPe8nahjtXzEvWcRtdBMiYQv9hX
jb5ial7UxoGmLcvD491xjJuqijrunXZwRcBqIyyz5UYskCHh8BPmkDHEqoJ7
OeqT9v1GxWKFQbKS2VY2PA6qXCpWZ7DXOCFCTffjTuvykWj0xs8+eyJ+Qd4p
2WSP37oELXFlg21QwLlu4G9+76XbotRjtPliY0wudKcMVxFQ4mKk2ksTHyCp
j/dutOJJikwUdmcbtg0B3bCxs6iA8CKs82fty0BZkUB62fqmm2nFcum4XMkS
cWOPuUdf4iUw3nw1b02P0K0Oc/bnLXKElZehTngPIACBlkf/ytgFlaHPpE51
JURMbMa8VdGozqHD/8LBU+KkaNr/d35RIhEHJZ1BJZepdPh87J4waz2umlMX
lUtshgboJb3/AWcBydkxfvsf8rZ+ub1AXRG7PeHGFxncZxZ/K1L7aThGgYYl
Qth71Wzm0Dy6/GbqakUoSHB8aMIT2FXK73CaFhblXoP2sgxvPnPA95z2ewJi
pU9ox3FqX7VrKiQJrgK9WEeJjqBuL61hfG0TxU4x8ZwIrCq7OSJvap0n7fo4
2BoewM7rsoeQCyPFqA8hXLqTcdzsoD6s5rrXtCM2quGoACzHIN4HJSbXJTBP
gcl4J/xr+8Xzs5zjrXawS2p3pHXkQ6bUULLZQ7kLR+IjB2nJKNrxBJp0PvdK
np0dh8HWjBxRWOxlJhsByZuh8OdXO9SjTXNNPkYPEMF9JTaEmOasKJcBC3oA
KlWRVJPiSXdVVnjVTxImhs1YD7hqTFShpuMOLLFRBb+hRwmGOuO043wR191R
ZAKFMJrdg5qa7xKctzVsgQjHJNBayH0qreY/9dcA+IoIfiHRfdBz1K7QxXKN
+451xeoLR+Z2k1eJWofkd47+v9TE4kTGZeSWqAeJiKidfoxC1Ejf7zC7vsE/
wzXkJmgjmH8wuwmIasUEqeWc9RKCGQfVHfV5Lm1QlKXjfFijoVMe5ZC8DhdR
kRmMmf3Cxr06nTGn6d6OXjUC1O/p0/RbV28vTxP+qXkU4BPJaOGe1k/pQEe3
v1Iwb3g840eZjbV4i+onlficFQZBfdl6He0VZWHHno0Mgt7UpaHRsj6EOV5y
/5bu9nukj2qHyI4kdStAagqY9RwsRF+SdzAZylP3rzZWIrREMOrBZPtrowGL
Ad74uFOEpU9GmVZUuNA8vFl2rFzQy4Ss3MSIRuIIIOYgReKN10WHxKtw0/N+
B6cfA+eFdcc2ZqMjEawxo17S9JgzjAyAu+aJ0NpXk58IesrLAFC4wKErJlym
w32m/C1s/KgmD+uQVZIIrmuhmn0pKG0w9t+mFU3wcQEoKf0SMkZth6Z/VIBg
EAZU6t/+yt++MFsKT+QSdPVfAGWdB9IO+W3bPtlt9eewhnVFYqcaAlLNQQdg
n2hCA5xU5IgZFXrlDdRlzW6R684y6ucGT+DY/yGEOIkNswS8HzEWk7FhGp8f
/4OUrxgyx+4DguC3imKpsLBJD01w8LeOkLY61Isf/hASDGrDrl304TDGDQcp
svO/dDp6buhmixmSukLAQeCnNGdfPtGqaVtnUw5sKCm2Jyhs3nfeXG6HDD1h
odqI729iJe3R2EfeMThScp9w04QJMuLqgrVMhW+UBPwHSNRXin91EiBd9p0+
mnBYpsOfvV0CMLW0k4TmSfJW0Cry8VGurHzuhSfMnYgPBxWne20IGFrkflU3
d+zE53f38zpL0hX3VWl2Yatkt/oKJg66Y9ABSd38kuEq0KCPmX4L8ksplYis
fuDZvMW0hBjc7rDjT5TLKBGONqAQ6j0zPe13mHdOKBG3qajzfI+bKUcFxg0W
GQh40+5fQ2HHA8eWc3DLklWS0QG6Oj8u7XhXc4BwnB0VHUZKv0a/BqAr3P7p
vxVCz6BOogpRKeONbRt082JVKOCPhRWemiPNCT3QewUxs4tCXGkluZkL1tYQ
igyX5KHtwKDgTdCi62IrV9vnjirRVBt381Ueyu5753ntdyNdqpKiWqfFUS/R
KfYbUSIB8Y3182phOyI6uJCXTtkrVgDjNn5ZecEXeLvA9ObWOdPYd2oRU3RP
npuogz3v1l6THq7AgLHP/Vt5Ru2kKgFLlfEti+Fb74zDRyGVvL1GuDxoxov8
W69SBgUAsW8BT/sjKl6oGaj/sazcav2+yLWdAIyqMWoQn3x3bRV0ULMS3VxO
SgvdZvtNrj/IFgUImTz/2jHjndb00aptOkaPBi7xbvWPSjcrJ96TYUJOqyFS
tt8Ly4SNGqP47A9BytovS1uWQfzXfVIiQ8vFPwEJ7BtBZfV55iqv8iUPvFQA
o+CZ0j0J38gk3OyfbvMg45bY4MC/f5B/i41PLunBeuTmsvsATjnwX9fPxgKP
uPCHrSSJT8dZP6/8i8TzfJ13ntxqx6pk/LTQ38lYHrxT759VXQFaLs8/ZTji
dgSyRJ/IQ2za2drIaM1KAPqyyDKiLSfvQ0t4VF4LTdNKEFhR/MfXf/h1zUqL
SWrJglaW3TX8cKq8aX8jKzsSm3/4Y8zk8ztBQf33+somIok66uFPYE8KTF5G
LdYc58UxSFcCEByEtqgTN3MPDtObE2spPEIhuLbCfSfodES+iO/Y+ntspY2+
4iCA5JLsGJz6W1pVrz95r18aFavqZa1El971dYcZ8Zv0bGwMj5IMNzoEm2mI
7EumNgl5i/UB6+DThppE404AzOXgXPN4HYQMJjHPMQ+c/vZjsCohckg2TMtX
jAsKx3o37IDgxLHhYR/mNQFanKS+yPKg0vnoUAZ2d3On0pXPz2xNSO4I+BtN
wxa8O2OXhenXD/eYfichFMTJDtaaa7VpqtWt5ZG8AdvDoNtzp8XIWRHBv6xV
UCAuM6TR3SWG0fA5OFktN6CQUvWTWXsAWlh5khnkOTtj7QqrGkaiNAH8y3JF
47F/i7zpINwe3RCqAtphhUHOPFJvoT83iYhp9YY4kmSJndnepJnqAbYP1pBa
T4DqyyaG3sDv0aeO8kwMnF876AfLG7yVinw8Jyawx2u52vJ+hp3XfXVhEkNC
eiALmt+eQZ3JM7wHlXP7zoThhmzEL2dBDzZtv/HfzsArBtRwdRM9Bf4n9rcw
wn9cJfUQ5WSmxGQ+JI79PJQ0bczfrUJWQ0pXrvH1RxmcmGP6rW6G9SYuKbY1
I7NzSTa5ESpkbcjj5Yku1f+jFQ280Cx6yzKPj2ihtdGWveDUd82/On6+k7C4
deSsOB1b0/HnnnjbpzqtjzoTRSfKBbCpkJVm/bJgKI10kfL75W5qi1du0CNB
dTtduzWLW5qe7ba6zdprreaDGChZTjHtDFczvd5pFCwVnUlZn5ns1NOChrhf
qN9o1CDnS+dm5YKub8wkRulaTy+jT9l8v9tZpkU5QfROI+ukoSZEUyUYZY+e
ZdUkBH7Dl4Yeu8gOSNEkJxQQwQ9hhiHcAvjhe6n9WZx4un7vNzqRTM0THnHS
6WH+OS41juTQsYw2uZp//5OPhm49NmKJgnU+g3FxrZSN6FIwvF09ie0ZeC3/
CvAweGl2FMY53Sof2dGpbu38x4I6wB3jMcLMZo/vtzJNmk2v4SAwOCdJKsUW
9U8GN5thL1ITlbD+hJj0XnCdlMs6u2egttxveaY1AvENA5v2svoXOL4o9XPP
RMSYnVgkm9cdm8tg197zdp5B2HLFZs0Pye2bmhfzr0R12RgQIWh6XBUxV/9L
DgaLeVNEFX7aSpAIOqK6CcVtu1T8xJJbZb6ePUHInM5whbya69nKqaRh5QbC
dv0o1lT720jigB0FVLqJn5eZ0MUfcEb7tfMsdFg7V0CbJoC5ifZItDxqs8ey
5BaPcg50CPOQ03eqaWidX6N/6mwuqwk6YnhDNqEvctYRi0A+HCzrz5FKAU75
16AgHbDcB3ZE7Kvzk1jyTleL2ksWZstDE3xZmN6Lw2xHk5/yB1eifUFJXNIT
Z6KtQA8PJ/w3YWVxjHx+XextO1IbiWg0ngsKQkujneuas1KFyoC02341tvxX
ShdZ9hZVZtbpGSeGxDVwvXSeAQjNgtb3iaD06XbewKRcEUlZVsxEQSdraNoA
Bv+UZKg9wUyLifo1hu3s+wW+R+Qwx6PciME6Nj7ndGW3g3B9Hr02x7y9zQwP
19Z+dEcslMCWsVkYYbL8vSMueTL3dwA5Ovu2CPrVyT9Z3wJ4rwEFnsYDWn7R
dHnNfRbOUU0uk35fepjqmR9cjfjjSzUgu5tGANFXXt79T2DNqPYXqrUcH+F3
DyQm1VB2ToD5D7rYoOKg7mJUTzh3d/YOlWb8ywEnn0pNg5DmVViT83Bn8xVg
Ljo6j0WdKgmmc8GzB50XYohwthsoCcmQivRNEef2bFWGPoqqwnbj77QPmEsB
uLC6jq3LWk94wkfdvkvnNoqyZkBNu9VbMMHbNUC1owaXJpkjqfEj+2KDlv7i
iIagIeh0pKtom6iEwcmUk6ugIJdk7hoEWD7hpZIJV4L2rRlMIxHDuRTlbn++
VY+6puyRekWkh4AC+fGK/8uNbkNnpERt9WF42kLMBwIYNyUwj0m9C4EYeOzD
LA+aU55N0ZF7ZOpIRuA7cOSbWwz0ZORd9Rdt0NLu0Hz5DEtjh6UMDfMC4J/O
gqFrxU9W6K7EUfMdgC28Bsr9VGP2iTaO2T+qDHgWysaOV4hPzCL4wlOYCyK0
XK3YCzQFeZT8muB+KYDJleswOR0Uilf3q+/n0Ool2LgspN30gAjU23OK0Os8
5hoqagEpN3JIQlrzB7GfHi3H2dDG98Hozn4l++MuywYR5M2NIzmUetCXm7gL
yUXS22/k/X5L6xVlcuEueOQ09/fq/VOz0rgxT0UOBSpA8prKPyGfpA/JKwHS
9apmwgOMpGH6MfOtpo26I1tl0HU8f+mTTFIXyWHkur689br/GHu/5mYp5+rh
7JVjIrvKqC2E6owQTHCfq4Jvyf0QJ4e3Mbm4L1OjC0tavx7RlxZuoLOb+P3B
TCeAnTciWfrQH8QsWOSlQ8e8MRM5eHFxMRtuqaVygA9UIaXJfqTeKl5oQIRB
keKv19GzCddpsW7icC+GXvw+T6fkkte/YkW0PgUU9B8mETgKE2MUomodURGc
vEGdS8/pye0C6hRRNbFkrNt24p1dgqcX8SwPMKRZlhVlrYo4jPv/W0yZHAEo
JzBYUP11omPhmpK/RjgJ2xp93exgkea02npGZakmXDBtFT9CfYMYzELnpSVJ
ohWF8z9l46ZbkMFIbWGaid0bWBm+5sOnLtNhWpt0uA/JB74pe6qgqhrSzJ16
MgQStlz9Vd6+7vRppg3nNIu+GubCcY1vupxrwOpZiVBkk87GmilPPsiY7Zwx
5oicuEwyXBjX/o+F6XfgcVkYe2S8YGB8A3m2awBYjbkoKKhsQMlJLJNMocVB
NK6ev0GhP2fKH8DIvYvGKBrwXD7QVpsw1j7XTX2/vPzVELke8lCH2+q6zJxX
Ls6jPz7CSUi/52sBmJespa6ZVbi48mNSRdmwzFML5mXLnfjE/7kJRUvOtOVg
inp0fTDNpygrk12Oa7g6Jcm2pPZr/YQRVMzyVbDRYgOLZf6jzdtrjg9Gu6h8
gofGwVd9drYdnr8t5arf/cGs9waVdsBq3C+KeSf5sV+GstFWwuAxOdKtt3k9
UOHpqyZO2AfAIB+ZEHSBDw2p8OO4gDCqqv264II92jmqzTsiuHnE0wGzNXeI
GG0QfU2xmyK4gdqj0oR3iGwkpw5YBFZBtzoVAaytQL+XO2osz19WqzdMaE1U
v6hv4M3U3fqoRU50CXKXE14W5TJhPFP4yqrIJxa/OD6fFjYsyA3q9ezyvGBf
ImT/M0MatkKv9H9i7GQr9lbdVDlYcoRNGz6D2kx9B5XnKcG+0/uzic70OBqs
A9BEAYYLboMqUg2F3/bM9TxL1hA3C/XCaowN4X0EUAE87jgOim4l87ld6cLi
cOmbM/MvhK50zLwtYjzD21sC3dZpDdkunMvHvvNyp5vS8X2OWlAnFXDAef41
Ygsg+5F1EHioZbjBs3PBYBNEFblcJvah8MOcfQ8Yg0IKKllh51aLdmVbQuFI
9CSG9NIDA3RXgXSzlAqUCoRGW+ylAUsaK6v0oSGpK/d9YsFdghJJTbJZ3KLD
WMuz+0Psru/V/5G5Ky8tLZDsiDpLbUq9GkVhGIugRiJWZyDjK1slhNHbYlsf
XC/pdrj9Mlw8x+M+NKVC+ZQTaHESlFM+L76AsfaKEbzh041uVtApFwiHSdGM
HW1/zlVkpZB6Kfw2XVY+jwVVfLBfbfASWhZcMjZc74VQOfjv4qL+rk/9v1O5
/p2yWqbzbJ8HJ+n2XDcuMvTvvD1/JHriuKBTMIrDPtB7OrZGcVwbG91jxYxt
P9COgxOLor9InmjqZA/r5ZJjbFHyI8Zuw0pVq1fjqh2BklUTWIiRqq/XT0P7
SMGOPNsNxV7kMQVkS2FIIQptGlWnjlLlHYpkmKV/zgI7RqPz8btfvcDZQzxp
O6lHfLDHts11vB46rh6Zvx274y7hKL47+8EhrKXWGD3rYxiqw3hOXeR/wNJu
tOW3plHlyW5pC00ph9kf4I1FefwbiXZDdQD/I0A8V8lONTIVGeyIWA5fOnz3
WesToLTG99HSZ1vKnJwmCmkR8oYQTrl367ratE82kaFg2v086v4zpC+9n+Qj
N/et6AiUZ+lx3GGy+wvBHAc46+Jo9HhMKawFRPW5PD8bVwRdV4GMbIJi+tSa
G8/yAXs+kemuDm4pWNUG8UIaoxpUkmeXS4pm7usil0NQUBtG6xPtXsvB20Xu
zgVrKPtEVIZi1Jokhxc3gPnpmjsaa0BUAEVHVvupibgil6CwD5S2J3JBpyeI
EZ/a+U01YwI+onPQf8eOEGrTijHL4Zie0YtyRVopiZeVdFNAMV0uLmTzYToz
VFo33AXUHW3djfyCAVP6kYgEXfKMoEVBSM+byGvo81kGS5RnjaO8FPDOYSY3
yhDG3pupSJ3UPxaR0ZCqba76GbP+irGq9nHw36fXthWffOO2meI1n/2A/VYa
Sx347UmenypANt7yORcXE9Ev6CFWc1lQT/09PFbIps3NDpHPKw9UBc8M6NUd
EgwhyPNRz46HWLqWuuHOoNdX3Tn/mezj1OZI6xw+rHsIWj+0VPJQ415Z+cAp
EbNV1/4nhoh8qSvM4tAYXGmorWeBef/2MM2W2hGK62wmD1yOF8tfEjVRY8+8
3Pq+u0n21LqnHdM6+v43AQJwBB7VXbxCDweakGHT1Esh7QqxMPzeXU59XscL
q7GtmZ01iCrm4icNHnOgqv6KEC8Dnu8zjJ+CX8m4vcVlzu6qgPJb7gMCiVsu
irZOLbaijtmNPuMqAitbHO3C5WSGWBkwxJZPamjfJaDvYmVLsB19BhKZWPXo
3a2AMHLMs+Gs84huMp/jMbtqwyDkONdJr1GVl5QQGntlQTDY2RnH8pY3fZRn
s3kYYkDwOl1ccEoxGUnRW6Rk8EK1qbs0GZ1xwyRwgUofk45tzoUEEynAbxkR
p3cz7G9K5LM+ny47j0GHGD43MKIKnQJFxXxNHu9x9S0OdUQd4Ny+42cht+dk
ESPX+g62OErD8Lqj00P9F4l0FUUYZjxgRy/9I5r/Ul8tInrKOYDIFGMTITe0
u7Unm5r6rndbWtJ1f1pFhbPGum9w7KJ3DZoZck2CR/uG5h1Qcq/q2Ex1vPCM
OvL9sJtj9zArJ4Sq/J3BKSBxRoogzAXZm6Plle2RPLLTtEMsLTyB2tZZAlfy
pz8quO5AUEFOkxmiwT/5kW76NpTUnJ2btm+M48EMsJOiNIIe8Vh2NVszqc9b
tEcSKvGPwFqGsWLdnuvq5CzJeOGlxTHUjp2q8ZurASh/Gj7Z8CYMuZHaAYQk
ncogfwFuZkhe6UYNe3E0fAyzfD7kJOSNLnN8uhhfZdAqrZmGffIiN0tetUsu
YxNTCpKxvtwueDTHsAGWct02CF8NVkXRk+d8Jw2WPE1xtdzQFuxanHC8D8Wy
Eh3s8TfaYyN2wpXqnyfHgvw+xdEPjGH2u6MiSmU8PdVGF1wqNlzkegJhMyoO
iES++tLAGBNzz1iIfULbVT1yMVIsrs4wwo33DwUh8u4QUBnSDvbefdMBucSU
fplw2aPwDbFJPWjFBtBtmRq3PHIkAUrBQrHxbWvzkc5ziYRm6t/7xv3Kd5dZ
+h+2Jje9jXBth6mT89oc7/9shAs30Bj7ngVLSpwLd9rAbKzMiS52wgj7eTyb
mh0aMOPk1+Py4jjJ3gNGN7yF+h3zwzkcYlK6NQCjMaPcadGtt2VsX3wOSUk4
xxQf3SPfyp9oa8NGUJHOcTa9gvjzs5VCaFYGGwxugPEzdSnM61iDhi+oZBpu
JDj7VW0XOkui0XyQ8H9VaG7upokDLKkFwUAFqFhlNHi04KmHLA9kN6vE3Ivp
hI+08ZNFOgITqad7Tge32zCspTiPubrlipleNIraERMW5WZe1MDXjmmkcqHM
mrMNdHccKPJ5s8QY04ARm0dqdAJUPMjEGPQNM76oLYwVY68Cd++IvFcLjVQq
pLjlJ7nD16ITWmDlgQwN53jIKugxd1ion+cWI3rzPkMwnz3MBejzKfKYudjp
N2+3V02HUlUj4E+BHkRIZA7TyqGSyJDa5HGGbPJjN/hw8MgpCgu6lU0xkRTS
M0ZAK+DnKKnXSXUsJXpHGU0aKPlZiL36h+onahyls6p3mNt11RlNTQiCDadH
r8joVra0/e4LYwz1xmaKNHnj25A0GZlWvImFnrhiqTAidsMm5REX41E2CubF
YPIjYMF7w2IArt5Et/722depYKuvspOl116+d3gsLBUchJXk3lEtpgcJ2P+f
qNCDlQ3HCjAU76jfXwQb7YuI1Up0iUi2jGmIV2JDwrqzhT2NLAfbi1UUzzuL
Q1cl12jcZhojK/ifzwnvMm7qnAArwq1BPyYdrd2XgRLNZdTluyqvut3MJvvP
Ze2D4EplzF6oXLzhhYvyWhxTvR9OIPRKKSh/rH/KZZZVuYF0Rb9gYCtVzSRK
fGO/svN1+r/xdpWtMXr8LV8F/FJRjdq+CnD/JEt6i9mSphOUi2apj9QmwXHh
AoG3NojEY+nUgrSyf4kQGF22dOLjInMrvlUB8NhonJ/54vQtG6l/zq0BeYvL
+mdQBSBTJHLr01+exKp29u3ZYK9lJRPKi1T1HjdBlueqlfNZKcFbD+o6azye
SnnhzfXE0i0DcfzMxxsnjfOl6hFwnvWsYbASB9Dq80RTdDQHXJ3CsUgBXwAa
twJZowf6gP/aExJ+fNeKDI2cXUqZth2efXncBuaesg7wYi9qOy9bc3NDwEr2
l8V8K/D87gvjLo+EcgyPd/9O3rLXAD7SZEmbYMslmkoD/X/eOG4FC5koJFEk
LizEXQnjZgz9sloLVGCFwdZGXhgWnHBGYf15e9TNTp1Zr7hjrKILeoHoVMhM
+az+1Qggx8JaAVbZVBM0S/HCQEJma1j2qhig6iLGW9iHFOnYcvYbNLN8QP2Y
aq3p6F8E6MYbQ8Cn7Z+CK5DavaRWeIJGZijbZjIeHTayuJ31UdC4IaLTU/XX
DxZeOIfWJTPHaroo2Gp6PP7dnxdPA1KchyifZFEQi3EZ374Wb747y5rZcmfC
LvCsVZ3Z3ulLKdZhaS3MXWKZa6DRezBSbdcBtbC9Dj399b+eCN7mIfPkSqpG
ssEvLvRQ6kPjEBWuyFU1OpmJyMJoKTjVSsKN4jjZvQNjXOtR3GKrE+D6xbFV
ECUMnDa/tVlYkrRXeYyyfSySKwIP1EdtDGkfFDGlxwPQXcW9yVDb9auHrII0
SfrteuP7W+g6bTmd9ZXhvCSei34vQDBaDi7E8sdNuys6eWOuZRncz0y5Bm2G
cnbcYRrVDOWEjM/5Rit1G9Pil4Aexv+OnUGOulGY2kSeLkOqPOW3Xlx6uSLV
FvLM+J/SBmj+HnLNAxGs46OLK1lF4QooPDGyFuB3dJi4ZJ0xS62eRIM/Rwwn
87/1T7BqtKpY4L4Wz6VpShlKLE23qyrRd1QEx0iuN6ZwE8IWfNGYerk1qTjI
qdRdlwPkkFXVVDF3nDHJb8QRuSHBjUa/rBEx0OJ7lf7GDePoqD25fVeaLuDX
9AOtHwnQccfUehM7Vw4woMLsr1Jg89j3o5TFMS/YL146d/y+ENu7Egcm7k1o
bRQ4SREUU8jfcSjw7/vlSHnzlbCpUdbXoWt4YwmDE8YSJJD65lS4JUHaPKHp
QjKG8Cb3UU2G5N83+nauPb298fVpaKkU6SSZqip6hloL7Kplc3m0DqcldwEU
qWmR0SeP8eXhGu9uzTt77MMOo6owjsaDlBzUE0tuzf2dLeYJJpg7ojqkjgje
YYUy/qAmbdw4oiNP4CXm5nna12uANd4pU5SO1Y+iN+6jtIdd4bWZNkWX2KJi
vHLrVg8Tjwhe4BMLxbJfF+rU7ZqyiZGhXRNxryRBXgJ6CGlxItw3uYu/U/U9
TJ3xMmtU+L/CcBs4fGpCFgDEyO3McFWIup2VBlJHkditc/x+GfeCH8d/ncWD
Sb8fJsZMlFulZLQPsy/rlT0yx+57bebmzgxKETA4irXREwfgepPaMTAToYum
E5izax9q7Rh+KHShuRpcEmzfemY21JCv8TH8ApRL1A8RkBwkz33euUym4Mvc
vo9t+vx35mOu/AoMLfZFlfgmtivUmKAAjg0JXqef34rbRC/nPNOSuAHjTa1O
FvtXzG44Dve5zGzp7l100+gnc9Rgod1KQjEq1pKHeKURWPpyJccXc06E+x4I
rPRVinMwzjUZH0+nAmIZIC3PXVaiuRmTFTA6/BqMvAz5O9bKNhQbudEDFkNp
sdzVWr0qw8DYA4yySulyy7hq84KfmWueQDKBCaNEwZ4RanIG69lmN43xkAgZ
XErLkFydxjmYsQZY0oSd1GVXxwXidtDe7Ig8wqr8cULMpdVTQ+VUT80hmWcH
sDvpvo7rAS60hJ5HOWuUDjkH4kBoz6Q+zi9BslXN7DFhypgST7rkRguFdiRR
oanndCK8fRws8QVe7x8tavrjE7BR5M2pL9Jb4AHUd+LPCTVlNoPUfPeBiPgP
CCW87Rv6RNwCfBWXTI/ljrLvm2rmYL6qqiND/thubBAmtiEnZJhYmsjWNoaJ
tYPtho+URYsDpv9exyErdhdATBP8QX2c7VEoE4KeHBThbtZZRD7Wq7QoesNR
m7e4lOm6t4Y2QJYsSujAcjZcnNJC7VxXr180n58LvjtIE/vSCKZDkdYfv3WG
6Kr2Ye3MMCaEaVnr7HPF5oRCevGxoJY2udoTRdNNPU6m50c/PqVKBucG3mb2
JEKq6klAzU7CYhwX7LHGme837YdKxH/bhW7c5YYcsM7NNaAHAzRbdu3SA6gX
F+SijRjlQWcuCL5UAAe+8qeBZkE59pPpYRy54saT80hFJSrkUUF8T9yc+X/s
Au6Mz13Ep6ajOMFVwciSbfPjC9mi/i3pcU321QhScDKJ+YGywWhKOeJrNBFQ
uxkspeDk8fN1zldonUQHp8as0Wqp63KIRGl4CKmZqy+G2LwA1CI+fsSzp1EW
cTxb4eZgMH+Gt45DEAVDwoUJUewKvIR3WCmXSmfdFUPy11quYwlugxsmbHZQ
VAoyv+YFf5sBC9U5J9cC66CxSMGHZYUHdC1IOS8Onohcn2zbf2LhzP9FN0E0
TCSx1ylvpSRp6CvRa2kNXP9fxIK85Oc+KOMPDuGZix4Qx3Tn/eCpKLH7d8KO
q80znhshH5aoe5EvgdBAr8JBe4Be81IclxqFWvWsfEaIGcOOVmMWU0pxIfYV
QEnJVYxnu1vYAoa5w4ofYqiQrcPUgK/OtAxp3UBHh1MXV9yJrfDnpdbo0yzw
CXe8U8evLpC5mDj/miAKaWbhT7/U+n2PdCM2T0c7QxdPMWQ75bv4iyDTJgsF
Hq8S3xsXcCZ6MpcaJmElKXDGMi1MVkYW86KfEYI1ylRcn3W6mmtbbL5qvC2a
1wNVridscUTALpx5SiAgpF7vLUOvkjT7h5zLAyLWbnBWVRb2YHkfAJt27Aq3
UxEdyE7m4ohzqR4LncBcNG0WKEHGNsSYmSz5ZpwIX304WcC8BGYFrwB1iBjs
v8RUIMtLyKYw2V40yP+im8U8/fezQ2I8AYrLaVcZul337rcGQ6g388gZMiuq
3iapVyO4TKumE9sIPB2X90wpUkoO+xY+8D/FpoB5xsA/jH/3tg6iH3jobOxq
KvUzg/KrxcVOt+sAfuCGtJAubuoE6qStsdYTVVTl89mmUlB5mAxnQTSYCACo
IiH/KtnbsbSCfWEysp/xJwLfSQwlNrCq8PfbxQKFY8Or5Qz6XY9K9k80QY2L
lUIL9taNxirbDW6/dux0WbdAGIFZhsT+wiGfrqjInsdAIPxO7kNOfqdRR+ZC
0wKww1kL5EtHBLhBToEoJhBXWpOXAKuJ01GNbqjrDWYGBs0gGNvkVeHCrJ7x
IE2pTxiVmfaS8Q12pGK6X4++XvvtMr83UAFrN7akgaRXI83br2OBCfLnxJxG
k3rlSaqs80lQSXMAszLpDmj8v0ANsuRWUD9gbiGYPt56thuhIEc13bB94DIe
qpNTWSrE2KOwDBdCJFpB6Pdj3najprPuuBPKLf2EuBE35GGQE/lRlVpUoKdF
oSl4ebSSpnsySwp+y4ApVTq0poqzjw8S8Lg75AoB7Rbm4Hel0SfWH+pQQsHO
FIKKaniWB1pI6nubwDK97fqjXnqiiJvAkcpvqhM/YkgSx8gQLeX98pwmMpLj
FpP+hYgsU4GgRmhvDLGJS9DvfcGU9Ylb68wBGSbYmsAKTuUCxorDYVRYzf3U
cw+A3T/J3x7uU2xx/1NvcvPesL3GP1TkOo+rxLZeoXc+0l5rERaXHoZ+FQU2
lqbyDaKoeKQfz5zdCF//zWB+IwIMhnBVmdv9E6bjaY9mX0yZPB51IEGFEFZs
cfZcbwFm/xJCFUSkGKJUyyiAWu9nD+P74Q4drs9V+vjQYD78FZLDrkrND0TT
wxt/dQvC82E6oPlDdzQHDE/XamXwGMnl++xo2Pnc1OxUP2YUbHfFW+qgJzwH
cYdZTuetjjD93qy6xGbIEFVCH4jD3cgySbGZ0TJto6cATAz0h+OrVQkGH0C4
rY8bLaAmXbIfhsX4RByE9NcupquJWd5/UhZl86RIReJUbMx7i+xjNxAw/2Dx
qaRTAqSgssHJ3ws/xzrLbl5LwQ/8C/zhamFbbX0Mt6f++05s9+ZV7W46ALZA
9BArSpCn3MqKtCf8A7TYgIe6nboLHcwazxEm3c6fD0bJZUfTNtLbNldEIUyf
47F+y/epb9RD9smXyUgcaSfLaoxb7zq7AA5+ptKxleXQv6dZRglaNK7oXp7Y
CwdjNbj3P7PitYHEYS2zn7qHgQCY/6LgzDcXBYBGCFMdlTmgx6X5g2N3EbZu
rxkNHGlqs6EY2nIjRtbw2PbewoY8TAl4xPLMiU6Si4qPqWDWcDyxIC4ZvqLA
w1fiTdqN+JyROz1d8qFeaPHbqsbwisjZvdzyoHtIN2o1ppYLhPxa1LpJCZVw
TkUL0p+41G4A9w8KFDcg/xRsehuAa6E/zCv7HY3PcodN1f8yk78dFgRUx4c7
xg/UxJybbKqCHZmNpgBw9LfYVRcgRp0govn49LFO7r6fSuSfXLpONXUXkNWR
1slQz7uu5UthsQg5ESzqWHqu2EZawm37zMf1fnlPhlyXqgTQi6B7OyHyM/42
oROhH64uWXldrl8go4zPrMdUYIqJScPhRTBSQDepEgLdogfMSiuOyg5P5MPM
4SLckqefdeLb2gfi35jTew+kxR0PCaNkoTCYTCtg8LbEln5eK8IWgu1/t/7B
XOOKGrE4GQFx3rE1Og4QIhNKRmTeGb/Fb2He2OVv387PWq6Vhp2IdP9HmOkp
Jjf1Om3uTdCxvV5CTCNhWs8jOXNHh1A/BU50pLkNnrfF2+IY0I2rrQdrR05t
+9OWjwxSA1neshViBr/AdbTax6d3BcU5/FZ4kb+S0P7HtSgr5THdnUEN6ThA
1kQ8QjJiEoQJ1+qxa76AzRAJIu+WsusRFOislHY+Uig8ikzRIkeyGXn/VOD/
70mjkpAzDDy380KvRMLaI2bKeo/M+Bt50lQ5om5D086mlsDK/dVxjkxbD2rl
+hWBDqQXq+MOGk0K89upnLpcIxI2w4r+E4HVi1/whZyAjkBXQwpzhaWM3TGH
md7/AagKnitAI3K9CMf4CY2nCu/Aku0XtNLbVOvwv8RaWQKYd0jSPpfunSzL
yi0okEbR7lcRwG3Wfb1d1+oZoM9eNlU0uRFB0Ae+uABAyM2YUjKkvUCzjZZ7
Zup5Bd53HsVYDBXQjHXBZkZetkoa9gRx5tVqEg382SDnl7VDqHmrFO/OeHRJ
WKv/k3iUfInF7asNVd2t5rR9nNqqCgthKh2CwfbWDk8mW5uIKhHNOnZk/ktJ
UyhS5OFBfO5rTFF4VQpjn4ObmKqPp8QeT7pHVDiI5e6T+/PTL0xodQSz36zC
NsO9UeeDyvYbsSuCXqKIVWuB2LcMZvdmN/MrxktN8UdmiuGy4DTei/+ES14n
1G+tVKyWO7qcOj42zzkRWSDh3ILhoDezTWrRjYuy35tg7zCYNy2BIfq5tHi0
V9jDro1WjVYHCFRyPL2WgG1XPS5Py9jVDWs9+snfeMThsJpADmBJRsiqOG5J
oLtq5hnfEoU8yqEU04U8QPavPfYhw3VliFOpxLjyKHcJDAy1kOFy1i9NV3sR
SFtNv/4I81ZhBlMEFodRciwxPmCh5bzZ6/8kUkQP2+efzApkCd9Y3Mp37Z6i
JGY7dN2v7vOMYWV2SKsZjtmU9oD3t+Y3RRjA4pbXlc8s+T4BimkrcScfDRhu
sK6efIezIQeQWJQsJdapgefc4FL+zlWhs9G9VTFJ/tCR1MqMKPv7XCCoRk13
QTR+vdpwgYh3zwUm1Q971EVcwo14dP7ScrigOW+Ntw4zDWNADphqvP56KYw9
rucd6jSbZloTQQrXzaYR49QgaQ+L94jTTCvcYBwTcFNEQK90JaF1Phlc5AKB
SLPhZhC26FNWGSh6bP+7aGlHy6kSiUfhcHTts2pfdPQl4WKlyXFehKaxUk+j
ReBz6zrfz+XKsFJF4rCOnMZd1qMWWghNBS3zntafjL1gHkITr6VR4Rcdk7u4
ghEXY4kMcvxRIDO/aad92TFOL9vrWAjqkIqBaKqwF7G6hFSLhqw/2xf6fLHw
UfMEbbfZD4xljVj/uJSkOTtZTg9UwAtNyXO/ZmgbICn4y8J9V/MPkvXqcy7w
6YqcpwuO4zVn7/dxnJYEh+Mvk2AF8VtMDPDg2j+hzOQjJJ3c63LTFazEyjfd
rYIg4wlJp4A4foIsoLxvGsk1fALVd+vu9CrCfvZC5v3Y7BTned8SGBNPkb2r
gn/lEYS/5SDEfqLA0aGBEtqSZa6cucnWSguOJWRdyrxL3dBdE7yG2H6HPUjy
3VGY8ykwZciWhTbLAGWKAXBYQvaD6eyVUPc64vnj42KYmglUEJ2CaqPDn8HW
FWShAF0oLerA3jTV8i68a5soSaub7ObNl/yA7bGQgYBEq6sQ4EL9ec38XH9Q
46h8VbU6pBXFF4/+lPnC4fDUy/WgvFcgU4YJRq4v/pE1mzwsTC1l+YF5uUI8
RTRn4wzOd61gW9LqHx+eHAxI7YerhGQHSXC6jZjW06G85v8xtsGDt6svN9dh
YPr3M0w1ShcdwKrtr/bPcPKD7yG4c1p+AamGEIF+QUgWHlj7jpj7O9bctzOT
WVWKq8LZjFYFPijGg4yfciFWlaol5Rkb2FOaRvVa2ePzeKrBd8obLe8njJcK
NEGWAwAR5m1fIfGywRBADak/KbvKyOTv41EQCY+RZosnWqBvpTTIRJyXNc9f
S0ljObU9RMRxUdqFmmQwMl4gPKXWSV7iHB0MhhtKer/cVWwv9KGPIzRQxOn3
Y33pwfYRitPrg7ofBZ2vxwakiHdL5icmI9VNK41Hps+5eQ3LW3i/i5nrylzc
fkHo4fqbFHidyxPJDdGtiTMdxHENZineiMDkN+XX10hvDVXBKocW4J1DtcNM
u3l4PuPnOreysxmQJnHpLuJ+bASj9sJZE1GasRju/suStVOH6p3Q9A9bVEy8
jhItdJFbYoUWPF3ZxwB93lmh7YIaplrQrYTQOsOILfGo9QLJPszRZM9ZpKIT
H+gQ+BIxLcy9X1JUTO1vFOCGSJPpbGrRyeRJNMA0X++taaQY3EPUImF9PLyg
QwSmez3aIRERNzR6ZLa4VWHapmSTX4WD6HlwxPCmgZxq2DTt2/67k06xZkXV
7aJ3zde4baIhUjjdI3yfkUOozcMSyyP432YhsIYqKOz7fQSLM5RiZvjXR0sn
OHXOhxJAFE+F09ircLmxb/QjuByTRCUAHak6EpSL4TJSnZmfdt7UHD3eILA+
3T918hr/hFQHJyGLTZ+phPxdwkCKZRESFeqwHQT0sFQEwyWqitTON0PV/LNX
DiKn11bcvaWgoWL0WEVGd1YGHVQcj3Y7XfJYtwHS6qfX8iNCAYppyAJm/K4Y
a6abmkBYGSfgTFpWWvhNlVRn/914a4M3HTfNZv+49d23A5J2iJD4ySG6bcdo
BXBmHJYNwEn2gyKgmBJmrwv7DM5S7Z1/bYpJihv2MT6/Iw1C8NO/fm/rRSB4
X7mAN3NI+eb4MEjhY+srejEQCvPj7zcx1+K01kWEp8CEk5/4GuqP0DXFanjH
za8kE6IHvh2pCTuPUc8GYEWWwf9Rij4fr7K+1c4wZ4785f8+3xbKOkTVkPHQ
GrzWnj+z8qdrWUe4uy22+7N/OvOCaoqqO+AeUm5f3KT6QLCxnJ3jRT2WJny0
ZZWQmjeVjKG9uBhVvy1iIS5zfNH6ZAx47pRZM657JcEG9RMHZqO5amv0e7iP
Ay3cHybfP87HtC5MMgnM9WonO8nevO+y3nZxUtGbXaWW2IKKzdC1LWqE1/Vg
qFqz174oLPMBHgiQq3YzBGm8+tv85JHg1q4YwGm686XKpn6/CZWn47X6SJUB
idLpdBLo+kaWIswDjGvTI0MbpxC/Vzy8O00j+Vt+Jz6HMKqOUMH4/L1j+ud+
cwvvDQy97Hh7XWiwhpYn3z4CJP+npnL57dp8JMcFDeqYtzJT+mfV8DuXkF6U
KA7NiH3FSfY7Dpmoo9u04cnyXhBraaG0uKkriJjFVEPiUdafe0fEzJmffWOb
iVVTwlay0Iq3PlL69hIeuVaNHtZAQ8c+TFvHFVAio3iFnb5G3/ElQwz6COah
PmlhsM3p0iK1pIYXEIzGgtvN1h219vrbQIqikNkEow86DswbYAmEV2D+QZlV
TeXf9ZX/jiIAdw/iGYqXdttghPCl+3RmRHF6k/+RzRsBjbaXxRqxOPyKvAW0
u6A2ZaCqNWDJqH3YuAMMGD7Ye8ZkNJNfKdxW3R37tzVBlq3tS5Ga5o+Rk+mn
d33c3V4lClI+9S96Vb8jkLa55xlEGzKL6XzYeBUFIHwU/uqVwzUKWu/kSQP5
NF6XebFzkKjTnDIGAiFjiRF5hidaFpYGVjksc0QSshJ9SLpA4Q3AmCYRDaZr
btrB5Lx7a85NRQJLT0dZXhNvg2KCx10nkK+JNlZlHyzTgoWjZNZcuCVRnG3E
PqBTci9qAk6VbwP3rgmCw28SqkMTfgmc6wAHk3HDlNirV5HBYW1HC3vIm6u3
5npobxuoqPqcrei8bI3qWLz2/kZIli0Bija91sCPeXEr05NytEl+zKwOvYDo
2iXP7h8j9DmIBJ6Ulq/ApaouIu4U2wV1ir24bTqwJA8sjctyg9ALSakhLlKb
ZWfZy+nEmFrAONYEWEm390Jct65YWDFtHRxcst855W3Gdv+tBs3Zsc2IhQZY
xxcbb9DksUz0ZHeag7xsBoWRKZLSKOmslwEyOLhDJ06T3VvAK1nzwwj7+aZl
x8fvew/wNJamM2HE7UHQBgS0Ud9FPzQcA2MpIcvpIoI5/rEjeSIvva8nM2Gt
FVZdLAuP8USiAjCo3E1J8gUsy7rNqhMmD5G+scsNR0V/ScGfAlf4PHWODkxt
k0OnLuepQNih6TPty2bfG91FqXRDx0ctrv9gqnRGoMtGsGc8tkU1jzq6lEpK
361adn9Q4Y4RF48Upkf84/I3bnWm2S/eHA9e5qMBtamFgI1R3UTNKfVebsa9
ZEvKNOq+LUK7bHjJIJaYouin1LOmhY44n4O8Gd6lyAR/QmNH0ljJuCuGztCC
OESyUQ4nNkBSlWeEgTZHM4XU8ztb9dY2SjyOIn/pW0/y8kPG9ZA6NpCqvLUG
tGYF9zpPWoH4XxdOL1SL9Vvg2Fs/iPKY+SbIT1rHjlRb6QZxbTLk1Mly20fl
bE8PnmTygl3L3es5TFOlO0vNrB5WreSU8yXMypMkE2pTTFPmzYJjLwbjQihx
IA9wzn93xg9KXl27pJ0keWsSDBvg08pLQVt4NL0mBpT3iCNRK0SMEQQcB4z+
JyvGzeFc34SQO/dzHaxPWN/UqhG/RQoM50XDfy579doRoAfFC6dAX4TwCdvA
JoiujOZXUr0XAsR69OkQXUWWO9MkMLprtTh35URDqLw6u9ZsO+v/Kopf9O3z
lHnRir8u2v6Bvls79yFZtgecNH+66gra8yMZf0YrApwm2/hQISHI4AalYvci
AfxPKnHwzk5wmdZw17zzZ49qV5BzvKnvGbSziF+c9qKPe9HVybp8bVyCg7wh
9HDF4QVv1TuJ84PznkRnvWgK0ceKvlXyeeRC03G8fYqZEq2g0XYGO4QamJwi
9bTwmoqSIZWop0idujTd8glDIGg91xsOzYlsaZD7alSi3/Tq4ajAe/KixNPm
EhlpmGV7FxWaUgDF36osbrOR4kFervVmfQnka0UKAM5hAHNO2KX5I/MEiVh6
7m8d9biEo+4scGT3zDPnN2xMHMmhP4zOA2xNXdxVit6fW35jvPJh77kjTb97
LJJYsAOaoYbpWwpDX0oaqTqgYY7D9jj2t8gUUB3iuUW9l9E6XoHbzcW1dMeW
BLdnw6LYNvkmTVyvu677dnFZvuZLyLSBgWcdOabSt8Fqgsko5JRrd61UYHrx
ECzTQiaeiKsML5/i6pwWeWO27PbgnsShsTj+33R30ABY0hESEcOzmDYnYrW3
4WqN9ex+idU4HwH4sMCvVi5v3z/b2ol7rcFDo53XbCT1GnPqdDmAG1cG8ZzA
m5Sv2HBDBr3LgD4o4SQwr9daS+PiErCQ6TlHheNCTF1ROImN5n/DTYc7gbRS
oFfn4yMy8e+tL9rNM8FI1jym20R3RpvimvV4OvcvIfKuKG1wZreyj+bff8dn
xT0/fibv4iN9GmGyLCC1n++CH1MaOPyYWE9INgczIVFVfRrUQxR6ZkoWFoRK
ZqfYB1ub0Ro8LvJRTmsUQfa3ErcH1b5Sfi01rzEQuHlPW3wlqLRkCF3lZQue
OV0HWeMpe5AXp+8n6V7GpDxGi53HtvjgGjRXyex0T4wGoP+hYNcDR8Paf7Pa
sPfimPhxnaU7kml/QFLnBjrhQME2vQ6PoVlEwA5WIyoB92eQXiLw1miI068a
K+gg1ksa5SCly0WQc6H7P47p/JDL85EnYCLLln7l/RTJAkvRC1BwQUI/2SGA
9sJw04WOpJlDkHG2BYBXMqbFVbSBOEyxb7u/WIxdEWJkmXWGDXbS6N8uwsPa
L6L/OLsTCiXCiHnHG8D9yJuObNv8ENAferty1iRH/fr0tsOwG3RWaVZVmU0M
ehGCOOWI+QI1pBsRM4kkhMSw3vDIF8ij6vtOygn3w7+Zj3aXkEyKZByzuV2l
PB8h3ImifSAUryM2p0AwTzH78kglSGZQUill+CqsR8H9NHXH4FH55BIDIXOB
FSxwhwFLCQQZSWm75bjJ/7zivwK4BQHwE3uJ8ssw5fnPgdO59e3LIkirdY86
JHPSr3iv1lhmnvHxpY0Paxhrr9GWfYlV7CKClZs/y/5Owa6d9R6EKqRzpJgV
KUQvPA+xytoyu24Dm7NJmuRmP+NS8eohRWCqqpXadeK+BffIa8uIajZ6/T1G
fLHV7bIvAlN4c6npy1rcRmPhAa2vhWeILBPiNRaCjxrWE52wpt7fUJElFvP4
kSzKa+SYU1I5+7GWou1XcSSbFVAk95bOzzIiWzIUtHJ5Cp21N9fe6UcI9ScD
TFTX2fbPzVSYwwfO0x/XxmPwZiuWgnq2xwTNfFBl23QplBWf319eQE8gYUrS
ned9G5C6DyjCcIIaen+yiX1ITpEo3grIO5awl2q+SCalDr9x15ABo6jw3VxP
YM2kFrwMJPQ4K39NWz4lS0X+3rS/DI6J/hsvct4tuJr9IZ+BXcjeFO1pGNAs
zkKh7iDAjnyWesz6Wi9J/QQIqf0hG9BvroS7sJux3NlxEqN75UE73JB0Gk5k
jFB+rx3qz6BnVhBMrGs0+nX3iDoXA7uUb3IBYTokZQaU3CVC6aKLj3D6hf3J
ai7NDYiXeChEctbvR9Y6jkgICClakDaYFyz70BJ2m5R65T1rDGH4Fs7NCVeH
W1lQvVdO8PXu9aw7p7VYDTzkpSsW2isP4z7sur4A2ZRtWNU25NQI0BcvbPJG
K6Xxwc2sb8Vb/3jEamaIZwallJXu19gNAr68hG3s7V8UNfAJ9NdUG1BYZ9Qr
8iXJv211WmgqU8wktwyuh75yR+W0LI95u39nDxZbxbFpzpUPVc7WJbg5pr6D
tiJ43DZ3zGDjuMEf0Wdi94B3c2ZK5QAaudSfY9ZrbqNRURsfk5Lf7+J6Z33x
ZzJgkTNvPXnGnOh99j9J5tLRyw5xRjsE0C6WW0FusR67Q0HMqNJQvCu9fm+G
MkHtN2UU4vUc6LLUg2bS1nYzLpaFCEuw/oFN50l2o2uYCQffNmUOupI4y7rn
KM8GaUPm3R4sedHil6bWvWlqsp7ZzPH1kR5JHLC/WtEpl1pLGlYvFVxJZ3qO
ZWZsWG5zGmQht9IenT4+wcLT02VzXp/vJBxM9hf1K9PsLzTghrx+OdqpGLVz
Ul/LYSrAWU2OuTk+2jHPpvy6kd9UVqbO0yMh3p7MogLI63pLchxVWQmQ6XjT
6yIUlfiUNhqPf6+vtRh5ULuhrDgiQyRzuUIAmcqpOZ0GQFh7IpACriyiOeWH
hCFbeL+hlVRn5Ql8SlJV5oKbeAEWk7T6VSP2PvDH+BtGLHC9Rxsh743a6Joa
EomnsZaGqaGlWm21w5of8syA35+695xQdJcBw0rfWCurG/1c15EGsWZqDKG/
SIqlpaSEWyAZxuOzjjygOnmEP6cPKs7EM0iqBptCra7Fli/9Ta4doTsVgTx8
6/1dOLvaZYo3hPfA8XKi+HakDnaR5LUL1iAl/uGR35DabfST/QztRQ3/3n5r
lIkaEW6Q+5TX7AFXZGCNPD8azq+Jk0jUDz1gjjqqWksNsuk/DRJZ3e6WLxgs
YdBheIxKA+ImTLMxZ7Ik5aCDetfOXZMNWnIb70PiDVeZUlXI5oQRmJ16JKBS
DOFl5F4ccuRFxg5j+DUZn6bFTKOwI7tBCfd2+XOne0Se4HebN79xs9up9RG/
3uAeHIT7rFBdDbqMWmqAdaPuwI2SaJqNHKzInSbqDnqVnthdmMazFR/G3dJu
6gxSXdPMxaCoHv1DgZq2salSMK7GYF5pHow8ragbC2opdbKHd8e7u4g4KfaQ
KYa63FSiyCvTny0Q4hGen4JeBOnAmVJn/Jpym+5UHjjC2JscikJT7NoC6O0w
Zy6vb9hCxlvh2vykbQq8QUx6YKFSwi0WQRJk9K+/yYWg3R7HstzSo4xQWX/V
96ik/QM4DtJmN5jVq7udDCo76W1Uu3z98qnus4rU4TZsaF3unkSJzuoMxp8l
aOOEMmWNwUUr0zlIYnkhnad2ORgIC4xzZXLNVYouh26cTCkzV43gM5dx2cGn
/T33jnkOuxii/DYXSZ2q7zKW6YzrVFt7iwirsIOvjJ0/DHvwryoaLFxnkOYx
PTq80pcVCSsKAM0U6U3gpsPhLvOEEsmarouZexY04sEkQUQwUiZhZa30nBNH
j3HzsC7s0I9Ap2daI6kGhueTb3RQBRVbbCwO0Siixwv1FmDYwBgVbkQCCYvp
Vd+GM0Xujca3HkATVf+6VTiqMJSKXqSUJK0ZC2CD98W+TflfhRc6A8QZiii2
oAJX76vYtFg+7pHhNojEutJVf4h5fdsflrWSotitc0MOPQR5Edj53trEfNyX
v/AMXYwo4KXos2qFYQtVYvhdU/eXmZQrTc8uw90guvpMmEiw+tVQeP398sY/
FJvZ5B384/PYE7+XfG//V35KVEA+tcCF8bYIMR3uYWzioe0s/M7XftOkRPUb
rNJC/EN4EeCjikeOxVP1c/CWlVzaOYqMEueI8TxBOjt1Pc9/3k+3SFI6P2AS
89g6ldz39uiQykLTaqS0d38uHpNoMaGe03auPmnktQtMbnkwSBAnKE7YD8WN
GZbpUcWT5O8Z0d0WNJLh/yARCwfGdA+3uyPXUhvzb/bvXCcS1pseWXi5FISM
uDhc7gInjP4ioqHODEDivWZGncAuLeoOaSmc7LJdgB9QEcmH9MI82yjJNXfe
p7czApMbeecxajstx2yIaHpK8pZ/D0mmiULATUqpYpMx0cmqLUtpAenfZwQM
cR6lIWz6tdpbezXJ2vc3ajGaYWh8qOsM4/acmCaYNXTgBWE+LZUOQydTvbC0
wS/aa2G6/xIL3RKD2hx6qxfN2kmVOJgWz+AdUAgr2bsesXkLm9Nokli5T50m
VAai/crmJ2ogIFH4kAJzmFOVqE6CQUv8rO3MDKBzy18BHp4/jlaXKJH2vPf6
tev2m4n7+E5lhPB/t3DECVeJe6i5lZC67ZrOcupCJOe3zXpyuocfZw71D4Hs
ADag3YJBOqorFAWre5LHCl/yBAUA2+cOqivtODewqaEHYCM03yCY5DmIZQCg
ZOTgZL8nNz+JtNs0BpGcuq0sy9q0BaLS2iLOtSagqJoHnRAZwZ/ss82JJSSP
spgBqaycxFneF8PShIcaabit2+rKbqJGX5rQWK5juOWKk45g32VgmdCv6WWz
gC+186VKHRRxZBf18V3nm5y7xn8XrMd7rUBsmtWMTRP/pYuHgCGF3h2QMzmW
JY7wtybPofdf7HFpmr5qvVbJOXzNOxL26Et7c/9qtFuZTjnHXe08+cj8ujYS
nGAtaFN6heUA9Hv210eAyZpt8O8n+YqdnYasDjbJnyzOqjTcpMbyN/z/yM9I
uOs823/uPVK3qA5IoFDh6BsPOgWlE6z1Z7b3o8eC5EdljfwqXSXMhMLFyIP9
N4RwKIfbr+qlG6hiSRPWljUeVkXO98o4tfvAjdfE4bjhFwcuYqU3fiX3QYgx
zie1DMIz0tkkBlQZK6ofLuEPOYaNrkn4UH9kupvKSZeDOBSYEH6Ulbr/0qCV
dKcW6rrNDM9cKQ8WskIqNHXhqCOp4swy4F6tQYv7zKqIwzETX8NiaOa3zNrs
tGQrKvFQIyMu40Fl+zqmMY47+dvhX5QjrDTwxr1U9oEJbCCBwLJrZRwgwfkW
6NKqzy4sRaI0g9pt78DPx2AEezumdjL+13eJSQY3xeqhEYwcXqlXuI+GbJRX
BPQF97U87e8VMBD3MXIJPICWEKHJONuAKqseoEXbOW98/W4qD6e67+UyJaRH
/y5iZCwc4yrznRC6FALYraWly57Vn3V7ZenMfxb5ttNV3nXURuOm/UgGowmN
DeDx6DZAzkgLo9aEC5Qm1dQNo7XE2JctYDVXIDAiHkx7qXN4NlwdAwCxpgVi
/fUNt+gt3r/pHDwLN1+yo5eE43UtBk8sgN1BQGuTH7WzTmyYuKY5BzxAeX9p
Z3hyXTPzrw/DGUWtZVherJ3PP3kM052I7u8LubzCMSY1gytnsCLEGox7GMRM
eQpFVIwyK6U4Y2L37WZc4vOb/pmDPGJ32nGOyioTVVPqgYIifPcjf+dihpn2
bBU40jyEnUS7uVXXd2YgZiI10uczvgiVTmNPzt2bckXKnlqQyVA0RK1psGJz
NF/+q+5/PFD5ISEFqoVwvk96sAdVy7363FAwofWM6um4Od7LxKArAtYSFyPd
HxuMWSs33WwM0AmrpBpcg9qJ7O8Rf7YgzEayVGajjerZW/Bo9GOMcR4Mvxfp
2kyiVyDtia0jfmtAvwxhlIreDo/IwQ4zE9YPjxe+ZV3hJNtKbuf49QYW3PXj
TVr/J/PaWOKTzvT8m5mUavqSP8rRReKEaDfkgJD2Ip+O6fizTdVrJFJa3hgK
KHr9GzdCGfgHznegFkFN1HC4nebE1nfCfXf6juMv0O08YDrhWdr4OssYCuyn
iiit3kezdgcTkSxqzz0UuwvrOEMmfuPklCmDcHhI6qcKiA7UQyFqenOnH/tm
ZuIOfXprtewpkdOdmCURPwVKZKyGLujNBCw9HsGEPlNiQEsPTMHgX9yuSZfb
A7YBYArXrDA/O34KqpF3ubAnoXlL8hX0B/pcyRuS86yV+UfwyJlYdn7dL86d
YZPwE/IuGY8ozZg7pBTVQ7JTfwIdROZdcTAZO9xbWbZR7Wsb1UiQ7+28kYg3
6Ra0sQResVcA1D0tuUKAii8GALzyWpptCj7ggaLK3EVXuzlRtegmWk49937C
zVTrcxI33GqTCkCvDyXpUPlKHCvonukGH7Y7YSMwfpKhhOdcGOLmVLnmElIS
Qp9hF+Ggr5ooYCXhFAnPKFt7oWuzwwx++lrKVeUCCYgtM+XckQX5Z7AlgOhT
fr/52aJ9V0Q1StcLmJjSTA/m+dse4w17rTpAA7PPdkvpQyeEAF50WLj6Ed8Q
ipMQsXLwKkLgFYY2wnoDEsNXGbZ0r3uUCmlAIHGQcnxT/gN9v5vYR0aIg8qm
DmlcbojgeVnXo1LKnArZ1HwgmUVIvxrZIgRRkLB9L2YRZz03jitjP147HlC/
+XBimSPuZFMjbqHjUFry9f4+PJyIPaEcyR99cjZMjlUrlahGZMapJ3Y7yCNQ
f3nm88fIrhuTUf4TEUfnVUhtpTdyNDyPyoTCJeNSKxOfgSksCkJU49wxYo6G
Vd+dDVYWLJjNAmfGI6MsFCNfOkbYXHGZGkIMOJArAqxwgKPEwgpVs760zt/q
HUpg3roXjkwLQxXCc45MPj9Pqmp82gvyp2WTxqwaMk/RYl/sDcCMp4a9REGu
o3NueIUgY3PickfzJGU8+Ky+KurErB02NJKmLWCig+e7stR7Xai/QG0xz9Sb
1/Qw+IxLtxrymjIq3pqsMqjf28ZzIH1JOLv5Wkr2A03Wl9kSo28L2O0vnqYr
5esuLayb5/T+ow9VQWx193tXsDwxnZ6q1ZaXaxAMkV3qfdcePLtmhuGaiPJA
4Ds3+l2pQaUpKFFmkN4OlXBa8wyMZ7AHoNOek3oVJfVat+kxno1FkZEgoalz
Q61PSqJMMUyE6l87Z6DAwglXJVVmF/k7lL4kXtiZ5jw6ykyYV+HqHsgHm5jD
Gs3cERt7EkSQ9OWuG79wrPR1P/XtL0R6T1uLrNSeU4RzWTk44sx9jYi/fEzx
pJJCrUZP4aQPPBGhmbwQnc6GPiZI16DGzdTL5FNuTwtWRHZeNbKcYL3lXaE8
n5VAxvWnVb94B8VkhZ+h2vxgronAXVC/gTZ0tc3dtHV6k7O6nLU7xU40t4xz
vZKXhICq+vxnoOOxyLAo/bOtRr77oPMMPyfxFgHN69z56pDkP/NywuI4fPum
8Fsi41Tfc9lzztEuzTRwgfA8XsDZUHArjnm3ORB36WfYX+su6UaxRcxxPmMc
JfJUvSt6ItMkpnn2vFd2MZtQJ/w1PQcyaXgws8uXnDQDkMJY4r5ZjXcFdxAz
dyg2i6qH8P53H1y5WgXy6F41R6M2S+nC5aDxPgCAKfQIrxw6fxH32RgjaLKK
Wmt7dRihKLXRvww5BaiLffcKmyaA7BN9QNZ9GCXxpcgCABsLlcz4MybTWIPc
eBcZJ+B2w25/bzU1PQ+1vSrJmdLGr7WWMGDwSv0CyCh8qOfPrVTclbR1HvF7
gCsSzqp9nF0CTpwz0u/u2PBqlhgc+qAzRR8Fv78hN+x0FHVD38VQRKFbvYy3
AOaOw1a3cBt+HdbGDu+O/kNiEC8Jbas3ebm4FnH511IuKRoFL+uoW/hLZYi0
VgkfBEkikISvez+itC8orbSvrhp6OgXc4PgE2G+AMeAlZk43PodQow9cn/d9
9Kj1QPZZI+SqGuMPFISk/zwD98voU0W6GZN6OAbsiVjMbIcc1wm4aB8G2FTU
/qC8XOz053wXlgl3Yy7eM9944/w0O4tOJ8TVSOw+M5ouxvQ15bZijOb2bRk5
YK+r0fmAi8TN00sbLcdenQzliYew+eOnfLVNKp1msGlOT95Y2IcK47Ikam7y
218NyzLNdhiPh+NmfALg+RD/b5oBunWOXhnRLFi0Sx0K6h5wtn5R0lRbRV8h
/vVHO3adngrGtCWLMFkcaX97abtx6uiiwHR1NhoF/+nTK/lbQT0inisEmO/q
oGl0xWqcf7OeJPrDovXUTJU6Pquf20V4scXCLzpWcqrd9eMjzCzWiy/3UwAt
xqW3hghTOzr+1KfcRo5lTDwAPaVKgtpv+YBPRIweGUEXDHblZeS/ZDPf4W0R
L+5F3juKmgW0rc1GHwaJoK26riRSgxFsZJrv7+AryAqoY/l1P88ltxFHROSf
o7RbtLhicmi8wsfZKQxj/Gy23BSs5yxjFYOf/P/zY3bzGXes7HsksQz1FKkF
UfcCDbFmC8WrTKRWwl3pI3unUhRkjJz5tCebiYeIxe8bE3wt9HkoPOfxQx+q
bmnzVgx388yp/ZIEBOtKp5CaEAHDSHOTXzWZpo7h73mbVd53Rl7V3F7RIJu4
Z3d/UeTvD7VDw3OKnk8tw7fWSJmB6r7ub3zniusTghFeKOMf7otkpoiLT12m
JLaREKLmUGAH7XrU/Vh3i+WcX6qpf+EXwbLou76qBLRepe9zm4gmLeGsjF0i
+BdknLc8KVE+J+KCcVg/WSgYR8/uNq9v9J4F5OVmGYpvErRawZxTJfoifRMl
kqWDAKdrSAIQQfpaobFi/nrohrd0ubacUvw6nNklkUjUsf69It0bgiKtQ21U
6XnKKZoHtWVF0krkr3zsDimDLYsffFBos3RgD9BaAx6M7UNeRn6+nWxHP7ks
P7ABukzRgBYhplHM9oLWja0mRTMGni7XbyyrEIVxKH7Btqlt58pnP8CUEX7/
e06/9Nt+kR+QB0H1Mcg7FrCVojhvJQ5Z2fCqae81R5luQ5lvWdsdSmOGhpFr
OtAinXnYlPlnho7FZ/BF3BFYDGfBtOr24mOfQ4wOzaPJibfEB5fdtemxReCf
ged4tuMUCfm7pbXZZZs4f5tAz5v5JEp2UTTi2Xrse5IalGWi5neiOxshcsxs
vohNEAqa6R2Tpae4hU4SFh5AF0Mzo7Ml+UXdHen3IJ5jpF/S9FFMakjFEsMi
mQg3xQEcUigULrdMXlOhtE0+eIdMOBPx4s4Fm3aq6Y277uJqCvdaRasuVtoO
Dx55Yz++ET3k/9hZt7zb8Vca1+q608cU3ub/6EHsZ5yX+ZLREhHdeT0EqOKn
abrxmrd/8ijlEaDI8xfBXo4Gx0Y5J51G2LUcdjjC4K4pLeCizRgAYrcQZNpj
6a2teWde61Q1Y5/nNxEmQqNr01SYjeY7yhAdTDNc5DWsJmmJh+vzkObVNiDB
3/yEIn2WbN2mgkd+cMKyB/iHzKKcmmeTqo1HxMmvY9NWqu8fihGIlPZZThch
Dm5PVj5bjllQUyqKa1o48mQtRDnUJWMZLHTTlEvEOjGSdcU34/oBK+CekSeE
Dhn3Bi2ldHB4ezsznEFdYQ30S87fo3Gv73hd6J8m8lZGN0NUorm6fXyl0iNh
x+1yBZFhh6QXf5h4Dd545KWx0AzRZSWgc0ehglf6dISFSIzaJOjCV6UG65lV
3vMvi+lD0EtQHFn5y1mCJf1t7LWGEr9jp3ftDVKLdhTAeN65TjaJ0JNEFhAt
ga3Z8T9PW1tCGCr9vFTCnQcbmDYyIQ/1dMw8ksiDFPS5m2GtaOD2/DQkq1Qx
Pac/dshRdJnBo6poERIXUcRhT7tjX8TDhaUFhiIfsYQUpmozbK2EOqOPvmmX
HOkRuZzrXRq3N6b/MVHI4LyDOxFV2V54ZK4ha3SYDmW4lc662/qRdQiAmSxA
imgkXNlTp0kxJKurnacV7oaO7SnAEncNnRCQJOOw0D6qDx+t1XwCdZMhiJeR
9KpkBgKNBIjnl0fUIvz8mMIdvip6ywHZpjoR1QlivC4GeBEguzge2awMnnId
kjPUxd6ymnTxEhbOhL1FsG+7Ol3LKbuBEPbn47nsDzUWfA4OsYuUdbSGTdBV
UgZFInkL/onrPGjIhM/MaaxNG569C4c3XDjehpxpYt7hSKVm3COErt9Htr23
87K07r5VGcu6UhN2rjrRN3vs2AQjRQwbt2zuNbWiQ5m3kOp4Y56iKRZkwIZn
PQ3epDGwEXwvX/ce3Jx0QQw7c5AcwY4+xP2Re5Ne53cbw1zt06i6WYnnEBiS
vUeK7Etqz6bYyYf8KgkgoRbSQtOhyuMM2s1GObqwWmkQsaXnnwQRZUuyECId
IQ3KyaaljZ34maIPRKqPVcffRu639Om+y/q/M/bzCgfOX9u6uxtRANfyUlmp
E4zzPLo0tUOUbBdTanT/JNKtQDcbrRiS1hZeBX9TsJkhD99Sm+VK6HM+HRpv
rOK7ywG5R7lTyOxiIxrAqH1vs8xRH3YXFgS4GEBZ+ZVNWeZtdwPhDFcot1m6
03zyKCR16jNPtM2i7QQWRlF2vYGdX1HJ1sqNETm4RDgxZExO95pV5M4HH8Qn
VOJVnb+75vxLdcUwxEJkTowYt6zRQVsYHIMFCvpYYTv6z+CmhNSu3MhwPsE1
jp+NqLhy1hrmI2hkmrHz3q11vtb0L79l+KBZU4UCQL4JGDb5ASt5dIj+nF8U
UKIEuak4+0CBfW5IcTzRqgU7VDi4dafP2tLQVWBsdOPylmntErmPkNqf5D16
rhy6EZhPlK5661mmaQRtKfDwRfD+D1zcDyApu0jEFJEzjMKPtzCD/at4ukHh
PXJbY4NxgswhwdfuEqM+WIWU9wlIud3IxuzTnAXc0RqG6zbWL7h+HthWKsDe
Yh9O+KVMgPOCnacyQfFvYXvMpxcgHBXEXXS+4GMjJbA+QD6jpgeSPPksko5F
CuHwm/7jjv1f879HIt8KPqzKrkrA1yd046zolsbk1f4GCEmIk0HCqxu3f37P
ZNxE+5wFGXPMeXJXaZp5kxDkXuxV6CzMSsEbC2WV0D3UmXsaOHz7Kqo18l6s
Bw82x9mGoGwpXqjzJVI6y2E8k3ieXvBf5DElaSajjQqbOHH4ekmp6BRgcV6s
BteUZEF6Ir5PMfacY6KOBdpB64YWkTKcDA613CthKCKwgXipyzB7vETdSzsE
V+b24bfJU5BS6eJURnD1Vz6axMX2QyzpxCc4dSM4aWdqUITew6iD4nrO1m3A
xJtxfdp1SOs0NfvcBKtCmhfePeqIyT5AxV76uFg3DDRfCOFXQ7icmD0elIul
WlAdTHuOnVo+oLnmHktkfuhZfvzuYIXwOF4DVSKTPQrP4fMZZ7YgZLt1rkWa
YkyEN9DWe6Dznebik1ryAoarT+ZdZBtu2kJkSPJbfWntD4SkA/veNwEAfFAC
BNkSdffEAh8MHVUsqX/6bQ4r7vont+1IwPmh8bc0mXbP0jG9Bw6/+L9dTdIk
pQGKIiPwFDQXrIQV/NCBywFAdAdqz+brk2aK38ARrJifG7q9n4FC9XCT5TY4
U+NShFM7EIl4rFospqjZhMDPqmBRnjf5DH7jKnsogwYeeZ+viXw2a+QdlNx4
ln/UFH1vcMMGkWFGRZWykWrolFNG3rCGr+HG4SfiFIN6CIXOszep7A/92uzo
rLiINnqlmU2EuLVuHuQ5yq3DlP9PM1T3zTydsszcIHhGsbwYxlAkc5Wbrau7
XJCrKaFGEaqT4Vy/9gwuC8PzFa2zPDqZ3Yl4sT2WI4kQL+TpZQ0+Eh30BFEc
usyQhbfC08FXepKrT46HA5dc/HQDDPJkdzSM2bM9Ug5GlpjxlJle1iVVjWFn
iEZfUNVsHLeBjUW/XFnsUKvcDOYdsfxP24AfrY/8/wBasg3cPaMNSfxYmpv1
QKV00aIuNLei1einUZ3h5JuMVOfPoWzXl8WHGFLHAIhyBhDk29q6MxKImmnZ
fVmtYYkBTpKwM/2kJvV8dur/Mbp1KgcBYF8oXkTc6gxcbwTcbmqlWLuN5uTF
n10RjPp49TWiOcYE0QD/Xo/ome5yOKek0pKwpYl6OZOqb63CXZXL+UULRJ8N
+XnnhlwmgWkUjcPRY17gdzRF3nyF2+U3Yb4EJxpU9q5rk0gY3votKHQiAoE+
K68Mr9hf1hgEkxBSbY2hOW3bSrhAy3RBBDnTbCiHZZNeTkS9UEbnQSRrUGBA
tbeIgW+9yv3XjxGAH71zItRrOt2EMywxHHfK1UCb4rDgRzlDyeszE4dcbxVB
0eHrHuOE3b5u9YA1nx1lHCidiznX1v8Un5GMU1IIp6oTvN3v7AbGTuBJFxRn
ceKawL0ZqFSmgt9Ok55dsjyP311XD7QOIeXxduo6CnvitrYbehQeVkJtl4zS
99MUzuATmhLPFArIytmGhUi7lNYF3hfAtbzz2qJRu4GOzfHM/Fj41v7rIuqj
ROkp8PopdiJ8G+6kB0KrsTULIcn8ORh3Wo0DCELwEjNnWmyWQfu/dtgcyf18
Jx5UaNu7QxX0PPvZjUJHMDBXsg6knzvS3XfJSzh7YLzpliUKTRJmVaDwaUOB
nW4JkoelUzTMNGLyKi2ATV3FBO4wBGifqpvmXmNNm2dLquUQaLEv+nGCjQxl
ntEBVJb3ZBDNntnmUeu8p40urj61d3NxRpUxwIo/sDL4wOEPp9pnc5JCkVmL
jf6Z5BIhwwb84FPpNMqBZiiQBbJ9vrsPUPIGeWiv5U81yVG0nvOj9mA/LS5k
pwdr+cinXO4g+IAuB90z8KGGnXHpVYDWUFT8ufjyk9Qd/xnQJilxhjtT53yk
FhGLAMl4sL8dK6D9IsFIvDUNtdOla1UgoHdchdfwxPcIk0H7wkvSxxdddAXf
XL9zMXFKmCcqA4EhzCX1le89cOuzF2TujZPhE3pusXSkMlKdNALVnTT7HQIG
7wPeGaylUUKINjhnjKWWr+7h7Yc/R0MZoxS9QAkxPahNU3q+dHxZ84Xa5BTT
YFlMF/rZKCNSG90MDDCjJbNfYJjRYZjJgB8583XQRdWyQYbK/xmmTdBvcfih
RdPRKgJvjgQrZV0vBnIr9AJXMv3+n+cYJ+xg4XUmUUgCaoECcLpHcd3gfwZM
HcsOG/O+woA3W3U/ONwRlhGn3ETpV1Cnx21mmpNNMqMLjJWS7E7QyYPri9Di
Fcg/DBk558sOvwEcEAnhQOdAufQfnJqgcfqxRFC+QcTmzwRkN7mNUEQcHUVQ
eqfwsOcToSvH0pxaVGdG7y3vnNppqdrPyJtqKwx4ZtKT8Qg58vSg9TmAQDNK
BIDRV5KaVzvkonKK19klt2QSo1ZhkMlomJn3ETaZwtDJ8nOK3kij/lmXK/V9
p2VkYuBF3Wuae6oWregtFUxpSngZRRx6mVi8fxlgdHsRiomomeZognPYD1fI
+Kt4SH75wiybm7M8K5XnIhFRcYVq4himdE0wHAH+cZoG00/bxpNac0M3+pn4
T3r9+l/xryjoSMXuC/fHRYr/XUcZ93nEuTLfLDp8MvWN9/NpEcwaIEpGs3OC
foLjRh9pFRHBh7pm6hyP9vuB/GN3Kf7KRUtQJznoR4blOgjtRGyJ7snupKkJ
ztOPVdG1nPUYJmET2MslXxitDKpGIbFBgF1w3Jb817HET31SIsgoxeQhu6e/
k8l5LKaGrpqHpXaAHFKcZu2y2ZhiXyg51Q3VrFTwLU128QHCJfeA9Tpow7Sf
pPoPTWOafkAct0NL8uY1/UbrLMfXNTTUwCJPcupeC0v9uPxxZAYIKk/qfiLF
LQcpqjzz8wwuQZaGkMNNuHQHgmgakpam/PT8FbVvXoLT5HFl0DJrNol68HoZ
FyjrKIcissJ4kZBeLYgK8T/Ecbq1vEsqU9eVPUqOWd1DMKcLtY24rNtSiOIR
vXrofhDP+WRnEVN/517v/zAcqwb/lq1EXs4wq+i/s7j9k+vx+UiEpHi6viMS
cxoAyuOnDSRwBmsqeCVlLKafxWA4BVFS6ULI8LuYQRPqDRP+d/z2stRtTW1X
KNOGg3IMb6PFqO+gbGLXuNbUUP9AHVp4q8JCDqyzqTGg2EG2tL3LrH22REAW
B27AFX50cZuDa4Kb/lCv6QyCtb01EBl6BYwV/GlNwtEZ5hwtVdPjvk/aHVHp
wY4wn0mFFGFJJklbOQ7ryqwxc4b9h9QobdtKQHbWZB0E8KstmM/Ncput0S+y
1s/2xKAJHHHYK6Zsdk/2BiQGBP4f4dRkIKLG2aI5lRXEjNYwYze/wmFrOknp
Hb2iRVIqPbUV0KKJTmZL9xsdpxwh5tPAatbvQx+8pmturjLHeuKZXzbrLQS4
gPt9jCROHh5upzTJh9vWtBVGufcNvJF0O7HvW0Tb8lIW/aZ/p+mNan3WU/kG
+8tlUc9q4wMJM3E+6RpIQz1T/mYqMRVUL4x88lKVn5Iz8TD+XdgB+8Hspmrw
EQav3MSHyya6kBgJaheKC1E4ns+eb9X7Em7e1GSRuAxLQSgjLK6jrwOZ2jPx
oHC2u0jQNRLKA1koCsrEeow6IUIgiF9DN7rJe5UWBXOixJM3z3KMywKVeW/4
WcstN8A30csky1WOpHKPUlXUcFojldS+ojIhSGhQY4gw4mWKnNZKlzxEQrzt
0fCWRRTzxLq8aUA1rjYpEvDMW0MwBLGYcuJHrm3lfaSoVB5fma1MS3+zVIhW
VBoo3qSlgfa9MQeW0wubvkOV9q6nnZqmrWcxG4kecftZjII+GEw744iJDnrE
xjH+IUajvt+R3Qe5vv/mmpo1OwbgyDPOFxO2NmK5q1Bh9CDDYkM5oDjpgGX3
jBN35iOn4UmNlgV86Ceii4GB428jR+TOs3UMPTGP9Gqm3JgdkQaCsUVCvqBi
52SwUSvOsq4QGumsosLalT78ZNmkkKUw3iSPLnxNf3srrteFD2xIAMAGzZ/Y
oa8JMPwmHsYi/fnRb5oVOZQQQsZsEnAcJ6iJs7dMEEXspD8XB1kqdMPv8npJ
k/Ud4LPgEDvai3mGoiMTv53Hy3VoD0A7z9INgBXXZ5T9wS1v8WAmAWECwS18
hKCKUgBGQ8YXuGr2IIXsn/6K5sRrZTwhJLiM+p3eotJGlGqNX3OFnhGEjM1Q
C+3EdRmJEFdUDMbtwy+Gk6LS+80SFzqeo4ReXcP5vqzrNCgBQolQigdLp1wl
cUGdIqCx8RUDxpuAcy6y2vmD1ZdTAmkS2KVeRFYpiL5WcxjQNpFCyQ5soU9b
0ustzfscOxTlXvqV5x8xagW5qf4yvomiMUftIj04Od7eUVIL6LsRAZ0Ppl7f
/cEm9nyR5vobRCeLEn+Oh6y5F9ybYPw5fKVqz3xNrlyYNyUgHU3Z+igJhSMT
wfcv3b709FpSfAKqEXPNJMlcYPLVnaI/bgetiVHevPUDwZVqz1kDcNEMQ2Cz
EGR1KKWb+Dvw2OCZ3medRIoUXSnceruk1jBZiMjcwmExTG8X8ReNmJvC07P+
JY2+whfMn4CUvIwdOWYw99eI/7CfNgbd2VXmNuMfOr0lIHGbgSS/1eCkzDZy
sWAvuLKevsZud7DnYp2plXAl4O9ocAeTHqBCm/EDGWR2KUx3Jl+owJksOv4M
zcRkNp1QTEM1g5gJVCncPQN7cxmRyItlXrwm3s8y+MYv58uBopcdEsn6DEuj
IMURxuG3t0ehH8Dbu8oIPpareD5/bIRs/5Hs4IYnGtnY8gVa6FwjhfybEeqQ
UaJEpSOp/0C4/bl2wv0YfCAKh0ZYvdZY9mllnTrKpGPJISt32g1N0v79EkJj
J6iLK3JrXHKz2HRHgeMiWskI1M07vZTnq2Ws5pE10HU3Px7zQf3DuuN7iQdO
Z/uLqdMrFyZsICPBUZqRrB3LjGO2KN6vu502v4lDq6XiQ/s67ETnBaErrKrs
bOiLQ/9gnJ1Rs6qTbQ0lQCAWmY8+7LcGcY0a19NTacYk1gQo9ePtnXJw9sWU
dKqyfGn1BbfgKvEBVAwvXLQDaRbGMHlq0v1eYF4ALmtbAQFHTVaJYlot2gzF
f4icJikbEIWeIKjy4W0fUQiDnusrMIcGa64HkW/tPzheJDbCI7fDEeYZkT1K
xhdEy8JQZ5modkCKQI+e6MWFAQpj6onMErhYi85ZURR3PDu1DLDABpnSaSus
MsXuP9gqEwO8V4Wb3QzpYlkVPmY29AuMXUojr91NVYA1gfB/afWiFtjlUZri
/2LAjuglgTKmyobedchqDJCT68BfnipSJRtoAOm9/yopVy04DteJ6EVexm+7
8/nVvY8J85zOa9z0VD/AzDJrVDKWFIXE9eEepjAVIQsuw8SO/knD1xaaBWmb
iuUfMo+/8y/HuanxxIp8rPpEJdr8KoW5V6iPRPWm4aSqM2Abdlr6JtHwSar7
YxAhPblzmL3CHBV7XueGN/Ccf5uY/LU3EcsBj/LTpX1RH0mUQWC3ontpO5RL
oLo1U8SxG3FiqKUk4d6JH+18k8fNUH6HIGEGQgzF8/PZEyQB9bU0IsrpHe5s
JNebpXKGI3f8WCn0UcDPgnJjZ4Wfb+eMaMBY4Vryl29oVfH8s0hnqu/qlS0L
L6CqaeYUcke1pLoI/RzUyhIlaUCUuTPhvQ8Pe8jydMeE5Qlyw2Vm/qw8CsvH
wJEp5DZUDU1fUKtmr50GbM6zHdk8L3BmXg9h61DQYmv+b6Hrso/yDKE8OxJK
vHtlW+4FXxB/iDjf8cK67WghbJtZaj762W1y3MYB+HbEgWzCZtjnChlwVolh
0Theeq5WK9ArVpYn8gQycuqWHxAo9o4oDHjPb7w/p8K9j42fsa14BRDUbarn
ARrbNrg8yLOJv3imuAfBbs3AAVRqutJ/oukVHtf6zOVvWQiz4gxrqffcnccp
aR6gCAEudYXtiwrJjpo/5ECtW+4dvf+MJL8sbgDzGKIArvNAFAPgIrgYbnNq
STOaw0o30OAC6dIyumxOaj+Yr8LLBJ/A/mIKudaU4V9hBgRFim9NTAIzrswr
61yQwixcUFCr7zl67rrOGCrLrd5HRIuABJhq+267UOPz0+zbksiMY+EJ0Ce0
MQ4/nAkX4IceIr+Kv8cRNaysltFe75zTgreqpddlB8icbQTHigkZ9UZbgKm2
AbEGEmYfqEpPl64ijnDTqxfj8PyU3JgVnpsxKKv3vajwRbxLNJIkiaOh7xH7
lWGNMfwyHSmHehWg7HlVwPIHI1PXMSVUwOQOI920KGti/jRCCQJESo2nLWUa
tbIBto/4ADRfHMQa5jCt8JjbGBs7KiY2aW7wtli/q63/7BdTUHki0YjU1n/t
aes1GIl+J3318SexLcHAGAGWBeNLIoiWAWrIKyD6IMdgzUu5cUy+JUEmb0e5
TOqcZwWXuKkhIF4y4Nzq1ArEyH1u35CFv+deKPR/mJmOSeNNtChtD05WWX+m
aOV85zS5d2qqWtm7N/ZwCQ7+HmEf+Uf2F86uqwYayCbAcCVtGpl7I46/0kt8
G8MNLnj3qW2dxEPerA3i9GqnOU17AKapK7aZp5JknQtIwZOhRJ/dM2YqsIN/
+qZHyx/Upa7SOD3sY/AuppmfZahHKqGE7kLVWQtfKNtIyC3q2B8WYLSDRWXw
hEWII5b+JoZQMv2GteHtoQl+udPX8i7tGDzF7JnPSaMoST4itqmy239HGYD4
0NEQwbg/PKIdgfKFZ6dWDSzlSeDERgXH2HEIwG8vJkhQqaNyWEBpAXUIeIQN
UhQacn9HVBmY9EKdwnCk9c1zGr2KJtUFKk348yChT3QXCTA+mslxvZMoMO1Y
OMMHAwKgBDsEAWJGTfsZiCrjnNZmLQsxurbfUKF5hVNCegOSuL95pHiMLbZq
k4hcwBeMqxMgYECq3ctqHrRjaOoE6BrXLKQktX9Ekmqs67Dtn7KENs6eXF1q
B5hJkuW8QMHFmeP7LjHNkJhlpdGLbSn/pRdXoKCDUfGqmjBj/o2R4ypb9gop
TXJnmoSiRBisksZlI5nb/uOvicCJ0mlEwpyByT+49hYZ17G10Y6kJvNL/M+e
Ls2A6q5jutOjKicQiJaqacG+SyAwWPkMScDA3GqjC7wV/sw0RfmoCYwMVyob
kd8I2Mvqgu1rKtg+xnyRN6lYlDvakCSZwfDPmzmU7yl9osCu+u3Qmn7hyohx
pVFIt+ljLYJDWk49ffv1QX7A95ckvfuLQkJ4X0PVFQ4tcbSxSyeNFWR25m28
0np2U9I6N2EjENIQoZ2/DmqdcdY6dmMMWjxrwfxK/WIxtGNykSVeI66fsKm7
5N4nZog4vvswHHAOdKepE3KYEDssvOau1tE3EUrFWpEl7dM2tmN6Ew0499JI
Ns1ryt6U83U9PM9cvjUmPr5JbcEQbDxi3XyRIiG1E77O9wZbYVZy3LyfLfkJ
MI4H+tXg4wHNJjPRY21rr/lvpHh3UsjY1lx7fIVduDmQ3LJL0Xi54u+Phdq0
t+2a8sdO1HjWAd+TgLjs4isR5UAabdXk38kVWSY/5r7m/MBENJzoIg73N8ET
bin5eir8B2kc1bw/+0IpjLTXAyOM/yylkgIj66c3qXsNpP02zEkssWgNj0qJ
337GvJTOZT8e5iB1xsQ14VL5of5eLIq/vWL80ouA9vhmmzUawZNKP7eGSdcb
CvgteRIIe8tGpC1UxCMb+Sf+Gm8Ba8kKswZxKff7LUocHuB/sq1VLIEp4ca+
AZ6bkQ06ajzCa6oMi8DxBOYTuBv3pBZVQNP9nS3zAeAtgdJSHNwGT41reXxL
243Bfi+m0p5AE70iP1id7KVNO/TIZ/w6w8rSNcOMiHxnxlwhrTp7AZLEsiYs
lz6k8fq3GaKfNzWCGtvCUExgFvGZHMgHAuAxoi7QI+jnIFmn5MkELxZVjGnf
BS3kRdIjR3iKbdRVAFViIE9aQ8oD3eVr6EZ9ww5MsuWh+p3lHjoe0n9twoii
FFUXeqmXaWIpmTZ71PZdeN3njq5iYyuZdZC1KtiCg7ftIOtXg8x24gRroPPC
gcoAjq8o5IyN0bI5h3+3WVOaIQvhwjchn3DLTI/9DMnXGZVVvFcbn48K7gdd
qjshb0VcQ76vFINsZAhRp3cXnP0pKg6Jr/T9RDnPvySZdH42MOkOVT6q6yRd
ibvSheSyWvx1mpzN6E+gDCP3uEZCRWq+Qutxk7y3KsU3pGx8b8og2828YM4C
zOpXryCLuIu26mfYezirwhk0NwBqGpbDHJfxEC2NuV0IOxu8rkhzJv5veaKO
fuagJp79ONVQJHs3Ti7cLnpc3ZXcM9bugjrbvMfemR/oPCxJeeuEiz3xZxBW
BDthWU2+NHPWJ16u5KoF75ef5NJzWDpZtV3Mc4yb7shIbvpvUda2oAeHP0DC
8qTVS3gYywV33mqZ0xUpczfFL7Cm3KW05H/gesipKTR/BMZJ13V8iauAth4f
arcpBy+QbBG8/u8yWrA+1tUbI3JiI+DUYMEUeC1upjkZyIraDRpdKixNvjpl
4QtDdoQH1Fv6mE5RnysSXr2xruOPaeceb7iIf9emPDMQUFmv0sFd9fgb7Opi
1TW1qcRdG6Wrixvmr9JTfSnJvGnf+Yxb8mfgQNnnEunuxSs4VkYsOsaw1fiy
rMNNHdQhzbc63jImsDnUWESBiPQRZPXAKdXtdv0knTWRQ1Pczi6d/jpjk8pI
7l+GWyudOERzeCdPd8Jk5fDG7I5pyWRbmgWXJM2OnhHC93mqkOZkSBff5tG0
Ahn8FooVwI9jNrGiy+5yYoMAlGHaibMohM4jK7UxZWHLkAo7ignZWtZugYIn
kKuT+TPugFrDPzVRwyGUjfVMeJsgoJ1AzIAYVSVe5mCAqA7kdVFxmYC7BFjj
xPZD/SKEsD1aR8HCRGKE6vm/p8mzyoGUiRj7nFCTfuKa3g72I7+/ooNY5iLF
htLEAx3vAKOo+ZzsgZJPKu9MUgHZBCXDlFJC21SALh11frjSOiA9Mj6KxZin
fNXt62Kk/2mVepEcCQufd1WbvQprjfmUpnDEXKPXuifGS5Pvemk6UhREw0l1
SUjoaE7YvpDN1DtEyWn3mGqGJ3E2yNNLP6zTH1LcobB81qoko4rI0YY27TZa
rQ9YC7uxakRTmg+eJ8cNIiohoVkokL1L1a7wb2O7rDMeb2IZGQk6xDJ+tIgA
SEXA7azpAePxjhZ3tE4LtX9ETzkj9toIKbPmB/4Mhz6Im+ZdSruUYPTxUweU
4a9KNmWfdiRUuki/+DM547NssY37uyMI1poFQHLaa547Flzyte1rqjGMg8DV
QAQaLd/RCcHPCOua+d+DSe/EKCLuL9MlLOPycYYic+rpGzO5Ei6LywUCziwP
yb48awqQpBCJ1XEyjOdQkj8Rqj+63aRMlVTOoj0VdChombNlFSMauHHQ1ikf
NnMbQzMa47xDKsuGic5GiieAX8Bg9az6SEiFPrO9fVyoaFrjrBD0FWiAbZgd
3zHi6nPimmLCyHWryQ8bIWWkfedRMUdcDS1i9dMrckI02WyDb6y/djmst35A
VvxBNn/74r/clBd4Lj8+W5QHJ5J6ADj1aoE/CEumz7otz0+R3FL5bH0Z5a6v
/SFCx4S+agZktMR947YvMp3GteFek3IUA+4mWUXqmS8OlGxR22+uEj3eG4JW
Bh6cXp6Av5JQDHFzV8URxVmL/GhbpfIXQqV9nBrRxcHYLlMtNSsM4qrjGihz
KsDaWAYeEsd1diFwkKvcahfHhayGssJHRADRgG+K5jbhKZ2N5E0r0w0WfHhi
T5flQvzhtbwMhwky7SGd4AU8RZ8rAesBlt4WZtp8aJH7FRfjNQRZguPuHnbT
ZrTCSoIGu/BWpiuhSlfAjpim9eBJ86XURS035ATudL1KuflJG/k3kciaKp8G
xLE8IClLSydyMi4Hrhkr0EKA2YyJNNjOgamK01zUKe7GIDHOU0fZ8C3KK45T
28W5i1EiDJwdv/qjeqw3spSO7pM0niEr82Nhb5PraxTqU+hsqZtgaPpq5kpZ
NZGM0X/v1EW+DTfMBe2oHEMgcn3QG297hR5uigmN85YzOLEezPlR32yAFfNf
F9CsoxeRYfh4w4RPbIv073iEQAtJHt1/rRXBs3B6GVRRAfg2IK/hcVGBf7zV
ntf2ZTkbfexVM2TLNuPyry/X1kBIkAr1jVfWLQzazClnpKzt5G2KoO62yeAm
fJVN6COM9PC5NqZ/Kcbu+x0q//UbpA1WFCOeuF15z5bKw6on/dTr0336qrjn
juV4vmp3C63/tE0W/LDHxoWQIaMsIjZPzCJGUTdymoGEgZx+pBdfsmjjbmZc
JGP5URnWB9MouGeMOqCcGav6tSeSN1mZtTM868hPCxM0HWdjUcpd2hTuazjy
HKXhjq9o4ep9TkSYAVM4sTJLKWqvFgEbW0ZzpR90POh+Hm8g5D/362FhJodk
wXp3GxWMOlN22DiP4y16P7PbQH7GH63KiRBcoWo2RWQXy1D3Zb5NquxViy8O
HIGWMsdX/u50XJOy9JDROPa6fcfO2IF7YUDC5UkxKhU0O5PAuTJj/xFG6BsV
/GaV+JWxSLSAfXJ/sgKPYDPdqBkAaE/LHWIEwS+4vbk5tYfNJW5HYuErMDe8
UpJ74OFpAHxYzlJBFwBUzoxqepAX60ZcBlmWa00EjzVbVkewoSrEhgnUIX4Z
l9vSKXL5zWl7dsLT9wi4pqGrQiPbzQcWlMK+cJ7MrwL/1soXkZ+M9m1bxCtI
hgJm753/vzENSJaRAhTjlwUmBEUXSkJrBxEGszSnA6imsqwFIyKoXRi1ULu/
s3cRyq2GaW1apZLMjaySjVlpohMX8NyEN53EKPrRXzoJM4IZp7ZC+5Nln68V
qnu7E6pQsX1ryJmc/qZSOGPnWMwuxXYWIJm6B9D1SmQAzWkrQq8vxbgDOdhk
UskQ9Sh9xz6PRof13dpoi0dAxdR35VqiN4MCBKNbqBeqclr844ts8SNhdnnC
ypywpJzMh3X1jMrhebJ1Z8H3tIpRY2qyAyg3s3P22TcOSig05LcQ7lBqMXKg
siyuKoBUXpSSZbm4tra9niTshWu5ahDptoIlTLvQ6OH29JIT5WEOD94xQV76
DaLUkGpg1W8oRyGTiuoqV2LTsJ3WTfn28taffa+NawDJSxMC80G++RISZ3Ow
FE6gQ8zSWQh+PcvU7SpFw2xSsUGuC2WTMRYbSyhaa7mOhAO7YwFK33Ljo2WY
EeGI8+rShIrhrCAFa3KdhomUicibFOqz5DATzsPaJE8b2RpWvla/imUwW2Z5
25rbkOwpHEwAwa1Wcdk9BIxAX7U+pEv/m2DtRMyiI1wZ2NMKeGQwbpjmRpOp
xNUruczakGHTdATJPOk6NkDq/C/kY5jonanQ0qdZ2PKuZ0mgOliIY75fHJzB
aXPDy4rxFIeXocf2DAZMquAw8iBLBL5mj8vCUoqoCCMMzXjNpWIx8Rx999Hm
wuQaXjlevHPNUttkmRsB4LXOouqXdW6ZnoxGPfucRb88DCOpeFByzt+lR7VC
b13AASagAyuw1MfZtXypKYIHT53CWqaKkpD3Ytq50umfB/qwxN/GdaKuc+au
z/u6ZJ+agR6ttfrk8TXax5P58FZSfF5/v4hg21QtCUH/wGRXvPoflrdF/lm0
ftJkgeybIK0Cvf0IuIcC5oauPLMdORIPAXPajKkG5hOldoOhZ6swySvv+Sgs
6PAPhfeRDm8S3Az1/3vIuheNEDPI6hnIVD6CDwqGN34Qb4tTT0pOjL5RF84d
IACk+c+GJ7KKCiPM7NOEelvKxJQ2OJoTY2cC+JsnSOSfaGFbboJeGtBh40hH
NsQAK5J4fA+EZtkHuk9VysWmxltKap0leub3D6o20huhGaGUaoQMMKbz94ln
HymLrYcU306tEhrSXfOGGw7xm+NJGTY3Qvn9nuWePWU6MRRlLGqVOh7+pSpL
OB/p/SzjjrBA/hrxqFOnHkDaSMAo0TuzkvM3n/EIGzdDf7ndf1RGzFzHqRgE
nVdVPNvllrxMhi8UHE4+g5j2UA/AoRISawkwVY4yQjGDg061NUuZyWKIRop8
MhGNHdTHQFznoVyalGhPkldW5PyBIQhwp+PkhuG3RV94aFJpoJMSDRovOuTz
Ncq6LBuJdGdAqIJrMtEutXpxVdcyiLbsQKSaknwKtqqkSqbna7MucGh9vE5e
MfMB/C1UqpkvFCVtsMBj+U4Gv1N281LjQ8Iy3Uh/I6NJ0XcgLkQGwKHCQTos
3mUppZIX2TDjOH7RwBeVz4bP+hR2avDGvqgfselbRUWcaVokq79e2yFpKGPV
1+LB9JbqTkd4t159RVl713kvDPcZPKhxO3iWP5LjgF3jRh2FT88781VqeNTg
XeuV95HZ1nCudRwGFO4A+a0xHbhQd05f3Picwjjb+MLykJelTAm9t0Nf4FXM
x8VDfhaVVv9bMz5Vu/ne9M3+XnpwcEbwsZLmmCdIhe5uTlqxcGQjXVzHFiWV
UmD0ZdlV/DQTaY96NYwh0C0qWitVCdWPhBWNFF0BSvJKYuPkhQrJwmjsd5Sy
7v0I2h6FlES05c0oMcYbYUcz1WJNs+VK2sOoXy1bWw0w8q5t0pS5+tEg7wvI
oKkrkA5E1rmHUoH/4WFGBpzGn89g5/NGOjR4fiX71QN7oGOvE2ofkftORDye
KKnqx/YMxnm8tcK0xTjYZXY5ndNZOsY9nxAvbHtcllFW4g8oDdtGzSLsP4Yk
QtdJTwZ6GlyR6Byd0DKEt5o/u/w2v6i7NX6cZfHcbVvV11QjC2WsDkylnwFR
/XYuM30NVrJkpA+orHC2fys+GbXgOK205XRoldDjfeCEoQ0T2YfARB44keoA
FXT2EtBF15QJGgjtJbxjcRH/cigC1kt0oaEep4ybyrTLRQM3vs76/ltILAwK
8s+gmNN9Qx6yydb10kHTcgeC/6plDX/Btqm/saIcPBXYszHrBqiJ/CKqw5MD
kbxZixvZ2TCjSzwv5UikuXhb2/M2izUNDTtb1qXWRx2c3br88cPwzvyRvhpk
aHoBNK3TIGEB6xcTJJywpb1fJjb5GBYscEmEfwOPPmiDdLCyYXX5Dp8xQEpx
kUOrW4dlTfBW47vg3H50azWVPRyL57jqD9O6gMcFpEpo5AVh2zNXOk3g+P3+
iUv88n1wXDRJqhUcwZir5k/nHN+LBxbLn92TKwHJHvL4xL3A5kScBehg0a7L
cDhD063u2k/egOpFwa0IaInw7chj41wbnFwZ5PRb5HrY/ZrUEkKz/fO0aEkf
IrBKEo5ni26E6tOow1JRRgpI1rvF+9rx0VCwiHyPXgjT5ypvbCzfM9Ba8Bih
Qc7pvyinpDM+OuKhNgRdRIqVC1/FVf7kLFa89I4M6/RZUGhhHigWlPMNG0FA
PiqkI/IYfaPGkgJPnil2RDaFx7HVvU7wHO/G+6muo9LM1ei8RTg9pNw5XAfX
KTSJIfXGFEjyyvOovn1KF6ykIY7LSqHDIuAhjHtZJQNlffD8+pElz+iB7OCy
15SMCYMSH5+6spBGbQ5WdW9OHdnGgaTQP30HQdMLP2gT8HvzJomGaXmEu8NA
UiN531aNu3YYXJmVI9SzTzl1bePNWdCn2GNu+h3N2tPFAh02fT2DSFW1szvL
90kqkplfZFWsHmBy838rJ++wRvEaFmtkZ/kru5XzqhVxLeD6mCQ0gCJC4jU9
wYYXW83DNmorwofLRctrsPKk6AW1f7NRLT+5CeUqK+ZVsFPfwfgk/PCp5c+s
nACu2yQbh6VS0OuoaShnPTP7s11zftroWzU7DA4kwJVBM4jPGCcRpUZbiWRb
ZRx+yZZm8HS4ynEeEOhFwCCnotT2eo8N1j9iqeNHXU2Z6//kIX/skygMtA85
8IGoH3GvB79J/YigPqMKqJ2HaqTA6GipTd5bUp41PcF7oe0Nl9TI6zzD588F
hMsOnWCBsYlhaHTX9uVsQgkcU67JV/wn4wvOml4SC4ZRsZmzTRochp+Zpcdr
Jyg0nAOXl3+BSg2BmqKaWTgnbcCciAl3dzyomG7vaGSEbiRaSZdVH+0JZm2Y
veNuQnPSILmR6KzNecOQ9C1hA5uilK5/SHoYXzHRgzFLXT/cOLZDZc6b+v/A
qzMLLD6AKvSpy7jLxJvMuCKsb4RVxBqzJaKCCS2eDFRVPDrGRp4pPKDiO2Wp
AhoqXIwECprG/fn4cjEsZ7iSO80yxayFwOQxlJKmRurGo+MV9huQLmlGtCzn
Isn6Na57nryO1Ht4ApZg0Co2sJ0nT445Fwyc4Ow0drZTijWAEwTlJbBKiW46
u3AMK2fy7zmOPXgNv8TaX6mqV3lNOlidBrnK8KvDNFH3+hdsMiLG9jTm2HK4
9nBeOLffdTSZM8cq+Y23m/stawLiN+aNiNHxOY+SXtNbyRgL4vIa26lipTWg
dPkopjtaHahuUMByudTEclbhnlY0UQJA147lw5HDUm4isLzWYDDyERQnlIod
EtD405/NCf+4cH+Y3X8F1bSVO7Ps+9dW5d8tWyzelP/7FTq7SLHETrs5LboO
Fo0JELFyGZnvqpB1Ro8aAnBFovfyypX5/721otdu2pOKQM/JvKeTW2dLyBGC
+dJtswfs/Tx5ZPcYCokjcUqUMJRQB1ZYTcwKfV5aoCoDTELVrg1+KXvmWk85
x/HkebZu7I8VY+1YDqTrD0YQPN7fNRUpKlEAo7jTosy3nbIcw5WawHxdDa/6
1HQpE9oKgf2x+RWmVTp83OXGsu9C8eDyhvWC43Hg2sYzXSa1KEHEsrQgI2hk
CK3oaPKucfRQjYOw8B9dygZ/ODTt/142ZYGTX1Ng5b7Z5MIohPlQlXGpf8zm
cfl5TDojJQuo5Q1ZdfbtzTE8K94muK7aKE6oAB9mjRqxXhE37kH5PxUegv/M
900XpTAKuZZpeWJ+lX4+aBuiCZLp4RZbHcZkAZxFYPyRpCWPzKU6cOd364M3
Z21jiz9J8eqcULOCq0Yx+vYDndSI/wXffUzBU55ZoLl3lsthQ7Vuia17KfQf
jpZEDAG/M91UQNfMFaoxnUYoh69LF3N29PW11oQuwsrqmOHrObyzF36sa6O9
o6H7/UqsIdFZnPm45d7mbR6+BoULR1yfk5Ixa9/7+htqjDq06uyvWz7xWs6p
M+16W6JtcWeJ7XCLOtIQB/B+WN+gyrRZAWYt7CkeiywcAsG3gQsL1p40a7c1
NVeNRZZVcFlNg76tGLKoKasgGByoyysO7PX19wQ/cIYUr0XmvUDZXFAxTW3V
5I2yFb4vFAeyrfkKQQEgHV5SKUaJ58D4Tqbcqs3kCLChuAbnxVhO2pbSRJOZ
mg6cjuwZOuQN5m8vW2DYCiPpi/z67pCnT+tyH8EetJ73CnfwZTpBRJvrl7o6
5OITB1ShMXxsqivOzR03VIqaXM7q5Bafk1T6cq38z0E8FMUlabYUJQY+pAlo
4dTVXeDUeofoLcrrcxn2ldKiKUikPjttDiIvZKbbQmM3+Rd8eM7IhvHimMI5
HNZ0HfNHVvSe/YWPlMFcE/XY9IWc9N4LnZaQ0DRzs/qCctmm6PRb4ECHH9qS
7tssIjVhB2ynUFdf35osDTyvbXmHS5jEL/DtuhaGHMBnBq2Q+kYLKFgh5lEO
HYLfjqalgLcmHw8L7C+49smBQq1tY33r1FUTO2zIC5/RlHDIhKL6bwVPjcXf
pJKZOaoPZPC0tCJ8okHJNbr5ZFFeqgv3RZh2CVwj/ib2ckiXTpuCefjhDV6Y
MOPPAiUgyfY7xM9n2VCBoNSllupAKqht2xcSL4AeLB8VWO7G31k8P5J3Dgth
eYpQjV3p3rlCtDb3qLOhAtS7ULPGVas94HO64r7zCLkkrAI57mD5hvebW1co
x/1m4o/uOWzWk7jDaBg4NugMeUllDnOIee2X7uCy1c6RPzdemXaoN8BKIAAk
PBqWdsJmhLJEteydfvVY6INXonLvLOhAuFHJHAA+DEE014YdUio5BTbQGzIR
ZEp2I4eT/0LdxsM2YkZYC4uLi8sOyy41WkmCqG/E74nzeXeyRzngxJSHJVhO
eR879GGuzjf3wChlANbhOrIv2UzqOxgqeMW3RVMgT0P+1Tv1ZXB6bF0obEjH
6kQCbJSq1T1iSoW5DTFldwZ9x0NYfsB5c+UOi9I/5Beg1jGJ7yqujn26aDtQ
yS68BYo6IVli84uMXR2OWZ+zfYTAjbgV4knWV3Fc6xjzgVctN+/3NOSoixaq
pdhlLp/xQBa+fqZ/1vNB8o1qJKHe4yhb5hwN5SF+83DyCtykCtsxo18G3rjA
C8GxNMvqezD94YSSJAWObhkNTilJCbcf64lpcdR4iltPtaA8ogAjGxYZ8AXO
QDFr92SYeIFg6rdXXyiuOG8e/FIMJALIIh0UkQcIOxn6QW/YQrm6nyUH9guH
XA+mgcMOIw5ZhDcQCnPQx2EWTnBdd24Unq2yrIIpxO+QpZvCnEEwHBWiPGDu
vqs9s3urVzAydkCqZ8PKiryMSQbb01/B5EO96M+PLptmACXsXPAYkgVDm2QH
MpAJnDUogRKLMNKBBQgUYR/jy/sM9SAJMULOwTs49UixLHPX63T7mEVcHTHx
6YJnhtTYChxWJI7QUl7aqnkTlXTnJ9OynvgjfFZfEReBKt/c4lGFV+GGCiYP
ocOF6xQh3MUXbVpeETGGiKO1xjppsOYUT2iLbnsG4zqkOzPbSacIV8IPER8J
3o8f9nSqxRrPKKXjcFhyAnlVw1Y5t81YzHQslxCJwKEAO1KoKmG5+y/lEvqG
CY4HP7ZWPtt79AKZkgeHWkSJO5rMbeaLobnIvx49A0t/xyPwMpzvrJ2ISTnE
hrpgU/xz+ffSWK04xWA6Skvp/h19NNIatea3eWL5WiPi7vVc8O62uvCjkGd5
HmX9krx6bkS9R7ms4QTVfLoflwMmG/97rRO9lM+Q/e5RofmxZBHrECPav7LU
hUWz6LQ1daFs8K+wqm34ivUy1YrNEPIlVqOP0QvEIjTFEkmHjtAYZ4TuL2Ve
ZV5oOnJol2ClnJMjK50e4LSMh6+4nWa1CS2TVz2woygoUrb/0333jUTTswut
H5G7E7Gu/hqNVO2D1/XDu3RyeLTg00/yk7GIa4JYTXFpp5h4u9Df+QeqHQB5
4i/IZqxXDgMswPhFwUKHUMMRcYgp5g+0nL1l7TP8lNAjDmZWISrAMaGtD4YC
trioLIqLACf2Ni4SBEsT6PB4a450axs9W6ktIugoERMsgNwSyjzBLYmNA4W6
Gk43t/fqasWWsUFEyFXPU872RuI/oRCRc/al60w8qwY9x/WUIrfGWbWXMwmE
TT/HR5r7ou7J4zfhZlZy3ilJQkPiHfXpzB8BICURrR/8BqGOVJfWCNMHDQ7c
zivS22UgpnUCmEIpkZgps+6m4sSgW+wTy3MbjvznAAv+GcIySQCmrOXTW8xP
p2cDT8Fu1IEdh/k8LRoBVhK0hk2NEnLdD7FjUrH6otqf6t7kNt8C05/R0Pw2
NVizUQowwTTCMp6k/as9IiQbMggaptkGLttd3QfSfBMmY3nHwImnT+l98AxW
tipQtERWeLvy7S7mnNZ//2/7uTxzgGeSTtZOrNO4h+/RJWcEHXOb+cA+S5jA
IKlMTgPEOEtrlXXKf1eU3Rnw8VOwib+GcarhBOYs6pgUBBr91w+0PfhCFSDN
eJBX2Z2p8xBvx3SCSyeoKc5ihqapObLAfL/zEhnOsq3rEhkWpC0zZ4eVy66a
QodOYOYGW9JPS94mJYwxIXSCMEzDjMQ0sS4iK4paVxZBy7SD9eI1BGHzNixf
++Uri2U1cAYy0z8b98k9NjtaVxuSd/757b4++Db/HgXC9OU/uB45b1WR2F5v
SMRLVCqEZkx5GYB1SGp2No+VFFOdxr3KaAtLdZhixxEwtHEefdbsn2ThuYaz
9M26QW8YCel2xDrC8w8jEDTaLqFgms8yQkMTGtIc3M+KfLfjg+P0cErUOuoM
HFX873iB4vaqcdQISOSqyrv7jZ42/BG3gNPi5e8BbZWBSrDesi2oq+KcHWjd
K5dl1TAIGnsCuXD/u6NtqhKWuseWgqkmDASvXYor95bf10pI06rzea+3y7p0
vMVOo9jFwWJKphgehgoyrqbwaoANBJDW+g0Q8qwF+TMdYpilGZGkgW02vt0C
CnHL4ad0bwBmabGyrZq4GqrE5phcNyP07S3DPM2lo6oPQn5IqdInWbK9WvoK
VlEpktLsRaZqyeHmAhM8I855FPwWp4z8GI9xYzBtgiwJl5OaICyTLnxOcN7G
qcwDq60gXniAt/Ncl9sbDWQo3Fc/ZP9hJzQmYHhUOqWSjBcoX78bab4zWJLs
OnRYwD9bDtIa0Afh5ufB43SS5ZrFgUwCVF1VNPDRa22WTEoZ35OD95bY30d9
nPUWjJzVHx/l3dxzLv/Jk2f8yoZRYAe0MgwdMsE7mjmBbvBev8ep47iuL5yS
CwTSlqiYvkTgrdf89e6chbYz+bba2PhhBBKKWKdJpFJrmRWrvFASCtkdhDpl
lHAkmrw9QxUkxbwSFwiMVnN/mSkLDDOoNuu8zki/mJmz7wClXIk7+gGm8ZiV
znXW0l4QXiiNuFSYukoYzU1NfZRm2g7b2+Lv4p/WNF47AbRGzh7xlCwr8vYk
RTH1iC50gpUfex5Q09jwAXx4OsgyplPItG2yEzywkDzKFMyeLkuuJUvkQSTi
wn5Kpo453dnfOMNYVz0J4PTNTT27inT8vexc3cUlnqfDhKp5ExgmX38sipUI
lM9cW8gTKzx/wn54VyCVZr2OCmPrMlzzWrWa32uw5k5YfJKH7A7y9XeaV1D4
+nHK4ig+Y41+6ZSexaOJyDWejcuzZPJw3qFQxpWXrnHQ4/WI7Kr2h74w+kOZ
1c9QXuyhtANWvUKIom8+SEX3uvSj+fICwWep8lE5KGHCRTeRmQbnns5n0797
VXsrieXtt4x6xqzIjylPWIx6jCbo9lDCTkjIFKhUsDvQQrNVBBXDgDOWo6f3
vewE4Uq/Hbpqry5HPyYUvHAunxiBMJ2hjORbTvDlPYufhDGBkNU1jfXe7rtA
3NhpR7bkP9SYu/ckxgIVJ4bKa+zzrPxCknqwqGutTzYdD/srHAJYYQVpdCT0
YQVi5Txs3Edgyp+HWK3z0CFD3yDyvlui+PEQZEREkNDWumn3PYAB1vVgnxPZ
+v3SpTkSmKTaLKo9ZiFVx8jRVK8Ah0QwB+ft3a06KJMDLrv02EhBhuUv1N4S
jJLKieUew73k1H6aB8qcCzk2SKRTyP/DskwAXE6ehfZlOV4JS/FnpoE88x3O
l9s2LtyoIyew4vPlFkcLVpn4DXgEmUYAaVFEEfG88YQuzpAaHNk8kCm48O3u
nXQuBEBCtUOn75Bi1fYOatSne22i6hUerIGQkFJEnQOGWSEBf36QBEKNL7F2
ywhIzMBbgez9qSGesWXPRccxz/CHmVGUOaZL5qbmeZECsyGN6NSNbAAeHrQr
HMEKw5+ENKx5375Zz7+FEYux5CDBdy7l8hrIcOhWn6b3g/TbDjSXZlS4o4I2
jPGmuxB0GPriAipPgnvdkao5uXk7XL3lRrIDMpTlK39fbeBt6sdeBK9aFH7d
MR13MzyyU92hm9Vs3xJ6FOh2YMnlcdE+SWHTBQt5oSpGJCjUeOT1q5gK64Nb
skUaPWwrjMJLN2jdHuEZ4tlPHOG7OKH/QI+3z+VwXBDtS5umUF7N2fgwGuEi
LzQELBMHa01YZWlrVcpK0I+zYsH9h8Sl5hVNtqDNPTTFSzTRE5WUWg/ESuFY
y3Pwb7TKEGzOdrKyOpQCCPKWmUx9UeaF83l/vbKjwLK0Re9RZtmyYTv1OqqM
rvqCQZyNo3vJxkhr00Aj58HnVe0kQtaZ3g65Zm57I2xNrpE5oKDzkKgheY5q
5w/e0tAxTGE1fwcRJ8u0Wkik7dVsOuhSI0FgQqSISrt3a/noKN3kCjozvx7G
NM77SG6fpR+S11UzHm+ab8Ss/LWryi4K765iRhkP08AZ33QdsY7GJnS60L5+
cbL45hA+ONQaB5gMgK9Mjav9ErvVTh+jxvU+RtE8m3XBTfgX1ZzGmIYTNBMv
QAWVzI2c03I8R9jKYe2VJXxPFEZN8Qzi1menSZM7ZTvmzssOUROiL0HuW6oF
EWQtOiUfLmz4vMuFO7tvoPYVr0GWkwNilhdQP8pdETle7oaNemb3Q4gxYm3I
BvJG9b+/wU/Q/J2GarzbXhQxArroVL91yPtHtNoDs5jERJr2TfYbq6l3Qpdn
7m+HAa868UlTm36LyztsK4A17cXslp6NwosP8nNzm6YVc/Q7AahutRTaM90B
KibOUfmtNaYXQ5oFeI4Mkwy/344gZiqD4RZ+mNlmWCzQVvndDoscO1ItlCpI
OH6MxYQ49so8OuSF23xWMeUvpILHYxLkT0f8r3ksRLCyZUR9KnE9thTJXol7
oJPt7qBXAZBemoBibF0bZZNYpMEGe3K/faGuBWTH8cX1cxtTbbtfbF19+7Kx
pTjxsjW5xiPaJEQNlDN3OFdaoe/p6sLlvmJjGZEvfsu38kz/r+J8y4K2zA+8
ZBKFBZlsKxcqzHDT4GBM76a/YTkdgHTng/7mCZByDiWSENQofF3tH3GFqjb3
f1KgKPCqpfhwmq3Kv3oLIPI0wKZhk9ABK8UViGmgvK/DVMxDbeSNMHBkOEWT
a3gkE6O2qq8YnXUZAyc3yVvGdesKd0T0XAzxNdWet/Y63eknyMMWrJj+Or4H
AYF7g5fR5UreaaNwNAzUKQajTAlTdSr5h2FKkOV6Eei/ilU+e/uHxFae3EA7
7hnnKZYpG/+n3SKPZCldtAs7jcQFe6cc0W4KkCi3l6AQYz/UVa2BUCih24cb
OUc3O87VciZ7oLxXRplTaV9ij7uqJLmXj1tzhPjQUhNPiMdr5dznprQZIYqY
4O4owq3Dsq32eGBNJ6ZG9cT9AEJ1C5rgcFp5GjP6xZqOJleHcRBu9DkKPcg+
TpLehS1hKOGIh/yKR+UTz2S0gvR2pZPfNBJYK91C3G0NdIEzLhYCZs2uXutO
0azcSeK5qYIIfkgSxm9DhGCpiNk9o/saJF6YgVuu930JDk4K08bMfN6KKMQL
PSfS6cecBT8z+TI5mCcma9vb1lujmmgVromQL7/kqyJbuMWUs9TWhuP9/Gcx
2+iI0vpK+uNunrbSX8p1Pfg9DYihnJxC4DMQPvW7osEvp0ga7KW02Sn7KrRD
E6+5TGMvaAsDE6hq2P6o6QSpW8v+25669K4IQML3FR095WQdls7OcNjT1zei
kL1xUM0Qg32WY3kAwu+oPdd/Dc07rWQ5IL1I3IhWZOiHeXr1JEuJ4K9WVUth
g6cMX6dmOgACitI+NmzSg56EKWmZ2sGrMAwBRTkKlvDwNYpoUls/DuFvHNbZ
ofgRx7w50WlbGSAPgLQ8Gg51GQZuyyMj1mgrJlKNK0F0XGBk1ybyp8kmRZnv
K6Mz3YxPflKS7B2SKg1NneZdROQjOFD8yPZAMozs9qaOencdjiCoq3JvKPe7
CbFa5NYx7jyaDJxrdPC7XGF70fFfLS5YwqYlRr5JtUs1H/ONeeDd6jCLo4xn
eYS3DADppyL0V8CfH9VRfHZt4CHtHgcrF5xBjhykekXZe8SjodiArroxdsZo
O+Clh5bxkQNuDIRCmo+6hng15emh/9TloXgXghTVqoypTAtcJGrfMdezf8aU
576STySUjoDsY7CDT8/ZLYeswirB7e1Fj+h0VMsH7r2lD6dKUi+zp063TozD
VbZxwaktiEFVrqKOlUUOPaIDkm4fq4paUd/ocR7EyRJD2dH8bYDLpsE0yuwt
7zJW2xjCFBY9vhKT54hNpUh/oIo41NvRiq9LDA1Inr/5EcMK0ftLertA8+Mf
Mv0dZCZ5c65mz0XqOXFef6YuRSusoI3vZSfNk4z+ncZq5YOIo3C/t5eriCnH
ZnDD/J5z1B75LaZ/NKXH3tl00YqYpCUwGmVnfecL9e8u+ck/DiuR7BGSyAFU
dKJMbu6N7L3h+mtznoPvrRTZyn+Buc3vFIiQtnmP0AG6FWA7WT1jhtGWEPIs
0wgXkMI+bVRid0hjE8bKRlvEDPlEKzO2Fo0icgFUiRE3/b0h6fe5ZYoLxfO8
u2fdzxegs+WKuTsOR9LPP4sOcZh5WFFCoBlLdoRH+0wnW3e4UF5ptXhvd0WU
KZTE363rAmellEMHEUxBLA0ZLLEKq9VZb1GgpaG8IUbIGUjKUAipcSHRdjl2
DUbQKOC9dqQhDGNGRey7a7e0Il/hVhFUfUQF+1+g7a39mXNdv5Pz4KLDLxvG
T59HhMV+vkZD24BkUL5shaOcK4EJ2ihdADBVLuKgMdSssfuWmSN5VRJCAPiu
ux7rGoRXqfIxlxyEYKs0jZu6jkkaWV47xrFKQNiA6tK1W6hgiUEePR7/4j3Z
VXBupWdEKohc/2UWYgcpvgB9kzNvpUXR+0n1H2xWKkWOArGUjSm5LJKv5331
StXLFSqb474ZKj3PR/k2vneqAm0uQ2Hai8mOs7pqP/mToxm6Nv7NH8j//prb
FDxBCgRCjuFT0d4q4FuBO9M7ZRSwxB9XrbvcAX/dRA0RSX/znhhk5ANeT25y
oqsOweiwxASeKDliUWuDHgN+R8DbUZrYXFdlzNMmZqdkPPevy/mMWzUzdSlQ
c2WRYuUcFdNUhUbmi+c4uQFaSnNMclmUSmYxq1E8AUTUsCvugH6TCYW4DEIV
6OkOnGUKTjJ3Lv58toQCnaSWKJI5psKw7e2WJMt+4T/HWLqfxP2P/QIt7mqs
1uT8u6JYIJvMrX3fxspLIrml2QX7UnkWWCmPwhepTu7mucSNfjXt2h9hu+T0
yh/ChAOJTVSgWS5IUrNVsZvQmh2XK65VvqiQFZhktV+hKZ75ozFkZcHbMRoO
25kmkIwoy4Yk6VyQYF3pxu6ZuwYX2AZQRGrhrYSFFydoBUlA8v8zGGF0f+id
XcgEV9ncLmJIHxHQ3xfqBDsNuSXEyG7vqnniGWClWJLFnqx+bsAcJLtVsXVa
i6UjQw3pSVTyaRC47kyTnqctNFRz1VLrm2ZtOr2uyXjvSp2iw3KeEHJLqO8w
jsPu59p2IG3WjmLx6KqXUsVeEUNcCqvCVzIWPyLIgYwijI2p2kaMDVazgFou
eNpJWMUoAYk+Xvf4sM0RyQuIkADHFHRw7AG4bAnu+4GQ9Hp3YPAOSl/dbDE7
5mnyS5mT+IZpO5ubSOli3nHnc63xaP5TU0mvWDQ6HeeVPJK/Ika61a7b8k57
z0HwEa+j03c0cMylMMVvwLnvDriXpjdEWqxLJD2k2/ovmlptkeUSeNEGWycB
Qr/Sc063g1KNJnzjnP8L5IEcXVY3ZbnsZSMBJnp06pGhRjKf2xb1sZlvu5uo
BQvxysf7OgizSw5xSAzkDlu/Z9MuL/u7kyR1GlStIw58GWesaGej65oFQn1m
OdB7IedtKq3ZiRROAa+Qpw4wvGQ6rYq2qtHpWGn+aBRJj86iupNlH1i4+5Ti
U8WzyRf1ld5gtis5HN8nlX/7IlKgV3toZsvNcTt9NV8yrwhYH2KigJggRTAz
NO9IIZJg64zO5L3TealFzX9CCIs25RkKTymxyGJy2vVOxWLsrBZrHoIeoFh9
YUIfxTY01jx8M92pZ2kmn3ooCbvWYvsAUJFtXkH8RMUX1lXeEKOQfdI9tSOV
U9qugpeeKQP8i7XVjIdWhHLqkq3hg57PQjd2IUivqPaa52yZ3sCGfIb4Jkua
TInnvps0uMFu0YWdzWdJikWJXyZNPmnyU1IkKmp3hHCV0yM5/2waLBzplLzG
SHMEY8WFGxiEMiZQ7Vz3nUwxXn8r4uh/Wy9ru0NhyG57eycNDNRF11XjTb4u
z5B9brCaDI7qJID+BMd4g4P3LRblwnNYikzH3mxTQaiWtAwwwE+jtZcJnJFj
QzBB0xILT9gkTXAJFdOiYQwpRhe1GyvGl4l5Acn9Cc0jge8E9V/u/AhxZQnx
QlQxHySjbOXVbhJWag5tyhOuMZ6DJPQ9qsNdnGehqb8VCtFQyi4/sEA0Iiuy
+mqT8ogoARIJ/zuistgE9vYlWG9E1Y0riMg8nQIzohi9Uu2AC8LU2cyexri4
kSYneiZQRdnoig9Tf/N8dpGZMii77MRaZb5lHvd4VGftk1mdDlc62VJWeGnd
sbO5TOQxVkKS61Lwiq3zUxtCg0PDzAUUl8Pkk1PfPqj+cPOSHYS4dct3XI64
DkXtrbt5sTtgtoNaClNCh4JA16QR+D4kLjsiB63qojpwfE/bbe8dxdr+zBkG
3P/tyoaBF2/1JNHXHBfddnethJ+EUGynzKMEjMsUsEFz7gcc4K5VkWxM8nZ+
/Gslli/RNqs0tuU5F/0KQgQiFmR1fXUnSvaiQxZqMQcxZpTeaBneOoZ7wwSr
dGg8NLpE7QdTri/Kx9E+bgmpFQ3YRx/WFCR95ovg85kU5k7OZ/jA/nUeId1l
2gf+o3ED44VcH1c8EtXPGCyFvnRp1qm1JYIP2TIdmUKpu3DeCq7yCBIHg4U0
rH8sdRoLYRXu7MmPQzj6tuNL7Q+PerCjkoQt25Qz4jUU8e2M5IUYyKFzLQEF
y2U8l0ZEfI3Owk/sfa9uLmwKg0f2PWBWENYA6GzZshibrKC3Zef7vNvk8pkZ
Tt6GJ7+NH6Pesu9KpgNEk6OCrovqjmKvO0CwuNLd+Zv+Zx1L07xn6jMk5L23
PBsgLyFTYSyEPCjpiq6qWEI3QhE94TRqDqruNzhWSr9Wh2IAGs9uiHTdyqqp
het4j49cWHoYk2pq+QKw976yr2ZBg7tSZlAE2iwftX4stiGEIpWVuWJztmTD
+envlrCmFxegQitp8Zj471gdc+WR7VHrKIBOqEvcO3eVHosojZamDUKDW1M7
0+fubjo3uE9xixcIScWDcvi55GknabUIZTYqbxMeadN0E/GD7otFUR9tzU5+
OFg2plIYJsc2IrHCyH4ob3nkLxZTON8rM7F6olr2EpsfHJZK9bcmgltT76cW
meY8nB+SMvJHOJDXw8En84/S1aFhvaA6syAnnpkStZ45F762UY7niqZ6y/zD
5w4csJSiD9JiIl425LjVQK1pnowXcvwqa73Breo7ZMMOQlxOjUEbYuBYCyFE
0O/zdHTAsbMYMdUVnWobJP3k0YOz2CXZb+b73dMiQ93bl3ioVOXe20XDMl04
ViJWh6t/VHqlEnMgEKXgdn0kSMDa1jvF3vbnz+vle1P9jnDQfsSexTIjZ2Cp
ZlpSGYoJFwfwTLHktSbckhKO1NFMVsDuE3i1NuPySuns8IhEhoWTCXr1RgFZ
yyAzzHV33uPmKlxmp6nyg624Gj96GPU6hPyawfgj7b2DBl75wm28cUID/XUU
vUXqi3E/CvYbHO4oth+a5E1cj4Bhn+tMA7Jat4+2HU8rsarFNm4qBsf9+6XH
4sAzBXAe4Kv/TMQ2GRjZnzW0ScojU1MLrtE8atg7SVdSjlgrmfFa9uGBfRFY
tljTmzYGW2eAdpB+NMatVQ+0coOVL5A5hH5SNvd2xsdCzIDsazkPqRebACMI
YyY6+iTnmDSRSQdzlmIQT6ru98eM8lbK2ao+8QbwIdNSf2Rk5IavJeTIqTkJ
xpI6hBP3DWgeuj/MQP4d8JMPy0bdwRswKe/RyPxgdx2Gdme3bk4eLMZLpX4M
DY2F4TvId2RSrCCuH6EVAtxNq5/tfvXMqbA4EPI0lwNsVxT4QsIseTcQgIzA
oZuzffM5VlUEiE7icTuV4NG+vdSlRj6kSclYqHFW8ljm6BiUVGka7KnZ2M11
VWTVpsXJ1DpIyMxGjYANveMNB5hkqs4Xj8B+VlXGYD8P0j5bHJ8vwzIAiuwG
Yl0KNFDT9sj6ctbmz9v+8GMs+AbPFw/rp3ddImsE5TIbTOlTdVIKZFRvSML4
YAz05Yl/3r2qs37SPnbb9eFQVC0FMAYUdwJgzE1zUerZiH1UpADKi5qDj9mm
eKnP1izURG1q+pLbdeUmfl6HLgtz372D6/XHuAJ7J6rRkbqv3cQO9mfvaFfS
T4ql8gVTNx65OpCtlTZLjp8RcqiiqQa2x26p0+LRYVJo6119ZTYS0eWJPdIZ
fuw9LH+mS0FCaKqjsorS9LwWeqtJ3PUhHv65nn0sK+fVLHfuoeH62OwCwexz
pewOa6e0hV9hr+1wqEoMdz5FaPjlO74zmv/V4nfE+2cKrgjA3J9eBIr5OT1U
Unn5s1Chy2UFpG+N0Bx07ohafnxs8U2qzA7pcvMZawRri71Mw7Vl1gcBfyne
4IdvoiNLAMBy/EjAdXV65cO2DZAXdoMhgC/Nv3qKMxlkTT6eDl6f0Nw+daXK
mMJc34Rlyt8J05ktlSTbsvMrIK0PHcuXEFMghmulaDx4or9gNPu5XrDKp2Kb
yIK3nxMZeViep1Sbq4WIn8DbMW3PjrEgo/gUgPauTQ5HBFAaFXvrsvjNUXY2
xs/v27J2PTzgfLgHzfNczU9KqGzsCmkvP35hASqM2FIq/wMlY3OZo3SmHsOo
U7xt3GojqyMIkb86rvDwhqhfNkDAFUpl7xwKweva/9Ch5LG+pJx9UEDguhzG
I/vx9i/hpxTe+bMcUDpMUvcsOzXRzmpVcaytgVmYJMocM1tcnOaZ6DkUha9b
9/W2UfhqlUX9tj5/ppaFfv/ySN9tBLajs6fpTunyWw0iXbr0EpUa/3H79fBJ
ld/Ac9kbMA76UKPSfp1yo9RapsYOnlKXedNV9IYYofrfOLDp9B2JkanFjkms
9y5yWLhj7d5l4taF2ruey5E3BYym89t43R5ZE8OmL9K4xhMbqVfrhMYW5QYu
lVw7ndVkvYNhk7FxA4HgvDA10ktKYQI86u8eeXrkln+EbYzdyIbfnyGwEWEV
atkBGiiz+X8nZVlJkZ5rRBDNKeO+XMcS110pSYkLoplvu8lKzHncY0MaCeyg
eBjGBDfHEmYtB+1Uxo/26ztlhhfftvZSNKP4CRJ2yLlt1lf+NYVykyEAoj1E
JB6+1CSKEvG6nGDQG8k7x5W7AHZFYiyRs+Vdi3zut2qDqR8X9hn/zBhUsVaO
UgkYuS5UzPEkbCxUBwileGmH5Y6WBOOg6BtG0fndgIwHecHxn9yxQ3PPUOOv
Ywokhsu/clWXXfpbW+07HmTFfHabhrF7xfdL3IkgDJpZ/CoN/cemmxAAQixe
BkdIjofDfTpvr/AhPjGn3m1HwW/VNm2a0euSklQjrY6y1QbTg6BaS92y7XBn
wJEyj9YLMUHDkm7W7TmNlys33BqcLMGeZiK9cyPd5YfcOIJL5wU+twwPIMXW
nN3QZ/JZU/+0jj8ssOeQRMawr3mBixh62hnq9Dof+xhuY/n2gP5gL0FUEBAc
wSRtei0+erwW1CGiEVfwIhWGN8FfQ/aFEELchgfI7/euIaeS10H9r2ZkfnmU
tWEhYc5nGxWXzFCq4fQryH9ufT8sLfE1huQV48hSQGZSxVVpBfhl+MldJ6/k
qy9JF7upGs7jiKYdxf2DniK1MpUnY32nEnoaX3prNrmF/C5LBuaCIGQt497Q
inSPyIIqEC+JlELlYcfavcSfp52qckBiJAeSFStE/ChFP1UfCAjrBJC7BqDQ
DhIYLzbkM7hqggViqD4ARJo4/TOzQ90w58fyVHbIlczN6Zx6RVuiBUw9CTKi
2dUXCrqtACxlenSaAG/UJ44N8wSgdolUMHSF0UV8FOB8vB0kBfNVt251wF20
qNygx86rZ71sURumgNUG1OxzZTwBV9h4FYo1SN2V4/ariO+OZnsRmojfkJn3
u1OwjJGM0aw/9N+qviKko9ujtKLU5IuqhavqzZ7h7yaWUjFNr2lCx9ZdNV/R
X1pUvWn+P30wj7DETbXZpWWnlDa6SJl5pN0Vk8VzDMNrSGMU0I3ZzTjQgtbj
yur3Hrd5b5QqWwhe97FI1c/l91d7aLRsU9MyYTKw/uMzUa2LzQJ1RmoYielW
dNzZeXr+f2g0NPyhSemUfR0vH4SQf2zQZn6v/e3rcHNlV2UFUGj3ZOf/j/eZ
wvG+lsZPySNnOMngDFUTW/cNvYWF68X5/7rlJ+1puGDrolhWVF9YRz8scDaW
nWA5JCB6w/H4eVsuXjTRRvaFN87CCNN8cBU3e/70zzvxXEN3eENmA7OUiiiz
uczJ5U4KwMJSTk+NAGfqMwTr9w+Q8R7YqC1WPdTx/RFZVscdshDY8E+kIRN8
VDYvxiiBBcG0KC3l1p7KnT+xzqdD5HszgNvzFWJBHOaBJvTZLNFVnGqmsSwO
dv7Nvl78R09Pm1LT4nXWnhVX93LsG2Gj4CKA/wbR93VLJ+Jwuzx6/0IiEfJq
Z7E+F7ShuGp4E6Y2fyExTWk/lNXlBJjuz0I9eeu3i2A7c9Dg76AlPrOt4kTH
8cRvyZpN8GBdPHBHNh8bM9CT3ShihOkMC5KnXOYOy0PSsw3QPNUNCeVE9ZxI
goebmKKLrxDdevUSaerhXINcLM5QBZZX3bNm3v+VkK9OooK4AcHK95PSrhuS
eB2+S1S7c9O9ZLYj6XKbFavSPnhpxVYG07jFcj8oTi/e13U9m1QJtA8+Ve7x
3Gow0WZImtmEBkuz/Lek6rRNGgHIXn96hcIl5Pcq7rJO/TFhR/YEM9FhpZzz
BmxyH40rwAQAd1BI/ZsF1pVgZR7U/r7KLbAN+hyiwszWFBzZKtOkpMY8HhCo
T/7uRLJohi4T+ETyhVFY1yUWHHkW4SuJKh1Uw7aBRtzwrFFajunJOuGafQ6C
AHFcZzBRnleRAxusiIdx3HAlDslNAahrw9f7c94z7gwH+xAJ5/rREvXeKXXj
4VHGhTlPcrnQtikxItLqQnpo3qbnvflCU5UF7BTbMtqHHIkuJOd4pQw53L0/
N4aUa4ZpjXMG2iWmoVOOtOyErc8ILi3gVPn7S3Hq96qbXn5FrDPVDv7l7mxM
r4CbQeAQiLqeabEir6L3l+Y2Uq6jvhJE9TRmfP4h484MRUGgHoejyJ/xwyES
tkOKzZTQ7whtF/gPTVvsZ4kTZbt8IdfAclwmfwMBS8LO4s3G4QAD++3Ta2DZ
ePq048Eej8SBCjVdYdxn1q20oJ375Yhut6LdZqAxj4XT7b6F0mI8pQ3q/7SS
ohNdyoFu8F43sfTmBR9rovVdYHAuvTd8ocFiPiojSqj3srJ9WjmjXivpOiTd
tO1ZSVOOemRSeXDX2CMfGPnmqiCIFQ7fHFtroP0D2HfaFxiC7EzaKJmjhzzW
wM87CWDG0MfNo5Lhv6n6/BKnHja4IsKbCfcoRHmObQgMpUskAVYsWqNUUq1W
M7CuytDJK1gEWt4E7lJD5f4K6qk3TXGy3GJosX2WGHl8kaAqYb4fKmoKfV7I
GuWtfbwpnjF2lJ8k1TjeaWGs+lYP0+AB7AzorU02K/I/rrONgtB/F1/PCTT6
SfJ/NQc+xzwywyD5Xxy/ZyE9uTRz8CBWd3dZWzYQ7wOru4B6GH2a9C00vT/p
9XbfBUh5Ao9CasI17yEkppFUoB3N4yoNqI/Bg74BCkqG2KCg/rJsr2pNW46N
ZHeP6Zo1QquC3Rm2mldPYUiZn9pWm1JqF18+DpJp21TR0eXRjhlRyf7AStHN
rK0MZdXbSrKYK1V8bawDgqH+fMdAOT79gi8dNxWoq/RHQkcTP+7KWXu47Wnp
3XwDs2IaWoydSNgRXQKAj9WQD8aVTokQXPvCV70+8ImIYM8no5kS5vwUIu1p
yIqT8nxkxb8rbwMFoe3q2+vnYAqU/aPk7TdS+ZyxCZplY/Q5jKYvjKzSQjEU
7T6pqBWpblroiYyZwbFcsXUFou1zbV2EyUlmkNG+dIkkjHZkWRObEbVoq6vY
YflHdgHPdGDjOAhDFLHWxBCYExD5sU6c9m15NYlkZsrtXc2MfxJb08pF9aLB
SY+n/s6tnInXGhOQqlL+VzVPC+T7itT3lzjZWZyzb7rTUOiC+igWr+dkhLsB
iLZ3t354KS3Q6+hbKu0LiqYIetzXjE846KaSfEoRC0ImPGPsSc1ZbUKVhBbo
hj8QqXZH8NLFNBDI6klMJHPSp7hZbF2HTVoEMM2MzkSO2GIVTfEPxoZHKQqW
PcBCgiv05BKc0cCtahnIyburvOURVSZov24DAX6MPQjj9lotSlz9wHeAlg4a
tleo/sGsJ4yHM7DblWp1ucSfULYviTdEWr6HzPmbB8YFpkdSpBE4sDgX6UJW
3dWAQUvylbI4Ev+E8pP5LL/bJiqq20UVyYMPfZGFL7Rky/KTPwP6Ev6px5jt
Q2X6Vvw9e5RewfiyQGmu1GZi6rO8dzL7l9IPwqFKRYoLZPmWtQ/We7Mwe2I9
Wq6tJ299DEqNPI/KNtKTDiVEQoCDJY2ao+CBMHLbU0RVvV+Ss2PILVNudrpU
ZqbXdbKu53rTJcZ7B9kxkTdhfYTyfqRI6NZnAndVHomKH9Zd7iGhKYSoPPeA
Pfb2AZTyo1J/ATXD/7pJ5H8kEkxRrhz4msX2guUopeR+JNYY93v6zr0GP6ZR
Za97QGHmTk0Dzy0JicNuBk0YdnLD17mh9y06EbAbBP/Vz69hHfpHeHFBZgny
lA8Ekvidci/rLmsEFLZm0RCMFX0F2oaw9SzrTaiHIDFGQGCbetaPkQiya6JX
KvNYQNYPKUo6gzF2TuLb3vGs+5w8eZoL3/f14MCMuho8RhIpjmrUgWH1Ue6n
0GFppFT/u8lkob5NP4SoCRRN6aXXT/eXjGDN0xqRZUcvU2PEVgBtQ7KMPf9o
IEC657MHWvh0HD4+uzxx9eRC8UkU4J4izZssU+LKrChRrXK15F2lXUwerXuW
R06xgX4qF/TAGlRvAYVAem0hQ2cK/wyADg25fs72aVZvbpv2xHBPW/ptVCnF
FQniJBeXZ/xVRNLeNiyAbXGkSeHtJlSvhDLVyP2VK2pa4LLrDRgpRdnk97wo
rYWF/MQId2h1hTSBTz+EhruvjcxE769Od9dl7IjBKuFkrsaUdgUs/jfetjhM
rAn5YE/XNZggzJ73GPFKap8UFVwyUmy/hKhAteCHpy0vhIoL9+5iRNLCwnZJ
GjW8Izjf7raIP4btWFEs+KBZBB2Ae3fkcH7Ie08IdLz0eptq9wU4FJPIQyTz
X8AvP11yI+nWuuj49jil3ZEov98LpLa7efX40r5HujA6+nBARVAcaxy8FjjH
fZTbf4y3IllB8xlNNhBlitI3azjKXOiScgUek0lhXRIJGE0QLVB3lcN1Oeum
wnveTqcooSBXcN+167Fqa4A1yfXQixUtneIAt0nj0zIa0YDd6p/VDCL0N9UC
lMzDQ+sgfv/b9owR+fDILNWdxDNw3kPlYxPm0P5w0KUPdjeuPdbakCBl9Axj
iSw/OH0EwK0+rwx38edGHoXphHoDlcrXk+ClGg+8lvQe1T63XIxABpi5ugL3
rfUCHijjBH3W/rYHw4ePo7aHeeOImbxjMxIDywZIVU/5GaeGz+HevgWya3t2
gNZA9WgLf4ykNjtPrA8BAqbABJpY5iNGc5uU1QYzR4o4k3kxD86S/tDnQSB8
ohGdW6VbH7BNvoBJj3dTNsBWytyHojabSjwpiYXb53/6bj/EpfZLcZbPZgeS
p/IzhS7+WDSbL5GB5Kn7nwwQCV6ozicKyEhJdv0ydpWynEL69aTkQPBNstTA
ybawn1b6eF6c8qhqN8moK9imSJp3cNBgoJjxpWrclnjp7XsB2zy5ohWqjwJQ
JGXBo31F8CIqDLYzqKDo1PSDw/qs1ZVjjDOod3W+jDKSD36Df2qckNMU5svU
h11QRrd0jD/D24KB66f/PTS3cXiVtBxG6SXZnL8Yx3ZDPDHK/OgqIaToNuHK
uQPcGtNsTYljtElBX7KvtctGJUQ6On7HaEbjh3R2MGnu63gfRGX5ktTHq3rg
GuSIz4v7a/FgQoYP/QQlTHdbReqHgEI4PCGbNhE2cbRrLJXvpxxgI/8F6OyP
RnQY9P+pBWq812iZszpbcO/g/sJS/qoivIFFHiMFKSOAFYgviDTFJQeBCPaU
ky+p120hvHnKJ3hWtq0rXFtPwUTMFRqrzV8CzQibAxFcuU8unq12I0oGTZxe
AKcbDczyeIbmWwYYjCQ3iVEzpOs4nMJ38c7ZpBp6MSYNJUSKlw7ZPwRJk8uU
XGZX3prrRSUfc7TFiXMpLNZezL/sLPLkBEVHR+XKLphSD9gavaZAFGd8vHtW
FnIrO3dD6xYjLwNplscxXRYAeKcrSIvTNpoQZQpFtDC8kXQE61MTu/Cutl4R
eBtMhHfYATHe3D1cFxIHjRxJ72p/zHf9K0QOwibypWHPZDgHGUMX0qycGSfH
U1g+yFVE9bJIRQJ74jL1jS9CsKLkC2CQSGQpA/FVtV+rU7lYoGvGE2/hSrnK
ZnPF8hZWqlToKZnIVb5uMGgB170q2ygZpYtc/zbkhi95DKgV8rCOlKI6eQou
iQ+pwiOqaGVEX3ZmlrjsrVMwpsSwjgJiIa4y/sreImwEtYW/gJSX2T2DdJyN
J4SW9INjdG0scBzyw7rw6xfqQ9a1fzrQTUAQypn3+V07HPnHDOnw66Ppnni9
FzscBEbDGx8i5DG0qz0+6uwSHKOna71iaY+CeEKb5lcDydrdbjJWektOCnF+
eWO623QReanl6eG11PEjhPXRrTVNL3q+BX3Dr3u9MIUp1DJTAzo7Rkczsx9t
SDTW9NliQxWbLOLJ3s1+STTHd7szFFk3GL9ojgkUswrzcc8Q7wfXLF7/z2nB
wdmNdV17jbf17j32PPvF4UBtlpGqiboRENSMs6NCpdPul/nXxY1aSjI9aPfC
xyq5Bm7YhPiNdHtddQWP2U86G9I20qjYb/Tus8X7GppUX3iOf0zjMHZBbXJ+
BK+Qlt0wm20uV1earuT+9YLbyLbAgmTnZnGude7ijdXYmR0ZHHc3F6YotxVN
+5hMcHYPkcXtfN8EMEfjZratu0udeJujBJ0hOoMZlGbPyFJO7senJgpGZukh
xRC1W9lmlvRnpERavdJzxcbczheQl7ayjkRAL4H0iXGAnbp5fARQeaTRuLr+
GQaXFDrn6+W5RJXwyi2b/v9vddb1WUyvjSmh2T2rlx0x6xO55uKIQiItGBYK
QoIbyI2hE6Xq6ehER1BTasi80laRuF6vQLOse37WzAFuwJQSAjBG5RpJXNBq
yL9NnpeNgOd6r0JvRoNxRRZncneGUOINaO5nodKfOKMeTnNeg3Ej9AcLCbBI
HvCWXxqslZMBlPLYrcMl5F3lc+mfCLGMFdji9XuRh9UOelYyPTb0o3kC7Rpr
AaI3dRUyuRryeEf6frY+lrmYuI23GP01PT03BGsfG2R3WOaPe52VL2R2adjv
IFyTMlDMe507MkPUGhiOZYu4LdXn9cx+9Q3JEtDWUGyjFULi3tynK+P1vDoV
WPxQjDM35tkFT4WAgenY7OF6ZPwyUJeDPYqoFiRDx0PseLnn36sBbA+wMPHX
Bi8NTv21igLBWDC5JteU+OdNbUB2AmukJnnd/lSB9xJalnOMOf9WHzGFR1lZ
4u2Kljc/04O/cGM1WpBGjIzLgkRlqsykyE7YTUccgcxRH08fKQ4O/lczJgqc
PPOSCLy2IWWCvtbOg6VMAGNofwuxTjC03LsfvYK3C6nc8o1f/EspQyMW5WCc
AQeiosCbGCnsKO0a2qrkSCUtUb7XYZQ5eIhEOvVhO7C5u88Hu/Y+dMfH0/QN
IWlNapzrbrAUGcp7kRuImvrvc8gMNhhBII6tpRIPidstWyuguWZ5YcrghpDD
wnxZclSKSomZNjNYj/oLcNnqWu+zyoGoiVY5V1cCMg7Wqiwap3TaoVark0yI
gCV4N72qDMxO07sTgo/YdmQxFGB1WF8OtysfEaWMIxQXsL4rVPd5ypil6GMF
XNxMwPDAzZ65mUqIruNj4JwuIl4ktttViw8z4/ouYiBvH3/0/zMqH+QUBlsI
KmPbjHa/Zfh8OPiLpKAAj0P0rfqmWLOGjLgjIXMEEKih0bxCoD1svTnliLnf
DY1tZkVo/jEM6OjxQqw8uYssJ0bSkW+ZqSddZnppXMLEFEzMUM6Li+YBsPdu
BYwGviTZJWP5SxWTo8BZvPgHVAH5QOqER1ULf77Gc/2R/pHsB5imYa/PG9St
k9b0hcdvjebQRi2jrvS2umnaJvQoEqza5vB/nmzqyRyOB1ZtttzVyfoU11EK
cPY+ogANAv0Lu69xYxAo7imMx9EwRUNU41aRfEEAO4dhs4Jl4xurw3g293tk
4Zr6QzbKdmrhOA4OAfw8QDGTukzCcLT83E6OOdPSggAMolX+VXKEIQDa50B5
i+PsEfUnIaibZMxFWkov/3f1u8tSe7+kDGrX/GojH63Gn6KUZd052REgz7PI
diuDcB1F8qcBJ/hOWATorpgNJN86/RlUiI7OlZc55Yqg+/pb/YJ5nHzq+Yyw
PYalvKhN7ZKucXnmFCgRRxyJpb676fm1DxpBxtOL/MZmRvPLCvd0VKUevPvy
DTxdy9owVOd9VIoAOBD/5qlHxG/qPDeBnz9JkjyRdKIX7HSosHsRs46ZqW3f
PZZ3NiL52+HkiOhTIMhXKGFHOworEnkd85MdsBxAEVxHGodSYt3rAoNUqCT8
DdDXrIHzjlYGo5TB+GfpyIttWEkb5/aIgRyBJHVF6zHwciCo6+fimWqcBEvT
/s+iXpd118wVHQBtLxosIMYRwsXe3mkkPNqOZXOSxUdZBjnNp5Dh0dEoBpQM
t06L5ux/6+ZSqW10inWJ78Xvaav2uOEjNACEcrhk7iB3+PPBFZJuvX25TVZy
HtqY7GB7BTzFZndrCjeKjz+mYeZ/29GdJDooXsm007DOHzzRVwp5638wS0BE
EAnoSK2INws1T615Daq8vu4NsiobuhZkw5p2srzF4QQJQd7KWW7SWcpZaLGl
MPn9cFQEv28IIi2iK39CrulO9mkQLTOwF3smmxYPhjbU0iNRoQsltTMJmy0O
zQrgjN9O9W67lwg0JdhHIXKKCbydiezZzyV11tpNeP2FduXV04TtbBG0aGv/
i+Jsvzu/rLfN6W0RDrPcayxQetc2YD40wob2oirG4zC37Ip4y3z4qky0ABut
7QhR7aaycCJlYC3ZR4UaYvnhUC7IWLoqfOZUsNk9DMMZYm5BtzyHFczZeDzy
nP3J46PLD+A+kyiRiMb+oM82XSXREnXoE2ertLGmubBihpW2aBSmHwePagg+
IDFC6iQjb45OnDs8ASCDblzYHpuzPJMUyvVHxX3RekGNFm0auZ0CDUfBMGOa
3NaxSD3R/+G0zoEQ/+SgtW8cwkhnnehka/I/pQ/bazqEiiYXuMsFzbgTr+YV
blPFslm6y8ZdsVrPlDaLgDZjKuXoailG099GbelJDmgPH/PtWSxwh8QX/KwL
HWXv5Ns006RwW1x3ORmFvyjMuxnsOIRKdu+HHIgsnuRDtaM8bTgAVyOfIBh/
hg6k5ONKYgdWwU+sNVkI4m1DDKPSu5GXrUR6gC3wSQaWq0QnolLqSWicwG9j
/oeRGh8liQeu87eSwaX6eR56XfS41gJLgRu7qsIc2+nxdaPbKal+LX4ADHYp
DVeRvwSFL/geYRJ2MPUR/O3ldlNNTVIZtoSFKeEDQSCNT7ef5pWUa/sUisas
ohfeYyfZ2R8ofy6N98lQPd2bvbuEVtRdSRcw08KRwJ7WD8PvdgDUn8HeOsqe
J4GLW6QEcbIh8xtsfSYqJFr2YNgNSTCGEoB+LUKBGD3nYOkchE+U+CxIUDJ4
aQ51hF6l3enN+rot/JAqlcDDWeecFWSnVoemAY1iPFBYgUH1+SjpFVFzR066
Ij1+EGTnSHscgBxqgdt2YRGfDn/fxO7jK3Fy2dIOVrUrX+kssaMltRyAnCVw
hoaeI1vfjpt5yrIbj1ehOCHWiAdf9QvPa0jA48EgJlXfWtcnFsLvK2gQCz9p
EXsHWhca6c0FS4KUeEdiNmiOBg7CaRCJFy9fXWSYPpwfH74hViQrXOBUSDpx
ZmcbAsCMWXGCezhE3V1L25XZ+u3xwV1XwXdLdCznWjdKwcwclzIYC2q3o+QY
PDdNcvxFRGGm7vi7noyOp79k0XMdYJe7n/V7bGE3k8Nloz3IpI05sLZMJkLe
UthmXDA3QfCxCo4ih5DLlMpAzCQnfNQBzXZhYHc9V27hXclyhNP7o/b4cAhB
qh1QleF0tcrWXaTW3iaQNWmi13NfnjAxSaALmhoMuRWxY9O+o5rjDbH9ijfz
sD66oGq9e9aNtSWX3beTATN959+etXUA0AwoO+8nP0o7sen5mrYlL/UbUg7X
O53Eyi1V2UUDqG2fYjCOzMqdlewSXNoNMM1ejshjNwUTjEXA9NG+pgdhCVlM
FJ2PvSMqDKxn1KSyta1ce859Pg9R5+znBhto7QbO6Ji7hm6SocfJjla6DGA8
4cX78pVhXqn4NxcN0cJ1/u1TwBJAyTLPRPUZZiLWfKpjwp8tOldvZNnqYsOe
wcbQDn+zcApmktCGOZ4/3yLZMWj+RkOoBlWIlRWc3anaZtePRHiiHdMLGJzK
DbKHPGtZzfyFYDasfARpzpz6k7F0sVTLPnH2qxVe815OtXxejgbpRLK2/Jhp
QeQgPRzsq+8TPd9vc+toKFo8qNBMyXw0FFEleP97jw0Ix2JVrAhBUKwWnT7X
zUIyzG8JmKPjdCo08j1y5kH1ilnjgGu7cFpiZyXkV/xWju9jEyQom+glLYYy
RPdWnEz6AfU6BLBWPKWa6Z357PDWGXnJoac0tFNZ5I18Ah9Dt0yhtO6Qcgca
Zu8wOSS76a2BZ6iHZYZm6pMV8KoYyWZFYYrkrlDhaxNasGjtbRqz7J1oHMoJ
2//hS+j0Q7oXVuQqpOf8kSq3Gr3lYD5R9xHEAvqOXQuwusoApgIwZ/VBN1PX
ldVu+1Hw/JLZwWSBI1aYQReYrt3YIh23+kRMlWLbelLKg/eSvPkSVb7NDdBT
uGy9KbTnPZn+Y/AUCPqWqS9fLx1HMcQUiwbKkrJN4szuBTZZu8kTLth6w4AF
Nsu7aaQcmW3MDKODyraA95hnVfUtm6mjnA6h2+HRNPznVvpAiTWV21ARpdyB
tv46OyZoEkwS1NoqxVm7mGCsnU+B8ZXGTRr39UTcgj/mtT3vy+QsOUgva5OF
TNZy+pNcQCqI7AJ0s9FfwmEzYle1VetuHUon7REcUTGJRjIdwxWsIWjxpPuf
1aXO2Gox19KM6EwWRGAMaygVY6WSf9acVXWxvGqCYEN4h2R9N8X8S+ibfbK/
JjPFSGQzmacORGTAtx3wvI0MZcFT+YbJJWMDuTwXojlB1PVocR8P1HK0wIFg
Q5SU3YZmg969Nn+C/qT0skHwgVwGralGmlH/WccLZn+fkr6oG9oX7eRMjldA
XgEZmyJ72EnKq6agXxOywvSMjCFK32yZeAPm5TSxhoP84iDcO8CgdfCQ/YPA
AghjNBacyPVFmldl8eQrZX2f67wVKmm89TfPIisQPhgHYj4E/wn9THPhSfYR
HCoIKezAVh/6j31n/pzrE26qpjS12Ahec20nmwaT8gKQ6Z0r8QV66hHQsSCF
9AYTwkzlIKPMJ5E25OAfNThhDI3TPhneGuzcXrTFfX6N874/gi31csqNVw/D
3Zs32PfKWOO5IuaHvCOWj/7GKWOnrdf5UZRq4IRVH0fpKGIJN9XDwo/wMb54
iGkMN8snCsv+kYahzoy9Wt3FE93VcVfLvvErgYAkDtLGjP295xqXn1Kw10rn
Y02i4/43YuFHf1wrlp5Koe1t6V7VpJyonmOa+iFQoTZiqfXSMWQ2KbSqKP7v
CpT7kgJnutMqyl7cfCKBoltPRdEbpf01+dmRIyXcaWnYHXAQQbafKt3kna5X
Y1dodrbfuzEck+f9YcEZfWnehtNG4M7g0pM7YAIa21NjgjiD3+TsOwNZuD8Y
WrEBGWN91KRhBD1rjh3lrieriaeneVX4OD+BBg7VGuhWFC9n7V7DGLiJwi/u
vX2xGKp/w4dLeA50ocmZSLcWKsybH/NjjEn/h5hoZx5V/ZWyxa07ZAWeRA1c
A4dBcYk9O7ALT3SysLwLUuQLqh2atFxMWTxndcZzguWv0x/KKFE4biMFDBvM
2QLMs9U5bwL+lITNgQHwlUgAWNG0PpWU/V/zCbRI2hqpJQ8WHKsy4ewKHRFc
AaBOiBsh9+tb9yLpY0gI1RaU17QdhkgVG/46fnUz2BDvM02D8jKy/tB7yuG6
4gX1AUcBRWtuIDp87eke9RutB6GZSPkeDrE0RDW4fpHedA1M4qoLx7b3AWz1
E2DHUb3FzCm4ajwE4QUHhW+HgR2dsaI7znGglBU6qubsnJ4bFr5IajbPFOoE
XQHNiRf1GHfWPCir45mFMw0kMxLRb3hOqBKlVhJwWe+jwZQXwRmptrh/oQ+c
3qtsQe369G11x20ofs+HQkk5IkIBrOGG/wclpO86UT9EWqLiLKN2B6ztxS97
+YoHFf7HEEE3Pj2MIAKazkYpDgoSLBWQDF5Fl778s0k2w95nStRAkY/hBlGX
T2xynLhbNj3CT0ndC6IMUOHW1ZP+Gx9gbYjqlDU28Np3DjZ5usd6qNxOS0Ck
BsG6UtKba4ogLdCDfZiADn6PBBR8exCR9N1dX+mBaq1bPjehIe2lRmFGuE+N
JAw5Zv8MUzAXHuL7CzpTiZPmoApTde94atvTh9vzHjBfnQ44NIxoU+t0RruS
2El+zkinBu4XL3AMOcj9YtwOiZkqshn4kSQuL8HBpWVc7ftNTIQY4yH3gDcK
nu3Wevj3XyMK+W2IjBI/MSJMgvqIBNUFssrtpzQUW67caeOz1Ttk/GVqsi18
6dJmoTWxuhKcjm9Ub1/AsdvIXRHrxFbIZ1QNre4j2Hts5Xb0gTfV6YzBSSz0
2WbjtyZqv5B0vfSHePQUR7QieTmAo2Zjl/3x1mDD5dsP0xLG1CKoOMGaAoJb
SIMeRwsblDd9qJEITm6XWzRotPWP7/71kycDClXYp9T4CrvxlsFa22dgyFrr
V8YXp+1BaRqrcv2GVpRqA6MqZLMQkP61T1fIZx23sjNjR+AFmPXytgFURyVZ
kjPiRENu13imSGPqoAlchdcs1mgZUF5lYBOJXppwpBiN7pf8B2l5TLb5ddiZ
eYDbzmEjAh5z6VYY44Tq4Q3LmA2sAcrA37ZGMG8rAP21BSCrl9gW6ZZGOoHF
LhwEtI7YtP7QXcdCIeFtz/9CJVF9KH0VuCRipnaGghARHMPqNQbgx44yx94g
vOIDolxMJQkravUmQveLdgLV23O16hg8VO6h02rSQ9MLJt5+1+HAfaloNzjp
BFzy1/k4DEQZseIDAy0O5zDpkUsrYY8KofYOeubhSf077ok9Ozfqaa13xfh6
khV9pcWPcWYuohM4tx6bPNxYWX6H4kTViEX+xzvyGGzL8ozRAGf/ZEOqzzqM
lnZc0tb54MB75nODZffPutWxxLqoNfihQBPi0X4l7ohMDvBhZV39of/+fVgk
KYcafwKLI+BPjJislQbgIMxVzDM4yptNmnbrt+tT4YOxChGJnzIAYZXypzNl
0EFH87oL1ioWEt2cnBfoUQ/ot4I5K9X+u8KtqkPifoKlDMCqvfXgAfe2lJwX
s/Qv8xk7FPdRdlOylScMyUf8+3AajYVEudzhrrvZaD6f6rJdqDFxhWuNpJoD
gsE8pNu6CSdOt0Nb1rpz7lGuXzGkdWi3oP4izEAKr/2JUGhTcyu6EjDu4E2S
DOGVDPhBB2D2FSPQbMrNK0PRzWtelydjmvb/IwtDugoV5TZhd0T8Ejielhy1
/hcwJiEKNNsapeUONeg+ArJxwuFN0aaLbyT7gyVi/dKYaCQKj4LcaObNfrzY
Emo7QtSEKiivXWzt5gdmb83WSCNOjlLWQ17fAfBbNWr5TVQVxFE/NnR0wh6L
ZI7nVP22CSbjlKKwjqagQSSWCfzq3E2CXpZPWtUadhX2Ep5uLO+L1yZEvraE
WEQQAHaNhwA2jGYWEXmYBvaP5ZaUP8aayIZzryj2hTbaz4gsdnqoMg4Yk2Xr
AEdtvi2iuYl4Yn48YNf4d1/ztmk3yERUViJMO+4QOS1YTorjxU4mmuIK0wpm
lRTqZaHPV7nGjfLqfU/ExBTW3cLP6XZVtZCoYcdVE3PlKlM/4plMdv0S8nd8
Q61PfWkmXnDMoWHs5D7Wsm1PWngk4WIqpJfWEgBemrc0RA8AMiikjTGjUVkZ
9D+Cnx1e/S5UXiUtX2kMS5MjgPPKSOcNhfNlfCKbsILuWncohLNLcIyUnsJP
mi9qWcMdJSr1HpM4018yKSr/2/D43DB5AD1eOP4dfK3DS/wmdrPd51tkCg0B
2Ki8sIvfGDDweEle2tViPQDpVj1ubsIm3ADuoTmxaRBaAyxVQqBOAGbMwWx3
AlkbruEbneUn9KTpH31RNrc+IyA0DG/j0JUA0CUr8Ef2eQy7oql86qqFMkkz
6ej9eZCCNVy4j3iqIKVdfemxVuDf/C1EVRhZnIjRvceLmzDQQG0mwzPfrZdA
e6NE19SM7QKCk/6ekuoh1IRaf09HzkGgLvnbymhAy8+sezqwLd0yOrUMwkAX
hF/r/w1/jFErnAaUf1mXXFPMzK6hXKLa7dQIjCA3vHfm6hstNXIBtRwOLCET
Jnn3JJMqxTJMNoQQVFr/VAAodlXE/qToCWhnABFUFCTCwIgeSTrIfVjnSQ/o
Yw6h7iFt0QmaBDDZC+ob1TO8Xgj/n3TmnA79nbEEZtTKsxqZd3kFu1vHiA/I
hyUqzmYajym3pPClcowA2Bmi5Wm8EdnSTmHcYKYqA2MDESZyYVLqlsL5VXrK
K3gFtUiN/q05ZUcTmmqmNkQP8YbfNTFDX4f+AZqTKaDHIuLPYlCvMF+Y68fU
Qr/ez6phBSPED22qPNOUOR7dZ6awaucGVdLqhG7t513hZXOgiJq0bIv75alt
Cf1ONxP+MOcnWozExE3mHwkKzd2QdFFk7RlGD01PCZgrj4DdLdMRstz4G4Ke
ofk6Ck9f9NS5E+1MOXrfcdhhyYXKzmgxT0l2zyGuFGbdkoBUF3mQ6MNUZ7vJ
pCTdEHDNfyr+DJ6EEeqY7aNyiCDadeoIF2WIUFjHrpuQgmBekcgIUR7K+RBF
TWOORm2OVz3Gw5sfKp1Incvtu1OQx8v4ZW0KT9yas4LvApD2DympP32oIZsT
9sagYcd9hE0ufodxXGUA0OQJrwVfWDn8WByp2ODbrsSpSaYZo7hM+KJl+QG8
8suEDUxP/y4vo7j9kkA0BKCJanYRP9RYcI/tjfYNZckrX89kuCbOL4UJmbUC
nj0dWL8Mb2fAZEe3Upz1ANe4JHeZpoMVPP4ptlTEd5wx/PmS9dHPh6ZDQxfc
1cFa73KTRAUWRaTAB9rHWN1TXJ1d3vin2qLJ458C5Y9fFSNNPvFf8A2s5cDY
kkLlHCnibIIJb1+r63vO6zZ0lyAGQI2KaB7/ULvcHWLBIFOpOK+mL99XcvSM
PWX2l7M5blmbNPaKuEqvnz2rcSsMDvef08oFxvmuKQ8ohOudMmW4FaAC/AMq
4cod1PnPmjFpRza2XFEywT3pkAEjh41eijA85zd8CvuUw29Yk5FzatQnNvnQ
rHKZROM0wNtQsuYPn5/uI+vDaiAfiYFPyzCXfCWMu2hXqYqrVJjAJ4P0FuoZ
bhluMyF1awmZtcZIk90zzhs+9B3QI88HbeN0p6zh17gGZhSOG6l8QB3j3loV
rKZ+yGK4wg5nXDgRRG65R62dj02LhovbKqGaocToJeI4h+rMKMR5sKXOKWFN
ky5HzxjxJ9QHF/gvbXx+00xWcyevk4RhdJC6ZTHdammowkAou9jk9q6nN1tG
OFh68bOvs5ObCDiu89LxIbrn42zX/vXFaJMIwg58ADCHZDFtbOiqAijoO2IV
Tw91FR3EKT7lS9aMTeGxqydla6rYcjaYNorMSgaIW6VLZgWGfJlFri7KAL/d
c57uLJ59YAqfR+xywdTbKS7vKVer+uJ71OUGiSb0eSG/q7LBejsZ/O0wzB/F
B9VRP69V2LWucYf7l5P7QUs+46Fsc0mik5WMQiiXhBVxLlJRVYvLcuQ/oIw7
26SIXzsRpGI5sT0Fr2THfYllnxLN6rYMLROiQ91BLOsziedQYK7Qj3OzvZJH
i5nBOjEL6PsxvaT0QAxDFCO6eB6XgktQH4S7yCQnO90QPI/+uwdfM9EtXcv5
b9Ys0Aq3HJsP9StnUHpkKx6MMZim6PLs3ELJuJOJG9uSeHSIlolWSGwezDjJ
0ZPBS/D9x0/W/ntD2fLgF+0X4ZZUpW/5DGNsP3VgbNf/597P5cGfIDgMhK/p
XJKk6zus1T/3AxTGmPI1oAgM1v7q/tvsOegpciVefELWQtMUGF2M5XUSRlri
/yX2i6sFRm+vD4/JvQgDk5qh0Lb0qJeDgdy7Etb0C3E14xsSy1yMbjYdKEaV
oNX5q/idPq5fm2Ojn5ywHohO0un/hI1uqsQNLdXpxLdRjLTnjgTvqwYxThTo
lr4tjZZqiryCD0sjzNvJKoCuxKdf4STjsg3DOVeqnlyAwR5+4+6q6HyBpFLe
rqg+DRKKtY/5H4vq8xWIsLICBoQiggrjofibaygfwAE1JQMwR4CP+WYIZoJZ
3eoMsnKaxrPDo0BOl+94PXipTPgA0QT6qiBYgFUZ/24jHeVx0QK/DYwU/O0o
0FzEl8gRwZrw1W6Cr5RqwzEatdGqx45kQwR0phLdJXMpNqd35EHPL6oD6bYi
JOEuk3B/12PC41uJfTJuPpzvfa2FP70MNXWiQPhJDLFf0Jmc0vRyijXR2GG5
4y868yR711HQxx2mtAkU0p4QAB1GGsXkolI0bTiTQEn5lrK5s5jv3hwz1/oI
7Fme1qUvbLlVc6az0bnyPJbO9mTjMGK6DiEEhi2gOPzpW5QtCUnGRk6Enkge
wfvUsonZCyE0t57cx3Y7ZAKiZYILRfsQRlBXC+sGEIPsluAcKXkk+BT8yNvy
0iUGWzcfKYGQFJQID2X/3BC0f+xQTVtsGOWMfNVZLebzCs6JPtYlyvAZc+PJ
68wnjm3/5j9GWjG2m0yh4FuSzIqqUnQbMQUGh5FuqTnIbLzU5SfTT+2K12PZ
8QUnFpvanKGan3BySOaS+tWdBNlY4BRM11wm/4aHOt4dmAgTccVlZBPx03Zm
G+eyFl+dsAebQGlssY7e8vXcMiPGRrFUKf/Y/GZGdoA0puTIpVHwpoIS5Exi
Vkr+SKVuKojULfc7qoAUcWlPA2otAKm6g+vJDx5pDje/hbG5ZnjbeOpJl2Ge
RADcP/ughdGFJ8AJyXRNMtBPrF2UmAoaLJTZBnXsHGEM6Ljp53hJa7FthJ8g
ijoU4q13twKmPrsj/7A1sjPPX7iD4dv/fSx9cvbDDE47sLs2p78EdjHO1kLK
VJ4wZfspLr8Kraai3LEXR5XaFSCeAB90bk8+BGN4nj3Zbo//yljCtbeoKsih
JngyVxgGrRDRAB2yETsRnn/50g+7xv2MAGc3nIv2cq0CVTN9I09SGLxr9hvv
Zf72TEQKTxcf/pTF+ieigh5FhQIXPFLIGBl560X3ZaUS1VeGCEpvuYRCNIFk
cRuaOut9tAbUH9wwddDk18BEKQAbIV1827TbA+uCBKjIgb32QnSbQ3kA1S+y
XYk3rCexeab1H+1KGKxDnzZq2a6VBeGXFOSJ+7zMLDHxOca5+8izK2ebG0f3
p2wArtR4Vcn5Vu6IbKM0U8MgvbuzS7eGhLmIY8tdbWfATgfCI7SNH0OpTs2T
N3+0uOegVddGIZrpgtoVSS4iC+xLDzJWSRorzZzNK9NiOXfe7ESCEEHqwSKR
rKwOInB+RUGAbqlbsYt+al+P6FwQh7uoyHflgKx/R78kH0wJ9KvbBgut9IfT
1jIqRuAOKd07R9bSIL1PYPtMqRsgmQ9aMd0OxxJOZ6YCVHffhQ81QsaZBKw8
3OCgs+2WFWsKweg9T7DRWzd5kHdhWmL0/NZg0nadoIf2IzULf7BOWUCgNhXj
g0Bhgbqtl6lENfsjKsI2lEWLlTbUAlOK8Tf0OP4EwrWenbJcqcJ559xBH0JI
PpjhxuYpZwT2L0DyfWlbngGLCunOfa0SULHql3cFx0KwFfDU+sRDNm7BDbXk
zi5ej/lRtI3Mz5d36aSChmBHXzr79orY+mJ/wx7iysY2X9K71TJseXxBYwwA
A5iz6ah8W2Uxi+sNHCiHDotRgtAOPdKAZv9gjNQq2ziWHp+6zpcEkStgfDw9
DgaydE4LmDtal956q54XwFlzQY3u6Z3hnZckXmwYBh+IGbefRcwzjAfkIga+
V38j4ToB+Y3qgV7NC/NdbVddvFqLoWDmHw046o3h0YEY9K89apSkU8AAVUDt
sea/dCrDWJfwmxhhseKIVwXe07ZSdqhM13c/7rXsAIplkj/uUdfB+KaDZM3g
IJxtPQjm7FeKZjKRHWzTM3Ay7Y9mXsqz4ai2t95JrXHZB+Lr+mMY2gKTMYnl
DGlia/58gx2oNydL8Kc9S/PbGA87RR9iPm1Nf0uYMKcKdGgJiH1ieb7/AKz9
2Mq+l+yS05KP8CVSi2qbVQhOhQkUejfhRq9UrVi/CxWhYJcBqkwl8LsFVeYP
478B5E+GALpilNXTJC1CL4K0U5sW5d+xf5RpnCMv/MFusznvejhVuHwtJkAw
1Rws3Z3wSHYsyD3SZGnZYHrAICY+HiJaLAB2IM/NlQNZmgzM8aTOxyGew53D
cDxQ8moh5ovnDgmc1ha1Cq1DW1PaGazr/4rfUgycFJnB9ZOtl+JKoD0ENhCc
cOVEu7+kHXZXtjZr6LW/BfRlYH452Tc6G8n9Bpo2ieLoDXt9a6Tok/QXfwuj
EqFfmcgBRvbenr/9GBLiQ8DTh7O7Lh4JZ9ElfJzKmN5vyO9m2/sBfbNuXWYp
qLRoWeKRUhYGLIWhVfx4RH5tRmWdRARm49eaYe93rhPpAhjJsZ8zaVE7I+iK
8D5cINIdjdqMGpWQY+Ww5NjtiSAf0NF/UI5iWZfPzRA2uGX4alexOgjNBCKF
W9R0+3NBslUxGVj+SZL5gxqWe8JI6peRCLOaBSHA/r5Svg92VvX1dYrmO9dy
C1khfXBLcxgsV3DvjlqiuPisXphjkrzhks+dTOhfibh8OAc0yHIRJpav/T1s
t2/STDAdSk0EXUrnYGqecKPIJz2/UNjvgVomEs4LN8FUlokfEHdjQonNBCv5
r4HRlpbmcv27rnx54mQQDXqOQKBngMQXNoTQ7AQC4chwNN4AmYBLTmnEBl4Q
pV1kSKd3IdqXdqQV08UZ4y0mO4aij9pcp7ItVhHEVCFuvIzYu0mfdibBrtfa
v4AHtSremFGAaLoMEHC9Ez6bzujIYKgaWZ/pjBcACe7ahks4E4V9xRxbW1Gy
LI+P4PxvSQZQhkrCHmt4npC4kIw7H/8mcCO8RCWiMd1jtPRit8BbTJw4On26
432id6aFshJC1g/BHX6zNcCWhi2QFALUrVJWeox7gnA8Om3ue+ZbFW5I0Ejo
PydADfma2BlOxnChJy6z8N97FFUmPWUjwa5W+BVfl+9/MxJZomWKG/sBRmhM
N0/poZcAE1yyoPjq67Lbd9k4mKGHVCdGqg5gPZgOS6K0ZjSkeEzf7TbniJhe
9RpSCJHZQZDa/6+RCat1zjLC7W9O+oPOTYaOkF+MFwm2CCUt2DkQi1dMjgvC
7vkTryBvaq6kTex5jnXhYEGIe7I2jzkoo/RWN1jI4oYtvotNHMvAmZdgO8KJ
RauFAsNledA54yuwem36HscinDu7ObAHnKnkxWsfB6t6nTOenZj5ELTeZL/T
8DbxZr1vwW4HLdC+nxMYhE3RanmlyIvXocxCDiM/dYqwVj/aSOIz8kk8Tb8U
UMnzuKsSdO5wrIJMI863hRyUel9Ko1MwqFBuxrGNVjcUYo7WUqNZcmA/GuP9
jTbyivVkuN7RlwRTfEv0x6zmIBKmFj4ZKztLhBPyfNjIKjTqy+zlv3DrjeL7
u+KJBVZD1I5gS+bVt4peq/8WdPGPLAb3k5L5d4opjZgK4QldGRDIbX7g5hM6
23lQXAda8ZTlp2UjLL2wyPG3CYYvw2HkTRqljTm5Y43LnKJ1gHvif/svAfHT
04+S8yACgiCG/D5qOzC/ZZbhirH0h1cqalPyXo0Nl1Oih1iitM/P6PIHrSyD
rINCrXciK8hCviPB/NxE8kFtl6SpKvui2SwNFVqhhvV8iPia/NUEyLo+wQ1e
TyW40RJiwbWThX6p/c+y4Ohz+aqz3vLNiZZ9oWrsuOVn9AegyEGhC63mR+wQ
FXl/ZEik55VC8WmIGD/l87zf6emVlWO6jAH0YvCiMayfckbaPX4W++Rof3k1
UVYdZWLh6hla8Hy0+kLO+54DeiHW5xlW5LjHrMgEQttUrmuw9UR5sIKIqfEe
WRhnqryUlQ0tMyZh17sIB8tMrR/sj+MnD63+GjO/cN//SHBvQ8CRv+cFGfuq
oVQzhE96GNLIHf52PuwrAChY1/MARcXpEYHMkuif9/zK4dEM46zDMgrnvjxZ
MEEStazar/qMIo7idiSsWXfWjHCvPGBq687HwJR0bIdGoa1ZOJmloQjtx1E8
u0TJOswKvTNDNVSm8YG3EB9ptCsfTvC5HuVDs1Jhv865fyvvszdjI9BGw9hI
XjuHxZDPDkQtSMvRnMQ/Ugdv+0Ba6PjbhF36rJkK1gVFXr2S5giyBqvhi8oc
/i21KgT+MRFu73/ym0o2RXW/ITlZpyGXrk5zx2rIwtZbmGT3ZgFadO44wrZp
6CJwj5l+eHiG6H4gTcOn0NY8xn+a7GZGfTji0E/1PdjSNmpthV93KA2Bil6r
SFMXSs1nyP2pdPcBN3oD56lW5Z3zHN/83pbeEqQj3jl9kSDJVIvc8GpCKPCO
gRaohrDf+xW7aTdbZIvpdrj+Oa4nkh2+rHqQ6vnpb5+PQhBtaiB5PDBrDDlX
VxHTrbtCsxfaWDVbG/Utgv61ansHVqYwmLpoidKwJ/QP+h5okpG77YY42Ahm
q/QkgiaMuEN3CB5sb483E9NMWSEvM/baZ/FmWXof9itXF4iFfvWilEZTLyi4
C8p5zQtoUrXNG1rbtg0TqYABGLP9R4jH2MJPpAHSOueBf+FQOXhXznY8tSAG
yVPiwDN2CpyFl5wrsSmKXnhBaL3uiSLLO/yd3DCQh2gJnr3tbbl3JF8JJSJc
e96Y3cKGgc29QtAKGLUYhsBEg1R3sgD83uU8MUzfHdOttigbaZSgkPJCYm5h
lRDjDgqTcq9HmnWPn2pYbbFg+KoAHHUWxP1U2hxwI8MpbEw4Gk91KtBcSb9o
Z6ZPgZw+wSYTJArzD2pYsulkNSDBOsW49zBgF2md45XZROFl0C73Dhtm3UjT
2GjSRsboiekXt6CjNemHZ3AtaPTaQ9cuc0aU99RcUhpgLEi16KQ3+n3NLAPz
GW9Vrh/wq302M6+Q+c1xnlnBvybgemBiu931W5QFeLlUs/pSPx1UDuo+MLnq
SR3mP0PWzkfrJNbbOHECZEkJ/kTTLLrarZbR3vQZzbBm/zvhFoiV1sLVZFqq
K8ROUOTfxQAi1fW9/4D8cDM71FO01SQ+wKt0h2rSNv70E4wawiPdDH6NJGp0
BzEvmvXB9yngshdO3T0LuPwucfIDoW9AnXVyD83huYvR3YC5QBwe4jxCbojp
MDWYcifUtrhDTIEafz93JZkU0Aaetsn4KZMXZGRx0pw3IPsesQnOaJwPgh9+
MFlV3VRXP+F/UmrDsYM6sYI7gzfdl21XuRlXIyg4bM1Cwp8FHGv159FOvQiW
Bg58Pp/teoX11zL5bgoBvFvhxLwAgyXzx5hORHVWyZnIuD5iEoTf24hhc8oG
5gQgyEVW2bGMdTroytv3s5/UvOYmFv98YHzOleojDw4WGTsiOUo1bZAaPwcO
Cb4w0ru9IQYUxXt/sSDpR6Cjf0Gz5NBxe6bM2dDgkDOUjmL+6nBMIc3rDOPI
+6kaopr1hZBZU7qRe9/O2VUQqeLpzY4CjRYw/QbThMWl75qcFbwHw1iOoWoV
uskf8ilx7FOAESUaqZPFpzUgP/PkJXeQMbkTS7uWjkx+XJQ5hVhbSgBz62Hp
pax5KpHmZ6okhNKO0MZKsk2j4PwVktRaqyF3059kIP8FVZnYqVTR8ZZMXyxo
xxuMTMCkGdohqGOpwgLyMmslLwQFOyslHi2vpv9m5Rb713GdN/8BpCTVXnqJ
eqfZg7e3HxjqDxb8TKI0oN4uBPdVLWOYoYWFLfnFRilr9RlWe0BKdQgsKBYe
up74ZArAINUZZB2ULJ4ZHBcT/jGNqTJx3S40hOWG68usd2/E7naEe0DI9cJm
g6c6Bl1BLxy4eqEqwLsPamOY+Whmke8ekvrLToj3l9JxhC+ho2gvc6YvpQhj
UjAGeMVhtdotYq+EBBpnYoU5fsTTw3jcY+57nEQUQwmp22D00AgPC6B3gOCK
WNQHBG6MbFelv7UEsD61fVUNClkUTQBR3kXj5PngYZp8JBUDo9ZdJiwYPDCt
aSayM5rOSv/Ajl1Reb2dUeeRAw4BNDIyT0tm0UmmrAvPCj8w0wPCZT2Gi0HZ
xoF8ypSKxmrm+5JfYNY+tRCmpGKvhArCvA31onox0hRgXZJguVFoYWWByPHE
+XWnzfIlr38fmsqGwexzVi5QOIUL7mVwMBwJyBVVSCFQXkvmi7we7b1rIIYf
dsXNbcLUPjB98xsD1SkSDZ6gRcoChTNS57rK+8o5EEvpO+pY9loZ04M8Z3Zz
jR98ifAylLY5cXnkMyUtC991eaOeO2YaKmbPtIOACNk+9GKlL+YZ9U62OdeN
B+K4t1P7yUNRzIilsMVsOGOnZfnJCQ2A/kk5MKA2/0N0l1MPOfRPNJn4gM+m
FwxcReaD/QZBcDmsXrXps+cldeKcbUYXlqynXJTYBPtJ3OYVggiHiNIp8hTg
QXR9jh1JRqYwNMF8QKlzbQ0t2kSPmAIyx18Q5q3M2RloF3RpGwAzCDFjubKH
wJySYQo1TitKhlDxHi2afCcxQG/DQdrV5e3hmRl2cOJEFpCvJ2CDW75od4F0
3obS+Kg0GJbqaZ6zU380F/NPesrX8CH0IN6qBVGmXF+rtxj7V4pLZaUOAWZE
E3I8FOXF3DUnk6paJEogU/GdTxMApY4ojG9ZYBJ4e+H05NOtLKrsbvV9Bh/g
6ofVHSZllGsOqHR9mWWgShrI30KLso1Of32WLlcKM8XdAFInqVpAl0QeC27k
/uyzU0c79wJXXDw8QkWdmZYyV6Ty+9L/2btSXgEXSYiiej+lXGVPalzkHE2O
QeofM/vuM1t9VKLsjWr+jLAq+RAYQjAoWtFnWTF8Du/shBfPRayxE6AuzC1v
DAaEvjJZhaC2cgE9YamMvWqhbeOKe67vfIQL8I/ocxbS8DffQB/0SmjU3sXA
An32ofFJ0wdrsUMfhq/dq8ovP4kbJSlQq4GYe2//6OwzKtYLIH0NbgRe7iY9
Ba+U9Ogdr7mncJM8eB9Ol3hy/xbBEygGODKm/do27EU35/YyGZEgelH7gMUo
EukgbUF9aDgO3aIC4i+9REq0JVPQIWFQ5fMQZ8vs7XTBSWCc/rq4tPq07HlR
O7P60v6A1vrMXH6ZEQRqXNlez31ljr/G4d/UR8S5A7H1tKS9HfVpK+q3QbJd
M09j+Wq87eE42S+mQyZguBNVl+XmlwcCFj9j6nhDhm5hz/SxLOFTmAwB0IS7
ofFUOOAcMUtjutPm/Qj+ZemZWuxLFd9sa3eYN8zpF0Fvg4LOsMOMJI70YJMR
bnwIP6mKACz41hU0TMBsoygq/WurJ4B0E+Sf1ZlX38LDRRnGAjdo8rfBPcBY
PJI62XYDMcNYU7ExwGt5lOPW1mSz9H3zJE1lO+V+yVGiZThlwZ78LuChIcpN
sozQ1HGz/zYWgHZJKYo6D2V3K4WZYHcUKUILfGqX89iAejIy3jZFQl7QzpOs
d7Qis1b7bivpeEAiy6Zu+xRFLys1p35R8w5m8bws2Jfa4NDjkJyTrz7Xahse
ovs6ILNj212bVBwdWTgdy1ekiGEI0BozpPNiDrwAIl5aF8Ar6bhxlQ3klK7Y
4Eyf8DmCsz5svPF09pSyggExieow6p++l0TQlMTIHpB/v2/gmzcgBw4sjoNP
bEVH25t6pqTpqScy5OH6PGPNpHUeqAOWgYKVr3KChuh7KYdaz6AJXhbvVhuw
5BUBDY1EHTXj4uddBLcx/7/+myNrptiYs7E3mlmBk+gb+TGmcNnrkfrPH6B6
M1h/5cP9e+AJB0U/inrmNOoZRH4rnQ5tgAFyKBco/GBU/Aip/tXbYSjh3kIl
O5GaHn3k3/KKZY/BVE2XNlZObdvC3NZEc7xD1bh8kh4Ca4WL6wgwYTNKt85z
OuIg+S9xHL5IAoS2IeMAP044jmFfybjOHc1XFcWgphWuV0wDawMNwQ3kFIHS
tFiPXileCrCZZZgGwfcMAEumsu90yY1e0EHWs4jWitomUhP1t5iq7Mwb3P/Z
U7tah60ifcoK7sKtv1EJhIK3dBlO45f9Hfw2RMHBGFBVQiX9nrYeso0kZYsQ
otkdRWuSy6l4jcfZ7TIyb+xe+hsCL0wAGD+TEpWc0ln/rYuwwGrGCOFb06Rd
ID4uG7zoIvmdqTXK4MV59srFlApIzCiuK31ZB+3X05WZOKfzEjYNPcQ9cvXC
0QEVAAoXNLtV/I6OgJ6yaqN+WRbqeyRwB2BVD+63bvtaJyVgvrMI/3HOPCET
jmPlHR8kw1NJLGgpLw9BUTiPsLQNXBJ0h88l00uOIe7soh9pKu+bj1NCu8y3
CoC8Rub9pC3umdE+rfSYyNEVJBvyOzTWOEutu6UkGh/Tm/pQBL8Di4U3siCY
qmh+uePKUPplbB+KPWPF1NoOzmURFK1YFu4z5yz5owmuHnPSqh/nkn1D9GzT
aNNMReo9CYzjdaux9TPi+9nbqAeml6YEsBcRJ1gxnBE6cLRCbC3orhmyqDG+
MCinyw8QgK8pNzB5z4qeiQKQVJ9pLWA4cOFgdK/IL6iin/ElQ5i6q412zrG/
KL2X1cBcYLjNGuX2fPkAOkHY/UhJjKsJdnLy6LYNfW4x83ZgRUIfpTVI/79d
WHW7NYUg2KeNL2z5Mtyn/g374JY+dfVHNvUxCPjM5IKTas5B4vg9o01F+1m6
e5J+t3uCZrqZVI0LqjGmEfDV70zsCg3J1lsTzTUrcJcxslQIXU03mb2ww5VQ
WNVut6qBvvDMCPWR6K2eTlfvky/Z9pppzoaWmGZha74I+M7kh/7MQ0yMg4tZ
e7GsI0vp+1rz6FrMROia+QwS4leCeetMEcpe3FH9fNpRNdXWTaWTZluLO+9Y
NMgdUp6oFjJmHlpitdYB0s+steFHRpqmTKobCCnBfj3SyXEyOcLsaOXeagmZ
g3A/X8WKd55AiPut6uvC7RjYkDKIMtvsoPXJmkKUa7ooo2Cuw2mnFOBzN+pI
xwRr8FvzyGEK+3PQvzKItNq/c0XwLxMXwpBBi/v4CtntmH9sh/BaqLxgPCyK
kN+AmTGKc4T+IQaP4KUCwqEsaCyEARzxtdphCj/dpxufFFRPzpDHkv/CZewz
EejFB4mrUf76B4y3Gqk5ub4BtnD0QiOecvAAHf5AobGijdQ6444DjrCYsrbu
YVuVA8VkSSWERmJb+LEa45jk/PmLzKkCkPEm357pQocQcaBGvtVdrCQyeOR6
24qW5porosCLQpztrR8PPqGcnfRxQHO7MO08yzh9grXvl9dxgvD2K9GKhX3V
UxlWqoLp/4wfJ1oxnOUnKdd7xSUnGONLRceUcv9LnigAZb1MrYO76uKdJDKY
Yn2oEpppR810KkwPJd3KeWWx6EXVvSmB1gXV8fKQ1bjRD+qt1KYNKHGHeCiN
IlVyehog3qBkdEaZe3u4EPec3UOMJ8lRPcCq3M5Pnzo5xqe1kkFlWM9iPLw0
CHxSMipBBh3e4IB9T2dlfnb9Rkwaov+bwDOg/d0qmVN4aNt0WW8yvzrXIY0u
AOfjZU/xikCC0Zkf4A8l+E5DLm9G0+IKVjvCWuTkh3Hdn1lNh2TFwwtaFbIi
JZUN05GxBUQ3Gdj/i0z2V9EitS8DTXjzpw/6HAb47ELVAYx+4gtkHm1XC06I
8Hz4wH80cExf7G6sm2kUfVKRNlPK2NNJTtBitDgNmbZdnrsY/w5NMLSBvS96
Bs2EMhYOhPBZ4NyUCKqzFlAX41ok0FP+StZ2NxbJKyiL0SFn3ZZnA816nizo
hAHM7ms1QVA15sX1GuTcsXInhsf97cTf0AFAeEX0QjIwbX+eDhj8aFXMrzxW
/lHeXxsvXZWlKU6avTbDVty6iYOUVGIaQ91rJ+sKEA+RYg8lAH/A7FNHyoKi
Tn9iYfIPUnds6HU0BuM2KDIDKMiJBCCVbgzae7ueNbvokCxYSRk+Qj5uxBIG
ruNgZwp4+fTkCMH830NliutUTXwk6LGfrd9rvxfGEb5HHynBbtBkv9qoTpba
08BqM/WdykpbERjhj28tapgJgMqqqXVzm7YQ+OEoEQ4izBSd1vDZNH6GGqVx
zVeWje77Nc0ZEbDxNJ8FoYdWw/kLWDh6smeQQf1kdYAs4YCBjJqIOl+zg5Y+
QrxBWaabMAWNb1xmI8a8g0e9W+B1qFZ1EyLaZu0IqJLg7mJIoa2Coh2b+K0b
MjNeRqJu6o9X7VA/MnkwG4qcDV4w07Z8llFi41HRq/kY+wET3vp5xjaEmqEl
S4Vj22ljClDozX3xo1pCe+VySffEMZ/+ufsTmMRGsDQs2Iy4Wa3aEF3M6JXY
y6BAr7+gkWNemYOKggiHbEJRsTT8Pht8RU0W1MV+MxVQYWCjADkq4F3L8AEh
XrBYkCzFepp7dFXu8UwOkrJwEtSnvWnhdLZNMcyXVNcXpIb1rUd7Xz9sfj7/
GCBqjHXrAQQAAn4UZCpAN4hfw2D6jYV8+G0les9lW8f1RbuYZdc5/pH3c/w2
bODpWRNG4ibHyNBI08cujiGnsfUp6N310HclAlJfcpW6GENlBUvQaMNr/blN
OJ0lV1uYhzYig5+lcPazDzXi979CdDM02+cHi9dSXjTqrNnXMO8y2DRqEc8u
6EusSGyRIBCP4Pmu6kbqir/HXWos6pQAPpm/llc64BAOPi04uLOjlbMq5/Ap
nSJWTzl/Z0cuXCO5vJEg3RRyjvmzYoxa7B+iQYVfrrHLert4RRsl7jfYg6oz
EIg8yVpEQwzeKB6QFtAnPczvtslaHcJcARCxowqvLcR/AccrzkcWRSnIEcmk
DLuTsB5mOEXNN9Tfe4gquONtZAqqvJSOj8HKhXnvPhzo3qsXL0GyJh4FWOXg
uFrMm+LndodgAOrXvF4Y5EP5pwzs0YTYNwVhTdII6yeBX20cp2IoVdAHvG+M
O7o3Hac8dHFWnfrnuHHIA2TfUmMcLEbem8KInFrYj9q58dcTtbEeB8Ofksk7
3ugLiQz2QhS5muZ2FkJRUCkKVanptWhK0W46Vgn703dp+7SPVeY1WxKSN7X1
zTtnoqhtckPaFG9b1WGhgiUjvCtRq/vE92U8tK6sVovYfmXWGN9IXNwXmIF8
TSnfh/A6xdTZ71DOrQiw/ojwnQc1175t/FtupT6idryEYdt3jC67jGr5yvMk
GOuVYl2cmPMeLepEwP73/7i4GF7mYiYkNbth+WJmpYYkU4ZRZanjMMZV2SF/
uEWv3OOLLa5328uadMVQ5r1jgzCWVNaeKqBzNXGZxRn5ySvRt97qVAh3WhEr
c6g477iaOemkMr0o2c2Ckq4AnVHcF18bLyrkkAFmpFQbjxrSsceuarJBGGiv
ftfZ0FUdls1MsnIayhyeV2cqgUQPezPV61QE55CZd3y7StMRzVjUCgbSSsGR
dPumDwgE6FFrr0lz3XqwSro3wWd9OoQpqBLWoyBPuOwuSXxQ3OP/xj7MjKcG
YsC7CyJalj9u5mkMQ87q7FVD3OmDf6db1fn/UMPPRPjZdsrNCmEbn6HIvwTb
lmFjp0AGmDtJ3+te1IY9WHaEJ7Ja5nbLHhY+raMFfyb8qMzmQpitFqLzsfVp
o1DFrCmmv9KcXDpIowePkOiBXoMJ9UC4P17DtuwtIOwQ6zgz7yhFWbpxCW23
m3xAAlOZwaOor2ufD35bKdhONsp/7K9i47eW1pWK+aWitnWQVMXwRXZI2jCI
3h6Ierdr5To02PyHAn8jQVqpanfhVdiOlBah2LexXxYMXGEqVa+aI4FfhtpE
Pn73c0t8g1IH61v3dBizkRrr+iuycnqNfanp3YPzxLEEDp8/5sn1UYoKHTN4
ldyUF7mIZboc+1oDdk8Um8flVAsMAurseO5KzaMy0AsOANYmovyXDyFwHJ1h
k+WfsgN7J8scGKw2MNG6KX+uNJ3CHqnQcgLBeySeITIHjqXIdEsixDD0JnqO
AwUNuBxI66cHeLBCYiqjWG6/EG146ODHiP1AVtK+sBEhuA/R2SeUlBNcRzH6
/oVNgIjLdG2MpjynaZskx7CFmyfDdtqL7DuKZG7c09xMX/3KDB+oV/djLg2o
NZE7f8AHaqLloYPpwHJfFEYb+AZ2oqk/FLzXimpfSHlgie240dCyLQJypxe3
CFl7t2gwMokkmgNcuySPY82fBf0OlG++dAzvopOnBgwNDjXepopHmpbYbXcT
0rk8Kko+FReDdzJEfi0t+n8VNAnSOR+P8vUn8Jlu5eU3CvYdbxgA2E2Ne4qO
yC2AuNXZeHnd3qdA/f1neyIdALYb76zLnsDfHyGNBpJ3XT06MwsKOydkxjjq
JJThHChdATQSYiSFEQkR2Mopr6XUNPq9LT2d4AkW28t0EY2/9+AbJyhA7okj
yi0Dfm6gThsDXFfZS2jjMt9f4YquBVr5p4QVu/e7WduJOLLhBwSGg81lXN21
4RXHNOynLaxMtVpzgnWyevFr7tIDGt81N7BTSuhAirum8q/9M5EkTZ5GCuVZ
ijlvXdIz0r3wFS1kA8/T4DjmFG4uxXTyQIZQtlKdReLWT8rBl2rGEFiCtKWX
dZttir/We/WSyIZiqTtX6188w2p6CZWV5oFPqauCdOAw5oOgHOOJdm8zfTI0
p1K8+EDqpJ5qwtrJ8DDMQC7HA0txZ4oM+iiQI/gY1aT+RfBCPdPNKl0IhQ4P
GZphdF0OJ+o61FoFr5nQ54FQdtBe1BiTF6g9CUC/8YzjC0Xty/bSfGRuE3Mg
Paq1HXlXDn4ytnmiPqqZ7zgIqPxlgqWoqxYi0EqCbb/qpXggNV0hf4CFlyZO
9LPbNQgFF7YKUWioS4Iv5N944xedav4DPyGB43cYQn5a6JbWjZI6JTV1e1sj
LQZoqTgSF3gDkeoFC9/znxLVd1lOT2xjh3FXQTwRaFUtzr67VZ6xfj9DdSK3
gfSIf1bj7ii0vwl6hQIah4RdM2y/b6o/lmH+7LPGl3b5AJ6Yh50rwCOsjoei
Mr+Vp6uKCIqgmAGT2kRL+4VplZQgwy2UhPWdlzRnrvbJCiYYnx2v55t5f+hB
R5Fmg5Or4FWNUirb/W4BhvCzMiKk6Z8VzArXPDJw0QEY/w42kniKDHOeJI8V
n0EYzuXxlMwzZdLd7Z4Ba19wqL0dPgBc265YUKD3ZfnBHFgNIUbbTnPlSvId
Y1EP9u0OWdefRhGgveaqzRTWXGlafRk2WaWY+834wg5kIaqPMmaR74+4gSnk
/9shjfi31dkagN7K2T5Da67bPpQKOxkjOLTRqfXH0ZjPys68z/2jaE5GVcJz
FFfKCjWhzPekBl8t/Olwc8D+h3PZfIQKqXZQkxHZx74PMySZMQ5dppWrlayt
ovLFdnL1DfYz83r1+7f6Ii6q/+X54oKAj7R99yJG7V3gevzQ09+tpw51vRZ1
NdVCvS5Z3BwaS3X0W6KdvsjYDIugRiQhkj/mR9ssx9f4aJAqEGPd8EUOZoUx
V/+BBx2GednLjwi2V1rWIOOU1ohUDnOhrM2ighWNI/okNtBEsQSKYvoyrn9g
A+Z+v6tjh19pX9UVcHe/c0VVtcQ042/QIzPjtDGnc92EbSoTvzXI34IYlM3P
jXmrq6p0ySPU1BRgvIRLwrunAgJmJd+0oqZ8ksuMhPJ+Qx/G2ZPTCcGuIETF
1ipEcuPoaRutVKgzvMD2sa8YVTGdNe3jevUra9SYkXkeGUYFxafbBa0Z41i5
6t++N5OMhaJOIr3CAVSJvemJTX5EvAlr6im8n8q5/Tr0IVtOAKtK9XJOF5sG
nGBoZaoak2C53ZyzRCHGyVobchVjqILkCu+9G1mIqe+OJ71bBHCsd/lrTXQd
Enk8k8/YGJYquipR307uZsO0zweaogGuqlL8EJjbKtlX8dIVgmSoTTkPf9O6
Pb3HksKhlGsHuDirE8k1cayfABUYILenyEt1Vs3YYr4wSTej3lOEuUMj1lVY
jQHtg2hFhUy4Ikim1F/6axlUDFGS2kMCOS4UGYoviRVQBDuu9nfgNydQNvfc
7cYyZGRtuNaNPpIQl0Vqjci2303siZQ9JpNeiO/ailLFXLJxnSvnhVIaDFKd
7jCocKGSx9xg+WdY9Tqw8W001/R9TY/kxNS4ZP4nuu/QKPAfHcuz9QhHW7Hi
xsH9JADrur/slpEGI51P1gL5GkWq8Ilm7PlWsYpwyDT2O6WFeLwZxOcBEqvV
TY4GoAlTnUpF5i1KKhLsIJnEZipDfqe4D92TZO5Hnewyg6VFEmrY0Bo1n9mD
zuD5wmAKphkZWCOEwwzRzQiCFlCT/j+QRIvVapWHBglHzEqStkwRSUEKa7kX
cTkhSLoR3pJr73a6Twi9pJV38IxazpglHbZDbL05bJt0I6xptXvRsgukvy/y
9H/+7EZy0PYRTl7yIOR0pLVulGjv9zISUR9ViAOGdBLqq4hpVh3JdOpfBhbP
gWX59gep4vMfH9mDaATNtoof4vMn1sohXeLnz4kkcf7IBeR0S21Klx4aGJrt
pGEtREPMnVeK/2OF7jRsH4u80tIiJEKJTHNFyyBK+Uwf45fMrSJR1nGrYuNB
TRV7kWrwvNDwybdjIFre2sTWfaRIaJYMylkmUo99igjQLO1oBNNBy9njCQUt
AqX7bYzfBbD1xopYxMcKiCmFKa1ph3VirOk1tMOkLD8BGccly+YeTA6lvKWw
7GMbOeEkhNUTsyGjlYIQ6xfqR2LWJSDKjHp3BOK8EHvvwtgrypH38m9K5Kaw
DVm4HEgvdypb9f3YKCQi6CtcCD/aAfCOz2nA/VG2aSAyk8xira3xZZoi9EPZ
fIUCAuDcyN6xJc+2vXNIzGN0BrWepKSUvrgdsHCU7nURR3rrCcvyrfLTlLxc
vVogbE1UNMxtpZM7bDksPt4hdyfBX/0398Z2gS6d7933y63AZTUfznZdwHye
MkVWpKMFfLJ+zlLirbEs3KWxEW3v/+Qjn0sZlgUgoZAyJFmoOdt5Tqq33QHI
N6ifLADdGWb0UIvabpfe796XTaNMkOES4hkO/9CdUCb2OIzqxiN5v0CxWz16
l6zyhUlaP/Woe5EO8ZwGwGpUVVJevM40SKV89sbSkOfxo4D/cdDmUMoV1KnM
y0bIr7cytzy9i8mbYC+xNoWT3S1X38yy/x3gJYBRZzsOBm4+5KyR+SZb/eRJ
VUEtQt45oNEDotovseaWOI/k/0xfqfmx71xXE7IfG8pC66h7bkArw+jawlvq
f4lwTTLAUHBhIxq5RIJ5XU9mXFYS6u9ZS6gva8AbzYHp2QPUvZ5ktDWDGhT0
Q2PuWCLZNsImx22Rp3j1160KemC1QF97BbqvVZy0nzsfCuDt7WHCAyXklOO7
HcsCgF4eCWipYlBwvfXSbOJfS+f87pFzd4Dl9drAHHmapGr4f+bl5WdyBBp1
WwAB+rOsODafdijCaSAMRyloiDmTvnu7tVHftaObBRCLdtjrQ7NdOgcnzUap
5jHw8nVwFLzqrJnY9LfUaXyN4TcVEZnyL10RuZQKjJYkE8AsRbFwhSeprC8q
3YdwDiRhJTqdl2XFTU9WFkeDFtge+25VjuyzUIzSq7ondWoZ6zv7gRUwV23J
ukM9we2TYkS7wB43YChuKA/jlqQRWIOtdACo2rxm7sayAVJLTd0kbGhZcvQa
A6vI0V3LesBxIvV8yyXb1NZCpkMksdUj4P7O72PAxR9w3ceS8rxYVcih/fgP
93+i2kxfd0TDx9rPUwO+4atEyvVLBw8PlmSoQwRsWCEM/9A4WBBAD8nKEJgd
AsW/ThU46LADnpJ5YMkrVzKJU84C6w0EaYM1FEyRGlRGxOU0ywXkn9C1EIVT
ERzt+D7q6bKwvU+j6MfTeyJKg5p4zz8DE1peePITSVeU6lrwnuukfV92SPEg
U4vAToWIacCsV219G7sruJNaUC6TOXkrjaUoS7MJKBNxMuWlpow8gCnZdaYk
T5kr3Dfe1cFnJpDqK7bWsySnw/6h177CI+1rAR9ChpdJzEwFuJvqL7FMve8N
IoaD0eIfW7ZI6byGd/Q1uHFFwCx4nC/mJ+85rQN1obBy3AzPf85xLKNBgDVE
osb0IX6+i9cdRYj7+mXwsdtziRtb3wry7nRCgQZt71iRAMX4a58xQDWeif52
UDzXdqJxxwadcUXVmuezH5AIwkVJbYXAbFndG+V5zYmb5q4tjcOe161JzTG3
8y8wqHVP97JPBid0CdRP36KnRDmnoyQiu+mbfykitLAlCOOWjREimchJmViq
O4Gib6BlCG7F6scR0MSIkXUXDAhSlgqyrAiKIph1BUi+YhOoP/5rMZMKSMRz
WZ9BGy8+VwQNkuQWIbHIyiL57zIXVVt3eu0t0M/CWwnS+e5/9063WsG3ByfE
fGbJc7Fgck/Rg5igSgL/53xZphDI5mPxLqWykFzxEqDVRXmwzNLdUk9c4GG7
LoJeaXr3+BygiExmmAPc9oixK8yzBjInP2V1IiWV1aK9Q+g5UVMM1Z2CRaNl
HSks5ApXUOF9VBV6kPyB8kICkSc12mlxCRIVuRs9AJ689slE7oCzaTdDiV+b
AJ3Xph/RqBTGaW4qmMIdcTnBVkSAIXNvHsOZbsAmO1S2QuyfC+vD6EfMFMNY
pddtz0beNmkQTwJXLCZ2BNRoaI6KkGiMl1DltIXkSZfRanDzWVi4HrFMgClG
N5luWsIi3EG62spWXvctt+k6z1yZso77Matrmfb26dXyyDWC64C5+0TwV7h7
/TuF9Oz/DD0MMgU8X1FC9nfVoJLsnj00dmAvtVpkZ7bpZAi9PifyIzTF3eiZ
BOh0iOV+Qr/2N82WuQuYLK7F6el8wvQD6oa0p4m9ZO5XuN/Ff++D4aAqkJ+E
RoEbGnkznvoHwgc2HEPo0Nqy+I/fiT0EW7fmd2Y4cKzrfX1Br6lxJvnq/QZM
YdVyT1vjrpFH+osNN93G01CYNWX1+nB0uLg6SZyeaFyVi/jI8XgP0pbgevHE
i/0QuxJmLjIMBeXMVvmDOxN/tag+GjuovRN5sE96XlZ5x2Lf/M7tPRprx7Vm
Irfi/ENdhu3eHqs+wnsJAcjiziqo3Wub2+KlFaSSQV1ylTbLnDFkEnzbX93J
LnWNUbGX5/dI4HpJi76xHaydd9D9pZKemnG+eFUMaZ/oswPiDUaYDxR3mjMI
bGvvzu6vBs3ItHEJIBbOpbK1LiterWqm/uTThmkHhjZmjRCdch2bHZ8Caky/
DuqGmJ1SP4ylOh1VN1gAYWHhF9gdyrX0t1tWmzWP51LrVjUCdZKfQMyghfI3
JkwZpHpV069EUlz3Ud2EYzCANQK4OB66aC4UhMC3ErEY3+b5c0YQOFbEfUpd
34zOUCSonsWB0nQKijhkE2pLIjHr/PbpMhz+w84/cobnsXq3bTr9YkHywwea
SPxmubOsQEiA4FOA6muXcQEPITdw+LIBLeFG8bmZFVzv0hyt5CEwfv/TDPxm
Bch1QPUDpsXz3IYgeFQp2FdXiHN0fLlhcZvQQ5mT3yX42RD1Ynio8HoqYMT8
ik4PKv1CMSb5Cau6v6S/nzYcOZ4Qx7a4UdNH0F7VxXg0ubLObQQdd1boXnf0
iNdTD3sdFimpJag2IRNDSl/ZdGaAa9nIJenPDIqz/km/DoevQcIFfi5V/cQu
wTdkKFmaVzQVeV8/skVaMXKV78/ZbC/3uXX6ZFLyv8htYjDQeD0nWXhyxYwq
1ZULTUKiHnnq4H4Gx28NzriBDzC1GXG8ktbauvKyaI7CgAfqu5tfJVBlOt8n
613Sryun2JYx/NMayCNpQyARpwDsg5U9iV2ECFXFutaRZuZbUp/szg3rM9fm
+hscMOLZNIp3QvoIG0nGTF+8YY8xEw9Ko4Cdgp3Fk/tUy7WzkwSkrwhBEqyf
gTDG6lsS6PbgK6k12+4ewCVPvYh4o6T1KZ/rY+zZH9sqCKoOQCVSlEOCMFYn
FZ8np+PqziZVL3BzsM6M2c2EZbO63l90ZH9KITuTuUhKBFFi92XR0/tLKa+u
X/s1cPUjAeTr3PyeaJ+tlS10LowE9Sih1/qd74T7EYdVrg/bq5Y4aCaBitzN
IpQhwJCKIfk6nqEnMiHDJA0q5JsZc8zVEC/DItAyvp3P+fN0u3NsRkM+8G5+
3gvu/oXpeCWPmazhpBKDO+kBQkSv4rkdhk+krG1yJAskq3WWNQTx7YgTyOyK
9W521+YCiC3dZqgnR1HVbVO8WxWI5c2PD2yXFGexAe7JHx/K0x/Q0MaB9tMM
0/ZwbkkOgKTFj6tM7SSqbCVWqhDhXbZ+ljnM9Fi4qqmq4jzn6a6E7t3FsCzP
qwUjMjsTZITTMWMVYauS+nHHvYmtb2faqOq778q4JsQo0Etr6XX6JFRdnTw9
bGo++/uCizBcQxGfaAkhen1m8WmnHhtmokGA3Ys7PjiKkCEVJCA91jXiA9ty
G/AInhlN8Rb5CrXUsChOG5h9qsQ9szcYrxIE8sRb62+j8OUduGaR9aWu51Ae
NDaU+Ym3f2n82hQSzijqVVG4Fj8N4PMP7W8Qnnfn6v3b2UzqNbMkdGiSH7qA
PZOS2elBgfYYHyZUtzpKA9XxfnCCrzvcWATsg4lSQbfU9XkmfZWFVekNSRh8
kAIc///PkaxHHfw7VDGO4EPNy/C1bLRIOfHDDwsvA4dRR9CVVNAS1o0Y+ceS
6Ac4q6ia+SGhgNWBgOFrnJ46ESR6VxGawTuwJMZ4wlJj+kj0RXf4TyaGwfJ9
kfo1LKdU6bZXU829wqG5YE7Lc6NE74NSPOFkWmWtcEsLmEgyIWna7Q3dzhIt
WEgCWNyiVpHZlEvgUdpCpe3yK7ppdHA03o+gdl4YR+LX/2TE0906p1eBpe+V
8N+m4KUBW05Bo3sugy+2hojNMzyD/q4ADqKHeIqiDUKz0T6eEnsfn7Q0wCWz
3R1VnAkRpF2HC42BQDKmATssvJNiHxQGTmVC9Pc2FvQmQqh/KgDMADoHSsKg
zLIrFTTz1bStoaw8XxDP3kw1bZzEceL5j84Ho5l1P2efleHNXsaDGhaYTBNI
7zJcy+8fEfUnJm4a0KPuDNuWJXbyBh6NwUa4yey9cOS5fXTYhrabt2gE06C+
fOpqn4F0nBZnJZWY85XuTsszRiQSNujW+OriptzfRqqpxNDlGc72lseg/37c
azNiB9maerbsY1ut1lb20DR86FKEW18v9VmIArjTv3VfVSi4U+0qeGP1fxIK
5orKyCB5wX1tmmTCL4/qCPgnnbwM9KU3o5k4N1App43oGRWzYiGaNQY/9Lp1
ztPZFkHsaZgfjutGVtihczEKr63nZ0H2vSfkrVeb2k5PsV2jvoaIy3i4TdTx
JDmuK883dmd1yzvc4WZVmYR2L5RQZnAfl2b+uhmaXN7fonIMz+qjrPZCpOxX
FpbLgVfGL8TM9KQNPmkBqxvMda6VraingfUifvCgWPPrEhKAnMp88ZI+JekS
NAzcoq0PMSSZVlhPfBYL4qUW9rTmwqxB+xo6YNt6HsuDyKS1AxlPmpzmoCvk
lsxdu3DeLMNk3JDtuV7Nr8M6SToSLMmofJnaOIjol7GzK1CUm2ZoP/TKU157
F655D8hbcXGakYUklZS7Hj95FN9yGXQwBnlLEiYeV9YXa+i3e8WlBiquAK7S
ec0V+C1CwsvFJMtQzv0RMJl0szVg/ENxOD2oty9V5cWGsUwFdWIgLaCU0qM7
7ZJpsI5Zc/eX2orA1PV0OCpgA5eI8f/rdAB6tKdFeqF/uBAvxN+rXMpJMYzT
Q8AU0nFZjCX4+LNhMhXNVOLJG0Mkr74VQmDWsojbnFp+ugUxEuIrxyJl43TG
9mNTBKAwuSc0gfERoSHedefaqwYespE4b1CBrY1FSeWR4pC+WUkmRcvuc0uq
0OecXazzjTpioR89WnrBAv6UzWocnBKewNLjCTGCPUP68Rwceadlx5P46KMX
G8yB/BhsvRV+qV11TgpnkETbFVx5Y9AI5oLL/gXl+xaNTqNWCG2yHbMU50vf
IYDTXmIhK0gmRSMJ7uivjBBBE3aPJqfwNBkv97sO4JjOot+t8cNUPtRVzeVU
/XzBPBBTR9gMTTzgK+psj5FYJzJAO+bmkHriLrZlcQXvJ0v9LRP3l8EGYQWc
3+JJ2vloU1/ue/N3au5bUXuHz35Q7Vir+xR0zZBagoChdE84rd/y6vMA+okX
0M0agMcudsFFKgkAPaIKqEXq5vRx5keEDyrxjSntFeZKHO8CCZxJlQP7J1Lf
VyaHQ4Xz2JuK3WuSvUbdLoft4iEy1y9P6RoDswybNinBQNaJ5JO0KPAJ+QiC
iJvk8OPXeA30pMSOZWl41wp9cSp+S70oT2RRXrvuq6e8iF+HqdDoaol6i3qC
l8J/OKUpVEK/bwAL/HyAs2ul1FmOfuoaqnj/6ixWYbGBO/paJ5AX8SBNig9A
tHkhz1pS8CbdMZnoIJApk3NaLE6uJf8qe5tgXILA7VP6yF83S1mtLAIXkYrF
7IVg/KpdDLNSVmsVjiWLniH6fBlSLSBqGHASTAsO5sbVOI0v7CYij3aI7dEL
aBF8AjZ1/qEXXRql6SsIA7sLJjZYmJPXr/58KDOiFmVoF5xkYxM38uX6v8pw
OXGDBJP5mBcDH0aUQQ5k9N4Tl3x8EfjSg+bRzLYco4/jaA5Tz7rwZhOcmeMK
iiruidfkPZCEbBOMdKBfqWHx1ZRdGobhoJAPsMWYH37Q9JLKcNmsv9+ih/rs
yL44hniIoqcwTOiVNer3HXHKY7ovbcp+lvdoJmWf8MAyrteFCpvgb03/BVud
ecZqxe/Jm9GE70qzaY0Rsdj5XhzuZrC41i3yXRM3nuPO3AhbxNx7Ndg/IeA/
WVpJO+2uAYhUiNr1H9VJjfNG0m0T+bIi9xCTwj3Hp1gYnd4efcwB0bmbjEev
6FAaSc0And4PRafD4gqSwi2Ckh8RUFFOnzD/uRSQmdN3aryem8gY+R18i7Tw
yQSugpSvNj4yJDngwLdZq3BhvUbpctgfh9lBIORDg1yio5j+5vmRo4HB7knC
/R0RuexZ/kJLr4RUZANjG/Ll8eNx6dBS4VlTvAglHhjvQk5Ds9Y0F9Pmuo7k
VShyEA5++nWtaDiskqQQSpG6PP4jE3AyXFRquTZolpSo8Nb/ZRrvTnBvHzFB
wtfAOi8zD8gDv+XyPB2GXr7bXRIfEB9bfaopNiF5gEDtrU9rDf27RqKk/4ba
sIe2lFnb16PBDoMAj0SI59JKRLJdCnnh4WunrAWXw5ZCJJcryTrqJzmWxPCv
PtDePkWgsklf3nz/ycoSFYzpUA2yvO95dNp+fR3gDQvZHCKcjhlyiMS4kJAy
kdgxtvnpUTvziJnxYWyIgJ33Bsk2dm70cwXsBfvmncODj2ItU/Xvb9ltmv57
6/Ttpi07BeZdmH8LfGScv7hw2bVG/xmv+/UEYOFAmJra2VjfGUKIPJFU2MX+
pEidddhrPqRThlyLWgf9PjAWW9LRWXwRUacmJUl30x/AsFRZRlozWmY8Iv47
YPuC6G0y8qW8qbWYISKII4iAv3fY9XXpRYuIeno8xYaWFrjiFaXPFfyuYRR9
3B5nW/D9V4AMUd020VPxXdPieSHzekk/mEsZNjUqQVu5bIWKofbWKRRFRom5
8KrX6/elJclrVuY7QgRJQGtSZBw6DP88Ug9T1IrleUEDubslGxyo2c0QofA8
B28b9Y36d71wLuPzqS3nvG32juA+hhaMJjhAOXIG1Us3XwORAoQrmJTrJvbz
nIenmfbVniW5H7x2+DYNUSMuj32motKqkWo7sK8s6O3zZ2wVIl8nPxQ11l9W
TS1sSrNB9gwaj2RjEsM/HC1FCFrybTfKbYixhD/gVQWet7NvG7/ysOGvy0op
9KGuNiLSZ5SJU6uy9lfrus71YJc3hMJLqanVDf+t1yMg1eOFByvE3wgk6xlc
6Mdb9xrXJiibnmcs4fOS0OBbDb9Ug7QjbmyTzuXQriboo/kFVUPGd2OZkkSd
9QWSQ56QoXkTKDeXkISpjla3DwJAiaBaWpm2cnqg84sS3wcRcrDhPhvbtqGW
00D248M6nSHOyjd/qc4Hy5/FPZtOMFu0Hui+Pl/PikrsN0dbvWA/k8s5k+Nt
taZQraGVyI2YqeNZRucNm4MGfKrmEL8NQQAYm21WVx796y3RDBSaEs0MSCrK
abNrueNgb9vVl5NMSVDKU5cGOwHIWYjzHA/GWzVdmTdIDiC6Nj4QPs2i7VXf
7xQCx981smu9v/nn0nt1MZPXqF0+7qChlITC/5xFLMvRDHLG5OoXAjexjvUK
qJRyPypNAsxt9pxY+zAUTKaFSLXUE/ahGFGn+r823+ynWdlUZcH3fdhbZZqn
dH8aA3uEQoiGxjiSr/eAhuDB5zt/nY84ZdqBU4sfudeaA+p2aTQ+aRAsV3It
u6ww4U1ci4vqngYaYk3EgOUFAdakmKQBBKKel++YQMXFUu78gSCyI54mdSOl
qQHGEfkhJaiyi9oe8GTJcwb2IaK9D8SRNCq4QDN0sTbrmgf05EpO68QxwSp9
h0gn6B+hb3XFk87tVwc0+a5Ye7MOUnpkHVzb82X2+EA7gpql7I3JhXCqvEzO
dfQiByp5Nioq+E20ts+89bGdATY2Nyq85z//uwlF2EwbrvGOwLm+7V3/Ln0a
d3TL1v1TVHT1hSYZyGGkCx/ZPdU6L4teQsQ/vzn5RRDLLoewgK7F8SpWk6pt
ab03MwAvzD0xEHCWyWn2lpTou9WEjqhEX1TXV1PkFfxMQca8P29pbS5J9NHC
VV2cxcjvwhrbUXCbTWaylKOGbBA5osLzErp/8nG9wxaTi8WsjKWp1Xma6HKe
p4KuqD63An61B9Rsrin7N9dbD+gCxxRdIFZ2Rf4kk5nbNkqWrWnoNW7yA7b0
ewzW4aD4SNxSLboAVERia0GmC0Q/EGIapohE82hH5jyYwIJYP4+QZ4Bzr+P9
SZOAiEsh4Dq1mTvXNZ64/jiRpHTeM0skVmdaVqkL+lkywOUjpMFqu5rq0b+v
PAcIYz1LUVfFmYskjgsXMw3XwNMsP6YuKdwTULWOO8L7+/1dzcrVVYvF8EdI
mPoOoCJDFaU5SyyD54NJdoOTuB+6Kz01bOkH3wW+ZVdKAE1A1SLJW+Jkrz8K
6vbQRyxCsbZ5HrisJR1v6gKp8zDv4p16LNo+2PrfHembHnbWBiz8IYbuimas
zGrvE84TlAuzY9k837spQaDSaD+mbWcHmHNyj1pJ8/EgZJON6SLbPSsRcpjI
ZOK3yRO4gljTYfkfWtAd8qF9HPf+Ex4i+p1oDyq/MoFciRPv5LeTfKTj2L3N
HG2GiyRRCoN1GafKDfMdyf9hoSgLhlSyqlxZeNd+qiXZexV0G0VaRfAambGD
hpmBcpbuFNf591gfLka4BvORYYt74wRy87yzzwZ6acW53oqr8N91kYGhbfdo
M4am+QfTiQ7UZ6ApS+MVoeONfuhnWKHMC5N7hN4xlheudfv+S1VIMVcjPXWW
cb7jj70ubN4wLiAedaXyrjjxF2JfenwWGiq3FwcDsH+mRmEhDrcKjwVVggMa
x449RZkiPGhvBmBix1ZB8u6880w5tUIV5kXl9OApE+GHuSKdwAyLZu8JMcls
B80gXMFplVN1Cn9mHEiif5VD1FXtuXaugSjeS9sKekde8z1u0sHQh0TpQFWk
0XXQQ6bYmJnCvEvNwhRpmUobTv0uDJHI8J3xx6fDB/zt66w1rp+PK+ffAZ1l
9ne+X4k/ld+fvpGqOU8FdJt2ytb6FD19MlZFLKUxFvR1nC2FxORGfuBlkut4
5OchB+5vs26nWC022ueojGwEwtNs7iR2tC3gW2tGMHO0ZMhZmSw+kzvqm+C7
OunvfBtLwQNV9rn2gtfVEKg53Mwx1+/CIx2ekggXorX636b7j5s+QxMah7JI
rQq6V9d2JwatdepU3Rsd+w8aueep9ib4mdNrFXWGYw2cdWHg+sSs8/ePuJh6
hXDkmgaHH5ruCXTavOR0tjUu1Dpe8BUt5dHi9cQ6H7Gk5TaiOvuhFyvOvnEH
Mk5Uzh/DV7v8g5mOPrKj7FOzSwppY4vw2OcNnuNu1RGqqg39qL7w7osTtaOi
Q5kihiU4rGaDcV5jq1BtMTepG6Yjylcg/AGAKlGOitm+yyPumcP12yXGwf69
cWT6CnUE9XISkI02tlWOrdmCiAcPh/0CWCXXs2ssjDFAM0s/d8OjpwXtM05L
z3z5Ak++XKhOUYcsJyAVEU8xF2EbIQuwOzEdjFseBREXooU2tR1MQTZopH6g
35em19NY87MIH3k2/yPcVLDzl7qUlQCTIYaEU5la8wvyq8SOs0XLTvgy2HMN
G3VFasWVhV/Ddcxt1Gcwr3k+SzCIwrifErdcz4pNPIcRW4p1rc+b4lvBn2w8
RlE0Uf9s6Meef5FX8YX2Rbxd0clnEFbH6tH10K9MOXWX91WDyyqaMbULAFo0
5tOiz3Ckhbp/GEnCKQBv66UNpe4bs/4O+ERoN6bjp1fsr69wii9FkW84CzX8
xTRFSmo9Hmy1a3HgQsA7uzvSmP7+g64vA4jGKdyy24NgFFe3a/vTj/ER/cQt
5fIthxzoZ4rvMM3pVK1c787xlS+A6VkbAK8vu+rg0N7ALN5cZ1wRB6HAfI1W
hyRnEAvD7/ytDaV/sWc9IZ+hKRs0WmEEK2d+2xVXG8l8GCex28bJ/oMNKJj9
1iKWY5c3n/nEtWn1udT5IOUPtF3VjGzo+ME50cm5spREOVKoOfPijPSqSJMo
GtFT8nJNfK4pptsp3lw266VkbYD9GU5JJFzSfPd9jajT7nKB1MLEmTBCIeg4
7JgmB0+Z+CzNMRx99qui+i+ACR+YPxKj+ELJghRCTDSp6JLjXJk09d15Fivi
YX5GgPSXZLnctyC61QWDnEX5k08kWaZm0g9I0RoitlrPjwqrwSq2myRXdPlY
xwg3yI0Oa6gLyCYnlmXYcyV2oBmoT1fzHpcjO3A7lsZPRRvxKZxFSxw4hvdK
jzcu6nSIY/peCHXjGOZKsBqIxlDPCQG4Z/Knu0AB/iYNKiSoS3+U8yrsI1OK
Sh3g+DbdIV8c5ulLVIjVdzhUpn+x1hv6JN8QW0hA32u2DLV0+o2IVu8AWTdI
iPLT8NcvxTaGk09Mb93jky1ifVjLEUO/axzGZv8R5WwgEqvKstGYWLS/EeSb
V4Y8oUI6sjPH+dXSUglPWXPc/L+wdwOofN1cZJd2JAIUlg3/tmPaSPsgVKVC
hGDu3m3bcpoFwuOCVgGWwid/k7WMN6Br+IN9VaAciwEk8c6+8dOCYVzjZWUN
KdUiPqd28nPAHLxgV5RtimykOpZWUepXKLP886oTxhUqWomn3fX8n7c16bDH
8Dz+NhLt+hmSIPH0+rtBxXbqiaiAf55+ceKK9j/6mWkqZtdTLLx61wWDCGdW
hnFGpO4nURdVfwuaGCiiWYctrN+qhC7z+7NvCO0fypmd89VMNawllbGAjh0+
mmLsKvFLQzljDIag/ijgnrAqO3RTr4WghEPUEW5qqAgSp5171EgaZpuInRl0
jeZHJ8fzFBpQg0+bI6fLx0cx+1SsPHUhZLqxl2X8CWp9JaOppIbvdl2e8Rz3
t41d1Nm0W4GJ9RFkMqc0c5NUGI0s7cRYvoRETgv9NaHf7Tuy3EAyA50DsE3f
oVpu4+Aud+UyUd37GOALS71ja+Sa9FxPFcFuetvGeBVurz4CQef5wLRupNVE
l89SX9juxDuwzPo27+cquXoZr8MnAqFyvlfdTlLT1cw5t03JiBrkXuCo+Jql
Qr0W+NQyjkSvVyiVA7cDsAkxBDnIrGR6wSrFnLfRlG5i8Thw4du2hEiLa/a8
4cJcxbR30OFD/YdbckR9FIRRpaPKmSz+WWdoMMG7p9xhIq520w+EIUW9ZKp8
HqGW8eTVFAeMKxodriK5loCraCzSfaiEzkpcJ3JZBw5DBF5k9KK8T/bPGZt3
paxk77o7nToO10IYJPmsoWbdJ4weppyD+UR2qVk8pGLxsYlIyb3kWNUP6c0u
F3jdFRmvKXv4Q1dFl7J+NVPCz8cSMPnNcEBQGw3S9KrduCq2JA6wdR3XbciA
nt0aHfWvfNzVKx/7g3o4slkDK5I/eX3IGTwHGVy986XGXJBWsqOMlfpYs+YZ
IoWqrz7/psWTlZy29T7LjnkqRS5OI6f8uXfTrA9SbHlX/Sa1E4xj1ncT06EK
4UUlXh45fBgeV7d3vYLatJwxpOXwkWcH+Eh+rOSy912Q/wSmKMNbBH08Nx0e
dOuw0hhK5e3mTL1y8hR3ef0+8YE2Vk8CliKqMJvmDxylZb0kXjm1QISEFrK/
MXt2JCFxvn8XZBzYIRHCUCAbvGvD71q6yuLmonq6qZE66EGGZKlgMSYZJkDH
QYMaYJJwaHSo5PHm4uHZJW70+V/bFjAnU/+yj7bxRdKmwrnOZQ4hB9v+l0Xv
kt2qpchbrKZpRHs3eIbb5rGoSb923NFiE+FlaNg51nIIX4TrPvjJAbpxIzhX
9dP6HhGuj93AT9janl/AjgQUKqN2ifjnTr8BslVrfNabgDzhqRoB5j0gdGYE
aZwCH5daZ+W0q0HpTTK8czcVy6xnE9I3E2QdVrbaQzyriaGOn7gk6qI7QmPc
aF6UDaD50skzHw6TT3oDwxgr52jzD3a7CnRi0rtg/L+/wlSiQQa+n50dniUQ
dEbkzSEFi6QbblB0ZCA7K0am3EnR7L19xQuYye5uzdH04j5C7sJFH9rHXRgx
iFaljAk0ZlGOF0nj/kQPI9EuzwUhyGmnS1LkNqjV01n2jMjb7RfbES1KLA0t
/qvhJMJs+2/eF3BHYvmPWmVZybFiSZUWbxXxh8kQbXV7gMw1rsHPrXZIoL05
ydNQ5pSbvCmgYkmkbxNaP4uN2Z0R5oo1iUUeH+Bug7yflARDbYzHv8myv47B
c5B0VtXDpOsgkkSLb3NVObqS3KlMGLH7KKqXHNFR7+xz43ct6KQeRvB2FYqu
ACwR28x7s2vn+SeZM/g8d1CzAHgniM3vQIZPEuCMwPFM4m3IRLY+XB8IJQeu
g4KLobTkHh3byt883pE3AYW1wizQt6Sa2uBkZwG1z9dyWxXuLmL6oHIHaJW/
n3SabkbpsK4BB5fE6l3x+pOqoEdduB6jFs4ZMmmtNC2z5j/y5+KJcnnUly0t
C6pnOpqHTWGgIU7c4XLqxQEoCG+w1by6gId6DCSEY6Hhcm0cxvT7jtEXCmoW
/wJUQrBHHYk9rPKEL9eBMlDBHsEG3AbeXrVLePdcXMz6iIU4LX+LflaqzYDn
drw9zbN2KrIT4L5bFFGBevzvq5q1mYJthhlwTlaU9lqZxgJQ7sGFUk5r5//a
1Vtzrb8cdELLsn6unbSxFmrG8okb/nTsCclw/A5FZAUPlwGfuSrqI50pB01F
786XzPTsJjzRlpg9AovVt28Py+LvzyD62bMDCSX2oa1GB3dZnKw2RTU4ipiv
8X8PFtH6CVxbC5JuF6NCOiqggRkd1KaJLiTgOT4KuoxXsmYTYTmqBEtxLj0o
pPIOVwmH2kW/HvLTF0P5+lYajItzXG/gqPAYwVB4Qm7h0M8VP7mljp/VBIU4
RfcBXTOUr4DGKpJaH8BX/k97/zpyR+AVrQt51tZeYM0zmGxTI3Wg/W5qyIIW
mzsj1Sf9z6nzcSVgYjOTcnfwebOK2RnsNQqZdIvThC9p9EhXDGbdolAUPe62
ySANYiQ99Zt5y/ZU3xVcNhaFA3PnNdVtZahuS0s0kBsW9DYY2nVBkU1XhqIy
I4kS3tRF+03lvcie0+0QzRfRrzkBluW94WMwQ8gLaPU953S5qF8/NZkhnPzL
hR/OoKSOnZFU/i7ElG3pMZ1ORoOBOiUAFFw11EgovHARmKEByEk1r99jehUK
43tamgpXePF4ZZge6JHk/CxylZT63l91ylyJ02bH8TLdLNaYWip6wCELmhth
9hbJ48IJM0cuKRWhKhf+ZjdXEQCJ5K+rGUq4TNrgMmKXrP/9MNpmmRHezTM2
Lhr+e2bEIBDQWFehf9oUZIuZBSRxJ4S/iX1A5/KykE7EAa/j8iNPZjCKthdd
986Y+cJPByZb4UZeXrZmceusOQDMChbRQIgrljPNo8UHd8eRiriHUjSKLXav
4UspoGPgQMie3N7Jy0nMdb1f3dZvtTMzQaph2JyL4Z4EI16SvVHBjMW5p0H1
HA0zNFIfn509cnDGjxSiYPVKxmRi7hbyi4s/b0+gR/Uo+NIV3yw6nGWVGdrv
y4slcOLCnDUpy16ut05ubYJ7eCXuLMLXFiQqcOh1jQUHTsgm7unUHLyBCH9N
TxWfM8Rw2lfBdH/RAzpGUrkbLRCcZr9ULqZIEXW6GktpfdhpKaEQ36XKhgKV
IlHwq9mrswHDRju9OZ4hB0Pjcl2li2mnW/y/TDlF6+v+dK24gleYdJSpDX6W
wWShIPBuC1DDKjWnZ3K5Q2Q6+HYwqZaGHWvqqv/y0kVpTFbOv3wpCmCNwrwi
WgcqkQiMpt/cLpx1pvwO5j0bkp5OECSOp2hqrYzWUftma3dnUFBkZb9IJ0FQ
tvhOT9xyRzCW6MX1aM1nZmzXq+5RmELIMA+oUyXvzbcfpbib+UOJzBK96hpA
2bAjzcXXoytkuant3LEsLZ2ahjorrWr3VuJQeXA9K1dJPNk9Fy4eKacK+8FA
tsInZwteYDE+lQF58nkDeV23VMBnl5GiDs4i0zQNPdlKISmj+Ty8yk03TA53
YU51P0jI0XiU16owaWlMBWDEOb0HOokVNyYe7r6ozVhV/729y4XDNZaeNLrZ
Yv7+q1gHObVsyC8LKEXSSTepvOx1qt4MD//5Vr5uIRwNYClrljBCUPwOSLjJ
bcfsfQHknj9hZMogtlTGPKXd/aLxNQh8wumVW6mSdekxae+jXCpEn3bpkheX
TSPGL/Hva8rrGF/ITCzjfR5hj5fMNan+TWiTJuYOmqVPqBOo3Xdb8Ll4d5AG
OmXaxBuvJFx+6559+Yg5ZridGaHjNfm0arMmTID8yqXx2JN7QOAaz9qdD0vx
z4HNZFXGSpUMb+7yfS45+LyxDHptmiXNgvAnwhMkDVvjjr0OYKn7VljwS2aO
VwOdO6gtnC6jRrKjSaFg8on8xaitO34QNSKrKcNkgEAPFtApvT6UNPXSDWGA
nr9FvhGmgjjCurtaWS8QkUh7OB9aTT+xXHqgfLPUtYSRFP803R1nrY7ekt2r
77UuLOsBb5rQCjdwEYjGAYiAtFZC5G0sREYBYplqMPqO/PpNGTauybrXz1KG
N42jx+wTwdFiDuiz655elFZj1lsksKYRqX2eJph+rD6h05aN7zCflIGWDuXT
bU+7AZ6syeW4hdSShRL9sz3uT5dPXKhMQ61ITcCMemrp1INH4f9EdLTlmPrq
ozuB9RP7RVW9xxnhGwAPdbZhcIH2v6DaElOprxuDclxbIe67pLesn9Q7Uwbw
IO1aCi6/xEcSzDbTQrlnvwV6GtwpFxKb1WE9ykM0iDObKJLA2Y1/W/1Xotki
yeU4YCCzuhKDlXuQRFvkQZT6r9RmekSBOl+ecwzXdzd/4cqeNvGmEuBfTHtd
1hohG2Lq148jp+wROMDIozjy4AqQfja4pt53cD63w4zaBPeVPMD400cwJ6Wd
uqmPRdfbgJdFaUb13yx2cycDDC/rC5iDHi6cNA76JviEnDS1HY0UAxbC9S+u
ZyS626p5a8jhzbeZY7LvlpEcjkq/qrrDQ3q15Y9y/A424z0Qtn/XGjuC4M/B
Gdylelw2z+kJNJ9CdVW60TAKUo676SBD8VbOGOnAnqePdl+tHpl2GIIU9kRX
xOBE2CjRevDdg0yaapPx6DDRMsi7+bg5LMwo3eMXTp0Fb3EgAPyQcEQpsbjv
ufHPzShISpUFODEjhS4TKpEBub23EKea7X1petl4GkjxKoMkvOBJfxd8o0eD
bPC/nn+1JNf7DuiCwP+XijKZR1iFSOxfd4TJ0VF/QnSXaytWIuJC2i8dHbO/
hLcaxezb3nhl3XrWDF+FbxnWsdWncIDjHL9lL09iSS4TXQ/UR0NTDnG0dYUk
SBgsVnkLNGvFt2YTxXYOq0hbTSEYiZA07CU1LauM4QgACeQWVOm4WH8Iy33f
nWWoncgPjQHuyXNeMU6pM98NeIot3wlpNiGFQuByYO5PJmFSQW3JgoHgFltm
AaqfrAP6kiGjkxw0dn1IdfNh9Bj4AWmf3aOTFNDMplBl13/5wk91maXou5fo
Kdin9L37gaOGiCGHV4dU3qaJjE7fV0T3cn2m6velpYRpurGljo7MTAf0T9y3
UJ5QQIsWyR/K2mY850ECxTRtttyH8PNTzxMUj0/M84rue8AtgR5Xkcc1YvOd
nwTQqiIwvSZXytDshiHkIMfTdgEjdMteeUT8zdffL/qIOw2tVRNYZHANvILQ
TQ8pz/EruKtiyErR63XWfOxPMnOOspfPVywW/HP85ldYls/r5JkLCVoydfAr
OdctdqgLI6L+dKVMtiqZj4Bz8crjxJsFlnz9F5JAn5wJWDiO6wvBnbarej/U
i9lj2ffRRAR0JH2CAP21TWGBD8dziTHUs8Rfb5RAotvi5pZkmZUjeXVszwge
kIrv+XfaAC75hClKc9aQDBsgFa9hP/rZNzhqmfnzDDTVWEBYz3q7XDFgN/9d
bou8Wu1VND6U6p3uRgqC8fKS1GP6sQipS5YPRGyBLSXhcoATg2FjqYeUdUs5
ExRl724nK/ra9kWCzmi6akn1CQAu3hq0zGr6ysns3V8Z/06biZ9NuCv4xzMn
zSbwda+FGRfBZygfBJIO2wOGL2s7Ca5/FJYAqyeJgzxW4leiTAWkMmKEA51n
ucPl0hCFD9Lz+5v0ELwj7kapP0Yl+F+FJToJOaC0wfZM900+IHZcPfvqQjql
XGiLO/Epl9Us5a5sI+qY+cF9hhLvzn1LyZDK1A4lgcGTBhSB1xETqRAJP0lS
Frhll8UXsH+2n1bQWLR8c3ohrlJaw1JBL9MCS8EsRUgd92Zvi9s/tzAY1Lcb
zl2w0bpQu83tMewljU0rlReLiXFOuawJ4QocMBGQ3U/kxKDf/n20UA0SciZO
CYApUWanVX1z2we4V1RDc430GeqytxQKpGsS1LsWw/jgJGstOZ5nei26Mm8n
BCmhCsevGOt5/olCYY3ymjd3xQQarl0w94FDh+K3DRbHwLxPkOwiqXTxrjFt
R0NATzjb0z8rF0ZzkYzHtONnomM0taGpM0t+4NXQud5WwwJ4rscGzR8/d6TK
Stqs03x981PWNwB7PEBWtDwJoH68NieKkccWPaVYuzyPX0PJqhNyjkUfoS7d
9wnejOEcHHe4k6MaGh1TDMz3yZLl45iX0O6Hyu69RfNoPsdxzh3tbeDRKAvc
aKK+Nb9paVGIh9FlYRNGi6uazJfuSrhlo7QIpw6vo+E2CHpMsxYbGNJTF8BM
wbwkw2rfSLoYjwglZCDw+C7GUOSoJaZDMpt9qw3lJWyaEYsNVCeGW+zfA4kE
Zm7sg11HoXVVreJHiN0MvzY76ljQSZZUt/QIl8YPFwJVFpC2J0RKCXa0DN3l
oPVzYzqG4hUB5e/hL2JRgmggtahQ5aIGa0xeE8rPKUzBKDJNnMJvPf3iKRZ3
TaQkN7irs4+cxqW7eS/WgxrgpzEEgaJc5ByV9uAmydzqtLne4Wy/Wpy+qUzu
69HOIkLNBa2e3t+88qdO3QzwD6uGHfAAn8RRxm5Muui5d1b8CRhjSFcGilPZ
g8Jn4c85YY+OYf23kX1XUqk7BNlNY91EbrkbB7xNfJI7IKK7qO5NXT8vP7HQ
wKWdVruBi/isdX9BsqdvyRs8alL1zv8WqhtQnO9H1RFTxm7iUe8fKxE/McZ7
khcuoYDwOSUX5I1GlK3fiwJ4vilRXy659Rfv3nLzFK5sefGh6zL8DU1EqvrY
Njgj+39pHoPB4seTTe1g8fCKZfuw63vwmk7T6h9fcOZdmtf8q4AAaID5xle2
o6kHGC+esntcE8Qh3WWg44IOtYtfFXN7nbYr8ubX+qaQ35A7AYeoiaROlQCe
PJPWxNeIe2M0TYuH4qRBF/e/wwESCX5bMzsKpJcKlghua3XTFD43+FdpaOqG
QoiKK34bE7eAdow/AfJ1ELZRYlv6KhehVBv+wmQhtoDcSOifqexXWm1d+Z89
7gBh20zElg4+IrM8BdQQc+sM9f6qMBjH6t6Uky4T167WqiE+eWirmSuum55S
HU+Wp5k7ksP86+lLVruNLchlVUIlTm82upwbcparNIAz30xbxtrGRBXEgb3h
MHzQt6Uz4Pri+4GVtN7FfhMFTHUICUPInJZ7pmpl8v0JGZYh+AJPUf4rRDew
JNTZNlLp2fKOvVzHTvbUlPbjBITXs8GsPnDVzJiEUGNU6i0nP/EWi8Dl3y1k
CEP1TVgVk2n2M23nhTEy0/AzCoVCda5hAQFLREZZRTSkKpVN0ggAu82yd1OS
T0vZWV9/QbKnHM7FxUTYOhFiAsEVK/7BW+l6yTSI0H7w5YhEecNdL3T1DKO4
t0s55ZcJ3ir9+NYY0nzXjdlU+x5tKUW76rheVincL5CAiQ0qljWYgrOVCNFh
o1cxw2M6Rq+RLfJHt1N7y16qhiwTUQ5xxWaXxg3ymY8U1tqs3kKKdojvxYkl
bPZ8cAvC27/MGClUn4oyGhsoP1XwWBjazD26czYYdx0mpjl+UMqJgtgeb1vU
m30zBMExpSwG4AU6ZWIrfvaIKpQIFTI+pkuVk6NDZvcxCTNzLxYOmimxWYZT
R5vn6tM4RLL2+TbMe8up/+eDnjz+PD9Ukdj/sMeVbRGUFIpIrabuLmNmae8G
qFoobdxl0TptxelS+F3WYTKddSeSNXjI8pzhZ+zRXXgwe6tKBui3Ro/wkmXb
te/0GvGUZ5gh0H7izM5XQAz6PVtV63rZipPAFWOzvZlWBeOd/WSv1H4oCU71
2km8WFcI9xCSghDz5Blz78kLSbTr2+ZO+AkHxa0Nz3IiFZHp5PxIm/eTSosc
n7NV5bU1skId/cEFH6r9dxhrCGiQ3pUoH/J4i6zsqHgUwwuNZdf4DUo1gT6q
hPO7QflfIZMzLveXFKjBbjrZDzICx8IMrMQTMKz31nk15VgiZU5QeRJCbmDr
Qs5iF8llAnY8ejqYUpY6NnjEE4ciRuk+TA1Ry9r0ZUjIsRm8zPBPuklPnJmw
31ZLGO4fvpJnjoPZ0X62wZYgF2nBuis+Ec1kZy+bvtgZzAkY64+DBTmjSGhH
g0QgkFQmHVwWzkOB1qbm9S3hsQ+Cxslqrc9DzOwfBvpLkAXUYVgMEr0zaCwf
DXGg2+eP4WQWs7U8g9dia4zbrfDW2o8ntyjDwFD78BUMQVOaQTrf9nLpes6C
zVa5n7TumBwvYhW4amGufvXcQxJqi4BUp8YVgJO4XC57hSp0HDXwtrbdepcO
2m9Mm3Bu24z8Xdt+KHW9/m+LlzsCM9D2pZbbBvBgXGoqriAGYGGxIqRxISIk
f5ugt6qr4AD4BWCUHtiwnYHu6FxtKnTIXc9+xDkRiL2eDxWtWQBSMQnjhPWM
VjMzWUJpyBkZ3TytO1CH5gyFZsp52kOGy4yshF4iITVpcZ36kfDo/MS6A3rs
UIEzyLuft60evqojPVlclD5dkwODl+i8RFGjsweHis0bTnQpIZVFMsPeQnBR
g3Je3R/quj9xWiUVAaP4tbbiDuX67JrXF26DBI1X2GCK/dbeDnV1+ZVQKe85
mayDq9jQWNx4bYGwa7Cs2GANtno8BcuCphEJt/2u9vPyxmPyxFC2H05L5Mna
YiEFTxjkMRGManokTId5kQJNa+moqv+6aUm7+O2YyXfd6gSUHYVHLUAzBv0M
pdHvoSKd8NsRQM8feMSXjk+pcliQ7/If+oyzF5FHcbcnK8oim1UDEWmCLwDk
6rAcVU2ahxMCwcjp6agnnHMsq0+KLy9CqL5Yl6zc9xaViMqOarXVN68oFaRY
AYOTKB3Rv+B3vwJYUanpyOmGaeLjYaSnj4VC6WcqZv1YnaMMtsOEr0jmtW21
rUqJnA201aAWAByz6hV5j5G3P0cwOrLNqgtwoboUytpvsTOojdPhnCZHPE1z
I9vCDU11pBNS1HgklditpOfAhyD+ukLWogDe+WzxGly9Wa6mU8P09g2FGpdp
nW8jeY8cZy7YjZfkeD3LTc9H1TmiF0VUryAthZqmsdC8Wxi5QprgvquEmAD7
+q0NS5TL2B0+sYOaurn/DdNAcCfP68nAoJmtDKN1T7HMJNypzw1E3ipch5Pm
o/6P5ozKe+FgOo6O7gePvetqeawtd58mI/2VQt1qLUFesGecvlymeUqDN3ni
n0+y7hVXwh3zP1ogGbxz9Uplacku+NICsy4OQAaHgPxk9RRyZ/ZLlhmkiA3G
W80VleZHyCItwOMCCejynTZzwdtFmS9ogvV2VH3XHB6sTs95wXt3bltMQmYu
Wyow6b4O/Ot7Jwqv10Hlb2NCYbsYC81JeC1fgb0St8WEaYZuwUhhKFYRvDRy
Bh9XXmZs2lJ6MGhJ6llM0RID1yBHJQG6dlGoz1txq5OORiKWIhEKgYXaDt7W
EcI1jqk90eO9sA46Z8ejmGEsE61KwEV7DXX83kdo6BxfDFrTUccy6S3203tS
AdSoYJ+vZ1Twm84XJRQj3ubsEJhAddX8/GyVUz6zGmkk7ljohM40Z9eg150U
kggtCauSk1UxABT4aPFWkWUM0PNIefSn5ymGDse3xfJeh8itSYWvb5Dd06Rr
UHXgU1aTW9RA9BZ0bKOPxpgEWbR9zn2Rq7syo3X+Z63yI22jcQ/sH661a8lY
T/G4lOJSUjC9e+36w8hVVK859jyT3aHTt5VowIjZXZDWoweiK5jR1irZSPP3
XjvuV4+RA4KU6Kaa5g9qNatnrm9rb+XKlfQOVPCj9J7KxE+IrRQUQQFuJbZ6
hAP6tn70SSWKyNLnqp0ACppAjpgAvoYxRtH3dHyDaDLJbhBt9w8yBIh2A4RW
AFYrghTbhuxbEXUhUIeEHUgpoB4/Tz7vrxiqomAPsJ1gepJkUknxcByWiD+O
E4upmjfCjp7x+rp0Ij/Kw+L+TgJJI5N46Bs6IyR4b1xGhuvGoLmwgjWmuQ+L
15lhcQDOGhpSB3U7AxXzzzVijGHq6utWG+CIlF95Gpf5DCvInULzY9yz2Qcu
HeirPNJX2f62iGq3I4vpg1zr8pyLf/HXQap+e3Em4tos9qsLh+vf/8xko62r
q0S0lqjcOFVFmLjH6sMjgH5fZEfUQo4pTLo/qNS4A1a6Se0fT+48J6kKmS3P
1xFr7eQZV+1lktyMnxbasJwTbRbjkrGgb08ijpwMybjbPHdtFzzEqbTfUOhA
n2FXeqJ5wIC5rW/AVFgUQLAvngV+pwaDv9WoqtgVsBewKaLn1JAmFQeLNele
3pkH5WmcAzF70LrfzEizx0VWzkG4YO0rHOC8CMBHw9pvEjdqfZ8Z9bSfBC72
u9+3+ddoWJhwDsPHBluj9a2KTFlnJ+oac6KTu2REkr+Gu5o7q8BIyaeWg4Ab
ZSQdVk2OsoFQ1CL3g38k9vbxa+V4uKXNmpvCAtHyUGaNDQUEF9soXgTl3p9o
/Qs6HfPCoGgNcgTuKunSR1gfGfUUrB/tBIFMRYLypzxpv+YHDXbS+eXskFQt
2e38MBpmye4+Shu+L6+g3s0RL7OP2fgGqU92gmdoMVOqkOk4loateKphTkWQ
ll4s1xYl4aQwqMPCl7qogfV9YIfrE0XW6JAghzh4RPi7PM+IUqGOHGjBSBef
i/EDGRF/x9uKREht9SJJ9GaFk96WE4dqCb0fspK/PbGkjNT5fD7Kd8J2eBpE
+CdighMw1EboQtWYmUY0DTaPrWvzQRJItT/cWmU39KhTO1FGIb9AntGLMoaq
IXsu570y3TMHUZtzULUsVU9bjd0laXAeXYVWd2NP81TinYuv/CExfqqeN9by
+JqX9FmGqv3jEEzEKwqifEkWwO8Dd+oJf9inOJWFoStZY+U9bxaINK2lr3F1
9CHMvEHcuaAACC//l0IsjklRB7ZPZ/t/C6t739vnp606fXd1FGGTbB1UZYLf
YVak9G3eSAKxExwGE2CxPs2Kjvi/g07DvPLnu4l8rxLefmupN0EO4VRLmESX
TFPjDQjaWgVjuWtfi40bWo8g4MiP35dPKl8jNkVw6FXPB60st37074Em+ksv
ulPTwnp+CoOgNmiM4d2RcLUWD18/c5EAJmyrvzblpJA4YdErBLVovsVf5mvs
/kqSLDOz09YKCrc7Y+hmOO0ggNjN9fpcrfrrhgxxMJUbN4+824CRmMu6xCrL
68Dhpqb6393/UIirKkCaX6dRnQQgGqBYYfVJNPBaA58+16atqjKj3mjYVO+V
fT5Ts9bc3umK+My7TrNOUAsIIJr3DxTidBfmAlbpk/vmfj5X2yx77++jiLPW
GKl7NQBK8RY2Qi70dHelE6fuYLwrWDtMXeqVB9ioczVifVhQOeaPpCq6Ke8T
mkeULCmADgAx7M0CGqxyc5IFCRll8kYQsgmNMvJP9GoLMBtXsJ9YOt4at/i2
lPRgw2NEP2EuhyP9zhQAKR071+KoNnmfkIgJVl+44IHo3fukFnUn+nKew4Cl
bG+aC8bwP+WKlhsOzwDdz5ONvjxsswP+XBo6Ic/nyud8k+ymVU22LchpfqbQ
L2JG+o0cQ5PTnjmM/SGzUAFyyFL5F9mcshNHVSHKhCqtGqbLsibwtDx0dEWd
ot4uKAXJVaL4NrMbH4uTMzYh/ng9MkSk2vs9+6ztiIL/p1tiuznWzhSFBLr1
gpx48Z9DfkpzPzT3PH7TZfyNIte66ZTLf+e/eU4ktTPRB3hjknBH3/xy6l/8
K2A1Jhv9IHqMNDxsfrZM4Nq4G62vMiVfwLWH16GQB92giJSXG4JU9iAOzxyZ
riLrH1VZMUJYb3ziK/dUbnwArYx6uI5gITb1IWZ2aF/aoUEE10WcE5DV3n8I
3OBauhsYx8YQEeJRBU9sUCMeg0Y2nVOXXLrJ9m7Zz1bYeU6fTVoJFJ9/OsN5
noBOwQVimqcpPLcIOYHuYTJt/gqUBFcZJasHkLoORWcFnhRI3c0a6KyLLwYV
41M6Sq3BSYBtC7hH4Vf0OeWUQGfaPa8xgwouf3MMyRMyj9gLUKDIshWN44Vj
RBMLsgljshfe+Hj/+LWkng6ZzhZpO75n9TDEVjP2DmK46eCkVnAy14tCPIRe
36QgeqNc49ZH+m3EyT837kEQemVkilDw9sYPuVumuznc2r2qRA4D6/+AOzN1
x8sZJpD0Q12amhWdoit2kG4JGj+me6m772WYiPdpra/6MM1/fVRdLZCfkSuj
k06aCEgj+xvx/Q/Mc5LSb59cG1t/k0jL3IuJm81XfmZZvHLbiHroPFM54EKL
x5dD+4kKzMOnpiZ0V7qsckxjTKpA1kOfmjSC7wOWdTuqof9TyzxGR9MiE9yo
xz6W4gUxvqRuZ1kJYZ8Nexff8Sh8kG9RIr6FvxXAGU4e5qte5s7mz5BBhAZa
FJxhm2M/WL2YoO9ofWtS3OxM0wILr/35Cldock5z3SS5/6cIdxW5/FyJpnpS
TWjiLDb5p1kHVdqwDNzCr1IbMp+W+dY8fizvieBuPLMJWFZh1pc0jZvl29Th
lVf9eQZm7tvPuHOlgJRcLXzyHDm3I/zEfAiDs2aJ7w9qf2sUZXpRaSX3heIF
vYcdNFg7Kq8Mu1+J0GPdz0U/KeL56mNwTo7XpIpCpLyk2LtZHacelkT9WU66
xVxFmudaX6ERHxbMou4k4NuITqR6wRpgNlrq35HL72Kj9d3ckC5bhQ50RvTW
z5Ved/6uNdYNvRMUe1lh5r9mabtc/GT9sIdv8eXdq6Q2iLmzluO0Bq0ZYNWl
Lan3RuEkif5Xwb/85nCLxh/l0/outN3UAbA3Nynl0lf9ZDKTN2rCux+vwi+i
5sjF0a8ubl6p7ijoZxTDVCOOWtdRxBIZ1397obNylSXlSRPtZu151Nks0w/A
yFeOTH7W0KqGDMpzZ8XqBpaWFDvvjISe1ThriW4+bxNLuL4ZWXbiQN1Yu+mT
zytImrnSsLmr515DdRi/+x3ePrNtAhRWk7UsD99YMIN+2zKoHUzPHS4WX4mq
bKVWRoKdLerSX12tgLKNDaSVzZEMmJPmmjSewZ+aoz6F5GBGKuMnzm4Y5cby
CQiz4NV6YsEAT5at0r6sfb7SwMjRDRK8Dvcc8hmdVJ53os8Z3paFM54G72ds
MjQmsewnLii9enEvdsDa/sD6qXdFkoRlVE8YvDmBaEsEA1HV4jtsWs7MkKob
f4OfUoBSqGPdqcECF6SWLl17kAwSFpFkM9wN3biTMjgJnasB3Ez0s1SD3T1l
RAjztO3MWdPDB372UttEP8CZUxl4UcxKwR7/efxu/7Jz3A0uV32OJDYK19Pv
j0lWUk78rcM4blkdlQfN8uEiu2LwEpXMD5zKCx0eBxDBukJ9rVmDmqVmOCCL
PpXJWl+oKvJdbAg9Hvj1hOrF2Cc3ZdeBP0gF+fylgLYC2XN01mDXA0oTSXHM
k0TeUQ3qe7x4EVyB9PZozfFlAjRauZDollSf4O0RJNnmiH5hGcbDv69+bqw+
J9uLDi/2IlqUL5r0lj78isTEbCk7EdnJDiviC/bJ3UK3EpJHC/irdd+SSdqi
BmruKo360gGG85+F+jqyzf2UXgFS+zL8VZ0QcG52OAjy4o6RJY4fNFX2CrtZ
qNI9UL7RJoWlQjowCpzqjTCDCK+8KtMCUq+qPjT54XZS8buDY6CFaQu0l9Nk
7c8bfZ5WChXUYblAl5Wzps1pCv4fZssjyIXr6ANM3uGFDwWSJh5tccCl3kdW
WOkGzfn1OADzhtEOObLQ4OXanqn1m132pVQ0QahaFeZq430F0uRgcoWT4ad+
0VkkKimhHrkESQUYxbhqGDd2PXgNeq2IEELjE0Fs9a9cXoGHxqyUVAXINZtb
7rUU9ZqyEwWPUDrxGU3ZR9SltvBtwRO6QlwbdH83THcqfa2cFmIl3l8plsWQ
yql2iJNW8TRdzyVmrf29Y2aZbfjewM0lZQp0EYeogUYjDzRPzX+YvXavPtfQ
BNRTXi7ELsTSoMC62cXRJX5XBmnrZ0dgpoHrZA4hAyEPsch19ZTOkA9Syh0K
syq5FQraqptvUcdzxRA8ACcmWQBmPOnbKns59cFh6ENFwznGl5pZDznJNLh3
oQLa5Z9DW2c5OKrP+x2QvNpJP2TJZeDktpy3XtSCj1bwz5PKSKOzW1nUE2lQ
lQ3m4NdgKYDm+TOAHguZuKnJTgNah4tkq5Tzpy4bypLe5oqIwp81WP0L3P32
AVnQJOkmHgGVexIKkdhCHD58hRGxmFOTJ/cKr5OgAjWvrLYaQR+I17n1hKVL
KLLz1b+Wx7BtdZo7FfN1bf1iyyMw4DFBIRRvksomZwebKs6yBSX55O5eg2Ux
+8koMCXHOLtZgSychEVb7/yqRJqwR6Ey9fkuAcHy3kWJXvTTUn1mLQHx9+Wa
Q9JtGfxQPtFokYCVUUdNaa8b29eBlqr8U6nCO0XrCdsT9jeaez2ViEYSeIRo
LSrI2XnygvFX3yHiE2VHi7FirXLJ2Ok/+dX/BBFs22sy2hJR5CXy5VnsiXQJ
JLI0lJuxUpcQGGVMdoIg94pQJqVcGY64NMOBLq5m+hgkQEgeBfMdmOC0rV6B
zU/xt4S+KAcE7u7A0N8yyJp1MU8UMIuyX6/FwD2apZKi4SAcqvw4Lm0nAlMF
SA7qFH52q5BN7scp5EXlZTtFwcQVThbQpXCn/Slk8JyIQ6Z9xwcHshZ4qlYp
YUCB1UftaJykGHI8IWpNUrQbSozoL79vREsijIXAapPSVdiIC/HQX9smsRKW
66v+kyi48xZTN/GkdB9d0NYrJWfo0QNyIBvI8cRvrEATeG3yYbjvsKYa1Z/j
HlHnKQ2BcG1kl29zK3fqeadJ7TEVqK+4m2LKKXiKBRN0CvqX5dJPfYIsYkvq
cxQ2HYC3W5siDze8baV81qCaEfulNIMi6D/oTHtOcplYBbUTeb8MR1fYKX7Q
Z/sFE5RBRoVSErMzgfz0Yon4+kXD798GXSD6IEmCPaZ1KUVAxqYTCm/QGXdY
a9tOPJ0ZsrxKsKS++sylN8TpIXdczSnHLPSRe+QjSG6qrXJXA7mq8Uzm3dYm
Csy7e6ta9fMptKz+m4zn5AxgvE9ZXPMZ5XE4K0FhZVOwVHpO8GVZtwwXnzBC
SyGhIAnxbEXPmnTf4m08DQHm9UPhpR0ew78JAKaCrJFExt17HPa22psNpRl8
3nNEO5IabQCzWf+KMtH2byNZ/HceIl+tuYiVjTaIMdDttGXidEdGZufOAvfE
QkGqADEBEdCJRZTFUPWAFSdmNn51VYNqvkUlBOqowEtb0kAg/U90l9unTf/6
JqsSawdCkv68rdFzr9h/H3HxSYsVhSxU2SP4o9sP7gdJ/Y3mufWpBkS262bS
+BHAWAMK4Wuc0vAIBdLr69j26GxD0srPdMtghSKnKES7j1RPslykm4bkQn5G
iP8vHSgcaVT7FdcNiZItkBDC/YcEVcqTAGwf0rInFFFvBltUeI/TChqhIG/G
eHanH1HhAOo7yek5iSDTigqkOXPjA8r/WmgVxdnXiSi5YpXDMBSJZJ4cCmTj
FRAhdQYCuuJYEqWD7JyW9YLDnYR8A+y41pPKo5BV8KdI+loSA+p35BNIY3Pl
yr3lZEX2J69ZwZeWcIU4TlwWG4+2CNlyH1V011oE7MpNvRqG6LbZAEVzWZWg
+TEJzS32/E2cMbo9fq8QEDKJqy8osEioKkGfnSeno7Fi5XSCA+4LcuGOubRc
XSUJhUrgPHs6EQiSNSDNKGskyf/e813t4eBDcnSiAtRg55GWUNqcRuP1Gz40
ryMDC0nvAayHS8wr5GJl1VYaPEpnua8EYA8WGSvU+bUB220nq2B0idaSlZUQ
Nrk8scnEfN5nHjuznzxw6NLv1EDunRbF0VeE/uFJiDE5uX0agHDBk/SpRxRu
CHjSVfDtOx2jK0NwQ8fAEKa6CQOMOZEo4rZN17nF/vxO/PlgR2ka+uvAVcCW
+U+zoacUjshzKmV5+kwkByhBd9vmqy/G+V0jJMTWEK3eJ884zLhNm3HXmFeO
7KPWKKB31uDTLLnJvm/3eYHIe5ReKet5udvXogwNWeCmJBa+UdhZsn+Dnc4U
GV2JTUv7N3JxRTfxuBvHB80P8XkdbkeQ5OjP3gIsl/bwZ9F5RfNIT1w+fTCG
B6qL7mDAGMo8MvFp29HDYB0SqJwJAO07zSVXmjjTogHOVc6gm4gIn9M4ZgbD
MLwIk7pGQ6aYvnV+K4QWH3r/Ns4crPItYQV6V5c3xqFwE/itXq25aYuVKN/C
f9phi9b9AiRg42OKe7u/edVKHgg9z5a283H5tSeZjaCxhCwMeBOEqcC8Lzxm
4zrOZqVRi+6gG4jXpc+Ndsvk+LfrX2GFSs5gsR20qzm5JEtZOZLP8gdNZkTH
ydHRmgVCM8B6SGE/tRqCTDcUAY+7HfgfLDY2ReFeVOG8F7fzyhfQ+fFoaplO
PUJaHJvX2dIqXZPBP6Jz3WXNnEfVq/lNMxRMM8cHJ/1H1SQt2L0k6G/ru+Eb
3uddZw/BVTHH8qhvxwb+poeL7Qkd9LjczjIlYUf6KPInYGKNS57pVadyDIaI
97ctreTxopprf7O01YYsFK8zOIjUPjPJvh1c1c3LfLBRnLUd6gI/J8L1R06T
F9Ay1l8VO+WRkFBSvOf1gVJvS9+6lvLYR/OY0wDoxhL12oITzhq/ZF3/to4b
7QlUKzJmG1XI4b37xrZLk8ynT4sWPfOyLosXed7ngsCb0arEoonqj9wK5c0Z
/sTEtq58yHgPVkPQAtHlsRXtIxcm2YqiqtXKyiT184UOtaig2X59YyKqAmST
4117XvHPdJhw423Db5Z5S7vb3IsZFCFBbPqfHaEvyfVj1nRqdDlvIfGyxGJW
yeHEUzoo2eXbBhKfDnuz0zI67tyeh9KJ+RZ+nhUjJ3gRWPU4OB2MsyZEFrEL
v+GRYP32//kvIU208K/YGwdslpT5iV6FJpTh1k0bv+qKUi4SviWRV2YsvGEj
J4TzDZglXMAMFDvvC0Ki4bhHmuovesHMhAt5DL/IIOp8yRyZE4wj+4RjymZM
APi6A4nyLd+3SiOs/5XYSprK7w8p/HEzPf0ZAdbnSW2el3KL9Z8+dgsgLIb3
h6eYeo76ZZ8mm+i1hOgt/0Ggwwgowyd5u4IIyKr7SPZCd0cbhbD/JIE+Qbea
ZiVoEsdexiPj4goTHl4NKNMxacsn/BSl1TqnsUlvCLGMALk7e31/ADb3b8Bw
ErvGvXy2m8E1cLHA/5IR8Jba/LXyrI6AIFiXWWJbmnLonOOryiGWJWHYoIDB
djRlxoa5PBn0Ad/Ib//GEfcwiPlCbwVU7ue3bow7iNQT0uRFn7/Lzc8gHQFz
4UkWNC3NLTrdKpbtRmhn4nwYYji28UHXaNxqX1e7p0erQSLpaOvClOX3vMaU
Ps0Z0lgzaAsI0i2971D3IaUi0XD032Sv+gjS/D9gwh1tyu9St6Xz9rqEgXRa
NLDCOk+D/01as5uyPnY4NO+hLa/BxA6+yzKS4tApuRRc0lzMOKCExQjOlgJS
z/buUSAMlGlRJ6J3s+YAjHcS6fdzn6ap28COv/B42r2Th1YdbJvyP6RHgRC4
EHqnViKNisy9GSU5TodfBkTfPAyP8CY5dS6uIMR5Xwvwdg3ANeaPXmbzYFTA
khQ25einfa3spQkVvy4c5kYB9vcshNTHaiGuurrPlwlrKbDimHqyDiaB5Jy5
LI73BnwmiqQ2F5hc/Yue43qnkrw8XAEkhTrOEU6tjnIwq2Inq3HwJ9urEDv8
Qd7KhduihqrydnMWb+ZC8VRZ+lviXQlZp19C3Lay+oovSTL2vK0TRATWfeAG
VauVmqgFLlSAGxxIAG13mV+agy8jZO6lsPrlE1H0BZyyvDumXImjRU1aKScf
rV6Yec99cmvQlVTMzE1p4GdHpHy3X7DOYK414M52h0TvazRUQNDUW/eactlq
/EF6hp8DyVtw8lHJUGKuNnEBDrfUi02ij/xCi6743DygtkAeNSOmxEv4yOl3
Ib8kIfx7wcfnBhScpHuqXoycejarw/LnL9qNw05jW1afMw+UmepLM/EU7JgZ
rrbx610uBED0K7nOteAjK8/Y3APaq3o4Aa7E7m1YrZGuTtHRZ9ejV8bQN3o+
dBt77ea+KQPR1+ILwDLU84fOdaUO/SgGFPAEBu6bErDofNsVRNyswbx10lF/
AJGd7wuFiKbp5a796EDeBSvda4wJwR9R+KMYodt06S5y6jocL56BiUD5uISc
HVToI2gnA32jDdk+abbpSBwlts2tl4I6T8RRXjjgBoZct4JrH/wwB4BIcNrs
g+z5Dh2GYkRXvkj81DNCGlFzAEY0hn4/gOSdmJgILS6RUp3DnMPN6EdbWAc+
G3oPZVvmUBOE68VvtDXPbpcJ8uqI31+vxW73JoQprrkPKnffwed0NBzD2SzN
MqMjg3eyyXyDg/MVFIk/+IHEzSwB5gIkdsOyp/1PkGemQ7aVFv+9sahTbNKg
Bn+L5cDQgA3W1GVkTPFQ2ByxKZ+93vmkG96vEh5COhxkkQP9KExVK8zcj+yy
8uYtJwrGVa8rFJWi9ezZB8Zd23mYEjth0eFwk3Ah9gWELh7XASCfzJGk9yTW
tRJSM+wE4SSGAtixGdx0sDFDYNjMxoW+W2hK8/CvWBwGBg8TQv4HBqSW2sWs
EPk/yD9/QeDli4WQwANiSCMqryrOfr+/rCWjHP1Rijdm0FJSUttmtqrNaLQO
dIJHWVlaxb7bCGLFm/uNXD9FspB+n/WyRsDdFCuY/fpZn9pAYtldOEaaOBkH
mwsMyagzf1kLlNDX+Ww8W/JPU3l37YDGlHiiBhX8bICfq1AK40GSUgtqQvst
ZDOwuWqPf26VGyAudWIDGEWc2VGKvtm8LDqTvcqqztJaFTCKiR2pq/ggoGbf
7n9I0wJnd8mr/bq7CxQXHtXbNexmE+K4fwc1LNzMxOnEghWITpxIHilZ6T2t
hJi/Agt/R5REZYOdMh8iQprcJQDoXf1S0iNGQTcsC2X+mYoJAXTiWI/By6OR
x5r3dwlT9FUXIf5Oc3yz17JDjgCklD/vI8UjfdgSzy+ZOaW/uR9QZ3PKcpfW
HUlxrbDbZvfR3caUphO/j7vL3fOO3LdG0tKQi9WkvT035oTx6F49zR89Prep
RTGjxdxNDdjbjeLpcG1WliaDDuTvYSorwJLyDdsW2QRCd3G5XmRtQAsKVZL+
eTBBRbU28+3ZzGJ41hE/PgWaq8S/MXJxDKoYYUSszcufNgqJxnraqf6yBDIJ
sIxPXh5H31m2bIdD5pd3i6yLDnqFR3yOOk2JfZ9vueFTUpO4oG2uoXEsla79
E5DdygayvBKJNNCNHDTatI9+f9ouLBIcmpdkoKnYv6xu50XAfecEGbsIsuS1
ciTcc+AUb5qy+e65Yg9QYGGkI4l+ggBlq0taWOPyldpNdE/YgAEgd0yaHCEd
gSy8qKPwoZjKtbZrf0RTWXwsD9JXAW2ZIkpKCHyS3wLiuqjrQB/NNjysZjft
agyhUzY7Yfz5HZkzAkV/Iw8UCyxYHtDa35kcjL4jvOonpY9q4Fnht138WoHo
P5XPuKyALa83rRv+fz4cvGjIFEGgS8EhJ2z3jtO6gXu/kPvKJu+OUwNkpccR
C1tbhl0qy00gt3ESKTlnw7uFdcsvXX7E28EXMqv3etSzdQ2a32bCsVHFt5Mn
vwuOmMl+Ly1MRfhZHbTHPdfGaLk9/c2voYAqGLatgF8w9mOw1ZdW4XKSi5oC
lsIsSGDgT8DYx79JQ/i+GnNtJnw9js3iYeXsonodDSmPH4QTMLaxAkv+pRrb
gbKH+3I+VGmTQ3wLwV2Z4sxQPNHZSuLe9uI3DFRRUtb1XmVeb80xPv8uYCAw
6+1LBJ5+17WKxWUQHs5KP3Y53UKh1tmtpk7ycefLDdgZ1iDXTrA3gIIX0ZfQ
9PGueG4bjdbF7aBQMh9/Ttyz/U5sGFRfgqXC/t4sYMLxUTLkk69ByxKwZ6vN
9rw0RdMey/qJ0zxnsMTXu5pzxOUZx5bQ4L6AyDhcrhSNGdRJ2MJkq1Guo9cy
EUmwoSgs7f5/LkpFyqYKvDWYlTn79GgL/j38k5lWSgf5DkbsErLWUa+rMEUZ
9J22ulhBZG5cAeki9CEmAa4m7T/PJo1yeimlbje3iDtv12DhoJfGc9V2DMIG
oMZpsjYNdvchN01jfkBQWf/PwNGaxohunDuNgPpeWiHje/uOnGwlJyMCyf+E
X024kSOhhMfjfwkGZGoiQKiNYvGWDugZhHDxzSGDaaCoKn1aiZLbrU6zPfDS
/RcbSubRFhHE3r1W/nOeB4Muy9M9m/clutX0AVOvAZ+19c3sR8DdzArGb3to
99O7mumJtx12D1MreFB9IyyBbCMDlfb8ag6+SQhxA7d0cjAf1SoMXP5+BQQI
+XRFrWTg2O9VmKio+LnWbO6vxLFBttdTRou+Km/ltRZsjQFIUgq0Zh80dsTY
V4/1UqfGbdZd92h4SrWguqSCaA3USl3lvfeQoIpXczK8n3dcEQApTn6QcLc+
NikL9HSvaS9i6/NNzNYbiwdbtFdc8DIozGXMo8UnsU8oH0/u2vrl8Uq2y8GK
Vd7kyclyZe8zdZCpYqGrp1kOEo1KHo/z9LimpqFm22X2KaDHE23TZil4Przp
aFaYrySWIZEVwr2tbZl7BwuiIK1nRmGVGCM0lpCBK6PEnf94aOlb5yc+Gilt
3JqALB0jT7Y8ZwL2PqHzh/6w8BZcnWk6YP1unckDIvMh1UPzLNyur8NBK95p
Rrcz3Tze0OnrVTxNwEaFXW9Vlot2c9Vk3auzZoW6Rr0T+QdSClVqQta0HlwQ
aJJdKj8Rete1pY5joPzzX1wk8OwFT3U7t09n0MHChmeEN9ix/pi6zDQCGOyw
U6GQXkfxWhpkZMzp1yFjji01XdPunkgorRAToFyOucNcwZhOAU6bTJf0ZQzu
19IidsXEC8yg/wxiQsw9mvBz96IiFBWv0q6X3tbtzxfoJf2uSrVxBZ4IMEtc
90Pzqt7VOuvUdGiUADWc8iUGDDIsPnZXU6T6QDBbMKuUIJgu937wWsUIGTAI
eCbhpzlnSULsXtv8poB0jgpt4rrFPGeUfvSCqujTPIvhARv6ycYp2gJy/Via
e6o/hxEaWNT3OFQ7xTq7QK6k3QG42EQUGX9n2/pzJWm2DFmm1oLiVDEYyjrv
pofBaM/FViX885lRBilvpFR1tsVWSWI9B3mUfbpzSmEgXB7oarZoCDzqNju3
yYiV0P3VheAPe62j0smde4z7y8ULoAFi/NxdNwLsRomvBLX3hodvLSbqDwXX
fs0hDNNaGIt7tDmB7z64ZYXvTWtqaDfIypCU6MTyFGsFd6dBsRFG504v7eBP
f/qBkwHg35TtXPJAIFbxa+Zyzgn6U44yBQyL5qvhXybRaXtcn4EhvkZzZdAz
b9nqpPqGv63CMhh+MEfBWydt7Vl7y41QSYXSMtXKkZDy+A8dnWMpMN/WSr/V
zpo4nj5K9emfQqnIBTbmPI/5g1pE1Swih3fwiypGt7bEig9ADpcaX7dZnrUt
jZRjYpFRzQHM2QIesMFxp99SnxsyWxSRbbtkrqV2ty6Hi6kKMGFhOISBn0X4
MyCfhqHNwh7eFojZVvQ5KY2W+u2YuNerr3cjmFDVeNfiw8N5VQmo+a24agbF
6wvOdTuBSN5xV8U0PWtcAQREL2jpEqH6uPLS1SamI5rtstOpjGnbkhsblgyn
nvUDv5OV76YACTVm1XRDqolG2RjA/fKjmZaGbXFTPuWlaixdhAcN983NJGQ/
c4UkgcpuMZYauBrbopFuQz/YAus/M8ktRp0lOmD9OZzky5R9IZ3Flre7T2Oi
6y0ayZ48i53F4Kd3s8p9qzYysIokgudfVgpPvG+keL5JWZYto73xQMeSjzP2
K0jdQF3XTj8AwJL+aySNnR2VaOzTDDGR5F2Tp2atMgBnsOygGe2rS8l+dYhg
tbAQ60FkqgZtJlhRJWFwKkIoEoGINuIEMFqFUv6k5sUo9LAGH7CRCT3+tnku
dnaq/RXfQ4ZDmhBI8fb5IfLcDuRP06ukYEhp5pCxfbaN17K5tjZWcthwx393
JLeqQA/oRSSeltZVhezyR/+0Yk2BfRzDazfn/Rml5nzIr/7CVGTUwY4fHEZa
AbcbyZE9tm2+/MjH0fDuPQjlpaK6TD5BxQwQPK6oZTdXd+zqvWZWeTYWHN3+
gowXTBTeanq7zyLLW+G+sMJGVV70CZCSfLaCP6aujqFKitAHhuh5kB8gcVfT
SpctPiaQd851WjuQuESUp04RfA1su+njWmtiEdTFxcgdAldO5ahWe2s1Kp29
lj/eVEUuG/kJluK24wWspO3KwY+ApFcYcTdLUqdDyWG5rMvcJURdxgbWYFE1
oq0oLpekgt2hXHFzSju8w5Txs+jByNGq99A3d4FaJhHDxJM9zjpNDqHlLeoe
X9M4T7qKnJWYOQk63s2chzadZy3oe1smiMPVw1ApSr9KeQOpqekv+0GQ684w
WVNr5Zl9rfGZZoFRwxDSJdsXF7XzqkAs0sYYas0FvGUuQPeE0V3IlvMSvg/s
kiv2M8iCnZ+HJJMy83hsD3wRFOdDF3a4wi2grEOYwbIqF8zpEn7+bE/WjLXQ
Rgx4fIgckcifwXKeBqnDVeKC2eJEp3+GO01bESDXAvpsWk2QeB0cL20z/q9b
t6qr04qLf1gUvlm9zYiCUXCItjzTW1mDIyDKuMlVN3jKWPVAm2ymqLgCKe1Z
4GyIAz/pFELxzox7PfgNKhPAsAf9CIZiHLgHcaikTJL8/lo51FmNY2P1lRXW
Fi4AL7UkaWiVzOOLNVsbNF2X9i9k75KtoEH1KL97O/d1vEZdeTmcaMXd6IKP
S/+B77PXe4/tjFMIZUCySqGEQtua+9nsKR8SCgseoFGi1Hbjcjj/0Cf52Tzo
bXZ1M1MM9vHnel212/ojO0d+7ZstqnOzI8XParDj2rJLQLIkXTMz/8SYvPBB
JX6RcYT2zqBa4oLHqC1Q5DX48wa6RAeV0hll6fau+cdqmPRaMtUFLmwtS6sm
Oin4Piqm8388JcxWUHurOsCzzkH9AIE1iVSKbzK8sey4AA5UU4eSb7/Erd4g
dioBm1lsiXz22cOq9S6Lnxpv9FObtml+k3DbAkIugauEO8Mf8XlRG2TxMUG9
WDKRXt0a9CNCCDHTnOwg/VuJCDePpRB3yLxdyPtfZrthi7XOWDwm0lMwkw0x
+1sTD61nF/YSxnEv600bUl452QWtD97UI/nZF9GVOoUpSOQqDBYiFaUGzd8Q
Z7wZbsRzMj/Dn6N+S1RTvZRX8BmFSO3fIP3LPn4uvpDAl8+5e8RzUFJoYU1O
m9SDY7liVPIPk4Efo/aZjCI49RY/Y7n31NdCMiEhY4+Qw3gIdPEQIL/9vTUc
cJCq6G9WmiJJ5HqG/Si4YB8U1POCf2TpKSMCjv2Flp/ZVyE3+hjGPUeJLX9Y
xGBjKflQPXI3XUYWZ7ydaH9SxM1dlSdgu5sjQ75fqNuONmSmdz7QcLH/MBQM
NZ7hiAdFtDtArKB6Ia6F/lAy1XDYN2/Zcc0/XBFjZHhkzbAndUlsKw2+q1tj
sDLiZ1mqcHqirUK/iKlZwrdylYc84I4gxCmbiPdqH+SjN9hveN6Wd8SwhQQX
d16VdSWsQq8tHXRfm/UPQIo1K/WG+YVdZdAKn/0PcLTutRFxNqmRO3M1gJ9d
cpyKjacdIfheNcRqyywAT0QEoXBIC1v9UnnSCa42ytgOLndafqbNf9CLeKLg
Dlrr6Ihgq+tboQXoJRrrV0K4LFvUG14DS2hhwxhJNqg5qxbL6CccmJMtZhde
qTcHOyqej57Sv2IapIED0OTIHws8vCMbO8WbhOoQcKt0ymUb+RdtAGMuYtzD
c+rw/Am8gHk/ugpFMidE7o/RqB56mAjvgaD2LK5TODFa9Tf9ZymWPfm/gqr1
qN6NOregzgquWofKH3XiQRmraYOtniQ/z+Nsw0QVgi3C4S00bXc9ntSyhlkd
8VKHgHHC9RqpqGUnROhVI6XM0R0+vn5Qq7zDSIyyk/0dskX7RMzUd4AODCX5
LaoslfQxxOsZNBg2Uf+iArbOuFUoINZOuBmdaQEoGWO7BeWh1sLbQQYJPgLv
u3roXgf7ULg5qR1lfCmnav9YSMbIbYLkuiXCHLxuGmXCc2MI+0qFPBBDbF00
9e1QCaA8FpveJ13LwzWZOeNjJ+H8sO4pFflUFD7uJFDaxShi7eY5UzM2u1GB
/Cg5UzOy19q5NM04URO5coFegc03LVEMHt5hmUXMQ8O0Ae9YSDZue3ytjfWs
/IjHdqDfoRvPI4F2l+mavWJj2ITqG3DfUZoiQhbsd2+rmmG4Ts9b5RExdtbK
2Ok3WfayHS/emLdhltp7+rNstE1gvo3siwUSLFiGWEHEgMtKTHDljb+/bh6D
kPBb7ZxL7I7udaOGVbZO8eyi5+Ejxk51SJbomjOR48zrxKd7Zjlc1TKUw8Ik
JqEnQGNQNBBMsa6FLXGXqg1paFpgk4QXQLIfoN9CaAVsdjl2qrykcyR3q4EM
Iqb+RWKTRjEhiG7wT+QZ2XKRhbrn6UltItviDHLi2CNoMRO0bJxNJ8xBTJxb
rgNxO/XO+V7eg7ZP26AyYCsuLUKyV/Yw4llWXHHpXhLSsv6u/VZQj3YC5mm/
ceD/jfHXSix5oc2Dc66q2WBfRPTALtULsHhRK4uzCoVEzgC89a02ILEFFCZd
YbzlREJUXTVCLpJFKtwAk+qskXA3PRE/Y6/vE5l5X/SPYH90M67QiJ9V2QWy
KF27XDrKyz6ickvGrpt9zaZth6uvb+WrUVziLVBzxqKJiL77A8oG3RBeac3W
Bl/b5bZFeplbAOz7p+nLENao0ubNV8j3GxkIGblqvyuwTWFaMlM2PgOC8CTZ
f/BDl3OUKoGJDIhZQO86Cvkhi3ovOEb9CJUsvkUXKMEGtGt/f8jD60VQJ58x
qfmuAJxLTR/Nngt/eusDXaHpyWA7SI8A1zZAvuxinAkI4N7n8RuSe6vRR6v3
4JDGE996bRsFA10vVbq79QMKmMm3h2If/Y+VvDlbhqNeVZxVx6dV8XIAywM9
5s6xJxZKEFtyNCW8p5tn7yYwK12pWLnKv+IdCz7yv/xQpLzUdPngn6W7NlrH
VhKiM8WqzYgn/kHXB6RFjJTfMMq86MHrVevF03MJHqZ0NuBrtMhOhZFUO5Dj
zx/voQ209fhqtwdLYPQyzqveQ8WICH32nRGy/8oOENUbY922YnvPTBJoq15h
GbzvfXauc/Spmdca4xAEhMFruef2FknSF8HbwiDuRgPN1y1DPH1HpqoanKkl
+LBWJJHq+iMhYbz9KgIr63uXnplcY69F3akB519Ng9zC/xqsh//YM5LJOX73
02lMupHxLSBSKifh30/YUoQct/p2pvDKP3hnMGOPi07ub3V6/X261lFMf+BH
Dg1XkwVa/0ObS4jZxIJ6jX4FSTvAc5OCWvQyWQanDggqBHrqtUluI5YFSVri
8Uz5ECTnf3uIWLq5by9V06nQeYoWSKOGAw79a6i6vUXIwWBWUFtCALOjKKN1
DXzJzqS0BWOa/QiKLvS33XuhuBAWH7J0KVP8WRW1MNlD8FTLxZQTyn3IOHCo
zuMcIEuhbWMO7JKOkg5RZLFqyg2iQ/KvH+OS499VPkZu1pUGXcxIH+5RT1qj
RI8L48DOL5c6iIKqZodAT4QRJ/AjJvNVmlgA+KW14fraOrvfAdofmQeNLXVn
k3S0yf4taVpl9t99EvKjfEwMFxiVsfhT46oqK7rUq7/o/bK+LjRMQ2Z2uEtY
k2+7K3OQ8lXBs2EsLFMZug5+bBGAaj7MjWTkR6jJuYykOICbBZ7FGSupdaK2
tuDwyc92hmVjhiRYiO3UBI+XKdsUslTkZHLPt6vAvQzWo3W9YW/5a8L/4LpP
N40ZjpOnYhs7vMx6A7OduBLd1Bt9iaWJlPKRhAFy3na1/jfrgFG+VnGbDgDQ
6PBlQD0CymQzTQZrv4ZhGyE3flsSkToIcF9rCsYZscPAYDTm24t95u9BsQZc
74TexKwrrNzF+TpPTOCaGlBp8EHYgm7xYkIs96FizGVQz799Vl6KsDjyOqde
4RHKlPa+o7eQge1Jxi99L7B9hMgyBiioNnDcO9qYGblup4mEqK7Vjf1Rw07i
yk5TWz56zSdZ5YI081xiB1LCxM0n2LEkCmuBLiqDWCFT/NxZr35qm33qEYxU
7/63N6vyO9v8APD6vTso2fc0NBBITcVwzW4ZHjI2wqIlY+hMN4ovnGrlHuGU
6VyhGYkTfyHg4jAQC2RMQ/lYxWu8XQk9hFNnEmNoTHF2ApVogl3ZJDE27LYC
JF/uBHvZJfQhuRutwb4bBgqdzrAPGDrqRXnWt4yrOuZJleTdj+YFVHeo5uvt
lNTy48xmC1+VeUdv4ZBoUq+3h/p9/iQoI9Djrk10t37SkFiK/vJn3nCr/sy6
L6QGXZMejn9mFhzqoylCzgxW9kxUYq6gny/SDV//HgYNGs4AFILW3W4PzHgo
XTGE4HIED1iWh2Q/zsKWvOwAYz5w5m+OoRb7XvhtVtgxohk5fa3X557ENozP
gwmNzY8aNmY0Ek+ulH1izMgOcLxQ+LtrhCZBwt/DBompvhgPrSA+8XSZ7Uap
cRECD1DhIPjCi/gUmivvXZIKC5r7JCkBKFikyzHECtRm3j0bJpwkV1x8c2Ih
8AmwB0vjoBW+uD8UENNMtr/ObDpUBHfbEQl8Y+sLJSSPpLTfbNfX0QBdTe/M
Iwx4s16G7i2zmMu6F2hfGTVAAjawU44HznrrKSqpKMMap6lnPdJ4P0CZBMiS
Vpt1k3prQpGiled5c2sZbvdjcOx+BcjVnIbl6ObBr8ZfoxgB4sUUaaPgAXp5
lGQRR5emKrMmR9Ojy7BX044+KYHBontYqviet8P9DNAIHVPRlZZxhW49nLl9
SzXIzWJx2fTYjAOEaxZEGDptxLaqJjETLPvW9zwYvcLbBiJnBWARFnGC21xL
v69OWR/eo2k3kcdMkB/ds3cihxebFJ1EZGSi2pQQa3htY98yGsL235GOVIRi
rfHSLjGF/dSfpWn7V+3/QRn3Wyx+rJTP4mA/8vSHLcgpFf8yRelDOBnJFV2+
uDon+LO7Y2RuOVx2ugTRfndx94ehP8Yx20jkAMuV979fx1mJ6XYBF4O4U9XT
N0xibaqp2GjKlCwTQaqIFOE6h5f+++hOPD2spr6HOvs4nKHbBeBHUJiRz+FG
NkbVK3Xe68Z9MGZAuFdGnJDU3EuE593UWsFShFlUI3snRFx/OGFeStyb1xvm
89xr+XituhkBDeVRV/JVgWtoXzrhFe6OvSbnNycfclxJmon93J30tjnM3+ad
x0lO+DhJOQNpNELL08x9gmm0pgVw5jztnz+J5pZDaEpvPtdcMqsVg5PySoy5
fNpVl6jcxjxEDtk1pHxTYXjDwR7JA4jlfrdEUC39OlNsJ660cRSd5WWas0Sm
eEzT9FFl1YSnGgWi2gttRdykwmJCoc3aXF2ya4JV3A0Yx9In3AGfcK7lLz7J
/Leah3+hPur2CoSap47Yjn57LOlG25fr2QLlmIXRKI27OfCv8ySQMGwm+3g5
H+NfbPZiXwLCxXwrFi2hAGoPB3brnuD/vQbt2dOQxiMj2rR0OxPTSszg/lcZ
aliwNQGHV/YKSqsEfuPUVTDqnhx3GlDzYZaqV0G2CJ08mSYPK2kT0veMPSdX
d3aYJa0D5VqKPdRERobhWT88XpJTuppZVYdx20Zy9dHgT1NWhZKFOvaOVeK6
IKw8l4rqqmpLEpoazrwfnqUpwoYI5i/3A8bIAZLNyPQcinqSBBpLLAdMggBi
5Dwc9RI53GdX6GbZfAWeMhYcawt25NGFLFRQk7uiU/LTRwp85fxofvso08L5
rh3o5j9RivCpf/ffcJfB/U+D22zX3LmH+0NHpvJO/aodvMcJjkTkKER6ncfr
CjN4RE/hENHKonXgS7rJd2tve1uOLT6kOlMpfCNM7TuwbyXSl9NYQdgOXBEQ
amLnSTOqGGp5lIs6BrT3dUpthW/y12OmpBf0FJ9dwPrAPIFRQhMbedzijC79
jkh+/bKoR5NN3Qc9OOmjI1ed4sANHfa2MYm2sJEQ7RrCudrH60xjdOzthlR+
fUUzhN/P1AmOVS3fYvp6em99zSzk226SCGHdengIPOqqHORm1uYU4qoZSv67
qFbRXzYconabKAEY8yrfhgEZQL2mAq08XHPUFeP3rtEnQGmi55nrQeiJZBNJ
hZ1vH9bnBh3BtY4GtD/zMSRY0Nl5ItGx+IQIZgjqwCEOHkMWPPkX40J/fvJB
9kzV5+2IpvgbWt3CGelTVJNbcVw2vbWxryQ4LaJUrQn6IFd2mrOP1bdUqgHx
uXoVpAEqKI7PKtBVhWH7AZsVmtUEkkUXT2oaWoAV5hOfn+YRwe4+ufpyABAu
AeZdHMI4xTkaSBatmwOsWJ09zrC/nzBgGxZXWV36K3hkRglqNx0ZQHs68q3J
hM+8v0ZI9zaARF+UqGC6/JlD+Kf8uozymCMwoSeL7LkO6PHTHXZtRuETgwXX
bDgMSGsJoLX0Zc8sElRhZMlz4nBgAzcLOOLzEPnauQNGZ+SsBB684x/SgiV4
HCxciCtzI23ZwEFOyb3wjUhGm2uhQk0d+so4kd2ncOBLnTpyUUngAL/BLIZl
H6EWG/7bEKQ9CAkHI7VopcVhFb2iTHDahjucQ3NcMA26IMTvBAGsebCTExvz
5ZZ6Zf7uv9IGHMJt5+LdzY5tFXRj7rZAOmjLR6mvG5bTe8551U/WZBfHvKRM
GXbTm6pMRWG/PJRliC7DLEHn1Xzf/pXA1Mv6AcmM3F7u5xF5MTHjfVRtBeKg
obeT0MGKWMI8UhrqNH4/WDReaZZAbqS44ubmsUL6NO95k0YVWs2JI/Qj3/5/
Zm18YW5ckQL0L8g/wutdYV4KNBS22/p1KjToDUjYzNNk9hZoARvVWyJZ4oO/
lnSgwf4SOSPKBXnBP4jVCohLSOJRPpXEsy79qL6A/3mV8TxBhBlTO3+l7btQ
KSshRTd/Mh4kuI6uL4UpE6CJv4Qqse2RSmAdIk55Nv59hOevMv0/cbgzslDT
KWjjGR3cIoAUt6SodyvSat8NLhEzOEYDvP9jy5fd4ONiBLtPo0uRe6Aeb1CQ
lyhQjr9igmZhYo4gw61Rbxjm+MTdBgnJL6Iy2u6YPTX0yeBu5/pDExD0izzM
RfLHfKOjID8BMPr0kE1hOUUzn4fufQ61Wugr8xVU439sZ9gRaVd7cZ4f0YbY
FybGhpnEOhH8txTIItCyvkFpdz4v6R73UcSZEntrT31UsvD/g3h2jNHC2Suz
kRuLhto938XlOSQ2sOcyAe7GnJuPVzEaQ4vGuFGJCO5Cs8J3b60pE6J0GIhw
NFLByWg2AUzxlXBj+YPhzs75BELQIetkGfBy7NLOC7DgZyOkJ1sUGoief3Ro
hke/JigeW6SJ3ZVgUj1dnNVvjP/YuTX/1BWShrU6psGoxqsT5D4K5TPK8/zo
2Dy4VLhc/Qc4ehE5KDktNbV5iG3MOdcszucKk4hnxDtZwrv7mTz8ljzdIrWy
rT8NRo1L2O9AWgVvACNkWQ+D28Zs96H1lOTQit3M5P+2xGjINJ1hNL0ABzKK
gAr8Ota5brPwE0sh4dpBH5/a0CSzLmFtmF3AjL/w+zoPpoZJuJahR06CbraX
sp0BYlBfoqAJZhLh/bWU6PwVbyz2Hv6OmW4qHAgtSFSGV7nIAQqte2GvnmI6
5TyExgsu+6qmnTmRXX+EDFy4brMM25h6NfAlUzHazypedCzsDcBMrD9bupY8
whkUq7KGcMq9wu5SnoSev60DhKkODVVhrSHwpY6+Kuc7rr0GjsYDuffD9DQm
h1hFtYxriMbf0vCYxpsJKP9X/fO4LPh7RINS9C76lSKvj9a/74L3CrlHa4eD
WyOEGh9qikpqDh77AT4WBIABaoHALraXrVyzEjqo4iwmTPQI27XyC+0oBpFy
/gV10DaLLJBduTGKj1C40y+KVQDjTm4D26y47cGSY7pZeD1E3VnQBIVd9/7C
GqtDW3eVpiW5gQKTl72bYo3HfLDLbxEPsevMoqSZcy1U3Td4Swr8uysJhSj+
G3ZXOZO3OaMHGjHwpcbVX4Ie/+l0oVmGQJIzhvYjqJFevTuC191feCJ6p0Kb
Ifl3NbsRYkYIaGDkyUNCb+PlHvrairSj4uXVQgLsC0YiYVgQgwrblKi/XU1q
GaUJVmZhU49gLMYOwe+XE2cyTS3AFbFd9E6gnHI1lXM5Oxky8Aue2Elpyl1a
lWZPfYlXKk0qDeE9CjZNtR7tCF4LFr+WXQ01mGN3cutloPBTDUjB646IUPt9
Zntbo9ex1gHU4LHhu2HDd/tK41ZZCjmiwMji62zQKjB0k8HuOZVVNarHn9gU
nmmxzsyrCr96C6wihjasRzl5b4UiIWlNoz63YPgWlTZw0Nlz/LbOmbow4eJY
aV7F3PdThChgHZqp3eKtQ77B6c8Ab5Z3O5Xegv1NX7Nuxq30eWPAmf9HTF7c
wPOfP9JYXD02auNPqKH/96Sh5ERBbPzeb1GfzR1dYou5gACtQ1VcYoAFqHpt
zA8kIEct2JKR8mohVNaKGJeobB/Eli4BznSsq+qvXFJGXy9g+tBl8rDnFWtN
kskdEBBIE8ERS+KSPWu626dpRD5VnL59nRcx64RVLx15ZAjZMhtDe3HrLKo7
E8kOb4coOWqQA76R3vowRGo51fb8e5fIn9vgkI0lHyWYgzwbPImnOYkXanXx
OFQkkMe0AToa+Q5g7kXbIV5R7mXJScf0joR9K80ic1ekrrSx3l3fsz8rPkzM
dOCN48Fh5CW13wHUFQ805C6N1YhE45QakhPue1hVlWCZI2Z99831cjN+uZfX
EhcexuyKUydv8UlaGi4yKAUisGOyiTKMfyAiFAF12j0zqyJ0D5Ui3SNmoP5H
xgM9xNvOmg+KS/mBTCSB6CzbzDRFpXllq4zo2gQBrXWgOPfIM+DnAZv7GCqK
2/BvnPACqJNcTK0nIp5lJsGIOXlhd1lVBSzLwu5uFXij0buAuAivl66E+rPd
BRK2wmYw2+6too+i6+vfZjQ0EAfdCRhqBZ8YAMdWiwYgQ+bxhnQdK5Kag+k5
ybRPF2fVcvedDOC4M2C7O6zacSWF3tssjSUu3YN+GA7Uj1/U54cdobl2yssm
EIl5frBsioViHBRafeoTglpeXMRnpvURhcEB++pMLf4b18TC10TcWeJhO4my
6ZZ7mHqLjAY95clXgvvCeEzHBS44cwMrax4Aan4nr6fikwVdu9mvLl9U5W/4
uk6KU9luJmtNuvnm9nioqMZss9sT4V2AIBX0saN4yscY1kRW2F9vLxOS+59z
p5nSjNYj1FbzVVSkPYv9sDqd5d54HCDJYFlqw9tTgRnCgngGp29zeOJKUweL
0Nzr2TrUooF87lIhPVMfzeWTj6jZxxp492hYaPawbwvX+5FJ2mZKGLaGWceu
T8IMoc62SFRI6OGHklZsp+TwNnxaNDDIjiYZJVpXyTpVCGPCFreE7AVH80Ty
cBUsOjbUAuMCDXPvtVYNMpeDPhzEKoeMM/14ObirEwzl5VMCTHiXvARaYTbm
3umuoMAo/b8i+jRAjEJW3ZnKqNG5fpeJPSmzQwn/+dgY/l2JVPgiO36U/QGx
L6onR0Unlb0uWjr4/Xw6Dj5QE8GGOe+lfV0E4rk/pagBq5KBCmwNpGPIgqum
+HStZQCY9jxH3HLsYa0p5Bex/b13pmChwUpT21qUZ5zHDoRrE91ieg8ACH2F
A7OFXg7+pt7jdunNloV5z1enR5eWDDoWOIlhw5IiUVTpPfDBldgwou7V4OuO
pMVcqc0uMs0GVU3evXYkUVWAjTE+GH3rIaM+roFuGts0m4pzNWsG5BoDpTE9
Wzbgi4rIz2nSew4X4+o+La9/mFeNKyBTOY33PcHCc/XTr0cEYh91h89QPOp/
kRgG5L94GSihfpp7r1JF5BGOP4DlXJm3JjVhFnROoOsw+GlVA4FMqstH3UEH
5ITXV/H6pfLc4C4a3Q5ksEJEplEOXgENe6MKKv/pVofzmrEXTu3rwGBHidbZ
EMmFmXhuym1+rE7ATjMpRHsWekNrcjaR4wTpHcLrcVYu4eJ6Sw1yL9ZG4D/g
Ak82ERUhU0258LPJ1ImBUr9KhsiykUr3+Zet9rbOD8BqlE4Rbi7Ej/iahYU+
gM/BkWPLcL+pSteBnqwLRUzJXfHAvaOECMAJyFV51V0+WVqrgzEvZlKqV8NU
AT8I3Ci96i1VdXnHKUGpkeSoamKSI88TNvw9WtJbcJY5D/u5xijPHH8NgK45
I+pwFM8clYjLSoHDywQs7Zw3lXADSOVluamxMCAgL3CZrmvLQxdQMgtxhHRd
CV8qnF9EuUzEkMSJYdT1qD09YJ/sVYW3RcnVdkG4oKBpLLlm+R4bWJzrxymU
YYHZO8ThNXS6410s5KKKHiCJ7Z4hX0HaIT1eEeqQX3Sam2qLwDfDW3moJtk+
RTAuvl0XWw1s9duuUqn0NbGdfN3y2wUYR057/8HtaqaIUzm+tUuxCK1yKnB0
o71ZHOmstB3VWKUiw5BA/xjUjH57486/a4rlH/U68bcWYZZhhxitatYJ+T0E
wBrZBQgtU3YLjv2NmI87u/fDZeAPLbBvfnK+WB0qtjyN8afkpb7fb29rAmmr
IzYF9zGlmtaSAek9uTv3acKRyhf8HabQPY3oqtd139xNhsQ7gYjmJWO7cZCd
kOgKJ73ljVYPZjVS7R8uTn/GLoXSF4EyRFwyW7bQpS8Mt4Hr/3OLP8LUMRm/
wPG9276NQ9407vV8yEqpp9DiJfRtlashMvFi7CNNj9GB6jQVlpAE3SQchhFK
llUBcsONIdK6AbKcRU1jyUgSvNZ5T+4MUH6OupQ1HEwsryYq/A3z5nNvyiXD
bBmHNqh++y38YYbJm63XkonuF9qyIBsUc+Ao6jkxrMkjlUyoIxBHjnf/Wj/Y
DSfX4wHBvXgGVkesMJczzmX6VMeVIaWfIxLBwXy0gVVE/GHMp+XI8CD4RZnV
PYgklIEToKeLuPgj5bZN0swQn1TVT4qNeEc6Ej4oebCVzXNz4HMUbnPxNV83
PVhamRPDHqzUq0IwPIk7IVHeEPqzRgOgSBicoLXSL9L4Hg4DiLlq3mRMmSKO
ZwLAW9kz6BlvN6SJC05GN1mgb1e3q12VLjBZ6U5n8Esr8//GWgyG3tS+RBPr
OCyw4rymNlipFV2UlBwWD1vya4E/G+08e8YTDdKObZqAw7qJd6/ZIUgwL920
vgToOcdvD3jlZn8MKP8VocJ3cd2zdtkL8c5B6/8IQGUlLeJ+3ROjFaPumtVP
CXRd6LbkAk48H2L5174kl2yI7rykRBNtf6f3klJwBfsVne678oorSMvtY7+a
jw+Xh2+KPYf9FCAtcri5orTdazV0yG2+9clMh86OUsvnsbxnl/CgoEEzTuD5
UlAZjnj5sxW6YgxA7UjDfVl3taKR5xKPZ+kKrg1DxXpWnkzmZ3S/K6FJflR8
TMh5KZz6JabMBmjVFt76z/H0IlGKm27x341xXnx9duH+kd5+gXRY/u8hFHCr
uAaghckPn/9SA9W5NYLSP/W7f57amI9S4qfTeWJN45udj2fwE3DQYxxdvqtP
5wuaZyiV6e/vb/SmRJ+X0OC8EhPzKXTk3o1ap1SXHMdfmZAhGw8sZnT+/2l9
NRP+JLWu8SOQZuFymAV0YGSxNZmoQtZ3aO1+HYWhbd2BFjI7eQ/GaAa8y7Rh
HZcixD/U8yzlrKKxysj92DeThjn8Au/cgbhcsZLQR2UzcAJgSuwOmQhc6+m2
p2IxXOEwQz0PsFebgRKR1xtEK/60EVN0n6639w2eDDsLJdYfyVeamTpM9Io+
0OgTVSy66ToqHUk9lTn2ZNblnPBvZZrbYYZl4Xy+E4UYaktOmjpusy0317n+
kDy262hUHeqv0ojx5Rrb1Byn1ODwFzT58jGtmQ3N/oTns2GeKbzFdxhdijRD
LgUjLow+s+AePUA1JOADzcIfHzO6rdFzL16eI3vfjzpUIaU/zPMBA4v8ZVBd
TCTZPX8VGxkB2pH6QjfHJbNzkrquy7T9gjqExuM0p4axJCNISjhi0r5wPYQI
gqqYQBBjDAvamaW+QHzcEVR0UV8zMozGEyKteod4O534+TL4jJ008w8aIBb7
VtgBJVUnvfVVLfxr4pvH5z2degZ1oKF5OghmS/riSLY5Zv7mO65EH6oe/cCj
zJlVpT4fNUpl1j5WvS8EfUPsy+dByIXPBvEzwD4o3EaE4bTinZh/r1mYNr+1
mazoadJGX52ewdrVE19GvuKt31htffgRIb2tdSzM7j7DJ0niN0adoJFMrgUD
4Tj8Zxvy6af+wvoctk30W2ubEbBglCOgE7fJl5x+7r+7+pehrbJQFcfff9VM
s0gjTvitSO2iFRU4dgDlXESxq5WpiPS1TtXISgHbbpC7f2fMZSxEp+WLgFbO
/1KjeRx1UdLqrARCcqhTHrUVVCtmcTOEAWk5zPOW/NgyHlcrfOY6HDgMcSi0
hlvYphdFGrQkyVlTWe+qHS7IQW4zwC+p8nY+c2qw0VHacq6un/zOJBsssErM
QjUk/dg/YaAm08mT7g7yIJIUE7BjZ7XrP65C4hTqHJg9/ZGGTSu0mXQp8Sn9
1CPSh/e1uo/DbvKn19bGEf7jry49XEfD9PUsz+Y8O6J90pRQ8aVoDEYYzIDL
33ZyRT/4THToznvlSfndlTRko0ubd8oIJGerommyhqVmCHxRLgiCpD9JuakF
6757TVF9rUb3Lt/v+G6kR0KQA4reTYeyKAJHZHsTyib9C028f4An/26Bb12f
pKojio9YPnluv1eFIHjNOspNUPgFPcb57xnan4cTYvFNJIoegzmod1I1JTsA
fSTboErjAy+DRbePz+uIURX8gXLIc6sfkHDQUGyM72ttgvgiNWogaqHIe8oz
JT+F1z0AwIVtTot98ghUVw/MtjJKiob/dB1kM175q1fvbNAA3r9KMAQqVdQe
dIf3EWUmGPW+xa78m1BBGacThQta05Af52V7241Ylt1jGzNqGzBJdqDLJBWU
iLryGrpof4WEBzLRApLU3WzglPK212GE8Cugo0zfIfcH4vG3JyMuDGQAxv9S
xBJ/i8ksBBmHWEAD/CDpNz7rPO9mIvQR53twzxQJ63pdYAyC7LDtVdqxTtWl
PfLqAJ3NWPOS/uRkzeCJzWcB1STpCMhHj/FEoH59h3O8zr9tx3WpMndwigVa
nv+ACRsnf1HluTYTMBUbJEstvXPQoT84FVYtFdWCN9dJFqdGcI1izJ2MpYoa
wV5i1rGW2GKxsP+X7EL1cRImqbcSCvKXVrjBRxLLckHklOg/f/qFxWfTy9Ct
ftaoWHDBGx7XYvNFf1/eNVGjP7QSnVzn8eHePym7PNAuDaKz+LMdOnSMpnmm
6ebHPHSDTM/ATs05I4ofGvVSLW8C2WhUWw6zJ8PQVGEnGMKsW4YUv/+ZZ4jz
KFpwjtjrZbXp5hvZrMga6XdUpiKlF9DRu21UessdPlD8ELCxPsF3+Vh7RHdH
hPbgj9e9ffD5jJxMhwN7tDPagGXnLf4woeySDuV/A3oS25AWAwxwzdCS4tBF
xcCrW3+g2sYdY0G1l+8sdIY0W7+cTdVxY4AIYqk3llkLid1CUxpFz+nKT0sy
pQOm6c3zu6Kep9ArU0EANr0cu2G5FWfBgTn55XArQ6NZHHuPH6nw2GaA0Y1t
yDICIZZhuaJopfbqbjcMvwVM5a346vOHMpnTf+H2r/Q/d6LDjmzrBwcR7vlE
80COdFuWFPmEfwXKN8Lx0QXfPpFoHadgprio8Gcyp3k2zyr+uT8oBu0IyF1H
Jjuyhi3my+mTk88cLd6Q8LBtgX1HHwFZq5wzQ4DyJM4ockdPIuXDoU9zkPSP
YnbkZCdpj9/pQX4M+qy+BxidFhCliMNYO9BI2ovsbtfZUZW3Mm5IpM/ZiAXu
WLSXnpyGQQPHzEhbjR68KrS49M+HgX29Hj/MA7KLY5oB19VTDbaHXyWp5XU3
7u8rZl1ZOYLHwaB8mJ8484kcE9RVh/JLUeb8h30hdNf2N1u/Tf3seg5jHtTc
075Tg0lR0Fe/WpWe8OyJAhjHyIQCywerA6DppoNKeJOdxk+8ccx7yx0HxA0J
cr3NanU1fItZ2E8HkyjRwoWtZVsuCEIfrCpYELI+pd5UiZ2GHw2gV2D0vZQM
Gd3jJ67/aJIvQ6VVLYi4KX6QyXOSvwXCxS/oJM7hSBIe4nRAYfMSskcEaf+4
SZOicAG1aQELoICAzt20e64W3cqkU6IiDUhaT2339MhLu6ci1jV+HLvOqmUQ
T79Nm/ZcTUNwbLnotjoz9pPBVUAyUtg5Eosm9xDsw8Vhfvp/pHgmehnYC0Zq
INii7o3f3DgvwqomuPFkFAV47DzkEDh0gef50logno/Kn8B85I1GCz6DfVhA
qHqk4ADkx9Z/VL+9q1ygs6vkxqs5GrnuJQZQmHxpsIchhyFFSr+Zce1GPlB/
1meqcGpbxDMVCGEgB1yLg04tQXZgukMIIKZySZ03lexBXY2RhjbOFBtBy/MF
QOjLu8iDzvUwfza2oakCkGIuA3Gv0Q/xNhF6GGUEnfZJ1EVyodbfswexuIcA
qlFKb8WgbqfTN/Tjj3ElbhwyrekRKNGeTwNHVcCXegQoxKeP57oYWHj2lCi/
zLrKKBkBbfhGzWVTJQMFLUWIQKJStnZxry77jkrLCu45NWWtch6HQz+NcWI5
Df5AyOzrEQocNvZVkYYnVxDm0wPfHhs/UIpHCLxWX2UrPz/3A4izDZ62d8zT
wxblz26U5eSTSwWtXjjl/ySSmy74FZlFxMVQqQwJYYEjvUFAoahZqwcgYMsm
ARpjMNs/ZW2WoGy1xliBmOOPCM3slNejIZG73AyNgpdzSJk9P7fie9dN8w2u
l62ZqWOdxUcKCfS+vsgnihehfnOfk2qr4LPriiLkP1px3HqfJ75sAQbaPKMO
qAdHGDtxa2GbVPhHFKpg7SkQTr2ZaDtUWJivuve9w1aj5KX8m3kAJuEVx3XL
k5ovxro+NIPTdD5PAjLvFpBP+0GYTvHCDU4b+2zMeuIAqzwzdHnu4F19Awjj
nWC5Z31rbzHpDOPhyABBTNAcAgyqhlJXHfvJdEF5r2+0byLT1gddcBLy34h3
fvJJzKfzk9F82cdHxCitMTP7HnVqgyEqWpG1OWd0Vi9GvtU4IW4wQIsTkRX4
YYOYqKCmkxaPTUfR/kbQGQNIA5ueerba6/tZC9xuosGRRU9afgmOjvBqutC8
PrFlAW7QcU+GBq4bZWNM6B0aBqbzxFNKTc/Ybi1MFs7mdM0QMT7goKQbYdgW
qzV8y86zbtwtakaQwDFssVESQOOdj2gCn2M+xtxjIje/m2MPHZ87xIG46H+2
JaIhu/L2eIADXy/bBbAH0BF6qaeR46Ch9sxAlR0jCG5QIrXwrvF5Tpv/M6hf
wfLIUXCvzSIDkXuYg44zz4Fg+10HHPYmHyiWgIMuPnjrjAlFrEvcIr4ZHBks
AfT878WFRoEwLGns0WKIc80+1pV+zhx0j+OootYcD45NMylU/kVzF7TTPcve
pj+2kejQiIkxK4Wz8ZpY6/31W28MYxcO0wj9b/x35lRXA4i+fzHfctXLvamR
ynDhx/BVT2QVFsdNsieDcHqMs0CGy7KReLfFJO8rgzKfAg3butmsCCqtREwP
rV/Op/5wi6Qm01ElOsCrOUmXp6fOl0CVqPaLqNurE89SM7eu+Umfw580uotY
D6ZmgIpd9Fxea3LePfoDUr/ako5j8eOcCGXxdacV165tCFiCPTMUgi76J5F3
qBQS/MJarP97iDcXfy/5T2BLSy5vJfUG/CIFBipcwL1nKwlNcruEB70Z3KYM
7YH9Gus+J3B5PpWvf0ZEuRd30pbFeTCTSOwC/GI7V+fuhX+kcXobPln8+2j8
mDVwz9MmRg6hJ5ikeo/asQgSqOPZ7qiKRPW2J2SEkWGHcvC2gyePV7nDpjra
bfLkptWJElURiZdDleUOIGQrBGBQRQUS/hNB8n4VkQ2r4CtTRatS7uClRvQ5
LI5Vs3zhAAcca3y0pw8cEjyUJNXo+b1jEv1os+8dgvGCh7ith9Jcq50Wikwm
L5dgCAwAisbVT3BPakUpY2Ha60iRrTo3XV34SA5nnxOa5t3ZOZN7qb0EbXvm
6zhwvSBz8K0Ea+zoPpn2ymqmaMqLs15eVWHN+W/dUYxO/3IzVMZNbDlmnA3F
2ljxE7I0aQESOjopwuDlNi+NIXgSJY39hvalJcR3qA/R/KCyROTggvMaVmHx
BVXyoYrSpoNqtZFLwQZTEgCZyJIa/+/U9gwSSdJ8kHEYoJ+Tn6ZBlBu+tu4t
I3vwqBZP00CXnoSTkKIz/5IWCTCqd8Bc2PTT5mjEf8SCw2gEfHAIXe16KKjT
KaLCknz0Ir1rl6TeW+1VZBOrTT+MGPgr5GYRC2DbjLHGWEUI0TfW9Elzh8cD
NrOFAPzVVXm8aRNC17GlmopiyYZvErUs42cOichgSswLCMKafcJv/sXfz+dx
5h8BKm9ywIiqKXrYVz7AIJiNgVpzj+mJyBuqjJM9C0fjlSoispo2PitK1mKv
7axULxkSqUEKL/pq70Uc5D609lwXrj+AUu247qgAcQAjqwVF1UpSLSoCDhGp
Jz5uhkXI2OxCj1QyE2b6fXBI19S2m0kzMmaplf4Ap7+F8iM/CfUwuk6q+81e
Bqbhcmaigumcex3Ytp6H0hnyyA9vRtVLGjoGMyZ2XulZPKT2pWY+fz87Y77S
KyLk3FGw1XWwETEs2wlPq2Bb9+8UD4pqLqB2rt1pycOkjQNsKH1VVL+yrBdr
HkI7sY+m4VX7fIv+rB12xEdx6VZHgPw8EuTrxwF+vwzvSsF12gec0e01Dsju
ucwU0Tzyj1mEAKNF76Fdr22LfWp3jY/JmwrqS8ajvt5elOFuJkUEZqx/AWYC
IECsW4za4HrrwMkmJ1xSCeikEuq+IJ9OZFUyrU0QoVm96t/CRZ+M68gW4iVj
pEsqOgezs9MJl6Fvj5DyWUeK+UhzeUw/3YY+8GW5urB/+6DC0LWNilbCeiXo
IyM9dRvKN0g5u8ZCUUSwPbIt0EuKj/nOpE6c2bfZXAyp+2dXk+RqNGj1cSY7
y+3M/f/JqJw7wyDnhtEma0F/VqQlUQ6uQgegs6HpIQk2u8iqQsoDp995Jp/u
NF50akpAGqFEOkGdW9du6+zwW3IWSf+hgukU87jMCTY7W8RWKawalaeGZf2b
D0wt2mvE7aDDx/qDZQqHWdgKxrYssPdJi7jlmw9phtHBzHTf7qIgphbixODx
liwSdI63qqt1f2ne9IBpLw/POHe8PDoydOobSvbgtBtX44VOuWr3wYqZF3kx
koVboN19+pEuMu16Ite2xkVhvOkcwENEFSJc2wvnm7UcaO/5W423WrD5nfHI
jlAseE5MrJhMobQ6G3WbwrUzXpo6HldUOS39tpSbnSyMFiU+h84jKmcZs9O7
AQ2/tkB6SIJNi2JtcByfp+AssMhqynCvEM4Ig4oQnOWDICb4fnxv/Ogp8yCk
1+QdyOb1JBCeD++A6dwJX5wdst8LySW62OQrsWQ0EFdzx4rcQICCW8ziL//r
DM4vSCr3lH98IhWraXlazhL6iRcEO1aCh/cBMnSDD1V1zYJY3xsnexk4NIH5
4sWRhU3q3EgzU0HNbspGYRGM2yZWmD86DQX1nQcuPyRhub/4UUVJCQd0o/ZN
roA3eI4s1BYKyBKcbs+QvVYZTrbQKIZWd31lwEDpyUrVJ0BVATpcBTFbpVPZ
Ch6S6cZDj5GA+t44jVyLXJ2+tA6nzDeZg8hGPjMoWzzGPgv3g1AQzZLHYoe0
MV1jB14KyqpLrhCc4V3IYKy/41Visybpuw5CPyCuO5YLBcgwmKJKpSbhru+K
dXe4dS+zIClCzaQYYTN+YdtlVtZtZjCbXjWHsDyGS41KqkCq1QnazJsLdW20
5uaeDzO6ZET9dcz2whGu/vLj7mQKQKKYCVjGGhMPp6FpIGxOgAVHYP9WcAGi
GlfhKTm5xoXmyrQNtYmSM4H6PrbcFMorTd6DY/2k1mkJeQYe5nVXd/SZ/kIo
taDPdMDZOH9k3j6u9TS856iy/A56AjyFE0AC33BVKF2npLtgdMd5CIMOQqPK
yM3HcwKmJMqIh4AYtldkhHsTrJxq9g4uGfqa+vsXrPH9CaEtxxW3qr75TjhB
/4aM4FvkaxI1a1FYT8YPiZabkIDXLirtdOD4XnA+uHqx8Ne0axZG1Y236DYo
XVzgt+T3EhYcYSa0F9tuAKgRYD+ezPFquaNY9dOi6d0IiHABVpnM+piUzHYO
bO2RrZQT6FNoPqk3bHQUnnaA14GrXmTKpn43dfDDVI5iIFSBqG2kCWFjVCDr
bdhDunInUSiBLFffPpN1IO6o6eOx1jTgtCDBQy2pUJqIx2GNL9WROIwRu1mu
jfdr3iwtVGFItqLFgxxu4Goa9cSLm40Sydp4JPUfUJj8ywvcItb0Wi0+qyPT
qIlBhTIpfsQlhzReDK51rNb23XmRtHqcJRQWRvnVByJpjw7tFL5OrXiLCbn0
CvR6xxFNSjBmxzCoFO0Hh6I6UC9z2tqVPQAkOvLr7dNRtJRerbDUVWQqzzAQ
MNAQEqqo/1cJv/FNoIL29ZMFkB4awS9/GKbLmEUuzAhfh06s+IFjaETLc7cc
FJu2cauYJfr3R6/rMf2uCphXj3AeS78GjSsOguKwT28KNzDjtC6gx7xWE5yk
Qx0Hq/vec0Lonp19K5EYoTfegMIslJ8zR3p705srD56o3UoEfIiEgU1I2Jna
i4JnPOZNGCumhc2EmsLpiHb6e/YcYyz4xV8IRooVKl2teZOXPsxwYRN7VJny
FlzQJVC2y2vG2pp2ZDzlyadOrrv8C2b0oglBpAJD79eUuSx/hUzEpK/IWs4D
EzVnyV4obzT35UkFhBZJ2Lky41iIhfyzSPLEFZtkSYosPp+dC451nMe9pS9U
tD+ieDLQZKUqh+E6eKD7WFlPFVi4xbl6R3pe31Oo+z6N8CjicA7PGNdGQhCH
0BzQ+FmuQq0xXkN3MM9sMlzpGgCDTxtT3DGZmzZ23MHisamOSOZavPSIPAw4
8yeBj46ASF1rN5WJrqVqdcZUFAAAuOcwKJoBMGUwHL+gS8ru7jgfukdFGcFD
/DPoJpCIOydkK6MvJVo/abDcuQPECadP4dNkMKrRevX9ZbfXeTOyTjlq6+cc
6nFe6g/a5LVpbI7PL6Otxd+6frs7RvnVve7rTcOTzi6c3+e3tlYL2n+z1XWA
HdoupbO9cn+ZL4ZOp+8FxGXdWqgf9tahtOvvVcLkyfcQmSgIaqLRBAdrCqx+
dUx+TxRH8lgt89qgSVFhA4cD3UuzSH2YEqgro2eXCpKnk80JIqUaFPL+Y4xF
jqvg1H+6+NArshbkFL5H0T+WEPI54a/DDIczAzUU67u8XOV72px/L4wu7pKD
CcLSkuYoUkFKGldoSXPeXawN8XHdu35wBUuNjDgCA+S8xfxlh2DvZfjDyVdR
XiyA9zku8e6V4Ya6Zk2Vixsou2pkxjskj1EgaLIJwGEpAvOvlyBBRkrwlN0J
ATnENTESVBCm1RrqlNs1O/bT0Rg3lo3YzHQh3JqU7E1mO/qbWpsVxyzoSnJa
Bs8XI7WnghvGEgrt/p65voqUa9CahgcDOWxXbP7m1LWQ73L4aWMtQnStoVDL
BmxeUNt8ExThcB0HxQq/ZfXPbLG+PEZ4GYoQ/4D9M/HAPNIaf+SK+thDPMjb
Y3cQ+INcJ0V+krNC+RusXUm+uMhoQ+Zicr7LEzvmJ3lH8KUGE5FkqBww7cH2
dXmVmR57FW7fM7C3Ipev5ZRZWfuUdl/Z1p2LDUZLd8jRRuVyDx5uTGGQrxQN
M49exrWcx/Tl7qGEmWVJ+xD5o2qUaV2xtRRrM47SywdOEIZw5ZUEbnp3TYDC
z7fON0mfjAzjmVz/dfS15cA1855DMA+IZwQAJ5qpvTI6EorsBHTkkzJb0Vfg
IwQmFFedxr0JhtuI794MoHXlSrx3+HnkZl8fm8EPub5SLTpYmN/IkbT2fffg
STdC7ttOWmD1rdfF7s/8A62WYVpTEeDgG93p/rxWDGTuFu3OwXJrmDj6Jt0E
UHluacmHjauNJdsYb8ZxvxbhA0c0rjicP7jT+2VaBHIYx7Q5a2anTSVfkRgx
MJA8NjyyMiKKzcZOyFIiYZCbxlG+IrTQVFvboUB6vctot3QxQ7aukut870w+
//bMMcOPUgQcNWk/6WgRffsw/isIxHzOf6X/3uoTklOvF5B1qKO9c3ZmFnhH
QvOzFfdLSIKJCefLCFjE8wo3S/H+GgO6+0/lnU0tmewvIdF9z9QTzjDJgp4j
7J2rWoUyAVzSbhP+qcTe4fx3lppiAnYhoW7PYiCadiAKLSKbsUj60zX+vSeN
H+yZMjDjtPsDA0uvxLwBKtC63KDBlCFAtNcSfNoEsZsriRGI+ckBu02osf70
PZjoCP0dfBzcTeGLPH3wtbYBw8hTm+eTsVlEbZ8ghmaouQfYDT8TgluTX5C9
aU6ci7pawEJtuUWW7OVewJSDfBFoFr74DAGFKzPYA4Hp4BNdDD8OHwT4eMmD
O7h1aqpFTMKHFdiwGUjcMkoguxP6bWYlvvlLbO/5I3SP0IpT2fvZ1YXEtoiZ
DkLCRMHejnnTmtikJ/3q63hY2Ug/krj6H1K6dVaMXx0Em9dYRjXCHHR3ngqX
myG7AofhIbk4jGpnTuXKR82hgzz3Ar2CKUK1CcrUDV+wCrKd3eoyrHXrY6sF
zAKT9vKmH3V1AjU+fdIgxRXZ2vOCGn7aa1xh/kmDBK4Q8VFGdHe9otpt2V10
8Bdg2R2lSlc/0AbtrYXHeDn38imdSSjFsVMNOu5hA1VFkU1/9TspJUTFqrg7
npfpVC9SkQJbwRR28UUinxSPRvvQG1VcDu2cl6EtLGAyWRTsFLAtXVg2dBms
wcrxK9dwpgyGnaCh3HuC71JfvM1HKw1lHLOkrnmBumgxJ7ikQxcUald4haiE
oh3Sct/dH3Tfy7cLNAQiPc6vWl9SQhhhKWOiC2uttbL4ottLvxKe6Hc0DmIM
z8+BQels6SV1D6V47kekUMqE7PxD0yndEBG6/wFdgkrCOIxRoWJRGpbULwDX
xsDlsK/7n2DeTk3lVdcrY1eoG7HK3cmDnjfFdczv2+8+tfhijTMno5SDkxGT
ZQu7JMrpKKzj4QnJxwaqRQ6+jtSk8HYNwpM1cEvUo8loG//9ozd4ZbE96BDA
4v6692maWtTUO48rgIRhtRlbrf4Tz3Orav2dXIDLMlho0rlRljornusNCP1T
b9j/gBJ3GmNC42DNUrRo4cE1tdMpubzw1CZbkXhegopTJXFvCluNOty9gXGR
vSeElGQUhU+ImHvvJZNd2nWrggsO1g85n7TBxZVeGin0+rPfNCnpXtpT1Kxp
V75AqVWT5HA0vQgmicSe6abV17n+NJFpzAQAuNTMLe1KFPczWbO0vx5Lh6x4
P1r3E6zUu9e4ZDRRMmUcMmNUG+A9x9KgzNLtjRVrnOlUtWFvUZzRSnRVorpM
ezgSuXh2c+F854HFLOfQl91dLMo82hL1nCzt5198KiXok9UvWCZGDOyRjoPF
bX7IVhMWZBhLgIy2UDqC6QUaw/NGEF0JRwfdft3Wg1RIuPppCAVo1DD5t5Pp
E2XeGYf6VeuYTFIODL/+II0Fvl2twBfpaCroKYPeVVY/Ac8gEyinbuoJncgK
oULHKKEZwAB3Mq2hns/arBA1SQefeGJb3rw2eNIj4QHntYrc135KP4vsC4bB
UxiFCXb3w8zhwPOR1c2GTfaMFCyR3HZhuweVuVNE6TDUwQKcIBaBausJXDY3
0KFTEV3T6BzccIwOpSJLZuXtOgnZgRnsaJnmBKsKZi/3kUkWW0O9Ndn4TyyG
Ns1zp36tzHlOSfy2k6oKLhRHWM3fIUnToHcTqkbRxmlNtloViEpH3eBzRuyv
/uqSbwfg1sT7Ra4SHtSlxGkwhdhipsy5fzpEkUSOJyIa+DDDYxoe+m3Ybg2k
t4sqsQwviOcV4jtL+RbRpl+Y0+qI4MiEUyhVTB8PUouDvPbBr5LPmSS0VqUC
DI0AVDDL4uJn5qcIpeAERWVIvq2wNkimmEbq6KukayTXHuGHfaTxH1apGozS
0tbPK8OQ+UXigHt8rN0Nv1EancFDYAbhkggcCZHz2KP9WN5BnppHVfKy+6fl
8wlEXwQMXaxsy02/F7Tlx3Mk691kfQvBfdg7tNJNm7IOnDuKd5bZbw2s7cyN
cpM9jhyvjqmBTdkzMRDMCid9gZY6KsXZokr0xsWhptJtYkLbACdp0ZEH8Wh8
eLse8FNAQkEiQrbp/H81tWxebFvg2XpEvT6/pcbjjEM3TyQFzlaBOc9WiC5t
rh4V2WWecdsTFK+AUkVGYYcMus429+sVMH7fMZvpAAnO46PconyIMuqxfhaS
bW3Ka6L+YfUvOLmknLwQX6jmlde07rEpd9uzutFD6iuoEj1uEnH5buDFpVWo
rQIrh0RwA1WUnNcJnADVtsKqouADMTQd2uI2nLPrMvfHt8CNkEjK4shPHLPW
COXJFi9MOl2OOgEfXYyZdWxuVOzoo8c5JKhzmM9xGdU1fHEHWYEMcKo2UGdB
DrVdFVHmndY6LR+3BDSZg2WXUa+H+TGrKzfCgG79p9kPAAxI+jE0wfxu5AO9
9nex0nXwMq9lEhVmHdfSu/sr2AVsYaynL+9Q1hhyPP9gSTUrqiVxPsN5LVaR
VYz++RHqopYqDIJHR31hfqTRdp1JV9o7RVGuGwG2qKeczNU2M/wD9iIejc+U
pJj7PvyKKhYirNE+MV8tJxJO2I1jMICNsR7wVGQpzRYI53vmwNqzdIkQMH0T
fCkb7U83q7RsIYJefjHnl490XaFAJzhc5r4MA/+UxregCJpIpA5ehl08tRak
2ruJ4N3VxC7ZsUELh1qLjMi/D7mTYc7l0KBAZZ29YBTkDnGGtLVFlCSjFmoh
U5bXp+pMj9WuRAFr3h5o2KRHbgxEaFGPGmSmNVcCoIG8qa5CJWgM/go71yn/
IphGI0ysSL3zXxOGpLWx7XenFUgIzbsyErc87Lv3jS3ZDQFXGUhXmoq2e9A8
1tNPWhR1qF7Loj9wp48xiQyrOYnpv/BTpkC8ODHFkMDf4RfSE8r4AZjATyI5
i03h1gJy2Rd2wp3Y3j+r3rvPJAkQ5UrQ5x1Hthq2vqhFnqKUu1k5sJX2rSSE
oIupBaq2V/+nd4K0JJkpdDczdTSuCwJM0ECIFjIIU5tcj44bNEDyegWBGP7o
Wwex9aGGVGu+L04Mfj8a38cbDtwWVFsJ1PqFiMPLOni7bIdBscORN4M6R8Di
deiMl56yrxSP8LPECsfgoRc/mJS8upStfttOq3OiU9BCM62Unzxlh+r19Kip
b+IPOjRwM4eZkSBWntthtHXUDnw/BMQMY6TjReUm71HJOeYYCIqz/Ras1RFU
iONDKGa2t83Y6wTbkTQ3C2b6LaDNigd2h3NPMbFRulNIAaBopRzATX4Nrhqt
YZLZwNulSa+AWmas6bE96f75U9CZt6ZT6AptJ+3oiPQxOsAJGDAm13N9M+rj
+Am87Y+9KCezvqWlvP+pcn/5sUIHKHPaY019o9c4EuPuFz7hHJWDhy4LvEg9
sa37TTf6NqnQYlBVvi1AxLFoctuUfmpKlZFP5OItUn7XSf2M4n/7AuALeFPR
VM7y3SSZW3QWIsVyAB8wRtHOmv1q0p6HIpRsYZJCebAXpvoSZFGCqgdguwpC
vBYC1ZeJpl4ch/z0RMXTb6DtU79wYh8CKdQYPUN0oFJ3OC/Xvz16JY+CdM2F
/TmFivIBkk2aJwHWtK8oaERmT2Iu8JkshXPWHFSm/UQU5Ct1ZM9Zo/PT2L0s
FuIhwtL2nr42RICiCaUuFv02+hQdOzZsN3//lf3jFF/8fE6AihOPC5wuq3qa
TIDk/iEN3eLaK0Yh8sJipV74L+dshqLdM3D4gswQ5SEj8bvawwevBU1B5G38
Znd8sjXr1NjjLJr8VBjSXBW9rB27oQQrOQCZwVTBniFku4C3pEaIgZ4fw50W
Md7T4e79EbTb0nIucYG4j3z4JqexIIiBmTsLg2YxFJyOjxaswbPRezSTsgCD
OfIx4GfOhsUxYQAGarAKWnICD2bviRmG7lgY5+EgAslZ0V/wx1dHUJIsFVz2
gFv3OUXKPuO6cj59SFYBFnwdIJ2C02rGH1YDqKInSHBDlZaR3NQU7U7Mzi2Y
Sa3A5uMWGtn01lySNoMda9pB3cofY9wnsSgQ3D4B5W2XD737iQNouMsjCw5f
Hdta8WwqJ8+kZjB7zPIonAvIc618KibF6JW5rYTKbdgega4AWb71C/dGOSOB
kdqPsbgIb9+EOpKjBPkVBoX3XOGaLP9/OtGx3u7NTuarQMoZOWj8Js5vt9Mi
rQAqpx29SUUsJsu6bTlbUQT+/Uqtt4G/f+KQPsTAnkgZC8mJNq1ny2tBCuW5
yUMg4mh2FxlYCGTr25pNCzlgqLO6FWjlIPCloxl0KMLh+nMjzggluPTusqMi
CtQb9bacFG/F9F0G+U8Y5lSOQTD1OfFX02+s67NsRRsjyIvHed5SRrEYPWPk
w2saERxpdfly1u3HU98nWKOiLb7HIjrsC5nRgcfF7T2TlgNg2BzPePRyW0jZ
+WLS8SI2T5Vub9uoPAcTUgPlBuPhBwHwB/QQ6SN6SXqLGd8JmZGSvZY24hB+
qDiwaX1mK+DZa2u7gcMpU38Gu+pvVO2BEEHFK+gGMIalfFn0STOlkAuKIq8/
hlg75scexPSeORQOoINeNzVJzTbd0IH+PZW4GPR6ZgPxkYB+opp/e1SE9o7U
Hw43E22xciFqfOJgXBqR0YFLaB6VNUEw+pQSUPOBME/4Z9q2JMmlB6+RFcRy
zOg2a+o6RCAdGKzCe0+vpkxwAD/dA8YCeA+T1tzKDGQkwyd8LBKoM3Mbe5WL
pPJ8JxWQ8HKQyKTak+tOPVfOFblVOfIiV00GcxhBhjvhLpVPVxPqRQHHNyw2
TIxrOAamxualFcXGIf4ho/eiZoBx3615sU+2CAVnbA7eg4VQrwc3IzM4IE0O
YbChZVhd9ny7KcZXRfA/jqO9nSyUethpYbmBPqh0ngXJV29JHatQLnR3vzr+
Ny8QX8idXgzZmeOO5n3xndAZubqRWSwsOeUr8whZDkws7ftbjuZdd37Ssxts
VFM0mHJdrK+HYKzcf5szndV+n/05ccywLRy7nEjmY3ocY2UZO9czzI/iSlx8
6d7Vf4OzRh3Z1T5wwis4JR4GK4wdVlkg5y+Iy1837lmygIpCawL9LSSwyBmF
n8sOhYLsb3jwr/ha5LSRZOjs+RQuXMwrHaVH0v0DnkHrNJg48LHK70U9PtnP
AcmEkLMaNeRSM1L6StBN0iA+v/IPRZs/Yvgb/zfxyGuvYKb3BFJqUXaABwWx
/7W1wNndTgrJrNEwCMZrZbsztMft2+qT3WOoL8o10+wh9+yJeU/Sibx3fEnR
lW8rfS2ist/ydKcCDpBQkom+S/faLQZiPG25aTZNfy1LZWe4qm5jkZ0IumBB
+/2AlpHr/D78tsmSaw7NswmKbQX7GHHgaX5FyPtPqJg6ka2zr4/d/4EGagK3
yUZK0I0WjlzsdFxpU5IyPTjBlIWN10AfYhn/sr4d0yijpGtvWcWoru8edW+9
Q2NNLqoknKfKTfb0Gaxrx17a4P8HLlp7L7Ab2wiwRCPWWM5D5+4T8M9v7E/D
+Q1MbDAYcp24YuFV6vHSZVthz5fCHftomMHkaVIoXBA2+vKqUScIwcyW6t8b
Tk0a5iQTUWQW0uJixfYI9Zq7YCVXL1C6I6LfBh1C2WZDFP1gtvMO9g60YRVG
ybtYm/bsQVI3FYPsPAtIMVozWM0hFVMuO4OTj7mT6CIriNMcwHz4luzIJGiO
wwDtJKXh3rbZZjatmqOkVFoZtpj8Pjvt24GoN6olqbjxAM6gNirggKyjhpDa
KLT/nXc0Avw8jLeopX0GoNSlv9Pyt2txy3HomVvZdmy1ILJekBaLzifr7bZw
dcyGpA/ellZqc/yXnFu5fo17G+AwMNknRS+dtqHkWRG07kEeeq7AOcZjd2ti
jpcITuzXsXHc8NIUID81IuojyfXYv//rTYc/cEfWiYvBpj15Emxh7j13xI17
S5ZqgqEEMmtKr+k+7EkbjqD7YMgXz6zPyvSPbD5KmjyPYIPxGCBfAeU8eZUb
2COv+wqT0zwIO6KN9Lm4TdHqcC9eztYC35brkh0eZcljDGdhjUsQv8wjlnzd
ZXpVhp+xfif0tb6ZsMI7OpMPtf5NW+vhiJt+tN/pAXsKqHojXr+EfPh7pwFk
middQm9L8bqirQt0Du/kCIiJCcUg6JcD5QHxQmsn/iZWafrMpP4duQDHTyr3
/0chj7M/NRqdIGopGO/N2/YQbDMRwuLYm7p9e/70hiW7zMk4N7EFlpz1rbyp
HelwsI2ZNpcoKFaQdRh1DsSSwMuJ/Jx3cI7Wn2ZrF38B5SSjkrUuyipBhpip
7gSKFM+OjQ6jTaiiLgxlpjeLEGTAwR11sH7sH2+uQEqYlmZNsULA5EZnBxq3
UvAXDByV5ATrVkjWwvjBJZ3vO4Zu9ycDKSXxDw2ac/yhMXys+Lqwz+AJTz7J
pDodowEfgPfyfLGD7g6Hr/j+elBrj6YV/ImHRIAw+a4KFdfjIBSCYn5ceAb6
VkEmF1tHV2+t1xtWxrPGRlcjR9SUI+djvYy+8rwRAv2s8lEJ/UcQIP/N02G1
f8cTuQoB4SBOdffIA1qvBM5BeYJ7hU7Jk7a36Lj++Na9ZH3CMQyaFtssMO/7
qkwJN55bSu61p8xUWxYj3ctbbLQGF04qhoIM2wq4EUCLS+KsuUPOayuLDI/9
AFXqefLh/xmloEzHOYYfUbJqm5njU/OpfmvVJFF4bzIrkfdcYSnmsU+WdKeg
T7GbhvqxY+Y5LoOA8EO4fZ53+2aq5KE/cGSHfNkjXuSz+Mo+L9GuXB6aEOUu
gxWWK15vOVVD5QjrwSL/ORNQbXr0naJdAYvevs31WAU6bi43Zquge1tkHKCp
iZC7jddjbWJOzT6WRcQE1mge2bScgDlAX55Gztq9LdnwH37OjvBNfl6ehPlE
sF9SlgSkN6v8rMf27WnQinXhsiqQXmRk+USa+822KXgNa1hjgPIajLBcIxvk
/xm8/vnj7PD1CBagb3eIqEkKvyEcXOsnAjX0fqVayzOYS8wJ30+NBGal2W2s
/MbhQE1dCrQX2eS9IHmuq71+Uy5MCgxdWD8J67hneqF9LNohi+pKPBvZo9t2
VJqMt9e17MGpqgdKualwsLRaRXG5i05TtFkJCrrXWuFymsNs575/mUXVvEby
dwS3eGEM/EZLSdi86tqQOA+fPE8goGv9Olr3gfT9kgKRJ+etHKRrQGdGAADT
p8SR2x4ey59XDq+z2aveO/QEqwrc51DdxscJ0izck0lNO0AZ8m9ufwGRqKo2
3BeRufEzIM/N/eBKIawtTO8B02mJ2WS+Nik+EiYJJg0ZYfxTGSlfycpiZCsW
jVlCxJ+gK8Qmz1ajTKBSWXtaci3kgcZRQdSJ9vt186j23aEBxDNZJIJbLabo
B6iERuqHb0iJjJrkfTlOwEuOWmrj8Db1tQFPzC0j2KCBY6N1CpQ9zyyLy+Hh
qq+tLmXX9apYcRuti4Glni27Lf/RlzBemklxyAw6ldh9s501h3OUfZfuiuXd
h7akHffCCNdQDFy78VhBW5drFl2UddeYQrJWgHpp0qlmCeHoQEdGquD7oo5F
30XS7v0YFuasaq+PNfZvGRcF6u98Cq5E2CvLTURI0TqJOuHjcgVIa8+WH+AV
BSrKUE/ZBniW0tjsVSDJ/0xohZZp2x/IteGoJdrH7G3XAyXrr/ZV7R8VU45W
fjvne/1PnaAOlzJ+ZrWdIr1UVxR71h54Ck084PIjy+WhG4YZSiuYMNmj2ujm
dhTtAHZ3kgasxu1j3FGkNyDypCkTbZdyy2+LTMyR97bBDXaMm94O9ulbpu9u
Gi4kaF7AndKHZkErZ8yUqk0CWLhtGGAQVB8jgLQ0sD9QvlPni/nSaHfS9znO
YSMoyfF9Ept65dA6eT5h1+SN4mzDNtGtdW5r1/dQlaHu8UxJvcdn51q1dWEn
jNmOSt0tMrKCeWKXbFuiY0nIgCZ9IL1ENalcpnIDQuEUyHy2odobZWMEqDmn
RHiV4kfuIY2hfofN5CXwCFYUOwC8agl5Jl9k744aceXghcQGPGSFk/I1Fidr
sRqJ0ux2dsn9T/2Jvb6vyrXf8rzWkE0MQWtRFZMToH9G7r/eVIhgShNHL5jd
PWWmks3bsidHkUxHq2CEZkidP8u7qlm7OuO33HGGjuwLw6Bj8URbhEQkEvcy
+Q1tJyKuTuGIgdju5PkooccnVNhRcgRMj8OQvmxck7r7vWSoqek1k6RN2ykV
43fCDpAWKS41wNv6R569i/j7dWm7ykmHlBRn1rVx9YEForsFSKp4LrTCpIHJ
/WQHopVvUe5LIK7+sQG7hyPnhvbHHUNwYC/nU2egdX7RUihPovjaVTJL7g2L
vCPTaUPlRV0qk2YVIo9DmYjL3hEh66DOKIigs1fGPQ7itEQfiDp78EVaW/N+
pS/J9xjtwlcCMtewo9qvQFXNJvYGscbT5bHh8vRfzc6JAb/nXyw/Q2+c1HDn
MmTUWCJw8EbhUf+zC8E36FwLf9KlMYhaOg52lGoQ4Rcz2P6JsITuID09wcFv
whWnr0RVAnAyaAMnUVB0WOT/NPUACqIIp9/f7TNY6XVavSgklR7crhCFpLn5
+gFx2P9uPbnGYmKOU/rImuZVP1CuJjHH0BmIJ8x+ZQjyH8VM1dG4E+PMhqNB
Tv18o87/dy5FB/wY9qSiDS1wSjqFuK+sLsv1mMfpu7+sNxoFi7H32m71PuWW
VZ0Ocwjh8iHHS4UJbdhCqjnCmgX8gyl0OwPEt50GAEykZqTPlqHWR+5mqSmp
N0t4p2Dj93BOLAoeaHxqH/z54dLp8dYOzOqtlu/9HqTUchFmD63TheNdOkcV
YUod4OKL3cXdXd/CMt86Otu7XMfqifEHn2D63cuQijO33ArgaAO1nO+r+7UL
f0piZAjAEsiGN9pJKJ/cFdxRGFj6dX2aJi+Nk+SeonJrIS6scLXVDsCLH/bF
J/U3Ot8fJPMsGq7x6627SWyp6eYkkOgmLapPdTeXpJ7EG2f5nH7lbYU9Xo0Q
FPlyDrpbuP83fiazuEPD6sH/vM5m16GCAQYjjeXvicRbv2aWMqL0QQow6hbg
8YYeWd0ugO60WywwAffflMJolHpq9U97McuPHDzWafYX52WGUrrwZSPDSZVt
SHVLDX0ez7beSifl9eEOkSQPFKde+MHxGE5/d927gCaVUJhJM1uwfyw/MM25
lmPA+n2j/vBlUKOXc/2yxgYnHRwh5QqeVK9qmcz9RoETfmd3HF6vCvWGDAKQ
CK83AvQbObhXdPMokA0lw18SwZ5NHr020lCDee8tuWCjxr01iGpLiGGSkiom
G/u8n7CRcTYo7CV5/MUtbQAmoibCHP1uiLRimSill/uSN2W3vCEpTjygFnCR
ehbsrO0P/UZIhOKSd9mWVEifG4JTTMd7Dzp382UgR3nvrZl0SKYGD/se/4rU
MMhqgsW0Dq9oggeWWkNHZt49SRg0CEgB0AOXvoedxsb4igaRkIeUG3f1W6kh
b5uJ6V4sAVgaz/Elm9cdYOc0yyrt7KNArDGuUZIFk+D4JEYx9vEyk/SEF4xp
2Cjib1YxuTQy46N7O4FCGm3XVFroHQyKsrG7rhAVcMwOnNrY0MovlctJIJk5
4Iu7qWZxb0q6BGhUKSUkgLPZW6oAoQCECP84TOKt3YLx4U0EzuLPQoRWcayu
jiFtg5/eDLAVTeIRPSqQMSO00CDoU2ynuKyru9V4rDTB7VDiAYkv4YGz9W0A
jcr+Wi9Ko8LwhWGuLEqo9pElkdiksL3lBidlgKY6bePxgvnxaB59fd3dbfdJ
A5ncpk7uUfm2ejYno4AB/UGyLbAZqeekGQ+xc7OJEqzrSOlngck+qaKd9STz
Vxj+IRyO8Pt+pT5Qzo9BNx6pHwZQwZE5KCv0HfkN8XdihEaByujaMWHTLrBf
5Bv3wlsbAhP5CsNLuSq4hF2lKBWU6OkMsyK6pysKX6qqDYpD4qO9RXRD32n2
KEXZ0y1sodYdWO/MRDqu//ls+5xuoY37lkR9HBBVMi8O6XFK+0Q/Du57jS2u
BR5uXuXC4mpqAHSBSqPA+WPA0IYa6Sp/9cxBrT4eUqfcuqbMLfaLXcEsWBXi
kJPOiYisusoa3Z/OUrOrx+5jGA8Y5777UDjUBwwl4+4XptK7+LKuu3H1iUvP
c2E0Z6JKHrYk0nj7oZoSyD7Qra1BKLETvZoSdwxyj3cmf4yz4iuBPt953yjh
ZbOue/s5IrLKOEG0IgG6R6THOJhfZTOSe3yqCbo65zliTQpLGEia0R7C0Wcx
+f7PsDkPqehjYjH6qaK3spglV/mWgsC6GJvfgZ1q4ljJ7ks5z1jvro1ULeAx
ZePbkwEI6DYaKyr8dFNt+HXukqX7V7AyjCLEgjwhaCyosgejW4k8YF6WC+H2
E3rJV2zvTRut+YzTHdvAFUVugx6quoqZHNuA20vuKcz3A7aZ2mq83yI18Uqc
37mE5+RcRzI434eq9F4Oh/UlLdu0diuP7QWCvFxe+OZgNbahb4Lg4ik8jkxi
5ZdLrMlCuX5Wk7tdwCGDTytIP6sZhbGPmhufash6FDwPwYo6INJh+P6KVK6L
HpENBaQZb0PfOIWxw2Q4zGAb2YoZDRij4guUxdXfZw+9qw4MlkTFtHkRSOZB
Cv0lmKUAnv7er9IF9hodFklymQol1NTsfWYkNDb/9Os36y0s6CH/KJU16u3C
/QNuUAAjJmD4iQdJJi9Z1sJdJlW+Yl8mug/W/gkpwP3lfJNY8cyGNO07oetC
/YOAQv6+cTvEqABbQ1DNL40kJKowVKoSRKy6kkK7uwIYWPLQ+nq61f1SOulT
HO9TnPPnEG/HU0rRJfjB8KmVcQTmwZveOjrTaqyhqqtzEj18RpmJ/d1ledA3
CztBvRuvwii80dzuMTon+hG72jwlQaq3sPiX4hl+mFajtB8kqsMcQieT0tgh
1BJFmbOoVpjHzCelY9fLgYyYu+8fg1E8HSd+V4VH7vXLlsNfGhQQgupkrmWm
pxzFrjt0ctxp04SzPGBGCFwQ6HKB12Vy+Ml21rxR6ehaPTHav51SZ32d4ssy
+c+hSfdAFRdRbR4HIn+7v6dAf0fbfLJBev7jziRi0JcFHOH6MlyKsmLvcSNh
LTOazWTV6qg+YZ+S4OCM22FVlPGcgt9Df3zcKEE5KtI9XF9NlJsJqqS9HSFC
y+rEloFskJkIKzgtiqCICymmWWSa8x3igXLS8aT3/BF28fRV0uN2qoxHHU+g
vvG5zXZFKPP+8qnGEr9EJWeJQFeTJA2uczvROYWlnxm+sTbSWQTue19TbC9J
YfDN1cYDJMq40VOBf/qhwOr7PP1SpcImyXwIVswllSVwRnmZkieVQmSkcjaI
IDVLlrWikfk0Oir407PmAKFwSeu2xl0O3RmFPsk7gUd9OpdO+NU92Ee9zQLt
lL90fi73JG07LxtsUgSqmTY2tAS7FgEbNlkmESMwZMPLy+Ldel1vmVTouUaK
RE1KcNt4AG7T+1I/Q/UZQq03ftGg3l1cb93n+RX4Y/zfkZP4MvouZiv/ACO6
CDD1nRHwKIk1c0bqDG9jJ8YumDF3I8QmfOO8O+6HZe1WZa8HGt5Ys07vTlii
mgKuEhZOlTTOqRHIkZiRlKWOWq9SAwCzyLZngkJa0iKuhR3prgG7aguHETPa
gb1qY59X5aSAFVB9Gckwjn27AOC3PlGpbWN50lac1YwFiNpbIUsCPltquMC/
C9CPF5a82+Buj2ySR3p/u/Ka3bPxfUFTcHFlEerh49B/hhH/nBTt16H/UmSI
Jt9rQwRTKLMko99RGiPhghbrkAfdQ72Z1IsOZQZeRrN3cJfj2HjjTQ3FsgUf
mdTz6rV/YQHHt5D1d9VztwD0NH1at4eNH6Q05bZcRxxSblyW9Xj/eZTJV3AC
O1j3/13nCdzIKuI25EvFQEJipDjwQIgzXUIXqdeFAkNYIpIMGP1dS6O+uGUk
nkNzTIJR5VVRzZWNQZKzJ0JUhPFjOsyO/3Yg//I5Zppekm68gY0TFctWNwq4
eJVIOcrhrOLYasknzbV3LbUOnL4tZBS3hePUyvJSXJQMggzGdQF/lrH6XQcT
9RymCzUww0OMThXaMlXN11pT0agXM8JzPznYxI68U1BiGMjxFktOszAoM2zf
FoNcDYpxsJZIPwjR92K9U63TObMMYFcXHYhGSl6w4O9IopV+ck0SDszKsljV
/JBVvkChw1Y7XPo89ILVW/6hvGrj7vEBZCwEqm9PlnzoTnIYH+QpW8u7M+M1
CghfmiJMwplLQ7Lj9H82WFwzV4Fc9y1DHu3/9VR49r7JGbOMaWX8E9Is+xKv
2Tpxp/4VeqAwPepqPmAD/2nqCF4zshVjv9Poh9TMOz6O26TUqz3phws26J8T
1lrG400+KjnvA0qmzF53xSmYgtoCa7t48qes6NPA6BAy+OjopfkpCx4ggQYe
HbEHbBAN4FX4x/A0FCPrxTCLlDDbuxy5uM85OINwB3D58BNONebD+VbLF0nB
knFrdLP7DPFpVqncygAR0B3nN0eq8wwyX+r9sOLpoarsv0rvYG0swJFM/1rj
fu3HTa5w+T9sjQYpofdDTlleU4lx1bA/uZfao7k0zj7+fM1VZ7ir5g9XoSdV
gji3KNBHmlcq8/Yu4F5OuBKUmCSj0Tm1ShSXHtNT+TFAX6l8pRFfzTD/u6tl
zP7H56N5cx+e48S5uGXatu163864ohubOEfZnjiyvpgbrTGJV4/Hsj5wG/NU
Wuctt1I+aDhIYXnYigZbjbJKCOLZaFtTBWIL6h7vhbR2jpM/Kzzb93C8rTzB
l28QEl/rfmnos0+q0uCMTZqqiHlpn6BX2UX9b7L54dIfXglzvgMX/WnWryb+
xWU4j4Hm9Dn/1ZJEktc5Uw4KLP0ZqpcyFwB3XS/0J9+an+Fa+RBwzDSCKLMp
Iz5ppK7NExSvNmiqguF+PsibneclQrm5bi9WDp3jY+et1IFgLu+VY1W3c1DO
Hd66aLBR+I/TB+J3Rdj447tXsE9HpANjqovNeTYPnuXBT/+VoQijFCCskgGZ
ZueDmIsmHKSxJgkf4Nf197NnRRPvaPb3h4j1lCdqUjL6OD8ePevQYLduBcyV
opY/xw048QowLp12XJobTLKekkExhcHp0hKNrnXiEsB4rjpjFjOuHIvImrSQ
gU8sgMF0M/MtCY6NFIq43v/ZZK8Kscf2tBRmLYx3zDRF2awI3SDzYE/OpIig
3QSwG8ylSJF4qR4uBqaNEMavrYZf2+HN00OjhxOzQv3TC7SiJf42edh2RB8G
WJYLjOuyLoGESfqmlMANGi+CYfIgwhxMskk+8QCA3DszcGHTgLb4WFhGQwD2
weMjQdsYCFU2yapyr22C8OlYVQO1EtG7jUA8wpG7xQAcH/l+zzWLIYElFqh+
dLmpvkOyhRu+Cs6MlHR+uxjRhsmXIKmRt1q1jT1TdNd5Ek9sLVVX7Lo6Y8aw
+3RCHvCEbWYYdMvpnJe9/xhizmLRAVEl2SYhvxWPb43/Ar6W3M7MLlcIm2D5
xsQnPSvwvboDKKKAQBtcfj/sz8BHMBBZtru0xyz79yuw9uhN3fGMhEFnKv6H
mYjg2MiX3jGN5saPXDceA7tR8DTrzr9G5dITzK5q3ucypbfWB9ZYB2IyMfi8
QIb6HPY0qeR4jdQJaQ0KMhXLED67HU6JdWBtEwjXHOQMnisJcMKp1uXFDDRk
IaOl4msxei6O+uONc9LeYJaTvE4Irhakqu3ArrLMP99LqcHtZZUm237sEUvf
dGQFN9+l5ZEVYs2GkKHsYKrJTyI7zZeya7qtMtOB6jKmDzQvZzv25c3sf/Zj
DWHHmEWJJfNAaTen6c8gBrGPhUSnc/8d63SICPP6TIP1T/nO4w/GAh6hCuTq
fwxRHmjbbV3Rr+mBULOeBNQxfjpXczHtGoWgVl1Y2dQPdfMKsHdBrHAk+rpo
RgxM69h7w788B6P31iFW1rbaIK4mtVVeVdfjlwswsv6z3kWavNd3y72fp+sF
RDO/D8gdfkX7/+6WD5waOm8lA9uwW7RfKA+LTrLHs/t9VS0JXiLPh7bxOyFu
OvxAtGok3JT1yJDgdMTbTrobEe+bmDRCtPA62AuLDcPCeHVrNHM4w5hWyZ8W
Gg8qFmY+pV5NnUB3iIqplvZOGTwbHfvfKzr0FEkrVn+UjnD+eZXQWtBJNumS
93854yYvbzhUwQv1lQXkoDIbWP6Kf43QUotj4ed9TrMM5MfA47ZFO0oDUN7O
4VI+dl1hPr8ON6/LkK+rQ9JksEIPcrOD730R5xnK3I/3KwhW9oksNRvrjD+h
bfJi94p/HwxZT8RXs7pIyTHRXi1lYav745yaue6NxtFyRb5NtMbomNbtVo5u
v9SpLNxHON3WQQaApAUj21PitLTWOCnX50ocB8MlsKIjJqA2Szga3vdbkBfl
6h4wwA4T7XEjlbP0Wt4B5vvZmzQI0dSuNGYiPkcOVznX1zGIoGXd3tG89z40
DvivMbtq7gus9yhX6zOUwCjuPtKSafB75cLFys6m44FyDbPJnVesfSTMmXoH
T7OpE0ILi5KA9w/9LPD7uy77PvHQklkfDLbB0NG11QAUM7E7sRDzqGXKkFXy
cQh1WAYFg1XAAXy34/QIDd4BrBMzwnolT2mIkC3UhXW1Ps91zKIB0Wi/cJ1z
PnYsKRavKbzEgU9Bim0vKAeTikTRKJXqgNiSZvhYIgLHyecHSIampJavKDUz
TRaXxZPNJiN/5PVl7CVXT6tutVLD50sqZDz/pcrwPGbvtTyDFvJF7VLpVjYy
O9dRGDm5gaImN+hBJwvnX7pXYud7cMTIDEzzJsIaagMZr3aiWA7IHUlW3PmL
5/kPB2ljuIsJFbCQooV87AkhZj9p2Cl1+QXZ1oH3qy0QqOGc3w25CZ6goIkB
9O/l0A8Z6P4O5aGbckmtCPtQugD98m6/2XIKRCJsZboRl3GRaqrrkdtFoquZ
QaUf3/lRLPwCeHaBeaNarSjA5AZs6i8LAe0dPQNfzJdKZ9gC0qIOA1Iu8B1K
lbcFME0dnooYUm0Bd5kBRZJXNR2SxtKn8O5a7uohB1s3iwHyDFuE7S/LocXk
6ycDbdet14ciiYaodEw1qysctPYByo5YrLBqeOKibLIKKRv3j7MW2xRvbpKK
v5EllufbJ4BorpHaGD3Nhb+5AW6HyAZ9By5At0ASPJcK/14VkCoq0SiZRC81
FRmQQvyUy612LcKpeyp38xaSW3gIBbpeGRgqidjdbQd+RaTrpwHc2J83g4t9
3npd0DfKoKU3le9k/lNeTbUTXtklbAcTJ5RfFS3ducsi0H+KEcC7tRs7nOgL
K4Gr/oAB65WcS+XHKJj46v/j0eRDxmWqkIapF+lhysr5kAeRsbBtcm0FltbW
QlQIoRC/2APrP5qKp4pG1uxxapBdrDeaSLjGA7QXb4AKGrbah5MtadLY4Ie6
rffLwX3h/wHL3TEkEnbdPQb7KnAGRD/0ASzTMvC6LYGZH6qVDyHwlisUxMMt
BOdwRUCcMS8/45UAwsT21oXDfCyHNEKOCCMhncXFhcuJo1pRkNnpVze1e420
bzL83qT7eUs35QN3aEHckA4YfZjGYxCQdTFEmsE0Ihc81T6prrDRE/0zTV0L
BawYk4hAMbxU5A6dqaq7MiLYqDJ7xESrdExXbi8sRy8BOVuXuzMJziIRQ1gQ
3R/bKKe8cN0tVWgoxiyg3eoL6Oju/lfge8yyDeAFE2qXpmdj1PxeqOoT+AUp
mtZa79tTT+ntWN13pEgTYQznZXJv+mZd6arlloqX/7VlF+tskM/zPkI1ax1t
9oT09HdlQ9pFY7q1LWhKEJxceqMDhOvfKCkU+g5MR7dYqChCMA4oUEB9JO6Y
rUnulmAVslK0u6AJ7SudGScpMYtM7lLz+ZmleWNWBVFb7eiOWaw55XUcr+6o
+u+7sTCcDBoasEpTIUnhUUnzSle6XQlSRSGIzMnkrk+w+mrmeSw0Ij2Je/MH
SNmIBxezXiAyNuEs+N9NoJoYJlln+sKni5Umf5ca1J1md6ctdBnbsHwaYFv+
UVgYK59xfjOaje0Pr9aqTm5SN6tXuL/PtUYcF78n925Uiq2j/Kna6m0SdbNb
WsrEZbca2Qk21YrzrLDE+/FLfeERD01iBr60JAq/pzkMh0ZvwTumLFqjbe2P
Zjhw45U4XCkpk1deq9Ky1CgUe0PwSu7yoXlSKc3FbbwCiHaE6hDc4TfExfe2
v8mXDroV2ld6QWgl79mwl+dbOBDFbfXGFvFn+0X4rEE20Fclnji04EU1zfBh
TTp3MEGuP3fB8yLT7UXeZl2W2SN11MxGZ371QSJt2mIEhDcO/mnVOWqrIyf9
fLAdZJU8wm/+gmBNcQSx65alKPsI7mcVRTt3LSVDh3by5SG5RdLECicEOLfJ
NOOocnCv0sQN3crW4m6SUUw3w+gZ4A+wNzIYeD9AbsH00Jshfq11v0s6boNk
6nJiXFiJELx3etuIc4Z2H7mj3B8ndfLKF2i0v1UIRtyLIOYZPENNuQxMSdsP
uhDgLc6yZakzudZ277+DtubSYw7dLq7GJ41navez8pzSXnTBwBxN1bMMRNBN
JI/E9sAx3PciJpa6vkpXwWmM0vEcfx6UuFotjHPcxnuuMRAk+RrY2gS/2DOY
EuuElLYhy0SuzpBZGDdcx5/wN8abYdviDTPNrGNHcoAvmuy2vdf6f0er78O0
WzHkviUkUx+1EJYjF1JPoOvbQJsF8VXAR0ONUhmleo7S/qdH/CtNXhLDx/0a
2h8OOmzWgP0TV04w8wBH96p8Jt1vl/XtO+0u3Wmxlv3aw80p9V0BF1WHH8XU
jz0xWxyV46GCHgAuPUKgNAR2TWrf5KdDraD64ht+4zR7DjcF/hmLJrEr9znx
CBYK8YrKd6IU4rvmyZ5LYV2xTd3aC6DLZHgOj8q/Q+IDzXrK3DE4JAzBs7fv
R6IbrzuTwAcfYbhQ7oEtyrH2r3sJsKWBCQFINsh+M/3I6P502Aoi1YDp3H5j
bBAMDUyBzCMFqAQCpU1imwicGhq8PZd32UhI4yTzI52TyCSRS6yovPZ74NDz
aILPwq2QRkW0eKqYmLoUiWfAFx32M1x5Jv0DJhFiH8cJs3dzdA/WFbJbFcXu
HcljXvL9GsL2MxERINPGgc0eTbgr2RvdBhvgMYPJhsnDt1SH9/rl1MCujmMD
LlAhgSVPDLwt+tDf8sissbotXoIs4mUwKPaGGxxIi9OfQTeLc0mDAEeODJha
T3iSya3yxXxijJ+S+A/CK5X7iw+QddaqRakyvWrZZQauiLJBbNoDiCc0fhI8
b3fEeOO16e3dLRS3Klpbsi+KB6osX30kB5Iw3VdAE+PU53mtHv+7zmOOyAQC
F8dtf//AyrwBRyyKgJBJVrR6lYZbQsD/3JQy38/cKiI9R9zmzbZ7j+UrFk6p
DN/PwJJPkE4CsfOwsPCAnAiUIHv6E/PWVeZCvbLvLp1uOqaeftVwH5CxiYOi
tbmmYTOAzgyTo+Mn3EV9spl2Bp44AHeD/qsF+INBx5YIfU6pmF8rBy6dFulT
bHQ/cKLeMt+uyLpUPmPYGgKjJvSLGij5J4AJZcDo7qtpnWIVG9Exhv4yQpcm
SXxfOR3r94BTV7YJsG5hXC+gZJBVqESQRuJPM3liQUcGJFazMUpE8tFw8/qE
M0Bw6przocg3UrMWnQXyHGyokKyamQxbWcTIUV6XOy4KCQSZ6TFkEpd5JeHT
VyoXXjT8qN4xLUJAbZTmMIZbbGCjbcm+gTZBQjcx8/fHE9PnPQtrKU18dEUJ
zcgtfx6468Gy64SHQhUBgAalPLpVyWz6YPCjdToEYaXZRL9FIOvtsJvLK0mA
l19t+xaOheIFsun2YqKR7u4L1SMgG81kEsnUoQN2Ut7pu5qHPUkbhL2Lf98s
7MIGFVo4OBdePO31SpSDZiJPnuDXSZP7X4RXycSa4tJU37Hph11qqFwg4lVN
8HaKszRj3HfkBkw+cQOrhjtFUZkal9KWdcY8XA4yPE9DWaSmk7Xqh/kotOHx
0B2qvfgXHDOiK6NwhZJih1GZouV8q+htaV6jTG6KDh0srxBGqwywvEsVHMvR
8TcusOYqRvCidF/yyTeU8uSH2mxfnhPaZzehjiWFay8LcxJbe8Rlvic2f1vQ
V6Rr0PVD9o7GzdAcGvLb5MuMJBGpZe0O0G9x24Y/LIyNBv3APLiEDymRwQrV
OVtOnr79fDpdj01+ViWFefxLOqt3PgU3dz/RURjh6FMFJT+XQ4R55HyqTbvm
dB0aQU22JV+FC14DAHf1mQcxUoIRsOx3aGdAqVY18/J8puBjXlp5+8c8lE23
fKjP+Wob9MsznPeaCJPEmLNO0QsXWy45tsoiwREPTTi5xQtMl2OEgWhnzQ5X
jmD/VbQQH/q25+KCi3Qak8yEIEowef9wmdTLO3QThDNUXjdcjQFRoqh9OQzn
mwu0Md1FgKiX2CDXfNnbbKvNz4hTTpZaNjtvEX1dN52F/cQHz7Wwv7bayj7R
bQSjN3617EoVm3luDaac4wVOPVrvL/lGjX/lZWM4ZmdsZO5G/DZMnihGRpg+
ReDOedKJNB9jrD2NSNSRZ+5JOB9XMPPCEHfdZkkgfNVYa7AbJ9ZmnJBwDyis
CNCaCBEzpUctjTrahLrBpSVyFTYxZU8ftFr8XECOi9kJJdF34vjxm9vXeyIY
gFcum41KvmToZdP7Al/9mqsvjc6RhkRQE/LEnKy2FEHJUSQmmIKlVP6Xs7RP
LIqKHlMEkt6YBUnc9J1f0rMyAnHgk0gNIctJzEV5xEPWp33Oc7/TjrUHbB5o
zkFJMYaA4lSeWCKnc0sa+3dWAaEy0oCT3VmGAAvtm79/8oh3Xan/5JxYQsNK
W7FCmZFItAr7H7HyHbwCUOMc+WnwUaNvHaRvYXZDUsAv5Sgo3F0TQaQpJ04C
2FQQKbnyNJbS2TskQdCsZt7JXUaSZxcFhAioMzIQRcVZUI5L40fF0cZGeFVF
TMDshtuIbegYbUVcM5r3qXtMq2rlhMY5c1cbv4yELcw0DqepA5cU2XnaOn6i
v2uv4wS6YY2fun2VzLCKQghqjhCdML/XUw9yTampsyGlIo9IjGEZV7b0MFQ+
JxiiMjSH7Pw27zo6N6RHyLPOINOQGZ4d3eWJdnTUWSAr0SfqoROaTo1PxT/7
QDuGFCCdjrxjnFhPF6SxbOrPy5OcJRiWA/+S75PvK2ZRqTSI/ul13WQsQg49
mRv3A3nsqOKlTxOTgcU8YZaIBK7LLH5PKy+l0d7+MJQFVEmkSOC11JvtqvFU
svcEAfRrBUoleXXZACjrbzf00KPJJCl/blWrqFLGukjgYi7ShNu78myazdvn
5sVmMMgf1QSvp9YRRqxpgldtg+VgIYFV+XqsFOp1ibyF1dMV4btxWqQv80Nb
Vm+MV4WPeHSpmtQu84nPLcU3rM2ASKMFUxd29mQvmZ062wi9pjbPvoXUnXAO
ndBDKGv5RoAcqfKMcSyjHem8Dsk1iCZ/7BbI1kytTZLi6iKAQ2LlZ9wPu7L/
VsHIk6mriNtBQtWXO2wkVXk7HgZed4VofE4l1Dzb5404Jdku480Rrr7dEfDN
D0xQ/fUS+bnOuS8qlMy0cNdJj054aFme+d8+Yrawa7lxxzBjqMPUdt5+kC4e
UDGuXiF47vHZaFCKE1HXCFRKTdpYD0WPfGXK2RqTEtgRHSKOOdbglhVJCaIH
S7W7KK9Et6+sp6vzC5af8pJ2t5BJmrsCR+gQ02yZlxEqxcw9odgE5YNakFj6
NsGLI/PEWvvI+zWgkZd3PZt4SAELwm6wMJlA4KfRPxJwgqHv7SLrkembqGo5
Mp/Ks/T04YEIug71zXD3jKoUw7jVGOJW0zpQnSz0lBB1mCqhUwM7uF6hr6zo
KTN890zwCYPZd1EAFLPpDUIclLF3eSjvq5S+UlimYMLzVXcBo/E/voBAXVPv
IA4jv4nYK5pKa9+oVOkT8Fp0NLMTFDZ8ONiO9gHbRnxJHUKsuxcghSyBbJ0v
bc+TjyCDLop7hJERE9BjLY7BEwkMm3s4LYyZbvp9A/fe0XT/GDkl/TdEJa0f
FHhooxCc/Xn0BccIFrhACApxrZsAv7vPpIx0pzDWZ1LEhv3QR+KrH1Z7HS1s
bWPpRfb2SpdCMMGyo9NDL8EdiGdInaO8r2kTJhoPd7mgEPvnC1lFMX2nKR2b
CbQtoiLQTH4c0tVA+xRQ40XTMWFlIq+szpPf3Ovp2ub85i5pYw+M+oR+UL7d
CClLAMoVV46gRBaAvT0k1ZVCdr4YqEzbxttLDzVDN+iBET2YBw4QNC1TQHQE
qe+CrRqLCKMpgZ0N31/x7WEduVNZlm8EM6h5JBNu13ynxmvaZIVActSj750g
iKMTMw5CPmXtYq/S2BUtvcLXfyXorwFyN6eBizwF6grZN7D0jybD4xi++UMU
17akFCWRxSi0iFzk/xYkqr/q6ZUxkvgYOi/ejiTepoH2tc7enPBED8TUFYrh
Zl3e4hNf4Rg4Kiv1xjCZEARoavbXJcadq/UcfN70arXk7FfNnmBggFCMJmIF
nsz4TnnWuCwmLeKYs5auG7uRNTFAwO4wm6IkWFnoLp3xYyh9VbEkEFCpGqNj
4F9cI/R+dUHSZRmlF8fauHFjBKmh9VL5BE8ZDZXxf9j63XQ34yXc6mCejjIu
pUNIzH7+WobisRshwt0bfhEa3j+PB2U8LgnEKfVYdyUA/etYjOuBNJL1k2Fm
gTd6vIdHF6KPfSwGyUK6jOBw4Hm75thdvTxrIejf/v4CDsgCcy4jn3XrbMnb
mo3GQ+shpeSvMTBWCGkqJzggva8lK1ccuDS2uJy3exngaCRUO2GzFnLbA6H2
OQaE3ONKdG8Zq/N36la3Pga9Eg9m8Q1OnwGxq2WAajAyHJKz8z6uOI8OE5+i
fXi7N2VevdeKIKFMggGpRb71zBhUKE6fJWRjRO22veCwTEqst8nb9V0t23V5
BxiPVGCAup2CPSTcUfV3tn6G6ndU+0dlc8BOU+f8LJsqDukj+OE85R7osUxX
DoJa5VLwmNEEgj8hhFejnUqX4UJo+C6PPzMjVHYpiU6e3KY8CvxfPDYB9tri
5ZUG2npV5la14IROzz4KyFTFvwLmZsXQ8ShwQTfWFRzmO/NyQ3454SWCNngo
gLvs6qcqXM5voicqI+IYBjKcMIxFkShXk/fShvrkb89GkkENF3yLcAqJhVua
YDpRshjhYpt7omvbfPej9+e4ahj+eD95lc6rOz288RLDIaWB6eZS2d9klrPg
NjpTEJ1v7YneoGSbWToXAKJ7wXUinhFAxLT4CkRg3nAINsH2kG065zaVeBKX
dgiQCiHoGjV1J7rr9MGV41V4Xg4Lqo5CIg7wMlWsiIP52I5j05ubxVfyXIkU
+OaJ0X83sMVIV0US4T2nkYTPVQQeWYT2QET7n3CH1GtHbMQydcDZ0NPVAcYq
+hPBAufDTU2d+bRrXs3+X1OqLtfGUKJRjdWOR7nxGfidxRib3I3dXOMbj8WX
x3pisVWUozEyZmd30gWHrv8Jp3xWXi4v59mdepdc2pPyU16zXd4mbPEixqGW
EbCIBuXVevBhqST5ifIkz4wXfzOXTKl6RfF0RCI4CaVGRxC92YOqNj7W0yo9
IuftklvJz5zFv/fRK6BnpQUBTmFZ5u8+sAfZ8QydoLyXeGQHACq4asW9JgMr
HjVFRmu5U+1f9RA8kGxO8tX42vescx39JapLXafkAxzY1oVtlRFsFiLbkHBE
GTvD0YbLBab6i4lXOyLiAJfUgFHDD0v2jtTBWqtzqh9F8M+yB7Uqdoi+6LFq
7LRGJ8sEaKDGXGXs4wUCk8or5VopZf6hGo3xK1kZmnlUVX7WchexLxLJhXL0
PAMiN3NylG8jOsC3Copn0ib0t+wMJg2AxaIF++/jKGkvBujnom/z+aWVWROA
iGv2qpnKd3KFDuDrAyBy4Zh2hwbTAC8+IG01Eq38EOyk2E3y5snpiyf5ApDh
O03BdDAmrCUZJc8xGQl4FGR0ljLU4Zq46rGZZ9Ph13K3D2UVgPfkYsbMnm9B
dHwaNW4oHw2/laEiJp1YPPmj47hg0jm3PdtLIy/2InjNHv0CIliw7dckbKn3
l/8Iar1ffcUtjptblRNWumSyGofTTFqpARftp9DbMmWIZ2ZxZQl9afZa6LVB
sUb5MD8KSvMvaxyoHubc+ZW/YjihXy+AdWbYmvveSsk5cOLB/751ORmtnUJv
X4anxf1FoHdBxa/PW5XsdGgMPiGf6uWMKdcaf3ArMEFhLkEa2W768gddKaTN
Enu1ZiYnUOIhWiv2dqujCGaYCLyqkGeTODc8CMaPCocLAtCJWYsP5CIbM25l
LvQvsvVMNQamOKysx8rbL6ixWW45FjhBPXusdJ24Y90EN7PbfCdF6jBR3LvB
XEg60Sw5JP5GMICod56nkqQnHktcGSgeEyhGzfk+w4901WSb6olT9bW8fuh+
xWZWfmFmD6jJbFRm6/+A7ZUdToDNkasTE3kOj7MJR7XvYLRr3irIqjdAt4bF
2FBvHVni5+USYSl+ROWiGcZkdoxZ4+i3PSDvOJWiYWcOldEcfpuyJD4dsP7R
6D0pUK5/cqa/ua4h3y/QvZOV1jjMqc9akM8mF8py1ABlFHmpVlTH0p5wb0zV
YmLJxqu1QN40h9ph5cxEgIONquKlJgJY3YOPRDnAzrFpDu/nn/In0RYc3M9p
Ax2YFx8VFauKD4CbB5QtTUgoqT1pZYV48qvYl7x+ASso9n1kSJ5TU4l21LZH
aiYXH6lRxOaXgBKxOxLbL34akWGmBv3ud1sWzvnoiXQ76EahGxkPl2VYI5VI
8BK/vDDKgsgEv5O3wViMljoMimG35x0OIC+k313xI6xYnXprWhcBFBrt2XhS
77ugrRepF1dNMiEAYd6OZs6+9ex1SOtF1JdxsRZ2Wmk7+gRqJkf5J2zuM7hP
4LcSd9drcvbNvj3JRDblQS39YWZyl6+JhZfRoNnSMq0hqfK8ExmMi+GpTPo1
9HbhnuK2qCwy85/OzkUaRiLXBxHf7I7h8vb5Xvvc56rNE071SEF94Amxtfh7
OB8uPBIQaQYnkTRM1BMIzb0cYZAVWipCNbX/y/Hn2qOugKn8tC7qjNAcurGS
ZWUu4jAfWmzsRhBnTFdeTuvFG2ypuYcCNPkm9v4Cou7enWotLCpvbHnvlcfZ
Kqpb65iqk/3zh7KK0H6yOGdhsrx9CkaUfQuCREuqZJnGUVeOBeqnvU13aX5m
vMLtBwDuTk5cN7sw43/3UURC7apiJQNbsXUR5PGo5F/xXz2+BlYO+RUN4I9G
v89FEsq/k4VnEq3bmnyKDSngBYcVDDOOooJE8wt5m9a9tF9GG7e6KkfwUyEA
J4kntLwVgeaTDK1mud6gz1VAWMantulcOcSLzQPB2/p7tYw6o/vsOWFOjQ//
pxadoy0XGDZcEsmHoRoOlzCxeb64Fr6lcb3S70Qa5sslzVe8pPO8RdOMnAyC
O30d1YUwLzVVUT+7Of1smMxl4Iq9aPZqSk5QO6zmuS/+ziHsYJMtnKIKyoHR
N03iNOiQP0i4C2PFIBRBXTmTPu5VIa0Z1OUekWPct6vTCAVELtx3bszMpH/S
2lUNgqAJ9IgpMm10ZqEhUrDZQbfHRiiUJQksJuOtQ7RuUa4krO6/bP4VHw3r
uHAcF4eR79qK4koHTvH8IPbh+A+OaU51FbBxss7U73L1cxxUtX5WXc/KOFPa
ZvVoOGMMI+NNdK6aRB8b6LyUYynV3yCQ5+axwqU62y8y27Vsw398eZMQpBLR
kAb3gTH20IxKGx9CgzIUVeZ8d3CurDWQZ2gtdnjhmsh1/ryawZRrRpijc7AE
Iej9LNTkR4SawUy4d989kBnPgpb81p558h5zFDwRsJx6g2jEsCQO30EEwZx2
ZaOylbNIueITMRaBI0jf/7f/Or0zH7j6ve/jWz1f/zXwiK3XVBSWTlbXPk1q
qZi3GcNOuVzNwtZtLJoAdbE1LMJ9p4BuRdpPSzqwpetXaR5bXdPfYum6R3Y3
OJhFTmED58/ErXqvtiJk1cG7NK/X3fTuJQsIizemz1+9AJv6HUyYm6Eh9s0f
Gejh6ZpoHVakOHrfEaEXnZbMFfHoXAamznQK4dQfaFxDe/KcweaBJ/2HvNsL
BxzFmelcrQVSEx15e+SPCurFtHFE1JMVrWOaAHhn9ZF3QqLqLai3sLSq4xOV
ngKTL8dqgV+kKREUYhYsKSjAOTKPJ/LbgqI3FiiJJpq3fF9gsr4mBkGlvLjj
fhiBVmOgbSTUKn20Q/SQPurxrvLFzLaznRRdCbp5pLrHHAwW0HPKiZxNZVn/
1Fdhl4/lEDDhL2yD7F4VndUE8d9wPjZVAkl1n8zX5Fo7AOFNZRsiI7ZMANXC
HWf2Dsr18rBDbRzFkzLTiZXPAAUiTOnMoOJN4KRblPQXOKr4OyuM/AIBDB+A
sX6frBNARen2GBBNOcMJvFyuL5E+zWYAsMRNh+KY7+JVe2mRNNsCBAsAIuEA
fW0SkV7sCljYoGEE3BNCfUCzolbHv/zgH095My6fmM+ZrdN7UxicRioPx+SU
TA7u94jSdjTtKDlQ21x4aEmdiNmoSM21yF4bI5AjOU5etK3BrSAhoGmWUVYZ
3YOemZQn91z+UERD5fVRW3LY6FBE2LLv5kGzt0JAZKUPlFLsGRDanHX7Mds/
yzaaX5WmRc3oOGbUtQUggPqr8gjzjbHmEX9FFQBw9XGjZC7HsaT1kluGJWuG
sszyNc8oKQBR98STlhvnyYHZN7ojqpFu/12+wVcxn35dACUs1tado/vLMv1u
k/5tLWL4pN+ex5+aRdJiqfBpdr6DPuTff1CAvChJssXTeHWgwE7f8avME+9B
tDMXcNCwvX8zk3KFKIcPC1/PhNWeFMsbCcMf00OcAvLiOg3GuVKKUj5IefNG
cOWKAYRZTnWIVjeyfCNDnywQiIXWS/ptRu1gdqHLhbfkakYyVyNb9nwWOb54
IQHcP4UW9xBwDjayttDE2AqlbfJWtO13VrUpQ6q2hAbLGfxsF+QSkKP6ASpS
sMobTipZelYFxNUJEADGQ6uOb8U4AHtJmlUix4Ho2q7xGU2jGvJ/pjnuCQZp
2K/VFM6gPkn7nn44Gld/AuRFKzfjoOY54DItbfvekfLQ4SJQAFpeWXbP0y0C
H6r0rJjFPvWAs4Ud1fNk7xIulc51D8pDR7B+Nhp9F08fHOoRqnTplGqV4fxT
pYtE2Z6EJE4QL7dBD5LRlsAuNdfdBmNILtML6i6EMgk7sa0QifC5a8hQtqv+
9lTJG0lgpKKWQs8I6kd2q+R8BqHNZpdyCPJyAmmyJII1gX5VX7kanPFPPJ3o
Q6YWoBJEHtThV1lE3jpP74Ga6InVFr4LlbcNmlQfx3/nuN6ggoTQYKQvuFdf
kXv4v0gyHIxXBfiXnSDXsmLtrHUpQYH2IXR0hwDw1qnRumyf7EmTAaDLKqnq
Xavpucvp3aFWM7xq0JjhejXMwbCYGzjYwYaL5M7nEqEJosJ7st0E1dD4kp2g
GbmtJiem/dp9jA76rGTN+AZz9c8eih5fx4iYDdVR9go8ocQwxMIViiTblhBu
eAsUeIw/cj+yu7YULC6Hq/dgQjCwrZKHpZFxLjwKS5/vpL9i3xS503RiMvBq
gcH057KBh7AVKEMW9QcM5nZ1AYCo3ctLBKMDb2IcJs1UyJIFgG1jZOyoE43C
IoXPntnYImIIhIhn9J1klErbgRQP+CcohuKwa7rb/5CxSXdrQn0nBvqICBcV
jBqsZrfqvT3bDfAFldMezwuT9PUiNujkd/zVkSS7OhNmNm2xdMJO7qDp06Iu
6aqtWCGb2BoTA9uJ4jECU5hyFPiE5NfMLt3QpG0h+uKERYuwKGyfzN0Cxd72
0QIrUkcEANg7H8SwP3rSNh+i7MZtfNr+VO9cS7b5PL2wowMGCwux37CjDp/t
bsmHBrjfBEbuniVug8l0R86HKOFkIc6a3DXniTrfXvQA/vu8BhIMBFa25pL0
psQN3APAYh15ivVPVumwre44bc68ShXp2UGtwpOcFs7cBOmP92hjUW4hoj6/
fiqti/f5gvbzY/sYdO6PH6qqUrbZqNKFldRt5jR57ON+p0XwrJbLzKPeb/im
sp3YzEdkLJdlcwShlpPQwelR8/8noGBD391E3FuG4r6YNhPyJ1TfGSRB6E9I
nZ98iP9iiLhMdXftjwp6uri9DCTtx/vlWVoubgmL2e+Q16PNmdjuwzt2v2lO
XsQk1BjAzB7wLiMHavpNoyyHzxbBbzDm87K1vXJbOLji4hhwOQuOmyZ8nd5R
iEMaE33CBDPAlzlogsBa/3y+ge17gCx3snpv/9pGahmrmYOUW1SmWtII2Qtk
0vm8WaXBpYIUujEJxRhWrClZgK6ZX0FGLfksoHZMcuOvdQkF3z9MUdgowRq5
7qnmKRnyYeIBnKOfUmVeJOx1V5wZBPMzD1Dv1BuTbg+1tDexJC2N/VBORtPA
covY34gwVg1uFLKYRk1samb/EYKzuG7Pg0ntPc1/P/v3uOdaSDqJ5mDJu8Gb
Z6IOWlexGruPzJl/rdOluCbw8LrFZ2w2iBRX6AhxvHdsJb/rguhQc67E9VAF
ND9AXOrtSUAjGnWPu9ZborHYf98Ml3t2b51ROxr8/m+E6LrS6MRuKB9Gae9B
G6hLsl0vF1wSbD+6X9KXT2i1GoS6tDzDqB7cNKnruqTpRJtwJbtQoq+VU7tb
OvLqL2sZLizDlWbpujqVBmGL9CgIok+euKynpvCbUUYbdBZBa7CqWen/GJaO
Bj0XmWq5MQDeCrRBgaINIhkoYTYpSFhv3aZHY469gViMjYffLLwE5J7OEcY3
uFitUqQCKOJ8vO6Uf9E6g/7L3Hb1Klmqs3jO9ldCCNWHfgntime/Gt3GBJ7L
zmjydX9UoCDIaWBKPZXCyXx3O4NscPbgLzdhVZ02AtspTb12js+0DSLCmSZC
aexZGch1xzDuxXsL71OLb4+KGaXPiRyQj2CAfQlB6EeqQQDdzBHq7X++elOO
sFlU/aZ6geMaj2YWblooSCgOXdpV0r7iqbdG3RcWiJfs2ss7njJQX8XqOPhF
0W/xQPcxzQ+H9oiBjJ6cYDXEjGPvrvZx0qMq9Vqxs7jzicR3tMToGv5vobmo
XmfcEYD7adsKTLAhp/LvSyXBvhxtLSKS6AtggWM1Ik6+/GbKfqD0vmffPZh9
JAs95X4bR2YiBBrETxKjKQGuG8nG0Yta4/KH+UStJ3f5MNPrBRCvOEOCeKkN
bIAij6HKvXkikR0LO85YXCCPZYBWF781DEmCfbTqJHOBmDHmgnGa1i6HJMAf
drHFWALFzBMqFcMr3UAnnR72kvsECNINzxgzv5mwPjMvVaawp82igGX0QH6N
o1MJHJmAKExjAAeh2TYzA3sIWuDGsWLIf2DAqCw0b1r3DphvaTYaO/rdPqW8
WTdTOI9A3uU1klSBLXxCgw5VMDlVN1Jyby5lg2N1KxVmx2ncfzhXmSbUWfnw
LPAaRCtAxXGRN3fsd5TNB7x9qz4dpMb+805UIhdY5KaZ/VQeQVLCD7BW/Jbk
HDhYG/gwMVR5dQ1by7ZkgxLhHcRMUxoGMcye2VUngmUQyWAlJTBRj8fUjvgc
u/WrlSCWPmuxfwrz7gKKaT9yZ9BEwzpRVAPGudIUN1ljSxzgSPlbewEENegs
6GtiXLYfm7IoyNrl7niJ7xfwb5YiQE4ULJHaTOYfgTYcdQpn7k8cRBZrDWAS
JijPCMAPEM41M8qBpAL7c6D5dbOIKkiNIdRS2zfMha1Rjg7Qmln+U49aG0fR
4ytnXFxUerbUkZ2OG2nh0efaBb3i4T/E1aAot8yVcJOgWhhc25TpxLtK8HEL
ukc2xZRWXNsrIkyl0r3TsWCGfBxivvroa6XavJJ2lZZQR6A0cIRA1P3t9txQ
q9252GA8JlMiwAMB5upn2D3g9E0Yys66ymWDWNSLR/HTuRwXMZrCZFC9OUu2
YmFASsrCoqFyjxX+6nqb+NL2JdFzmi3HqHD28XmnaMo+k0RR4kHPCHkdPBfI
D4zXetn4dhbOsHjaaBSCQePDPs7f3HhRLaSGyJe8xd7xnhqjIQm/8m2I/9ui
nexQAyLvEmCTiEFCk/cB/mr2MFXgr3BGIH1UOf94LYYvasyKcgz4xLA/wDU2
2z/0vlZdL3MgcZPdjEvV2P2u391zyj93y371hTDfn9VL8nNao4vEVVliQWRq
M1yDfEYnaOkPncC7Sr8QZVNzRzl/NeeoTuXcDXBGlLaL4RqOPsPQzhWOBCOY
zBgtpteQ/ymWcNALH/EpqAe6wRFoxakcZSziGL1qEnLsE6q6AUX8+wJQp53Q
ZF+Vpi9GScRk+hxBslBT0Prs0ZoS2/EYiQ3d6QU/lRWFIAk/sVdwNzb2B8pC
bE24DK7KaiJyOBbTVThrTUYcIMp3hIjvMdN6s1qr61XMzhe8BCjP2grcUtur
CwLWqqRwZG3NzuYiKXIAWJFskkbUw34434Uf+IDmZQIBCOXyWftxIzVtIB1f
yfJ6x5BhBbyNf2F+Ui4ofnVFiLrGx4wMXBcACsguPmWwkM9fd0f5AF3XA/nx
fIF9MEJePFtDTjv2caWmuPoX0Dk7EnRWTzb04t7I2rNzVUbOKgMuu8BBf5xm
TtuxQX1PE3qusAhn+e2oBNs4dfKs4aDHkeAxNKywdmlIwOyaPFOL7Jc1Us0c
wXqwqralJxmK/MopOJy2DjGr9+zLKo8aqDTOptwQQRtR4FlpRgVaQKEQ/v2t
IIPf/WJomm3Zxi6iVOGNCDaBTkUprUDF2K5xcTxm+EcI032HRrMaKstoFHZD
90jvDNyPETrfwWrxTlbXJm1EgKu3mL/Vt0g92Lc2uRAizI/FukAmLRWrAilm
RCqMv+DTB6QeNPU20D8dHJsCf89Oya2USS11CUej0Zbu8/OFgWXLkCQmoIKA
MrhrNbjHLTwgP/fa3l50CDJGYigU5tM8XYiXJl/NtKmg27HJIGr3DWlj5nFI
zxmgtgos3Cfwf6HeguJC1J9butYJ+BdAG4o8KnkrPa8wzN1KgsmNB4pSIKqi
UYy43DP9G936VhMTWy6aTGReS/4cE4Lf40q8fFCY07D4lIzCsQXHOLCifKQV
ScmMfP1bP6llgS6yVwe5gY6lr1+WknyoBj+fa+qUZ8tGXzCn0MKNfGaUzckm
aQrnnlHAmyj0sE6wNejGitLUq+8ezuaS4NSJ8SAWBjy7QljUafSre89f1Jym
eIqr09g5IBR8bM/L2F8t3MwIzJ1pu9rUdWrr9L+TEbB7YvXdQTWZzQ5P1zTb
qhIxdu3UoKyiAvbXcpD6iP3ASk3sH/ptw+6nZ9A4lZO8HL1gi4/uldy7u67t
B/B6fi1FQmbQmjhnF6nAfXhl3TRtgi3ZKPph4cdBeOYmImo0S5UtoJxvpXBg
+QNV6VqBemhbMeQB00nPWrWCSYrrgbya6sJlBbaB1fu4dmquY6LJY61hbRZU
bAhoKnAr4cRLs7Gj59GUbxoiJzOoTGA4K76MjPdetSx0fhJvc1/g1QZvp7ol
s4cSZqcpgd7SRmn3awYAdFr4TRR6cRVbfG3DSH2EfqU5xQJC/ARUuaSCAljI
gNyQAleJ5RZzj88mDUUQuRQ1QmKCOcC7Nhk8QDCrSsj28o1uNx/+/1UAZzV+
Fkj54GCeSC1cAUcJyyxJYodGyKTfhTF0O6RZGigmTlHTp4O9bFdmhPxOjZxn
cgqgsZDkcC5zVMIRPzYCzHOEogvbN566NKSrvDxoDXLYwUxhXuUYmYSrz35a
mY2JQfpOQ7vuLTHqtgylmO4Vf0LQKR604lHYuxqdWLT3zm9mU9YynJWdVhdM
O/R3Uk5O14GBYkZOg7akmESOruTfTeqyxdXgyqVZx30f/yehjl9DSdvd9UGz
ui70uHOIkvFN4EeME+rLejWVKs6a/efgvt8Cy3hK2iUfRKGugcvG9Rcn04rQ
oX8IfoEcY/NevSC0cXLcvRScVexWLtPzIDzYY9Is7R135jCiwlA8zDG0UVSX
FwlLehqi+Kn6kLCdVYHen9hsaRg2IBxr1VzOzk/ySKm2UUo0mHDPsKoLXluX
W/BHkmUMI28WRfWti6G9KOZtQARmcKZD+R+5MzxuonYw9JUoK4QgVqi4b/qh
uvQEpZwvHrkydJGBeG0a9MdZN85fA2RE+juZUm177F/dDiqstIBt/5KxulPR
+ADEv7SIn3isXW6707WPSfifGTphuGhRlqP1wfCqtZdgpzjtnZ0RqSJaUbUR
zWO2qXbaiPfaCMJakxysR2gzT9xlv2w7s3c2dcLIbqjeF/i71+csYSU7LwkP
IM7AJdrAP7JTKUcFwBa3+fhmqy9O1w7OVZ+gxKO1WE4Jg77xpAcgNbBxgjFl
NgFwIp7MWMUNmkcKs2HSXMyy0HdYGAAgUXmc0bM2Del/K52hNXLRw1Rz6rSJ
/XmZy+j49xfTiy5CEyLSstWn23TTiKfUPB3zf1i74tx3M6wFh37JrmJIm8em
13fITr9Umt3m7cZBg+WRTtxMWUwPGEQW5DMsA2Xslnx9qhtltNwUfGCMomSI
rvHF/xbGeobjGcUkCdeW5sbZIwjnT8xLBxSN3Pt3RIH7N/ei9OKw9tTH9Sb8
ihiB+p9rYkan8t3SuwGzYUYuFOBJnic4wLpEgdxJeDNyeTMjMix9IqEdGHxo
KVr95+3tQlo9xBRIu/tUpsuq70ueOvoppxyBNcRPJ22uH6lkFUgRNjOWTIIR
ado4rmns93wP6k0fk/2wkBFBiOA2jBvacWGzS1+CfeOhSUe+nrOghjeHPOoM
wXH+iX35wRK547svPYJzNpHNz5YAT749f1zz7YpoJM7Jg9Fc7sX7lwZxa3zb
aL7iJls/Aw+VCqPQRGS5s0dW9xp0VXck6DFwsxKdpnHglpikTHRaCNk5Mf6X
v+mUa1rLfBNv1kdiiMqasnGUS6YYxh77QqT5l3I/NVz2SwMnttomPqWixer+
mpMOBTeRb+1lOuPVBBoiwPsQ+cGVLDIlds5RGmnJBwN3W2/0yPoNTyShN4wg
YV3cOjdeEJLUkJoQIA7A7xRHl2PzbMM1okcg4if3WqCfru4nrs6P2pGbCScf
4pZ3/Bo2KXLcTQFGkz78UudRs4g2oZsUaYe6UDWGuxarIGYs7FC2S3W92CVS
gYhWlEt+p7dN5reKQ0HbFqPwHNCx3qh6u5zXKYTr2hRcWJ8at861yZTyBmkL
+kigkMEgFumSEixXamIEJPuxXamm5uzsDMXhoVsMARP77oZThQbhA5ja/Gwu
sXhgzNtSy/gVcxp89v2ZK4HVHVBbHHYFQalrwpdT0l61GhwXCOkq4aFiyELo
H05KMs2vniswLLVh9zhqDHxuqJVL9QyOhsrDLWx6DX/fU0+msqgjh7sendeq
MdhR/zDiIja3RK0/z8DhuWUTJXL2Yufj6MKGB7CXFdi2dFtZ1hBi1Wk7Shzs
UmVvB51cID/TP1LQBL5wCQLPmTMCNrHktJ8lNTn09gwxToK5uQnzZXJG6UVv
atXv0LRiGAmNrk+FQxVlyL1FYS7xuWVqxcf36GKyUbbjQcmFwFZabZ98sOAv
VECDMu2nvUuekXPsa3BZCn6S7pKnpw9yA9pROTIEHWE1Xhp1eAdQ+p/zrZ8P
rjrCF+YtxV+C3TjneeNj60u2MFg8MNwTp6WLzEjXrd78Qvb31IWA1DT11jbC
JYhB2sSjMjXr610YirZ8ZJEHrDpXD02YlDpxox7moa4jeJDGAV+idrgsc6Vj
8/ejWixwjueKaNA/lsd98y2vQ1n4FhPH/P7V3KKIIF3Ye8MKpbK1diE7i0nW
pJCE1IfbQHulaAbjAX9rmujIr6ORIgL/gtyJggLxRfHJ4avqso0XoH6+J++u
WmcOWjhv70AlOiYtpiG4YWt9IUw3JkO4D9Pp2LIsDebrPEDwZnwHoKGXA3Gq
zEfHaeLHg7FOKwELrq1YZWYc3tcz8dAaIcpRECTp6R2YLxYIbMGBBMR+HlUC
i/8BDRwMMiaXu8xXxdPEoDqq6ed+eRGofKn7/lEdNdY/I91C+HhrrKnpCSOa
T4Z4Y4bA5eEl69XUgnOVk60uo7D3zI6h/PxEaBkVNAnx+H0uS6pFPhZr7LaP
VxErf9uMCU1dqzbkViD/e9+eLvcDHXR9FFrUhC0Vx8OQqIPHhb3PA+/vY9qu
wYjFEu4EPNwXlitFWKyYGNmo3HMOzKcXuSypecG+AgOO9R0PC/TqqB1g2TG+
ODtOSlWFIYTPdPCQLNKp4kOMn2WVuU0KZ2TWuFIA7WvYw9/YLKFlSo4ryN+A
pjAU7kH4j6pkQ+are2rH86NbN8BycE5BL3/8Cq1/BH78yRYHz6pXcJIF3p27
MGERrVIgurST+0Iclo5cz3j4g7dv/rR7BTUJ1i8Ycr9gLSxqENlGHX/k52pm
94mlx+BGblixsCibVSOdWrsBISnMugBDZmFdbosUy0UOTxU6uHAXFEA76HL4
tWhWNVAtLcTSeSHE6/CuEX9dGcmy74ORfwrx63tOSKKtT2P/pvcsV9bSLQfD
sdhlX1UZ/BBWgTk/cMC8vOgDZcXUEsgja2M2X0ddx5/EbwMRLcPSTVXbUm7B
Y5jYSlQaZAtU4Dz7PXOgEc7DXqSWuL9OpaiLVR0bxqyAfiwTmsw2I1kfPWOd
1ddb7JFxL+KgwE2hb8bEpBvteP3TfkI8iHa9GZf+cqbverwBiFFVD5YcIyvf
MQRTN3yK2zV4uMdEOW1rkk5+M3iQNs9MzO/4LoiQ4nK3WIUuT+XVZZNn20iW
6zfh6tS17bWwOHqehVwtLbeC2wajPNmA4hVYk0uODn2TujanRWIx0b34H4En
Ab4N08g/2ylLfPwAINz9B2jukRXgT7yztQ5ibpBPm5JQ0DC2AEu5IGSWjaCG
jVi1UOExLiLW2PIxO6Nv4AqNaoC727D6QRCeDupCVzcne4KGLOKcGCmArDox
dgtdAGl1UpGfPRJrp61AfNW/swfp+mlvzKLOzUV3he3tVnw7Se+yJBonqCwp
VSCPnIPC6NRHtK+g0F+tcCFZKrkK26GTqLE3qm20XqlAnYQY2563uGhafv9c
46vLtXBzTIDunyqj7iu2CUH6oGasft1uihOKCZTmFySM9KAG4EIxVU3WkT7g
xVPI4M4Rg3r687UNetJByBMnJtEIptyq9y/b+tRRDOiUUeom0AsG/rY9qc4K
xMP5aPV3RWddd0upcflqf8pzneJAprnNgTv/j78sLqGufbQvRx3BiUH9Ec1x
hSQOM6V1Q5aWApgwW5SfK8Z3IF0jWw9VPRtlNMwt9RbG5TIMlAvqdHFw7/Nd
rRmj8Har5T20Y6UnXRHwMMrkpdU9P1WYwGsxTNPaWEX1F0UsC/+ayV8L+dUB
coM4d4sQfWV16pZKNL92oV3uFgbLvdL9+xRk9/LC6gh6fOdYQdopLdCkEciI
RnL5BF5SRWwiftqh6lKsFesMp8KiJh5PP0OOJ4uuCbvG5l2uoNgBMLOl7s3Q
6FyU+KrVZj2h+EisOQg8saqErudgsVTEqXsoqmcuIy0+ccCcNWg71yYAGFUB
IKz3JDPtzWb9q11bEO71mGIqjnmKB7RTWadb9HQMtsoDizhzTS311sLYL+me
eq7xV2je3lMnPxnMrxDmuHwWG1BtvAh3lCJKrQ53Z+tOkuOhLqXOC3GJvUfc
LSZY2VZLkUZIY8VNJdUhNBAR6RDiaV//yaP/OJbWYfPttAdtaeFYBZUcjVFG
8TWDKvv9uXzCfcItIF1oLlyyKHkuCZn4vQJJ2dwc/2PX9+y4sss2nsaw3GMd
6AQQwn2ybQhTTaTkMmW6t3ic5mCamk+ZVkAdUrULUEwQaVgv1QQGPC2bqvdi
fFi690qPOL+Hf6i3qq88DLPAki/vBa8J7c7xVYT/Fbff4Mnt6B9vttcyVhsq
di8aaQNUNbpbmrmNdbVn2JegwEFQ6Yi9otHvWgQvnQK9iVRZt67nSmQynzew
BajpdAN7Vitg9ZlklhFJYRLi1PuFxrSMCroASDdOnjdngtZeimoSiY8dzL+I
mlvEjYwiw4ak2Aqdwb2HaQrmSyhID2HbZa5zP7Kge9E50b9uh5hMnnKPv1cb
w5eGAdIZqwYjYqna86ApLJLKpYGqibA97+BC9BhVoNhTGiOsO58NzSS1vYfZ
WX2NzRD9BrmNfhGULfyvtY5O4DdxW0DQpWdWgIESm13P5Ef6pWxTWUXmNvao
+oui0/CZ3HBqQmWPi/tAHbBmlzJoodwaIUMMGVX2DU+LsLxZ1xdAtK/tEkM6
FDuhxs7aP485J0VnqRimdU7JlTykHv3XXwp/LQvvQN9MVcbo8MCAyOeBBmXW
oYuM+TZ6HhMELLSvWFcQ+Mu+kZrSFIRjcwX36Fc5Kd/HksEhAHd1VmY6BrPK
6fmyOXPpJdBI0rmNXtH8dSA7avEkBhnqU2VrCPP+dAiw3Gn2L/2bSPdZPh5C
JvJF0MxNP3cuO9BuTQvz1NDme6VGnX6rtd0rFy5Ax25J5Lxc2cT9gEvZkL+X
VTlQUiUwQEyOG7p5SS24dQVSrP6CBj5gMxfrE9jmd19PdY2qh3ZHE0DCCJh1
MClvHKM2Y/u22R54FIBoaOS5YS7LzBYQzdJXpFb9Qk0cQZ3K2ptnxmPrmqbE
asMGe68nJwaHFofvGd4MzNdAgMFWaLssz3hwnBrmvlNWc6gp+Yv2+vvPPONT
qvPbjCmGwRjn8dKlx3A9emdlwn41lpqi8lazDX6VsCjdhvi/yYbgCnxxNtvP
CvmHdeLNWGgYLr8uWEzoWFrhOEBDHhxoHidRB9fJZpVfPQLa5eegiJSxVgtS
uH2eFEbmmGaO/iKHrx2nQ5Us9HzTmb8/MS9gtTa/xPDFpshwCLtMo2o18poO
JLNUtGNYzxw3bpNJVKTP5u7iaq6VwzXx9kBD5iQO2CwJTToMWSPpH+iXwvP9
GjDylL46dwwpjGji29ceuRoPA7/zFFI9iSH2ehYQGlC9DISXe8Y6qXVVoUWY
JIj37hWrG3RfGfoX6Q7sW/Ry0n4jFmXRalKJ5Ue5lDoFxmUTz82Ku4ACO9Si
vP08pHFpxqrFbLeo+RZ/LUJQRFcsk/c6vRBjte/jLzyXyPouvrlON34AY7hp
lVgfzAe6j6Qoz/MtDUTMKTYGUYOP5RTEYy2jOzf9w40s+D+uHNn3fjQ0uf4N
wat0mFBbLd0WVgzke0VjjXgDQbZuFz7T8ShPx9ZMsWBExlMeA/rjPGN8oFsG
rL9zIXraMjlDUHFRFC0fOelE2R+4Kq5KgOcBR4NELQLcsWy6PQjIE4RMuluo
+HS1dFTRcH02KEQS2jsgD6LSu7tuQdY19Y6yeOvCqmyg6nNWhooAINvH9wRS
ZA+5L5vgUYTsU3eqtuFQJx8KDBcKsH8LGbx0xn0w+IoR7UiM2vpeP3O6iTjY
ng3FHkRUD4PRvwrxfFnmNaTMxN9nH/Dr+f0JwxUXtGP0OEsdksJ9RWJqgFe6
EytcZsNWSBEfGqq69Y0DS9doK1pXkcrNIPgCbUpe3FjV7B/1aydl8AFRHe/E
0qvQGUqq+33VIKIM6LgKPwypVodd0d3bPILyewesC5dhFQZiR9Mz5H05ViKi
vbMMWYmznQ7LXtC/moLE2WXesKXaNvp1ZFa4fIi8Bslq4R2yGEKktVvKPQJN
z2+AJchUz527M7KauZVdfR2aUakRRej/9/uQEGhX2tYKXsiCfxMiFoWZ+piD
V6KFx2sRSnDASjHrzs/rilwKk7S+4WyCwDAR8Ql7idHxmvqkVwInc/4yPvT8
vRJrP035q2FG+D8VlRzlIjsCb4lXfvdViXYHPyoc99BJUpj1GFphcsX6lNd4
BCF1tdtAytzZ7zXClcsd43T1ybSeRbVEcr8TaeLsh2NQAR9avBj1J1REsv7f
cQLY0xCzdgD+fpeaVsjMnKgwIK/dF6FpJTki9cSITu5+96JqeO7TV5APJKVw
LN+lF4MmjWHRASUuflwkIUWaqE1BE96KPiGIzJ46kourjdaNMw7LohTg51S5
a/sFghQpObCMivcnMa6JS9yV7jm6VDlUplZsFZd//uZj00B6bX0K0+1ug+Ms
RWfWqP93xlNj63k5R4jbt5T9Vzz+znsD3BTKC43HZmr+/kubmDjPNqWeS2gg
i+wfMXYVr2OdWDA9wjNTKUm1IqcQUoV89LDPbNC3Tw/fdvuKaUJUSQuLkIL/
182XdzdrlxQkX1e1CNlYd+woyE7zsHQnHylIZ5OS395sZbgtV0CaMokdRlbk
tso8a15EPVlf3cAEQv7nf5HhowJpi1Lm6knliToftMmXqmFctsjwbarVdd5Q
kTrxN2ZdBT87sXxgBrkYgBWYLF6+BZf7vO/TAQFz590ksmrH8Kw8Q6MUxx4V
H3P/wumvaakpLxng7mgrFmJK6m0y94Jxq6aXx6awfXWvfJc+r4bIRXLkwyV5
hP0sBQdFau14jqbf+iyCy6BnBX8EviPYPgjej4jwjXMIj0mps1fupgCixPOQ
AduQGBnCKi7uG4U/w8y0mrxEpgwCT/nhDOrOu8gRoLbz7K1pXw/5zRWqh8jb
ObyWt9NeDqbWDOapuXxsEc5hUBQm/lnhxpWjJBKsfxovLKAE1WwLd4KWj6rQ
Yro1DERmShp5nFk52kYfuL/5BHVOHfvzCVoVooUuGiXZMCOsLv0ME2RBdm/c
dTxHzXHLb+FYMnSNy5xugOQnVhe3q6q3XrU20wdTeYd7X5rFBIdUZwkTRhSY
HpjYLSvkgnHIfFCdrwe2MaGebiTUL+6EYEekCVScAfFLora/JnXuGNlwxJln
84ce+f+4EPZwhNwnUmm93RkNzjCU8JqBOLXzh3aRjBMmH8oGAAf3Yl0vbtAm
hu4hochq1DnDpfyPnBPWGB/m2TkrivX3hx5I6ujJk/PXs/dDLUI0T1r877zT
dbaMKM+Krj7wMPVvJh7S0OaaHb9OyFw2ifBy/uHL3jtZd57+QvJH+yXC3mhw
5/CeJFzXccHr4F84dKfeMG9qkk9HtEL+AU1UHX3jQvBgKaUGSdpPWpwuKD4X
QoJP8Cxl2j95wJE64P8YBzrjQh2VGDGuOHHByp5FKig9EmTL+gQP2UmDv/PJ
UPKwy3VEU0Bld75qn6rB4OkqDWHa26Vpns+jwL65CamsaJeDnx2F0yHSAgH0
BkMcDGCbztnxow8x3Eb47jWnH64a3FIjqGxcjZuJ8ltRmnTpMk6rtl9guTth
eEi7uRyvdgVW+dNO2tMlRCT4lPoMj+q8P4dnP3uWEsHMVbEu6qV7gza/eUT7
lZhO12KgneJeWDHN8ptGY7BL1tM1cdiU28mYiKxhZCei/YgQmt3kEpFV9tyX
kUgo6Re0jqRd+IF6EtaYGnqGpTpoCEOP0Uxy9mAJBDyAbK0rwqFFzzhKAUgt
i/75GzDW9v4gEHOXBk2gqjvrXfQK9tRoEPn6zlwEZjUpnLFii9Q3XMsbNfge
agjW9eh2/JKjKyLleARf++iyjDdVSEWIps8Yg1lOaV3pc2h4ICzFVeE87Wrv
N9NlpF0TuMHb7zxj31UpwmkY7gF4KbhGQU5fsiyTwNu+GD139zKy0Hc+I8Bd
NkPYhqn9llWb7hAyi1buxQ+ZMq6qF8IQ++Pzcs45fBuwivdDbbpwB4MkESlB
mSmgXreGjqOxhPD5lDRyKvCAtAi7O07NcPPjsG2D2XEVbbtN9y8Fn5/t01H1
CPhcQSlnjCAe21BHi+wo2KO22ERxVxLoFB1z/lHzFbtCzWYKi4CgdH0vxybt
xc+Aqopvgg88/7AuC/kir9frWCDaNTFp1m4fzVRUo3SifORIClZEppCI27Sb
8NYOxZfAlx5bgfNeR5LQjEVa+uNi1yqHCyLztZUBPk42oefKp6f/Z5ZoWD4G
MpXmdo4DX0HW36nTbcWQ9Ks4EXLk3Jjt6fDjzVl/AAHRFAUp4QcVGAiBt7Kt
s1Ocmtbn9t3bbSSjWM0d7x3Z4Bpk2LUi/KBtvbbpyve9iE4hB62/pKsdX5uw
JeAKTAXYzL047uDamKTY7zfDCZCuC/+qROvYR9YWVDyXrUPB7eZl6G0I/TWL
zDj7XV+jVQ4nwp0CABHOhmVKKd6A4ZNlzFT77APb9SmbLs7XRlQjxkyG99Kk
Xq0DLbGWsNc2Jt705Uv7VAftiAeeT5epjlp8y/FsuTB8/qtKV50F3SJCmNu9
sytH5ap2lhgOH/PVUkpSosgnH3BwMIR2/J+sGngsi8xQlMckGr9vcEvO7MpF
+QWU8qTLckVMdAaeh9sixI4Sd7YXFChXM7pCzcgjX8pLTmk+RdnlLQDVn5Tk
/Z4oiC5oIs/Pa+huoVX2wqeohyI7egKxJ16YyOk3RWpY68Oo0pNdOlhpy+3G
101aZK+KBONcvgvt7oWf32rvdeVr6dFtMbB9wsVyEMlcf7XDVCkAlhUJjIQA
J0LEmtu0h89N5PwwhAvP29AOWD8ImeVvRoRf3H4Uiz1ZQ0kPjXlYhZHqlkSC
RLRPJor3+keKIkmS4tVj+vzA4MfWYykFoRqgSVPfYYmoLuLsqJNx2ozc1NpT
VFkRAJygvD5eX2tY6kFh2IJLA2afjCgvnfEz1gz948Q5IiVDwsF1C2UX4udM
RwuPd6wV5iFWPwQg7g//sVCoSyOir/6lM3TFMs9bjbGuINLD9Mf1dY24p74u
KcRoNICCJSopb76TYPvWecRfuMVGYX0Qqyfw+ZTYOOwjRPYieyaBQkJs/PRr
KgcPrAeqAknz4H+t/aVF1md3U9Osc79ThPZfCxfJsfbfuk7mEU0yzvekL9W0
Cq4Yvwqg8r16XSp7zECKf4nNfNB9IpssURPsCk5Hk5JiOu/AniSejF0NDQ2b
7uWr9Y0OQa5I6PWi4n2rblHLbQjbj/qztBxy9lBQS1ay+j03u+FY3fiCoCLA
2I4KWf+nLxu8EDbMH8zatnC6E1Dgi0F+po7/PFXVrEmUAS1eEWJCXKZEd8C2
zC5YDSwhj0U1BlXSZ0LBChWASjcB6CLFtpH3P9yZU0MAoUMXTEv7hRiu4n1v
wG0mXdB5HGDfF0WM1N3Ckg9h1ekurl4hFWJiQq+SajAgW4EftdzcL0EicR63
oCxKHRIYL6cTscX09nH+db0xvjcq2vE6vwcubf71WAkusuPGMRrj2RkA85bw
SXM00Oetaz8Ydw1b5ulM+f2rj4hMtnehcXjmlXl4jtve0gW1x0utwXMyBRR5
v0cdIXAb8X5DKI5MmUF7LpOT5MdTde0MzVVDn4M7gfWr2+8J2IsqCMS4Jf/r
JfiQ0Hi4Y04t2wqr5HicfjBgzywo87LNiRYSnx96cSV2ntyM0RqGyz4fPy/T
bVKabCKNMGZH40tENRqnikMaFjsiq2/pZ1h8vA9KbMgBbU9ra2/4EzPt2/do
sJWK9z4wrWQBGjnlz0WxRG8HfHKP78K8X2Hf0cLdTKwsgm8NCsOPiojRHc2O
w7f5Qr0louwO/sZXIgzwSFTVXLCxiCleQrVWLcGJnKlQUVQw0vD1xJo+Q2N5
TVHx+iNm+vUvYV2JIW/NVJ5iadVQNE51IQUsZK9+Mj4yaYD2dcTqSXYfzlhA
r/AKg5EHuG1o8DDhDX4nYKDRyT+cS798sV8P/aO+JcHuUSAbUoeaT71yNT1L
uByMg2uwfj8EIHuWWoVjM2AlZXxmDl54du47kc62v2YgewXI1KxSCq19pMTK
kUzDf+kTSBce9T2okLdYmq2A1e8WDWlQYYpAtJx7ePcND5VBLCZuFAYv9dKt
yejAtKNvkz/OjF1Am3ZBZNC3yO31j/JYYoAha+J2nIFVt2yrpSKKIUL4I4yU
fssayUmUqZTbLxgsznl/emITqEHYC7pg9MXbdWm/XW7z+rdiTKMibYito3IW
OJHmiNVxueA/tYvmpm35aNTcro/sPvEhBqApzpjkEojiHdtT1Jcslf5U4EA1
20mQKFoBSLbD9vjnyjPXri6gj8CD9SPtj/TJqtCwcWBgvyoHA3gO8yR1c7Yt
uN+1vAYREmuLfN4jyIqKzUKzgkpqyt9oZR6uMKkV3QmdDXqzSGvihOGh8ljf
hEqqKPojAv7VlN2jQmSaYo7O9ZNPC8q11YvI8DRAS9CAsl8x9yVjOSW76sI/
ZYhx7xS9n1WL8wXVf0JnHGy2bMQMf5eItP/pUqr8C5p9XRSZQzwn0uanIlyM
rT/6h7AiLo3ZIx+HMDke10pK/WO8AUVJ8AksH0JqrMURnX2QHwJ3UCm5kV10
2n2UzmVXnCIR1abuIEa43zhwuPCZs792WF/3qYnRsL1Ncfs9kw5mGTo9oHUz
cW5fkqx2BokxcAd7Or0Wf2ahR+6SE+TOhK8Wwf4kwshirSq/s+WcMYTZODbW
QzaFa89Uar7SSn91X15xzsCTfJgb3HZ9FkXaVSpNW8Q/13YnwZNmcJi2Qqr/
TR6vA0DE5gcGFwjXHTi2Cld2yMpLtfaaJbw00OIiwwhjRB3lGU6Q3B0kE75U
5H31JgxmYw4UtHnxFoRYa0xw39SmeWZe2O4p3owPq6ugWATLsGRP2Pf+tH3M
sGqi75KaIPje9/KYBTLKT03PdX8p0vJpY3pWSfO56h9p07ge+74CIr+90Gcn
w5nUWnq0L8Th/eSV2A1s0ZQ0FK91DM6stIz4Di/668dNCtoDcVQh6zJVbrPp
yoZbZ1d0Qa5NPKMJnptWRsFtTjvDZ3yIW8nSHstg8CdSl6RkuoYcdsf5zODy
1bccaDZjr6TYVKDLv3g68rks6rU3PfUebnYCIQuMqNSw3nXldqlvOD4dJ5hB
S/i5fqxljifl2C+vbkQOjfomL4C5HLH/MddkX9uKKJZDkeqZ4OgPDlNhwpTo
/1ONMKk+HHnxTPF3d34Dsuek8bUaeglDmPliMUVL9cxekzRgJO7qkd558NKk
0WSXOY/OhRKnJR1Y1wtJkBsGNSaKh4Azpv7z0RsxILZJenv/shkPcwFtANFN
ogycCvjTHNyXgWg8hmvj6t5iTACAK8HIjafAz9SQFf/Q9WLysajxqC79sNXz
3HtU98WkPo27N+6RFCzak6Eb1wUjGNX4OMOuTDdr5gqmjQEN0Am83ewX1QxR
XP04IWaR5LxaJi+FLPdzifnCVPKGIaoqZMWYRhEZ/pDlKomgsexuZLxdVOtS
oNKcP53f0xugSJwkz9/+RiVjo+JKNBpV/e0WuK+lKL9ustvht7zA9vLzAe8Z
ScSjZMUccm4yMo9NZeWOPNmIGqWVs9enF7SsGqf0KisvHXkk1vDmtHMUNX7h
x5PPLiGDnZEoscsZqCBQkDYGlhAdXUTA4LLt3JbH/Qw8CMkRIqEXuxb+Tx+W
V8Q0VtQzzmcnkTA45P5qo9KNnc4jLKoLlGhfGrGRs8pvUYaJlhtyKd+BFJ0t
HvPy8WBlwU81Lam8VwyYHXQzZEjr2iFogEEs8UmtlLvYhsVUA0GO2TdjMzsU
ZRSAB5XAU84Pyw60do1uEDrfVkK/qjkYlfqpE1umlkW2QrYsmyT6zjN1ghbZ
jVulZ/QC9GGuh0xCha4qMbxmQ3qxKGO1mzADTluGDpFm0t7zUKZysskDfZfn
w+jn/JKwIRor5cbvcCOJQ9vqou0D7ngyu4g3wmZiBdl9b8iQQVNMz/Agsi1N
cIUqhDBpIc8YtYs5oUqN2xE790sjgummPVsZYynxGo3/ihhgYXCjUQwOSQUs
fmiX9PuP3r827aokgSYQco7JgB4tm24ROoSNUp6Kr6le+n+kRZsI14I+EyRT
9i5smsI2NnRD6d0tAK0JWyuko8Eeg44O6t8aJelolEEVKnp3vXgg4qJDUid6
xFk0CFwmoZb9WMaBCOrf9B6M/zfTBopJCGNHbGq6b6fphBrUUnKX/1DMAS1L
d0j1bq2d1Im1Is9Ws2tWeKIwYEWrALJLhqhlxj0rH6d1nWjM79dF+C2v02QR
Ek4ENuLVbMC8un24FAbp/7pbtk5Snj/cnKZ5H6VfPKnkpq/1mJXtrlNRz6gF
htCwGJqQY8Jbx2uP1LBtaW667eLeV/slFg26wN2BfnqIzQ6XPipwjFw9Vxjw
QxGQNrAPz2MJKqcB96lEjCJMRs0zNu6balxmUW98SMBouyADd9zrHdVyyR9g
R0cvsjNsAyrhKcnm5+LGeaStmuQKsH+XfNC/dfqVgTt4yMv4BSWk+wurKBJK
y+W8qR36XC0j7L+D1BBRg3kj/Kx6imWuvMc7vFFfTWHXUuj+A4JWIvUGecMg
Hcrb2hkQp9ZKhrv7A/AU9tYXkbP/LYkMtzsVHy72IfGEUrj+ejoyfJsic9zK
EVM17kyBZczahBRPJ/oBfX5Lvk0xxpletMZnniOdOCTkzVRYHRcGC4dqwlwO
xuHb8XGVXb/9/BuGF6vXTuK6WnrzX1J2XE8Gi69NBYIavF/S1lmeaedvJ2Qv
ZlpYoqpZ92oLWkz9bj1e7WyNDxlq9GOC9Jh4MZieEJaX7BMmN3wPju2YUufR
xWlooTocI1QuLyPOmYyU3zldTUdguYCoBEq5jL5ifIUZezkSAikkn1tp/Shg
PogNi+Nd5K4NkPsXaUxmmrBtZ2/hnQDvu8SZ9rlzW3smqJSl1IJw1VglMHAQ
bASRMv3d14LsSrSm0zEqp0As1yWIi4u+vJd4eCo/xMja8ntn8s7oEPjtTGCg
8s1mjagwc5XV+RCvdOEiuW2STcU5E7Bx3KFyqbOIg1S/NQE1LU1VBRAcbcN7
j4Q7qQRn5SXkPF7oQyqxBcVwbnLy2JPMu4i+1rcPYVphEcIF9PElBA7LMBOR
lMBH3koY1EUqhMyF91ccmlIN1sF/G6kZ2ouwy2YETaDrKMMD3Inm5fwD2kVA
wrDoVf9pHsI2BmoMrkpKrbiqBP7I+FekK112p3jBID9xq5WqJMz0mS+n2B1e
7QrmbGtxGE8nLLdsUJXTNszWUzcMQTtkdvixmX09OZRZ3ajSAXmsGLg2lLU3
TnkMv3H3LlQ9qlOx50O7o6lfJxMm0Zrwa+1SyU2nOIrU5KzVQUZItsx0kEh2
d5N65sgouUqjTFxv7Au+j2pJcBFvmKFSqgXHC8CY8GpeAWgzuBRQASfMSifH
SX2flN89W120tEc5ClD+QMVHZWplBVpo0W2AUWTfgBGd/XhdJMCFAKIsDiln
1oQX4/Gg9OKzWu46KOXMjUA+zy4v0WgEHzQQ6XnPxgF4xpxTymy2ZoOLjJ7P
92VafV7x+MLN7iBwWRFrwCbIZbld3UGc4rreFLjuPpLi4LcNkdFcu6U2ZR/T
FBBeE/K7CwbCcaQ3qFU5Nclh1laIdoZceLrrT1nmuwEDE3tOjcS/HT+dCyLH
xQLuLwCtvBvZflNul2K32GFYzLfn73XxLDoCManelTiQLNDVwhEwKn3OCQii
JhIwS0I89O4as+iaFgN5hTOjFFWHx1vjieRYqLerU+QK0+EI4vcf08c4YWB4
H/oNz3nZ26ncKqvfs8ANKhDYFk8hsOUoquEJapxefW8YQDJathMbJQpnhe0o
keNEfEB8XvCPEEOcF9+qOXHWHMFcjGb3dzg85r0kTNjKqeUFKtcd+uh+QRNm
kIH7hfMRpauqkcCQaak7CmIYmjLO0CwXNWPwwcvDztwmoNmaTehoKx0Rq8WN
bLlb5GF4QiyXfDNtr/ybGyQSqsfhAwF0hpoWfb00LAxJsdau5YRlSZekTXtI
X72DQTcBVJelRRc6LTsGk0mFJRuaNUU8RgsP/OxbP5K1DQqOqm3NTE/pRg7J
o6DvstTf6MIa3+OwyVZt1sVnsW6GU47RSA6DDIA5v0F6+SaTB1pQaS4qAn8A
EW4g/uB2pVRNUAOiXHQzvR5OqUwobSdpDz8kXx4tWwF8KTux+TDCJ6PNIlJk
qhcIhzQv8VMZdyLyyrwD1Psr1/TbrJ2ji9Mm7tMYTHRjbqKOB9DVEg9NWpuj
GS1QlgoDIHE/CFmk5Zp24hpHHEpNFMK61c5Q9ksn8jF40mCCUDPsa/6eS5La
OSGFVDURoR9NhjdN9WElfcTwdKsikbeZa7guySDpmC8/BFmv85NP5dwNtDlh
ezKwMfIeGiUA5w/9m3GFdFRdO5v63zASpfTssuexUQkW1d0b/XwHAyEgwj4B
sb5lXPxer8+AR9ehGgHTqSzGaKufoDAuHcYZq15/1ewxPPH9Mg4D7twlCAsd
LYZu73T047ozeWVM+n90x9SDi0buThZIWMkzPu4u25bdMIoXa2OE44fcDG23
amSEHdO6K1X8ItznXzdrXRNZB6bb+jicAAT/v2edE1gmAdA1eUQWIBn49J1e
vp0YhbXNQBqk4vQ00FNZ4yQf9YpQ4o4AEKQa1qPrBpWG/SjIx6kqnm2Kp8uD
rqUcm/F3D3Xx/xFXFmoytKFqoaHhqpddR9yYwsWSJylxdZiYh1jpJX+oqF36
3Qps/mZ0NrRe7XkiWcQVpXGAcJTxoY5tQY+mSvUOT2+nrim6G9DMQLgUWugk
Scu+RrwcAWlQmB7wK+eafZSk5VigZ9+75gIpNb8EB78sbwASUKuxvG55u2NV
OhsGff19U8qD48p3GeEBMm9rorXFZCXN6Sw28PhicCiTzGy2hXbctSJqiQZa
rnW70YR2Xgz3c0hE3tTxve+al5T+UOPVQ/UuDGoxoMBQychUQJ6h+53E7DNF
vXpCOnkg5TuL+WpEtzxYTRFr+vF0R+8L8ZO7dAhI288QHVqia3ZYyFrzSN0g
oWLdTDo9zXZky+EMSbaXzM1KxFq+Qfol46lkK2iyESf4rCm9U1RLRfY7V9YV
sCTrxoSzWvVabbN7PVmNgl3YKWgIPbfOnkvsU0KaaBJxSq0e+SyFWypgGuc2
oecNzpgmyfg2/wsl4CpOfZ9sN/3WMePVf+JsQO3AEjAx3YeaShxOBmEPgMMH
9o/2hCZ69qxdIF3gpeKDfDnOAYAoG69SgCV5dFkvzizk4jDQMmU+hxnsltGJ
nQmg8WuI2mINYpBMJG/Eg5Si6YQoPnn0T1xeTnCC9dMj0MEYTeZBssY9ypWI
EDzYDYPQ7lb3bfRiWC9o/xF7lomWIP9gD6hhrGmAUhiHCL9JmpWj7/eYBuCp
MnKXm6c3ElEmdYVokB7nBvrpfj/y7vDVMCF8Amq6h6+WbkGsX6AHWSanhUXd
xz2qhBwFLt8fQ5D70ixbxBDZHfY2Q+N68I3JnSKR+5BksNa/DKa7Y6ml+zZK
aQUfa1SrjweSRLN3hGPNCNw26cpq3oS6wgwJ1NjPT0iLOQ1uhRW7Nbulz85J
GbpNxT2l62rQDAl0z91yLOT7puTPrRYoNSyT8IduQW1A5GXDTAQ3T6mEBuCm
ykx+I/9HtobA3mCmx9PfNzZWbl19Yj6SMe/XGsIPeUNKtnUzx9KmjYav0nCQ
mUyYwk56uJakcuFsT0oMmQttZsJIrn8JpiuI3HNNtfCggXL8fyqk2aixJmvz
By4G/cjt+qBM4lYHlKr29aZXZmXTFEOHh+0wRUwpJdIpRzFq9ivjF8YDEoWW
sk1h7NlNJzuev5gGGu1iQStekkgB5qPD46xI6L7IhlGlyfF1PsOkXMYNY6Sg
5lieZ4kDxucfQDnmtWlgeYVUW82/aqHYWzNbd9GA+rMy7OEu8EqWS+LarXS4
a0ETRluo/Asu8rkJNuAuPkgwckY/4qq+6tPw3Y15f67nd50FGHCn6aHhaUKH
qW1xW8e9A8D3fThxnSj9klGZZBnu+8s8nL3U2+wPY4F8zYeTNaqrmxoHXTdh
TAJ+1IA8ki7lFzVsDTIyLEvkuyesknXF7u8/zrOdRaoC/c+l5k+g50+mMnPB
3I5kKJzFEhoj1M4Ph2aBE/iYe2fmnlstkQeD85+lTxLvRpYn/kDxnTfvu+5q
8Ig5YcmXiCzo7sBDkd3xDo5Q46Yf4a0ZUqRoBI9RvJvDnCw2CG6FBrYPeaW5
JHFxNNUUuIWucb8Y2TCOVHx+1hJpkODC0knyXhJ4ZEEHu4PYbsDqgSFQQAqM
MF1M0ed3GrNKPuWVnqyvLL2XQ1e0NSR23uF0fs2erdl210Re1txzCqv6dtxb
9j1EgQsJ77uF56EZv0QrRUfvHh16D2ISe3Xpq4aww+cxA4AJmKftrqEihv1h
GPGScOVY5/GNb4FHLsei02gxJzFY8oAS23M3k1bWWfqQePvgdAix6Rp0B6gT
zCsMO4v6fVvEzaa6irr8KqUPY7OJNXSXvvck4B/ol7t/H42Lp+Gib1SM1pCI
KjMdnrcDKzfIxo1sND0HE2n5n6b/53ikNsy/S/5TJSytVJFUoY5RqCvKac90
lMjxLKwYDC0W5Pub/LT7g4GP4qJ0bS+y697xk8h507KX1KamgJKfHMzy6hfK
gvMNNaVAN9TnXcoNHgltM1Xe6C11sqf4GeXaTLgssrOwsgyAEfMZdXOGPFCA
QIZj2347FC8OLJjkA8yIZ8/RTNDSS3zJIPj/zlSpXN0OKdbBpu7NPXjNE/XT
bmZfn6lM3/yvd7fpzkHNNljpwsRrCBvHrgk1lN2mTxO6K7NfUxroiYn9t2ax
OKG/30o7ZeVkrkTeQ9RKDZsg5YUJO6udELVnOdF29WyEJsTk4UeEuf/0FfeS
VxZQieHiU21vYFvAluMlXbE8ZRuqoVn30DMO2/dYmXHpLWQQZPKCsKLukPcM
nH0XogefWoKaFFZl08ulgHZxVR+ZvaiophYO1XP0J9Au2cckz3J1kBSb3kV4
ui9i2cGfjgZTtS6A9u1+g1+oUlo10rG1qtBx/ebOnjn9z+pQ9WGLdZbSLy+i
NGsX9qYD2Yk7oKjYoyb4LvMlUIiEEdegGTnqpCqMgCV146qU16todPByPpm5
eABmimr467CcC/sUxE9yOcVPDv5S7PW2dzritNLzDpuibP3rMbBNNaDXef4H
GWJzA2WIUY9+mlT4EX6AspTppz2Z4jJGx1eOXbteyRP6m6YK3Ad9wjNa+CMo
D8HerVzAMyzVihkwVt/APwa3ZMRT9aRmuAvea+AnnrUtDBdk2W1A+E5uH10F
kyaRC6xMo3mtMxKf4f8k4AVNlSuuh+duSQ0mC1bcHA6lKT8Ov8vJcK6QZB4l
lmkcRr64ia1ZiotTD7MkOZl42NkJdRwTPTyLmiFEP6UabAx2vgdyRI4cgaLP
B2PaFd3uVdbmi/gdKKJaleKF96zRfQP8SsKlSp0vRfEXdZ+7KoWlV99HeHkL
D/8b+VRPD6jIuGDeYPhJDkccJ+3pTo65Lo7eKhehazQEUE9DgxZoveXFhPwl
HVthFqld43DM4gHXvJC5/A1eI5klzg8UtzFligXKlQid3isT0F/pBAT+DiSm
wjtkzl0XqIVfSyeKdBeC4XeZmP3Fpg2nsJSnHzHm5yozZyyUziEBw8GoigUm
HSRlRhwDl4+7nlcuATPmqfD5Uc8j50sJieoCIVwpEXpZy2bC3qQcvLglZUsc
Omf3wKAQxE9lHczmheF9agldmMA+I3v1JFFswfFNEoCFZlnAArZT/1tyTUvI
Vn5Ig3QaMx1aGm5Nwy6xS3zpBYPIljFghS9kbxVvRpv7qkaDgGUQ0I7Ds88A
/CJ+FndQAaRQRFxFfnvHPCEuihUVCrRtj+/EG7cBXHKY8cBZYreiOS9rlmJ/
YwhYjvDRkRwRbuMIvHRY6e8pK/kQOn7CeGPcIOueUfEq+jwiZJ+r5R8Y9F8r
c/sZnUyAovkDLDJbr9gCsE+y3HipGIXUklGHWlyU4IAweN5YP0Izgp42gxpd
BhGUQUyhzj05FUEUv054XgYnfQjQWCvMkblikOma70uKDEOtaLen0BICkeCs
yj3JJFSq+OfeEh81QIQFUfuwmDHkvTIf07xowqsjgz3o37xZAEUEsJy2ytwM
r+uzuekkVYOaCq1BSqlNLxKMBYcSxhaFeL/im3MuepQJ18HTktZDP+MSR8Gp
uuQf+Fa1bf1tsxLaC1p+x1+Mq4o78kbhpDGOA8QRn1MqLf+cO3TPgZ1Q/wZL
7NRoNhsSF0kdBgNy3TqQvp276dtlRP3a+VU5S0hb09qlneDSq/VyBYjZvEzP
GG7MZ5LUd5Fp6oeCTerjoapBH5nLO4geeotMsg+F2s7Q8lwSbR/SU7lDCJtu
6nMaZ/IN1CqcfuAzKvyTrD8KItRa7OVhTP/ei5l+cklvreG0R7TCtb+vlJNd
OIsPeKxrRL87sYy+z+9XDkclDdrX4QO0g1Y92tfOKS9Bx//HNUzaLVue6tuI
fXi+llQGK7IrQmNXUvZkCLwunCWmwSia2J6jUgA+lm//5M7OCPUFhOfgq4Lj
FEZUvlLWXBjmrrnu4tmlKXAM8dHTJcQAecH+xvA9j5S0zTa0yM9fWY6+Sfwm
eXC3vFze9C0L2y7C6rYdnzjNPBjP4SfbSeDShOV9aSDkoFzs77xmrad2hRf4
iuL78mHm5Kff5NeorVTCVo/3UpPYNflAPZmgiy/BuTLCtz/rXHq9JAbKevbI
m1dAb/lFRI0HwaVJgnvRUb2Ti5vA84G+R2AHDl4fB2Vyn+4Crcwy6uLNAn66
u4Jxit9zyvWR192lWxyMaaGdGwBpbLY3/0QIsjIsNBl6rXTCpKy9c9uIMmCr
E8mJvctAaiW7uQaEk5MS2vkv0/FcxKAWeMDbRFjzsc2cnAll3j6NFjqeXO7R
9vvgQFDrtLPpodnQMPytOOq7nRRK1z3FfeiN0S9ObZj26riqON1+6y16Yov2
CRJaZuaJB1R41hXQmFK4DslpHc82IpK6A5JQAgUGfpTIbb2aUG9M7jJ0h2Zc
856yXoU8bUcRdHBQPVkSJTUybmaBxNewVbZCf2+Pr4WmDcdrnDfoVXchtVBx
KW8ffazgSLafYIdsiUp7cGo+gemPRavgrM0pR7QLF0OsKO7GTWVZZ1Ry57TV
V89AhP4tMukBexjLpAfsx7AGGuLArPfcQo4tqaLejiiEs3jhtRdqCjP6sO32
H/pmbTFxL0Em6f06UDmDaGkjnAJF5RPaPUK9QihKaLCslyS1lEfk/I+uGe5X
boNYWWXrB+aOyo6sLSh/Y1JgDcLPQeUbblcT0RQolpHlBc2AQFpP+df5O0PW
3vlj7NM0bWnkVm/hTaOsla1Jb4+Q20YPcDxLYHLZUkbBxBoQJkaX/FWVVjrm
izHEerHeNovOEHFLiXFSApgLGKQfBvVDqYjVsmOPWcOhH8u0CYbXy+0jhV23
qrbRG4s2wfGk0yl69PYVeAIBigXd2ICWjuhrrv01gkb+JG5KdX7krtfMRNIB
Huf/d/KQ4cz2VKVIo2iP6wBb4Fdr4dC7RgEgNLuT2rI9eGC0YV8ZPAE/VihW
SLtvIP6uaepCVE2Omw41guaFv5uesMeEknK9EAROfIQQOCwTrNOWUfe+/OPe
eZW95TRvTa4Fu7ua6wA7c6LBBx+DrJ5r+cTVeR2irIOsMBxbMpIvrhbNoTIi
bgMA+FFj0omzQb1XyJRqKcFnN3ficxFJ6cMdLVll0W2jvIZVvYqpe462JdMO
JxMlS+dkhqvXnaiuQUExsNmdFD6NN98g5hvb/7Vbvx8eQYuCmxQ0BUWYz9tZ
F+tabtiqRCbvd0d7AxAlQ9hZcS3b8TDgAZpQpnGrZGq4sgiB2N+QZIPfxHzY
C+8vUb9V2rwpSBAYmbfHdMHT2MlwrD42ZkG8tOV1ukqi54bFjVWQnP6MVPwX
1gFOBrnVUavp1Rwv8uFEgOWscdl98hRWwN+mT+xR0M7AHlBem5kPptE6tebh
cp2bVCYFjUmtLZVprvYtTB+4blkCgDQAc/2tAW8U0L3bh2yMnU/JGrG7xD48
xVAIdGBSPBVAMEcm3Ne1NWJd/mYmZ09T23jpKXCApLI2ghCsOmCENsv3lqFH
P6+PfWMFdSjRTfOmY/v8I+H3DP6SXPGM7tfOJaz5KqxaWbVggi8PSa/iKnS6
dLvUCZfGQPgNcgtjActl1OK7wEu184cLL3jlJhzkqREKFPBvWd5HAaMUIaoA
6/O+0poNMkAQx5u/bFfo2bGfKKxZcOpe1uFuSrnArmo7jZE++gSK6kJ4Hrcl
Wrpj1wrAy1n1EmTyzg3ANnsAVymcOdwSuEdYPfTSnc/iCbV7FyowNvu5sQyj
YLoP/md7SNgx9HVjqYZv/NbjZjMA1Cxbc+mWAIWdaWuKcsbuT2ZRT5oYS/93
MLALqUtrNjhZIZF3HX0+cWnr65C/pjgRy8l86uyLj51RH+4ogUYAIaNlHCEz
ZlSPcAwfRcJbIcqDP7K+cquTCK7TUKwm7OKs4fhbC70cZ47bpOwUSQv9QgD3
Wy+pOfPG4zdYz5eJxKMWVvrERebNH58D9MPf87hA2QnDHaHxQOBjbClUAgWg
/iPEJZnWLOjsCT97/FHIKVYVt9BdmrX18tRazNTwVOxKDV4BgjbdY0zU2acI
llbKFNrMN14V6Uzs1ySOHnIxEr6MBj7Wm9wmHLkPL2lWdzIanpciXHmL2iz9
fETE6wf2OAkCf+fgb9OU7PQTjv8rMdOD+uV1ocsQHOQcGkt+jZJZLy2Jir0c
C0CELPI5lmOMw+LXo/7POiF7SPJmwGLCDQjjnwGMCfkMJGx5P55FTZU9an1H
ENwojS25lt2iKwgTaFNTsK1vcFKdr4+UucGmOCN1x2pdO+h/EFGmC1b8qRtb
Nco/MnOHXNMupT1WJWo+CvbB1Kr6OrtI7NIaCN9/+bn5ctuf7j9rNndmjf02
VNZIWjiVK1Y6bAY+Qfvs4BKMcKgFzBU7SxMIM6NxY05vWWVKl3dlYTp66/+n
zwRTN6foIKM4c2o0UAZwi6qGL2OFp9GnkxlYwm6p36TjuIciq9DmSlvsh8m+
HodP6m3Euk7ELjftTshllYhTQ80/Ey9e8hC6kfRTgcjYMgIqLMnIgGomOe57
xZuVKZG/wuRUBE2QlhfSxMry1/qu53oYvx45uRP1L8ojGAAWYOFRzpT+CiRD
1/KmxzLQiu24Ti7DRf7fDwlzz1ncXlwjnd2IiHNIG44Rql5RBigwndstIont
tkYWPJJ383K+HnJ4iTiAaKaXdGy5gvhULPKJDDiSu/O4g+ZksJZXbizb2tHl
2zi/L86wGgLNSmdwOyQ3mBd/Ww76tEXbEFKlJRvO0qtEeeJWtrXN1ibE7UYY
HzFGJMGeKt+xw2ic6+tRDPqZrO4n+6P2VbpjG1HNkHW71hwVbMEppPHVDFYI
w/MfX0CAFmEiKRddk9fJlurOdKdwHhLXgsURH8Vxri0LC7JYjmK6/p5RiWGf
dNnuMgnAP5a92iMlJZR7ulW7fKOEUcsTZQAo3SZZHTDZ77LWWROkIv1Mii6f
iklaEHl14inAQq1QBCPPT33Bs0cFKi1Wyl2nkEUZwsDe3yR0f6sECZVeMmIi
AZE4mP+i/yvwnYcFw0FHGVzBKXNSRAj9kD8Ea27j5r2E+6egWsbQ4vEUvQVr
qyRHnAc+fLTwzswe792biVB/8ydrTmUcGlCLLcL4QDEzc4I1G67BnMmllRsL
G2SQg/Roc5vCODKPYuRi4TdbYAUrLw1lKSCrbqIKYOifGaNBJU7+RzWOnHO1
4rFAx7pfaGtu00VrzgWZbirnX9sVxjXa3GH7ro45vJuQvbxozmrAYnnM6kZ3
fdC5WOhyivRhDrNxnP0DFJeyvXQjvqFjANOcFd+qHq9Ql5MIXr9L9XqQr6+G
uxLaTT7LT8l6I/dQVO1OKPoyL0ow++e/Rw1T7uy4ntCMmEvYoCMRxM/s5lEX
S0CIHMX0V/qXSXbuNkfNRA7Mc0Sv/tBdieQS9y5i6IGz8YlntI2sua8fNkyP
52ZUi76U7ic95VO0dAs81zH8/skjZ+XXA+DUNyfVR+iERLk4Q0nAfuQay9yO
MSqRW+EsuM3fxfngmoXlrBqN+ffuIsHlEPqKeRRXhmrF+HdfobkBuY4ymW/a
F0ybbIuLJYuvgBishQRBYt1tBT9TBt00LtetFGb/0XlgNanPLl1gGjacSSmd
1GrRgnJZxibIAjRU7/ESPyPDlJj0e1ZZ6TFr/g7sSwyzXUUSe918MfBr+n0a
gCsYKKcEMsRQ3j9qJRMVGX3e9rh1zG9UsHMshhN6aM9JF8/VnVSoRU7Tdmlc
+FG+BnUT3hdN0aDsiDX0Lh/UCorbrepw8O0OStnnuz5fAgyzGrvO9d8BFWVk
XNRsuOk+XHDz+N9R8xw4+VoUkFSPSIlK/FzdKDhRnK7q+UcJD8cUpT7JtEGl
ixnoOCZVgJ5paSAcckDvZMc5Na9m+TFq1LqhExnKrXcAPGcashqkx9Bs4qP6
2/E93oDOoEUfsKYxdraKapVERWuOCxMIQ+trJL6GESNi5ARgd2GX1hET4Dt8
55+mhCSFlhVKClZDYIUqurJi2zXJfhs94kn0BMU4D1tCJHJvP8/WqiAmTZFg
D7D4x40xSGGzgO6Yye0N0H5Z6CCHkrmHv7ch9/Rqwo6UV7eTFvQDPrekOMva
4aIOOtflfifdPgmtb3YOhk9LWZFABEoMnEpzBEEzKXqGPyU2Ehz28TroTT+t
Q0IJAAinrr0o1Q0rcsRbbHCTsPnqdWJ2sSfkSVqL+2BNc2uEbLpCrZowWB6F
t8iRakOynaNVJ5gSrHUMx+589Czjc876t21/fy6g9+88rNfZ0goysbrbZuK/
GO0/V6Z5fIAScbGJUlRO52d5IinZaDGBZrq0ZyJpyNTH4pxj6OM/4uBXbHf8
5TmhWHp5UrESKa8LF9m3ojVtUUZq+Vam/aveu7an3rSOMhIghmJBIFrOfcl5
UY/1j3P6/2WIez8B6mn7g5ycvaJ4/uxv8ytkU/O8k4YTP6/JMyScfGpTZPn5
r2D3ucaCD2NVLvxNiZZL4MYtkHPaZRYo0leMfCb6REZsgwB/c/3m6s90uy38
4Pkmst7me0OQFrsjJOk8sX6Z8kCmxBqwryA3MEqnFLaOegfzh+owh9ozIr+d
RVPFOUgH8KVO64FHCE3w3P0mjiiLQ+EEKFjvh7kvs0MNIJaw8BMGSoZyKko+
wG8dw3jCeOkHDpqHg4zu/qpB4Ta6g6xBZYKlintlrM4J7dO7F+9cqN8oPa9N
GevJSPczHIvHqp2ExOxHA69rmNaXQXDPqzSBIFESpCpz8aa1CYCQts8xT0DE
cwjkJ4QU0fQuhQMzsXw1bX9X4QeBJtFKUXVE8Z8Z4rIcDJx1u+gklC9LUVI/
o1klURe4N6TtzE9CU5ZrS/b64LRS6PKn423d8fepBgxqAFCUJmRslZ43wTXi
zmBJaMrwFBjWy1ejT4jmEGkZ5CRhzgjz2GUxGdqREF2PjVMl4l9dNjf+DopX
LE9hsMsKPy6yXo5EDjRYYZ3xmTESWcZuo0ygNRMZlVL1lJMlQx+o+I8Hrumx
zsk5j+GyYDjBHV8OEPhCqY/ykrali8eY1cGtpFxpHtsSbDg7ABoSowdh+7sN
00QXL7sAuBahAJZ09PxZTf9GeyXIqbgkpu7P2MJ0gz8xF3DCXqESv/4pIZgk
/Ll1FEPBw7NmI7dhVkX3XrMw+5FDvBJo0lwzcNuiHOou9yhAdx6SE15mJVfQ
K0iz0aOAnqGBOVLGlLi9eBtJHwJcLUQbqJlnFEsqJLoVnwbyPf7DA5GVgS+U
pcxDrmlBi8srSgEMyf7EpL4PFJ80am5Dh1PbePRBZ5oIlTkEMGJHLY/xZD7F
P1pdjEscUnwb920bf9AJWcKj1cA2IRH7j0dqK+GdyQ9l5IYqEXKHEbk3Ec7F
faqPMPo5h2MmjcTZp/f0yE64p3VNvNBmvtwud9p/QBvQ1aSyMTCcSqXDt3RY
8qiQT6p+8Bmg9l6k+5sXsIikraw8JfokRDFC0AaiICXjnElnPfDrYYPL9pGM
g3nhpOPwxYEAdHdLpzDdFiTNVqeExnPT0cAlzaUhDsQ20o2np/q2ldyw+cBH
nnFwp4k2MN0FZ28ub7drSTH6dZczuE9m0F9M+P+foFLGw80ZErMZu7AGxyft
20uoVPMPti8rz/Bn1Jlm7XWHXcmU79AMepYn6sxoY3lHM90IR4mUhHScU1IT
hH1JscZdreiX5oVWLZj+emCZ/rziyB532FqQvfHIFhKiQQUSCWLL0G8Ha7fn
+WZa1bYMuPf9XpGRIPqxteEH36nRw6lITtpYtasXboTMouiS9a4pI9iW5CTd
Mne093TjueeFOfppbSXaJouST6F1hdr8HRC8jemYNI7zLLtvXVvTlPJgSx5A
UTzZD0C2vvJ5ljb7Tzc1YVwZTMHLg26mq3uejmWFJoSusWPjEFAALyF2DHn1
XvThRg1q8CGooiMzkmFbzNQpHKRG4R81dw2a0unyF6dDtftZYTM5EKBcMi56
A7/plz0cSvdSZwvGhJO/UKvi8WbXUdrQKa46ACxQxNY9XDfmls1d0WwOaHMA
PMjVAr8NE7XONArdWx00h7J50C3GwjKq8no1IZZm6DqOhn3+llPJ8EAVDVWI
shbjjLoiS9JgnUpJF5E2+nk2w7l1cZ+VXdRDfJh0mbAGvbfgthW+AGz+ung1
git0+zdUdWSeVRPvKVC133D8yByk717aVOR7CdBCN4CDVHvG6WdZcmlCk1gb
Wqf91bMSsw+WO0poEgJbiyC0O7buJP4Qj2cR+UrtkNjD+yymeeZHtljCWRUK
iNjBa6c3diCagPazIpgjWkXhg2pe24R9tYDytZwhAuKNLp9ejs2fYeUWBN+Q
5LvXPaLzXXS+CH8agjm1zoNk021T4jLQXnTQ+l8RhIFFfdL2v3up1egtgnam
D7jQtU7rb+ivOxdkq56oAvPxppbWt4vNZvqqeK2szpx6dY0xeEYVW+KbZB6z
QI79rGSiz84JYZjwuGw6B3NtW0gEqwiQNM0B5UqSjud/Bi7JoeSyGjxmEaFG
YZE+LoLB1eNlWu1XZyoMSOwRMFMgZlrQBtXyV/k21acvhbNFMeU5vbi6TBSc
pcghM4d/afAd55msCileZzoi+poegrY6Yswrl8drpkwBGvndg8ychkPk9UZ/
nCCsuxpkjuIaSklbVX/1i8T64IpqfwrbqzCY15rCjNInZzjgxteiAFApzR4c
u1oawYuL0BSJhk4D/h2VBlG0xIQHt+zWgxg9LV3MDl2r4fJP4WBOIGrm1EdO
reN416q8yHmaYXL6OC0GZOshx/RlCrVpYbvHZcgatpimv7bnrhYMSemkNwKV
iKHLp9SgniXujiUFddHTsl5/aGeCQrebX3GnL7UDSvIGXThM80mli60L/Zr5
+y5vhvPMmh0ePTlaVFpWwZxMJTQPtX59ojb/5RqQQ0d+ZJNykY8Uhr3eMPIk
vD1hSPqAbT9/kaJpidu8XGYa0aj3q4FbQ2kTIBL05Cb/wBCXSmnJBkM1CCkR
tmUAFBU1C7evN0E+pwzoPWTg1alFMyesDZ7jQH41/j9XDLeNNQTpQ9Wwr7JV
POxyqCeI1xqAKif1wjNqwrlQuNUuXiSlKvct/oYbkL2/CBgiuNR6oL9fKNd7
go491019oMQxcwa2EBAvLUxSnGG/ug4I6b2WYGXt564YVTznw0VNcFSK3zgN
Uph/5Zt1CArL/DHQ0OiYiFEMPoDuVayhQYZwn9HTvWOEhx/Ivd0EZMWXglYN
/aEixvyRxhfJql7KIVkcst6JjWJYiSgNndRyoJ8YVQWKjslhltn6S0/PNUdM
t2za9lcYieTiDTLkp8GM79d3qXvTj7CJumxFl/Yt5HjMhtqedYszy+kUa1e7
LeFa5xDz5hyg5gkDU+vilQ22kmfnGrMUYqapTvtfHWgaU2BHdzhLurjNXpnQ
5JSl5mVAIIZ3ooHjcZJSM5SdsCXXAjGo+PWtnb0+fYZFDAiKIieU6yWIYsVC
P0EWaR57ee+Ay6Vxxnn/OuuRmq//NEMnL/uc1fddT+hFqkz9Y967JbxKLolx
wWCepm0GzcWEgO2EpxSg5Tk7V1AS+H8t2AoybrqW6XMCnwt7FurIUiRYCrpj
o4/4ijhS5/payS+ZC2JGh/ZfQt7WC+hKUYGlsH5ZKAri1sxaxe3k52jq3V91
ANXHSkAw3D3HO9a+hVTHjOSRBgVmz3NtuJUCsY6Z4VEmI/zQjsiYNPSFLVI4
6Z3sMzAbwLf95Gyz6Mz/vnH7QPKCAPRoUqdApX/AyqL2Z701nmIk356y/PSt
KXjqPsYnV1/Za3ijrcOV+qD979ES4XQMTKEP6QSPB7mI1tFbilvogScZONWm
J94isaX1IPuHpnus2FCZiQ54dDvcyfjdgL2X07X9VyMm4B294NHkVfP0NyFc
cmZAE0QuX8MDMVVhxKg2WX7qILN1ty4vADzdl5F8fXCGIaSK0ATCTZ/oa43e
d+NmHyPyDrnAeoiquGOtakkd5CB6e/fcr+Sn9JWvgN7NQ7luYfYwXALAkT+f
MiqeeXuUFfiew/bfgvZ1H/BwLq51wpy6PB08RglSdL9NgX3U8N/ubwHwTeLR
Lgcu5eZSzexbi+YgFd2rTMO7cdc6QN3MnkFWco6RAr/54Lm88XBOMKPcHbKb
Jr5Qb+/hZ3xs+Yv7V32EEWRoTmNDJyqmProCReMcWc+1NyK7rs4XgfzZlJX9
rwwPesJTbrVNNn+xemttgz92ZCq3TXh8XwXpze10fJdky/y3NlqhVnXERYSr
MlWeHT15M8N6C8v0BN3wSeQynIk9kPjSjnzjdRNEhv+qRtJn/WQAE2WQ0sCG
u4j8SJ2dEJbs9F1Hix6XGbSwdMH5eoNPqL3+D+lwRYLLe9pY6x65LYS09Xmz
dHyoV3VtsVtUnhtZlDfeL+nHHK6upJARtUK7DeiBbuPs2v+1lLObdcqkRHR6
iQI6zlXXFMfMSlt+vKvWIs1rHyk6BGrLRWXVw7mDOSB0ccjjUTqOECYER6A/
HdPhzMQx3nZs42KNRsYpyZs8veAx+zjzk4TvvDLLA7LJidn+tJ6urJNgZhkt
W/NZRodat8oVVtC1TqWNJF5bDTo+4xm1lB3f2ymwPfr/tIiM6AoGKPqYQqc/
SbZMJX7MISvfcQzcdxoNI44VmPVs4Hi5my57yDLkoi8ONKGpIKhPmFeoK83y
4XA1EW2GgjbEyFgCMD9Itt50YVUMn+Mb7JUvkGkiRwoTYjvOPBeutzAXtskr
l1gtBFrF5UsVnh0w6n+wj7v63KkFjwqtH8ZEguCWR6K3lPjAp89oZTCTtRRe
J2KE0GTcIC32goW81ZHgWassd40s4GdaMd/XBKyeyfflc5apfn5gAjlBBKn7
Y+ZD/vN7SclLAC5IFrr8z7Q0eT8lugmRKwEGqlas8VmDVYN45sMZ7zncnWHi
H7VeROI1AOmS/aytQBF1ldzOY5lpmwIlnR8mvavKgxQ+K/VY24RJkDP3MhJM
YV+TJ5wDujwI8c0O45s5bCJagrc/9KXmrH3HT/IjKR5TU44l4AnTap8pBr4r
5Ty+W64Ds5VTK5MGvyJhLVy5cFf1PLC2KQvH2oA4h2INxXekybNXbi702DMN
iRkbOSC+uiP6nLOLlx4G17AR5SxAFAT8jRxnjghwUIDDMOiY6tBRktChoQzj
0xqn3dvVM93RpOg7aA3dRmqD1FK+A8wZebZTewVUQBlBqw6Irf2rAE8j3M26
STjlmk0T1UNAgWeG7qzUKWGr5ktW/5cX3gzpCXZUqqMUFpm+cHX0RkpIkvxc
EM+rhCk9W0ZaxZd69T2aJysWKrX4WUGCoAD/hsaCkCoWqixqyVJEzIYX2jQo
86MFJSY47EnTPhmctFtPSfoD1JcUxM06Ph+3RiMlAUSM+czOIOEERMR9FL2u
EzQ/HbIYC8oNfsnNzpALc5emGf6l3cR9M0vByI8KMFlRfR75YmbEft3F6hqO
kpOCHkuwUr8CJ3eXKluIl/l4XKlCXQj/cbwfzyDZwALbdAcRRvRk6GQFQ0D+
OaFYxtP173FslwQCCiXQEWRIgNokO8p90Nf/ryTNOkGD1KqNGPJj/3xDc7/C
Je5pw+EhEe039/FFO/gm9BRXbYLLoq2dvM6Mtp4P5am+zd5YxZR7oxKMXWLz
8KEngok/y83zv8mOuWa8pal5puLpNrywCBHkicGszrpj1GrzNO6MUbm0RUpJ
Gw0TC7L0rA4G8qp2BGr8qcBVqIynASCbxmTrtA8L/kXUqVl04Ge9/9PChsE2
G6fuj0aGfzltYhEVPImba52E2ynBbiuK1Xe3X06KymGPYXMh6rDyPwy0qeOT
aYxZuJx+4X7mVboSVWvErt/8SK+LREcqR5mTK9SV0oFx6NhSCQha5uOLfsuE
2gIBlErIq0ZZzlfzkNaakKYKzeRF04iap8AeH6YRe+AP8K6cAROOI/X9Qmhf
oHNKIiNjNEeASURTTGVCyRh99GtOJfoiywV/eEkMRpLuz7eBBG+0gT/jcqey
ykCJFTJLXB8UYgY3Kp/0qmn8ouVgsVCE7/5dVoHHRVnDip0aEgrIH+0PDLDs
E8zwQFgmPKz05bxk5vGRV2NHsEudTySAZ73/00Yux2x/PgQX9GcKnOMYuUr9
g5HY6pqR1l23yG2AKfPVq6uZgiz4PyB+aFoWVuOutJlTAHeI+w6TTol561pz
iAj5xF+n2CwfqyGW3tP2cU9sLS04rV4qKByKYNmsUmbUsiEyHtff9IiWwaUG
lyF/c+/6+1l2v7VtXF3Vj6+Qo21lqdtTI15Kk+FGjh3gL8LZML2YKFxFx4tS
lY6Dslz0sCoOZD9gyvlENFHAYlE+GPTA4lk9fYBDnpXmsV5Tm9499LPczmM1
8cN7Mfr/HIbfvIQYDsZqx/D4gFn/rj0svDy0YIlfZgrMyLcRsqNUpML1fSHo
QgDR0j8f4hgOLY4OPZseyPUV+Cf2HvkIFglwUdj+XVvXNI3b46RLUstzFflw
x/tvD2OZHfyywPBChV88CxxIli3EZIeHz1sjNe0zjRs+Y0VoAyHEQrpAuup5
1Ln1KAIgddQn2UYj4DyK4+62vN5NcbXr0mmPVIxN6WD6rTtHshELuf3bCE1+
IMzv2IE5thuNqRChL1WC6xOUymMLeRCWVTjc5hvqNahy51wwLy2w7Zi2YfSb
/STr9uBvBvni/7h9ZderLrroQfrKsIQ3lhmuqU4EAmw7c9LwuEdpq1LCHsE+
nC1V5/2oPX5JfITflFu8m+29Dw7dtQTFIw61g2poVcO/uihZktwJn0xGQxjf
R80/r1SARm707G6Izt3yg89B/knt3yP6FwqXjfnaUFgKexnM08/Dmuji/l9v
qgoZt2UPcie2P3kGaff5UXnV5fHefXR9NwNyeVDGoefKUt0FBoZNOdDDaAyU
Iv8mx/KWNjTrOwc4Wk9TSt7W+1fsWfw7gRDuTrReeYWPIiH+IPZmdwcrSElZ
RvmXxHnGh+V2bsXJ8eNRBwgwErzvFjq7TPOxdkSBcAmk0MpnP/dCIy7G7043
jxxCpTSWqD4xQKt4+jE1pHhfmPAHt3x6xj/V8wBGXD8MybyhoctZfsjgXuPQ
z/p5jILvbSnqPONpdRc7lkunEA/LngU4y2pFqDPih9Se0d//ZeQKaHUSrOJq
OCBJ5ZXqLOy71PaiqNPSFh6a0pBbntqYvOy5L3UInkBHsbaIYtw9UJw2hkNP
l9RtOd/N7FVG9ZyMRlCfnbrABeGuhyQwsL3xHUtHfs566ko8iq8nDY96hdmQ
6LIXO4K4t1Q6fy2KRF/LvyqyDmASO9mEsqJBrkRyCKAHzLKFR0ih35tl1dTH
35jaQV+GBAtjidOmScagebUbN9j1j9YT65K5BFXadbedgRpmHs0dcSwMp350
AiUxUSvg2GNRT2wJRUuLFBit3RUU3xG2a/mc2o6Egoss2TMjCTVAfZRRnjE9
6KOIvChFn9mTsgnfsgAM7M7Jp9/OeK/3NlJ2dCyCCReMOUA1Wxr183W5Qfl4
xRO7sb/YoU+Aajry2efZBwLJiiHPUJjIZ2CcFIfpAQyIVjduxTs8NSvWbBmh
kFOVGDqowI3DcGLib5GUMXGYCgISORxaCMn0eg06AQaq5Z01QixwO7RRFnlM
WcMhOx79ImYfXX/VRCm8VFwc80NvD9IIooeAn7cUNL699mJ+qtivmbEoIHH1
4CfHbN5Az+FOx7MeEYZq8i2MeUMVbACyvkzr3A+1rPqhlxN0R3KgRoRk4oUX
A2SQLGpthvytu7jwe9VI1W4rMOT//1hPwm33N0K3IXnWg5sah1e28pWYh4RZ
enjZl/aF5f5WUogy2tg/V1SOdSx0E0xbSPXfRx/3venJjK+Ra/3edxjIC9gi
Yokp96IR/4NtTmyfAIY1rcMvFKQqO7ZMp2VYFPsCxLfBfFq7VjJvFy0iT/9L
V2uK9pyDB8roKSKY1+oKB02j7h7HkbhW2AZOBumEE3M8jGUkjtIhul0YpZ7J
lCLfuKjcCQFBoq/4NhqDH7eyBW88IoeKR+ej13f3WgW77WKCaxx7sa2VoZOZ
OcVuDYBayyCHOLXvc86llbYOR9jkGLk4f0F9P05wXTVvs/ZoZCB1rhYN3OvN
2wTMVMaOaElbACO2sfkMkgDfHQFZlYOWU1Zts/V1P0BYAyLXTeacIJfy7q8h
lvf60V8drpQ+wrKB/m8bsW6YiPZRYxBrVbs/h+gzBKUsbe+AvV8EOTDQzowI
W5JQ+v1hVZRhRmrwVXjso9hNT3PBOo2P2kNWEAxD7UTtgGzbMeOnqgQXU+JP
Pdw4owCeyaisGedHYxDnRF5i80tQhWvnB7d6jVevyJWdi4eSavWHVk5yTG5D
/jW3NXrwAlyvDQlya9ZG6sdjG+GYt7/YtfbQWyQFGqEuqLdN8n7Hq88+fKaU
TWmrUkmpaP6rZ0TAFVx2QNy9qKRAmfew2jwl9RkfZz8rGSaUNpoErIWugSFe
R7/hLYNpBIZqL3JOKQIbEQtUWD67Pk8MguWlsbA79ldy3eQfLT38KDH13+Kr
wgirErp0TPsRlrfem0p4vtzVg4gtzbHDERD6o1t/XzdA9OWcrBjesrt9eadY
DumRgwg24FlmRxTSm5b7lrnmpJB4bvImp2ipL0yAhzW835lAkicmxxTgYRqZ
l68BrgHOZ8WQABOsnUo37VzJbpt6V25h9DOlinvjN48JP6ng2QWHybdx4ZAW
f2wxEDIAOSUegTpm+lVugpAAcgCxLbCWUoJbX6pDXkkmEXrey76zbq422Z6V
Vjl1t8FConRflWkHyLSYf6Tweo5Pj+h6mC9OYzVkD1osNZaV6ODUqynDaI70
00wDNJrkeThcYI3jwt00HWemZrzE2zY6ARfyEiua+d0ZXSaCvmKRgJaprkAg
8QoSAUJiP21xHT0T9lDGVOSZ4/Pa5QmA3K27cywiI3p1fmAcfsIZ86LfaGhu
5rAkCYKsWccDNu4DOmSI+adQb/TShQVRAATnfdzUZjbeU8lpBTx6AxjrBOlw
XSyc23DpOkuEHeiePsR7yC8Bf+rElscaOrpJ7rgxQzRLVFq2omXMLEMe+p8V
L4LKMF2TpW1QqTHOKSKFFKbDinWdtsJluzm5ntiYndXw21U9JXeEE/3+hLSP
+fSK/Cct/3EzlMsYQZ9UDG+HwiCl84HDfJP91LgRhIbkHKKOmlhnRIDBmNcm
OHl0R+lQ5ce0criHFujABEOz/4bvyXw+J9Y4bZe/SUelNZpK5XNMz5load+f
GyvztNXGe3qo+N6cS8QW9kl2aKLx1qwNbc0nPKoIYBXSgZbvKexsQ/8Z6xAp
/Rxq9wxlOQ1dbGkvi6gfjrRLMhCsWgOKjiEw8T2YoFvsWkIUoyM2YMH3fm+C
bKH3WZzXdTfZ0f68zermTh+uHirORZiChzYypQAezihvmt8W6YTUefgaSe4K
oHWv9V0RbUy316QiU3zSUE7IxkGgktZJRNyhqBQ4OSZqNHg+d6dvt0VPygbc
ZanqZGpZOG1kLcY+TKOnLCiYZrX2FtZNnpUNOFptYC4KKi942GuSw0m/nEnM
nAY3FVsFTas6WyRgBWFCkFZOabDmOX0cZUCeQX86LtynpMvapULTzR8uiGHz
Jnd7+AH95SB5inUA3hGqkFyDsSTn0QZjoMeQbKbcvb4WtJmslLwOM80g4jOe
OiWWDGKdYJ6xraHw2ZrHuBz2di2TpgpGrNNbkoDITNscd683T9aUIsj2OZSN
xDCCxzieRwWSFNJ7tR/Tf+Br1/uSDvLe2GsWrox2b76eNcgnQvq1ETIGCsvS
p7vK/nbpKCq3qKdVins1brxZOZL7eLn8Mu3d0QGP9ZW4R2twhEeiF/dIAsVn
M8N1COJG6Sm9U1IdDIw3zzWO/h/okIFkn6vBF1GrjF+UiTxUl1Y6UxcMbAzX
42BhgbdjKjGy1BgXBsWqy7Yv4jRteEia38wc2scTit+kwc+5yjEW8BKJxfku
kNLXKCRis0oyiBg4cFKCgqN61NdqWRqyVmnq3606DP6cMYB6aj3w49S28dYH
CDRN2qGX9kx60hfkkRUwJxHZTtJhMpj7++f5pnrUCzxKmMmxYazZofVTsxyY
azq9t2638H03BYuglG5bmFFdUFGqbrJsx2bFRIJnhk+7dSp23znaDfCq1KZg
4zcm3vksjW9exrFY1PCo2sRpUD18i3z5MwnQ4NsZGhdm0zoOOZZm9vvPJHd0
ZTxpkhVA31Dv6V9Z5uB1+MDwjk9sjAPAf5IATcEhMkujMABTNmCWtMgkAKrL
j0vmqAtpaQpj1JLTH+SJ9962fb4RFPV7WieRcrGSa4T/HtVlfO/UMCv8tnTl
G2bNiu8CIuSk6f+yJ/tmE6FkDQ0TGn/lHDdkflWpcY/dprG7/cHTHaWHtIom
69x3UECwWqffrTts4p94BoTdgMjR1f6no8BXIkIKo/oaCtNTzeglXIPmnyZY
+DTgGDYNEDZcfAKXrzZJIpT4RRmhP72eHt5yu7bbsmtdbGJQTRUogy2ODP3H
bOCuUAtJf8Xgd9uVpXDqABsjKKWV4LFe8sfZCYd7D4s8dLL99wq3j9D61jtg
qQRt8xYrueqRx55OTBldZa6MQXnWEqHxkn7xVC3Mg4NYUeXOtyy4oKo6lM3B
k4/cKVetoPuaPyjlw5EIROV/M8UlqWBt3qZPl1tc8W6L41+TVm0J3+kgXOoT
zoKgvDOlbHkMHKATpxQWNqzBjgwM+I4qC5ehlHglxClEc8IEMo1sD66J/uJS
XQYojTPxqkffVHeil8I1bATLX/JvtN3V+HMFV3SzpyL/j0DP3x1Y5N000WhX
34sRZgLbwyU9cfffvc8mR8Bv1u+HPlB2l/gIPb1AUPgN4gokwGF/UTWEW2zf
OcTFKgEu3ZBRleHBzdcBtr/TXCbjouYhlXOINiunu1qWSeJM4Ted6cpizLUi
RodUs4buK5tA4fEmzillZK0DPTZQ+iNGSfPgOfv1+2NLj4Erg4T9Hu8qaz4W
axXCpEhg/toCW4mbr7bwTDwlsjERshqSF9g9L4ltI/bDZ0Jw3lnnr3SgCrzc
3y7qwn8vf2cLQdl4UimI94Qo2JOWRvaT5CL14oMZcn6r/ZWvVbmvk1uH2zD3
nOVD505xVa+zfrP4JmqnE9K0rCwMe8it9m/BRziKxysDffQXHC2KsiQzaUPV
sqOUH3sAjns5hDb9zthQCxQlS3xdhdnAkge2X4IB5eLJaKXZ9pfZ3WlRkwsL
zAA0e/y+3eeT2o/5sWabIzaeWvDzbvLrvnZ7XlYPAwm4yplYOPD5vduXuJc1
bcTNHyVj3+J19Agr9zkxvLpTiD3YC8vT/XxgRgde6keiM/q0L6b65+AgmSrl
FBnFTdXTTLNVNgQSodMVLyAAteTt0UXPE9axU83SQ8jjme1qL+R2l9+LdLJ1
Q1iWPavskj7HMCskh0yo87KReYTg2R8jpvO89MVnawcLi0efLA+TsEXgQrnS
SgOEbNZRmXloxAaT0BYaaJZjtBu9Y+DzKip7/pVBml8TvCRczZMwfIcSmpjQ
7utv9h92ZxvQu9WM7zByTCFI9bWX1Y8LK1zCC9WN1sLNaW6o8Z69f4hRrRd9
hXnjiOfqTHg5rmMMl5N5evQUwuoxYTuqj4vsXNqyCY+XK6TvGPzpxIbqG6Tk
rBFfmBD4/ce+6dF110CQ2J2FV5oiAOTuK8TAeNR4VIwco6QQvgsZjWqA1tqz
1oYAM6ZzlBRoOUmbpPPZvkMimDYezFM3uHRfoj6PRE6o8y7YzQz8kLJ+Dpj+
4TXqj/IDG20UL+U0tFQfQpuAZnPND9UahTkiHTEgRa3oi/Vo9JrwEvKGWWZX
jV1t/gOFXjmoHWtA0QuvM728Iyk94WxyN7JjZMTfwcNV6/89x2n+PG0w6NPp
Ky+1WelxquBStyrd/lI8kStLG799LPVFk+GUetIJSnWvRjMuO3AwaV4hdXGR
7D+wcDrLoVJhdp3BcMLUosNx7hS8mvHouDvEm0AhN0JYXoh7sMrWbX6tEO4a
KbsK890Vzt2nY/yDZJ93OH7kPRaP0olFs9dbJz8qg8+cunLcvAep368PKEtW
v8UAA0n/PEfptI735viY6/KvTrKtVrH5Iw79BknSUNCtY18jor8oIUUNDFbr
hUwHs8M2birD7bOdA10IqR7r4nFO13lo5zkh0rnCu3mNjax9pG/EesgZOBlG
xR1gNhwKFZ63SqYT5Z01CpxER5aPQQVUdyUw9L8lgx0kqTQaGLWivrPB3ADj
quriSg+zN+Ei0AiiWHJVXyKwiYS40CL88MjtBQYlg2ZVfvoZTP81/s69f0NP
zR6N8CAF3kKuBxgxPceaveyfjdkszU4Ul/hCYpU9ovVul98cRW13GF7Mhhai
yoqSd/ysD9giTUoJbgSk7cfG8EjI6aeObFNwxbYwG0zPbuERRVc//1Y9uQCX
0pkvSaKkqYR1VWAgJ71qK/WT8oD7OkWApn9gq0hcC650Sr4JzqyYlEOGLYuw
UD24og8pCppkcPxWHS1cND3sxjTvRP0xMVT0Mojks4VuuMTYGnO/AU978uNQ
JySO5HWSYJPiDLQlmujX+boXGEgc2Qsy/O/1kni55NxOtRRvTTN70EyTeaPs
s+3b18mSOQd3ef1D7FqTtoqhAoplDzbalOzTwQYCgjYnjwFLEJl6c58LZeuy
7C4g4WEiOzfDFYgaR9TPA+U9JzHNOZpHB37rx/iBC0YIHTQe/XEZS0xHfVMZ
FxWVthAfy7OGHjUWceQ64rrQlruROMm54gWdPZXX7TTnf169dlM0dwLVVSym
AB6Qxass4EoNe5X40HsQrGedPVRIOHLQLeA6mdj0g1GzWjd7KuMxtYP4GZcA
4Q7xtXXHK525usZRjvKulrYZW26qL4kbmqwIFhYTiKF3YyEuk0QTBXT5AG3E
Q1pM5vEdDk1eOdsujY9UsNNlmwaX/2wGontnyOMbgD08bxVWkAeScSqgU51G
qHl6tt+mY7HaQCHcZyUhEkvswrZKzvP8ezN02e8WxtGZC/lkwsgazU1Evz1T
sXngbVrKcmtqPL7qMt//6Td4G4Kw9+uhMd3hFkNC1DLsmReFyU1nbcmG2GRJ
VUHw8xr/Rfrc4URWKvMQ0K9gD+osLYBnJ2v/M+inTlYMdCn2oD6tTVR8eFTA
HGMa6e0+F+iMzlj1kqZ30a8tjLqYXhT/q51wNR0oM1+5wazkaA8pFBxwGnFO
j2wqP+xhaeZzB6gwfetHetYl70yc/1Fe4yxDqUqesbwFRgdXsEmzKCbTiYJj
/6w2gqXyeO5H46Tx2gkUCMTSCb3CSyoY4zJ4LSiwfxCZh3Pe7CZbLdmJRRd8
ZaK2bdzYiIe0YYuEtbwp48N0C7MFFd8CbNFB+3qawLqs1bup0yvwEv+666G3
4TumyVsRc0b4SzAzoA9V5rJQ1dZ9upVrn7WafYvNuDnYw2aInJv3Cc/FmWaY
AZ1LkDJcrQUAT8btk+BUQthbCr2wZx3at44gt7BEcSo8aD44uhOvrmWo8UQi
ZL6hkiuCTuhfdm8uSk6xUKTUFBAEH3QqWpsNiCq2fpqg0bXObApT1bpWdMuV
AvYpbfqEcemLx48GsSUEVfp1OwhUj8J9jejlAHBWSbVBrY/DbFkYRsfTH4Nr
Il0h+PSUI0BLPWzIK5lB238+GAN/P87pKGHy2cxUhF69KmCeT+xcsJy8uY8d
WMPlAsv0W3r0FcCvZjtZQXTHiSxftZ7/wre2xYwuoCzkcpdt//zC4tWAMDdL
tuD2OmxtulgUWa/leTOVjYQWNfHKOujUEDNNcaZDL1bB5g4vLsUaSs74qmRl
OhdpzSllXhYvHVuvp6XUM2UayfRpbx3atEZvfBWJEHuvAea6cyCn6Knnt1us
OJmJnDHxOwygqB0VsYIcYlufiNAOO5wojhM0gCevjLU9NZ8fblhjfB9oJ90s
wfrO80SQaCIR1Vpo6TGluTxoq16JEaxxNmVnZmI/vhPiALoUkfkfMTcTlb5s
4nSj0rY451vEm8z8Chx1O3+zZkaw8tDkwouJFME9gUxLYlh9ZlTrIvWjhmrd
vvnYDuKvAPHq3sY74G59ojXrY6Z1zBiE+Xr15rGJ7U1bQxZE2ieyA7l8ir6/
8vA7wb9ng8Bg3zSWT0jP5k37wlH/2VEktG14yZWr65iIeNCopXHxm0xfXQyB
oUQRsVfglPy5D20V2JWMYpGFthNUcHhzUWcnFQq0khrKhm5+4hKG6SFtj8TM
YHwy8B50WPfVUG0OiYiEMzMMjQjdFB52NxtwP3FLCX+kFnrWZvlrsHPxeOau
aLDD3M9TzoqvSgpIgS0lFc2duQnNK3q+D8Q4nuCBVUF2RYHpCHc9WCLZnPyT
BIqZSPoQ3+inop1Iw+64qJOgQbuSKALak/WaOkX9VVf9669qQbG5L+Bk5HMP
Y+LlvO2rvtP9pg0a36uKVzW0iRzO5O+b4gBKB2rYCasu5/igYZ501RXsW+gI
ZsNOPamG1tIQEYt7hjZlwp/k1FgRjoujqF3BC9DPMzXTT4Cyjzr5eR92jo+K
K0TaNhWP2lvQBjvZTFoPfUQTcYAJOO7Ir/OvffQ6TmCiscPbgjzQKzXkTXRa
z8ZL0DFwaUNMtvTDowRXzZN5U4y5rLB7fQBRp9YsZwVt9XdgeKiWjoBdYwJA
do3XNR8mk/jI5TqFlhIpcPbRkKvHUPon7q+AM9KufknqLgcXHgZFv4EEKko/
ndveQJijiyUVUxvHUgzWiA/4wuyLWzonr3oNu9em6G6C6kspd9uWJogFK/h0
LOBHZQ6Z+GQ4BS6fJ8g4q2vj6kRedTS81ZI0qBZoaSym8+bEnH6Tbo5aqlVl
LU4WxY96qwgbBOh45Ibnq07fLNb7pThHDK8aCKcqzo2LXZp0jmRvMJ+mYKRC
XSoog1cGM+QgCrjriUi+Wvu0BUiwFj6mvDdzaFalla90XFxHYs6j6AL5RUi/
tU5F5Mj25jMVc1iBlpePQzaP2lqPnWLVk1rcox6PTcFAMuVkb+cj8du8Qc1Y
KrAfnB3Ju+EX8YHZEAwJTuWsfl+vAYwADmovxfeVu4pUSk/nY6X8aRpScL1B
JH6txSh+Xq7wzins3dMAKziSkz7Gu/oE88963Apj69d71fIjw7FZv2VNoyjS
Zw9j2szUh/KiwgsxpwhwSrEfk5MFSJfHQyp9gRy7aJwo8afQXz4rHg/p6nEZ
PT8x0Mh6ZEG8szaOqZrDP1fGIcBvSUL7WcdYjrPYY1GcsWgSmbjKDuFLWvGH
y7MfbnOvPRdXYpD8Lo24vzCtwzEBare2F4798CcdfZrnfcIlrT4X+HAZIahp
9DkVxiUBVome2VJIp4YD3iikDZRWS8ZYmVgiYr2z628eQ7rSyw6dops/OnoD
Xp1Hbht1QKY9EOWvKhVEAVPcskp1HIDYVhjsMellQTa2ug6q/Uv+6km9qui1
YO5opiCiP+YFQ9rhUAzqwfbbl+LrQA44dKnWzRr0ae8ziZpareL93jy0G8A6
6BVmH6d3jAzz5no2ZG9JsEBTy7hG3H65Z9DWLE4tjjE3CNH8JjzjTQ07ApIc
00KH/3oegZ1mQKeUwlIZkuPmqYlcVHoiTxzdfG4hGLHVp+WDWXHS1VU9ypAp
/X5RzR2Mrk9vIET/Knc2OE7isrlor1yQoeLT9T2MygUzoGIWHW4Em6RvwYHN
3S1RNiKumL6Fic2MDqFdOG3OGtuQZ78GwR+7KL3Mhh6vJUwgoerxpwQH76vQ
V++zr4Sc2YtcrikrIzXWshOdxczXujSJz/JD+CImV666QqxhN+LDy17lndBn
NH0TjAWziXE2aVTJtwbIp9gSmv4aEhkK8/19HUmJJINt3ru1awSi+gEj/rZP
DhVzeTbzHLw7X+Uf5ec+TqhixugcfN88IL+EM6rJxGLM9ARcehIjLX+CCHpZ
S4VLMmBzk1qSr4xI3af5PnKoqpB0/q0Yt26czVFOvb71K+w1Wm5mfp/IUoyj
0VOrQ7EN+f2kuRoXGEY1Kc3yt8hf7OkNemf3G7MyBUQKeQ9ST/vvWhP4keT0
XY+pSgf/06ILFPpWwgpkEpwoygEiuDg3Es1LARdC3Rh3iOAEJdLNjR2SgzUx
+E18KZzcYl6hxdcS+IlWnAvZd8yErhm/6MVF2Ou4PEJK4us822gN+uqIzDV9
WM/nBGHsZ43gmJXHfyWlEAhCBfmPjW5GPih+L2Ag+qYo6zdGdHM78Ej2fdwS
okzAi5mS5stjKi4NUogJ4pLLDX71IR1BrabVSHC2mz7OWIGL+/1xEAgea0VS
9pxdPQDbMwZImHAZZo01JV+tZWEqxpL6cfgLc93USZHX5nqfgAY7Yq6XA+CG
NFz8vGGdHp0Tj1O+MUOhW/LvlECpJdQsBtlBMUKSh9jMmYR09adGkc8EGMfy
SVSz7YhRp19O0qwHFRcX0ZCp5wNKbuwfuxgPXPrLiqL0onQC7C2TeNrKjVb8
5/AAjQSNNMx6pivZOsfQWe+lkDETOTCGODQh6qxVxM/B2Yh4rwLQbxZ0rQUx
Q0Md2wdZmVe+W7lHIMSmR2CuBb3GmpNijs965xdYgU4TAPrJlAw+CfKSLzhC
cag9lZt0qmRUlv3pTZBDDfRrGxgUdJs9LuuLi4YfejRQeBQlayUPqcgnGw0h
zDXCzM5LBbOXSTlgb2BBC5zCehZA8U0/x/1eQ15avA9pKdhYBjJ8tY4Z3tsA
S7dRRQNOHeuQZxrGzPpWuuh+elo3ZeKLovhUv0+hwQCo4KjCBnaeWCvpUAde
tUJBgauBCc/I7bqHQadMRRRVyhr/8McVzsbne45DvX3e+fIuIsh5n1x8oEBJ
BJV8/qp5/Cx62drjPALWHTzig9+Hwad29cSEW9uKpslUAnFZ8ax/kz7ar8sb
jjETqU3DidwF8+sZMaGjAYTXdkuB3hL4q40azapk/ibv9w8EJyob+WRZA7V6
AKWt8WYRqz5qJfToRZOMHBuphlXv1a0dq85X7WQXWz4bWKfOf9dJSrJJ7aVg
zV7eNWYwvL5tgCOF40chr9NEKH4ahwjJhOwL+xC/4GQ3L+gtJQNVO/CX4081
3n/0joCKWH/IJFA9lmDnq1XI68jSpRWfqFWIWFZjnoozEqk82EH/vKSUH5h2
pKGPu2NnbgdL16wY2K9T3aODYipqKoJg7tU+HxgCQkrm9lXBJVwreTHRtMWX
79qxBVapK1wrrBEcydqefmzeROUYl3nO8GPDO4oz9uIAUuLWIGKTbmIMT0JN
9Hxt89QLwIu0H+l/GVBGVYnXW6uFdZZjqsAl4j7Lrf1Bk4sgjM9eddhxb8LH
EiLbCltsQXMpSGxaqPlwtamObq7BSgnd27mQGwBc8hYkrVKJhsonBrRPAAA6
pGSqFDTg/TMPblxbdfM91j+CAugfuZrkmVksBeLbFU8vogGChzxNRsThhTme
DnqOeBWwQu3/zdZTjNdE2XQXlVY8L9kATMGbK0uwPFAHzTXbXjq609oshoJq
tZmEVBsXK07zwv43rmn07Ioahgvt6pZZslUbP1xQ5K0TVcoght4Gafg050/l
7+Ebj7iP19A0RAziuu6qiQKKLsFfo0hBk3RAaM6J/Uw9roygEfw0A3Dw//3x
KI1zoF3IauLRciu9btuAWC5TnLJkxkxuzdB2jSPk1AmLxHhUcaKHg3fXyGKU
YzpfoU3FqkKFxFpDxY6+bXfV6cwSLwDdms1jUgI904SJPzszHu0dad6yN/wJ
2QLZj6GNbeekzx1EaJi7mMGsXUdAytlqlMtXKYgB7B2/Vk/LnV/alewAovO9
3c53JAGnvd3YtHBKfl179Kq5KOBxFM8au6JBUY4Ko14NBDUufwIAS9yDySUF
jf1q+6cxlxkfH7EsO2II5NU6IGJnQP1s/sFzt2fmsWnr2glZ7Peyd8GPNuKd
83OqLkchag/GUY3AwxaE5foOqjtSgdTE2hMtw/TV0dZ+P9uWDjgCCAhMeI3P
jBKaLUVgb9Z9N8yacSsFF50kpEBDaf063HD+80MqbQCeiOSyQwNHsHz3A17G
AamX0oWtXOhoJQ7DbChXvwBWomFYFHPtLuqzpSr2oCv6mNvqV0OShiVW4WUK
sMvXv6nRe01grRGGmo5Ce5eKNqVMA/D74Asajowy+fmMNvH1sU6EXUjFuObR
eTUDsScoZ9Hp8Qlpp1mfyYR/BWyTMqDvLzQILI6L4DJnoqWx8GsZgxCkYADR
X9zjzAlxd7oaP5I+tUDoV/ZTeyqQ/RamehrsCA5vIOasDG7r4ZH0YVebIGpf
0oSyX0FKSvRDCBm5VnzuG7UF8BtrmMHcDOmpinbN05wkMAMDzJ7VQkF5srea
d99afw8lGAi+wEWHZie+n2QAAZySS5oyVvYB/+5gHuLeWukYWiarDIlloRwW
OLzUEe9L7xwtgaqo5oMUWuR3FXxD1kxa9Wystu1WjRIFK7rJ4CfutKGl6d+m
pdu4oQVyE3sGIXFm4yf2I0O6WI3BP8ydGVCfms7YrlGYwlh4MVndoNcV2kn4
KbX2kCSukMySuqm1iz0eSP1rUN7EbNtPRlnyQx70bYiRimxFLJ9uGssPwwUX
SWXpmDbWCvDJQF7bzfe+R63YW63Wh/j7YxbWmokqcTViSLGYWf+nFeyj4vVt
Qmw8P+xSczvIPsGPUIuKddBiqpNdH7YTu7ndPgtTxd6IGg+O+DhbrYc1IKcm
rOw/ONOwko3GfM/WKFYnkXSs3P/F3ZZclXMqoUL4Tgu4HaDMf/sYMimKeEF3
zyv2c+18Z3QERHFg2kSTlN1ENdRrrj75820ubOWWnYLkAoTjPnsIb/sHqisr
gM2x4QrUefAlhbzda1Mt0YaAMrPmNvHOw7Rz55MQgL4lA8ADsxTgoCoLcpZF
3kWJE0k7OVspJdXdc5uJ+p5NEMs6rHoV6fnMifkcmR0+6WEg+wtTYr4JvieB
aChSJW746VvHhqQP7iIhtzIqc2yqq5n5S5hfHqUdWJQT/+QCLd2EQ0JIA0Gr
odRH9JR5qBzXhINuCV2dNYbHlkhXXKGUTt6lFG7LUrVDPutB2rl6RzGGzgnt
DRQl92ty0c1mwBvHcIDYafAmRGWKjWEP6YEknvaCxDMVUYQ8breoICJkTMiU
T/MZCLBjugZLNcBHtUhMIj6FGeyBToir86l4fLP1rhvQgunHmsnfFZd8QSrw
d/AwohgH6kHK/7mBbcPJr3pTw6ega6n7rXwPEF+ThjkdzVmsZbs8qxPzRCRh
PejOcuRE1MY3MLoTQBKyvFO1Rz6Bxm54KDn84DwzIXZLZnAE20d4ZOgzlzDO
AuTgf76z/6bldOUwgXZlX5R9GjqGtj4TG4KPXNo74zRfJw61cmekP9j87rhS
RcqA1psoXJVsqFc6tDobLq3OhlPJLLjSrm1NpEGIodh3pbDfLzZ2VL3ItnMb
55sanWmLyIoXPdYl3AopPVrg/rM4XGoO16FfZ4sN9x/SGRjLCpO8+Xo+tO2q
dMzpdUuehaR02kNIvsvXFzgZLN0jIvfDLqYwMkRE/RV59OZ+NywMci2KuC5B
l9qU6Johj8S8TpBrZOvrZgCbL51/5MfzmiHb+WeJoBr5YkdEjEIx/+zZobob
o6VOooM9mn4pGiAM01K8B5TofB7vGJ4PB10x78kah+zH0HHLGO/h780yD5IW
MA7xSxhxNuAUp0C1nV5RUSeN0szHus6QRwP4Rbv1kBES5PigJA6p60/Lv6Fw
mzjGXoMMyftbFJTdbUMNy0R3CVosxlVTOiyQ+NROk2eT9jjZaXIyXuEwbhAH
9EDjdaYClNNbPivTLsZYBU8TKQ86GYhPPRIMZez7NAgNCNFvwzCvhAnPKdus
Z6XuRr40PJevMv4a4sGCNME0LeCuv00qnmNRcgmQ/YJFj+/nUfxeJrPohRpV
5L1vj4wZeAaa0UVcaQoG4VFdsy4oEz1JgL317XqdPlBELtWDgC4xco0rqRDB
3bgTb9NVHtxf3E1So90kZ2MJbzMluD+emuvKihax/dpls0FDZUY0OoLOOIh5
RvzzCbksmP6l78sGEh3NM6i8CF+8xXUb1KL1SFiluFDKy5MLfMYFHA7zr69p
hYekEcztaOAkFwg3Ee6+oOfqivZP2gR6hoL0HLEBTodysXGjhBUGO2zmsGAj
cG4OyVCWoKJNshCjNQ8Zdj5oGY7P8eKpKdiPjvncysIgeNn3GsU8m/ddWFDB
MEshNsbK4K8CiBirkLgtZkG4nzAisQaWc+gfa8i/YzIUSZ2y52y7dNS4nz39
kgcUUWZzN3x658NaMi4P1OaOW06RVQdbgbajyziD35SbUAWk2bx+VGdiVl7V
RvgEQP3kXxuwODzYylXHMVeMTuSnYQfwFd2F9Ec8k2EhkCQPAtne4gN88nKZ
fPDym2HucPmp/mTI835Tf5avqFYqlPJew9jc/5Q3+znDZi3tSGF0VeFUbuG8
Aqjq00YODJ5GiwXMFgnFdTu9TzGLyKamKwwvX/OUxiHKsx6KlgRj0s0shUIl
BM1sVWQXJw4y+dyWkGHK7N86iVoAE37aCkmmS9NUPYV95X7TFy4/nsbVGuoW
kHyjWQMJdoyuqEQBEhyU+1hrHQ4CBrxoOdBNpxbICKMWw2RQ4QMBgPaWN8+h
E7gWwooAGj0E2PRpH7Mriv6AXgSLARjlf2Q7TSPK64T2YrH23kjOsO4pyo0m
Guxk8Fji2YXM3CG99yJOOiWd1n76MjkuZQ8/dvawgl5N6z4+8b922Syc5rhs
c6H2f5xN0gIINyEGxtFabEJzuRKoClF4Oiu0d1zulWmtOGqYXs5HCREsnw6j
Pjf5NFWCSQFxNmgNK7ZaxRXiMcrjtpDSFbe8cur/xxCzkLRlcfEC7byh/Znd
G/l0CRSnTD9XgPcQZHeDHufE0lr35atbgtQjdqSTPIDJJALZoUDe8Fmx76BM
cEfu/0RqqUthzZDMLUl35yhWfYyNS4dCWL/0RiiMAJISFfF3DKslOThpbIfc
Wg0slgdnLRm3q+RY9VExT/eFPTHjtb4IhfCFkjVDMb2B87bBazAD2xfZdIjy
5hMYTs1CO9HL+/ix+RQ6X5av5stW3OmaMVE1xcQZJXcxvhKvCzPn3aLGfv95
TWBymXSMdh+HajHhew1Cpd0nFt8By2OwXAJ8/TdtI6WK/XenouSVE5YZxHEd
tCevwvs3y3BJMsTX9ULKG7VRL8sOM2ZBeXlAM4H3xksgahFAccPS2Im6TboZ
otc3256qaNSGh1dlz3pSShhGGqvs7DCw0wMtESlu4WbXMc+Fn8drRif9Gx/x
mV/xNOz+ySGM98oJBvVURv3MqYFnHpkBNWnucrDr6PZAyH5J/17vJahHeA7h
Sbm1Gun0itg+xfnkzRCxbWsWW9Ph316iS8uySRNGapPKkxW+Py+lfL79F5Ca
4Umbojj8MAnCRZDdxIuiqanGaOoFm7qkFEPqM4Ea7mbYO3iP0eiw8zpxTT6k
kNLFpFdKGK2Yxg4gQZikNSvDw7vfhDZu7p50ty04bbBS1GMIt59f3PooY0Jk
cTE+y9Vdt0o0B2OtQlaxUL3yfGcQNV2qRC6yWAlUtJVsW1EIcbjzh0ha2tp4
25rM/bjteY9wtbbGyfYJTOHS0RC16vsu2icD1dN4hJDDKcQklQWmo2x6I0B1
2Lyw8uMbQgpoZc5ChhoNPN1d3mCauNlXM8WLp+YRih7uQfO6w7UOv5mdK9Q4
VGbO1k+1b0yDVCYkozaUN00lagGNmt3Khu9ZhqCQeacV9+TnfNZIFxAqONLj
D8jll6iCB15SN4JAr7HBHgyFXzSQZxZxxxberEl//KrelLKenJRhLePgQ6wM
8xHflwYMuYvUkmA8VAKqHnhWKvv0vERLOnXx/zZS3324wMS+TwAsCDXMiki6
GlV/TgNo18SpGPDnHUrNdVIIrXC018qDiKuSDjFv59YQcP5b8NeVxeor7BQd
SOZFTViuDXcuM/5t6VRDeyiv02NWKfjt3DRkIVTE35GNX/hWIQjLlY0hPccC
16C20yaFiVpizHbZufHBctW0oJNfRiPYsedCqejOOo3DPpXoWRb9FlC//6/e
tAHOUaf5+gA6gBcXKddqcQ/jAw+X3ukm8mxtFM21WmNVuiCaoTpdjeYYI5gs
V/NzwW+f4kdWjKASxXvf7f1Y6YvgZFiqV4eSMpSTEkAOfBZWAWgDtSUVWtGv
bkP9SsX/LuiKLEGKOhTEVc7acxw8hlyD+8gTV5XuNdlnsc6wQeLLI0PmsH7v
Ts6dn2WrbAOFwgSCwu20Xi0mROkdQnM3jAZs9YtUTUQfUZY7SOe/ueIVkYE1
XGwpdXAZPguYZ+er5e4qT1T1hFjizlXZR3z0HfCUavVjCrpZNMXYBRg9XUA5
4i3pVrJFZ6RVcf/PD8yUXesc98ZT48LdOsDCss2rGVzQCM+hRn3sU+iEeOfN
OVZJDOs/EXyDkJhn7Ax/qEsUW0MJeCqBCDArkQfqxGjr3HEFmWWZJmmI6kVQ
CcTb1lg0aAaBLzY4bIgEQBBy6uALrhPSdkHGDmnWgCk9lTuBweA3RdjfgowM
29cFSpXrkSEiZmnfXd0g5wlgrEIgupLBQqoUZGZV+LGbcu+sq0iTlttfsZI5
4IB1e0grH8+vg3sppKPvtemMxv8MrksG7sNHys/om8bOsAOr8bENV/PqWauT
XFwzEPH7zk0BW+oAzzWydrP401vkeyl4ic4qOd4NtdFuv3eQYAfvUoQ6niTA
MN9K+36JBxd3ppa37e6Y1q5AcYNbGytbYIjGygJyN13sPn3rfgRA2ZskLSrR
TH4Nq+tj6T/SryhIehiT6TPIthRERemRMGBuzs/ajsQr50Qc7nnzpbCPiWAh
ZGP1+QJ7tQTiDJSnNL9eA7Cye+Uu8OwYI6d3OJlX/U5isrYUFodBRIHWuyIq
GZlUyBkcjEvfh/sc1WA0ZWhGgscSiPsrRzkVhMDWfW+RvBkGpS7q9UPGfyVX
LHqJiGq64dQfQsLDgSdaYLIwukiA9gVuIXVdNxXXkbcRTow3CKIlFXqtsyXI
I6Q2VsEmdIyru7W5BsGuOEeWr6eECn3REu2Ra+K/YyuVMDrhNj4NrgLZA5G+
i7zZDMxpYhX6PGVycgUb8H16AYVVZ+jV9jJCTcgFdx1hQY22zfk1jiC1uO4/
qK9ibwIopT2nOgLh+WbD0AABIGsxlXWWnd2AhZCkfVQrDkzfM5t0q28i/onU
0jSkqR4f56VSwJIR9RAZ49v3TLj3UlB7nQrbawQlq5xD7exRtptqxsggy2xs
gB3b00fd7tYNsS9YtfJFof8X7U4zkkVFttZKixysQGTnh1I4Uf/d2/uQ7o9w
QRFlpB/92GvCZ0yf0kS+ooLbpAze2PQCyz5TRGoBq+Q6/b+aPxdFCq5YlxDu
KH3CoAFwE/SfM+LpqXxhCYY+NDn3zya07xYyyodOhuOqvmNRs+ejL6kd3HzS
530W/Z7p8vQPBr81G5im7vjferl4/DzQCLllpDvVyZiCljP1O2s+vuMT4t/3
lotDIKgphZKrwZOuVmbvzDFJ7EFqFvHfgTC+gljxkkdQLYHaZjWzoCtVmvAH
nnQSuv34yhSoNyGKKsdOtU7xe9AupkXvAS00afxYTHj9aNk9eS3z76I6SFx5
VJHHVo7CLd6JoPCXDPp5skWtzFwmUOt95MoLvqgU2bfUCAR2Tv1PiL2/8vBr
0AMYzq0Yfq96LNTycQSCb95oxLOPqmhZs0OelLa8CByyaWYW+6bmajq6lo3F
+qiw1FsmkTysUVqlujjVr0z+gcYcsqSc11vFeylGPetfnOevOp0Y6lVBm/16
sbk1L9f5ToixtUupXmA2wugD1mDYmea/3I3NRqL+c1+Q3pSX18BdZ/ubXCR0
bryjt0YS/mW9p+4Gy+goP6jHX1F9GDSbLYxaOKfifqFOAQMmt8syYMkZ+h+c
jml93MJfX8kij41o4rJqAHyKzl+QhBs978SeMIezDJMcNOClrAKrUF8ixplj
tIGuvjPBKcRBgvjTpFTxYFb3tWWM0UmZ1vRw0Cbtrh1gD7ZhDaHaCMvdHN+l
4HbRC242Oqo1dst8ty6jwAEfr1OphMuB7j45fhJSrfNDVa/pZ0nbPvZ24PY9
B/J5ZLh6HQSUCzxDx2XR84aAMYTuXtPL82icMJf+ooCzVPvtfQF3WNw6esOy
hhnmuK4pnB7JkA5XlkUvUMtCpgkh6BN6a+8gJDoM9JwMfqsJSCCSSp8YvAQa
TuMH5ENPYm2KyBKzBJNG4TmeWLTDY8vLRfSix4C3ZLr+rpBkPA3WPUdbg0qY
VmpQtciMwcLfGEv8qlzlYEyxZq9SbS1L6bO/XzzC69WqXSjb+rlLIIbj/LHh
Nzgjj9RdHlJoMgG2Iz6zHGc/5gw1YOgzbtOgEvb7RiHiAOYfoblQQbKF5uCT
QTglSm7/mKY4PRVyR/02/aKt7Tztyj/UdX0FPmPUe4H5eLy4istRsLg1t1dE
rw5Im1k2i5isUGEQWJpo8VZHabsXsROxC9FBP0kvVT5SX44Jyk/cnWm4WJqk
piADT42Dbuhat4dFGx2pdz6mhl3c1YWyaCo/BAZY3sSt0C3i3PxVzJPWgnOG
MX44aKI9RsaGZetNCoFKnL5OLdGQR7T7LCM/9CzKLAA2PJTRjTpqE3XNKGcd
+mKEaSGhG9gql/UnQgRcJFSbXzTFdIvUm3mJY6/VUJ06O0wyzkeRoLLdeZDv
QNy5k+y1mBaQaDeuxYlBZD0/Ih74ejox0eNqWb7gbS+OohrhJvBHJFSDmpt3
EVMr6Gu5lPQLm7O7a1rOwYTV84P8jvIOcSSjA1AWfnJ7kLQQO77NycrnEHVK
EtUvmlkKRCflRi/SORxBJrCwUPUvrd0w40/q5iXxqBFZqp4vpwFV/H3Q0XWH
n0ncER6uzl1DcJd23townZcrPZKYFFBrhvhpNMz5R6QHmuUSeJdtUa8piidR
iq57hZ0+lEczyqC3VjxMbKR5HxCKHed7jDynncQLwopTh0vXL8WtDN3SAEP1
PwtPP20Pfghgu9cBZrMF/b/k98wW8lv35GnDYz58IxBSh8H1IpKrXOp2fjye
Oas7riiyzEuTcaGc651p8ihp8zxlYlRH93/cZl95t2yU/RtJw+F3OXxc0092
VR2tg6EWWZeXX4/3Z+OXOFKqBRSA84NEV0ygkzF1HZUeSeOF5HQy9ARVargs
EvZpdZ00u5iea1ptZv3lFCSWlYQiCax59esaiQ22xi2gKIUh7dRc0q3n/KRw
pXDoOdT+7v+u5RW4LL3RR3tUuFCBL+O/A57Ttof8GWD4Qaa/Jrs3oFBEVwM+
3ng5Wp56hFVixBjEJRFxOMHwR8PxQ0qaLwGtIpovh4WQt/dPEJ8390OWRQHp
1r7RxbikL2YdDZpgvEuLinytb0Uu7k3ovdFrfrmMu6Pte8sH2VhmqYFsW0Ff
l8rSV4MZvePndSvxk9gfFSqlyAS/9ocLd1tcKdlF5sltRjbhkDIHOSJzJNpY
llC5ljqRmZi7R3R8z/ehMjCZXKw3XzCQsdltrANg4TiirfA0HBb6Qyi8P/s+
NsaLxmFWMBm7MaRYJea7vhySVmSKuToGR8hPQcDoy+C67/X3+JifimeKtDOf
uXFGRz7cuJtepuTnP0Ms4kz0iFw+RulGy3wWBYdiieCPVAsatVNk/qU0IMJL
IhvbLFYak8ZHec6ObLYxXhjyXPBBr+t7eADbQUjmzXq5/kfB1wNXXyNoHb0L
6ci5l5MyVWwItci+rnPldeQ0NvIJKFv7v4aBn7BH5ClHD/WU3CKOKbdMg3HI
FLWVpsXyz/AUHQM9Dz0kfT3K5W62cYejEjqP4A1oiwxEcuKvJpOKF8IvH5By
PT8WEra4aHK7sz7wN2j4x6UAVN7g5clEpncY+am0lzqmYLlKKfiErk4oZ1tN
RXAq1mNkCicZcTEBnaaHTfOyeiM6karzzS+HnsPHjscCIZIvPCWn835mMAq1
nMZakJHCSuoVytYQ9ucmuizouZGHD4nDzFQXc102OqlyqnQZXpUdbmdziSIV
MjQS2D7xmHMoYp7LBHX0Ib9ZGDCM8Eb8hWZRrdXnq4LvbMf2bUnPwl8OMghV
HpN33/lXq1OL2Ripnr6CtTnHVeSQrVqM3gpe/UvznncgckegxqUsEmJ0Dk8Z
1gqzOLzax96scwUwfLxVHUar4chRWaQpms6cihOscq7lbw8P4WqBYFANA2i/
YrH9ZrKYZBgxQ8O22X5+PHST0YI9YU40HJ9i3mfdIj9FQ6TPZBFYcdLGaCJP
gSbz0yPN/Lec+fV+IhfbSx5nRFN7RXAMPIe0Tz9pQ0dlbXEVGG91+A4EjyZ6
rZoH65tltMPyM/V7O78M7ACjsko1JdCOZjZQ5Btrz5UUsRRqzIr5O1FNqwPS
6PNljphrsjBcffH/DgZjB8E6aGAbYgtZVjgNnbe2F3+ULlyeyibbKFn623pI
DIH+u3f/IgTnmIaRFG4qQMYnvq+I+O9wOrsZWjNAm6D6Jqq1WIQbNBqyYBWe
7BwXGsicR6l7mxtWktFG6R9e+j1jmh58DnsU+wbSZRe5y1gYoGk64i93IQS7
5q/kffbB1mZzcaTm20W7IrWlh/RdujTtkhR/mWrjE1BvE2/U6da5QGPLaqN5
zGpQLMsqkNji/o4zyHGRit75IZTmue4DqSX/kmnxuzUr+kEyGu5Vcppm7i0S
b3zMkoa55Ace0T9fNlKm+tHQdxi244Br1C0vKsYWJWd204Wf+qhqWZa8mu9d
eNkptFhrk+Js2uPOPOOGmRwkxkkCmPAa6LNcm1iP/zUPjhZHOq2jx+wBxdo8
6im0PKzDdlR5OzEAwmfTR8S1s74X+DbrzBeuh9MhXj1l5PCk927fTO8bQVMG
gmJubJh5vra6WKgs4KNIkt1VtfsuwfK8sBW3PhhgvbwX1hLIgj5AI49nOzVn
VxdD3iMQC6DWHCP3kkpoEE5F57+aHSiHzZu66bR50cLzyJYmGh/d8X5D9FYC
H9pzL0zhnXCP6UmSFU7W0VQtSdicObmJi4uAryJjX+mR8ehvbh45v2YXFquW
LefCdHsUBMhm5+rwitcap1QsrzVgC2K1Mac3CInVsIhg0fPzrhn9wsdwxbYm
qt5cixDRA7r1StNG9vJIt5aEaIl/LDN1LhwrK9YBHScnPLv1wdNvcIDLO7JG
eZhTTqwj4j0hf/x595BpbrFqmzLIoM6Le6hkA63uA4Ql1euJqwfGvAhtiueO
cFxEOIuDZn68ksml7wYVQjNT3PXbh7UJxT1MkElpFBUNcf6XuKgBiQPx8Dm3
7lj3GZNU/DBnLedEXi7uSgyidPD4eMjjHJbVmbE7daVaN361SNiY2izGLMsY
KnwIqIYGrJmz+/4aZ0vN/QGfG88H4K20pSv0o+1eyaRiYWzE3H2fWwW/mLa4
ji+CR1E/7A8KTXvu4AHgrUftE3qXTV9loK6NjeKOdPM3Yetf+4aLnmanOsSb
5Bd9OPWIKdPo2ZfjDQ55OFI1QdiIQkGpoi2Kz8tHdhZefv0u9mP+xN+3/SPv
R+xBtfsnp0Djg8Kw7TbDZ+765VMoEss/ccvvDrWAtrzPwz8erHCzR4sovSM7
foxMK/qUmNa3p/9qI1DY1OyPh5v/7xriNjUC/neKeg3fzkBZH9O0jfAsYZiC
wUYZo6Om/ahdRtITMJuMZfppTmXKteIEfKJ7fjcIdHoMDxhenvuekvJ70YCN
VuCcP5/7frCxKmKcSB4N3YQTWQgVeq6KZHf9YGEJdci+9hx80drgFqZ02kOZ
+zawS+G6K6Qpu0NINY2VGexaMoYxQlzYHGrHCy4a9P1vJYoW+2CDnYaiIy+/
2Wlctj6krcD+QGjckDYcqfIyjL2dxnUcT0inkbqJJVdUEA5mB8p44O2qQFBw
N9TLJIYqR3X5dZare9oHBUee3Wm3+qfdUFhTo3PeCZltg4daEkYyHaTnWgYW
xKq69cnBpeXWme6Y/sjGwJ3xPCxmjPLXuu6MlTklJ/ZLHkOlWPIF3AadAK/O
kXu99TG5/gYC5HgG8m/8LmiBcFBawUeT4Hs0tgLk6ObsQ/8gKynAxd7z/sA2
WADY8MbNpCo773/rXMk2Tk9x9tBaCYidFtiyfg0Z52aQvEU8pBNSXzaVPUJ3
BbTDVQfTTbfcvG5bob+w5KUdTgjBI7mgxx4tHP/ks/DFRzLrF5UO/gWyAmYV
ihP/aKbh+809ym9g/xMjTbesTDj9eokhVjpEE5cYEk2pKm+IjUX52lbqPoW/
ZPk1TrywuAaNvUCbF0QXS1qqTAYEQzTRYWqqNMiszXQc8zhzXtcyahERXkcD
7ozxyVrzXf6MSDBLXGoOT4RDzO1is0MvjsnFz8gRXMJF5CVZ7J+LQnf7MLrF
nTgqjYvAdja0GU21e2jXbizBK5gCw4C/fug9hYPQ3d1cUIb+Q3txrNEPVOPA
GjdpId4PRERKczXhbCMif+614dGLJRYycjZ7IuenJl7R2G2THJQOKHmJBJaq
qr2xMtZWLut1mpV3QxVl5ujwsiaK/wIekGNJsOD0J012zR93RtK5sqhJYXUa
APqudXxL+t7Pw0+vgSaarwLAmpqvCtSfSID+MRhtiRz+d4eEq4D2kmRUDYPI
lvLXtVbZw5iuFH7Z2de/O4pMCxSpc/zq7SLpNQ1c1XYuajVW/IVHzFpIzyxQ
T6khiwNMfDcysmmsBgP9vtegrOTL1OBhBtkSUdWMexBoLLwLZ2gYQGN41NfM
+Ga+KSfc+kgbmypg1KlAI+MG2DACcASdbHrYxb8vLHvD5duGHUK8BCmtyoG2
n/mfERF1g0MtDwZUtK0sHDfWr5ob+EEOIbgnQVebutvDYYvYR1UuoQVicP3o
GlojelWcGvN+e2eTtY+z2y6oXL6xvVLIBdQYAcI0AGu7M7boWw/yoaj1PGKh
pncWggwHR+JCptJEmXGqWC97L/qLqfTB1bw+UIdRWlzIHIFCibp+dxVq4o/Y
coYtPWtaRABe308n+RjqNchirQh0Fd8zT11ZLnft7tuN9UHonNwBqhsuiHTc
KS5k0wZr1wX41H4s+b3+qQqVWKNEcGozxAbGLHZ+JJpILmJAKymhlebm6dUb
PDBB2nb7waVgy1wgALWXYirGWc7BT9q7DBlPOVLDWuqWIf105GLY1SybF451
7sIr9G6OCHo6qyjto3yKmprA/OcStRkdKp0qsHLkFzbNjQo8AD3DcYibb5fc
7ADXvlzD9D+93ObxlFqmJmahGfBxISUVZQVwacC70NDRP2AlG/fdHCx9pmDC
lse4tHnh8bW4t8DIN7D5WAcoGsUWFjlW0jzCupG7dXxLlNCflxtsymkkOTST
8q4p2OUR2FkAYR3x5oNCWtYzEgph4uXZoEs96GRl4sLa9boLlHQpRdfWHJdj
eGHV/oZywn7gjnuz6mvkGmMTP9R/++g3Jgl6FSiTt5St3a6FQr/rr9HOcy+9
lPjyj2YOMHdP/CmGkX4i08cA9w3Wu1IKXrxFbUv6ECYoaUI5XrK/7JpINJRh
LrzvPisREGvhtDSs/6/rPSLFL6UVTCp18T4eEPxsJvOsfljrH7T+ug0rz5/F
4FizWbiJGGSO1/Bf1uhM5aNnfolHqwBSPyMJZLSIyzsCHA0t4KxoQ80JW4iL
i5CzDYwshgQynIEW8lYqv/TJId5gAe2xHiQY44V8OrvsViYjtCVmdDsSeHJH
cWHDbSE75aFp36Bho7xPF1RZQaecbg6nUTWwBFudHmGB7RN1NcSkRQ7aK6pU
UpJDaWbAqKBe/0uYeMEk6IRi843SOaUJRNJx/jYHp7J3z8hWQJfiIdb2XDpU
iYEpitdoFlOvRd+zhBXqaL6YiWcWsnB52SDbftskClsqqTM8Yl4OI9xAjb5o
SiGlyvGKbnWY4SJDuWOyWENhw9Aho3LGTfKTEFDfYBU7KY3XuSKLp095rTmI
qbGSNDjqnXxx2jpwf8FTF2dVrr7gpGHqJ7p33KsKXMvKYG/ZR2hJgJvlpnzv
tGbrWV5oub5QBBrDBmuZDrGbFzcqra8v9I+KsOfdtgOkKbcgLmcpz78jGzTk
f+mlZJr4/oQioUVg3R5MHrzq29ejI+TNOJJ2PGKhV6E0TcNy2wy2TcY+TmXC
r9b2sMu6/lkynPsZGn6GthdzIXDZLp236A4QdaPAwohpnRmswzCOwCpavmX2
UcmoGB/3/G9Vh8K/nqNsvRyP8AUpAkj3M93Lkk2qfkL8b9NUJrZyMHhLpMIQ
ceZGO85MEG4a6t59h+6nE8Dza3tVItvReHDz2L+IXHiEjxKwDyGuZpX1ki0f
3YYVahajxvXOOWc5YzwPLfAwRdM5kgj6pfJlnJTLjkEQtWcOqEnmVgTKqczO
euGD5UdM0LgtaV/UYHyUcniu4VRAJbi0BEtrYPwA0Fv/kCh++fCZu3Lg9gXX
t3SxCdOKaRull4ZRvQSgKIrtQ+auij796KLTkHGBWE7yy2gdL11HXGktVvpi
/etGQGAMHPZL4Q0QLkyXDSga1geCPiM8e6s88PG5cdbV5sc2F7dSQdleG7vl
3aLsEWyf+rSFg7fwcDhgpeJQriQh9Qvxa0GqG4qCpJsM/8OheQL/Ygf/tjoL
yAhuIw2cugB0JW53RRSMvUHslRNczcvV6b5uXW6/CPgqli1jLAIhAa+7Gyzq
FC5tCCsHENMaydYWtZVnlHdrN7Q2XKKZ3336GNnAv4YV2cqIf0OsCodcoYOc
aamz7F2MbW07hU5NdE4DurC1sDzPmRxLK7VW7O/A/22bP8Tot4Iog7BqlIbV
nxsQSQ7eLQNOLMyLN+FKziqBbzgO5xlMYuZVqlgwvUV6hSscfPbP0pVLPI7W
TZmh4F8c4oUCu97seda+iP9tKQAytBF56owOsK8qAIh+D0QLigOEYDrAM/qS
2FfeWpCTyA1v9JU2cFT9p7WlSTOT2lBDf/Sg8jbP09Kp9epknsBXEaOaoaF8
PG6e7oYJRRJY83HXV5usgckfZEFe0vD7bEB7WimnpTbU+RDprNPD0MLJJguY
kpWxbDWg3mMAAWNO53IG88w9VjAt9V+sokMRNWuClJxJ3/x3WxfgQ2p2/Vsn
uGKMDD/2SMSIIiGzz5/FiOW/9O7a39X585+0pBddLFEP4JaNuMkP6x2rlubq
0/DDUNZm05WQDjqGxlKQgLLCo+QDVV9FrPFOG4WIf9Zix/kzc2Z0DLPUJaDG
XL/CyJ5JZk3SJxlk5pCjMfiAKSwwNNhehdK/5hSH75UeVvpsglePwsJLirpG
+TxhnbLt3Mwfaa4t09SHY1yAUelkY2MSymBD5PlI4slq6QhY5RvhnFkMHt4P
bGGh+wksOXpm1chZiGSogwkWFPzPdzc2zzBta+3DyWEc3B3ueWyjmAw21TJ1
2XTv4Eej6eBy0MdGxjpNoDY+UvbLVem3PjKpLqMfLapeODwZa1WUFwN0ItWU
CG+7vu5YqKneZAJIDNnZ32QvpORpPInqQlIh9DB6+BqXNKgzOx0DoFnLV+k4
a/JoSJpFE9ldoZS3dRww1tvMzIvAw0sEjUVCU6tmsu3/WPT5cTswlu1qFEAV
mF5Y1t9b20N1D8i3L/RYby7bKniJTcfwqQ3du7nkbDoslL9w2MjgwYUrPGgf
9F8I1J+6MgJNTpcEYa6U/BY3tycgH80U9TUcausmXzCg4JkQfq1B8e4+biU1
BAwoBft1Te/I3EF8lx+yWWEj1doRGWAe8fNGw4QO7Lefpt66O0MjUgV4ZEGK
fL7Jw6K5F+2h0GzOtD4A8X+ZsmfiIY6PLP6WgViwRPppPpHpwMFoUcX/ZJm5
sJTCO0QScIvrHTst4pNdjI+7OVtfYVwst27yPvhW3w8zUsxQ10LkYqB4wCew
HdIPvrhgrTvb3BohIRLR/jotqLDOYDcjpS5bsv6iE3pc8dO1GFN31n58I49p
6ls86rspEcDU9mmVuCZEbsmXacCmyZiTi2AymF22X+jvCyv7391LifXIsDcz
H+neXmklZBpb6RGHp4re/9ZKsNmv/Df1z3Qp2upOtUe7H54/OKkRK7NErpZY
o35FKl9FwW6Nubyz36hGQk/V0lAD0uL9+4LRpI09WUuC/qHdagb1WnEcJPJt
wfNOLG8NbmmWEGWMsLtK1Pr0BliRYLXZpK00HXFMp00+Bh26mKtV0pUJiGYD
+PJfFI8GaedUW1LOok4jR7kKxJobnFKk5prTTC1gMPVlGi3iTEnvfuiYNYil
Kc46/eZmy49oth/Da74flNKIbU1TYajLuWomp1Zv7T+zNkKYXImtEihuGUQb
4PdFOV3Mjb2yTrwc17Z1i02JbE9IjAtfNxTrdU57Cxc094B85G8WcIpf9JwM
idijIvnadAApgCDZC24CQknZRSq8R5AfOPvkF1sRbpPruvmSV2spGlHgJsqg
LsxFC8bg99KP5XU3jp/5gQ+G1y+Ni0XXYXBS0unDKCFUzhpkAIdDkou6eL3Y
NqBGHX44cYXTxK4m5Dzuq3yrBbticoS3NaN5yF11962O7HNIN4cCoNBk4NkN
eRvqtXz5Za1p0+O+q02xhEP5RkCxYH490V7keUtwPLoBWJaEFmBuf9jOY1RM
rSy9CARnpZGbBYCON7Rabhh3VraGLwPYxOsZ97M17YXXiz2ufK5A8YgDtuhi
lf0XlTMN/gHgOG+SU4KmIUiZbUVtp5BKv3/Z2TcmbE0x58k/JkwgGqusJbAP
RbP374EO5s5zO5tQWy4PW/wHT4Evre0aZuINA+57vIrvEay4il0qb2btC84I
6MPPI2190Nd9REPjuawPNIPaCeAww55Pdb9LrSueRX1HAbj4Wxuh15PQn3AX
JGU7eiv24d1GkVPEEQyIumOku2fGxaE0I1jGKXxZRbKiGGJr159yXbUHPR/z
wMCzoZX/ke2SlgNOyuLdsJTMu6ZfuNcxCIYS9MG0jjNM9HnggNUe+80GZKCj
DsYC+yP6+QTzd0h7kFYbCnhjobeLHplU7iv+YFwQzX/UMxD7Cz/gBa1baFMg
ESENEokHFTuyw0y/OOpbijiw+dvBn8vo9VFZhWntE0G8JISO/UOZ+RaaX23u
G7TssLUgjYH5i5x4wb2RIE2adpKsJQnAcJj0kzccskvyHvWBMMgTpl9xy43j
0sHFj8OG79o7QWWoBVUzWbBk37p9PMPDPwQ7Yv8LL2HJuBdy3XTi2Rylodzj
uJaLrc0XXfflHuRWUI4ouNlcCoRlRJuLsxpTHuDdOMK25rXA9B4pZ9/JBTaF
di5uvYaOMiE1aKwPl37ZykL8rm+kvC1N5977co7qigBmVw1gwzUml8zCaDTv
uAOje4qK/gXXhdRhGYyiBC36ykqHjQi5xxH7XEKvM/55uVKcX/wYSyTkm3EG
ThGv8a1LqQl2URYcRnycouQd5MTxNAcPIK6IP8VkdMEdBiFx8UxMb5jyjBmL
HTkOYfcCTVgUC6WKGNEy6AyqVuFvj6ZbKFXgySOtkD2vVomNh3wuz6BOIlaf
yIct0DHJjXMfwIbZ/eZG9JKJ1bnDQMOwpqQm8kBZNrHIFb8PZEv558xBIGLN
Gw6SFVVmF9naB9oRMu21sqkeserWIiM9Y8DpX2L7eh7GIk6MwM2o5tX2179q
hGWEql6VyINxiHsXgyVF0wcOb996OJF/mQhsesdZ7FUnfxLEUXoNwoj+iG4I
5B9sOeQcsu6X0hOA3yp8rVR9ekobl6d72/5bIFByNvXgk/Ej0Pm+DYajlalA
iiiVgqyggO7ZgM7mJ02EyvuTNRdpp3zhrFwsWY6q+gw5mKFT5IYhEC10DwWe
Ppvwe6JQJNDgXcPYBnj9j4BL+EEsy+Of6KgXbbI6nOGs/SVS6SHO1HWC8jFv
0Oo5J1jqycDoDeBdMr6CcIpmplMAHkMA5D+Z4mWOBF04Pvp8d7kmh74/3s0p
yKaOXYi8nWHTHQcB1EyAo9td4vDZB7ljLNjG6hIlnoHh3i8Ktyi88rfvf2eJ
S06I67v2g79PSZMKVLMThwtbVM/j2dZk7QJmKraC5lGrJnwLDTQplXFf64F7
FOViIex8yf8V0aR0iiX7/CPU/33JVN+ne9xNT5xFQOMDjA3jqPKZgwHhfcxf
2QBSc2vPZEFtRCW1re2ruX0Xntz/qB3pXCXWBAyChtHW7pkGRvKFkn+8FQNU
T73P3d/UXKZb1E6QEarh48s1KCM7M97KLxFb5z//yQwcTqMoMoFycApGB571
nRDJZq3tsVJXhgvaiDtdYnDD56WFq1oR7rojAJ2ZTaBPW4UnmKZnAxKCvD8F
FinMTK9d0RVNHA1DV4OWH1adE485AA9BsOntKfq/HV3lgeyIPJbMWMRDAB0W
uPPrMsqr6cNaDaQxWKPZuwfs0zq/kap2p+TO4EtalQkbcJMVquDH6zO/PvKQ
fiTGvhxOMcUcUv3eeTgNWOIYRkWPWHaRxnsZwZTgpzPVKRLyiG/rp77QM0Dy
iPGpiwAoBbeHRAGv+qu8i2iBOsXttAeFGNDO1pTqWBYYun1oXscNIwnkoQDm
1I9n+0Pnox1UzvMjs/uj1P5GsDL3Tb9V4NzqwUSrJgNjr3PnI+A+HKDfNaH1
ZifIi30jcorJu5Jf8WucLrNVJv5zAPxBpmoeBP0vnxKfIq07mWk/4EOOMeFg
ngIyuXW+Y16bNVnGSAHu3y8YZO3mTYJknM/JPBUWkQxv/oc+WKzB2eWBp1oq
Ed49xhei3aWXXgn29CCNDYgITQ10mUlfz13/izzHeb9reKUUUUeoVxKYpnIV
SXIOVhxIAozlhi5hmheIvy/PmJa70Ml9VVVNilwPkUhIrbYq9w7DHTSqCjMH
DfH+NY48vCxY8nlu15kmKlELR/QNxMoo6DDwPEaARBY46d6BS4N28CV1KYTZ
qJpxGVQuwso/kyepdlAl2je4VZhcejsIYbz3gsvj2WFKy1hEUbbPUFlV+XjH
xvruNJklqDV+HpMm7u/ioAWa1Q60O6vNJrk9M3R5CJXEkP40lEJhf/3etYcF
CTCSrFP51sE4El2ztvFSt/dNLepkY9WaLIcQxr07xXS7GusSJAlZSNmpwOzS
jbfZN534o1tCetROwo3dkwnboJeKTto3kwvU5ENPogVtKJwpc4Bc1F6nHNu/
x0iNgbm5JETcwDOe8yzdIVbb/fQVdVYHMyLRCTtZwo+5Fry3KdQJxZOZfQSY
jm2RH6v15EiZs3Z+end8s905YA0ijs+xi8y9VPF6d/2Z9Q7v9BDrBKQh006+
jEisbf82rqNw3i3jgOlyQ9ZT+ox5b8PdfC0JVyIQ0+N7a5c1y9Xs6XQkk4hP
j7cbeQ03Lo5wWop2dYvlPG4O42TCxALYa76YjjxUYSuTmbwmjC1srwNNlmDy
VKIsF404j5njQ2/j2CUWNqjyjgyWGSmZjf117ahkDUIXaEMNcMKLGY5gv5s8
6NfTWIzn99nPROcr18Fdcj03rs3rXDp2EI+rMTmDwS6128ZsrsZ10/YQQlfY
Nd0vK+5igwwdjSqzElqBg4j0zetqJdK5ySIkpwRDShqf60PYGHVTHu9erom7
LcmabdmYsVJvWLU2Sx4l2FXAwjIz/KWkHmsGOiBiSbuxgrsr6A8T4/3uPWiQ
h4WhXTmUaqO8htvQ4caZMiuR41Ai7Y5p0S7p+k+flt80rhW7xPLVMYJ4smcU
FV3WlPnclm9GC9kFX3dzpzjV7pN4a2Oi8skm4Nf97qEWZ3pNihIkBz8GTSsE
+SeWVS+4jkBqdr3mERz+zCO/lXgtX1z6uMGnNXy1G9PyYwNzyImREkkZ1h8S
q8DNtVE4dmvZ7g0cmE+WxPMOOAGY66umxA32AlkeCCnZwBtdkuBx3Yqrdvxg
sN/REQ2Tv2yLYwyncZ142uqzRq8hjG/bNYceJdXGk+qa1ckKeq18AuaxHsmX
FGnRD7BI48ln+s69kp5DRzWQR/QnDrp92lj9DwGMlOGV7AWyLxxSATkF9kYG
Co1rr9mJghJoHgLHm71CJ9B6KdGJNwbD8IjatlZ/6AVdiszSxzSYxsT/7yTn
51BVTtSm4QMlmMYL0AywtQAtnzZf6zHy5Mvv/MhEr44D9NYNKRfzwbw7pNA6
6x6wt5Ouzzj2Zn3IHUR6DhvQc7M2jITOc0r2k9hJuGTCRNTbubRxLv51YuSG
DDGk+CJnj62U7e2GJywIEMfilAgP487G44LnCx4ebbd90sPgN9a1mGcI7I/J
hBCkV69LYiYjo9OYl+ptipWOwqLVcDULPgM+5Af/EnYTa5zVhZdp9xEWbNxW
hif/XHlNJan9YCVv/VeusH7HALNqPXYeiIATmIXCDsXH5LauyCsGe0chRnA9
0AgYs54JdxsZ2Lf0AMLatvOg3iNanxA/hh0LDuK6/PItzdK5uhwz7gUQ2aQX
J3lElnos9tD6VGp9SuDPMcV/2Hx4xJ33VnZ4DGx+UJle675fw5QI051ekr0j
Gviuf/SFY8FrJpmw6uy/ZgatzCvx5xSxv3U3jEFjkNZYA0zEJrLsxR45EX+1
6XSi+g2CxyZclmu6jgkakKJlR9edf4b8o+DG857PLadPO5eS8/RdMExbBr+f
9H1jSA7Fh3C0fnZEVtmjpwVUojvqwVwFRw1XmxRqsT+C+KusWclbov6pKCrn
/IHG6I//5+55gGq4dN/mqmDQhzQRqpLo+3iHkkpIFOaCtQOL1SCcGgE9KFGr
AfmY1egmoPh1pEpo7vttHTsdtY19D9k5+SB7RHDVAvk7oqbgHBrCAKbxof/Y
URR7ZHXa59rIgyObWSvD4Slf+pdhB49QH2VzVowcr1noo+2W5tYbVwQspIQu
1Gz90dM5uRzrMF02SGRpExly0y7PVcI9Ju8rQsCBAwGKLRIqhJIxmaYy4I2x
WLoAEaql/kWg4D/uOWbfM3rz6SYrt9sDywPlimtf4pjRIKaUrZTiXsvM/RVt
/mXsPFIFZBuoQ6ozij8bGj7WuwTmzFcKU5yYlW9ZiOsSCzlACBXNlJvoz0ZG
+Xaabw5PKnfZrMWSX5AJDLpEDjKgjr21Rw4a5Y+tQ8fnISU5JsCKvQIVQHI4
S9CpPurSSyUdcBbcbGnGGYkDuoeuXFWKVnzISIKBiAEndpiRCP94gnG+ZjBl
MSeOJBG+NQRvYhZyJh+HKYe+JmgLKRgcSF3QJrgYuyf5KfMWBbMwkaiopBD6
YfzcBVMwMBYI7CQMqmi0YtilO3fiZjS3CaKsdf66Gx+y0JkStkDSbEx0ZWFy
uhO+jMgzbpP3ul3SLk27ySKRaOJxU1T93g0qZSpmWMGfgVR54QIiZCM8hpNL
2iU07Ml1ebAfHcQcomA3FmD+OKna5Edg8aqwFChf1kWYTZyTpcngB9tm3YL6
w8ixfqp0ChzVQr528jFd2vk3vRZxMTqL0m9UDzqdgWBlEsDWzdTsnBbj3Wq3
UT3Q6p4zi6Xc5Nqb4lL9Us+XohDMOrmhd0DzVHxdTCA3i+6wKOXiPNNgEgul
4jrEq54yLI2I4Zpr084IWcDlHg0QA5esQuN0LpkKIIEFNIAiGO/dEmOX72zq
jhBa9D+IFaFDHT9OuCt6I2KvIXS5bnY+R0PCzgofRo8FOjUdsfuzxDN41vxX
YfmuSsdGXyzz+s9YLxg5E/EJcA8q+ZyavwjgWfnKldajRm9PG/SdPsy2cXIo
FZjLCX9gBDR4zrRVkKZSjc7v9phYDx9EKCs7AGgUxloe6zB4pWYcaaYUMxZh
Sl5KTX1DA1qvzm9zVzDTQ6ffOwt4e5rU4cgnp/qh3iYA2LL6S8B0qdgztg3/
FXoSDSZDqHlrGGsLs4nl7vhCSzzOhrFdEHweKUemqb5VzUbm6DbTRWuxfgQ+
zKQnfJ8c9xrG4Jzh3MscuRGv2/akYPqb/++z2nZFSBgyOEEY1XwXH8F74r+x
3fcNj5UK/Yc7fSszLhPfBwZizPVzXSzjYBVljsufDYkdfzipbKnttDH48yYH
K37PRmzLhEw5F/IHyqADe6p9shU9IR957McccszXUMjnHs5Ra5BmwDG3RghS
+KIv5q6Rxer0B2LkXS45RNHZRlHJcfuddziLLt3ZmGJqXjGwQo4yfVworjBH
2yPUbOVV7d68aEa2NWA8ctpYxUd58z6AxZsSru8BQ5oBp47HUYjWYlqYi1Yp
4bFCXdWqMvO9pQJhCY55Ib2h9sPk6fiLZqmWCeWctvBmS8MiqlzxblUjRZu2
sM2NE6WfGpnFU5yU9DFHcZib3GoKRhXfuHgFK1p9rntd4fVQSgoqJ8RhOMlh
yoM2H5FBlZP+UAJdeDbSAQohL+5am656Hc2B1LNSDh7wreWUEV1auIyqFH0S
W5UoGjkaeynbU2L/8DfxDpjlCj8cxSQSbXY4uAPWun9oDBmGPDFFBMJ441/d
0qMJAha4+plIAgAjhDjym928tHdp7rQu2+HHXee+sZuAI5gXdF71lAjZ+dpU
oqKyfkoEtWtc6siIDZ1GEeMpkGm49XGra4VfL8dwh0yt/SRlEC8IbRq1e3o+
NkOAFmcYknnXM0AvaXZTuZrjkcHoPNPtkhakQPGwdZYpgcr9otBaoWRTSUDb
6BB8ywy8ZnD3cU187mu273CspHflzOpgLNqJ7l7gwXBzWa9szd6RJZLxMQlv
EFXxMiRn0cqFuXiKNkG6UDvWqA2AADj1r/YLAK9MxMhynJ0B9yz8dOPLRAnF
l6cl5/D9OgRGZphfrW5INoWX2fr9Gi1wOlUqoI1fwas8FxUwg69NUQvO+2RW
2ElYkCd4pDqtQfwId6ruwYxYPik1KANt1Tc+yNES3rr+6fhtNpDpTQCLgYmE
K3F0YlHVCyjBlyQpYt6dGTiJtRCNH7YFCmnpcwnGDWFWA35joprDqYKSerDg
QSkA7I1rjdbQDTUUihc3LGu2arW/8js3y+3hkS013K2VcdS5kdMOSCOuw5Ec
kqnTZkhYnA7mPbIptGxqmcBrOAxtLKH4HjwM9PvyvROt4O+3Z4e/Vyf7TLjo
Egk2Jn5AcJLWy8odmFi7fFVmEJbdafrt42bHFBLM/F+cmvy3sLVp09HyfZiP
HTJBdMSo65Pns7KR+jdKs3riQqCwf3nkBxXLzS5abFUEPvVhpjc2jZplDCrU
xtduEb5gIUpuh9IvR260qFZ8g/INhZ0pGaU0vUxVscDkUmUiSg7mNkwNbQyy
owT2HO7MHIrHJ5ItRAixuvPXv9tWlGNpNxw/DJ6vhPu1m0I049q84EwD1lbr
9B1wGIk1GfpRM1Da0lxcz2JxI+0KZrZO4sCi+3MFVgDPGpYaiXjunkMogLkg
fxVL2dYXIMhQ237NVihQMpv6JsGDyuSqqMurPNBIu5ASgtazHegD01Lf7nqb
1yIwvyEBPj65TA4nLOLJTarn4GxbOD6xZc+GTeKej6FL5iJ22l26L980E1p2
qFKsoczDb4gILqDEucOV1ayWUAzyi1UcyXj6Syt62wxwtAPeri75MRcveaOR
TRObaCmQdveVh/kL0uxGCZCCZCWqNiEituBZJ01XWaQqP1h3pgNJaT8GNVF7
0FHgJhtmViQkYkan5luP+9B+8+zFpuzlKD9/0OtI+yD8ze7X+7lNwhCSwSWK
+f2Nky6RhnTporOINdE1ianTya9BdHgtOpFwfwSosD7M5I7Hm0pclxVJD0Ka
pwxEabyNzqrm6ic9D75XLTMAC3D2ihgG5Ef1xpTIQrV1EKEfvQIKDVkIF3lA
8gzZx/tWJdR5Capj+xGnpyeATyYTCp1FaeicqrdQHm1OdJK9zObqNq7araGW
RY5MC/g9BQNvYU6z84nQUIUuN4V551rbMcvKWrui/hPIuslG/YPFbt6lua40
wPDAMGMZXIJ4M4zvMOeYKF9KogBtgLNk4zr/szv8vjN7QGMrAFzMYQJpsbYh
rg7gwT3r0dI8W4cloZTEn1g1k7yylxVZRwx8rmfTIESJbxX0x97JGQxUdFVa
UPG0zQEzxdAa7ggankZ158iY9TnqiT/baIW9q62pN8ndg+b4dWS/LHGhaNu7
KPid3tyGaUjKhPOpkkfCCOnO3+AqsEkMQOqUNTDsDBOgcGjit1DxvpllQOwt
VvTnRU9JfXIYeRGyahwE7UN8z9+EIfMX1esmzZu+suze8KYwYCQG0koZFLUd
Al82g8UGbXFwpdQzv+BwVYzCEU4mYqC76mHfEtv0zD5JRYLqDr1YqOGfORp0
cwKwK+rVmb3EQ63jSeGlg1pY4vmTq6YkWLunIBrp0ZmfT/Ce+1l57o6mBqFG
b1kiZtsUs5TKXRoV2NIKiuTS7qDGktiWqfWixIjRcdW4khpb970GyfOlojbl
LHn9ORs5MUNIlSC1BNHtSI/06I7c57pKVwh3pSuwBgi1acLmaXn2vgSeywiW
56b8nyqTKVu9ipqIeJchiwZBghfjRfHpUvVsqg//HV0i6NAWOtUHWGuPgnNC
5/ux48rXOnKigO17QgojhiUYuj1YIvnapkqJElk8kdOTnF398cAlHxsef4Xj
1iXRSqfWrADuAWvI7bxSAq+fUBJIB5u1OWndVXZRYsgTr5busv7gh6C3b0jo
b9umAERJ3MhfkcfNE2Z9xixyOflZ/KhJibi/Ol+I+JtddDcFYzrfyQaST2F0
bFPZx/JfqSDyyNWbcts25nkMVK78HqJOq44/YiyJyXgyl/vnyj0hqN9NYue6
rZNmJVE3JyEXOKkUy5WPLPCU+EjYuf6ySDrcGUddg02tQci9tOzqtA3P/GEA
KMWmYIe/QaOFEehe/PZiGRPvBGoLcecxcrc1FQ52809+ZAYNk7kcFeDI2XpL
0H1MZ1bfKYRYJ8yguAAAUYPntnrgLKVyo7bKDENDZkHQwLv6k5Q4W50X9GaV
wiuGJ6IPC77YwdMcehHFBxi7Go2gXxVNNoAEZzwHSCISKsu/AXMr2v0wTkzs
pkJ7RBuYO0oIx9BGv0/InScv7t5pvFw2aDAczs94ggR3xSVMFBIbEKqSNuf8
EueszwMFlvoAVonJugu591jRNmdN1GcAA2ykVKzgdMNOBPJyFW7hMeXjazss
WQaoF1bQ+V/NmYiSZM2gEUJSWHI2rc4K6vHdeXvhXpDjLtR1YZ7EP7qh9rW1
e4tBMJjsCLaU79MDsrGnqqrkQnRgWCVNRlCTfdbDhtG8YhEie80bf2ycj3Er
GgM94hatDC7/R8vXGaXmscK1p2W5G+OtWOAcUkdU1pbFTLuB3Y/DQswPrj4w
0gSbMOyfnysGNKFAQBRw4e1RYe5unwGagTM0KLtltJxpYx34rxzE+rC5+qqf
zjjnNFzuKrlnO+0FKmkjZPz4ucPjegvs30moOSzShSQXqRd2F+l/hF//+opi
ELF1rcURCQdyA8I+Vh8mhisiuhIiJccftz5En2PQwWew6KIhjoG8lQdJNP6E
1okalaOt2mXs9KGEYepepxAOTwJHSJ7iymwjQd9UXstoeXQf+yMGbowFJouM
AjKMGaxVVcOkW/igjmreDLbOAot0pivVhSlWCSwmhq67hGkhMxELo3KBiix4
6HFEmG/iFC9stPNR5H5Bc4bEWPUNe6AT8Tl0evM05caMFlkrG+KDQj5BED5x
YITFyC6mGYZecTWCW1r1X9t0xpu2YK3k0mHNdhCf9IPbI1A0xabMU7ynZq3I
a7H+ilxUIh2Ci25DIQ9NesZwtzPb0Oa5LnJ0s3uk25Od7J15Amw2Rxq14ZK0
HE+q/AfSAxoEzGpzcWQVqO54w9ZPDcgo1JmFui9O7BudZqw4YKzFiDobMw1B
lDisqPsau5aD27j3kj/hazDoC2CiP/1NsNq+bT8s1uzSpkVFWEt3Pi33+2b9
tzSyzt6dnxDkDE5MbalyMUXBJI0yhPg6v76JAhJRP+u5eVVOFcMaqkPcNtqI
8iKRIEcN4rcm6ipXw2kxdfiCaVN5ao8bCONFvleVAkQMhku32RVh09JOzMhj
Zi1DMYWp6KVkAHZzoMyb6K4we5rr9HGG0iP09VmLk8mubQnf6ZUFqmgLDDd6
u/Tj5/BnJ70bahDTHu2ScfD8R+HXdUxvhK+zxtWI08ocFAclFDyccACWx4Ec
OmekzqvMoq5ElBeBM08Z7PjP444nF9bXQYRMtHqwOcwMkV2y/AyHJs680yjg
dFKBeDaQqF0mIcZb2lhsOCBJrjdu94CMYTNJLxIGpXrOW2IsFP0EQPPqdeCi
JNCbIc0BRSVBMaPy9jox5A8e/Poqh8FmUF8U0+bMIGGg/OHDdOmHxBJOYfnd
5rgtfkhASiSX0nscWOpiDhirS2Hs/8oLpuJbglN4RfttOj9TXFqy7lZ67vpZ
muHRVjw9G+uCHiGJSRX6AKh8HeKi0kO3FuFKVWlm9pZa6T6buitW0jNJp6M3
F/HRnBDzb+a0L5ZUtcqzI4kloD1PvW1+Pro1Oubi5HGEB90gCqBXtq/RYMgo
+9IvJ0qGPDs90B908Ni+4arFdry/GRqKnjtDOCgLMmEaRW6mQGWGhqk6GlSM
tawG6mmSnxp4sGDe5Qq8tBYIRNB4OjTn7AFDtcPDxADaFHXzlBvsNEPSoJkO
ZBfddbSrdYw3g7mehmmfxi2OWOXdY4thTPWDA4BKqk4DNad5Ab1bL2Nx5W4E
vyC4yBtEpcKDDjEExghx5B3MofKOLcSx2wzJrISKHBWYiFbnKs60vMp1jkVg
MwyT2+j0m4CROAnE5LlSs6uiBhVTISE6ctpzzGIsYsZocl8NJnP2FuzlTe+F
VdkSGtoL6BwrNOGOk2gKs4p1q9CVe1XrEDyTi0O8OqLGCmI4RH9/vEcLzk1F
8W1ca1dMttHyuI5zsmzN4toBuk/tBNeecc5ZJnhcR7VoCGlMVR8/IjYmPYFB
uF5NTyp5K53jzBsNE6a5eN4/EmaaWBsQqFGl8vyy6ZQg3kFIhVVO41Fekpcg
mtC1YN1ya1dgazgDvyzw2zXcrJoVkLMdqhl6G8i5YuHCxvrqZZ2eiNbY09cb
qPgBZ7HGSnwWHv+DxjkzYkjKmzYDVA66hyR89I3C5xXTa0dBKgDf8JRkKKPj
Qko1L4t49turw80fVdHGBAmxU9m6nNO6j9IMuLuBEbzORoQdRmGXdPIEHbKZ
Jv3ZLIHziD/+wYoJ2Af9+rcdTenil9oVqgkMjSNWQAty6XFuJ8jE1wFWjQAh
pst5XmzhkGbAtqy7WzvthKiNrHSvXjnh9GzwGutGVGqj19ORCh88/4jRZx02
SlgHggE1GBLwasch4MSnp19rAPP3yaDNREVC0ZSzptLRgbcJEP4rQnHzS3Wa
crxikVyq3Dsxy7/zeZCwAvxclK2UUuDj+6mSg/3rhbm5rMJO71slRaVTLHVg
0kbI3lDkzzDAYEKeCsXIDLcd5hHuGz3bXHHY9LlWg/mhOArKexTkCy1u85kt
iodfMexFF2tek2FfDGZERnRr/qZlexEY/eFlV+BU3gUruFe3BWCxNVNha3Kb
GPtXQB3EDjjpleNlNbV+r+PNXtXwAH5D0JPibsAF7uFRMJnY9gxzQUFT32L8
QQOvOk0+apfyfF/lo7M9Z+PFx94ZuDztsWPAe/MwE4KEb9ZI7PszeeqduEkL
qzO3dn7FbWJzGduCnpAGikKklEaV0EE5qjbsHSjwZS6xM51YnJ9nIsSA3I2b
nseMcPt+U64XUnhw/YsJWCG/LRGcJEVUdWHxEwUStlqI2aPyuefjR/3kOD2f
4OnmW1x5rS206/NYZIdj9+WAo8HLW1k3SLmKCx36a7Ob7G1cJERoXda3nK4+
UeQYtnqIm5PmgWgSZN4J8PM7hetyIKBSt6UvZ6T0qN3lmxZY1vyqo/Nw0p7l
8uqM7QZKbOk3HOSL6YQMlHKUYPu2VG3l6UaRkGGbtUQh+WCI9RSdPY4AfCti
WS6moS/b0LdHaZUwfUQU9PU0qE+Te+HOrqrZm+h+fe7pJ3p69cZuOlqjxTcX
m8zQEsyoTmB0dkXX3bnMPkffgdEis7fO5wMCOCl5Zq4VgxGbiUr6l+gJlVY+
YFFSmHMkzwO5Vfre7rLw/3iajEtkE5wNr3isn/fhxAt8GKhEToDkbCOi5HCh
32ZTOoGWqTK3vcZ9cueyZFmcy/cB23RT8g5LphZ9OojelSsmP/pzt4ec67gs
bIBnw9BAVEbfUu1WHUXPpWQSh3SoK2cDTcIDuDRm0zOcXBa3TUGXEBIfXkMx
yvg+Se2Vycv6lUgR1x2Akmak+05f5DgqvORCbMMRzMR4BNgteNqeGAd+P+l0
s2AIE8L4eAmBlWDY6aG1Y+41k2RWmGJOuAYa49L8F/5iQGjgv3bXdpEvQGDp
ScknN58lUZfgQ/w2BooCrDk1WlCss4GGTgcBh5UYpK78xPpsoJ8CM/olDxTs
QmsSsuQnPFZExkyXAYTRMA7zF8IsgHT9uOYZDSRc/ZiLajYnMkdA1OuDSvBc
wPSSUf1hXVbhlhHtZ52qSqnJ6wbw+Mo4l1qFJgFOPF0n4Plt8ntlXL6PhmLg
mX9E6DDmrJiK9w+Jh7qhYRjYIFpLpKhcIJoVwX2/YPsqLPOYjrZsC9Od3c9I
SVuytrqKnzT3AGP7/s+MqW6xqylUk55tAjaXMb+40NrO8xatFeKph0V4YFDa
8A9HpKscZM1R0C71L3TLedOi9Jd0rMI1srMH9a5q/e0O0JVpFs9sMgfg8lIc
dcCroo3OVYsRDI3srWUyjYsVJl1QyHgL/z8CG8UFAZbHmiy2eEA9EELQHiqq
9+AOsqD23xG413/aQGAfeMZzszOosPj2+xAQz5sPs9V5nWeEmY7mwNTbe1KC
tr271I1egasEdrYMFGbWhdYqlyCP3YTIla3vao1WI7lAGzRb9P11LFNBADxU
aQ5kVUEdRRXpySrtN1cq0VAomLK8QKWuDXA7z+xyvU1Xkz9/8owh3pFsCRTY
IZUezjoH64lmlhthjJsdFH5huthYl8HU4CJxcVIVfoQfWmNmhNOP78zcNrem
5wLR3rCGyxSWLfm4WgnHYiTsgYTovEQFO3YGqQEyswcRzCTtqAotvnx9Etwq
SXyXbvPNKzqVl2Oh5CBjbJcErpQsIPrAxdBJ3ei2xNSW7TBRv50IK4d2QIOa
EVmiqs2LQkhs3dDGGJ4L0xNkgk7W57xDeTZMJxd8eUSxqsGO/7ZMvnu5T0p5
dk5TkX9me7jVc0GTOg9yTLQ7gtoLCkbyOVQs9UW2/5ZB1qtMK99E3cwhKSEU
xt1zYNvA4VpWTfbhE4JksHn0ZXnl3ZWVziXO1blmaVEbX2eS+rY5Y/JqVT7Q
RTsbQvn+moBGMliyFOlT89ipPWo6/HVRlI3axMcjqKEV7nSLTnVLP3K2lx6L
7U8Epws15Te3YwR+viSTE8z7Z9Yer43pFQCO6/EzJHAzDEdI9v87XDh9L4Bg
22gghmdBP9neAHXPGh4qHAbbC7D34mpe9Lgfxb+0yWU2UgIRR4h6phF6ET2W
ziWS0Z/6dQGtAwLPAa5yThycvF92lfU5/aD8zOoY+Rp+lgjFNJ6DMQlfLXzC
yJ4dGErWSvwI1V2tXIAXF9sh/JrZfEB/dT2GyXDDSK2gHe3tk9TIZtjX7sVp
ZVlZD9hjKYZEvvHSzrC+8WcFdnMUh5Up+PbNHJuVLicrbSGuyNk/y2XHqte2
jSBJeDTYi2qOh4IV6algTlfWzKjnGB9VUyySlA2Jgw7avyNld2FCYTQcxaNi
ewatd1XfYIBG+evcmftfBHJdJ/aDcPBggaugO6Gf2qMatRMw+U3+qX04rIjM
PijBnSuvZhvaxSZeHS5e0EKLmYghSZvk678OEuDvxW3eeCfn/FUzDKuYoqbL
zl/X3iFviiR+jMiiXyF8kScZdB2r9VkzUqzUzGZoUESonUSJ5+dw3jEQMPE3
rtOld0elgVYHaLY2FgLv2cuppkYEALkimubp0GRZHwUcqeuXzdyTg7dFMhwA
mzbKMo4a571LRl6/wN+/QiL1s5Z5cO5khVMtkgYzBD8HtQPjBS0IEemvWiL3
8YPMrNI83zphI9nK7lHvrCOxkqTdeJ7Ez2TbS9fjG5JgnuE2Svc9gIASiQtQ
cdabbJa1xIsrCBYg2tQcGvRNv6rgp0NMVyMj1FTy+fix9tNKwoYa/E0aGv+Z
01Hl8uSULRR056r21eOJ1h983HiBjnxRCjFCV3oWU9hVB27KzcMYOq0ZAvwf
uRucCsG+ZAq3gGjWsLSfRHeOZTsd8/gwpDeTvxyi4WgjcQaKimRX6DxhuYB1
WuW3YBQDfLECCna86BC4MUMQm5PrMR8NNn9UQ7gtChbNd8Tc9H09Wpw95LUY
BQm5lEMZC61FOHxEnLIxXY0fdEDzK7byPjWCFYc111O/+PHDorwVOOsCpig1
gRgQYe/lKaYnGTeNXhXt3didz9n11FsUxToUsBInJbRuQJzx+MG1QvwRaUIh
xh8LL6HozI17e6663zd52Ag0FBZNk96BLBtvYlV55LklCz0Vob4v3BmHcedH
l35Pb9WyQRWAI2Ky9ZwVO7HpPxZoMMTF+o5Gc4JdyyKBsFe3McS6NiaSts81
o9DPlbVMkYDdYeKl/ezCyxYp3QVLd4BGJmq579ElzR0Tob+chJRrv977YSyL
6f6rB1CbYfgbaHrTL9wCHY9sHwY1eR5Hn7YNVYbEAxS+wjisKTYEbAuQglq1
GZiwkhbNjOSj+wpwaeJ/S0aHiUuDMB1A2uXXnjSR+Wa+26PnC9r9/AIZS3NN
vhkm0G7sthr8EXUn0EN42nKb0KFpVuIvjGHBSEItcMwzh7uahYuWMQfttJgm
+wLA7fLGe47355KgWKmLlqFawxgJ6LwvAYYy4khvihlTm1pD5jBTRr/BUv93
R3dDkxbb1MVEmmBuBbUZzsIq2GaQF2vYcHG0zYhSuTE7yCfwjfiURpYFyTWR
+laneX/kh98TCUz4XiDhi4h+WuzxdB1YPPa2GPkyrnGKLw4b5PF8UVTHoD33
lbSwPbKCKj1TYNr++wFGmbASmSJSsFuHAEC40lFUUB4LlAb/UO8jJYn3T88Q
R4Luph8yIKAe36T+B3KAoqGJkkVmdBc3XjKwDuIi3OcPUC0fyWTdtkID6L+7
ObkOCydbUS8nbbqP87YMbxkY4FJlMzbCPoPQRhkxif1O5czho4MgV98TTnXU
nZCVtXWjsMX2h4JZ6JDaf/nfUCrKwAXOnYED6epBA1yW+DekOtG0QRyrjVpx
m0gaaEZ9pYoFG7RX6dHAGIhwihd8GPww0e1kOTysDyLliCHCUTdnPYPdr8Bm
TL4XgEZWcmKAa+HtwVi0pQI240gP86aGGYcF+tO/XIlScbi4wd7U8SNvsnMs
nUpogPe6CXkgYne68nc9IM9NDKGsp4c+XyO3j3c2Vv2xeCws1dVHDVJFtz9p
UxrOcTBEOn9Ig01ZT5zok7evXMKqICU/vSRze6+PhUATSqvxWHCMDZ+d29/c
M/XvtC9iy1jDcEMSJfLQOQ6/lmV0X/NHJnz+KDF/NwKoUulxQvGWnmF4f7Li
InkNXP/y0thKzL7YYW3gowaWFA1up2oBiJUxFFFWi4nahrgf4qD+HT8mZGoc
latoHvE1xBcqH6N+jJU6EHM05xs6Lr9ZgNzlw0adH+YO54O27Fz32S92KXFj
O+lvwhsI5mFV1/l6XVUg9Nj8akeRPoPIid/nhjg2NbXzKmVqrkVWaglNnJc6
rYg+4nI1D50VWW4DVuc4qB3hJ6f3QP6sLbJpjVWiyj8+fyH7heXrUQDEu5dx
EuEXOMkJzceknkrmOsB/k9u8YNLWxOKhXb0i9rbZ9i5mFSzYOif0jul+nWb/
C665w+AopTtN0shb6khKwXxK/h32cP+N4FkPcm8EnPXDw9Y3EBcPD4lAD7VH
T1g6iE7OHeFZLUTDmAdgAfCOwaG8R2xzHMPdu4g0bPTboyDnhDEKKoZpfDMi
AFMdV9oZe0xnJMnmtFqDzfFjyTYtN4DOWc9gC6Hz4IB0DWmtLS2FbsQDpk1m
i74t7009awi1chrtQ+HEV/8VW333Rz7tPzToxdIHCbaRJXsvFjkh54Q9b6hV
egtjd1G1sGCiMQW/7k6C9aPwcm0vj6KXzX55FBL67epaiGroshafXH9voE8T
s9JJ6oApfibNXnhFTtc40gUG1L3eSpSPEbCy5IbWiXAWphNvrQVUzMYXMDh1
tTAxlUSNevJcjHtiV/cDMCgJjd/IpeMC8hsBj0/gebblSsKdyc3O7iF3Wbk/
iHrsCgjD+w7N4n+dXbJ+KO8qWIH1ah1mrKZ4i6z0pLUv7b1es/RHridJyN5z
dmKRRSsxaYnj9FsHsmJSS1zrZDZWZOKj9JYMj+xIv48YWzUAOxm2SLNAfF5V
oqe0m5ila+qYzzLedp0yoNdlH261uTMuf6nOc92fawqRYK9u/YTb1L+AKxxQ
umCuLq01KWqQojhMHEqPOtsxVBTkWIlAbxCS4MetHNlxa/YuTh4Z3H9231qm
+/OZhda+c+mdqgupVfZ+c1Q53cgFvkRtRuyQDcuDZHsYO2XoQuuRPDkKgral
iwoXMm6qgUjJCeQgj8P9oBnFV+K7Id+1cc47s9ZkAMJLSggOFDSm+LnSOlev
nZa6tXSh1Yq6YDxfBOMdRWQUotTVq/KO0GCyOUzS1R0xELmDN1grcbzn3v97
mSWqRlFfzRIsAyp2Ba9yOmYM1tiemstsiUVlqZhVQ6jlzxfLQRb1U3WmDsa4
ksGkn201be7Qe48rZFomDBE+uB7bMN9mmag8HhRnZvCa89cfEBJHjvyphryK
JVhKbsfYn6H/EvMbgqaIuS5EFOiVD7Ty7DfabGqCO29FpxBqzAQOxQbfE85V
ldr7PhpBiik0AxGesYc34E/BXXaVKr+cSNWpYqj96ruk/NIDBPSn3VpTtHcu
ZhM1SveYiMneL7uLe22j259PycOtla/fE/dr/5gRczaIzAj5WzkZl0Oy96Xu
wRBwcLKSJ7IXZd7X8Tjj7dTQMYobpJemNGSz5bMErQZxVTKUjAnq1mhJ+rnz
5El5CkcP7zaHYoZpyr835fl6Q9mMQCxwN/UVmQgIuSxi/HJczdPH0/lzOnjb
9V0kcyYvsKt0m/otibL38CBEFoEUOeMHF1S5r4FxM2D7vloWmw1+j/8BYLZ2
6d8RX1aK7DtMfuZIMHIcrHZh8CnBzVSKPWdXLEobG0tOHoDj7QYZeUmZYwsx
oq2jcOP4IKyrtA9N11Ud/deNhhGIilSyWPbaQIdVOa6tqxmqZaRopMrK9X98
A1NFbj+/ulTBFwcWyPLfL1qVY0J0sIYbziMIL7Aj1Rq5jYk7sUoqa3Lq62wV
bkL6lV+DKt5eLVMsYIfBr5oTzeZVgrXBjtFeFqmT0F6AX+xGwTl4YUngSrgR
YtL43eveZFprTdNXNcC2xJDmbosFoNaYD+PXDdJYCO+HgkfcMmu0Kxn1xl5e
hEP1glzXyCeIxeF3OpQokquoGCY/nGzkj13uM65F8g44C9L5DQOPqAwe8o4U
ez/9Mw6uycf//m8Oj08b1veAaRRPBCsAxnvxAzrUF+p02xu//Dcel3B2HBzF
ZX57un9sRqMFpkE0xL89n3Y0nvYwzgyeTLFCMfm3NbwoFb5MfQF0VV48s4P9
i93OXmXd6og2AcNWNVHuyEBu7hcd3g93Pnlc0+8vVS1nEV64BNQ4UR2N3lwd
lU0Ms5ioAklN6ZuLpXiVwgdKfDaLr019WDImYkJITukkMZPV9cZl+JGmteRL
xYJa1apAjQ3pV+P5y9Jn2ncigqub4pgfXiEZ0WLTiA/b6tCF1AXDZWtFDs4q
+rfZRo+ZG0ut/WDCGpNowely6SAjOK6fGg5nWbi8ZPHRNJ3L7NdZuKMTUX04
QQcyywR9tmxSVIBz3VGJiji1fYMiSNaPOK4fUUomkbkkKBG0rW0iBq8IuUy0
uGnR1r9tu3b8yCjUuvU2/R1VdtAhw9MbuCcRFafL/LKdbfXeN2l8rijO4BtS
DgC0vlcdk49Dfxe1o/gr7DqMMBQQyFcA+XniJL2IVHWwtIzeSxu60yC72klp
uhv69sghLu1Xus8vxrcby8dek2ygSX0W1PPYd618kB/mL4IVuD8+9dwkL4gj
ho8YZk5K+uvh9J9Yl97rB1lkYGTZRRE9Fb89Vuol9QdzDT+xt6kreAox/sDL
bQxS9JKTKHMmjI8/hh0mRazbl3NgXzitF2rYSabwv/Vx8fPTb5lvK+5t9KLY
7hR4JAbkUJS5bCCIznxwXKbGWhgT0PZgIDbkUdZjvLP8IRfmQu3K3ljy9yC8
770oPu9rV2IYkNOi21DLNEFfNRognohB8UZfwsU4JHg8U/ZOJMv8o3W0rd1h
GTEqxjxs9zGucUEgKDhtHpfYackO2jTGBWEmHBaNLSqG9B6OUWKTf+gCIWMv
hxpHIlDF90OuwD6Dq5uhdKFEV1A7ZbtClxKOBCGP9IraY70aA0EPw2TubKXr
wqiE8oo1m8HMqZUwIakhjHNeMbPKIdZghmNujOpZzi8BCTVDVUrc8SKcN8J8
n2RehCSsJnJKpwdJWM1t7Z+rF1MpLAifkEf0Wb/y8zbYDiddRhek5wH/hSZZ
OFuHYuqi+MzRv71R7cgKSnPpNFjjEUCwWCw2g1dWVqm1HLK0VEf8qHLamqqq
c4Zgdnaw5syfkPDAD/cejAP3+TYwNcVXy7mq3jKdKE+MM3t2wzHqxerRRyFD
UyNGRrXgLOI5GSu6I7i7eY20je8hJgxRxNSUqjYK9pfzIL4kr9GQBZWQW/Ak
+7Ic6HuRT7JGE9MRs9HdmPtDWDcX3K2sboBA7d6uyCWEsYZsDcnvDBApmWQw
7wqAXYYERtuKqdL7GSYVD01jpVnKz5b26bfNt0Z47iiuQfr/DvicUmtN+otk
XUg9IMxv04cDZAE3UTgeTAB9xVx4IyS9/YWXstaUawFaVmzkW9OplJ4WeUAa
/lWSQqKkugvY+tJ2/GqtbjiL0S129Pz6uBKzrLxsgYxM7r/AoS1+GdsYliNY
Nx7EL3IYqNl+x9SRSu32tA8wR0Ji0y382TYoQ9CwV2m4sc/6Xx1WUGQ438Fg
IVWkUUXJ1uW3DTtO1U9IOgrGKGBfToYGbrEbGpmYxbjNIGjxefb8ggwjqEcG
uBrMhIpBzI2G3nZfP16E831Fr0Z4TaX/dF8Psnx4WQF4jt8nIbAY6WzmAD/F
TNO2FMj4yx6QJWfv9hX8sgrMreCEWN90m0V97yih/OA1CukeP26EicM6nJYe
AevCIpqANkOcjQEWCz5o6YVJgQcVFNzmt1kyF0A4LT1OfBncdW03VlzAFJuI
CNdvcAsMc523jZpOvHnpyvCGxBU+saGQyQspIgM0htjUHvcPlCvq/2YwB6TO
+dtBsnEwZh4mulDNmFaT8gE3qMwJrs/EtKtNx8uJ5TABCW4Rnha1daBYzswE
w3pHZ5Y4QWYapV3w2wXeoJ3iRerkr7Y6oBg9NHMAuNBLNt74sN7YY4VdqvpC
PYo68kNVuU1vpMnHm2WsR9W4p3jjzbTv7d5bCnTgMRm53tR7+Te9kGrByxWF
f6dQKQyxFRxq5HgI+8m5LRjZzu8Di7z4iGrHlTbDd06mAaWNGUhhrUm+LCHb
PTEkzDM+Kq1lJ/Gq2wW5c+5KvFp9A9SZA/e1lcqM3dAfkSEl5a58iS6xnn/J
cUXnVWyfr+TU9HqGjNUTcnhdcXCV4p/ybqT+j9c+aNE6OYgu1GfyDMIaFO8D
sT3P2aH7LiGn79qRL3xEKtnKqAjgx2GFv8m94u8zBDJBl3yQonXtypeejAy+
86eS7tHDANW4y+a3bwe6ai95WZnCxX9HhGQmYCLrTJLl09EuTknezZv2UOIX
rdgGVXhWNVW6GotUklzH4FnDz6+JNogzEtMJgDSDJE3pxEeiLmoiwGKOkNg0
pAQg0JQJrPJvcc8UeLNBc6a8gZiwnd7qj5ygyQLzX0hib2vVHK01U5xwJOZX
G+To1adqtwgW1OEO5asmwWFnQJXTECIxVAxmHWCgTb7sqZY7FyeI7L/25NOg
onpqhyv9p1ALBUfCi0667QDvs/v+HrcGtAUUzMbBiVmnR7kiW+4IdXlqrg6W
/nR7SiAEW1dPrg6kvYA1QHc4D7UyjyLSbUat+NkoCPQiKLUg9CxCjrqA7xQ4
5sT46gghfnG9DQdm+yfbJySCLGzetE8oCM+XdQApE5a6wKjdAQHZBaIbHWb3
vslaPZJoURFUK8R4lrlt8HO2MIwTGfcNRHGNRMma9bH0ajgQiL3HTBqjD9sI
YF2MbQsp/UwaBcGhEYpo69qL23FBy9V4q4lYbJ3we2fxz+ub4nuFjw83pVIF
aYdD9RsbwYKa5+/SEVyimAlOieIphqzRL2gMmPztHxHt8JnNJtlLFBJjLJ3t
Tbu3Q0t9ozJhuq+OCXEDYF2hEUdkDcY6+cJKR7R/3HQxKpfYauNnPfNLKXs8
Vii2Y1P+tu2Kt5yuj+C01CeqrmHMiOUZkoNgngGbyKX4oVQ2FCqyvaW3LKE6
qPYXlzdePDqt/ySfxBtIWW0KbCYl9m2oIeFINzQGBO3TWCpvaN5U+WfkPgBD
ZMgJuFqZ4h8NHyHhcN7BppYs2k0ZU5+aw26bTYHwDQ6JQ9VTirQgdjo56Q+x
dMipKRfT2HhDgdmjRozoK1mYPOz1vWlNi2F5ED+arZbgYpFgCm8dmfcDGocm
vZKldXyVYXRlLlnqEAM578QIIE8GIB7IrLm6qK6cIVgV+NmSSndhWzp0GOHS
aj7eXCcvEHhCB7dN+oShNt9Zu6mRk+2BBYh4Es9jkxZRH+NHn61/CmwqvaJq
RUVs6s4BMmC9HFOoM2qhBHBWp/caBIwqSaabvUhUgYYVMjQc1b+RLkKC0Gc/
tDH8PQG78b4frLJ6gMa7cHuqELhFRmz/wL7ag8KC1l19u55hDV9nAiKD5PI/
ual8pGc86UsrIop4cSInGwRNdBvTwJKyj8+mfzPg8FNZbXoK4lrZJORipG2V
VO6pyHtsHliwmcKK31qBdH1eXslHCZkNzsGhizR7q3ZM9zvK298/Sg2U5QkI
sgzLAUtDeJaSwPTEupBCIw8cB3/tU4cc5mtEpMcMXU9/+l/TQQvq5R7fFXZX
Jz4n7Oq2hlGoRmGkJYNe4Ey3lPjW6sVe1dVhqMksqn07xDBoubcZVTXSIRw7
7iVB+ge9nUwNSLX7FkAS7pJqrHQDlT2g01kL8cYQQFodOadrHaFSL9/509wJ
+LOGh1vC4sBbzsBCQO5o2HhABPNmRRulkBdM9EfN2E7cW1r2ojOJz8pPYDXb
y5smdYR7fgzp9CLYxrF0Dp+2TAjn1EUvCqJQvLpQExMTJlhCvvpGFUbxhBCN
gR63uBG40+z232XAfNWPMkLCgJ5q3L8k2OdtIi6+Km1sn6hiSA9s9LJRo9nu
H3rMbyUDQ02yglzy3IodtTUpZDBLe7ZIdbNja58jma+oz9KrjqEB0MzeQE9D
J63lDoxSeYikOOUGw5/zRQkYt9mxpY1ClOzcyFMPD0fb1KRrYu2cEIsMgqY8
bwomKK8m6Wv5cANqKEi2ZtgbKFl5rRXjst+sIDSQNM6pZSeOb6bb8NhRokUr
62p0MzGyhK9sA6uoywARx/qXeMQFF3wH6P7G2zzfryZmZuWl1Z2j25dR8ALL
n8G1h62luD7mEL55OF4K2/iW6WYCCL9xFBKEItw7JnB8oHiOt87YIf00TWwr
nWHKmG+YfMkLsa7TapWPTEmnyV9fqE9w6lijOgm2YZSWC/ynXBe5B7xi/6YK
Fopy0XKbwO1127vop4kds+Flnfd1DPxKAU+hYXqUFk2nVFdtJe9MpJJDQJ8J
PtLdFZtYS2iocF6h7U0jsKIABJjxBq5PTSa37f8/NGIJcQH9pXQSXiEKwQNG
6pREdN2YEPUd8HCElIe1grlhQsCsos1VUVD6R4tOYKnDYLb/vAvznpgTu/nM
Yv/g9NCoZ1x5D6CRPfdm1lnROGUR2NlXuzv+jrorqU5oE4awobJXG/4nvuh5
U7CQH1X2r/yLTq5jIdsEG5uINztahI22NsjaWg5uqFknxzCLgDEyCBNEc2Id
6Il04+KlV2s4VIcauaDCLtDkeWeH0a3bn+oh8XFU2GymJ7LnMD0yMddiINzN
Zu3z1sY7eOvbjBOB+SbXJyJhRZZH/wgBVkrQOv3WiCW45O5dEQ2r6ckP3mrT
77RObkdopcbvmLLzVm+I+Q48y2l5EgM99dtSIVKZsHBzsnztKLMAMblwz4BJ
LE2/lYhbPcAA6UZsXG+j/7GEo3MaDEv6JiRDfQM5elzTWEaprNNgaPLI7NEl
EXDC1gqMMSitqdl7I0ZJ5QZO6mu8Dczub6d20Tcg59ncUccIR3oyb/INFBbC
LICUb2lO77f+eDaEmpQ49a32Tzju9t2yrfXCcHbgITmq7evopiMlk4l6MHp2
XQZYaAErqGd1Y/kO6jvhLfSD36YBciBwE0I4WJci+JXQJFl9Ilx1PW1LkaZy
vK3aXOFctFrRI3X4+cKYKTPbE8n7ynh8avNmmic6GWgNaFMtXwsAD0HE7eP3
jEldT8htn0dMVADY+a6Fj6vuLVTnW6fWJOWjbgwhB8I9wVi9ZI4HLPrd8rVT
P38UXgNsTTpjIyeHelhd7f5YoEBfifvBbvlYy7PEIXCbdRU8PImQQXP1Wzt9
q8d0w6GXWbB/y9KVBNP1XaI6dQQuhVsoa8TKItHB08BQULRQvcVQEdKlr2bU
c7VMRXCY4bxn7+vYX1Oqq6bHV58C52fLn2ogND/eW/WnellNILVFm36A1cA+
ZlvsMebFFqaX+BseRdSv5TTjWLTAh96hoTblFgvf1+mQBct6dMfwfg0dE390
qGtcugpB3o0jAXxPenCcNfRFhB1I8mChmYVXWy9RvoYig9B3fd0RrGXNkCxx
Ip9uEbq4HPSRcm9diuyYqgsIQRT3RX+eq2d4PurutXMjFUYGkxz5yjajSaMs
zFrFWqMdKnmmVb/WMHRiAsfEtCoHPxgq57qnGNGluk7zgd72YxTHohlF05aU
4PceaBsL1AELT2mR60E0ZIMxvUZCeNPy3Rf/Mg13p0mZBdsgAtaqgwxnFk3D
kR5LZ3qD2uMMm+9I0YkJbAUTT+G2yss2A3U8h31fEcNhRhJ2tySpMD9L4+ho
K1iFFBncmdc4BkBVpeHq2Xm+0YSmCG61M/TkdkFT+rwQrL/KQLLyoLmTBU89
iTekE0QYfOLuhtawHeIj0uqfRfhgUaQ24Ng+6sseGKh4bvurX/uGDbNuSyW2
k5tDs1DsFrMzKrmaFqKII4zEEpoTlLk9BZGTFMVtepCXd0igyAUafEPFWHJ8
24Ymq+vnKndntbPLqUbLqlysOoT+RaC9AkjL7yDLdkRvxBwCoEA9Xqbm9+4D
oESrHLA6CAhJx4/uMR/oKTjizKegthzhpvy6/15pxleTSVzGx6VkKNy6Yrby
j23Cq67LOowqgb1T/Ew+emngWYCTt8FH1mVayaBoHDZUx836yaMhFw/ZO7xc
JuQVoYih1pyv81BruYsL7Sai2IwYqHe0vQv6tP0PPgbN/nhMQFW7BnbEOKN2
K7mAgUYC0wP3+xDOpIUbnM7lo1B16fjDoJvkDoA4+PfCmuynHF10F16OE5b0
pzhtY6StL2TroE5kwct9uKjvDSLnlKAJB7K9BJAK8DSmlexCdYC6iARPB+Qb
G7dMBm8J14aRy539XbQoBB/jS4tuN3NSptm+Vifo0uXUBDpZoB0uYKZBvBiH
w4DgeM+wNjbxBJFylxfCGiMef/+8auvVvxTuaY0nPS0cMLpqwoPdiUCFRL3c
1+C3bK5qXS/Vax3KEIhQP05COioJub8JIFhwYPH1KzFHif5lABgJD2m0nQkg
He9sGreT5A4seDtaAIqvejzU84lUq5dxqciImbluwhUKHC1o71XowE3X6a+E
dUQl0jBivQgVwEu5uG1ze7DyxXA/+dGjFvs5b1FlvPakaRrOlioT+sJyUpbG
G7rAPIbOoiwJAtfgK7L08pPy3Am/iQAuBdwGcwyK9WKC/3XpBZuviPLzIwaV
AAlnSmwHjIJnhMFpot4YluWaHTDON8vnJ24LEL8fYn2CUIxJh98MC1K0inB4
BIwbzaGpvi03lpkImeZBevJ4DUqfNjIoNedVE28w/tUjZc99z16v2bT4if+Z
RubcpHJ3m76DIE1Sxb3K157BNK0BXCoUVPhkFiOOVZnjIvQM2HpcA1ahZ/9k
/qF0BTx3+eWECCWm9RTfzUXNkIxmVWIAZvp5vMGtrrkbCTZuWHLFuhtwyHGP
I+eNA43C5zc6YtTUU7Z6gZ75ZySg5S76zmTwHriQPpVeQ18gTDWLJULPio2e
VYXg+rZQ1WhKMr/N0/ajNW9W49VAjfNBahk/ffmnvFkVLJi3wZDlOSLN063U
2vnZK27j6Pg49Q6KbniCJpjWFBh11MPvM0mxryaFTLutN+wl1J8+SPmKj+nV
HHUdSwSNQhSvZvQToXEmIVD3FaUEm+tK8sdtAlpqvNTVMazq+uzPlk6RiUn7
dX4hbF3W00f4zUN6nwlob9sYcYF3N6n5EU+Asz+3IKzOuAs7YrKA0l8M8ICO
2h7OKC1N35MnallyexUYTzSxOWaa6UxcWfrgazi66PNTr15fiYLDInvi3VAy
1YMg6+DDL3T7AEM+MQ0LzMYOUjlVu+KmHvtqfhesUyHpM7vdDU6h9l0Z0eNJ
lSfO315VW3UJd9bcj987caElz4AwPkyeWmxrySr61ejIdT8gqy1zZdUN4bM9
4pDDpWGmlQ9fDhuNd95O3h8j9cRZyzx27/s6wHQbabdgMnEdW1OneUThaozd
isFJC6kfkpDE2f1aM0dqZMFcBbs74fcRQqqbFAjIok7H6KniZf3mges7nnLa
vEU4ll/6usEOECIugW2Zd1xUBwdfI1Qk5MQI/9LuRdnNMhPdjt2DdRzbYAJO
yccCAdg0NorilO+h9s0+6hrXE1x7Zz+u22Weq+F8iWStdmXsI31NfM3yww11
MrRRlbVDZswBX2rJSyOJbPj8ujBonBtPs20seMiHnujUoAn/Ss3LSpe51DRO
Iaie50F9S5MWHOHqDEkCfmXTmU5m6rY4NJhf9FYKV7v1W/vDTEae8tctQFcc
VMw/o80TkRxQAhOG4Ux7ddfOOwwZuCZtBKe2Ir7GPTVku788MgRXTzuNIm2b
kAlwovNEtWbHx7lq6vzD2yWrmo29U/05EXORJabxOB3G4PFJS6eHB3G+t6mP
h6YLb8wur5iZ/qHTYZNvgPGFI+EWIyC58Rue5CL0qc4XkKonuTKhd4Y5V+0c
6rM/uBEcaSmjG67Hf2S9GhJcWavemGmexrqiNBW2QnSfQzQojhW0nGffxBdy
HN5TB60n+Bcttiq1XJTmMX8LzdO7L2uW3s8WPzYlPsckZe8p/gjTcBzt1His
nq0yLGE+yiseeiqE4KGl97U2SzOhjIkD/YGThSgh6hCoNY6+zXr1FqOQdrtQ
f7vG4PHPQlFdMo/IlnVH+WTy6IbJ3+AiiVZS1EBNenVyXAp9Z9xUSdkP3kQC
e5VmMFZrA/SFivXP4PADns8VrY3nWtwDYou81+F7LJKyjG9fDAjE5L23VKJE
TlyAhywH2sDs6l+JaqkcmU/irs3hb5Ic5s1iEM2D616LZ+xylcHtrb97Y8Em
Hp5l/7WBd2RPVjof0jC7xrmbSs0DIKHehqoe37xt8GFVjRl2yGThwQXwPUna
gWIW6Hw5W6PW9KIc2QugIvrA33inz7gCwzUa4zsaE+2jkMarq/Fdx+1ebcre
lzP6cY0yIqczzvZrN4jRbRt9BtBLaipwym3JRh5uasLJeiVuiW49KChenOYS
mmlVotgUGXDiErJNQrpfgZvBlC5L7Q6a3Y2mn4hTsC/nprOQvqBtQKEaDd4E
q8wqR6WOZS93oH1zws4AM5Cs5KjP18kXu47IX+kHXhaN3MAGLoa+KtM2V2UP
PZp5hlHLqeoxD6SLGROXgsAZPXMiPStCdizIaDCNHSbEaxNUhFIpw0AR1Yd+
5vEb5rfFPeJ7PLVxbFcQjfJ+32ue22QAj6OVxtMTHAfD+D94xAuEmPsvsFx9
s2M3i9stIzZwWUh3ja1ce6pkjlkGOR0Iynqf77TxQ6NF3UG5P9MjaytVXRhV
rZaIsDdDJc4GtQMqLH5rJ7Y9sH7fhu0WlQcBi3z75LgjZiQ7xdjIkTrWJYgF
9ExAr1wU4+4oNb50HC56uED24fHEcYY8n8TyNdXC6UubwBfx5X8lBoF5P19i
FPHM0ADBiQsrNVU3DXWPBnBBAH7opkuZqIlBOOsmZn+knMmdFjF3qvLBXgn9
elT7eJsV9ZLynH18Wto1lumzqe2bgIHqU1pjxbRUMp+Y0gK8WjIST5jLAkzL
44lVmmt9SUamrUn+HVun4dI1hu3HRjg2KDj+sHKbcyG0Z8mon8UBpAp2WaWQ
ytLxiyHafW1il/yT/a01Em6UIwymR2gpY+I44q2A+5cye/UlqTOqgiClFrSF
WNbSQx7huSzP+uMhGZ6I9dwbDtAWLO5vMGLVuOQ52BPe3AmJwUiwzZmQyloo
NgEIbfYr+ZNG+ARgYigql7NnDlgLynLkQF/93gj/FryWGJOCbVnRfK2es4ID
umbwDaxMVkpDKSdGlrcT3QBVurR751uLsKnvsNf3hwKP+WaJnqsp3SM16Gz9
fO4Y19VzxlMoNCg03DG1Sd3nYVCN6Oia99S/IvlwR3rZyMjI5jCj4RsuQ/uL
JmFPn1WiU5zzUoM4l9Qnxv8H4vTmL69eZSFWxvc7ku5rJEeBuaAti+6+sH9t
XDwzkG6GM636/Afd4Wg3xmtV5/z/Wslbtpk+DyQBBkSCZDa/i5svtGkMZLX7
S7crdnXBNohIRuA3DLFdZTyOUa2ZinjAdOzMXSRQvHSIjVxG+VdzgJq8y6X3
3FabSul89myvjdMgz2Gd9TGwycPdvX7GBxptCv77/3u7QixPldtA3hkeyuEp
/Ue/IfI2lXZM7vCdRtWAULgwFfYTMYXn+ReV9UmibO7B3P+TAvtJkcpz3sJV
GU0f6aCOVtQYrZQULDEAL6omm81XXl7Xn9MCxTQ9Cv+75qR9CjpwksdZE5yA
pzyiaO3QzOY6F74FlNAAhosuC9JFK+GdU3eJrFDrtvz0T4/7CpJx18P91NGZ
FZxUYO0AFybQVbjpLk015lzOvcLZciSNwr9IXGoUg6HqbqzF15m3PKc9BoqH
EBLacCfQOffZ27fqm2q5QfJKOoX7meaqr0j374ZeEXQLHmXrvy8pgyrCaX/8
n1DgltmBm+FUIWpJ2/XjMyps8ID1x6cOChxcc9MqiDOW4RzPMJzF0LFCSf0E
hG88GFLJ6mSBbYOX28I4ihM61MPz2fY+5V9w52xlTv7q3HR/q3zWKvDy0cs0
tPrQwH7e6i4U7cDFE0vlPi0mVGcpzTscR9/xn+Gqq51HDbC1UQNt+BbbM8Eg
pVldRnwEp6cX+5D6LjARO/SxAkcca2Xy+iyQ1TKeqqYb7wJEpmUMtmJbJvee
calC7zQvO2jv1IW4f/lgrMvcJZ6m/DkaA4U0kpw0X2MzhuKnBCSDEhmv/6/R
WwpiR84L4ZfyFvSkA08odx0zUiEk9DMmAJJ1zSeHk7gqAQeYulIZmsMfBSiY
cEzQDYsnMW+/s6Jq4oqalVY8vyMIyEnDTNNYPPeV2xBwVvACTQ4T57jA9bL7
T6DG1VpvAiSDTV4wOEVkpqFtcgCAJA5530gMHI2PVjERw1lNp+Oh0BNQFPQF
uklReE3Z15ULhd49Ywuqur/iOQDTVVhsRbuc7WgoT/nHy/EJnqMNvUuyTXUq
suaajQqvQDWo97OolSR2uModDR5BTFGd/vuyEHACu5fNDUnmqSHCYk4rjUWX
yMHs2Gl/WkUNkRXuvZtfOOIOhC0b7Jl6oRAxUnDPOQOe0wlJ1Vm8Z/8+cBFU
BjR8gHcZYdcETLjU6kt3C5K8YXwmYaFfRV1OShPPlbAEYN58L2o4fRzjDP8o
9TZX9v2bjnWranUV/D0VyfjaI4nr4jZnoMhMj3QRFilDpzkNNeVx8f6FEQL6
XmCMcjNaYXnb22JHcsOww8HwBvQPfmIXMxPWHh5FFBlQsEMh6eaye2lQhO9B
Qu4RQgg5MkSgsMIxyPGQTesVKlZ4YGVH1HBQ5tc3+DrDssXaEOKPFkYUGGnu
ggu9JbK7l27Ho+9L6gPo+eIFnuzFbHeA8X1ZARH7k+7jct9qb9ya0xPHH1RV
U1jwAcEhs+q3Y/IoA6CXuKz1PG2e5BDNXbk9tJEpKQWtjvYY+fW5xm97HcgG
4eF4o3BrROcf/vf5GuivFGaNl95AQvSJBUSKyhtGK6uBe0/wV1HHgX07+pcS
psVOIXs7eAsRRBaH8/o6B8I+ujnSIpNsD9NtR3NAPJ6qoPCoACi7lZPg1XhR
pdMx6T8y1LbNZ2iYn17UuyPv85TvEYNeTtb52LbFneSD02/C7v3SluKRJeEl
mG7nhuUQEg0enA9M1080Mxa43qsliN/XdbScEk5J1vj8oeUNw/B9pmJOGV2Y
YtkdoFWZqTtSNd3AbvwCbBpuTXfKfM4Gm5KQvZxGaEzDGsHHlHO7525rwGCd
Et7DDbKUCTwmqOu/LZZpBnRwtNApzceKf+rBhGTy/gW2RWA2igpSfqay4TrH
fBgLenXAce9sp8sJzFvp3QZGp8ofIyw4Edf5Bfv6vRV8r1gzWD/xZfrQcpVH
OFZWs5vkQs7lHZ1FN7U9kK41JSdkzLDD/j7C+eFE9Z55mn8XlxiJtjiSZH62
JBh39+H/Q+ELAZ1DuejeCCFQuBYhlow8d2MFaB6DfcH09WjOaRuVNr/qBLVP
NpdNHYq5bU6f0vG8RxNR/acgT69MoR13DategNB8MJEe4BKRMwAHAm5WFfe+
4UXrpflzwHRaPZ2afVeJFBjXRisA0kCkvKHiovRMC7nNOD0gaGfQTdj9W+gC
NcbSkgbAL1ewW1hvzETsMOri56FiMWguPEqpYVcoo+MK8Z21DEq3dsprA0Q7
tcUcBK9WXPUzgjZbCKgSKzN8CKhLF9wjNTZifyZ3BR6MoMMAiPnZD1dlBghm
qUeI9m162drsj6IwP9h8B8m46PD02S0e5+ZbcbO0OFlRoyVzD1u/FU8f9ZJD
dge82OCc+p/k6+mLxEyHaPDwPBX5dSYDQk8hXKFYv8Ba0fOj99hdU7CPGNfo
VmPlNH9l60IHzMS9mQJOdyPKQJoR9RS7RebafsJJ9zzRN4uZNypxUJI4a/9i
1Qxa8ekoUe24xSYtAKPHmRxITzCidOgKzLbthK95nA4c1Zfyb8K+NkinI90F
hm+cgR8myDAYjJCGdcXD12uqaA/YjiVRQWdLxPfjqhsOfQtmB3xKzdnU+x1I
u6yf+GoE+8GWARwa87IIc6BIULCPzR13rl3EwH07xs1mjD5UxujjjCbvmxtK
seUU++N8PTvejoBlVpl9ORSP1jWxyjlVmycVWm5h9HquqSqCwycxUOIsH93z
wk6kYrp0GJCkLQzXrEOo9l77/MOKjaMbtcZrzCvVTXbWqhvZ2C+gfs4GMg3O
5gdLWvfDTN/iQrYSwL9gQP4lQ64tobriNIIPU7OMsWGZAHf8F1T3+L/9iGeF
f4CyXdLpawgZlDSklrs+FaM8I26V7qpZIZX9XGFXN5U66mPTMYmTZWjNt12A
LUjKsyc51XLCNJptlKVeXie63GDd8ES+ynSMFrLMOFzfyCyLZg7m1la0c9ga
4NwO6yQfrlYWMjqu+UKvKFLoukuCtCaVI1qIr9/VqOQv12X1iACkB6UoI9X6
LGuWYt9MywGVN5i0Th8xGoSxJMbOYXAFMpsj+YoRHwMMLeJnQofTjy6pwtJh
Qwo83CLxmTuM3Y3Ya0KrUbiPOXg1/DQNnil5KFcyq2TrMjLriu8j8ElB1hYW
xUylUsQiLaJJmVf5uam8SbFefzFNP4J+j/BCagOTWDmbjYqw1v5+rUuQmvyM
mxyFH6cdCvZLew/ANUdbmSXJvcPlya9pMFgMgybwxTFfVBkaSQ7Na2p7Zz8q
OZqGnFSOwhfDM48RJY0TUgxEVmSp4dOQVTKsPkrAkC3+aPP5GOJovh9Vph5Y
w/pT99yEVIWgWuUAoMI3hnjRz+Kn+nWwRb/7Qkw3HXbHusr3Gf/ixGTavA4O
Ta4eyJrT7u+EK+jQUGctdkyfjmAYrEjPvX7xyh36cA9DbdoYoie0codLiB+A
2fEbSZeAfrJfjmt+yHGH38Q4xpPWXtwrBYHos1468Gq5wYuaWchy2K5ojOvd
LWFf72bO91UTUBeyqNfyJXlA/r33UdAzhbYawdpidJOo7GQFPNL1/TtMC1N3
il/lVv+kwGBEjEY4c61OKvV7vPNRVFSMqJr0U6T3ZaHjrfwHKXmcCe7kj7WP
TBaD7Kf1PvnWrZMBZHjoC2F0vzHIj9gL9Bd9y70bZm6/Wsk+qIV3tQg2gBoF
S1DOydzCq3b5trEFtWgPpT8co+WXHdSgvxYXzA2jLrzciMqQGSXqTP9sM0US
wQ2IMnmROJNcayoZTYCtm+oBoV0dMIJmGMz6Eum10dYvVM/m13LudEKpIi20
Fjyv52g9KqW0mKR0zvegwf9Wb/ELiriEeRagHPG6R/grluc35JKeA1x2Dmpk
ZNFDcU6dMuKdYltmoCHfwIiIGMI/bmBBfK3mPd2zHFb3I2rzYfkEZ9x+JyXj
+2CjLYP/8nvIBrSgsbo9R8I4CUckdWDUt0HZnQqwNZj3385wmb1i7xcYmz7J
ub9FJ7GVc6OUGOmXimGa7jj4z0V4FSh4TgnsX6xv7b0mKO80VFA3rlofoQE8
xa1VBp5VLseKO7VmndxldJ2b6mgyIST7zGyl70wEgYyd4xGi+2xpFblOaaHU
7yw6m8CyWHrqZGPjhL8RHYxBbRIAII5Kvt7MPHtzWbmBLhHHm5bREfNTUwd2
PRux0QeLJh0SCGqBnIHMbNSg0yW9Y3nucGPHQpgq/wJS5re/M3VPVg1ibWwD
0seYuSniE1yOk9BuYwDEGWJYrKPVdYy41tP3VbZkzYIdexQsmCfUVo0NIH7O
QUKO2kJdyLANUyiyWz3jxQsDM5f9dfZeJe8nyVtT6ux/ZkEFFJOoZb0PnESE
eEHjfrtOTw2IP4WaYnvsMyWrHTgrKGYH/3uFLk94T04bbRJVcjm/iweJAsRc
wsTnQmc/ErAlFWWWr7IKlUMo9X+aXY0s7DDAVJqC5GMcNh5pDTzWC1aVR7un
0yv/M/zxdlKJCyT3+JAgE19cvOtdrKdQz0Lts9zurCqpNQkr0lPkZbuW+g2C
hGg5OHX2L9cjoJZnHfc6C0PYUiXrgGHaW5j5Yh4LCWxYlfvNPaA0WtI7owYf
twiMqubUgreZjYrHVNY7vZ36mTYxDPhAjeJuQauw/Lb7RfeCvUJ483JuP3fh
DPYLugzawvlQRmS7Ltr+AJEkQWGDQlTaWrtOw037wyawidzCzSVqo2iaPUdZ
cQeFE7cNy6MRmP1M4e1nbuYaHP1GTtfTOIsg0SkIxM0l4gJUQ+sxk0njB0qh
0kAyfjmGPs/5bWc21W3/drfdl7bNTN8iu62B2YPW8V3pNw+goRMMKlzQlE/D
fh/Tjd3CDU/AihEFfjNDo1WyWpFF0deozLefnPndxveXag5djeoxHK5nlbXe
z9Yr3YSHJ1nzcfVnbnsYxiHAIYKelsPNSOL8oQWeAk9fpHJi59T8P4mJ5ku2
ScPTe4w0w99paYzozywgsIjI0YvYdJdBAOuBUqlKCGHeCOUIxkBDBivibBKb
pkfRXbZbexof2P8oPRCssigF6GKZcVy3yQvIqS+sovbIAEaVGC9LiyksWRxf
FEYEIyv6UPfhbTLRmjHGNiQtu5rn9YaPuVQ+Uq1YK6j4H6UVdg0qX5K4WONX
UouxKf3OGuPovGjZc6gcX2Bk5wFGlyzzViuqUxWowW6WwuQYAmQLYqFG7N8n
EBGEXazwc6KzUO97IHP/IetRGadqHsl/FLKHDw/AuklQKHp0JIhvCnxXDAOs
fb1k6Zqhba6tad5VLdpnQd6lUt+O0Qy+MlyteBLm8ED6WDpOUFn7VmDxY4wY
22zQBVTmBFXvGGtsA9gQsdv3FUCz5Aw8zufWy0LnkFHpL3Jgy+dXvpg5ecYJ
jOVf50KBOytOjmRtzciXUyEuT7einZtXSpJxO+dzDAliy9OCWskWsMcux2pI
ue0E2namRc0KZ6SuHDZ/ctLHVOu1iHGRR/SZLhNhsQ5S8/6KE71HDuwVKwpA
7FhBjI5wOFTrQwapkVhifquGTRO3Rq9hiW0AUsGK1tSsaspXVY5Aee9rzjnM
SA0QuFzdWjI5zP/3cqXu4MOmRDSHViCyoIN0n1biUlbp9il7HS3LU6GcZbNH
amoDNijyCRmhyuyBHfxaSHV9qzndDdA76/WS0aTTdRbNTrVUHaa3cFp5uOG5
t2eYqn8S/PBtriLnmh4p/hLOOZjeSDqNaviM6v6ZxdBIsxjyoQWsvLKfAL1B
rdEMHRz5CHu7+8GXDLIlCq0kEcShjdaMSUqP6GunowOVA36XfDRQQ+ob/yp0
JtlIrs3K2sw+ltUyGmm8HMjnLYVVBh83Y5XzD5Y8YvmMbPWOImTbmzJuJftq
jsC4pK3CnU7MX8PjM/t45QsitCtNv2BwGRThVgkqowEf4eBKTTEzx5v/Vr8Z
AUOi43Wi6nZ/0zR+RYA60ZybjahwoUpX9gnA0LAxUjXTsntOgJ0tQnWJFE3A
Bb6LjhgVF3YWx0AnPjSBtN+lIiOSS4ePKZPjmN+NS/iMMqnYCgqmH9b93yvX
zQnFU9bbzZe1hWkAFRYGbHqfFIX2AjiAxNxmg99WEhJWDg44IBqPi7e8hrpT
txsZcBIqllotjt4jz22HwqRwV8h+JzgAq5lkEz/J0LjnK9BgEaJIMXpSLAIM
cuPQVskWmhTxW6KocUHElvINj4klMvLojV5rdt5ZSg+YUq7Uu4ku5L+IYB8k
eMalP8pq/EwUR8l6Wmb49TyEgeMwZksgMjp6JKTM1xXyHovGq7UClQaHMNqX
ftKlCqzojZ9y9Yyv2chqYPN+EyfyirkYsycr6XIKjRJx5/9A2UBwbQpPHFcc
1PA0o11/Pid+eSQYotcctYkheauRFzXRWlNKij9DTUWHgg3IxHfPTA/izeNs
6NoXGrww8XkDyH4wNTuuy5lEPnLutgbehmS6y7SbF1H09ix0Ot6zjvnJlFq/
xHc5vsOaAG56Z07RMPgHv6nBWpcW3ZbEkF//ZFXWrwIEakDnFE+BdDSS4eAF
msj9Mzvf5yJMAPf7vI2Q7K79r3+fttQ1GA/1EqtqmjmoiBL4U+ecOqcn6Ewo
py27n+aakJJONi3palBa4aWc2cYaVDjTLmTyvxqaWtI7bL3cxwCuZQCJEwUQ
V6FdXi45T1P7EmwMvyaZkoU6RcbrYlfOvCaRpV5o5bIQTnPm53Kl8GvGKBrt
WCZZ3tPcoFXiJRhtuDHR6Ym/Nvqq7xuBJRc/mM1PljtdYSNi/67v7XVCa0nM
Tw2hq9G7dHp+lAB77SDrRFFbDWYYwQVnBJFOIP+FM9LctkHO2qHf9kbpQhY2
8ObeynuPikBbRMx2U+iL1bwnO9Hva3PnZRw45jziAiQ8v+l1deBWaSEBd/Pa
Qy3JkMkGW2dChj4IGLKFxfzfJRRMSlZ1g+5l1TzPjQPAWlSbdiyeok5ppVej
pyjqEoXqASl6+4pvpmyi82nknCdDCQ6bUEqd1UPGtDIS7uebOY8l+7cvsMbI
o65le+QGPEuC/Y/uuHlxVMV4u22nVjk3Y0OQPUMwGc+Vz4mImPZTIrvJvcjf
5zZtlnoevoKjuLdBYSkQK5UfswSQqo5x/CD5/+HTL1k8c80xb5zzERkS7DeK
GA7VqX54Tq8w0KGPLWXsYxAahZZoXl0RXPWbVIxomD4CeJirx667QWvwTcPm
JW/BhSst10PuUIn6U6CJd4lqZhDK24Pxg1XH5aEGFx7oSe2anfBGy+48WLyH
81OsFK/zCSabotDuH1AnVTE3aPsVWiBE9MeRx35Xw4zwo6wT3dJXP/gO3yUE
sGl88XVPnTPg3+ZVj1dctUsDVLnSLzaqXlLu8F7vDZdwFNN12R6aSvsZ9Auk
5Z+cnWt21UrhQXBw3pNk4cap4z51kW6qKHIlDSlmBXNrnCT3B850mvCHAx95
pXH/hk98p8Tbh5SuGtKFKZtDBOXpts9dZzt4qypSdemvTLXDQrLCud7fPP9C
qMr4VFrGBX8W6cJhz1PiMmJCheq1AuvCrBBIspzF0BcHEBJWcM9Ql+QPEg12
UdAypNLA3Oi8jeuWIV4gHjZBH/bpaJ9PiPNJOCy+xLdr/YuDztaAfn1hq+m+
tsZdxu7P2TEEzEqFkzEAk5wFIBYbKhfRTCB+M/BXQhUjtrITrvsZx/3uCl/r
ThLNmAVW7Sw9Mh6jiMnyQT0t+3aoPijBWQu3CalOXykAq/o0GXe4cjCYuNrG
pi5Ze9uK/N2KktqWVYIZcZWejTchhfAUuUt9H3ZRnYa1x0ApjNMyP+JQqFaN
BLa7cYaT9V4Oo3+FWswUWrWHznGLqTahccXkKuDtrKMe+GoD9WCBxo0ZUSa2
UGDf6rqZqAmUIm+nrAfGsCm4IuclDz0DJ9vWtxYG/SEkKvJ9k39Eufj8RAt6
qxcW+aX97bkZKGqNx706F5AZisQ3HiaRp6cUBuf1FQvIskl5jXbJfy35PLDN
tIVswwu7+jJ5ZRzFRoEYQsdmAkT+Bvn2BxBBQ5Z3jXrgzzUCldiyKciIBb52
kv1j/jUOXA5m7KLYsI6A7H8SXm+B+eubkNJOWr42K06ic2R2GmOZvoqCRSh0
99Vh0djXpz46/qU7UjNCaa7WOY0UBQ7KJHgZMwgSc+P+QMFHqRgbhScUKLsS
gQ0vfB5HUlWagqrRHe2HGz3J+LrRnkAXZzPVDlFODukeuyAtVtU7vCnacfgQ
UX7YHlBOPAyuJfpMbPn32y3XiILdbHPHC52SgxhPamLvwIFPaXySxJ8f4Rz2
TZMv4PZPh+QlY2SSVtOXbuo23Vr9btVh4tZgTKR6uE7f86qO4I8BMT+5eYES
MwJthdhG97VhVS/hyY6XzUv+MTkElZr39uPsh3ta+oIVrQdWcq1XL7lP5HN4
SkC8pBsSkY/v5xsJU5UypGcZG8DHfFZX3nxmJO6cV97g29UkGjI1mySltihM
tVLrCjImxyA7uhSb9BzdApJSlruxJqyZJBhYt2XycqHoSnCJkpcJvjAQ8tSx
DNoCtb6gBnOcbpXht6pSWLMempnQKLUTYqu9M0+PSQp5nTAMd4/w8i9E3BJL
yVjh91VCFwpbiRlQoFj7A94ZwwWzDpfunCne/oKwfUeDumFnhWQ9+qqtTrpS
W3n3fuARIXu3POPHNdzTurShl5eOhXBQARCqzxWoEYb4bKQlD1+sDodVeZeP
AGtnyx25Jg1OCtPtvzS90dZ+pkcD9GiX24eLVVWVJlhDKraCxIxQoKNYVTgJ
60VDCH5LUJWbZX9LsqBM5FDmOe6njIF5PduQ4XPRAagWVBDldvu1Hu/x0H45
vJHfKXooJh10A1s4t7aIb10H8nWhrdW523oqeOfjvHfbOvEMXazJeMOpCsuh
DSZVy6aFc/dbkHSIZFD7tXhQvzYa/oCAmnUXAqqfsR40aa/laOuLdZyoOt1n
wPDQ4rQnHn3Et7ztFMj9ri8NGaK86GBIOYha31GcflWp+cMydX0djhza6u4T
VcKlVTlat85k2RHGp3eCdAmK1Akm+vbayWsUXcNam4asCLpTdKZcEaLYLJvi
Oa2Asr6Zn/eoCSc+lZ9fcsB4pKuHpsXtWKooJSrmYNH/20bcVs2b6dCLRd9k
e3zqmgtkieHlXSWTqyX7BB9Ch1JbiAs9Q238OXVV57dhtmWsFqv3/bZ2HDOt
pdVZ1HnzN46RWTQDnRGl4V5fp0eOW5w0wXJ4pqNtZl+bucmMTSf4bwgfGo6D
qUz3Anbcf8yx6ZOQRhJo5uVCn43UJNz3FUGb1I5bv6gt9oumDixTIV5G+pli
Uh/1EVh5vg6LFylnuitbaxyzcxb3p2iCZQa8uHOk6zSA6t/hbf4hvEEkSaX+
w94usaNgqF6JC67q2Irl7EkX3FA9+d8PTFeuvtxInca2WFPR7vq5FPV3GDJN
9DcmHtGJYrtAAxfA3xDG8jJniCEkFCQQnKvYniqdNXVy8IGXAalp82ibF1BW
KPMGGP0YH4INKG0qROUobf4QD7sDMgIP9rNSgBKB80lMESNHMG5eV8IctfgQ
2ID19yE1TU72qt6pvltJUv1v51xbFyzjGXSiCOLD7u5I7t5KGr7l2FxcCpmU
8FgbSB5jOik/+4ruXmGkNCYTrY8c8s/6FVHD+bC8MvsjEI+eH8L+I4+GA4IM
/9SaH0D2SEfIshKIzO6Y/Sqn4aiFrTqCP7Y3qVDP4Aq7rYJejRqM7uEkYlGU
65LULNul91LG1ZAOujiqRF9p7cDRLMpwaN/6d9Si6rSpeClBs9lbb5Hi40hx
9OzyF5cIy2rlyQksFg/YURpgCZPmLTlBURIoWdXtHu3JZu8cnVees6OoLWCe
zEmmdTonIoLdoUNGOligDizJ6qnJJjjNeiH/fXMVeRMCVAxj33LZMNh78UIO
bbuzDG7keZ9aphxOEhd6YzzaSvVR1gkMnNxZXXmMKtbyfD8/+hQTA/BZo9e9
wuFkB4avmRT1JDwnc9H3k6kv0kvuiIcINf+t56tUmnGJ0h1AitAA8Axnud/q
8UfUdfwtvTy1HG6KmlD+SwAG6guU0FLZ1qX3cFcKy6rTo5Yyga6TP4dzprfp
a3JRCzOkeyMyolBnMeMcjpFj6De3nohEPIboTh+oKvejU07zQfesDZiq/iHf
Gk5iNmtot9DNJOruMWZdDXQUvQ8W87UlKFDBIwbS3V392Sz4DHaPBUuyx0ME
C4qt2cEG8xO82oRkJHZ/h3OzpYqPJTzrHA5LT/5MZdXzprZMgChQWDUDOn7a
a9e7Vdnvrjxt3KQwZ6zqXJoN3ci9cJdGbIsC16uY/yriVTwl5P2B/71fgSGo
XTo/8A3Oab9S2uDhpo17QlPl5sAxJXljA8H8MXnTNscI0NwzSZEGxyVSSWD8
5W4kEfljCWjc6hU5vGxVFAWvKxpvGIIkMhGFW/sh32dSH/+uYc2DcFzoObCF
Kt23A23TaNnj34yy+hTxZlWEf5kyP3bc/4AW6vrkEILzbx8JCPvKRvNJHCvW
1cCmfy7EAtSKtGpgXDBc5cGXGFWpMmj8D6l4klDVf+FzYj76viWNhtygVNah
dXYdRA6XQPv07FI2Nz0Al7QrPAczHYkw36OOPb8coke4WTggBa1bSflaN0BR
zzg3SuAFQVWC2wL9i6fphskc6sWtbuzJVYOM72H3T9kfYdRQDU+O9h6DtDYH
eOxVG3WxdRn9M9nvXaSdJLPZdVAS7pQG6EW9Z9d5Rf9NrulJqml0lYf7UIVw
xbm7pGhOkcpsD6IHHfRv01DRLHmstAf8HCfvfm1LFJt/TBzT2X4Rh+5o8iT2
dj8DH/eSMnqdyk+WSHXz2y6sI+RZzUpCBm8zHdqV/H8f67f2wli+lFTy6aFw
szb992v/WJs1M3nuAe5TeTxDWmpEOFTNBBhXwDqXcE6zLhuxRkBkEZNKiFJm
Kd3XIfh3eU+1+bNrE8G45ANP8tpJngbKi7PJ18fvQ+xAP+bSyZgeXkivA7lg
6R3rmdzvbkR8uJQJkgdKRn+WQSp0UwLlIAWA6dK1EFsQUDJKMY2/uJB+pv7G
j/LrSFAzHi/8VsGa+s0wsoATrDAVTxOgeupDqtZ/JpRxxpWzT30qKuVe3w1E
/xzZ0T5EVqNTILjJwcDwBamJN90Vao9QIri6X22QloSOGGPmC+RpcoK8/1pV
+MCvYlpxVw2sALaHC+y7DX38/RWcTMNrS5KQhUExi3hWBoTfMnZoE6v0E+sT
miJ6Gb+YkOySO15TGs3HcWyJtLgeeKEuB0UvTJNOOHSqSA6EmI+LaIJWBKWS
iKsmOeU4mCfPyReQy+GJszZPXFkTlIiKLj4SZ8TkX3Tbf86Pw7epzQvKFQDW
+e44OersjescLcW8t7Zv5lQOd4tILtYQCACCaBfJ/ObS+sFpQv3N7lFduZFU
iaMqO/Gpb7Slp0xD97ZjJlsszqOVDLHugo2Ek1O7mdl8h6G1A+frrt5BHEI/
/EYqHAQ84VYXSsmLx3lzsKEq+QIchC5bez7FhI89ic2pbEpYYe0wv8H73xNZ
i6T+n70UYY1Fqb7rBQsiDXlYrm/Pdug50BCvURFTngbyCNXDdCG6Zj8YVFJ6
nrJOmTBBVPDjOJ/MnMVZKyj+LubF9ldlrGXudBt8xizic0rwsav5gF0ZKxB8
e8fiB6ylfmMYjPPTi4bfJ8iUyKkSOIhWVasO2Ymvy7+7X+9wwqxawbQkbU+7
kKY/cPdMEVRzp82TkiLyrHJeTpW9Ldg/lBDHfgt1P1e27OxkhrJw0RDaHzeq
SQTAzeKF11KxFQ83/bKswvuRWoFmzMd1hVe2RKbb89p5ZjGI//dl9pY7oKVQ
/dzE1YNO0Ox/YYcNPxoyFzBUS05KEzimYnb/aHsv4C0odVbCM6hj+PdSZQbW
lw9JOeUTXY9OypRkBHze3du47Hy/UqRmpbzoxk9xvPO8Fz2E1iJOguCG4PZ2
2YpT7y8yxsyAzEa2zGNNBBT+CTdh66iV6kj7T9mFXF+CimZWMD2bL8p1gbgo
4v+c7ntin8dAPG+C+wVf77T/d6ng6JX/SRvafxTMzoGIqWh32RIoNw0OA7uk
0BnhfwWBmOvzdGsfFsgWtAIyoa4G3SuR2krAIJ9fc45qt+mtyh4xb2tSyRiQ
76Jhc2L796wjOR71I0HdWW8H7SXfPyKhgOeyPPis247Tnp/8OmoLWVP+lMNP
+8SwAcH0QNYbxkJdZJJSHuJXOyBPVebt2LzkbMue404gTarUvLhf3ApSq24v
gaWxnRFziKgAzvsVM+lf4sPepDL1PrUVEkurR40kDleA3VIqaO/uSt7P5L7c
7VDb9bDho5wvbTAZx+BtijDtHVmqKrmvq7tdyZyCnT3sQrB5qAqRKGW2sV66
dcCZrbM7wG9KhW/U0qpkMEKnmLdWjijEIy0L4mEUG5fW34CB6Jv+99oXB8e0
yp1eN3rG3fDMyV6sqzkKM9SOZNi6vMTrtD2IWtc1yyLF/JNs2XooVKRDxkRD
eYzLb4zODlweC4BUmVfEsanPl0cOju11tKYJNFF9WPnSy6Kt31EPzOtJEZ76
DJujiocpDwF1rsGyCuaU/aHbHdwt9eNh5tAkpQlcghTUfvVFkgAGjrAz0HKu
K2H6smyBSLhUwdd58dZKpoe4RLQYU8laWkO9Lr0kLJhvsUTjk78jjY8rBdlA
GSVI1TU2FqG9LRsvBQFv1Er1kZOn3z9LfDpSTMRC9IWohvfhW8YX7BeLlrE/
hbqh+e2XPGBIJkLx7XPcMO4ktEI343vD9kaoTYSe4gbabe0J78VG9ss8L+rn
njL3VLDTgOmkv1tWKYrEEaYulKbchDh0vjYoFc6IT14PiFZnaNt84h3zjyHW
g4T6HC+1SGkzN1cHxPdbZ4Nm3vyiJzDsapqWRA7Ehlu75iKnXlEAFm7Jx+6f
J9ZRjjxrVADVKhgUfVgPF+PYRdcX+834omiNMK7ca4lYhqqV47u8Hn4vX4wH
vaRo6QQm48K3EDMSUMPDGj1YNLU9WCEJkIXXkgMrOAS9v0qzgquFpRbGAqvq
TkrOKi6kT7RPGubub6ADVvKv5cCEAolwHXmllRIi1nYDu/Q0RmcDEQhZzFKK
XZw1Pyr66nOBKxQDIC7oP7E1YlbuRkZNqzmKGr6IK/bcGs6xhfpz+tKj2EZb
q1clNJCpZC2GSM5Gk5bYSamJH60pntokOMwH1E+4WPaQfPBDJOGRmDmteZ0k
GzExWH+mzOLAhIh0iBE20bVwmjvdb1jM7kCsb/8eQShQKoFX0UcuorTf/j5u
eA1eQiNl2CBFCgNDT2EjnB8L4VAWXzJ5k/3kvFEo3qUtWkoBZ+sEhtvhmGGM
36jmp4kTuXg4MvOGP9GY+w0HSitKwS7wFyG/b1gBPAQ92h0V01cy9WK1uTy/
raJFW9Y3vJqEwP36k1yxoHE9KhH3gvLVUQBsrD2nxjbAlZIrwtdACYRQ8hWF
oifIVNifRhL6aIO3AiuPJsi2DNk1qz8+5h3W/vvVY4OkeTEx7wilHmnY6JtS
Z0zx6GItKk9O/q+nJ4iHCWL67xueTMRvWXU3xE7BBn8wtcr/dp279bEVXyqT
N88VGTLvCpB071H4NvKm4d53yoblVjAiG2KsxYESYqhzFiWNqR3TEiLZ46dQ
riu0+UDbvyLxJYwmAohjfV57FgeiOx5o+DGIoTaFjB+zIBPbqmVIJcDebCS7
1nYGl5W6YM3Hr92ro0PFfA9V7K56aVpJneY4zlpp13umgZJX12IvEAcl9D1j
t1YijWJu5Z+kyy0MWFxdc0fL6l9xMO4saMpC8rmiBHZ322cdp+JWjDF+CFUM
SmDHN1arGih8tyvlJ5YwKbgs3ZrBQwP0q3HPp+RsCrHIsB7Gy9j0Bl7mUQHf
vTptLYDqyf8MKgtguCEoriuHzBnzX2L4XOlp/HB2NKKPGl2dzznM/kQqbtKI
oVgjQRT9/tgsVR8bEwVIlCxB2ky75lO6d/swcWdAZova3uO/eUKHIZb/9y1i
OtUTROpB4rZJYDywCsWeHSqLfmSNe9vyr3xLNmLaQSlRyE+bdvjp1qxr3UtP
dhRKekZBPAEUudcxKTgnxFeop/V0atDoK8tOcGvKlB3tzrdM8fLyvOkZT1Jf
KcdBijMNjh+ZZUe+hyI+UKKVu/kN3UoJ391sMw/HfmPSjxdu9j3ygcBn2c1/
LBMhCJLGwcgTb3mrjgtI5jdu6tv/1Hhv/eZpwfpbWeWY3a4/B59Nfw3vfMAF
F4IpdNUmBlzrsePNfBoxsIxsfU1qRawW/54yxJfnWHywqvRdOZx/qMh4zQmF
HI0WTayZXkeR02K+7Yv7hFlFTOh02qQH7Auvj00IvjzHlSrS44Uy/AwhB13Z
hygvuJRhLcput7kjsl+b1llG27vTiE5X6wZlvh1K+a6e3SIYTCqaRi9uuhoq
owtsQBQscBYyDs2f826Dk1tVSTVGn9TJ/0rMjET34CtdLXoW4jCC7DmNIFIE
m11twVowsrvbVhB/bj8oSKBKV5gOOJ2F8KSRDifysPjENpM/1Dpw3SVS4m7V
yt54kwj+avIkVPl7RebQH2DpoPWlu+tQtM1//XcvIY0AmhcFNDPxSxIhs2bW
HHlHgDqrsKjAKSCqvlsrP3AebLooErAHFXyzyww75jk+Fu5EkHDg2Ur6F4D7
m85ogWBhAc1nwBTwLG4F2QsET5meXyFJ1eGWi5aX+6iaQZ5MQb8NS+4hKmOD
uqqy0wU/VR0h/WpcCzuTkW5Qo6jJOtM8qCuHwJoDiSJ1rJ2JadI8T+QeEAhk
fgOBZcfWVa/fyZrJdXJCtIqEicl/OVzxVa8YxqhCuMvOpEVQ68Xp6e7mx4xb
id0+Vf8p6tt+mF7sJKkp0JK/YEmICm8s9O+DO3Adqb8iSMhqTnBSHW8SAhMT
1m+tncTODIR0HYLXxl/EYOfGsE/oFQtePqabjmnP8fu492z3HB0LU+QDXrxk
xT/c9IktMlnRM2bOSyKezgAwEgEKuvtsvYvGd5/zPsqucgBhlqmLrELZSUx/
84zqZlF8C+so2chn7t83SSM9SQgQC31AD5tZ7jQHv/VCoYip2v2IN8s9iEkG
+bk5pfmp1pn3GCsI1Cgmqb7kA9QVrpmNJG9SdReK2Ae1IbUKZ1rT3wYhV8Wv
M6dhegfRmhNzwt7+nYmOlJV/ZkL2u1ZJaxra4J3pPRECKaeTfPqFKfbP8w7t
i2EiQ0ebCbdes3KMod4r0gW/1Az9sz0drAyURsg+PbLRfai3GnrAl5SgDnpL
Ss0locolWTchvpaOEqTXeJPPHTT7b1avcbCkdTPetkdbVcsSikgXS9RsjD8m
moUEY6ScP7iF5Q3fzBulfifJtsF1U5lTiy0IYaGfrJVGXOtW/wdRtVcxEDit
v12HLt/5rHfUWEwcUm2GhPoFvkEeqDWr2A23iH8JcOym+j8IVTEeCUeUQg0m
ZlxGgbW46u+Ur0aufXuONd2GzMBVHFWLF0P+5S1x8X0MmIoT5Vuj0KBPLIU/
syeZY74FjMX9q2uD9CvsRiPn/CkkV6KVvoaQ27WOUfbhQocb6TwcrcUL40w6
F+9mZAmer53dqkyC+3p+xbD5vfs4Ktev7U2cnua963y7hZ7ifj7NzPJxs1js
tbtHaI6IOs0HPKOrIxOkidPd71ZblRxNSvZ/bU+qk3RX7wNJ/ksxC9A7Sy0O
bEelRgyr0/X+b7gEjb4jnRG76mbzk9k3TFxhdh244csUN/HwdocCcA8Ifm6Y
33+eOLl0RU3yoH6UDDIthsSKT5rh8YfMvAmgl8iqvmR8Dc5a2ilFguuJp3uo
9GO6kuCc6hP8HCNZ1RU82SQmljl0VgYOC1PZ4NrXC2/mag54ihI8KS8u09Jl
Gbhn0lvntBV6+vGvDr5s+XDAoXIM1Sk9tsYyg5NCJRUmQg+yplSPqTNCanmR
N29fpMS75e+Amb2mg1VX0xdd29aodD7DOuQ/Za5HnPO4a8urrts5cS+qWUgU
DWfMFjBNHMWyz+7YwfBMA6wP283j3IaZysQzXdu3aPNBO9ZgwJAdSIhkl8BT
LsVri1X/YQM77uhZ2pKdQcXH7VM7+DjjwPrF7amqQyx2qGtGcMi8rfqDSHRX
1lh7DSTycqiBzXveO/wYPUpcz5Xmwr5GAw19BaJMbut+xAzADzvR6f/p+QVD
9ADvkcC2DyPWRhjl1x+CsXSB4MlS8VKFCdmFk/s3O3VYBkBsjw9ha0+ykR9H
4paFHFFBWlt0MR3xRQ1A0e6cSA8qBYnBcRxkPQ0DEVn7NBITRm70+7uGopRQ
TOycx15Tf5nRkahgy1oxKjTfqYoC1+fiunwHFBj2De4RvZV5/rRYUKZrf3ZO
2L5r63gHL4Hxo5B2Hc03X17qkXkSw87C3Be6BieVYwZHepLpOJXu75eFkRjk
jVHCnWbAZAgfg2bICmTKux3sNyh/sZtZEaYDBRK+gEJQ1lNif5PpkVQ/WIJa
xi5q935dwITTKRgzlFLTe+H7RCxqKkgo9Bi20Qk2WuaFVr2x5CliRK2QXXFM
AkE1nDIVyIbuSKLD9UNnAmS1ATog4a465qdCMEKEVn5XrILuPYL2wEuxY3vk
UXrpsTnTc+dJL+gHaJLuS9E+Bh7Xa7nawoyejEcNIiIwTt3RpyU3eyQQ7jFJ
mNZ2VyWCzjqCNhuVdIJYBSXoaqBl9ZCvnFgMsOU/gTYbXxf/2nUMjB+Iana9
ItSkv4McZEqn+D6f0PfsDALqrmzoCIlrXsPyKTZDeTABrWiluHckSb1AsiKW
dedewfeGLKaQPZEzVSP6IH8cOeHt+k7dQbjTFOVsBg/PFghw5CgWgUrGUJuk
lTrrljY3GA3ngR5FGmcSwjtNwGFx6bkQVSzSNr0cvbdilzPsjM55+LDzMahB
hnSqfZ722sxdKdaCro8KcdQ1PkZ16e3yAWPHEabATYwFshWsblb/PhcfonL/
+TYeyBDqaTmso5fgyrYzQGMHdDpdgDj1tP8wT5ANREtNGCql9gmQEBkO16fq
lGbmxr2Givp3TYMtqW2dF1a9UeK66t9XY71/D+5UBt7+uU2Zxw+iwSOzj4WG
67kMSuwPpy4lOgh5v/r8usOo5LblCWanIC4HJbia4HZvbIeCSKByptidbpvC
pfkdfyqU4OUqfXnqUllGKCMXnEJOQqOVfH5mXInQAfuIFddGshDYsNzki585
wDclT+oC/W39vKgivtSSiMU9R24Ep1EncLUwi71lPetrEwtHld/nh3cdHzZ4
sJzVQTGH69l50thUis5hITHoFJ7B/uJGMjQwQ4nEYIcBZJWlLdf3jMSR5uL3
zdevuuEMog0dwi2kqDW1St4OSbrqEHI1JdmBCScXJoO0ktPbKsUy3y4Kxdb7
vqXzUs8N8dv1XU01KgxHEFR3fayRIQztMtrGpouMxfRRgfhBO8do+gJ2NLUB
TQozJaIirXE1jLugg0qtHCmjhtTJX0b5FHo5iuZiUZlTSOUv2z7pDDhj4pwn
+4qC+kLdNSYP4Gb7zLsgiAqo6iUfe6GqtdvWXLCAqAEtqFLxKyRvT78wKfy+
4NdZPdivuDtd51K1frMOUp6UyXxt+NqiD70ztAUeER4YfOFOG2mP+MRg6cwf
CvN9TQv6W/wwUxBxnQFT/47k9K37hQKEO0PZYeUjuOfnOpMxlDJKugH0UWVL
yTGUw9jDUaX4zJTWpSFIhE6sOp64DzXE4H3apLXocq1qXKkuuIIQdpUVSJRA
frRH1UK54/6CctXjD3kcS5qXik9d/fuCCn3i7hCvHpFOzavjXhpnp619SbQ/
s813Pf0Caw+qHjYbNYWkit7vvnEKfpFz5oMVzogyrgOIfv1JN2Mwe19A02ym
1K/aKXYRPrSQx57Yjy0+/rH8HyM4H3442BPEUmg38ya7tGd/bKPO8cZUNB2X
2sKxh5EcaZNmP1GfcM+BBqUiEY39LKkDYUdpycPD/J17o+C5T4WRoogk2coF
3A/nz/FxMWjYad/kjW6uLBIPnHgMx8NV/CCT5gaCxz8ylKtyOhS53YVNrMvI
Xq2zwP/62jUrr1j+cO06ZRXW16LKf36wyrgquIu8Gsp/VWiP/Og6hP78aj9Z
dVjsQfRNoKSzoEC7dk1mdUj1Q3868GBxwWkg15VNEzuIA3wBczz6l7CKM4YB
EFppT/pppCodvKVsk/AlI1yQuqDGgKk0i5ZbODg58NYVZNkY/s42LNovwqwo
6XcNZFPzVhtkay6PRaAc4KO2oRZX6Mg4Wg/XLiTO14GScbuf7xWOqPBvr6hi
vgg5QQox1dFdG/l9Y78qVGXQSsJweJexgfZeLJlx5N6UVb0scb0Iccvn9b7/
WWQy/i2lhO3GZBMTO58quaDLml+0lGsNIYvNAH+hxaKV0Z7P58VWFZIsMg7p
WVVR36shKaRdH9IylaAdOKlbfn311YE/VnsLZm6ClXzs9YF7/tjJ8K5Icxw1
gh+ZcybHURNkhS7hnJrxuHJUkRHZjz4/ZxBfcVrR00DEfcSSSIrSKMs6JvEw
+g3z5kfO3j2Fii9AfEfTYE2aXhwMJ7yFTzH5uCA08+2nQXBeiE3OgPHa9TIu
7sgPGLAuHA8MpfYsRJzXjgWZhq6vh7HCy8LTuzM3WtnNQJArQORJ+ABI+Gzd
WWGNO35WcqcqdO+LS/sP7VH0skyiVs3JejFcMfwOMDW0uYOALzR6LjeJdMlu
hyw7VrpZMF5cI12ptxs3r6U+wMXCFXxCoJqelY8QU3Uhf2XBwNgDv1ZbVOM5
YQYU3aNTWZpLTvykcNcEEkINJuimmpsC4uEN+t1omhy8xVMTcZ6qS6cI32uI
1qj3mEE5QYWmVxXImNP6Nk4ZfKDB8+Vz8n8RU148tNizVjalBYwCwRB/i256
phXQKbykomqPGx7DzKCAg4+uEU++st6d/wh8exjluuQbjSqw8lug0quXnnL/
aoK4PID8wcymgwiO4WdxaGBnJxInRbvBfjQca2ZK/YRmuZJOpQQrTPli8Pqf
PDF0KAYS6bTsIy4oKPyMicFcCxXGzrun5DQLxmRPgRAu4+0azhDtVJNPXx5T
orGDl+mOHYKOYlwKA5vtG6JU5nlMt1atH0zC0D5ukvcbBphwuNykoEHbhLus
xKkWeWBn+VwP5WfJZ3/XCy4ibyMf662fre/UQYeYZTwdya7RtUfxet1P0Z31
nA6n2r3MzEaKfYOrtgztbUMlNuGrYxdXa5L8wqse48Foj3AhsrlPntD3ZaAA
wrqrO7UjgdNaNzyNRGP7ByFWcdV2ebl2fl2OGZvShE8Vq1dKrh2yYFlF/6cs
mRQOlIaJDdlt8KJP2H/nEm3aDAvU/C65KQ7XXNKA33WoOtvSfgXBwFmsqV6M
Zvxad0pzO66X88XqNoxxKIQhNs7jE/rv2aiHMdUt1O/bX/eHwiVRyLBk4IYs
Ymx7VbP4c59++TG0hkIgue9wlJjEwSCO8yvjK0dOAd6hlyCwniPVGVkgzK8C
2U6zUGSGO6mRNrBHbJeN+N2nIbuDFIpIoHkJ2DFcCi6zkBNHC4SlszBAiiuu
0ic5ZikgBahFdrxRNqr0vuebJWL6gby4KOBvt2hyy8WYEw9+xeQniBBYHn5j
ISKwxu0PFFC/23b3ei9RjFnhbNwOYzMGEhvbWlmj4Aqli+PzT0ApxXFjmKoc
44xncubdZhs4jUg7t5yi78rHZ6unuWOii5vQuY8TGGfKxQrceSLupMDrepsD
dpZ5oeaJQ7rsfbTqjHyL4vRqaPhOJLLRhCWv4ChuzJrljRxxUF4nQWTR79ZQ
IXTz8cZNCE9hBaRsU8OdZ7448BmmGrZN9BVcx9wnx8Fd/ktRAYDlHKX9STTu
T3kNFqqL6rUGkIEVe9i3Cprn9sJrBxDcy9oDjANlHUtoPoXjXgv/YIgR5Bnt
/PFS/Z3Dki5hyLGm7AfGcsgeX98RMaoFm3y81c8+P1Ht8I/9zQoxehKvOyXW
lVuB1kyurOOTpEWtb6AU1ej2/CBhr6RuWBBtQQwphtxYyzPmZbfHKO6v7VuP
e6l3MfvGP3ot3L6yy+WLJyqV0lhBB5A11W5Csytrk11zz9JeqF8zwbOh1Y3t
inmejqHYMxWIfvIr5i1ig8LW//4l8Xcw/gPKT4XebylL3aUwerhBm2KQ/j19
NcW65aL8TSkI05fOVT7agmpriye/y6EqsuQbgEzOqHZS3FxxRDLuhgMRUjIx
3OyCtZASajPcmyM0jrhF8xREbY14GO10zsSZ4dgLijRt6VZptUKMF50ki1EL
xlAZD1PFWKYcOwLE7jYUxKx3QudECcBnZc9pMdyafe7I/YdV67wzxcFCutgJ
yOD6mnzvxJK/RYM9I2sU9HXdPEIh0VWok9Ofybugfg3yATPjm9SBaSrZ3oYn
8G7GJRpvsWGSKEgRbt2XxATNfMJciHhDk/XZBiQVnmSyrZF0nC9yqS9HllPA
DITbBbuWN0lFvRS04foJwzh3axNnP5okA8sYUYxqSnoUC/ZZcIbA/kqBIiN7
Suxkd4fsqvrk24NffVY0/+pk6WHx8j/OgbrVzHGK961sslSeytWIFPqVT8pC
NZR+RRWBlJJ8LAVsi4dnnoB6OyVibVVHqKpEFW7xcFDgqRc0Fz7fRU/4buLj
aQbR1EQOiU9KBJYFuRFb2AgYxY9/711mgcgGQ0qQTrDancxa4tUs0at+PU5N
/Gq1hu09F5mhgJ+tEkciBIuSuVYw9nNXuAQFCxyrXT/xZYpr+b0vdbJaYySI
DGh1dWKnORn6AKGNZn5vQALF69Moio1+fyCJpWN3rDENQ7FpRCXwyQMC0gNK
jT7VZK7gAyjcYQ38atGLLuqT0LYDY/PbpC0O632urvv4Zw6djaXh1elvghjV
yv3Cj0iCCopK6JCgPU9xkHZlEimUuPs8qhP7ZuHpE0nkon6w5TPxq8msydKv
DXcCvYMiUo2gzrKlra7lBt4lRjQWYKJle9YpKUADeZCBGVOW0Z+5phtIhfjr
c0TjM1wIrQi5H2rhoIMs2BmZA/Imkniw87J0PoiI7HDM1GQM+qvYpHYb2mM6
psI3crBGf97ZZtRuF65JANvH7WhqQi8CLcXByne+vTqanSq7SMGFOdUQpHyj
dqGWqseWPuWRYgdw1glJvuEvpgfhvY3Rt9gpdt1Ss1RKekVadjFFDmvIB5sK
+qikucrvTZHuUdVxCISA+3WOeHfW88h8WdGx4mrsSLhzsB05r4WJ0OZkzQbq
b6dU03Tq4zHLKVQJw+wMbVTURr4GwPUAblSW/18e1q+VoUPcydEYWoV8pjZ4
3uXD0Va7XzQnPrd2peXNcLmCAZyEas7sccHKGP6hmQI0AH4bRo7AVTN/WADu
BZzgNRALf0qEvIkkkktC5uC50B5ubNe97LxNFTaYT6xMrW2kX2Czl4kWv3mU
1K4sqaHrbYIW/Zq4+E1gqLF1kYQ66mcTNNQzrK2sbhbOrxTYKDoeg9iUaLuE
2z9ZqbVjjIXYPvA6c4W2Pd3xyRPEk0m/QvxsnRVpjq30hi5AgkV+/VBFg6FX
cM/UbjH43NYbjl5mPFMK/ZWN+G1p2Y6dtZdHqV1B0560or53Kzh/n2JMquL9
e7BFgrCP5j4nr0riMvAgBfMhqRE5kJuIcmxoeHLnqweQFWS2JkChxYVS1tnp
fL3ejTGPIBMOiVjTKNp/YcEGL3r/kaRKGnM7A0xjX87y9W2gEqfUl5O+LM+W
pq4jqCs63N0nG2JonmkNdIOiX+YaHCCJBLg3DUNh0GNrOsRiVJ38ai13RgkV
klDFlgSQrlPiai3exF5pK7dho/WGmd5VRdRGN/dtv0G4BXpB+HqWRPlDfqwD
rMwXs1Q5M7KKvWGTzhGbA3t1W/5facq7g1PcSEw+hR12zlhnZIpAncPx8SRM
qJK8E84+K1KAzo919ny9WD9YVt2OFyFLuOuENlPOLnBKYihyRwbXik6CrlXc
dM9fcOtoBVv6Wrjcgrl1NmvC7R9D4f8iMJGVooeOQAiX4r3SraEdJj1GJEA7
KbR4vVzSTI44EaBX03OkEyNBA+21M3r1X1x8r+iL9xsqIJjUim8B69vYDskC
xQPHwplgSAxvHHktmsrBlo+ckud/oW9cQqJHttE3sEG4+ioZl/dHlEhTiQzU
buU6oDEjbvxRP0HGzvsyg+YYfXhbZ4UAlzT1WE0gQCU0Bk+rj57RN/b1yO7w
WrqkwG01fWHPC9qo7ARsZeQdplQg5sLsggGHxGWz0ipNW8j/lVWJzJm49qsc
bJkL5fcCV0SASRdGGtNOTXdK9n45nUDO/BP/Au/UdgZFk+ap5kL89voFHZ9Q
tZw+C42dt8rFNi2RResQ8dnTfAJCAsMfTOwlZKZ7rnQYUctQiRTIzfjnGGed
qGQWVGYbEOW20KICLDMgdgMqaR2Cx/3eekBHtKBO9weVgIp1fw5RFyv8siWM
ZaUzrw5jTXx9M9uo7oEIhqul5HoIvKZVtUHrj73o3gcZzEpjHHrVK9l359vo
w2y52aUAefA3GFyldjmICFGuNU9N4RVSmGGCcFw3mn8Z0SHZXXzpgqG/yxhe
t32zYdRlkXQgC/6gBWPXukS6bFICE9gkmyDak1IHXvbqi2fC5/uzZf95vNZS
hq+VHGxccMzGG/zmFhdd5yMSw6ti3EXaof0OIg5KZYfHrTtzCVFC4lEKEoRC
x3Ty3hRKCvuECJYbFsBy/ZYdJ0Z3TjG848QwCyUdVMW4pAC/39FqOyLX14TQ
V3Xo+MghPL0gIytz2YIQuwWiipDadW5TJT5bLuo+2Kdo2nH+BEn0unuwvlmM
uYPBWVh3vPS5tOT4IkOO2MchqmsHWg/sCJIVD8sCt85wSppzbp/h407xZUZO
W2Bx/yXayqiqDcH2snkZBjhPe5XZBjihzS2BnHEcP8l+fDDyLfwWi0Q8UQ1N
ifR9Xw0DL5fbKIA6CPGt4PHasi2JrSPjp6YQSFj8YvSQLXOkYCQi2WKvPDUs
KsrGprAOOzeH850RkyaJ6qoKSZMgh//GXZevuG3pZVTdAATq5OIFSXxb0JyH
WMgPqdByhTgjm8vYSmZTHsFDwsgnF/eN0gvy9++PPHRWrlgqqitjY9Hyco05
2BcLqNQVYdiIAe+Hiu5JbFvS73o8gmElMIP4E2lRDSh+TfvC4MZdAmhCSgi+
L54w0BvTsLWFduLIL7CuLaTWp3GRk/JMVUGVVYTG9o2FOPqEX5ngmV1qrr3q
nfEDK1R52rSfyWR9hLDTzcfKA/O+YoBadiO2tehSRvaG8e1FDY4h5YEqUMMB
sutqD4iXBcDc9jOW292fhlm04JccgLmRYv4Iu+ciiPgkkJxfZwo35Kj0oyNV
cbO6Rjw4FTVJSg6YtS7xQnJ+B3O6352ylMIijGsF0/MKfbqUMglGSsIoEbFO
XLB53bOqIKT0ijpR3VnWa9SiR7vCGJVI8skPUrFnfdTzWrNIH4t4Thahg+xf
3pyVhK+xF5odUStY2v9+9GliYbllgDTaYOe4w8AD9aZtiwByXm/dOFQdmRvr
Qp7ERe77OiTrYLo0T4mrL7KeCrCF99K98eNL6asxEIiGaBg7QMpwUJxhvxaz
QZdY0Ngy21Ml6Jjmk3+7rRUsp52nwO6q4VEWeM30PEM/sKYaZMZzpFaxisRu
PIaXI4a6LcwsA3Fy0FDeRhn+dabzNaTPgExS6WCcMPmvy4ch0x5kmTCr45NS
AmXz1Mq0AvzeyOOalV8riEEeC/ucH7XT5wWBzbj3mJEA8pX9JlGprgq3sfiM
rJMmTu+mz8nJgqZclE0qcZbRmTjOTLp3/DoM/Jdt9QGooHcRczAN1cQrMwDx
qxEOadGr9srVKMKd6u4XnO6GBrsNkgs+QfbI0IcOV90akBfIOUUu/NWDUrn3
/rgM+yBAaRBemmOogIqAtkWK4Pr/G6JFusCsfLlNnUFsd358iRzHOpdtuqx4
CPNgoDTS29jP94LYN4fUjgcxeqxT1mqsMcTVexJ6SeEukMhh8OHjWBDmD80U
MNY6Kj558whJSrhhtNiHSjw1z1/8v9AlY+4N7/P4oVXcbCVOncbHP6rYXCKK
sE6IRx247S9urwsQwwEczVEgsijYmG5JXFf/HhWddxKohE8Fhr7UiavjdEF7
xET8Y6oDpAQcbu6efUBCnq5Mx2YM7Iv8J5ThpH7yohuRBMS6GQjt8GuVDalp
mw41b3a5NhNRp4BqNW4JW2F/EkbeAbVtJ9kLAUezZC9BPjdKux100KfrzJVR
NptQR0pApUWC2ummPBGE/K0FGkvqkhFkr8SL4aQGZoSlfQjOg/LA5Dqyw7xb
4xcUW8mlw87MCj/10AfwQXrgkiTyr3Q5BhMsh4sOY6DgWWxdnqatzE0REmzz
lMHETMUE1OrvUXRbsRho3OjdUOu8I4Qk+VfVrsPpK+MtIgbrZ+XIhMonkypQ
BtBtBetL9XmluZkdGacsSN612iR4z//sTaYkOD4L7sV6FjNtl2q4vo6uFxed
GoUNHwMY7YCI1+jq8Cu/crv84JZFGMV5piz9iWjoB8s6VQzoqlZS74e/TIqm
J6BHRfE6SoZ0OJh/FFZ3Y4aQto9cfqvs8+ne1GzGngEpu6M9qyUjfcg5+BxR
08v97IpiQke2h6Jh5LZzxlbRlAAs2OF4LdY+MBpZDllGxVAgRtM1KJycUksL
N/n/Zah3UMU8IT/6Spy61j4f7YVOZXN9PSGigZ2g8FMGipWj4sQ0xADLwCim
ujhbqRpzytM4UkceKvTPRXOg4dD5T1U9DxJKxoOMcWdbgCZVRKKHeRwtmhdv
yFbr8dS7+j5nkIcmQy41cEe8czNk8blHUK0cmPERYJ2pcJYS3xaKTX60rBpm
zQRrgPcKeb6cCjgLKksg5Lc0j2WT5E8vfH/JNs2kPlIkpkwqPl3C+PF8McvC
k5qIpC+kjvrU2XF9gtcJMyeOdToMrQeagvahTYMngJryMnqqb3w+U30OwuxG
hnFqgPKVr38KI/DWycmZ3xTSv1iTwsIHUeq8KHPxybH3iZMW0GyQGo9UQiCi
5n/yb0SvRKsYs2d4JPtuKg9rcNfcn4NBn9aPUOVrZCoJFSMFKC746C7hrSWK
3UHY3A3vq/GpGzcNnmugPzYPRaxKEhHKaLumaP4jDUz59JR1fn4XcO9TVYFQ
dmMqL3od+twhVJSPbgxG0KA3wpTsQsJywJBYrMZzHGO9s3blMsWB0Jr7ebuv
Oa7FuetC0Aam8x50BA+RQV1T6O/e6Q69WW4ed7D/bBYtebcW/M60gEWp/iqh
wtzaAxjorzCUbP2n+PzD9Tw36P55dR+wd4RQO+ynYVWw6mX2Mn1sdlrrjp4o
5Y7mwJ5ajk6/rvZZWPQD8IJvDWHBbulf0Cwwuper49abqGElc4upFKexHHYL
9zsUplAveeMKXbGWeOtM+HhvUo+fJlHMkOJNFLFyKrIedrkHxlLLpfd3SapW
l9nLXJoAkOu9xGx6IN7Phcd4gFC2OEapcbud30TPYokvONzTH8AkYKN6a0kc
ly1wr5NPEmIhLoqGAvTWNF0iziSnfPRmrsSpZJ2E84MWZIJX+UHNK7YVuf3Y
Ivnw5AgmCtjeZmzFDi6bYRJjLxgD/ZbPkgNGVfH/Fj+7f8ZR/6+5pdPepYUI
0njLyyD38I3ceJ4eUfoJHz2SG72wdgKoIewN3uC6jezSdXPRPQLlEpJ2UmnL
z3tYzn3dJBswpMmAEorQ+PGX1B4i7AHhQqaJs3MXhWs34FUq8vOjaTekHvL6
ww8AevwTCFfmzNXt7Pnws575XEpfruVxISgbqS5MspdIeW5g5sZAWfvSQnxU
kO27y60FSkm4JnQNKnsYN8FnE+f4hqKZ1TYmbVwY70PjZ+5O8murOsw+Zf9e
RgpiEiKFjr2MgtnC+eglVWJLx0EW3XNHlV6ah3rJePseFWq3wE/HyiaL/aM9
IdQwnzlMPQl974S2l8d1DM2nkuvlzELiSzhqe0CeYVwg1L7Z+/g7toIcfMIM
ZziDSAAd0XZPHeqZhPn0mfeUageUFPLqzNixk0dgk80UZaVZ5IXQN/wVH8oB
7QjBkqQoKC7WERKO3TztI1sjUoRSoWUHCj98+z0f7XsGtwLq5o+fWrGHGSRC
+OEGEpNavfFlwYda7qYFDNorVz9BrYbA0jPfO0teWYfkm5MpJtaT06GPu8Ti
sW6IWWZcA6se1oDpi6UFNUR9k3g7KhNtAA0U0TUm8jheaAH6SEEVTFmkK7A8
dnyOI/S7kP8zYovcEbUD+eDRvJHs1SPoAeEQX29UIgE+Ssn0ymiVyvldcfg1
ySLzORiXp/xrOpc2OrJ8Da5qEJrb0KLYfJNLFjII6H46cVyfoD2XjEm0wwVQ
Q55KnPnCw4RNNOgL7nO/DFQUApEehzda+AEYyv2ernLi3VHR9yBAIP4iNJ68
GVHwxK0YT6rV1ie73HDUymeHsxLn+e+5JY+qwFsWIpJFkF0vJgwffpTr9TOq
FgCRi+MbvkfRDBcr4g9ML+LNXnUIitAZuyvnj4vhdEfKP5P1EOg68tWIb+Vq
x/aTAxX1xKCNGBiK6ZkzakOK47PEjASZi6OfEjTlhXY8GD+rvxe93+tHC7Tb
mEHYatMS+Wd08apDgoL5djC37/sx0Z3H6bSOC5Fce2sm80xXQJB4fCYOzwKw
hzwSVuOVJTNV8gTNuM//ww2sRx7tnl6WvzQuC8CP34xlmsvGbD2DhhSHUwfG
IXcH2VcJFrAfBzeS4jn9D1t5IQhVZllRXCqBHm0vqlVg4MJu1+Dqel2XIKaA
iHaPAXzWH/4O5vKKFfMM8OZRieoNrBWCFUzNmwMFYdZ8Sm3oHRCE/AxW2x+G
NkA+yFJD3ucaOGsdvI4oEGVdJdwSe7OwVxMtiHH0KfTi2erF3Y7+pTAxyi//
nmEN9C7R1xiNcnZdXJjhAtxwGOUm2GQAsTAJs2QBG0AN4aibDQL2FpoyF7cW
Ol5bkN3ZbcbQufC2c4rvfjCXHwDxl6mwo/5ei+iSpGFUBkRCrcJ+wfnGQZK0
aTIH/s1Ncvh9NNpVBu1YmjJJSAux40aTwqACSQo6bnrZIJYBODDcNjuRbY0S
MXDvDQx5MCyXDxeG3k9HVYPmA3174dNMPe7JFUHywyiUGtpaA8f6cS0SDNpC
wZtzjxpMfHPEu8nZyMy7t9ScXuFnhuSLCyLEEEeS7jKaB/K5Eo5Trll0g2PG
XQRqn6nSqJ1Vi2+EIGVlQdXOHR1kBezuTVtJMSLK7qSezvbv1z8x7IiCtQcy
rb2pHfjAp46UcEBaLis7PSYFknk6gTXSjoZC7yJq1JMotlyheIcNiJ9wTs2H
vvqFYjKS3craPxt2nsfWrE9HON0bpyB8cIHQ6yAbFmJVBRnnJYTOElzcIMBg
iitEs/gxc4OSalltjudDkLLYPsmBdXvHe3r+B4Ta+7qaz51fA8gTkh9Fzw7B
LPmBbpBffLeeamhGoFCI+G9kTSZZrZA5mqZ67SbwGTgh4SLyKgI6nlX9OFJa
ZNn1Q38nKqFCJExWN6cuP+mF2Jhmn8VBWXgkWnqxzqCNn2TDU0uQdejeh9r2
pP14ZaZHILIXb2Tk5O7ystbIKRgGwVUqJxEcCTUAjgYQLx4xdkqJ71mCECvj
50eA41yRmTeIMQcW860LdtAPq+kYkc/xg5MCT3I1Wm20ukxXxWnnoqTOFeiV
vcGhoe4GtOdki3RIkh4iT9qAaqjy2Kz69y9oNDIKjGb8co2xs0MdUv7yxAPJ
vQVKWlpVWlakjdmrp+xPQf6TAWVj/IBuj+aWab775Chl/fq+H870XdoWMxbi
ugErSFLhtNsxJLFT2SfmUMHFqaLb5pBCU6U8D+FaX9DlS+vxBamtSXrBIAWG
TyL75BLLvB2IcMdBL57IXhPcBc5i85Q49TGWQhrgaPZGoZpRR6ZF4+LYjxPg
SPRXspTFSjvTUVOsCJynyC6p0pMPagBNVUmqb8kUuV20wuz0BEN7MgSDrUav
j6/Xsk25dock51+pGV6a90OlSQZDKaxqc2q9rVbS4aXP8q6eHSV7G3QydCJh
6ejuB4TF6XeTCZTwmsPo1APn8Fl4Xux16FCQ+bcY7tJo+PBK7FOXSUE3zZvn
y76Ag72z8J3kLUWdkicPHpg8SuGSo0m/6yFGWvwRWh7v5OSjcZBdhRKrx7aJ
so0WNTmzqoxjeB0Fwx1O9fGififVNqESJKJbdgtQKzLIZH32qLoYsFDPI2bx
kE+SC8ie+iZVrCBW3/JuChrR6+BiOZmSOSPjBax8SpXcGFH7PWqADdXt8W4g
eSLv3e5d0dj+yyjsSWGDzd8r76yKDNg05liLXzWSZ9xUaBeNWE7oKtUxj1gm
V0hbleN9luh7qHa0g8lu09a7rNsYKUoPYoQxNbHSMFxWABnAhTiVci//GLFT
ou2CLqKQ2rkQ+0mAG+jFYcEHNRo9DSva4Z9OnknPocG5GZOoUxsa/0R6LULW
DPp1vfW+UkER2qHFbbm749gvJykIefbhz/YpUhRqus7V5/k6651OXLr51SKi
aYIXLloQ8BmMGrkB89dyNjPuUY8IuTzgVNcwtRCJ+GK1OAl8PdUyYEQqMATo
oA6Eyor4nCmCyaZg/vvNdQFDAExbh6IlC1hzUvfPMz7TA1P9SS0Xp8W/iqtS
Nw6JdsO/WO3Z7lRIwEe0Qlw84ppQthQ/TNjTYErVyyecUPctRz3E6H8Fr2X0
HLtGeis6dXLxKaN+z3QiTdGux67bMXF8Bpcs1QIL8sOTnEvOktdOSpVT2/Q7
LJeFLFJsh22IqCREF08Y9RINLp+xKoA1vZtgXhZlTvVrbluRrLDrxtSWxZnT
Q1xsMHPQSgjr2nGD2H3Kn6+FnAeVKgtP10gkeKn15HKoyNCwK4smJtigURQ9
6Bim0IC6fiRr3N+XY/7LDLGbQ97FFI7yjOxPyv9cCxLgHxhrSRfDDi92l89T
1zxazdDsygX7Zp4+JOlLcpO7H+ATOre0kzwJJcGcdNq/BE/qz01zj59WZOVF
YsZrBpmLcZstxz+hb5dpz49Dcj7kE6zS/QdhpYMeSqIvstkY2cl0RUS9mi95
xXpJBW6XYH7DX6s/NjROSmDgvgAbT0NYR05xX6ZnWnuNi8mfz/acaIuAhKj3
S/X4Pb2lUS0TulohyemmnwSz0U1Px7S5kvj71Gnwl83K2ucmTtvLk9SU97XR
YWUsxmmbbLYvAPIq3E2y7d9TADPvCMoUWY2d/0Hc9usM9swI2hkUajenGO34
7oWalzPB1cNNFQspJUuF62YaSe+X2GJihvg4o8dz3lvHI2SCgyYNSGcZX8c0
3pbG9eh9Pa/zpmERrTnpoIfwjkjIxYLK085f1ml81CjfGrsM0ZY6dIvtPufl
SD1uDqhXVgEJBMTcf16b4J6K0NuXflIEjYBd9tWQa6N3sYK5yrMQy+ux8qbo
+Ws4+kvsqIX+tEgyV7f/NjCtx323Oi3xxKkmJuZftO1RpiR6DTkTN1RWYw3L
weYWeBflLGkQwzkDO8UsFc4v9km+tAsJbn4/gLFb51Cvg354AKsbCxH/rFKa
V/PuudJGm0Jl/XJPsFHbtmXKSg4/v1NC9nvupJcLbmO15PX8sWn3goisqvF4
QSR26O8OdrLFLxc1rj87uI1M/LN/sLjD/b7jFODdt/BN9oUiCDvJktKliSQf
pQBObsekGIjWS1k+uDuWeM3GxOZ5viRegk44cmQpizhl1iLr1XkiJiTqVJim
+jceH15dIgv5QheVvMQ9v0G28p1craW1lkfWDLCumBkQIKL//1v/SinA+UR9
/wel+Vsmx6nOHmPZuW8qjZmwc4fSq36Jwn0J+/kQlJxCw43217JbM1dmg6xZ
/7cKTomhpYnKmMvjRXXHNcMXa1DiFVRB+xZ+lo3KO1L40xGbC4HanJvQhdcp
gbPepnSjwW2kMRVPXL6lvKPWIO6BRyRiDEVekRXEDGEUfCbfYtjqT30KB/rj
zDpjXO3Tq4Gr2Tm4g4yvNGii2kv+hXicxhVjijyKxx8x4UWC5+ouE14Vpj4D
MTrFWCv2cSO3x7/9kTULJOeG2BfIvVFONPy1I6CiprfD1UvzL6qPvmtZ+O3f
0qDgeDLvd2RAVX56srANdjQSgf4ghvzVTCgMEQRqpes2yCGJxjDh3ZKz+EJL
mtWcdeXb9syfhPRc3cwRLJ+Nje8AUIfXIeDpPetoQCwvJfJt2ADuYDenjzzT
Lo8pi8myHSEeuvwzVWGP7GCwbAWo3/wuUOh10EoeInGqTM5n6Ul+ejbj3b0a
3x/NydpX6eV9bJTtey7Guw3LhAVmlRnj9lYUEBOhZcsE6JJQtIgzUAELUn86
MFbgkRiflfHzPwayAzSUu9m2raBpcb7OJsbuPKCCnf30+H6rSbWXCllCAwAT
PXbH6exs9SF7sf341LoiP2Sp5AOoDyCTfTzm9IuEtZf0CUA/cg0k6aG0vd8w
KnhxkQfZAH97Eld3n51RGXJgR54JfT9xRoL34hiTDtqNthSUI2hFVRKPcgF6
paQeG1ktX1dVvruh0eFBHxlbJsP9Sg/3agxh3aP7X6bKC0wlM6rlW2mvzPYb
4RCjDxYDzq5HzZNcu/M7FhrMZjpCU3Kb4AzkibaOxLyYj8Sr1n0TrDI72T2a
az1tmEh5PdmD3iowbNGSHmn7gX1q2M/yJggvIH2on6CB2WkRy3dLstRXX8VB
7nv1K54JkxFlFgmkEh9RfI6aAqjR7e1b33D1oRDuwT5r7KwTBBPxfljjVZBs
UmLlXGRxlKfUCP4EnAydl7mrnAbsnLqleQ24THx+Be/9SRaq7mK92JVA4XcK
sqzOeJTrQWGV+urVvEpNIUMryTrZLnG8W756yZn04owiPDCRWregJHDzFMCX
F6+sFa1KLrj7vHv/PZ2rBynfpz/ypHXvTusT1ZKJ2z8s6DOqMGynYrJgm3xR
WlbSDl6dL4oN+md1c77GgvtDVhrTwM9Ui0lo6jG70mtf1mAK85YqIvoerlfa
LnDodaEoaRtOnfLd2qcZEkEv2H6HuQUGcoM4cV/j3eJTWwVhI1ahusbS2HWQ
aQ/KP4g5OKaW/C2KX5f6MsyrOVuO2uq7QPAZzb9qZSY2usC+dWrKahQAVhse
e9MRLWh1hWOw+jVFW6Q4QBy9F7pyv6LioqOAGujaeGMJzQI5fQehEzD3Jpnc
x2bDLhCa9KJA8N1dmR09UB9UTeJ0xVlYZlp778RPx9JKQjkFhp4KirbInsGb
OmFaJGlIubAhrWW+hiTo8Twh3tvNiMfRojwfploMMmgGWCzEgU4XhO04mfPJ
u3MTUCXk57u+vT9jEG9lbmqd3KDUt7bgXthjaJxgGCyMTVh8ht9JdTOcEcx2
yPJkZ/zAxkmxNwbQ6SdkNUChzTr6FTJc9WM1akO1xVl9DzkN88eKo3+Ac2lp
neB1g+JB1xm5hyQX8YGtxVUrayYAxc3UbfIvykODxasReyVMYK5FRSnkwabN
YglsGUmTnYJ4/tuQ+qCucFvXfgS0VKP72mN8yA5vU8w6Z4GjOt5ImRCI0lVo
cTqLRecVQ5v2SmgdYoO8nFWJKlLE+72mWJg6uoaJASP58skkABPq/fub3GWS
uQb8tN9b8y1OLj3s82ufbMurWWmPWuikp3Dy2XewMVhp4TQ8zsf57uZFFjfD
w/tV0T+yKvJaI7Tk+wn1eIpm7JAUMLN5HksmUhgMVRq56oGrG9rTOvAVv2/p
UBxmjjA/WLVms4JP0wUB+G7cmuBMH9a9Cw6caHxFmDd38daKxkPYH1Qq9JvX
kD/crUZdsHSJRaJzLfakDD0lEmbU1ouvB7EKnXZFwBalQ+T7u8wY0eVneHUI
PO3xER7jXI0hfu5XBRG6SnJapZr9fhdArFU7KrczcGjTg3pVU4Ofb+ZrpcXe
sOuVTPeiezXWauSvfSDYzSRQKsclVw4/wYZqAAPpQTEUL1ZSKE8mo2cS/A9x
Kdr1X4LZ7mQyCpF16Q4uNpxFympfcFGjpZ54eXUqfgkBvWKWQ53MtS0pWWMC
ZHl2VjxLnWxwwEEJ+IAW5NiBv3J/eEC3DKWCAUIVDyOcOx5/IaXU4SZ6J6/p
MO9G3EIR04l5r1AdVymlIVPy0oLQtL0uyhoe2lhNcZKDaK4LFXXcv8DYlOs7
O0VnUZ6LoVp/GC/qHsWSSfsvtLF8hz1547CVw6VrgamBkhdfX439QNWkrKCb
Nsh0GVbcasbnmNbqFkifH2jQK0Xq5Qn7paH5bwAv5p7XnKTXN/Q58A38FXLK
J0D1YIVnmRRC2ghC8WRL2snhFJsTIxcYpdw5aDdwLTIJiB+TVAaSiKR5cFE0
CLrOGXBWHE5Loq+A8JPrkYIF4X6eCbJiWSyIRvfBfThIXacQMvp1xZMXnISL
+n0YZnUn1I5H1UKyzdLmMe4gCzMlNu35rd/w61mCqG9l1rxG8ekcb4EB3Wap
WTYE66iR9hKqGWWYkvDDqtIRufUa/7UKmZzjbU8B/FLtiNe0kILvGycqVwS7
A1YEjPf4y87ojSQzwSRsfu9dwne+ur3VEUBEKoWmIGTz8oEaWJmXPNVJ8XtS
/kvWt58wH8YQMAMTGKy52gxIX+3qPRpneAHhqZy9+8BjzESG3rgY7EpSxsAh
dKFrTOn8xSuId7eg+4GPz6+K8PNgpUJxf5Ysk2mHvGfEY5L/W7T/O9WFoMyb
GKvXNqKBrvDgjA8UQ7HrxWfBQxYgxu+hk3fJomBV+sYw9SopK/rrjAFuuleI
jJixT1Fn3GqUG7TZRmXP5ZsD0KLnBpfKL3cttGcBFdTNuFYNFv3TLJJnZ/fc
XVM318/oSC2ZHOt3BcbYI0To3YlOJ4wb3rZ58NGdw+0bkil7JvUFZ94PrCcK
m7jso1FNldzGeRm2SL1yHu0HhzRaaOIKJgzw062fl80jibbrsL68LNgZZdaG
TkpAx6WcZmqiYG5IV5KZDRHofvyTUNHq1khiX2p/Mt102E5gEOo2ij5583ov
OJBD62hyGfTPXZIMNQBCw62R70lXYh7B+Qrw0PQuv4gHarRiackPfmpmeGxu
8YTagg3+Tg6Jl0BvAx/MAQTrg0BOYJmaFLqzRDQyPy+hllD4fw5W5gJoQwDQ
zaoP0kayDHSUEx+oTqEBTMXMWZ9chaL3wWqu6yF/en//gDkPpgfnafA8I8Ab
pxMkwtnkrSDNvNSnNpLG+aCPEtKMZlrz4Bk5dPqOoEx3glFq+wdF8jhNo4Z4
3HMyFxcH/4LHAY28PfvLWWXQGYIQKYsT22rCrtG0BX0x4WMa4dpIpOQSR813
9Nzead5SAL0sVLgSVkw5csqHdjuJD9S2P4Lkmf37p7dFSbJAOURG5LYPzsmW
MRAMCGuhbV034BoD23bTJCkfbax6iI8a1UQTqTZU2jYDY4ngDDdo64bQByiZ
J2jQoJru01Hld95w1//vRBkJP3pqz9BRBEZT4ozCQokHS8Pkr6RDJJd1Kta1
tqS88Qd3+XkZ5bYPJACDdu20wf1Xvk4gUUZIijrPuMbkjZpm0YM92TrM465s
c//hrCp8iFL/RLYoo2MY3tvP93B2JSYas3arCaMqdrFnq1taz5QjrWx7alfm
KgaKRU9C625VBa6lQuug08P5yhoVWcq1PDE+teaO55shnUXiVY0Ivh/IqEq4
Q/mRS4OeGyShoCxr3QK1vFotq5IEX5Jd+u4br9ufaNHWv9ZBLshOxpO6JUnL
9O8vnA2E0h78FGEzL5hKjL6JJdgdb9sw6aeIY1vK+6jB4V47stYxJWNHGMvb
i5QeKUy13DNDdmaV72as5oDIvsl75yx40clt8UirE3umyMJCqVP+PRSc+aHt
OaNXhP7m56Ef2Y3zhF1XFL044p8zamVobQbv1uDAh2A5ahfa/rLIyRWPN9vQ
W/mSk1MOItq9ULZ+BqcFXcs0GuC69wMS/SXzSdsipyCh5HX56SU/v0bgINGK
WwhFFaGcIbyPUHXINmnHmMxcV54forky7tNfoadXFjA/Nzhh4mEYMSn5DhmC
nZnKSZVnyUzRtTHE0avhdI0uJPUYwRingxK3wgKc5OgPZe9cYhAj4AZZq6yK
uMQRw3XX8tbTa6uTCLjiX0OB6vvHmamxvBTAxNBqKPEnwzlpEARVltcNYMd0
hbZUiMhd53J7ugbndhW6Iky4epNOrdZqrmREh6rgE81OlhUfpKg7h+USsjfh
IRG6X38nhhAJUb2KL0Ft+y1O2ZcydhxR9YHoosFlMwkstiBgb9LaR+2P6WKe
Qj6q3XWTJ5ubdBxSgymVvu4z0OWIvyMRcA5jklyZms0oLpKBpiFe1RsdE+HD
cKeJKEBXmm5arhgClH5RGRmi9F6FIBQpqTmLwIBveCIKCEyinDudIC0Gyn9T
UxdzkInp9aT20JDq7bfA74eWz5e9pW+vPQvWIkDTCtimK/yNDdrXPwUa/yYy
4HRL082RcH/L6XIjaz0Zr8nC5tP10btGdpVgyJQjGY/Ssbj3TbZGy/RGuaal
l8ckIEOMvXAdRiRUKvDp3slFXEsYKCFmeNjYkFKkzTFPkdkD7uNhjMQp6uPC
PMthuRrY/mMtNdVps8hzu1dV8IvQi4l4JtPhDalZ+37AND/A66Z+X3pEDXiw
zORPz0cgFR2jT388JtTWwBPWCPsAOVlqNvHYZ6XmSBKEnAnpg6XLTvEa458g
ydg+6feNdwHDVQdwpKE6EgtOB37wEbXtiQ+MaCxZSPzfJLvaWdB3DNozwGl6
+dZaNVeyVY2nkoUGyRjit3vpKp3oEHNfBW5gyG+WVB/8GfIYQfigKyXuVFT+
U4v77TpNMwu+vtgEJEWNwuwEFLOh4JDQS3Db0LfZpQyAvQZaDGkkjm9oNmGY
2qcPWGZXmN2pGtd1GWHoc+YXNdl4wu78yUdYPQbEpUC4ajVc1Ix2BP81WKHG
m/3KXlyOKAEQXdjdzhO9uRXtWNooom6ZaZTEZ9o/YzQXYRE11FN7iUoDgvyl
EJ3JZB8VyiE9l7Wfel727GrWufP5Hroel/2doHogC3Dg7z11lZSaDCwrLKKO
wkNBdaFKhoUThPVVFrMRDjEdyFCTF5zSQFASRzu9sL/XOA6dL7rIh201h1YR
gbHxDnS4ml4yj0fnav5h/QSOWqpuALx3tg2bCMgpg1TLj3spowD6hkJqSwdu
fgYgPt5FWqiZuqnecfSAu/TI3uGMKs1Oge37/kxpnvPVFsIgyKldaAaqPKoQ
PLV4bd//0Ee/lyVcA8S4Ck+J1fjNRKx6wlWwcxaM77KezrsJdPawlzrZftoD
CcB5o6IsVoCm44h214V31jQFncQ3Q6D4EvBikw1xMxpLAQF1fVoCloCXsaD/
4lBPQzHJr8cqIhEOa4bDLzaDKcqUw7/TCsecMHFT82Cz3+3azBlnwphfSoHI
4kP90gzmWfwGDmP7dADJlY556EFwiFylK42h0bdxTO2s0cGeytFvKPQ9Ews3
sHzz2XiJZwjnwEYKhKGyTNOeIcWexcQO+SY6d506wuCL6FNyNUZU2ZH2Swtx
uZr9OJ2KCn/ilp6m3cASUh0zn0R0PXAeVNKubixY21Pf4rEDJO3J8t67IV2k
4EsXNRzY7/T6PyTf/AorHhSH2YXhe9Q3T2Z03c+r1pwFLWPv0HW8vVxQwIf5
YJlGPYRAGXJdOlGkh0tMfw2Otyu6slv1JTHnI2QR6lNiAR/HSY6lbnRydM7y
16fZjQaCHY4+TdTMJyjowFvjlJfIfRy5dzJky3FzSKFXLLRfhX2rZRmNKjLQ
Rf7hBNjbyMj38GQx6vzuviGgYNTE5g8wGjYnm7bVvKjZjCGrwxjG22PYnD8g
YFumWOR4aAnceaQf4J5gW9ICni5w9SQw3Wer71ZoFbf4aHwuCGHjoCxbUX7g
4QZAfd5fSRxfzcNLpmow0FLi+lAuQss0SM2dNx1X2X4Nm0gOKu9WiNmNVzuj
JYPkm0DxSa++xpQKwB+awZ33IT6hmwuwjILAmRrm585QJQstSuXTITwZi7YW
w6hrTVIq3O0lhPKXNuO/5cFu5aj1Nbx7fpw8CcHo8T/MkrBv0CddVsEJ8py+
BKGJY4/ei3Wi2zPEmlQo7fbEIvmEK3C49VBgMvcjkX0Q3cXvIb/OYcWhSzKK
C6A/TsDWY6rH80ZcjnBdkXaZLAHt2DXDXpIS++MY9Ql5dU1XMGB6m4qVQbh2
6d7lEm1j6nq7CF1rfL90l4DFhHMx5VJip7yHu9PQMTY8XX5+CtyP+4fDumx/
KfEeXSMBIvUo4ABrKQ+xoT7zmRNsjqysklCoqpTlcRl3nvdLd1E1l3l8IJTh
5hFfUmQBEDR0RlaxZd/gmBgxwfcGjiEwqeElsVazYIBqpw/IrpTP9B2XTXki
EpDnLz8+SuuQeTX8LZdCDljGLnoZqizo6URKCxcxcO7dMimxGJ632dGjO2KP
BgEEHvMyQo0P894c3hZ+quRsCaFQ6xVnLP/kBkNZ36CeQDhhqM+bTGkIKtx7
0hkEqqDSo8oMC1ufr4vgGP+ChOoUuDr/zZFNNL5O7suyeTbrbBppA9fTNcQG
pIJEWpNEk+SxMUPFvsV3FRB48B5+/EojqwRSYU1a5KG6iLyRDIlXipK1ELaL
RpGIKOVZs+UPJEdWU9JRzS0Zc5qBqUyKXLGO2u1bqOyEeFpqWIsGUKk1rzFn
w/UlPktUXCBmBhOWG4YWsDzf0xv48dcNeHMm5ed4U7uTEL9KuqOuzqwt4jz3
4OFAs38zF8X8TI7xeRq5gAiWz5ucHkKrOzHKZU5tpTBQejY8SVGKrQwojylw
HwdVxZaahGGMsUQpfMIOIUQpjFvHGT5ZN4MgZZhs0wC1GLbB1Ab5zlmiyz1r
t7Lq3zUtKs1urAOtDee1H6Oa4TEjYzGGAa9apamWLw7AzZ0QtIRawpXAjNLj
zG1RJ61vW2rWvDwXmnwBHXeXUyPUCWiCgN4nPgGVKEU9Y6okuwtI2v7HA/uR
QzGNAnkDGLoU4dc0GTwHtv2jtM72xvMBnasNm3k5UJ6kDGEKr+j+qSrkcKBA
KXnZsK7Uklu9dXEGNTL5/nLe6wyaNa+27uFNzKbTlzc4ftY52vVLLevt8K37
IGQvovw/Z7/zlPQoXTY7NEL0oZjz4qWGKkeMzOcLeNHwgd0k29Q9JFf+f6yn
XWorvyALM43Y0Z5bfFZ1hWWBoUstmZmLkecfqdfJlR8557ecFpelrlr+bUxT
SUSA89VaV1Ity2ZqknKM6BcdsM3oVij+pp+Ce+x+ztBK/Tg8T7+XAhNrx2ir
I7JlKk4tpXM0WmespB9L1fGNSDzanb+lKBv8eqFr1zsvB7Uye7EJFP0+diZL
4QOF0aRgwkYdGg4qiuelRGYc1i9CyzoyG+jtqqICk+nSEE8GRupNjSVz5XR1
guTFo12Ia8rKXz0a/gJrdRbFxK/ldyXGea/h08hUb0PIqUD+SosycWIJFDJF
MSsCazSmD/T/IrIX9g7sG5VRmZ4LEj63gGheO0L0A4pbR0Sb7uHVs2Zb9f0b
YjEKflp6psYcf7kl7WCloJjxk24SXgdKVaGk7lWzbiIHOiZ/rcWuvqgjAyyT
TTMqxCgJoPJFwkZtXcb0JsirL8R0WOZ31GofJGwj0p+h0PgZ/qROlWFnW/wr
Vco1otttzVFwioOLf8Sb9S9uz/V6jbvCva56XFBicToB/ZfW/RxMX1iiB4fv
cPurEGKHyqlu40N8pzedKiCm2mIMfOPWIj7guwlDgjk1LMa3/l22nzM200UE
CHkaODYlhoN8Olm4jDle/iwatNWalF8W5QTzmvx9qK8Ub6Vq7RnuoaOyY9W0
F7aJ/dm3fl4ynMmRs6qklddzLCFgcRYmbeI82cKST5hU+UjcDApQq6kJc1TM
y5I1d5fvTnBDREsCPCxMT4ZmYlK49yRtSCtHkYNoxeNKl8b5P1fv4a+++I0C
Y8CjK9C/vtLS9veqWIdnaOYP09fULG3GgGEfst758Lz53ayXE9MKdPmJzO8d
t3bUW+6HnY5SW0hMqoCeWZLhPafvqjg3RMMNomSKCJvjW7+GkAsKBrYOXt0N
OEQMn2lLYCRcWJg0sjD1rpkVHdhbQ5SJyieNEcYSV3ok4cHSZuxf95iMn9IQ
+ZjUBzHVA4Ph/H5O/hu1/zGerYZ5CrqvfqpZcEqNXpEI0ErumPCgjtNNaRLS
g49iwH7zpFXKZwcsbOhHjxhw6txMSUNqwAyA0AZTDrxEZWpDdLHhhlat/wnb
dOg9m5JRR676i3635Tsmo3XCFGVZxBKUzcqIEYhqBPTefnzbX78+PLI70DuY
JhfxKAPUPuY8cS2vYg8l6GfUdviobC1o3k2LKxPX2j5zfJEu6rOBh7kahFOO
H7d9Xwcjj4m+jfFRuHXoLSJ/trgiC+8vJJDUKqeFWijL6LM5FygkI9BFgJSz
BjpvAhdk0Fwj5IXJ4nQFR0d/WBeCYTdL3uwLJ16AEzFft24dHwqjOjLWIaiy
DKeiQkJubnxIeyHe/+naE0Yui0wi4dlCvUm1/TJssZ/JDIqwZAIWWC6jZm/I
Acn/lFTzSv5Uya5IhcRv4uc/kRacKaigjipJJGlXv2MVkUydEc3qzbg9QvC2
ByFegTeEhh4Rg0OzdPVaUnlvsEuSOJDz4ljpqNXxDaAcfYAb1wpYt5qEqEAe
F+FpeIbPGY7zYtGCDziYzj1CXrU00By57zUlhOU9h+HTDs6oTMYAX8+nbeM6
NT9gMdStV/QazAFO6tMeG/N9+ERNjuUT6atcq1sHS4q5pFeRGEKli/X5Ik7T
d/xEJBeebDuv5PVQ8NE/jZrN7KhETERSysFZxYPHZut0J8f1m95BCnPDzLDB
BUPijkm1jOJWPS4hYedEZi0Muk52J5/J6eRwjmwCg0gk+vBzvVDVOdWoB0mC
QEWUUA4TdUZQQdTStfJOjK0dDSVuantwhmh+5xNLOYuC9Y9/aGPNeQPIPAoe
qNEfLHhpBqKvvcFRqwl7ORL8u33ygJ6fQCe79IsGAC2u6ZnbeZPY6lke4UgX
Lg8LiGbh9SFCccV4XrVSUPhwyotBn2DlA+cHt4u0p95PKQMdzdjlPqAikp9L
CRoh5SgtkS2LHBsjt7faqj0RsUNwYqyB9xHfqwyWkHIzhvd1US+xAVv2HJu/
fml5RSAHvui1UD/esdKahjWxj+D9j3ByhToAjRw4K6S5izcoJZNNY/Cyrn50
nhcNSC5gGOl729nr0CEr2ztrUfgrjMoAfDi+kbw3DIXMmJNLbm3Z20NMZxl9
uAwOiO9N8jii2r1lMJjCmAe82RJaxLvHmSx3gDXNKdQyuNPFXanDTIegNfUN
R+hiVad4tQYtjT6t2UreClpn6h/IWpdYd9CKRLeqnOXH19SuT6pk1I4p7vAB
KFd+J70P4twYDdh0KWzSaOtKnpZFLePh9paqSGhucw+4iucwsWJ/WaiFucBk
MxAljg0eR45NiBOvKsDVOKQww3O7HMpnm2Spx5kpHv2vXxTtKlIE4wDv47le
TP6rPnTKDW7shqy+42C93c2GsHO9IxGixH1T5e/Oi4oPWoINVK3CrCoK1jqe
jqxCScX+Vtlam0Rahm7iudTiYBuPBMP0XFGtKgci3Z+zTJrGKKhuibg4x348
nt24XIeE0pLGk2UaM2Pe2Mo/iJujMHZPAZTRbyngVm3IkNC3Wv0dL4pUUGjE
cRg/VFLZTiOeTBDzxZGfEaMdFFlXmwn0vSrXTvJ+LwnEQ9PUb2g2UYb7kiJ+
5wWA4hSF/8lMz0B5r9FP19lArracgWEXr8g2x+l07cIVqXwsgEHJIstPIhTI
X8h3UkBb2deXVWXELhMc7oNkzqWX2B/O1zaf7mU4YGYQB2O2UfNjnsHKn80H
pkofE3JmbdlSgAcxB78uZ4Nk6kFKODy1OWtR+IiOD/+5a9uRqZhy8bKzLYQl
vKETmm3aBVmq2/JbsH2PM4uYeGDOoAqSInWEXp5WkZQP++hl2xVtFiNsiqwV
vTQVARCR62URq+BwUl1wFpG+cIGZHKV7rfqUKYy68mekEcDHQhIA+eeJDdB2
/v95R//B1r7hhlJBdRsQzQ0XRK8kMrtNYR8LjJtnGs14EyMmiod5zWwE0vYe
xOn+X6vJTmBGT7mlSLGLMiZdsQfbvmpgffAuoICxdBKD+PKc1azIfPfjzX+G
1DBa1v6K53v2T9rtXMHKGWcF9dSzWsM9uK/k32Ipy1mubBPFw7AyE5OhdTvc
Kcnm/3X+jOsY6TyFaYIiTRRVWEXVpQXxkt7hosoc8N5zZYWH+07fCX3gDP9A
lvvf3fGrKP8LW76rOfUn2RJ72qNGhNLPCQ3b2S7WXkrcpZ516ykR61FrGgyw
QGPCwtMpw7/UodHmm6LlfvLwHjqqnG8Yoz0XSRlSG2OrEChmuo/svsRlX/Gj
VWS7vs7fvqGt/ux1Spbfkq94f1IELiIxaK80FPKfzyXEVZFeDfxoCHnRM9r1
AUe3kJ/0xq/Bifv1QqaZQBI1Bkaukd9weQhjQgaVbKewuRi0biBYLxDMy8bi
12kh6b3+aPjpU29znhJ6RxtevEdSSpMFAV61tQK060zy+z9837kZ+OETSIwq
aOWqa8LPau1uqmCIVXF2oOnRnUNjY+0CxTTBSoaQE4b0f/y0FNRa3HY+pWa2
md27C0GDyZtTmYQRDwVgN7I38ocbnA8pYRbiMlqBgqPUPKBoR9KDV3gPQgIX
nPgxAgkqCQBszEZg6Re2F9hD2dX8j1Ymqnsa3Kc64z98Hm/2zKaG6ZxFhTh6
GDY6YA1gvfEOjPwPcUIo8RqtcoJCo8VAoo3rK9PLqidc1jI58kD2ZC1PzKQ7
ITYICWkV7exDHsyHdZByA2kT8A7x6acWPFuhUaozzI6AsBzpI8+ACVDIqqTw
m+LmUyDt6aVfJ5V087VDxPVYbFvcoQFIfql6UqAW6i4Cg7AgF33ZvmMzw3al
Lnr7+ThPZnX03J72jMQXvgcl7LRNxJf043f8tsLnkKF9TYusuNIa07DafGsz
xLoGYKo8FTvkXIn0NoKOYF6FkOKEblhkNVEZu9oflvEtTxZM0zQAqXGbZwwq
4NBGvePasCK5X5KJFIVRp1D4C2wBetzNXOjpLKrx9NpPvZHKqzM+uA0PCj2j
txpbCIicdatxLQzn+jMWztWZZFZsLysgg1VoSZpG48lK4BSxO9TCLwGvHvsg
yY/0YfJw4DBkyi6K1qw/ZHPw4sZQmwLdRLrOBWL5fOzvcS+rqxO8x57HlutB
rm4yA0DCuTAnpIBtzRw2HIz7bVvPJGN5ZO62jDOGpFzzG7CRa7lvY2wr78Wi
A1xRv3q7N3UrYEUfz0S+5pHfFjfjjFuxqRR1scBb6Pmhky1NcfDONuBkLFHq
2fDtKgHxE3veMkw79CQ/f8R15VAI4jzFZpzdP9kickDNSk8um9Jz6+7rJT4/
vdenu702qYzmWDqcHozL6RwbRC1pO37jA6FGs5rl4dqhqx4ViZvpQ8CQpcDH
lTM8RFR03LswpjyCymW2jt44xEUBWc9BczGFMPkbWUlZXL3gpl19MiDPk3NH
f2jG5bPDHxHSS/XPG/31SPiY5tQM80dIOkgIOjBuM4mkZWqlFBEhA4GGhK9z
Dm0ZvHEPIJcqA9Zmxkk0QVQDdVp8Kyl/MYnuMrdJrXkEUbFKgxaASfZBzkFE
MB2wkdYOT1UqGyxLexmnzfWkRcUI+CuXvG6lFxKgPte8OFb0dNoKbwQ9XZ6u
SrINBVftiBnfn89hV9QRBryO6SrdcV1PUm3sRHJsGZWvmeQg6PrjF5zuaZhr
BXdDo5+mQBHDozVDwUHtKfyshVKhm0rrfBh3l3V/pxkLHU8UtDvgww8NUcFf
Sdsa5E/11NL4VZOdNu/tfy9DkACIeNnuL6LStcSiNzudQSmD4Ue+yfKaB6LR
fT1kdT8BhvpLfQdThsVJW4pHl4B4qqdzklcDek4cmuqsj+kLKTK6X9eBNF1A
R54YA0bVZCun5bN4C/DX1EYDeoRaeHEgy4v0gEnX4WhFbzO2AYslvRnDOAXy
bvSCUBmjrtKLpbOHonM8oE++usnivoBigLmLOvuuQ1cbT3yJ88M+7KGTXg7d
ZvkokrbXwM0MsHYhF2/p4OpnygPSKerPNfDCoHb/wqB/+y3vcNkgDhkg3cpt
WSjVuAuRdLzXWkwQOPLmPgPUCLQcWfyddAt9uZMfRRWgIccCJvipytg58r6e
zeSJiYxQgQ1Qe3FfaiICCI53sizLjt5PRufH3RvULJlUmkgCIpqjufeevyGc
AthZ8jiiokcdeOIfAGnOpz5dBcrlLEUt9QGKDXyCCu/OLFpt3Wz42LSIWSSm
PdWAXhL4oaojhWijlwY3TKZBikvwIbuEuw7kbdUrDvVcGOnUub5ITGirKxFz
Hek2rC1LKKO6QPA/XON9gwaad3v7jfREw1U+6ZfoBgEdkf2k5oMXPkFKPuVF
9ZUmS4E0FKWpERVxDUWcOVxp/E1Fe5f2C9WPtScsRUt2nn1q4Bvn03iBMujy
8Ceg1Ed+qQ/SPcN/gbkojy5sN76rxhX5YZNVlkY1VbJXJwNb8ihdTLKxRu0U
8uE161XPYByhTShvZ+t8MNm3qguhDXHKcITQj0dxZk7bMkn4vFbkP1P0ptxQ
ibNTmQrOqVB1ZAF6QsVKy5F1H7zHWsgL8K9nCJhRnMTX5PUnXlcjITN+Ssoo
Dnw1d+4L8bFhRWUy5C7AztrGnZgE6PbnNU/lKAQaPSibkdGkX6sUzjZEKM3N
u7vrO287EpSFd4MvQYy3cjMYu3wZJYDO0fETamdv7NJHjp/fJpYWrFZaUsR9
NCOpUgqOQTW1lEIsdkn4XU7hWTqQuqqpd6NH4t3s8RHdVHz7lpcH6GH9IaYj
BwoKQ3VvHFN0G8Qk/NiaEPMCKSQey6CcEEiOrZjRFh8ykjbUq3VgLMHZLVYV
+tXf54YzkNPImGn1kaGxHsb0X0GKl9FXAzsX7+/OkAqcktXKBeA9KTGVp6j2
5BGOukINgcrIqfL2sH40Mjvx9q5z7kr6fv0S8BUgv6TDOumRi7a+ZKcMqXc7
JBUN0S+4207s3fIMdJ0+r+Lc9w5JCGEhXS0Agbp9C9XBHL7guub45h9K/g4Z
ufH4xELKF1HYMBXw5XRC9wzwt95CKiK1Dgtw/rr3SIkRlGV/4VPiYAZpJYlR
5CZ0v7cgR4w/CMPG6cXbBfqtBMYu0rgz1MHPL9GtypSwx3BxfnZ3XQm895pt
cVaB5m3L4+vmHZ5OoMtU3dRCAI3ZWXEp6aE+Jur52nfOFA438uOhKZlteT6u
sqEvoSn2VbLdChyr2hfvJkKSNm2+PhfgHI6LvqmqmBvaMK++5vt1Ts4Sz9ek
xK5IHVkjUTF/8uljzf7yX1UZRK19dkWcWfCU6MT/vJO/qk1uNzDFs7//D3bQ
1Nnp2Cwr9JQFpD1zwdb8d++hqCHuQtldUmLz9NhaEIaBnlGXrltgmZE2Gpqq
JG+JCK/u8x+dudM41QmMefFugenbnfYX36m0+l61Y5IUGFm3PpWYTQ2s+e+n
x3Ef8YAdXWC0kGK3LB9pRUE0lo9UnD51fHgiPqynB1oTeX+pV/8nNLLI/1qt
lgiBYBos8JzzpjgosN7mjVsM4q7NvhP5V7nxwG4XMvzvkQFO1wPkYrNXGPEH
qCvMcHuNO4Cixj8f9S0rDHDRYl4hS9Mpk5O4DfLRvxg/rhxC8gy3WDT6yXM0
Rz4jyEysC+Ws4udA2fA8vEfZajOLbC0mIoozRRgABBd1OYDvMcxlJ91ry4Q0
rvw94MHiuXyveeMd6KFBNENGyROPkfYiTMDGxBqqI547yIDraOJK8agfoZ/z
TLTv62N5ZLy/XtYeXiH8fu5DJzel86wBuiTmFMbTxybUdDNoQBmN7r0zvkaK
b36qILX2jeSg/l0bXqJv+PpaK1W0M8TA006w/2CvaAUG+q1QPSGPdYq3BZsF
9lqgc7oPmCoeZWVboH6yt8Ic9pknVclCtB8H+NcgAmoFsH6+tL+vs4Oko0pO
+dISDj3eNAv8bUSAiDnrZp7nnJJD4yGm3EzUXxhFsMh2qPHeAoCUJHpZBNze
lthRQsaQPuAyl+d0w5VEJdW7Qn7rmd+WbbZtI1hyf83J/GzqijD8MnafV+zv
6VgGb4plH+nYgTs+ZCjjnbPTso6JICRm3qhjvxVBQHqaLeDYI+W8yPS6d6HZ
4xkO7mlRosTYJx+rZstGePFM2U5Uf9caAvH505y8g8/DM995Tb10+eRtxdJw
mJ9YRrimAS80qct5n3KOo0zsdemDP9LgpIEwaSbG1WgnV4P42wzuxXHwMgCC
7Fo87G/XJ5mtvEVj0kF8V3K7Zyv/n+Ig4HrUi+11tnfBfODGtRPE7VmZ8KCl
2eOh7NfF4vHpPCkCyanO7HYt9p+uWCweSDDAPmVPewot9szxL8cHNDmOoZ9c
5aWzbX2zxIGpPvWvzqBzTp34kRJJkAmkioBQA9DfoRp+CJAAqaUbMBYJ5GXg
UZxQ4PrtUdO8U62MU/0dI2pC3wDIlzFOrMUZTZ5FMSoYjzqoT8Iq8TiFQa1N
a8TcF3oR/G2Ay8AfI1Zo9Bdw2qxchi2gfR4PJ8ixO6prqDXNZ6Ilmgb9L9FU
uyRre4AtKLT+m9YMsqSWN1wgTLGf65Grdao/DiFzLXA49p3dhH5zhdsstpmB
tg0ANGmkDOgi6xmxW0EPE0SsbR9ZqRvOeZEGqIg7R7COBBkqidgdru6dpjli
7FFHjk1CK1xdcjFD1VTGgxz0t+Ft/UJ84JXHcKZ/i0aXSXSIykSgDirGTZ5r
f7G8/Kt8joJ5OofFxZY4jk4W32resC4pyIx7mn2dBsI0eVTnqUoj6xdlksMO
9Y2OPptRk3GMP2EkNQoXB9bHVm+IpLh1IUyfS3O99mLCEyzYOQxgrKAODz7D
ft95nfbm3+Y3y3BDzXExb8g8x5PgnkfHJgHDJHflWjwFPZz8k1Anfk+8WHD2
EU8guc+/nKEPoQSAvXHhqmqT22mzwUFSHfPCFDJa4/cNQX//VRkP0BKU+W5f
/D2b+jQrrXoicjM0Hsxj7ZrMX/aHs4aJIqXVSDu4nIsNDUYS5eaXvj3jZc50
VINkGyxmzsc2jLkticUopmFcGjPhWF3bzohkQYCK0nPFDpDHaMih6DOMzLu3
pqBd0hN3BuiwHBqc3cvMcc16OkG28LoUDDddMUzTOiuWN0Nri9dJ4zU/9TCz
/JeYJ92wtfSTHRipRQLZ7kG2vgIWslxMNza+/OLW2TZ/mm/YC8JxchizN/gw
EzSm4wXGezGnZeOpWPlZ4bsRk7TeWmkHqYeDsdpTlSBaWCmTdbUM2y6VJA1g
0fzfmy5b5qCcOc/ZiIFFkbRUSPBhrzsGrQ+6bG3+Arf6ugaw2nG+0UDpOmqb
3z5IaXPD45dJqxZhlFW5nykKdS/ccjq035Olw4mY9v9TI3xBHqf6B6eyAxeK
fZIOrt277ZREHf2qv+0DInGI2cwC+XHtpdExBAhHX87qKlTVPBXQYonapCgi
BNr6JJOg+asaV3HtLEgi6Lt8QQ38VB7Vreg2hCgrHosXKkSSd12fsQXsNwWI
hDaL217KK85hQSyVyTS46sUWDs87+Dnd0xQsdqygwwtB33yJlFNsLug6BWeT
kqywrNryL6OEMkxVwidN2W8kDIIAytOOX0iuZTfU33VZui6tZblpWzKYWucC
onhFehklT4GHJG8XXlUSaehgUM45WF/SZM4yp6u6xQsadX1z3RouDNijlgmk
0onCtjOG8EgOWc7nBtduExtleZHcSjjyESd+CeSt9f4V5I6wM5YzaISuq30m
h1+OW3BWzAFP9IikDqOV6PFP3hdvC7s7H8DXvpCCfn3yI6k3aUruce+uX9BR
aDetMsBV9wKPnI7QcmQyL5Hg0p8sSsSouYbGoKklMt/cPBryiewYCMnyhkT4
C0vj89PATHHTxDf8tErr3m09x/J3+1achpe2xXJm6/crxBzjeSpfYhcZdjr7
FHPyx7oGov5+C3L3SXeUZsEWrI+d0jLQeQmzcGYN93XVdig9X8s+faO80Uho
Vxc8Y7ovUFTU7CC+HoHhSYsnp5DSAUCQqHDIPmf8spdhkHFc234CDcWodLo1
1xuRKCE2kA9n9vIqK6uK+U/mGK5hsE3U8YrZX/pK6ZWWFfa+dXWOnrzx3CyI
XCB2SGeu8OCijuRlUjRhAHjmAKajceL+0lJ4i0uAHJlGW1ywbL2lerBqISo2
WQPkHBmKdZ1XIt3kOGPXfz2rak4xZ+/mVCJYzytUbJsG/UnNqWZCJ2q8MvSl
5UoEHpYEM/fsyBgKOq1qDxx57+CkkAi0s9L8isntIwkPUqshtofcBE3gV4T1
n2InJD1tp59kL0r+WEMs4ZVKwDebJnwMrEvzX7I7xJKHgRBxP0uCs21kFkKO
Mn2CnLhTP37hhAR9IyuYxj1km0ldoV/p4b0DYLQOgueMOR9kvjxtdK6GRtM4
SW2hQpko8eGesX79BswnUv0Oa3yVWCsVpcSTDQeuym9P4LXWxRhkX86EOHwi
p6vvWc7c5Hpoqa0hkvqjZP0ByP2Qg3A8TnBxgn2NHSlam7XxCE0GHiQBGXld
gz809hPzOFvc40hhej80zkJM3n+kixRW9G77iWiBl0CQpZVo/R3HSXaP/5su
kM9MxK65/YY48EXCRQOM18ZC24sBTgCLNoSyhVp7pwhDJhXMqC4AmcFKtCqq
Gabmz0WP7ZV2z8yCD93lX6k75lqXO+XX3UmndTSt/ncLWJjM6+kLfPAJGomB
NBLpnlE9mV3meGYbuR1H59ds+NFAXJ5fA8Tr0mIGu8wDxaAFaxrWOWnuBRT2
WAhvxS+XQ/TuMR0vqgl3IyEq4GFjc3Wo0PZwZxKFc0dNWGVAxrx0rYirdD7l
+LdlOfmExWd+W4do7BGyBjY/bVreDMm+lDCxXRMpIYQ+gy5o+EezHw0+S2q8
r67V686ThtA8Ww6v0kFQCq2dxWzJHv2L8jbpGNlcU5QWJDIh2rzYBMZFtAE0
KwJozIDYDvVAe7bMGfOiQzbVo/ciwUUPIzKWg30g4aYAI+a1IHMbUBs5ulIE
L89tNh/AcFPIKvZr+IXfqQu+hIBRFSaqkVr8Y17ReKvG7hpOzy1t8kUoFiTr
tAlhZlj+flCueMw0+mjEyKXZugvRptIdI/y21ATz7YHL6k82S9Xc3Xs2T1Qw
jVf+QHVXd3X46oWzjLKfHGQwnNajQOSo6ofmz/6LtbT8peqrlvy61powPzZu
hiZCmu5l+ekbM5AwqLbWSlvLEcIpXo8qOO9+P/8GeRZSXKAbQFwIYABg1QGY
ivgc4gpH+NqM9qiW5BJiux+0CQtn4cScysSgVwdnCBWrpWp5EJtf6OrsQ2N7
rWbiFopOaVP6xe+mbiYFvy5RU8qXzCey6QLX523jcH97fLvPe4yOoxLMocfQ
2YS1cb9e3QXhgOow9zPFiOX+dLqqzTfKdQwhFKMb2eTITHGIcip+TDPXnOSf
NRhIUyjrrB+SunVVhyj6ToLLAEoLHIfO4Ba/F/7Fb8+rYiHZ5YuHh68FLFk8
VwJGjEdF1/ZFA+oCHF9SewkI4hUDcIeFRZ+UreHo+QE+ExYLob8a7mFRIyfa
g5KRV9RTTTvqJ9+DlREDG5n0fDtyMt39Uc69nuiOENx8xv/zx2HvwfTrLOjD
bbOFukO6CXakueG50GtJaOG/C/+5UBSIZyBFoVB/cAhOOIzlPzSh3vagMI4J
WV+P38W8xyDdq6GhKrVfzSywmdvkI1sVYrFrjreNIK2emql6ZLfQZ0sM4qeh
rAnYnuz8CRKa8aItipFYA0Ku5WFzx9SQKZdDFaMK2jG6OPsw2gf/KI03nR21
GM0LJAMP15G8CaUHuClcpat8OIYSKSl9CXb9UkHTL3J+jDcygyhR/nKYuYiZ
O5WSpYFjQuIBDc/fqPqKDWGNAhai1eCwKtP5KeBI8BOJibLVzBLGERPwfF+6
zpz9ZNTpBqb0FGniDOMfUoMYOX+BQj14jUjS0oRWJRg6vH1xGE69N9A+lyKw
Q8+nebyXTonfxrT41vz07y7ImTqJ3wqU4YEoipjyxnVRHx66VXL2Brv4Kpkd
bzYFoT4NtKZL7oFguNcTG2wjLBbn9yCHA9vGDGvp6j9cfjB62SeXnLf5b8+5
zz379lTmbUFDX07y70lbesLAQeX9nGC4x1bt5/3rRZiAqygDPbzCmzz5mu7J
IfrCrl77pMdq2Y8Uo6sgT0jOc83xVtjb6OVp06/D0nKM9up328abXLUU7NqR
MR7Oi1hysj39KcSzChInwz94XYHkBJX3lBUbae8D8aDn2oW/N3hPA+U66NvZ
wITwigkcgny3vcuy16tH4iqi/yuxotZxhN1DwWuZ/zg+MDhuFtvVTPyH+q0X
cpGcMpSUXCVlk1P6z2i5WW5/Z7+W09bObR4yg9P+R0KvpQmG1u8DEv4dXqXg
iD4f4L9jLpOmFV7BI0ABynNRpQSCdNousbYWU1DzvT6WBjTOdwRgHngLvCL6
W2qRFRXcOyvoSjvXsYDhTZ3jE10mBX15Uu1cHEEcxSH9AlV5l6Z/rMPqyjRy
8XxKqFisfZCLEHkHESv4+LXhlM90+iKGEWpNJ1ZyUmyoUKWuY7uDfDDS9MuU
pBjqAgqSZva0w+xLi847FmlmKdklRsekQpG12q/4zyw7S7gLF7oN2cFXbwFj
m7q0Bvin5T4oQVaDPJV5623lbrrU3CYoCgsQnZvPXXVsFIz1Dq8sxtOiP7eM
K5/Vcwsse0zx7y3QXw5RF/HSz0+Bc3rvB1pn2hJVJ/o7ROH3vNAz9b7jKO0N
eEqyT1NgE/yreF6dM/csHkkAvZGuDg2tjdG+Gt1GwTIUGjrXgVgMqGGmMl16
h07fZEHzymmJJ41gLtN2BLePc8K+IQ+sMIX1I57yOW4mgeuSAmn+8naezXEm
5wbxjPDdv9TGjtMOX0OB/WCoa5NyzJ2ww2lrME9S58QvJnz/PFSR6UJtXfXr
5Fz222wpWXR7KVMb0mQElxOtXtI/lxqHdIYrLQbw1u8TsXZvIfId/2QvI0QG
jardAybQUJxcqyNkx/RzkmYJcQLhbYxlTLeoGCTIKycVYX7yaDaLmuNZXdas
AWd4AgpOp/VrV3Yie/b+v7lhWYdTKB4FyKbc1c76toFgqRfSIplsC69XBoFX
KN1S5O31xL+cyLVQc5tOAZ0+nYPYEXBJzAPsh7qnjO8St0GQGqGHSHF8RbGs
jS7Uv5iNz/RVVv2Cd+cjLwXp8m+nw7ggtr4g9rZc202sk/VFamI0rAysiaYl
r0zWIr7o8O67gnokavPFjQt9FqzCEHw43Q+QZtIoaVZf4WUsSBa9SUSCR0GY
Q1byUKKZ1R7OKZFw5OtQWwiR09/DEcPJA/YEJOFO4jLK8XkqHxDr6d9ZZJ1x
eZECd31qMUKLIwlodlROfWdjSyy/YTxvJqhQu5LIPxEdyY7pjtVaL/gbKrE6
ppBnxzF3JNP9kNXmnKE39boggRY4Mm/G7aE33vuIbE/T3D6ny2VgRIM+l2Z1
gvVQpDDEpLdGi3fBFN8MUlAyS0WOv3itas60D/pmLAn2Y4taaLLNXSlfcwB5
EPKitm85ZCAy/1BSfNoqjAQO2WQUI9POzPPFbzTV2Ir2pSNkAwSCsVge5crh
OfVspRAra72rQe88BEefKpFX/TjzMxyd6HAGmPl5+LnyNipd/OU/zrSyy15o
MKbzkhHeOh3T1UPjFJAPITf0ZBpsS35YmvRT1H+Zv5o5Evel0+HZufnmtbwS
osNhFLAcjeEx+GWVGJErSAyzC69pb4pYqFG1cMlePsQq9yZQ/Cen0uMcdzYP
xFQ65M1lJuKf5sMjp8HY50I4adjJoSWTByrKxFCA/Ofuh0Re3aUSjGnd7n3O
6METRxyFCN5LZx7wS6UzzAXhHfrDs/fNAnxuKVWH5D6wmV3YQf9qNOve0ME7
+C0WsACcmRQS7gedtvqifKV+VHQK+MQApMJOD2Lbbh4MvnmupYysBk6lNbq/
VQ+vQzWjOLNamEt6zIsl+9/0AZbY7eOrwk+8Y1z56e1Zh4ThhCTXcT9y7/De
a7jWBgkhh4Jbc2lbUenKkSITUk6OSE6w+XtcOfcdRfuOZlB3CUZ/fmXEGcr8
4oKEpB+AqeE5kAnrSmPvsmEj+jOmbEw6dlEi4ZWDT8bwsc470wl2THAxmAwS
LKPs1hFAPi88YqCAIWngSffLrDDhVpzKNZHq2s+qLzR7R1RX2vtiBADR6AXp
F9446lOSHRxpeOnY+jVGVOowFQL2MwEeaKw8VBhiXj1dI3tjumj5PgYxoAOH
CL3T9mBIg2YBmCyxq5Bon6DbhYh8MhHeC2vWHUCtEx+riHd8GSx8porXoA/V
ZVFy17MMgCIlwtph15v3kIdn+1t4bRLzhjcIGk44QrbLQGXoKSrnOWIvDsVC
QN6oOxn46Hzsm86FQXefKuYBxXRuH849lDzQIOwweYhW9yOr92tM9wfT2ALv
ZlpuW/q9uc+16Z8cssroMmyfINs4F+w111ZENqN3ytVixs39UsTnCiDLHbPO
K1rsltiQpwtAIvvKie0GbaS/jI+ov1fBoqMDI/I/E3nwn1C0jnvpBJVJVeAO
0UGc0OQD/F4P7Qv4QCPyvr9UcYrbR3zI3TbRySzIeJQjP7xczRo7FvgKt3wr
I4dV+Cwbcygr45wirO+VQQqE2CDyvg5w71E4ecjMkad7B+NXlBdT9rFrabW6
HGHtTPpU5kcg+CbAdEdRXEKF5qGJWiaQTmBLIzEdO3uS/JG5nsLoMLFB12Kq
pj3yNt13Wy1BTuJKl2mClBbIT6TnFAmrYZ2NiI1NVdK8nBU6WnKiHJ+T1dVC
9XCDoafMjLji7wnzq9JWyLL+EhmHllEqssLlrARjLBXAIKTMCmPXskbDH2f4
2TYx+EWjDYCw+lWVCSlPSAstVjdLBIMsAeXT5KY5OjvOqguQOeJKWd2e3sHF
tnLeEbSKRqBYEjj9kTNIrJi1G+e3w9RjxPgKX8IDvSAxppLgn1rtUwH3+aG6
VRHv4FMHUXvYHsS+chpK/9AEcygDdtJWJ2dcWbrBcpbBKglT4FrmhGQIZS8X
9D/I87i8I/FMP9GyavfAN7jbkOa2O2h260Z8M9UOJPM6x/bHHuKWqjmC9pZa
lt9FwBB15kEstWjcsfOvIEZp4b0esNItlxkZR++65ObfOP7UV7Wgao9G26iL
e1Zbf+G5TjPzWcmNXGJteL7vNig12Hiux3exEtAzEvUNqC6C2F6WobZNlExO
OcTqjAfpu+RyJSttlgqOu+5q+dLLm994fmIcdEMw3J9qIuuyr3pwhH5HgaYB
2v/QU64+J10y2S+vOsJLPec0nmODnc+7wa6jbzsIMsdBMgwlgIfqV34OkLlf
QwF1dh/ly6R1P1BIaRIvw7kZ7lPKdZZCIBdV7Y2Yo3w85tj2dckwT/d2OuZB
Ii3vXTF1Slxchrcr8rk/Ou6sC4GouoSqaPGzDBVeUYhEDpcO12iXiFc2/9Vz
zKHEOWszjxjW7MOxlQnu1diZPIya8utCkuw+mHfwyhoOgtzeHISp4qcFoOek
ECnN5rSF+v0ZkHSYW2rxY11mCCM4buP/Y2eF3BRlhJzHT/SI9less4FdBjX5
WCbwDsQjhZ+jWw4CcOSNgypiBxSC/s7gZJRUwhOhSKNJBteD2e+hl48pW6mJ
kUbOLBQJabXvWhlidvT3p5otgu//vn4cyxWE13D2fM0K+TRaRSImkxU9t9a0
a+iAOFOm1seqraKm2o7bExZdpkBNYIxVgiQU9o4QJju28qvM8gLmYEzLFyw1
JP5YrVij+pFMIpVngvxn7GMc/eahLtMnl9oaWQ13I+HU3/jzGdejCWrn8ypT
uv6WpYzSw6bGnHkqQc91cma/Mkvk9cqY/i2QKDLFbOFbipLJgJLsAFjIVHlC
BPWf79ZDVqJW9HKw2FG06bdT6ncwY9BGs02c/k8oavAgDR98+9kY1m9k7JRC
pHYZmYnpOBfC9RK4zyZ0B4mOPLkuscchkaA0Tcm0szksl2p4KX7pR83mzU9A
xC8wLAba0ENoEjZMfadp3S30znFQ+0KFWLFM2HEXF98/32NDBoxTF9NZDo1U
aRftPJgwTKD9yEXdO270coRq7tmVEdsuVbNNnIYAFKsrGdxSZJvSq2XaGtoo
7ff0WoD/ZVLN2QjuK0qBL0Bw6KN04gJV+GiYX0FQ1aANXd6ImFynOS7/jEns
Ev2O30gkYc9sokl9jmTf1NtOTHBk5et+SF4SH+8Tw/Cv9E4EwbtXT0QWTY8M
SYJQDOJS5ORjufxkEDygSBG1nboUxvFiqkg6adpx8uH6ndt/XRcYfEdeua2U
F/BEtql9S2t8HeqMTquQBD2ntoKOOsoacuIyh3AhdYpTX4FbF/+rxAZfF/0J
AC0DReGCRE5d+e0NSLbt7J1jIOcabYitOtsbLxqnTWULPDUS7GYWU6I0cpcz
5Diq7F4c+smnlSfklJAO/TXa+vo9ZYmTbOv94AmFlNOabraYvJWS7bZOSByY
xoi5Yeae7trQGqtI3EKH2uWVLkYdP/MJsX6vBRzjv0CpSwvJZznpyr9XzDIK
TJfiLIEvZ8HYdTIHGF4gzfhBk36nL6eIMk2WYftfhzJzMjFwqyg8MWmlxIw8
eq0gUPdvijaEsVCPjzwlOz1cCA1wlRHxCHwZrM0tLwpHyB2ntJ731ufLP+Mt
s6SQud+hplc4RhC11vLFWUxl9CsU9kmpzp6DGN8gh/SfePWiysYZ+3dBYyDF
MvasyrFMm3ovpnnmpMIY2gKD7uKpQIf8p+VbeS+s3Dbaw6E+5/0Fo/moSY4F
IlSdlcuiQOWhYbdm14nCcZg4eZshpsIZX0ZzPkQ9bUcs3zyIWUFyyxe+nfFi
WlboOXpLyUzGeihk3suYHvMNcnPBmjHMffnw861gv9fpdWB0sBQpLh00XlKc
izo1HkCocKUtfDwDTqf4FVH2jb0QDuLgb9/qK1KKRTLf8dIKwxFOMvTRo/O2
EaFAiaDpW2KjVSMV6YADSpygx5UachT380hz/deugwjVXKU9PONeKU6zkWiG
kwnnFy2TemErbFjj26AOZtfCXTs1L1DxeCMvmDwUEggMkqsYBFg44smkDNG4
fbjQ6KcrPYICc30Nbfb3u4m7t7NN6xqovik/kZ2CG2YLxtu2R9WRu85Qt1GZ
U2qn6wpR/ADCqTzt99dOMinUdTyAniEB9QocDAI0hTtSQ8QrLu4ZHj6dk3i0
o87Y82ak536xhUyoSJKnXNfijIb2m7vpT7FaBM8+0gI/4vxS9zXNmkEi4TzQ
u0szf4u0i9K6k1AC6NZaMS1gTwEfxmweLMV10OA3wuZR8AGpngKoQr80eqy5
csoDHkt2I/sBY2x8d711oJOrtgN5qlFaxB64kr9Dlbga/7L/G6VjUpYdHPgU
y+Ra3e2SK31fjmoTRVRdJCuAClb4UN3BWV9ijq3ELaVxCr0sX4baU7QkVUDb
z/VAaI2Xqppor1mVRFG1S2/kLgCd6r3d0Wt0q8qOx827UIQTni7lKvmq7DsE
GTuS45qISStRaJ0iNfZDLXJY4+GxlGlMGQbmZnAmSKrbEuMzkHRyTiXGDVsy
7BZ4mwbX8iFGfNwjyDjhyUqA/8BW7e97aSR7cfmqiatPrKOpA1euNkVU6hqp
oErjwohBwn4NOoGHq04XtCJSfvY0bm1lScjJPmNDlBYc1JLBGEa0iEoZatZ/
cjDt7Mf/mSaDicXR3cfM5HOCgrA7ZFIxUfmNvu/6+T/RXZu309lEJv1jtC97
CqTUWY9VEM2dPz8k8BhoerRbRt0R82O9wRGCnA3qov3Ox9SW7TTpZTOgUdMx
isXYsO1hHd0QgyZazKjGj3NfzuNTCqPv4AIz6NvedsvGhV/50nx33duEqKbQ
n6caR1HbFlY66sJTGYfa2FIdA83dfKu+rSvQRligYgOhi+h8kIcAA9QYnBHu
KgtgBDqD7SsGD0IyynMuCPXM9d5HKwzGw+9IcZyN4eiwXLzYFZ92PmH/IwUs
AamaL8Nu2WyMiz+7KKGjvhSMzra9ClePL/EuzVSmABl/+1L7MNCDiWlgqa7D
waDWQ5uuGx2+6iKIgQ3b8RNV4Ye6MIhjVtYBspiAapnYsstH07mlmHPRJWIL
dDhfJhGk/ShncZohxw7kjtOCe6al3ntUfyR9BhFoxY/yjAb9hX0xuaMVadD8
iKA2CxRrfiLJTy6A4ZfLSzbuNlPGNg+WnmW2g2x7cUmF9vEuLyt4tlQCLlMh
vjZZbY00kMmrMvZXXZ3VS2YCa3Ef6iU4e4x/CQiVIHjjmHTMX8k6nmp1ri4E
Y4Hy3yGY12t2RkRGpXaAaJQjEtz2V++TqtxRVGJTcto/4sHv094SLIZ+5wLz
zoBHFfxKGqL99e18objO6jk7uaMdAS5AumCFSDJDxGjkxwaEN1A7hWOXGVlZ
8U1J6WSmUc3QQttWlG4NzdPf68NxwYEyJN8s6k9Lza+Ts2gx4csd3ACoOhQf
UBpeG0ifqG1HK5rKKblEiQ+eKCqIzywQpyi5zz0IZXNUvsdjRZuVP1bwRf1S
h/AUSqzWrXuxUTPAk9C2DaB++DgDeNRTY6Ut6F3nfB5VIVZMRLX9Zmjw3UrT
f37+LGNlbv9Q8EFvhxOw2JTZjjfUNkBodE41TIM4BZVVg8mmtpUDBo5tvSSU
vobQYjhqgdcq5/uXkgEI1SFch7W9lg87LQp650Kmt6mmsvH3dujpXG0opTPr
UI3AqAyp6j76K660LmLvqHIbRfSZ1hN8/FClHxIV08oTaBAQzj+NgNDOExFz
4s3u7/2gb/jpmYlOZgxD3UO+ZWDind90Q4WbAOVbeJXXfDDnOhWQX+2QT1ya
uBihFCdkBsWpla4eHzTqJst/UQQudIR5N1ZxKbsgoAHZoakiXYj2Zy805Tn0
WeSTyEFSQAzKYJvLXdrCWO6bKlCxSkw0KYIkzzH4kAuJV6xP4twjuJrJt2+9
kdImIagOwhXbKC1Q1HysARuv/cJaJIpKi7AxpjfohK5g/oyJ4xFSLhVxDpkv
cPQ1UxW73Kx+eMh8jZxXvBUdFZaHj0Z/q7Kff5aNoG+8In/xt+jcqCu2zHN8
larDZH32kuMwmxTXZoQojJuyb+04ahPxcIWczxcqTmpQOC/TtNnzmVFTz9Fe
XJajgkSU12Jn/TaVnyHvxB+2oG83IuC4TlRD8wfHfs+Uo2FI0rHPcyZf7tC3
EKcr5FiL0ZuKD/0gvUc1a8eldE1AD54NgKybSQ2bwGmKhJHxJuVsyvqwQFWa
ATOQOZVI1XKXb10fCR7pyqK7y44R7FJxRBO5wKG5jPrUHG354EWn/0wPS979
PM8ULs3RRp0ZbTi+YAGYeg1mma7JFWOVi5YEARh+fGGMYnL8XgQvrcW52Z2i
iOsxzXQihGeMZPWUrO2W0mfKcO0Mz8shMXqCmN2KIY+Ku82LbJ2adEqsHCEN
CFCGJdesX1sShpf9K5PUpTBCWb0D+g+FOhUuV6fMoZtLxcHRuYIh285zNSUK
YAJWVu7mcEInWB6OgEGyWZDJBd6SU0CBVaFVgtWVFd1W7qWtOpJD7nNvsTT7
ArU5KZ0iIvtZDc7TG8PeYGiEkso+zRsZMjFBFhnu9fIHXsN+5Fvge7H138U+
EERKI8qaNIu4S3fq+JPJFbAB3D28eYGu6SjHZX4zjgDpzhKUhCCUCQGqob4s
CXsAqt7Om6oI0ZfU7iUhkre6xXDznFUIdcmoIEPkuhwwqEIxoL/5V5abWnuv
dWCfHWw4YjkLteQtK8t9A52xGhWHATijcG2NF5wkyd/47DZL4MuKitvGlMwl
h2bcLs1jxTO16uTzLuzL1cNZS0JAi1G6bDh1Fw2azYZO9mSjhdRwnEklSYKj
hh0m9v1T1OFZBtYShTlLphZPzTxjwshXNy6xajzmSPwlSvvIBAaGW2j0h3gq
x54LBSxJLSRh9UenQ+NmPzwRMJy1AOM/3cCbKW3v8rq5RozEEwhVR5kEbkxZ
Wp+M0MpRgSAChfL/2OA/pHTwpFC+GyDhKgAjMBeytClzuUPVOe3ZjcVoY9fi
qlgWcRRV/rRTWwLBrH/LBhQNSKZXNim+hvN8yXPfBb8arX+WeJilKE8l0f2g
sKHt3focmu4fh5Z5RlIcGy7uq/jXU9iD+G/XI+DIkWczyR7JIUzQbe3Il61P
3AgG2RdAtGas81xGicFe+btxij8CJDjy5LdYpN2KNBv1Df4Gx7NnAnBI6tJ0
fTYYN4VNl+PDTpLguDbAKSAnYsu/v53BNEWMFeA/afPIshhzBIXGoRSeMywj
Ox++W29QJm9Anvd5hBhBiEKGRWzEDp59JMU/OAzy2sf1z+gX80JAhtEAQp4s
vGIZE9aA+h/9LJmpsZNNOH/hpVR54X/OcGbhG0ovJxr1gvQXMsPxF8FCGq7s
leLtkKY5KkxmeD9eu0WMPYjQkP8Qr5RdPNq+T/sS9g7wjC2fCHtF0jEMx34y
Ur8rQkdwKzdtMUpVzENf037qotNlySab1T6vdsBxOlxzJOanobv9E3Rf3m2u
amJ3Uu8nXueS3ITjyo5RyptF2xJGtR1Ed+WE1RtDuy6cXTTTpzng2VK0VN0L
giRVRxmJg3K6xLxurvvAYNjrPvLG8gcSS4tOGQFzwxcL60BXSsWyaQwvCTEF
JPcjb2luDbR7IB/+TiJ4HpO6T8UkE2gFNZu5AJVJHkXfo60fd3hoo2biuAP8
C1mr4Cf7TqGmbJnJu0K8O1QZCaDIN+zaG0pMX9DvKtIG1l8ZdaZrMLeIKNz6
Zd//4iQZXRsCfBJp5nzwPFM5Xn77bvv6EdT/BWI5kJ0AKrbyED3BIJwf5lwh
2hgjxo5iDWVrymCO+KyDPosZ9Rw5FR+4wfe6bhxndnVszb+RteBEFTfyFLic
86cYjbEAdOC2ISOep0GLCdb2rQ1h1B3pJsbVvwggWyVqxZdd726wmcvDy8Bg
WpeY/Slo6QHdEwqHSzZsFJzT+8c7QGXT82vgmZcMvqT+zTYuy8dX7dZj+1sY
yP07Qy7H2+0DgOlfPA4E8Pz1j87Svp5nCBkmJQe1eivGmiMq2yZrWP0aj2a1
SMnE+BYVHfWxE/niIsiOqollQCh8yaLzOtM8SpHM3xh8NHdnuKd/Vo+2o94h
4XN5l8QLd8I6iq7YxfgCzJRRuGx06T0KUBpyMTHFXXBhSWTKvaK6GqSdQpjg
tlr2r/elgrnpmog2hS454UvqLCTDc2m9nWlYS6e/BfrY41CzmJoEY+07pAu9
LVSXHDv2o5h+mQ15/y4NK9wyuxnqkzHLB8TJ/G0n/Wf8FFhGdu/j97TCuCX0
mDVsdbynZvmYM7plzAoKGoFKEEIhVrnryVzrQHmxY9Dc5RjgW49GNSk+VBQp
qlhv1dwfJWJ/OuKcx6jgyQKFgfbgfooIVhsSXFcFNIlB12ZIU+ra8yOmHX11
0jLoc6QIK8ZFG7uETbzHtZq0XEbCco6oNygQfRAu75mDEJC42bPPMh+U+w3U
0+T6KbheXCEb5qRVHSDuL143hatkO93aYgWi/dQbymH9Auiz+lgs5xug2wRR
WMuAsg8mqTJ4Ts5pkk7Je9Pq5Yttv2RZrhBdK1aHGfLv/Wg4PU6ZzDudVA3G
11AvJf0AImJu3akd1R1wlxkGRzLO5lzkQd49skXDWc6JVa+SYNUD1f9YJJUA
1GPTeRaP6ovepd+YhB4RHQ8V5lMlxKVmk2lhgqoWky5QVCWcGbTJ/GLflTYu
KNh9Lu0g7OXgAHI87LredavaI2nnI60BPswF9cLNeS9BtmcV9BkR55kZIxjc
Oqlch4nPCZHa163HR9GVNfE2XPnaWryQc+adKxvxg1fb2Wgediyn3O5liBc/
NgdEWFqmUdQ0RmY3VXFzB67AUNjw1dgga0QZlK9BJPqlKGn+l+gH9fkPmkPt
pU4g+7iXioDftPrdONm2fjL+/t36xRFotaiY7T5klNk9R2x4sOGibi+kM5/7
+hkNHJvWammsQTy3Cez0L6v2y1PrPYW7DuUPfjPVnr5608JdXum4WH7UxcDd
rHwmniEG1+CmzZkSEeyvShGaE52VI8laIOEFC/o/CyCgjU49gqL1qod0j5QD
toL3m38jKSa+MPY8bhbdnhEns9CcjaLCtxWDhCjJbEYgYUMaKRX0UApkjwI6
Y0/pNI3IpOyZ1Xc6mw/l9fCRDihHMEi4eNeJN4HNdHKHt/Rz6JB/EqHLKd4Z
Shmy1pOah7SeW1MoV/LEx+pf9OmXhgRJXmzSma2m1rfN0uE7KHiOA+kYQu3d
ha1sepoMNACOzw9YGJyGL1byenQmIUS2SMjJ/b0mZB5RbU+qtjZmfbJKL5/9
ei9W05nKTsxIpVL+32NDRpKDnOldmYFnhyA5y7dGaWcOW3PFWQa5HDnu79T+
pvbC9g4rIxFNWxegc/SDBcf16x7UK5Bv2Gdx6D8tJGQoHngdns9hZdS3V+jj
048gsbgx/+rGC9FahYeJAumMJAu3vsHGk4jI4a7jBt53i0fTVSB7g03dZ6Om
d2DijFYd5g3ArVPxHLMiSTRRjyCKluW5IeWxinZ1AJ4uHOet7+bdo/o4UsnF
L4p6HUpElHUIvUEFzRXiEv20PfogGOwF274PITrDMAYyHHDMDkgozZ7eZqzd
aoBgg5fk3wS5Ft55ngyFOYj9PTEbWmnZKXPfPdBb4SNxdpCFrWVsVF4hOoG0
vBlElKgcutfkLZIRX7nv8Gx2/nlFCBYqAksD1AunD0xaLNGXcF+JiXL38lPc
cQ9HM77895Mp+ZGqoap1VjsWLuiAc6YeyKpoVW/TmbbqiTMPtlNfQdGJZG2M
J2rcs1XCrzzD5VTbigMELabK31XlfUMfsSOSX0Rl6rmndT7pUi6gkd7MYAHt
7qTMtCDQR19q8Tz6gPJAI9LPvTI4rpCOwpv5vuDgRln3UGwdm3ym+oHCb2Wb
8dNvqqV/jmgbhUhn7ppE5CjI55shu1ZcYe7miHcizyc04rvvGzifj68K5jF+
Sx5FScyD86bFXJnEuC1N5g72BUcAjJCYQICgRjlJGPzDKqOnoN0xcdTxaTsY
iWZMEzU5/2xErCtw3muCNG9XHwplL907MVxIR/JW7cztZA1gHYJNoVUPi9Zk
pmWEX3EWpcH53YvTtRZloZ0Nn31Pjy86B8FSkUEI//AUxDQayD3QkDAvA85u
0tsM3a47RZ405qdibJAqvB7CJb2bB+bGp5+6RyMLQFqQcc+IEfdj1BhG9oQK
lOHgZfeBBqwAXwvnOeEzlHyPTRx92QA4Rfeauve2+VNumzpD7cjA5Tn3fOig
J2gIxibjKiMkpnfvunSzixdHstDDlwDhlut4NT2R4UwB2MUWVMQDv/vYSFwV
up+72kZPAw56Q5ZSX2o7pfbS86J3jYvRJ1b8fR+hHpAphzJmU/8g7nKcl5sw
cJ74ar+4gyitV/wsz5zhiHW6Zr1YgD0sWxuH6BJW2Vg2Y2qIWjrZZ+LdI8as
OcmDpkv7TogKYZRA/8f5tnI4CnAYM3gz5KaA+dSWQxmX5/2N0JdjV0isN1JR
capsJijTHfYmwZKhfxiUm7IIlX35D8/p05D0x9GBi76bNnupXTk2qQrpyup3
ZDVtjdIh25GPyGEy5PCvUTodFCGN59Vx6+ZNjUSiIe3ez2xQpDx2BF8+oJ6u
5zOxW2yJWZbZvzSosp+Nl9BlqPc/i9F/FRAC+pxQ00tJgsF4OzGPjn54S1RQ
11uSmb4k/w4fp7OHLJSqaS9Fhm9kG3YjIEuJRJZyoquOhlQySHNIaQPTqsQv
SiyF8UVlWL2Wc9TIP2DyaVFkCJ3EUGSmUIYZw2TGmdZ1e2S0oVB79e43kpUf
nA9wfY0Xhw08UKc4TpfV5ZfUpSwV+eJup2aRCLwc3rOx9Rus9zzCOdvDdvTo
z8XPAI67BNl7oD9XVH0FhcmEIHFQ4tTqpsIov/Dlp+YZPfEBafopNRrAjixL
9A/MLP4QJTmhonYuDPeWwyHYoKDDk4343ligjdaG/eiWlWw56rEddzeQh/kq
Vbh55W7/asZzdmfM9MKPThq3rF+TmQUzZNGj3BDslHWOAi6gJOGAtPsqC1Y4
roBvs3N9zeUFMBxSzChaG78bQ0tpPZZWZRsD/GG/OYmU7r0shMaP0JijjKPe
Zwc8ypbqyS5T8FfSftLFb3WNOtMkheyItw1OK4JHz3KoheRH+p/8eG6YWQyT
lFbFW66n0zNRz5US+zs3onryH65AE6iG28gmFWU8VpywBo0tmm1tSv03agRM
eVImUhcaX1Ii6gUt8q8vtOxyF5bRC+AZCodhur1b4qB1AouFGqbCersjstOd
yaNtgHxWvnkaN9Csw6ECS0ISMCVlPY5n4OiKXJ2BaV6tf1Vqhlg0v6Qu56e6
46lj23aKN/xzOqkwqapB7XvDcAyWcMF2J5EtJMsWAvwnpf287CI5QvafZPf0
QmufJV73LROD05FEFTirLMeCDBw57/CFRi2aYRHu/UIpmANSu6eAB7ElYx9o
vBTzjmU85oOeoGy0E5oTRr29hxbLqDdgIGpGYOyadsogYqQtcpl2ElVeCOlf
SQBNnmN5yBq+b/dtmJSLcxhLpvzxLwDcQDCWUGqS5s/eBxTVWQ8oTZ5raIWW
lB5I/nR2EY+GDFkZvQqeJle0CWwI1yjQTVgcUtOVa0F+eoJMylgtQw64a/F5
Ng/Pk4wCj8epgVpqJ9Tll/b9DLke7n2WWWnacTOeDJ8BpRZzjlAlXsmlLQvg
C/MjN3elSfOi36tWBqKza2WTHjSYvqGfNV9z9aBd0LoNtLuQrNLE4K/xRPR5
8jXKWWU5f3U7yuv45DJf/27x+m3g2wrHFY8MpjUyCqfFToMN6ow1fMVpCXkw
mvopYBWfxXW8I4moe/7P133YOfUdJJOqG2eztTTPQllc8ChdLIdNzPa57pH5
BUz4UrlYDU/1Zc3U+FhAVIfadEj0jh2ytg46VSmKUaJ2IyDeBkI+vUII8HM/
eVaSIrOFLqdsXo9jv8rDVsu8JupWoy3sw2ugkfNY2RqSXF4t8EoPcgyqG+eI
oP/249Li02B85tZjBfXOPpuapJFISOkYtywN7DsPkI6RT3/aINaA+JOcKtVb
eLSxSektmpI9GoA6J9A1EZcqkN2+e0h++BtAcfMpCKaAl2/r8Kk5ab289dIV
NOURA27+fcmpDCaB8OAcFPELJBOqEbbUyHOGmG68iB4bKY9PYIfhLtHNY2fG
DqWXuill1rwk2LXdkuECC3OD2yy2IkgXKGHQ4KgGzH02tXlhpQ5Lns9fZymI
8MgkocYZdqxu+h2BN9qLJt4FwtcZQl3y971CwtuGmMzuY4fGKorgM6nuEhMq
kSkkpOLpYIn/JeNq9Tued+rr1X7DJj0BmZgNnE01Lxb/mzGCE2csHCz4KsCf
ZAMTqC3DKJvuIyBPdRI/KEPKOUtHhPjsXB3YEZQxl3b1zoxCqqePfZdon1kk
BIWQGXMzJuA5z39XiYkuqDJZzt9yE58H03JZVPtEP7gNtRpnFXUufQiAOJNy
y8K5kZ256NfXG7nrn00ZAhr/mGTI5Mw+rRnxEyILrX+o/+sibc6cy5Dtsaed
WvcFVdcfvARgaiL7/pyzvarK3+iRrxclbGKvlX7wWwQzFi5AgCm0W4C/Kr1Z
KuCobXx8BpBwta+2LkzU8pSwNktHGwr2BL79fJoOQCJo6FXwRiIepHYd4Jb3
SLuAgcsqwkEesNDl7aodk+dj+0P0YgohJB+rpWOJax1tOcOxqfVUdeS8GhRL
uCVW2lhyHziuXFgtqA4Fu+KR2vfMxsXjMYISJ9mRJ+MjImrcM/8k248bnFFz
vg/JXbqy2fNYjQ8zJUEBpm/FO2csE+H8KFq4xWrkfabmTQIuUbzWdq7bxiyz
x49uALYmOKk0IAbZlwZwUXndrJAKi53VietIope/0f4sQ9y9vHyr6B8tTFsL
qFnYz9c7hgvF5F1WqnCMKDy/hFPyFiavVvwjuWlB2WS/yBK0mg9zYGZW/36e
8uWJ+F1jzBq257gs+vJ7/aYjfPVtwBgwoLWDdmZh2p8jI00HLMlb/ryhRi5Q
s37xcWutr/O6mcHbOMk31aFzhEE8An/XTusgjR3lfcGY8a12fpRw4zGJIcQU
p79WHPtLNZyPKnAsGMhEIVFAPuzhSgTLfHwN0IaAiwgON29wwWJw9LZEUx8a
Q+c9i6nSFfWKaRLY038YBf/vy6dEEaVhKtqNO9fw623mBFzWu4Pai2RYoQjh
FgW6M+4p8zQPLZp/QwZhvteXM8mZbh3rHyAZKu1aaQPEJmLEoeZBC5p4dE7o
sMNxFJkvU26boXkyA4PkXKhkgc30hs7olbzCHDZE2jHb5wGdDXaOdMRfjtV/
RUIBhNFJYaYo+pZ1If8+Mt4JbVvHsugjbENs4vp8rBVMk7wt8o6d13vZFqMs
/Q4s5nsDnzsS9xeusJ+hbxq8i9+BK/KByBMN8bOrusXIte41E87G8QvBCT9Z
vRC7xLa+ph/eYMZE5Bv0qp+HNTVnqoU+qrRLq38SrgbAEId50oMN8XBofZUH
17ugLylHtTTp2NuaccNVJo6A42mk6JZXVSlazP5+DcPhB2oD/iTrtNCEX2we
71dWW6f+O1uuKU/eZHk1JvEJu9ugZcsPXoolbu0Rc0qP0qWxbcEZKddoSiqG
paDKYeWNX9OMbP4bjeb8fvwQu2HspoVQTUKQ2GtLb3zuw8tZDZFXLoyR07dJ
8hJkdHE4pcZRt6m4y8koh625tNatPSHLb0duOt3YF4TbKFJ4Mxds4qewbY1K
aYfr7x25g/C6WRAZ5JBV2DFQubYgnYTixTcqalrgVum4He7Cq6L2v14F+sBI
nQHMAPF3zz4wzTzikVWjY+cu2nZIQxqsiB7wpI4aNWxuAJ9MUmUuQh8rrJcv
CXyg7O6wDA27VtgJrQa1yIuTqrm41n4EafnjP0LPWyaURlhydz36yB0OnYQx
5LnyL16HmIhIMdW80hQi94N27ONwjglbziDczAyCmGL5AqAkYS2eII9xgFpc
5Sdp+cDSgUCaX+07lJegZSbq3PdxOSmENrx8H4QHbiLCFQAv4qB6uQMLmsLb
C0v0SSnIJZPtkltHanxbG6+yWPf+0jo1k/aT//sRhBvYZSEJ2+MmxuAc2lpd
Q2Uvn5jtslwmX0m/aSdJBR4ZcDKpk3IQYGME3IkSGL2gjQSJTKydukA4wLCM
zDuYl3luu7r59ztE0yEZAKJn1GQUp1y2mSwaioa4fBiNBEwMjh0bP8Km6BI7
NEjP0UELWMbeWnGtM4bsieiCtmj5IcoE/OeM7jgpyCCofU5zFi0qg9D1n8LY
+vGdBvpBUYDhh+jYWspFNvavd+1iolOnOiZi7BT4bh5jxAFRpnKqhpx6+zvF
Nuy9GKvMjyF9U/fGpeiZhgUFpMZYcFhJcOgut5T2d6FMG4nV4SZAWlALGStc
2lvg8S+Ka3DMTiyRijO4gn1wSJNiA810GXuGCr+jcXFLPxsxH7P79dvofAl6
qshFdCdKYGOxu0x/HsdWy+1szA5ztekMHjTzCHNk4slmGL7W0Dw/4O/vIZwd
BaDJW5nFyINlhYwSKdysR4x+HjJoriRC3EryGiO/H/iHv2LMlZHp2NPlSkr0
ZJBW3l+tqJXyIjAZOnXFa+QQH7Q0kxIf9vXEDRyuMXKs2p3GWDSr5Gz2UzLB
RDQAWOOTyv3guEgqMjyA2PkJ+FDu/v6AKoc4O+jzhKv+dWafxSHm211Fcd8v
KQWuG+vCF+LatcNJg1xY7TGDn2UVzSdVCCTnqdQERJe17CsZpLGDJuoSCJy2
aZXBxH+O010mhcGx2ZqCvl5sHWpEd3X8EbgmJTp9TJew4oqEg9DwvvyFlqUn
CmQZ7wKSrE5hFVis0xHKuQENRK7AdPfJCrJBaHKA2UGaJ2w2//vh7BQRjA70
TResryvIPVer4iKnuHbJN2vRMzfyeNSs9TfKXETaUHWA/CEJTskWGrNgpMeV
yYa2qfMRhKh/fjYrMoCHuwLXD3qNtZNWDO6pnsceUD99WUEm76ATHjSWlK8X
uhTl4eREWbPi7pNgQubpikv2LNSj5ud+eF1uMzgn/mF7UJVFcEo57Q1ez4z8
DwwfIE5py22Zui5+bPMXgVucaGbSDOrHW43ieVRKHfOFD0l1Szlyld/T7EFO
W+01PzhUZeyeziLE+8P+cNqaeFr05cSGe1Dv9512jntQx0gb6KA/CzefAPsF
89aBeOHOLm4ZxTIkPNeA9/yEnxkokNk8C8+MyRVKdyiUoreWrS+CdcjgISP1
OhK7nn842wkM+i8ATfKAER/dUcGHphljW8ArCIXWn/nKjHJ1SQFhXC2bFERG
8y/xVoYRgWgqmsMuv04vY8KpR9B7A0VpNjT4h0uBNRLMUVilGFVFPJv1CBlt
jnhd5nxg740EXcFkIODwEEoi+q2dJi3DZadN5/ITfkTZj1W9o2paIMhoVrwh
p9y23dprJMBhRSEOPWNtfdRCGnRbaIxrMg1QEJf+DPESGkh9TnbSDXVprnFg
WjuDzIYhml1CCI+18l17MG7FJBrdwUpB0Fb29Zv/+cZLL8jycJvq0OshGk04
V0eMnbWRULMm98kGJtdvejHpE9Hiod0IzNmMdfpHVObKwaprU/M5Zk7lFc3z
/XSVULoDK9H8CczWpAOCJSaAqsB7VuBYaF5eqgRO0lTuCMWFjYY9h6lpVelr
B9ssFlkYqLPwr6+OAD0KGCMaO5x+X8LHsS6eT9hDutaoqzO5tlztUu1yk3OZ
zocAi5+7Fem0idLBZVfLpu3e+AJoYj8Yuh4exSJyiYBHz+EOX0ySrBeThmB0
Cl1sKiuKa20pcQtzrBAlFmHQ4LRbtKqxHsCljAHaPugVwN75bkHWorCT8aVt
wgftW+BJTHoX8LDPWU40gUdgFobpV7F4NsU38clxe//cR0fmdVKTSiIon4rI
q9sZqr6E0xAWQJF2LnAU3qLppDjvq+TJhecRCgD0qnu/bVU31fMsnSnwv3Gv
l5HNvMVOlFW3sfxPULiivQL72n5H3o1irUQhxmerr5nITXTntmSAK0cwXGMe
FCuQpk5bFwOrNk1yLQOsn9WitcTgLDb0vyOCP2uKyShFt1DzVkSeC9H5zOwo
w64eytebc3jXLdtYTX4eTN56BmDt5MVbWNtcQCBkjw+W1jZrospymEXqjDBA
G3yM2RCknh9t1IwFbaSyZaNYJYhUkK67d3meri/kQgenhpU6S/V1S639B7MZ
kp5uRJVhT2AR3Rl3nV9dKBRhQlFb0sN3ZMRWv4Vy89z7f4zdrgTfe60em6sj
JuGAbC1N+UQ6LUk0mYbr8qEx7ULlRpCftvMlHTDUgLjKKrRtFa2tD2jCcTb7
DTly7ah5EGVeI6LTXPPdCYfqrHha96sHTobnApiO8fgaFd7u5Zaf6NV8eot2
OMYb69MfRvJMTD4xF+PaKUJYuBEKE5fchmLwrpe4aa50j+y24sbwGMHYQdh9
jvwwIuU3PviTv6a0Du5zJliI8z2AUwXE8vlARK69NVWUlxd6ZayDb6p5ze+q
kpYZXWhMm5N1f+rqQ7lQYyaNjrv9R9yCuMvGd2esdEe1f2rk0LX/ED1W7BPg
tsXHxvwNNuFjoKB7zEqbRwo7vxhUv5uBTjxsJGngri7Or8MBZgVYLfPmrjFO
rbj/gkaSmUFPUmOofnwPG/DkR5M3Sl64xuf/yLxzDXksl9/ouW4j6ZEtBmmT
JEIdaX3cm5n0yqXGvdUXgk6f7CBDrvQqP3lf+PajCAmVVBLNfGoPo/ImbkiA
H0n14b+FAr4S9XuyqgPkxZySt83n8Cq/W3mQva8wrKDkVLnib9XNQPE9Uk/G
x4tLeuZG9JNffXtEDT7bAmQO85zyponIvB630g7YC0dtQ8P3ZPWBO7ij3OE3
B9kwBzdaP2EN9VcdiUT7xjjLl44FZpc2/zl04DaBPc2niqe27kI7ggwrkPGw
1NE3WdADY5DPyjLFRIzxRDMP+YeQTZj/QI4JO/8In4yW8cjHSWYK+TMRUp3b
zgVGQ/plFDSt+888T+fr/GP/Oi/KmNu/quJohVI/ogPe6JxULnq6YW2Ln9N9
UKnw73NLIo2dp+AwWc10If8uX58WGfVH80WgfzbbNOEoOUcnT36SlEh8byne
D0kiMlftAYC72f+TDdzAj9qMlGgxYRz+DN63BCNgXIH2cRwMkT8g0cfpdbi2
39oM0Kxv4yqQ0hIryIMn2Ysa+ySjeFrPmWgRlrhQLwAE8cugyGN1yVDdflgx
2c1lWkT/je3ssDelRlk9SkQf/IYTT0XEvP1FhfMCPTchGFvazEWzh+ukIVIB
CDtaiHOo93Ra46tGXfvYrfXf45taOqF7ZttODx3fs60jvy9P8UfPDn+VbG4U
+1TCKMw8Oh/yl1g9KwQ4nn0NYO05rLUdpSpGiYLrtiMsPUmzhjAFTiUj2jUW
SKSBwf5PaikG+AlFkFrFfpkTUI2VTUhUf0Mt+bL2f418jTNkgyMqAu14M2FI
ONW8I1t/59KPo1mSgDeUlTeoD7CVBTcnwaRowOoKvqxXfFV+zu1XJIG9lK90
iek2j149wyqv4sQ+JjfYUWLzI5QEkrpNWF9r3j/kNXsMDWDCeT7E2VhPcSe5
4XJomiN3hCrVeWtOplgKrGfJZiwel3Xo5m2wxSxwdpy1zhqJykZNyRlwdF5E
8ICeChQ746fzZYTx+L3pRz3PO5oEGbY93Vwixu6luDJYgPhlGzd7qA4C9xWd
uiMLphMmrMMsmrHKCaUUmNtnxkDT4WRkT5uxhfO8YWujQmLWrOcNJEVCOUAm
RIIdp5y8kuktHigwHJEAwEsvyYptd06yS/Nse54zbU9thHnbuXgxnfg2K+PX
4nTylfY0Nv60A+297Qov3FKwsBSLK38b15i/ySHduBz02TJTPjYWKURg5aqs
jrdVzvvB/kuUyERfrkx2xp5GBLgk3Z8Al5uh6u7VaWqfzIVkR81Ue3YKtF23
TGv83tKQGRNuXVYYLKpZFnxzlfgHyepz4/LFe1yXhoSr1HCRyB7awTg5Yi0n
0VxQzaRX9zOViCnv84LLQsgoF093Y29DVtp5lqf2kmiom2Il4J86x647JHvH
4DCED8ija/yyoud9chYCVZPyidVZLvZ3kE9RRAiA+FpJ3LmF1Q7QXtJXkpJa
yAZtNLssS2ZRzXw9Oi7Bd1RQFvxoTEbrcXPU72T/foGPDKr5USqIRw81OHAD
J6bPVeT4ymgPe9PBHGpFWjonx4rztk9bv/399RqjMsRWwhIQe+hU/eSqfg0h
Iuz4qqUkIiGqiTQqEjOrXXj4gsIYoLh1aPBKVgwC/IL+GAW9Wi187AnmsxsX
avpBxj9djFhSUJpEXnor5q1cWlV1RU/HwrukrUhey6ujsWkwPqi0fcHeNnu6
fDPjkVzH14iEZtGZz0MWBvS5lRX3EuGhfQY8kRmd3aILViHA6UI1sLvScVU/
AWE1brUs63Qz9UBJvXFNAa4HmJ0Z54tY1eRJlD0qGfljFnfd1sem0UQlcwUc
cLkqWFm8bZIHBmj+NAocYINjq04rC4kGa4Klt0IlusDSWLR2Xb6IeuZ32U42
ahI35DcUvUvQ69rPosXB/pehcXEAyP1JojuI4xhbU9nwhOOhX38yzgjZJvch
RqclsVlVsOvinziSP0mOwToOSAYmQmrEFQ5d2orXh/uVhX7Keph/lxjW9z9a
4eSX50kpnxO/IsH8Y5MWDTUwdpsvaVofm+wi5lO0YL2xkolpRE24PE6OSUta
k7JSdDnFS1qFSOSem408+RV+BHnmi7FaKTfL4OKR1bpDSXDrUcJbYqE2aAfs
gfTk3HBzWc+YhoisyGUd6XGUByRgcAl1LLW4ipA5HikRm9/2CH42d76HtNso
is6rHDizkXGolXlk3XG6VX2zPbhc5jpxiynNws4sfENWsB6FeVusSGOpBBeX
7R5nygKbllWyMnBkB94WtbFbb/FPha/PeHjydh9+Le8bqALGuS8H/BuJS+NP
GY5f1aATospDr4/iiCp0bYR9OTaZiRdcGSBeBaAJEy0KwGlStlVaf1d0TMuB
0RbHsVtGfNKQ/Af2IHwEG6OVLOtId4e53418S4qzi4Rfa6o26/pPTk7cG94q
bz4YHB5+p+fg4CBVKelWmJhVn2nQhcUJuNCliZ2JG4D1NdlO9ZpN2WW1fyM7
28OVNQwmJ8G+rhTGv3KJsxSzeaqEw/jWpp+m6AWlR/S9UvHok24pd3wHchjp
Dc3JmPDx7VA5LU99AdPh+xj4frwXj5QbNkpS14sJVwd6cEm6PittJk2cPsxG
74u9L7uDqgXvU1MIsd4Pe3D4C/3peAaEu622fmeMqAKLlgCULyRCy9pzfHSW
Tke76BDJsxGnm/vN8jow9uAj7H+U65tnArTWcXJrxgZqFAlGF0kQfnf9dRTo
ID+pCL3Wff2wlXcCAuNlmdiQHJu8DGfBJYfUcmt3KT2csJwbtMKcbCdtQmEr
kUU/U7fp7Squb408dq1tCawA0jAclGnZ+7agEJZxVMwZ0I63x5axHOKhOAGF
j06Gc4LyeI/g7iC3ebMuk06f5/PU/HQqtU/JRGh24NVKKcFLQ341sBJ9IlBt
0NoudCFpWruP4Xn+uidPc+2yinETMOWADGUBE9kCM/wVwU/9Nj1jkNmkAmwM
rC86u68BbsMtWzzTPCHLkOI3sTwDcc6C/c27H7FN1Y3FG4/13xf2XyrBo3tF
NcJZJ9l/TvCMgupk+T6i1CfH0ueK2i+3vdoXxUgSJM8qWc9pgshq9/Sv4ApK
baQ/MKDO/1pUWYFKxk+KCep+jz1ZvzCMYYheCV1Y6wVNmHAGsX/2KsN/U1Gl
qnUbJtHK+L3eOPYeIfdNeXy40kee6J+Gue4XxMz6mlA1joWpCOiUb5Nm1PJQ
zOns/s8k61xp58FvvwEFH/L4CJNhYwbJb05dDwnKOSYaWgQL/K6v90wehOJE
nmOq0NJg6QBpEzth5CjtXhddYatTYdNoCiTBPJN77enOjeidZVVsbl67YYpY
QaPuD/j+HsWydIcHVAPuvFjUWihMchSJ24SFL9bdGIfKYAJDHHoB1veSmQ0w
4OS9mFRAUXEIHkvIwqNbB3aw2dLHtTywbpusgTyi3qVnGm5oXm7juZmL7CcQ
wknfX1ySRHVy/FGYQclTjKiXL2LZwvmX1tPguS8XUvjRL9HxLtYuo/1ZYCWE
7a0efu9aubMP1dsZT3ohPxD/jpnH2zCuw8+VrC15v7IuGd4BaakLbUYEBUOL
sbFKW1k+IpjfJGgc/9MoPE/ZPiSTVz1pPOJ1dx+833rHc08fyR11xFF50QmC
lt4M1H4/hDwoEQcuFqVp53JoouNyVxxA77Gcb75WeSh3ZnJKiQTbG7BcAcUM
sumK8xP4Ol233D63zTvXMOvpIgiMzuLDgrKDinmMfVHWphZDv40Ffob3gRYs
6z765t6CXKR9O/7gTvhMZU/pANh3qVK8GKNjfWBW6SE6n+NrC440iFPVNV2/
j7n7JOqGjWHnz15+3EEMZU96LLFGhf+B1YLmfsA+m1qNyLMXC+fiIB2GMcTf
oT+ygu7f3+BZBLv2oBT6jpXWc2a7qGHSHCa7LGTcJa50BQ6JxAYozTih+dpx
hURwQY/dKEGSXS/PIl6F76XMe2hK2e/D7mjzCgUKthE1+xVLRT2SXNmgvyTp
J3u2QYfVub+szrPKfCiraDOQjWmpik6EiYFvBPXxmkLseGOvGURwil9RvWUY
Mzj2QoXd7VYydAt2/sCLEUVBPLa9FcBcV01+sAsAdMzhEH1GFrN/EbR2ZwMi
8FRYFjwIrA6XG8c9SzPm8GlunG0cMkzgxcmEOch5NGAwoIkyfqkN7g8cPgKN
ogwuaRVD/GFTgSubMqSd/hamyFzWtV+eSa2/k44MovcZxUQEyk35smQRXfV2
XyuwaZgToOdU0dqA2ueA/yHwKzpxnlQhOWM9cRjHey6v8nDU8uEvvWjW+np/
ZjliHBmU0x1PDO+VdwJhhlbP76RH+mzcupkWlz6jxqigZO4r41g23Jv8+hJf
zs0IRL5o2uGW7XZ91wqB5NjnEnGQqKAd1Bxt6PGnYhe9rfglASOpYDE+ZH8k
b1xAYOPbGnlLvy/RVVXzTAu51+/rt/EPU1dPpe+zQOpe9/SRqnQp7eFdoZ/a
A5KX9xlLLvWguA0r59b3rTiLwVqPMvIbWPRggitETDKebcGqv+haxN2BUsRr
kr23pZIvoAMnHmcgo5MNvD/lJF7kFMuNf6FUeIKFZpmTyrsFBsFfJWlEGaO3
esDPuKPYeFiARCMXvu0DaQu6TQRu6b42uCgrcrQsaaKyjtl/2M1UiQZjtxq1
hW1seRyGbphzJm3xQQix/R4z9ZVvBBcqBiLei9fdraDmIdO6tx2oXzmD9sc7
Kx7YbIMWOBapM38x4CmtrdFZa+YX+kR/FkdC+/7pDLZ/BULsr5merKRV2ZK5
x8r2iKze7/0tmIORoLK4PXJuz6PZ1qK6p7l0aeJiSoiPjoCHYJcbNqxZU5ld
ERTHH/Nby9rLclFKZrEkp3/9wE6cz60mmCxo3cmuBt9qCjPxHisGDNznV6bP
qETMYVaaJeRsBuYAr8OrAu/xjXQiU7raJoY4+4nudYbwV0oc3zNcvNH7FeJl
YDbuU9tKj/vZwt77l/GDLywtuF2+y/dsV+6V3g5DEnHx3odyat/YTZo7tpPc
1BcUTXTHgvuDB5lByHLzE70vHD5b950lqslzxvPWrfMANVjEZidVFYNf9KZe
EUNPCCVKvsfam6EWak79Zoc/4ckHGGntfzauyXv/nUMhOum5BCpN136Ys1WA
RXJxpk5EZ5mLkxk0XfT4DsJveYNaS3ySC/1DhZiT9Z21GJhsIbS8CVooMy86
c6bgNIXw2ExLwBmVeeqDGvqG7RrBgOwLBqa3GY1XKfay8KdxzOtGZngkcPI9
ugo09k5brGmekgu5omgH79DkwVYIqNj5JWS5nLNLbC2+ePsrM2PEMiwOL6z9
z2fAQutj9mp8F4oVn8ttF8joqpXCPlWDJYblN13/n6oJGQTt3sC+hhzOWaUq
9yBgThvFcWrs6v0D2S08qwaTjlhTmFgvU7jxE0fR/KAcSFib42LMRxAs5TVl
3dfPuRZ3PoxmsNlnUa6WtMNQUtz19HPySw6Sz77guheaPEwXRSyYirnNDoRU
bD8/EhS/VO6i+kCRzPbgIZ22UpxoB+PwWHVAQRBIChYILXvd5U5JFWyriU5q
kdyUukPpq6MkabSVEXMQWO1IZop3rbLpm6Z0mnx8zqmvhPe1VeczqS/uT5n+
No3HMpm+tztCTDtjZdQ20a5Fdv1Zyx8W7YMui/rERyID134HgdrNORd5PxD3
Fi8Ja6derFUXeFszFLJ7kBGBPgtKYB6ekMdBGLCBF6aCCzODmdYNuR4cyE73
wAeR8nXYwEyNE1Ulm4cVW4ecSVVLmdcDUqFqdArK7pVMwiWZyQ0Dtptit4nk
fvtWV03nUxErVsbKzb6nNlVIPK8jh2an+BDA2tgGP5npFWtxnqSMHabMVlkU
DSGpX+hFhHNtcNAF/KPpuTY1PLOw6ruvyAMmEN8l76BkeQXrTDE9qbjbN0aU
mH0TAGbrtO2lSvbo1btHfpM0qL5GpZZ5lcydKQn9OWdEbYdWMOyAX3qATBWr
kyi6M+89BfilJyBZhynrp53tTugomHY2m671IIqudYrdLrOA3RAyfJxBijBc
Jbm+b60bxaati6in55y87d3i2KNIhIDUVNAFIsyIls0KSPwVrZzixN02ykFD
aP/ZbsguEP7ZRRUif3sh0TVp4X0XGuYl0qRQkseS25/0UeFIomLbxVz6YB89
O0/LQescM/jVJY90cEOeO0CfVLiZTuYaI5+nHjjSNNBpvQwzlsOMpnpJr8dN
RAQDunLicx+zn7kprtarlDl1aSBDQc/hyAyUygr7/aBpckoMslOkMqhCwSBH
epmErsvnH3+wBWh6SPg/C4CSCKQpqN+cIkoutmK8DA1iD8RYTOIdzB5ec3Ws
XBTHl/oToY/rNt4AYDULlqB9M/u2xf027UbEcoU3enhcxdajlP3rp9EZGh4A
PDPAOlNYlk+xbaFOgczIaOAlkRTMSWbICWTCahj+m8scQcI0duGhFSxKaK8c
DZruZfsLt6BiaTpU1T+X1Tm6H5l/m6y3iuL2W2TuTjqLrpfV5aeqyJzCL5t0
fDIV/hnUmhKM+Kg/MgVP0MhK0REZniZAF+W3FlDCahJ805RRzRn9ZL38TpiB
eY1obb4a3mCXid+JR+4HKOvFwbxnZQkukBMwmLHA1v1L45d00nw6c/4bjJQs
vFrvs5QGWXNi+huKmHVAtQi7WidX6dxnt4UcSdyqtumLFFJ5SYJ5B6yUMXyF
g3m31yIUVs8Eqtd7E4j5MfjXAoQvSLQnNWXGRZnKt9XOBOSJWzE7PEhsVWzY
44RfineC8fvjBgYO4hlCo21AZZ0l6qMM7JcJ38oFKRZzOsj3UsMFaQQHh0eW
8aA0AmCCC5eFZRfJJ841KnBMKhenlCXR1KfgRZiw2/3rJMVcGfm8Y6IsiyYq
pkf1y9hozD8/Q2kw1DQauStQBg3GbOP1E79F6phUcJVwnCQ4ay1Or/N8BCBY
M1nmbUqA80Y2sH8p99+OV+HW9XGgJeK+JYfT5BK2Eo9kaE/datyVyvI+ZX+r
0FYymsHOpfCYfuxTMrwIhaG0OHhJL28jevc0g+N1j+j8FLjX87JU6KYzs2rm
VuPbFIOyeBYYPUzNnlbCyzjmMX3ejk6Jy/qKiPN2Uw4e/JpVtX/v9mXDvBBq
P0e/zSKDIltFUTkiVXBmLxR28ItH6NHBiDYXW9UNiwgq9aNn3Szorgd181YV
MCQC4eyBb6y4M0ZlgUnrQ/ry7xWa0MKX7rNcuNAdeffgedAvOt2jNciHzmPK
PYEJpIelBkaUf71VFnLxznCjcvnJljS7tslFx+sKN+RiK7ioWJXyeiJTjlgW
Klb4N8i4Rql3hU9c6Cxx4I8g/Ng8WPnAQQpV+oGymXpSiveTQy1ZWa0w/CMg
p21pJ+xqJ2rZMldW0xr7kHs94JXyL/XYsQhy+daUeL6ib8UZ6wtOjHPXVsDS
vnsU429xDMgIiNDbC780CpQxQD0EyRVlK6AixiBJjUP9uYh2qmFkKWUCMvT9
xS39MOPYDmxXoqfK0Ja8Vp7Xh8njw1sdV3l1cV7jmoAFKXkAfvgidT0iUpIk
wQS+2iHYUSzgA3/x8ZEjb5eAjEv+zxSslonceHAIhmZijUV1N7IBSR4oOxil
Dh5bdJCmCslsOTj452WGZLi6Zp8j4wPB1N5ezba9sjDT5iByusAoUkgWdY7P
9k5Lv9G5sMprF2hL//klAvMqYNpHBRXkYfH+Kui3dktSCcvej+JJgfBQfhg7
SyUTIEhT1hYAkOPSYGvwkgNG6pOd+EaFSaiTRSXSan2zlnNLGapeU1U4aE3T
UBW7X8/RVL+KpiGsioNsR6ZGSXsD4BmWqgpvV4hATGIpeIG17cPvaUhlcdOs
m+xwToI6ch00woj7+AQcs8+ZplpL3VmJ9BKiRN415nGh1kTO7TqgHMWCHY5S
cnCn/5esNips1bK7p55PRjvVjk2LIfPcR1DWlaonSt2niDkyZ0AC+SSbNWa4
v3D1R4m1Zee+WrOKLTstGAIMTnQjrHXM2LM8Koz05pWDr6zXXBOlTfPEXolJ
2Z/NFvX8gQ7ny8qA7w0Pw12LRgcDzeeIh6I7hEv9Oqbxv2TeoZvfidv8W/0F
X4HVnA3VVMZSKeWkaKlIEFhFDzaStcmivFI5VSOoShxKNyV3ga8wjhQGiGzG
1NUUpdP5e00JpqQL9ylJfowcL2niIoKhdKTjmIxHXyp25hX5Ap7u+zjAE4i8
QS0PEXGQDnOpAXSwXmiY5QtSh5uNIRTkmDC0Kl2rDlxSQqQfVBBbPGoSkw4j
B5J5+FgqWs59rTWdei0iDQPxjgu3X+seEsT4I6Xp3bnXzfLgzDHEKtK9S0Ot
Lyd2W4whiCUTZZnyx5+oljZhURrJ4RfyarV6ZGl411yg6w9RGYsqNGnnZCRM
Pm7ryPRSVih8A7epV9CJxtsiduTceRGNbldTVwo6RdGPLXC0UVxDn5JtytFQ
o7L3l1fsEbhsmN/ERexk1zMND/mGycpXhGzthIvsB1zzgt02HSwSFDRntdcx
eIdxL1Lg8HsOZg5DAuNKYP715n5nFdYfVfST5yLhYTpPsVzWg0wIHmvgsicm
t5iUxwZvfnntYbJm6n5WBFNUVoqFFos5LxVE8PIxcFHcrli6YFe3/KF8BNyh
hM9FXHrLVtoxyHlOKp1z80HxrO5rxqTp3WpN8vix7z12NFj2UR2or3s6lA0q
48qFBrXDy/Nh8Iu9ZV/8g9bDpthrb4WZIbNIQs0B0cTA5YPAOeuj0BfvVJNQ
8HonXy0kDp0kNM+TYUvvzcPa7y0NK8P4BY8+5TxTq/CgcfwEXJIK2UXmRViY
86/btPkKaCjN3UekZ0Hmdrtkor4iR0epldrZ+61wtOSvdUulaTBUZOpABF+8
mt46Y6dcetR9HRyzQJwRFERM9hqOT41bNYKW8N4wDf3ahMTZLw/jcqJfbBGu
LE+wqDvS8Il+/cSXQy8YNh3jG1y4obnTs0wAcDBIOtURvPU6lY1iVIJjj9sE
jxtQCMVasuYtxh0aI/crD67SvPN3O4BhGxtVv1re8fbeAB3f/ddH1xQz0gnh
14xtr6jX+llE/50/fW4tnbqWhzWil9sqELlVangilU/3ZYY29IJ9YKNNAKPJ
dAvUThD7Zar7WHZp65+42CEPmo0dlZEXVnbnNJNwvl9JmjCourvN/6pfC2jd
dEMWQnmuFglnm/u34S1FxcvqUWoXyu5WGwhFfVGgHSIbKz07c/qNNdNdhs28
bDjOuu+Qfm7fMVF0MuCUpIEHGFE/NWpK9ozhZICQ3lIOhfMq8kGxzGrckkks
liB5vyP3LOk0E71QgOmv0nB/qwL4BfmH8RPmdRlpbWiOHPAqcYBM+sqleAZD
TAN879kL4s5V6hhs7fOlWkjSDrE7un8zLStjnIxW7G7DnjgoKbnk6rUf3myP
eVPjWj0UpDAQiK03AbNucc9rWMvDfLvcgYToCHSy9CzRi9GGQc2nBFDY6xn0
bG02TVeC8M6krhaTjaRT8EFeWssUojJqR7epBoAMm5SioellvV7opH/HSfRh
rVkc44pD2mLXt39kvSdLSrnqjs2x4s63rTCrtDy3Bd4kO3HeNkZtJIORYHsf
omr7QV99vkz3trodr0i6GWA/yzirL54U/QUTTiBvBgQ/bBDTC4PFRq1OuBtc
49oqcqnXQ0qQ/BLRqlQVlnypXp58aJOq5ra2C5dislZCAlvO8ndzWlXonwas
idMvKRVLnxaY/tRrtRB7F5OryXX1Cq03mxoUMvrEaguUSzd1SmkqCR44Z+5r
XNIrMjlWPGkKbi43XlN6Yme1LM0Rk4B6Hvu2j/5EDL88URTSsNWpHwcE8j5o
i29pKK41sVmuPn+FkB7Y9OIGgVqhkvdEDy6Ts6DEwmv4zhkHXb2hreBnSf2A
3sFt/h1DRxKBcvJs5Oqx4MFiNW8l+8BtLy8OJEvRhnpF+TR0/2LdAIJ59BzV
kfG4eTjv1iV0Td24+yy+7EBrfISIR2Vd/ojkx4l2mKk2KHJ4ZBh5OZAtpcLV
jAaF8Ma/JJIW/rIn34/nsvtQbW/7Q7+XsRVn8PZQa86XrhtcYGrk3k1lL4/x
vAyGeDaw2EO4RW3YEg9qenLnRTR7sli/Mjk1kJ+IxNfgZPX1UTwprnSl7nXc
Lm0c+Hhaa7f4WmHkrnyfcDfmKNVFfidwFHM2M+B79CFjXVvq3MpqCqzDIq52
391g/lPGYmQRQzBVeRdF0k8sD2deiWbOIIyEaFa92w8LWgtEh7Dey6ZQzY5R
iNCg9dt8s5WTV3kJc+Bl6uadXcVIj65CUYAIHGOvlmgD461fl5ld7b8oz3Xj
UE9pR6DRsHdSQ8NLZ1qixV6QkHKlKM0TXk+jwH5NuP15F4GITjyKJU3mqszG
YK3M+TilHWY6kyhuuxKdqpoygz3z2QiGFrJGiW17wobDERDCn89UQrAabCBy
44DVBhCLzGEJU3gsJKuToPJ16VZVPNqZFDQktvUEXayiLFaZWgnkeumfuZYU
qb+mwhscWCiIoBrDYtOgTo4aSmpyEj4hS2Ugla0k7T52cWE2jj9TFhd2WGBN
4R4ZK/2x155EYObI4wFpTb7vfRdl/bd8Fbfjmz3vI1pv/KNXmRvZBcQjq5AW
FqvNMF2Ohz1jKErBzedbvZu1uCvZppqXF+AA4Ng2r3JuqlSn21ijbFWg98HS
VnhwTrtQ7vBiwlRD6t411V7IOesEFbW7P9FF9/LiXvw/qJWyXIY/Qxn+o7jC
h41jXpXe2SiC4wXtHmez0ck/BldS6p+w4cK2d9tq+KW0laYh97q+Z0Iv654k
07Y7sYi1cHRIlU729rhjYnQpy5Hj0LdYU8MqHWhxXPSVjITXov03IkwpI/sG
stL1PY7P8WkPuKg685lKAuKyJrRUzNIN8JM31DLTKis5fU77oswSJWqTFYR7
DGFupN3G/+GaO8fD2G2erlj08/sBIRm/ThTZ5irU+05R1gMm+hiurp5mpp34
Tz4vvc2bpXxY6393BvrOlO45kZoR8OLyP+KPSXS2T9rZtnW0r+f1lNmT1rep
KNC5SZODWjBGssyqzTWx52lFb7cSG3GcmoL6+ulrCK4n51nDisuwrTv3nauO
CnWi1IFYMgupsTyqeGd5sKkyIMgG33TgG+yhn4yqr2Uf6su86kdkTw/rJ4D6
ZaoALNbJc7THymRZl9d+lVeY1M5ImlptjdbTsHpL9DKLMcF3+nPJF08OAeQ7
W23w8Ajjqb+KlwDn3NG7OHg877EhL4Ti68+ukXx44iOEFVQ3NZsSeJtEgafJ
xGkiAp/8tZcGgfMPpwHFdDQdRi10gYaH3nsdXyCR+ojrk3eQSk4ILbFIYqzA
Pw2ZZq1DGF8JRrVpd0nSdstJAH4d/f4g4DAusO8+T/3KzzlrH6XE5veLR01J
RcVDBYAefHohgZG7PYDhUtPNrhlk7HJcLQICeBwl7nhHkRCRkqWd/lFsHsoL
Vka7CPHKzOV9w5w9hm+dQgy93vfrs8RRx7TlWf1MdfBdj/xPwL/sYqr8rNPA
h4wcoM0WBOqbcCTxc+WnaEGYamYU47sXZmp/CzLSEUAy97ahCWAZy33/TCaK
jy+7faoCNiOCbKTkgAle5NovoBhwxNYIS0PYlauhv7n85OgeOXgLn8E3wXPy
y8BCG9zCA9A8REogL4bSTJImtAPA59sO2M3k0d02gdB1eaPavXRl0DXcF/Vr
xWC01zxc05cN9BnuPiXswjQgj8jfjD3GzgsPI9rPL+Ysyu4fYFN524GF5pA1
+TnuvyJ/uQIOB0CLjIhF0CGuD89i+v+AwNrh4eEsS6WI0VkNxC/OZV4hTm2t
0avV+cDv4XFzTVQTmZ8t/q4VI3I/5tlVX4UX5Y8jQhJETLcNvnTNutSgBqCg
GMlA7OVOuhXeUD0RCyDZRqgDZgHbn6SyuyWcgZ0NDsIJzOTINL/ZcRGbaXcj
XnBOMlmC3soHO4GcLiOqheblmpoiKKF1JaxOExbHb3F9A094j0XiQ+qNBfiE
6aVWgY4C710FLUHwvstAiWhhWUIVPtsdEc9NhP/AGHEX/moZGGEfjkSln595
AkEUXL8QhtPPoSPZK6yIqrW+CTH8+gZIzR6Z0zKTRfr/kocycwF/cqya0cKK
fJrgQYFudaCrY9exCj9ZgXJHK0lVBG9skNWpmkwNyjHVwZuwy019lsbZH9QI
MGLZ7lHUAe9Hr1c8ZO9qmSuszG9cEudzNdizBGEk4Er55CspeBsQdYqKQ/Z/
Zvm6YseAv1nO1ForrwbT1EQ2TRd0C1oGkcs4HAINytslB4w3OVswkOQGuRiO
2RcJ5FH+aseRMjYAIwfOe3nxFa9NKQ7nztasSC3IgosUWCzpkrtBMlfc1E/O
0Qo1oE3axXlGwl8oDUxC1STUzlNWq6EL/uP7N48OEgQNHOTEWMhobI+QbYig
jUlMqYffRo+bvfVUxUCLbZK+HbALp8C9hq+yrrWmFYSGSZ1hhFGzVh4w7+oq
LY2WyU3GrTmx3ccu069ALeVOLF0lvAIumoBuFmC0hdiMm9tOEAJbjuRpEia2
q8w9Mp4kQsmDMADgUZq+FMm0/cGNIOxvxvsSRmXmmDphCloxxcEzQuH3d5rg
vpk6TVDejwXGerDy96W31jDexKhMnVb2gNKFWewCNY3Dk6WihD7VJIFkmfhM
a8yDIlnThlm2Z07lDUOYb7FPc8cteZzKv+6bB07fi8qAiNm33RPgvyKJLotJ
zemQ9YTX5ekjQL9wHi/6FysfBWXxyqmE4Em9QXyM204O9VbiRvbIka4n0rpA
4saHB4dO+8EiGTZtOBW3GKV6pKD3KGgCwGZmNQkZAH0cLqmN2N6aS3ynnF2B
JpRBwSh/zNP7OTCHceFfJqk/mcfl6GZWh00/NCY/3xnMh+/x3CXpr6p3ZTxd
NuqeODnPj06aIVhoRIqtiU08SsTQbXL/1nEYYw+fKUCDcrar2xWZuu0MyFnO
ssCHs74nggKTsb+yoDX2+b9NvX4dcTLKAmVEgHwbc4AqmQ/e2OS55bNMRN70
p9c4yFXAqEHb1k4mhZYhW3UHSFThapr8dRzEFa8FtZC41LFKWeizywgnV2z1
qOOF+CFFc6demBhU00dscfuEWyBoKDsxVSc9c5YYrH2c1RIUXTGJ2bLG98CM
jNsHnBhbaWEDMBfqGpDuwpyvDQRT6zLjXXy8UBVJ8XqKZEG4UdvejjSL3+jE
zCeKRmkxMRQXrwFMnxtfImSptjx/ksQgMhaBVJTgb2QVNnLeWZ/C8rQxL657
UScwXIhNOFSYxsY0ifOpcaM0SvLr/JAm8BfCJqzINbb3YtBxP43U0JK8kapH
S9/fy9cu52DDoaGMS+HiqWlTM5QAa9x+tUfVz+fwgDtF73y11Mu792319Yes
vuggenfjNXqjECF3+ajSE1XZqWsQv9xqSEY97Zny+Zimu0UF0Mw/Jw3Moza9
N1peNlveGJn+qde/IMybapQlrmdN2HFLw43gHTQy9nTcKZ5qjTUsS0fbnQG1
eK5rLd4DA4zNPO/qjMhiZll9xc1J+NYeddUuez4vKoCbVjBeu4/worcPrBYh
yNVIZt7tooq4Gc8jWPTgivddhhvLpoAnDVPZFZXN2qnuL78f4ljsx2TBwXBW
s6RUjvyOjAQtdA75Dz53wpRrCHyx/DoJ1+SyAgF3mphP34eYGs9JUaqaCldN
Xz09h1ZdkWuH2yKXrh05j43zD9elm+X2i2rAPxqkVgSV7Gn0LAE0uGglnHD7
h0ZmlS3CGO5hurMXBdQ6niVNBzyokFEHzVX4ItBFzqicG5aVC9j3XxR8G7kL
Orofnd2ZXgketQspfJMejh0z2DuumgDSRZQv9S9jpRyileWYw+AJPJlShgUJ
Eow/vuD3ziA5o/g00cDJCxO9G2HSxU23Fn81mW94uOOTd4Cr17PH/dpvgDzD
Ob6S5UZUOpJ7TDAbboQ21UHRX+VxQKXeX8sJgKeCSXvCSBRkomsV7ORNppM/
aPIjKjjM1wOogALzushEah39k7tx8vB9sli9HrWUjKB8HZ40OxbMxCQOvbTR
esP3/Qutt4KVOXGu9UgtgrPVMxfwO+htdLzRp7B3mPNeTTux2oFXpjcG4nhT
zElOHf8rLPgbimNXF2oKdQ6yLAXAuBy/LJF49Ps6OL2FkhetiOrgY0hzJn7f
bXHWTXp1LEGE5QiAaqFw/ei7hz32nUpVrWKct2S3BpNH3gHenAWqDwgbGxhT
5uqey/JCToxNR/1t40D0EZjZchie7nupm9i0tumfpoNedfRQT+j1Vkw1Bm8/
1ZTTzfNyF7tVuR1ZFDjTrmDn8ogtWvoN4BGvL4dUrFQEquSECYrpowHysCcv
K0cZegpkjCipm0NP2zp+2n8G8tc+O02Yfp83ZzgZKI2v7viqZpMLO4rJPe42
lVy+kaH66dX6rQzBn6tvLzHkwNpKYNd7r4IrvCMORu/MLKuFRDhQtP3tEEbR
N4hoqUKdcc8PQ6skp5E0iLuqUCus8Xu6aLhCw7wUerCSf9GpmVlY8RUfd5d5
tdL9d98O5pHlMB2LEoGHfpL4u4z6bDJugNho2mdfSZS1ciXJBeiB6nhJibD5
y8jcUkFmxRavu01xcJOqlwge7u/jaHcW0/3n5JucHux/0o8o6ksfa5vZwT1f
FQFhS5cWKqOlqRYEVYX5ity4zVofdeJoYFIyl8iB8QGEArurrECRZ8Y56MqI
adEUm8YfvxgG1pqJPrN5U0rQU0WEPa4QDu2EQ5Gs2sklc1l8gOJI3T5JbTjx
U2Q6L5p8D4HlbhXLPbHSyy36bipshWxJp40kog9GL0eRifxbEZn7m5MlJpOx
UD7fibbonFaB/8d7bW/tgIYYwIsFPUUlnTcFTgAnJe5Ts1njEkMdA9RloDKB
cBmANGRm7h4DT9B9c0j3eZ+ADYPxW96AcGzRPhbrP9HLxlBXQRFAIZETDZeG
u2+N8aQtzijBBFbtbngJdDzL1c4xHqLXE0hcRuQroXUaw+n4XoMETBTIJB5N
fxOXd8N0yJxjmSsOMrA81te+xZzO1BxDTfhc+vvigcUUsPUVQL231SFp52tG
smxDptIM3FTJ4//4ZZFQpl1WlQ+cEBSoLH9zFcpqkSkxuDuvs7RheVgRAeea
FcYtJzQribfP756dt2NcUE0hOOJgUGX9KuvrHkeKXqYv0MXw0tlmCmngr9Xy
0rBBItAbYPXkBVYbMSJduqty1iHCAoUcxrRFa+SaybNfI09Hsllb/Oza4RQF
EN3URObnGESZsOTwInQkS/HwbvEVQEGt2ADG2yvEvdXwBpE83M1Wei/SsRip
E482923jc1aC2Nw0RlaRAW/Wjw1y5cuuHb2ASTJgHAr42c3fjvLdQXR8+ppL
QDwPHgPcK1BhImmMCEN3RhOOscAEsiu54SlFUOcG6meNTLLD1cTfWWsWcqZy
S3Zr9u6+qmXDQ9bN62DvoCybk+aiUheKnT4SZMISg3nCaAO/hlSro+HL7CGJ
kR3Yl1TS9XlzTrmeMbaIpeMb7Nx9DvJeakrVsePYoNIkwZg6kdQw8hMRpggC
aGDEN+0WWHvKNQI9n5Z8t4PfpLi/xrF0hlaNPGTzvlXlwLT3Cq2tMbaswWuE
ja2ot0PkJJqeVcWMB/zT1sGFgNldeVfHD94pvzEjFihu6QfDBlS64Og1Wi6X
pORAWlUfWin89SujySIn88nKewzbj9TKSyXWhVzMXQDYuzH+N+RpXLoMs+2x
yGl/x6d4829wvd7i9HAUukK7EqN20/Nqt1rOfgCZ45kwefq4ltydJuBJZ0E2
J24yBllC0FU2exz8g9txvlpMmrbnJVlRLoIc+iZ69RkViMXzHg1QgMxULjyC
rWLi0BXuFJMMf3LBYEKgFGIGtSxqsg2vNOU52A8b0MUro912ab45sdAfF0Z2
ScnO7WEU8IfAbJK8oVuMuiOB7TStfjAINCSFxew9XDWXFlDM2THI/soBZx8v
Msm3LGCzwR9YeEaZUI7+kBWAmLq/Uj7gbbX6MV3zG/+nP+NTycec5XzIl5ce
kl0AO/kS5lr0D4Z7ohEjN4a1WbY/lqwkSfC+YlmG24sIb07If91wenidN5zM
2eLVjMl/mn18GIUbbQsoQOatvaWulKixL1Ee8lAEGFayM4NlvHha31Of25Eg
2EqLjyRSiw0INpCepLCNtRR+avHvRLoxyS+OOG+5yIUflhOjXAzLvwRFZ+7i
QK6xWj1T9L93Qk9X6AxV4BJSUzI5unPiU9LsfH/mBFdQG5Uws5Y1sj3SufZu
VmI/IaQ5PQp8cxeb5PjZ6arbzA7J+MqmQJm1mXKXaKVpE7ky1fv4+uUD0MSA
C844ePQfac84pgZVstAEKfv13rRHjec7MaJmKjBQjy5j/MvXkmD1KxRZwx51
7GPecCkcg1vm8jEBt1IcbdGdx0au9krmS4YtgB7EPED+NQyvMdQqEUke/R9+
F1uzxh15AWFPoVRzGBPAbCK6/Nt8wRk9yH6buLuQsnJpfnO3Xlhp800Pmpi3
4SkkVgW2gK+OboH+wZX0c+dEtRhJ/Pb9ZCsoNcokc9yMwsHWYd9WDahCt1hg
ThUUcWyTRbfo2GhEAk5s7IT7gQv8+77QrueyZAfKosQ1V+m3ShXxzOqr/YLK
lE4znDYk3yxwK1SqvfSK/uU0ParxfrTtKuT3RKD+HFeEyny5xup8Ai9FU489
huHqCzLn3hGuMiYtqgaVaAY7tNTDE2tiBjvJEAjMX7kJPPScRPCRKvKJrhCQ
tFBJmNE1EZ8oe6OXqYXpf3g4qLD6DfF5UxXqm0BJ2Fcp7GxvlctbBS/2KlaP
f0QjnPtjA/NPFJ9sIOkfi3ofkjRn+a8NKneaL+tMOmsDQ/ytk4++2KhRDHAH
yFeQZM/B8x1a20WVdTMCYQJq1qDXbeJL2TKjteOoHZKJc6hSskqJ2Mtn6byd
Oo0y2Yjz4AaybjEk2JTCqgI8IHUheMcpdHBcD5bdsSGdn2cLXbm5dyZT+cEH
Ygzs/Dl0me5cywcFaqeN7uUng9FbcLFWX+K5/dS2Z2pFI5sRXy69wVn3r0v9
ZG8XTkXna/jvMsNEzhrl6SOQXHBFbfdeV450CuDgLKXh7+nkUArOaNgfvwLe
+MGCjRGUMGqYQR2G35g3Fo6zlHbaJNxEjD3Hr3VIN9iL44GQ0fDqZuItjkAK
YR1mHFi77imxQ4+4KZPPihZoBPTI1wR21600bKBlolX+6yTVe0ZtUQx9f3JY
R8Y6WDQh3Z8AzEtpw4iU/8tnoemA15Umk30/O7GrLIaJSeLWuzIeUGCfc4OF
NBBqKw9eF6LLl+FNWqiw/HnmfhFaepIxD4y5bxpitZKK6r20qq34itFBkPL0
7Bk/7O+AYGEr1YxFEi8rTyEf/QDJom7tjFIQj2a8sEWwkOYoT3wa04WjqjUD
HViiLymO2/1DAbBU0y8m7tiuZU1Movvt3Gy7K9igb3tqjXqJXDpX2yZXjyLi
KUSGc7CcUfIuwksesTyBs2C4Fx0WCl/SfFyxan0yh/P7GxAR7bCjf4lWqmDn
VHLBes1pQAwL4kmilKALdMYkF97Wpn16N1S99Po5LsVuui9QvFsWuRyIaI+w
AMfaf0ZZsGTg0iG5gsjjscSC/7vy75uieR60QQHEhto+PmUJCuj6wK9MBse7
k8aAUu66+2CqxaBhU8Q66+gmBH5MxV7ci4THn0TOpJX3jRsBdCaO/HNvMuiZ
oVcybE9cdYa/18URDT49nrLFCCYdE6UMMw12FOuYfs06j5Bcj9UwzlJ+PFDP
rKGJrVI5OnLB3HBnsrbCcNz33wB1UtwiNfBgQubDjK0WzghBGFxXkICmtLMM
zv9hhlI8hn7WPbscxlW/xeKUvlutfhoyTio95lkJGcmfeCvyhMLTYcOMGCvX
39kMemT3H46WgYS5+K2QsLBf9IoGSvUDkr2pvX7Y+bQnXScXF0NmtPqv1fNF
Jysit13eGpzG0Asn5KRRuK2blegWIsZCOE+Y9qtmnAZftJp7lIX/lmHUtl2K
c394aapyhDhUtGHoFRjb34HyXJENkqtZ1rtDaSfiEkzKtWVI1+5oy0y/vfEB
rDt6FqygnH/G7tuytpTPgGSfZ+OLcoIIKszalKWp4b4JcLT+iLxoi9rIC5U9
TESpfTdZhkhJ8r/+hPg0UKNB58GtMqbLXxC0KAF8dfhtYQHD+A8+WF9h5bs+
8hQjji/pZkd0CY7X6tP/ReiOoBaO53tTDpOyQBLiRwSC+lAJiTo/LyseGcbU
iij4LFI5QWVyjwzTPmCIB2P9re91sBA0rWYTwaMmJf0so4TI/N5idbTApOt+
5cZhH4KonW4Di42mq7MAfKz43u5Y6alI99W+EabHwjwHqWn/jdvS1bIoSCkh
J2fevjvuppUsAIwkO4slK0HYnfUcup0BT5tqHipJjHoH6wiHkqiftIrYkSxP
ac1zxgS9R1t1ICcceDEOSRqlTLd5fIP36CUf1I/R2vuFEolbO7sK8FTif+iI
b/73DJsfnEISqOlBY1QY6NvYxIRV3fCjNw3JssksOj8Tid+LmK8WXU6ZB+MK
86PJ5rp/KO9S5eht51Bb7j7pK/R7xzY6dQfg/wuz8xUjEJYz6ceiG2hlOyDM
OSHMwC6FBbWyjqJ5mJXyiY7FTFCN08dU5e4tTns4t6wNTq6RgOn22vKoNYDr
kHSEk4hO8+bFRm9/4GkG6kzk7B33LgVLystH1RwXulA7LnVmIt4lWWoKriGs
TnuB1Ip1PcbWDiZQk60Oa8upXeK9V3eloOGPLlOYasqQ+qj3G7rGYk03W4q9
NhQDe2iY4vrZXWq+s8hMcwSxZI/4DqEk4dbvUYQlmZiak8+v8MBNo1BflY/g
a/B46TaYbImv7ZXKkVDRZVJ9+RIWZlBhX6dPoY3595NprL11evG1AkDMGVBf
VVUyLV+vZ2qykqauKakrk+pPDZBSJqaq57jTLmCWdNkoGnpAwAuVWMIie9gA
g6ZujroL519wQ7lkl77OHV9aqZuGr4Q4czkR9lmJGKIqtPMIhN3O+kqVRBK/
akEYRTz06oJPdK16tkE5QkR2Ea8vf+tDwv0JbNzEZR6wTgZ45REyWWZr/vXF
C3Y9s3sgttsPvB5/A01LYvmCxBVcQN3RS1JN0QIGTHTYT4/943LeV/Kcu2iC
zYOkDYQrDkOtrHCnCs0Y0uHu77X6YfwaDzBrsrG15y3BVXpmEr2AaISb9g6J
lRHEHs7pYsfY/xiD05Ij15dQo0t2vqo+bGziGc/eGjj9Sn8e7hY79Zr+F+Em
lUfcxC33fe9aMJZ/LH/xdrFK5X2GWWPlysjflRvwub3TkWbPQMJTdqc2sDTR
29ekjCRs+mfDAhpOyU6yCoOQFyBMWyuE8Q0a2Wg3KAip1UeXhZul15BVMRKd
DbqlHr9kVK3zwEsRBy5tSjuoek61o8gkDkbzIHSGWf94YR0yIEqBZj1ijDdI
fCq0fTAkGAZ1MqzC7t33OQBSj9hmI8U4meo/DoN1Nw5jQIO+sHlASvnWusFI
fM1viFVYV90w5UATifU3fwpHtaAgOPUBYxLMjfflg4CNIDOxaXiC6mxpsQHW
FhG5+DDkySnTe0A0zhHCmbDKuqbn9YPLOuym1CVZgrqD07E7MBnGXw0KZJh9
BdWvvx/LBDUkB+gAY0Rro1eBFH8VKfVN09LZTc/rDnefQAWgmrDAH+MHDHR9
3inmBAeFsJz1sPYoG3yJKfQl8oX3uaBJjIyaPTqNrG9w4UwCD5iLasjgv5Ur
fXk+sILJF+2YrAKMOKcg5kGO10NT31xq6ANYJsCFe8QcqWw6fgd1uDcSHiI6
gCoiqtNBb9+JjIaF0PMYuW87HXyR8UL81YHd2oDa744VfuERaMXdx9nIFDz1
8x+7w3gyrkammerLx3DIL8ZM6gibJCBVi+D1jPCtKGDa0l0+xNitjoPJYlG1
ZdkwQhFKNgef0QK5Q8c8Xm0tz/P0zY+rmqY0isXDtZJxemqSvl8nSk2zdL5g
QUmpJ0wQjAL21XXbEFEXnCGQ7pBJue1OjZBQZJb3EzK7FV2IUThml1LZGwau
br2ZzT8Spqwpvolm4hl7pUstSuPLtDomXAJo4azaqSYfwCqpPAtR4wbv6Aiy
9ruFkwH08dUQ9ja/WZ94faNVeLuB5VYMPloutJKNcq85kPS4GTtOCXMGrE3p
7tQUQKom3SyxfLEJ/amfLsYfWKb9aZ8VzdrPNisseRHxap5w3NmwBXPIjW10
5+Wdge04BJBrm3KpIDyLcU6dFIbFPbeLvcIc05Cph6GfjtCfHVIsZYe6BuVV
vtHnWvLGny/U0n3r8NZElvfZVDB4pH7lamcM1MkAB7Tr5kjD/T0My3UWZBE3
icFkf2DI646arf2xk7g1yI9atyxURWLLjQwvG74P/0e8kNT8AxjeIXwE7o7o
zI2BZkCXlLdwHVKQfp5suefE5nwEsH5ht08kilxZqflyU4iGz2UDSoGhc2Sc
yZ1N6q6jfM7VOQaYE3V3yJgeCmbadZv6sTbbDKfmSuX4FZlhvtOYhZ3IKykw
u6sXeTppcZOWFaTATnQFXCv08Br0+VbzlAHq7ESHOvV7ElP4keG6Wzg3rp91
8Mjy+qSeIHXs+hf2OQJFpk91/+amZVVXCmhPbd+qt+8l/GOjJgaDlV8asyuu
PvXJl0euFZ/0AewCB4eCfRByfkReyl1XxoSxRqlkVG3PRzaHE4alrg7CfkoN
XMBnnvN3ovq8BdfmQRwIw2H/N31AQsM+Pf41jkcfskLnOzz13zj7M3GfgybW
/yYRqWdsBvdxm4xFiA/Lc3/BbjZ9muCETv+NdOxFFu28vBxv42xGK54HAoDp
blA9rZv5mJnRqdHWegfDu75c0ZdHdlhZ4YuumoGkRyQnuTcYKOrV5eIsh8Je
GLy2WzwEHJPtBfNmPjvFVotfMbhpBKl+RH6pRyxDbqjq3IvPiL1kqNAlsA1H
kQrUhIYzRmoP1JEDyhjiBgIe1RWdNr0fGGZ7B6GjfEZQhxCA3uet4DAztKTS
dRiFLgp53MS85R4HHze82mn2N/ItWfGXlNhhormb0D4r5aaSUfgIzhMIJnhe
X5dnlX87Q59CRNnBniAoOCV/TlZ31mYUFX9OjDFMPY3N6pPIXXEhyUvo31Y8
pCEaHx1+CIecc3PTi4jGymyC4otjDsyIQVpVvCJpANB2Jr1Sn/3E+fg8gNEe
NRQsDhTOiELRwmYnSOSBqlUcjQC3qMRt5DxUFPi4jUMdHqBRZiose6puvAHO
SwFjA/F+Egc732Spfnh28ujfXp4+p7u10bqxflxHVMmceedlt82va0VqQ0pc
t9IDFl5Iy5ScVb4mZzJEfhyBhdD1TMATEzS2FfH3YP9vKRFhsLu+Y8yk3Z2d
WJ0Du7eji3WDLXrnI+HsFHmRLVEyfcU5J24+o9RS1Ny8Ucp1IGb10hclcqDO
jyZqCFNchu73pdUHCOMGA4C663D9rLx0xJequSyUyG7oHjnINtVWRY/laiZH
d7jANzf6zjQc0B/xwYpGUJyefK6bemB6cWfnI+msuuinaBRQu0GPlm1YmOcb
7V6pldViY+10uHx4ZJkNWSpV6PnGvoIUcJOtKn2oCbnqCkLr+gxdankXRul3
EzTL1kWZl4H+gsn8kBwuabjiViU2Taa+py2yOLV0Z4d28yqz5gx0wQX6HNUF
pnl4TUcrE4pGtY8HJm2rrvHfFJCQnhOanv0BIZ4vDdry2QjwRZGJLSjudJAB
ppxCHMi20vPFTQDBz+Jx9NKYqp7A4IgXo3Gaa4AY9gtaIAdebA0kSkVU8USL
Txd+kfii/ljGkiaoM7FCffx50r+6r8AgFBHIFbKCiIdMbXDI4xvzxXlLtG9E
Gmj9sFRRTf2008WcS2nzAJsKPkmLjlM1oUbD6cRCctOi6gZ0NRsFEgI364CM
8r6RWtHpBeWZkvJqOMtSeBfEOtoiPkD6oEgk327hRMupoExiOCjS/2MIJYcJ
cxt+c04P2RDtFYzHipq51UormL7N0M1lcyzPjn4lvqANNZkOKY5flH0iaMZS
i1OakJNz/aSVs8CaDw6CiOC67K5KOBWoHtOaP9GDNQlaQZRDqx8tVMG4WkpR
3hmFikIVrKxKQmhPQCPrF6DddaX1r39zJ24x14rpUJS0B/gks5a3NRlSjMuu
UkIVmmm0x0PZdjYAlUI5hmxBLs0pBJ7YArdBaYxCrBhd5spY53pi8k2eO2QS
9AxeRP4jotm0+INjv1uxO6krKvJ/f2Y1TdV7bQPpmWs/QKm43s6EI6OLOO3H
IsGwKBH5rDaOTL1vtIHiG9516uYxPjiPolGYWpAtm4TQs5A3JC5cutlKpc2s
LWF8pL2VAIaVWEJnnq2XrZ6Xpd8Ze6Bj2bGZYraAJeccN8aq0W4onRvwt8zY
/kd+jxX/S5eJZbloQsifB+kFbXZjCUfmiaJvTF6hcyXjQNDfwIyyUyeV/dQM
PNnoDSUSX2Rnnm0LuHPtolQXDXBO96qRZTks0ytx92gSWWWHWmT4irwuN9k+
BFUotgud9FQUZ/Kx4WIH7pCpzuAVlnCpGNTqYblleQdkyvlnxmPk2+9Ooo/Z
yaGj2ZlGQLFdgvLYvizW9S9cGlLVY+l77edJY+JHIxbXHxBHrqx3uIiaVBST
qEHXyzQEJESxBFLbwxX+5R8ypEf57IlIrylILKsCnBKDVfAM8Z8BcJhWtg4I
QEBMGcD0iOgfAzu/52CRcUVE89+fU51i2TmllDyuKAqdnGCZUSo9dh4wnBal
FNnqZomb72HTIwx6GuAoiP9eAoc6mQStlTD4D4TMHmXX4H2PhbhuxNkGVMSP
nPz6QYNGBz1hChhiNZTDGSxjPAKhHuPr1sgh/fNx7bnUK1dzVZbDQR90y59I
7GlXo/Wb1ZL9iscIStaIMax/bpt2NWiYKPmqPQEYD/Ms/h+enY4HWjTZxBDZ
D+CAunaYZCJvqmPBOqwQK2UoPeLDFee9of/40GyfAZrXcSsW7LONIQanfNnK
kCnRetpVMCqAR6RHpQaQF0xyvGH0AuRbOPeXQbNRF+K3YQXgtOaISyvjgW+L
qp/3LhmuDDX7iGobnDjCfhiYYDE1ZtRd8+SJ4SynMO+mRRIAzOLIg92pqBv5
IMiLbE0bnR/QTaJ9ns+aSNfrlexKKfbSCCFPDH6vr9G3cjcv0meUngWjEz5r
vdv4YCuzn1PFVY25jVw003rbEujRxtuuUK9sTXOV2F4VNNF8I8QFO42Ij9Pa
DvTHj/A4ZChL3c+lD7vMiI1QFB8op4gw8WQatGrvHtJ8hlD+IqHXfhvFJp4U
EDzDvshLJ941Sr4mnq9c3GvK4lVpbvAA0eF35KbExA2Yxm0MyPQ8yGzLw41y
60u3jLGjw7k2f4YJkTc8eFCchS5XF2o326DsgG64TuxzGSW1JFX5pQDrhNT3
x9dPwyIMfhsHMOFm9PGHtlwjFZxIXRLmiWtKqeOELRqVe2uenl3lLdvb53hS
/PCkVhngX2fWPjNXsdI13akWvID6zrjcKVTTUa2NyZE50oOr/zYygTh6vsoK
CdQhM/5xvUYLSHaS/sIEzMX7qubsXYFaYSVXshrUS7ESdOqrcJExVlPGgnhr
9b4JIBxooHpEKMgDUs5SyXSB0j9q2x/Rlsq5PqCx4tCWNEcU0D6GB1pVHBSq
Hmmj64VxPd3fMq1YfVbTGkiuf0jzTwub9AzETVT9jjhk5EHn7TpbwNznDpdG
rlPUdKjHnJZjlTm5UgZwIWSf+A7XOZHZbBncAlhSTwBkMim1LZ7YfgozyPNN
1+kBYhWzVygOR1IdUeX2myQfs+8PWv9VA4+i4AJFFHEglJtFGeumVmmHsBOW
PBdPcIledGxpup2S8/JjZvmM1JQibDJcjflUQXIsHQbqy2V1K1hLbFGYZopp
dau4aswhostnuEtOqFAx/zcphcn6y8m34wkXpMwoVPTeH8+W4lFbAPJByS5h
+8YVrEE3bN+ThugcYP+PlV+5Ww5Agk9pMx05IBaX6PFRyUoaPKPk/7fVnyci
Js+9xnTOPoErxzduDG8MsFMCpJu76SPCk5jwet4kZYH5Gh2IhU7RryAtKZb2
nkB53YDb3eNVd/g2YmJbxrDVzgE50DWtP1UX5ASP8x/Nfmu/Nh0I+By0Qp4l
ZixEst+zvKslBKmyIttS7hPCGPv2ScniQlfT4DnRHL6pyo1fbUvVSJteA1M+
qbeAfZok8RHeTowI2109IKzjlxaXDr7ctW3qUa4w9ch8aVm2vwn/J8aB7LPB
jS92Nff5cu1SniSnWwt7QyaflfKo23VwGDDkCozOsypmT4fnOL8N8mGx7i+o
9iG67MNKjzb/a1goYXaPEh3cOM5yX0FTuiERk/jz6u+ooF7aNXS4f15biDix
9XnJItQCX5Lko0JFcNJwcUDVU/2QaE0Xu0Ugrgxm4tiUvr/IMd2ICj/rjBwN
p6YO5MxZ6Ro3WV0HvuUTQaQz9F30qxkomuLnODz0gdySKzitva4HVq+ok1P7
w1eRfu64pPeZ2zIRPW7jBQi7qMpA5ffL6coFQmWuFHrhpU9EQ0VI97F4dG5j
HkQGJ0moIPrE3Ex+JeVo90GQTS1zJhGD8z1i1/wZLIds7xxnUnkMi7HD1Wq8
s9UTnh8oskeg+qh4nlV6DogK4JQi16W0+wIRipf9EmcNK23LmlAdViTEGVTd
igFgmnSLc/9leVgq2RSIFsLoQygV7/GTp4tlVl9t13U+nMQPjmkdU5TBYGdg
Cyh7/K4J0aIO3YbPGlydcwdjuHU5lzXHf8EVoDSPCnMqzs1sDYov0W5cMxri
XA0yhMHDDDp7YcOjfRVIOl4GxkcEAoSEtK5QL1i9s+1e47uKHN4E4LCUjLdY
SENQZFpw0rLnZgF/rBE2p473y3Cd5bOC+uJgqfCgVf3USua/IusmMQJXnXkF
SYW8rEvhh9zzzn7xcZi8tSns59td+Zr9eyRiqqRpeQlaTLrEy/UwQDLThiWo
ZQOTFw6wHU7VL0T9ygXIfb4x/7M9CqqOrB6mwZMDrCRfV27A322ilAhPXFXc
32YF9crHD3nuH28Etd59MW3lSfakCub913t7IzYYXQwi/r8XyCtUGeCxIEb2
npYVmTvMXmBHyihGNYLDw7vR5KS4aYEai7LGwZphjPgZtb2Q0t72koUoFOoh
gJwZkd7JfyKYUhrCZebzWkSWh0KWWRy7gnGf0qK0yfCuj7rcSL/xftW8H2IZ
PIrfX68RA1srSL3PJAiMGwkCP3AqE1My580gG2gyzTXMCR/HQVzlT6diIMS3
GkunMvfzO0wPboSTA/ltAuSQeVbOfW7/x3C8h1SlNcAh4OPqFv8vldg85SC5
DfumKtFC7NxeSnDpvoTtJ5lX87lyiqiDMxby14HsyzJRqVdWoo1hHdTBYX9o
cjgTy0ZvHAt/Vc5ZgQ6RbMMiVqiryg9dqEk+DJaQwDqnv3rdHX5jDlRp2v0G
y/of7DIPq9GJvrvafBmBe/qSIf2AiWOfMnoX/lqNpOS+d+YEKiu1nk7M/XvG
a64Mc19fx8pfH9eIpDTvduoaryQhuYKtcZFXek986w4TPTUEsVVfTyqT8agB
Lw+ogQWyKHZ4lofIifCb1bYKROvN1qkvHikHw+bvBlkPa8W/z5EiizhtGgRr
JwOQqeIYDIAe6Uvii5Vgmu9f1zKgNcifP/pPfZQ3S/mDStJ+Ex310RIi3j8r
lwQvhZtV9Ismw5gMl/n0bxsQL2EYSMss3dSpvbkrM+X9DIbglDJwxSnu0Rvr
gTPoQGuKGLIwBmXmoPPqCfpnVZh0e4ZxVqR3DOH/vdFXVJpeLss8sse2zedH
ceaSnjhKo+CXecWKvpv8KLAoVeYBj1I/TSyIBNnP4rUzwc3stbmc9tSZvOA8
IHCIC8LsTVY3dVcSALmlByfiDBCE3dyRgMyXDu/yc0bT78iuwYy4aV95U2Di
Yklk5RT4trgXvEjbSpJQkT5BmQeOlxJADrpsreKMWJU5fMkBFb1itDYx7RFO
8snM8hRvBAfPsEI8pX1wD5YnytngLAJFMP3y4ZVNaHOEidXvg/zv4tdIPnyD
F2cQysBIEc/HKmM5/7Ce3cl+fnc1O/G62X5EWabe8jmCFFTVZzskXf53V8zm
4WKiDAAoRxIr19MwucnLiooj6EtBGN4jwrHzLsI4S1FeGIktVBavDST3HU7O
XQTzznXq0yoGxwEKwpwaSkJMeUKthNpUQd2Ltap0yGZJSeIxRNU9gfiyLqWQ
1od4XRqUxOOtzUE8IfWhbV3JN5aBQJC6pQX4wmuUKA6a0i/KpEcZejuJBVYw
dDwVUt3j8b4CuA7V3U+S8JG+1rQkbLeY89+1xTCW+wcioIXSVlRqwn1Tp81c
rwvHnftw5vPgVhDvb+tPoXTtVIMUomafs7SP+fbuCzTPbuCKwXqKfofVsY/N
GDJAPBwByO2I/EQNIniqnsUx86M/p8YIbwF0Pu+C486joghmRiEcdQfRY4BV
S2xj/Uy1wbrMSION+G4vw2hhy/TrLpeHAMgllvFxHZ3A5vvGJ2FY7Y3vlQUS
kXW/fcmylHz2RWk3o+pdwwpZYTaTyfekQwV7XaMtAJK9lrB2VAym6nZ0ZcDJ
BV9nNhqUQ2+em8IGKxF3zW5UHKIqmek1VpPWWQb7gr9MAxRAc+0h5hRtffXt
NxdLGbwAqmuruA9xzSZfULFevsdln1He7GJQ4tXSizITvwJGZjc89bvc7Lqc
yhnaFXm+OM5hYGOVqD3OelREOfb0PodUJ+0OMFgutBnN1q2O32RaY2D/dThE
bcTfnKPCowF9PwgrI/FldR2Qw+G4a5Y5/jw77yMAa4AVbAu2DDGCiPrkO3x6
yDn26hDySgjqiMQ9offSB/xhlrjzo5gcrqkcmwX8O9N/QpHKbEW0I5ji2wRP
kO+mYKsTJp4VfjkzUWmnm3180XknmSu0YMuwhUX2FKNEPgGb5C3iFS07Gr3h
YSKotPahxj+2/LltZbud/yhOOQEP0Q0ezdleVMymI06Kq67ud/dUnHlx7xdr
gTP+0Uips+zMEkPa//hJE9U9i/yVTlu15rdRu5oAJoiByG+wsG2jwyep/UO4
sLIsEi+c+ESQUXxbyi8RLGNkgmwAHxBfuXmO3amObZv2yeHK9eOABBQGgVEZ
jIgLAA90wsdGz17LBt7FpAwIVnzfKqfqqkxm1hK2cWgIAmjXLWKrl9eqCvDl
ESCoVyU+yzQ1QbqPy9XxUMjUyK4GuLXFAYKSAVUYYYLfYHzbO9o23O3g729n
gbYMhOOI1dCgw8MS1NV5tjsWQhEblly7hCcLJzZiRFSD2OsBVngAmgW2o+Gv
VPPJ2tolFOLIVN6tlMdK+yXQfDijnMoo/tEgkgTA9sxCT0QI0jtYohQzwwzb
U+rJqIBqnijy4186812STXh1MGrP5qnCQCGcb8zGphFJyKXR1Ql0pCOMlzq1
OkidyHZL8BYuQxOXGjvO+SIusE4QxD43TKC41pcPEWokspYFdmEsk11SEFHK
VS3Vq0qFpME/O1CQsLOy00P1onY8Oz+pe9L3qJ6/13E9l/lkpOgAZ0GhfUnb
A/BN8u7NhL6BOFIC6cJEQDDu5iravEmyCUcsEpY6O/zZ2niDSj0gkLcSIaDv
uQfCfO9pjrg2XLChn4+O8/8fcjMDeqk8iBRFPXPEjIEg6ajaYwJzxxPhJVg7
Iu4pS3AykVC1f+0+vzM7FzvxvcpiCZATunyS6y1jV9j1CLLUdBZdvORiJTDW
TnuMn1diLUWutsGL6aQ6nw4uRxn/5QTH86NRCmowfe+wBwN9UOSr56H+ps33
o29Z0s7W41p3RJivAafy0gQZhR7u/Z9qEVINDv2z7TqwwgmKp4yG3qu28JLA
uTrVG0N5tTdIvxX7OrReY8jQwIq7+ZwL6PIyNsoLxwiZC7lRzC9aCccBRCfe
b9x3kZqPyJtFTibZ2EOsxhCjriFi14DwKBsWgJj1pp9qmGJ+QNFo1bCivIYB
LHJvmNLrJ/tErLxrnG/WwmChpV0QRSOx2Y8ls1zg6UkBGzeyQM1NcG4POkPm
1zzlmB1P9LHZwCMPGz/DasERZQr1IkkIScO5jSP0uRAgquMIQHAmWiMYnM5r
RluK87ouJvFDbZSDA3EdidcHn1M864aernF6pUC9OiM5wvUxmrYCHHJu5N2K
THyfesm9xgDQTZoEeamXhXbHpD7M43P8tJEssWi/2zmA7P4/I0v3qrprqjsj
fOFNY44q6Pb6cl75Ulc1Pt0Zn2XZdWxvn1M/LyZYUKI9CIuPp3+4XIgghy64
cr3LYsroHMu3vR4GGwYoaRBR0DDgLR51CsDIiLtor4iMhikOtk5js8CqpDom
nCECYVwOobWOKVZ7bolhu8xayAlFqo4dIjAnoE8yN+jUkGQ0tr/RY4DnWaN3
4ZrkCQZtbGRlbiTwEitNCBFYX0Va4v6KrppWPSzjgrRjwT2vU778zyGloTlY
+bmpNwA/W3l5Xy/QLrhesGS/IxJ6hud6j+axwrXNyK4cf8gVVkPZDwVZ0nFa
OB9sfwlf2zVJIoPVDjuwzjxypmbdAi0sqgnQ9/DM2iFP9OSRwHOlbJOwEKW1
iXyyUsoPvBke7Ey/8yGV079wSHWIaIBj9pqiKVlDMIElYMDY3PxkbXjgVa27
Y7mZF/RcS3ufnwPIe04to8bmvRAJ3q3yB5Giya7/v0dXh58GS2UnkBR1AmjV
qP3oU7CHstpCx+P1E5dSsbS6HQn5i1GF2x4pB+xpkFSoEyXj3ADJgReEg61k
T3kdW60M1LkRhVJd9I8+P4mPVPnBUitp7u8jkhQJs/Yx/xhLXTe5GdmtHwi2
L29EvOLEUO7H1lPP5Xq1QtZVrbFu9kCBRipXyGI1CinQX7UXvX5uh7Uj+II+
MNEP2/OL0Hw23KoHngoDf09Xw1+k7ZFMiRLMIzbcwzOF+ot2zQ6EeeoaYGx+
KGUGESpjDbU02iYjUU2NodgztttgZ/ElQzbaAbiuTQjf0F8oUTISdA+1ZYFM
yGNak+MR/rBYnNQ6ZTT23LvQTX1vf/3xMpKUZpYgnLavCVquBY2G+Q13rovF
WfXtZEF8xmR5lxdcXre6Pi6EwHfiqEuK5zbbeQmAakqAFk5NCi0pdQGKju1i
0FKPFP4hJccep+gyGHhzJV3HTr2h11lLpiq/mtf/PThV31PiHDb8RjPQ2HqE
UBoVuGf32ms+ny7fp+whIchMHiDCTfBxjbxLGEllGJYksL//mD788zyBEkWk
4j5oMXTxPN2vRjK8ewUnCWUHVrj37T4QKWutjsAdcJtbiZw/1EJZMZsrYtQo
vIGz6F70PYLw5I7eKodLyVei9w8Ef3LxoUuDfOf9/2QiawMUWGK3ywgNJd43
jKDpOCPEq1n9Nhp+o81IPVyKmcC5s7564A9zqgyZBHIUfBHxlT9mw7/XnWbP
rlXtvKd7JUHfZ2WHrt88bvobfb/phsOsvjtcW52jNfrdKtk6p1K/l4B0yh+t
qDsK0sGrwdd4/oSltVqJpDoJX3p8v7iXmunkczS23YGSM9DVhVgUTDetA0vN
P2ER+WGNlEPLrBxPZVZzJj9nHsa88n73JiBCEVMi6PYWM9C9mZ92OrG28QPM
JcyLIM7I1JlzYgkXuXqEhBN9Xg4nehB3VGQnKbqnDB0GnesPhhnGozOXvLOT
+wTiVeP3yCOOsbwr8tBFZUgg5eYcr3NycbLYz8TEP7Q3iLXHdq4zv6JXNO3J
+aJpMOudl/WoplLrQ94d8+Lu7W58H4SXw8GHK/wgBrbbkzO2P4Nf5ZQmYwiw
Zxzcuffg3H9HbgmgQAnT19d153DAbd3Vwy7GcXyo29FvJl4KlQBWrayFK4iP
PHVmx/3Spg6wfQD9cdi3zDu8Y9qby66mios/FuDfv0Dxb8qH5TfqInCKKAQZ
dbnS9YznQBIHGtBrJTko6Ms1bh2vDJ6JWkCVGKgmTvlSnazRh0h3J6Xh96aG
DuVhGTeLSzNxQN1HAiOmDQNGDVp+BxhBDQW4HC+X/LaFdGzxj1rOrQ1VpVge
JCQ4FIT+4LL4Fx9DpI1nYBuRIT3SkBCIyvGzqjKBlL8hc/D4HbgD4C9IGL3G
0irZp8r14ZTU0V7fbjbhIXXkfJA2b8hQkMR5Hcoy1fizZubBRLR+iU0zf45X
Zlbh0aXYQCkcAF0ETi18EKePbcv7TWW0WWBeUh/vGTRhEvSZdPzxJJ3G790d
u8xlBoTbhzBW0N2mlVXGd7qG0QYcXtTJZtL5dI1oo4+unIVzAPiwMfYoIXTk
QqPjQv5MFlum+fbOWhHIpSF7rKWxsOtzsqdq/ZM2gKAxypBOajFsEcCvm178
1GYGGwhcwDenFGsJDSyHytfAKyLfeqyyBamQvABxznP0gmGuFdT3uWn05E6Z
RiczC65tEBOnnI6rNMk+ExEaUoxNpw98wjaJnfcaCQ8DCc0z8R6iL9NbTfAw
C7ulvWoJXGKQGiEM/PBt+t1Q1iuoUOJaQhZQ/X/am6WXKlDVNXXcuLvbA5sO
F7EatJn5XGnO09e3M2Q4Fkrnj0cebImufJh37EBleM2Mu6QTFyMftVS5cYc4
0xZsiA+nE7EEYLH3gk8rUYDAb7JIY8BsSk9NzLf5S16x5IORrz0nJJvhSdrQ
QV8mSWju9GCXRp6V9kg4QarwfVFicxC+d8pm0K/mgPWU+WI/aib2/FGKAAcN
SlZgYnsEvuxd/a9bO6iOKPZxWXX9MphM7mPnJcRt+eh8efv1N0tjjZ+1krVs
KtWeMzVUyvB9STUEyfOClkZXkUpRNL2wnaxXVQRsbhuyR42IlBjqVGKSja90
SB6FpJMYr/r+0mFxB6ghXTaZcCvH4cnYkSjEcO7Ewzs+6/1OyYbofRShfuzv
ol5vF8+GpNA/t4ymBLUt36PDFitxCntEdP6fYhW1XkM8E23QWndUUlqBTYUn
hENOY0RO5SNEhD0JJ6SgSW1OsLmD+FaIFvrkiuKR6RvT8u7clKdyfFkxNA1B
nFQkXOD7fhcnpWnU83lrSJFW0E/rkMR5r+e3vxbjeCiqCClgbfBWku6VZzb2
gsuEQ9roLGhQNuZPtiNYiy16GQ++6b3KWbXahNLsFjxGb+MzY9Q6AMlEL8l4
fjmHkjldbUYzrFZO4UuEsuDb/u2W55ylQmCQ+rWcWkmSGnS6h+TOI9iCoylA
oRUGG64VER8HmHd3dpyjRLrxSD/4Em5LKfJrC5OYPVcMFu5/SaxDwVfBfBG3
mDm3pztzCv4vmcpnfm8InusbJF4Wuvb+6I+ys7SutWciNOWoh0kIGlHHFjsn
mdej7ycH6a1bbnWPKQcXpcmHqReTUhHvhI1ZVVzh8DCTYNuzDUy6QbiAlLfm
0DSZHnm3EPxUtM4iNqvgERYXy191yK77GV2I3giHtw9bZv5cvEDmPguMqyp7
Zkyezzdp3/gDj+gaZ4QdUW7tRPRNMAUV0taa42jhyKjB2lVDXAIjDBiFdl0e
DJdDPnDyjOqEJrqhUfk2s8R0LNnNc4l4YoE+UR26k7dNVV5WOjw3V+AvCHuw
0e5SiziJvraHHNysMBzjEySKRvNyJoui8P9WTFMA9lf85zqJrmPYZys7SHJ1
U/S/idxfRXQ6dFhQ5Y8pU1DtxSDhfzquhR/iFsARDt0emiXYhH4PY+giNxHC
7FmQBEQ6HgXNNNwfB2uYELaL++TnZPLqpARkROJ2vIJYanTgLDsbFlGC/Ng1
i1B4Womr5akS8NVlGaFvuv2Bkrj/iW9kP/THBhCiPJHeG0uMv2xGwfHhPTL+
l3kZ786KJgBHpjFqcOBiwMW4T3yoJh9yVMRx0jXoUMAe+OKIVWTZ/YB/ogiU
jaZUrLwQy8hupRzbWIvKUm3OBF8mkr/O+xCMx/WlyPRPLM3x7cR7IC4m4BKF
QQcxKOTEVHOsfXag4J0TKaf/dxIx0/YPQF2N/uLgZ+6+FmYP5H2QJDiOs+SC
CFETHOfd2eNBuwVUbdU3MTHT+LU21ksDGhPJowo1idtPJ2QL2m3ODKCO9cAn
KTcoHWPH4XnBXk9Rg1+VFnKnez+3LpYUO6EgNAKB2egm3eQrqVgBw9t08q/D
nHFSYyHIHV+pI1E9nC8NXs4iE7Qf0OCIL+WTMZPvkoR30YH0g7jR/ixUKCn3
swTVR7TEVjPYOCVh735QaBGzRbEry6bbyC26PhXFrfxbGUP2i5tVb27PGJCp
XcRNCsHeMIX040sJmQQI8YGbTVK1zetaGStqfRKG2rbgNiaIEGMFpps88YAm
wMk9/Vm1f0sGRVmYzk38W72dtD1Ed2xrt+LcBKpsE4GB0I1DbSpoTGcinexc
F2xkGNGAPPrp0+kFJromV2PGdSNqikRp9MlUQoUWmZ5PToxW+Cp2ZHDZY4lC
0ySghb95/WydGcnzMiqnaiDUjqc9upAok3BmU5VDIdM8WLxQ8eppo3EHwDMn
v5HXHy/MuzqWTCUYpPdYmxqQ+bSi6xjVsZZ30PptKx5yz8qLorRkbkIXGH8T
0IUfo3TRI0K6jObCUZynKnuav9mhrBpwdxYqHuosPtje4Pay3R5dr85IJhNW
U6kP2edpnDuMC6rKMnDJB4rW4/SaavYBkSj+BN7TtfIWW640p66p2IPsu5b1
U5GjyP2ScL8m+d0SKXYBMJOEa7SMCtOBPnHHp7C/+MnBu2T2opqN4687c/t7
esmZZZkLl8IWH1YOemxPki4zFwY52DBIFXUB9WtNDY8EQy/zZtUBC5b0Yztg
VAgET1xSEejupEAxeHjBDo4peF2JkOrqn5oHJ+SjgOy/UIHbBpLR2mKTLMnF
D/Ixlv2+y7+qXIVv9c4jIiMYmBOpDiWi34U01rRNl0zYZC9rcUGgDYvOVkYG
OBnkryROIGLcR/HIsHEun5JETBsvRGyBgsoyaE20mtSNhJvHy/DiSf5guagW
76motmTCIJryyky2W0PovMFVoF1JtApvWi6TaPlidFlZTPiRnHV9N9Hp9KIO
zyH4F3W0hCh8uSRdvwxNgc3j9EeaC3ayqlk4Iub4qAoF6LIa2F7FmZ0qS6xW
A2pXC7BRXwfRNFv3scdkjOHL2XCJla/VqmKKtopuSxMX1iTKmufDVSaWdjZM
syV5bn8xOLhNdPw94gWNPQ25sLp5qdeQSnmMxHY4Q0Y/+nhBuhkV2+kHzI4r
BmqK66jOIAfhOMTGScVoL1GvZtOwIz9uuaJS4FpEqUcfKQeHlBZoDNSXbHLH
dXfcO4x2lIIzVuNvx776MSad2hL+8MICMqXgMx6zZLSaGaJbxnhG+ktOb/3C
h9pOFp0uAyCH+Ye9M0D9wP4EuTPRO+Ehc6u2UoyQdhQ2rS1ddDkiMwl7rWkI
filevLWaP2sXu0eIbzn2XwnWzLAtKPWULO0P38VPmoz/hPl7dyu8kZSt6c1K
jm0nUGITTvWMzpdrzEo+vgyQm6vCxssmeCX6yaqR4c52s/lfFmy9DJ75apQu
gewFf/v2SFkxZZhHAN6UyqVEDHE0U2O4kKaC0lttSwcS7YL230oaMVwpgigY
Uz/woExryOjtsL+VMTAadFKxAw8ZhRmG4Lz7WkXFRJBBovYEiXy3vSTr0IGi
dY7zMqL71meHmjuXQLEA4OMeVmVPcwdjuiOLr/c9vmA/gyfKKJN+n3UvrZOx
zKdlb1XzC0zx267GZKGkAPkt1Qxi1yzdYO/EW2auL6CGCpz6b8K97IabPK1Z
DAAqZ3Z/2Du0RTnQfvoNuLtBth4yEoMpBzc9gF8PycEAQhkN/mTB+29FvoPO
0KTYp7hIzyP1WZq+IwpxKC1ygegl8VOaN4KcNM6cnvfz07+DwcngX9LP2EQd
LmHJh8zZvgeNHYmz8R/TYg5OkBrTSMb6/5DX2A/RQGcCZwzOXf5PfNkiF/l9
3zvngZL/2F3NPQfl5ZWC85chcVBzqg1nZvwPugaYtMFJZDD70olN6KmVjdsh
V3gjW/Ci58U9MeVjAeulj/PhHYvLgkbqbbvGo5Qa8ahSLe6lKDhLFd8GFFBq
h4NOpBID5tmRSjPiFcKua91igs/HpYchQ+e3sWhhqmLpDLKC338Wi+aBCkMk
ewTcFVvAN+4C2e/G181DpLOsMsn0EaVwmRIZMXwIRVjzbF2Wiyx+4VWWL0Gj
7c5qnaUmJpCvjhYa+TfHElw/PMdnCoRpqaR+2uO35qYdcUKo1Q+lxXKw+Mz1
xeO/3MiY5Wq17aGGRdNznxNB/kFCG82fcPumVk9+rmj0t1tqEGO6yiMqNVxW
oW0FgxDHCu8HMaWQuSwgPLTd2UAh105qgxx28AdFhlJ6NmTrxa3+LYg8L497
5Q5UJe7tuiE9i9gDwFtl/jM0Yz+0TvhPg4btEZ01URNYWBCGbWBRIGFjul7N
jVxnvXQWjOuJWE5Yyq9GtKt5lZlkP2EPGsFZxmQ4r8cFRyHKpQM1VZMEzHSC
imUtEUMZNkXVx+7wEsGuJ/YM+Yb/P/yoRneBGbNAg5r/Cg1VeCsf+VyVnUDi
84MbFgt1i/OvhdRtQq//lpvJzAUQszVe3OqImbMhZKGzke4ycDQsIOzZ9w73
L1M2miAvjYGNm9ve9ZFVDEezu9e1YKehTuAFebMC6vSj7C5AaKfVo50EQXNy
Gf1DC1XOQ62Wyxqb+Q6PT5TI+QAB3atrrpMiqrpgSDNfXyA7byfi3/vebQnB
w2IATlCd4pmFMTaMZL7a3Y1wnoG0bX9/Ne2o6kEmKQNmzjZmWqvoQW+WFiqV
Jv7Gi7NwJ1QgxIwn+i+f1igWqR1Si/TWTdeXY9VbQMCHIgWTScmuio+0fxKx
5GwFMVV402ML3SeCNaD8hhwobS4Q/zUkNYIia8KNb3jgT48xdahv0G/hkTo+
24dZp6nIX9DjXlPF+ZvJFtfPwSinoZxoUs+DoAYqvJR9ho6wP8mQA6ChUM3C
zVrT93EG2wWTMA9Rxm6TltC3kjnYElB8G+8i1A/PNfrqA9/GPDG5yr2SkZKb
9rJ+IxEFk7m5ieLA7Znk9PHM9+Cd8Llle5KgJF7xGv1S4tkVkgOPGINC1C/l
5fnLTnHFwtiicg3MeXGujRw6UW2iXv/nLmk3b9Na4RONBkSq5lK9j4KETSwT
4AnV4bbscTLXJoKxaLDS7LLCMk/NKQ85/KCxZav/ph7d04O2q0XlqCwzNIhv
4trHJ77tIi5sswUpgMLVAJXPBCszR4eB06M48cdd9wqrVqupf25+zUVWufFa
Z+Xk2jForNW7GExXgRPWZVbmTdFgwGmWGTzArCvTntSYZlgNfAXJK0l/PoZX
3pvnHXN6zooJq4MwbhZVHUqCUXwz/6DpTDn+NHa0lF/vpMhurhFSceecR2pE
S8QNUykQIJDIwcX0srHLstwZR9Mr0D3JDAg2syCXZl0dxpPFes4U7lv2fHm4
twPNoW+HPzPxjlxcULigOq/tLweWvQPBZBwBhqydJhFZKnLh50qpDYq+ej5F
dJNG/a2rzeVnQHOVDMSvvpiuGaIO57ZQdRU6vnXuaxu8cVK7014X1H9sQbb+
N1KyRoag7uk1Dj/DEupFcskJvUs4NoIVnPk/cJ2s7TWAk9o+KWbxjkh0kawD
xW5m68bp1TiCnSX/77INoAVMch0bspZcnME0TNxVRf8vyPbYKOhnoj9/U76z
LpT038JuEdiJ+ziGfuAvgA+pISP2dhFb5NRZrf31i7UogPi7bnBgt/vHUPQ5
8UtauTLDDddlOFmaOZIqfJcOti3HCjinYo4VsnI+CA46sCxI3QA2eIKDiX1O
zRcyKFroV/oc8UruLM1/7S8OskCSGrJ4rEKLShWqvsV5l7oNh/CehELdbhq1
82bKEcEVKbrXvbN6WJpW2IVKcdmTgqBIxmIPOkmTQOQwphpLL0iKFLWZDafs
05kSfnH9ajHdJcUBnnGwmYeIdYIC/mh/9EcGOMQn0SDKoR2gMToxDXxnaJ7s
RxzTdwMXtQ2U3IIv/3v5k1VC761KHOxsIgPN58DRXZo5P2xhoM9pb4UEAHUu
K0wp7C4HW9SvNGBt26XHQgyEq90pgzm/9RP+PnEbjS3BrHuj6K7ZmLjOP8Xj
BMOL6ja3cdFekybsPHNGg11sfWPAPazseIn+OMbvDOGxPuiJMdzMMLDYtBQt
eMJpctkXALYTWou+TXZd17P924Qe7rCudLml8cDukxIYV4IatT0nAUkG0Vxx
3ZcFy3in8HnnAY/pxgFhnoyfU3ce+svhEt1UgftEBJKEc6zJ5jTJjh3285+o
3q1nAQ9UuLVwHRZhklSIpupwdirdstZJvxQuSc+8W3MeLCzUjHpfrkqfpQOl
PHr0acH0XzlPNjbz1KkhcqcLxtFmtxjMVy8IzuhoDk0OW2/DybB58GjFz8Vs
XLMpdYqYqWbcW6N0ReTshIyTLhgfByIMu39EOBamdl2bPRX0LG+X2XMP6aPU
eS1WRL9Dq9WKaFH8GzZp8Nw29EpKKPVhIk8zXygVQyrpSToBPWxxtoRvZ1Rn
KVPy0hDunJspBdJvaO3zGAmBFCfc4WhJgFCc9tTtwEN6V6M++ZN33fHasu4Z
6fZS5phA/l+8I6ceQbjnuR3jLDSdZFVUyytDHGcYtqvqn6+o/dzrp3BmPjH3
OtIly98EwnwFf6ThnP8spZrqWt6XcU5Xnqd6E4KTj8LXc5BCJRZr306j2u6K
uaoU9SkhinwtXFcxL9k1pccpTQzUMk+mO14JnTKjKAKW26ElCfdoWyzSUHA9
G+lhczfAXXFwev91m7Z7/MdD4xJVrdrx2wMmPhnHLfRl1m/sRyy9J1itFvKz
yn6s+Dm0FBeF1hPakTRVUgAv8owoO9HTz7UYmTBAuKRrPLIvYGJ5OhNS9mOC
wih6LBUGjIXYJeF36em6ASaWar5QHgXE5kOrnmGXjWPynZe8QeB0rowF78Uu
4LQX200WILHyERvCJTCUVw3Ku5Ad4TXxlefaR3s1nQbFL0ZbOeFrl68M6Qzj
WWhKORRK4Qnm89chI+hVz77YYE8hFRpOY8tULkBkRQXhrYu9FsmmBuUoow+P
Mzg/vZSgiA1bmTUpLryBJxTXpJF6gnGkRqeXWN47MygSOh5YaW73gnsruoK+
5KiBNo+ITJBWFZov/PXp8XQBkGpDzbMP4lMNV3RCS/SMiE3Yno7H55pv42Sa
jRa0TgzAlvBQ4D4Zbqqlhm7/e6uiWsYLl6x396elMPjUHVjTXlScXHSmCJ51
IGBU8lGtZoR+AtSohfkVnQVTf/UzYJb+e00gqCibJQ1e3SQMK28/J4z/VTek
U4B9WeUQ8iHj+YlYmEPqTHRUEqjI1Ri4sQba4esCd7M5V1SuNgfhJNyOIE8z
5p/0NcXh5yRCmp6PtisK9PJBNGeDyghwif7GnP7xkMp2YguRZhqIxnTQZst0
hzUnP7H2cYH1wQ9XYg+YExw2z3So/riOqdmURkQgxgyPDwBWgk1eynkYpcp1
cYTx7EKf8s0zdPMt6F+0k5+1TXYgZ6lMuk+iS44YGPL4C8pdpJoEQRDzP80X
NMzNG8XjCu8jkxLO0NZo6ChaO8XI5CnvU8xM2KJcQzkDLlFT/SGsDwyCqAAX
8v7v7dm3HulO5hEpIO12NonmjJmIg/TfG/Yiwm4r77Rmza/6BsxW5F5BoYMu
OIxbgRQysTAmN2HkY+b8KIIPauOPCoxShhN1ddmPYkqndoSxmzs11N4fO57A
+QsfGC9J9XDnMvWvfu9FpFkVOZowkLGLMcfY6Bcpl+wjaI8iL9bje9Jtuyj+
viJcjy8wkR0SX29EdhlyVr9U/QQ8qlRlBe820QDCQkxoOSXLUanT32mm8CFv
kIOPrYGeoho9gypnErNYH/e/LenfdhQzuUtXGQQ0XuE5Njo4EPt/Ik/XAuUj
q8vFEh8Y/qxP8rjlYEikJuqRwVn3MwcrtYiQ8NDygQR8oY9Bz4U7PctCbyxb
HTlbbmKiHH0Vjq9v6MzTn9RDPUdmAyLTNt74jqvGBcn7GHjY6QxN8GuuRNR1
jnrAhCrC1PyQivGOipmH4JU5CeP53HNPw7EcZtphAG/bEtuKX5gUn2hxPP7f
hb31Ka7fefYNwqV/tBF0rW9G5XRYw5GYD6sAqY3Irp8DN62+BgGDswqm2Ft0
mz/Cxy9nfyRSaBSWiB3S9LypRmmhE8onL7XBXMPUGATZZJRB7V9Je91PUzjx
9J7SSUmKVD+mk7k3PWFVsAch4pzKmAYNHABQOkwqcWr5Ngh5jlb9uGYBsLyS
KekD4KfOIkBNCsiXeq67Plkb2pxgIBE/YnLzfXzxjOceFehJFjJH8YzUcQ6Y
UuYvgKnlSuKlNWAyJkP8ICo61NU7XxR4zsNTmv7QPuZ6Ep6vwpNQ4zp1nbIp
F+TQOZqMpYYTWDkWRN8NI+iIRCNm43ZOyJjKWf+Q6FpBauB1xwVJOqVxdCnF
XpDIHMBGqcz9qVK4VlLtTKjr6kfkK+nnJiOyiU8z7zxgQ/5+ex0ikFSfi0Wg
A0GJ513GjbK3me2DOymErZH/U482J1Fm1T4uQL+0gWYC5Ztg/qHIn6x+7idD
aGQI3ZUHcqHkfMti+l69AQy0Hw87ki0dw01qYkR7+Gc4/cH6uplp+Qln4HLp
eFqwcTu5eb3E7tQ2Qz5Mv3j/9GC4RyqvM9qE36tfxPSR+y5PGT/q3vA5n698
lg+WgznkjoeSx7Y45+qjBP7TupClCCKBTeADovZPoBQzKdAIEfk7eZSUmg9m
4CMtrUD1hGADfSUSQDZ+HrUd1KnDdEZYDncYPqjVIn5FsxcKpNaYau6uJ5Vs
1mnpRwph3XUCmeFYVkJNVIPaBaU/oDseH+ChwuDiVxBUVcMRFFL2H8vBxhnx
WeLm4/4TYdpF+qCfR1UfiFnGv2beYUp6aU702/Dq4f2ozbZw4uueTnZRji1w
VIFCTQZoOwsW37LdQiwEqXJncOnrFBoV5TSisiNASc0nH0GUODdSBl/DuvqD
q6sNAlt8taArpuJEDcK4mCyF2+Dm6uNmuShu6WkO+FltQ8upr5VgfsWkP6Pw
F+CIJ+C5sRkl4m/YvnKvTdI1zRtjVHu6xsCaYP/zVd6J6npQxlIUiIom+5e+
aix45PFZ+O/VFCGJ6iM41qyNs4Y41Iwp+JqFc4Qa9I8Gm6BgISjuWW5wMgRr
GHZiGEY9PDZ8xXTQxSkL3o4o6fdYq8kRksw5w9/Jc1c4UlQ9nhH1JA7SNal2
UxVMDn+Gt2a3Y8nGWGZkAyuKXffk/Rj0MHLUe5s6czUoMpxXc0TRHMIpjGIS
dWjcJ4WmtstYXl0/aZ0ku26r4dhoLC1wcYc2umHNJnYXWaRDpGqwbayqy37r
kJGolRcsbfHQ9elgCdYpEWYc2XlqkwVX7JenjRWnWIA9qPDXRypX9ub6aCsR
CwJoVdvcw8qWKvL6d6J3XdAuPsqenuCkutAis/kFwp1X4Q9prL/38YUIRtRt
8R9VuuuZjLqYpWRqHC0RKTIcDHg59PqYfSbgsXVOcpK8ywy8YTzjO+T1LkCS
gtmorxw/P93ZloNzYorLeKhnrqsAM1QdAtGpUGIT+KJfbJdKySdCGY9gM/W3
uqFvhSYnI0tvkOviljjEzDg6Mglx52P7dl3qgsp4o9IcakZVwDFklBufXpxo
qIThW9jqWbuDZoGS5KOhFCdnBMnjUswjaNr1FKQp5+/ZPE+AQ25Lzye06Pqh
KizLMGAOg2ZKl/Jgjgw8b1P7CPIJaSVaIugt3R9SAWGUkCYwSA1pexmULf3g
+GA5XeSQ5TN7IdvkqsIFKEp6i/U9kIaiPWMgE3CtGKx33CjM/EwnAD+reL9B
je9151G4u4w/EfKVGvg5FneS6hrHVOEeJOqVO7bX48cRbMzfG9gsBNgA8oR4
WJ7oe5+xAML0kW1by8SO7Qh7vMPNzTVGHq0HzxLdBYzI10HyqNwsSI17o/Sw
788I5WsEKPorPnGH9+u+nwSRRGoIL/1NSocCY6HqvbgaKBvTK4f71Hi0TIBj
6JFm1OPsO/btOVWfU1wDSMBJZfA9fmvT3taMUAOCEmdpB7L3LDWOBv5dYkn4
jMjhst1Y5OKMUdliy5YQhYTlyvvj3Ee7uM+Wo3GB1Ee8gnUfbXyxKeXBQj38
GenTF8X8iPAVCJv2Tnhcvk0f0h24cMwPCjuj+F74goC8IgIKRqiPgKuHEP10
bLKfrdCdx2rTToabdonZUBbR5pIA6huXrwwJIe1nwe7lOhgXhqg/GKm60h65
7eCpz8XHhPzQ7goROqR77H3bze2wBkeJwaCxRG3Cq/Gbywj7btalD33IQRrs
LSUtYO/i1KWaHyKW2MbXl/GzAFu8UBFytLC9zfJNwYKV63ECyfudSWtpdMUj
JYHkY2YuYzCluL1xPiqumxAky+e9xJTT2hj8ptculmYiFCRzZX5q3k5D8C8E
JyUTiFm7lRgADSu0zhlm+MuMsZ+nT+TMFdsEQu6oyjZJ70lMNZTC+p92rMJf
Zry6DTpfRb79Qv38SvAF2+y3waJRvQAUETAIKvPvkKRgf/0TaZ1j7X3Rvn6C
pz9vtrL4fKFWBLFJ+Wt/KgC5dtz28tnAVd6sCOXjGuPJhayrKFsiqBpiGAyR
JX+CaKOj6esTHvj10aCTIHuWJEV99k3sBmQ0zMbTt2hnIwYmDtMVojG7r1t5
fJKj4g1qaKVJ1j9SZWz1KGdkm6YOo+SXoRoIxHY/+2VOmQH/oBHfg6bTeW5U
KVx2x1KFBWxlFsAwUw33BFp0ltThTeouFRyHLXRPiUDmwqMug0KVQGrSpCMO
P6OUjT32tu+JCPd0WLdsQKsvKmI6b3YYqmfWfYxGkJR8+SQf/oTNXaZ06LnL
AmWFXFxUaL1TOwMhzYihRHCyTnu2kRUUbB1T4oNoveyhVA7mk7Srk+4q5GLh
2xLD1mYlKWSLAMUeG+W2xGfbdDwcusRUygMwrM0GkLZzq2knFl/KAyXAMgdB
lKySaTQ2kiHjD9DKZn9nKk1Ju5Dosl9P3gWT8xyjEqAMor5AhgWc9mqCQpXV
sbXDHZhpE/mTyQOotYu+87GX8Jtsktb0UkEytzp7GdOxEqE+6PXNBYe53DO+
F0/NOsUdgsfyq9HUonv6zLEcwgGyZRn1i4ew3Dcrkq02rmc6kP8c34JMzfKH
zKBqtLZEFMNDJhIfnDh1fNWxN5lBKnbm8qVdjF6ZfceMTpyKP5ayrksQVTR0
GMUkiKtBKzfLc4U+KibXOVjc2dFbHytIMzztAPMUdBn6hPhKzO/7mJY5VFE7
kgWYZJQZW1rF2WwlAKzeHOtGVxzohV0wikSokqL1HZ22wzxvmfqxe2NIX7rS
1rbR3+t+kIFQTwoP52w7HinhDcI/Y+iJeIIikKrMZasinVja9FkSgZpFekAG
Zj3daOC3gwf2pPUnHEBVsWkcX85enhAljdxNrDEpfZcKmKltQwHOs2qe7DXA
dtKVWC9nIKDWVAEm+ABjXuS9r7rnq4AuBmIF5ASvQLXfsvUrT3YR9U2aqmIX
4sPeLF68wN93Kpaj/i4M4wM23jzjXUxBPEbHJUkgnjS7WW3c4o+U8Wohk1nw
NNoXNy6xx1cbefEAkQNhrsFNKGtgLxUe9NkSdFySeAQOlX9o/kYEnLX2VqYy
+gcWeQwBG+uU2+2193ruS+BO7oXk8cdS/swFwfy3zcsLdYRuUxjFg058h9cf
m2eUXVBYRvhv/m1WOnb3RTYx6mc4VDQo/fqfTjxmF5XCU7eOJTrU7DAus3he
9Ee8c7v2kEvc7FDJtLQpcopsHkZYJfqMggGHUSCUe3UMQ5LInFuBK+BrGkSe
x9Nv9VvnJm05h4S1n9oavW32FoeZzzgIe1ssHQIESJi5Qv1GgY1KBq6Au0FK
IYYCOksILKOCs/X9dk1wgxCmc1ZL12PnSMzQ+2UaeQQW+R6vBBqXQLgk0Bjk
1RPA189Ad1IYVjDs+rVWvs5sdaOhnhW+s+7NOj286kVVEXaGlPgvtcOFmL7c
4ikmZ00+YfmRRTfCu1H06tnrGNQG7tCIkOJ0FcBzoSu5Qx3q8W8LwZAXCHEM
wwnoXCPjjQulYL1PjXTL7B1fX1PlmH9i5UwOMWd96hTRWLKbKuP15nxPRDT0
/+99EXi3aI3eflyHnYLYelgo1J8H173khSpF/ouNhgNx6TJ/Q/Aj1BW/bjAK
eEGqeXaJXxvY1CyKC30Dxttt4i3rCpXv/NQHQ73KH68KjsoVKpGVQVkB2VDP
Xidd+BjLLiLZolj+ds83RY51fpXBHP904vAaPLdFC6vvwnWqPrYU2OD8N3JH
Rd0P4WSA/9Ifvo8ibaHhpsN8trwqDwPkQ7fFI/QO0ftfcrG5JKPB19nwXJ87
T66CvrSYYK5+Z8lpPxfH5w1ezAa9WQCevckjTD1lMz4BdN2BNSDRmMA6Trji
K9N+doHpuKaLOq1aKOmnGUsoIXX1ilrRR9AQU9+VTpBRkZF8bZzMcoctPToj
Q03w7C3ljO1yhIGnv//jwccyjR40fV6JcqfOH9JLQYEhNXrmxoIc3xbRXEXO
lJs/HtfziDBfcr7pVBYZveOiwoPZK1EApnr4WcJTibOf2ICKrE+vP9gAuvto
wv2KrBbsxc/yYv7yxvr1r/V6KfAOmWXdXNaS0IA87ZL6ZYrS6D5uYGGBepEz
Fmup7nWMa+sp/a+y4siCufVVgqsSGVSnp6WQiL+oTDsYNx+JEHGQdmA8MNi/
7jxvIa7K8G9d5j1IaLMEg3S8YZg+mjSnn84/3aN3BX5TGm95oRh4cTOS5wOF
JXpz7570Tik4kOCFQp9UZ/vZLFd6RyuMVTDh9LcR3sg2zLeqrRg42kKLOnAm
eda8hl7HXuGjSuo0ZKf/PbmePlUEUHi3vQAK2cjWRLRsJPlSDVUk5BV02PB3
a8pKqURXxteDzI53gNmPbaNk/rNli1kjjRAraWd3jI60TqA1iJQ2ikhSEbxA
b6dtzt9HTUEPHiFPyIa9omM4RXT8Ubk5o/pA3aHWQ1Zl9CqIM9QzjNqUsjSV
iC2CJDOGr/ZQcIz/U5a/9nbdlOQbYfCPf9s5dIBh51VeE5OGthUgUv/SUuOK
Te9jtSHmy676YGutNhsSEGV6lLGZ6Vi+IEpKlCabBS5XKDPf1KEOhn8WsOGl
ErHWWGRURJADFdmiIkvNKXHbMFCdcFwSgF02UDfprl/ZGMaPiiE+mt2pFcoB
abwBa9yWBE0jGBS8zDZt33ymiwwqIGE+sdNrPNHF3wQIME808ur1b4MciBLb
GT1HxUbnDphWJXDptm4hq7OsjaLHwdBhqut2lwEXCjUY8fyNrrvDswbn2Bgf
KaZ6JrmXztRWvTt87iCjhwkoUKHe0eIGtyCuE/y8/eWAktwQboqyxxcKW40D
LRv22RiWLQDukVr5M2nrjNGdIzHD2q1Zg2zHrYnn4fFEv+KFHmOLWgZMCpDa
s0R9a8xPxZAhls99WQuDf2CCIQMe1a5OkD4qc0RwdsXSXYc1X7OR7i/Qc0ep
9I+EJhEmlfcNc66Ndg2Jzxdbcui88KX/FsDMOc+GDuy9ZMHTtGtdRJocRUmM
DhyQ94cYzLWvfAXm8zIUmKrZ5UHY54AxWshlfHBCYzZZb3S4p/TKXJumYuWx
+YXCJqBx8An2oel6Iv+UAYRRUnK64QFbB2Zi849NHKxwiBOgba9erU1s7xMu
a2OTKKJ0qd7LFuysdonrp1d+mWi8s0mItwvPMKUt4+FX8LSgTYUZczpgYGLp
TxEjTiwfsM8zyEMKjt/UeYswhKYZMlj1uy/c881LmyI6pzg3yzXvg79GqdiK
barzYDQUEzzjn22SsYROGCoL8bSftB49/qRnRgPkDG5zszTRsQVOcKlUTO99
l6R3w6luXN8w4vQR7r5uV6KiLMJnNj/jY89hTwoqXMVkAixEM51RTKOfMe4S
z06P6C+gB6ezAZDrs/ttMuUZAL1OPvK+8CC5ovQs9EhquZr2zFLZ6e6kRMEN
C4SdkbhJitcexmilQWcQKys8ENnZP/KTC8kVp1ABeNp25p4UdBeXKKksDOcA
HRYzqpC2jP9YuKzqDDkq0/bgZl6hGUYzg+X/0Y1OQgbLtAS3u+e/u+O7bmUN
/YAyG0WFXJZzlgJMxrKevuupmF64NKUzcN3Mqe6O/ITD3hhPoUU8AiPxhO2s
CW/PTIW6fZD+mdWlBUWS8qtuHjgEn83aEKXdQODufb2g1bXgg2ID6iCZl0Xt
YkxcCFgCZFqcOG6bLDxt8uqVxrzfyN9/08ruEOThAWc20TvMKl0x15opE0rh
12v0ARR5rI434YKEkcHyQOAg8+xVdmek0Q496lAw4DDvhrI99OqXxm9EqAaS
hTxhoCaTPlgyCAZtOQhdLQaSQnI1K0okmaAmh+LO4bSAQ3tl0NsHKiCMKuQb
jSQZW499qc7cczte1Vk08J5iOLlVosNTgJgk2ksHm7lOPX1s8k1eNp1ZxPME
hX9iSQEgrsB32ThvSQYQMTPvxT590rppbCpafFNvtuNV9H3USq7AexKIs6j8
G04imh8lIdFzUf1KliGAeifE22N6R3+xoBaAg+bfnFsib/hy5przwrULsbpj
4xofEjPmn4icSiQn3/AjEg6pGUaV+H3Ts9l6v7rLrsblZXY9AjoYnU17kOWg
PNSDFeV0OsKABKOaobIKMvFLkmvZX/OPrPnsRK+CBK1G+jsQX0G1IcfpH+lu
WfRemh+TDeeL3agB9lpRJCgDq8HgHyxkc6VleeNRpk70BF1YVeeN+GCcvGX9
KQWzV4BOJC8rQ+w4myC1BSQlD73nMLhnKDeDU2RKyCnUFnv/ps9ykr+7LgV1
HijD/QTMPR+gH5voXHlruL2hhzEMB2MlFuYXXWxZjXloRHauNLiKLXeOZNcT
vVMIVTQLbycbpXq4dv/DN857YNlY1PcEhKxacMUkVq0j9s3MU3XDxNg0XsXa
mJBx2yd+LmVlwSB2feV3/8QuKouOmgAZKCp3hB8kTVtsU9ur2UShZGgeqgS3
qo1YwrX2vzf0+32y7GL2xQlOwHWuqbXEiOmFCSUnNGxNLceEXaAEvEW4uY0p
W9oW11sibF7X1GzMuGLooRc5InfRLs0AkzXZ5wdXXM7nxj5J+CmxDWTT6D6g
3P2EIrYsQOtEYn+LIdvnN1r9PQoQsryxbm1zsniVlTfLdzRKvVs6z0OtMUVi
AYKSSu74Xprx/H4f5pUhjcjLa/y6414OV/Cia96b4iuOcb0OskseBUprXQdq
1kEY9IEAB6Vb6xbFVYKjR/oMD8AQwgSYOTiL7qqNWRqDCumw3Dv/Z9nQ8PqJ
YKX3IiBeXQezdhlsU1ClMcI3LilZ+ZwsQj/9DWlflpn4HPZ8GmbnvsgyCE/e
4mpmQIzWakZnUbjhbZi5qssvLpgXOQ0Z3H+kMheZSjLbzTPf5bBAJ7kaLk4t
rMj8Z0hyeMnI/I5mGU+h7KGO/6elFlKP54DlHQ5DS00zaNaqs77MrN+otCpY
uqW0zIqOn7k3LJ/hAu3KZyxtVB6w6ID2t/fvl/+191Kt6Mj7AxX8d4heCxdi
J5q/532g1DpJc7uWWatWErzyXy/gcYwgeGf3lM52m6QLuefQAFD46KgRXy1k
RIJJ60ZGLMmKZ697VPX50ANLPqXilHYA0qm6rNOO3OcH7lr7O6OXw3UUlS7l
tThZtxEspQ4HIob38ZnXTACQqQrIeSl+VR1yVjj+himctaTJyhPXT2wyln9C
nYgzt1cMfasymldIGOxmTY/TL/NWsi4fdFAy0teCbwAHEB2H6uMFjkjy5pBS
LsxJbXxGY391469f0mAe2uxtbpYMHkM+D1CMfmmnhmWYzDOLsTrDo7ZdDJPw
emdS0uKeikqaz88+/dSc5BeXCZOZun93/1TUk+0xxzkKKZmX4rZ7PIXsFJO9
QlQbgxn6VKTUYYx4m0XYPimhCKdv496Tvhaspm0aKcIM7yMmS8OjPSz7t8vv
MvX1XIemV6ORuB4A/Mrx1t9CWnyGd0wSinyichp7xe7STbE7zmt5BWbrnrWX
gpl1LgzeZn7A/a7aP4P0Bmuz/dEmuiYrKlncKITnI4TObrRAKD1LbZuisaxM
j7Ellr01RVqiwCOQ3lub+blrQ21yaIvjJQezSVr5mWr5xIjJeQsmY4Nr0vgd
j0OK73QmjyYQ4Ldrcz4q3eSrP9mTU4THqhIjndX7cZwrJaeYbvFAfg2UlS+a
CbQHIYh8rUdHcsJ0ZOOfIjEAgaf0nONaf+ga0KDXPZxVW16zAlPzj/32YWf0
A49S6Ccih7qLSKQCXemjgvXILhrACRFOBUGPcjDWQnL7TavyxQs8SDVaMDnF
SNL5wFDXEo4CV+8Q+2Kn5/Om1ad/CBgpn7F5GpLINvRs5DZpZ7xiL89Pqxea
WoCWVy9WJD4fXCompC1KBft326KFiWyp3xNQD1Ni1QzSMDUGyWnGYxmmxsfT
By3L18cJtIsMMa4WoAZG+8G9AfsanUeMHNI3XtdFu38S7NiZebCa2rAaIKqf
8RDvDHvoAziw09Dkof2tEFG99SWlR1zRFIG1+3UEwT4NTylaWk2Y8wCNg5kL
Ck4RVhsq6vB6S9nB4ZXjHkj9KYR07a5cv40pKAZ9SstK2mj/ePNzHMPKoay5
dAuksHsUfRyY9hlfglB8LIP77z+QkJeg34k1VvSqb8qIim6N/WFsCJhZKQnY
bY8mf1HHE/jPLg5kwFsYzyvidolgcT8PL1r8X/LTzqIex0VzxrGKiaTvZCd2
PqxPZdLPTXPedK/NTs8fgjRvkiM1+I8BJOHZ4kx7wVKfN7pYEGtwG3B2xVeN
9pKrrLs1oFPP/c7DJZlYRFA6HYBbyNui1PwCGMQnIDmim+n2OE784i9yWzoB
8G6bIkp9DDUlHtIvnm6E8a5sRbKP9a7wJGkK1LMpayAoe31WsKXCKTGGUkEG
aUW9PVjAt3on3E1HaLAnlKGExo9kcSj2Ck+FWhPs+kyrbMuM6UMF4pm8Gj5y
uWW/V4Wl5OdOv4vfNjTqbM4xlWSx/7qL9KYxiZ33c2r0enXH6rW/BSv0sHyn
Nua2las0lMIAGyeSBlJfGWqI5EllpS0aIwk8LS1RhjIhOkocs+khjdjCdd/5
HCeRSJcu33UEnR3i1p6FQLLdg9nC3pE+Vs3axnHdutYVQE27pOxadjRB7Zmb
yRMc2JTBmtsbKmKd4I1oeA5KbNgcDA7c1MD8zIKw6RHquSX0tA6M6vPLjInF
JQmnCkmU7bM3HSrEW/3IaTlxkL7GtV+jBm4t4hiXCA89PaUvQ5M/DRfEUk/t
9fpSFyqPIN0VNgFZuXaJPxVZ4eGe/hngjznSjC8PwLg0SWF6BvW4MBOkBJWh
8us2SK+QBBB4bTzCmVwkEuZkNT0ZTx9LSK/CeTwcGEq2L2kEwkwnuFPnBaVL
zqId0ZHC2uUIlxd2qQh8eE+4xXomwKMv4xMAN0uE7uMJp/zqi0iaq9lyHfFf
AX8U+RPhxGWlfkve2pDYjxvGGCe0aI2S7RBo/g9UF23rlLT0MG/KA1UcW37R
c2CL6+fcejT7aJxRXELeS8LOJtndXMDXbj9ZEQyB5b1UPc3KhlEXuhfWjLKr
Wz6laGa2oGF6vPAE5N1oaCmw77YOxc2SszzNgTFAmEN0my/6BEDSjj4Mkgp4
b4VXZF9PVp7F4/5gbIzNrBwRj1hlR/e0Vk1OTyTJaKrphF5qOum86hjECEQU
9joCcVbOGfdMwrhR9MnS/b6IdTSjt05sLWvvI8q+cHPtegMYqpBUVynN870G
akx1DOXE2tAahUW1Wfvyun6RwVLQkzg/Ib/nfN/QetjnEDje2T9qVNlUg3tX
fYg8Bt3NUMq7yEpoPToAMn4sYq2hKxhH9BV7dBlmnnxAfwNAPmzVEZW9oomD
PNe22uT/E61KFW+Dxs8EYazBRxSgcQkBqNCMJHy3Zm28LpwrwneVJ+C1I2nW
O9cVhLOKR/TkI6gK1Ne5tvXirV3J7mXaGbo0GCJok3mzPvI4t6HDgV7OCf7i
f0DSOVdWw8O4tl96VQQCV6jICejaWr7xRm2+EoLW1Tno5PouWHmI+3VIHDXm
SMdUop05oG1H3w0LOLq6BduI/r0E8DEozbQG51/LOU6Z7fI8mvfopCTbXIAa
RaGbAqZSmKGDar350onYjiErN+2jLMyuKKjZIvvQm9M6LQ/2xtyJb1LC+qEy
+LGHvw0owB3CzHFaPdB9tfMz5U0EDQokpA3ZSNTHFoit5xWLCsWfkVIqSqvm
HEzLeZ2BcW0IkJS3CPfiy9LNp8O22Rf9cLUb036UlUiwUNWVDuOvGoHLN0I+
Uo280lN8lICaUGCaztqYLyiAFGhCSvXc4B/CJfaHs7gm0uE9vUzGpuFumsnk
F0JPiEeG054TrcSZmP6yhE5fb1hVU8CqbQ/S0yO2PTWKis2lPwXsYN2EtVi5
zLCuvvLMRk2VzlF0E3BiXPEMhEFvgSdnRBnDP/TK8jr+kq5wwIS/sjgHQiqF
nxfuc3Ek20Obt1v1EBctUs0e2khyREd2P2zguxCCjNZhlR6qp1g+zxtvPgc5
vZ9Wnt0v3GEEj9n0DHtMklU6AZmcaI5LEd1j1zklksFiKOYDuD+RJaxfoy22
YWmRP3h8ABui+L7EJqAdIO0v2kHteLutx7I8YpqYEluiLnkgTawAnXI5CK3X
PlQ6sxKzE0y4tzLVXoxRTkIp2epwNMb7F7OHvydhLTKbCMPL/3yjLgl1XfjG
v9ytx3wXGZZGqMnIpp7izm5+jbBURqNqB+LkSAeOugILuwJGcwVG7j85cn0d
VFUAmPEF9enE58is9wx0teLibcH2f4QE45sWcJIIDKhRqh9BDe1xW6V+0u9G
POaRkIukSJwdvX8fXo3mF23K5u41swhfL5q1xx2b9273rEhRK/P3klRj3RZb
2+OOBax3opJd2ngidhIoLZ+AqNckFaZ/DD37PWu4Cq3sYj9aJerX23/LSz8+
xZfNcDJO5yqA2cl+77Fn6mYye/LTbqwTukVvZfMwQaQG73H337JJCCRhQbJv
jo6CIxXBUgmDtLIDhoCDvxt+RqvhOytmLnWUe9YUskXQg9Jc5rY1/PaBjmr5
tCCieIeheYtnC2mShiGefi56gzASyHxXEaa5ADKywRa/W0LPlw5uWaSsowh3
h2uIFI2PxqwkPH9CKBojH0qmhLRRtYvoguddbL6CMnHsrwoJeUGHdbmvvK80
fiKjngllmfpEB1ESF9Ltt8wqNMxF5Vk9nVpolYkr55zodhcJ8dJiuG1Wk/EN
374MZKu+2Gxmzai6imGQPY2K8jUM849DMg1+lT2uzR7Cey5tntIYpoG3kQkr
VeTvkkh/JFJNLxtGUt+Smi3Ec1Ydd1U0VCNT+0aosBNLiYjerLw9BY2Ezdb8
aGJf5lHXoyQSjZSzXWEEYJBeC+Pz8rv2KyYBv6yp5jL9oxAlAk1QPyABQde4
WBEic2FigOIA0Dx38DFhPwvv+PNBOOImSDQ6bDq3KjscVTtTAzIMjRHzJ8QO
LkkeCEKclYPfphzO3BwA0xb9sn9cvHvVEPopfvR8evRP8Jg+xjPQ9ML35tFu
rE8T1HnQTSsUfFGVxP0gnON7WIOzEw7Josdi3yICG8g1kc5LgrzMXL1Dawc+
Yk3Vwm+7v8yPvi5a3jI8tWb+1qqegNq/8nr6LUALP+Dt8ekCnUqrbugm33S0
VLtSj8lNY+/14TkamtM+H6gwxujVe0RRTSH/n2kDMucfKMMNJG/Y8DMNbOrE
Qmn+ZseLchjP1sx26Q/ti6RXvfRKGYSp0s9QQVBIxpmmC4n2GJ0rIZY8jx5b
n36uwD6fE7WAdLXma6fTG5XiIx/8YESWDUUWMJQxIH1BxMWBoIRtGszDojmo
JAdv5ANekjbUzR2vXfL2FgBWIuUPHt0UGHkizKIr+1tvTM+FqIUex+z6MZHP
HGGLxQ0OI5n5hng5uBSaEbqp3RwzJxD33Y6V3ho98u9RbFk/ui5bRB1zgPOf
53NgWSCOjMF4PsQ6dsTMO+FbngM9hF38mPG7nI7emzVOUzMH2g2GwUJsqAoA
p/D8lK1iQEcxlK287qYQ8YZX5reKGnGW3Ua6b1QGjR6WzxrQTf857UvHZf5i
lGdWVfn+Gle4dSAoXp4wynwmZzOgd5ThwOZxpI8VMLZaQ2Pns5v5yXKpva85
UQUx2rze++8B8AL9Q4VksOTV+Vxfw9xP2R8Yc9aAE9l7s5VPt1P5uaa8ftWu
H9pulrGM42dy6vdpm67jBaAQVBShWseshJtXZezUxNHMqXXdi7HVQnv5v6w7
m9GNcjWV/uZHXgv1cMZ5bd5FN4wcNuUtWhVDmVe5mjKKQtPqA67fVKTsNRh+
ubwmdb5QZHjX8V0wkS2OJcDCzLxCkD7hhXAUEK1h6NWBk6u2N5WFfVvtZCoH
angIbS9qB49y0+ctjI8UlJYo0jcIiHxLhCVGvZihSLXdj+IdV+t6HoLfkiG8
sV+bB6Pdc1tpa0zarud5+FSK9IneEnfjS+h8yP+XeAIaxj11vm4bX5NU7lrF
eZzvua7o3aoTPxDQEyZ0xUMNxZNCchzo+0M5jqWsPzpArfxD2UrHMkLGB1Ay
aqoMCOzUDWn4Z1Req8qCo3kpQ+SlFl8iiVcBNrUB11m9WfAwYhsmvQ1JHytE
Mtic9uzxoijZnABRAcbMHItYWw49/InFKQYqmhMbxS+1iqSNvmTdWy5o81Eh
BdY1E1CsuBrwaCc3hQ3OHjWtPrAKzYlNEo8R+ZgqQ4exRwZHcZRlGI22YVq+
8f+MGctAz4os9LXz7it1HelsNGmczTRLR+Jj9kJKlHam6SzaSXfCH/SmLMa0
OubOtISs1Y0l7u3ppe/+SBUx9dhbe9LChl2c/80E2kmuFOVE7UCsuM1w2/8K
YjivoC1UREKJSMwEdiuyxdFCBvxHBBFuC/daxlwp6QsLAYmqFhhj3EIX6upV
EAI2sz7+z14BjmvkDBI4q2NZP5boiCJqLolrjmr+xQ/licj2EMeOR9851oj/
Dwwj7nnknbcqa6epPxtpb6jSEGRwklmMU4t2uTCWIUh3zL11ACYuqUGSjL+V
hFVzLDzM4cGWDEfA2KmhPl45OvPUZkSh8Of6p0vjPSRCuqqB0IAEvRO9vWGf
saYH/iKHq7PrfB0xvV/4urbDB34fKaDiw3wQy+7yT9cdeYbqaljI30turFR9
a6WNWYUnYG67H3iV71v3ZNcuIfOBCgYeosxQShd3gBWIiwD1azfIC+gxKSlK
/xebighb9WXDdtT6YOpMVuzrghh6LWrhPAhbahGflaNM8gIpgAfdsPh53A+p
hbQrcbLS4eI+G+cPhRE1RD6d8lyVv3RjaICoaQ8jgMtamwo3kUuchUKQ2BKZ
Viu+X65D7GaNNEiFhp4le5K7OxaWkLSR2Br0mW30PzKVPdSBPEqd5EQAlH4r
Vk4sBIJKKoz5XuHzea/3tQnOO4mJPYk1oFi/BFJHk1vI3Fyt58JDux93/OAH
cmqVRTREpRPQ3/FaJglAcOQS0zWbm7UMvvZxxY4zoVqbxBS5UnbTji7sRKoO
IGJqKPXmWEB/M6HEzHBmp8MOOngaIU6BqAe/W2nIOeG2hCz0+ezuHG+Vz0lU
SW4H86mIE9eEwczr/hMWzF+6yYrGwelaj8jw7z+LygZgljukut4xmCajvcji
lTtQzI3wNC1WtbvC9AoSl17gVmswTcPRbu8AIWVI5ul1GrgJDCAzDpFe1R8L
AY0DkX0MC3CkC3jO5luiaiWoIWMJ+UdibFXCgDSn2ROg3Zp7v9p/L18T3+y9
PeIK9RZfUgfYxpW4Ca7BT4lvAkKTxYvf9kwaXEMQfuxU43mo/FB2pGM6To7S
yrhM4IYKvbG4lH0eSoFX3jUuYXowiL8sTQbTDOanGFTQ6i+DX35Nq9I+qEbC
MlEwHZZr4KlEyvqaBY8hhCcbIdXjzszSPm9p6vABu4arDTzzLV+u2t1EC3+c
aMX5G3Yeoyk8XF1ucQD0LdJiBrxCMlqwyw/bmlEd9sgXHwO88b9VtviCP/hW
SrZGScUGnXYPOkoQ1NG7vp+/RNEkrVYsl/aUlc28Mye+M9IMq6POxUfMxwQr
wn/y/YWSF0++cutvThd1VmqLd9A65qkPG7PWG1SBMaM55dl4CfjlwT8iT0Df
I0pDBdh8fG4h7j/wzgTYJrCpetMdMyQsym+3rP+WgPtgXrQ83EL2m4pa+aAE
laMpo5Lk38msOniBa5oUhXNSjokv10l45mL2udUdQPygSHlcVNv/4JOwZF03
LcXBrw+uavZAJrCOxCV06czCIIqc5a8EgpcTn4J/ma0fUTlVyES1P0o3Ml8t
VBM6jOmllD0cP0E002Q9VHgUUiZivrPobXdllXrl9TOKhLOj6a+OHjLznBdK
JpmqVqeHNVmHczyhmGNOcL5ylQwVhujcpAHEWV8iieZkj0QQxUbgwQcQ6LLG
UtwpT+goZOoDvS0SMPBqKyS0gDbTf0S2rX1SJTLKXP8cPbOBb94igEERg5Ov
6RLfEliHSO2LXZEN3Sg9ORYt4so9Wy30hli0HA15+OX+d3NH+O9MzJMs75J2
4oYZjQxOTRWW0oZdrqWhFe0kmY18XC8MQCtbpHeIHGDUaiVLx9QObecr7PRU
YLbc2ilCU6Kvh2VKSTxYwQPioXANVhsHwcLUT70280K97Onc4EqneM4jIchJ
MsBiTa0eHIThQfEc7ffaDlZCvzYEo20A1Gz001BsO1blIiUgbXxkrj+X+dXd
aiAmsq/RyGnNkyIXYV8cM64eOMhJo/AM/0oHoOasDM0TbJiXnk8Nkd3QXj5d
49OVLerg/IOO6VB5GNIifgHs5aKHrsTRT9pxNenWcbY/3dCIdDwS0S6JzUf7
82tF8w4rT17MvErn37DCSHrO0GHNS2GiJF+4+YWq+se1sf6M9dBA7p/lQWoM
nQ3TByjSZ+kUJhXVwDf14pSGFBLdOtRAIQLfQlwO2tXLtChq0FNirAEa2yPc
1XLoYfq91FcSYNk268aLGTLfh3TaKYsABOK0ylSjuo/tMyTB/AQH/xWVsU+0
XyAbyNV2vaFkiEIr5weBPnyh0PqPLwEgsHRTZM2bU7y1MBUvMEEjSkNyj7vw
OsNqXDknkMY7EOMS7ZS1p7Ym2Uo5dv1m8YX36SUA93UPHwtDrvSVX9WBz2k8
AvZhXe/VZQpNiIq7nAa9kjreXJZWv+fHtLBrxRNFX5BgovvJX3HiRO8LsIK0
HPL637A3sUnM9HvZHBdiO11paQYasOV1PcGrSbipW9oO749fXmZjhyNoSyfo
9lKpaE2IIyL+c4IQZFIdCyjOyeYk9vtfWD0HoSzoJmGyr0c4WIkPdBHvXPUj
4sKy3V9fz5ohR5JjjZYW9S2YBZ6c7UP9wlY5hR1aOpE+7qHUqN9eOEd/CXTK
M+1YdsIs3un33ekMmHy1ISenqsbadAa7U9vf6uUQcXcf5NJGVkxNwHKkqn10
gEGjLYSARD/bxyX2gV47lIyE0oMTozSebeifHtBVqBhb7Kh6Jtzz2nElfBx4
TUPdw7llEmHUpo0uMLZU9au14pqkoaxgdAA/3zvsagbJ3CE3Fu5ykvKxXyt8
HlaWd9dWH09Nkn9D19jpZR2gtoedvuYN2tO14ADV3pPNMb/CY/Xurtq51n2n
lYknh1RgHTOqHVvqC037WxNqvjs7m3UhadLgB6U5AO0hOyNAA34i2e1kUP5o
F8kqxobT5EvttMURAOw9S1yjBwFXd9bFmbcjCpoRTOX3oh6ZV3sHuLLKJl0c
q4eiYWoFuz9SX80FJKMErn5Wtsbl5qRnZPSlqjM0BwwUnAeC/goL2DR0FPAD
+NCeKWpaCcgM/bU5j16W4mQrZM+7Me7KoMfARfBMDGEggjN4i8vV7DMasB8C
P0mzz4WZe09812XMSYgjSjtoCUnm6Q5zEFePg8QagLkVf/p9O7VGq+xdaLJM
7SjWfvzKz/ZOHovGGakXmJ5Mrp9Bl/xcJvBbVwVAVVRGqqP5FCu4CRH6beGk
TWBRm9TIH4m47UohYUfBSryUIB+6Wy4HQipto8YDEyG2g7oX8egx5o0kOvWb
ZGwgcFJJUnsB2CmS04Ben7BjVCD37xqUSPx5+OgKgwZ9myo0/WJqa64Ix6TU
DDbZcAApqS8YOpUHTojLB8zTlGKxlcXVcD8BrF7a8pDS+y7/VN8rwlvqRtu2
L8x+lfC1vgw7ogzt7VpvLwhy5M1cwz4X2yU/oHHbkfCDNQDqtUF6A9SFXiz/
DJul30y9Ff7XANcg9AMXhpGKwy/lNzNRdOrOnZEu1CV3nMkePsAEAWh7OLFK
UvJ5tGpDBsiQewAkhI4/1TwLx4Hsg4TpM3q7t9dR3MNIBc8Iv0d2nKjWwjaP
Para9nXRpTqeXGZqAvu5x8r70+us8iVfGsfWoWjxkLyhVbkhreqVDthYw+Kf
0+kvprzdxBV5CGD0ZWcSz8uJpmr/yV1p1sYOirdypfgYwEZpst6N1TlwNAfQ
z0KLiF981RU+NoDx75fRC786+ehjVUQe9kbIE/+OoUOoXkZ16a73NPuWW88a
1gDTf+DtBnTE2Z5RTyfIQGoq+4LtXxZHFNueaPLoqDBtnXYY38iUrEOn01Yd
8eqyfsdD/lW4dGE3mallJHCOfcT7FQfD8VCLJ/yoLwM9jjcUqqnhjlu2W/AA
4qMKyHjbR1ACvRew+Nn2oUIrdU6Zxr052uWMLCXcIXs7qY8mnKsk9eDMNWqM
pcUYVfLZl54yQeyTaqRBW57VwGS/QokOkbS5ChabBDkyWPjMMRG2tETdvScH
YQ+qYcv8cbE0eJ1RBVTfcCvWzR/59CLKVbP0NC2uYH2HNuZE4EmD40Xoxqdj
lww8UIZi9asZoM9Jp98MN6NAAar8eQVzX+C5V8rgWa8/CxDV2y9ahP/QwBPe
YhN0l0ToQ6DAenqrQFDXmWvANVumC4o+vUcq6CIc5qQAex6vh3Z5J/v14lkj
GrWDs2br9EM9tzP39wM9fKEnh0oBe1AlUsPH9sAPOCtmA771AxzV/aQnv4D8
42/s/mSDqaza4VkDrQ+YoJsz5mT/72xpqvBhk32xRtrjyUXEEMs4plzjob7t
TrwIh4GML6xQPwQlYid7pIXN5LM8Kz0W2eiGe4UW2ro5MRsLHwa+CEaAwvNF
JnaPWHaF4zjHzjiWF1vsVKT60o4+5l5rBfYvnR1PrQcK+An4rM4miXUqrA5u
H+Wa+e9IdXzjzwjQqx+G3Njs3z3r6+U+E/uViGGD1P6f9p18/dskQaP89yj6
3nlbsxn+VffWUqB7V2KfLheNzI9b4YcgO9+vOnYR+m6g0hPK9YiG3wcStgey
+RzyFPjBhWoBEZKnzZNk/YZQxC/ikNjryoov0qBxrA5R3bTnc3zW7wMe3FL3
rkSefcA3n0+tcjPuhU4RvY5w5zNyqPGZbW4ZpWVuwlnHesu7GhpZPh1nSXOA
j6lkBd0yY0j6nnDfrKcmpioLPp2SyXrS2XFEYgzsfRVkYR8tT2B+7ehKD1Et
e0gKifgYHh0SxRCSvNGuAIMgbPW6Ms4t25yIwwStymweFrQwRQWBG8HEKDe/
MPiqoVazo+htqYIDMX3bHMdMHKhaH7UiBo+xqhCNtzfGZ9G8CQZc5vAsP0za
r3VzDET8zcSEChuwPglvY2jUkecYMC49hQReWe8Rohue/DEqyUWNWOcIE2bU
w+1889wSUgo/45EbRbFRzet86BlJCAmRiD7snCCO8q4lklYFgpAX3oxG82Gr
AZmdk0QhujpHdDQHmE8l4gxIRTkRhuwK+t0kZL83CF4aueqMgXRYzeCbEis0
h/f0oyXrlCnTyRQJ1+eDrFrEwysU2l56/CN316Tucr0YOx7KxmpTSM0bjhbZ
RFdEBEg2nHPBDBD0rLyKulI1fDIbScjTAFO2beHCbZVv6IBS0ttiCIT09809
nElyIHcG2A1sCNkUgWhfYq6oYc4+ECm4qTlVvNWauizhkhYDj4cKhCCA6E4H
T/9cmtp6NM3ZmId9vQ6uas9ubecrlEbH5qgRKit9NMYDktAB6M/Weplj4yNk
JKyEXr3POf1t05p0Pykw8hFysKfCWOBHns+cxL4kF08bB9pzP1dY446KKSZ6
78/8mwnECwVgnK0Qq5NxYz/zu33lrs912DqUaMbG0pSRxg8YJmvpY0V8Lzut
6hmExAchQnC+bUCQpEC9nkYXL92lkCEhxwU7mURhJvofztCq5rdIu3MM4PCd
ya9rCMw/3qfTttP2lM2/zSKjwrPKFdEoqF8KnvkWnE5nDHyLNpzX3REMosDF
f+QznH5NjMfwJYHLVtO4cksZ9Y4Fc2GiSsn0MDdK2eTVHERTgY1CiNGQA7n9
FOGb1J12qvAfcz3c21HtdUq99PA0nq1ud1nJChpUuLaE+vcmzfq0Zgh7c1u0
4N7yLpzISRHIgmmn5JmP01Mg+kTbdVsCEcxk1Z/9DRX2Iz+IatKPryBGUyyT
ODuPUSF2jdMrWfesqMv4W6G8/6KGG/2ecjJkG/FG0Q22/rlE24yn/SHg3aEf
O200kNiT29Al6kWa00krJW7Y7HCB9fYYSxr1DHA7EwH0qD1WIBOLe1LACVAc
ut2vZNgwZT2oK8D+nn4zvhkwjOWiKTgtGMMie3DHY6BUNssG+xK/IfkoVdUU
Ie5aiK77k879WYww2GNpfDDXLVT/zE8NHs9t73FEL1jc8lteHk+Rzf+7eu8O
GF+qS0Kh91U66AGNrIkYDd6BNigbwsTg4h0yFF7Hoki1DjzghOzPh2TLINxo
XNcfuJ3w7vG3HM1nSIO2tjunGympfCt5H6dsNl//Qo2os4/5EfB/e4JCSjnY
7b8RJzfXCtd7ZLJWFcQMFbI96X5wLaO5qSGNLiISpgn6YUvDlQe2K819luSb
eAXVppdZhtiSrJhuidhZXdKZQtqOun9JPkD/lEb8UBENNLNAMdo1rGad0qhP
Bw5UV/hXa8l5p4mt5QAGhibYdLiVzOZ3tQUpkroBhph8H8v/6OHXOAgFxtlR
S+UuVauDuDXd0lkYH9T2C7hoMl3sgAmm0VyyTR0bBDRokdoBFiqN22KD8sGu
ISKSgxoF4YMGKfIeL/28u9QCan1ACbn726zI/pKvuup2kuz1MfpGb0XdAsBl
1/mpTlUR7DGRX+YnWhQp7vZDUg6scEwuk0FmqFZk7vUWil0l9Io7hbcLAeJI
Gzv4JrZKDtg9VvPwGrnhHy3He2s+5rqeaK3x9NfNWwJ/V1Nf5NBIeULQ/RFL
+otU52cq0dBpoVzwBb43s6mEK/85K9IewwYL4TnguKWv6CtG2qCPzrozvD8n
qGCVMQdXk4Jph2LmDvzc0OWLH26/1/0pYKwXq3KHHiaCf5tE58VjSI+Iut7p
5+C8aKnB1Yyp7gXWFu8zkYuMt22g6tLWker25Nc7P+1TB1vE5Nhvmb9j+AbA
afLNi+lFsU4ESH9d0NhHZqbpmQxh1kvPW6WEXygKWJ44qCb9oJ4ym1DcTA8V
oc/qaoPITlq/ygRaqMK7I5nC2ysMQNiw7nI0eF1oe0H7yKqNhSxKeSa0u00H
/Vr9XgFPYLvz8mQriwcb6pseQyV6tdnTbkebjT7/mw7Nr/w5g/sNGnZrE5QC
uH0Ddg2gngeTMDpNu1nnzSoj9ccfN5ejAz/N/YfzpB4fc08JtMXxMTCB/YPJ
1itJxcrhGTqKylHTSPKDWgAc8cF/CWUbtfd1oF0/Q4r87jlSCGcOw3v8N15b
KdCQ3eaxwj2kJ3U8LlmQixtiPzmYg9hVqm16d9Vk4LER/NOg8MrLCgFNm4zh
8C+rCuIWswCMYF+ntsDRBJdh5sjcSvQOaMh1UeR0q/BUmqZosONB55njw8zk
k0/jwV+zK9MXR7+eUiDe+vF6/cmsf+zdh6QUqj2Z4LbgcnkYeyN+ZBdyu1Wl
mKUw9Mlc5nAC6/azI+oElhlfwXt+XXnS0e4586uEOAsTljUXyT3YK61Q16P/
0Ee5KtmpAYO2SPgkqDAXtuCftqeQuJ5uKPwoncr2iwfbCJmVg9Fr5SCQKVIR
a9z5H8h8RYB8TlSKvFa4KaS49rweyIijyR3h86j7PjHaQQTf9C696jPZr0yq
Yt09aFxirwUb3OTh3hlJOdYMEq8kUiFBWgfWgnI9PQXboFlY2QiYEiP1XJnm
vll5EAeaunPFvvC5UYmdFM3tAkygs9y05stc3/0oHSVl4pK6Jm96C4poQPYW
63+CsFKrMtV4xzwhlEqnFykWiC82yrylRNyNUpRrEvQHJlHugh1S4fbpnj5k
n1In9xoVfUdYQvJ9APUCBPQj/DomeseC6auTTLms4N8KZ7aqIhBAyAqPjKW1
A/n5YEZm19fs5M9ZHZK0FBb2xvLhTWSH5J2Z0VYc0iQBLeQBALqZhWH+1zE4
/6iBEDbiOaIULaq3mPPMtdeVWR3r/LlME0VTLvCoy7GUtxq9U+IwY5Cgx45j
kTiSRxOUCYxr+2jIFoBZgdNk6q7uPW90vYJSxnH7swiuF2mG5mYsE3lJ48Oa
icKu9hLvZvOiLaZpctqaOJCrPhlYzkZ68enHHYqQfRFnvFNDAdJg5dNge92q
sjSkbahvLL4BviLzVxTvZ6lW0j3ND2RXSOV76nADAufOxKKaSxqcoYAqKdS5
vtOhIjsNsU+53THnTxstvuP6pojQ2mqqe+8NYdnnt3My9trTbFZg3Fpc7Rif
npq5uGvIR0nSroWo9SsAzS0s3Sv7LYYRVkm7X7wHe5xEbE3Z7+GliN7aqUMd
EiLQr50ZgYjMyjONO5+TpQxl90K0iTj5pYT8zPcFn3EwIvS9Og1uLoroTyHt
+fDvFw1Q620Ljn8m0/COkfAtIiPTWoANv+nClo1z1yvUb/ht4J6Tnvx0ZTIB
0RdNgj2ZOlKMDoipL+uf9cLH2z4eXGBZxaQavBakbQEmKZmPv9A0PEBcCOBV
+7zyeUhwx1GiDwgM4PlKBz+toRm0md3XQyyy+RjOAwo3CjwZ2wDEn0BGDCPA
bvdm77aEmPPvDyvAaiovU927T1iCwJRvlBVQSwq+hrf0UJ0HNQOh6Ka+M6Qz
APXb/zu78rvTQNER0IVE63kxgRZxfYaywd9no82Ju0eFILzS2u+TN86OtEE+
SGk4J1BPbuZw0WsinxWwQ0dgdXlHDBD8ip0uMry7b/3p/IMF3b6XObBrmwj2
MalwiELE89fulj+RfcJPl3MXL6gKMuiuM0RTc5Fac5jurQC8Z7FJJ8Aodfxn
CbdaPRvhZXcIY13ucWFL6KzErV3tisqplunqUhp4s7MsYt0v4qt12GSVXbJP
oPZt+lbobFyEOK5ia+wGhd+Gwvm5gg2TKfGyeMdO/406teuhJYBuGIBhxHIO
wTzvRUXJD3cszCLqomM8E3t48lz5xATYxDQGoqtIw3ciwxZfmPfQC8GaT6KG
HJjgPZ0jtJjFYpojtbXyN/tVKNlv1ynq3RNOANV1/C+xaZCAp9fhI/b6e9Kw
ax7GFHzm1pDNosO19pv+sMELycMdQJjpYcATMpVomvYjqOOwpcpJfyG4XesM
6CkooDo4utAtUuUlQP7DVcmHwysb+b2HTitfMPVSi5WlbVK4dbQn9DJ8sMUB
xbMKIE8PO7an9L5iYS4HxkxMvdgCFaNNkxOat0oc7NxjnHleCVdokdHf08LX
GcvDdCljspEeuMRgZ5ZzzUVYvT3HAHWd8+DE6LE3cw/Xl4qZonddVAGpj3uP
UvLXvD5IHefhv3mIDnuWb4wvlAHlL9FQJWgFRTh8ALS0a68lVLfJx33zy1iZ
kjd6RcIT22Xj/+w5EUgDCI+fjsmcvoG988W1T73zKaiY4LIRUVLrpiMGOr95
eAjQr2XksueLfTkuNPnhOIKztHfUIPPQbvNGNjMH3LpzY7UPH79s0/8zgzEa
8g7TEDgtsR5TNGL4FC2e2q9RgPZcUm0COc0aHIQyxPxDC3t6ZRUkh1p9uzAH
TYqh6Y7D9tGNzN5n2HrUTxLy+CQ+HMHYo1LWHnBiJbS/3nMf2jxZjmUoabhU
iqH8bH75JUwpU221wemLZolDQJ3hfeUO3kB7NlAMTDK64GDUOqZqblkJoJZg
Cxhj3FSXYGy+m59EzS1sPRSlAqLfkLynDt69//XHFCzlyjN64uZ3c7WNbCIX
k5C1L2oTsAHir2eOZXRPSbLG9g3omz9pg3qdTvM+2xmKDlff+P/5dClCj1CH
ZceA0h+dTqr/zAJ9ezkQVCT3K20Ydel0yZDf3rG3KRiAhau2wrkYvi3hsLWp
x20ESCLpSWnODuEQ/zAUMB29x0TO/8du6l/UzLufEnG1bBSHIT+kYtj+LiTU
clZ/ELB8c0e5Fmr7pqRJyw/g3gB7ljqMQrQ6Ls5OmIE0RR0i4MxqbAQ+8Ehy
tJ6y9TcYcarct8MyIBxzqKUnQw3kO9kixldBPdSwOizH6Ir40+UpBphzSrwd
IYmegtFhqHYGuE13P0YHhGqHrPwd0EkX/QJwHhRUqHBxuGJytqqXP9IsBhTP
0EsDsQd7Td4aDB1nlHjsWM91dx3qKFnbBsnI2ivgXC9ujMZwrqhaI3OtoIwg
hAOVxy6lCcCRXb/Y7p/4KO4OfC5eHVpeyEiJf7RbbCnS/CtSb255n/Kgvohg
NplAtAaxYmbrxQ6hzH/rucmBR7H0JeWqmtix8fRfSaprYoeNNZ0cWgYzXA29
rendvYXIvPZEwDBBZYctHKYqSfXwtw9ybKAHbd9wpocII8Q4QtMbbI+iiEf4
qRlbnBPYFZLAdS8iklML75X3G90FOBXfUSJxq4WKjxUbAf92MEjhH4zWHOX9
9yD9V3SI0jn8V0RmhAlwQCPpFsXrd1bvN1PdqhyOziXR9KfAUUFWR07mePKK
o9XYPwnwtoqoQCd+TPzeB6lgyyhqKDpgjObgFfJpqtynxNO0Rf1haeEQ2f9J
jEss6fLpbySqOVDzvQy5GY9qUK+2MmXLQIhFOtqqHZGFfS/AgmJnZKj/rZgM
RUMzMLOGH03jT0X1sbSF/gsLJ8K9H/jQF+KP6hPuH1dfjBgGz92v0AocAmaQ
ndSkMaVnk3L3VCE0ko6aqcFHPrBjeZqOEedTNPEOidhYQZ7tH6qzsY5mddxy
6zC/cavR5N3WG/Ug7QTJ5AjYben0mLjiTbIxqUMb89nTfcYnxXLUc+xA9bLT
dKoeG4tLO7s43EA9Kg4ftJEabmjq1UWC3vv/Lk0L2or70P+KB+XmqDL2AQDq
zLuVq6PvSHR1DbIlZ6aepRAyyRXohrv9QMKOJsD2T4zIIY/UzKZe7p0DyjB5
T1HFf/HHjk6pbJThQ4RxR5xUpw888g0yKSMWLOTRJSugZzWRFGVuihRA63ER
8642l6SEWYP6s/FaI8AaWqGWIbJJaK0Yb+gMelxb1Ar0QfUKpjigFxtgrvQ0
4gUDRC8OUl/YsPgTX1iVB0i9oS4aLgeCtVDDceAA+a4GXE4o3QDVRdRH4333
NnSfBL7x9CkCW9eFZyd29VpgLEzpTG30kZbgjMHwFFMLsbPpvN6Lnj7R8vcR
iCbbvPLVYDRybh4Fqo9f6E/41S1Om2gbc3yhFlU1rkGlk9Jq5mrsAY3S9Vuk
JjnXr92V+X/3EROFl8gQqqjTTm7AbcZ12h4bBWmGFRtc5zw7amIxcI06pO7y
9K+fGjsUEL/T1I7GrriT/UeE2ecNWZ583gK2e+HHDQSpSrOkpAYdfSb/XsSF
A0N4BjavQ8gaU1oxN9Spu8kHXOitEarUtJAEdhKtRvyFHoHbQQakeXyM1x2u
jmkzvsLxhYwiKEoPjl5XHN8I83JLh9GxLW/UbHRM2I8CKbnZAIDplLceNeRH
UW7lVWyof3uK7SZWAvxmMWlHYA7lMobkWOkmo/GoA2uyfDzDZUC7IwO/xKGf
XOPY1BzdPvHBAREuLha425P1w+eRnMdpFwrxUaPhmy0W18d0OcO+4ve+mfyD
GXOc4FXeExS6riraW6QnQP96lvrRZZgRcwq33hiUmfjUZLzCUt1rByD9GEdj
G0Beyxn92TUT2O7IV0Zy3wcjqzrG2JPH5vqH3gFO5DknnQKMlRly7HI0GFVe
q/UZbfHi6D7HQKKo4ZRnaqaTxilakcMDTnhF5vF7FQtw8ymLndAP0RMP0SGy
9dpzB00M3oDETGnXuppWadMxwI8bK3ZEhosE58o1ac0h40caxyQgRx+ENV80
fK2NE+57eo7W1VjrwZRf9M+sM+GKRUByAwIF6FSOgubi2w5w30ySupmsYzFc
rrE4mggy7+X+x0nqvbQW6/rR3KBGwZMY385I0ulDyXRy6GsZh054OQAwqHw9
cFcYPzbqSaJWCNHB9u9d+UxqxQuXvLyRDSZhAKFC9D1E3cj+E3vupHrUY2r2
2oFgzsbKPN+EYHdHyJSCJy5GTBRW29DLJ2imrBZlm0vKD2nH1yP7g9MhoFGd
w3snwoIzLgYYyxe57yR1/V34euVtIQ5mqHAJ27KvDURPRYNe2f1OzxyRmHz4
ZWaiLqnCe1UcQqnEnFeZy6IQCUPYivGQ0/1FqhbVt6Cbjws1I5ZbklCzhATt
55OLIONMIbkMrj5OGeNtltBgeOofjwkaM7SIpwVzAeDaS2KlDLuLBmGt8McA
1g44uVSi2siUI7Ylu5aFDjeKj/NWrymDlJcZz1KOnvLulb6yZMmQAGOghOif
HwYpmK9nLuMJEqNW+Hq250C14kpOFR/XrTumJaAxiTZlXMOAuO5SgoG0EAlk
eDP8iChB3u45wHnGGoSqnOcasyxOYkvDO7iMjaLk2V1embmx6TKyS/UVX++J
DAozV/RJcoDZvrW4Wk4RXqdxiWnFmrQLHngC6EehVMcqMClqwWZhwmbRGb3d
2X//aN2mZ1hnTkxi8pQH0giogmXSRZB0DgAnvLu2wS94jueJHD5OHymy4GHm
ZP9xdx2xyjIGtl+8ACsFKemdKClaqh3FDp+VzOw+T1GVDLL+VgcXICSIZKlm
RTRsSd3TleblBaKdhSL6UkolMCPeJyxnbkVSsxlWDYfJtMUHSfoJI9fQauDA
r/+ClblWA4yld7EvyjpRJEA+1qmCfE/IhjyWPC0zjpzW6e7tI77869c70+c1
FhjEO7yhIjNF67CVJ17w8+CcHvwLCTFtT+kqHNud8gELMDxN+IdTp7m1RyXI
XSVCWECAFy9jzqCaOMJX/jsqTIQ9V5tagNJLjFnztIUHfnExzt0i7rtdKZqe
n/9eCICpafUJ1yJcPStV0tLeFsh4Qqmy4PfWFzImnB58YJQ9OJk2WUetCPXu
s2Mgqv8Ld9nF1cmmIxV0pcBBldjqzYrzZ1y2VMTQ1WoQUWcnfKdUfgSD4jnl
qcG1s0gKwCCrKBHZ+HaHuf2DCjS5QXgrkDEXe4y4EEcyKopqgCeZ5etfqhvQ
4SOHiCBMQhOMSF6PNQPj8f8s8a8vZLKmZ53mhp2JbVHGcJqkzs2qvVGP/DaE
UtI0Mtq2J2cdHaPZxU4MmuJMYhXJZuqxuWU7Ib/DnoVzc2ydEBK5LHf3jEg/
/VsfJmXz4vC3vsSmsqttumhNkZbpLQ/zdU7sSDJXWYULPeBUDG8eK3KJhZq8
z4zpUh1THO5LgdmlqSxUfDGI99Ms3S39L7Cf5yalTqFxNwLJ6t0e9AquPH2P
3ia/MY6QCP/IsRS6/OzYfO230stbpeVTrk3NqZICzehVXUZbfoMK5GgWA0Z9
eQeuUvPb9ua/L4d6HBtow5wehHHuBWmfcUWY3EvQ/FdtwdTUBqRaHpBGQ6VF
gxq+R5iNtNsyTf8iVsnvd24C6Dx1TtYEShO72o/krAv2wmXXjiMuxfXGVCQe
C0bL5MhtxXHszGWLfCOUaDwapWKEIjEPNoa70FzQP9gz+ASl2LuDoveyssAO
D+F5oL0ee6aDQcGjNkRWyGil+PJ+Z9jVHfGfQRN7xVGQnfxy10+h0nRW+ZDZ
lNr14r+FSVJ9Ty6MeNl+ZYt/Bc09F1t4FZMPiOpNPdF9X+XtUzlotdsFxq5b
yjH+1X6vjyuckaI5nh1epAufd/PjnzJJ0Yd7eh3twoq4vQQJcoVfA0MwV9K1
PLAxgSXRmeNdgwVrdPiaNTsr4Q6aQJkgQOa6Xaku0IFzwzHhXYmbme+FLGT7
Dd0hO9VHHMaKeQyZpmP7D6YXep4w6RK9QYPNkwnsdqgVOF0B+3RF9ztKjieY
VnOeFPrwHxcbyVjXkD1H40GFh4mZDsa5e/KDcNBafFBpvqg9iVhuEzbZxMaL
4eBG1GFuSGM7f8FPXjMEUC6X7G+unB/+Ypmc14UksgJHpT3f+a6Ez27rWQyx
iXeRzZWQ/JttAPM1/4EzSNyBAxU3mH62lt1InSSmNR+K9Mb8dJJpysokFaXS
rLbBhqfM2TdJpAU5SCojPMcPs2A8ldpyQ8QaHr8EC/ckAUry6S73JFC/bFbJ
OI0PRGaPyvi0J3RC7zmOd/NN4afRe9Z/dmjew2OdHUYfWWsjpxIbs5VVWAaJ
/5OQ6tRaXHNMJYCotZUmEboIXB21XvXIiD0pTGUddV+uaRudV6OKSSRHI1wj
rkJfXh+9eVkkI14UoxdZoEMpYq6K+oPXfXYl4UmWbt6FyuPy31vam/jyA9uI
M62XQNfy3aXayYRLcndaYrIBNFjLE0vCuTvAU1a3CaDmfSz1JF/Mg2DyIdVQ
L5rkimm59xNOVgIHpyOyz1S7Radceeocshx33vCzqJgu7BGZM0ydLfuGX5R9
5schv4tPq8wMt0q7LnkpR/Q1K/hD8Ut1vrLThaIw6ImuTWRCqsmkI4WhlJy5
u1jZ7saihl3E80I1ActFotWxcz00xX4eS4lefxMRHsvRONB2Ats/20FgrYio
ZCGPcBKskREOKZd9a67KJ0QGqtpjoW7hGIpvOVrLcEjMUBVnoMKpo7u+cLjy
k2A+qruoWY8V0ov0UCdajbK82BUIRVbJV/dswhcOue31Y6a3ktKt6qkoxrJx
JLbJYL+Q9a5BXM8UYzIbbK5Bb33d3CsLPkBr/bdds3VbAcK8mfgoIjFhMc59
vyvyqLlbM2qWuqSphRfXEFjpFMSGW2mo37XMg5xix3Uzxig9kd8qunRLiEFj
zXHZtvs+hhVdkNY2S4V1TRGo5TvyHx1+471hi/bfoQOztfxCKb6yyF2DFi5J
wEOqI9Hky5ho5YP8HhkSib6cJsIdTTGtL8Y6LjtrOGqNGZH9LMuZgc23Vkxg
GfH9a/0mtltMzP2g1c6gd9AF12o7k+ZeYXtvCEmUju7NUGuEWltZeLDqWnGO
uiF0ic9WxJ5jLcgCXjRB/K2pjinv4BQwD74EedZNaGC0O1FRJXNyV+YEsMr5
ZszULFCG3P9mJOxn8lFAgVabi8zPiVlmfO3BXKkDfajgHNYUpxH3MxeA3uAu
GViB32HWfdGDOAgdkyG2CXxxeP1p+81M9ofGE5YYsl90ELVNHtoXW+PLpiiR
X5PKlBlLwa9eamhJ4/XWYtzs3NHyOu9FNUAzIKpMZxdiCjH2QG73KcQcZOiZ
/Xa0HMpe3+gg08nP4KrOtS7Eoy1gJFi981QpKyut59Qn1eYxltFvkNmgmncI
Y+9F7pUr32NpQo5SX74jYd1O4iyZs8NrXq628LQ9oEVgXgIcDOkUyDuu7+T2
cdTwIpdODKU0NM2OVNr9dlD9OIoCgnJNu4pNWzdRd3LBS0y5ODljcBAYg0fi
U8gabRSN2LPrTTDXAUCquwsup3PGWHXytVgnylBLU6Nq2dHL68p001VS0gdy
vvjichIVFQPD2/s/LzCL3W/RYyia97zGHP8upkaCOuzR/2CKbNV3lLwEK/gn
8XJjlSOUZT2gFUkdNt1vcO4kLRN8BqG3etsIwYJzHVtZTkMlu6UOLqnAk796
i1aQRCC+A5nJ2+B9H1mynVRzKDt/2BTC+wsDcpIPSNBZ5eQg/y0TZ3C66cN7
fYy8/XJDzwUCRZTYCARnnU0dXUHE5IB1qiCsYYD0ct4tw0UiLFM2AtFGs6yN
eEZ1keEVl5AuL2B7+RkITcKvVzWiS5tZR8SS3wG47HiNhwrXNrHJzgZVW/4k
IctDqvPn+3lJmLH6i6NEZXCpzJS7J9eCpPSHW5FO1sX7RvPTYe1Au+OaO8No
NB+tQKMexBoeGzAN7JuYCI6tVFzmfEVrANQXY53vWvKT/G4oUbtedlIzc9UT
oYfi5xRfFGAkkRDgy78mw1FOdjilDqYej5KwEyK+EA9R8iWIDGl1PSppp3tL
sEE7tUY8LjysXCmh3tXSICGD0vhXgSdY70wdMvzxyxz87sfB85EJlCUtWlLM
QXYlYfrvgKoiP6XOgz1XvbDMJFJ/KbvsDCcafUnXEUeROKUbLzXGEk/CSCDz
H96boKI4RqwXEElFHYa9ke1SQFGFRKPVw5iOMi+ivc69FXkABk39JEsoeQCe
ugK3Ea+IDAU5zNpP26dqfKbGY5SlSUduq4Mn//ueZ5QXOk1fQ9Mj6rrLu7vv
uXdxrMu1Nes5q6enkkqYaNfJCBfgFrcf8gig7ZCSeqRB6AwMp6ZiN3/pmCW1
1pdsm1x2b3GkJLB63+PQ1uRZOah50D68XZc/DPLK9qKG7ws1aN2LVLEe6Bci
gOJgH+0ubSLnoBc9KUexYFYwh8t0DPzmlSG7A0Te7o1BTL7R5LrzhXMhJD9N
pwWVr0Tj15/zZTx8LduRHjDOiAzC7tSE2Bo05oDj3qRibbIgw587lNeRvJga
9M4svk2zqM/f3WsFc6ijUyrngBjWbVAOMrpvIvM38JR5ZM/YJv04o7RRNLBP
VF50sGz3fb9MizZvtLTY/ZoLydRJgf0Ppa6k8lDIHIQebbEkLpmcNXD71FGr
pzBN8mZRY2VraVOR2KmEji2aBiQQg3ZPQftqBQ4sXjDHrAfqDsmBvzir/bgf
2qZRnCD5qIOgucB+sHXyCYUMM8jPHASX1n9jCWjUIeAUtHc2HA6CTkg9+SNs
lyDTwCIwTvv6lpb66MFZNtBHw/bjRjc3FicrmHFiXeRNuwyl5Av4D8viQLn+
S9795zwEYRRczLKHIU+l82EOesRTvanRlP1Imn6O9I3bksDhj1Z3/M/2HpTP
5GYQT/lqzg7VKHuWvgAsdtcihXETShbj4iTswrPYpx3deIuI+RtVhh9ydjR4
DzWAe1sMnyut0NawGg+RkQaZ6vPpyZQLjsK7rM6O/jJPjhHt0ENeEaAnVr0n
2NxHEkY2pmq/ejPd+KV9g+FORbsx82rBfKljZKFeXd/LWIZTzfAaM5hJpiJ0
E+be7BvVm7tSMCn7suZMD0ttno9ZrQuXr0LhEaZVT+clcJQIrMU7ksYi/83d
zSEyxAgClvRTn8p5eWzVfaJiNbs85wj/uzyLyF9eGupTjBDkurKGzZnu1a3s
89rzRV0RzINNjKQ2d3Inr7c+OcXXLhl/zEYs015Qh8zT88kzYCrUT4UPt4kO
r6EZ0HC74WjusX/c7EB8MmZQ/gYfU7/OvOsMXSk/QxBXh/ehgNtGhN/g4Jq/
oZwCtntevJs4w9603FCfS1d6HjK14YeLz2WHrlzkkLd1p7/dqSWkbMWB4WHV
NSYXFIV5yhfvDk0UzpA709vAs+oG+K5YVgLZqlQYFwbHREz58ld/QMXxeBNh
sbeL/tzWbPvLVddbtdlMNsZqP/aRRlZ5lV99+Vi8oph3hNOqpAud2yBmG4Dy
NEZzrGB+/RiTXsdRtbhggCaIDMD8XMs3QjbE2D3tCNuONn0ZOuPBHhcxdAtV
xE13/g0pzZJkN7JxCxm44bdAuY5b9nUINVcV7xpvPVZ6f/TMMsnzUkUXt7Q1
wLxsAsiYbFcI6AYbTNoih7XmDRpNv8knCdVNkTqWj1XmKAW4nAzYMLf11nFN
ErzA1ap5H4dBlZ70KYrRczrBN/gK38exONRHzvckwIbcXoCgYGYLGh1r1lyi
GG+Jbo4hIIiVhMlPOzDo5SyEk1Ms2uE8wY4Bre0OPTjf4m34d+tMXLlBUHmV
NiQ+94P65ie3+xq3swBnO8z009pF0Bg7LOgfwQcY3HhLvymWhuHyDjvnWrwV
bRCE2+O4P7HgemU9gxhD087s7t+lDb6/+bEY8eYEKWY5Cqi30rrF60AN+6b/
IlpR8txFR1Cl5wawHlICtFtFtykwzgLW7Ek39P9LLIw/LfnNpFOgWI6YmRPJ
vdfD0MkdWT0fx7wGVoA7qe/HeST7K6Y3zYNcnDMHxWRPOpZ5RoSMam6TWoGQ
mPm0XH830OYap50xWpB2max9DuopjeCGLSwZpiRx0hKxu487aHola1wv/7pE
Dkv6I2S4eEa/V/Hrr9uSwuLYZfcjFzxqCZx41AE5t8qcUfDhTrS6P/lqL2lj
NTZTFlOxojwXy1N3pR3HbX9lqUSE+0Rz53x84CBH/T81mRCpmJHbsutIp7/V
pOTQpFtgTrMWkHBtQ0RqmR86aL96SIJdZ0GqmlQOLGroMfSbp1/SxJDwWowt
wQ2+SjwhpMm5UF/H2fzCelWjoH1++00U3uVStvngnUk0qV6vPzOlrlqv7iGV
KBqntj7nCE7ojFajpGQzemLD9WOHgoDsGVizKiYv4l6Ntn2sWYMTEbeU8+rt
UyBojCYl3U39PY8lbll4ASzkSrIFc5elmvg4Bo5tkf3O6HCJ7MlJouETN8+o
qoVa91DH1rewY/jjoH+CuhLkfRr/LjoEZaxsQJ+5cZmmwbvvgrKNad6t6JdH
sw4BKJBGyqmIySmgH49z2jOkZs3qafv9onBpQv1STDYMU3KE6w8LZkIzYssy
rrG2Ol3EzdZE20XEUmGdG77qsymdAXi/4U18kP1A1gjubL6tLApShZRRMvpo
nYrHA/+DH6MvRlempi49Jsmq61/teSu+l4Tr0yS0wt45VDzHPfe4xtOLQIYz
UZ8URzLhxQsaGSF07oLK+MpuM3e0vdxxVQI8vBaQr4rT0FBioGOKXkpLgIOF
DQ4CH4SEcP8yKcM6hKZXHZb1IKfOzn7Q3bqMZPg4OIzxBH4rJLXJn5aoChaT
tj6xYaD3ILLiG4EfpmEdNIKKj1otnwCqIDsGX9TuuWj9JJqH2FobsjdMLu69
97IID8YE5ahECMlKYtOPY0Zzkwr/JY64vU2zrSUjobBai4n1jC05UxXFx95g
opPOSvKzj5Kw5JZge90B9QzRwz1uHCn5FH7J82DVdbfX8WzQZNPMcxQxyyQX
4zCQVDVE+rMFSxShTL3FKqcDNSk1b2CqhRZ1nsU60j7Z51Yq8+dVGSPizKZU
Q+ofQM10jNNwJGmydZ0lCROpwuysNkdYMSy3zX2mrdlmDzlqZEKueIIBoEIC
PEtcqpilqZnismw3F1nEaG9z5tlqxKQ+fCcA8qlu+I6m/wau9DfPxCYl6tnB
sgeKnNXFqrxRRMs75dqwvZgf6ZiFbev7kv4Cp5oEBZ0lBJcsWiioTbpyO8Op
mgn+OLuWzOgsfSTPdRlOtbEF3W1vICeIpPhbsynKh/LM0LlVuXfLOBzbmzT/
GefY56LY+irIJSL9chI5QzWKPDmjBAuZs9VLuU4XRTTfv3mCfTB1T3LSuFB8
mVoKAXfy3CqvjLg6gC6rSmYSVqK7WBC0+L5p6vWmr2CCreEfAAmk+x6L3Qew
qYILnAks5o482DiAedh3RDSEdeyZr6d5KRUuTXxN96aPginmQ+n+D9Qw+dCs
rtNtdUQJKDUrvcstoSPazzy1dlL/fAS6RD3fpHcs1Tmdr9HLBcWZKR3vhTqW
GqImprgRJsYM6wRMzPIypYTn37jF6tIehCxsnjEJNYnGiwxtHEZp/ZclNCuo
bJNXAAaV2svknNQmc2sQeysucAXRPJR4XH42uvRtVBuX9evMIdO7aO61QBvo
nUn4Gwvg16d2YiGtnoAqgmwbleKdVCfTxjraFgFaEfGO3G7onoFf/rIqRSCf
c2eUMBWxw3GxUbPpMBfKWI2Fa+K8XOQqSrzeEEDVliXczRQ8h/CvBUj4HpPf
34L2Tm+fRw2XsJUgwA4k7zuqKehQrM1Be2B77uQa8R16atDWZ4TGlao2O9ql
ftpQtUB1dU9LuobK63t8s0mp/ux+ZAIQkWrkOXE3tYT/A5Dlv7Btk4uylnys
g9x2LO+1WhAhNzdJRKWk3Zd2/MuJ2fodfwS0KwEtd01OwVQzJ59WqypsFldw
RrCBnyLiv9uTU1YF/ASC3Lws7ApKS7abASfllUjYq7XRkDYTPPjPvVn3vzCr
8zwjkg0Br0rMnqBrk8JvCzdpfY2rZDF3MjF1BTq+9PDM/Yp+U/llvgv6TPyh
lvQ+m0xATHKdRI7TK5mkzHLNv8/NE02nZmgf027af4u+A8l9udMQU+kMsN+W
7tzsA47+eXjDDs0tc5DBB2itZgbl2UvMV8Lx6DRNcKD9RKEtJLsXpE1qG0to
GJNni32qnlD98X8+9ULDQKByTDrNbuAxA8h5i+zmwtVCba4WQdkxMs63JOAD
jyQh6QSECoeZTlw6MRY7NOf3smLU4gqMEse8lRoTnZO9wR1BC30F9IqARIom
jqYX7gu+izMAx5p/PXCm41tD/HYXvWryapIVWurGRt3uYYWwYaqzFfDSF2NR
T757T5zUXh1w1DW6YynbKh0S1gKyXKjR2/S4qTRWfKsHalCsg5dUFc7jbK5Y
xZ4cFRIcPkmuuUkz13Ghvsght1FJ87MCDFBuPPqHhowRL/0qzMA317wueV7v
LhPx7qAfPnXK+Rw+xAD2hyTskHSFLuPCvjk9A0ccpkMzm3TUbRs3k+71a/FR
W3JgZklz66uf/5LtOQ6bwE0AjIF1PTIFPebnfLltQv4YNm0PnYogRVapL4W6
EMNjomYD/vwbi14Zloilx9OW3Rjhk82HEX4RBtZfqLPZi0pIT61pdFN6p7xD
707bG0Hu8W1oQc4lMBHiFc3HGGQT9YBqqj4OKQ9xm3K8eJJzWq7Phjm5EhON
1dLUZiD+ZhM8VTcEwC+OVgj38JlrQovF10SbGAPkBf5c+y6XSQmtbWtYiCY9
hMLIdSq2B7PUXpG6Wt5mxUYkSPC6UnMVjjWB/PabAlK5P/zpenO2YNQHZ54d
ajYqi64QDrWBVuJvEifk8rgyhIZkjFV9It07aSDGMY589R27+RJK0IYqsUj5
IofCldom8KrNurwH+sQEBhjVJ07d6uLMhJQ3kRV6A1/ddZI4PL4Hn9d0Y4DG
NN/MhRmMQgOBNt5Xp/dARWwnXo6/BvU+EmEr/L7S16Lye7lsVDlboNmJ2QGJ
isVrTFF65WLF3hwIMJ5d4nXRIYqg7eYarWoHWL5R/HseqdSE2JsZBy9H/+vV
XngWW7q0UajR02Ksu33S8d9zgVt+RhaqBMpw4kVAfPRKSWW4VKTuq+S3d2O5
zur6rVCzc67JT1ZFIqlFrTffXXg77ev127NOLEUb5ena8Lc3RSJrg5/F9loN
0lSvQ1SabrBCJLybHR8lmYJNpp6dJJ1UcXJV0yAiNpWMMnVVlFfbjSs0Lt7v
68IS6U0yJYccaS6Twj4ibM7xAcnswHOOFgBvx7Gu40GIkjP6Jav09h6pJUg8
TAonQWL6GngXi1OtTZWKCqDXNP0rHI3BcVhDOyOW7AoFyucRoZGQK+0WAnbI
ELt/Oisqq+EhCHrHhn9GHl8zBmegWqb04AAewpVXZp/diG8LU6Kr1X/Lk8lj
GdcNcBT+mPRTE0qJnjqXK9bQ3FzH3tI4EqcCFO4kUX5eU4qMpf3KCZf6+5yN
IsCot2UV2N0OlZqb/GB6hmRjn/DSSaYCoKwYiV5kIM5IG26BbBZqbrZ54wT9
TiltIJpxUOKNpeJgyDRd3/GwTJ2hU6XR6URcUyFFEU1AUsrFhX46hNJBYMOb
KZbJZHGezctTiXc/Rn/ELE7VnBzbSSUhsA9HRguGTrpvU24PTOcndNBT2vX7
FN86BHAkEQYk+Z3J3awnrpzNbwbAXDmaVAbLhwvMORm153Ys7qcAAyc+F6LO
EiRJkKRUr9U2vhp9Yyi39SeKFWcH/FaPyccNmETeTTgHlGZSo29Ped2klMz0
C09aPIf3WSjsKvTCT55qyXnPRyoxr2Ku9Pc3qQYF8QYG6uCELt/wAPEM5Jzi
jslK3rGOVCKVNvGwp74h5meEy7bICvb/4kvZSIpL9ESlHBbW7cxRILkaukUz
skvXusLB1OiQiuM5UWU7CYh5PS6aT55RrmxghOB6Y1yF6qygIPdkwwBfdjKP
lLw4e1VUiEYW2A1VOx3JhxjzcanyPEI4971VCszZLuISNJIBu3g1IHwfCo1R
LkGN7OU0oRyig99stPazOArFBN0Q3kcrRFrsj3UlRMMQUmNvK+mJthA3NNbS
nINOHPQyW+zca88VY7H70pr0hocFgAbKhVbrIXalrQ4gJDQ2YjRg74SG04em
XqKhdwFTnSt6aVxnYD90QoQ4NK5mE5Cga0leXJkPWTFfCoioQTpxM6AFE74k
VUGOyGj7QuoZw174Jc9URtvtz0XSQXCpwg0dLe7t9cuC7GA1eEUd1rRRYSFh
da0nRgXCSdOTwWaRXIPjHwILS8Iwttkd3BXyQXvXg/D2DR2b0aQp+hGpzGlH
z2D2BHWyo+zsQg/VFTjzsZo+EpurGyDe11ah3Sl+QsslwMH/nIvsxfBuLVz0
L7kev2ATcsb4ENGOEWQkOQ2w2u7+FY3gCEY+QCsu+02BrMqRTai16yfDHTei
cbN0f1L2h/BbvcQqgUBbflPgHZF4UzpbMDkppPhodhlXG0Hz3oh1I5yrCjmC
uwsV//KSQyMhUGp9qspppo3wO44FfbmOlmSQMbzReghE/yflWmGy/9oRSxPQ
FbVNur1UyLFDEV+e/4lrTK/t2P4c75eEETI3K3FiCDhhg9viGwhEFiPqfYu2
sD8Dt5VZdRogX6L4RnaGY9wL3KlguOGXTNtronUbYqM1AjayVMXEuCIlZYgM
Ec5kX/Sp9iC0Jq8KYSSjtbr5nb0Kuu5ywOZpSYyHtf5Y4Tgm1l0a146fzqJE
wh5wBL0wwUbx0P08tAvVYcNcHb05zWlZCj/jybHlauzrPPQ4udxfahl9pDdh
gvGjGzSNv0fUsms9NGxe4i9XfWImjihMF73RQCV1T/0CsXCEIybF9TrOi8b6
wg532sRQwO21cMkrNPIWdH85DwzVdZhkKyIwdifZRz/sCknOA9PEuI+5PBNN
uLPAic6xZDr5xgOFRcVx+x4p1LNzoMbM9WI1+bhvacTSDJsI8e9YbUPu3dnx
/BcU5T6hys93oB/yB2W0az3NMxyhoUBRN9k+zK/OxA95cZavX7nKzA+DcNsL
0w5vj/i7qgu96gEB2EXI944bi9bZmESYju8IRZ4GcpHZ2meebXSAw9Pk35wf
kk1i+IJnZIoHpNoqjgZnJQel8OURqbsYqZN1bfWBvsA+uSK6ljSqnM0PZhqu
XWDzQbHmtwfu7bgoIQH6hzVvLD5qdYOy/5n2cDrN5CNzas1pBdB5h/GJpNEC
EQEMlN49mZv0+pzysboBk+iB09PhTaf4ymtTQdWkSYNG1xYrR8KhnFVT4mNF
VeZvMvypL362xpLMAJ3Fv5SvayRAPRXfUBOWL2Mi2ZJT9y0tMUeET+I+uNfo
bM5F7UX3YBscSB9wRxO5WuWqyH1+7aXf0U4BO2g4VsyNoj1+7nbzSCqWDjdI
AcYU1MOg/KOQHlx6hBR1yVWqxtGbjyG0khtE+/SIfNJbkPGCzJUHnxWvoXRa
usrU0Hyn6iGE66CqBasjhDMOOAVUKIULtxRPF59BcMRZgYwUwTRVFxAyOuQR
6DNtYEnTx5KBAfrfYJ9rF4Xf7+xiOyARavk09mEE6H3+nn0j4adFsOKGugX8
TKcLZfqhQK9v4aaFPlWjRSgm+F5QPtQXep0YoSMeLhU3e3iUFwPf/5vsm+zY
54RKY55r2zgJvTTdxWkkj7x7LlY8FIM4oT9d7GjF8D94p9frFi0Gklp09jBC
RclupjXRD12waQeYH9z0x6ZbEXN1dfFBsJK5HyDQI2Oo/vrWVnRBmi7WzmDV
u+9SOCONyetoHanfp+8rRpvqCBow4KG2nBcCiXoibDYNqI6tQ/+FmSLG57LT
d0DpxuvTSHn58O9uRDlRRyibLgHQhELqbjzlGmkanx0BgLHjHR9VOV2BNcfD
7lbsbPKTN58w3UJ8CH0PemxOpbP9MynPpvbCYjUGtpHeFpq9fcjDIb8nII8X
I6RNQ143w8KmBKKSnluUkhU+TYQHKZ2PPz+bU7ehwyJ3Xhx4ccthfzaK8mDm
TDFAX7E6IZNz8aerws+7JVm8thY0UovxKohSPsxJ/G5Ty8Fw4J6o4VH+SQCJ
22i06+CjlL1wG865Jr76TiAGc1KLBIZ5FQLQEpz8fri2ZXJvHeAbVJU9R5c7
JmBxqAQnBMc5M/plKNI/OISCh/kvm9RMM5lmeCUUYBe42f1I6oyFBy0ip9xG
SN5jVqkYFYqQUSC2DUtpY4TUX+LbNr7XusfRXalHf8BvPLz+Nhyk9j4xB4Dt
pXyvp0E8N3/EOtoFnMXUhb6FS+XmV00jEwILP30ZJhV7+Gb2wv+GQktKkORV
zfdFHqWvuBNGzqjeAQSOIOBdk+ZxcqFXvDujBe5RvmoLrUifcOvIHpRrlLX9
FlpnpRRxE0XfSGC1xxwZwlZUc0dlzCdsK+U89s3hN++43LEQW7vjtWT7pDsn
S4U5Y4/wymGpoDqrZzsxNUXm8GZ3nRF4qZj/n+2VauMwnFaYdHygStPFyjVQ
DJdJMjAKfEXQtoB098mk5YzFhhSYL/TVxZuH+ciHTCiIavsJCaLgsrYfWsZn
dPNo+eWNaWNv2eOwel3XPwTBJn6SmfbwM+LK7qGSDJJMbfu2AUdaTG3uXZaz
8vbDtJZne+eiIGTo07p59wl+aLwjqCvK2XgYi9TNEEqA7AaDg7szad+CygP5
HBHBDHZKx0JvnrMTgasZyqMERIBJu8/MDHocRTMjAtvsPss+cGKADiigArWH
mG6FMGcIXha6NdmTjuEdPtcoid2jpirXdb3CWEfkl7dJ9vInJgjkQKSzW/wP
bM7ZqOJmDkiUGy99v9nXU+l4spJLHluQiDgctosTcs6QEzKb5Gix1rsd2lXb
tgwFoHo6MOKtKaF5kNq9ID0IMHsLkhf+MUlVQ6qjakZc1wXnLa0kLE5OGUid
HJRkhPxKvKQVvWazg94tmJGl/KWwUkmp/hDk/PwIEy81W3+4Q1mkK9QEU8ZE
xHFoJMaIkpFgGsUXnUyhTwFKdp1PuoapJmD/Bcf3FP0uLb1tJZgxqEkstIFJ
Ug6Mopgmy6uBoqjFhbUf9xr3+Hhxd1IQ33+4D75dDECFXyxvV3SU/WFOonPv
b9OWCgecSLtZL8PoSz0/Wfd8a8msbBez3eBZ4V5W76t0r6fGLz1GDJZAEs2w
wmyVO+VX7DmyLNOHcAkwKC9mSavCmiV4mYCvpeJInqt+i6pKtqG60yDASpO7
4yMeUQFF7xtXtMAFURMA1EoPh5qBZ5NIFw2uj1q06roHETCNgkOyhxriwsgJ
RCdvEJos6qsTAxXrrjhXKI/2XMlsf1Cj7rIB2kpTKDvB5cy0oXTgrJ83azzT
Usoyzv+iT+OepYsX0UqYSfbfCA5josM5laD/76o8BZiXYGcpm2zE3QQN+uwa
Z+UscHoml9DtSF+E94CxKFFaB6UA6tOAGqPbPNz6Nf6UzvhHr6J5gGKkTtKS
pUUnCbpeOUON71Hx2GKQTfBSi8G5ICsYxeyzZmo9LTSn5S0v3UVDQ1dcfFqB
LzzoYJeOMg0L9q0E0G+ZmoDOu/LYES3BtHaMFZ5AWk+vOxp3IDdSizMPnhIZ
VRnYOTl78N4JVPTQOiNKjQrLreIUf/KFmQvfOl+YOh6dIxSYmF+19O1/zaBZ
PWo3zXibBbHY2ZiOQi21apxYtDtUsXglTQ24XoMJmO7AUSd9m92tQzRDhlct
qUUDORTkandpzR09TO8A2IbvrWKJGXL1FqbYAu0XGa1S37lh9D7Je/5rLViv
aSzPT45PLyrsTEBdPH/OD5Vh6WI2Kln0tNOQvqWvyLm9Rsu0qPZoWNCRkEKJ
l8tw+57zYk5vEhdnrtsDaJ7QPXUCXWJrC4JdQ1R5XrPbEBxrX3JrnVSivQ4M
A+6BTXrBmQqOgRZdTfedt0OjrWf6h2AXPXPhdjf9GjdGsA5KZGxxaO6tC29w
f1rPjcqFC2d2rmmQXfd+7ebScXHxBOEPKwOIjC9afFq5fap459aVUPUtqoAM
XABT4Q5x8+WPkiqiVViKqv8B6NOE6u65IRHXVKrw7FQBr984X1y306TKNWDn
VJC9kGwcgU/Ti7doq9OQJdk5Z2l5KqG9UYs/ldMef40us2Zq8gEUC9kFoIWN
J7Z9VAbdx16qVw0ucovggwtOxxTBuBZ1Vi23/wvTYgYtcGyAg7HPcWooTTmB
RWra+SNp7mNV5AJ0Cpbj8g4o9jYHlFAImAn16qnRZF/Fb4bInVgAjVX4Hh7m
ajbpX8+ec1qQvFn4hkGm1s4+iogusizjS/CHluQWk4erZzEfbD0/4FgmZmkG
A28bJoBMBh8SpO/GLPmBIvSKk83SAn/Rd1fPHqEIqR65zB4FZNgvCASpMBgi
e51yWr0uDAT91ZLs0tDZGXvYDAdswel/Z46MHQvOfL1SpDJuEv141RAD+/go
1dSNuLvV4S5oG+4o7sOkcKu/1NrFIIcDj3fZBIKY53HYVK1xixG8fy/QTjOy
iGejULaLPF1Dr7yPlP5omLxYXqQ92PbSSmiuuQwEZ2+hSkPXzA9NRTyZGpbe
i/6CE4+Mn4wqBWbEE45u41novy0Pw5Wn5gW0XFaV3FXwvKve2QEWl4RtKz6K
FZkQXjYuG+KkOHMuZrRiTcBZoVb1KNl6k+AV4PcBQjdO2sJVnfTuYZbYWm2m
U9b+xAvYvlLnL+6UetYbznbcjVUfqyES351ATnHi3ZN/ZBSFWHBnQDYPyTER
fJz6aO0BSwVfnfR36QDCJx9oN9VFGufFpuig193evcxYF1fheTz4Z8E67VQ+
vGmWgg6A9q1xKjos4LwZrMEqVpP1u1ntgyxbXMXTv7rToGQbzcx4D0XklCQ6
+xSH42HTJd2zje46xGiWjzMXyeZqqJ9xPLF4sLe0I4B0U59/hsIo60qN237D
VNbsqiFOnw5EzzhICDHhvNcU7pa4r9/RbfrPrLKHq4SchPFfJ8h23JygwY4u
H0HDV43w8zf95GNxi6sEpXuQO40gKa3SOW8Nr3w3mgOuzsN0LVkeibohNTiA
I0LpUgg0S9F2sk/Ykj+WwnZQSq/V9RcAC+eVRy6IfICJsVUGo91zvNixC8Mb
XKoV8XRnvvZ418HAUXuS5ApP714+bDzVuQtil8Gnxp3mHresECQRamEHFB+N
YDJ1jqtuZTWTbEDO74gOgcSGNF7Uzk2QdmaqxsbtbnpdmUpIRHkYbJegX6DK
L7vuSAIl5qJ081vfmeHjNXD/TC4HX8Ii7tjuNoaFduY5y/lHBHOiYUJlGVFh
qljEx1eEBddamlTgnexkqpq+FwiM3w+6mO3zKNyXUId9HmuF5apMI4IHfPQq
WQ7MAU9KoSr2hEoN0ndnC8G55gD5b7ybGw2i9qDlKW74+utnkK6na9cpfVen
1W80WTT98CCwKJ8O2Q+RE6Ed8O+OhM4VKZEX36qiLSMzsiJP378+3vzLCO3H
p5G83qDQnq7IwvjSGfH9rcekqMVWtiZVuSnR6WnrCmSujmSNTxIBTY1NsK4G
Z0DGRdGxHf1Sithy/5nGQFxs12227WeHETonKEg1PhkeGhM4ruyMxxoNl4x3
OkDlvHzrvIBrxXD2QEZoFUbJKyi5ut5uEsUUbm5kGZ8y8zR4C+DEOFvW6aju
lras4chmyZ6MMU9ZSufkoShuDvfCSzgIeNSK0jXiBe/BN6CW2isbZhTkKvEL
hBMDphQ3KpEaFKUIzMJAMKNLRNow9u7NghDK9k3whoR4UYXdLAXgPNeQAwjN
XXC57sHx0x/CaNJFf0KcIX0izz3q9aDNxsXePOHMkNoEdWa4cIezXZuw/pJU
o0/qNELoQUursGyUvX1OvgKF+2xkqDEbpkKzGjT8gNBLuC/CvjNrop1Kwh/0
lnInCcqkJvF1pGT7m/eHLKNxofjmNjctzVem/2pqxADSqVBpT7u6/TUFsc9t
IorfSKx45QmREJAU+i6+9QWcv3wZAKc7+WHU9gFGveKfgU+BVOh6TTc2yEvq
Gx8ugfumri0NVEIAO1VAkJpJ2R3oulYQ2brHvfzfJW8zBtQ8CDs9/duWMjFA
PtAzQO+DjX8YDgzOwKTsdpkT4jeaomFg+JAJAHsJZxRM6UY3dKJputMixZki
PN+17R82QxKTUVWsZQHiMjqQikUzriGcmlr1L+DjjTFmm0AMlRpr4h6RhK0j
2Vn6C1Z99DbWDiw0hRgKw2aej98bEE6M4KY0vksaCAtcXLC7UIxnBiH5Fqjg
DUNpK8IDReRxiOq7Jkbh00QVNcOT7jJQsitO5YT1iobmzylKwVhwoPJUUyaS
Y2apPhinwi8ur2L4/bD8VTMiWUguznMfNqXMGLTWEU5RCW5MGRJOIOKFWzhK
Y3DYwz2dqoUdU1Axcf9cezOd57Q3a9ZUOnPP7v13nE5/pV1+ygkA1rak44NR
8x4xVHP+H4KCNZ4CC/OVfj/YkT9TFEVpC9I4mbul3lb2d71MMUnEiETN9IvU
vWN+hmm5tfTSVXV4YSLJcCVxUSGPgk8E0oXMMe1UZjje3MUwt6JhfCnrXSk7
RxG6/VNT55TWcBmg/zldCSEPdji+r3yiJYb0UQmijLS3hTUxV8DyQTXF3qET
N8WAasagcSyTs5pe8wH2RpnvqYEi5kJOGa5IluZohC8wqQLm+ZOiM4BXzj+P
9fX2DSyjvVhfcUgMfrr4xiKQdwrA+AS1+MMggiBg/4MK2o/KkLg1L76M20p5
MHmYoAyT4a2pRKIVzfaTb5QMdqGBjvA0jdl6g3kWbIZcwhtfiEMvvc6unkU3
BmDBZh4q1gFR/8Dqsp9UhLQoQIIeO6vEDKnyH9HH+vkzFWvGQYHN/4uejnJ4
gpPsCarCCTOM3KmF1yHs40XAg4JYviJnAnjIHgRCkEuyP9WPCJxpO/zSd/DJ
SJzp5EI21obzbnx8rQcCVea8ZvT7DtWiefxOThdi7z8x9BkZJgLQi2VhETcN
NMs0A/m+1CyR7xEOUoW/0gEeCXVp0H8JIqV3xSiCYG9wcmRCXydAkiq3w8if
lxs5WW0CvNvPbKV1yFV2rWljCgu0Mbv57j4tR51PhzEqJOB3NDagfpzLAaOz
vRPm3YK3UxrE76wQgeDTqcJ8dwE8xWsxHtC3bI9ZJV9PWM5PblWSL5lE1uQL
qqUsj62S3SPS0DEpqnjxW0xO0p+Ta/3Ork3qsVgRtmqHm30kIAzGYykpfaHe
0XyMs+ApQD3eUo/2EIjrrHUaOgr5Sv7WPbSZjLCpSyMnSUcZAyx3hT5D4Qdn
PGEu2LsPuTKqR5RITmJ5TvkWg2vxtmDAjgi4V7yFL+5FyxhAzS3al/Yemdc6
voUUG4e3zL3ZgjsBVVHxazOAHnJRFzn7URgEIyzprUlNGwvd12d5bcsnQDs9
ljwBQdwzqAawpMpDE8b1eFWVSb4IC7f/gLIme3EaiCxgT0e1mBYrYt0chETL
WO00Smv3BjoCPhxSqJmWGIHY9fWm6WE7dSINYKu4XUGJ70USqFozgrRhYh+H
5PzwCvV6+DpwCtAHb+3B5GA4el4+6XFMcMbB1m7SJ/z7uJdDRqQWnxZTMG9k
Z4HQCZTjJbe+mmmO41o7kbC421Sju90/UyOIVCbOxOM6mcTWxS7ulmXDY4RH
nmf1XTGC7ePNQ8QJWJmC+OfG2hjYp+ysbLFAN0uD7Jtx74Ou2TXzm00kGLBn
uCaf7lnnczNXR+2Tw2ejdQ+gm/mES4GfzzNb5nPKEVjt/6AXx8DNAl7DFavf
dtwNXdXOcsIcpl3DIzRvZW9OltPUaJPOBlW7S06Cb4lmzKfG6ndSMs2kzJsW
Sb0T6FLo4EqIGNkV0ql8jxhC4aNhtIKOV2wcvFMkFGsrKYvyBV7piSYCgKMZ
bo1jL1pmSMy+SBkWdxBfleJ1aAXSo2ESDrsi6OU6k5p8MgHkMFWRk6gFapot
IpayEM/vO5jcd9KFdJScBf4Mi0weqjGfG4egDSfg59ICtUaBc8zxLwa6a9Wb
lOwqQ/LhQ5lSkw7njCj9ushzTOMJRo8n94uP30FUE6SPjBSs/Xa4ju1zkI0K
gzTOc0Ot2rhCj12c30zHXKXoxy9lTh6umwZ81pzdUdypWiKV0siA+uDUR0WC
ks4lif0WNK1H5sFkCbk+EqcQ6gEJ8OuaCFhcJeB+jdalTxRln67/wMC9JU5c
DldrDjzbDIKFqv83dErSi85xCNo1lVkIZgC4iQ9ZXOyXcpa7NKkH/cH37Dej
nQ9F9ZBXPQOKSYzemO2JmUJMuZCK5+6AkiczZSB9OIYq9WHjfcSNbTY4VqKz
pLLgeluphwdbYMA/lzQz/HSEP27+oaR24GeuGb9g3FKmRCCFHJygHsnnLW7f
vgARkFrRplPFyP+IGnYw3an2f/96zfg9KMyfEQ/qJtWpIY+G7urhNoudusZ+
SCOPYJ5XaO6z9yFA5wNlphSpyxFsY7Tkg4TdFaT+kQXXErSC1wMYX0UxA+ql
WOlvY2iSFYYpCKelbK2hK75tTg9To7Tuic7Nl6Cxwmm3BDL58zvZmMIVEPD6
oJ1/2Ik1Pe1TRyJtfHpOPlPHbrsDLqxYFysMTQnILo7GJooqt5Hu00HFKiN6
wgAN7tnGo6eKtm+5W6ruQn1V+1oqakugGqwXscLgB6rW1D646ach2ibMhBqn
ZXgcRjPKCEtcbPLz64Jzn2cwNlcv1JfyFWFS18SQKiWMJBE854AOvLbS3a8d
8zhbt5gWD6KbLBi86/AQLC3tu6iEJXb1enTJA9Y8fI/z5qtLdg/1QT1DL5q1
D/HB8mSQwyNm0pwXcYPCLhCuVXvqMdB7x2aQE0mLURDWjG6pg6STfk4gR1k/
8cCC2DQGzqqUPQ973ADlXFz3wp7eP624jo30CjD4RVc8IyzPFxAbsOuetYZX
TIcorEm1w5YNkfNf7J6qeFMiGDF6ko10C/Uz0FIM8kI4d9lE1/6qeQzrX0qd
hKPs1PCKqkJrjDBkCgPKO2vzTApHt/rspspirZkopyKwb3mgVeSkpNBOBDRP
5mCXB5I2sRMbnfLBMN290lr/+9ujaTMU6R5lRLdoGh+TYJEROiEwfbeKbigd
/IpLH2JCvuLPQIILUzsloT9SxM6UneagCrbl78t8t2wCFSv7FST2AfIDd+f6
7QUdqfH9QzZvX8xZT9RX5Qf7NJwIlGOWleJSlJTnzUGwQg8kLyYsE0gAytKH
UMvz9lzgkkLBoNV4tAiQcGT8GmtgQNN1Vhc4S72OYXqA6TF/Mrn6oBCcL9ik
McLlLCvrwC+6xneODH+P4+iRz6uCfuvKe7l49gIr9UVVdnrKmhgzrtOyhppc
af8M6LjxfetyZa8/qfYq5OZ9fGakSv4BDlBkuT90k+I5+TQIPTfbP2gs3umO
Jhq2OfgsFRWRpXfmVYWieDgstVXq8GDURNEjjzC5t6VYEruHVoG0txIU2Ohf
1w7fhInd2k40hebVyEQ10QdF2LzDHxzYmlzeF603GHD5FPtwhZJP107eaePK
wKXIKpUoOJXv9EVvly+rvIrQ625/upzYr/T4NVZ/AVG3nep1ieYDPBWkSAH4
ee8YMY4YdMeb5A1l7VueMNVJiwxogttvPfBOz5Mg/Yq90YL+BRTs/iaGnAEl
TXpO2Kn+flo/TZpXBhhTaPEsOMZLSuGUSk1r4MtaZmUF8sXFNP6SFKqy5JK0
P2A31pvr7gZqt+iaqaxTMI+t9LP7x6okCywwCC8/NN3k5DD+I8E8J8av306f
Y2M2RIIuv4G1YkoARfQi8RO7hEk0NYaSNkrh0/4yqQ2twOe5R0RcCOwAIds0
SQ2tXOYu4mSOIxrUjSOyBSlu8/CWGDr9zPQXRJqGlN/kwlRp3qLPKi/Gsu7S
C0ynkem3Glm36BGKGPPV2az9ANrFB+KJU29VxxFoUbQNUnSCPXU+FBtrjvBx
3+V1bIGNQ8hn6PsWYWzLkYsjZTbPYVd8Q1B++7NhaSQMOuFP1nyRDFpkRalz
2/GsUwYjYHzvpZps96jjjxiSkeyhZxOuG+gYWKczsJzsX84J/6qF9/Rfmy2D
/yqbrIii7/Hn8Re1x255EqAA325EJXwL8asx7+dB1s1IUCDg7/g7FCD4tJtM
vCrpvlItvDTd5RJwJRIjl/jO3N1g4MgTXYE63NUdD1H3+Dy2Xwb6/b+JJI3/
xiAQ65NJmohLDz67ec0bF6CH7afNzjK6POcPBi62gvd9fmrCst5828fxiH7M
CuP2KkeEgHPt74x67Rv9RQU+C51EUOgi79yPUOVIEvj2NTErBsvmJdbsEZwA
pJk7gBr5TyXTjQ0zMMYXfZOk0h53QXBq/L0GV3FWFfvCOR3a0ICeQbmbaVLl
25lyTVYE0N442EZhaLhzbuseUzD7LwRs6aHD4g2sQwVw/dMw7VIYMbvud/x9
npk34N81eSy6NSEm/PcvBJC0/afEDQaFHki+xaFTRgY0VDu4w7Z6KDS74gNl
5e2lkb42+GG72gY1Af823tfkXLoQkTz/xTVFi221xQx/+jFLxRZt58qFFVVn
pKr1wkqe23rcebAxHHH3JImckL2dsYJzy3teY/cz8qbPSmw822bEro8k6QZ4
iDepgiEzRNVf6bjZl5Wlq9HrIL6cNkEXd2XTbCT0qoV6g4Ltu0YysUKt44IP
ap9TyUFwL3qIlM3sNWcLRU/cQLOZpt+iyFa6KpIXg8HUYV00f3/7tVnqWL58
nXRudLOr8iyqQsRB5DGlZbIKCZFPTHYt1dUZuMHTtWc1J7c3DZoVkheZpYQb
f3Fc4Fh2tGrMAdTx3BCZJAxuaAu5f2vLjrNOkxiXh32r6NyuKgAP1PWITaWw
YgiLnmQHVF94ukdKhq9nkgpMnIPL04ESjZ73BLxFfvObW+9cWEJxfm2PzWso
F2XieoCVWt1/5fFK6c/8urhg4+ZHNbtrWNCt/XV9LORTCSuffWkjW5sf4Duj
Ik4Kc95Z6NoyxVmdAeId39FLv/d3w4al1QaP0D7djQ9xNDI/B4xcxtXYlNtb
VZDG+mepbrzdlE1JmNS7Uaz78DwebYbaFW98/lj5TGJ1HwpIo5WEsEJzCXjo
ZBpnY2WszhFI1zw1yOtnBFqWus9ecuq0WT/i2VAy32InGvA2hRx030ebBufZ
DU8Gi8+EA4Dxw/ovy7BYSVxtaXTgTmT6w61U99sdGewW1BRNWhlbf07QCPkw
xtJaE70KTqL/ZkMUi5hqojpCP7z1ncIQQlEcNVJkjTUHpsuf30RPfSz0C4Dc
agjj7kGYcxcEqb1I26z3aglKvFST15I0N9FypgyMpBFt6BCKmk1Xra2H4rcY
qqCAYm6wycUHQEZEklmzcX3FRkrRMDQF6QrhhpKsjG8nmNW55N8Svv8L1V+J
Von6EhH88sPqDzBDX5iiSCQUBTL3KnkUYRWjGVvOFSIMpJfwf6X34r0gYQro
rguB3KbdiZeE8PSX1/LelKL29O2HIpu6ekJ/HMyxpy56RgFOkdWi4m4PE4of
XRpK1eSHCcCsDKeUKutDtijTsY5Tuk0LtTOwIsug98U94rCO/GX1eWkTlcG7
4AEmoXAOfk6QPnRBKNCecrDh3Hskq2B1P+SMCxtYuULQpyreRGNoNNskfe83
4FDBk/u//XmxPdXAln20hiEgvGTM9LToen70ihulJil8smy+lJAiMcdn915Y
V6Ry7maqBUizCQiokxu94BS9FABINXMXB/E1RT8Onzg/Vs9tCZ6tjpu7CUuW
dLk5RRPfwqG+ILZB4EPaKcySlbNXw7M8ullwWnFjdel51LTJGYhZnxRwnPRd
3DstNkOPx1+eHaITLZ+3RpKVbIWcL2XbNiAw9uSbpwcF1EF6NF7JbC2AquOg
NCjV9+7f0ec8sFuvOVXWjzd9ArDKzZCPQj7USj9EfBe1ER/ruXtArbusGjQe
XR9u/9x4hKIIzdLm7HPpN6dohXENJIDyBN17aXD3yyaJo2GIiLD0YoSmvRlJ
HqfA8G5zvI6U+ER5q9SaU44rbmv7Ld/VeGJT0RiXiX1SORDrwpNYVzESj2J/
j+e9vyCgFs/x73Rn66rVEsVtdLJA+nnUF74amBcQvuDvgwg4FCnGTmd6oAiH
HrKRwx0kk/+2Fobm0ScfvLDCOpAY3B2gtn8XMZeTeAz4VPw9FfTuvmVk2n93
SoRPaPCR7WXjOG09L6Kr6cAVfMNvzUjs3PsVRVJTeqVt/IqljJwpnMbPa1+0
FQgspYwBG8yY//oo/5cPsRzxMGUFXHolDCRp+6NkKacgqdR58lLYH89pH0RD
JnLVqTVFpAfVanu7Q5Gn7qxKM9hoW+/EXzZLI5DHZ9F9FhmUG0+NTjreNHFb
zyILFIoaj43XLxxJZMrKKusf/IMADuDHOFWzctQOSUgUboNiKdJt/UaY4ZXX
yfP21+2/pl2nM8DWbQovqNjQy8+BlaMjQbv/BzISxkqiy9j+QPdz4AUn5Jz1
CJ1C9CL45MKXLdRxER3fgAweHeF8yeH/HNnXMX+Ro+Y+tDFOheKJt15v2Tii
f+X8z2VntFidupHa/EaKL7QIDw+CfiqSN6WNwNBw4GFLMfcNpJkakyevNeda
2IoSt1YIhO1wht6sZxa6tFbzlku7VTlqXThYLuayfTaKvqFj1UuJJPOVXKzc
RJxzJW+QjVcNV8OnBHPsURxbztiTs3tcAwJh3TD/Px1w9MACNukdD4O9Jfo2
bZ4DuLSL0C7cg2s2Zgo12HyCk+k4aANTdACiS28D4aDBePpFaTdAGuOWyizd
uceFD0iRRAwTYr/W8b/7B3/ozHBEILuijR4OCaqbcF+8nNhABVSMVnF7eL9N
6gAx3uzzGhdBHTYWY8DfqCAHb7CmI0pC/0JjDvtl8xLU6DgADEvsCIRe9roO
hZbIWoDaGDHYF0mLdRIW8PmM5MY2J4S6PZERqu4Xe+kLvExSon6JF7gTzwJv
U6HfbjoHSIwW37hvnI0r76p1+zmIUtkrhqMR6WQAxsAkp1HwCeYjwh7fIU4Y
1EGtOfg+l1DvRRJ+XLg8b5gLp1htP6iNkHsNdRT93yhI9zzOsN9Inr6zZ6/Z
48MOtI8X5rAulYPZEWPNOURbr2yVM3pnGy+3mII4TZ8zco2IEDmMH+3jEUNx
OEfQyXF1QyPNLVZ8EmxXeKgQJFFgo8AvwmKWrg8yONpnCQrNl2crZXdG/1J4
oqf76LD4iVQMvpnDUjAQjMIPK2+yBwf8CFhCeqSidLNsbX+BxG1Si92IpTZZ
D+y8TEbTpQYI9XMd7h9Rhs2BGrSollstAIyaOhT+v+gZPJWmEqKQvXHjqaEU
Dh3Ex34AxIcp1N3QGUg+3Wc1sTqihp7/qj168rQvVExeJeLS/fndFHQj9CE5
M07OvZJF2ccKznthXGT9agDxDwVEz9h5XnQiL5bNXEfJUVZSlrAbig/n8yNS
okZoTOCTLNMTfS7CVVTxYkqb3WS8TrQ+klp1FAtVDZ5hgeLjia0R1gmXeR0j
Ka39rmz+PpVibb8lTPh4co/sv0zrLo/PnkrurTpxN+/izPgI9ExDjlyq7UeJ
3PWm6gz6PIZgwGkBaQXqLrYehZYGObUBIhmNnU3VCD6iBkqjrq3ku8Vop5p6
8ojEWOMbks6QF6hsuBCsmGLkjL3ZLV8eoirOecTEeSg2rR3tcEtul8sZXajv
lVwSaGFJ1E5w3MFuDNe2GKUwD+cWYiciPwq1sF5uow55isg9oJYpsdk+EcgM
V/JIrrcYuYgAcwvua5mmsVSuohLSSSwOPJaYmKUwv4fYqQmLu027D0AR8qrR
Ox8lSROTbRwWB/5EYm+eN34kAJd0pp08G8RGWh3rZyLA9DQ1iIE3xuOgfOHU
ItjOUH5DZzZ5LjBWzIABpiI50f3I67lranVj2P0pfuzkn1qKDzvhu3OxXUdy
dhB6deW+hTdBEgf1JOSywISF6yy0XA9gZOvTfONirM1qgVS+M/qYqBls0qGv
AQ4wN0pT4K6rQ2cKqo5nmvY4JyMGdm6FYpW74Ie5APXKKtpY4nboblbzvqEn
v1713r2gG94zRwdytczVjaxzBfurcjmap815k/l/86xnffkNsV6VuWTL6YVT
WcKxdjOkbvy3q4YtLK4igbJ0MpuVms+jU1K1zDY9HN6eDEcM4jZxtILxc1Ml
2SrlX+8+SiGH2OySwT27aXtCsWuGry3nAnXWVEkVTXXZPXCbLlMXkJNAPS92
Q7nh6fsB1zBaMBZcDBKIe27y3mNpmuwIA1rg5W0UHlqhT8moRoC0o4tHX6hS
/j1TuShQvjznBFkYkwPN/uVR9UQen9nDJkoNI1rYrXEnWSmpNfwPNUW70v+4
1k2DitKYt86XK2lv/KQKH9JXe/bxsrBi6vHcyLvQ4tsJFpYLTXeu1ZWR5jdn
0TivUTY/xWT1FrF+OLT38iEGH3RbRrkaArqgAAVOdKSXM9/4MkyuqNcSL5BL
zXFPTz0HdI4wYHLKIdxhvcBm2Ivpsz3rD78f1apkNzgf+KvQYnBfOlo41ZQq
u9OehH9uIQxJ17L/GgxYDVxVfGo2O+Pk5qadCo6i0YgNp2gPD8HrLv7Y97tV
e8dNsrhc2Wim9NV7fKsu9pUkLB4cND/mJA+pcFJszmQL9oRbzFQ8l+AhRVgH
3YD1OsK98naWTCEIwWHlWarhiM0+n2qXTfzzbfqtLlk0mX4sV9VAV/Azdg91
0WRakmnH6k6HkzE7KJ3/nTVAM+mwbvX9ZCPE/93qCGaPL5U2FNCQkwl5fsVI
WKEqJOjFk4GJX1SnaRbTKRd9ifnhqZSz+DJA3dGDkyrEZrJAVoZasmxs4vIA
0ouO4DyocKMRzzOu7hH6iLHzLNiMMy2Ih6ac69Z5ObqE4I199/9SF2rUCv9s
cFIaNjb+6bFM8d2OfATzysqzxhpVPxr5JFBPc8SJL3CCOBfyWADsFtpwEDBf
sFt4kwkz/pu71tYu/fTZw4A/toPigG+ef6GI2NpxL/n/+T8n70DRniHWu9DK
WdcAqWcqefzzOiS8JM6BQMc1d6lei2Oaig/+wlpd2Qxo730EUx2FIIVpW+py
fVsRk30+DKiaeFjO2YXBpfO+ouczbVA9tUcQahFZpmqbWQwLJgt27QGb0352
Uog4Dr1PsjiDiDdGWNApKDUd2TuH2y0M7+vtUPU0FbfOzprNZGSyE+Ei/xbn
ffvBaa4IOWhvcjsPEKtRkERVUqXpSeEAeQCMlN0ONhH9Xp2vnA5F2LiMH/xI
Tq3lqNRbB3CRuF2nXpGBoFO4LEazWYgJ0XGptomPZqXbT39fEtpbYjGIP1Sw
3o84fgen3kIXkWAFyHhzgu39owFVKGPRWaXK53zYcj449plyHUfR8w6qgd0B
r2NkEb+sDeVBXfmuDJ9ce1CbnULUGuKvrQENf0ft7tJUizXk41CxCyydIjdj
/H7vFS1S4qWTcc04z9TMxgXzmDXauq7oCRB4YxcIpCw+hnvwVq5oyX7oN/i3
37zWPVNGXiC6FpB60wgHsm1hYip4GNPujzdik3ny0DVLFxEyz0uDxmWTy3pW
zm+8cvPR16jSGwDdyTWaWwbURzXFmFeus4cAwcxIeDb0/a7pQpLx7zgeWFFe
4Qdmlxa3bvQ9dO7TdsLoCGJGTmqA0mFhRIPFHyRKmJ/dFpmT39aVxaGml+ie
3PQJfGjMzJGykTMcSkQsUXoAiOtICxgxUqoWB6nys0m076zLxrgObHd0hbH4
GSmTLZr11lPL1pYAbOwerefz8JIxqwdVbaGV9rUUUXJ/CjerXb8/yNF4otFa
U9A4w0GtLT8GDe7/m7qcC+KyIW+6/FfLHEYTAjGvVgb2wkZFRKeO5wKMoP2R
GWayDNdlzvWHGDLTnoD80RnFCRU8Qyb0B41J/tLciIuz0xyIHR/c/ZnjM1re
6PM8vdSzmzuSPueVxnIia8Gp30xsMHXxqUFGum3Ln8Uzjn6Ch0BpWManJ+Ag
jOXe1ukai3IUG/Zi7QXx2LHUCwV6sQAFelH7dkahqfpltFRhEeDjJqQEChbb
VPV51xiWNOqpYMyuhJAGatxUx/J2YolDBwCLsaPlU25HYkMgyLFTJPLvbZPk
s8KgVQqW+GKMlIgtJfqwHLQnfcqvYAox3ixxpQ0mvPWBaY9Yjxl5SFx9UEA2
+xg3szo7Ti0JGrTNoiAgZ5ncRHmPBqo7J2yxP0mIn8fRYJcgcVfngJvOLFOM
tWpWuse0s4FLT2gi/JUgL3kdfvDW9WvO3/ZFAYN/Px9kbK+uqjU4cFGZmUxc
AAkHdlxh4hfKYv3Y/cDs6bHnF6BRjN6AFwGOEK5d+/VAAO12vhwzd3OsZ3yu
cPCTCC1rb0sVE0X7Ff6VFyvXfIN7IlenfcgA/QleAk63lvW/e9yHUy0qeDJO
kBy8hkN9BdkkLx66e7vqaAQf4nFjclopYtFjGlO824sVNMetb/Zpx4xUzqfc
9gaM8DPggUVbZ6zLMZTsTnQ4EBmRjDXLEETLPiczzg6Uhf9jJaFZSvnPIHn6
cfqZJOcJkacxX95tYpZHWI1ixwQ2Wu6wEKFktaVILl+cCVJ8WuK9Ibn1OOA+
oIDCJ+E46bDj7fKuL/pZVnAoxsjiUoyES7HPaKsvivFBaC+QlWq41qeu36sN
CNo2WBLCszaeIf0PxurV8vRlqrq1ls/lddD7XvXEUlQG5wgk3QuPqmLLTCyb
PVZJaUWbS6f7PdA+wP2/l9Sa3kWkkNmxpv0dP4ko5Blte+ETie1icIEQ5oTp
wFcOU/U9iPrhuO2KrNprWkhBq/V8fpj3S4qdn5gfVD8kNNx9tx7rGeghnKPb
WUh5zcvqlSCP8WHC1DxYMhTictgc73Th9214F1RE9vJX6L+ViMH7JGOISSkW
mcGp6ekwH9+wKM+sx8nLHYp6MdS9TDqkAxdR1wI3T8z5aRP+2R4xzfhvwFWQ
xmkMrHaGQTuKjKTHaR0KOV6ygWWhuD2WLwB/hjnys9iKrHm7++ANSROzQGoS
0+6YASR1EYuBiKBw+AkoX+WdoICr6S7fIj0QY140sy2yvESOiWU0ClUENrgt
dLE0fMbZm/QhL+4OyR4mUVAnRNQWWLHO9pvyfVewL2WB8/egVynkT+6VfdjU
OpzFxD9Uz1zf3Nl7ljuDORKaueAvz8R4r8Js7KURCVzSZU2E+TUELKXAe21T
1HaQ0rjA/JE2mFj9mUjTCaSAinNFnU70fH6hEwyT/axGF846G5JpoGP6OWNO
0b3cqFKcNrp6zy9feNqiGYlENSYFWXRmqXywTBWqekj8GqvhyFnkY+FZVQEz
QvNAbK49jFp+ZHR+dQR+TT60c4FXBs58SfxtrYh05Rd9IJX+y4F/bRYBKi9d
sxuC6uKGO9AMFhzvmNnh+MIQ7pwA62cc+J3lGgFJKMHIqJcddDxXYDZ2Z4Bu
w1WB5OpU/IJmdiEm9z9uO3Yn5svajWeISpsOTKMxSEBKNveS0MvapMh6Nqoi
82pWZXeA0jP6DXWDx0AKztVmW8IwqNjK/XC3wvGKNlbhRH3tteEf7VCYJOw4
adOAbp2Y0vkguOW4jFMHsrrly+bqH8DJPpKcHqdimK9YKGhNNPvDc4m4qmko
8pSs7alojKGUpn1+7LHVRR0YVMpq/IY48Gt9FUqZNwvz3q6rnvSlOzP6Y5aX
NF9zdHPtaabBGfK6aO9OP5c+4PAZVBXATuurU3NWah+Rn4hJ4q4niUweLtR1
Ag5NaHuYkWwNTsOac2opG+zKwfTPqEdwJ9tO0YU1lqumRnz/6S/qaPBgFXRn
xc6SD6bOqwUXqADwFVbeT4YpiAOu6QHh6VqNd6h0OxZfxmsFFhQvKaubLY1m
n+C0VPDGgGaR6vMZuR7bH8nC+IZ/NZRJ8Xuf97bNqtzfwE+JP0iVulAMqiJh
MrjXfGjdjCtudAVYVKG5n0D6h+2kQO/Jj8YMiXTwu6c8W1paHGh9H7uR9DAB
ESncW9cEuDaUvbG/Z7St8P2n+XhrzXSgji0iR2WgXbvxfe7Oc3CnQU9vx6Q0
VO82yGGiZG70XN+LHUpS/3o28xbaOok26Un945aCIHTxWKkq1vtn5UY7nxIq
aDpP8xvEUNtDst4b2OtCWXkoeULQpb361cGjNG7eETDJMH5mHhiW1TfBspsj
JsEPX6XmU7E+5Q5zrrYLQ7/rOVDYek3wn385PVufaEoPMBxbd07ENdq/OXpf
3Wr5XFQflzJzFhaUKp/1IWL3eFDJKGoqgi7tb01JEo/Uzn681OSJ+IZ0ghlt
9TDVMa0eQr+86AFaCxigcIVZeBtIccLORe3BcRKrgydpSnWuybSgY7FoAhfm
mUFBzoLVohgxk327errbjjgwMP+xVlR3Fy1hOApF/GfnwAoo2ED90E+7fVVC
a2N9vzeGWwGI3vWRVieGICrnNxbjyyQynsphntG0f5A23TfuDwvef6Phbo9P
Bzdj+k4SYdyBsxldrE+MusziMf77cXNNW/rKdtqshiilLyMSHjLeHf/1aITt
5r/Iu0p/kKqttSHtpEd12yhB074c3hOUbKlrLfc/agz32C2Po7hG3vbSFYuW
AH5nFFLgocgONF28Sj2mLBSu1bY/2fx54HBlcdme611MgQQgSpUwhBTkbztv
sHkI2TvRNkUJ3r4vv9EKsYoB7E0MpteoMK2rz9Nt+CphCC6WUt+DDel//3wn
S/FPVm3GuoMtpkTh+Ro/YTrhhWqa4y2NcN9qr6zi/RFBEHBq+ixJgcu/2xzu
IXteKWr9YCjBCgRtAm4qGCajQr9NH7oZfl9KwVZgg+DrDTj03P0CCpGe4+om
vdhh0Ta9yrGPti5turLMd/4P8SbAEMD+JSZ3amwSsSfPkY6uvsaqQAJn2o0D
PnxViw2OUhph6r5NibPwoKLmyjxzSMZYddnRvGRh6rJdrIbaiP+/CGJLP8Qa
FR8Agh6TQQ3APfS15keZoLhtYx7pr1ZOMuvolx2Wc+gGfP8hEBiFgvaMTSsW
Q07/JtDsHrwMJ6OcTxnfdh7Xd9Q2EYuCO15dbqdabT4mmnf6Ty2NTwrAM+5v
IEFWI8noyMSPVh85lB9Q4z3GnksRngZXSaZL84Kx9nByfhi0bX4ZDYV42D4k
wl1eyQ2Fa+ai2ABRugfUNXuD2I1amdxhJdr58CWn2R2x+jXwOdvmeU2+3pIi
wq1O+22Z+4+vBopz5RSPIroanpETjXz+D8u7UNYNpxzyW8zeznq9n4SSa6FK
T9bpU80P/3lo3lzrlFm/uMv83W40J+lqIJUsX3MQbdqc/LRBmYf25D6v0bfi
ki3wdKe8ak9jaNJGRiYMJvsxUwkl3wtSp1JQ2bqApncDCtVXBjrHSqcm+9E5
RsFvrxiYD9G9S3O7KaHPhmzK+FYRXbUh5KNzDllbxCcxhgyr0LplkZLbOlEw
G/P+a68LqftbLjQ9q9Lzevc6uCTff/mTSIcFZo0KcjI+J/bZtE8qxubrRrb+
JtnW53atyS1DaNXzvODgbYNdMLmE5xNEZeYfCE3vuuyT0Iv4zr6q7zsHbp8S
dRALmJcDTKLQqPH0Iw/oo+lXiBnfj/cwqh0XKMXgMf0t2S2yGsZBfaU210lq
mFLtdJ6rW9UyQ3fKwzSfr1+Iwy4ZXBs2urT4qu8CCK2kqWz7YM5ScnK+WfVH
O914RyEr+p8iX44GkKUMfeDPzunwncxqJUN8rYsckUh/Vp6V/XO3BO7C3s6O
t1NryvTkVdhdH+3ziVmv6PcaSjeVqlKv8BpA9kYkwjvfF4gtFwVShtH5nnzF
kIrfbif2vthO1hJc21OihjaOOf01W5w20ZoVmKQcfvORtIOKL/MmvvYbtKC5
MUpvDfymtNonQTgECv4lWlxcxOzHqZQButBzebv67lb4xEv7ojARASgsurUS
XIpEHo1CZ7gFvru5jl8W7DneYBRyQN1iAYHGk0DCwwqVh5xAm4r0cbsKjo67
7IiwkVBBLQyu0O7IWfcuqAzq1ag09OnJHZUjyukVb+/Ao9QC7khGSVlUqMMx
cXgkFMrmWhYiCDUO8VS4JQCNZNHlFVLT1fSUoBZWFqzwzILnSYauZN2i5MGw
BW52FyIZJubp7Kyf/ZMrhyqpH71JVYNQ6wQdCW2xSrXxkzsyfjzUrsd8c34t
ibbshrpSwFZUJmJbvpxmYYk23mDqWjXnVaTbpxzNB/OpBCojcfLtXNBEmmcX
LN9j0FWorM1lhrfNR9yMIe1EFnUUlrYbVm8NSJz7RasHDr8EE/g0iZ3/i1KU
bw0sEa4DQ0eSa4iwZv8UadSNPiOZOGdOLTgS06NrSVPpPo7lR/nCxpx86iOk
Pp3h1AHRd5sCRu03de/W0D/7Pg/okJiqkj5McgIv4QotsijeeYYX6tNdHc8c
wXXrbJG8dvKOSExQugv5yJaLRWbG9k33ka7fOdUJbWX3JIrbCmvUol0K4tsG
MVIIK4S6Ik8Rb0vYu7Ym+kxmmWpXRmQDK2ZSB5SM6aDR1bLVI35xwO6Cvcye
MiyAGyP3ee5UeX4lMnA1GIzh7Kp+RUVoJWnyc6+T9YJaCM4Uvr0Jmb7wTtPo
VVFxjgDs03bJpSKshJjFMo85xKPYIF/CRwsXtMrMA3UaRomNbLVZjKMwtemF
tFkCInuz6VNGs4dJP3bvJAk+DXiy2HS61mST1kHa8OQTE0L8xqlGi/XlIWsI
+Gxd5osImDpEXOP34v7DMaLU58QS7y0f49VhU7Nsal1vVxTKn85kOOpY7h0j
H1H3k91PmWrXzNU+LSkXnq0LaBv1gV6Gaj42illVVvSdbkOmwRYrWsV5TCTv
nQtBgYFZJq5fzorXCXWBguGyvz2hAnUucg+N6ruE8URrm8Mf2yCFCsRcbyc5
u5Zp4bt2xhDOvytsFIlKzLoqMBVc7SStPNpDzs4ht1NzDLFghQBb8TBFeDyV
j2TJHtg3Uwjg/AoPNaIFw5uhLYNDLmvKKZ3bkEF1MLKxR64QSL+IlAFp9kFX
S4ymOOSZxWl4y411/rd3LXNZwX0ENDZtwKd4fhn0KRy3qh12J1sPhW8+jG2i
hMZxx+I7l9Yp7HHsSdyFXcxO9ilJtgnK0k1HWoTfmpCjP9VbuL0Ns2BumGR1
rxjeJaDjWUI+fuGeNfAnY00WRdZTA5UZ7MWg/z8ymMM/JK2F05+UlVk5Oz7E
pw5DogDIWoQhDQs4aVAKKWfcrkEVY0+opC7Ke2ljtSou7kp5qutFYzUzpp8K
0wFn3+QojOac4XgWkMe9OgYbqjs64ihaKNYFYMR8ORPdzY7J/RLNEB0Tp9Dq
QKEHFhBvDbC7lglMI0gbkus/1xe+LC2Az+qxPwpHWZ/ugQLQtCcSNoW0d4AK
SpcSJI22npcxJwZ9Mb5q2oHa2BPPb0RJZWGhEFpcm9urvGtmmrnLjtddVUDb
KWKR7zbiLsnbqywlVTpuggVmcepBcb2rHd/T16WZ6k1Li5lg3zjS3g5EV+WU
pn4xw4RfiBUBXKw65kap+9sWP74caUqLk7gvlZ1DT/2wT0K/8hr/leoRsVCO
BbB2Ax1lF82fzHx69ZvbDZkLio+FlHI32/MkHnYSaaOmMZDifCjzC0Off+k9
R5NEv6YgOVl2Bj1n/WiDauLEpg96sfFvFlDSoFU6YI7Sa8h1P5FJdDfkMmEB
2bFblMtaeADKl9T9mD8a69xk6V2j3QqfTKqKtRCwDOLNSK8zwIX7MWIQiGMs
p3boPKWDbBA6jn+Sejt3NzPxibmaBusFi4AVGTuHQ6n670Su+bhza6LrSJoM
eR0Seir5Lee9sWLQRUexXaVQx/klpqEBmXRGqS6wre98rMPqxXwFsx8hbFZj
Zwt2iySaGgwy0PfzL+OkE67NWJJKz0nUSH2kY/BzX4tPpAkiQXa2QpI3wMBj
PD2agKBiwpsU15xmzu8gxYF74JYxiacb3e8WaCV/u98NfJ90q2bppoz7anLU
EZlFbGKLqRjOQaWm1Vzx04lOIWA34lMYNZPpoKSlSytWfwhXyGQnJ2LQFGoP
T4sM9tyhNpauld1h9tsU6wjUvbm00fb6koDnp0to2+y3tLTER0U1Nhqp9qVB
BGZya2yACV0gG5p/zsZ1HNVUscZ9wtkJAZPUBve5uwYyiuIw08GFMX6TJRQL
oCVupPqZCO82fcL21Xz3OqVWPhkXdSRXa/V/vJdy4CX3gzrGChFB7/fNeTF6
Z+OMzSlBXj2SwUSLL+nRY/Fa7gIJ+abmaW9LGuFYm8yJ0nF5nZW8HRIbgXCE
spzncX2el4jSrjQ/r234ChdkKz3RNA2hqOwOMaKH5RpLsxvwc2Rp6/Es4O/3
bLL7Y1jiFgO9nWT/vCU8uSZIfAAOPOZX59WVdyLrUX/Gnr1J+otoITiFISGV
xNNdXDiGx+nkayfKyEQg/ghFlOorGd79JduMw74DvS4bOLVqROZjlTKAzG5X
ANDq7FQOkM7hSnqPxZFhxq1LBYDOEqOQjguJcsJ0a9TlXhrI9u/znTa4K+5u
df9CbCj5P6H6NexJ9HVrRfGrAEq8nRpih/f8Ry6Pt9walnARwjXkrQP/HIVE
WBngRWAdtqQRgZzYNsaPjDMviZasC5nxqC71zScBCsouVjWMHgsFvCqFy2dW
g8jxT1//eN9VGb3xISytnQqLSp/i95bgybFPZ7wj6VsmciehVLxEHJrYw3Uc
aHQdhnOIV7d2jOe2UpjvSpa8xkOJf+smW4ISqGQqGT8CJJU7DJdr86LElgJh
dtuYbX40B1sdDt0I2b+RrQe02mwof92HB84tNcdCqbA93pLwCEKxxT1LGRBT
T5XbFjaPrr5P/VbPTK4eDXBc+p1TTdBbEQMcvJVJ1/kbtacGcdBKBjcQWD7y
jsBoeTozNJ5ULl7aiVhA0EcTOXGx+v9Wb6GEqmMeGMHHWmCR/pbiZ9Mpfw2C
DpRtpQuiNpYgJXH2Aj1mIjsKUxNcpQckjcq3Ump8CoEYdY88ORp3N2amrd9X
RlG3vdGwUrrk091erJ842HLb5kQ2VrV0MSh5efWiYOGYeJuKvGSeg+4QtS66
IGqUk5I2kitPvWMI2PKNqDED84X4r6CRGDdR/m13vAh87U1QKkTrXU/393QS
JG2bTpX+Hm45FUzZPpcbK7XtLfdeh/4TbksOZ3pVMa2OdK9iJuSLq9/67yZ6
7/GI972Ehh1G0oQImdaiQafEoUpVkZGXPjWFE2ERv8TI6ILS9qeYrGzUjzt7
g1rIbdQGLmnNDPFiFxfrZ1yAoXzfdOC1YHW9iunDnx4vAMhUaElbI9p/LTDu
Oy3onGJXX6ctzAtBTenuH6VmqLsD994tzCWs4KjQ+MZ9HHkmhC2NzmFK7R6a
jjlMkk1cJcd75r0pkttV9nhN1hd7hQAi9hnt3QZ4NYkVzOajQnxu6W57xstz
cIgtMEcTa6fZ7YVfKpBeDg4iqZDxUhPvWqXk9nnK/KyeHpOlE5P9SZX2tpHR
kA9yMoyH1poQHp6uUzGDo+3k0R8zc2SAHwZryFwtreyR+6TUrnDf4qMYtLRc
OJMknuK+8a8g4RiIjwJlvl/7V+vZpJWcWSOD/BKigc5DlYBRURnBelFWoqEZ
2J20+kx6qI7M6Nw1R7CGAEEHgo8/kephAPP8V1Op2XYhabanIFe/nXqZYGQi
SMvzOPAqe8HHW1SNiOIAdnIukfoCgsVhH30rhN2Clh6Rimjjb0OlE7S0FJDq
ITPfWxGA8v7aSKyk5PVhdzBaQpkcYrOWbaIGZkKbNHehbrP0iEKT++mNdJ7/
rjBt6tRpRfR+9cpHR1oRjHxHDV3hY+mZpmhnR1wQFaGH+RigCzZ1gjFZfFC8
xIcXIn+WGUFrM78bFV0ElxOOkZJN04vUp0qnuRvzp8zvKYP+VNsa/mxtkwfn
fde+ooC1d2Irv67vX9E5AcJpUpgtbeyfktO3ve4gQqHo6O7TuNOfpqS6vwdd
7qZ9flR5F2bpbleo9R9LQEO7WQUvKa42GUAlAgAC1fhtQTti3O9nwPFsU915
gCUI3rGsR+PzPB5kB/m0V+Sj93pFWmXLgSu2lgVBX9WsjDn4KA+9yMIzThdk
WSbDmndek9sZqU0On+4zmm19Jk9U/qwyhI7XeTcVt3FMc/CtWxngBI9HznIc
73+jphJHuGGnBH77KAah0Fp5AC4NGgpLOxlSWaeSYqpGkr6A9huixWuOeOo1
fXQdNCoIyAgIIsHfPnAGk2Q8vjMfKFbFJ4Pl3bpNuEvL8S289FlfXHyVeZlp
oUVgLmCr9kFtf3Jlh2w8auBGH4bnrVyHzn3sesJiom9/RrYmhI5AugCMVQV4
nTls1TUuDiz2VrVOZHuGaUhhhyyr2Q/TfcfFz9xZ1aNzhw/NEmi4E3VrD3wY
ZAmJsEvVnn3i/4hSY8szQGbBkCaG9+t7waoc6EQroY+aaDGMiIUqWEwz9kh8
zD5Rim7k8pa0FEXaHfplbsPnuUtoJoCz1x2pEqBc+PoZ5UYojTmuTDAdCsQj
7DmIpM7Bms4LyG9A8HVFoNVxaVCj7bOjtFjeUndyuqrtV3GTSp50r03wIndM
BJvNdiSD5bNWmb/4IjL2PQOp2Rb2bgSK+YClb7/2TW4+SIBMmjLY0M+gk59J
Wvq9V9MHmmr+H+qdEt7nCaN9EyBmbGX45JlgDUAg9AEkr472i8tBIYu6m9kI
x89tSmmjpyLjDtDLHdT0se+v9vTpzSB2+HOu20z8vaFUTK6SCNCLbekJjLqw
eF1S4VG8/88bnNx3Z6B7uOPF0aelJLQaRJwia8WKqknUdSYCyoZBUsTRMIFR
AmosGjf5xMifSfjvVy2ICXJsM4idi5OadInSnX8kYLRm+kwfGV/s6z2kdpVc
KxAyD8NMRtZQIFrshoMCySxLyGdsGIdukxqRsD2Jtl/mgIDhQbjGA1pCabl2
K/Z+yhVzFxqbkLopsY5XDt13ToTyWQdqZ/uH9JxW/stmHHgxdBTuOhP3BLFz
AU6cmIxlxiG7fX4NiI80WksQ43/exf7VyHExBCHwr01uZCATvccloHhhOrmF
Xw3REfzSA3teOE7NO8N3g+lGm3ETyJu1WuzboZaoPfISSwCm1nJHk0P+ABCD
3hhd4bv2Dw6FuUN4U+N+qwOYa3Kk92ETuyxbKmi9cpXK2ydhqhPeTSQAgAZF
FLDSJENnHkRTy2luZx8V45u5ULU7aNfsaoJrCktxEURsc1S+2TBKvOS56xQu
+UrW7sblXIFAfzdRLDEMPthxFpd/66I7kB1EeEyqDlHnp4jqI+Hcx3E7eZkS
VrwqAnNt7v0V/TIvK3qLhI+DVwYIYfuHSOQDF1A9I0JmfIdjuvZOiwRUlxq9
LAmeTHAkHBW3QlxchVjQI/o27GppJvkIDJ4uOclS6XupldHISVNpubKq3pbc
Vw7P/ilIa2tocW+izYHzXdpmGyziqjTjD8oUoZEBxsdTrv5wSO9Op6C0hWKM
XkNCv4LNpLoWNk9qg24lrn0sNLwGtBFVc9CC/uTxovW7PekeVZ51a5Gg3LD/
EfVDArRKEHEytaXKNlzJe8SMSNr3jblo6UFgsEUOQ4hHYhGetNGhKC8Xx9oo
PgFKhnsc6rtJQbjHhaYfmPsfkV0+fDMTqPBT89x3ZPQasztHQwiObWtLcFCH
XHGhO1lgaC01rH99apnDvP8i+oHh7FJKD7QFWmFkmsRopMVyyA+dIGowTkEX
TGZDuKpk7aSDxHgBwcPUpzbzwEl8HtJO5BS4wmx69BqGQlowXn1c5WbY4KAb
IyfFFHQZ8GEgRXr4fjOJ5f74IGOwbU3UycaKw8fH+/C5tWsDo1U3h3OZ8Vxq
YGCkpwvxW3yM5dCFEcvR95pG858BQL75uRf/9xbeLrcIKWj3Yu+HhONsw9Lr
jgexoEHIHBd9XoiZllGnLOqG6D4dNLUE5hS7/2SfUVHtJCXu+j45BMNr/v18
fUoxCaal1MCNLg3Q2xcVMSmUjHG5oXLw0m//kU51ml3n8/Ly890sJuwE8a19
R8v+kN9mgwaxN4/xtUIoO/xxZuR0aTBzdHSoHSkffEMoykzq4dJxWh1MF1Y/
SFHrZ0878z71dJyTciceyzRBzbh7G7JudkmQkRxoe5t1GIZg96R93ihPP4pf
Cx96k0Y5Ah11ex06DECKk9wtTq/PFW2civ5x+xGTXjhEsDDrwGC/A2lviuFP
edzQkrzkUD6jaBMrwS5i+crNAji7hm7AdDobdwik7HbDLUlb++cJU85YJttx
XzHde4oXxEK/kuZljeEwIKmY6DtEOsCBB0PT2m991oHWJhxUUy2chzR4sUFo
9QiBfOjEROD8iJV4Vje3VvOtVmEj3XLkFnfPY4pmFRfKY8WP2OyiyvsQQyRS
YcnuRIsdOpe0PFH72qy+HmEWPr6hF19Oe02QbM8tFoD9Po5WRXfgOS05M1tl
MPy+fMBBvkmOpBsiWAskXtpU/TcgB5Xe46O2Rr114SBebeQcycNgIRuEgBkc
Jx1l1Q6NalmzfhKjorymvTiz/rc4XGT+esJcC6WB1DZuJ9NbzpxkEAlSjkVK
pFAeE0KlynblyOzlFWpVTxZdHFZc5gnDrorofgsZJaUmA1E07xe3fCBpvozi
rwkylqOupXq25hgUw8gk8c6H9X0Zy0CoxqXvfn78Q8Fn0TJLoKMfXSff3IDB
HutyM5KT4Kcy+gPCfVLd5xbVJiALmquT+ntF4j2HzdjxI09hahOXo3OTUzHu
Dt5KwZFnk9jRBvFYcWOHPLhc8RtGJDeizAimYGUJnGxhrXabjfinPgwld3nA
BlpJ+ZgC8Yv4QzIKPnxx2LcwOjmAx/4Qs/OcRPzC/S46tO5hLGc0xr9UYdp6
W5NWevb2X7+m98e9Dp9ZXBlqalvHNOZ/4mcK6dz28WCecmOUpsgPJLh+3Uuu
zjz1Fi5xqmiVO1RpQLP4VTS7jSqdZEakQ/JJ3TFVQ3+O2JjOaQ0T6AG3se9E
teJFQEpaqQasFyk6vjSUWVtu7h7QLSHeGMIj5p/fMapS9OtXwffJmANCcfcO
RrxxSSMP+cyemxD54iTzEHQa04VHhywTERdy1ajECdwfzjRCBjTYntLub2hV
btQM2iIRo07oUZ4EpXA72fQuY5XlAkiEBvDRZI4Tg3gGwhV+w9l2jMTOMvw5
hCiqPVqMcl+VMeLaTp0XiblmXR9+0ENJ3CxNR7+AXykFjdEaJ4YW0tyQ9BgF
FPrauu1ZjEsOUEqvPnNdSnqZWt9R6/ZGu493iOPPJrtAWO5IyerktP6llo4z
C4WbfazspYu8pSIOUic1L3wWfvAIkezoHX0TcWTuh7pxvwRbaHmI+9Jj/IGe
CsYq2KPZNtd533W4UFOqqWr9IsYRFzMm3pUOFtxTg81hq0PraAnz6MqBmsCa
szU9OOb1kYsZg2RrYtgX6p0bA950J3AOhlzqrZimOth7u5X/z6GG+q+nUMl5
qh//5YUQctG7khQ3YqN/eGYv8WfPP+SO7npcuutfpqhzP8meydBrQdJ4OPqk
u4L0bhxrpzAaxJ5D3sDZ5KEIHSmZEB7hsSnncHljynhLjcMp4A3jQv12wYjM
yKBXtLvpnwjxFCG5DKDM44qmGCkokbwKYOFnPMLu6DDCX5rl+bpF5lfy63kj
X/XVz69Hb5oFdvwzx+8+ZaJc2gx7TbE2a5LsjBPs+NbUgEgjxFZpX1MhxTl9
E2gV11xJd7pz7D+UniCF0rqOyS/npzJdg5QHxmwFt9GlCPwtq9KwQUJTtg33
FXKkmtwR/kKv+pM/yeaamlxKuH+50NlwTFnTnPCOpdTr7k4quuefuQuj6jzZ
LyjQAWG5XwMw/90IpW56HfIMaoma7p/L+ByMVX9wNuc3RSTOWQMCD81JCYER
xtLEAeUlGDFlZIhnG0IzBOgi6G1Le4zkhmHy9NCaUSoxFwaLEq1ydAeoU2Tg
iSav2HE4qNEwQ46O8j0Vae7HqVZwn4/lfNXJw4Qqa/XTVRum9q0PyRRw3o/T
2EjEnzTBQA6JUD7wS7ybIZOBeWk685QWjFcSi6h8e0CiEg0I9xeX/tOh1pIs
3v9IwEuO+UI/rJ6RCOA1nfY88easMpxqDlapgrKvBXWYCkB/Oejj8K0xK9xA
aBqBsMRk+fU2M+aGXAXhX2qrzim4S+RSd/cwk9NSrhbYbE5VDLXAAPl7Avee
235zGuHCc7sJXzLROgWLuNUoVJfCIwxnunggv6yvfQRIqf3VtA1t4OLMLn/U
f7SNfs+xdy5pU0zhwCRcCyNbvBVCqPJllvSTynvpELrZm7hUoR2BiailmQmE
wdWCFFqrN+McCwie/JIB6sSQb4F4eOEPHlCMzjVxQ3+/QOoSIv3EE2G6W/W0
oKw8R1fZrrg4YZUA9gvMUrlOWNk9zDmvfTIVEyIFLGqJC214Qdhj3/SS/udA
EbKkau/8NR5J2o6gpm85xA70m/W2U9CqmhN2zJrMe7RQQEA+NjfrnGg6P2p+
ad1iXmcKI2HpzV9lg/EbezwupOQ8MwpyrcvnfphSRYhGHdi7Nkg6vZEy3W39
NTl58jaStY37DKS+Bl7dpivJCXJfjlcOVXNyRMw0wKKBkR2uRZ8bPcoso6L3
bkqOQhzIUxduWyuibdhfZf1ryRHXQO4cjEKkQHCRQCI+XMf8vPOwG+i7yJVl
shAmWAB879U/H7cE0MeMV/vQyeuAEMPRCLBUm8WaDSRI3xUNT24i3ZlWT/N+
eCHQoKrZHDQVHYsbgEzJd3TbWG4KN0qAdkxfS8bp1zD7l+IUDjOI3gzXxWBa
ozU+BWWoKg8Nq0L2AgBA5LjSzL6LCSK/SCfUaQE5a4i1t6QavinieMoiycxS
eWDxjMwF1Sh9dcfa9YkJ7mVYTtsHUJKGThdTKJDbstcCkEVR7K8oaHQ+4/py
2CCsecVNY66b/FY8IYahAQHSuRoymsApa0RoJtqLi5IZj52y9SC7b9xsf7pN
UAyhJJX6Z6QsIiIb4cO5LqicobWAWiEouv3Nuj6R7cpTGh3V7pNjQ99nfEAv
0mPkeRFqlawP8R5fp0PlK/yTfwc+zK91lJLSSej2brzQ9UR1skQ5QuzYJrol
PIORBZj1eSuaprkSDjCQwcAqCEi7T9bjWHPco7CN9+9dMKo3OJgAZN8PhF9r
tK+vZ1G2qJWuLSfi2Vq/Jd42aoeP5qJ6V/z6mtiBiJkh877DZVRA1UXwWLpv
oInDvFfYsZxL8ZtHGmTI0gWkogaThDngAFQQUz90yEPNMWR05xSJucYeqD8Z
RWgPL//cHPP1kE4hGTy5IWViHveTXzXA+MxCqRhcyRqP7hwZw90k2lXyFPav
RMnpyOgkXelGI1eOshmgVGkx/SJsWxUu/Z9z7CEt9CXUB1MJQdV0/uI/V1wR
cMFOTaa8ChkKV2R6JVADk7eqkL9n8CHDNonKo5ERTPt7Rj5H9e3a+BnZQbz6
tl4UCa6oTLUKoeUMpy/8y0XXSwepZhGplUsChPtVO3vk19bgyukaTENjiwLZ
Hf+48FP9l7+CJm7Lnxzd7HsK/xhmKHtkdTjff4EHZ5ZtVkKwDGM14u0Tkhnp
X3Jf9u9ZFoMK/3uMyQZb7ER9fUGkQ8pDCHGnv5hxd+4ksZ2ch401KxDc2R7Y
SQsaNNvlZhqenAps8v4o1FCM6cOzirIpxm5b9k038G6GkULz1RpJox49R3Ix
JehK9gcZr3lwA55eSzIvKx3TlVZORL1rn4mKI7FfOv4JqD1ennMj4itq/V/+
u2/1poE0u7Cy6xLvDWgAsXvzR0d5T1Ry+Ae75/NBX/Tt+qRFwVBH40plpGJk
TM+QSTkF1YUhRElCs8UPt6LZYGXFJNYjU4yjOi7l4CXh+bq0I5Pol3SXQidu
LeQqQD4AosW6tbdUGQendGcf4YmEZxzl/OZjtjPhkmKfSy1XIB9wVM6v3bjQ
JvGKcAKclNvybhwRDmlRKwD6cHIvQqOPrBNXU4gnReUxtlGGSFEeIfHwS52/
VncCT4N2tSykHExcu3dlHHmrUXg4rRvrdaIwlOa2QmBaO+XI/4jUDqHx4X2h
uBUExVZ4TGnawAX5ZxzyhjI/iWUVLEE2+ZpSjeSSoTQxnagmhaJNm2mj0xxf
mOrud51/k4zIIu53pUeYOm3rhV1ai2sbb8ciRJhi3iMpEi4OpPbfUAjEhWPE
qJtS4s/85gT9swAS0nn/6/SNt173TLBPtbKAiQby09Vtf3Z+BWZixxrI9yyD
tpSgGEkXlYp+hWBuRoVfbvGMgb+pdsy1/PHFrWbSYyGkX7PSwy/Qnqz3LyXm
yTG7eoe8yikIT1ND0DLpO5hgZu+nm7nAgjOhXE7B804/UiCY2qyHwpn3mHUS
OmFq+NCDK9chm0deN2nzhqa5c69glMLflZctOjvDaT/zStTQtbSGUdGoPLVD
67DXC+/DnHwD4F37Nt/io8CHUH5pSEtz36PrqDV9Bx4qnAYJTwb6HL3/kn2P
4EZJuzSw6jI/hMUyi7QkpuaAvb7h19K27FyyB5tEKHeEWwIS2DEzjCsTHT/h
UtpHNwU9uV8A7ySksNDOfUGtoGhOIc6D1Z9if/FLVeHITdtuhPMZnJDrqSj3
A3CMWc2Cko+yCfDsPcmchGrMUGxtgzz7BnKJUrfk9a2x4cRN7XIYcPHehZ5C
7TAjEpv35y+Rpnh7/KWl0YlDiXCfPATmx5gIOeWktVb+cHT9/rZzaxkanDeC
VvhyE/cL0jZlcQqOW6fso4c814Rq8kwopleGkGo8/yOruHvu3eWOyvYrTewe
FzT5CrfHMYzABI4E3pWQn7oFRf06rYLsN3LIGuRi994QFVqIb0r6UtLRx6Hj
SPf/W+1/nzaCABnDkig8yrJOF7y0O/PXDao/8KcmijraUuWv8JdyGlMrQ9GQ
2ZlD7k4AxQpa5KExgFThnYKEcZHIMZ6tcNjyCdBiURIGDT/7TaNOZzm5km80
6zW5T7s6z1AMdFrjBP3kc8M0fu26bYNBE8QCh8KpbHbB5pkFeXxfkG0ZB6ra
/4a/av7JtatDFCiFC0D4eadRGYS4sxwHzSMKvbrKhSgILvyFdvVhRt9kbn1e
IFlcmRW8XjV/UwJReC3uWgImEv8NOqDixx8iYzknTMsMSf1Kvgw4/NBzBRKG
7l0MV01Y0kASizWcx6W16C7z5g3fcU7Nc5dPwF7/bAhB/CIFlzbqonRb1Vod
3Q/N2dBx4LASpFZITOa8Gv/ugMptcukrKduzSUVTZeGwBsbRek7kzSkMfCsW
hYJJeZRFauQLOsXomXppxifim73KAdxGvRGyTBY0wg/2bYsMh+cHe1CSxYLh
IOMahjRtwHeYsDYr/3Q9hJHfFmT014icgnRVgIopmZLI729QuCPFEY55bVfX
vrR4Lws0rLUf7u7piO6Bli0WlOcuneqLmfGUqmGKUhEDm0Z+foFztPH9kR4q
yNFtd+gaxlcOk8JHEoqHQN04NsQf5YoF53rBMfuwMk2QuPbzLV1fUloPhBED
zhkoQ2WYOT+C6OzzfL95NFIQje/kAnz+61wEjBTiY/HbfvxXKoRMc4d/SO+g
ZzjlT+nqGS/44DhetB1cgUMQY/pv0TXbE4hJMWBVmCFvq9DYPd6Bq05Vk97o
WTQLG9fN/xN15MJoU5GEHhRh0TYvyBVfWJN1LwAjcXXDd0SeAcBuWaTFzsPD
142u9zKaM7fxyHjZWRB8ADT87QySys42qoF+eJZ7uTmbFqDL7PApiMp4hpS6
OIxh+qxiP2y0qQ4LX0poVW7UDhzF1YszBdXOcXJloVksr3O8xoeHQQQ7Cpg+
yha2CQg9nU2TSRxd+TtVxVR6AM3tQRY8zzs8MCP2Xd5iC3sOx5XOWPuvsKE1
EpcavwmDQGJXcWZdvXSwWKM9TzkjfJ/EUEJkqB68TMI1i/drZuf9myw2gHpH
BwuWdHB8FqcUbXu7krIk5GNbsA0dGDVspM69Oh+Crd3G/7GQi1OQRjjvlLj3
GXphOZLGpAqCTgDGfL4KYjOdcHNbzuzcEUbX9Z7XSnJos6x3swf2jug8Arrg
B3J981j2ZwOkR0TVRHQQ3hQ5iEqab4MZvIIaibwQjTFbascODbmzI+t/qq2l
E3e4/V9a9Bh9X9AFtRAM1pB8MpS2CPr5blga3WCNqmxLGDaE0eMJ8eGAye8h
7e6xc5KZa7t5LT4xMhhzFOwbiHMsZ05aBEPrzpwQ2AcQpkOESIu5rzSQ+D1v
K6/Gxo6r13D30IE51dLkYGkaUD/0bhT48mF6stm2jIUA9X+VqkLGjvlSP+e8
trkhmGMCOJldLs4KH9PlYEqFGPIkIKGQ51fvN5YSEDStHPRSfGcszsN2KWEu
b9wfqGuVHHNETLVFLrXNXI2hTAXlkcUwkWtgtVENTV1F1plltBVSR99mm+2i
G60Rhj5HVCt98RyBmQaUarAyuXXvV85qkFpqTQdgV5x0p9ulgcFY2WNeNjYS
0273nCYB2c8sQN95GYRD8ZrqukiEdPZiR1aMjvn0Zue5bvqzQH9S9+pEc4xW
ACbz+8VbO0TJPL+VRmnzeH6h14vCL2IbfObPOMUO3ORibZyh5ZHa256oKO9g
gGkzW8/oRtLPukC6EIZkdevEG49W5VQhZEEXegZHcyPEYD59jIN9cNKVgLDP
RIR0wB+hok+oiCqmzvT74eklkaAkQ1YVQ0X7pSormE76Ew8I/uTVlg669CKF
MFKDTLGy2UjKSOU8sUUzbxrZbvk/m4SREvEQly+kh27NO6CbeW/m14eTU+5R
TrH7+olZm7YIpH7QKphWqbs0tvLjG8Kte4d3PhqSI14XIzvBz06QV47qLqk4
dqSJlT8fckK75NvZyreEtmbUSjQ055h98qhmkcV5wrXHWZ3ub8+AS0aTs6y5
il7sDoGU66WVEkt/uqbeMKvQtmLx/wDwdPAqA/D66xdqI0bvwV7vIMeFQR31
z5vsxAYm+QbBUxF1a8NlKXgfS511mSqthEU/4wD7svB1KHShZQJoWizaW9Ma
wAdI4UWz/yEhjbXmAzqPTsNYKUTWVI9rdzhnDEK0MWSL0UaLhWfDgT7x86qE
OYQr4s6ee1bbxRNPyr7/GqiuarX1OlefPI/Djj6Yru5FlHdsTMxBmSLUGGa0
b1Q1WbidBj6+RISEE8KHNH/QhC0pjc4xT0rQtGFfN3ALGa0F4dFcZcdNKgWN
XjsQYSGBis2oXvyOlUwY1Y0xtvd9Guv7ER9++baRSBmijfCjCDtEfkDIq/Ly
+F5lfd46Yy/VKUXuXFKS6Bvy9FtCfL4HchJOGjXypXW05ATqNITtINdQFIk7
naWtzH8aP27P2A4s6PKEmQaBa9if0MTKuh0otzLkh1l2KDVuK47Ox3Q18NgA
96eGwLj6SfHAeFm/CEomt0FOeiISU9/OTuFUjsQwX6sXLrNSRcqwZh1MNCpR
JVGE34Dzrm6N6bF6qZHy1iKs3QggozPUaUUPOWz8sZsEr7v474SQ7qAr7eBM
w1q56pGBXPMt/LfgHcZu/ZFlmTM7T1z6jSpymgoIvweS7e1jpmTyN5fHD8u8
tL1crN8DHOsuAbOpGj/ePEtx7nzP+fChCqLpxVN5GAzHOj0E1/jf67j377FJ
vxJp7wywtFc2TTIIkoysLINjrpHTFOmbpoz9cceSJ1Zb5aOtmKWFWTHeqUDc
OOLePXQS/lSUJzhHcNHKX7eji2AsJ0yzSBYL0JBxCQIMb4gXnFppZ1N3J2NW
rGT2JkmTR52gCaBxaC9boGi06/fHT98C7+ojfrsZRkRPoHjj5+mWYrWW1N/H
/uMrxOsTnFmC7s9vRM4wgSugJZxR5arYhOX69sBq9XMXlXj6LzgkbRsjOpJx
KqLfeicUfhY9xeb46AoTzx5fR+xRMXod2huE2A7giUfLHqdWS9C5nG1+RDhD
Wzo+rmer3RPfH6NO5nbiCW6U1LiF4OIeeZ8fmLCBKTTauiYXZ+WHMaNn6u6h
xECwdIWv4e/JpJlT03Y7e2TZ8na9LE2Ow7/UEJcQ5BC+MhQW9glmrPVAtcwa
+UGa/QNSvt+91FrzZNIWnWVP/GRZjT47XaJ739d5lD8j7o5R4x7UXSSM1KkB
gMlTQfjQsIYovSNFhqNF95yCwo4XVzksbFG8LuXMfW5s6fCqDE4lrKW2vPqL
7MCe1VYinnj/sx2ZWpnF3DfWrZsPF45337gl7AQ/vkqi02LHnOgzKmvvaTpV
L4etLjmVyIrw9XBVNEe2EhPKdhH0Co+NfR/MyGYzEjmbk4wtNIszSq1bQ42A
f/wx9vmWrrOyf+meBNwSd/ksBIlHPZ/KOTCFh59wAy7i75keo0rlVLzZgRvP
tgNW6CAn9FanvhzA3aHKPSWIZIcM60SALuTWSJf3OnfY+Nbs3iOWtYlfbeuB
KL6pd2KdKzoQpiLmTrv7mR2nPc7FdvRfEOrmPF5SyndrbQlvRoucOyZ3A+jh
b3eD+n64ZrNIfW0kx/3pI5NNVWM8Ym0HpOPPa+Kt3ycurSxF8B82yQoonJT7
qOtk8G4qQvoYDqrGL5hAj8h1epVV53Kxy/1oZmnvECJuOWXocZ09Op3IwA86
xLPaCMlZAf8A6jivQuKejdJjS+XkEauW9BnyQLjN0L9jcvUCwnsiR5zO/Xtx
MvAhdyvGnK+KDPKmve/ddv/A/AjX4NAWG+LsKA46mzKVyzZYetNOhBHAH2ar
IfS08TxLCU7HEMjRfpZqt2vo6nT9Abui/W/uNHCygZtUqXSaooYPFn9RNHs6
KsW3i9mfKUDUrFphH+ta71gZp2LpHKh8MbnMGLwu1r6H7u+vht+yoXdYG0PR
msurff509rVZAl2+Qcwn/0c3Zu2RuAdaBbuQzIYD13xBKyCjg6j5dEngY6gc
jiDat4lRUs0qRTkD74ZMwjvLhPfaV+k5bwXBTWiPPn38g39Rg7O6BIHcHAeQ
k6uFSOmlHIdC2ZQNR+RrnI8WKuwoUcc2WN5CyY66cUhEg4t/CC/R+7gscjBp
SvIBuX4zmehe2mhcItGmePSGstFLfS9BDFgQa0sbto294HTbtiX/XH64jydQ
OnLitsglGAiUi3QH2JjmIMsX0/u/B/ieUsUXWIX99t5D/zp6/F9vNIA6t3e0
6q9dPnIqvbUU50XM5Nt0tljuykm27AqYdgXFZx7xaivT2BUbz855LIazP4Nr
okZTasN4SgYCnbu/Qmp5uao3YoCbAG5aUGC1XmctkDUg2iXkWywDcDvC+Syk
t5I8RPi5KuwJIqweT30x4TNieL6D/2OdDGPVv25e4Lppe9cQmEcOQhe+yAae
bavl/8IzxhQm7gQ9UyO+6i+8IiBBXDpfDrHoUiVRUnsmbH4nbbVwrr33OIIf
stEI+3InNLix2y4Z90V4iiv+ZeEKkakW5W5J+/IrTNJzPZJnt/J1KQMbpONM
JPmirSsYSkGD7s0vgJm4z5mj61ai1G47zeU27uZWxY3iORijfVwGAQQQdlSc
D8kW4PpN5loa/W5zWuCc1QdtvfzCzM4TbdRtApLrwgfQrBf1dPjKe65fkOoj
ysyBqWOHcpD3aTzllFLNBNWXf0RsbnIwQHZ0a31qaZy3bYAQTs+0Wz9uyT3P
eSDpxds3iTxcWbHKpwFGNhRl8EnL59B+BoJtfM75Bb028F+lsyTl37zzeJvH
PT52AmGob2t5AsEDYmT8NOWlBPsIT9F/8mLiVfcY6/FqJDJ6rZ0shi9ZAhs/
zNGt5gOe5k36aLPyWKLgNkwvHazqH4Lmar+MMWINim4TVLk1hqMUn0b7ToE+
tToelg5H8T8aTef7YdecwmCp/h+SDTBPCd9kzwHcwzWssF3wgW5+gY33/cyP
+c3dPMjcoktwTRaQHYLTIzeIqQsORQtuss7VVvnBxiZ6HQxqvOFL9pSXjJ1/
h55TPatLrpSiTCWCWyxKToELb6zHEFob6MP+ZYPTwZU3gZNrahVRKmbaJVrV
wizJD5+Qs5OQ8feZEbGOeac/ec14pAUej7swrVhmwuq7C4LSPR96jlwR5+zl
rY1hm6N2cMIWmwtOgGYYW/5Kfh6m/3KDEXK3QGq1rpto5+UHX2jXS7PTgwbj
tui964zhgHvdTgGutplelt/gHCCdUGA2oDsXUD/reYVnYo7KpNaELEysXls9
z5yZo9GudwUmbwrIsFtrRsVOKbvOJZKH2Ik1PRKL2CtXVOqONjC4nPFX66VV
ihEigmCyxWZbhY99GzAirOEhvhKOSErrPU2flfh+ZAUANOgOG//aE0PYXjSU
nfZrKmHscAAZWFuecYxdol/9u8zXsNO42ecano0WupIdMuy0C7dCeuT1uFyM
xyW0uFM2coH/NPLeH16EM/S79kGtPfdCpbu/mER7LN15UyUl5Poute0DSABB
xxZDmKp+JaYIZmDBQcltpZVBd2dIRL15lpBNheI1dvKWKq/z5APvuqH5AJ+U
Eg0nCQ2JkTFpcdBornOxxMU1yXxb/N4GFin27YWPOAXm63aC3R9kfDeEEN5q
EUnqzkwSZFbifcy0sNiZ2kV3h0VxgE/sk5clglTnU5vMH969YdCSAh+OcNW3
c5e9FxOyYTz05yCeFbyOgCRSDMha/5ZKvsuuYwRnS8SDv+5HBDUqbWw1UCa/
cWNamxLswtP6q0R3NBLXZ6B8Puqjmngcr9IeLJaXh0bJvN/dg0UhhYayhbN+
vXFBkYSPt7W1VAblY6nYpc2Tk9gjJLfYVGhIjUSeUW8TSXJ8mfrws1wVEF8s
kisLa9BA4G8y4pgufyT7hV94QxeIfpeTz50CH+4AD/+fM4ekQEkYvjIQSFJ5
DQWMl6jGthN+l+WS+7Uybm7LrTKEv1+9yBfUU29OW2SdlV6uDjYjQMwd7ioP
vn7sCMQViPIMzktOyzSEq0iNC1v7zz7gYcXS+vNftw5Hr1y27hyraCpmN2hr
h+V5KXZYQs21xd8rSpI+KykBqgblPImddtHaJR0svIWMfWGOytqVPTMTz4+4
zrl2p1tZ3IFtJvmPFS0r1R/dqObLf3FgT0QQxkR7aoID5oiO2TUjdYrbWBPT
l/PGbx9DSLzeNRKfkiAGmWKJ4oy+7NpbM0WdhpqlUSYHx+ccsUDpivIh439p
a6ibt8mb2e4EA7wDxVIX1k+zqDzlguC8yExhGeOePIRadC5s1bEIQeZRXRb6
5mOL1Zo7aoA3H0q7oAF8oszPgC+E8FEZmdAmjMVcivgWSHWk/wJKQ3JFQI4B
52mTII++7jA9UdvSJschwbWBavm2Vq5sOr5ul5xgYYE0WyxLpGSjVjD/guYR
T1W+7bemQURMJl83f/lS4CZ3iZ4jga3PhEZM5DfjOn17Cvg9XJF6IamGN7eY
b18x+iVuNsEgd08dORbFlbvj6Hz3nsApczC7LG4EYs+q8TfAoCCOv0CGuk6y
1w2h8EmFo8y9piom4K08dyvpF3XH5LA1DSs9HcwRrmLxLWKsUaYS482B0F65
xMxXTjfxw24ny5PEBfUUxAhMyI9CCYG2HZgiysm+ZcXRf4cRtbqEUMDKPw0i
fm6hUefn9zXXzxTu8/XUdHoRCHAej3aSfhmGAco/zZjszyMOLKxYtxHTmDb4
YK8VVj3UUbIHqg2yMO/sPAPXC8TBA/1RPFnNRL3rgM0Gi76XMSujgYiXvCVn
XuWbdadT6TghjuBryWt2OlSbgzQ4Q7TX/ZlXJ2rkm0ptXvYq2wuNIOR8W2x9
z4d+SIqA9efvq7/HMFkkYYuN9+qrd66D1DY7ezd/Wi9HmoEtLpebowgzY8J1
IakQ2VQGdy5/7LbWvyUIWfI2JH+0Z9cqpn20VtXM8y6CC/NJ0hzt2Y0q6Be8
IIZG2KYDksxpi1crCY/nobykilAZmTtnFB5K3TLScZnyVONmwmuqeFQcllGM
nn92Bc/rMLYv/Q/m1PgOqNXWERS26SasRROgWyD4ECAsMKcocDwCOp5S0Dni
kfWW5mNi51oZDvfsa2gF7yTm5hmxX7PKMfH8S14Q00FWfWQIgTH/h6nUpF3F
eocoI+1Peye5JbGaG2+xxndayPDgzxub+DLcRgcojl5o/eJppMzOn5nd2vD3
2G0hjAWvWrnmaJrli7wyKv/TwrpaoAliTWdAUMjpJ8M7Dyf3IEnU0nnyrhMB
6kxHAyoigmUlMqCn5VIujrjD1BBZaylYYTQGVUX05uZIPb1IOo4VXEwbfqR2
dSJPkC8zebdP4DhXiVV2sXEsnLDN5XqTJthxlDBMvtx5M6m6kbVgtgM61C09
jRXqBjcwGrnmUanu+zN6u+qO5ygZbFL3QyF9/cJrJL3ny01TdwIQ1B7n/BPw
slIi5LcdH7yP7KLKc7qmTBqvdnyuPaAQYNOA+11mGCjCi5dhM4hFhU+Kwult
BTpnpvPheRFKdp2Ih0tBQArtJC4LdJ3uF+7runns/W9UXCZWtOqCS9I4bMLg
zVauWNMozyHs8GozTm+ZjEQlLBvtg5n4JKPF4pKyUFNa76TWbWb1yA5ZsC+F
l53gpn86HXGZ+86OG9mfPEDEL7yMrYr5cwuXxzJXf92KgnKKKvxj7BNYH5r/
SM46aS1mbQo33hiK5QioOb269kydG43itvgr9WjHwDmZiBZEN76aMXI4Bt1M
wfm0YCiAWWPqk2BnaDi6h3+gKxBQ42F9u4tHG3I5lfxA+sghVkpGq3wLTgPQ
LjlY21OkLiciHi6LmZ5M/gNpBA7ZNtvV1bxyYtqhw8aLpjfReWjyIAZLm4Cq
zgRJZ2k0quPSfkMBwCsYnpVEqk8WIZURyQO8m5eHsTejO0s0cyLLZ9To+T50
nZOyzPKQHZ28V+QnmEzMkVd7DO5LaGdYi2P4+LRbSO3ScmNIyKgveHaUAHmB
SAvtdx3OTlb/vE6wFNO4tlVWnKMXRmrNWi79MMjzL7gVXnGHSSx4Dnn9+mEZ
GRX2iHhN/G8EcxKxG6cBibHmOUT7MLP8B3/v+IMoBdMx7srUtSJhap2isWma
c0kXsaVb8x9N/1P5pHeuB2QvnB6h9YM/e+YG6nO4y8uZV4ZXxvw0oOH4CKWc
LBuoNs7ccDsIRqVJ3qZaDKaRREtiIrET8h8pd8WM1m3+fri3Gny/Ht+lj/ZQ
2KIav0SRI2cbIJWOtRzZxcJIVmmJorar5ruhLjMUFj2klnbkinGCXbLhEXze
CoVG10c5NblxHsgbQmeean3WAcwQvGQyltbsobyxI/+pZmEfoZpwJVCw2RM2
sL5hJaZBEP8dM9MBaLRJzqRRUUhK0Iygtob+CtlbiCiiWz2ukDFBqz4o5n5I
pitTeEO2tvgCYY9oMnBkNGmM/TdOEd3gkb0sAq+MnBJE8n8hOEVITq1vM8F8
He25x/gVSpoeILcJ3d7GSmKHKnPPRI2fG/aPeVFkuz+KIxAx5OeoStwuwZR1
xe8y/n/+VlAvlfvm5NLdtvAPIxtFcCykPT+vSeOSi5QeWiVrdb5LtiOuLd4I
oPcvG++GZi7y5X42jAug9XEwALizrZeCozt2Q8uqLMtdkL+YFzKnCyTScX+S
HDxVsCwCnYOKpI76Y/ygKHtufYnM7kCNhcK7EsJebwsG6Ux2N6n6hvRECIOg
rFSPV3foHHEO93mnjQVAsrsZj63/9/0xkWLugE/TkinsXDY3PnOxqRNo5DwT
Zt0c4fhP2jv1U8YgBhJprNcBb47FjI2VTfWTM3OM9ldw0U8lCSd2RDllQdqY
JpE/qJevlnMF0awsFmLy7qa4RUvJ89x3IR287q3Vf+ysmDmrlz+Hk69WRgyp
kwdi+KvkPMbneV65L1hL6C+ql/896bEv1FbeMn4DpcmHa7pCnt/Wn4ogBZ9l
Trz+bGQRkXvB29IomQc+nDCKjXvuuKvAsX7cg3l9lQO0hs4k0bzp3ZtViNnG
ohxeR9YryU4p1LHlhzdY0TS4TPqo4Y1W8/+zQT8ZygsA2PubrIcYnHCeLSYx
RHqx0PNHejqm5mARLzG9iE/8FdYc+yBlBip3W/3sE3GqiXrdVu/Ojd5XsmB/
pqd0upvQnucEuzLe3yrCX9J6LQ1nbn1+BUU0gb/aEdoPs2oh5yZjMVPINaYu
cbDkLB4BB4m9M+7s99/L/4AoYBMMpmEv/Y4i6InFdyDNcIXtgYELhwOa4CKk
vc51NZX4OXPSUgOBwcqT20fwd5w60xst7eW4lMB9ymZNVk4T0ySo/1/Ym5vn
YPv+l6dMCNP0vhR6feNpdQa6ybGkvkAulX5QU8rXFWH7VW+Uert7wWgA3PJz
WFR9hGq0rwzdpbBT6WI6GkVRTlm6it+UI9v8VHewwfBZlCAvQPKd+20jDS8n
kwCE5dJLw8nJV3ptdX9WLmJA/MvAXkSxUma20Q3yYaowtVE1GCJilx23gFgK
2r97fWbgZQdvLMUP9p1tP/Trs08qElhSoyp9whP4Q3EoXCAZMJGu+/vfIomm
JuP64E4kI4cT93icJA5fGA1H60yNTc/Ue7uQGFy4ocB+LTU9f/OKCSW1LoeV
F5F/iEPz7voQkqgGIru6RcDoX48aIEf2CSOECSPrFIG5nvsNDvT534soaq73
yWzk++Eep9CwnTzK5fZfzOxelYNwBdzs+GRwQEBCNZCRq/U3p9+vNuytXZ7n
uc2uy1DvLNLxE1lpiAyNALPO6HPFubNX3CxqwkSa4ik/DNu8sF74Od3HwORh
AbADHzaf6S5gbmr+b08lJ6Xc9/RdU36Y5iO1Bi84I39eiaG/F3G14HB5Q1Vk
4gKTqYyqLlk4LE48568XbQRloHZ1dQys5Cxz2O3vsQerzADz1kQX3eZQitMS
c6vcgd7uynGYCCHgLId8X4x+8adwU5dZDet+76GdcdF7/eEl/np1CkdGq6B5
45UFUlbs/W9n8Zvq78UDduOD7LN4nxKpgluyvKQxF6zjE8B0Kf6R6DocB+R3
jhhOGLjpzKyGYyjJUgDN5DlAtUn1A2Stb+oXwLt1hqgD7RbRDtQUCtoGKdsY
qhAZt615JV9dshkvvBx2zJ+/CpXqc/JJcEcYDC64tHLo7PIfnHd1WevA8rqT
VNbOIkpMBssKA+2MlVxnV0zlZdbFD9f0C5mJ1YFIj9GsT8SUiZRZ0j5L77VB
/qq2GqtcoFy/M+81C40m8vp8dk/QdQUJygiwneOi9L4ffRjACsrZoM2sJ3H4
8Q9vbKABM7b24WFJM4kgjYDexnf7utkoDxfceos2ubV7LQWUXugJkU9eTMjt
xuZ6bb2a1U5P6uSdq1BFDSXd5DLXeNsDeTyRV0g4oYwomKplu2S7gfKg/+DW
lL9/uMPoPRhESeKSzFRp/MdHnQzO9tEPfx6pIPDz+hi7dKTYOns0iqAF1cQg
2hzywTq+csT6tWlLp2t+VrUKV36lLjoJawPwjLSeVFC78vwobwdoJDqdnm/j
qGBr/vENHEtM4udkMZqYT26kLWIc6C6RI0zKTjtEHEdIrwfnLjjpIZT1b2d4
fCpb5d6M1+nqogUarMbY8xcwuhlfgAoZMoIqTcIRc5fp9qyN6z0PHpHhdILB
H6ojyuQxEq7FWz/OBrXg7qtb3OTFlVdu4G5jgrNEVLVVeHp22w0Dg1y9hoyJ
CmqqhGEHh/k7eFBGBmrJDhgsQfnpzSTcpFBiGkI/qE2IU2lFyoy467cItmT8
57XnfvdZV/h5DqoNll+aC3YIGCQ4W5HcRtKHnPbR30VZX30BENOFnqLOmGI2
qVuRTDNwIJZbpzAQ+D7crWabOG4Xrkt+fq/WAs9+gMXoCUxx3otRjXaKE56P
NhFO3XzggG2MAsNBy+XPBO/mesS4QnCfUpWX8FdwMNo4n4CKIkQPHPwhi9rj
HWvstMayAiP5HuEJ31FtFZ9Ir0ggtqiOvvudK5I/5XJa24jyxve1Kaxr1uOi
yISangtn3T7JCXeQ9n3yKWTSfbxhVzn4oLsRQoXBEusuRRoDPd/QGYBJBZ2f
Oz1ALhtl/FRPfVxi3kl4wxWldV0azs3+BJYFnBTMQb3jVoWtUPURyaWvwCUI
Gkk6Lf8E5DcVAAqLXTXOKK58Ur9A8fHWNfGX4M2zfQM4Rrrsc7tFw5W1j9GH
nJwBwCjflMRwIKTm8eeiJptU9kIbJB047Q/+BtzNZoPbYQLZp7v2d0Ha9s7x
4ovjoieMknv95SSs1VsI/NTZtKtyBCdyo5nei19IeX9CdPBOQkMa67omb/pL
8ody9DLyqdPrftPNnjZNTE+Lk5M/l7svb4cg51q7AwR9SbRSDaD0TWSa8KGq
UApZ0JwvlC3ygygYhtQYM+UqP7lyfbJE+UgHL329Dq5gIh41TQ8z3HImc7cy
QUt+2PtDtQOiWdkw9PgalAbSYAR2ieb04o1Ul85+Yo0P36Ixg+rCCNG/EwKD
dcEyax7Rk8hIks+Oy1eVyArR+ZSfxfhNCrS5kxaz6IRM1cZXOFdmqDjo6KTl
OZYqbRXEwlhmEV6OK5oR1IEJ7C6IPCOpkauZbfmySxAvun8Q53HZWblqT559
uhaDyleTENEoFypOwiNwDamrCclwVR7FjLvyUbLh4Orze3POrL6vpRIKPNHF
DkzqmxoL7xXN6FsvInriULq62/mHz45CS1hXqD9qpx8Q7Z/gqmLcF5lFoIug
kEdkvJmmZLKyu674wgevy0ZrwvHOKn1yfdggRHxIM1jd7APn2NK5zt5S3c4v
RdgcfzFZNpfHbIQ9a4GIlNhYVzqEAWk0fUbUHaq9PwggNS2kGryJWAMlIozW
6Ae2nJzlBZQ/e7U7xR/yUMdSpkcNwHEswGPYdARwcyHxSWO3pGC0DzBDloig
bqTUpeE5dNrR6czxHHEdLMq1I1pWncfQN5ixXRUW40gKjJ4zOL21+NfBiyye
kljTwBCiiR5g5bHl+CmElqkJYgzkbldpQmIfQLQfn6EzBcxOmqOtPGfbv+6R
/MD16RWJ/YQpWJOiyj5mIrerIjPPAKon5ri9vxPwrLqiHN+8YlbhxVemjqNN
NW6zDOe0VDedhsMq9yxFq605J0RoezcBdjpo24HTUQLMtqh7s6TvOyrgtMj3
W5TxtqeeVhkdHGv9ymIWl8V0PS4oORVKjQDiTv05XiJJ4exnfpHfPZr86Hjh
2RAJreRbfUKFExf1bE00Tqo6/UeW4PnV3wOVw6KHsvi9uKRfxPnCoR6dtbbB
sMQQ9wfLZwoWSOmBCyUYoV3BUptZfW7Spn5Dn6iqBxCXugQxBn2yt0OM3q1m
VYBwBwNEfhw4Mq3txy5bYmmfeNiuCbjpl+OpTqPSvmQntswaNIhj/g91bbK1
THML9718CAJa+JXXl2/cps9zYAnXLAyw7mOoteg9cmJ/aZI3VzlPRvpPEgUI
WjHdmuEL0OYDzjlDsBmRGjVbwHmUH9vULxXU9Z8wwmceKfZzZkVdw1NZUpkW
TfbXZ/nStjPTccQdz4OQaIySJHjLI0hM1SG4wvjhoZaYS5r47sF/kLdGnJey
ZzrT+KNeejoZocTbyG86RAW/PPqzoGgfe6sjk0KLB7zfBuF0QdlVDSlQg/d0
RSGz6uZeNgYpqArk27TNkaEx3UPVTTOxe/a8RPjvp80YV9WwYsLM+2qnwJeW
MuQOcY5k6b/1ppYbq/j6RsB3f0TOKkeS/sT34eBbksqzwrXBnlxVsuvqmdng
95DGe8CugystGrZDwMEMN/ztJve0QSCXKvVTTckfUlYz6RLfuXooERqoVbfb
3UMfMAhgoq/ePBbf22xckHj0X5lyL0RwTsk4wxIYY5ohRbcvZtotSuAamOQx
VxcaMZAk3fipLH9RVliHql5swJ4tezF5qOS+iSsJSzu/sd89SkQ1swPVMfqt
nfr6D6znQve8OUcbdZHAxW5S/mc1/oOBxrZGtOtRJ5+I6nfhAlERlHsrr0TF
KMFpEaJq7rOwEOK9oxkQGimiMCsnGdeRd6d688AWh8Y9CdPZBSJJbgmFc8Dv
t5LaVk/T68J0XNsjk/oNn58HY65oDe9MXzPkYVATdEOrVBINvZ+qpscF3I/J
WAwOssX6Ts0z/oG3iTI/yTQjdy6JxfZa1Ncqja6Djy+hUya3UXgTpSYUE6Eu
lalnyTLC1iQbodtwmXQhqHYbcEHiDwMoVj2qCqjg1/vQUaN5TZSkBYO1c85K
u7h+vAzt0rAiXrIUKdr9cQj3tPAfIy0R3s3mbUGw0DVMME0ITuY2jCXal7nN
f5b0abEYSrp5XLFW+KV06wcEeYJwRS8hAO5X6jdPX7jo07VLjW+1bA5IiN5l
ZwxhOyRy+rtUJ4anYnHt5IFU+4XgZVpS2Q/JOgGZHSmvrycxQaceSHqfpzFW
FC4uxhV+dLMC8Hh/xe8kNOK5BhjSTzLfbwMz1kOSlnJQGNKbRdPTcltE7Q+a
vUw0AskErRFyo4HJOq0jj+8zhKYAibwnrbNvZ0l5G4lYVjZ5FmCr7n5qJuso
FTkTjySIrHEF82tZCrjtALkO28xU62lveMebqaNmORUikoRqCXQLpPVPScEw
vSiRXYMQCFC6BzhdS27mevUWrOMlHA7RJ2JPhGdlOMuzz/CCaaytikkDyPkq
TReET2e+h22WNRpOb0BNZeEgW7VFXF5rffqhVoAixtoRy2TP9YJ0SeHIKyxF
qCLjiNWmPmgTNDagUByk4LMTueDVlhNNzcd6yigkSkxZLyTWeGB7lJoutSGg
HUyZV3T6sWS8Z6djtMLONOAYfBlXlhCYGN/KrXy5G/2b2eT89HDmpYiBgBCH
RQaRPC/FonYeGdOvPuIup7ILZtvMF3Lk1dG3u3YbrM0tl2/K0G9MMJolxU+9
Ocjj6vvc0+00yOSjUh6AHIuK6a4wD2L1PGIG0WND98gmnMkWgMVbeDOl3P14
7IjdpW20EZHLRFR/Ayz8Ihmiwe4WwvfgzCTHO1zzJLtJ3CHFDKmfVFDD6+B/
DAYTHhXTREAjakDP0V/8YgQoipZ75o4xOLjkdMWL9NIITKApwhLHEuwDLUbG
K/fBBpCT0Cc4hZDx05zCgGRz6Zxtrjoj+uCXQZvOjkdVQ5ftBhOZ94f5jluO
ReyOr/AmeoIIxIEJGlvz/NeSBL2SsLCQ3XirO0Qlpt+x8KTOARB52hFG2xpM
B3bcK2S6OJ24WKS7DBNJPyyU+tDIhpAB8sJIGY7ZVPFUcPKXqQoSzoj1Nt9r
S8VxI99uvzmVsAshxFQTh3VBxkHQbKxWbLJ40W8S3tHm7qGy81UFOhTiH3DT
/VJq1sf3V/exbVIxGSSdzm13hjaO2+2YFxTuEbq89XD5Jep+Ze7KKnIZ2qmh
jPWHYLKtPjUI7kGIlymKKAGGslPy8fEUEuaDTHDuXZ3UnoXEY+kFZF2LklAb
IObViUQjbW+RRqLZ7bsp8/D1jGU87EeSp0Gwv4yNRrCdXe/nNyHPHhnGdREB
m3lh98aXaJ1CXQ0TPv8vC5FXkcqiQkTne0wewv5Py6upky+ksujU3P16FBin
hNFdpYx5m6ZfvemWcMsrbP2LP4dWQ/VT0IcFNeYIdn094qsLjDT0cYx69605
jh45y7FGRZzmGwgRqTAMopGnIwKzAg7qH2f0CHLmJgR54Llda5QT8/L3CQu3
YuaXghbFhjcYvEB0wUmYGskoVJB5HI4Lgbjiy9XrGiea4ue+Qdx5uHaGAsFi
QYvDZvcAc3DqZmPXtlMOx309L9AbQICJuj4RbZSuSADINevVCR4K2rCtiAER
ApuXDZU+T/eCzNcA5v0f0ctH8uqrCIWqMSpW4hxFwLj21sDHQBELZj3h62Ws
3fSZyUKVOi30H+2Jj410irUBM2UXIAwvTt5X6G/UCiVQdOdMQOzuqsS6qzYr
HhMrnYGDcp3n2fn3MotBFQ5+Q0L15O4u2zXpHh8kyPsQgcWMbzyMxUWLiOre
8QvIbqgkWnB517JVhFqQPRbKrzakYZFwrY4lK/rOM83i26v8ME0ZF1qs+sfs
RqdzoOxWmiS9IMJFHYbam8MexIGK/7BcZz5NUyeDOehBnrJ9JP9+vMWv5jC9
+VzjGDUjL4Za9k0X8xiCZsLW0UeeY/rXH0VcUWl5O9EYxDb/t4X2gn8Su46D
S12Ww9s1GlEM23Fx9KY0NJESLh7+LfrAL5j8O8RS1J+wRrwF9PWfnGMS4tS0
mR0ePVVM6i0A4f1/JUw3wN8WJ6tz9ZJ6+VkHOhfat6077KWzkYLLKgE2jvZa
ebFpHSBF5ROpDHs0La2o6dUW5Qkj1yegASZdhO5kpfb1w7qwBTzesQxN6u0+
0l8CAQcFImQ75fzupsWsFumGtEIVFdcsNPqh2mKZLRmZOsAEEsN5tC3z7nZF
vw66eKftbh4s/+gXbGLI5Q3sxYrTwe/mnwevHiQ0GNjxukPFi5PMpitTKYcW
ltLker6KgObWM1hpgfQlNxKSirhRJew+Pmd1e+hg6bwdC5QwK339zKslhmHW
cXjzRoQrr5sQ2lSLLZYBAJoc9m8AIyrVpbCzz4VSz4PMZN/sAGw1iaEb9a4L
3TK/JkGmI9eO3QFqa3RTZH/aTDic2Qi1hqdmU2yJ5YD0s7chzIgKOVZP5LbK
rz5zWzQy7YUUOAhnI1bQAnaVVf2rBlJEsl+ip9J/L5PrHma9cTEMEKytrfbj
R3uUciOW/ZRaFWwNASzsDjiZfRJ7Kh/Lp4NddiIWgIbxyy+DBxnPwnJzH6WT
byRbM90AJsIPNCETrShtCnKmWUKW1CaAz9yNJ8lHv+GcdLRDSVUenQipg983
GHuolw7+cYEYTtGJI1iqTVn/Q2kci5xfPv1u1z3X6ru0dxC95d5/neqaRL/i
yfbyRW9YPhMQLgNBnv+seNhy+NLz51XJD1D/83y4Dk4YXgoGesbLr8qk6CEw
NUgwvra77uQ1vAD2/vRlXUTKmvSeaNpAHh+NFK3PbyQrKDoJVxJS8pqiS3PM
GbhAQLXUMHiVMwQuhe+jjCEM+zKadBN5Itp+z5QXXKxn3eDFY56oRnZYMHuZ
HDNSJfg1Dhzv0ZnRTgQyHh2NGpkUB9SZon3eshD0h/tSa0GnMjb2VVkBf1fP
NG0dExrkbkzg2HI3zfMItV4UVXUS6AgaUfqT1X7TIrSA9YTF/E/P3a8CS21H
NkkraaGViyqWslAuykB0Y3dPea1oeTWqH7hHskE5i4hKR0JFDdMkruZ4idE+
u1T2M1iRkKA+/DiQVcL6ndi0pPHUGP2kY4UHAzSYnJnnXZ0I1w79srDWbx3k
Q8qlcu8wSs2AArEyMT44nBULhC8JLUbeQokRKIIA5KYDqe+8FyH6hjagcRJZ
m5ERFFurm1z3+UZBN/ZHFSfRUBh+SBNoVW1TZpYyQr7+THJmGnrwggAc7qT2
oY/H+CH5OEUo0m5IBCBMb22PSjqt1oMJeT62HOBbbWEnBadr8ZC574mqDbXx
qLh4ttCOThpZ+SPFv9bib2lawB7V4qCvEkGMVtLN1CgAXTcHttElVZaPJ7Au
W2Oo8BFTkMk4U9n1tCUyZJZqHLFKd77klvQyKrihKpv96Nv12dwIIAqvIdFE
2j0WEJqe0fgAdC1r3MvoVhhLKamgzW09dt9d9Vf/bmRDXzN4n9+F063aKXxL
EaS18I2tBNUtZcIwPnv2NC33rCtQWH10P24qjmpWODS5s6a3NukJ5a3YsFS8
LNBJn430BTf1fIecZz4Yi8FiPZXN16wz8lJyWQ5zDXNp3LkjIBfK2uIcv9eL
VfKKYgIAIIHnpCvOovecUKpv5prXZlV1Euk0Ip1ly//3TEbK0uGwU+8ks7Ia
FHj2grR5XN1kosrAi3+B5U5IABl5sjxwldUcN/nRzdBjXWP6sZzb9oDCjmf+
icBa+e7xUpGufbDXfEx7ZJiVnvXN4fM4dD6VXy6QUnDYxT42wwJNJnj4wvOu
GO0lBWh5LghS5T8DGVHimnXvMxQWhINZGvWkcs2WYxYeKLUtFFGnzW0mNssd
Bm7LMqU5z/NuGzsRKEjt5AzWuu50u5ZqEYNGTLDa4axNEwdBWHYKPq7rInl8
0rg2XpHqv0KToCjfJ7ACHRSGMzEAmOACJVagQoGCiXHnV6hGy/u3xt1LYdh5
vGNRQi6xAInWdrRMMf+MGzSwD2I9apY8jjup9Qeuv4Mjdf++Gk1tU0cspina
BR7/jeuo2uq5oAhxuCGIlhmXKjkri93xa2d6I64c4wUBNHP0Q+QoNdhupVoP
GWqYq8pnWSlHW8+boAGXeUVCAxe3Si4GG3xKoGA06ElNJAwsGAqBIbo+vHS0
X1ufR4zd458qx0XVks1tSuEy3o/qzqKUxYimMgt3GLvzMqIdbYqsH4zuAp1y
752Rc1bFPkhtr8p4kFx4iDGuXJlRRALqqAcFn3sE4bm5Qf/uA3wpcgblj8iT
ICqeFx0nWe1PLr3x3kKMJ7aJR5Bg5P9ujOmyFAG8knjKIwJgyUCZeVzF0U8a
0Ydf6FN6u3IhPu7bFO+hrC/aRJ/3jX5nRlEOne7sJgyeRapUI28317ODr32E
FCfbhRE5EYyHl52lVmdyBvtuhxRxB1UOzs6Ij6Ded/VA65jOvVbux2TXd5db
dQSWifkIEvLUO89ufph3B5wVEn51MPIvR6PMiIIS9Bj863uzcL8J7uFdGh7T
6+dmocoSUtOX94rSHyy7p/eO/deXRN6VgyXQ53vNiM3NSti9cbOcFcRQ51OF
0yhmk9CFZaATgBM/1lfDKuSMSYE8A4HWyGoFsF86k08uRZFnogzIt9s46fKd
R93xiPI+2lj1XkXhFJVVp6beLpYyui9frTfXDNP5HPskiObHs5TScLNbyX8Z
DmKgp+0EVQGH2NhPTtiMlwJMtpzR+h8nD7Sm4W4BPKRVAvX/kA/oVNXk8mld
jKWnfh5sWgw2YPbPnrKUcTV5sx435oMsU1phJXHrBMOEVRHQ3MBI2FiiVzFr
6/uIbHMW9XT5ezAoGkHUNADv8mso1Dm8M5M9wrZ0/ViKOAVEN4j8Tp3njAZa
QpylUuqloK+Z44bpJ0Qco3dAzLQSZNIEf6JOWfsPUZGD4jJppMTSFiEGw6lK
L3VogYi3LkAn2EsPLdoKWrESXkP3VRGVZLyVWKLfU4gtaGJ8IGOVjGFm8Qdo
UZOcwioVyE4HXi8sF/QX1xNtCg5xb11CF6M19foPJYq+Mc9Wyy6I8NLpN7ON
cr7eotz38yHkIkeoIMUB0CchR/m90PsVLE+LUePz1BwZQ2iZvxt8atOuPo8V
CJc21yxTXLhgdrj6H3Bq1oC3+DJ+mU4CyYu5lGn4Q5Q191vTKb46NqAEG+DT
mp/hjQ5SR7xeF6JEI3zznZ4YuvC1Gh6O1SwPTw2wc/IWc2bSvrH4d+8tGMn7
4l9oDC00+oLk86h814glFedTfetmcs77DsxsQQOoaYSl/9onqxsgWkNStsGo
r/k2hc/ERR+mFq1gkVSx50KfPkORUoRaZCnPap8RIJOvXbgTbThviR97qJRW
EquwoDgP/CdiBRVvyNwEx65howpH9nUrXnqUODVMYxJwQY6OUa8hYTdxRTHX
ZOxgSmP0wwgdZYan5+mvgFZSa0tEVyOA9Dhynr69zItrIHqKOaUXARtSiAdH
jWKZTQjEYWTYS0tp4Bx5PFqki1exOakYuGh8nnFi0PsWGcpVy1WK1570muW/
ZE2yjhWmvoqDbhgArLJ4TJRwO1eRci/cISmgZCfaHQb9KMFmoeJ0e5dVDcql
x4/2zw9eBdhvmoNW78u6rwE8tLR6mZKME6VGRRjlEx+HdZiEBRqJM+tPWuJA
ZOSRLkdyyfcY1ph0yda2QNox422fGDHBvljPYiC+hl8XKGnMwzrmTIZvelSo
pNEQb1ak2Vm4TyT7p+cCDz/7HNLvK0RgSwjHPonEz+AT6Yb9VAo091ZT7OzG
KD1NJsWwMOJoFwA5kXeke0/VaGlmUbxq00brd7QyAtuBxdp9t07Cz5I82D02
DE3jHbZ4hf3EaKricpdzDiV3fSXamzXLb0pisDK8Mru0jBuWXpXctukSsC4a
R98oxp/TOZ39K7H0ZdR8Ct+CsPfTWT1bVGbH++3LOysujBXd6B/BT4q+WnIV
YeRZH867sz3eVR2SwCVQdt9sm9MdU/qs1GeljHQ8myihy3Q1CZqaJcvyf1JN
gyGSpO/RyUcfqwAmCvnvffVbxSauA1PGRSji3i5L7pi/64HVRitPzKUGHeeh
DqgbzQfg8dijvHTPViFRCaiDnrS18zqBd1lp6iVArRr4CZyw3hcZsm/qszip
vHyNmTv51xFikeblGSgV5HlfpEEkBr7VjTxxJOruJOQKem9v5G4Oca3agkAx
HhsSs8A5x2NBBqk0DnzTGBIhn0dtRWUTI/awN6ePiQOht/gV8Guk8QhMUkpz
j1Dhn1uZEjTqjrV9rKAulspfaTUJ/64DiFFHciUF+2PxvLUvR1fWoEctcfzb
4Kvk2YeqiHlfpqD97Qab0t0TXsU+yQ2iP4M22LBgHcbfzUhTGEPD3vdFcfnA
0QV5XJ/1KXklJiKMOTboQviZFHB1NRpbNl7GQyFcYyiSnMQ2EdQHSasLt87N
1RoeHX7IjfimIKnrlwRmnB/TsnhiKWZyHMhhmTwwGnFhBAAvzs5HDwa92H+Y
ktKMshAqmvAXELVQ6Zb1YbEeSl2abAOfHt/1vOytZdMZo+Vw0TB+rK7DERN0
oysgYJRM2SajQgYRviSjAPvK/wcI8BPn+nRzR7yGlxGb3fgNwBLDskzRt7Pk
F7sbacdRKHzIIeI+j0G5ZRKppQaxprui1ysODtfmpj8FmX4zz0NH9jhq48uX
woSCR+7piRPEb8RJ21bNKA8Z/NM2UCUT81A2v3vRCnvAncMLLNPN/eyHIlQS
2fRmw/sQFNZ2422xOz6LiAogWpGF3B2e98wpxIp/wiZ9bhhRClAGyNDg2FYP
y2bKlgcJihuIGGXCiyCLnBrmcLKnm80BcvoAs0NFI3b3GzKm7FSgR9Ts2CnB
bXwNEsfslXPyw8NVXPl3UQLzhW2taMFOXmdD1Xkq/s0b2B47JAlOnC5bV+oe
T2+AoiO6+zmfnM2IA5KxTH2SMAixduSoerSPzskvF96j6c9qV+UGWkPtb7Ao
IP5HRvjxDt0KRSZZaxcBqAIHO3mZNuSV9x6aQ2/amsPMKDzc0AdNQMF38z2O
3Qp7FZuGAa8F22Hjy1+s/8/dGcy1Xo2eZ2oqPbOK41qeB/bIAReYPNUE+xHj
gU66cb8tbW5njHfQ0t2or7XYYqjqsqDLHfECcxLU6hsFFPdWxWSvhnXEru6m
2k/ObscBocq5ujiMVykwaptznyIyfiOJqJvkk+S0rnN/C4FRb0H6IoFC8AJm
ONXotWM2x/+RO+2oWryCBFsKTTfQBNtERlT2TIpJjOt8lkZuhymwZZjnmzja
VSmi9JnVOvcjiUKyNlJJn/Xm6svMDa9wGmvKIev4LzaaS8bWbdWSEuYLcWZC
F5qOxKlvM2R+3p82+eloOR3Os9AKQ/JkRL5Jqptl4PV4JW0H8mRVF5Gup2CM
pM4snBdC3Dw6abnbNDPgzrfNVKwkQf7I1q7uznG7TiOXpczJX4q03JH+BbAs
bHJM0LyxEtVFMGymWMFPTM3iISw63KY69ZOfHXTQKW+uDn8iuctj0RtxrZOQ
h7Nli0i5WMwM+yQvDXUh4g4VqiypeVONhOv5WmOP/UNpdGbpdkLmQ0KtKoZx
gp3HMUn4SJqCeFdJjZlct/lzkDDESxTiTT22HmMXxH0ElXRONiW5Xwwf+Cfb
wKXBG/hi+p8AOmFPfNxPhMnjOm3Qls4Ji9zc5pv8loJSWu5ndjMT7TuO2X8H
/SFpsz5emFpV9crOouvBPpYv9uhfgOzWN+cqnmocvA3huknENZ2uLpTXh+79
rRzeWvrITsOfUWnjLMPusE69PpeuKfftbHoufNzwyF2pDXc+N0h8rBJ+mqeS
r3CwThjC4xzbgilHhmsQtXGdB57NR0oXc0VLE/R7eM7KX4dpTtlmZ3TVJv82
pWYEMLMxJgK3rOeZ3P0pBH/CaObhRXFuFBLu3A+gush43v7qdrHYURImDls0
FbSaiAH9lbbZDs4CF07v5mPMbgWzSlwHrUxUt6hG4agCYjgwGcQV2a2vvXoS
rbKWeIuXJqSsyiB0C4frXevDmdJz1ue2yiyx+XTWerwHUtBleB7g1ipsdoNS
rVCEtoYcQXt4Ed96HqsKNjZ11XH6mzK8opux2WhqrAgNHBdF0DWQB9kM8Nz0
jDEqVPGU23Wjl/xsWfEQbZwJ4C5JiSu1KdGpBrGXRc187qXB8bk0rlTLaR5n
9je0xqiR2Q8eAi6ygS4s7a930pHD+9jYlBkEoiKq3hezTVraje4CGtR3tnjn
r6NkoM3tiDKMDTVzHCNOLIvUnyrtv3aQV+RlZtC0itV39rot/OqZHepFPCvd
FeW4R99+ODFSIYsZX3A5yNZe1IVy9o6wE0d+mgQQnSVYyy6n4XsXqwuFQAKF
8HJ7N8tRcyFO8v+7Y3FROKBujAFUJTxWQTA6rCdd79dkx++4mn/Hzw7c+2fA
BGbKynrKLVYlsBVjWGcXJlxR+QaSwJ+TmHN8L2PywQ6CwL4nixJKla9gdrBl
3hBuTcBY6S5ZLiRlDOOaSl3XtoLWC5/VSOK+fuP4ovtCalq+IY2V4TyHdmdw
Uu7D7bskAzAqww0dFiDzsSU414y1oKDQweNH/EFL4IXv00dYHHf1+k6i/if0
kvoM4B98HCTVjFZBPKaimaq5FuOI3bl8MpnDUnutyPh7AEXnoS37+QA80QjJ
QEUEhNiO442g9L9fWszPNUM4H9/AaLvzM55LLIfNvkwpO2AeQehwXJ9pb8ZA
/J3wmbzze/GHEl5oilpo2zG4CQucp3jgYAy+fFtO2ZvBECBtlAH+eZuuuOKg
pxQ8VmTE0SuUjTJ9zKeqN81ynsgnB/aE9UW5ysibENJv/EKX0aCGRgHkz3PJ
KSd50GYwHtOSm1aXXsaLLxL0as88WgrVy4whsgyiZVgxgLKC5q2wA+D2PqxS
ndoiTZWH5YDbJKA2pl+AFykCn8/YQHJ/jfpLHGktZPm9DNlfq1K//E896iLJ
4v37xnKdkCN9efn11Hx1rbJcqs2x0pYv2YI3/HW9YAOByauU6vZ0MoT3PyKY
YRgoVRf12J4qNlx3GS8yg1Fkla6weVpbhTmJnSIwxHb0DzJTBPE5e8c2SkfQ
Q8qtRV8Q6RgZ57E5AKe7U8xyeITNXC6ooOnT5IsO1hmcrb0TzesEqk2gNP+l
SAksnPn3TLjqNRVQo4DiqG+7zGTgUHDefy0VfCAJfZIFkzC1vebs72r4t0jH
p1H1m/n42AIAeN/JkPaXrrxX3bmx/1qI2XgBBqaUtea+KDoM06aNib9d0J4C
tJC4yuT6ty0PjXwfakKzE41D0XPMysC+4L4/Pj8olaoD6ZTVBh2xoBTZXVWi
ijg+kymG9608Tzodb73EikpwEHuYJjXGpXB89g51Xd5cSe5Uszc1/Kvutr9O
hIhBohKOJXjaic6ocIeyYc9hCZEk9IzgeVm4R3UXU1Ppqf5rdvLcKDxtfVTO
00zh9GLyJj5dtEH5bD8D9ZyOkr3du+lcOzH5ELuu0hqDRzcjLk5OvTexAieN
0PTZTtZED0L/zjmXKWLKwHWZfanB/Io0eQIiysRXcfRMM6rVXJKr4LJRctex
1UDfIr535jik60+0Jti51dfblVBKn6qTLfg/T8hY7PKXIsqzng97J87HfGEn
RsseqdgAdLVJFW7ZKVIMbKYYig/POPyVVkQJ/kqM4GmTiQriLeUbByG6cSkv
dGfKmgzGEFUC0k/por/lC0fHFVyQlzExa44bk3HDcVFw5aPjPhzxrsTkEDmY
ZxdnormUBWccEeWmXGoQsGehpoRHRoEuioYMXPsvTmOdMOACeCCIa19o/pyp
ARCIlV9SKtynykF1ng5fzOj1G430bkMTjjkMFE0glCk+tll8VHbLo5CJXNJV
wmjDXMcDkjQ7RWWmEUQu7mb91Xoyc6B2mnQxRdLkgEIa1uJCOgCvwgPVjduY
GHhPvCuJZp9dhR99dj7EH0U3RffuK8kMZoWvsWg7ZMY1QpxlUCSQWjtS7Iu5
0NWyJfBRQrT5uzU+qkkLj4KZZJph6BQ1mccobIaE1pGMTXrHoYk0/iug36d9
T46qIjdjiNfF6HBQSuLpv578/UhZKYOZndQTsuKJ50IfkkzrpRHoEAs/xpVG
ehaL4Ih5jc4YqRLE6bNFRL8BM8DEbhhuwhM/wet2eLyQ+Ul+40Kw3jZagy/Y
TWu6h7czG36NS/27ZZFJ7EUGG0FXuqySD5AbXlNYMU7XXbl1T7DD5ZLWJPc8
7Mcc+VIm5h0WaERPbq1aqieY7zFlFAm/xQHMhZ40QqpLdPmgUTQXOqRpR/Qc
ghtGd/xPCTkDDrDndW+wdi7QtRQYJLRKL+ScLUp2/fhyyIkW87G5qkyFOECt
Pj9wcY1uWYvo1u01ey5aPBWD4n1IN7UOiI5xqqZpQED6cCVd1V+RuVoAifG3
yNXlP8UfMnRV2Y2JRjfgMtFDjuBUbIBPi2Ars06mogynDs0exjaHEFLjcnCS
eDsq8GBwHS2pUZAG2qLOqq1855bYgg9jfnv0NsXrPiJpNZNrkCsn1sv13Xde
I39IkQCi9jWjYQYsSqZ+uBDWBoKHzWhZ76tHoHB63fSX8olf2oSkku6777RC
rP/kWssoPTw3uKAYR8O113HJk3HKdOtzhP4A13ffvf8xviRMq0vZA18+bs+C
tvY3xh1hZR7cAmuBpeqdSk3wNx4578V0oSxnBMh+DhIZ7pGQ2u6Q00Onxm19
PIra9ZzEEZXWdn12VMkkQoaKlHbxhODv7vIhlGblsDi9l0ppHmf4J5tmsCuI
bGJX8Bjvd37EWJ+e4Pvo0pC0ULeQz1J3cY4omM4Is9JpxnO7D2e/CdVg5ej2
f9KXWGd2rmk23YFDJ1P/SYYfBk3iYGt2jdkYEoosJy8I+qQ7EFz/xqPT2C0j
3E1+AytxrX88oa3Ew6xDm11gO77XgeBWdwazV6HaN8Md2z7ynV9Q/iUhIUEA
+KpXLGHvEu/ibDKiMyN8KpTRIoJWbaxZcVkIhxkRyxwcYDEcETmolC+u/IcO
5f5C+DQVYuUIYtVwADU6mkpar9D/ZIVUJXdP+gj1T5CJ85d6MXxFYEsayKQX
E31hY0IsHXkLRdO6j8jxqNnlMOVCcaCiTPuNvHQrWA0VSw+dgNIq+7hil++H
8gnq4zf1vGsizW2yyMB0ylhKaBxqwiucsCS9OY/nPebUsKdIY7UblC0MxsAU
CMrMmY9V8Ctxw1WsI4/zuXm1lDPC9mUSAoyId68G6a6Y4G0DrwdnIaRLftYQ
KRE6eyAu0MOo1mu5e7UQRnh4AmJw4ToaS2mayzoXrqusevT6pu/gANEjeNQl
JvHUC5WNE5Bsy601kfWzSKEAPQ06fyOqkOSfgcfUOf/kxiYUwK5gvK5THCsU
E+vi5E3JiSqa31M9hrrw0AvKJtyTP94vAhBFZ6mfgWPYbJ2oHV41P8CMgas/
gv9aXcqIG4KDxzCLJzrPLtZUAwKCHIMVKiaxZNNVr3yJa9soVjzfsIhDuepU
GusVRVLEGrxYyPETrb3QW51AM/h9VH+29Ks6Ky1rBj/ZQjVOEGJALWWDhZX5
VWgxjAsgkjvogm+KK9iSzl9tNCrKG+BmKzFBftWsvI6OPKRmEt4mlZzFO4c5
5Z+0qOyJgDQizvii2t6SrdWlD/hQpVnhGqeeetvuXrdrSEq7McfLjuiVcCra
APcFX4U65XG8vyAkRYUod4mH1efIjlSLQQFh2c5CJeXZKiF4uzS2sNfsvy7j
JZ/zO98rPF3cfvZXmKm41sgQDBGq+DWfJ6dEdtxp/I7bxmCvrYzSRyCtiFyk
L0wQKU4O70VJaZlSRpOEhRwNGelPKEhnYgrApyCEg8hIpntbMIQnHK2uXoLx
2P4pNuL9MsHwHc0iLopDmYuowPP8WaS4b1vuAGWagiIOPlVbfwIJpFx2qKYa
OzCPLUlG0V9FKHSLVF6V9FJteiSVVhnhqZd06CXK8DCpmPOeLlJkrxtRV3du
JDMKfX2Ts9dyBtd0guWUAGBkdI1VS0jkNHKg2bIxF9tr+i+4QTXWUZMopmty
ZsFC1E5Fx+ejWHkhrfmZ/OQxurAfEKZ+qOWoQKlx1Ao7HEbssQeg4l4TzzyI
iHRw+OUz+qyk752FiUvAfVHC6Wf/PdA6NcZdzSgqO7s7kGKTm0mYifPDXXeP
GVtpU+8LfQYHqJnmfRX/PHSkQ9qMliKIC/gLi+8PKagQL/6ID2RnzbyCD/hD
rGZGwDpMLy/L+W+f64IIzvmhj9tWgcaDEiOEao8vezFT3ylC0pj5I+73+Lw8
mXw0ZHdHipkv4mwy58sM8tDI8f5cljPGHKfWYuMXIdcGLGwMoYX+44ZVJm8V
nZ84Zx3h37EPsXdaqMxN+DGCkLEU3QZ57QGxYjslmt1msHI/0J/hvWa+HcAJ
66iwpNFGfQAWeWg/xK4m9Wdj9oOWBD6bGD/VZa0SQVfQzfE8Gp1CGXS9aGF8
LCnobLjO9PBRuXfSUGzDUxEdG+hdXF5ayjAAaUKozpMtMm+4FP3gg4bQRBWH
eXQ8Moa2lPx22reXSfrVAQt23Hw+3ckeSIwSn3j+wsDzW1fVLYa8MBrfBO9G
VMucZOV0Z4MkgheTu4SdUlCGhhR7QwWmTNCF0Nf7UVigaAlxnfTovq6gP0wI
ePLlakpXwrvjev5Q6bZeoQ/HeCBEYeJpPg2G2gdNq2sPQ6fuY/qvmK+Sxd3M
g7ZVGJYKWlqgLYo3aotriTrrpZsZ9pGKXe5jZDTyZz34EltzDHHc2lWqkBvs
UIy4lnJcPI47MT7Yr62mbfpy4Jb6gZm4ikkjxOmvBoFs//ULVtrBpZ1ILVVa
9yLqLzqqOvGbYAXiswqyODT4kdTLJ4u8MQObCKV9g3P3odHTbp3e5X6xvMdp
V+M85p1+Fzbd+pwuqdsI/eBrozNRIYtCeHKKrBvkNk7GzOZpuu+zJhkBWEjE
kYzMMYTk5asecEPAKYiNHc/SHz4f+r36INe5E1ZVKAL4JFs0cPJEDnNgfecV
F1KUHorFTaaEL9XR+tvnWxGvcuc5BU9rNS+lgRaAsSgG0wp6gXbKHpDcpUqd
aMyUQuG/b6Nmm+68MPW9+FQdV3nuWc7d6zvC/En6NhgTaJjKM6ffEs2vX706
gau+woZAaXOPaqiKUYBj+MBpdWoG8Y12DuXhFzeJ3X9zZbGlL37KDglJdXjK
SZxJuQFI10GelzSNDtsNs63sPD/hAd4fA495/1Q4SCgFoMUXosumigZJ8dGY
yzHQWxvVMNstaFTowm8a7keCiacqPP4Aib1bQU5Xu0+KAtdGgi+LvrG3OWLi
fh+HOCUOdQThKtvr8EnrILOe/OhPwkCQiGs/07A0sQWvWehIEPlCkO5KzEXR
/G8X4nm6v+86AxC6IGX1L4fAqq8abQ3TCO/OWLr2ELbTDVG9CuEMx0O9ePMj
17mJnRyHdWxmdKu5hFuFb38HM7Qbvfh5fPCnIq83pUzpvoOXmnjurdaJ+s2m
EI4E3kf7ZtNu9P2AdBGTe3zVEzeK/vjnfesRKEPbxxazLDckjcmzwZr20cG7
8vPJOrkd/JbgpsAL6vKtWIPIjxfTGcYNW0F+ZhXAS5CcZp6uRODHp7apn8dK
kQiRfk4S92h9ANGxODe/sRGGvzDZoOOTRgwd7CPaJ0zlqmv+5PQi17+NcC6H
AAzBbm5fxeIwXBUk/J5bOkY5qyTJDSq+hwWUihNPT0T679qS5ox1oYHU+AcQ
4tRjcGOZYSPq2MfBmCNAIydi/uw55fV/mRGPUlr7uYLa1b6gi3KTkO48Qsfp
BEF/SVdOxuWax69x1oeKz1Cj2PsK9cTXy2MpbT/iv9cbPjq2jQ7kpcseVQKQ
wHCRS2V8McMR+YCSquzA4VZgUFO1wB5EWyCrO/2BC+eQ3FKi2anFJt3kdPHo
jY23fZGDwGcpB/GoVHcw0Bh/SRZRJwmQQwIg855pauttoeFuAhf4JTtLYjEB
meuRr7XyKI+3y7/+ufNHvoUhilOynvNZQk9Vq62ngyH5rG3kV7PZqqc2qYjg
gzaPCi1wIjFJsQlg0A0z38eC/7pEvuZpooX1SUtZvAz1KZPvX20wEFW23j0B
YDWfBtjK5YiEa/P+pk8EsH07QgM0ILaLGQVTfr3BFW3HpP86N2E2VqnS9wg6
1tKxGQXzRfN0S6+EpCgq3t31pAyMGoSXI4QsISAJ+c+V6U6HInrBQuziILEd
iwity4DP1W2WjdlNYPlTt6IXcvw8iqWtMOASBWjVrPh6mOX5/gnwFv0YodHF
1ZpGbmooyBpsdcIROBZ4KPwYt1iOUUJ3OzM200DNMjlluKAh3HaA2R9QD148
x3yOH1/olqeILwGiULaBsKVzeuggayqVeIqaRqh/ZaCQycxP4Uu5KuX0mDow
Rs7mwrIFrMSpG3lVYKsxOSZuNpaoo1Q/jo4BMsf+9lAem/PogeVN6/RcZDsQ
/JCWtp9kdgDq3EXaoo1UeGsZPR3mlp+xggN9sAQyc4jIyZVp9r3QfAihRQnH
Chp147aGTkmCzRSB7DXmOagPYV2p+Sny7a0Vvs4tM5/h9Hx7BQC93TinAeun
Ss53iEeI8BE3dJA1L57w3jItmZqOTKzVrEaHG/In19Nn+X2ZaK+PvAGX4CBJ
T0ScFqflFrZs67QHrRiGsyzQJcvoRTwTlY1yzYCxFottbjlO4YA6LvLrd5Ep
PVIBHbjy+IVICZyrrGjTPfH7rWmAhqDWPYSWoErNZyNJqHPFSh2A+aJ8wW7r
a2ORqh5HD00y/yOygtrRT9YERlInXYG5SZSewh9zh/LE151qOSyePSpe5hoE
qMiIgMclBfZZOw2JdZNmwxQqpTUQ2iVRGti4hffvUS9RhJlm3rf6IipLMyBg
W5phrvGi1Golbuk0+Myd+yN3r5/eNiBc/TTXednlf3Czbm2eqbWpQfjsA4A5
bcHKhLlk0JDg/WbouBni8lF0SphBHiuC9E+jH4BN8X1wWhw+GQGIZo2/WqtQ
zgrvra1FWa3SRmxHoRwg7PxLOciuWnvlZ+vZkxbzya4/MIekxH2KYEPqTsRa
YWVGqBlGxvwImO8BUAu7jB1qYj0zfV7Ftm8SiapyESgtegY6o9waKOT59M/c
pM3TW4/TasalLarJVwMg6DL5Mpun4aIkhnUm1XR2sq7dPHzd47AcgqxdqDgu
JvS5sX/hKuxivA6tDrdpe51IuyNQWiv1NHM2dHvi821gy4NEikE0kWh6lHrL
q3EvsthYZrynLqktQoiJCHVGGDKEZdbrBh21sWSW7bcLK/QeskRGFPzz4yWN
qaAo6/sGc6h+eRXfTAk0uDomJZmeuJ1dtI/zFvbQtiU55t7RznslHT5abIpK
8MGoN+qMX2OgX59eMXPb38Lf12Mbbgfvj7MZGLfsNaI0svq63LOiEByPTNJt
+dt/2H/tktKDmTSmLDsqKcLzFCgIHdxpUeAVd/tqxX5vOo8MxqaJP/2YzOXC
B83PHUGZAacR4AtHEln1hDeqVC8hpRxcqF+1633+39B1Gv1GpKsnP68kntkY
PabtNKoXktCvZLycJF3djwkoSPs/IxDLXXKe31MYigWjzkZc44MlgpQY+Dtd
ApvRHXqpNpnmy38yec5ZSUErJiNude2O/GxS1IjA/CWiSQFAu4GZacuQxKpk
a9Lw79klaHLkCretHN5u3AdzEO4iXv47PkyTFB8MkctNbHJPUuUKqD4zZZef
k25x6jixlybWl+1KfD4hcuPmPHZqg2GUtqm8yyDyZxBXfe8abf/XvayWfJL5
5XBXW1vNuPpBCNUXDcqeQbVaGk4yGohZVHel7eSoMLKDoUexCvGgXEQtT+5Z
xXub622Rbwe9pGsmRPPQ2xMz7ulGDQW8KN9iSKyDNMucFiBU5T0QLD90vZyN
JRvPoezAyjxPvjCHYWbBraUoMCVlbkGEZtXoEelO0UH6e4KtrGpgts99VrQ3
Wj6RstCTL40qNyHuXcPvGBE2jj5aq9N7/4bGu9WO3ixuBhr6+aw9U+fExixC
u/bbwVi4DTYNU6Ky/Kqgx2sOX/z/55GiLvlF2Q/3Phu6x2Wm8aQIylhC2Es4
QFErYZddyylxIAp6SJhq8emjAQsiAHJUz0dOxhjeuH7M2DFTUN6+7Wcs5agJ
fLdlAHsFWBp28NI97Yh5DUFAD8q1Hc00p2LXwBhzjSB+Mx/q0cd+WLeelcFV
AyrpcNeHWadJQzpp8Kl+uYhyO3kX3hn4m4tjHpLvEvIU/TE02RAERxpJw4OH
D0matrCC6ogFBXmFdr6J0KeQUu9NNDaT1JB7VOD+kNTs3Hw2jqKd1pOKiWXy
tCmJWwAYF/Xhyjq4loP8+gWbyLwqkcqHyvYf247Nf+armF5dj1M7F14E+v30
DlZ4+HAYxDNmBY3idQe4R4K7cPC+LDs3KkCw15EtoLFgkPWZllib7CViS5zg
o2Qiora1b+s+rWJyl4PeQvrqv1zReQrZMnbQyoNym4g0bjzvoxVyicW58a0Y
g15H1ouf4nO3GGCwJbuL+V6nVSsScKMclTuf3qps26ZK75MK5tsypaVtoTCh
oWPaFymGwldF+6GXRnxlvG/x7JmqTZ9+TcWpIECw3rhkKk/0/gP/atuLTbrh
uJGmsMOw+S7LAKuJfT05eoWL9XM7v5+kVjMMtaLRSCrUXEqT3A3qakDQyz0n
ZIpr7kb8+7JS843sQD5MPyVeEDTvkdgpFLF2Eg0e94abVG0WAwxyWlY836FP
STiBFYGmb9zwBnAr2EOjbPNPhPV6AL+r6ufggwef71mT5nVIOM16Xqt9wHcr
O7c1gcQLO/0vIEOfJF0bszezLBqKi+eLoi/s137sFoxOFumk6Yfmr/w+SUea
lb15VZn1gDCTGXralj09k6Zq1Szss3crbfQzU3jXjHnrvguGP4BVlXC9vMiD
qjbcm+G6bMvLcck9b+e11tmdUlc5AYJIWruSsGRkfqRw1EbCRpb0m2+Yhi9a
QsiRsqufSdY6YpN9eAePNfRBglJf1htPCNaUXKD0JK39tEoUZrrcS3Jyl2jz
mjj5syPviXntZnCGQ+hmajwKHeKW9omzET73XqAQF8ie0iVX3+jD7q4nuWAq
pH9ceT54RmTJXw2O2JIarkkxwZnb7CDYvYPaURtse543ybtaEYCBRcltMyGQ
bNuZGTktVqIXXLPAgO2Am8Ezkn0IBvzxrBGMhnV67FqVsg2ygdPQ43BUfOUv
uIDG8GX7UxaSmjsbtIVQgqGw8FQcOoorczxUDnv6v9hYXFj9sKGZl2vF61Jv
vJaMZBCUe8sgAfrdmjGsPBLBk/nJxNi9kqEH4dt3Px+zCCvE/WjEp1FpZO3t
t1NyEh26dgEvziTN1TY93vLLPhWSuvawsKT6vL/31xtfRqhkE9Q0GuGM0utG
Pd7+U10I6kmUNs+p9PLRZ8zao14URnKgP6irNDqZLn1Raeg7D/lYiEHJfp2l
fsozU2qMIlvWDOm2hneQltmF6ZQ7/TUqFHDvOL5W2ycn5UqVUeVBiRW/WOOq
A2UC4/ZytQhaTGC9tPCF5vy4J7qlKR9E8qYS3O6bupeQp7DyDChznahuX7ri
IrUBrFXnnH+BFZXSVb2pf+1s8fembe43H44oi53bcVbnAbh1pJ+OfVphWQrB
Euxu52HYelHutR32aL9Vbvoq3d8gGkjkI7LRQnkMvGDDB5BpCCxadTwrze7L
6rpah8dUOnn58Ierj8ZR14ntcnZb9ERrtoWUXpAZqJFBxMd35WQcQWOfimL4
3YhXqMImq9z5UMgRqNAE9JS3sFQeLHmzRciM2vYFMAqfRLoeKuupdwOyuJeb
QcqB4N1abQkRZd3DgNxwcWTzwsyhSTv0EC5lbTPnVcJlGhDoyq9BTdy5KHQ8
ptgag4IXK2+bazXJH7i7Xaw/gsCE7ndIEYIZToz2xgtH7Zak1mJyGHTruVNL
qKY0zR/xG9nWDrACMDQaJYZmVJVdQa5SFTTHEi1OGCYRJXxqJ9lZYuxOFkQr
DorQervMvVNkQYKgR8anHPqJHFBacW2aB384Qc9i1f8Ou0NdK4AqoVAW9ZOx
7X0pj4fWQbpM3/uG8eU44lrgicRte+Ym6UbLeBt/ifnkXxZhWdnB64CM7R1x
RXYTU6ZfQyYY2bkXSZymJK+bhxrVRaX8PGOIRXL89bGf1Yz8DS13AFeKkTvF
FthCiELYoAWPDHwDte3xaqjIQIgOy5oSvuzxb9EmZVJXfsEQ9pOkTN4M24PK
ql+w1vl6r8FTofe5IRCiH593wnd285Vj+9ed5jvE3WpF727uRm9dPE5xbDZO
NuXJxAJ1D6xxQciZePgdfhU3oP3LGgFnYRgwnZYLqREZBsfm8r4nu1ObVjtR
eNaepzG7kCyt77rfx0frqR8+XgojJDlwY5IHqJwgMY0lDy1PQxEq8XdgVBFg
6HK2Klg0VARa+34YBsWhDVY4SQIpUq2SydfDcOPUsEtXVehS0VUDX4cxAg2g
3m6gjDJam2jiV1sPre2TQcCeEBolwh5YaSst46YMyL18LdpVBZlzjJn4CYGr
tLCv305bLV5/JzJCTyrYDB/TzIloO7WnkcnsdxuDt2sFrehvsG7ZCPVQ8VVq
tvkM4uAHvTtoj0dUOxg++WUeLzjaaiQOd3KiSW/WC+kTP9xDXSOu1x1lQx22
tnCgYije0ymFQqiNbigD/WbvrQbVDuu23dmV2g13jUj9cXUUyMxD6qjPRK8r
gqNVJtDkqH+W6Uic2adCyYCFHZueO0R/KGuJpLWOtyNNY+dvS9N4TuUOlHet
mukVkQAV+P4XtgGTjL8JysDAsMIr2fBfZDDlheAIIMSioHsjRN0ZxkskXXNI
50PY9L9o4xF1c3bc6WRDzDuFKz9P+TBV4OZ82gckhGk+lB1n+EXxpUpG/AjI
lc8H9audcUSOXAvlgAfaFt6Em253bbwNOcVaseFbhc0lZED3tMy6IFB7fJLN
zfr4vul5qcdJxanXY3QZRrImLYpqDw1vTcNgWjmkmQ8i9H7S+aMzdqOW38hB
c6hg6C4gw4c9UD2KYEdE3TlFytQdPJTwvzYIbJczJnC85IBFbt16ccnu2a79
RlRBRP2I3X24qBm49+/ZBdXp9/VWMUS5CNRvOOOU7jduHx3sqnq3zcWLZIJH
4M51SRdJlRx7Ilz7Aj4DiSknAIMjdVeTbSBagbM4ZtMYYbYspXI/WOt6Uq+d
dnoe0REV22MgK94nhOmq/GwqcoEmkzHawOl/o+eeerroaBU7O/ZD4kWt2tj1
l8HYnnGlZs0H2bNsFEE0fTFn6o7qrpEzFi0C4B8YsFWTSeVcdNCHpbTRMynQ
uwf2kPYpwvMp0r1F4E8aPMY5zpJ+G6sLZY5K7+FVdeu+XSkhN4Fs4GNalUIl
YvBoOii4dKlSUb+gxA+prLLfmADF/OHg67cXA7clNTUKDOneuHinRkdpMmoV
fi3Gles7sUWS66hE9oqmYhoW0NghJTgQ/mw7Pl1DaKMH0nvqWeyr78qAlmtS
ClJnPkCOYcjieLIioWqWgjID6u85ocI78G3ti4s2AYCz/UAhcrGsx/FvG487
/PQxCrzL8cHitqGjKknT50NqRDUgTfUDemEKaB+F0yPHbYIItmzG7yX1nCf9
/yU93c4u3b0Q3GB34vyS0hprC2cuUnosly2udQZsMrFVhz7fkzcwaiaVJrzN
GYDBzIcVDBY/uNi/aYURBGluSNKb2EIt+CByVNtB+E9w6SqYIbHC0e1XHUBp
tXHx81fuIsBTGUPlaGHgVgXX0gq8ozxZRwEf8QPUmTAwjtZu2Lx/I6C3tNP/
5QjF8X20iFBNRObS1hy1MAyToK9T+BiXDnvDKdKN7PG1eRfjNvwDkJKqTcsF
dMLOPNhwNFYuFRx3pYGuMg6bNxQhFtU284i20KtO1bxfZm20wuqG/D5eMj8K
2IHqQ+ATRCMLuiqzgrZ9lsUQhwpscLdipJGde9GHht/ASzifuHs1Fuc0j+xQ
YtQb0X9bKse3P3lu0hShlEeVJEo3eGyTHW85vX0C7/9KfYC855G7OiCyTZLm
Bs2nPwzj4GI8cecvqsj1RAo+AKlFzxKnUPXE/iIex2TTlgPDiHo7gN/KkeNX
vTmi7/hNIYgNqQ5e7YsI/uYQLyVE/3Nrp+CzZi851+3mfx4AJNC68UbWNYlg
fY2R8MjwWyoRxxA15r+OyIooDqG3/YoNtfQq9BaPw2H3z6McxH5pMsOgat2w
PXhcQlanRoAkacO23YXyZyXCmZiMfisZ3syuzhJsT3B2GNRMPbjClYeZc17N
5dj5JvWxW8Tf2H6LBGDZ3JH0ZYaGyM7s0dZLewmFuqQg34zm2U7FqzMuCg+7
eaQLhf+vFM8JAMqKbKfxEQA0pn3b3YgC7JXgxr7+Kc7ADy7oQfogwNyksCd2
cOMez4PhKe8RGgHdw0lF0TyQKllju9eRwKJ3pFD9PE0CbK0aeurpwXhU1LuW
Tvsi3hZtl5kCRXIk4HsQicgDLnGtIT+Ffeaz6+IZYhro4joyelk2YcPgWtUS
kl5ZUgzkZp8Q9yOThiWR7DkolFp+UiMArC4CGIkRivu4JQ6oL5oMs9gwzO3Z
Em4BpNcaj2pCygS0lwWQuFTtQcy9WSMs2v0cqm9+Bj2/A/TmpIHUKN9OcFw/
LTHVqMPxV5ZLErmQVkyGDMqETGpiY1TCHKrID5Y6vD/uYZ94j9ejXQtiWri4
jpQHnXJIK0va2yyCmQPSHC6Y2mvL7RSSLAJabbvh3qNdhECOlM4rpoe9Utd4
H7GxfvkPAwhLZ38FzJgq/Y/fQIOPpXiL9JXDSuomLuzA52iDLMVCPTNXMwk1
ewqIcHh+xvui23OO73OjAyZ+hK/+NaFN7EVPxjZfwmEkxl0YgL2JImD8zEgE
mD7MZlgfg3Y/MINce5DNNTpR+SkL9sMjRjj4picZTxpRTy2WeuVl+WSzfopd
ehs+20YUr5SyS8HFbsKCFPj95Rb51iG7LVMK3x6OqXHlipQWbfbxUo51tqZR
GeiIcmfwUnSjwLmEvqeKQ75ecgNtNac4gDTXVqJVd5KFZvvWg/6yDKdwbOA+
ZvH+Znaxy7RFHvWhuQG07rxYHlMDG3ngrSP1xPyczl/vnvWBHcYXdtLYblBV
4wdvCuUcNW9c218+rkTfMmF6mZRuS46PlrXQFtC1ozfTiGoPHS7/6DkzXnG5
1nBa+8+bCchH6GXvELle4TM+4QFbFkK6CkGpI8VVVLQpn5Aj8YFO5ZABa0Ww
F2FZH/u4yb8z2QdCCLsX7Bt7Vdk2djyuBMTkK0BnUPj/CcXdnNN1X7yY2ook
V9ttXLA/EvtFLC61jIvOfIEjiKTfNyFVheWdB1aMTWiiXB2aCSlb8G7uWJBH
jNLNojdBW1F9QbnAf0FF9o+J4sn7XIizXQ/e6uUGacGaK4fMU8QrHMFFltLB
2u5HAiA/wQEtYB9nCb+2IcI62No37CdKaLapuUQbu9sg618jhzXk+YcbPoTs
ydVifwz+hOIfAicEEPm3OfFwnLppZkfYCuZBnXVEJIVYlf5qB+bhD2Skvk1k
3+GbI2bfPo1JSO8Gi3vbdUnjW9qbxQ+vjGSuh6aR/1NpxzZKOyi7BxVx3Kuj
PuQv9+kabDQLM4d8Hc+ZKPAMSBhEryihS72TZyOeWxiajNi+G1iAX7KZK2dI
Fxp/mQj/9G6hf/dMMMj76lxZBIghH7eBWP+jw9r5N6VrsLJxY1AnQEdlHeQd
Gu47f9uoUnFWrRym9F3fqZKdo+scjLVQ8V0iG4Y1G7wal1TgrTVT2bISfr2G
jIePLR9uoJQN3eztaWvnW2Zjx5AnPcBNdQmj0Thc2i6nkgweEwJDlSDd6A/h
hOP9kk2OYjkwsqfKa5VitjaPQL39xWeLp0RRcdq3mY7hxsMYlKdAumIYNrKf
wUol+tkNDuUqmQ/dMl8/aFkKVS1jVOo5fDJTjpy8mAbkNdsqIeK/sMjZ4Mvl
j3J2poWD5xKnJhsclGtoKeYtOSa3DK7P3wy0GkRBOADbZtoXj1Lw/evIXPrt
6hU2GAnWQUXpFE3Kifd9m3ZgfXAXUcCLdoXHAWq6htir8budanHKKE+f8wXH
0+XA6mgJ9aFf1FYE4TV9HUyReTg0It20TsZmCSyi/Z73rlyuqLmLsp0+ejnq
VwM5h6jLq7EU+yXc4t/UcbjWNeuOYQB+QrZ9sxBv0OLMvijhmEcEns4AY4hQ
SPtuxaD8eRbyFAm4bY8DAQz275WS2QkOHsn+WjKHNZlFFQfaIwuNbyRDCrtW
Sw8BjSwqRsIgPua1EU3MH6qh5NGTiyAmpOyQXOAlJF8DNsJ31XA9Jp/N8IC0
a0S9plrAiQD7NZODYmifLi5mL0ubm92fLdXKA1pXJ2J1KZfdBqFISngryQqg
qKN3fH/BuR1wtzoDLfFE//pAdxmW/fXi1XPBI5dieWmVWHte7vG3IADRGs32
X1Td7q5e3ecRviTGHeQCU+hmBgyTbNUEznNA9rS7VHThRC+grXb3RDbSJRRa
xlIrQOwooWdhK7HZqY5RUoYOIr/oX33CBLgi2NQqYzGo7URC+aBXU0DC5zLr
xETn89xTdKMS5H9PU9W73S6eNATA5hEK8SDDN5cwV5F43qHf/VbBa09gznfI
URjHVPoZduVncsqLMPyPHItTRl5Benm6RHuxAAsOMhPq4r9z0MqKibVPES9E
4RyweLEYulu9gc/2mjVRp/Bn5G9DApAfhfdq/LLaHzqNxyDq7xm0VzP69F31
B+4ESMFzZ5b49JsdjWrlZfnsjQx4V/5/rs7I7K4BDCxeAi9hK+9mMRum3pf2
k8NcEPPdUyIlWvP8zM80OeCcflYYzOi0Dq4jaYQp5+PXL4Pjxyg/I2kgo1Nu
OgJlhwNd7HaYmTvSFVPeXnhyHrh8eKVyshsxYfYobHNEGnTwAHApYBY+ou3t
idZkDeNcbQtiUWObwH8lShSj8Dn8Q5Owmo1qJTUqnvJjipIgs1gZg23WJYU3
FCeqjRqDiXEr30HevpFVZNz7ZOr9e/W3jYAqNqomIVfGSzJFHyFeVOMnBM6R
QC67c2txe+BJ3XGrVHSWYrjyin/HgVuaZSTnPhtqAbH09N3DwJMNzOf8MBKq
MqWk7JbRx3zecpHCv0QcxsXtVSEkqrHmDpMB3K3hhdRyWKD9NrmlgtD+18kT
I2foQs8PCsOWotv525pQ5eUAKOnB+FqALxL970k2lzpU0JD+6pPcGmCosvJu
p9uEAE4aw58haHJ5adJYjg3W3occ9KvG8A677YSYAWXGh9avpF/WhedpIHqd
+VYOslwqdGlPjjkYX2oZCN8jKNO+TinupBA2ZH8hViJ4IyZVxPP2YVxjx+aQ
pNTDmqOufzaLsG7D7omfy81/CfQs71rG9Nj5uZtZRwrsIUgMX7wddzABACRE
SdG2PqgDVN5EAVzFJaPvYKWKfyGUBqtr1+3DCYU/XNSqWdNes4vUGXlZ+4o1
NEXPgSGOAePy5sZipLEtp8PiMZYg3tDc3J4xNCzIc+RixN5c/00f+SpfkNe1
k7qNMvkpdf/D9BEt+3/iD7goK5TCo9lvqCYkHW18toZeDgtmFpwyR/TqwrRE
He61m9eHqm9Rv2ayhsMzxBL3Yf91EXU/jrov7+impYOjAoTTUVBI0zFogI8R
e/dbkd6pio5hus2h21Sw+a0M/esl/D3DU7qlqkcN+YH74L+n6ti+OPd+P834
52y7AY/fE4cOWbK+xSqbMuDJUu2PYAgD6Qdz9DKfaoBo34kxcvYYD82VabAc
TBf3krDBB6wYLC2ESveECnBCOGyKXHTj7njxkbQoDFSNlWRz1RRmx7ozhomT
ezTkhJw/VjL3KnZJc4bl2jUMmolltjIuGmwmcfdGXo0+N9eNauCXxcEBME+e
WlHw3cQmo0Ru1b2qakwOv5Uqx+Oout7xoBcdfPTNWdeA20fA6eeqf0Ej9v91
g6N3s4tOceCfLwzc8rTHluOk+hGpI3yn/CSOnhnMK6OJHE7xTt7wgxFGvzBR
+2TiOUmOPrNq9LQ73GyPuj3TFlDiHhfDTi1J4Ai8pOTp3EHyaZPbtidmWVqT
GMClFqQmSVI+XjPSZA46EoUFFvkH/A55kWM2LKsflWgEmzCpmjyuMYQkmPLE
X/4XWOS+k3Nmg/+qx0c6RTWZQE3pK8CltTpArm305PECMhfVt0JLD7aR7yJ6
snuhYPvnXSHwFfDZqJYEjqQLFx9Yzs26h8ixWSb7g1wYyT4SwTtk01bmbEbY
CqaFKUzmrmCtmk8n71iNSP987xSGj/jHAwnBNV84Vxiob9KcCXat7qrCsTh/
rksJG9h2zz/ppVqF3w/Y7gjOZDyKnMFv2PH68WKiayJ4/DPF+Y0FdciCX4VZ
scXDDkktLZuNcUCQNVB3KU4IU3BcTBoTz2kYCOlR6414/z57rdCLd9cpXnZw
pMaQ2dk1SSbZRS5HqZn+cuI6nAtUU38v/kQoRfsjFoQjy5ymHigU/RYvu8ss
LU9KIKAxVSt8c4CEmNNHvoBIYMx9sTX98aXqk7F7vhm6a/eApkfc5xGOawfP
LeqvPEXs+g7eGQTWbE/yTGV5nivtJ7DCnkMyZn6Zr6XsiGKGLkoKRPEwUOtD
uOYPJbPXRuWy89HirDJFs6bZS4kyEU/Nu9YZ2C6BR0RocQjxTQrdUijileUW
N0G1io83OT1DiJ86qsU+CuEa0q3AxAWUtYFwrrhR9v5D4/fP26jtc74PHOc1
24XB5AoH3Bn8t5BCMpGHUCFMo7ZpSswhpwC2GL9M7pfFJowHNOjSbJWYCcTS
LwW8p+HkMHYo/ikpZqzw9q4Rn2DyNDti7UaNspvu0X2lIuiYrfZPWDb/HKmW
gT3K9qpno8h6LE8VBGGVlWc334hAU4gG996LQAWOGKQ48P43J7vEG7Bi5Ob6
pku8xqkBlyB1Rh8IN1BN+igPK1pjypvkA+E7juxm3i/miFzjpcQ+tu5jODmx
wdvoL73rW34lEVwExLasSGxxFq12dJRtrNstTJgUwoPAzG7FpEnJq9wTKnla
p/HUDGmHYsgGQv0k4AfTvylO+1VvTvJA89aA9HiH0oHOngFgnqqhvXCFNBkK
W8lFP50BQuw0g1valx9ZfyYM+BwBVZ+PgE1kEFbMS/Tc2K2XvkTlaLae+n/w
Hi1+XrXaMxFk6CvFaE6XyljNZaYH+2FdEn/xT6gUNyoW0IdJ0PvFfDCtgMTj
erUh602iexWIT92riVBzACkLosZSrVZr5tpDJpynv5DgcMOS4YlXG1we9V0l
eaQIRB1dgBs6FHZQUMxMDvfnhBubnf2oNnXXYdVSSB6ckgLd54PMNi/nLDnW
ZqRffbUUUXfDLoX/9/OvGX3W3X1Ajt/R5zYgzTGx/xt2B/Cb3TdKkW2+rol2
Pd6/HeYhMACSpG8dsdVWmUgdQc8IsV0vp0GSmUt0kqNlQrxhrvgOXVdhCMs8
VfFzvo8u9Qt+WYK8Vp1njxa72pZZOWC2RHqN20q2pMN89dsggdR2KNp1kc/m
fKhI35jbmehBGBHDS5fNLs0mM0KwsT0E/PoT4uR5oq1dBdKDHK7yW8H3c1SD
yhUV3p3o0TFAvjajhMdpOljqYF5GOBT5hScK84gPmASw5D3TxXvmJ5HUdwyp
1CY4L4x9UQZuVPyx5G25CSwWGxeXAMfHbL/BJTG5K5goL2o7Ft5aFWcNDnbu
nNceMHdOgJ9Vismbw4Ikba4GQd57DvirtPCooPfeqIJS///IShlucrxfk7A9
R8R/VN9yNSqrKJGXNBNzy0LanOLUsa1d1rwrwiJwIbBqzVhC/Z0CkCg63eKu
fq9vzgfP2hsDWiIW8A1oYyxCK4qh5ypK34tYn6rky0/cDSyEc2z0kPT+mfQu
lZTrYyg+DCpviDWMqrJdK2AD5Opzudj9mwfgp1teqW/BsOCl6IDOZz+FLcCQ
f5rK64CQQhq8LB8przgEW9LzBUu6/d5rnVjFoaf19nKDw0MzrjNDbPZtZ5Pw
8QsbrAQTvoczZJCREPPqyrmFegeYzwY+O8OMSHfI78HBJcr8g8h6/4WWMgHR
jITc7ArqvJ1Xv+qXVXcCJqNCTfR6q1ZdBX7r6Gf9KxYKuvsnZVEA95Ffa6yZ
EZQUgeGqf97bSZ0nJRJGikl6npF1/wmX+/C/iUxdPTVfgYGUhsOXbPKr7D2Y
9TRkNGZN1dxMe9u2Tv02NrtsiPveXepQiaHawox6466b1GQvMD/upiwRdNgY
Y4rHfgsahF2DmMeNWQHR/3/cf+mKxotX1uxKdaeRfLY7+mUGdwowIiLM3+bK
9OJ/N3/LmRo3j4lVj8RGkx6zQYKr+s3AynmR+tPG820eCzsXmYTKtZRjfn/K
1ck9fbybnyc+aKwe+AhF4KHbpPCh9W3guIzsT7VfLa1QTrm7poHXI1iwBpMi
E52hXB236H5McL/0S8X7ey15krhGP0JT3WZEP66kkpzh6XA4XbkxGSGBe5zb
EzuSz6XobDmdynY6a1Krgx0v3IHklqnOIdjZj5KYFo6fT8TLKOyu13Tz8TWm
4DnnIvHpFtdIgXZ40a4KCpayMvZz51HQmXFdVCZkwlvw3oithSLyEjuJrbYA
+6ON6T67c3eCEtQiFosiKNnvGqMkjFO4KICF7KmZCGHgkYZSqsD1Vrqxim6F
zVnJUpULlMBrUSf0Pv61CgkILmB0ToAqry4Ts7W/CdyKXkikoiu9Ea6aSMZf
LX9z7/W4Jwk87dQElON/rji27f+dpilcioFnZt8nq9HuTEB5VUPwrZ1m57oG
b/tQNwnKJcN+QVExcJD8YZvMP3V/V0RzZ/ffKJu/zrqb75I9LkjT6XNqkdYi
o3HZGCOk+ePrStkNh8B0g9ZjqSorXakhslkYLiC+QQwyCuU0HUM2tBkPavvf
YbcV+s3AENfi978FUrLooWjY4T6EKcXltNwfIr7K/Adf9tAcWh4cmlbJHy64
sJ1OSGFZY9jEpvq5LCp8oexH/0ErSKEt4sgH0pKdU4IQymSxqoF7T8DoAOJF
vnfeXZH70IYMAZFu9fbCr2/Mg4K1HIaBKz1PZAp6zYT1sPSiOFiyK0LD74qb
TPYUxaomMO1Zr2xyFn9zEsNwsFM7Y5eTk30LEKX5y6efQADOtaJUC+MN5llH
pb4TkV26Lukn8fTMVzWG+9i+33c9Q7fFLs0uEd5LKCJpaKCm2bfhbduT0P3i
cQH+y8hvG5uIjtfDHR/UWf8Kqe3CpD9UPU0A0gS10I+v3C+4098W0W2j0q6k
Lct5KaAtY3gerodORMUFHpkeq+LBx5pJRyNEqczb+MAd+nUOan/FcdseRWJE
lG73h6AJ48yIZb+pvUP2vusMHVP3FI2GsXTNa9AQmfSUcjZpFPFhZv2lnNXE
P42dQkxwBWUzHHMLaqdEsEzUC34e8o2XzxdRmLjYpUdCyKhhv/ooLpfxKo0c
Pcv+Ce0jhrR0IfNe/vs3LLLEn/83UpXqnosRCV2mxhzqKzKSkrekNUWzkWuc
Yy4Sx1eGBIncOrXJr6QgRxLEqSPpIk3917ATiBLsP9fk/zvanOusuyKtCvDh
OIH7kI91ryEVoz0q9iKd1+cxc6t9PCWVI/8q/yqIiADDtvO87MjmIEHYKuDy
LzKh6a9G7xZU7fB2d2vPCvRNt0i8DFO/tdP0PPI0v3Zw557Vi3O2OWdvZiYI
9nbkKeF/j2yt3yMbcJW57JIc7aP/ig0hp6//gBMFa/nEmR9KxJLHyyJeBXmB
IO+05HzjJuQjcZvYE+1A3zeWonvU89ZR3WwBOJVIwH0cP05sV64fcHKwEWOW
CiuDl6if/osQwUE4mOab1do1O/2MZ+sQw5LvGcvRt7DgRTjWWhKM17Iog2Dk
N2tSDO++zstGP6SmiI3vY7omoikEQ66fSdgFLJJKxLiaE781EzHmgH1/LoFP
mdx6cFLTR2SaDersMJwnjRUYX3WTJTF+YgLWGzM4qqzGNdPyR/M6LoUDriXj
Xz1dCDqEPORrrU2I8a4B3um3rn7kDeZXr816oHZjwKpwdi/XFwkD29w0KKLK
cNPfs2tx3HoAkKdEEQiKhT5jKTokTs4o/seWYDsqSovaNc65moCMixjIj8cZ
byeiDP31LXcgG3dDjrSv6LgInud5lpm5ZW7GQT7Zsz0WU2y56FSdNd9nLA8Y
WUwEHkFQ2NOHxCVW99WusmadwYCAVHIklrwdOpq76yhAMQeqWwwTBFPdY4Fl
WlKh/aKqd7cKj6Sw4urPstAHgM99sr0eERyFAC37DJC63IuiD0Wic1sp1Ew7
MWXc53KiLSMmRwoACpasDrDJ6T8U2IV/C13iD5S9lH+oRaAOXuwzsST9mNIm
XNMIg1g+vsTZtNTNoKIEZfSf/xGrNm3KO8VjaZJrN+2DEAQicKAhc5MDYHQQ
GD6fLQ3VZ2hwCH2cmFIvkkEQs7niRaLcVgRf1GV9mJOTu6x9rvNz77D1AXRY
SYZicocD58Nv15CmNg141p++5gj8PiwDS3XdlMj2T5f4L6LkHIjlwm6HCker
Z5TTORYWjdqawZDVB233yKndKYXVUkuBDdo4LrMqMLevzOYgMIME+cCME5+2
dJ3Ju+bdoQInXm1K23OM7u07Sw2eCdSJf/UUoCuSgjivhRY5+iuPyHKFWIs9
iz4tveCzgGEUBiFJ9+wJbWqZky+rDpLJtqFfcTL7wbDYBwIuJQhfsgNKfPrA
mK4K+fRANU11hI4fLqSo5v9uX/C4J7KRN0iZqPs8YuTZWFav9aJcYd/LnvdE
xNSIDgF3/qyAwo8o7YGX0aVcsgsFIlVKK+zHvGfz/TFvxPMbO+w67rvBy/JP
8EBb45GCq9M1jqPT3iwawQ5kxkLUA2sF0KPWvGkzYFYOEJYava236OYjkeAd
nW7XGtpEyncwj+8EE5rnJbHVh3RQ8auLyyfRnPOp+O/B74h2NRb30oMSqbuO
XSQRNuQC1e4madYtPYGUuN/PrHaFfLlcStSfoJzQzN313c6wwHKwbkBown27
E/ttffnYZ733+EWJBz1tMxZKk4rN39a3jWnScUDQNjy/wZ+FJY7tNF7tFICE
aIsBRsCcRrs6Y8XTpWtsz/jnl07CdkOheNxhn0ebeq7hAJsWmMznI1M3ECsI
K/8u5D04VyxEB9mxWNVAtIVpWpFkmEjfK9rXjSuy84BMI2T7OhkV3TscnU/i
6OIlr0MEpYKBqnWt+M9aEVKazkRdZ9LVCsXw1dllvlQoGU347SSnMBgMLYd6
Tfb78SEqlsJVGlPou9FGRhQkykgfesfgTRkgUHPVJOEPBFPbFNkKj8Y6vlHx
+oyqyiGH3ODmKUx/VW4/ugdAuezFK4ejqLm/7+aE/IypIf26pkfaf1EVIQXT
PldjOUPTooEt0Su7e8o+ELcjC31iXdCBLhV8DGWQpC4N3GEesqz0fbYu70KY
7nCEWi8Fm4nwjhxce98ZPYqC8cUzqV5Mp+DhqOhdTIEZ+cGxtO++kau3LNjn
YFoN+tteQvH/0EA4ucInIiuYP/NDsyrbbFkU2FndRcuQzezmMjwTNnyW5nAm
qolxRHdXAq6mvVlcTM7hQ0wu3A1hhCpu7hE6MzfggfbhFPSPz31bzBCN24wx
JaveyiGhS2UASSvfHRMZGypHKx/q1fo3Mw3M2WWV3E+qbV6Ok0YFsc16XRVv
1NHxDw3iPH8yqvQY+VbaP0qvChU1Key9L871IumK3fHg5qAprpbD6K0iRaCr
7jtj5pRdQF5spmqP5BxA7ZlS3zzR7tZlWdEogXdsWCr8gbkX8F4+z+do2eGQ
T1jYCTJXgYS/yTw2XLnp5yexmB/nnZsakh6NWU9WAPFfSoycVaBeqp05H8da
20BQCAhECjnM87WyQbvx+7OgrCs4F55rTNzcuOAz0vFM5J9dFv3LAkN9L9/p
LCHA/9qFd+L88I3gYeB+y+rpDyZKdu0JBwIcirNsA67C+GenpwegWc1AMUYu
YG08/HVGs1gHeyz1Y7IrmwmZCN+qVwC3ea8cqrhoS827hsFLfV/8+ov/2WfV
PZYDrH7WtqsagSLtp95hTxdVtrqJB9tABm5LFSlVKNBPRZWrziFABT1DFCP2
r28qjDqTGiCnz7gvAaS0bPQ6USRxZpp/6roB9LBmx8VZzfm9/PEfIZKcvALw
F6k7dE2F7ureHjRjsc0NpErXRbs5UiuTjWKZVAJXzvZ1oLxRbpNlNBP/t8mt
xx3kieVpGhUe4GPOnz7OHSbEHY0C3+Eum9ih18t2VlnMnQaa+ysWue7yYer9
rJzOvGWB3sheSjlpg9IlUv4Rbiw93o7W8JxbKReyuHJ0ZXGaLklPCu2xpNZF
LP/+W8pNh9QqAQ4EuS67WOKMQNiV7CBNdNV8jM9nUOSfAAw3f7b3OuiU1pK2
hVoKdk1tkgjiCkmvDPQsrtaxErtmYiUA8Os1GrozLNN103PJB92015QtTHSA
5r9p0rHBeT/PiajMnQ2s3QXLX/ifCqpwibhY6LWF0AYswVlLXmBPbFg2WgE5
dVduIGui/a4yDLHOT9JsLaQeOU5apokuebb5dXCGCWtZDJw4jsXVVmuEBVQ6
JhibrtCMviMPa7X0xQ+kmLzigDIq5io8UhS7YHsL05zwLjtDOQnqyUgljHli
Xjct6BlHu81pQ8NIEuVa4JOmhvOANqVKrPPo4GnHSUFx8ncujW+khXOwz49I
EUeszoVcZS+Yh0RjnuXtMBgEbHr7+AMKZddaHXhqLTu5xm5DBNDoyZMf2ZVS
D5BpEN72hwFDO6TLmFswyW/BBz9pzpsQ4AJv3LuBGzQ+eoCqs/TWCY9o1Ckt
xGzFz3vZVezCqS7km8tKX280el4/0mFtVXHZCCgqvZAscd4rvIT5bwFoaMe3
4C6bs2EAiQJ45simDYk970QpBvhwZmkEdXr54B2aKsHYa5lSnuek49iwK7Ou
wYbd+hcJaBuCVeOXQGVyXWh5uuvEsgfaY1+V8NT1u5Xft8PUxBgsvI+AmFKo
Bmpg5MW4uJwW33/Y4hG6uT2nKV7FhCXU2ck6yVVolExXoxoTeSy/Gx6k1Eyi
6pbu+ybOMTAl0I5n+YpMzLmCbafB/TLWuHHbNxA/zxTMzgfULkJ4ab8y17VE
jdGq//Fe9EyhdKaqIn4iJg7aFPMEKCqLoMTpCJmi17qjymQ0Z3KRLLtjDLbM
2Bb0SQkzjxcW1fGNI9FcuFjaGzpZAtotzUao0BwllR5oabFQUOe+K4A0kfci
+04UacImnyXGgJjTrOpO6iuJUwsfwqEh8+gqJqj9gpqWfVCZeiAGO8RSjEre
ofqKEiXTM+YQltmUc0lX5GvpFTpvBWlLAJAkaKhdRenbgoEK1S2iBMECKnqL
QuxIfCUb4zRcmOw8HxTw0bjtmeI25/cRSaED7ZV3apVDUJye36ltnl9KjU9s
/heX1GKzjDrs2dpoSR8AWLgx7AvyiNp/FDhoDYuyPxRMTAKdkp8XOgl+9nFH
sPWsL+G/kEJRBNlD37SpmMDV28DcMLiaxtnU3m2RkG8gq8XG7bB5m0D4ODu0
UH+KmDUc70CLGXzVOAjY6bmAGEpjH/pK1NP4LTT9NYdoRdGhypASD36rOLZB
E48PRpknzfoR62O7gxSkNb1Ltd1CVQvPpOmjhzSasQQdk53kngYKDOm9Fvdo
b4NGFlKk1L23WLf/e90uEO4sLa7gPXx7axBEQUmwws70HfW4vmQHsiNLeryw
DoOkCW0HnNx0jn3/2NDm9fSaAs3kfi8SMGFP1+OYS9iAS/WT+zCRFXY8fubR
dBM2g7wuL2mrnojc5WiePl1mzq9YYqW39fCwQX56ZOL9vVTx8Kv1Cz4W8Tm/
woh6LF5SYEQ5oiLkomfsTCpTFWXtl+D8dNPbrpcdyrHwsOu1yowZqlA6hchG
mYIJuJdfxEuaQdfW4Z01RC2I8a00bd5+eBoxpucEJ96PC3XBlLPZ17qZ9XpW
Gy13pqCvDkpvnj/Bw6CtY6rCf8jEDPTfv+758ScrB4jgpDus5XQYPQFsg4xB
Pu8D3b4IZd79hq9f4AaKDZOAYXJaySVHtd0xNukl9VZ1rUhURCEtsJeOdXyk
WURD2PIM/ldDm918S0QI/QiRDxupNBrRDhQqYgBgygk9ZK3K1qzSaDIN442R
BIa8PRiN1UkwTDYshWuJV4s96rho4IJ+Ymo5wHpme2Z85tZa+DkVlLHcWHBU
6khjklHlq96ETxNzZilFVq11rbJOucm/g83bKsWIflTqnrIGhCs/VLizldUJ
UD84XJLjhat9njuE5PW0tlHoGFBtST8BHRl+9IfbRHz/GoB7NNL2Bj7aUtf1
ZY1Jt5anaBowwF4hrRHDTQLWDdImINrSkSom13jrFkCsPdD288tln/WySG/2
O4nXbVODbcorZJ8tYKXlcLFPNRz4odfWAb75Nxgijo2fEoMpmuqUgkjmtJ2o
gBWDW8hoPju8Mib2NZTCzmtACT85PQhQqR65FyHXKdrS1Mh0m133AdsnNcdJ
QUGMUs83qs4qOPIoih3T1UmO5+3l1we7w9kTeBUDCNqgRy8DMXXVlWp+5x//
7+TT5ASsU1nD2qwjXbKilUrwV1dmg3rJVXqKZMRfjUKZ8FsF/meTJI2KAVf6
biD7svgCBoZXN2gSAmEXFs4Ltm/GxfEYIOZ+w5Y+Kpt00b+gmvFN4hK1ZOJT
IO9Kozs5Xf9UXtRgYIu6PfhkVwPPWSn4OZqmJ3zT2AL9rzvjYZXgcc2u6CeV
TuFrAM91uQBQdqcpYEoa0MdQ1+1Cwj7ZYNT5zd2rsRRRVcLcf0rjSwCunzh7
NquE8PxcC90d6ZurzIrufuBKqe0wWn1I0aVuKUxdTHngMm/GyxTPF1n5EKdA
n16vKk1foR9pRwGSR7ya2oASj0jjGRapkxOrxluSa+6Vsf37zHqbxBQ5dXgJ
nHlbuWbZ0Gts4FsEcHuAvwr1B8fTx4Ta4YWOZXSDJR/0+/SdGgN6PmYJqJEr
KWenMyRPVKpognImi1lZH7VbrOK6uZSv8YCWt0Fo4rwiN2IZcg1ZnIpUtE0/
pDa69JzsNdUELl7Xl6maGQnkZb8nTL+1+L+FQuApGLkH3cuGv0YMu/wpSJUE
WlRxr4cSPedUYd/QIy7LY+ywttAVMEZGCRX83HLqPZbFiJcpKktG9BGgMfP3
AH7Gmo7uEC6MI4Pc+wQfY0whaw2pxgnLUDeHAcooQNTH5kSfa4W9a9aUk115
eP3htS+SMjKUbQ73w71niGgSH9qQ9z9ZmOSIlwAWu3If0DtKlzNGyMdQlqpK
P5eG1b4YjrdQ/vsGmFxb+0i0lrNxZBHnVXfHFv1qD5Ves10uQ97yIDs2Rrso
qBfzlPuUdyEiy6mENgntOzQ3m/Hbug5hi7Ggkhp7l9p8MQuLB8gZxoM47Pjj
BNFAoCRlfZXA82E4v5syTjeG2Gh6j0qqi3+UkBlP4kIS8nTrfEd8+ghu20JH
foO+plL35CvuEq1WEPARcR0gu1DZKG5S8eMHJLJ/qLofEKxB14lvBlAjTpST
eZ8lHT+QqnhHU8u9LddHRrTgIn/eQ4+8orV0tCEoFdlaIvmmXctj0Qm7CjAm
wLgQ7k0QK6UGynvRvVgaMrjNhyDSJyTcGQ4yEtygN/xgu1lRWhCeSJmaLEZ+
ruW+etackbGn/7mAufuY05ge810bKhJF8/FqAPhcV4bwfxcttFAwWWSJ2aGB
GY0E6VnQplaeO1nsaurBK3DGi1E9Lxz78BJyQTGwG/TMiJjwLOThgTUJC1eA
9UWAU/4Tqe2qauJT3XsT439TqujVs6P6K3Mxs//dA5zUZou8+glMT3DDf6KT
qEImNxyoFiznnzrgzfqzheIyUcnTetTuyymwcCCkcEjg4tuf23DwzY+r7kwf
FvlLwow3N4b5QhYx6UMSvCnicPZG14s7eoa0TI1SlM7MxTmuZnR+m80eqrSM
ROj1CaISgvmL83FRnq/zqbmdnEUxA9xTXwRxnvURzEzy3RkKVg9By0/7wW6P
nZqPpKIeZkFZaFJ/mcMSapOqfk+2CiMbPIENjpq6/nSL1wIXWx9QBsG8A8SX
s780jHQtv+sd/6kaBnoBq/GiMjXqEFWSeZai7iyO4nztzUODjcOoivdFDDJd
m1oQB/oMYaRO9k+Lt/dHzsJ+1JPk7zsPGkK6iZOzUxR3sqnMaVQXSnOZi6uX
9ahxahPh8Np3fQ0T5b+IL8bBhgO8ilyLXSp9eRiLBdUwy/PYwLUABEV7SOpH
6Jehjurl2BHlkT6poRmLZf/EV1STXOSyxsZsS8FLDg0eHKHn1mMQPaXlXjqT
NUByZiaJ+KZGkTDqesZd/Eo+Rr4HLZpf7AMiRoUIZR9cjZ2Sb9bkv9Z36gdv
L7+d5cKtwGn5MTlefWFlaLDKj1fTl5vAQlYv/sM878TIEpunSJfrMuPbAt36
KtF5+FCyWDhcX8KXnzxKdR+fZuPmKGioJdMI0X2AzxqQl/cZPVw5N3i5VEp/
IiFPWMFfPmEvNM+R9pNJkZJKHdKjeasexCLZSpERznEQ1dOmuqlDveMySvxe
dXXumDYu8pUgc7LOBYeOEzkAphEavtTqSlycb7LXtca9dAdMcGzjUReMER5C
lZch0Kk2/vmSIo5X1sJwyNhXNjsK5+SsIJoJuVP5KQM1o1IpO2NbLF8UKjPl
rn2rEIwC9dDQnAbORcFrAK970qWmyYsszcq+Kz4LRUDZahxm9OAU+IEbo2k3
GBFMItkTrTabOAuy4i+xJJaCdwQju0siLcW/uG1eTAux6CnlQlan/mp03OP1
5wV+eRdxVk4DiGkiJNG2fl81pagR0yS+p03vTdHKV484QizgRk6QlUwsqDtS
z5w9J72FklUScht6F+QYZyFOg1macG+OxjnfuyXOtJA9j8I41vXAv+Tzus3v
muydSgRcoxMz0eHPQYo0f4jtEdeTIHRGQSmTRP1N/HxX4nZRwFrjUqhvUnBZ
aut22kx6crQwfb57Dbpjct177gfQI93BGD1OprjClWQznzBgxv/0tvJXfG/I
TKlviWQUEgur66CGSuEDrygWlg9LnDCwMLbhfrmMrJXNbUWUjcayMQpd5Qpq
EHD1wM4XCvoeeHF64UtK/Fw4bdOQNp2O+/ncVzQKEicKrNKMjEji1l0oESr8
f2i2g+jL/XX3X7zqKKCVTkK9nLFl4T5Qo7aZljDjNV2rzBq0Ckbq5XeKNIHp
ZqFZFTGz8UBixVgWq06QPwhjrfWaV1BRsyfLPQEFbHt8izlgpODQ23MOwbDK
RonMdEnHdQw3WFYxUyrY/0QxPBU+8TlzK7TRAKlr4KzshDLkx20S+RSz8VSv
mF4j2l62/5KmFR0zhsVepoP6uPgjKNKiI7qU4oF+Nzb/T8s3rOLNFEAbcEhT
xgt+GpS2PvSH93rxoSfUGJdOXMDRzX+CEOO3oHqtJpg/D4R1zbJgbbvA/fJp
SCFZdnATiLUcbQ0txGazvuMOiaAPH9U9gUQCEuSN00u73qcogoWYKM7i4E/j
gZZWAPUZoTOa08pD712+9l2jWTFHDnD/mAr1Gd2s/Ir08iAzHKrvTL5DCr+5
CfL9GcPHQNiGYB4tms5krc+8UGenb8Yzq865EoYRLv8mM2cpK9W4UaOxlz5H
jmOGkhZ9MYnSLJQYQxSf3RhaRKsewXxkTXK+3TlG7IUKOKML6RyQLyFk8nfT
xRsH1LzxyC1J6vaKx21uKKSl4g9Ik0hE/Jo5Da+VpxxVNLbtQdvNTXPfxCr0
oTcLVZ2DbVbbJic8M4J8Dt7nSAMlSQKyyIcWA5trJ74M8zrtr03d47hK4Eoz
Rt4AJz+vhj5g2U7fGaOWKhGcmQ1X2la78bDKYvcHK7dUQSsXBjwC0ONyjo7m
dlHO9FyRLwqaOhsEl652dwZpBz9w8fvO0TIEAJCboKM1AC5Z9HyA4WbnR7K8
05Yb6boBvG0TRzk189gm3R6I42WzRkP3xLvOqpQb9L2ApsmICa4p/jqXEoO9
47o9WSjyTrZpDHXGA4i25mcGDFKJSinl4aFJwmGZwBeC4K3tYUrkWsUD4LN5
m2E/1EP4r+nkKqfwxw7kSxlN6cltjsBn6e64/aZhXnwWUx6sOyeHwA6mP7GR
IELV5VCtkeMGqJmuf8iniwNuVB2etOpJe/A5y1wlPXOt2IPpdSlMv0YFX5Cu
iL8uQQiz3H4lLmSyPJS5MlLYuJinVDU3zrZbjYkHJXbOjewzgqaz++Hp5UPB
JrFxXl5sgncKmTPNMjvHQdK7ZctIMDZjelKlLSyOOUv2nCh/2izFXDh5+YpS
VaHqA5LzLQjbSRyn0s0nogk/jWjUxVEajRE/Zg/eow8Z46ZRUKIwXN+feBi8
Api+f8IluBgmInhT2iygyrQm3DeTerEOcM6fWQaC8NlnHQ6jXnDn+tB37dzg
6ty0FvjBIWHihzdK1Aja070rOPk731UzJ81+vaWlyHvZROMIHvKp8PJ9Wkss
1yOr/tJvTBb4QkkUeHwtWeUNPgmOSnnvzVBPWmRf2pJxfEr2yDV0fFTs3tcO
nkH/MlFdzPcUC8DWKZIej+uvGfMSi7Gs7v1eKCB3nGZ9T/AdhY3C0UunZvHJ
c78SdWC4tVY7Wrrx16a7EphkBTUt6J5RFH1FP2J8uXYmrvIf7om7DWTDrKil
jbLxk+kyAkW9RQlefy8NfX6lVEgFDSzCBtfJD4WpSfibrzDqysfKOTAcneMw
grvBfO/DIX+Fb5yFkio/2X5YFXuPqaEh0vujFUK3sZl3eVXB41oxi9FkBu9v
lKEJSKbAsJATCfo8FWCxF1dk5jTmS4qRhDdPB5vAhxYpxLjEik+liOSEdKd9
sR2a1sRCytbKoSU2X9IQ2WQ9lsusyi5IsH2o8uU8b0pBDpiJMzRcfcnGYuQX
U+Z/J2x+D9iM0D3ZCSUtAAgcc4HlqhOLviQFFU98shFI67OuwHafgNtkMSWv
Jvuf+ckxDPkkQMsQ4y/mLWamS8WYb2upltAnJ6W031Rqfy+KIFxHKBqdz68g
dCgXLgMuJv3mH/bHLanx59WtH2KU566EP9QM7NCjQzkaJFPQ2Gp8FW4TWIvI
NqgptgkY/o2VoRqtt7resloS3SJAPDshVeEvoGluVzwtmA7Mt/9VxxYBT/7t
7jFmHFgdlzOTEnDde1exUg8Jar1eLm3wtKJsKyTc+pZlx6EvKjij08m9JvBo
uLFp8fH/FmP+b/BAFLPuclra1URubjCZJSR01U5/7YU+pwvyf31iZLF9TSgO
qYhQ/9T/bUMOFz1Q6egGpntcpOM0xORCI62a/vmfhQXHCU5E7M9igQFMuXyd
J2ioD+ih2WaNlKZ4OpUpGi13mkTV5OOIIvPjUby6GZN+MEIh8Tv+hPo86uLO
SkvdpmdMsJ0LURhec0osx1ZP0HK6YuxJak+oYQqxHZWB81gmgltJQsfIcvJE
kggelz5arZsJffu6+QGJVA3YB2EFQmEeu/AWzhmcnBvHxk+UOATs3QTzCuCT
bB6sYnkHOIeyh0k+OiwwNNWZmoS8gXRDTecp8LOhmEYKpSHil/n0DSHSu+NQ
hQQyCiO3iV14Qcg0O8DUrFJyRoZInF84ranJyBllPyjuM8mANcQ34syq5OMr
qSQSEXX7ZbDtYISUCFtiHMxFcOLZ3M0Q5zvcbHouVIuW1KRyxI6xoiW9ZO30
jJP3KXQpKMn3j9qzpLZYzUtlEY8NNuWKCld83aHQ1xx6ztRiC6YjUrPuagEA
oxT9nb4xWd+q0Y5jCvqgLtUpyzZ3byceQd0cQ9Efg59Bq6E+4Zy59C6G7Sge
vnYxAUUM9OkKbu57ieuh+9jP+jOY6NM3TJj5xiXRn+43b96S8DheOppAxRdY
rETZX5uPL8kzV5A79E9LFVdMdIIfQkIFHFhaDajHUrbL+zv7Ttvai8xQ0nvp
I/Vot2Jb6cT2HesgZM3PqfKtgHVdLMSynKEnBWmgdYZdOcFx0PQfUMGB7yza
snSRWPOPivVFqXiGpnQNnxVEVkuDQHbzBz9jIkl1Z6S9G41CNhiBvJ1vD0Vz
6sipfXlIwvsyYLUPCfIWPE6oaVJwH/Kxc+7ScQ+YaI+rewEOyg2CuM+FlceS
jnCZGaSxPRGiZr8MKeaSp3vINhbPtSTk93JLEICkJq4JUDNU7AMG1/fejPae
9acyUQwpjRLUVRfaoUH3G86/k0zfVTourRxtbz2yKqBhSjBBHpkykXaUKCMW
yglASFi1nCD4wHbnoKW+K63VzRjaWTVkybxLE1Q0r6T40pU1bkUiAm9ExNkT
DTJy4Amf9x5i5hb7XpU2CCyZJnihAKZQKSny2X3ngoTdIiQWfwOUxTodOTO0
QF0vu6VvNvJ22mQjqM9VglE3e6/4MIPGm0gTJNVLO1IdYMKJ2apEYUsjGRQR
0FQKewqQxiaK1lBZkqjUwA9BDiM9w04le4tS66Ai0wyBrQv7kjp5hq6461h5
vLOiNa1n/gaqgsQzklRAOtl9KbZa+kWTPkd+Z3XE0W6hbTNmNGwZwt0Jchzt
N/2m8JrLz4XOLMIR3KKAEjqgp+hiLpX1I4eBzdGE8FfyQ1wq/LpksFkzUlNO
3P3BYIr6VkqeMifLgS7pfvLFK0qaAYEAWeY8dXaeTJ8GfLZPC5+IKNC967QL
KLm3KJiiVoP4tq/tYty7LoAk5HUCIc1O1003NGJCblcw+qC9EWa9x3bArHBn
gnHwStVSXGIDOQXPTehK5djyyBftG4sxdsC2TDxN6TqZoBPE1EK44PITYhLX
6Nva0RIKGTADGkMSFu40Sm9dBTitaLvf0aS2+kQGh+0zbze1oFV3KXnVI6wn
ZT63hLyHZnWYiEj4HPNLjyKKi+keW0Uscdlxjv5Z4kMEA1slx7Y8pWodCe6P
kjXteZARlmsj2aQnohWI/yOdPDpO0/ERhI4e7QSg9f8uCgf9WXGCutaHM2HZ
tr5BdboaTdqFno4C02dvt74hVdFUdcasBPqgfDpxZ0KogTiJT+U6gvUl9F3l
4lz7I9aESfvmazY6ZzVDe6bty9fxqg5G27HHZDuzqMkF98+roYreeI0s8oZV
Ahu5CwAIkBNQKmj1u5OoYcyBPjqliyTWZ0Pt4H9hSMJ0Lmu4/lzLbO0wtWU6
yQ+Ub/4WC+GxaEb+Hrk+mMNhEgR1Ii1Xv9LpdufeVdbhA7FQPP8lYiFPBfwx
9DkY9nC4PAbcgXx+PwybZSJCH/YE+sGrInTMMUxtm86wjRIqDwjK+/xlHjyY
2ITXTrX8uUJQeV7K23f8MXOyffYuDTkbQHmV5LdS2YA6h36s7cNNqUomPHNa
9Bl3wCeBSscVwl2J0Htowf+EVlAxqVggL+nk9UPq7BnZgjsqDMtAKAVsc01i
fgXY3pA5xHvGN3oNNYmZYcIJgnzDkMC7n/D0bSWnxSCLgH0/8I2ze2ngVofg
dSih3sy5nGTshVowzt//MIheRAU7p8zC2V70YruXEnW/eqep5oKFEqX8a4ID
H30CKPvs52RY3ZkdGJLZLknyHPHVuvZGRGCyTa81CynR/Vo3mPVcxhPrnAH7
Oy3TBrI4LAtEVFKGnzeoqHRn0m0sLW5xwByW9lFA+iwIZeVjuu/gOAsofH+G
cRbfjsc1W9SyQDSeGFQurXRfgv8/grI/jF+DB/di/fYTXzTS8Xk1IrxD3egj
EiBZhi5GCtwgNOzMCGlMsc9s6MEzP9YpT593/o58g02adOP2L+d801f7QKsX
XXB2fN/bhIwGP3fvdCnoNLRdeGycswQRMCvoRmZ7r9k8r9LWCe68Q33krBbk
MsvCxJ2etecH2DmFfOhSPZbx4B8wMaau4i6/5bT5WcQNJaqh2FRYhI7xm70v
Z5V6/AToWVBj9QbUBxDhSPIZD4sA+lmcIJ8cbALKd6LcY8n+ZXLV+9O+5PCp
8FULLzndmG/XfrmreydyImb6LuvGfxlSi/szNweQBXYvookdBtUUbApl8aol
UJ+DmmnqKPtcZPB6s9PlA8vrpGQO8Onph8nQNA4P2zuYjMxP0JnFuG1P0mXI
q3RxZEC/ruXReS7rxHG0IOavJuaNFkEufb9No/NSJl0K00EpmkzUSThH6POr
AuOccdxs8sSgTgrsFcxMyo3qTPgnV9PDoHPwFl8o3NbmxuTY56EQdR8iasyr
WidFp2xGz2nbVuVHPOwR8WOntlVzYEtFbi+eCWkDVoEb2XPIzm/RuacxTrCK
sGCVosPR/Jpy2FI/Jws1oSvumq2+vHcm8hQVSQ1Pa45FZDyx0oUSmzpZV93r
ix9xEi7D74ueMmbkkwaIGJwKQsD4M+xtCzIMYhQ7I+DfoEeyVUhF7lJ5DhkM
+r+f+0U921LViWs6qBsLciBLaCgBy6hOmC3L9Xjl5dBjxQgclB2ome4dIOWL
+mkxz1aCJSsGM9qq/N9Bd+AoHE1oJNaB/0TJZAPXb0QAwKVZYy+QTAN8Getd
zpGPKa7aS8ZU2cjbOgSTvgVJpj9H7uii36PLZb8wPxWIgQY1dKWZZ9evxdvj
3oQMixQwkEyIWg4lfa/RcQ3/LvyE5vqrS9RGhi5psJ5vZg4EnDXM1Hv2Tfm5
wKJVthhWcZDEjw5GSkCOLAQLRtfGfqqo/xegCYz734YzImgLQa3UzqDP1eyF
+19FTdHW8FeMB/1xwIMws8iFBRzprHbTq1FISbdGKdrLespylkG0oXb9bFPh
fHsf89wR+OyBrTxAUT8hWs6J9bTsSWvGyUbLX9eTqOW1jie2OhxHVA3acdVe
nRBkUl19g9zECJiPEoRpjw45GOtCWNar3iPqBFudFdI1lc8o3g1BC/j4Q3Eg
Q/XHHfrS1oItmOk3PrXYqLC+RzFt873mpHhbtdgVsFQmgcB9j1oQ7vRuNcwX
57ZEEaHRlYQKUV1/OJ1WfwHiGOaOC7YoAwohzCmeoS3Z31yqUWB7Xu2T+Hqz
9BJRVqKyu3HyM6x2rKYc8knEDI8FfMPrFYG2HLQuk1HHeoFFQvEZMzWawSnA
t4mH29QHQQ2yY7wMWmhY+GRHT4vvU3AG9X1qN6QAQ7DQoKewQpQOL/A+40Oa
D8QCTEw7SYxX+noo4KhsoezshsL4Mv396TmxvmEC36OP11UhFjTvw9u5OKBu
WFeEMtCA7isJYc+kLjlpEHOS8X51ZO0qKg2BG7Lzzq3MSf39E5jgB2Oeq/n/
HumUByroKumQSGaP5cRXEpPL9FSximiPHvyJkCW2vL9sTMGMbFYLG9VcfiCY
Uwx4wSP37AhZbzpEebOSG9TDPUE/ks7m8mRejkqKu0MBCQ97vDjDhU5ahWPy
hxW0vO3cDltmLrmrLzzCh4dxxGcaqWSBNnVcgWl1NGi2qu6hQxM1cCoMJj22
ZnPJybPQRV8AHCiPg36bHc18GdAB8ujyBE2oMwBcBsF2NvcYlRxvpPPIzRVw
kZuVWnePjMbtfS/GxPnfcYzv1gAEDjFxL1SfNyuSTGkUclG9LSY1Ggc4SCcp
zuzcRrwRAtNFv/08f01lO+Ogwk0exOk+Urkg6YMR5xYk3DpTJPnaNoYV+MHk
iKp77nb29yiMkXxQawMn60XuKdHVvAVpLud37C3dPem6fFK6g5RAqKBhhu0T
2njwY30WKE5my1RDSwVjxq/5gCyCw1zo6fHOZwUn3uvrwZ4+pCxLfIExq8z/
Hu8EgBZ2sAR8TQYifc3Rt37B6xqpiSYiWRnsg/UDkgcj4Aavxk74/cBeqwUN
IS+SqnVXlsEdq6cN27gyPdd9QCxJMeQpYsnjQ1yX+RMqaD1NsBj6HNowspDE
jfVUFhuPCTDhphPHfotUH2WIoCi1P9hvYRdVN2ZPmjLuIG5lwV7n+ge6Zjxn
qbItYkU/v/vb2o63t/wiqK+Z17dbd+L94UQlI0m/9Sl+7+YDiW4RlRhQKqA7
MyzWNdP6b/HxtHjXFsXWFSe8FqUFnMQR2vSHVKwKEgxY9fKmIpznY5y+o5ME
owPjxN10863V5GkzisU49pf3qlZ22hGrk/T8GjYb1wsNZ2wOp+6suoggevjF
/MaeLxfhHsQ92Ve31FhrX91zfkll+Dx2yIXR+FwKEmWJaBdKrfoyJJQAZHne
y2Y3HjkKtYaLOn583H2TMve9hU/y0gyH7iA2eKpPKMkwPuqKZvm4yhOn0iNA
uUx5v3pUMwsMu+45YUH7Z+2hxtZnUMPjLnvdKji6JTkXpuUaokwFpOzMCz4A
Xg50ottz63mNnT8ou4sIuf7zAmD6Bg5QWD4YwAD9pRMKvEwDMWxIVeJv9kui
56n+jzkW2LtdkyZ5vRFkjZvfP/in82KSAVTPyGYTtqWaPVwxO9c7fKeV1w7r
XKBfDE6PxLGm+V8UNIeTV/ijuygdrMznU9fAj43Mc9twN+ED6xuDKXI5Ve82
HyY9KJgiIyK3QKrjwhjGj9R3X/vSU5hdrA9xdJiqnw9/T1x2QeJJJAv0QLQ/
t4G+rEl6qCmhXNAVchT8h9jwNjF2IsuOfPHHESAU9cQl/mLqEz/RRyI1JVMI
ofZvCXwxXMnbJRH8OORDr4vtuoCnzzkrqrZZxz36P5huOWJgg3IfgxYksCoU
k31o0EQN2fTdZDdmaoMs4DTMc0fF+j3L8k1G+svye5a60Kyt4AeKt5Vo6sjk
MOgICiClwz3erL0u4gz/ZxLnjYSpfpuFtK//ytMzt5Nga/OyKgLYEjb4Yur+
fXJdrMbIFPAijeDg+6uvnKDYvq95IuCv7IodxpAY9mrUEYKk7Kg/FQvo+vyw
6Q7Wq5TxhPeubP+wVZs/1byvypxzps95AJPvPU7TTKBVD597OFbLCdVD22qD
dw8cx2pivJcITx2kMJmC7ZPg5VIa6EHXQeQwcc+rtmRbsTu2JawoaO9zxk4P
117Hnsw1PwOcKQZO9X60BfFP+3u2Yxm7WEt3aSvK/8PGHIi2FhksvE0AwAJv
pbYbkJ8Bj78+rhX4PsoM0qgaqY5pCoGZA18vSKikemor6dzpGdwmdUjfYO8z
PPGjeOC0N3hXVySoTyGdEzfHpmHN60Jk75V5LV2y6scjnsmg7yclZ1kBsLEh
Lo7p+jXikhaAp4tKAfpCJUtbyPG/gXpVPgsk1mNRU9SJK+CQUcv8hVZrazkF
PhI7ANJzSKM+vSqQ1Z2h/98rrEKaqCdhq2ayR/91yNZMJaoqXqbFmcWZi9xf
t6Z/XSOWwhsJQC5FAyzFE3zCFGwhO6qPzpIJZGwoojEmzGVMXvJ3SN485Fjp
K3EAEI9KeH8zw811+hFsKZshc/0pCaIhp+UfjyPIVZ0AggI8loeWHCKqqrav
1MQPWlnUNmCDPQgOGMKvZ1ynR5mev7MpWEeGjGh0At7qX3KBoOiapEA9z/q7
7XnnHR4XiWi2UOI4uDEhuJHYSd2BmRmcAMHQ/8+bY+l34FbLFD9ipz4m9KVQ
8vXt9oS7sPU0NyOTlwfwWhd6W7jhGX8iL0u6wJD9R4j1qVvuF72g5jUnoKpZ
2u/caF3/M1qMeiC5XaA3MY47H8/5U2x0E9MRUN7Sp2RtrtTXnUKdgCbs6+Dd
FIaHEOnC0sDGygRkLwzMehgnNNarXwXpNwjdhH6dEFeVrCo/78NctOwi8cUU
oUPhknevHbY9W5iHW3ZD0vzVQKCvGWkAEnNtzJEBGYX9cYO8oRMLJbGtwQkp
nwStdjGNA7mK9B14BRz25ALms1yYCMThDvxCNJk1c/oMDR1LIbfj12BsYK04
DqwcjE3crYUKGP8/+9vKEYfE/uBRREigAAQ8ShWHapT/VVg40/0HmzXSiSbu
P5VWtXQf9mqXCN3bMag0ljmin0NYRDI3z9bGzJQrP5AIUVwgyQTpssxCZn0m
61EJjIstCXEOr10TdPBvzwmUt3NSJN7LgGbRDhM5zxEzOBDSfr75Ggwqqd6E
NqxTq7OJeRXMvQtvAMDEw/pbCEBmUWsZyLTZtGuZs0dwvIJcjXJyf3Rf3Afy
fCH9N+gIoKLmNYfbEuN9J70sn41z8f2RiG56zMftDuYEVrZ/pF+yGzT0nggy
/6mQjBK0oz582MnDVVa7VOGe7C9Jad7df78RoMUOPVs7O1jEbqbv/oF1EfU0
Tpb5dA55Cjhss92nO8hkvXYzSXMqZW8uzpXiHhQgw9sAlVEntHXJZUgbOCcj
gw+XIryoU0edOVLre2t63JyUSE/0l/BUWep7E47e0brbxHJPYik6jgL5cZ6t
WHwLpYMcrVBNk1yr3XbNN1znrFGzI6p0uQNadC1oANchcJuqjk8E6QNV2XKS
hIgOoSCHiWzcj417UwOMjY9Ojh1+uicDgPVVZsg9CZd/3h5sm1YVAfB6/TSp
Mp6IBEysz5oyXPN0HzzSfrNjOovzkyVslzOdWYsDSuJFrmDVim+fvxFFJ0JG
DkbESxcz4/tViD/ztzMkDm4jicyxQ5F7jlV9VQlaOXctOSjmC+3bndJbT3Tn
SId6hMeUyYea16O5JeK1bAu2zjSqh3ypZMMYK6FwqWYITRu9N4AMmu2F3Wb5
mrZqoQyQBrVJauhEQ0HkW6BNJ2gMcP40p1LRc90Tw/ziznZIZZ6yftwSiY3X
BMJgSMv4IKKnsySbZHZjMUSovPnjlhBQdO7a7YO+pECS6oNfYxMznbffQ7U0
uQNuv3a/p8ZXAv+ZzQlU9f8PsM50Sv/0eLkz3N8TkCjrYp0oMBNWAl4IXwju
y0hcDmm1z6+B8fT2+niY4sIUftZi3+eBygVbluEdmW0QqjPUwiMMilGe9Xub
6VnhJ0jLZyAJvLXaS4+bnqlHwhQXBpcY87F4fd1nOfrtt/zTRzI4nNgv6got
oTa8q/or09RnIHzrplFWlYqrf9Sgk4cb4iSErzTYqRXwaZZ/J3lGAp/Yp9W7
kPTk0DkFfvR9ExT6l9Fnfi9iw4WzS0ccKtlnBJCNc8tsGAPx3T7zjB0UBzUV
GGh29Ek8plkT5uSACqDDt1KAieQlUUDz/9k5GMm4BSqo+VUmks1IZU1ROaGz
rt/Jh5lvEgBqk11tjyadphDIOnvUPyOWudmIH9CmyNsBUW09JK1BmhdcZ/oY
hxacYkP8zKgVxONsAehUukUirO7jIsGkx5n9Aizy2tT9PjbCwK0wffMO4AhZ
d/nQjc6S5Y9zTphwOCkpP8/0RU72twHj39eUBBenk0fFE64lgmdxI5AUO5nC
mCmPrRTxBgoMjluFQ8P13pfPhbn2sn2wbwR1V7KxGiM3L+VKQ/wNkrcZcST2
MA14ZwwVcHT6j6FiYgIIM3trdZMmJ+zNY5TBuCd9x/KBPqUNRgVubZULvgVd
nVzeOXXIu36jiPXniLA2BjGGbI6cGwnUdNKXoydFXBMzWPYkk6+wcwsAW3Iz
JrqTD01xO7B5HhcOR15RMrCTu1X3rTQcmSm6C/5tmjEbQqiUdo0FFiJMGCtj
DpxGTa1cythjW61edMZscQiH6S8MHPvGqJVq9JBUOfYuB0Pf0dRPpFTHlzzd
0FSDtErjU35RpekIlGVUEM7zAGTPLiHK8UfL2ShCO3tDl7G8wGbDdaus6rNx
wBbapY5NShiwNH3YqgluvYmtq2bY34DTdm67BXDkx3r87S5OU8XGSXQABv3l
39OcYY5pDqLutKpHTNv93X0N/RE5cr5tkzOg7iIeqofO6QeTqlZ039jcZDId
Ff2Er+iDez2pGuewABFNd/1xwCICUFMAAJanCuuhG9ubM8oLjuOwTah1o5qi
2+HkGXDoMs3IpRk7AzpFfmPXaRsUooyaF6RKiIjB76xYiEFq8hN53H6w1BDE
KhPxbTUqYlCQHYSr/pyONIdnWRp0nVasmYOKhZonP6Y72Gye6vYN/wP/drqv
LNcAYSw57HaDhKbOKGtc4MgMt07CeP4BYXRVX3pC6GJ0+63iVlrX3cVMrP4K
GWlw0UTVcnmk9xjEuoyGBA33AWNekKPENe4NH2/ck4pBBdfL0H4KS5ea2NGz
b1/CoeUfxAGxUVhQw97Gl9QzKa/xO9azdh/cCmI+c2gtnRHjrD0FZdYR6r5v
ebVrDj+KYwNpa+Zpzed1vHEPVbMTR+vKeVeWqtdBetBsC12s6T1zUew97xSC
AjMxpdMx7OnaBBWa+rh6zE0z0pup2d4+0DC5vJF7lOXx4uXgjp4udBsI34vu
4f5wjCJtlvQ0dtDpssvl6ST/rYbsBEjf6m/DtARORbaTpT2HWHumAh4PjFuh
OEhEk+2titKSwxTj/Ufg+mFW59a46qPxS3yO8nONOMlJ2V6znCfh/snD5pik
X3EJNbFdlSIuv1Cb3hbkvNnd8BDEwPpuUcw2n84pj314pAPv0DXj4ikzDs2W
+wYgIIy3ESpeWRc9+YEPdJ87dWqgurU7VeCaAehFLrK4w6aC092j0jlyU3u0
2oU4xSSDYYgE+1TUv00sgKJhaO7Lc8hRl55uSdFlo+7HR4qrbdwlNxdghaZg
Oh9XlptEb608N+5Oy2XcmwYYzWJUJsb8QHwdctODQqfx83+y3k2rQv7g6F9L
OmR0wdmvBUmJP6egqgapA9dnusGqrPQwYARWCfCWJty2pXB7OK/kvhDr4zIs
wJ2dZGdq7aucgLvAhNKXNY3JxDCcbYdUsObBnLjBMt91aS5Ml1ayAJvjf/BR
FkM8OkrmEcqo7B0FpRqwh7pezVoGVTbdl7Lvs3Hv8dP3HwhQEZx+LMm6yZ1H
dvzG5vxfjLwVOKzRigpRr82IgEihlWb1Eltr16DtafAtmbqvKFO/1WT1kfBJ
cpq1fY+jjXW6a+jSKLt/k35imXI2kxyFuaVSZK3FnDpgTMjk5/2nJ1y+JkaJ
dcOZ6kJIVJ4nLxy3YwNvOofc8ZKYHv3ID+coGFKRtHFJ0ke2Z2C5rLTYMVcv
pAasSSZn0353e5xd5Id4g5AIScHkpQRiYEjN8NmwvnXc4jwU1uRIr9vuhE7T
Q7SvygaYHMAwd7tZ1yVTu3RJ4LsMbjaqlq22kK5utXRQZ//NkpFqRYeQlP8p
GGRwPVjVqse9siN5oumYzB6qfNr00c9mTECNIZB1faK51zd8+6yzFaRLBqxj
BZyNdvbBilvsWA9Z3Ia8A17od9Q6Fes9zcP6SFrvgdW02onv0m+iWt1wBTIT
2mDZ5MhecJBk/umBKpf7PaarlelGqGwOCbwr04duvJCsbWjlNHtQ3mfvuVSp
kafmQr4lsfJZUL0/z8bBQiO2fcRpSHceevFntww0wMWCGEVSmfYE2mZNbKvs
iftsZhd7fWwBtgUx3y8ivqOfcoky0ESAJtF8anNIHSHcmLHGGCAB4MpEUYyA
v2SoOl8/lCRBqJ7zIt5IEu74B5rWkQgS0o317AacPyWu8vNLNIzKBhISGCm6
YgiiJWi31vhF+TvI6XRf0ByggKJ8GQT0cjddB1XehN2r/St2E2/hJ+q0HxNm
Qbi1vjYkm2P/1cVZiRcrWtYg1z/Sq0/1QWzDi7ZtsoQ3jznOTuL+w8D+fdth
VehhIGNi6LHg066ZpedrOxue1lD6dvBGM0En0KTde5g7dq2zAKc9HH+4XGom
J7nWmQGdWpb5Hs01mXkOyCe87yTfpVBkC3j/KPAL/TSwTJzqfUTF6XDNKxM3
vqSu6+0W1pZZ/V7RDUm6Trm69OZz6MJPe6qxwkbrzFzZjC/ibnYtc/8i1e+p
MGW61M058RzbIiL93kvUwBAZXeptoCSRRv/meGvOF4ddIpTsxV/o3oVfQ3/k
9Ge/saaz9HVT5H1l1+cdpKKc3WV5RHULNpizhMfnRH4vaTGblCIf3TJCWZH/
3glcEwKOhUqd2gSRNeOC6hmhZy8UxvqeJZmX/9AIl765aOR7ufHK3fsvuKQK
FAnP5jEskKQCDLFihA/RhBNLCUWV7LrsoiRnw9QP/NlRuxPInjlZ9odkTJqE
5zX8BEX34DJYx8zlXcmrfZppqqmW4e6RMPQBDleWBe3Cu+CHSCrm6Ma6VYtf
e0xtb/UDs73qJXViiKT138nK6pRGyvKjhBsFtnfmoz6shs/9P7xsSJ90xroM
r5XXlOAoQtGdD8F++MBT8c3d17lN/fA7oBFraxz4CahBHtaXD7aLZrLEMoBp
EIChaygvhmrLJNhE7fkxA2/8Gi7USTV1n+cF6tVjdmlBndIHGA+qHcmgJd63
UV25tQB4n7YE8MjUczGgCkONNEOwBZCSbbpvnW2rA37H81JyZTkTlnU3kG6e
TSluCnnjPHr2bWew7HA0WF9/9be7vbhva00weOh2UcBGQUxvhBZSpNXsjwV1
H7X8jz/ZFjKd7ST4ZX4rmksq8g5Q25o8iVDazX7kX3+7ZEdbHVfWm7cgCEWl
u9AkS6FusxpqU8Kt+Dui5SDg9NFQ4jG8h2+33D5yLF2eNCKHCczVQCigV3kw
wiH+Y6s65gPnJzs/473KM+bIheORdXRXpOh+J66ixkWyzHZgTA5O/A52d9J+
naUw+5KGTQtEWXLFLV4N4T5KaYgJFwwgblxsin16KbpILlvrr7gAe7UVuID6
1HwDqM8QLs49cxyJMQ/LZQXj6IbnikXr3hHF6RxocJ4kn3n+1XvtzHic4Eld
PkSz3RBeDtDO4A5zJK+eZ7fzTGdMTOsPykx4IiqRawO4aw5aL+UMp2ONdkMy
BHMEatJJ0Vwvh2b2Yt1eU6MKOaxDyddEeuuxLZ7AMceFh3KLYeYO7FJzMWxV
lagxUGlndfMCqM9xukL/+UrDk5gCQdIp1M2KJV9jw2bLz9sqzTJ8NdK7HZ5E
vEpeX858GMp9eWrRCitRJ4njdhCpT8YTXrP/Oqu1z7erE7TwpH2/TFJXcc2e
YrD4ZdAcJzDD4DkUnGOMc+BFRSKF/Io2pK7QECmpmybgQ7N/mv4Zc/bhR/XB
TsezHcKYPOGX3mFKbUsjtfbjuaVB5oVmor39WdubvqGsFQzzvXrM5qxtzkO2
YuPCeakUpjOoaYwvkGooAi32jAtUM4yMoSkhG1z0NnUy4D+H+/8P2DKBuRTT
1O6cbK7/aaZuVwTC1NWGC027a8RvO03YpWktFwm6OTEld8JcuRdMCGEt8b2U
sctg/0d1CkYxD8PjgAdrFv2ws1bP2jLq8nv7kpwH94f3n9oNGX5S7efpE+2v
rr0w1yvcqJcaHFjYqI92E8/ZPtZkiXL2mDGyb0u6OCV5qF4qMkP8dNDaTD3V
vbte2Hbm/TiHWReVKD07U7vhyNnKmGya9s0t90EEuVW6DHDz28qk5qSxJ6Pu
VpUhOGMDV0Hjs/lsmHlWrMb8RCGuk04EMAvJOJfrbcWUsgxvYd7gTh4ohG3B
x/SjvMoWHDUq1jHhsTw5rTJDrW8DRW526c83vxvteMCdolBeuiAcRveWXfjK
Fl1ER27Wkrf6W6HZcQ6TfQ0VEbP1x0hZyDX4g6pW4HKYneTBcgLotZWydZNP
to0/Js4AjK8LBDVpm7L10/gij+/bkLtouEV0tDJCW4N9wMJIzDb2muoVGARN
WG2pWn5gcLln1oRTTY0Lr0L+r29dARIXprY5jxUKM9gvBJPopcHwSLy7HAXl
J2A4mHmdgTWlEDszNI34SSLtqaMUvN7j/H7HHliPpA+1knXqV3GAIB6ab+cB
9YJuATPgihU4hHRrL5ha2/532NtmZr1eJUl9Z2xPsT3ft+63g4WZokdHoueD
pzlvVzMidVRV/KByCZJyVnOM+3sKW8q4KXxIiJoW0prnvM6sburBnGLB8fDZ
aZTEskDaa33Va0DPC2Hd9EwFfmYveko2P2Vzbct82rCSXjDRXLgcFL6r+myd
2iL5uDVjfjkJfl8fInrtTA1+GEweN8pjtzk6za9+xtFMkLO3+mknd0hBFAeZ
p9ZP1ezduqFLR31J1VqU77oKjDrYjbxnXHPOxEHdMJ9FxTKjoheZ/FKpn/8L
Daz/y1EcXPtiGI9ZCa4PHMDQi/QCfcH2n6WC5u2L6ZfngBcERz6VVuu5IiN7
alwa5hUzYoINc3wkUYEijJFEGYo2nHLo/2MFh5yRCvapWLyOp4lGipw7F/H6
ZUyBX+Zy+WQceZYV5Jt3t283w08wS2NeDEUa4p717ShWTnXsQV5k6o11lEa+
qVBy+BzKONz/XwRkgWkbXz+MxykMRUyo1IPHL6QINmfOKsvhFRPXi+9g3Upl
TeGHTaCdXJqSk7sndE3pAJDanQfyyxA4gdwg2jcbQBz7ZOndJuT9yRsdo3Je
GWMAEtCVCkyERcuQoTc2O6KWQlAxIxk5ZbNbl4g1F6RbeKRJJLLVuyZ9ECek
uCwhXnbfYQ1un/qZnYCzTSVSklLeFW7HQatCaGN/JIwlMSxw1mx/cRU5MTlb
T91+1UlDR2FG5xaWxQtvGZ3fTVWz67DdXEVAIgdCIFzvuFK2kea/LtdoEn3L
Fw6nu9K01D/3h8XQqhARv/rH7tM0dVwxD9krzuB/qIkRAAoxdRx7OX8D3gy9
sDhcWEz7PEG1GoPlXjZiPq5LSZHF2YZRXuVtufwOwZ4SDIS7UgOTZZpOqmGh
Rpnf1+lVHKbArFYpfzYw/dJtezbypycmtriOdzyu6M0ttPEjnXiieIATjpU0
7b5mvaQvWruVyAQhZMyEkNviLmgtUvVNZq/nU3AikhmVv0p+LOqbivYKjNNp
NZvp9yEhq22Ddlhdpafil4kWiORnibxhlzNOXBLHtLJFeJeplyWgFXPNVkLD
ztQogxPZxFAnCVsn9Aq2TsTJz/1w4JYI/xv4lj3klPfR360mdgJzdkXfuTYu
eKeEgA/TNksmC9f3ot+gBzGE7Ixdpmx+FtH9CD9fkFA8z8A5ZfZAQxCPtBtY
cNa+/U0+t/8E09Uh84k4OU1mCo43hDFZX3vGY3tzXZkhL6Dm/bTNytxuooiP
ayfPsFjl82n7xz24/OIUx9gZDgcE3E0iShDEAwH5bImdhokGYn5iGOPJ9r58
/LYA7hk2/Cti7e/PvT3ocwjbnPTIWH9N2tetRYJ/xYRfl59Zd8cbM9uyDD7L
75xkZzV3nzbSC1f/89kOXNaP0uqv0YLMCBadSrGgqR2qfwHequSFh3/5q6W+
sDf8xxQweIvBFT6TXSese9Kcv3JabZVjH4w3DsVgbL3817DIR9RuNzc7GDnV
+3dqLnH3h1KsfouAayfgVoKNM6dqpIsrFyxsYB8e13pVydHd/xeF99GAaDFO
O3Gobds+4894fPB8Ys57R/ZF/3vpPUjccBhQBUN7E1gJjNnfn1jUcyKOJQzo
FYPRAVxBjQpCYsbxYAIw9XSXoqfKzS8wSPpDrRqyUhG2V/DTec4MDc88XuxS
eb5T2iP3C17LHFCKD+p18nF1ibEhiJVKdBDVk8zBQUcJGdOb6lBJIxo1/Hys
B+C+yfq/gFjVVmXl3h6YyHEdhI5OHNH98NzwzsbV3VzYZvPiJwh63W4rPTzG
yE/evqXT4aFzwyVJJnS43EHDTEAQ05C88j0/HkhTRhF4HgH5Oqu9chbeEJi5
IliLOc9lqO2RuB9sjcvee7AF5tyugq96QL9KJZWlEZk7WqMTuGcDOBpgAPCj
vI7LTI8dXEysqyBke6qTRbUHNmaVZxsz0UfkX8MLmFHzWBCggU4c5iLgmzyU
bu7pbK19O1u8+DEgfVmZghPpmTfvmAMa44LCJaJUNd6lPV3pDjWf/onmqsPf
cDWqTMbAB54im2rFZpRARnALmLSOWadLBnsMKifkQPZSIDETZv2rSMO6Sn+N
8hCYtE2p1FDtO/Ar7mF5UdrPSgz86xeXbQQiyn23RqcnIRa2sfIFeSpGsIYf
wWvJds0ADjEzXux/I8fuf1V061kVYG/0gKvfFB2qu2RaMK96OhPR6D2+cCAC
m+rjr/zFtSNGprJ0j9u/IlbsfFn1aWOrDTyeWQftww3XFDcPMdFn+jHzigXq
H2iWe0l2YmC22nHt3BzVkhCPp1AP4aUULdNBQBCc4S78iGYVwjKm/srMLYIu
LIGfWrhKhvPYECetAAp9TYEYARJt2IWSxuiJ1QdOXh/hDLWKRk8qUWOXzlNP
mE60nUmCOVLRnZz0fyZbR1DTaz19ns3OTqcmTIkWEoWwS+VpWDZUPMPQh0to
0iYwakVjUzvfGy7ZPqj9o4Kivzf1KxxIj5QaqBaa4OuQZLt/kFpmS4ZPnoqn
6A4UnVLiVW3hkUn1R321fdyxiUNBy7NF4xXRyRjLl3LmxGnYNL/0z6oUL8wr
80fn0EZF797MJOLOE2aA6d8dPkBgzytPI8KMrQaZ/V5iFxm7UU236eiL8Dev
SCoDTDejdVM/7mnEbK9dD5Pb8lhoGtefNEyLTmh/qZtosicz6IG9Suz+jSa1
2x3YwhwAMtR4GsF7n3Ziyei83FFWHFd5tglwC43k8EaI18fcdhbF9bcnDQs2
kqF6eB4qwOyDm95A6vny3J1chp+67bDOfkVb0/eo/hjPNWErtwwFtv2K1mg4
HN5xnzobH+sMCgaiiNB8124LFrdlJ+CDpEGoFx6SpX7KprH0tX1Xf8DioQCu
DE30zG+PkjSQOFBOkYFeWcgO41EISdTrKNTOSQrup1lmK8Dsm/jIG3U+SWxk
qt1L1LtAa+sw6XF5hwIOeb2/lcFvASx35DnCSwfzFDm7vZjHoRtA8Kq32z2J
5LN0fHGlmHHtBq3g6WKiECPuuR3EfEOg0uviEsG/6nHJKMNu/Hi72oduUCkB
u5reT3gy6Jtb6fnjHG/1R3EAB0GQvv3stJyztHOHZQnMfEdupU+ItDQYVg1A
J8Woe+do8RBsJwfTd74ueYtyZrbD7ipLIlF3XCGCYFzfl/X79+p4ZzF5TXHD
eqfXKtgYzRC2XUEOhpHbXOkHixeLVohlAlAn9VPonVLMO0wPi2kDlCbyMFGq
Iev60nw0tcS8IztehjwOMnjyHv0ModtmPbaG1DMOpP/x9UYtHUDLGBzAT0md
ocXfYNbgMpSL3sF8Qj2gKFItJV0gSIo6cWsE5uNke/Yx0B8D5O40Mas7k2yI
4OPwMSxzo8dQzE9J6zXkOduXxaNq6I7elZygrdD16IPxyzVJC7L779p+YtgT
9ibYGQAcokdwU3gvP8JAphzDcA8ZtO/3Z/0SB25l2DEEA/KvFVzMYn8Qs6nR
4oTCS+Fty61WItXnuOafhIahBZc34NuuTO9QwB+sUnNy12tZlVNH85VFdzsQ
CjcE+s+3zWr3J0ac9tUK0nhnyIO1fc+K5AH1kCqmqRSOip+RFEBnkJ6DEmbu
UpfQ8XYXhrYxEWX3ueVmFZv4e/OG34aeC5gdZa8HmKoojDoV78tt8PsQlhUS
ptPfU0Gw39ZJEz3U8NZ2+vNtbvOcIBaIsZGzhAKc8xTE9v0JQpYkQCG/h5yN
/yCOxdte6rk/2hH1oA0KXquw+8QJpe8541O6hu1t8BA4XDAjxcOXVE9TOWsA
ZuoAdgs0tV2g+SYJdfssIt2QFDftCeMHeadjDgC49tNlnaromxrn0oNo0KCF
nuIiqjaiYLeL//sWIYrlwJ2qZQn9TOecaHTZ3j2/VxA2HfG3/SOSy73GRgZZ
nNCbA79cmAUbGaAkY7ZGvAJa1BNs5NDBh8UaZvSNp5HuAHQqjkdOnvULhF/o
L73STD42tUCrzFNS/QbpzwbteXJTrMVgzZwhNT6qQieH//+1yozc8dIp75ES
eCbncP7DmsAi8/suic3QBdQW0CIZRZzVVuFEgT2fLrnv83q29b6pnLkKLpEi
REJERdgVhiIjV96WTTxIbVHAminOnnVedzHHAHeh6hE3ddVtJ/bfbYXkEcXp
1qnJ5AWCUFZy1ZyZM03Wi5uamRBkMp9J/ktELQBOfzcROrNqTcrP3K8NUdx6
eqcSgbtanPItrh/oMq8Zi9tdbpX4WDM7V8R8M93o0MCOOrUQSjKsZjVMywvv
UAyQPKlyIXGcAtsa2kuC+4GAYJ0nlf5L4YqwaWzDLEfux+M/I2LFk+laE0r7
ltkSXf/WIZssKp0Ss+4chxukYHJgeT9LdJSPu07KDUp+GTKl9SkgZUw9n1JA
BkU1qm5/GRnzxMZ/VgbwHyPsiZ6pbYQzuR7DyU8/Jr/ZbywdhTWHXxKooAlU
HtRMPPVCx3+3NpiDfqTF7QU6S/ktqJi5Y7VI2YIl/Dqj1Xs8WceHCAAwDAIl
sfstf60nICr0hdCs/p/zssXrZuQvA+EY9iVOZFIOAF0ZemifY7PPYCDFU+B3
QISbyJnPirviowlpz/eotWJgFPjptbvqC6Cq70A5YeJxo4tiFhFvgUMV1pCg
CoExcoDvAAsrOJJ0y48p8GOCyutj9GmRy6lzdb5I/H+2//XgqzbqpNZyHnVV
2cpru9IrA4p8sLMLQGfJaUtaETaNvhiHJTCzwCBu5/lSd1+wSBhTE4k7pSrT
JLTGOOvD/jaSECgMrB+bc/fGMKlWVqu9prFoZ1ik7NZ6dtR6PwrrpxjSxbJW
AlTCBxnrwyllbqWZEH0kmEboZO8r7wVlu9OT1Er2irrpnSXe3c430Lmh3W90
pcusm3r1IcrB2eEIi7V6Fb4KSxz6/rPRkfDLhGCLHJZ6ntCsVmFbhTQwrf8s
y8QzJdzBuQBhvRaW2s+5n9893EYZLyg0wbQhU/hdjWYy7QZQ9oc9lsNvNPOy
DGEyN3GGLS6l9mkbJziRPi2Ip6tQ0DYt0kml9cMzeil4Ujw7cRFIjDhkEnBO
PH7UtJlsOKooUxL6yw/8bV5s0H1PUnDqrHu4YcDdoS6WDWxrAMh0sd0NQcoo
ESRHoMwJhRwHAXtuZtJVQNICPbTunl9MLTpc4j/iJFASfx89/sjImPPT7jGe
4GINa+jwtsmrwWiUb4HOzfJ/0SCG1w4VXpBAWVLFrYtvG0AfV/SS77K8XlQQ
x6oahajO/r9xqz8S1Yimla2N8A3QNZpS4J/jFsYRJWeSb61EVuPJSDPvGLuQ
VGDWnUF96YN4gMuvC2JQMoJgkXnfmZ3XfW0OTpiTb4tGiWppGDdNtZnpwjwz
Y0xkIDKFHToMyyQJex1dgpk62C0TbTGOolyjE0nsLCGX06cRkw/S5g9kcEnR
ucHTzOKDAdNMd7EwqIpNWLTMyQ6OW5+14+1Th2Uc+7tW90/ToGgyfso/CinF
MVJnxz0qdRdVd7miQrgLeaxtyE0cv1N4r5xM490ELWxJYkDj4oRwE28LiAkT
IkdvYV3sJmIBWZvFgeTXZRRi3uIrQ9mCLbbrq7jxTae2c2y+b7A1JJlTZnIq
hHWHIAz7ikZC/mVS+StMDLhy6KrfJ853k8ZdePeDeZ0DMdM4JVr+b7fR3Ius
b/RHIMLYLZJXWkGleaPm7hVQsIq7Oc9H6GAkcOU/avYGn5652ScQIDP6eppj
1CxSuWR8dpknOuVgAFcW7bCzYctz1d8Xqg4rEPmftrYyVDs/xh7lLk+XbmCO
Rn2mVyUj0dUSks3hbmtHfViprgZyvmsc+e0rSq6ywj/PwUXjIOTnvpKwHanS
oC9seVY5GkJq4xCh3YDoP77p23i5s8GETy3EBbGeCKLIAG7aaKw4qLmelXcU
ILym9puaYIlnqP8yDFIczKgiwIy9e0xXSQTkD/M37gFHWVWUsPw6NHyhIrp/
i+2t5fqIDMLBoHzN9TgHVQp6C1s0MdnVVMzYd2pxdZUd6AJT8laD7CtxSWB5
KfnrZOYt+sp7J/a3Dbk9CuRzTMrz4V/jPPqb9bgj4k3TFpnbSkuCM3N+xhqW
FYFo2X3/c0I5IZt0TVhzgh5eZKR6CcVdNoITsU2XGALaw2x4c+76ZFL45EJg
OrV+dU4JZQTa4OIg81QytUYZHYwoX0kNGYD6nHfvyStw56/E+wXuNL53jcVw
5qVuYXzTcFfPQW7kVoJ20z0N7CTCTd4cqGYA38E7J5MYmIRc+fepzuNtenHm
GP88PJYZGAUQAG/43//S790GHGqnOSWthD3wHeNHwySnloeyqdMsZO5nqRQ9
/BdplrNoipzzmo3Imd/YCsqY/KWTRaUYTZQCaYqerxg9ouFHdSA0iIiNK5+w
DpNSTHcFIBok4E7OzfZKKdX7bxMLAFkWRJFPTcQxrpWlc1VqHnMVER36ECGp
D7A4B0RxzTqaVHUzg7AZ4EOZCxThnr62l1WB7dPYhipFmXEYhFjYydYtncKG
J/1lMiok0WKXrOC2Bm5CLy+OAj0VzXKDLqo73strMa13c+3doxLkPu1a1Rs4
mO4cOzroeG5B6tCgAGbXpxSzmJ6ZsNMte6NNtsspi+lSrxLYpZZe9Q1lCCHc
TP1TntoNfLpXlBMhmqQDNpossQKoKlZl7eUfxORNLly1cZGEgAv5WpVMOd5H
E6HEgcm65TAI9DOLVTQiQKq36sTzEldT9eHYXfzjERmDeiWXZiNXcAebGPj9
WvmhgtY/Jtjkp8tsg5r6DtGdb7IBd9AtDpM9cDAG0iKSdyu7rmJPKm1oavpI
iCZQMkUbQYAwmzjpMW+zqTz/fZ9zD4IbsFj3B03JPZEyaRnA61A/S0bz79Ju
TLKJeZE6O61HLVu+DUD8qH8gfnMH52oc4VG7c8w9cl8lzrqwCMXyg7EvbHwe
AexibqXNvJbYwGLfCKiSeTZPDy11gvGEArki6fJAyFw/4WKgWAXmKhIQspyN
8+RIFvFdvdNptkqjvCK9TqPonesq3NrjmibQD8KviuNUJHYkcNIpiVgklsgJ
OWiEpFaox7R5+fZlEyGpIxx481XCJJTFAYnDDR2k/gRQnAip4qNO3Eax+jPa
FK9SNSX5FOo/2q9dNdZmal8I96cQtuP3WOO8k4XRn3fmYfsfG3NEBK0p2b90
YWAcKWWTpAyjKP2L5L2+W6OWQBQzk4pPXG+H/vTPJSvJFDesBkO1cB5ILKBE
B+OyK6uHyA1S3dVF1EbdOKaCY7IZAlxYsoDe00DntbPDaJSjmY6Xj2sKjYJF
cVC0jPo1pGFCRVuqYmxdoSIzfYv+XtiBekztrFdfFkqbQpXWfK3BqoSDWB7w
DpjSZ7PWrXsDU98+JiIRpsJZ62ZEDcwBZM7RW/x7JME3RpfiTww/5AEVSX59
IhqL7b8e1bDz9BLRFxOFIn5EHR1reyhAO5R0h4FID3EW7HD//NDtT8baD6RP
5edt6L333ZrTwXrLk4o92C5RuL97X6MB7z9czflswufRjZovBItslTJkW4Ll
2JmImfRmxb7rrhDVH8nNeWbS7P2/T0dGbkjKG9nXPV2aO7+4Pxo1ZDkF8MV0
L3pnBklCIQFsrcrxlIR/qN5NuopbOw6bca9OqiN4ocUeMWQ0FslG7Tb/gXhP
fOelVu3mTayiqbKt/JVZZcwE1KOwCRDMuerc9qI4Hb5+315y/wdEHceeFaba
5IHRers3k4oLTzKZR03Qb6RDOjZszNButL9znIYAAWcgyM/LYhRAVsTEMoQg
8Rg56B6nAc0uf/9gOfCeT4kJZ0jZqTQUk5Mo9U5xBemcAqWhd0g+DnW5ymHu
7E+hf0//W4kX88lBBlHydoaGNlZnScXRd50JVqbMNwzGqzoLAFhdMFWahbqv
nlRUTOccNjNzObFvy2sfQ5REYPH/lf4q8OflZL7L0QNBvfOX4eoOsLJnQLv9
zG13kBqDCBnLxmoOQbEY1epsGA/HRsZQEDyHdiNKJ4cGd9RG0mj+OJ2fi1V+
SxmwQI0rhNOQ+KhAfDWOtaCMIedRQ26aZdEuwVKFGs2kiw0oOsLIZqiGEEMn
xzcMrv2hSg0aDZqHbDnn8aIYL731GpcI8rSpyf45+su0Dd6qeWIKJzcvZphL
G5zifm/xNNJ7CTI6cfnEuIrjpYExpNf4WRxDaoZIQRAD/CW4CECs2KZt3EjQ
PlqJsr5RLSIEHBf87DstHrhAA9QyYalIlW0smOiwZX3KlLPiIY/0tm0M3Wvi
nYrw55TdwZ1Quedcc2jH2RhA8jApGBF+cC0zhDfDnkDj7WhnwhomhUgNflSG
FnoqNRVRQSzEbF9das2H3Z15+hl65qn7t86Qrcb/RllSVdr2tfRJN3Z8JrsH
axOd3y1hPtgSUHNEwN+QH+cyLeSLxq4PhvtrCd7Mo5yNIO0e0hPuk9j8G+Ct
zG5rN75vIJoSoIGDCMW26kwRz0VBsNSdRxuYOc89IZ8O5ppcvzVdurWeNDpq
I0biH8RY6lBrhewgJQyC4nPxTXIh1rHXInN31SwpC+mhhq3HgA7fYlOeNqtB
e0snIcAzXTVWrWY18nclntYcSVEspvpP/YvXqHNoCP417EMIuOhb+J+luYPD
u5Z/V0tBWZthNlRtG6uOhYiUNqb+Njur+Up9blDux92pu/Tzj/+9ImqWbbAb
gXiGAiy+C8jug+8SjOg7v41rBTn60fd6LWtlOSJZBhMnnesPyeyPoybNp/Dd
96ujmK5E4YVarWQQeaRawUuphQjwW+Rsm62aDbw3J4HVBcLVizU0F7JpIrk2
r2MkpyTURv0j7+EdXMMLHhGu9uSiSdMtfKbhtqMdyzOFFyhXL67QeUq4SkEd
mzkYf1DeQkU0IuoJeD4qXjLNNGAV3S+nQxSUnhfsBCRIuMl/NQgWxP2Dmp67
dzUniEbxVD0rG9tPaawbtgvpZglTeQX5xdpIC5n0P/9R+ga//m6jm7Ie5Rad
h0o3eaDuh3d1U2w7rcz7eUAz0yDDN7bCBWU8yqDgWt6ktbgDnNR+xFDV7QGT
bLUPLdqi5YIOPv1Cmlp1g0k5C23UYBccfI8x3wvxSpTOGUY7gf0BmAD0ZMcv
/sIuAFw/SSZe5jBGBm2vuPkfGx/im0rPl53QNfVUdLwVKGLrbyOS7byJP+En
WxrDRbgTq69jcl3dXThyaz7/vqu03NLT63To5ukH0mQatcD0ybsF8yNZw6QJ
Fe4gCGHAANae0HJ/25WhhqLe2WrDAzZWYQqpKK4L941/AJMjkhmD4poV/wy4
PU776DKqU08OhsHOMHCpx5FpTwrm+9T9BDhHcc1JQyOkbbUE6sUnOJyMehP4
E8QWGX1BJ3Ci36v1SdvWyhuxS8LLzTjkaypDdxOznd++NIcwzZH63Z62azv8
a7TJqqiYiMIX3SxJToK7Ga6CvSA3Nlvbeghh4h8tFseSWb+pJu/YQYAn71AF
x6VGb0JVIyprPkpZhU9iKfjW4JneS9vNG7y/PXYXhCQOt6Q0v1teZeU+gNqb
iPyQXqO2QYAK4+XtjOJ5ozMU1ntBjFeAyc4417axI8PKKdhUKVvPx7snBaBH
4YNvqEPsN+9tNF/tgbK/qOqPEM5oVKdP39bGR0V3x4JXBY8fR40s4SWR+XLa
64I7mTVoppcAbu0iB4V96G6J5r9E/PYCRABZzWYF90CLGdVW6XO4eJuaFbKC
JHfVoz0VKEF7dcr0FMsX4jrhbCxj1Igs5MsO3eDlnRYhGkMJ9HiqLSxpQiCG
rXxucZ9PGxK4DhyP5SkMJmFfv9c0Be9CDsNh3dxHRphOJHZAgZmU9XW7LsEL
o5pWGx14hAC2cHJONgUFhgDU/UegWjJtL5KD9Fob523FvhHokx8e6X4qo+sr
/rdNipFXYyJf6Foq2u2hs/X9hnmzf1bxkm/g7T5MkRUrtjnYGSvFbRmASjwl
GVouQ0rNmQAfqV6SoPMFDywy3ivZxr48yRJQ9yON79hN2wvdy8HaxhyiSEWV
hpbrreKghRHB4GAfA/DSgI64VCNPT0M4S1qMihjBmKGufn+OMnYgpYGSm4Pr
wg8qIxBW67lOoaX+yDkJ3SPWOtaUOV9PAu3xoaTET7phwM6ff9GBhiNSmrHL
myUGjc7P+15Ivqrd1aRifNt8RVVtNHeEPHQ2dW79IC3VubNqSJrCKEBRhMeB
Op0nqu6CFJBI1Q8klKh2GZ7c0xfaE0KxwPGof+zR10LwrXJi+vSapCvfomRL
i4rSO1WML7KmkbtDzl06Odh9iymCcpAYGwuu8nK0oQLLw+OegfqhDFSmPO5f
wvfsn9aibS2NJV5h81uXMfFcc+ZvLvH2k8sAy66qoMLN2z6UMT0bT2wwMYYf
i/5Fzxalv0XMJTulAxHEVTXPq/M+tFaFoKvYiK6SkRP15RebXosdVQs9/Y1Y
K2Ak3pHHrERmW1Cmj0kE1qbjXq1LLJ9KEHmCef8iiHb4neSBGi7ew6Ko4xy4
J9u4GWM8kH1AclF3deusNl0HnLULGwqp0Af3mifsSbnF1cTIPngJ4RfoPNzd
MdlCBl3q/a7FLmuSWwp5k3qutKG6YbsiZuzjUAy70YhHwEC/U5Ow0W7QRB1R
j6QcBfxqLnQrka1AQEG0qWT3ZSwjzIoc+dqKz9topiunzhfy95zP1b0ygfdl
z0J1JDSk7JjdkC4mFWFek+9HjwAU9OW+8wJcT5P5kCs0372O+vzKxn+v7rNS
ZY2h16N3ZcfqSU5ahRWRnhEVrX1gT7F7rH15c5qS1j8Fg+5GycqeWpSlSwre
F5QiUO0LXsqFBurBm0R1iih2ZyXExF+UmpABWMJs0tfRr/fVn5cdkTOMXq2+
WO4MidFTCRh8nhESL1p5eETlFMDcEdZPWew+J6dmRLGGazya8BqrutLxjGdp
grR5/sbj3r8KDJ6JviPKxLdWkDd7X9T4zmsTPLE7t1kK0W/ZHq7XtjNwksfh
NhpTvPjFMgLg02Qccm0FViXfe1mcuiaEXanLWBMZvzisv2Tq5+klS9O4PrID
Xq4Ew5lScOS/18uGzL3Lr36DobmbvyksCh9dl94sTJ2pKvyWWkkowbfdxNd9
bHJz0fKPrpmD4+U+G31+QSjdz3OjsqHExTZrKLeRGJLtwkkz8o6nnEVoRTGR
Am8uDl2YT9lm+b3C/8l3x8aRu7uM/gryBQ24v5VSLsQpMH+Fbese2EEQVcrF
yb1vKgp0dYQ5tTygmOxyfUsOC5kdNWsdPIYfA0Zdld/obe2mGq5xTEkLUfNp
rtqNekY5MEdJtLWKdReYmBIJiANBmyUhC/H1Do32cFXCdNOeNqvDdjDjNWbY
arPHOygC3c80o2C5QHU6pexntJ5dQKsbqQrxW6wbuhFAmlv97ao4AduIsfvR
qlZaE86P/a5cSGDNzzexxwkJ+09EzZNClJYivWA3sN12Md3SYCHnSw0GYFl2
57dkIkw1j2Z7k8xWTge/f0PtP37javoC6UOlWB6Yt1DNxo4nSvyeXPF49Rmc
94LxRR3IFZc54/n133cOpBendkEQNtIlX10jMpkBaU1yctB/JOAJIEC/4D0s
llb/3Bkx6Zj3F+r1l52LQ8kHvx9PVkl81XbcMyTWtNY8EAUugLZrIdrMk2/a
NPSUkSpHTU1ucDgRInzYQg3FcvmnYOoQKYGLtsaXOie6SvGN1/77o0F2glu1
pk431TRI69FsiWObrh2p+NAG08k47ueF2BcbRqq8dG++HwBD4s8sGtz4Ac/l
ZBILB+AJGawKAVRrDuXKJyRPcvjwyvINEVc9Zdry2AaOIiBNdpefLRGnsWDB
a/mJdlkamsiPohv4T90/O3HEWPXGkFQRDazGn69NkZCPl3KSVtK7ea4GSqQw
i3+ImPEr+p+E+7lJeWXkw9zo/VeGkT7u7mulzdbzLwWPVRF8s/gAVmgKwKAo
zt4xCw5QMxOZp9kMQgwQIhlVz084SJ3xYCwoktYLK2H6Xtl83q1B6t3Gv+/Q
DDxOv98ZO6IACNgRupDGLNWFzNERmSFH8J5bKqF0zE0t6wts95TKL36hUKTG
224NE8eq6ptiC92T/Hx91FHZewjK0SuGjQn6XPfVvK8yGqLS3eFmBvI+zh8y
TU1K+OjjoKdeYWwlvqNOvBPQe4kiR1EgBcw71YqpQPnHrJeRjM0VYfdK+mzW
6xkLVQiJvlo1bdrCTQCSA8JMcL9WohxpWusvJUIsNN5rUwsXHR1rruwO3fDc
kFPmWnZvyaCpzVCm4d4a++btHGKKVLb6+Y6b71Whq+9I067nYMOfb2DCPXPi
9HT4O445y7kV1lkKiCq466K3v5HC62nZGD5kKaKY2qhL2/UcGf3gNS/QdGRt
N0MZTt0mmtyMjewldtpyouFW9d8YRZ7LLY7YEG1VxInsTSyCXDP8Ir1JVuIC
WlDQiAJUs+Fg+jZ4ufoucdmM7ldZ1Vh9aPyeoDJJ6VbBLVM/3lqINWHnMEvD
Oy0DUcD+/pFRkhTBWRqiO5opovWxnv4GqrA0bkqTc0ZtXRIHy/QzqHZc+F/1
C9Gmvt/tpEyRO4M6h7Eg9lWi6/E1xsDFqUKZI7h4w2HE932ybeTNcVOWDRT9
4hSI67uLWOLGcpDN363qLTOeqyssBRpb7KZs/Ar4eAp29mAS/oqgbpNR+76B
X1QSDifVKK36QjmPNmUo65/N2z4JsUgLGCOv7Wcf5Lfzj2CoxHHLG60nulaV
6JJtWi9xvDjBoQmo1ff0A8liQF08mYbsLQhAu+Eonr5oTFj5UUaxiNzyMIux
38Cs8awjqn5WbyPh/VERXwDl1NSZYmSfsNQENecw6NJ0iDKVZAPEaZc7IKT1
JCrf4CT1gWKBpLgRvIdDbcXihxk5WsbZ2Q78FqPh2hRDr2mTL+vWAkrNuOSl
mnhjsm9zStIBBF0IjsSVyCbrAjcUOa47EkU2PQR5JYeBfMcHjaRWgUA4bZYi
qG4daEAIhRutrxpF/rmZWiEhlCj9tzGN4ygHbEFCL9mRu+1xHKcLj48p5UVL
9A+/xLYXN34hTmuxDcBCUawRNYd0A7ALUgmreJKkoKp6uknh65PX4GJhBqHS
dxIOQTSYW+QKDaEmYNPOxWeAdYyqbcIeLNBs16bn3bBAJ5uTVkDZUBE4dJfG
8Wds8hXxhbEv+6OVRToZ5bgu3H2Ao7XnEiFgw/pZZnjZGN0x0HMzb8QpNc9S
bzlGcelPaQqN16FahhPkt7YVFvKueDNgN/EIH6STdp70oEFCdW1uuOR+cdZg
5HN+HoJqyTY4BblojjWGKvUAbgTAkjyO+jEZ8MPpb8Aij1PjDnAnTmli+Ouz
uKt9xCXoIrGpUY9guuRgzQlL5tYaPqDQ2wptJrfxKbCZ7MR8OITr6eQQ6B5O
cAV0fdn7gy056Xscmu+cH4IabKzLC6Axle2uP5ySaZLcuxzwfCTFwSK/rYe7
nPxHbr8tIhx3vNvu91JGsMo/rx5bBbVD90+5G8dlZT7eo4yA4Gl7V4lnDKw8
qjc1qp56RVpLrO/9uR3vt85uaqNVa2CZzAgxgQeeDS+URBjGA9Q9/yQ9MBl7
i7EGpGtlTDc4Cu+2LUJNZOsOr6pcURE+NqRVlC53hsoy/BNHXMYuaXsNPqSp
9H9uHyqtGy7UoYefbk52/uneMzZoVxsUZBSs58EEiBFMntnMXNREu21Vxgq8
0hXP3TyKMo+CV3Ve8p3cDhTt5g5K+JYIEGSSzed2nKe8KSpYdAMW0/RPSjWl
P+Kk4YGy8NqMG9ewq1ZVaPD3zisXQ+dsky5UAsMf5cUGRASR8fjjRm/twYLt
iRRq85FXCV5HzGAl2mHVBYWZIqMcWOBSI89V9h7FUs9FOnFahe+tNCS2lKMK
y75oZf20vyw5ulNSPXkNtNNmOFeM5A2EmpI+c/MZvANWChtQkeitPhVsuQrs
8YT73eD6fs2tl1VjjiynlzVbgnLOyda27WOBic237mdnpchtd0oWfYjSqhAK
T9xgNgoAhUOPybcjV/F+J+EtW1kvZ+Jk1ufsbOcoWxO5QBf7Ww1SzAadgnal
byl6BBO8K+uyvzlVME9AqzG5CD3Flz8u2S1TQyIapzR0f9uwB98gNZabhCHc
vLSY+ruij1hkubysgi+jTtRPH/Yq6vrS+wgziZmiCKeap2pCjUn0I7D3XGSR
TPy0u15y6kxjWJ2AXhArUFv5FfjGBVM8Itgc+sESFMKh3/PRwPLOjQ4LL14X
B11M2q7lFVYJc6rdIPN7BdysovtHfTCt0Z+qijoxHJTOOBrAiBjzRg5xXrzJ
9j1SdgR/sOi/Gb1ZiFB+jT/oIth9ID9sCPTN76z29fHng2JSADozoa5saPZx
5x7z3JfqjbVUYfd3wVE/h8w5IBdsWS99ujmEUXw86EefXKFIbX9+TX7YNgd8
3/rvL9wzWMQcX5PXl58aGXOBZ4kd5Rnuv0XBiv9QrLBJNCCJVfczYsf9PO5N
CLhNn9xlDtEp+14vRLnmG3LQEhyz0I5lPrzjmIImTQBdG4jZPJ3omIfO2d/9
KS/7mDbX3AqM0wr3ECh4RaWRhXpw3EYU9nFJ+dZRQy9DTsOrol7Vmt0718M0
UJEQhSawZaig3V9q01poMIfxToTjDWHs6igTMYxzDJjD4xQDx0hNguUepPve
491/G8gugIjz4Cgj2JfSBAM2llt0LF8n//vC0i8jcitozFSx0dqdHbNp0Pnt
gOAC6zMWpqxcnBcWi9OdxC7xZ8eqwJRY43H02OcJpwHcHoTvKVwStOxPS3G6
wrv1Ilsh26CVKMEG0EdLMpehZK0xBqjgVUAQru9ryYBTTgi7UNgp2VNXPBtv
yyT+2QiHXHUOw3PjPj4sN/s5PpRC/caYN3Po81qrNYAjp98LbajHFzIp0o41
NsVAhuhp4aKCuW6VE/H5S8107AkNj8D/7bXzuYsLJRrzHqry2FeDX8ZZa4lq
ZSq4LnsYPpbaW437dzx8wI3V7N4JxekdKiowpKmb7YEiPVdXBbRRFdtcIuAP
Lr2yf/lQDuppKXb+J8OYprpN8j6UC5l5U2U7TEi8pnNVKShsP19gAFn31+QI
FxfUCu80oq9siRSwoWgjGLMSSovZgtbJNayPZScx5Ge6S7oG4cjHuBsx7DmY
tpfxepCxhm6RmxJqeg0NRbnAVfM8kfXfhnp81uOBNVFuPcMDwfMVj4eVqBoY
rO1XGACgWyY5Je5heZkJR+mIiHSs8EPM2RVF/SuWcnhJj6gJzOSRY4qJXCqv
vU02TkxsmolJcULGvH2kl7jCLtPs724P3j6rkVwkWCeEfZilFFR3SL15vAhu
g4XW7RMxLYkZsJJN61ibQCk6DWq8o+ZpQm/Obhk9o2JsVQj0xEdkc7YQnhaw
O8ijEGtaluYYnuAm2OXWl36TvMgjHAO4NYUNr6BwtLPIEq4nnzLWbP44dxjy
vmoJUhjwQJxpOsNEv8PwNdarLU5x2jyyEAQsGH0KfF2rqz4g6fyMDW777UnX
OfPkDf/EJYlcyBFWfaAtaZZRV8+ujVT/OnsfXVo8SGtjI6RxQIOsQVE8jYF3
lRK/4rceZL0Ch5Mb9aRsLH+NrJA76Qz95aWIyJG7R54JMRyFEhzLormlEpYv
7rGMaN2FmSAXX+GrxSQyQv78o5mMToInHTkcgjM+JEuv9VFFBG2mfdVzmb8O
qVnbrVpnETpVfKVEaclrdqP7nFOmzR3UWlqUNZIyY44DVLJnWS5tb2mH0eAT
BkT1xG4Crrsyz67FY/GhBoxQo2jW/fJHJ9Sjud6wXw3z78Wu8zBgLM2iB/t1
O02TIZQPL5StW72Uz6+4EDW9fq4Enm3TYIrxZSNUffZDF3JcxQKOjqtzslDs
P88p3YzozP22GaI1J8o0wm+efPfN5CVZP+92Cs6h8aSJZhxraOCdMGrYqKy/
OhgKYt4tTvAYr0EnyMFVrJtKWkUSgHHHpeoPv9al9u1JwAErKhSCpM/ZH2PF
BCJXc3TOoGjIU1Bhm8+RusjaP9EaWSSLRRx2afzBjb38/o0fFWnewd/7Lz5i
6IGg3HhrrpfhLInMQXWYouEioNltklhtap8S6g290uv+DqPehu0XkonvB+qs
DpxtdxedkWpHHGx6O3dNB1eshH11gH4u0YopMh29CjCdlDuuIBfWfWX3d2y7
wZ8pIbEMUE36bhnBVR10mmntGYU0ix2S/GkkpIT3nZFhu42HTWXo7J/lZhs7
WzsG14EDcSbzJij7KeAk0mGT1XJLbjlc9+5vmT1+6AQbTzHAP0o7grrNotYH
tbqCtqL23ps1Azz9v7cvt8orpRnVZlE8Qvv8sKMfdfDM8QOZCDfv911SKC/e
vwc8s6lkPkPELcvTrQCFUqEiZKGpm+1lLbb9ar15Jqiyi7d51rCuwhFzMGaK
M4T6j/d4V8WCRMud3KDiCuv6AD5KZF33FP1O7FenMieSrqdsJcisETU4Xvo/
dzkC3205jnWxw1aoV6hpaLa1IEDiTdZcE6z/c27GE9GWT4ojELh08OIDpMvd
F4gnyVrxgHvrjc2Q377NNOLQxef/x/vr21UCc103LGwDV0sYuDl7z+itphmX
VId6Q9XB4xBavLGpunc7pq6dg6PKvVTs9g3IPxQd3lJQCuGVzQCeJA4uPHQ6
98Jrp5VrseLKPspeX3m/qoqp2mjliQ/cTpRg9Y2PGQlL2hSDaT3+h9icfCBZ
xabaqmvBJ2IN8O9e4Mz09FL3Dd8FTbI857XuOYCwRGYum058am+khjQM1v97
2Z9EREStu68ohcK/geXsr+D1leP+y6hR0mfhRGJJOiCuZnKm1cx4EUVso8nv
8U2JOEkG7rXIxM8kKx8suTs7IZEhbYzJqxa2SQfpexEFKnzmCSfOOadw4iQV
Dpw7E67b7trViBtotOqPk6ugoyD3GPBznXW4In85Dd5C7sOOOM3W2Gy4JfEs
1x4uDEsrZQCwj0tOErwotUdvbpldtbqHIk5AYP+7YHN5lPN73jy+rwMWsdXC
5TUChaWFJPmr+Q+tCpWVv9J8nQVxGQiKXGZAq5WFhmmcsI3SUmFrcOQ6CPMV
t9oYklnUr9he4M3y85ybodtShkNH/SxUCzDQpsGWAdWZ75ZJHpaJY17x9O3/
gyamjuOIdzKZyaGolelAq94RQcbBu9UwUMANd8zcTfc4KukyEZ2XqGv2tY/N
8CbKAjenYO0XlhJ4zMtyqXSqiRGB8wVzZKa4J2uUhYxjAd9GemCdN9+TESY5
ChLjwBXvDxHzHlOJlW2jHdEKjjq7SGWDW3f/Pr093yf26z91EKspJ8Vng6Zg
Ow8l/YC7VNPvjeKrVlcocrUPlU4GH6qv338jEwKKxtvWvOOzFjjXNCS3bUBv
9KcmA5qHHv3N1l9Rhzk5Cy0Dd17s3QkjDwwDMHjhirgb3mpWab3isklz0q7b
M6UiFlzUyRbkBzGCClK4nyvNx1zNBrD3BxtjcAGD5gY5Pqm09XMYr3QTAd6Z
K8d1985gJlof8JFEoh8qmLT5XtnLJEqpiTke3g0NkoeSx1zz0J6dKdL8f8T+
8j1VXHZbxXAaF7jBlWIL5B2/o7Q6jqpKbAkV3v1fT8oZ/PeO5C0wAccDkWV7
lc8qLChE+KqlxOwCIvMJFhnXvTbbviLxwLIxsAhXx8hFa2Hwf5ZH1zp3m3d3
HSMiHvbpRq9MFiXByLC4edebIaL+iZCCqkMcUQIS6mEz8udBCntdKLDOk4AB
av40763187SKgY1J46EXESwvDiqVW5VFxGUJkUNGziq2v33rk+9Gm7sPlPKM
fB9OTg7hpIBnixD4lv/wtiRENIDITLj53PPm2+Y+5kUSEAedEKw8MAefeqxn
qqMrGR/qKbUQ2SvhaAXwliTnV4qPt8/o3F0RgdIkOsppI5gRkTiG3+opqBI7
2P6exVy8IaDe5jFFiey6JSNGOcIGVlapJ6ryPrGQcDCEI4vTvSHsVcGaX+ZX
eUsq70+pWYy46vMexT30ek6Ep6y6aFjL1Pbpf38cSur+9bq17nxQwD99CBVS
WWxZFEfj7uAJwokeatwG7GrkDgYkeU/GWfWTdZCj3bWjbGXrB6hwKEO7+NtN
0h0eLTWohuEqTa8tfd30EkSc/7sFm1JpROKXAyXpBciKJ6ZU4bQLi+hEFdJc
ZGYyun6ns83SuYNmHK/NKqlKuhaONlgCiszYwDnItUFbEoHu8Nx1qZI6njwr
GbwjP1CwmLTNc5oNnTKXx1NA8m4oe8ES+C5kSzOc9lJEJDLVh34khVsvoKeM
Ia7rdPQJJ/PWVpzQKouQgAA6aF9U9aE9JfRCmtTaH5w8KltGov2f0D11QT6v
qTrPgSniX3Mx1/l8rhrDgG210VpKykmLUPmgMGLh7Vitu1Vos4NE27Ejbwd9
+WdsYorldY8t7j4rv/Nko0DnApb6+LvcmQisRPpVSWRj7JqxoxzxJX/nGt2f
ChUnDTNUAJ6bS0YdDbdsKmEhAXuwpbuaAQ++YjjicwRDYCQOZoITONCyCIwH
h1iR1O4Y7ZBIdoUrHw52RDPS1rbNHarBCUxrQIFNsPZusBItQU2ntD5EOt7d
Rd/GE7Wn6NiRrLNv9gQ5A8ibqDnv/SjxrWuzj8uE70QfCWgxVAv2LzNf1lV/
kyArfjBTJJuYSjRFSZE650d62uOqXXy7iKhu7l4pOJHWr0ga/Ew2mNCpZ6N2
QcFw4puh3jFYeR0NMVvy4DOAB9noRw6iUyATP87S1Pr2VRuKhN2LGUblFyoD
BFOf+VUf+PaoF69TkU9lbfMZCkAHNLjeQFFLhk12VF8HZxsGcyltxM06+wnD
WLE/HgQuztEXRM40YP0g51h2CSY9Z4b/oyEA9spgAj1gw1oxKpHzgPHanNQh
XrMi79Dmd9uiR94oRFZlTr/oClnn6cFhv5KdPqsR5f46GlwTTxeeuD4ZMFc4
HIuTuaPk7jMKrA5YVLkbMG52HD3ZtHUwKdVfXeChAJNF3aLY6XF0d07OzsxD
Uv+qVIaEyBZCrMvRy5RYUlNEKBiGstW2ETAqKy82E3MVR7rnEDFjFFigW8bf
554mSGJ5/Ig7kLBeaqj3FRzG/NkBQvZbLFCBP6Z8S/Krgl6DDNrTDlGGeCle
28mmTYiRs2C3WCy3VWPKkmf08JCpkyC6YpA8ROy1sARz9mXJx9UlGo9HIEB9
jVX3oTLKqH+AmTslbpTPL78Cp5Q8r7E90vCZNcEp9+gsg6nr29ySLc6gWAFw
/BtKLRTB6tKe5QfX3ZCDz6vDv009VU+1q25GwDX4dfWIfaRKN09yB1fFWCcp
mB39g4S9bbA+ulmgK6S+tzSAEgMSmhDokYDIccjrx5Fy3lJ5N1PuH26CXITc
q6gU9UhjuN7tEHE9Z9QFuaAMbknz4HfXmqcku65U91suyXIv66cz5Adn82i7
NLvreOWlCVSqixp53+XP4a04lAc90NGfbPO8IYKzkB2EGk+q4hM8qjVxXXlh
TD2TNP4nY0O0ICED/+JRa0pREZiyqcVvsd8pTbrYPRfeeB5bt2H1v+dbndWg
y2EYi0bOVs63NFSdx42IyFCQOEYyHV5+CNthyf8tSw8y3b9GKvylj20ildMz
0qGKn08AwScqy6n41XtDsywgglVZ6qLkVx99tmjssjpDTpMwobUMcG/QCOFY
hs8ByW+bI4YRbgv7omaRu+6047H0ljX6TdT1yPB/zeJLqFj3Mvd5L3Iy/BOJ
IKs13UxIhVoxey7NcBQkNBZ8Laf5S9oQI04ITReFB+H+0HZE7JbRimzvh1yN
xudxWT8nZYgbSFe2W6b8SGg1p0rxySO/4ZQtGmoRgAcyTBnq9Fkk/Our1FlV
y9K6gGLoOMiGdChh/4L193iTKeedIlOyNcJP7LlKNp93gxmZ/SfIvVtsTcZ9
osS2dNmxS29AtDpLUe+wi0lqLeApTQ1TNDVQ4KtBXHz/rhYk0zA/bfjo4b6H
pkS0+Fs7aojbGaOAbB1pqglxeqJ7XKcVDqgQTYLaEasg/qzfx56ady8yf5Cz
Jm6T0qp7QRLYmsRxLz5uOk5BCn7EYlxAvcN0z9t+wgwG/mY1sac2X0jCdcgr
+RjYut7kji4Mf44wBxi3JaT4gra/qzskl3WzDa1qc5U5m3LAqOtfH88kpcX5
abwufGper9kgQs/oPOaeDRHFpOj3Or5oznOgUtQMVLlmCk2TAbHOxMyQrLJM
s81+qGXMkHo1rl/y+iu5dEPmV0oVp4UUBNimShPUW9ES/Y2dKdgVG0m3m+sH
6SB36w+/Q9DmufJKw1TmcuwoRHI3dgPlF1d54zxCUJ78kLvFt6CSj6lMmzpy
pYRh35T5znvPeP0v7+OgjuMO9qBmIQ8nthi2YocGkcaS45cXSAr1ktLDx93d
JXPWmziFkLui65ukUYKtq3qnHUP+yIWwxR2MNY0Q11G+pJ3nOONZf8F97hKt
KCXRKdf1rTbBWQ2+Ew0DrqNwio1tSvFaGHkalWX8XCkosCNwIzIjA7f/BtxX
FFTkSO4A5pYoJuLEf8ZkwoEEBxx6KTDw5ZQxRpBoWXgnPZrqN5cBCtJ9Y6Qn
vhdLvV6XtZVjA2DQA5+RZgZLQNa1OJg7zPuIh+GMifHTQN+7lMU30rcNNgCC
vVtBlqzupr5YLaZO5je0f0KZwPcxV5PZzsQcyJwxpb1u48JfKu7xPepBUcI1
t8WdN+EobmRBpwWzr/Sxt75VaT7VTnEHGJIpyAyFCt6HxmvVu91DYVfpwXuY
GO8QkiZq71du0fLkO9RmB/x7tQMQgPJE0uUsDahtK20WwgmDK1AOu/aQKYtp
v5TkFtN88ORsOU6lpxufVDc8NTOKItql1Y9qp0BqXkYOBWP81GstwieWGC+O
etpcBoL2NQypRQsJuQMca2mFlsCzrg2SABfPvxTDjrnapBo4EMLWk9Hxwh/Z
csc6ZwqA1BdRrqVtHZt7sBnCBRSNMC9PwmQTLIWTw1xSc/xhD6dJp9qHX6lq
86TYNysWFzkUZ0GcifN1+4y2uKrtEa/aQZ75Ga8IzM/v044Jjxpgv1dhLPrq
/BUdUB/ugVgPhq0ilxTtOTPmqctTycYwVnzvoYQDK12jKRFW5kq6kkWEHFOE
TtG6CrUaTEe1+KUXoM85N1jvCxBSbUs8pwNJMWi+IiHTCieHi+k2ebx+GOgC
3iUYCtNsyuDlUKwdg4+5uXlgQeHxiu0UU/cvR5mpMX13blntq5SIQ/9F4C6s
4B/n31KvYyIKWaVO70M5VNAmkfe7KkeY4/oHb2BDeCwRSViU/jD1iXVCngKw
g4Mkte1ZtzDDcjqWasuQ2CLtjpqcXdtNyaAqWKLJ9gofEE+v0PVDts0InP6G
gF5yrniOgxZK2IkwXEX3avnrkD3Ot42sni6vRSs92SR8xJEO2DdcsvBtD7BI
pLPFx0zRtvAUDLmvvkMUGkDWje1MVvfCmdcD+yRJ6/BwjECQjEE53rdAfEDR
T4zcHwnM4KZsTA3CYs/VEnse+bAQOybV5oxrD70FH5lZs64rE86/r/yahkfu
F4cSp+iOI8V7LfRHdTqOGAoUBa7DilHXsbf3FSsdn6KVaFCAvav8Le5UyycH
pFBq03nRDNbV/PM0fponlY1XH1jfW5SYjTgG8TJmNWkwdkP03GfzlFezb9J5
td3kp6/BUdW3+bPzWQg7IuSymtJ9VIRfvJAxrYecKpqwh1O2R4O7x64+gR11
VhgJBAO48sKT+o0lDe+xI8WopXeE1x1SG2pdayNrpp9DUKZaKTffkZCa22YQ
Zd1ReKwrHLocyedoe7LhpOZ7yxJ3EJXUl3DjWCaYTiVk6oYeLqHgJfp5xAth
YnH8MDRaIOJzm9mtnxbN5ry2JxJczJVhI6wvVD+sAUX1ipM6xLylDd6rUdwe
8Am44mknvD6uRr4+4XuCe3Mm5Y12a4OKntXuMG9e2PfvxUjzKKTO+a1UtjfA
BsgNGWO1SgVey9lCwqao8pzFTCU8bCTdnM1iJWL3+VfMkkQU4Jtp+tA+kw38
Rbwz8dca1oN/R9NXqoVvjVtbzyR/P8/4xS6ypy0F1mcM3hMBpEVbaSxgOvnU
XxEJfmDakvhN4HIeXpI7DWzYxgfiEM3wvZ4temsbenQewXjF2D3hVf4HU7BH
8gztZWYZYQ78h2WY2AQ9vVIA9Dr91iNv1ImxtOMWLlxPoLO2jiR3yZa11frH
O67NS9/vMmiNJqQHTM5sCPIjdc95iu5uetl/AYl8X0xjGaeOxTy4Ix6EYwoP
PPJFFXtMVh9s0LM+3d2Nl5ye4tE/fec2nmaP+XMJjC3yqFcyHPx40wIDGUV2
DA4E9y9quIChO673IUogLQCGDyw0KwvNVfD6nzKjn72NQUOPEuhimQhNOohj
6JwjnDifLdWdqscpI0RNri20ZOjUNEaRAxFbu1db/nQJhVbxdUdr8ubEOAwj
bCBhbbdsbnDgUnFJlpxl3rRotap5AHfm+HJ9pfOPd9J0f/fr+eD8jKKI6Xkv
+2OpWBo6oqFaRXV4l4+yknHvkBkRqKDj8FtKXGjz2qIhZL+XxWD7DwUhJQhu
pGie4PQAXqO6HVA6BepteoUkdaDJg4bo++QA5OHHh+KO0/2h2zGIv2kxUMUX
9a+He49mOXIwuMMIAXQW3WeM0v8fKrKS21R1KjY8GqqZkGdpF1RqL44V98sM
gyNKaWte8AuT1GM5g7F9h0gm9GNmkK1Ucrxx0qHC6Fp/b9zBmpHKdF3uHO7z
dme7BPNs7usKDe3vJWrcWI8Kv48bXXVseXTXZyQlHq4OIlYV1okxDlGW/CEN
9B5wEDYnjM4jMiyRhln/+oeuA0c6lMZxdhyCqH93uJZxQPCr2sg2aKyqAKfc
XBPcJKFjxjJc6gY+/tL/BAEVqckcO1p7h+ps55D6+6NjHru3BL+BkRh52ez4
hA0Sg6I4Fu44ctzETaFZ8VaAz/6AseoKSgXqORFWjzVnaQFfwctgrjjV5fQg
cvl18z4d97Ce4FE1zG+NlWdepz6wiKo4zki3KC6FiWqay7QVGsXlYW7O0kb6
+9zaFJYVZjuhVTRegrrP+Hew7mp1SJCl/DDwIoBu4tfivgQKRYOSnf0EZzvl
ikQxCCl+y/rLjGePkTxh1G2hodQE8e2qIE0gDkd5zfPW51JHrYcmoCbHKGss
H4zgNawgyIyqmGKxSF2EVMS0/uTvOsTB6dlKm80GHHg3l3CtYp8fZYAoPsTY
53bEn2w6jck4Tw2IezUQfMAUfe+sosqqfdjUY5lLq6IuXpd+MGlM62twpN6H
/faK7M0sJMGW7JVYDbgguJfp8tTXWjTF1kcqWi8XrGlPup6wxo4P+9baIP4Q
8Ck+ryWNUq5zgJdTF53OIEsnK/Le6fuIjpwCsVpwHxQQ4nTNkG1vYKTCxzjZ
0OrxF1eu4VYs1My5juUHTkaTL9h67SSt6pyFuOn9lGMZH5cz2YOk9Aw96m5K
FXLn8Z7E5E2liFkHfGbcZyIvaIKlClKJuA3BpU7cjvLxZmWWpmP5NLHNLE4Z
TfaVC7oT0MrsdAVW7+wn/aXFf32i1Ji6eWl1iGHHzcfqyRl4bMVu0L2Pzh1q
r27z38Gts9KQvRT1m66BpA6C5VkYDqtnP2dyJbbEegxd7YLl+ggDhBFcoYpR
XFFCb3ls26qybs4mA7Izp004q+4B6oMR8+zRJjSp5h3WP0wJqE4fidlj4qLS
9OXmROlct4cpFdy/SDq8+IyVNN9GvUVsge3XOlrMU+ZTQEskXE/re45ZJESN
bIZOnJW4cxtaeQkUlP0V6V4GeCHTarumYKzB4KIsTPn5MCKlBjFd1Zm1xJXV
u8Ld587bwuYVYECqpwJBmP0n/gz9NcXTgzTaFnBfdO0iQUgkOIhPU5gTrPfS
LJxxbPCxBLymcXbVu4CAjxvT9RbWieguxdtHNUOgdE8U2gFQVs91Hp1XRBfM
E2SAtJJ568BmjhNR8z02HA1QIwV87yth3nCfSPfs2oFIX5E7xNCACk4s1ozb
9KQo4yALsYvFBlC8YrWESwP7cEhyIhOLy6uS6AkjG/WRlVExM/y0R+sLqOlH
rVE6+45AO9iRurqS1ZEdI8SNZ0Mejtal7Wc+ojxbQ/WlXDZf9E4AI5+STWKR
F4yrTZGYNnEUAR07RA79Ib8bnVKPf7A+knAQtFU+FvEXAGaVff5siOkNfTLF
pCstmVhx7GY67o8hdgLA7Dyg+6vfl+NWkozXGPPGFCC4csZ24pCSU4REUL1z
dxskkQ6+2jh55df1+aLhGY9GGolvKT8lq39zXElawb/6H9Apn6lBHjyu1efF
hrUE5c+zkIbhwMhyUkZr9NkxcbqAm82SS6cgDNWLlGzl7m5vx12i9TEwvnaO
7MWQkPkl3sdW4Wy1hSCvy6WxtbbQ5+Nvvih3O3JBPjvsfgR+gQCr78xODNO9
IbAgwchBIrKbCw0yHLfGW73gPiFoz8Jdk75fcwctut/qpKKb4LkUlbtIpqtD
d8i1nXLouUt1BHo2cj01hxguDQY9Jc0STMLqwQKIiGrouNHjzHjyUo7tS+22
4NQ0GSP1T8n5cMLfkyRH55CZVoPZmQhyRr2s4HMoSANMNu5hXQ1QP2J042f8
IL8/fEQfYWAU/UznTt05O2kYBn9A7v+OVu7hsVJoKtex0htYPbNA+t9QvJlR
XgZPKX+g1fTLlNmsfCOlkKDi7nq77xjOstROKNcMGSOKfgwuNxFdh4S04yYa
w2HrWEVr3RwupX75eLtHkyi5oMN+piSN+HH9lMnnNUrLyWjj/NCh+8N7D9Rw
rnACFFUiZjTeTz6n8CZwadbwj9+/GeBGhgwj14898/U8aUtEsaj7Lj8bpcai
pUZpsHnS709/JS2tfou5OhKBD8QQqk06baUOJWPBf8WhhIMil+FIYFKL6Lmq
80I2PqUZJGagQUs7nU3CozyGATAeBfjnemnqf92MSeSk5BYQHiuDElvqJ/fo
8gACjU71kZODctppIW5/2FawG7T1T3cVwlwtLe/y02KejMd1O2przY7FHw1Z
M1htld3icLrXn49PXt/JlSYWtNfkoQWGyUsz7gPHe0uOjJxkczX181s6hqSd
93CBPvkjZsgXj7HxxsgRZb+tYa9cBmf3vagQEJvlKRpsAXRYNgemXcC8+6gx
KkFmLOk78n/pjXs8XCMFtcznfoZiqVWUUYOJ/gKC5txOcHeiR80nGKZpRU4Z
Sg2MDNbpI03hlofijUqc4MmzOehN+u1DQ6k9nNWQpf2yMaamFY8uOWeD4N1F
T9c3nFbuiHaBni0tbaES9ltHlgR/xyoEsz8lN6Tw3aLwrBp/Ol3KAxUDaFP7
2WDE1smuuk15oW4K9d4mLRDSV12tsto1keVcOPjqmqEgFndktxaII9Hla0cP
LY6vgp/X+T9aYTIUGYp+zWTmkbG/HGiA/S2jNFSmQ4xTIGAAFchayJARyK1i
6Rb8b/nRk8dXa6GCBjIgRY8Xol2i+hwXnYpFyKzHLgOOMM5oesXaQPzZSBHU
CzkOf2LB7EeSKy5xp5DgizkjuzV6xvXntp5J64yBfaVeCbJOajFHFVIMQXNQ
CM8HD84zQtz7GIe57ocLIxaUBjbf2f9xUdVQFNm9TvKwDddtD60GBVQ7wAje
9KM38rZ+gRIIf0Lj0anDi+tNFw9zykTEZHXVaieq1w3J5ap15z+qMMPbEXN7
T0jiol4RpLRVwh6IqGnOXVoquqcQCN4/Yzkjf00p0FxRJ5Vf2QKhNh1LY8Cu
syel5XJKmsfrE5ooEHgPLfpt3TGnwQP2tXsWPzhcPVTqlHp1ktmUJmpzZV++
NdQ2ao8v9oXSPZs6f0YS76tgR6FlioMgmopHDqzo1muOlYVb97RLMNDwHpXZ
YwxHQIuCegAzxRi5X7d2kUC8Ka4VnVmvUI0LQXZOwFHZ6QPotMtLbeCnQsAz
cB1Mc8eqMO8V+rPQ3JIpRP/gwIby3qL8lrrgC05Sf/FhD5vs4uNJe3co5/M4
N9s9Is/AZaA+l0YYLzfRTDPaa9JHxj8CJSp1+mnZQtlMmYoNE4xVzkAij+/b
QpYntmxXkbDYF8a6i7Om/u0EqFgQIJ8VG8WNHfwgf0kty/mNAmpuYIkKD6yO
OuezMHbvSWT5SemMIkrCDxcwmwiOCp6TTj64xKzD52gfgUcaAWCU74O1S1bB
g1rpx0tlqLlAzRVMFAFuUVY48ZMMRM1r7UAhaE77rQlzczD8MlDPy2cw6Kn/
GqmeRCHEwPaZgjWYUTOAXIEKACjdtxM5cpeudkz43FG5qQemjNSShz04MKoU
4DHZe8Nxn9NMnR7Bt9FquBPucqC9BYF10naGJ3OJDGXeIoNZ27RxDnr52LAt
TDQuUpf2HCLVv1yGjoK1dQdHXsedTUlUld6/7qYH3eGV+Zzo0+7XvTUT3ki1
xUSLi2yCdRESaScXu2dUin7msmDwV/KF9lDdUdpEYzkAgtWrS1xrN9shOowG
5rr1bkVEaZvje5VMvW02iRC9FPsDJOutY5ixyk0JYwVJJQr24fehj4T2G5gS
W7MtctGfDjPR3kU6uRW3p/yACjm6jY6G4V4t8q09hBxDNROpMY5TPTkXkBJg
L0B8T/BVask56mbSvGztyPFZeCzzj2+l5ErCAfPb5BxhDlRnaPj/lTgEA1UZ
YzcCYOSeSgNgUSRAzprGW3XOdsIUdh/tjOgD941Q+fDCQgbO4FWQrrfKbINA
YDOLfi9ELYPZQC/mv6XbTMszevo00kzWn7IbgCuk5lVV5o7qhhczx7jpOEEG
nIZZwuEFw2ef/7rJDkjwieemGYTe1lJyK4lysReDykeWZkWHMJZNgLBbzULX
DLtKybmu/CNcKfTcFHIY5qocLRG2ZVcn2Fa3FGJgjYg1jHVuYZM360YSwR6k
DAoJ8iMOj0vylCrLFKqHL4aT0r2AS8hoaxCmA7uEXjHp2f0v8cZ+JSSek3LD
Jg9RjweChTrfA7Xuu6WW7WjECDaEGeouG7WP2qTnKQTchoZdhZkk56aAw4ku
mua78b57G8ejpFbTITgGxsPQvFyv13lLqP+exnGw2hUKkoG/ZRJ3parHxzz1
lCUFytxNK/0Hc+3+IgyHfHUSUjal+oRPyvYVbKfPXE0IW1K+/L6e13VIbwtl
r2xQ6QnyEJxmXAf6kY+C+kUNrXUn95yLTcEukKq5mwF9tOxP9fq6hdbvAUJk
sd60xYtak0Ot3Fo46iA+ycj0SFGhjvGgW8v03Z4B9UGZm+v0qWzZZK0hYAo4
fkHf3AkioApYf4RJ5u7bx0FQXhTJcWsSu7ffzmJfbM1Q+TzLqbWFQ4Lw72QN
PMN7IZtYUZC5sDf5Eq9iimIWG7QgYUPK56pvXt6Lino+RLFrZrRCQ5m//RVp
l+rdJBXK8Pt7LjEfk2OwwkSq7SI2qL+QttY/Y+GiWagcoSdr+0jOINdP4ckU
AQrSqA80G7bLGaY9C8T1KpoXhyt2IvQATNz6dCnwZenAHu9YsAOT5x4127iy
B4559AiN9ZTExW5nXmwEV5UcEehMbUuxU+8vxkM+lmLo7Ik3UStPMoGe/55D
VElbWvBP9dBBebSvXoLGwVLX1CCAHrX0384mJXUszX3iexrKJ+XT/KBXwgD8
nJ/qW6+XMDMu2mMt2eHtJhnupO81tX/I5YrhBZuru/idcKP3G92jZhA67enS
LqQZSUwbDLH4Lpv4R+pRV3oEihU46cmIj2QCHihvLiC/XryHv8kn2ovw1/xT
W57g/hJdj072AUOCcvesjVJQncIhPJFb2cYtxjFps2CF/aj2IS6I+o/zUjAv
TEktpYNICYjjikyyZVHYqwiz9x31Tv/8V9OIVOc07hdo2a8L39XTmece2ZrR
OhoLp5zp8Nx7IENo40lZ17KnnjJ9NGu6SFwCLO5KTCvIlxRU91ARgbMXYRAu
CHRYWxXIVOaRsrN6nXJrJ2N5RL1sVvxkCKe7YBvFQfnk2g+g8WtIWhd309r5
UuqeQch/dULDLtQlUekewbbbbF129WAGuNqPPcoIc6pjou6UNPoObDboxXMM
MDTePja6YHhOYdO/QgME43oEoJHEZCgkeSZvav+Dor+tyD0BrYzXMjGfePTk
LEVQxD91tnikavsr2TdbD6yEs3N4oOS6x8M59Y7wkHnS4WE3lXjDeKHdYV1m
Om3NZtIHkUs5rDMvAqZ5KxaHIpDdxfOzsnwufKyb9ka4H8pC1ylB0BQDeYmq
dXpA9EcnkIrsyFg4jfjKeBjbGJGYTqnf47HokL+wCy+E1SHjmYmv+FWslRgs
SxQbl+I/f2RGeziiP2qmmvCPssNa4YWrv/+uHymPHA/5sSUDnm5j8YsaifrL
FS5CjYd/dl4JmY18ANxmHQB98yFH8jYoC4M8oqjEEZTzR+vw7G9yE/EDoDDK
OlO30iWycij08p/C2x1d5HIDhMBDBCd1ns0SoQsT8sv2nNZA/VIRTUnEmn2v
8ZZlwVof45+FXhI+eujGJwd0zWYPh0eg8riCTyahLAMPRZOOrhQVyVBoUhvv
fkTcX03fAN59T1Lzv6b159M+mvdFIOU8T6bWhIkmiNuHNEZXplkTL54CpY/E
pTdPOXO30TFTLCqisQ2BcIWlJlvQBNQ8Q1JN6qtm/ugaFsp8/bPBW/NKjGmN
WABI4dIODdgfYmrtYjCstuBolMubBD4l0vwLeImou3e7epiRKPHe8O5PIEez
QA/Tw2xuRd/7IsFw16s7ScQxmuBYQNt/jgQg8bpMSCM/T3Jh6NBoIHITZzYi
MvJlRiN2PB2cbJHIuDRT2onNJzXkiZ4y5gjqwaiKsHfAFjdaBjJBlh87w2W3
9YM1WGDDZTrDNMRMJ5C8uzHM1HBDUZUDWd2iEzE4PH3NZtAvLl9IKyTMX7wT
A3UCltsDtV5gBVBYvNMoCWbqIbIv7ENyVDKZkuWAT+5YOQ/X15+MXMfd450X
4K9X/2S6qnKcSAX0njQPz51MVc8u7oBqWM6Wex8sIBehjVZNrDulgQDKAIXc
e6n2T42IOFFy+LcCwM2P6TLnnxmQ3u87Uq7k/3sW8IkZysGGgXBfHKinIzK0
NIv+tKhMXtvOMJ9tpENNfqF2ytIGuO/ES5LA5AwhMV2FwuXOTyz9c+q4hEt/
KXgv5Ssb1CG6AbYT9Ow8SUaH7zoyaAVO30xbRusYybJ8iBBaP52VaVF1SVF/
M6n9Ec+0d0SF8IsdAROQmtmavI6rmxwIPdDfUaE8vNsF61gqKqDnWiQjGK52
JnDPoGpLJKzli8j3Vff/OwCPucRt03OQ+xJ17t4wiFQVDYeqkte+Guu8FKgX
1GDubSQ/YA1X8KD+GMp4OHlrrShUbUO/jFEDYzIJBHTMHZ4NU4e8eOHzv5vu
D8oUTc4p2IM2alPJsTmNHFEHblZg3gahpfHJjecuUF3jFjYIkTtW/EGH11Mi
h7ACiMeA3ZLRIAZEsfP33e11IZUDOhji/GIgSawyy58qomFiSWZRrsGEXHQs
vK5cwfFJOjKdX2TfX/KmXFbTSbTBJ+YmE0zdrg6YxPrgjzyaKTJvrd36IY4c
PoablibYqh2DYU/RGFekqpd3wegpVjxqfr0Z9df+iOgOxe7APtoksQht3av7
RkPe1kXvKcNdICaeNj+T0gDcxXokQDGfwYIPsw1lDMdb3rar4mSBZKHDgGgS
Ki0aIYQxShkCvn6FNCbkjun5G22i9rGRnkLqGuon5iC/C+omJb0+hTlwvbcg
82zm8iz0Df6naYCxxY9p6y3/S2N6vvwznIzOc/Ik20nDQlMQe0SJ0qs5fgDv
0kAaRPwIa0YFVI9Yz1WPiv2WegmNe4pQURB86z5Pvxfx40HofiEBwWz2hWvk
m9KzIYv9LYSmfti7diehVTy5pfGbXhVbYpdpgEooM0HgxUdJKgrjcZJ0vEV8
wjHSzLs6EOKk2YiTummh/P+KuKj3f4zPykj37OO6zuBxwFFjZ+vrfNuttyfo
vwpQDVVmlGgDRq7dWTcgtrpw0L3UGNoaQUrNQUC8zRVd/NF/K6fJzCAQ7XiG
65VBCg/+BEQaBGQQ7z2+VUhi+dchDcUP9qwtQQnyChh0iZFc7xrxIInEX45d
cAcGy+ikrGfJZ4mMNx/1qwugwGox94zLDjdAi8dkvB/gB7qBlUKxjlTTj0hB
bPnNSjq9IPXfDfg3pHCDmUaeu3+gHue6pTdPZtzSrQquZ9fmR0vll81olYsl
hk83e8A3uBlbCglvySAkAGnk3m/tBd8FA4X37j0LRB60+ENbpTJOCeHRtIqY
OFAS/ZYNGZ7rI5bMB2BDt+DfRUXajS+A3u3x2iLSlpLnL1E6+z/Z3Z86d0ML
SmHIsspwpMF0xeVdu+jreq4SW8wmp8SHCEXemrbQuU4xRRsQzTAFTRwMT54q
DbmRnErKsoK8IthurB2rnyTURYgTbjwlIciNJ7jUeeqUzYmEBS2yWpXrIrPx
U1Vi2ffglMCZuY+V4Px7ARf4V8lhSJW27COYlAG0TazxoiFzFhRQTi5WViRZ
9070viNRyAFw0a3x5A4oPYirOr6LGRsQOGVLh5uuvxMh4ttOX5Dwr/MtxDKT
PoNJLXt2iy8Ein0ZNTEzrerLDfjnUGF9k1/V+jXegJ6Kr/2xJ8j7qzMahzHF
o3EqnFzVaVakO6eIyX10Bej8eaNGZpWdAb1pC+OiUPeDQsNS0SI4UL7Ye3OA
bVUrwpt1pDbpfIwAlWc3dTt5CBo4dAFC0so9VOTWizGz5BJljRqYGPiHiMUO
BnW9UUgir0Zbsqqp4aL5ASNoU3GC3uAr5Ek6zOdTkANu6KDYT+9rAVHOsQ2+
OzKIqLbfahhKl52kraxxttxf7LhzU0RVIC2lyfM1mIzJy4AmT1zMA1NJ8Q6F
4uuGi6m3pIfEvkctuFgxv+wrFwyHOxOrl7KGTutAU0E04BPrf1UmwkgWJ3SK
gRmfRSvsUGdjEB58Vjpw3csmLRwuERmKDwz9o4/OUSfnv0CDI58webxGPd7I
dT0sh3vK6uvfZAsD54Leo7XhbMGDiucIf8d8D6MF74BJd9I1aMYrtBFOvnKt
9qGgrbsVWVUgxi2IgOAxKXIRZkysFK4Nj95jxNAeL2WQvOgIqV4s2XM9Ltca
42mOdnlOc4VoK/IHxqgRmzBmqhj+C/A4ULOsBH+wsc2BE3qy3014rHtFJMOr
PRqVZlHTOPgGNk8H7JCOch5iv3xqqNfI0o+eRtvtcF/MPkWj5v1+bSlxX/BA
w0JaYjMeGXM/QBcrvwbVBZfyCTHzqrr1rDNIf34oTlJR8F76nE8d4TB93tgL
YrdIrgodMUKzvGsFhlDyJ7ax2+Ce3zEvF2iRn8tj5pYvhqzmsf7LWGM8LzzT
ii4dZXTUv385UGq8kYgFR6Fmr5NBYyAkXlqaZmAqrO7Uh0r1ldhGL5pu5D0E
G9dWlAaGX4GnBHE9nGjZoIquyejDHwY5XHhcfe9nTa+kuU45agx8Y29PA11N
5Au0ZCmQOBlMK4E2GHMhXS7FSiZygmDKTtMVtEarKeox1Yw43AtWuy0ka8z7
iPFST3WkoYdlQ0bSAmJFuKRHtmmY8u1kEgFiU3JPfr/93LDuEjf7JOn12w5i
s6KOOQDflziXLnNaHHtx1xe/u2lNzLJGID1h7hALzhWiNKaMjplzUCIqHblk
8luJlptQOInLLvBeay1xNPGs96ijwhsT4JzEDXmQq647VT8frPS2vaxePy8U
VG5rSMm/T3jRn1beEjY+V+2p+37/3DV1wb1d91z8Y3Kg1GveHrHQ0c3rFz37
da5M+ahVWjKpzbWxMBqab3EHZItadX13rS2zjod/pumcFlpgGXa5YjKV+Txx
ymvM47e4reSfwwDwZQ3NxL24DKm5YjTdlBWKz1+EXa+nmH83gdN/fLRtYXDg
oq1SKa36lSvmwt2ppmx7I4TF0GU68X9HDV+BPZDbfXKoz3sA5Oo5M1oX4QfR
7q2IaxewP/sFAGl1NE64IyHADcv4+bf8K35wAhjKs68XZKFNtNiXO9w0GOBv
g38+/ev+V++71CsIFnbPf+9rqPuIKrpfv6cygK82vIL9mwxs3t54tghu+4/M
8ARMbghxa1uHyiDcv5PZZ1nTGbxdQUnu/GIx+cvT2Eo+Qt8rZEAfldsp+xxF
7r8WPORqy7YY1ZoOVXZ3s5Fp/ItaPSdYjLPT+PLfeL3tQvxzVFFy4iuzxY8/
PGT1c4dHu1KhEf94N9RmwesaKuBz0pBymm4SxYZsbwv+AbQc7itBba1h+rYG
TaqoQ6Ndnbgq6ibLnxx+DHv6icOOkYFam2pIpjcqkGv2EwV95/vBIT0LseGj
vy+S7fALPMb9CW0ycyJSlB9mmvIAW0EVYHnrk7Hpx5wL4oKrOOi5+YRsMZU/
TulHy4zwsASgGPF5+pkJkU+a7MlSoJAQQYBFyUOTGDRnjD/d2uoGaeZ3ISUB
xNeTYSuWE2+RWm3VCkD2fOC6BvGZGertfapS8iZKO6TvDdSt8P2nIqGjcPrC
wzjyXxTL42HTiUg8s5g+uuY5RUO7PmoemHSx+TnIUpZV/H43XIOlMkfhYtlI
LV0q//4dqQkgG88lu6QOylg5CphPDYIoHx27fwfHpbUpyXasbOgs1FSAYvke
mfYhC7K3t7dl+s1gAiGXszmL2/aXt2cHMo7JVZ398j8xnhuZ91O999nOiVFl
rxW/STwuXKRQTY7FtjDskAco7muCw+qBabPKFdKNPdmtihVAGhvfuEIj4Kg7
hk04XLFbCTMEzc4vdrt1A+YrcCvamhubaj9qfWVqZgfHoMM9v7Yt1v8VLFOQ
uSppBoYvm53B+Mxm5aXLTWu/BIY+sGrDepCGusrEbM0gYSw359satcuEFdL0
4JaHfC5JVLkda0YbQGRuTnbUVU9mx+A2rpw5RUyRZcXrfCo9bYFz/HwU7bRJ
E64hldMdotE8Bj5B4B915XKkQn8KRLWjSlgs21wmjx9YTA5OH0i+6VF6a83T
JIFvO4tXpQ/VDUi9eHxO0f0gfa+0Y517kATKgVSzbcInsmK841Ej2n14x8dP
+GKAbwR4YG1xFBr4jBjQ7IiqglXLeLGmvtMedva+mCQIxqGNNc2E5OrjZxvb
tfNEiJPm+dre9gOO+MoMivdsm8KVY160eI3x4GTHOhljCJDnwETVEqvltdhb
5mj8OavkH0Q1J2T4/MK4xOAUV6nn5nIDHZFAm+3dA1Stvcw1OloLFnSAq9eT
+SkpDYtmv9j2XaJwY/wM9cvg4VkozOPXheN43DbhI+rwI0hGcN78Q47HuvE+
JU5u/j1meR413E0EkQw3DPDioQ2smS2bajPiaHi19/R0sBDI4Aq29nA5aqW/
TPNP2E+Y60Kl4YorfnBhjD26I9+0F6A50rUbKFCXwUjD9JH5mLvpp8MHztCm
J4TpVkbjm3fcnIhlVTG+MiMyuiPJOCFyEsowRbx7n4FL2YTZix/WbwiP6zeC
gkgqwQT2LxW/F58RGgEcb+Cf5rnhgO2d/A21QmzDpStwRZZMUTtKZBphCVsv
3YW/6m3vddhFRuIalcgIA5KVofRMZp84Do6dfDyr1l7cMO9aYDIsVfNF9Gqi
IpOCrlFTYgRq3cJUps9Dkg4hP2xfMHT5FEjoPnD9lcIThwbNL//s9XqcTMwk
LimCAy1+fWh+o4aY8bj9L/Kmgx19kq/yW2rvFVfRDKMY9XpKxTuGfqm2SqcE
aoIg9LZBf3d5y83mEOdedHAwbtiKZ3mNIKwKN9peIP9740MqutyJmfSggRS9
Hd0sBPCf+44JzVh/LO8qyFFkkDS1xxdFhob5o8GLHrR0UFKG36dgbvgNA/r8
61famFsfQRQd3TaVT1hXub4QcncnhfQRz+3DKRkR7X0Lwc0Kmgv3G6A9f1FB
VAIYMu813OI/LJSL+KR91JHbG5TfUrGQpt0IUh6hVg5wYTpHxNCBz52xiR2n
fvjiy5vFm0ft2iQVXPoOqgf1Wm7a2A5qvARjCGpZNxvdfgoIaq40gpFhx7I3
jhd/A8vmaLBm23DiQsC9NCFvQAcFA68G6qjB2d606riqryFFq1CrrMwJDM+/
bXwewwGAANhtCtAxUNsXbA1AYBgFVbE8kBWxyUB2VkaWhb/14s0u4t06fALg
qTMWGI1Yvz9NtRo299VC4x9rL/vt+Nf3fyI7vATL6kE8atjZ9KuKfkoQW0xx
VWjVFoZifSfQeN0QQx/bKAm5xgtWRcwti4RhZl/GxUV522ip4TBmgJESedD4
Zp0dgsoTus7LiiZ/zW3VRSwdgCfO6Js5dfrvcPL4oTJfH9hutW85wbOFWGYE
KfTqM+MOvlG6keMgqnDndJhj0nKFDg672UGGWr+NwOv1pSGQBjjmM8HqsPcu
r50bZSN6pFVcozFwF0amogsNyZJJFHxaY7EG34ok7NzShSsWr4DDmzjTPbXd
BhXiF6MZtFoE/eKW0kxBxhVFkDvfiXBXXDzSCtUk431lWfZLREepTDRoukxP
sFGyLpywBfLXa4ADhQsXTojxuL+u2ARW3PwYxMmOLT3hYzxJY86s7ixiK0ZX
kGxpClcFNw8GvqnHLzFy8IMC+ehCNomCvSrHufi832F2xvdTvwK6KZ6vICqG
uAeTmjm2Fz+PkUI+jmgvMqqDWgnQz0myh++xXbgbLul61QSR2Ou2pKc4lcOA
d9utgeB05aj8qjRw7JjZ/WwObxnhDSYofb8HlxgRJRAPL1WhbbOZKRb/UBNm
grxGCXLOItWeBMRBJnXhhxX2Oyf81LAC2bcOvg/+nIhO3YCUwpRaeryPz/Ek
ZTsp2vbiasodEhQtZdHlL14UIokfxZKSfc0p8vMro4+9W/bncUnVP81A9UwQ
628IK1CpdMoL52RjOLsVdQBhRM006DeZh2vhpkrh/ZKxths++IH18Q2Mr0Iv
XxBuQTzIbkNVG/AYWflxme3BBF7QIRbioFvpq2SbDTndLl3v+KyQkrLfYM9B
10gerT0X3ZSEel9YPnEMpGmCsYOr1PtV7bZb6gLR+ZghlURQR+hY1eb+YjZB
+TlJN/+XzMkMnShDn/sQejPxGevo71Brg1S7vBkwWBTPCv8LhwQIrXnpsCox
tUnPmfGogU0SNr58nC3BOporfPu5I4cZf0IcjDFRGxOp4XaDLQyiLAX5ojM1
ySMpXvUUytGwq4povEuZ9CTtnlGIWtD3yg+cGYVWKiIkkt2uP4/AgmwNVq90
nBme7DIsXcH5emBPq6zlMmaq7PbFRMaSHAVG+MqToQJnXsFsX+X9F31UzI7n
EclKPR6/R6rkxapSfRnaa85JVJDNPwiFmyI14wu0v4qXev/LjqNBuFRT4SyS
9dFCO1UiC8GYcC9tsTogKxdLWSdZTMxc/nj8tFye1MDRf6eO0M29C/B0l1aZ
vVxZzIlfMYX9NLNuxUwZ5Z+bZU1J1LjOj+yML8MTR2qvYaiIgkEFLsR5soMi
5pL5dz56SOcBCmhFDOuJc8y8/1iHZJ4l7WH2O5U2EjBoUg56XVt+d8mVi21s
aN/kv2Wh29fEId2RwRcFncA1NDhRg+KVOGIJbKu3sUsy3a2TkdedSu8M7Mcm
RerXyyRwD4UyJIZevRoyJBrsmkGi0AIuQcvMuFvVGKdOh9DyXQwl1nk0skmg
9Q1V78DwYx7yPJBn4Nd4kC0g/AZDkemM6aOuu+sg3+o1/XThbJDa4VtuxNDM
7JrUc+1/CdA/6MTlRdTzp34cUSg4mWsBNl6WDiCxstOvco+SQEiihJkZpaMA
Xvx2kL4eqHkqYl0cGmjfmrmKUiyEP+gQn4E4g+l5AzAAs6BtDoXCVyaFv2V1
VSg2sR7BKYx4fkqkC1W9HOzkWptB2FCTL+F4/ksDp+p1QkYQxGN4pa7yksTe
KJlvC0a8aZsJvADm08NMaIHW6KKrVXsGTQr/ZYCWdJLOmhs0RanX+Kv9vwOp
O7ahjh40zFZpGipFeQOy8bwbTvwWzWRyCFpbiRkJJiN08tCb8YAwBT9vcWQg
0g36k5dFLZiXcy/PPEJ1TB+XE4fkSDXIP2maCnzPZvZjGKmkzBChdzKG1ho4
H23FnLV8Ph/fsSM1RJ9W2uYyeFuq4X97LC9YRVlnMQaMUE2igV4HoYwsHBh1
O82IE/oisImdOEnR19f2+t1Td8jI4/Rc+d8bdOPNsUCRpm8tlIuXghOkTkWT
i91LaKd25i986Hr+AnapDxkIjy4QdVZ3siUcM/SkfLGRon+iAduyekbusIg4
ooxx9StXBPvBF9Z1a0F1QsMIReyIsIu8RwAwdLlQThS0MgpGCqN8CprZhl5r
RFoWoQCK+mDYK96FRa7F6qhIW1pXqyWhqXZhDqSjAlZ9t83w6sgv5+AS1FXn
+SJkHjFpt49dnvAhiLRIssU/0V5OXWG8QWb26KA6kqXBsrt6PwLwR7ajNJ8L
LC0Xnvnsc6HLAebhDEXLsUX/KDR3b1nYm60x3h/KMsKd8dJJn85vZa+gwqDR
IpIhYXchDd3I7u0KBSVqMKhzYzfqb1CrOSnDOEuSoXoWy3a/VHQ4aaW4O1+R
CrZrwvCiJ4goKNcejp9F7t9sYMmb9ltUWgvkke4x1yCjf5KYpxnxrBYA+1K2
bWohwUm/p1yJwMbj8MvZNZNaQ7sS9QgH7dRnG7Y1PFsHlDGJD8/b3rbjsvr8
YwZpUdvA5VeVU62GVa81Kys65Lq5bQ38UrcxEsqm28r133ZKTkQ2VKn8OPKz
NJ03lmY0sfQdF/kDvDdnvOOIncUQ+mDv9zR0SNgzwg627wVNFZJLyes3ztiF
EG5YKYsoFHVQEC3s5bZs+lAc3L8JDa2A5JNf62UoNxk7OW9F2n/asRK0exLX
7BjV3ogFnqPoW2PgbCVK2Yu5OVqBdAxolVXZRFcvmAYBd8GQLAfQb47Svorq
zXtKaRNXSolKNqLJj2hhT8f4E6s9D+mEJquyNBnFtEDym67Ogi45FC5YJLss
MPNUDGGU5PTncukm3ParNlHz1girevP0lN6TAAUNU9zNkpvIl/OJjuURgAKu
6bWXpUQORBesdXf7hWgNJ67mmARRc6G6ptmkTkEWCTyD2OpTZ2lg4KXWvZGe
kvbJgsZJ7Ew1YasjdiuGjbCBt8oL2Ne5mj5SUL33192HbcylqNSEhsGgo/SC
F9/AWYDfPPIu1jdwGNOa3jrYPZHTLIoyIQaEcUa9pY14vII03CF9VjLQlGk1
KR8Klguz/yBrLcqsx1NzqwvCe3PmD6HnvVOnjke6+fw3jA7qgybZxwYls7LP
B/JwnRSxzj8gufD/RRPNjvJhsy4zotarWmikOwT34nixHkLimbSrCJS9iojJ
lSXL+1dvza65wrSMSC/WQ1GxDPz0paM3Sym/WXqRksJFfrajlBc4Wr0byJ5X
7CT4H23UDokw976v0FsLf4oKniqucu1AnvNWbvIsbputpVXzfsb+UN7y8Ibp
aCkYmqjzMOdoGlXJcA3oAUA07ZWqWcidTVVd/8bUFfSc0sB1KeoPeAsi86FP
0bBqbrWhlhBRytMmuAHOvoXfcKLwCviRJ3pdaErJGVjO6w2LmF+MzRuoUnLk
UyiDvIHktvJZXZxcVjVXBo8GjkuziiBptnW2MHbSeJAB/1lsyxPxlfLKOEnI
9zSMhUPz+TEI86FoFqym1ZFBqh+OaIZMHt+BR/sOfh6ID+LRaed1jlScxAPH
TN+/KgAtCV//Asx+auCV+w6H2RfUpI0XJgKg2qLlw3yv8QSDMu5FXgk84Syx
JgkcC+3tLqoNqfCNrtAtW9L82HXizleixJ9tMJL43wmBw34f8RkkJPS0UZeh
GzJWoUY8H6ypZdIOWnFz2q9P9y8tRQzpmWFPKEc3oOQiM/q8yAkdqVZk8HiO
BEr/8KGjsr0OQiafbVgOxx8AGoVSQZuPMtT5WYrKaoHgtMwlJhnd1xY2wp2E
GIjKw79qc4eoDhC5CzD1J3W9OSh9ZcAPhH9X16uh1oEzjTMnE25ulA/kyang
De2jVw1Se9N1iS3AOncOpUYjOHv8+1Uz/4ok/nbmEFSUebieDIpijAtKsV5T
kV+iOrfY8vVarp77QLMIzzbXGIv92j1My37Cg7GrvwK6EWodULsCz4hAFx50
OhrNQk5Oj/czd5y/f30CNPWipInesalVs1SuAtpwHutkINWjH/pQ8xDkVKxA
o+1tpL2uHlkLTbja1Wsg73WG9uepjGFR10gLoLCFS1DHd+CSpPU+1WYphBIM
QCfPrBzD//RaqpJ32wvp3Vqo80caj0S59YU4wRLDQByNmubbkk3/gWJ+9HEw
r+DC9Z3IczsyxnmT7B+uvtt1Zo96eM++WBmNluT0UpKdYhqLmSPDuIY7hUHF
6CYs/LGHiKjrOq51g091xmQrsM33sxwCEtFnvXf0gtObq2AIiE9Yz/NpE0gW
c45akpvDG/I0Ur7Y+f8K4UeAK2k7qpvMJz+FnwgXsfzXP0lHnAW3FzCaqxZk
/rpf3KMx7G0bBFygZpmPssx99mVFOrsAI6ZMliiuUTO28aG7DRsj7W6lIany
w//UMwGmjWw3N6cTiZ55HHBjXdJK+LtKevfAKDLHs8XLLgME1T7+Y2rTi46L
sMru2m/QgL5/ewF1GqT+trEkHZ/a5KCRZ33EKF49hQPG/YEnoZfzglX65Gf8
TH0k0tBFRXHdOuSzGMa6dIRfF1k9beqi94qLKMSOsD4tSTA3T5Vq47Vze+vA
BFNzm+/lKl4bUi7g5oYh1YSWuyge2vWPvko296pQaRPTqCDO/+R5C5DCTxye
AazVfAyn+JY6Kq5TySF6/Ge+i+TNkSzMIBJEnAba0adpTZNrnLDyimK+mfMl
JzttKnQuWrnZUBHzS0BFzcyARF1LHzz9Z2Ab3DczQBO7olABZRbA79/Q+aE5
j6TM4WyD6popKop5ETS9pbDwDsQXHzqPk39hPrYy3nGb+SpUF2IUyr1VanJz
kxRW3tTfq26frmSMbwUwwCei1M2qV/Xu5DrgGBj559UrRpBMoQUiQlKDxl20
qUMTy/omXV3vzIaHQ+pKzmEO11AA9XcfQWpEbgGRp5RGP0oUiI6Bo7+tBEIR
3vBpmyXW/JHvPIW1YznLtP1dyFHh9YjFHJrYlZmb4/HMZY0VdW3g+Ay6Clo+
SdXUGYknNKkOHYwXXDPQsnf7Vq9cXwdJdmsh82KacTmzFL9YGzk5++5KHnth
k9Y6g9wz2RwxHpMG7xatnG2gCf0A0gKlP0+7yZjmN2sT0a7JqN82PG+ZYtcK
fUnus4fF78Zkgon8MlUfDmlneQ5e+Phq/y/C7nkSwahNaB21jeY0FQdMu0GC
gROTOc1ahz+Y+DVlpaghO1cZqElAMviHQHyd9WhK8v/aIp+XXZOTpPiKys4J
124CAGIADM06Iosj7/dzXZMmptd0qM6xJCeycV/fQNv6hkvCCX+IAXBsCu8B
s5IkLkj8G7maJreW9Ppl4sWKAY2P3cQLCauNqg17+LmTCzOD1b3+xOj4SYsq
URsX+KzcFkaf6VsobreUnbUeumgZ+gU8i/mEuAm0k1k6NFv2GvYyGbRkeU44
ds0EGmValGfTzvlYttISFm0afGJVJw9MHjc294JNQmFKf1C+HSvGZxFbDjmz
IUKZ49hgcqjroFxCm4bxsZV6VBKjbhFpenCQrF61jELVInLIDDqWxpbSHfz3
YyWT+BNJy8i6MGQW8YcSbe7Dz6xHSvkv7Y2H+xlOiXVEJwnW7eG1sNoQNpZg
aDGpwd5GRues1nKZ7qOimV8cBthAyMd8FsLsx16qyrYrfm8a31BE5tohYaw0
EH9wq1K7GFtbizlCm4NQFo4eQO1cVLZRrTDbO4R+3s9n6q9GPw6K8qwrFqrF
t8sQJpLVrYoAcg6yMV0RsWLqcqurz/6beeqHhIdkQHWCpIQoBtWegLlMnBQI
CTF4/U9DsxrpBb8Ilrv1hy5PiEv2jlNBVXWvssD6O4AGKSYvI1a5pG8/B6r9
gEQ8VQ32d1/5UNtvt9Su9G0W0+S7LOlxlElSTIVd+um9Tpj8ylbfKN0FTvNk
SehffLt2FyoHYx9MaxG5WLUq+AmghbmKwG6wgmUrgX+Wjc/49qGewW9ovObI
tve0MiYYv+3wDwFipTGCwDdzsGU3Jkw43/J+ioMG0hGNI9+7lds+KsKwWiYV
rtoXr/QIKxfI3iNi07VFyiby60x2ij2L6zScmwqlsZUxdE8ycGYJgcmg32ft
PuYHbxirvqX4NaC66f7lcSK86udTH9/8tg8Gw7MSbrjruajU2xQWpU7lIQOn
j2buRp0W0fP1P3eYzI3oxi8Pp7qYQrqexw7lalEOsiVQtK1SeGRlNWPdv0Sn
afIcLjQFEvsQxat5LKvSGHzYh+5BvGCRLO4JJWLnrflz23NHGP9lCl5v/XnH
pKgdjg4pwkHL47UmMbAUKaldgAY+dtQN1XtFQ+ixT57QyRwc8rnjd/BQpYE3
IiKuYbJK5f1h8XG2M37qGZOEZ93fFBN12HIrgSqWROdOwW7w/dg4s46QT5rw
nfEpUvJta3xJIPDjMDBT4XO0QojomxMNfdCD2U2RY9vGt5Ct3bqNcdr19Xvw
i1kbFZPd4J36ZMotuFSD4ZIue3baemklmb5RvZ4Bog7M8aGweEqI38k/VuN/
hbpW1oulqnHZKsKyHyJtmyjM072bwaZcf792+QKbrTD7Z38vau5B+qZLJayn
1KU1+9bXy9SNTDIsIZfwsjyknv11g+SCDE3elKTgCs2EnjmFsJ4pwalK9mJn
j8q7Qs68JPDEt3xz9zTyTawBncg4+5W6VX06RoJq8gY4kcH946Aa1r4DfKJo
vEz9ZTkJfmIiKAgHRP0dZvCLJtHqBHxtaBXyRY9i2G/NeLyJvmV544R6Js1n
/WjNn6SkcDemfqW0kdn9TZlBmEGkDH1xjeO5WAk4r0teKUGgSCwBbectzDyS
sgJ0qbNt0T3Gz1IuiKx3Pw3GguXeFusD0K6/WT5IMG/EDs1wpCyvHp/lbmD4
Bd8z4SvUmmCfqbp6Sx8jpE23FTzRODU/0LOnbxsXiLSDX38Zdnq4S8sMrvVc
CKTaMpdkKON0zUG1qGg45fDZef7MIA8VGPgzlsyOPyS+yXZMMINSzC6skKoM
jY+ewhmE1arrKQmkeNpvgcUz0fKy0G73dSJwvEOHQFEnKeXkT2CKXnTW5U+U
tJ4NbGIwH8kXIRNsGxFdMp0jM1h7OW+dMRNpLHPHVcAVC/2pJgoKx0zZLDdr
Kc/R4ScAss2DnpRXXhERx/WxhhFdNlYQ9/ez7JW11vG2EQ/W4BX4fB14NbSy
vyk2nFEXM4Wdv5R0lLa5yEpDfaahp6oJriTqPWFyPpEpYdylNz/MfE9AjKUC
iLkkC539LXADeMQluzDY8tSQt4PIyb+AkWRZIpYdhN/SJYyNlnDwA8IlVl4p
yLXilf6BTlza6GMDkR1W1Q5VHElited5gwUBXc1HNGcP/kUIPn1ZH01oHYMZ
eGn9Tan0Enmqsg6IYKXImCmm0aK/sgGMgJCpy7B/V+vFUHN1maN3ltNNjaiz
ZPanE4STOwoir41rQrIPJkrsRKu0YPHv7CtX+3yjQN44RDc5AmGIYx5DK3rE
NxZq18c9zv5OhWG9Xjw6NNyp9hpOoW2fpqvTQBU8krVx8MYVVLMOPM1JbLbd
fif1k3bv89zR2NCO55/GXE2znBpCUiXCv5QAaJUXzQ6PR8LcjyM0bT1b1yJY
K16YcWF3fF1F8zfn++yFYrCFVkYlXgXbNSetvHMBP6QTVsu/H6cP/m2z2Jyo
vmY5LxAaDhN3LofnWXFfudHvFalvj0ChdHzQfWje9SYM4PeGpOv81Gc1E9Vr
G6eFgyc/fPgmqdRrQ6aI4R+IszV2jUZrrQdjx224wa4o3S6KsCLboPHK8jTg
6O0zCs1vAR2STe0VPiAyCSvBH96wHrUHoZ/gi0IjSU0GlBbmg3SWcL1kExWL
pgYpu72JakeiWrFj8Zf3SSjg+NopIPGB1Z+rLCeKpisq6/gqH6A2WyKu0X2o
OSaetVcmkmKj9YQNseM64+c04eWTxg/72j8MMl/Jtsg/MUBqgxlIoBzorm/2
Gv/dGHItwkxMBsh44C0wXY30PjlQKlvnmhUZBvDj5y8tlylNcAjGcmE8OmIm
AweSrB/UxXybri5pCo/wjsKDctPI4gCe49q3G3acL92Nz72HOnlnpOAHEJs3
6uAM0+GPX8Zb4pQNV5MvQUtaj/C7rK8+2iXdaVF+o+gmTskUYn3pTN70G/7L
90mvLesBC9g278HTFdGZndM+8r/32n2Iq/IGSSI+x5hKy7umUw5axtHDZf58
Z2x2vb/gv7jdcL4aekRtbXroL5C7rTKG7wM1HuMWbfyS2vVgTl7Uk9rGaTsJ
QKIG0biUCkAEITkHRsUz+e27tBZiPSow8B3JHDxwNoK47S1m9ukjTpo6AC8D
mJ80G6UWniBD+OJg0W8jdJQlamk7FTtkudddH9mtBdxvm8gs4r4TzTrxIaB9
t/XTKUX/YFkqAML5IrdVTzcqQ9GDbTp+KxjUCEGd8rCEIANCra9UL8YR23cb
Obpuh+6amVgqH1MLxVpPHxCJsui1dJvVHT72qZg/NT4X8GurJXJHAQAS4oQn
kL0UVMHB30RMxB81s2z1IuQuMX9TXlLkdNQqgDyYQou7dt6wWUPYrAX2otWN
4LdSDVxulO/IqyvkBRT7cnEbke8CPFFP9UW3/WmV30rC4hRKR8auWhQDX5Yb
10yKm1OXUDfcUkOF1Gn4FdVGRwqrfr/MxDh+ZEJiBHpwp3tVq0dkoiwxI1f6
6H15BZ7Jfp70ZL5+/yQuhREuzIfWqBnYMDM26t4FgOR7zqmxhZSg3HBp62xr
y16/2iDp68mwqgVc4kdz6YVXvrJ6U9M03Jj7HGkTZBtdaBmLsn4AhMPNsA+2
lcPwFGlisy3dzmlphsEbWa9DJQiXXlLOs+3wrf4rmcW8dIFMSyXBujGxIruD
dgqhePh+w8TJizfnDhWpApQlljoye8+LbSF8amKndEyHhUrYSHgLof6sNqQ7
VDJLXTra0I430X4Vobmu9+xaMG4dx4aBeW+ZdXk2UFAttd9oCUqqYSGirFOt
sBk5iQvkofRWVsWKuy+eNuOoXcykNTs3y2anVfJ+D4JZ0r5ZHzGZGamjyF7l
CcOUX3zDp7tVcwC10ClxBdkHSbV8QuUPs1dyfebt4luNhcV0KHrnJIlG1CAE
WQnOQNMM90lNeIVu8nZ0Tn8phimsAKD4aX3yHti7hSScpDc97VY1v63SCGbD
8WEgwscHG5hJN8DOrkdsb0vcd0eioZr9a/KpP0j4XT+FJ9DgtW8K6AOcxy+i
hn0OmObGGLKJuJJSch7/8/QQAXVh9GIF3M3woNMxp9RVy36aPg1JgNrSooYp
tQAi6XrYtqK2tJulYg5G7RPt1eM/L4+OCmIvRJUtXdWmrCE1fXxkIuwAR5Nn
cu/0dZcBf30h1NDmoLIVqSpTU4iblXngfjXhPF7UQ7wvVpFYfZKLtBHauZkz
hnMf+jPZX7IVv+a+g+mKnqKDL0ePLaQdWdUkSuUvsfHqwi3r/EIcwy0sxGXI
pq3yvFryJ62DwzLweAyo88usVFFfBGNjnYEzFCFSFAY3E+/Wq008NyedYYkw
9VNP7Fu7KnT/tNKkGGFbtz2fAMYiQeg5L+3/XXb0BvhMmgZoiXdwZJX8sHy/
buSSkjVN3WMXG4069RM4p9ZQtQclSI7fVlaP9An4W26jfrWvds6SyUMDUUTP
CNx3EsYjExHhHYqQY9VNODAbfMH1UjgYMW2O+nStYiWrezVhYCcr1CUolY2z
Vb7PTcdiITgwNijD6ASx/OkLxTwq3tt+oHiaxQVOaIpFP2hU/bjRERKXneu2
qD5UhQnJu1RXF3omA0Nr3TKoRxOeh/gCrQ/BV1ozGxOOpRq27p8dX/k72ZSG
aiS4U9rBNU1fiNIIWIM8Uuhy81orRYG0MYeQDyehJx9u0+cCI4GCyiM/NKW4
OnIfW2pVX3Ovi4nFhc7gSbNf5dB6PvKw4Hs/34kaDaP2hdFCLSvr+bGVuMbn
8GVtmONmW5vzVkH7X4v21b11bh9O4vCnr+szaWZpy6t78ibN6J0jixGRZnY5
vrBTn9WT/qGkHPIAUKFitE8roNw49LQNaMRYq0P4JsDQD19nhhp/+4F/NmI8
YnAwfDBAya9qHV3svkE43I8jZaPQjc1jo3gAWPgW0dW/REUIxNlOrGbqrcnj
NRz8PRfy1qYwr+ndKd5jkSQuaZwseOsD/uEfOP5TzvSb2eyODnaqQzsRQt2Q
IBRkX0ZDm6QgeoPisE3aE6OGwejCmPEGRnVKP7zie+14ozPTrZ1toP0BucV8
Ow+L2D7smVAaQGD3USPTEUNgU6srWd0XMo+Jl4JQmlx6kAHXfpzQ39BtYnw1
NkqSQ1mPGm111STMAbmLzAK4AiIMU4am5NdCRXhqJvjR+4YlGlnru4r1WK2C
RL//6e8j+TPG/GMR4Yriu1jpJ9cFueli1vZLDUR3LS6FELTc4fI5dLwXfg00
BmOXDHmVZrTUEHWa7T6HC0qOOqlCW6Gi/WaZ0/siPZgxWcdVBChtu7SYZU1t
mWSK5eF4yrdHmEYhCqPPFg06kfLWxJxsmbm0BZ7/BGKqC+ZNhKwbB+Aok29Z
7J6R0qQ76AhrPPD1O+619GgL+xqMdURIera5EU6uzEImWMHV8shUTYAN8RoC
9Avua8XdM/W9NgXQwVoN/izLY3w/tHv9/7ambR7LnWpJ2zEsDao+hcCAwsWq
ShEY7BaTWX+dzLb1zWYpwT5VhAd1uE0IX+GZ1YpMFBNIAWoeU87+Nh0wHEjc
i4Jd0eckDgsOhf+W0IWU2yB5ijsMJju33I7bJoKAAaBtb/+ARbxVU0FswWCH
h2aHa6SUgsSHPJdf1RfoCKdciMbo0A7Q5RMLn+LshzdaSPD5fzoW/MBtJQa3
Ujya89uOQFcCMETxW+B5b++IJgjFuIVYs4rj//XbFcKP6FXqjNltyrzAvAMk
D9aqE866v03DFYhsHh+6vBwl3AYVlX3cdXAo8aZATJgmt/lRu3Bf71VyM0o7
1BfqI4iLGLyRtfizvbCt8o3mo7RT9KOaqI15ZJyIDy64kImqb+DdRBHn/7YW
66fSy7lCHfGX0wUqmsEHpry9AsBA+bhFiG6i0B0NTb6+h9Iu/3JSmPMRAZpI
E2VZ2ccy7D+Fyk0n9kJwTcv5sWiSp5sZFlv3BE4cE5vtZ1jwO53uLs8GQeWQ
gFgMWFhqzQjgqXUEk6x3iaXSrb19WvPgnAy93RWvhSBuKRJNqne2PkPTAMK6
EI3v8rbwptP+VWZd4WlGlevmXEgHF5r5UHsBk4DOCiLxaB0xjhUrHuEZRNB6
YEktWJzn350gcDLvgx5sVRldytTBQqnM5C4ZNxEE9Qf2nj8PwpPeJ8zJ6fZs
XEtVjzz1HYGk1hYMXYwjUZeqm/+LnnhL+ybPaHSlZLsPnITnn5LP7pYJ4LR9
G4Pbd2uRIz9fROMMw9YwGr/oU6kK7Oon/4H6Mu0+Mt4xMa6yPu9/78IPF9p/
3SyxfJ9aVQlHBk57cit9efE5UMA1poUw/smLrVJ3yeBq65k4vuUoBJs7CIcm
yg3fyJkrdmJAYrztaLDlbM33qORsafESRlqOJB3I+Th6gRc/PbtcrOFY5OX+
nG+ihT+WWjO+JIfx6l9GCgW7RjASH2ESZPiMhXAId99Rg7XmfdPvn9i+pgd9
mLTbAs1qbOlUTi3gM1JiuKd6X62aQgrhbaj+ZMnYZmSQWAb1vYTmBN4qcq6J
p6Po0ca9h/qk5Udf9h5kYAYaLv7cOcnV6+RXm6p8iGvURGLzm9KFnZtkoPHJ
4gTd33CaDKId4bv6/sXc09TMDcCsVCctuZp0r4x2Mk480jY8O9w8Hc6HRXiv
m6jTrsOGRx4j/NDU3c3lsZSPJhD0TWwhhQ5+YQkJAMOYEMI0XO9yGO1ReXjJ
VXlXV31w5Bkswtpi8itw+7ZK8sOZWGkpUk7cATvS6T4yDmZEwyaVWW0EPn1Z
E/xgvVTycS04+/ItL7BMAEglANUqM9FRaWzdQrCipTfkojfvUDqDQnrF2+V8
sySiVLoGdn/oxkdxrR9KnQ1No+Fc6y09/M7Qb9YvCr/Y6jIJv+2ip5bAX1ea
Xu1wEZXuzX2xryoI/H78qnT+Vt8aumzuyPeaJoqhMd4bTk6zE26HKH7jXu/D
fN9fcLJcHIYzb+rrVv2ivywGz6P88U3oVvhDkIktMiMUHQhdc1fMwFJixRKj
L+QR6ILdJsHpHCftA2jvE1cwAphMaNmCZl4X/supV7tYW31u5FbCaTNDYp+t
5Lqr5x5Y1iH4875ua4+RIdV8ImGrS7ZChGvLUe9IB01pO4DFk4cpTYt+S7fA
+Bfs4FgUR5+5WB0WOhjxpcBmDUSe6BVcd9bMtuMk0OAPbODtHsk8wyiisCL6
lpEuZndiu6xPglGkUsEIFdw16shW5GLcxyD2rGPu5dk6L6mjFNhm6Vdu8Plp
yLsdKKwGUyfsUswado0iVWvrLR/MY+NWOV9dcGUZk+CgX2XXISUEeJTLajQj
pQqFDSkH4fMc9l5eKYrZKY/59tdiOzTJfro7wmGeFT2UtIiF3jwD4ScxQ6px
0Uw++Sez3ELwVgR+WeL5TQ8YFaxBVEaBdjD/5PqZiFaZiaY2S9KE+THgqDtP
vSjFxmpCZvmkR8SolgtiJB5iyIY9apNyAZZNRlMS3ey0EgEXNzg0mL8grKmo
IXoNKqc9eYT2hjlKLi5DG1AN0GJsnmzy3/C6nYeXU/0KI5rvJjQtmlX4/h26
8qcVFVrcyDDR/0DPJe7fHEirlDBuRuWHbs7ZdyarVXL8DaPeDfmkftt9XoJq
4vUfY3h6srNciWVrDC9ulbo9t80ZNWcpC9TfQ9Th5uj5YOE9oAigbLyMh3D3
/73vf3SGR1KxAYieVwKd68Jg/3pO2ohDKK2x/RCgMMntHkvyMYTjMGAIZNfr
3QpKeK2NYovxo8SCe2hrC1d7zI5CpEv1vaUcan8vZRp3MXhM6p2VDhaDrNK/
CP10VIbpjj242u/ocrVyZUWh8FV0Lk44lB5CVu+hmHqN6wAXUIhqBfuAtrXK
ms6VH49c5AwtJVIqJ4hFj8d/LIdNjB08Io8WP6AMz8YswA20SvkXmtKhOiFq
kEe0Hz6D6ztbTBwdi+L2CjsLqDS5UPXzyTz+eLkrLpq03dLe0f1+9BMKsP1F
S7I7vfakeTUIlHDtNOBkFTT/cOGOeEOjFDkikjl3+EuDC648twXE1pqxlf0t
hTJWRnGrTJXKnpdD7PUnlvPwTMoEI/82clKxl8eOXJpSX1ZVoUV9RZKObYBX
CdwU7WBgT/NTYF3BK11az4kfN2icIe0HQ0Ip0WKYL4PbH6yVxNS77tB3kFkX
edtw6IcNBmTgg2p+WRXsXjvs4WATTkh938O2wURyExE1Izrcw96kTMU2+BiN
KiLc2fl5M7L9KkYNs9GSPUawQ9jd5GOIKikzXaSlQIpmF0/Ki5w25IBRIAgd
xLxuHoA7sidY2IXA8Ml9Wx4iYuFhrkHc1SossXzHaXav8ZM9ZZVwGcC7d9Me
lpRdeG2eFrCfLTY//nGdcySO0dRF9D3krGDdLbOQsZBcct/piBHWFSZgYWAE
/hPZlIhFozS0uSLCCSyfwZnKSfOiwZ/GKlI4AUvs9PKfOcUjX0aUTRMRz9Cd
AbwRWSg1wgR99ItN35+kWi+W3KB0+aB4lNhWCNBobrS2FtGQHSd+qcOD4p52
ZVdGrpAKoSfge3wLXTxNV1a9E56fxyLZTvGShik027TMkfY58vJ+5HnSywf0
urYFMwQkK6GJFT4c1LJjRuIukOu/ojlMSSi2Wb5TnekQf2Jd5OPEGR+2yL4R
wxdVlH6hLH0qjxhshzWE2cXZKiPmfGhuo8CaKFutbEuZAsgLPxrj57JK0aUt
T60jALc019Hyv9KKTx2RWp5ePlzU+ldCFK6q6wrKWF2S+IChfEnp4bOhAUYs
TzO/2U6v8p27OYYEtkcZ+hy39uW8iwNWntdsUjKS0NLUBFpl1OhJAeoSi5PA
9mpAbq9fw7VQLfJngISKuNmFZ43fi1k6zCHz/Hqym4Gr4laXvfTsSSFjuTDD
HtMrbAJpKqNY3l8VzCS71XSMv2+n80DLFvvxthzvSN8BkP56+v7lQz8fVdc0
M3EIxBmmhXpJC1PLJpXPuLT8NqHO4BYCVvBrfayi+kwI8liHKbrJmCNUtQ7W
4tft8S9+utzpuQcmvhpter//fS8jymlx5eLqvEhbiKUp2SqIFbLeYgAkJC2P
icUyw5RPGHRtCBGALEzgBp8yIVlebc/FeGU4dimWZTCLJDpzhiNCa1Auv8zu
5KBFz6e2yb061VvICwov4yx9f+s13AzCxPG2OMFv4rVz+t5Y9Uotku3qogo7
M5uaJ+FSctbH2dqcmZOO7xzO92g01GNoPyK1wD9byy6smylf13NbkLuq8/Zt
E8aiTKlcsRrAp+qXsChwm7DyOQQgzjBLzkASucBSA+Wahyyst+ib5vDDkZrT
gPvH3SjRFslnx3Wg8UaJF31bgdqHY2qAdt6HHYTN18WKqBTcVPccYP2yxIV3
DDzS4pBlwajqVY/A05SbAH+yRH3kf8p52+/j4EQtYFjZEsfmgstDbRQ3R3Zr
rgwgWe8uA01JkciQUzEWwPMXrCdbjht4bN15hCwViruddk76w76AbYS1fYtn
wTrrXjxDOcwa5Mp/7oAfiq2tiP69XbbenQ2NdmXkYW80oqBT2DCAwZXjLGeR
LLVKVxTbhEGZmfKOAs5oopGqgD8wt7DebNSHYNaWKhydx6j6G/LdVx5w/0QP
0SwltwWtpsjUjMizNWg4Tch1K1kBxli+qnwi9XM8wbTyg9EqFll4BKLugkKs
wBxIpS0ZBoUuMIX/Ln6RPzBqawb4lJ/CG3yvLD8GAhJ532VoMkQXo6aR3H8J
emTIbcreMgUDa3Tk5MAw0yreSgV6Kqxsg9Ie+aMajD6pfQRYTyYWl8WLCaAF
Mi4hlQG5aMGgPV7DqUh4AKdc684udIP8BdcNVI/p08X7Dli4FAikLtPC+T06
hKTTR9dE1nSjZMCXyb9PeY2UjqrYjp6/cuHXO0q52ea6yfZv0Kc36A/gFMeU
cUFi4CCKDGZ0DbHHIhJOpd5wMo6NOujYBwyp3Gscjc98xkfE5PWzziiFUWGX
DMMs+hMJAvgU1f/CiZotb6XWy+JFwi6DvQp3+FNj9yqD9YeB2kzhCV/CxTS5
9W2EUwjtkAT5jam8jjGQvXjL3DNyuoF4yURiECooaVmvGTjHGuQE+lLb/vxC
svOq170ZubAqQ7TEATBXlzKB69vM45/d7v7jVLjJjO3rvkxcQeSZu9WvaHFc
9uQl3NtjxtdQc9CnzWtCsYtXbajDCGtegl9kcdFB5atOibISRjUtfnIluEU0
eummFci4DhNbZafsIGm1+K4x1RC5tsXIvX/K1m1KiAUph/CYR0VbtF2uwJEh
1nuDufRSNCse3rVyOcM1K9k/5G+6lq4cVViEWGGayh+J7J380RlXFuWlCh4j
cJId/q2tjqqq7932+BzSmn+aEUDH0C1dB/T5QEJSQa+/qmRsv787rbBEV9HN
5Jv+v83XJs3IR4r7dZy/GZd2L++CuCBsV9/QtpZ2YvYKerjdPADTKAqjvKJH
t+xqYVfnuAkTKOUQMXeHDLpmC7KT0oTn4Ui2HWrxMTb29KVkN8vYM9KyRYPV
I8yIPDDbVjq4GCBViNtfA40x7KzGO23wlag1wQ9bxrT0kpvkeVz5WiQ5FuRr
RDabTLX3ATLKwC4hxKGVsxlWAJsGFf0Q5czEzO10fOcMOEzFI4oRzJPiSKsN
ldiHDQIsYuOrnjeuazOcK7nZ4gjJpLMabD6tKdDPE58NfgKuMspKyZYerWBA
r/xR95aCC/YcbZEY/eJ54mq2omFx8RFjSyy3Qk1F+1UbTw1tLAFkkv9yB4PQ
txSLHx4JgYIukccNEzIfkPKbmQgyOnMDjg5gMKpSkSfMA/8r0Cf6W2rcibmi
f+2sok/qZ8BfQfCfHFyI5znZZh7z61B28TiTyM2HZqUPTzFm75SyUne0I+MQ
CvCTSoz22IzMn+Xmkm17YPE+BGTK+fFUlMhpMfyoD+t04Nce/YcYIppxuvQm
zy2ZEv2GWYLOkzD3U5dLo9hDnGz5VYB6Lc93/I9UxFxHSoRXVyArquXVxtIJ
NfhYHUSNFNZj+L1BviChh+zLMdwhuffRIlYVJnccKmxLmXM1BH+Sv3vNRMyZ
gfgAqy+am1Q82PE1WAbzp6hWbBKbAiAxz7s9F+jgMKt18HLnFKVH17VCW1fh
MaqTe14yYK8QaBUb2RKDMzE3Udr/SthnTwKk6IvqZr32Tycw/RvviA0QjSDs
+at8dD1vgBwfz5Rr80Pm7rtkvdLVjOtgZT/ottWJNLOhtg1U49a32Iiuj88K
cEJKmcKHPkzxj5dMTkIvF7wSuabCrrUzV9FBLhaPVj8frGmgzkS+XptSjxOS
tVLbvBL6DeM6LYXtlysTx4KimHqY4Uw33e63AxosRcc4llQXIlr7/oS6gdkB
SsAi9V0MapFZTK5XAOIPvG4PnxaZa8sB8pgsWvQnH+mMgddU2zjKBE21HyFs
JRt7rQnCOdPfpb2HXLZaGge1Vidv3XOBwbTyGtqWLVdG+e4DJGYSkHunZJMQ
iccQ0vo+/m68i8fUWleRSULVWkXuj/6eX0lsmxxrWf06bZvp9E1tl7+8ZAKy
pO/IlT4F0+j4pSsJIxAyr5K0R/HKyS9D5EYpSURBI3QyiEj/UKaVlnl5wZ7k
KXCCWGIlr4NWse9WfY2ioApfvQFKrAaVUahtyvJFT+TSSbZny9JEdluSCDKW
z/Lr8RvaiWHMp7cN3vs+U3IKcWo97uXjya5jzmCbk9dT8ZVvzMzAFmTRnfKm
hv6JLh+wySZKSvZKoBpmCswQVEwzGrGztU5fs8V+gbwPkUAByFBfc4cNreEE
006qF/lrvBB4KEYzN8HWKso39Ip+VH6KyzrnE9aXwKofq4QftOKxN0mAi7k1
tOvr/TrGG1Rf8JlTd3JPNjEou2sdkqDKndSCZEko3/S5yEQCtHb+0m938z1Z
QOD1bYbiLvxG6ZzM8HKTK7nmGZvBqNM9ncmRLEHQsyKTOb7wWCeFqoHAZIC7
21GygmEXgK2nLjf6JW7HGaTzTHoa3gZC/l7HeA1gxCjkgFM3TSF2WXKZhAbe
FeoDXx5loU1nW+99Ib3W+uUPJCm9IrYKWpmkRaMDx08lgFxRqDmX2VPCrqIH
w5C/mb7W5o1vv3rmJDNdiu14Abu1Eki+BySK/4B+eUmgNnvgDJDr9+6zgl+N
cxY/JanIbCoBlT0+Tm21F8xrkpUV1rOiXxaYT3qkm6q7K6ADN45FjuLwxtgP
KF+nL+J/4i5GlCUdTgIWrfq4liOQ63LUNMKPyuwZ+e9kWRJ8otXUh5u70Gph
0btW+99VrQ9u7Ge3NqCfY+5nZOmafQr6vOiHaTWtIi2eJZ8ehd3viBnarWjI
EahjPU+lg9JTbJTbrvPj8lOw7MhtTbDHwG8zfFB1krciCPNhpqn+kHn0ywxd
JjZmP8/sfdi72nSzgE8lDtZ08097eUCZxO6/qLU+/lHRf6v47fChYWDx+CFb
C+c5G71x52DHsl1GbWDd9M4hNz9TUkkU+UbSuuKJ0hZi1cnxAQKSosdPz5uu
5BfbUul039UwVPCSw7czgFXpD05D6DgJCt3DoRhufkaxW3pgtgrRFesz1PMH
aiDnP2sGyi3I2XFzaqWFTdxGaV0SWWf5zT8Ij3LPPqyVg4Krj6Ll5++N3knG
LyM+cI7D+jRV0c8HvDkYR8mXVii/ZS9T3OBzv80Hpf8TjpQx4T2EkKW3+2ea
nKK0ylbYmUb9IiOOgl3OZTw3OU2sXGvP0WiNyjc7eAnbTk6Lkkw7Una8KJqk
POdv39A5n/1z1Btqp741ikkRH8I+LTnJx9qLW2UNO9glC7nOtXuJH7sBxlKt
5pE0mUf1/uSTmG9smWQ2b66A+BNWaMtYBk0mgLq8Zq6pBM8vff2NfUc2PIOu
VM96u6ufij1FYcX3Aaa8KQ8ki95pw5EF87/h3WeIxCjRF6JZABv/AexaCKa+
IH7JgOnJPmnu8Hkzd59Zv/SMEL82E6Q3VzVgIxACXl4LGIoKvH5v2W1gVODS
OqcWlc331c7DuU9i4mUoIkiiaCcDkcEpd2yOmBwwF5E609QuunNYsqJy3LcA
VRuqab2nl953hAAlh6vMaZoD+Y2TY6tVeHUqjsp2jNkkmt8u4Ofkg/K/XcF8
w5K6+oMd30awYyTt0rBP4h2r/jvuBV0yVPVs9/Ozuo/b/GQrimCZv0XsX0LM
5R/S7KgwnVtrpklSakvUL6ZlrK/vYNMylF9cXbNEqK/PbUxQIPNxWULPQHDM
TcHxghkaT0Fc/P8UtfmE47Pkz99TkluozDqxgxBsSBvCZPvZfhQWcyaJzasb
AlhxyTHMcbfXtzAsN8P6qUoInXlVgm0xKYtl6td8uSoT+1EciDu6ZVQq6Hoq
TWVZBjb8QJ1uixoqpSDPwhsr8Qgef+DwDyZb95AyxHYemzCjleea13KPXZs4
1OG7QvGpfsHwy0T76K4/BfvOyFdnCgG40bKObAXbbCa/dssGYNWFzBXf+CuF
+REriyesvTJ4bcNqoRqXLJ3lc6znXU1Z73zYl6F94HZmAJHhvCLDJmWB1+Z6
JEDT2im237J3ZzWHkwadqMCzUoYbqxhMlePGYM2ohJEb6BRD9CPX9etI8L8f
dhSQuXggyMQcQp7vdx5uAvFDnJJ2aC1NOEMir4hHyP6Ll0IINsgL6k+1u6oH
mYK0k9dbUfttvCbkQd4qdLPkt7Yn3OjoM8gN4OYsDhDR9O/kCfHe0q4FlOO2
xWahohmfK3WM+dKgjgVZZ1QjDETSZK6W0oAN1YZJuH6AqAi21nSEc2LySwWM
DxC+HVQC5IXy0dLikmUlsE0LIAuYVBheAP2tGNLISw0KPp2Z0th9tmsYv4DK
xd91aIUKPIvvarFj+WZ+sg/BOAG3mBqowNci0Uroz4sSyhn2aeSf3hmnVhp2
10W0RL/7YkXJ0IgPzXzuSRa92ocJde55l3g7CthtW+wjSc3FppCQOaZsInCb
KCukSsflAw0uvHPSrdKDvuFDAmW1dapL+PSIyN4MbilVpfL8jDgUU7xmzMgQ
oulXa8z/aKTjU4L9Rhhe8xc8TGdIZdZfkmFhmgo/IlU0kcz5aSX4i+MPC9F+
udVdt/9qxMJ1VZY6coy8RFLvNz42zuKsaPfmFlZzztyZN7ysN/o1QOfxARFL
GOSNBytiBiayx8CiC/RAQFK4xjq3aj3HtY6EiVkResV+/wu9qWaFUCuYj8/r
U3zF21i6bdM/GI+kUmI9h9zGQ6hmSHzMFPFjHQA3QTwSvMMiilyzJjNPdXH8
bDSX0csOMMQDyf8ZeSdsMb5Y46edMSuQv7yshJTeUvXfD5y8wzgsMF3rk/tt
KcdtIjR8tAPg3gLwCywAMPz6uEUS8NVJaxjIpjPNKL9UhvbecXJLP5FD+ASv
hvpzBzLoTYekiTGgxvo3lPs1niuyjF7ztUfE8poK3dxgvHeaoVmzXogK6MYp
Qp8o0sF3TuuQzCZdeecwqM6fdS3IhhvzIoj6ZDtpAgPsQTlqKo+jqF9t14Ac
iUnH26eJGa7KdRAAT5YGkVUVpXxmpaq20U3sxRNCoN08aMv4hWlCn8EVyIvX
+y+nC4xwCHdnUWzuCI4Azdc7gkUyrHxJ0ZiKnKXuHjjjiotPZ4FFCREvQ4mY
FyctFg7I99gshxchdXzyis06yFptNwqNUJFfGTANldpOISzFxtCEVYne9Sfp
LW9EdpLuoPLCL8DxmGmALZuBSwjpHqrQCY1wQvLSniHeiKcIn/fr9UXmumjv
9+yT7YQl2yH4/qTrB/xuko/MG22Xdws9Z1WZn824xYyks4AKXER1htVgAzoF
ZB1sCiQGvfMMKxHzebDOzRuYcjr8gCuoYgaJ+lEvmhrnDX0RUhCyqZ8d3mar
i93HQDedpNhvWZy+yzLl5hSyNTM7KlBKG7Jym7GKNDIRXjAH0k/7s2eiu2hB
XLmIGO12HFOupgcBtGlXzhyzDo2eyUvEYGZG3Ai9TDPhfGr75ExKxcX2BIbR
6zvvMSr58zR7lfffEEczIH71EpuFIfZ/gJcXo84js+gpZIp4faGUyrfgCxsM
tpQKxJnWXEEDZYUYoE2OVCKQ2ljrXZQzBtMEMpd8Cq3diqy3kTCigAFaDHnA
ICo0atjhXRsi0wwj8yyaq91HpqTrIgor+gYo+59g1MhBNdaL6doKMfYnG/mx
2Q2Y2uladnk7/InMdxlqWR1RKs+NitwEdVz5WORodXl7PHQOkNcFrHJFeZ95
SJLPuFIgXiNOSC3DEZ9YhMQvTlAACkF/ZWUpyi6SbSQWVmgYBlHzCgRoajhP
2i5Y1RJgfuRLMAGEaYsqLflQPxBaDsuqDe5Zr8M8igv/CrXbJpv0VHNHnuxT
FQsVv5at0dRACmkYCEQwHvn2FqgFNbCqVc3wrCDF0LQLxgp9HVozuj83yvqH
SJE2RE/dM3cR78mhXwh3DhyefTQojvAvXAK4cK6qIU1sl1clSlClZF8W/7W2
Z6+3UjgJNC8fe4VEV8reyuHF+RhJHgjflWdogtSg7XkS4Up5f+UXSgQxZJAh
S4b8zJ0UuMXGvtzPQEm2+3qbmy7poShykfeffgH7onjtsk83YCnEw49ytsp/
Uadf3dC+8lvkm5AQTAQ9vuQkB4niEqY0kb/+D5i9LqQ1LozKcxrR/Kie+pHK
tc24F64i1ii7OUQpI0empZVebh1c1mLqzv2dc0C6ZzGGzZSyfOm4ByPtTVVg
0+qKAGOWdN9ifJEZ+zg+Br2BZxlZumS8Q3A88pmBRX5CJEtJII80Gt66zce4
80WVJuoE5XFmh1sM3WWu602l4RAD9mtSa0/X8xeUOSd8hByS9bxW7UqQVR5/
cHC4zTcbToANHim762B722EhAgTMs6YhQ4yc4+c2q383s7druhhWZr/K6DoK
WUggfMMRYT7CmuMv/sH7odIf+kFnlLulrby3IvqV/AEo3ysN1MAYd9AXj7EC
WMdvv5XekoNAP6ZrJ0xAosr3r30kLf27i0CFotZ7F8gVeBlFRtYcSQ6IOH68
iEUq1JT1MKNkg6bgJj6BH1xnPetfuYcIBtmmAXwe0wWrsrerghlQquVyXwPu
jdTfS6vXlOM307QP3hq7Lgu5Olk9iV2ipybN5rQlY4kLvkvOrE9zPPheIWpP
Q7fIaT+9E6onsToRuUy82gMcs0EXl0E9gJ93A+opifddIjJPDwF+tf2lBoPD
yO01yN/j/wJGRjX7Hgyz9Mo6tJ7aw54EyBZCff9mGyTQbHfUWFVECvk8UlL2
E9ScHrwP08595Idz4vUSz/6PZTj6L6LQ6Z1IPI5PD5JTNxl2ab7EC0Erf0ap
eZg/2k4MbaMRlgaG0ROdrjHpRUVul+ACNIKKD3yuRyA7o7B8VyyNbw4C87O6
xWo6HePUB3ZInJbI7h0wfV0g43uUiJJeyCDLHpSUPnkaVa1mR7vujHJ5EM17
Hkil2b1lAV2ChWz74CJhq2XKS47OqduhKToWa02ML3ke8YyMheZuy88T6Hkv
6WKgEIRTUt6RN9WXHOvSMsUqDLs6sO4CSHuceHPnyS3lF12pDW6bsgFE79i7
tQxg2LQW2ZuSyt+nKDT8tbxmQZ1IdhyamU68qyGc0Zjx/hpcncUgyFr9ZwBo
X4uS2Qt+EMw+9ZiS/QLa94sXQI5hCdzRU4gBnhRphqT9l7/H9OCayviPTVpd
wGy7p9Y4tNVxt16d+yljEzbpVf0SxhcKnpLjrMkl5+FXcYPxfyq268bS1+Qo
OnSXzwhQtfxCeZxrffjXvKMxZrNxB51imvYwg2pm9PNtS6SnHOyrdNZbIxsx
qYeDPkYFhbR76/i6RwTOku/P+wpm1nVbA9KTGEhfGh46yBGW5UkuUTcj0kE0
akSECBo1hQ5887oGYWDRCg1KOhoTQqicooZpPEg+SyfpDZ3fa/rPFV1DdJii
BtDmjJCcxg6sVuKjGS/oZWBt2njTH2g8znUbIJy4z1PqN5/JGF9zavzUXmum
hhJ+9oz4BVyNYpsSnZsy9u6NRscTwjejtIjypApwu1oi0oP5MzP1N+nYHs14
0CUdQFp+5c4QQXW9v1r+UH+dSNBgZtHdqk8LTrCePhD5mYfYLl2xRGu+ER07
CjYdJIxLQqeUDtgq/qschF2EteORakIoEEg8/CAeRn/GKlcVYA6L0A6DgpzH
2l2JXe85cmG5m+g0Aj2bhBusLQGOBWfeTD95atpWXYifdlz/kh33pGLg0LNW
XAjnx4B28S2rnSpH3mSGGpZgkScAURTqkakWaeBAcun2FKTI7B9SQzxmsdU1
8C5dHMjuKBcsjp4ZizcmKtzlCQ6KKPAWLZ10XbEAGhMNJV3dwXVlrQxuRQFG
iz/KSaH4n7j6lvBKsdtqiwEZXVxkdjkPUVbhldZYl8SqDZzXB/OeV7q0avU8
A1ayrBbqDitohvXX+NQ6oyxeeXWwCrEWM+zYamnvJXExf2NTITexG0KfNm0r
t/1fQXxxDvKh7fzxW1kBSiPQJvagSj84jw/fSBTMj4kcWVwCtLZj0AK9bxn+
hZmUcUMsk6Rh/faMQIUZKHegPbgQMMOR/5gS8AwIA9Az+Ob3wuKj94lorfzB
NoBGkn8uFH7Eh7hkJAIiVUG6pyDLyRxEP7DemIvo8TixDrQLqc0qNStuUl5Y
NCV5EB2WjBizKXierV+dYooeNc4A7ine4z6j8laaeB9mQfisUL4eSlW4lee6
MmFPGZ4zg6Nkonm9ww84itk+5sspVprmrmRdWzFI+x9lskvv90btewI9DQ+9
OPnqxDrUT1iV5XDxRSHdoo3bSHZmZ4/soqFRO6JsUBkWoH7V6VI3bSe5mdpi
tM67MuotdgG8P8cMS8ZQ0faW6ywE48+6ctSvCi9VoOO0S90FKU3myFRk+zYY
7ZeinoYazfIqbqyUuLxLQnLU9FzlzOMMRW8tQLG3CZhG66GAGWqGvHrfyO5h
zjtlhoutTZ76ujLJnJ2XPHQaictJGDQR4P9+XyACjoHJ0AQRmmW5HYSIX1YF
UMqH2vYiqjs4qJzmNH1qstFAsAiP06JcjWp12zwriFEDgy/McdLreNima3F8
g7mOBmh4Mzhg46e19D2Sg1X1sMyzx65GlM6TCbHKYX5YXahM/kCuUAbBh6WS
T1Fl/qKMnuL1W3Mt3gCGMrh+a4HeWR4LN5GDYZCQwcWZFqEsS1+SXhFo45XM
1QDfRPprauC3aPZSx+NT7BRAQYHIyC4V/bvub5xM8v3GTiDW2FTiByo65GJr
y9OT5vpqHZCsK1uEZYhNQXADtLt+w/Oq2dTL9cv3M5uZ8umtWgQ+DXQ4etDZ
y7VCCgIm5oQR7Rb4r14k23LIZkGxWLjEmEQqF5iHUgose1oOgofp+kY0XZYw
M0NxLpBV8VolaJOxCuGWVnMJf9N2utdEJtJ5RRqszKqPb/Lfnd6O/CCbqRIy
w3Wyl7LpCnO7UVtqQU1ldjzsHmhNULolEoGr1ZWiQ7i+wm3wSp9TZyeMyEKh
/Qgadl13P33OgGXw/Sz7WgwXH7jxtUyafnIpY161dXH7KKdfX2BqHraMr3kB
x2qshi3lIVXIjwRy782gAEANvhou3cvN88bx/iV8V+UlNSltxKUVUuQvmvS9
EFjQnNMLJU3PUs2cXBEOYHr0F0aEiWGE6YfUOh5MrBvOUghWsk/ZLj2LpUGT
GjjSHtIqSwyGqORoWufozr46SwmIPi/j9dg8o+g4Jx7Bow4pCWTBftQA2aqx
wwzC5b5LP4u5jzN5y95b4IqYptqxGB16dMDZrxbX7ppZ16vdY81N3rKEq/E/
6ezLbZAOdxEamt8vCCFuQBv3iVskhac+OXbl4SydyRwwzwBcbh/zoUiUywuM
zlItKljrCqnusdTYSbwkqTi7kzLnLl7srLaTBZQdf2DEBjMBna69NGY0SPKW
mcjFT6YhHO+uBWh4ACoam0I8qV/W6A1h4iPryBJX1TSAAUVsgMs6scxNJjoY
twYADTm/mZeGCyhxx3/JGhUtvoEKY/tbOg8IlAAh3XAaV25RN6+cpdrJ+zw6
l2tc0FINY43i72aKWXEKFOC86a0B3Ib3BpY6JrRQ9dm/aqMeXs+aIw/DnC02
uS16wo4UP8qqKZMo1axIc4+a71PEFhMKRUl3U1ZAzl4rqM2pUr/BRIMMDpXm
Rk2OAA1y0xGTcb3gL1efkbERpf6U6WG9+SAWgs06d5jygXcN9k3oWJrvffHV
rX3mZaCDup4YZOzbM0iJS6FwoheZXK+RN/4NLdiAtRdn0Cfyc0OEVx90T7Os
cKbJVnQu6UDJzFZyHadsoz4bfY/zh21bXE3dKF6ubmY8V58b4Qr6aTtaHnbk
gl+V7/Hw42Mi1Mm5KG/gbDZURtshf9iNSVafRElxZWjPa4fXEIcBVaXSaO39
pwAx9NZGPyGKwRTQxzxZ6Rea6kzeFB8qooyWTLiqSzG0yCb/9x9hM44REkWi
JMsKar8ph0G3lHYFoRHjWDH26pdr67AhMvXNvwzlbDDkPJ5y05Xy4SM1xYLF
4S4O6FTTo5/SBy7rqKvL8qriueUdZtf8obJGhvEIfyqJ1ZBsGv6egt0rApsC
LT3c2NCNmn130IbenXWEUeJEGGiXB23fg9b1r6xnKvdEDTt0ewLPoqGe2y8a
xxh2FBX+dcLWpZGxS/ix+kyKMI4+ZXEt4Wy7WVyjZ0Vz+nfjwIzGep4A+Wnt
JgMaIcofvi5btn3er6rHqhsiUOvCEmx2WFl5ydSp+Fmfs3HKZrVmoC/St9+Z
r7/PQa37TIheTu8Hv1SLusEx+ZgOFvQTZ1SAsZai7FhGwbzYmSxx7s97/s2Q
3symAm5eLXGITIYtdZZTJaL28BOEuGoZNPHSSf0W1VBsXKNN62zXl/AUJUYL
ySdduTXjXGNY5xSoa9V+MJfCnLiWbJFhQheGwhfQbNXQ9pxfsD1ijMRlrbgF
QH55Nd1zUBOaX4tds0Ti/RFCGGdV4XTISpJQqWS5Ed+ap1ypvMT+qyjwd2x+
0WX+MWPqbfQutYx1HMsGzmjphyGhfCriXzEq6Pn2wBOEBdq45WDSoHkESCt/
dlKywIYUn/z9zDzuOGinQUNQAQox9OkupYSyBn2eOILQWvIXSgqML/1BdgGT
9VnIkU0mcZ2bVhHudDykqLJLFXSwBGNo83jtxWmsU5Kex6UImUl49Bsn92rL
tlSk84o5fQo9bb2kfRUsSuvwOuJhhetQX+Jaf6zswirhFvqZ04nM+pHSEs3A
G42ZEqP02MbPUku4snVLbnnSOdY+lJw1aMKUYUuaut/r0QBdX+b87C64jerd
qxKD1n1YK/mCFMxp+i/R5H5k8NhbAMIZXUeh8iWTKR6Wobh+f4hPGuuaXH5a
qLPz2NL9zmz7ADNEHP/aD63FBytDyw53C7WtfU31vNcsEM+ivdtLECksnDbK
SsTAmpoMqC5YwObUdt9o7al9vFeDHQ9j9ytXGkNSKZ1uDshxG2t/JIBOkc0P
RYLGas93u/bNjHizPyD6sy04bWfgNKIdYIeccI3Iwt9ggKp7/zAdRDkab+sC
uRON9GtlaoGEoWjA4Uz9nhHgB5+Oz+kLgQLWRYlBhhR2iu3f3NHfPr1bOoJ5
qtilyuvv3JV2sgVJjWuKm8NZ03EuuhiggfRTmpqnEZSJqqCK7pc0K7/1E0Wm
g5bV3OKzEcWY+WIk7VA6oM45VxMQLhixx6ds33XXU95DXFYgtSlW8NJw6n7x
gQJbt110W5c6KiSKWuiYTzaOr6qbw3nmWHthaX/LUXddT4TM+HM6NOQcdJFX
qM7Hgln/uhTHz0PLSqCdX2oH+9LLNJZmxKosUEbYTHwHIeYaeW9v3pF/bB/T
gHkKUVlUIRHxrgI5dN2hBEvJkVfvDxoZi7G5iJC2LCfQm02/xdBR4XvmRAU0
J9JPxW77/03vM4Eeo09faXT8/iBDML59u64G1AnnGr81rDKzDhT7BeUZRpCB
cqPABf0vsC0eFTH/5pu3c2g+5Cyu/yCOMqL1cSFZec49itbJuEHj9pSrs55G
kWT5gElF/AXF6JB8WvFc7/R1BaXPYaMSOiD69J3AZkpkXMcAV8bi8G+SOao7
j9tBDDRb8PAdWIqLAdEeWjJB6zNKwwvpsNFLSKLHBouWTwSvFcIm5dtGADDL
5zxrIlgUNmHGn2W875CJi8CDxquJU5vM2Q8W1Z2fjLnnffeTGsLpAhK+CMS0
BKPUo2OAawV1O4BsPQ9P1TmOPg/LDPUI/M3tNoV2LDuZoq0bktyttxWbWsTz
YdrmEBbTo9KmGOLLvoLaELl5NHwq1FcD+K1sgtGyoDE1F2TtnkGlziCjOioc
in0M0SRI49PihuFk8ah2PNeJrB/uN99RO8EIakUmrf1/YFQ88T3Wz2DfBpq8
7pEh/DgUvUnXzK4e5POIdCEjoMslH5f0QxKgyMkpiiVTcL8Dlf83MWP3GRSK
hARPuT8X6QkFyknyoljWHxqKTB01AveJ6d/jRVNkWQqDHVXFoRxUFC2S8sC6
DqeJM2PFzOZsKPYhinQoA+IZ79lum2Me5hDt5Q5w6Hrud5I9pYuBjleAJp5y
EnSHV6T0cvBFssLJhg6YzQ+/FlVaIqh0PQbnBEkyfqqChJQYm3xe+1MSCpCd
ozrjs4kS7e4LSQJvsOt03xGdXkFoQSjAgc88jM2BtM3tXddf/U/njIYJnypa
kpOgaCWH8Bk/sFQ3BCSEqMXdiGHlMCMfw0YYarKEKNynW2lKOJc7IpZCk99f
1Sw1uMje7UsXJHJ88W4cbR18VihNhFiGzxkskBtSxIft/6FcWr5Iz4akonqp
YfnpWfDWSZmBlJ/rqQZp2a6aUddHhWfM65iQjIfW99yE1jSnsTLf1AmT9K3a
r6RzNkqCsmVWvOEEYwl4fQf3mmtHD79JP0mwHu5NZ0Sd7+q/i++OECff/2tc
W/Rwlx2mnOxoT9xatf5utaqFb303lFahxKJ4PK0hiQvYBZCQy732rS98ByD8
UIPk53Dk3vqb+N4wIZR7k5CGhY3EhDXnMTA6Z16ErE0CwPfaj/bnsoZwZ70D
MKCGFjMbWvPaXqK0kGXsvKM3o84YfYs4ii3Jsj6+BuFTcd/A/jSGwSVGk4aU
ETIBkQwt590OtiolY364zLqIiyIqxUvcnOixyDfRy9bENumNCf0K1MtP6KvC
AnlG9XFUhKNruo+9UtfV8juEJhkHTQmdtKsJFq9+pNcpHlQ7UkOrTVzH5A10
HnzPdALlCG6yDTaTQIVf9+aVutWfZ0CE7NoPV9MEPAD1uSm88672KwkouPKL
Clf3HHIj2sOO/XLyN0Gx7FlDIWy6CBZMew6bNRb0YmJseETDsZQrnDXfKFbX
SR2bar1dbSbQfKJv5I+5OsjMC7VdmIhlEPkeTFWSYb6Wrmno70zyFN1d40Oq
MTLRghAR3mrcTODDvywi0+B1AZfpOFn/ihPqV3ZMlfii9sz/KdPc5WBnPGo2
uETzD54LeXe3sLYXKF1xKIDQ/2h/CDvxtOhZMGkm6A+cadTdHnYgJt0DEoLh
p3GYBYPhE8XyNh5ughYy9SgV8/TXfFdF7CqPMi+RMYM9f2FhyZr5gxoPKxtO
UugHjTWVYnKVFh6IKreUA7o7zLl/d1VycP2Qez3uV0tswYNqsTELyepGjOt1
QpMm0g2olLiaH/6MWvO5tYNINoJXEvqftJ6ofKZrSxOHIPCbXU+jxKV6urNy
4ESstHenQ7HBGTf+3scb/lyBx8Q+FTjbGX2nO9Z7nj3Qgi9hwSTqOMH/xiBO
PqqMpeRkjvRdv25psnx7vWoIJPRFxaLNK2MHwcfyx9udJnE5BNRArUTo2sB+
lWsPKZPVFKur+AZSHWRtPwpfFciuvNvXJZwdzdoSdNinlxZHECi7+Dyd3Fnt
3r31UyRMa/+QxxjNFlKbhw78f5EsAvHglgODVaSAl8sW2zAxycx6N/8wCyQl
mDMJggdQyth2DttWURNPiyCO4tA8xrNZfyujPlpGxCrUWIESwvrAcjlZRUdy
BsU7vUTEOn8xiaDRIKH/7AOWg4oIdJSjGgj016dF/Y3FgOrqk+wRcV/U/MAV
qw88P8YWlU+xj+D6nB50R7KE7ud9fOsM1HhIka5eCHMQCjs+umN7JXXouVMH
1jdBrak+YwkMwLkF3KKJEOnNbuGU1PhVfwJHIU7Zf6Na8ERzKKnsw6dkxF4A
2dZTXxrTcSVhCZ0ektC2qzWv/Cgv1/eHH/lVWhv8LTJUSjyanhjb+MYCLUQ8
txFJc8XI+mIr2GgpbWZU0GZiAjLVPI01b41mGmZ9I3OdLF0W8u2LBURDtZA9
m9nFEdNOAzk+H0KT80x6V23WtLsTsBUdyGxvBJqb1fgeb0c6ofAGcqG+Fm1m
C27kvEFo6WT3V0CqG8/YM3yn7TJ/bVS6CgMCb7PbuIyphOiutShHQ5Zg3HaZ
a2RWzhn3EDV8JwYO7pLI62+1it6G6Lu1ic1qKozDnqBpUHYMU/NSLt7y8u0+
MZlmTv0SyAa+GrRwk2wQn/hrAD34tbqtuKrJnAB4eJgvMYe6Zmpk9PhhC0hX
+v/TU9BYshFczTpcDdCzAxx669vfgwxbfdv70FDTsedQn+vYY65y3h5VS3Ex
TGWfCF6Ao3qqIVR6EJYKg9A69IbhL7LpsZBzog0aKm8TjsfGTq6YWAXQVovJ
yqg1juY1wMs+eBh8pW9FWsXXkv9kd/lKNn0MYYJEhi8KhxoVwZmbzMDiQNYZ
BZH1lfx563UnYGVEUEi3aWu9CLclde9dwYW2t3lnnb/VAWJ4+Dvc0tXlW/pn
MaW0TtgW8ijV6Olt6GOtPBa7z2p+/SwZkQ+bo6HEIl2GaqP8ernaha4L0gvB
zWd6WoonqJuxK++hpv/7yexGZeCj0cr/MOV9JF68uK5tfRLzZ95/Mkt+TkEO
jkpesps/y9VAFuJ6XRDipYfCGXrRYjHI81q+LROW/bPWBI0yQQ6GK0jZXTtl
1IebvQSIxftyR4itL78DlZnYCmT5sZfDDIjz8Nu5/k9xkL2O2vZWbcLrka6p
iRS0++SU2V6nFbYcKG7mgZh0wsyPGWciIPSeYB8H/lTXkoOiOKGShgyWYTqy
lL87nRmeya6AnSauA8qtnXlNk2McpZxc11nv3NpJ9Q3t2UH9orjJ5IaZT/4/
DwevZ2aOCjXlbLFsge00ysi44WsW8giWaapUrWyK3r7xY539PebIhwv/L7Mv
8b+R75aSNBqdeyCta/k710gsTdv5egI8tp3V4HlmpVnZ5nst8fK2NuRtCf9Q
LAgB9UIA42C/i6l+T7Z1lTl2b8LThhw1Fh2rH6fLd8THGImetELGDQV7Foeo
NV5DFkDdlUjX065MczcnbE6iJ7K1/a+AEB52r92fmvx6XmAu+NtPRwDFZtyu
D1BoEaSShlq0zKX9Za3R00kB3S/hYfqaIBqLXl579rijlZMKS+kSjxBCnwre
ElRuIhX84Z0E9rIC6yH6vgo5/I0RE10cFFfByKqJ3THJtfVKQ9nH5CyhiIpF
LzmyB8mtc1dp0rTzRNiVvKvCRt5gJnkerg2j6jmJws4UMeQsFp0R70noPImY
dqvp5SK7g+Adsl8aF/PSQGvt1O5ViRoyb9Xq6KrLh+jbEtbBOhpw75SBiDW+
ik/Zzpv9yxcN2uUkEbx99A+BAcsiiRQZpkIB38pc2Ud3C9VMFJQRYqygQGC7
QNqdcu8m9Td8SCzXT0U0p0RzF4ccUi/X2jOeVIjxSG85GmRYW1nDsWsMiHA/
7VIPKO1jZrzj1JwPS5OMTCf+jDvgP6KTlEQetTmEIuLx9nyU1OQbyW3I80yZ
rJ9veYKgekz/qAVs2OaG0SWngDCBSczkdo2PPkzIsxPcgeHmVguvGytIgSfU
7HBz09A7obyjSx4+9c80scrulN6i73VjFnUKYvGCVIGjszx7/0Z+7xM9w+NH
qHANO4KtgAbFaZ70qsN/ZE4z/7mQ+mKizsfn3yXLoagi0DKhoU1XIDw1enrb
VMoqrPHgxVvgGjbIJ2ytb4QyjAfrg83xm3GkJpyR/Zu+vaMLHbvlA76ik7gM
3A6p0l6JtmRVFaUO9zIwW3M9aqZVaQF3m4+pD0wTg1tFL1hSXHdx8wHkwF//
SwTOdH/26BnnNeus24ACN9mHge7sO5SowsXHBnkEgncniEKbc8VUC8ybQx9B
XU4WR131iIfCOIz6fObsJsoQ7iWDChGS9O4o+6NJGDphWBexOAdE5u2Echir
vaOpRXvN3adnpT+aIngwoFgmku7AQGGSdE/3LXKCBi1J5igfWtSoC+U+Akef
sRkOvVmHFoBDXoaE5NsjgNnsjk28vGr3VRe87B2yGLL7uYzeGEkElSGcVOrZ
Y74oIpkmb4gonNPZnhDR5TneeUOznwgB4CLq9nxIxjP3fIKQskh1IxkHVrEJ
7uI9h8mtNYKlZQbRA6ovjG/QJLJJhaylmhAA2ZYPkwpGbxr8tb9Cr4SWDHcv
3fRPZD5PlEPs+N/LDuMstzwiSy9ffOLYNhgVuc1lKvMkpZfhSCiR7TH3va7N
T27Nwh1Dx2iWpdapmM/myeLCZI1XKnOQcKkdPSa0vkc1h1X2NJK1AErA2okE
n8dstcyfeUQ0kkG7CKh2iE3KjNaVxMJWJATzxNBtFDCMPX8l6VxN1SaxXdEl
KLyLuGqSKbW8M64bEOGV2LQ56bBEfIuDGoJSW/sfroECPCmafkOOMvVCqvpe
iCQ+F/gyks6IQh++7faiQ0VPsNRTnaqto66jDnY9polqBQzzzxUs2HwUyr/W
cifm1c+nRLMTpbgIonq29jyyFFO28BGQxSXTKbvUg89HOmT9XN7LcQNG+icl
+To7UpDDZ29SrJLYpRhtQzO0Vo6JGlshhA1+bVwjwayAE+b4OHTGPEFANq7B
AttDe4ETaXq/iYsbVkTYqOZUFkjsMjk5QZNwUaMC69cjC9ug/diu3ApM4i0Y
KFlvTJldKeywItmdJPSTwLc8of9OqjJhJL2q4MavlRKzdh5blrOLJ7aZHziP
Gtp7GvSbV5QDLKC6HfyyfVM/TZMvsI+J1HR2ZXCjd/S4/QL8NgqeIM60TnQT
Jw19WgTUA6KxNJt5e0mpmFyw066k+DGQFTh/tw+uYwue9i1MPVF/zoyZcoz5
MU43EKRTC0GSaGb4oQ7kmy+Bea58Vh/jJDdkufugLxL07cqGlGm+Gc7SP5Kj
ZEDFpn00NgJWvWbzKhl3n5nENgM+Rpec8x+WxZDFi0s/tRtT+Gy25OiKojsE
pv/vYz7pacF5XuLWp12rS54zoPOM2N8VVmATFijsXhdsprA2KrbDacyCj6jr
Luj8Kg04C2pXF9AwcWgfCUUFZzOnQBVdDzgMYUQhIwaCdOtNFDmnuq4QyslQ
q6NFswcG4sYQnGytKQdeUR8i6UrrbEjE543hJir3y92JPW0bjiNJ854b56xM
uAslssEl9cWKdPsY6mZy+xJsQdCKGKoJ4Dp7H2v10tRXP60A51eSSV86qUwQ
dTu7SBgqtZHllMVvpQUV+yotxJBJTCgavxqfKHcz19o5t8pQ9/4cD68sfb9R
CBcNcMCjhzgNBY59fXnfLEn+kbHHHISJm1uZRheM7Yi80FKfowDFSOj+0OTa
n4wq+6M6NUL0bvDPdc8uoLVBuJqtMasgmHzYT0XeNO4WTVSYyU373uEHbvyj
94zlEaynBbfhsKJFzCOZPy+JYjTQqX+w/ld2DTSD9V/Np8IieuUzSWjBbZPI
W7pjkA8PojSWG/ALZukCum8vSPhQul1C1+p+b1MB/LPTsSdtNh/YaR6RVKaW
VO2dgCuEgRDxwhfnTj1oyZw+r5mzLvC3wmexG/qKFzJqp0LArRtfwHndyli8
rDYmD2WxQke/IP/kovuJLKzDVb4W/KSShEx92+STFB+Va986zzejAGc5p+pA
Ek/2KGQZHo85jiFKM4XvshgdDJ5PPSZlbR51xqclmdc0OZMkASNjCiblWLAb
5GWF62IW75wwvO8Uh62Wb/h5bVDKw7KjAioJocHuQpza3TEigud4KuPrOtf3
b4XJ60hqLgGuDE1OSk8YhAq2GXPGty7Wtpidi/hxRkK3OsoRnxCy+QnJ0ljp
0jkqDsfzC9Fkg7kYvBirObSV0BW+F84SkHdzYh0YkzDzXR3gmRBR9dkYHa4D
9e+twjzMeGp7MpoPBLI2NCZURTQDgfIfj9STFfLaufG89SvylREdtrnEzzEv
/4UA2ZTRcLvTZxsTDabOVAJqbtwhcoIfd0DL+notYU+FkiulMoywpcAOtu72
SeB0Vrb0RQsTLRtnDhwN6ftzCKZvKMs1hc/NWnm7QubW9OBsrz+n51ONP1hR
yuWwlaO8HXX4qJsADr17aSdQX9lI/alQI0XBD8eCFvr7aAGjC2JZ3ejYBRjC
I5sT4/KV7HetirQ/S0pm0chaU3tf2ZSJWQ2woale438iuUVR3u2+Cf2H4TFW
2MDukmOB3cdOFhWkl4Vshh1CmTKhH444y1KE6ovZ/qe+2ShRNkjtxcTM/iCp
0Ft7fz9WYsvv1tHN8L7bLYgN7QSZ+S8g5SDHr00QV2YslPXMAoWycpnmAvAA
yyhDFUHiQawyKalFot9p+VY3slW7BS1NsAZWZ+ehAZIQTBlqK2MjLTAv5mh9
mIBlBCFJzifhHXj4XueipgE1bnA50phPbY/7WNHXklEowdtj6HeRPQqPw2Vg
NbYHNzJdWcjo4H4b/jFWPJo9HOvSfXf0zj+h1uH6X0BChQs6xuX7ZYOtFKki
VEPJEZi9hkmn8sY/8TRKFV7Vg7c+RdpygV6RaIFVMmS1oQpsbJnqE08kGe0Y
UFvLYD215pRpLvVZB7WJfB2CxOHcG1n4dRTrxKx20LvFsH5oNcTJ5dwN4qKk
CjxfTxB/qKgiuQgJhq1V7/MSStvl4zjdyXw3Y5ABn0QpfA/VQG74jCnHGrNy
57jctpfVxrWc4sKkNlaZ8hYpn/j5gIwTMWe0SVHk+6/yqYSSKVvWSeO83ZwO
F2CXurVjnAeJ1D/BsEVokv3OcELzav0D5jJqMADeoyEYoKTx7R7JI0Xa2kbT
6A3z5kQ5UPr4ZmZ3SdbcpV741+UTWgJHp4IndWmYH2YP+hPNyIhKcYsiQsuv
RQpzQjmdxnhxXiLTmw/T13dtLaKEeFSzJPCSDfhvatwQfpX28NH+Tv//zBEP
50bvocXkc/BW5yGXoWcl5g8ncgdkc4ocHKhxFNeES+fUeVQ0bsG4LNTQ4DFD
cqQeIAoNEDVbHNHgcCS+kQf8/4hmXcfpFO+k+lsDjBUUoKNWe7Bj6itxXMvq
lMp1fkMqUxS+U49JQjufLmTqDy1pqja/ZPp02B0Ogtd8q04uOl9VYsy+0Xkb
i337erE75hAO2oxXLxD4994iT5bF+B3GRig4cH70PKboJo0polEAeICiZcU8
cmeM5jgCWNtCGzW56SK8ZvG3VzgNALB8g8sNhDabHKbcbSMkn7p2vHdRuisA
NHSoiyU+X5dTMXjVprjmCw/weDTiRVwNvkfiwbgt9rmOo4kyoWoLSKURUGHY
ERKo1wW2Wk3j8Zq7WfszUQjAuemwwr/ktTVdshdUhPIxiic/TAtrkCS2xHkw
t0PFmgQu59wCiQ0Is+Gx4BxOiKytK3Z5kVmL2wm83p/ksyOahBTIo6Fw+FWC
1wUZeQldwlggTK1KzVAZfspuw6q7vmdQjPjR4NYjRtuAR/GbEFznWfkZNs10
sdS02vzSeh4QvslDJwhO1mi2KfNRJWNCWXR8I4vvKmAEXNk/+1rOCn/Dw4Yp
v1nOFugaB+qNXzjxzmEnQMynu6rKFp/CTCYtFtlrTlG/874oQ948QCISzeSG
YNiLtt7DfYEdEacBOWW9cV1MVIMEz5aanOglqA/cSOqPujrpAjYLTsRFL9LY
Tey6vtg7z7R/3fsgQ4rTsuV/b5j0QMpghsHSyVj056cCQMJtUuyHHa36pRsI
hRdn+Dm9WzjTtBULRvNTd7GGMeDFAHeTtuRrGUdX+lqXOc+d05T7vLXnHsHD
b0KUbKZYPBx4c8Bm8kbTj1dOmpjATE0dUFGfn3yZjL6suNdPjtME98Jap1a3
M8n8mpRCKphFpv8f/mKSkQtAiks1mD0VVtkTx4hlRd8ews7DBGe55sa1axlx
25k6C7v17EH+pULtA0Joq/Zbt5ybnM/vRlqqd2dZgoHlnJl7AxBcJgSb35uu
VvcQni/wwcMgbvyrECbXHUBy2jCPDeh1A7naEzF+pM5HT04tUVwUiEEQ8z0d
q/OxJau85ippeGIessS+lXHBiGvEnn6kaC8zEMsX/IQvgYCenjHZGMvApHpz
vOSkcMnHzcOV3R6KNUPKyK0lEwB41luCWEiBM1k0hvfYu2/Y+8WxZNXKlNIb
3rynI0YfKOgMCy5RueYaRYEvJOM2Qhl+BaEWF5cvm3TnDXcjvA2lsPUZtmvA
aMTPbtl8RSIWgeR78yJ9wAVa0MgTZebpJDZc5gL7hrQyhRmA7pKbtOKLT/cH
o4s7JAI0OTRsuutAdnlQQwmquymxplEen6qDC9gJqe0FSZkOyqaDLRvJQI4G
ms+sg1iOLFxKK+fWFz8eGvdf5KqZNz1PHybw0U3rGQ7TFePIvpCBELBv/sxa
QXd3/Ydz9BUYYxcFiGAMoVFiERl6K0KTnqxvwxcmHuIlZAcIM2T2Ay7JmWdo
MCG2kj6oc8ClwFjzOh05KeQI6x6UObI2K+VpC1CWRfuYnr3V4JP1Mbzp0Agh
Vi0FRCiJX8NPKZLDMun6O6xv9ws6UX5zY4JOx9RaeQ8D+MTsKcuWc/+v3spT
OY+YOuBT9MSzkJaSGnrETZei3q40gcFlV4mo5SiXWP+E+r1ymg6P2ztC5srD
exufDUF32iuRFxw1TB6yNmJtP/kepPRjV5YKZDed50B1Br/h18vzDadyo7DI
S3OiJBIdt/FBHkjiHlRUd8HO5T/zewl9rrgiUe82s0lnGON+C2OdNt2VTqLq
WYQ6gQ7BvyrfvZx/I4GduW9EWduGLZXUB7C+AbqH/PQmhWcJZpx/58OuGpbe
qiiXQSCxLNLd5TwAH0+T7FAdtvo4MgD1ZXQEeJm7nAm3lRLQm2r5586q7Dcb
sFXEZamiXX4Ob20LA+lTVM1cNMjO4LHUfmA1nM6LB+lE4sO/Im3C/M3RoOEM
GB6AbEMe+12Wyw4ggkYzQ5PqeKu44s3iZMunUhShFKxBxM0gaTK0TkTmqkZi
fcIQ6rr2iCjSQOaUqaHvc6pr/wp19aOyNQnIa96wtstIYT0UIQo2RnS5/Olc
piwHQHDUSPEtmcGdE84bVS2s5f2+SIh1utDKd+Q1hCAVMFZYkjK6S/3T/OAu
HLQP0D/lfR4Mjw6N0an6ersj5r8iYXWe97Q6Dztfvg4CY7HSy/tfswh6zBpM
mLnXw3QtlGW7Oncjl94g/wKzgVdt179pclGuPqloJKJ7b4hXFA+VXeGifH06
Ik8w1JlYsvrfY3yvmeq8N04Ok6Mh6A0eFF98FH1ZCumwe2lEG3xEojo+uamm
jlr0hhDMWGDNhuzvSTl99V2ldS3vp8oQzJpQo17BMTAIbDPMkNTIe0VOovEa
6N2i6UpO00P/UsX6hPRrfI1hXUvnqD+/rr1Q0KAee6+3GoKzCFQLPjxRuYGa
DqnGwSHxJiHNgItOYtFhVQ2TbKnouYqO1deL1fgQ0t5ViEPUEJB/HVr4KdI4
1XGQi4VoB3SlXNm8XRk+cC3xD9tGiiKpYyBt119PS9ciR13/0ey/EnU773KK
g3jIbSFgqcn5uCMLh/WgRtogNuhpkWX17hzEiyLJSDWgFU16jhc2J7orBLCr
q3AsJNNEbQZ0dpSbrL0GxAdV+TXSHN4Qkdc/0HmNeoJuO38zkiw+z9brrfee
weLYqgPXtSSuPuyf6q0y6/8HZKSC9uF7FywahPUWTpvfLnubPenYHPqommRR
QHSXxTPL/wzERYE7giXC/IwJ2StwLTynfoshrd/AyYHjjL/1zErR2/GNut9c
E0yRUiNu+JYR9H8WJRxW7kgwzq/Wt667NWkpBcKxyNt9g1MhdTEda9rKtxsW
A/x2WoO+fOswTyXbgIr7u1TLaiTMgpg+p3b24v3yspy4LeITusA1nhq5zDA2
6pSE6SDMejqMcZDdSa1Fl/lDCFcMDcTfeaejmKcekASGJrqQDydnuYikWlKi
SQYZYtUTOdgmh7zt7PwE9L+GoV9NhNFDcCbw0izmgKUP5iw8wO2OBW1zz7Tz
gBjCKvvkSN1l75yiFaSdIVrksXS2c/8wCSsVDQuVBHu/lENn2GeKUbRyvoTR
l9oNRqFXapG1vljN5QYBf5hMz0DZrOE256fG9g90z94ABk/nDQ7WuA/95r8e
u2fZnfHNoYJF6Fyk5eNUU72Tfg1YL7WZI8n01/Auwz2NB3fQ8kuj8qjgC2O2
3u8KBrsUd2F74HkA9iTPqeuIs7NZOoPpqqINxFsbHBg6MSFKDMEWV74wkBH3
z/O93zr71PVbHrIN6HmQ7HOw1IEvqi4Egoqm2krPkqUahpLLZ0YqQ8yUrSVN
KAgZh9OixUuFimegjsHdXO7QFGRyI4QV1cGHeXxGsBPJu9fD3O0gXOMVnB9Z
jiVpgVarc4q9dVGtorJlTqzFdVQhcNvrnrrGj72hL23nqpCKu/ByJJ3DIgMl
zTHnVTqCIKRpUGeMO4XMyc65NTqLUiKYu5NxiHsfFzFkDANvDlkLVP6Lo5tA
UP/ewqLA+AC7R7ZFNueCFiRKIe6kr6f2+8JZ8VWK/UwstjrTKd418EA2adtW
4oP8ndES1CWz6nQ38jsjGsz6uLVuMgiqAAyZFzRrmpkjP6qMUM0s/1yZgVgp
HYq4d7WRFUNzKajTpXea6yH/hWaQw/6vpaSyFSyyUoK/+24cfAbi5RsHkbXV
rqxYto2DsjXClPH/NvTzF/9SYtYXO5IkpseBLIbTI9KMjPigvwYVfZ9cYXsT
LPND9TI/9bZsnmdwQgtfdd9mvlIEagOTzcWYv1VVZRhAJTgspZ92kTg7moNI
d8bDyS8SPPtJRX0i7bf9ZqsCE7suuyRIj7NilvU3yHpXRxITMAJje7ibb0Ss
OrZiTEHLTWQCPYdP2bvCvLhHVT+RjtHoGVypiRB6c/9kHYLx20C31gvI1sh1
1yl4BtCcVMbrKUQGbAwvepsWIZDU+EVpSdlKrKw0evyAqQm6ighgC12HXGJj
kr9IQTTgQ87ADvPAIqvpfkt5qxyys7nfnGHVmA6zIWODSZardQb6CwxOf0R0
TdbBDNmo/7jwcaSiGFS/GjPR1dwRzbPQn/bboVvSkeuisJ86r+WweKVY4Ze/
uKE138ghBpq/YPX8rpvyhFQ7d4rlU+aZOaXCz4hx1QBUK23EgLHnHCKsgs/e
/TpbbphJ8UrkJKGfcx5+ETdjo69fY5L+Q31itS6n0q7XPuO5/4qvVU9ArZIs
iUQSiQ7M7zDuMXmh8RDTtrLL1Ru8P60+gW+2ob2lX/Thcti3yjD9I2w0Uypl
v2o360KYOjUEFe4xLSrdR339GVM5JyPqqH0cJgmMdq8f2R4qP8LMP4gxcSYC
XVuVNDhVfJ/5Q94pf9EEYGDRrZsim2JrXM7Kl1SUDlJIzDr1h8NrD4CfBk12
jdiWAj68ICCX973N5SuTPtkqlpxX99mGc1NXLG7FQX5m0QWhR3XZfE9JibDX
Z2wt2S0CayGbgpAPa3ncKJhvPALH8j3yYPkHg5mpITYibjfONE5vfFcS4YRe
AEG9HKso7QV0kv76b80ljxzKIAWHZdyqyJ9qYotYqHoiPnakHhB55ArhBCoz
riBLoGIhnoW4SmZdwIvrGQuW53Lyj+7gj5boCr16gNzRo6NpEKNVD6qS/Vay
QIRX0AbuuzECoDUQ1F6DrVSmzv+opn4ashs4vvBhL9XyKAZ+KXJ0naWQ8Szt
1OMoDgthblM0cLSQm7s473OnINZqWrMI57dH3xeCekkWCA3eKR6NSnCABeiX
UNClTJ9aHvZliFsbJEn2MGFxRfARgskREWwjZmBxVAruPWtd0imobd2Fu02M
boNT8etSKZ/cke1tbb0ataObyInI/PEe7ffX4k85pYrwlocxe3P0qZvxeIes
EUY1956QbLAVLL8kkYbUDvnV+KwQaeBBS+CuYVYoT9ra2NBJksmBRdXNZZeU
+CE9hy2en+9WYR/zu0AAthizlOVFP+NkX7/QArJvGCHqQAih3XsJj0KHTzMT
H/H7lG6c8b+wquFV70lAW7j/p52PXToEH2l14OeLvRO32nhb1OtFmq+TAn9R
slUYNrzoLHOk1Q4Selb6TNrC+jOMCISqs34Uoxqp2jAacvJUo//pHEKmxs2u
Fomzj3QsGyRUguDXLsP61qt7dibh1qNhst4ZidHSGjnzPjLYsplxAijqRfiq
KfNB0xuYdKcJwaZKsKyX9uqTnHvrZSR1frG7eNffaEJDXEeQYJik5QkyvRXU
CrGKQ1s0+5PsdJX+iarSREPGi9zi0so6jBu+c++nLfzcslxMNjdY5brjXU+P
tD9k/ZuYUT0fx+JuvRiW5DCkl7SQf27yKqBDyBp5r4/q3zFLJjhDeZ4iDaUf
qhyH0cwPSCrqzu4hKy75GJkZN09cZJh4XwWoeRLarfRD4Ulf1/6aD/e2eWmZ
P6p6sUqmZMtMq+b4etNXH/20Wiuh2Y0q5d+W95QOyn4IgtqsCJrmRYODHzSz
l5l2FPeMK2tiUBgfDQ8Q4mkOPspHn61o7qqiK+aj7pYVlj1pAQzbDV9LXZ+Z
2ME98HRuyDcBhly/3ZoNsMp1EbT4sIxUWPY0Jd7nop1G04KGn5f62rFvne5s
Q+iZgcyxzatEEKhnl8cWA75LmXfFdAo6vBhJ2fKDQvQEt5btk9YIWw2fc/HE
JUgHq61v0gcb0LO+Ac73xP7fnX2Ttob8FLJkmKcuC9Hajmp2jR0sVjS3gNuR
pUEL9y3zmDyHJU0+mcEh+TblABxGcpHEjFuDjJ+rZYZ9/PvSlVb2bIBYY5rW
VGeKqpUmnDcGtpKX7IfMUGnTekp02NwibAJ4yeVf2J+nlkOjR4hFddu6OpvF
OsBf6bZkmfWJ0/GovAQPymD8zmu7yxQ52ixTX5LcQTV93Oo4I+g4lPD66EZ6
avmTPyR9HRvBWiCfGSAEPQHJHddWrG6mZXwLi2pHphmHHx3x09Zt5d9+3Ti5
Rc6gnhnCtY955UAvpTfxm6YG2dfEyFvz3r/oHdPmS6VRtCJfcNMBJ1FcfzhB
+8cs7+/BHx+9TXJmRm/pPIo6XLaCYngE5pU6SdYwW2dcnRT9EeKwLQWmHuHF
Ise/oBFZPwdq9Rz2Ig2pSy3jkQRGwIEdI2ni0cAZ29sbhniDk0DbeGelHMK3
5Okjn+ObCQZGnmy/Q3YsotwEUBZ9novZDiEryDaElIEATlOVL7RiFm38qI8z
eh/WGkaKldzuCXMAUDNTMEwMpkQ+oxFvgeU0BNHqnUf3MlKr5Wp7gTepi3Ty
Q+/uSeaGfrp77TBpjOyojwd4HtH+kKv3Ki15FbOCyI0Zq6UQoLgVsvV6I2T0
XA+L77aFFrfwHJq0d6ELuQuaUQXXLBnR+IGr55TjLYa4jfGUoPAF/KvDBNin
Y3fGyNcfQaHTPMv0fzWt6HbtaSSOPsEbRBHpRmiVvKpcIVjPlbAW2994/fb/
+ZARDT9tMO1IE8oCNkHJIrN42/w5J0HDsm3Wj6VsQX56f7bb17yFBGJ7O8ud
5sWv7hYB/m7lAC4GAiF+O0jGsRSQaQr6uMVcxLeV24Zo+aGMFnq8wEwAkkHq
rsyqEL4cBjrJpeZDv5KR9ES6UuCDpChnflBzCnugOxaspbRgNKL2g1tKg5SV
KIoLxnh17DCdhEIqzmAF+qQIWGWzeWhTeoMccuoV49ZwrREIiYPjI7bSq8WE
R8ZHmv4LX2e9MUEWnvOViMjhUGK9I9gxbjJ/yyMlIM5Cyc1chRaeIoTItJVt
jYIvGCjD10lblw2Pg29z5sBvL4AQBeuXVmo0AWfIFgIEjLdFMh7vPh+byWoB
riEa0/RmWPPySSP8M8HNlkrDehQzmVV5MPjwWjZyTwZ/TuE2dIujZ3BIXkKN
CajiAvkrgM7YrpkJ1sQkD6Zk/OmiC+Gvr3TafMuNAODuYk3r8qaqOMXhw3FM
XV/daJfIqht2lOYuCiiARYaBRdPty8vYr1dHPKx2stPIN+5uNLsR+jmf/F0E
YN8/S59lDWJbLivY8j+t/vmK2XxR+T4iN/88e10FCY9lWLaj2Rawq4XPszSn
f5wwTHDbPUzWUOj4xTpdQlFr3w9Nl7OqPJS8qpSISUk3CTEqvq86n0sAacMX
N+kVs8C0JQdZV9FTNZlenl6ewDmWUyKL7fgCCJXSnNc4xfKAOJ9+MDWETX2D
fDvHkN8syEc/Tznx6dC7jpB+v4f58YdO37PkWWURJjGLA/zJXsYXnKWOVElt
GinG62E9wX4JCP5A/VGzGT1sJ61uMuKXzwQi/5cAoohyMvEePWCzoEoQfYF+
YdBPJlfICmYUqCapaeBQMH+mWOp54dKTTUonJ/rRzuJ8G5bhibFV5foob5UE
wQ3hRNJAPPpWBK1AMJEFU/VICUzMRMfNHnyIoquhrLJgLhLXCTssKHIsQjdt
hpJr7JG7FoqD1Dc7yWvaznunqd94pqAP0uLiQz7EU5G6dirkPhLIgQnif/jP
5NbdcbxQckqLPopxanLNvQBAh8RjIqmb+Hl/gnM5maCNg9ZltSNXFPEW4KQY
0yOOpl+SNQJroiCLhzJUS+tlep0RPfyqc5ZIFJO7bDFZ7Gbg6qCKSnFxJv7h
koVdlhOf7ZRDSy/mOnq1UunV4hP5C2U5T2E+NGpQVh6PQxPAIGgg8hhzObXM
kNUZ4/bAHMxjBNolUtl77fJo53tpXh0CpzoOeHBdA7jJGABH81Wjct62PSzk
8dczJYXZ6PWVzSj3m7nBulAsjDvnceuUUh0pPIiPGCcW8OnJ87n2UR7Z6gVp
QT+M9LcxG8bsyfEpLW+e32KwfXas1QnbwFT4Q+pqe5EObyp+3xwz4FNcyw/t
L5PSxblnnVNNZ9TPb0GEvZc7F8alHp9xPryVsNrW1LK9PMJ5qHbuiw484R9o
2a3ojO7c31esQaMbCXJaJ6uPsRAykckMrYNavQ9JJh9CgfqXuE9tI5b9g2DQ
MTX4Ox7MMUnCoQSjlZzaSSWC8LM3AFTczPc8k8n5X2bQNf+MfGHiq1MPHsH1
6mczZcycfGChCXO2cvNbDc5uBn4lx1yoOza9kJDjJBeOPU/ldIPhjmyn5+ML
UI+kd4sNMk2sFF/ceoxITSjRhS0RWPmHG+IVSpJ94LbBwxE++hNo004qqCNW
dtZIZw7GbCLV/mkrU8jYZjNHMOkG1xXeWdHzmg4IVMJs+dLp+fqlUBMPuE8J
2LogkiAiXNflxXiiXC3qHswbz9DWF70bnGnKaDCLUQoVWH04oXvBmN0pFWUS
CUCD7qpkYTlw9BG/I77fgfLotdCxve5DsbtM9InvhItiYYXSnWxCYE/yZ15G
5go9S39Jhh/e+FUVTZ68XEd++KS53qonnoTwXv1/QcyaSe7MDS3ceQMBvCe2
zMMXUrScO2wCxNIvwr8gZoBZaJFIKl7MhDFafq5oyU1w9fWOFfkzqXJ0uZZ2
AuC7tAnXmbL2NOKhtKEavhClYSPKsxMf1NZgj6D6MsxWQXEmbgri60BTujVg
oT8MvuCL6NcWdM5g8fhMZfcyys5RtwDDMcom9b3/z6FgG6jIQPm0MuAWi8Jk
W3YAl5pqcDWiLXv6wytyaz+v/1sfp86BGAjekaHHAWmk5j2xoF7D1G5w4o6p
PIC9td4e6fVAFmTOcDAyp+QPD0ciFTwzsICdM2jda+LfCrah88KXnhQb03QL
SnlspQfV6Z7bLiSwz5KQm8Gki10PZXSy9q7qslRm96jBwkRFpDzYN73Vd3+u
PJldV839CNckZUqKm1tj/opm384u9WVKdbj5fYHFTrXZmsGI5+qV5aMq65ne
Zp2g86eBAavIFds8x13ND5aqVSjE0dRVhbdcgfi61D9/UytkHF02lX9WCNG4
DYXi7wlSmLoYkZMJh8DoiB3DtYw0yuih1GuIHFqRo1nS5XdqeZSd/blVRNNJ
7XRB27KQwl5B6pJVhii7318UsGHTCyZ1M3VLumSA8Js/GwAlHkwZePrAszE0
Wm32OWvcFyzqZoMtpU07NRX7if6gU+45/ObNHau/gQzf66mKKw+cryTu8N9P
FOGZ4CWtlNuKXwzSrVFZe60VCnhKEGYCq4S5XY/JYxzlaZf7O4qnoBRZNTaA
hrO4DcgxPvMGIp+hmlqkmOlza9eY9QNnw66f8HuNrpzASsiCodVyMNqMpwI/
qgCueWmaKP7upx9skMzMQ6nAYevdN7cvTZGkbyV7GlnNmMttsknt/QFPq6S8
8S1Ajjupioko1qEW8K7qtBSlwWP21pCjcbpRXkbm7Fox1Wb4qX7VPdcLxJjF
LmFNy8BpyRIBw+QacyEAl1Jp9L0ijhqYxwIVNVrJuDqEdML3U9jQZ/No7egO
uaYyBWOw7McdhzkjJlyqpaAXIMzVeUBI3sbDzczmmv5r+sNApTj+NT3VRj4g
VKIGgZah2RJR2XLnMLIbJf1Z0vTC3IgH+fivzzSFbcf3YBZQfGDfJynxhbbQ
5ibPpbZ2jFaAZhOAg3ZUR9/cMsYMp98GKqwNPtndI0OOEFVywfQc3eyTtCmI
mAhmNC+kAbLMG6zJPdGPGnSCVZ4c3vvehbq0RTAFjFO+kVFxYbu5Q4Yen4J3
fdGU2D6ZiNyC+cn+fz9ry9draVpkAoUIlPKe1cgJVwSGxZK//4H/Uuq+hkg4
bcU1VNCW1UhgiS/sgbwFUnRxpGjGMjlMIIafkJAeRAALJ7Lhv8VMUkfTT3lq
L2ZWJ8OyPFxG0XV7m508f2RWKWIckMyELgUXUwYh/Ckaf7BHoeiHyZ8ky3rO
naNB7ONP0jqDmITRrgPHLjB7Nn+HU1Gx7MkVYl3SrkKNa9buOeQLXAeOXZeR
JQfi3j2/v9n7FRURI1HLf1HASq6JDMJdAhHgwKWVDjhmqGbEJXlfpjjDSiA7
JaGK4hINkH98Bl4Qreb+0cyvqcztMXOx8Zr2zxZQWdkzD2+7rwOSymFha927
BO0qXpnX7P7M2XlkLzSHnXl1J1L38EEyY3TriSq9jmLrs06D/UDMOSkWGRMB
Y1/NQtjaynPSNXC4DfHz9+l1rvNqd+0O0Vz4Go+t+PTLy3fcwEGopk8sTc77
9i46NFgdoJFwVMC3zf5Aas4nTlbST/4CK7as8umXeCA4jaDNrWYdVaicMYkF
ItBHp84VrSo1QAIiZCQOtVCbSQpVjCeRl1cuWakQlrvJtWbogBJo7ETM57yr
IO3UtjPZYCgv8NHt/fTZKxVivulXFWnztZp5EhzcUWKmkSaaylyKgqhZOmfD
L+RZhTvBXBOOQWeqrF+Lq+XUX+En5+nRG99emKudBsH8C6xnP6B1Tgc66dl1
IkfgMAtVU7YGZ3OqOaAFmfQ4nQUyaYiod8oxww5uAul403ilrN6Ma3enWd7T
NsDIDXH5SXjChFV4gP7D96843NFNXugEeM6hPsJOw8VoDJ+VVgsw3UiS8WR0
4nr9fV902Mq3jH2Yuvh6a361judWrwegxwLzumWjrGWvdVm/iZchTngnnUjb
wtdELFBciWjMRO5wwvnaPRpadlPlSj0ymLQuhfnHVxpyhEe4s5/Vx3VRt4BI
Qnw1tp+HjfO1NUh2TVZlZJoL8QBBGVjDgPq8e6NoxfbFKcLOJEOT4Y/ubsSp
jP3mtQ/ZjV5oXovKu7zx2wiWuqlGMx33UsCB803x3X5+nW0XkWxnrk85Hmjd
QaQIK+DtE4BHQ/5uRgy4c/kaCHsMcEwlcVUjr87OCJhEk4FrdilV3RCCddZ0
PmTxU5yp9p4RHQkC2IAq72u/9UlJOnkrvENVVfq0G5XRqWNvmPnNLwPrmRcY
5C4mxd4dm0U+i2h/Ht5lw7O0YtJn61dZ82nO7Gqju3JFLyGMrLrkmTpBV7nl
p/bSXdCae+yMbFm1AV/wO4rrgZGKul1vHcE9gtPvYn+OH41yUsCG0jLdh/Lg
PgsdVWvF/1fK/y+t6uUvoC7tizbfiU/LjEuzci/5w4zMfI7ruRcaWiUp0l+M
+6oBflQaq0IxqQ2wTHELX7bePhy5pxW/qm2xTjiv8nS6t6VBFVCLD+vcaQEa
NYRraNd1bLCVGUOttFAbqKQTn7KeEU8QWZre5S1BsSX957nczkL1CMsY5xcC
0DBmSo71fEdOCy+wiEoZAYy42rD7j4/LgWpWcvct1ZyHBt17bBKnobOIOgxA
vhgNyXvkGd1uop5M2SLszcVALXTDuSxp3/pBRYcAHPvtyKfVEO74wPg8yFDU
8RVVqUkxNNvEw8R67IJXVjkYNYBZwOHO/xrdggk/OAzdCQN4POlkSwZvP6Cl
ctOwc+3RrZUna+y7LzeIg7ovfTVnzBjW4sn3gxLK9XzHPZqI362wSqA02gB3
WnSGXe4rNHJjfuvFt9+ky+GmrYeRd2h5BTI4cffAQO96xv1O1Y9/P6F+7iNT
tk0DqWg1HJpkElEJwCTLJw4McyP0/YAHQ7UMQ5AVov45rqXH9nQcdLAI1EFg
QZvEVL2pNg9OmIN68IQKWBUxhOR5MDJ9hqFUUx2hdgbxHkpEQLzvcc7Rk7+Z
4P5q0npJGpZ0RYRAj6pnJJjCigU4CTUAhXrQxC0kKjLRzSg6HEX9RZYpuJ/K
1ImCbEgbmSRRvTxMF1HEZGZak8koN5TUQfWraM/RDaPLA3M9XfsH98prnqaH
9ZJUGVO7F0SXzFJM5j29v7l48EpRiTmeONzbbFtWGNetXRGI6QFrlggKHj6T
BKb+7SSWPiYntpnkJEA5za/LZnZbpVto26k7LM6r5FjEqXf9i4Hx4N497ujh
v+omAUtrSp9ubC/LhV5Ca4SDDTSsrKdO/kBxfQ83njbOyfN4esSyFEwhV6ew
KqrmhxIS30AJoAOuRRhn+MfGsypGDTvx2sCeHM8jtioBG61QVaJQSq5S/rvs
RbQRdGhgSM8Iw0UC4GF4qik8DJH9QwIStGQo2Vqg8H0enDVSS8oJnYP/jGvc
7WyhzhThMt33acXpggOZwOFxidlvWRSfBfm2B3ckcNPjRda7XWOTZVzLN/de
cOt48LV1vUnD03pfaK8fIynDJQUD2jBk5sNuzLTCf3ej1NnmFRSHn9FqjLiH
BFFMUo9u1S+Si1yQAPuxkxQeqyWt00/jeXPz7yM5wOkYs7uPUQWqaiOGLM7A
yNfh7pOfEgzpQuD0VrDb1MASIKHOm8wAPDL9VhTS1z8rNvCdkSk7QDLum0GW
weHZxQQ2PklvqozdG+vwQW+9oelZDBcC5bkWH2srwOLaklGZDLRkPyy3YQcq
S9sJhDeduUJNDslg1tTmPRnsGh8++7nV5LJuqcB7jP5XCfJGsy9loGtR6f2P
mDJ6dt4MyLEqn9b3aLraz/5j+QIYV3TrFLhmFRcU2S4VofVAZNw4JcdPg8JT
atGi7h9Df9LruUSQDkw/PO2tIZ+vNZ8hLS5h3YLd7fHvA3tXimd3RWJB163U
lODHx0BaAC0UOnZFMGNrqg6Vy1gomBYynTAsT0SunrbqbvtsbR5oiHGkxEMH
x5+0JOpVZzfkykgRREmOS8VyE73RBAafKD1rW2LpJSUBBi2MDzOsv8w0LgK3
IN4N8HKrEalNdQP/iR9pm2mhM+eT7Ieftihc+QUk/wwjnuD35au09RcU3SD4
iARVPr9PwyQDldBRjKDpM8cka364UA0btgAzxCqJOPC87Ujm4Fr7elzSDywS
CspsLIKml//+v0WAo1L8A0U9ltEJ2Zoe9LfBH5wbnqDV/9FepgJK5bjLFOVb
1sRgtIEYW78ECYPdTws9//3xpzaUkqk6c2nxzVQAR0NkJMAVSBDiQhudF6Wz
XH7UgiXjGzzXii4GizJOT1SzxbpmC33T4/RKTYwYRF0urQE0bv7Jmn3CNx2n
G+PR2bhthlCuTnboLNh/6r+eeN4NIKxDwLtCeXK0b4DPtKl1JMk9WcT1oqQN
IE8Mds7tU7+bZXSOZy/Asdsmqdr8C/aSiuBR9CsY9TjFObXyRMrbJCBIBGh9
tMLCor3Y7QQTkAj4pJ2dJMQ6tUdlT12FdZEaTVGw05UMXuG++KB4LK7kqZpj
2C11v+/3TTrTT+8fol3UgsTIOPSQKX+Sw5GFULMq7w+jy+rvbzxezm3SvBz9
8bIGwJvIkGw+bVuz8j6KN0niDElvdvgrkn3vc5YLcCofQ5h+f18tnv+VPIe0
j3xYKQOlYWC/0m2joeXPgDxdM9UsWpb0tlCln+NNZQ2AYo1pCnxhTErVgijR
Q+t2cMSZxvKSG9lwGkTbwfaFeJILAAZbN8aqsxzzRweGqPzQvVxcRk3T/ruR
p3ysRAl6dqtaQ22fU8xzDLCE2pSI1zRhBD2a26WHx+0DnCq3+G+6C5L/pxTx
L4vlU4/cxgeKUOe4KJTssPkz2JXmzQ+IaAWcrR896ycHEOoSJyVVUeawFxjO
GwCYkoqbmWhkb83f7PnglszFKxKxjCCZ1aYuMAl9KTDx546ms+SxgkNlqPEU
P5aLgps03HK1zXpaRBGBWdVUKzlLZwYUGHx0GUdO9V0uKl0Eo0ShqaO2dsyZ
gi6P5PsniUpaF5xjZbPKb6EFzz+zA+AmDVWKmXDI9+5CbB+KUurFg/I3bCkO
Sm3sZ6hSnTP1yvEaTtJdTvk8D3VJ68qMGcXXSg0CTmbyc7V/YkRGwRQTz5Ev
Kkp+evIGKm9iTRwvbOSJmxn++eDISN32vK8dik3cgImOi7qLw2bCuEAgT6c4
FOAaxkYC+3tZzRGTtuSo3yP0VUyclblqVe39Y+eU0YbYmw5N8Z9czfdqgjGi
WSlIo+PLJzxfi/3h6SOq0draOrERy72Pxm4jfwylAdzc2L3bWeKnjfnSoIE5
DSxKwP+4TqHaJ8JQgD8S/kPiBtcSzAGVwGN/l4R0qaZvq4yfbbAyIgeALYoE
7DJUkrGIZztlGsZuB2SMgZameeeS57BSHossSwvurRSDBpltSm6ksav6YS9s
ICy3AZASGoklu9nOSzOs3jtn82yeLXP4cIgVijA+h+vPjQPLHp1BeL3AX7o9
b5ePIVegjtsWV9kmz9kNYT1vWCHV8Mthko1bUsQzSt7UVcLqa/64roK7JMC7
djV1ghe5ozYRdF0MHnzY78Z92yYzlt7WQWESBJjCpDLtST3X0Vxylh5hCalR
g+ESNwswYPMozKOzMPi9uawaPZVeSQA0Ro63bLZAiKh+tkNbtYTt/l0dRO86
WgEnNgynKlTwTQ24038vM9L6xKSVbo9nOILQd1fc08o8sXtXB/1Znq9SPWbi
RdDTqc2rzydDfFlt2PD4xh8PqEMQ7dmBA5zZfbRLK4rxCRgSsnr+eJ8pE46E
PqRFtdxLoU8elPGB6v7D5KSZnw/RcpdoeVf3d/T2X1Ml1cREz1PIxZ91OWsl
dyUazVPHaDUfJB8seSL6CXZWfLXnP/Krd46WS8SHP/IfhjyM5v44uhgaOpQg
FrA6BfJH9ZjHH5z+jCCkug1GERkQH2vbv/JFQEaVhy4eDzqoXuBDzLPPR4Ba
HAVkmEDuSyo51tsp0znFXBd1qZQkuWqVJUijxdJiOGXIFec/oPC+vyTFE8fi
hJH90+z4xqpEntszyjAVukBoLKEBfeEHUxvbYTFKhhV7TgZ9ZHRiHVTEOr/X
uCQt6v78n6HoZkOUJtSwKWgRBfH43RhCqVqtKxyarVT3jjqQ9UGSFEM3AUAP
7P2tzANoazJkeABQZDru6T4kPbHiUjuKcXNl/MrtiKSbEjrysufaU/mjmZjm
g6U8SCLlUyv3//3OvqH0dEZMqGg5x+M4GkfMHZNzbbjiomlnIXCm5eXigNjp
ZElrlGW528JWPjIfbasaBpIV7ZLtez76/ShT8NCN9HnS2z+k1PXFsWASd1yt
dK1Qwlz+FlnvcV9t/25fZNIKcz1l7rUDecQHwNYU8MbhKvT/CsO+1nAt5n6s
kqymqUe6t8i/OU42tjdFTv6eu76SLYt5IJ1qdzh/Ign1JuEQYHU8H65DwuS7
2ptaGK7uXGtRyb1/7HxBV+uPgs5G+Y3ysd1apPznG2T/0LoNxvrGwshlRiZ1
MOkgKc/JrZ83Bv8HjATp2IV37gygoSvuH/DkAsiEN3u60VyazMxmuUKOj7Ef
rrGgJ/8fMDijI58YXJtF9ldutqf9wobxCijy+EJ7xEB+3YIItfargMgp2iM6
bHJwl3iI/JC/KisbZZr568AyisLTEQbyeciVHQNSR6gMCMGA51mUhNtL2brs
tBsM/vfw8WDMCE1YY8Rw/2Qc+z++7RcNpXH81IHTvyJbIBoBT9dd6SdGwNt5
97ksIGI9lvNeLxbkRNRF7nHzo1H5d+DYXqHQ/lWVxHFSi+KO3E8jNCBblpDT
rPVT00qN+YTwWeqGALX3rhsmI7s/yzNF8UUBnnk5qQO7egtbxKjoqI5v5LYG
xv9h+mP7kk/358ljER1Q74mMB6TkP7mMHeUWSFD6nhY0H1Rx5b9Vl4pdjmvR
JC1r0d9hM3/wGA9+AWHOFZURuE/fQ5csH3M1G3A1FTOFf5SwI7asMRi5exQT
t33byjRiba58fT0zoGimuDCpwNWBHf9G6KutAAiGBmUbbNOtq5PP2Ue6hZ+Q
LV6AIORhpUoVY2fiMxVqoea+j4Z1LI/tOxWbzbw6tNlrhbrXbTA6vUEaYv64
r4225ohqjen71UtQ1hM0V0NXgzuQh1+IZ7JPnmLWxXtvE+SJqwY5Xy5Icjqu
LHMDOEIDwfdGSltJ3Mj0Dji9Z/GohZaFuf5xMMDguO8wOxiyHAAtxk1apMyx
Hxyf1TWN9VUx+zDwZBC7OKYG6F9PD6SwBNXzrL3GeCjiaQ1nEz8Lbjf0aljW
pFdLJHAn7W0/MTb3/92VOo6gpCliwYJjb2Pos+O7w3Pf1/HsABi1iAsC2az6
qkSgAQEEAqW1CbKCe0Rqyil3Vi6MnOLRdwNIZsNKbvbLr3YP59lsBoZb1bBX
uluZmASbLWdpbWJI1t3hGQcKDMvIPCH4jyFi6n47OUxxaGZ3oKkg5p0A1Hct
daBV53B6liYxCJoMguodiVImvBlAFWYtE2De1qSCxcrUn5kP7ZoWTIzYSmVp
HUoRSUfZYk2OE/IwyCfaZuU8t8rQfAo45YFXjbMsJk0QNWawQ5ybIhe9qnDI
FKWov1bgGoGQ288stnAQbSuAuRHS+v5UfqqWNgellTyuHhArdEhkKsGFnhPl
SGXC3gl/c9lxZxT5nPpRSoFYT6jqe2ZZqrXBpz9PPY86DA5Y1Qj6pGDXhHAC
Z29gvzIXZ9Fcnox+uSDChEpz2vH7TcWYbRToXplWOPLRzUm9bW3HDRvntvjl
Ak+9xt4uPYJWQaXmRm4tLuLz3WivV4We/aIblu90lWqbcQoVTaqX57+aMDca
ifWzKcWw8z1OpwyqL0YElxkTDJcwJUpg6nZqENxOXE3s3097C5Srrr+S04ar
wLve+NMGpRqAqH9g6hwv4YSJCJzSf5+7EqMNOZ05COM9WusK0uC7Skg4hvd9
hHCHf14UB/qKc+PFF0OA6KSjj1DJxeNptoNGwt0ICdm2Phxff2mFfTSX8Iwj
61zBdJ5DfJxYahp12K8t4T4mj+2XsiYQKfsRgLbMmSFiM7OgIuZBmr93aRPP
dZQqx3jl69Mo3Y6bpPv+A9NHSgsRRhN0VY01SgpTIM1s/PfK7FymUWGkLwkh
kAmXK/L1aEtuIfD/v/rUbqQxj0I1PH7cSKC4Axx+e5lBvbLDo5NYwwUAJfcv
V2xVDTn379zyRE9X1kwGIspOiIVZviUawZfMYkWMMCvdWsat15khpzD4ZpZt
OMdpngQQwTCcXtLxTeWInAYYWWeR7cQre4M2jn9CUCqeBFintYkzECqm37F0
de9gwjiJ9qb9IYw8rxI65I0DzI8NJ4+nVcNI0Au+nrwVYMiLKxKuO3Gvd40a
2gzXXk47I2uznDVG5ex3+OLpgpYkR6LLs4mrboGtInh3ZZHBeb1y1PNm5zLt
+3DYeoa9eYNe6BQNJG+JKknE+PAncPspvG/jbOqj9Hpjj852YocLeq0fUFnI
/AOOOBlRZQVKXgozk2pNoSjjh0Tm0QGA/kRX3mKSVJqeKMYRMATayYO+vcw0
V2Pc89tSrHhZisCWrVOxP8CNgfObYcBNkM0Ucb/jbW5C2Ra7GCQzC/eMKXL7
zSQxYNIkmdsVeRSZbP4Mkok3R3iQZ1mEZznKAlaoTvEMZzNwwnjR6/5v4B7Q
L1d2S6v+eGpwTiHW2XTcTqP753mSUyu1PTKnV433Kzhd8ASL6pSqXLm+yWDX
68i0n340345zunSZOUKPF+7tmksOLq1shwhdMPtCSbVzyv1q3wcmS4EJB4+w
KiVsSeM57pGtsH1QlNUlSQg4eIK/HMeuJb8GGiCbZtQpJhar2kCbDi1n0jO8
weQaML6kVNeMCjnCznGtGHLnvS9lijAMOv6YNk9cld8PWVW1hdlAhzqIYM8R
G+EFgcbFHDH80QJOKv3UelQDObQ2bJG69mslKwvAFWM+eRv2ohQluiULWAYN
Yh1wJ0EiR4nCyIS8rP1ceHqlaCPE8bB17K2f1oFjNtXISe5fCcwx1ZfcPbM4
cYmPvaBnwbhPEzZj0uSQ1CAC9VJOdaINGB52dzl0cqdMtEgFj3bIQD9TrMt8
c88nPAeoGYOcC0Lo7rWpYR7PK6vwi1xLDb2SSYhRbKoFEfXwmCr7somO9w62
Bp35NN992KS8ZshSX6cBjVkozApzh6pFwSMhWGg/1yonMIXpzWQAT4LJUJNy
70sVQJCvuX9aUqdDVsH3PrHrXLmqfjhwF8V6TkeGCNwFMHIUWknCSAxZk1bc
DuwxfQNvVCdL1uQCfHqSbUy7JuX+2GjBlsJUf4eVI2gGFe6dnoqtfhWpWXgz
ZIqtQ0c8dfaj1b3moV2Zb4pky84Gmsj91xSQNps4/yr1YmlVuw7BqVrDsnrd
fIzmQBv27kJWiwEzuY18oK9Gk/L+KE8W3FxhE/OGj35fiOXfkn/7pQ3vNL8a
dQyUU1iAB4CeWJXJPqJfLRdBlD4pBJnmH+jGMLVjSNjHZET11h4eIK4AWjIr
uHG6jmrrgjFJ9DZi9rIaLa3FmDUB32UbuU0+L/EYG5dDN8Nq9czUTYbSCvZR
otaxDOJAq8uDgYEIZQKKxUZLx93vWvqi8oFaF4EZrUFf3Bk/LgcNVO9+DCMr
leukCg7XfQw7e4z3clhPodQ9Qc1L7GHPteCxEDS8EDiOFUwqI6prMz0CMOzq
IO+Kb6HeI4vz8+wkQR8r0WDSv32DyQiB+P2Vtue3ABIhzc5yv4zLQFoIw2s0
v06o86ljIK1h0q6HlQSS0k3dpItA5XTpOqAQO8JNOsiaVPUCXu0aPofq/xq6
kD/3VNM+1jstTwNERkGJrcfwY/tmNYK3lMIDg6K69xwzNU6CJeaNvAJj9Dsf
bXUaKaPaN1O3CsNC++FGEUNbXhMMrVzZ0cRsZz2GdcPWIFaqXOf0gU0ZrgD6
viyeUYXNe0G0TWI17B0nFwWIQ0Ue5mgllsVQ/LHDrANmoLwhraPkzYso1KeQ
AkXnSKn1Gvwybia8Vfnpd2h5334PxpMaE6+/INqkXp6XLYNLkLCjfOGRAVuK
csSvwhQlrrlpBw/qdnU8DMLnqBaT8DcqhUPtMDcGZupzLvcTQzzTQnO60KHw
QTTJf0/3Xc7/A+UK0lEziH856Pa6Z7n+tIKuA+vxAif8OeNLsmjFArKOm4HK
G19KdE0aeIZZjYx1C1K727CoT2nnxXB3PMVwPanK7tD7UnXwvnJBELpg1dD9
NASAg53dAX/z3hgWVjVkIf0ha9PnIjDiQLfscgK6mhQFXCEOYZFwEx70sJyG
rB0WekzGx8pFoYJonfZ6OwLcjQos6CfeKoTNZWxlt6Tw6iAZPv955xq0TMGP
UGLmqUuZvhLo/A9C0BFxuepu7CWcY3GaDi6/b0lI9UczD1+KyWNO18hUUboV
fCM0odx0HNtvfMy1vJ6yMPyyUwlG5RbGe6hce6n+CretyhJsxqst583OH7jW
S2R/lQybx87NaK05O9MAjM4mebugvMdYXt+psf4zLOk1QxjNkYpXDPi0MWhf
lsWQtdOnvicJaYqD8h/jfo84gxnxapz6aC1yADzqe0rZDV1TDZfi4YfzNqoJ
CiOr6VfACbd2akI7C2tSKaggU1sOo/MfnUCIU9KsgL5YBEuaKNmMbNXO6EQl
kTYAi6sNaFbYPDu1aPRwQpfHhcxsWF8ovI8zBi4npV/2yhALKpfGBbsUPFD7
titSnGd9sQKVhoDHpb4elpYbI1Ti0AoBUcYpBJDEo+ly/vPQU9nCA98wRWIS
Pi+PCdA65FggbwyD15TD0zpHg87WAREo11faIG/XxnMeh0S1a2RSNQ857uPs
FsnfGaWKfZfeYj7zraqJTP6nPx1PYtNJyAv9NCXblBPI4eGlBDEThiD3u2yH
Yy8Hp6pc1QGGJNa1CKon3WmINqMaokCGduI2j7MLdHGIjU35U6Wc2E0wYz8q
NpV70PbNL8M5Pe0BmhnZjEBTHHOSvFMAtAGBRiCewT1ZMuAY6pWMWWdrcEKp
ZREtXgn+36uP3tWeL5jouAoWjeXTvOxbCZhFaj/w89P2/dUxXYcYEx6oOc6y
DGMsjq4mavUrGp4Z3FHpI4WtelIV9PdFO64Sya7hSk9DI016UHVTgWGLE+54
M44ehOOYwaKS0nWfmJ8uEqkb8IJ3Y5lPDJ/xyboJjHu6BXUuOL3XX+ZRm8IP
moZ/kHjfdOEAJJqrxE5b9P7RaGgl2sO3cbIq6BMSPUbRTCudW6r8a3QNHNjV
/MjRQZ3k/PjPoCGb4TFAuZ3ah0qM7njNiw21DHyYSvmdneN3rx13o0XNH6fc
yAtFK1SnCbp4ZS07mbvEUlWPcanUNwU/7cIVGBwlq0MfB0TDCKNxcbFeAers
VKV371dk1fqlErDdo1M7wKHTI6JBQGajf+vVPRuCQP3wwPojQpHrMIw3wCri
7OWTXy7EJQCM7zufFeJVLv3KFetu+LyeOw1v8z6scrUKW5DLmW5YfHyKEa1M
jlOzf/19rPAbTbGXbPMNbq4GKLHAHOm78EdB7DLh+8rI4xDe9+OBA90s3+6F
ADKOYlciYwkxpfVWuZaDUQnXm88Z8iupc9XWoN/dn6+Klzr96HsT4nIIVx8p
zKLvSPKQHvs4WfABQ6aJ7/4Nsswe4D7DnVLFvjb21ztibO50DY4V4Z1Xrlhb
n8s8w+gMiD4P7JIdH2RbVK9gn+SIAIGlvODpicYh7y0MIqr5EKYW0Ksz/KCP
ZzRlwxWCfrOXhcB6HI3Lia5lG6I2qdmYLKVwG+sGMbfEZ3wuw+tVtFluD9hu
QoSB7pJ44MLONvCJiQ0JqNpfmlwuCnfwKKAcMHj2HTlkaeJ43/N86rmGqdXf
yIAr6BaUtXIMadBwSX6GMI5TeRHRkYArYl0MNKyILXfFWgxwmNOnD6VqXIeR
O7ZMP8dAzjlMAxWMTplpHUFFw3pTD1l3ldZTWTfS5OV+usQZKhxWSh64buW2
6IEFBYF6VyABFOQG0fANjvlx/2rl/BJgMf8Oxb0mBmxdgssY4mcbQuoljiFg
o+wq0r/q5lUKDHMXpSboFxT1GcvDsl+C4vwC++I9GvOnhg7rMINCvlpNbtRn
yrH8w7Nq3szTvaY5yP22XSPXCZL/DrxWkwgx6Iyfqpj+zbsC4lXW93lcj0rG
f9fs5G3iJHHHu9zui7vXMsuMHDfT1ywr7AszB0qUlk2zNTByKKYQk36E74W0
HL/+S00/Ruvm+V7jpIS7dgnoNyDzXeDkctKgY7MryV+l1JCC9PcNhOqJCR8n
LQ1HiORF4TWrVsgJ4Qj1JQ3PPr7AcK+G2dlaEy+0LWecCyEwL0WOObOnrUXX
TCzYmeSr0/rfRUtkSE/DaSGXI4CSD7/e+IoKZZIgQEufPRwmWiaIdjk5Qa+T
52IUtsQtvICBSzxsaYGcprtQXtbyv9gVO2LJrHDbNc9Ip89RugI709amE8ZU
j69xhSY2sgXUKad8HQgKs8ojz8DXXIp+zEBot+6AYWGmnx9TFL0k1Xo+9COq
N5jxn6WOwMoNvin/LAtNQa7hZhASz9M3ssDnIbNtCJ6/k50TOtVLumFXx3wB
nZpbChgRrVm/kFRAREt8NvGqGY/bCisvKkLd8RFfuSzuV/iqebzieFpX30Os
uyMPsXAEUEPN0nA9jzimFBZuKWNctrGs9nufSXkVeALqFwGP0oW4BsgJxSw6
BGVC0+CMK8ZzC2tjITY1hl3GwWi4eCFRX3/d5eu4Qe9PjIGhLqTRbzrTTeQw
Ojw232/13/wDMHTE7oZc+Ov/K0p2ndh4pXdZUjqtz2rzfdGA+uQBdUL6fNIn
5USGv4W4jw/FofeJ5ZZeCVzZUTTe4QNMHHJq2tg4qM1qynf2CntkM0YkPMDC
apu3NLwtcFZLOCCX1q4ApibujD4LaVKSPRV77g/+8uSyX+g0/Jo87GWstfo6
FUTkEbt56Ls7Jml/zUUj2P/vuzTcobHNktxd4lWdXE0eWTO7LavZ7tYAmc2w
K10x2OEHF3zRArj1yk2+ZzddF8EEbv0VFyCdhK6MnSgc/uIJoM3EgTV8rASJ
Kz8trHhMHJtOmrOEZ8Lyaq/F62bH4V52qU54TMmc2BSDNv+p+sme3cXQuMgK
srhCuqutlWUhsBn/XBQyff4tJFHndHI6xRcg3eEivSLJJit+bj6FxAVe2dVU
Q2mgTe+OYMN6V8c8GtVjutKJ//5A4uVCBr8lT/oxBHVS7x1Y2YSTwJPmue6A
AA4S5lmIhfzhgfDgX6kIjwzHvr6x8B6j+qwNJ6rzoqpT4V1s1WmmQGZeWN3J
P8ZfzxD5M57iYoFZRLCD2UJ4uT8nmWPqC0QIWOXDlqyTjWzaZ6wCO9BlXndo
oksGrWuOAwmz2QRzAJBC4BV+BUTxa0g3FzYQ5uphHruPee3JsD4iZnRPy1Jc
5/yEnpPyiwR4DfR9+w1tZeezjwhgkuWkVS6G/NLVc2E2U+VrrvLsY+CNwLri
fUXfRGX8L+suMZz+zfll0L2gZdCIgIJG/rV4yp7EkbWNV/2x8+kTJj2m1IBv
NNfoLXqkBYbdD4KHdXgacdkmxPYvtnQ7MWX42kBEhPpazEgL8bamTLEnJTBA
GWGbu+eg2J4tfy3elRQSe15j5BVef56g5VSP01K0aSmkgcQoCOcUETfnsqYw
Ek4Ec5T+nxM/PiHJlTNE2fbO37aMBY7mXpz0cUNLla/9y4XSb8DboMRKZVmu
5u5uXeMPXm8CUnSD9segMmpE25QzzdZc0YzRGRC136U0EH40eEBon1+H5vxB
Wr78/VvFAFmto3Nn3Ley+9ebwG24a0sau7CpLiURoGzoBSfj63kshFFuyNK9
StINrJx0YqsQFS5BSZydOpmKz/dWyj/8mzBaJEkh+Y6Ei75PWZGrcEBlJ61r
xR+P44PRD7c5Z1qpVeUUEIYwZTcCAIaDjYRYacpGpiN/fFmPkiJPGBy+Kefs
GpISsPvBzWtP/BN900yH+kHRaxaA40DGnZwdXptP9WtmKEAG7wuKT+212zaC
Y/KjTUIZqknB9YwiVjWmoID4xTLuuV+bqdWdGdv6oIiO5z35ZxLJcrODbPUk
yLu0cuzUaXJrLUXpgs0+fmYhQotoKB6Ca7qPK6t+XvX4ZrAx/tblzSyoUn89
EJBfffd3jKvG2884EYfQvX6ZadCyufJGbZKIMVGJ7yavm368IFU8ZIIaUouP
9kPWcKZ8jZ05gfr8dLixhpaiVZW8D0toSwdFNbbkK6dogEZhvbT2kLVZ/aco
5EcufzdveY0zyIslL1bwjEY/M2UpefMJQ5toDhuZ0f6FzPj9cljP0t3UQNo+
smwTCLv91b5nsdm9eTlJIIvsDWJDZnAxz+PJWvEHtwIiDi1MT7r0aZUfrO6l
jD9GEw8n3EHU/KR/bkjBKcXuLuFFgCS0CXeKBIJVLFwnXSTw5BZnnJqJGLf0
Bjdx/N9V0ChNqFgXXMWCVCB7kLXplEEInjmsuWXbhhCheuhZtVoL6fy3kk/s
5nTiz5PNSb7+9DYkWnL1vo25p6LjDsGNv+6mIKmH6qMShsxqyHq9w49R+uzU
6AtFK5NS8+Rw+evfCTRfxdF/0H/n0FFhenwNwIttxMQDgO0mGhX9xFFgtcff
iEYrKLylqv9zUY7Qp64B+1zD4UUfXUZhOu56sbBFLfAPgE8R2mJezagx0/Az
2lsztfgblWWrBd0i5TW/PZry+dhyY6NzgeVam40iDN4akxy+ATzL6CqgJsnh
qwBnv3bhUufcH7n2zGFccuauEU8Goi3DD+hoiqWfBTegL2haqHX3aXDkAVtR
YdQWtbLkqnKZ8Mb9/xvqZg/6Eroic56NC8CBUzGIJ7jeh1AsWnW/tSAf0XCS
6mWUBexzbkDQw2DQ2l9kRx5Rsyy/gBQHoVOvZdc1kvSlkJl7dqhfPoDgQlNL
0JcZjvyU38AlQPqbQ82xCLvvzuWXdDYRi4BoJxk6+FY7NTto4NgIViaRJl+U
QEYY2PfrQepzReYPd3l1IxHQ/23kwtc13UXadEuJAmC+gt7GPbj/Rt0X6S3G
4rPu4fcmF4+f2agB7dVlJPB6LMCqOmVucu/GfDHjNB1GbeHX0MlUgq06VEbn
tU98piko89b9RPu7lSA+jj8aCUz7yDfcdcAIIJVIMpB2qBjMGCzLS2EuMvLm
3gzX7rtnPI+d1iO8PX31cDzzX7RDwkWf+qSojwbcSMPcS1NDh/O0LEA3DaGn
+TVvNJqqrwOKEtBaAtza4C78ijq3vqDDTUy7sJ+qdIrGFwePua6gpVWs0j5I
y885mHSr7jRaySK/ec8rI+G5SODZtdaPipPeUjq3Mgz6asAmjksIU0tqzd1F
Eg2HfvTmqHLy5OWJlRKlr1DGoSWZReBhegJ3h7yql71y9sUXdCJuA8RWUCUl
7mS3baXBIBQQgJIjIEY2L8e/SAxXCk1iI1lHZV5IiyKoOIj29kDopL8CX7Jm
3+TCYmTMm0pt1Z8rj2708q3d+DmUFXq/LfNRtmV6QNUsRdIoVLzT3qNfw347
+xILfwQfoIc98m2HdaLVlgL7K0rSx9SrRMTlZdy9e2TcuWUfjG3FAPw0UWaA
6HWEnm28J7VIvfWMeGeX7Dz7wWC0fjUGrU6u2bWEeWy4rQGK4MOYpJKsDn/n
9RFytI9mjOvLrO6teMlIAl7Bd7XJpfimV2/PYQhV/5/8ZLndwDeSbY0HMzp2
QaxG69iJisPtbPYn4yO0eGWCwCDr269gfDcB+Yu6xBq/HktTacnYBO3MRf7g
e1K54Ky074xfhBh/aEC+/SO8B4JewZUBlcw24cxIs+Mw04Jo1bL7/2acvtNv
Xqc6BhP4E0UOzSMkcIAt0dRE0ZxKzU3rrFdxHF+yJD3MG1MqGbFlWSYb3k/I
G6lBCz5mz55LzzkV1rcRSWIXeB9GLJL1HtDQErsbt6iVTKQQ1URutQdIuDY/
2LpUlT1WwtRDL3y9mkofmtPZhgOcM0yGZo1i8Bv1a4HTvDyHlVCcwjyTFhue
QV9BPmz0hsS7HS36QkuucJRzYTYiNjRMb7GgnO6mNfRHlxuvpB9DFbJZ/WWL
0+8lzgegFTTPxaKy16Gctmxa+oyTjhgbpuU0O2jDDMNWAhbSI/MePXV8V6SH
HxdGuZeTF6c+wI2fLgPBTzEvCei3jQRzGlUlrbAdziOdkHqfmP4zsLaXQbNq
vEuN2Vn3bwaIEKu45p+2+zBbjU1CecHnhikGCgaZXC/DwXABBmzkBFYSEjMl
QWr/fmYBwqdMUaz916P40/whJkKKOF9F7pVAx4uZny/6seFeBhEIB61X/rIy
dQWz1bK4erM1hIP/rPvmV5PQdJPPU3HxPaDIzjgy/NLYqrjSBrBt2kMLdSkt
DAlETBszHgV46sMbMJu/qJsA8UaF4bK5lkTCrxrauo+re1eF/9PKIl3f3m4g
kdjn3dfns6qNsqSpn4+HYTzjCljtGHUl5q5DDreEfmLMJrHQgDLeZk4ee/dQ
Dvaw5U6xDJcsQrM2qufazoanRhZ6QPl0l2+Ud3RbWOJHJxTiV45Plue/6IzM
sAbY1TQ078VDZHs+w4OJRHXJY17PPD3PdxBzq5k4F7hYdVubbxKaLWetMRdT
YbeBUEx9SXeF6GhzXlv8tO00p7PfSCktQrBKtMBoGxh+oE51WWG0FtPIAuSR
qO3tJ6/Q2PgXZHdw0Xv5M5Om7uTFx++lyc2+JWE5fD6p21BB5E2n1QD84rIU
z5SC9VNPsPPKlZ7zCfEVxDR7N4iq1GEtjkYKh+RVEe3NB/mdkruV2ohBHYQE
JLZbBfcV+4t8js0kKeotSn3NT8UQC4Nmn38KBFiqhF1eLlI43wYzbPjMa9m0
4DNLXTufkY8XzaSj4t/DBH23PX2nSggYQEmHJe4ENUllcRHKCLZSnnFP+eNd
6t4sIvTpR0x8P0a+X/D2aM16+dUoapf2WXz9vlra+ZLmpo0L0eOqxUh6nw74
S+qQjPEKRMLYuXujq8rqGCba0FH8xTPfQQqH35/d1DNeYWFOc5HrDNFv/vz3
GYdz99MfQD0RghLBhYZSdueJtTFbeN3CrEp729y0qf86B/KaEV1CMcfyN7iA
ek2EFy81e4qr9vGii46iTRR5/L2M19apFAy3bDKnv13WQzV+45Q50z8ycpzF
lT69W602yoBrTIOb56Rz6aYBeHQCsbnpciQ5LnEmbdTMm+vbz1uzcRYq9rFm
ZOeylD765qFDFQZK/f2eo7fIfgMAT9wA0qdK4D5ki9MXcHOeqZuQX+GhAiQ6
pWUw033OnTXGvomQg5d1MgrtfrBmDNyGu4Wy2hPxbRoPF/6tt+ByKImwYft9
z5gf5WYsvjidJom/ewn3L2qx1sXyvsD9tWttsCLcfnrOMxSN6S+EJMlhz6YT
N5kdQ3hZYndzukkOvotTKTs2Mg+KOEw/BdsMfB3WVDWG5Vyk7YHDK+bQxIpV
sXN6bmBeoe7txDlxhCqtIPTkbc92NFWNq+QQBoMSS8lR2U1NIdS0+lc4N6cL
XX5RXXrLbgMENrPaLtJ49MR6FjQPoc+/9jNGHP0YUGAp5LRiOQFNsqcYCRBe
ozWQt9hmOFiSohVDBZry4jIcogcxiv2zjbPwOoAvBZNGxTmGIZxsU6ZqC9aK
+res3bOLwhHSxJEInoaQ2kpzDJ23nJk3XiROZxRWjS6wKC0KpktLV9Sag4IU
0OlUSSqOr+3/c4qGuNOq0cohurOQugYs62hhoQ1+MjijXfB1EsBcYFPw3mwK
mYdctLxA4vlrIpcc+w2BVL8xu+OInCuY8c0fK3hrRP1Yo18P5x/6cgrNm6+M
UGmfydmLCgXUWBXa5k+f+snfMgujOpKzffywYuy2KGckat7itbt1ZLZv6aJj
v48sZf7iy1SSurH5XANVLqT4YsKwwA4oJTuDvJ0O0nF7xVVpX9ULzUHLip7Q
lvXBFqrE5Ym/E03+OHHia0NVgTKDKS5aj5hFfM+2rGcwpxwH2Ks7FisU7DJ7
dZF3k8qoCzFFNUciV/37opyDww02Vf5fEhl2v22G1X95om4c6xAjyhy+KRuO
8e6xXa2reJKtCIhGR+yKlRu6vCF3dN++fcJ2dTDCTKtef8lve2MWDH0nX2o9
FiwCsPvuotX6SmTqgTwU1+x6xD+2qVi4vX+NiYc3BCubUS4zhu9yQPAUV6SG
SFcIiTDhwGi8l3V47sKbih3wt5dcYKgrWVQyXYlrRi5w4eGRKW+87BreWJPh
YMLH5rrW3PK7wGdZUJxcR+zFhZJl19Avlu9Cnxpx68+4rM0Xg1N64TUhAsNd
//GOkOqeaVfpIa9F8Eg2KMVd5yitoHe5OjPsUDrTyh1bvlUGNS590hRkkNTT
6+vaICK3YVv3ZDXGWybOdWVpHDaDox6cWD/qrSeZ8rDjVS5eV8ILAt2zvhDL
sXhnYkJ9QMc8nvpnR2+/Y65vIMgJo4fqQLZtg92FawOyuWmaIau52pA3AQVs
Pet0gEXC/67BhF3nOY4J8rIp9g101w6r0MSWPtTmNoukmmdZq691ID1Eb/eg
WPnG86lANDpbfqbyhkAvh6VdEzoub06pQeeOC97lIy8DH+lurQWUvyaaol9j
o/stH67X1LB2pol3QUSQEdP96K/DHXT0WqF1YD6Gh3WoOKixque08Xyi7Q2E
5A6NmR2x1HnPyvZjY/qByxXQiaKUZzfqpH0bVR7eYX7D3v4mpc1Ny3Je5RXm
1AB4GtG5vGlXDABu5/IfIVsB1/Ia2pZ3PBCGpU57qpNKrAI9JEaQ5q1cxtNa
gdbO45mhiFtIgepZ1NJxwldgZiKYWxdld4jOgHWKN0MqejN2QEJJDpzKGu31
I6P8b90nVEC4Rn9FRQ9lxd8n1O7XaRPaaUjhQD0JgcJ0iJwpGMAIBNqxM9rD
py7cRG1D4Y+33XJt0Zuu7AqqDKFCV3WlLVvsyZLC6VkRb6vwKRwIafVxCQaT
IGf0tTYIpHovve9jxBG370mqJ0UV7esAMYm7iif3+tJfvkURnNsw+j3Aefpi
LOV8seZB4wyQow6bwGf+BgDS9a+P5vZ91AUW07KBF/y29PtoK/FkHFeLe6CH
x8clPQJ+xEzTKZId75K5ivbeOuMUp3YgLLSbqpwzaNgBly6oWLtc0gHkdWTd
VoynMMyQilBG3az3BK0CBkeadcy6Jb9rVcBrOjciMox+BDseMkTlczOq6/NE
OzSWNmpXn24CAVrgFFwtRhIgf0X6f3/u/NZ/oXoLRQMS/avqBy0jk0Ir+fUl
OuYv0ISw7++AlO4H1pcLvq2Z5u90mfQUdg04gdiJFaGtztfDPuDZ8fTw9Tyb
T3kg+rpra25uvMyeTLZ7uqfysjHltlsrQ4ehJl+nleY1Pe5TNDqRY2MXAdzF
d8CuJ2QXpBZVfWJQBHXIJMG9rlnI7mqQjgbOXJdzhb6n+hmsx1Zp5bC+38D6
wMPY2KKdZdOQPh/t+vdxF7GStoTWIw0sGmeMN22qLgEy/cU94/D6xGc8o4MF
m8FJf6M9nLfBTfI7AzaOBMtETSnmN0zq6xzu6dx1ae1mw27VvSQktK3W0w9x
RuZyitrXtMMSJE5ohrRDFpeisDfJJdJRUHgF79rJPxzdWAd5/5KtYTzcPmn7
L/YLeehH8CgQM6Y/JACYQeySQFzbEmHNOshTdU8wiVXGuOe0+qiR5oVcx9fK
1mhiF/vnOhx7ZExclAIyez7BVsJNHZ3ds3dQEW7nRSZ7BDxwTNFd+qi6JLCQ
lpVtt6UOw6Ik6f5WVuh2Bc8egH8TngxnHiodj09aQHhxen93vGPP6nMEfYRY
5oyvOEX3Beu9VRf71yU8rVaG7zFwqD4cb9Eir1yNg7fxn6jkOtOtAXCDMfTz
PK2aBa3UEoSRHa4Gi4vrBhSgDTSXS+gXIK+EA9x6rlHXeKOdKg9g/VWBYMOi
TeQOoOQs0W7Y1He90fJy3EB2i9NGtfX+p28u1s2rudofG1JZ/WZKBcOzCAzW
29d2JUnmpVH8mRBiRBBQedizJcJrNqkOUU5l9+IAO2ufYzN13jMmMZagC2h1
1cNF0CJTq8YQo9ONJ/UHldEQA1pyUeQS0jsHwLNhvakecWc1njipdDxyRylC
WFlhg69kvvXLo63ccde0JIF5EMemQux5kJ4Ubc+Y28qgGQ9jxwQixk05DG8C
hjyCZxFwSEfEpcC87FcCX9OR1R1pjcxddJJ11UHM1OuLwb+x94ZFNQIiwQTP
rwGz4ha21lJr8bEewumrfO2Y6ps/CmxL4rdvYV1fwF/fGf3iKkl7SvBAWeLb
s2X+PxRhS0mkjcIdcnvcGJYrZfSvT5lAbV8P9rID0sC3humAQqu1RSHiY63V
pg+D7ZYdd2sUpg/gtJRdA0Fi8X5FhWvNa800HtUY9yaN6S6VzWLvDFzUOPI3
PhopNEQz/aApu6nuPXlS3tyTDRuW20nYqi7XpNnrWpari/8iIXvE/mBCbMPm
OArJVVBbEtLHGy3v9E4ziRqkY788g3pNlgoAMRMX8OiRiY+JHvwUh/aAGdea
xBNZCLuzUx3Scql0QdDUAIJPt0zgqQDsksdU2mUSZTm0FZxZm2t+GIZn72NP
/EgdJ7CCalU6WTyv2b5LzNQMQgDKqYM6V0lroOv/CasuCyUlca3De1BUC0iZ
sRHxdmo8irn0tDNwKIA4NIkgXGJN4KN0kJH4yTGo53JNAFlDQT/mNbM7kKaM
hsYX6kbcNPk5WbL04PTlVIsIn9ZyzrIVe7ulVU0GbsUqUi8WcjGLwBw9VyON
wh6b5+kBn7BY/5c52qsqESAY++5Jmgr6xf+BUBv/7i9qqSQKHVDOTvJIq4o4
GZsfAu1bcmW7AlSw2BQMOPxcPLJd2sF7VOaePJp86VbJrtB8aMlTjHwga7NY
+ghm/aDXJyPWF7coBxNSQSPxK0oQgZlIOhKX35Rhrd3Py4h//JAPnSpSvTSW
BHAB3a6q8CjPReYBzfpPrm1XuHVZyZvxYgSLn6trT+NKh4icgyRDZGw9Qb5J
vHT2mr4oXWqybovrr/8ngFKeZAYmPsNUpmWdahXDQZVZTe6dCyxWMYMd6qrB
K4NbZ7/4iKUNN+ZPgUooMlf3hghG05uUYrI3lbDYbcgcorIa983gzDWznWab
nnZ6uIYSFsUAVqWDyMeIOH/EoyxSS4dwFfVA4VSDofzc/3ylM5Tn7upSJ17L
yuWigGTAiSX+bkp2zQd1NmD40czpo1NPodJ4LUwGxFIKUZOth3MXgStHdmXM
sFmTKID9+26BIcixNBZqrOfJG8BQ3swEBgxC4Rv5vW95NBDFRik/o4VUNMGk
SdNY2GiLKSdzHCQixJGUwtDNnoPLZTnfv2eiETfPVCmmBQIvjnjWKyONZ28O
gGI81Q/cgWlj4dN+J+9YNcSmI7CQxtWu1pPFi8AmLMcp7U8A1SRfFbrZCA2c
XD1SwuBkaGyAyhymnEPDTsMMHJFl+mwDG5w8oAFTekGQDHVghYJk/+rHs2Ls
AYZX2mR4sQNNB3nhJfHGyZGW5UeoPFipI8LTXThTcOMMdll+gkH5wNxUMqLx
9oV4t0PWaiqAvpwXBFM+G0sNismzZauwq5EMpqnTaAjXm7FromOafdzdSfZ3
DfM600ZuN+McWoDXPXyg5MtWmQZR5VtOmAFoFJVI3g9GYG0OVo8dsVRQxM0P
zmvVPATpoPwqCQ3DXcwTDNPsMLIDsrgJf9VJiBl58gVAFtKUFPnY6L1EWWrL
s4Jbbfl24gPm91Z3GO5yy5OTjGhTinuUVE65iwJjkvC55UC6vLcsvPij8QOG
9w2A+gR7XyOebVwhs3yTLVdT/tjLUTgV0aGDs1Ll/WJtA+vMK74hnqLWkyHV
BO+ug2ASLBmj7UW8T2M7Av2xlfxfOcVW/5A7us6v3+fvORVkb69Z+jSNg+PD
8GR293VvExGlnE/Le6Cn8MaPupSJGkpX/JzLqmn3YO9f6PIRSj8rFxlp0YRU
lc0Jy7E+xIGVkF0ylusWcTpW2mq3OqBI7vMzCE0HrIR1XMoK3eTCHorxaDK6
90gTWX4b8cwmUIJxUJnIFLmDTSUz07pDrKBZDuk0jPFjta5KXhcu0w2N+Hf7
CCpvkiwhePSLkqQYk9JafAErdYE0iKICCFeQmT7VCmxGFxXRq28mt56n9Odn
vjKMdDTAKlgbQ2mSRaHhtqJK2xteZwZDUnWAR2nDHR5DCr2QAS+TsijVX4mE
zguXL4FdmaXvZb6+96DDZuKEx3fWptOKHekx1N9iPDxENJC1YcEvR9I2TVDU
u9ftjVZmPzkxTN7ZKNQPEknh2bIgtjJbzjVAZU7FAJgieook0nQrzPhHKLk6
aIc7ySyMnAwLJEbaRmxX/Qto+c9eqO0EJ6LJhK3tS4RwCKOlutm2x0yVHvc1
Q6xZVvLF1XdxEnBuBnCJ7NF7qAyI9fN3bzdsCh2OwYvQ/MyAZdsWuKhwpgiC
PN3Vaky/Wpasxr43RmiSrbmslbIqPf5cpDDXVVGd0xcwAFvrze/DJbeVZScc
nACi0dVtBugr9CaIfzOR/Z15PxVvMcK8fCsQyDfU7Kj3dWr1bOyEHfyZ59Fu
Bu0sa4V9fUP5kzywFG/UNT90sf95XsIRKjqC+arY4Bfd0UE55VBaJIfW46GT
PQhmU5cpIjeeQzNnB7VzMOK6eNXFT2YnRR8jtDxf14JXWrb1FZ9wJO0QS60E
pkOF/Z7GygFiY2I6IX0wdTxNtwtI9j8vcjHyftWh+GQ1/trhf5sQDKTvoBih
SgNdLt1cg2X5i1/0975L92HGp/WdLOB+SiVYBLm0s2zQ3kZl/27Vz+Cau95+
LojC2C+ZNUZnGre8O//6199GzXJKRgOK9vtVaqb8D6JUUrRmUwbxEGEWHNm6
JFsoSqiWyiTvI02penCFi0oaJzEBEVmLLjC97nIyVlhNVnIchyJHLTwb1UBr
c5oBn64L6E/L6C34zegwKATFNWSb6JbKMZz7VJEgb0dtGmrh+dYnHYqTVyPi
eqQ/AkaXakioRx9bQZqzMQHrrP4d2hVJaWQJ4gHxMqfJ2Eq2DMnsiiJTi4o7
dvCHwMpjSsjt3wqSJsbPInzMFyjljkyCWnBXwihllvFOMXbP9319x7QIOb5Q
2W1kTZu8PTWkPJsCmlfikvqnVe9flnBe7UUMlWixE7HTsE9VJUFmPmkExXM2
keqA3NkDulR3RQPJ/lSC4OMep6h8P4vsecPq4cDhOX+uFzCmDbCCcg/F0enw
VjwehVbpLIvoikurvU6TSHH3oOWkJqVuJ5U3vGxbKvShs3hnZx5tfv4JosJ1
q8KrGDEi6ny6w/UPfdcPhIRge6GyNdVbNZ2Dpw8v+5hdhOv/eEoqKUnMvh4R
VQXGQvQLAtW8ZZSb9cZA/ovPeDZAVLJIPJwuLMiGaiIevre2qT5V0Y7asXu8
KNoHd5pd5FYbl7sajcr/jSzIsox/Yx9bmS1+ZlsYFSRPo8ehnBJAnIlhleAS
bY31z2s+qMmINAAza22SbtEEsXrORuMwNUyV2D8QjtYW76DLXAuLlrf+9iZs
4IT8dxQAVcVtlLOYWTn8NQLZzDcpJHaCcE34cd5BBjonbUW14PW0yxirK9xV
yb/C0b5l1/DiQS3EDaR7Jx1Cy+7pSO1SH91Mtj/QCsz3wrsxfimgSdPl1JOM
rS2AuKHZW/ATtqke77MK9lin/SHgEmqQWVINxzg6BoGeirAx9xK2UKttL3/z
GJlSt/d1QBqlSlyzwNiu4gSPgRmWdwv63KyTxkwffL6/6Q8xxiSnokcwg138
aaoPr3O3DGs9lcGbsqBVAY2TlV9CxnufXyjS2q3cZMAr1r3S/16YLIMX0Omw
EjGT/z3FXAsfMCQDIrIVv0cmNQjmaa4mNBQTaENB8jsfAjKd8NZe3RFFyuYY
92eVRfzfnFKMzG90oUV0pM1GFhtc69V4Dwg7IvUWt1w1EmeZ9r2xGNYYG5jQ
PNdwc7fEccf9beWbEKXLELSRsv6jzDtCcee/UKHgVlhmeWKPaq+CUCqIEk9U
ttq5UtxCFJkr7EbEU2ZZKjIA1zFuoStPsAdRNZXCQady+BHgxXMPJdyViTgf
OqwAsd9uqQy45ipLJvTCkTZEJrQ5+xuOSj3jOsxQOLW7HNA0n0JfybnaY/Ff
YlqUCp/w66hcN2qJIsi93SlzYXYPAHI59aT3Vm1XQt/AJ9vgdhgXcrbAOL+1
xIXN8m6b1q+g6uSohnrf4p4qL+458+JNQPC/YG3Gmxrhv8oD1yqW6fLahI4l
4+NSG7TCnEqRxA8bJUfUlfL7cEBGUnL4CWKfNfrT117ROpqbB9bovW+Un/DP
qISCqrQehbFiwberHOdZTYrEwS6QK6Gi3y7hPQlV21bzyFhfZ1Tq2FQsa08S
eyxLtd6HVGxCTNKrAZPIMdhvmSHKg5QCep9GF/k6clf0j2xC1U8p3T84hnT9
dIz1h592hjY+svTCGF3F+jJzUvnvlfKdGSw6DsarR0SfAbmdGAw+jUyMOWXq
7rv/YxHzv3beJT7Wj3hkvXv2mz3qsM4MA9hFmEFhz2NuyGDS6H1plze4dcYd
MyG9ryzF3Yn1y8ylOvaL8khVZpj56Grx9ZiC86kQkruWLAgM/UoB6tFH6JL9
jXH8Qw1gaPAXhSwoUBrOkeOL3gROJ+/sNnAUT6PeR7eA3iKxwdwmtzG59Zwk
EZ7H3f4j+0AcTQZ8E6esHmIObw+Xe5E3JLLxkAW0UFIukSrkSPqhy8LoC/sL
jHNy4fCMXO/A2WaM+W7v3S/zXUt5NW7zCanqmcsyfHsy8QV817/Hampio7uU
6ap4DwX+VQ6eCrVxJKw5nrWaylejutgjc2vgT2+rxC2rw8McJCHqpSxWe810
LKZemfmJc1pVO4FPrVPabOmwa9U3o9UnwgbktCTqoiJYftdA4oinydlLgR6K
lrMpt16o0oIRxIsJnDbxOrh1LPp6dPR7U9b+xJh+LPEWJIy+QIhrcX13S78S
F64UQSKNrS//NJfiTxowsYtltG4uU2Jw3JfC8jobivBkRSQZPyH0OZ6xIgy7
sfcXM1jgb/Vk0t0oYKzIS4mdql7/I5W90TEBwIGJdgeP5YDMR2ztfzqNmgrm
YwU6qwxOfuKT6ZbeidFbs6dprxl/YQVmCuoYaDwvXtEEXMzHY3z0N8pl2QBt
khuq0pr5d+4AIuSATMXa/MhaDx+lOTXqwlLNx0PjZKvCgY4WlAvzQ10U56ig
Zc6HmoCPbAzP5rHiiHiCZ+XI7gAEwg6tDxe+cfAg6M5Za/qTflw8ksY5Cuse
gbjtPldScumhdE1GRQ5s5R/v6TIHHsUebrZ7CbmFmpil6++k8Z8ZNLgVOgNB
Q/XtSmamlf/NWc3COxgga1XN8fzL2of0lS3WhwWlS8VOdosJx/8F/89fKKfy
5/InH3KlGvVPhzHZ2AGXZ5hpO7L/dbzyUJzlV0hdK8mApioU31xKfp7SdeDy
tY1AudyxYBb+B+FltDKD93xfDvFrdWD1FtcQdnY2YEL/zbOA6fpc5ii3IqMO
WKHPugTKI0X2NsPb7/xXODVM/9+kfMdj+ZqrYOD4AefrG87xBLLdWKqfHbGX
1y1WrakQLxkPwoE1w6L2aOcmNKFdUZCIe0nNybb9bYTE6gTuTaaAoFCKVE1b
0PvKtastmyCn+WWkvESw54skxWuvoETc9El/CaWhtt4+ZQVJrnT1ItQMGCUj
6f0DnUjedgFI1mniHs9p2ZGfZ++EvEja+wIlIQmBOyv3dJFnlk1ajEk2hFtJ
uiz2YXhyDnuQuw/PFS0LBmtSddXYgq90KF5LXIB3D2k2cx6F74zfz+eQTXR0
qI4oL2/P8lqHBt3sS2AmV+ysDfE8WbraJhEhKbzFEeFMRgNJESCXcffbuyD8
vUQXQ/pEcsiN7pBTzQ3OcWMGCWDsWqxcy8Y55LYXSDmWzNoP9sjm/zKzjcbt
qjh2XmZgmUVhIWPS+EqBG3rIyI4nzQhdwJ0FGkkMLcyIVk10fqoWaxpGXzqh
gva9omKh3i/Bv5CajO9FinxcGDx9A0dKrwt0mva65XLQ43ILkS7mMU8BQUpJ
vQtQ0yY9h4nLIE/zzRSbifsAn8gd9WrdYudHku7tvCvdWqOl1uqZh8hMG5b+
p/900xc5VTxEORNiaDQjerMZ2oW1ZTism2lBjtSL4Yp3QULOeOS1ioC+JTuZ
bgN0AC16N12yPpUfWNr0vcGVeABTGKIQfI8i1wI1sCDdkUUvkFJnY+zDmJfw
UHEdYlgtRIAGAXGAehEWxizE4aeNPj7l5aOpgx1WcKMXvqyC6F/TeXbBFW5u
ReaFJoNu54fONtPqpaVZaDscs7igmQAtkgTAv+3qP53pI036A6t7cIITXqof
b78W/dJaAhKIHhsvrKTQPLqIrA3cV7zQkmG8FJhprCOl+1EOd9qomh9bAPgQ
S91WGWzVOkFZViL45eiQNOR4HQ8FSwVJlIU5JlDg0vHF3lIjr6duxVl6r0NS
StH5MFvxDysZvNe/JbV8lEiWtJ6qvkbmm1ROr98u5nO0B/2eDRf9RouVihC3
Du6DB8OyeVH1qfJtET47CCyzHKl1AWyA65P3S3sP0B5+XyxwVyXnEQNTHF5E
Zbuq/CyHZtn3oRHoxs0Q5PKb7Kh/E9hjDwf3W63ENplDJT8AR6ZS8s3zMgic
CCPAchMWPwMNDR0ExgCWw6bVnSnWOX7x7aFiJ8PmIvNzoW0e4iUg7PzXZgnw
dyptz3dssUgtgqJSy29J6vqYEOSG5ysXGd71RjGllXRCept3WEZPyJ5jVede
Gw1kPGkVOub2Am7JQB2FZJeb62N5Wwf15rBYxOgLIT+fANR484ijXNrRRuuE
jOQvIN+Und6Cb/jLKEt4ck6rWKLSfOcdtr8FXCSP9AhP/nLpRPoatQzBBFcg
R7v5PIueUxUmbuQIG/tNm/q/6GfvIpLzhGwga8dvfNXWLLpcUQil5VmtQ9q7
qkQl+aM+jUv9Ivm2q2xnFN9d+/+G45x92CVhpKiKLyKIbRs6xH8yMNkAsUte
8Rmj575xKv7ozMFYOT79g8SaRE0H8zOsRwpLAGGCYDfzLv3vcdkZYlV7CDTZ
ieZoQ/AkwAlodO5v2A4vGLtm8lOlLL1Y77hresredoTvV23JnhsBdPbYaNF9
Ez4Ie7r8gfcLs3XOVTsZdUCJeT8BvJAzr2dgw7aaGooA7PDGngUkLtBPbIm1
QvmRds+lB8s/4JRJIJiFYKt2E2XFLUv6B6pZ97JBtRe/CkPBjOa/rVTkFoUT
9nrsnUpqMNaMHc32UrGD8cciw0sKbtSuupEJR8gmfc8BaFCCo25iycF5q8oE
BMaV4E0FAAxTmPWQl18a4dIdnKXl8lM0JtJz8NlLd/BjD2/tt65d0G8MxjLb
LL2Yh43zpAxf46PF4rKLZIbLGBPdrmCWGaafcvVQQ2vvHINZ/avfXZg7YSRS
8svizNjvfV6ng2qnynLgp1r3+KSIWou84GkrcLkF38EdJ670G53rV7lcnunp
+SESnpmXjtmx9mIf4b+EhA+6WBosapHt/zAVvr+AuQXDayqhd6sm2QZtRzIy
w6WtjMx7RZqkR2Iz787vfT9ZVmVG8sxQrfE3nLp0GJ/B7uMmhoj0Re+g2lVI
C0SR6c9a3q7zOmvtxW9Ef3XIQcdGF596577dSmfz2KrCKSKLmrmo8nTuIq+Y
br9TGoQ4zzt05KKLiEHfB8gvJQ3QMtzL+cyhtm3hIH+HBoKEDnFi78m8BHSJ
MAbxwCG81vSP6ISP2jTRdW/lSzZf7Nu5UIZW8EV8zECNa0vZ0B6CbZk91plT
e40BPWMOojdOs2MLR+bj/k56qimDKKYaUxFF/WcTZq2kVGbMWfYml8XIDVs1
8WbfTCmuc6/1mJ47no68Xnyet/kWyAswlIP5zEgTp8ojJTjKIAtUs7fcXTRE
EjtEaRi29SbYV9ABMAoKvL0i4QLvSoJSiEcsb3UaGDRHKJ4OHqjzzvsSAgo+
xZeF3l4y0PR+bXHC11RFvVCS93thlWOJwZZE6cg6kqM6yPVLyVH2VcQBIvqT
BRNFOWr0IowMqILuiv71xOruJnXMiRYp6du2AZC3LySpYiKqmi1iR2ey9alg
KOo1iYrmvpzB8UnTq5X9joWS372gdeDrtjrJA1ho/jmAYq54LbGdT8L0lw1b
bVW9UEpOtoxBNxyssfb7JtKU03JtyLhZDp/4ZZfDOdrPRgNymfJMmo6lgjDQ
spd3SzkuMRRZvCZ5LoeHl/kcVXF8eamsy4makzI3JY12jvvSTo2+x5v2QKyb
Q+S8TiJV+GVAXzWgvRNB6DA6J0DyvSOVlK88SJRxHl/c9bqQg+26AuwGWOBU
AVd2ivgy8f++LvX6fJMcixLl+gm7MYurPAld9kWAQFwlBRO7BwMY5tMV5NHt
6jpQ66vQd4Shbn5J7Rrihg4b/jiaGBPnE/80QtY+UrQr9v+yMOglhWz7hq6U
qh191h/RMjbm5ysMd27lTIP9Ovb9q439smNtElhNFsRY3YZ65Xi7J6NM1+7N
9kJuFtzPtNvaJKccZ1Y+h6/N5I4g+CV/keVbDD3UdvBADpybiEvYPg50DK9I
lpFBlUyU3rqICXW0lfx1WDVbM3jyesYBgb0qlLE8yohSiJPVa9FduJJngCVo
Ze4EfiX3aGCLsYtU0VFZij6Xe3ukAUz21L8J4PHStHvKaWuGc/nCIKCZe+aa
EwD8VyyP1/4NsiUaiASZxdvSBkaaJqzaZjob53kN0AwYSuZ0TNhQ5M6OXc7R
NMC0ZC/ypj/ScXdSfZCmYDfhPg9P8zKvPA+ACoyH/v5klnuFmat5bpAxaxPr
+9EyDWQrqllHvmpvbuLksZ/2sPH9hsxXcBpWoVV2Eagq/0lyf2/pkNA81JLq
65JqWE+GSP10hnJcbyYCEUbQkfKdIS8VL9Sg1HRaChYygTcAi/fCSg90HaQ6
O35dOC5dy77pGvafXmUCQ6OgFRVHmfgioKVxo1VD0wicoKnnRWo8oDDVRQIz
iHIONJ8PMH693cHk4W729BbVc7yhg6BbiD16wtijfgGgD3lVIbQfP20zuhVZ
UvPk1yjO7nXpHDQLS3BG56rBCE4Ndcu2atHqZ90qOHY4FDd8zdLnu0h8toMo
T34yP0IBrXzooFL1K9NPuf3ewZF+MA7wXlMLsdJuiVyB80PYO3zUQmq8SksO
C3PH5k/c223H2V0gOQ1fMlQ/9DZpVRqgNXTnLK6Z9z3XP+jKSGTVrwv5fHL1
2BNieIX6xGGjMxhshiJ8cve3vd0GQ28fC+tkUIGRQmdufZnMLe012H0j3L3o
apRZYdG593H8GRrWRSlCqREsq2YhmNmMjRLoFfk1og4h0sl4iw/c6Y/cMIh5
G1Cc1zzqHJMT/pqq58H6JflimN7kpz/USoqWGB5JrZI+ersIr41ZzrjteE28
eSQuTrtDsCBElAPUFGa4pFkU16NoxM/iqKJVtq/FoPD95QsveQTFa/F4kJ+h
SYnMFtZwyqRBzTlez24S5OWTLOtOBcc18cFEYrgUYLy9bsQHMPlRpRkZQQVE
30EqrUD5/rHjlU2rTTGmmdIJ99Lw7nZL5U26d6RAEN0VteMc/5JBnfgTu+GC
hRFLHU/u3Rubw0D1PLoXO1RgUbKAYtTeSTEYsSEdH2Lp3SYA8Kvdd3hQtM9m
PjaQHdIxs88Osg0TdhABEck8BJIxsZ1nLHxmUfo4kMJd5SDh5DSiw808splY
WqkBEUltm/iupsOi5WfH4L9nZH4wPSMsKSMLZCh1MIeOEO0A0B2Q4HiS1bKt
FIY918749s4eWYb4yFfke/32/nMYGV5AC6KUcYxCfERyCgSq//vmUxsT3jzJ
T67iT7L1PJtBX/Hrv0gyuAbOMysVne4utKF6wFl9szsV4uO8LXT+TxduCseE
VP/pKTEDRgNFkMt+LVpoMe1yRhvu7m1SZ60XHgUfU9SAFJHAH0ktNyC3bhYV
4oj1QeJrxUFUc86AwLom/5auWwTSOUHl4+dEINvHLY7Su535XXyCkzHRP5/I
JDJPF31zHxO20PMi2klJpOpkfR6Hh/vnr2P1ZQfHjJhD+v3xXlBz5Nw6myQK
PGS42fzbGoHk+PZRtaHvmcViXuMaPHbDaRygw9dTpCJJ/h5+x28YckZypdgT
PT3ef4NnZFkMiPNK5x8HfQwWLXQinXIRsuTs5lBCgnurTOTTUZ+eDBVU1n/Q
jH+w/XMFltzzKzBJepKKTJKpYRVdgL/3jvIs7ITIDexNJSZLEqE/4XlGjsYc
NWzqC9bGmwFTRsYBA3oP1fo8Z/TjnQKTAyeCcLWYFCQrcT6AarEACz6j4h80
0TDPH0QEOcSjGTd3APRZWfcFydBSl8BQCjIsbI34IV+hVAVy8rwu4PylEpod
GOScOpCdqfoRCn3Rs7zJ8k/2tLfSzxjqhiGPlXg45+DI2D/ixWQ1X94ig4oy
0MQl6/0fH0mBdTOzoD06KmwlB6Xr+C762cgOxnQE7Oa1OPSda71JSgL15/Bz
phDQZsvFLZ711Q0qoKA1kDA4tomaROw2Pp+tXTiblppqRKl4N2UVAf47Zlvn
oyzdNodQN7EpJpV5xGxbI013d7nm8+Vs3MDkSuMnjOKzZ7f8vbK5sxZsMOlO
JrtrIAhMBIz0l4CWgPa9NibemGkor7cRt6OIVIRFsVFf29gUaPD6E8AX05r4
xodeOpMswHR+mJVYjbTWRIrcYER7Jw4XuA+WwwyAKrxttl8bA5Z3V9nuMbiI
paw3xBYz5chfTpT7jbr6ZTDNYjxRrmeIYCBKgipdNgDO7vLVzHLIKwAJA82Q
9eLUfca85hD/Il/rEXDu5aSNMjv06LMRLAptlqNk3MtbAz/og/i1+onbnkID
+hptYn8KwitWM2Nk71peelY9C+A5fD0qvQTBzhQyVhETKX3B+yYOd94QrQa+
eMFbcp9D75cb9Sq6GKDTbyt5TjBaDtCr722Om/SgivnQ1MUQtr1/NJAXpzDq
0Tn2U8QkstppqqEPrg92kq/0R4t6S2Wwi9rTHSSkQe2BkuO8BGKo6bJOKdT0
7B6dmR8WLfv7OO71t9IcNK6fsuOb63bGB2FC4n9/lWp/Gt+TvHtwqizovPMD
DgdbXgWYCnsSYbVdDhQx7jRmrn8kxWKfmJ4i6/S8odqKEo5LPrAPFadyjzZe
EWmf/Wu7BcZEzx8yAqiXMBM7o2s0/r9d/60ebM/tToJRF1nMv4w72RphkfEv
xTS6lSkfS4chpi1gXeaDbj5vdqhsGl2CAnSvnuZDFJ7amtps0d/tWv71EeWx
2r+54diLpWpyUtCQg1rgU2bsShvm9WU/5vfDg6uEUPWzAZvQFdWMELrL8b+g
v9s0PcbmfmIe2VsTWRUXMpiGHBmWuXiVIoUFUKAt1aYrlFWJTPANev1PglID
SlbhPYfDrsi91qtOrzRPmwiXzMVowA8Jo4LqebGGyLT6P4bW1n7g0R2qjqgd
QcuMnNfzEZ5y7cZj2c+oKCznt+he8ikQ5jRyc/98pDBv/keHn83dlpX/R8nF
ZEdRGq9o/Djf6qDAOnQjlOPwR5wXg2ERkSEHWBgHy6A0q6FubXnU4gS3MiNa
w+T2FxGSSbjqwkIq4na7pKjTmb6FbNEsN7BptvcePd6VY5P8MZddtrec55FO
y6xf6Hcuv9r1H1YGbOaFvupQhs5y/iDZxQXrE4zFW4S7IJFMh195XCRVj/Hq
Q3thr0Hkeu0qtf4ou5VF3sfTA44WYSAZJfasABS6rMsLS4x+sNIiyPxFDAmF
rfooecwV6FSfU++1tSc2EI99JC2VNCvSgDIucs23200Oi/9TBfIAr7CdW7YP
RYgpDP919cYZCin4YViSiolSnSF6GLFFBiEc5Ry/N7TQhV9vuebb1y2O1Lij
thNQbzooXag8chtzm4yyuDX7IMjIx6oTvqUVPW5pL4wPYw+3TqOFspVxwt3b
R8oBHR8ZvhQUHbJ6f6DeVG3q/KVobCwmjC7L/SrRr6LzFkQBdugqurI3+Obl
NQKlgbf0hyaQLGS7UjF+cERzwiGtfiMx+nVgxImq4OlkhL0CQCAyblwnpczP
y3RSP0u4hGLpeWzPOGMghVuFAA0WCKN+qNfi1OMiKHVETJjp0+v69UBPYt0c
+Gm8tDwQ/TyJ1bmufrTMTHmfX5Cq37TEVOB+li6CoAmrd/Ly+wQdtzEyhdin
oAa75jjxmrIrirR5EaLBEN90xb8h0h1TXWFH+/1tCbC8O06wJEjD0cA6L0nO
xkaFFNGdwjklV+BpmRq3yKy1GKpo3aw2Fn+7but+D68YRFvTCieEzq4ssAzw
vGo9RSX67yaPCAPO9+N00hbJdJYa9Yx1qpDFzZ+oJWzqZ7tvowIDArk7hl84
djW0dUavSYhBnQaZYqkswEEWYNB0CE43h2gjHT7tkGSXwYG1uQH4ZOl/2Pix
KCQsa0SoArhrpqL+U7CpBSJ1utLYDgyzV5TmOr9UVa1PB4IlPrBXZwM5WHzW
qc5kjWzi3trYiFy0Rox3Ag26138td4VpGW2l5xaWVBElhrXHr5Svkt41ibFd
8pXcX/CVV+9bEovk+kRDOkFC6apW8Aiplsj2G110KiuvjucuFbseERzJe3pA
plVhlvcHI9vT5sk0itSQng/swht++Bl+ElT+xV6SeCWtuk+/lLTzbTpdjmcS
ntACL+/e8++hyqE9Jth28OUvAkzZVualwSR7flUi7pEb/Y4OLM5Fh1V/lnxH
sL2nRl5d1H60sZm38GrkHZb4BCIuJUN0Dn8X8wpJ+ANXB5ZAn+KZJUGBYvPF
dEdG0W/wFdi3MMixiVCM8fyuYDSB7YDWiV/XQiwfNzHdvqCK0pp6DpRTlULT
5OAf1YtKaGpxcOVHC67aFeub23G1ggcDrc0qugsB0pk2+vvJ35+biGQrWzOX
3Ejhphw0HjwOMquDbSvO7DW9dNrq7GrNArwDZ/6VmVoIL4HjjzCsBFHIcFQ8
GGMUgv1QcRAegMt9Eosb0r+QvxmyriDRxgqgNkRbijHC3Pvp4/Pleqz1G7Zs
o4qr3h+p6hXRM30d8HGjAxppK+UKJm22hyNB4irr0XoJ6NmeVNDZM7QG78Ee
4MBHKfbrvy3XcB8UmZaL35sKFGbWEqyTmXrKVWirbl5kb4t5bBYXZa5cxYPa
DGcacfluEdPRDMN3WpDS0XDcbWj8rNW53azruLBfxeIWlVQBJCWJ9KJnWx4O
NfddHtjhrqrXH7DnH69HjiD3OSVo+YdWdVfuwBuYMUg/U7/rakbISxCZoEQV
SDAHYg3gsYCbSVbEdBVs7SRjf7pin81gsp3ha6+q90PgpjAkwAqVjiW/nQ/1
7yYO7UXpfH1+zMe6ND6L5m46ljVk78mE5el7Y6XlNstjwiqf3TcnbEypBjt2
s8YdQDGOKsLU1d30Pv7I+fGnPgG5ADWbi/UmGyHubwR9BhXhxTW4oTiLGSuN
uMw/OfyBcmw8AM5uzTIPjufIoywVnUP8owoirPk+d/QhGlsCmtsFv//wEsYs
2JHwSPif82zdACZOzwk8nsRgtyusHIx4NWNJVMp3sZwh3zJnJg2f/6p1siEb
z61sIp+6LBSUfd+7KU/t+J+vHoGWyZI1wIC0FZCeKSqZIh7kGPymGeIpHm/s
sHHwas2qO0VfLkpO/W+1w7qgsyK/zrWAkUrzZ2Yy05X68R4TzPMw4mr5WS3G
zPJinN9WX4imKyl9knrdBYZUQZ7am0ZZffewyd+Zo9lf+6nJbU+fKAb2LvGI
ncYra/O6SdGUmdFJlNP6svXtVzhEaqSgnvh12rZ1WiI08yRgZzzIPkvLKnCB
x9iJDSBJMhFVlH+7Y5ZHE5T52ywiNUJymnnJ092QiaB4GZTRPi41nNpdOXUD
r7Xfeg78s6zP8y5HQ3ZXNsDvLTGFmwO48JeQVa15RY15b18fB18FAKTjlS6I
FIcKZEhJYCPR494FOZGyxfQWgdsru75BqqZMnR0D8qneUxXcYVT7rgBNw+kE
qjBq4ppN0yhVfFSKzNYsoMJobSiyUxQ/DL+a59SivOMIAw+ueRxjETdlHxgL
j4I5Gg+KWBmAn+clE8llxcOsMN++aoICDcC8eWKtMSLswFHUniS0am23Y4Ak
ao/9sYLfgc+W4L4d4QRriGs4f0I4aqjL2i5RKQgIh2U5s7DiOejnT3ct4+r5
evZHE7p1mT6sHm/z5cCyjXDAh6V/6teBHelYbb8CKLuBhUhYFUdyoU52CNZD
xAvI1TTpTjW8HuTL6foUAXvdN6pfVXx6UA+dSE8y3vOOgK4FcSlSMQBOU820
TQ3B1vfsmehLomO/3ODE+okNMNIc842cUjmQa8127dZ7uoco+dDDZb+8OUoO
C8M9yYYIbFQgFZzzCkoXc9K666LR6ISW2D5aqIRnna14VZfUoDtdYogwlSwY
YwgI/j0IKMzJIyyckKYLcvgMPEebE7leRfuHcCQeK29rqkl+aCUE63Qd+4Q8
36RWCYMcihhCwiiSBeLT+yJdHkNjm8BHGJ7J+3scOvRd7rgLf7KZSjDfTqun
Wny+eAEDgiTUm64GJNxCMgf7cPdgwkpjtwRXVUBdoO/llz7nsc75QOSCDjbH
HKrNJpE/FpU2qjX0WPVrkbScyioZsI3cUswf+DsKztMSZR84FgyWwNJX364g
XHlvk8LfEhLbioqE4fyo/7tqGaCVG1r1aUF0vwelyverD/5VR1vtbZ7D1a+3
vbnqdAo90TMcitzweOvCKPFSl3oKoxCh/VghxGnzPBuGD3eMnDAbtmSFfJB5
M4ZaIsUkngRuDOcmOYCLd/Us8PLlja1SdpahrEJJxgkfXRnR4Rvj3EDMWc9A
iz3wX1SyHSh7IabY56XnG1g8ZppnHfvvm4gk7AkOTbBlcaR1rEtaBEaYJ595
DVm338quppiSOH0zt0tkdWYVLswGWajmGOqVfsWJQqaQdhb+jdLn+uVaVW8T
S80VM+p1r/JrlDdK0prwFOUrhBTR2iscJVLUHQ7bZhtzBHwrm6iQGyKynDTy
uLfCRCpv/U+SK8fSuZbxqUW6kJ85akwujBeceXwebZtYRk2XrXQq7h9mFbTX
oFwRrGtu/C2QtcW2XoGQXzfIyg75s9W/56xMmRVkBaswC14U7VUvshgoBlZj
C6N89EZw+kfzzwNNmNXOacVMhrMDtoi1eVHF8eDm6z9Eo2Re81JgZwcvutJM
2ep+clpNa02x/n78h1maB4Q/XJHkmeQeh8CBD5e3+YG4N/vx/I/y+4W2GLaX
Wl7qlscU1uCv1ug5dTXhlMk7Rfmh/DEKQCIN26ztwt3lWU24dfV74hesdVbU
QGWUU+cP7j5GR4Po7YC+xzTHWS6Td9dETyHxs6zLRaO0oeAov4dPcQrcj/Wp
JZhopy+9RQk986dIf291+0Cet8AfJDiSKBN052dT4aX5ks9oyC5qui+5H244
R4D+UZ5Q8PIMMFd6Z/6GSHQa4oVuxbsrKmkQam5wV+B6T8Qv+WcOpuPK9BsF
rOMPpw1i1ETb17F5LGptEUicc6AzJMX7BilrsLi2rUCIQrrVQepxZ8eUhIIa
u+8wMXfzA0xmB9Gyr+Npem1NXB451callKhUdGRNH2wHWL/KKPxet2Sxrob9
TKh/Qpmdo9SDDxeNncBMD0pTiXRZsPOjl9eXn113O+dNey6yI47RXM1yTf6m
pedk21lLxd4nvESS7J/AZyYMdeaQ9BQWY7hl41WiN658uS4hOvjZHRqoEmzN
mV0b/Q/OlFJ9tdgLuOku558hclSXQmB14c+ui0Nt8u/+34feIAvpmO/XJEZS
/ooK23lXJFmgT469QBtoAMNb/hKNELJyget15z6FIqCy3aDbpM71xW3CzJEN
THTn1d8tRWDVktgCPKJl36cpBGnUNwWpSNKBMRLXEjJlUrfLSMgFHZjMsALv
DtgWnogZBXZqJ/hxMXmmQ/zbVqZFMbKAeM9ZcSdXNNLa5rvPe6G03FJSkjFU
E+pN72gTRn/FXa9+wAWL6FzH1Lsm1+O3pQNrdiTSGB1M3qfHwcg/UDMJVugy
w8QqMZv9TuBXspepXp2Axsl9mhjWKla4WrOTWdfcNFcB+G++/muMIFwJeO/+
Lb2Egi32OcK4La1PuwH6iBpvmQdVVw7yHvYeutVYAKD4uRt9gzjyhFGgMDuF
8lAjWbI9fU3SiSSpxI23lbXR3KPPXbc3AiXJQ/l4sydvXuNwScyM6N5pzde+
S2oFYBHhkr6LXhKg82O0ZtpTE51GzEiR6gWMXhEoDthIMQc7HjbJwDOFDDnm
qjE4E3dLMUeW3wyPljfUt5gEwxg6l80vJTIf9NNdoBe82dTBt2IZgnO8kYZh
7wBf5KgKGilBVJhgGIU37xjRWXWnDWt8MR7rQ6uW5EPqAnSvWHjXAqTUKERN
6k8+9fk8k6ljdKa3U98hAWUi1SJAR27jCIPpBs7H5uWGY0mKYZZHSIV6JvA7
rIy06VmaOWW73bTE/gIAKjYb0tJWoLF5oSeN53NTaGhwlR6Aoqi5EY5yRa4u
Lu6Noat2ZpCnH8eWGhkSHTwp9hyh0oZTpmw0NVT5NzSeI/qmW4W56DlgTNwg
MbZ0EsmGq3XwKY4AubTVEmvImbXe6gCFuvmDm3Q7TXZtV3nR613Jq3WcWcA1
bXd0Jho1vnEfWEDr+IPpy9DusWt/NDg4KHMGtkP3zYBcNRZJ3l/VmyOsebOY
zt53K9SyZcokE34VXRo6V55bN6yPfSsfbdVIUqfS2gHkCvb8JoWbvdZu5AHS
2AwlUFHd2409wPo4HZjQxBiQcTzZND7hOMJDk6xG5N4jo0Vy5jSl1gto+MUr
48E7TrX4m88GvZA3yhS+Ltq4QdxyJEk1MJf47sTZFu4uyXgA/TzAYoxJYKA4
T3f8LpZanQ2McgSNntN9MUuHTH2MrvU0IVoqMEZumnx6eOnS9VjYCuzYKGMc
IMYiY+Ajf24e8VdeAQeGh0tXDOHYQryiaW5I5f8wYXR8DtzK2t0mW4TVBDM3
PpUpxdE6CCVX26tDbwECan09UtSiR3cVzx9VE3XFilok/+1Tr/BYbhi0ChVX
040aoJlpxoWiXWkzfGUO9iJFkj8D3fNKSeN6N6+LXsxTASo4tmM0B+kSmotx
ZpXayyffnReefKOgivHEqzOh0/882TW9f690ZZolola6l042/hHnvG5PQjM8
Jza4Mz+NJuQk2lfyMLuRzfuvnvOkh97CzpkwaQHNXJ4Zy6YdQeWoC9ywkA/Q
N3AP2ySdUYIekbLuLJODgkSFx2oOPBQ66w9Oo45jaNliPT45l0mqA+Vy+x4C
LuTVCg5BquaV7PCMGLwxm41rtyAAkY5IIUyd9tr0Fr+WCKTqrnUHdjki0z3I
01+oMW/9oirkXKIEccOc/T5nMLgnoEhLd43cBDS6EiWSxZ3BaV+z1s7O9Kd5
zA6dl7hr0Tc7lZCQ5kvEyB+uDipYEjHWe2ARcn4lXD7EiVk9g3ZnMUaVwkZ8
f5PIHuhyPCDkdQoipwdhJn9MyMomCDBuFfoIA+NcPDDSmqmlcjA1DpIMCDJH
uKuGzDMyfnDK2BgW1nWihLxoqLKU1SXYX3dnVurWXThMaFQhSA4qu4kqqj6Y
zvXwztaR1+Py3Ed17JqlFq6ugWQoUh2llUsklpxfZx8rzxuZ2iM4NWR9ccEH
f47cGHMrlsZKEQouNrd0uxrkniNLTwoVGDUfPRmYILhashFIVrPAVUYg7cbZ
VnDlmrcoIzAgUY6zkmyox+wlv3YbYw4lnV5p4xVOuz6vLp1PCICpy5aaoctF
6drvrQI0gXj8pMpolNYZAHfr16PRPRBur8EDBzf2hjbevzGhGwGy9GuAQ8Fd
khscPskoQ9vfRVQ6aocrL41+BSeE6E1ZDvJVGCZcFBSn31hvz2CAMrZOS52b
DqJHi4ZHXj6uY1D87INZ0/2Z5vUl9Qvh1lGcRpQP+BA8ppofi3VYu63wGXIw
UQmHl3y+yw1L/TQ9i0ZSjg2vvd4v5B4BkHFSE0HhIw93dh19PrKo8XprSvvq
E66kAvGnDBKEsCMDUjB6pG3dWzKsQdsUixSqex7dBrB+17Z9NvW6HuO21FEh
ga+qQuJrTxuQJrax+qZCJevNjyOyhddM6JyInQjypTjX94zIcsxr2IIMEfuV
yx84WTue6ENZ/VgwfuLH066ioI4El5d58/iNivnAmPxpWZljwR0XvGiFeRBX
B6eHTFdQqHUzixGztmEHxKfvp8zEFVKVtXkFdDriuCRzWlchXhoYm4VF2sOK
gSIkueXiSpuXoAVJT1i+ToRaR4o5pO/9DE07U5T43i/j60zLw4fIP4tmeqkj
/TQxspDNTRNPSGt7iajMq2absHdRdbCtblCTo6VSOLcItLQzGZJH0BTL/uem
ZTSXDgR28rRTJZe8oAYFfwLKLo69UirnHhSBfypuy+iZ8gf6YEbNlBUsgb/J
gbSkMTK1VIFLQw8pv0/3rnBxPFwNhWMvO8YFTOsn+NKrc9CPWkZrbADFYmaj
0THTbp0yOg75bTVZpRNC9bUAORa3CqJyeOcbXguy2K0MNNDI7Qws1C2rYmDS
d7zWjPxdiaIICWDcjTw3QsZ1g718WMR0C2tklW4LuK23HxekuWrLPYSyiW2w
EbTDJHgNkNFa48eIH0x4NzsOoOdzojDopq4Oi49J5d+DdiTRVw1XPsNVsDJ9
nnjLR3/QvNE8kEpq8YxjW84rwLnGyj7EeruP95kmWY7lq/9ywsTt6NnbpECY
kdHomV52mXBxacxJAc2gMHI/2TpOUWXJkYMMIGfuCUGRStN5HOiPqviMqAwS
Oj25vsiUDEYzBCcKPM7rK76f3xN5v0OLqjY8T8cfNx1z6F3DrkSxiE6fsAm4
FO4uNZ38r/Bp44zeMxsI5Sood+D8fyTQqzRy9uopzmjSvUpVy+jjL/cywtYR
rfg2ngr5ln/SkrD0WHWzgSY6Prl+lDECA11gClWyWJ9fYIMVRr0nnASGV2p6
XXPrL6M1tHiVs2jNmo0g7XmjYc74hxar3mT+SBozUCLWiZQkwAZIRRTkdxmc
XTgVPBLXyzpWRlkHduzBXviRD+e43SbvyLS7IPYbQkEoXVLmXoMOiPO+d+fV
ZgQ6nI5Kds8sr2bA7HjG0XYQ5G8QU+3UISni/RkDvxaYmUimmKvujxSHfSNg
w6cY0iQJv2PCAIbM84K3JdeaF3DUaju0V+Z66AiLO/DwcaAzCBrZwlld7ciX
kLICymCWGIdsLf0HGyd1qlXLEu+RmH5C6pMLLVfCJowk3fx0lGbCyatqN1Gf
ij9yxraFimyc9hcYJ+3dczGtBTiFe6QVDSwVIiaPWOuf9WnINmrG1nVWGJEr
3QnBvEv73Y6Ns5uIMqMOvNLQqm9Ds5eGQhowBs6wCcPOrjLLCArIx9z+SI60
EyeGrqEjb7eS2etImiLXLK0u5Hpd6u+q6WemlRo2OsM0dZbM83+g3Zji++Rf
Q0F5iZIH0COqpEziK02aIg+3Vvz6bl7h4vyQHtb3PsH5hHqY5Xjt4ZOdsa6u
pJSoewQ7O37b1//PsAY2VOGZf+PenJNgwIA0z1iADF5gfC43J02CmDbtIXrL
Qbu1Cs7u89VcAoz4YwnDic6t2jUBdfiv+hp3/bC1CH4oDjUD7iKzO/NoRSJH
SPvhrmNvXG5OL1Kxt0hF8MiMYd+iwvGRO6RJCbELTx+cmwtgahCcbhHnc1WU
tmQrkDlCAQ4Mn0vEaFi7lnFC1YKyWYvbrHT9G1HPPl7fn0gpEnBO98XSM2Ka
Nzg5hxN2rrtpU23fVTYFEsmYhmrxcB2zxK8Idrpre+y6UI5Fu4EEOlXHDE/q
1gqvSnob0xW0BuTrXxXgjtupQarvBZigI8iTulHR7LUe5RXh4cfLg2Z/2P/U
Snkm/0S0kCJYwIZrOwGAj9jFJJnNJcd74l30ueDDdRIg4juxzR2c7B+vM30X
Z4CvrgmLxQ9sZIlkEZELXrmH+352OXktgZ6sf6LuirzHJsdfn+/72rZXBF9e
krNdMjGnFDf9k/DUM5Qi5JdeJyqEdpxmC8BCqhJ2C7EVcvMZ900HICVHwgGq
Q9AA9IAHOfYAzwuzZLRLu8SK4bz7fmvGK56WYJ1z1Lv/wik/l9Ies06YsBWE
gFfPLnirmzeVAq5v88qS5/lvsIE5Q2YSMRf/SRSxi1tV2CbSiTBe73X2nrlq
8WI8O5tz2424R3GDGnpVYfOPLQJWjI5ijo7f60B77hX0Xv+N6R0oN0vWpHcj
FP0wRD2Z0Y2p4212i4+PTx3d5XKCS6wMRftAIElnc3D1bEtG03oT3MB0VGm4
OeD1zdGyqt/UW3fLTjEYwI7Q7oG7cMXbE6N5AdXJhQx44GhvrRZ3IXBYnDa7
BAD0bpZdkOxhry1a1Vbki/9WNsi9ansUR5Mjjd8URpvHx93FNM/MvTwDA9Oz
58MgM6sILWgsAgKE0IsCHUhbQcbeMJqJC2it0j17cCVZpd5n4k8acY4k357e
rCQEAZbOZb5v9KhLzfFUFQ6DE0ex88Hms8/UG/fFyHx1a7oUBrk1coJQg6Rb
H8omTgDr4EtTAwx2Z/9Nf2xPJYL9eM2XxBhUjI/80DV/BBCwsSlAwIcMZWiM
Q08FK/05HOa8aIlHNqfXZeVV7JO9sQ6wEmAMVhq8nQvPykvt8HgWh2hIlhwO
A8Q1PpWlDCzglTfniYJTGhHQGOrPrfykWe4vw+fwaKv2OlBCrFL6ZZzcPMOf
CaV6Wb6hncdNv7D3jB3ZgESDoY7ZvvJg/Ii/tN4KSdESAABb8VkoHcWWTi7t
tBzV7oPSUDbPwGvOrxOWTJEt6891RzLX5Km6QfzLy75c8+zYVLIkVnUrEpKy
3p/wPlrEck8yvkCNsP7TTTZyPy7YdIZNt5Zxa2YoI/HY/YRJ96Jkl4u60rfP
VzTlQ37+9Xlga3Yw9wzK4nzQMSgfyUeeU78r9FF8gRs6BZkgB2/hm5F+XGJN
IGAasIJFZDsAWDxvLtkA3fNmKuAREzTEqRItozQhkWEY5981JIpRksS1RjxD
NsQH5CmvQ8mMvWu17EdwbVpIsl56gAzDyhp6LpFhMthBxWTxDeECOTNjWhBu
7qPuakVEJ3SlnkIBiUm3KNp8Desp5Bi3lcme1H32h0iEiA67gT8segWrjZK3
KF8mWYdIW+mz3qWaWLiUvDh2pjAWWYVfVG4JHpCFtz/HFO/virCyE3iKO3E1
7dK3/tU+NjpcRAlfy6trYY8mnU2cIn0scUrxosSKyS80eslyddKCkmo2miB2
IdSEwLacZDdyViTnIK4inTIQdAo//2W6+0lQl+aNYARF4IRJD/gWQ1CVQcjv
rKPEpwxl/U7DLa/2OF4OdVxa96iX8YXv2Gyknw67swmGIPocEE554WB+lQdR
pylP5Yyk9caH7LYwAYVFaqO49eJscl+x/wTAcTaR6preSN6jsi5QIrv55aY7
bBUiSZW/E6m0LauotDhNDef/xxy8kFnhXX0Tkv2x0u/4hiMIHatQhynrr6bz
i1i+Y8voQntcGa/HKoCDllOA0geLEz7Xc4liGbnK1GgEu2OsoSBr+FZcDVXQ
jbOmH70wq/UdhrYsAn62VH2uyhpvmqvdE11v4RvdLqDAyxzq2VjI+46fEJj3
FGFeMYhZU6ZDPQeTKVWcXIMv9WAic40LhxkSt2Y1himfpC9ucaZmuMffHsYR
cOxd5/eXatfiVM6bdaWjG2M2oE8fqp6Gx2tJLmO/UxdplzLl5G/iYejL99I4
qX+hLlCYmkEhVZwUqDqhE6AAJLqSShpjCKbpdWat50el5fZF9DAZM5e7nquj
sBlO48g6i74Ts91J6M1tj6setGUuQ+P2Sq6/AsB3y0df47J0fc68z5hdN/9V
Si0Y2oL2OQ+8L8F4YZ5Au/aKxZXErJFUxGdEMWTgP96Y5Hndy6Fuc1WeHSRx
CZ6hzIE7weqQK0p51okfFUWnDLSSlcbUzAJH3ttbJd+etC1+O1cCH+gm0Id7
9vVq+FWcYqkkAmqAlB4ODIS6LFUVFviHTTXnWqiTbWrAIeyOAgDD9FvcwZZg
KyLVHP3simihyivYFzGqt+h9mRpBunXuoI6VTupkqVeZY436aNRBd4MQZvBP
sOBHjjhd8Dp3ny/vIVfslP9KY8+Q6ArZma6zt1cHyCEjIdfjNxbRfJczL+Cq
Y6V9C/yYwAcPDN/48x4yYaeJWix+moDJwaBJu6cGCVY/auny3+w6XXgCCfLi
qNEzTwMAiAK80sPq+QfxGEY63N/5SZw8Lrql5xp0a79VQsiOkOLrgIntRNXu
fTPTP2GlxDU6ms7TfoXEEaqWjHIWoiePPzsNfQq5Tpqg/Vvs93eLJtBXUbSo
QgMQ95vd3h5fcUKBUBIZWdgk6fMUBpJpjHFFBN2Ds0rC+JGUPvcNj0q+ViDZ
dhtkzy59ZDndSFWUfIRLRWRw/5xHmZc7PMjrf0+MxtooDNqssnHgYQG0bGmn
zob7zn3V2eF9FfLpWCjCESR6SlTfM9cGCXal3mGgUkJr+lgPvTGD3G+tw9Ms
jTb0skdwV5ON047b74iRd8kRm03iMVHH8WqaBF+9nfDJ0aH0HqNdqwMbPGmP
/ILGka5NaRaHxnPO3q4u4WnI/s80TajPXmClPVK8K63YrWw+yedpLrVDyBks
mwQ/go0ynwLa/5/8XkJfjqYpX5SP68jzrNGDm/WXUjrnrocHVEctpkHsZIQj
qGNTr9T9iijfyrMmev0h9+3b3T+tE8kZkmhxmsqJ2btlwxJZrkl7ETs+SBTO
HpmNLvw5f/sfcsX7oWc3c36Po/bVndWK18skK53xsXgvY9W72QbNd9IQ5J5k
SuCN6wZXNO67snXivhFB9IwR/1hgnYOd0VniShS2mV7i5r1tVTmflDM3GYGo
vBSV97yBG5KMjFQB/y7cJ+wHlxnWhmIugEfAeEF1O2P6fK4OXfgfzm1kj03q
MnD0GsIxshUfJj262x5LuOPccxGc5QQOvv/TlOTBBDAqNKbh1yQNYFWh/cSf
xtWZiJcFA8+ikRCDURf8JO/g5MJtRjnX4c+LW1bh6hX4K5R8ETearyfGlS7F
DlyztEPFOcL0q3Nxpc72uwq7GFBWv9OkTD4G+suzow4VRfw/wk6oUPj+qTzb
AKo3C69+qy4I06kXZ3TQiV27flTBJfkvdWp7yhcZJR1601eBAwvISt/FqaGJ
zXnWEdjKjPqRDkWAKUOA9qIAMR9Ybwg3nzL5eHt8hRFSCrpQkcW0HosaVk4w
iPP6U0eTQCzIbCxoI4FKJJAIP3s0LhvdKeRan6AxcGhlQSny2tFzku5om2nT
hUe6Yhnj+opiQbWyKiuk/qBH7VHe8OPbKR27w8EjtuiWEljNSg82c3DQ2zTH
hMoAxmOrxcKnCVEBTfKI3xjIN7ZmG74wHiIuLX5Vpy4tmmq8TufBepvvaPzB
KdvtrwIVjoO33R8bY04T3pZvDAhaTRLqwxLYGO48t8G9DGInnB/6emrGVnVg
FzYQCeVgBYYIQp3eoJkGFYOx7jfi9M47jiz9pbctoH6yuLPylAExq4d9Kr0H
sPXJ+MRuX40B4YFkVgGTQPY8R5DHnc3B623g3B7PhSmZqeaSMQ2e/O95Y/de
iurnWJqy2uD/U4soZre8YXKwvzo1ltiwTFFXI5sZzYRLkADqni+9/DuuJZdZ
lYELOuO8/VeBKrWRD7Qz4TIOe5I4zdYkESdoWkGfXkBmIa8FzU5agBM5gP0M
N3MLS67mJ0yT2Ry141lN5b+Wf792luNQ0jPb7i6ppa1eo3wrEZy8K4arsA4+
P59v7nadWYZJLrBwh6aMtcuRCgtrRqamCfIVhq5U5vhQ1EWCn029T1Oxv5fN
Fu3nh10p/I4ZI8yWQ19kbisV2I48ZY/5hgi0oMqky+Pf1DXVwvBLrDqAWhgs
SauHtcrseLB5FaeguEkWpX3C3sUjThYyLSKlJBjf1Hbkpr/kOmBNMIYtz8A/
y4KG/Zz78+QS+DQcwgKt1yj6kX7eWZDYw+zKfktXO7F2lsArImJkGrV1KCK6
U47+LeTPXJIT3rmIjr5nVStZyYbgeu4Gqghxbjopp8LFWB22n0ckscQ+rD6O
tyTAX7DcUxi+r6meVwIjBV0Os79pXZoNOU7S0ar4fT2f1PymasWNAyXZw3oi
A2h/WhjF6pnV7Fj/It0/ZzBMdPXtHjNsuG4GCuI/4QyuPdj+iAKSMq3Iy2DX
HjsWPMkQivAetgN8pz//vUJDo8IOkzuLk/P5dg0xqVEFHhEhBVPyTAgSrXS7
TKmglFlC5zTDaN4ZdsXWK0GF2TOgYl3WbHPaKjXFtLgVlDzegyoJ98E2V9iz
/kdsH20H5jdOqa4DTdH6ZbPbte7IzwFlI9RbpR9F7vh5IGqZIut4FxjrPEMP
RXM6537/MssPzoJkEof8RJqHModTSeYmWAs5WNbohvSS0GHOfU3z6ePZ6Kfa
4LGuLORnio9U4GdpZFtN4I2ty/I2p4hsEaiHWJkf5eD/xcmcB3Dw2dwrv0bp
MByxDzidVlJyqNCdbcLJ6sIM6AXqqJH21OwcVb+7L5pfo/4jA33r+sd6RDwm
lTsZ6XC/DDtlomwgUcbZUp1M8X3xt4PgcNkn7JDY5FC6+vgr1yNRm3UuqMEl
vJ6fVC+KPsFT/0sfFpN3ZXibYrS0cZIlYnENnI0c6e6bCLtetsfr+Vew5m+D
VF1v47Oav9q/0yjG0vJ3FAlciSEWy7S4g3Wi7KeYgDUClmst40pRnKxpdDcT
aPHn7VL205dQccIzv1C9yeXLY8CjLB03xdBd3ZMyWCeYNDBFDMluv54E3Ivz
MzZqo+L49ViKRzHQK4L9o7yEMADd3XY9Eu7nmlLcQHR405FIpzoOdGUu7Rjr
v7z7ooYEtRf5ruw2AaaM8/xaFM8868LPVb2H0LitI+k5JdbYwRarS8zch32u
jQt4CNieepWywGbe27uM9LCo4zsNyyuEwwu+PP+jVKz+eVccCjvo3jLeu2wf
lYEvTEYyrNZbYfE8ToCedsEndu2z25zC/y28D+stPw9DkJUGLPxsEr00OnZm
MXOIdm2vXgpCxJgLuXFbdrRS9j0/8nWu3ejho2x4Ju5mwBWH5JTDGy7e5vNm
GTKRMLKGyr5fqdfUaQj3ZfMEUEgJoQK7loPGBw68oV7MYFuheKRDkqZFyuVu
lmxNaim9gkO5VBKtPHNM7dj1dYys6eS48AMRfJnlEbIXvDE+qDabMAhCKHKN
klkYZk0KfQbVL7vNjdjvw/zlh9gSnR/vXv1KjDH2O9tTw3e0soXjouZIEt+l
mFOxIDE1CJnW2d2sHJ4A8EK377KK3X8nGQTKA/bSx4qpPl9kGF9weAExBbFM
t2up5yZgv7xYcEM3JwGnFDtEfU4yf4L5sUfYlEIagOLcmYA5aUIR9kvl1o3Z
K+Y6CY9TeBLU6TPbgUwtIuCRJAldpMeKJMet8MMRvjKxwCDNXNsblFwQQ/ly
gYxgJM07NhJqYcJtGZ+6XkrZRMOzXYLt6Yubp9vMX08D0W0Wvu+yBY+ZWgDh
7vXfMWPRGNg18vkejbdWUURO7DR+Gqka8GsZejx5yLxFkdnavzLwUYOHLURz
C654YScvp5SoCHCd24QTEWA7lCJibzKb7WvPJk+LsyBZSBmBAkgikp42D1M9
VpkzGgc1G1ZWZgz/tv4c1l6onZG36acHzEBF1WKGrvjTwewpUV4F0I9Z1BaY
EdI+aXDA3GF1t2UYgPinIuPcILDmU2NXjey2fb2EMYYO98LX5ms3+oo1WJ0o
z7v50xBPX5851z7M/NFFmdioL6DBGjUoMoragw/vQxx5NvFGKXExwVJ3qCVh
9PfwGEmtvZ5FdffCsH2ibVeKNS/aatiWWzSxyV4q8ApQPEaBme1MtmgM/VYx
Fp/XGBuN8WA3ICKm0FjvBv3iQP1PgAjsW0EdpR1nTswnaM1iGrQOGj1dX2hu
q4WhhVbEGudE7w1FJu32jrWgw+HsOo8T3m9bm3nzX+2azTLVLoJZUFro8CYc
7FP5NceC+RYkqErWY2pWv+02trR3gVczYtL5EG8ajn4xrMnNy24QJAVnOmrb
zV7qbTjOwkxRDQD2IJ9qkUbAimZJgAVsveVqY2Xnw5WhFPHEamuDphM1ymAh
q8goZEkIibpvugfOzcAeeYbMGQnLbDutkCd/Acdc38v4ce0DiFnBw63G6Inx
SvdaehSc0LnRtYV9TbOvS/hkqNJpIDDyD+y5cx1VWf/8ik52U8vdySw9XrHj
fGQ+84NxwOifmTZxwpbIoatuqwIbwp4+D5ty36OlEx/Pvv9d6WGZAswk2Xqn
KZtcZWtnuHZ7nUSGej3mIQKV2xistTK0DQAAlq+FJ7GtQ0HLaYVcQmt7zHUp
XoogDyKddtUYYpbRW5wI/q5F3MCo08oiPlqTMuUqetfEzvGWFtyn6ebPfLIz
K5Sed+diOayeajcQ/+NCSK9MRRsmdDMGIPp+iP9wEA9tR8wIfhLLtuDp0dYE
pmrViKFkuTEPiuFjacVi/g/9Bh2QSiY/5FleGcRjoubOYqWld9qR4sXsJkNW
6E3XPT5fRdnvzgCXy+zNfa6hivhQ09qsXgsBIkDhqwOdOHd5FQlw8c9dmMrV
zH4Z3LLApVb5fDcxaeq+eeH2c79obqKQZL7xDti7n5kkUWxCH9E+gke4HfRs
aJPZNvZO+DgpyK0x0AjtOvuOqk86i5ovneummtE6PTp4muSeVeTeuXvH80Uh
lcKK3LtsWHFSbEBZFhhQPwbnYIviggDKEykRfV+AeAB3bQsBSi2JbbJoP5fc
a6ORebP+9dkTtubz+D5mbJP8Lgt80VSFFGr/wgTn9U8hk1z1VKjhIt/RDmm3
V9RnFw8zmUVIeoOiBQcpSaDP1nWnX+39y8/czTaGBI3GMKi5fxrw9572E2pO
hRCMiY1lgBklnsM38DP/8b1cvEucye/WfhqmXGhv78fpaLXc6wALIiUxEk8M
D0n1vSYb3/N3JMiB1VdmcCwx7Fw/9d0rvGt8K+L+rS0lcjIjw+WpLkWgt5VC
MmOftLhQ/PSTjBWyI8EHQrg3OgDRjvYSEcpNnW+PawQYRE+unvkB1KJ9WtRE
7rlqS+MmXGYIjchn1heR0wfO5X7Sfv8ajjc7nhO09KpPKDRiYRUqUOVxABpv
Y6wo1RNCp3m5nR5kVyrbIDnr7XKnG5XHIUfRYP48r+zCcOBVv+HD3/9HLbuJ
UwjUILkK73sxqOy7u03hfwXdIYZY9LFKYkvyx/EUkGdjklx1JVIkT6yuuJJ6
qEoG4reK/H0Ixh+alcYFz5AHRHDBnnrI7e/SQVqbM8UnOkSs3u78+dU/JJHI
uOZJeKkTi95EffyrEK2DDXDF3lIYOLQqPMbjyDdZD7Fwaab7ZPzl4XWDn0xM
DfAiFb151OKme0zIXxvK1/j90Ogf3/p9kb44yrV6DmITCs2F00cKU5Wj3rDS
o6XqJZIIXI6T+TKGmaaeCqBfz3evBbvixauGyWGEpmulIA6hfhHmAOxRF9FV
4Dxs0MWP1JNhw5+j1DbwtlqXgkjCupKNm/OxpmEq9qFt5rpa7mpSDOMU1/IF
+wv5LFJ8bZz3Vx4xRtKv5B4qLRjuA9p2sqOPshLtmWNxEEbtJxkVVJYBzFmz
QvZ1j51LDCTjwErVHlAaSJ4DGlQFiui+Mpy/+HlnjWxGG9i4NzjQbOsDiJTg
Zw98qILKAix1zSTg6OoAYA/fvauSSLRf875UZsR6PqqF/Wn6z2Zkf8NLo9Fm
tadSeKN3dpXVkMeTXL87FQSy5tDjTAisfpNQIh3Y/Kv/RKJkKSWGEE03wrIq
zTo0iMVyqo4kl2XhdHcLynxUd1e3Pb7gyrtQz6Uq3LMcRWj7a/C8xY8ep5qm
cfkJHuzboCpnMH3kH2lkYtQNWSDIm5BICFUHKVhoFtw0K2mWw6P5lubGom7v
Z08VQbLTiao69jxdGArgCZuQLsreOgDF7kC1psXqI7dM7z1CkOlYDpycvpgI
18TQo2d4V3F7WnNzhLdqMTTEuHzXwUnFq5MneLTLtJaXqdPGPSwxWrpskC07
hdqnnUl6/owN3Upnkl583BJ6EuNDdR6GrXrxKNYxjT1J71eeCY0Wi0Bvov2x
ESTSeOFi1+Qce4fHXjy2ooxhyaq2srTU3XSGTwE/cjz5EbWCIthEfFvtEVYu
nmRwcH4vm4dzFMhRt/kHTQTcGHPdwQeDRadoNak9EUfkFGSwxasgCjwl4NcX
clzgHfW1naBVsFZgIu3n88iKtJg+QjEXZMVSLrjrfSIQSAHN0NbKfe1I9Xff
NaocQgn3B1VLNgRAUzss6+YYgH/tw9wXSdpyDDd0seAoePMa/aHK6c8peslA
XpmFUWXD8q4GqNs1BVGBHDnBmYYZiFAKY7nv1W7XeGdy+vW8yzmoa5wRk6Wx
sxH/1xXkVWmO+oxZKbNVQAZqGRIUAfSQE49CKghXo6/gO/xOXCR9fuD7hey7
nkCf58RApVVvU+A47mdDu5nqrDzZHltjR1Av35ijlA33T3HgbOpIMzTCitop
O6+rWoU5UduJaOKwbWu7mQplclZXt5FavY5mADDm5zaMpTLhYaJgdYpwdv8o
5clFE8EEdRo8lwbFNBceuoYWnIyt0PvDpH+CvOvoGsq/Hy6Nshididi3g62W
niihP3uTf0pquHv3adSdyhhtG1RSBW6qcEYDAT3QpY8G14GR5ke8JXLJWpbL
jQNLrS73SOZ5izOil6LTja/W0FZY+anO2eSS/m7rRq5XHX73b7jpITctUkqN
n0Usl0qsTbEbAkFQBTdcN7qMoWeU3BD/E1XV3DiRNlLzdH4Kinq/uSxQSrrA
KfjrLcIUPkDSAOXqKWkRggw8hdC8ZM7/Pud5qU8Hu5oO2yslUHPWcNY/vkPc
OKzcvmxb7uT7BfMBoihuRyr+hw/pd3t9khu26+NOAD1M/VYWLZ95mDgtCxBY
M9C47u0dSIO+WnFmUJW+8fM1tUJpmioKKTXrBMTvIg3OWsGGTWd4yU+ZabQ3
uzGNI//xtW1+BlkpCj9mDHvZ2T+5gZkARWT/L0vMnq4G1y9wbcGuPNRo9wc/
bB0jsWgM/Gusf7bR/2MrnmOWYXzH+g9VdOZCU1Bp5yCLHRY3qp5Pty5f0HvM
egSc8BK+4otChOA2+AunuJCcMXWReGEtjOMeir+9OGr//l4BKfbiJ++j7/m/
rsLIjXyYqiAQWXUWGqHLilgFqSC+Zt4VYBgnJHAP0YkxrTACkKxaC916Klre
ajXZORa60it7MijOybUaHEk5qnhv2ovcGqtc7FFQWRICNJIRF6vU13FaE14j
Ci7arw5tCK0wx7wNiil9Z3jaFWrBwUfnCUgEIzJ53Yx9Bd4/1pXuBnidt1nL
YVioXDaSzrCa12P/JtfbQ5lHXiIl45qyw29doxyBmgQgJgWzCbZcE78Od89J
nii8dg98vMyE1u//n+J0gteZllmgHmpC0QmO4BA6pDsP541A9dgquP13mGOX
cUcRuRm6MhN5PHVspZbhKxc891Ww2GqQ5nYxi4lKPbZyu6FaL+HswDeKvkKh
XSo4zpHtfc0f0SsPHK/zNmLOEiuzmHnBPZlQwxhx28VBolw3rnvSk3figYOg
e8JyprU9EFyJ2rBpyr6Dg0sFY46VIc9c2Uv2HJoBryhE8Lk/Ump68U3QSRU6
Tc4sFDCDBUNcqMcWs3TWAEMO27Rch6wtRrPru0pyYfDFZCKvrGtklBlGNqga
2WcekEbKdbhpPDy3A1VvQpLPX7vrfkhOOBGyqf7JTgEvr2Cxm09vWtf3t1ix
sQEUk/LNCwawS2Eu1fQB9y1Ys7GeuutHhjqXOyGDX5RSf019dU+OCmbkQMWE
uug+m46rIuHPBzfXp1aOw6ukfM5tNX9Sc8igisO67u71k7xMKjN4Ez9wFUp1
+EL2eImHb3qoHppHb9Q18iU/XNVRo9jUGB+LM4FEXTFA6jM388+7c23YfFEz
Wo2eDgTTUOeOksK9+V15lnMP/GY7byBUMY//nP+3eh7pmc+ae3EmGe5RnaN+
WdgyELgHUl9MGbbv9H3t2N1af48A8cSzZp982gJ60MU3AhtVnWS3zvhT+AGZ
pzBqJDsjZtbw+IdoCEe37PbcyFfzqz42auVgIKEfrwbclgLWUk6x0PtGCvQh
Jy8BkT1MWWCSL4aTqGGhyB8+o1Qx3MB4tQ241Rthk4cqDnDxGvE0cogjFHdD
E6r7G4OOV1atSDtDTLKX75ZOBA24PsDNA6y7PDzzgyvX2emKk9XFaqRaix/k
U3Jq8M6wnS7enOTCqYEt6WvHLZeOo0s2X/YPj+i+q5WGxTtnvmtfqH8znN4h
4KMiiRvnPHNdnsPxJgbx6I7m/hvPIi3kc2DNhAGwlYEIwfFh+Nf7q4a+kbsl
ZUIxZwfkn9ImY7aOGR3tCwFgpchz482BPkYEgmqqQMKAURIgcami0JkC5UYq
ayojrzNlYvge4/7s59lzIakTNxXHsuOFdBY+vvY0Ig5WWt7H+xNGIAGLI6Rp
0XZX23yRsyPbfqja2/rGwSQDzWCa72B2skcqD5TFW8XXufSd3oJgj1XrEQ9l
HRdOictbnruTVIXCMmNGAAleUXOX6BtlnTPSd3gcrcXPfvmywX3X3e0L9wh1
IhJJt5Ma36sqLSddZyMBaORNFxrm//NH7mghpVO0nFXZ3fWH3nDmRkSh2nbN
SxUZjJiykPsw8nTxpTsG0nj18a1oZnaFmCh7skoGMCgRBmDQfOngCIOZii9N
7D/ngCVsbwSVSxgcPdxnPPv0dwFLp2EMEtLU3M/fY/dzJZmAvv0Gif4fyH2B
UDEY87N7AxSSF9ZORjDIW0s4qWAEyfJ0DH771lz/hZ0QbLx6aK6Wn8EI/6bK
uSMpzSegA6mEYxCMX1t9P6rZbV9KnBmTxit2mmNst4TTny+z8zfk9TFPz58d
WNi2Gb3pkmGOX3d6NqtV1lEjSfZ9jyZet8ekRdsBfcxjNAOT4jmLx9P11K0K
QbteizNd21FCNSwScDC3ayOUB2DPsvwkC3V54SLv/1ecQA/X/GlMPZS4yc8m
wpVx8Myx3umsvyIfNymb/TpTYPA/VkrUBsH1Fjy+Ro37QacRJpqc1hQbetSr
u/w8NHGZmeg0tsiiiuRg3OfEG/2iSdOmUBVzQAdT2cmcLniub3XV7iwewa3q
YHdOgVm09MqW0cstJyNpCzGtkbV+lh+WRagx3dLOQXQbUKX/dFsUWmBtA0wE
oHSg1jOPX0x4Pm+QiRz7xvm+ePIizQUD9QKxFM3EIgvyaDDhti64azgb3e6r
wd6JZ3+48pCR8mVTqObF5N0BwPDpzPm6HcLrLanwyIhzrNDL2PapPfvuPOKC
MJi6CxvxtvFSGv3pTBGVp+ILFkQ5j0JkxCmf/uIX1yuICMtCaNRAPRyTnLPT
64y3Nd37KlbZpJvqyA3f5/waldvgdG4gI0+haw3qBIwd7rwk14I7+WscEcu4
mzbzZ/CoiUdvM31C+3fEZUNgXWGQLb2fym2gaiR7fzX/WtDcJNt8L91XLBmE
516/f2WOvp8VBgHgLvH0PAp2SEfKmHGISh3YSkAExvy0KlfWmPXSi8nTVg9d
TsH/b8+vwuhFLh5/AG8p5LO6ng4q+6nH3c9ZMA8IqHGi/B6V5wWcTygwmxFk
4bUPMip15ivavKYh2NYH69hjXsayXSrVb5Kp4IrSodrfKlhmY7OjV4O5nG6O
UnVMBYUwIHXrkFeFPzPVuWu2vX7ji6QRG6Z+moOjKLkT/h07YcBBSdIDfJE8
mVBVa2QHvz+Mg/qshwMK66UTceFR2Px82eWYdZMiBbfFJVHG3i+cZhX6Ii4E
Ioovon//QJvd/trDt78SwHMADbFvCRKof6bknxka5dwipjNLaNcNvmSOPHuo
Vk52HYRDvMHwzQ/nbotJhSR+KTKrGgXj20HWGozbLEprwOmP0KlZNLbu9wjA
/Xam+q/NfCsLY8X33FVLAevhAfhHN+ws/qB1p03mWhCg0xSxmiLyMRNPWrfh
gPbPV1vx0dS8srBrHbM/RPEEcc1TOxpcxJtfyTW0z+B+bKLIpnEe955DbgXQ
sBjz4vj8uJOzmzeCxcIn4bI6i9U3xNbvOt5waSajzz04rUWImuYYxNkWn+Mo
EdMxV2lXPEMjHg04+1r8m9b8iwq/Py2TjB+y/f0degcEmP+bw4QpPxI9CcPH
YxdkP8pGBP9I4+36423D3uMZNZmOBlHujR1CvnasxgsVTepML6EzMg7IahQM
Tk8ufxaE+BrF2QLqugY6dtxXCvZJG1i2fs5VbNhVB9rmVWd5dCYUTA7IClxe
oftWjJl/93VQFbBttD8TGS6OE73vW+uZtaEHtzzlGsuyL1hcWiCa2hhYjQDh
fNHE+1fIRCtpNG1fQfhPK1KiCypJnHtL9vIk5dgC9vKI+N8nt/i9LEobXj3m
6E3uKAdWVkbDPq1BwId9l5jDLRLefgij7TCwA2eoMZt7ys6iJRevH/LCBBpq
2o5QodazrbZb72P39aUy8VBU9PQw3eSSDd9TqvfFaRqpV3zQFkf/QzXA/2CF
RPjjmlu55erQ/pzBd6X6HTOUcUU/4Q+zrqBO/J15iRuDVBDwlUnb6RKeVuzv
C7anvSOT8BmvoPS4Q4GIiT+1tdcKLHayy6SoZg+hAk6k5SplouzotRJLN0jt
TkG3f//muQZmaY57TETkz9f7F0n0TwvglULIz7wnkGTRU4svhW7bjVeV4O/X
5+Q74QX6zbwvWso0ovVF3x2Cmiq3PpTNXDWKu/LC2A7DCanlDuJrrkmDzBLr
HoDVbnj+bQf5eupJT5eqmtrZO4Lz86mE0ppSzo2fdPRrOEiVBzjn29K5kNJt
D1pCbwlVVEdphARpVd/sEwYf0onJ0rV54r3dS8nM1+PgYsgGDHxn67bqAJqm
A3ZqtKxeRaerXVGup5USobO75yjy3H8YJq3t7f8IhwRioSSRc48ZQuzx0bla
bq28oOuUcyUzvuAJITeaL2NP0MPRBe77EXz9kGuhXdTZpSd3jvsbuTMRHbem
DmhTwDef+FGIr/aG++TYgsW2AymRivbKlLKLmuejLjk2k5c3a196XYcbWEQ6
u+RbhSAIdmuzjaQpvLDrD+PNo986bp4RAddRhhSn8z+hxWU8UGTkqCrhypFX
ScNw/JUs6OAt7/3Pn4SJ0vJqSiTKmOpyKfZG4zV40pWE0oZbUHkjEMowL5By
NXDsjHKCIk7KiOLW+opKRlTBvO0542LWVbaOxU11gtWAXgUADinwOMXNuJpm
ynKrXuufGZ87H3/3nU9GUL3WMGy3Td8sH6joknOlsaUjtHn2RJ47BpMnjV55
ltp/16x8Q2cXx81uSxOMCxpewyloXqqMbuQ8WX0bcosSHP59AI/5pg92wrwW
g5kZPr2SaiECPgofHG5e+zQs9pe2xcF8i/pIPuV0INr67afkuhDzzHEm+pdC
O9JlvCkrGGF1xqxl6aLNtMzXXzplWsHGy9l51/G1waDXJK0vclL157gA5eRa
t3iR5iKv+hUmBqDOGohYFAB+relQUnhL+jN9SuMNcKZbawJRcZT0ubN/y6Wf
sxnTJirffX4gmehVKWqk3WpjMtpidTSW20e4yjdLEgyd4T5CcOEoxgpOacN1
1ebdxrnCI9//o74cVhd6y73KnGrkWH0wATB3BMnJko1/Ov0JdOlJPkJlQDLu
6NbWs04QMOcAMJqpBBjmwWS72a3fqtsooTSabUwQVsaCqiWqYYGS2R3hGqG3
mA+77dUvKob/Wo3eaZ+UnhLqdHjtjLyQ2N0pjqxo5qSICH7AydDoqwngFfcw
XDGB21U2j4UMzetIqkqPpFdEETSw1SwL4MAas5PZ5ESDVeq+NuYKr+Bip/hW
vkhdXymPh0nh6P88q+O9MxDyBHd9srNAlcx71ox1QuH8tD5a7iNwx3jXSNAR
8OyqjZ4Ok3HnSzzrOfNIaKFB8tlE7E4p8Y5GXMKEvOPHg3gNxRd7iaFlEGlB
cxolGQ6nBV14jwiRZYVUMn4utUeEgxJ699rz1H4mmblC8Ju91QCKQWCwwZ9p
1nd8SFtWPh6Iu7EkEZTliOpLgyXPEv7ZrKpGkhrXBCvZs2FGyo49XwXwRDYS
ErsEIfS6I9kIlWhSWHbFI2jlpZuknO0tPo/iQ4fgyNBv72pzeDcpNz5gZRhu
VPXFtMSuxj3giw35WvAtVbHIuzl68DLgeE7TpeAnZuLXSClaTRaaLWKdxam4
r5a3k8QWVT7sMbGlCpq48mlerbVVrvXlr0xnBKTIvM9EYaEXWtV55ZFpOtba
+hUIY0T8No1XWA94d5ZrTOp93DZ+p8hiaCiySVIrF5+f+p8sHCv6+Pd3NBK/
pPKG450Yjm1tXRz6QLXxP3upUmoReWO2bff+S5QzAX13evQYasGAFjWdgyEb
dsFYjltycSMsjE6WZlvkd1hlv61eQSm9aXvg48wWApFsRUgnw5jIhL6yBrWP
hn+96rhTwncoNUtraqLZCptK2Gu+uIqAh5wguDe41liaBS4iLxfb4pDB0sl8
TdBBVj8VAhilIAG6Km2AWDMoOYuKQKjBHdQoFmXuh4LgM+M4kkCbZpOF+6OW
uU65mlfCVPEVGIB4/IFfIq8A/e8H0Svq/IN2SXeaGdh0BCqk9eprWpMfR1U8
RhiKrt3uj4UJ9NbqADc/Ca2IRuzRHYfak0yq3WpU6n+oYFoG7zIOCAfOSV9p
4DwQDt836V5xE1Ng+S+XgdJCJ1neXjGt8CYrq/1xPl5Ao+s2bBmgalquMkQU
OIoSjJLV51drmVZ2bYuOakiLM0eCG6L3MzsVzHyui0qn0zUMY7o8GNmQgUEl
ic93nY5eHPnvBxtuxIKeUBrH+2kYAmb4wGWGDT4pugVc35FybjVhGh89G8bd
lbjg3HQFugR6/qaQ/1hH3LTsidcn9HU3f5jBvB2BvEzeE6MusfNXeWhCP9rl
2rQ9A8CyZjVe+5wtmVTrDGq02SdXirTi0KI3DNy8nY1BatoT8Hs+4AwJYoTD
yx3XQgjiGz9TSWKcCa1aZQ5xWIAfoadX6WwI7YQssdHStI00Fa7ftnn3hbeT
myyeUD1nHuQSXFOKajQdkSx2Ocwq6soFTbm9lJvgaHXbUWLRCWmqg3uK9VAm
O71X4oHmI+Xpd19ZJGTh9v3l3zSD5bv2Qa+TJSISxvI26sHMqrENzmf8B5AH
i00CJMlWuUJ3lf60jCqRSOf+ZjhlImAUwCRonERiNNRWy06BEYZEIn1GGdOq
SzOTSZs3szWjZ65pWz4Jzce5BDRzTjFYONFCm69Of/hVt4Nh/X/sZF3vlwuN
pbIsQ6HEKr8FAl4lzpykp8SV0Cgg/3OHPsZZ2BFWky4+6rlhN3KT3wOtKEWb
MbnHeBZcsNxOre8ml95/9Te/cNAOPv28vM3qToagFHpJANnzzGrCbuuXfSty
2K92hIosLcPb8RQFi/gxLhrzX+4UVkObXsR4PYEVZxub10Ecw5UeuvzFZl39
nDLp7L9mWrX5BUqxGWBcp1icvhzjQdbTT07S2IpL1O085Ro8VOs67mjRXJyZ
EsVG5iHY+TKHryyFAzBmaS7rN0tob80vZIPQOPZsVt8Yucc8Dd2mEwMHy9ro
Cs5uV2cjYAGwMH4JNtHHX7B5uohmd2s+DjRAu861XL5j2X+Wq5hnn/6RikEj
yH779RChi0awdwM38Q4eH6LhzcEOCtREZ7ki5MpCqaODsYQXbAKt+W5Wi7pu
IB/mY1gSMOYVev6eNhv+1V974kI0PLCq0er4PIOp3IskgvLD6jc92zvEVQih
uL0OJ88PlITfsTIbvigqBrCQ8z3vHm/fIl8rtS5JgZyMbtdv0/Xhqm9cJRkK
O6mBZT3qUmVi8Ve18rudo/yoL/vFNi0k41C4D2yREgHmwaWoloni60/r9do3
Gu/Io0lTDVwhSUQeO3eLS8YklL5GFbx+aZFSxES6dk/+oCMEz2wgigt0F3BN
Mej48lEMt6Q29dBdjdwdfjnAgJeYtADZWqIpXZSU/V+Kvnd3ygK6Ocegc5vc
WxCC4vL4PPupiNytT0pWJk8JL0agepozwvyQJIAgmPmEGMCYuSy+tvovm6go
Ayn+XEzrY107FI/DgFWQNXWOJRs4ckisQmlbapnLiWcQLgCdsj4Hizal8GmH
slOqoZl06HOBKUtd+bGRix/R6taRl6RWKQ+gbcBYWSF7V6vG88QbQVrOU0cu
qXI+FiLIab416fhkLcTYJF6O63HeBBcCe2Ku83xJRQ+5XGTQlPh2yuG4VdnF
xxC+Y79kl+31+GBo46UHeKBQ7BsUdv1byZscSRElxY6fK6djH9S8G/wVBA5s
J9aG+FYxI+YEDK7xfJSYHtSndRf5nPreY+s6kUSKGz0liLuo3XQCf4iV1TJ+
/KIx7ka7YTNuGAnLRQS5YkYWNTHjuYYpwhsdepnIuySeYNmT0PIfL/oabcAx
cZ59BuP0HQk24rtCmK0fkQG+BdVFGNH/Fgf1HjkQrtrV2NX3mkZKjTUeq/u6
qdCE0kIqEk3umKsHMUt9oYKYYOTfS5Kc0J7pQWFw1ZQ3EeZn208/Q182mI3X
ei6aNh8pXk6gUXKMRT+FFiYByepNkKkMwkvyquke4PX2a4B+4yFIXcEy8+Xp
/DwZYx9DPlrDpFnwkAClCvPRhi2Fky0Kk0H1S/4fRAf3Lc38BCbPZ6yk6msF
7k4Jv864R82JmN2fGlJkLDxLZpJZ8EfY08my2psKw8Gs3LKzKt1Y4k2W6neJ
/vYK4NAEdvISvmPrGfnEZYfE8S9hKu1G1I/rdwx/0GH7OESXEOBN2PbY5wUZ
O8o7V8cqZ4QBpc+vJrjcDW5R+XQAiy7EWxKlzyI3hJ0J9C54u08zSG5hfVGa
LGgmLmT1Msmsmi5pVIJAom+zVaRo/PQ6d8XY7x+W9xBsVcT7BrvmhKB7XBNh
eZ+YVKrX+sCv52GIVnL/RdQN2j9jmH9i9XEFyHvmT/ltzpTiPEPHPDw2hg6f
NBFg1g7uhRYvLfCZYtzmuYAS5xkS6WY/XVXHhMDy6LEHxdUVCRd2EGPO9+LE
NIrPgqRFp7bmiz+iJ3U6KZaMgoGthmN1puYVxrd3MYmxarHHb+EjD4fFB9Dg
9CGJdkm98qlYXTVtg/LZtUPdFffrxhQyZxZiPUPkk1juHCRGE7dTlqld6Tfs
pZcH6ixI/zWuHvypZTL15KuCOP8mCpl8fmZp8s9jLFtbhr1wliGfl3oLC/jv
n0DJD0fXBcTFOIHzHFQ2gv9JqmOqMOWttxjeNJ1PIF7kbif0LCJ0oaHUNzCm
gU02vgXJt5bnLFqtZ/E13DJr0xaskoQEsCxc/jfpdmc9v1dzL96J3HZWmEll
9jGIKbRAWuQKs/lYcusNsugOm/0ANal5dHD/pj9kkFQHGgEkIY4vLolewOyq
uvbtVLIlyQwSiYkEOxEmcl8sk4RarkHAJmAhN/3clyQpNCRdwmaSDIk946r/
ke63rijiIghxYXL+qEnTihha5jn92eJAE4SgSvUHAaU368ckPpGWYb0S3ZbK
DcfIRQOHKhQKMaLsBVERXSyMzrIvdZyqsxdvcWBiGquwvyZtLL+xEvP3aPX/
p/U8pGYDEE+NoyBBTGE1eGPaVYQsdjZ1SXjvSZMtwT5Sn0xjSX8nGeTIMTdS
nXJwy5YolUQ4NlDKnyVZWs/FYECnvl8qbR27gyVAJaalTuVVsDkbjOKCihY/
mVwX1FKtgIIFYpj7LcmhUb1cutYJyCx9bipHKVFr+svhN6WFIxtHdY/cXO97
LgOY8Rbsqgm8fgO2rtkMN68MpgDK7VJlK8/O7REYgtTWUGMtguMArDuSSsR0
d15X4MVxxjxiyGtPKvmHiYqMf/zbcahryIasNIoFv2edJzcB/qFRdIq+oRuE
tBHcWLC4wLe9QJ3JN6zYSTgpnaCffnJGMS50x3J0G7YRCiyd6E/QFCyIOE3e
1gxqt53R/SqFskJAMhLbWsBWKIZFqa2G4LD87sweEHDUV1yvcDFuJ5wzqLrI
onT+cOMkAkT4DI+3daUcM/RkG8pzOPN0nPps8kzLbKraaqDMwKptj/YVmV+M
mLyOait0GGBnzKcHYkz4H3D8u4uNAoYQir+Ie9t46rHIkjIli8hpDaqkVWPI
jZyuh/D+DVtFswDxySJbIwDexfJmmYU27WD3BWH5Mk3QXAYDBtJ2RezSXyyo
uZj44rrkOKnarUeo6hdrb3rSfvs+B4Y7e1s7qb6S9WsiSsG7TUZX2b8p9/tA
eFeLAb9Nbrxca8twjKaVj9zJYtyMJqwcck1yD8ihxQwmeD29+sBkWJKroLAA
TKo+m+sOEmXnlsKJ/3PdyvrlW7vTKq53DL9+OO/5w36qyWFF4l/T6fd36oJ3
NLk0kXMrYS7hvPC5TNJWj4iAbAd1PNxjNlHvhCBZV2naGI1XUAx9nFShRjpL
M+slg+vP+3L/Q0c2hMBKdAb+n/MtVFz52arMoIFtOpALO+E1CHjJ8nNfLTLE
TmuQJ+4YnmLvRhvU2ki4U+a60vZHnQLU5xGhCs5ZTGnyR+6yEr5O5wz+0Uh5
WvDXZkTaHwOttA/Nl9s+t7UZBMygBk1T5XguFacbbmvdpy9P2XXC/t8lBbQp
INh3WuUiZBEt0X1oiP48Av+GhTQ0akIfxwiHmlbNmAOfgT72BpehayTsB3Ml
hl/B97pvHKmdsiCPvMoJNLj7HUIpSq6FTNRQ4dKmyC+5u6n5g4iHrpnnmWi/
cKcsttaHKdvDNuGjeMJti1iSkg0NuOWrOcvWLeBq3o0UafgYZ0WuyK95coy+
DZIRVZ47iwd2+vUOv4EbBsJgRbN1vxzDC/eGkERpmIZvBqZ0Nc4xcfiPqG4j
xlF6wI4hAtX2yGD10QrKHGltJOy7KcbdzQsl61VD49O8f0HNCjqS14OsGP3Z
ZueXnyiAnoIAmtRd/QOqkOtJ4FYkhFSEwifyEXtC1z8lLYLQjmUwS4xcq1Q1
ogfBLo6PukKuuQ1kCW7+5auySA52S5muD0dTck7u+NRCHjh4G2Y9vcTxmwcU
3e1VCw7Pwq5ddtL+AG8vhAwtLanAooGC0IkJcQN0fBA4UCy0aavTXrHEQZBl
XaqHYWYTfdSrak1ZRrnB6lmtdgmQWprpdBmceXR18fbbm0l0czHfuOKQb7yS
SVbRScTrE8Bm4KfeqWXu3zCWaUZU3E0gjk5KjnJR2c/1r4PfcIXLo3HOWixd
mlELl8QT633MunFAHGsEw037LGn/tcnOdDxjOKKr253kLNAsdXiDivWY+VJ/
WbzHEGJdr1+w6yNQEE2f8ONzqbzJpeyPb0/p193DCDhgEN0FD+nQ7Bs7mWzx
RcvsH+uX24DS6XKY+CxEkoAZ/oqFv8pv8vU+7smk7+7NmY8sEfhPu+AyhbZ/
8Lxr2aPoVnji2o1OdJ9O84Ck0Yrd1eTTpW07autXrZVYBL/MUEwEXjLJKKy/
SAvqOyCWcCnwBEceJc8OuOUw1x+70R39JLp5gFDDX9frk8hwknKB53+sV2xv
7gRU4wkP4slmKEvVdQ0LjItR8r5zpYpm5lF2j/dfA2yufB3mKgtzxhN5scMd
JsM79kQJbd7n30d9Q3OYnZjPpO0oNFp7vJby7I0u3133WFk379Tg8UiwEHcA
7M5x17fkopNSPLzT9pfDdt2xxSaS4xChOAt4D8CV4gD31ea7Lc0TDniSCKG2
fk4U27eSXCNmzoN3MLAH1ovqY0SXC2bEoXj3/iWE4UkkxmjoFkzFWpJjfokP
3mbE2Ogn68SKDQzkxlTeB6EjhnaRtNFhxW3oOg+VkqM5ua42od5R5vRmdEqy
EArvHWUI0ehCGlX/+0cQT8l33iSNxihZB1P8+eouVNOr9/6NCjggllXdcXTc
e7loaeIXEAa2ac9/Dxt6In3hlzFGv8d18kajmyxRVAQYcdRq+I+owY6Cg5AD
5y9/0JlgGyTAVxDnNnpt4oBXUBskjDa2v2Ux4bPYzZWYN9KXKIOeN1oK87vf
MQVxJitBQ9wt8meD/Zvy1BeBliZzenZrpmhdbX00zf5jU7UdY/GxVbIBVqkf
VDnUjJiom8QflI0ffWdM4Rt16KeVJ7DE0EAgLH6LpY6FInYLZAObxPL4FHpX
nqLDBshHB5FqbbSIseG651Yib3qcHsmLwmdYGfmFTxWAfb5/t83nQVAR/cGo
Cq8Hm9N1FCSkB0+rJW/pSK81PeO7UCSAzgJoiplS0Tj+6pvDO2OTL1Y2ZSNT
H+huBQTK8yguNhw3/FVcEg+DNCnO5A85I17/4ekVzxJuOajVaOE92vKaTtz3
hlNin4Yf0AEHCGPf2jGAYL2JCvcUa0BGANGRbF/n6coj2IxOkk787NXoPh1R
FJGxFtRo46wcdil+caSrYKcthtvdAAEx4/k3LUpt9FG26tPXc2Zc6B8xdfS3
GkVp5g1RO/95gzmpVaFV3yz0NZCtSJV2+y8DHBvembi2z8JRRSn0kyYrrUXx
FpRY3k7FblvHe2D4Z/KGRlj2k6LZ5k+5MgffhBDlrhMHuSKRB1SEAjrBaBDv
2mUzeLXZSE9yE7f6/8ZZI0yNbnLeVcV2R0vWOiJfk7rwIvjhhNOD0gFv6nPC
U2tBteSAzKeQF3z4Gqi2u9saHdA6533vZdd3I9MqMgmQBkH/WFdGnKHufYaZ
VM8qhApCCBlWuWCnmqpOAriAoW36hWhjO7wROgYxc2Mi5M9ZZWFYcvE3YE4l
+8woQb3uAtRhKkSHXVlsg4qpxe2XqFQvjzceLbc+Ah8ANYzDrAY7OzCWTPwN
OcATVftCxU3cLbw+jf9cfHEaSdFAknQhCZi65rcffkODvAUyJlhylQYeo+P/
FfqE+Iiw2q4rz/kWP2ED52F9rOL9JMbX6SI6h0anBdipWf1iPr7cPiF/5wQ9
Raueiat+izDIiLKhfj8pPjR6xk/9uqT9Znz5cCX3qM55rvDoLR+4zzFlJEQs
xpt3z/AkUYEsOdxc2j8019ySh7Ppb8Hd2dM5vIAERnaLB3/X6gC6v6K4Ewbh
qRxzSRX7/q2yZvqSXCsYq4EEvqcI16fej4ufKCrYHsrwwkzlyJ1AMxvogtFS
05F7dNtiSKjzZpYQgdc9FiMBq352rwLd/lhS6ISM9+ZtCqK+gzhVPrq9mEcG
WO7kMJxja5zzPCUU+TmbOH+PIHE4YV/3xmtXGpGDG89G9yBn3EjbK6cUI5mM
VfcR9RW29yqnET2PeiWTDY1NXtsDKmN+IMENJVtI1XxDe5spr3ARyk4BQG5X
ugabdVzrWP7+7EYiqSPrhjbyvSR6VDEhS74cl5YpKrTvxOgzk9HfW12vOa+D
chpj3H/ldJC4xutOProriPmA66mk7qRhx/2aolfHg+gAaq5YL6zTD0QTtryi
JA0xywWR5kNzUN2l5lxodFKLh8hThpnEryuEJun9CxlEOhNVnKI4JNdf4xCa
XjHtJPPYF71mlyvP/ZxpRpMgQeckjtqfTrYtyzv44ZmBSV2zRBvtSsqbzxEk
ppjWW8kLyxERCZOaHSb7ljqBbZiNOcZm1E0fnnBfgryNuJuIICc/CaFtubHd
G8igGMjg1RYwko91xaOWKy8OJGlZYll2z3zbq2+Kr6cjXJNcJTNVO2yAhh69
j6EkPgvRjF+WATusO5cHYcOSQntpeT9fEnz6Z/iWsLwBpcFhXxbbS7Goyhmz
7bKVdCL8srPBuY8kThhB3hbyW8BDv8xOgVtEqpk6AF1CIh6SouBndvLoSVV2
ZU9HAi7qN1NLB43tXLkf1c+sx5rGqKVyQWngVLRUPMPJyaCKiCApmSQvxXfk
YnfR/oEYOjBzZIfIdg3A4gIZLqaDq2DcuCMqOGtcnWD5VvlCv4+9Gi9/bbX6
8SAlcfrD7iEvJk1p/7+UsELNJ0DLFcxvRgdIs5LEDJnEuK/uEzZvaxxPnJpG
x8Xv0DGKp20rWJ2OXUvM2G1Pp6lE42gUV1V3gV2NC+alBryZmxqMjU9usgh8
2XMMK1olnzPbbL9FB0dbCz5tyNBKB5Rv6Fb4xQZ5CoNm3Vv0ACQU+Y2h709H
klT0Wovqb6/VnYWjCjSBIGawDfaqIB2MzUBggkWEdBrgbmHdc7Oa68PSIReO
TRwM0Srt4/ci72fAVLn9byj1TQJ4X0B/gT4JOMeEHxZQgJSIoTJgJL3yhL4R
sq2ytPvepGPxAcAg0Y5IMdX4REG5SFjBVqgUmSd2ngxyrxccEsW3dLJTJGAr
r4dJIrRcslzG53uh0WPVQY6JeAbzUEqgRipt5l73PHdDVReH1EfpXZncOuf4
/JCw2r9sgefoDMH8d2v33cG4cBuBhoMIyjwtf3Hfgg6RHwQNAe6sreElakmo
UzDiPKdw/1NzcRBnZbJPNNCtBYz9Cd+I6UkqsJoPBJicW9eLvjqn6pnWfySQ
0XBQJvqch7ePsuRFHCvGDefys+9MqrZNWW45FrCQrLEGrFJRiYUiZt/MEvnA
WOkP+j7FygyV4fVsFBM8Hb1jV+fm0+7d7uSpaRFpLSiSA2h2gBmE8g6RClAM
p+FaB/+3IxwT5gl2w3TMtx2rVDOt/HlaZwmqpUxPZY4C5vhPr9yh8wn1dAhc
nfMdB4nwdMZc4sREiGOZr/ebZU4PENWsudbmTjQUtqiKDf8wphC05hYcSqfv
kTybxQLhzRJ96UL8wmS1xY7JhwVDOpv6vcAwjIZZ65weJ6LkkiXClbV0Ezx/
rNNjHWf5tD2Yn6umA87terdGXefSwsAovufPhbCvpBzCaAmXkQX1ZWwZxuo1
x17hoS6S7/E6Uo+c1WiEAmPArloZFfsXQC4RLvE7nVou7GK1sp74BbU/OEmH
53/JeeQVyY+aGybU7z7t0PX8Yi0zZr9eiQYVmSODULSflgKCRDHQSV2rA5fg
P0DBASrtkv0vFNghsZreCYVgWc5s7q4SAU3oq0oilMrgI2Q/gmrcsdh3IbNh
EqYoqGHLHovB45Q807Zn6VU9OTVZSNb2dyR/q/Atu4w2GdxatJRDrMav0WHD
/R/Vk5IaV6U/QPU6EBeGEV3+DgEYNlNUC5WjntW+0dG/izvID4gVbwLEUQfS
V2pBPrFowsVg6SUrPJ3EbYXpbKk0/JBezBKuzWGAkDVM0+xkynjB4pG7cU2h
GkiSSh3jCV3UuNhwJzXowfIzW7mstXM6IrM5sskpKvGD52E99vDSE3wVIYOv
IczpL+iIvXDzna28JS/WTmoNk9wE1UPVbr09imhwhSUGHQdKqnIfW1Ft8Q/m
KY094/evq2enaakNXjgyoGigX4sX8uI76716lQWbAhKBazrXYgUHcadKk3Je
ABo1OI6FW4E+q8pPCFrTdsXQC329XKgOfqvi/lfObAlFGmSTJbFNj6VD7fek
84qb2TQiELNvTSMvuidJ8ocQT0wQXWZef/M1pPhFlqoULq0WAaBQPb5KZAiV
jLiebUHJgSYM5TnuWLPko7EACfOQFcv4Ne7Xyt225WAIPqugAtWUd2VHIhkg
FiKY+7wVUUjf8g73IRw0NujdXzucnYP9EznY2uDo7sN8W2wHUICEYvnZb7Mc
NlWD/QijoPyb9JT2NCdGhJP9AavR2vR0SmmCO1B2hf2+lfo/JT5QdMZncHXu
dK4tpZYH2M/6d3X5hsBoyjqCmNUbiKq3+p++z/a1YEDf9xfmL0tEr3NXChUy
f5/D3b39SB0lPhuAUFyB1/iealCAnE0UOxCuNyD1l2eEsyGubFVQDfmdKTXK
0QdRor66XGQzVdXoNz0orP+MRb8bzLdYTlW0UMgmXuB57qTUeW20g2Ikh9aj
unOQSnBRUuDSGQyeTOt3qyBSNVFLFYJU+cJ0Ttq3/rcRCjMf4BB1Z7w/rAtT
D1mtreM8mjbIQxSiXVRkpvRZ2LX2dUsbEv7ebHZK6R2oAAhY3BJWxFNNd8in
5DZxUw0KYeEoL+65fgUfWh1HlENhd2BOztCsKThM6GeI9b37vHvIkVo6fp0a
vHNREgJtBugmZtuTANhuQEC8YCGGomYPwRHSlT0m1M58evdUTb+xBN4DhIT3
wPQh9zAbblaPA+9DhjK7P2WENq1TVLBNtXIupt6WLLyQQhVyEud2xIkNCMIS
3LS+4vmR0h0VEO4J0oUl+h5sjbMqeGk/BgSgXIAXk7q0GxmrGrXdifnA134d
zyeb64rywmnII9ik2xqF+TZ0rZFltT52UGu5tp9+V+rH/7u6Af5gDIwyv1Hh
VLkRmyQiPqY3JFueILQpvbHaDW6wGy104ErhFGliDTjAgCK2+m4wHgwMzGTN
QcCFKimXDZWeXw46NjfwS/V/OiYulxNsUfh2y+kG0pYMU4/WUhflpgzbwSHa
olcU+ek0K8CYy0i9oeHGWyoewN7LWR/BmaEoLkBntaBSibyqHI7IFpn+27AS
WSJhYfsZj6ktB6m8Nxi4Iw/MApmGC42G8yz8jEi4bgg4UQUuVkv5rH6KJ9Y7
BXFkiGaYYTHcLOGpo1xSVy068beUpjrGvgWN09eXGJOr94VwzJDkB3b24VoU
6guC5p+QUSLjU+sIKBc8G0jQTGQs/CAPzENO0uQmgjz7efuXgfppP4qXDOx4
X5OaTC4DPg9NY95Webbk9GAQDBNzt38idtbO/PSk8QZ7zn+G842uk1CCYRs4
uu+inlUr7xXewrfeKRAJfTaU0ePKepkNs/nofQrTLHktmiyoegTw4YlmWp+y
4qietQaQl9N7cG47/Z6cxNqFbbtrvaHBi8sq5Ed2NTwu+QlH4/3GN6DQJdOQ
3CulKgJ2Gi5mxkhKVG/TN3hLo4vBZ7/u/3jfH7OGqfBKKl0csQGlC80iHamE
mdtpDn8ca58svPr3OxDOtUDCWOI5K16gJ7g4TmBr79gTQmAq+GiGnikg8kCX
N7/j+tvZIxivg1V9f+PVqU6KDzn2PjbYswqHmsgtktrM/1kNKLUpi1Roc1Gy
0XSzOn/6nVXrZK0yY8VGZnHORGULlaKSjamjOZG+W9zg3svSmk+45V1T5xtX
5FabrtP02RPVY/842nGE3fEngoUGXPSWekADO3ea2oK2iFhjFwE8Ee7r2WXG
JFcxTd+SxLklgFuThlZuhVK3dq2xxA7uMcMBpxsITDIWmQDFuoWh8V8xuidp
oHkQLxvIZ2WEAwmVX0UtPgyypiHhMR+A1HDq8Vq/3C6dEWBQXxqLbRA7NhQa
yOXiupEKnLo722lEoHIGhzp+g237Ip8vik6cMqVXJfEp3p2WqAxsE9Flawvo
z0JTlrT2fPXg+he1HRcCLXWkIYZUK8Sv7zhRdir+JcyihilNBHWLfjEOiVSh
1aTYE9pUgKWZAcsUITLnMy+N70zoFmHzn0jdkVf3sCJjM6fcStpXSqXE/g09
v9mLJg0h23BY0+QDFHIn38MiLOZoBzfRdKwDnnbnCB2u9fEyfiZEKoCBcE9p
/4CAQqInVSD7uPAwugLUiQfjtQeGFAhrsDbguvxP6thUFlz4tnPKxyiy1LCR
1mivJnxKOPW2/Qo7/CceuywtuK2+FMAyuw4cSUjQZn5abp1q0QPSLVW7USy1
KD/78MV0sUbVTUyuPG6tR7gf65AfAhwBTfCWuQjefcHsTs41MJ233Aj4QzJY
r8op590c39pNitXrpuH8uBq7P4FO2YhlkDp0BO8cwbF4ajbrt7+jY6ezWeR5
BCxh+VRoZU+Kg59zDOlvIXOByQF6EOpCg506DAUUxqQJrkODP7s/XMfg9LV5
YdOevZZenQI7m2PPc+v2xGiAm7kBbGDf9y2ixHkvuFufYf9uxIMH5TeYAP+r
fXJaVJnaarbxfXTNQHyh2KLqc2l9yQLCQUWb9kHFMh0PuMWfVO3ADHYiYyEI
y/JG26X+hLNoeyYJOjrQVe64ansqDk9zzRVSmTaihe/KGjK0rkM17tzviRNy
emSRUBvLnsETAIAuQiY5fF891LC6AecERny/YDwpfFBsMeYKfvDYAWKWuyxe
LtpwM9jSoFgP/IIphssudf1Qzn02EuQm3W1MqgN/KDM8nfvDXXG+zPJZ+Em7
RNToo2tWi+XPLpQGomm5+uB/RbXXO8+C+XLx4DftuHt3XhjOMRtGUApuaiVx
chNFyapOoeu4a3G/la755VwoPxn4LkrpiBA9gx3unhezqweKIg/GuF7UVgXU
YoXMfHS/2lhASZsllVt1qUjq5tyxt/yJ6943gOUE+iFOiAHBVJja/j7umhSH
w9xXVHTcs81nyd7MjCebUEwGFNK2WGmG5KOc/UMmYZ8Wmgr/3ZW3F9vOSOYh
5kvYvCr0bx8dxDDRtr8CpKkDeVIklZIv0K+IwUyk0bOlSTFf1g6lvNnC6Qzy
L4kytLrbIj/MB57DAC/IUugNk/gU0GvWF2B0HJdbDYj5CGV+JhezMqI74ssc
rYlsQuGyAUvF2iNqtMiVWm1VNmkujdFJt8z4Y+QNN+sfG+lUsrOKqXiskIFw
M6x3ePYjJlIpvBwc7w8rSwq1OVEHn5l7kE4Ra2XZzfDwWZ1lP3A1Q1taQ+qe
2hD6EeIy8xwvICXwX+ZEbXR0swBv/qFSFAzGpwR9KEVhZoBnoQmcq8dzmnbc
tPj789s1FIdLtw5aItZ0ocUOZjz49wXL0l+mng2jap/+jnBwRTxRljaZ9aMK
n5F9uaufHXlraaHhWynNh36Yp7lHt4RseO9UxTLeLOphVg43lPjsk6jXlZh4
JV644CjJK8OM/wLcZxb6CCi7x6KlqdU3Qya0x9qNCbA624NqAK40aj58nfc3
VHPwC20Nol7dxNOzjDz6BYmUaeEMbjkHhAf3aDI+xQZNlfZPxO7qeBbl9/CY
XfDUxO6tRONyljJO3rKYmSAk2t58IroaqB8xMES5lvOsjz4cj//eCQ9lH1j/
DImsar5sU5sG3oig0ixG1Mr9usj8CTTrhBHRhfqfs/MJRGOZtRW+CH5nXhib
wMEA8qwQJP2FJjY/07qv6NOYtz7bGHLBjTNTAX0Q8Plit1kPj9PMbrhVP41I
m6l/uUzuWkgcZ1Ifc38Ct9PiOCc05ig6P02gMTny0IP2xSAgsWU+4L7Ofn1h
Fzh05LDaK1vWbeQDTFNNhFJQdNU9AIEp/BdRPI405PssFX2NxOI1t/2ygBPY
MbqWMXmqWnY0l0fGLrMJuMp3uqm707360swdR5X+5EFP4+iboCYRUm4dg4HT
HkpeWdtn2kU08Q1A/z/3q4R3nYTwPzhe5Iu6vOM6Fle1hl9X9XKt9KEVz9Dh
3h4OzIiRUFMoAASjq+N7i8jQoMGdPwsjSiZ4DgBV4GAy04d950iHyrBeCSU2
JfB5bc+pe6FGZ7ynRO78afB8f1bYSmHy10fLtS30L/sEhYQ609xxAbmpMJhz
YKiU1XZIqKhy95CHd5cnCRKhfMMa+UZawhKKsh7w90FghY5MeYk/e1Pq8UMn
RR1VY2aeLdQWEanNi1boJB+n3fbaM2KImTKfrr8TjWpbt86hLPmBlk+NTk8n
C3S5bD3kB33CCGJhgxVt6huBM9XzQZNlNSrZzUFqT57Unez5msnKM+9lLG3a
jCzEclq/3QgwAoVWCBE7XTZE7LXtuHzvWUX/WS+xCIqkzey+vQ64bFiki8NU
OBl/sWE8b2hNVRr/Sgl/nzS1btoNlKLNWEErZrqDJCA5dhH8ro6pZWCEw1O/
pl4PDnaVuILkTaNMmflYE3jzbqFeALbZwsfUPLSd1m4BGC/xgD8PgTuyv0+Y
dP2BDvwmA2gFAvk9QwPW/JvwQePm3HKm1cd5DD0wzfaPLogRrms3ifRbeUcl
DmxQHlt9Kqj/SX2Gvng7MP/D1TC9MfSNH08buO+z7WcVgA3HQ2i+uK2LFmty
cnH4ycO+1ZpaTmzE7pl/Pyriwfuk1qYXCW+syvh/VNy8Tlrzodl4yHvVp79h
jcE5RcoG4e81U5oyeskCstOnHWc39t0ned6YvBbzAejR5jP4Zm8ah8HnKU2L
Kpc/2AepY/mdhsnQSmmL4vYbQpw30QhbwX92L3b8Ww6SJs2lftmjouZu4Chn
5bQcm5oE+q3MDqlOVRe025hmWqg21BMiUj61Gid3euJ9JO4IHdDQh4eJmXkM
wQo8YMugBH+hF1RJwXidpwqt1QV6mzPsc4oixXa/eDlVuDSZdIbfoUGiaXrD
qZI/NMR34z9q8DrsbNpduO2g5cf6Gy3rAZkRkBlcvXwE35Uemy7NgcMYWAdu
2RbccBNHOxrZ0Qn7gJYTLlMP+05ZP7RBJ+pTk71xOByIm2S02p7hCZx3KGXc
51wV6AXioyUgR8aGJBbc1vyEfTlp62MfPYDXf76KhClhwdLKjjO6gVPoBbU4
cp4+LzwUcZPilSekgbzeAHED11y3JZ02L9MJ+9GlZVbyyr3MEF2yKMhroTH8
WfCKRLUrLgKRYTvAa141NUvy4+PvU4l+91R8lPZNTE9RSOjTk37iDisRKCZQ
odn9AqB/kINfCZF5qQO66XlI5hUJrzfYdsqXVFeVEjfJ3fNtTBMKHHxsZGhP
Po/N+e+mPWBy9w/cTms8MrEn0NAQF8F793CipEuA9qKAaPFWL9cj2NTpzMGF
wA52No6X/3Wu4iILx7s/bZffmzkf/9Uh09gSo/NpQsDOPU7p1k3f7PIaBH9K
KDflu0WSQCWA0KOr65LyQtxzz6lbPvrPmZ/tW+5nkkF80kZxqeyJgV1JWOlp
M9bAjrDPH1KsB6XoGQ2J4N/UxLIKwj99W6U7b27ZUKyYBc7a1wMjuSpxWl6g
iJCnjdjadRaONmdj3mHEuaoySynvfEfg2Uka90c8GU6g1H3E0fk6659LflGx
MeFKHfi+NZOKxSTfdgPSCUQUDWk0gCSBJ3SnFk50kH42jCCf6l7ze5BtoXzZ
Up5SYxUVlqXmddvZmg/bUYuNXauG+2WRQrPH6R6BuJQIITl77AziU0hCKwlf
q2badqVHUx+DBydCmczuQ5v67m+L9Vv3SDfPrYSVVJlEgCK+27pK5EMURxBF
BFF4/8sSuNm+1R1kEX5HlsGaP9QmMVh1G4C9N9VPK2J35j3Ji1CCBXLnFjjT
OeDnPS5b9qEwGXmj2v9xpm0WsWEBX+tfWMuWhtHQUMrmFFhxrejkSf8UPWT4
tpX6gVSWtmtwKKHPxgHGEIDwoWddBLzPUU+NBSJxQl6Z48+wDm66BPaMqMDS
NM1bJ/QwmkkYvcYVuAIpBo56B5r7+KJZJTQ7zF9/+QTFvxZK3QGm3d4hmTt+
TrwYnz+DKWipLmdhsob3NS3foRsh3kJq9IvnU64pm/vPebwH8t9GydzQKMRZ
A3WUCDg1vkMp/CgCuo6BtpUj9csmuwaBrjrwtHXuLDY+I2rl2iGoreBSLs2h
A1NfDDehvcQ4/R9uqavrUzCf1FAAnddgfx6iyaP88og3vQ4Dz6WFm2QU28Kq
HwcX2w9OLLWbD4RdiBJpTuU3sZRFGwa30PEmFVt0jGwV60UaWB5iQbxWL0fL
ZD6UIwboyz/ZQGNNuA+nNrVWuaGVe/yHcQU1K1Aat+ICvmggeI174ChX2G0w
lmidy4EVkA9n+Cy8qDXcuFoI/2Cx6ivrrCg+T2Jujn5JvGMj07pAlFHF0C5f
PyKqtaVwNWPJH/uCLER4Y4+7Wsotc5STfHvq67XC1moBQvroOfdH9AznUaW9
n+aZ7QSmtjOe4nfGEg9jQEZdC8sxXkJaSRmaftvnBevIh+7RWKSfLvVcloM+
/nDIW1R8z+JTaYUmILhHCg1XNlIOUyN3B9/erseavnKkkWds8Jw14ptXNwly
vTC9HNaaOZr+UMNKTJrwRq90iOybbBg06ftn3QyCdlHDbRhkLFLy8wHuGlvI
l7zeRJAF1VFhJipubSW5f8gK8JE//nulqnE0bEpzbytf1Ge11fn/PksDcwxK
p4yYaOHYCoyYW7GIFl9A/CS4979x5bmw142Tty17lhlvjKJnDIy5UCxPoz4u
+9vcnBCwoqS4tliY3Hh3kc4Ih7kpPSDzTu85I5B4scMlM+W8d8dWsch5jAiX
jEEZjClOQnhVkNDZyb3QbMVHxGcIelyAG8aIuR0y0ad3ruQO2+eM+CxbkvYm
2jGjovsSOD2KKNkLrxh3q+FhvVyS7g9wMbPwTN/YHBx6kpskE5zRQOx0Jn3D
zNmdOVLA7pvuAlTK/N08CANzUkWjHgcwjqEDZiXxVlbSnqqzl2fqIrBj/pLC
42s41Asd1BrP/UUKpPXAu82hai+pVOsQ6pzxgC6WC/y7E4E8V4NxCpAgB4kk
tM60gvgefYngRNQUMj7NNs6ygp8TAG2bvkL1ApgAD6TYYG/DkHSLTv8U0PkP
4f8c1XyrIMu7XUBYhTJAG16+AllcNXE+Y/7+0Fkz59Tz1gJP7ti6m7CvPave
0Hfa8GJ3dNRbcCif01JaSj9czXm/UM5Pv4YzQ4h25R1VyetKqtOD8/L3QNqz
I9YA6TK923BHp85rixBmFbXMcLTJ8QWip075nDn017qUkr5ZQyYefARDIHeL
xtXTboRM6e37NP4NQ9G8Yke9rziEWMJF3gB7NBuuFu39ujWFrqBz/5RYcaDB
Jhtv11VbeIDiYxaHEiXRUPWMlXzgZdl9Fcoc+yycJlDkyif93++fIbHmv8nE
GliHhQsYmRP1p+IJx0PBVzaa/iqs7n4yqwt//iEAMvUzb/youz9QIC7tQZDo
/jWJyUV7KEfZ8yl2fZj0jKxXUV3ftAyYwAP9usfv1BxMqtn4tFLY96arYBzF
sRrqZrS4QhBQoLSEy4+YW+ZGluYltJg6nJh1cgBHlA/Hi2Zkb1fRaEQoiI7/
srQSeGIZCdGF76aPqqYNFV2kMnBZITKHVjLDBrGIQrNdAqzw3ctCwhr+SLTR
anhBK7naqJkTu/vKNyUK9s3qTPTALMiiT0+ng7KRs9+dUjBij/2D6DEdqmOx
xPzuUkoWZAraMXdRTv8QMR8uHRoqOHBQMsT9jqVJvO1LuTkJ1HDMAywbCXTQ
fU1l59Nrljb/socY5TN5r+qFW616Lp5CpLQabszLWBtyxeQrZW7h2lNYC7tX
RLhTlETl1dDmAeJBlv5Voq4XmoXWx2eriyh0508UGcF8jeL9Hj/M4d4ZkRml
7YuRoXfDXbzQ+eoweb1beRFr3/C4qYxMDDqnUEL31N9fUC5VfSDSmWit/Zna
dor2NFEKZAlp8sBEyqMpLotSB9sozdGu4YAuuBAFj9Mz8Ueh85+CEkgLGjlw
HhDKxDJohScm7MZpnJoVtmU/w3sHI/rzLf4Lw5e8UK75npTvBEbTiHBqXHhG
bQ56pk5Ww1lvp6hmo1pdGaHYopN9pwk1nXYHmC/auRHZ6RHaMH7uH562H33s
TXxXysd8mjgkM43GRoHqbfJY6qcQm7wyi1pIiSlH0UjgAY+DLwPwxUO8PO76
gaHnhwFNWSZtiur0Q0c7uQwl5n41Q/8+4LhyiFzX+A0ODt8Qv1p5iFAPuHCf
SOyyGveeUqlxasd+0A1UyaZP5yT3Y7eJaAVedH5WNk5G+adJFKRqljdHloV9
lbSj+Mzt0kw8U6PEpdq9vH1XRWJF/6eUmE7ZUJCG7ze9Nix2GU2UK8arNtwI
+2rg/dh+EeLg1SbRP7ihCXkolnrU7JnEC/nr+jHWCX6I8IBk0cXinlNmnYsT
YjF1JCleP39XP1np4e9r+r+Cv1roiRtQJaoJ0q/B2GUC5c/O0F0bkQpos0gn
a02J3i1Ohdit37EeXUlHJi/DL48a/qDDAwceMRtBpz/qy/HzhvPKerUBzj50
qua7H2cKeblaFfC5MiRZKgs5yZlM0FF8aEXIdtNPfitOjjebIXgpecBbss6/
GrP1nV3ZTTpG8UsOVcS4ZzVMS3KQBGD2wsyXOGta0UDUsaeF0CCAF5/pyaPg
VfNB7j7ilGbKYpzp/9IMe2JNcPCzWA0wTM7LYgYGzcZ8GeGzGMrMFxb/sJXB
SVzXQSjh0E9gaBtsYv8c2BpKSRNXBJUbdObjtHCEksaGE//FzoZWrusaFcUr
Syg/BP90Wu7I74BRDEG77e81g/qEaemoGdBmEZEqHHoYImGPtYC7h4zjVKTL
9rFKXepYAsyzNxrfSDnV5regqWggLFjvRfDS0lkAhPG8nyV314CO54WOPrpk
WlmBonLE7MR432pGGkT76rQ2gCFugFnggKNnQtwPmdSd+HEvr1KVVDgu+mfL
Z0fOGjCYEAywLT3pU5Yi3F0SztVZmcFJaRpaHRmPkpP+4VJXSJvGZNsX3ter
3AWYxxxp3f+ZgXshUJwIJQKnB1DoQ92G+MOgpWyZm2smqHT4UTVmgcQBNMe6
M2qxNVOUgtoEtdxV39kOxAB4Aa0eOO64mWc4FRmrjO9Yl0RCAGfVMTALvdMc
TDYpq8dodqqSXK48tLl2UWA4rGisdVWGvw5pB9MMhLw6UOrixYW1n5Hr/og5
NC+TFY47AhLGJaYzxmlxpl2CI8WndNtJqxhcVRHX6Wbochii17duT84rzlGh
we1SKBXQpXA4ijRj6dk+T1KShvIKbQDTNKYulQbJU1gkfSqCJ4+HGOhMHDcU
oA1H/gRdMsnlsb+0sbzb7YkHfpBP/jgtarUOfOwvHGVvpavaevCsJL7dbkS1
MiN61IXXQ2vCG+9t88mJ1YeE/tHpI/BptFeqfBTddLfsxCPvfN1fhRIsi96J
cOGR6Gk2HOkjpc50Dx+pAWVhZ98yjBiRB2/L7MwvNAJbQhExmJaNTZ2rCqV4
fsJYSWEUYIh5jy6gDa1lmNrO+kCLor6txWjs2r0JyjOQonvUdytS+efr/+qr
OcDqZnZsyjFovybECV8VY/AXe1UIODtfPf2JUTTjZUJgzfzrS7Ax0Y1vOxDa
UOqTgPax1GeMj7oMziDLblWhNivBu9pTuXltyX62aIcPb5N/iYniBqjTQ/LN
QrZPh0pKh3XTdAgMf5ayhCVc9j3CZraKDcDUpqLpg8Eov5H16HvZE/OOk9NY
KV3qvhNUHamPguKnFgeB7t0mdlBcDbxEGyA1oYconlq5VYJDvA3dPbO14HOM
cyey07ELML4JiBpoSGA2P7lb3h8JrO5mEHbyM+mcDoCvoVMk8U8FZAm/o+aD
llBCgEkdmZgI0s5/2XONp6EV1NXacz+2xawKkVJ5H+aKf3dcCJ3U2tkqRkm9
zXcz4uAvIpfevAadbc5iy8YzrJeHV0tGvAIq85cgaiQwL8UkYD03G8oJAEek
JO6GyPO/cQok5rZjm32vk5AawVZLclfcdJQO6qwHUaCEXqIN/zTpRUNwRawT
4jbFUSqU+m1Bw49KfhB9ZxwVQfRJd/45AOTL32+THkxTYpYR512Jf6xKL4pz
edPEo1oljoQj6bCGjnY+qIklEuQLFp9NcSB5LO3O+s4n2sP+Y7LGnb1+nhFO
swmi4FW3pTXetCzBlBSKyIJJQpuUEkqxsCHfWnVRXQQEe9RpE0TEPIh3fM51
empvH9MGWUSUGlqXWBxPpBXL+MJ/g29e3d2xjSOoa7rBnEr1ash5nnZpEy74
3orP0QaMWRQZLa+NvhkFIbnHeWsnA7cn1fNQEsC8oD+lkFLf0jdJOvgku+xK
Wiygzfi5+bgviv6XkZK5LFrxzp48HkLL//E7Jap5P8xInHZ0LMqpA8cmj2YW
inTo7cW92CYeQOEeDjB5uRqKaImHMBUQntNMKSgKTFW+erMPRQ5uktD/gZCZ
sIfhTseUwQKYSVWr5sVe2mo26Qi8Q1ypTAo7OPWbu9lgWATFN2BLy/Ex9hTe
NKrr5kmbZjc0F7FF4e2xB82WOw92brNl0G9jXpOQJZ2BO/AU9rvvtxWBLNXT
00D/B0K7fo2FVxvy1pr8M16d2gsWToCWWUtCnHfxmP7jvyp/bDr90Z11r2s7
Pc4nik0WwxaSXttIOwV/MQwQ2Q6ERH3gvvuAmx9TOJI2C6LMjFQJrSocPSZl
huuWtwxgAE+dBhX/68PH8cZdSkkOGqbTC9niv3EEOmVwZQBksNA3H90dVzPh
amcPzG1bQ7PPt6Soe1TI6KtgoYtUT0Q1R2r9amDIb21zFWy9i6L9SZROVSPm
w+mgFL0Z7AK4ixp8na2HsybxXb1YWTkhl5XU9VQOHriNUD0J5fnTaPE5zU/p
nmTu3Dvy/aHH4y+ZfSX5jWtkIlc0XIzTc9FYhoivH3zYKUNqIyqxnrxsoEZO
9BqImGHLVJ/RI/7nOeG+9r2gelNQCN5TBSx0+ILckj/UtV6WWBXwktYv47px
PHTdc/bIhEer9N61iXqIAovXpCtPKAFbFoLRra7ePY8p3Khmci6NRoRyizip
utUZQpVi9vkzo7TQ71tEb+l3W4FCZdO/VAt9t3/orvSWB0SBFRgxLpDSWJIk
C4hRhHC8ldylVVrE/7kVIRwn4ru7EEsHaTldtnQ7TNALTnIZsVM5X6wst7iO
z+jPV9bDLvhRVTrQ3/crRRpDLZvqnZipspMhYN40cLovXlnHmU4I1/3t+IbT
HY4fg5WClYs8Cegxp4rtT4Oka6DfWQuU0647ONFZvgT1vnn2VLOqLg5BK5Ut
vEa8b7lg/6iaWDKXL54YwxNzDRVbKTuFt1iPuKuBI0l/QvWR1a8oAy69jvrA
SJ5rzBGVOXmsbgzzfnZXpukApmFg4WUT+zwu0QGiOFYVGA5uz26yHgitBtQK
fzzmTg37Yc9s8ZP32+faDR1lBkfS9YhDRQSbiicZeT74JlNP0lZO03JcxGdN
ZANpqVD8mVZNe19koHInCpAgCgdQ0YmAJPpS82ldw0k9gW2rO6HUyON6Oq6G
zsuFJvvbZsPv9nea8lidHbZhBQHwl2UOW6CdpS3yPPnsBk02vFpANOS1J7XW
Cr6U0/L/reecUdDKfV6UuvJT+WPyjKHHZQCVEQUhAn0ThFztq+Zm+9bxlNqs
ElAg/MRTpiqT3HHiBeTG8jNoKvXp81n4q1MJEfT/28ftGKnFo73J7E3+784I
/5hMfDLaxxPV2+kcTNJ+MGwzEIl+z0yopo7APfHWid9P9SFWTRrNmUpLg6lx
8qkV5Lz7w+qISSCotnp49NWoPY/n1N76iPamPxaqIUNnx42aEJ2NhQWepKl6
G5xkauRVsu4nFiH6o1pyfElS2DvlCpJcNErVyC5TQXgCCIuoHn+f/8WtLrh4
B5Oay96fT+2UeWV5BwJdEgad2gD4R9R1o3DxAdk6htkdcE0x/VKwrGoYiQ1z
zSYk0TXD5hw+3v/Y2lCjYahkEelJsfs3+2az1YYQF9Qr/o7SYg9mQg9G38VV
7UJvLIPTgs+ddGMMhWlqtfG4vIJG4LMH0v/9n0O3TAJv9RqFPhWthnM9uXyJ
OgxCObmPCTGIjRqGTeAn2YRcBWOnbTrhC+GJovWWV8kQn0Ebj0TNNNRwxUpf
dm7qbV9JwJ2v4gdp5JsxUUFZAEi/HZD2LDUvY5eM6gMwJPGgXFmZ0c6Bij7E
sjp49UI9LjsTW4DCL59aiuumWUyxX0DPh0b1Cseg7dOV1/33bGfm/oyRBfMp
FZ9NuVzezdQJcDBrCKvSoOrBvl8oF2GzLhSbbn2oQjaJBEjmRLi1QsjoAduR
5JUJ1VJn7Gj1/itAWhUy8GSu3qwB9YNXbpJGAONrM4hju6wxzpYJSrW1NXo/
5zzmA+JRCktGZ+USsxU9m5EsDYI1ppaQnyplJ8NmL/3+oDqKHxPP3yTI4k+8
QFQztQ2b8KfpEqcMUZH3nvpculcDHylWRQhl+nkNU/4PuB+6I1SWoop/F9qF
EWS6vjA1CDwenzR3nTxCoTse99iXw/dXKMinIb1SklEdzQUGiGmP02UjwHFA
cNjPUuH/7cRgt50D9rxc5KzfM0OWS9LTAck+4C5P6wsHNc4XCj577/cZ6fCd
apd15FskLBS8KkQ01yQw34QcbK2IoU34BfK4hcfdybwnqUv/5ZKuWor9cyNr
kut+g2nxSOd3w7rkREM0L30/9pVNQglGt8XgAqdGIhp+Q8vBzaGHFLG3qDWf
uGnzVqw2/RTWWht4N07LdsiPRyh2iD1znPti7eQAtbUVu77mlhiQyJILiVV0
hlPDeIpTjtstPrU8TqE1+MIHoPjIWBAxmtpBHGT/FcipUhfYRe8nEbCeY6J2
HZQS1uVjPhZnQywGX6k2vdTV3KgC5xYL8ADvqDkr4bEMa2lNmn1Bmd9somFE
8UVsGKKY5Km+voNHU7qyjx2hTptmDQDeucAM1SrvASY9H4moMbgtvl0PXTjl
0jQq4iGJ2iAvzX1uOYrWX+7MCDBT8h9UjU/pkJxqsc3MwPQ9FlYsbjsRxqTu
XAlkumnhTxhiaXlLMDT5TGJp/G4jcb8Q10w7yp+4gFRX8I7ptUJA31T+EFZJ
EcXpB3IPy55YoFLLNDrnqubkn5JqY8ZxW9n19Wx389zq4myLSORroiraf3kc
7y68ulLj6iWdoD+cbUsvSvnGAOgmYXboV76svwuQFtyVmXDUQr65OKwPZnCA
7adoVxSOEgHcIPAzqEjlZMP5ZtJ7U7i4QfOaFm4FRFJbX00nDG2CjBdypK/W
X6Kgx2zqXv1wA0FTmdk7+7zaEljCEWpD9rLwO+2o7yL+JwDAphQgj97rBCLc
W0+pYQs5mxDqIMCrcs+g/TyNdpIsHKUFSkWkiklWOOWc5HlT76FGIon+0ZfR
q/1KvcDGA6HAk472161TPQ8YUYoc6Dl0O4jnherSIg9EXS2wgYK+7m5VcNNc
HXMFmZaNFMvwvrGIxPr0T+vnKo9vP86Qkl2RAzHtP9AUwmDyzNMbaUqKCXJW
KFfQE1GEaf3KuoWUke6qHbV9v8XVfx3+dcRsnbxVXEYuWkpzYb1PACyS95Pk
+Rbi9DAdr8zSlpUdpn4MeKqf7XzcqeFElvIwqEUMpV0/ShPMX5+5Avjln/8q
8IDWjHltUpURBbWi5LLvH1gaAWkE3Z6a1am8BXqHUyCt7kkxXxF3WW5woFf0
cUsOeRl1JZVOOR0VyQfOeo46fUmw8u0nGLmXT2S+/WR6uNInpm2bb3DaRif7
yzDXoK44S6KrywUu5CucMJVt+wpwSH13bL1oo3+zo9vzU0+vZIMJtV/jtgPq
QJLoZaO5+/4039bzyEBSXPCBwTUTHHLZbPj3v3/jGkcbrXOdvpL9bkwHKECg
vPwS+lqKh9XT1XtpkKOYJNH+Qbk30yVOFSAlFq1A0PN7+LDhter0PaM9e6Kn
QDHvDPhX6d1tVGh/s0aSIZTzPP03Iv685qzg7whtGPz8Tir98d66HFbajrdQ
i/yXzaD9rFHr+mog/Ik1nxW5j0b7mpiFIVsPHw/1juzK/GR8/lPt0BQmI24x
x02kAYm52/FhNGQQowh+oaDvRjR8esJ6DFWp5hVzSo1CJ6BmWg64YJyvNEda
J1bX8JQXWO8/gD3uRb4PZk6blmQ4Nekt5j135yt0D1JANFwdN+9MOoyzApt8
+eKjophKH1wsQUC3Orko95RyqSlmsoldcQi1ifCdDHNK2M1zExuMMrAyUdKe
w3by4CbPnUY9VcIu6M4cJ3X/yfCRgyBLaGBFiKu+NvuwD7H9Dag9f8OXPiHG
ODxQt5GGNWB3LoaCiS8cWZarVSPjNJerwDXU6xssO2o88q9JqV7Ej6Itcgh9
234P/lD8QGjVsVU3bDWspGmc/GTXvNwu0sSE3nOpL38p2qxph9QxvK6foRYf
R8wwwq9Vz87qPlHAFtIkLHeeWHoAQhhX8kbIGFqvK/rUlLP8CaGIatQ87Zrb
pvUrGxhS3Ng28fDBF+Hi8QHT6y3Wl+Kf4xdrTTBha1pjF7IqgjR3ZvFJN5sx
uSO2iopNGOWpKHMTVH81QEY8tW9ES4mnwnsEBRycr6pT4MKqZQEckUd6WloM
QXd/luXQIUilNxGfeJ62t/jUilGPmEsaGNTSqMRMMOcjkLCkXIf+Po4r7bX6
WRFzSiBi45Lu76suwVsAhKOUs/p5tIesvKd6lQ6vLkdnHRltaytjktQt75wh
4nLYxDPN+9DEunMm6MzMkZCJP8wB7W5sTcAs9T2H2p9n4Dovb3sp+j83H4LB
vxnyhByBDyFDk72JFS7Wr1F7HvzpJ6O0FZGJCR4Khl/tKKEcGcCE3xxVlAhc
L2OEX6is+9yfvUYLLKfhNQB3ZjNgVpZVligvNo6x+NXfVl31WnIeeOMCzNC+
IvQRlaY1W3JS3+wd/7VH5qGM7C98WGLLomnGS9lX2WU704zN3fgXh+KUoYHX
zii0fl7u6NsAKnuixGCXym2jTrKh2ZUApAWFRGJ5Ze9WgB1h6Pa5OWgXNdoD
6LsE0uo5kksj34cCrABygQnAORY+33L4ei0KYCdCPTt1aPg5YTPKPLvUMHN/
mEFsyS1ZaAIT3MuH9G+E3ZY5KAD6pgFj8Stpx+d4tZvajXNRLwjLR77hwzNA
kLPYXzKNotFpl+GIKU2ZudVEhewMfUbMj0kI/laef8wAwWYJ8gLj8qc/pO2a
3F3m8Y3GAHPJ8B1kPpNtr2kerlF+lOJZ5Y64XSsyRygno/tsfxIz2qMbLvgp
zhmpCJqHLqHJBDWBmahUlxVLzbgOFJ9MYve4nBGZK/9YhT4XN39GQg9QUzNo
EZJ9qs+GhUokRD/572dGiIQMGBp4I4IFjnM3w4a17z2XxZxYdWtTPFI8kCI5
zf7Hjc4O61gdQd19ciKeR7Gg9qxLJfScGodCPZHinybIdwdK9QNJNp9kR6IC
TEMNG10bqtNvaVLpXWh4DKyuk9KqYYK0fL7hmdFecPDqQJh68zQ8F0yCE9Il
c7WRb42AcN1ykLzZLmE8iynsXkA/T8GKgHMzi4dewTZnBGwqPAIfwqR/J44U
A5RiFBYXgQLybawiDt/38U66YfrOOiAbrD9nx19AHFC9p04xLzC8iQFzZsUm
Jywi1Y6lLx9+YhYReGhre/VaRcm0kDgvAvYVM4mAGhAkkih6tPs4P0oAexcF
Jto7Uu9f7rw8Oub+p+m2IobgXLnX2JKnaRsM2nGJ62qWx2W4AyCOgiXwTzfz
3w/3z+n6cCk2K1DdoHqBoQgCKRpCbI/sdDOsOZOUggVM8vwsiQP2jddAjNVm
iavsBNnlXGMO030ZuNqk15Oa2aZXPj6Sek88Skq9hLYiGEFDIe+fs54JsTxg
y2zmJqAr7QmAaFpmu8Tb0VK3Vb3SCfJGDYqZH38hORsLhpwmBv9QZ3rNLYI0
bYfjOiQ7S+AgO1cBxnc1E7ZMvBVMq5PqZs7aUCvzo+b7Jzy8AgJFjB0Kn2vq
1M/jgr2WRfo/c+jjU123rbUCEJhcwjysQJdADK6UsSGER/xCShNCkkIHsm32
7cb/BlurLFGLD1/HbkPPK7do37/WA8eW1w8c5G38oHVfedsLrGun+8vRo9Jw
wXzKvGxPVDmZJU8jBzXC8eieXc1zWA20cqXnzvyHBDRdIdwBOhgiPNNFZ4X0
zYpthaHFW4S46K6/Y4ZqC2WN8C4434Tf9H3GWtbUfpEoWqGbYN5iecmgW2Sj
HpXwTNwtdivR0H+sbhl5HSTERlD895aQG8j4ivKWFaXigZEP51D/3+ZsqJIz
5UBLLomHY9XdImMBMh7AcDTxAmyDbdJGtjaneD/o9bRo+NcqPNjPsVMftXRi
Xa2xBFCyi9Er+oHh2aAGNLnBn4QtE859Xv5kecMKlYEQYNulAF8xIPROrxUQ
UH5f2TQCyXBYK9AkdODrxZGsZorhyutc75k85z1htbKVzVDkTGafi30ohxlt
cJX3xsWQCV8ZiEz31smzx2c2ehnZR7+hAuLcuFqfMT3eV4hi/p4JLqHUev/B
i36PtK/Dr0r0QxDnE0wzHLfXuEPYUMErQj/FDogbdsbN6tC6Vuc0lcJneVHU
oDOoysEvCDeU0J7L7vZxFhgsvm3/313q3JqLM6xBlWOwZPbwpuykJqMTzljS
HbBwhvAc057JE8SHVWAYwGa1nWeHgbBTwWbmvyKLq8/hShS/uZw9+NaeFEcX
0aT1loiQysmgsn8YBFKUKvHgCBpDLuzGlze23MRgf5YfuQ2Enjwdm+zEt/jw
iIQrQlAzyAjvgkljcFwlxh8NXB+oQZtXAvpyxIZX5mdeeeTzfwbasV+Sg3ib
/EZ4tkkP4v0Rb0layIYQjAr2em3E0r/IP8y3WRTLG+QdyOqm4+k3UoNkOIdl
fbv4Pb7W+95qIX7WRrmBmTf1TWYKI99+5qTmDHqlCk9lzCMlonnZVH9MCwRX
PamzFaK/2W9dJaoB8rwsCAfQR1ND5Y5AmVIEr9MgwyiixqkwU3dRmoMZE3rX
TS7WxTxB6CzS5EKv38190ZTc3WydUKUdG/EerzANeOFEglTczZ3IeXT+GfBo
CGhUmGdObU1wPX/+GfbXj9CM4JMevXhWAvV2ViPumRHKVAWQJSZN88CU7G/h
DYsMXQJPSub4lgx+J4qU8ycXxe4KlFrmLfx1GVpYq3pt7UHKN/L3wPhGvPvf
4qMhd/On4L2DzG8TTNDr2lxtoyp3wLZWuLWExKlLxTNdV5ZXkmUWyhJWWtVs
CcXBohkN/OcUQH6Ea5nApUBvjJlkGZ4ykrw5Dq31lC+KSmGfY1UDTholruFi
4LxIfA/h7cfzSr9tFWcZLTd94qxfUHUNKjfsxhsWef1MciT85kcNq7/Japgu
Nk3A0URVDcbUvnMoZSmIyTVW9DOhrF981/QfTI1GQzuNjy2WSOi04a/QGrTe
ftvCsEIa3UO0tOovTMMuq0J9y0dn2tL3yTGTamw1hp2p9lhgL8v7v8Rmcs6e
WKse1s5W29nb5sDfOOAhj/bvYbvh2Ba6dCv8oBSh4iv03RAVUYAr8Pv2Uf/M
+kfJ9ht8JUoCQD+OFACL0lo0antkdT/p/qYwmP2WisFVW1RcDdy9IaimvM9Q
kN+H5yZDoBKy5ok88Sbx3Hna25MR353HshlKeuwZBRomnhXdj/576IcQAiRK
MjIr8e61htpoELQ38ePESwdxXo+Qk0PhM/aQ9fgO41YbIDwGeYQdiGgJSc7p
QAfLsw7BTgTu88equ33wdDT3W5ZQQ6hB96Pp5eaPP+9U5FLhK18LqLfPpqDb
kClThuBeWHGq5QgZRb1MTMD9ppBxGtfKT+0BsLo2R1WP09TkeU2ea4bb54La
JrV/OKz4LP7fKotuOcQYIJj0ptFEMZ3zSpNIyd49JGjkiUdSJRbVjjsrEtV2
u9gx5TIOHTsMdURhzx8HlA68I9lPB/HDiKrU+4/YuKFpSTnAv2gsCmFcVIxc
0YTVWt9gtfn8yESm/GaG3eB4bUWp2tuOi+4asNX2zP3zjCmqYzuZgukfgxUA
gBWMtgRYfr1hf1TS6usTvVEZGrEjkHZIM4biHdyNCKqci2LI1YdQADEVAay1
ojGQH18o2RsawxO/ICh87ZymRcZJjRxCxspRidIcWycKLeYxLbwzamMqiuDI
C6n0AVzGrDbOul8n4zH+dV0inQxHscyuQHEF9u+7qM47KhxWPKHmBN7LxFxf
tXBiXYK0IfyxQBxF7IsBJU45RoBaOe87grZ2t5gXbjnZL7biEJFx1WowVGDs
BJm7d0TCJ9kgC70uCdWDYkrR9I+VDnCeH36tjUQySjlPEq14S2pS3WG29gKn
5SdAMS+88h4gPSzS+dI4Xoc+bAruKWdwqqNPWJQGmz1lvU+aZoCgps41X++J
uJbyhiShrCuRsrdRq9bVpmD9Y9c+P89fXGcpQxJIOV3V/vY9xpoBIE3BivUU
y697SJDJ/VqXBJJ4gsJE1TmyRjysdude0hsJiQlxg2BnLMjHj2HSxqvZyOHh
r2jQ9U/i8BSD5YPYaQMpHxGVXiU/6EQdKo72Is4lAriikeysH7ehsFeFoDMn
95WHjSLUa8I2Yi763p7W4XqtO8o3jeVbrctEuJ7TYtjry8PYuxrOGPsW2RZE
M1y9lPNTOpe9fRI70kK9KiF2+5LPMpMb6Kf6trx8uI53PFUmJL6cqxXAZJrt
6ADme8qN/L182A41708otJ9TUg4NktO1/wAwetGHsDuWFyqOaJAwc04xlDCj
rpNoFax5j+jewrO1gobnFaxyguLMBh8EGV4P/A18cpFNkZ7suR/buyHmkDkS
jd/EPvWdtrpYRIvIO5nnC0cFaRTXaajrGkUt10FxmWbsJIsOTsbH7NzYeJVG
ls2VHxvOE/dMyxkJxp+/bqo0p4sDx2Kw0+zXvgL95/bVSG3AjGGEEWCyOxte
lN9KGRRjfBV48KVxIjic2x3Ugr3lWy+Kmk4tA4NrjjQdoH/XKGJymdfPj9O2
OSNcSNURuHogzpstiNZoKnWQSwdpJf1a8PloCGBD8vIdvrsd1mpvPg49rjG7
+zj/GkKE0zffPI6iIkUhEnlWBWy/JPF2BLHoxhrY9yieMLIonAyyQbamQs9o
VaPvj06NDZh9ZNgkPQSpJv7EK1wTa7JQZxI6sAATRwSPYhO5Xd4pAnBuHKXN
ijO/u3wWyTS33C8ZlSwJs5Vw5b7ecaG51zRwQMje1B5ib/w49ZqlstTBoh1b
AZlhKGeAjAAZ39gNhQJCJiWiiOQkLEDTIs+lh/iImBYqte4h/9qTO1afZVVM
d+SoqObHJg9DdYS9tZvS8zGFQ55l004jPSTrfNpiHz5pGMHdX2LlH/xp/NfD
y/FrljDbL/orKqOWmv9JeH2lyyJz5wVlMMg72N20oDNYSeu6J0N5bWGdHbUh
lAblY9JprwZX2ZBMhA+6ZQiUZ90RCKFQPxkT8lTv46Qb2VlGxeUBRQJ2svQO
8nkTN+3wLDAtXvizlRO7rzLFSbIyaWGp28t6CCPbDItHbmGbkiyRSiZSbh2H
xRAlOqJG5ZZLqxHEKy4W31z8Hb60vYV3ZgnRequqogPGPz8qzwXP9G18/Ut4
VoP02jMA0R58g7p+S/MzLC2cyn7vJj9BUAAaCgX5q703XA2FnytOsjHR+Xl0
mOdYtwxXCB+h+2areGE/eQWM4jlMy/EgkJWG7LUwtJ66t1It81nyi//YE4q2
iKFDXTy6RwW6nXZzmPcJjVjvOFl/zkMQx6fHTt/3bPY9xeJE4IHd5jolCfQk
MS4Vmacgs+LVLAW8Q6v7WItl2OHZ7fHls367sgELk1kbIzxqOmd9za1CW1ut
mfC8KsAGAuTSZ7u7+87FNoTqbVN98kaYHapMksH4Ve67SP0EtCgFsc+tYyAB
aPrR0U736aWP+hpNDAAF9cLbpSZYFgihe//x/Hham4VSJM0sUhuGw+6sHGsM
mWNcD2p2SrYPEFVXrIgJQ33nuNs7pqAgzYluEjmqTgas2MBZJHe37zgv0BbO
BD4p0osS5VBDOAX7n8kXbnEkm4zh2FAUAvnRvPw6O7Xh3kueg2LB8nUaVW5W
8xXkZoRX0h5RHzlZWoMdg3MW/Nbanla7G1GntOzOY3qAhjnaa0o6Ll2tTuCF
NdI63uWDgP/jiNtW7KPYCx+NpcuC04P9x/qePPu0xAN33eD1zcBhBbYlFLnv
gnbZ8w95zF3ezHxGhU+nQ0G5QS6wbyBkQiexhTu524owcPsTeMnWpI2ExyEy
mM0h0ThvjSA3Oh5QDW7bbA+/jYnHnpalpDdmW5LR7+JU6S+0rubanprLVpvh
glsM8Cy74/e+TCRIsRXh/46s6sCpXSE0J4kFBiwNAP1+r3F7KAmcFQw8jF5g
C24O2lVNGpYMwD26Gz1O8OiMKG+rp7V9iz+QeHVYMhyEWEnvuBZsfgBg1hSz
l7H+XyalpfYt8DD023dQRQWkpbhEv70sUu0CgzMz7nyKT+R+SVrgAOjqctdD
Pmg2HV1c/PQzBqsugWerHBmEpltL8/4oUvibh3Am8pXz5NyNZ2oJKm6DiD1w
DmErMntOqSZzTW3JdQDX7r4M/bx85gpX7pFvmNHDjL/LqbhJVyYJwtY5qrmr
7VIo77hCkn01dUKAL6OsdF2DSokvW5YhYqCtkqQjjkt8BzWgqWGAmFjWaUT7
VgBYp/EjYqr5mT5dH5DupRXUpE/8mbfBqkAy32MJ0xaGacVl6pQ264OMSLeY
AJvgNntPgFdrFWlE4A0Ct6t/Fmq9MJKO535T+jNPXEry4PglCK4NySSb3QB8
IKeunea5aKt+0oc03txYad3p4kXQa7rqdTlmY7UzdOxDdNohkK/y6isCeDQr
2zNWUxGfLQY/y9JQHm/CdGaHLjPcgMIr5ixZPmq1wuYzgYq9TQ+8CCoZvpGd
z3muuhtO+MnOwKMB7pP78tzM079EQ7CzKOoBLTg/ZjiVZXtICvWoZJuK89Ks
D6kr/bZmAqQSXPl/cGEWPF1pyylMwdC5ltl7gu4rdm4Y0eQA8pIrQ27PCVMR
vHApEnLp7WvN0vtR1Z+lgonBd66jY+Gu0k+AzdsI76RQQnakc6GiEOVQZ2/C
B4bUF5rVHOHbVxMR8puN+Sjig+MJK+xIs5P5EsBqpR4945XZ4MfR+6XE1qMc
WAS4mZTTJ3rJ0UeBvEjO+mVxE51tH7wwlZ9vypUuq+vmlm/0K+l1QvDK0cwM
m9s1oICCU8hKcQC0cNCC7RFQYglx+c0V+JXoQRZCP0iDTi1fW++O0FZaa0su
MjxjE4894JywwaO0qvYQoXpoX3hjcqz9TYmkLOQOoHCITMjKumKxhmmT2UhM
3IGiQIkaGhuAYol0a/hOfmzw2vs9thAiJfJcMbkUGjjDHKrdc3r6Q8gDFFkC
4XgEuUKQa6S2BF59Shmz1LIH8GH8AJnjMH+OMgRyTiRgwxZpPhs1qWjR/Ar+
CJT5jklzJ6RL+zczHqS9xTKBfvvh0SSREn+GvyT6nNmBzmn139kNRApLuo7i
JC7HDC/8LLFy96MGPrpHz2HrULzu4F873wM/ry31HUhMdCdJQ2CgfKZ084Y3
L+FtD6sx7ZHJ0n3l3Gsh3KVHqzaWAZj7kHeGykHg0VcHEOFJhQr0Xn72jJTm
Qw6vhO5ZoloaYaJw604YPmJBtgSYvxFtLMbRza5rz1l8z/X8mzhbd/hpqh3k
lgi5tD1KudfT6AtS17rYM7E8QBlZhRfraE2d2QJdndAZmkMvMrWlN0TChyPY
OfWNhKMU2VCbvwPZDocS1GPfR23KioFDrd4mOJbSrY/nOMbEiZ9XDPPWu2qV
0ColDinsMOem7i4XFAoB0imzAJSieJrJa3Npau1zm+R15+tgWeMPPdWciAIL
kG9hmLuMLwVQM2kAkM89kriuhOynjDEe9kgYYrcLP0biHcvaVE9jcf4BB/kg
0cMGmbOF2tbw10id9TG4qzUcf1Qszc/c6KPnLuHI/FLIO03YYrDP9cgjidAn
x8LVMmabVRfUefPvsSeFU0RPl3BLhptk99NoE3wxNgE7kFr9OZM+GYeNX+IF
p3Yccla4rBn4atswU5VBWPm8hsGNV4pvom7L8B7W1tkbM2uaCM9gCtu/iHXq
ueMlPSt89zFyY01XDZl1oNVpgtJVxb6B1j4/anlOzUoKgnPA1h89RYehtGPj
7bpp1nCAumPYEvVZCDiTokDqFXZYI6dJ5CMqTzQzXb7zimdz5JrrenTPFciY
qCkSeEq6aBEIiHayZZdVolJPR3v+1WCwnHFOz9Pl48ZEFUjSXEQIYF6+6Js8
fTWbUFSEvwM4RwhIgFYyFs+8he57NrkycVv5oMzKtKF5VqLjlqufQwainwPO
GMreF1J6n2L/D4+0wvkHKRzkof+Zu2R7jMKIW8KhidphFh+3ZpYG0nn0/S5Q
KA5HtGtClTyAcaXADNlz6hUelJh5gkriFeNS6q1/BYdbpwvrA4BUGrlWig+F
SfUMknNAeSNgT3OQONqfUYaxcfXy29wKhRMeDWykSrNlp+YqvYcV5AwEa7eU
lehNf1HRFw4Mh+VzK0G/1f/ExpROdjXkD8NmpImAvDQHWTMSRi3B/pGFQXvw
fB/q13BlBhWxigN2HU+8l4fD6K3Cqgsv+nANspfrlYtflgO93otcF1xayToL
s8iN66VqqEoE2vBOTI7ItvzxtcP6Eq7t5gCAf4W8sZe7AzimSZg9ZJS6i4hn
3W/61l0YLkC7efG1KtdivJyrcgEB1pHuN4bXk+KujEhvHToSTKgu1ivdUvJs
QgNaC5sqUP7zyq2EFvsyKMeHj69qT9uUxg8duZFT+bmGWt+3SJPU9Xw827Gp
V4RPA47XSPMACBKLOxcNnjExePypoBufrPiV6CVo3VP994TgSfpjVLtBfxtn
C+bqVz4IPka6YzxyMViZ9TNke0fYg/68VbmmnJ5zMtrfmNeBIpJxEb0WcBtk
TLnsdtRaW6PIljszkJ73n2smTjtuNyfp1usEK9Nf6xb1XfX85igeb8gIDmck
KyuQr5YIJ89eqZG7QnMtp8tZKmJWB30mSSu09XMevC8Y0gi73IApqQuXoCTV
Z5PfxDeP7EP6CDTxZJMbBsbXzqCFkLweG6BcuBbp+/uqxhAanvlUfY2p5OXL
j3k44B/ItI7iwlA3fuQJWwcpe6xEhWjmWf0l48sYPMkWMf7Q0xbfya2ZewUn
LgYu9FbFstaYFOxpAzFpyiqZTEBkqcqv4lwn9GM2/kyDxrvyvHv7DEfZ58E2
NC+dPBqcCvjQCpKRK+RF89ClPrDhRRLvu9Apzgx/n4kXAU3ofEqaUxTbgVQR
p5nwJJLlOjv0P2rehpUQh1HSBuU7hxy37zGlgbShl/jSPWzGMYJDeUKMoyGV
bjFRB1TCLOT+q1BgFXErkv56M7BYo2L5wV86NptDuG8Rhkp6QwZrnJgHnSLR
fWu4SUpzxtvA2hde3H5ZTPNdcrLoY8TugU/qfOrimNcuSXSho06SVO9pRd3p
tv1q19pqEOqxoPy/AK57fWN16V+O2at6JDBviAqh9Yq5SxPJcqOZzBnEeydl
+rC14aFIFuqf5aL7zIn6tf6vdnw0tKjO3I3MbFTlPhWv37L9bDwU8JSvyQSm
HzbNTL2tdGcBggTXXpZRZS/xiOCke5kxJ2NBbCxMDSd3du3N6IqF3HuM0H2O
eUdt1qrMIEiQpA79ckXT7ZdkB43810jZWJtEEj7meuaPJtLoUPY2M1p9iksD
4I92ACpJ+eBMC7aX/RbuBIsqMMu1pWVDIwJIhSrmtP+Hu8+eIHU63yvWZN0L
AwGQCI/lx6xOWNHJKomrtyOjEX73t+XKoqqu4DhJR/sjaSowmEOo2+cl7zrc
jatqyJQ1SBG0IYO6TEEXi5mzwqXVC6fFkDb9Uh17VKReJPWtPuqWYYu1qM8X
HSi3sgtXB2/MI62bRG/LiwTPx3x+UJ0dNJdQMxq8MfVtG+MB7/PpqUqxgtT+
s8cxDYIABqH13+JXSjYYKViBhKP3O3Pyx1o/tLLc2nLkv+lTmV27wjosH5iS
wpyBVNQ7T2DXEN8UuaOhDsBuFGlPEMnS8XnjiiQWg+dULVDBzd4HaneWm+u+
xNTkubSYlBsHq8wh13VIM6L00YLONM2N3huUgDRhVq4aA5WO9BIH7QIAXQH2
xzyI4KrTqCV1B1XNNs8S07cc4Jp3MW05ndB0g939XAfGoOer9hj22KhIhdt+
Ov6LoYPqILMcMH1qIs00J8u8JTQw94+cPsUIaWptVlmcp0XjXHoEgChxeaFJ
4/61GaarmfxPjKnooVUl7EespVEKiI/Dlz4ZEOms/5MqsJDyvB0ld/TNh8vj
wG2kJ8mH+UW4Ceh+Rvwa3Yxj3sFMzy7OPUyXyOZvnqlSmHW4Vw5IckUbQZZp
c6ujyYBgmlsxosaAHUsCFncQa3suMaTueSL2o/7Fg31XHDxvGRBC5voZG7I1
uplX8ggBAxKsyfNgGulqAw3ZGvNRaospiJH71d+IneIkDg0i7GGhh7c3HsZA
qu/HoQP1J5m4IcuvxR5oqLxq+CZPRI9qCrQvD4BCJyQAf4ZdALFA6FgcTyxd
2+Ud4KdufDnnaDpyPfabN+SfL4rD/uRe/N7+21qDMQqmk7jRUwoBuYgHyPV1
O/JGNjRjGOnHpTRddb6M5pULY9SzMrKAKpFUDtMdF8fsXwoFH1dFLiLMxAwv
Wb6ZIbI+K5Q+ixO0RqQKpv/WHAQISZOJUKD1X+SzcdEJI4GNIr2Neg/XVcKl
CyS5sqhxAcoL0ZOv94gwPhgOG8Q17QyQWIFK9Kcnt2xZkdf51FpE/5Z1lK7t
UUfhLhUUFzZF1m99B4qcqJn5maRTuwbWQIN/81Gu5Tu3frF7UwL9CLQlJt7C
QxH7Vs2DeX+Q4Z7Oc2CbEygVJXMx0o+TVf8CI5Mfh4cpUkKNK7Y9x6Am9dCE
cTHm2SrRlGWPygbTzKNVBocUVLdGEREEU2LeSOTJdK2LQ5bR0+Y7DS9Q5qgJ
/bGyvVJoGxB9t3PYopKGGs9VeYfnQapSQUDcXjiQVqKb47T8pJyU0c/LxMxL
I5G+KG0qHbCoFyTRDvDcBXTdspUnzC/6p7D5M6ENVFiG1fla9kjRN/lkbBkC
zBouUSC8JIq0NLWJzE3KBhF8nMDR4DGmPhnL9y4dRpMgvTGh3eRa82gdDNH3
l+rywwCvWdIv+rMD0H/Xu/NUiIt1sgU1i3i07aUwxopNq4S2N5us2WR+1yYD
3+8r7cpw0hShInbUDXg/u1lY04p7gi4F5TwWIxTt+3Q9Xhcg9RfVKVy3go8Y
9qRdgzXTNdYk08cO67GkUMS8tZkc+8EffFoL6R7WVvJYlzzElerQibS1AEv9
pux77MV5eyC/RcxwTImeySY8hUVjqlvaw+MgDVvt4kmusuKcadRTz4Fcd25w
LoeIDjgkqO/2gR5gGGhHanYeqHtXrs0RUprwGaz4zCngVTureTBM3EB6sbVy
qsg0lzJ93yG0KLXFzekxE15HxUjtMew6HbaTxtBciNpVICYn857hauTCBrg2
PylEEuqm69tgsxeqSEciKaG/LIL8OSuROX2Hq3fM+NW8HxMU5xot9Rz5oAJv
JMWNCwHZUUUQb21NC/yBQOfG+w5o03wHQo2X/e0K1P1IBAmwbQ8nO+9PKPEo
TRqwLhPKj94z26/7crs52EGzLKVBboEsyHC+7q6sBtWBAEMnu1N1iYbU7FT4
LeWpyTx/10HAf077y2cpgafgxhqcy/xnYIbF6a4oAQwRb81F5m6NwZP7T3xC
T49RqRx9oOWeKnU2nXa9G2tfiAXGSW1uMvSulb9GzlXRH2B2bBhxuO1lASWK
+AkeljSL4bEbEjrd7saEVt1a0mGD+IbuAUUy5FQU9+eh7XnOsyDtjf5l6I2/
SL9XKQcWa1DTiMbzay3En1X5lalaNXdzVEQ1z90Gnsm1gdyz9IE9MgKcWxXk
c5FyH+hV5tFjTgjmMLXRNhAkEljthndJU+0HyEa+Kbyx56qV9vtUzaNd8QGj
LuuXxUd3lH+yn/+N3raEny4gVNJOUBJSnn2deGqqVEnoHXQbWhKoldgA4AYq
qUQiZkFsHI95MVc1MkYAQwYheHAuhgNtkxc20ehhu7f1C43hTm+NZZrabg7n
kIddo8yaB0XP/kKKz/aWQRnpgP7sFCCDD+2KnTYFTpWUSlmssmPf5znUw4Cd
Qe/u+H3kMF4KKr7Yi/k8oPkZX0FDcwxaRXpXUPpzkvSTXzV0ekQ5fU+AWpsc
qmjTq5eKEOAjh6HVHG+Xs50JhjCHoJL1N6uKIWxjldadgVFnOUvyII6zJRF4
95A6UbQPa7qp9lvgVy5DDV/3oUSQqaZIN86ILVgPNoDQRMSbqq92mbrFC0oQ
7IUYTehKro8En8oh8cc1FivEuPtP2ICVxY8lJfeyMGhft1INA0g9x39V2D48
87xRWbZEeerhS62t353nnS9tnSRltEuvOTeIlGVqrlYReBRLa3cK1FIwkLpt
hWkXYwyEc4obC0YF5tVnqijlgivoIuJSs8oSzncwgjDxvkO8juow+Phbd1ho
QctgJTac+P06kfiTTsC6fV3FlNy6tNa2X72pqn/ViV2XYCj/j4KtPjibz1rP
7MhOBhL8tzRNAvlDzKgbqCN+yoE9lFUJ4mWFLhu9di1+LbjGG2XeZjGA++I8
dT6ux10oNsG2r6AwKPLwOcHUqjR3fed8XvZh9oGpWnUx0ofiIQ/WyKL6bRXb
dhWrJeepYA63qey3z72GyL4Iiohf67jYsNSZERrN+xgTmZw6pGlEbdWCxf+Y
hfxg0irINvZxSVqDwS7s0/ZMLp3yZddcMfraOUtM0qgP1t6Qy5RPuQxQsyxu
73avTNyWlOnigBFjm/e9hWNT6DvQz7HpbnMNVi6pG0Qhap/diF+UByV/Gc2u
k7APb4FcOqrKND3N1s4r0Daak11X4RfGbT367Fyf+2A/Lt2ixLNQZzUPaIx3
qmmZS6z6lprOPXk7T2Aj+fti9UDDqwNmACp0jdkX49Tqm2OwJA50CE6cgdah
ULUEbqFLYIyi6DJlRwQwH9RJDmWbTN3OaJtZbW3rxPPguKqgh7dbO3lAmUh1
iR232yafEPBLOZ5YujA4W1pukFH6K7KE9kOiPcaLFenCMQQipKTGJb8xBp9P
wWpUnlN38FTR6FmTSHej4JnpSUOViNrAfMhBxBzXq+Xn3G8VA8M1Mn6eGceC
5jNWYTXA8RpaH4VmT2jnbwfP95Sq3A4kafTsAMQXzZIKYwng4dPtefVYj985
hSlNP9FmWoImNOarXMLoy/QH4r1BdzNyoEzZujTjEA/VM0G6n63vfSRU/rw7
18Fq4mfYs9dggFVfKFTIdsPNGJrIyVAkSNXcXEpu13DHIBcpjNTW7/fnquJ0
QO3ckuiVeqvoHuFh0WTmaflimsh+PWPnv6kMzItOdzlFJXTJ1wKQ4VPChVLM
mkQJ+FrbqX9Neo7TEYiYyl81qIXXbIQN0qMoCdtA07CKnv5WIKCL9zx1ZyVe
GLzSIn0svWJiz6BGYISoEhmdHA6qjeiP6j4+JDT3Yf/+TCAM3PdlhBiHkYwz
bUn5gg0TeDZ5TH9v+zFMDLZlLCqeMlZ6hk9b7DXzeUgJ5jSAG7boX7ts5IS1
jLz+aJizTGSe9D+yl3htypFiC5e9a2qZOfJw6x0FlfrYP5kkGFEuxG2qgNBi
wAHJCHO6HRG7yJykMA5C+Q6/UNUWlJCzG2QSBoYCRVovZEFY1ERchijSzlZh
vbIlp49rK9UR3//6dDO1BYE8ML6lX/BKr3oRp09JDcdr4RDA0tC6d1tWn4QE
dgafhOWFjBFJYcNPxYIXWezLy0OopvvNASiCYq3CkYivs+lKFbR42hYS2BoB
Zbpl9rVYuED/aHv3JSBeKTstYolxGH+Xrkyv6oQX6ADQ/JGqj0hpZH7N+RAQ
0MztG0lkVQbWOqr9JvZGoIixOYZR+1nhEBm1ZM3sTiFJgzp6LfH074jvWDJ5
YKcqF0suVx0YXHffPEwUUhIv3vO22jqOIwGobIQvCaKcqRHiYDOAMwvk3gU7
mAylFf9ThtIq5XJs9apI1GtvV1VA2VyiYocdYHoUb3SJ8yHKshIOWzbOLx5d
Dbqb2N6FV2GydsTVwgCduPm1MUR2y9eRwSdegsajqB00dcpkiMb8BCYbInbo
p/maAnmm6pM4MtGnGQdI6XcmOyRNXjApZ1FLbkfKgoVpHRNk6qHsIm62DSDx
W+2qLCyqXHvAdWfQFiTb10Im/q/CHthCIRTOr63NU9cf6iWBI43zRFrO44lu
TeJG6pn2ZsI+l3+DpsSeIyFDs3UXRFQNhzSK9iht27WTrscGiFSEdVddcqc7
iMxJniuwW3QyUXW0Vb4zvXl6vqsdLkX+w5L0AfDuX1i7uPBT8e6hCjCLrFrn
LFm4sLRcWn2pzr6f8uYYfW6T3FDusMw10+MMUQ5a8Feg9AqfGcwURFZzbFmW
4lU4MDXPcI4xjL4K6nSOap6iFZ/E1zi7PfFIxMc8TTmz6n6tsMysXT4lUzrW
sCZtYT74wyDsEjy4wBvh5zqEQxBiorT0vfYIqVs2NP3Dgxwh2YfbgFeH0DhH
2cwsnZ/NE49AI+qSd/ZWyyPlH5jjKglCpg7pG46S+Ro4oW22aekewZ1OoMkr
6rzQlOBGEFGLKiPjR3bfGcta/Kl3mvi/RAdSxNr9JfqIV9jP407bySp8hkvk
/6Lx42RrH5j28gItXYQcCCL3k7cMC2IjIiLfKM1Lq+POVBjF78EKhcJUtLlq
FSCd1zXRcy/1z8Lxf0/dzpzIpf1jDmylVEHlFE5/PFT0UImWfTtOTPIvLqtj
+/066TPH7Pf6adfO04aQBOKwT3Vl3rZMGRdJbO3zZ6MQzLbIYCjD/u5CRY7/
mYVuG2h7eHRRZ2k8j1frfO22azS5BW9FizQS8073GTzFDZFWys1E6vWdvo3T
Xi2I9WdtP3YQyUxJFY3/00lNaR7gy1OYdafgNrtqatT2Ifo21cwKq8PDC2Mw
bgb3daDA0g7sfPlhZwio6BNqxAx/Auk2NGNASMvbF2dwJz//6k7/x8HWZL+/
vFTUY98Al1fyCWrWSJDcVk6RTU6+XnQPh2ASZoj4UNKsCOPueihqGGwCrpGE
7Nh7CXYdCorvTcJjc03GctZ8v9NIbZBMtYbD88CXwSIqxg9GRNWGKxJMWJql
inZmnUk9BF2ItsydJFY2SqAxDT/aNc/N2mnsT5xrsVasYZMLiXq9X6QhWVl+
LdH2TZjHfYTyLAmEbrJyKYQZaoXcpNIlS8iqrMJRW48e9kqVSh37vunfCexZ
Yz5jzpproRUDhfLL6eBZxULgXtLpfqc2UvK+jaiPEzcfzbD3E1Jdm6CIpr7J
eUGsI2SPTEaVfIwLag+m74ZmdZc93g7DVrPnAwfzRPCEUK/fjGgu35pBxkzc
2ERMyCHfD65v7f9lOUyyshdu3d3gzhEvXCFJD76wgPMuJ1e/z1K0RjmZPy2g
uYLpllV5jkINsOyrwhexMm5AFdHNJ8URR04cntG1+N7j5ZKSKTeAWdiixXHS
9Sbd0duZXzXJ2A92sWgZ27hmHOn+oMVw0iaLnYJUOOJFH/8ATEqH08/gO74+
5mzfHSBzG6miP3v8RDR7qUEfTbMu8rcAULAtSF/9KBsyE6/VdRVvQIPxmfg3
aeQFq2yPGIaFA05wyWLB2bRGbJhZqsBPbyracdmTzKsejPTcl7JMDeSQf8/0
qwIKKVkYTMyfpXUhadQztCXVIiQdCdqOLNsjZrzAp/l8iiS1Qz2PkPRFx8uV
09bVgk0s7kBBLVvFbCg7+AFOOOma2ZIIdQ0DeUxl+77BNPmSj47sAhV694kE
q6NWmgfXQJr7enRSjlNBKFFGSZYD7SB3zDDuQBZB47KpiEsojBdb9brCmXL6
Mb6fMfWvwRr8tk711qXHxxrmuCvpgA/sKDxEKHZbL+pNw1XDg+a1mJZdNpyH
fgkXqTwiCChB5uHWm3XP5kTCrPTOKwWewQGgX4G2sNces4pkrmKS8Hrm9Gz9
/jJIOql2X9qDOHnfSU2cPChXZd9BifQRsQppmgQgaXV/I6GZIZAhDVNIT8qd
KLPYz3j9rEsMzPSnc/VWRrQzgt0ncf8h5fsZ0KEpwd85lUh1+PL/jqRSXjup
+MpqOWHgqaCPr+yn08nImJ2BZG++Fgrzm6HgCerv/Xn8eXfOyRtDiDl8Jp+n
4GO5zFJIWkxHacCZcYupKsnxsTVB8LjIlW5Fj5GomBIm5KFRJbdEcJRlb+LQ
GzY6bSOG1c/4q2H39NnLh53cZLcH0Zuo+hQdUwjqKfT0T7s1i2HCirdqPP57
pmbLFZWYAZXH4RUTsB0kW9hLxD+jBKLqwgaHOy/P/fXOOiXhBwFelz8JV1Ii
ObJPnlSzm67LPmG7fz2VDzr1mxksut77Mrl2BXjFO/OgTBoSl9oCBmHuQFeV
7/FWBmgrDuTDcALTmqY0UZ1duF4raALb5W/3b9GPKxJUu2RIIXjWl79MfuCz
TjjWKdeRHUG0VrBwvOtgFifNFdMoVNWRT7GmYAEO60OezFF1vxCrv/Wk+ObY
QNBgfIELL2tSoS0POfVew1thFp76JWPhbrjuau7lOtYnWKnpOE4HpgIda1iu
wOUH1h8zePu2MErDReyJ2hmkLq1VFOXrDZHxxjVWZezQIcCZeJ3ssGop+nUz
FSPkoVe/5KWRYmpQRss1Sozkj1X91RVMBANYxrW4fmKq2ep6Pn0c0DR8jwO3
pCQ8rp5aaVIFElYH2Jby5a5R7Bx6hyQbghk6k4fegPk4YxDcON8ycIcBI3gI
r6Cph12Zpl1vOE9K4IRdlDQ9Z960c6reGHiRODcV3FAh9/D0RZryHbeMo02Q
1DpYufk1/EEz43r9O1tyw53PI4tt41Sz63gVJ45Okbp8xPsW32R+t6gBJq38
6AhVELQMwmqAzEsyF3SzXFISVF+VxWtJnAzha5K6OagSVO8T3YK8XYpMl2UF
Jg8hDx3jkbcSA7dd8J+MOnrwAaNicuhxhzp7VXgeH6EVS/FdAaoliCu4K/bN
eXy2EBGhJZoShIu2LYKM+KizHkXYxzedwrxBQRsXN4jN5uugTAW9+FM611yf
ZHy/xI1UWsjPyb6PCxYaM29UKPDFZTpsWto2608ZZCghuxyjRULCWoE/ar65
U/7CG8M/tSCNPT1Qyc5bLU3ZiCYpGgEGwA8kd0K0vQUTNGNXyf6jUPyDmYuG
uaSE4NinKnkiKcQvqqR5lEDcuckokUTeYI5jfDcqiHGKq9J6VS8RCqTTk2ng
I2RxuHiEETzGrkG8K/6jvZxt9X/PORg93XhNLoKwUUcYtnkpGuyIdwyzqx6r
b+He/yzMSLNHNeXP00Tfqy4/2goDTh8HDyJ2YCaL5pIjnUUVatsmuAKpFLdz
dHqErAovuExJ1dAk9HOavW02YDE1dJskHdfFTvpSdu29nixTbor2Z3Xn+IIB
A4O9AdrK8aH8OpIHYGPKFyWk3gpoGL4dyXR1pBHpMnV6vJ5V22qAFsO+VNP+
ItgclVcdCkl/bPTQ12yg0ZJjeVbP3iNdPUh5gYEW7ZwJxmlKkiUa1oODZ0fY
S9Hy/jTzxOT88DHAQ9pqJRlL/1M/4C5KbAHExOuuxfV9nFEAy7r1f5Ve88m8
Ms4DiBzzyQS+gVkS0Yw5rQufVoKrBuzaThmk1laOQpq8qoiT5d0OB1Ik0odK
lYb5DymVWUmFjrg8eTpd5LOaMSdwh7dkRdRnBSkK9IWCKuIbz7g5jTZ7O6ir
fUhbOMwH0TWepWNsNcLJ/ZDnXZfI71SGzLTdaHHfvKuHdpUT4nE2bnoVI0uW
pqhXhyhce0U84ZJ1FFaYj4b4TXJeL3JPq7E4TTlob6lyQ+kmGU4+dUsgHeNY
WPySDyEd/qsZLPjXf5Ft63cTQ6EUK2SEk1IZvkZDZPjWlsZsEdJsT93kbwO3
0FDFRRHXB55t19CbHpf6Da/UZpXDI+/hIokJBVaazVWaoPYoJBomRLCwhaTU
H3f+3mJCpPQuGV5Y2G0k+5LgCI/iDH8TAI/mPzGyFGLsoEu9N1QO+T+YTEao
1C2CCisP1ycTwfiqKcVbE6UHwzHyABAcnn/cEePfjfyAcxpfhQ6QbOZASHIB
9RAmvGQDnGSRhL6BU817sBGpTvjM0ZRSiZykFEZ5vp8RRtQfUhSw1YkWmoM4
bmTbkixLKcx5BwI+eY9fMAB6zGRX8gH69GRLL6M9tzuVySL0bcVkC+0L/phj
E5zvEi5sfUlYIfWvafg01eJld1QBgLCrvOWwPQDwQTiO5X0svboG+83C3Kmg
KG/LTd4aXlyNlZYz2e5EC7h1x3NHCom/HsfqSB4Xulnt7bMT9yv99zYasae5
xKLBJcXCQUd3lUu8MgieJM7GMVZlfLm9Aca3wLXeUET7nwIjieccyTNxjGuF
0ZoG6R+UMWIgUGIlFQRjQANHQaHXyBdPHWgG3/4sc6wFyO8AfAdlqmaglGyV
0FqA5jJXbG9lYSyl2vbaM+Y6St3v+XDS+zRjGcjcNOn1VAvuQ+A947Wv5NPH
nHwkkgULn0MjA26U4o3AjsxJ5hYP8oqd218JyKqfiHRTYY5PNCW7gz1HW0HG
jEuhRn0A4jhpD21dlxpQzb5silLWuwADb1qyGIQYmhVDptwEfbhZHemcSmnp
C2XdaeuQSnrng6chmt/580uayrg94AAhLmxl3er286PzwuSQqSatiCetknb2
1eDNd64CsFYvwn3wn5dor7HGT1FrdwN/LBCkV0vnyuWjepe2HwCscABGwT5r
/Ot7bEOLsjpxwj0dko7m335CaFnam/Xh/nRAE6vGf9SvtAGZo4uN2QOZOugC
OcrUHyUwllHTtXQu7DA+ew6GGFFjYBF1L4zAq+4KiAY2XFcrqFbMFS+YJchH
DMs8mILq/FdLIPn9CqxiHfnIKstcgxu5eQV1CkcO3a1arXanjLndgGpt6+fz
z5s3xgySCnPAQAfxuLQlPQTkv/Y3+kVexXidQIdfdlnaqlScWCUmba+zynrY
VhXINH5eayGFIxXgkONozVsQDbPftuIjH/PjFBdqE34Eaz0km5D0H/tXtlw6
ioHLN/YX5YnDwnaGZAF53QwkHN+t0mX9GCZjqmyzjUCLH3/vrGTlKP3+UphU
uD/qaPeY90GBTnRfzu+3uxkUzaKxcMsmKIrnUDEnK9wKK0OuroFDy+1wDNim
dJpA4H0aAcRWp3fCCElHVe6CyMerIGkq0L6HsAO4ykvbQWf3R2Ny95OrC7dT
7fnHl/if/hGtqS1UAB2k7dTZr83VYuCIbkkTJB2Sr0ay1zhHCG0An31MPVE4
fyAUgslKyj1zAzzmB1yZmkdHYNIgEYOsgn1SvfdNVeoTGo1s+7Pk5BffVkMt
r0lu9YWH59DAPdqxZ9TIohN9wdeyOoI01Juy5dVqAxF/RDuWnwEJHH4v/gST
JO05KTEfBAqbrZtRgSWi5JkYD7YP1VGhrcbfD0GMgu1mNFzkSOtThlNXEQCQ
fhcjAtD1GFXGtQ8H0570gvCGwEzVWiB4sjvWXMbRDpTvd0B7wOnPoZOEO5Dh
nCLRR/mIrocYmdXIuT8YPx6AApLidMxOgNkmwKPcGr77IwB+kE1QNIfRb98y
VXCdHtue72BcIdhXLK9x3yrZOFgM/WhQY6T2RV811EYVOCb67TuLzhI4bpX4
NUUsmVw4YJGe7pdqvO+rPtf8BuYHO7EuWqLyyw7uamNTR0cQwFx5GmqaxiUi
gP9uxrDODRB2A1JCSq8Nf4UpnwrhMqSiLamKVHfwC5XaNDxmIvVy5h8MVj3b
+65jWvAtdtj+7jOBlIg/z3NYe95170aPwxs1qWVU3vIKJY7ugberEnBGga6Q
H/x1T5JpkgCyE18JoB3j6+boVXwKw+ND5fH8lG1rOBob7fwL5hDnmMJ8fkXs
lTnDyV+M9wY/tByvG2DfzNx2OHufm4Mn2Ry178L9NN94gOsP4k8ycijiaOJB
Iwy/1YkRMrvk9MmEcePrc+Bkxl1Hg0to2EEBZZTdY/gAD1nc1Hi23Dipsui6
Q72kj2BoazDukDo3P7vgF16A+sw6D93FAoL4N4GKadQVj5h2wYc4gPXD9Rkv
fo5qKMS1VxR/bb7DyxX48C3ISq08hYmY+lnLVAKfk826AVq9hofH7PXvYKKc
yCbodk3N8MM061LFVsCHEuDnnA1dZQTpOTD+TP+84fgCTdMFMqldHBF1Q605
Xo10QJXF6FoLD0pKC+gviG0dhqbqv/1c+u86JuVW44LEBxcZYJJB/R4mTele
sJaldeZzcYE7hQSZ6n1wd2wT1LbijwGQWXN56OhBxi8FWi7fvJj/nHsxijLK
D04JiOuRQjcxilTQWQ0jF9bgXufxEWznCQSO/fwDyszil7XWHzrK1NeF3vD1
ukjNd81ee8xh08Y+SRFveHgzPYqvAO53Z8X2BAQhykEoq0E3juCMRBJNhBzu
xx3l/QCQITSCaDuOmLUpdcl3RXwbGADDjMDmslpxLK5ggF1l0vveo9omCrYC
9H95UKWkwz0UaAqHcvnh+kSFDi8Ho+eNza4xSp3/axW9MxD4ohmRbkg9KSH/
vWoxxjShp6zNOAoS1vI4IduOZgjRqh3+CN9iN8cnaiobgd1GWGwFgjoO2Zts
fDJRzbRdvk+HMccolw8GJYC6BMslKfZ33etF2HThpwFvqVlZ6sB3EGQDgKUf
0cY3QNTqYScJ7G4oddQYqiL1b+EczGVayAeSD3yFHCe0RDl7fPQzoy5sTkHG
gB5diV59a05j85znUAJuDCdz0LlFfH1ERGo1DokgqfQOlTiVvLDIT1/wdGV8
a7iPrx/S14r6B/DodSTjmhYx5bBY1UBwynPG8JGZXqwIvaNhPp1zfkbuF7FU
UXijEu9ZD6M/AKpXrREb0zhE3e2osmMcqoJfXqUcut/qgmUNiMXuJVNAeAdm
OF+AE8XkKXy9LSlkrwKvIyd2DOnj/LECX0fC6rCAIyb9W6xLA8RW8O2ZwPVu
8FFrtvvZl2pzGVwBYOKyC4yK57VcirFkW0t8ToI17BoUN0CH8V52NDKP7xhV
CtFJT+e2Pvve8dqn5dITwhkAryAE27X61PqyeuTsh11jfyWo8+TGAfQdgddr
vaXBjSR59DEjWW0NazN8HeBMQD6CtQQee2cpguxKBtATd4qLSZ2vlwL32SCp
PCbQ13HbcAYMaxydWzFNS23Wi8oJlZzAwpOiel0H7uHmnFunoV1cbIKc6k2q
v6L7gE51HQ7GzW2QQ8cgEUmijMEdji/VVghwG4ZI/C17LaXfLj1jcKYv9tVt
1Jx7pJXk+fX/zloYbYLXxgAmHyqwA1RZ+fd7rTGOckSoy/jXaX59BN39APAg
EKLA8FkzXYf18+B0e+sv7QV4jot6o3Z+eAwLW5tQx1gEJHdUqFvvrvXC8F4n
+QuLspK+L1HCaz1Z9xc2EBjvY5smTeT59NUgBinqgDYB5O+m+zwdke8Q4ZSk
secaI2Zxe5q+LUyccbjAmv2cE3FY21u5AxVGBsQKVsPiG5HkJQX6CkNlxvTG
GTmlm0A3nleK0I3yqTbLEtiaVIhLOrm8tImn+Re1ZsDfjAogHfYB/RV6JD24
wOEd0jroDUnXqbPqEEz+NkW6r6pp6dCRvbsLwrieds0Ig2uO0U0pVG0u+dqb
zRe9PNksbS3Wtw4nm4w/M223/1+CV0AIICqqyVQsbg16xU9QYiipbAWWVTq3
OqP3Kfr2Vbi9JsSOCXb+A4D2UQjIbjb74ERyUbQbRRANKsJR9hPc7Eynh6Vv
2+PWfSqHTGEZjhXqyB1BTaji8sGE3+odd+02hWKYUapz0TUb2MQZ2A/ozaA9
er29aKGkmxF0iXGTKxIQGVPLBsmZ1Pg6yh95IdynJwYpWyz/1rfKQwaQFCE3
qBW2LmBjjK+A4+qC26zmwm6fx5kH7o72nrwLAZfK4CImg6QILvEqugys/86Q
QtLmmPItNV8vKkm4URQXHxUxxVpxRuaszQKyYVQEh+BrmmPFPt63rthCAgMX
p9zHKdI3BH7NzKKA/zcKYo5jlaNFMgd1DQKT+MY6pzANocDkZ10Sjq+MCF6A
85ux3B2JnYYvWfnr/eSzoLfhcaS8GBJqsy/2lfKtWvwmpr13IZ7xl7gLfFBO
h5f1TVGd66P54xEu8Ki+Ni3wzAv5/hS8i50Qa8QPUZZtUhAL4ZGWjIk00otA
VTvQ8krYawFxnQR47QHeM4P+d7BoBUPi1NB5eW8pFd5SiVM7tLxx2ldaD+nQ
VuhPS3bpDjAMPCzXxXTHJicflQTZFf7iRpb6IMJFwSx5pBL0igXjziJ7ypks
/AvAmLo5IEKmhqcTpdXJghowWwciZZmMtMcgSJXKVutPvYb3pJ1q3lu85bFp
ZYVLr/NiKLE6hmWgZpdjT7JgovOjELI7xWDqK0RAE1Yh+MYj5lZ1eBg/X3WJ
STMEHazjDPlJY7DxWLm0s8Xkk1o/2+0JhcUdjRGd6nS9rFPJddKMoeRfeQBc
Ok30dXcjmq8HVxLJAs7PMtP60+jt59zREVxFy0CYWKrvNWrNVw+8T4vJDUKy
5LtS8j4ezLhN4j0RWi8KlVJUGOiIjpqYDw7fPUG/YKOLNGBo/uvA65HNNqkR
sQKle/rsQ7Ix1k3n+ApFSLBUujQEkz+Hqxfd5LCv33Xn249f483rt08GyQ7q
+mF4NbXIAvF3mi14B7MPfdku75WHYeUYZoGoQonlbAovAYA6mFVy32Mpbgqh
qqt4K+JXnUDxKJsHGrJVOIjoIBM+pgXKpus/I/k+T35+vwHdwJnlitbKUnvP
2oOiyPYwScMMJOiQGJjY/0laW4mRiS1fs34M0/TToCxaO2cR0DEc2Rs1F8y2
6zFvIEJh+LUUjKJuAM/2wgLIjGkq9/3PdpmOuda900qFkKMrJUNmlFjf9a5s
JKNuzOff5wEHe7X4UZVdvHmWaIgVXlsbvt70AI7CJKJw2+uIDKQmRaxBE6KZ
OAEY5tdgzJP95o9PGY/1bct2LEK9qJL5jzulIBM6CF762Mcz+g70onmLTe1P
6tnkogLw61ZLRiLmNJT4W8UPAqOgcXqFXScOqDtB7QFr5MQdo9qP1clikW5q
PHHzGZQQzPTn9vLk+EfuJuxgOKtc+aWslOQ6anqbrGAWIebzdo8swk1eICGi
GM0Pv9SpeN/6PNHfO8EO9jU1WFiPbFCSuHOmZYAAlwwcoLI1lXOsP36fGuYk
EeCmutidDZPZtTOeSpSavcSL3YRa5iAHaONurRsEO93x4u3RTULjoG3JgYp5
pSCE9Xs+cajZzMjaIUn9VZvMeWcLRoTXYnEX0KX3O5W9/2S8hXxfTVgZnCmz
+Kh5ilAspvWIobHP7SfQIUTzFvbWSB0D5Stu647wadC48HHxb/CCHn6dpcz4
47xzYDIc3iirfyYSrOI4Bmu5NVFqfr+K0rb4txEscwGy9odb/x0SorvqUHpX
x4VVWstEvBcp6JH8HlQI1qXhHVAQVFbr5V7eM4oD0nfHMsOHhYu1h+XdhUsw
PFAm6cP0Bx9m9WJhUEXGWZLcV62lFFyVWjWl8tXTUM4W7BMwHdtR+aRsXl/G
4vU4WAdv7BZ0bPgwII6ONQI/DHDucFAbYlz6kGwH6pXx4CfghtDoydcu8o+y
4AlVpbhAfuaY0jqOJMZYcKBBr9FOBmPq9MBQx0kHFb0Gv9Is9tMLu/egKyOQ
rPayOzZkI5XoN1SaA1oIsRZw6UVpxdvy82v3CL9Vf5aypGE+TSOlCRMbXHHh
R5Rb5K7UYz4Bycs1up832pbd8jH2765XMrz55cXf0E4nu10Mvq8+b6hdcc/8
1LgoFsMD2+Nbv51VbA8wDqrmJ2IMJnHb+kHcYBSEAR556lvZtUKWOt+HWx0i
8baiGd8GUKqrlpLyvE7Z7Oxknm4pVa1nFYzNQS6FEvgBf9dJQqjAwjEI4lcL
PBsskL3Ph5LhwK6tZ7EiFP2GKkmoIUMHIalwPTzlponn0zA1Jg8YaimykaJq
U3jXq4zJreEKNTLB/FI3e15eqOLHCeBuYeMXaCQntxFTRhI+lbhbRn/iSCMd
APDqZQqgG4YpjVJ5+nGQSUT6YirYrVnstanx1WIziUAI9Y2JQ9CW1vrS+gnE
W2OTBs1mcWaP6lUvfTIyt7ZIEbVTit9j9Cop/fiZzoMlEsGWDIERsRC5n8ji
fXn6N247U23SH8k87Wl8r2ien5dgdeCer6Ja5TjuX2Vzex2H9DQ/lQDTd4rL
yXkxRA3FYkUJ/fJ9SWu8RiBOTBxzMA5nlmnow0ILYdWxVhDz/pDsSkik3Z05
UrGiGUDfhEeXO1Ga6Dd8aR2W775eeEevoeg3IUYrELoCHL2bsf2hslffO6rX
Jm+ugyYGhqVVQ/Fr/hdRg9323hyS0Tp/2n6UZVpFYBDawf/UU1QyZ0ZnVxjn
bzSU7ixdqN7Rz9K7f8alJG2EuvP/dwNRhBNBx143jqajOXIdaFQiWT/AKE0t
UqQdCNh7BUM4tusgIGXebKeclP4iG+oJb2Wkb/pwLah6d0Dx1Dn/ROXmW9hZ
TLITBqGHXFmvkSDPYLwR1L+A5VVrZzuyTCdh0VTOlIEd9xy21/wV9lGyq/In
2lf+OhAV4oMWIygAcT2iSUMyc5e9Bu5nJwmyzNJMP+d8Az88G6PEfjmzeE7O
cKPEn/Y7z+hk42xKrthaGM6ew+GkM5Nbhk2ml7WJBlBMd6j61Nou8lgy4R9M
O7/oEQIBfXDwR0KG5zysXyWQ+MXXPzFxDuz582NkdwiDWt17vPUNrYSMIzfh
ccB+p/5g+jKGTCTnQvr8vauDTnG1DAaY4+ZsRIV/ptn3bbp+PfHQyjuUxOns
1BRTxHJvVRDDoYlrg55/0zt1G9x48Jubx1AU8zUYuFQgTIInVO5WN1Fi+Hpd
jlOJqjPjnNs9FYLXUY8ugshgyZrGsimFRsVtK7BNJXEhux7gwHQ8KqeTP/ah
UgRLFe+j30f5JeK+QcrqYu+QoHSgWKnjxuhHXB84qGY8thx6csQ8Cdf0dqBS
SxQH7pYW55LUaGjV0wqHrw9mG08em67lUNiagTAUUVpbioS5vuVs01FRpnxs
Bly2wDFDQLjF5c+Wb7agOE+8o9SNtKwy2y2FaWsezlTCWfHZn0kVbJ0ZOFdp
PXIwIrEWP0gcIosnKCPie8L56zZ47hgSZ+wiJSDmdVVhI6AmyqiY8FiamZ+0
fLPRIoIkSXeoli8eyMzMeLh/3/KSFeewc1aJx9u5vQBbCDHKo8zlN912TYer
kT+p4HWWtKrx3G4cre4b6tcv4y3jelkEIVKfRqHfj8DxqdpdPeAxeQ7wL35/
j7ONv80F7/1DUUf7sNnnLmnytb3UcF76f7kE5xwgQfdDNOSSZfMpTr39qsfL
st/m/w/x8OnX9vFzJT0ulPm8qknDj/RjcUo0zgBuEcDoxkTRQ7p1H7+dF4ca
623OvTN7zvCDphtCoDB8GK7QbZ0Q1wV2rm5Xn5dF7tyCVeQXExj0dEhioKCq
Ez4W9ov8Er5K9pKmUhcQVCDIgIDyMZd89sngf9nzCtFwPDVNiWWQPEyCN4q9
z2yUo0+MInP0WFqDJf8lJwcTRpiAfIFpcbpolwRCO1b/+YAHAVoCam6sVH1j
V9S0NzImxU4ts8uh5dgmmoXbOYnLbMGWrZVd7g4lWZqT4IJL7KSqRFHsTJrw
SUZqkgBjBGsjf7JVHWtkaC+NJppbACz9QDlF+bMYy0XS8qxBYs8Sqk4kAZPF
Y0SFO7IkWdR6eNcHL+A8azDMWoYJSRGrVyf92WtIWa/foOkk0WJUkbFwxgsP
0ELatsiFu2BiyQdpS6RFP5zllZuoO25MQEhgi4vRz7P8HywYcbTNCHEPriQ0
Zx2OvjdeWbuTovSC08eCRVVIYPY/6rTuxDOjKe5qZAiIGIfHz4EPTp1lz8Qe
5fEPaBu0GGCuPafJyPPJFthKwkt1tS0r0QqfE7e/RDqMaaZHCSCqdmwrn7nc
4P/VAJxgOtePAesm2ZxHooA/UAuXb5XoK3DaB+ie02O7QenN1RRbl0CLkQoG
b2k3VJ8L2cmezcMm0b9wOvynRxd4ohBqM61+kqBYlf74FjL5K4iAG7XCZ0bg
rMO8tTgIuD50cfWtceBz/GFPWCLZo7LeJDLXfByBj+IeWIWmjBX7iriiqW+h
rIZkQwaD1kTYVgbaMPc6D6nu0V3Nstxr7gPP9O/21CMLY0pFc+kLzpzKGnu4
VCWeD5bfkVGt8X21obCgSTMseBiBuOEZryWbrpIIPBNjbLJCV3wKCl2lBRId
q9cH/8hPVDkUJ3F5V45gUiad2QncH7f1YRnNp6J7ep1uQ6E+39uEF3SU/XjY
lXPiDekKT8U1m1HjOKlR+UQ1neFDox/jUiNfHyodeHbgfZgfejrvZ11Vyrnb
3d/SlN8VPKLJmg0xw1Y6cVrefRE2lJF5I8RS80IgdC0XuPSA6Mim/V9adsVh
naf849IC9xWuYdTHoJTnubMfwZqh4btrVxgYbDeDpKxTPyafqUr447SxpOyr
J/9Afdq+OaLcpEvPHNHXfMa4kM9wOcJ6ER7JMswyCLN4QMAx8IVOF2kcq5Cr
Ki5++tluEcFpRoqMcv6YvGTPVoI/ZEFxMNP6YGkJFHIt21ydf59uanznO7I4
c2jjKxHXzmFSGz9HRd7Lc7vlVNyV/UcihlPgpFYnMibD87F2vw9qWu0515xl
WZsMdm7zDyfoHuK7z9i7m2Y2whrqwnXO0MZSw4Js8WyX2y1AIKZqvI7wiYpF
6I3tNBTlEACCCGV00s5yti8NupTWJtdWdzExRuhuX7gG2U4hWVB4Cj0bZNei
EctrgWrSS5E0hiJM0sZJDx6n9Ax1t9BqXMdh4s9PvmsPYsXZc8BZSQr+pQJD
Hdu4MU30FZvcnL/8rzgAXI3n2Ch7ICzINwBvVuqSWHUd8U3LQFwhQCOukDMx
bjW//1+Lmwx2w/BNBR4BDN2/FU7kaaWpcXoA1rzf1JHtbODERKKEjRNssA47
6nmYIuw4Xl6zRXMzdy+ozdWru4sieNSLMQG1neNPlkzsTkwB8yr58o8fSUAi
j7Y9U+QnWDQC5rGdUAs/0aRccQmgyUlT9xfH2Z5vpF3lvFTzGJHaq0tYNmo/
vpW2SkO7Ge49fP219cEDNicWjrTHjQwEkqEclyjfFSBiAnhqrwPj7IdJi3H3
TVEb++4W7/lwL8iRIjcY1l6pg1EmE/SaBiCmFEgPkZBDgDm5bbmct10PKxC6
4CSnC54xSZGxuI7mjfsKB/lZwCJkAI3qH1XgcNImSvB9PvAy3NtQFVzFZLVO
TiIp5kTUmRJV99wF1/pcKCzoOGfMyaXRnA6yjhzgh+uEzllMaj4D4qf65WLu
Au4EY/EYckJbkBj31RDKbEsbiM4HnsowW0PcEohP3nppogLMoqejz62Tmw7Y
e3nHOJUtmdchEzq8B9Y4eLckvc0udnEZ6LMla5YEx7twJi567kt89Ix+dPqT
vxBY4xW2FcLJd4un+/9Q0hTaGjFFGCbLWFPoKSY2nyYTJqPDRfNPOCjjECRS
+b4YYItWNoHisnpRFtdJWjBr/zzCQIpHBa9wF+CVigdkMsx8ycBkavARWLZq
dLGifozcQqqrG+O9b4VR5+e1QzSzLiuwZADaY1kn1eRDO9E4JNM4rEE84Tat
UarY1pitkkaAj8qnmtLQJU7XueKIeTFSpfXxnYtFrlwEVZ7Q2lf7+RpCTgf2
4LEGRMERWEx/hx9U7d3zwXYyWjL6DFmRB+VABFXvp6VUItFwUC2ctOBbCaWM
wPeKUdX2orZd4QnKtM3efX7Me8cN7DbKlOkXI5dRmxyH5Mwd46NsEbkjYu5E
qyscPm5tonYRT26xHG8zVnz2kdZRO+l7/8h2uwq80nnpDlHNbftElRsFmC6Z
M5016L88RN8baJ0n8AUf5Xv6FrJVAUVaXRIMm5TXSMggoCdrZ9ldPlQ+QjO/
WTLIKPQKTkfy457khPgnrPBiqWOXgiZxafH3jJj3icTZdpxLPcRPVtU2E094
Y2r3hpwYSEB/OcuKeIXZcsCW4PJIOIzSO0VhyAXxGuPZ+kTfJc55CmcU6rjB
YD1PcKEUjMtRlcdaoEBvtHzD8x2AsU2IVCR2pJL4RdruAcBcx9iVFCL9aX1N
osNXhFISOJEyUsCOGXtYcbNbw4dL8QHElQnY0wff9gBaCbH4FcXZc3r62Q5I
6+KTgWbA+hnegzcEn5ZlUmPwAedVRgp+jZvgRMXG2J4vQGBkKL+VznJ5Uv8v
D/EUiJJsMYeFwbVhU8JNEjDd+LetgKTKsMaJf9HrrMfmXDxKU13wrpYU7Cn6
naRdEGv5w8j5ouoccOwAcqGlhJeqkVCzx+wiYDM/i0aZoUx45BctCPhkaAQy
a+1Ag/2/L07KSBDFzSeRk19WA26M9BluCy86XbLcR0EO7jM44gQx06lhC+GI
JLty79UeDOPKYaaNBXY4Fp4C+eocgbxK6Ag4MZXCiRaYM472o/1P5k279UVa
OqmM+zXrffgr6ONsEzgW71R+DgHtf0YL66rbjTI8KEcoQruSDUeiAc0fdlGz
eTTRVuuehvs2XNbu0HG4RshuEY/i81dKPLVHQzwxaPw8qEk0RPEis7TLCqmt
EaH9YRmCc7LuaXh/gDR33CgynyGoYcgRVu2JaFwOZVWNy7bIOx5CukQdofUe
AvJAAuHHv4kBgrlPNZJndJQXnNbJfu9G8MP7IihwwL0gnUQkXcxpPbQ5wuNH
fJzcCHxBDHBMWcTK7ZHo5ebJ2yB0NDOx3h7mBXPZ5Zx2j2TRlirJDWHZIWXf
g2oHS30BNATx0q5f8t48v76wG/veT6eDhj52cJTKTRhIVaRWTE5cF+AIiebe
OgIOKfnvb0FlfGGLKtjdWxxH+1pRxkgghm70RvATfTMMk3R7xZYepLbJveVi
wqF9o8zHInaxQHbG/FtrYI1n9vRu+n5WwYMldAsieFPkYLXCyE6vqOrzwf+w
n/dOQyxF2OMZRs2xsKXqD3hmWjb10C906Yo+AwDQA/IeQo5j3mTMbLuo1Y8/
HzXebtjH0PVpDPAZNjguuHZkt/1HaI8b6BSUVaEFPw155XCSgOlrF4uzJ1n1
h99DKOFaJMTvHYBPX3n22Af66T3fcBovnV/QVgNA/B/19KW19og278A83yia
gr8QrEPUZtZnkmrajyODvBSj703rzJo+IdaO/mvbPLdpsCTUT9Ytb3UGcoTp
wsycS/nzvhfQ2QGqNW2UHSuKqqBPeXhHTwFgKp9BdwrHRiUKpCNBrDfu0SOs
osab87lABC3gxZ3yyiAMo+hbTKZeWvDSFS5vqiF2TJOXJw1n5rjtoA8jdKxR
4uaUzhpLCKCphdyKgQLQ0zKjr0ZeNGm7XjfzmUOnb6CpE4Zgfyk9d+hLN5am
7t2tORJIBQg22od4FdZJBqDggUr+DAWHrrkJEWPg1TQ5dSGEVBj7YCjDVJdF
sGkUdPZF19hNTDpBWjFXqh0BJYnjE0jNgznVo2PNsb9/UrNCBVSCjYe0K8Zf
rElkTlZr9u75EsH07FNyMCnAf766XrwtjgcVWDut6Psx3qB46ifPqalvbCyX
Q0Yr8/VP32LQAc71MWgDwtxC7FMsBokGRiUy8PK7iMzayPXWsdHf3sMli0Tl
NuQHP2G65y954LG2vMXN2f8ZKHMQkjGsmvni9NCHAyp1PrIE7nmDvDP9lVCW
m18Aa1Xdi4e2EfotULmbBxsoNb12fFj1qKkte8Mbm3SfhppiGUN5aZXfI6VB
D/2oz0WHEI4YkoYAaTyqumZzIgeDWY/IBh5xjhBhNeiFlz+y4Ipx2CxagzO8
3Oo7dh+31dsXKZ8dj/UJzA/I9QPk9sGR2EPxfRX4gFT9FreKmEB7c/6IwzF/
nEnHV3ZYoLDWvwF4j4zS1uCNMfAOJ2VZfdZyGowwTUurnBzjwbkMVJ5qi31B
PCsu9dK54nOU4Odtq6RxKCdhwnG1Q81tLGWQLDB+PwCqy7vJfjlylDQSKHVl
laMc/RnMrSHpJA8+UnUjRbNkrvpIYN6grvmOg54VpN8FoPA1w37tva5hKCx+
rcjIPySf+Q8cTakz8I1hQ8HPJmcnrGLcwGqmq8l14oF0lQXiILrbAsZYgNma
2ZhwyeJjU7sbtEUKdtE8xr2nEKg4IN3jT9rLR/0NB8sF0w1kUnvXRFLcMj8h
0AExXYE5osqk+V7EdUsA2gcIM5xhXG7HDE9uQULhF+X1C81V+zNMHcsOeXMp
iMEl6I4YqD3gJYg9QbNyGI70mdpAepq0UVxD9p/4V5g76qxYTIHpViiUMFqi
SYaxEYJyeachnxJFffilItdLI4nq2LTriPi6dEAKZ80caISmy0kXgAdwVUSs
eP7r/MbGgOjRid7sReSobfCZHEVCAlWhQMYPDg2yjgQFVNLyNA1EVsNnrpPu
Iv0gNdvBW65yqcF/QnJHn290oTz5qSkvyq4taK1gGMnvWz2tbxm2Cdy6C3uU
o1kBGujAMVnFfGLAgbiczBS2yyZn+eNyO8BmPB07qgADfyddPxDX3gE7VELw
hznPAkCJL0FlWHvWQANzmBPyLrSiHTUBYho6MfzvdigGWA4FKvHcxyn1iwQR
sfzWrxw2tWUXTX8jLi+XS+k7XGzC2yBcz09Wjr5UgaZR9F1UHJldJfjFGs6z
RH+ACR+x0SjmkRS6ubwoKha+ktjVLgV83dQQeBn7yHEqDTwlUBrmJ1wH3dP3
s1NT1ZBrTBhlAzFUnkscDGTkSSwcgIohvTNQOp7AOLXoHBlfbHvZSJBjz4hf
4KllHOq465rNR8U5jvqPBjYDO5g2ICE8KftJJtRPAh3Zfe3XwXWDfmRI4Zzt
tQxTN4CNr2WA2hm9kfoATeq4Eu0YFNn7C1RBUGSRwSdaK/GcGug/sCsezXxJ
9kfn4sPqP07dk8zfLUp87YgEf77wNe5KaL4R/axAwqbCq30WRI6+PLUEkTgf
Ku1LOBSHFUvVeeSWGuQNW9L9iaQfPMWL53Hqla/RdfHPw0QlazJy355rHw29
yPKgP+Mr+rvKBpaoAbwuRwky121a9NRn5SADqDWHr87YbC4CrmYIxv9ePKK0
L+MK42E+YV8S14qVmgeXt7DuKHhSlLtbMiwW0vJPe3rXIAdhZ7hRJBdh5gQe
3ZqJqcA38ep2cnqMGzMxBj+VLVC6ZrkpHoaWbtOG5PhlO7rnLhBByGL6j7IV
FCkui7bXm3PyEyxRT11DVU4NnYDYHQvA+UIv2snF7nR07zg3LwH9Yv0JriDb
ONI6byIBvN6JONGxc6qiSohqGDvFFX4UW4NVQis26oqkuTIXeqqchtpRNpYa
K2B8Bk7bPnKuUCYPgUZPdHhW+UOi3x7JUhuPSUE3m51WU9f25v2uUbi1bzCV
dXsfg4YGMTpfsjVxwUSfJfE4PdK/wJXUnWMlstf1NicxBZ1YGMlflpJctr83
ui/tzyb70bptqlCotDkmNglABDB1JHm3deZpXrFaE9ias5+aP9QnFXa9n1//
1S/eDaXn3+KB6b4eVGxuqhcHSKDhT8uDWNAjD3p8VIgeFhg2riDDmLTGdi/7
+hzS4TV0Jmo16QrEqeQxtKkMIrue5EwthFbq+E/7CGVqqDg6pQKA3BaLuzLT
Ufah8q4ELOLx57fWiKrKMtXCKTpUJ55/SqxBj0msDAaoj/B2D8oL61Q9KjgO
+MK7KvqCRfMwSYo+fSCHjiV9kHKKtTHliEfzPIPrD6Go/dpRH+sN5si9RVV1
ROV2bxJWboB8pc1k9Dq0V+JB3HNFrZRQ1E2YQ4bXjVv48tJGy4FRzTb7IvW/
2XTcKDxMaGpRKkA1Rfao1X3Uc9bSbcZh4jGA4OTIX4NogcGT9eRnJM7uqW7N
/0QEl3mzp1wnE1ggjlgYtwJxiCOL4xmBMqjK9pHk1JSFjZzlCfDZDd54ev3p
nREHZbSCvCG4gMIUZlpHUj8KpQV36qYSohLYuGEwzXocn5pgDlgPqpzG+/JB
wFVqt6V4LOCmdET1uaZMCc+6VkKIm9bFjKSzLS1EVjzgZKpSNxbJJD0Q1woG
F52zspsluJ6nOWcF5YjzezHhYosZiXrv2cJN2AiyBo/B7YpzxGdxkO8wSKXl
ORpebXPo1dfIrDjEIZOk3lahHkeArOJYNujSoVNk+Hi56DPmo3VdNlSXR7UL
p2/wjGHeIDFeZS6xoOk8LoDLq82P0vq02lrSrnKfRf8EftS0w9hdomX6L4re
peeYHdiNAuIhxDIZLLhY4Ei7CYD/zasgoflLn075OAT0JvRg2sNP9NmzqJTG
l0WUZ0wPQp0qSnysMDbmWR5Pbh2/v1N020TX0bJKXKZSsVkSTJIJSgwz5TTr
xOJ6owr47F15lbJKqllXl5CABg/bitmOGVvxv49K4VpBULLlQVVVBJLFOZWn
nOKfBW2iXiepCrdvGDujinp1FEi2LgMGnJN2Iego3mgnw5g8lYrTtCCE56u4
Qd52zlxsho2/7Z8Df7nnmt2s1HZV2+ah5fJsQCn0sVYdBPpvptJsbHlvK7KN
Vj8W6iNKrgNREafg6/8hKU04FkN4qTwYgGl/EAVJ1o7dNcZQXmRNvC9a0xjo
5/erTga782Vs4Ea2XOXhU3bK2g3eKmXEGQ/Fned3buuJWGAP+imSCcEZBnzu
F5AtyISwu6ww8hjJYOa4awKI2Vub3cAAMK47qAYUWQa133UUFJomZQATCuhQ
sywfunw5wMAbtRGWJaWwAqGVnCii0/KLTze4OPvArzj7o5FVlt7U/mZYcQUR
nIhOC5uRUfdNgB/FcSEg/8APjw6TPnFT3Nzte01sJB0TRGhO8PN5nNFFJ5ms
RiittDprlUMPIqbATypDodpxbxn9mWk+/a4f27o9fwiQWB1DHBF1oSUABa4o
FtK2wbqXJ08ZJ0rFmGwi9EdiKOrHx2gAtsST3k2eZzKSvScUae/aJuiVENqp
cNC3XqesvnB0re6SrwPqDTeebYLZVkLwF5lr18DtzIknC5y6b4MgMS9hElxC
sQPIyqpedk+Kbq4VoHELIXceM5u8keF+G3/hVJUjqzP6QSu1We0jBLWI0EFN
VjsD8rO+E5gE3wrcOlr5yUaTKmhfJSn28LmEhnWmqG+4BoxTPFMsCM68drx7
upT07msh7aiJM0GoLeJXdNF6DQMvv0PXbonKFLzrpgQ7sRZvFkU2GkT39jnp
UhJ/ARB+QglQ5TUmtbbOod0/dYmph1Rt5APcqbumagS0Y5kPpjvo7fVoUtGe
6r/pVZNvCheHTGNJymyQc9ZRX1aoCfrTGxy23P7E7J+jDCMrZnUEASwJvATK
xrAEtac0RDEQFSZwtZljHZxexxwYhmsAccqWwV5aKCrp1GqCc7MOcs+IE8m4
alsUbohLNG8o1ZXJkpqQ+LZlKcu7nHCZMmDFAHXBDsmnPRnrlzGPbXSIQpi2
XJZVdWEFh0Y9DtCLiJRoVvHpyi6TBBQugeCQllM/RmzUt9CSbybxh/gK7T55
zz05ZKvE2B317R7IJANamYgZi1KpV2yi4g4XKI5iaReScnZ//EDdPF6QqWkl
G11sn5snrkqueBSSc47JFGIHOK9fcltnVf/ldMgy8mLFhrIN8jvzkxtlu1SO
8ZZut8z33+psktm9Uw56/8jpHTq5xpd6MCSYUxHu1bdhnY+PzUtOPU+2LoH6
qfu/Uc4V953vvTArd4/UQprEfKvMQiohuYpYmmVLKEdVC9jGASbDnAFfsWqE
ObzgK+fcBq/7KT9mgQhPTLFVYnHkNU90yPE4FeETo8qFfuFhwpEx3V4kU7eH
NJ4iaTUb+Yhqkuuy2DUBouczRZQyA6euixM9l65oHsU7ecX9lQI73PAtExjp
YWpJQcuY83oTyLa8nTNoaVfE1sDp0uH0FQMPEko4sCPN3ZmAlEIV8jA5XafO
GRyGR//pcvfj6vLLW0FFKkzJysb4rQhXF4nq2kpcR7ZaTcM6JEbg6QzflVnC
l2zEDUlHPtjrMY0DlD/GDvM0ClXaqeV5++2+m1XSpVFp7PQ72ALrK2PU494E
Z+qbBAWzac5GegDdPfGuV+G0W6AA37aRmptJU+XJqfppre9HpNB+P8Zb9+3I
SF3Pm68ok1o8RURlQUl2hWWAcbWtkqw6/cWoq7CLqwckKPs+y5fZWDKmD7g7
0Qk2NW4Np1+Dtxr7llwYMRDOID8rE87Bp3MOl8mo0VqW5Gpfi+/wN/mQC9oN
KJMAYp+9aJAqCMynm9aiO3sVmABn+lUsBZqpgfhL/TwiOygqH+ekz9zpkshm
riquyRFTfhFHGgWcw7hBTNJk8Sf969oiBIZmdwBtgSvk+Hk6fgyvHBu2vEdR
pOguzCWOeyCEqk9lx1TcmpzQhKh61zTWNbCqFriEhiVCZZHhete++zqHeBqP
AoVF6318N1Gz1blwKpr4L8Lbel0tM7NCvSQyUbKBxnLNpEPDGG80ENJO/qBU
PKVgC5FaPMeDW0XlM9ySdyJCyNOgEvB11TbJzbIew4I4wl5K1XJV4gh34IPx
UWz0UfrNcIihFiy1NUSENiW98vYYcwyKBOwDS/a469GgFIgSk36ed2HCWivV
M1NccqxsLsA+BLAsJs7vDTz2+g28tYkuWPU5yQCJ84/MT5LjicE4YabcMXUl
PN3lKTFN7MhTK4ziQVXGhgvbNmi7nWNG1YxHtjpQwjR32M2/dxMpb9Hq3Q/Y
tdFMGjAELmFOr/n9eOAKTQWppUWXo+OjoTz0TihUMhb3vcsrJcRsiCruQOTL
Z9vxsLtteLUVIH9oAWNXFUMQ0AqDgU8zNEL0KPkSHQJMMw4Lmg42QEZXjAoP
Jj64RT6VnOKOGgAaGLog1QigjXxkwf+fuGP62UvDDDhomRNLrVVpDBrYO+/4
Q7Qgd+/wdMyi1i/kCBt+NhZp08jBkUv8/m3WV02D5tGWbJwoidN49ntQIcGa
KXjjosUQ931IFaphJ73z4TtkVGIiNfyo27nVxw9AxkMACM2RHpau/DkPYfK2
Fv+NsYm6PkQBPuv1Z2CRg/FPBcZJx2emfGYsDNX7fVEVKOukBiaNvnY3xvjv
kvt/o2vN1PXzKU5mvye9Nzxkmtl0zl9T3FoYB6UK5axAF4nVXmcaaaQnsyWl
6vw0fYiL+7dCjKI8EKRal1r6so9T1HMVvUEiJJcCQsrP1fTPNie2pVcqfiVd
ADId/n2dapQEQBGjDWjCIUlqubY6W7AJkUtyHX+41DjuLRjDD2Z8g59po57L
xVF3vOOSe3hqIPRYQoh7FVk60CGcAfAzaCGKNzM0mBFuFkMrH1WHGArB5vM8
Y4gx912ne4r/cpxUsFb51J5lireq0norBv9qhUyO2iZPVvm1o03hmn8MchZf
Sd6AkFZXv1bfVV7Q8kMw9nFHEFcnAVnVfL2z+QLy8ERCde8FHuqVrqvMKb1S
vl3+OjU3zu3RybCAJNZqPlDPhCW9AgeAfJzRAWhxeWFvYbc+DvxwwU+3Oyzo
sQgwauvSL6rPXnI5drvyaTneAW5+03ZO48V+bGcrsA0cfnwdJv6dT6owYhUH
r43McdrsjOGDoTDHyHWGImmfFEPZCsau1YHtSgIPGucP3H3aFUffhJ4msf4S
P/0ynubjZ0IVxO85/McQP33uRAlMWcMrF/uVpiGflTtg+Sw2HCNOcRF7s2c4
ZJ14VSwuHliOgUA8Og9flYxVeKgajjl6yk0ef2Ly8TWYsdP6ujkaIffUaATM
hkq51GI75A5CjhdeF3O1B3+byJOlFZA+i4X191gtoFOYIkC1DHeCwbPwqJZx
P22tmt3uHkdiuqttpgRWDboJq8bUHlK3K9l60jUkRFt4IyBrSmRnFTOEt9Ct
K/OAhATymZIdhyl9G9CkTES/vUd/5lr9HoywqFwJ7/CYrUr3yEtqSnzZ23SC
K/3hbg6G7CxNvuwbSQSJaoy/bznGB9AR0Q4hr4WQhYb9kUviYfw82f8Aage0
fNG+WnQp+R71j1gr5zi31ihFUx4G8Gj+Yfnz2g2pOpDTBjcv2lCvRoYWvFM9
BNjZ6AW+B70ZRF3h/c5gHGiDF8bMDmi7Tl04TLEuOtpy3SvZC4GamLpTOUYw
zdsTDRjOlZpPvYublu3cqihz7E563HoMsBlEwkMTDymNEdKVFkEv58LyPpjc
3g0NBgkwBy5JrtNVoR/PSxLw7jErLznN8hq8hfnCIfipsEaZZZwP9yCrpd2E
/E4ZxIywR+1chmfjAMYCiH0KrElgakSuRd9/JslaLd3qUifQbWwfCzTTPrk2
ops/Dbx65Xa5YqwUntgxaveL++0LDXbw3ne07m+1czjjW0Y6ZUuppb0dCvWc
o5/HoFEwI00gcOtARNZ2DfKs7TnlCI1U3lnpq78a1njt/lwUKcVipLCcKD6+
dlZ5tye0Qc16TvD8ZPmrCtQb1b4OJiSciGuC+q+gJoMo9Ik0WCrugSaOxjEV
Qit2tiHjnECy93uG8tCl1/knEcMS17lwIs520Ia87dPfq+79viPvRTBglE6v
8nCVg4MUp8OSiFkZnT4dz54sldRaX4RzanS3cXkvRL4eno5JpTW+mOgXvLsu
1lm1mCugI50LGbrDh95V/TEoO3bTgHwCF/W2uACqerjk/GAB5zsRFyOC7PdZ
nTYm1OHjoK6ySVMRFYZP4rjqDNZ4gwEglCN9zAfdfnLb5jMlgXkk4laAoVFx
yMhehJdUmpgxJ+urwgX+E5Ldlil92s7FE4waxNsCRRlQV/WFGtooAyqpsLvK
cgrnnqKK+//QhDEA+c3s2cN9OID8y774WZ9VB0fE5krmjwND7Pm7rD0Rjh32
lR7cmfaOQVzzEjTREI33e0rjDmU+QG60Q2BNWTmI+UO9PAt+VjS8yL7aJnCJ
w0DJNqnLCs/PkLLJWhqlkufGOsxHgplcOfFjyaWYK3HJ2ulG/AhRbuZk/KYf
OSlPvrEIvc3sRu5yEBQRfeTU2hDQMMXi/1VjzHd/XSpBXBfM0FJzHfZ6eh15
OGpROj63WbMixb3Tld/X6tAr3N+Ht5QVigX/D47YLldbVIuBRLOfEYWMjLIg
zCugbDkIlyRcvJm3ePn1zdKBamjPHTqrDp5eLaYLmhp/5/OEu7Nr2NIl3R89
shvYOeU5IxDysMbEZEWmQJhY8wItH9Ilf+nw1EOpzyN0ykt6jN/VpZdyz3rv
G4oyaqMHnEwB3ub2Dpd1GBWdI+GoMbxJBoiFbrvxjzljPH5BFX69lKHCWqn6
In8HEB1dHIJBHkBX62ukNKX91MGm84uSj6dIgAZf+dxRbbX0cr4+Z0GoKz4T
th4nLx8z0Oao6OV0NivoL6QgbsbW3q5pIc6gZm8y/4LNp8TxM9JXn3jJWb1B
wxIbIkL4USd0qtK0I0hejR3XmC1iGfTOXUhfzgupaZaqWfklsWja/1qeE6di
MhIbZuUA7Ae6fflbtbj9Ew0ME+H9vKVlVG36P6wr35B3C+gCXdxsN6RgOgEC
68VxFDadP7O6yt+wktGD7khk2kYWhyYkgKn3UlcWrJpA8m3aJSeERZ+MJsGa
ZIswLlyFuS60alCYT8MW0SftRTN7dG1b2OsaJ7t3dUh7zyvetq5nkVWP7BUl
TduyI/A43gocam02+5/TezztwWBawTmVLxEjkRdPtwyz1nE956Q+i3G8WoQr
mDD6Q8qC/tgB65y01giGWgPtlIipedWMRV4PUqoX3lKKB44bZIw+KBygVyZ9
q1VJ0Y6BX9ej842/Rbf3G8+xnc7m5YcAyiGXlmSMPx5HH1INOfTqWNX1ft/n
y1UqoJ2En5X935c2207k+3Utz3EdfQIXtljLiV/2UAH5OTO+TNg3AJn9y4Mi
8G0XbE6Ly8YLJ4kL2XAh3cdVw9f9RD2+rI+EyxCqgBkpvigeoPsIa0BMxvwE
Lz0t/l0qehOb4yusnJUr3Jh1qKKNUN3kCqboLuKGJWSjcb/X+SSuQqXvbFvR
nEjgk0rasRv0XfbMnfnbhtmugPEDmot9uNxI72FTuiQzXUR85qXR8drZocgf
hxZXK5NmoEHwprSsP37O6/WcQ+PZ0CEnsxGDCMOJGaTh3Fyq/1ahds1+FpXH
+r7lbKs8S+EJZJO094qlk6PXTJoeswESDNLEhYbkDSkZVqpNlujYLPGla5AP
hcM5NhfFXzD86dlkKJdLQ3tyQm1C+ADZL1g/mUrn9ugFb3OyByw0CiNdxRns
0Mt+aZXB5AzTP6jEC29lm/zU9tl4VrYMv7GDJ+fcU17tJp0Pw37g/Ov1ud1W
1n/gzdo9s6fheSynA/24r0jIODUSjHS2DjcbK7yJsn3EpkA1ppKGl00Tcz5n
GWDBjQHFyibs/Lx0N3ULJeuOjIJyzhKk+HQjgr+KYw/lGlSG9A+1HIaAxgBQ
8d1SGvwveg4II0t+YJvccumpMDi+0UsDD2jwNS8JlHrGE0jbHC1uYsR4sO5i
tqdJg23EFjnPgWjPAZ6GP8+nmrjCF+hgPK71ZKL2d8QIGXtdSC6kbP9kpD6s
UiE8yVcArk39HU33C19DNFZCwcD5XyRvnauGBJea/Kq+HkJTMsmebLXY9GLV
18I57w30INVv9rylvnc5xzzPtVAUMupetijw3vlUwl2BzAMuj+9+WMF/OIc4
qPz8RCVwZ08ww/DyJEzADZV2I5rUTGSz55PqBiFr1lJmbjZG+1+eILMHysSz
CpbMRUDSFwgL4PuPmaSWBD8sGX+wk7ZYbZF2zb/PIZ5e+D+y8jO7hVV6ZFs/
mb4orJ4h3Ji45COHeLsfniNhkn+ywchUknxB+dnqKXS9Qszo8By/frcNHU99
+pTP6xfHa8B6HlhghTzCMvi0+d81QQ1wcqO17c09DvW3SUuepI9sknLEP+Tf
Ke/kmwbd8ebO/dCC7tWV0nllVlMkuk/+xhgtm1/odeLCBDeoe3mf0Bzjvyjz
ikExSDsj62l/o1omzIYxIMVKZze7gNlK+Lsh+qHwz82+N6PzWdL6mOyyla68
c7NtMcoxV9+E5U+jCDGpZs9Djod9d+oQ9cU6iZAdD9EM4Ql2WebN2n5/TfC+
RZkTY5LE9i7suHAra6nzHnv9DL4lFFd9rhk1hQz6Nx6c+RC3vBDz7nlXbsFz
oIju82XKAWPs40cZS3rYgAeuO4IFXLoh2yqysdkQeMAaBmoY4qNoM34plRka
WoFVTYp4ilgrBemdpGPCQHgFqCWt6/dE+h3yQEaTj6qSbDcUXWxRPNaZBMgm
o4XBeECrLavnD8P6QpK+VUK0clrMjn4v8G6xW2vif0mkQy/qysa6oZ1VbB7F
NitvL/DMNs8nbM0JVZ8ZmoXA3Z6zcKQeouFiigHPehzOdonzI8/KNkAe1+ei
CKbWYEE/xtxlMu5S21rKQyFn7+ukbRKc3IrPBMy+BIUKXvjAI2gj7vPeNihx
QZOhD9sfR1Ojavk0OM3ixaeXEBBuxiawRf58YACKNDrbovlnLYOqf9RsCcfj
cCf2xEwjVOrnTdAWrT5yryYo5UVAZ2mmWVuFBwaZtGfsPGjU1ztKYhOKEhRo
vhxLOrj/rHRdkj1hm4VMOyMx8bFt7FA8pPmKIoFrhKgcdmrhuZzmdcq3hmna
+ghPGZpFB8v6NmGglAekeJgZOY29D3aTgCpSMv0u20xI1hIs2szzmDGXMdoJ
jruxGCEg8uUzFFqZfPYEnj3ODshosjT+kZvOzX0eqHbqrIj6FTjvmy+kwxco
RYgr28o038x+n5NZ6rW2FO3H3dWdfNIBcYP6OB33tEIyO/Hnfh9AGxODXFDj
5/n5SKQiwfKKbWIV7dQKLQy/6EXfXhMWDZjw/b7Roi8tixJZU3OmaD0AfAnR
GNIcgYiTHKAzagHgNjbL7g+jOtjLK1P85LBZO+crfIYjcgWyK2hb3bOy3aiK
MZj7l/QEgNS9UQLNyku9mQW3bkqbQKvO+X3F/XOW13gjYdfiGMg05kYTH/xk
RgFmMGgBCafax1CH7B3aKqvh/groujNc1S73nW24F7P5SOeIoOPalSFVVXg9
TKUCjxphMCHVxJNTlhbG6xUg3UT2T6xm2pS4q4EeXmEHPAbSClm5kJSRgWPb
tbGzOHiGbP1SYmt9wtip32f+dE1z+ViUAxattduQQwPMNhEQBTc1W0GeZOmH
E7zzahmMMpqGliu1ZVhVQIwevMZJB5ISreTl+xxFRjyVASjbK9JHX8MW5Y38
yY5isKE6YAcsxG39lBF0NNbYhTn73LVzUnwK8oIBkT/Zo7t7dnLzT2M+l98D
xsnl2lrdkbhna9q7QRCAp8i5kAUIBYZDUIUJ/svKanUubPaORGFabXnxTSpD
PFMQ8emh1jhcEMz79yKtRKJLQMeyvMQzKn1ye3fNR996PHkq9jl9gPsmoiOw
xE3PVvwO2qO86EGjmS6NUUiMLnPwFJJz8rhG7zdDpaKlqWI59lKqAjWwnjtk
kYLWnsuG2lactW1EfgxqibBAs7xeXEyitmrpUU9rUPcczAumzO2XFtwxHx9c
LjdRcqHZd0gidFwmU/1JE/aBo3gOSa9pFoZ1dm7TQlEmBdQvW0fXkLR+wuaF
EZk+Il2Kz+IP+APfZNcV28zj9wYI1MvnyYLkvO4LkVHN99HnjuUemFb/LVxe
JeZiFNaoKyZl6bYnO9O07qfyamGpXI/iJ5TtEgLVkufT1GjMjkgQvVdtdnYh
JvK68xxbRCkncvWFxJSC8pz5WgDDxLsvinS5sXzJViW+VvP1512n7eLdMACC
KGHFfd2TxIC6EGft6a3AU/R42dNt6RdwvH63v1A5ruOeb+AjK5pDBPcG0olU
KOeOThhvG1A5vDHQhAyBvBKN5FmWxNKK9mqFifkkikMlatq6XwaaUMGJC/vB
weh7D2AXIe7QDOvq86J3fuOVOReiLrEcSHbQfoYG9jbo7gICzVg1nXz6LVk3
jKfEnO2RHaY8jf2SNl3tquaB6sFmGqGQQHBISCq44GcnZqNC6hVxawbUeg50
IB2lB2vFvVYbbftTSjyqaWWG5Mlz+8SpIUjXX2IwZjXnYwMTJkZg7Io8xQhV
qDSNu3qtQIBHS0bx96XXSZjqhg+eLRpBlnD8cf5fg6c+UAege0zYgdqelZP4
H2FG4R7WvUu+eQ9kP7IrRfte2J4IIzu1HMKfsl+dBbW4htkGP5+g7ohUNCZU
z9qxo1DOvxXczZBP+7J+Jd7iWtJxhS4o/g8hcfkpyWh7hJXloWRNrpdG0h5e
RPyr4lsV2FusXiQzCfHyL0aBbrW9fEs/7TZzQeuWoMvicRxp1ZhychAhyb6R
ULcTlvULxQb+dGjyCjV0VdQZl+Bu+ZN6ltQBkK4nB40FqMQvZ/1BLdyJL9Cr
ygR7f+Fbwd6kb3qIvX4Ag5gxbeVSxwt3C/MaUWxVJb9t5s1AQqsn5OkFM1P4
tqL5L7/D5KZ8Oqp/8YVAXXV3nHg6gKr/D/M3JDa4LD1W2Vb6F38t1ZtvWqoi
xSr8IsVe5k40fuosUcUYcTIoGd+JU/ylToCA/hw/L0jld6WhurPJZBPA5BF+
OGK6lAhH5c5xFbdSXnKgbfqmOkLhm/PJLlUg7tTSeD8obrXj6bmxRjwBu59a
3cqNtzv8fSd+lhamdBHaM1jS+1O0oxWpgJZTzRigRi/qGKf/68XpecaUJJoM
TFNOfMsN3CDyuDTQuwJMGzrOpHtHEuY/2dEAHKYbuDguq54HuVHOsJ7SmPi3
A51U1wwswK/hbk+Js+Q1HLJu5ypA4S9eb/UdkpRTuLyEsna6p5InlhjtimCI
mULAoyrj3qDr10iv0FnnLkw6HwGsaAQTcwMcgS8+hJWTRosjurhdUitMzxRW
0+5vqlzjDQL2shT2CIK8QPhGfXkG8EZDAfY+ScaLIXt+T7yupGm5PLajt0UK
U995rH471pVWnvjKRW3YJRbZceK15MA89AiXJ3sGXnti6MJWnLyN1UXVFU6H
Ig6ZmoPwC6eUQmrOE2YqWY3/gTnMXeqltak05yujCCzpPOkfB7lvInT3yJaG
ucVXztn8HRBynDGDxBuMpdnjj8+3iUhWDBLTG0KpyEl2SnI3KyWdndy9cKxc
f9vFw768uye2BFXOvPO+zf/h5vAxNI24EwpZc917l4eW3Wyer6+NPL4eC6Dp
6SPSRJgbatMv5gzdv6jePedojgjMxnexwlEqe+xaCwa3Wvex8zyHlYLzEkus
4PsG5TesgmWDYL33l3AH/3GKnIiylHhsmaomf9tYEHvm6QdwOcpAHehh9vmO
tPKrL0TTu5f+fCOql9fo9wQ7pDp6nFfIHexOq0AsblQo66gp/5+DWdi7Ou/8
fSwA8gs5FrltJeGcMWSoOCI4yAYicGMq2Vu6ZYUWHhgT/aGimaZHtJfuxQ6z
Ua8ySIUvOpP7eVNHbuJXiaZQprOXIEvix+yo9GI2zLRBgarT7zBPTlpS7wyF
JJSbGot4M1EGp8LK2PMyLLXLYrqSzQ3MDrJ4lLgWAB4jlZBF8odxbQrvEB+B
2/U6x4Fihd5AC36GHQUj/G8KdOOzUgNjVFDPm4XRsjEtz37dCGW4fJJ9WvcC
1f/VLew9sy3xmhnaGUMOPtWGB+P0sUgOH63gmk18M1gDnvG94W5iNf+Xt1fZ
JYiD3PlxFk8X5vC46oQ0c3vRMhO19LQvtOz6Tf2MZfRmuzSvbMk+pqmRQDpj
Z+kxdb7x/0Y8DKn4YHKlKLcvOUXN4Z21BcX9X0NAUtQqxB644oBesPDsF1UD
M3Kd4e2A1kgmQA52EMuVv5ISRjDSJIiKdVbiCTYjJw5xY1oRph6Clq2sZ8ry
Vd21/SRj8tqvreT9787t/Gbj3eyvuTJi72VVsLb6TRPvwnOHZcRf5vuMpA+z
nEQipJKd190lRsnZ6CgnLN8BNBKuBOP1OY+VAU6pCBRKIjU5oOD+YPf0uLev
tJW3aGr2tWhIP4t4Z2yq9EjrPQcLqVFZbpOXJmGVvmiPwWfkFlCHoeGyxJSC
SFIX957AdfS539sC650QX95I5UtI21q7/iZcTWkbe55PTYn777mDYynsBpeV
jkJXkhMc5FzrF42LloRytPy76G6bi4BXLvE8vZyZVTfYZa2PiM9rlIXfr7rL
n6Ij0LBsBhZGdhf792PPCmWjnbocVH1mS9M1DPuUUZDtsaKFBAcbOKlcOmvX
0lec3b6qwbh4Tg0DZ4mju+QjDSqpfZRyqN4lrMdCZzJvCJpZNaCRtxiTvFMg
i0qoAInI78WfbOdwtfJVecS0aDUC2X12KGblj9uRUGb5AoVx0RNPh5o2Ukku
0eH9lXwr8uWsc39r6ORFws80IEsQhmaKUj7ACkZFjAb8UtV+XXj/BK9Al8DK
20IesfIdvAjnP5XnwACkudOOIIRsH6PxckczNHZi1/UfmxLXXUoynqzm0DYt
aSZnL7wP1cedNbJ763VDjUqSMEZUB7aFNptTX+8vrkHXpshSjR/TWprO/ffF
lkAJFjKcD9CFD9JZKdPC8nHIqFQO5l6mNG5ZLjMFsXH8s+XxwSapcLRt0xGd
YZnags9oYGlbf/M+7gGfOohNn5NCdvwm4ez2/PbxZqXb/tZJ5+YKIsARKW//
ae8/5TO4JUyO296NDvjuTe71KqnL5LBqke/3pprTShe7RSHFtQ4Xo14dcZ0G
LNDdpERSz53rFC430Ar4Jpy6I7WIvS3xVWIysjtYOz06LpsSwtMJSh1cZqkW
LWBM+H6DydIRv/gBcTb5Dx9dbwUPAFOIxtLw6QSpUTVoBmrxMLGPoRY2ibGf
3Bk0GeWL4jaU9x1fJr+GVKePBPE5EtcrdCkbV7kBuL+0QtEL/8k2je1uuYmd
UfjcEChFC0BG6s1omPcDGDzEqqELdawbAIGWjHzd2p6zmAj7XsM+mZrDxFc0
mW/vZd7f6IsPuedTNyHEYGg6TygG0u5fwJY7WqPoy+rrQyBTiSHOHABs8ZVb
wj9XMXmE2yBe0bLYOduK+If2g7CKjXiNNhvUkdBqwc+Jm/AHNyJ48LG8w4rM
7EPloN8QbvVZiiyAW4uKrYWdc2GGHLCeB5uvWtiCcuLdvNdIUi0LLJz+fqDq
y6/+UdaPiZAK6DMmOWB98dY4i+5YVudu1iKKBiGmv22+KLOnWAzfsqaRjgHK
gPfc2OtlqgZuZ1AZIGyjbiiyR7VQH3gdTqztLPv2t1FnPf+cNBbdVTzPub2Y
RM5Ev6CZXZX3GyrbtXgVIRqql1Y8sBeWYTpd4QAdHeT6YJ+yzONYSjv46t4N
SD4tDLvDxMAA6X7wZ2gjNdgQn1Vi4FDZc0axwwRnDklkzLVLDsCL6P1SywN2
D8jaWrETR3fJjmB0ZFtGUaVFgt0c9Ra+fWnTvu56QtbyeeGqvufNEj6SZkvn
Z1EQnEYorTowFE4f9JFhZ+rgjN6BABL3fS+8FfvMl8TTtttjLPN4S3cM+R07
epc+7dhDi27bIaUVQ3xS1Ai1fKS0igSQF9IE8zM7ShxFUjhNkP6+5O8fh1OW
CRQvKHUfVsnpxF1lUt/uTC6/ykTuYObB+erYpd2zAsL9EsnyQ/OhFtVk5Us9
h0eCO5h2Px6e2ra8l8WLOSL7txiZQTjY5LIQkkoBvOSqjcpqqfbc8o+AINZq
THMm70CDtPaLr0NVQPbs9FTe5I1LlHo6JZpsOjFiZVI0WFoG4foVu3ym9P7L
h9dRz6I8zCtECtrViMDYVw28zYnsFHSSFI0hmud/o39TZCuOK7qh/wTz2sVe
p1BSxEjNIBV+Pj+qs+gdDXQwdZsyWdLsgJIV4OHQny0v8FhL4OjRzbG+50n2
slI6sM+dFF+oECBMQzdJAyvYM/MLDlqxrd2XpKHpbZKIVexW7j4X7WyIEoBC
crkxWXQfieYGVHtqr0QIUVK6L2de3zXaI0frsqVHuyxJGWs3c0tRrx4/f+L8
nC41HgImfE4r2uiCPHqe6J5yRloeJkFX0B6LMiTgpGonaYb1+y8aJdRYoCEu
/R8EIaLaClQaICUvWQ4pWHISoMVUq0tp/7Q+5UIj/jZSQGepdxkq7qbwn/zV
RcM8eBBb3KoGnslWLerfPrAX42BQQmHoJHrB5E2rfOiKPUi9Z2td6UuCLYpc
UqlcOvaPyNlbcJUGQ4waRCeetLGyf3UAusOw1lpzBEqjNvwnX0jSwieHfeEP
a5gSrevXtcye781KOPdOk71mC4XmvBJdr1P7M12c2ew+22fvP5Q/ghUKdrPK
oDEzzzajWusQg6wVSCfBv53vN931l0LGWtYjYBUakbT0mW9hP7UvOkDcIJXR
A+IWDDUcMZ5zjx275p50mtbLsrzM+z2X5NP6Uy1B+KNEQrMTp9koXHsDNcv/
gs+/VvF5E2QnvdgLEzVOneATSps3L1QVjJ/ujZANFdEjClVVoQ/s66gOxE2a
XpGlHwx7uxRo/qSDg6ZSJuZmEQ2kgz6dTtVunVy0cS3GW53qdF4O55KewbbN
j6QrH+4nEnmpFGIljH0PYsTDKpz4IkH9hAs7RIlwivlgP0qnZuCWoU1XVBpy
pGgUvCWJ6/5bfdM4uEo1drEzmzEBDcHrq+h12WAsUyv5cnJ5uTMXO9/KfjuC
TDiNHtJZlkdfaO5RBkAOuKVcFxdYB0JgP9lFEs2rmrXywhfaWN1y/sKBEgOT
NhZz4C95mcrveRJ8TY+J2+9nZnBrAnZbROa5yacGGO1goOacuEeVAOZIuFtk
kt7rPKzCdchqomGC69uFzmuwzOuxqppdZcXGofBcZpQlhDEFu9dxG69J05fk
xUOe06SOKeqEDyE86eu4ZHj/uwqrk86+0AXjVS+YTj/X221krf4VsSLgsOIL
5ifNpHOoZXwITXmhN221XewMbHoIZeHPX7pTnuM2EqJDzFKWvxF2td0/u6gB
+y0H5ONry0FqybFSjZqlwqxRt2N129mu/vA/IMQcpBLBTUCFPq0X16QRa2qD
KiO7QUOJfzNafOOeYog2ZAf2amloRmog8VwXu1/M7vityu9Q7U3fPJdsvcoW
ng41BGQZDD0mHJD5tENvKqw3/KzeDPKvE79pcmsWL9sSHW+FtTPmTL7rfhhx
VlglACUfqN1M+BQZXwvd6JzeZC9kqtcReLP7s47c9EXZ33GwTw6g6VQ4SQes
7rTLMtx47j2hi4jnMEi1TFV8ItdufH6aLVC+YhbatntQcpf0uEX7YPSEsRKx
I78KmuIx5DaHuIA2tD8Xb0iOApYikyP09UHFZOiyx8LRx2mRcAUlKM0Umfr1
uHIhp7Jw0f0jD43Pl+ic3WrKkPyxyFDLGFydZoAo4qq150fNB/mfiJX1y8kj
TA93lfj3smXewNCGdLn5o+iVsKt5A9hUH3gabGUb5z7ufJgoafaOjnZzAtvo
wgHxActng0qNaH5NxWsXB8G9LtP085dOSyLz9PgWJd4jsha7IchDVXBdLvsF
qpkuNaaZDQUEqX6ZU5quKhi67JNFqOgbFK+YzXPqqpL2RvJmSDmkNNU+BhAK
kXmK06bA75nsA6/05DPxiX1dipo0rm1+jIIymEJpiRa8UuQHwcqYlcvKV27h
lv29ikJmcGntwf47d+clH/RIvQjzhRbZW112tIA+///i9SxQkn4348pKUQYW
03mECDx/yNSWKeybLlzti/dS22jTflmGhRE0Bx3WQfNtDkPNz5nARJtsJcly
DtYGVUpTDTA15lN0g04t7zR8xjLMRF9CBC6qEEqt0rnEOMAx+QXRPfDiaj/Y
8wty9P9iPxuBh19HqlTZzDOxwbJeRKE3o8rchooq3MIWoCXUkxve4LV74xjj
/b+CTGxIO2wtY/ivvUR/e6rJQe0/CGSDAOdU9cCA6o/d3Vj/PeJGnsLVKWgV
C0ZypFrdjPPK+adPDJwrR/Dey3S8t4DPo4cfFu6xr+5U7e8b/j1y2/qHr3fL
eiRrWjAfErF3LjADACGVC7VtzC3v91pzS4B+WjC8BlJcz2vtZz/bobwGTjcf
wKcTvDpmcoS13aU7VRQkE7sP+YZHZj+Q7XuMOSOk0bxrC4piebE7wLuPYwCt
lsEdPTcVgPgA2YR4do1duCMvoeUBJxoOvRUxwrhbFlwT0gA2AQqk/A0cLjZu
O+WCMnUN7hKSe06YgioLcGsYDaIyrq7Cdg5Pkeq3zw39AKYmWR6qIeo3d+9f
+j7OetZMejqOVuma04a/cV8jUe1Aj/G/TsaAp8sKIh3SIQ7yGVMPVGKFzj1E
B6gisJNj4oKTT+R7OlFJPovstvKmUqbnuwgf0wcQUx5DIDhIAJ44vOmmib+J
hqijbKjMFQ6q+ssWkzoWE4xqFhgHjf8kqIreiahAhrTh15ph02QkD894FzPr
0vDb8Sl07PhWFHUQ0JJpe+9/BEmjWONSvkQSKr8oHNPxp/LS608KEUsl8HmB
arrhmU5PihxPMXfGN2gsHqxjLrmIqVgFcNcICtH1zwb02YLJmC58qfiEBoVe
+azhVD3W1zqBJpGUDJW0oC6ZVWZez173cqFCl7JRorp8quzJMJQ2LCAhBOel
buOxHen7WPk53ApoMz3p+UZ5k6okH5yz94pm0SynrFSkqLDWrJjoHsXAZYIg
3xzAxnnFaX3WNJS24gUrwD21kckcQ/WaKXnToJj/5qU5PpxkVOKN/Crtdp+z
kJrt3ib0XIrreHCWvwVlAl8wLvPWh+Ng1sGb9IiEIbRM+GMT6Tz5n54Zza2Z
IxHgJw02pCtTYhCJ0AvJNHg11wjn5Yxv2rNRVEh2yjT59uyJq1nvnZzhJsOi
W9DiyOi+/ZM5C16Pp7bZG6GEikc3KTM3V8X99qDzfEohxLdlY4O+0kX8Rji2
ULH8DDqq+0sz1IWyefTK1hdh4BECZNEBA4/DPiBeUtMgbPTzljk1QBrlrf3w
BjnQmiYQbhWjfIyhr3DLG5QUgpgJ/RZ7HTikI4s1ch4zlwtNI9JEQAx8uOqx
p1kqrqLEan0AbvDrLXyUip3lWAgribFRHGaVt+UDS6EePXEc+kFDZLIHPxEg
74JXt4+pKGTejqFcj0AmFluoPqf9684I4fdReIV26FSHsQOFj9HXNPAjyE89
5n8pubc1Tru2WVeHqnkBDZQLKBSZ5/4dwWpJ5I6SKSb35TQDVyomK2TiofR3
wgRALt49Gd6rEfkSjkuXcc07qOBf+6BBw4UroFMDXb0GdiL3whv38NdJliTS
zgQB4685fT+2xzwxDRfOFm+7EHRoC3FyxF0qcxsWtFpnqxIje+xLEbrtaSxJ
IzdIIqWKF35v/dJNub/gzp5jUPQtI8WzhDndEUhD6rmlROZ4D0F0pMxV/WVZ
gSy79qPY7Acl7uYiNP6RiApEk+LNMSnpUP/s4pIe9DUjk4vAsdil6pz8F4nw
cJlLIAVOzySjIQs9G1x/2XRwlT7uCLTJ61aDk34+DL0B/itHfmTccoZ5vRht
QhInN6SfIGOCMDxArqzDZb111GVx2N9CooGzvigA7m9OVhlKXKFMJB/ePOCy
plyaLSM6N6i0j4RVTdotpudhtcHqaQqI/Q16o/x8p3BaINm5wTCAg2FoXDGy
8HiAEVR5CjFvioMzU6kRKlQt5r1IiLMu9OcmobTn5C0BVLY9PSKFxyN8vgwH
YDEd7BLR4WQGrms8iB2GLSsqrBZ6AzuVB72rX2r3JMOcNF4ULfIJa6KHyiBr
ztsxocbupFhuRciTDUiF2Oh5HliR2FiYjR33yiJhxNlA2ZrONMv2Hn/BBnyG
Vcb9+UmILMaXsSG5C2zalBRGpwFlEGyhQuVr7JqrjctE2f+f6ieLBcefS3rt
3e6a94oYQ845lxkDixkZ9mgr0FAmNs/Ei6mL/ezPLekUmWxASKwfhPr64ve1
+Kk1bEF2DgQMz5R1MFcWCBow762UlEvtHUrD7OzLlDAuRZmH+iofSXko23zF
abME/tRw0eULJtGtOaLl+XsxuJFgtkHPVPgmgRAfz+hFUbeVJjn8grJsagnq
9fito6Q74PzGwn4ZK4STlNcFDCsX09pbDJYTyjNRcx1FyKRmyQB4XrGaTEjo
OoHrDto5vsWyVlf2MGwGza1F/Xac3nTwKra00DGgv/Du+++CS4rGg4Gz4rqJ
upr1Sp9P19dJ6M7Xf4NFkvt2axbbzWz5nt/ilobVV3JRcOeGY81PIE+uXYop
wYIrEoqK7fk4FA0zC/uG30KIrVyvuqgoZl5cN8u3QVhRZDWXjlwpEF1pQ54p
aWppSguYc8GdDWAyOKHM4X7MOsRyxsSBgDehk5urkFwUXNem+PNmoAOFfMtr
34l5UYtcoZCLg/LWiL+Y9+dMvm71qYwU/EkhiVMANK+fltQZoIJo9BpThuc+
+vOYB98IChPIGd4nXCv+9APwVuwDbbK/ALyWE9ral0HMKu0Pad7FTdFz6ciI
5xVGTa/BVS1+8r0KFs+3jwif0QmvY2k0QcYE148bZa5YoGc/aCOU/sbaGp0C
5MsONrjaD5nwdrL4y8sdcVpkqbr+TfkZvuxmuA6yn5IvL7rK5zNNTTEYHkig
1Th7MvIQ4vjhgJk1QjmbAjTpKFC69xE0ZSB39OvrqbMOOWUZgro0Eczfc4DJ
ZCcyBebq7OVJNGwRwdp+Q6P48Z4g3PELkZZm6AkTI9lr1VDkM3L3cbPIuWHA
juCphWPSKFYsC0VJaMHR5cE97xYfQDU5viEl0vsofX2HmaFtzlJGmEmnfwZS
vadTCUUnN0BlUCChmrTA0Z0TPjTvjgq0ZvfAyWPErfvdRN0JCdsSorxgAplD
YYzeQxCHP6Vuy/6JZUGMepERTqTQ1/hi6f94K4doELuiuJq3Izs5GRW3apSE
c9/hGXvRPJEJ8eVJDgkyLgF8XzvSQuu86JXQ8Uz8ER1LGz+eNUfjhz5/5swK
J5eG5WOTOSoYvLF/08fHet41Kmvh4pmOQzXz66Jdb/om8+UDlA3ACSwSPoO6
cUfoL466KCiNGNp1uOlW7QR25h62eSh709ZIcJeaGTqqACRYkevPNKK1C0zf
oGWurzA6pBqiClrEKtv/84PlswhlGY4JAPNjofm/vOYTvfqEJFWylbbBpsmZ
VqtR1R+vG3jjy6HlojPOw+tMFlYKOOeT8PKkEhnWFUjvVCXO77I0aSh4rhzo
jveXLMiZHzYV15h3E5tnxTEEf+5pGQmnO77gHj2w1XWBAnfMsuutlL9wZ3kx
uPAUrM6m8HAHi2lLXEVzMmkOLL61yJ0yZKkKTLk4S2aG3tG52m9l8RlvkruL
aEIT8t3eOUqS4aOdhljj8uPJrf/reSYqaZ4DB81Z34/PivAGT2nrow89B4Nw
AsUT8C+jap+vu/t0jefdWdp4QLt4FXUaZaVnsKoyOIR4Yl7ModiyxfJWMwnh
C0DiGDNxBczfYeOt8IcorRkm0/25vfeqVLLPlOCYg9Qek/d5qIGOgxgWMW+u
YbUh3Yp/kGGfxKHVb0FTvDVlVkN2MFMnoc6S+b7o4Ye0BQZ1EZkiSeEOaUba
E5AOQdg4Lwa/XXe3tWLgAAI9yk10IdrwI6CkOyXVSol2DllWszBVLmpHC8Vy
44Y33YSlrJxPj7q6U5aY2eCd70V2JSZXEo7UaRZhcuZ2XORw7qepZFyT65iC
Vl6I7sPCEsCV4sBRfo4/VIGXkPFC1clWkFSyRwVM4tXJ3gdbhbfhWYpORvst
dcd5FrG5ji9q13i4PI7BkD44ypiVUyNBZF7Ek1PVTm13KP4DnoVPokj5lrw9
XdYXzjxUAlZEX9rujGW4r4iycarBDeSHpGOJR81qnbATHMrpLAewhk6EnX+F
6rIjOsgC7uIdLJ0tS7FPLUGHOwn6vOrzRjm4fByvk18f4pGXxKminHF3sFPP
H4wfpbwdOWkRWv72P7AqRTAfIuAyoH8jrCbQVGCJs9U3G7/+tNBGnAdX72Dx
cMHXMfCEskzA1dl9G4xGtmbuqWGzf49hO+Zvg9Bltmyodeim2K22vk0auxt0
jEfIHRg3AvLUcL0esx52iRKIxjEfaZ/2jnri8Z8DeKPLZn3rjkJSSIwrNZEy
/NFI2DMpVDM8ZlXsqGbu7fBqI/5SfzCGkuf0IOyjYz4BT+fqEQfBjSLPV/LH
z7hyzYwQsXF8klORVMXMEcW/w4qAOaBaHc+/nA6HwrBBqUVD9WjH+QVnLsJC
1PbWO/v/L2U9juVI6kMvkN5PGw/hhynMklfz2vd+4p1RQYkYtXCmOmSoLrRn
CkARqOTnLHZpsGglOEf3Sr+5/irUX4KOX0x020X5xvKX/isJUx1yH6nw9nmL
t31PpfCfluwTbR9X1+ZeovYFgzs4TR/K4PUvgzlzv1cIE9O1QDnGFv9mqOBA
1J4rnNJzkI6pSqXJPSCM9aZNGfrRkHAavS8QfiqHh8kwy7eREp9+6k8P5Vs5
UhwPdRdrQjPFNkn13wl5MEdOeJiHBOwYUjWjj0Mwfp4PV1w5SeO2UkbWU7Xi
7nLrS0wFeJkIjmDf4IIGOf7vBSZSeEp5avtbDECwb2l/Xf7hihhb6cf7L1Ns
Hay9e7lY0EKzuVgQz97goS5VWwOMuYxXjOOlTUaAOWbFt8JZ7+Bpyhurr8ah
99J4/4mOvaPrCMPmgfwyS3X2kXdSvYfbYSYpApr/hQ8LkozuX4giXZUeBlxu
DwKfIvnWz6O9Ckv6qOaan3yzrLuaAkwYEzz0PzjMTNTma+jv1p5faVly/Hw7
VeJgadAsulNUOp4bA+WlL3/AdW+dUcSjNd8p8ezSHe1tEvaIzeN2/SIWzptR
ztH1+rFc419f9jg2HDK6dNvxq35tXZneuPuwVWsgSkgiBTJv5a2nRfdolTek
UVhsPWwbluJUQ226J+Z8ySZY7/ffLnI5G2Wp/TZutf/LlCDcGJ7gs8kDZM2O
DeG3ZeBO/LijUxmdPU7AiMf9y51kzonVAQvplKcwBi/EoMikpOK0VqwXzP/M
VYthTXJ//G1Fy4wsIcM05GojBQ+TNpNUpFNnSz5hyHOuzjKCz5VPehJewgsa
vwy/Dz8pWtmvffraMVVBPW+8nOdKKCgqCxgMk5C0wJJt+Y0UodCsj73YTYo8
tSu+t8hrnnHeWA5W/o5/M9WCli/m8319wtd3FFF/NGYz5KJs30dU4O+0SIhB
GY+ukPFznRXNN2cW1hY9VRCguOXUTgC0xcSAGfaqRB6FKQ7bVBnAsWikvL8L
yOfaymErJlniKc2Cp47x2a/7upmNlheozXnONDgtDSM4rrtzaXjHX73TBP3v
SuBsutdp+z250TsBVsS6VMBMikhm7j6gMtxsUp7KNeU6mDySiGpfguwHzvvH
cKcmhirBZ84LfG2W3m59OONkAWdqKgc5wufGTHp8C/LWRQmS9oPUYPKmRgUR
Dg5y3zDhkaawFcWtdCQO1xQRJStaZ5W3MZXT+V9D7MtBTC4tUgo63UnS0C4t
U9uIhajOAfUM9cXf3kodTr/QQTHTscU6pOm3EnSmJZ4sXUIXpF9cezTQvNpa
F9Elt0bBDQt8DAqZGwufjrL6SFfe8Qcb2BJyP30WT+d68ha0Lx7M4GxJjNYX
0/4DeKMVq6MRRA/7TzzctiUq+6LNz0Up+rJTfF/U2OBAPZp0AehzrfIS4yQr
VS+TDcKi5FE4I+jTWwpaXysqI5+auujBSJXss83K+qQX1tR/XSpmDLiMhj7+
Z8UVHjk3CgGThThib8QAxH5Sv2KQ7etxDPiLWpNE9PWB9mg3Mgs5R7/pcJOr
7pyxoeBrnHRV5Wa5W8i5D9g/dmFUyrxdTrk62q5KpiL2bj+TC0fUh0PVacCj
LkKP9mPuiJViz0oeZ+SKFYWXqUvSyylJ5minNmNqR7HG6nGXFjQUmvveABb3
EYPi7Iig6GB6zt/5+p8JYOU/TfrAAulanEENge+0GVf0QM0rR8V55qSAu+9z
3nDuRD0+XEdz4A3c08vk3oCr5iksvv7AiHfBw91mdGROjWyMeWOgTM7/xJlf
VzOS5a28GOQDIzkMfYv1fc2CKGAEK/yCpdmGNE8SOI4KruS8bKemO+Jv1Fml
jNkReGOS85zR4/ioahC2dkxzj2m1OCmfP/xxDyl06JuT3oSn/Yf9ovlcQvg2
KIbeew28sB6hf5HYvfDqF3TVdDJh3aqa1/fW9vMOn0DubskvX/qa/OO9DPdy
zuKTJxmL2h1EMcjvk2wynMRWu+huXbQeMTOEoiH1BAoKhvkA54LbDanWEI8z
wcjVXtSajH8uFJKGBcE29/VMsSPQ7d1dEoy7XH8TzD/6OveV6u1Aac8iwi74
9R/X3T38ijDpPvJMaTVecAaEy6lEuU2F+NwagvzybF9lg+6aNZXSVsC3+Pb5
jib2YUrsWniFN5xELBT4Ox7ten/XV4xab6mW6WOMA/bSMoqaNLrtnA/RKotu
g0fKGq9KN5gMvg4dFlHmzdZxmVZkbuHG/1vk2I/vfB9u++LUVtYF3PBi/3g4
nyrX8gmS42sV4d5n6p0dZ5QRNVbG2gFGtSVzWICh5IoRNWNvQTgN+PSZQFk0
/VxwXJTBgo/jWRuEt9+7GHWwz64PQDK1kaL/ZVNFxI/AiF8KjCYe42lVlePD
wTPtLwIkw3zhOcdGPh1MbC1UeHlNkBVMmLuZRkbbg19H0Z6kBMUSbXh4SzB8
TJ+o6DKXXdfGahjI7q+WzTorIiLQjt/3GpRxTrKhTsfZF9sxiILrnZ9HsV7b
+hysM1ClyVe2KVfM5NMxwMRlRn0p8qjzUGILTnOW9FiEi3/AepZuPoXlLo70
pO5dfWhtupJsy5b+G4OtpHuMc9WpGjeL4SbmieOYlDwm3br6IaekcN+zhQHz
4FwZrLjCuf7i3sxOu9Kb+Vsym2OE9cwsDpTkmiu1wabiOJtdY79kenYplJVt
kb1Z/3IbXBbGuUjzcdS5nrS9AUC35tkcChfTe6MZXyeEhNODi+SOv7wy8itV
2L4NDFvjNyrRmNy1eNu28GDQkGxQ2FOq8oyABiZfj92SJl0CpMmDwfebStrB
jeL87HW/pZF34T9XjPZ7CBIuT0YINnZ8IgRb6qlEglcPPHR2f+b5ztmTbrC1
DsY58gHRnHFre/NaBjeZ3JWNE27w/5gaXmPdpn1G6avDi2O2tjXWnIWKugU9
Y0qvk9nVawXtDOm7Uobr+wGpHVRpl/esDrxuDwBsDiiO6jpI6G2Zbgj1ksGc
9LjDyswUtUX/wjmYPl9RfvDjMws4isOMnLFpOxfyDDiiEZGYTahJFZjo9eCu
6bOxfXbGVYZg270T0f+a9E98n12qfb5FY/wbXSgmlYBONzPPv7/sfJa2qGNB
rJT7VGpbXsii6F7ktI/z8kPBqXLrbOKj7JlYBZfC975MvqwI6+moct6AxueJ
oqm1nzOiQFevzaccoQtg/akzPIkPULzWBjnM0p54TVHOQLuVMXGee9wDfSzb
miUadeKyVmomTf6rM64QHLG7oeNuMJGN+9vgibv4oRbMFxxABuBIEuzuJl+p
k9DhpBjciTaA/bmevV0uPvDXOG4/55NPy1KK3pQyu5uai2E/Ah+3xNaRqkce
xFX5VZ0rmmZa948rVyvHypnu61nid0qczUZF4F789bh/YyiZTE2E95dkllkF
gmZ3KW7uZ99jKYlL8S2fKEpe7rHHrz9Ht4P8Ki0m51oPNcuL50YYwN6EJ+Dd
m+R4HOZX4M56/Tl+LF0sSBiIbLZyph0R6IMlJE6tuL5nmWiixcAG2CgWDCRb
z+HATb8AMGEOc5YKDfcTorjE60iymFPhlX/YMggY9YOhwnXPfQd7R7qkVoM6
oo37V7kbVsp1cpl6EgpwfZioQo5opLdNKQG35jQChFBsHUb8eTzspOi5mn5I
N1wpoNQ28ud7hTOsC6I8K4//AxxwOW6fOv2VWZNrN5NeAP/wFQiSoCexmONs
haW/wgAxG5WkFIqMefA8Z8OJtOEfk3I2ZS65xnVyJ3LNKHprVrB3e/0KwtY0
qjIUOk/V70R8z86U/TxaQtlZJ1lRUKgjvMlCVkDxqjAPi5F/WMXCEsaXJWtz
+kVKBQ3284/EUtFHfHlEMoU31FfbJHKUTCVYOiaVrJorfuogHDYpCcCLZ5nP
MjJStbssnvigVdMCYz1d4a08DZBQxfeomrIbmT71l6ojhW6JN7colZg99ETa
c+8nHQyMOWvRqjgmHZZ3PWFwcl3H3rV4doL+fNJQthGLGGmokBSJvUbnz0os
g8gMb85JUXos3+jTXZHnM4938dmC8HtbVos8GA78EB1VTC0cnHhZXPwNWUfA
KGEQEqD+Hp1E34hd/faUju6yvotxHgmeVsVKTm7Ylq0j9WBPZt+xDqcJJW2o
Xd+NondFM1Qg0YOwGeaX+Q7FOSyhnUh2/nUv0IcQn0OgFPU727HKZSe+uUZ2
NPWTxKTIwoftZkBbyUB1BxAc8TO5uY9N9LJopKPyVmgeZmq26cKf3q51UGpc
SjhELP+J5stK6gWPiu1nATr7UAsrXde9R3BZqNvKbr++sPHcOK3e9R1WOg5R
Gv0KM52qGgCzDfelhvLwRw5F7W/QMXyPYlvUYAEz8oCuPtMCy+2FaA3MSvbV
8SW9+yQHbnqj7CWnEhyy8Lilgh44a2JWC7oDrFIzjL43j/rZoOlduTH9oKQV
i+OCQwVPfEfdqsCsvLzl1Z04OnEC2ZnCSCOJuF1D3790FK4LXz1r6xwLagWz
an/fHN8Wc/twWSMlTu7zVUM+1aI6abPtwHdFPZvH5j3nULEleK47ckV2IfSh
/TOU12BsxO/bCwQt11V3FZ8vlcUalaNmoyTkkvrZOqGtRqqdnLxWYS5ozwue
+l6x8kgUNxqQ36odkywgHGz8bLruYyY3mjQeKrWtR3Qj1xFgy/DWPISP9gsP
URJcQsIKQl5T9nt8W3YYQRDwp/6LGA6labLwqEusin1aT5gWuQlj2xDsf7K0
hqOkHhOFtQgzLVmcVx8QiVtePH6zr7a1xLqIfwjuagLPbmzRBl4at7mixpQV
hQMih6fh0ywjoR1MbwiOtzKQ0jhqj44jWhX3SOuZf1qd67cSKjPLzBegEpvc
Zp2FRK94+MsYz0wWF0Q+UT2YPuxAr/zaL2Sase7ljTFQFwdrGBihPT+1F+51
2ybMfiKlakMJhn3v9slkTCPwrRBYWsK8tZ3Z+0sGuKdYjUVM2YpU6ms1HLMd
kYHodoeX/yL0hYUF9eMqxgt6sLJz/XjUX+K3NCsnO3JiptkNvF7Tq/zac+/6
nMpcCxmg6hE/Nmu2v9ByImXScRFWvOYmgk9b1DlOiBwxPoBtIgYreW+bjR0f
k9xTqA1qe/kknBcokoRtkEkzk/fsgwf/xPH2vtFd/2858YeDBFeOUpd2MMc5
arAg8l6P97eARjvCZqX4uU26iB2NNj6ImGjAcbile+qccUCjA0ZTYMzZWmuh
VijlwnIuJo9VKMc6uI8Ejaxnm9wg7EnjMXyxujUDyAlvKjwvSEApM4v2nfRi
tae8I0zkQ3L5nPbu6udwRAMA4WaX262C9dVfX9rkrzx1occAneCoMTzpItPd
HTTq5nZ8VvFDzdEw9G1ZmG2drh6CskWIL734FmhtunyLxuASJ8adEUAMkZGX
KzgpTKI4zHoRgeI+zA1kwHuNQG1e19LJYt0y/TKKPNQuPwXCHbEGNk1H6pR+
sDHIZfr2En1rINt7gPRMudjSjxxIhrwYDlNAlwhP3LVpAc3sWzedbs0+7mNl
yaCS75BuvYau+diGTZrNMyjmBrQmBemCLBGMSDy0fnPucXiaWpVNXsgZ1Pr5
IJNRmzk6syVmf1OeQg9he4Ep+hcH/xeCjeWIRyVx+yAfbCYgaOTYoxQb9di2
8W97Vd/AC/HHlbJoO3Q4gIRL+U+PPXSbhKp9tqfmOAVlficNDODa6ctvBD7e
ivLZ7FXq5RsXLFD2QRAkXjqRO0sHpqv+W64GdwqH2p0u/w14Z6RZYH+cS4aM
CXJz1eNzK0J8JHjUct9VM41Ta5oWJIosSQE1UvXjfH7ZLq/qJOqLzYhTz3UF
RCaHpgYNJK14XV+vZKsjvuFT0Di3/m3lbj5F8GVH60nu4dWcaY5IAq+StzDr
qVQXpme9XUEsKCs2in1xOrff5lkvbYNqGRWr99dHLAo9iV9hunTxoNe+R/h4
cXQDoSd9v4cVhqAO2w78eXBVGTbWXd2JqnpGA3gK7PCXd6dUIui/afJvn79o
Vrr4XAPVcEhKNHcBC7le6wh7blpn1kM06Ehq6aKFh7quzy3TZOSfe0Vu+Twn
E4WNb9fmlNiDXTjrcmGuJUw7eNN6iXFJ5Zj3RiVD9K2iAOe1wNliJgVbse3a
OMutBK7z3op6dA7IS7nvXztA1bOOrLcxhNF9JHFde6bJ3VDFFqrroulyjKYo
ayX4JC3ZNa6JI6EFqOP0UyKYYtb55uyUx3L7XdnagTREh//6GnelFAdsfzid
pbxWFuzNZ1l2ZC4QMc219p0W0WD7EgGG2B7gv9eBYf3eX0NXHwreh1CiBGca
WZHM2Z3anVPosF+Dd6RjgoecCe17lnvYFJh3eCIrAa5Fu4gRz3FwI6LByQEa
G0LTxrVdPguwFlrbEvYlU0CWq1c+jRqGCXE4jrUjYvJyMCG67gURvYtlzSkL
pKBs6BPUc+bqFSExUaLBjMLOK2quR4RJIzk2gH4ZVmYP9mNZfwWt4y5Sv5gT
87WzRxPDtVb41SVEEGR509wYEuC7ZmK2QaeC3pIJ0ON2o6rW8nQ3B19Ghrnd
UWTK0KGY/LU6d1tUidRdpq5X9VfdH+5eNKQhQ10V2NTs1lFChuUkuqj9bHCZ
ivN9G8qb57YmJ6vJGd9vxAT1Ybm5FwFGxV338LuWBw/RJXKZ2gQTXykpoAWm
2mFHOGYW1Hf83zdsosgm8Mv4FBuPJv82AAwS29HHbHrAs6LLWoUps4eVnd9D
1HN+CUq8+GtrMdyceWtRehPnOq+c/4aWLvycMTw5rzap+FVg15KS7SW8SDqm
GIE1DpDx3bp5n6W6DD4zsvQLdOlQNy6v/wDbphednZ0poVLvx3Y7A8fMQd7H
8tYFZTJC4pLPLoW2//uj/mpsTLyi3jv1T6vyGHZJgBZsrm/UA4gRUDe+5Tm8
NtemG4ZRDHLwW2/4ws1YaYDy4JchtwkCGZNK1nLBwnneKSRsg/LICgfLk0pd
kaJ8P1PVn7Rr0t2WmxEmSIlJ/obNCVoXrDEiuSYKx7aQ6kIB8xHkvkvrYy32
yW8VSxUwhI8qcY5qVCRWcW114+cSQXE5uCNDJxiiK0qSiAZ1aCcTHQ6Jlme9
Q7QggBjsTh3TCJADl7impWnZY+bxx8eqJTAvmNqhIyxq/y6WvEpTLh3WyDYq
WpHTQs+F5wD2F7uxY0R0KDcYsy2fWpqJpZixQVeLYr3PJMnE/HrDmLxJODXS
YnNuIlSH2R3UJaMUK9ILzTisynuaI7GVGQaQ41EYqpCXQBQGfc1blA2bP97I
KCKUawan2l0dzL4DJ5bSeAsA7Ctxwp3MbT71pRBhCtCJrauixee8S/DuBb5Y
fhfNfaVzdymQ47yeUc9nZthswI04ONNK0w92ZWRRNWLLBdEI76TtMzUDoC0G
SP/pRi5Vyn0/2DGrwVLIs9dDhNUMhYar4SmxM4RC7JzoGQuAfOaCntLPE9I2
Je9+tlviAI/DgI/bRTCT9zTqLfEnTU5SX8Mt58KP8EklrN5NPFXqZqHi4fx1
BXrLBvI9NaTsZ5g2kRWL/lzKcQSojt2L8os2IFblVj3Rryser/ZsIRXOKnBd
6rxHHlbmK5C8cNf81TJrH630hyDfXKIDN2HmLlxR0J2nCMDb+tml9iXM7B6z
BAEsplr3aDjTHOhEKfo+iM2TEXaHHmW7wf8abGzwJZoBs10/arvkMIAcLK9U
JcvCLEcvlflyfZ4X8onezJ0l56Prp699nn7XtzsizCesWS1ZRR9es4T8wzPt
uqi1spCIIn9kjj8xQuYuHqmCI4VMd0CBwRFU8eTRqkiP2izVVRCqTSxRD5U7
0iG9HJj4MAKYgVfR2uOEKJ7fWsw7mOJyefeBunHQ6C++xHZX0w0OKpwN2hoV
iMcDP4hrEwxNZIiE7YXYwXW/i7O2N0/ZYNbbyDE3x+htC8h/ojwAQCIR64ff
SJC/iM9okM5LnAbjjQ4bBbhOgpgCWIOzBdcK4dPzLzcBqKt+XMIvjWxTRpFU
q8Xqr0esgkchtUMf5TNsFXzPRnc/9lv40aKaE4ltuu6EoeOxk9xWW9K3pn6V
BFqthn4NEK0Nu2UkzgIBEFUdhvR+BjqFbDK35kPE40di5u1jd4bhPAVCblBc
p7fUMdPvChd0fv3xiwVrztdsh0EYNioZ/SV/vbgKP0LCSXlVxWd0OCzav5Qy
wlDv78TYdAUPcs4XyKni8IojmO+tXoGMt45fBsjoTVFVBAZ/BHyAlxOTnCsL
IqqvOLaFTTUhUgN8/NzyQ4X+sNjkDRdO5b8+00RB7CifPE+PdVRdfC0qLIPa
GXImtIu5h6P5pNMxJ61Yw75C7tdbt8oe5VLv0TyIqXAP3DNOBpiJexHWABCk
lzjqLcVY9GtJfsvTTuBGTmV8r8IxPql80KNxz9IyrWccjcyXJro3+HPihEjt
y5KE2i3KP+hkNj+Rdzqvk9hOT8+bK5mn/CSIxy/aTsUjCLvA8PbMkXep5oaO
RUt75ll1cpfFmEwjSOpFIbZfgHT3BFdSLW5mbijqEuzYJ2SpQILB4UL22zUC
tYIKJA8fDj53O2xtKGIxjpxUM7tHShPF7/yQ1o8eGLrr50gEUgjh64Mwrg/f
mr97sOnSCrxPPSPWU/g4YmFJIuSU8CXlMNKpEZyrlaEvPTkI5MCn9IePGwW9
FeENMIm7cTo+Jc1mn5PP2Y0bp0DN/7K4jPrtwfw65/sPuOpy52OE/E2wjhSc
TBJO/hRU14KSDp14CA2kHXMB6ysXkwPM8Jgvk3VRnjdxHf2JZQMS2RLR1TIY
I+LNikSnFhCMo0rGw2fVVtlAtZGIC/b0cgQb15q2mwUl6kslPI6NaqFd8AHj
RqSYw0KApwaUcxlYvweUeAE5ljVmXG4BjhNarvB3zfpw/r6MTn5qDL05kH0Y
49g7DGB0CZBM0L5LQCl/9X7bwoJPDBNeldft92obp3pzanrperm7vv7Iv1vJ
txH2t6qM8txWjX8MOwno2BwDPLx2mXwo5CRkZ5eClgKm/mglVqFb0167Cw8z
YrF5b6arJaPHfXVSnpicPcrCr2ruL8RBiKW5bm8jZTvJOQWwq7RpNo/sszkQ
wHRu0UHGS/QKiybkcqt6tnT+n6VZ53izV9+8c/VAcMrhaWU7W2RgqBXahYr1
FoeB5u/1n/EFJVnzH+uaUFLUHXAZyOU1IJ0B4DsFkzVZs5hPo40OShwSs0Rx
R1WzfE6KE5SbFP1cPJmuchVx/Ge+JUMcJEwUN2GZM+5hdvpum+vU8FdNnCMH
9yx4JFgbi09mEp8Np68JCvacbDVMtnuiCqP8liEHmrrJemZpxFFNUCWdqpMk
7FSWLTBEBGRgfPgE/AcdnY1gHLqz643l0/LUzGVoylSRtE9gJQeolfcbmcQd
LdoNyGmEAmodjgIUpJVSyNHUqUXCsRYC63o2REC1TJe4vsbxYjAve1DwrZ+S
aicwequT2ZC45fixnfMrZYC+E+0iv6M0T3SrTyheKKTAzmvErwxQR8I+HeV1
7bVUAzIe9bOU42xVTOCR4nNStQMK2lDefNY8KG7+4KlHAHj56IQHK7LRGoXV
d3u3v5ECF3ozKkpBLKqPLkwIr0vQPyehEhOMyrQDjShmGTzazbGrja9WsW/H
ocavdSb3s6r769Hl7ZLEKENFEMTSjt2Ji2sREnavdGnOntZFkWYwKhoUj+1I
MTXh1RAH7h+SPnsALo2kBFCoh/s+Rg5e08XAKW8LvzKw4XKF+mzmu6zLOp2R
JabcxFRtU5ECWJ424bCPkkFEU1rzCs34iq+pLbExatydRMbAxA50cHdQYYkW
uDhA+o8b0VdnOD06EA8W86eCCcwMxeLKYue+uFhWuo1xYvAUcpgBcP8DMRJR
rtaG05Tws9NCM5gBeWsNLEI4yRGEOylGe8lizwFwJCjyV+JPoOQvp/MINVS9
HHYO298a6kB2trlxz5XeALpV4qkBBSp5scu65OwPmztUTto9RR0dl1nS/VRB
khqiAHPFLBxauJcLAEMjay7wFNJ/tgTLRrMahlQhMzfO2DHNkbZTTI3g05KL
CB5JHPuQf5U2RBRHhfw1a8iYnE6zQtDuhKvJXwrR+DV2zONBtTtZfzN6ay5N
1ZxygUTNk186f4/dqdevlmTZFYx0walaawnfkgvG/zQuBZ0r5nE8pcxXdQPV
r6sXc9MnPJWLBRajlz8utulosB1SzgBDoDpS5Fh56lnTAsSaWHevDhDUTas0
ImROwgji6jA1FbyTFirzAhfsNSJ2f2OA6dwQHN9b1n9MWyu3Pd0sT7ffSMuK
JPjUu6Ji2S+jsCBWLLSb9RNwN3uBEuNoal1AAywKE0GnBUWCJ411Dl5LRRDz
zYbaZc74s6ICg/kS2vTfWtQ3SwZw3yVRSGxZyTyObUiaPYl+tSGkLMJzPGwA
R5Z0aBZB3AM1nb8ViCflGkUA48XdgaRZGlC5VG1lQjBrodZSBD7YxC1Ys07S
lK+tMOYUHkwJfHg67s5OSMZ0y0ljdRmdTsm31dGv9HCE9SdR6HPSyJTyhOO/
G2YzzXtOxW/m/H/GmC8vj77yKHLn8ZuKGq5e4LWzkThyK/OOfu5cZ2WvwL1i
4tsa+mVDuWT5fwF/suRZVMyLEFg45mAmDCZ4vkTkjPXVV292ePqoeMD37Uu+
OcgxV/Hoz1/ac0b8OqOUHdsa0QtU4g9U8z+Y7auZ+yJriTL5zKJqxxiwU9JP
pl9/T4d8/XkXBBE9Ks4YtRfBlwvpIj8WTRpx9CQirKjKZy6QIlJzD10fvEgZ
2IBfBOVibXjEFFjsTv9LAd5ohabelNT+CqugG1iU1nb6iTpdMkMrDb/xrS17
6t1lZPG5zui4ZDqzj1SKeJ5AKCOl5Bgpes039syKKTLtqBwLiExdkk/nFL1g
Yz5uokYTj/twS1Gxz9q3b94X3XlHPpeOdyEv1R1Mg8n8a4vLvoKffRJIxfZW
hUKI/LG7JZmQafWxLfgHR5/TdnJ473vobe3IE547Z2cXcv/r8oQl/D7ti1xc
xk2Hr8T7bB0Fd/e5UGGAqh1cxJQxdXH/8jZ9Uga7IA7/hviqmx+RYLH5sArB
Ozzf4XKwooxPBSXYKxdSifPaBCo5mLXn/E6vJv7n5vKw2PbuFE1YP7mRJ2da
l+WYCnMW0NYJ2AKH9Mc+a+FRgAmJCGdHNLZKY0g1YOyegkODgPp0JVWP/aVt
/Mp6cqCL77Q50u3ypty6UBX63yq3hytfNE7M/QBIKmB1IOn2JTFPieIJ7Viv
x+W0GfrM1QznrFkMcclaA8RPyMkObpVhk2gDoQR1hvaMXo7f2R6UhTl33kvw
GbazlVgalDa1GiH3wcYXBDem+45Pygm7tynh9eJe73RjNQ3OIWO2z+z342G2
9+NQ0vilQ7IrsChtXnJMv65l6VSc4oTjV8eagwFsGQKw56pQHlWjfXkwHeyM
ewbvW8RgWTf2DI3YRVDo3e31weNCXycj11ktVwb5rjMJRPnUVPr0RQQFP2gX
EAOviYSQqR6s/Plana7wkLtORPTYcweJXLeZHvb3wdvADFOvsUZmVHcNLxNg
6XcZa+QyPbfqUY8N/eC6Q6G3A6oT1ajSVLpD3E6xXsMs41hHDOOWRQhZqLlf
n1JuKMSF76NVcxhxOA/sDp0ZFjXNmzzdymgnE75orv7OSSiGW9e5K+2cKa2y
IhHiwnjVr+q4rSYEwAPlIs5ulYrx+rWQOQlm7WmInNgvQM7o9KdKUATlRbJz
8FvbO4nUNNx/Rt5XxbOQBvn0WJFgb7gztZybw5K9V9jExqIl2uvT7BQY2R/l
n3uTnh6MoSrXg8T/wc+T7uGJ/YqCo3PBZGSU2J7uAJaPkL/JjEztfPRiKKpH
ICRG0hHQvwWeM4qR7DTOdNCOcakK2IO5u/OL0x+dHZMXy1sSkzdxQ9ke2MZZ
fWo6FUr24HB9FKEIuizfF1svZg/V0J+e9TBgzDoooOpRs/ORRBulM5HtP+xC
fMBe76Xei9hf4l3stMIxy6WdyUfwqsAlTJ4ZhBoSowWZ8NXMxVexUoSBXVeT
ashGIQH15a5iQeCSmKYZsl1lc01wLOKuDLXVGqRGIW7wFVaoxCVx6y35O4h2
rzS0EFdla5lXEiGPYpAcID6nv5Id6dopojXLWVOqgP5r5UHnVszdC0ytCP3x
2Ak2ONV3v358fILTdmK87nPWwi9ptDgtGLzsESvtIrNWnuGJf6p1WQr4zTVy
1vT0CtRSnDYF02V+XkMw/QeP11Au8uOXaFFat/SEL4IJ1F2LAdY7FS9gLn2q
u7oeMepMZrMfrkR4ew8+RRSHr3DmXrvW6DWtGANqxCjQwRy/e2GZw2tNE2Fm
FzFtS4+S3hUEWgakOmJjJ6jBIYh1Mm1P2/MJhFaKyZI0UmxJAR1ODHXcNWLQ
X2wfOW4clcYvHh9kTQN94WxgdA8JB2Tlh2HXKkizXfxivLFRBnjjIzRcvINL
WBwkwAX7UVRqBlVygs0ajQfcOBJ97/sZr9YOUglDY3UfitNr5XVUtqYRNkhK
Ozu/CCTMyLcnrClsq1ZZp+wSDW6cbD3NgaK8OV8bl3qkNnXJOzhqRv7jBSgs
1yLwtCOeBfGH8J9fBmNE4LIfTIEEb6JKuPPg5CP31cBwMkbX3+5cHWbI1lpB
MpdXakazXBjvefrpX4aPU0MtNurP1YQl5QEiC8sgTcuKmlVE++ZxdhyoRbgS
XYasrYFOlWrP7sDOeMSKsim2Ek8x7Epq6KVOzu5n8TlW0Dws2U+zV+NhXzpE
m3lSFoY2MR2FSmUP96j9x9AjgsS6KTHoQuBEkM7hU9mN/1NYpaOny1IN9Viz
tBwvDs9gCI5nsMluIeunmBsnU/X9QGf/vbvT4g54o1MCUIS6RLX6LIP8y0lj
4fExQudPVS5G6yYfmqcuSzbIVAXx2DOLn12dYb/TO8uUlOS4wNiOTVnlYuSO
TfBZwK4eO3DzH/XMUaxhYeqB2eNmP8FRVqW6ntnMoaAe1Q5Js6S3P9lADTZs
EeHvcuun7KWXS3zgrreNEAQsOywTIWXxOXxmc/myJ2LHzkQLLfZIqX35sZLD
KQDAKCE1gHXIs6kaPguDdzHYHLWxH0UUFyOQ2inNx643988ltFDbZTn8D+iQ
NJEWNfMnyXLKz1K4bdTLf2BSmRUaAERjqkFdbKu6n687nTzPVHsxLxqFd3TP
7fSys/5beprpv7vQPXqaGzWlvzK9vdr2WhiRAZaPNS+aZtEFAlbH0yVeYqvF
5s2f38heyXj6rM31T+Eoivq1OqvD3RzQwkt2CpcH5wpVxDqyjh2PDw3rKkcD
Ft64DSQVd/Tk6KIN9EAR97egYt/XAigPto0LEyp3iHS3gMzym9rVuqJBR+gK
ZK1Bm0CE8dFFRAPoCZH4irslJkiW9JODt4XzXKcY/kHyUTtsQZImgb8Usgw/
3tU5gA7E1V/z2ssgfNaFeMBz+VhypHboRpjcuEyifHxUR/9ECkexRlhpLBMW
eud1+VGhlyip8xVdKlVQ2CpX+6sQN2IDWTce1thm+aGo5wwyGVwRyYIShN8d
dzkSYfu9xyxRq1ymXr7ZcrLfHaRLHfkQ5rkejRR6JXWky4xAPhXxDcLkIC2V
uTMk25oocfLsyhoQ0BOsLmzu9tNhMPDW3dbgLH38FTw4/98hSt87n6xdDoCd
AaVNIRWA1laSkg62ycVpALgBD2RxK+2/l+pI1BNUAN2l7/IiA8AJvJ//XXB8
Lf67xsUMy2+IZXDQcKW6ObSPF6CuQM6D0XpqhVWmVj5vuL9ihZcXMpl9eU7J
d/YEZKjIFMLbzH8jr1Dw80G3ZI5Ipm0TxATw+XvC7IESc2PCV08D+BndLdQb
WCH95b/e9iY3VcC6Yl6GQoSHTNEeNXazBblHRdvkqn5HZ8p66Qm2L8t63zC0
m+jNbzFP+HywdzctygAuT8t47RSuQo1dL9KrSqa1m8IvMVb1j4n8ZfJ/3kR3
Ka7JY9pALxsTk16hoNcg/xyjFISYV1GM7My4uNm62J6C4OARCBHBU7+eenS/
b2Kp6SC4X+pRcb9d53I1WTHjxytT/0v1WR2k/yLwnNae6Sf6W4TdIJEOXfmw
KRd4Fg3jDjKTw1JLl1upjwPoINWCUglGCymZ9C9YRCY9fjDmZBbXJTtUtmi5
QNfxXocGSYamr2PR70YxujAOgBqXoYBkifis5MRFne+PZKaPo1KvL4rUk2/O
jfeb5p28KpHspRCG/KyT02Omu0F5FswGtMhSM6r+DfJWK2fIQAkgWrt/skC/
VpmosBtUTvYkcs7bYfzY1/WGp+5Q9KzQFqizJ8uyQCvpYbF9kBoameIjKDVR
9KSr1dCMhswxPjG3xJdi242Hed0zdZDqppclrRJLszxi4BcfMaaFkL9ztQM3
HAwn8eZu9DEkG3g6Wqay0vSZ1QJVVALQ+CO4cbXdE77706pMwkBP+gJjsXK8
DEtA3t2Qwyo6tv1xlG9jcrquIC8Sd85q1qKmA/nhT1kpHVOt23K+bvF30dNC
K2CYfvZ4sRGEgQqU9FHTevO+dLytsAXAfltMvFMg5NcxJedUF/6qniRuTit0
JaNvucX4ipcEIy+kyeiq27g11e6s49qvds4AMbL5HCxQyrbKGku1xy1SVeCD
pgevVWxyS3ppkvf1HzwE434ZPCUVD8WfKf4FQ+7o4RTdfAUxqX9CwAkq7afB
s2WDjdfmbuY4QZIL8nF4BPCfApEVSwGzt+wFE0QBrSxdDXznH5Y9BCIa2rNm
DFAgAcKqkgvYLah34xMqJ9C/cuTi+QmwweFquEAWFw7UWikWLi0wjf548z6r
bbES3I/Phx2OJtFnQrH4/u33uabemM2Gnk9XcMZWZV5Go0fKZ0A7pZaW0yQe
YxwgciPJj/djgasRLXffRYDXX5hbd1PZVgpkwMF5eGWkmiiAATRbeR0L6TJO
fOiEtmfcvkJOPcPzQex7mEExxLMsf/GFg83EKtnMvgl1kSsCaS1ZxJzP4cEe
NLuPcunjjE+51zbOk0ig/zk1vaLvzk9PRGmDUlEw3WJs06wYn/Ci3cY6GsRR
ygQ1eXoqzovjXN9z8y56AsmxLnp43EJVLb7YdDdvBqBfm2CeIODt8Di+rIdz
U780DOhvTvnOHe/9+JT9bpSMWNWZhe/AJYBsJlziOD6fg/wK5U6gjFjHNGdb
Uz3sy5VF7xpNRPEaTj2sDGh6HpzYpULABbs+trzduFLTJCZv1hG79yMzm6Yw
phqbQWo5siq58v6lNCbhs0pGAXonUk5sA3j3tUdDPTpoJWrbf1PjicUNpA0A
Xcheq2hjcfP0hJmQCCObb3OiGOXo4SCxHIFPTSGlixwnMXuTZAZIhV79giCU
kox1xnbe1AnrqrVc3ppW4lVjyrQnzGODpXPN9sRJgmBUUYsHdtLaTLumOcxA
MLBP41QPYaTZL5VeDhQoLkQH3BZ4oDoxbzoWL5Z9N4Gd5JwENNow/5WHRy3U
HdzbskwVUA1xbSOz2ZMQJmuHru0Tmr2Fwhsy8QXaRH9+fxe1nhI5SlJcROun
aNqQsgW3XnmQj2pPCTkJFQ/aUdWFZHB5RuniKFA/iw7bGsLcbHs9kCtZlY4O
JouEhlx6QQdg8ebhNeR1Up+dq/doUbV4jzTiRTGO2Lhi3TveYB4oUal2Mpp6
OF9/I/d9pFQmrPBG6VS3ZO9d85QNgF68N4cA3MKydCqPsQXRQ54kk4KCXvES
h1z+/h3WLMvwyKKnkdsyDtO1TjC1scFyUaiRCD7B+KxTTM12c+drOf66c42H
VuS9eMWbtn0KHph28+vESyVvQ5OtVISK2ydqOqyskLMC2xdPOihSIhoTm2Qn
NcDaEz7lKfxMI79fm4NCzq0sSfgQqTK+qZSvND2TFqkmhewB8PxX9Ifr4xeL
T8fw+hEiVG94l8lLD/Mi3cgd1HDoW2DDpZ5sNx7VJCU/6mz3EgBqlffvciQm
Kl3EJflTo8dlwo/Tmq2Ud7HUmp64cK/0lS3lgG6+DGtXRt9wRdOvJ3ACZywd
Q4lR7OFr2WXSLf9ylzRvCUfE/KNXOdHYnNRUyQm6nPL27Dk0OGClOucCaaw8
VQ4Y9ibILX+9xvh1iVp15Ay6yiy6DEjXF/vsf4+ZX4PEJIxsolq/t0SId9XC
8BrU8WJrGeOeWrHscQ/kRo5XdG/nGzF37XPE0KIafh3xvoRYcsMCxB50Xkwv
9nJ4vC/7uANBtSX0CwWuGRsZ3CUYE1LH4BO551SbOHPXpqqYi0T/snQobi/g
QswtZ1n2xqZ4ZyHL42IUQ1rFSmcxQ9phaZkCzWLBgW15nChJtWgSqxea9KnD
rlfCo173CG6wLTQVCi/EAa503FrbMo95JE1rJo6sXG4+N4BJ8jzZf4BY7Dvk
mX4ke9vvAd6+92o2HfVaFj5YlFkT4MRHCcYxwp6IRZxaPPo8cgPRBe/ZbPCe
keGWp/qSpJNB3MTMHonM/kVpQIyE9csl6+0YSwwc60O6QF9HqyC1KUhkkCvJ
aBhqGV104PJB9IGXormzznn61htk5TDHwtdX3TnnayKBFvTBHKmWzz8BZ+iF
Un3urzF7ytXokPsCYGU2uDl22j9dgYh+WzPbv76DTWenafqalBR5a+fxD+ig
slb/cJOeUBfAWGCYJtDn47AAjW8nTh0LuRaHFmuE+zIRgyld7cppjWSnuRqa
1BYiQIEOidwKTP2568ykcqKCSUBYlCRt+Pd+ttONE3/3xfwVgNql4d85QI1K
9FklaUzxphyV+TWkXpZKUJd0zqZ1OrS88of4uIo6kifbgof7KcSNUQ6dArka
igg8C+Rfeeu4ZZ5+LrnElI4F+wPMu9VEXgHvkzVXO1qGRuMs9VoEjjS2rxco
pcg7AiITxmyKLN6/H1nvs9IDVizq0sYCe6crxiwBl8ZPZU0Xe4gdj21M6pZN
83LTLbVq0bZybGzLIYmC5+N5fU134CnbMKlaVeWYDwZ4pk9btoU2007XBwHq
L+H1licKUkwSUWWSwnEmeTW6o737l50I0NxKbcUAQhLGWVeauFFLOJPVwQ9q
SWftVMgGAGWY8rNuOmMGrkNh9cZEciJ7MH9BtS2Nkotk3j5nZngha/yl/+Ke
0y9aZxl5a2/bn147wVG57x2oNBNTL6hiF9rKuvIbrDBumie0ZGuIMYc/DBTP
iRA4s4u+5U2wvMfodzY0q9QmHoljX0mShFlbvHqhvBQKuMBNUpDqb7kW2fYY
6aDC+YmFih1lJpg4SisbU3K9jF32o67fxdyaGW2roMBx6ODKysMxIVz1WxDa
yBsU21O33plhAu/9GJWB3c5Bue+CMj0rftS2u7ocvWrI7HV3ZTi3PW8112Yo
XSLLYB9Ibx/IuV0xe3tv4pwOnxq4PcZTBzNdGgH50qVr9K8lWpjogqjTdFPO
J5DP9QXITajZ2pMF5ixaWJxDrLCwYsqVZcy3jO49uhuGOdgkQ19anRTq8RLz
ElR3elaDj95+4NxbyC45hrLehQz1P9bKqr9viqlAG8h/v0abfw7N6XVJIDki
r5o4H7OAzJJuS7muEV/fT+L3SM+VUifwrzyIS+wRv0ROf24ajHJt9ZXefvnr
IHyEOKDh/SR4rmtB+AaXm46M+cz6v0n76UvFyfMP5JnstZg6f8Ix3x31MxKh
N7xjC4rr8v8/zKtXXt8ocpQJDKfupX8olV8gm51gaZ7m0GFVT94akUS4zBVd
drKa6XYhL0/DmeW6wctN+tDcMoRytwcoiRb4F1oKBtFwAoKRWeFZuk4RoaS0
QlSsisB+TdYbjwQPJ2Fwwr/LAoF7pBUMrVZ2Gl33TaqzYrxgPjGDYpAboruD
j98cwo7o/SeSzeFjyCUf2FnSsqhSeTdAYvB8obboWIEVE765etDDLtbBE1hp
oXVo70hKlINNzqiBgX7+m2gHExbeNIKpH64eq4g/2flRSwwW33St0+xFBSbM
Qw5Y0WD/a6Ob0NCcZfodGTkXi2nfCYOVtMdKFw4lUOeg2f44MGDdS+eJ9eGa
DRpQQyd7z04QIxetFh2GjMFGisBeDmoOCGTsE3EFqJHMuTrVTBLRR26xcUI3
g9XatNtJAaYq0Z3rUQlHSD9yvUlwsxpvJecC8/4LKkGThYaqDK0tJdbXUyr9
O82Cf2LBWU6a+NLrj/4I9kpz6tQL2VKk+cBB/Pey5cOVrAUmROKfCcJ5rt/e
Hdqkrl/h2lLKUPpeWvTl5Xok1aS0lAEu4Lb5R8kibgZoD2/RScOJFktfmH7z
q0QN69hOJOkpaZoD3n7PvUJJ76mfUSdlLk+JdhV2pGxIEzlCN+Cw4M2PtXFm
aPTO72sXVXNmOfx6aBrAGBI/m/vnmSWiQnW7t7/uq+2Ysy1eL9E2/igrWjAj
a27c8CatKgliIQYEYr9KC8INZhiWQ7T4phfDEgxtu0HGc5EZpg5sqGqY+Q81
MjfuWn6rI0jYN4dKwKdXSuAmj8WAolqnq+8/YAy/6iOqn9HeoK0g0PxR4x3D
SH5hxap8UkHQCmkmPmnvZ7xmlkNnrA4dNasOujA+ZBaf9A53Xus9ketGQEMU
mGyrwmNtm86M+LGoUu6fUO2Xw2uf+AMwxYQ2SYWmd3mSDd9tzNIRiHbfAelv
XlqAGqrIsYJFMwRVr+WhmcVmJ7eUXnWOND58E9jJdNYA97kxjj1ItLF2arT3
105p2Njm2e8in/WfBFrgdsKkluhyY99pvxmPjw2dMmWYfu9qdUZbL2nqMnl9
NyduAlTupnmeNpUK7t3mTJtCkOc/B+fmkS9dZjTdOdipml0xUyKqJiiSVROf
6e7a3gowHrvwRC+WLSmPrZRps/BFkz+KJmZoZqM7rnnOUDfVnL/caAEgYyHQ
2mF2VeMBdIbR9UigXfyuS2pYNkKkwapa97/VvH5t4g6Xyr55bSPVyaFlmeui
B9W8gN+Su4DZ/y20MHSDhTPPkyplNlafS+yy0WRzhNTvh96EBebpIM06gaoO
PuKnuyJnkhB6195HoiEV58hYaGiq2OdM+CoJVXrFWRyvDGeskKRx/tAtMlXQ
Q5435jSJPwD+uEc3Owe/p4DsSK2NbgNPuqZEjEVk2vIW4LOneGxusOoWHt69
lyNB9H5vqbqMVOp009s1N8pRj/FGtcEhwsUXgEbInIUYwWTxJnbUAzUd6tXw
JGDGjZE1duGSPzEUH6V/ffRh8t3S6DzLTxJQ240YK82qltX7imRNyLZxIHnA
pwbQXszdkjow25FMHlDL5yn2vC1KEb8/LihOVAYPdNbLfQo31vYtjqes5FfA
EDbBIllke5Uilaud537rCEsAM9i0GeakS5l0J5UUUh9Z0nCp7umrRj8CeWXQ
AF0XTF1pHtUhY+ILiCZpgenKi1bydNF1X6mfz+RCAu7VK7ByM9+MzbwjuQKj
zYJ1xx4gL9TEyoDXfrxdbk5wEEYcZWb2Y4xXy3m9AFh0ZkHlWcppA9C4KvN4
5s3mFGVP+FKh93B2k+NM7agd0VgupxaFsUwpq4FtnHB4b9ibkchUdKZ9//+T
gVd1Bbr5df3GfMQRx0F70auMO+HxMkDW55ZEkj4DeOwKJp3J5FsWNg9ky9l9
lquNpP0NEg1HF8KJ6jGUyJXspiufRRe0jTq0uXLvJZ/cquTx1CH8PYqxjOES
Zl+Hsyj/pfHozomed35Myw3UQ7oOcxKAvd1YbOs5ZD33H1wrUdGyFNEioxNe
0jGyMwlv8hjjtpq2Q3LvfPC+VVymly4LGdh/Wb470+Cqerkxb00fxgtp01S5
wVslhUNGmxSIQfevaKZG1tNj93NyrRCO9O/uZdjKazUEYGQo3x3BInG3YJA5
Ru8KnAxsmXNUIyr2OFc20J6xAaDDNwVXHmtrM9grX6ZQ/kKDeuJ7QPdo4iHr
lIlyXhVtRUtXjNFQKM2bI/DFB5+qJDnp+iGKRFKjNFmVlGiok5PXXvScGmnl
f+ArlY8PYS83vzhKMew8fL7g/WZmQuYQsniGIB2RHi2Wh5StDJkYEXQShfKU
mLJ49XBQYSFHLEVIKYzLqF7XOKQf0ytnDaLM6bn/GnYEUIWzTB7l2WhveJGB
HFxAorV0Wwi4+orKBouM4vcUEsZWu+7SnMSbl8Qsl05U5D9kqijIBXquE5Y2
DqDALmmE0gdw/gsUTKRF0jXK4bweLV1lo+5nWS6IKqs1s5yMoiEwqBUcjGga
Nka+zMYfsMGqMZc252U4RBHAuk32q1SWJ4+kSe9tVGv7ZZCreUtwbACMNkgT
LQ4H2FHZWjRCrxqfvty6DEjzj87IPB6m7ePbP5JQhBWGwk83cg1IwWKLqMsv
A+Hw5rhv8XsxaiWY9iE6RBaKCUYoSZQOm18pAytLRyK+ReGT0VUeABjYIHqs
IkE3eMWIAr9EI6RBpDt5etNJSYrKf8Uiubwn0zS6lpnVThLmILq1X81nLTQV
YgSU1RTzg77+vzB+CjUxXxRzJdbTNhm/GL9JM8ZjJX4JbyjZv4N6U5PUfdVV
qjYtBAx9UBcWN4cppw3lldgUW2B53SwuHlkJJZgDH0a8qxDpV8wxbtBoeK8y
C/s6ErIuV9YPcKyBkzUL96OaE8r/IyQGdj3V01zKuPGMZl21V89Pivu2uAuf
cNtaRSDxDYq1ree37SfpuBFt2wRYMDIprHUvgEFi9rx0fBVq86IY3uo1T6eJ
n4zCJJ0ap/dxVSzCvm5/Sud07UnRAMPD1bs5sBafeHWcqZKYxeYRgGjaUsIB
VNq4TuUL7Fc5vwpkiGPUmUp4Kiv96OYJ7vqwiebsAaFLicTpNOHnRZGrdqcU
astacZhoePNIokEoBKXaDo+TukBkpmovxgz6i3+zYuX9RtiEsBE+LG6jZMdO
KeVSnvxTf5ybjhoeNxUrD6OZu1P6GA6vdhITsae8EJgJ4un0EaE9glm6lVbT
PNJBbcZaHa9vVa0uYb6sB+bGKLZKEi1yxvUXpg7ErbWHburUt5FWgd+dIpG9
/DSKeh0DEohs1tkm4Vw+AcNS66LX4FzxaCFCwO1LTyLsc1CmEJNtWLMT7pno
y3+uFz46CJnUo0O2RkD0r3ciMI2VwXbIGIgmvQV8HDFLSXPEg81Nbp12Wtze
/4ySMdLguuhq/Xrdf/flCWv9oUtahEZhCVLOGY0gkGjki0N6BLpIqkcg+qJj
KWoZ46hJI2wULJrHn4zJ0R42aDJarQKo8LLyFt59fTatxzQOZQbAnekXCRAG
w9jRSTv4+KkBXGMKkRGTM2A0z1nFqHuNauRbpQqt6z6NeQZQwKaTSxdJfHQd
eWLbClngwnzTKD50le4uZfw107rTQ1M5mcEB08t3vQhbjfHtTwTi8FDVJH8q
v9i8aKev0kMQyNzrlYBK7Jl/fQiOtIwwOU0nSj3hMDjZI6jca7UOdsKk+7Jk
FL61664lw2aFX/lGJg9DtQgJ0HUXwvHgRPdDnMCcKRYXHcrkZOO4n4WR6M0F
960xVnO/63S1tBnROlMr5GJ1J44ktuSdRJLLW1sPsm8yWpetfLgTgzFL8a50
FSS1rEesHjLGxmtRfG+aClyKSSgXlQ6hgx/VzyBCoXc2D9YD8E63RpljEIUg
KxrJfF7pbrnzcRSio9yXD6vhtUHJVkL5wqF7ojlVNK3V7uM8SnybvOzSctNq
V6puAdv94aGA6ko0qOW49tJN0px7wNC/RSdoiK9BksJiaox5aTrBcwgZkDTv
8dy70AIvUDPjjX9fJyfG1zTiYt9L1SHGz19w4VuOnZz8veGzIeAzusFx61sO
JHK1/nIDk6/+9cXtaP8YpQrI2nUgQaGJhDAmiLLVh0o6DPWQMrdrJdM0qijb
7rmDCsp0Td1D2r2ydWN9pmNScLXLP35vZMJsf+EIGQD6QHRwEmpgAmCU5Z/J
gTL+5ZijLrdoEbhS0UdFViS6HswlNe4S+3kDRiZ++H8/0hyQ71jM0MgKJK4l
QsQKNU8OWC0debQzeEXaVj8OAWc1LrreXpDmNEcIdTpg7ti9q/cOajrlcbhr
5/01YkREAj34UujN6GV4yOIMVjuua7IR7hZ+5PhH98VeFqKxm1uJZZ9gNs1Y
Ln+/4tmrUEZ6ddsoum+X05kcCufhGhJd8GPgbBLH52jJxS47cS/AVo+u4EZN
9wzgxhn2Yk/yScerFjd4mKGAe+q00r795V66OR5+zR7/X+Li1Z9Ndq1IpgSI
WAFa2RihhlLKhPF6fcszuVrEZEf9cnKsZkOaKEa+T0eO2SffuSqkMUPkJfLp
qZWq+o/Q0+K5TDl2uAkwM3LCEAN9O99Xi3mxh2tnIPApIFkhx2adKdAqyUFG
LjFBakjtu2pYOXNAx0110VbFk6czTUgSNpn+FABf/gLDlKLwwzvrxcodKxwW
9Xy/HjM48qdxeNv7rR+i+aTkwmmIXpjZNlrejVEmwFGqTJUhhVDo5sQJIv40
PDY6xv2A1OICBkOy39k/WP+SLHAsk0UCUPI5NALT+qncyUvFkGAO+l7wwGII
505Uy/ITUanvgTLyCHug4aGMv+2ksEbMFB0JNKBg7l+drAQWzlrF446TxExh
8I+RYrLJF+TFTz7876dzrzuheczUpCcOhQFhJ/H1/XyOpZRDyyALNKs+D8qU
5+xV2UC4VhSs6sp7944oOYrRupBZMD9XYBA8txdzQ42B9OP9Q95qqmQgxN1U
TnvANhSeXN1vGVBnuMNrLIcLbI7ZMoyj4YFq61ku1ptXtGbpp6/1nBt7AOfH
i9QZoZAe331NrERiNUxzhwcCeXcOECRCGabDoKGylQA9yS8/SxvLfCLlpKWD
6eTLZgqfX+khtoke+f9WhJHMoeMS2IZeh7flIAoY7FiWV3EuXwrPWTv9BXt8
/1OSs1lsizGfUyDdTxgCHhVOz7ESokBllShZe4uZnaPlnw9q4rYEFohsGPr4
W407ntGMwV6bZEEVGejPv6RL2UhDTikM16w5NEi2q5+0huW88VCnHnXIyLfe
MElwa1XYMRDnTtLppoGAzyjCV+zFLi8SMr9XqFHjiQGXfHhq0o7MJfbTDcsw
W5Tqk4KcVofm0ngQR5afNZtXNuyxuydw7rIz3IiFe0C400e3aCYHBSfTB0S4
BuTlMO0jy+hXPZ+0s/8fKWWsnHVkDDN5W6fVrIc/QwKQbFfpOhxsC45owybG
Lu7LYX41uXDRE+ITKiBFgb/wnHFUW9uLbW/Ovcs/6T/3/hSGaxym99XSzWYh
StHK6OzTfr2bnkJw+MaJN13P2Sw14i1cx6K+e/Z8v+Iu22S21r5wQNNeQ3J0
RScqv6PnBGEL4Pauk0kinJZskfU47C5jrFDbXUgATpfd8JL1F255OpgJJOyC
Wvq72ZXt0uO7Byko0VmMfG+RF9YY1IFfHj9If0tLxFyJ2MEyP2VJaxdV6bm2
QUKaP6GPhhbHnuobiEnucFxPjHflSU577+K/Qk94I7sOb3Fgy9DeDVlPzzyZ
W6JvdaDvG1e37XkTMQ2YfSvig9RyLEqbErpAZ7wrBCMswyYuxrg7TgN0I5IF
VZzIyuAlu6R3nn9yG3p8x++ePobmViwknlA3wNqanEQ4XrGgBO0svA1K/dyE
M37l0gjhauIL1B+Vziy9Tz//uV//NUTFyEI3XvoBSpEsrsFPvHo4GhbJDmqH
yhhR1dtr8LDnbZI5lMGWE/rAofQRt1jGXG0RYpWiplGfBl55f2gQizt2NUld
q0eskAKSkuzMhFJZZOCwWJWLYX+kZbFJw6FajPOHN56RJqe/Jn2LHvRd07nD
KQzAtuXfrEao3hUVKACO5osyU/Qp3RM3hLy1IMPvi97L4DEydv+JnKiAxwW7
a/EQdDB547zjiK25w1E0aABRIgAwwBtPSm+S3/dSoVevbzF1SV8uQhlN04QY
xoRCjw2Szqn+hyw5vnRG8GPVBcQPCoifknvMRFp0CgyrlRyVf8dFUAbUoEoN
2Vlt1/j7by4MHIXcU+NDElBCtPjWaKmupAWMcr+LZD1lgs88cs8dL9HO9tAa
qBO+IkbEpf75bze7DTzaT8VkrJORSqomfFegXMH5Pw0PVebpFi748KgSpSrf
w0dRUI4BJlCrQl6SgbXoscQmpj/QB6+RD7pmbESiBTzCjiqQTlDhcB+2A7EM
bbb1J30ZdPa5LfMMP7bUfkIyMjlZPCxMX2YMYVkUHxm5Mg4hsd0bgE8iw7o+
P9lGssEPWoyXs2NyqwFwH0yOyxKGp9dCOczOk/lo4eTYwWg0HQO2skjU5maW
Z1R1XUT34RnpTmNo+u0OxsPyXaCveQ6nD9QQupfPuv7yZTSVjlPm99aasCsE
ZYyt+I9780iClHdIqF/e3vs4xZ169wQCQzFOpmUpmp4cBu8E121BcIS2sFNz
WJr9rqXVNf11VO+F8JHYvO7ssN4GOnsjzg6KMXHrSTuiFoKK2OVhX1KMIcMt
w1jOlifdoLAIdQtasj2Sta1t/hwpkJgTONtmmQoCJYq+C/+e0wS2d9IipO39
fulAV5iRqOjEDCsSkXFEHVgol+9ILfASCx9wHMq5MP5NujxqOQxLD/aBABop
SMPv3nGHDbUHszL6O7AOrvWa9tqsl7r9VItHiTv8N1NguDlRgCi6zj+J5isX
uuB1SVFKoRkhbdENsunX4wCGUVOaReeJrWta8kx4FSKoHwWyQTAa/b/EjoVQ
gWmcORmWrczs9zGg9/MdFjav76vcNj03ta1q4sZc+VdLIKuivzWmuh3jodCH
cORUUy57yHSSh+ABvh/3yAakcyAJTSfQUW7K9wWPzvg50U9mEZrIxuskpWyG
bsoBUVqa+r7xAW+fhzTC6pJqE5T5M7O6JmNM4kXQWyfT7IZAmK1t6odGTB4d
zoArlJYg/SSg4BJTSXFM3otoo4Mi3WyUc6uTq7viUlgbR44wLcI3Ea/BdGHz
udFT4eJmv+q2iA5C6HdoZ9FNkX1ZCyCqa3RL5b3y5To7dCid9AGOddEihdhR
V8GPthy5ifXAMq7v34A27PNXNmZT9XyIhsIv37U2GC0ClMW5WSXAHd61iV24
Q4FbnHp6tswF/xQr339CCMDS7rKU9PlC/i8FLKQgMvm9+WSQQftB6+RqHazc
+py3pfCHIAJE1cvO1NkNA/oogP0ua50RsDci+sl0VQS7799+1W7QyAruCgdw
YOLv01VG8JFUuHO3CEPdYM1XfykQZENh0YuZlONHd2L1jzrZsbFUY0rlaixy
7X4a0Fg8x+lfHF7CYPWZlBlCP2d+PuqcduIH1iy5UtXb8qwdpciueOvQpkQb
Lkm/6pTC2GhEaNxGYb7fd7dOX5rmeBtUuej4+djwf1EiYq2iovgMtHl2NxF6
Qe2WbXurEhEG7l+91H30DEQCMp7ADM+sAmtcDNVTiQpU5jpExia8xyB7acu5
Db4ZYcJHtY71ze0/c+mrmpVVbZLVMNUO6bILe88TDxueDtCk2MmWrbdg8LZn
DVblVJEqrKMxaX7cEv57YS3S1iopt5nuY3ybmv2X/F87eccSKzYYhEYpJ8+q
yyA2al1DFcqzqONQpUd8ipXpBYFb7Z9WzpfNYj9upmGr3xKvYCPLqHEiAEAr
onDkQ1wFbStfy/E/cT6mARnNoNYaxyEWvxaxwCvkB3DUg7C5mIVjglYkhJ07
GQhHd6S7z3oXvtYJtnTViIQsGsqP5huqSuT6cocJFVR6WCxwNejH72vm259l
/wY336RwgW0GQYd3YsM9dUr23Sp29WMQz+XaoDOPSjMui0djaDbebYOp1Lmf
62GmNk4MK4vSimNrAgJE+xrRW2o3cTePWkNG0ypjIEeamH+wAxqvZj9gObTB
/9TjwAZok7leRBz7198jvO5KckfKQYRrCvDfbD4yMmIuCaWcdJdmVc7jrNt8
gx1kAIRIXpSQHWaCHwcdJ1PE4w9JhxZvnm4sFH+222o1bBzZB5GS2d0z3kzA
5qOxy8ETgZguX+HukucwmvhvF20TaU1EVMxa8cEG7QqWhLXJjf45AzoEh0LK
KH0RQIWjKv06bl5ipSsXb/2bDzMQEcOOnMn/dDcyakmj4PJZZF4kfVtvBUai
e7TgoWhQhRRqSv/HMhNv80RTg8JzZ4+4szIJ0OVuvVJ5tNwiNy+wAWKyYOeR
SLDx3yPKusulPk9t9o/GXMruw98qUcck8MgDw6ElQ1hcQTnUg2HD9HpSU9kJ
BYX1ovAO5DCrp0trLNOm8Z1DeVT17VHJg4BCYXQz6EvtGa5wbSxo53JnS1Io
162WlJ2SckVtg1K5KX/zitoX5voNxoYoRapw4+oum6wHW4M+AgKabBnmDVbl
lwHd0naVdOGioG8l1xSJjOkCNiYIssg41DcGtl6O+F/q8vgcbmOUIU9l5BIF
6ckC02kQUOPy58OY00XM2bPayUjvSRM1g2jhnGxZKUwQwzQQQx+ppTCdF79H
yTCsLAbOpqzMTt+lCZleX9Q/Irmi5RlfvUBtvXJ8suhJMGYqADMTPFnA6BRJ
7E8YBsXb1rewngN6M+b51fvknBuk56TGe9poqs/PUWxTabvh3/yXrzxmuj67
rz+w8P1Ukop5dP3A6V/uUCSRgk+KoeGi0kzHA1M8q6ZRAH5SdmNg9mZzoT0f
n1RDaktFjv/eMgibP0zYQspOnjosmCDLeJHxkT5ivl89bNQW8n5MVndYYWzA
IcI/2c72/HCAT6qq6nqifDKJXtGZU9wf6k8I3Zi40B5fCMHiuMesJtDXpKzV
HrZqe8xb/D3wB4pXqP77sP04QABHeGW9a+Q6fHjr3oa6b0g4W+S670/GiMvi
w6KBGyzPJdUZ0bXy2Lm4dA3M90zjdv1IwD302xlxAqaHdNBjO4V2nlfKlJDA
MVp3nhQ2uq/IV1lFHo74nLoconHdaz93TFknRZlxua+gZT7QA11/lmIUwtIc
vbhdUuW6wl4ynRN4kmRKwnWTY4DraXqQ9AIJ+iGNqgOedp4ZJwqga1S4y+TH
Zoo8XyH3sg7IIiNqSxImYP2jrS78xeXJpEhQHA+YnC2F06vLVt9SnO4N7SqG
/oJCmnDqn3s0lphlUFPtsoHFekwtg6zVKnj02JOsSYosIMfVGzuzpx/DXaM2
vfKQjQqVh9syVZVA1sQeQb0qrLRMRboaVknkSJECL7dEAd75/Ph7VhYyPNxs
4BH924Wmj8mcs6dL8dn7uHDLiLNGSSAonBqEwlM4aAC2nxhnbAaSWiFX8zi/
YxRqhvH1jYE/1UyVFvG4ResFsF54bcQLrEklCa8MnjO2Dd2aSjjoSUgXyTHw
ZClLH21ef2SmLtLzeXCDBVo/8Ccw1U835ESIX3VSrW8+bYKOI8IxS0NGj+YS
UHN2cVrzZOFp7WYX5qMsWaf7DYJQ6fjVK1FnC8VnJ3AZUbzgpv5VBx4kWYqX
RChQVfkGqzimksezXhuV+7SJfzlmBNyJ8insuJ7BADdVk52ZjLV795o1Odgo
he8HZ0WWHP7iLO2d7ZyMDSBZEwL7zPQzFEWAdSfVi1khBPOQNLMMo13TwLB5
VSdavh9592931TAOrSu31Z4xWmhkBTwevh6z+E1EaTc7AwEtiTM3toidwJR2
WqVulDZ18/WDRHxET09Fct1+acJgJJpltzLPGM4KCOeBgaXZ9tcexZ/t6hAv
XZlxFtmNHxmvOfQXnRdzKJX4XHxgcY1A5qCNde8OgIeTV8SSgbv9M7kx2itp
HX/9Ue8pjG1TfVgo5Bxag1qGywU7F99Pqkb4of7SPmxBC0FZDlw+SssEpdEI
0LPIz2RaDWoc5neGq81XXl9gRfMKqhNojmwtQylFOUk31XzIWlkVQkuPiTaT
4ejpJXFFEX1sEWo3a5H5sLfJp73wAOWJ3zsLWiVdaNO9tolg1hnnPtXG77dj
W28gHPnSkvrNnIkyfwiB0rEpzVTV1O6/kzbTQ8NYR6wx4PwDTA4/iIGZbExS
yyYHTnPDKExbSuXQI8fRuYkY5Zde2aFpknd+jSqvtMwR7z+uQKMCcLc46sfD
56Lqn/ktr6o5P674dFlQXpbM/I5AWSL9N/yyUb00kM7IL4RssM9gKwUEOyMD
7TPuFJ4FZr4JF9jWeQx/5YZ4PK5mYBjK3+zpsjR8U5jbEBPSaGuiP6be2/w8
w/I1zEvnfe/MzLeMAz9/WxIDfANitfUMkaC494eRdjeAyNk6P6Hi83oaLKxm
pdLBxCXSWxOrXxRVh1IC11gozEZoHTjkX9Sx9SuO6ZNL4EbETphqVWUzNDRD
P8il/s5+VECcqSNnbp+J1cBbHW9BfBzLVuXj4YGSQ3BhdvBF5yLvQ/76WFmy
/0kgWrcsKPxBQP43+ps/Y/Pm/qiAETWFZPNgG33grpsJj294NVeqFdmvGweA
CUkXAJDWt3wmRu38xA2OlTuh8B+BHQAiDbeqjg+pdx9iNYM7cwxjTebf8Hgf
WXy2WWlPDCibGyzQP2DnUxZHDPXVprjPciF+twHaa545FFSTiBqHXFP4wIoL
X1DEh6xqiALyiMsVmeV9jjJ65YoNhk+x0SZJ4pNpIlA/wQNSBiqw1G/vrW26
JT2z3bjoxbDsmMwQ7NEtPUDoEboCMs/85VpkBLMZSK09+2bAks1iZE72rRtO
YXApmAxZFwtcgYq3SrjXN80hCl1xBb+zwwKUgz6rt/bypi6SkaAJFYRFah06
PurRbNTyzR0TvLcPCWfCZcjFqOLlVJPNqh68NKk48WbZjBqJLlwTge/ZzsTE
srv4UFG//yzMTGsUb5rrwixth0hZ7MnDWJuFSziZ+Vfn0fXMjVRk74QVw8Hf
lT/nbSzOqu/8E9zAP96b+MvFeUjqNJBdI+E8Hnf4MVHLPynvi669dkm1r6os
x0qm76DB0MfPJ2q1EjvGDmR95hgBLwZy9azZkjiofjLoMaSe//qZ3S38DbcZ
b2bdw43+/Qjy+jsyYMd5xTdQXGoUuVBHSYcM2Lcm7Fxsui+IAd2XW1rNNJPh
zmkvA+SKA8c0Oz7jEwk65KEKPrXfexvUq2MIpeuq6lTfo/Zq0bM1z92SIfrO
8JIc0SIqa6QOuuPDhxDH9kyBT1dk23wHt7mudpWj2UPU/wyUnpc0Uevfof/T
D5/9psb9UdA1B0w78mPCT+ykL4+ITEGJ2GzdfE5VGxWdMThJDjNb2V5BcBRm
HCP/tiyZKeJrBuHgIIABWTq/wQEu5rMUIiwiW8quflUVgCbdspUt4UVCmRHp
jRjoIrhqV1oDOB6Q/KR5YJeVo1v6ICAjusZ63uJQCkkpDqWNJ2Hr87h7WAv6
MSgBe2sK5vdAS20JoqXJhsJhzmNdXDbNPG3nkJcmk4ENxCb7m5OPrjkNk/Ey
VDjrQ8CcLwV3FG38fFkskzL2936DWXVUip7ppw0kcQDvp0R7ENhvVd+Xthqv
8BmWbgTdEWhvVUn1g/j0kfH0G+jeRDacsV1hc7enJ7f+f3Lm+m2UOrL5E6zN
/BnBjFcS192apbRx9UJkybm3CtYjFASX9zzYQ3tRz3tEAUWBlNUlpUTm7OGQ
b8ziq4846CLxGCHrTTew2IYpnSJPBxQg8dJMxCnvL8Um95x4Jj0FXbt4AOuJ
6V2zphAoaS8ulgq/tFAbZRkjdkan8991c2SW5UtjDzJg8jkJEWST0uU3eHwF
HpwMx/7yejAlQTGQuqwF9jK1voN7wwzL1aYr1Slj39fWdJLZf8cGfJ38NIz0
fs+yO/R3ntJNbI8EJWgTPIw2AN6DHKFvpIecsTN+F9sSM+/b/3A4GUxRU/x0
qMOB/ofEi8CubTa0ynVLioeZUBxMKa/VN3IPHQ/POLDasX97jnZ9k45VFHZD
gj8EgnBPIX0GKoz+Vex+ETqHUae49yeSUbWzT8w+W0qL5PknJtDqQX//Dyzj
fB3QHqnJheuWjSQzUyw5usNVzlWhw3JynXQA6m9utSv5P0LIS4qihsylbX8n
8ertAc8elK3D7AdEIXpocxADLP+U4qHDCUv5X8FVU+k4rY5mFfc/JIuqO56j
FhA3E/FXb6QE2ZiZ+Spqs+CaxjrKZoI4PYCbjeQKUFYKYz4sctUjRry1M3kN
vZrO0L/lK91t1q0fnMA2PTs02cHe7hRSHH/2zUzr+Spm/f6lDTLKS4EmecM2
B6UsgOjrnjSYLQuUJjN4eh/LHsg2CL1wvqbE1E1Z/Mvwu0j7p9ZWJYwhTPTg
xIJQLTAr5hea+heF4rzPCSbRvUXA4WTwkiVqzPJUuu1oZYaCo9yQ2KUTtbTK
EvQMjfSc4c7UKm1WCBH48CF7x3s464Licz/U8a+AxBRBKmhJdVUDp9Vi3Qpv
tT19cZMzI+mCxZ64LqEXmCoQRSAECH7bNJs1lDDAtr4uUeS4hPg57Rmfdzlb
nEUD8HNzRQgayOX9vfTODfCt2bb2O55SYKgzku+rIXtsxAUPlLz1PVtuOSZe
eE6H9VnxkxKSvLcyp6pyNbYWuPabSxRU+bAXuwGgBn3tMdecwcbd4i7IxNe2
a/q7EPskp6u286tlc/4qTNbkLz4BcRpGC4yNGRWD7wZmv0W2knSXbRUIqeEs
1pnVpYKZEB+rVXQDmX1bq240pLb9qXzg6VDlCZxZLX0uFAcfjbmjxcQAzPyg
/deE3UEIMu2+jjwL2t/9GnzD8+6yya5OVHw2JuSORjmUtE5FzxTYbhBiQKfE
gWtY4cQ/Dr5bTSx3CE4TFK9jdygXyp06M021lEsQukdsbLC5l8eYcU2jCOk0
KbFQ3mIG9zsU4croEsLikwpgm639JkKornNkv2M2wZB97uRzzMcX8L+3rTmQ
RMjL6H8TsOYUW7X8fzfBOihDxzN/8yCCS/VXcDukqKfBBLVtHp/sxdHVtu8/
KCRXCqo0wIvUydZMwwTU9Y8hwEXot6BNomeGl6Jtf6xkseVZL7aVmSlUF5Ce
zVMIvpYYnn3G90yBm68srACM4Lz9oKNb2Y7aAKhVKhPWr+KYqxZWPP3GT90c
0o884DKe8rRI+9OWUw4LW2U8anqiKID/mPpIihhz3DVv1QDOU93ZN2sKXoSe
rCCi/VMPLEoDwSyPE3KyTHLIfzXJwkv67rh7QrxxcFJLxPau4UbUm1YXjvza
i1qGdUS/ed/W8Mg5MrK1lVCSBSPl35PnAUHNPz/L1imhAQ8KW8NY3Y44n5Av
jWu0BSUfhN0nTylsz+b2KzdkcO2l7Z4TMJVwxWwypkseAtz/dZnMeSa//sKg
eOZ93I6gfwJXyXsys5nEI4ofP5i07pTDFaQuryhFg6zCk00t6NStz0yqrsrW
axNfv56MQUKiGsNEHJnJDtqaqBOF3+eft8W69RRdyo9N3MFGP3IrvxHCbd7i
6nWej6bauWEOlEn5QA7GZymuJhp+EongMLSoNt8yhc21yRma3uortZ/OR+C1
wWJj6u42DmOMHpBYoPcRXpK/CMV/8AMzgdJkMdBli63ZCTyPdNQeTsiN8dbn
jeXONFWmXq2dtqOVhSG49BgisGEjWbcpzW39C8g2mG+M59zt0BczfK7ytThx
0o+bUDPMqR39k8LAQ0V8v1O2NmTU/10qoqSTlvTLtp10Cj0983MHPwic3OQM
rmrn3avpVL9rwZ86KSVmzhLhHthFZTuO0ujMzqi+5Sl2Hfb4/ZOEhTtQcWtY
LJN0fDPXQRH7iRA1xObm4mOsyLeHT+xbcpYf5Ca4gVVUp1OIN7avo2EnLT8S
E9HHa06iSqaxMl/e1z39E5pLoOZV7CsbkFOBpLen2KCh8E9qo83/DWVlJhy6
54XUOtgwC0W+cpDuohCObxqWBDN6rhnTUvJjEyNY0Pl4bUwWd9pd7BjSRT4F
rZ6SQu3H4duxL752vOS4w4tRtHbnSkorCGJmjQHtzlYjVfvGFM9jTQLvFf11
JJ6YvVBCwu5HVjy4M7L5/l5sVM03ELs5eMu07wSUy8NJP3wBJxLbTk2Z+ADQ
o3mRmkuF4+VmRBmuDRKqLq4ElM2Gtmi4gd4kUAdnw2TqsyNxyjaa0zIE40h4
6rdG5vyn4A0SNxsk/huV9p7Qgw16eDFsQAHrzDh2HLbjLk3543GE67iD8E9n
m/fD2RNsa8iIBDb/vcXjpxjO/HOlf1AGrmMcg7X+t9n15nl7eZBAaTZlMksa
S+0BL/YbaTK5Kpz8GQCxCL7sYeVyXvQh7hJ4SM0PRQeC/J98QEyNVgdGeLCK
F9VArZhc3Gzfyw/o4UWd3vV3NZZ//SjYLbH3XxrUdTFluWUP9g41eeL3y3u0
hb/M2t5zmm1IAgTiRtKYJxd1qhN0IK3kQxXQ0ZHvOuZK53Mb4BgYeJKJWQUR
Vvx8j8luzzFwcF1WWRUbWKJjE0hLR6v7BS0vfuATV9eGhCB/P4/tt6hn8qg2
mtAamQG7FWRsk9jDq9b8nl8O88ooz8jq8eRV+a6nUnRAZuuApxGR5LDh3+5o
XQMZo+wdp+pBgrbRx0sDG+lAM0HFWj3t7jexTO7Meme+zdelzubyMwAL/cB9
j6jht0F9sYxU7K0LyXPsgs6zg51M4nl6Rb1jUX1wicNNclv1wEIYnn+lTVTd
Do5kkWcsUj5GK87TNsugZO38ljTxjfLxkn8/VwlNTF1C/h2kByESC4voBwEM
j5CmXV99fJwkh2u6I7t/IOlHHe0jiwBkKXA74XI2ZJSEsAZ00FGA08s242mt
XCSvcKIdxGVPpugKAHb7MMRnstamT1LRcl2Gq60b7tvllI4C3YCvM+6NAFuM
kYXY1m0ZYpzMcAWmkq30cqZYRkPAruEE56vxH3Jy1gLkhYntiNbcWPPfFKlQ
+Drs0WgmMLlB8ZszsJfq+CraW7HHwYMxRa4/pJ3cZthj2vojjd0TrIOmHuwR
r6hVSCyxxjhrmmifvPuJ97pOnNBcJWqgiB6HVLSD+f8queOFPl03K80+2DGN
945NH0f8goON/MeLYmjKlz0X+eG7JG2RebqfNxX0c68Z2g0XO1O4ewe7wvzd
WaCRcL78Nb+xSvLUDM+iJvRiGVyT8aRmZWrqH7HiT+nlE/qc2gD9IlW/wX4g
KQrhb203aZ8YXJ1Eb92OiSiWyAjf/bW2Yf4BPG5sNlzq5OUpnEctBEjBk+Y6
zciRNJ4keNUux4D9zwiHBrtI9NeUycdBa+yDaeb7AjRkCpKr/O4ikDgJrhuI
BMb0Tfdp2BhC4cOdhavM9wUZHefCorXk2IiZOe4po67QO3ph2Ttm9rx3dddu
1H7UwA9csCA3yQgGh3zVJ4C/Y3ykiWq7lTwHLvIxpM9lMVXcreU8AzXawSPV
qxsydP56LKukN5an7oR5roL2FWPfAONvMj5TdNLFRb3Rz+gMpvf8H6mPMnJO
TjPj+jvTHJMVewc0ha4dDDaP5Gxq+4DSv6+E8VglcEuq/ay3awOQE9LBV/aJ
q22trEUkM+DC1S7A/wjE6nNqvthRPqLC3bEXDb9Mdjm/Bh9H0IRIghjY/IKJ
OAmUIAFMz1/q3UgAe7LF6aCJrUnfQ4LrtyjOL2jh1Nz8V+NPN10jQA2pwNAz
dtolrg1AzKNBByd02Xj8HfgF4VGCemvrWOBr6iTMUMRpvbYKBNyBoACEOeu3
EEPoVxvuy6mdrI4QyQZPgi0IzBYbLcO3IBb/0urEA0Fnv80RL0PFMdshxUu1
bXAmHGT6H81hRNPY/YyYN10l8IV74M1vVPOap+83Vtzn1ty7EbZXbQTYAqUx
nAXE/u1vdsp8K+X9GKlphIpoL7TK9pySUWxBZztpx4vFbcBflr7dc461Vuik
VZtgKAm0e3bXtad1YBdGxDrRI5sJVpwpDavylgWAlLusHnxlLDJYA+tHSOkk
EgrJGKBjudSWW9Ry+aUALg1Ogus6tYielRZQ+AqehC31P8PjARV05KCi0jE0
E/HoeXqGW7qo3RuezsiGPcUXu5Wg0/sM3f9R9GXLJTiBsCoS95jrNszRBp0n
KVdOECQ+Azt5Xz8/H9mfZ7xLo8Fc2NWHcOzDsYqtnn8O0/MrTL3n1ey9V2vz
qtbAGHK/bmd+edUmZpXgZbj2qmOKqBEXGdNxrdNc/6laqWLHKDZSSknng1vc
/yv0xz8M4b4VFzhQiRF9ywSjPYNE8DiSvrFzM3Qrdoi5FecwHyn72XcE7MzR
6hVeITBOLOLTzpzcYp2LKP7hV70UHrHlLZlx/8HGya3zmY0WM6/gJTInn0sM
fNIvr5VRGXLHp/hKQFyb8Hv+K7VHdH8n6Uo6Xzx9dGiQWoXRgzqGpEPlSFGd
zmosnbIVXdY+duIzxfsNn++xtb6WtyCsYAw7oqzrE/b1o5NCqkMojWJEeqF/
vCoYtqENhAHd2VRes2sPbXMDcVrdRtTmSgzlF6LJ9UHUdIWOfM2tM5R5/gju
u+Tjl6SeP/KDnlumqaXkMhzXC4OCyShqo4cL4NP8byeYc8/mM8cpVD1xSeUr
GJ1N4r4S40CZ8Z8RRRwrRyJdxgn8N6ffXpVx1RCOg2USTh8AjBlWYLKnrx7X
5J7WuFZt7LoSYNMqXULH2eqOAphX1JSr/Q3IcRnzEu6xhSj1HGkhtjorJ7DR
dtASwXTEFApZabsI4sK3rUgazVJ614bqAt2r5UQaEXleOm8MHfIjWA66SsQi
6ueZ4Tz/WWMviFUCezJuJeE7hKzL3cbeXHdvmfhlV0WpCqJOjhubgPo0+yJj
7cbJlXaBH+o56b2Fg6/JHD24K4ZHO+ccX00f0KYRfMHCiSHQdDmn3RZF7aDV
HKsr4OOwNnOPXUFipRW1SJ7TNLjytp8zgvgxuUC3PvnwRlQ1qqnpSniHthrX
2iTf7ZAhj1EqbkY10j0aqRJoAh9e3Cnvkrtf3JtRWB7TPFU/qBqUyudYx7rb
gvYt3X8AUVD69Tqs9H+ftlJf5dhBZxiHrkGB+USEAUeL/Wa+6WnBvF8wJdnL
B73dVZ4/QAHldLHMB4FJlSYt7tF6rbqsTSYgvACP2/94qkjOYawYHpv893OE
tosR5nVU1EDpEWt6sCCmsT6r+ZV+BbzpHZX8nykTqwlJeiBzShhNthqrdjTJ
vP8J03j4gztXe0FYok6hJFTr2pyXSeGY+mqJ2rrp3e/y8I0kvosjrUF9VYKp
phVDZ504wyAY5x/dAfx0ieCB1L4dwHKcJHdonLvK0mvnORWhn8/nLd+VjvS7
E2i/3PN9pIQKlkZRnxx7I1B0xoeaJEaHGboYX0NR0RUYem8km1qmuzuxpKUz
k9Hmoe8RtJ6MHs9tR8Dv5FYp44dJV37l8Dl+Mmsnt1lFvzwJW2HHlcEwMdGA
SnMQxoVVD3AV5sG1az71NP64ifTNl/4BSgF7Xsi6KphNOFqzHHCCt9tQPzcA
g6Gm8z8EyxaIp+V3hn9wwXdT/OvKNGdgKgpEUyh1AGMXv1TZiZa5ryLzmBCi
4CjALtqrsszVgGkB6OmwGkmIf6D0aUkJC2rKaLLLiQWQoZ62M4aIlVmk4AsC
tffhW1TkfNBpptoOA65WN72pMBEuXzkEB5LQj9thmqa6vMV8VIATO6dw9jdk
Bz1pnRXnje535jz4W3FdEVvCR61BLq89fx8vB3iMilE8P/AGM3mYULKwqo7j
17qwWWNvHTwWDChyrksZz+GyKmED2uDMtvA45G4X10q64MEzQEZApkDGiFa8
kCNIjvkoD6hQJ7aBl6C3EsvA7pnMfbqQ3G2NSl5FR9AAo3CKS0fHHjEIinBB
ZuGRvBR4ziz5TeohnT/OnJRMpN4arQR+oedC5s7rA3TZLwzoahlHSeQSZo6s
fycHXundMJIn88MFchlNOYJmj0NZWSXw9z49bW3zUvbHi7SsYVc6RJRvTFrX
1mTdSZZVE2bQG9s7eG13pMCLadNzjy4NkiOMgUScf88cORpSDJ8szzIBgc6E
YZ0w4n+Xqm6rVEdhQKJ/egS2xpE4P8YgH/+RtFbA2ZrV2F7KnzitbhxOO8ms
fj6hkeacs6ZnkPrRKFS8R5CIribp6U+oqz2Ut4Y8fcZRZQiRPKziR0nUZCiy
ZwBtjL6cR6mNprSGnx0J1TWeX6BxIPxCGW7I7ISWqamH9p3nQ5XXZ1M70VqB
SQ75BvN7bS8RuuldI/fPAvdVw9/mRbDokj1zF7pbO9uulqq707ZLUfauHWWD
ENTsX+/vEbJHk4y1+IzeuDgbMZNncOq63PizSgM1QOqf6IhtMVkFDXTOEhE2
z5a4ZpyPQJEXjK3BGIf6fVbRSMaiGXcTYFvGd+LIhAM7KjqtFa318MuiwY0Z
szVNnU2Ra9krFoSsSRHMQklj5fYHAuPlGyBj6+/Yv6EpOhKrEm2jSSVWKTPG
X/5SgMved5Fxem3TkxjgSa0OJYGeuH+wnTqO+39BnEjrmfsmcQajQBNnH97d
iZWbFAFlHAFwAMC08C/pAyRSlcP3BJNRn05CXagILNT1gDmLzNgMWPnjTipm
EiRztFEiKQia6M0UVnkb2kLDF3V+nVoNcK8SqTbSoEsaLb5fBEzFcpfvxRCK
JUl13KktV8NGb0TC7s7XiQAK8onhokeKjQygbEWd7UgegSORn8UV3c6qTIkO
m6l4hTLmlCA/TCkzDmkRwZi00l4RjgdLtjm7JvqpRVsN0QAzCK1CaVrBcSyy
qS3kcTAQj/clmP/R7uvM9VbvoexR7bvVtlW3TaTDPDDEG++SA/9LBrPSPFuc
NdD2Li2pRDaswRG6w60xu1GvyXLY3Y0iC/6R2RiZ2p7k+k95CoMkUIk5MzJD
A5SpwHGolRyqn/gaaZ+7AL2pBYuijw4IndVP73DchJwFOQk5nEraxPb3yyO8
qtLBfTce1X813lnS19RFCOkbytc9HRw7pjxSXsR1obvLJe7g5VXwhLmXnDwa
FHW9qwInWPZdGmb1ezcQSplfiRjp2m0pHYQXZ/xrDdpYKHyIoHbDXfDPbK4r
1YTi0/hlVqq2F45pLIQsjBHySAbR0HtS7br9+SaMzKxdyWZsWqArWJOzoFSw
EzW+MEbHwzpCExKVOFTtlG+NwCOJtHsbzrVJkagv2lF6Yu29C3m3sG9RXFk4
vwJhhmD0u9RGTxulxzTQOIPjnllIUe3U4GnJl3rUOr4Zq3+hfCoRZ8dG6X4n
ilu2mq7FktIZLYNBob2c3mL8GxqWZXRetB67Jt0VDQ5dZTaPCEf5dm/EoX7Y
nZy+ZJi3liwYAk/RMnQQXtA4kbTzd36ciG4qBHUNM/BM+k+y674g90HaCD8A
CVys6c4vQmTwxWq3fEjx3Nf/X8+mcd3xJqfNOB4LqhLKM39XrG1UEjKxV45I
vCKYJMM+I8YH5G8tKrlTK147IrCJQ27SEip8kx36duX4wk5ooHJ7Y3sTnkEe
+w6zBzOhURw/rhEJCVhezky0Ri+AxSudkhZ5plPZUyixA8VDBTwvKNiHbKOY
b2ixD8jS8eiG9NEIJW2bcX5rhWU+/PsJrfl8N8A81pCrKvkyTYNbIUvqaVBR
IlkVbwszdSEoDXS9S9FAy1aNh59TPbpYTlv68G0JnkvEIFsdoMgiXV80J3la
AcmP/MMTl1KOpwnkqA282ZuA74Ckdr/YcTuPy8jXv95uffkSmPB5hONJaMtU
SVY4QfCcxbya2WdAemtVgduUGqhcYwbnD5m0QT9XTq3kXRujho2TpmuFNb8j
MwBUJrdj8nCL63yPxD4esbsp45zKtTrkGfN8x/DC46kk1TgrlRs+N5cyRPmN
0fP6IgDekqh1nj9q1pif2MJid5E/28u66DxluRxeYwxYomYLIVD9devaTb/r
Vu7rZM9r2AZmk+OaC/gcPik9rbvLIdS5eJ+H9Y3GnPo1sK3Di1PQdHMgk0af
0SOQB0yU6cW/VV7z9orpHR7gz1VjvoSNIfYoYzbs0Zpa1A/hviPkii0sDXmi
1o0/+ORBHIdLFtxwvrmqBN7Sfk4oKkUKR/Rd0ShIRQ6iHB5vrgHO14vehdMY
QrqJW/TTUtrn7t8boUaRlMIowPoOWa5R9sJbNx+80lLG6wZz1AgYIdXPAESL
Txhf79o7MDUUN6yPXywpTB4fSLuoLOus8T5n3i7cmvbwCppyE0Cv8UhRMAVN
EAmPJFrHNpDsypM4WtnHQMYLwNkVcwpUf4Mk8JpBqfhqF3bxLlPQc4u9WPYV
HOiewTKucEXJYpJyWobrN6uJKwzCXAStKhgvex/YZ2EWOdMLfx4uvwKwYArE
aGTVtqMHpVvuozk31aAMChtwBbY4EfG8UpwvWEHlOBmYR64HVzZDorIn3mWb
6CpzJ10XI9mpNshuPV8j2zZyvEE8wG5J7YCL+W+zyciDC4kw/tlB3T9WZ+Ks
HKNjCVfcZhJWX5t7DyGVV9NEeVNHqKgIkfv49RI4aGWV//6OQhnB2x7OoO/h
ANlWsGwLDnEtWH2VAwmYYcB9sRma/SYic0k81ecuN+/nv+9uDea6w5Ms/jpu
tKpHDXonwodi45+lKY+lmoLSMiBuzYmYU++po7h83ZfOPvpFnPGsvrCbjD17
TSyyPsGQIYgd5kyvdyM/1LAcXgUzG7Fm4GLCy+sduiH3j8x2wPgT0FIkEifs
hU+TbLPsiuPKvbcDFH8f3yjrm7+fH8eArxvcGNSRIDMxxIytx91fHW8LQQ6f
/0k9dwofqSi1+WoQJ06ifau9GapY14mLMtxV3QsvPVfTpUs/rcJdPNLrG+8F
QxP8GEh+krMAVzUzjDM3qx+vwBf2V2aExJ76oNIFue3nOVhq5QuHtDNfAOI+
iqSuAd9ElEv4X/KtQho/3ewLC8A4kHBedsUYEVL2gjw8zG4tFctKZ5EB/Xwd
7rzC5vmcrdGEX63FKPtRZlv7VbyH2rk8fzdzKTW0DaDyzfkvssUKiAI97MMs
yOP5kwk+xEkEvEujFUoEKzKEaI7N5nWsPv/29jlg7hwnYlbRRYKlMaeHWoxw
h/Nvj3ZKJGLspqdAHOjoxO+PTM76SvNH5P9zH48qbc/Xseex055Z+Sw4c4V3
LRo9W7N7kgEID8Ak8v/o88PsF1bm1R01ladFIV6xvIM6jev/UvnNalbXS2le
SQy9BDPWXbtxAN9NuEBZx/hlc1pvCP5DARMdwBmYWbs8BS0fS5KM0PeTxFNY
BY1ZWaeuxHfUXn1O5m0JpFngdLfu+cpx7QrjLfpMSYXLuPkv14UsSd7JLrP6
tTWQFk2txALgjH+splSsw/ndGi6IbGPyVHSaH0Tjbzv3fbFoRjDwukZDt20k
5NCqjQ00RvfV3eOzPbUDbASik2pEHftYhP4gBwBe5+40Dq5d/VGjOQ4INWmJ
FjcVIe7nVOkPblJlcRW5ah4LGBRnNLiV7ODtTx4aiegJ6wzT6L99lLjjLOQz
xrvr/Vb0XF1XnRStXjnKt3ZmgzWrcCXsR91jlUWtCMkEFERuKZyjJcmm2jA+
5nfpnK2C4wCuu3z/MCJrW7XA8YB1AapGZNuLWpANYvB4z1OF0HbsTFHSqQiJ
Rjfba6YtaZ1U8BLsneMoYQuSaTgdxiqF/9AK1/z4rBkmtUBoPs2nQkaAaa7f
NFctEn3gIzjBtrfMqgmOqXPE05b1AP9v3ayNcZwgL4POyiA/zvc3k9qH3ghI
/yL2T5G+VZkOhNIjh7OZ2Y1rAS7R2o6qGNzXuVNMjuFCF0EJ0BN4y1XmDrvA
Gx1qpRPIdRsga7nlqTu4xxGMsjz8sH0u8gmpzaxMOHMPHsM7vBFlEqDiMcaI
RH7TP+nINI/gt/rwea3rJUSj7DAtY0da7I8awJsVLDrUZ6uzQL/QgmSSF5VK
yBBpd90mI0gtUgwpb8Iip6axKNSy1LgU/Lri5h2sm5P5KDBujEZ+Lc3Oygfg
2DkGQkQXg9MfUzth68Ncli8En2F42VRXUnesmG5zNfp5KOFfEXUNNRClc1Nn
kIF4+k/2ET9fJjBC3R15z5SfALH0d8h4iUPne8twC2ZWZXtfvqFNisfrMwnE
+2LDc7e0On2nfb5RtblbeO/vJAQQLmuw7QwCzMyZG2G3VD9BAYU/KAlFmhmi
6Kvjy6nvLU9M02Q2hCrv1hMgG+b+L9KqLGWmp8esIrRIFq7CQt+Sg1YaJRY3
KWL5LP2uh4NSft+UNgAriKIlGTI5wOxtODVJcCMShsjJWhvGMdzX3sK+lrYa
ae3zwIadL3bSdHREuBd0j51SA/Dxv8wS5lVub8ooL0Byi1JpXH+olpYJQs0U
eLmZfL3fsW5H4wE5DALa+39UfF3uz6dqUPiLp6+aaRfzDDs6QQKFTwcAryMC
RCanUEowVfYScmAUwEa+MfqQiSsmhdwAKzLAObmhAZIHSkJg/iucqANAA50W
e+0Ke+QyYv/unfEJdSCSFk3U8uY5vKDVYG6A6Q5okQ+nqANiyiEnJ3gdrIEA
fj1o/jtmcnMujI7uh6bdHeyPn4ZUiDIY0x1uobHjvRQYslw0vjLWtoUiXBeV
yvSzD2ecpnTqTc+U5nIqVjRL8UVE1abXKihgLNgF2nMN02/V3fNi49yXJznY
5zgdGVvnIBcM+McMpLWzTWQCAHs1bfqk+Ums9FcYIWgrsIYmWdq2YiPUcPee
4gJ98s49PIFgyxvlp15R82wANEw85jacuqvE9szZ0xY5WVyOH5asAHQsw2QI
1IfRlSb0icfUC4y8xIuOdT7JVRboEAIfflAIrWf9jCeHwlwAoWZvX2el0v3C
rMqeo4DZW6BuWmvZ8SQBtF4V/1/QvoZ4nLrgxesVjUeapzieoo8Ah1wDmNMp
lA4mKvLuTZinTC7pPyLwmWRdmSB81+afbgTWFxklHFwx7EPd2Xk6y9aHliS8
vWVoP1+MWB1W5rhaebpO+LWqT9ebqDH43f6Yob8dGizYKMxXR4vLTMYHs01Z
dEc8+Os7N1/Kbvm08r5VgmetGBoFD4eq6urp7CA/oXXBA/VImIflmxklsLoc
wDvPF4RzZb8WNchHznP3nvC/s+ACs4SrVGNLKv14B9JrVpRd/AIN1+0aTqrr
zVbDl5pqUx0r7pg52zSIgQjwELxGfpeKS0hwS2ERUTutIC+cYFHkyAVJGdTk
evZl0M7vXUzWK81cbnrN4eTzZBxKbhEWlR3j09GTR+yf3sfHxDKJrcF1DMbQ
1aaHfkQVhxKbuVXfyaQ5bZF6M7FBrByUFN89fEXGigaD1UfdHJOftsDy0cFk
j1SNhZMOTbuDJ3xfrjeeFsH8o0Z/Yy/OrKzP4brm3Qm1XSq/WsyTQw+mqH0M
nM/UmsUtzENZNIJwNQiz4PuCwqdnUthq8+5ck5G0TT34oINlyBiKZ9SUjXQo
3Gh7+7iSDXZ/22ztXqQzfBR/QPxO7m7k/yefB/sl9h7/1PBsmq65Znov4LNf
4CbGmPJId8vag78jeXf0q7SOqQuJLKFaAZEqbnME77PoA/J9kECViIhbA/7D
jnA+0h/nLOzww0rjd7uxGSOd+5d1341pE0mnIxuVJBb8nxmAVBC9VS4g+6Ic
qJMb2qrP9h/cTSZNHx9WPxTN63AFTRn13IYXtuLXgrhmzybhzJBIwOb6DT7X
LydtofC2PJbDeqq7/IYToeHUhcjBromxEeriqk5wlQtsfz0DzoCRY5a7KBSi
PsBQiq+AnqZMJfMqIGAYzWUBZ2j7qntz4fHR64Z0haH1JjC/vG8EMA9uemg1
/Yvl/y0sAhvBP/Kly8YlAsFxCaxrMBB2oUTbr60GtaoUuc/AoziX2skY+OdM
9avdSgAXyD3QPazXK2ZU8ZabgdYmYLHszVeNxKDASmwOc6m0r36daOMMEjgV
ECTm4zdupPrx160T7gCfsEyqnJVN5+D5W6ZH/LTyffTMiagouTa3tE2Y2sCt
JRdHmrjktQedCdprRgo6KyQapwKCPbneQPmJGH1aPoT8VdMzVZSKI30VKiTC
zD2JFQ8giBVxM0gLLhl7EHfPwXbF4l1aL4qTq2PJUSE1xIXXANsxKP6IlgJM
uuP0GdL18I6+YGaFlRKFff5H4dpWIO0bWyp+Y6UJGxr8VvbrCOUOtM19SPV1
y+vRGjt6UP3vIkOXz0sIiPah1ITNbCAsuKllE058uCBMmQAGZLqr1qvIXa2z
s8n6XfrFkBoN8bv3osPJtxMYyScbLvnUpmYCz4HhWG0AP3UZ5JmcV8b5/9nC
D+8LORDL8jIcKuFuHP+3I+2pgdjOwlPuBfZQGfCoI/K6wpwy1SOj0l4rHBEl
llOef4RI7C/wAVquh7N9ktW43gDIYWIGqKAe0giqHeV6QckJC7HO/qOhlZMy
IA3vZUeGh350ONSg8LFctFXtLYd12rUjMv22DsVyIhExL8nWmw6qn/JUv9r9
RuhLZA243YuTx3scD8k7JissAT4vPaN34LogVeDgLcuvkqY5F2vDCNrHEeSl
oRcJKePZ67/Z1ku9j0mIs6rQEcOkLKx9G2FPlf8VDk282P02jC0imR64edjD
D4Pq6hfo7ZSQ9227vc8IW7xmbOlL0hTrpdzyDISWwsuQzHL8HlqiCmRGjFSz
oOMBeJqIL6bokZlemnoUdYMVIZnrt9O1ZvLx0QkzB/j530xI0pQMWCkNIVQS
aYLXXyLhUfBX20M9GQ8UXR3QoG7bDafm0EkuBkfPCw3Jz3PBm7Sck5aYUwaW
Fv3d4xHk2++x6PV4V00RixB2zYrVGooSuV4l0cL0tD2fErB6Jiut7BLMyjBK
GIE9Xi24z8fL0XJ5qwlgCnu9r4WP5WTd/mR+4a5oKgVQ0k3t+oCVSt7mgyj/
G9yPEYCUGFtjv/STnCJuBa+oRhXAs6aeNaKy6Wy4zhhNQZ+I30XbNyGEiQk3
FrJS9Gppb9rzI100b6TGXZE6cSODfR7If9pgyVOMcsYksP3CtTkd7NPatwKv
AuNdGqQhBoG9Etk1NjMQ81hno2WXU8y2A+zZ90kUAGou9hEgqtVTzDAJXkqQ
Nh1IzbsZb+ORF12QmhcxyhQ9ZC390xD68+XxcA4uBS+KLCByPkAG1t22MhHb
211/2ili3wxRvBmhvgZ5FaH/tLdh5vx8VqCRGq9rT0L8Ihmm405szp9a4KGa
oJF0+NCbQWvmBtTYWpP/tq27ZuPVwCIcWwB5wadWaEYKD7ZMoSDfCIJGOkEK
liCnUUZNPfMoAsJH6OuFWvCEpG7ttJLgCYTjfIi/fULhMfJwXuXbY/Gibczx
TtvT6fz1TBKIoeUnEPReiFATmq97gYVfUgNqpkhD5bYCeHXsOeTqflrGvpJB
Y6hb1PKa8B7TrbYalDqIzHbhLjJs+uTXORYiP1VLu6Au9lH93qybwLsMQcJE
qOzKm/ZKUB90k+RdiylMnbz7ZaTmlJZOpaLLcaGfERnHQQKCyZHZEKZd03sS
R5p+XDD7WuNIZJNBOrJM7PnIJSRZPUCFIjZJlLT7L7WVMGocoAmONNnqqHRf
FGN6NIN7OcMyvQic8NZ3lr53TXCXkssD0ZV5rd2mHaTEiyHopsZ0CSid61ne
3t3oYpiNr+kNx0SP1DCUM7P1mdB+vH9ChqcPYSN44ruwlLkmf1IJ8tEwXHdj
QT9MT5RlJFWGj6HWRIdpb/C/lWNYr3OUFPvCop1YIDOmL3jtltNdA4HLIDVc
zptoYLdcyN6aH6gUYtp7BQb7wxD/4Yu5K+y1uTr9TTqOYraGdnwhIVALTALG
gLnQRqYoSsng4Zl2N9i5F+4vknlgHz5BmsXUaGeoBLhmOa7Rw/1M3LUwLqYq
FtireLOgzFCmhD74CN5Fu8GxBlktQnP1mKXuslwOBW88OkNo6M4ZM5Mpv30m
wdru1ftomuIZgSTqjM2EHTaXy0r7+b+q/J3rj7pQo2QE1EzbZT4E1uUiFUuc
vF7P0eDJtFeC8sID+Gie+CmPonyQ3zV10CoyRM581hfJrMYQPcuqF9jbo1pe
XBqCFps+x38sBhEcE5X8AV+/rVMxIMdNg1tTBW7CTOq7wKNW1WdzwqCrRT2V
fSmrPCvlqfFsaYstCyXX91dIE3BDfM9SEJJiEln+y5Dk2WSMXCXLx+b61PJs
pvIokdAERq/oxMEVM6BDm2bMQvebLSpxRK2ubY1rccXK7XeOWgCGk09ZG/d5
iIJbfTNqDM7Nw89arQ+QAo3zowiNTnTnnpfLTl4SXEG70OnGtimyLnRgk7vJ
lrhbmTVJgE145foq/9McCDxNLe8gM98ll4YzasM+arfRyLiwB0GimLX1YVho
yAaR3fI52jwFmoEbLIaKz7Bqb2NBLGC0zywj7cw6gPocLMc17om+o/aYzR5g
9wdjEWG5Exn5Pd7Ykm2wj30F+LcdERp9lansxp3Hh5UGLfgECXUDLVWk3cZH
gTBC6KlxFKoVAxB8vIqu2HRhhfavJq+e9XUE1Zr5WLkzrwWuDUNqLkXy5IVS
t66S7TnxuyNqGtLZcpArIBR7t/lL49DbtUSS01rPRlRoPmE+HfR6AffsPnoD
i/ioufk0+Z0vP2liWD/ji649ZkD+w81DgATKpiqW9P5y8YlT/bSVUbA0DYkB
oYMPS25F0p6qXFy9GW3lpukFI1mfiypte4XVSJuGykBcVO+K0fTVSnUXAhHl
rLQD/EuUMaC4XQp3YGb55LfjXSgWUjJCUr0Odsts6eL+yftVE21FasrX2eMj
NnyiNSsYpRy5MTqw+GlredmHjTYr5Ed7zyfFbQ5cgts4P+0Cv80991eGw+aI
2A7k7UQS0xA/yFxHmr5Y6Y1OyTV8Bg1GmLUzq3aN+o+qgdEXyTYHvdQx4yfI
AG4rrMfd+W5th2tsYFwdcIA5SxW7groNpE8Q7U2PpJuZvtNewNzuOj/mesee
HhBMTusqPAZar26DzApsnO8eJ6KL3HDKU+OdWYA5G6iMyjDHh//2dKwujzmF
9wYbUKDyxgCcRgvxhIImyU02mfzlLrNFf9eUKBD9rfZDXHawVWoL/Y2UD8tm
Oj6LCHUaig/DapPB+pCxT2law7MSnlMfxGT3GTei8BYP84R1hG+hK3FrQrk1
Eoynp+GPUpdxGlkzzjh8YPS2225my4VFvg4VpnAiVoxtaa6ap4XsbXVWClDe
ryMqOMtkjCy1PWn3+mvnoimv7cD04NHDTDCem069kPdkJ+rBLU7JPhx3bveU
TWk7J2FYMKFfLWFpmgjJdYcZddUI7xEyJcBEC7v4SfA8Sq9PEcTRZLIJW5tL
zLki/SCmP+tQLAIeh3Kj76QR14tLiJSkybm+iokAClIbIFFTklaweTq+tEJm
OpuEtGRJ3oYjk0l2qPLPqThetHSRjx7UTa4vno86iMJ8DX74LU5mQmE7cWrM
3MUmagHhUkvuVYNIbl8xq7Y/z/YY/NnSe8JtY5DI3710ZNBlN5Yc5xnlUQMy
gywQC5j/ep599nBK0LF6AMbqkqXaGaDaTm4CDbIMi2XX0wfyqbZtQo9RQJvT
cH3yyAhcjHF/qIPykD8UG1qaMZLzEB/aXvshQpLTYshi7tPa4mNX+E/dVD0d
LXI42QArulXr0QMRVbEiAlXChDPpeUKBSQ6gNhQX9YNH/iUTNUDq8zsqMCNl
kYQAP7wrz7Yoapbyu3YDvhFTwqE+rIEKT4Apz2/MAmiSwjgMnZQutIb9W+1E
ZGK7UqX+OpCOd9bGKbI7+y1U8XiksqLl3M99ssTZYnbrHkI2b3SVMtHdXhod
MlsFCU6zMEAM9BJIfQ5lPcAzs8WN8ZbEqhwYIYj4ExfBDh+wGWWpt++IjS0E
CioEVXd/L8zMGL0skM4oGqUxwWDqRWsSbOZt2QLueUFYcwi5z0psBSlr48Hu
yN7I/mtl7z/IF0yZMcxv6eaUEyS6QR/q5DNKzjtiGo7M08GHD/sdAhYYjt0F
v7LOghw4jIn8TdYK7UZvDlEA0adKi9OIe4SWCqOrznvVWTFjUAL4mbefYWJ3
HCeUnpnjagEPXUh9UslS8cqz6VdJGsYPBXqJ4BeIYLamzLYmPzo1V/oS5jO1
a194NmJVX89kgo1vIj9d1Ox/yKMiRropyuQaqk94MYws0YwMOHbMUfbP7oer
Ok56iNHw0xPn1Fl9eFmesGqpX4to47dag10NkUlSUhVzIZUYuBgF/UG1LDwS
QUcqASzgiDsMzGFDm/MDgAnp0zIUbk53lim4lDST63rlObjpj/PfX0ZDmPib
9GtBZYeHGTxWxffw2rzBUT/4sSi24kcb6svLmeHftGXQWIeYGTQ5+6SwbEM9
0ocGq1egscP/PZGu3uXRkm2kV3vmYV9LXbMiwW2OmR1UT36Jgz4fEvEzzeFO
VEIdjeaO0CRBxc2JHzmlxi3AMd8EqARpGNOC4RDixMkYZtK/GTwIzFy8JaRM
BAyVEdf9TevReCPSyZM5DY3IN6TQD3yWvClkOTZ2hUGoE6yByV+iRGlgEed4
WSl47vxisDRHXVEIJh+bRvbH1tb4WooQGfjKU9B9JeJMGYYqirW26Q/eYZPL
waEp7wdPbClByo1oNIRnnuO3Dx8gXYFeFhzr0o+sbZrTpJ6sAYs4C02ILNCw
tzOsgKyZ5Kt86GOqJs1TOOyvvB5kimC4uv3Y3M2t7PVqTuXnFoZu46vkxylD
PoZadUJooElOQi0T5dz+khB7L8J1lnDG5kNFBRSjGVDpPWtbzUc965PZ1ziv
cRlAjpK780FDKGgchRAKPgfVSkPygWb8+Y/vqQEeCo6pBmSPY2ACT/fJEWKA
y3+JuNpMQaC/eFiN6oSJEmSUeQ/Gsgu2fTqgGqqJPp4Vy9HqDhGKMv4DZGgi
hXIDJYRnh+SGguotgj91M1yFuYLdS0G/CtLfK6OIAVBUlDQhnMFoDQ+P0kx8
Bzv+TNaH2xkOte8PEr604yaQvbNGxgUYuQsM/5zhIvhhDh9wlXwnNiQWAiDa
J6tvP3fgZC9r5WQg/0J6NQQX08FW9j5VG2c0F7UrD9I2JlfwHKZChtJcJWTd
83Ti4LnJVfIr9KVZj5i17cGMefgIoxco5r+6f4y544m81J1JuhLGVamLnA5o
4yCrfHkd+B0ooBNYD2WOu9B9ZZ9T4eKMVbgLzXe3LrpMRF/C+K2VqipKV6gg
4TttkPI/3q0KGnPgEEsOmL6pJSZocU5c96ZH92PtGkLU/ODTtrztwLTJrDt0
l3ByEgylKKHVwf5NH2PY5/9PW0DDmplB1glXr6yXLi2VhuujpHfAolJiNR2T
D2CQ32PdWmr53fqoAhGXh7uC0lts9BzRFrRM08WoLW9/6FaHib95QFbXpkLr
ol67y5vMt5NKwdHi+2GeqvTU/wn8XFvWEe3tHv9hm1xPhVtpZH8zw21YHAkB
OlwlJOKGeHt/+4C8xoNrDDsxvFwnOZD8Pc8VeYOPfMI/zxt5G6KiJhDsoSW6
EYzcD6C5J+2ixbuHGg0D9bHH4KX3tNbkPz0MGz5ZtUPekQZrbzGdeCxWlm1t
r+MqYrOnQOgHL8sYKIw90aTYVl8WlgYWGJ971LZVaGVlp0RMTN/YOUgCBcTm
oQeQb2SuSRddHuvRheUO7pIQBgtDeRgOh6VxVyPqwogDxMihh/Eh1X508g0d
lJ1OcgGsjr1AO445srkn+uUCGnwxnN7XQVKRD5u6LimCAksoXvkQwgdelFxN
eJuy6o++c7+W9CCzTJ1471n7Wg/Xou/POjKyIDjwf7JPMj544XJNHEHDVQo8
AdEkZmwKCrf7Q2V40PxHsx5LPts1sCqlBdvBW8nUldpAhi/iALBwgmTtzy9c
DLhfu/5Xi+96BiedABhzZGQXMaIr5PZ5qOcdbia9rjbmi58+y93dMuOIs93U
jYETW9gk5aFi+UZFrXiz/nS1Jg39LwVUPnsINBO/4bVxYBJHC4kjL+CHTW34
4VojfFsnTxFn6e29D1kuTrYox99m7d0mEMj+8gKm7P3IBkBUgWRszgwDKOcs
daJRhv9qoigfdTBfqwWyVmyUzoUSNlxsRAmZl23c7m98k2GbQ46YgDbk+EPc
WYnktB7O2LYlAM1B9nLUI1A9vPvZEoa8lySvhOANR4Nnni8V/7/OQEBvvgiL
6gOh7AMl4Zhgd7fxGpYFgoT3HprDQ3/CtgYAhNuiLztHfPlQzigSGBZeXJ38
khibsqqs2PZkpXo63WUd7EvbgK4q/KoLUjFVix4GR4lOpoLsKoY1d3bqksrq
yKK3aFQ2auxo/t3VQzkNgq4pE4f83Me1ujJ2JkasylmUHMAOTBqhRbCF4h5J
844gDpAc5V0cR86WUoUvvnEF/DLt5VcDlBodlXF7n3V3e7hgChfDwXggfvec
BDEnWh5yapzTnhWOx30eRmiqJSI9YPAKyrfhLvXUcy/2J4/uI0UNT/5x7vyy
VJ5G9oyj6VrtQh8Zg56SKMoak6qRV5GVkUFE/1W5A/Oopg67jhpD4i/Lhu3J
tU2HF9C3Wd+URLwGOpmKIcprW85hIPTzJXaOiE0TuKLmQo4avC6qAbVkJJhw
eP0KY+ktEoQTZSHDmnqisJu5LfP5cYWflDB9h8IF0ZULWEytRZNsXo1PRKIf
6JrQj6x3QSLTNvFUo7seA3oxSle/7O8AE4OsNF8yf9zA/NG5YY6onKxNixMx
7GBl8I/EDwf9CQV4ssn1O1C0vfb/AlYzGWO93Sohr7/yJNhbgd4+NZYXZSuW
RJCsaNVw3vqFCGWVXmIg33KIbvM6m/jZ+8GmMyQdK4R6pRHOK9dvp2UH8Bik
mSMps+SeGuzeRsTNKA2TB7tlRJaeumfBziUjCflQY0kdqE+eu+zmOzGdRHRa
lEqKkSbJSqk0CCnn4Uafm5ot4G1/pMRrrVfw4BoddSlIKlwvHSflTgA5vQIq
NCmByoF1nmKcydDZZHLm22QwDzD+WabDH70ItIObRMMPTZhCvT+gb/AkD0N6
L82dReGz7NdeLIAVS9G66vyBMuVj16xxd0Ch6ixTc+8UsyY3Q0PfGzIqJVHY
x23BqUxXNNRbSls6mRX9zIMoPAX4vD9Xe6gxX7UcqlWTrPJKED8++gYF0DUn
wjO6n2GiUFUc4ueQ6gA/GHGRjlDQ0rSgJ9C9XFzD6NWw0nLODQiD2CtupSG8
jeM6zVbMe0y4Uz3vFq/JKNL7dpqHxi6AuLenMcR43VdEpF4pIq2LBt1tI+g1
/EAONO9DbPUmi45JI0f1C6eIapD9/qCKQkA4jqa5TD0iTz9ucbxmyRwAWURm
k4u0/LrqhxOq65E0kiFJp41pg/T5rdATsxs5yrmR91H5nXgGK7dLyrbPsPN4
Y/ufEzN6niiMxzWVfTU7ffpysq2PTOqFF9mPPmwdBTx9/Y3ITuU4qDGPBus6
0RnIjZ5Oj8716KHFxRR04+degfv+mZq0xVEsXrApZV7J6lOg+9fIcyxnY6Mk
IpGmXHSTLCNph2iSdq11ac4PQ2Fxy5SCWGJcT2blc9fuHayH7QAyFXZrOLyP
+cjsEZyyQj6gDLraK06xjLaYRSiQyVT6peK3jiike3EJ/644iuUXYW+dPWrB
kbepI66I5BLPJgd5ZGksIRA6CuDkMW4FKWvmK5vqVBi4ky0NqGMRpTr6CGwD
6pQJjwUeqOtBTbwKQsVMTW5OxSqVxFck62E4tVymxYjnokEbypo/i5mtPSrX
KbCAi2Ie962RWVrfPQ6HeJReIJ43wM6iCsnEmdv9IpgN++ZLKsMWwx+/j6ip
ahY4KZDP19szvSc9IqnU6wSeD+n3gc9oho9z54RhcwYJoiiwvLmblhITwdo1
5ClsYjKLolPaj+Q6we9AIevEFiPqyvBbAPsoJFM/hyDUeo7DEmoMf+JNXBYe
F0Ssp12SyBLGEu0SomvYXmmtQrxKjfOwSy57c5MHUXnEd1cEYBspGvjrx4Qm
zAm574QfmMzUEWX5kEn9OnjUHqpJGyIAB1GoXxvvxxVYIfGqEhkiY/q9lktJ
WKmZ3by9BZ4O/d75/qN2wxBFotAYQmSJkDW/HNmOiYNvrWOqcJgjbHU0nTKo
0fraRQ5pLvMovBDCHqn80+DTPFk3wnLlN0ItziqH4tlYPHdY2Ms12w+ADZWk
kv9j/s/vD3ADHRpMH5gGfuOV3X89iYEsqntIdSrfEVZMXWH51eA2idDFX3b8
CgRRHa3OPCBrXW4mTPI1JvFf/wOA3En5ozGO9VSC8MFE9535ks32TPa0gctB
ZxfLqbgwS/J7EBtMNXmMTGHPPozuS7OHUm6rlUCj+EQfDG6vuhzkbV8N8+6u
uiFacESSEWPuJRshoP6bZkzv4t2ND0bY/2b4SZdQ3H9icv5QdGOyXsINdmD1
WV/Ktcv/T5uHzofecMdmwzSrw5JxbL11p76lY9O+oSTK8FYtGZPWFro1+QA+
EmvuhnR/Zn5UKeIezTuy7HZVB21KLfw4yZfRVrs5vGo3i3Bfx74bcRac+NuC
s2L1FF9Y3j8SrmEI5xmWRgxXrCCsUVBndYCAZaAgbfdM8mJsxvNXEG01HtRE
+SIY/Fev4jdy4mJsQ05oEvqMrB9jS/84t0phpYOaj8vRpDgHtno4GNv6gH9E
A1SCBXY1co+aBR+vWY0L+G/OsZEvbtCCpkUgjZwhczyuteNzzh1weej29/G2
frQAA8fcZ8wclfusY5m3GCnpC6TeiGN8I1De0gIr5pZO3DpuDJe4K9/iy2Hh
3IuAHw4UveH2+0zr46O3MHQF+pRse+4DeI8UyIQYO9TzbEYoXTkMkakeDG4g
AHUodtIbyd9VSk4n0DjFnjcpiwcmfJTfNwoyGEHVKdAulqokqayBhirO7GnT
E+oqEsIgq+m+7OIEofa0nUNLB1N+yTs45QGVZj/RqUJED0Dv5zH9CO3nI3t8
UyIwkTZrR2mb6QyhkwmYHLlLiGaJ6fWpyJrHJEwRptq1jjGIW2hU/RZg05n3
r2DCXekPg7hm3F9WpRd4thRUSE76pkyN/U7ZwbJaM5E8cAeNw9cYfGkZbsgq
N9+YFY7L9Moume+0Vzk+qKHJZRwz09yAHG/1/5DedPV3Xtu52MNthY9opIIK
pBFqj9xUBF0WbZgh9d+Jc6nGt4FylfpvpDgqhID1ABVfl8dXCx4wabgWjKjl
fN4ssMzMkQ/uUkL4547u19T4HA8w4kHnyd5Hgw+kDNaZ1cZ4E0MypZsrKVQB
hn/orXs8H6yi0/zqzar0DRa3a62opanCKx3EsUZv0sqQ3JasEYxB76+IXf5F
9B41QPGhQV+Cl4Ex/erSkzkQc7lqsSqfZJqySno7hmsWgak6Gtw7irZtgK8n
hGJ+ozMdqKvbHhzn1/ebHYYqS2k8ES8Hg5STiuQI9iGqi4FjkoxsO6rTGr8h
8+vcLhMbRn7lT0sTwY0KbsaXS/PuaGwO537Bgfne2yNWw8WiarHvG0VPqSQP
R+MH20L4I7lBo0Wi4ipUR/ossmQE4/ygspPmsznF5yyeF5Bcwq6s6Jg8eQrY
+Kqyju8WZ9ithwBDsY45XD8fDKV5Hfa+Rc/QRGPnbKZSJhPabO+h114b4CYg
zpK7lpI+Xg2PIfZ82bR7GnVZlvygBSZagN5lnxfpxzyZN/1DvLn7cc+GONfo
l807otakyuNqYDOUTiyjmemQAhnqy0vFr3i2VuG+J0Xy7lZLg3J/J5FYvpWZ
0tIQ/MSPmB2pQOyf9ZTZ6/4w+x9NyXf2wjqC5p0F8F/x92N9a/67L94tG1Na
WVFpzm430MCOj3B2zJpJNvprSoq7n0OJPE96Cn1tHRZ5mqzrN6AyyKI4aXD/
jo6QHH0hKeLh8l7Tu386I//YxYBMG3RRpj3zyW8JBdqALVrIB7Isf2lnw8fc
FjRffIebQJFnWkrHnArPaJDU8SBD36nsipgQuTPbCffM8catXxjt7jbauy70
DuGOPa4Dk6xRFSMcAqD75iaUHAQwY+ao6Qqk9cIIJ/mQpLTygkdI6VS/94LB
pWnyFlIYZxFb1HDWDXMCfHxxv/rZCWFJDcU1uSiEn4WDfry1sRA9AJe/tf2l
94iocml1nedJGGmx9NMbm2xlaq7U8yQVWh5qfdi34C1/FL1nVhlhwirEOt3y
SvOaZfE/NxF5cTy64W3hTH0XGlJt/Nrr9jyTO7H+W9OEnf5Dc9G5Dab8Ttvy
DcoesWZXp3UAeybQc0IyRtPXrbEnZUjYe0jXOmqwLnKTdLliOKwd9DR/QgUJ
DRw328A27yHFmTScoFVF6AnT6jlyXTQ3pVI0E8Ga+UP29OqbN40xs8EcmuNh
XspoeloPvRFZlFQ/xOxnfju3XaxfAaKM72Xj436QhmSV/n5Qu3i6TmTc4IB0
VNd9NlcuqVD9hdJdaykbnJSj1DdUeacaMffQzrpd7mKCKSNCVrVKtW/PPU+6
btDleQ3r9hLmXjBwoG95aRU4pZOUpK9N9mT0yPeJqgrohPUKVTGstB4Fv9sO
h+mbq+4UHjY5NEf9USSk7Iyw+j2sf5Qc0qkfN6tirzAKPoDeF5rA762Yw0J7
j79bzSxfCmVjG0GVYZnT8YMlXxV6AQ054Ys+Bp1mq38ThmfLT/6z0/vwmBCS
s+zJqmJc58cgopfxIorBbQ16z2jJP1p+JbRFUdk+v72pMtvF5PsO0VGDZnId
UvkIJRykm09UO//qxeAXt51FVlejqoRbm970zzyAtOLKkordrnxIdvsFsu1I
2qUzdfjdUaAtCzuB0C7NTbk2SlcoBC2HHrwKZ3wOxa8jwxIv9YpqQAIVlmkv
aJBT8OFuCP9F48nD3cc3F1FGWtapF3Ehi6CQ3DZaHE17fXCTsVk7/2fp/8LZ
Xr3pnjb8oLSHL6dVkR7YQauPnd03AXUYuUyzPK/yB23/asTh8Ejfpkuz3IQ+
yyY+zcnc3QlJY9fE/nqVvQtZGihisdpkIRnRnEe/NEftIOipt10FyCmNbeVp
PKwt4qM+ZkMYrfxRfAw97qXzBFn/c8+x1mv0U3G8/NPSptbqLYPT4O8i4QI0
CvHvuOnRggI3npklR/aHts1PabByvmG8Z559S74zwfDlQw47rggsRpHHl3R0
NcAJhquBj+KeEaoiGWy0k8mbjMFmplJI23cICJ4ZMtE/XGvrSsYPPMitsZ3y
Ugup/k12G8G2CVfXbTZCFa1JT1a82maZs/UUmj9yCq81eryA7pqB42bZI1fj
EOFt9AgdaImxVG/RSi4IklQBkVTYVKNLbfV8bQBZ0Ui+yqmRepyqEdZom3B4
D9XIONXmeJsdxkz0wcCclw9iXoh0KtXSCcCkmhBjw+BDTkE6OXoCvapMI3tT
Mq/DTQDMsSATxxw9pTVFqHxT7mXYi49FyQ2+s6CCj/hLyhy3m/qbhqWVbbRi
OzIceLqeSbuNQxZ2Af/OTmE7XfpOHqp/OAjr8/fUh6sniSX4FoKW8zQbFI7P
x1B4oQ3v54vpGtWPLotgk4VUowJ/ac3ffRg2MMiLxgM/C3vdId+D/aMngf9/
mbxv4pwyOb1aPbxYdtW5p3gLwn6OcX1sqUCDtjo+4SpWa36yjFa1DqSZuY6U
+wE1CKYNQspqb4RKHF5UYr4TV8PyEBkfS6n4pfD2JQcngoUoM7O/Nx6SfMEX
j1ZUwnlq5kAO5o0HED1ReZ4QtbLzFiMTYfncsD2try5FpN4PuXUEZXkgWK6v
drXpVnelz3T4KFsqCyTqcxQ082dP0m7vNXuZI5q+lTAan9gQ8EOlgdQdRWBo
VUhUpehJULupp9EkO1/pR7R69Anprl/4v2aar/vaPCMHSDEhCbIkKn4LODPp
qylYmV33BsKb1AikL79ZPRFsC3DRrxVnrOifnty5B0cgp6D1MrX5rprsIDOj
qd3mY5ZNtZCIdLbTCtansDARQoJd4lnitUqf02Fw88M1LPOqIrh1L8qrCrRf
juZl0qssjH/S4rRUSzqczdzuov2GgCy+kxjj2lmiskE78+NSpFKiJpE0ruEk
IuhX+ElpkZqHXIXbPuRIUlYmhcTejf5DYK1kwMWcRUD/4Mi5d4IthA6/ZL1w
Gbb+06LOpBbXCbc9ll1XzQQBnGzOTjPf1Pwlq2TmG+llLQeocWk+zYA0VtLC
J26//aqOW3bBbA6iFXYw92qCLG05TFMi2+uP7d4r4lYajIDeU3KC5Xlc+j3Q
H14HWzVu/Q4PtpDJ+T6HB79xaBNRf5d4A8C8eVKim5jlEmCA0KwKQnmMQd96
q3PYXCHyIfqQ1SiRqLifapLtM8sP9BgSZaRMRICSe/ejLgdM3ZauMDmRDx23
0H5VdeBNcgJAp3gm0uaPVRsPRmNvBPdandofmkfLtL043eTC/VN8xRsDQ8An
7CsFrEl7hN+pVMoFda1Psq6oVayf3TFushOYcIkngsipd4X6X8shSybPdFSp
hbEnYt3OVwzvOv5st5mksdm+Rky2zofsF7pON96liZlkE6VtY3vVvP5ktyhI
JmRkxr/azP3zoVlt2NFbS7Q1GMMG+OeUv/xsiEYtTC+V08Si1Mn8f3kqLUrJ
r665goF4VNbts18gtfxCsR6VVKYOnwQxh8kKaHsAqxIminXGCHTiwWPK3G4A
RI75yARu4w12acYyLVeyjR80M9DMYVEWmFu57dSd2t+GPH1L8ClHO+TwwOY1
Byod9DfachyrTZ9zu9HnbF+I/SIY/HtlXO/59deUGw/8rp9c/J2hwBYst/76
WcoIKIH1+GzGV+QYJMkC5Jo+59SdezJSpi8InMxak7anoEL1V319M50smQE5
N+YFBzCqwbkoAFHeLdo2iG+C0DLgiRbcnxR/ST0KXmAjNMLp5V4QbxaOutUx
KM+TTXhcE8oI7kSEgCvCHMe4X17VPArvrbQEQ5Vrsb+nGeWL1WmM0HzopL/I
KzCw7SujVWJyfR9u8qKf+e9d08mQbqp9s7ufJUzfltKTqx+CEIJmq0jyw04y
/Zm3BGSQ5Qzb++toQGTVDXZP6lWBV4xqzV8E9yp4g628olgfth7JIrB7wnnM
EihvUNjdsQeSaFgSaT0E6vFVGSmEANM3mEP99cdyGTUOrY4har9XiDNIMANi
wYjNAR8F4lAnjvFnp32jWo2YnZlNUIeMQMk4B1Zs3WKQC27YJYE9fOQuTu++
dp25lklfBSojoq3gIRc13mtcr5AK5QmGpSSFSYaUSePbM8ePlQEojMVfoc9c
X6UhTc4WGgkWdX8/18Sgvh71BipM7kKq3Um7twuTXScLQ/zSAJddtX3A0zfu
81BCBsOPaHG3gpLfyPU7m2F6ShBaCuFTGa3y2O2QIIKNqllMGJ3sZEyCvIaO
pNMgjoTWxcFYGNkpAPm3QD1pDtY6os9XAjt8gPp/Z8toB4NT8/Ittt9mVnMP
lK4HOKJ4SjDkeCySBtbylciE20M5vTD3vayx+WOVkQYGOVKSDLVMxDHE38q5
upqInDkPcOJIdsy9uQnVcJZYZRIpdw6wlBWgheIgdTeREiJQYaWXb4bIHSaD
eAHVerqDmO6qqPHzNYpozto7bwC6PW/YgPT2xrlIqrE6KXmnPz3HtNW6DuDh
aDMJR7N3vEiLWn4K6Br8kzDxzigaoTh8llMnWTNHF6TbIzmOg5kZqQPzKVCS
KlNcgwa8K10wcQYSibelIjVnPSKyFSeD2h1NoHUgnmlZvXJoHr4PwgMz7nXe
VfL9t6O20N7AHA+kHNeFZiOFtu4fTItlgttfXbVKlqA07E90coMT2meZ49K7
a7TSZwcc1GRIXtQdqPAGmRbvHJW/jFlU1sl+Q/ttZvPhyeGQNpkfbAZRshV5
CpNZlNHrv5JklTbZ5BYHI0djKmJWZhF6B99yRbsaffcQpgjpOvuS8v5mpXHp
nu72SuWlLVHWsdTCYrUUJtBIEaMIF4iek4tbxM9Uw3B8MZ6erRKvGnQlXgDS
KNpnZ+haWQupTS9uiq7sCc6iH4RoBCM/zUI4m03FQNV1quSjuJLGUBrLhFwH
lDyXDLQY/bmA0v2ubF4QfTjHV6Wt5lFcm9PxqwVOmoEmq36z4574BNKnjD7B
+DuUPg/sSkOw28D+xUnfyi52xMXImUITpanrkw2iUYna1XfL7upfi4puym8E
YZ7IGN4fMlDR/d/bhY2PLY1xfFTvQVg+fH3gB2cGVihJ+jpPEpAJ3x8FT5Pb
Ri9RQLQVpaW4+UyNDStv8auKwt0HrUeKpFBFT2CCKPB1a87UY8bmKXsPikPW
5SDkoaA0tpdCwzPnTyGr+d849J2BKLdUBvJrkrA+JyF87/xNPZOjOGnvNbtQ
FqJtFApvHmvahifRPGxb+9pnbJuJDDerDzNsqkKvIJUakRFU+UnOMWmXCX17
9rTitUrVYeahCc02IDZfcMUvxAmwU1ErooiRcFH/qXVPNaVgidGo9hrj4GW+
tuqv3jA4xT0yDJdtm2u+Y21lVkVLFAWcSLLeU32eJNvTgvBN1Tz+ln2vpK3E
C/0kiKTEguxZEXj+lHRs7w6S4G+AQDP7apikyQ4Aj5apfBkrtvUTj6Y7QFUd
B9HzyS8/rdny9WTwCFRaAnZmXXOfL7NS/XbFZ5kVvOg4+28PHSax6pV3kdcE
+gTViHoQbQ8FfWBN0htOZXCcAVai2MJ4pidSapMauABKRLUczP1O8nRpxCOX
XrVQ7ncznYcmMthrYoD1yRVbkB3pTxL9auD6ziyRpup+NbveYdO3jdBkoZq5
jdPAwSVqIU22ONAXXX8myf63RLkZwIlj+HbpRmVTh+jtws0VC3mR4txgLVxq
NNtX7f7oU6/pRWWDnGMqKPOE41JfaJtBlTq+jPTZNZluBadoF0i2688MC+XO
U1rGWlHj/EPjf4hbqH2xOkoNuE6YC4oUy7T6F2iLlv82zn0AmF0Ij2e13VgG
/+i6fLpK3/v82xV3G4GotTqPgwQYR0AoKkRDF1rRdmebpOkNsd4Cu7+NPio/
+dBvZ+c5pbmj7uxorZfGkgSnkgl9V7nKwnSvif/d7JAlIsiYixmEVAN5kDAb
rpgDUArHVMomYOVQnB876XE/2n6cZ2RDe2QJpD0skVW7iJJvlSmL8btdqXec
oetlQBloWvg0fJZvea4NvG2/gSvJmXc/i+BXpH7LyM+dymZ+rOKzXRTmUi9E
4AvK3ZF7uH0c0wOgc/ymitGndaKPqBIdIeUDy1kkvb8N1FTDZqFpzqIFzSLK
0+VI3YkAkDDfbeeawt/m01i/fRSm2cJzO3qNbaIOrTe1cwIV2CyVVtFh2ukm
wCYCaUQyW4ZP0v+8++9v/pSmPhRQhGuwuAGuCMNL1EqCmQUF+BvOH4gkPjkL
XtJsHaGY6aFbxRy0s95Zpxb9fVycXvDAaUw7dqos1MZG1eBDjyDJS4UlhCah
r8wnJksSFEOc0sczVCqv2aotGUtX5DIV7MaNoo4SqfGh+xj2Qu4ZOuNLI3hA
OT+Mgu91a45KrxuSp87HGhgJCtaWbJvNyNAU1iIqFSE9elI1x1DyhijdzUNU
J8KaAdEz1zuiTiOdl1zESpdHiXvXeic9JtkXwsAZJHftbP+TPuHebDnfNzNS
LBXAggFfqmYdXlQR1xCviapKn4p0HCE24ElgCcJIgYLhaUWs4DE6P5Oopv3m
bijlSoB+geKhSvEdzmGnQ6z9j7l34joOgs7QLfc7DFRrn7ttV68jWxtPb/2b
j895GIcmhfIeX/CsaTXJ10A37NLF9xvziuZH7g7+UKgpluV7XRHI39fyo4Ju
sqYtgD7vMm5ItOGDDw/Vwy1lxGvvI9duTqEsWBrxu8JLB9qK4+7IpmPRYzv7
emMpy5/oKmsiucJnPUrEV9mPdHb46oGKm93w6uemi0jE/5XKMdrvbBrL+cbY
fQDrE0BdyVGrFENjhmwusbzBGDsSVDTms2hDxzOFg1mndrt0irQMWLAEVU3X
FLtn9qrDZJuImjDKSvtf/yBSW9iJVj2vfbP884m+QpDMEelV2Mo+3WXkfJui
+j41EORfwcJNFFq4HJnTheZwgU9zgo3bFEOTKjG/LpYauZ+TO5MaqJI/z3sn
5kosu3FKL6Jug85Ce4c/+CBBzz3/ubIqgP4lFbAcZGbwRgtZYQvEowIKtNLd
oVOeJY9E3BcVlLOFpVui9OFHqakzoIbll7BW8BmzhDMb0TmAFOr3/5hsMw03
ilq9RnKiFKu0q2qEgM3HjQyy1KKRkJ6e2kn/7tvt6sYB1GlGW36CDOWda0NP
BNojzoq3mlrWOCIKh+0QvZRTGhN44iksJ68wY8pLIvxyYIEE3CYm5JsyaOpF
yaYllirTWTE1E79Vp3QHcWrqwwjgAEV4EKHPgL6WE2kBDYr+XMU4Ypz3XyH3
zjW8l36GxHxDeTk8KgN5yviTEK6uvOmomYngmszbRJCRkUqlStrdvOHcu7yT
6Pvzmpmhy3kJvBmm/Bs9T9mTpDbovSVXbUHyb46pkG8diCgqavSJM8zqRzKQ
jeS7NRtpBmSNcm3nyaZXBwKNqb9/zCK3OIPgpy4Z8VZ6Z0QYvNohXtuj52pQ
a0yUHRRJBEv3+uMdDbHs2DW+U/7/EeBH8aVuXp8ZMwHXYx9YH16iFJE8pljO
nLiosez2Tauykttp7Ne/5ULAMEvKsdcOxKrhzik7/WrleA4E4AFihZcWNBSE
813bqHiIVY8S3PHoeqOVsoXfFIruHzNXRrJw72DiHFoydWuA0TG4X7zTfpsE
il3G2mV6j1GIjejNmvhBKCNS+oKOB/7Y+NeauCbbk75i9ztdyrfHcGDJuIIy
0RKZVqnedROhBc78X3uv8xLK5PXT2fGHN8ykm5XrVszYeyHDkUNXLi7h8nDC
xaLeMhN9OQf3Q4uWjgSjtqcfYrd9eqSa9UsTlf+nKp4bI4zmVLPpS1j+HG1z
Q/Mfseyx5o6bpesr5ubVV8/cD5Zpzy5h0zYC13BBSdk/yHPVPt37glIIA6rF
yUhijPbLnl89wnrfiN5AOF8iAkwKaNQsgAbnWqp/V5mxtwAxWiSCypob63aH
ddtwgZ+0/4nGAi3qncHFf1NstRjFVdfC5DfyB+00eFciACjsXqvC3AgH3GZQ
Mzc+SbvWvcULInOGUUqAOmfg5dn7Ordc5qYXGEQ5e8KlkzTSZwuY88ej0ILc
EBu6iVUMfanwpDJy0Qv3n+rN+KlBYarj6Dqz+oS7j0OjLxpuykJcvcCMPzKt
0HoUcuEMb2epq3hQhL7AfvwsBEIzts3KydsfhbRPlpLvlxMox/LPUJHhoE7T
RL0M3DOf2hRIEKAHFMpqU0jOc5FDpbkJudBDWT1b5xPj/6en9L5TX7vhqORe
CZZbz1Q8oVRabwxs3geo90TcGwCwf+FcXs1nvQFvEaUav0x6qoNNm/bF5ZOM
xHypQ7D2sP33tgHDipzbP1lkTx7aD0L+TmZK8ZJk893ytcrK1BHzaho4i37b
EBCDUPaHAqQoZ4qwx5vfHmVQErWihrpDlMRrdpR6vjnMSOh5G+X0YBi6Gzl2
3rFIgpuSQJREltITP4wLiPg+7AzbG3M4pLD8U36S7AQbj76kCAbqjeB9Cfw4
zCN+SS2rM6ZcHRSROlHh4oTPIIgTk4wpFh+KuJafuqBjx0rvOjw1HMQ5gX+m
aHnS2YvwUoiZj3UggqrJtZdOxxyE2GaiOEanCGDTf+4cYloetsNA8W5dz4Zw
3hb1t4K01b8XRxgihR9dVyfRalzg5b3yNbWJ4aL/qfrrMnskSYlSyeuujdAm
S7Q8XvdK+YEFnmfXcimP23ER/Kt6zgYwFC97SqOKouYzLxmw9OGc+uCbnK3d
QbXke22TkF17wrxPZOZgFDCLLSLekJ6JszX0TkTlulrZHvpDIrESlJeSSS/v
q/bkUu/IguasN/DL0WMWQ9TcL9P+Mqd7BtIqP8BbKoMc/75ZS9x8u3OcR6Bb
Xy/2oXETIGhTnT0/coBdxTkOW2xlg4JHV5vywdDcd+49OCvdLbh7qhxzWdQC
1eZtn1fk7y+v8x2yf7mIw9P9y6M1pQv8ji+PqFWahfCqk/j913yqOtb/8PFC
3P9BbgfkqGLacM86BiLkFpZfFJH3JK2tT44uvYSJOnlffpyetQHd4S+0aPcz
4ZMJL9XHSTixstKSxVWKvokVvn4FcfYIAl6wLfN2NeWPOPFhbCruxzkfW5kA
ds3mbnEpI9Yir3Vn9h1nUk7pZnP1kwQ5FyH2dDD6/2Dwc173DjeFNY1NKPaX
8i2+jTpMj5q9gWg9P0gs77QgwA1z/yJHTZLfrh4xZY1gGu4piPL7jh3d+38p
ignk9LxguxtCEv66HymAjQ5ISAbX6gfZ3q/0C4J2/nc+Gg+l+Qai2zNgnGTh
R78h6R1O1jMdOjGBRtfDv75cnSZ+H/DFK0FPR5PXtw+bqU05xbh919sIEqOT
FTFmHvZJZcWXhfWFwlJbAj6eE2zCTUAlQ3I5FyWX7hTVdN6N0eJr1mBVLdDv
jexTAzEnjPuyywN3kbZh43/JZYn88D8Eupb3SoG+//Hycc7Pw86ueYpLC0J2
nVnMUwIe/T2hjnYdFti4CsX8V4/dsLEKViSqLAChxovXPlphJFZEuAOCkids
JUpjGi6G0k1rUCOBqTeDDuhdcwd33AvsFREQLuhovz5ow9qOokjeqAf9Hn3y
uDELiZWZtaqnpQvNsk8oI5dDdI9mkYKoOz5iWdyX60xz69+3x+VSqgims4Jx
wF43wXThyH8H0rNl4m1bW2XWeOsscuPGpPIZOMRr0IUFeWpOTgE2Xdw8wiIN
zlqvw5zB43Sw6Me9pRWFtr0fXBZzyAomq8Nid9fufPQRrHl4Hb6N5RGLIHpD
YHRBNhYcX5tSAr+EteLUuj5jXZc+Wk1p27gySlz5mvIMZ7NOSIXOjKJ7n9r5
dQsMtTUIWlAAaR3wt20B8e8INmr+VKa0mHChRdZ+/vyvUAk4endcZ2jqY1CC
1o6dM9JuvcM7epgWNgd09u0Jua/oLHb6uNKJoTNl1rKUUMxxTfM3ehIixo6e
g14yJD0uPZ4z9wR5mIYtMmsIzei6KW2GvCcQoR9AFGgLwUuS9rZedz4tqf1g
KA/9S9MFHvI+49puZKCJFGcKoLyvH8LHFbOo/WIYJzlOi/cgvQjmaXmArflR
J02+OM+UFbdgbzfCWHY/OCGwHwtDtLxBZvkken25zIFgjTQLimLJXBJga3pB
GGCIkzAKn0RDwq22NLes92jHIvSssM2jko1TU/r3CJ9Ubu/0Bwdz7ZK3nDAs
LL3MXTVUg4b9o4z3eSusV8N+mJZtU5DdLm9CIz5tOKRK/WrOMBd0rI0D/iOv
BurBoZkXk5HNZa0j98BWeDU8XNWT1n9yp5dU/Ddj+ZEuNBm6crgnN18DyjYS
fUyf/I3ExTcq63xWxWuHImNemcxGAEUxlb7uAYJ1iQaCNYjC+I3zKNuUVInL
Bc0aRMjf2fCYXmnMLFuJpM6/rPqC6xDxfD0NPZyehtvyFP89X8TwhFpw3oJE
Abk/kIimQN4PArGWYQkPkek8NJ9pYRfahUcYB777WTkrvULkh89LRdRhsy+d
jxKgi+WMqsq8MYiIQTIjdZN22KiX0F3qGiyp18AC+4Re0R93IxUpGCOFmQxR
1FGbxP+tG5GuyNVMuKhqC2iTLeWJ9a0riMrg376Up1v/DBj7BKTRyjGllCtZ
YsuUhVSRC7SCsz/+7JM59tU/6ZeS/w+a6tky1ow+IqfsPn/9XEYUXfdK8JUo
EOIaLyw4Mz2nJGAMErd3YmgT+fAXFDKCU96qZxCUpixexCZ59n+IyYCic8cb
qm+YvPiwbn5DjC3P3ZYrrPJfNtSHwzYtzv5Q4zx0F12BXQsg3pVAZBqbgTaw
10z2hjCbcG9Xhi2TR/WGDHxBcjUjwU289RFuyKujCoLC4xeb1M1OqtrFvkgP
ylZ0qY8xqQRsO9+R34MhZ6cAaXEXeW2TSjXvriHtvGVCGB9v9E9a3rZQ/MbI
5ZSYYISJBoCet1R8DrzXnl/VHnqCtT1mQbBlrtohpJ59MGPqIEEP4PFr5f1L
kCyBvqebWcLUSwrQRxxjerSnLHqd1qmPjoDItDZhCoG+YPnGRZ29STUs0Fba
yk5WV1H6uBhakq+MA84dZhaqtFPXJaSPR3BTIKwn/yt8S4Y+lglgo1Ojxob8
YHfa8NXGFUHGYMxRFoGNjAfj3M+ZmgL6CEtWtkT1MFV9oUdUwzPbocVvpwPf
SWR1934QsIoR/l0tvtZU5o/K9SN2J5id0lXYyU1/hEuhmurgPfIaYr2BUPrZ
CpWSINf4svPHrxMdWH+8ARi9NFHn+bWmlwloyDw5WaigU6KeaYUnyvL4cKO6
a3CFU2EptYhwjabc6+xGlmf4gh4ORY6DsaY9vvjOLsed+hwmJCFFCgqI34FL
2YCTzs+OBbKRwK6pOWLuYKKHaiidTUmEpxKkOS0ramp76voXH4gWPfGG9RmL
a/0LvuTtcICGABtPtvZxGZNEk3nQODFoXESo4VQN0KJeWDMiVw7lQ90J45t4
lnLXeCcak+0gihRd2/chu3IVISBAhDz0uWFbzkA4/IJXg1b6ma0kwvuCpAW7
VFuk8DmK7c9/1YRyTL+SWnfcH4PhaJcsoa1OOgvrti9jZSZNQLT+FAnkv85y
mZuzJBURH/FVjdgYQgMAn5gpbm2gzOzkos5LLfElKDk88Hp0R0B6fBIiCmkm
73bUhdMVcFENK8Xxeq2TY+nB/ZySV+uvSxxV6vLyz8CJsvt+uCDWmP0QPBL2
EvAW2KeHfspZVoro2+xr995DeWV9Rfgf4YIJkNbrULaa8NFO1k4H4A+12mtK
dkq+vV3c1SDzm0GxRec74Pb8h5KwKRIojKd6t3zjDbEj2BxhBcD0GvpkfQZz
NagO0EgNgMd/jKsXNo53hygxGBJexcBE31nJkJjMaG6J0fPLcGThYrNVZw9h
dMSBrOWZ5fOtCrokrchVqCx6VJS9AezzIJYVzo21XY0NLn5FGIMJ2a+EsEll
kWBnJmKHXm3AV1QrTxUcP5illQqvvhaJNlQAfyRDwzhtEr3N1MzRtQz5QoE5
k8kGOAfak2kyeE4JpIOzpoH2YqPoHVIehc/XMGFSjiQsvI5rYMIZmgWBzWnH
F2AhcXqs+P+0vYVOqJz4sCZeKFyrIoFaAGDbQjdjEdFLYZL428u4DPIWnk7t
TRR+ZE6Di9o75ZS35UrR+ZoKlAJS8vV7WXh3ZrRTxBfhiIg28AOHNJZvUBdO
S5uAwRxrABdVgq7a+oq0Ozr7Prm2JsM6mS8579e8DYXwBg3QkY1bdu1f37nY
lAuDgcn2+ZILSNQv1CYjPn3iBLf5rLjJxY4FECWaWHpZ6sdfNRyTNRwv0SL8
rdMRMHsg9J7U7p42wd0HA8F4PEvK7D0rEC4wcQdiaMlx1H1hwvq+UWqpzshu
6x5mwQrZ3sdDDVWybElk4riT0I2Qd1ruwjYnmVlIMjndLuXjWp+yES0rznDS
QqL9QpTeT5Nfo2RKjzztPPi6oXEYJXDC//j3b9lzXoeR5/pCHAYN1ZqeyX8h
rk+TQ41Xb/B/GnhydSN/v6MNAPt7Gi6mdCCQb/JN3+GL4W9pVIiaWDa3RYL7
2Ozo+/Lv2RSqnpk1r6DIq/ztIiWOYgGBKj2+7Yr7+ok5neBi4AnZbldFarRX
xEwxwi/XWauYQmDbcfMbg7cAdq3xdCV23oxH5WEZPYB/VrnfFlTlMCQ8i40Q
a5jtCzsSi28PwBMxuvVFZnRrmYqBUXqraLSZLPS8Dz/v18U+IDu5x9S8euSs
JU0GHdShU1jrfQMbRRV/abb2uQ/pItq21edOmcFChAPy/MwyzGTH2+FNX3YF
YUtld9QJNAOojpK0zycEbfECOd1DA0bC9dJ13h++mOMqBqdaJ0XjQ0dlWp/b
cyQQ4jy6dxhfuYQwotvxmp2+tW6icr4calgTVIeeiUbADhB5vrIZgRUE/0GV
sbdjT8pyVBnBGqcqt9BTwvTI1s9Az1Y+eibhqkEvcWBupTwe+i9ayTX3pJVt
NdRIFDp2YfrYCZSouSFj28WwtNsP/6hu8X2l/GS5CdivcJiyn7ZMXtGp0vGQ
UKXQfR5lV7qhXlGOX/iGAqRarH1KyVwOR858QNgb1p+sg20mJSEKxhPwfzf+
KYb7N0KwRABlMlxo4rJfEiiNM1JT6+OwAgmHPetJpIiuBpw7BMm7Lcx8a2Se
vF1mCviiLV6YAZiEPBTrY1DPhQoo7/3L9z/0zV1GgHUpXBOJFFr69kGyT75e
yKTrKAKn0525RQnUY6w917x8AN2etr0CKHBi16w5+/0tOZZus61qO/dEes5K
/lJbH0h1BU4it3AVoCXjZ+Co1vAx9+9ldZluBQ/LUO+JIknD4l8xd0NQGXA8
RwwomujACWBhx1nLC/ynHMcLolB1mCSpA76vOvCfyJBqTECwBMAixch/9pIo
66WZ+Wnm7PVORqDwhFnoLW/1tk6W6Zwp7Tcb3qX4dNME7KjgI8w8KHKdkqRM
hf3zH5Eq/RSKbz6vaQMjMqUc3Iz8I/TBnI1FAZuSV7Xy335CtkEe0tZTpK60
gTCcQhkEZPDjRUmxnURQJ8EGoomupWNOtOUzS0Zwd6TDhdc8CwZwWe4RRtsg
ct2jr+hqKlN62ETPMHnD0UPcLOFgtofJU13olz4HcsMpp+mEGJm3VwoYd3Nf
rlCrofP2kbG12ak7Ee8giHogOE07zvdyCTnk+QSfDYuyFT6MnzmGvOpso19w
R0EmNSrgiUtT4ee4ZEFnwiMhbK2zen6rhJjheBl+L0ERNpOehna7hnEw78Iw
EIvuELwhLUzj+q8ZjtfoBEt6YfR6OyDFptO8ne5t/z8THXRfPlPgh5JNvKqZ
r1FLS0K0wHHh3/24AwNS99WBw72QJQzYPOTTaYAcWD57HRWBXokkW+r4cghY
jiD0YjjiCLk7LtxBO1Sgtbjzoj5XGe36CYDYPSvqnGKEbVdFFxEgJvTr8vr0
skyvSnRmVFJChMWsj9jr3pgHNMOWzgZHCok8BR4H/zO+ITBLLBLGv4hUuJnY
fe/qsyfoOR2h8CZ//kA2LIPS3tePkzRLLoTOow0NP1oMaEwa0XZPm51HWnXI
5lB4KG3IWostytHYMcHMSOXXlAZdFp1FR/oZZJPyHrTe3Qx50IAztESYx//Y
jEyT6Qsgx7XV2Km/8hPpx9DTcJC1HFev2MOrNdc2nL8AzXE/Kc9kw8LMaJ4x
u3NDgMUm0FyMjyAlqe5mepP2fvlzOvXHkSKKrtvGOzNqHWnbcz4dqkNgecmN
UT3lfTr+QGHDdTCinMDmUt5F5pMigt81JjMmL/BgLBnzsGWbnT6hUrdEM0IK
ikr4vHlhYNcnp1pY9UMnfJ9A4Nd1mX/oKvdOe1Lwvwuuw5HOp9Y4uAC/pNV8
wCcSqkQLF+bVY9mCCyCWMtF6ZnqgDbm71+YDrTj9Rj87uqvWffctpgONYkfD
DlYjvsCSdt2MXeC7i9QA8xzLy0H/royfE+upT7O/TXexygWiPg4Y5RhHWha5
lrKkh84ZG6mNMfAQQIWpPfddp6bKDNfq9TrU52ZOQQhswWST7/xgEOG6Ddks
/Xgk3IK+zs+rxM4d8mHKBmYyQOB5cz2WZjI0Sx18QJU2ZLEHHU2Oyq/0lwgn
GgG7fH5ZRsJkDia6k2u51M4t4MMe7pglbMesbtqcmgf8V4sBWHduFsPp591h
Tniwsd7csQ/iMBM0Rm1fyWJkNe/UOdbcVleS8z/qYY9lf3ijhQIYdvOq9nIe
JzOpfjWgbrQ+xnlASKuzmmncG6yv2CDfEuASKXYQMlkQWLssFb6eT575sDaA
GAvdgxKEcfIUPDLYD72IwsHzZgnsSNjaUGN5KMthwMpqB7z29LKzMdL68A+k
KIwn194cth3fOF7DeWHxSNrpNQHwdop82jT2tabA86MjRwIoATYMsUQ8vGs5
jjkMsoy/Ht5cthv0q7REEezJQA5BdJFFdQafpi9M/ULrQy+N/g5B0hRPiHa2
iOSv54Qx50UIrgY3pYjzGtVPuHar/r4qqnqi1+5tqwR1HQzIuwM2xSLHOcJk
ExZxCqtCjACjtuycSirT1TcKp860LQ0zxsDJSb8pED28SHrHuhlTaRbCu20K
yBzZbgelNUXrVc6TAHc19RIfXKXGHynxD5zDhW/DROEB+C3iiMalFLc/MZAd
jKipycJgMwxybk+svLM0yEriMukWBMiXa16dsMUBdcCwDZbkhk0CrhQtv4yj
1qWiB3waGAWFg4oGUsyL7KbRXhrXNmKE7V4yHL6WZaziH8Ca8vNn930Qm61f
yxZYcq7GSLPB8MWJY87qd64YkenPD6qvZ+XAjomyWL9DcTnQWQm+irAI4LhR
fOv67LupdMEwIKwB0zJFue1XASvu1cvHEbz4n5vQqQ2wQBBbS6OXVzNDvHud
F1AcMr5eUNx96j+4oRHvDakSpj6eEZqrsReW/58gmFbyYt1sDPA786I1ijcV
uZffInowe9KDwi+mp/3eDY9ip2OrqZL44+6ywiifNPVFnD0UItIdIkZh50tW
3t1GMLr/gpinGeKWwuT1ZnKwCDu54FQ8k6oXMI/CwCNUMOjL3swl4Fdk+ith
AyDqMdf7laVB5IK+3gsVvFpAAKBqhWZT+P2hNEE/xAYCHJnrYV7Cuy1w/JOl
Z2geGFYS825+MZwI7GlsybOsfthJ5AxTRe/Tfnd36ICMpbQCY3GlxkT3IZd2
GG//4XCzLEbWhfvPFyDqPAJEobP2wk289W+pU8UGwnpJv7IsSpi6olEnQNKF
bBnaU+bcZpvdNLD4WFoF/u6LJR70Mzi4inl/9RN37Fq4OtNMP3dxaKY4wxGj
bT2uC5ahvKt4pgy9yUPcJCiQUZ+nwxJ3hvbnoKf68OkGm1WJpO7dWqU6G9im
BkWLnYDXGEY5ge4cKQ/tGGK342nXk3hc6NiaGuizlJcTwuzZ4dn2KA0OLyko
AfPGA/6P1DpSGA5oI9ns1OjEpfnFIRec6KoKBzROh3835OLAsk5Kn/IUX+PQ
IgnphES68ej3pezp/LlThfA4BnLZBfmIhoJMURg6nfK1Y5D3qb6YyjTfkqp5
A1OcJJYdzDzGD48oCrsqiM7c/zi5iJkBfA4d2Kb366uVQdt+A6jz2n+YDR5n
1azGW4nCuTuinAkmZn8kxhSgMO0Qw/hk40UYwm6XNQLpvSNcIkP/aXSnjzHc
4MlF9X9DZYVhtBvWON/em5EFrj3qYfpVFKxey0rmNbw6H7SwD8yogYyL0WRs
8HZmU/Czxo5prayWTXXsymDq70q8SjA8fmWBH7QEzIC2/2KV2d2OTOf1edve
p8J9CsAvnJH10+TNVcmj+4dJAXVx15DPEwVBh3B6/HpZnW/p72WsFNXLQNhT
2+guM3ur32r5ftTV3ZCVJMtBolY4xZ9sQQ3yqax0Rj83q2ijKDc/C8aNdbEN
MchexQn9a/+OGSVxrs0xCw3E1nL89z986TZUxB7t1W049Mg3Rt74wlO22LZP
+AG7+X7vpm9F8yl2hZwnQa0Z/Y3TiTNv/IXEmrdcZsh1nL5tim8r4EsrWEa3
uxfOlog9cyFQD+JBgQlUve8+0ev16ODThruluqWlD9JKxKx+bso2Vipue33/
4RlyQsH+as3Q4/ZCLAxst39c7SEX08723EH6GznFUCJEX2UsS0W4bWFBQXMQ
jv4ZhZIBlLbWFZ7hvgoTadhGVmIvp4diE3m/69djqFtwb9QFhzYHZlzTJyyG
nfFkW9mRfPDR39OIqlp8wIwdL/JNs+xKHWinrA24Kj/9JZMHkA4CU0eKNMH6
8Hr9sDS5ObeyoRq7Cfe6rP2eEVhgpr5bT9NKyxZp0z1yw9ylsKbBqL7tzB+D
pht69iUyreOchYeu0qWgVRkx2CzYa+K1NTmSQHIbVFJqEJZTwiALY/ljlr3Q
TSkAXqP9NtcqWfH6NWbc3rT5dBB/ib0h2B0DoiBHMbQx6JzQePf2OrV2lN5t
yW5wkFYl6xY3YA1ditztwdPYD8jyHN6O7WSMfXDHfkWEotWiiikZ5wEUcosh
KK16MeLe/QWmP7S8Vg3d178hvDhxm8klN6JZkj6WOsbWZAeYVDuKVcO8CDOh
cXVHUfaYPJRiFja91AvG+IWmXAszNAiQNcTFwxl6FOeewTVtWx3/FddB1uAh
O8/OhDKa/Lr07FsKHXBbBk4fIluvo40CSw3ENnD4a9RvZmic7WnWau/SmCW3
29oy1AIO6eiJShIcmSWqnObfruOg4ogZTHDayMIKikpGBNG0insXelsgz/T/
spmIcd4zqD1IdnoxDPU2uqWQYYApzN60piBiyFQRVBB9gHoMC8x8sRwkJ55f
LfwJq8mGf024TNi4RM303KEe24tnFkYeay61YMKIN9SjBpArfie5BDI1WQfX
fGT4IO9hV8iBQEByvgAIG6QazoXdk8Oj0c2Od4av8jXkWoryRBQHrKawoPEf
PI2zgsfOFETi3BrTVS6A6WzIdDOr3PPAcfa4aDFgNmcVO1EX3xVVtocj0qFw
JhHOcJdZ+uUcvV0yOnvtf4mRyImxS7yL0IkFn1rUFVCPVBCUT2KJm1uX/Ie6
xXCd+74vy0XzpfPWFe2DyE02LHDB1djM4J5yF7Q47b71tS78W5PanWO3U0tM
lA1FQf4Me5tl8LK0LhNZHCYGLUnqwsMzy4tfM6q4LMyXI9kMdNm9yZuyweEm
NVNkB51zpbQIIhy6LwRl7E/d+8ccuPxozfCY7BmywSdxs5Jo8UZUBNjKSvIH
LCi9FOmDXn/Yn6GFllxF5wcbiSSteTfdZ+hh4vTqTZOp6rjUzYG5xZsebaPr
MU5r6m62QLRi6xCueL+hYcozKYNrWKkr865wYylLBsXvpthFxj087xQOhLby
gpeGcMQpTnBUkwAAtx3IRc0MlcU3cXB0+cxXVQx8m7VEh1nG6CpHbRR5W252
yZ6YEVyfHOVSy128FifWJnAHfKUl79i5hXUlpLKpOJK1rAESqoHzpEPH1Vb7
guc6WFdSgqtQ6mViHA4OJol77AgB5jgLr8sxzj2+ybq3SjH7exc4HYT2E1h9
LjXl45kKTBrwZb9/1bmbku10XadvGmAk11CWXOii6km1RA35v63Lj9o8Asl5
13Q4TrFrLJEmsaBxF07tXEAx6VX/ioCDzPUFH3SqwCUTUu0pgTzvY6pEwXje
zPD3bYaa59aIME8wmjzGlpK4x7zutwBp8/OKBe92lAyft+rtsoOVsjjzoocM
+ipQ0/fXC+mqx+UQsjs6CqMpTgO/f/Z//1Yq8gZSFjMYAFhs/Ag4GwU0NvpF
7azCUyqVc8LiFW9vxaCmoe4RqfgUQjOWqF+fZqsBWXOapBYzzfY53cHrO5pp
hYzWDmfz4ORpM+n6MvtusTFtnx2yc6YziVTYwJNs7/VbBDCvNdXlsAmKYHiv
p8F0h6thVnjB0YQm3mdtCjqWURARu05kYsnNIqdNvP/KD495xCtK6w/YeWzR
kmV/X1tXovJPHPrwqmslYsZw7SUAX1FUPvGzqWUZK3V82zHS19R1MG9hy0ls
J4ixZAsWGLWgIs5NkdsJVCUWIvTF2gQ6OL27LO8h1MkHkutbUgtr6BIfuoXM
mDaVBwgYTpeW2fpqGoXbvis2JjDcC20/lL0sDcNbZZnzLq1M1xO0n9xbFtE6
gQyivVBT8118gZzYf4OT2LfSDzRWVWMVQNr6omJ1S8x07QR8380p0hf4fWNT
qXkPeRyUSaox5lUfb5AZLgeDkxJsqX89yHUsz5R3c0/GMJgI/wPRB7G2vNFU
tk7VukbbcF9gVjpDkqUPUJ0RZ/kVYihkDT/PPN6vuNp2wjUM0WrlJILX65gg
MCTfsGKAoS+yeYmL5NRFdrhC+OYGADyit3GwQpnd8MDV+7vezkXFXvQAB2gE
L75ldBxbjmQwQA7LOtF1ZzADLkQ+UcshnRh5GtWT/AwNrh+mYe8BWgdthb3R
xxlpr8tyGdH9+NuSEvVjyuaj0YllNgjlHFFe7BvZEs8PNNen1GzBEF4JN28q
TCMxxOeyiVSIFjXSUh5U7DvFqveROfRkffdc9+ul+3K6gp6fbBmKj8G20c+L
CZzA3AT847LV7zM6Pii/dq+yadDE3fOSSDzWXwCq/tuB4cMHGznlfRHHGiKf
P+nVLxdIZn8YI7lAI5i3NEv5ffltO2tx5FwNy5YWkjO5NUfcKpwe87gvvIe+
rjAuEQyVOsagm1rP+7FT0Jh7po9IYvXqmElCCeN8y8+KgibZruAglbDM10D+
y45lpTQ57sPhmXoHk+13TqctIuGgWiPcKIhjWpN+7o2ffa3sSI2Q5QhzNnt9
uWPGawWhmIF6RALGOQTWPLgJ5RJWS8XuwbptX0o6u89sI2Esr00UsyV2dacV
PUa7Ox9yk7krMau6j0Z0poPJuIU6MrUU0rR2+HVkxcFAa81r935GRP15T8pU
ljh6SfgEbL/Krl+yjL5VFCUJIW2MefbmxwFjThT6M7yZtLcgyIaKx9SVS9oK
qlwHP8bvJwHHurqJFcZpJEtryMFqJ5YJjQd5gvmGh3ubWmTD8WAJxP9wXKOt
GLVRzA3V7auhc7FERVBNf4bYRoOpgiVnXQk2hx2DpHLjH//a5wicFmEos7Ya
B8IinuQaOYkQJz84lJII3+urvvPO/n3gFyf/aimuF1uWvnCVPtiD9FMjeiAy
v056dH5mBsrDsgJIwby/RzOFNP+99yefVcTHeRrUo3EAqB3MKvf784d/+GUQ
H+qFDY8e/8BGpcM1ZMC2ETtQLq/KiZ8NAV5kN9qt239lSTljSwnvnAvRnRJs
fizZ2TcGDk1PtM/Nve70sqRj66OT6aylXrTK5yiONlPQMntmQzBy+bLOc2do
VAZws0W0DB0jMOTNq3Sxhbs2ianaBtwcJtKmc0DNCZTK/Zw9xC1zlb9YwIVR
xXqHspsRRb9NKYQBDd2VrrBRHu4a7KSxsZh/FKyuzkIXCyeSQtIG9wkdjgOp
dZePvb2U4kUMixxmRIhqbce303n/pDqwO2adQAf8lUuNe51jaIqdisUzr/w/
GomnEfUbEuP2EgwGrXUmsLXJHskVwoLopv0oZ2NSRCm1GFFpfixPDj1SlbZ7
K+tKdx2c8vet4raaKUWeIr3xJpX6R4QyrmU4ayNuE1gPEhbBHiLN1ZxiQYwn
T9goGZEB9qTP8vAJ7KBDxb8qPuo8+lxolKhxnVyXBprwXgR0H4aJvQFnr/DD
2UGiPwK18Z1NqSVUTcbiqUHpzZeC0lVS8j8GympzTEC90gEkvRgbvO3J/wxT
e5OfRUSQ/9lpkDA2x7p/z/QG7dYjym6t2tqmI4nvlcwBPE0EebnAvrtnbGGN
UrCs8mchrn+8P0NkDbD4p2Fk9KbXSAmBIid9VHFenT1za+CPnisbCTZX+SxQ
qQBY2fM66vnzR6AZpQgP04QH20KnLSKfD+IwjBSzrvnf0YuJ3zbLXATjsYky
RkwTbo3B1w+51LO+VcdxRldioZEWsqIhL3OvXiIEyqc2TPpWcMYZDe1Na+cF
Ps9gjcSX3Kx7SjDpTw8qay3MtIxrjZprUpccJKZpZz4c9/qthR5TDNL6uecP
9eDLMJA6WeUc0sBGXZvsgLscqWD+8ycylzlXg8blydT/NP3G2l88YRRDMJLG
IZoxJphioNHGSUiedc8hpC3Emniv0AQCneKLlNbNZ6Go7OJ/bU9RWEKHLdmj
l2sR9SPBJjxksviJES6ZeceQoA0to6NJUn3khPdcpNkcSh60BhupNfh2xeK9
Pu36r/GXyFnadvtbeYBd29/AxnOLwXMAW8ja2rlPRJu+2Nutofo7fICACVg4
ZcQ5p518mQ38ub/VJe3W6P0xjux5zbiqwURD5az6+ZyLf32/aF9Bfqon5WJQ
cTmiQ33VheSR76YkyicTstBK7HqKs2+S10N3u67GJtu2t3V7AyLmfXhp33+Z
y8ZLzLr4rIBv6SxMJRnzb86dfchclhA+MO1UWrrtqZqv+R+kVOsz/KN+WIx/
t0Xyx4KRvrkhDb8b2a6GPCdV84LvSloosn6l+kkdKxYgQamdOzoM/o1guqme
H1Hpz41+ACRcnqt1nxKqBzz9jbcZFYY5OUJ4BlC52wuXmbwwOD2KA6an8YIE
eHhvewXPyWNk25cr6Yxm5g7mSgVCg+gE6Qwyln/g1wW+N7RhPZkpRxXpXtTr
IF59dF7GI3uf+u8koU+6g8EyHld3eGLdlzJEFVn81PA9HVVDnwmJMZyRWfo/
Sr7E1YkQKA9uDp+Ni13wpdqsCzbMfxNZSRUReX8gAU8y2VVCiX8SisyL6SN1
p68uqaxA2LGLCsL3Nn4R3xmYT6RPHzkRxKHmIGh/v3V2V8DiZrGLk62P20oC
evkinvchUArtM0XUlPF7h+ulB8EtacJ1oRtFOB/ns5dAWvvMtCIHhVl3+mSm
rd9hicdofI+aaCgDoNGDTQRqRi1PIwmL8zc5LjzxwW8bJj6GKFb40nGwqmqo
f1AVuJwTp4v3GzvyoBtNYRWuYgdyIvDIdR0U4khA32/7uJJNTkA48+ZzmF26
ON2NLRPJVW40m9LkNNiQAK4H3G/UiqLUB65v6qSjCns+i3VIhBAyHqbs2Iz+
kKGJGXMAJSzo7HIzuIvtGTRGOMG5sN+YRwYfKvzmHhaxoOprFrCtVubrvRkL
o9LEaQw+XmOEWGmsGw9IdNr1hbdspTsxCabmx3k8cr+JougEwuD4Ypk/u98H
O7gAHir4m/tPrO1oiAqTKHK2UzytrEqxaABuIPdMb5dy3f/JGf5A4wKqsbI8
XmhyYEUkhnt/YeGAcZkErk8c8oDPQGe9fP/vOElt28UGPfuDD7OsCUgE6g9Z
Qy1IzJiuV0i5AJGVQ//GKQzEsdE5DkazPWg6bGrpDE/WK75WkFTWpEPR3DgL
WooaohRED5HmOOxj2K+GMcof/Mlk5lRKzSkKUm4lkhxbxugKOmmUSf9LSJOu
csXlZxzbKuC1hVjZTmAYrFFS5bJQA42X3Cdx/ocTerVwPSGb3p2GnPtr9IAg
nYFBs0EzHp4bNYtiM82VzcM/0YtQsID78lDDNpMdKoVUygM6fec1NRZC1K2S
ONH0qOp5cHGHxOgzAG/ZC2b7vYW15jNS7XU/oZdZMUuAOVJLVKC8RpJDr5im
SpzspaqJNlHAC7onoaBRSy6E8OpCL44Iv4e+9ung0ZctFy/9KOwFYJOrKdTJ
Zzq7w66FWZvYPKWKap5GGLvN/oUGjIeqhR7t0XN4CueWqGRIOa90HZsktAUD
yauokveJv7U9/eF3ZtP6rH46E0nUo+JYVsgVSo+NfEvKtvRwDv88ui3UsuDe
0It8V7vXskbwU8jkW1YTzFs/V/yQAg4aqumKeyZ7jbUz3hqe8HJyTBrejCM2
Yg3dQ8ag+lnre+lz2BM05ago2ZefKYUt4MUC18QaiFgKGF+DqbBFsGnwFl8X
neHZoVa9Lv1dVHL8BPzoCdWFNisAIEpsXFFN56i2K8EXhmrfbsk0Tcry2Ia8
0YdxwlpA+xYwLHmBhwBgHQMrvgHY5yOxgP7BXmVgQipr/kNJ36HBuH6GOjcy
oCRZgzCN9+F1MSIqfmGyFbTNIsUWgeOjFqQVOFGsGUEzDBd4xFVv8tEHH2SB
wK3vQZl+4WpFYGW4qbQlZjwNl640wBZtu/q7g48yngRjqLhpmLAVajwd/XDX
XRV1/b/LQsELTkoCX6iW7JPLBHwsT8SRKrJitcf6xNpotnElJ6Wmgx/vX0gQ
1Nnoc/cYh+5asN/Wrx0Yd28WeRH5rV3oxZQWQAmYn1MOycVIvU610lnGAu77
ZhL0bljAIV6XGhuIgCr3ua9k65YU0STVRK8B+H+w/2myMBYLH0dY5Tag5/7K
ape8GTDJzXI0eJGeR9SbQ7aT6oKoot9GMXklqVN4fNi61LYRZAnOT7gU+V6K
WO7lIorhbvMZTobkd1ETmoJEYJJdjxs8/6mYyb4uxBFQUPoVCjAJpWUqiwNk
7RzOJeldCvNo4HzFpNjc/9CjS3CouOt2dVPoPROuzAi3sBv7zgUxs2OCsPx1
mqtzo0MXBEsNJZB1Q0o11QuA63SOy9RcM4AQzaDO+A6Ynsm86pb5cb6QQT9u
LKENeFhqETABc1ZI6fuYYNERidRCcAyPI8SqULJuf5kS1AO4MUAfjmDBm+t4
gG3zwjXui6GyGMCov7mttoKxeGMtCbHRd6iK9Y7+1m7AqQjVq/MGIFcEBEtE
oz9pq2jHOGZOClQHygMkseypw+Z7BzKKxpilpUekcB59EPyfpqjaBsuC4TpO
VzNrGYg7F2bu0qps1212uTHswezCCzDHPzgAoTuAUz1WYOLjH2Rwj1d9cwHq
NB1KjZ2+D7ajTeW9KNq5TgJR1PZkufWby6e90kKjMmLL2GA+4HPnyMGiSOv1
RSezHhJBNnBrLW450Vj/mJAeXPbwRUYvDN8pnKHRiiUZJJeViVZKq6roJVE3
ih8ElIQaX7NmwMLDbN3LTr16yrkT68+dU37HxyhZ/+BOziA2wYuHhgNHmMs9
lCtNhx5EZ5TcOdFaluzV3adsi/hC8FR5jBS0UlQch7r98nMwti/UNfjOHB5S
tJYcpl6f5DTSI0tMf7fIBPEKtX/C43k46/bAp9LUNersMC82vhJHxYZ58xWe
9RfbqsfXRK1n0lBSUPkPySlzeAU4KL+c52tEz5JEtha7e2ka043g+8CKK4q4
bzY1ITeJNYBuV+BPlf4SDVd1wzOZqPEM83GRxTxiSaCgXdcNh/HgTlfJHJ2x
WC0aYCULrjoOR1aH3yxr55iK8l8ZmSyAVw71lAmxcUTUAY/oPyD8b/11WKeR
PVFCIFE0jhru76SNQ8vHBkVg4/e+L0bG3vMIok7/8ClwWK4Zc8bPXjx9GNS5
MKKnQQLabU4MYvtoG9OYXyaFucxF+gYVzIJO5XZ+GzfeQgCs+6Dwwz20G5vE
wZ7hnq4Hx3nSDYa/kI3J8X/TXlYuyaMxtTht4ozIDOqLvkfxms/qpzmOM2u7
l1NgHrEjud+0TzgHfeFyfZKCgXxbfxuv3K5CKKag5mb5EKlUkM2t0GBzPU4m
L8NdfXLP9inGFAl4NFcw50J4t+GyB0nmT3Crfnm8F0WlTpmrISk6d2CJb2O6
Aj2khZf2c6Uy3JYQUWlzIoK0Dc6//MD7vO06feR3whxl+cwCJq0visd9uM33
Ya/4zDRG7v29Hp5w0z/B2CcV/lyC4rYjUZ3VPg8EneudNcRgN0xNKU2G8UWj
jbACa6B8CwbSYCHQFhlT8PmtIsvFcKzp7bnMKCc3aZFOUzznrbYMxytLH2fK
0S0/0LavoJyUNGKAC8DW78Q2ZDJg+BwDVu3EQHO5k9305QZEljaKXU65ivDZ
H3UmCltDxtSw1115m7z2AMAhqzVN548KXhc4BQcjq7O1pEE9jtXRum5ELtfX
fj+iSNbF0dFAqyI75neOWf+ZnlHyQ2sHB4nwlKyIbX2WP9mi497BxOlkP+nk
xH44SbBPxAXYvnBopiE9u89yTXUGWuew1TomFjrzaSFvetJxTG31D7xO43Nt
S/iCVxjNSGFbypbwSgznyIPtjXdFFKkXXyl/NQtR9eIrlpuQx8D0z9C4leXB
l47DX15o2vqqeovm7/bqqJfnzG87Bk2ube1ghvPC+NA7VL9gYPnkD2+KXKYz
RhLybIvwS6BHZiIYw/WCFGChy5EZVzQcbSCkz+Ua21mFQNukOR7kkMEaXoan
0orJsu8EgpvWUPaZH3kIpmtNIsWpAM4MwvUfGUXv8/1zRu90m4OCz/dHbiWr
V0360sUbmyZu1CtR2Bzh2ZnFcQUrBVhxjxvD19f7LgUfmGUw7HgOI6egJ0+W
z8bnpxjdR74ZH4HAN14U0CRiJOql6C3eq0yorJBALSNPRmIYnX/yFODyokcS
OP6sjBJjjwZU3MErAqAV72vPWcMQ9MYO3D+cO7NlUnMWRSoYYJnR2C+55fyn
8dhfEzavTCjMS4RASf2Q9wvmIVmBwgVbvo7IvCFTLmzDatEnVnKCYo4iBmrK
ctbKs7OyEXDDbleOAGrlNdgXLH21jUxEeu3VaPNIGnPFqqEfIG1bAzAX7B3Z
mkvuBOX9thxka9iPdscXgHV+sj94aUUnfHFG9PvHcw0sQxcZyv1B2Nh6RbvU
ff93ThvG5DG07VFknzCI8td3RXqUc/OFlXGWJAE9jdowhegr4Cptgvs7r+cH
uGH+ioDLePJeJOOoZJe2x47Dks9TI82XYiHIWaT3Yly1uw1CGhhT7UgH7+1k
eMoL4358oHI0yBV470Hf9PA1CqPXOpk2+lzeITZ10bmbuhq5uqdX8oGt+1tU
wayW9GRFAeLqd531+9g0cTPAD6qRuHF/gDYIQ5B/6p1vzw/cZ2nBxUVp4Z2k
rkEkb5IaE7R3N0rgZmM/EXpbG54SDbJYLlKbDFvy2V0S3fkCNvxWZjSGjnqA
ZKHHTQHc2bUZhVGrmqHFnHdp+QdhvT+0Zr7Xvpf/V8vHHfym/VDEmbCTeEhb
8vPM/pBSS4/pomaZMMKsnpFJ/8aZd4l99wpbs3xmTffeg0TZ3eVHAMTrgHJQ
nXg7+SHrdwNAaef7WwPWXzj3A5I/+vHZhriov5TEkYOzTfYjZgUr1V1RqvX5
dS5IEi989gf9zHysUvooMYO4lotT0F8FDD6gB2sN8cjCYWhjtzBcQwtpbdpZ
QOdE9LybeUIUJyuMhtWiqeEL7zAiDjpDsQaYxLjS5eenZMxGj1Kr1IrxekA4
+5sp2Kn/hfrGyOkio+GDE4Mzs6bNqKETvVgk+1+vxNpTfy1BeeW6G+m4Xqpt
BOqCVAkdK8j+Z9iIuJJlzG2plmF2z04VXBjjVsziV6mlDnfatjh6QJv+HNM1
OPEKstOAx2CmzBVr0upbQzlZODwrwsOgViuRH7nidesFPMkLn9XyyQNLpQsR
ZRx85DhPdze9j9IqKOGxRZ7sYjg+Zt92FHsOMLeWRQy39WqyjkyFFtIQ04Xd
FdDRNJcads9QrzJsv9tnoVevKGrKUKbZFB/f6+fK78C17d2+c9jCe16hsaga
Z7GpRfcxGU9Tnx0Odm1Se1Vx7W3yHLJr6MghcNbXvipj/aPmAXj7mCc0r9f0
Ppy7+itbQxmKE+fo/FNALbK8Tisp/zHkTCVCX747Z1Lc//Sx/QUSfgEFR90q
jz1aEz+/y6jHbRdu/oMCLE7zompxp/i7bZ0TBdtH7QwJ6VM9eFZZUhT3xIDm
B7FnOW1CPkUIPZcEIF/oJQp/dXTOL1Elgag2zvnF+4rR4Sli/fLpm4mgGcrB
sJF4UTq0fS11KzBnPm7UzMPKc0muLIBD8zjELVOfHnhxseDg9d1WT4LXyEGi
pJbvFdERW8xkrz5jk5xpxgXtpWHki1yrvrvcOnJA/9Q79y514ER1RKWjOmOl
JXprlIfcNSQUAW7BtwEUuwrEbkUUc25WqBRtU0VOo9rMpk8WLwqeRuqJKPse
BxCtBhaTMHSxzaqA0ffT0Radtc0Py4d6bd/ln0v9fQUPkdijuJYcx3/VdY9k
mLOlA9Vx264lcG5E3fgP7XoQ9wrcMbmTYD8Igazp2nsyU8wO7J5vEif8D5De
jhgCYai5jBR3vSaFiC9TlJB+aiXhf46KHxDaOR/wXzc4NIpwEl2gRneBdtj9
eJtBi9057M6nwrLXCRkP+D/KWJReo1HhOcURPWhHSQs7uUYYKcEdg8sC1LvR
0Y0iwPLMbPYZIkyiPvQSi9DhRkj9jQVN+k4mBdjUAW5U6x6+b/LJbncAdj67
TCMbJ/dOUtPKhGcs1SjxkudGSISYLmW0q3wuZKh0/r1Y8CB77SeG+Cvf0rIc
RXALJwINhief++dW+8pi0FDbSVFS8tsHH/J2b/RmcNYFXqOxuMcUG1wp4nCo
X3FlZM11y4A1wjHLy9LGZ8YRYGwh5TjGm7Uv7Yh+Vr6Fa3bwWE9JHabgQWx2
bIghz03RXN/tfQFy+8XNEhaQOsv7V3gpSGBzboC+d9o8P1bXfpAQ/3nt8MGe
O8ZkbW60izc/Mm++4xBy6ff1rp9L9lE9oV5zM/US8q8LK5deK8cmAw/kGarm
Cs3I4HS1mjGoQh1Y9HjSTDKpqJBEbQLJy0mzcSCkVLi38erWQQj29HJs0D1W
PNsRhC7NSCzPeE6T+7iV4Er0/fe3z1FE0skz6G+TVGn42/Cv2qARuGL6Hlnv
AwVo5RWkZj0navuA/kQzKRKcG1fL/aUdvqttIHuK3H9c5r0emS0FvT7O8VXU
uaD/eEbaDvspjcXO4F3qtwlrRKuRuVulzNDLDoxCs0aAe0+i4aok04WyRb3A
R9DBmye1jRMJ5+xniSmeVtJcUExOmiuwn4nPwC8gx80f3AmAf+1QBpqJFXZR
7gFkPu7nQlOXiNcJj51BiwjUmJasuKLlYchjxqseM0xj31uIXOK0zMKAUGw7
3mJIVHQ6rW7JDeNAIKhJZr+A4PxKpCSgWsKxgPArFS/8M2qlqk+9x4GWPZ6/
RjbQAHOPup+LjL/zP8fn5sAvhcw3Pg0qdiJHWRXO3EoUcYVHlU7oCGvDT6BG
G/x2DkJLzwOWRfWSXl6ACabl09YJ/uqEiXXHlLZiIPsXBaIFEbr95ilznA06
iT6Q90g0V6lhhZxkXO2kwdsM9D1JdtxGrOt1oly7sy1SmJkauTtXHrMT8Eza
8sdV5/Yg4GB5CBZCdazdiGfn7bUf5rCKnrgAUxOV4tJ9k0ZqRKSde9z+lg9m
jHnSlm85CyChNsnXHfMRO0ZlfjnJC3hgDFaropwD44TXmgFd+a/aYYUrilie
wWnxZgZD1dRiAQI/BuJqglyIdu/3WrJSrUH1tgPNsdZyMD2KHiX+z2U1wH7/
Bu5oTJlMOVCrNOugJzmbqWWYxbPOn6MYe0DQkHwpqWlIdTg5kCORVeg0dvxM
5zRwjFt+CjE6xGDjuS0lDnSK3RpuMs1JHfAZjisV+FwmHYG+PK2hHrRCatQv
WFCC4dK/z6a0+U3dNFAoTrOwMtunY8oy0zm4HgNMX9TXkoF/yIV4IODKG5w6
AU3oMJmhu7q0OPhjo/V5b1z7+9y5AIpCSgN7iTbtAWzwRfSi378h9YrhKjxY
5BB97eLapGHBbGg1n3Lio7HpSNMqCpLocV0S7nkaiyXBBqD8GwgMHfUQ3WhU
XJVfaQVUUkI1KpqjmWEqwrpN1QApFBycXEWrauKHy2NGL2nRZEvT7GOyLtSg
WVX+NRvMrYhDKPebMVGmwH8A3iCaAMjYRDlvAheMAL5XEulJZbjirx1ygeq5
q9Jv98vGtAzDahZFjUhGsS9UnAnn870WeEn/oObgNHR1IP41seBcu/HT8u+5
a5SiQaFm4Ewaqz0rH3JBO5TIxD2hw1ZnxhVtaJn60snqGqFgypzUWJiBmiAw
FZSCHYFmW4gF+JgRSSXsbDj6mecy+DlDNV4iSu+Scms4BuvfLKaDKIzpM3Da
rq/kUsGLIbhoWXi+c3cfw09Ru41bnsvxa3siThYqkBMEyFGHFrm3hE8GQ/PK
cnvYysOylQQYjIzAVbvd1Rw0p6bWcXVvWQXBX0PGkHfV1j+s9wPsY/ZGKID3
lsgtMjjGfWY56GPe9cIAqO412bDnXwJaSvlJmgtxLj98kT7AVyXv4JWAjPX5
kAhq8iowNHR3bDOhzhN2Wb/+fmxrMe4KZ8Aq6xMx4CZ0LMeRLcEtXang4tcg
nqtMmxDVrJgc0GGNEVfjzzKvb5UApc9RMBTJhV2bVQY1cx27SW6N7KMCyiyv
ThmGdX71u8quzteDwR4aFYta/ThLkl3r4bZbk4upjjSsbQmUP8Sp9bMlCrj3
nhsxlWw4hXHMs/rantuJ7Wqy66Rm2WuQO30MnKnlcu0zjZe3lMEJ8kO395Pc
B9DpiGMBNzBDsQzbgiEh9Iywf4XMIbf0xpTdwZOO/5OFoGrFo4w1DYnpnOZt
6g0xDREv9ykKIjVxnEHsrTQFr3dy8SxLzdYV68fogkzsz+v2Op8nzjCR9njn
kmWGlJa6gmeFJ7wuhL/SS4Stz6m1gkALWN2rBHw3OaRSKMm2d09xKCNtbILi
sLUGhM9zxYVYKPbR1sIBMFj8/oxQbJdQ/HB765fknEOutgSvMz0MXD0fGPPg
Ah7EPuqj3Isa1n8dqY9Jfsb8cPhE7L9eVzfMp9P20W7P2YORLjKpNLB8k1oY
mDzVf95qorF5JoBDkjIxzvhVa6a4SpCzuH5X79qHPSY62pvf8a+/gJrESHgX
qMx8/FJS5/phUMnARcMvPJfTpdNVOjc5fyaMAI8NqwrSjzsueGP8WByvip3n
rqyUfkSVfUC0VAdRHwX/PyumMOuXCtry9rKQJywtS2cNtVh/O4JuCTjkyFLT
A4Am/uZPRBzHQDjpMfGLqzTjIrbEr9mweXMWtgmyciS+6VzFfCBpwChQB2Ld
WbMQ2IVAhqlUGE4ENiP2sbIpepdyXuJVGxiU9HmBlfwgHwzqX9L3a3qK+YEW
IqjAjITQzEDaiyK5pr/lhtA2RqgXXqjT+DM51puytbjoJarGsqvecGUN1aCZ
7KkZZJRza4lpiQeZd/Q3rlWEXbpkM5zGIB03T/8zqQ5j4xTZxHJQCTgGgO7X
04jKhbSLBUvfxc6xTUcExfSsIlSq0hP7T0OIvRdwzENGHQyPxUbHTJjkCND7
Sh2tfpdJksPN9ZI9W6aPKcq3GU1i0hDWovKcEoNlJkwbUREB5z8YX0JavEfe
BS5w/5NnOD9MPkgaoVh4OntsRkWgGAV5nhNhK278QKKUb73+YozRVoQfFEuW
BQ4iqQ2eYATu5jXhB9CFH7S+msZKI2EVY4gCjM3LFhxNApel/fZfnpmUHVIK
2MZaLo+mXEaQhRW0Z+MQyqkhJ0t8QLIlDCik8IDurCjnLNLUgM21M31On//M
KqbjDDv8MPUEjFc4pVVNLQmx9VJWpYTjZ03h7vYrl8xcf9krERJE/ez1uo77
/Nk1pJG4SXM/6qhrfPEWg9oj789VPlN83zX98nedcJHldPPbCWPhlVLHKHoa
wUCIIjXuKJuY1/HXGKz0qTJL3dTfxojyxqKE7IOdi9Y1InDxwV2UvnuCOL7C
dvYCx/MJf5ObYr0nzMx+MNR5TldL/rVYzBA/HN6C+mDkAgDc1rFJNlKoYfqC
dp8/Rq2l0r5nlwDLKYEQEy7mUullDiI4FhFyUCuRARN8Dkel6Ux4E8s0Swcv
+z881R9XKZ6Y5o5ILqfaDJo47SgTgLWlGBkkNanwsNloyi1PlUyhkIXjdaqZ
Gi6kZOoGZwAM7eFQVtGu16aURJMwM8L2Gzv2p3CQ+iMxgcvQqvKc2aJ5HHqJ
6ThUdLTDC+I8ggWZK5v16oA2AE6EPokq869GnupcV9lUUG6jaqc0tHszockd
WEyq4udYJsUtj/zzO1iBD4VyjfPpPZMSRv4qNyb2Ovg2YISnDwCNkQwVuNAp
rJy4uGSoHtgVWWUw/a01l6Q5Nf1Y/ys2+5Fw/en8Xt+8Sd171jW2qadGFlhm
6xk3QWsADJlR6srubqoqivwxu8L4QAs7fGEInW9dRzje7m1VaJ401bCTHbp6
L6vM53j+f+6TB4Jg9gL0KYHzIcl6PMyB8slL9MG8PSvCoyIMnmpXyJ7js1Kv
3j6MiJ9M3ATFgv4EkRsJCFVuJ/utxjb7jX7oe5rV2Y1gaGBsq0R353B1ocXi
aNzRma7N9cxhho4ai5VjpzVf4RrvqQgkZICMQMLLXIVkHiYt9+28fuEeCu/u
NEN/cWj1XHVYoCEHPsMRG+Ac5XFb0NZjvHoaYvHjFlxKmqRwt3LHIqsomVQS
MdNFAAuXek5aCSdl0VwOdkBR1t+DTHvz81LS9A3k5GZ5xo+4hz45u+uVFZ8J
jlfJVBuDS1rcJ6fbzR+FAuC7es+Zi1N5NW9zKGX8yp8rLbH8+qwHN02wadHy
iy+AX2mZgcEoLxPZEtXwoccT2x2XtSNN69/UgOWH56G1/rydobDWYBnH0+cd
HrLBENykG2F7QCmRlrAcVnlAIJkS43Td3CAc4sJPXW8MQw2VWvxxf52yY6ws
qoKguEIS8MvTOJ5zPzPbi10x69pO485DllhjADQGMaCJxrVzDBVHhRzyqqa8
OIieIsIllLscEZw9nUb+K79UHFUlrj9X/hWro2o7MKpD84SuS4ccFiibDKUU
01XzHR9bFXuDw119mjjEwGwTywi/CGKBZe0Ju8osVcbhoPDGPLtTXN3/M/j8
qsW09RsXXA940HA/05HtjDI20FLdDPF0gasrDhOrPgvEWW4kMO2Y3x5FZPCR
8BMmGurcfNMVsby0Z9fIL1Bj1gcgwY+9k3tocKDFYiVxZtsMD/6X7xq+kmv/
SxE60AXaT77fPxEMrwH6tS+LoUXUFhVwZh5fJexC3nspmz5Ca2FAyJ5awiSt
KC6XB3tDLM5D1mluLIJx8DPB61cZKy2ykfIV6O9aQ3mAcsgxUiUKSLrX88yo
8opM+BOMgk5gHeKOzPsPimHXn0pSzsLicA6IcL7oJsNq4B8ok5G0aT/D9iuq
7xsXcF4aYLE3JHfSK0afXVQTcrJ8Ir28CNzdJlKaiQ2VyFotlyZ7JHEUKfga
T00uJhYgo8EoCrR8DGE1U0ju75BoOpbOC98KvW2ezrVAbIZjMSHbDcUypwNP
9ZHD5N2h2tcmNzeHSJFIZ5oLp9jqEyniioVv3rGBch/l5H4IsUNC+G51xXlp
vSD/N8I02ETfg/vRxBRj1yZiG/U0fstWHjgZe509lAcAhlkgzGCo9qacc5A1
XrkyO28BBCt1zslxvaTltG/U2sSq3UycnuW6ocZ8TSnlhv3168uG/8Z+rwR4
jR3/89hOf4mKPQQJjg3yCdDf+DjuvG7BqLrQB26A1rFZzyu7fKjrgQX4hMsY
lzE0iH/TmPd5vghOy2mmBQBeQFYlA4IWF4I5T4iVjgLcx6jfD0/atMzp+ioF
mZuC+dGdS5l+EdjuF3O8C2JnRgc9k1RRoZWQajo7FyRtAxORNEugXiMKJkjf
nX7/roSihOj4riWPkm4JUaBJsfQ5sA1hne3Dtp03lltsPjyBwsv1rAgEIHTD
GjjV4Mqz9TKwH03ZCo3cJ9FRYlJ87v2EUjheLWfWyS5hukazufX03Tl8eUS+
K1xtLbKLV99De2N7BWBng/N6eP8phSCsmvp7fiQT4pOkdawtBw8udWtxWqaL
JPGCLFFEGfhLvp1VCkJsuawHUhTYbghlAEIK0d1CjE0go0ajW7oAEUe32rTc
5FG+FZ1PZb6Fwsod0IPs67o3USC53uelEtPHbm8a91dM9hcjitkEgVQph7WC
ACo+TVpeQEJKGlcs4krohCHrsiLFeHimQPI43frfIAI1zfctFjhmO/dsKALq
fg9pZkNKVne3Ne7Ro8XTL3xjtMJPM/ahmilKDM/MHiJJbfvhjV32RLBNOWIi
tZ66I9QwutDjOsP/U1rnG9uZ+kfPvKZgTmIzfXZjzxqs0GE2//wmvlzGIRCe
GF+l443CNIb+5yAg3blZ/c/QrcBQIMJUWj34p3Hlt1U64DMGiGpI9I5DZ/hB
IWqZjD3Q+PfSNDqK/V58pE9ctRngg++DKKcnASAH4IOW1J3AbAl2TQXovE53
WiNYmQsyNWXfnyBUU9Hjd0FmPaVajKneDqoI28iicKscpae0jeChEv3enmrk
MjZf0DBYqKVfK2K1Q5DPMLjaMqDcOniBpyu++EQl/GMdYZ8SmK9FrZ+Gpg19
gda1HDajG9vSAiPUZb89R3/cg/V90mLmuXpnH9+WBDHA2AEcWXEqXaIKd6Dh
xD6PeJ6QtF64w9ZIPYWJzJaTEIa2gp/xQr4cVDpCHc0Wr6QyFYNI5cqolC9y
0QM1qh15kbtMCsF9SeZPu4Z7I1491/Us7ebdke7Bmzc59AQ6UF+jJRcPlYhp
CZ9MuAXPP0hPSA6/c80oVVBcsP2qbYKjoztEPJbANSpBwaVU6KBuGqRVDt32
TWKA/dBUEOA1o0akkuhPs2TifB640ZGx5EoFjtAKpAEgZqsLuDb6gzvrtx23
hE5mpBK4UUVqRF6wLzFlhRefi/VMSOOh6iOw5y2kIQF1LpR8dU/Shhr6gPgJ
uxL+Ad9GMy+ttmW2V7e+eRPJTKq9R8PfhJm+CzWDeomT89KWZdtohUDHAkQy
0S94p1e/QkaR2nU6E11Ua1YkGcFsDlMjSpQuCkfVxH4ayZ5fQRVdjl66tI4p
CIrPwcmwkT0Ql+NL9WUFcAzV26SN0BR2g/Wdve1JFb2SSU6tgg90CO6FhT8u
f9378MtHecufqz6G94SHZcL0Onk7qXIiKfnvlvWDnvm44L304/SkidsEmEuf
rFm8jctJDtK0ilC68axiehimgrnq2ULHctthSxe+xIcqBJ1BblPGbwbWkHo1
l5QH4UdtcNKF048eppk8s4j/V07WXUnq9wXrakty8DuaUhfQMxDJY5tQU5L0
YfrFCfV8Hjwz41JwrvrdwXfXuKbEMYszHTk1rlZ9szZaTGN4eJBfI+RXtS7S
AfYaoMpJ48GXIff88kMlJDTUDmSrEhyIzg9+aMLZjJl5Hy6JQYuoG9edcVCJ
GidzeBccWT0l+YwsDsep6M3y4G8mfRmLm3urLjTXmV0D53Xzx7lYw+T4/t/w
2oVgzv8SF9saeWeFmnv30TOif4slJQsqVRrqCXeVXUO/eCI2RQxW9ZVHFBq9
wVu/YoNUuem+Xqoj7a7USvB5tg5GEucXUK2cTj+fw9VCDava3wZq7cQwCI/7
55RItpM+WErmX6FtaEZC2ceAP3J/T1Z4ujzjqfck04S6N/h2IZiDxicPvaLa
npR+lsWTYYyxP5clQYOLNpUBDWmoPIUa7t/FsvHgIDC1NNIDvgSGOe2Ap6N4
FEQYYcVggckA5wlB47v4qqMMfPKdl7papFTvPtKN/dGfIkdsIImU7Jc7qv2w
uZ2F5Xnhz1Wc/z+3WOGKVq0N1EhqUov6DC1LF8sHECl07RBMXLwWFa3eOqDg
x/hWPa4Qb2EL9PMJOlWR66VEbISmAevcFaP0E9Sm+MA/V20gCK9LXITBSgbP
IC2lQrYYUtfHC88v6BoVYuZ0ml5fsqEp4GTGEUveho9KtHqgdYdezYaD/wm7
6UDXMG6KFLJDALzf8W2l+ekwxXzgZE8148Tff0sjkYm+NRWiVxpU3sf1pi/U
3Pyeu2oXNwIrlCcYWsBFk9cEdjxp74aCVnkAc1Qel3k/9wFK/gw9XwfwQD9a
CK9Fkdpfn8pxecQNEpBgCEH3YEa79QzUtXmSadrEAqS6I0Dz62l9ya+VsevM
6ywbLNKA3hESCwv7Cggpl5nOOtxsy5rTdPGI6jSFgCHwEkzpyIe5O8fVGgeM
2uAqmiSzMWVmAcsWv/NCFdJhaY9ZwBnY7M5brc0WH2CSJ1ciDQTukjpp3aEH
qg8l+vTzxFdv3Qgb+qo/8Q88YYfaMxfAPmdePFxkAosOGWc/dxamzZ2C5f+w
0b7t3WzB5B25u9nYj47Cj3p6OZMW2WrqcWBi4aE4ghxGah2bjqDAP1WhtRcN
nzbV96jWZSzlll9Z06ebVa2ZHJ20pMCt9pr9nq0uNN1rCsWKHhiW0/AlnjTJ
O2rscoc3jDWDl9D14+HvXgw1HlMxbibsKrr+AgmOiQebyqC+fRTUpGUwYOFC
o9H6gL6fg3qpyfOF4YrvhsYejaDmhOMpTNPgE3AZt9gw8nJ76taYjggdt2pA
2RF5bidylOkJjqJvr6isTo0QjbAbRkNQwC0vIzzgkyi+W9HC/cKrORpk2ZHy
Orsd7TsfJdRsyhiVAOhOOhD0huO5vqXJe2V0tBsANMIobgnljy/blmSZSy8w
bCjdc3EvUnd0wG6c6nGy+G7tBIj/4SHSuibvoLLl4rNBFxKJVEl6Rc/bAvFZ
ubQdek5Pm+xYEtGQP0wgHdxUWryWioFQVgoWWSh4HLOzNdMhVrtLATb91X5c
7ohw/rwv6BcyR31VZoFuDrukJWklcry4mVOySD4eKBlfy7R+vrdn3Yc4xBY+
XU7PwR2q7BmRz0hnMjmPO1JEAeAfzZUUqi268/uoFewDelowyyCsDYKrNilK
17VRtC+zP2hn2nuajK6uWV7pkTTf1WUQzTYtndCyHUcMgmFePvah3CTPJFti
6xzMcpzIf+aoSWM3YhOI7tTKhEELuRmnRBvLvLFuUPb1qH2Q572cA9yqaOvy
6rudaTv9a0qZq/YJzPxICx8ljqBfYFlSr9XHPrhteJeetvwF7hTmKEtZxEk8
/dv1GrkKQRWyBB/9BBGyerXhlhJUTQoMdy+rjo9mJ4niLkQpZ1LL2DzKK6hi
i7TrButwmltsmtMhhcKi2EUoiqinbN94/yAU/0EW7D92OXBvWRcc0z7qQ88x
U8ChqLeOpOgQ3c7WJFc7ZjfF5bT6AHVPW6TNyKS+iFd6droeAE+vve1e6/8n
cJQTfcxpmV1YTrP0aERM3p1sEArzgWNtkmv+/4F+v4vF8lpN85zZ/uZfttpy
R4GveJJL5+DfpZuOM9ItZNIp2h4wRqQMQsSvIVa1GLjMP/p2KWCKMrtsvwoX
iXmBN7bWMBATv5/YY+/UVq53zTUAYJrHaJ7/Cw/PIVJ/4dTTNCniGd5Zk53K
H3qSmdvB6q0+GoSooY8WbyojW4DkbF6uOi1o3BCdYo1KDMhXxb8tyIBvpq9K
3tttDnc8s3JId3KWwakqUVzuwy9V4pkNnqQ74Q+DUZOkSuW6/EPdLU7ewAdc
PNT7f0lFpG+YUohy5BzF+8yldrdE3MTEtMYfkm38+QX+vYSX4StaAnlmcZCb
hTYs3UrH4QD/ky6j3xEbKVN+oQ490tIK5s9FHF2Yv9u5+jPdFjTIs29ytOKi
V49971m/D10p1DlmD2hB4rGD4e9L0x8YUNRrl5goEsmyV2L1ieEKZekfJqcw
7g3MPGoh09dZ90dQ9QZ6vMF/nc/BftDHCRhK8aB1cJbQKL6WQQmWVFs5f1Fa
dpA8Wh+9FzEsfpdliRM93osAcY5ElU7cs8DfWYfCWGN26XjUN5RHf7HMhVZ4
wQKGKiGqZlAm0zf4peFC34bqc22QhZBG54VXNqYyCIl4mHPRPbSTJ1+lawJY
KLbRI+uJNVbA/RTDU4TKBGTElSMy4lpDTPytVas1L5v0HTkziZgmeOUeBXJI
r4GMK6OgLmgJNI+bBGtCq+W3MOP/W/mr/aDY6mkNWbWRW2+NvCBpJx5Xs/e5
Q27eHlJqR5buUAcqrZV2yyfKfaiaQLhsQfgF1yx9GdY7etx5GU76IuEpWeJJ
DZu9uLrMdsKGWxEcbQYyCALmKUdtDIbJWNtjGwaZgNkQzf37qYMeKujqpQqe
cR3L6MFvlmoT+IJtJqBExtM2uSMUDGxLJ3yVJj0XS6aZZkpRWjeCaYhu6OO8
vn8EJYfCn4Kxb6WqA8yCsRY/F/FVxDJTa0U6SoZdTJvSdi2p8e1jOg6+5jAe
zGJaAPFH9Y5SsVJvcaSkmmETR9b6ahzyGTI8qvFFNHiV1WsRpPyWLK+RBDF2
ezhm/zHDMdnvDlnQq8/Nv4EUlnSy2SMnWdNwEvs+dBYclFadtRSIm2cSGs+c
kPrCdGPQLCj7UUvcIPkroCUWsILzNFCXz13B/7QYHT2Z9fkUp2iwTykc9ZhW
jXTKD/i3RdK4QGrMxQgiTmuUEJZc9iEfuJj9TLBFBNBVOFS1gMi9m0UoapRR
wdUWCQcRxjVGSVGQDgMlgAqc1jx/Hve6vUm+jZXW5/aFZQGLZHrNLJ/cHHX3
r+AqbGUyHcBV7uYGUg4JG9lCibU2NKsSddcivM2e0wXOQ3Y56DaO69L+zpQC
PjQ70SSXVDVGLh+xSYxNXj6+UqWZeMm8n9yINrulLO5cBXX3gI7bRRoqVxF8
RYZWkY2XzlPtKTRed+3IvSXkD2iRXnPlPDiDto+xsHWyGydaw3AG8tqAi4le
Hs4LXKHCBG93GNVMxaAiDKt9XDBbAWrDT5zP3HoVUIfW5VVuTx7yvBCfC0Xh
rJ0q4epdJNtugUxvmRUR5GfqMdnQzUZqx8aab5CTknVmNaRBHc2XzUjENVt6
pMvpw9LWo+XvKS0FRGRZ0YfMx9jWzisp7eliB9OuGvNKBe3iDVa7RwkjFuym
gNLNv3x6WhH47xXmwk5ut6wO2Q+wijOAh8tiA7AKs2NeoQwFdaLdEnVJC64D
joVWD31yRTDaB7nwfe0QASJY2GAZ1R3O7rwv7ijJZ1wFt5UATP73m9lwRxuo
w8fJOrDp5BQnDlj/wIl9JC8l5GFGzxIjF4NEkCgp1GTxfjMSFzBMK/A1YUUy
USv1WOev0Oh7KQL+jBxa734OHa+zQY5TVwsQZ8DcCq9Uyum7Xhhli+JGQ0xA
qNwyfgrbd+mZ2baHt38F6CcsSRdq39Xk/UrsXMQv7RrUcNsJyT4tLFhJZjEl
RELewI6h0DERDNLQqSffejAaQNmeGpv2kkYJY7zKKhDMruUtJ5q6h7aGwlpZ
sMF7z5kM8e46kplqGdlg8OKZKcG4N8K4s/4Bjy5+8hYL+Jjvrw3hb03BIihG
R7trXi7lvIe3+bpPrUPueYHpZitWDxmbzlhHNLCpsDUMYd5Rd8cqIBmv77Ro
CrJE0RTR5lgRY4N+HvQb2B91nCq+/YDtidjBZ7iDOwkUIPmxolvH+pH4zESC
PF0dKnKVTgXG3WAUcjHHWRfQztrd6dP8SfUTYjKt6B1cVCV3Ny68THc9wAbf
WH+GDCDmUJxjR+nKcO8GRTR8MMGau1QbNdMxVpAipoWkLxrDE1tsn9Lbzs1h
vGcRiVbXi4DdV4sBXMsvNCUhyDWXID7AaYpyyVysq+rVikGkJ3pAlzsiiW0g
faVbSnitZk7QDOoYRrMSBY+lFXlPrL5gG/0R9CCiTfa4zhhqEIDyn20AiIqo
AGs6EXH2UKS9V/LxA3h29QxIQUyV3LATNaNiat0nM1LmbGzouPeJdwwWUqic
kaRGPR3PFn44j3B9dG8yojH1gDEF6f1s0W2p6ZnaSvj2rPb1i51lHy60ZANN
srSo1PqeRU9E/374ReqPY2AWbKxU+uz1h2Dl+AyG8lMssEpiLcCTg22lBXuB
trJOpLran9rf0b/fcuNJtUjBPdM03uIkcvY1cUAK0z50Vw+5l9bfAAvNiOGF
rRxQ7mTYLmpDGve6hYr/GpvyJIjtQ2eJemEkuQDwYFh2KKZ9mwRO+apSfVFi
XofAasXDSZsspofIK9J+tuoBLxlmIJkpBqx7neXR5rGo6cZtiWtLR/LkHNEM
2F92Zu5hiaJ+SsyYa+JsfdtXnX5I3HcceMiSU0ntHE+6jhcqIC55EwZ8LRxA
K6vHib4QENQlXZY4NyJz63GMYxn7KWpMA0jlxILtuQxkhRSm2gmxsGG2h8Gt
gnvskpsDhb42PLbjnFK7MUIQwieDr6vYZbzf43aXKdI/itzepg9DMjz+h1m6
HValmqdJFluvvAKGrQMKUI8YrLjUAuQmL+uhXarzv+GBk+zzAWOvz/SyVEiV
6T7OsF5dkJHgpq1JSHZNE17qI2PTZFXA0tn4dFoV/BATByyw6G5pL46+awMu
KY8P6CFY1g0pBT2O6M2pXqhMj4FgXFsfyzEcMZh+PW0Pek1sOwg0c6GMf0mV
Z7gC7NdPjCJsJk7+UEoaDwL9bMKO3iQluYgxVqpDTLr/Aq/hMpDnmh7hvp4b
NIZ/dtpD8aYHJrpIdwb7H61RmMxYuBZwl+fPy0mRXfAH/eA7PCPNOcNRx8US
0l+Xh060UIVsNYjErdQ66xcz12HJnqgD2k7K5PTx2lTWmCbMDgYei4zu5Joj
yeLeBTRo47u22ZmlAlSCXqZhEr0eop8JHFInAkL66ZzwFPSiXFetcvv6OGOQ
3kOt/N23J9MB/0cv4gz3KtiVE8iGxyxtcGb1Cbj/GXbIBsVHR2IM+Y6IOqqQ
PIu8/DhpmbtUYYd+Pl92U97CoAaf/FT82UPkhn0b98GKtQnG3M6qFfjXy+jV
WlcBzXJT1N4ky7TWSQTkxNu/cof1AtkpeLiY7Ema8YNRAfZvQk4wppGwUs/4
Un7pztkC9ckeK4SD658zLOVQ2p7G6D9vCl63/Wy0Nbrxz44tibXBflL05qzT
tpxCgfSKMs+Dshzk1cuvzvpnXHVwnRZppT8klks7CSFnUJyLMpyhmtxAl5Oz
bu/3pscsZi7DYlrfWtM18UC/nlLlsq7Mdg1MvuLjhTnKsz50tJ4fIL3092Rj
JPqxDPlNJMD32liZreTglRjdWkNGG5aTWuHioO6w7PxxhCl7ptChuw62aUh+
4heKtja6+QUJ6FfFDPfFBIr4KpgjxXVygiHak4dPWYjR3SXuHpyqn6fYQiQT
lZpVA8Af0gfdz62BiSLaD54CqbgvfqxgAnuw1dZyHXfUuCfeYZ3QALcJLpwt
R1RetLOg9XLLA/owd2UGZkitLfVwBkVkkQFKn0nCUtAZNPI+KmK//PINtXMd
AvA2bTxByNm4XVp2IBUcJS/EO0NBXLbl5K4xN/TEgNNA7mO1yXF1BdkIZhvr
r8eBR5s1YItQ8kMD8oMwfGdAglgP7oSrVXFXkyeLEOShCfk7Zwna87X1MWrI
Pb3ulkOR3xl67gBQujyLB33GG+NLDaehtQ1GBQ7ib0gW7jYSbwSMWdTEz9AR
GLMQgc0WEFlk5q3EcK8VnFRDM5Vysotqp0hqGhoxCHR+G551ZMA0f6PWoFyy
s+p3OQgCbbV4++mbL/YrR5vZY/TSfCavlxOvyUE8aEnFDx3tnMNHeXyd8ZSZ
qXtNXlwetmvLUlhE7BwQyqEPz9fh3R2NIRJ31A4fK2mMWGC5jFJBXQMk3ZWW
nyxsnD3i6FB73o6vLhJIi7cyi5HBjqik3qv6zT7Sud25bcMZqKL4/Hayn/KS
b4c5DXUQkFTHub0Z6iMwE/3GD1k1q8hSdV7EaLwkol55c+xwNxT9Y3GocJHG
C60bXairu4ykgMamvdWZdak/VNe+zjyRWbwMX+Xvd5//IEvpBgd/VusmrIrE
uffpsfyXy8LQQGa89nWHaqJSqwBUiTo4ikBcicgCVn0DL+jFH1Wt3HZv/7FV
SjCJzPQcMTcKgFgm9+FSHn7ZP05m8iKNmzlctoJCbdorWc53c9d4Oy+dJAqI
kREWGz203uCZeSos4CvLJPCFe5FT2uhvLzERoIRn+mreTLtYiG8yAEeumVew
nQS/cJ9hc9II+SB/8kJJNMuCgW81KgdflBIITrDrwYGSTTTArHbQwTL51Esz
B2LEuIPBontPhiYGmPimvdbDoLRXK2fYvGRuQ1VOHNBQ2an1a2XAH7One8PT
eOUj7kBTLdIfwbXD+NW2Cyjsqw2QFnK1cAzgc0ar+RGwweFinKW9W062OE2R
g2CLcd+hJCQVSZmSuZlSbn1nBvoAT/8KBHevmAPytLP+gmYs2ntlHbiCvO69
8EznXsE4v2mHb2v9x0eYTirMGUW4gigEtU2WOjiUseRMZ7AqUqKQSmkkHgR2
1c5IQzN3S2bwGJvjMhezkZiovQXo0OkMi52YqCEQAPWVbICCRd6i8BKDp74Y
+gl4IsDODVmiMlgHJL0RuUioTJ5DiG4oPBZtFi7RygDYhbSuRWzpaE/0Pd1t
t56xAcLr1pAyX+lKJBE5nokHxMcfc/G5o0D3SZ1m5qFS241C336pD11hYbV6
19EOUnASemH3OZKj1tNOnVeltC0FaloFG9zCaMEcoisywAexyAsVjkOSfXCJ
uBgX7BKY4/EPGhJwZ0AAFYMtjIid3fEaQPgsufhP26enlE9aG3xb7fhC11sJ
V3c7jtUH8d5IXBg4J2ar55lVwcmE5+quvKcx8UBdYft1jVdx+m1INwM+lPBP
Ugpo+vDRnXVI2ENI9Rw+/UQV3WAKneXEqLgstFNBYNM8HSxegwkkUofaX5TJ
q1kRbr8WdX+eI035hd5jV2tc4Qmsd02HlyU+oEJ52fpxNr9wQ8+ntrtSVYMy
0l0UjlIn6QzOTdEH/95oQGQH/2xgWS29OQmpjYTFNm72p0aHvDrjiSpvBVDM
8hXEBK/owQcyL3g683ZfKep+nwq7Yvtms4PJPcksqK9ZLe8XMTqnIOXxLQcK
WovOvWKxGOF+EwLM+qxmz73cUycRnrQImoZkWVvMwqDghZGPml1sQ4WuibDI
RDLJi5brkdTmDRPkzQuTe2KrJrJbU7+ZShC0BsIgjvWMx1xNCfb8IZ1wOBRb
jm60JGZ/vCj8N1O/fYbieOzHK1GPzJ0ZAtAnZ1V5Ep0yxYEdOzO0tPNmwG9D
E8MFeQhE9LnYvaC2hKBfQoLCRUE5kmxBESVdg3Zh2neDmHMBNkyH9UEf624G
RkPPrWFD/qbNBZpdBZHnhlbkVzvbNZiCb4dzRcVtjoKjhn2iw2RuW/EQzbHp
AL4juqADax/QQMaTScmhPZgf2PaDVRyIlEvNujHXD7lhznzQzKVMZeSuTkaK
GIUhV6p8aRbs7rxV8hrXHw3YZtlouMgobKi1/zsd3ngfJKE9S2UHcqfnx7qV
zeda6hylJupsBmpFr4+9rfffR+WttybLUVSkOennpvUJd5OoCBrP7OJc1mhH
BSxJBM2PLsAdHoHEPy1Mod9Z8dfnriVDDY2kgOgy22+c4U6YIW7iunzilLo9
j1oTBP5K5OUyX1DCRJEclomSxqPs53S6LhFr509eYISysjW4YT8oHsHx0WwX
EVP2BHX0Ay6uTKONwPz1xCnlYnCZv1MrCnDMiBl5sIJShLyG+Qz9Tij/zwVU
/7bMEisv5tigln0PuYJ4oeOm5hkGvngeXnboRKPOCnTyqovme/VTqVQmqGF9
APjhTj45g474hjY9u84i/jabFXJ/lScsFt94JaRlncdpS7pJWZ8HX4rVUzTT
miNQpXZkQKesm/gS1j4uo6rJkkBr//YHEUB230GwRzm+eMsgJ6kM+ESrZqtM
zb5gix83I1ChPTy/R1rsqAb5hiuamThgNTKlBbVv3AgbQpeXx60zToDtuSUM
btbxyd1IAzmsDHg7v9uwlsG499kVxSYJWMlx9cWtMw/do9W5eqCIi1s3neCG
1QW1ntWn9gopXTexg0U5h39rYAwegHqWtbD84pqucAp6mO0QYtuWUseLpQ8p
2AatsTxc4wmWReR6SUaLsDigPoGZn8yWdc6wI1WvBxx4E9FNKrgw6IYEJaPU
hIo1yFvmlH0eCxBFciuQJWPAaDfB8MZny1+fpLcKXltmzjq3WqJJPkvU//JF
7JNu8LSNaFMiTHR7DCL2EnWNLwxTEPpIMMjut22GavrOhI32RbBacr7y7CcJ
7pZKcHeF0nv0GYdS1/3naGsi8OszvQM2P5SGCzr/vSHEdXgKPoOaeeWSv9JO
IxetXmZOT9L7bsJOtTPMrRuCJIsmMqR1BeUOOxG168C5XelB1fyEmc896Ue4
Y4LHoalFI0LczR6TenjgKWHAwKdGyHRj7ggFrGeUbZpzjXmMlvB7nf1vSm0L
u4i6JdFtdLdLXk86x4x8e3BUDm6roKsYE8lt3u0mvv09wNH9jx+QrAtCIY/b
NKr5y2CRKhZ3JXiSqUhVcu3jqIxfybPSuohQ/Tri7fzHom0JKncOoC6eH+T0
ATX6OuPAahJ6Zj9wN/V8nwGqKh7xrN/f9DVp3BHQVL/vhHb3O1Vw4IiHDIW6
Qb617Ol5XaG4x+XANzsLUS/5m+3nJbYjXOtRK9T5jRhnm4+p60VZwduTSV/J
YlPFVCaGAzkk9r69SpL0od4zhqbHx5WVkaCNd7IU4PuK8b+E7QM+FjVkCjAT
46ZD++ErWMkVrn3Vb1J9/AhYEabnqSn6vJMtp2Z/KZGbP6MGyG/4kof5jUx6
C4d7RSav9I7+qsmzsLBrSwVIKCkWtrCGTA1H+IushajTsCwihApeg5jrNR4P
LBMwBSdWHTEMSCFjPIRcDa3yuQBv7UJ7UCvYnxqqD8R8O8Z8cz4FgillSmga
E7VRIGUBp8II45YHMeGyHW6Y6gN8HWy7uy6tuZo1HsKQID97vVxIfP44BLwH
eKo337jytu134T28fme9+VDibFo8BiVGBNS82vwoOgBmJXu91tK45sBGdB18
j1OdvUFAu3sBpIajnuVmHwTJY/TsvwY/F1A9Q5Nfz8P9aVNtg6jmo5G9n21P
S5563fmDUV8HVGcTrSaSXdEEqqExMMopgJJwV+EeDpr0iiA996pB4kondtj4
cKOK0a8P2Mmdu8w31GcCA5uANbbst4mVQtq2mVlZ4eMtU00cn/zddONXp6so
SM5fmc25oGxPXZ/R0/oQbpL90glkW+jYGj8CyGRl+9RIsu9RjIgxU56iOou6
NKcQ2eJ8ZTvJ6Gs5yNTnlniXNaUqe4Ybc+5E9jG31w+LsoU2RAyEXs0On7zn
9jdt0TDdrmdFKu4XKJeGOa6KnVNGvsGVEx7LFZtQgJC1s50Xw1Mlz+D95/4X
xM2oG1m6aPF40bAD5kKOQwJnjubOvVxAk6EPBr4Hz/Oih8TEEVr15gRdpKL0
P8oEOnXtXPZvhwKNCQMoM/GdAJWH3dx3oe9FlOK3Ee26d0lxE6/h+c3EfXC5
ERnXgTIsMhG47fMgALQQ9F56ClaiDI79l1YbO/28mnVrLaDHMZSkgUXv0N1d
IjLJCmiUxpZLIXkWzNc/brTSDiAFZHMA4mRRwxtfoq0qAasXx9m8MdFGOaGf
CtirphQKXlDI6Hw0bmHvB0ydVHgTazeZoYEZInPuJLnhuB8gLPKKbVH/CbAX
R1PchWv+14LgUXepGXhQBqficoGBxcP6vefvcQehE8GC9xgdiFVKPOkuPpe7
7ekla+YxnMgMysyBJxvZoI1GwNEk7jtbacgFDwcul2/cBYdDAmr+3qfLfPQz
xj0Dgc+PFnmNbdCEdbE+OpZiLAhmSbcuVdx8moq5X28wk0BM3uSLJMkxF1R/
P8nzmK7NQuXlV4lJXOOBK2YEN3SZQ7oVIK9ayow4g2JGkNCSAdwD5YDQWN7T
2aSzvR3NnF3/8m6/RbAU8SJ0zHHuSM3OvAJhVmZZf8usdvNny8eigoRNoxbn
BCyWBlxEs5tdvbjOB1XHU+y3Qqz5LRpWLO5OLAe/TJYRlTFDEcha4GMQGzt5
l+TT+a0hQp7AmE5erS6omirIjv8O8INZHVR/lwqLMDRrHYcDRr1TJpsjmMR9
bn8VDbLzT91umwpjiidYNo8lxef9ggyrOevHOSWRSqGR4yDR0bVXTMe24ydn
/Rmohv5H6G61YpFqGdKn+ddsVmo5h4iptJTUCLTWQMKHUY1Xmk9fUdvnU1Jk
h4aAzIE1bLqanwhqQOCtX5sBXnhxxAin8ED/JzSxnFzBn4H2Q9z4Zq9IK5fN
0fnPda6ZzW5z9sYLlFsxTyOPUtW79AT708Sj9V8scBfGCHDj112MaVQuKfwk
tqzk8D/E1A+B91eZvHKUcVMhFHumE4cWNgQJDXFEcYZkmb2t+5yZYFNLLCp9
+1agaeG9sm8iKgGRh47zj1vG+g6Lxz7TOxdIvO4+8Mhhgz5yq6+0YMmU8IrC
Aa4SrufdLdx79dUBg9zJLlSoQ1NDGKBEGm4BRpHa1YT5y4VYHhHWQf8iEm21
XN+gpvHT8Zg2gZbiisGLSIa0XVtrU1iiRmMAbHnkgXhD7uPtctgX3C2nS5YD
iOdbgv+dNqfRyI90xefoe/uLz1xf85sQ0yj905H21MyISXUTtm6SlDcqMNfR
8uK/30ESxpPXBwqXjHZRu6egl6SKgoAbCbRj8Opof8wQ0STJ7/FE/MVc6mgk
IU5z+vUzpH+i+pCFr03gloDZIbJtql0mj1FqI5mNUUNjoZMkB5y3TJQZTFkw
s3FB6Gs+L21RaSNE37BrR12QYk3fcRxmMdaTgLzP1tiFcile4kAQotXOIbZA
7c2c3GNOMhAg3R8Ff24NaIjA9KbxY/ONrEL91zDHMydHKt3IaTjuoPluyvfF
e8MqWJsIIZ4rC9mWXLB25oVsIW0+sEZ6dEkjYWIk4JX+rz2+vD6K+uZ3KXoj
Q+mZ0YOGBwlhy1f/oElC45yTaIReZTrTvnitK3V5DcpqU5oA7tvd8xRnVkHH
cTGd8lI5JGerX/7JIhnWn/3yftL+3yNDhRgGeeVlbYSxv9SS29mtSh2jubYm
FJT+gyuXPDEnTGkzkh761z3UyDfCePtz99LVFwPHoRMtPbquHvPmZEYDRQyF
Zq8Zwiy45cWSqrckjuJd38+cqoD6wZZs3Q0lY2tsoqM2X110mFtcbjNJKRiM
xIPrJqJb8dAGt0NTEE85HSiMjB1BqLOh53FIrictOOzpO8Vy6cb7GFwlV7N1
o53L6SYeeHjhkQJlkU0DgMBO/q9SNyh33XQw5vfxdFTCix/OHKV8BICp1tBR
ElfZAHK9R0WowYWCkEYLkWwu6gMJ4LzvCoQUq0RJ5TvuQAQp9SflRlNoykGs
S9VsxnlUxNWWVRk5Fo5E5JWKheXLWPTgmkNMw9yWnyNA+tacnDF8DtljGW/d
kQtIaup/jG9XeduHmYecMfJOE8ryYDpe0RkLYMsN1PahnB4eILC9WJLL0Dzi
hK08eL1xk3X5H9LSLHZko/z9C74YxTiag7xFwCi4JuhatlS0rpaDPtQzrRAK
NRAOkFNiHAZVT+1FUkkJl003M0j5DjE68XdBVrnrxLu8PtSLd9Gnt3ZtZ2DY
FGywgxbc2bBWJ7O+/ZyXX+hUGG6XlHC5JupmhCeW5PPBelW7PTFr8vFD/1Q4
1pvnsb9moLm14Zz4TPiYYggxvCXbFAl11WZmO9dPJmHyksBseyYe8GWhxRgw
bRirZCyL0cDi37BvrOBQay70ijFk9XLIkNV2yQeg91Y5BBMRcycM5nCewYG9
kPLAez/tNhnNUXJ0eeMmcupTAGOhAb99Kbv2cj1jqsG375eM0cFijsQ0aI6a
KzOwQNEvFbntZA3Pu1At1POIt25EzxT+k1ouPn0++ntpXbwkrnteyxwmtmpV
ItOScfMioKA8vpuDbSDzqSWT8YUZIZMceCi7VLULif/GvF6nv+qY9+t8DBDE
Fh0Nz/RCx5J4oKmnHjiApz+kbyl7RT/8RoF8lbVum+QsI22tQhQdLLukHzF0
e/MGyEGCPbFrJBDGx0deYRlYFtdFJ2QJYQWfJb6LGueWSrYcVnnl8LE14/C1
iZmeSagFpmBlvaMpQ81F+fUUauPYxzrpG4Bi8WYgzT4/BJUgUcHKj9yUb6Ip
7x3Wwibj0crQ2uRvq790Bhby0uZSkI382XFJQ8TManw7P04o9BYBAeS1Z+xJ
bWuYzxa4Bz33gNxnUtV9TAWWel4v2zLNywcJC6WUocXFOmwwW9J9jYnmU1mT
tepO8NVTQyAm8crhC9X1PDY+19XovxhBaqVau5jVR+dF3wxuYZQMCe7Tie+8
vkppa85eEcYWEcUyCTUOt0Z8IMLJ1eSHTAs3MGQIIaHTUNN9ORCtn1H3tCbV
BMcJCM43EiQCmGifGidnZqTLVPU5lFfmrrj5o0MWsMo6FeFaRVgRTXzfh3K6
g4CPxXDRHGGfW/V2/yMdfsOhmmiAkzEwzqzgwR6x92JyNgN9ok7voFUaKnLg
J0DdLnTOHQ+BRzTcRBMWGnAGEFTa+OuVNXMXuVf7wNQYjX8BCph2B4cUYDpB
nXrWpoKBmtsMiK7mI/5lEKQ8BaS3W1VcwGml1wJqLfL1KqJ7Vw9c5ZKFQhr1
xTKgwiyrDVzz76Bb9wFSXVMbeVo5LaPmnw38H2MzMkhOjvvCYON7azLf+z4X
GrHR7VPHCH0OD8sqrZJMUjlZ8B9vKEhnGaNuMOILBQyKTq3WTeo8191SgyD+
3d5TVWcqCB6ZY+EPPoqvLlcNXAxrIknPN7DVJ5w0SE1Q6yiMz4xgG88tu9Ca
BbXvK5kXivDMAD+jT78DICcb3jyYbiK8qhY0oyIlLSaaMXQZgXPOiklIOENh
Bxg3WPB8OSA7F24orkFVSsPHTpqBoPG4Kxi1yCee15098Cvq/B6Zd+IiLHCY
0ppXGufBTJNljsTd7ECEHRUSpgK2zs/TlQyxn5WYNm+POdbJdcMUsCIgSMp0
yodFk6LtLxBvVcfJzxf9yrRn3Mq9+1Y6UpVNuOVfhgi0L5X73zypnwF/sV5t
A+Lu6nJWCIOHPvwS7Y4DqIuX+PHdsHzBmKZRiXW+yk1o1b5QnUnSye8xqVjn
67MubgTQ5A3lNopSZ8t8vcXJ8I5PhEeEshOLqXGWbPeSCOkokOcZZHLGxkdh
ydiciZyO6dYuhG//hsTbvTSgGOjrajLKmLWTmmJ685nd19Het/QG0Othm75f
zS/4P1C9Ih5UjBkJntQ82v2DTX6R26cVXeTGw3WnTyPlSycAVDXbJwAcl4T0
MJnNpzvdBgMQQsRXMXYScPE/UUPywqFuNeqW9k6xu0ol7LRupODJUUyt5j1I
WJ2+Bq4GGfEQKJzVcqbMdsZEzstnEv0aOSU0QGgFycCGJsVo4fcc/75YaUhY
t9VEYk9e4/jpHlabaFC93Af6NGgkW21Zd4W0R4xM3u6z8MiRWxiUBo/f7Cv6
TaAzPve6Ct0OzG+WGVqCIe0zvfqSGgoI4Y2VPEgA+4coYH1zEQMdl6ZWlG/6
oir1ChR771armK6WouFL67izjpsHwRwrQZ43E3oBbImI6NgznIlj/L89EsQC
fw5YT/yuQu7qC+NdciTqYrvLvlurKmNDYOOBbyS8L5eS3zuHWJKq+ygsq0bk
6gWZbykwYD0Wk/tvNRP4eyBXCU0lDiPm7DqrOa/JHurDgry1WtCbffKHFIoL
4J9gg8uYrZZlcXXLiK90mTjW5U+2+d0yfLJOEanmJnFKzwZ79NUVUxWbpL/U
C8RqG23VYEIPtcanaSaBfFqE5/BzRz0t9MFYz2IxpVsUnVXG+DECE1jnLtAq
p5vVqWfnSugXEEVBIrlVqgtQ29DDzXTTmDav1rbjMUsA1AMJxA2jf9yijhwt
QmUddthKWlMaY/ET4OEydCwJbtLnGvjrN8Gyk9rcLEoNsnYi/JE+2snO+w+t
DvjnHQz4Nw8/3IJJ4Cmj0kNKn9hkF4yc+/NRAmQWDfiwLpdbOp5nSbjiW0dG
cpDI3U2xNszks+U7bwtc6cZIZuQpsAAMDbUrzHgf05AjSPSYYIo0PBQn5nje
0RRKgHC/uRnox+T94Ow/7hdC1Z+owmCFl25Bpqe4IWAVtt54Ej3+tcAex46P
7vvxsWXvXqp1s38SgzN1+JeKWkL4H5urPzYP62z1qcED4utZzhqhvgdALnqV
le3aBUz/4D2iVqUrDGN6aBA9ddE17/BIWOdR4Hq3fQU903GDvQDFl+6bxN3m
hepe7T7kr+DTc8lUuHind6S3hFCsp3AmmdxJyNWWfTB9sRRSiATfxwMoOd8J
zqf0B21ka30u0qrDfyMl1Jh78ogD4R0w7pOX0aZVI8zFbUg3btSFMcd1zn6l
cWpcEMnCP8Ca0qxI/1lW7mBDyvwgMEnXmqvYCJCXbxyi+Q8ki7zYzX3WoFtP
y2BaenkRjcV8JAijZPoGzVK9HHP4aWe/vww0dbS/hjhTBhIUDkOe+4KalEMl
+XhjfIWbYYYKaAv0Oz4dlIbm5EuKsriTsO5BO4peATHVqWR33ole8s6vMlsF
4V8TylsRoNddA86+TWuXuueScGbsb3iLSoes+mZdY8f+kG3x525t+ZCe8eh5
Z2PbVVWwYdAUUHWsQVGvPmnasgSPQwVvebou6/fwNje5CyoxuSAeTjwz8/dT
/X12R0KH69WhFniRfY+pPWokJdYVLWMqa4cgXcXnepJTJJtYsgWyXzYkI2FK
enuFZU+3WnaviXkUARAWJr40B/BMLS8FiElQqpFL1dE2eaAqS2ijZOMipCL6
Ar55+Kg/WbSSVtTRPuNOXVkkWgaRLMXZiK2/Atrqfa5xjh2X8t9MHDrA2wJs
uZomvnFe7rf0rovgVbE4rPCqNARJ99j00SaqcBBu1QLV3Y9wbG+eroJP87zW
DNosh4y0wXjZtMj0qmYKDCIBSwMdAa7gFhwdkvjIxweJ8d1C/hqYylTfad8T
1rdmaBwp5o0HCdCVjhUJD2G/7TdJQOZzBPwpecejIeU9t5IEzzvX89e1JV7r
lt4kPBEVN+0BPNzu80B4gLTrnFcG96HplkII9wSFWmHS64VHNC/CnS/lQqBk
fipm5FjnShKxU/QJdyHIFNuUoqatZ5ENJHqlKDzDjphuXw2F6dQMwQBWl8df
p/Yps3d3RLXzWTMBeD1Rkq7fpVTMJCmEV3+evM8UtexHu0ojGY8rPsNAFnW2
FCF2jejxVK1I1w7qm/SqM1OvbTySgkVwgmecuvcCGtSe0yWQcGOob+hMCEnP
erQ7R8e9NwEtP0exJdFaPTcahxuRr+KUJkcRMX9P/jhNb4zhl+aFw9nHanFL
mH+UxsHdN7KqxD5cXCAzmkeZk1sFcIsacohEVSxPmAKo8q5Q8STmbbJy86rf
Uprllql91FxMSd8McOfC+dMKXY+hkVt0ij7TNFf5wk/Blf/9MRW3+J3Gf49f
QB5SkbUYlItko39FokzbzjhFNhijvsRfJuxH4UPcwosgKxe6vBONyMrODzuQ
0IvhyDW3fU+g9D8L+XLX89vMth2eC1PUXLvsHDh3U7JYW1hFV8sQsdmjJAol
WDDmooo27pxmZ7iZ8U7G4xM8I879W/x66ju9T6xRXKqStcBbOQsStCHa4tKz
TfoU5uCvkAe/FRE5+h9S95BCe65bqdOR+NWMTSE+7HH/h9c/Rv08EKIak4EV
TxZr7cgPgVKixkikgYzjbxKpcYb9Tkd1I+8USFewiJ+ExeMOb16hjDy9YDW+
eBThRAwPu10kstrOPbVBXXauJQylGvUw7uW/fHe/7waA28TUjDPGFnJQlQG/
Q5IdFwkEKsv8K2g6nE0i/4v/5V5gpsbFS2Ift6sUHk6lCXEuWPejm0Ic0Vw8
FK7sJco9vv42ZbQSd5q+j0luf9lpfk3ZQVqcis65+sMh1m8ntJg9UnW67XjS
EmlI2Q5gvNoUqgCbWHxmk6osZ/mZaDDxx5uo4JnwqDOMgNum+rZtWUX6/xqT
KWRxciAzShS/i+ZFU45bAS4fcmcAK7kMrnWcdA6/a/3T+fhtrw++QdZWC6R0
g4Tjo2lR5JJN6o7q+bXiOlah5j62BPLqhfEtTvdL/GZZw+gneOFoA46xYoEM
f9+5yTW/yZJCp8bhUaxIZcVJ+vkhdE/FUEtMi6KsgZyVA40uW0CVVALfmnk/
SbJ0l9BJ04NB9zgG6dt2Y8CWhYufZW1RDvhOlF9wkmt23Kg3qGC6QKUJEJri
l1EbbJcb+Ezdfp9gZoAbn7QSraO0bhLGqN2ioLA/CIhVhkCwHKyhrawzqTYw
y/6BAkEshlVZYJjbgf7L0vJHDIwO6/du15/dxzp27NGNER1GCxEmqKYlBJev
dix0VbIhVWKmgkLn9iJ5KCJsn0MtGoAD0yQ6PtultV/3xxVagD3UovCDCLYe
w2lVu3vP5c3ryFTuiW5gbwRPixzgQQf/BgDTzhpuiNgvzovJIMHlCMK1VGMK
tGdy1FdC+S36s9SIHMdjECJEQJHsRbrjA5BAXfm2YkWMHqaSzYvO5vg8NzG0
lL4HpXn+m0xVZC5ARV1p+ot133SOyfHsL1CCIi0Pj9qAamQ4hkrsGRT/6NWs
0tChpk/y5xLMysnGBwOSAxk0e4IDb4eEMIgoLsj3cpGfcDkstAcctCGSDebZ
beZfSXIb0ccrZm+DbaVI35LwP2iTqjrPbFS3rB5mmsmHvd/DHea6N8JYlJSX
gkiFxRtLoyRFb4K1SVHnhPvrztapOE3ZaD2sRk4mzxkF17AHsK2bmWVdqDNh
EMTwAC36hbn3CJx7ufRk/hxieP21blLfpGSnyFx0xWlpSbVnIiuzR4jlvbZ/
hJMHZKe746y7uwnwnmofuxYl5v9BVfINzLkDLw/9VE0uO8QLN7FBMVNk3Ku8
kFpLQjKMBIorZIYtO+KyklE0Z5b71+qgoB5SOa5h0O0xwjdiK+KYJ6ead+hE
bpX/bWcZvZIDCFjCSdvLNidsBO37sKb8mxWmx3Co46hekVA4pQV06PawfLRy
sjPHJrw8cZcv1kzymoztHGhYyelanaTm97DTia0KtvKwiU9WfnUuabWu/juV
jG4cOFKJMTPZZc1gTKKSRYpiKpOw3YxJQyjYJBfh+WGmVLjRSwXsHTBJ0WFb
FVmYQfNmOh01E9PRTVNshOR2d8ECTwvxqGEyzFKYdlEWqdfA6CRgVpIpvjoM
2sYLRS3VyhGLFZCNXikT/M9hJqsLqDzHoERiNMxU7m9ORfcGumv7PMGYTuj3
lFhPaH4DlSANR+PCf/NU9N+6a8APwVepvvtA+MDDA+GaACV/ZHfd76Hmbv6v
KsW09EwJrX2Coaoy75btDMNOGta5eWTfcN8JlDOZa0sXjsxCEnSe+/mf7UjE
7PjSeVJTdQHd6GSllcOOBw8cltbNEi2DDnLbW2DPDsILu60AYUGlWTDGbRNS
O62oim4a1iIwZjF9qRgQlmP/2igJ8e5n3SwVLLOQAoQ9PrlZl1ty9br5084j
OA/sQM/vDJMdUyonoeTcszKnMuImoJMQfzve9efSyCa4jlq0ir/+KUQYyW5G
h5c/SQMRj/M6StMHfWF7zagnvPjCCJCFc/o893Br9E95KFbsWxRRXNtk7FOv
a5EOcaqAxLNN6wshGBLWs/pQ1adMW6PLF9gRCqaAP/Cuk/rmYFr/YUG6nMFI
7LZiFMgMs32GuN7VuOOcWtYuV9sqaVNtApc8r55/KUAlYwcZboB2+2o8smi/
4jxPAAeRYvRwY+q2Ddnq7AYgZgYAvgc+LNSzreEj6GdFQe4+tP7f1drk6/yh
rAlRenla++btTBeXZrPweESUyNBmUTCwz78WMcCsG5s8nznxPa8gOLm/vvkl
SNPBUukmp0yqy24e7Z1bZKC5fiwzTJGnFIh6dJnjCMM8yB3CQG/WtERD7ezH
ypPrEiI8ngzN2DdsogH4rmBNzh9yYaNxpZsDqKcoKM3nflraKB+gRLZxZikr
FmHrTaoBtk327DtMqmuJOzTkwx/q35D+VKDbDrfIh/sFtB/3jeUwTCS4a78j
9ZHRUtDRx5FZQ1830o0CNSex/+ORI06yT8J2d3vA/4vNcLu3BpeKOBCmrws9
J6XSK5P/uiHDupmL6POElNRMK6I1UdR6W7Uz7Mql973X1xLspfFWwru+o/M5
xcgCd7tNNcSQ7vdLn86Ks4nljq7UHP5Vb8sXZiuVDdniX84t57ybjhOkg6ZB
2ueIlp3caweGCLR6sKdWVzmaunkJo3sjcTcWW5mMM/e26sevSi5AKbNiGbrx
SyWHhVTd4vWuKr/pSvUUpIAr0c5zwqHi+TzOVTuZ/silfJry1EDBGjPRJmpu
0qxgpcjL1KiDq2qtJGpxgYT2cT1czpvexCNAyhzK9ImXKb38TOuIpcQeeGhh
xOwfwQ8q1Tjmk8HuLF5Es5TZb2c3Xscsd9NAElFyO/KboU9CNDwOJKOic0H2
Y+nYjoAV54ynHZW7r0xSfyXVJ0YPL2ypJrsvMJb3ZdG+WbfqiDmy/xWJTYvo
AqbL0t8All3LFTppgLsx1stbK2lIMVB7wv952yelZ3BBvtHFTG7/tMVxZOjX
xMG5jgxakBl+WhxqmSzZBfwo5m0MjvGn01QfJ5Hoap9eXEJT+TyaTt/R9VQN
gNS8cKrAKpWmULWmst77aUFPJjfAqt6rp8JVLy1SNeDTrWALs4hEJtact0y9
pf9oTrs1OHESi5i/cedlLCKYbmHtcpdA2Bnkl7OBysSij/IRsQxQK4ShF9tP
fbYumfh9TyjdUQgAyB9lCy8wZnaYDfJKWz8VT3v5+aOsENrzUZFCtpo7fsP7
E4itjLQNWWdShYvq1+wBDxwR9AjI9MGWn4BM2zV3qKA9MqyPi4kscS46B4Ed
duhGz+alAIDqao1tBSKVDCI3nQCS8UmzU23gQOTs88BNKp5Mkrauo0noucpe
zo8b3jYa5Lj6pehy956hcbCncqShyZ9+dwERYNAiNUeSVwnbHcsIcK8c6AZ0
mGUQjxm/Um/cY+oATa8u0XrrinBX+xOfX1eYhZp0ZDjX5F59DTVQ0rbv2r8I
8qTtzY8e1pgQWmP9qrgo6rYeU3/2yis934sQ33lj4wC4oBzNKaXsyzHPm1EO
tj2eRZAnPXa68Cn4XPGtrCIa4XjQufhgvKvALO+/RRaRTJ3OHde1/ZDViZ0u
Dc/g9s/YgtCOKe+fcGFXcQuIk9byPa/to/fuc5El3vD2GndZpqqr2UthV/k3
tXIy1T6tMZzC11RiCqzPhoK4Yii7mpH6NGHJO8zSlOwz4GvzZS6Tl3ytIg04
9esd5b7+ukD9l5X/O50ac1/1SFOKveyzFZB2tXhX6mcDrwVS3oLH1c0RnaiU
slyiJKslAk3a4IlvjSkLnQnazQ2iuar2Zhr4NLsrRik+tIuSXBpcTBdIT9T7
veWAb1u88R25botklphT3Q7LO6mZwf54k6GN0L18ZFqG6aVZuAi4Cymahoj3
OgN74RYksdJVjgxL6z9/iDudvZMF3pFBuYLCJs87Wr5DriRKX9gE6IXmRXSs
+C1D84FbY2kQ5SAy3mK9Zzpmp0932r/LFsJyz6+/z7NHUZITI8ciE/Uchm3T
8xcoJyP6SXxHS7aKnVR3xfmOriCv3LBHnu+xR6fCwdAKDhFhvgZOh4x9/dyu
LMwu43ExSqyMMjnxezD4Egidei5NCbYfjbnIl/hbFG+BletpToASCqyWyLKb
34Iaitm+/bOmeiX6MO2UIHNh6zxH3wOAd4I2nxhnbe+jbqC3PZYixBttBubU
78yKpoiNkV9nM/h/Qp6HQMvEoci4j74uSHbt8rF89qH+e8IzxHcnOJ18OiCG
1VBZR58saydJPrs69YnMGDe2l+KHpze1GBjdTrq7HJU69y2wlAwQzxsA/UTL
KUz+kWKgSY4opPPhSjHrM//HZLe3t3s6geHJmmASfQz5E+IXzEvwm5aL2/x5
j08uLF8cGrTxRt86nyoafk4R6tSIHChSN2xyyZyhkDzCRtVsAPrYUHn4m0yZ
tgTKGalFA2dwq0I2moQ1wrQT2VtywlMI40Lao24WDCvSOc8P4WZ6NWYUpSfa
UC5HcwMyPpuPwipvO4EdKmYjc2+vbOHXiyJH3PHUZcYs08iuK68n8ygR0sfe
OywMgEdhVh5TCY36Mqf4BLp2FuTBJr+RzZeg3TauBzEsjBGT4E8sYvNmiDZc
8mcgbGQRm8Mua5FmaJxLLbN59HwgH3B2HJ69d1ZyZk9FeFuvs7CtLTFF11UC
EPu7XYY2dJwKciX0R7yYxppk+3MTINF5sZgYJyBgmbnaV6aSta0MAtpObFVl
TigSMlUt7F1DBKZb8vQjrUQZYBfzUaHAwDhKyQw2DNq8y2zW93yLA4DHcnEF
2oic69Udqxbd/fCF/UyuQuozcLakVWkg5hQkhTOREuWqKLpq78syxYpCSZTj
7jCnfZvBbJDI0VNSjbvHtitjn6h2x1IKhJi3tJvahovw98FVAdLt/lUGVKuP
gC/PRU+sbTCN9c4LZnH4HgKtdAtENF0adPjU9tgeP7t2cqTetRoQ03pHRIvb
D4JFRpf0B+sP+27HHfHMBvk6Qy+JcBPIKkzYm4pMm5z6l2bWmU4xRG5rDhGc
l17q9aTVDduH6JF/NptBBwp9x6aCRp3UsJsPU9xXL3YYuMLTOaxkLDVstHWE
3/C60WdW4AmDOvoVrsBjqwfktnd9KDtFM5bh/BC/zZ7Ybxi99l5EBYaUq0p2
q23gA9DczSFi8zNkbnyX1ieL2kSuuGLwjBnqOnCG9TnCJw4aESJ0gpH/8cTt
2ZXbUy9UJX/ox8gUoWfpwNGZoaSPFFoFc/XrdJYe5Yk0c5fNV/ahs4Y/rJmY
4bb3EmSrDTPRFdQo41R3Fu27hXZLzFsVzAL3KY0G+3JWYAkR7XOuMvbaMXqW
y+1GQl3xVh9pQHvYlEy3Ov5QHUJRX66c1chqgzovTXFjPgYCwYF2hUjmEfP7
gOAgoCXXYhKuJYbLSgrfmGCKBdZsROqJckqYVBYSP9e4gfmbMmQ0mv4GqRdF
3Fk9fll09Fg1TpKxJGeifTZ1jhinLk0lZS8E3Rs7meWtZbv7lhln81aqo2mx
J3gzhU4YYY0VOrIi3Zp7CCYkw6JB2nnOc2VPX0763T3qan4V1F+11khdfwbY
Qos2Pqfc+yjKrdWCOqj1tsVesU5O8GQaWNnlJO/2UpBFToK5h8tGeHvD2evi
TvIQg5Q5Qv066G8hWYystgA0gfona8b1SUUii8BTz1JXG4JKbWncX8Qe/qnw
vPgur/0M0mSrS7E9X8Ke3QDNyUoaF+Uv2PN2kbHsRHy2vh/VBvbdi07V/lLj
XrYumYeVreDmSYsJ+nKSQws3F/9zsFecNsyx+EDUlZuJMHSV4UfvrhHUGvDu
y+p8yXC9hnrBw7XTAuxztV5Mi7VJLadrKRrPQirWKIS58Iil7jiOIqf8UjaU
Ee9oqI5zTZF6ZdFqTKb5ud73hkospZLyfV1Co3HyM9lW9LEJ+DEI/JlS4Zd0
51Ruu7IOz06NNKhCEpaJ0bMn5a213Mw1+1XqZGTmBqiBQGfB03yJYoEDeTTc
ZYIdk1Cjrdmvd8be/rxoZtmetIeaIl/4Uz04tpsfohPLtpY+t8AhaJscIFh1
2IrnK26WPZamy253z/BXUu4w6wv96ebB2PJbaVnPhjdu5S+umPLVo8dXPMo8
N1zUyiUMj1yVY2yqmpKW04CnfzKoBRGHsytGLcFV56eIBFMOFXyH3NuhLNSe
Kh6zkElze6Id8tvoIrVuOATSaV60xmar1Zm1PDD9DZg+jU70gHUlRZ/0uYcO
tzg8EJRDqqURCcfnBvqXfsbvMRo3bAfsCIBq9qMA9l0QnZ+2QAvAnoaWn6gR
RC6N8WUYKtMEWKdjAyydeOxO/6j5r3bNdKOl3AAV81ErDEH9bDP10DuOaaA6
gYuu54DPnKVhaHuWSQsk+oQvWvD8g9T60IybdC2m79g6I4xmhNttbq2VAvpz
JUkgPgKbiimUl1DjEDhs0ACkbWJMbIZvXINLqFm/bgh0tjIY6Az7kD9wol/K
2kWIsIfXKxleWCj7zpyAVSlaWgU6BFnuc0auDTAET1Q8Iug8wLJm6mRTjEjP
0r/b35BXWYEyXTdSUkhumo6v/1DJRQnaYTTDTZdzObcih8wRrbW8FcTksr48
YKJGCRgWD7mxkhBlkozENBWN5W5k+YztSgoOwbK8nmhBP20gjXsCWOlUKHjx
CP0T21AXJsbbiz8jFxJAyfnHUIuPuoQRObGzRN1d686URG/mq+7ru/l2tV7O
VK3nM/kInunEwmVNRlaHUSqTweX09Fbbh/DmW5XlJxGlz/kZXKW8wi5YCbYo
v/0BWCFSYZPEjwtrQiz9K6ybquS2kctG/X5l/8vTkn2xo0X/Lhv7fO3/8r5w
FNReNKx8LGQe2OAXhDkkS8MLOYQ4o1DXh5DyM/1zUHLpOfbnkRo8uIXAb670
dcC05AwyIokmpV/WtstmRnOZA4JNzOYDeI5nQRH5zS3w5AKZeadmg7kP6toB
PZIg1QIzkTaRCR1yJbnBRTNTUE6G2zuxLzxzwtSBSPBswE1u84VyIPe/0jnN
x3fAO9TV2VyG8iUdxtBkVq1TeitY3NW5tWp19FkNFjnbQ+0WKXminq6Yos3u
AazINHDXo7mlEUIlM9TEFwgBHm4nIydFTM8qziu5/QAn3J0CWwM9jVn4vrzN
hc9Ib1S8WY4uSgHMwkk8sDyvJ5UgK18ODWiB79Reog6mo6n5WinZ6jOWCYUG
AvY+sBEAjFxOcBD9n4cNxTieN1nc3HPeL/NxbGM7AycKIFxBifDk3Fa8dRRd
3e3nblYnMsTAZSwmatYIGPpqBVe6cAJ14elnKcdDMYwmXWQZ2MoqFGkRWkLL
8G54xQoi2CygxReHMvAaEls2RQbRIVN0ur5bm9WDzKDG9yQWEtVW286TrYFH
0E4CuNGOL4Wb28ZiQ9ECAFmYdfMBgMPkW90aZZPt2xuCfVVrFIC3RFaAZurU
29+HJaNGDZKdQYHfnu7pjHAHSIN7rT+8unZNp4BkVxz6cu20VnBHxB5JU7S4
bhsecVixQasY+btKAnfmteSD8u4QNpCHKD/PSy5tszmmOnUSSFrKeOhU5+Ul
kNjXA0OoqFQI+v42vxTiQkUXwU7BbOfyliAenxWH0XT8FC7nQ1cpCuOhhPqj
cHGwNJcV9WQ20WZJZN9rRXDi32eX6iC5pDqomezxAqEjE7qU/hK9A74jtVIp
ODpCUSwV2o1GTcGczu6N2an0AWmtmvrv8XFAVAUt8ngg0uIHQYlv2gXopwcU
i8yH+dHkHTjuFj3bMF9FKZTyI+KQcBS70Mzv15OtUR7lxuv0T5JkggIHuoE6
PMLmC+PgbKtiQSjKpxh0DjjzrIXV47pAzly60jiSMMr1P+PNcxipaV2BgEmg
EEejOYorD8nw2xBwR6d1HCWOvu3dv2AfgQZyCj5jpTfFN7XvCmA2G5P6vvXa
Gtaxei+meID5/gn3d0Dw2UTdXaGbU8cUcqg+3xQ7tUAojJ8V20gRVP4k6MPX
lZvUKoiZUjoWQxM+zN0WX1JCvIHoeVxAaKtJazNaJUaDpZ/oGwt7869y93l7
4RImkCd+DNaqTqz6T108m58eEWLXqkNyxvAVWc1w9TJzFYQKrDmnri1+Yodf
G01El0YcIs8LdJfeKfK5vEK5C6WPhOy/hEgVy7yPQFx5k1G/JRABXYQ4LtX9
/RYldZ0N8qRa2FlxE0D0gmUMh1/CwyggoQde3FczsY5x4gS3hC51oUvQniym
RyniQOKtwAv4P6u8JqCEzQUkYaDH5hAcZLpXrP4Onr/L2WbRhfoXPO9lC0d1
/Vga/u3DFvi6qvuPE9B0oJrtJvHCyPuoySu5XA7EGtNQPZcDCbWq8iNtyVxp
KnCQZXstX9WMsxFAo1y1N0Hguj5UDI20GMPWwrzpu7faie0/CUKk1qecEAOk
zhAE9G/t78i6OnEFAwCWh0dfp/0Hexteo6Fz7dnHz5pQe4BtEwg71wOct6Nm
xDCqrnW+MkFA57askVdT1uWSJbspg34ou4f6RSNnaHTuRlp1tFboqkd74kEM
pxoFsByM7aPJ0ehi4If8EbhCHrwMhsaWTvMZ6QSsxl4VDWRRnYlkJm56gk2A
uKHaqMqrkuvt0b2AUaDc3MKkhDapqw2f3+hwVwdPB/RZlQWBO0jGFQ/Dea9V
v2Pnia0WkoBt/Yo4BZYYrgyXC9CNCbFWzasqkp7djMA2dbNx/jCkCAEJQ0mU
iGhKr1c9c03oe9sJYc1jh7m6jk5SpTgiPpQapy1syOH0IFbtnJytSDxicZzj
fJN0OMyFSJ74ajUXqyhol7zRGnb5rLjeDfIQbJYn+xiDuIWwl389gGV2qkmo
+s46FOq84GyTxpxhwYfzarUKUZyuL9JQ1EybfAznlPmklmTSDnoAVKgGadGl
yBZB/FyFTRuXSc9NJtYAHeYjAba4VfEp0Qn4+1/kFOxYVIqtUzk69nunWM4z
CjMdYbPgXgoKf36XkYeB/NMNXTjjNNp2JagnZqj5si2O7za2K9V7x7enMva4
Na718QMme1ySjXAfswfOBg9bm58etEVA49GlhY3HsQ7WH2hcEnHHKtJv8Y4E
JVlL9FX1qZ2SS6td+OaCZKD8w6w5buTBzFUCDP1kNdVp5Cs8bgi1bEkbkbm7
ZPal/u/bhgsYmvluZvII8gLRA6fzUOrS+ZBJObNpSoBIeP/NkOgCtm8nrrXB
nURsK8mekg+Uf7vGHFjOGyFY1Be6/4JWrVSkuNZ5SaVtMjBCzvBRylQj85xG
RhF1/8ic+IJpI/xJPNBj/YaaV72Brt9lvnf09AJBPeV+weBlr7vAWItvy9Ue
oSeS/cjKehpUnd/jUjOryLdMTvyDVqnX98OQ3qoAw4AeXwz+dmbwYqtfiULH
+QRHOXV6NxwXWvg//zwGOQrdZp4MdfyiNcY=

`pragma protect end_protected
