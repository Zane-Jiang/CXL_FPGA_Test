`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
PlqhHZ+EyBgXY2QgPzS3P/bEFbhSCNsRw7uGNm4c1SkeNItsX2KCHfmdNqU1S5+3
7X2QLA9y0HzGOg6y30wlKOXaUTZ2+BWp8eOJ5Oq8Yra7+i8dLfl9WWguJh2Z8NQp
w5nPvwNlJl0rluVgqPu8n2aAINU3og0ERVwET32duVg=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 7488), data_block
Sayhj3VWvlNYvnrraJjBdq2EdFxbFKloQBo7rpHgQO4chjCzY/mP8GGv5NMLwJ6x
nc4iNQ5IEBY86RsuarwgLNJKJ7gNzAChA+ZlRUKhEM+0gcweoTG4dt0RQw3EX3i5
k+K2khPoKpWqdax5iNZ/qS2SJ1XFCfD8NvIiJX5sUdu8NoNmJQrUH6Mpj5mcCpw4
0wvcdFjq0Wrn86O1Efwn1DHI1r83J/71h0TCokcMD2+3jiZR9tCql/wbdu4Oz6+t
vujBfLAgyDH/77jUiVSNwumvbi8Lo+sowSMy2xYKvFjHDQxLQIEN6IKPxFlmq1Jk
ro3iHcL2QGSYpWaDDAkVOW7INU/Fya8mhHtLP6xoMiejXNqL01QZgrKOrE8YgBdt
WKCMfNlOsvwkSp8fXrwHF9g2GtzwREgMI7Pp3rtTdJcTB0BQ01oviBgki3xJ6r3G
4HC2xXD2yfoXLXqfyqheld6PlKq9U46pMZHB7lhwLsTI3HqdD5wK9Bq942avP3TN
MBJhwvx0YkuD9fIuja7XBnBZjlinMN50vRKiUzCIv+DG2avt8yneQgbe/YOTDCTq
PJXjCQl1NpHU9BbsA+ljjd5ixEe5x0Pki+eeoCh6/P0rzTfIKQ6UbBNvasOwXJXx
txuNeJCh5d/is2di7uel7sqpR/UL/93eNmgCH/0Gd91z3lVm+rRsUGRbXMM6Ae6D
FS9ajA/wKD+5orkcTqN6cstmVRp4fNVXmNGMc5kZZV/YaWLn0lgZL5uns5H/EeX1
su80QYRRku8HsTwPMUDeYOCeSNKtijyz0aHH4TRxjAiiZy8ZZ6+aNePgzmMkfkAt
NyUoU1+rq1frzwlY/Cvpyx+Za3AC75tYq9wMuSnNhSYWzFtLRoPkr9hN44tJi5JA
1AEBWeiN8fDhckvaW0LSou+a49C4PnSIana/fVnWMp/hmQFs29fYwYmYLiOrpX1W
8yBD9zvB6vep+ZZZTakbCc8hGfOr1h+U5qcdTzcAeuaMY8MWgsah4eI3nzGVZslq
dSS2w/CTDBBttKWfr8P6rq6FsmVlkRVL9gkvX0W5nswZEXGBO2mFFW2yowZtu2VK
pjqdBan9QnIFhqNQHPxKTWT8evilT1uk9fT8+ob22JmzNpNPv+XruBancAfApmm/
9S3DW3fkNbFTiG3iUY5ywelWNjniPJBMOEXDnO8AwiZd8twAM3Cz8qC75aFjayMM
FQkkkl8+Kj1Q1PuYS3sevDihyTxgfeWyPHlJQFw7TNT223W6DPlYGizfnMQFxHzc
4OWaEPvGNYicoZ6GfO8vm0i8uNmnvlheTx0PdRHn5MlwJSE4KZsgTJoOBMJK07uL
/KhRJEgS4ZdLf+LsKCIHLCPJNrs3LUM0gxtWUkte2p9S+Slzjovq4WfykdeFTy6P
2b3xwbaJ6z7GVEkNDvKXl9NM72tfLDaSQ93pkw8gXNTL2Ju7GpUDhvEPzhjGnJdh
qrYs01+nxW6eKujng98UN5hCUrWEzpv7o7lDGnWFzxxjpEHmejkq5AGCy0xUymBV
3z2sO2kG3U72ZIev/TqjgWpimknF+o6J1PBNTYjX0YIwmKKIHRoMlLW5l3OzqpFt
cKI+J57Rc0dfrU5Wn8+J8F/5mwMv0gPyiLsIm0Vp6Hm9Vm1e/F1MjKxxRf4HKuCu
mOSE8QSSf87Tyyadzx8gj6+He9YNVAeQmnhnRLJf8b4MFmfROQE9V3we4LfK5yWk
c5cX1i9joJK3B12twMkv1fghlAJb3upN8jCYZTNuuEGToKNlbSNI8Ft4s2D2nGIY
wY4q0wBAMUHvtRLPk4PN0MKCCjdZtj99ejnVx79SoK+g64vlfxNlscBbGS9ohSOU
oCpyP0bkx4yh7xH7qa4eJXFtgbmHQhqp/FLchseXriQiXOSxfR+PQ+101CacKuae
VxfwNtfzcql19sPh0IFoGTz73QnOQRJzJ241Ua9OwoT3nK09ZJCR4RyVDI2tKbBb
a1dg6B/ZAVsQvv0/NKuL8b8oqGmC38cxDF71tg0VI0BNYxAVgHz5ZUQiSk1JbDWL
yaBtRFvVLehiycXDx14Tjy1ziZ2y2sfblj0Uf+iwddraEouH8RO1yZn2dvmXT0tc
fD9fQwaxWcZxjZC6/0W6/KeHHBKYYnUFHxothmal4Qw33ho3HtMbNaZF2TDm/RWu
82DpT1sNR1/eiYW9Xl6ik89UnGZcreOL6+wcvQOwWGqORiRYPIUw3xDmHDNtrcBW
+5g/AVUJdWkxIlvLRFQ/C8MsVs70IAhfTP0TZkgbPq9EzrrFA1L68U1Nm6raOwTO
CNz0X+wojkipn0ixoD/gJGZ1YrZMg9jLhqnAMIdBYJUMm6NGOTZj+rcDxQCLUqEQ
mYd6oGrfmb+BmMw8fIM56ntrMXwGh6uQU6si1RG+KrjAWry6EUrk9nnuB/qa9qMZ
pFJGCF7whA4gmA+DlQhZApGncyeFcQJPcWYIq5tDs0kYLvkDmQc112P1LVkuTQlJ
NHnPt3RTqy3zGWhvdYJ9HRRQ0B4nuaA0L4bsscoWCPjISJPzqK6DIykrmk295wFE
6DwpBcsWPiHOqYZ5cVLZEwgnpOt6r/dlzyMF56cxJ4kIA0x1iR9b1RVyFkToHvBX
CFv1SajLcgsUIUtO8Gm1nXLen3w9GukMmGeiCn4NXQmwgswoO4q8ncNWpY/0kDYd
4S4uQrN7aCRxMcemK2PLpM30qiMJbgRPWSTUNiTYG4BxYF2DVqcH10ch4IRbDDjy
6w8r0ckejyAt/Gv98sU0qxZ1tnIjdgrDN71zW3ZLYa/DePmBcyQO/Q7X4PV9Yhk0
BO3ddyk1GLwEW33KZ+6fLPhxz/UR2vYnRlEfn8CGS48qFvy8lth3TpWzBrCTV1fF
OAtc7N4+ZrXk9HW0Ackr8DsrHpWVxNCXU6i1FvXO24/gz/wyIcXaRoCMf37g1CfQ
WCFFj13J3P/y6RXN/QEvzga19HBai5h4kPSv+W3f8NXo05KRvOU3RMXBaXaG9h7T
WOfXRVLXsQ191Jdkv7RE7+xMFKoPyHEwlLXUTGTLdG0UfmLU6EOO9WkqThMpnRKh
B46I9Dxw/xlbvZcgBojhCUl0ym6MVBp9N/8cfHhq1DsXaseHuvKWcjFEltYscbQ2
5+Uq7c0c9rK/lcYiVOiqE12XHB+xZzaBUmMUKXAmMps2Wau6Y5QL6qU7l1lcTWrk
RDW/IC30WQunbID3PxU/S2+NurSviNg0pXTwiwCcLK6rYHgpCDKzRcJBgM8SZ+e/
C5Z/T0t98/ozos8FQwyV0+odzSXPZwyO0s2hAAidqkdwuIqHRJjBOiVgEXtzjrWs
syZF1QjuSSNveX1nR66bGflfElqj9eKhlDEhIFkorLpr7fywVslV/FAs9zY0g8S4
70dnIED7ER326tymmQfDLrtujs6/OX9T7XbhKAQyac+5wZdVRRCsyHZFKbAMvlNv
LgjiOcx7B7dbYBeKaw4BGqyaIqFi+zl0suqccjn+LVA47hKBkrOWjiKiOzq/O++w
y8DE+eqYKfCoQb0S2god5TzxmpEXH/UDDxuzNRVFZzkDfSFh3NeAUqkt49F+2KiZ
4CbiJuISI+f6lMdlQv2nwKx0ymzu+S9VTjP1rEcmX+gpyFT5dUelt3M7rOJ0i6ld
JwjG8uVvWLcI/LZ8CsWeDASMsUcWOhyyZD+KjwGqO9wdF+bi7nhCI9Kl7MaW1odl
xpnh6cjLscvvYk/cQZAvcO6nPwNDKQUxFdjunFuuGZvvvBdoWlG3wz2lIrncnip3
fwJki5EV5a8JHL0ctMOCHwttth6TkRkP4evOBwdlex056+EdsCpeQLqq8/y2Ko9+
Ml0Sh2WvFwPa3rAwWgR2v19/ybiXe4YPLsMQOS60ajz9f3Ml494yM3ySzHpM/LBK
4zJYKeOgQB3LAB6rcyf/t267i4XG9W9koR09sTRT5U1ecsXuUSbX5ZolzRArJ0Sz
jGsAO4IggRD9/aiDAO/y3eshSXdFQWQ2jtKlck0LwH3dPks2bv2s/hUkY8eWMM5s
wLpoefhTdZKyCPqFoQNDD17oMkqOORH0xnBpPoTPQjJlNks7PYvkONHMf+mq1NIY
ntKNrJ6QRrnoYqwwNUHHu5up6+MkmNLKPuf3b6eCN9d+KODTaZPoDwSMqG9lbbQT
cLKYHgDGtLquLUkxlMmqtQruVYxAPGiyKcKWiR+8sa+LXtI1V0323xUT20C0O+Qr
H8Fu+xHZryv4Ofq272hRknCsr0iVK8PGO6UuWBkCVGjLOSDo0ulxf+g3BApPwFKq
h+zW/ZkZLHbuB19wuaNkhXu7+IAnQ5ZLvfwhqhwXpjATCi6FUWPE1qtw4SSrjhxZ
MQRBMYMM8KVVQlUnuswWgx7WGv3SrSuYLvs8EbK+mu7CDdhHbRVZ0MPwiGOrJ0SJ
Q42VeYomupJw//DzWm5R+44CVWv2UbJZCUWE1KaDcBED5UOdONcxCPOqVc4143+X
S7dthLIVZ72Dy4mrsGjqtn4bnAWywuOu4bcQE22LfpNG+90F6qw5FKl1sJ9H50hy
/N22eKZd+gDrNH4W4MdT6qr/5z7WmpNtK2NDpQBornuV+iKWBx95bPucSoMg8e6d
Yd30x4VvWC5yQa1xCG4BnrX4+sxxrLC04e+0j2r7VQsK9Vvhgdhig0Tyi0dl7n2t
/Y6hOcuoXBdHDBMXN1Xe3mjTa7blT8WmebSjP/1A3EnrpfsZgcodOKQ2PYLMVVee
w1M7mr9yx0NZWVuVCGIERRPcDBtHzUc0XtaiE7ccHp15txztyTUtM2GEBAFXzrYu
Mrj5dU0D748ru0tWnGPGBoJOai1MG6a41F6y0rRVxKBPKra2eLolHjp0bBNmcNsA
JfS2SpnBrxDNuw4Rz1eWsFV17M4XbHDd2jKeiuzyJTDFjUVeq5ePU3maQjf+dOnE
WEWZAhjPapwyqJrnZPJqxyzynnHBaG/lMok52fejlLkqz2OMaxSgZrNjun4vhNqq
C+hctBUNP7SHHvEaJcDgXqQOEjg24vNtYZrxm4szg5bxvTjd8H0wH9TNwtoaC59J
fggYryesVczmPUJZ82DGpjXaC1taUU7LMJkJeNxokioE35HGsvp8pAMfKTzK8a/J
KgvOhj0f4XiiK+mhURMIHEr6/AZtsc7g7ws7tjSRqIf1AYxrmCi89EuKLv1rPP8o
9hdcvCvvGleevgVfEX4hYBHYUry6spVFrL9BfoNPCx08tpcv2br3iRD6v8IqrnJu
8GVo0L0j0WUX+N4Xqtsf5rij1oranVzOTzmBwroOV/p7sxxtHu1oza5xJdw+iL0q
YjjQiJmKQMdvHQARvndYwN90HtUQvyA17s/Wrv7GC65QyUm49WdEX8kQ81Qi7U35
qDQOTI2kyaDSv1bZqa6qIUYCLoqNdJoBY9SQlam5v9bbfZqQHSqqSLN2LAAd5Q3Z
7Rd5Abj86nChuh+PWNz04PZ0ou207KtGjolAVPcD1oI+1euuyB203hHnGr4HDzgI
NAeZGSFp3GRlQT0NjFKDA0v5gwBd60AATSzeYXUqTVtbr94APdhWpsnULL8kvIru
pVYC/wbb5ERPtTt7jUbLWLjIXkdCP56h1qeqP6kSXbVTxS+fsoxvZfWSsyunILGm
Zct4DKxfkOPsRj+6j9YpbsoWQC0zx5PKb+Izr8cIfvZQHXl3wM9zM30iQeJI45Rw
MfHeJjFkjXNSMFZ72DWfEXGHlpnnuht9ORXgRiDywgbyJxXnHXD5DxK+A9ZbN6bp
7SWxlX0buuXrEN1Sf9RQDkrWDvevSAd4LgtuHkA7Yn8w2k1Q4y2GlLbwAkZUGqzT
H0SRKE0dJ2f7qpPJRN1LGHRFPePOqKK1QgaBWPmy9/T8m5NWYW+6rjT040E19Qud
s7yXsrBeie/bSMGU59oER66v+GSRfQ09KJd4KGZWbpkPRPuTC7dOrL3NPJHhHJ64
FrGzdqQ1uBKagtHw4vfXHAKKQHsnAcCWbAuPv4rYjhLdpiBYhHBBVhdrhXd6E+XI
GzG3OkFsTl29NWso02BD2B9L8WofB4lMb/FvvakhXJ4rbaQofFZhwKeZdr/bTt0a
+no+zVCttWPLVtvx7txzogVRS1H1OzolT5oOdKx9dzTmZmLGiztGx3CeK5GwEABm
Sgz7W5ZA/vcwMRzj8JgVj8zNeEubB7IlNdb+wlripsYJ/zTF9OA/AyFz7YOiJuxR
nnNFiLkHKxAtpN1idCFrG4pekNI1ZsvQ8yDQvHD1I4JjAfmB/8FFgvxlAJ6GjVcj
eDdz8CgGdDrQx9/oTJM8O5K/al0LWui0tbrlbfJeEPktxzara3/lA8d24bW7Po63
NOB5Ri4QP5rRkqiRDPqhyaR6FRY6b8R0dz7RJ94Wgegqa3b50D7xUgbyFTiGzQtQ
KJcTDTo8xUMWCu4mKWmnr5sqmxwIaGKueQc1c16EKSYb7kJyptuN283IsPBx7xx1
yxQeOfWHY5MQcF8JWUGXUg77sRgmi3gBw4jw0WbJsP5CQI9fPTEluEFGejYGZ3gn
NrZxyiAS1iueSkK7KZ2Na94Z1JSg8l0vyi5rGzf1tDJRaTKs5TThWFHlTKIowRU0
lkFwNqev6B9TNKXkv5zv6Kmg9lFefwH88uG2vQyIQ7YU8z9kF8VFiGR0I505z25b
cN8BA8MR1ANDUgvymDO/EFo/9K50WNvRpQx/RDFwd6XhYkhhq2r9tIEg468kktXc
JBkFILQUCXTUicOAaRA8SRFZyrJdODQxFweRtLDhEZutwBEPekeH9WkceF+Pj2AQ
4Fi0z62i8OndiaG1o60dASEC/L227m/A3Wox0QlkxSYwk7KhPn3KYtLevrKsEDDJ
FJZs0yHTAGJ34499eAPs7XL1DiRsMxa4Zp5GI/SsfPGn3XBlOGeEkQ0R4RYzibW/
DRtDC9ce0jzDgIiI3deYdnsjLTnxoKXpiDIdV/7ji5RV0BB31w42kKmLIxZcV3EG
ZxWloCDRLA9r5uz597SB+pdye0Spokhd6/ZmiHG2dRmxMtkOtVth+z9ghS1BBy7s
oj/TMo1XSpOAmqkJ2waCP47Htl0MRT1Eo+3ttlBTg70XIdrQXAMXtZMeLcH1rhgm
wttF8On4f/jPllXnLuHWviJNXpEV/21jPFmNSsabdR1Ka8GmlAv+iMOWL6krcT54
2vHxQQOY9ypSpD+5U0V6BFgJ3tgWtTQ3Xa7CBmvCywECPP27J2T1SZj73POGsxhV
sDfEa5s8EDX1/cwAawuObJ1XLKm3KiXyW5q9UdEhu1MicOXAfDnCkaSS0NMzN18D
7Oa5kTkayOhTvD2Vz0MR2jHgylD7if5feeJM/f7DsbUL4pQZ0YPtvfTdBWWvHVWs
OGmx5rLQbCGYlcuJic1aaVsvpp7c68/Tk3KKWXfm98PdtA2KICRsP/ORzHWkxyOT
K9PxKeGx/YPG7OkajdwZn8vf3h6mo2TwreSoAZHBZ0QXj+EhkRyH8DmRJlwSyIQ/
PLYsMxlwNuZHkx5GfP+yqVINF1DGL+rTpzAdse+2RhQ+KF89BtktB+DgAwx5ztV5
DvgJlUYiEf9AszzRawEOYJhN+eKvwAQR99D14H4sNeM7HsdVcWyj4dNsGlKchxF2
y17B8upeZiMbpm74JBBlDiwuFWlbfbT7wsOCethe7As5sQHcHn9/Ok8/CB8onyc1
WdKBwCHhryNhKxtvULntFMrcQPmeLSiX1GSA89cFd+HSs9+Pljpo2OCh0pXtm0Ep
ysgMKHR1t4v9QZAhLxklRTeUa5gzUHxbihf6VzwGkDbrO/mMiCy0HtfRZuFSdigL
cWnF6BtO/5iQ2eKP8FVwB5KfSraFgTRcLnD+hkUewWkSrAI0OIqq93xXjmvyJGHP
E7Czc4Coxffmus0Nlvs/W0EoGVq6Nwnem9tbNMOapEeZQb6HGtcvIjHtjAeIzcxB
R/0PWvLm6QcAkOS53YGijAGodW5yaEE3ulfcMkVg50qMKzQqZLkqTx0nUJzEr3ru
U8eixAn7bq1+E/m8Q8B0kHEOlE7aTo2mDaKarO7r33IR9+n4wsitleglsnfShrml
XS1Gl8CuFyj0hJ+/YL3kbpZul7gKQBJb/fRdqT9j1aba/OYaxxBj+3OUeMsBcpZI
Rm5+XxTxF2U1/MiA14bKP9C2qiY/ZOBwhz3C/VgfKlQ8UnShHyyTxWgzppfmsCOr
+1H6RTP9101Oq7KFEnonhKly/DfV3usRCLkr/GC3YbuvE/aNGsI0B57DYg7w4w7Z
Qt3mAggV38hNS9OcIuggKUWu29C2N7mte08ImGrkQK6aVs42EyAwZzklKgB51Y7J
VAyU6iBK3b50xFiyDj/tfLo92jtWh4qJgDzJdJ/mL2P9hyQQSYBBbISoDdrp48vU
gyu099KiAtSRA8u9f5VvU6F55K79UF91SmdBeZn8wC9MAieyKGb0TqyBUBdklt92
nuTkWf+bIp5TdkG1dL/7Gxu7D58NSN8rZOFU2WHurt+norXQZ923CsSoeFGyfr0x
l71IjMB4mUJWiJ5hWMjCBXBff971EWSetJAqfo1C0tzFf+3LjdD0EaIYnZKSWgA9
MQ22hA/KiPjxsspgXu/mqXxjpwEvCs1XpJn77KHSPy9oi4v3z9hX05T8Jxq42nPo
ryZ3r7yZa56cjFF4yhe8F9y/fOB57XuRr0i+3lxsLni4Z85VDD1qASplYpgoHNcl
7YMVHzUHwre4719uI2td9y1YbPadmj+o6xvi2vMKK3wCaMbFiYQaB3DSnb1XGZu6
UEL0guPE//pS4PZMTAyjacviC676xiCPAXMUZ9g566gU1MxSPB/9iGY7rmu9EZ3K
1XV4ubHOrvIRJFtO/JWmcF6hLH2w5BWvoQyBccv/8etG7xHAvcgq2o7X3ucH0VC7
srhcUt9cGCPx9Q44hYONPEv/tN6bIyQiyG0VzOeiZX2uu51jisYO7Mh4V270cwX/
SPXxzMzBxLj4uH9cB8G3HOYGhxhA1SwYJzdrhcI+9GJiU0TxC4Y7r/Gx61DadVjp
nc0cO75AZdGgsVa/5/aNFyLAzAIjDnMbN0gylwm7haiVGyWSR/WvI54z53pIJ7jH
7AL3MeqlOdFTJEogkDqAj0ks2BMnQGPfqO88wDAd6jgzCHjC2vI5OcrMotSJz3Wa
GhYmaQEyF0d0R6YE1u/1L6FO9J57rGHBoPY+zGqpGjfx6SQU5yaYSGP+WOrWEpej
T2qKITKuwRsf2kdpb37qYpfiF/ED8Yk3NANhI65//ZMb00NV+Ikul2e/c0/mxQA6
aIjU//7jUwpwN+bXocU0/kU4mGJ4pfEGslImhvRNIesYvsFpiwxh9y6D625EtEuL
q+Bgok7YjxkJMPl70VwxJr/7LPJgRiCnEIQpdmi+0u1u9RFVdVN10kVSRufshH4P
jHEE5i5GxC1yKFW/5nchO8agT2NgbQ5uxb2G+ItE7nSuNk4GdFJTmgeih/5HSU0k
Z7xWybVmKY+X4QCaeeCVk1umFin/FnWOzuQ9vDF2bR5T//4UGc8eUrf0s5flwV+J
eosXENVR7BEirZoMHxrBMZktMRgHcFwu+st+vwo+l7zeidbkTBEk8nNnlLOqHMz6
V+eogzq9lYleW4RAXP54h7HDbr7UZZMe/LDVK+4zAf+dWP9fmrZXb4ZGo2hST/dX
Qr7TrC37t0Eh9cjvX4dJBE8MYcDEBuNl4oUjpXFeA5QH1fLag6zMxklDFMURN3CN
6WmjdDJgBTaU/U95pJgiSkOxGE2cpnWCxTbwL32EbZwPQFMD3aDOKOGPSHwIR1+2
tj9fe/asi4TCiFV/jF79wKIMZFKGjWXXfDTtURNXON1Q7uyIGFBiseL0ViggE7Cy
IIP3bZ0rmOYTSvwj/FXP2HwH0HYCSmFmVplzjAt4Ns5xCwTPEy8Mb7sjcvYNPx5Y
2L49tAE+UBAD4BvcnQdQBz2sqN3Q1Do27YeyS9jbyXFJQg1SoNKVamfwySVTnRXW
`pragma protect end_protected
