// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
htLmwdP1jsax+tiX5kh3GEBotU7PoYbBARqIQihX51Skcjf3yj24IkSi9dO10dQM
b9IfdB7A2cujrcNR4ToUcF5R2WkpWbHKiOnfONS4Qb3MWaYF2msBeBJqyeQgK+eM
iwSWzBO9r4Veb4J9eK1exnMFr7ldiMDL7YSPDdz2u9Y=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
V87oLI84gofAN8Pyl+R+KIPVrSSMvZOn8Y+k+1azbiIl369daAkiV920r+afO/4Y
GlKh9LfYHljrxcZIBeVpBshHRH8G4yDp39tXqGepNYWqcJv5jXvXAGC8c/Yg1Tfb
mSF/rJpGogn/tHXrSX7ET61wx3Glo3vN489pRZ52prxq250QPDW5sOtWCt+LUbiI
nuzoUgL1kdUmcoeBmjspgT2SHTi5HcIH2kkZVxXM1d6KVieHAKxD3SArqurWnvkc
AjixOs1hlK7bDtiXKTitZMRzHgIwzpOOt/bsF0oD7mEvMtw9kxBc+wmWq4YvbA58
RCKJ9FRsZ/FZQzButgZsUu07YkaJB4PxJFDsr/Z7jURuQxJGvidRoWVAa3m9U+9t
P5hAgpPt/3FMKRVLVts1bBG1jdgQuGo5ClxeEhd9sbmE304TfFAx/0A2oJ93dMTT
EvjawuWX+Ha4cfiG6AckrQy1eOJXYVCuzsWst+4fMqVDS7j8oVswYmxZJPsSEqMl
XF610Uvofkv0GDYGdQH2lDA/trWIDmml5Vse8NfnwR7VISFll0BR2RsBMI8pW6WT
t5OpPMTOs4dW++dMlEo+h9txF7NLoJ9NRnmvInsvRm3fxF2F2qgIZGBjtIQu7uj6
iUd8HJelkH34wNYKeHbAIeuMFevwtqgDO6pLZ0iYbu1wDZvmKlxvQB2A0wfQ8rjZ
ktP1NiiyH3Y5BzbBCpHRJ4Z20tJDXQ7bat7PzfauvNgEz4HDR+IILoC9nT0FhKvZ
a7GIYPhlEjNsJ/4f7bFoy7yTd8pJZAsl1A/SQVbj6/lfFYDcqN0fTrxno8LE526p
700nEWbsd1Q//6NNiKW2ifnGHJMu5E6WgIH04XUT2aLtIg4wA3lwojEF3qBDz78k
ItftYiinrkIRMw+Rb9iTCOAYEIpF9eNSpbFeDj3AMW1A1LUPmyIyNuYd96Tdu328
0MLowJ1OiL8xwbjGkWEPaeuGaIHu2DJsABXlxZRSHF/K3BCbsJ7qHZhXKJmq1HZV
BeMRzFhO0zwv2PysUJa8Y3Hmn5idpOzhsETgP5WibHx5Yj1fIppXUz1gr1qxzEeM
fuDHfagb/BvRGVIVxKUSTuYS/eikUoKgcUwGxgsgrLBAxFTFz1mUGurgKH5sgUKv
lhckPyGM5CNufNDaygnDgxJsqznr488O5DXnYOICFSk/2qj0sj3EBACpw/j9LkSX
ZtNWEMS+QyVrqEt76tY5w3iqaL2Hi3Wb04UsIIgIxoRBpIYUYiLxcq6EkVaUPtRU
ICGeJk1TubRBEXssHW92vFuk/dx7/qPAR2L/kvsz9xXIbCJan4tT+iMrEPdPX4kR
qsfxyxYuXGpDmAG3g23N53NJMEnfbvK/8SoD3dw0Ua/7CN4Zu1oNfcNgjmFjevj7
6L3zSZZBpcIfSq/pijFZq+XBTUJo5lWmR4xQYKbFwfMINAZwzrfNoMC9HbzIOU94
wENsxPxFR33RQQ19Nayu5QnnT/fFcTZhgWZdQ4BXEr4SJ+nVxafQiX9VMBfuy9zm
jf8Rh1jLVIN+frTsLgysBX7sHVJWDfNyU1ra/hfueOMLvxRjRt32+5002G+9CrP4
4ccwlJVCC5htJP+mvY0yBY0gYB347Sg/vNvC/vz59G2acE2qmuPbTtoORcukbx//
vn59zSbcf03YH6mzYLwxs6dRbxyPoLNQHKGTyR2NVzomLbXr5gazlDOW5LCKUznk
YRoNJeDUZdmvJGBRZGBD5DwF/fx5uQTJLFbku+YO2BeMRMzXcZf3NZ9LxEtCtfZX
tBnS0EV4kOOq8FS/6maZhLly1c8WKX/Qd01daRuq+Wqj2CwbNaPL2Q4RR/fXJXkn
pmfW4vit3VEYT8hCmHupwqwbMGYNSeX+SW2WEGowpJxRZnvpKKndCJbEgkL6t8Nc
/zCCVYHcLtjZCygzMVQrBgocqMfIvgiZDoqdpRRmZz1uAZhXWw1PmGihGblehFRI
p78GFzrm4kBrCsbfz0RaHT8CacnrSc1iV7uIQE0V16m5rhUsxeoUNuT7M2flHZ0p
Iiz4ozn3OHLHPXAYk7HqPbdXWf4/dXzHYNTvvagzlO6G0oxQiERRBoFNHrM9RRe0
dyIegjt0nppefKpK9W9TbVKGaKjMVniJUkvGQrMmXJ5NzdRNt2dE6pJj2X9DLxML
HnYo5KPCnUrnix+ja4fmcKtmJRVOAIp0eLve3h/MQphIEKNJdvcntAsCJhEUBN8H
GdhcBHBVD58WwWBe4WrhF8J6fgxSJlS+l/mrsxZB+2vHmhg3fy2sci0hAQAJtA+f
Jv3DTREQN6I3nnVmO3+593/ar67muARU39uvkhDPfPDKJM9Y4pSWux3OGwmJ6EW7
0MDjb1+jAQbwQjfc5C7ohakDmb2ttpSfYNaLqqZzDrKVcr1pHHleRvXFd9rWUh6P
tTV/dnu4d17SD1MmNzmaXFX0TfQYLOsgY0dqmS+amYTqBeCxjoBMLCAPe4g80iOL
LOMTPRd59VPpvzHg8kpDYf2MC9LedpuQ1cPdDYk4SruQgx/vvhLFCfAC8YGFWkgF
orbSTGZ7VxXWSq8X0Lc7s1NSJexLFlFkIlaw4aOMQzUyn2DjIQvxccqjJKSKF9e0
Ub8FP9zA18mJjdibnGgcR5QayLYk74JO0DoQO5iY3ws+R2CgpYemjoNArJD7s7/y
kkFCSLn6klP3Dzk2Fi4fMD7MlV3JdXlhSEC3EnPXPJDcYwhGHNLUXGOZqwZXkwJt
tJhqwWmxZjJV+N72vHVSMHvd8PLl6l1aL64IgOqYD+PMhA3+fiQeqrE1zvC9be+o
gQMe/mWHH8tK9zKbeiuqXhGH5OfPnn3NkPAau+wmkUEVDTDrua4ScSjTI9ztxo0I
89cohfgB7D1CuZksxO8NOZXpoyXyYQxRGOWcme000g7x7ZIP09Kmqi90ppRE2L5Q
pmVKkCi4BV4SlWjxfx2N1gZkkRjBNbfpQAp+sT3ffgQdyCBltouhWtBaK6AazJeb
g2k5q6Mmi+Uv7P8WcNheBe1FI2ji1FNly8H8nf0ZGkTO1TWnVm4AZALY0xVS7eF1
NJyH7nsJQJ/htgoAhk8aBDdFZR+HkoN1ScjKNe8f53iYb+9MTpYI0Ed1I8+42I5V
+3bX5XezvSRh2f3VQqMo7RyQrI2e/CNhEDySkhdZw2URuSQzyfmyPmQCJL1+a/42
PndKynyBIyZ+zK6h7xh+qhgd1r82gLk/Bg+gfHN+KKonZ+bncMhBPsjcNoLtfrRi
W5+Nsiuuqf9dME5y7ehv+oVkYZMda+LufMqocUzxinvBAz0nXkEI0aZ3CNS+hrf8
6srNx7AdCl+oB6o2/DreQxJX0IbUrNzUrtXktHiVzcs3sa+Wf4q+bfKEljjy4U8B
x/PrQZimxTGcYFmtb49ZdL74lMT+cxqFelIZl3I/zNhYadDBJY2vFbzv1ibNLO5J
SpeX/rAHUPfrIIhPXH4b/6TAOFXw3NrrqK1mERdnz9pYkbhORibZ+78166Za21f8
3Iyvb/rH1zLsQmjmd0/L9TmxMow0nJzOm5UJrDmmxY2DRex7dGc+XRfcQR2jQgpP
79RRWJFeGoQkuos+1bB9OELnK3jV9bU1yghHwPjPOb2XVDvoMUjt3nD6MCL1awtZ
Izk2+zA0IWtJCzL9QcVeoz4bjXm2yANvzhk94sKIAp9bqWE63TZM778zMWKIQZpI
Ix926Acb89NraPC4uvdotR7dTPakAvIQXkeBZtuomaEHLKx4eBYrauh0P1pni0Za
TrN2lsxW8RJ5EtaK8u2+o5fzx09IeuFRMedLlBugr873dxEFrXb2Di6dKhNTAoef
eX4uRKBJD20Mn/FWThAhE12yi8bpOHYS52CafnDEXTEZCI4DHAL2LFzrn9i+0lok
/cBidATeip1Y2cf24SwO9F5xkZMqqKIje53FVk7plHvBKgRp4sGznruDjwa+GN6W
qdBBMRnWuv8Q3jrwwRkpan2BXDtUvRhOgs4xwoBpffEyf9sCZeBk2ojiTvLI86a8
j1rCIIK3kZmzRxqtko8vclYWzYeelMg/AS9Y1Ru7gqTj0HFWHGRXfRz5OECaIbnr
3Vwvt448bmaRl8a9gzlSScAaz3NGktDqbs5Br5Bt6zSGBtaMQAkq/ypxHjn0trjz
7L5CnIHhPrRM3fRuWWetn4tJ+fZKbjYFTsuzEIdacfNXfem6M66Gq3IfOVgWdDSI
nk/jtInn8V5opI7FMMo21ZYdjhJ7VuaT+Wp296sNu+ZNv8M0JuPhXheqai0oZGKO
2Gatou2uHFxBEO3/Lh6red5MxTmzyd+1tGIwwvZ96gcG8OljRrmtcNrJ7fqBG2Lg
79fONgzKyYQP81LUMWUSwDl8qANVSMecNgjvUAhZt90Rlldde4xY10JPgFHXMuzJ
UNkYCimjBQytttlwxD49cXAsVjadei67S87focgyeSFKCCLGLX0WxjP9lpKK2lYD
AO5oLdRQry1onrzJgj2ba4EB0g/5FAbXAWaQSd1MGEmth+mgaZsw5ixqgd4alWzw
pDyKuAAqt5vEIYMRewjPJtklStg3q27gSXGc5q12MaQxV5/mlm/5WnY/QZNUJHKe
zd1Lb5jN52NbCwP8t6NOgxx407A0RsZd5v9LpRq/BhwntGen5yjem07K+5vKczKK
usbBDolrwmLjaXkT1JC8qgKl+QyyL33dV95JsjmhWmeH7NvaqwwiVvgEcXzRByDx
Y49emrV6GhnjOr0ZvNZPnAGsL17MXyXXRatEcQoVcMQaOc6UOdKb2rOZBC/wZy7U
MDauzN5eO0wVFj5vsxqtEH+r6QC8ACgbpjeam4xNmHOjB6zOTcVSJZn+z+sBgT+p
MMc1HSW0VIiimiGfRHKTX7tM5flp2vxH3m8jFp039OciEpUhZHj+n0IaZ4xkuDy3
yM3bUaYeh22pzzvjRevQSs0LEvNK6Ch9O9CXDrhb7uZGmGyXwzEM4JQcRdUV8muL
CZQaB82SP6l5P8aB0az9semq5M/6owT7B/QIv/7TKOoNABgEsFXnOBGUjcY4ObIn
nPl7zmq519k4XT7wZAi/+/td0FDcmICaeuGhiLhzStw0dA8nJ1XZJ8UNRGEzLxii
jjr1iUhyTKB3S5RuzNjEVdxntkiCSbygHyCJGXN4YAF5akjGLi5P3XOhdoJsvdki
nGCczUbzcrJ+RBXt0gndf/3ShM68vg4FPa8wnpPe5A091+qQNrvSkKw25XxuoiZk
4Ix+r/iXERj3iI866L7fI2+wSuPw6RkHpoJ+nnVs9E6qKh8Ij4EKTGvQ3f9+igOD
pe/2XQ3Xz9uHnZn6E67CPAnh31oqHo7E0ZGXG4WsHDOOaFHFR5cBft4hO+IEQOPb
cw9k2qmxO0yim9j1hcRtQPX3f7J+swYrnSTS9UkhJ/5B66amP8HP6ExpW3UWGKEJ
J/83/iPnLtmFda5KYGYM1UnGKIw2535SCWYn/Jbt5ck8nJhGlM8tDx6WHrvY0x1V
QIoskyLboo+Z5oBx/2jKCj33uBENUfT+tOjVE6THHijqBagTIPl1Yp+p0OUnR+hi
PQB6GEhsDjtT+JM5HP3ePZiLgEaVKmmIhftvvpWoHihgKVpUwXfu0hxEl3ifJLZQ
3sye8niKIm0LFSfdkQX4Myqap0dlCRxsjCzx99Qs1NIpmU2DrcQmY1eD/eR0Q1SI
KczFCVXqQb5xKn2bD2+enALo3Bk4wyxwDVqkDdQpOGAz4tYDWvENHaT3LvUusT6M
Aq3jMTVpAQ8ibA+CfusuB0GoKp4fIJLBOZXne9os+5wBMtqYEOSrex6yCD18t2rn
iDJQSZjnz51ZIlvHUq6KSOB2LtjlQHo+q2wXdsnFYgBbKqANL8qGFcbYQqQNg+SS
Cxdc1fs6ZFiTm2Rgyht3/1Bbuk9UJ3hKxDAnM6h9JUdYjwBpfOwmuGx56ry22BAj
ZeiuOi9W/826aRkdUtn/u5IxDbcpCyywBc0fwuqQXX/+2HhPlZpBqeNZSwSEPAIz
0kSDxSGehAs4BiAnCf2Q2PaEjEwV9j9uk07gbCcSS7M8fIfVGLo+q03uqVhdR9l/
hMiZpeLaqh2ngCihRPQbjHesx7G/rfQaqBcMIEHODadpkKRtYw7M592KmnNL+hKC
C1HNdnSI0EfQ0bPeT837vuHRJg/cZuBP99OyNSP5aVAB6HC3JcCRyKVlSDQ38xxG
yljf1dPSY944AnhUPiM8EUY8ohfGQvvjCJ/U5G2gRxV6LHDUC7TCnnZuWTAvWrgU
5S7ANuavrKSdwWPRJqGTxVYbVkl+VBu7iCQfrdYkOiV3qh7bN/osn9AU5SinCOWK
GhjgkdeLuivqou8/cMPMEDJBYNEqqUBkZ7BUQM8UsrbOUlJ/3pNslIWguCR7HAaw
CUkHPoqGUBaHgVNVS7rtt6Fyk5jID/ridE0bdLDa9RCPoTXwlZoJTug+2eMa3qkz
8/exDWREJPhzBp6RQt9NP8OyRRNiWRSd/XTCfUq91TSSrJ8Xr1p0maxVOIGqKZvw
u/u9wVTEArKKpwq1N0ICfXSEFKfxbUoN4Z9skmkD0Vh5Sva2C0xFhdt9t5iwLjj7
vSFpU+5s6CGjpo4KCJLWcJzl+001w8fbph59QkDJgF0RM86pfRLELtu16KofLraf
sFfiY7YkpLePLYRyJ3dV9KGxSGdKFh9O0fOYhyPbgyNTkj9/yOLGV2E4RM1xGcoi
Py0l98fViLlv/eTg0AuH1vgtBXoyqvpZMjYW2g0L3NkQ9z8GH/A24/iN3RSEeVPF
mm4pptnXSX8RPzLeVVj5hvRDwDAeck/iM6gf/bpVTWIeYn/oHbv8n0fJ3eTEOUp7
YP2xec2C2uPyPsAecLfMqpFh1AuHyst6kmlke2JNP8mOmAJA8vKGL6vrHse6IvcM
RfOVGCT75gjhjQS5RyZdL4h6RvYCv4SJYM6GtKHJHgnqMA3tyqtSciJHPLh5B7AH
Kh+QK8XEkFWkvfBckIWUqTXkBWNKZNlqmhCo6StcYHaoJHBIjz9y2Ymx2T5ma8vP
BitTyNrFOY6EUyKGiH39EaAJYQ2YMSYCUwrphvmOgBR/dPcD315u8idYT9guN4AZ
Fak0FykU5AECmlWFgokKnZJ+e+sfLI9TILksavfvsFOweeB5w1jcmm7va8NreELt
Vvi/I+EAwwxQQCXVcM0I5ViDLXSQo61j2p2qdORNMwkWS+5gD7Sar2wPXsVl0OZC
JrKt6QVOgdj/pLrFv1DW3bbILQl63/pkYjBuJqy9SG8dTp8M4dDQ5eYmzLYBoMYJ
0+FPTj3Q5hoyYmtx8TcC06wEokaaWdhtRJGXLGPATlbg3Mz3Hs8sBNxbLDLuQQkd
UANKHZrGt3UNCD5Iq/2wShDJ2I07ZsQXPM+CQ8Quz+jCbMhC9Tv38RwWGo2Z3wOk
JDbKvyH4UR0qaVapiwxpAFHHDzB02dMNi3SXjhPoOo2rUlLYwFOnSvmP+h8f0TsH
TEiU3bDJ+yk0EfJB6DxpeOO152BgbYpqU1I2mW4jTAc5/H19WFyOI7TVGtRqWQwZ
eWGRF8CcU/zoTbr0hV75RuuCPnfx7FEzyFHSoPnCUMXeUNSKU1IeiFrerkFthCJ8
ovk5NxIHDFEqAJ0aVcqgs9V+vIv+8yOstvBrYLIkFKr8amkMQUROd47vx+xJWe3e
c4KApne9MDOIJZO0OvWzKjmxkTXLJaAeFC/a2xpk+9DPHydTe4OMe+LXNuoynUxU
wPot4GzPF2X2T86GdHnRNWWaMlAhgYLEk6ZriMdn9QSmktTNkirZ4+clAwD7GEHt
Q9wwdjnk5w3jG0+wL6MEjzJVKi9jB6M6BOdMJBwDrmawyelGK+HgybDZuQITRk/s
2OFzrg4N0m7lnBFOLEl/psmrCRcGLOLxUeDx1VnveC9uymcr/Ubp7kAqNYL/1l2M
XnsU01rgjMer48v0HtFw1lQ6Fr3SuYfytht5Tb/f07Hz1/XIG6U/irX5CHfNbK+S
VqouGVM/bvfQQYEpvNguZs27KjEaPZLZdDr/+NBdlHSsl/buFPrsn9tYQzKRUcmA
nXYR5GUfd/gx0CeNVg1QeN5dNo5tJfEQuxfT8b0ppOCfjU8j+OmSr9tUs9tPdPP9
Kdao7cPQ3HlgXHAZxl62q+xZM1Qfg3PF6YNPtn8ZIY40wseo0J0I5lGVNs3RLnPN
zPYtHq2lWg+CXAiBp+EhxZwaj8uXpWcR3wrhGhDv9P379qXTBrmArJvOq03TYKcF
/qEzL3oeZi5Eqyvi2IEzO6zWwbloI8sNh8hB5xGkA1f/UpOFJfW0rVSbS6nmaQBj
mvuGJtRfSKD9PJQV9dY+CEMwMOu9V6vEZgnsnKr+msIIsDuE3kAHmp076fs2wGWg
TF7J9MvZXVy6ib21ZA1h0abrQIycOWptBuOwBlwyE0Tb7l49gnvkEcruZd2Y2mz+
YTKvnnpW2Mkwje/+7j/m1GP0sAH1p/5kxI8NqegrujKxnoQpascdTTK//VM8rEre
Ysth3e3Z5ljRVoYV9ncKfv++EcRmD+zCYJb3H1EuU3ldq+ve3R1L2jzSo8JgFLa4
kAx3M47jPjSbvZsdsJAt95WHU/fKQtU9cwR3vkZK130k6oOHt7UqzvEvCV2Y1+kj
uZX7SqMjM6+STfF/hhML5ehOylzWqLSpEUcpGB56/8dPUMPyVk83vt7nw6lp8tqy
Hm7R6nE+i6IyRgmpEyloL4JHuHWZMwWpD7I15064t62T1SSYarSbKqBJvwj02Hnf
vi5889RKWBwEOeXcjQaSWhYxd5SQABPNMPb8Y5vtqI+5DfEMLwXwbvMtqu7xv7c8
QVHxDkMkhRrC94in3xOMO2thKUDoqBWaPEp7PJjJtCKNU3PDX4MMabxjyZGLLDxT
4iWFd2FMvfXwsdsjkTtXKwhNB6XlP7CEu3+5cVzVg73lD858msGpDK9kG03I6fyy
AXF5UfX1DykapX3UUntR1c+q0rETtHUTyXx9grjXTJCg4O9jZYmrAGIZG/RIxf3L
OAAvDpl3Nll7cfvJ+L56KeDUaCEj0fDo13nYN/zf39Qr2YfDUPYuGfzfqcqStzxu
lme8VdyPJuoU/84ZIPgkhBBc8gT6Szs+Aj2XtalxdAoy8R1orsGyPUTZsXkAFOZc
kk4DxmOjRJB+ruiCcHRXHeHy/vWP86U6b3VCbZ/ZtD0Nq61RIdPAXRIP3gXhUV3H
twHHa7Rh09I5stRyOf9tJZVvRzPL5RAghDrv5m4tKRcS9tHCE7CYZVg1rm5VeuxM
Ye93kqelercYSv65AjQUQ0SszDiulkaEU3OvEtC5y687ccQUnplO/sTQoDtzfePZ
Wn+jCLSyJEh9MMBMhLIN9yCdA/ig5olufGs98jmIx7dI7Es2rDGutubBwyuqE2hX
QmraNzFHPhLjCjKiNmFO2O48F0Xk9vocQcLI5lZyKd6yvNnF1kMUm03YH0KMXmSf
toVTGjjMZSOeCWjxjeBDmRNJ2ubuWmpT+qSX/U9gs3GpA88dNGnLfYzkTqW4LU5Y
mvXt7jutx6tmTKc245Rb9aQXQwf6Lx6ubKLdR1RzJiZO6HJTtfq00ABhrI2XysLl
UWjXd6os6V2kJatK0WI9H5xdX9wIVjTez3yBsKGoTJoEW0fwN7/SOgkRffOQ95PC
+81VeTp6xRJNbD1gC0J8agnXvTAVXD2GlFsH+TjYvTSpaCBYOEKK2JNE/lDL79HC
edcW1hCZxeCno/MAvqzlX96BtONi/e/qQ4wKPdPfSOI2NPLkbDBnkmXoIwL1MOes
2KyQdVLMY//pxzwC7HEd2uEbmWhIKbGAPfer6Cvy2wKCz6xrc105MHSGmhM4xPxW
l/8VVap9ckaLoZqyvCM0kqL/p+C7ZnTzEHvfluik5yrSf5OeFnwyBaq06C36kILr
7iBL8+0pO7WVbq7RWKAlHWo5jBzjAg9pTyPfCzWiDoFvSaqG6kYvRt1HAhdaBz7/
x0faOcaUC+U88/mpEuOAYS53jy44R9AJXGW6OqjfZMBFscSOaDMvU1ZJWakxCScN
mbD4S+DLAqPl/RvYqIIEX2mNSL7ZahT3XQc/PQbb2KSBmsVyN+lPXB5L/2zfN0HW
kPn2DMdspoIpayg5gc7lDIWaC1ZeDViMY9lgqLDeNp3JTl3J7PBCZw0Ter5ePnAb
dHPBs5EMr6MC9356FY9KnVgTLk2j2xaO+Xw6+jgG++NK/uTPlCOx4mnH6msAnBp3
2wZig+IXZauU4ThyTvndtDEBhZIvSHVVY/xNaSpNsftd1ZraYsmgRmf+JM/W4O/C
sDXe+y0UbnTgnhvGq5c4ANNp7bp3leErBZvnQkrh5CYZ1xXj2DR1ymprvrdXIkDJ
lgCLWYaFlEP38tol9+VLyWCLoXmNGp0KjFEokWtfUqlo2cBMSb9HnQi2ctD3kJOA
FgoEZC8+IH7reMp4G6dFzoC9suXinD8CH9zo+1A4cceusoVe4fb90IfnI0aGXsi2
8UuJnEnG9D/HvJX86qE006uaqzJD0gsSw5og8DqGn9zOlIJjZi5sdVHUNZAVqDSe
9z5K6sbaIi/09ToKUzhaJIXPnil7LboUUJHRaPRcy9RqARR7GYCn9dlIF0SX99RC
vWEMfsEcN9mt/o9PEag98DINkmYVOb44F/H0IBPvDRmSA0EPmPpE/DgUEkmWJ1kh
ZarMDnP8SlBQZyL3YbQF4mIuthg+zPfASrhy+OvW+RCyrmY5+WTDih2zISnrHMWw
EcgP2I9fQcadrs4VacNlKXck7h4jfHaFVwVCDGIksdQzHpLXXQ91nYBTSfM3OYG+
rjrB8a1Wzu90kdkvTJlKRki52UfcveOzAnc79hJ6ILiOJD8kg+qvYzL1jqZOVsPv
Sdocvu5GyXp4NlOxdyw9zxA6scf1JbX35aGxi1ynoe79/43vYWrVjttt7C/THEcK
fM4wANpileng9H6Lgrh9RDnqxx1C2qVEzllWnAr5gMNPfq6mtfs1tkJbpmh0zh0q
EZZYhJa7Zn544xeuhfKpysXgoNndlThOC7BYSZMoXlaeNP8HZX3MVFm8GBgWYED5
DYbGAn5q7Pu9pXxNzK+AtEAk0YcQqsV4KHFChrJCySh9jQJQ/T0KSzXrmB4inmnT
tgvPH+0IxOh7QJVzfQ9DV1DWhqiiEMyVg38lqtx9ODp4Yp3ZY4DUIV8SDYCexiHm
EIUk+XKBt4ylgHEx7GQvNR2yUUocbeOoMFyAHzUMp0LC4pB+KZo20hJUmKvwy6oI
/iKrkny19neu+eEod9NlAYcasSg/LOSs2EUaIXO+o+GkEe2n1YtDb8xCTnenVYW9

`pragma protect end_protected
