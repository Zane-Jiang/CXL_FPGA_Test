`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
SXK7yDpEI0f0xgCaSdQc/wEpiT0PWvSKGssJlbMUMkT+WfSps9k1L4h4+cOYroaP
ikZ5PkwpR5cRhhJ1+2s6uI9FaRiwS9npZjTIvFkZzmAuhzpo0idHueMQZwcIdvpQ
N/OoyDNc7ARrOwNrKM8aq1u2ieTwZLGLmYQw3q2/z9s=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10736), data_block
p37BmrPEemKWM01cMGXEcvt5KFN37qK4ezPspcU+sP/Eu8MV5BqHVHDAAk9Ty9Uj
M7KlhvSZali6hC1kAImNfWx+p6+mse17/MOWBw/rfHII6iqVqq/8D9z6Bxpcha0F
PExgVMmPVGPmXwZ1Rt9GH/h3aOfR/0OYZMb0LFx/F+PuX9ySKF6/movJqPTnZ9zY
O/iNhQqa1CvkfLbklqgU19+voBZLbrLASU4fMIZJhnP19NpsBF0Wbj8jScvuPSh9
i6DGHCeNzgFxCDGiOz/6EQnZjeouWkgKV+uIS+YLSoV5tps7N/DyNxLa+Sc/cxKw
RkTQ6TGbuQowiIpsxadeh0Agc6NPbXwRPyDUMf2/BELpYu260U7PxEWOrWphEUtZ
zMwrGO1toCN9jXYQyochaRF9rL20JUwvPBhjm3ua6eTUFcqyWSh0wAxs5xp59yBh
xAPYec7+FveiRbPgqKcP1Z41wDP9hOrSBunaKbMc3/EDla/sKdz/LF/BMm8ubrH/
pnlsCv4PIftD0CrfhbagOGEKuyla90GM1BlwDFNmoHTd5FEAuzU9MPAqO//G5unZ
RZCpENuhkf06QrB+WcYyHExATkOCDsRSkOL/e/hiX6ZKT8p44ZaRCiouMyo8kM1N
YsftdS4xqQFKS5ALCXcjd+MSeMdzFTupRoqJlaq08lXmLxsJxCG8NozAANchc8Aw
6Kgx61hxl9kxezRYD1CGi1YoxhiEa2VEvLhzY27iXe1JZ2Co/HAxwTrd8vXieGhF
w4L/YNUNvkK55fU1z/3QkDLHx71OsaXn/bZxDyItSEDxmiNDLs/J3siR5fUFtnmM
L+9dUjeUKnu5tZB2N6uH88171dN1WunAuZ6WkyPE8gn+O5QaCWKXkrbPFOIuyeKX
BizZwKELODkDoj3Pys2usrwyPT/JgJjHoXKUc0r3ifQxJEgg9kQc3xQg0dc81bAq
Qof2wfiJFlH+IvgiRK8yJ9jMS0gBLMw57WMr19WADQyaWVWhi3deOI0Q+X3pzpF8
TtDYRCJnKn/6aImGvb2NGX4nYUuV+X12kcKWWK0eC/rXqFJ+6S+t9yhnFtIz4dtO
lVr9JN2M9F1TOiyxmuTbjQzXoLK/MLV9fW3qcX2FV6A9MelrvF3kcdpQrvaoZ1Xr
s4ZGTWKQoWwnRuXJT7wEvVo8sB0IT3LT02LLmJG24HQZJgT76pe6LwyoB4nU8VWb
oJqnB2JyCUIiavO3zoCTfOwYa3EXV3Q2CZ2GrqOZJ4wuDCO8q0xn5U7jOHJ0rOGE
CifGoIypZ8BhKYnMsz+IiOJQdDY0VN6feXEt3GzJJmyUM3kuVIz6ykWB7YPt1pAy
LDY3EOAHpDoxk96TlicPefC6LASUF6vxPsyADZq9KV8RTaXD71CF9Uc7ocGEUwG7
y7zBSQnnMm+cn46+u67ihwVf10a7XnqkAP+GvOm5Lw+YDc11xtRZAfaZ8+tTGYp3
XnRRTg9LQUUrOTM8ClbGwzodNG2+GIvpyP45qC66v4sOC85umJUEq4D7WBasFgxQ
HH0W3MbBU0tZQ1cSuzKSz6ZqIDMnQgJ3GuHiLipursjzXEivN7RsUbXfkhhgLJhV
yInDusr7qD4vBPSuN5tC8i7AwO+PMQtDHI1TSGPyqvzOOQnblWUSSCUYczHtCOSC
jynmtxQez66lZZSqs1JEx5Vav0P58sM+CheRURL8iA7JI4WVtS8v2KkTYiX/tp3i
82PHnpdqqULDGyIyiW4qz7oljEgg9es0pYhXtQOMRPtlKBXiHJ5Dodpq6ytPGDuA
VsJWH27sZQTQ78gwmgtAncBhlvGjG38XdFtnH2XIL1rk7nF9IHosJYxesRX0TTzr
MiR/i4BtUf/5MGyMEbJA3idUcWGai5WoCtexcqL0Ij+fFPf8urNgeXsr2Lp8sM1R
yALwULJh0/nqT+mu4Fg1Qz5lnTR6tDOuX05PHgXIEqMrOferuQx2L7pjn90D9Dil
JLma993H6Abn2CnxDTiz0WN1o7OqoOF0jpdJ9mzQmlCO/AX5QjEfW6/I60XeuBF0
N//JHSYuDTv0J1Dtx2HeXdYz1W7JVvN0w6tXvTJaD0paDhpTfwydO25aLaHHVc7E
YYcAkdK4qf7h7f+7kUA3ZgWvpo6rkVtsvwggZ8dFD3ICXCvhB8zoXWydyi5k99YS
mnHeZp7tFSotTjzW/BeM5S5x8cu+5nGAcTwc1Tx2Cnhbl86WQPpKjKndPyOxPr8D
J7sbx4k2Vk8d7nqTkQyGhZClcm2yh9LVhaKNok1vrrhfzvBHdjTZ+8x9G9O8zhXS
qZ545HkG8sGKA41VK6ZXRbIjf9OQs9aWKsGeDtWasoJrt4bgcQ/jZCu7jOLyOJ96
b1kaOr0cGODR+Axwab4oinWTagua13IyoMJFQKKmYIaJb+lHWUhqEE2/hKR8wPLV
nvoTTtT0qdxAhNLUPzPp7obqMXDE4/wJ0myIPP1vdEzWEszJwjWnMfo+hr8e9emy
KtgswIs/H9lGqScdxsbA0QwULqXOMqQ9G9vIMc/v1Q5UQrbv8vKsVDbtZXAZlyBe
6oIYI9B8t7+OquhPTWYuXoLJ/efz9A9h0AMfY4lV0MyO5i8JdB/Yp/unsNf6TxZq
uKh/ZVJTv9XMS5+mkrBdGFx6WoWcEfsjomraINX4cluh6CNbpcZa7Afg2w99s4mA
1aJi6nUo3vtvLQMEDst0l2i8n3buR/YIqJzfwBt7ujCGsEEss/ifHoV8t6r+4nJG
TlHGEWtI8l5efzJLYN8z1MZvAkT9hLDd7j0WzmVQ9jmcocdpN9L5/CSWep68Ax0Y
NzuFAG9vTWBNFkyVPhCaBNQFLECd6WSlx4nALdnMLnts6WHq8qsbFo1YosGGxCV0
XKeEGrRz0Yp3iecUZeVPN6D/XYDJ+6LEcEkWZMGNbDgQuvu3ut0i2Txi7GOIS9fK
WF5uLLSQ76lsm8uUIlFnsawIpDUCtmgWVKN6YdRe5VLQ5KWSmn+XBlNBvcVfSvV3
CnYfjEi4Bk84+O8I8S0pC0uQdsejpw2v5Qu4K2t67nsCZ5f8jiGlcG3TtRk+wlKz
Mmbn1rWyljXjeYSSLENhepdhQLuqO/BzAATyFRWaCbkPLobzBvrlZ34o7LtHqsY/
b3GnMamAc1eXmfJDoxoUgHOIS2kk+BVxGqgRW8i8k0KeaVDsT/e0ZHzohqXgPs1M
wTAUfxuoAA2eNtMJR57HPRqzvk8WILD4GL6ZubnFiYIDNtio41b4GB5E24JFbSJs
ReNoJ343g63jTd7ggM76lBof3iNlfp+zfCeash/CTfWOuinWI1ftY/Atu2ch0UIV
ra34nLZA2qQsc733pzP4IeRrFmBCS3CWH1PfxbIt98sTyZs+E06w7ME2KRfmAwv9
1mUSWz5Xjt4tU+nA5Qk3dGtxGlyhmgTjHubNGYCk7M5U0ubu6cFQcOCziYGzH3iv
itlztJlua/1wORqGvtQ9tmUX3GU0g0BJ3wGU0mK7KAMoNaNn73r6KTUuWRt7tS0d
iSAeSk/Uu2aSkLq1gbx1ssyGJuWFhm5X5rCPA047Y3RS/tr3FkseF8vIcsuifrzU
Lcio5guFAZaK0XGzKz/qQF1XtQMDFFp8YYQT1nmLzIHV7H3v8/rHs5N+n9Rq9XJA
n0X6n/Cg5POLu51QLV/opc1OcuLlh9k9YyM40KM1QbXeqspnUFW3gy2Fbb5+sPwO
9z7ka2+dsdmQ1MIKr4jjTd63oyAcfzj2DhiA9C133gi3j2cg34t6GKX9LFkTr7TG
VHu/p3MHRJioqc6ZZBsQRpZ57wMdjT4OkbzsFDZ5j++my1g+bS6QPvYa3YkY8sBu
t2y3oKJeItwwYHV3hktg+C/lRf26D9zSJhYVLS7KWwNqp5QP7AZfbkateOl5kMp3
46o89b1f0s6poX9LINO4f9DD5mHONzzyVQsBkBL8uuQH146IqKYUp1caxdbgJunR
zEuSOK3clnh0lgIg9TiX/+aTtmPdaCg4NPAgJ4Cm1Mj80OUu6pRrPQmtr6jxCmU+
e95+0a/goDPg84+1lveVCpLf+VbVeILWeBqZfkGcqP+Dr9eS9oTESceXYC0k6gjg
CU6UhyZDx3r8cXL3kzx+TQ1f02DjF5H+C4XmoQk3CLYn7vOFrmN8B2hWpPHg0uVF
mck2pY81G/XldUv+I9NjY/HEkq6nL+jzjrEi+LBatZyH+FT+9gNqHqHFcV2Heiet
BxXY4k2e6iE+MYYDSNT0bOReb0tDb+CoGZqVLf1Zz5OCQcQFmVH9aywvV3lau5Gw
xBjuEaCbnD5gKcLYX1u8M5FQzJAlFiPvHbbtPltid9/gwBe36EAhU74BCkZ1LpKk
GPUvuEJOH0BANVyAnFTcoB0Ev9I8V+JL5yIp81q0e+mYvk6wO7+PY0I+GhSmuPcJ
989dwet4m8dB63j+yUtB+Kx2fmriyQIDWqQG3SSRiXBE0q35di5SAoQhIXvqLUUn
2RKZgDU0j0LFA04S8+6P817HqUpxNuzaBDef27B6YwxOVH6Hi78ENzZHI49g1Wm3
I0Quea4dMUenJa4K1RCI8muzjRBNJoOMerRXNm2tdC9V/vpWAbtWqgLH7YmyWNTR
7LpkU9oxjoYiNznzClgkeI/sPQ1KbZDnN2WWx052iXS/wgsVZwfNATzDwFxZ6RTz
jLfqjBmvjtivHD+IdEvFcm1W1FXhZp4UISwEWh7qGUnYHKyAHmarJhz6leOGW8hu
SvdkcNx1F1N9fHHvr6DnXo/2bWHxSGD1a5skYF9C3lyh5QcDoyUUiQ4+l+S8mE5/
H1mIu5O844oKy13iOxr8UaECLSNgi+ocx7xi0uUCdkS0Evmmcvd0ZCUy/zeqXqvv
FfOMNJ0DJ9jYHPVD4NvUpr1wOKpNHyhAD7hf3zCPr5rAXmUFPUVsG4jqHSxmxYRu
o/EFJtHGLPYDFNrFu5QPe/13Qoze21YsiAy/wwHy//zI/sxfhXpW49vy4GarQ3f5
J7ux9dOyUeIa/U/xOFOoUxnJ3Wz7gwdQRJR1/g4XqNB/t+eOyuAoiNHcDQ+gTPug
7Rxf1DP3LEye3m7JMULyRD2pt501kwyMpQZemO22vnrRS6+JNknGK2i13yYTCX8t
6vgUhJfG4Yl+a9vyQWkg3yAUKq7hRWypHou0uEQfF0qy44dp+kswymW2fhsEcj4D
+SuqIJWExd8paQouyh3wu5J+6hbhUZyY0wJ0xSu2FdjPFh4x1KfjB7/kFPenOvgi
magPKP8orwCZlPO2IUd8oL/dlDorfz+2E+T7+El20PihhBRmJkoSu8iJW3DKdlIv
CoDzadW49O4ka8t6pS/HYmjz6grZqBrfPn37ssxmDcB4YpY0Ja6faE+ibkSplzhX
5PJ5Znf841qg9yjGQKJlzfutyy9F09MFIjm+AW5LvI254ygvQSK63jOKaE6DkaSi
FcBMmugPuwJTgTCkCvkYMqfzEqLkWuAG4uj6WDurRzGI9Q1OJZCdLu1ZGNMBgy7D
nKeFUB2tOCoMoSGX1kHmIEzfm7qNIcTDhPw8sfgFr3WUiwZfJAIa6SRyT1HIHFO3
eYbE7dPz++1mm3DKKNdDe/e/ZH4T5jTWAhIn3ps/iT1cW8ueOnaiPcrbBAQCNOJa
me5t9Xq3yQsADxaK8kvkVewLe17CJt+q0CUxjwM4Ppd6b0WqQmSUUB+wiaYh5NgS
5ivpa5Q+t1zYqJjnqc3dJ4pH5mW+PN8TbazZNH63rx4ZqK6EV3rW70agy4pYzziQ
tpyImc0SaI8TzjCr7wj6LkrP88OEFGnFxVNytXci/00j92W7Fkyk6QRqjpKgVrLw
4mGj2XVTvMSqY59QpRuHKDWep2Q013w45Sg/+3xYfHZxrPvxJr1YTEbCDMFGTEMf
xKmGpKcHJuuc0HcW9H40etxvqDydJj1rceSJRVNzxI9AGhr+U7xVxP99xjcZEbBb
pv/aDpJinsnBilv0f/x+4M+hsyvDD7ZijH0jvd0NqbQJhf4N7BCQRiNF6qdcJG2r
rG7Q1dPtVgHvxDwV9dv0MwXTYwCYcYaJezyvOOkYIHH4C5ka5wkzgEB19WGtg3gs
Ly/cJJp29w29R8PPj1GYsWPUW9PMZrxsUI3ZX2Z92KtVOfGoHt6zbCC3oAcr+fkf
bBzKKMZ4mjtEtpC8q6Qnv+MOfN9XDpnW3FYoXg2YF0stWhFU/CzukXDlls7wcZyZ
t1hu6aGUS/bXhRHrYcv1AiPWdhHqboPP5CgVEafRxZQA9goRMJZ3ciblA/CZttG8
psbdl4QJBG0uYqSmx3AErBacBnKLW2KoKEIHJMCP4BfhokjlZl6CRi4S2NKFeTOY
YBGob6HTQXC5VE7cNLZYHMRUnOlCYFhfXKx47Yl/VmtT9Pf8aqwttXfv4UYMclP+
+jqnR4htfYmo84dHD4/7+byGzP9zrmdw/J0AcqXdNnYq+TfJp2v3R4VZTZzqegCg
kkAatuAC6H6o3oYXgA/shumLe5X/+dmyxEI2P/dK8p+c4+80jzcVkhNetgsFLBMP
O/uZ0g4z+N2I1OLdnUu1HEa4q/OqqvRKHuF3ZJrJlG2N1eeriq2ELW2bjUQO9/sy
QrNrqSqhdHdXZWTtpN9uP1CpMv+exoYvH3RIogj8WcNgoJZr3APkDlX8FPLtFrxO
VkeryZU/Gmd38rxqXMqszMFRkZp1z6YKKtgraysVSmll4j+DPdMJYKAE7JLOHujw
5NYIuJcnujUtwOaR+iwArnFZMTA6NBU8WIqFSKqwLgre4dgrZ8P/kA9EgQ3+n7yW
UgSa6WSrf4/BQsQdC/p2K6gqy3tX/fobgvP3dMwCCTJUr/2CqaLwvPHPvbd/1zbF
0sIIpPDVlBrCEWCSEuQ5TC/n6N0jl4HOHPmbSAntEJPgkt5UU+Ub1n1czrM8pSyD
0uUs5L+CaOMpmk9f4eu5ZFKfnSmiYlrlHw1w3KLzhmiD6wbcDV14c4a4dZrinCOK
cQoKXPUuyohuxkssc/zJA4K/iu2eMVBzi/MRYgFFKMkPAql2uOfxT2z8ixcR8YTB
O8axX/1XNbUiPxSEqCitqdOvsfGLTfd3ht2A5vnuxn0gOcQCMPMjqDmAS0OGg40K
vyy1EnWZ0FLrigZ/GNAUEv3oVRZBE7vJ4zR8OC6GAVYM+922/GWwsWMz0O+HDbPS
+zGNYIAwtyr9UQnyCv3rq3j9/K2dmkwCoqlWDmVdZPwxsYz4wpZGncAqB1cpjahw
tCcFTVuSPTOaJ2cO5fHsAmgZebIRorynYRAihyFm+d5RnpGC7gl3yoO31ahpW7kD
5g8gbZgh4kUZBW5nLVsxPagq5GCspA01CJNtR5luP9wEuLQE3g7Frq8AvQHoA3b0
njIICZObqYwX8A7wxGNIbkpn8KMx7RTpg7iP3uzuyzIaBmhpepRm2QhldMZu0ZJW
49t7SK3qJXQ7me2nD/xUHnD/4Ou0CRtiAQWaWH21Pqfu74bEBii7XMaUuqf8wvgY
tTHUBxzeoFUH8G3YwTuJOdZsqEyTcnOFneQE01L0LVmnQ8PybBbGHmFgPeen7S8i
s2jfB0fra4LtecAXj0la48jsqGmvtk8mVs46mscnEw7195BZuqsQ0yof+/aXC7sa
s3GXo++uhYfFEz79lHKzocdONSLTwu/GIP5UB5JfkvhJwKLrvrKJv9oqB9ODdgWN
JKrDWJqDA1n4tAOO27ICOSzjJaeGD0Qm3cEOwvwoBWDA6e7jiJDK2PFU5s2gp3aT
CgyudzxGwdZ97IK01dGe+ufhXiVXdXpyrRRL8rNM97BSAR8/YPz65ZinJ0j9wixJ
SmcU+CoTq27vrh2RfZJTS4C48l/i299XG7JCfo1f1bqrOL5e7uHG0S4VizBCDy/4
+QsObDRu2S/Wxt5SbfzgUM4I/D5/Hm3nTVjj75aY8my0vulpRR6prGPlGTPDXXwY
liwKk4ItUDz0WF7PnJw5ob2j+ZdHHrdm9qhOKpL/Ck8gymL/wjBPkZRvjXapzKDG
8oC4Z3nNMd9eKtf5ZJSpyjOKd83ECOqHZIiXFnHf4hi+CBNt8c4UCcTsUZyy6jnx
GFcVae1iyOWWNDgUEpUEWyOqoss4Ife4dJgSZ9NBHunfgjM2sSY1+VCWD5CYBSL7
nCIupHRLFQsXzhWd26/7DZxLuxbiHk5WQCp3zx5Mp7yK+Gazunbs0ZiTRvt9olkU
R5PQOuyXNa8YE8Bl91zAdepPgf0YWiVTcRhH+iXXos4ESaeMawFZ8EyQLBXD5SHc
P3p4CM0HgdT0ulOEdCvh0nH6qabseEsFy8trESiwDpEyoaDngrEdMX4XFmWFGXgC
zFJvkZ0AjzHyLzC3w9H9TIqaaWjsxcx1BRjk1b5SbH9vXMCKKl9N8TdhLnn7aEjQ
Nfk0oSJZfIZIngtQh3HCvU1u9ncoC/S+B6Su6jUtQ3XQSrZzPYzcq1SyCKX4mGNo
NHuS9Kz33/ipuq1ACrKXSdqCfM6+PFqi6rXVGtp3kG4In5SEPfAGwWKQLnDNQ4lA
hPKk2bhrNo3hFs5vLRhNolS+g112qgkH7UGEqHkRlC5Br+q4LpTLo0j9b57pKHiB
EXnMCXcifoUndofu+9Cgi2rb2vdaz9mi/f9oUAQpcJ9EBmn+f6AGA2dr8Qke8pPS
2zbjQLniVIotHgrWSA9Wma8ZxENtYAmYdUjYlt1tiAm2EmCJBVxe/jsPKzjipFvn
7e9FvJT457mcOtprR/aukTK5foxWrxsvWmNXkCKgKA2rJNCpL1vmNtHPJjN5xokW
NgKugB+bq0B6rVCl3etDPqJJGBst4r7bdvTQJ5TgU83gghir92WijgOe3UuGSrKq
1/zpmjxJKRxbd6W19lMJ1VUYh+B+PIrHWRhNR+TRj+ZYEsx7iXkBndv3sX+UTw0i
MWrpFNmZOpbdzK2d3iS3tUioG9Zk5beZEn1a+O5BsGawkrI3NMvsCuujcWjIlR8G
liV63TXID2/3Q6A2dNan0TkZsTEWCo8xcpfrigblZBadb+MIyCZxY+tCwySXT5LW
EiAi+vnZaQp8pEOQ3Jkyn1yV5qwdj+ozC+9jZ3qvEEorXXdhTsXpH6NHDUahMJIH
v0xL8gH6M1IC3u/sK/UosRXlAyEQ8slVTZMRbf3jl0f5kIeAp7P/ywcrklQeCIn1
fHiC2YMngkPGUg5zQRbAjNEPJsGfrZpnz/UsN7HKlaTpN/Bx3T1LTCGhpO85QdGw
X5POVicTMsP6cY2jsElOscpv1cp61WpFYNXxNzFt6032VACWZSeBVnokuVila8tM
v/934uiJyvz0hW0Pbg63azt/XyG18KYSwmluTUM7PrLIl0Albg71LfWODpe09h9H
ArAoHlVBUXNsFF3yZ2Fo+vfpAKzHBiPmN/+wx4fxAUIh4oxk683Lt8Azcmw7dgBI
Z2EpYgRk+lLxoEKW9qTAd0lJBW8dRzKfe1LL+NlcAUDV9TOHj6tE3g+3A+89DVNu
OikUeQFb9tjalC/6dOGwnpzpdhdjzdaLo4177yKlIcAtQIRIquhjci+z+65T0Q2X
9lEWTPJrjgjHw+nPKUNHycTkJMX+BZb4N5RcDwSNCrEIUAoDEq3zW6ktF40FDBFs
oLvriyM7j119YVNATqPmm3gKT2iba0YXcbld3Ic4vQsVk8x1zGyzQG0or76+SKvr
M/2GJDxWyy5Y/dk5dv0Tf4Wb6vG5sM+OP0OevSRvGIV9BNzIdjyimwO1jLHMpWpM
MNacKBLDDQUPu6sndWvZakMz18akCL8wuRPItjIYVAroLuiCarnRjyaPeyzUMGtP
TUvCssYTrQtO14m63x5Ps720+69ak4djojcH6CUXuHbYH2jhXfIy4BgfDzMx1gQA
vEIrXvoS64Shq27BTC6QC4vGnCDCHm2LZO9CRm7LpCsePMaWf6C8EFk05IEC+Wdt
pwymTT7Y+K9Xm1w22uD5jwpXPo7qsMjo1ikO9FQdZRqcMLbJVy6OH5i/DjTlK8xL
e1Y9VzoFU0pQr3iw3xYi5jhyd77VRaOUQt1GDkZfkO/vRezdNBbOsVNNRc6Ldydr
QjhwBZhEW+u0toS/PNPHg157DaZdGu1VVqPFg7EwjeGtSpFPhVy3ggu7u32qQdho
QIjgMQXBi188SnWLhBNNSawAK3y2ftqgb9JZKW940xJRy3APmAeWr/r/EPRcEENf
69wt6rCAcgkW719+3kKhsloCInvH/dMVcnwOaXvLZLG7B1J2ahfaW14qx7XB+kB0
Gi29OzhI4VLlGj0mZBYrcabSVmJofGw0hPTdAVOAgSsKcffYOMXTgsiP8ek6gc3w
mByUximOy+mPRuj6Go3PkZhUujwztQZmL8yLQi4ioBzglYGlTSKgqCV5Fa+Ik0dK
9eXXf0MjIINDKpDMAymY5DDVpE9Rg50KxN3S2yeyNWtq4ajr8rlQWl2JrIqvYAtM
qoH0k3cwOe1mIpeTEtaXxQ7y8Bu3YTqGXMYs8L221LGlm35YA5CyjNdIQlMVDsFh
2yovnivwQuhlvGWGrPydKu/3fDWj5xbT8tdRg3D8furGMMPYAxweqhMe5Pn0IPhS
WlGW0//lRJNV83n8eXLLTfQ6scTVAzXWOQAi5JfIEikCsQ/vR5978VoyzhTX0C4X
NLd32fHp+V6fzwumbcfeaEPV5YPGmVVTVt6uW4qDLYXaWNEAR2I+uPyjTSD+qyxo
kWskEbRPdngEG72jezKL4HlEE23/ICtrtV7SlSVkjRPbvFyU5jbxz4ZplVy6dkcV
uAKoqdGoBo4I5mUzDZacV1X22hBPDZvSYJBoW9W4T4c6I0Aj2+xxtVuO0DegTHoq
W79P0BrNin7BjW1Aqvov04+XSjaXwNv9kXrpuSuY1Zo2HglEc7CTy/nhFUJzWHos
bZB6UKaEMnGffPSD/rWV9GFSxTXJf6dUichS+oTPHzdeekFACqPci0WYp2GhRShY
S8sEc37+XACKIhjeUmz08thSBbxRHRXdx2xbZgHFX9CNLy5ulfOg3oXisIgP/ZmK
QT36BwXf1aT+ca+ldTFDGTt7Yg5c9USdRR0d36ZIB0PeFXJf06AWgm8l9ufqNFeI
y6gBnmBEyfYvp2be7ZfdtuyXu8LqBkcGejSOL6aAvvNh9K70QGTqMpTHXj2YAK7d
3xNZqvLqEt2V1EfBlzgIowbBMHvCGuaYGXW7LN9Cm+BaEb4oVnih3X1WmblAOW4E
LvWo0+LbXrxjlx/xGwlaNlQn7IpgP/TAI5qDvX8qKQ52tw7BX34IFffwqTYIJbVF
/vCzWUSctI+1l6J6U1ZeOWNvyTgm5lhxPYHIcrxeZDl+VrL6gAwgnXlhEIiG4zJ9
WCDeadrzhYkxVjHYhoVlW/bI6JzkpJDJBj2+EjtmQ0KN0IGvAn1xLYPOPAbnOp8c
aoi1Mmmo0p3gCWA+HBGb+N7HFmVKLtcHTLKli5CtbMwzxDf2Nqu+M2I4TQ18cZtt
MMPhrkXxj0AcmheijyB23DH8v9MzXR0DV4+GtOA3fgtLKC0EZzEL9lxq9rpVfwoD
lZlGYTQt3pTLg8Y5PObXS2Ebl9sAdN4V5NPYeh2IJAoMOMI36aOUQmD/11CPXHmo
8Aumgk/8iwNQ6jN7q31NeXiOIQC1AyFrHUhqZ/OspsqFCddxooowAMdKr63YQHzK
wS7XyoD3lt9CvQFJXPVSOJyiOmhk/klxafpI+e6p9WNVdBpgtG1mxEd7dW5tpIAh
OM98dUaHxtQvrHxIKGu+BgtdaDCTjuz/2itr2GOh95kyXLmQf9218UvOevGblDwv
/TBY69bLWsmhF2pY0zbWc1zq7hjwUZ+an2MNN8gDhmEt/gmhNIWJLOKm/ZU589jh
OR5uKckg65lJKDAZldnQkS6WBCA3fCu/xcdLee4X+r5ZXY9GzGkx2yOvfm+MB67e
npBixl1M6e4iZa5pXCf/W+85Xzka+QiZICQUeOy7qKX4c8LWTJByIIap0o8PTY9t
iD/6P1EihNucFaHoeWMOxizs+4b2r14yEn90bh3ADM5fP92uo6XJ4JLrS/2OWmtC
vH50BBVubUSW8KPaawN4TYoCaQC5aJQ1TfOEUX7wWLa4l1cVm6CjA4zN91HQs0Kl
GnS4qmVGcM225Xq7SQjmOfMXxuMMgJhcrF17DtWAfAy8XC9F/p/btqBFhWumFqtz
eySq4mVaySY+pbrsrgJJqxudSDF8RN2yq+Y2cUAu/xIYQEH7rSCTyg83hMUCUIBn
UJZV8ySutOeJOuQaT87hKNAsQmEhCUuMstd2cOedRqr3NAnnC6vAlCQkrH+oHuLP
wHXVZV7T3Xv6C3lBBhuMBmgNnJ/X734MMwbpCaEEPAl48MoHL6wXG/DpATKPRMlk
Eqen53wz8lz1997eKoq2fcqg9paP4ra7GWucvKGDtzYGDayJguFFeOTCd5qlJok/
3CLPpuIV47tyTpGFR4LFlnPNzuso5fV6Anc/evHCC04fV09nYvqx8eLuWpxpzobo
VCGyv5q8URHq38AMaXFl2ZcU37lKOFNqPby9MhZeLyP/ZJZ12NEmkh8YAZ2hwWTy
2OjKBGKZQ4lDWHwHXyaLQMAUoVdA2gcAWQIQnuzGnGjPReURt1o3bgYBW/1VftsK
0/dEWEyuTxg5GEWanKUzPnRiSZ84/VpDB2xetXdx3z1a3Ibbo8luAEVjxkRcAVKh
T6xGaaI6t6a+c1r6zWmnQ5cD+2iN1Y/GEGvdyuwBGVz2viBTvVGXkyvVxQBunIF0
+aECDHKC52BYjJP/ueIVHD1ZqQU4ZcrOOZccT8AGGaCWlhDjQJyN15svElGHNwj3
kLNM+vj2CEyCSATGRzHpygKAYBqR0Nd7JbMWbJVc9wds2YF03QMCZbnaG6dXxNgM
VNYiYhxAQlZEFB/InN7UFSZRrPvG4lDQ03dzAUUOeBzbyR5VLHW2P3i588BYjA/R
xtncR6hZsxJ3VTMVL2nx+cuxYpF3TzLWucjuLNC2o7ixHOb2ZAiyRe9tVJU+cQ4o
KgwSKq+R8hCI/osSLBHCcePzYMUjVVzcMR6pNeKy5xTjpZ8jlbQ6agmBulWWECI7
eNZEeUrgX6rjTxreDHyc9zAJw51EQMcGiTMVs32uCYaoC50Hb4g21W1qzF+DpH7J
w5s6KcMTxfQDcQfSs3iJH1O68DnIrdUlNeL990R5kbSMdqLeswK9YNWI9rLKzLHR
TXJwfGnrx58aQyN0Hjq7M+8QApIs00e/BE/+WII4t+x3QKik95y/j8eDYGZyQU57
Aoe4k/0VIZ+eiigNAcgVBTad4zPnle1mCoBB23g1Tl5dtnmjJppZPqmSSQGZGiBo
39Rz3NPiQmopoJrgaTx9MDqemEsnjxGvoOeE+Ux8PZUQaFzRoQo/Jq2KOoexUx7Z
kNXD/ZRr+R8Fab7vHqwInVKBnD/TUcnjUnpzbzAfe3YCFU0Ix+e5Yy6NMG1ZaP5A
aHg5M+26a0wOr+g71avVdc2tTWcpecFjlQkOvEX06olqII13cmUYQO9PvyKvNvPY
Pa//lw7nPAUgGhOIQHfiXxBdHhzWOBqCKAvVKaXx/mMGBiQLT4Qusy6ttX4Q6euf
iM6ST14ByZtHm7MsHZIN9s6oNvLa/DVxZz5bJsOQFk+qjvPAHbiFQiAskLIy9HG4
Y7Sb1l4xDZyOFRUSIq14IwEbFG9kOa8oy56Pz9Lc8d7E4IHIzHaN2r0iU8QJ0egp
hZScjst0K+GAjcnUEaiHs1/wfkqzo5tu0zLzTNzQZW3Ix5vcKDjHL8VGQHTxRF2H
3wl6j9K+jB00DqEqo8kdgH+lzIV9bsbE0Xwz+vMKc5QyDsPqHII8HjFe4ABy6mJw
vqPhhdaG3/r1j//gIy0UJg3DBymSBrd8I5IzpERM9o9mdMeZhjZ3OmB50txO4Ob+
OXR2lqZdiqzk5yD7U1BJ0kGkOictCzqooAqi8sR2GUxZ+4FTGWZOBGKRCs3ZoON3
5Dflw4QZnYkuE/M4COAvwHSEqJM5ZjWMhT3GSJsNu1//EDMbcswy9RK3ZnLOHvyn
WVyIE7HVuMc9WYTTPWPvsxupf9ngoQj17ny1I7/z5csm4cInJTMg8luq2sVWhhaZ
615gt6XU4WddzSlQWQ4LQW2F5PZLoHjgVezj2ilktXtvmtaCqDg35DLs7v8Pdk2T
cU4sFgjO+oRKJ85n3lsn0Gz3jot61zZJi0HT4aqCierFp9yflPbroJPbpHdZpkIC
EyNGTBH7CT+aZqyxLWzQdxDswzAzo0sUNhpHhWsLplH+8OhVDpqH/MvdL8JCi8AD
qA5CLrKXqyv3rDu7XNR+kP9GfB88SpehvDifs1w9EV0=
`pragma protect end_protected
