// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Hc67KKPCdg10uszpkAkfQV5wpKHjAyMImmeZo+5raIjyYtArk69rELV8ZfTL
EA0+U143WLfnIj4mYoItmxqDeo2LZNQDB6gPqPfJuMfOns0vh5GtO1+X7wFb
X2XWJyxKPlsz0bLVIgTGlX+ax1Az7zDlNB6oCyX/vuYnjXsbZZ+B0oZQxMOh
R90BPZyURTzxAwkyEUwVnJXs/Jyt2WFT9sHrZ9iauTh2/WDhoMG65OmCWYxI
NY2aAmk6y4T5wU2JmfCWz0vcpyj88RJq6l8vOoe5mqN7MRI6i2jQwJvEDEqp
7X1Us2on/iEpFvGqr1i0ydOcQYI3ILPoCAFXiBzS1g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Z7DfVTyAVA8nNr+llDc3iFUjju/qhpZvefHcfoA9Xgmg+K5SmEbQis5Hrl+1
0CfT4EP932sKJjPGVf8st2gHtDSfWFeThekLwBtj+eMo3OHseusKBm6iSJmU
0hYEHz5MsJ1GSoGZGq892DEsVrxpVToG9/ToBvnNByvrsFqZD4yC5YRWvnnc
Y7DyKoUVNS8t6nP4ZzFZKQ83TO4vhGifgS4sdBCMn0ypP9HQD2ezbsGzYgOZ
T32KDrCSrHx9miBGRTuSZ/VYCRWLzVCUkQSBeiWCtUBQNV83f+ZGoOkRaCQj
A8ABi+Fkijqkjl/UvzUJum1S51LNbYH3rK//LrfH3w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fr+bgMgWrR6GAEwpZGF1aTPt5Sqct9seOIBY6r4ZQu8skT3fh8u0UneQPXer
Wtr9XdXIZUyKaY6qMDjz9jBkDFFAgfAEdEk7UmT9DM9M5V1FzZ5G7UYjfBmY
3Gn5qRaP3VEP/EV/z1POyKCcQ9g0/me3IFXrJRPJcCLT9saCg2fWdmSX7dkf
qEf0v9eWqmyZgJawsWz1SVfx5CeUWg8nv3+3MDEl4oUTzw98yq4eXj3af6Wm
kwG3nuVAh+M63FkzKzQgSsQCpGO5CXQwQ8MlUKnjSlZLteBSLgUcUIR0WE5y
w4Pzij52pamwjS4yxr4eUAHHJ/4U9XT8lvAbixvozg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JEurxLnf55Lp58QJ+gT+5N6CluOoEE4zJ7jVbx4ViMDBiBISm3wt41hrRx9o
+ipHEWF6awEhcQ1H8eVp7rywOy1F0UalFXlTi5LyIMVR3yCSSaLI8VUl9Vm/
xora+Kh3wZvtnCTCzAGIEGnGJ5TRDz6X0IWpFPlicqdbruPEnF8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lBaQ0lDJnJDgecbkTI6fZl9cnMDJ1XIVyrX+z3dXMzI7lWY+ENhKIGhAtr4G
KL7JRRyFfKaKIVDEopzbPTmY1LiqnXStMC15U16/KZarp+nvpLzudUTtqWVl
GEmBdKlwnVZirirch9OC1Ir1Q19nITRCrRwyDvnshmuN3Wvy3LmEAXh6py0R
/qUsGvVuGAkBDWjQohFfK4yjF4Bm15gmwxITaTJSQDTqXxOXA5UmC2VXnyxf
MlicYv5vKRA43Ix7JK2PhoFJ4dlKPfD3nHeKiufM69rZNL8QdAYtkdZz6Bij
EGm0nM5eYN1FXtMarXVlDfdbws/S7x2Om5YTjhMR4ieaG//cdNBJTBaci4hj
aLfEF8SiUJxoRwQ7UgzEvQAylTMTABTZSwbRlf4N8O6VVn+XDmJ/X/NGcZc8
DoDIwIMRrYhfhyM8Oga48IZkWTeaOglm/UOxyo0KuTygk8vJjfFqfoZ5KtCF
FpqZJxGab90uWHq4FZbwVpSd1VPQZA8i


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rMgVPY22X7tF5hmtSpHM8vzyI1DgS78RGVuL/VrJcl/tRu9nTd4sAoKeYEYS
FH7QMmSmiRg0Y5aUrASazWpsZosGFhUluukJmSrXJuzgQeRrDNfusSmBDTMs
cLUT15UMhtIowz9J+ePZzWtZbufAWE7c/cgJ8lCsGKQQq4IHsJ8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
brNwA0LZ9vId9Xdz1uBByaioBLWHoniiKP69VppkRFWDH6aYzdSNETiN/Nj2
89Iaa0xXipKY21gAPsZmslKKJBw9aDdHwI8dMYFuJwNAzg2ua4TXpeMWkCQr
F7L4l62Ol3fmc2hdgT0zTMZczhQmchPxwP7UYT2QeeQEvc+3eLc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13840)
`pragma protect data_block
gBQhgtWP6WAtgvMm0iObiTefkQCe0QgvYNf/eqYRLK6RRkcNpumBPbTC87BC
ln0g+oaoVDJ1Viz2Lib+lV809ttTQu1v1LJ12SVgYGKjs7+f62+dgSqWJxNK
ZDdw4cLc07qx9gUwGGuByuqd4yx4PT7UNTMxLB2PID5GDmwMzX61A4Ra03gX
GkO808AeMigxBXurSHq7Y16tZoWsanRKtqBBv0P0Bejz/GFmU5LKHQI0WsB5
l+uL7/YC7KnwX0iCsDKW5qHgYg8PKuCJUjP9Xf8CHVbS5CT3c1tL4whd10EF
IajVvVWfH/Avxop5jJC0afmrfWOTmnYgx+stDtrSq3DTglsAG0yIXhnfF87k
P30USWLgYGPBds/FpRhNftT8WVRi2nC9lcKUWvKkDYXzNIf42Iba71l8Pa3b
uiRTHOsP2xpP0teE6qghdcwTgaQF3X9lnMN5DhLkDQUJ8uuWlIeV9+iwoypi
GbJg7uc6Cg5IR2FDLWYHFhU7X59G8DfGzB03Ip7TmBIdgSvkKKThs4ApVpRU
NED+sWAosJsmUHIxrgzOrnWEmaR4mjGV1uAx9QLPITTAw4bj60zfWeD6vg1i
32+SEgEBS5qbBatMxhGFOwO0p/dkCaW+TN+KJSc2kmLe/Fpm99yPfQ2ercLZ
HFSm2a6GP4L/3/4mxLTg8cYTGu8FRpoPWAR2N0B2SLyNxvEUCEZGKf5pIFGj
SH11IGN5jMYNKElRJMPJPS6YlHJps1P8zaszQbBgZBdRu+OqPFgFzoSqY577
x4YsgvKrDxMgVtd/XQuJR/AhECZoZyy2WjnfZAG4YTZwEPtfaVSPzLELuojq
Sa2cdDVauRY0hB6BHpSLB163/I2XmTU+unzzwKv5/mjnkX3MvivGKg8u7LQA
o7NRYdJHc/H98VXkVfPqnFE0mDB9h4uicR91lcBaUfUL7TKPCM6BjVsIyS+S
Uas5eFTTicnvDurfF7Ha7P2KYV0OjVMQZ2DjIJLei6QohEvkvZG5XzcmXjsT
C6exPXBkRGGYGnoNPDyg0vxi7LpOWypniae/k03vd/aJZlg3kUUCiqP6gO5V
uWs0+lg49041KE9p04CcZn4JIVQLqQPtu/nK76lks2c3a99y1cMQ+/VcMvdL
p5DvOn8dNcefwTmR2F9v9jJPHfxBOLNZd/gocX2bAOYiEGcCFnu9+U+rYkvT
2ZE/s2OjcwPA5YNLcXtdyam/fUgh7ibjAuaQNMw3TI8nMG3DrVJuDr05+htG
HY7aBo+ijTyKo3s4tRcdf1PTIsGR4cjnVM7595rHODuMGUgQOgKtAe6RoSBr
yY86WduvKBZpj+Tcl4s8oT3kCZ9/AIRVCFt8LvdDi+kNX3LORTYZGv1hRC3/
RV2LUrJPl/xyNA/G5T7+8yy20P0jZUYtC0CbBn3v5QFa1ZI/SFRXo3nQ13n/
EuKpr7EFHdts4PXe+0btg07+INmKlmV+Ra63ogAk27FVJDkkCb0oNGqD8vW3
yAnos3J38vB8grJnEamVG9zXFVSIUf7PQdjj+PYu/q8otDqXwztZ3hOc5yKO
+XdmJeAhdBbsHlL2HbW8LZnlGQDk/NZp09TQ8W7fbPKAb8+hi6bY1FdB9LS7
rXthgvTU2ENZR45fS/7KJqTo8QghDhcrsDLLd+u8j0XLkvPRiy6/d5aYpc+T
8qhwuue0hommelZJh9XKf+bR1/f3VOcJQuE6kDH4jSKT1XZZJO7knDbK1Ict
rSKLEJlL5bQWf1XbrbxhMUzycH3v4jjqunox+KOmDXANQUsPEK/t+9SRIAYm
KEeHyPw+bxKbPQncVkmQJhprecOqL3AWngV2fv3DeWQlfqyEdZqNTXQsiU6l
qXU26gwdaLd7TfN1m20tp+wne/B0YTwPzFSXgXiPdkAVx516NIQ3Ry8d/d5O
ETNyvY2+P5NyycNdPA5EaPujSqrpxSQSt9mOt5nNCR47mzduQ797ikqeuXyN
+kEd/Auw9+rsA1F9yRJIcCkLWnvnO3PWYg8Dqk4vAMVQrUQXKuTu/Z9g6Jch
n2HgHb1cG3YBAGLP6ettgEmkDPU2GeVpQli/BHuCaSvOG1nCInKUR1j069gX
mQ/RW36u1AkTfv7aBfOrBx7Jqf++GwAdn/HYzmteHWnjPM9klCdjpC5bnwtc
ZQWJlptcn0RBtKQBytCEL6c0Tsw0OaM1Wv82lOGIOIhMi5o6yITQSdJSK4hd
IOBRSBPTzRhe7bvcyygkr4r+OL9p5RLecCyNjQ62UFEOiAfaOEvB3A+Y19HR
+6Jc/gzKxA4X5sOkFq0m8saZwk3WNF2Hs4bewxkq6/LHtoHhD6qPV1Tm68tp
N87NE79HX02kp33xGbs2qaBw9h5WxCJciXmAQ+UZayb7P8ytTm5JTIvhRmtY
NZo7YNN5pnUTeBaGVudFuh0XSGC7XXi1Q7U0RYHaLZ3WwIxe1NRsSVsKegow
d9c9MqNwkB0g4UHXPlWfbZJZSLNmV9I6gOqDnzCREm/9r+2io8ZfKBX4EUQO
OaVPR6c0yqFsOrt7xXsmnBYp9KuB6HO+fAT7nVkFJsDcS47dhghynVVvT/wg
KjQZEWOcocnOa2o1nbZZSONfS3v8hUAqEWoUTkqyvU3IJOWjGnxXQX7AGAjt
uaQ27lb4QfhylDYkbMYgHuTXjalEeH+roKY7BumTclguIImpOUe6D1UP+zoP
pdVwtooyd1l+32UD6YZeZZU1yQgO/O2ZGgYDqfqbpvFxY0H48BVqKoQ/xp7S
5zkX9cSO8vzGC0BRGqpyJ5JsB2Ei+jAxjKxWa4+ovjKngz4K+nickTBC2wVW
s3+IfN5znLpbrD7iRGGK9wuca/cZxEFvcFFQRGkkAE4dC6vZg7tF4XIQAPm2
DKq/jBNICY2TujUH6N+LPzbEh3DNC6YBnSSy35BlWFShd6NUaoXe+8vVHLXQ
Ne1ycVK5T5+6p76CYina63A7Egl7qj5zA5MMeaZH9xR3OjG4T9fiZ3apGL8Z
7R78dFM5wTfc3bP1ulPVU7ytzLQ3PtAgW7qT4Lb4MhJAMRfGLRbc/Jl0jNPn
uSmTuv++663cJXdM2rzvBBEzr14yziLcCa/P0siX4yIaXk1X+aNLHXHOl6bp
33WtPQNAuFM5eUsUwEgs/d7Jjcxs+pg5itFI2iAQyTuxUA9/YCtMUjlKamd3
cK6FgCcpFTXZYabJYL9v1+1Guz7bHtFATXVQ/GN37AXQHwQ4kVhsQb3dPWdI
yA2UqVYmv8y4tNMahHfpuZB5KKhLyARhwoVupv2wGdxjeaX5LekyAyG++WIW
TBjnRcrjgcZdnQdzPI7mvz4rspJz/GmI8uGr6wG1PRcAg+F+8Jn40Rb4Q9+1
eKy9zKq7PMBRt4Bf4PP3Tmd1n30Y5x/N6ZdF8Pbu53YxXegMkszs2msAUkG+
kiz1RIi9qYRbPOMy8tXoRJLBDSVz/v5stk7Qz9vnRhAb2NZHDijn7s7zYQ4z
M37QzrFCKZxOr3Wi+faZCNowSl7nZy60UYzjkYeoNqmUw/Gm77HHvq0gVz8K
7U/EesOMzqQht6Sx/lETPqbo3/y/uBDUijhaCfaLymn6giQhvxtEUi1K5gCb
8E55JORgkRpTbh6KZoRRu6MTrP1Rfkot9N6nGcV/pwAnAJHcvghzT6nkKI8o
+1a3KfOzp/ON9Ov9O5oLIecCmwFZkbewfevbKlt/ZUImQZyxQtB8sMLmnkmW
RBczY+3QUgfNhZ519LdQqhmAzuOEFa3PIO6MdLeXgsdyEciL5GR224MNtJbg
h/CMaS93vP71ehjcK7RUPNJziCP8mwPZbcK8tUvG+BAa59Iib6yvh49unJxs
9MQyIdcFBSU1GNWeneaHJY0HJQX80r5RQQ8tRLP4lIgwuX8agcnkhQwntkbP
cW77Gt1mit6YGrrmGwIdyuUzZDq86AtQ1pPyBWm3OMKlD5mUAxs95acs4tEM
lHw0TKAQ3NBpm6r21n79TD/ZC05CY0eyUtJXqrxAjud293f5k2+ML/YhO5TN
NOlfC3mXXV4qGKP+WYRUS3snw9TVHoJ0gwr+UN6wtU21CUUPORmobPe8L95G
WNk3YNnJHA1/4qPhFkBOEKNr0gRk/dMcONStnbsOBxL1P8Cg6r5EJfvoaRjQ
Fy3xQoXSezuWO8NndT4gHaQevMVYggu3WeRc/2iiJG8ZnJcNuEZQq0dLJCVe
pjFReZyQDhk6UKxGgAPEvT3i+2yMUQhAq5JV6QIcN/mDQxfmF1o6nERSVnwp
p7kl8n8okpc56Z/n1nRt2WDavCKQPxmc7vVmM2MnPmRNFO9/HlNcS4X8mMfL
tQSnFtfAp5Uch9Tga6igBUrSipdgaVT7CHI3Dv1uYqBlEu4CdW1yIwUxd83q
Pk87U0gzqhIbWmHETkeJlYe4g25V4Jh13PVgkACiHCtCX7dvKVUlqyOTfokG
PAItPuDgJVkuF+OR+Zj5vd0tRyO15HZCdqeNhpjwhdYc0Vrf45HPfJ8OpJzj
NNdO+8mvFi2XR4DGagLqr8rEkGh3bTrAw/7H1nrXi9UzL6V5tb3M9wVET2lR
PERhd6Qj7V6TICQJ3sUibAMsQqYeM4MaxLIzLmslBvfrZKp2OpohEjIq2+ag
ioPJric0N+OEoiM9meNGTwBwHUybfMQOB6HSAa6ly+X1drAYxOBGtb4ADVYb
r9ThreDw4abPjcrTgBhiPZCtyYCQR88fOV2jOZHJoKIdo861JdK7T1bIFuDo
tAHlQDvhr9SPkxzugLyPkiVi/9uNcPSUWlUGd+lhs+V2lwGsDGl7CJj4Yf29
Pq8XJvGu2pRRMsfnz4QmHZ4Nt4T3zOJil0oUpgxXDd+GF/7SMp0Prlm0+Wch
ZCwK+ybC0TVx4QnHnHdbrYke5CCzW1c83PLr6X9zcsVZ36yQls9FaOOaWtyc
35RR/UHLKbUdX7FaXjAryQGcDjkcr+Pg2QENyzahMRvNMKqro7RCqW/fx0G6
RVCfqZqktvozm2PBvrBov2eIT+TCcgJzbeJ6K3JvCUkLTX+CivGNhqpdzKCA
BJXOxORr0+dIQEKuDdmK0a0G+gcfpM9+hojhqANUXDs4pZF3keZCIjmQk/3E
AOu/zpjHVNUnIpATkr+Otmho7HBA+BlGueo/XnlI6WMI+b7bphJh4EavzVSE
FRttOEOUc81RqsIyjtfwbQX/BkNNa2jpTPnmOjSYLYhcGbveQ1R70M+oBP2q
BYV/HW3fxv1cvugMaBaNWPYMY5FckYzboza5eXZ4NX/LHdaSEqmVm00i9cpg
TM9n+0KqB5HgYT+D7W4XvtvPLA68BX8OihFjquQmzHlj8h70SAN12W8AJ8IU
SKk4PPwNCE+JUVChSCynWPgm5mkEHoRO99CfDUysRFwfBFL9FuZGQ0Db1BAa
irVrmJoe/0CXzzYSbAo4viy4mDyiUt49T1fKNrFioCy5uiwRBwIIkjTyK0b6
OIRRfTqGmWt9DYKGmyvp3INTUACBPr9jFrrzTlrUTcbmUbb/z5yHDpIAqfVV
RIEa/OmQ+q7WfvAseFndzK1cCjBZLsUigEspqO/GbXu5zykKELIZ0f2xVwx9
o67KQDHcEBjtcbXSWRCIR4QQuDwWU2FWk72uwboxS/Zc6zhI7tNywfPD88Bq
Gv+HmS5wbLs0mQAsN0oW8amVTlZblFXFEJr9xkQWvR84Ys6vZIBvAqlHW6t3
9LDFQeO9qeBeLAs8juEMMMyskl/GRl4Df4NZd+r3clP/zKMJF8RgF5U5Ykcy
Fb7Mm9UZTIIjB4Gsft8XCc/3WVvag466tx1Nczp+CotbdBibH1i3z8yemTy7
sq4YN6QNrcCriFajPMhLa7LMl3vWcnbU0U1vsrPP9fEc0lXMGY3k5k6VAfLp
/JDjKqe/7o46T3dr6w5rG2/i4cCQQzF8+TzRyHet9TpD6p8pMrzmKdqd3FAB
E7Vaahm4QA/8G1WTKibCkJbaUpFEyhUe7HSLDBfjjyBnYbwIIIuncazgjaE6
YcKTWajVkpXHSKKnlV4gxLmBpPa+OjfZgGo2vCbg9IW2V22jyAe29RCEZqdx
GHtRdHNNnjznvpUdxvxmGA+I33j1chS/6J9qdlbZWZgTPdvofmCp0KIC8OyV
g8vQ4YNeflwdXFJ5sQYqu0GpO0GsM+ZS/7CY9QpHME54z7oA7imOu9OHOD6k
wuacNijpEZ+WKWDthulxFsnyG4bKtmdfPFWXE+YKltnlI/LWw2EkVevbgbKt
Rlh2ii4AXXQU8ccjSonknJZO+SRHK2kgAYgWpFXShXGeNdeklnccTVBEbEdQ
Nb8bXKSxdwWfDvjaKorVz+D/m1g+kflCUFxcCN7pNR5OvYB9z0CzG9yEQkTp
RsdLAjj/MZRZbjz9INSCAqf5TZcRHnDUcUs2htO6NTBR/6Zz9SDYdQ7oao1T
lnFjsrzJ2OO9KRSHfS46ZDJG/+7XkpHdD5wI6DGjeBFSMVpkq6JUghb9GuOq
QRGVWSbJIaVCpWghMwfS/C0iTwO/R+ZeXj69bYVDrm04UJhUZq/6e/p3QIw8
cJ4VnZVQrCjv/D/xAYiZi8cW9mydUqqVXCr0WXGjrXWz3N758kP/BqQtmgcN
g9xBFbwdDWVaYUdiyjmmPYJsiHM2DhQXcXFkYbU7HnB5F5xWXwDMxGr4z9NV
DLBpE4oSpXlHihn0wYghhnkqNJuCq70DO6/Gp4cX762tCzImbmbjLKAyFpmt
LW3QovyUkKRJrRskCJtqNEtkj50oQ6gBU7xwjkPnWyVgLqzUR35Cc+940AyK
qj/sC8U9xJilD0/dnkGICe4lAwfdlSb9aZD0MM6R3B/uaZ16wfc0BigCDBes
7S9gJe9YrQw0VutawE5qxFvsdC8dnBI2vlUZrs18kSrcn8l+lAOeM7qQYtsb
saGo1/N8+8jIbKoRYNu7oUNuO5NNzM5HC8bWAbWT9yIy7dTC0SPjNEHqsaJN
+v7XLC0hA42M3uxcpKjlQfb3/wnjMys8+iHjqNE2CNEg9Jdi4BJvK7l//puh
/2NanUMS5Fp8YthYujRv2XVEK0TeNkVZZMp+2WavyV8vIEDxLNbTcdj/m5gN
h4wxy4O7mUqkm3ozAlp5mDdpprbelmENwaE889tqBeecFNG/D2eyvJ4+MHGS
CytIEdx9o+cxP4VTVDt4e9Om/oHrMM+1+14++k/Bij1pA2wItFRFr7KyOL65
IAjB2VXhvAaNAkIIZF1btxPncMhc8grp+aizkfhBSEOpo2d6jns0T9wB3DJJ
5z3tSW3OEPZYkTVcB/o2RzoBrmsItnb3KPgUEVJKud1KHZty5omNp2xbRuBB
/05biR2K6NP2clqQJya/c1RbtdDhEjF8oL6cm5jMMhbl2o36e6kydBSt2GIf
i3qhc1RLF+fweqBQrtFOSMrg5TOQptT8oLNceoF6/sYvr7lVjLu1Otw2hc+O
lSWa9IFmEUjAGp9Kpgkh5YIP3yWmYS8ABgHTwNinoEcg/mCTCgyywZx+FCAK
JJCfWPbbUFnq5EJD2l2xx7n260KPemNUmBakzuRmo6tcl2hKueIUnfMcxxBs
IAXkdeyKCkeW3XYQgQCDATpdA2hhByUWrhRknniFJws7/k6Lg9mBYh5e14Xt
kJ1W5/7Kybf04HEwjnLquRLPojngRNVH2cwgEGN5UoRqHckb2FLjSfKU08GL
cyanPE96kC/l+/eVx0AZ8HdFQ4LafwTBCw7Ws1gDRISHKZLDm6Gme6xj0M9v
fsQY6Nn6eeC9CIf0iWOmry0dPPrGkaebBrD/hSyBpo/5fMklR3zyMT0g1z6H
ENDage6K9NS7fEsBzw8RHbjDNtYqczb1AhCmIgjR/krnX/o347QoTo+MPDOa
D7XJdJU8wUdWyOyDErG9Cu2hNQXwG50GEhipk6NSQ7fEKexYFQkQSpBjJJj/
W88qBkCoGH04aa+zw7AYZVT6BFvaosm71gPYaUXlT1jGEaokjIXUKXKVCUXv
JVZckK5uKKG3bHEbeNzr9Syy37ytvi6zG30HwTYubS6RM2H0Oh/KCUTFNc2m
hpsIrhyfQi/JNbuc2hi/k7MiXYKY/K0rP6q6OHwaU/Y4+wNYHkwlI3jAo2fz
JmPLZ0BNiWisCS7OtsymVH+a4B8sfdeCw/W/cy/XjQPqjAklVUsg4YV4izyu
r6jz+YSVBMlzxK6AZVveDMG1m4vRk4NSkQl6wXv23cWBqT42HoxowGSHrtEa
AboVhslvR7Qw/myxLP1ub3/oH3g0VhWEypqYnbfjCpYozgkprplUKBjUM2/X
9TkAdfrLvBrLeAFCfcUD+v5NyDe0VRyaMBuDt1Oqbu4wuuCTQh5DWp/c1Gw2
84+lDAzIfPaTBlK4S9cyxFKAlCIAXybeU0IB4y5KmxH1gsDqX6ua2N8InJ9P
V5EP6+e0+Qc75UHh6n7Op5VtODRPyX6a9ouiw5av6nSUBwUKW4YtSRwsKeEE
hKiI+5BFfxJHvitjgB+m7Vl8gZj4g2d2oKzwOae5Q1u0gpSCf0KsTlM9pLeF
IjyatFUx9iwGBCLHrLiduAki1XYMkzZ0chyHi5CQ5TimpMegtpzGEF0DJkCp
cktj0k+zbvwvpjFewj/FjaccmKxkdTo94ziRut4XzyBeoQH9mn1GzSDhbm/z
JtZpgIWx5IK9YtYwjTywKMGhMtfNDOKxk+MmyVk/hFaogDFuhhgJ8OMrhnK1
+a996k6Ogsy+4lfQfNApd7zvPdwJYzjGalF4j0VcXgI+qKHQ/4xx+GAeMqMr
SmEK9tSFkr9y6jphUM0eTYqBwbz05X+9kTWzfLcsD9tl39/M/XehB6pwrdo1
sGLD6kNX0QDaErq1ZF0hvkXtt0HAd400iamur96S2Bs2NURydwGcD+S2OMOW
ey5arGzsYeFx8eTwyWFcZMjAZU1yOTj/H8ilfGgDaf9KEx4w5+5+mGmfNRke
ib9q+rwI5yF/4hL5eo0zROGpGbI8Q74u6AeHXHPFzykaYXJEbjzGoTHfxOwy
V96h9ZlC8McUEe34V3qDTgCDabrzX0Xxz9Eczrcc2gLYt4EtC4zbEdNX9Eoo
myeX+zOKJZdY+d5PCVS9vc/4cQirgD6035w92XgB7nkh5EZo0IpwjR5PLA50
XJ7bS/IbO1KNUnB+TToY0znJZwO5kPEna1hYmZnwJDU29C0KtoKSGvmjQXUJ
xypxJ/lau89+dfYSWcoopRnN6eV2FLUKJJQfYtfCVd4Lg1MeQ9xyiBpnVNy0
FMfBe7aMAPO96gFeNScS+DJwPPL0NqCtxuEEDeGAfs9MgkEQlG7DQBrwNauh
10w5n7vk46fHamI65/sy3HpHdZ8kRF+rwRcatzU/uCBAxC6rb+zxLmsYa9Gn
/0M7dF9Rs6oQNlmf9ikdt9RCFq+SXP1AwC6xw+KT0rYbvSQfEh3Nq0fRw9LQ
KVufcqJrT+VP7KJr++ytIdKPOV0w9FECsZL8VnVqLpoUy0OsCZAw6eQ4cZEs
jLS+VPiGWBZ1L9umpR1DXg5JufjLDTKEZxZE7FOT8Awhh9zoA9605K2LRRkY
mtl97fkNOa/+cYmpl8VBg7m5vVPuO0SYh8RjpFpbKxZ8xk0IZKVNUIG2JCKf
2jDQgU6090Zn6wUwhC79mq2TIx5LCUwSiTXqMOwkksM8h7Dd3F0y22wHqJie
e7dgLJ3UGBrNKbISDVCrqAMDGcypob3Wi0DtDVGgoVE7tr23GnZjeTdBaQab
Qj9SFfCj5dySHfpyb8EkyiIuGUArtKZkreyMtpym2jPVmClf3lrROVLGootC
MkdSxfGi78fzdrs685YAUKAjaNtCsML91bbQB/hy2frp8xvBkCP9SKFrVJ4a
614BEYBSokCZBHjTCHbfbtEYaRINTh6n1onql16eBp26lZ5y47II2pUMIHpo
r09pMdK8gQGQS4dn6R0fEdUhf9KUm9UlOn9loiegX1tEl9yqBnXEoyrp204c
FGqMgJkRQu47GkBzuSBniNqg+9yt+17FIToV+nuJxzye4DP2qvUGX6b6DaVu
+X3yEBGLTEq2sRKlIBEEnhJz1FUFnUmeZvpxsfr41QpaYyLlU1o4qnDuZZ+U
XDKTC2INt+BksiU/1/PhyyC2EAdLmni2gCEmymvqex6EiE90XfIeEJ4jKReu
cGBQh3wRsLEptv7TNrzu4uR3z4KdMNo+hGgI3+6Ws/Nsw71kOB6me5ZcCWNr
f1g7GVPxzSiu42NlMus35TTST4mt04nAyanQ1AaSTIojTG1I/FBzkeksb7X8
VUxE699sIORDxa/ml5Xvb95vgDKqMfcH2uDB2JW5oBtdFITNvCbOMeKrq52S
o0/sSiTYG/uIlogyjV1MkNSvzmcfWMxkEEh1fts/NfH1HWWm2mEvTs8iL/Jj
34n3JhJ16vZgS+RS/2UkT4oz27MoUIf4j7ztDx8HA4AK0rYduip8dNeb8q15
QzpjJPoy7znzFnl6m8nmaJmtU4f66skC0GK8pmmto7BB1oOc6nx2XFxzHJ1A
mALsJPMv1FiAAo/7j833oJ7RZeeorOtYa8daCvS9v1y9KzBI9SaJRMGTU6gf
TIwj+natzUtcR+JvkmncOd8NtGDQsTzxRzlIH5VEfbKz6lv+xmkU6xRTR/ZZ
8X2nOKpMtS+qcLfNS3VxPMDFnRiIXkcmuwOCNXovL/r3Q4xvhn8Lu+K8g7UK
UE7oNZ4eqIzaD9q1ggWzbQmQYiD+rEtQJJccLjOILGwsrfSJXzxia3CxAaBB
sjcen6emLYMdEcBdENEdi5e4MD7oILxr9Vmx8XlQE8Tb0HlfzWJLLoVswhfR
wSB6HhY5Iw9IcHEz77LyM0vpNFgh6o+7EQOkZjYbyqhye5HHrs19cRM8Arml
HHJSjTivDzBK+yvcxxnV8QI+lnpXQiIrSOOVR8D2mj+AOPz8izyBzkPuoQxI
DEobM4/tFYEBpzik3VAofk3x8mvjNQ/UHlQnKTeISH3VY3onDS7Gid/hLtEY
KMYn1kfV129pJ+/sQQY7aDjXmf5wQR7NnrAKHqUdgiriKME95MGazrU7f7xQ
gi1bsHUIGO3jrQ79cU7bTWvv5QkFYleTqVIH+Biy+nLT7GR6TbwzzsDi/JhN
dacHjQmGAh/QIlTQRZfvmcYGzinNgdYkkYyBvzsegeVz+IX55RlsfBu7LwmA
6MLBLstGxA6yig4EhuZLeLbiz0kPs40gG4k/YkHKvCeUDztnx8wnMzDVMtb/
BfcGJ864kYtL4cNqr7dM+SaTHxnFaagpkcrvs6ck/nuNnqePflQMHGUPDEl4
yKV8AXzC1lD1bxdfVnorkuVGF4QRqAjJ2sl1FX/wrvQmOwqT8D3SoKr6sdY0
o0z5BV7qKQbzePb1ySlSG0DfntYUQCfkrAhBIPjWeOqemy3aDurFQSPlzanh
41foGguHwsc4B38slVoMd3oaXLlIj0U4ATm1KcS2uv20KGv5RDLvfktTw+cT
W1bSLzgRWi/XKVHeswWPsASkSYc48EdS3hUipXkxHbjIWc3EfHXTMEyHUF01
zDHeqK/S/wzwvnU6nND6we97dgfUUlUsXCsA0Ym4SQ+PFE3ZFcLmtr3lgmUi
9pZxyIjAm5mTpJPWp91E7x7mV5TeltuPu7PsegjsmW36qz0v3Yt7giXOxq7D
e3PJ7GLwcHRRVkbfnB587j7Di8j3YuOWoStpFlqq9YM6gNLCQ2KXymJzo+Zi
BRgKn1/Dgy2VipVeBfaqSgaCVIPCajMm2MHjDazO/b9X9OMoFh2yKNP8GEpp
uFPnjSaatqAY2DFaWnt0zFRylXZlBG/TYWgukp59TJsz2exMbeNaHapcGWzT
hD4R7ohhMDPj4iCivQn4rnddHm00JwjrU1IJP5yTkduCQshtzx1SijuYCb9S
vZV0WbCwy7CYxGmQ32+vVnCPJSOIgMWhCJjJ0zcrt0sXtBDi1P768u2/5ywz
q3NWBKjumldlBS349t5QYcOdpPR4XXpRhy/b81uzi44qsNf9aAUd13cXw35W
9DaEgkFnFoKX99m/imL1MkCP4b1z6h4ZtUtl5Qj616yaxIuaLA7+Mlo7JTWk
sa5HYnzuIgZ+OfRHAikPudEdDGWIQ7DSMnCefoB8AtPO8Q2lRQPzXvepbwSu
11lJQLSoa69WSLI/aPRZiw8N2MjtvvcrfhgB4ykwlA5TrW3Qom6eHS1d1hH7
+2JKbnG5QhldCdtX2ZRqKPhaoghnQ+ByvEmqeUZnJigen/ozzPHQ2TYDJ2iA
4LbaauuCPI+yxz7lmIUCd4+YedhHljYSQm0r0k0wedyXPiuQSUYwrCPK68hW
OPN9/IR9j1ib9gCyn5/8+xpIwDqgH9fdb69odIkaZgQFdrPTp2cMV6+YEY6E
L35NnzzTinsjOBTqhJS7qvTjYzLErevGXihIpfNFLxB4smkD8fwzLmgSgSKr
b5pwDiOfI/BS7mleyexopfsEwJd7GM3zBuZvg3jbS10NSOOWnhyjtQZLY6Yq
0y6iqsFO08lwqYnxsbzkCIB6dYarRW6mtBOyy58VrQh6TsWdr6kXxDOIhqt1
HOnTyhBJqdvoamCnY4thNp4m43chzShOu2zSJ28JQChtPKwA053O+JFP1Fgs
Yjbslbd5tDdwgSw4dii6Ts+rV4FW0Qbl77ubrL5PbXAUNMd4LylcwpTSCr0H
Gz2GCFGvqLz3w7mk37VVlbRstXDIC96qTAWTLYAKvG6seeW/rJ98e9XP6AlQ
L4o4xK74+7MrUz3Uh7mWrrXYYw1VfG5tU+Fo2TdHIy4SckIVaVS3R+ddrlXO
jsbdjKe7AzLEncLRz1xlxPzfW2tqsQrnt2G4HpWkvQ7ka4xmnAGTcZ1rmVMQ
JcBpE68ELbeBRQINMeaHPQqxCyjqcsAoIUiPJs5onjq6Z/tDobQSP/Y/mRGS
0oK21bWfuPA9XpCNDIGwTAxbjKhGlnUha912IpPcykSrwXElm2URB6Lp5lUn
AATNZZoYiCaCqM3Xp80AzqsElbLd8iRrTes36CunlJ/qmL4qphH2QrDWljic
UlN7/AQywjgGQgfYtLqUPJfIRRyI6F0FjaPjis+rB62x6V1c7lkHYmjn84ws
7W0ivCc/x5q1qpUnUjFm+T73UBKa/ehJwhMnCkZh9u3yVwoxIMm2T5Rp9LcQ
7jvm3Lqk9LHbGgA3RK6UAxUAdef7AXIyu/ouPri3YIcPbyuFFO5crDDtdEUP
8Qsqn9fTkvmYH3UAOJC9dKgbqJboLRZAxwWJKdkXz6OadiXgRAZXKjQkOnBo
vW3nEd2Z4djRFUMSV+s48KfjJHZ3umZJvraZhhkUGtip6/3kkawl9JC2auqR
aM0YJAAUc3aaWmFiAViSm+uuPkaCBNvqSL3CbFUYiiKoSOD4DnDP2C2N8yc3
OVeBMz4R7Q9UMWsWeXoQwHel+wGVQ8MW1Vm61Dk0rq3NuyfZJhYrTY24S1BA
KEr9zzbS8pKah4wenAyLbgRjc5Km+GYKtqHlVwKUU2lsETLlVFO6oDvoBxE3
iUBvGRKmzFFy6JqRtvvtmFPK7fzQTkfSINDWeeOKd9M/6QCwhxlmakKSKQgt
AleN2xktJdpX1RD8yNqeq0ci2OYXVwuXovO0nhOpatFl2pTtaiy6sTDY1MCb
r5irfCjgSjLvckBoMoPSgGQ6+fsTbs5xSwDbaXaLa22NAlgWSE5sbHkMX/MX
nLI+y7jFK9KNykOIUY2XfaCaB3ApXohrvh/+a7M7SsfqkV3uredtX4zgNab2
KbNPP0CJnnuUfGtmewxgnipV0HCCKQsNXud0UjlIEhUPR70okMjPWmd6Wwrs
wZoAfCaYRnXQKKpVcipHn3Qhz7HT540SvE0EwjzfdYr+oCw7sNJHpvzaieRs
mrAvN6CJ1NaK+wYa8VyPb2h0I+QGGGlw61BAULqa3KRUurZn+HkcUbzKfUqj
NdETuBdfKQR7Mv5MU9xigldmC8Apz52/RPtMhGdOfbu1M/v1pl5g7uKTpdiq
5pjv80PTagPxxHGnSE/zCv0VZYfGDUx2OqmlrdW7Otr+9PnWki1Cxroyso4R
UxsdmsmXaACZBBuzXwNXVSJypoBinwYqFB77xhLymTeECqMGKt1Mjp/tjFNo
zasdlff416BD7J2AJkrnvSKtjOflpmjR8VJL871aHIKebC+FMKUZz5tpNj2+
5qi+AyIuUhpg6fS6/7zWCgA3zKYaMk3yN+/PfUc66YKdo1t3poWvzoMwOOJp
GxWo3Arz0f47QDfEFUTA6i6MYuCoiVfvvxvODeORy9nE1hcp+F+wGt3u2P21
Cq/P3ObKhqcDm1YK2DPVw4pb3UID38PGXSdqVBTY0ijML1XdxlaK15aMiQ8i
1ylHA5lYwuReyUewVd2Ugomu9115ToR3OC4am2KijWb6R1Uh5qOmFBEP6dtM
mp4SEK3uwlApcw3RFYjy4hgUaPJ2JnNGlJlNu5ytSKvsv3E8PSQSl99ZQMRi
voNfHXS6nQzXi6wvkAY1gfi43cA8nxYVrGu4+V7362v5BPHPM4YjR60hagWJ
L3GG0ILIqPz4q4PGb3va9hu4fE/KvYoi2+jfmsxJ6nimIbsKHCuKOpQRHi1y
+r6pEIAnmsKU1uGEs/vYiaNFEK2F2CPC17Y2AcnbbJND+jUIvVd8Hh8oSvPB
Wr2XsTKWIWbkbUI7Ew2I0HIUVpVeC5txyySdpcNi6YvUd10wyykpHGTBUx4L
jvJXH4PM7faG0F7RRq9mQAvgho/a2oen5KJAIGDCE8F+5F8KHy8uwn8ued6b
BoGMVuQxcI8nP5BQLn0i8bzuhxvFFPCFLoUnhzm2du4M6iCM0YaZkNGrMyZd
+AmbYVZe9VnKwQeiogx0vHvd3gISt0HdxgAniLlVri5QCuwNb/18Di4PUEoL
r/PbV/qtSOWPs3j9mrCV8J5UiWYc6C5WNLV2KMipej5OhnZrtlJk4wI0y/AL
LqEBZV6NtvuJY4b+7wJcJWxlZfue1RKUbGHVgBcNWztsuVQOBIfMOjSCeUWx
R45guZuDBaVo5p+ZJbhEgASUuSXNZDyOkMJb/q5dk4TexD/fldsjFoPTxoUw
/Z+3dzDFuzPhJFy6azHq2YWhxgs4p2WA1Y0UoCQ6yVKvZUGY8WSKiL/m2DiN
MaQu4B1UHQUUN+bwxuQXQ2zz0jJRautxwHQEfVGQRsy0bog/+kwoZSLaMlEY
k2eg7Nd7LikW6H/8rDFiSRKoewT3bY5StWHHoZF5YBiGQ8MIeg/mqm3Ja3BB
5+8Q6Ofvgai23OUpdEEDDQIdwnO/XRSrQ7+fw7D4tWBg4nGXC1VC2Ks+oK6i
EaOdR9N7zHmsoISXFzc2kmuZ/f0Vgvc9KXY53J4LPYFqzth8JOtK7Ihz+C2J
YN/cUlZZIifxpxmOCncWXs7V2ZC8vPodlKgx1SHADenxys7IplNBGYpnDqOO
qA1n95vRLC1NmhdMK/bJ+9Vktj6HPXpvgMAXuQrxJlXTY97Ze91Wf72zsQLx
AbATHtZYPBzuZQ8gvsL1zLChCSejXfGxQDCV5hSGRBrQsevOBBtHXC+ElF8y
GAgv3krxiBAdaZlXjdguCz+GSaqtz+16mhzTQHNHnicCRoLPi2VvGtmtY+/n
rdM/bYCW29wuiTDBuaThPMxha+xu4nUvZh0YpmyLkwiKdnsAWyWY8bXWDmFJ
Z4pprEc85/JqaYuxLQEmZyXRKUTvvedZWq/NLDMVgRAuOACgGNf2f/ok1Z19
cZFJg674SlFcuKN9QApHozssb+3w10vHxus8dE9NP6ubicVf9BGd1DhNws8O
5fKnUqGszFL+Bez1L4Ye9lvrfE4/7k1FqFGo2GG6WOqCtWsVUbjpQU0ovn3j
/5Ae3ROeX/Lo9sGIkyniijCp8Lnkhp2zGLG3PDPGCdG7+VfeHZ3o6IrIcMwj
/CWTl7RAXVVcDPD/wk8/tDT3wZ/h6tt7U3xhT7DQJgPqQJNyhKq9gkWnw/Nq
ariHXQ3DN3YwnRPvE6cHFhx20B8s/O0UCypjSBMDv5CUUYPSIGmExShyGxse
0fkZq4ZiGVwLTFZzqIE+Os5XerZGAX+HyA2qsYi772XQeHsjnsbRmp+TMczF
MH80zGSOQS5qxMFqXefcGK+wvrGqhGZuumKIkGiGbNF1DPfyfYFuPKMBVl2Z
qHVvL2Z+x/bi2GYG5pQhP5twn2e5wS0uYXpfM3u0iQs7BPvSqDsSxSNVb3x6
dCm5yNidm2iHw49J5O180JNJS1lAsSmKIVpYO/zXp/URm+f6m0UxLt+CpLm2
yiUTFYJP2IH3tFjroOBxAz6KYBbocinCZXJsuzNpwYYVwI1V8xSgCxqJ7ERF
+R1jvf3/IVeALlGX53S1Ur+MkCOt60iAQMQikz02e0VKs4MbJLTtOqpNfmYj
ZwSCg2gQQrFF9PzZZ1NxS0CmD6fir8GEz6ethoxcm2SrFPoU8hVNf34bVV4M
QWQl1BB78T64c2OgOqlIwtAoL3MhN/ppyYRdo5LI2XQ+3dHJZSVtPwA+JIDi
TyW8fQ9ezi7zRmdQ+iu1pC5td7EO0y5tqSs0ck6QYr54kUXfxU8sEs/U3k7D
7rZh8rnQQWHR/f5kjOsa75XYl1I/ZM77tCRcE3E9g9NljAzcfvxMWs6XXU8m
mxEhvq+j5Ca+GZ3JKiSnmYLC2iEeexZuOlVqbFkxiU3n9oORmOfiomMK3NUC
dhXiQDedRg4ML6lzf/rDP4xgKGXsJBd9IDk/qus4oDwfXjaUtt1ckIcESPOF
paC0V9R5JvpbDdw7TcEQhwHjQj7xolcfOq5sJxu4ivCBJwNqTVOvFM5YWFuP
Dg7aVMs6o4EKA8cJwNo5ls4J9QO6vCyTEEMIpLudb9IYwKfnc84kVP6SB9RX
fdPtHxjPc/tr1257T/JrvdB0iw5c/7ZUMoGIy+EUGiNxduCyUzVlXZMW5zZJ
MUrQRqF30yndmK/jjr5GP8FV3Pon8GZvkjhmVqAUgEYHBEf4RxZ2whAUEZT2
/ElJ2PpyhwlaRi9MkxWvuMql3oMnFdWXjPc99xVfdKax3729Qmpzc1udGTHX
i/6uFY5YgiWVt5gYJu3B+FsanN+Ns2HyMBWUzq8dZFa0kwO60fEQlcggIQVl
6VQGYsNbEcuochyO2R7//O7RGn4EHX/gq998+yxjFAhZt7VIMy8Vn1Fkl+3p
ikARcKfvCsoleSYTawdzIaPyAtfepd83AUcEArOJAI5pGduc5ezwmPsApJGH
fD8WhcVYOIs1i8tiU4XdhxgkPA6TMHkYaODHmMO0ftP9ViRs392OYJeFVQ4+
W0jtE4wewlVQKMXXeurQX0r2SsUDZQqiF3T1f7LqoCL0KxyTyPr0zEHZgXQw
klov1iEmsMHbWxZ25Kp6XXdnQdz6OnFrSIofyyGn6uLZF311fZZD7W7z9T79
PIeUC/r5vn8j1gWoB5ZwNIu2vD07z0CroLEyC9CGu+ejBte0kbs736WvFPHt
LN0coI30/iqv7+q+F1AOpV4dSPEBOjC8H4EikH0fCqt1KM3Ci56Y2AFuVk8g
afu6cW43d8cwJw2ZTSBU0TuMAthEdNBVv+06jW5hIcgW4BU+OG0EkSXGvGwk
UoY1omcFKZkyq9tbXuEGf7GD904jdWV5DpoojAYBbho2gkvAJXqWkW0k3QrX
vGU8fEaY6SvV4etK+6XLo+7JDGQPECXUiCo8Ip8elhDoRlXRAImdFtoJQ47q
InDGG3qLrLYCXeiWj81GLErVXxHPGYtf5fxkPU54lIkhHl3K38GXj7tspQtQ
b8rAksCxaYF+ua75qKXwavse+eVhLyav2foYYD48i1Y92pSYX6YJOGYTnT8l
pRDaoyn4GOq+BnujyBKXwkTmUfYQoxbmAHhxb+0iNeeXDEtUtMhbilktTAgK
ZFPWy5b6yMwbAR4okndpUdWxfEElXoQI0rAaBpMzMj3auBMWeXTAQIrYG1tT
NWRwix9LXPvWGT3sviQW3wqEjxGU7tsdcRWD21TUev65X8/rwEEmKRw4Jlmy
FN3BSOCXB8731f/rvXcYgqT8HgAW4uc7s0V2z/HXBDETcACBpQoHBHcoa48M
ksb8SMj9/uUtvX+6usIDCaIZ5r+V3RKley6D9Sz+LL9VHa9LcqeL/sO+HT4A
bR7rGZjkxqHrxyodgC2xGcgIQcZUPw7hXqC9pWSAmS0+vXgUBc3l++b5AjZs
6BicROr/GNihgHL53Ozk3fMRt3/cG0I7tgSUklurr6xyDKtoLo8h+0wwcOtr
UDCpz2ho8W3DFPCphqC1UHLxkVpK8T3xM8Tvmzu6gN4sLlQ3/2KO6WI1ur7H
u0RCvPOLhz99d8LwNR2KQxMur5yOEaK6PuOqAT6l+rJKpdw+2djX1BVTU2iy
UNE+EPDVWWUOJUBT3/rDZ4ErnjEt91v7zVHBi6wCAhuAHt0nQRr+USpdLDYM
ATiR4jyEvqSgDs7wcOzReMLywvnGtcvlgQ==

`pragma protect end_protected
