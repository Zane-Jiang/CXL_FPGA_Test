// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
K75fhqwT6+KBuONLqM8suPyMGu5OU1VfN/qyhCR2VhyISwzvkE5TdsQqNmq8GPfe
TG8ol4d7LN1ex3vesXYULr4dOBeBYBNbifLqNYPVRtAZ/bzhpnluiBx1ztuO4Bdj
+LN4MhpUbKbquTsZdtyJ4dz5oeqI3Zlh2d2o51wgmSGsbELr5MFRMg==
//pragma protect end_key_block
//pragma protect digest_block
tHx58+uoeIost12i1dEN39HL7k0=
//pragma protect end_digest_block
//pragma protect data_block
0Y4IPMCopk6EMPMq7jE7g3Abxo8vfmsVL8KVNN2116vxwdJW/LvtT3mnJoiherJR
Lam5+m8FJlXs5AqhG8DA9SqRHGJO106zzn314KkU4cTDn07/eXdv9CBhQ5IaVWdp
ET4HH3BBQdmTOHaDDIJRxPkXar3JTKz4648GF5neLaJOF1vuqqQq5zgZFzkP7A/3
BMHmlYzpvOIURmPVkwRnzpSPE0nkQwsm6sStHPXrumXjk/IsEUAfyxE8Aae71jUG
SENooGpqEsi3QjIaU0HDg5pAvZWWL5XDlanSdsTGhVmy0IHH9eUo1aBXa67QjIYG
sy6cGqpXzsAKBh3CyV+8z/Q7CAIzGt/eJ6CIxcnEt+Bnc13lskuUjroezcw6GTFx
unualMeMiZYgQl6unZPrabG4iCMz0e/46NYCXKYt/9lIU36OJTk/urec9FkReFE4
RGmpwg2Gn1yiicvegZFHXMzloBtDZK5PESIOZmvky0RCCbPKrL3jNttoXIKAI84s
CvIXeVwhi6ez3Q2Dl2FMT+mJAvu2mfULdZ/IQjcOh+vZx65ZsOmXN+nelpWITZ99
LrbC/hUW6Dpcp9sZD3dmjGPs3wx9w501N6j30Q+4YQskR95y3iOWankcHXEiwthP
2TH5aHCT9szBhlPFWypbFzkX5MPad4IKwwQnxWfhc9CSY6jzPqFUGhRWYmb0YgV2
LMpgE3AFtIPWyWygI2Ft67cz53sIJNeh+NBvXAs3L6D5oVshroYhfTZdeGY3ZtIe
CO7k5RL5SfwOiAC4A5e/0Wgkyn0PgD4R4r9op9u7jkpiOKiBlWyo29KVP2YGg5S8
yMETebYGRa8hc79m3XbO5vmfeHsyGLltAHWOZ4PizhZSFTR6zBLAYlrJEDjGoEK2
r5GTMa5K03B/KGFidCSXb9gpbsK6ixsmQAI2PFIUA6SEhhjPpYe3PVx9qoNGvvj5
cd4ZJcstDCKLqOIkgOJRPco4MXNV6bNHxxJBZiT4g1EkfipUBbqDpomHsC7hYQXg
0kxHQ+mUV6XqJPQA9OjxAxpi639lUaMkL9lTMRv9v4qLSt4l6GdyVBfEhIIvHHqN
Hdo9DLJfk/8tR+sszWubwiZ3s+TotU7I1af30uyVA0mBzPTGTBUyxShUt8WEUSqZ
LcVBFLJ2eSLFlf4LqgPuu0bCrdSfvGzF+oSjm8UpyUqqZZM6T9smQwIhzxTXE6UL
ck1ErdG2cbloYPO3uiuL7lTZLJRxYKiZdtfdaP2MzCv0MMF0gCwHv4/GkpyfJhAq
q6xCWhnFl0P5SW9eJ//SGjFVNv0RK7N0A3duNt2urImNhggYXGSvovxz7nGwGdLF
0O6vbCL9ZDDEk1SrpgySBGv+hxgyrGx9Z33M0X4TCsWBWIHAnTWiJI+kieoITarW
1tVvP1vO7WlG0e1WNpuyQZTd2ra5IgFqiyWgQXqqF39DIlj0fJ9IkbXp7hPNlZUy
+B2F6oxdZ/Be/dSkPq+7eTk1zV2SQuu2pP05gWtfAGatbhkIkPDvlmfvmFi5BOGn
+JmJ65Wg95cF//wZMQi5AL77zwsuFqM4Xlw2jhaqEm2PTDYCzmgfNlBrIJHFCNUR
5qpjPKVtBhWzlAKRJa/bhCxdaMTcYXg3D7Rbi80t43Nos9lPTDyI0Fyimts9/LJ1
XoKAvaO1a9Kn5w7g4/ASHsp/lAg8SjUKqzG0enAsisJpfGq2Pcqi5ItcjEHnOVbe
yOf/ZhFrW8mIqPlPdWs3lEQUMFNPqpZ1++rl0tc4Af+Ft1feltQXMhSGteWujXLr
dagfJwQFBjgoVHNfR+FtFWhV5e6IuJMNEJiT8cbBEIY8ncso042WT/VKQ/w3pEkR
CEz/+f5Ka2dTX0VpYImBT3oVKHAMQOXajRNKzW4Nl/ql8/aIyZe6uTk7lkTzV8+r
K6MwJABoEZNN74A4eONyTnBnJdlTAI4OPyeb2BmVM5aISVGkCKY3zM+wGFjb3ScZ
XmdaQvCa2pMzeS524KUQVUI2TXrrNwc8lx0AD8cHshZvBEBxHFCY+oXJ2YuIBSpw
lXEl1YF+sCW+z1oMUkQ9Nee/xNtvpMsC0ODCxQ/NIdkztzK2m/BJAzk9UUht18oW
Xg2ZhScWLMnmMM4ba3Y1SqiiVsGjrrvVma5LsNxqXWly4BwSwhHHWt7lsoxCND0z
Pm7qAX+5ur+ETQV15rbjKC4vCiv1FedcTroRkjlau98Vz51TG/wYW6cHTNo9VSEs
lnMvHaPdblNWTrcmO+LB8pU/a6PjSHZ+xgyPEIVhKZ7YTGxFXtFixxc1I6tEXV0x
8G6A8QOF3zgUjtaRo3h5XdqqNaNjtarwZPv8ZCX+Abkxv/i9JjRd6muw8HBqk6ao
dGxU9xb3je6UPbNrJJsp/8PRmRMv2ppqOeqz6vXceQCvAxpXRon86mnP01S0/MSk
EFmXt3Cl5mcrUsRUSznhLTwSOjNz2V4iOCLP2cuVhswHptbYoteVw3WLtOy+gkaN
GO/HVuIC/50djY0WkYj6oaqdsFnZ3Eem9FUq/xFVsBs/xtH16TyFtfqFwp+p5Ok4
RI3S+6KOrQSfnybbSZ29/rdjOYWJ1GD/crB83DhGAzmhjX5NcQ8+XiD3xLYy4eGo
kq0DL2QiPiAB/SZBpByqZUgViHPYieS3nLFOd/NeIlXn4DJR8yzlWLszutp5obg+
MCES6MgUS4EwZ3+E+AtIBlY11Goc4GmSIaUEm4WPGOrCDCAzGKF5xKEfKZjrM4kP
PmNVfiO5+CKtHGXzoUOZt8DLuRxmG4Gya3LDfDD0p8eUO+suc65Pgsrv+MipOzw/
z7EinsSZ1T/uH69Ns6YOBohTHdIS+YLKg24Z7t6l3MbhORFNssMPOPEhfB9o6EBg
9Dda7LPzilfYHFuoDk3vKLVe+RNB0O2onRT6sk9HHsbgzpnMqpOs/12llVtfyoTD
h2aw0yAOwkQXrczxl/Zg7bN1b4dDEooXwcAEY38XGQ0jEVM5/KkyTxzxcZMGO/eg
FiHU7zkkVGCdRghyqHdFWF2prAIvopS34S4ukfXUTJvD2tZehbrMkM1SOAaPlyPf
fgoZTGzVzEFQT1CAdunpG4utvhVw9XgmDPAIVFoVVrgbw7YJUYlGl/0NctJIhoLU
96oj1O7CP7RrOnGIJQuDRWHWnoG/Fe1Z+Bw0+AiXI9coQmiyFreUr79cBrSHwIG5
sX+K2fLq1RcSgUqTclK1YMYgfN8ycX1+Lp8sdLSzGuCyeKvJbMAAM1sqN3v8tPqs
4K7BfRIhdPgRwf9IHFce8pNXKOxxXc8z5g8f7rdNq3z0fZtOCtEUZmjAzyn/dW5c
i/r0845Y7udfNcIQrNQvp9v5cKE4Gjj8QL4JkZ+JXUwLN8T70K3NiJEI58fczyW+
1jiPeo1bPIDQebv7ZLPPN7HtcnFUIayOTy2eQVYC02E4Cr0n78gyOOyZjtsNcFLi
iEDG95rXl6QN1tTdzTznbqwCoENZMZ/LXkCkKG9jwUpObKnRGJyMDJ5HKnZny8sE
Rb0uEKxvhhKs4QTedzKe74B1uS6mWvKFZG5vDryFBXEODVI1OCk6oQL6RW5MmiRb
brDv8j3IcjWp58A/c9SuVdwxl9MVnPk0kacHQISxgllCTRFjoxucsDngCekjmOan
3e6qx6/vffCxVv1I07989zief1dJUGpExGZjRhVNWwnN7RP3yGsyV6a3fA3K8YOl
XUQ0ZFh6ilJ5nPmfNNhZcxB4dSAINpmV0gYr81cYa5AKw5KiLf0ejDeFtuFyxOPJ
fHzbCnl29q4B38PEO7esikNo4UW0cg2J7a/aZ7IViCddS3a0WTI9JDFnQe7Pdmmp
o9upLigHpvGrTn5j09sDcPhBKx8bs3Ps12IGl98CpfkX31CdmBjY8RaeerV/7RD6
9yxfLUG0XOknM55+CeVASY0Ets13ErcV8GP7TUF3JMd2Gf5knqJ22fEm25SMbRTp
vTwS6anl0TH9wIxk9/CrWAJux4Wd6uUxSiHfpaGa4RYsZiBrU58JmF1E1nTRRiVx
I4+E+rP19KtoTI6An1NCa7viI5La1TFjakhfGiSx7i6QK8kHihjGbSrqLim6oQCR
jGYbEaGH++MenwJOvE8E6WCrCuciW3Jni1zQYLAToOUB/qTupIRrAHxBdcF1g28d
RR0xbqMS8HSlSW7k9r/L8JzbrjSyfvCIn5/bYXQUJeIAvNSR6r7XP5lUXfkpnWTU
qwTl0SNkZeL+x3j2/z+3ZftKwnwhIOMxD7cOxtu8SsNjvQnRMXxa9Uq6vuvcMohm
fc/FIhG2EkmW8rmflHRqg4aajBQDjcXZh576/7FEtCxkHwNWwrLqGhYP9KkSk9sa
Dd3yyW0s1IbYRe/0jV+G9WeCO0L9/7B+M+MldGUUh+AJqTC74YisP5aqCkjbPa0O
i2NvVNueekKC6JRt8DpRtELer0TDIBVTD/nju6qJDsQFIp+n4FoNu/JM0qujeCPe
HTTa+eBDvOtVPxHutThxvonNQO1N/4dliSrVkAss51Jv7nDy6FaXQWrDnJhtZhBA
0vtUxhH+UhcOxtdr4MjHAaLsfoE6SWAd7W99+cTHCRmVQMcO20xT55GpkFjMRqYd
Hph9R3IazsmOuH58k+eVwwRpTvDAzB7hs023QQw2sSurDdPWyh4cEir0K0eiQ4dh
BEL0yw/xL8OvkY96fYto2onsaptAmZfF2+4pb9vfbGmOD4lbTKmagkLDvEwHZdSE
Lxox24Ir8GsHsD+ciT8D/4stK/nZUfHpsVLF3FhcXhNbsoeLQVlz6+Bsb2WFvCvX
8FJ8PwffEHqfunB0BGj0hCD4NRNxoQZSCafCy9rCAHF6wY7HkvAo5+BvgzvkNqOt
kxIRgt5olZP1ZF76cSi+5dsPKEexRTyR1ghBLxR7+eLzwh5en9YWMrApOEbIuPq2
xYAN8St+pZBSZE6s43jyjXtm1xgSAl/iOHVARX/DX9mJhVq+hxAFI8WM3D/U+QEr
S6S9+haXvgkQh8KTO16D9jgij9qEPZsL7MZGEK4hfAdp46dGv6XQrjdsFg+7As2b
1RxH8By9Vjr9mZSy5yp1tTskCJ86PUXPqhL8WdfvZO/nX/C7ka2PkYTLTn21GxRb
TWP3g8kdS81iwIsIET1XH1t52v3mcEBqPTppnVk48+ut9XI6Xf1aX6OL6pDJh7Hd
i7caKZTG7mIN4uxNTdZGgXTjUG8k1OOW4+Oa9BjTe+ffnCIphFDlFBwYf6wrJzb/
OF+IefZIoZM4N52RtGaSXhKkzDnpDaDtEecwwjiWDOEU6llX7LzdOytFHwFo90GO
YUXQ0IaHI2DnejfY8jmwnua18Wi/d9q3zIXvG7LCK/AWAE3Q82kGOjgk9OLAfKs8
Gw1aKHfGDcKL2/hPBQqDqvfH2MCe5oP+qJOFfhleHuTkUsqsY1FzB4Y0A7WN6Wzu
9Dihspw/fNm/OCFwlXat/4qCvxFJ8zFI/sx6fZPLO7XM0It2V3zB0zOX5IgpyYtx
N4k6FPCWjOtMopovYvQLbN4d1VU17LM4YyI00qEKO/ZMO4Nkf7WrWofULi0P3loW
tJWnTdABik31rtd5t0HCXPQy/+Z9DdrqMTFE3lapVDxGiQqC9I6QTapPh2SwnL1q
Wb9D1ZAWr2aV/2C8tKQ+lXRREqaa26W5QxAEaL7XCD3zHmq2DFch0nwt2x2chT8k
yd16Fa9wgyQloCRZ0/4Qde6kSAQ5GfouI5UYSS2Vd/5io261oX+4hKa4tP3VGeu8
WkR/St9u7AUg4Q5oHzcUiaGHwOwrPTIlwgOx5rsQxmZRkyZUN4elFyY29j/X34+T
ReA3LROncJKQFv1ngqvO2zGPcSPrQ4gyBauxv9JW0j0WUE6RhUanU5b5h5w1MLGZ
0bbkQE1mzI+lDkNiOS3w2jLOUD3TOObT/1MnAaFtLI/TRjs1EBfkdYnACq8WLnVT
Sr6hJ+AeHnqolQj3eL+mT4hnb7apVICp3PmqbcwlChvAGruHg47VoY7vXDIXseAp
FU2lcew3rZaAlFp9oY3w5NcIunsOIr7j6/ebYpIDK6I3w9GawFh00vYiwD4Jqae8
WYKhk6VtIS1EcAhjsuzz9tEOb+NcQR9ebZl4Nhyb/f+4s0lfZRsKedfTp5TqEWT7
ckk6iR9i7uSppNYmmDfGF+IQBFrbYJYmIyIiWMq+61D77P+6adq3qy+hSge0dSpJ
/kMOwSOlOhuAueF7yn4sbHhOmjEdDDKRnU3mCsIToZlP2gZlZGYT8v8TAdKm4Fp2
BINZ2XckUl98JNNRbwLZi0knnRod8zVgkaNS/8OuiTg0B4VlIx7+25V+tQfO0ehX
l9mBzy8AOPuHiXQkAwArhtpbX3lJo+aPag89qCdfLiwQ6vlvb1XtVSn4OVxRnTj+
SFEE8Y2acgMTBvvSlcZWFCRm9P80hnpo+MMcOpi4D9jWNKOlOMq7N361VZK+P51F
dcmGFcjszf2ib6ua4UGcMVmKr/3ZSYF1SNpyW0S93FAr0mKRDzYDrvjTHc00YiWi
bthY4Xnvi53I0ERIWlZ9sAIzWTV8CrDmdVNqCtCE3122Lx5ceZr4ThWQaP+1pRDa
hncJg/jEmVWjfgSmEGeOTuO10aEuboyzCi4NI/AxsN8kJtygaBxp8xzmccMLR15U
XfOYvzK1bPfGBLCNHa5zitb+2KToyd76HYRIo1GRctkSzL7ciOzIzJZLDBfQsnzP
KQqchWc7oKNtpDgRIvkHggXlAXnpzEF4OfPT7QhvMuZQCufFpDUNFmgcwrB4ihlo
QvQ/XgbtK1ayJV1tqcKCTnHsTkrC8RcGI4cER31pvd4nSV+3/0iNSJdizd+9zOc2
LZTzIAgPknd3ZxvktK2SVX8Zk7Vr+84X07AbjQMxDuHqDDjVc6GGO8VVRwsZv9ra
njPI7+0b2LLi8lCZ9xQJqMIjwC+F440A2nmGGrM/51l1w/85Q7P67w5LmiDINA31
qrCG2z2W/Tfau00yjm74KvfjOpAqgtpC2oYfgRMahjbjfWV14EFT5Zqvh2e2f0ec
0kfoH1Jz3VqRxo8fwK+SFg42kziop5y/diPcOkeY//OyckQln76rew9dQKuNsR73
DuDFmlBngAcmCCXJPycBKvYH9Qhr22caTVDeDHsDDY3icAPmX8jQ4nqYQqypApxq
TEW6h+RryXoBM2FQwFzFozzqfmX/W7+prUEI4PvTai1dTtP5Brxxcd7SGzpcidto
NHglG5BrYXDY6irVwlfQCmueLWNopnj/ue6N/AOo0IY4/0ESfGf1AQarUjrzo3F/
tEiMjBibjtgSOnePqdLKpFD49sxHL8xi5g03IFOz5dg/voiTCH0lytM3HZIAoeyr
J817ytlNvA1MJ7cJ2Udh8JriHs0HzNz05br7GRDfJFgR0ZU04ZiTGGi9wOiUBqeP
gNb/FfDnFrAeiZ3+YEr0HtceIjVqeAS1T3MLwuOqarMo7rQL8GVogPnoN5sK5jiQ
gY2PSwCNu4QzcuGd9sxhIKOr/ONp2QMcJ7/RHa7qgwk35+ilAe6M9kzpojoLNN1Q
bxep8srhJDfrM1jJ/1PjtEwemnKg5hQNxlKU4RO9IoQ0Sf+svjlpjn7iqyG6LLWL
6/Zvw1Ms5frdyDuFU37uZCj2HUF+GYXs4+y6vDZunFPhLwo7VtrxPd3AYztE7yUv
jSzPxEyJxTm/w+ig3NHIkpI9KIfG3+FZnOaj4/TSQDra1g/JpF7wAmkLeLiqmrzl
icSq7jwC1XJY/YsG54dksMW2bmtN4Fk7mQwP30QMkkqEiii5OF8KyyzlRbypEJOt
Lki4Kc70qfKUFoBuBnN7yKEd9XeOJrgeMX5/aTuvwXDWEsuI9sBvCg83v4XdAHEE
YzpZdcs5k/7uV2GRYUxDNb0f2ir2z5MXSkXg17P2rz4SXkD2wNTmrnA4hy7Kc8AY
NvnaWxKF933Ystw5e99Flvuv2KVi7BFcATOlM9+gegvtzEqsXksU3ngNHiKEgjMO
oVhxIyjngUV0XzKEMpvv27ICISfDgUJgr4gPkMDttxZtCUiy9A/0bjZ/4+YnXlof
YG8hO0oJL0S3WtV/ALZevZSSbX6Sm7UJhwGv0Fy+kjbo0Q6BOE2tzl6Z063eimyI
kRSegM5MQwnyGRiCKicJ5TYOKXGVmDZp05AfUxBXtDdrAQVC4YEs8hKBg5L/bQAm
QRRr9ZeDpMKyuYZ2IRwjf85g1jT8RiuEkbiC3brJcBgTCJMxe2CF+ZQ/8BOeKrNf
3BXQcR5UPtk3x36kAUoZyuPfb0eBx6+0U/8XFK7mxLeE+DclBlh81MOWNcmzAo5w
xd2Q42dVU/fvPWWLHwiStOVCb1i+nD2OYQAtX9sDkDzSE/dPpJKNsnkx3fLP8M5I
U0zUuj0IkYO3mFdMmn9fqrf+M53C1GAcpd3bIEyrt09NviJDsfZKhiLLzN+AkWvJ
sKOoK0vwfuv76fOsg243vClCpeKyUz6+jDWBGmB3X9S0wHSGFnDVXlEbXjQCoHr2
oqRDXW+p19A4THlmwVsQ1xESJxbgLwK0yg2F5/0jWou/NR3Rye8rdCmzSSBuAWL1
qjDZwNog0Z104GO+nA18xbmC/Dp+Z2VyQFNMvIaqAtcT+G5WE2wqUyzpSqPpe16J
YaXf0sXPR14RbUXp8qDkG4c1wqRkH4hyBpvq4ri55lKNQj2Az8Rq7ww4GmXksAQO
CBJBALNd8OCXjtCiRfyM3QBZSoVrkiAX01EN5GlaC5HGiqbZASxZNQJ+LCSp4xJU
bFGaq8RC229vbjYwC4yvD8e4kxIhDpa8tWyK5pg6dM0mMOWPEj/g/m9e8AzWL2fI
uxiGmmu29q9vHsoFzHUU4KzmE7iq1UD1BOicJEXng3m4PFjZBND1GN2l7CtvShX4
El9CSLYb/xMwmS2/bewKBAT/K1mbVPOhiN4rpZQ4wtUFmigP/58xsUvuPdRe8/G/
i94NMdGZH9GInEnqer/KQUsSftJ3UPmB8pZfe7pc/SjKaWlOysDdgdVOdCLdEM/m
lKGQUZ0Px+Ie2rW2FVNbtY64KMPTOglmmg+3r8JKARlN8nf8PiralGNreo7Asl+n
iZ3ciijHZ2PCWNFMmVxku8Cl5kg0tuU/JvOjitoNeQKlVMlJI5evzFsfd3Sp50Kg
vmRLWGPt4hRLZGNgkdNSFzFXFTbKF3mrIGeqZlw1JG39xrP1zViIFArs2sio9siQ
TwZGL+18HhE93GxMxQoXdkJvz2Cz2SXFb5Xzau3hacqCHpPDiCBPNVlAtmMpyjZK
43SzFVcKrg6eecRARo6CKMox1zvgQBc3tPtcpSEiHMd0M6wrKFrbGdX/WGVhw2yg
mH+Z1LMnTPTcUmc920c8Id37moiWhBrND5txFbPdZTsZUgZPWCta+pcqTeXLNKog
NZOk+mxXOICqZN2KMcE8WLOcnkY1Sm2gLmXpUAwPPST8/XDz8MLo+uPbWozYp1XR
wn/61X3jxTZTzGaWMo3zdvurvyV3Nq9BTtgYtPIWSHfcKY5ORA6i+ErhqboczZIW
H5DiPGcUZsLL7RSL+HOYwKeco7uZka78vsfTxGvIHioUJx6KGb+Tc4neGEh/42iX
HhET5dHWGhIJYPYUrh5CCvYAcoUJHYMBTeP2S0c8sVJbM9ZenRBnwejWCeh+VwMg
LqzfAYt3HyuKHpCBjNs/76qR5atfnAwEpGNKIlQEEgoqUZkiXXnSQM+SEfIYXxNS
ASdk2VUHmzDml97Ijen1uzmxYpleD0awTJwbWN6grTTSFkoHG7KLb1EueaPm+gKF
SN8n66Y8cOA6WeTP2Xjl7jaooaT7R5XGJmLpxgrrXZ0DjyXyo68AEclX8JbZ4SjR
ggEozjczFKHWIa1xY3ZUguSQGYGZOEdrFW11Nb4arfukcMTW2M4rfVFJiyd/3u3o
E6L8dWU4Zr2rwuUAb8xQpfaQuWwtsLa0N2KmQWhVklXvLXjjq/g9TsMqWrH4byQQ
dwL7BT3CtzvoEQiAex6IBKyQHn1Q59nSMYWYpTBWIzy/5WH2G/htCMHtt0t1UyBw
9e0yY7gUs7X4Vj09wnCrQOfkDHIv53jxNnMB+tfJJZRWZg2PcTajLKAioDum7kdg
Q2OeWM9D88cVh6pFcMHjdCAFRriqFVxKu0uWcXL7yDZiJ0J/V0z9hq0LVxuTXYiv
LObP7X0Vs6KD3A4e+T2I/n9oZsVbJgtBiBM80lpZzTrDClaLNEffPh2bxq8hi1wm
bY5U3zT+YP4jHqAn9qrKDQi4xM+1mWIVSuat28vqwh2qHAW6KNKXPu6AItYeXAVV
glPXpusLsyx4GOyaKf7glyCrqrGbucBBvIF9GG4OdgSnaoccJLUaeFwy0te2QS09
FWBtw/Rbx0Vk2xtHGV2sOYZ9xb50jEbnV2pW7DjtWL9coSJrAqhAgwL1hfV22v4I
DmpzOPJpc/HQxP+N4OOyH16F+bHPGNT6FF/vqAcERnR5tHu/ulE4TQnVkFOinKoW
VqdXK9ONK5GUSFe/P1drvj3sLQWxAfipioOaOnyxCcKpwMIp46NIecyNsR8dmWzy
zO6sgH2vbWlwAM38PttlRTo58xzEEPIUKvy7w4lSUGlDmdBWqfgJAXrDtB9Xv+Yj
Ci/czIgfyfTqxqTwp/rfrymU/CYCOtPhz/CxaGGhddM54GHz7ZTj3Uih1A5Z4+95
TD30BcAl8sx9d0DetDFeYpMqd/Hvh7JUU3W5j7XaoTGm55KsX5p46UIt0gKeYl26
E0V9WrxGi9zQsCI+tVWoxcimx8LbZWt9MTb7371LPR0nkN5V/q/Lb+UvATQZ7RGi
pLHhH1Zi6ilTDIRAlCE2X5zERqTRIE7MP4C1kBizO/i5SWM9Ij9elajg6cISolxu
XEBt/IGQSx7KtScEZ8N+UXOehUPjr4RWc0S+xGWwUJw9+B6Awmshi//41wMwvY91
Fllg/9PfWB1veVaA/StAGAj/br5JLYI+a7QVz7/dM8RS4MFf6wVkUFTzCKoNb+vf
VqCGJpTIi/BCE9i6dxjyFI+N7GeJbhRwRPPw16kUIc8veVzh3BB8ZUmyxy2Hy95W
BZF8RAwbtLRBRkX3H+1j99d/iB8a9d4DhaZiSP0SGEZjl+2WaGxeCQOCQvW/KmND
0D09h1rS1yFw/lnPWFbGnB1nOKKrCAh9l8vTwObUVDZYGrEwAP+HzC5TBX+FrpCL
wZ9EDNRTLkDu9qT5dpHL0a8qaV38wluoVUImQTsPxgWRt1Sp7kTbiU06ooVxqeRi
iQuJYNR0lrjhAoimpsPhF87qDZHTaol4yjcHf50wKkcpzRR5AI1k+wHwwiUcHrWt
qEVgjNffhjOAyegSiVmkhJVou5AA//pnChAZPeaDwrAToI34iLDMRO4g01fd6RZW
HcExJVxWW3uRFHj+BnTAlzH7fWuLiJulARR21VQi34+yikva1E67faZ6hzm4viDD
gUfrWcC32pZmRfN6aeuQaASzLWF/ByKpCBjAd7ILNd3AFXGQDSJD81fnzhkJ8ZSR
uwCabkMZ9lTmsl9hPLBW5SoN5RmjOxsecgNYoWxG+x3r7bPyrcgfxOB4iNWRy/2U
e+TjQWNe+AhTATQVcOo9JNewsGEb5SwQJc/Zv6wyjgVuJEqPXC9qb9rAwllQn1P4
LzFKMLepnKgY/YUpuU6dnAUd1510GmqWNqS2QhkPa+Ry3cOA9fl/MJ88mgJAS9qn
6XBOmBi4KNjVHIH1v7opPc0s00gzGv+ieSxvXXS/3hThz6BER/iWSkSMcHb29EaX
ZYEdKhHBioibpZaTIPd0fVQgw0tQYDl5gcD4ynf3HN432FkWhqkwOA2vkb11JXFa
KojYtsh1lo1r11yqjzOapbdbiHCKiPD5jTFfqO69cV1c5yPBU046Pln4C37PAXYK
G3VxbkO2fO872A9KaxtcreMq1QIC79r+l08U0VONF/7AIZ4wRQw9qTMsM+sE88pk
34n0GmIfRd0jiKrFkI11SFxwHzaEiQTqoZ4SdJ5RqMi1bvNg93wMkUQXXWeWF8Kx
bIbnuuWtKqTvUh2Extfp0ebRDN2DZ+52aOitn0Tit89b9ZXoqatruikoGfIgKBSz
lAb+vgE9lbOAgk4LiS3yLfrkrTAtF060SeeJB0oRDQFwSspI4+i69TIxbj8qK3XB
/Jb1570UoWCOGJvbyaPiduGpfH3ggbWslP579NpkwybLrdMyKfMC3ifE01nIPQjP
AuAwEEHj+9azP2wgXGvMj3bjbmQ3UODf7jOFtLXCOFDG9urXZj4yvo438oU9wIzD
tzpH3/EtXaJV4aEEtHpnGfZ0gydqUYsj341N9+Y7YJLdKNSiV9zMwRVOcLHpdHAP
nPxhh1hCDWvbObYab2tgK4NtLoMNwnOWIEowDg5ANXi3S8lmjL85yc9kac8Phg7D
/FrRDxpjXYnXWa0N9TS/rz8GF899aD4UUlMs1Wocd0Qg7cGQAuKGgiuy1iSwpCDG
pQlfDH1cKt1rfG3herRS7Kr+UFRYkoCex0GSJQZLyOgB3cknZb/Oe3A2y8M/LRqv
UPo+0Fk6m6fRP5MtRai1O29XRZHFcv0fU+kYnw3Y+wQcK0lRefphbyCdvop8+bdI
9GpYD3+xIsS6xp30P/BG0AxihMk2J/G4fZ4o1IPJJQ3ZJQwwUX6V0REKS5C0irmW
laXlfsGxOqUEijKT7Atdmd44rA9t/V2OIoqv9oTTR7yV1X7exovshgaZxKTYDOwE
OQKEXYNSe69TGIWv4lIf3GlSvihO8YdD/5QldAk0lW5nt2my3MpNIQpKlTn84OLw
/2KiRgg0CKPK+2FFk7ZlN6v8aCrnm/4Tseqq/FZPZKSR2F675DGZ50+gW9q2FeG7
oNv4LjCjkMWVeu5Eggx7/zSGCYxG4zO3NtdgKKK2MiDhAS1ULVxGXDZqu+d413wb
uzHC+70EDx38pp2MnrK0995IEDSCUxSWeObESZLyjWMNToEAFX28t1Fx3rDhD1KZ
lhJHCqGHGS780OAoF0mBR/Y68jcd/NpKL6FdaDsq03E9zV9i6l4ZHCNJr8IVHAGj
HUyDOIGZS6sp72DHWrK6/UdrJMkD3elolTdwHyWpafbAqR7Qrz2mmxJB/oa5N2+X
sOvFAN/oUcR9PknYJH98lBFkgzfDJNlHIPElPaoDsS22+s5qHeUFy65RadK4gxWF
lw1JdNcJtGjEJ+pt4c5C9lzWle24YVpRm4tIm0O5rTiHDGBm2cccTiG2bMzdUDGa
KdrJ4uLBu7yVwj5ot+tGVWOgvvg3Hzzd7ULzPpAyj5ClzBJI2yAU1BGYBJEeQPvx
ZNGnTtNiE2ogi6PUegOvth+VMndO9QT/76FkOVK8+8+sp3RgFOpo45MIhoPndokt
yPzT/R2POoJv0G1lXSLHB1mRZkOSyqcP8gd2rWZPsdzTxObdS7JOcZPTxmn3PyQo
OeJD9LvY/UD15a+5CB9pzZpgM0nAItdBcc37oPdRUWF9cSOkmwtARm7IgC8U+XT/
iBGJxKFMyvreHfm+oUI4AfZ1XvNf+HUX9fgUmYScoGqcQ5/yCdaLb+dbMCXl/uGp
Vchhpq5a9wRZc1jTQxCrTJMtYacaCNqUi5qC4XfJBQet2sEuB2x1vS53JI93aWFf
NGjuI3UXo2YVaB/3eSouJqa769FAWsEhiF2GOp0QK1wRSeLHOJtQ7+5/DsSlgNjz
sZP7zJUXkv6nbaFiQfFlzx1WEBN3WcTHFVH2gnORQys0UaSizdXA0sPZtGML/Nnk
oCFQxVXtRPaGL59K5aEA9UYt3nvXqmr7a/QuIpWRusVOO8liuWAbcBZM3tNf4ERX
UGDbRVuNG1Oxwc9yRCmbX/YdfPRa6/WgG/9FBGOIma3EmkDFZ1q/mueUGLkIO/Je
vuYXECcsro3EPCZenSAF7ehCzmkTMsjRM3cv5g3jtaQaGcyuTjEe/9QAWhDTUfBf
Cgk3U5u11OvWwISSlEE8S6fsMfB43rMosSgXaLNd19SMi3OeLhJ+0Pb45vq77DMs
DkXwRWCRtzKN4ngj/GZ95jVvALkYcmU+DoAc0f9nBuL1QP4MfIgxBxGSg4EmPyUM
mrPEsVZkOJoQ3nPjGUvQ68AUOPlAqDzD8RJb5gv+vSgSVoeiJLx5cCEBwFTfiYow
g8Zh/qONJZ40gCPKEW2aAuYi6NI4xLM/U0IutYuBbyohReoo1SEZbJlvve9zM5mo
4D/gXcUB6w8o3Ty7taaTf0f3I7eKQxAib0363xyvkhYIO7Dg+abCj44SyouVvU/+
4o2z/95Ew2arHuqM1V5vNGXCi/X5sCIPOpnz290qWRjeOwNSFkNlOyt95APXKAid
9wSRflTD7Tb6KVw7F7T5/xTXIwgsnDZYtWoAi4ob9EaCUYbBUvxNL6CcVsBqkQ/J
PWt87MaJMH3rCBiQcGzDvUKB6BbhLXXMajr9MZO2Fy6mpAcahudlw0XjPH2l9yJr
1iswKnMX1r/v1WnF0ylLHoFgv/i9iRCCB72pn1eaSMM5Ch5ec3f7i1Om4Vxo9MLD
Dn6ps8ihZ0+OpNkgyp3BfeBk0OW2pf8a8V9YR3vSo6crnNuee9jqcwo/IRSrcPUd
mjzRpOma2Dfj9i5IIMIhdsnDhacjXF03iFeh0RMZwsXc5RBr/8OE7+B3qnLAq2p4
s9Crw1nF3BHYZcDHTGRHkj/9dIt8aU8XfHic9NRObdElOQg/eQbbow7OGSJ+WQcd
WaED/mGjufU9kVtl3Kh+K2vWBZogzfJ6Bsf8wK2n5kx1ylHexI6+pD1sAMaHcRCL
SIkgbrceRUPzxNbDw9hV0ihMpjtHAEJ/g47WfFm3xwPj1pyN0g6mkfbvWp1vwjfQ
hxOqLGd2N2VXFn3ASaDCtWp8mCHAMxtoeB8jD9tuNw8ssqwlDiz0kwleaZKX659U
LQBQKuyuj+/z2z61hkMIQCgL9j2I4+jB04ZI2D6TsLY2CUqr/76u3nfkPtpWizg+
LTOyYzINqPSGwpVxW1Ry49pgdtWdV5pnv90+AN8qPnq1mkqjOhxaf+NZXYHZVPyZ
S+mIzo1CvqYs+R1kiLMAe6+0IR5+l5WqOTzR5bWcLUeh/B9vLL0+1yxeUJGRVN+W
FaiLFn+BJfjBoRgZU7pIOE1gdBhfN/G7vI5eCWJX9T4=
//pragma protect end_data_block
//pragma protect digest_block
M6/trQhXA/k+lW/svb0UccyWJmM=
//pragma protect end_digest_block
//pragma protect end_protected
