// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
kqg2u/vrnaHruRF65L3HZOVUQgaFNlHdS9+bAKvNJ435x3TomrBV6zyMTrjZuqD0
LmXcSd5a2USVGX+3yEJP0DW5tyxojI/YPl9IdxzuQ86qoEv4fkNgZXxzIpespclU
4fRgKjL7xYAc3iXm8qec6uYZtuxxikpxBUHJFdeop3U=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6896 )
`pragma protect data_block
YQWBZVb8HcF4y6aEwUrrfBXzOzxa48XLNk1sXkzskBDFRsk2PsW9yjLK9DS+DNH7
jh24OY+IPQhZtF1RnAtNvdRRGW5h97lbjQerwL5p3NLGg0NetH0anxyqjP9bSFnZ
S4Pc6tgYkzI4xuOr2il5PFeqvGgduWeh/vNNAaSTX3x1+P8hiryNFkg9n8Mco/+u
d/Qvsuyl7Bc/n5cXa+MMRvf2ewYw2Fz+9B02kSCxZwq9dOFfvdCJ6oWCZPLIC2fM
daYzrsJq07rAJJZ+urkCQ6qp4sW0II1J0WHb3zyeVEkxHR2riQr97Ei9gA3cGERv
heDvKINMsU5VrruwUyAf2OpgmNqXB+3PXlzFRVSN/1xhPyd1BsmYTSjwgxE2Xu3H
rmwYSKomKn4jLYtnV8U1eJCDqPeFgpVocdbrbbr4pH0lJpLiaC/mLVF5sjQrpfKV
vuX1NLy1P6X7maMSnKMLnIPTXos2XIQ+NsSpQ6wS/Dl6onv6DyWOF+WeewUm9rok
456SC6doS1tLKpjjOivjIderdGulddJOyQhHExwHAcPNUKkaqjKQ0Wzz0Y2n8b2a
ModLKe/4U7hwyma2X/om1vt9XbJO5dp4Lgz4H17vXq4Niy4I6i6PR42uIr7L+WS0
lClrod7XdBu5mBH6y5PvQlAU6HVV5BkUOMLauaYnfPuQVR5ucbNBvmqcdBLoQgbw
ow9jJG+VOuJJwtx9H3uhI2Z7CmyaGPxG48xRChzzDP5NxTdmmE424RVN51lT62ll
htPrFmfffCy5ie6VVadF+gyZam/PSQXtHFEHdflurZzrIzc00BYeDxFSPQjrDVOl
zARXs/yd1fOQDc5EWwjJ1OkjuEtehusar73nfjFxzRLiDkn519mx/cotrnJTUdMR
c0ZalxbXf8kG4hKLkafW/MbgPZJdgK0qd1bICQCyFKOmA+hMCL72okYF3w/mvZgf
tU4YLaA99UaISU83b2epZnYzcmmnc4HpL0AkxazyjJOxEoauCckAg2I/mSnZt0bQ
xUBV3zkc/M5Cm2YvI0cr+6e0klDj/U+mKN3r+Dac8nwbEHTHdcuSzKb5sSIpsmum
wWGLVKICDJ0V4Hy/adyxvMY0+MNwstA7mROJTwfMOaCcshXBtdGznpXh8goYsooD
kHgzzWZ8lHdxPc4H6ozzypfisOtjs2vHI3xSccfjH1befA5sycJWcLH++OXFz7TQ
1V0DU/6Md3UWIc0XL5o9/1fEkiMB5jNK0eV6c9YLLMmfm8nBUtB10Sw9od9tLBxK
dT4381pDZuURSlisteCV/4ytWj/UpIcdSwo/TDuVhE9vIbCXhynw14MdcSxvZkx1
WCLy+rAcaj/gNt/gV/6O6aspIh5kZtM7w2sjkUrpfpPqSAKy3eZbeA1HsbyuHl6V
ICxgleGTG8XCPzuTtb8dwJ1h6ZqwzYyyLGSUn3BTaibSKsgRKHy9qHaArI5Amd2v
lsBGm2QKqy3pDw7Zn1k83/eYOMkkr45u6XDKfE630JwYNvZjcxzYN2XwXjd9UlCR
MvTEpg/CaRZulV+2wBjW0SQSLnZQPgyRxiNxflTbk4mwg7Dm2SS9qy6oRsKv8LOj
UtPiSmpZbBkJ7DbLuQ3Apif8bFvSeYG3p4lHpwN7pZKZ0IppnWZlCMrwcyepIN0Y
1FVpTN3abhgjZ164q+cUzy4yihFe36+IdzfN49rH7i8YsdTb4sV7Z8iPTEiXD40j
tj1lMNXwKxRLk4DQsmbUAXAABLuX8YYi7taFtCXkGiSb3Ai3ge7mLFQ2pchz9IWY
D+sJ+ueMbB0hizyOP4IeXxNFhNS7BXL7QfbAYFZcrQOjDFu7YvVeikPsxHEq0MMJ
mcD268xvxeLJU0BZkYum+Fb+r9KQH9C/5gkxEwnS4uBJEZUS71Q6jKRbDGhrTghl
CUfpsUXGXHu723wV8EDS/ZflXG/xny4fR76fDA3hWTxYM8uxucjxzzvl8uXnp5fe
9zYry7RXri5JY1UCZ7e4vnr4KPU8/DZEBBvtNH+tYkljUaKuMV/2JXzJbL0E6NXq
E6FCy0zwoDnMNF/fDWExFrlICnwYaTs73186KjDUUokM5oIPHOUtTvoFz5xv/7nD
FI4IyANGrDLPn1zamANWHOz8s/D/ZqeH1Wnia3eZzpbpbOjgkmMsmO22vyIeDqpr
xJ7K5BIM7fFftgENbZ3k8+tjdzdlNH1foAOCUNrFZmgTPd+jjxIjq+yGYb7tzf2o
P5vbVviGS2kxHvqtbMXEYQYp86vJxdNjHIZsFwgxzddaXbPaICU14RO0Qvh3Z/lt
GQTUWLZEXnBk0BxBiSj6AikpknTB1meeUWs0LIyvj9Y5dgsJfnTvgLU0GaLrFM3L
/aq7i+XkeCbgLdEY5t04GwZ6Y+oBEMpkkQyo5s3WKOMySDKAI7fQpNP+kCRbJnmq
c/A7zrPQOzLOx7vdRwNpXvpNKGW/kDipgqO+052+qSnHpxmxNG6wwP5Yfeb4z2tD
T9iKfaMXm2leYC8VmmB7fG/yxpZCcn4lXnGaxu4CqZIYWgDFvMFjRy/DdeWyn/7U
ulL33q7S1/avQTJ2Gum6jDwctQtTCeHqJ+Tcik+rs8cL5N5P2mjvOIcb7QR8IwtT
WQ19AOpCWFDTLQ6rgAmVIignbqpDhrdatBZUjHDwY327wEWHT++7O7tNVNbjPCrw
ItlPwDlaA5YGagyPsfHJtNa9swfv9sMchF4yrbBQMT41rueF7ijBgQNQOg3glNhD
nflrZYc+/B6HTKrH2I7R4GptWCMNqCKAty9jBceHgNiapzxAs/0MGIU7QeC8BbF5
HEt8gtd45OquubcxXDhJBOIhr+2kfglZexqI6N/BcsFkz606JEwHiXKEskHzhhOC
rYenBLvQ0Hs9sUNkeI6Hs+c8DfplhxOdTOcTf+QDTSocuxQFoJfr9YCKStUT2x9Z
EmzISK/oXkI8wSKnJNGzWmFS+0uxsw56r47z4SLwdVbPXvaFfUgZFwEidYNwa1wp
RH686k3Q/5SoNQgfxBcPvf2lmkkHCw3WuUmTwEImpxL20np7GmHqdtUAmCnp4Nmb
GxuEoNqavv3FjpL1FhIf0hc3eAzpug5wdTB/rRPJIK/LDigJ8JlZNM8pukbFo+be
7h6jY+hQ9XmWlqhKWknbAdlYIk8R1G3lnZ+qAWc39lU93+DAQDqJi/ShW4Blizc1
IBuy5dqWf2RAn1SLrUHBXbLh6FpCdI76WrB8J6ft/DE6wK6RzoBuxY4vSBtWQUP/
gQUojDL77OqOZUPcdccTEeJJB/oQAKn5FE9PnQ9sVDOQ9KO4r3Y6XDG+ebERwvzM
txBZBYHu+VLoPa26kBWfKactXfxBrX+n/s+vBVDZ2j/fklJBIJSWP9IaPX7ZN8JE
1tTSYPNPPEMyejJX5PdERHPdhyxBpcvfLPRNxBrNQ8+Zi1sXJzVOIK2n/4QIPVZF
YRdwvzCpPo5hEM3p3NKq2iv/uxaJk14a10pQ2d2l6bRMA8vbEs9Onf77lYQSXb3e
wIlLt7/+dyzfZj8aDpkNmvxVHQ67b0orQ6y5F6gtbOBtlDzMx021e3aRwgSvv1Lj
7dRJIfP/03ZBu87vGOVBzWP+/ExRgyyiqQdHzAzpeLT8xSXBlMf67i0SgfnE4w+H
AuSnsAiUCfkTK8qK81M7odSN4lni9itxj4o7r4VNnW17bvIlCowa1e/bU5mh0IhN
5K85NxXVQSyEyTvTmLagerfYyJRisBubNH8neC/OKYpuUrJrUZC2x3vkLDRhsRJD
2J8UutvpgZ8OtCJ4zY4gGXrlbc2Ijq4R+zYAOQh+5yArgNcqdExtZVl2OP9mRZDK
mI8Srl6gWSAv3jUiVBmR0G0gRGPXPdGIXUMJVnVgnsoe/bYuG1VJ7U4n75luGgXH
CzPc3J0/5ro1sXNWoB/HkJ/LeGYhCyHJbyn8znXvKe6cfgIVhLaKXqLFrevKYQxn
fRUktfSUUeDqZpPS0wrsLkfQ4lbGnUX+ON715zuRy/lq1q+HHt3ugvlD9EzW2R+b
/kbo6hWWaDzv98WurIysi01uzd4Nc5Tifh6WPAQ6AKC2OeNBZShg5G+3k7nuM3Q5
8cQ3+TYNnCkOp3qBMpcNarnLujS11yC1O6bNOk5bVx3AeN3+fvB/yBLwRtFBt+6Z
Eg4buXOnHARPXzGKQ22RfdvKnFtrfWC0JgBlQpoYDOItfQn/0mhAWpL9zAiimEpZ
3skbwUPgg3fy8dn3W2w5WNC/qHpXaAD7j4t0YZfyCwscp9jZ2xrlNWHaB3aF0Xib
UkkSY3uFOQz6GV5AchyzrK6HEQOANkyR4CakAs65/2o73uRr+pvOlT0iiSuBVB4D
4giXHA6q+Mgq8BjIkr8Rwc4dDa4gukCAB6PhRvAxuoJgI0Jj0/GayGBKdzblzIzH
xKotdjc2z1aqvAaHr5ZA4AGPkNi2z93WlLJ6ofX6UBN/09TasqB7du9bGcQGZOgE
ssTBl12jxYwd/P4K4b4LmnnJ6pmPmX2ffByLqhobNjOsm3SGCHvlaD+Tpy44t1Cy
kdOt7bCxDRA02s9lZ3DQOXRK40iP47teo1RpnTHzLUqv2ez+Kh7ITtg1Sjr9wWFp
NeystB3SpWJEa3U+AZ/GpIX93jVrn9ezxGijQ9SKzKUMvQDvgMkVpMrYkWhqgp8H
K6HDTbTsvPzA1WycnWTvkQiYDF9AAfzpik6/fCqN/a0wf5T3tI1AyyD9aCLjBnPV
sIka/b4F3YWS6WPahn3G6EaHTdGiiI+9438yNiNY8y3xddgcRTS1OUuOOWkyasK4
7njmHK8OZW1SSNFl2DLEN3hXSOX9Q8PfrPmm9YAIZXyUPMf9z1fZTuWlWu9FxRfS
ySpfvvkBuCNn6za7Tcbqf7CvNbzuEvyBcedcwQIqJU0QwdlWVr+Po511znirH1vC
R0Bqas8dspCpKb3nmrU8olDK/WBlp6beuU/hPrYSIZBsNWmIFaPyPnM326JHHRLH
MNBuH7Yz6fufwcz23t+5jfwJsGlMB4aRYEv9heJGkRCbJKoooweC7e07mnVIeArp
3ZcQbOFNp66eADb2bfhfiVYfwMZ92VzgRxXt8Un22OnlZ72j3hRbZVvIydqoz+EN
7rqhma8sc6XGpmYKfTpKAGPQ1qXL9ypF6nKS2mUU9y+vDPshR7wftuUqhTBBsb7A
55BzFTtTdcR+Gq1kC7ICe7ndM9GtwlIpKvnrfiuaHNA3Ti96EasFf4rR/kPzIvop
DlURIFirQP+FanGEHHuvdYmb3n4mspdFN2ZL+Uug+7q5RDFx1S+BSTxwLH5/id9g
YUb6mjuyvTFK+AEWUtNX2xWW+NcL3D2ReeEKF67cs+fSWmMotf9ruwRnBxpZ1Pj4
Roiywn/PD8i1Z8q6dAKIILv033ePZJb+IR54gIXnhjFFs6AubHU8wP8gVgdTwySj
jdP+YLYTZ40W7w12atyIP/8YLXRdil06ERbltRdsrOcdzBsUp8WFe3QOTWbjvPcz
1eHaTQnWkZRObZazVShuTNYw860VmbjrUKhel+heTJm8Ce/hXbR2oHqos6uzQYDR
+OjZ08I61ZiIX4Jkr0KdoZLdD0OgMwcE4THsIRSHC++On28UkSX8Wn2B8Lgd9NF8
GX8vG5/Dd3MGxjwWSzoHxK6IqXc/w7i+4iIk4YcgFdeVDzuU4nqfDgtY+4AA+BPa
HrE29CYwDum0AgtINmmNavU1meccpPTWnqgHSXNobT4cwHsN4U030Sj6c77ROEgT
Nnlm8cP8iJzQkAE2isQvxF8gb1JaFNq2ns7wLw1hBAD7nxWGb5apma1RdHcEEVW8
zafCbQVEEs972nWp97FFsNAB47u072OuTGBtyE70ayxUQldkaTUr5ao3sNLqkPRi
6WJQBXBNUivIpV8edzMjb+rW3D8CtD1UfSstmnRCpoLSM+OPKEIz2LoAmdMFVdPd
Lb+gv9NNB9Wq/yi+kVZ2fY9hddWuKDZwgLgPTxabhWNPz0bN7xbgVzn6c+x8DOh7
a04YQ3MpZXPRmWskVGkseokGJAhumK4CiKuS1PTSS0IWFVM/iLDw3wxXfKQCn1uv
wzDs651lsFWES0iUIt9v6Jhrz1ngGPqW0ubOhkZgg/5EdJMia8PzWmE9ZCVJ7gaK
IuvJnvli08/zvdqLQIrA4lSWtNqDgeZQq9r8a/Iz3xtE9/gioXq/XZbpHl7a9pAB
mFeH5Swz1X/ENYE6O2hYw6HetBVYec3v3+GaVsK6Bgrh+1PxFfCi6gO0JV8khOoJ
KUZoNlKNQlfnmo3Avy9iwbvyZqTT6hvQP0gcYqpVLW3x+C1EjOURraGBRpO3AIsS
ptObxCz3PYCRp4X3aRAj0kchBBf2dG9tsUQs8FHliDciHCWWEPVf/zvVReaPnP5C
xugswOhL0VDXX5nLv1wGFGJ53g1vnLOUx+tU31zl6borTotgdM1OodG5UOSS3tRN
8Mn2pHuEvrI+xDRVQ4EJ7J+kzghzdJCZw1Rmgn+k/LMEluJakSrSOwYm4cIznWJ7
vdKT9QUvxcDv0y/rQ971Zg7pt23G43FxIWjy9T5eWWtSCvjF2N7eWFzOfFiccjSF
21DlbkyF+Wgs9umRoWFwFMaf4UI6cwalaH4CbuXvo9smevEXG/x1qHCWxRvoVwU3
ypA9wr02ygGLWx6WXiqdcDT/Bm1tbKMDIP6qWn8z0rkLDWCQY7P5n2/ckkClUPMZ
NwFfMCvfurmnkgJMuUGsx7z0sKJ+dhSowNYVFNvh2P/IZaVV1deWFvJzq/Ty8sX0
TdVkJrvtDwW5qc61M3L2746nfCs+tT4+sBy5eHeznaV/duyCFCiovDKE4qKZqrON
eFPNFDELsGGaVBJfQzdAW92eJjkGc5gokazN0pP7cUehu3+evuHBk93jnmUgogyu
SCJZ2NzoTc8V4TFxSukgpuvukhqU3PxZC12bQQ7vykh0wTP81hMt8yw+sr/tHTFB
VGdK5bKPsJo7DQ2LH43Q8FgvzCzW7D9lWcH6SDRcHKZYOVW6qFUcNzh3XbaLt/31
B+WrdkR1hoSIGSOulXVyU0yOYNT4MQ/Gl0yi0VWbiCTwLh5DelbiFwNGLy3ghjgI
DG5VIw/E/QfGeER0owbfupfdPwkQU4HJiljlp9n0gKStew3alQkztBuSUWMGYhTH
DDcI8QaqxPCZfwJxTwrmafiwCZMpLNVmYYnda70fAYgNL2/bCvtI+Sq8J1DbpeQP
TSNynW3FEA7qJsWESUPinIktET+Bun/Rb458jY1URT3jA845XqY5JFoO0myoBpjf
JitP+fR+16xd3FSDxWHqhONJBdkEGUIutC+2a3rMVa5eBNohFpFOVU1qDNSEgiAE
i9nv7s/aBtdN7HPSxxAApkyYKEjxH2dg31UKIM1S7gLqeoSjdWFDZuDoydkvng+i
GsOiVhBtyJQyNW2BVt6FPH+4rFADVg37CROiE+UAgbqCShtoBnEqujuo/yL/W0Vt
/EW2h9BX2yMJKt/5FvL1spmxrjC4pN9FSBFd95jRGa6dYQf4OhRoEjY+yhy7YS0R
AHTxm/S93A7miJXRzZYIqZP9JDwKVg7lMJa9IsYIVLf2x0J2/pH1urOQFUqxIGO4
1AUePzxCtkCNnJpAerZ4bhDJU62OR2fFdYRLzdxrx5W47Eq62rxNLFbIdHN45nmf
TjikSlKOWMJ3Qm2FnuF/uM5bT5mdSfyPGe5w+/hIauSLDHlJCNuVoaDHt+bflEgP
xamlhzfLP3iTS2Pi1lkauezOgfgPfLr7uUXr1GJuBKQ1y+9lJlBvqcjiF7ORawUJ
oAQFdSZS7rx4nA79SDtoxfRR2bQajqLxB4uYvwEq5JoK9So66EPLQ0pP3bky0CX/
bxXsDzoxC0qypqLcRwdW9/HDPUJoLJg6IEZgUSeg/KFJ4VnzP9cMU/8AMHCXsqSn
SRw93CYTKx4tApoOmzFlDmPNnvQSUgd1slx1Lh8D9jOXaQsRGjYFNDcASuTKO1h+
00hYC6acZ+HMZCn1hMASFHzTSm7Y2j06uiAMgfYST1ysC3WiCp3jC8Wr+6ulZLS7
I+DqcRdxxq6h8gTeHm98yIbrc/ZG3Ig2FSH+XRfIRh3FamK4vF0KQMw8kd+Wz2vj
v60Mrg0M3pokOD8tWhsPCsbb2MrrYaSrhPbilOQn7z0rG3iPOCgqYzHqFqWqm+99
NwjLl9el/2zX+Xfu3fYhWrkhTgQhdiRmJ+HVjIiwOqzPVz6YyLZuxzC9KzqSmgr+
5Jt/mISUc7y5K2thurEnN06qZGWRNNVxBxhP4uTf3Bfc9UIS9Ju0OdpiglP3JPKt
XkrbMbgZ3bduPS8I6lTBxK0iL8P4yT2p8gSRet+wW/QvR6IOgAmt2DKXs0cgR9fG
YKRp3H6qvG20kyoeyiRXnSJMr6XAKD3lkwoOUBXVwKgNMVeVbAXJRG6JCr5JkWS2
oWCghovQHEBUPBNijN+/8LGCEjNKaqVd5aB7Z91luCLwlORiXEhn7Qk5QCTuJMIr
RJxRgrN+la492R6rxQ5heJpkhSYMHSCaE/FLSvA/nq6zscEYTpAm6ABms0GY55a+
l8PZ0wgpX1WsgdZu/CNUAQ2o+lDVO1CibSw8I9uCNLXn95uC347guGeX/9ES0R+c
U5ULW26wsARwrayDxtHPnQMcG5lf6zRdd9yVhwv/eDRgNxB+C3GQhzTR9pCQbC8c
D33mpjScTKLHE5ceEYZLECweZcuv9tPqswbV2mqTxQof20WbYLFDP+DD7lgzRPT5
jvT2wqRRoLh6+/yPtEJ2g+SGy2AwM4O8eclqC7j0yuChGpPQnwShp4ucfxpPU8se
Af5wQ0JWj8MQsSFZIDaNEqog9HDr2y2LQyzzylW9aw7WhiZ0mqIbz/jm4Q0o0yj9
6W2lAHWqSp1dlEQcFZU3gB7ycEtsJJKeUkJze9PJxwL1kj3iu1nalnRIeIr6PaAb
KPURr2eRu5bmC4SBC4H9GjYbzounI9lL2RcyPzBxYI2WuT6S7yhU1QauO5CkF+hC
1OPmtZnBsm0RFoWQXrS9xprkEBuPB5FmoDP0X0wtBK7hkQ4tOuj3KZAH/U9SVzSK
xQE04O8mVWfPlPBFdfnh8sSlcdxB17kGjTouQq724VWBQ0FTIs7k7Lt+kj8DqJ5e
3vee5igRY/x8OUbAZYiQk2P7lA+uZj8r6ISXjtTs7II=

`pragma protect end_protected
