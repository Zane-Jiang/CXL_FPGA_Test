// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mfgElIqbYio8I9m1Oa0RYg6shlkyFLuvUaOtZuVERiwjY2gibWHdbi8zRE97
x3TRkkQUS5KqCqPB3LkDW6dQujDqnlPL2qSFzBm+ywrP7tqHXhjEzpuXDYhf
0TL4RQuZXVwJGyXy9LCdTo2I9Txi7z+/hZ499fWPYzHj9lUM4vl4qsOlyQZO
HbEmWN38GkNVKtCT0rIMmUmpmLb6PmhLA7s4pSfA1/EwGsQGV3kdpF5gAPby
A/QRsRjj6k1VPEucaH/O91/1TyWWxpAUCN4wMDHn++QEaxfyRyKCj3cYvXhG
AQZWefnVwxcggWSE8VXRdvH6DNjRGbSI5fJZxly5kQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gzV2699w02p4+I20Vvv4TkrTfWc9+SaR8kc0mEeQ+AZmUn9/yq1ZmjLX8i1d
JpXe321PwgAe3gCpz7r8flnxWE6GBxwgZRdnPiEgGJ/vkaGG3yQzwBLMQ21b
6QL0YulY7+rNYnV2YV+J50Nb8nxZ1S2uPbcbJW6PiGvjofhbrkGrKzjjM93E
0YIu1NGiT2fQSDigf3qztE0QF0D80PbTEhK0ZtIMOrOX3rPCCrjl1zAxFMyR
KbBs3YKMd33AZaBgNXIHimUdF6yDIpW4gbdPSnzJwyoS105R9QNdbWS4aI2S
cl/u34GOBjGCv3Xm7Zg3ti59CP+/P1bPYPodUBF8tA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bAwAYag5+S9NPzx6hBDlwjngauAraGjhaKCASRnTDUpQc7fqRStlQ+a0EmMV
gUNmKp9yZyS2Hnw6spwPdP1etP/5BbE5DDg0A+3piqXrvroYZ94iZbkrNwAI
9o/4KatIQ6Fb1on0pU5PJbPnF/8n5EwVuUw9LBT1O2ERbKmbUttaY8XqeHLC
HKnmgUIlaKHk88z9Pse0vu/BTBEqQPGrpUwAuAqWw2OClF34bDyVUplXNTVH
4D3dnFyNH9+J0ofFBB7c1VkIb3p8SBJS4vduo5gFy13Ne4p/uFgiIKkG2OaE
4Q1uDiM+slbGHmCeY6FRlBSwBqsbvBsNXObfHMPTnQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Zq8pzKfBtOjYM4OPInJd3pWxI8ty16L3qMHuPLC8VZX9zKDh4rDETZn0en8o
MfyoqEPZ7Rp1Olr36Neyb5UHXibwPR/XYStCu2Wv6rUeEv7RDwd69bMS4kbt
nmn9lRk202laQSgFTAispjIeVipHKQYbgq8R8ELTVkUJtXfhRg8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mmTr6Q+oCH0GlTS/CxYXMeFyEqAON7WlLIVLZTrcaeDuz1F4V29YI12ib1jY
f/WdlacdabMVR+l0n9eujU5mBQQW+Oe3PFrWL5dMneZIi/HvuEkWKZGSuTVJ
P8lLCNmXKOFKPTLaqDxr9kSzyrAJOR6pd6XGZz09gc1EZoHfc6NHT1ciNWOe
MdYzSqMMNeRKOPsus8sy1N2So/E5qBZlYgWslUZffefDMnFj5O03fmtXT+gE
Ri2kfMzd9a1DAqPXfnm5/9PGnSNWBGCTytVHr+1TkPFt093lOJUYfXFsYs8N
cGPL6aYTHrpU5lOs79fteQX2hZr6MGMVJrGfEAv+hn7crrPXwGxabXZ/+sG0
/V12NdmGSwYL5vg+piKpjIee/Sb0bQFQCdT+f2WC6rhDX1KbG9mViUKXRhUs
S0uitL1K9VcgQEg/jSedLNA6x5WsRBRFnr8XgGfxpmMUafjjNH/B1WxBiO51
sf/NHE4VQjY/wu005520upB+SxGqUfCp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gxq9Dk6nsK0Mn3awL2ZCqQm+dLzBbSlt5gvmo0V0ayR8n5NCCOr270AwHE9X
qMkz7D8t7h4dZtlMM++XIj7fwRZekQ9Svk2Wpqq7BwDRFItv+muCwlDLR+XJ
GDwOefkDOZHscKSwkLRppEQlK0jrSsbail0m2zI95GsWRGfaFqE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eLhy42rwnkoXVnDVXZHXz3BFJ95cWYuu7h1/RE1/hJqcyAjWPYXgxUF45SC1
kqCPWmiynY6Ycj6aZf42OiGnQy7+Pm1lotlHAhw16+0d2u8mf+X1Y2rAfHhq
YIEo8JAKcwTCNCszONus9EGVVqJmT5A+gEOEVUvhUxgw8pJOXO4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 924752)
`pragma protect data_block
i5L0U/dfoNNcG+kl6RZkkxahmY6aZmeeTOOlPmWJyaavcLbIn/qkcabL9zOO
+nFm7n1tqxk5i2WKPg8xvsu8N0qDJT2lA3VypP5aY3N8CRR0kdNz6IpFU3xO
2nK3f2UTYGF50AssNVKOGcCKtcsoSZpDoS58aJx87A4bIhx3IhiSTjNvOQvY
wwzUjT11h2b+5l3Y21hUc9O6uZzbQt85JcVH2k6WWaNueoxwATbEyIGQYIKr
AQuO1zQlUc6lasIDdKbQwNWv1/J4FAVJlljsWwaxf3bKdYciqWva0/CSNpjd
tevE1cFTvc2TZBPpFMkOLjV4Sih7qPlIxFSVkXxxQN/2LMfKv7iouX+Nuvxn
jgxpHvWVXMQRNylMTzTarpr1Jf4ZNCN3V/BzE0afdCQEs2XFe487CVjVAkGQ
+k6VRMz8MFEBX+4Ifc4LxwlyU3B/VW5vvaAe84V3T/MS3yuZI8593iE3ypxU
ImP6QpNL46zp6CmMQft0caq7pN8U+OcGyT9LO41IcFq8qoo1H/YAs4642Kkv
sC9Efak0f8buS+6uGmre3YtRcGncLdemXVNpGiC5fOW1aCrdxRqoFLi2uWNh
bs6yI3S2lWTXo78/kHqK6meEn091hUIDa4CVxNTsaAChQlvqkzmEPfmaCWTt
+S+4l5oEY9LdyJz5JstqwBHbKL4eavYaaVmlV0HqDHE6Bb33lJiG1EFWmoOn
b0h6JR1Isf57iiSmarH+gssiWOo4hIn7sF1fIWR4+psXDkXOYzCovzQXuwoz
AesXmvadml/sb8uU7P6773TLKNYTwK/XBXdV3xYda6PawOZK4Tj6TUv478i+
X4NN4MLNOVOJvG7NlOdUyjj8jotg+5UxA1YECVY72SbRjIHpeM1pDl6gvbcW
BmboVIeMIQ9uuFZj3gkF2LvbQe5xAiZOSYV9e/r1aRN7dXBJKp4iPz41GH8L
Qzqjh/QjsRc3JyJAoC2qiAONeefVG3Td4dssjynki1fp4+idiacCpPlUf/8j
uGoJzx6lCQeDcWF1QZxgfAt3Ye+26+kIuM1kjMNYoZG/Jio24Mi8a9omzNoc
mQrKMLxComXzfX5Fmav1mQgGeIz13JlWlvkVDaVCAi580PbujrFZ+Y6zIQta
od6iWXyzDiNUWjsUEc0ZociyytYouP8lWJSbBKuiN/zAS4r8OvgBM6drKuT0
otRSd6dvCNj7UzrripGgeODCMbyhvwvjgiwTzI5lpzUDLEUi81euCp0EjQt5
PN8L4hat7sbon0li/StzJJ62wdsRio2nSIsqdVYTZ2czDHexXMdsI5BzF2Jy
1EVWRNqSRLtBYOD3Vox79Iu4BKG0F0VtkUYJM0DVJL7UjiJro37Ekz99ieK2
xwT+xGd12LMn5DdQsncfHNsVx2d3KyBc5nzwdpHR8K/nCv74tnCazDZaULOP
uyBStiq9WC3O1b0DD/UzDW2cWWEvp4wiKMyRUE/nMGcP0WexA0eD8yYMMm7X
7hI1BO5S4ntcwXCnJcMXc/MdKqDR3Om5InkniRkw+kUHIa7Ss35/AABfa7Uk
z0u4z8wKBKmcobcxq6Nmt3imXTe95XF3I+3jH4+EGPvr1SIkQbKgV+ey+hM0
VGIDagdNcSY2oGl8+DfKlbsMDNnMPi6mWrhbqnMb5Jpp52JZmdJCKkF+tKDb
hIjy6Fzern6Nmp8cDX6MN8QACJGX0c/+p6RlaLxNygpNOLQkw+oQkR4KVoeJ
cP+aFtjo8uDPF8UdcaeqoQWDc4oc99SraqFYWn1UwcIk1neYo76NAjmofDGD
3WIRvryOVN6EB9iAGFT1O8eS9i+9LgahnWejn+4haRZyrXoV5bRiPhVDiUXh
H6n6aH5h6FwHuhKA2zWCkCln/7W/N74P6U/6c4vVGfCXG05h/Cp33sb3wFF9
vQbkic45lZJqtXTSHn1pdOuUTgOQ3CjHlINgJ2cy9zO7nGvRTo+xz3lF3ps3
r6zQ0eNvSlyJnTTj1D1UkK3PT/bXGOMWey+HPWRjdac4Lz+kQDcbVdUPZ95Q
Su3fTvY9lj8DwMMscMcVVpoVTJcsex+URUxv+xow7jeYlrT7lLRXE3wIGWAo
m1nI/HjtiQsZKW+6oanqLydR4jl8IlUl0BYgn9zFHGiSZdFg0/6EMMjPktMH
ADKFQIB413MB1jgYfdJuA1qYUpvwM5hVpod9B4kH4G0Zm2O3BwafQNjFDK47
FoiRuitGNAdxpZbkR0BY2KwJjPAwW+NbKFRhSTAA/rqAq+idQyf7XvEo7vEM
yk6kuvsKjmm837bBSsl0FSE1gJQfXEVKU1CSdwurgqUY+yvCyXyF/Ctq33Aw
jhYwI3jBnzZqH1lZj/kj/Q1wf9/5W7P3bcpOTPbXgzha4Ox2zciITnXOlWvf
jzmHje7QgHc/XSUao1XPvfLgN6a1ziHKrEQIPqJ3tkIQ06CSfUXJTBb/vPc0
frWrTUUljW9cRJugf9U9WJoqNCoqOFsfGJMn1FOHkznarvA3+mljm8TSp6S2
LyBJUMCprVBsYGiM7KTPXeUPePfa983qJpds68KTbzLK8YNU0zljnNLzm7hV
cuchAqPwu8PTy7XasrpnhLZKbiuIoM/3EmmBuO1v/42USgH0vbeP6C0XvYtK
PzfmGumOrvUhq6sSuvmfje3nVFbuUoPqxnlSbhpp2e3vxaZtG9dSaL3c/P2K
mhHjlFWA1+5jyPGsMnSaYV7pYDP1tZkzZ4l/LFRFfJdLT53cQ85dyJ/1oWuJ
yllSg/QzDRWWZ/K9+sg3ZMt5d+8HXBSxAk2ffw/fwa7xguBCyNoLda/GO7Tm
vG3r04OrP17tzMBzJvwse45xqY3r6XhThTs4ixerpKWcijuymkna1I9nqBfv
mbWjxlILqAUcKZqAp0l12lpL2i9+4mZuokFbtc7tXIykyPdhDwfabfLP15d6
hLmW6v55hgiFzKo0A+9oyoxB2vvOImPmvbRvDwr03hoxeKoUm6FAOFi4Mjeb
p8k3uXvbdwX95hEYsNCBCWJsTfXtzo8YlnNI7HQgeoSHfUfGKVK5202gjvwH
NleJMb37u9P/GLJp9eUVIY1GNo4bljIJZ3K5ZiEUiky3lyqvfJTW8VtN5Jfp
4WuxOvDe33SzmK7huSTtQLNw3nLjfYccbCy/RJiB+pplQhLNNAhnyT44ZpX1
kR8NWvsN/cJduer8fDlvmlguHY3YBDv4EfT6OBZHRww4p4vnFkgJNQazv1uH
1w2KyYZvJJLjW1SqmZb3zYgeNH3tRva/1AlBJd8iA0NA5WGIO5WmetIO7NgS
RqedkAzOWwLp/0+pG0oCKyBVsuuS8rYA8gRTrdcztHiQDtnqk3CPrunhpQvp
hmOprM17L50cOfluIks6wOPBJsHcEWI7PeasjMa5YhORPe2bh7dioblhVfa6
IfU6X/J1aE5rm6z4VyY2ZHh/NRL6veSJxSXBLUZmGq56jkq9oy0VMEThY4AC
3zwxx+KmlMTw3Y0XHZj+Vw9urMBsLPrShAjJ2s0t+eBlIElY9HO9T85QdaWP
1q/q37gxJW9ywLd5T+x8xcg47Y5wQuD36+Tj55CGlsJnc1cndxDGfP8dOrdS
y27UxFFaEDJC/752ta55Fsd9fXf2qShAweu3+fpHVZGtuE1F9BIarcnC16bK
aumDDN3hCgrhJRRSSRgP7gO06Q/G7BqHg0YDKHL2St/DTc0OA5Fz786aNhxK
8f9cRdziqPB+rZ7Pwhxng4mXyy6YnzwrbZwwwhT8yXMiqF3JgthPXjmDBHaV
jB/5EDgXs9kUhw3nTlccVF91QCNxJfAZzPq+VBE37AiqhKX6w7guMuh5aS4G
9BLJjkpbgJDNcs6reFyNywC66r9sCWu/B+1FOci+/s1ccjE9lcAIEjODsAqX
uSAhdowvXcjLAk5Of1Zv/vEb+69jPW8aAgbF3p57kFrAqHRVs6G4Ty5+orfK
jEDx7wNYh6z3u6cWLmrYh7WUxVpnyivJsMBt2sM3AJElfpRY3ZUVi1JSFGxX
oNu0W2mfIS8HnaMPtubi3ty1COp0ArJinlgkehG+Hu+eqyKVv1TBsXcyH1WZ
kEBGmJSwZjontm1jsXiEAibfw3SCTdYOx8825ViKeuNA91g5X9rMzYmeVS75
t0UP8YGIg7vuN1mR8J4pzCYwpxxGWfCyJK8/TSPbQEtsnB9TtwVBhapxv4ur
z27IsdoaiF5uv81O+Y6ioBATkAvWAh8GhH1bUfBux7nPwhbKNxKSsDW0sJd+
d2OY5XeuG45u67pYSU9bDJRkwEyG31BMYqzL0fKGT5OVP745IihdSnFi4y4W
N+EOUxVIA84jM/T6vVl7PAMMraytX2bPZp6e+glu7bcRk1k6K5LcdmSs1p//
sRy/9/C6avCnvWuCzCpx9PW+pTDsbLBkW1d0LdAURKy7rjsWIQLpHycL84Yx
ZXfxxcVjDcPAEEBc/eebjUWQLaEDu2IOoVkrFdEUVOXR97pLyZJhY/jVjJJa
87Z0FxkVd4/Oy+VFi8WA1qnEJ0YrrNKcWZmEV6kP8ERxeu+JUjW/t4uZYAoP
SHEwfHtGdInWifv9Ax4Heeblgk4tuOKNy4wWwZMggln94csQ+idxUXCD4Rei
x1VMSDpTAs9LzpT0jmE8gNa+aA4ATLzwRI+bAatG6MazEllHr6Iddjj+LTpr
L2IppS8n1wGGfQ2Ob2tUi44b1SyU0pE4nJ8yGZiOEZMM9HmHOQ4zjxzg3dv3
2mRXcZWZ4ebOQoFW8ewLun4WadvtUsdmYxesbir6Begbn09RNVtkTabqYXQ+
tMHNfGeCAXQA8Pm218tCv/6gMdNCZ51a/OGS4GTybTI25JVoJjSz9MLKVEa8
sn+YRf0JhqtA7RGWHS3Wv0Q+QWfOHY7bKOr0d3EAIqlI3EEn/98yOjbAzGPa
lQJXik5EfW/YXrywo5kms/VMdp9qFoItY2gdnDFQLmkNmU+5oQdcVt2Wsn17
jUnAn8Tx93KW+ApleQ6VYe6c/4f1Bmby+l3HObjisMZ61sCNgqerQ2fWqtWW
KL9saWbwqGNwzMML5EVFUy/vTcRuA3L2S4R9gu2SfTNB+37DCvyC8Qc77Mvv
scpA81ztihgHvQTqDe3mfFsp7+CyW7OIYQnJTBcfT109ikEEv0gSO6hSg9a3
5lRCQeehgI1PWSEncDa/piT6w7nQwisWCC5LUjl0AJH2ZRJXK0HczJwjyP/j
JDgb254x767W0YZp07z1pmklajJNTkdOOSJiuLkp7v+zGP0rtcREVF2mHZ/G
X494h2UZspTS4Vy8ZjugMaTrQLvI1pEMJrYzR9wOdcb2+yMyBukGXMcL5US9
9fKMVfoWNAFWpXW8eRm8wn8t2r7/4YZY5BAWvqkG4mnNtz3rvwr0hF3AZhz1
KCWVrmDUQ/z67YnH8nJ8UWpAl0hJU84QFYD/tqT29tnYEEhX1mDsmw1pFQNc
PzdvQYKmoBKAy0tUQZO1TxxW5ApHtESvyNgzhRM8lcocVTks6XLMbDSHY27G
0sLqV2bBmxdeR1ZfyE8PigHtJr7L9ppdYzm86DaqkUJth0S18xsx1pPWqv6W
jJyk8VvIucpI1xl9ugI8GqiUARKtnANHgf1F5V2gibNZvMWTT6HiFFNp9SlZ
RZYPLUMNCG71ZInKnxslws6DBrTPbIcJne5vDuTAckoIOhsKkNGXycXqE7CT
JRaB/j8BBW9pCA8GlKwFQGmzor/9NO6bkB7nr1KsiyPDQaeUtueu1KTrX4I1
cXrQw3LOYzy/8VSafeTduq+KG7Vy5PgH093qHjwt5GdQqDmp96tCWZv7uXaL
zEHk/2w+shXs6zc2z6xlhERPxnik9d6siMd2M1l/LNFl1Z65KjtR8WGdXAGW
Y0NtTONODfH2n55qjIdm6mZRKtotmA2ycoljnGNrtnaMuYHZz2BzmuU0j7sH
+ZxMz7ZgCFKa6F74DmixuVZJOyzfNeQDvdbxo0SkCaW2Tn6E8mxnsKSCqBwB
+fGwE7Xs7hOUlZyoQ/P3wjWeWfkZv0aZbpMj3vxGUfNkAO+Wqcbd7+gZQUy3
H1h376FZu0BtqFblUMLliHp/f9QwK1blTysTuyWTJEy4JiFagiMEXMGlJ3FI
RV9ZfpCAOuIk58I+tn51s4PS1LrKFS4sNqauFOmLzuo2E6haImBqTUmvWPoj
HYXUhqZYJF8VHwIrMLLtbBjUpHmT4h0Y92S/+/os90TefzXMPorjLJut3T5/
zy+Phmetf6qnd/PUYGD3jSh5j7N1NnHxeRWYmFM2OwWDz5z29JwhXfnB2LdQ
P7Nq4UaMHEEfToyU/o4su+aXGXuoJg0zqynKCu7pZRiLT4aqYLovrVUbjHvj
EDQQfZgRPa/I3SNm5RCqY1hBErraflqqF1qwEZLTJsKmIwJ2C119332iA97Z
MKtz5zf6uJBfPk6ZpPC9YPp2w+ANYmmYFafzDdOEFncQDslOs7mIkuZQKTXC
+6CuT9E38/tzM2DSsGp1/c4CjKXA3Gc9bA/jap1kqO/E8aV6NvMiRaDPEhB/
/zx4GYSt7ZVLjTbJdGSwqF7kL/0PGKA4HW/JTVi/7Bf+3+NYhkQ6JXBDenve
jYf5EUCTy0Hu60NThIGIQg7thv5FwtAUDhkmsnX7fGfDLJnYFhvm8+AdN9vA
+ZdGo6RMMjE53OOjXHoSNEAbEcHsPnH2tb6zlnkC16w4UMHz0oRWeVMLEy8c
Ysla41YDazTEFXGeNOg9U0ko9VRlJ/JaY1Ipmn64UvIvUAV13ivOi49nfnoE
kT0mooaetTojCq/CB5gBgNWsPu7qgCNJI5ypIFrBRlrmfeLn57C8qFxexRmv
r/8CYAjnl+aDPAVI6gkApr8a5GEax0C/pNCVuw2egRg5w+PnLs7EiiSj+F38
5grzAr8t5iMbQgsMUNezZIfhcIW9Z73hdS1nMIWN/2QGIPt5fwsCNXDtIRZh
jA0YG72IKunKC5FDEW4qjNmPiqbwcew/Z1h14XM9KVXcV+rp6wtYZirQ4y6R
jzaFEElGyZDiCEDY53F2Bcx2GLz9ZITCoCIxQNXEHZ7PfY8zjjYOw/UWbWeE
ZSBrtTLd7b4OikE9ZhgIkGeZWNscGuz5AED4PjK+whppNtsFV8F9ckMo/2JN
G0FWSFIng3ot1s75szin1+ceoQFCEwDCa2ZmNSmiGmk2IvtSuc5XhQdikPrl
2P9EmrIu5oGryZtl7ZXQeFRrYUUvELzci1yD4KZbIOFJ8IXnyZ55f3lbb1h4
hIeQO7bwap0LgAttZBFjWKCxOp5duTLsb2XFXgL/PYvo+//lsNZbS3ccujkU
F7ApeyCF5jzI3E9/2aJdalXomnhlpp0vzLo2qX+42SI13A2BMW7VKPl96XbV
WFQ4YnlD/vtVIuDMhSatCeTw4stSiXFeQibyOvqfiu/aIJz53oUmP8REPKqY
EcVEdQLd1HcEWIJPJqZ+vVof+X9YboNAEYGw8h5JDR7xT1xIg2snRgIS6s0H
HUuQqJmDJwQ8fCNsTIu89CFw43y1e7drZhJwZXlaPHeFDk0JTFCIwdEvz5l9
oo5WjgdWF60mA9LLmHYMUDNs/xGfZvht2vkwDYVEw1qK884vGrH79BGWYLWY
tCxgAWZQ+29DqS3T/ofZMoe40Whzhi9mwp6Ehwy2lvFyYwPAzTi8HruRqUdN
G9pkmQo3A1EXiNokC0pkIrfUq6th1l7dekDANcJmJne47pptk6hId6eYfMYS
1WnzgOvLo7IlUxp6Biw+g/FIJDbXNPZkhYhlQf6YzhtnowRzR4EhinN+sE4b
bcb9/IkBhOhQnRQe5gOX++DQ05dCGS5zLhUHTI+XnDUH9d/5Tc/FDviG0DTm
y+xxMdRfjgTSHDtyvjA1/8RlIa5RGPkOU8hK+6/nywJNDqQXBRPX56r7ZGGe
a9df7CwkMBXRs11aiuMOsaDPId++VQbjfx/kcCTAkkhxCrJUq3dn+zIFS1z7
ENtN2zpnFYoG9XWr7wjnTX+UVD6isbHntXaM4QDwiccNA5izhNXigp8Am2Y5
Xx6togGyJp9SIYKkgnhXgtQiD1Cl7M82QaWVV8jKke97pyGajFEKzX2Fvu0K
rvT+MlPl9gimtgLGN/XYEURRPFwjp9XRoDRhZKGI5oMV4jF6/1QKwXx5xH3F
ZCDti/NmD/YKOor/l/6CR7R/KoYKD93JJKbgdWp/3ICWCzadVR4FciqIQn8c
GqKtsGogNjF8tZcifPqrkuXC5HlGOpvweHtZ4js8FqBOZ3Js/HGTQo+uHoMd
7gX0QwQGocGcD9AzzMfalrL4P+y75mquFHFG8JmB6991knAC83lUZivMhPKc
418vdGc9BfhQ7xYic2Uuua9xl/jS+V4tn/Xt+N5YKx9mPMI94Ywej8kLTTiX
xBnjj7z25FqL//E198pCWjCSvbT9GB/uBRdO4vsoCbRFOj7LaNv6xoM4szXo
Nh1d+FdpY3Da2xah+DW4r18Q1fGeW/OsYsWF/bJJnHGr+iuu7Z4Jld39bgpF
mGBb0uzHIvXDBJA+QXZetse2Vc0Q2oJ2ToMjCxCVM1IWJ3Z31MTVYiYvQPG9
oGlpMRkXUR5YcuI+YRLhLKCGOhwamM2qcO3pQilGznleCrLPNZR3+pRcMtdc
DeB3UfSRKXNVtZMlvF3qYIsh/z8gGb3LVhBbSk+v/YPl9Fy6NkhMUEggAfqR
6FxFxOUjh7CyrdwdPiL5uAF3WmNHtPPHaQ7aiisjeyXSvx1oDCGn3WNqquYz
MnkJtgV5FjRmgXdGhBrCa1cqMwhntsXHPGFpKzKf6EKzoDloOFzBo3mgUFEN
lDJmbaj3nWwnm2UqpW1Txwt2rXp0eXnNLe+FY8xQEkNVf6uUGUKL5vfoV+4G
aGIjVw+tycd2yed6Sad8GxsS2qWCFEa2SY6n5bv/4UFkIZIC6tQVqPxrhSpc
LGr4+mNQjATmdDkKtChwSSF5YNV9VZtCQOWAqPFaTvXw2mk09mpt0e76amiP
a+JnCOEaLFuba2zbWtJvi6TiCK67pC3o2gdBJPPtFMqBaD+fydlmqNfN/bSG
V3MafH4bZwOhbvaXc/KvD0jEHNf9J+xS3cRHhSjHTpbQygufug7SvCeFFtM4
Sl+5j9MKdIKG5wWzhH7jXu/G7SWB0vsFyuimyG4QOaRdddWClWZ31eElH01m
o8A10LCXbX6lWKRAW04H56gLw8hSSM9J14VRuyHdGKMsgC/W2Y0Hm7aD2apJ
UKxRbnHhiEvOrI7767BnP5EgEzod35sO7is7i4Hslu+znjP0dVBfdQw2bdK4
8iHm0Pjce+rQDflewZwuMmrFKdcDcg80wnPXFvrTZsVTLe9izK+hwRUeV2Pa
sLwutV32WdXunF12Iwk7U3lylg2NWub828udk5pI72sze6vpm6XmZDNApFai
ja9uMjs5S0IKLoZFV7vFk7VZ9VkRwVx+fogxCV4/I7RVjvULwCE6aON806ps
LOqlDuEVw/FqN7vPi8ozDHEkM0TfbtBC2IfU+pk28Lbe6AcdqjeFRMrmSmO/
ShaeakWQocTOHFJhtsZD1xXRKRWHBlbGpaXGaCoKB4ZXI6KWqqqYVHURmb9H
M5OpjBl8e7Hf8z69ps/r0HC/Uv3z8hGYpLULWqbW6o303MfbmosecFVnRR/D
+3vg1t3B1GyZeIaiYYuhmW9YUKebPHLKB0xUh3QX7uz2XavbrsgfCoKzUzWT
4paGcw5Fln5whexlbKyADV7oHkm2EjSZEcLpkxjKoE7elhw/4q+YNkHKWOup
PoqTDDe/R1Djv9z4S9ah/AsYapCOk1n0o/b6cz9duyXWQp7nkxxYkezLNSgN
AO62dQaDdCnMFIQdgL/sOly9WA5Dy87vj1zzl/VItBEx8wn5hC6Dbk/ONRe9
EdF+tzblM0j6OIcp0zcTFFa0QkwX/irY2ImYjj5EmysLL8oIT5yQHjaMeCAo
kYw0jBLCOFR+RaoB677xcNQRd/AlBoFaDSxUJcRBGq6I8i9cDQ8c+0FZvKo2
jxIyqW3PKkDiGyKL4sO2OR6Jd1k/DqJda7ptCmd4et1H3+C5gVnK+Dh9wwh6
XDZh5h0vr1Yhw0IbAEj1WiRebmcU6OamZxus+XWOLXNU0A0RT0UZSzjkiiWU
x4L5iHgYKYNbuarJIEGAmlI8bm4eQ6cjc7tgqG7vLvVkAhZzAd/E383PzEIY
axRVTUm/1Zc/SzETeR0cUrIHus4vJloG9xpIDIe3/+OhoFfLkeLni9SLgD89
Wn2DqBdzryiXx81h85pdJklYUkDt8A7f8qmxWD46Hx+NbxW/cI+oFF+vVlMP
nKuI+13ei9i0uRVwmqdj4aWCtasaf/UvtquKiIlTWCMGlAghtPGwJSoauQM1
UhBXwd25V9BGWTGBhLCyAoD4/H1szjMQ39V4bvuOKPwI8iEWdqiKmXNnmLqi
T0os3zO64okPc1XbISqLBPg11vn9lK0sLW6YVR2F06L4CVnpAgM36TlZ11o+
Z7C0T3V4AQuiwKB/MAiH7ni6EbrduAnwwRoOmyX4OWw2Ab4QhUHb0/oVAaRY
W8nTutEUHnFHzAXoUMz6Wc5a7/R5njJK3W7x7mHVlQdeRAMPxukky09j4XFH
V5PsAah/hgIvnLeb8fYg9P3mIGkEAtDAaNy9ndCv1VbF8+PyDtGE40QVsUKh
mzsRiGaVdN/YvuuzVWo0jJxUIubs2wPq7S5Z8KsUWMGcmkRKE8Dso07TUqR/
oujpjtJVdafVSZ9ElMJ8BlDAAg59ZP/CRcTe3Efn5O0N2F8ZlQguL8532U+w
6fD6ZYPYdJppPUwreR3jBAACiJyLQWgtETols+zPGOE0fsr121FzGC8MoWcq
Nm3VPUeExJSV/XubTPm6dSRlBRZ+9tfYwWuzyBxvYmfXqe9y7pziMUNqCNA5
wB/02FTDE9XtbZuyjijbqLIjRgK7uCp27SFL42FEpdNLTr83VSedi0BPK1oI
1yE55Jb+4+801pwAGIbt1BE3AAqtY3JYRY9c86serlMiEcMYE5//sV7hxpIN
0gC04sLxKyrsqr2kdGNGhm/YtiwNn8P6D+bd2avHTE+r7Ldq0zo1a5eitMnq
4z3Gs3OhKqckhIJ/KtkIorg0qZlGsf2PU/jvStcUVP5B6ySlQsY2nCqCSB3i
CyUnklP8RGGDdV+iIW7U1bwghDCALyrDsxw8QCQbrokeH4N0S+xJvsD9fpRv
EBx9KURYU2akl2dHI3qZWzznNX9hbiwQjmIVz47Fg94BkzwFN4CHiFzUoNpD
0rqJyrcoE2CBZIDM3g8e6Q+gA0Iol+Q6mig+TH0B6FlYf9YAM/JJ/RmA8jBX
cMwTaNNrwf2A8+gyN2HF5ze8cLKGqrS99Pg2vDXMsqdiFfeZbTJAf286W5ot
RIiTsoNeiNYG0ZuZZYt2DMMeVIEh9kTLArNL2nlp2X0WTWrFi8jdUSDLGqBy
qEdotY96jtZgn2QZ7lbIQyZypD+QPKYU8MOcKbphjBVOiVhQbbkpTtlXaIRd
xjBvCJdnK8/VXCvBaNlsU2rnEn6hag9P1oyccK9sZ3JkGNniI1Ob8d6f5VOe
wjWIDWlUwN0VFAm+XyVNJo72hus6KPWogncJNthq5NuKsZYDHRv83tDLuW2D
wANFXvqMbQHDAQVSTeWkTOm4GbgMqt8ABV3jiN584g94ZAWHuw4/88xqIWs5
sF5PfPwVftfFXtjdFpYEsjAa5h1/V+DBxvR9+3i0zFzt4PdbLJ5R7hh7hA/u
ipvFL+OTyhgu+7ippND7YjbnKiICj5yug4YBqqJpBhodbWKUjcvb7gMIcwG4
Qr0K5UFc2B0/sxTEbumqi9jVRONZkI0ZB51UvpwPwEIb46AyqoFMOVv+c5KU
RTD5j22G5lMgzO8NgKRYvQFQK7hOmsJ0Z6strxT55CKuwbD6wNhSi22Oo3hv
4c5p7BE0OthF+3MrbHzvvEokmyL58ivi//L0jbRfz+jEhrwKbvbVlcDNERnU
aFbyXGWQmR5MXJfg1TIi05SbUECCceehdZKPsAOFcuJgq5W6tx/zZc+Sbap3
HTedqrBl4/n4mbOn1tCVjzXIPadoZMAnyGl0De2OmBIlgJl26AYitRILU9JU
DYyumU2bAymaSlWU4HnwmM3FtrD0SKml1X23rWvkDbD+8CrJcC8TplsQvvbj
fjc0QcxRC2HSxgiG2gPIBb6e00+Iq+HuOVVgoTiycNVTqFg1sLpAToODywBb
lIFDNEC1eRJqPhtEvy7LWTTCf1ZpJiW6FfYyIAukkG7Ec//0uU1FFC5i9ZHd
CZunjTS+M/4FBiXMyxUisnQ3LgXcbTJrxCwDC7z3SPu+QPdFUgyAgxSqeTp6
t5I4bqkIKP9j5O1yj5ObnQhU9VtZU/5mLJT3k8kR8/YdbMAhn+FmbrRTuBnN
+UKnhQ7Sqfh5gV21vf/p1y45YJbOADFLe08xL+2ASagi/OjvJzfZUGM4dMJn
CmAP5FSje//SwLBTkrI7NuMCqO9uNr8+3y+WiOuygr/iFaFdeRQ8xkGcqwVc
jAgHlBZ7GeWLHQ6Zild13CRxVFMoVTGb5PYWLncI0kNGqVTF+Cd1ZXd0nCre
m88TfMsHvGnI1F8R10rBhlpsAcunHbJ9H2CcjTi1BriuhYJaGAjXtPhCTx4/
fEeqzMfFtSK1PxkpOEBHK/OH11r6hOR6jKJrJS93u4AijSX+kSntRaedeuZ8
iuuz330GnwDND3BIT0W4BWUKWJQ4XFYvQiO+rVEv5rMHh8L1kXFuL8ovzOx+
PWvewZvspemwfHWIE9joWuhZjjlLV6ITnYJdJkZ0I0TDVCys3+ZpBx4SWgPA
4McimsD8BizUPh4S/+pStVpFh/lIynrAJsKc/t3FDXKj8RTfW3+co4HwwOpw
zUeC0Gdz2ZESzksjxd54+uXQG6XDF1kXCfL7BNLVdxkkpaqj9DLAQG7Ezkkj
gf4EhTG4G3H4tGYnMBb+ephwP+R2atP1dpxUJN69RzkMJx9Ge+qhExrm4kRi
TnZP5jJ1IlMuaVA5MB+FkrtXjbXqzsYjOLMa6xRwdvskBO2E720zV/KF6z7y
4aE8aBVmT5vAumCUl66H0RCodKkpGPDtKrWse6CwaKbes2FX6wsH89TngljJ
E7VXv72tH9oQehBLwbwXdLXTRXh6+6LR+HCxicLpdFVjCeYBj+m12nOI0IqC
QCoavHlfBsIt4ZI/GxvPcDmb8pD/uaUnjFTcAa3J8W14h58c/oF1PTidxp98
FFZyUD5ceLKZ7xP4cIBntSCFtOixpFMRobz+3lCT9j7x7hH3vBJft8GA8hHB
/B+YoBZPb0bFQEvXqT0KP2aSE+VgCHs8MAOUh9GAEBIEq9Y0pOP1ve/NA6/B
AmvlBP2edMgJg45qFTIX1zanNmwS+WwZg1sJXLUn/XbQCjgnWgqqKUoauXdQ
OZ/B5CNxyrBq0qGDgS6HtuZy5oonK1RaKu0RLM0pUa4vhe/8KBZLM9KkDo4B
0yY5FTrUWqNPjj/75emip4bXG+P6AvhwYif9qgAo5xEdRe0LuH8zpWv9uwKi
97n52qtd65wf1J8UGCjOfUu1FNHkt5NYHt6ioCB3NXJ7UK5XYlT0WtTPeJEN
RO2x2b68Nc14qest+iADxPpv8xxUmnlfkusuSHiVY7s8L53qtkm1g8SgCxKY
v17odFmKIA9ewJ48ikkKS17NQP2gkDVHuC7TRvkz7OyxfPcLXzWuwfRo++5u
to1bdCiN2W7L+91GWvMD8X9URt5Ud8vwTy4b7IQ13MLDM5wKyrhxcptfWnEf
VsosYQIsgrskRPfFi7IMZfffUwoTK0vtz0q9mm4OYblgaDKcCwedaJBYtoSs
r/BXR2rGeS3iog/uubqQckw4Je3SBOWp+vXjnQXbkXqgn+AOKKv+v5fJGszC
5dLgPpVb17nVnRP3tPvNo/xSJPBAKq2VY+7TGhpQec3DDxu0R05njNO/VH91
QEg5k0eIVWe216WZWqgoIyYBq/2NWKKMxh+oo4maN84uzImPrTu6ocv46ZJh
BNWV6gq2Nt0c2vZYPhKdmHYV5MKvfpRcH7VSwZkPGWtsQZSWM6eQYzeqq9Oc
ohuWtR5Q+8DAAZRB8XG8DrbIkO64uNPnIfSb2wbf+HaWQPW2l0hncBj/pYWC
HGrwv9NY9gqtjcTH1AaKAdMg2IefKnZi8TXHmpQCw+qImq//cHG8KKl/EI2V
aNPmUu66jdX3wut77qZTpfBguNT2ULVVGQySKMxvNEeTbKMsB+JcFe3HfLx9
tCiwcBYSQOUu8Z7sTyCyS1yPFebsBNsg1YwZfIrPHJaMF71i4C77VYdqm/YL
nVE1e/6Br2hKb82KZ/a7sG18/T+slmMy1V27/BXsM/qgIYzHU6Ta/VFuolGU
veTIauny9i/rOVM8kolwgJFDMUoI0qH6VHRTmzHc/LefKe2JUK6ZDY2SpcS0
RPNDwGfIFOBx3tlRISUectucJRh6e8TMiTESzYhLrw8hqA6Psfd2L9cyGG9e
UWAo0pCcof9zFPrs69KrJBbtx61SFYS4+zIOKjHxlvJDA+J8uq2ccT/DUhWx
UQ3gbEylAH2t5l/n55ULfHZEcdGusp/Rna5aXD98AUNVShw4Qb3kAzeB2GSx
tU5gVDEDNzm83K+XhkeuYCYwI3E8ctlFPKC9HcNVqw1OLU0Dz3nR298ycCvx
VF3UzFmn1vI8v588fg4MQmRMN2fiO/RyrREut/xb1vL1e1AaSKoV97Ti6TPK
ukm23wC4pJYG5xBywZd3nA7+mLca3gGwnDFeeODAX8UgBLerP/kXMbR4AnNu
5oFbMCU4O/TqBtwY2Ot2RpQs5YqLzmQ+ri2rJPoN6DlsnQfa6Q9r5mnC54rn
jFzqOM39/7NvcP5qW+Bv5B22mk29kM39m5AUu3AYrsIIyG454B7BewkkADRO
5tO1GU+0UF4rZuYnBy48I9l+uvC+5z0kv8ZcXipW7WOCqaQuUcDxReUw87EG
Hfst3f680uzjaPV7mfO7HBubE31Toa/FLcuXDXLvYbbYdRrIzGkEdIOXx5k3
QEl/sBuRJSzqwfMLbEbPJfarJ95cJuHoS86iRKCVI50phaRxZRLVZNUv+BWV
H3uvI7bQBRKBOiwRmO0Hc1kFfxJwgthccJf8LHqBtFYitFanU4YZrBXve1iO
QHlUSM7FvJ7zmQ0zBynQl74nBu+GbsdTVRbOvx+5RneuL098nYevurtP5oKo
tD6+0FPoG7LA9yA6ALtrB0Tjtc/zM8SKZ+EBYLGdIijqxv/iS9/xQrKgMMGS
aNJf7NdYP5v834ioq6p2GhgiOcg/8zCfJ9BkVrKIcc8PAC74o4kPpFY7ttiZ
iYwqoufmQ/oYRRfXMYd2gNCW++oQ0D7XZnPUy5cji9tJElsr1Ke5UAt8NrO+
yzd5uoyzX/hJzkun1LcsjUYgt11Fhb/OviTkRQyAJyjpJrb63crwTcNIV6DJ
KNpwG7NMIcv2VwELipQrSbHiSfjO97O2ixtbutSdwnPZ+DzG1n6RA60xi73U
XdnSwJSnHhp4gQ0PzWHWwDjuMDjxUdogEgHaR1KMCJCDw7cKl8av1fBkL4eV
udK74V71TT3CURxkWy9VJblrmRB7J3yR3467aeX3iDublUtvdqJelGfhcKVs
15o6hlNnTyazOfEi2uxu7obdQ8QA/1VQVLp/vNF4flpv7PgFMFwE+9feUZU3
2rIBVotBZkitkT/cFm9AZqGJ3QP7xrAWQsxp7nC8VobX/D2Ds9rYZ9Ib8XZQ
fOghmru0ZQT93U4VVtkbw9xyd90+V82jhDzznPgOm8TD/Hw4lN8EAgbwRqao
R/2QVIh+steCe+vsX15U3C06Jk/NZi1Ylk+AKivYlEmv0n1+aNdHCR/TGh2A
RdmCETYyaYE4h1uFmcTqB47abKNXUFDvJ74WeV0IQk7hrZ2sMpTsf3s4/Sie
St44rmZ/F5F8sHhPaMdxX1bAR0xDRl2jsbgAQjWIIR02OpFJ9eTdaVdSn9Jt
4ShVizCPDOaGibixUY3FcAtwhEH2+LwflspcBgvL1zyXzc7PjxYbr6cDFCql
GpK8Rpp3bjxQRmNLwEBCpTxcQIDH50tvIIczr4mggL+ns3Y2LKw1wawgkj0S
HW1HNXnr3lbR4HmoPMsh32+vb/UvuiEJmviQ+WSXIZzlp1TeAsNWFXwZCKKj
sF+3Q8JDfeW14yoZxCJn2e61iH4Z6xL3/QOs8ILiqjD+SNt9s85aLkoUv7jp
t9BNmKO9quU/d6yyAGD9lJSvnUWmGD198t7OGXbKRY2uyPWe+kzmlmLF+Lmo
nPoVkoaGNYDEtbjat5rYP3Mdlx5pUkRzjxRj7TG0Mh3s1pQ7cf1GZK8DZL+J
8Qi9vJ7ZS2tMgstwJSp8SMPhSJAz+3R8gqkESNhRKdzz9YZjTU8R0C6s1bfj
aQnGCfixwq0QwVI734+yN0sz5cxcXVXnI0/IS50Np2FDCwYzERGAaaND4Wiv
m7N4C5gGKWPABfQpaa+xJw6dm1oQYz+tD0uP/eUPQCt3YN2G+zQE/ABhN/Y9
vj/xQAip6xIZfQ/Z1Fah4dNh8lPg/lV8hYzG7SV2Cr696Hl4uKOIA41Rdvcr
C5cpnfP09YNTZgVHQfwGgjnqXAaR8aUn50UCr5DeQNuSACy58zXGbqlgPoRh
uWd9kVqttmmgknbv3d9slODu9obVv2A1ouJqmAPupnuwV3SuizIa6iCYJ4hH
YJH0RLIApEv6pXL5dTDA0pe8n5OAVjlaRbsOSQzRqORko2Nv6oh50ZEHsuA6
23hWh+N6EqkkTzdA7NXGKyHaTl7YAc0aNmmwQXz2lTHAWj6XyN7O2Tl1U3EQ
u80nAwGEQG4xDBaszcfd38KJ22DRtsTu2bjHflnDD4nXp+TcD1kAfkI30rV4
Ed4wOTtciYrjFD1mFT8UO+Z4bYtCJ9dp4dRPIzeRXdwL1VsYCbOMtLh0qibe
YtG/QmSoxquQiUn5ONGi2NZm5gLXLXADXiFcMCMJTuUfA46Lo69Fpr1QtNCo
jWm6X9BOmjHIJyRB841/QEQWK0VvaDKm1ZnXl8ows0adRSAovhdQPkn8V17T
DJrq90VTHin7HFzEWwiLsKEwlJqxE04WoLKztEUVPwxzBR4rg256fIG5MN+A
bxU/akhsVlvQR4wM0Ucy+NtYqRd7G6usF5YpwOQjAgO6iGLes/bczM4eBhf7
s0FDx2TGjGVuH/Paxwewin7CdvFn7B+iMYew+b6nNITuHyvYQEH+iNsbbXX5
Aiqm5JKW99qCK0GCfLICsviGlsvhLzcchcrSSGde6K0Bf5iFiU/gaIS+GVyH
Y1R4dsshRe0/4HtVW2RzhT8fNv6jWDq7oG8EIPgqj04nRoPgySCykUVMIbya
rdgGj+JMsg3vNqYYc7wsSFipms8NzvaRqSV+hDOFTJZWoH9Zkcn+VluXehGr
Ks2f5Cep/cfMagYZUYHMnBApJkB7yfC29Ed/wgjT6p5C7GzGPAOzzaObHde0
NrLRrAT2gJvzzNDNVf4IeslefLw8+tpJ3B+pg8WdKfp3r3bU5YTTWZRtNZ2O
f8zXff/ELWejObvKaeznsdBcjUcs3BLSvcELl/Yxc+BTderJobvmMu7xMM0y
usGwHKP9gFrCw2YavmIPM+HG1SfBxZwM70RUECBltSQZWjBIxxwBABy3boxE
aBBAB2arS2WqsKkvFtwGzWRTFHtD7RE6rNr9i0T9EI0SIx/I7Fns4pIB3TlV
S0+WZbtg1PLB3DnO1zT4uef0CMcXSBFWyZ/rAB2P2i73oOOfhvIcVAgMgZac
yIy0F3au+yuH7u9RVLhpBe0EaVNXDzRSJtV8dQmpG3T0Z9DBAvy2LyJ8iFXj
ed1rANo3YxX0pu69c3jAffdiAxkxlJp4x/PGdm4KSFalGRrkxkg1/dMEFesV
0SKt/MPAh7mQz//S7OFJ5F4TUr3+nbHiTKnA+cDR0Q5hCtA3JwCJ15jwwMsS
wpiPR4G9JixAQTWdvhuNeeOy+A+dFOMfvNW20jXhC1F+0v00w46akO644q7A
lELiocgwCtKTucfXZeFHteaeMGPygOylWO+LPRpud3F4kM+mM0X6MNlCTGor
6QzJAut0FKfBXzKYTLYT+750Bok7jcC8hTro1hlaquuvruV6ITI9VHUG19gF
QIlhprTJYnurvGJZGuA71nx4Qa341IFuTBHF8wgCBxmE0Z0nxKFY+gK9nPEz
okI0DbBGHmgX17DzPGrMH4NBHOVzxGnUTKvAKmTiH2s5076nANvdHwFZr833
KrbujXZvq74JzRw3UbiIVNXBoHZ6JOPyOmMqWhOSQthEyeSXdIpC+v7MTT1W
Crcucy1pnpuk7ItTLhxopwTgQLxNT4uPRQGAjuEUBSakALaNx8Cj355y48cj
bbzgC3DKn9DVkjvQcwP5gqJNajhEk3hZwffZOYkFPwftVrT+HaybBY3AXT/D
8jZ3bF+yAXD/JPVdbNdeFtkAPRy/El6nM3YVkepHciT5MGIx61HBdfiR5a82
p5iEVPbGQiQl1g7gS5MpLKxbO/eHmW/+jxxlhrPn6ZMPkQjMRJEbPGpp/Ru5
H5jQF8yJaf/mgenS+Cgz/c6LaGnTHVq6O1Qiz1Pf+lO8cImmzoeWNT8S+dGr
T4FPbWlR3iPSitXeReNw/WstnLpfx5BT1BV4kH3mtiCqq4QeSk9GFVifznR7
RdAvoJ9l1J34Sf855mAeJrzI3OBT0YRsKXtKov7Ay05ext2f0XSvryQEX0pV
sMdwVjScwNgKveTFda2HFI9ZzI/YP6OtgFgtmcLEXH/scnnlHOqJs9QD5ait
u4iLNbQKp8QCnCVtB+d64RIKW20PpJ2PKzMZf5oJEzrq8M1sWGiOZCahrORp
1E+ltm5r2qYNwZ85hKwC38tRlj3zQZA32xd5cR9FZiyWUGEVT8cn5l7BRq63
LOGIcSDFnJqJKxZGr3IJ4rqF6VOvRBChxmFJHiCe/Dnpc8MlYP3IBnmcVm0E
bk/2ifZuWLu4aPdNOFYouyg2t0+XSlQ6URm+CI4zFeAo19rXQdNUP+TNEjcj
hjGswv4PZtXmGg4eT9ek4n36FXJ5d8sbUk7w3vAFD4Pmt1ZB+iysxfMWvieY
8xr8dBzT5PGaX8dcFZGZ3gxkBEK8CunvycehLhkp3HcD56/WDdvuFjLM1fAA
C7/71+eEhklELdakjEKazLh9ady98/XQb1I7SN8Od8RLOGi5QhVr83u0CNoh
h7XcM7pLy0T18cEC2RbS3jsn0DKZp+3nGA8x0te20k3dLGFm/f5jaxU8viGh
Jgm24IEb6aIrp9fe9a4DR4wfScGYLkG5SKdIKUvXO87T2nZuxFbS+NEctmty
/MZohWPgW/i311JA7DeJ46RqNYJxYvjlwAVugxz5Ex9foA5YK7wDSkNTIkkX
8o6ChPMA3lXM1j879/8FmojY3rstkWe+48jgR0fsQr7w0/vwWIAFh994KlK3
eoszFHNnDsqIJx5edrOuwxyY7I53J4KO21HX4yxF6ufG9kq94elKUCSGSLQP
FsyZFHQlJ4FmusEcQy9uW4+2Vwwt1e4BSFIt1YGxIqk9jpYh+cUMZ35u7zTF
ypB7fBsyrdeaccdREODMJdTLHYAUH+p1+Ls5JZH7i5V/uazkE56RFlUtvDCp
yDH/pZSFtppnBSUqZyU+etf+k93b3mhpo//x51W6xTLMVacv4vy3yKhTamTh
09JWk+g3r96gzDP6R28tR/l4ULphrLOl4LTxXTlkAccyDNYcO/f83qH9vA3P
phGNuYZsfbfg3UHly9Syyz+SMOpGTI+O+lLdZl1WCbG9LwbX2PPunSz8+AAW
wFbz9H74jzg+EFhVcpJo8QciI9g52NQN9stQ0Lsk8p6VWV528IWR6KPW763q
9NfjhvuMUTchiBQPFHrEc/xxCKW1sP8tDx2sOeHZtiyDj8I//0YD7ZUQ+nJJ
Yxi1EW6PkST5PdfPWfZnZ5wzEYvH/BTE5wTONJAbGbTpcWBk3gJ9QujrVQ3k
we6pXwyCQz7x4Nmr1fC0b6M4kcKgPOd685N2C6rQHvp7v40Od6mnmJM/8p6R
d37kv1Lhd6cxO9UFjPvFZFmqZOHbRUWfCueoQEo+ZroHk98ajKwiZHm5vIse
5xG/rp+gGIJ+8Cy2EBrjjqALygilyxWTxatmj1EAwJiCBNQToEdXkGljnVmd
jkRo13aemFw3YfY2miIEkZ0PaWorBiK0ykNG2V4bIkK27s+Ek9WBiNM7jMST
ULMyM3jRnkbaV4MhnUa+PW1fLD7Mz6S3OWI0aNR/+W3pRdxaV2wHBivB4iAd
S/TfDwZM6afuR7FMtsF5+gOT4g1/Qela4gSU944Hc+FxkA+/Me477GTZFGBT
WkgACVl8ZCafh3C/7YMM4xZ/Jt2p7vXseo7NeZMuZ28U39cKCoVD11CmJwm7
uzcs819tNGYs2JEFSsiDOI/XphLydddVdDR0UvQjaqWea5j9fQB0Vsd0KzSd
TCEmMIotqcp5G1o/LBKQW355OOi6P0m6ue7j24iTCs+3lpBt11MgRAeKtxW0
XimS7r66jNQjGvoyiyzEMdbzBGa4ycUhVOrka8+hPapUDVq18PJ0lNCrhiBm
PbL15NlLHyYid4l0Q2fIRVfPvB4Q68z168iJdi3nJHfHHokgR/9RriCciaE6
lPu7MNq3UbGGAKnebFKRRIc/v/2N9k9jVTiM0b93UQbtp7dzdfQWfM2V/LgK
7ORZUk1waWi/AKrWgfEQCGKkW+NJE05F49nnO0ZRq8D7oz/hDtvMbULiBh2L
tfzqPk9rrN2PQ55vQ6z0ew5wwh7cYzvWGZ98JceD/qe8DEbyjpZgmpGwF0ea
cwAR/LDi1/3Jf19e4E5s5qGxKq0b4zyacBqqewuEKYtO+MeC9ozPgHS3Hft0
w0MA9WZ1PTjh05yZ+Fcz0umVaL75BwPTsnoz2TXIp6FedVaAOaIr+KEBDHNV
5CPj+q7A/SIElF9vVeu5YPJDrz+B8ZzVwzcaPigTrVNPDl9jm5lVhhPpHqMj
T9S3kqmhQKL1xU0L+7VDtphX0Nk8MyOrYpORF2KuNSJU3FOTua4Fh0pmO9JJ
nZ+fSt50PHfnBNbVy2rfDpBt0BvDDgaZV1XP9er58jIy2WCBZBBq4NZ6oDIp
wBP9W/eD1y6IW8jPzpq9m0XQRKx7I7+Br+9IhD7NfxCXcF5mdIgKa+0xTcXm
jtMYp07oH59+sfGra0JChoAbtirRpQmj36FQhqKHb8X6gDuFOU2sz6kVp7go
Hd37pPJc+gtDgLR4qMer8T8YK7snCgwB67lRPz79CAzYwpgui39MxWkGr0gO
iPOTtdMbM2Ows8W7YpDYnPyE2M4xczTYEOwuECTmsflRrnMllSoxfyIUqTxU
tJ535eflbVQJNHDJwh7malmMZTMig7F9imYwwxXJagk6Dgw6z/R8YrjMpDKq
Ur2LzJkC9LNFy9WUK53v+ARZR8jBJJnbOcjZtoGAdbH7Fvsg7U5F+lLdJTU0
Q2xi9MdVEAKR+Nm/g/PJ68W0GQqq+6J4i5DSS1wSVyTXSWv1WA5E2+MS68HD
Uqsq2Fzm0gmwjcO6sqTI7TwX0TDbPHTZ5/NAfzo1PiChjkdXYb4h5JJ2LLGg
LkOKk7CjtoqYPHU62AB6gb1IInM8FeThG0+8N4GOyEJ9sCtEL2yTxaFq80hX
6UN8nKYHzKipOIzokkk0OvxCvPj7iagsUteb2j/mkCICMkbpGrdu3s4eHbg9
wzsLBCekYsnURERlr3LWkTXPXePHQAP2cXc6RzMgxlNDjl/22KFwZ0p6ewXp
9shfC5YF4MxuEyCAVzFS7XUXPFwSkCfvujMJ9q0w2SrWl+fZg1mGdUMnDnEM
VoHi9FQMCc9NUMwiaRWmvfcF/SE07fY3gvcF30oCSZKGw/bKFZMXxH70afa0
A0AC29TMRzk+BmM8E/KSiImAcF2wrTQ1DhNPNhd1/V3KPA65z9kTyckj9kgO
nBmift0ctQucV/RBe0gWUV/8qqMCtnh3sUE63DXNn0nHuU49Y2SzXnSeqhf0
eyPwmzaK4duTayFm4j5tWqpmQqBG2bo9ptpD7hLxRdQy7Kk9X9kxl38m/YNE
hWLgjaW0JtANP4rPXHlJDnaQPzIGvNMPro1eml7JWQCfJdy4BykhS9GlicNn
jlPTws3xF3od6ZRNP+930boNToIliMpF3Y+PYHvN45FzLhqsQn3WyDQfTSA0
zXEMFcM1pZxiFOH+cRNRYnMiRJXAFhCh4yG3MZVbpyEs45hUICwQcJdyu6QV
hly0y3sS2utKHV6JehBvrcrBy0v4KLwx+9KB0dDEyU2gMZmFgru3gsdVj7JB
sJSMSHTQVbMCaX3ThJe7fJSwtllXACWD9fhZ84gBaWxC7AAzEWQtk5micjBn
mYdv4d/3FB7T/Jbyuzs8bpYQf0n5zrCAtqAAY4nJe5TTrMFar5DvWRATPRKB
yMuhGihYF02ZXNM4tbNF5IQZF1w12BX5Xs9QFLemsLZlwmF1a1ae/JVHJVYp
JgBJirtZmwN9AsC/kpHMvrMHzmM9J4ZbuHXThywISdK6/S2G029GMf/8fWpI
0mEIfJGqwl8DyfL2G0jo4CRHA9nbC36DC2F8E14HIeP+D4cVSDrN5pKouw5O
ulY2FMQ9PLBu4K+OFTURipk/6lMrCRD3/LNUm2oxtUJFTEKZTR8YBvB9pCZK
yjwSJgwwixRhPl+8i+Q8f3xib6+d4LD4D+2yALYfV4LlA/cG00zC4d5i6fOg
EJkPrhxL9Fy++HHXKgRHWDtZJpRfK6q1r6cT+/K5nM1L4X0EkrKNXSkby1so
0HJ7BdJZZEGFEBM1Xh1Di1+MrDgeRdeFhHKFVHggf76I5Xoodkiqfs5D7SB5
Xsa4qg26zdHfKHwaPLdM0pWFv6fdazmLXEFqOhxyakozM+Wurxu84+zknqup
7zE5SBH8ECND6kHr+jJz2mcpvLRlWOvMdUtcmy54zMkKaKMoNcMocHvuCESn
7GOpgMwp8vpsiM5uQ5J+pt6Zsx5ccubh9AbZV8cUQhSuUygfNbQJaM2D371T
/OOfEaC7eQ5vxS5lKZj/4+8Yp6xr046zkIyeMZcTF/QjeHP+3CbmaJkosV18
SLRfK+PSMLLMWBUPyDvpUVZpYBlCftj5rVsWadEcTn7icIs0cVQ8rmBou4Dy
l8LsFGj0wNSD1MUlf86s6h18rJ/Xld4DXm10YU84XrKjGtNZ+qq2RfGpF4Zu
nRCEcgAkciWXp2m7dmWNROF9DXOMDu72M2wOPF0afxkriTrWQEAYOniKRRQO
eOIOQoHlUJLzYwy/Gdqc5C9LBgtB7YW3swIoihXemZY/4XDJN678ogRvnR99
71dL3mCJHoWRKzPDwlRPPP3W+N0lPqXspG14BjJ/MwqQYYXf73+7jbzL0Vtv
NJ+sVuSryqm32h4AuxVDCsp9TWG1RZLhUrAssbOdOBBHN23VlaTIIHF1BbLW
RvRlDcvjmDf/XP8RZ/Kd1SMI/L17QXDkT08AJ2BXvWP0yMD6fg3ghimzR2BX
QGBxgu5E1p3X8erhC+E/mXF4xcTE+0aY/U4JYJuDblCQ4OqXG3QydwthA4GE
X+pLkoahyktEPNw5wg8n0vGeHzwbfKubyzC7LIFpS7u63OcJphNjAYea1Ygd
aEgMDRGfb5SWK0yuSvCdqLlLp58KekgYZ8f3uFHDcqLj3vihWD8I1Pg+THT1
XshnDU/i7nOWTTe9M/dVoqT6b2sUnAtNPcVl63ANWIN2nEUxgkh0PJGLy5ew
awDvFf5Y4Ug8060ldTfngy6ZgrZ7ctEdvwWd7r3JteB3mDpQxCKRvYRuErbn
mez2D0HCMF6x6JweIyXuskDIlGk+lcOn1eJLWx5PoBE6H67VE8fWXcMcGKpr
00GfyQn37waxM3vL79Ccuhkp971NzM9BeWjy9ACSU6nuDY+ucnig0gso59Ue
oOa+pvBuooRfH71k6ki1/lu/YOJRX73VSIYSr524I+wa4qkJTmtlTu7hEY0X
lhP2hS6P2HV+/KMT0SJ8+2wF2EzZM4X3GwFTPEpl1hWl4JZu+Pc87uSo0n3j
9f98D1jCxLVjzJdMi3vLVPAc8GD4PdpVC3lZOHfmrx9HsW3mlS+5HBGPUOQV
cej98RGCPpW/K5y1WW9fd4coi26nTGkLPUHdcm/+zIvR0ZFPM72t6WYzTZWq
TqDkARZKhJN3o8lCQlBcXSm9KCqEBCALT9go55J74vuzPZgu8Y+KQaeA5bte
A7rQ/IQzL9qtv0YOo6qz5OzI7daiFU57r5D12yTIXopGTewaf9EP+hZCxYJq
AAZdj6lUxZrOqUtlgzjUVipROKBSVyGEfvq/vxAtoI9WC+LpJo4r5yFhlCST
hNXO8lATpJdOCN476EGiiJpev1YGdfKcZGC8s7vnBYXxOEGvBGF2V9Z3tZth
EMInN203L99Dh/vbX1byaYzv4LAeGeYpciAVOQhD82r93bjNb5CF0zi97TH6
EkxmCZfnCkais1+R5kQ2s3T7Qwrd4J7MCUp38+uZyOp21l73wWunVjPScAIE
E+sLJjU6Aim2Xb5XQmqud+DDi5/6emU2uyVpFi1D6S5XuXvP6FL7nQFpkLyY
kkUR8PdH50xsHITQsxEWcnJrb4+T4RmMjxZBPZLBueTBKqZG5sbk+MaFc8OK
FIPvMVC9CQF/VgGbuz8F/LtFmo0L0KLsBnw2hRoUnUBIpFCYoS7CNZY3Zude
zyesTKbiDCjllv6/D5Erz53uU91FKWO3b17oX0GbzJxdzY9az2DhTMbvehNo
+w396z8VbUo0ft4hOGmlpHMpdw2PS1pR2TJxs+F0EAvbNnB9wecH/mIAI4ZR
bgNlcfr1SGJGkOdxyKSg9Mw4fM9M1ttG/RvbwKjlzMUxuJzMKsf4wiRwANfL
/wfLZ8Oc3+3ZUm+cFHdbwSjPW3JpbiX7NIIskzisJwNoi7odX+XLCkVlNrvU
2uVVj7oHWAKlo20tve/RJAac9u/8MAdCDK+8YobkLFdHfExvm02JDo+jajVX
ThLWe0MPf0pRTd/OPRvUayBPY6nk869q2RbXTyxTN2dfgg2FfeVfJC221okB
a1AgseBINELHKlonMqV9nBza7rbCMC5333YGVLtWGTUllOFiZQKu4If+z50k
MTetUVsZAWKrJcHvuy86yxWfWCeGLDcOCza1nAK3ZwlIpoqUIN6f/831aQ4T
KTullaRhyQnhXZgZJV9ziYMm+uW2BZCEK1yBIlTcUq8dSolFnWT5fRtkZUxu
cHPLxz2zsZUBxfnU7A0fkk330wwBD1c4i+Gr7MeZJsbdZyICmpETZcaq2g6u
2xO7odV518sXv2YYZLibDKMjI+XlGkVWJ0frGicoE9pEAkuNgF5PRH2l/DaY
F+6HEYtL4kY0Oopvu8MyUBD0v0+/D9jrRxHZr4gCuC50Unqy1uVrDeHe1Fjm
cU141VXhSqROe7Y3yks6m4f6sd1fUw5Admn+yXk2z8mbP1rW2RQ25fi/uNls
pGUEdLnap/dYCFQbSqbfL5mOm73qIVAy7icw/q6UknmvBDHfZryGuneLmXi+
ZmSy898m15OpS1Qqdyq4BF1jEmGUe4urX4RaqBBTuuVHSCAhuui1gmI+reSC
Q9pLPHnsZZOy7Ozc0Y5e4j0JXovXcoIkCtCjk6HfpDI7Gd4c7jOk/t1YuozO
O9Jwk6jKTkYBZvvUyGzZQb8r76DSCzL9aZQTe5H4GS32J/7gdbiAG04h+Ic2
1+V+cdYr4vjHu/DTmxSM5ASIPI47twQyNiCklrGq2aMYC99meYAhH+FeY9Y0
QMsryJ+kCDpsXJ9+/Do20JbZoQu4YCyFRCXS5MkfVEFfYuZuEs96vbOrPsHa
CFowUmmtPo9HCynFjQXD/wx2ghkPQxKLuIZjhBh5J5pYkOR6L7ozQnHG3WY3
hip/W6jI6zaqFb5QLmSpHmM3NAatoIqDmPSutldMLNMM/5nC+8iKik+YhFnD
1yB9ubyfwzVhfxtD/G0IipcY85B9eu+P3S8isVMK7OpEnql0VTmwimgwxqxa
3uOEJ5HCE6tzgmnB00s0rc2CY16mhl+56+yA+g0cWjPFBbX8HEpolSJNqYFU
VapPWbwXXLpI+iovixpEnAwX+YTyIhYXd070Pc57PhYoYKk1sMigMiYe9VTV
lyJRCKuOcL0HyANSm4DBaW0JC4V47ZUdURBXFmx6fydiXiyXCo3srsz0EEAS
jh5ztLop03fxZu3PeUlto1YokeCrJlbgts+TSTKLA2aPxtRBYBh6D7251akl
I1hacz06pKU0imJzEj9Xrg6cIeao4gHjPmqXVRc/r2FsMhBUsp8zIVf0u70U
jeKuSA/Cad80A4wbdivQrRvpdJR+/wa7J2ZTKH/KLnOm/msTxPUUfyyS8iTd
AasMH13JDGokP750FoY9CWqVX6XbFvS+SPBoPggqWUaIzA+t5/ZGduQ3m1c1
MxKLd3DkRl9UunhCW9MF6SZ+b5rQ9pHr8CfMy6pMFBJECgYOPQR77I8UFdtf
OwWuHXA6a5WIzoEfxO4e3SJIAwOr78gdcRA297ibw+yrhhCGetXCCAKySRcI
q45HQkdpYOZilCJeg2t/DcgCVHk5Q9kTO0zQIkHXUIFSluZb6Ad8rAHYoGRW
5A/JzAJVgF63W9vDpKig0M3HdBumgozfcQMn/8ZLhcUpmSuWTpX3u0osPuIS
LZFZYgVU+J9rAkHAu4YolEOcWKt3IiQUWcvYns/sER8niHWIqjI9DtswrOPK
xEyjgsVnKyAUdGApS3lZ5fMIl1AlT6G+aSZ5E2UPb3o4KxKwbPvvP7+frSz2
na25NPTrjMG/Ytp/wg0UmNt/YFq9B23Sd9ouqh6IK1c4GEYYMwADC6hLyyyd
aVnVTdvlh9PRW2Yn3lnXBIjpHDCRyeUlFc/Rk/0VCJ06C9QrztNczbQ+ep4t
XqSMfRgkly+JZnhO+2hiDsnMf7fcR4yWtYttS7/5VhhMpJZDJIdKlGwsOh1Z
b6Po5A4Th8SJaLr26RJQjNDrypLj8UilusyeJ7mrFo1lxE9Du6DU4ysJgMjQ
znsSsmwkpjt0uekzrCJwNnibxMF4BjkzKHHtYELMK5ktqFElc4qvQfS5XIDH
kgqqiYpc2pER3f28KDa+o+juKCg9UlT6QrLAadPQynnoMUhacWzIa7WykCg+
J5nH91hctIVzYY7pq4412eT3eI1bjv45Ht6qhOAxKacHTB42sEVzNw+bma0q
aa+7U4OYQ+i9k1OOlvaDDBfA22Y6KhyFNxcm9eft/fzMf3g1CxTwUfMyWcrh
SiSRM+7jlzYM0Oqh0U3CiBW7/d3x+ej6ULlnasQBS21BXr26MmY/zVJwIb8W
pClRmxFlBz139xLAEc3OeikQlXntVt8ly2JP85N1tu4pFK4sN3vHowjAGOH2
uqHcMwSWd8fQSKCyhXT1lTA1P1/A16VYpkqT7YqUTY3axQS6Vc8WrqZpJ3xd
s44I5h/WDrYXNzOApRkH3eYr9yLKOh2kUFKbq9EErxItdUgVg72LiRCxMZge
iBjSroHk8tNXpHan7zGJIjdNdyv1MccWpSyElpP1k3ujNKouNyil7BX8Z22Z
3KvJUiuBqGeg87QGfcJKohuGjVQA1KbgA59bh1G0LUUGVnC/OlMW61UqZjGH
7KuH5rpiWUM7KoJMnOGcGHkANJ2vcn0U47Yv1trL0DHbB0VqxFmMDQuVKvN/
xxVEpY5RLqXW01l3+ovKQRyLLMk4tD7Jv1KFS338ows/wjsly0EeC2InutZH
9Ra9o54BAcXdrRealWQPwTdsq1WEDP/lkuZla1yxuxi1hKg5tFaRCcrut5qV
DNSKU98SGy4RiUFlJ6K7dp7ZUzLsxgaGQrf0kwlAtyuK+P4JYr3Z44FJVqBm
ktm0Zov/gdJpKywxNYVVgjj3RicgahBAm96PKt5oSEKNYp0DiZstZf24ighQ
XPLGOgzb//OoZ+CbsHtVzKT1Li5EoYL9EgS3mnO+txY7TVBVItO4I2Q+Ucnb
eC0ZUQSYjfJaW7Y982feeSLjDbKC/tTx5+I+E8PEXdz0+6lN2P0qEYTFXFsb
IXc5o8zifPAvriLRJndc2uxBufB/PElxlA72dIObJOFFRz8DeCa0g12JcEaf
/76EsBA+hO4P+DFq6RQUjYfrWF1QvTzpQcHg9rAemHaAX0SagRLMPFWDFJC5
UjPnKqturqRNuYsxLmwXrwk/T6q50L34cnC3Nz3fHwAHKqY56+obWYVyboBb
mI+GZwj0oCCkLAWGWrybkn30zWTASk/np17khrZhC70wIR6b1CWx4NLKITwv
SCrKRNXHzNnPQtHEHqoBXY7lQFSvX6/TU+d9x0LNpKyZLW9VJ7h8voNrYc4U
DicWj0eIMPXqD7AcwpWQ56LBOQ38qA8oCbduyXhhPRJWCj7Rcoyqs1wY34SF
XScs+8L/YJVsVKM5Yij0hGBH6iGPL6uZ7oDiTET5Lc2++C33+0hPzeMryRgP
fRdp03UMnNhoB3Qb7o5/BT8mcZGx+hThJrxBRzztQhxAkqVaWzQWKf1fiPl1
hCXFQB6aBtHBcmhNyH5nxkVTg1nlYUwtIsbYh4+KxLF8CwKdVQLSrUQQBoWm
M8lL581GlwXgLVzXjSDhGo46iY3UZRcKDSo462UdTdt4VqZ5MtVUbJI+WxTk
RlQg7LCT4ZFdtkNJVbV/IFzx69HsG0tO6ML16MKiaMJaEQveJOSkgIjvC3dv
HOreR+TDecrVi3e+TRTi8CDA7gLl5IM1zrKu6NzV/GWPV6cidgE8SbCsRZmB
1MRY3SHam7xZ/R/uos0mzP7bDHuU5g13GI4GwZtkpm5dbAnA+jDkAnTZCo2C
6NV68lwF+IezEUlImK0JaTw0FSXR1KrarFVaMv3D3QtFqtKtd0liHd+RO/9f
yqSy9H/KFgWpONjet6mGtJ0VSCRqS65sWl0fwpJ9sa9T9EJoW9pekC/hLp5V
p/UB5s0v0J6T3MhFN1/93s9V9DPXOq3cI6QpI+HwMZJqTP9hiu89dhKBnNVO
NSM8T6chf4tn9Fjo7UlYPkVH/SIy98HkaSOZWVuwBbj0pyAVeG6+0AePb4JJ
hVieZoJ/ddpOEhTyMpbewBwLnWIusFW6C9FDQ+azqVsKXh4Rst8kT2mvOGiN
Nb/1N+i4k1ZX0GQFaB4PYE+1dHzinyjmIrGcP5BIuQAAvIyjVjsbrgTh0/bw
l2M3bQHzdNXY/5sYP3Zy5IP8aALzL43cCtDg4A0+cfTvwVHTr6IzoT2NMJJA
0ccylCYoi2GhTFc8LPxzfWkdWRALkkgg93DeZ5CQTt/HJN6P4uFZkb3T8Rpc
8yenm4un45j68Pa+ZYA1ITfs3xdBI280lU5GUf8TUx+BeJW/JfnARccNecKp
48P8+S8HrqIRfAkb3Uy8mrw/mAOGsA3fCasx0HntumR7ph34zd8FbVxy6JUA
tJToNmFgFi/1IrpP3P3jF9NUxGuRfUSEcbidv0EjvFADGOPycSPlP4nU7MOw
ZwWO9YkNQCmqZWRdfj98SYzxOvbFzQ/Ewusqg8x345gHAI49QG7vHTmGKrvK
nm+thWSfQqZfahfeRocwmhV6IY6/IfDGg3WV/VMginwMfSmuLc3vmu7RMsAC
J8/CiHQwvT9M/3OEta7TiAWQRdPe1tYvF3f166GE21ac1YgNDtiT7VYA4daI
gI01xY1F8pWAIciARLF7wwSqnH1J84TztLtAAvp3odsF4HmlqqJpWXVrM7lu
kyD/WlEOHc16l/vs/VT/zowKY6Xp1IR2NnvCE05Z9hMCUB5h06QgAlVujRQ/
7ZFvD6sIEbijnZRNnELeaQzPhvaYDGh912AnpfrYHUnCV2380nTsV908JCLn
xBstQsPHsCiWuBDrHincrAOpN54aMN5Bgz1aMqxktiEa//78w3zUntxUlphD
Ehl4hzk8MWPV2/SkxnHnF1Yl/iQ9AqlWhfEPTKWxdsqkA3bZ3RCkLiwuqCAu
EY1a8ZVCEoxW8llDGdjnr+ktV4TnurhHIdwtYtVr6Aw58A5Nxix7tLZYqj0g
e4F+VfFFj4QlEEtEymegUwDZv2iyrZaEUiB0yvGgFpoFTcvQ+2K37gmO5JTZ
0FauKC7hZuilfzEknGBuQVfJo+/2L+EV7kCLhAXSe31iIl4L+1ZY1nOOjnyd
hOt3aTdCBY0roXzGN7/ehHn/qXvYDGTL7usRdjiSn9OE6FKLAI9+9C0AJH8j
egBqq9CoHKe2RfGDC6fpr3uLrYknIPj1MakYs05+MzmM8ZRveHekte8aABKw
PrHEMOTlwLGG/R2495FKQ1thUfSI5Q+W2lriFpocFUkNgnFJ9kP5tt1WO2HJ
eoHai1S6+ctdaRKpQYvHJ9s91fRP5AIkXcoDuTS4hH2XFeXAZgn+69b7b6yP
myGdM+TMhyIYJZytFktCGC1Jte9dihfEedmz+uNW5D0ZyLAnyniyCTZzvfvE
yQTRdlEhSalZ4byf8wlcs9Og5GuFyvQ+0ZL1r9km17GlYtYZsM1Y1syzC8Ze
+DGQUGEw9yOeJC16suz3wChZW8tAa1rx0xornFGb9VkKigcVKR2WMgrMdspT
EXNbacTo8YUmToWzrblmiWdRHUYXWDHIsM1tWDbrWonm70G7IVJhRm/lDUIU
Reo2+M0CPeIgJjMh14sJbqNbD/ZQrBnq/Pi7Eu/oV7HJ0fhFNY6A3QVCQ+RW
ri3iUMxEALWaA01bcKPvEe5PfaO6KrC86w5/ov/e4jKLjDa1lsDAv1iW0rAo
FkqGJvyHYq0+K0Vtu4hF6ttMsrkb9awx7MRo33fWgUqmyaHIDNNvd8HKuEn5
dagy2eyd8EGneVJrVEdpiMR5MjZYCuX63nYRsv61CEgQFF1rFe709Cpl4u0O
cmCKqzridJQTSm5uiKoOlZ9/UDXGqQdgohs+dBT1xIQFzn13foO3XFstrPvZ
m3CJcEmtKlQ0w0OHJNrQPNcWAJ2xbKzu7ggSF1S36pNsvmMOFTNuu07mxgv+
zWN3qbIfdlwgdBMfCQix6vqip7an/b/PAlMfM0amkzJ372PbHYPrnLa6T9i9
G0GcOjbUkH2Yp+AR/scywPSfw2fkA/k2uuLc1dETH8T0MAd0pqT2XyUwbfl9
Ciwow7lbz6KKdjUkS9qaR9s5g5Hin9DRRjCkbB7S1sa8b7mgLoHl2YrFZJZf
s0vyUUofUbhW+dBkIZDj+eiOl2msF3chCD0e0ZCp6jM7spj7tfGynXcnnWQ8
VWmMBlPjiVX8un88Fkv/FCt4upBBy+ykwkELCf6LUCjdyLTCiVzURdNhPFIa
OUOgkbCDyA8uLsx4E1uV4yMLPGZWsyWy9i8oAUSIdwwhRpFr6LdVB6lSAaSs
2Nj1RwpSNdpW4WN6Pwq/m7w/dGhsQPtrQFd7fIIKIkZAyOiwNAzexapKMITL
nGgvywehbaoawbQvhE0udWZIpib1LYns7T4lWOz7LAnnojpehxM91d6OTof7
U+K5en15/90Br5J2witLRcN8LtBEw++ySL4R1eDPbiPQY3QetukpDbLxR0j4
LA7m+06PjEx/aVYVo3hGdVeVA/yXy0TK4SoTc3wnvfg5sepgEmplkOpWu/Gw
b+W2ZCS3lhLF01/rLQbH5qKlcdKj7jqX6/2Eh3+UYzu2nJxehaeoZ6U9a8EJ
hVWE97SvYE2wUeAZ/L3HqsJghtPX8nCEfwPIwLwrUq4ewgD9EgivVmOJqNT4
KiaBrj3dRp1rwdMGHLOwq0T5t494bU+J/Q4Eofi65fd2e/RgQaRdLKI+PSo6
A5tWQyig6ILx9Vo6CaDULOo07ZwNN/7FqV1KAjqiMTsbsxJwAIZdCSkFWhlD
PDTfLYtsKfJ4vYPz7SrCTHqAlBm6xhWRi0EKRoi1wZj4JmiG1qPhYVyEmDCi
kMW3YqjigttTxyzhRqIyuC8OJsPdO/dURlrKpsue+uN0PIsIJW52PBzNl1tr
vAM9nHhTmMsjz3tW8yggC7O2CdlZQnstPgD7OyizXTHeQ6QYksxniVas67on
FmZRzrrH1EhpJJb8LejEj5ptOgtdMb+fpZoXw9VsBtlfWBe3iJOv+EP+ntKT
c/nRlvwFrUMEJEaoPDlHAaGbMDNHm5Zf2p+GGb2Xteuo2shPrWXTw2/TCZrt
dpaJGm6YmACOBlEUynXyp3k/zI3j1xA7h5rK4MZPo3lhJNZXJ2OMcsZ1QJbt
BJsEoIZiOscVo3Q1nc6v8xs4/u1RSYT8KVpPhFxRs3yndZTco/xWMznQQWxX
OgNUoG+vImWeG7m/APhmWqmc5LkAL46QaOmny2JgWjGmFaEzQiGPKTSHJHuU
yv3XO0FXVPWsWuRawDuiyAjv4fItZvUYO/WH+hS6mtfKAGGAPLbrg8Z10A2o
eHtO51aVCTSz72ETGqK9frHTCn0O6vVOVGRgBDNbMWCY81fAQdvPh4Te1nIV
3JCo17TtVGH1NhHi++Z5bGIuFQfCfQruwhPkR3s8zMTjDcz5ShpWZSyfspbi
gi6Iy8gBfSiFA9nyihPg395DBy4DTEVOerdqEJYrj+9QXTzbKqUwn29yTshL
dUaMSyMXOAuMRTnbouz+dAwOi3p2rraSHbM4CaokJICrcU3R1qshmmaQxX+A
Jk6lK1AElP+2fmfbeevJNXh277HwigL6wWjXLFgOE9FOAdB81/F8qhEuVpsh
jicxDV9dkJZDM6C8BSxuH7k9uDVmMXWNXORIEhsJ/FtQGLP97vqNBZ3ZNDYj
55RloMbXponOy5mbcZa2I96qXp0Qqp5/63Uk6gpSE9Wu32FmCidXvQz7aUjr
U2zplxfSRQhFyJpCPyCUah3/AkAq7L38HcSSiNQaBPUswpGmYKpv84xn7Xv5
RF/nuSdM0b40RiITT5cMQLUOWpIip72jPVrzMzoYR2yOci/vJs82fLBPhmNn
q4bTsT1ENfEtikXI1vrNbm6u9KkhyC0zXsJadPlX7SOTMgGki2HZIulDNkD3
ai4Hr0LqV+FU4hlbOTPB3/z6mAOm/2NtTS4IjqUOFBRAUOzPwRo4eqVPokEe
oLj982uzOVlKkN5a0lFwGh2sQi1tJaVmbIDXAynVBOQrQ1dKDMPfcOt6L8jb
y6ra54y/qV8FRIznH7nxwzfpx7xGKToYddylpN30Qkxnxrp/UTIBTQ3uUD2h
3CSbVDIcsZPi0YxZ1MZRA+xf+cXPxUKilSrQ8Ngz5Jg7ICRGY67Pc+URwaoE
wkz0hB3oAB4jeGRsY4eS/DFniwbYHJ+TEPKF6q5p6wqrXq36S9TuTJ8vIeyT
P7sSNtWE7eOhqwUMf2TqWgFlsrAG1bbNmemdjVI3fjHpuDmPXVeNBB+dQrI8
0+w+VsnIxAl94MsZ6xk6SHtpesv9bxt3g+WZHzh9JuJEquGsKb+CCQEIzKJw
lidW6Uqt77U2ygOV0pKm/fEtfGlpkJSTYecL/w1jzkM79ueoqIKErDbZmc0g
5Axq9bP+j9tNYyVroCX8HfrWAq+znzslBpWHyFAjzS5CBB7kcWQLlIaN8MbW
rDnaK1KiCZIgAZlJf1lI0Mx/tJNoBbygn/gJZcXRqIw/5LFftXbgefguiDIJ
sWnUV8w5H5hKMNhYdhDcFCizqbGzzV0dDOcfbZbvCxwaBBXNiD+UOSUPFOvI
uXf6ffqIRO5HcXdev67KEkYsZgMlAmpyE+aVh3kTPlPHVDqrLaIpGo2MJbFJ
nlxKGX6kFplZJ1vfgSOI97dvG/IbrINnrN758RNgbqkdYakXkTOxB5LHr5wW
3oaZrBBX1NSKwxFOy3yWeq/KveXlkwsKJf5ibklVKAwftesc4OJMyCLQpLXr
CTBhCDjuoGJf1atskkX1FLPCEdpk8Ej9PXCQqXnh4uF2j+k/54D6nCU/P4A2
bQ9I4ELzXsstqpNMTpSRmUQl4LusbHlKbrEb+l2SBzxm6ZvpDquJ6i6npIgl
AVKg/tSM1/tOwBU9m+Dir4S0a2qOyWfGJqVo4N3qeF3OLrW//+mn1GPesziA
8oDC1p4Rqe4dp16rs0RVEPTS3JnSt3DZfimbNA45BhsZL0SG1UxDwwfyveL/
JO0SEglxwJRp9KpjOZTppREXY7kyd3cNv8sdoxu67OUdYQMoEOQPZl/g9qeM
2iTzqD2y7t74CXjEXGRnQcsgA4Ao33FaAHy23Bkr7tezJ4gkYgPP5L8wRPC2
nt2lfTcxMclcmM5cNcQlMNwWuCQ7+PFyUdHf6wRFWU1BtQWHUZX6YB6RAh+R
vs7HxflvowpZpYtQC9QigClwY1NHMK7fEW8A8vmXtahxb2ZXOShFCexVbjis
IwNhLUqWTOtguGJsdVA6snb+x+IFnrvjunmyt/IJFgK34p4dYgxDxhmgDgDZ
VzXKS99sCOWwA2kwV1h0mE5kF5eWpZviyjkH12taah0isP5up/cI0xksjxeN
P6QYV3YnMrJkeLvomfyQLMqMSJrPSh9onwrigKh6R4SPK91wx2f1/iwusQ6w
/W+dxkA8cxUsQPO22lBn4MJpMls6Z5TZek2g/v6s33fgFbFLZTPNQxGeLIrG
40M9t3PyUKUS4Hh1aQMDt+5xb10YJhA+qVnN/6nuaee7qg/TF1R5IXFHt3PW
O0DeNzyp6GvzzStkwXutyHsCyR5PA39ivmCBiFZLcpz+m7i7mZ7/XFrDfi0O
m2uxLcBJqYGv98O4P/7FWRKVPwGg+So2JL7tPZoGkaPEUFz4C22/qbosOZ5e
awwDgvVpOpmuuwp0ExPnRmyLxQ8bdPieLWcyG4Vk5zO7pw+AssKzhSuhQzJJ
UQPr1StLsLdDUJauMpFBtXAYRuZnRd68CrI4j6S1FtSUo34rhRMN2LvcBP4G
DkX2ILBtTskfw98q7Kz/bVQfk6F3tsm96R2xgbroQo0ZjIkqLh80oH3DWp5A
n2jW3FDNJn7wbToXZwB58tmfEhRiQhsXi7hf6qqOY1OQWMLqKgzkAT+mmkXy
oFu+GyJGBgFIL2fBtqAopwR6UerKWs+sSUdLnRUP3teE25OEd90ASczdSUx2
xu3XHG9OC/ngySCoFq/pkvXPilUudzWbwkuJ1VL0RucX0Z3qbaqMyS3cKu8w
HnBM8Dd+HYMU8pJbMT8Z1TBAjlqwuy5ApMDrVLtXv8jpTDAMYZldZy8Gf2gf
SStGegTbTU941Z3fJA6qOlMjtUmzeR2PxjOPxhdNrnHmVcqO8nfxR+zF8+p4
Z3fOnbCJIiWWxUhDeXEVwAYom9hkrIyBbK6aS+Tt0kOFBa2TWuNP+pncwiBP
TrNF8dn7VJR0wpxsSc8bmtqPxJY4bW+Aw7qKEqqprveHNVR0rmJ8J1CT5RDl
U5d0Fm5ao8ednscr2ZdjNbLcYcYXfWsYQzxU/uLFOYJPTg81jsQvRRDCZ13m
UWFmm5+NAPM2Y1CkXCFqPUHmgnhjiYJNPUWsHLAjXDDOPaaZeu6WxQb1Efqp
xKoG8IKFVQrriMof1tiSh6i5JRKPzajHDt9wcA7suQ4OjRERnbsD1lguFkZH
28Mu44rXuJs/isILgkludM8+JdLLnip1FCTpDbfkr9Oy+2FL1zKavfisvFSm
7MWzgGqe7rj6DCu6t3jNl2/4nrlZHFVqsXykacXSa3Bb0IFI+0JxCPC54uvj
hN/rxRKlPnezvzKQlLxyN1spp8hMhVCC2pbb7k2Uv9CO8Y9uLHBdjNAfOPjt
HcsfQLcvXkNjkmu30Gz6wWcSHFR+9eyFnlWRdFUzxepwCRgUDF8li8CNgZ0M
3QHCmhxxW61bmI83Usq03aPNRMIP/Zi32oLwKoHUp7I3aPYwuJ9POl3okO83
PlRHICUSxcoUDrx/LCJ7E6e79TfPcrBm3R4+gBanKcdwZqbnr37/baLaQoeD
O2U5wBjdAAqB4nF5LhaQ2PvwrHydyc6gk5aGP1TlUbGw2qLnr0UshFXai9Uf
kuLLFUSwn8ladNalSPDZbkSRRss0bVoU5OBiqLi0Z0OEfJIdXim6JCvxFsmh
jsD24V/izpx87vHjvUYkfa2bNKIYZ47Qpd0ExfhpzxRW23gbgnbAjvnhnaSV
EKLKfF9/8ASPX8l+ZGczAHr963SQMoUIf9TU2NuECLaprXCfhIJ+vNzBJtY2
oygx7TZb1jX8/3T/qXNxKDtf+afH2gLA48m5gLXL9I0bAe5iiHe7y0ST5wKb
XvATZpy7rMvYoPC5r6r4ymfi59cALhY1RQWVbAy/+nZgM+xTK8hn5D1CNrcN
m532MQuKp48BGx+jNbIgDUWyZf6UhsNi+FQzciXJoZnBvHwvWyCiMqvWszRS
NHnVWSk+Dqpl5HIs86MqhAs6T5JMo0/RLab34kKfDmpTG0sQiq+NE84QX8C8
n8VvBqlB7kycFDLj/3aUTcnGcvLbblnsBGa/wPxznLt3IUl2o2ExZHTe3cVB
yhzGIyy77p1yOnaTEOs1h5EWKFJ6JtAncDps6tdPcDAWFRBVJL63X+42HePb
7VvJBwwKxHopUw+0e3CujloQmXxoF72/w6Gvu+0HeZJXscSI/8u4P5SDFSDG
TfuEHz7M6cszDL6jn5MAGhpgIqdtEVRDWlPSdML1ZQXCcS0y/hSf58mggEQ7
AGsJYWHbaKmVLiNyESjnymG8YMGgvNB3NEYjbesQjynnGtLUsUHgkhaM5Nuw
9fhzpfNgCmFCpmRf8fJr9cvRnySP8LU8kBG2tdkV7Zb7fXfAnRg2RQY8I+Fx
jNutcMy+nmXbubE+tj0cR3/u+Hbaw45ZhmS35WONeTaAGpuVEg9GaCL3hgLX
I5AeSDGDZgw4pKrUJ1B+bt1dQsEK84UJkTpol+HI+HVNCL8MqNfgvO1Qd6zR
j1776P+HbKmbQs/hFNfePyR87W5Mu16p/8+t4f165vFEwj7fNh1M+OQcjzVX
+A6PqUVWNCyZYGF4qphvfpLUUNB2BKCKITr45mb4Q6htc2Ih34RtfoQ/d7S4
kAn07BhlpB7Oxk7s8CAdkNKjTVKSelloyFyDV1iRL4eRJ9ECmt+5SxkJ4X3T
QYXJa2pYQ9DfG5eYxtKLmsSFtq5tfSoJQ1uusJst/dCzxYP3yq+1b1xGXfUW
W0fJNo1VnIyfsap7GxNT8vkiCM0a/5YAcqGuNoyhBQ3y4G3SqGD0Esp68YeY
LacLSsobpteCKGVggsqdw341bJlabdP0CR7RXZGBT06jok8e5kFVk0N9PA55
yy4RYc94tV5tZulEwqkaZFIgBfT2tpt5DMFo4GYwavBYGIk8et8Zmj9e3ZIt
JpEg/uu2fhL2vllEj0SZdkS0BZzD9kkfdWoKbn4knVZcVnn5SvUU0IHj8h9U
WxaLf/i9OSZv57bX+vTNbDsyHWYfMIiMPuONOS27rvdwG20498X8j58Ac/5U
eFoPw2Hk8/lZQ7iccaOzRnV6m/wLBHZjaWNZNvEubNFERKwLoWw35WUsBUTe
vGrFdgONJuThOqsJWm4qUIALbe+MpWomjGcaiMuKHO7UVNeNc7rnR3TDtk+s
KGCyb6ZtwRBqoIomeZ2E2nD452UMqn69ZDvTE/4sBQngGAiHWLW21ASEPg8q
GVgDoFnpFyW1vxvj1RfIdqcMti2gMJp3Xg+H7esnmWpFEdwTuQsDaG4RIUhB
f72PWLfB2wR8nKe91PypJC9edO/Fz/BibmqI2bKDgW9RR5ztNKTxZ3bk39ei
3ZqxYADoAMSYGAeJluFTaCuO+1ptKa4K11QZc1L7rQ0ZqyydPzXSb8tK2Rz/
+VsPKYmD9mLxJswUnwSr1wySAWnDYlVYeu/uBwuMQodtlOqCtxsFcbfPxmAW
DO/m/9J6o3r39a5nvMupF5a17+qSyvXvn9/4ap0frfDD8a5qnZSJ5DFP056n
e2cUfjOGp89t4JC2Fm8GxnsUrfI9Ef94zaVWosywYALfcYJ9lxpZbEPlFahj
yaOP++j9wLlaJyihgxWxDPUhTkpAzwE/3a1tNgxe89BF0WrlEMrpV3vhusyK
MNrDHHezJcsjuOcZa3rv4raGaVEQgXtbW1TmAG3JX62pIyCjFo0ug6LL/Y8D
5uLCCOhcBefFDEKVJL6OAYzmC/usVTsmriDNsOd5B7ubZTXUbrmbDuNBMllV
6O5WluLzU6RnEj3gki3ZjS+SAZGsVa+n8fvHjvBU8lAYui7VXtGQP7ULJC1P
FbJ+a1w640uTt2HJxOmbezYwlI+LS5KDO7ZqVIgnLFW7aJ1T3ZRA80GeqFC6
mowPZ1/XrwK9NkBFbEdUGm6Y2MU0tRO6m0pxuSbekRi/xzgHRvyFAUi3jypp
vv6VoOmfF4EozzkCvAhyxt+J8r1xMhA6VlHmNYdlNu42XWFCU7HQT/eO69+d
7oEfrQYxS8fY290OmYOgHDbS0sKMy9RMFap8KCxFflUJfSrT4NT9gKzU94kC
V0smhB8LSzYBvjaGcZDoCVlFZxaPIuVitRl2ouyI+DHeK2Wv58WWgNpw5MCI
XQOykaXMTSMqMZ0YYgWsXrFviYOf9ucglt5sZ87AQsYCBh/MScbm+yi5nI0W
4mUVQKrmYwT1EPWGWbUBSxrNFSVRRQ9zfQcsDf2E8IRj9w/TsbbizhRxIJCa
FNulV8dl7CmgB59UcxXdaaozw71lCGHhxF5bH2DtjlqdTaXlxQMlSpFnSF4v
77TBh4qmtUjb0S5HYSYbnrK6RwxbLMnaK/EWxpg0ZEtqd8uklv/qW4owAkmz
oOrgEgjrbBggUAnr6E8TB9E4lFjFuoNJzV2XLLW9hhHWTV7FVyYNRQ5ag6tD
GjCK8ZxiN4jIZfYWWcm4WjJPdQTZ7RwSOYGW9540cP+UpKXMg0Ymx3fXNKK9
tVrxgDHBLVY82C98FAxlAYnZ7xoTjoeH9kq2yfnV/QCrut4Mzdf9drLUP9+E
HFcTnXAip8JajVFhvdw2+Fw4oz/eLDHKM510rfkqxBNdSg+keWaNqGYIdOtU
QxZox8UJQemZLZ8sDwC9GSujIekh9OJ2sbcK3lGfMdolrHfx+nfOzbQb59qF
p7yMdODns0Kk3dJ1Y2LsVX1kgxsB1vxRdoRKSgFfuabyL0wM5jyNo+hIAvFu
FA0smNJjct8agitTb/GkacWYDAd1nLjSRiC2HMevSjEGVYllqZX46CLL+X46
Z0hXzMbyLw8YeWfh+vRhH1OfTLlLrhBJKMqBK+kmkkcOuj8KsKu1a3b09pZl
JfFfMkYZUsRT9E8qPxk93pWynO7BC2MDpPny1KPL+WUL54FnIUMifOM6M4Fo
VrCqOPfPHXJjquJ6/1187r3xj3DI2+4Q/gcuvU0wsWPUZG7/HxrRb25x5wfs
ldtNJc+nQ98ZaFMrZ34EVo+ydupTNi2vyhZLysjT6d18K3S7ibb7xZeezQ+X
Z5qNYZ8tSKDkSrsjNUyMOou9XEmI0ldYB96ml9oi9WOtKSaLJiTLLM1cuBDC
rHlsh6xNO2Yq6415b6LNUag5rLVuxymBhRTI8oqtKFinh+3/XTJkONBJoZ67
eWJAQocO0f+oWvpFR+mnjUa8MtUwSHwYOgJ8xz1ZIM73MsBYP0nxvHUex649
cuLxLBaWjjUOifObpZ1lH44PVBntMNFqK5ftnTtNezquT5//VGaeuh7UxX1F
3vOEDbdNnezDkB23qMKtEgOq6f9kvsFhdWr3cg33nw1I5YoyVPj1fXN1PIgR
mEz6GSzOlXh/8v8l9Z7wCt78iIVY6AZkQ5Q/WPcoQ+5DaMDC/rPAJP2T8dY4
Gwe1UsSd5SO/itJuMMjM3k7mhT5cYu1Pm6yn4qH/VJEqBSZ8jDDbaXsCE07D
vdQvudbGh7rDLu78Hsp3fCjs81pC8EQIzqP2KCkZV0wHteYgs/cm3fl3NkEh
5SiYT8/jFysnU2f4TC305w8MJ5CRCcH09jz4UV/ertjedEZ68CKYVeUndU1Y
o32XNR7a7eCjqLC37b+IkY6qxszNquuJVNSyYb5eSLcfYqxKLzVIL+Np7hvi
nn4G0WLX7LCnq/mSxl2e2mO+lPhD3Wirn1yfwRNBMWjkMasW5WoZ1/FGaEYX
HZf8zahtyUQZUz1Pi36uYJgU2XuHVKpJVNnNfBblYuZn/tKadby9/NsKBUfO
CGF69EDINPvxURm5OUmiwCwc+3b/wXNMr6OK2Krq955RDwBEKUMbp6IO/rSq
9uWe4XWZoW42UjiFrfiyMf7jrhHIDG1CON2Ai2B5i9hEYoVGMUMObhAW0njB
NkbtNpoF0SQQA+D42HusckKFft0aRB02Md2Hm5IqgvZqsxJOQYnMylH5EOXe
2qjh8lKzoqwFiMdxJ9TTylZaYbd5DwhinEtGQpkIIl73og+liu53JqxYl93S
VbYijczcspPm8eFmbLzfoYtUQ2d1Hifz7jkLvgU3gOw5b+gU5Z596SG2Tbs5
fNzS6U6dhJPIGLmJQXhGl2Nb9kew5JdVd3F7aVm9QOnhildzmdSPSm5M7GcR
u+Gurogy9lJyulavI+mws12oUoBfYqn1UT4AoUDypmErNKCoyHu3e2XdQwf2
Sk56oqC2DP5KDqzV09IyS+5qBBfvv5tJil0rnWJXiTU2umA3M8N3eh3RGNAE
kTHFvqtmqohzz/Kd/r9kBdpYfUW1pd72oPzQ+CEye9ImFY37DTstwO2C4kXw
t856kI3R12OnT2S+/zHzYprzLYFD3UioUpAg7j/OVS5j3woj4nNFgj4NyGf2
D5A9WuOYMikmeCBzkMx8WblTYBeuGakaYeGUo3SEYGbJIjCrTm8Tg3OzqajS
n1PohF915shANC8Sp065ENKIMJeG9du1zTD5vOINOqMZ18qke17OY6youyDq
p9JW5VgEVtLtxqbwYYildFZtw/Nb6juOpHcK7H+nRU3nGdNX3dOgjT6NxXF8
J8PAh6VnXoJLKoJ9vJC9k7SHkvjorxYjGT6DbCIEmNK6AfslMln64bV7GGYU
drq0KWXnWJIcYd0byuOEEQSGc905GJMewdXtCL8WCdg5mkkuHWRnhq5Whknm
8VCmJgz+31Q6+JvNJTor6gCjplfEEvgf2dyifPHM4AZFZaBqsGfBLZXSU+5A
edyCd51hCoSKPuORx4Zq55VmNTgDv+cAU7bFDVN23u90T+qfvGahgMXnMbAC
Zonl4Ey0t5sI46MlEK/VMbjcYz+HBcmOvUFjsKZWfys6pwuUWE684EaizmRe
evJE4+5SUqiWsNJT/MKEuAbh1BlKrlIj8HFk00vAcVMoHQUIEsAl/9YcTAnE
rs/rjCfcw5APHFvVt7DZ0qxfJOZdUc+1+xB4YFR9kIfb5oSQNpKwgUrqYSat
6X2MlZm+dcu5NS8SVsJ4uYwzuGlcxwvQT4eeQChplL24+v90qrgVcj/CEHGi
2khp9ns66yj2JRTTNYzLRBZ/9yxOh6WfBx0aYDcTm4llbuS84vSB6+F3QnHC
09QWyLqLx16BhZDXnbq+9aStZru0o4yKNCkRFd5F5dsdqlLaiRBe+810XTMb
JycWkUFuGTrF8Us5PXwN7pSWK2fWhKd1q8ZRBVxftCf6mZ5E1ZgekzBYI7D2
v0AFn9xnGhCdVClWDS+5YarnyurETy6Yf3Q6cRXSh5KqKUYIVoPW8+a/JgJR
aWE7vrhrgHjMy9Hd7EJ8au7bbNvyfT6+hUUXaj+7wmRQV0Zm7zdeBzIjMczh
Z5BYsgcDcls/3rCoGqBpgUiWZ1Op/2OZzTsYnpxns0UjK2B6BYaZ8FHyHZRO
acQ0ICXLeFJz8lhHSjJZ8nnY/WzQuk2rwkRMvGxtviGXKj9GP/zRxES+MAtv
4SW2wrG0yt2HtLqwYLzS9HmG2+h3hefEoC5S6qUDrAGEpNN3hbP6ZdoB55Il
E5FsKglBIr78uCJN7FoJZsz9cuqmpm9lzgyqPXfsxTyuch+TuomIrir6HGSM
D1vF9Bv7isqu70F8q8fCyxpurpErHXWnknM61BvC8dyasJmcNb5iiC/rPOhI
asczKvAwaJcuEK+S9lQE3BsWfzKqJ8VRCaDDlofyeR5MnJ72WQ20YC5MU8xR
umAtweh+GWz5OIdMW7hlDoxh8nAibBNN9DS0LsIcpHxK7AAdeB3o0S3udPeX
0vUBAAzgXMTe2H2TougWLCHs21pR51QE2uDcwEDjlQ7vWUdewo1dVwbfyJjL
VoqF9lVl26jxeLp//cJ/jgJx7fn9PgIyGNUXmbP9nKnx3zagUL+qtcXQcrJx
nsluzBogDypkEFNVId30BHNCZveStlrNd+NIMsAyoAOb914bY5hfY1dFRQ9X
LKg/9wopR7R0RME33Zlw/RCyv4SxBh30/b3NrgYp48ZlVevmakZeDbsD+ANj
tZxdqZACoMGWNkUMkhsr99G+3IqPUzsASApzruz+QJA7XJa/3LJT9q3XisFh
PE3pMaCZdANgzkrLIt+uzgbJyPmB9NmBFIZVv4wdUWf4vPbTW0ykQDDYLElv
5C8igjAI/VDOYMxe61zy0lbr08wgeQX+/c50YKK15bUfglIGCN1BAGxLC9y7
Q2ZcZy1nB3bP55n/yqEJnGnDNyYxGvsHhWZldlL6spr5jc4El/FJ4i0mrJUW
dCSdY0JyVunW19fTA3O2u5F+uFTUZsJjUiXz7xW1mYopdLc7y/LEXmjJKdvN
h+FitOlWnrmGnc44pYwMHbery2xk7EIL3VQFkuA6VKcqyoXRt6Pz3vU2Urcz
nr7LJ8ZuKvWOraCGUHZdiCcPF+SudnoPvNZ7Z8Ma5uKy++EmoJXhYvuc6Soq
azQ32kBaXmyJhlhpAnjrfokGwLhHtnWDpJq9swoWz7vuVeTPFNFrKi3TZ6tY
OoPsL0O97JhPw4uzojJDRiDqdcnYykPuVN9uUNXeqXYpA9ZrOrUeFXNEf066
XzGnSEsDC7T/hBeqHSDFeX7lKFlndg2oqj4RDXCO5Vu78lT/cqnvjwoXpEqs
YlXIOhutnLjAs//yu2v8lrH1dxrZmo/UjzWZXPOMkOUcwd/iDGyP0TwSqY+/
obKkCTOI8tPnaS6QJqruSKdR1qnSUAX6re8m27kny/MffOBiU+uq8fRbW7+P
ic1iX+JTo9MnV8he/+nh5TEZxT+yma9P2GqOlkpEQ+FuVZygUFwW77Y10yET
JZgukIu1aAsP2iHwmX+ZCd/jI17ItnUQW95jpig8ANpnROBfHHJHy/XQIrue
fMD38CoNms9WwiVze3S5z+thGQPdkVMSHJ4kLEcVssHWNUpsj9HOisZ0DKQI
m+oRb+LNdytAidET61B7gIkqfeg7Rz97KVygHlWOSrip/KwBNUsBeKWUgsSs
Q18q/OMbbMl1wxAuN+IXO/e268IZRf0VT6KWdBRMRKk8bOv2ZQKMVPB4No9h
gS4f1oJ6j9b1BpzclJKVSFUaxjyE0SaSXtX3MV9SGpP8n0hsAeAGwZ4t226D
a3Re6NW7R09CZRrXWiPjLMx9Bo7eP9Jyw4za6G18Bytpnx8Ai/hUu98xkyYt
JqLUsB7U+Ko5P8lz4Jk7fiy02TcH7RDQ+Q1X2XE5vrrM0Vz1w7PrP7g3O56j
OPQvl6RVixbIVJgohcT2FqjDkV6/G5cUvPpOGyi+UsBLyRoH5k/Upblx2tiv
3p55JreHcwGObO9j+1mtkoQrmL3c+1B2Pq55eLbLaBUoAEnEDUsgAZ1B8aVR
h/8hDvGD6epwEuA7g5EvKTlP/5LuUbMZdXnMcL0+H4M8Rn0XTHyn/G+JAhL1
SVoamJPo6Y/8yQZ6rFPAwintsJoS00hQwTPuL8b52MPPqkhP/xW7uLlCsDS7
iG80HvIvzTsJnFusInsLy76Bj+TepN74Mc+N4Psh/X2pXEF6Mfyju3poAZM4
Z8gaNmlObAUmnqJhpRYiRwQN1FZWj+r6idG75vEE0yV327PpkLZpgpqLs2rb
eeYOgiabfdsCayqHdH5VDpGCd5F2Bzadn10jZDy2CsSfVl5Mc0IIsk+bNUPJ
h0jKK1DYBKkFOYK09ilsCdMxb7drP+RXnZcmxc2FhGDYQQXr0ZK6sOCVaat+
HBAn88EajZju9ooLPtu0TQACIM1gv7O587HY3Gnf+95d0e3zGO33Z4525wgn
gzaYelcRAQxCbGvmHJsm9vMcHXuvo5G4Y7pO9iVKAVhfAafqDGiDh5p4JfLC
1McJATNFzWSRMrKBrpN5tvoRtGG20DKX3b0vjfwDSTKGP/JPxFneHNQl6bMF
uL2g0WvTdxWioESBFVLOPEUnbV4YYzikbFafG9Vux4QOYeSyUhk/1dp+NP8/
XwcmMHDpEA4FgGg0hfIH/N5zp/5rg8yA5Pllee4W1PJqwcVzN7hvq0ZENTd6
5uT+6DIecagdZpiZHpyuJ9isYkTRwAIh7snMTbMp+tDQTL7gYbyEMJznwHH1
Vt45KwAgSG/1jHHt7OkdeaW2s+iMZjpNDgx9RtxC6xMqiPVu6xtdHcWC0RoH
HomAYQzhnRuCedOtwGzvfTLkdSZIEYWKWhhMNHon7M9bsfyNTDOL9YnEN//Y
0RAlGadh0OIX+GwPAGHGJz9VKpUOTuG4HFA7MCtr2dY9rAF/SWPn0NArdlA8
qQMaPde5/wwmBJ5J96NhRI/CF72um6cMK8R1e0MOZn89Hp7cN5CwyyoR8a5G
nshVBAO3t5lIqGMeKFffgV2S/VXF1IY0/r2Sejb3kE29xpHXLJhJeRIIzbPo
AcwER705GRx+uf1DSrHpnwj3YRCwxa47yMOVi8Ldzlak4jsI271fbdc6wBqe
wYJLynvISx8MG1LNuq9nCUGjstK98/IPDVPPqMNr8j/BubEpI5pDa4qGctiD
aek9WIkmFdGx/BesZwEs77QX2/27O7NU/nSzuJObiojc5YS+ew+3ZoGy8mG3
oonsbiOCOBw64Zwr+dksF7d0XmTbQj4FqDnUUH089Mqi06wWPy0oojWFxlTP
kyy1/p/wdAeO4cffdacErCLB6MswlUxEfw0g+vZG3vUEeM6wPXw3VumSHI0C
i6Tpdmc0XGf+1tPttERufAbnAgggt8eZjaUWesph0/pRXQQvTN88i7UoD+dG
G/64XMV5MuQhQrqXTOKTZBbxQ00Pkau4TysdZsOpl0+swnFKXpm6pRxO73CI
t4APD2oRftrA/45JFcgBExLJ+ksZuv/ABhH1Deybw1w9r3JocqEtrxy3NXTj
d/68oSauxTlteJZS3VYcDOuUPhFX4bRHFNoD2XSpdtpKUZiKxC19YM+9vtgP
60FxKw34lubPtHocd0HNBW3e2RkpVqgGVHCK99+ild+HPLL28ywt+nqRWZ2+
yIPpc2WkvAShp4bEs0mc0duYRQUG1LgPUKabhsrdK3TaWFkFH7I7yMgNh/Xw
URuO7wDPirheyJ8JxCjomEPGOLiahI/9mRjtjUsLIwD5Zq99ZscwTQQeU4+S
EVvlWGo6ojVndg1JOGFcdZq1zobfQ5KPkthfgDPfpV7mBNdYUNDHsWaYTXqB
M1SEj/0FOYwd0tDT/uVdCjJORAN2Pnzk0pVRvV+GYXcvkTwxXnsxEFsIELVC
e0DYcAwPegJm96NYco6LUDXnMmi5B2DQ96BcWSYiM+i+20tnK0UidgbROpIZ
k7awrxRYRAq0kg5f8rfGi6e8ZAHJwjngHWIXpYFzAOcFv0Dis1YdTeh/JGWM
yeNSmTsYKaoZ8+qNp4d0YQCa+w3vXyvwmpoNa40tNcziD3v5J9NUWS0dpCSk
4S5TMzRNlNyHix5kOny0iZw3+B6zVZEFsAEAMGjHJxaoWVmBTCl+P4Vuvrv3
jCayY4azA5mMEIDE/YrAWdGXy7ymo/R3/KI7i6ce1J300JIhpN0Lu1ijG/us
ieA5A8VgFHYmJCAFRA7xOs+hmVdnCldEnhpnu++Sz/kusWxIaFdFcNfvhy5S
lLJ3/S1AUJ4GrvSrdodJ6mgQBj/3GXh9LTE3vCkog96eot0JgiSzOkedOS+m
oMcjPOJW3zzdDltDYAdTPcTBxTde240lLHM/6jf6r8p2KCHar7ui82Brb0lD
QASyVH6iZNcItdV+la/e2phU6zl6aTisHmtsU1nRuyu7oPBVgLTfHoEWvjwe
AV7N+/WXrDkABva3ut5TBY8JAY1Nz/czp7SInd+iU/P2HfdY9Q0UyAQdDk8m
0KDKxCBASDvLaRpTjVK+x2JrH+BMNJAVPvq+szZSu+WvsaKzEBTH2Tncl96q
4B1BvtXKPEIUe1WHJsXIYkF8ucIvAYXMaVGWL6YYYCf11jZmX6HFXcYWLYhf
xQxc5BXKwFGCpz3CgX1wCEIxV18XBTIN5NLggZTzIZIrOaOmrYEAyrH8k36p
CdXKCBEEK32BgDi8AAH/0q2YoXKhr/M3AWoZCDZ3JXVkdRKgOG2Aup4US1TH
VBgRxwxPKm94QSskhBdHmtMkeIqb2K+yZq1kA1lDvlRjEY/21BSkDOMm5sKS
CU7EoydX6wJWKfxyb0qwuMLhsKC6j1gtsvcOZGi2JbBsNbs2QXH9ykQLFAmb
5QJNJSZmvY3t3L/jBpAZuwtyss5aKSSdOVrI5olE6+0YMi1RF5bPGqoQko0b
FTbWE1iN5k6W0/rR9N/IVvyvTMzsiWOLYyBljZw8gd0Hg+mIqg2X07SwPz02
qCmzMe84a4wuvZ9C7Z+TMWSb6U6Qapa2f+aSdKNqM/Pijy1KTogxq/INxT+1
U+AAd0HK3rs9g4/+zaxKeBqXDNKG/HO0lwbqZJzI91sLbmAtU6UdiKN+L/rr
njUVysbEPRyk9L5k1zeZaziCF0pVX8j2eD5UsOSPw81CyTmN4BSRJfvYzEDM
bkdvNeP1PovRGssAiKjGMuJExJUg+o1617OMjLjMQh375OU2AjmCL/0yjA7g
PtfX2NSktNpL8Ha8AoV2x4Ajfy0MdLqcgw/ezXnIKFCtPChLuNdh8vlpMInc
98heYbbINo+md/UhRc+0dVhhSgljcN1/UYQjsXw7qKLjywWM2lKX1IeZzR15
TpKDtcpgPtffHwVUrbaYU/DbJyV8zWSW4c4ewoR1oLaHRz03oO+Hy1yGViHY
EFSvRiz2vrBNy4If3PvY5sj6VywbdpodKspXkZDFBii1yQRixtja+K6iscJA
RZcHYvSxRZ6v80vPoF5eofHIVE6SCLncTcDqzcpMUXW06qhwBC1SGSLq+IaL
cNmTofBkqa+dCt2sMQxv3cuItD0n19Ucjkmq9gUBU+18W9R1J3Q4AphZ1xXa
DLyovGbxz0JGW00heFkuQfkIdB9axxwLZggaVrkJIq5GvmxFO1ZPCdKfj7Kx
v+RDXLP0vSeYiHIhQGYcDAoj0mXF5XMILzObPNAT3HE5kJ2E1UE5s5uvADjl
/ZqGqCrPynHdUMByk7fXMjJVaDwmpi4gIY6OTxn6nXOJgBDJerMKWA8duDxO
9KSdnx20SICf2EHsy4tASYkU0nHVs6sMKSLHA9SDHsVElHhfsCg5poKZrjH9
h26qpNVoHLRLZvWQSFSD9BZNctSFcsfNBsGSu1Yxf//VeLKkAyIEpSifovYv
RUEt+eCIfY/PGOvJh9E+aavTxDRMMrmbwBRt8aWyGuKQXJZS7hyj9G79l+Ea
uFxB3HcBt2kTRCDvTdWdWfSZ4I53YkaZMLk9aBryp6R5SHGH+RsH2umRAT2v
BTUgl3UnJhqfnys/RVFqBmUFikBBVb5n6a105/vfTAiA+kvqTmvqdVPtUnqE
7KR+uKiuDuhk3m+GzkMOucdlXw0q+EeZ8MYpw+Zg5ffHTt3Y5rf8KN6vprfP
9CLQziPSlF4KZVi3hxFIGsE3YWT4my5NkZXCNPkChufwR6Onr8/EZiIWqqpw
DlzZSFMyaNCqhP45ukynB5pN/aJ8kbPw3Hgrc7UIEv3CEQiNTJdN91UArB+R
zmBb9pZYjp1EdPfxaUFwYuBZEIA9mwf0ziB/XLK2jKFCAH4aHHg4VWMYCYpQ
TOscMCfU4MQ5DEC0Km+gt0cP+lC7uKOkN0BNRkBjNMmQBi0xZr25BtaOmdFN
L6APo4DsYHn0D3wQ+8RSIWTiAsXur21T3HWra4g9dCEsWPrEqNQ0uYTd5RQZ
v1Qu1y+n+fP2FAZa9Tz0wC8U5ILDINaTxMUcWAwTu8CcWCD8FJSTNmWYlhMm
pH/T3KMD9f3NpgZc5jJbfywy555ywscNIeZjbks4aEFwFYWwV/+KFb3IUSzu
lDkNNZWouQVgeuaLb49wV48M+bxFbVnOv4xzflyuhgh/4jV3gxZPrr4v38wv
ujywGuzrbwCo1L9FGDKn8XBSHlc7OewSotFBL9mcu/d0kL+W7kTBF7qhn1uf
WmZqBdm7zZWApMsYdAHXDZ39s2UEqzCz7uruR+N6nq7EqxvO66eWIhidpaQD
z+Jro4J3iIpIk50nv1IrSRFsZiwCco9GvMw7iJEWCH1vrYDY+GTSE2gDReD9
38uepokyUkmnKOo0vKV4MFx2D0IbdcXweTXWbA8jIxuenkq3++gRf69YGJVq
qOauhI/jcqKIMm6soAApfM1475wmVIflGiL6cV7KEbN/jj/mFUOLR55Ga9kp
2DubpGeiPSn51l0HWCYx9MKWWPM5WKdDnpp9/Pm5fGPmWCV+R7Ij9bwJQB0x
gRVRMetsEI8QQn6oTLuSzcwaAwIvtOp3VWdkHhfjIJm1WWhqc/vLcNa5qNR3
dNO+yWXfYcH1wudtSuOZAczlVnFy9USyRvRY7jCRbzdUKcge16As6ddTtpNY
uqcz0s3AXJ3vB8h9J4GTzL5f1FSx2VYPVdx9dDqeurR+5R1Q7FTri1snNCRT
tg15Oq3YQsT7Ja3KrojlC3/N1uoyBj6MxvND3nSmYUjBjjhEpDmzc89s603m
29VZMnUGumx7eY/gLrr2OSy6I+CGVGBocklqkVPlv2ZL/Tfa30A9xR4s3oRz
DKpDsUzmi/DGLlH9dkXenxhMuWmFXKLAEKZZpYubiqHoSm4ocNvgHIXpCr2l
LzTiVcnfS5iC9xZNzwoSqIFS91fdpw+KZACvMuDPIKNRhTgD3MlI+Jh/oS8f
CNjiTx4BcTxbNVoKxn6w4MeJZaKMNyRFTgt9zwUx4zEt6ese4b22UsfrXpAx
ls656eBmkS20E8ZUhd9nJGiXq7zghfsLQe0Utq5NIZMJIQlPLrHe2YpMtx7s
jtvoZ6ZpOeedFbh0mXesLXuZr63JZ4pLcC+RM9fME97bHBljXOx6jMhPbn1I
eZrphvt8GT0JkQM5BMqNr15cKx3/FDuLwBWb+axBkkKlL757zJdJaeTa7gFe
YeBzgj7puueDo6UkwXgZ3NghpJxKIhp8nN7Re9r8Vi5ecVkT1es96tt+lWEM
XhPE343OF9aEkJjXZRZ/kYRCvp0dRDGIBcPi2hJlwQl0J0TOTFWkkr4iD176
kGnCog1RTmNUn6wYkiK8j2Jnev+dJbYMvsUUelIeuCH1ewN20KctemIOdhoL
mzyjzlfIH6LjFmFI6/JZDD3fS+IohuQxwybydBPf3Kx2ADMche/IsKahvGyp
tmxphUIlvr4HWYmJc/Gh15CYziCP8D4+y8/xIFBmf4f/Li1+YJKUefer4awF
ZptTKwH6+SZRl16sxI9TWgNcoutz9stq+dkCucrzpdxOdSkg7/Hs/SCHtGPP
Vib+FjY1+Wtbx2WFva/Ro3d9DQYdgiy3+UicRdkbmVj0z2fAKf1gj89svj4E
dHqfWtbK51yxAudt6CGmpk9VbQOnh4DstyDeKC/vJBgJ9mnlM1b3bVfXIcDl
XSt3CPI21zmxzBuPFbaVHVt2GZmVaitUoVy4FKbkzucs0fYBFnDLsSrCz07Q
01vk91+3BS+kdkB82ErXEClhBAUfy1FcehRjOP+7krHRIdMFmta6wWk6df+S
24AmFZ5xtuMp1OGI/rzsxaT3sMoTbrQairqE9DOamOJbMr1Mm26hrndCXyD+
F6BsN0jlucEK5n/A9ITKqTU5X7gW7k4r9AHCFVZ81t+PtiJD178d1qOjkD4j
tBGER5JsBwAEm2oZ2VxJVTYvaouY9hR9gONx193/3XFpBnZubddSFFIVkl/b
YPdq3kzpTgZwbdpgBi0tfyRjI/8BU3sef947ngvnDLgYf0HcrJZ+UdlZUZ5b
y4WDSWPeZDYVt3A+fvPMAokG/DtJYsrLkEMmw+JAmN4eMObJTVtS7GZ5LN/s
6U2TSNOb87rAYA+rQFiIqWh/VwSzfimq0X83grZZAiKFD1kjiT7QblA9c7Om
ciV790prMMbJY47G9rjiYyZ2sln6MGngIjrMBq7wnegfS7ia4j/CbpnoNx85
+z/Uye9cYnL/+YuSG10b88Mcry16AhGIOhFMf/5O6A+iYCZNbdELbKAkfg4F
NjUcXG3fc+oSLYepFOXeT7Fme7tSZQQ3fLNV92HHz9Y7UUELVy4a4/MdSkf4
8ULjQ4IYJyEbdfxWt0pwWowHxoZjJZrXbjA9TXqKvVYdNb85G8HENZI88KCb
XC5z+DlIVTWtaJ0SDKnpUpNNNQIj3M95UdHG8MKtQIASH3kbWxcJU+SNcCCY
Gg6TkzDJAS1pmrUbZaDoaeltX0NvXTp8H+Ox4Mqsw7bVZ7NQSTmL22KtiLnQ
lNMPF0XgVdwR582U7bFV2hlT7QytV91+ob50yrxJwnxjhDjpug5izUQFhLUS
UXcwvAHIddDweYghjeDE0fyO8NdL6YbPUBoWD5CPg0wdIMlAshx+IkwEuFcp
EcSSGx6Wj3uwYKCvn2sgeSlzhMcvgQFLyF8Fh30lA59iWVhbmVmxycP+BzIW
Y+ZIqXQ6qUeO3ax1Y+OlEWszQob5Y+6PfiDsAykT6EkndDkMYth8bWinvmGT
Owthn53LqF3BqfmJf2//oBuE9wU3yKCc2PtsKAJgknW0ReFtYKaGaZdt/gBc
IArB879w4n7y9aXtx7MfwBLINHMosEelWAXb22U9iZsm27xhD+QK2Z2HtIzd
hTkkRjQqtK7uQTeRylt/ixRForhSrHzXHr0OBHRMIo7sOGKcJaoRLFeguwX1
CJZ5SelGKJJdVuFuInmbocEqQmuGwTr25M4zWuBjHL9jLbKDzPdHw48FxNK0
zsVXcPql1bIAYpkebvVpuYfkZarZKBLIEpEoFE0nksCfYXJg1nY33Zyy1XxR
URzZZZDzpNj/rr68mDi3jMJSkszb9SIKx4b3gVxrpQ+F6kprM0HaYYV8mKym
IAZ+1vGY6x4by1PM0N5ErTu9OkJak+Rj3VWOnYfbqC92m3vpJj4jJjWJ74VU
Yvr4uac7wc38E9wkXNKVoPgBZdheoY3BTuhS+yDmuJ6V6bT+/J1LUktB9g7V
dusVJpqG6I+miLzq0QD4n5CWpmw2GejkoESygDCYYjMEe0TeL7WPyki3+4vw
BlSAr6+eFwOtPx2ZRWc3LaSpZqPxt4QAiYPkN1bgdnqWtiCwvV77B3lIG+fO
Glny/kf+GwC+VtFslJ2lIYfOt1pyWKCFSdpGrOapfe/+i+UW2jOzjm6zpCER
NeZES90WeDxa7tbzs3MDc/iKGQ6kUhiYJ3QgJBPQjSoNIkjPlRrhFYCYFuzV
n2MaINZP5TKIp0l/fnprkRY8H0SMkVV/94eOUfQcM5FundssnVNkhGq4cppE
6ZwzT70Fbe07AjjK40nrQV1kr6MA/22wxHWMZcyae+k3mWQXgb6dLACaWcAG
w/huXChuWXJXgjm7f1HqIFhRhL6eYKSN4h/rOwHGLK2bEotWhk+rHjOlJCFj
FCuVsskanj9EmZBygoRdXRezTzpDEMYnTzNNutO66EcdX8jnZqMIUn4vPh4X
KL5wvbsVfb7v4rwZ5fSG8FqV7LQvZ+kpnZV3ZILVHgVLGgeXTN2nuYfK5LHG
AxAvhO2nxyzntSgQqllKZZvS2JiVtRwzSrKEYx3eS9Tn3giy5c2TfkPA1bDZ
7/mRux6lhx28IByLnshdXEUWcjkfWnOWSpcu0wP+gk/U4B8fGSrS0cbTA3PH
aNA4rNkGJbEFSJpWu1xUskiV6VVCJEAJCzwyiuSY32eP/+PdRRaAnE2K24Ms
QUa8IQ9f6e6Tkg8ayYJvEDm5UJW3YuPeTjTRYpKMjl2TDFwDsWHUdvcf1T7z
Gcn/V9xyOwsyhMEELnMvs8PvxNjbZfYLlA3AS72C+XkBGc4+h1xP3PKKTd+T
cpoOGjk85OkUlDHjEllki0y8Skot7Q5SOcX8iWJaAKhoEREYV3FIu7WUXqXK
x5LjlUHBGgiZuatPJb8z3g6NR76EdTqHfgquCucx8TtbZgoEVNVw7zNgEeiG
/kQ0R2sKoU4wzi7GvQ4Nz79Ixo9pjVRKVlKkdI8x1uRJf21qjCB9Lu4CU/8p
lcWLmr/rUS6TjloOpcHlQFPJNQBRS3godbF9lC8neeb+OqwzpqjpPiUdHxg3
1B5SHhPwB8pVYQF7axTdtxTxdc5g5juckB+7xIAJ9Xb/DldXG/aZYgjKPbBa
1pcho3yHAw0zqF0rA8HLUkG6Tzi/1MUxrHyF7Gq144C3OJwsy+Nbwqja8OlF
BMysX8QYk4KzMwtlPReo/FVQgJlJ6TojU4kYDTDlIlbt0R4/Ws3TIJ7zRxtW
Ieiw1MGGkur2e49SC2nXUxaefQqRevOCn0lcUUtR4D4Otrd240kDGcmDNPO0
OaryLy3vaCQ6BgNMzC51k3Q8bo41dFZsAK5Dq9VB60ynzQM+KIa1Y6HwUL0R
mPnYttcsIfXCN5QzsodULlvbTFB/nK94+Lw/OksruTMq/jESRGOTfDL2oJzd
v/bnKYvo59XKS4MDogp2nnwwjcbij9R29ofa8ojlXi+fI8Jc9Th3HDidVfbt
dqPFC8xaAs/YMQXPrH90KwZ15l6l4gEycs1IxCMcgDBczGBoxMz4q84mNOXy
cLvICaKVnRVGSc9n7FTOQLkgtIJpaBWqpS1+Z4nT1yiGy1FvqIdn3QJdqGZI
uYK+cckWrcniAINY40ZOjotBLwXwQn/phPXqa9B7dz9Vr4WBtqNDkhIuZap1
k1v5Dxo4B5pFiUWeNshEn0eKjAmt+oP/M42V6sAohdVTHLYoN2kMID41IF+e
D7EdY/wUU009FXbuIwxzvsjsUfhXIz6lHFygCEWG+rdWKBr2cB0ZsYQnlCdt
7WiXLuxKYseu4glfixhhZ/9kM0K8PGS8792VbrpkSsk6tXN+iLg6E0cxmDYz
yv1RkUoD6wuW1HjwX6+B3stHfUaWFu0t57n/M46ViJM4DMB4/Fln5VabkcnQ
YKJoOFstbx0ZPlUuwFlUSLahNIS6X7Uwx/ENBK3G/18XxCwUMkEA4SlrepIt
IFYS91LC2c3+PmWfkmw43VAE0EYJwePdXpiKQByBAJFWfxu+3KoSHP1queN9
+DoerX5kb0S5yXjOPl5TtaNPmJzqhSKTRT+/oZMSNJS6qHj6UY5cyv7Klq7J
EUBQU+qJNWwZhqnhP6hJpI0Fxa/7sLolOb7f6SM9AaCg/arsKpnWu25Hl3rY
Tvsfotyu/ymUJGS3e2Ls17mMvAbDvpR6ViooEDlhr6gfkxY5302vIwz7q45q
WxGtxZwkT1L1J2YWPeDx//cjkHwM3maY8eKAI6rEclsfhoLgDuhCt0W/mnTC
u2hTA//8yFd+le9CLLjo6u59OMI01HpuTgwkBSdU9qD73UMK+QfiiazpKdmn
ubzrIuiV4aCYFP173eG/Jk4O+soPOem9MIr2iV0dNEELOiWGBnNiUN9zjr5O
2pVvE1mzqwAJ3K1UHRD9ZGOpIUE00jImSYsQf1+cFrNVW41scOLeR9X6Yt3Z
XSNIHvRz55soFKIsilutVcfKPklZE8iEgEL74efbLMCIBEZceEOQRJhJg7UE
ML4YJgSp9z8OfHJyuOEyL8GzFCZ0UyK5jafMZz6SRJhwmJjiVqkqOKVT5JDP
FtOP6pTsoV8XQ31fsQpOUvaChptBNBQEzCz7HL+bOJp0CwuMu8WUJY59NJYa
lN+xXjtCKykKBxfszVcsyXq8t00WCg4Ezc5LotDBtjIeR8JN+EIzaP8ruZPR
VI6XmwGgZxZMn6rplJT3kFfCVUAx089YxCrPa6q9OyM4VrpPMBfWxqRUx1p0
dg1ad3lIY+3TtLSnVlXVvGfU0z8zQ0bFivh1ipRVd3rpapHQgERnfmneWMws
zJGbwwVMpb6Mn36ZKzl+w3fyLqxH5ECrdDKxWqHYEUgHA+Dbc5TekBS9TRij
/RR/1DlAva9VtPY4mYTTJs0L34oHNJvqb1LXXlcYLCUme3IlQn184QQokTcN
rYA4FBOqClSJIq/FsBsW6QVFfdKFTpdMk8RZj7ORYFM17N612epsN21CRZ6k
gVu6nB9ONPKyc3EbGh+XmvJblhkCtJbqBWEI7ezkDAJ6hzSUgise8JQXMG9r
DdodPNsKsrOVJp+yybWhz0iq9gkPkecza2cxispBGIVg9i5tG5QpZwGZeiaQ
HPkNMqxrRAheEJTTpqge2GQR7ZVUN7pZ3W47PrAVNAMbVAbE4nLP3hKqqe4c
+guHi0K5dVOoOa2vfdVUhJymdKRez2nc7rbd8OljSVv6cwveJXsu35INt8IY
AhZ/cLKUqW6fdMa3k8mXaW68B9EeuxRg1h96Ozun75PlydLL5Cjey2v7cygF
R1tO864icyZr/lH4cRu6wGkE0wC3kTi/OqdM6gL8WzWNkNoaCVWftuU3p0OI
5A7O0S5WO05q/eGvyRYZdZ/er9mIeeebmMaZkJ5Qjqpegt1LJFMGx+Ey6CI9
0we4Hss8boT5dXjfLHZhtaIOEdJ8O1xt6NPgXgcjQWyfXrdbQGE6oKlrWi0I
Id5+O1iOxc+u+RMPtBclSqxCi8STIWHNS2+NCegJuq0hVVHQ3RFOowF6u6a7
eMzxErCvE9ZOTqaGpfr7xvbG/MCUYhpTpQeM7/LEZRHiaNHNI2fCNzHKh3cL
8m8J4r9W0qCHKAYFdeHYo89uGCKN1sGRHkebT4WcaJttAoEohvu2Co6kWqgw
18ujVyYjxk477+Swz8tu+loEtVFWnKHmJmDeJZRVyiTBZZ+XybLACaZJKWk4
wKIgO/GqRljPdTIOkv7hW1aLFytXvn6duzxvN/Hy7kDkeNCkcmcDjkFfUoMo
y/BcaWMxbrHDHmMAmgdXiaQMeDLB8b8deJTEiYfwsUpZlCfWWhGv5l5boUkS
vN4Dq89p7VSzIsqfsk0uUge6DPlnslHhvg3bwf25JztRAO3MaRlDHGz1Q+GL
C7CfGAMZ3QLOm9s04CAWJ3AQck8EEnJ3OC6fMAKux6Y9FBw5cgDZcespsx3U
lPpvci6BTLB+ZeiGmcksnXgxkRQ9IfJS4L/3XemNh7eGuXd9JvPtrtWm9sQb
FT0ncwWGgezWmUePiaLhHNF1o7TRvSQpbcCs6PFQ8tjOkx45sHZ8Z3OB2TO1
/auFuw7x97OhpM3m2Cl+iu9rci2bgCY9wVtkPxb2ZtbQCDRfHOZlHb8j1/Kk
JGEyz8i5Yx0Hv4pY60v8TR5myClISHOHAkSc7+L9bIvG1UNIQlH1gu3FIfnw
q2JtWbZaRuRuv92IHPAYLOHEfl07fYuZ+hUWG0aTBDbm1Sw1WN3l8rnH+6aC
T4lW+Qst++UyU6/yc0aS4aXsX+l/Z9BPmhLi6o3dfH/W+lSGyq+e0fHIm0kY
BwQrkATOCJtWUloD3WNJoMPIgj6bXnzm8C72VhMOi4ZIQg3Ljbsch2IRmK/P
6IkwLdcWxzbcIDg8Rt+/C0z3n2kC6Yzr7psYUSjIsMUgYCM/oGx3hQj8slLx
t0F4O6gvrcLrorYVID1nE3vFGJLUYuGI0kcgznKS8ZmNQTPbWXgKKY8xW5vw
xTgxuQykwEGdwTUI8ktdepd8E0FaYTlDg6S7KBVHeiE7mZsODunpfmiR4Dfs
VPAMq5IgYxwKYL6SSA/Xd1DjtqPwWjI6HSU56ejUKdncjaSvyJw1HqqdAOZY
WyR23PY5E+AkPYIC9HhMqoUa1U8G0o+6tE9QWrxvdbnrXHIfTUKwT1xOwC6z
/GX2kN0ylsm+P7P/7GqyY+eFMiWazuhNV7K24cLKNHGfrwRIIYbD4N53GkBd
LSqOJPdNZOtzWrPJ27VbXHl8rRSVXuROSfiD0d5Rz/TJ4lrELmBkT8+/cpW6
XuqRrhuB1Ku5khIp8zNTYTZ76C0JHoSX7yXbO3HM1hgXlkBzC3sHnSrEPDse
zer6sGlyGQRcRDbOz2ezOXK1V5Q4ZEpzVqzvsS9OqUFuhWgavfnvg5foWqwx
ZZ2MA6zyG2YSrt4p3vILadyAF67peKuqkOiVITngMDwrAvzVoPHt9Gm40YZc
YQbYqGxdUUjxOsbESjZC3eIUQY9OMT3vm6iEhdWEnSrtTu6KE54khQlqcc/J
gTLAG1cqSLC8BxkNv0rhb9Tfo9x18LheeW2SindGe5iwfeMIMYZqXTlLNzws
8XzieXGviMpLzuiuzZOKMFBQBCbZ9yvXkyQ9FXoTwV76XrG6CcX4qC5wV9mL
50i4hRR6sfYhkaj5Q7IVz/Icn9rBQivvhTG2+HcOypsnvxS9K5/KUlQIHYXg
IlvOxHhzN0sIOxhbCiKTDsQKlL2/DRReggUI5PAeORJ19OaEtAYWpSDbW62b
GZvim9lUoeZOhgA68H2o7B7E+TU1g94OmIU+7qnTCrH0OLOpOm86YM3jDGa6
r9wCiveydwwLFOEas17JSsbY4JUqJbcLduv9uLpLwHY2uVU2ppgRx++pDPFe
LFaGaRjwbxpOt4HiDim/6BTMxCOl1dTEjn3F36HauYQebj4pbUFaavKsn0sC
1s05XCMoJ5ySZjXrZF0sm0FrWv3ugijIQw3KAGcOcsMR3hIvKsQP3KmrQyaE
LeYKvQxpHCiNVQLxB+9vbxIELKDs1DOlM+28h31kdPmUWGdRtKcPKwN50stW
jnREHOZZ+hnAXtsGsMJlFY1cNvhz1W71NjktS0EGG38ZuC8yN2yUgtjBNJgL
k+WkwA28DO8pZSBQWnQjEzsbKk7ndUIE4rRqXyDdx10CsXho9aRXLUjq0A/n
pscgmuL44ouMsQsQiU0ak6lQFKFwixidbkfzRhzpVR9kjMwZcC7NS0Rwd6u/
bHGI81EJZ02gThE4JRQB86vDeVJxOQFCH5+A4hBOlYMq3nNWySaR2cdlRdAI
kqOvsxRtjR6VQtrPxFE/weKocuFAGD5N0HdG2fA7g49JvpNjfxbMkrde52yc
y0m54peutIB2rqAvqNVYA//9tCQbDq0gEPOMoOOCH05WRv81xb+P965FQc7N
V3KcaudCrdzcP2MB6PTVEAVYKz24YBH2z7TdVrCkTqcQN1lMZrJAJj9k327A
nYPxM/iRgrLuVyqmsOF7CENdxdpNkkhMMOxEbldE6OFUKfHhZWj9MDP5lkHI
kC7AxQXJMR04JEoHDxuuXg869zG7r5OevDJcFtziJ4XeOrigehegyA1pf7Vw
KHgeoy+JWXoUZv5JAhoLRbKWyQMd2tWuVf5c93eyhhuo+3kX27igGdi5Q2ig
fDbMci0d/oVvVIjKWjCIO2S4xbfYTreOwRFJuTuwu6joN/T0Hf1Ok+baxT7L
bRnLv5e6YBjf1rTzCUJwqSHAqss9O3gVZbJfdWjzWa20BxdYS4mWs0URu1y/
moAg2Z+p2Lw6pbM02MH7YlB0St0hkJbO3zFBHLjt7SKHOtJ82PnxN4dGgfTv
fEms8pGqjPTFEUg+yImUZFQygMt2Y/GJQS7SlpJ80A2ubC4uIjp5bXlaprkL
3tyIMhGkykwzsUJ6cJMnpmKxkqZww3OUEJvh5sA+yGDeBnmksFfHsn1Im7jf
mxsV4qBk51wCUVd9VbJqOW742qYcHJ1C2rlxSsjU4msTA2K+/rYjiApGwtiX
yq6uBq5IpRkvHgfC3RmcGeyLZy+i2ktzGtot+quyQGvHcJ7itfUj5pB7sHe5
jIi824nGB7Euysmww4L1/eFf8O30KDK9adGKXBwXGcjMxSST1F3SyauZium8
fb95g5we0CpzR1KnnP7QNsm0o4Yz+e8zUo06PRox+babUqfugVhxkwGnM43C
7KaTRxZOy5EtTbQMKJmn2WLjGfniBBvxcR/Pbwn1twg/dFMYQzMd73d0RkgY
OOKyXIwG1SuYg/rddqUco8XyVtQa6d6plGcSH/0dsKRxZUKrscZ1Ca8PejLV
0LwPNC0HnrlNck5GLfsxIBZkAiD84x6qZuyipkXwRTIGfMbNepRaV4Qga8a6
EyXVijOhk0ArZ0hCV3pKu8huNf1OrlXZ+X2/fqhlHHok/UDDtFezPrlyVBVk
YwqK9RuFrDU3lAVuYhoz0BBdN3jhV7emPzMEiLIWwBirrxQyA+WFq0MDds7D
r+41NakfCK0nvUxQ9hePX+YnEAI8Omkd67TlL/fJCotpjC7c12v9KLz3x9aE
fhXw/+fMn/QCBjeWFwIy0r7Xot53kMJginhS2pxbwIp/MQANMr9e1a+mRVM0
oZVOk57CoUI6v2IGvGjSlH8JGdQZyBpsd0569yV+w1wc9k0s3x6YNPzydrqh
2jN7kVxKC8FwayxReIYR0wh45xghBovIJg8c5GTSmFmKMFlSVUiX0yPg4xRf
DL+HMqCKnm7HELSC1X1uul9QSv5InZbZTwjq3bg7ViMr5hvmRa/Oa/xRjUIV
mPzqbDQTXS1JxkCJPm85FyNDc7yxZJzl9Xw624ukbpPjdMNnazNtcQppCcC6
CqSqYr15Ah39+serxPoNeqR0oK1Vc3WCguqJfu1vSQnPYQcpWd1OS8cZPa8U
jEU9zOxcGARnPJbD/n4i/FIUkx4XwkNrStHWVt/ic2AaUbkCZRsHkGJB5LYi
mE1nqcJS7IWob08EqZyWnKeo7RlbkZgPmttJ+j57cGUZNq1oOqSHg44nFguE
v1n6y93F7N3+PyWIq7ymnCToOQv5mn3qrRAk591XQlVWMPxpu+MY+/xJRNAh
XmnSYeFtQclaN1nzbInIQeRmnF0biAjPvLrLV3k1mpDM0k04NXcWdtetidsH
wuLZS9sP5hZtk4LwsXKDTtVE0m0D8HTD4meiKSfLi2GUs1GLMJR9ml0lUutG
Onq8WunY/BgIIBz27fhi2jD0Lmyv+yRg3iY96gVr9Y+LTO7X5i8v/iPol+C6
qXfz4Jjljw/9MeBVoOzaJ/8ZVcTxD1iClObOnXbieI60N/sQRNaoa9PC5cvS
v6JEUYixUJ99EwF8vc9AMnJpNHeBOoC72h2GUpYNCPLGIZE0KE91L9RfxruF
FkbesAUXaP91SB7LXPDjCPbHHUIsTmZu6Lf1h/GAJo0+w7LH9FhmrssUR6zd
vax0NypoApK/fBkrLjZi9bAottVwD2McwHUniUp33za05ffv5agDxHalkdX+
OvLSx3N5GqpE0ko6LaUnLuxsoNTcEUyjwtGQZd1j2wsCZarG0tlFxsK6FTwa
5c76o/o4w1sS/cMM9lU2DPaRHFn98NtX8sDx9Z0cAv+fJfXnEZcWUapSfqyP
3mO+QLPy3anuMOIhGlqx0Dd4dzSs9HDEOqdkWi3AEhNQlSN8cldut+3o1DI8
BINUGyKecg2W9OfMi3ujHjLH73Pj/eXnY4L4uC7saunhRzqFzu9RHuLDTq/0
NmiTaCZC9TOAZheG1n8YUsB5IiF30x9t1MywQLvbKuF+q+SnY+nEiJBIDZpQ
nmArR4OR7bybZpCX5aEpTwYKv2NQDEFvpqGbPjOucsuOqVtSBhNz4sZJ4Y7Z
7kUWwedMFOalszGN2vaVaYio3SIqjU676DXjb1tuHg/iRhamUF29FBtEf7Po
9iNiWF+pewjYOGu4cutlADtJWeRXWM2UeqNhmIECl2NMsCQPMEkWu9YaDvLE
vGmsplwP7dESW4XgbZ/F2rXTekO54v5FnMsrW+CEvTb38XWXidqxGl1s7bSi
LGD1ifpQRG5gOJSLFcrE5/uH4oSQWUauoxMh7hrLMhytXMQjAR6FYdlpk+ou
nnJU6C0I5q2gtEQX/m0EC1A5bx95h0aA4CCh6MYkRJUcI2uYvb6cfxDUvTbG
xhxjBkp9w7VSa/C/25g8ze4t6wOpdL/BY/2MnjJHf1wnp5ZkILOWUEcOwmF8
mDzkjJZDmJctj23W2fmUNibFxXH3uPaJVE/1TBY+Q+l4jJk5nksu6OJJShOL
qeWc8w2G9VHOnodnEdnpDNy4j/bRJ+60khxc5oNB84zlcK+g93ooulLpG2CJ
bWtPUFDD9sJ3KUDuc/ac1U2fgxcwjiaXsUM3NGg3jbv6fEd8/RhzjqrG2/FS
smpHzeGww7AjX3QbXa/+fTn+zNj76RoXIWVCuYf0Sm82LltKm0umZRi4FMf5
n06uDyEdcqZzGJ98NXZb+tS7ZlKjpOS2BRmswx78ZpgGFux71p8LrMWADp5p
FDN8F8+SNGrpCDLJvSu3ut5oXQBr7Ekn47zYRWokPUkuyDm9UCNU/kt3soUc
/fuDiRSUd9mJtySYdpNmAIChK96WhzWcaH0MDCnzc8jQCX8eQAYf2tYUt83J
bZriu8JCvZwIDFT2pQVVL3jpjRjSdyr6BfibtVliJXAx3NDBIEwpVh7XBFln
J8qGBfa+hNmcNN4hOjD6+IA9gzjFiesPIxhQR/CJKQcYOXY53/79E5vzWuMg
L6LIz7JDNcAnj4VugnIdv78nw+8uIgRkwQLQDVZGcDUuOXocBbgnouipCZ0o
LufL8YInsNBFNs0Yolgsazaf1g+mXsj2A27n3aoc/w9gRxwLSU9kOzEGswaq
h02b7bpccloSdnMh2s36tJjAp5jg4J+pRFLYCeFUc2fFn8llBrKg8INT0xeO
oIj6hI3Tksy880JQq8UQt/fcFtv3oAa48D+oAzMgQC2V+9d02txl8psqTZ7C
0zg/CJUlb7p5VQOMfB9DX4WyiHqkVDCA2iSLZmnU3TgqFwWXUHywDuZxB7zg
20j6rjsgK3Ut56s4rb36pOsDrXy2M1wcJkvD+JIv9YW5k202ZjAJ/sq1DiR0
/N3Cq/1/g9EBR+e04cG7qvoKywaQOoLkn+1kQXObz3fp+xqdIWVexOiIl1x+
pxnzc7r/CxFYM74sPUZwYRvcTm0nYVP+OVLpLlnLI8H6gJAPvdCfdEAlRC/1
ELhwk4Uw5S7mKoPr/etkm6tbzEzDrQZ4q09Zy2wVOX3fS5FhXJHYDSP1WWGg
ViPU70Z3OUX9niiUGDAqnDoriiwzkBDNmchB9PhIRU8BPip+5yXGfj6N5HqI
pW4794fWVxeSBozBiGSE5Pcm4xJ0RwVZ7LcXe+MBsAaZS76LJDqnWLSwCa1z
Y/3gZayLw3fCtLbX+mCjKOw/uUOqa9BYwGACakHjBluAT7lUaMeFilp+KDZZ
xMt4TQxvuqSWuJkTaLeZ/wRBvq580rgXKFu0JjwFkFEPNOes0dUZxhVXpGPg
jbrOwced2wRkRvSxMs2rQswvS/NC2ui3kzJE27PsTZB6aam27lfoS6qLlJLz
EPDi3ZFppHYwVWd0rIuJepQvWjJRfMZQoEH9DdljXJ8JRbziDxaXCxA3yYVq
dDEwR98nEOVBwJgMYL9HPX4it4urdhyootCLmIFdYua+Qm6TTe7H8qYwubtU
p6r/1VU1BWY5R5RAAWbLYwa3tbxv9u2QQ8E7vTbSU+/FAyShHlEZCa6LmBAw
WeNnxlH4IR91zz+J8v9JeD4oNUgcz5wooMFwm3Jml983KFJJTg6jh/ZDQWsK
LUf/Cd6mPLpVQJ31CTFc8JPAz15OJ7CSmk0RpxGxZR1b3KnKOQZTdDhaCRxg
cpJo95DIVadOjyVPGtFLRcNCTgsjdBKTxRQeZYoh9gVc+cofFKXKuNdwWnCx
plAMBOsvvysrpi05fR8LQ/5Uc9rbsNWzeAe7w75DBs9k2ykRHF4lqDzxoShh
H0A6ve40XWeNt59mbzpvyy9hjLb1Vx8+7C4PSb0LZjZCVV+0UCn2Xl4MVbQ3
q0+7hk7/zSgc29fwtdSWVP15QOsJzq9OSAGh+aj26z8mYWVfdtxVeDfOEF7D
Qie4t6ij1Bwzv2flNt7fQDj5bRUOy5Tley4uTBrVJTmBOz/5ORMjCHX11N40
Y/3qhkwHeP0OHrY2uEZylIzIQHYNDWNw+hTRBwldIKFOsvdLSLHcTJ6Ab9Jf
8lDvB0NHTm8AK6wdI9FAlo7W0mI4mWSaA7hkgcPpOz+6pcswZrHQxDT1bLKZ
YHZmlD7mihrSZ3JfaHs/waG72nf6hvaftg+JNX2dByRp7hWqDbX9Yml0YWFf
ELDcTWkgYzwqE4szsYU3vrEiP5q7P6KK5axu++uLypIxT10xnvrcpUNUyxXF
eey/oy5h275IGMX/nrGO1DN/nNqeD6Dke8BwXtp6M7xMgZM/ESnskCG9COUd
FeeFxpOgc+JRxY0eMGIBUHzwzhChnbNenOVJcE7q99a9SlOFnaMBNc/m3A6Q
BGyGUbJ6rlSa7ARilFTXWaTtyi96BSnBJbGA09apOSVH9G0THwUttWeSNeJ2
g7c3bRE4AfJy6rebsqpQL+QtbugcdEHD4+tMeM514s1VAx6NtewbgTF5olVr
KeqBjiiB12ndzXP1vQInvlqG35rpp3Qbf1ndawaAl2uBsYjdzM8Rx+LyBkeX
8NIzunk6zWyC8tfyqMo5zKmYq9XxZ1ZiszDOZGktmM11fqIF7ULp7/J9zMbR
9pQ1i3RL1Je0TivL+G5poDWap3RNoSvUVjknG8T5Pon78yvR+xppUuXMWwtm
SqUQ+oihsQ60RBdB7C38/4YXenxoC/tWw1L49oPKD/4KncaN8gvrj/eesjqP
+Uz7guT9rMUUU2Djv6bfFEpHlxdOnXSmttCfwahF0E/oAxtahpYh+Xzsp+ye
yJt0Za5LKPDwwJCgCZIkL/IZS9I9zjW3W4yqmKiZIyxfMuyuFVH1dTFBpyiH
yhiG+Rb8ruMzRzPR2azHQ9FBj+vNbsblgTph5NKEIk9PtpNURrMSm1/bYnxW
ONeMu88ZpN09I66r0dz2EiHie3cIL+HRONmu9BWPPMPsfK/F1PE4bA1dE7Jk
rm0dKERht0gIs2S/wpfo0XoS0JcOdAikw7svnXtYYhNjccL/KNtIc/YP21t2
5hGvoPPK4pLu/b7h+viSXFBQUInk2aMl/22A20mOHMK3JKPeWNqt5uEndgs3
FL0JM0HPIDtw0Mbjcq+/2RQrCA2r9k/ua80cHuPBRsAagOomhq3hTHGDJrKm
8D8osDE/oS8cfACfYWjH9MORCYhJPFX4Ibn/BIjMC5aqWKOY9OdOY55kfPrr
MyfzQSZqAO58JRDyOrUb8GfH5hYbe4SEj/7CCrYG6NyDmaofZ0eOA1EOu9QG
Rqb2IZICSX/H7OE0n1dJz0UqHqYI+8eEfBwpb5sHxd+GUAZT7O+dMT8MlVmx
8Tp5s0FIaqmY9eDuFz96FMnb8FCxhTuir7x3M1pTtqMmDJ1mAyQg0bYlyJYC
2DwXVe69nX1KPvvP2cgI/Cqzt8agGMcXO9bd6jLGCJiMa05AGCN08Rpmcx9c
xvto6KA1YxD/CRwQu537GQiW9iHZ0BcAuxJasfLH+4rutsDVVl/ba3Ab6zi3
Uxuyd7k/FOBnI3m0RW2bmWnfrOhL6R77tVptwPFTan/nSaLlekxK62fxPv+8
r66OaNpJpNd+dyOcju7iOp+i2YSHm6mFyxcIOD7RjFUi1pSMCZduVrVFSm04
hi3fh+E9MKeC5m9ejcY2ixh8FBFh9gZEDmUf+Q49JlSCQmnX7LUEMZ4Y5duq
bwhdLcDRE5+bvZjYtCBH1KeKrI0mP5xpm08OOzeB7xH0dqlXvom1Ax8jrxZB
CNpBirR4aTn+ajBzsv4allriUlahRzpy1SaItScTfvDd2EoF861+kPMtZNyK
cqXNGtBKVyTQbHlAGe20S+SccpzQ6oAY14uS7XEk5jWJ2SFOxChe2crWLTgM
qrG4w6h+On9PFjgrGtvI+QRqgfm6sBGlZQb5jRRmVP9Alae+2qgjy8WqoRFp
qFQmRNgR9L0jyid81ovLkicbk36aKPTzJV/Pe8nnu0AwitL5vXjXcOTNR1lD
vuKpxrG+J0//e1gMnmhmxNQSleUXCkG34lwdmzGRAuDF1L6RlPDnB3PidKQL
sFsfBjs0lnlOgupxxMtEBR2Pe6xGXZH7Ov5aDinTDQD9OsCLLyLQCDziEul7
BjbDvKq9SQ4GguyPUmmbor13ObgojOs4s6QlZWLp7vp0lOUZoOg+Z7qtqGt4
ZJd5AstJim/e+tgAuTkGMbTZw84UtXk2/nNAoJaX/7QzHt6thuFQogUU8UXY
ciAjEkVDRhJ6WIjCvXV5j78f26w2u5hSJJpQd0e1Jg02dp/fdwfG6FkEEIPi
ycpwURVBCIc5fn5p8jNuKFS+GFx1NcWXIY8g5XBnrP3CprdsQc3w5QZq/UAz
lqbVXXRDKX+wAZDVvXNvvwQlCEULTnXTEz6JiQgvlgqOoia18AY1Z+RCGeup
wSwbQrByo7vJbD8thDV5m8RDUalLrY5XdeyvcVsbUPSrkhs2eLsGHveyf48l
4wIlJTpNfgjP6MPQTnc8CLcZBlqknGxVNkQZc379EnEgyerlxQ3Zc5LzbzXZ
UvBEFIyYZePjBw97caZxZM/DVsfcffO8x3F5Ia8bVPfy2aszzjPjpdstg0WG
1A1ZgoJ2fEzAL4AOGxuFgLGrIRCHaUHpZQbUsWDHt1TXyH37QJCBFyALMzXo
ImbwklX4ZnHkZAthOK+40ssabVzlInyZJFZxNl8PWNiewlxhemd5FLyUqx4R
PeocXS/OwfTp4jBy3ZW1I/mOBzObCSuflJR3YD49oXWcpZttcVVvcKqDY7c/
MYUb+WMOhPoeLUh3vz/L8WJBXg8fzWzGi7PixS6gGZwb+/T7kp2CJ/Soj48L
04y5Y+ZrqZPNmaWzSNYZA6G9O+4t8LOskhOYC+3nGWJG68vXUfeABjF49Qe5
fzW+UCru7heNjgZNLKLy46UkEZN71gYO+pZQjSjEeEsA77B25p175srVhHue
Y7rD1SI4/Di+/B0xLFUh7xOB5Bxd1vaZnyc8pJyqP+Nc/56gfx42HC2X+96t
Ok1bXwmIkS7EBJBrAqgl/dOqP1JP8W+pRWyiF0Z86OV984lVeKpUYORHodhw
JALOkX1ik5//hoStxQ/tuXMSbYEf1d15l4oBWqZYLi4gcdCvPWNHaXptrVbr
dYVqbPhYd4S+af/1MWK2J8FGXEkzeVeyqSG+pRuMRlZbbS+2oDdB+cO8Eexe
Qw0NlQDhDHdZQpQcH9NfklTBC+AXBKSrUwix1GPU2f5axkYS2UJORjqlwXCY
aCMCMaEhY2nMWCquntlhCSsDj2s3dPHupyVNg7VIhcVcG8Oy35qjccLQVkAL
DCmFxbryyiQw7u4LAdGpFPyGP1ygaqhJurYYtTl2wvxaHeBTGL/mA8gwKNF8
VPoAaNCKDpi+Wgt50fW79uX5+ZOJOJUPUKMtRr/eVrRi/7rkaCfFT/YBeZDD
KmOf/Wl/UJWMTvWaCNFrAoYW6iGZHDlweQF/S4giFusJx/5j816L5vuBTY3/
otZ7N4FjcToJeFlTe+DRPqAYFVeXenGAkCDDdHv8FnFUe0XtbCoH+GwKUI5G
iz4DOFQXZV4fn5NCCok3C//CFznGkepKT0LTkMkOLSFt3Xtsc8qKhrrdT/d4
nLyJQkofqRa/hgw5hj0k+5pN2haduoIzXPa1MKdcsgZjHeuM5Z7Ak4nW9T8J
LYTXGEGBink1mzgvFMGNYuvJqQ/sanC57p1iie7vwQj+03ojeyVnuLT3hF2L
1I2M22SAyXhZhxzRnH8GSGYMbuvfpzDy1fBzv7pO6E6K/s1rUjEkrITUT8oD
tQCvkslvgMVCjtFZD7FTphCV7SYfN7E1FHgFY5UUW3fYHlaxk/QDOQqfIfPP
07+C6MjsGNFR0CJDhgCnqoyCmRd09cspa9oRP49Vqj8h/tM9qX5xWfXT/V+P
yIlBXrnQmYQQDheaBqOLpU5IVOOqCv31hSUoySEWAWArRj33OAftl0wgzR/P
VGV+jwA66gsJaQ1PKdWPJhbuSxNm5bRdQIRUB4epNhYTJn/mwv1sKATYsr4z
nL564bu/kWfTtq5CWdW9+SuDJ6tPx1g7M4oNOr4b2JWT3mG/0XIPq5m3E0oY
u5irheesRXajSsjigapFmskkqcxUErNCQUrYkPpC570Mpb0MXb6SYO4JuE+R
ZbFHTI3H/ooaXWBd3Nwo3YaLh2/tFrp6OjyHuQFkHvL/FlqVy5zV/7P/Yf9k
7FGEOM2vyfKo/lRRKhzjz1kZ3mBGUU4+hCJIhX7erJ7SZ0eL9Swhga9Z7OrD
dEF674mJ/uGks4SOnUSe3pUEBx/m95XLOwYYaYNCjRdwz4miQbfwQIfZJvlX
3zyTSkl9t3rpypSMnhpo7OEmLWEgDjUa5Z+OSwSPcB/WZJRO2PK3eYcKDurO
G7ew4sDXRr6iql0vcr9b9ZOBH+M9YuEkBfopA/smtdE8ACdzp70L1IbU/jcv
vuEH+NsE15rAwFv1mmPlJX/IhNHZStBmxWDcyZWrQkOBFRXAukjNFo2Ad5lm
xJ3/k86gN/2PknTyd1RO9KMcidjywZQGbnhsHwcSVt/5NZdGqcicDd//JSel
6NgmV3r230tzISus8x3LTcDXVThZHdvv12MvgX+o6w7fe4kknKcB8DBxRHL9
VRfUFm/RbSqtm88KkFDCqOJ4pUB//O78PsDtYasc84l7iqSHSK+6gT9shAOx
7Bz5+gxwTbjmiVT0zB6iDBWNepTCYMNOEQCy2NBdXxMz+hB57p8WQ/QYBOGe
jUJo5lb5THps+zOQ4TlrYhzQRFexy6ndxQtXV6ivuZYCatBvXOB56jAXduss
DkPGBMQb2MvbhQciWgY5CjKcj7SSnEudUsKrkFg1p90kFIZEcM1biQt+OrSH
iQCC9mJUcUi6uJPiuNbQKX72Xxc0fLX9Qy+HSpowrlioYzxZBRRbV3cNovY3
5ieXE8hTI0TGkMMzZcC6Ea7koU3mYLc5jtyNJkpzxAT1UGLWbVf4q+sCL5yW
D9O2sUbdNnDNF5sBdkeLD24fcwB4rySb+ilDPNV2OPgTQSpRyQNWX0yoB12K
cw4/3OogY/MVBBHSqwitgO/z0pZaY7hjaLmcW8PGAiuRMpqeoNfB8IuDZHvw
8+4+n+KfIQmxcsKxGNp8UjMzUpQsIx0cvsbrwziB04qwnBtqZT5mcBnu5pAs
AXNwLjrZinYYTQCOTq9/m5OwEVa/BZVa3ss/KkGpOhCDSMPTq8rTEsOCkWq7
bqEpFG3RWVJO6R+M5ER4wuLJKHshN450pdRX8c4SYw/dueXe/aG5pP9jcSA6
lRATM25Ijsw4sNJoE21uRduA0BLUg2otAdjVmGrOTHjXzhIRnhm9wu0JPAzB
GVj7vWnb0qE6RGie8yKT5CjS1fdommr7t0KszYaMGTOyBOVQYn9PCuEaVuYm
iMpbvJESlWblD97WOOnFOaQXaQYhsA28pQzxNTf1/ouZyT+tIjucjxvjfV5n
LlOKKwp71GyetAW68GvjCpqs+5H5VQnPpURXJ5d/yOVt4FPG0EWKMPQF5nC8
jbenHrkm6/61SoH242AET/bzDQr8G26WsB6SHJuExpgnCmMp8s1gYE3kky21
5LuItVocOWgcTpz74MPK9ZRGliZPmWLi8oGEtUDcBfK6fPCCuxZVJJGiofnr
USYqEHSLtO1V3hxKngOllddcep6XSJaDIeMAqqiutJib64B70HSpKCjE6QY+
vnwvPBksA5uNtnFdr/Qzhl9gzJa8ecG3qZaU+ZHFyYnxbl7VCUb3SwkOR1fv
XH1lE6dK9J1cqMBsEhcPMI7fjs0Bef49PQcODuaruDzQVqTiJ5YA0Yrlb5gv
lr1Um/yHI59VK1sQ8TmbvynroqtJBg+FpyuLqokFnNjkyYMWSSJvc3xxV6MW
hs5cIyB5Z5GtDcFpqq4gb+CelzrxN6TZesE2QJGF0bDGXQxbvPezk3PCXOou
Dei9ok+XcDbNVKN1wqU76PafXuTo762B8bbhXsHV0su7bg0rzrqmdv+Hg6OQ
SzHpxopp2dM+vj6wjKGNzED+jlGiIi4OPFadz/nSK55JfqOtjf+v1Ok9aSyP
KPwnOx5bugMywxW4ly5BbrBeR4kk2YHNiTdteMliHEJBYs62rhpMD9ooWwbH
VJchTOiJvmMyZWlOXKn56MLQRjez3DlBBcPKkeiKgCwbLw8w1TBXWrEBINWI
noYIZw+yxC+GKmZhC3scYJo4DW+jmEdsqm+7jkZYDZ9Ih+xHwJDPUJcQMd2+
l8lubSoOkUZCkdRqWffG75gUUHVQVCMZ6szrh40jvlocYzvc0nvt+lZi+Gsm
nUR7INxeLhHu20B0SNfDdHXBDbPfOtlOk3OHp3HaPOugapYF/ZtZEDBxmGN6
CLsMgznwdRfVkCubMFCPQo9OgRXbBihU/PMkGU3xEoCNiGF48dGQ5I6tMdwW
7jcZnwIqK90yKnlIKIHlOZ7DblBL6cT6OwTegMjQ4TylkMnnAV8L7vyOgfPt
WZCzsnC+pJFrbaLU7737V1qxfGFpBRE6/4iuJFvZkH5iIl00rWB0vyhDOugw
tK/emiYY/f2ZMuwzopbmOdu1IvS2zif1/A3aKOye4ubgDmmAeAJvlTwDGEnI
zVFGyanThz2A8aI6WiL9pOWjsYSq0p1Ztei5S9Ey1ErYh3AmRmS70uDB87wd
KwKL6nJsz05gkcHSd+RE14hqqjR9JJoegjWmO/TjLsmVjZPemyWJpYnlriD+
Gpqguz8KZ+vEcZJpUE7TTQWCtC5L77olTQvnLHDEcADQwblTNUfcpCzFrYJ/
0NWKayLQSMQFNWhJpOTveYCrgm7eeqAgYzTIVt4jGN7BlysT707JeNixsFUa
KgdO1b6le2i93fZh4EltQaxhY90lWyYEKqYcYBVgl0yEKfMMjjHvfJ+nBiwI
z+LQqKwJVm9TtFhy7f6jXQAAAGnbneZjmYuAujmC3BKEmCUQH87XsOwJTGrg
wLBBK7+I6XY+spYNQex2RFwJVaagyECPuMKQb496OK23N7Bm1F1+pMTHddwu
5bo0+8LlTrmPNP6s1CXzqG7mzKDvSiFTLAPOMSBsCO4gFkEGcu5sOFjfLjG/
ykwIu1GQdKTgMmCVR1AilTITSlAByQxStqsp32f4FeOKeiRoEHgqxBY4EiRp
BqV4BCGuoD9V8SYDjMc7wge2nHBJAC9NCk8x2VIVTcj+TqKm3OUGiPtnmUP5
zUJBLBjRz41plIJgCxCrVwtRSP9e8GGqo4XUXEkXWbIIoiuk2Dq4rce7nXC9
dRZmrHiIoObvxO5pYbL3cImBgN5krMKtcChD1qxcRCw7vzLDyLbqB88RxYCN
gzlCGQ2a8aQn6UrW4WdMqtO9BCCDm3KvGWPis6jFFNfcMc6VYBaodmv2qaxZ
jesKJ6xBfwk+dE/UVrb+XfNY5g6BNF2tE4ZLUUxNnQT/vW6cX+XZU2F4SCuH
N5dd7rgUTA5BP0akMqLSkUNqvY0kFv7LCMwFEzFqNxIyGPiXiyk1jqyMoSQ+
c9N5Jh266fxnMBOwrFuuu1Bf75B+QLgB4aVE+4B0tfiGAO6csZzG8yzyVZ9W
kSwBvK5SaWsBwkRnraS4H+qx0OzPmh6+lSBsUCyT79rbvIk7oyiW6FwjcvsW
BRfKoZCasQfssLYygfN31QG0xMzCC4wncZqX3wTGUy7OTh68AAx7QMnk78aD
SE2FnYv5h6gs+2D3MFao4AIOAfWpko+6wPI+VXFXi5+IG1BrsD3aMgZDcSOS
xhyHTv20X9zvS8IdoAAnU3qiJLMy6mFlTB8dWjnyPrM8zhUdVRkZTRFMs4Zp
nOJBgF9c6BHlcb4i+uAkb3EQ3qp8w3dbhO9VRNYSJql87bWuDGjHWfeydXcv
FuLNNsh7N+FltRorBMMIJfExY61KDxAkk7jyv1phGxR9V0BkNeAiB1/j2BYb
s7OHUGswTb3TbM650SqB0ZnIx++zD6lfLtWL18+rMcb+uMXPGOnq8xhcKZY9
IxgpeA1NElNPOYvxq2S5r2hjWKfEmF0uXA27ZnQJzmGwebpXEn5EHylDipN9
9qO3ydYtqe1Bni6KLnmOhW9faU/fz2UNYdGA3bPd0u+oOJ56GIz92qPJpr+8
N5MmZnw+eeAbnaNM1iKL0R6OA+bckga/xPK+w3FfEIrcoq4jBGOKSpFhgIkN
yhAcJfl7Fe8CrA/jkXWX8+bWjFWCYwx+pl+Fx+AGWoWevceUTJdpE3kQomXl
hlq4ue5QMLgVCf5U9tKBEnm77cbvXgXx5JilUqsNdnpg+sgtqyBuqxzG+nGh
YpRPjhXvOoGqcEj/UFOJeAl8PuiJV14Ufm1EzQtN6LIXO/rGIglYQ+C3Mrqb
3/NEggU9a5Y0vY2oc2alsfSr1GZ9yGU42R6yO1+K9P9w9Qbsm+hymV6ei9Kb
Fy6xALgTnxXDy9JTEYt5KBuSgvJnE91ZUca9lv6BvTn7BUVRxgNnoRRhS3Dx
emqWzwPfNKO6gUgp5b9wMrH67P3qUDpxEUmQdH6OBHafob4yayavEoxt3N8n
nnJZYy3otgC0HFu79j4jF2NVzz0AS1/t+ylZhG6P2loeYzLXrE96Mnd8PAEf
4nyWebPsiOiukw6A4GwlwovjYJTwlhg9cov/dU94so7eRIoukqvYLDbqk3TN
Ce3Z7rOaf4n35Jp6Pm+7ctBy/uE1qVBzPP+E9wa+w7GtrGfmZp+6Tk0XkIlj
nclU4Sn9ggC736xOaBa1VO0DbVo8JzBtjj7Hr3dY9TsZ4eTCg4OcWN6oo13v
echsuDnMyQH1TOdKMp1BV0Tl07sJrNKmBJXXAGEFCN8dWUXpN6Bgs7ZgNCKq
xlqZLESMza4j45rPmo13BKrh7k+HVm+ivoar0jmGaJDLMIABQe64MLDtUfTU
0qGQgJ1q1iWHNP0sCbouFuzV7VfztNQ3ggmVgFnAkiD5rI4rJb/Hcu5kpMEN
kV+jszcCc5lWUr8cfdUhaC1FvqzEk563hD1JR4MI4gXN/hyZEZ5iN1m1nVje
zTnFKgican5btxA84wnHT1Jj9YTUjewHWPP+l3p4v0HfBP0acVB0J0FNgeCl
mbA9Fk06uBZ8fEG2X8RhB3Eue+eZ630QGsaQR5AJq3yNiHTSGevogkZ7u/JU
IF6N+0ATiIcTfPaDB0fbko53WzZRat7MXYsbm9XBKiS9BrABbO5gyI+E5Pps
gImisdnj/XoHnkN/1YwmdnHsFLPhyxGFBOtC9C01Fck+ox1skcPMA4P1EJQY
j8knqitNJdBlF8UId38DiFfd+5wQThuNxEj+rMjxXcbmBM1o/AVZjs9sXD7o
Mvj4puW2EWjWUs3v1jMnw4sedxtR7QB2KcL6eGMgxArZnotohz9UAa3c7fuK
gihagcl3Lwm+HqN6m5zHqEVf5l/XjnVBJycG67DcxnnxOE5PhnYjPqNG2ATO
7EwyrdVni0x1aTbSaZx4w+L5SBIWfESnjM1jnFpdLwWCUuaDGuTx4C4v9jIE
SfHZ2CRrRIxMYUY8F9JmL8jFkBsJn5gMLipbfQr0Vp6uU8CcCoCBu2K677My
axmd2rZ2liuWOf2iotCnl8fZnwt+ToxULWnY2Snj6IQschsEcaydwiBHFjqc
H8IuEQLUjiJKOEd1W5NlUNno6xdaEik9NFWlB0U53RkBMMh2oP3bkF6Yb79H
FWempk1d+XebcZhTA69NjWTf9xGOD2UxFcTEpxaan/jzIoV5QZkpUaG6Uz1W
bHZ48Ek+xNAmpBISOzBQsjjB3vU0YaBvoJdC1f9iAyOWT9oVI560hGXhoQtf
BYpXR7ddmRlxrUlfmCX2b+/+axP0/6XEswHbVMmfe/ewX8V3FuiIqfftzy98
EhxTkWetA0z2YEHeHTOYVgAdLM+AugwsD1JQI+10a0j/1idU6KXD5ebjaF9x
yzQYdVtJiKGxQxtkQxFFny/FPaTS/1fdg1ZoWokZl8R/ytluRqGujnG0c33P
bZz0HnhzKGF/hc51ckP5imwm1gDQTV40oVwl69Hgqx0vDQQh4xiiDyrEhkP9
KOnKQRl07A9F0WMaK6t/4q45XYOXlP1A+PGkrGx4IQtTl7djiCXEdihQaFTS
2tanxLI1PAvA7tcxOdFR9tR9/YTwdSs3obSk8HfLIWmGYR+cw2bqIjfeDP/9
mpTYu67wv58Ws6c59bF3WdMuODfHdTZTIp5KiQG0CgFw1MQrkOACupmHn6nV
6iti8tkOkoUTlHVzU6OCmy/qv07T8hqgJk2p8O+AsoKIcNZnzc37lLoGn2/h
G5Tx9uGlI3H0FtTl5Y7TqlmDceaMF/IXjeV+LemlTt05U/ZMlvxtVBwXWJBu
GO0lRePcawIpDRc21LtSCLETGZv3AmGaZqSHkobnGl9iL60Vxy8YyNw4d4eK
aSvj4bywTA3EEInOLfa0oiu/LqR2Hs2HKTESD2FmlgwcC5ex0gHdA5WR84y4
y+d736Ah0tGf9v5U7ijBlufGqyO7AZa6ZZ6mCLAgXukMauNJLIaiNqG2NsTB
/caiJV76+t/uHz6OY4eGrplKawkSw26IxDuTWFX1vZvKgWtepCnpcULq5atU
ES9Wznfd8mIa/ApjqWXyMPW7txIMwdWUVKj1pcez+/wdcpMzNhTV3fL4yiLR
Bja0cV0zOoIDkZURL07kBnp5xPIF9W0wqlGzPu1EOkO8lXQgRQHoiTdm6pIj
sl3QoDFrRszdKvRG7gLULpKl02UCoyghySZKaYbUnP3gsN2cJ8yLfJKppC1G
D1NySKWhUxeQq//Pt81yOBmjir6faNdhPjVMiH1Ai3D7reh+g7EO063slQ5Z
UHZLqXFqRJDIcUES6cU+l5D2bXLmLi6jp3XZ4WoHUWc4S27gPUOejdsnsCRd
2lr4edchLNHexa88MrhlmpzLuTdm4atGUIub+CTFSSRtb0VYBd7npltSMkfk
go7YdghWfAAZC0v5zfvUzPq2RsWt6o0kQssCgWn02fLdnwIOH3VPpR06nQq+
3RvF4pUqe3BnKhYVwr8vUbpg9g/xNrdjvmwFAW7ABi3iH25Sjcryy7QVyvuW
LCZSeWlMCAmtM85U0x2aiAdjKv1rsR3XK02aSWhrnZhGO9gMoiKC3LIwVUAa
syRPI8NPqCX8tsDUZXjcqt7nENrDZRtURxT+8iTnnGy/H2/8e4ExWfUh3xv+
r0n6LsDdlvc87xIZoU5ey0i6yRpNp0rHoiVWQEUIz4B6QbPnqWAiKohgiqar
in5VGHdnUbicOT3WITjZiWJceOkM+wTLUBBdDHCLN9GlvLSlJeOBxgfoZPfU
MLicIZRZRQ33v4AUkEes0KitaNfrzzAI/Iv+CQD1Go17cZNIAMwWyxBGI4vT
2ZFKBchyFn9eB4M1u48+r602Q0ktyxJhM6o2+mAYR7TA1q+xosT6wfK/Tkhy
kz6Se1XNa/D/NWsS4CE7ZOC619OSkgEAd26d1vQ273fM2/FSck7DITAO3EQ4
X+xz9j8+dWgISBcORUFmibSJv14tcM58G54opanoQpdlZRmA609sbBVaMFXh
I7yXX6ZCN0swsPC/eK9cxNzmJbZHm7Kvry2YGmfhxgBP9TXdLZgzhIEeJrrS
xqGCEaM9JDxUAoAVUN8pNKPnDtdYbV7b2Dfg0kL23SueWbdm5nDmGKuWbKUR
gFD7Hl15alZF2czaGfQOhCovPuHXL2LQCBitCBFl/3olgC1l2i5v2LkZmb5T
LJOk0GO0qq+/1fzp6bXEnr0GtadohE6feUH/N5cOs33aLV/H/jhppRPpali6
907fxnJ8KXsuVp+/8QCag1HIrLF8BtHxKrhx0Omp70JcjqBCTdshCQywZHV/
9SihIwEwLsFELxav7DPaH4+wo8JSLJXoHKwSkl7JrQmz0dymklPTupE0KqFG
aPRjRxyF+MqXpflLLEXWI7OW6rWOl+t7ddsInpXoEnlrmghW/MRkhVJevcE7
6GRX4kQme0J0HMfrqgfLg/rY4Q5bY9TGEByH/Q85LbCegRu9URpcy9AvUDtM
M51IOJK3jkRxYH/KoNHoeF6fjvLH+Dbafvk3yk4aeAi/EKkBQPWMo1esGlAQ
BtoaUFcHN/Vs8+3hP49aS8Zx+lTzwNj+ciKUdbmg1FrTKf9fQUbGWAicJqw+
JBwrHGpvr0VUEO6PnxSrhDzVd7NlWb5lbHZ4qq98vjPpYHdG2JlTCnxZFFPA
/447bguNMrCsudRZfJpRHhaZmyS7itl67qy8JHg9azgVBsImNsnkYtc690/7
C2ud1OmQ04leScWEcLPS0BYDPJpq8gqmvzBFSXkCdLYof7fq8O1VG7XRt+J/
aH/DoWdjnoWmiZGupg3KRsM4PMk8ityM2UETW+JvjwrhA9vyuBvZUg0Uvde8
acSq5m4hHTKCQFFsWnxO2b7wmyNlPJYCios54h/mLy0Wf6+yzLv6brStTszY
+Br0sPN+G6yG1tfJEPa6IbewjP2vsjoKzWG9Hyoqi6HEWDyVCpQAVv70hnr6
2J5u5+0oecpGBpbjiTnHTNAl2yLL9WXbLT4ZpmZliGqbHUBJoHQ6+TFCoYwZ
Qlf51v6vID4gy1XOFwHhfSSiutoAgYXPdG/EwMTqMJCu5ufENsD2ztoeT6vK
PpuA55ISyTuD3t4QtzEwYFw829c5HA67+KyzjCwKVZyv3XRrdpANocTz0fpi
sQlRNsmyEriMI8oYpI6uHJewZjMtTDlvGPlwHWZSc5FbLicvSQWQ0TH4Koj5
PC/2ZLL/QI2S/1oMpgbikwxw5ZGq7x592+AD/eBvyLIbIdoIIzIVfzl0y2f6
lGX/Qr2HYdIQVlsvThGUaS2nvPadwpsyIHd8MEbsVCBZknEUZ408BIS/8Etk
XWviPgrea6iRDJxF5OMphZai0BK3vc/S/LXSuyKgZ/2koyC08191PP9HtUqo
GlaZM9I6wMuSzDqomsWN1/6N/vVlqOO505EoSj5XN7zernzoUMTKqHbCBwJz
r70nfeXxQIsEFP7UgYS0VKkk4jUxiM3BXFaZotUBQtx5cj1ch1ImLeOY1Dk3
Kkm1WA+3y7JSLozOsxTQfZ01vuMIUPJTTzifmcH0GFuZlRn2ZQjRGBDQXG/U
BsTKLatOJMiSANqY4rQI1XMt1KoyOGDm3ag/FR5JVpN9R5E6Se915NCId2kZ
YTN/MP+2aoCdjoIivc6IOFyK6EdPpG/5oynVPEcDBgcXnA1Le1LH+qaVIFtf
dIVcVh06LfAKxpj1TvY29DkkTIi2xnvsZ4kcM1BKXg+9XFZ04sp11OH6s1dN
ykaJdPnj3TN8Uy9RDdzZ90VfuMooKtgb+9DcDA59DHuwX+q6E0BjtTVYkisV
SgkrhY+VC0JE/KrYdCQCT0UlMxXIQz/9LKPXhBeAwSIQDl0CJjAcwen6fk3X
Of78EL4O7Fg946gH2XL5wcDtr+CpVGTVbHXlUg/v7ZAjxgwbcAlzqOpdNy9O
zInJgDdtm+fjJvNngjHKVREYXXffg7LwCPhK2Y+A8pC5qEh+Pja/92XHfwFR
+C0Di/e4fBPk+k99L++prCkHzRmj0bi+WJg2YNfO8RC7Wcd2VAUm3CrFGERW
rrANiJ+LxYhhMubGhCA9LKoYZFKT9/NmKzmLp2V6zT7QQncyt9QmgV4/0i1q
HQI9HRNMU5Auu5/JdsidBDMLcA9Q2T0qPa9MV2OOyfX/Tkurm4Hwh4vh8+MF
Oh/KT65AyWXPUIlIFh2jabcCoYiEsb7qZCokUkQxpN/yelbLeKtO0wxtybFg
4pCycs3j8o9h9a4+q6ZKBgU2k8spJC2bd21kQIjGYPUypsUyzIJYZLC60Bl2
goLYukEQy8KcjmDdK8B2VJGTcIaCf0jM9hGyw/gBFnaqzDru0vFPIV22lisZ
o/KOd4g/oFRUdWgZP3kDCiIIleFyvBFGfuoZM3FCWVwUXAYvx2ox9+4mPE7j
p1RZkcwetg0tZV02aFCsYaEj3N94PByCf+JWEFCabPLHQjnw28nM+Uc/YvyO
Hvw68oLSUJCBrfufY2D/Z1grpGzv/BM4ujNwhQeDhytlEXEyuoVGSPuJ3YU9
/Qbw1Cw4daaYlT8Z0fNnV0KLj+nSzUeZ3Hhn7py8AAs1qMsW2o06Cnu9cDW8
Ak/kFwrqaOGNuWhU6aiVKQUO2n6BZLrUKFtWE4RY6wmMuG4jqDRMrf3p2Zw+
ZCrfFbI2BPYVnnZX7ozB1hDp1Fo530CByfjwfMuLeGxhoU6wlFtQImM2XR60
Dmb5uCRGiuq0dkjF6N+LF+S+DNGoFuAP83uKZYO581Hc9TWlHyuB90Fa4cE+
yZfi4g5ykXeHnzg1OsGvLArxf/fmRGpXNNi2qrH6dI0BtouVoDcf3oWuYOEG
QkZVCmVIBkseQUkYmwpwLYNjiZU4Fx7TdW/DyX//22pQJo7+wit8/1PC21c9
D6NOqWB948AXTsy3wGjgZw2uySYCR25mxYd0SH1i5xf9r+TIvdyxX4dX5V02
2TP4yd4QaW3c9FZpVxRfebrx2qTD7p7v9E8d28/PPA/sYvsbGpdbm+9JsDz1
ONnMW0i6xI2KpiNalJCrq6mCecMrhHgXftp/nEFCh3eXAyP77CQ3MBFacMIy
uX0rE80LFujjlPPR2gA6REd0G5sf/BZX19KLnLOGo5WwO24X7cQNTAs7PTLY
2rsdVI1mz9u0fqMoRFoCCkSWFdgT2ZiW3bVewxN4hYWigcvgiM2UPDfZRoor
4yWHaVD7rJThu4HIDHdVXyuSChc7sXpJ52IpC1VF3Mib/B1v3NXlS0aVm8Jx
t8nB9sBLSzbp5sgcX5iq79b65Wf6lgU8T5jUsfitqexg8pjEkAnepTx1jPqt
1ni9IS//5QwwzLwVXk+i53VYEo0cJshHqZiESh1enD7CygHaJ5sfzgHhN40m
ss6W54Am1Ps/bYDeKcih2F8C3ZTAM1Tfc1bWwop6YB/nICEbZMpATnpaLJ6K
oWc8ilmBQhcx3NISq8+9pycoCuuzkgvQUbbY32FEmC9RBE6qQbTFBc3KAMaw
pQds4ABf0wl+DmLZXxfFMLAbseAJ6BTKG7ocsMKHy58In4igGLBRiEGQ5qL1
wLDQ4JgFn2RnRkegGvthUsnn0igJriF291Zw5V7Alc7Yu9nqqSb8APDCnl1R
ah1rnwm3YgmpE45cecLXeXeEcIc/j9UOdYSbswNfepAmb4qvzP5/Xc/bqukv
8i+2AdVvLkeJBjeOexfbsjxFYgZjNHoWvsCsqvqqTIWL0fKpviNHd5WoEtMg
0DIq8Z2CkTY/qjYRFuKInGj+q6+hgSbgVyuhAcRFSQtgXEgyjF2Y5TGLgW0j
lc7dE8aH9JTKv0eIsQe6ox/OGdi0oHahAoWS2gMbD3cDBfHTSAJ+Eg2gqVE9
bIgJV60Ej388SE2sfRBoXoD2fc1NWowJnonkv7JZchH90zBC9i9x/kAg6HVp
TIPw00xKWR21lUPD6Z8HeTjuJ3Izp5CxvHEabQ/xkeUz6CL8WS4y1KA1ULvl
338ATzXwffoLq6bCFuQRlLx1EF+qGKk2vwounfX58DwNwqtJPkKB6bbwDGyF
kHmrXO6ydvoVEDzN14kwacFp3i9e76kVfPKqBFicQNzvR8yoAOqQ8ZhXgdir
+vUR5UM0aGtuZ25b5LrXp/3JvrxH8SCF3dtD50peKotSCapAZ0MKonZPBFH/
BYW/5Mzrc6esPpB60Zvi/OXCATXYeKRV6DlGrku+HQZaFJ4Cp77S7MjVuYRW
OnXKr44nbEvmwSD3fTNvhWaxlcMKqcyFx6j0yZGaLXJRvk6wp6/BT1ckbULr
ME23sqKUGy82DTCDIu8QYQ8bSKoLC24YfvY4E8TEkAtFLL7VTUn4gyjEJvGM
NvGQmcd1Cz74GSBYVSZQO7InbiPTO9YKiyiYBM6+UYC7eFOyshff/y+o6vqF
PwR60DRgpCv8xMmyuo3mOliOa1TG7P5DGkC5RZveiGC8kLRn98ZnYAv/Ui8v
G/Hz4nVICEtSz5Nzp653c2QjxOUsmVPdOFZUCntxCXZsVnq40KzwkyHTZhzR
XdevMCS2twuPPEfjqUEeii+WMhq9DgJvNZ7KEgKibYuf8m7PktiC3RHiHTcX
6VlvdOWofoT8wMPGSMjmx3dbz4c5hNgf2idnqdxn4adhc7IxOMt6PyZTGAHb
f9RPPbG4bAlg1cOpxF4THIlnmcbOfykoqGVRk8hZdZRFbxA1DfD9M7yIfdZB
dYzu+dJ6IkUXuTeLH9WDwuwjuJoaqRXlGxEfnKZn/znOgsCdKhr5CkibBDMS
lm74SemKWrdiuXQN+0NFxxzR+PdubBZIhys01N3tW90Z+C7jRd8qCKxcC7Lb
2UEyrqqRSYPl2e5UTtUlCqONC8QqdW+HR+PbLw5J/Ohm+K4O2uRFlJMrs5eU
56skPtKBET91vodC3/1kKbeoAa7MLANRCpYmRd3UbrUFX/eS6tx5CkQUtVWk
FveIYPV1DnjUkJOqqHmYUOe9A+6wYlLVhaj7eQcW24Jxkp8nEtwXuhr4Isy0
XZ7gYcdAD7LMAipCyV9x6O5RiYbl9P4qOJL9JIHxo+fOWldjH1IsYHSkhmPy
Wja1DDeE1lXF4+FfJm/2i9SuyqjcrzMxOFSwno0XVoc0a8/uOkYGOMQj1m/1
HD7CwB9pfuKmBHeQMN2y0a9ZYHAaBXXk5X4vwwMDcSTTY/CZEmkT7E8fTIWO
tKt53O6WRcZF+gm5pKStcw6NJuKaws5dNSImUVJgpZmUsl0lvYDlMH5W+GQz
2XuNRy48PTiAo2I6ZfWkceWcwU2GtiHKARYpTMkn7ASYZ0X+J3fcKftXkspV
aBdqWzdlmjzFDQoZcGAqXM1Bm0T6DxBQMShrKFqNT132/Gu06e/EOK61e0DH
fd203IDQPGqi3RYgwoVxCfpZ1V97iczPlAcZNgVEbL8CoIN0t5FlJF3TOZPA
gYYLUFt2mTJBCPknkqWfM+kpXaUSoABMmqBogC35sD06kjNRXQzS6iHG2LLK
IUU66ZAP1Ar1WxfGXNdwXAO5Z9U5rxdudHGCGdM5yUCXD92xekzJdEa8o+dc
5H+q5pw+ii9JKU2oLW5ZezBcpoXuCcgKOZCHG6RNlwnSwIjUGw6eErCB1k20
Ly6E0tFnbdFsMc0KDLwcCcmjjxs5dtKYHgS0A9uHe7+6I1WAto1+GFzFjDzw
x2ThpB8cU/md+ySGgzD06ZMjgs9yKzHk5O+jiAriuIwNspYQX5sXpDZjwyHi
cbXcNm+VMvBNqC9DczXgqykyufnET+f5jBJJge9oiQdBaZ9Os02omwtJnvLs
8BvgSU25jLGZAQ+uDQxgNNmoVc1m8WvYQuip+q+W+nm9cKE5mkbOXl+VeqSD
S/QFOqT/T/4LuykcO7G3BkOSmCNqmRqaEwnQP7hDwzZ84lFh+zQ3YqMnAR1y
xDrhzuX3dWxgCn76gry1ZkpGfEpk9DKcOCLCQMGnbUO03XO5xAEfQiTYomx0
awy6LOamIfk7tnXGEemZBcy5ov1K5NPwTQLLLu/ojwLKLrf37xP8/H+/VXiH
/JWDJSkj11opG7CAER1EdWKO15GBF+g5LQjgh+8mzOjTufCzbUuZ3O6tZF9C
HbzmDogG3RJUoLpbohNNLMPf4hGLN3OsufFLKEpX1LfxOu0/zELgMzKXdINv
P6UEyogmhbD/vi3IgcTQYTeVNytCSVgaz9VlRAlqJEoupCpMMDErcfgujNMo
JpnUoYGf9jQbO2EbqKOqIGTlxH45q7Ex/KiiVi0vsbyDygzJ1m60zHaq6RTU
Xg8RYFZ3h1I7/6J80UHUQN/fEhLGot0NCmxFxFI417Sd8DKcDyinCk0Zr2MY
zswetx1xPCqmaX56KOaljqG19+sytZ/3FAc142yyuH+Ks0s2ohO+oiu0pbtT
DBCUYezwhtdl9NEvtWHEf/mPFzyEl0o6J2Sqx7AZzVnL78TiGbccurUyViG/
ZnLwMJoAjHXagspzsHMnIzwKljXSYMZQdQVd6NQzkHxWe9Yj5uQmwLgiX9Bg
Gmqh0REDohT8N+PYic25j41PFQJLobFeclZF0TAEljD0tSnVTJeVBfU27MX+
ehv1z3JG3EqKjqGQceo0rRoDE2Y/FY4Jaw/eR1dhxJKYoj9Bne6yuYYQgVlV
dG0xyqPxxUCKxPE1E8BRP59d2Lax0krgCe2Ys/HUp4bs7IwT1XwA7nElbAqn
SKL05W+srkg/iKUOhvBsyh+jwBRJWDEixyRFkhTpSLB8iGzOf6+7XVAutw3S
pSeVdzl5XhiZQTIUihh49aJtlsxIWW/o8ap18VWYs9a28/C9ufar7L5hOKLc
HrxeOE2HkZq5VMYDFJAfu0aNJOsm/xVhzcmPK85wKr1EjgLycKVH9ofN/vqf
NKF1OAOzWdY9eeiVSlrQeZ/4zq+8kiAGtvOYAeNXkpGLLwbS0aSWLDE+51+C
WkdmKcGrWqJtYLw4+7coZgB63fN32gyw9hyH9r4lGg3HiRvBZLqc+2JDG7Qh
uSQ2qDBQZNXKUa5g1UpS8tJny+30FukxidDq+19GzobDbmtPRFhEQQhNzRWA
Cts9ppjXkrtf3+RdQElpcKJEGLOb9B+y7d3GAMjTb+Pgj6pkknZ5qDn0sCiJ
ilUv9TnBENNkSCs7DfUB7YJIJhfOfYTheUAlBbfPhR9ggstCdXymJH0f1gtE
m50nBweJ9fJ/smALytBpSQj+zIh0fnc4Lkrcii2Aee+JEh6D54M/nqjjG2cN
7MQq+p295RA0fZfCmx/Zdl/AoERWsj2TX7hX1WuNQbzpLt92tg5g7O1De3in
+l1yzs7eltFCctoRm/lVuS7RhlIBeDEyz7J6cO1QwllL4o341w4q/71H/sVl
E7KeIlQ9p+kgFBTd8nTgat0V+uDktXLFZWA22YPTakeIAC954Ng5UMKJHq5S
orWZqbtnDcW/HSPN89Cjj9Y69xmPXnhVlkUeVIoXDUHB4LC/OJREtogLIs/V
wH+CTcscgeX6xen+P3bubCuw71q0uxh92Ns2h96ND3Wa5/uzFqDHszBWWnoL
wWKhNs/K0yToxcfS+hC+to6MGU7lv9M0aKYPluF+LWFPKHcyuie20Cd0bBFC
R9nw263yvZBv9ST4Kh4EGrA+fDjgFyCYiWgldsj9EKFYw9uVepiSrp67b+y2
FfjTovpzBZ1kTZ774S6g1Xw/Ha2dPFGR0B2hv78wDkqGoBSQjQgvZuk1nvwa
y2QgLsohZoP0B7Cax1VH9YSLc76t5ToVhCPtxHZXTJWgFHFZN+3I+ge4XoSU
i3q/JJmfe8maXCEuxPeP5oXhl47lhzvRe60ynwfZUdv5iuXehGSuMe1yITa9
AouE3j8fRpGVSNj5nicruLr/jnqvDwX0ob7YpLWUAf0pErRQMoxIssSZF/nr
sx7nhDT9xbXKUkR+/veau0BnMiMHkjkMoFXfbFnEtnBo70jYUEjO6/sGeFIR
SgwKGR9mGeklyWku+NCLUqv9pZvViiJELtUwhq4mAvo5GxmX5E+BFsG7GVeI
PxCjp5gHuOxtPqVufB2IfxBTU5epkRIkVOvT8QWXA8KomvE+HvqagN1MhwY0
zBwrip6DFZcBeV4HFYMfX2XhkG/91vupasyLA+z1DHSOLEwX90j9YSs8Caeq
mWDU+M7mQMAiEPUfKOXWBWjSMy/SbSeYVPypWFgwFG38GDD49UmlBWv3o+U6
svzKXo5yABd2coviKFXMTHIyIundV9Fo+OdGfWtOO9PbqI3CEyR+RqqndPgx
x9I+SuIUxLJjQxvGxD3MpmEMmRHIFfR9C8rrIZ9EJjtJbazpmsoPf0Y7B9Yn
gx7NdNFvqQ7uS1MGUvEsS35SfAfh3ejkqVdCPdkjwLavOV1R7DI/vONlWC+7
aUvq4mdGGUcxzgnTh/22g0MTZRErwIOJYQ/6bxKNwzxN590kMsEUOigjqYcP
YRA/3lL6LUORzeHrjVzwT5zwiDxbDsnTq6jL0qikQviRNvi/T5UnHQ56OEtv
0ldjBxwJvzauVesPy6GDZDl03nuE44eWhpr+ep3/sz2L5s+bCWBMB16GOgmQ
nlBn2xnTEl7H7EHIccd2lpZchkqHBNTbpJZjjz+0UyAfCEemee8B2R+SyAoN
bFybe9OeYXcpjFXg3o0/+ocNaq51nFHVD3tCq3VcAdUYkz+WsGbh5icRMM9b
/zjggGfmURd1lR5Xsk2V42PCKeCW0Pc5kS2+bOzxIKdWxN+zL81BCfUWn5sR
mcoxwLq0otL/kMFe7XVx8LMUdRDjDaGBiEBmKD6izVSKjHm8dsue8Z92AndQ
jAAsU9Sgmpz7UaMFLk9DUHMu9LVm2mzV2FgfxJHJkWbWOJ6qjBFmzqaUqx67
zMtK9lQ2ie4ZbxDZdYuvk5XQ8J7+LwhM9WS0aOfsz0QzOSoizQDSQGbRI/bN
DMKcHSMngnjzACuw4mI9g6K597mfhnDrvDCNP7B8w7o25xYbo+CMnhGrUqWw
fFzGjCNc3yERb6L/KmzlwvHVwuUWgOv/Ab/sU6jnrYVodh20dYPLhWlHlZXe
vI6XTCzIvTVYRG8dDdeea0AeGgNO65cDs7pGaRUeCcqs+23dj5jTZOLvUm0j
FzjUQc/ZZ0kD6k3KdXuQG3FTQ6/TPVBGIKUVUkurI944s5Lk3L7swmErKhwV
Fp5o/Hp/Ve8hQA6Gu4Zj/1u6hvpK4q+T8cFLcsa29TpBYtQ+D23w7kOc4PPh
9cskQAYQP0NWGR4MgijJU5gcZTfFpu1puLathBL6G2czVKRs4XWCyE/k4DwH
Yt8nWWomFMrEzhEaQMFq7TuXA5aavomjeDGOrDFvYU6v82jIBPUEGuNSliUT
he/2IwpoaT7fyWEziT+qJ1KerGqDMMgMQg+NZUqJHu1SOjHkeu0WoXXuOmeT
hksbb4qflTtGV2EQwFjInh7/B6lmaCGw/PzPUBtiVMHUv4EcYaVsvyfHiFFk
sCSG/qmIEtXVWThwPEsnGvyZaLerjU29sY3GdqR1ze1Tx8hQuJHmefbLpfUU
4zXnZeWvKcducqdN/N9lWCb+hDx+E4g5qaU1J3Undcn1J71ySm6QMmkfKw4+
8NZHgPjrmM0/CswwzcEZblBxhSfG1YGGVIUllcjKsSjf7VUGw7rKVSmBwnE2
ka97jlE4l8G5t8nlStjbURk//Ncbic7oOgJUtvV01585aiNDtIpCL1Ol1M32
/UUwPjAyCMVfsYKF7JEYJcSnd6fqk0klFLNJVDoiwtgG1kc8Db/PE1zqxdoG
UoI8rtf3kDc27v5a+tFjTFNn+78Qg1+oWQCmqBTvBIGCUhpTZ0Cr7Po4K9HI
eIg010/APNxKKZNW/5ToeLoIByR93XcZva8j0ft6Ty+qr2TWyRNxGP1rztYY
j5CiLOaC4GgxryVRt5O3lPMFAVnztqcWRo15JK872r2w0k93rbaraHEvSA6o
TQI9c+AA/NsFF7AuFRbvyMahSTChye4SgApWEnUA2bjLv2knFv/ifvkvmD/f
yli/lvTq1SrZjyIN/1u18vSSskbn5gcd+6JVIIs8b+RmaEk76sfQSmCumv/V
ehBAHX4fgI4NZdVWQtBFPcW9ZAqd10r8ow+G5Ue6y2niO4YbGrRFSzPbTJ3b
yO/lqrCUQ1rD/cootuxS82AyDqWF6qMhithosJu53L02rscaVmdSEbFLFF5i
5kkkrjwAntm9wG2tRXRnkb+NtHYs1u287BJ1w+C2anz9c+4kyRvx9CYPIoWg
C0w/bMbvNwSPayjJNVH35eE+EeWuxr2QrMH7483GIAGrb+ELuW5K3bj6sVMx
L+apoxfH2XjnCCSuAMNYmlLYHPAV0T7vujGcSbewnFnMGsrUwRwR8rlmIcFs
EjyI+spausR4Sred5aHKTyCQapZAWMlEheVXEuHcHh8Vbnn8Bci4sfe4ECja
8vohUWfR9m/AceUuYssyrHHEcDgPpLgVvfG4n84o5g0BmLZYDmgCyvuznm+L
gojghLQcOXr3kL5QiaB34cms170OmMAmNumj6PuqKxwW28MuacJQgiETwkZ1
iwKLZDlC4mHimvTygoonPsIF+Tb/Vy6eXMnpmuSg6CgqT4qGNQ5a/Q3E91GG
bVNk8na4GpEn9a2JjtKMbjaEvxrvS3N182OCLUccUTYRwxTZRXfN9XsY5m47
kGQ4WHkf3AXaNZ1eUqoN1K4UBrQxQop3l/0QpNVA7M1N3pVZ9tFmzGPsNLV4
1ELvK1RcUdVCAGXpeJxuNtTb2RxpzLXFBvIhNjx1C0+k8pNbP4HDhProz7/W
rIDQpemJnsrCLnXd2HfRQD72cLDCDElbGmr3oSFN++8TpiUQW0BQfqZGoIXN
AW1tyeUhCpg8csz/ZpLM0p1kZTVn+gTeH8ev2tGWsFH7F+TVbX4f31KbksWY
1x8K+I+TGox/+IMlMi6rnsfCRCVXuxXdZcS3Fu4mwRQC9+oeVarVhInPPR/1
Y1bGdyTO0jtBwgQC4zrYnxhD77wIZ3F/+OS3Wv24GumK16mq+jDg+QDTTJsq
zJqtrz/umKp/TMiO6MKdpT7qERkBY78Ois/ymvxKEo8+PQiEQ4bD5GeU2uZp
/Psf+qkkqCFDrVai/XBOn1BjjbbdX2sWtdIbat0FcTqcykqTfTLTTqAXcf3b
+12qbe5cgA//giAB/0OSfOxUFw+ueNT2RyRU3A359swfp4qV7KtLcoB2+mxv
GA3x0q1Ygmft/n3TBjx3UD0jEvugabb906hKdd+8euhoM3qFiZKUozNYt8Wq
3bpi6goqiA8WsXo7YNmRzpj33DxJPvtyaTY7lHhMSlR0uHtLuFcsyxUXYOls
19BfL91s0mreJoWuz5koiVuayJkl1i2NB6AGwSwMUPJL56LEMhHOSjCUalp9
sT7lLjhJsmMTQTCdSDZl/JcjJ+ufFj2A9/yBNKbssIbJ5bqy87Rhgjw0wEvT
bivxNCZnhPxWtnDcz/hw8vpj7fOjHISVHaojnvKWZR/SHzbrxtHa1RSYUpyw
Ej0okX2fx+HDuJ30/X9CI09bE6Z9DowwRb+Oe6rm0NyIAwgy7p5MlsF8jHkN
+rYnksIGxZN/7pnE/scxey9vJjGujiVrFGPHOkbAoKHZPFGf8oqdms3KqzgD
wFhv5Gy9mV/jLqnM+gtnD4oscvhnjJyAcnMLhlr70ir/Qag2qaEXAu7hfpSn
utw+8CDjb6hHw3PZbg3iCH/wqLKlXmlDXk7aIeQ42kkWmtgz0XYrxC4ctWNG
/hvt/gwiuJGH+q/PBFb0yoRYJc5WJeuFNL/gW5jgruSFN+hyGbd90eblsEs9
AVRJCZ2nv/C/ZLatTv6m7NVdahDol6v9CpEHamL8tzE56SJkFKCHxxXix9J/
NfFbnykys0CmnGtVc4+jkk9IQOC2oq9/Te/9pjErH6yGaFPgygY9tvwO2gIk
zUU3BJezzSVFD7pM6eeHCunD+cEUltVZvdEPt0IYBV1Y2wReKvEY812k7jSo
SXQVd45Uz7868luPrCSuvNlaBqJhoc1y+/1yyLWCQhBfMQbPa7YmsEW3P1Td
AryqBWdk3SXvuaHIugh6DwG0nU+nQKWzx2dbM1BpOHvN8VwL1M8NCYmyDpTg
dlftNdUV6VfiKCFTgYy/O2rSW6Mh7vHzHZ1NKKnaVAa+rCy7b666RFMcKHPP
dxwHo0BIxLIObWDZDZ8F4mOg+LXyprRs7E0iEvyTEH7/tcl1ULinkRY2sQfr
fITuM2QN15qh80NCjGHEkFFE63Om0cuLIgrrymDYkNdhQyb0lS2fQBwPrKEW
vm8/+LRODg+VRRu7qShkANApn8bSxOtbfcj5AokuvvsP6SAckQI7Sqgi6Yfy
gGhmCr7aWj9qo8LObUpaffJgfRPnY1Sr44CNEl2yaqTiPepkcw0sFbnf94ZQ
lyOXR0hynxW8C84DRppVaZFsVavMV8/Y0/jgtdv0lrSC/fv1Ov9GgJCBxyFY
I23gmA1zRgsVMrQN2IrjF+0YFe4kRTx2bIOeB0iw/Me1+aonCxX4vlyjwun8
pNYrq7TaGuhorL89MSbk8TEhBTDecA/M1sG2q66YjfilOOwvyEUQec9JtEme
Nf/58hmCobalXs3qX6xDgQnPDksfaa/LaPkZXl+i+ZPiSqb3r4iiG3LP1Lir
V8Q4oQx6Wg3V35QFakoB310qVUOCzwZ/6dNSbSGGVvhZKH4oQa0vf6IviZbM
xVZikXSDPDdOBroWqITENGsEeSTfJpXnAUpEUKLf2nUOpcnHSZekuJSWkP0F
YWQ5y9IcZ7We66L7/VCHGewXHpe0OVf+2eORIk0WlGNApW+Iey6vpX2ZBprH
MZCWNTiXVZPDWIK3TmwDTzm2WrMx9NrbMrmqzQjE+nugPkq4kTb4bIbefYsg
lY40+oOdhuC40swO+05+lGeHyJQdlm5V6wJwYqQT0Rgo48st4vWwsdR4JPnN
Ff7OaQ6Jh6lO9KSpI5cNhyBXUpR4QkFtdBku9eaY0Kte6pErcUMDGg82LYnv
k8AHARdQ84+LYtAo1W8pZIQ9YKuB+N41NrfZk5OYrzHiD/+BN3Oq+WsmQ4aU
OF5Yzid7k+4O+D0n9RorB4E5NIFlRC1mFvZCE/dT+C1ZBXoL26ZiyS1JBKgB
/9Khai4UEjLNVAndHGPCvi3MTmrr4W3wCX9gB2T5HczYQhAe63fFAdRym+6u
4N70wxR7sepoItJP7Jr99Vh/EARlHdNOAI68QXW57QaYd7ZjpylMiewNcdiZ
cSLiwDaoiS+TlI9HzH43q3MqTY97ph2aWvVRk+EApQWPgilnMeKCK4nw31G/
8iptd9nPTF2vlcwNRalLJnQhE1puTFTH9wVm/AUBOyivrK/odMevsTzbqDig
e4WcfUdlbgfR0lWSZiKIYEdGQ2quofOBJAyQXJ2hG+lizrylyPST0Oh/h928
OaFC8XwY/jjoZ4yze7h1XXDScH1qI40BxmB9eUQ6dIyrnzlNKS6CGMvaYqjb
eWGceqzwmgDjii0V3fEuZjmg924K41x5jj4WXWeXeO+VKxcm/rboXg3w2Qd7
bF8k0Pqfc9beq2vZWAJ8PHS+6a01jjbSx8Xqkpd9hUW3qMCbNuiFPaOCJzn1
JZ8wYEnV8he2iYJ9NbHPx1uXgjQmq+jR3N3qgGsQq8/56+L26AhdSLBKucBn
rfRSWPc2TU+zHEsNPALh23QUo+SGTrjC3pJvXMixbMawVsq18O9sRu4o5Zjd
ppsszqtLIJgmJ48vFh9cp17CnPZO+55Jw1A4baVWl+HX/GlMlalJ5VkdKKEi
WN6MhIGxrXO0iGQWp0mITceao1+JVZ8nPvGSMRjp8LfwqW3ibjb7ZFFjSN2e
oJ1XprQ2j6kch6E6NV1ldXDzFZhr3+i/EAdWhi1yT4hyv3vAeyjigbVPRYLM
U7JNEx+03Biqk1g6KNCeFq+3jOqfsDhjXnrPNnu0KGX3West9VvqTpAgLJJq
H3aGcDYFafVZ57TXC53+5bZW7UtxxJEj0h48WARI8wLNap7GMjtNpMwKXO8i
qduCv+5H/uHF+/R0b4FYv5edDcex7Z+QWGdNQuIElm9syx+bHgTqGsXKdSzI
cQLOu4B/jZg8Hi0vZ7nR80TXrviJAuGXn45830BodLNuSZ9Hq1M900kQ8tVH
gB60/sucbwBjKV/TqEzdMes12x2vYIBBLjndWmHIBAhw3DF9S2Ity5T7T79j
0PwdUpLPrTLDlAc4eNd/U0Yp0L08sT/j6SUeR6ytwqLS9erl5Jz6f7kG53/i
KkN9bh0zg44o44ySSYTGlZ154aODxIFi09rAQ2ZGsfw7hCS25AgfKmAdul35
vVbVgPs8fTlQkfww8IdC5dZ5h6RbYouizuOCO7TayNKiD8wDoePD5cveHefg
ukBI8puKNJtL9Z2gRGk6TyZY1m7CgOnlHpTGGRDQDXgG/DlJxXCg841gI7FA
7uDBW2IwzP49WLfp8QuXzaIb76hyiKisRVWiMsuyzoLu/3Ligpn7n+2Yk4yN
pFo1rkqkm6wQLpU8dRH1sg88NQ2ELOww6dTfWTVy8Mgzvdvj7jSsSSiosHd0
OwYqm5rEy4QR0Jja9k9XlT2vCESMW8gsZs+2xjCf2+wBiDn8kJLiGF8B/qd9
VfS6wiE5BJF9X4h6qORHZPO5FPntMm8tzFdLyibf7nRc8qFUh6+zrums4cd6
1EJu58DtSOxj5h+mWuTWJDtx/TXHi0n3aAbxaiNjxwO8NKia9WZTEDFxK1P2
CrJ+LrstI/r7WcXHGRYWsi8IbH/9iWdlLCNdyoB+/HqPgstpitWi7yD1ueAf
NPXU5nQZvwBtd94Jqe4NIA8aqsQhNhAr9sImBQKawv/ejjsSGoMxSwvNDSPc
1drvFVQJplICMl5JLEWJOHoRg3eBJ3I63AwSq1xE9OU3EaNKiXr5xAkkhZFv
CQUa43E3BU2T1nKDPq9f+1XLPCQ2ZdrlZHrZjGiIc9CCmpqlszCtyNF59DQO
DCp96VlfnDEnif6lZssZoROlIZM8v9y93PzXwcKuFkcVpKuRGry3u/KkiRtd
lWIdzM5Oc4MU/N08FbHOHrJDZFSAxATsq6YpvYrU2jd7cEBrCVYv9K7HsCI4
W8AzUCo8aj0ofPY7adFnT7Sgz5FtDhBWSa7HZhv/zfKqcu73/ixtcaAL9Hv7
EPIytL4gjhPSqk5o45M7odQSzx7tWIYgAuCUcZI8aoJkULWaWgdDygespL9Y
4O14lVcYBEbYsbOqh37W2owhprc1F/bliejP1O3FEv8htqqVVT5u39C9Jfug
YmL1vuSN3pBltlo1ZDmTP24DcObyVU1T1PshbvA583xF5hDZWzAj3Z4R5NOR
XnDLYsx+QsgT6381YlCPHk4gxlGVeBHGbWfe1zIlOpLru4n7gnkgpdRnFJ/G
XeQmEHnJdB41hnvOFddYolR/Kc2uzSwc4dfReTuOWhA44HbdZPwXotgukpfu
4HLwKEHE1xb/SOvkVZQ/cgiVKuI4u6zhDvzHwJjfnVmRl+P1xoPPdlCojk3v
zDDiyduq4oqtKnYjgKWHlqlEz7yYTv2thYuD+rlxmhwBZbrIihZbahedMYac
s5R88rYKHyHMztPN9yPdvHT2D2ofHDxB0XLKCOlT95Os2ZwBG/ehcmc3x1jm
K3etgL9jCBpv7CL741TYBYSTeDpQ3qt2YAV0cpoXP3gRrb89fr38kkzqhC+Y
rdRokEAbTCHF6ZXPGHf3JWUP5ak6NoGjDLkuA6kya6L4nmU/UH2SrYyKdw+K
R9RtFwNQQUIn46DGAUmMAv57VDg/G5iLB48YS7Om+I4XUH0P4AJ4gjIFuO4S
XeYKkQLRCD14tnND1CPa2yTOsgUAt6pC1PHRa36HyyFPr8qFnJ6qimMEWYOE
SaUXRnPkf2LC25QyN5tm7LvM3bHcp4bSRQword6rKo4ZjcrCTanHycMeaZ9V
tmkgrOi4dfF2zD33lCPceT8ANYc00nmt/wJttZRxq1G6/ExO8Z8Z6diEdcwD
rij1z/XmePRqnjiY74cGbIV7A7oscDUJwMgRyyei32HTwJI+quDpTv5TO1sk
YPasSyn2W/Di+K+U+5c/s1J9PjGe84WK9XCI9WCiwgLkyFHIjb6dhpvktmDL
pckhk8EG6ijz9PY59mK0LoUgHA3pQgV5kN61tkrEwu1YHIANHzFU76hsK799
JJgnV6lRg1aFFfJSgygyygaj0DncvOQtw+0kIs2PrscJ3FsT39bJ66+1ErSk
JE/jmMKA/Fvq0z2KxW1yiSWeI/73VfaTvsiW3OFYJR6TN3gJ5VdZNHhWNPF/
iICuQhDEnlN62aXtv82H1girYSAX/qESOUX6YHevRidOc98IWPmNDFnC0SDC
NsdGNCGvfaDnwL0sWw7ATp3RrCMmYhbOv/s0g7uFlyOWZC+TVgkrviG6aLIm
xGnanXx2P6QwjP+SsteSbiunaMNNL8I6Jdoq1Z8fxvwCbi2zpxPIoClmx+Ni
wqC6e+SAo5qQ8L4CWytFhYLkFB2CRlEUOhGjZcLU+PH/Er0i1Wn1ybh8Lte9
DhzSmMcfaWJV/w2OhrZOZ0q+EsyYa7NGQaZNwDEySNawVgTaREYIF52yP4nw
poPvMME3xV+ITfvO73oba8UpJkZR/jTS5vw9zMKQYc3hsBec3n/9/L8hmeAk
My/p5C44N+Qt24q4kdEcEt7l83+dOMYUL6YswsTEukqVMw8upDfiuGxCi35K
iZtRSFNkig52L2upuBZcPaE/JQ5SispmdpW2C/VDuBlZVe6bJSq3fLLRXUvc
9aiy1T4zTbQsGL/nNOVON9MYAo7Bvp+0jRE6NfsACThBv7b/q78zm2iHwSwi
XRJeDgfqtW45mi9c1mZSWsU7igEfCNZzl7UZOondGy4edB3N7A/AbeWZzrsZ
Z7Ns7NeoEzGjxzDeSCFtmDQf3oAve1zPMnRykDA7s93vOt+00Gi6EbWEHK1w
/iTEOjt0JdtOKwmWWo/bufV59FoIXZQ9Wg7xNVCR11JTV9x3seg3j76BqEoO
w5oXHDMJusGpj2IsSxFfJHDlh6NYXqucVZi+MIgQuHePm4kr9/mMngoY4DTR
7XsXmPih6peGkA4K741D8UuaB5T/zunuKhC7clXN2oZYROLdTTCMv5y2J6ZR
phHk1xSeLTokBSYlJ7wYyPbgz9hZ/aRZZZzRfrmFfUkQcEKnXppxRc2v3eGj
op+ZwTRSUXMx8fIXDZc/TeUX5FM4EHTGbqaCO85VghkXAjj0p5pS7LzDLNei
esXWUH3JuWDQC7K0bev1Ps6vX9txlkBOeH+z1os7xtLRPsKtrkPDnRti6GTQ
1ZOKtGMb9hKm69/6xDSOAMD3U58zI9Zfc4cof5ekE/BdFNxqVWf6r2hoPHW9
JRthvuqknwNL/cnGCRrTUBr3z6vhliiq9APRRnCMTcYzKx4ebtFKAvQKdBxU
/aW17jqnSIlURsaAvPz/ZBhTxRKLbBPqTHZFVKBxL9jQZcusoq/LMZLTHztF
qL59itmFxjG5GFL2ajOGAVwPT2sAeC3Tl9EAMo76VVUr36Xo4l6g5rYeN6kV
A1G/OEJHBNLeAS4bAojyxXIPvCXcdmNOELrrYHqk0kw1HOKw7IW+P/EQwAKO
EhzGhrQ0M3EBI+HgsVJfJ/C3eJYtGn/2pWvMfOYhXS77MSUS8+A2gedq7PPS
1xVbC3wJW6Xs6uybdnq1lrnvRd89CM7vLqSYZKAKIDSIYKn17gQdQIZtBhxI
VM6OleQ1hsNgkYUoTgfMjfBNbNZJ3aEiaR7abtaUs6x9c2xeByq0t422hyum
9i0LxyKAiFvo3aoXxBIvvQT2bwD/Rdo7SxZzykh6WB2K/+4MKpith5ykfU4m
V3GzmxLNQRZHukjIYs0m/8mwnGmK6LCfr2FXeP+MtpVeatadAr4rU6wBClQu
xRmWzjbmDV9NGjbcwz8I7/SfNBlDiKCilzB8/D4xn9hv7SwJ86QpreKU2UYU
oyzyL9XTuykrGPA+OTmdxsfh3bIoqxzasykKuuNi/UjiVBKhODscXrQU3A+Q
gnTKUMrVc/nQTd+XK/zG/kQ+hmqOidJbxqofvdASiyEgbNdXGrwxeo371hfL
VXpShRlZEPAEg9AFDRCrJQFRTstzl+mqZB2AAw2orPTkNqX8XMkmbO51v4xC
zS8vQBWPEEvFUNFroqMNUPWezT74QYGysC+he/geHEXpGaBh3bUA+Lt8zuG1
CcCnazDbnfN4YIRviDge/dVbwPZbmvcplirWSxRB2Zga/EzySnnmphWIAXJT
TUmRco2+Xt+QEHe3/+ac3yCf6RTctFapzPALRCHpIsDZq5rO7gHTzvdrNs//
weP4cVPENFinjKguquRI7+s8h2kB1qPBhrA4nfwAID67CJ6XsAWMHTA+dEBS
kM+gFZOUiBAqDLKTVZQXner8edMD39+7cyvISqQuhprRsE9Q7jEGTQkhJrP+
8OTPMgPbXyro1QbzT9qjOa/+PplZPGFwe2dtAvo/k7Pvg0RJ0v1pnBibTJ/5
zUUXalBEHWtZD+4hd7nYuYLM2qpvu4f5FmBe4O7DuWaJhA+dkM6Cl7p9NY9C
0zeB0VQdCmnz7bFH62uU4b3lQzT3g+p/iqshhcpauqEd/p/P/nDme9fS2JxA
2Cr6rmRF1siKUbp3FNtOFrcaFSqWCFnJrZZtxAYtC5ESK+ZiRYlEID5ZD5H4
8XcBfZCL00HuO/vVNk7bF5oPlUaLjA3WuGxcbwZrrUZaeC290p6/8yc1DouU
JkPev5no6b63RKPG6BFiaFHq97s4amscMTAbu4d5jIOB+hZEkyDepgoXSkHB
9q14J8f0ngeZiIiPJvGodKAh82vjH+xuWBtjM3w/oujqwxSDV6xqyblXnza6
xJaQGQ9NpCP9jV0FhQ2XqgDmY/20aIF/YajVndUX8RX/Rho8+zDZpBAgSELx
98nbc44J401dXqkWSs7oGt66+gP9T3ljOIZsccToge0pEo6CgXapHfucI6Pb
SdJq86F76L8blOwQr0BEdJBQoIrNzuCaltxKHogP/bXidn0wXOr/tmBYQDEH
DwV21QYE6OBCfcC0sO7rlutQrfZSXAK9EimQFSNmc4Ffufd5usGxljwyqHSM
QMWC64TT6cfhKZQStlm0TyuXKXuti/gOBv+2Lcc//KQRKEbKAyRuQ2VZXIpq
MVeDKOFVs1UcLyoaOKlfVNf+7G6v7cYXKFnQAQAnpcRx2XqnyJp/Wsceo6bG
tRua9UvLqTeFc4fKktY7UaNqtGTTJpdCf795/6KW+ZsWAZHyKamn2nqXnyYx
sEkKsn6pMDDVBRs8w0AxeWl8LMegZzB7xrGhu6LMmOLSw8HoBsCxZ8oQehRg
wWfEjeNya6uZPrR8v2ND8i0GXBhQeJ67R0o/x/KHyQXPSuFXFpFnVUYFJCWl
iUtRbj0EG/xcZFm5ZHtTrgo9OC+pLcCYwoAbyWe9aP2fUsTEKgtt0uMmxIDP
K5CeYpciBp/e/a+JhbTK7ezjfWU5wRZhAVSJvqogN/jbmBvMaBZjmJCOu9xn
x50FFO/WZuguPoP6XVGr2FrR7mA6nKZLh4RvVN1miAB8BhY04/PlJyiIvMhg
qpDhz8pPC3NGGcwvTIi6C0QsXbZP1sFSsxaH7vmiOiv6+hIrD/83Z2ICLW/5
Yc5BECzzvonVYUFxzaZQQ50jmtTi4sFyALppbiqFVr+cuXbZppZ4rAAKOwQp
yPoXdNfpy4wsUks6klPjibALlCeCGGbYhRRS+t6jLCKqmhwX6P30CmVMVI/z
aXhXp5hYXV9FbO726Fy2bG9L0dvx965YxPsWFDc80Lm6IeaMAtP+jxldmLAW
FmNa7rlM1HxvfVSC8KH9QaetqxHzJsWWuYYdCh8H7QGsxNnGKfQrgrTmWZw5
16qs8pJhhOCKhS5KRd6O9AKowL+i/F14dUWg3UWwC+/r4ag0J91zrz5vMAHk
WH0TUx7ZcqRdYiRqXaA4fL/5MK/HZOlj2KNmoOOxArUAhc0AdPSH8HlcIoZZ
5yXGu/QPVpdMA16V8EX4YMzWSRcKm6Bli7zNqfHdljoApyr6ukPholQ8Ol4E
h3V3RUJgvDQaLI+4In30N6yAfYiuFYyaG+weHjDAJztsgRsI/y0tkmSXNS5T
LA54ubjvzt6IRoGRoq0kTXAjeMzXQIdDf9MYj1qIqbFxGTREuqWg8VZEITYW
O1kpixMvTqRAY2AD+X6i3Y/osz8jun8IpYrolgjeHufKh3H8eYvO+out9Wbf
6egNM18/3sxv+qc7p+7I9WbaDGKbiBWjUkAq25/iB8kmHT83w5Z9ihOV6Jxp
3qhKpH0sj0oRHWTJmPcK/CY0WzVbNUq9Xip2MGJ/+L9O+/dM5IFbHRqMlQHV
g1K42YVIImvgMasX8/4n3HWn5y61Zw6ojp5kkEcu5WPEQS2cxJgxVHUPeIy9
mbzS9Cy2V9cfWHoNVY4+yX6BSGqSb8O+9RSy2FXnPcp5Z0oBMuca1TKEqz+V
WAV0RE9dt8OjFvwDqdF97p6pYv1ldk9tgBQVggfaROq/7qyAhNsEMhG3zzB7
0BTWj5adeAh/U+kggI3+xC4yhJq1kZHr0n6BN00evgIVrcub1Oki8/nGwJ7l
RG5c7lchgdvu1Se9MA93gQNFG7tpsltqvtQLPKUWl5Zqxg6frGrUO4Y+nM7J
IFJHYvYOPDbv3j+dZqKzxOYv4FMQU6MuL62DtalEcjkc4+Ake+Ba4HDnPgp1
+/niFgJrAXMT2E8epJSM0HMnInJXHn/xhL1YaREDVDxp6fNxcxtaVtIy0Zid
P6ws1WBo5T2RAtFWgMH9xW8wCIyBADxT/2N10l043oGWiUWFpXDY6QUOMqJR
t+dBqjDoUFiAOaQxqeLlAqeFXeVmJJPn6g+ETGUvIUEBcHnTnAIkSL0juGWt
J/fDWaonBrRp1YpvBYE96d6jVhtScpaOXcOEknVn/HS/1nwwybzXnnq6a8Vj
X5M5Gpd+r185aam39KAZSI2KlWXjtc6tnrTiEyx9APJkzJtzDWQtJcsEvJae
ecPeUlxUKWmj3jnBrVHzoFIydbLWAuMMzo+B6IZOXkYT5hmwAOqdmWZNWeiX
ZI2GPB2sWB8ZfXn33ZuW0uBQOgM8mCHhRMaiG9R0hx5qvLBLsAyqsGWcayDE
pyYUOheHvzedit99lz4llMljzQPxJSJl9wWoCwfkKiRPpEky5tmccSOHdP9u
mD2c04DplPUfknKU7UyW07LiL/7zxi45jl9CXehEpTeejIowDir0fGWqNSyc
o9Zkd/W07EjK8NLSIX0Xe7Sin0CISkwdakLi+W/D+vQc2GkNxifJD4MszZZ3
5sATFG2KN/wobDtzDm2qydymU4JhakadO/iJ4021ZvqYcbrNel5B9UEQyzHm
eUmfF9NtO6uEX95gab9YLNvPuvP8Zs2xrSlWaY5C/uyK5PChM6Ni9rb5Dxu2
2NDrVS5vcNxBtJ8lbgVOs3QB4TZlh7gZ16VwNp5ii5XcFOChilZsnazR4X97
GGXe5+M4o1B+XMmUX4uB6NAZ4WZXxjDNw8PxnvjLwaf5jkl0YyygBpu4soXq
oOnRtb88poYcvrPOdaxGia1+GP2/VyFRiHkfQuNiQlJmUFjAI1MDprl50mEb
57j4D8pY7Wlz3Q3JiMThxeL/yzHC7nnVqLpT4d8NDfnA0z0rTCWoMQMCK22G
rYpx1K5H/dMmum33U6UocjZ5OYDYXRHx2JRP3AiqhV9pOx+4vx0Ra9JyDuZI
hEovsI+sAoATHJqze5iYXXDu0ari/Zq5b5E5pdx4HBQqaY4C9lu7eQUWAvE6
P7t+9tNLCcvL4g5ddTxOzCWzLxuO7Heu4uqHm4iDScvl6PVgXcmh4Oerhdhs
AxDAETHWIgiQTjyK44Z4xNV+AhwmNoDh62/csFpezjDRk8YqgIeLMhxuNFrp
ZcF+E9cwCJcS0YtnELGuUP2oAwom4dE+DKsHr5rtScOsRm1KXqFUtBWifEdO
2euXThRW2VRoHgqYZ7oWieHWimSnMkG6oatJlDUYQ8kl58067IZuOXMQKbot
7jCO9VzjYU3MGhmxEjJxphjOsaywwhfI0yycZ7JLSR0ZWULUzwXy+BAZO/Re
jCD3cjJrXmjahQip0rGsSSHA12Jxg+fWm0EG1zS+5Kp/BuUN6bqPIcoJkmjK
m3L+PvoD06/vXRKGR4ZEFjng0vwU0/YEIg9/KVezyxS/zBZCruPfoGmO5u+t
J7QSWpudiKy52JkrtiULlAG3A/sGeTM5KehwfgNMsQVT3CtlM9PlLVe5vN7S
yAi4+YnQwgcOMayVwLS0izgjj1WtAUwAmUgwNNsfpdoM4E97Uvt6IDft3m6R
vvr2Dg/kTAo6nYpAY6+ZFq/St+pEN5P/TwmUnGqTSAgNnnfAIsE1sy7j9dcf
6BDWsD2yYsLuxE8ERLXFqfWzgZrnOyuunEdtX26zX6/FTmqlr7IsyMqY2niL
5Qq5JDlP7XHGxc1pAoW2A/LDNhCleh2hJRUpGR04U349Tn/VJ8i31U+EmsLO
pQBi+NEgE/iWuS+/lo5Xjbd//wmYKQz73O5pZtjtnPjS3TB8GXasSe/8D7mO
nrhRaQ71sxrfZsSnJcBQluMVUAQzrJpkPuR6y+MclJEpYyAU7TIDO4i9k66Z
awPLNbanPxdLvmyK7XzqvIvYtO+d/ClWzHFwTZg1QxOmupCx7ZGgXVPvFA8w
+x4R13TWJpYDSIAzzDijzzhlwd26dqXZAYoQqLE4LpeKCE8BmCDZcNhAADkz
yuGDhuJL/9+zezkSzgk0tJulI7Z5SM7679ZYS00DLW4H05CkMEPbSpYe/eQX
3y9qOs0ZGDt8AjLozf4hFS4uyyZayWS1ce1/3HhVugZXG0u4rHOSp+gYywR8
KlO9o1QrwnlD9+ItDks/PSJvMmFntVGrz6gJqYeAFJOUgg59dnBTd8KoVRAM
qkeeZEMfteil2ELiVF8MbpD/aL0oetOjgN8x+V6jM7/o+3Qq8y64ac6eZd8Y
kHiXhJ/AgE8Z9xd7J6Ry6/RX6gbKGYaNS7rTexqRHQdPXvF+2nxpsBZhG7iA
cl2Dgbex/B9POrI38Qk5iManK34Lqz4tqD3lfDokU3q+29tDRrOhW9PHS/UR
IcboJqqB+E2u0QtSt6trT9ty4K6tS+D6xaXwgBmd+oKxULk6j8Qc8e8ZCj/W
aqFUBJoUi30sqqIkgVhJT1URry1hzw3FLq25jpLSoKkoCAiiWX2neP7ywB+R
a8rxtK1fJW3U04Q000TS8qxYLMEemdmujnbKyDHe+y0OA3w5ziaO3ROgVi4f
be7NnpZgxfsjljwN1BViwkTZdzURv2TkbgNXp25h8wa49IBBNdiVCAASYMp6
rHwyb3U338ks1RfRDuGUT6QBNABthPrNg9p/+M6UbjpWqxhnjwRgWR6pXFaE
pSB8Pd4YuOQA4lP1vaqmUrDyCp/4kMda+zhFnXth5XhtNkNYgOLTPMUgyqaz
JvwIbi6ZtsCNZ5BnPl6VWaHaoe1oNrxEBJF7RlZRsoTxDvFtJBd97ROdSpRJ
JP9QVwFmnay+YwoSpC+3a/PKQ8DouzL5fx3ioOOHgjiRE0qL6gh5EYpmhyVC
5gX/NvjXtS8TblrBnM1QoylOmPBi07xOxfjvLtPDx8mxrkDGTOga1p7k1PxA
TEeZ44DQERyjbY9DaowtR1WUNWPo8t3uq2qyFnWtuEZxwoE2FviwZ6Ei8D/R
EWEOty5V7lvR4xyRU7V8eDwChTBB1U04gxMRQhTQTZ1x7VLd4vcMNaKZLHL8
Bm6DDlLb+6xzTG3i9fGmoLnWQpXF/CcrNZlqozpMVy17KxnDYTg5rHrhbnAC
SNREDt2Jib5QU3ZczId4bj2mh4+OCl1m/MtidT+Dxj/JkZvst+3QpQucSmmX
wCZ1PAmEkPPPSwtkV+5F6TC4xPX4QyF9yU9mg266T72iWAT9wDtqnLZrQ43r
FJC4H2vW4kYljePfIqGkX4HZrPocWFOoNtZZE8CeLHdxqqsT7L/GcIsmwK3A
tFmFjo7gFYds7uAi8p/IWQxJbu5LPthQ6JR7AOSAu44Sdgy7hJDcIYySN0hS
9ZuxfBiGuiEz2P9dM9fuJG3bVmTL3bqGoYEa7DeXxQQxFE/YIglT4kPxdDN1
CZIrKA3V/KsqBHRBMf57YLx6em8zPsssKYNMeLWLy0nuLp/7r/+Ke7cS3Afh
mEEtBHE+C+tTc7TjiTxwoDJz0uODdpq29MCf5Owj8hAIngicQuaEx5ud9XcF
6eRm87ysRPVSGm4Gl0/9bo+mKrW6gJC4Kp8oXt9z4vpRSwXwoQ4PbsYPnH/9
7HjtGp0GJjbRqwH2SQacBDyKNym87stTVJMNOQKf9Xy06Bj/JRndMVmaVDu1
8nTURrOF8tD8ycDH2JcIW2Jzm7bx2PiSuHsbgVYc2Wdfpefph8J6AZ6VaOWG
YU4S4ZQrM1b0NgbIQiKa4f82uYfuIJBQW3K7HStBUoG+Irdrr0coBwbGSAfe
p7k8AD0z8vwOxU0Ix+YX31oKKfRhN77q1Tmi2UhvG6fvvuskIKgOLRYx3fI0
2JzR6yPu8oE2kEvBKHKV2aGt1yyL5NsbIIU6XOHlOqSlyaSzg+yAG+xf4VyB
3WxCMhlnIulKK/gcxlaaTBhdCTqQKrbjvkCA1BnQhpEqQDSaZqsVyzEyC5kJ
djO+tEUjU5xXY2yXu0fp2FcLh8UHSOxGhrrcWgJJXEjyaqUvcDxw3w1TlkB6
atlc/ahRGiue3i4EvuB26zLDaJ/LRv0qD4imgjkqfKeavEC0SiqJdoZPIe5d
0wxE5FDS9jgwYF7oCN5Nmz7sUzkmPYr5bkzHFiVACuHbBkAHF4OqpJZx8h4K
85VU80REZHQ1rR+bU66sDH9CUDG7bfeZGytpQmhF9grRroLP2fT5qClK8Sp4
k81xFPAHvab1COi70bsOdhOudJBDXvHKRFDNkeDV6APKtWqZHatjUAl4IegK
Z0KdowuaPwO/r8PQscwCbCWruW6stBwyq3ibCSC8zh5tDFD2bFCRZQ1+Xcpe
4RXwKvHYk3Wdy3ae9ciOEOacYEXEeCpbFzpWlJ+iE5MYctOZmLZn+3umx26I
Q15+QO3wOOhCg96acCYiui9rn11aHPGBGGBOscfYu/G8PtBL8xLjWL3XfBFz
lwO2GeKigNt8W2ju5KKS8v1kzeV4BxShSEdb4BbQjWIEcLJqTZik4P1w09lU
ExdDhQ0ZOaxao0RgHA+pqYTN4XmWsNHBg7ctN5wkfOmne32z5DNinhoxPT7Q
R9g7MuH8P6MkicasTVbAh+yv/Ujp7vaObkMmnXSWju7TQyqwjJuV64q1sdZy
PbcrvpbC3bhx7BctiOSIP+Y7G43KEYM90gVhz4XNHNP6VXAnziLHrJRtkeCq
+bxiEFK8EGHvdEoBFAioVNKBPRfgQrAOKM+VdFAVcuTg+NkrS4uUUCjK9a2M
BZvvNlycqg74ZAAGjWBr1V7eD3Hanxj4BnFDh+2UiWRtPvuKRVBDf8qF3R7j
DX+kcx9E7gk8WeVcalaV+VSqx+mEVVFM7oEi7V9etD6m6rHIODWq1RclpYEl
4vZWCkwIn9ppa5AfBWsiw6f9jfRB5EP54T41r2WEkYlbflAYRTQSSFNgFvRV
yM/1Tgy2bJSxGUl163pnT1lCebjZrx9EMy088iLQUypFg40SpScjuvhOuFyL
15/XjF7pWLyNfw8FZhb5IQ0k/5M7u8SKdOTT9RqWteIAcvAe7eU3Hqnofckl
ki/BOX2Y3kHkdZpni/rB/vKwKBUcFipxVMIzgFH77MJfBzjEZ/LrXWBuNs/6
1SNyR/W+s/JGFy3KDJwkGF9vuJ7tHMClCzlqshrFeWu71UZhb9IUHMLE6jya
vl//NAnQnLZRVkNlftZrYoDzSfG2x68uMSjTXtQFm4SGexhIrF8yvUDMlGl1
scTh5heQmdAs3ZOQ8TdhR2aZvhidW0JW4W4rm2tse/Akm4T6ItWvxSE76wn0
Q+q+LDG2fJBz/yVLMLfvcr330btElw16wQR/i7bi/Ymm+0alPVTyNavfOCp9
E/sMpfwxvJ0MuycVkwIxdyaDwJSEp6GlFhJ3bHixnxh2bjngHnwttL1l8KNM
QzULrqlKkVx5imti+LPaMxFQRL3enqOxj3/jn3bguTGLixlMiHEOSq2tyGRb
rwIV9xLy6/5PU2K6MX6dmNyiIrNCa0lK2vb+wQme/g8URoxiiuKRKLQOmdET
e5gDwLRdGQkN5s0GII5j5Vu+FO1SChlUJs12a7Mjk+FtdAreYDLp1LRXvndA
odsIeAqjwaUGRpcv6yWqijA4r6JzT5X/Avl5iTShG9cce7x7U4S7DbI22IWt
Yv5g1RBHljnfO02YTaEgsXqu9rSMvDtCeDqyANzCz8de+AEf6brFgjsEoDyo
rPSQffdiMyXcB/L54LU/3EB320khNuNfOo1aIl2pPjbnRFgoMCEJIVENKpF8
b2c0a0IZPtdKGBBX399eay396aRMHDpCsX4qI5DA4Tubl6V9ngl7MHqDoL3C
+O/9tS/nJvNs93gQxWKLFFzfPgUBv1cShC5b7JN+XvFnMKc1p4O3mtb/FogA
wr1M0QdXG71w2MV2cLju0l5SlB+f392qGTk7ksGuo1uk7VwVL2Uv2HfMaOi+
BTCYObhEpRrqEMbupDd6d3emR4PU/766+OSIW6gLMRGm5wZZnqXHiPI8oSr5
BqaKocmUbw/n6Rd7IsGfbKKj6Z6+O+27X/dA4EjxadYw6XrF2kYog5e1att4
0uKhpvSJIksnTbnkAA37+uSmCG5/LX34AyLJjhYO6jgbZuxqxJ2OROlIEaas
unxwh8g/gQGZ74C3XfYFPnG7gzm0YQ28Sq3DyFP8hL+JtiZjQU6s4WfLrHFw
6HkwOvgb9UH2Stc5sbDmfDGXfzFk6RCa62mzK5ysj2fwvD4uJotDlsmh6BHB
4NXII4w3/KZuHykQ2SupF4Qze+8p1MOf1LCFCVA8sDIErQLsahc37vMi9lyD
f9qPEW5r1y7uU/wCBVBeQA15ZPYjVFT0SOU/Y1HUAA2CG68c16GHj+orNgHC
Q2OCk4mCCQbGDsnpTvgk67p26O0KmbT18GI8BhlKly9TMmL38uaLuaPrrFqY
mY57wOoP18poOXFGZ4E+fkyVY/H6bx6/xi3Td4YiVgequ/pb8H3dyAfN0Kaw
IwTb4lKUUa4nqKW9uCpeG2iHaPuF5MAEaXS2GXap6P/bet7oF0YgdC0ew/k1
pAKZEFAAjaLA9Ov4hIiMvX/ydxohFex5EKnIQVLvRM1LH4/abkD6r6pWSt+k
n1iKyasUysfdBo82uISpzsSq8YTgpKiId4j2V7LiK6WB+tx+iE1GOyS6penz
T4LHHb2pPCfDpdX9YWFJzz8TQe/Tuh/gIsZy3qlvvxeF4DUQCGP0YyYI6NNh
bEIA8z177KnCQDnqXdNdoVLw/XZRGrFi81PI0mMoJ9RTZ5GPaW2vJymH8C/G
Hu5GE7mDZaocViW6y7HIDhH1qL6tq/SJg6ZFDpXwAt60/Cwhy6zKtfCm55JC
OawMVpyEylW7kPnsltp/fk3Vhw4Xk4ym2tFuIjsoR0r5CquOUC714baxj+BZ
+AZ59/98mjiWb+e6xwhVODq8tkPTWgTleGk4TUVyChA8z93L30/dhbdlF36Y
tZNVwWMToKMta2j0M9/2tqdl598TCf5wqRHzcvnTJ6rNgIIXx2vceWAsQnaT
N900ESI2bcVgdbTrCjEVJK6O8+6sax+c9pKOVaRceVNDknItO3byhYbZOSGi
/kqx6ig4dEce9NEdgk6SKW2C3+66RwEq1Qj9n8nnEZG1u7XlbSN2QxASGNL0
MTUNrf81i/gKWPbR+ABfzbVSa3FyCGih2YAMf4R5cSJ9GN4JKZMa1lZLfozq
TJI7zW1gYxBbF4mbN8t8NoV2wOx4Dii0WA3cVLNjS9V9G74nnc3AmPuKvbpa
rrNPWx3dlsuuIrbadxP+QKYRm71ICeK8RWGdJ/8stXQg3OmS0uWEicb2wIXS
69bpUC3BL3HHNGLYhrXWIIgXLRpfcPy/NQKkp6KFR/2Nvod4DeCA2ZjBCLBS
r1sRvRzHiUVgKuAj7ggcr1lelnkVJAAuB03ClIFMInC4g3bfREvJ+XlhbJRg
5ag4e/9In8YnWuiiBDnvajf4YMVWB7R+mf4N6C1XaOb1BTMDY+Och2vPJ+3K
f9D7uNC4Fp1FGotOTBeiXPYHvMl0ikig9Gy5oU4cU9lH/ME4J+CD+DnboTPH
kSpWBcX8U43xVxnSWcBdYvamQDuVsfHWf2G/8ttQvk7gyqr1dh1iUu8jL4eP
lVKN7RzCib8uEcD8xX2vNVMfiDNH4Q63jrwJLrFBN/DbB8f/fcFboKgiUVMX
e7Xh6tkgh22kJ66QzCr24IXXCz2f9qruDLJuVSUb74nM0m48g11jpt6YmevW
7a9XIVAwTJ06Xtbfvl5/c9d4ObDvuo96scetYAg4B2CLBSkLR4K6xn7UjapE
UwySkw6YP7467WMDMErtP8DuVGjmrkwmnzwkObvyvq41EgeSdJbv0X7DJBFh
IZjl3wDkN78Srb2dgSinlRdqw+wKuEWSgvFdPwLt0TtLYn5fpFmyXPkc0W8b
4Aae4A4teVlJmPHsbDkuOJgsIsUl2VHiZRnIUV9fVzqn+lTqH+uzX4Qd4ksl
flDXLKdWjOq51tnukwD76b6Tuoj4t1iIRJdK1ftS6JA5pYPXeAglEE+K+2Ax
H0jAbEcS6W13l7YDB6cEjPk1wCjUx0UXyGG8+rbxEuMRI1diRtkJz+5VZcgw
TH1vLbdGjxO0wanLYgOYLzodJf1do52HdfgheWhQJX9Evt1Kxkj8xqOeSezs
/i3tWXfLJLi9hC2fptLdHnRjnRKUaAd0no7CmkJTlWbP4kNRmBCYqkNN3EOI
RRX6hlHZUR7TobqHI+Nu388EtuG368CXcyc7gXRzFNVnd/eiuM4+oxgdjY3l
koSTfrs6sn3q/KLmB+f9PZBcC8dg+QvAWyx4jE41cNua+K4AiJflcagzF5G8
QMJJV+kZf8rcXOxnKlgrGEhP8iVB7rl6Kf3A614inO6/SMo00CVJKbsl6SBs
8i1fktCDplt4JGFFdVecCAsyOQMh+hkggQx2hDJWtZ3C6GNmzF+7wAHfIzNU
mt75f8bCUyJ0SKelXEu9y/PJVH1BbtCG4WQxYyG9GgmXQOcn6bCjqCylyDXA
0Kn2ZMJA49NgWbOopCMp0dj3Sc2HfuqRV29J+p96vqsbwTJXpswNc2NciWw6
9j+omKO/yZuddcW0CLBJePKO2wCNhJn4gkI9fJD4kG4h7ztBEtM1CJNvDHLB
FwWa4YQ8HWERyPSzeRVu1hsGiPVn/2Z7ZBxz0L3ShNNeeAmBawed8s73l+Xb
7T7nLcqqEjL09Xrsj4G5f7nmzWO/9isOA1EFaq2lyPs6hDkOJP88cvKMUfiv
39ONOijvCqC7a/P847eXjlERiWfxY8Wlu74MqjopYJBi9EeJHCaBkzDD5mSs
hv744hjWb8gcdd8PwyZkxq7uV8b/K/djixwadRfOJeUpA0Q/c+nGYlG85+vG
I+BLM2sYq/rVp/z8UZd87j6lIoTTQ+4LzTd9emWGuaDv5pjx01axhndqte6N
RTtByYKb00qS962qc6tnGUMzW8IHaZfuELYNxrYHS2/uDi+dBjhiRujSI4Gt
QPnEAp0TEWq7nSoqOPQLcI1yxFhOJ5twr2EYebZenacH1/oWl7+LnkAMS5/f
2TCay07lAIOSh9v8fwvi+FGMIhs9B7geUKjiU8pQW4I90mCCp2wfFMm4yfzB
UnFg2xerq7KBqc8DE3wFZ5rQ35s5R5kXQ1rjLD4RP1oDmLwIF8Jftc++mJ9Z
Lw+KoyduJfEUU7eXMaDNqJ8cPKbJ3UcxZsuUuxAgovVFrXCrkDyHeRu90ZAM
HEwvPzbE/FRSIGfD5A5xoyVuMaJF8c/CcxIhElI8wuJwvD36cuZqwGrnkk68
8/BYz0WAKjW2OB3BpKG0lxTmutoRi6HOr2UfnkLUINSogQarMJ+/LPV1zCRm
eMPUE2rSoRD0z4XKiccOd8O0Un2fAnvLZ4rbbaPiemQrhJ3Bs5UBa9mbTdKE
0hHtiGLwYf2ZZNNy0KwcOmQX7URJmZF79d+5wwoKT2P74zspi4rJ7Itroxf6
SU0wLL12h7Qdhz/reGN8kCrfULkt4JLMXxrGWpEh02+CEU4j3aDMtzFgcEEN
uyLm+jfaEJXbzYOy1NWLIWSctDr2HAlqMjMJnBSxyS3wUxEebije+PziRO2r
VebfJoVbXfUDvLTGk0i/GJnsGwJFue2by4N+2hdGDqnouYqdK31q86+10vcA
KH4U0zeKAlMB0gCiAvlRQuphuZwl3KGKBnpUo06iQ7EVOqg2LZle+Lq7c51D
/gvS/VuzqAngzywDNSoj+1XSFDKe8T7iFfafMCGbaIPV9KmxBKuK2FSdhPUy
k2uaZiFINfHsgYnYgTfVhvKYlLnpJ6YJfjQqJyP08sFzlAzVWA1vBhfwrbHs
IhOzJBGOTw+5zOh9Pu1DpxbE4X2FQKu6X7RdlUguZbuUYW06fBYe0yNylqg0
0dhVbtssbPwzSh1e3IuBXlFCWBztcbPbohCa6fZ2TmGNALExhcs8hhCNBkBS
YJ0VGu4k6R7CoOSixDH1Nfw/qFTBbWLAFk4+UWfbFQ5oazi0wuY3/0aWciZy
iHoHWygLSgWBcYAYskQtjgXyMO9YB762CqCDp+/MMDh6bv+5rZzd+xti9147
aA+HcW8Eb9jR0VKYklOOmxPZueNUbkwyMzSnIWX4ASBuDGRhduhIChuUCCIC
zT6vIBATx2IC30CFEThbREp/aZGGUhk3/amUFG4PySLI5EaqSvqOZ+mXCKmh
cgmQuulbTMO0rC5PVrtvMi20hnqRKqWTh5xrexhCynr3av6dVXDiIyHBPVCj
W9zvGK/r41h6/FEJHoG2QfgrF3vbTrRbK14nvd5j+zkrV95Q8ED0O4bkVhZN
gZk+gRo+UdOnwksYlRhBfAtheQqGLqUyY8rIXqBxiIQNKl+TSaseUa2Jo62n
Ccc2cnCd210xWLkwuKWO3x5cAM18rkWlQK6xjsC/ImzM1SEVgyUUxKiMX6pu
NaYDLwZ9TZyP8j9lYRsE8Mfh9xURlkoJrYzomLHCK77fkxaInkI+60yUVMBR
4XZjkQh6SwRGo7F+9ngISn7ZS8S1kX+2gIrCSqPiPn2lKvWgWQrcIKsDXYmr
KhQ3bGR7OOAsZhytlikWfZYrQui3SOrI1uCyEu9fuu9osiVSELSvso3mWmcd
T69EMOFeJ8jMvQCLAVdAzoTLrXiQLPqqVaC77lIcrcpkbPzCJTuRYiFrYvMs
nFsd2LJYX6yGkCfyu/m73xL8Ax5niyp+BlvUt3Pl3mW9AcXuqKdFegZbap//
nFjzxZJHZWlJBi4rTMFijFsPKpAQ+qzR5cd4n73jUkDZaO0rNYvVvxATxa5C
PGxmnDfRufJ25RjnB1iqm0dOz4yQR2rWu6JR+u0wRWHTuPgsbMDKRbHo60h/
1VNV6hqsCL8xoh6VtF1oxFJtced5I5AtphSc94OHQrGyAjudQWESxaHcb3fT
nn3V7k4msNOWk8nhbXAM+4IVilezFO+WTB4YpHaduzekIn2fWsY4t3+iqTTF
onTV4emPI1e1wIcUI9Ny6ydOMdVIOSsAZJQx3LXC7CGyeOqsmVUVQc/rsCL6
3ow2+AYoWKrKQWE4rQDtfjklgN6F3qSaWFJ/W5RFbSquHk8s/MSPiJA3dseA
ADojU3mlc4hzgWa8L9v+MyNDAORug9tfXlKvuI1vbySQwDN3gz90kHfF2nnz
k9OpAhvpd5dbrr+i5AaLeeYliHKEykE7uWJ6Y6hinKxrR7D19fzgNcbDW55b
7r9Exbq/CQ62z3tLDILRSMfBrKPWARj9BPg97HGviHJPD8vV0BQZ7bCA17rp
27RhfLgcRjxSxVe2L/noAYeO9OLI2iygMNL+zz+hQbz00aTtiiwfICecB4nz
4+tG6whUVugSlKBB99U+lB4yPCo9Zjmc0sGNs1jhIz4r8Nxb8pfPLL/H2xDW
0IzOZBy+EJRPD/k77Ri73kRoubxgUyVzsxdLiAMvDm/+Gdg71Kj7PKz6SXfS
x/Pacs7PsQP+h9mJYsKFaQoXqYF6zRyh9noleo/9DtoReNcvX8P8luFu8JA5
WrsR84nDCZpgd//wT6+5VVi/UM6X9IUNLEqKIW5oc3OI1e2yEYxDIII/IMxV
qUbPTBwSjLEIau8Jn9w+2L0Yb0sEevFQmBMzEaxif6ucsJq1g7lUnLMhx9lE
WcsFsYt+UZF2uGgtccRn9G4kWfJG6Lt8vWl/wVG/5f1tq9wV3HaUu4iVyj5S
Xj3ZpKTlCfWfHgXEAjwgXdbyuM+9aXlT9/bIflj125AreGCa+YZyp0hJg3S7
ptlt/0wjShhRAKYJHd5XU1a6REYMu786SV4vqOVAk13NW6n5dYqyjxiTHWdG
l4ijiVeRc3PRrtYCIzRE8VzlndKkpws3XWlZsYDuawkT+mSJqF8FSOgR5tMH
2uRRyH3k4BfZ6YRvle3hDyn7+i1QEOSTC8IqggurW0NVyGJH+m8YFU9X5Ssu
rQUSmzMUv+/MLJSd1Gc8vGREejxhm+heSqHknS1xqcwaszY0stIZfC1UkwXh
vQbr4atAFxOb5pLt9ZVR0JKAJK0jWJJZlmKSIoGeOOli7uwNTAHGNqhVSaaP
JHYpwG/mWNjH0zuITSSdCFQa4t7uPNd+Ml88G7I5CNTbypwG1NAjvo4ukYXE
Auu4ib7bQXSf24xz8CKom1A2DE8YuTt8rnRuayN1L9AotpjIE18WvLTuXVba
si3Dq+jYQiQeAU7CMwOAZf7kXmEYCFK8/Dp/gUAYMUze/V6tLt8gcsfoMGq8
MCzaOg7kp5bu7XzecyboOZTu0unmN7YBaUG7F6BvQDxSSxznGEMMdFadSXUW
Y+LfUyxElD9uLvpEF/lgqqBIjZwr4tRzd8EWrxSGcjBkH27j/EcwL6SZVlfK
89Dirnk3+y+AD2dNTurqyYkEp9oPXdft0WJJIVBfwO9Tr+1Oxe4Zqkn/qCmy
j1B+YVeuxrJLyEdbBMwUnPpl5rkLGVodLHOymYU9hRHlnDxW/TPUThn8rV5B
mBCMHld7FBB0EXfV26JhvNqJXLCL0dFqTU6ISg1oo5cHc8zngEr+R9hU3cIg
hWbgJxQMG+hlcolI8TPZN3CfdB7LCgyHYhxyLVINPFfApTDEPZv0G0rLtMyH
+N7CTqOGJZLEbA/uDz1MwNwONmASoC3/nR+iKDlDfi9uqqCcwD/DOjE3jZsU
IcJah9IjcJdKB2tibduiTqlhKqwZjK1tW4VlBJOG2s5s3BQkVM93W/Jdxgx4
b25kOk5fqnzcK/ePyX0VY8+ljnYvSCr/N3J5a0xIG772NyqI8KmdvXBbN5he
BcW912MBa81/lZlm2Gl2RpL0fTTs4tslrS0dNuUQ+vd16VEDr2Z0b+0xU1sH
gmgfjAcFkjl+W4S6VNiQpRyNKC4Qqiw5tgs46df+hoFi7pejKfh99xyL6ubP
a2VXpm93ZuHKc971ulyswKKV7KFYxmQvHs9zx8BDZEfQsOwWJRRFOdx2nMN2
wN1kCxKVZAtMCJjQHLQpblOxpsUK9bA0xA43zeZj9IZxdDmaCD3ypXQarAZ4
v37ZiQZWE16gKQb5t3bIkZAnC28pgk4cSM6/BcI9NO4EEOIOsiEp5D4teogM
n5CafGld7VMy+DuqZc3rQNQUcTam1BDgLdjEz78lY0Q1/sIaqbOn9OSo9ohz
6laTmrsp3+9/3N+Pi9/ARSXYxj7mKC9wizbjiHy0EjoJfjEFyCrwQd0v9cLO
eMFNwASj3hLmyR6Jf1OMhVmgtM1iv9Gal5wHXtO+VoinoU9r3U4MqGAyJ6LA
QXove+VZHngiShy02V/hLlh7rFFyNfnbNrVvYTGtiS2wicKGwsWgv5wbFfAR
u80y7n4PTwYTuaU0z4l/jzOia9F+IwVNdHl9AOvtU8arq2IRo95mKtnD7OwV
q1sADQuQAl2SnsdhULPkw1y3yz/Ehv9GBx8uSwQ1ZMW8Ph99GoCg+GT30p4J
NGExA1rX/z5vFtl1iE2f3JoN4j8z295u33LgazZUr2zObod3+eu3ymYXQxa2
D7n70BtWtc6Qm3Uc6WYn2M5XtHF1WC2C/LGOG0vuUWn3XUtcfMeQ03syogfS
lZ8YJaNZEtRUKV084rjAANdZbxhgSSJB6/rn8NJqqgp5JmA8QyAK+CdaBDvr
rlwAaGrJcVrNuwR3mcHOT64HsqGY7nAX51nzXHV/sCvwhS3X6hH0ahuxKDMz
l33PfSoNvd44BijhcAzYS+qFIrJIyDOcO2QjtV4dYUpFr6pA5uk5ybzaWNRV
PPc8bUe9c/T7PyBnhEjJDwvfvdS9DupsacAVYs53QwXP+Blo9neWHIA5PXb1
mxOU8IlsI9kmdacZ6JrIvoqra+x6V8DLf+D4uoF6Lf/8WHExOMMfZkSX7Idb
S1gkAXwtjXQMLJI/4GQVee2/SnPg8poKZ3isiAcK814BCqvE72MVFv/D7u3P
KFNx2khcEELwGUD1n22lHIrDk6G/iVhZQ/GOxrz0ni6CzgSXTpS/BiiMGVf4
pOa6wQBuHJajcWZ8rYgZ0NKNPzo92UpQ7SDbI3FX+hH/o6QukFLTnNGxlVpT
Y9pJIS0DMpgeDPZdt4LWluae2lovGc1o/sFtncseVEi+DSY3O07FPCkFiTup
N6Ow8WFKyh3t4JsXngpuNjpIViIKUlFbXjmziHOP3Q4ihDKAJHknmD/iEfNT
jBa5rDgATR4Qho/L+sz8WYir5apu01LFU5eqwEmTq0XdNi4dzR6MbavZFaWM
mQ3uuoY5bWrcbjm5FR42ic49PK7LByGRFkmvpdIOcGQr3XZBbODNA3jLB4gE
xW2N7FvoJbxk3v2wo+pbuli7uBQgjpuLPfnu1s4Ac26oOPK7L+zAtbm7G0O9
3FCmozVY1d7LyEyhcIRHUVY4hTYg8iOHEe9lAFPTC3wD36nePc64WXoWvuPq
QuGZ4WbdILP5JIzcKMWHMgKgBTyms20hgjHtut/4y1mZXD/SQjJzB2AlQp7x
kfSX222I4CYwqaO11YWZvyvy9/aVPISpDcu3HE3pGZjRdo1yHQgg14b99+YL
9J3qqyg6g/Oc+lIPmcJqo14exU97eB0cr7pTdTZxkKRpuRuIALzwKhhJJWUb
my3g3vDvTF8F0saS7jiguNYzZGfjJrahNfg6ZRyuPzZRuSnjJ995KXN4ZNjc
f9Fq+EsFChpjXnSqxiM8tlK4m+4b66v5DiMhgD0Q8lSA7+Bs2LDYpHtYkN2Z
MOrpCXKD44LCtov2VovWaG0fAGB5aQ8L6mN4Bfu95Wi7hNSVQWb7b7yANhWS
5zH7ii0foxCZ9Oi3oWnRKn/r9IsWfhsSmX06cyjA7Q00Wn8pcph67BnEqXtY
YsBLubT6QYni1a2jolMIC6ZNgx5iLWW53KU1vWVIZ82WBM9TA0fs/18GcH6w
pUqQRPvxA7ACRyZqTWp3pvXxNqK4r2DiiqoaOcdRR8pjq/SLjfGbGD/ktzcW
iapuwg2Rrni0yBZw0Beeu3eOtKpMEbZibpQviYHZjCC7VnrzoAW9HU87ulyZ
cXJQGBtoLUP4ANA3oxg10LLX869fx4nt9HoeMCCgYPFSWT45G2LQXP2YO/iX
K7XIbUCdKq5gkvryw3RCXKf9EEAlk/9VDWHSXLGHG5aL20knFlVu7/k71qBb
qQPTPjprkHsS72888GXiN39WQIJQwI2Kwj9ro7G/mnrK/noKRal87tqbwvR3
5xDZvsI4Ty7/ZpJPDoI4hv4XlyPRwjYrJ5kPESU+WpZIAPsxXYIqSNLaZkg9
PkBb3UpJjuk6Cs75o4mnYOYguLNxE4KvHB/dwSaEln/AW5QAeX7kU1zzUnOP
87Hmi/zDtlKlCILq8DzJjWuGGkTODXAfY4tkDNWkRXvCPWuk8UI8qQcoGfw4
cbHR20fR+XKjrPZCqUfAkff83bbhI33KC5n12oaYoAXznfGXvnFwYIOXxNrv
MdvqTNgLDP2cYSplYYLYeA5eVJ9HBlr5/Fw00ulK8rM3M5GJr/F83GIAy8ME
H3SQk1qZuzw7ZW8dP1sH8a0P77uTwLm5GZ8WEvACzcx1g0/QLbTo90w3Pea/
fjkqvIDKj7dxMzm9UwDQLvdqw2471THowJfPZ2vfMB+r6fih01cO/EkJKFNZ
YuEInzz5Y0FbsYBDi7LdTGV8FSEHgXw67+uJjR1Wrgsiq2nVhH1MdKRw38ER
a09AcYMU+dp+YAlDzaI33mxcWvXI/BgwXw4lf85g7v0d+iN6xK8Bv9Wr4f1J
54p5z8SvJNrG9/dZRSlMHUC3svAWn5YQ3HqNtaEv5lKFhoj9gQ5dmyJ5Bqvc
jsLBcg1bBMro3WjbtlPT9IHHhwMCoJ0ffPYRu0oUYts2lLwlSMUZylalAtCB
dyu4ej9/x6ZYFaJp/Z75pB3A46G0aF8etG45nj0N86KvpRSSpBs2omveORX+
dqOZkHXY9KznTyPgQzx1BdxvVO0XNtzoCDVD5wgMpDSIZ32UBpG82QQfpzVj
8i2sIoobvzpTTnwR3DLSofaUfCTD1DgrP71rnzxFL+0rnYbVdBD4z/o8Izms
jccRVm6enW0h2n2Z6IjgcxnTszWCX7HpoynarPNrBGCQRtY4Wfj+gp8MA8D8
INygN29+4pmAdNkUtRFo23KtGJj7OpuRrZZp4eOazRfGnWJcXOse5VguFx+6
nilN4988QF7r7igO6naCHHC7fXizurjNnJHAURo16kS6/aeBzUPNrCO5J0ey
JC1LxW1TpkShhs/uRJk5FAPacH3kikIw4s32z4irkV7SVbIVpsLKY/k8SQ2F
cQ2OnhIcLxiSELQ2OAiLi0XAk4QBum5QL6b+8UvFuwwgppqz3jGUBi7Q4eJI
qr6Ii4QfP2xJStwyVWBlhAjjcPpHHVEBJAR4DNyz46XB3vAAbBZcdcButIOw
d4p49jGhDW14N5UV9U/UXo4rMdisI/9P8LB++B3/TzcMBT0gMyUZNPmgUUZL
rwXr9NEt13CtNe0nnlZ06pEd6cc4ZyZuzKjHcs0Q+SuhVfMpqSfGaWkz0OFe
ZtGxElMCmiFS8owoG4XkI6+gFSZ3tFpY6gaBTariSuOrYGuiI8YJrwYZdGIE
/G/i73fpyLt9D8p2yhwshvtPtisIJrHGx+R+mV5j5lcSFbC7q989YREylQeW
M4BFxo1MYVnMRPbbWR6CJzNeXm1Axv+SrPJIPm3rFeqLImZO0RiQTvgUGY5l
SqRQC6SYdDSWa1CL5irCsuyYjvS8OHU/48nxz+iMOyI0vv54sVQPPb0JAB3l
Od8AeBQxgp74Af1ORDIOq8DdCmBMcGuA6sutgom1LBhI4AxOUjNaiLPQBsYN
ugoiR0jGllWlb2IhhpsFJJzRcLJE+We6l6YOZidmigCrIDj/MDTA/53H3lUH
u2aF3T2FxuFiIOCtv7mFFIGGhJDXoEJasaKlFJsVBP93Oszw7w+IUJ9XVAyR
lLwJnV6nAqhkhqFsoWBrXIcS4+1+yVYVYwpk5q5e9CefqFn3jJa/D/Kz3bb7
/8D79llKmnpu/jW9Ltt18YghR1NR0YFQjcMgqXnEwrAkGk1Vuhq+0hDVvXwy
WEADYtTIkvBp6PPCWEluqCs5HC0pETTWKqaAfSAkrecgqMbP9cyfLwOoEvlN
erHuwY/yy5PolqllDvlqjV3ge410AzcukV63z85ITsk/CD9aLKisymQUQwjJ
nE250mYgwnXsXbWtw0c7WriQait7mkKVRLXndwE9pvbYmDuRtjgmoj0eU0A1
+bhK8dH8HtqioDJOrJOWDUkRoqwiUsfCtFVPrcP4+A8mRSeTRPVSKvjYlZEs
HyFy2h9LzltnWgaDbTP1F6ssLMfBKoWXN4Mx9yD+/YRajKwFeKryr8VVjI8r
o9reqmzFrAOy0DPxN+cv5thugWoSMnfseP6z5pqZOQ8zo+7VlcWKFNlac+7a
xYZg2F/7TMvvbsn0DfbLz0VOpME+f36yTGSUY+HMyP9hH/h9v1WHsVzKGR1x
s2ji5ABGBet6eGeVeQ1RL7p8btkwvJmILrCZAdnG9xcxKHJ2MV/0qh+rOEei
FHdl0lD9ZLl5YyycPSTIkhb3EUOwID8SzfEgDgeNICisqTZOH+XwosS4Mu/p
NrKYVs2TyF2TvENLAPmNkJiaq6x76XfkARZihWrsfNTmjIcHekIZ8kL8t+/7
jFVYXgni3UdZC4nG4SdQRLKQmVq/rAckdgX+YsHfs9XDj+t33j10X6d3NOkS
yjW0EdrxalBROkwCg+6Siq3YAbrpuz3wAGaj9eFcLR5NmTCy3sPUGO3pM2Nq
/x3kH05lK6dESkuYPJ33NlXX+/3VJsPg931XRTgRIiJNPRT3KKYfCWtSuLmw
ZeBVyY6RnNYCg1bmgMERvU/Y0teJzD8I4kolT+6D+B+j2xQSbvw9VVG6Cxfs
F0EorIs+q7vjDCYFP0+T6H5eYLRzj/bGcUHJoFAjZVPKcI4RvsjPxCF7qaW6
aaRQqSm4PZNbEymY0+eXgPtWl5bKdIu5JyXVcKYKHhuc7wHpgH03FAUB/UEJ
ppBg/FTQplCqQouARMsHH902yGEsv3ar6bAvVDXKlhnIIK8cPpglG2VJZeI4
q8VMneapgHrNf430lUwWiNcLXCfDNS1L6pQGLmCEQsC4tnNHww69LYSejSeH
eD4yJUntpgIxjuaCRjy4eRRWFJBTEVqn9XVJ9GhmQA7tFkd2BVW6LiKU6+Lf
yjOVhj5DNZ09jdvkEl/3QHHkIDDQipL1plm5TBSMZtalol6MAu49HhcbPZNg
PfwfJkCqGTcTNupFcN8KFZHTh6kEz6d7Jfi60uOpwGmpVhkgpDey45Cb3kPw
oX9MQU1YuZhrC9NjdpvdPb/ObE7tCYbyysA+xzIKHdVY7TlCi3XK5oIwMldw
HV7ypTs75ZjJfC0XXNM6v9iilXMd6VuN+vinTk6t4NCqwxjj6fxDPiEeX9nK
9pI6tnBPTQyA37rNZBFmECXpUm/0Lz8ba9p7ZdA/71op91QpQaQ4Bl04r6jQ
vYp1TcBgMKcgNqeZY57JJHaEYpRhXoEtNsFgP11HsJZpvDbI/VxtThJaeADU
2ypg/wBqIWyE/WtirAG2MmD7slP8XwaBn9/G/9rP/po77rrxZ5aKmJ5Wz54b
bS3i1lJRBTMoytGuchEcig5k3IfTMBXj3IOQEqNT3mn18M2v+B2ybHk50Lh+
xeAQHwDVPu28NOenTakB9yvcohWcATW47LO6+rudfmjPaQDuhVBnwc4EL/vV
m5KSh7//LZssi4Ck5csi1Xx0ohL+Hhzt8ArPGZ7hJY9ElaIbqGoQ8/uJjE9b
J+9/3sHO+wcfT7CoZmIYUbhYTSCcCzTRJ2cJItN351JvWmb+f+sgBI2b8QLX
ApljeIEuVY6QwEvtj5IlLgX20CMMq5+0xI6bh3uAloxxDdAUa09LJKosgAuY
N6ikXOr+omZMf7W0CmvVok9GUP59bFUOF8XM0cfn8oPcy5hzdJFvLhQYUmD3
1eopuL53odFtXyBWP78VFZQCyva1Tnh31dG4QgH2tLxfwAx2wuA6HkoNhYyg
5I6cR7YpXttAOgfNqgZ2tyBAlFMkn1r29FM53oscWYQaD+4DO/xtmi14ww1V
aHSOe25mzrje5wGEAV+H8lOy1XMESQegYb1exvGOHFW+UWBgF/AjXlYyf7pf
xZLtlq24hxRLx/jB20CpCrxhN3kNV2h2Y+xqVN2Iezlkrhc7KjHdZO09F2P2
DKO45LnWadYXQO2OomX/4FiQ1RrqMFSLdPc69GbOxCNsR9pnt2su/TpGVZrX
4iFB8Iveuj5iUbyv61OiJa3V592HsAAO2ZGOLMbV/Wpps/CjiDpre/VxPpn9
ddJ3p3169UoRc2Bo9Uj4w9Qq2eEZcV/1nT6fWyIioeXcW2VMexpABZrz6JvU
Jm3PeH02n64/AHp0NndtPZIUZTGTjTv8artIDxXbr2YDIEyDk21i4BRD/bjb
wZcdra8bxSRY41E3fSY9O8FJeAcHIqQEK0CxUIlIxUqKLtD4wOj7RA5Z+Inq
VeYjL+12R9cE6F6tp+ocCUJnXuLVZC520SUCJHcCJlsok9ZxmNpgj57jQVkp
dHOmeCrK3V8ec8hNZS7TUzF6Y1VnKmQLGPbcPn3FjujhuAcyZ7RW4lcIYFVH
nxLealW7aeIixKpOrQf12vw3GTjHqwSJis5iZHmhuia/WXLH7g3wwV/mHUdr
9URadzh+KcxIVFO4SY4zy5SMIn7gOdFYjW7DP8+Kasx5Ojsz401/g7gQIxYH
hElGj3R+ukjBn3sYx4Sit5BfE7Rvrm74yOqW3Pf4pvN//Y9gVyE71kJ241zY
Mq5mfong9azuszJoFawc0LLn1aV+9/Xzovkeck6BBdiSIDdcPlH4yVc1YMRW
XABHe0kt4IJGAVg8J0iiSMgK4kmmLsEu/Qd8ibd6Bvx3n/Z+hy9sgXD1vEHX
WFOdt4O7suq+8dBQUZLnXAlUv/gmpHGuKZwUHQL+Y7uqbbzON9//fHJGLWaU
ioXYCv0GLQ0MICklXsSY/4xHI/3QalzllTOjhcIAhq9BzzwMpwWycfyVpIjN
Mc2CdTElJTM9Bts9lwbEkdBLfkwed7T0eJhYUzWw4L05iImpuSMLsiRyq5AN
bROe6lxxmz2Hel//nMsiJTBAskKUnTxayGmHO3PYWGOWwEqtmGKkr1BKoJBn
pa0oI0jqMPdUzWChSKEyoAnZSOebAWP3qbYjtnZ4iO3/j5usChelrftI4E55
HfZQ5skg4THtZokHso9rE8d3D6unWNZn76tRirrx0+bAmL97j8xpBBlOAfmk
03dtT0dswkAn+l4QNUe7lmXBaHHhFtG4Tz8njYaOZaHyhLbirLAGnVVhrBoP
98SzW+XLk6JElwidv3/3Vb09xZUCiqlFx7qUih5B7d8pLsYu5gB/Vp1rhOrd
8xKulLAN6vboHCeBX/tuOFH6Ke9butD+vibmOUQ4PAP2EPOfoVhEgeY4a1m1
VjrH1vubv2X+i/jXGfvUx3vtGpMWG1oHcf8uy8B8rJyccTh6VhcYxxafEDL/
KLjBfZv8R+3VlYwvjpkR+QO+ceYq+b3BfccQwqAQJ9mh224qx76y3vPa+N0T
Q1n6HwxBTzYM9bRINXg+II36jk5DNivCoMHs/aVSZSPjfdWcM381LLIpfbhy
VYAR9RS5l/ZpDL+jlkHqxAor4xpy/9Oo0blh/8MOF6a1zNDzQ3rdgSA59h2G
eVqJCa179rIzwJasw2/hYCc4ytNB2GrcHGfHzhWxaLsECoLJ6N6QaOQcG764
+yDJ6aDHadWc23SSCNWCwIOgrbrlAN/X1Jazy1rLPkA6VAUCwojAneZBO1st
DrgV2f7NgVzR6BERnvqMQYDkR+NonslaEw9UCzQ72xgeCnqSxV1QXThAiUDV
TamHyla90Mdo1HzrTfOXPG8GTtECIr7tJIrpY/aRrnptxlZBv1PyAMVktQPn
UkDZHs9DIz3kItIc0VCkCCD6IQ38S0u1VO7qBC0ABMe5IiloL+EFc6in0Gni
DrGGOL2e3vLnHkTIhWLzcAhZ++Q+29NdFguTW9oqr3/oKG2/5rxAAmsDZGcz
xwJKYJIzZpFaBduNxVQsJ1Dq2xKowD/5/MpBU4b3xsreyRHxQ7FuNiAyGL4P
J/WyICaPfjALe05XeE4/CI1K4ReGbd4J1rswcPk5rbvAxI+BINJEfXXzn8eW
ICYAbI/7UzzMOlQ7HS5zk1fPwfDq30iEaCKQ2mMMe9jonT/6mqomLDrKXTZM
8mdaNjgG7w9odeKzejuGuUuIE+4L6evL4p2S1kJ7CXeDR3hXD1sXpBofgkMt
ZBHJxE12EoSz/LJlnIFZOgdckdfm6nrN+Mi1qQ6uB8mADgjbNvZIV7NPakKR
EPBdiUftHsDmCeemZevtmZDj9+YQDqH9BpNTTPYAYqJKC8K+y86gbF+4A0a7
bA+pkIgK1j88G93ufLB4/bssMKA6b890NaVgZaiOnwPMG2QLg5grzG5W5sr1
qoYTWZN+Vmfi2A/edkIweVf/j0GFmhWwyr1pCTYbVYmitiSNRpALLOKMXlcC
HNA+V8vXxeCARACeFvky22wi0eReLJAMXc4OLJb0N7yGH48h6tHip7kR2NvF
Gfu/8fkrLxtJyyTr9MYfHAie8XYM5PVsCAUqiRef+LacTagpTnHskfMtvI89
Z1o0rSUZKe7InBH0jZ9tMH96HHGDsQ+JjdFo4/9K9JGlDiwxOrxh+iOdm37j
FCsiIjmyz/WPw8oOIGs9DrjNp+YkI+/tcbyMmy0xz80K1E/XBsxBsGqpGST4
Dql7xh5mq4bUhi2y9iP9/cbvvMT3C4C/6MLdLnpiP2Q67K/RGaWnDGCRp2n7
U9bcrMmsYLtCPA/WtimSozQDl/zFIgWr/jpsVwKOlgRnw5hAgXAis59u+dm3
R6dOpRqMjIyCy1suY5OBUY/2Olq+JTkXqFDy3OcHHijEqIYbBm2rW9STn7kx
dK07fPozm13rv74d15XqjvmyYMtBHN90LTMRE7+PX3ZO68OVGPB0RKHNcMf8
f1CEmMxXp6tkAldPlKuAuCvULRZZZZIw7aZKSJPb19bTnjCX4x2Vt9/7TDS6
kQJiEZWMaHlf+AmR5gnyfc8IJlbdaHZDOtm2lHZ/i49xcIkLj3Brr2n5xyrm
VbUPCg3JpUFyHp6CHvMgiPdc08KcZoz+qHXqdXUhfHRr1NzMmrOQG5AaTvBc
f7dB6VPJZLizH+KBSIyXirVwvKivXTglZl2cinm7mgBFgbU3vuXlltvIbBp4
6jYCEffKUNnKqGbC6w9PVYWWveU3CsJGcSCvhWSdRPI8HhVKZGlmzcoH3EOX
RLL3F8SD5j7UEAu19PmvkXltpFcubrn3uIYhN/i9kZxgrExprSNByCVbCljf
GgVyNdfDktS41RWvkvmCYaMIITBZexVPlfql/Dgr6RWaeb39XxdP+JQEU/W0
0YydLNEiBfnnyReSTP312t2D6QX193IPhXAyQGE7NZqww+JteTXF6vIO3aLu
IURJU2dsI69O+e9eM9OfPD3YO6VgDkGszsKexrj/WRtZ2yts9YTIRekoXCsf
LaA1CSqot4ZV9woTxw6vAaFuUwZZgicdBq0nI5sWF4yWiEA4m7YsynRpcaH4
MDJ5FhODT//4MZ8IHhppnZrONLn3LMA6gKMSEkKR+fOnVZaznQnrv+GC8h2/
eNTdIOLtHuTg2s+i3mashKYFPsUM+WZ8DwQyqjkoRMD58rEyO3RTXTDN6oUX
DGEYo17cVlhq2ddoGqa/KiiV8ijKth8Yn1BNrOcnfw7iVLp2dRty2G2vehkf
9JMmtzT2FpCLH9Tg+JVj2lwNrsoCi0IOXLXKqTLCjhmNf6b1Fw3Ot1IqxcpJ
E3g+jGu2iQVgH7F3GQTgGAL4X/3mIZf6/KEL+Ncza+agkbgcb1VJBu2DZgBr
6l+dydWcivzhwOlUyu61zftK1kM2STsx1UsqO8T46virARMzhf08g8AC+L1I
VmVKAHLWChT6XgklkvcyKV+9/uz5aAWpqe23j0MDnS7XGS19yOIxeuXRTm5U
QMu7JnebAKtkHT6IzaILx/HGeATM8wBZJlRAjIGZE0hQv4ci0DFqVjvuDnMN
/CuWTSYYCFcCYTGfkY3QSoCs8CMf9hPO5TRIz5b8EI9HawNHqkh7g403cXz3
7d7n23QSVSz2QsdFsYDTG9IJDiubmswqjnPBPI9y5HUPAwOBoWyXo2D+eP16
eGuLQNFxDZrZzvItyIlpAfduNClNxNDcEAwGeJ9zYXvByKaQcXhxeJPaeS87
c3D4NqW4MB9MedMWlEI32LVia/yfMqOSwtWhw6srsS4khs6CDQtSyT7bZW3Y
iMmrIH99otZqoO5bNgBjg6bww+hUZEi/1c6XAR7iNoKs7ARgXqwBtn/W8F0k
0s8SDcufQ6Uuu/fPvyfPUPYD1wSrwh2fnmZB7TtGb69gYLzH+EYmqklfS81p
jniybn1xo5FkwTlwLyJQIfSYflvfWjyGlA1udEzYDYeXYO8Ox9Uoa3R95FmG
1h83FXDR0htnE81kEF//aYdr1BLykF/PMp26ENJShqlewTtsodXVFgMW03oY
b1j0o8743NUjL/Sl94owZQXnMpTGZE7YVMoW7KVxJkwGxuvhJT1D7cWD2XUU
JDtNKlMFb1vqRkJyqZBmD0SbbVFjmRIxrsJI4z8OTJpLn/sWyXLIjE665drp
7ATE7Kx+q7Ew8CUKhq3OO6W9wceYINt91/HLQWQ2Rrdl3YdAQ1m5/Mw42cMC
Jbp44fG9+R1VGt4rJOPjEcqFFFJLOzPjxTyXOd2I1KEcyiA5nOYCEjqHzJj+
q4SRu3O1AbIhCLDoTxG0XZIqGao6F/GJleM6CvesAmYLO6UwtM+xa3m2YAJb
SdEQhGf+DkWt5GdoPD8qJOqj30Ue8LPX+haYk63NZubXG0SfHJC5Bznvxj6i
AO80BWpGsBv/sZVkDzn/cR+4eBeYtNKwfFkAD5jNC5uyNSDF3LckCWBE0HAt
JQnBYOuGCVoOpk9YwzDioIggFAD4n+yEVXX3d4J8G9ZqizA/sR/emOlYCblw
PpFeuyGphiRD/IIk1oX9aLhnX2PNktBqBXURu/BmJvi6fwDngjys7EpeOmeg
pOHhT2lxLySUlnTHOu/g2atY6GmCUleXk0LEBc4TeTHeAn1e5j1QybdbX0IV
dWb4Z97ySXKek3xkVwV2NigVThB2RgITh6CLKz3CNxz4/ngeSvBICi8InFpU
pG339jgWXE035yz4P89jqhxKDN2eb13BhMppdi4BF3MhdXOMtHlOqaLHWdaz
VXe3FaDmt+h6e8qDmN+hShcUH/IOJdql0RV3zjRCXelFq8AMGohBL79gEVeA
D9XmVtzChQdCu1MSvktqt1IDifZUurqH47//2BmhWh3iBu9dTR3gkeUo6gxQ
Z7L3nLcuYOmp1QBDXsQ6T8iCEZ96NW0+B8UelhFcIgxZNyiFyMYxG7ON7uJM
xz1/1rRqS27ZCnk46yfkdByI9BPIlSRLSDVlqLJlkmcNrLJPHq/TKGBYWV2U
7Juu81zwRHp0J6feb7IahXYdEEgdSTxHqVx18qgOQCwxB62ZkznTFsnbM8D2
iFctsL2hKvWE+EjvKlZ7dVld/O+7f1FLOEscsdYHColSRsrJ4g3eiEr6M+Yi
AoWdFad/tHWugRb2C7XjvIJT+3bN7hbC6XFRwEC7KYB7uWTG0KV6DCzdnZXR
MGqKRqesGMPwsFbOKMQhrauGoVXy7EDo7gSiSP+QJoA+ZNia9aOpHKWrqvWk
42BCYDQ1jC7oPZZFWV5qpY2KrYwUV1RJU465T8xAI7ZO/zhdxtQBU/KN5THe
SStIcBdD7n5xVWjWzzoLKGHsnknd1/cNqUUizqvuVxeXDzhlyHVrpMRmx/E0
o+dupe38/NZlE2FBW/Ws+rAPHB+G38T6zRijNurAuaO3yEVJNJyN1aO0wV9l
/j4O9uMJSkWZjJcQ8an/lucs9GbWKfwWvP7e0uAJ0ZRZLlaFk5wHpd9kwBL5
p3zjtXroLRqACVlKNtdt/LnOmAQ7iXwPcTs9vL1pna9OEy2DzHNhOLhWeuqC
6RcuGCUreqCvTahk1/61zGw5h3Is0EYe0F07k4KvyP+nH3jiBwB8RUHhoFKm
vkqRBwrL1NfMFjpJhW/f7JzAmiFsXi09jnQy/S/w1mh39pdZI0dW2jRDKdGj
TSoicVQxH/U+URhJWqkhkw6FrEJvxWU/hypZhfZQHbPpbJ9lifOwz4gU6wXO
lSLorj248JqgemnwIUUp/cPFfVPlXCxnAzJHO0z1pGLaV/AgeN1OsxJ7d3EE
rX9VtPSb0jHjRdGqUKN9+KyFjZmj1lWvhp0kq7vox7Vrbn9ZE9YvpCuWzxBN
ISlKYOYYckg31b2+ICOnViYxIVEMlbngSnmzRc1S6P3hzJPqkdBPrvpMiYmD
cZ251+2krXqbSMzPKSNDgWiAJFNMaqnViKqhIAqfkm16An1PYm5J2PBKMaEh
CmUayBVxILOltVyfpbYPa6jvO2eQCs7WPnJZKI0BGV1aT/4BWj8f+lxaTTGo
uEILVrK5QTtSlyHqm05PKVJ45VddTEYuOGCBQo7ShdZN5vIJfTC4tGdNgmMr
BlfRrseVLRfDYvm7M7hJVn6I9MNAlld4iPXgBZ+2f/ch6tbyIndGzYq04WRt
Q76I2XNvvselEfYpJGX/AtpCIKw2Gqz+02qRKNbnQFCipdPvzYP+2VFxyeT/
OMLrdG6Xzsdj3gm8LeJy908jTmmIs6DMvlKlRPnEuvngxK1FkqKxGNRCuTdm
5POphvM1/LJrksJRjUFmhrzn9w9L2YyZkDKZmt0xZs75kqU3PQj/I7j0dDP+
qH2/7nfFPvMvKYoOIPm59yVyKILcrek18SXGwvauuVNspuQb+Zg2QH47xkid
/xcnxF9yowQpbVGM81eSsnmIj9ScKJac/86HS7AeMalSkRjhw+b1Zq3RqcTO
KmjSDs/zCPrbSfS1pe5C2Wi7GgolxxEfNgedbY6j2khmbV1CnygmteUObOtR
CK17kRpKhIUGIls+6+/WDJyt7WksQIdl/WNbQ3zwOv6XNuR/apGGsCF+xRW2
Dty3IFxPJFlavg0bfwWojKx1hxLbHHelTegapEC1mbMKDStyGxmRyEib1ads
xcPyRm+sraFr7d3Ny+xFSpAiBdJm4N/IT4tYLgK19nmzwscbduF8ub6Z4gu+
c//Z/aWvdIKAQK4JHfGfbUb0jsJtQbtd33xDRQS0lYq+odxMAqzhX/ImWjQ1
cqz02icxvnD/uVpev2AQtQsdh5rhhbsc3I7FoNee9L6PloXg2UegZ+6QjfNG
gyo3lT8sZg9Xt4mPDk4HIk/ofBXztBPR6Pq9aEhNZ039jCSLfm4UJ8nIUuxD
AOySMEx5zaJBuVbIolUanQtYnfCA8lMTvNQxYTTUDJVIrTF0+m2JQBod2kd2
cRTErxHTBmUGu2cHeNFBuEz3cLGA3i5+IIZPfS4a5v0iwCAuIZ0S+WP3D/Ae
fPZ0Eqgdgly0E9d2SuOvWpdeMlauYIvamCO3GQdVmvPEJmjyYrb2RSMvpxWA
JOGmU9CjW4DezHeORLPMaHyhFfhNL97ahHpqe7X8FOVpOAYqzw8yCzgGCT9f
9xhFpkDUQYRpqS/an51QmYmxPQ0bxq46BxfeIKWx5rqBKGu/10GYve17Hmv6
8/xTzI88CRpHjM/yQkp1sXOmBXo8yHtACejGPVV/DPS8AkyfQo3ZmuJXGTZm
9QO7EOnKbCLIcAUe28RPXVdmUu/LC9tVJZ8Vhf2y3yZsNOxlHmQB5zN4Peyy
8Z+o52ThrLZMsIQFwHNBUvVIPWlVz3/doBL1ETnus8F3Cnk6pz9FZCXPfL1M
fn7g+XCyisC9NyOoNKk/of5DtuNf2bqWqJ0dAlMkuAFiI002V94vGkvNRN9o
q3LVkjvyGGFx9kr+sIataB1vHzlc3pugF8J+vRNT7nSfOVPG6SADpJbb5iwi
0QKoqiypEVDE8HE+u9z05dUDUoq+ldAICdKAEU3Qb0Xv8PguR/HQPRFyhA3Z
J3mh2WQ351Wy7nwsHoV6JTBNL9+VqQiJ9FUMEdxxaMSYlEapoM69sc9qblSk
bAETy1NdpESSV9RFpuUWXwhUHaWqqChcdjpaqbwSJhBxf6u6qhBiPFmrYa+X
mNKYPOfPIu2KNgBVnfErEEBWbCP0T+ofHVDT7UgVcbtIOMvv5L3QjHrczaKQ
SaML3SW72dX/5SacIo1QGQQbejHgn2GqXCR6DhDoYR0MIJDQA+drzyL3QCiP
U2os08nOE8umJrcVot4MG1DkvjE6363lB2wFiCH2hi8natQGkOyuv/thfsYh
LkWDJaXHF9KtZOXbFL2prgCSdVIv3MKAm3XzaE9oAM3NZ6SRwgwBgG5oJru/
Y72LBKVjaD66YpBOF28QE/S6sG0JXuD8y/yewhEP8u6ucXnN4Gqoe8Il7IJA
X4tXlYUMVwJKDAA1MUdIwlVMem+jWEAV0/3AYglKTa/ASETKaGvMJVw54kYb
4COGwLmvzw3qoJ9Wn0+UKv9u8I9wL7rHMw8BSFvNWY6puaStJCTq5pJS54sW
Iz+bFbiTQVdvbhfOgDyDodeteV/NaaKNCRsSZpqY1LvGe0GCsT9JHbBihevi
rqlY5FnK5vKpFtZuZ6m80RU4h5KSGhIz+/SlAh5hk+zZGSLOYJlbtJGoK3X9
YBw+tQgc6yipwbV4XxxOh1RzLwMTuwEeYmUyuZaBkLNkuLZiXoJBSWFFhk7V
OU74xgySooLE654/e/MEkke2ZPwa5hYfyf6XRBrwc2E/iDxIhn5dhh+QuPSl
BvfyBbqDgqAtnCLGxoOK0POUKnld0QFmlx/Sp4zqQnvjjUn2bM4B3wyoYPhI
cftWHqsuAvg+3+5i3qrSZN7AG+Myalv9+H5d3r/qNbGBdc+08Cp6LZHF7UB1
ClmEs2I5soxdRbvyHtvNVLWfUidC9WRR/V6Tgwaygp7/eqQ8PHaZqm6sTLyf
HONaEIZHz9ZbPqxxF0kC1+udCqWunh/uOAhRQt8bAr82GcgTSHJFKteQ/caP
ekj31v4b6AU366ZhhA/N2hYUskw5lpJo0txtIctVomfSfo3k2cLTM3trbvvq
Nhh9FVe1h6deMsW1TbG7/FnCrpvESdnK4zynUbfXG2bjfmglZKNHUxs/NZgn
rnmTIRHSKKhA2S1lSsDc4mL3ME3ql7VdKGZW9Nw4u7U7LiKKA71amZhUDfCu
yA8rZlx4zIJQSbA30PsJO2Qwp06jBcbrX1CCpmION6OkvHiCGQwFgZe1jvJr
n81hbTxIjPYzQzlQj9Q6WTnQgXeNqphdaY9ZWky4968p169YD0ivkGX75baf
sHequFyaBn5u/sJD55Tb6OqMmYadkZC/azP+R/VFeuHSPvnmzVEizBYDJpBE
OlU96k66J7X9HdfVM+hH+AD1zeUnwSBUU2aa97ps5VburqNq2PTTJw6vY9sp
Z4w3woruOZq1Y6IAanw+IZzQnPCThyC7gJUgrtPXpQtYFXcBQImt5WAzdVos
W8DfXhjTaBw9claeRXCV7VW2P4BusZNNYaaSN7oc7gV94fiN/tl2CsLAqZXJ
7JzP/IJv12EAgDv4uynFAQCp9sDoituljbKbqHOrdl26taWHcqdiQo2seksG
2ONhuyRBch89ImTXUj9Ly6btRIgY2xCzsmkWhiQVNOKMEc06SQ7gGTrqh6gb
ccfpa24qRgPqMN25aXhiaARlRoeOlmDPxrwF0r15pg6tyRtAzz1RdRoZwXGw
Hdwfg2V9+xcpZIV9Zn48a5EXXe9ozLAUStQWHbpACPYabKmzXE1+SrLiAKf+
P+NYemeWHlIuv8Nj7wPvMUpO1VpmpskUQgHiXgDzVq7tnmBTy8JnKOrw8odi
3rJ8EQtUG6sjLqizigzKwiK3gEzYxm1z1MYrUZrO8YeE9Ay0dJSGxUKP5cOz
0HRS8kTSAUgKynMOk4GQCfHvb9G0HdVE0WfjNn+jAGKZLZy0SFAsEQjOTrvP
UD+s8oblKNUAdUCAwIeKXK4QJccH9X2DXb1HZmt0dB7EGxbRhGP4LGGWWo3i
97SpwKqZHdN/if5hYGZXVJtpubg5zBVAAUfQPibfvGK5zL/PK68O9ElzVyaS
H8vw/PEHKWRiRb81eDhg6/sb71wBL87h9Go6YXSBf6wcBSk784pxCIuxK4Sw
M5fEtyKIrGBcUjAA4imkCrLRIai3zvt1r+1sqmCDdFlKnFoxtJkt/D/sxa0R
AXx+lYaIX1aNG13bOKnIcPDuKqQEMFh+12JzWkFcfj3xeS9Y+sy9bUuC9Ae7
Gnq2NjOvnIq8R9alEFoTs8cPJ7bgnXYDniTbzPeKiBzWLEeSqSMcDILBRjwy
6Mz33ugddAOOhTBRJfM3mPxRl6O4ov+41Rve13z+TdE1zAwkb4BsLbMm4EZx
cH9SzX5OX7bsR6O1Oc0vZYdEgmMydtBAQVweTqMJXvuugcLYGNt8mm30MUPM
dlsllYoWra4sjPG+h+6gtl2xv1hpoD1riykwfSeHcOeSxl1J7voxVoOJWxbF
7yQTjHOmhFr6klO3vbe60WnP122958sRETwG/U/lAzg1rg+f1kFyr1Py1NnY
g8JYkf7JjJ/VB8A8hBLOou58m8yBRySd7ux0F1wf5mXZPLkBXuzKKPorAN57
FuGkJwb3skk2jJiW6JK5iElndmVnmhi3Lv3ARJViz+EIcCdUlz0BYtaOHZMf
nXTz1oB0NWmTx9V0sIGLD9Zp6/ualusyMbEpmpY4FVUToCleYJEKvoQzXY2i
tISYA3RWYXPFP1+ItQK0ZHo/fG+V3IGelBcL34ofKKp2nXkaycuianrrp9aQ
iDps2fRbBa+JdcOH/ZRk1LppIrzOnfUbdu8c6Pub+C3UHx3p0MHi0vQWYvpH
CZKlRvrg8AdUb09fvseBTXOraJJN/3zrSS5YMlthgW9WMG9L5l3UEl7sOGof
4K78J82FISgPUOA1byIFWXEDN+KjpPT7Sea1GMSGvsWgQcsJC1tJYHLuMyPt
upqylNBirtdv6DBU+ntSHMay8hVThl9lMxWgT07JH9MIUhfnHD2iZERxV6YR
Q1/znqElViBXUmtljY1Q7cwGcnoArYnLNlGKkCfgKhD1w5GJwfbMVXkYN3gi
Ih3hlJ8DmXdCvQD4Vd1mVN40YFLKA5k99X+vF5y41ftd5THX46b6+b4mqPSk
Hm/dlIiKEDFBJRYV6JAfZRpqIHQpBSn9KRgja6WP22q/But7JUGK55EPZFBF
ZCg4TlrytVi+vVKxQxbN8AbvqFIgbZDEUfAGSLc7IUr6X+0ccscZDNmyzdBA
yyv3TEfKUs98oph+7keWm0OZmUqOFwTU4ZGqIXqAM37D9QQQHM1gqBuH5ZJY
5rMX2RwLWeJ2OnTg1cInnBSYxaoZxBmb8IVg1AEeoSv4A6QMPzyldvvNnQ1W
XNrKVIKJ4aAE1ohhfJXYwSdzdIZlPiDVgFIoowwpoIUVOo2ql9p54lLGvJdZ
F/CK9jHf8vLIhQUk+NKdiQYhVC78anMkMkYyteJC5vMqF1R7jm80WJnti2y0
ZIn9HDQ/jY+tzjbF9LRZ+jBazLw496eA5uLhSV7UHLfdqr6OKeIEwV3jwI75
pj/8stYkbQsvYaskVG5foQCArtd79AOLZm558fKFbd55334/1vZTjTGW6aIo
R+emzLRuGODdPcojDndnJMjbHN/a0GqJdVrNPIQ/3SQBwXkP38gm11HoCYDS
jUq+ruIM2IbSOYY65gz/ybwfDJ2ZSGafCtEsYbEOC7DUpoYfGX8qNL2EGQ2d
9rNkwcPELZkkI6sy2uRNcv/hy8ax3nQlMfav3hPEwTRSL5oTMK7Z3KWt/VWk
/eL/gA2+2dPljunx9AX49KG/TeSZzMFB7JgSCNLYEEmpKaywwzEGtmc9SqL5
NKaj9E9f0GSs/gOCuOCFc/TfkN2CX7GHiowRFQCrdH65XqplEmegisq5K6nd
wDcdgDIgMBN0ND3k7LdX4oXIooMgVILx4d4uYRRT/H9ImD8zKNDXfovXWVhy
AX8WAVDLVuH27UmEQ2UZKH17i/K96bchT47zYmaybYNOxBAEXns7dKRlMqky
H9S23rB/N8NbWLgaXJpwMOexxL+de0RpD7guT6kFSFLs1O1C60CatHduL6pz
/+kl/cHOfsj/NOKZP/Zk9tn6p7fQJ7llBGezEke0Vne8Yax+d9mSRfxRMLBL
Bf66/8h8vL3S8HYAbv2+6KX1vZnQ7LzZCbIuTzpNLgvX7S6AwuAHQJyM0F2v
ztXMiPfUJ9rI2EFnQq9SuuW/snEHhjRgKeITUm2YIAEDUOEyFk4GO9lZTu+g
XX75VqA3cXss3mn5SuDcDIO5f5t0syfcbEcxDBi7haQ05Zzyu5owx3hg08Av
pw2kJATqmkIdOsb6dkHzHEPNwRa8n9esDp5ewGxz8oIPUsH3HMsNMnMHgRqO
q0XTSjDYCVmAMaAcIQTKYgFHtHFaALkDDu3gWM7kdG4NPqhs7LryPygx5lkc
CtBUYiFGTWuFTuk0gFxtCEb/LFCfhtv7HPVtVU3LExF3+AErP35eKUfcFHw/
V4Q2fyYmlQzrS+DIfsceDSQFOZS3FuFyaNw73smmJfYgJIBQDwI3KULATKM3
cEqewoBrJXy6YaOZ80jyovFw52q9UFhQfj2gWwIozd/tw6rjsmM0E5WdfXrp
ZGI+APpQlRI3e60+tT36UEAsiJgidccuRE8YG81tLsl8iGnQPosTa6crroQw
XCk6Uu7MUbHfECQ1TZaAI2v6y0TbcT7DZW7ZysCUZOMDJVmaf1JkFr999eDk
9yR2z9Z885VsqxzNioAViYn5i91DVBUqskiJEj+gPuovV3PISduDpyFC7Vxm
xbBquEOY/+8bCpZThtZ09mhxfOUyUn4i59hjKpmJ6gJ93IKDcDbxhotWa5OX
BKcP5aGwwch/4wDdh2ewIzfbbsI5e9VbJwurekN3z2dimcHdUKMu6QeU0Dlf
85f/fCTKrD2mfIFM4DG0BXdFpY8opcYwqUJcn6dC8ftMuw7llhUXS+v65Ed0
+39A3lNj6B8IAUU6zl6AjKKImdx0ztMxbUAVOyPLzGXJOTNpGvEkdv/4Tz4H
hGfTxckOsRZi7LjTjwuQOjy86a9oMULHbzwKOME6pvCFOE58T99orDZq+AyP
LdSISAZZZwt+73O+UHOskpKbmy4+oP+0ZbTwLCXmGgqmwUMGndTF5EHY5GbG
5EUq3nac9DOxqfGPIUq4do+1lf+CBMQUzvrcuLeldg8A77nXqYJmhIBdwVU8
NPbqAEP3/0zWymtjmc8Wi40bcUGB57FXkZ8Er9YU49rduzcPNuKa1PJaZk6n
qyagIhGXMZL2hrrYsUfoelxS7dn0mUIOjlD0qiqqZHS//HY+4PaQYIi8uuVq
jawTNdBkGlnnuS3VtQOt5otBG2XEKvzpSE+/ouH5t/5nZjIN7iH1p9s/WgG8
ak091OwuL4+YCip2CKY7PQIo+9b1Gyx1RK5WZoxCHlmO1OjdiCmtXdp/S3lH
JNY3Am0xPbzjxZ1LYTU7VYxj0T8POsS+KIeI4yqlBXW3VSNjqSKt1KDrmDGE
QSGVQ5yCzOEeqkA7JJ70/mqAlchRriSonJEbYFS6nhozxZZcim2vwdh0dqb1
eyeTFzTEBnQOzDoHQt+rsXGtoTcsrRJUHQQw6FfIHTXrfbIUvqBk176plnTp
PnuFPOxJDDT7atbdi6hwKsYRpjiYzV5D2OZN8iCfMcDX3XUhkKuDBGXP4G7R
jxCdaSazMxRqKcO//pM4N3k2N1H44Nat1f4L+F4IDm/ajk2jL5X2GIHPt1pA
P2TamvqMHD7P5F2bYLxjGZSnCZeAP60yT07vsbCd9Omnb18L7uR0JKaCccMr
BHzRyGKGComCEIEoZvLgSr7xGRSJeWPjsPOvaQD1x3OemkWaaYvX8pdIcEST
AfwX1NAOphOMk3Fvk52EdBmm/EYR3q/LUtDTLeG08shvKuZEWX2nhi5WhKHV
CA3MXQjTq30NE2YK8gaAqxh7dgHTXLPLaqWiLAVwyr94K5HODMqI4CtVowcK
f87vRd+Kr3jmhq11M6thCZdG8CxngCBavMH+3aCD3AcjRVgi/DpxWhTPwx5W
Nt91cCvbsiM0GhykBsHReLxbJuWsUeUGpxiuhI2DBWkvvMpnHaQgR/ojYxlw
bs2vIe/c2iPL6BdKZKRvf4jiXMo7CZTEMHBpz3nvkVQmfzvzxJTPeyOKsoCG
MhiUCt7ftZrEqt1CoNEN3NhY5PMguBcgKdNdcXMDkh8eJXHdkg2gDQ1yxx/K
COyGe4pssC1SgGrAS1bwCsHah17hfnuxZ1cSnhJ9U22O23ZJFYwesN/xUyJB
Se6GWcbh9ZE2HthXYNpV5uOQuBPL2TYEjioNPfcChmYnT79FN+ks6S937I9M
LpKuIg4dycH6/wh3Fd8J6mS1/aV21xPmUP5te6dW10b0FIEVMeSHTDuG97G1
Waj0QJ4PdeN/MoH1+5ovsA8vDrhC3b6ynp+tE4J1QSSkHqCJArB9zAIhCxd6
EeSmzQZNSrogziXk5G8Rl597PR28HGhDuteMOH/zAh62C3oeoXVqri0GLHxZ
RnChYNlltNFbTbx78qHIR5/DKEau9CWoaS0XRoL22XkfyrR1YAGlmJrep5kl
fLDDkzipqj8qZJW/UOftmTFeZLHKLBM+Z6h02oNo6xeXLYcb8ZjGK17JO/gj
NPJh9Z6KijYnudOyDCSMRc46Lu/reJLOj6w2L0HrMKu4jZAD3gyXfxKUhShZ
OijNATCjr4axHPzfRpaNwWLlyc+aswTIBwJfIqngYSnKp9QsFiDSHGtn7CJj
XmZD/UBi1GoX+0RPUY9D2XXsxtK4TFcCoYmDiX0tKFBBlM+k9bNXxRJD2kls
kKRvfWc/lWHyFhKoYD4TMqFkWS/NQOQ2AamS3Ii0+GLwgFlzNSs0es1J7ELm
FoWCZDY7B2dNqGOxbMQ1yRSNygnTQh/FLxnzZG51viUY05naztPICdL3Pjtt
3/Yurcl+GgS/VbIJtubnC1I+NKuIFw7mHH+XBEPo2zuNRGOPgN0l1f3UDV97
9+U4ajnB/zBCX3jlWK1AJ4hImkLWgjMUIPTKi1+TaeUtFBQOuJSjMM586/KU
rsMstGUCMw7JntjkuwQwHScEl3XhfdM7y8LRRF3MoTOFoPfrZQ1zge+BursD
CjOEWjTh6mcfowFTZ4giin7Qi0ULVHxzIF1IRQLNKzCghEAvV/lM2Lpiyn5u
qbpjd/pXLHAQ1cUPhJAlsg3m/1r36osWuUIot8HSbrKqIE2TwcVziJFNwYBo
whM4Qjfb7i/9VIZIQsqyllF/vdlJ7poZWmFDLilxRbpggFgwegqADTHCnRd6
XU06V4ks7dM+zlGXvER0uEvBP/0qqk49vXkKlY7PIwvq50CTGu38AAqK3znT
Cc9lfUeJVWl7B0F0qrIJQGwUaihPsAoTrk34JzEDtkhuZEJbJ4jstwearEvT
/dgG5Pm2dD/x6sdyt5qfQcAjliDEE+0t+KesD8hPlf2tO+TbO2YOmGu29ok1
zPEtBIUEyPzCaLB1JUyKzvcEt4p+/2bVglWCD/sZeutjPMPvyz+AW/q9GdK1
TsYmoFyNlhnA3MSsL2kbth2yNdNtWLc8feNmGnJ9IMOkMVP/e3/urHGsz451
GRQHl+tXgMPX3FFafKKZjBH/0JI0QLkKMJGwNbdAOqGzu24mpBYJtJvxf2BY
ljtR6uCqc8aff+MlvARx2k2zRyW0ZwIUwZ83/omVLkzInaXixxrZDCkRWu7V
Gi+bexZZ15ee0lJjk1tx0w3LeNPPGwU0n/5qV45b8WyoSP+diIy4F/YJpFhH
t0D340HXNwogJWif0+VQQYVyb7ZOtTuDAuNzoAFO4G23yPRHq23oMebl41Hz
XKGp38fgc+I2HB+fwbYVNfD8T8EXdNRoQyvtT1+Foq7Mf709lkcL6pDaidpd
qAhQUTryu7N0RDH+veA5ZmUOj0EBXXwATUts1HeZn3Sttd91S/A2/7fBMw7C
guUXduy26Bmnvuxf84dzvIC/9phdhfSgRNnCjCGkpmr5I2s5xOTz/iDy7oGR
SLeCI19rpJCwSZC6nRbNA2uqz/CZxmkwPknToTApxO7nYkieYvlsLeLlEzGd
7mZbLdZkUuyRcChPv/MUcH2egcPB0WdW5yTD39+VExzk15H8m83Gxr24Ypet
yhwJM6UBxsAAGoQuSiT+js6utyETD5SsFeKaxrEEdk0JrFCuw2Etf+RVLlzF
NlzLyLYujVsIkPSjZpOcC4JrqNbeUVmQyIyW3Y3ZFORS1D2ZccnA9hreWCSR
RzhDS4T84AlKdT38zrneBWYjqoiuQZXIBY+iQBSsSWRmya3pmDaURScGIn+i
1AlyECeohEwGSmH2VI4u5UEyHgv7TgDSxc3NLqqbnPptDXkAFbhtO8wu6Bc4
Vsmmya7rHlMklsIy4SgIHprLAG2t+3huRFJ+S/20Yw3SYHi6ZQZE9Nx3E1fC
2LTpmdqQq9D/ft5nOsAqUnGRNlJSu3KDPCpGYZSKeSfzlZJ4FxgZKW9wS3mW
hRHG1ECY5TNyAT7EglcIZ4wWHolCJgCCKB5yftnAG6VJEuGN9W5ZO7dR/YZq
Hxon3UD2VpPTpA95GshAN7DY1P5nf7xXyEIw/aqrzIqkjxAZmuusLcuHne/p
PTvt7lnODIx7qrHe1YjirKo20Q4SMKaQXTPUlcxuUoB/GtkGSJfEY3nrfipt
zn80AuPHxs/qZfzpnpBqduzk/3sMy1lYG06IVEWNmaopJEkqT4iglU93SyyR
wKSf7o2HG8KnbBI8SEP4IoU7PlUTfmQqrQqBVZZE9qzCOZ5VwVDoHxE9jERH
Nzm5gd8zhLR8Vws/cMdcC8SCYHQQR1y8qu+zoV3iIYEbpCXsyMtJ2BeDStAO
SXFmzAoJwV8efZTh96yDLK9Io89sq1Ff8QzOpjEh/rLgbWLpnPfD1MvIneUo
XXRas7784tKTdapKX5fZo0NInolaZ62ym93l8uGw3oa9nKKdUIZ0uMgRw5P2
a2I9giHiLxAn1/RlpwVAEGF1ngpIDpIiV7qFUQbiCjWKBkO+3nFKCcArFN3v
iMKBAwSFRMEF30rYpmpWvKsq80MmujKnvcpFHt7u9YuKU0M8ZF/bcpu9xMqU
MLsce1ooAwSQCp3yPSf2JBpWnHtFZss15nQso7xP9b+ns2rCD5G/rkLTyFmD
qfk2pZ0unkON6Y67ofJYJTk2XajZ1OrpYNysZAHTE/SK1YJvgK283n0sHFOQ
T4aNu3quPYJHaLcy6oo+qceikXmNPGPuMDMpH0o6INVm7X2AaLenXRCKySqH
JEM0zNuidQDktifoKqT5uf5gJVPUplG4KK/cWOwa/1rBpJYrwdclDt5kYaYx
M3aSD1xLR09GvejLZoTDzAmWiHn4AKK3jEvUijaqlgoBGMtcMWrEbrjl771/
48LYrvUQwdcfy0wU1RL60aFXSzKj6XXDCngKFShU7sUATj3kkOW4cB/w+usI
wIOUFm4iZTGRKE8AtrxvIuDByfpQo/EnUYS4BbIkzkt6htXAAb8D4L4rGMRC
ZOQh57gAJCdv4TC8oaGZf3A4wlKHTfln+6r348XNAmt7z8DSBQb60mSa33AY
Q9tta+GqgKdDU7L1oExSpHn0OiqUCNjCWQnK3OJ9MEDIHkj/kS0ojAFW0CkO
aYhOp2qxpi8H5eIm4XhiipAuLo//8I4Ag7WcA4xqkrOt4YRbryScKiz+Qd67
jXAmJDlIN7hEi8EgdDe0gLmy1cDazCeI538CiV7h247VtL8f+/uVx/dcu1VP
amvAs6GO4usFN1AbIYK0M5AwklsAVbvT6u7s5U1cVkxh46OYBXtyBM0CJGSZ
WnxA+6NdqESlTGOj9nM551iT+LyKqxsQD9u6McQh/sgZ6zV8ARJl60GX//wR
pQxl4XMdG91MTt/vkvsKor+4otcVhkJOd6m9LWdlgtGP3XwqWIHv0i2Ug82t
ypjQ3BiNPe9gwDJloeL39m1Bb3m9XOsXlr4PfYR3c0TeNyX8V7LE9KW+Pz4p
SkZELQPn8P9vmId4+uc8JR7jixaQYlJx5Vn0zLoCJ0TkMUQutjtR0VnfHUYT
n1fhPfxw3UJQZU4a7rrpSUX1aV6l6RxO5B8dJXYx30XrX3IDLQaCVNojJjt+
r6cmuVGmkMMdA5yzWbOCfdCPRXEWf/5YQ3MDhNAymZFeewcBvunl90fq7ZYb
PxSq+Zl859ca0eT6wYcOWrLqT5q1y7A8STern+4Jjjin7axkLT7gwmy89Gh3
7Nqy/tA8EZ/KoIVJUwIY9jaikIZomzK8yM4OTxMdcaTNKjj6oKC2+W4mPNMc
w/Wcd2zro/znYSGzt1RJqlJ7dOvwhB3V53nhErpvANWq15JtMVA3KCQE3Sab
eLYNxTvoV7vaCo3rgs99FeIRH0y6LYx2Tzf6Fb6zXkR0UpjqaBDxet8hS774
YnS2zPQA2jK1rTvTOQAktj90pMbZIv1yLOc4VyUFhyfVE60wiSz/zfyf0b/+
yqATuMs2aocJGkpFQEBzSeP2H4TuggErZAJPTU/Gfw/hy72UEi86ae/z6SFq
I6avd0v2ms+MoO88UVvInm39HUnkRrL4sK/HyrArxcBl2Nm0Nhql24WasIBX
AKYuG7oNWsPYSAXU5fdjokuM6WBzZLl+bqrPgrHh1uex4mowjtznk9sQWBbw
XMdfM+17tl5rSeBZ5k5wMBvf7RoF8hN9wE9MQPA1H/S63U2VSFc2DUO+Elwf
siG8VhEKgbg3xwzJk7SPP1ufXF2DUtUzdwZ1LqkiSc/UKT8f+1d1F+rGV+AK
5ksJ34J4jrobr81WL/UeV/C7eFFNLjboNVN3Y2A36469YZAIPop9Kx+FYf+7
lseQiZlup5UAIXDe6Jye0ZZxx8HqgdLjX2bg4fLqpzU9hx+8wlEb7izK0wFd
crfLvg9ozC9JaI/r7tONne7SYqiJ00tfNND679bUSy0eXS2jx0QGLcpN8+nV
qdwef4+++6wj4fty8afPy+W4nM9AZx1RHuCqR5aiUxo5jKDcCf/9DTCUAZtP
ZNn3J5WzWmsmgWRIuK7F0Z9FUV9hHJUNLIZ5zJOgv/dNNalklRfzilo8GeMp
T82VAZWMAwNikJf6rjGMYunAXxGsS+TxJuf2Y1hJRl0eYegPweJkuStEgs3Q
mKoNe32g4PxsshHuuf2F65ieivAb1KsS+rgOrzdRq3FWfR2tp/elRH/r388F
wnvTYfx474B3SqqWI+B1yIbuGbykZ834auBDqpcoVubPZlKHm8Eaap1IQxf1
JqRpffmMUC+nh5QVEomFHe6iVJF578l8rp7uEbKW485xRDemJdh2hF0MacHs
MrrHpD4ognpvYhFhU0Ho51rcFLK5ge2t8/eJ5Zfid3RZiYIeWxTGTgFQi2MD
PqOsWEoCsgKuNe8AYvkU55ykI2rwhBtZJfTfFeP6jitRovwwjih/XKYJpoTm
yC3THIKbIBtRmKaSkw721ogY8roDhpGhlVEkzZgQhJ4x1M2wRbYpy1bZaJup
mcTl15W9dG65ZyLodjqKSie3pofhGqKXGWEm4hXhJK2u2967gtXNe5pLsavj
UJEPSWF5bv10Lok2r3wZN7TLn+addC+WR1w8UGNphDMLNr99w7GjBib4XPcV
m5+FfoLFH6CqHq7ZnEhSvoNITzaizV6iv6cERSILPHPQ5U5vyO4KAmc04Dkg
zFLO5mF+Wv/U8oeF37e/+0Lrhl6YGsF+KKVmHuDWQRarYrp5K77a6tEoCXTJ
P0Sgrp/wSzIlIoV6ATWL8n9s7xIy/HFHhNwJO/gvKNPhyvNHqSClFPcITawL
kPCA/J+RQ/m7wXgZi7DlqnyluYVMuM2mNknXmjkpP5ReZ2Tldyg8IHgG8Rqy
jH5NnYw8XWM96nTOqDZj69BM/1SPaSXJPVVrRZu4EjTBOFfUdRkNasdS5MZs
RpI8H6EKqp6dgzpmqE8u8K/3cvyuzDY8yBv/N8Pr2eIoCIoo78XT8VNTU8bf
xGrkUPZ/GbSWiheIOWmdNz820OEVNRwhbLqKzTyANmWZz2U3eMIo0HCn3FAh
C/WKcE7OQe6LOR3kPU4acBf+R3h/jjhRjqnQ5Qh59VFEpFwedkKCRs7c/7Pq
8H2BVSJLgcfbb7wcddjfUbraMR4BmqrweukxUL6IVZKA/ERQXOVQ727+qcbI
YfQ63Au7eVbx++2iKse8ztbXrkMPKsHYN4i+BN9K9cStsb90qiMQ9UO/wlD1
nl55+z7nlWD6gCAlYQDBgEAeJzvj71n+8s3SiFOWo7f3EtgVJ6oPNv4fWf1q
8pWX7w6FoFxj2XIlpL4rSlV8IANKPV4TU3DxAoVzx76t5EF4uUYK7f4e2ykf
kkOE0uUYmmO40spOzIwRo+CGECMCIiqmz+nVAMRHlMlPdZehwMnw/wHOdRwt
Az7s1WkzS7D5owOLkOhCpIxJXAeQAKKaljNUXBQuZd6+NbYOm4h3tfUW6nWk
9tFSj0p6UzpafV7wuToYyo+TBzqmu8oHzbAAYoP6G3jrXXEPpTTUDhqpU1he
uOYY2cfqy83LMulagYk+t/SQQGZcDtElbTKbjmI8OoxRSXu94/KUWr3zIH+H
jrOwS2L8h/P/48C9VrG8r6zIX3Bl6uYm9PVf9Z4ASStaXgNZgVec2wdAPHyI
zi2pIc26arXpq7gmfXB7Pzv7vefBIXuZojZijt7MUpoeJYs7bhJp5W8An+B9
qiqEmCHfQywS2PPJjR3D6AiMvd8uLP0em//nSvInm4KIbie44CYzbDeo4JUF
qt2dqa6VUhmbaMUCwonWQVEfRFmu02yBH1l4eBzqYTnPl7d7oAyRNxCFEauP
VraZxQhFjE/fdzqyw+Ob3ckfrrFKdW7uyCoV3aWPYtw6znJ6kCvZWH5DO3Ov
LDPduaeIvW7gNay1tgHbRLn7EIeWAhNMmw5a2twWSn0wdVcMEKSpjz7g6ysY
OejL4KCUq1jOgMrgCG0k6KnTTuBjIZ/0YnY2tNebasGu5W/5YTvOBkxQTuh/
2xrUvp3hYkQ41BqMA3bWghWvr+CHFUct1oarn5ed5s+Y5K8tSz16R3lnrYCz
dwcktkpEH7mQ31pPC5CQtg1BlCG4oSyrqqa0lfbkjb6uqeHaoK1PRE2QfY4F
16sJzyVId8+ihTuep0Fx2kLRgrj1IyybwWW1Bl/0/fgzql+FaOcBJNdk0vcG
jeVMx0j5RFVX5VKWiops2aXKU1zerj+5AE0qjAKsmiCXkrxUp1YxekTUHsxt
S/8W6qB8YH0sf3fk0LbBObOjD4qqgbzm6d/VBhxifoBXL3qmiuepT4I24nLw
dhR09f5KvByL/gmePR82G6pk6RmANMoy9+2/sHgWGNU7Y4wzLQel0VVWLFtV
u8E3r6oPL7CDT+ywCsAmPNEPD95C0QTg8yAjpXEIFZ8ob4BUkWZPHSXwMf2E
vaJSIh93Lxi4SCpnsupjF3wxP3F4syDH7y3nhNCt/nXjoMI0InIxbf0Y1ZfJ
E+sI9Wpt41YQKS40E25xJjy3ghFF3BkTbtQKyAz6gE59L18B6XQO5p8Z6O63
6Gq1Zkaio2nXVyjdXtH0zpTa8a4sHDDZdrEdF6w5ERb3HUTbtzt0HHwEHa24
3vfhY3MWGBlXB3ZvH8xwbCKC4Cxf6VU73mj/8j65T4L4UZOR+uc3ghn3HVek
KyyKgjQUPQvLrdaDz5Ya9YmULjLEqlUy7f7znKmf5M/DYERWWX+ZQHuPmw/O
1JPVGk7hYiO9vl8sdxl0TqcxUNkdkEyKcZSzi8ZV5/0z+NJEBdhEhCs+9MCm
YtJ007mvWDcPEhg3RUMqcuaj4oVQVghcSkpeoUdYUTmsEJV4hy91cUZLknLu
dSQeC62czYI3QaKXbAQbvRq7PowzjpUlC6J1vI2cTKSt/yR+0MUlYXrucQ96
YUhN5o2PNlp+uwxUkIWaGtx8z9QgGkuGVXzElYH8WiRP6HjA1hQoo7nKxJRu
fLVF+qRxnuXM83T6U1hGpztbHReL0tEgWeqbKEuu3qENnmWvd3Ii1f0ke05M
ji1ePt45KeitL5/zN3XER8kwt7Bx5NkDJvC7ayFiLBPCFK21wUvvE6/LpDKj
g782xY3u4P77r5ObDhcLXcS/8lKT73idcew6fczUIYU6XbSY1C4Y5z94AYCU
wLPjuoJxzhAx1RI/g6XKaqoRrqshesXMk8/jXcAP6bkHJSYxSe1WBrhR5AMc
PfhDaS3f3RG8MYXqEx8MS/+5gt9l6BXhU2X7Pcy9JmgnBXEv7/rZUpU6SSW6
sP7VjE2gU8XjAYk1Zz0SK56mfyZsPVWxbXxRLi3IuBXbJZOPmy6KQ/ddiIYG
avrYAKEkmTRVh1talDZ/nROT7kxEn1FUxPxqrc+WFN+Fx7J+oxn7dsRjuBWc
LcTGEc2At3WUFUsGOQVC40dmY9z5Ro9JXRo5E26eQWXRucR61LCqgvub/fJD
kRmQDksF10GSdt6CKTBEh7VFEW1zCu5Eh4Qg+i9yRdpMKo5oqtI3g5STUjiF
ZazpyQhbo/5ovcNbXqjEeH5oLdV42TvOYuxIkc2MtOGp2njlRSJZkgtlCOcN
wQr6so7kp81ArGvYjRT8d0hrITwwrOi8a6LFUy/c2iJBj9ChPd3kMpXRd0O2
CeWyRB7Xa/BHvqM/nt3Z1afus9eamlUOswsSlAEv6F1J83T0uIC7PivUSBkm
ewiEfNvJE8mg2YklhXoEJpRQhNCt/190WhzyReM9pkKGGZZ8fuAGKBsxEMCK
1oFYvZUw0fjYxbakrSuXVUYVFAOxgSI9gTGVrcF+hRCu3D059ME3LQ8Y5Pv4
9VLAlhxpUo3LRn/8rCdTQ6rTzAl7pO9ymnVRuC7Dd/JOT+DXH8ccovW5Q4Ib
h44Pnv6aByTvEE5Kh3WltTYbf9hF2crlI/3WtKn9U9NYJnpvVg2KOA/vEVa0
bveQUV15QNB9kKAyISKobrB5ofb1k4Zfjo+BubcBiF/XqLfsrXv/pK1KLtUh
nSCdxuACI19HBOH02I9Pju7rO/cV04oT4T0S24oXFV0U2jkEk/NXrEIRb7+Z
5pHA2VQlZQLFInYfIc9l2K1Kg+PqEj226fdgb8JAAETATA6uRZGKDxzLNjKz
4nhztiGGIhoSfDHx4VxO+XOnS8gEo52jjCeILoP0IONoLxFRQvHYS5puLkWX
CcKWdIUfyrO3HQ7HoHkrHvnJ+04ug507bKFw83XVWD5/AEgdJOA7PU0XE5rm
bO34bPdK6W2yJaSMJLHLFy1QJNKBI+79aK80DO+iVJndJVyiz+o4nV+mN1/K
L/l+6Connc1o2ArHscsCWcj8HFxYL5JcfO7LHUmexhkyptJt3hFvJD3yxVuB
s/7pUbAyA6a2p8rc/+K0H9oNJ4BJR99TNFyIUp+Q2WSrtlfmLdwGpcJatp/a
jzZkGXudg4NB+6ju8lQp8Zm0rZGXQI9OGMCR7gSxC+wkFZLOsabD3HqSvLK2
terDY36KDCSLHhP02MhzmUxaXjfgDvNTaNK7p17hgPLw3T7b85wdwpEUwEeZ
ZBa31Xhsyg3rfcZycgOU7hpObqzc8vmAxDCXQP10DS6oZdCEgYXlnVMo+uLm
A3r5dJNV6U1RcRTYLtGhB66VasQvDdyT2mIoMophDRys9qJLz2Cuv66/o/7M
LjRsmI8DYBy4/RaFHKdhesRUruXUg74mwXEwqibsa/cXMO/COfOB4CzVdBqn
uxjt19lH74j4mGYRiqU6usumQlf8PyItcZejJECGBDZKFf++qLRizNTziR8n
V7Agn9Zfo+cpi2wWxWXxNnXZ8ujCHhE87YwgqgpOXpkwnaAbJr52Eg7F6tkL
IUPgQ/pO3I+c8LG0ovMtKkx/Gj8VrJQDloYoupBcOPiMBa1iUeL0O2MqQIKG
xX/8IerzBXXQSMY7Z0pJrVlX79Lu8DWYHpe2zlWDy2Ta4kYKSbEphRBb+//f
Dqfx3CgG49gPcMU9/yxYEPw5lg8raRW4c9+UGRBbJ8t73uBgsl4QPZXfkvzc
dZCzFa79wjptxqhX3rVuXseSPYO6f6mwixZsoUYBLDQu3hnvxdIctyMNTckU
YXVWB1be6ZpkpVQAs5NFNgm5FjXQE3H2hqrOfZu7rWwiefWB4yTVwTKRNT85
Aa3btnWreZ+YqzgShTCArUoOECRLjbY8sngt8n5JR44aQRNDbhWblYCER9at
Uz0a8Z1CY3+QPH6dYY0Wc+klA7dDLKO2fgkDIOEuRCAfQBm/zKzJzsVX1xMH
98TvMOn+5nvr/uu1HwXlTNZ/dREt6ZGPuK21CP++9/iLZ1UEMCSPQiYWXJmS
MD/rJ6Stm0bleMpon7dXyVhZXJ6LuU6Bkx9z1+SlVS0y4tpKboUbvb+dbITd
zvHoYjfcev03hvgNA3I+AqRcgrDS4qh+MGR4oaBXbmG90LjW2kT9Hl8ZvQBk
wqmc/WUT07egYHXkT9AfprF8QyXlkZ+tJ1qtratGw6urgjmAe6DcmdWl5SPL
uU2eWM8MCe9OofxUbUpfG9CKkNziGkBwjOnDMICB3kVMpNH3+PorXYnBZ9+P
iRHEjMzBvbXkq2RI5oNV6LyVKQaKdRQy4wAAsR9URmkOIo1jG5TmIq4a+VyN
MYZdU7rC6bylScRpoHw7Lv0oX3AesFvESXgz/9socALkeDWXsyAWzGJ/CG+V
/cs8vIn2B/z95G4rPJRngK0m7hRiDe3WfLt2LCk7ylv8L4JBBGX+6/Tbsr/w
3sYrGH3SkBNmd8ZKj7Ux7Bm8z8rEDmoi2ibnixohrFMAn6XK4r4HWXkXs4fM
NzhZZcEtDBNg2vAfi533zDmnuVjDmezYVThIL+aJc6RmU2Dp02r0Nw2TDs+t
0u8C0y/5snZpVdViowm0wnv77Q5hM0vKXB44BbjD2AwUb1KW0d5U62nRoTJP
jRWokrFiQMBnZ+zl0OD3V9NfBpmwFIiEaGHB8qNvv26twB3dl6MXjPxkgy0X
VUS4V49WDqeVCcJoq7s9jC+Ko6hsZf61F3J6YoRyLXx7xZH3Seo6Hf3lat88
be9NIieU1hapMFKfwfi+bb2V4W0OUIbH4rzPPBgppWSfKxkusYcXHkVaP+wP
Tb/rxlTEWD2V8ZkiIgpqBYu7o8KZ1TfufqRRH4OmFoLw0iXL9pJDLTFOJ9gZ
4lV+MLYp53MRx7OrNwTLmYpphgQuqYTO60Kr1kh3/o49+WWUXsrRZzS0UPII
PwP5O1FhULfqS5KA8NS6tDpY45+cwaZ++k1MUVPN6+uOYjVthCJfjhKp8sbL
Eqd7NQVRp37Z0f3ETo089KyJDJVdVUV6AcHvNTjeIsEZZTYcT+u++/7OADUn
VizZtccheMBXXuX9NTK4rbXL2DmeIbsq/hfcC5klGGgWY9BTCDXXAIz9+UBk
cGjUSjTyB/uBhx1WMVdjsOu5PGdgyn9uWAyBRtj5sr18agmu9sci8fmT5NQi
ACk4+rucozakb21RGo/Z9FN1uoWSspAh+DjwTzN/mju8e+75FkiRrZXCHQFK
QlEmVdiJo75DxrFlejn6cNTt8L1hTdOu2qPNyArQZuqQwRQEMy8YUFd47syB
UNtflHKDcifFsxxVzRohEo5T1Vyr5exTfiIWnsmscMZpX7yFN7uXhhhn+i84
1H+9CIIi4UtwUznV+3QFm5wqqA9VuE+MbHPnfkqB30bGk0KqZ0f9J6VF6I8V
efCxg+60vT1aNHFJdhEkwClou6iIcH4OM3MK4iv10+gsBvVC9vW25mZIkJGF
Qx5Awhk7cDCVtJAItOobUKrB6p0iI9/uONwmjHJvhJwaPXS2bSu/7NVHr47u
CfR570C2wppPU8Q9Mjab0VFbzo6dLK/lAUbLJ3GStlrtaqkYzVoCHW17pylO
ABuEawHfZnxz0NPzRCyM6qWfMU4QcwdNRg+1295O9rT69yVwdPrl+2jjuQJZ
F4UbZBtFNAocfiW2HL6s6YEUScI4C3Fp3F06QsL0jysN3a9tpQV0Sm7K3FCr
V99HLJjwDXniKosmtvXdL5Oq6mfVx99YrW0QJ1xaiICIcuV1q/ifN4K0cQrA
VacazHQQCloTyubaKUfHzHlzFCsJ2DiHexrIqqqOXQeSbwU4ERjQjHYfA+Zb
hMX5cF+T0BYnNIa7pbH0S/bqJoWiwV+80oLiGJ0axKTe8MN7/5u5apUDXOTU
xwT2KOFaA2ees3qNQody2Zp+9KMC9sfUfaZWHU4ROVH/vTW7H/Po7Q0gF7XC
E7Hq+Owy2hX4hvE4jA63f9oAG7YlaNqS1m6Huo7WQJti74jLKs9oprI2T4CT
3d2cvjdoThK0IGWx8eEgO7QTFhtFDbtfKDl9rHaZDZH4M30RWdIu5ewYMflQ
LRSq9mvoV51fsc0CghqwkV3Vwivzw3nz/cUst21Fb7+eQOWvWYsSW2OokW/W
r3s8y7+dfMVPtVpeAqI4E5JXkZLi1X/vdkdifbkTmk0OzB1bz0rC28dQG9M1
PUOp4TpIxNLG0qQF7l1TWwdqCjZ113sWphzDiByFBy/fC5/TwoU1ie9KExDD
C7GrW751jMOpqK37J+8DQGv9iEzJ08YdE7m5aZrYrYjycCNW7xhXOIcSatUj
eKKGx+ypTOvkqao4dgnLCnwk4qbdW5JQ8GWs61B3T4Me7mU7bVw7J1uXmPiH
3wH5/ZevuoAA05MrxqYdGxW9CQe2cabASt4wD50fIKJu1iw7TMXVeQrweLfR
LDg3wH1YwQGcgtoWiCX1DnFwdolhh6FWX7hBOJLyCmvtLJaigmfl4c9mIfv1
QifmtfbOUb6FQDgM5+GtWQ0UBWy5licLI1OiBPs9Eb2FbDniH+cmVvSKW0tT
IePqVPXpowNc/XypeFZXKGptVoQxBlWwBIA0RsORJy0Hn7+U2sMBqiFOOAXX
b0fv5qm5+OegUljF2ctbUd3alrvsaJRDJbb4qGbdc4PtX7NJwLw+x3Rstyj6
fJ9IePz6WFjBLKX4Zqg3q6mrP7fSv0LfarAK9Ytl8bjOYhQ/wP4L30t/fYVW
bPgX6a7khh1wCrxrQN/OER9ErcEVOV+oQlLHE475cg7tpMD3oTPfbsaBK7/5
MeUiZqY/m1p4AZekvukkaUSVJOWARSXJMN2JFV9DxbTy9UIVKGXFjIxggHiP
IDnPF/rZS1dccZCLHeyZ9n74RvWXNxpvVWxvFMsVgfylein7+cBqyj8TCf/f
bfgJnAPYcTeJ4HbHvnxvj0q8gMg0dh/1WGD0La+xXDtnrEXOFJpup+wSu9nr
iTPU9WtGYIrExPG89Twk8J9TLyB0d04POkj0hxGcPP8oLSuV3afE/4wAW3sW
nujVPS0/87+ZKZGQqZJtfWT++BeTTidFhetHyRtz9gMb0svXxQJPAJlgWLp+
hMn3UBBnQ2QB27fv4/Hnnt6TsA9U5SWVuIewhbGtdAsRnwZvOv0z9K1noW0E
P7UVyQQOyIj8Fj1S4mp8P1XZEE95RdSTzFbFbk1B8UyeE8Yq87SY80MYRER4
4uDp9pKbjE3Ce/Ounwvt1P5zHhaWjqe66A5H2i6Gnbb3CRUeHTDwFg6wuhgk
Z9LEd7BCgeNBS+QZ3WILvjadMwgt0vkFUl+pQtWzPkVx6WiJjSYIqP4kCrRp
s/Dqr3HDCRQXufz8/NgIO6qne9lVDy36KRs67CXIjnDzC3U2BxO1a7nAAa4G
Qk3AzXsSfLTjfsS4UIgFxidjlhiCVfTa4f3sXvL4WLsVH6YGtXhqe0KymiFF
wd7LsKDQUhIGZkR83ahf21ub2zyVDxeTbf6ujB36/TDtY/vfNbGVhy+bkjAz
S8xi/rcG9d0Wafox7dSmpoOhLoiNxXbcmV0nGNvxHWhfiWJELE8pgkRQWyRX
vzfnUnxKp/HzVJQN01ppoMV45PW1u6PwZr0iq+rAz0jv89Ln/CyO2I0gHwXO
IwE0NUzeLskRsshuFeh5weqaW1+J7ByZWy+JihqLy5QIaDfMglAzNhlxYkc4
KBdJ7WILb1vi0c+/jNj60j+qsH7UhFVTABUNhMP+D5Zr8DESRST5BTMrHr6F
ljiJUrBi3t1GqKCeZh7nXtgPh8KukyPVpz/pOyP+u1FIMHztFc2+mKrjWTVr
0Jb3I+b8ukfTdE4T0iNfyC6y1zSJL1XMj/m263zBgDuQPEj/kXOd6bAOklP8
WgC39+QYmaB25pP6oMaXmY3lzGdxT6+7YVi8B+w4t/WF0lRbPffGyIMrNVB8
PmLf6+z9sSpr3dvxUCtN8/7RWO6xBt/gwCKkLXQgpWylqYYRQBps5AH9P7B+
XAHyCrHDtcM/leeTFgPJcUpxtVmaBtF+pTG1H4svwtJUCWTJwUdQRUrUyfre
KVYkmhXMf1pZ5Wi3ujrh2UXnfyVRygKc9Ctp9EBR5bJ6J2pMAHdO+0Xrbi4T
5zgBfpNvnJcSwaSTabcJppXrbTI4vJNNp2/HfRG7KaklC1WUYWJR48jumSEZ
lWo0HRhlFt2zVUop+76OASfMY5oXJKF6O7rAk6k2oTOIQUKxqWth2xfcnScp
AS1sblPPFebJw+sv6t+UfJGjvQk9gb4JROUsctseGYNa1a53rpibQaBp1VMO
neGNqoH7uMHrWsr/W6O/0U9JxQHmNd9mv0GBdumN2RmaBd4fdRG2sbjhyZck
uOMk5wAT3pceaCDQG0DK+IP5Ecdh8goLE2fvX9SyreR6Ig4bIg9dQuIqoUGF
zSQUfGyXGSuAtDgEI5NFqjLGwW/3aLncgCRz0D8VMYS/TNfKjj/4yXmsKszk
v1SPZbGT+6rgFK3W/LgMKBjtH+jjT69W4Q13HVRqw69OroF+wC5qsMlN8YcF
mQsHGl1zM/jfZ3u44zScmZ7Huj28Xj6PwICHZgI09OE4d+oetuYnDdMONzuW
OA9hbv/Ztw9NarOuapzyBu1VWrq19dF+QvNJXcOSSbgxQM4QPDqX6G5M7KiM
ZwcpQC7Ivpotpm+h4jbJqYPVFF6K/XsW9tiy9KebALjOMwO3vqaEttZDdfIN
aa0j6hAHZLqjIcncrgTfp/1CEMAmI13qX8DJw9Bx2uxityw4VeKNERDI7Q0s
QYFReh/1dLnxUN6t9D2wAQDB4WRwJIgEaAuA2LoguR5BB5MqcfZq71MadqWT
Dm4lk2+2yHNf3V96U8dh5hT/xpOZxMjxt7a1S3netOaVC3SeFLclHrocpHGV
vNrA2K/pg1kobSK5joKDejLfWftdiWvNtqLwtixZ2EiVJW1hmjcX4+8hIA6d
xAykcAgq193XpSskCQpnS62Ps1dpuJH1XIzCVJ/RAr7WNt2WxKjN/NhLY3d9
jUDncErMY1scltLx8tTyuN/P8ZjkjLoqnf0qFWq2ZWVK1PMPnawqpe7kUh19
UuNUoa9F3WaQcP4Xk6XhQVog68f3Jc5FgnY6KA0jLiCt6iow95qz289WbFTN
HM+lUjnK5XMDuIDh4z+zqCiL/Y97t1IXx3mPdH5Hq8SyM5tm//SKm1yd5M4u
7XHzlOsnnHKRa281VcRUUMUZmaZNkstfdZ5bIkYGy7LKRE9Kwc8tRCl+WA4S
HTCUUWelz1kN8lGCv1tEAjQZ1HFuNja3YwiR77EdYeb+58IJEvkrVtWwYo1y
yFY0kBia5oNzPGRWTBdrmvbnTcFMp5/bl+lWi4E55u1Ybi+FNAjQRoGVQQ64
M+YyiqyVgOq9bS94HGV/W048iXYqTB3RP/GfA6yfnvWgu8XMuzHWLiPjtq9y
3sInpBOjaj/Ft5lVHiQLAErNlbnh0hDwAKbc7VJfNWyPKoqWnsjilUs7kUK5
0eo/jiSS/gBE9DV5Y5DsX+olyDdxjSCipJ83I2j8eO6tHyiFa3i783OK/4Gj
/QIUJxHuKPeDwVS7pftTjuFi3HodwUJlDtCclwnULZwu7+LlsgTxCPptlGBG
tYoY1Rw4qd7k8mh3P3H1wIv4A+/uFYzP3E+kfE7I5Shc9AveTLa5wwXm2EBY
uj1kuCAk0Hs6Kykqmxe4LuDq6gVs1uufJyanmes84ncw/YS2RY2VB/yG5GuD
TYFPcTd7RAS4tg/M390RTbSPlMQJ/duVTAPiqXIDT2GKnj4hyKTe2AcUhSjN
FWawy14IQGvFJquiaHijBzIRq1HL/FUdM8g5H6YqsOZX45QOUMrJT6dOry17
KXCcFZ/Haa5eL/rCAyy0narg4qbBM3N6rV5psdgd1Clg0KQEve0/op1Y7gFg
zBdUxJ1g3VkEakOIqeDCcOYEwQjfyGMRAaSot6AU6KAZ8ll63030nwGrrytd
Q4/S9IUF/W/hqLG+clyNS+N6e8Po6VTfA4wZX7Dok7zgsPZlSIazHx0AgWNt
AIAOYUeHgJ3x0ipyVbc2jfVsNPQAwuBV8CToFeFDf1RM74OyW71PASYkbP8l
PaytmfgGjwe9FafWR8P9Gl6BPWmSZl854Z8WNnh6Oj/9lzSyUoN2JgQ4u+1S
A1WLFXRgK1+EIf7AKiIj28bmLWDe5OmPbXjaowNuuE3QxygK6r6JzP0M0+bg
gc200VWUccf1pSfL4CWzgF2Z6SCq8aE29v0kpj1A5VE1kVIq1MlUI7tAw1n0
E3lrOiqZrIg2V+UYI2FAlnGdNM4nFydgPFQ7ClIaBaR5Ts1UPSpM2IMOSukQ
CmyMTwdEzou3l+M/GcNoA/8M05C/GaKbHxGFHXGo6td3i4MEv7fJGqPYWR6e
Wy1Cs8pugRR8MbeC6t30LewN0EyY6ByyI9NpElSfVcebR+TWwaWVfJ5TyPW7
ylgR5FShf0wTXeCYrFPlA4jeRizPpuY6oCykoIyWcVkKqkGfu3qxSVk1ZYOk
DztHqhzz9ToWvOPpADMxBkd3k3Ky3lrMtAVzedGC3MN9D07O4dJ0uspAoCYO
4h4QkJIjy6N+UGa8AX1Hm5a5MtyXmY9cjY0uMSU8xIYndujrRp5z3tWxWYvS
oxPeQ+tIrS1jvxJ5v40e7AicAxHIRjpgMgrLcL6R7nmb6FyFGxBqDKCMgRFh
73Lqj+YrVQeLdYhHSaMqklS/YXveR6NIQbf0M1snR619S6Rif/N4jdumcX5p
APFpZTKIS0uM1hYmInFmVr+IT39JRYuRbZAiFOxyVG1ummbHgpnu9isKhbgZ
7D29AQastzjDoTbNek4coN7DpVovPhFDFDyK2tGskpY/2E/tgl8WfOB48Dfi
VQOBHUSn/FSP0yAKdzalL1rYXTscBzpa1/PSy+cEEU5+eeXOygSmiT5cjRrg
eUR4QOrInZXRMJMORobAfkaGqpuIXY7bZn68odlX+IpeqIpcbvDgunXM2Y13
VKSHcoceBjJmn1N3hy5vRHHJqegG/hb/ah3rqSYYSHMs7pHoQZPPef5By6EC
ByovUYZX1HDo5ABPq80oFicp27Job/ZxCZmkcZAcb1auDH2u0dEWltsnMluR
M/9HsDkv6JC9Z0v1vbYdw181qtyVdLONy5Sej6VT/S+/KTSq4TNzbz54tfSg
FafVyiUj5UnXGk3lRA6LXbv6xBvFcgRCcxX7AOFdMeHAK08bEi+iCNQtm+xs
FbZwPS1/WWo2uuR9wRHdmf298EiHvI3AWCNiPZhhtZG2gnQ4rub8ONFHmCxY
At880UBx7SpRVLm3EuC/4IGLNSbYdgobnlyJoNu2uRMZRPcfJTt3pUbW1tyR
8WMq3iHihegZLbN4/IgtuVABwsU/nG4BV9EuWjmxOfYE+Zm/hvtBT54bty+I
HFNX/R08EMBYlgNPnNZET6+aSKOPv6sawZetWwvnsirso/uqJkKw0OGez/Ha
2dBpWNFh7XLDX2L8bXNNaRfxZO66h55awM2QVPkg7AFB4lhNPAX6/p0clMEm
sQRdBkTe22dNqs8Zj2v6nAT3E/4ERfo5jyEK37yZg9If24PaEYOMF0yBzn3F
0jolrGmX+YaHnNIr7aJsblFyy1yNAOiBPW32TJe4b9mcPPDUwnCKfV5Rk39n
M7mJhb+B++X7Qta6qwYv44fCEckgFhcGe8xs3W7TrqDRsn9d3c1helQiLzdt
3W08VhnOu+aGi/7QRSAT2zv77JHNzojqRWKL7TGLpZfUJfgCknTuM5EH6HKu
CEGccIWdR5iX7awf97Q/uRhnkPu2g7i7HMEi0gMLpDfyb3AIUobHh+RZe2bJ
BU4wmTSdtdV5jbATjLqh7SjocGVe8HsD57/mZBIR9DhT70Lk4SV0xYW0jeP9
aFFKEEIefO8QUAsAbjtSCuMTCZXH8k+E9qxRpk7wKd1MMUnjNPggbXq7jpJf
uVpDmZsErn38xTSqulqhagW15wlm4ZRnBxy97t+tr78hdw6lGqPlnsNPVLmC
AJMCGiQ1WWhu+CH3c9QohKKINY+9NPrKmyfmuQcA+TAflfHvnczrWXtenEht
QgesgMtwGWcqW5E7Rewb1xCt+jkaKe+4XbuoBBkGvHR0C3SVbbaUZjz90ncw
BG06OSKytU8vOB6goEtzCpwUdTswKQ6wwtCMVa5XTLx2VUyEw0E86fNA7sBU
hu9hZgZuSbhLIUqe965PUOfDGK59wwvM2Xaz/HPRphkn0D55qzxzqdd9ITVy
EHUX4MUP8WqdQ9zAiY43SL1lNtIGpDRBQLMbbFJw167BogJyr65Z/AKakqU8
qAcp2H3KTrkqkcGzSYxNCY1OK/ZMqpWx++H9hoOCa0MguNHnPO5AolkQlFpj
3K/cgNVmaQxORTQTcPxZ99WXMzQ27oIE2s7tGgZ/9CSDncHSYGUr3PzEn8qX
N4TPKnfpE7uyhlC+e3fYKUSWyyVX6lzxSKtjzfyZ0IGCTxY+gA9DDIKVpyvG
Juf0PDt8QcHcsBs+k401xzBL+glBM5AVSJIPwhYk6MfmqGaeTE9+49ncjRL2
fgrX/g4gwZm9+Cl2AQdYKmOhhN5iCpMqdfNJmcRsBzTK+II+aPPEoZciLfpt
GwBp0WQ1GqTQKUFnBKs1YgwmAvtN3P12DVpOUrmdEZNrlSc/zuiUtgWP5ZZJ
IXDj95yUjyxaSIwnAA6WktbZe9wplQ/TBX8LNZOmqoXFwqYUDTOLMT4OIna5
cu1JoGegoxzxL5M6LujH5m/qyfwGW+D32GF3bez5TypZCnkLknAAHh6V3EAb
sU5+LXodKrl8546fGyEMWD7Zy/s6TIbmnwJ9bzcf+YprQtREYemX8v+zQbc4
7q8eIyJilKjNXupPuzRTgvE9LeY3megmeXqlQjfOPVKxpGMeHSJ3Rd+wPC01
kfyvC9BrbpJr09PLtR+7Wm6allktrIORzLIaSTArTgwdJkPZ9UIwIeBinO8W
QE1P9ySAxVxOD5Su1hyauNHVvDgDkWkv+1HzuRgAjwDK5WI4k3ko2tMbioA7
bQ4ee/lqm0h/pPZ/PeTRpYX6H2TVEPvpaEeuxqxr5ASeAsMcsWSh++s2zKUW
rXwaLrgdg6JKPfR81he9jborBj3bFIhtgQE7j6N0iN0+yV7b0PCXal4aFuJB
LdwhVokNJods4+nUYz9YeUs4Lxp0xnN4qECoSFnukSW9E4rc6mV+JL0bsRto
sAQxLWrGNMjxxTtrWaoqzyDs18YIV4Y8ItVWCdkdUyeBdWiEFk+H4tK2tu3K
sP4YDGgrCG/9aKJhMVUFeI2GWUUa4gZLE6J0k/6LPxGA0GX6hSx5rVUGOND1
pLT/4O8wG7h+K8agLMl+19iH1xfjwxf2DOp/HNa1laW1+Bx3JHPcEDntmshl
dUGzuEAvn8YitQPlZYDUmtiCxX23wqcRZHmhpzrLO5NZU7PG7jReE+l+xN6j
eqcdCctiVfihOiJHJHCkmHmgrUz2+0ZgeUZTqemT3M6nZdwXHMawHoq8qMTK
Aj9f1ZFZrukyJNGQVoVNGIOwaCrXYvEsl6Voewa8roGWv4ycea/lBRhVfUca
ddgG7y8PBSAnSUQFnNaD/tzwONi+jaqwS6hT5N6miHNdGwJqK2pilkYQt09g
WRfXa0QxBp00fQNoo8LvZEpUYyl0ebY0+DSXcN13nvYXdP6vUB++BEx2GO6B
X+ZJuU175IJ+2iW10MmMKBma1iupqMXYLLnXu2GJuY8CDlf8NZCDoCj/ScPw
0nGl3pa8ndd7BOslnAIg19qa8Hk9Bg2C0rhKoprN1W3qImmJtbijsbkuJDXC
AH3tP91Na7JU2dIaYzfa6TF5Nk2g+rivGSfUYSqd8aneyzFelyFy8vxAdEdX
JLPsuXSDnlZk3bVr6gKV4xAevFELW/opgAH0JKZ0DEUQDo0MDYnQIqqCVsAj
IrO5Xv7QOIwnzFhsaWWI4ltf654GmUYdJouy0LdS6LkjiP2Aek5lbyy2Zuhg
UwViJ6Nuz8UA127xAGJKYtT8qiU6GhuB72lWS/kLRTLimCjJiuuO3iXzpWc1
3LLLKs2DhEmAXJD+dSEW0bCbeZqGVpizhskzkk5l+qPHapmZx4ieXffA4R+A
Xd6nnvoQegLpUmtk2Ry3qDaK1nKWlJRTcDd/GuZ/YiwWVBCpCAVXjcNEhkwb
y4BBxotvu5mO2pZRyoYQ4qzOWGrV87t5iAokgf8Yj+9H1f0K5gTs4affAlTt
o5at8Lo+LGnoZCFOKijSW2XgZ/I1t2zpYhKHCH8oXSOuHHgUn0ghrudQMkPQ
SADn0CG0AcQbeR4Oo6FQindBcGB8I11Mds9Pho2r0DGiu2HEABlQaPkZBC9u
1sXATc21MJIj2XS3Icvt1teYY4iZcYr554eMiaGUQgGsc7H3J0W6l3I/O+Fh
48UL9+7X1RpRcdACsQVxU5VzlmgT+paGhifwE7GodWuV8Agr4mJ+uR0VaFRv
Mk7mHgHbVLoZrCH+pgF3nv+OyU6A2cmyeYag/LR4joJdEwiMdxAtLfCE4e97
Sgn/98gvJHEqhB/zagvm0xIDv/5CYUovZYm7wrxUhL+r1pJY2oCZvxNDgZ9O
NzZ0Q4RxDnoAqWDpiP5psz+I/vmjB0Ws6eFlXN5f3Ao3pGhBFDFzVwT5JU1K
L8K7zI3gJC2AkLSAVZPQbJvXl8nzPSA3AbXQY5DEmsvlKEO0MEKyaLwP18QY
o3F7BGnQKnU4LPQgS1EqKiadyb8aEHsoXwf4FS+iCQwrjDF8WS8c/gvbkK6K
n/bOp4oKhh0jR4QgNQxmXtuMxPc84I1tfJKRpcgZWcg3ePFACokorlaoTozr
gkapuWtjqCCZ6wvUEYEO5I1BBFDJJendToiiUaAyxt123G4cWkkbir1+09fs
i/TCxwgPxDe1Dq8Qe9PGzn8x/MqqVz+IdfSNAYzkPKgV19SgLo2pZH+VwELD
x9UYunlVdWGOgz1wSltdUXVro39Be03+QSohF3P3DR+dp2QDim0k2rKtiioe
B4O36/hq2oGoR9L7aNJM1xPxWFLs/DNvvvWjgTeZegT5AO7X9wJ1HJMDVyT9
7fyrdIyuqynyXBHZlsLweMKDb2kyJaIRqNNNhFLFpx79QIcW7MnXoDy53ni7
4/rigmgBY2cuvQ5GEW1Y36al3rYhgbXq7oKRB6FGbXuQWHFM5T1vmbDSa5Li
wtLKNAkmB2Gco21Y8F5v3UXXGTiCtVAWnLjhUPP0dbRa4JW8jMMg5r/3d6bj
HxgAfiElPzd622RzLovnyCR7N03lUJna76DKfZ7qr9rIBNC5zK3yR59tL7Ho
AmcfRAfMmHay9FXZTtsr0o9Yidz2ovUkee+Q0AK3FVgsSbonQOL+g8ekAhWu
YV2Tn1D3nvbpm25MEboiEqw8igOX3BbGq5m1tCdQUYkTmDP2SfTuouVPyZ2T
ZGPnZJbR3LwlrXK/p/NKgvIj4VzjvL/Dh5vjscJ6WMCFYbA5/HRyIqIcXaiZ
qagNhb7My782rvNZEyqGcU2ACUAY5q5/iUZesuWt3d2Ae88CcIVbjT5Gh4hJ
TFU7WdFQkt9rsIYMt+RkLJ0YNkMnSRsjzlehVccEBLGkGcYkYOyeycRfMOEL
3UgzS5PJknn3YCLNERu4kcPsKB9jGnfS+7E4KQFCAFQ8Aw0WVMguxwpK+I9h
iwEi+7LZIOl/GUKqSwqlos9QZvHbWNCdDANBnnPiC8COH7w9XFWtqilTAVV2
/OyaeHCTrv+ujjRtWuiFoKQJsOWHGTRoqsDvYbhOCm1SZM/0uBu2bQdvxNH1
4ReQ8j2bgFF7QTHy+5CLYqwTOuCRdNYJw4l8SYYlABfjSO1qhXSYkTAD4sm6
g9ID/c91tJ/0cK3j+DKnCVyQd5qkxvtYUhod5jdYoOHgkzWLT9V71Qmg1Nr6
3idEx3OFUarBzs5MTH46cVuTtwqMmgIZQBIl7MZezXGVXlTGWU16rILiH7Sf
dsOQ7KA9+W9WJpx4Focp6ZyMlHXd6ox//0eprDrjKcaqE6CH2GBszlsvLOny
peSA/gj/mfXkvgZQnHpDwgjwiQ0c9IB60PU28nQStZLfVQUjQfJcEwBYnf9T
bTj0uEVSMR321HXVzqsIqSVAcYtjXxNC34fCFJRF+WwXfkHayPupjysd5kfa
TBMc40+KnfUAxHSvy9RDVh6M8PkiA+x5a1yhi005SpfFxzlztYio7mxwao7f
AeL8vyqRTLAzTskXG2dQKKZV3XQkLdz07Mc2R8sCIu1sRFKJRTcQxtsi/sfI
Hw3QRqaGjTVSidqS81cU9b6y5UNxSrqFSRmPeNs3Sxu6jipSnL4Js0i3AEnK
iVaCJSrBUnSluRDQ82Rh5VZBP7HigB3HWd4YfHF+nEENtycQlR+/wGAYs/Ue
5L+VFhZafngwgqF0VtXa9XYDQde6E1W9JlG8bpDr8HIxZZP4Czw+ch3uns0M
0MBYIKAmok5WGdnPfbA0akPy6Ewy9CEvU6gGQjEXCFWVK+irI+abB3QOwVhp
W3yqj18Y76vtZWwl6I80U20JDPDYK5LTO+NH5AggWhzNQfwtXwBHqCvhNi4X
Z4urECsZOrwvddBtWB3r4yxeWr0TH/rriAj50ldPwrwqu8WF7XnfEYp8iocd
BT7y1mUZbDoMsxprIUs1MmiLTVl2W/u75O2F8MHpmyfl5+7zsKUY3gxN8gzY
V3z0jwoZHVeRXI2D8uNvshJqEkw+1VUwsxMFi5sL6TrEJQ6hrt/OOdXB/kLd
wnlH4XQ7BKGI65xmLncLUxORA/vJRHCR0F8c3LeEHBpk6IFCco9cIij/UVXS
nJQmzxY+6DMXTl6LtsH+TVot0ZajzfwoWwZsZSshas/bjUbaKiLmPeG1Buxm
gtYZzn/NWFd5frOA6a7kI+jvfm/GRYy142Pi7eJreshI0rQ88qaBcYK0y4Le
AiVzjJJofCjBJb4lE5GuahTiIFQ5LyTvoTCYJ8fp5dNh4xrI74jSqpRKzh5p
kSBwauNegdM4bmbnwMCFijo/JW45Yrj4bqP5ysY6ouuN6z4Efpj3efIpWNdG
THwNuflCjv3B6Fn2KfPHwOTwJONWUc3e6nNDGJilT9xUaqz1lJ42edkKvJOF
Alk2PXsgpu5+8gCNlTKJEqVmaD+kFAaTY/EIaYxp6GoD9QZILKFtWPKfTdI+
Q+0G0vsIx6h2fMsI5K6u4lpEZ9kfhjng0PRy3o6OaqgJQkU3Mf3kTdLXAo/8
hTIyWV44uXvyn81XjQ7oQINUGSHYqRmmVMX/7IZXNfS37keb5/i2Z3lqG1li
gBtDp8PAYweoe4MLmsIiCVuOoD6lhIoM2G3Aes/6oZnlTRQ8pvebYy0dR+lz
qUFPqrUU75/IPdYWI884FpTH9dlyujhAH49+c1t116pOPda4mCyQk86a/p6L
YThfNvLKHgR6EeFJKm9IrsaM6tZq2qWXvxDf06YFE4QOdM/U+2w6IN+EE2li
zdcUOOOPE9dJGSUThNaaPvRCFBioxVWRpKhKxDyCkKzQOvEu1jnSDAiB/S+T
zFlu4LIJmM94eCjdaLnwqdnzt6j9ZTPQu/wxwCiENzqF3wLVfHnNQvGYUZhH
C6HX44Db+JGb6su7WFztlGEpatH/RBAAArT4I/bBmk7keAveTNzmj8KGbbW+
ZA/ycPti252X26/JiFFZPoOxrTMlgMFmS+3Ca6FUOjuY0jGHM10nII7xjSbk
6ZSyD2+wZoEKUHLOVJfE40aBdbyhRkhsR+EfefXmIzuamtB8IEJlHUk7ddno
X6hu8JuS0haWVwFeEyG8774K7naRYdbTEiYPRWZl3HQ4cbHgzVqeT56AqN4c
BYK6tddzSoKPLoB63Z2JxKg08gVkihDuMErJ5mwZ8YltRw3K88hQZKlm5MXL
UdcqJSmiMnx4N4sCN1AsiJ7wXAamxJuJgENapEG05x6oWha1CMptE+/w9tJs
fet2TKeCXWYLqHXZz3cvWxmRxUnGbPt/ITqQCZwpHCCImid1z3n9qRAgyCdB
948Ml+tOWNWtFB4UWuJD6wvGoOJ+7+By5UiHv8m61M4VxZj10svIdAlhbXE7
NHbE4pjYEV3hFjD+Ge2M+oNTPQEXvEDlYH+fZJ3CvsptTqxbLQCHGuAnNonf
MAWFBp4PMI8wYNMBboioJbDjg6ooC0xmuIl7KviX7FXURnivRzP3DAXiP0OP
zFNHH9kdoHZmxbakP1vGR2JnfFtJrWAR2crDUGfKFnpRFL9L1djzsqQdbw2X
CtBscPNUXRWskozXqALlzsHUKO86Pw5YXcswCqtzjEZ4lSSv/jIcdO8qlNCD
I53NDUvz/UZdYT825o+pg5RfRpPjKmVExGNLjdhx/HKdmx5XpWBUbQ+WnmWO
5f/MAP3zwVnokuUmfzBUAqzxVEslL7kjLkHuY3lfUoCVKbmJs4Fu38Qas8oa
2hXwRkvdASeosiDJKqu2p0N4c1AaK5oMFxOMGKL2kjX7l737SQj5yGWOFoip
blew11F9G+7HLRXuplv2xZMhuNnEqZOuClTsQVqGq7Njrmo/9Iagp4O8BaPo
ti/4c0ceJ3JgaIrn48kFmM2AQu4IEIIJVI8ucaBEdjHyiSHTFYI25euH8Ag1
2iwTVo+zM/i5KGqJtm+tUnydXc3nGcGSbP6oW36d6ndWZ91pJ5kpXbASME/d
lqb0iET2KhYG3Ma19P058QIfjBHKCk547LpcWafJxZ7zwRKgw7x4NZNz3LC8
R9FiL1h5PCEmOZl9nJTMPEKAMUzoVC+x8zQ1mWtHKbKGApDbqaoGvt2C1As8
RJjatwPzfbSW58H/C5Ax827x9CosFq8bpcMVkpb4aiJd9miikvC7ZiCGmYyE
dMse0OfGy5xZ46sBRmKB8Nk6+Eg64DGjALWGKeWZtV3nLxNsmnm95BJU5kKt
yF8zquOo/ZJqM0lWdNMsEAy88UnvCW0Jbt++IoZPkA1oA2NLrVq5Yku3+VAO
qs/YAXqnLZf17OWTmuBN08HkNWBLgyCdo522OR88Obtn0YqdAxmCO1mDcZFU
Ps8k1BT6spkdIWGIpjC3OzfuTrR6cUYgleTWXxa3sVuyQPnB4CQcEFy6sbos
U2b8bocuBXC1iePHx4/SEwWY4vaJ5L6/W9jQe/+pgkBf9vJFPEESrdbqsNRE
CkXiTQPXMKbBeEVJ/iq+TbN4Wj0PuWJEYy2uckbFB64tB4cT1RikDSMBKi3p
SOQNPMdLgurGTg6ZdY6lxNLbiFYopzaiOxOsS+kPj3PRm4EbQ2XI0FaUGrHf
N3KFinQ+/bEaQp3F9LP93OkbDa41qjuK+vyJxfZjllpmQywj2Sf5odmzZuf1
IAFKyQq4mjGNnKX+Bh/+AZXD0CCPxxDTR3WdRZC88qYgozk3fc/C76pdeSjj
pCQsy3KBsOXCX9KmFLCUUnKLBSlSUs4hLEALNN8lmRuUvoBEiLi4923A2Axe
rGQAViRQ80LKy63i79+Vzq5PpoJzlfQbcSMOKPyshcllOP6l1R+XHvlYDdz3
BbbpG0/RvM3gT2o2eUKqQzOvEasS4QSgqO02xcEFDZJ2YEB3Sv5W0TaV/62U
qtio+BrxOLnXYS6ITq+2ULxi3Q1Syz7otR6kTrhHVRrJLsdOL/1pZgT/kJIn
YIa8x5+Q+e68eUqr73Jt1F4V0IUOsqgq0rOyzI+4nxQHIsmqHN4Y63uF9MN6
YwTafWj5qchARAreDYV/Dso+wx4xyr5Jo2OlmJdz6k9xKnoNOwXr5xmmMfRT
9Tm1jMETOrVOEHWYnkk9mxp9VwHtdvh6vGG8w2aZLaqxGlZjOL5Bf4ZF9CwE
6o1xecx2sRbX303eVutXusxDVchOGyGqgy/AGg2Ior7glWrZb2NPqX7iZAQ9
SLD5HYD9PV/r7m8Wva/mUJviNOXRLxxBOyh1o5WAgVHkAQs9PN8nycyPlvwY
QcM4J1FUmEtjsd7FJWcO/qCjvIR8Ww2UuUxhFUFaZxrTXise6I5DGjlZLoUz
y0xjmLZ8XHGPwIU39EQZlq71peQGJWlnBIuCQf38pE5RIRxRWlAXogUXDEJg
3fSRgxXIfo+uS1LhUJ7H1AE9kw5EcON/7fO2B18JvLeNQdP1v8SuT09fk4rh
w8T+s13EwMkU+2O56a+AQUoVV/gqq2/CCoCtoXM9dXp/BDwyp+bGjS549+DX
waEdTYP728i46pzwgKiGNSf5PlVL929MRilqfaH+7mXXrG5OT0DCdDZvtRNP
fY+o/wubqkHNZOv99WRepT+5hnIWCBUXWaziJ7k5LOAzONauvoYj7ADYHGvr
dwTRWyWYg0tUpN9W3QHk4J6BISwgai5+2v0QrEWOqLsoUy9bImB8fAvc9/Rm
LZHnTCLxWexfNahoOk3rbaZ44AzitEbV/Ou9BHqheTWPfG66yQk5LTwXvSwx
5hgZ6+lS7BCy/dsQHFxLAxEaK9yfqJUBaMaXBsJA7rHw++I62g4aL3cbHVZQ
LBwHx6i+GHhKQkVHHe2XWNnbHsOsGRIHE4KHjOPfZTdiqfhOU19tadEvRVFN
JZJcgR2pAHbB4V+EdlHl4vo/0nRoze20aydBJTj47Egf7+n8pj72OZ9UwBwX
zuHMfWDkgCw959D2qG6Rsncm1W6KqjGvPdJcrv9j3mEWI5eFQ6W2mAxMTDjc
+uVja8NMAWGOQovNEqEOU+mOpjGgnQK2KnvFVUkK2JxoF8bAwTxQtW6BHunJ
zjzSEdTLK67kaZbifPAmaFC2wJnyl3V1sqyCwCJYHuI+sFrvWcLT9nagveD4
9vr3pR88ORkhmTJhxlhFytpggN6hp+GWcofARd6tRgJ13vmbxxsFt0wVrbMM
o/ocoa+3JyUOIA/Ly0j0ATJGZE1z9W7SmMWCuXhcyuSBjMbHkXUTcD6GGtMS
rJYH/qn0wyKePsPn8ilNe5IQGw2WcmdpmIHEGY/7TxajULyVqOdE+HV5yeT8
6c6ZdL65iFLZnM0phTmVBPaobpvMv/WmSGHd078vK4i0G10X5dDMHC+QWKRx
SMJ1g7LAYKYOB5+2rUxCsfEOPII/p27ZVcGdTxSmrrNKfiFkGEiuo2fnnB1U
C/SgrjNDpzYrygc+x/KFfCP8FoYzpv2FBLz0HDyH1xuinY+ES3j6s1t2YxmY
uYxDMmFXF9N9B8K+lG/wk49wdAM4/164+5+GRqfVTxE2dnVlqjmoE9JqIZ2o
wmO1DuiIxCCs2tLLUUlb/8VyuXakNG8m5c+vs8FInEdT8TaqC5SLvfeh9IHp
S1rJpQc8eXE0gdQPNksujkKwK7XSf8nzyOBx0iCOOApceJSAubkpC6L/fPsu
k1MhCUlmboJrXRSccA3Doj1NfivfUB9pmG1GnJmfRdew4PpAsM7FOOokvNLJ
W0YOCvyFHaz8ZVXTHyGIbcDPbom66QPoBvIuJClIqyWmggM4eLR9a8Y4v5Y7
g+eXOzjI8XTd2NK4VpxzE0xcNKBRCZMJ0FbPlL/R4iMIYmAVF22m9vI4n5y5
q5QZ4CXwt2IcceOqcQHK13LgrW3ZqR5viYoXWL/sFkznT5vV7jZUD8F83Tmc
kQqPyJ0JVNdfZ5NI2i74aV+bvMHNng4bb5n3Hf+1KBXRgEfcX0X0raKjWcDx
ntvsBff5rmlmWBRn1m6sNOFLp9tqBii7IWd+/vemHHsjvujLuN2LV5ccAldP
oGlVQOn1uPJcjr1oNFPzpdpkZxLUeatAJR12beM/rWXAdCqrGaFe2sWzlUh1
HqdV3uhcyYWNuIo9EThlY2MiJRcMo3tareUa12BDqGbmQ+93Bz0bcCpiBtJK
FfbEktWc+Mo+KWFdpXW6+I4b1c5bU6lvGAs8yij0YOkqvOsyDfR/odwRwZNF
YP3la8OLnZDhbRuRmqjwZxIl7rNOAPshjH9Bqdkp6JeferGDeWxEpJQCefRz
G3zYbE1qZJd1rQxuUBxEdqDnS7p+ki5dES0gE0zSdRwKrvnKHw/b35NCE/yY
XVnJaQpcT+wOCmGaI5FpU1wZTlTSDb4LcI8pA9HcyKAIERHbSg/O33jJmnA0
wZEt2S6IOCK+P5D3EF+M8kwapEX1HJSpfsoWgRmkqcRJe8K0k+0AP4JdR2sD
0IR56wMVzeYGgzO6aG242s6+A1CV0Cw5Wcfl2p0yJFaT6nYqV4VY6qWRQRrD
Da7Bp2p/TA3ByvYuJEONZyiagO1rPA+3xtuvjiaoDIff/WOzzt3V2yIKrU8N
HgbMuyiMjUfjQsFWIVz/iqLo14jm6a/p4yEo//SoBDYboZiXrrlUxg+cGjqT
vx2n9/f5uXwHc3bB9XVUDdEEn8mR+nVqzgbWFIbHmomv9CEESsChWUQicW0c
6JVgf44dPJ1TwqMTUGqlw9zeZtxjAXe3iJ3EQili3PAq32X/qnnNsuO7bnZ5
zWcwRHHMATJPGR0YLRXGqkrBOq9CsD3wGqRKtL0pyNekKIDX/JE5fKeZWvMs
wknSOCtBxrE97eSkMjhGfyhTWQWU5MoNAZBF1cXpF3P7GlTDWn+GjhIIFL64
t03rk8Nv+Ak+yEr8pjZF52sQZ/ywuvHubeuTJeyUEsYgcJAC1EEYUHR1NsI3
BgfWt9ga88ZzE+P4RK1j7GlfSO9JgsryDn3z2zkbJehQqWt7Vo4gg81hBOMZ
2LloKFx3EXwc9RPE9NS7UVI1hLx0SNnilNqfd+RBIwVpq8K4AOT347eMjKC6
Jp/0EK+enAeFmrUGRKWPeZl1vXOvTKIMRShsPEYCkuESgxhqjZDPWpLTkF5d
cPV1RRKojKXTCjw1h3xiXgjun1j1jHmyDIYZ+fNZvFxDThCWWjY7hoU6DRPy
8mWOheINGCYw/tg0dB5EygZw7NlLMXMlVfWnVw/2x0qM49CjGp9L/Jl0Bfmn
Y+0LMQan7fHkGzwHZ++HPA0AUas9vfie5ODmqnnGoeYvyCLYihc9R/zQr9Vu
G3Zau0vZ9TEtk9CsZzGTaVZ7Wbw4kndkqZNq2WmTP9STchmVyI4FhuLrxnKG
N/ZUi3HC4imN1HDPexxi85tPK9fo9mcG8VYXFW1GyE+Y6q8dPaWgCnTzy7BI
V3oXvtjztEQpNF3twM9RF/wZo+AAQpqhTOh3H9f4bOmvzWHoJZnv4CaCqhIz
QDyEbCi5ghSXac7vLUtMP92S/ksyYKmNRiLnii/b0ks0jrvcu3h70vCHLn4/
MqTp3AXXwew+1+9AnsAGAS4SHWMYFvo9TWR0D6qXggz/C9hvkmeAq68cyPaY
ZxQqk2EkwoeJbPfCSeob4eoo3zhKFho34sOCWHGAXWwhLm+jhqtuSgzMo4r8
BHMWxKBMh97/OYDSMsMn9LyhvyctoibycjhIji8wEBtWIOYbzkh7RwEveI1K
Hh09JXKDZoXtXS0ROIUAjdtocjffaRqJV1jm8kXE7Qu9FEf15AGOvdI6bevA
uEnvt4d6MGaQXSTa+keuN9M6HwjFqdoDdDPT7C64265zUHKsGP8EeDg2iMOR
wx16vdkbfXbLRH+VKHYBve/M/mPhVWrXAjYl+Xhi2DoOY9khQRxaQ9rbdVLH
sBPnNsDQ0RAlaJ1unVarL9CFTgnndZ5xj7gpOsPeHdBgkTKcS0gf8v0Tbagm
YTUgxWupuNK2lVyBnXBe8EgGeYcmaA+5DhgtNLQYdnfA63W1pTjU5sjF1Nm3
9MeUvdjfk2REQUAcwb0PokKERi7J/+ILjMRnRtzYanVlx/K9nmzpyRJzSXBV
bkAMEvfRyd2apcrF89N+hTW3xRFoCPAnqQsa5plLkGEmCMK6GDGHSbsn5uWo
khdbk4TdsUfXerhmZfyHRBMaX1EjZ3VMqD9JJPltwYx6qlGxMt2T0s2l+YhE
KC77gSas0BdLzuSMGMOMzQA79UfKs4QXcFF1AKq98tae9oEehbO6ut0QXPpv
JcQyIOPXqalKuuT/266HJ0YFUXW00U/Q3uPdhf5qRxNeIBJxLaglN1ragRrY
iWjPBbneX6T5qMpGYMjtyIlYGrddZS7RBRM9WAJuT5nB6Dra9OLU1EUXVeFL
VRsRPVZ2cMjpbsUXNn71Rnm4mCw98kr9AxIguM/rCqtJHu30e9ei1Seanb6n
K1TGe11F1cqWjvsyFZyKQp2W7XflxBJ+GsI1ec1KET3FK9FeqtHCakvhawit
n/d3z15lzcMafAn2ulA4ZPoYqxlQUSzRFEHn1/vk+aR5PYC7n7gAr7wR5ino
UfXg5iqC+TOHghf+ULFhqEjxdUC1gKAdKQvmszzj8E948C6Xbp6GzKNL0I7W
xWN+agRgVxSk0N1F0cp86HORHI/EoeU7x/JUlA5Ey7JzDQobAZebjqe/kuZY
NCPFtfBZWppqbrQ5pBGRYlr8ZR3fgTqqFBjTuuiQapgCIzH1zUVwaUZfrBt5
Wt+FLa/bN2wIhShj2sghSwtDBAApaDwVkqeJnX+iT9OqbWlu3eyA77JYvMva
WGzuxu6azJwSi4f74VIsgxP45ZdqjqQP248TqeSD0Qmhq9ZtA97qxs4xRFy3
W60reM+TxvevLd1oTEnJfOuJHmm65sMswSiu2j9K+xCHNaf53ry7imEVeAN8
mb56qsThn8VEU3eiExwASw9bD7elJVgP4LSGTmuOn4nX6W7McM0zI6smEBWT
r9mmaBs7v49iYqg/ANGkzxb/Z1gV7jLSlMO78FtNeFEdnOJB1PmQc5nV3NvZ
vGtwBMyPwtA200x5FyNqSdkNHlEf8hcEPZWaptwPM8NEyvMhiXwYSxiCb9Ua
+T2YcDloIOKbFmudg3rpYjsXrqvQ7THLsn1uL1RCmaqhCimlIyvvxo3Rta9h
tr09M4q91BWX7sOtd2xYK3bHUiXHoWbTahVjxC4vrjLLMhL4KGxzGdVpCyT+
M/uKObwOYSjyb+4aWrDRz9aecTJ06r0NCP/c2QjUDlEucaluOnRCP0vQ+Hv3
57IZQBa3BDwx183fSkrw9piKchm17Ne+A337rL1DZbB3WPns6FdO2MXeHGpK
BPA+VS4Jmd/A7294YtJoip+XJyhudW0THY2V9q8vvIkxE3viDeQZuBlAb6PM
mtCJkiLuUJJSbHrl4VByqL+tArveN6fvkGKcw8HCvfHbXBebr8mkWWdeROwR
1mEIepI0LrHUQc5mF47UCnqfZR4GcLxPmowaMGOz5EIL/WwSFDKbjglWpdjq
csXDznn0VbJm+IZA6n5clTshHfMHNvPbBsno4NbYRSwZeqB7CrGPJNDR8xWN
lWYypNO8jF7YW0a4tT35gMkmNkAzOrcK1uZlpw2bdkt1P+4dkp17fYcrYgsj
jc7TpXvgEWaa4lCXPziZipteBdRqTIDcmz97VjPhPLV6i6hDYJlELglbfkUj
36wlqXF0O21CSovn7UbvONaADCXsY0K82TWSwYuzgYvOcdchojNrBbv7mTEn
Zfc7gM6/GjSntgrKXZ1tnrD/fgp8/KGuyyPxqa0SDjWgRwIWMJDW+6b6bKxW
xhbtqS7xlVY1XCFFhpAniJO1pGKnM2wFD3xAoB/EqK+dGk7ujrtRmlH+uaU2
wzRNaKbVEo43F+9rMlqSbUPDY5n2gFcCBCn2zgwmkX5dtL+Hpbo6JtRzr6HA
dUIvBgUePlDeMcHpxO6QaSeCKE6hKWEpHILv+IV5X6te7mEWO3zYimsvh5Kp
XouG836h1kDmQ4SkbCp+kyaEiUJzhg9R+1OD59FkEX2Od95taRnulbHjNVU9
TLsjRaPS4FawBUafUP86LG608Iuzc5yFf3MAu+HWkLckiYL2f9rr/xJq1o7u
PBgg2/As6GW6rc9ZUAHP0eUvLeHrIsnH8KIj+sAdZUAp1WhaeK2FU6McgF8Q
c6ZqgAh93tipVQIohKszkL9E9IWOiquNgHcLvTL+VgybzoygrjOWUQtLKKtv
YyLRKTK8wNKReekyAtua+TtBC6QHxGCNSp5Z978zrobcBLYnNW3cESDdpJDr
hkIXjSycua5XVDfb+eNjujdPz7+L97vwhuV1T2s5NV98TdbxKCfIRE/vvZLQ
tbqUxx6MDUMb9kCPtteGk0xaihRmegNmqyGtlaFQqb7btHTHkhLa2g18ETY4
mN8iAU2TA2AuQIpyKWtGtYm66ImMJPSZIg1O+ijH5SasRAgXjNnlGSeoEzJG
yixhTCb+hkGv72aroqsfFZ4VrDGyuG8mLWoClWoPgB0oiJRhljgLeVzsxwwf
/tQAYRyHB/DRi7u6EFHVZqtlgzFZmxX5cBD6HmA5pY4TsQCe0aotS5YYTh5Q
yjhtVL4nLkoAuo/sRsNWkhwCBGONG9S2lf+Mc8TZA6lvc9Xc+aob0URGlj3k
LMPruz4aMoUDSDO42Ued5Nn2ra0gTwliWkYCVfP7r+jdQD5rD4pV8j5rVqnv
fxL847ySrucidBcix9d5+dlDeyZViKatMAGyz+VD2vgJCqek4e+1XS3ZCt7k
KN/LACaQY2ahfnhz3puSp6uVuZTgFKSKdQb8Xez5AEb1tjsYwDiKcnDMc2VE
kXRp1aJnU8h62LO5GDY7PQipXT5y+ERgt4e+JizDoxkgocbSWivlFW3axLQX
mEIvZutiy0rX/zVgsifs8FAcE19ajUjYo0UvK4Jrw942Rl6O64nZPCq8YJg/
cRbpv8aSxyEQ8ObCNnx0BGYAduvK+f50XGa2SA1s6/ASJS3uiCJOYJOjF3Wj
wlTHxwZmBL2z90HW6NYbA8a26J8XAHGfeOkfTfJVyLbBzV2q6ysXBsieEBUh
K7sDHUW8ZiOvacYo9ivd4d2o37qLq/AwgYSb75cfW3z2kbf4Kb42gLQ7Hd67
KQs2cVyC3I4sL32ki7Wfl8vpPIKBJeq0QQ5TRouoWbCzDiwforDa2tb9qECE
HSOZnsuwAF/zpAtbiKzXOI54Nv4TU31O5R2Xgr/W79Y6ijEPkAqZfFKobpVZ
Fqh62YGc+AW0sJAyWJ2VkOqDa0JGlROY+J+55wRnOmzgUGGvz8KOBmCFY6Uu
yKpv8YXbqbR/i+2bOgBF7usnWk6NOH8pbtq9o1f3klzIFbyDh4BktIG4fI7Q
jev2NWAAmSmW41x24k8ludOgDlPO+70QvgAnQIGS4DrBhQ3sV4wX0LpeexF9
Mbv8n2o9J8wGzdr2MEmDQYlt9OlvHXCxT91smC/ibrM4FlMK9afyka70jyu1
Ud+qaYnKvAjSkYVMjvEQQRML06Jn1Y4REaakEfUT4kSU+03dYMTs6Ju9xtsn
+TgEiZeLoLQi6qS2d+yv74x2B37S+wYx2N6/u1mMCYJNrbuXWQabC1aiICJk
thpN6Q3u6MIRV/q9xFH9LForxxGEBifrIU+OHB6h7CemzM8U3RJc1jJECc02
l6kI2di5r2cn+FcEsE10v/9dvPeO89fJx7jJSfGqnRThK0iE65/qJShTcM/q
RshhGUYY1oJQJOjxcgYMg6pqIZ96AZn6cQNh3g9xbtZZNBks931PilpHplo3
LLqbnuK2taVsE3DukDYnm+4C6F+PwH8NHGSdQPP4HDq1CdVX+zauD8if3JFj
A7upwTSyqVg41a5xj/zdnzaN2ohi+f6g9h5gya+w0JdJEY7nWRqtEo84ASuc
zkEAvUX2PvkJgjukfbsZb9hfi0fqCpI8XtwJOSJzCJfnMo1U34GlcP/1ZQkx
Y+wU/oXQu7P5TzIk9uILa8MtSvzuXv1JN+0ThTtLOXWqPj+vmNIOVLytFFL2
vik7sJph5APe0NQoSwZZOf1puIdWeNjVGW47f86Q7NUwb2rT8NDXZEe54JVj
FJrV7L7yb6D0FDWQZijcfXwJhMImgtF+v8zYWLDsLiq/VVwpMQ0iEERc4olk
l/SPGC3iMljBQwzAT8wDq1aZBYVvdQaNtpKA5VEGix2sDPD58vCWtB0NKcX+
3PlMCQrypjuF5SQUAEPddideWCEcMkRwGeqnfBZcNbVt6e+d9gsqmyFM16bA
g4tYWDodmnVy5nBF8O8U0SUForYKTo3ZsOs6D7kNJSnw2DCjS3fXOeWfcsWz
FBTpt5nqylFWp9VcR7wQo6q8TEdocpaRmzzTokPguho682qlMEsviP1y6uc3
Zr8B3Y7Mk9hJlMYxDkRTjHobG+iFB9UgNQfH4IjByrWIklM7k5oUG8tVSuHm
L/5BZJeWfur582+Gumkz2vRCXfYyHjBEjnFfd07S0AGZ08wAJ7wCFql6WS0W
hI0Vc+R9mc3jRlyhgCCl6+PBbUq/WwymOeu16cD9293AEKouEjBjbfTd5tPU
hGTz2qAqT2qMojUGmn67Wyci2Fy0s502qeJWGZwAa2H9sB/spCFtTrPwiPSB
n8d+Vca+j/eNFxuCsCwyouM+Yc9WjDEQ4W6v6p2WQP42TwVCc+DaFCxIg6ib
u5N87V5WxvX6qtjRtHIKiGRyAL5gCj0bsRlUBB33tB+BsaYFUjYtA9PIrmkx
V2GtrqxmtQ5Pfx5blmZArur7f6Z4y1IHqYs41TDesNiuhO1Z7o2fuwPzJ5lh
LS3T0KpUVb8Tt6s8kRNOAJMB+oMCbmV3JkFVP3R1sicBbykJeHq5+ahyKtV6
dBK39X+64CqW8dAb2CL5aStkespoONsZAplE7/IuiiLM98/guZ222e3+uwN2
lZu1B61Zo7AjrmFcMCrJzBVTEsiJMZUhonLoqQwjixBUvsqpCGnnvLenvxEs
hKOGMG9oNDvAAsTF0yecINUrOnSBxrgUrD7tRxN6Vvz0UsJcO2gpvK3XZ7MT
2w10HZ7rSPFWTHo1XvkCLF4sow6ng3mCdXoLNNwda+/JZdeNjra4VovVp0gj
bee3mgwkwnScpuOzXKB36RRJ27Vid9sygXc9m9kWBhDeOsygobFOP73iB3lZ
AOx1moPUak6k3RmPhqHDKIE2BzQCN/0BJrk9dX29OPOr4/J8bVuCaGQ0HdiB
fVtv9RICZuJciY8ioHcqjh97Hc5ubZvTFIKeYFhWoosSLkfud2q0xR+38/Rb
wCmVEkEMSitiOtT6pZEaYkoYkSxr/j+hMd67oQkK8+KeWeZBfZjTuNgmG94f
iI+NvjGK2kuRV9VXYlnhKb56qkENQhDj1cgx54Nr9ReKQkOJ85ohIKWr/Sy/
QhWwDIWPtzfctIyK9jgZvWoqhfYfKVR2qhZ04myzO94us8TlhWYh5V8MfE//
0n3bsrfZZCsC7jr4xe7BzNxv3Anu9W5+4SYuVKLorEC0sVbaMhxZtG6KCfzf
wD36PW0yAUSBg48ieg4ny7Dm1In/XgR9Ph3tU5423QyQF3usCuG5aJyVfzJC
UTF3BOnkGGEr0+rpsJOJJPd+7jrYQQj62jpwYtNhqbZt1CaaYrgqv/dbBGX4
wlOdbnQdqJiGA1ZKWn145K3qZB+AkPx3UBNNAGkTBJcrBLs5Nqj6kHOlkgIT
qUAxkECfWVIYxhP1FoKF9KwVtKNBuPVlBe4DBendtr2IYsOFRREOGZmjhdYj
8GORB0HYI7RibBdNNaHDIYWz38zhpld0WX8aqrXMeEo25W1pi3xQJbrgI9T8
Yh6y2BZf9r33sy3w5LBtCQfYaoieFLHZ675MRy5+pOoKO0Ls+wbMkxsFe597
dUPO0ZdGDl1Rzj6cvs/UjuyI4auj8LjfApuUmad9v3jD94Z9aUNNbZzfCJ0u
ZHizXOFi1TmQloC38iBnc51+9H0urkNihHNBeKGB5Etd+C1II0z9RludUOE4
W/ePXflJ3rKuk8D/DU8r1zUyT8cwQkUpelkhh32EY16oEE5S6M1CQ3xSrUTN
GZaN5Yfj9tTGIR21pA81n/DZ06H7fxLeIEpgCv6F1kQ075cGtkB56lihMvap
Ry9D0zTdao4vd3E7RBroH9YKQi5Q4DSLyDKC2CRWie1AK1VaxzrXb+1GTgBB
X+XchJ/Q1kWgcewnTN755MyTHdDwOMg+OaCbtmEnZpa0DXuyR/R0FOjTmHKW
ty+wb8C3u2xodEXqPpP3PZKth0GLrHfdhBwwyfvCkwWOJVqO3vryPT7wOMlY
1NO5nRVe5HEmJ19Ijw2Z0vr/QV8gDUFGaVfHgL9EKPXWbZLDYd2PDHkMWq/x
+fBZFUeE8Sby4BOdrdVwIl2QLDfHWBtx3GtqqDIR+ZJGTp19Sem9rr37qIpw
X+CwnOJNTI9nnJzPEmbfK4Pwv6xOBRN9iMPfvURbJr45t03VNI7Zx4ajVZZB
DoqzzNB816e9m2P86M+4WgA2kixEiZBPsVUrcsOnMT+a5d2D9XTK/O76hzAM
M8vK78EpCoquAxw6tERVL7iA2GrCNmqkUJ0exJNx7NlArYaEVC4wmmZUCtuU
fu+Zx/U/O51+QwcgWmFmtFjfhdl/zJO7BNw0heFMwCyniJHlbCzSi7FwSIZz
HVE4cnYq77ZkA0eP6/HnFhpkewLHYUaXJA36D3cq0osM6WJ5S4yvYZ+Y337q
pUw4Z1HIwHYHchZNrYnxSaTcYwacC7af0KV+ndW0Ng9DwiDZXB1I89Jz3Efi
jv/9uUrSegQFsZzYhle/NcRMqac/SKFb+gvAJH7EwSlZdV5+8GAx2PTpJnqM
cxXflH7CK+jxlaD7DvXf9sOZ/zBOGhGnPiVBRgMi+EYKhBdH7rCfTFePdlA9
OmKr9JToSt9z4nC0uRNnKc7Nc5i4wb20HQofbJDMFPiGT/666nrLVeC3SQ59
0nUcnyVNHbU3G+zMHtoUD244EtVRpy+3X6lvtNm/FcaD7SCj/9iPI75ZKuGM
GjH9u35/Hw5N0K4kdEB1al2+dNXt7vEX+00CKch2u04lp48HinW3tUclT52I
fYCo4NsvcV4H4Y1dLtvJhir6YjMdqbn3OK7z3wsgJY0yhaMoW5US1uWEQE00
W67yfmXudNVF0NN46oAR+EG5dfxnGOFwmI4D8G/eKJVA1I+S5hC4LE3bdf34
Z9U3/WZsPa5MnEqz6K6+WbJ3qN98MtUtvtUpwyd+i+zKmOqn0ueXFJ3EvV6D
spoMwqbK5G75iek+tB6KCiPpJhJymGk9LSMoqOb+AEByE4aH3NGtUuVKjH7V
C9SPsELxZ9OP2dfZf1w5WpPDstLpRYRvZtT5MzuRky46YmNIjOwmWPTxTMD8
WZomFsygjO8S3jyzJJHfmDpKblDcxAEk4L3VGI/VvhKAznkUwp7ub7zC7gj+
cl27LyMks3m8qOCjh2jML6PVsM2166/6w9ZY9B60h3zxEaMMvt9TFqKOn1Y4
/AV90QwiUG+/pPHVyrZifIPMX6OUXeQt81hJXD3w9l3+lg1BwcSpjQPOTPdg
z0SZJuSYX5Yy42NbaSM7X5OfFbi6TNh58x0yKL1N383C5s+QL5p5J/ibD/U0
SDMHe3OJ158LRvjD+YcHORFk3eZ2MR2P8FvQs6hil2IFfUWkDx1NhqJeLj/1
kt4TdboRD9iIyU+rMho0ByUyy6Rv9IJHnmW31B9StAUwgxcOX6MKAh1F841/
Zkg/43mbDfPSyMvzFndDdHWoryVDQsUgZqB1yvOsgL1cipAwainqEyAJlmim
bAfRfu65/thZJOdPgHF+QIDy+be1BH59FM1rx8wopT/LGaBO2Q0TS0h8E9X9
wvKcReBpQnEu9jKJIAhRUpx+mEmM3rgzPWo2ikGY1g8ppts2zOhk36SbHbEw
LQ3O3S/UtQUWcmr2Ydgh2EcweEExoE3dpTu6+JfshkOZlKCmrsa4VRBYmAOC
UuAImFfWxKJyyV408nplX830X35tqmDp/UsV7So2HDPgLSINg/aG5RVg2pCN
bVWSXbGxelpyHD5ACFicUoub5tbl6OycTJc8aoHGDNMkOp2Abwtlad4F105/
JpD5Wecotq/HPCiSTxO9CdIiuco2A8nrLgVVOSWdiQeux9iISKPLxNmllZIJ
LOK0yrYPqeQ0bUnv/2gCV+H+pSnHRreFLI/JNM617ss2gGhYRglTzryKZZwY
3pnA5BSwzRIaKjfo1yP82ymA5hXbQKxxgl5uNolqc6Fa+bx2SCDGFmEgQQfv
n5+aiLF6J5orUyijT1KCWY9GPPGte/9/bvtapPO8VeFWqSk6vIKK8ABWapL8
TsBWOnQay/nuXxrolZ51CUI31gDGGXejlxex4i3H6gWURAro4rof3J24DESy
nZqPyH0CfW74GTs5UTP01HXC1d5/CgD5Z2mqJV3eVPtPPt1fZg8qz/i0gZes
IAZZkCV0S4zDBA6l54UP6VvPt8oVvHCrNJjzkxjcODOBeUwuRkmGAlJd2fCe
LXT+XEj/Rzu0ewIdF3s0XkbdfreyIH4e2d3bt5XPIUCJFk/RRBYKhOSin3pF
teazzJQePqjothE0eKbesHJGSKpYCOfoE+ItnqCE3iHJmfqLZHDYWnGXE4zD
/Uv1kmpg+UXmbVRkfoXOOVpA7qbLRMo2nB48TRa24+GgV8mULCbYE+itW7ik
83kDcrwWZI/I/fXOItWVXHljMOKUfKm9alQnlEr6Xq5rpU9QJ0Vd0LMSsdSK
8U6R8ux2etWDsx6B3pL9JME+8631cY8z5KvfZ0SfnmOHQjRTbsKR/GzCCUrX
B2JPLwe72J7ocC8ecQL+tw8cMwdALmtxYlyrbOmWkog5i7To+1BgqEuzz4OG
rudCsJoz/MvvTeTSq3YjEom8sJyPn7nrdyRhB69h+HNoC4kuLFf66gvSydtU
If8FqmSOu+2sT9a0RngXfR7WvrNTmV2t1jD08ob/LwD73aYbAq6uhDl3PWsv
GlTBfZM1N5XRI2UznDF/97QGXJGj67OKSFJ6gQS3/gHEe23yraN9P/1Y/E6K
SfqmACmQaPIRjQiSgPSTNMvBU2MEs5aEMyHioc/5afBmMtIOXZsk+QRPW5rN
VIy8VA9dJfT/ApvdC1djw7pRn7XqVBr2ZuNBbdGgPXUkX3BLrbwucYDq7lOU
SxhOkdAxGyc6VyB9bzleXkf5nmSXJp+kVGw4l0pILodLzniFPZi4ljldVqYY
RIPmzrb0Il2nEu0amhmawzYhZ9nbkYX+mF8YnWK/6TPX2F/eyBq5RqfBTDq/
I/EEYHpr7sA7YeyWwJ6DEMeVLgFcLiNG7agbeXnFsePzXW8mH2mb614nL+ek
pKWUfjGEUc85gfGsjOZWiDGq6m+HNBxmCmxbKgHLofTTryZwc58r+XY3fPzc
a71jVyYyIiUQWmNNevqdK0LKlg/SPogoF6FUt4ZOwfosJtvCLnkudk0W07Zp
ORzaNXlmFNrXJc94iNJPYN5vq9aqpkl99XOB54Rdry3KCX99LyXl4u4VQqs3
+K9Va8vveYm/fAAew+MxrlYx1aN+YY4CzZ9ZRT69nr8XkMCAEc/+Dso1yvMF
VEm91XBs9nTdv099wcZGtCZ7vLVCfk+MeeDWpVUc3lSV4XE9G5EFrnowGAkl
niKJR790em15xel4YyWxBnXE8ssRp5BYl/BF5mKRQ4k1J6cXQ1ie3m85UE2f
vAkboW3e++01HRZ8tIn/Hbj1QGaOVOjCdiagRdfe2aabTg4BJU7tECt647JK
Jh8z9vOzCaFt2vdJ5U4kArc2GNSWdYToenhqv3n4SwtNQAULmVM8LFTSozo0
vtca+aLh8icO25tX30yyae1awOm+vtP/1hSVBQ1sZ6ifSUZU9DwpRJgkvoAq
oH4N02szYwD7XZ5fQWrE/yi8BOWNBkAfPl03VxBcA1O3mzghYa0aiqkrMBjD
JrzyNqNfzy0VQbRXokuToO7KXIXx8N2uiEKrTe8dEim4rKn5Fp3fSwD1tEli
ttdYR9lNKwzeq6lT02VCcLf936Z1MJSW3LbZxpHxMKKVO6eZa4hZVmYzI1Qa
kzSTFg+JBza2RlClev7xSvKo6MAvZfeOeXjPNRetuuFdwdVF+3pvxw1Dt+uR
JAmN3+SVqWOiOforNyWMVvcxVAlS9PPbZ1oajmSmPPE4HqE3DTGx6mHeBJCX
Bq461+NnEjhQCJ+2KHZvQ5A4N7E6OFv+1g0CJwjZ86FPZcSmXMeEBuhmP4Jr
Ptm5nN5n8/duWT63Fu+t3NnO+IQjovRkX4FqK4Kw09mW1FiKed+rgvWpQoP3
EgW8Oe9V0484Ay30QgKkRqgK31Wy886Yqo5y09Un25sbUvNB00bJ51qd4Te4
wCIUBJPfg92loizXJStBE9qXJVVupdFvrHaboFK1MnS5WeLlYAQU2xM2Vkap
KjgG4Q22b5+GDokCGELsiVnU2iOryliJaU6cNhexgBrJwMSmWOn0vir3urdR
O520Hb7LAHLXPX7k9J8zHl07QS9zn/psv2paFxKgzg86N170k1kxkS1nK/GS
hBQTa5fUx+hwyaHnTwuraRzN/rpFOF6O5tHJo/C4yT1VIfHCPj5lBgzCRAW3
/8fUxE8M7Dh9QOnrjxqoEgA744BOJ7GA9dPqs0dgaZwcyijW4paCKUy/0ysz
vESnvBHhJ/NpU6nFaosdzS7enyR/CerrAwrIIGLhO/wH+Xr0Mx2MKr43QoUS
cXwKWgEGRt7WstAPt2g/fbBY8zOVidiNwBDDnKVZO6GWRArxmP+jMAkKxv9x
H35AEqac7IHeabXqR/d0cBT1PRsxG9CucrVzPVfuH0IlLlbtTNUWe+ZKPZ2j
epcwJl1/o2+wYT5aVQWD/Xd66Vl59xE0oGSEuEAH1tdL5i0W8UVC610UytTJ
fxDWU+n83C4VCjF02MpG973Fdp7sINfSlglxElg2oZJ/j4KKjzste4wLd+sX
jvCRaAXYxvPQVP80WUz4KZjs+1vdraQa1W620qvshGO7AnqYMCAR8IOeugKD
XlXBIBQq2gMtTwZMIgo6LPWDl2N424wAT7SYByJwXItrwFtRFhGUb/D3+ulG
6xiHN7qH/cNYyr9fVJXjUD6aA2iucNOZUfks9ygCVg1ddkzJOaSTtd/DV7e9
rrNTINOr5FX49zZipP8cUx9xrldZrg/9RE0cUoXok9Xk97qTryMK0dOyLj/T
zWhBGpKtaOBg2Xhj1BgBl0UFBOXjBD6vw+WxWYGAN6DtlZ0hQamshz2Dtzq4
TSE/5X/txf5ngDiA5W5Ku6M+Pk4B0k4fwiEGp9EBZCYzFsvKmoq4aALoGv/n
vdTa1HN0V/Emp1jWEqO/murMTDCMUv3mFyKD4smezLazN4SsezgteYuHmYBO
kT8bgUhXYSBI950sDwUOLWkeaZP2AiKuob2TN79QMiqStKw/u0zhxkr+6UrT
If5HBO9KA8cRtHdA/rJXPacQ6UJdsfeAybfJsOU3e40dBwAQQZHqzUduccwx
qzDaN2RCkbAsB6lOyUBkYCyMeoRdOSQrg9e7FWZOlb7VZUuu8LC7Kz7BiGBl
vrB7jNLzdlrU0g+rU58mPOztCVLs4tIxB2C/VUZjLybbjbj5OjnpEYX3QMix
TUoZEwfrXwJ9N6ukeQu4KzemMqn7vcIaAkOsQjm1OlnepLS/XajRFc4rbEX7
XdBP+2ln1EFyFw5egYadIVWY/BmfpflKDg9gvfvvU+yQMiJgZ1kWHo5zG6PK
nvDpf9thcsGiAMO9zgASPF6UrLItMR/leaGJvgVGOHT8MiDyIEI18nzxbiF2
Yw6oineD9ywieCTTd9HEQC5yHfYkuAJNEp7Oa/TTYR/Zhxm7abGHyg6pvHxX
xZ/q06Zh44gU+NhUHe/58hPeswW4VkSedYkriSr+Wr+aUrhti1zIsCKyZEd7
YSa/RMzZuszIrIPTf7wNaGOoicQ+l8NyPWfP4P18NvJSVcSZWPh1Dylj0d1W
pIokiSpzjvTjlfkq5eXGcnjtu7IwrYVaZu5pUk9Bz2ZyPcsqTcKT/4ebxnTz
PSnnNDja3Q1XwK3u+zUH/WEz5reV7upcJtxbOyFFxYAnXXrU+ZLgvAJ1/r9Z
SIYBcT5QVxV7+yk0/w/IZYtCgwWCrtg5YCfGjaO+XJczvY55hmpX2/kqtzk5
6sS48h1NOI1QHMucAWsIHseL+ubjM+feP1FfwPvGnL9rVHpCpYLml6eakby6
WV/8O7utnrOUAEj7XFcLYDeZmJ/z0jM+1sYKZLCK5qJ5GQ5yo+GVOya7RtsN
TTChYhn6NIJtq9NK5rTOCYHbzfowgx3MX07jRRgaq1LBObhfpqMKjuf8UIKd
K9KZzJL7E6Ly/rgSG+7MjskiIbu+k3wQQleI7TApbU9hNGh4mJJz3A6sBYKx
Zsdd3S97kPydoH0XfUc9xAIIZp1bGd3n3cSyUA8ufRa197p8gkOHYZUJH/WH
CGN8qdwITdlTIm+242PiJc5E3rw+6mpsIjP6hykulKKT/oBY1W3SKTVkU74O
a7lOL+gbD+zo4t6Vh7Hr428D2k3q6n/+vzfvxi+7lQAz+3dWj9AQePnj1B2P
2iAqrBwG+bDsW3hT320IqLqWJGTK8L8r03mt5twQItNzWcywIhtKxK6fQTN8
6wDWt7loP7cC0dc1kddvz9BYTZYvyedgN6uavB0cwR6YxFdbBbRSbftozGeE
+biKk9FEfv6jYYtUqsMUBXBpT4v6c5e+xg705Q3Tyz2QNT0bZ6SxoeYyPi6I
5eXmsLqW2vDiwXXCXTQ7bWnP0uxFOdpO+bvAICfnlZf7gOCx5DwkQbcq5vJS
3eRzvZoS4WwYrQQTJHyTnwStPrUV8i/+zjrMI02B2gNcwdtXysCn3qCQYGY5
4Es9fKVOMCvVkdJ4+gzHtKyfX5J+apleg7gZwoGe9PX25/YVPKZji2hjIx1n
qv77Q4s0n0L7UdzvuqFSXtvO7NnImB3TVWtg9v4q+3upMFB9CnvNW3k1gX4J
BuGarchsZ6XrcSvFNlqqrjHF3sAjoq1CC49YFjS8AuoEGJEVL109BQDJJrfd
FaZK/uBoxVgy2XAyMzK7ZsjL45K4ahvKULLnOG266JmMw1TFwIrHk08tvKjB
KE9W9xGqh7D2vPkVbLLaKLBr+5eMJFHuvJ1GgUzR0v80EUH/1R44jjd6LBgW
9nvtKHsfDhLmf2pOV3g/vMRo0TlYI9RrMWwMFG/FkUt7gYE75e+5QVZJrqG4
SYDcLmTxGhv17YBDKR2ZojNjXpCAVY6+RWQcwMFoc02+vtNUSBvMK8GWBCz+
FxaRcgELj6CQddfXClqEe8/4bhV2MBABm4vyIXXbmHIEDyChY3f06SDeBqDt
EEKdYtzzBYmRcwxX7g0RLGX+5gdxuCHETdbHwe0wdVeK4dCanKwquYH5AzeC
X5Kaa2NRdbcZni1gH4CNsJmaMSpzyIRQB28TIAIxzZRA8ogV2JTY23AlIkMJ
Y+/xd7JozytV7aK+O2ldoJ5tHzO5RGx8s41tUfWMCESWAhXOxb6SO7KIvZzH
uC6Lo/FHdhBZZ5t08VTQe9GyI35TWPDswbG1bKUGd9gOC2elbYboI7QDfprB
UOjqOkQH2k4X1yV7K31wVcu3tzHE8yxb6cpcUYK8CxE+iY0jh/yeO/98TzXm
JUqLJS2R/ttX2wZHBjL3pSw21wSnmourcni0yhFpJxUEfo1mOtUEqEsUIi5W
4rp2Dwb9MpJk7hxWy4ufhbN+0jE3tFBX4MgXBVqF6jWZ5BlOjeN3Rk+n4LND
16hkYCYd1NWNptsJcmL61+qR873ve4K0Qa2/fI86LXnVChx3lDggD9qzI5dr
dFzwePoIkQ4ibR3ITH8NDCRd9h5GHoEB59WHzatHduki2JGiHUS01FFfLdto
x4OdhpMNp/D0B5gVKz+SQQKLsPPfFK5fPCrhEUTR+O9GY+tgQSM7EhEMHlkN
GVJomfKsOCZzxfE1VfPuQPBYfeWI/qqUTgxMXlYs/HmfYEy1/MuKACmfx8j/
3e465KpfJ3hNpfbS9zpLEAMW9IYfsjhrbifxXSkSrK8FiyJD4wYcwwz06Q9X
Fzl1yDFOrcikeM4qt2TyUQef4uLrCcSprTa9kYqwS0l2LYDUdlXyHBUqnEPK
y/fFyvP07yTstv+TR/CxSotudIeLLtie4k2iIZnvDd8ntnkmNQE1I208EfgG
0zl3jZgD7Y+fLApSxs0h2GvGLXL/xfsU7PXBUAKG1bGv8PXV39urtP+mQ1ze
mBdGmM7jtUxJ36u/ZIHUOBD4yY12fY5CTbCnDRX1i21/AtQVcUgpdO0Qw2O9
3VFMfIQ/D1+QJaGKxqJyNpUL59Kk3nZg5s4uymah38WyxKiIdeLqwZL2aK8c
N1Jq7XTxEaoZL3nRED1XLXMc18q7xK01H84AMxBRkvX6RbXa/TXuBK72Zf4V
+0WcwtaOVFJ2rwgJteGlWKdndIFxALhEtcMNMt90mY1CuRnJFBWS25FqqJeE
/Hf6kaVQ7aHhU3aLrl0Amee2AHsWc1tnWRDcmZJBUs3V8VibqBmEwT5LjLcC
rsXC0c4gr6qnKv8Q5lvT50effGclOB6u+CpJUqIg6fXmKn3q1sm4q2bNlaoC
feufrseHse/YXGQ8gtE52lxltLT71h9uJhmwzRwq3t2HDhVwDGxasfRic+V7
6q3XS0aIRvoG5rWLMQQgdvKHy02Wai/MYxWlWXEmKFUEs9P8z2nwIZDBARlN
lOfSchC0Nt40UNEb4t7GzEl2HKcdIqrsxjy0AlqtRjq91b8o90sX7GCJIHN3
Oa1XYsKhQPb6DbrIb2n+2ptkEtZBU4qD09w8h5dasnXG/tz9jagrf+NbKTY7
VnYU6anrn0iqHG+K435G7djgWwqIQ1yc7l0T68l5rWASOrvr5J/ub0p58dAB
zYzUK8qfQIXft71C9dAz0neRJvucD7gv4Np5iyJca9SaUuxHa/xndGEryoEW
qdxqkQ2c8JsWqm3ujvLO5AEJ/Wm1epG6ctZ2HVX4IFkG0K2W0Y4EtlHSZK8G
BuPBPK8NnzsaO27rVWZD5Ijj/4hEEDD9z8mx4/e/J0VMNJiv/7HkqrU/PnN9
mKAVN5ZRgOeof0YBV9xJOv3LjFx1r2ONS6pm5Pz+dDF97mE2weRJi3JxVJHE
BWrHB+QNyM4F/7TdETcT57gsnqT3k0eycK4axADhVMudZAPS7BF7CvkI5Bg0
2njNxWNpLgxP+wosWbrI+HArsMM/4GTXLtzTG28d5qswL0K9CyJGr6q0KRY6
VmgkZoce5tkJTOMPSQLQIMH5SscGqNnSau5zje7yiLmIS3kl2j2VApSS94aF
dySTsACYiW5YXh74gu3x+kcT6mwDUT+KjuX7NnvftF+pQd+igikD9xvWxN/Z
qc4TnrojNTWPK7sOwkPQo/XEjYEgU/ZaH2FfZ0Wks5RkIPruaVixgTqWm4Q1
UF4JDTcM9iSHRiZ8WJVPddZuu7vLXB1i9Uoo35Vi2qoD2jHvZ+/a1qsE0UQn
BSvOla6JsRyqoobBhHjnvoLjp0kXoHI4kfSdLd7JGv2DaBwOwPP56nJNFfx3
vftTksqKEQ1RSMmaz4LidTON0clXEt7aD25kBwJBNVejlrK6Ng4P2v0hiAA0
/WzqRc5e0bKIld4Au6mQ9GKCc3AnJrXBVrA6337sN5///JZSy0TuLPUprr/9
gZYVDa574LBokDPueZtfVlxJI+av+un10zcBjjt0Ps16CUwAVjH0UiiUlmZ2
wMLC9Sl3bviFJdrSHB5ctrn6u+GocNNSfo0DzCD9t8jf+/6abeI6L9xJh17A
BfqVDMp5tEHLD729ArLkPSOfUE3aRwe7mWhogezKYkQ5sEt/+Nmyl9TyYdHZ
SMDS96UH8XH3lTlrokLS9qMjwucCk2ADq7+Dg5hDsOejB6YtlYwQI1zSxL/z
3DLeyGvBqPA1Q4CwkltMYa4Wj/m7fVj13GMLGkm72KChhYLMZ7djjPP902QK
5OeFcVUT0BsnCe7iVv91Tc1si7i/eJVdjXs3hzMGukyUViSX3cYgnXIgJy/e
bSIx0v6zO889AcuXXI6dEZkcfAxoeA2NqHZZNQaz15wcI34PoniHjNcTI/8D
VLQDwC9LGd6O2YMA/VqpIaWIz7MXFZlqChcMqfK6kndH3aBU5QQlQ+YaKFei
Sr2zZfhchE88o4fu7vtjGG3+v7Oi1bJwR+PxP/Qo5sDVpYOcSXlb20MFeuMf
tms20v9uEmY8Y75jpYs4jlh6thJl1nrTVYi/TbVG7B59L53lGS39Yb9hpxQI
hhwpp/I2BBZFcVEELDK1gnNypIT022z8I5zvL8E9QrXZ2mUqqFygRe505Urk
2dHznlRhxDYoyI67e/SYtV0cAby7ZP8Ux/stycOYGW/AnujdTBDK/XEZ87/z
JHvI379HWt4oEksHlx8mKbysJOUqQrG8w4hnGISikap1DU7F7CuB4sheRP4V
f8j3dPJog2wF1+67UIXvmNN2Y6SLDtqKX4X2sa0ivlZqEiwnqgAa5k0lrmqE
qK7TWEJBwCbCrxZFF9d/aC65MRQGJJccLe9XLJU26b6Yn8pPVuuGjLlesV6j
KNoNNk1+W81/W9AGoJwQsy6rvSRycaGi6pj7NvyAyFjT4TQsN4WRstry4jic
GLqLAFz32Xf165rqT/8njeB0DMEedqqOJi3gObtXWG6lluSJ8Pkk6v6xfk5R
NwF3DD3DFtIX9JN2Rw0hf1rr6iBw39/YRCbe3BUf3JcDuK+FjIWxg95ZbyZ0
RwnIgPhidj/v0sA5F6h+6YunM0b8sN2eApKP1nSB2iO9AAtqMAex45AnDw3k
Ro8RVqqkZR8LK94RcXFxHNRjs7PjMnRiE4QWA4DSoPnsaTHJE3n/ebck7WgB
T9R1zgRB3KpZ78ULgufjwKftrz9RYKw3JbidDyEXt3XPSB18owGzeAT8CaSg
AuOHt8cv/uOuvBvOIjFqGfAWEVlOqY7GT9FaRRP2aAbZG0G4H6NFMiy0KiZZ
6yxmQPZXw+zxQvXRUrNIoXgePCL+tHoKS9CBboaFgG2+zJ8Ad1p318ixTW52
AOo2yzP2fT19FBqkt4KR9+wa1H/2tuFuXhWYhE2FKUPhsM0Y6OGr+6FaaK1K
I+hXQksHZeraSml+MJC2eUs7Iru/SAT9ZxZmwjAA+2E+ugsm1wzRtHCsJW7i
Iwsr6syNU0EQmydqVL5yVdDPiGwNhH6q1a+9SAKnNFlljUoNs/kydFUNnVkQ
qnkf9Z29rhlaS9UckYYp027Q9LePNtFJuY97hlauni6xTweUDJV+xkvF3SfL
ikSJFuAXwitQCvuln7hDQzbPELwJaYx4ki5WjwLHVWV1+1HEk4VXC4R/yRIP
Q+MguQXNzW39i/O2JCmfRkur/aEUGf4sPcrneMOPbWO53c++Eucu/uoM9TSd
Wfuoir34PMhl7nF77JpGGb1RYf8HzVxBbna6gjA1FgStbLUHR6UMviAY5Ijl
IcK+VKlAQdw63f5bIYBkg3+qqw0lDuzzQgzCshUq9oHCJ8WPMZOx5c1ZIc2q
i7qsSU++QElydkjxeVr1gOzSJ2gufGRu8EN3wE4ScBClyCDOh3UDE+GAIgiy
fWmdfqHt/UKxRNxsCVJUSDBX9/34wrF3Jnq7ziKHVMAdxyhujd46NIq7t/Qe
4EdzAf7xZ2XNB0qxevlO9Tt29fZa6ybsaW9T2wZjgxOAS/KbBSzEMPzT8z76
sdC0lSfa25OzWO3hSyNPlB2sv9y90WwgBybKn+EYOIhvAjtJ8eqMQ5WJyvHx
LlMrLyG2AWhZ47TF0UXTQyQOLHR7/iPMIOwOQoatqXB6mKLzT3PZGwOARB31
QejWXuDwLB0NXbotjwAbvylKBLVs88p/3JOiTIriYj7wcgqRsimKh3cMl1oD
rDfyb6tTAgdkVSw4Gm1LvsJPZBMuXACpYY/asBuq8kuZ7MalQmzUO0A7aIfX
YT2D4LMGb1frhFoUvcUyMIsZGTWgWjVH3tMyZQ28bOZrdEMhaDiQpp7b59nj
p0YMQk2f+m4K7Bymd2Ge3dCufDhPAgMZqdFI+nrgdcHghK+3TymJ77Kn+6wk
aFQBTEh6zogsieJ3IZpwxAuAnltlUWTdTHd2Ode7Yp7JQBYhzP+zeTjqgID9
SNlpr8SpoMwthXIF2RBNzgyrOlbyiytMKbnvT5TjGkU7sxJRglpUHj5MmeXc
iplEKM4QlG6n896e2uGnCwr4FdW32NvzwDFpKvSQh2IsrwEZ6wKzJpuZkBcW
HRlsCNGQvNVg9rl9q7BzOIiC51OWFJYUFOdeWQMxKG+CwTzbmPkeSEV5hqyW
OlHj16qIUGkwzKXa8H8MZPOcwUG89XRcgyNO/dgQlsfmFngEltd7Min/+JWF
89gCDlyMDIylcZnToJNJmRL6By4ADo/wywifmbrV4vEcSvhhuNeel3EJxCHO
r2hKIhBjnygEI45JVb0/5mwLKzDqTEZBXKHeR86U/ra8lCBijZqH7cVbQ1K3
PdTWXcWayNZVEsilk8Y8SI3ZkJZSmzxTw5fCgO9JGRfFml9M25Y2OK7gPW0e
0DmzufGg7VLWXH+b/m1UQTmnUQCf82iWVPBqXEFC5njjpMAJLSH0gvm89TCD
eZFDbETcVZXl9ZIr5AUrr1s5eMyxhaERxP2+g00EjYwSVVlZqm0qTGG9FOhQ
C2Qem377xgZGOMU0YUpAS3HsMDFeGXiC/83ByjyOcBHYbRcvQzLW1U/BOGRv
SV+my8wbpRqyISw3NSWOixxitryKJr2m5OlAXGfnxVPPpHrpWB3PoWIe8KeM
G8iYDwjqQEtN/Sf08Bc0+MwBr0kUIYvojLRgjIRMBK0O2PPSlk7Wp3LT84yd
7NLno0tbhzlpxENW4dAwLPhCmj0XF52nB60RAOWEgVvs7A44fuXiCCQEgqB9
fE/j6cQb5rRk4FmJiMXBAg+8vY9NlhOZwiT5CokCfAjrBZkpFhMpRvjeai/t
k/KxbyqFysIsJzL283IJV9TVMoEoKtxnUGEcWqs96PtwdWIwIeFsR8kYaaQA
LSHOroaWn4j3FeYZ+sa6B3dQkhXfV9dgXCNDxhEWclSy2+Uj9VGa78YQZJXj
QAzTmUjTtf4UfXFS/uIT98dOgxddRoi6bp1DazbQuWhEGFCtuK5mEcDX/UR9
RrUDOnFwgl0WPEGH4DJqla3B7QJ5v1ltl1LoUZnGgSX2CS1qPrCbsHp9V9sS
mK89qFPrGhXou22kO4TbI0SO9YwTziQNYMRKoredm/AXe1bOk54wNPlv3xIp
SFo+Qxo+x7FFYQU7XZ2WRzDrvBtl60smZYo9cugA6OvZ0phmP5NUZPnU1VTM
88VYaO60TUD47acZVIFk2crqXSGaSBuG0FnYZr+/OG1N4k5PZiaYYxMBloXN
5zjFI9+bogOPpcDnP8ZO42yqqQQXf+jtW9MLFs0cfgrO7jxZQSL8A+1fM+gP
xfRNZ1FWSO6GJK2BMVUt1so6eezNcoZ41886Bp4WRDf6yO5Z3u+JlByt3u51
Kv1/PamosqB7tmJLZ4T+4qFvlr/YNPNUuyglWIm1rCDj/uB9GDocO1VrS9k8
RqTOfodFOySfzpAFUWFXmwK32sUfOXsyoHSmv5A+ec55xYsDLgXqVTtDSBmq
e/WsHUy+Numy/K4vhhWlEer6OeMrCOec9J3PtR1hdgbDUFPQcXUI6X0OtjTK
xaeJdB81ZsbXWW0CpKacpSxodHB/snC+f+M4xk3sbxZPFhnnsLI6eydhgp42
VCUhOux1g/BOPRZkDtJxLF8mhWgTBN2fFf3pU8/yGq0TdUWpFnX7jG7UcpBa
EklktH5oRgxs3Q1K1WhbParrFVLBLxQsjVS+Nkb1wncTzOUsP5/R1o3ngGtC
xm6npWt05mjwdU2ueba11DtN2e9q3UTJjpg/J/nUos4HtP9hZsgj52RlATf+
gHkUyFPPz1sPtS1cl03CefDrK7doUecC/VxnUSd5lG2aHhg/uBkMU00/LXyZ
iPGAdvKotFq+RCeHwLOr9HD/PTTgW6XhGBZApZBdby4+UMv3BlQ5nr06DxQ1
xtLy4apN3EUyeXhOsGeuyLCarD3h40pOWVlz0qbL6ZLHI1e28cjWNxFPfl7+
TD2ttY9vvlVVEINPEITXTISn0ySuM1gEWKg+yAAwcjDMeownAwCUYbYZBald
bNQ0oVgm1x8HX6+AhCs4EQE8zxY6lZbDu5BI+mjkUmBBRQVyXxvX3WKgjuz2
2Ggwy8KfdE/kgyGdGuOvnoUStv2a+1TisdZ0OpiECAWnlJvixqD1+K0ACegk
nTln8ebwdZafciPpD5zoSje+2jmdnZyuIABImScTR9hz7Frnv5qVG1sPVZGF
F7YiOg4W/gcu8ladSpHxonW47OTXC0/wsIMN42Jh5bRlRdlE2JKp2WwYhcQ1
KwSly8a27TeWi8HY6ZkNbkynN/o0LFqpt7ABKuVp+wNtr+3eL6zdVgbRPkrZ
gw9hVr5gS3RuiygyvEX/tV5NHxtXCCSoHK2EL0BDPft6Vaoc9mIxdfAE7m7d
VSXWMzFfRoKJiw51k4Q5igjcgAH/jcH/kVaY5pi60BESB5tqpIt+m92fNnSe
12WNzB+NeetMTh76BmU1sh5dp3wwQgA+NOkBxodLAnwn79m4y9jw1Tg0Vb3s
CKvPELe8fB8bYKjCVHbjPSgSfkcmAijQ/XBOuMAgOxauuTST/Cty8GMzpCzX
Q2ZXCV3VkqSI74yzeB2h2mkx3PvFxcMhPk+CKOZ3g9Ke5LcUWk24SXbCCAjC
QorP8HKV6xVUHqBK6vVIY8QrDqDy4ClgszcaqYW2JrQYktsgqgeMr5I6vc5I
hEajYo/TudKJWhancHUjxX3gNXXpmFbz7AujfGxvVOJ7QMqpDn7aVqX2Qeg2
mYeh2/rk+Wryxg3ZHEPq4uybhaLbRWXGWrJEEL0Pq+Vgq2bBc5PG7no1sbfg
mZSbm0JTGpYz3JAwOHPdEfPwkNxUXpPb3LY7HICf+IFio1ps5vblfSFp/zku
FdYFucoX6lF3ae13vb9EWtM4x1JA1GIf5VTBAgTeIwZ5oSdMlg32ULKYsrKV
HALV2FztwnVzG6Sbiw+1xOR2p36YF5soQfOCmfWhNJ8XD1pyS8uWOf4uINC1
A9DCaRlNjVfSPfe02Jf+KMXGuRe1gez7r/+PfCIGtYpqfzcJxKedrphJW9mt
k5UvyftSHMSGpNm0XfcIaPq6UPqA5tcDARsUAh4VdoFZHYvw14f2iv0y/5nC
FMZni0ibMoNYobe6mUCn5F6y8TFvvUMMFZSq+lNRT2VDtITMdFfyfjg4eXC0
8qoCSGHPe1asE3Y2rz0s/SYVBQpy/3/KfukfhXrc/gjt/W+JO51Ihu132fCe
/bdSAIO/O1kp0tn4yobfIn6s137E+rolBAzVKF0XT2i1e8D++5oLKjDlxXnH
zIxbe/9wSTfHAh9Ah+8i2zJ70sF2CSWHi2Ec2GEDl1dvST4wqLKNSC8kh8DN
P8qtS6/S5ViZmWPfwiBvba//NGSK+y0xMXhZ8+7vYgOkyk3vplBU8mK4MI1D
C6CdmsEkEO39HPn6ESgdxF0cohoHAi5lRGshISOYKmE8toKUC8c+30PZmrtJ
uUA9R02UNtM7PZDJPL1+sHf21Z2ZDHsVoVWgPYeyZyuI3vZOeYBk3/n28yyo
wuH3RHWxesqHvJqh1tq1rU4OZuJIuqmcBh7Vcd0uruSMmzAl/1/KEAPu8bFG
wSDMqMLuyLH0PaQ5S2loZqe4A1sjlnLpEulv5VOt07TNVqeeKNfbwWiebJkM
NqRdxGg063duPPtQs8TOnsKBlMArEs47Hz0XncAdsi+cVlIXgzJazBl6n/WF
gVkRk9/dKOCFSM4YEwG9/kcjFmb1xcQrfFRrsi7blyBMdPG1FyKRaZydR+2Z
NycdgkR4pjFgWOGnAqiF04gf7u6Q6rAvP/WX11P210WkvQwZ21uwQcn80Gne
hYc3x+3B42qb79H4nyOvmawspZkoUl5dcn6vcErXUUwIrX2aY2NNfjJqVh97
cCet+tKWlceejWgdLi3Uq0wJT0Fb5TigS+OKYX4Q4PyhSjt64QQZIzcWFgf2
duHovYjGVPh0IGOP/0TNKFYoKr2WTn6bsPz14HaWY1vkg3/ZS7aMQBenoEey
nTGOVcMN+JRa5zEQ3Z7G/FjYBOedNxuGbfAGaXuojfQOnDr5LCFUE7mWguyV
p/TBXZwvLpZKYSTj1FEp5Xm/7DHPnZllC1I+NzzUU/aQhYECofgxsL8rwwUo
+waCp0oLfVqJs5n5m7Rn7OKGQ9pvG33NzksQ4egm209nqK0aHZt08d+M2zv6
FH2NSC1NdMccybaQOWgILJQcFBqzYOkKxsAzklVN6QvIUlqiyLVPYHltk98V
QIKqaArSf/AjywgJyKivzeaYRml5Xdcur2LCEpRSSmDKDDr2tU4Nonqyq3hq
7MHhAjc2rBLeIGUvvDBNzjW+Mm3pRir2x0pVb0tBjTqWcqYb2zwL/IoxeW9s
CxvBUtrO465dk0aoYkw4xyosI+JwtX/F7ynmdb0WZkE8P7ZK84SJw0w9inin
zEua9idXGkk9bkq/iOfk4nThLBA3uMGPtE/LSMt6gyrB5sw5Mc3nXviKsCHf
h5VkD/6awjnxql3CQeuYp3zLwecEnC1Xb7/U5QA8OYUPiVi7tu8pQ/GCFxeR
2q4PoGTbtKSQfKQ5orYcW8yUUeyzdSbW6Zjso8PKEOuHfb/X6bxwLlQ5hpw/
bidB0STSLFO58bXxPz4veyl3Y9dGb2jCRpq8Cz/99o8EGvXQxNCCzk60JS1G
RWo/lKbmycT8NNvaSnlNma0H43PnkUvzuviDhGj8vpd//2kL0MILu1XBqAhk
4dnSpXc8QVHu4ZZXgcfEn3sRr2VuNwlft3dXp+KzrzB/uptzjxH5kpQmto3f
Oms/fNK6gp3i1a6cyKjMo4eQ1YYclIm3QWvtqXkDQ3d091PrQHG/+De1b/YQ
vKwUz5eAr49aWkDHm1Q+rRC/PC8Wvu0EEPKqqHWrStYHS0qJTZZeQg4VD/DK
eaBfVlGJtyGBHnlJ3yglxwKWc1hcO9jX99kfYgic3Z1F68A97x5+qzhUiZd/
dCIWarHRqel89yyyhUa3wZi/crNty7xHMOA0Lx8f8a3AKH3+M88iXNIvXzPM
r9POOvK3LonBrMR+P6fx8RvfL97loMp3qsdmT4zdHjFKsKhTGc+Jq9wEqd7L
l9yo1nD77v+b9AOa4LkHYltEcDAhuAsr6q0k6pkYiJh8sBlzSGnM1T8K4un7
kFbLB7D/QzNl/HwcZDmA4ntnCIvj9ro6eszEzY5HHL9x8DebDj17EIZRdAH5
S1iBtRnNlU4TmifVOApaEAfu7t1BYaz7SG/0lq/f2m4zAh41lBGXjHnm4yAt
HlTM5HKDtyhYcushHDMpjz5w85jSr+t+4t8v7Nd/gB1nBSUJIAKbogRxVqrE
ggd/jBuJ8qVH+ll0XybLojBCpxJARtCAdRA7gWHSW/HOJWUQV2XKuuIlvCM1
+02Rr93IHV+gIT9VunR/wOrgOnxFzUxE2Aw/jE2r8Z4QaeowOIUYatlFxd/j
L839SV8AeAVg2J2askl21BAitw3fHBkUpZja1UfjuuhRyedE/r5Qw+dCKd3A
/EBUGXNOSIwAnAP6gCtnhAe7/OHr+NjCgdxb1tG5l4Yg5ZWHwodSdaePs/MF
9wHlmQZgiLgCQeljCCeZabyvq5nw9QOUY8OGRBtlLJ9BpAnn8aXBGDi98eeQ
kC86zoUlsqpXQtKV3rvoHRoVgIaHJ2ShfB6Em3DDzAB90qr6o+f6IUdca0Dt
YcBlLx0D5Y/+iO3fmquShblAy7L3mH6wPUFYUq1ePjCmxtdncKMu2yjPj4L5
6kB7TC3zzTnk6IBcJhuvFuC7sJ7Jfqc1TuCMpCjC87lrndwcEIMKmriUur5j
HEb26/RXB97+ZkPBz9NKHGdtwBSrda66BPY8t+sdp+KiSJGCNRRd9/B2o/Wi
Q/H9VNOiJgk+o02di9IgNG38J14x9lORQDQDPTY7a9AND+015LS/MEfYlNoa
lNPEWSPVY4Jc4HM07ZCi2dgELeBKTYS+1CLlikW4odTYP0+9PfcfLJa1oyEL
jCG6JKI9HmqA76puNCzbkaVF56/nysrCC20pByNrv9O1b00bB/KIJCj10xcq
UXCOcjfD/81OObUMK7mxbd8Q7z+6cmK9u51sFa2u3/Rd7lXVTKGIy8CrAFzy
DwoxPkFlFtra1jrXkkrp9WyclW9BWTm5TY2vTLvVhzsoFIUL3bPTZ3evfrms
Df3jWQ2aSKhfPjNM1BSXA69/sHjgcsaDpMtQdqO+ZPUjZl32vbnXuUfYnUIY
+JlX9Owe6ycCCyph2hhuxTMB6HUA9ql1br/aNCm96RahyVIoBS3/8MlGrzdN
JUXbXas6CyAQdTbBzWH6mXB7OL9Ltfg8n4cN6tYVZFe2b1UInaR5tCTXjAld
+A6v0qt6B5Fnu8Ydu2U+cqypJIkDxUWayLpu5hYII+TJ/CfSrypv39DuGiSN
V0hVLvkJ2LttNNIL7aZx8+yQXLUOcKMgtOr6wcs/Y2TL2Cazq8u4+j8FwYW0
QLVU3o2FIb6d128tXb9VXubHXmw5sQu4asGWKuYAyesd+FUyTdtnO4uPqYZJ
BQfuJ7rSy/S80J5KolbibOZS3w/kZR4SLUNC9OwbiZ0i7AwW4oDBjMrz3pK8
RnOx5Y3XGbidr5WrXZFpRQYk+DkUSkkYONVUj2qpxLNtRuzitoSTHqOLUBBi
EwbEJF+iZA7Z+arprcf/R96kxaM3kC9ugck6p69pO/6vi2G1i+Bmz6tZPx9p
yyzKpKq50glskVxj6C1ifmkBb+ogw4pkptboTL7dxiuBUsZvLH4gMjIHpj9/
c+ZR+912tyhMcpu6HRx6TjHRSTLEJQGI0NlQuo5gorVZTBVfZlo01yz90RXe
EiigVJ09X4GCIj/XuJ1osjEs9PS0hjJ2f/3HeDpzZAgHqnVfj5iMk6pxuUm9
DiHrNxQrEwF1oYLcnVlYqS2vPGX9TEXvwF4Ty08KIcFXpwMKT1tO4Zs5oIbj
YgegnzOwh68OS8HoXvHPEVaZiroz1AUjRNFZgjQz5trPHx64cydLHq09Cbsj
Cj8790NURak6LNYrDfvfiHIfk7jmpOf1xzeAY/HIZcAitLq6RArN2mOM1GaH
OeQ4/1czjrg90mwgeN9MpVQCvqoJ/NVCEEfXCXASvDBH1Rew7xFBIorZQgkC
uRTICBblEzxF0fiX6N0o6FlY4rcwQRDpMFtFSASA1O+YRZrOQ/z2f7YzVFuW
KtatwERrtE4scwftpLb2U2O3ay2QQgQ0eOeQ8vDO7b+8AoqnlX2ikLHD0nk2
eSxdN8nx9JFG1Fxs8I0stnJxjEjIwQnIVARvH+vPV9SuJ92bthoBITxlC7zj
C5FucRE/HA4Rxidf11lSmc1h7nYxeq0oM8QlGlQXXYfPdxSYkvsrmWc+y1r9
XhGe7gamHqMW9SEyxuSahAUEnjq5gc27SMB7J/jvw8MoNzcC5VTdFSKfpIBw
MdxFfoPrb/rkCum4JGP4zjcV23zuC4ZGwZZAo37j4MXlGsvYVOjsDgXENAyI
XlFRp2rstJSuxVyhxvgUhFTuvhZ6dYgbv8dgFq91hLaXJwKoFD5vGs1qot0s
n+04LQmhIXIeklxU+dQhddx9PoQZY2DrALC46IzwJbI41BxMauQazT+kVskm
SBzXxNX9Q/MjfLAiMaC3fdn+ys+wyn5TVQqswEZDH8zYIo271yFqt0M2eifX
JILonxN8lIP4LsSL92sOWU9CFThksefVNSq+hE28ZvX+/znHKGFhU/KJAH1P
IyKPR8FuCYAzkM1g97eEJIzuEpzcRXc8wAQ4vAeluQcKnNWzavVKRqosfIPO
jpFaHTNa2HXU4QtNqLRaVCcayspeWEqcDSMhS/nO/iS1cUiFV3yh9Rwnu1Uy
mlXBNFXcrsJS66xfYqr8a6t4rZXb+LhpnbsLLpIhfdMSYnr8jl5u6qIGgtWZ
wKVijHXzQo23oZTBJhsxdME2kCI+T8AgHulePqpWTU1E4rnzQSw6SbNdJ0KW
v+ek8ghRyCB3fbOlfulQu3UuldGOYOpW+DS2WuQZuk2szjIG/iE16LwEoy/h
1U4zlvCI6ftxuLiHuOxRFAJCI5lm4OGguajcEfkl+l3lrj3u1+twh9NL0McR
ZYaCX8XngF3enw5cInBIaMmRdA1s+Gy5dFl3KVqk0tlyh04CG+tlK6+LVQsO
Hijie8ZLFPMUI6TDNEoHsUxmKPTBRjHzsdECKHYBOOMBbuX19JcvISm3C6MK
i0yGBB4Hs+bZaHFgclwwFyCbGnOd+3f6AFY2sKSU8XQ3U0m9FvTAcwforjp6
sxt1h3RB43VdY1c2VBFWf2DsZqlVkbYCleYUin1Co41PQ/Likm0f+bs3NH6W
k+iONshr5rA/X38YsN5jya98v21zHIkXvh3XQiTSm2cRqA/CQHrk1MG3Hlxq
ApWparytvOlgLuYYpFGD5ehMKXPz+6Klgudi1Z20PjQHBO4KELxJe1sT6Hcc
P8zE/Cbs7MMF6JJ0JZf85/2LkjlRqJp6ylzyhgOllv+0UazXOyMz9w/JfayH
lZsowPByRCnys467jmP/UUsUQ2P3kqLocC9Ima4wLpmxSGzByVwGOorE16i7
XGtw3h7J2WD9gVjQtll1t26jSWzh5jG/qD8ggIShCnp/UjQ5zJUtgMufh3A/
Rjq/pzpF/T2N2QkkYMFpWCtADLNSDzT97ZcTHsjM5/uBfYqO40Z5KDA+YiI2
06XRyEBJL+C8WVKdLR9Fe78AG7djCaOBpPWy1nKmOHgATputVErwIVDZfGlP
5YRnRWwvrbxCiZoKj+H5KvED0QSxVGXM5tOnaNwnUoaUhdtrYaH3p3ibDuTl
6yVe+OpttypCdqC4I581bngPCt6tUQ8EyScyEXge2tptee6Wm7a5+XpivfwO
/p9/WpK/M4rTXQRaSrEsmTUoh7fFqlh8FXZk7f3hKj+CPFNUBH5kPSoWCPLT
RcjpeGOLakR/QwB8dhMluy3T9e6gZR9eseVVC2fQ21aU5A1mwIRL8gjdgfuu
8W4fcLuhNRBUVk1sm1TzQBryEGgYwlXm6AoRX6qf76dd+Ve4gxltoAQYDHeG
iBL3n7ATgrDLnNxMw/HonfjMgrxqheRYAKOnlbk8K+TQj/1eGyGDZLbjaJwV
akdELr7py6UD5wTmkdG5u/92pAnlw1Px2ZG52EezofRX4J07pYnO+xQl0+vk
7UI04nPnlRwzroR+e2cG7DQepTOSXE/T5T2HzbxUyRZ5tCsiDn/BPL1EM/ef
g7Jhe6BR5qRq1eL4Dd8r0rs0frnUN1PygfjnCwlB9xwVh6LkBnbb3SwxL9hH
aAkvIJ5Frwimc5LVettTDw53tjFwyTui8tO1EJ5mWoRUDmGBb7mEq3XH/naE
e4vFfqUbKpWkM3cFCeauScUWEM/5H6Gzj+xAQi1MceYVb+evTVuYQwZzqgXo
RmeDfIN6IhiazL0AXrkLpdO+mJ8XCg2JMHVU4e1e9dKI1NkVon8+FFJWtHmm
BIQyteNpD4Yl7pQNsAlE5a4YEjlOsZdak3FngLMiOXMpycbwgHY/MOuFgBWs
WX/gHFel3lvBREcGmmO/Jri6SVwy6Lbjq2XRQq0v72zEICb450l0eGlLNUIj
j42Xl32eUbKZ+MkhTcCi36s5cyDtDi5JkFZFijCf+BWN3hIKzn092oRAQzGH
GtWyVn7Dbf3uoH5hynaYMY84lRVzPiYn3aiSbHP8m+U0DDiZaMsJobXeXq5/
UY/VeTePWwXOdQ0s4JacoOKjtLZYFweyyEV3tN4BE1WkpU2nP9ZTBqEoBKJn
1nxwBOZ4um7f4XeLs7mOA0JNXLoRRhLcZ2+6NGFiVXN4mPgHQAHbwH875ReD
QJeraUSxIcFpid56po8UU+mZ3178C/+jhZMOMOmlyVsJZnhnCbZoGipOrqJu
CN0gdHtEGFIaFzZXkq1+1ouX2cyTwWI0pcV/GAv5NOhnXVIQzOgSf2Z8HcMg
95mptPJel6eeKwgYrWZSPjCa7++vlVA+kdZD680sIc1raZQqRKDoENnm/6n3
xaNdSetVaQ58bt/ig4U9iflWtYdvaWNYqpKWTdKU77Mh8Aiu/AfUdoQ4x7Gy
JFJIw0pcnVz2l/2d5Y7PRCQGAIo1n+0TVELxYlrQP9bUlCF2EkMWvP0YQWRV
UBRfEFdOLw22MoMyrASpIfzQmWegfChoUZUbCC7JVgwCu0KMW5J17V/4kFqI
DqK9yO6YDR9KMlcUFbUE1U10itlVPeyKsZtW2fnWiuGBydzWSC5KX5C9nvVq
2oWVnjcfwo0uoQEWXHd5PLefNA+VSikxXHi8aDEZ8aWbdnPg+s82Ggw9Xbtp
2K8gBtJC/TtNB/TET+/GK3//XP8nSjWpRk4wwIIBjf3YvibkPl2TodrycEIb
6i1KZbfU7fs14Sfb4LkdGHFsaL7EdXHXvMkI2v0RW9ZZd53Oj9s3rsg+T/S4
PXjTN6uyY8Q/2aeZepMdxLcUSQyAOVgacDH66t2HQzOhUSg38xGpVGxQMDxm
8dbM11x8bmRKIzcjirMyT4DS6xcsuwJjG59B1zwCO6uibTJstzS/Thmw6wxd
ByfwzWPZRFaFGQtR784tYHU6TVQVYmqE3GJ3cq7nx+j4M57U0AofyEJn03R3
b869ys2gyW4YPUkcQICP/YJztR9yNeQ0y3V9cpNFsc/1cpWutHmkWk2ojrzi
+DP37bXDBLG/LY5KEW45o5M2Gcotjlt9fs59Gp1LudpJYEHTg7jw/bOvr/su
JHtAUNcG0zNtQgKB5sWx2Am+uOqBsSKblm5utD0zYXBB94jmr/JUMb+5s/O+
t7xPZiggjSunQxmjSjAUBL6RpEFQg9dEKexXNZCn3p8vpWJJaBBO7aiIoEBV
7zyL+5JZiRIhZMZPmCTrTDlAGgUaz+rsjqSDICEDHNoDqydS6QcpyB3iNRYq
EMZrfM0vkZxidmobiBzKwt/jkt0RjoizhbhR7iJDiEK6h67ksg5Pz90uOPmQ
1QsGGTMI7AwOo9g943l3fX+TKlzI5/a335b6HyOHzUOnezNUvAAvQEZCsui9
NlfkvWsyVVdhOqISohprd3lJsPlmdyQSY6/91Iv/fiE8gaUd2rB6VeUdqpHC
rzO4O4H/vwGbeWPlQ40p0GQsVfSrt5Vvrfm55yfEdk5Go/zoJ0rAdH1Ck459
KorocnACdRjVaiD3CIb3EWBnQQWF4wa0LdynLregmU6Ov4bTiZDD4Ahcb8h0
QZ99wnxZ2avzroRcsZ0Hsz0DgQJz7AmVn6/UfO81R74qM6Bg7fyonuNbR4kL
zK8qOq7FlO7YjpHNgngcjUTWx4C893HAwfcIoCQxFi+c7wC3jwf6QDbFdGc0
Xgo7Wz4xKZa7IYeEWVVOaZyitIXF1Oo5zjEE3DVgJi9g7A7LFahPP2aNCpvZ
OsxYZaf88iMnSf6CTnPZE7DolXOMdctYjBVPRtp6PlhKbWlVSHB4O+wCjp0U
2sKH8rahumsMMHPC1WgM4Y17053Q/lCwBB+xpOGN+zXWCkjYzDD2wrIh0QQj
cpDXvTPmYCxzeFvt0n2xJcDk6sYT+eW0HD7LOISXAF+THdNMhmyHgyUcro8w
BtKhXbaX2IUdNQ5MyhdBwcrww5ye+rBKMHtTBVVRCTObwscWYBHNGoUXnZ7V
sQCbr5UYKYO55LhnzZaMluyaP2mKYzmLnganxYsqEy+rJaJZhxFmyPTV4cmn
YSOk2Pl/b9K3Zv3Zhe/ijIPl+fGYP94qEDfJdzJV0fTEhYfn/UcmXDjmklgk
zv9HUdRhhohGy2k2O2rb2QzpKxLffPGxBlw686g0k3p2rkcL4bSr4pCb80+s
VHnn4ImdleR/aQ5oiXjl3UaqOpGW+sN5AN5+xBC/rC3mE2pg8q7t128J51QG
hJ8na73rYaj/7R3Ch8dE9bdf2ifJA9rclIw9t5NnmZH4d5ZpgRyvZm4JDXUG
zuydM3o5a/YEHeVh6I60BdQbCqErH/BdQ26RQSix72rWNoXrjhAwgOPq/iVz
9F4DsywSah6cyHQv3UGJ/Jjo05tkAUoro+3HC/z07Oyd9Gwi54aUGuE2oVCG
uNduSxK7ijaxJdfVy8epOdb+vYXL2jNDzUF4AjD+Uyx4qhRbB0qLcsBfGrfe
pq452Ii7XSfHcw09fWXywiPmnMyE13VeFYeRXcSEeNqi8XYyEqbf0/PbiBGm
Fkon7nolUvB4qccLYG4Tt6YvDkjv5EabXO3L4FzeNfGO62F26BsPJvY9apXi
VFIcDlyHGpl7Deqq5gfi7k0NtOwmc19iGkXCrHC1qjZmdHLo4wQEKIlCyP8F
Tu4CNfbJ0ptEEuaRo4cKKomyjwE+I2IuyncwJCmSZMmFh8y3Gh4lGzySOzBp
9t+IhIPX0rtvL5cTu8SehbqfylohN9Ra/oObzg2tWv7nbRxt81O8LEeKC9Cp
/mP9jNeZsro+Y3PLHhp5PMrlWN6YP3hnYiDIZjByT6qiVXQO5fEx+s+qPvQH
S4TR9GfqhxxTaYF1sLj2SckeOUh7Ty4jz8hUvY5u1mVvnM606AjFsrvoOe3T
cwV0+R1L1m3FjidCo8c8QIt0LPMHDJ9jFJXZV1aROJIW5Xberj4fVd+RXFU/
DCfDiPbNowXz7C75hoxhuY32LqkmEmX7NpO1SlCq/avx1LMMW4FCHT5eYRMV
7tBhNcdlyy1k9WotaJh/sNuw3W7MK9pRyPFro/Sg1hDV6O1e0VJKa8WFiSU0
OBcXPAFNLuYyLfyyhfK75/zdBfGQ1Jl0V85e8ctmEHH9WVwystlVrg9sWU+8
UAelJpu9f1htmPr5n+5t+sWqa/tRIvwA2nZkVGxPbsn9ehFPV8nWeucLD7WU
T7XcY41OWDFuLsfsowp1q//QyVs55oB1SFs3UEjZGXA5KC43oL9W3PUZ7YV8
WulM8Mg2YeiKC2J9QS5TpcRosksg5yQqlnkFS+ONW8bgfUWFLSQBmv3j+oWA
hIbHJZPfvnfpNCqOWVUtvr/HztPgvg2CTzKFRfOwwEo1wRwr4J7Z2d0e/woB
I2BDAGFxHx57GtKnmqs2+64Cz0MgjBxBVMeJOUfI/Z/KBu6pnNNt1mpIRWYh
fHcCpFF0K0cxQJCDTRoNNLJgs2Z3BpskaZOrQYodQHn6VLXyVgQPL57TYm2g
mxCuTKDT6btZxzq7UeUDxvlo4jBRS5dPPV9eoEc5ZKtNPrnHuudoSMca6tgM
cditbaaP0LDsKADNco6fJGvADrSW8qH3RNdzldNO3boNJJERgAGyiazCpVRh
Vu8/+GVDSZehZPeOQKKsDnZ4E9w0a+GDNrLEiVgxz8e06G4yk2RVFgUKR1VK
dBbutwZLtSxAf1CmTti3KLcc+GcaSs9usGYXYBRu4hnIKgtfA55WHFUgv36c
O/eq3cPzDRwqJme7+/3QQrwcqKH0sc0TI4tWkH0sMhXa/Tl5KEYAxirL6T1s
5juVPBJAFdJtXjiPZDjenJihxssKzLvmG/Z1LMEWMV2etK1cfY2t+cF8Mxp7
m20ziljqShLgIv5wHttoweXNLOa5tGYLWOwt/QfxaZ0MVtNiXSL7koJWD4pI
QVNAzHaBSMWcaSy5zB9qpkiQwZjDE+Fnv/wOqi4KZ58Kd58Fg9mCgrJVj2te
aU5k6KbK5pZDErOiPyQpx755LyzKNKuSeQ1IMUhtxZtjKO0mn8zcUZTI8ixf
5q3wm4gDEc3HxCtb4GVBtUzRLVegd/bARBBnK1CwWwmoothxGCwN48mbuJkf
4YXwLBZzehkk9S14ZjQypYO2lE26xjtC1yOMzrL26wLDuXHjVv8FyjPAH4pQ
3vhw71Q+aLbiC4HKZe2OWUghFRqgLnzI33MN/vzt3zyWiMrUjja5tXiTRM+b
D2d37SQ0PWqJGmfXrHfkjiajzXIXIHtZSRDRT9DF9KBGaFSBXAjmtM3gq5gv
CmRYlduR/l91W3dIDIHXV58ZJjhHihImLY9X3SuOkcDD8uzOTASHWmDZQRW1
XyPSQ2Ap85AdUUG2FumYclT+i7B+/HBWnmsbjL5XzCJAYvBLMjife7gKceE4
z3jtjrTfict5NiWBYfrAkeqBbIByxfgp/Y19ohh1fSiWdpB/vRRckJ26BCUw
RDr/KrX4uRUZvhNl+G6QX4iqcgctXrJkXcex5dAer4EPwUdRQjgLrvHHo16w
6MSqtGkLcdRmvHnYyHZx5lbOmbfJPhpgyXEecwTimQkZkm7W3+m54wbwj0Wb
OLqQhUZVs134YlnFlD7hg9cKEkyhJfDmTXrEM4avjH3W5EdBxb603Aiih7he
DE7No8tWePPOXATnSxNnfUj1wlbQHuNTYeEEZzHjeRg7QvI4Ik97YSVqbqK2
kx4LeF3sb4Rbyp5XAHjdFElLJdf4o5RNVOetTQv1pggNi8WnGWj38b9HxHTe
wsL6TEWygHohNwSiSEhBadIXIPsioqrE5aqDOujL8kqWeS0B6SY8s0SxYIfg
GDrLpsyPnQBYxK6pK4a8Fre0GRHttCbzH4xixZFbYcPs/eWSg6FUuRzmKX5P
KBn4/7OAYauxDE3sOKYPzxWT0kqYJ4OefBTykSpBKRf5S3+bs71G6PNTyhVn
S5t0DInFn3D64Az08DY0zdDZlvGtlr+qP5uSY4NQjlUuXBy0s7UWVG65x1w2
C7PyJBO/wr2RBKo7NGk49dEul8WJ3XM0pBAaL/HxK1zXILdXkfK6LIr3lKCh
lGLtn7KlKl0YSYxrSkqAbsQQtMkcm832nQEpmYN7qmq3fE555fMxMRH24AUz
J77dZPW1qdTYINLaVpybOln9o/sk50yFBtVaDzuHbX/zErUW6pTpn8rTnw3S
dA9Dnszu3/Z4F8bBm7i55/MV5YYCaIVpUkfUVCBVkC+8TpMZrHAjDRJSOm2g
4oIDTCv0juQvDbm7lbZgW6Mx95JJvng2Zvw97Ub7s/bHxOwSmouqpdQSMQWH
7veexKdGSJqv2kdFy0+ztRykYPnM55PVtDRuPul7fH84Yy/I02xRYoyNv4FC
DG3jm773rkNqPGj0oee/oafyoG6wNhLZpu2xlyvhX2ppjAXO4mE85QbjKnfB
1x1Zhvj1+8XCv5+kk0R1ZVLFM09KytCP0oaRKAZHM/RmEycnCCg+TixpLwrT
NxO9ecc/E0cg7qBcMMGOQ+m2/KQIL1WJksvQoio8OJMXNfFzDbGiGRP2PIAI
v93yJUwbzNoFfNgD0rM6Eo1gpEF2yRkpb09+1Nvh25tJcc4tOJUD+4QmL+St
w71ni9uWwpSTpq2/j9saGdfQBUbfq4xSdLTHCJTRmc1/Adt4hpTFRJM9JuM9
lRujip6Dx2Q9gOHVdz/Bq6M8CMsQfuuv5urK5ofkxsjP+ARVt7aegxNo+/Ec
+LdGqfrWzh4eFTvqeEDsGwWBXOP6xFHosy7xjyolCvHCurzQsgmXLpBeqb2V
bZsyncwTaIx1g0X+3lfSgL68aQI5giUEQ9Fk0yryh5F3zY+L1rX63cIzdisD
kxkmkKrihKa8MKH40ewqCJ0rlHGsvGYhbWUrJ4k7YR+7tyooSaBDJGkllbrG
A5WCZL/dtgIGVz4hjV58GHQuXkhl4wOc2gzsdiNrAhJ8HcJ1yh7rF9MmM7MV
a07jab3ywPp2R041M1lm8iTbK69gbvizmaucJ19A43s/N4mh4Nz7B9J7IIOv
UQyqWPLscG7bq5pyPZF3uh3OcQBe1Fwa9BAP8AILIT5KL3/YHLTlW29vPLWP
pEfoelMCBf5agg174wO63Y8Xj2p61SflA4lry2t5PwI34aIRJQ/fpZgiCJdL
0qFcgoYD0qN2d2SQaiHTf+k/sBzcMvj9T73DyJ2aDuicFACAWYEo3cQ4DTJ9
O6eOhPIH3qyeqJndWnlK98NltPwPBhrpt4gcT2zed105dtokeysJoIu3JU5P
lzoegTspbSk5irYCF8JiS9wHbSnpkECAQYSt8Bh0bBzl3WYqTiY6cygIUeUc
6808s0GX1tjWEkNx6qJxl+C8+DLp5dG9DOAZ9YpACqrnuQRidvda9TFnl+jp
CrcUBM7curAwnfu1aC+f5J1jCfdCUe9mx86dGpMFmJk6OdF8vy/QxqZgJV/N
cRUNIde7YYsyAsWh5bzcHjEaFRSOC3gIiWleMCJkQ6LYXuH28kXd6Kh59Wmg
7gQXk86esBvznc2m/MUYE7Gh+kmH9rZxptvkjW98eLYroad9gRCA+7kWcMTu
C6EShLZFsny68jFsPYx5YAKC+zoK4riBP4Mpd3WT/jq+Ca2c+I0TrrGm+vMj
Ulq40yEga2o4Nz/sGzrkxPWOxhxDTBR7J0LEmsSRd6kVf/xVGr4DQrri8bi0
pJiPiCKA/EmO56zclv1M3AFyGScwr1YkX+3LOpyKsmMdr8JM9I3JqWUwisbL
pq4ZBsFAJ5j7HqoMsQa6x8CRkAn1ODOzmPQ68qq80Eyo5LWRPc95T7Ir+kGX
0olPeE8unTGQ9Gv94EicNawYWuoxy/k+Gp1UjKl8u492Z4ZRdRBPe3EM1XoC
OMrjWaMRQ2nOvDOy5+MAMoUcRhV4jbRnz2y4VtgqrALWQlFqoRDXi9phiTLD
vRHnWx319lnFlx/YUz/BGWy8MvriRJMvp0IOw1PgOxHS/YmEe1g4IrHok139
sPzl89B6MbgukGG9zNwFBqrW61aXaRjER6fRAlN1T5JH3kSmQ+uudD1chE9f
Z71UZ2SRat1Aq7bU/N1MSCEiRVZRbOvE2FecImEWdmoRGpD1XZ3vdy84ywhk
WbrQay41cCkHH+nWNRigktqu5ZK3vJtigALnNmtt2LldSfmhjAzd88RLYWYL
VPPk+5kkuqdxws/AKnhhoxaJY+Q7/Mnw7YiCrvl1n/1gzg4wDAcvEDL3iCQQ
jdfLJR5gENrNV2uCP2VEXej0ou9bczhYXlWCOpP+UbLuPFoSKIKLNsbQGzQ2
EEhcWl8uqGPAvNruDPZ3x4PZ/I75ReNFKcUnNgq2Rp+gBF6TDBI9wW2lr8p+
0ZOmKymbE9WFNzrTh/g+nVVjhDEnonbqp9ThxXrxitOqynCPlMxhPUTA9Hig
69rS3lvh8w/BzqKbSle5oXgFIaxjfsj8H3jz5mVsXVshJRDF7Ttpgv+SuVs6
GAUL8cTlokQyLThSSfTgEvJ19ZIkodgiETFgVdp0lOROImjecH/sKLBIKbBG
3+NzQ+Rb4fy1gCLqO/6c6/3soh2mtlZZ99I8DQ7Ga+ONaoDYc9taNv50swUZ
VfJACm0wQGOPqOw213h+FbkMlOiOQJbkNzZ68sjgMR7rkAq/vXBJVOqrbtuu
sHAK7rby1xrq6c5IsHa2UhPusiE8xv6R+wx5GnF1Fc539RwrarCShS57ptkR
6xx9uZxXc22c94tzMgt6+BWbwUkpF5+cP4/1HdRf2NoLMavtdzoPHbFjmFT0
GZqkZP0QEXI65eS4zdYzvDwCzeTsXIGKhSUXg8fob5+xtfBMcK/lmlNalt45
SMIagNHQT9a+qKyk5UWwllkru5G+gq18OX0XFKFUh1dnbwZ31d/Yobvn9qhJ
klTK21QqU7cN/iDtc3YxWnSVSYetf01MmStzod06s3uMFsrwGSLJKSVUQ8hL
QNRRvpVhvxxW8rSWYcnWncmTwT6r/3PQaIyhoGf5nGEPZPpMpmWm3LsxuK6W
eErk+N9RUWLB6TJtoS8AbkNym5UxzweveeSdil1YrFE5FNN8pUELV8Z9djO3
Vx9q5ncfx9ZFP6Hi0Yo10kPqecI58lUoIkffegVZ7OcwegH1AZO4IowWqjr4
aHI3g/ZIFCJI4qnaK0IcSq4D8ChKh3yo+gM+HjAYxsBeBHyLTnQFO/WkfmQ8
PGjpuOGTSJdJHHREEM5iyrfEJYwsYThXNz06mWA0BbJfOtPVzZN0mXjVART3
QtaYJXvtdJRzstjJDkT8WtiF51fup6lTaT63DVYg1rkYA/b0aNsJD/+pos9D
yTq+NoNqVYt0pSNjaGVHH1f4F1JaPhDZKIYOdcSVx87XoGPiXQ5eAW4YoBLb
jg4hW8NRLdcZMU4FQrADoKiFllMQ6Kb3U+11Lgf7P3qi8SrxF4OApn3JggbZ
bxKkmilNR7YBO49X6agKWra7I4yxhb0kwU1LYL/LyVoTivy8i7iGolQcESD1
SjSCzU6xTDNJqR+VlgaYW7KASg5zWy/9v+DOLvGC8/HQCppS3V9jEhAqPAyl
+4pB48gjiM2UsI0gy86Vnut9xZ8z2kp4kIDmSKJGW72IIglaifxaTIZyNgxm
+6eLi37y9UyRPiFmBP86xhPYLMmJ7qleRmIguYkVLZeqS/Ga4irFXuIx2Q4a
ADCoKisEtRbC/G5npG5P6mEQrjNa88euQJlnsPkrVNf2MirKqGK3OzqrkD5+
GKAg5xjv3WDkfbrcEguFRlllO553O9xzZFBbxotRJDX2BACM7/XznwtZp1GT
n1ISdtFlYu6916zg2fswQ+qHPFNCeB0cl6WsbLleanfFVdNCxZ0EG2xjRxeA
g1TszCt7r7tGU4sMYCWFKiQ66l9wxu1diUrjOMlT6/xH5TzXQmrEs1XhB42N
RIAlEPVJ/unKZ2mGm6CXWvqxbRUuYvOCWIMAwEoitDRVBvsserAsW59kj6Y/
BaVsoSUvQ+n0PRzkwu7TL5Vu/CKw+troHfkSHSVVXkSTgOMa2TiACIGWG0Ao
Fog0+SMmm2xG+XNAg+/azMXCdYe3iPsUkjJxHZ7RO715zbkmanQbNxqiBjYO
ThIS+Pab4UpZhIVRRsHBSb/eg3ki1DA9jgAqEZDvHehTd8GH5XVrE/365C6F
cTlNWc0svUvNIcqV/ldL3LTg8Nr7McYX6HSmv24oARFf4DF/cFDD2+zJwlF3
Hov+0HStxXHZJOTmx1m77qr00KCzEx+bhkn7WppMQIBbkSclPUT/cCdqJDtc
6XxzPhwDFfcLnc9JIS3xNf51B9M2HuMJQS000DbqDzZkYaa71YdDFSdJD18B
d2qGoftsanHV0+XOEe1k7aQ0mBMiI1Q1iyxRVBmX5ZQIJosECxEdCLmH+fwO
TI8RXzBqrL8I2h1oNF/IsDpOG6/1Un3/Pr38BoV+LXPWCpQvlM2WjoyBGGfA
Zq7um7FTDZXa5TiHRucZ9CWn/QDF6NSUBC/FI0oC+HtKVwkmyh+Unyqin/kO
69U6g5p3DXQZsSTaat4FY8FIxc7mkZ3m42P0UF6ioAH/OIoWkxfr63Wg6yxC
F6uRKcZyExW4KLnv2gqJmJeG82HE9EDwU2s8bb8ZDlegsSTMUQMBMV8n3gNm
gfn59H+KKSEH2fMZLYXRCQ2F6qyW42mIZIXupmTJ/lQ8WNPnOhR6MMfZPveZ
R9CK+RiUBlAlZZUdCGx4/0QQ1mpuz9Oi402HlC5TlCi8iYBPyq+FF5AZ6Opa
rMLECpRHwCmM1keIEIxc/49CZOi/LI7pYHhSFcTiAAlKY7I3Eeo5pTwLynwo
hjnPMtbCw0VxLeKp4YJh3LhncAUDBXgAb1rD1JEP0q98R86HxvzHDOawisDP
YHgFYaLRskm4IZ/LP2NcUQa8y4uDXEEHkhgLxaxC/VP3HWFoiSdAL/Bdm9hO
mrxId+elJ33WybXLBg+zkebjFIijzbZEfG7rumlRebSRcS9YwTRULWQdd4sh
1n5bGQxhr1IRJZpGgMaLsbXf0UNm09DGfhiqFKeMdJh7llWYHanZh76HPdlR
I9fm9jvcpwajHyJ5HL4et8bXiWTufEwF19D0GHzYCgU4mtTOQEz4oZbAk27U
3M1VsZY/J7B07KaLXpUIxKEPitzYCn0YewgeW4+q1j92+x7OGBnhx73/jLHX
txcZGvutucCjG4d44WcT0NBNqlmRM5qTXNglIqGsFhRBDQIXCH+kTOjzpCgS
13n6eLhBgN/fiU62chx3HdDBb3f2IR/5IScXL+Y5lYvT6E0St+1i8WQyMaHh
PZWHdrN1qP3+GffzCtyjS2W3C8e9iHlMVSKRSyJJMbZ22/GSMa/8axBh58tp
/lQ7WoqYHYjiUEmpzF1Dl87AfqeYCHzkDBK5mAgOIbT7Ph4Ml/KBdT+z3YNG
bNGn7Jf6fJRx6pmqWiLYzXJTCGO3IzoMrh5Zvt7aZcAzZsiGaEiPPuq1e5N+
t11ZUbhPgc2qdhIE9ECZSm0m/pC6fa92oqwcZQ/ty4obvsODPuDYJTPid4/p
HSshQs3jYdU++NGqm4kgeU+xCIfNVwaqsA6aTTzJTAPPPZJiX3iDJWlOkSIN
tzei9bahcrpjJWBlDnEbesE6S96DP83B2i1Gyq9J0J0kPuIAmmxss1RISvNN
FU2Ng3dJgP/WyQNENO4eI868orYloyZ0VOTX/TlKflW3YOjWHmQQptwx2fZt
owQyYMw+/bxxZ4IC6Dv6Oh/ge0tWWbiP1nDaNSBvOgG0RXMUpldkMOtfhlfp
5GScrB9gxXJXc97vMx6s7n7PxtesJXGkeLhrSRKSSnwQC0ZA8nvHC+2qgN5R
2X8URNlMzgQrusHiaaad/X91/T5Ux/XjStOYu+NgMGWruTPpfxTwPQLBIKiG
yEcZ7OK1aeXy1nivqls9TvtjldALLGlFtAbgtYCckpugN6EK8AY5IO095JZr
ZhtJR99bFkzZ9YdKpQu4swQV16tLSDi7U6aI82WvuMUSKo1Dpt2SiPIEH5Re
ni9+goiQBP9qRlAXgD0+6exmE9AjyQ7gCqW2BjLNCO5BFjkzDYwKWJzBwmmv
RRupRecMkq4oluVbCsT5JKaB33RwAol3TASMDMwvmlYRsu0Aq+SkrnNIU8r/
nODtjDMc9tdhZZq0/Sx0FI4mvDqtRCHgMlYBzW73rkqSgBBffhgJxIYNjB0b
NAamutUUBfsftBUrl+UtkZfamUgjDhxodm3M6ohoemfvMzwS2S+PHTWy7dDY
+m5DrH1JybIKz/Nd8LLqYwmzM1mSffY58xZ/KdnB77A37zsDhSKGiJTkbDe8
xMfBHcWPWDA6O0QhMdvqzNDzjdzfwb5mM4SmHHeY5t9BxvVybR5EbQxgoXF8
GNy8IOyKqVXPn8Y/fDJvatF/h1JaFPU+g1iEhgSAuEL3f75focoALKwqAd4x
S5qJoyca4bEz8jIMCI9OCi5XJPbXNgpE8sjQ5O0179IQo+icX7yTNlgXrVf6
5W8OX3ht7xkg0nks+Zl4mHi9aSxaz67TG7LmvOzCZTNSMxQ10Z4y2CEVEY6j
IvEJYlNAFMbeKogd/wmOtULq7RQV4fMoyALG/RQirHufbKSNW4O6zZWY1ANI
+LgLpE/CjY9fMKNIGtsdmxuOdQZmA7ZUGEZ0pmQcPJPGjoGfbz6SqYmPrxDO
1YHWclgOIm5ro3KZoDZgatvcdpMPvfDUGPzGHhrfUCA4Zq5PDemmA0qFk2Aw
afazZbLQEfMeefh8aW8HRHK6O1RnUn3w9sPFKBJwPHCsMXaXEk52gXHTvkWI
cBMUvSc/nUsqFj9sfJz2UUFrKkSNb2Xoc6ucXGDLQlRHF2vWFREujS+eJ98D
WcyyQNvD3JjesJmg7vcBEEeIJ1rc3FNju957ZvHquk3hKl/8N+w5kwuxDO6a
MkWPVS4PzbrQqIbCSy3YVnk7Vrkwe5bWFRB4fVPWTjDB0FGe2IpB/23l0NfL
sLAOgrb7fd25/cKjCelFJzAuzca11mmrSjXf5dJPFzrYTOZsK4GM0j3Ur/RK
FgQYYSWG2ocMeCKMQGHuNn1hr68ODdZFG0j1SNckE0DQdIBs6j0MFM7SuYSo
sAhtyJz6Wy5il9pZmxFb5PbIjNpownDXzw7tMJMDp8mHO8oiJgDsjzzPUYeo
Uihn1WoIUAAoiucAXtNL8xZ/oELCuJ7MaBXivDHpBFbH28b4VDoWPx0w7ihL
Y6N65fOUFkwBWYrJ/9VSzCMIqNlAgPNK5RZuloC8h8RQnZO1VEi9j80Hj9/D
i1i9NaV7NWateAihQAPf1hrBhzI2y7i5mhoV0jJakbDq1Caxw8i2kvN7GAXJ
DWbOHF8chDSgIk0EMkYzs/GCe8ODOGWJIfJV1H+gVjeGln5iVFFCznAYzJI9
zSb/ha1wvhD4efL1BbTYzrm7YbcO5yCrXfSYibuIeMymxXVcPfU2oHAdNw4+
9mlTdjx6bTev/WL5UcxfZMzHyO6ADcuPw5kLh4Z5or2EiE+4n4bIEEoB6Kek
7/tgQBk0GA73p28gJJeSfNB78oGLKiYQCZxlg6RCOIW8PkUlJpyzTfG/bw9m
DEPQW/AX0fssxHBHxZya/9iMXA9Fu8YwRGW11fL1qBHls/LhBMDC3ta8JKBX
nrlJP8niq3AjnAPHXwoBQc1XZSfoFbrR4xv1B650H8gzmobdgWplSX6rAXWM
j8iPW9W2aI6V2iBFaOk1XQwcv5Fp0RvvdSNOAfM59kqtuyZZRtIXoKDb0DRG
lfdV1axTC6SkuYgmczFfLEU0uLpB9+tjwEeVK49NIM6aLPjwUPe5J6zWOuDS
xr2SdTodzWFJq24GOEgidb1qPhGGJdRmBWMGV0LnMani0Brb5c1sEQSz8vQa
BIOWoYN6NJY7gSi3YKTBnGu+c6M2zqHu4QjxcCwpRd84cZav2n8U3j1Z9kmx
hMTxIhtnKsrX/8t5BNbRKkyPE5tTPJzSTIb9HUPF31Xszi8gg7BtH8XcOC6y
Yq3aDhPNrNboScCzFlQ07HcRBqFHNDIa0D7sQnefsMq0powqrarJWEuMyrpK
/yT4JHxXdBS7KR3oSa2WdxsYFZgyY7cr1Evzl7dYixU1cTCC8WFRRNDFjbq0
kLi1aCP90tZwjyotwT1UeXXDd68ff83WM6bbOYI+Tx3+l+ikXneNtC+/24Sd
Q+9+9vGCVInd+gtDnBt0mYX0Nlq5fLvcfmYFkHs6JyNhWU5Y2NzcZeBJWM9i
O41AIazFl7w0S1I3ifWz3gA2mgGo7V7Q7vaFSNs1ixjQYpqKawP4WF3x9XKf
RClnoISFNAMUK+4Iflo55MUSjA8Dl/IFYlgkMUwY4YTcZ41LpGoZ3xdG1Nt/
90D9L1oyldH503iwfgEuJKSKzj7BEsZGIjFwOonL7/lNJstkJ4/CJJRW9mdy
1bIgIH78qkyrHgO8n6gYHc2CwmDmYuke75Nrf3yLD/QopWd8jRg8AR9XQmy3
n298TQmQ8MC0VsgJw8872KWLL4CDeaLfHAGpjqiSR9y1sSblTQ2bb3NC3jAj
4R4oy4qf3+wJpTSH0UWWL8/Ukz49OD0bCHK9C+ijW4xgcE3m+iD93crxyZ5J
zjwLKUl/ceY/okEjoE1gUhKbGauI5gtBS8LQwBYYheV91Uf848Zpo81ZTzxk
OS12xn1RbVrkyR5Y/KzlEM0x/HjGvXT1yMvr4f5+DfRvcMcLoAb1Hvu4R6Qf
Cs2Z1NOBE7dDzMBI37qBhwt1Kdi0VNvIyAPw3wCg+DsjrdIhJfksM1Jc0tIV
AI8mTcCbt/lk3sBSeIh7nyVu7Nap/HsBL9Z1QxMI1E607rE7DmLO++wnr7uV
+OMABZV0xA1M3o+fNPij98o/13bq56Vuo/1XLp7EPsl7iojiILCABYLeXFQe
Xb9sHFYFeFvkJk7Paq5G3KZTSPNCzHZRmadHNR5W5GbbzNdZo60Xw02SYyft
egBwOJPAI7MMQLjPC2WqcSWLX+/A4P+n+I+I2gst9sVM8AWQ26mHy2jiPdsh
mLbWgc7dPb/T9XgcB0s1VrOgkxfpVXLBC3A7n79lm43bwICwQ3vEFykyYxnr
dBZbUBT4R05vHUhkjbSOSat/cXkv7zNXr/ZjTFnwN633DEO78zn2bXNFJDi7
wjnYyBnX9d2RvSvURrRlK5xoFQMT4/W8Vov2+A+FffhkX49vIU3nNFCMPQyJ
HJ9ZqylYAPhP71lZv42t8YzykpfrBRGWwe1gFuqTIo1uExcu2F5kggqvAg0e
RRkv81gcPBUyOmjSh/fx/z1S9C8Br/SiWTzLnUN/nqXH4Zu5fbJrhMNhTN0q
K/yjh1U4RxLgbTAMoFBKtYgsYDtd8jLTosN7qGEZl5T2ZcPV3MO4A5MRTFja
gbXD3zPwwcweY8rq4oReukwTTfv4P5vwV7fm0mzO/tLQ+jqmu7JVYQ//mWIX
m3xnWJQKOr/lgU/4QHlkIbk1HhuWtPGoKkSROBvX1nvo9u0GtVFUdlFkiTND
qt/6DUdHKCth2CP83f+uDA1rfw0oFzZR+CVBTcyEbZLmqAwrlSVykUqe0sWn
60bbpPgJEUQ9HjDjZEQCJalysF5tF0PP8otlq1tHgL3GheoCztlGFLM/eBXG
iiUtQdSbZiSMXHE6mBioJ2BY00Unbcc8KoEZ3CqfV+LlboG/rbF0Tqqkn9PD
pbLG3mAUuZ6Nka617h8Sw2UaeXON9x35+ymAi/6qpFljFi9Qwx+sS265S+pk
m+J89CfdhmX360xHzyI1J0yWZdeylVFlPY616mPNOF6aA9aFYx8KluIqrJk6
TktFFn/+mbp67nvECtLNXqZEknfga62fyeivzf7XZA0t4d+KTYStZKf+NimG
lDNSKEqja0XtiRaKkMLXn/ISnIRplxp8zqZA4KS0Eg2RSAN0HZxF2ypv7d2q
QFSpuZr/l4prFN04FI2wOl2jX2OH/mSnrt5WmzawD5B74oRLUz6kQgr7OdXc
nbnR281L25nup4gjZhZGj1LKxcSr5SblgL6oHUM8UtBL2+SV5IkyP3CVzkUO
17qGjxkF6Hz/ovYBficqMt5HgwLcDXAlF3SgX2gS9E6ql/GRhD3u0mqdaLGY
00m3AiLAPXr0eRc/letKmhKNyz6upnNAZn9Pw/573iILZZrhu9VzTH/R0rlb
5hj5cTJRICJuS+zUudxUK+dBUpzgSM0oJvxDafKwEJ3Gz0FTm5VpWdaKH1ey
iD+D0sxVbJsNAjhnROWldEQAO0QOduzAL0Rnld5+EvQcld+ZUuD7nwvk/wjg
/3XlXwvlk15nm9M2U9l+115dOFxBt439VF6bafBdrkgMFUC60RyTLF9V1SWJ
F2H7joXl1zap+WeQUjdpr7kFehLiTHEp2+CcHcOjAix82wBJksYxxs7Wb51Q
HQd3dZpak66WevLj0farofOiJ3X/Dlg4u23WZDDWAOkPfwXRYnusGq6C86eY
bfCHLVBIzxVuGB+eqk1APrxtXdhWRYKObtDZoaZfxge5e63B2xqYQNCoit2K
D4K9cqMiP4wcyAUFiapq5c10ZCPNN83C6H5waBShw1vm9I+01jyOR9lCBIbf
KhBFwTK9XMPOAfrRN4gQPU+KPtk1uqQV71Bqxb3szXyEYYvxQiRcCMw5rtyd
PXwaM3FwtGSlMR/qtNs1Xfchh958C3H9Rb0BDxmoCFkefz5jYEPoAir3qtO3
yEXkPJPGUOKUAkaeyinQVvIftE4Vy6wh8Rx8Lvszs19xc+xDufhLaDkwwjyQ
SzdxBjcq+oDPTfYZ3unJT/XKv5cXSrDldebqqH7P12aJb6UC5IqTpI/CEQTW
XE6zzZ5SSsPULeoa9bEpFFPKHehjv66GWSPUiM+LBTVbxbWiFQh8jvrlBC2M
zU0nFtYZrdkazoSBfihIxIPzo16r5L+pKyqVLsiSJF1FX5LlvevWRRqLY6WI
G7F94R08D47WKPzAc+MwkQXOPBdMr9Mmc82U2ZOP3m+4GWh7ryvYQxCG39dL
wb1axKmLfS7fo56yAWyiAgjLUe0AQbHbs9b5nHNxtiicraqMF9YYLYkNobOV
i9Ji6CZTe9I/7EUu0xJxim32dG0NvPpVjN6eLs353xZ3jQ39Xv861fQVZF5Y
UV6sEa/Vshj/LDjz2kBtOXP8wSLzE9D+hZ7NQ2+nJPlbbyo7k6DC7A8bbuME
ImWATKjttAZjUljKCJ23qKWtJ2EkE3seuCAMafBTyCmw9UW0dlMNhsPEsRnI
+S6v/NV4hX0qf2pW8Eivsy4eeDEtTwgtU1oOWh3AQ5TGgckLuLDcdWZPrl/D
bH4QFcr98YZirXqBmCemo0f4u60EK9mNdPkxvsZIxl4w3f2aSaDbDNa7Ij/O
RbjvL8u52BGE1mG6EcYOy1RPRaYwkVNyOGkm9Pv7Sikl1a5WXozjpc5HC+Uy
9T9QGbGi/DIblnJ8dRdyMhw90I2S1c9t4pjoZ2AopC8Tp+vmXLDyvbAXnxO4
Q2km4oMTHSMgJouqoiZvV7m/mRGDUaavbXkdl/3rftwjfTJeRhENbG/opMxC
rePxYKkjfI+CTETiJVbhQnuX5fQX2IYNqHNtqGDVU9um7Qmg+V7i+bp4Aol4
bGz4Q7VSfK+wOz17JY/IvKdW+fkLDhZqv5/fe9pei2xMeDskfIBPy40WyKDR
gM6DvSAVOuBpc1yKHMELN6vnc04g/J+g3Dlw8XFLZiwwbqADEm85a/Gwc4+x
94lu1sBNE0z8s4hJ2Jrk493RBFatWyCPf0IoLPQ2prgzjL1jCRyUqKiueS8Y
dg0ZfGKa5KFVz85da1jyxaIy1mAWIR1I4GBwwruVLfHqZnGpOVbh95gZYRKh
NDBTkFA0JJ0q0T/V6X8r62GDpyqdZHYDH1gkNpfaRyh2iYMt1LtUiBJuWYgO
ZMvMEVdYBZvFzavvJQh7i+wnqapTV2nFZiWK5FpYR+hWnmVOVi73qIj1Q89t
gYC7A87jUywH8s8mp+EV7l96XNYif2oklzW0kbeAwsiCLxIgtcIe6Dao6iEb
pmap/+YXe1LsMxGM3CcDt2Qpnb08LOUSmZfI4vKgZQaU7THOaN8ZMp8vi/5t
+0HpHMZL2gPCv4kpj/J0H51T8BzQR1CY8VEyqRXA5UretaLQ3zANQautUCHf
QQKzY4CPG84ZELz7tNj91j3o0TuxEG/AL1mGv9wraWHAhnX2J9MqsYs4N09J
WWIZvguHpReWvuzKfZilj/vN6Ha89YTYuqHsCiby9mGxY7Q6GPs7+F6QZVJD
y4RIJFnFACi3OcajFtKObrlWFwBboGLuj/txt8e+bql12TZRolH6HizhP9Se
LCQyx8A0Qc49TUoimnxFkq7o5ytkoJj426KaB/6eS8PQU4jdOFDS8ACI0IT+
9+F9kM5tmTSv1KVkw/q+zSmFUB2SresJeUwU/1fLQ6NVYlMuQElvJCTwyw2Y
js4KvMidMtuWWEDZzy0sX2mGKjvOi1T67vZrXMGPS8CQXbGMD8IpKkgAIht0
2+zHykuISfllBK2DZ1VSRPxC6xiGj1sPHq5scoRCQONK2CToEyj2mpfYETmQ
5BDdzetvFvUe7/wXgap7XrVeXxKiD2xrL0lK5SKZKEMYw2oomXtT0WQ/bxP4
1PTpWrRsisrA9ZcbgcUXj041QeYN9fRxRjaFUiv7gyM/KnHAGto2BLSq2mID
rAFwmAItyixK6oA/6AAK0OAguzBWTl0xH+LR2WgjTTuFR+FZyTqGsBBJrI/N
0FTfNW8qkTfE76AtCeT97oQnselYCjRQs1khJl2SQxee5cK8AjZlUnMcJwWA
X3aVlQlVc+vnXxLZHBSeq2iBz1nS7+YZbadDazCJSoPFfsABXyjesapRwVyN
7IxfggGDh2RLXlCTExv6Qgnbb44EUNIwvKvmDjiNk6Yu1uxiQIgEyAIh3lJO
e0kqCfIZDDgT58ujGeIhGIzALUVBTCI/IXpG/7Oz30ls3HO3BguPCR7O26JS
oMrU0l43UcobMt/K1DTBWH8ywx+AzsVMvEWv9Gtg/289q1Oa2z5YNKIbkEaZ
Xj2KD/Mm8F9OBRUQE47IkDHagZJVBjLztnb2UoWLL+7WGE7yY3xEMdl2vS8S
1WxOyyfNEmUWqkHrdKGpiCwxV5a+z6uMLxQv0eb0ctMwNlEH3zleJC4MDVI6
dS/K9C00YnFm2IzvNbulVD5VEzfloLLLbfgOUbdIIZsk+1CT9uij96Q1bh0r
IriOlN9d5UMpqlnXfn+Uit24GYTFtNvhhXM8NTvW4EAmBXsVo5LYzNJV6irB
V/PkDyvufTQmGzgJsmRgwXq9XyrEj0DTEOW+TrC3enlyh7lH6tLlQ2xC+XvE
ojRTrpFUAds9Qc4kcS01+tIGZ9OjHX9lApWyLQgP4Car5X4Gd8qWbq3iVPVk
M4V5M/SKdVGhXt9Z8Q3YkosB07EnLItSclajFpTP/FRdB1zVxdjh4QIJrJSY
fX1OgtbeoJfw3xGMpH5hgsSFwU40YcPeugf5luOemDVzXWZwEDymkkEaOLr4
tsn6+9yCg1PuQhEDUxeixVUDPov3o0OBL4AUg81yzWWUMjRvGx8mFj4GA+YT
NqWZPA5jjgbQnf+zshi4N6dZ+rKIEz3HNm66f11sHO/sapdEjB+YZIa5+ctK
gpoPHqCkVUlEau/moC+VxGNpyD13MeQ2oYfv3oqlwlWZOelnf/uZ1uR0oqWD
AVgpY43SjQ3mVhD+S0iPMuDxUFl3bWSx91qv5VbOGjp94MTZiqfMeS6rqFlA
E7vSkl0Nl0naMPNkE8jgl9o/sRM5IaDh7Kk+b1i+gCZFgbJDGNVcQo9gzTzA
yubR0bC6kwbN3WseldNjbX7FRxdpaa6od4aSjkQkbI9ou4ZXDK6fGrZRbhPY
8hJOeRkwMdzrEj+7E83jGEF04re+QxhJOfvDlgne5sViiRbbAuJ6u/DLAs4/
bb+TBL92ja/8wanY9UYKF6hiJO/x4MaeespySu8Hk0Rweqd5JIye3M2MC+pC
arsh3qBW1OPNyqdz2KkcI/Mvml/u6mmVv3d/VCqT3H4+Fy1DnPPCzn0ezxr4
xBZX80Ojfk7sKcZxp9V23Nz8dSTmMVTRKlxuwvps7mLMSlxuY6RMNE+ovXXP
YR5y6INE03868INLZKjMMjzvD+60kAUqlNh07N8cV2/2J22vd4tLkti7by2v
LlJ7TZz7AQfRv0neXBTxu8YsZvLeagISCGZNIqGaT6lHB13NDTyvhdZuXslY
p9wg2slJetQqf+ynOtM7FHZhKOM8lRVWVW1ec/WTUCTbo5Nn9VzN3ZUq8MoO
pU7p54yjD1s+oM6QZ3oeOEywFOrTaLAFU6FdeAjmk6T/Ub6ZFldRYjGMOm7e
EiTFHv6PkCZOJ9QhiJ7xaxh8R/RnOPp4QGUkPQqo2LhEqqQKhfDhQSLE6KXw
ebakoGfgHIJb6hfjzUw4SQEdzbZxHo7Q8SmGfiATujYaijlfXtCB7wjYBY3e
A6oFxwubTV9K/75+50kB/Q88mv18fXL0j/UFYRnpkNLp9ZV0NIXW8z0vGpWI
p1PLwAzuT9htoVWl58Kh5vV/1c7pVj/qVV7ViyOWESU239iBIWJ8k8clN0Uy
uG0UNPgDT1/dsqLTYfkeEDA/hsNUljJHxlvcM4DcmnzreXKhIg1X1p2GY6nd
L8C2T+c97zvsrVvQHxeZ6xmF5cI5JcSklEIf+k+zeZHsS0zITL4BDbw+oGyY
VmPcmdw2zkaFdV6LQ8Uw6iW2hTBFwJ35Gi+BfxOhS4T8kF7nzhUPVihuut0i
RN9RG3rCOf/9keG4/HoSC+kuBHYEozJh8+ft8GN/tC5lq35fI4+YyLzYsBBH
sL4IIvZCIh46S+f7WL7UU5SogoiChxafBml/2iqgtH4zXERFFucwzoKad3g8
ob+JeiwbjyyfxZ8i+dpNwd/iWCswcjWxWkH9I6/1ikaWuseQdcpSihd9wc8Y
7bawPkkgsbpReiDz7u7NdG1XNq+7909UhftsFwylRCz268BYDAj2M0Oz/Lav
FQHCPMQNS5QZ8EfmWHTRPRUdqiSNtbzg6QEyBP6eAXFlZvCnezzrTF5O80dU
3DYa6s+MIl9vCmV08YhhYRz1g6WS2XBXtbiP6MPPVXQcweMKwZbKFVkaUzDb
suUaicHuDfbNtM7nyw+055ws4hUAwhNokxtghM7q1yfVZwBTE77VgZFtzYtI
FqgtWbQhMk/Q8iAz+9trabfH9oy+jA0H7OD4KdmPNHgXUal6jsKetay5GykG
XFn+9axFimro0p8nyExtU5+bKRrxllK1qmcdVApNrqjX+aX7Q1fSnOeGZQsz
sTxjTtmjkGhcZQgZheKf33aUzHAdLm1rVW7L2RfWwBnbj20+n+lllM4NHXas
QlOP7sioYPHF6INroSAWkOfpIe41Tt6hZ4L8J2yQehs+SgCaXVZRtGrAsCYJ
80MC9Qf7VB52VJUBTfh9QwjdibdoqYl6wbLxWvQ/WmsNs8ffbrIAugQ7zHig
2VJlPRBhtW0XOam3QtBdwDozoru32ImXBu8R9niYXKC4KcBpeaZQ+V0ppno0
oSW8P4maFkq/dGJqgAWSKi1Bn7I+I1rCnFz5WF1izdmwqsaawRFxdKVzTQFo
u+YPNYAHPlqa0dkIe+2rakxCX0IKtHmECQYyD4JxHdycx4eI/2LMFrj+z9rM
N+JvwITMh4CJsSmA/IVqFxFCe5wXr9sdnch0zYmQa8QkE6MTTy9FZjrmZ6Ht
CtujZcUALoaXzcbLkwNvrQ4TgJ8jXeYyz+PHFlmvl0Nllkg7ZHyL5YpI41O4
l7nczrF7DgvGnJgHbbp+R0OqREFF33fwxAQvznOJGYC6WRexSF4MQkOSSGKh
dX4PzirnZ86t+7IXYIvDBDz33inHZk9wBoUhSZNP418zCziAoUcFhowhPYCI
MZTJj7pgepyP06taz6C62lbXbciGkppYJMKrTyVJUw7tLh3HtT2RopYEC+Ai
9o5FyOgnII2lYtoGtXffQgDXiYJz1DkfuMYg/k+/tzB5XI9oeYK79ZOiBFjK
xV6QS9joE0q2unQis/fqrj3uKZmTjNPcw3eZf1sDFEjxPojq0lIhyLPIAbun
NDDkBE1k1l5/vU237ih+KrTzfbW+3eamdkmc1VqZB/dicOq8HndjO7jJ+04/
PTGaQuPD7PshpevgMIdHD1vcOy1TiOjr6+c0tzvG1CZJThVU6bp2mI/d13rX
jIUphadN/SCTJy3uuinZOVUhPNnxdHbZ/2rJDRoJeoIcS86BwZPfYddaTdN4
Ux8KGihHkElqGa/gBnww+H1brN+Fz5cuE3BCQNXkXBBj874GlRllJWCb7UCH
JDaORmCHsEoqy4eGWnzA9doqEvYdrDpCgKICMFrNaJK2RenV9ZeLiw/cuz/g
7TdG54bHbB/jipZoJVKkgA90LUuiEB/QvCHS7ns7b1lxz2yv6w9Z1QkLmJIJ
kUVCRTi81LIxTb9lMTNV6Bm1AuU3Qa92VAEVDpriLi8//W/TN7UjyNJ2ur4r
1ysXYXhCFqe32t3ezZ1bNctVxSC74bfWFtJgPVdQ6gWqUgFduvw3jvpBqQhU
BnjXOH8xet+NOu3Lv8eVd07yZHBDD6JWdE8ojN0r26HIuFsNOyEMZBDeeHb8
Br8G5P8dH4UY1fa1iMzXNm5x7giwk8STtBci9juJiWv6j24xXiXytFWhGlKy
9OgZSYbbWda8HlvsgjYhyMHZr4Mx7nu+Z76jypcIyU6xusToG1dYnkvRsG44
QIv0iBPkJ862MVO5W+CDe6YgEUXcRdzcGLlcBUCaWCTe/7RXCj7V7nupy/mS
HwvPMr4HA2DEXcZ2yRfm5Q566UslH9fH2NzW5uhVDZHYuepQNVQ+t1cLEeIq
jE5xyM9dtmBKCgrZ8w+KJXGSUyLZpSmp6WS+w08U84TQEcdUAQlsjnTkENtB
MVXMNnr/v3+nwWI/oMGaKQf7use0TBZXFA8M8FFKoPqvTYxiMWZ7yXCwQpuP
DP6u6aIt94+U4npZzxgIF35ecIFTTx4LqG9s28bbW0k7W5UZBpMYFd/CU/Dw
XO+t5GkEQ8HhgrWBigH4ITmB7tlOhqH2ErtImJ47bd46m+fFoZHQjqdVn4Z4
jvpUxLCTVEo3MbPhQ/mVo7KgGH8FsylkGYMw9YxpHhSqhiDthSQ9ABI1Tb8m
pdd34LRX4twXo/dDpGuGZ7RUfm3yAxS0AM+UkQ32Zg3LmyVo1XgiEJTK4HH1
he7zeJCwK5v8+ITOSA+p3LhWW+HADNOovo7OtAPUN74X1D4VukpyBwutUrs7
Z3q+9O22BvoV5vjo2Je4Y9ypTYuWjKSEHUjBtohLOesdam7tESA7ckLaNr7C
CaXS9LWFLIaLpcfRD2kBYDA7rPIAjl9uTelsXVqdOBH/u5lQFyzrsM/ys8fI
L21tZsz0Hr8M8zPMdW11WUxIJc2Sr2a+RD7lwDrgrozfFHVqlKxXbG03dJxV
M7QArEUYEAcB6w3fkGzmzwjDj6K6ow88lQUuUOBW9i3ox8AgLXhaEowj08XX
RVvFYBA+7JLu6Dzyw9BRK2MBnRKeCBkrNwfLplVfl+Rjohm/tvMZ7cOLMBzt
acqS9WKOS5UPdBMU1WfzskQgblATOAqOYyp/KtFalFYrhW0ZBosseFeKJ0r5
GipG22RLUAVbiIiXjq+loKxyn11KPE9rII8gqyAjKoreohgoKXOX4Y4Pk/lO
ElPjJ7lPNQJgNOJUOg+YEpCyfPJMlWYYKkSL8Btk3WHK+EJnOmUaRUtHtmGt
6F79AMLiEbQbwwTpD1hFR1fKBwVh3KI8Mr2jaTwn+ogNPWj8RIfqIVQKYf3V
cCA1zTUgQdasF9jJA0of9uM9Vx94kwpOZkJgp3ODLfIwRITxxOcIB2Pi6eYC
jcGJopaDzSk9jtLSOysyyB6Nw5YerH8kIjnNBKwKAqcL4jsj6gZS7nyxSWxf
S2imsxum2KGOiEeQfTrP9nDbL04+aT2lWKjS+83gWX3PUNwHRomd17vILFd3
32A2BzqiIU0nvFreiu9SVoTEFghJbaCmw7AZPVLemjXPbV+820Xetc2LamqZ
az+PjrxdPwhmWDC39bHKrXBcGJP8XKX3M43TwF1eObC0D0j4fjSkifNYi4fm
CDXWo5+9ynmtrxRFvE9ZkhKeSWjhuL0g4DO9P0lEzbjxIVwxMCMmaWamZ2r0
909Lf8uTBxk4YxyKouzAKT2VBuX7mud00y5xcJoCVNAgTU3rQTGhlF0ezITT
xgT/VnVl/Fna18AlEbwFry5ya+q7PjWhmAF4GK05WJCDtmBzOw6KVV+2cFRB
hd80mik4EhXqAcaxrQlLJ54es/l6i4TPv2Kc0uy3Tawxo7svqVjyIFAd5ty9
UPUiRTk9V+xoJd78IaBDP1a1AjWRewdYCnBEM3M2FOYNR+2bD9L5m3z92Y2v
zf7GeHEMEntZtCRQ2QCjZSQHdsllGDOLl0DAbuA4f6L+7DPC9oYO634syJP0
H+2TX5JyUBHg4oZkXVfJwi5G1witI8zY4esLELPa9S7I8Ma91Y5dwh1ApEst
3gPUCg7QPNguRSshYOo9lrk+EGpae3IJYRSy733taDB4lcjyNEvy7ot6oKCZ
HsxNJ3jShOZpZyMB6pnymz4ORNj+gF5UWmr5yNTfRiTbdvj9WpGBtSTtAWwv
99l2kAxFlWMj5j/oMwslCk3/Kv/VPN8xgyw2PYw74Gi6aspLyUERmXHf11T8
4n0sQ4cViBjL/4Tnm7snoi41rX5ocMpvRznEvrF+ND3FGSRLcq2cPrUZ1aL/
Xrva8KXzrKHeWruIguCAUCCGWKLBfNZG3QlIAhi/WReAP8xG4bmVMU47X89F
nseT9lyhsZvJwUXF4t0YDABDvgnZUcWzLaeMZp/mtx8MOMJqa01MHClPx4ja
qmA41ScOCNDrMFrkqGKcXJEVfDJlYrHcFBThMASwd9fE5WjiDj2Yj9P7zRYT
B5MkiVDUO4NjpCK92xDNo/FJpEifJ8DW6ooprl6V/qq4VucSG/kfDGhKu/fZ
hw2VKYFUeVOie8TLqlRSfq1LEJ+lI7bPiMLGoA7sPg7q3yIEWou6wsFy++Pc
juk62viEh97yHyEi2xSDoFwftEVMIFmpwoHAR3dk49VNpYa55/Q2Q2qtX4bl
3CxQ8tU0KbCExhXZ+YTv5tvX/W9hHKxyGetjpVCsy1NV4XqiNW5qXr1GF7ad
19td+nVf/rUUY1A2nm8CGk1SBgY+v7LFserGxqkRzz1Ypl0AUjweGppUcZUW
79a4P2EKJHjHb+Mv3vUs97/XyIByrRt9rRuI1JYxhblQF/cOzq0Ly3nG7hzF
udyS+BwpJ8Ta24R2aqXy2z9iSwrnY8j3CIsjAwp5L6B23MRNrimup82UIZXA
UbndbmKC9eA2LpDT2XnH8oenssZHEPooS2TN3o2cjWIMa+wKT/H9o+9JbaNf
u9r+sO3IX8nMaLRD0KYs/SOlqITGOQq7LQ1dt2nHEVP90eqqdnbLuZQOuOzM
gU+EhTeEKpIjbNx7+Z+QOrfaNYSMatnPnUp3PM61mSYKhOgE+1Szh0sC2VO+
9scfXh+/TBthoZegEHmN86TDfCgJAyxFUqIM+3uvq5ir+zI09A/QXj/AdGIk
PX+3FE4cs+Bz9CIMYVJHA+NZxtD/+6VsqVYhGtlaQCzVuSzjYyfaqWxVKnUj
hHonLzeVueg+sU0dvwe6NxyQQAs/4kX4Vw3HyrP3yEZthm8g3MwweUdythCz
awAbJGaJdNU8jbX9hmmCQKLPDHSokY6ZF7+DAyU880xKk5e/UAp/lk+NTlRj
EAMVEliFB0i1pdR6AXFORLyK6modHdlcc8clNJhQkNSBGly8+qmQQXNXZv3y
5XzkPDWsMi3RRv9RaACX70hxMMuCIjM6HynfNxleKgMXJ4vKgBNVplGBAt/X
iga3RjfS0T0DujL/T+efsuLT3EpdKrz6WFxdwamO4z8Al3rFsM4jd8nRFT/R
E7NRpvkS8g41vNjkqFPGx8LHfuK2beQCRhx1yII79/5glygAo+Rn7EsZU9B7
CFcU15fBgnIgyTDStbjO+KEK8+KK6EVGNChQSeL3AKxS4MtSS4u+n+wCkRPC
zv8dRra+9JS4/NNG51Pt92htKvorl1Mp5/5uohSl3aOSmelo63xwyOura24u
rC2uO7WpTO+qHKsd6SyFAZUlCtAhucc+iPNF0qt2VAYWGkQl87X/BHJB4sST
mAz8Ru0YcFvUa+Du+l8COViSk7QolVBWD9iMF40RuRLnBDwjY+rook+93AOq
lE70M1Ky7rsVGHULIi7O6yka1FDkI06uvdyEcs34ZIvYCTVXahgmOjjxv4XJ
QO8axrrnsPPmGUr74ky0yAuRZHmCjyPjIjsbF1bz3aWE+Ja3V+n0WmdysNLp
b49yfpN++oR7kQWMQlEsCSMfG16lTdNVSkmMg8DxqEzB4HUev16DzP1hQvHA
P97YNX60++yVtPRPtzXZhdIp4pKaim3PmyR7r/dsTupO0yfrH3B7msIIDnmY
DZEgoiQsp3YunCraeCk3GunnpQBfwbNBJUpsgEU07b1RpMRh8gvdS48ZBwpE
tKIlXcomafal93mdcW0uflQA0/2tkMH0tC06p7Se1aVp/9RdKeE3icyQCrNk
NKa1Diy5cS9weKVQr6/bp4BUcAMDTdFbCREBTVqb5gSdiVIgi2OMkUlY+glp
AYV15AZEFvCa7vldufw/YJ+OaS2cDP+MWrthVYzFsc1RmxP7aQJgUnxnmFZY
v7iajmvilAAxQczOWtCn9m/lyOS+kIicpBnw26kg0hJ4tkL5TK0RUDODAoNZ
FhBIV0q2uQS+e5F1osBSeVCACXM1mDWU3nI1dACLEvgbz3giFN5e1qIHns2s
d08dGfpFkYWIPCM43zGoBLZjbliuDCo9Efj9ip0B0AiP5tA3Djfot8STMgXz
/UXBuy9lJFgNraE3D6CZ4syHVntL/9Ts4FduCA5SXO3oZvBrPJMJnbNk6Jd+
5CoknlOqwY+O3WzNvbVHc6BHGcsQ1j3/wo3EA5RTgUu53q4SkK3itlyGRgHc
rfHwsGtsY0VXU95Vj8HEVIGZqYmesd2duqENSOkliEnWLxJ604arytbaq9Ua
x/M0SwD+Xsa2YkwqgRLWx/g4Q7hjVmEaZ3f/3BBjV7qAXtUwsRFXD/0J1NCt
zeR71pvPdGz+lFnxaj3+PGw72jTIjS/wqIZRGLOgArlw9WlI8NAi8VGtfiej
gG7Ql+hyvQsP9mQ9LtXYdsfvGKN446mUclYUH90eBvEVN27pEWyUlGUOeKTe
rcVDyKh4Ru1ziwuW+t/oXgAIrd1XhNPKC7HYNHVXjuAETEq6mjoCIO9lXhNs
pirKhcHsZstOmCKdIypB4XsLxUslu+m7LBaITt85YKi0I0fYo70NK3TIQXWV
DSVzN2Mqk3GuguDmlwfILiuikjcaWTWR3Je29uPcvTGCV6ee/JcPx9j5yu9C
Ij0/UEWqGsBn+9m7ZJpx3Lchf2d/hj1g8G6Lqm4oVtse0ZszvHu7C8HlSw6Z
tORuwvik3gLpw3OXlpeVHHlq4vvhvx5CE+fHru1X9y3omy2zuDRjiCoJUbhQ
yOo4/AK3L8iTAtruvkcsim/LDBhAlWUT8J2syP8morcffYODsDpatzn08gAg
9FwaGACciaOq0mhEOKkIJe6A3yJcbBam0PEIJsqPQn4C15jgSVRW/QIBppNa
LhfAAEumB1ePFuKi1sWNOs/UIOJHQT8wGrkSvD8m9dkt52ArJRiCUwJ9ZveY
BUgJLu2gSCXK22LrhpzzYtBJnzZAbDHZm5n23bS8ytdEvQzqCUELRDqJzzu6
4CnFKfMx5zNZiae3StOxJzFI/9ALA0etd37+IM+5lwWSkdYxfYwmwiv0wWOK
kqmcXk1ePr2tkllqgob97XesKD9TSVtWE//fzF4pQvAVktYqSmVu9ZI/gTXk
HDfsM/PiSrleML4xSH+4H7ZOltc7FxwvRCLs82WZ29q75+9WxgI1QlhhG97y
Cl9vOo8O0f3SsKiaFePwgUoqFKXVM6vzJsC1yI60h07m5DTYJfPCigc9hLkq
Pa34pyTOfF1PwqZw6V2XvDIumL++HE0KgeJIgkvLbsgMtSJ1Ux4KsU4iA6A0
GPBf7eC4WYYtFuK7hbhTsQnf+3GB2t+LQfIgCtp0CHRzZHG1kknrfhkn4rQc
RnJdB2/lHWvi2tkLldVb/uOnGU0cXHOmFrxCNPkHxEK6gBG40LB0NdvJCvZV
oJ4/1G+hzn0JUug+6YsRFQx7TDjMqRNW1c+i8n8X3/ftUCQImdt5Y5G9b9by
4S9mUlXvqBLcXovvu8dLepGLmsU77fjuP4FjjQTa8NVZ7EC4vKBHNGEfwsKn
kKRhAflSg36rdX6f96JhEcLPxj0eSUd7vMoXeehRtIAatuvRGxxZ08Pbe7et
WiRxW4s084AA7JWxxUWg+1N8jKKIVCsAzttujCCNYsor3YUm4ZSWIM32Iejd
J1IaOYmP/0khV2EvmTOvZ08Rcxo8crfZzPKcbcgOYu72UB8ECDJ0ZXDPTGcj
ZrFozkahSNg7QzsrJVefYoUsJ8M6SBSf7toO6Zm7uYGe1Tr26iN9aELmsAX8
tdxEhT35tocQu0CFrKzx457pU2nzFwvyZPK2wlkkxHqllFaOZ8wCGVRrJAAg
/46SspGEVow8YCj94qZTocfIK0/ABpwd4C4aSteLZ8VlpfmOCNEHQ6BDqAGX
qh4iiFf8OSNsMDhLYTTVcsJ9c7QTmuKGwlLoTGJb0FzyNzN2SU8F3AO49CE5
xAB5jcT8OH35tPDRf/pmcDpgYHUf8CWgPU5SGbritd382EiitGePErViSwYw
/dKCzQUwbP/E05tyodWtckxXLGLbdDuVybBOU/qAQuP/uciu5HNInTGYtbFZ
HJC0qX6ABAARliqMrVvvLU2F2qzRup5pu13AXMYUVwl8Uq9khTsoaNWJI8HW
7Xm0cadIC61m4k8AQ5Db3Oq+LDOB4y/mlyIrGAp71zNw/4d5qHfWK/Rolvu3
N+3WS/jVJlGW5c/2pcvVhCi+8sMVhduK3P/zX9DPZK7RCDaDv+qe0M37yBEm
cqG9MOpG6OvvUE5V69+0I5mh1oHxV+IcPUuqR/DulyoEYx0htyiB0xKq8amk
gnS18RnZzwjucqC7IsQ58E+Jl8Xj82AkiYn2IRSfhnd9BBWRU1Ni5moqct5l
Ibx0JIgOoEbyL/yGmTZmz2lVQ+513PAcRyhg3vtBFfx/RJB+yWui63uI3CjP
p9oDl2pQeRByQZ4+LzOePS9BDRYvGahiB/R/syfGd9fWeiZF/1F+ufriUs0Q
WbyN0pq2y4Vlx2F4YhnNgDy7JOpsJ6WFG8c1Zlf+D6pm+FO08NbRDPYtKuLJ
TVFYWCzBreHy3tWLNnKWK1Lvd9er4boSjTvmjsPuJYWj+nUdzS1iRPzg5qGy
boB4esg015YSx+YusII7FPpZzI08N7AuWS+XQFtCUGKpxdL58D6L0W8LrS/D
34SEIy+u0Jif4qRw0MQbZVCxfcYAb3NAlrrfUns+JK8qwG1zLaQdumWRIOiH
Cky5pbQqF2FymCTdqxCpbN15vXu02zg/NjLKI2SQXQLksLnT4ZiziLiIi0to
Myw2m0GjLq9eCCMx8dFP5aWfXsRjs5b/v/88JKnH7hW5Sasp/L/rP9T1CO5R
qLyjOYfunRE3+KLJ9MC4WDRjsHe+EN7lGzt8oLU1+NzfGbQwer7/lDrh+TNw
GTf1iEDh/+Bpe/6kYeC73+TlCNyGsEOW2HnxwjAUHdkEFfPudQqO8dGavSuW
/s16/vvKMRAMp/TzQ8oe1hPIwSj6QU6dDhRt3lcLCbngnjXGDsyfrcY+atoN
OMc6OXopKIHrJjSDAk7A/1Z+WW9bqWtoUB69b0/OR8oeAd6OeLUzNS71p0fI
HppsEGSvMaT0mjFEtZZiWuGVpW3Mj4Jn4XbgDDHZSCDdOG67VTYyvCZOHtxb
7S/LU+nB+vp8L3uQxBskV9TOQjui2zMpk2KOFkR5uTj4UKbAxBjTWHGnMKuK
56i+iBuXhQB3XuS6TJtimoa+lb9NXZ2Bn9wUngqOoYTN7tOkScU3CB6A5uSF
j/jTNXFNJFwC4JWdL0PGN69lJhb+WqUJBIgkX1KKd+maBvibsqtvbwTGVbzX
tqahWJHQ36+AV1MxsJ39kY2g+Q5W4pEBrxO8ph3ZgvyhXlB48EiOSmJvluRJ
7Ea5AfgX8T/+sOc3SkSU/qVidX5COkyOeNH/CMRI+wZ5s+vEDyRpcrerK8pJ
HoDUY9je/Uep8q8e3VDOPHhtZT0lT58tXnUD5adRMpznLqdAQlk+dsy/VUPY
AzvDdeCToGeVND+POx/P/LH6BUPeWCJTbT2aeFUTzgIonmJ9w49gn7jLu4cV
s+dYUU50XKB0N+PewgS3rnbmHG2wF6F4wiODGM295jNESbDTXDZ0zeFLBrwm
1aEEQ8TYhU7L+mpxBhdWnacBhBtkGPsBASTfaH/WxLrAJMVELPbbTgw41Wb9
ORptlYuuwPzScqwccB8wZ0zSS2sFac/Olb8BL0VaE7Bbw5POKP+AoV0BXPz9
GSeUVjvxcx2EChtBHspB1CI3xAl+BXwKkGqtZi/KybnAzRjzY4qNdwLFIxvF
Urc9KgW27wFUJ5gULVdBlTUsTRpHU3lYR1M0hSM6H1o9P+mMIeixe/n5geGV
3dH/RO0DwWknvwo+aQQ3BHjpHDB9whChmyLgwEfBcwKDS68cTHT5NQf1RoxS
Zr1wFk84VG8hC8O7Lua2j9xNmrd2PQWHXI5AbCQ5KvpwXTDPQvjwot1n8QvG
kKuCgf134xOL0jATTK9Y9mTJyRdRO3IlLjA2XgwCjp+0SRer9poRV6cO+IoP
IWxdkz5j7kNWeKt3VQmUdve2LhcOyH2nIqHjUlWqz+J3R6GKnPhfxnCSQSuP
eBJ4y2jum4f+IofLDnA3zHO1CHd0GwOrM2lNPi79xxR0eo5Fc4XhucJEqXXb
EgFugvMUraUHaMCGG+r6PQqktIdrd+L/+5SCKMDxLxKgjEWz4jXEcmbrJBkU
J8QcTpOqLhruifTq/VQ0D2leB8V8il2Iaog9qHLq2Vuv5B+oqG3kbXDMcAF3
uY/ise5K3R7txnkQqCpF7JX6PRSUmPlLczai/afKEbtmkktZswr8Q0SC8hN1
quDrg/4Uy2Xu1nvf0GrCkDq1qbZ68fvTCFm5RpZyTz2l5w0H3Rzc7Yd3mJIh
9dgdGUyzDBzKF6QhoXoxGAJttatNDnokvOp1pUeHAjQQGjV/BgRENj2RR33t
hpet7d54OX82FV5I7kSH/m4G3P2nOlo/fAdk4RyL0fEqzaWpzI7XDX0TNxxq
mNHkt4fpB9UKSbBzGPllR0VuQ7BJ2CRRIDaAIFhP7pM8JFuyzhR3yYXbBOGQ
KRaVlRs8vODtFdrOWsO17voSjilY5cYT/XcnlO2ZHeHbe1Hf3S4c8RNa3S0v
XPqfKFabSOdKJ3B0rJP72Xwde+ndFNd+sxVI34CJzwrtEKuxX78fnW2S4Xw+
vTKR82LWdaT1q5GuUSOy6ic4Mh03LNwUTxpfimXy9scobBW2P0QuTuB1IsKl
J5INHURZJ7e4gpQi74lODEg5NqpoasSO2LMXM4Lfzjs1dgJq0ytf8amIet1p
EgVAbUUrZ8ffJ/LfJUTqXnIDPQP+5OGQ1FFeYcJiwU5pDlhokERUaIgshei4
3lwLi14/3WNDSGzb6nYbYspMVjku3UTimmFlBeANams9qtjTWI6k9B6KJ6vo
h3RkeJzR4kfRG1W/Fxl/m3s+EU3MoJHQ7dAY99mHqEKhv1/Gt1L0dKR0bYPT
ozh8wL/DlDk56Zgjqf2k9v7jgW1+rcxZdibqYwt22XmwsfX1KTSE0VN26QA3
HzINozYrNXybe+a9ag22S5vyMYEgtkfHPfBFP7T2KQ9tfK7VLhgghVTuQdhZ
kxjOdw4E0XkM9qLT0gz5rYbONFLX6kYOArjHgD1GuMWWd/kVWKqvbRHlWo3Q
QaC3LJXFQIyBXan3lYbhNY7Tv9YWlT4fHfWou5DfnkLNsE8AllwiB0+w70RU
DHwSTzNQTgL3b3nvwjrsguZdp5D9t8LLrEx7BHvu9TTPK1d/nbt6vvo81cY/
sSEOmdpsUQ2C9Gsj6W/DIR5+9pq6kiKXA2r7t490n0DSKQZOq1LmXRR9NB04
KW8OBdbPdK+10EyAIHl4iKSMnHGqPL2c+CyGJBNpI2yc+H8vg2wqKMFqjKJd
D+xeUUGTjzFglcbndAwwe49UmR4MqR4uxnHVXuzqdcpxXhEDSGzvCplmTuE1
J44zhzPbiFYmDdPRxgaSOg0vjMmrXn4npKYT3Wiqt4jZp8X/Ibni4PjKS3ES
3x6iVWkjAC984yqGR/s3c/zAWgM3vJcI/1n5dQCwTsEJYtGHiW3FtR3LafU+
FjWvEr6s142MXzyYI1hhBYw5yGKYcW9wVtWvSq98do450W2fJ+0goFst3xqM
gtuPExcJZbzTKiQsZw2kM3ZBrcU+4xNIoKbQSNNu+G/9uyNfBglHxyBdLShY
Q4e5jFAMCieuajxyNYkn3JiJpHvtUx5b844zgGJ94H2TQElsLQvsGuZQPlv3
Y72686UMJsKrpvw40lkWfna/QtQxJPldzQJlIBcDT4a+ajzawjHllu5LsEO8
tDTfqlKQ21nY+3XUeIACmjq6vqzQg1vGiK2BD1uz61SfV20P9FOHEDLKcfNn
qKlXT3Hxy4gb+ZNJYSRJlOnE3hfCnxEmARm1hb5opKYqGgCo9VXTc8le4zEI
HRkfz//wbVU+HzjNQFOcm1wqZkbVXZb29iB8MbgxQGKZGk5Pv/uiKEaoQCIP
GxSgJoHYAfjpQeQZzrep5Fh754TGuLlkwqz9GTE1AQQDvBTMMLLl+9KkLEJi
TltcwiHeOKik2URN2NKfedgid1hQ7QckGJC2mGGRvDSSFLcy2MmiBBuenjbL
iDsdfJZDhtpdMz2Pw/17VD2cFN+9NhGqKVH8UXxl5R4V4rapeUeRdrmTsJsn
In9gcJGZzlk31CLlBsni2BO+30qqS2ZpYNvDXJVXkwMrCUNXh7XmerLgh1sM
NTGWTBlmKooEoHVFySxnblLv69uoI6/cHgNXiGlCRQ/lbd+X9TmL8ZF1KJJ0
lF1Fs8oRm8S69QmN08IVKNivaL0Mku6i/LgpGSe2ZqEZw9DcoocGEBv9bFXv
O4ln1+TnlINd9Ojnj4BBA+VkoVtPGbmId/Wg521nr+rad/pNNaBlLHgmVuR+
r/bZQ4fBq+BG0jWJPRRsPBF07XU6jNkNOjkNdB7M9h/SqoKc3pJ269ptQFxJ
B0m3yNA4TVLHnpD0fzsE3cf+fHOhV5xntydGo4XiAUj8qr89SkQA1U/DrTwT
shY7lunUCidYnrHfNtu4+9ysg0vpwMI0gg8cMhbpgesJ2QKX8RnYTE4IOg3Q
It2Un33lAwgh+gqfj81XpCZBokfxIn6QTt8Re5A0Q3pfH3H6+oI4jRSnk2M6
rTPkdCbtD9qYu059obA6Ut41YeqVtLSZ7DcG4FwynTi7yXOL5VHspK74iH0S
Vn+9gc7Dw1VoMwQug9s0tVsYbqr8Kv+RWMaC81J8IkKlnyiA9dmUl+TanD4I
VowOM1lt7SYlhaBuec+0z7DVyFVMGKp9mExW6zDNnScdmOB1mG2hkw2WrKGA
EdBtSEomeKzo6ZqGZmvQx/WMs4rY12mGW74XZCV6PmyqXzGS3jnFHsQ0pzEW
8N8gW+aL5wVD/87OEC90Vq7TJ1NcV+fsGV8wpH+RmRbm7WY90OPW41N26jLY
a6Z+BWNtVv3cTuw7/Fb2SVQHaQYCTSBLp92ew9cNZgDq7hKpaxvjQuVQQN8e
HRRoOqK4wpQ3jJ+HoggyDOqTx7GgdiyXXdw5cLtxX0C/Ssn/vX1pV0Xg0BOl
v0+NqotSQoGyw/IfxvcUk15nnrF8J5mGSaBt2WyYqQO1dy/IxKxfje4m0mWZ
LucI39AekKK6eaM6KBjexulG+nzlSf5J03IQqCUSmIZVqzsKNL1Yx4XlQLt9
udR1UnXnKekBRzMQx8Z5pC1quRdqPCWmCC9BQOgHi1M1bHWpCP/3zOEzGwzy
VZRonmH4LwXkNKxIPcOT3YeCPBoDFpHH/1PW1E9c+E79JvHsByZH4jH/glLd
l7mafGds2NXGTHUMXOu6S2nFzgHkPySoHH/406qriAd3MTflbmq5NN708iWc
4nmNglMbth0bsDL+F+aRQ9Yka7jhZnHaRTxBgbyJybptoeyaznGOroWypXJU
JDpu6zwtLbntZr5SsLjb2HqHL+C8AO2Fhah6hK1p2p9BX8wZGurQ+xTlUQ/u
tLtfm4MuwiMWRKZOI0paPe0BoTFX8DhV8jHGnbQ6xuw4txKj1x+AmscCr3j5
0wWlxPpc0JbSXNIqojVER0vz7SbJIioD18pHl0axYKznCkpV+w4WV7ZwMMEL
vi+uopOddiL+HeYhNpgosuRvWHunLUSduGY86Q2Eu7hrkoDH+e/Olec+mvJa
9f2Xq2IZy1lmlSWgZq4u09V1yWeaNLdqcALFSyFFVKdCsyYl9HAkoBU/pe+p
BOVD4OTGG5eOxQooTg5YIsGIijzEN9Wx8QJRW9f41DmyhvWOv8t9P5aLZjb8
2mwxPxz2mHtpkpRIqr0pvwHd/9vLTeYMO6taaj5gMd2pD0l1C5nB9tSqAqq7
vbG3toCZuCifKflXZ+ttbZz6aWQRmTi5zQINo/XTa+O/ga8wZLDnJHaOxNF5
O/Gad61rshVCG2CtuorEzDAZ10qHaCb+rqG9eDrfbJtAp6UEd0bU5iOuESuj
XUQr14fbE7s5yz8NwBFTFr0xfYRUrmkqhit0spFTSNRGgno6KM7yW7KzyUB7
PDRZtdB62Nvufuz9I9HzidPWv86QW3XMHbIh6K02fvmecmTtNscLGRzhhg8f
iPRJ7wohqfKcXeifOeEjBDmla9OU52KG0gdPQkAYNwoY8fHdymcf1gyBiiEa
LdvdbdONfckoUAOWbPBtysoUWDww/xPbawf9k5Vsts7uLTlKaCEeR2jHyK7u
IobmK+tvjFnqsucOACJ8AnE1nl+mWBMYaux+oGb+SxJWJlABfRq3Qep59nWQ
jp1BiwHtg2fvRwvTnrbBiow8dLhZ2EW9n69qPc8c3p3wVbNQvEQkN9/3r1zk
QqvUD3j5Qw1bDvTDOabMaKt3DrO5n2whLITflWh+oSrNc96N2nQ1Ti9OsYwn
mabsfNZY2T6W1F2WfB36PZ8w6l2iug//eGoLlA3XtH8WIcdz5GGkKu1Wu9TN
p2BQjM/BNWYDZMh6xBfgiF1NafIDDCGE8mlvTLlR64NVWDzofR9SQqEC9zgo
G6U7ZVEkD5l85zNVw9sPnQLqSN55M3ZwuSsdH9/IxVn8o253ssmKizdO9bjq
2RjCsimzaPEF8dREnaxdL+Fkt/GMJ5wcHPXNLHa5CSw+kBV0DuXHb5v2QMKF
kmP4L/3qKIsDI/8/fHBN5tqowjw7FeADaDUarelZmwQ78BsfrGxbFaGNMbl2
Hth78a3r3/+MadvI2RtDTRDyNdJLXBR8RL/z3QkJORQXChcQERgZELzIHnAp
v6isIq0rfdviD9jb1IdymXmW2eBOZDh+d9O5DaIisSr5xOwFHfZ8GhGwKCtL
Pyz59ytFQylGrCekojrRiN4BKmM/RszzCJ36N4F/cXUSE2SXW51Sijt6hFxj
fgnFKCJRsnTpZtwzz4nn4RN+n297wnSskrXqV4+e5KumEXpS7olLzJo1XVOy
BmKyI5WQMsVTlz+ybMQ9uICEJIJl4jkADRRWF/i4xfwloes37roLrmKtAJXF
p+4Q+xEFpw/jkwZiPU+YUlVnLfXslMJPMN9K8hRTWLynsV1fifTSzvn0YCrj
bMvd0ioIhsgw/3OU4hHZPtP3a8CGq7S/olk6WTkjOLsW/Qu0m0g8HTndqjje
cwl3MlfOKHDnOy6yChVnsuTuEts5sCOm61T5kVD5nnESjBodoviXQtqVyTQs
YUxnI2Ar8k2RsCVCLSSe1/15AERwvsk02OWjdqtLPkvzEmXKjbT1Le67zUZ1
VHlt/XeFs525XxcV6RPHAWzl3pPA2W6dC5A6mPPp3Gj8Hqoxx6uVX7bQMsAU
XXhtYaL8l0MwHNnAi6rq15Jdaejrjjc3oDVMMmYsgmm4F3j4apNvhXivZrnQ
UkQkf3bBDM730+YIvCmKTkXZCNYaclmEtTLkGi/DUM06pm+QNunKhBJhunvg
UbSIFU9s2oRLOq+Q0NVYyT4gLuF4j8Tj2+YbwlW22ryTKUAtcMuz+bIMc2F3
D+b/yQVj96BrL0SG/Lg3E4g3mt4E/MOLioB0Eme0I48XDeHFCnNd2SfFXOVX
LsYnTESRQPgZV0d4b/NWlmfyfMQwhmfQ82XOLzUicEGgJwhmBqs/tksSDxgn
dQI6f1TXubVedF6hcBd9knZcXpexJbqFEAxYCn2n4mfUfMBNfAn9XkkX9OQP
s0ET6EJKCfZlecs6RWVGfqyIz0EvjSfsK1T4094zSpgdMhJ8cFeyOA6a8Qgb
TaKhmCe3o8W1Wk+M+gi9othknDkzvYl9v6IGo+Icq1A35v0FR7diB2jyV11+
9zwoLj7t76EK87PAZ3jqgu3tQ1NwyzbodC60kZLlf7DlVfYRavasJ1gdQxEQ
rCyTdLynKJSmuMrGUGKd/WAMgU8Va/LC9aFMvc2MosTfWzQnLC1jQoOQ4oR3
y6Tunnay7YbI5BHqRNtjJQi5GkQTgZs7nF/nN4bhjBAq+UUczUx78gmK+5pT
VRG9PBnLu4zX9vRJQEJpBVyEujMTxGXc9vg+L9rYgZAe38PZf7LRHSNdaf5s
s/29mQde2u32gUpj90d5nGCufVEaHq4M2a30xq9ojTdAewG/WQQS8muP8JbU
aDh2QO2mXxzSaIICy3W6DhWWgBp3f/9qH1oBsBEGbkf8k66aV+OwcTmiO1+e
O387qRtnzeaVCRp2OO4MYyO6Q8nB0WOcEOh9bpVZ6Xz/RuMTDWMiS4VOq3VC
Pi4ID61o/FbL9o8WDy01H+uoSp87VhQkqyeJSD+P57PBda1T33SG0dsW+2OU
oEtknusSIhEpzuCKsynXsRrEebKwQNySUwGFBiSFiSD3vUHnu34k2fws+8TH
n5SGtyjzRNoCulJZC6KR7TJzmKHC85XXDXcsibfQjhWwZFlH3gtTCg8UVL6Z
FGACNq9z2mzMTEBva3tvpz+spyxBdHSPK872saJYHGc4EmkWsUjYWYKcPuHu
YVWHwjDTkSEg6IlmEggGaClCv5gJ8q6Fmplc9GK7ciqZHkilP94oADVpVb/i
uPBdAZf82pwT0wL8d6KTpdXfkuLLuva35vNCe+MhH0wGGgYNX3NI1Vrre8h/
+L1pbzsMqVkWlgLEnUrtHVKGHRr8kCZiLUsBLAZXfUakI1wzjEL7NTi6Lxwl
FJBkFPgEi9LTdlP5InemSGxPy4DO4kVCIQHAy4A0xGd9Ty2Rft3ED43+XX9u
hFJSkQMnFGwlepEru7C17Mj0U+IEQF+SGbeyexwGczeb2qXMA5sbUhrxzbtr
C/pkL21xszdPpfCMPN/2eew/00aKfKrTqGTulIdpgPV3yzzC9AY8eVxIVRQK
/WDrqT8ViggZCQF+fBL7aaN5yYqL6ZLzmrKS3oolLSRNRJa933nbTytQ5V6Y
sSTXI/FIkCRmDLUiAaagynfDqsD4zz4e7Ip9GY6kuo9UB/s8TdhUiGfpqrap
YMsM7yu/qPsRpB1y5AiZq0v+wICG+E6B6JpRpGp2vRm8H4lBs4U50mijorzf
fQy3yvDo+1vOS/suBg+u4yrVf6FNW5gtlrYK3r12Dxv/1etpsHdfO4cMxEHp
CZs1VxfANrCTv4XpFZZe7hAlkJQwWJkzICsQVB5Wq5vx7YLTd6tSEfrsXV5I
aP5a+HW5ZFlsBdmzwzPpEYq2+ionudUJWalfZOl+3b4IbhFSNgDlfUN2yAvY
qZtVN7Qw1cw953DHATjFQ1e+bwAzLpKYuRKINXr7d/krwm8Yk5Lc0MHeO6Ov
xlS26PsU+FTtGV4EqAuvU62jnqD3rW2n0lPZiCEnkoxcJ18NDWjHvocqzrOq
SxZ38X6s++JoXqtg4l2i6VWsbmJynNpPE41MM3n5bt9pOQEIpi7f49ozzXG1
KCcyAotfY2sd62XcGeUqWW9sJE3i1ImpdfyTk1U/5mlpM5ah0PLRcbvv4nlo
lEP9g25Hxst9wDCWFaYfdxLziVHk5K4JyQl4X5EBGtqsnZNqC2qHc2I9guMo
wrl1QiR1SOST1hO1QYf54TTacxn7f+itwc99RxW6CShKbGAaE+oOJ+sDHZ4w
eaZKTxijFDXQLK3YsEm1OrD8x8dgnR50F4ZZqmADY8NeqVQKHnLUkveZSkOI
7QLdDbK4KW8N8jnLfUcIu+gl/vnlPFoMIAogmLCad7jNow9+ckbB56TaLVRN
vnIDI3aKFiZ0qZIBcTe/0Qq0xAai/s995ERE2q8uBkd489IkrTPZxSVuxoJR
R7zZHdC97CQyvEkuWl+GhXGfd3sSNEFlK1KfYY7SWnglS/mlSi7aO2l13t7T
M3G+EeOkwO1pdcDEevkzBqgDxR5cguOb+yEO3eUcByVpoqml0n49YN9h8wWI
bdFFRf+k381MDsMuTzFVtzeUseTp5impbRnBzeMF1fIy5ibCt6/8mbVgePLS
oCcCJQvHTTeEw8n4kQgEQTdi6jF0+VxArs2d26E5VCIuJPfT4YCZ2H14CfrL
EL0A1nAV9X9H/gHrWsYnOGQ2IWB57RhP4v6uylttVUxEUH34JaFPy0iGvUdX
wXlAaEkuivWRwirQbVeCSHagyG0QBqN89igMLVZMekhz7PSt2EFA16uAd1Qi
Paes1qSBuMOt0zyrIDrydz2qS2MYmqkAs57+ZH+xFEW9UGO1yoD202nfSY+9
f/yPLQgRvdJTD/LYYcgE5K7dn3VRA7MfUxlv5XVlx7N5ueeVYPKdVRXfkLgZ
ApinnEQ/QYv1dSmuXFQMnFKtFq1K2LmypSJaeIlXxB4m8yAdH9JYjd0U6WwR
v8PgaTGho9cEPaNVE1yEr7DjGaOJzV081TZCfmVBLUTYmmika6uD6dSQon+c
mePdWDpoMepv3NDxnQDTeDwtXFNt3IdUNiAZOEodbjNMb8dHkqE+lVkgAH4y
+iRbNN2XdsFZWSKL4IMKMpzZotR76/y8NnXXsCqtkNU3Bt64lmOkQzZ+jjDd
lPOOnDCak4UiTVapPVHR7Jjkswu07ayufqmOKC3kZ+7Nzugaw/iObVtK3Vsk
1ev6EP58wICti3gllHDSqB0TZzwokTlVzeyJdCyovYOOhpRG52Qrd7XbGz2d
ycdGBYlGcWeVoxuUmGntkLEaIAcigjsjIH0c4xLtxDCGxocoBLUn1C1KThI0
G3mWpzP9YJVNujGPYxrCvDzqre7ZfbRSnV6DJOBEoTdDuuNKhS2BMc65pdE4
nhR28NkantXhU2ugO3/xZ90mi6wpQ5dj/8hHq0q75fWZbfTuEm3LMkZ7PIDN
nprKfJ1XlXCMScjve6aLhq+T+UkzRa90HSJiUudU1qzy5WBI4L8SKtsaTWsy
58x3/c/7OyvpLpqmImjdOUGqN58y482lZq7LbkUZEt6M7Qiew4m/XkPw8piA
xIx240zNtdVSebApbU2W/DoECuzyzZfJjyvyooWcisEl6EqmvlQnrQXtz5zW
mjHgWts3rPAcY41LWuoDqJorq5hK8ezysHvMhMLuyt2MTVFXJ5NoUXaasNGz
jkEVXeP33Ppcw+ZifJ4vug8a05hzx8kHttBmZ2n0KiDzHnomlqL0Jr8mgfjt
rUuWnFQdwgfV+FSsiKk5pUL7sp5Y0oJ8cjhNt10UE6DKmugdThT1jX3eYF7Y
Agblj7V+OW8+KVFYbXsh6yC7rkCBpgZLII27vxOS22R5YchVRjf0hW7Axorm
/flSK3Qbw7bdtFI2VE/hwnPfazhXAx9Dm7kiL/pMA/NkA7+owEa/fET+TEun
VQUlYIP2OhRzJo4S2nYwgKphKN6NDZcZXI9ayMcNk1GSq9n9RMoposPqwSuX
hKa4IoWEhaJBUo3pKj1sfDP10Z6JSn+cu8zh6YtNw5LcV/QPG7qRHE3ho11v
bcAQmcrCuUVx6UDoWCY4lAwaQSaPuZ+/jcixeC4VLhilJ/FLNUVqjAJBQ6AX
DzcDXmZj5hjcxwZuhcg45TNSzo5DPtgZp5tCXezMLf1u5/kWJZzRQnCq3+e4
8a0jjG8cV827QdZzmlBDiBprG5LLPQXzgholMFEX8QsB9qvAKPp6KSw7RZXo
+w0DXrLzhg91t7uZJEVnqkZS3AWRxdLw6cycYrOK8KkBQpjGup2l7zPQN5xf
SVyuWSitVQaV/xcnlvK/jfDNBeI0XJcuqKvLneud7viIeMpaXiL80SmdlNdh
wLJHZX7/n3SSooVRG6L5tpsMVOvMDi3Z72pAh8zZVpKiZQ03moCXexcTUO+o
tduxQNV/xVx1y6aFlhfOT6YR+M3j4136IRT5DmlK2hp1l1uM7JMQvuc8ckOR
sI7aJo105iGeZxq+twIYh2G/MqbYgk6CU0YMFk1TiXW8xTVmYUvU2li6i9DN
ZNmQYKAAcbszyV5blvn6ukje0YlUfF49QzJL19aL412TZgHNyzKP6ugYMo3P
S/Z0jVFd7bOzTnLaJD9uwWWv1hoKFNnWfMsP1CKPC62ZwYxBJDyZPLpTKULS
Jz9bBOt8+QTDOdkA0zNhxF36jzJlt2O0rbvbubWugGDtCKRWAugqJpQe7axT
XfWPPfjWdpD+rjO7LjBKt2fN6OLbCTmPApfwhwP9K+r4lXDe0yDtkKuT6sie
Dlm545Wyt1irUyJg3IF2sESDFdzvZiZ5Uk/mWnYOCMdRkIAJVTXvywsBSZ7Y
eOQtazOfJKYMzDewangiihe1nJEAkWYObw+JuMkbjER05uojMvtOoSvIzFgh
yLNh/tkJvkjkGtza7t72gaZKeToL99guPqXvsnENaAU6e8oFE/IU+IdCe1Lv
xYefDAZUm7StfPFzUNPGIwXvGFcuXx5+849BVFM+XucfsE5UTEymygWelFlZ
G3CDdd8OaichVrEM2vVnxNZDltE6i3wbjXEBnm9jusVSJLe9/JexVY0bdZo1
S8IT7KoknfYoKuEUjrDgTiV0aYy4pfQGF75bgQhh3KyMl39MxVYd1JzJeWys
2x7q47WtrdZK6jvHgYd55fEDuYDiPN7uD+AxiKfkSs2645xsD5OUWgap3FY3
MCpCoqeTXe41i/1OQlXTc2nmHjaoLlBcvdKWxvVv3J9GyCAK7Qz4RTMK1MlY
O67vZHjzueUOFr+Y/mJzJ0y1WHtrV3NlIGVmmsPyNqcWxLfZRJzMUhbn+Qit
9WwvNkMDJxgwtbbwur8o4osY1hKsgkgq/mw+Ai3+xf4raLfQ9q6VFmXVfZN6
redIjDjhavu8iYym/J0rD19LjxUxS1a3SHiC7xHNktahSS2i2SjDcHbG6GoA
aqcmdAIRcHtyo9w2lZjCVdn7KpEhx+QYBPr57gXZ43zlTUfWnW1TQCEGc0wS
HEbQlI5cMMjJsIs6di1jtIu6NKLcvNeRcRnPfMzXkVV3iPrIHup6bb1WaDEP
UwBwzE9xZuqWWEZmMBnHokhwwzEQMHbONnmTlUrDI83o8x1ij3iC6R6J0I0F
FxGXX+Abeg7qe5D01ywZS3dYDyxNlieABhcyjR+I2q9Ald7dAGv7YHZUFsIM
WP8lqL+ECD1enEcn2RxFduqSCT3hPSy930Vvy/dTIhfxU8/dZNtb1TvdmB9k
DPxAfGLyxtngM4os7QO2q7MAGq4XSFSYIkpI/nJPYS7NnryBn4ycgTY22USX
gWTBrHTlE8Fx94oWiHVwIBLwaSiX4wx2N5f5bJYe2wsOeKANr0n8ETV4Vv51
RsDWalfqKMUdIhgI21IoJ30PlM5fY3nHdR44w2Fh7AqGhwy7vYN6AK12QX0K
/RbKwIRilU/qnUuMr/GKTRKq/5JnZHeLDe8TmhLu2fbZbuhwM5OzK3SaXKPW
UBBvXTDoh+ThtbeOTO1bQ1rC/9HYuJy7aqFC90P5BxHbHqqqd1Z8o5RDCcKB
Eq+MSV9zLl8IVBXaEb6mzPDoSZ0UqxSvJhNXPZkK0duEAJE40F9U5l/jppjl
viU7rIGPPp7QryaWrPIAKwX4YHDcY5equdNAk16aXAVsxss/iBXGr6mTG1nt
A2iZiCGBDJENtPpvWifvJkaQR6GBF9dO8iQHF9cYnMHNs+QZlSQOWHD+rH50
ECrMUsixnzIKhwdwd8HivUsGdId3d8AM14TUHKCbV9zL7waqlQsEJLXJWxL0
Tv46IFRvYfRZV4MeLzu8GG/ppGJ4iISjKsCdv3MdN4Any8omtL7L0Ep2yoww
WEFU33CfLrThBkCbf2YxFAMlMSlB1PNSouTgtxjFMA8cUOQKypIGM2HUzDY0
HuHPAODc6FIweSPBBngSdXodJJjVZolSBuRIXDbdyFDDjtDFwEmPDeMK+tnK
QYkRtmH0RQ+ir4vqsWvMg95+8xqheazTPZ1qL9Y1apJsBKLDkOQTDTK18QHc
7TNfz3E5KAaahJ2oK9RXKjOyfNTqcmBspY4cEzbBllIdA6QJ+y/7K4E1Y7jN
VF2e9rZcUR/9HxuO0LUH8JBLZxUEg7NqkVstGtrjvg1xqPPMsFZEc0uI3DXz
cxeyhDZ/+3v3Jbo2D/b6IccArhe+IcID63p9lwxdLhcrP5odfszCTKWieRMj
5tnz2QH5/ql7oZUwHo3DHYtzX+xufIvfpDeLo9ZJaRgGtHajeITQqkHkAdIy
6V9Ul3uSSB2ERhQQQqfEgydm9fJ/aVUr2YZBhS2RmJVEt24DkSiQZ7tF5RZZ
m2x2WoGGITJ+8NPSINbICucIPmGYHjsYgari67Jl/m+VXFKa/1CxAdAdAVMy
FKbZ/4rxnI+pOBbKnJ1P+3MJ1ReDXfQsISBvC67v55a9mK7W3FFZiD1a83Bt
KRiEJ9KVx8N3+yFotEIJ+rCEBf/nj74FYGMGYuboIJR9kHjaMrZgokpvJjvy
a2bd4oozMB86pn3JPDgNDP2EX/DNOQ6K7he+pQoiwwTTUr+ObBxuSCJa8T4k
jfQOW7eNAKjWG1PkYNmHZ8qZGjMLpzrjcfjjdHRfHe9uO8hwjZIxjnVBYyNT
vfWUbPZSVlYWIH8mDCIZ2bI9zLzAEcv8/xcz9AkVeLl6rE7K9V151LgvIT8a
+KRxI3pQ2KEUW5kFIcQIzKX31arIHQjttxgXKcnA+uNGO3pFMdQuTjQNJ9Dh
YEW487gClbolENmtcwwYI7tEIuOH/heA47Y0SCyInv0M36YrB9tyHINtavjs
asG+UV1wRBD/2sq98cryNeM+mqlOsujWUEviWARJ/kAYlHvUz0/AbgQw3JOL
ug8YRZGcJMzIphIq2py4GxTxI2F5JObZknSlWhj+L2sIq6/wibHQSquedhwh
W4ycO+ixg+5OmiHymID95m+1MfFQlPiFVcOt30spxHO+nWYNRp+bVkbruWOH
SZew4E2+WISWf5IKyPMAn4WxJuExt91bZiXeiqxlsQycfJ1V62T9xXtgxxb3
V5yU8t6WiW4c/WV/72zqPAiC5pZPFe4dF+kles6WWucRvJs/RTvudlFN1/as
sc7n8Er2sox2HGXE06HDcYw84Cq6BI0oPxNg64bKnufAQRQLmb39vHUSm3dM
TbZCgSZAEN5OJDXwh63p8apRYJ3dgrwIS89mHvSzS9iEV+nvN6fDoACYr9Og
Z1dBnQhVFnnFHTszX5gWdLn6Rv7S0QL2CDEGT7kX1bXok1RxaqIDMQV3wyOH
sZLk88bkBBA1WUdgaiONOWAPJ3nvN+ldym40OovFX/qMgNUTjzFxb9eIM3mr
feEbg0yRW8T59MkRynsocIEaVt+3G54hgOZKMWomPvErsKgP6y7OBgetsHtU
VswGnuFClDMxo6m9tbp4EItQBFqJ4uQCizSu83ROFf2un2YGNcfTZ3avpYJu
ianJGhEcxHjC2mpuqinlwGD51ypNR4chRuNkOZO65WAu+9luTrB3Me2QpbqQ
2lGaDXKwQmVt/0Rfd150jDi+afTiEEOjkvWhjEhAD++ugWOmSkSx/Qpww2b/
oib0s6TklHAkIQUh2aymF++MFKshjSEv5NT6Lgxuroy1i33ROdzME+OczHLj
p9x6KtyShRdkvt7D+z5iTxthp5PieJPN6SjqeV4uOZGKBft9tseXQHDObd1B
r9BLowGBzUyN1X/bbQCpZT2qqRGE6IiE6fT487rwjRaLBmQIGqpf08/8Cd9T
UaRm/ghjpk6t4oueCwlZ9MlpRvjwBn8JVQQGFB7mehc8Os+suoxH61739Juk
KuH/GL3VmuDNek4JPGrd43wvhR/xuH2Mi88xhEQ+yvA1E9WtQ8n5/O72luCW
eh7z73Lkc0yl8x3aWzzXDD+scsFzwotuYGWVJo1x7pT9TVa5NnhG5KB+IA//
mqLeGq/gSBoPn6Muxmg7lM13AcDeF7t3DU9eUrA6/pZ+JxwY9gP9Ge0gZOrA
t0AC88iwuavC2p4oYexMIeEWrK07x8+EgNab4kVod1VCql2k7ct2TAaAGoKO
Po1fMGk+/yfiYnyWXi2QqPYiKDc7cWgL7mt3t2VvW+SVeYJIdw+zWwCw47S2
+wk7pwmvkP6QWQ0JmEBcwlZT3AQ5ZwU3zoSkvgyo6vIEUTdqcZJKN2PC9sZO
i8GiQGAKi1zwRfKsEpxlLK1KaEq6ozUS3AzsWK2xK4ESeYga/35j2jCzsV7E
/CXcALYMCokdObqYB+gypaUV2XhpD0WGxck+pJopuaxGMInVOkupW+mx628C
NNz4z7OX2I0JsxTQ0rD+GsRYi5/Gs+nZwzjKt+jq6wU9BdWb4DGRBLDNNtnJ
SHs27DeyU4SR84yjX4uEO7Hl1i/D5UFMBo5Uqo1DkttWq0V7BciOgZLVkv4G
smCVDwiZM41MEur7q+t5R43UWbT5knw2vnufoUzeazCBtf3MxDUv4XUdvJBN
hkC5pxt3/CNLj2cvSF366mQQ02wC4utKF6Ky3SyZ5kefTKGl7YIJ1yWBxg/M
MeJppiMJBTGldlfFIdW4+rL9s6OVoXc4i4+ZS+nl+n3H1+Pph/sA5BOgtHff
z6LZgaHYVpodjQFrP7d3Ch7KF+7pyDF8/nd6GIU1W21UP/z5IxL6IIjM/j3Q
F+cvem6yNoVOGctK09NjKF1FAfpfhck/thNk8FlNyw/pGQQ3LgI7gwDxQHno
++jrLDS/Pg06gVZGRV6xIjaUb0uIhS1cCe5EroK0yzq/Ivi0MWiU3WgsYGdp
XmOMd2XdGqUzfVdMafdz6sm0xiZRL9esUnYaLVb7I/ilDLUmlgd48D9nLr1G
p7h6o0+cl3PrvHjsxcjkzp7nvLeU5rOjfUlkHFRVevS1CikZimFocWqtJ1wo
SVC8mv8sND8IPdyGfDgqSruivRO1R4lU1YP2sZn39p9VJ24+1SpS0t5Md3ZD
kOgGhLz+yie4bPmHZs6vjDnp8FtNNDyb7J7TxU0qb7R/4VbqWcj8ZJBNQjJm
eoGt6kSSdkIzxHn1Sl8sMK4/CkKjAKpnrukKnay8kHBx+HnpI0rDMO208H/2
l4LU/4O4heY1Piv9F/ZF/ak5i6IVXBAiyQV/C1zP/f/LoLwXhdKD75EbiY78
wXCMgXZwO3J2dbglbzZv8FtkjwkZncRIKxM2KJ69sh4tjjKwjZVJkpqFNHTd
tU1ntOHG3Ps5Zfr4UF5jJK/mu+/sdQ6NYUg6DtDcpGOf1roaFedNRauOQpYp
xviTQViJthDZ1w4tQNIV5TT/T2alZOsfJqVJC47oEN6Ne3ZHUCwYmz/kxBwW
Xdag6wtD6VfayvwCXSxRUvS7/Ww+8yPwkrpy+rZH0ZVwHu6OXD90bAxJ3F6F
hwkmIjt9PEoZP4Prb24BA2jbhxxsAYoq88/9+NXkkbngqAhEDJ1FTMb4vfZC
35mH7bGYC2CndYC6lNmEIlPPXCEhKYGoN0TWjvWOBLOSF1+bgsvyKceOAQtd
6dHxlDZyPAJE4kzFTM8N0EqzNPIsi4NLy2HSGR1+hVNZcNt40Jrf+sDPuhUg
ydQ+0b3Ot4fS3Gp9G8jcrpOs/a6S8dDwyiPEUdsiUjDBDIdL9H3B1LGl9t0G
yc9deAc+7ggS8olwytOg9AzpM4lybxM+oO4qPE1ljMrU+dLjLu4I/4yDdMeU
i8YxlivL/ijNzGuS0Nf4mX+kd92cBqd8vsrSc8XTDo1d3EtPzKXttVbSkLZt
o6aLH57yr06ZwDJnjvwtvrAX+wQtDxWlFX1nckvAG36tPml3zpNoG9GguUp+
BnNQeXcSTBrx0JklOf7vKRz4ZkY/H1d96ZVPYxG6MSceF5ZqjfT7yflH15bu
hqi2YtPoETxy5zfPVZ1QzJoSKrFNEIh+dK6yjU2SRo2ur4cta1Y23HI+mlc+
cHMdWRwy7NRRqr8OjjLcy7jU2i7SVEtTYZiJKt8rgW/+Jp3tLvfVUkOC/ec/
Nxe8VqdkXsXusf9g8vz6bTjMoPVHgSDa2BVRU8E3G+F0ZoNOsvZMU3Jrhv1H
SwS8V4+SW1P2Af/uckxDYfvpnnq/+TwYCurYiLWB6pd6OMu+9jBNQvN2SD4y
VGlHbt3FfDLnl1ZntyyI3atN5yX9/XzFOPNeRJxkAYnTfT0lxqPso/kS/m7U
gL36HeXgBGbdRVXg/kszl5r0immOPcmURIMXDwee0eIj4FDNi/HNzdOQRXKp
NOD8Ro9HEgyXmlpnSPkH9bdhCCx0MtyqBNJPSKN2D2KWx3jirSotlhFXG4HX
0bDhU+Lws5Gwj8m40S6apRbEVyAaQ67xYdawblBukqcf3shFPAUqGX7F3PwD
havS1fJeIaYdLiBt17vx0plaK1Y9Y78Czc6XH5yiObXF7UgfIO+6W0uPJSkH
sZ5uxdVUmhghSFTcFXwW4TsTqGe7WmuMY9YGLcatGW3issqjzr12YeAyB2QH
QIJzdwsjb/Y3J3Sfndlsz6zw8TJGEb2yEaL6n/8tP+sLhNlFTUkckAXIkZfo
opMsSIrVM0dKOY0/iz9TGq7Z/lrwGalaBqYPV9A1vttvkYX543W0y1ie9D9l
9yI5HTOCAFvy+8wqX3VJXYTsPMt7rfMBaZ0YNYW5Faey3bEUdsYyGAB/mZWi
Q0g+UrVpArRU17cvlXxVE87RsURNY9P+VSfkJ8HPBMWT5mWAi1yC7aUUMR8H
M8njH41AhVLb59C3kTXptFJit9sdBa3KzFKciJadC/5pPsAbVWg2Vxau2KDa
kTkkQBlsuxuJGhbZWEEgcn1N0dt1H+eyKHubjTnAqdRHBRcxcU49fs5HD1/R
QB6FUysPFM28klm2zHidM0lRixSUJcM5YcWQCqOUsUDyztxkJN95Z3N+X/kP
r1NCG4uhMWHymaVAj+FCVugOfLprO9ho1+xL/M5IWVnbiWlPvnAmmROtwG1J
/bRMuZ33qt93WwE8A0nqsnh/gLE9mISNOWuddxUMZuLXQ73bF05U2F44v7oc
WuXtOWAiO1i5aP8IJAGIiDRz2uKDrSTb2pMbl/4hqFt/bLA0FrJGbJ9A3lP5
AP/t30tZ8upWWDJpAMo05UGI0a/psAw7c2VW/8WcFcVwYvOXpIU8WERergGQ
gQqyQ1YaCzr+5egAjhCtPSx6TG+fCRdAjUwxVeo2TsM377GbjegQoTwti4N6
T6XfQeqqwGBDh8giErTQfQXSd/rX7B5ku9qizt/A6GgBuutxQ14x3D/Pbo6X
hD/XrDRGKUiqPi25MdgoXReQXhbpMQippw74nMOCK38Qp82TMm1Nd18TsqbZ
NDBSXupGPwjYdxfZ6Zj1I2CzXvCz/dSXwLCZfdBdpn9+wRSicREIQIYC6wMp
/WSFKqXMCcFi+PAtw5JJaYQPH4KseSm8Ttnr8mHYI8ykVzn2gTnIDiPQ3VGG
wQmlOGfLHdz9RM7IiDgBcd38jy6Q4iWYwhjAba+jwmrK3TNJ9gHmtSR778gX
8pENnaDYJ+CoNs3JBuhzA64PBgBCb6ekSdYT23J1NVUiEhkz9SJHoE/MhYbV
hQThD7sRwHrMM98r0iU7NNnCEzvj6zd6gQq33Q0X+lXgGBCwwFaOP3m/hKeG
bjymafcknOpGkLB+NnflmnUY1yZNASUXbB0IsZgASpKWHnJkvmTY05LHUXYM
v2O4Ylx6ldlyaYcdOdw3zTQJYIXqKJhPCHRAmUsGhrk2pXB6U3kIM3Udklzk
dYQ7GUG/IhvDIXkU2Mc5GaMJp/l4TFMr4Hgn+/7lqFAjUVdaPMp1YHtjDnib
nafEYCnPlkL4qVE8qX2GlVKvZTLx5ovk2XdI9d8I1e4ETUNOFtfapqlute+b
TFgC8EXnHH9da3Ah4SrcZyPuP+19VUUtuEsZSc2hFG4kCJBlk2g5A17QUAgb
Ai0JkmPtudndiiSQMEXZWXjSZomc1ZCZi/hbHLzLL3UXpHgVqS70nDLEtVfC
ttSL74BN3nbtXCDDc0vE/shWcmPZIwxqiuyHgID/ZDSW2iPVL5wptTKZKjcM
oYYNZoH34N0aNxGNzCdCVp9CvXoYvH17lMHMqpsd1MNeok/1wmTPNPtFZ7z7
r1pwYhXRykwBdivrbwHbwHdDsxJlF7wEk+Q/HTSrqKjZS6zXT9Aj5eGqQ3Eb
vLIdV+b/wbg3ZYFw/M15ZlR0L18ngZfhQYVvRINnlDWrfwKhu9VBVVBV7NF3
Kl9NiZ6anNtx6uxdDAykbDdwkRUYL16FivzS6hLkcXBA3B00kb6F95yZwYds
n3x7fxMyACS1u20it1bhksG+s2+d8PrqB5v55B7nkZnzVEKnO31AgSbmT1Kp
CyNUS1ffUCGTPPjBdbgQ+5/9RrVM51LKana3kP+fEj5y2c/O7qNRenaifugu
1v7rgYoPH/5bFrBQ+7NXsj08WNMpNvDQiqsEweLS9gIBa162+yNphLTS1LQv
V9zzNLHh+MvzWfZFygx5CKxZ16t8fVlqPRoOZwav08MdrqMcaSz8ZmAMfABc
dMv5byEtvT+/sSa2CAcZhLEC8GsirhKvFlK9WHNJyTI0U3UrJ9ZgNpr3x5tc
pz1HZFvPX9ZNPe+8B3EBJia2mY9V5BQ7ePUDCfuveLXF+ajr/1pZEPZtBqgZ
vY5OXeLxAtQuyedQDRT0OHfZ4Fov6uEdMQokhoiFxHzPL2NaYCkbGGQbGw1a
7IX1OSRZTd1zzUp2+Bcx4UepcuAke7UlHlvM5nEJYgs1TFcEHQwJAGuwRy5I
Zwy/Egr/kvfdQ6RAdb2f5sZJ/7OZ+ygoIH1tUskWRvFisM+LX+9MPBiQ8AOs
WGPAcwuONH298RPinvXbRLHCwyTg3wOpsLCzg0HMk9AmAxOWS9itjnVi6BTQ
Bfe06+rQH+OR5tVqSyuJKNNykwU+I2g2m96Wbsbt/ValnVKlulogTERS27P/
tJHYRpGuf0lwJeofnvxipYrEFbkHHK3t16TunD6i4BuMiPTGy+a6qjnQo5VC
TTh+wz3H/GdO/kWrCz1UnG6TwRsBZTRxA1jqcldYoPf6uq9YWy23+zQfmssc
juIuljLfACdxiP1QDL9ZbKmwOd2ZAolhvH0VxoSDuLAh21yDQV1PRGYDpib+
bN1fMoxhPg5KIdVBYUxdnEC+IZJAnpxKtk1STlNWtryYhZHdGBGieq29jky6
D00vwB44wJydintJI/cgfQv2echVHwXXG2RfO2isDzhTP4l3w2HXDWSF+WCI
8fZ+iBEA0WX92dHkSg/jDMtHO6HtYG9JDorvzs3FhIV8aK97XHAFoZAn4YgP
PQk5uFvLzrg+LmDxGCIPvB1CzX7NfQBfBtb9xkwyXsGgLr1u5ntQBHslB1IK
5vGRmrZv8uaPpL5dBD/rPTaxW/z0S5HcZNaRgs+vDibsl9gWtbOz/n5YZVwO
1t7lLJFOMZ4J7hAoVc5aFbyCBKgEshLtG560FGCGsR3f3r4qz6QOSXlU4cGC
fgmiQPzlsSMdHBnAJgULgCEqU+0kR+BFxi90ZC+vUliP1pHSmBuApSjJFcCA
iOccVNbDZ/NOpiQymdnuP4kX78VzNHpFPsxJ64AioCS6UxuxWF2BKmw6JGiQ
vHCYF9lbraFClyJ2NK1OXjYSBlpOzbEamGSCL4BAZWmqSXUURKPlcT1fzzJC
d04UCsFcw5x8tLHNEsiuDhnfocyIitTHshs4EnWgiGUL0Q3aT4og1gshkKSO
z7z+FKscVnlO7bx4yyNSrpOaecgyUe99Gr/6h2VDJgEvfzIv7or5h+mY0naY
tvr1hhrlhD8jY1U1ff8vOq70IAFGfxVGX69MM9gwCPeeCIZrV9t/g9Pumw56
t2wSLCq4NtzSfJ7v3baEvVLmjIUM+xAtUwjvlX0J2s7u4/C/k3rAw5IpkQTP
Q9MZDncdZz2ttgzJwmPhw4o2fUdhzBavGWPll9knsgTksGqffk6149BgRF2O
yw1Luf88ZxafmJOBMmO7Hcze07uKe4MSTcarP/jQsx1XRye9lCg0h4Oh+dwt
EZ5fPbYFdRDDJJFiULFlUrWE7kai1gACwUx0UPJaPiCv2m+aHzSY8IG7QyyA
uQfY1JJED4AU4It4N7QxQlfgPgweJsFqX1V6RQHAYxCiXbNXAfC/WIr7V6ic
vLDhEwvZl7mzb7Jq2HZB8YcDndtOnpLJoBdiIIs5TZhykcb5lDqt4vYubTxA
OfZw+D/roRsPsWpUPYsuaqhNJtX5oB1As3YsvOeYebOfOFnJwrjnbog53ERB
AEtHgSMbhPswkB/lsP25vrveh25WUEq9GGsnKFtNWzNPhNQL0F/8wGuO3jG9
3s0TvSkuQZZC201TDNssKl2UE9j5f43uX1fLNQtfjyVcRBG6eg5A9kfqprM2
MEuSIlePP/qy7IZkd6UJ6ukuwlnSxsOVFm8cASOIKUn77uHhsJt5bthH25cP
4S6jTVQCtrNIBEgEPuGHxvDKkn4cX5ooJwg9bO5/Ts9twFxm7LX3hItLML1i
xhLhBeuo8Uv9q81guPUbXs8gsKoKpQBqQgX2yruhPd5q3rMItlaJ9dWAbrjW
pdEfw6PS1xpCPk4M8UUKw+ZaRBengvQVQVk7tLkeiuxpMsLoYLB2EaLsxScY
5MSsr2CCEJyKG2cZLcY1Xv9SHi8Y4qTiR7OF4p4AfF087tYJ7NjlYUPY8TBl
gpDsfQsNLplrErFIHPaQCpUONV/Fev0/ihWmz8T9dTmFS7m+XKV0COHjDiZa
G+3hTtegM7bjRXuOJ2NWcnN2GA3mLAI8Uh9NAeXAWoDfgU/hX50WVa/8ZK/Y
LnM/grkoigQ0AMqxj3CWaDSb2k/37dW8j4S3vKTHnIvsgVT+qTCD4rDUd3Ac
WSYa+G8lyQkIXUtU+Gl9RcJGPu4FFtrZi9w9kN3AQJ4SjWriq9yuxSlXlo+r
yTLlasGlh0RsTgr7bCQ8GYgx46LFsYwsA1g1DxVhl3bqh+7WYUxm808R2raE
Al5OFJqNzvDkFXaAjLnLRJOrk4LfgVo/D0f+YBMgHvlfEr+GJik0l/g+87YS
5xq01sBwq1IA7OiGap98JCBDwgEG4vtyffoI74ylN3UC4K1nGoJepvZjwqSV
KVlYxS1w+ZtI90WdjJa2baPgcCORDzW+j4eXKp/ddjsEXOGyHCuXBbGpd3dZ
le4i7w4ne/lb38+Wo+XGWEdEEZY9Co1vjs9MPGlLH+CNj7ORbBw7ikPl0U93
2tCIwPTgDLND3Tr3sAF7/AN1Z/Fgu4f+0AgZJYtbaNu21GUEeaZv3SiLLSH1
2Gq9Lo8+8fFOx3/ugoeDr/6AI+h2Kd3hPzJef2mmNRqSuSrghTqxtY8kcCCL
pqpEFR4mReb6PwMTNwueEaQsF3FM8wk/NLnB0xbEBCtqZDjBIq/3aXyS3QbV
zc/9Gw7HIvmfeixc6rY8ZsN1R693416EGvDQzBt4D8clWVGnrmsmGJea8z+k
4xdpPOtuqaW6zekWP7RmSirRqm7zXaq1RpAgI0NyGtfq67TPiP19EJanmQKG
KPiceLK84iZ5pHgHwmmjMjcLTv3+KMhbLlyLmufwY+c1UhndoQBenQwaE9xp
FnToVWjGWf5tadlG+cdhMYEqh1Cu9/dRYPrIqyJT7C53lKbIwLRwnt4poS7e
dgEYDensy/A/gyKxsvQe/1y7i6z35AxVevy39bTW8Vrt0Z1Dn+W2IsWXnwAy
NTEN4D37sJSa4e673uCsz/YT+QNVAj+lTFwWeIZP/RiFmP1+HqigVAAD8053
plMFyqQRxbdi6SjJfE53zveO6lYtFzJjvDj06O5Pr/lr1G0MvVf0FnqXXob/
vXP8i/oAcJ9IexXUOsdaXZHHHQTeuzwZ9729MoGIKhjFalUWxRYaJq2EPNpC
MaR8AJP3u4TXnuIfHIKk3bHNr2uLRBcv1/dbPDrdGmBVNBkTMKQzgvgiGbxG
885n8hyqT/Gr4+iK6gVvTXQ3Jl3QBcfH8HsORh+TXLZmx3rcisIC7n75sbXw
eedypVZQKfuxAcf7Vj9grjVr5NdtdkwzOj4ifgMAj4qVZlG3mv/bA/t93js+
3Pv6eUW1T2k848iumPEvDkwkrrXZeRPnlGw1tVlF5JXRNsm85+Nrvk8kuBe5
8Su/EKm9QJxMcE7YNAITMJR/QEna6AHnm+REpBOTM9pWQW2wpAXDXh5EfhXG
GM8JqDq1DqXiEcI17gNyPyKBLe8rlNVtS7N7lspkfYbQnpSUpLYs8EWGRoeq
e4qDtguxxCwi+HsTvf6gdCnoycw8ZUThKBZaDqHvObOq+OIpopAGSIaNU/dl
V6rkUDkY0X2Dp6223hRUG9J4HO0FZcSJ2XKNor0xn1xdFC5PSw+SaeowyZaX
bRYbKKw9wZHffddThXdnB5fWKLLTPUV0dNiadBrzlQptFa/rf8lcZGklvde5
eMQHd/K6zDj0iOOYDyMi6JbcNHiTI1fWljAWl8lHvNcLBxQImFyVxrKGu4Z0
9PGwAobX58Zd1v3eSmwaWAs/Zl+m5Qsnn98+2U9mV4dTDAQ/ENhr/Y6BhzZq
MzUKXIBclOYfmVVO0VB708UOd5XlacpXz6FaXlqGsGYpMjI/3te/fcfKptKY
ctCvtgGTGiVqF7l1UWg54AM06/Nw79o1m21Xye5pZKCmV1QmVZbHpGium4M5
2JRxCzTiH1QESCnXxq02JEjWWT3Fnq59WwAATxGKj3UzEGT8v0TpTbAquYUq
0AGjcbQ67xOVGi1KVdznEEfd8SzYL5L6E6wR3YEGayhQ3+mJIsePEHCKtDAw
0kWluwGc/m+dGdHQ57+/8soDoGCsvlxm2R6n2UUtUQOpZgNRA2oS1AEi//9W
yxlZJ/Kv6j1RlHWP826ZUysD5/Mxq5w3i1dF4B/E5D9tUkdUWhPy1ZQEUuSx
qSYp/WHTYyOJzO0BP2Wl273m80kLV2UL97lAI0QZDwIyfUHWkrlaBrQwycN3
k4p/xD10Tow+JWekKfLWyyutJf8X52UsSaCVLeD2JOvGiFJFS0doHk8mtNFt
4eS0kdZH8ukD1lL0Jg4iZyZG6g54W/Gt4LJ43ibr3z3fAelrI0UPM/9C6KKo
cMWXWcprUWPXAYeFozc5FJ6AcZLqaS5R9ZKHZP8v+de18nVNHEFU7py70zr4
lVobgrMUqIYjm0ib5ap5zKSuaRPt3M78rw02eltPEby8a9QmRxTok4gCCJFr
/YOw5AS/gcUaD9+UAwCIbZ53pPHZv9Ruw780L2AF90+nGya+07nuxDi17xxY
NL7zaaWN71M4cvPIceVCEyrEeXi/YJUBzmTgS4bbZ1cXHif0kbFEY9H81Y4P
zUd8fvC4VjHCSd9tkY3xq0THkVuez4dfJ2AYAInvYmvkWbL14G25Cn4v3FUy
kjf87kqFZYq9NpMm1CRhOTTLyvJ9J4YqpyCFqvOSTjQOfBLgkPAFOb2rM4KC
rgF2Cr3k9tXx0Seqzvpqca8L14PEu3T8IV+ZSzULmNvetrN9yuFmk8+Sni/D
6RCB6M4IpBVpsLcfguH/0SwOXqXMibpQzMpuFTh5Jdt0i+7WPxzTfcLrrG6h
0jlnNpoEPUeCj4xiM5+L090JV6/XfZpE6Vo5G2KaiDGjn2MfU3+X6zx8AxqJ
OfWFJqG+DXgdFPjkA/8hab3BTKvaY6cH1ktjkOVdz+K262qr5nrtBYDw6MeM
qL/QsoEluTqO0APiLySRrSeoZEA5mk4AxjVv6NJ9q7YzhjlzAJE1jNcFINzq
ZMukaCp+BH6okfDT0plAlfHbjyrBOwoV5PjTeDRYsm7ilz5mSW9qQZ8/g9IX
4HZC4/fYspEXxyxd2fI5rVMM0ZlKPADI/txPwDdRZxrkBMFYKmKsqkuRNNJ/
bot3x+8MTeu7z4+WHwi8OimukdQ2byTf3RsaRlDVER9xNTkafp0PMNnbNiHw
HlSVpM6CekcA3qRGz+/ykOg9zeTODE14yOzlywoxp09wO7nHVYYGehd0Gk/N
zrrfHbPPuWP5zJIJ0dRVknI1AgXZNMhZ/RFH9XDZHYevp4viaRGRWyOa0Iok
Rpz9dSnEF3iwyk+82ay7agOc0pEYXf4qymw+JkxUXc400Zc3F+TV9VLCPg00
RnahMJEgx5sJi4AAgBoIyRBYacPCP4LyaJLgoLYnuNkv+jkwRfEGdUk4eMLn
NfldUSoLa9WY7N6ruY4jsKFE12+kXzcgBhGXkdEdX8oPfIoPf34FTvJjB4rH
anH42JahDYWxcAEIGc3c11l56wAQuxR5j/3H78rSOWztkk2Y4fVevBwqC4Hz
TV/YgYQk+udjuEejWebSWuFpsqO3M4g9El5vZkKVxWeQTmR7oeuWasYnpSps
WXO3RjScmVzky/ooZUJeyqzlJJFiUoWSL1/MjVH1G1wqo8Hw/mJyQFhtIFgt
FnzXI4Xwn1BVd71pFAnnE4MYLpZRn1+tQ7m5fGM0jJ0pPlTEWxvCy8ENtHem
NBbzmaukZgRf+4forKLK2Y4K3prp+8qSLEQ3bDd+7BsVcq0LDizYSPwtQkRb
XuCdK8bRx8gtyW/6c2skbsYrfsxX8f1ROj8K4rsBTjhxAVtj6BDESBBE9wFx
QgeELOVKyHrRvwhOXQOelbKXuBZKxw6JR7ZioWSYYZnrcTRasBKJ5X4CX8mK
rR/QnJBVa4QV8B4WvsxDAHRA/8AqmNsvBggbyAnMk6kC2gIkG/+MT6lPVTlA
pMMpTY8aUD4PyxgEUN1VOBTKP+5nk72gwK52tgC88zpsQLsZw9I1QYscdJQe
Mbl5EM0myIs7iu5m4XxK4KGIhcm3iUivHCXfZD4i74eHmHiN7OxpZo4D/uY4
T/cWgoqRePi07wQdJbBDDXMhSiVwk7Cx/VVHgxTwykGm1nj0ULpFtBS6IkiJ
JIc/kwItbOjiwafz35M7lATM3VmKdksbTPgD40QVQwUGGxgIF4YVjHUOjROk
sqCQlxPFXWq/hgKHvePFAZc4zlc0Ztrsh3WYRlvL20KxztWjgQoZrNVADkEQ
aPAF1NQpBmtpqCn8jeIf/UQ0JpyTM0kgeS7AGi7FjEGs9F3DNNx0yvyk+jH8
7wwn9FiXQO4dSciIIH568K3OnnjDu/a3Y+qBMOVwyUY7n9ej24TYjN611OPu
FWNw+ghDUrt4dK3LNO+Cv2mr6NBpdlf41vqetcOnAScFcOUnLBtmbEMCr8Z2
AFk1E5+fKWvBWsfY8EHIGZsrL7TlGTT0QMWxPquYy+2kVbsKuNucpejZUVOr
s5MFfOVIc0+4P/XgD4dC0ypg9v/cRTYf+L8hP5n20juoN0QxOJ+vF4tU3exp
yePrrzYAKdGyvSpIhtTdMtGY+933UMlcFB0jV+REUEXIF8PDQfthn2PZ/4vC
WT1pEqTJ1VPu71TXkd0tiGCCrh3ZadSrPg0yoe2Kt2KnOsDgIyHYbd9tDgzc
jLDEo1L2BgVVDUFI9sS59JtLZ+nMaYn2lGxSRjQBhEJB/6eDopksNgFmwFl5
MIzzdtB1h2yYD3CWO7mkFqjZpLmzX1F68+ghLu2upTj6qkxZrgTPjunzKlyj
LG+k4nFrWF/I0ymohrNa7ZtwszG63ddiRuKrWK9uvIGZBmlVtFXH5Q7pkIWT
Alj2PKaMxbtZEYnSSdutC/ny6xN42stowr+wemT/YUVVjIV4MFWlnh8yL9b/
suuzx8vrqvmqRK1SuRPFVrYkWawE+K2EKazoP774MEr3wMHUf8AJwhP4JS4I
brlkKAgnQ6eLQu5vjzgNXqUVlkzi0Jb0sXfqG9eT+PizV+P8dUjYpkSWSZpg
Z5VirX5HX5LoJYExp0Esz4oJ3/lw8235r3KXoPJxvbkkLcAbbpeP58K2mpQu
uXu9o6XIUvf0Pm+dw62hldghApad066Y5IDtb0P2m2ktCQ51bwi+ZuZgicYz
Aam8332JFLN1Vf8HVh+hGs/m0dukpnABbyks9SEGeCKZHAXnPMpl6q0MKj/e
tLIIPqqocwT8LYVAFM/cfN/qF9tD8vDgx4TcYpTwJ6vrtlOrCb2Bp+KOZaE6
sSMfBP2/wX43cZY7Mf9PTJv9Khe5chLrqR/DVQhFXPxySEiKHy57Tch2AWLO
MVoI/eKeNibIJysKQGzDSsY+wQLCXO64hFK60H+zwDmxVsElMQ1z2DhAPYeR
O3rFfgPSrxaOEJo4hAmR0j2nFPe8nHF2mLLkvfd1uSjSisIf0seGYU4/MpQD
quEti1mZokpGhWDQ1qIIVNG3uJYDsi+tS82wKmKTFuSkJONO0ELpM8KFD7VP
3LVn+9mDWtU/db4zSgO/cB5g1SQFj3pFBMiWOzvICrW08Ml2VZBaXGbrYEGG
eIsw2wwamlPVeffRR6WqpLoDFR6dIFm4EfAWDFEHObfGkaZaeWx7R87LGFzZ
6U9xJfowIWMtSGCk6n1750WC6DR0UT0ilLih9olkwzAolBSHMC1KDLUxtbJk
Z3oNPIyESqsIffoyLvT7jRJmUmRTst27JTchU0yrEYGhdsxIk2WeT8mwYSR0
Uq3IiYVkaauArHBE1cp2V24JEEH9WbxIeVP4U3zfxY7Nplg/0SKyhmRfs3Gi
wR240Zbj/HpoMN2oAJz2A3UIcpmSh1ld/haKi87woXo7IdGSNUaazQW9XE4q
5GaknmEO2w2aVco3Gxf7Ual7LFROA4c1CIopQv0ccRXbvvuhVGuWug+JbqQz
0RZ6GVFAERc6SkYLtHx0GRf2MwBph5xT/MNAYfP469X5XPLsYOmHVb0RN88Q
M6ZH2XEzcoPJknsEIMTaU/ZF987twEhla2E32PIF2oyMbyKyCdisJy8RxriY
R6CqaFhYDJhxGTjc5inbXauqi45kK7tx4q1SbwqO/mvagckhM+W5Jq7g9NqD
Jl7EoJfIWysEJZroSm1yH9vC5ksJjUmvXNtaFJLPJjWnQ5vFUhT0Yudu0tjo
Zu/uAlRWrw5no1+OFL7QMDaLdjWgqlZE6N6PUcaBU5lS0j0undlWh619k88S
/iruwTLDa2OmaampZNPWJosCvCXcFZZKb/ktPc4XTqeoN99YPuVPZtQL4EIY
EypBaCuecHytfeOr/nfA2Yn8U+1wJb8SUsJMn/SbE9f+mcjAnPlyg/tTLNKM
9gxDGO2QJfg/W6lplYqa8BqRf9PUQjaSeg0/qG9U8da/CcdSfxjhH+EVss6g
Uk9mCgrWTJx/WIAsS7era3tFfGTvePlfgNFAULJW224LcJFjPB2usZVzv8Wn
rQIR3WO+hYNtviKJjmic1figd1/xyEBPO+tooO1qqQJ0TFXWj61IQY7il+0d
cHuJQsnMN8tfkVoCJSxdtCoiTTM8/Adr5gyxmDYUJpC1RggBPTaZkwOGEPNe
gMYb2xaYY7D4O6r9Mv+8+dBpCePHxDZeqNINSt8F47cl5awgCJQ7CVrkcMDR
BWpEe2bMUXHaCikZv9S92s/HPj4PxMputLuIRXEmxMCzQJeNhcZrZfJ/fgyW
b3BQqAAd0/i/lfsfhCK7CbB9ziwr6ZUgufO/q6FzkCmk8Y4wxG4dVTVHy/7D
evqKYhRkec/iUrfJOQJe4Wd4AkRY9XPFIHwmxltVlW1oNkhUj5IjEagNGFP7
p5rOH+JMry0XtPzxMaWMEqLkeEITWUSFWnyYfUkbfiacNjrrH1/iTkaZJZBg
owJEUPQMECk5VcPtOnqryZ9EUwKvNI9MjRNu4WfD3nBfv2kIUKRrPJpqbseI
Qwxvnm7H2naBuO/9igrNUF0VMcMA4zJSbTCwzdt/RNzFoetLwHNQlGUflAGT
1wWtYs9ubT1oWo7hO0A2akCwxOv1HHKWLHqo7zyj9TNYL8CdKsBzbwSJ1fxq
O/0Pkksbu9OhzsQXrM9CnHM6lluJpyyoyGcO1iwzH+qfteYNOv83B34FBiV8
yKMuv2rWwiHPhT31w/hoI23lvSeXUAZafTQWXYIDvZhy4kxcRl+unvC4+VVB
yC2syX3Pna9NJLexzOkE6eGpRcvHqRzJSbyBPMmw/KyDmkE6BURO8LQtKUob
obY/T1IFh84sXgpsBp8Lio5zoQUhGv5usGUnon+iPFIKdFbDN7N9H67ScNod
4Oj3OKpKJK5qQsDFAz9i4mxoF3wu+ggLtfMpZw3PTgUUK7Od+s8Rz4Vy6hKr
tjVl4vU/EEsXvyHXF9nyYZdBB+Qhm20W2AB4TbQU6WIuVdkh9U1ieL0yO4f1
e0bHnQtLFYXj6xa2gXm4ulCQpFezcP1wR5fzA8hJpDKV2vo7TenDpoDCvagq
FOzgE8Wd3GjK2oMucaVeyZa13x7B48jNLbMbEC+xXUKH2SvRlhn2qf5q8GyC
iTaGa1jXeyCT5+sVTIszs+ojfFrIvJchZ5MUS0Qo0BYHMbomEmRe7p8fMXWt
uxEuI1YNO3Opz4oqNYkbdpS8T8UzjwhPgL8Upuoi2LVIt/j2fAfH8zIEoFCL
18esJ0p5O99GRQYoHLC8LD53zIN3JT0u+zX4toOfzuMo5TAMnskEVskCVrAc
HWI2vO3CyFvzZSbcRWCm2IodbO5Pu6mgx9miNv5biCw1SYxfTKr6soToonO8
rLa5hBb1tc7HlgDAuEn6PNJiyKd0oYQ1lHH+h5ZjLn1LvmvSbY4egbCIyAzM
goCMSbrXT0p0SEFbiuh7gkGXMLQk2VeO5KlH6w+oNtUdVrzLXlELaCtlH2rI
8CZjoFXSK4UjBXX4RnkUz1ybAgMY0SPDyI9385Zt5XtH2UXY5TWGJgY0WY6B
r1ynltC+w+EUeSRTCF8XB5iqO6JtvzA1CpxERAoNydLD0PVEbJVCdMRzyEHc
2lV3+jZAE5VQEhVJxrFPB/QhRuD4/NGaApdPuHC/xOPqP/i6T18cWwvVQEmY
y3AXfcz74Tl4OmGr7CggatUakT/80nCP856bAvWqNxmYi5bGAUIs5Ld0D9Tc
blrwxLkOdsgxir5ny2/sttGHQ8kBWfIV2Yr32/YrE+bdNlCGaef1NrkS5J2g
/7W9IfGwcz282r+flVdottmy80fP9kO0sCQayWjN67nc1kAfj2c7CDlW3jQM
TW3WccNPMAgQLk9Y+wiNZQXHhgsvH8Z9/7TKplxyh+Myp+9yAU0UdggQzna6
Sz7FnGJle0lL9yZjEKXXAjnHRVyQx9tWKjSL3Kcg8v5WrNIuGdaEfCv5MdPB
m54hCsKtSSCojjoJ5VZLGxk7zAKVrcSMxAwvqNhdDp3fekruI+Vagc/08qbX
N1/hJDc4jK/2YCLNoUIcy06K/EKNbdVejEWsi/puaPQBSjxdE4xMnzW52dl0
dYxASguYVZ5gXp7tis8VuX89C1emFCiKNOODsl7BknJIcjmv2LxMMt5+AsEe
Bd0EjYU3VgFV488fEMOUO5cqlCK1m7361770HQKv/QiMYQe0MXgWMugGX8bT
Zb0RVogX7fYhmvw4WoJZK6XgocLlJJzMShT2A8k+Fj/VSBdq1+YttWlBxjQf
XNdnltaU28Ey22u2M3fdbS4/R82WSGZVhPAz9PYnJBVUE1G+jZkO4srDQ9Wd
TU7dl7cGpuk6KvlwiCZUCe20nOvpYEJ92AFgeDHGRyafEqNIVuWLar4zqLcT
GrNedHsDyV3t8BUg+yjeR6RfCRCRXW490i3YwIFpNPpAK2kd524L/TJ8NWye
3SA/CxqPdk4xykZqdnBOBn7EV/llrFLfvlKPNsk5DNom0GgezAcxhWwiVVS3
UDLmZX8GYs7UeI4LSv784saO5GNw9olYgsg+1Sx643i+YJOGj8dAUl/Gr2Iw
mYTWLM67lMmxU7oU0KbmqKYGZtDdcuVJ/62bow9Rf3rf1FC1jGIywR3/OpaV
vc9PR7NwfEH0HPEQsITLhymaCEMtZ35KlRAxvEjWAoubGbcQZ6G99+n7RRtm
Yn+S5C+Xdp5q4xUNFlOe2cVchm/YhCkqwiAfX1kL4J/qSmoNkYPwOyh9UuQ3
CllKKFyzS3tV+RaUKUo0EJSGM0fKwNkDBVYMPmOWN1xcK16MXVoyUdusNwX2
X5V3BUGjj+u9tneoZux53BembdgDfJX14fdQ2rSVdx6sH+lEZoRt1iOOvcwS
dqvO3dRYxgCRjGJv+22/OnbKw8RxDQ7Ptmj+c7eDw9D16w0tJFR6Lrhn8Afj
OEe2KmIpdbSIBr2kJjR1liMJNPIge+XibhiA2usGqCPEwgoTbbz5TUna2hGG
SFTE9a+drdZFjOe4h82Rt6aIl87Rnbz9RAQgFIriFIQJ7w4VgAzvEAMQMYVv
VoSw/iT0ruKCc8SnvgWFGgvCaYVxthVlsO4FhBzZn6cDONMsKR/WMOcLIwB9
SCWXDqNhO3PwGKzcB+ip57Fy7cWyZYgRJA9yfbL6+cjEFBJMjv5esEIdTfFg
EzC4on72+yI83cmF92wIMzqkQvArhuGsUKS06AUql8uBV9eS35WJimXrQpaE
Or1GxSma1yVcKewLRyzebxfvJJHqgPd56STK9657yGvoO+u+ScqUehSntM6p
gSqiuiYNVSG0gFNLDTUjbG8eUnmGQYEOpP+V8TH42tcgiSzUsGReRdaOKHMj
+1hdO1i+cLB4Jt6qiIwqKBxQqmgdfMXug4MXu4os23imG2meyguueGm/u6+t
Z8rqu/xmKK/A2CWHkkfhqPcbsBvYjYXqazOPNaKAMaj25m5dDOpnn2xZZfEQ
AjVRMi2FZX1dkX7nhm4VmFXGm0JInw8NiWaWzXyXQwRDOtD+NpjnppYqoDLx
vJVcVZygbVKQQsEZ0mO0seR7R2eNw5Q5lm1NIa/O2OS016fLt4fWuKoSqOvf
sPr68PkGzPEksc4jHqnwm8VoP9DEIzMXYyD00WVoU9uKP/UKvYm5MtSCFu4k
BzXmM9JAFNdcYUtUkrrqxgdnVH60wZ1n0FypmDH3nmMAkJ1ywUg5QuiNFxnu
w8AhR3uKgWsMsyuiCNkvaVVZseUe/Gvep5/lx6NQD9WJ84rfdln4P4ZRVlNW
4iSrXNe1M+dXIkGloO2yqknyGp3/FbL04QDS7FYhmq3r6GlLL7f4wMqLa5bU
XlQz//FQ8qY7sWD2HVjCbV2Oj6bsHdCH9uFxbgu7YjPeoAXQOEOjV3tg0Gsr
3oLv+dMCttnQOEt3w7zOkBd71WOLNgGF6oGLzVOLYsEy4Ci9fLg8ixWhn+JI
667CwAY3hEZludrHKAAWQa0ln8j8fqdDW6oXxFGA29cxFBDEuE1nNqousCuR
D/9D9Nvg09oPK8w0reGadzup4ZwzTUtOsKIu59ZBs3HDmEwl7RA+8JBs/wjP
fWTDF2YMSecmUdFYeug9NKOa4YCOa8k3kV2bBNK6gdexqZZy43AnswzAZ3wS
Q7NnXOK3G6PLOMtP8ROHAutf7UZAFwwzMD5/7S2PNTfK6O8cD68+iEfrcWVN
iPimytI3AOqLRXM0N/jIrEpsvaVokYQcKkpoFGZaeEauZ2XX74KgWQ5X+QjE
AnTt4kWbw9VbNkADJzgZ4839bm/sMKn8gkk8kcTGcWl3i4uRJTVy7TPBc1IG
NhUw8IY/Dgm4fjToE+Fl6nHDWWg4gNAgJ90jkAKLMXZMSShoEo2fcYXH+QM2
0oUVdQ1oB7wuvjGdliBUt6rOyyDpt8xRmG3xZXHEEx6qXnLPhVEirhKKttyA
wJZiaW9DWYsQeNLHyI5+4zQjPX3st7HWBSgrPAokSrwpLGaC9MUkm8DUNmSL
7oWKlVrE3XG3n/yAIUkG8lrq7B84WKYWa60atQaMQwZFPl/7OFOKAJmxUuPR
yo5pLkXEC6JvCdn/2nx+Z1gNWZ2U9XS2oJsT4XDd1eXP9noZ/bILqMt/M6q1
zeLl5C8ffzf8Yn/eNf5uEN5gg9wwB2oDvkyhvgPOb8+oVD4lIGRZRx/dSyxr
qXIWloIqBYAgyNxf/VVM+YsDY9nGVUiqM5MNJil3rqrWGJr3HFoB6XI969DH
wc7sra4qnEScooja0nb4KZ+5GzzVHdLXSJDeHGajBjX5MsC3joW4l7qV0yZD
gl7BbcY66zkoVBoFnodAVlyAqg5ET0wG0FuRUZvDGKfpkz2Nucyycq2ZhbwD
ZVYeKHZWApwwiU512lidPYdIkxW4XtF0GjpSPM8yPmJiW0LBt7L/d+C3ag65
n2tqFw+ye/XvkEzJ4ce3rfxh1roZLkj5w75HvWYJ5U86vHmE2USGahnCFGo0
UF3GEF00JPpbdIq7cgLf5ZrFI1KtLAqgTJoYekAYa8akTb45mbeScVTBjWxS
m1CACNh3XUbLtJj+TkbY2M16SYnry617jfi3PTrGmoiAOWWg6k6UnHrS6ajp
9FKuzJZPHLeIrTpDyXcokTpwzqN9btM7IbmpQdX599YAHcOhNqrr6WgBhkT1
S2LhR01Xaf7x9c2+8qmTMF6cvBjr+vmim+PF3CxWFoWVUMKvYsRB7NPNBO8C
FBV+eXXHAPqYsuZni2fCxsXEmucBwHcGM3ptbp4U6M0e3RfOU0uGg1cdxh3d
Q2JDpf2HjdfQf4XX/7cZ6C7ah8vb7oM+QHxLCW1ZWrAqfP6Obv1UOLQc83L4
+94Lf7WtnLnBSyntYPuAfCbpb0eEt+usKLg1M9G4MHvQIzBdyo59qBVZDQvY
7I28rPk33rvuR9ZbpYHhLBH6//R2/DjLpb2Fs0iQ3ymAMMkANWaE0PvAS3Hl
ctdd2rSIccuX8yyrPhswY+o/8DcudYFpE7KPErzL5IEAAnhPKTxgvXk6dB00
Z9S3g0mpFEpm2/ET4g6bH1mX2cnmG0WOwd5HACmUjHf5e/lxGT//L8X2PFP6
OIGJZUURyN1nW+sjg9YzD9vHhFInhBs3BVB8gBUqwf0Dicq74r8S+fA/HppZ
LBWqm0dCo46teoVfyZQ+d32hRwgEN1bMmVqxAomyoObIW7YZUDDadO8uZcoz
A5BCInJN3/VZO5RaWM/BPNlQXHFZO3IYPQ4BDvS6w6IKxx1NlS1HYBBwro0C
0Gb0vo/VO4cC/Mf3be0FtfsElJVtZMB4gnReN66Z8xydXkh9CTlysKAjRUKk
lHDY2AssJfIIolmB2CdJICwBhUFIJ5m7ujO9XrIP3sM8lUonfCHFwXZ37Dgm
gdjJF0RVqyIHj8KpOWkAFrFJ8g4h+FzAXc+B/nxw8IuWtziapeueSFny9IyJ
afVxN24b5Sgi5WvGGw37Xh256YOzvQtB51f309WwNoQmj+MuLR3sA4isSw8Y
OMvyQOzJrktdhy3lSAWG20th13ZjwhjpkW6pMqSMU77e5dxdOAlgmi+1JeNz
/82waL0j50DcPWUR4sjoIJnQoIKHtl4mNeQALkNR2AVoy4M0qQehtlP+ovq5
1eeEgNW9CUBY1GwaNOjpA0TRcAudpx+0vhYhcBelsr7O2Ni+b3S39g0mnBXh
uYrklbjHaaHI4Wzk8XD2Y2jg2P8hZ7YXPYSPFm57PzJdoK2N/cICrYiALbhu
SDb8hNGUAFTM9uTROLMgppWByKdTLrqhyD5npd+apba/6WaPhiHSIbJ6cfxZ
ecayQmM6KyYCxwlGY5zpRSHs1J0rurx6EcJ5ivm+gOA4ARFK91r0smR+5p6m
Z1Ch4/jMB7RcC+L/5lqSpOVcnuT1f/pxofMJqKCU98aj1+F65yHnBMnXRj7Z
kG5rUEpBDwWQQLappg1PuQ6zMiOKyddXbMXEipUkG3XGmwjH9cL554fw5kc1
8UpiEv4bp4ZqUzNiiDgxzjntw+woJAYOeVEpTCa+DNhwty6lU6YwkJ2YCn2C
YAFIBhCQv3hwKYv6TAmphbhU1byrYR2A+j2ai3FOnbCNE2xxHQ1tY6FBrhnM
TypacRvmQcI55/yxS6LwH8Q3XN/5fE3ulaWh2xVi3NbWEuvFL5xrjK63MLve
fiC7Tc+et+pGhoH/YcDTCKM5ljH+ddm2xbdrRtZYTZl47tN+mHJmxrx02icA
/ihLVdUNixmsA4H6Mhn1wY5R0LJg9fqA3hoS5gGNbpDgzj5v0+WvNnN+wevr
gkZWgd5mUFyGkmtAn3wx6Qs5IMTC7JNbdrOeVXaY3KQd6ldkooXkPwSfwr3E
CBC4x/8eqzrnDFqVmq18IRv2XQtgQjUvXfrv67BuBz3ktsqBb9WRb1SkEp1W
5R7u2buMWIJX4S41DSXT+aU4kt5hvSFMzY1xnvqqxJR75WM+4D63JNuMDka/
bwsOmzsRr+FpZfMlnSMWQBGx/0CEgD0oYBP2qVjyCWUE+1qh5r+d/Gy+Pees
XK9gYoVFKyh3SpJUwlpOrg90sIu89/w/gaJvIprGrLLA2YOAFzGyOcfrK76J
MX0t7VEi8q3m6qc45PMT7Hxzdx4mNG8h4OSKl3FCHTt5bhJmpxEZVmG7bMpp
p1DRg2ddMhf90DRL1YTpFQGcxkdSqJ9LFIFYVCIPcbdDNhvoIvKCoNZxb7Dm
STYE+MaIj2+VZy2msSuoAKvmFzMoh5zXDmGUJu6BgOjAYZgplXGlCONVCEXW
EOzTuiyFEBvbHUMXrQ44YANQ9Qeyq18DTA+GZIqAfJ6LVDtEwNAeQKOw8SqS
AZKZfqlqmQtmmG7McHyshQucFhKkZwrve3AthKw25hisDUAOR+QEU8N+EclT
PvMmXN7zSsj0wuxU5GquQdktYSm/4TL3cmUTfvXJoAqUI+uYw6gi5CFN/XX6
WAlNNK+GmanhtsoywVV8+HnAX3uP0V+DAvHUTMwaFVxLHz42n2e37Gv/EZr+
pP4+GMg7TsH+Wh31DopUPhNnYRi9H9wIcWaFyZOpDrfGLiNjpmvLrcrha53L
a26G9CaWw99j2u78N2RqGabIExgXg3+zeaI9AEPidlBG3rJlD1IHyaK174dc
EYIzRRAd0KH8NvKT7mShNLHhJZk4jrsIxjyzD96o44VLeL7lAFbnVggIChJK
IkH6lgrihQqWvr1I8e1xpSDRcejLsswa6oDV/s8OR9WqXcPeFvOpLibnBy+x
oVNnZoyjihlx6DsYGP5ANTTyhJx2RD/qzQ/olJIoWcxhANEkKDEhMDxoi4Q3
BK2Kb+/uMlf+c0T4KdrJ+sxQ6rvmVPyy/HzcSba+poZe9AFPncl9Y38rTl6c
icenFhKcGJyjCBEJ179OD0r6+f3msBGw2u5HtJ8VFVNZc1m/AGo94cdJ0lGI
fPpSt3edLeIsGJA3RZi4qtKBT88eOIaXtB/dia2bWwM38Z09mFxaajf8nTt2
ZPMRYC/xGPizBAkVs0sRMbFaQ+v9kxIlAvut7DWfKnAcAD7Heyti8Y3sOOT+
CETbWU2dJhPeyz+nnYnl1hOjN7DiIX0VYSP4ttQG0Ym0cSOwSPcqsyGMQHi+
c6EkoZyau94LPSNgZl0kcQfVTv1N+j9bWToGxUMJUedEk9Bn5ezbTzbTQJrr
xvdpAJ4O49Kl2MexO07+8dNwTAnxhTil4KBsNzpxNK7nR5Ek42LtiWk6NcN5
WrpmYi6JL71u3yCc/ndgS5CPEtDjxv2Bi6kEOPr3J3ywOOcA7n4L/PODmAVr
x8nMPDu9TpVxfPq4lZ/v8mrlZ1+yyWmOkpIxA2CoIYI0j26dUlD6TCHlVGTk
DrGDzOvSUpAdKjXZuIxyIk6Zww4ZwG917zH+d+L2MNlwic3zzs+Zbhodb5/p
QMIWhhqDZaL/eqym1vhH3QOQsR6p/KU8rAjkYxKewwum+QNuT69+j81K3QUA
6Te8zNV5mfxyY3NfU1SQwEHfoqXuh/SMV/4Iub/a/JLatHT+pOSyc3p6VBe8
lJcxP2zf8mPflrUpbu6xo57FSxjDK+mZHEOyOfx4IzGXSVXlfiDcKjjKz3xT
7/heimBqVLbhL3IZ/HTgiJawSjvJPma2lNQQGIWimaUfZef86Vdp//rvfnbh
nJBwrQYNcvyHEt66NSwfULqGhRdapX2QZ331yml8XQ+/YIGO5Mwrn3fKAANZ
jVePQV7ei3c1fijv03sOAm3sGnvgfbXqLbuEMFeOVxlbrzT3p03jSDaH9CrD
qRujSx6zuDxk6XnuA7bEn0KK5qxaPsOgVcKK20dlOX5CJTkkm41eNaVLKorc
W8TpihgVFXwGxA8qUgExsnNanREgM+aWINIskc2zkfwf/Cr4D9HOqBWg5wYA
HYk3/2tpdUhT9oDMISh4Gep1LHceWwutcuKP7yDefEKMPBeZpTTRr/SzPsiA
4meL1TWbaJrHRHzIQl0BpELgHDF0CkpBr/FaSoiw6LUomLYQlYJDQAwd7KA5
Wjir8S+bpT6bIuGWypIfu3K7/eHuYhHunLtxTd8IkUG19eEgSrIZGRZ6kwDh
Js8gPK90Z0U27mhhoXGHDg2tQeJoO9DBbUO2WzgxxQeiEDtnc1tFOXT/9lF0
z3y+VUOxWzv26mKnvXAK+c7gA2BzHZlJ5XSWIcOgB9D/9NHeeewPZAqyruR6
Y0WcmGTBILcd84s1GbBfodIOwN9O/hnTasTkZgFcCyJddNNPEmAq6HVBnd/v
jq0nEssxGfVx/H2aBUurRAa/TVN+clLX4IUREedZ4meP4+OQQmBgNQ0njyhQ
NPFYaBNRjMrC2vqPZ/Pn5MQduMk25UxdbsnV1bWyQ1j0uPiYbMWxneBtSzHw
8ODqLTmiNx7O8e7F/4/C1AlLY+sYrvo0kd1Fu7qgfvA4aQ54WA3hS+uKG6Mo
JRTrVfpEJMY9xMA/NGug5ZZ9te1WlSMjYBp0yyUAQNzgrYS6l4WvgaRANywV
LpXbYE0xjUuclD2Alo6JkyTdjEPUEviSfZ3qMgWD2TbsGZeJIOgUBg4n+CHF
bcaIfxUlfxDdzrYZ+sv7CW9Jz0Ii6ov6IK7rPYrCSh7+IjnybeGnbXn2t8Zi
owheODno9/GB2iW0lSo9cq6pwf3hpmZ62JlmioO+x7TzQ0Tc7E5J8yYhZ+oA
upzmc68yr3odZ0bRegv0eG7SwdOikj39wwur//s29YZFsA4IEPAr1IwjxMD6
js7vUetx1Ec355Xf5hqfcYFei+V0b2LG4n4bCrdriEapSxqEK1w4ucEHm7lJ
4REMoKMLFPucycuZliF3aCxjFFdPDVceDK4bsxrNJMOFJkR51ofgUYxw8hOI
hnzwSpROWZnmM2b0HlAUQK8CSvrtjf4k/WR5HbD381aAv1cEnQ9UY0hg7v35
j2kx3FWuaw8+0fkheqcv7uZ6H0Ld7QYEnvrAFhv2qj9QOlOY7+QfMG55Wg4K
6b3L08qWgMJgvflx8Duo4IjI/sMr/YyJVF7GatrvPjtiCZpmf/R8Z90TCaBl
txVjfG/hRiRvUfFXvjbZKwnKZNDw2CJf6/866BkTBroN8nc0q3A/L1b5c3RT
2BYKQEhdWeUV5P6w7PvOWKj0GSPjydli5AsF2zrunseDry79SxbcYi2o38UZ
0oRxRKlDGnyX/saAunApnuxf+VOJWnuMTzj0oRaM0qGGxvNYs9hTfIj73SrN
BIcYyUdO8hdHg++3re4Yd/AQHcmdhxbULc1Ckg2ZzDVuGokHLJ8vO+HGKtyZ
iZBQZki7c7iS+Nct0U2aqgI1yBxiWnOitjnX5bY/jZIlHeDNMGRvA7+OYBfY
IxZfHAVJhsb4ta5JpmnHyZ9YaoiRqiYoSMEz6P68OxXBNSl1bWiRPJTwqvKI
9gZ1qgkBsg+k+j5tQDkFm7CA/jAorSZGcEHnNO/GhuDnzj3GxnEyf6bQF39M
1zWP36sgl8RusoaLKqfLeDqlRSToglYsFKmYONGXCQdUn22Y0PQCfQaAYgCA
sEPDyZ8E5E0gQEfc7UWN1/DzKZHnVM0MGzvArQmZnzsW4ad8Liq2x/nGiCnI
e6QjzMpcpQIpe8fdHpAHkPeA+uZ+hkMv4eal310ECw0J2EweoqKWvbzxHOji
4qSfS0AF+neQR+QkbT3T1AeZkIwSdluPHVgWT5qHT8KmHKKrfDAFBPUnmQTS
oznC5ecNA3sUrG4Jm5gbuBah73RB3+g39pkLwcK1PjRTZ9OuWaRpNMEELSyW
3g8IUFhFSoByTZb3S+wzXY3wtZJM6IYi064T7KdJpo9+zC7TdY0w8le9F3Dm
/OjVI16PBTgdOE0wcp+PJEjwfbLWYjHHvsekQ6aMC+FSaOockOCVIQtFcPug
Lge5vQ7gxifodYB39t0anitSrFCrzPa2JRWP7xf8y/A6DivCKD7Q1dd1XmHZ
C4pPXziO4wSkC7Z9Uc/zJKhdcAfYddS5/Q4H49V9bMDtuJhC7Tfy44Itwz5K
z4sy7+BeT/AVTIQfV3rEY7NkOUikQr8xyugZhGzoH0aMEFjeW1uM95J5G2f1
V9qjauVzF+i066ukozMILhDIkQ80gVYzKfuKgvhRf7EzxnwOF5lAxiXZ/4oe
o3EGKIrR4PJf2HUWiJsuCAyqahjG8rE1xby1K4W4eqqf/Ckg4K/OnpP3UwxB
vcxUeU0x8BKYjOvw183KtzDUCd3H2lCkdcLwrNsooMAlcVzuKkWFm1amAuYu
l51nbBUYU0v1MH2ej//CuPrAvTlCaFNJHZTyyPLoGfcTGER7zNJUMJlki2/F
9dpg/ypoxrPV57MhG7gMuxXMZKm/KukOQK3G7jfkPzVNZal5/Mt9BLdpHtJU
sCXKRkdnYV+p+ZWgmDB3pcO0qPczuzjwsgDrZNckKVQFfIAvo3Iu5aHJswU4
IEuJYa3eWPjahbF9p/ZFS9VdpygZavLYzmvOCfySvEvaPW/gwbqtwUqdtKGa
spf0FDyqDRpyCckSYf4XGo/qJqtf4d7fuUTDqb7FIj8VDRQ/6R4gkX3dhNhn
0FhHL9fJIWYhSFSz2td7imhGb3DgHcWDeXfotAFmTRlR0kKb6Se/gzGuuXwb
e4GP84gfDHCkPxX0LAzEjqXGfdUEIMQ01wvveF96DlNbgbNXf1zZiOOg9cL7
6eRDAmr/bHsmVjuu7GqE9XW8v2aAJ887oJjNK9hESbdnKEHbAsn2RVTaHdua
frQCW/G7wBU0y7+wn/lLp77jxVFy8o1+KuoFjSGrSieVlg7fw89DhXSOYbTO
K+nN+MW6MCwNrXrQZAVNzqg/8MWoZzybKugjC5fkwrGDYUjFon6ul43Mj2QH
qzGDkgJ+W/Lrs1Tm067+LMTLT+EEiTWnoLc9nL7HAUFnzNsWB7Gd5qiTX8QH
HJAwe7gCnKVc6Lc/SfpaC9rrzjK+OI9nxo2jVpze9dv4kgciptOW6LPuOgep
SmzbhypsCjhJ71gahZEYPitRk77L/wKyvsmnfdeClHNVKO0FSB3G1o8MeckG
nWpVWESYwUhGDJb2xVGqRQ1W4G5+77EEyxjQIcoRcA2cINatAxXIeM6jUf58
m/8E/87sQY2tAoOWG6qqtiK/9lGEH70Ajcfd8uA1eDxkD6tuCZDWuy6/2pQs
UJEuAPsJ/pyCrB+xIfuDlOolicyony5mI3YQQt5DHqAOKGaZWPK82e5tBD4T
C6OKygzu3YnVYQ6JTHqKtzX5J3fie6Mj5W0sk1AH6l5z+ZfCgAcZaUNQpsVn
EnNceJJhTEF5LQQhVeqF+TPT0qV1Y6rb2Wt0RGU46SAtKnvk+W6h4kwjJvuj
FyM+LHjUX0dtugvpLW+maP7AM5WG8JU7p1L1PoHc3kdkl2WOP0g5wfkVaIeX
1osaIYDXRIWO1vb0j0h214OXc4UgqKJWANezo8mUIWpaBipJAMQ34pw1JNxH
TwVh/hXbM6W87Z2hRe9wfbehcqKCBMLX4VxWfbk8QZuC8/iCdiJv32y5vzl4
nM8QPVEVZ16kGTwNpGc5wOHHpFU0uZbTi34u6GIpIPeoqpSaFCRgi+CnF+Th
mWRwp+I7N9xzmnFUpFk1IbaJiy9YZXzwYGWGreuJBSFr5sk/U2SuN+GMBhFL
c16lKKeU75XHrQVJpjGgi0oGHP5B24+za3irO9vIsulI/A5aedSlvEA3cX9r
y13l4N+WqwDIo3nKjijFIjnjZgZFs2n52BEpLY4koPQs1N1AKHZlr/xxweSc
eCuWVUnWSP/aBeQxcbT8aOTwRyRhbIATFhfDy02jJ5/jtveAdFSoAHU3mfKz
7a+YQ3ccyPdk9zxWBLvOl/bWz8XcD/Plo9+4Y3ng0P4gDUkkQNehCpRlachQ
ibzsFvbtJzMZCDekoPAVzJK8iBjGnd7XkCMtrMyCWFoIYd8S5llBtajYj0GQ
HWzkqyExpWPwGPNnEdZqrAinhSJ6y+g5NFM5izHV/fiy1FcZqRGn98qOTN9T
N28P9fF68THdI5PUAQL+OgyoH9+IdtfbcZwQxxpBWk2bSkZpTotQOZ9hHQKf
DXP2cpEAnbFuh0eRGxaNYjiIjdWZJqng8+QLkkBEiSiwckto9IZ69wsGaYup
kweKStha5HIGBTSyq2UI01xz/jnJpwgj08inhL+yKi/Qtho9T2Pcoo9dR7Rf
8uyz0tcP72YSq0i4w3Sj6JxkiPhprjY+0Bqay9Yo8vAnfnA03plliz3X8ZWP
4dl+JqBUDI0uN4odRJzgW68aRc+wZZv/bXzlIiKWE/b8b7l7m6pXgdIFpjMH
PiCWI+OJ7KXfIBEuGkYKIXFTbINOFvvIncnHuyvknwBInkS5wJL2Baxj4rFs
26f50K8Zai77SpJbYtrcrPT8yOMrrN1PpsGkCpcnZPFmCDfZANC+8BUF2kIR
IcMj+AbEqpMuYHSd6+ozFZukPH1FazykSjwpo6myNnCm7cKIYUnLoc0X51yo
N/ATIsASxt01mmgM0SutJ7AxE58Q7vahTm4ycYlRHqWMzJY62YehJCGXio9l
zFqH7SA4BmhrnJekDeOEywpfVh3ipBHnwhMLdQScWBiq/Zw0N+JkORZLgYdY
P11g6SE3KTitsI+H49RV/fzTWFJZaSmru6S4j7ZjQwklY0SDIG9lUf21q+Vy
JM0zZECH+qdwixW0HXM9D/gVPz1hSnCKiC7l9Hdu1Ca8umDYW8n3xZo5mep7
XHy/YFbtAxjJDPTURBjtqxUlbb2ry+dU29nRIfbsNRD2+KYpnYVL/817yGpP
2z25zTTOXVANz6PG2rZAWOY3fR3nwOXWcDtOaDt2EfnCSH5LGHN4u+ggTRuf
MWpKXJhG+Tmi3lu2Vm/46QnXSdLXxlIqcB1MzbSLNk9yVINQm7yZUw9Q1dBH
oLRjFC5h5fqXRUHln0DAwdOJZZAWwR7A5ExNEDVm50UDUtW8mcGVlX33iKaM
SIbMRzeW6lpF5tNlH3cgpmoNVQnK1NQpACFuoct9/66/NKHl4ThzmPIMXNuz
ygvQscZwdS8VGT7lvii5MFNEY6FJb93aZNQMAzwF4eRUPo0qtTaHdBIy2OI8
HDgym8juj8O/dyYhEs8c4Q6phbrZ6QD0aAtY0MfXlg9MZnrNXFHXRF3ybpDX
mE+p5Ty+N7VCm2QLVjnVlZURYHwW5t1+QfF2BaCf+P5qB4oYXAwvnvg7ddEs
kMdrBIwfYuC5vkbmeqY9RNUdtb52gCvpPjRqeAEEKLlIQdv+aIfKSIBzSYDZ
C1hM12EJoygBFRaWtQw4B/z/VPrwq4OWFAMoJuR3EToyLErF1BaahUjj7D4U
J+3tkVKjfA7E3cMBeh1P0BkSp4m4otR7oSaSTLmDg+JTHb5AMEYeoeQEl5zH
5yebDtBPtFX9evUFeAWP0mMgS3zPAm2IPqKtz5XKY1xZjAqBPUBx6JrfrFvJ
O+ATxm4vx6JU69UOeOVXk24L1LiFjjqVotPsVZLefd5zqyCBTGK4LB/nf2cv
EHnfvA3/ksEaLAYW6P0x/xPyR1TWKMHeZhjP/AcSqJylFVpFRCUzVhj6fExP
wG2mwfIBRGWEFiF2/VLqtnvLMJyGCZsE11nHSfKH0D86z3Gtsz+16m4MzkZt
4NiFzAuQTLlYxn243IsvlvIY0zHUmtauVQnGjWeYttV/d0qYIIfEsQ5Ph/oV
CrT2+C2Y+8aEY8pdPSaBLerqBRBX/oyqM0ztJ3v9RqYICdd7V8ohnBWC72If
OnrWjRyNlgdONIZJW//JPIuK6KvRPIgeq4ZakCW23xCeh9lkQ82FOikKy75A
kzoKICDLV+OeoBWy3KRyiyZyvxA0fxjMynyFB92+YKAzVHIDRtPsnwxpZw6e
RzpVNg7Fkug99NFvmrEU+Yqz0Zg3LqQIfA9eNOhb6UPKA8Q78cKZ3TWNmBCB
IpHSp5kglfxny7D7P5C8GFOCLp+vG6EOPF1l5CuKyGKhNl6hj6q7EKpIDj+j
WB6VgDI6V8cBQBKWEGyt8bhezWe6AV6E/yl4srRnqOmITy/egDOW7gWOdz6k
t14fhwFQeE/qvy3RpL1XZ7tJNwg2mcc3n6+GbtiVN6N05jVMemDNajYKRT95
2eL6tWXwcSyuNeRY6k5ZfFNAoaHmGniukGmXJOFo1cZyUAhBClMQLFm9S4an
q5VbmEXfgHeSjuu4ueFkouxyxy2QE681Dwcn1UU4Ap3iQw+u/r4WKaW+8pty
yowfyDVHhB6rXKhx5VB9o0azlkakq3e4mCat5Xut38gU6YweyzFG4xb/BtCe
HN0ZDkoO88e3pzoOknFEe1VemWqJPmEK9Z1FpF5XIWeZ9X00MLKuwzOXVt4A
bufxIresXlHd2RtftM0WkZr58HWxfv4uMaR15N8d73ozrW6syIluOLFX+tAu
abQpAMrCc/fFVqP4r14AIqhr37dgz4zk9SHYr9IdXejpDi4IVpJdHXmp2ahF
7WCviwiWJ7TJ8l8aQhqesB5J4klA8Q/0GVXMMac/NcRED3B1eaXti/h8gorn
v5naHwdNWH9G1wJ0kxqMdi/uKt5eC1eAX12cTxegImn+XPHRjyfsYanjczSB
q5fAn92KaipSSiH/pu4H/txifN0fILiLgd18/0uMNjs0YeoqMui/dyI/F9QI
Zk+CTaYkliOzi/8KWX+BvmwmlRPreun1RfXc1lSNeaVbSgcVfqDLIt4utk+a
E0bnBcmPXVTvIJK60Hdzzpe/HgRAl4rR0jh3mcUiT+eDSxNwVwDT76PY2+g1
yo3OPc+ECBHPOhwW9Wu7asLTRsL1VEQx6BAlbaRAG3vLgYB9LpOIVD2CMScp
77lfsS+/T1UqYDxPjV0B+7Adm8ivxe1CzlGGV1KngdlzSG6BIVQ9B/GJ9vzz
YqeH0i/Jl+tgPTLHJVnY//g7wAEDY2g30n7Z2Sjym9RR7levd7VhIKACn3PH
P5CIwlKKIlontz026+xDdLRbghfK0Lhgthml2izXyEDjONoMLz2HzVekL2L7
OLhCssCfYxAZoC+c1OSULlByWB1+8GFeHu+2kWPW2TDmKChjCyz+Qjv38CvV
SvUyR3DOLEO1ne7vrzvBTaCcCm89Scz0wCPkZwNGksTCtDedxbRaR2VXSBbD
UKnRCk0qaLeGbyzrUHOR6XT6dwBfTNHjIC3LyFi8TsNZ59kxs5g2X6N2lCNV
7fYTAwZtAA/RlfSUW1AeNW0hGGfuJADlQvH+SMVhy682Ss5TncUPPeI2CC8q
1S5Jpr2WxaZLf//UjYRniS7dbTxlhYF/exaKoDp881RxjMizkWOFcHn7EeO4
D8eM66boTznP51npsNM4/tqyLKK+zaAl/6N5op9hVDyqScpZG/V4xPt9L5yc
9v3fGPdgg4W5/sLEWJ+NAPPvOXhXjT96QrrvkVquVcxt45VYPnr8gWOZ5qqG
NftXXiWRXlivrJGYErbABDpBDIr6HsvlKKjBqrsP+6RCj16peWPU3OWxtQre
PVufUh+bMCiPNRFlZL3zNJL+X/LsraIusjz4yfwJysO7kQ/cbpheOzcrki5W
wMbWY0thRKpsO0ze1rRE6ve3+YqBx9+AQ8sYjg80KOdyUNahaVp4v7TMYwks
t/SrfArdmUZBZpWCMMM/18ZNCvoxw49FLkRmZvxUCSucHOz8HXlBleEeyU2W
kEs0YfW9FPfQz0IDLaATxh9K4GRxyJs34dMCGlW3Ob/d9FeLlfg9WBH27vPt
2Mb810f9CTs3Hg/ik+ZsYJoum5/YYtdLYriBHJdpAWnyxDOV8YoQu+K6xaZF
klESlZcHjH+WJ88XFbb/lR9Ie3NItmFoR4yJiAI1Me1aVdTRFt0XcG9hVuEu
IBPmTQHZvDAORQV1/B1vswJBCVFqAQlhymh02imDhpFUW8k9DmQMJGtNhltu
8N16skOWVn18YuWGV+GA5NigxuuFGAVR7lMjYeHI+jmE9p7RtDRFCN2WyK3r
UtNcedi8WIBpjyIj8Noc1P9EDBRgdHLERNz1ZtaxhE006AlW5zencZUe6Ano
LvyNXKFyjHnk1q8dXxwwPHMnArWxjDY2BoQYgCiDEIdu+Id+P2elLToGca8z
13L+/6qntQMjBGDxYgPQ6ywuA0gj+ABOSZY9eXljKkQGtmbup4NwoGzT+yHY
M6wh9DL9Gn6PKRUY2YXCvEBMrAgBCoJzHhZKB3l5h3iGqtSkeszqquSCAblH
KpUods2b+fFMfHj6GZpio34ygrE6iRXmA7+TBRFDf2/1WzUGeOs75Sn+NwVf
+DpLJ654j+9udQaBa++Lxigy4DsLoQDpNCJ8WeiGdCz5iaYj26Vh3Go/EkMW
d2Y8jYlLdle6NlvHw0a0MjQ2D4p/xbuktP2511ofHRuEba27bRWQth+OzzSL
PslqN26G8JD8YQpgPC9dCnF18QhOj3NPu/+Y1KxJFK7JXPdeYUF3INUehIFt
abE1gzOSi7a60Enl8kxoptu/6SlrIsrkofIh98Kb1vB36/zgczjDQd3AOCDr
yjOWBsr3Im8HN+z7lualbYaWBMP62mzJB0uL70YfOUeZ1atfzDY+SbMN+ZBo
KlWTtGMCxKyPOIZiCz6+kLgEoNA3fegbBYLrOgO58KUI5EM4Z21J4HBuLLCz
bM7IvYFA5nMDOneBNLD5APK8usOxeOKRDKTsazxiZX4U6XpH/GAfjp8NUKad
7Rc+i4bbMf5+opc8zpLGL345YtCDAqX8OaeISiy5IjAzBoxzAJcsQ9MZJpgw
7lajF2RQJsvrGO0pXohfDBJtm8ariXkCmCCW/+iwlTTMTlroPyqWYM3brdNj
TF/o0tXKBXnztl43LfN+JPmPZQle4uIBSvgBVdEI6g5DY5+/0rIYt2D7yXHd
AVgBx+1OPV46tmZhQ6yhMtX4C7w/7n4tedP0es5iCH6OCNmQbdD5egyLYRwG
Q6+PWZXjeHABl2HidgWLQrB4UP7Inllcau0xvZCeC1aMkDCvHvNHXy7WYQPn
bkbE9jKw1pBLm1s1ld919iu+wTq+fmk/hSk46aOV1A3XJ+I/tnrQJGcA9azG
MIHVVH4y70FBRJ9FtI65vitmAfTl2EQfigiD+6KUlK0VyoASAo6oA/JSdp2U
49SOxfxyqQhzhazSdlz4xbJ2vQ8+0u7SJ7+MYD0Y/Y+VXtcvDOOP9YU94n9l
aJ9hSE+o3xMSVdQ5VBzo8EGHuDdHxTRHerAVMwdYwI2tOM4SGMyQdDndagh4
P3zY2PhvaFAZ3T5xGAiBgh7vtG66dCkvAXqXE/kuyPsPALgUF2XMBSbOvjqE
EyrkMok9v70L+4+H2ymLqx2c5TvDlfRnkT9hto2doKkGlgguuvRjNVF4nCnh
JYexdkGNfZuVD6hdfNjQ/kaPMlKqcnD1DQA7gCRWe/LqC9B+WKfZgCiEGuvM
D265mKGBqxFaof2AqT4FJyDtJJApt4qvnNfrfB95KN7qyWPQAmMf1k3E0Cy6
cMgSZ57Ocfxm4vB63V0WlR5gMPs7t1p8Nj3MSr9N+0t+26Gw2rVx0/ewPjmG
9KpwXjyKpynFRXVXMQMvboSrvuiPYvItP2VJSRy18rJDMTbr7KEl4wA0LRg/
36jq1Bu9O0a+0lVudWF4RCYQMqye8wboT+fURcbTFYbYVJIzt3UYbgkADgwJ
pRiuU5dqobpmqO3KQp2zQOz13OMw2Wu2/W+DnE8/Sl0Bp5v3u7EZObu0bL2I
RR9E7yDSDHMF/mJ9sLQKFgpGj6ke/fRBUvQpGvIgG3SnRwVGsU9ak2WJYAOX
qjr5BbVJsD8yQ96+fie2URWoehNRO6QTVzjMqQ0FLpDEGURNxdbwkedibuPz
z6VQaMGxnbVgydl3wa8EA+UUMj+Rohqaitmmwk1KG2cPxwuzZnHGW6cWuAiy
nkWhF8YmwdltW+pfnyDUKpouq+tUExVWdKMX6jaaqi3VVZhMcWirqbi5nxaM
vTYMpiajhgTRpc1nGr59T4KoQ/Rn3jtG6jWxWoMPVHLCxVZcHsM9rrZW2k/+
JXtf4PoG1tDHQH9LoRUtrtR+bx9vbpR0KvPk0Nh4eY/mEoq/xI3Veqm3WF1O
mRHdjVsaXnOiA0XlFte70fmJn9Qkvj8crnhEaoJvlVhezsOyNcmQA3OLYoqM
7t+gnEit6vrBt9CVGYN6tig0ZscjL8CwXJnyeJOVhPjgr5TqlEFQqolHr2Pz
Cqy1SiZk0PkFgvuAH9cEmX/ic0nja1pzbvK06AjbcC2robGdkw59G9pxzEGK
3q0K5HG6am6oXd4x7ZoWQQIOnkTGCiok2qjnYtv67hf9wAnfWPxJTVRZnl2H
nPhV/pyrsPY8yqUEPIjszrKRVsOnaDGYn3Wy15l/lEZYsBX/xU3nkkjh9r3s
P6OSdUT5Y6AqcbGJHFFWTd8Ewi+gbIxEgyqFXsEUbIgnTifLpDOgxatOcgzz
iVW+MTAeetrjM3OdzYV7Dr9mdixLVL+4KL5rWjKbOhKJAnaFP6oFYG0U1Vr5
8eBKU/EsVxgzMs8S/Bos+Zeg3sr4U+I6BKyjVa7reTLmZErIGfebtdxGHn2w
M5AlgZRYPQSRE1yHcm6DFI5EXDmxsRr7P6nRZtSvmGOK9vw445WfpnrY4Eik
t3N8O44P7nThbwqYEIWnhUT2bQw2x7aw2JWSjybiztVivnwmM2I8RqM28oNE
4lk2SXWtOjFTpKaGhGT7FqaOnNzYLsUZ7PxgqNbQZ3+IbkGCalSXzi/1MM/1
jb0fZ4o7r2cgbyAo9/120iTiIPBZ+iFVv+mq7CKbEH3HsWT+E1Medb06FqTp
MrJatW1GZDv6ltzKTdwOBvU1RtYsJxefbfMhYEw3Ld2hMdWrkMViTFmiJlWh
ZWsTu9XNdUI1ytIr+9sJK9Fi2MxqBp7ohqHA/A7fLKAys/OnuCIxy6YJVe6A
qFwy5lc6elmmdY91hLIGIcKt8T7FbwHC/PiwcGeUrwo2ngKLQxG8RFodHgNY
YuMK3LqEEI8G1qTlkPnVg3DsMYRf3BFWODD0Lxmuf8KUw4HFhf4NAe5o4cQI
p9PASA7FPN/mO0M6Vwz/rSyY8bgA5MGEwQRpyLL7NJzecqX905nNnJadwE3z
gICXoumpCWDZZNhvpQhfM6URUBT08ywM5S58oam8oy4stLkS79bWwH215DGf
60lCRJsb9obYQJkEtVxuM1rGPozdbcbo0imjeC3qM/sS+XzVV65/BOp6Gkza
WwgvtuRtcHg29K946a/M1XvjiYY3PpRlHBPv5XeNDrDi11ODRj42SfBdbpZi
okc3K2SbEIWmEDJCpS02VJwJ65VGRIVuz/0NEE4bDTclMAK1oz2QCp2tWFCZ
cZKb2RgQz6IOsTScNOwDZeynP7Oqu/Igs0aXG6y/EtaH0ZWcE6KtSDichcWD
X1ugbTmYYJQ9+t4Dh+LQTSzYCZqn6O5CJr1KS9O77NLTSHyBaH0z26AzTIPh
rd1HaIthTifnXCi4eX8aOTaBEgQuCbZwF7CerUZQXIU+Cbv+iDhJO1Kc39n7
qG+DRyTia6P80/i59700y5BM8eqcniQAv9nWSJLdLDz+bXun7GVQ43U18To+
2xG87CdOX8YzwPxwYgKbeDbyOMysxJDqmy8b/FR/Vn+iwKXPuBKwG0gk2UAt
U7mOVwbdEbvyasGe6eGfLvRIt0N3SYQwAmdwv/t5mSYhZpsU7d1Nd37cY3Vu
4mv9QoXfidHku8Phlbo5+LfIwvbi8ojsq7mG7SdlWK65IB2uWOcv4Bczmi7N
dGm/nFgWc1+XpfQZO71OwpRlpb2MCQ4UxgJNTVEx//MZtt8QhZKxBLcEte5d
HeMo8OFQl3Z8Iyf+z80FEUev9n08ACbEP8Qn5YGhf3vgDsW5FIQ09SyGlTA2
nNpuEP69sjyFWNWLcxrSUEsEt1O7uFutHOqCn+l0iMENrOrLn6Pbs6j1XizB
DFgsI9Q78Hhud6XXAaNpR6HXAYEk9HvH6VWH9DTEy23Nt9dstIU/32E4yyZS
C5hRbvPmFmImBHVrcERKntCBnJ/CUmDU6oskH7OcnjK1/rvywFZ9ONcQxCcU
w5uCAlv3i2/jQCBWR4G8/vRe0yfKWnkwU9r8kw+nzDPrN9O4Uuq8OxUmYLM7
N6MVqvF/5B0uqcNzm6mpc5cZr+IkNc3e5q7iLKtNKYL1lBu2U7eAyGRX/ZUD
bW4CwUNls+e6X0fddlVqkwGaDu6EOAenM4uSp3tgsxDG1RP3bkmrS6EFLggv
CtyVwEbqtoSVRjB76M2B+KHga1n8KFw2rzKW8rjJmQ055pQwDm95p8X4knMu
EdJ73LUNxfzz39bE123sR1iBvTZVdgDImhWDhLkgZ4SyKMjy0N3KveW53ciP
OiHiTMQv9OlpCyo+vicYDcrTd9/6UV8SdCQOQtnuXI2I/o2N47Vjv5SyZdRH
kyLWthZEBjjaTsjKDsLaqBJIX6ckH7oRrrhhg8OjBys4BIjsxHtq0ZDqfWoN
qZsNwsrM320zGsMNEIlSWiWWZ155Yn9CIMSS6UCy8pFFdQLCSiCr2QeQRLsr
qcxAO4D5fj6ednvdee59PxaGK//TTSLkTc+DnDb4RyKeIFz32lq4bwco3ZyH
Mu4MwGvOUVjeQ1+o8S9wKb42VdcjPEQWSaui2K4ZrGsMf1XlZveoHRu0PN9L
GmeJuwSdYPrztMRXIrgqpY1YWbmn8UXu+KpSFobzC2DbGXL+4GNhhuj2drrQ
YyGDAkg8yrUbc8dLdC8fNSYqChFslkaxvrt6/OCYVAh6GWO1FhciuqTk9V7i
VQx3B2OpB2lZ9+YCafoPps2jhXkTlQ+ZUVKf+RzuhfPJHQN9WbjJBpBSvfSe
vsQG6MtM2QWyY1UvDdyfBYhZRh8JNBeWN7wt4W3pqmhMV+NW9rANpR2elMFT
O+nduCLt5EPSJaewVo39AATuEdrhpc0SVh2TvbOQdaJ3dI8bVfVQm9ZZXtfd
8SB3ReWAvptqzjyP/ji6Ayp1rnotvdHyO3GtFYb1LASL82hiL1CYM12WZl5c
oYa2Rqxy6ovr/IFjvkr0vAefG1J21JbP/S2dX4EyFmqAnrduDaB2RM7B21e4
uM3+d4bMbwvoJux8PqUCxo1fM53yJcza7geOKaqkIYDmClBlGgOmMTtKQ4cq
+evX3OKS6T4F8a9MXBt27K7xggRViTHvD5rMEFva27IGUAyuNK+inRI2Oz2K
tYl+S89a6WpiN2JFMNBS0BTmFjvEUqetr5ZWvFR5g2GL9gAqpUMYEYra8Rij
ib3YTOBVeJWXWGPAaQqT5k+NYSHIzW2PTgw/ZGdRb9cEAC/Lh5JuUOdt6irj
T0aFZH+wkk9tHHGXgfNcE1HyfSNoDLRZyc/s30TWXQXCj1rZov90BYQukHJy
J4P8MWsm76/z7x0nrrOF2yEknlD4fo92jmWt8+NObxEOCYZpfhRJsgkrZZ9R
uAVSdYXf/KY7QwlwaQWHJtZDeOwIeQ6GF/HMqHBWEh9qqOhg7Ih9xddnSS11
QFeYLT12heNcSkJY+VmreC6vnChM15ZRYS3G8BYNNVbz1QDvvZojoAK2EEa3
LUiExJzwobFy56izrytpTmtk1CCBXONY6CDw0b5Z66+658zzTyow7Iy+Q7zJ
wHea1deHZlZ8JAnhtmHbe7wkWraLMtQSZ4SwzrroTkMlcLAQ7gT0j4KWBk3Y
xzB0sWWlxE/pVW9BahLT9lpHLFSki7iM9fZDCj0L9WzARWCQ1SgXVuxypyq/
b6WrL9Z+m1vXUl0PesRpGJ94dnbcgYRI5bzjw1fT0hzFViVaef6UjhST3cbs
H5imT3kBKsBLXvk6LcEp9n8eIBn1xdje0bFC5SfYIue1OzdqeKZYPBwP96hH
02ZDmFpk+0VgtUClzLq97FLecz1wv13k/SkaRhfIMKv73WcCHWamtFOIo3Zk
GJlMqTdq7BUOB3nBa0fp2QEJk6YF3LzjXbcSQ28LN5ngLGObLmMd+6zLoaqF
odMLsAZWkNgwldFhcKPqLufG85p0x8My9lWD2gLzO5Gb7hPiUeq2x/6Y3Sdr
CR/M1X0KMYxaO5jcJMKP516L0ISIZot3h8tG+s/6O+rXPxGCZSOyvghfhHak
1YaAD0y9uLr7QamIyxZBAd8TlmCBDtrsChNO5rVrJmscbGWRG/FsKEfm0EsH
mHIk7IZMjdp9MLIoUibNefajiWu2yYL6GpzRSXB4u6ngljELSjXSzgNqyQrA
3qQSXDFu7zoMvseMxbcPCWO3fU5rTjkBazjXg357odG2n/YSVf2HsWBAyjgT
F0+GxRifDFXolTztbvrspkymE9xtOgTh36Hv/HRmuTul1boxlmACfXlpQ33m
l2/lCmdffo2C/9i+1LngapzEEsVmGD6ETpvUvAe3JPlb26Ms4V115HwN7fP3
aMkw3cX/BROatIT46zcXWLBwfkENmLgFZ1J3iAv60VKNXHX7Fs09ShIzjRJ9
nR3wKKw4CdSJtLVhlyb3znk0yRtkPWFYeGQ1txz5+oY/uDG9F5Yabm45cf/C
09AQEEUfT8cPPMbIaTulL6IZ+IVVa5/jVTyC6E7KNVBuLfMkujb4u2gYrG+A
qX1GPrNIDKFIgEmn35KVhDTSXREYFFPO0YO1SAl5bGlt6gbvHdTv3S1NCgD0
maxEFlLTQXsLuiiUrZvuYgb0BgUyEUQikhIhyrhBp3TZZB7mheenPBX3VxaU
7+4IrcvqPjTL1Mp9gDARFqKqm8vQrAApQnC5UVes9hcqXQBVTmyfhSWDVOTd
ejz5yDk9SIi3dJ1Rk9X8Gklq4OPRt6UU7Ea5DNDGZW57UddQfGc2pi7ZkOCL
aAH5YfI7vZ9wMvZC2rU2Ikvw0yGXA1sJfEY5cF5x/mHaaoHIt2qQCtSLi19K
skALXNJ6zZ22hTWQf2ZDvqZsN3lgwINEdTqLn5T3GtLb+sVX/sarJCuEoemF
xdQARrx4x7m/Z7mSPmQRn9E0Fq4bHBtNsK5KpE7WRKmAgS7ie/cVfnLfgcf9
T+qwPS5YOGs9d8llAUZX+bhLcEm96vbZ0c0jG5oJ5jGxm4vBFA+XpJoAouNS
JElb4JsOTWudGnzlEybu2SUfDuTsWvuxWZIRRQkKwoc8EsrErzHEkKTPQM6O
COldnDkbem0jO7Ip5dug+A8QqlurBHVKLgcxwHoT8jYhGyMdYMPjY1xSiWim
DWRy/jqJmP9Ti4jrnihpKTCCV1U9ELV8GZIf+5FvqwBPHwfsG5QhWELYlKiN
9ro41c32o74yr7/gU5XfrIyvoh446WR1SGrG6whKpnvD+f6kYZ4y6vPS9xIA
N42yp/5eP4dEmAEnwBLYuHVzajH0DQ+cyXgciSjWBVNlt/P+oIJpeoT1dt2X
0d9Qz6cwtytuOUs+RdgcLdSzaI9pmZfMAwLQlR709QwUE0QssjbXxgQZNPLt
aHlCwi1JcZvdJbBReaDfiJX5Vq8oQAteX5Kv9VBAYPl37Gy03XkyUHP0cP7g
ErIKBIZdkcP793mvEQ1rdB2hIpIr/jfixfGtJ9EYpsmuRFOaDbxmUFSUfXfS
2LASQuhsm2un1KpebHUAgS8chTCMkFGd+n5i7931ol+FQUwAtrMW65iGg6sW
pU3HljQ+fs9uDvGJDfMyLJXGHUkRGbridc5O1hRqNQjnW9he2r6Lz7NVViM/
UmaP+5zjCm3gmfr0pcjL4yb931ZbBGejL9wYyC894R63/KRoSKfKkDPEMfJK
dZjtvbp55clQyVM7Ft5gw1xx8Zeqq11g790x3OCDD4WXrQoWANLZ5ismT44j
px8PJEhTLoxCgtrnAZJbwbUAatD+0zAiiyQZO4pkJupkfYaxjKCOIfK5jYie
Y+Cr1isXqyYWJ3l00f6zrZWv+HKErcy4oOWmd1ZA1LOJL1CY1fyswmKHTL8J
Lghbd3sV5v4rNyW2FajrK6cTyMUBK/L6+FmyBmIUcQyIp+3G66sdTKrCr20X
CfQgvK8oHJuObJgMXvsed2yFTu3y0Gu+wkRmticmFfGwbJjH9pBJ4cRsKgml
+8o6Xj8xJTIkzSOJawZa28kmGol8t6Avt5JZJGzPeX5769x3CSe5aBrxNYBP
0p1uGpKf9u/gTCS45Dn3R2ygvAjxk9vQev70WtGOic2dsogGVBUjN18iJ/Vz
lsXoGhh5hCOQRQLgiJxJfBWRPifjoyLxu5PtvDerOsSYh5i75we1LK6GFrPg
DLAQGHcNLbHDsTETGgJb3CxB/mfYhzJZyuS7wsxgPxKC3sLN+Ph1ZzfI3JSM
2B57yXpvLGlkLt2vlEnDyR4D8kE5TzqsmiZbE3nQIhIfhulhFj8xMI21fQ9k
Fn1qBYN9dOkesgY+PT7d7aXeFQYaBUtCsWPRRd8nv1Zqqokm23ghNeQDR+76
tpHpW1q7C4yCbcf8fDr0qygHogj6aHL0zO9LqiYGxGxuplNYzKDSg8/VkbDa
WqtwL7Phc7b9N5HiyYlUhDXGiN7LA8wELNdfL2iV4RjM5PT5dw8Uh0asJEum
lpR9FdNeqrye71iZYKaIJ/9dV+NpeHgEirVhV5Svn0XHMzq3VxAiFJSjhjT3
ks94HzUPyycW3CWzGHeCLffbup3nnXUOdNEyVHUdg67wbnHn/3fitMFNJ11v
hES5CbVvAux/zg+88M8Ln57+j+sUVJ/9fozbnI5+ZttzcNyt5GMlV9cJbf2B
qJ8VfISi17qoBBpqCe4NC1SnELaRNjC99MeAr2cj4esB+BgC8a4mEe2qXqDq
ZMgV+TCa7+p4SkGp4OtScw7/rjbeIaZYDmGHs2ZQQ6sYYrk2X4PmpIdsVFhE
VMfspVO/Uwpn80F+gxWXuGZfW68JyxpNkqdMmi1ZbvZuInPOGdV8xm3DrmX2
qdfGRwMXPhLrNaEo/iUmgfVOommh4OM1DEHMcjLOIx8Co39+bsOaM5IPAYt3
44XkDz/0UDUFgKf3wOJ0+Yj0PU4oKkLdJ1RAfYpyDQBn6+XcMmCU5nxf8Hm1
rLNqbsm53+mJymOwg041R8CQ45cympAPYGRLZy6cTa71Oze8pXonoReR7cnI
y2FdlGIjKqY1d4Cdcq9N7oBpgDYhVqIh1zYGm/OqqENjUgwxXYxNqF8/LsKb
y1lYzmlqLdTWr/U5xg77kiWNmx6u080EfljTnh4TqGNcCViDDXzopL7SK0di
HHx1Me8aBjQaRxnRUWkPeDJsuqNSdnafFcA79llXHYj205zgLRz91UaLni7K
JWRpT5+0hbeYKNNHcm7Yb6MZpcK0u1q9Pr86z79mx0LHDHkatlfOjXvR6r9l
C1SSm27sLV7v8O5Kpl9N5ZJKTMSr9X0Bwan2V+518xHFdwhXmXeDuiGq3+1O
oqnlFK3z7BuiHz9DRbseQBymDqRql4vFvOvEed9lEaS0ThCAfCzav3m+wyZ8
0y4m/VVCyX5EAshri0jjcNORsNqmmjnlr36dgpRXqRweMZRle7S/PuhwLuw1
Qk12miRIynl4NAEUeJfaV5gyEXr8jhOcVxqk5SiJBve4c7Je9pmij/iG+ssT
U/NCghrK7qQkME8BY6smAnanlOt3ANNM7/1m0Cg/8PF7EoyDyzKFUJhA5YTc
n/HmFzTHFfJqtZrbFC2kbZWmz5VMPBLKqTgEMK81LfqIxNCI9w5+lZ6r50rP
uL3VBHVeb5hj6oW1ytSt7PS2xsI8lwQXkrpqE9OsIcUPzANgYSOlH7HBlbF4
Gcmq1IbXbb/GSbP8PnElOpZeWpko2wPT3NneUIDfLr1SxESXYyRg/OdXUC2G
YbEV2RWCT1BhPOKXjVDyoG27myJVJhYHlOwXe2gcWYdBtYDQm/QVM+MjQp5l
vgZ/XTzliR03HaWOX/lmZg92lZl58WLgWkP5sdlFOiDYF/Kw8ZdNiHW1WPo6
yQzZe+yHwoizOVgbAS2OD6zxluBpxN3PF3u9W/B10V+35lwi0ll3p5AHPccn
LzGwrOxVJhyqeRWVGVDOydUe4CTXKm3vJ05ghRSc7IGzyCl/ktZM4DbedkI4
SiZCTiQhzEQmaeKHv8f+udVEnIi9aayau6f5rC1BsaOHVv1e6JgFKi5DyedP
3PsPoC2z1UjTbUpXM6uTLjFfK9GoA9tj0yQxhYkaT69DlF99CykQ5jy9K6jV
eWR/Y+qp4dGo8rnV7nURp4iM4Wp35CG2xqMOQkr3WhbxfUfxcRtttCUNf8rH
S+1mCfVWCRnnXzSnUIFZrZUhvJ/XWlqSFpaLBavkDt6NB8W73J455o2OpWWD
/9/VC7NJzKumPo9pO2U1lw3w3Zr4+fIbXTQWFd2cWSzLy48DeriVwkKIIlNq
1YslyefXzhUcUne33MRAXP5AvsM804by//sdWt9nUdBL50BJBv9negI8DkfA
Q8/VlAkpl9z4f7OepuObGy2FwzeGfR10EYLAhGAUAf+g61tM4TnH5civgcCW
Mc9VI2wlSqbMpxs4lIROgERUaSkbEz4COcd/I1O6TEMc8fcgwl86Fb2JX9/2
Juc6Wld5u1C3fvUyYqk1wf5IppOflq10u57vE/IyyrGBTZqfrAHbpvX9FuKf
tjusBwbAHK1+fi8uaUkUa+2GP1lwrqcHgN+hOOxzfU0r2L96rZcG23QmNsJE
y8dcJNX5euYqhGHB/HlBuBpYBNVcqUlijPgqzfNNKVrObgObqkBpKilXXisl
eoe1BWtXmWiynJoKi2Sqxj8XIpBp4P900xovIa50SHiohEghLmD92aKy8Cyk
5r01WWujCKwao5vaDTXQzwldtxLWUNEt01OdRD6Gqm6TfvJ20qLW7i39kWS4
6Fa0SsN0M6wDT4dtTn1M4FIq8sTVWfasPE+FTPvfm7rdaJd7Hckx1b7wyCne
sZuxuTaUQl+7c/IjBUNTOvw8epioNAhCpHEJtuxzx+M/O3L6kVNJIQLNxynd
TrDK3f1VPqGRrWlU1jKO1lbed3i6FZABvg63IP/ZI1hw+GxTwahXXsDD4+fV
8OVOowTA+ajOvBsqUlpGph4JpyyDFBv9GN5hb6k/Uvs+4Bxw4SMMNbcURWu1
pYmhfCSSpXGy82v3gWYtLZO5gm5ngLB8AynT5jbX06/GTqL6WXc5oii2MZoq
5dupYOTOCJqfH6wwznXq3Jq4+iI+Z27OoIMH7WS6r++p/KAOXnhEhdarw1cr
u1x1Qn1jdmGmzOuVVRgh7YRwLDEKUZvXqAzmPDFvlwMk2hUipmoxEwRsizhk
DI7SXdZ1fUvWqSig5niRUKluQTd3xyR1jrLvGGe7Kfq/AQZ512NE50JvwTbh
YYEky/CUmPNfDLb/SiyRUi1U44rrm0EVRB3skC9gw3rOpqrVORVViDA22LVE
jyOp2BXioG9K1tuCuLkILoR442VzRh8b7d/zZk37IhmpH5cI5YjtzskuJ/Ke
J/LRWDi/xsKyZUAx4hDo70Lh6qm/KpyDBo504J4l8tvkwkesOOZ4Uc3ANHRq
pSSAJeOeqVOFue6dxcfIOhOIgf3rhkY+U5pW9VYBbUQX+bnouI7Qu8O2CW8D
J5qSpZGfTNefCeblNpUG6+KWyQToHCFbQE9LAi0RkOgCjg+JMCwesBqZf+6H
QSXfKQnrVd6jyim8xqyWlg6Gv5FSWxPWQi6AvhptgMTZovQdIUKzzK0o4pZz
2VLTYyyNe0ggSm6fdRb4RZHdAlvTrEuIUj3ihdew219+vCW2Z37XLxcpwiap
ZqqU3zsM9ly3Ew2JGDTpmPE4YGN9UFZnWAkauyxnrT4xtUnAaoNwhw9xxZa3
KsOP9Z0WDWdxTPMKOiIyGDXdMcK+EFMhgRGakN02IvsE6cJBkT1DJPkC/GwV
RaxxE+fQ8oPpYlQ4ZHuws6xFqr8VYr4wvCnKSmBibtQtJ/DAXL7V7tSE/8Qu
mTo1CTk1Ebpsy2e+N1uhxXuz/NvVarIPtheNqhUdKTHupB+rqWw5dCdUjk4B
FgAVfq5p6ZDBOZfuoFxoJdlQymWzTezRMPHhQz9frBe0yGEfLl+NDWM6dHm1
Qk5jT38e9vgfwfQ/ZhkIGi/MnD21vcrjEOfU04D7Q47jMteoywOuiyd8YMT5
vpL73p9wonFsDeYqjH93q2W9KgMz5Iv/4xyT9TFO4/mf+EUdKH8tRvbJ82Sd
Na/6Nzx6fG+bLZRBNrfg0U3UAXExP6pGIxGdgTEkZuZn+Udd/1Pi7J7K6BiK
vVe9F5OJY8jnZvjbPZAsQlygAEWD91lQ7gYhSoMG3ob9Jr89MAdW25LBr93D
V4zpJrVAzU/M2pg7gkE7kOzBUOzpub2gVD5zKgn0uWW43rA3wESAyx+x3hl9
PdQn31b5l/A4rKcX0wCo63a/LJkPSocTBUqZA5znKP53b8NVhRTAf9pDSR2m
U7rF0h8nm+jIi+NDA95dG/mDCtdSuHCB1/FsC6SxCEqe+VWIaRvpz5PtOtB8
sv0mMoRlWNxBCwgkWTShzEXvAowYY6and6UNUc0lVD4CvQteY9W+1BvV7rHX
RPGDZfGhariEIhpoPo7wLO0Iqp75pGyz8QtwNFaqVqaO4JBX+EL4EkRYBecP
FLvBsjYPGPfcafCa/LvV491Z34j8b1CNjTxenFURYdCik5n9h6bDXdUHtfbf
bZOFhqiUfpZ923r5/WTUurEjo46Fu+KTMh9qb6dFIVgw/gITU3w2rvcu43b4
M4GhvMRBNUj9yMt8CC2I0YAKyq1YuSoUWbz5T/RYY5pRaRlufRorHNS99vOg
V2Cwigtp6u5yXgc4CglasGgrWTMyjIaZ4oBimDO/s3EqCkSef3XTSQxxA+Jm
bN87gw2YwXvSLbMA0+H9NXsKyLCag4TwnBddZWUV4ymT+E7GtGfmFn+TTLHB
Sj8T30YwLr0ao/OvzQ7pyi7YqUsvvp9mfd/rU2rpTffE+G7s60bef7s11vhj
OdokmjhH9COO7Vho2a3jOnAiqjYwMm8TpPtHnusE/VBhNGYrBjDfGGZZPuZo
ZLBwWwMXwfszRwXkCGpFwxAKd1e6Dq+yfQqqFymsR5nkAsWeX6qkPedHnung
NiRnyxzQbQYgXgYcgjT8+GgpaV7ZAVsdlaaINXssA8SOxqx1tN19M0be4u3r
TFoKT2zsSGdlse29kvmn9+eyQSJ/VvDIja0rq7PyAfCVAwOG3JECYO/jNUvI
mjUGWHHjoiLYkTwBlSz4l3dDXNETuFCGl/A6rJyEnw155SAT3UM5NuMZduL7
xS+ki5J6bNFK+lbBz5j2mXw1yMeNFzYKj70rg7qoI+9XKhwvnAkGdXBtsIsf
2AiWotY6aUu+lhwy208LsO+TPEgODBuh06AD5wwicUGp/77Ycn8NYaJiV6vE
IWi0gno4hYOXgpCW3mADcPQKoeYXnIS1A1vsqgmv3k14fMBLy0rk09BVdQJk
qjZtqHFGGMBFwSvezzaSJcoFt0NKJ/RP7garZlrOoQBfiWxqOQrGMuokqfxv
fEwZE85eG+fuW8TV2FbiFTufeT09VsWuzWrTFkH2QVHXx1KI6MIBN6ZhzAQp
hHGwYpdfQAqoufkSj+oBa7BCih5qVC4OOXsNaCyCSnXNDfipNNp7nfS7l0pr
qLKlcszK9IGFH18079ba6IIve9h9z/ZNhQlTWfrS82gCBT5xTB1gXOsng9ot
9eGLcagxRVo1RSHl0fXFWIu9rVZyqrfy27i2ArgOMa2lp1kNqEqmcE38C87U
lNGlutEcjzZsQZ1XYUIeglo1J5m8eAhzI1rvjnEidxZnvQXZyAQTZf/KDD31
Mf0msUY6byMhzuLfZbCS6TmYDWGtTaV2XUNjHs4uCg4TE3lzfvEQ/+NzAqhN
bTGlCXmamTeQpBCTf0KER2sJJErELIcbu6o9Hje79zskZpmjB31u5FneCyb9
gZmKLy2kUXHo5BW6LNPozQ1yMfvgQALx4HMUWOoDCsY2pC4+/UI8flCbljrJ
r+O7Dk2hDzx5Wtcrx0wRmmlrImU6SzkY34UV1lQdawAme0aN1UIcGRFrH2zy
vJjmQ0zrwO/FSB3Z88jVqaJDL6ZWzwNTulI8Z+4vW5goiAdtSgPUjplj3SsG
H6oyLFYyexqVq+S376mDJARuzAkx+ZtTtXo+s+GIs5ZP44sAwz1zoX1yxuXT
Xx1zCN3Pz/z0nSS4C/igFz3IuUvpjHB9FyeVlTZ2yLdVD2rjvYc7dcaxX1bO
5wElzPWRHX8fwD8lnx8US/8n46AFHYMvN4+YUsc5e1++tlaA1jdLIaWWhD6G
rhtTgXV95xvn5bFl32sHs6imtq0ngkMv5KIWi5wrpp55YKRTDlvmYrX5lfrC
hraCLuGvk8pCN6uRhgPPkhQLzkKi0xfhmT8wdVWJv3vi6uRmDmRI+NTtD1vU
xVxTdgiyIZbGhuJWN7n1SRU5VtIQJOPvXb5pqtH5GbEEEYMpGy7nrskntsHz
qhYK7t4uxWx5xQ0RCnIgpOSXKvVaK3Wb2oJ2Z7vMAXyT1Jv6DR0uqPOjEVLs
VH0ahzBT+wS6oJFByxXol9BnFUhIcPzny0T6Ct408ttj6Sl6ielnYvzJGpH3
jYuj6Jm7LC8iLmizRJaNPw7TgV9HCS0JctelgBNdrQDSRW7Ouik7+L7pVsbR
gTwuG/N9KSN/z6xuwh554EEvq6LVyAki9mRe/Qjv2iEMt2OqvtptYJygHDUw
fp7FvhWsRdzlIwGt+UwkMdVEbe90zc8lqL65izRMZ97vi3rlsbWi51CKpUu6
ZYf5EJEZs0+EOd8a9KORfrTLLe3nV9JJRDS0kq0GZ0CVRjpjVF5Tg4S61OWA
Qr7aD2tNL1PtynlvLBUE5zp/Qc9r93BBkZYLjENiW38g/jW//HrlSEjLokfO
iNMPm7KiW+q845/sq6uKAc84Ah7VynnkdxbgO2oLMBaJdlgFEdwzv7Bl0bYR
raY5B0/trmlujLFKU8UQq/E+I5cL/eIlAuyWndxZMGmqF7k4ihPAkgX2+gEp
maOreQWTawIbCFvnMb8Hv6h4ULGmnCGweAq1qFO3VK/IW46Qw2/yx9ap+lX7
aor1Vh4Qt9KgeIhWXFeM6SJWHyPkgmdqwawsK0uG2x7kUr71A/CHZz7wW02O
KyJbvh+PHRUCMWhpaFT9AJvdFbE2UDBXT8U4T/zsH/U/6k9ury4tsa3e5BhO
CoycayAZF8YHH6eddhT6TutWJpbJgxM8ziTZR1SVAaT6A9USAvCcS5X8ORxH
Q5dc+xwvbbukHubaZBV79JViwzR2xklTNffcIlgu2lG+A97oR8F7pjQajo6E
XygQQPiefiKf2Stz4t+AlbpoPVELoZI2vA8G8I7p7l97WguXYLF5JuxGplI6
lvfilODSHJ8jhoclmuF3hCQuJA4eZUdQqj6N013jACtvZDJfIbROAJWhhmEN
gTy+Qc0TgT8QeRLFq+3dILftEEySyEhE/N0w1X7chNkZNSxVI/NP5XxPwYuM
TvUhMEpbzEdIc74BnN7oYGLqa+1RWPq1begaB9iMI23UnV2y1eqHmjCGJ75k
M6JYLWnOOo2cuIT3MS2uWOgCCsiXf7+YJb9UNIikA9kfQ1tOTlON5v4z+Uod
ZXZGDu3enxDMzS6dB948jQX/df9MVGFPg18u4+Wh3iA8j0fqyvIpzcaZL4cW
oZCceFonH8BYA/su48fYEwsi3+KGb7i7zQ5lceNNx0CYi/qZ/7sWxaxwJVbT
a4pPgmrxVJPEZquXtkzXf2420ke51pWsBechPU5kuS7ICB0ijuu4kHgcZHV0
zsLJp+oxNxElFvstgC8q3ethBreZcC+4pCUA5dO8tcppmDB8ex6Pl4BWBNPg
LyU0kMEcWQ18MkUHCM+aZ/DI25AVCpzV7R2eX9FQSpiWwuWMxMDQz/PNQNL6
ZJnyNg9y3XycDUgK0bYZ5kLl860SMtZYfkf3pMdARw7eG1xF2wsrf4WfMA62
ptghih/sO0BfnN6O6D7oou7qCTmsSWq6E/RuN/N/A1NHF/xdLqsSpjwHgCXX
5hyL2VQOBxclTKn5RyPtCodbwRwCkgsYQg6OSllclFm0ODwHjlIxHvh2cBxG
eMfK+bS0WkA8RfQAtIYvvGZY4ll3ZGlVDg2r+IN8ecco2/8yzr7DSouF8zFh
nZ4OLCxTQcy51EvfyQDCJe4Xko5Md4AfrfvwY7Rqz6spWst75BiVxXbc0FgG
mmbXWgrZJ8b3bTW6HYl1Vu3b0viI3M5g3vO/VyAGdIAjEIndQmW+KaB4PVkK
NhubJjtK7LMoNjphAYaFyNfxY3YnOKWsi6gkbE+aiIFKpbU2pKXQsOHY2QrN
pq7CB/2ES8TvM7WY0CsjXlPAEZy8PudBKtiUva4vFOYQLofM96d0N1vVxedD
FtWd/UvY2xt0NGQBqvxjdP5AjW9LsAZJDn+ldujdUtH96Gx3aihdgd83NnYx
r7B5LQ9n4ijTQAwrLVqoZANENtOzvHwhuBXzl9JiMcUcxhArmUBpmGqLac4J
rTSMMKbWB3Oxp3aW0j2my61A1yf8qiHirrtpqxOFU5aDvXvxhcJVw1bPAt/S
HY9ZRDIRPQleBPQqzjzjUft4VrCShuYdY7AnZn9Nkv+E3oL9aDc4OBCbDVSt
B8Chd4/NUCvonw7vCBUStTKUeEoOU7/PRBSvYnDhDE3MZF4ve0KFaD8gdHwH
RDQpgdyHnIpngXD8VyP+g6NMFtOEQHY41z3CI8z9CJkAjHcr6sBZZ5FOPu2x
M2Aozmnvv2t/CDcsTAfHTvEDWvuCPnAp9TlWpoMJWQYHWfKWVInvixE1XcKQ
K3Im/iLe++2bYj8Ph6oO5+jrbS8SGayvaeSEIrlfn3R97eUtmk7XMrW5WRgp
v/wFnkn0Un/PlXUaE5fBdk237Q3bYbh75sQnULRDtpgXhbS4pNc7ZsJanP7V
NTMEl6q/r63YmjKl3NDBGydv7OZowSfhtplZbjtX4K/5kClqqCNt5cM21dQN
saMRF3klvpremg9h/0l5Ifd7GTWRd6pYs9ABBd1tqn4zyPjVrR5VWtuqR2WL
L+AXgygkqLTqgTPUNoC70l5YMNgR2ZAJHLwL9InTPmgCOJR5XSa2ipnZ0g27
WUcTMbLb2cM1F+n4XFIhNWXbeHaZ8QfmbmKiw4mIxlIcu7jc6y/uRU0nDABM
0clxAvuuN/3BWbbUYNzoJAPM+RUDoOPNHONZX4CAUeCxzKwDcDFOGqhMbeXd
F1tw1QwDpT68W+W23agPhdGBkFvWNQngHpCZVFLkN++33CFbAs4f/ytYE+zX
ynx2EZofYtceKTg+adXiULf9q0HKoOClv+mu2dvQS0zhdht2Y/nMF+VQ0pe+
gAMhHQB0UT5w8QpqGDdsvpeavDW0DBPqf4sqjYB32QW3ZWBM0xTz0wsALMsg
kVVc2dpSHi7UkzV9Tr7MBrU+uI7IddgBmK+h1aB3r2FQ6uYNzrWzduVZ1GKh
0XyBry8epU2IMpLbymd/GtJBEJhVGoEV6fq2VOgBvKbA2e+xHf7Psk+gD8DF
+C0zr7F60+hfT+NEBEMmo0GnJ2eIIxyraNhxyRx0rQRsiB35Om9c8Q4eF146
O1NH6x4srKLJ4l4f3ipYg6PebrwLR+dSfHy8CdIXotEljaVnqz3PQQjzYg4O
41N++7733J/5ZjZJ578ykw2uxsIrZTSRhC4txwdNS46n4rIIspXhGjXKMYL+
fS1FMIzIck0jyAtNEhM4BdD20rHrqCZ5x/g/bXhx3Nz7FML6m8tn/SGd8oeQ
nKhT+2MkKAXA1QP8A1YwWCnCMeGTRHf+EbsuKRwx6/EC+inrg3/B0Mjzr4Cd
3DYK8Fr1FXzMkpyzSh2xAN157zKxFvqnGtHvkA9lLWoHrmhcrHLdPF/HfWay
RygvGVkAwkkCzf9WylulSL29H1wcTmZIlo+DdUNMvZJgGVkhNyUj9HoM2iTv
PFR8fnXZ/lKBxuIsOtpQl4X0fLETTP6YJYj/HUSj/BC+w20aDRFJE4u366jb
eDkZ9U6351F12XWvPPiSFBK3dGCsLM/09//x96We/M+6JWTVIAN5U7d1153w
sxnt0mNk2I7N1R91erjYKOke2N/PYZf7Xl6RtVYcc3e/SO6RDQTAUf+Qqoef
oWs/e3I8IDXO8E6hPXZdJ1CwjWsLDavh8MqqvHh2yuneVPETkITiuzA3OZ4d
7ukk7iRPuke7cyAzAhA513ZsSrxuJZwF0AyFXiTqf+3sNuEuCS+iqOtIwi0m
DPrkYQ3xwQpkuZXD4SUoOdpfxKTp6TKIU7YdcAz1TOX4rQuYQupT5FPBfwI9
T8ySvP31HFTOcwLdaY+fxwZZ7RhNdk344zVDdkrcakQ8cH3DOAdx9LEv29X/
DjdqSxVnhvG8YoLptsaZBj2Aukmp4TtbcZFtjHD2fCdwpjUE1jMg00/616W2
O3AjCs73d3m7HnhWefSDW/Gv2f2BVe5NElgiNLjcFxDWxw+ZOCF0a8TUvB8X
m6fW7UEBtHKfOioU4cLiGvnRwpK2vJ9lDp2iOjs4cKH+xFEkvwaLiIGBD/YJ
p+Dw3OIprDSV8ZChgXckRpOl1UO/iFPSEEEUXvdmmGqfsl1kbuBcDIzt+zuM
fCe2/7D2LfcuDvWISuV0E5OPl/uOPsqY7E15fAB8b+Sf2iLINwcWeie95K9q
eubL1xe+ql8HE059lrAVR4GI6TiEJEhqlJD7Un5xg34yYvek+Ia4yA2iLm3a
m4KLg5eJfK0H0FC8lhUJnjyCZMefhoORRWg0QBXjau0lXT9XLsr+L3uM3eZn
z14Kz7YG+0oU0AKpUJbKPg8g4RH4ILj7IpukLubJ0BqROhazRpdIxKffNNe0
2prZJjDyAcmKg6jhR5kgk3LlgZLS9xogZQYo+c4KhM31fZNQiyd9t87yqOkn
4Tu/xCVyDcGIy75TApq5a1mzLF3a2xek8+GMqOWs1dnqVQfx7qVz8cxGU6mR
ugmq5Hhq9KoArGIgDjfA2Or76M+yerSecI5Z8c6Z+GytQ3ySTZr/Wjr7i1ko
Ppj3di6XvLCZmcTLfeUMhPIZNd1Jny6IqOVv0oDWY4FboB9ofwtDGjk/vgbZ
+gWVATuSCxqc3LXlqzY1joHkqqSZKMACgQfgy2T9wt/a9PmQfJYK3l6uGUSF
G6BiNloM4sngSTW7WlQi1AT6+KwDCrVNYw3ky2nkbQaPwlZcd69XXKVQ94Gi
xJgnrhl/+dcnEfAcl6TfdFijXy9FmgwKxgMhK8HHX3ZCeMbvwj+0hvcYhN8/
pg+BCIewgkpEHvlGPixj0FsZnh1vYG76Pdbrl+CV1AflQvwkyLxNOQT0VnIR
UenH5Yy94QWPoxbT3EKcZphfHcAiF7JwUcC7shms/RuZv1Syko2VXdCkTiek
kiEWK+l7gMe8SAEbFCUTCOxom4fdstCkhMxCcy+yOhM04PRQbgIrbecjB302
d5B4716+LRM0Xgtyly9hDv8MDLlRdNoc3MTFXHxGJwnrO5lBgxUFsOQnnH7/
EEbjtAYXOjMigshE0FfJbA5R2uRZ4Y8RWYSvpUBEXD0tvp5+73oJlBkGvFK8
Cb35Eol4OVKCQvhUgbbWPf3X0Ifz3yqPqtsxMYTr7nX3KbYldaMc1E06gk+w
TgifJEfbz20jNnIv3ckQ38XMA7+pgBAuYGPbMk+JVfNWYGwoD0va7H4PxaN1
0dFyNds5Tvmfdho7cET2Kczs738NkE8bNj51BO7aM9EngqXmMbccWm3F5ln0
vUFjNfJYQCM7jxgKk77Z1/gOxgYws3M2018rZMUX7RNWnDqQ24SeOseDmHX3
n9lKLyMkIbflK/Fm9s1WairxZBuECra0zP2rVv8ZJD/KcqK6tXKZXLQRx8nE
HTthlwFU9LPGqoCu/MdpSr+9HA9uhqed2X3O2pQFTaWSwNA2mfPjZOm+i41v
/e86NJwGPe+PbgNOBlYVmaz/bvOEG3bDxPpOxpJIC6r9GqJFYzygMevFvzi0
OKLiul6t4wF3/uu+Dy2eP7/d3AEDnbX4Usm5oYEK8P+qXvtwauAcKWOkudQy
1meMIgoZX7whhZBGrieSh98ZnmtPOK95LI4wHF6mIfis/ZPuzEu43C0UFK7Y
4NN+CZU1PXr22EGyhIb/vZiaGwt6wv7piwLcGeKLTCdBuZxqm9kaeTnSoLDr
woUlYCIlN/cXbU5KuIUGNKkswsKc6+RJuhuVM+G8UUrItrReLvmki2vDPChj
W2f1c2m8TSqlM3VoP9ltBZ98oPb4+Gwt0wboJOB3hJB0fubP0neyNk2XdN6Q
kIMytBmji58gfYwzT8+WLAc7tg1JSrifM/9jE9LXVseH0rE6rb9LRzsSATCQ
Rq1id6QyI70nBfo/4Yt/mgwrHnO5R29mkXhH1AHVts4rFbmAOf1g6p3WWAAA
1D2ZRYXqIxjTfB7xP9vggCq4s44qNEBLs4CiwGWENKtCsJmtaDb2XdmE7UCh
12UToqG2f65Sv5g5Ypv22YC0GNsCCcwY8tTNZQOuf1xZDjxSPzL3oNicJHoB
1AJaMrcLZLvnINfITy0ZaXft96Qmzxrzo9pk99+11Ygg1WbgC7CxO9FC/tQx
c2hcW0Lao4y+l3tXGuNP9aBvUA0WiKCjQ0iXIQk5H8Hc5+IoUM1bobpjbS8H
Iyl8DZLuLsOcid2WPR8Pe+BBHYPZNJX3BgXIpY1DzPM+Z6YWdQ2z+gajwLME
unFAIpxGyb1cyFP86slshgue/Dx+gM/6oIm5cF3HQSbSZ5grhY7QVwKs6IHt
R49j1zpSR8udiHIy2rhZhkirEsYc3ZbMI6WM5rK3M+iO5B7WrQM48kVfucq8
71Xss+eXTA0NyfSehAR9UHtQw6VDiGUx+TThkvZhwZ+BLilFhkfkeQaEmQK4
D01beDqJwOvWrU9at+JV9B4RthfFbmwo5orbjUDjKsRE7ZmrSrZvd6883xnL
h3fG03qU/9Kt6exyc/rPTVBqo+TJWWXN+h237pdp1J6th+LxpVFx8GLX0T82
ROVDMvSC6PL5ZjopKlkQMTqYGlGIGVGX40iw13jEwG90r7+fq26wTQhX9fyK
t7eJU6QcDw0DjgofMk1190IRyVxo19nIzuN4SzamuYlmHuEmK39nJan3nFTU
1dvkWKUbpKPIj1+wBKbAAX4bVaGHuI91zOk97r04nfaGPgktXHvhN4RBn/iD
jxlrqlWcyHEqiFtzD1OGt20ag0fM/oCMjMv+jKos+70rvXCL9846jlGKhE2D
LQUrnSIMXdzzr9fMKcxdS2qzT2UNokmHug968z6peZ9SQbc+v1yW+Z2m4G0g
VjgwlmNmzeL/vnVG3Ug1EpSqlZx0XywPKx1J/UCM+8ZbKW+0QClG8/8kTyno
xaI53kcGXIQUFSNiJZtBuM8MfwhaWTmcrXL+4fcDfjrKkCqvc/AxJllSpI1C
lRRpZgFM8S7PXtFv/5X50gcyUNvQbWAaXFAgMg3NhWVLA+Ea64KGIAzGFOXS
sIhns8kCwPIdxK8qsJC/yRxwFsgJbUDRv2Ep1mntktDUOiEwpMD00iqh54l8
wfvZRXC9etE5yBT4PqjH1eBNWnwi7Y2AeR9KPw5ebfjTL7kREFWN/TYMLV1d
hNhvqeHu4T5fc3o0D9IxvjUfhXWunn8zu4Yh1dYXOj4Z/DjloulPXpPbsTmf
lWN+wck7KVMUAwLfYtXFCzwT4ZNf7sCOc8yabUWFoMf35oHRvriTxJax5Gih
ifkQDQh3Q1ydvjRYEWTJKC3hZINCn8RavwSF11jlJ/CqX3wMy63bGFnrQ8fw
M6N3UrJKj+r6CmsFxftCv6zbudU1Vsj48tsXzrPQNwr+tAA0lkvIrAVH/3/+
xN8su9nzPzyTlikqd8fUppK8I5u4QKDQ1XKX4WNNlJcJUQDbXWyF8ESGXoJ5
mHCQa8W6zTG8XWV7QCqy89NmdrUsDVGtMJO6rdmP7pCQSlTTjNePltGcblSe
AxCb/6LLfBfJq6dTzg6TgoQYke0p8uFH6EWo2+ZeRzGaK2pPdP+sQF9jk1w9
0yNv9ciT4gC4EOX1RQ4V/seDK2/HhQ5iae5U2TOWd2MxCWjlUHTrikx5LeN4
lFI3CkcCT2+m7NaBJ2a9NECIeB+b0TOYz/wF+xmkTZ4RA2cAr/7PtyhhauE4
oZ1PmzQrW0m0NkBl5iVWgUrbSpP4J+WTVTgKKzKTsMi1ih8h9jYdWrzuDwRB
tZNQwpJf6w+IlHgwUHWDFtOusmSBXSPPfijwYviwbT6fTDcVHbQXnSqlwH/d
AWGPCz+fUaNQY4UMl0CqacQowim1OH5204owUKciGFm3Wu19x46gFtIunmst
fHH81cH38xhk8F0uEEKccJ2XD/MX18fT2D6t9j67cIl3MCjRMcaqAAYVYuB7
DZG6tizFCeNsZlXQm8wcGzK+55Ot/Td5ex1IVy5Td6j4brDikPzVUxto3dBr
NyYV1jWLiJmfpNqfA4nGI+pxnKCCscoHK8TJreXD9XJyyoPXOdBk4wu4CAvL
fyR/nlA9WLyvI4om0Y2+IvtxuZAOVn0PCMFwQ+KzaLPgrtwTzg94h7eTOtrG
JLvFql4QDQifT8NKAQqsIrxbzDcP+xSxf+eYXSjXEdiHw7ueQk/15/chdFyy
XduqzsTA/VGWUFLQYPuOUucQdLxT8zJqhqvF1u+wKSMEvGAgIXMV3Z4gcqRW
uDiPgcuDCAz2FZEXzJI5411riUEnNqPd7bmsci1Ps5LPSn+9QVJTFI9zph4f
5tUgydh1H8lcJ+WHjHyZDCSe36rqGt6guNs9Vk91frM+eJaMjGiSP1iW/96F
o7t9m7E+nr6bCIViAPRgKduVUzQ5FcF2BueKrek+a7hywerwOK0x5T3bG9rl
h3VcoXXrDLxBudQSi4Iks7nZ8soiR71jIq9DboCSPVaS/aln78cyuK8s5hp8
BinddNIzWzR/LZ21jbL/ihlq9GSEleIVMNGMN9xTZd8G2jV9s+J8FwjLVk7p
oOOJW6PsWZKSAgn1WADqPYxB0IUXCYje7gHSVROKgo4h/Myc8DhQQqh6uCMC
TxG9PpvoCE1vg2qfwcAjxtK9waUU+nHOTYiwin69VAVpES/lk+CU1H0OHZnU
FA6npr3+pd9kTrZuCmsG1ZcjumGBHEa/lHxHAEd0AaFB/XbL5inZtyzMUR7/
1PDT5LYgcLekslsTpqd+iwVHAoVsoJ+rh0vNd9ceZ1yRZIdaOE6ewv5WU4tU
JUXg3fzrfIqNdjLNuKPLchHisa2IHqj0aWrBigToB3r6YM60zZxIBQUEtztf
DfgPxaNJc+T2N0eXpRUghPPD0Gx4+2wKTnckrxEBUZXefVy624zuhuU5PFU1
JodZos/wsoRqB4XlhYbQ7Rjx7/Qy0D4cq9g2kPHyhAKuqyrR/qZwk/dsrO/I
kx0nDEsSWg88zBG1myKkjjKuto5xQuxskxEK8L/4nxsn4ab+dqWLOUKVOHiA
kby4GD097v2pEXgMOAxhn/PbJ9FXdKs7vZmwiQJ5cenjATuWeXcZovZkkRhn
Hzs/ffk3XM/FrHWlFke6FRE0roVvE5/yChGx4HG68oneI5w7akwmBf3e1vCi
XZmfn91aSY/l9UArqKQDUXdoD826gjFJGGHUSp9GCPGXtkMLnRdsL0exfMJI
uXTYsn7Puvsbhe7s76QYLRdB+m1jQixv0sCnnMnMEP6ohJDA47Ebs8mKoXGp
oj5TFyAawgkxGFoKcYvSlOb8z6Mnc58qGXB3F1Vv/TxAzYYIMHKPnj6I9wo/
cCN7UFpVhxkRuzR1B70b39HFy77q0c41a2JucfvHOdfOOtV/lCQ8JEwuWFiq
7a1KeQ0fNNyYEOyiPJ8nTZYlNKNp/4RPqhYLaumeQWfW3u0Ofp2jOaTvzDQE
2AwHdF+fLVuJopH03PFH1HKgBcxOBewxUteTwQRHPjPOyIx9xyn0s1mjbmvz
2bqh8m40D4VNVBmVwWcDCMjpZFp2C117AiFiJCb3Y+dvS25XZ19XLh8bqWXN
mouxMAGuQaTpI9mnAfmIqi4OV2YW26MHFtsfg/p3O9+PrRtyDLNxCXufd8xZ
uARDpw0KP/d4Sa2sLvAGQMtpPB6p+XqfmBZurzX4CqRYp54lZkdTqA1rCWtQ
4DVHpLh+EXjV8DWAjvjadyDf2MHflOeBoKZ8H6/flm/kW0vKInynw4mn9ZjK
6teUFwU1/moOGobCNu05gsnuoFSU7WjDfbyJ7k2nXC9nqn5UyJBqLnOS7tOB
qI9WYRsGGYYhBdSi5WhTtRSS9+2xbhrcVZ4AJscLzj+hRDtUdvgo/aYs5WJH
ziWxI8JkPui1h/clyteYPiFHUzL6KiOkoR87YgukxSKy35qmUsOSc3aEDuk7
zGckW2hrh8fPOjh7MrqNxbfGcVv29ajFNR4MQTT/hladallz9vQck5cWp8Px
1YcDOkdFb2ghFstWWlUMYVu5luz2CYL91Ml0nuFwqBqBSHrcaiKgmtf0Mepc
hYwuLJjgSRhPZSmAAxvINRUZNinBdI44MZZ4AQ08G7sG9GBfQASZ1qVJuWdq
a0AdIDKAeGokqsJ+Y1u15UCVXUKUGHA8WTibZ+C/yBDIq2jTOQFvLsRV5vQW
NjsTf7MxHJIaERzZxX6K5WL1vibcWPzPe26CyzuQeFRYWPTk4mhV6f+IoF+X
VDv+tHMZaqXQigRKecaj6kD1gi9x9BD2AC0Zia+bMiJs2/tQq322svJIuwnk
J+u/4p/5tfQe/gHK2k+jAHrPDTGcoBIdHCuuC9zXHbwz1Sc4+s36YBQIKBDP
q2MayiO11YLCsOOaz+3aPSdYqBKNNIoiM6t76CYZrzN2jw0asLvsdQjDbSN4
Kmyebb/oSTHKcVB87qCrrTUW0Ky/9iA35mD+Ifm10tpQPxRssAp7pJcKnvZ+
BCAE1jTzGbiDsk3hLk0x5RbV1F6P7ohkUdgjH53W/XaOy3xgNNWXbLU43iPB
TAJw1VTFshwPcggmY2eAfRkTLfBHGodjlqQ27Oop7/SSTRmHfuj4/Q3dvZhw
OraiGN1RE37mCPzI2fZm7qNt61BzrYEpLwZWBIheGswy1kbyAyirE4nkteL1
Da7z2MDIsO50y3z+M/hoRVyC6cD+fRli/vuLk7fXw/xEX8/V5WRT/FdyLWAk
ZJOxAnrizKKwZ7row98wRrBk7frQ3d+bQQGoldl3B6dR46jngEEaJrGUvgcR
iiLOkkd15RPRDnxqPeqnJhBPL88vwDi83CGC07gT7FE+rgXvN2g75doV3SaZ
a7b9QXAEFGiO9IuTaSZ/a8xTwOuCUGIDLMgBOZZlLe1GGC/7FqEqAFX5aHkO
tK3sABJnoNEbuwKFMrFV7syG6lkXOqYv0erNPJk4XgTtgJQzaLP1Dvfxw8DJ
sGfK6f8R2eZC3BUH+PE3Ay9enqcXtF3CHVhitzaPki/muX2UuOJAKHO6Eij3
hMac0/IQx46bpM3ck91+l8koIyi1+IXi/PNNj/pSoFPSAJAnz2TxfAbhTPbY
ntCIMlPo0supuaovio4aPRewTS3GDo5wGMC1BV5vu3OYE1HVAtUALCpR4Nzd
HzBGEfYr+sB9/MTv6XeyP/BA1aFp5EE5UDpxfutrpXt4C5tvSGz4X1Xse9qn
zI9Wcg8Vkgywwm7LiqNDm/OTfpi/+unaQ67HVHM1yZiv4IIyV+TGpad+KUsE
D3ymQ/+GvaDpQTaesKZ0eLD7p67z3tm1grk8BMx+tEuH+76hI/1fHunVct4T
rRAvF/yba6ADx6Sz75JLaMZO0rAkc5qc6+QOvCajM1EpSJpid/BBNtcbliR7
BgcpGHuHbym1XmQyRihW5+C4LoPwhl5LVB8VyqARuMtxLV/agqKrZLHNAl+u
9MhJEqc/PLzJeTbbATH/Bsfhjz21IBevxeTb4ca8reKfXHR8kCrskCLDbrHv
eQy/8TsLMl1jpm4zPigFfS3MfzYZXPQaXcadfHtroJFyHAXGeV2wveRkeg84
lXZYtgH+QdTDCe4uJ0CAds4nN5wZfCNX7lsXwsRTVUQnakNMOy+0quxNX4hz
6D5cW4gQ2HVSEk2MH/uwwsAEi1zguZnJQkbayz/NraieT9fnqnQzDnmTsOIh
MMRd+6nbuGTTRZCPpE1AVVVbdlQT023yGi8AA0mTBea3NHMrLtjYgPUjLsYE
mGlDxOUF9GNIVpSWEx3eeDPYZDVVUnvPyeRwM7zrKeoiYaHqb6r/X7qL1TPb
8uSe8dWYDtM1GWXGBwsR70saomKh9W/5OzNK8ZFO4AA7K2QRlpMzaxzOgAmx
9y57RCNaB1dNMs9NwHmj2tuTipnV7Mv/kboJir6Uyg6KhArukzYvIYOxASmM
qJVoL8y/CIGbzRbl0ZraTOySTP7+VtKlpr6aofcSTpIGrqLqMjtffsEpCoQI
hf+kWGVEP57Umt+gm0E82pU3i0eFpOoRXGerXxP5z0fprKQW9ZmPOOOp/vQW
h6qeHu8DcoEzLmhFGMbZudO9cWtetHA+Pa0N1ZJ2g/sl8o7c/Sp9sycSeiav
lnuRUi4+XTTHuYwuaV4LW+z9ZUGbJWCukxi/5UyuVNugATtS7zaMgv9k8fcp
JP73ZF6W2ZVbkI8VrF8dUeBlqBfiVmMmt9p4wrDvy2Pikg05UKOZ3l2pyts8
Qz4MMITRtiQPNcBbRiFLGsrv5rQCSnNvbqDmxG9nYC+BxNDITB4DcATEUgOm
aFgHombZkzfNq2kuXsUPuEAvWPkpHOZCywCszUJTtLlzQLTY46o0MUjlZhMh
qZUDuHm1yja8N7mXVIs+fZQeBOrkYdzL+Qfv9cQVf59uzBiwXuBPxEoEc70n
dnoEd06xwKzJJV7krOFErJeN5tXnZ+3JTPadRFs6+NeKCcVTpFVpDLgedc/b
2ouDAQ97jDOtn3nX5/a4CpqQqThvX6jSrYTb0wE9zbX+7bZ2vRM90p+QBB52
5nkOjD9kSZ0gw1+t/2KaCzbjW/LNrLY4mVF1fPwjeCieorNARrVL6F2J4QWb
je2Tm/QgcON3Br5y5ia6cHMdVcR777DD1X4JluEzYUwRuHmNRj6R/zaL4yXM
uVU0cFgvHgOfNSLBiCnlAAJUqGF/V3DfdWq4ALeaoNVIWO2DcmstgAsvMK3F
0uNonP8m8Nvf5sVg87Yd9uJM9+si/wZMWBHNmg8QLGTsIQOA4ejZWgB+fHEG
6p64zsWq7EEqRVmsp7pNrlrHf5aZdtnlwnXWw1Ri3oZSHGPNgn4VZdDCUF6S
9F3Li5T9wv2QXzRTRbSz4i/4R+ertwzBbsrXecFyOjF0G5oT0x3ly09n3vIN
aXwa4gJ8fPGGjfIldItkAO7o+HRkVy8Ldok9qclc0xP7ZyDRHH89qH2Wly4x
S+hrvRclohsPgU8Q5AWvqpgLOds+EwwMjL5fEgN+InkeGXATCTjyyC1NJKQB
NOVLmDTufeq1UTMUJ/Q/zwvG8zlX5mAl70HfK87bKKSop8LqlX+9/W1iPVW2
0DRzQCxOIRZZQWXYm0ZxGtLfHK+cH/Zy3rRzQOsC2tBfnZe14be5nj6WXOGJ
o4qTmk+78vvLzkj50hnTSzlzu3jXgs4Q4pvx2FT3yLbFrdgSO28ZlvVMbW+g
guYb3nCFw6NZVnlFFqaHjTT2nqYTOBKKxalwkY7G0fgOznZ1vlVq/YUevawq
wqGNvzocYVtnq2c5ftsQvkuh5awSEepyyUskSI8YXtUhq9ohYOirydlWHmod
IwIo/CGVYK/5dEa3NsFVwb6bIyIYgOjApEprUyETQ4QzQO1AoT+s9ClaDOEH
RmKaeRy319p4aC4lHnltbthYj9W3G0y8/8dRLSVWycl4eRf8Z+5XiKT6cK3M
yptSZUu3fMG8+OgXGg09ze8PrPykBVsIDnbJMyvo/jDLPL78xe1DELFQ+H7u
KbneOQY4LAwH6pYyS7hHKPcvOkiunrJYSqJBK8px1yQoTZwXWWkmBMnexdhJ
XfGoABHrOhrxzpzeAU/96M6uqfWAfRNTTrDtJfcdAm9sTl8O+H4uUKmuyoEN
oONyIWARdMZUcXPdNEMVvF34W86IfM0X3raocRT6FaC62b5a6BHW3NYcfNeI
Zcb+EJ80SFD5zYA7aJ0AB0sn4/AvViery6qEJBLfqXjykeIW9eRrwng2Cr5p
7D106sxuw276vnPIZDR0zOK8BrUMGTHEgLssyVLvM3ZrPU614K4Vk22W68FI
+bb7SNDuXssKiw7b5NdYnvdR9RpYtlo7oJgrERlpSSMtGq2lR5i18jx6Q542
XpbZiLHeL1faev9JISWRG9aiYMjJIOcGBJv6pv1TBS0FPqSi7UUUBP/pLs2T
6mmZUE5zFfNBq9il2nVQjrUxzYuocWFqSWulaeMHiFByW7tE2wGPX4JIGiAT
VOCf2BfMzh+C58WrRfHHCnwqRVWDvWDyJhZmTip76KKxeIrX0y3XsC9eiHno
kufnaBTGExn1MVAPs4e9J+g3rNT1s2LQBT2jXc8bVkLzR4lajWiNG1Jlx2xn
O5AbUiA3EPprt3wGXKr9n4QPZXQNFfN+nFPqJJMmwsrqKWhVs/RznzqwticS
EJuwPnhtwgfSZiNcNMGN4LAGrmsFOyo1ICL0MxlFSjsGFOxbOJgNnyv+vta9
GxK1EbtqOpUr8kHuKj3D3jPKH8V1olsazUmPari74HRa0z5hlHWAUedz5e2g
BJWd9dULp8giSBHJWY7BCpfhTIUaGOFH0VadH5MenmkbnEAHffVGu7AnZaUB
SF1eJfVdcJKMIcNvvBgSGWK1UEs2FdGdFcQTZkj5V1VuS7eWyqji4eXmV88q
j2eiDxMqdUZv347hGGtCX8bz+SV1oCRYPp6pklw/dQhrFjdQYKA07zlIFF7t
N+6Gw5y+6Ybw6v3WXP3RieCfJzmOj3wuZAx2QbVZjUPXbAQPC+6MWZWiKhzA
eJgJudSeCCwzj+ILEehbz6bCV53ApqTlEg59xVE6CJzEYvXOmo/ov1ZpVNxg
OPkhw+tqwWLMxolX88C98/vTp62mNOKD5aabPqtWNy//bbzj7tjkSFnh6D4A
KKJeXFkWoEHzmnOAR9enDgh6/XrlTy0lE+yKwinHLoiRocccbkNhhJUDIy+2
w3dRtooMeI6Y3azK7MtsOHtxk1COpmOZ0s3sH0rzPRQ8Wrcdo73U+qWq7gS/
w9kknD2tDqRYI4QxlrneNw0ld08FQEl2LfR1oDuHAMqWjoiU/RRfER0Or7ND
xqp8gtlC7/gsymr4jA9IEjBI1qBM8fCgQfHp69OMDnDoqyQJnxmf4fTsGo/6
p0sYbHjm/3R7kZSbI6ZR+Tf+mHHSz1REGWPYLrgMPX5H29Vt4d67YSKoz0Cc
xbkxwrXnTT/zmR1TvgAVy4VvegP7AVPHsNiW6uzcWbQ3ZRzHejw3mGs0cHYi
E51Ts2zLmV1rVLoCm0vz1B2c63Kmt/gZSIxaijzkQAEf9xJiG+5VhcfeLf5n
dh2ph4NT68GyDa99SXIBY3th9RlstZljQTy12Wuu8wNlvhGGVmyO+9RnbsrS
dkKI3qeOsuH3QBsjDLnf0XENSKbOhzfXu1uRCtK8saip31Zhxgb8OKN5nG7U
Xs/K8eemgP1wYU3IhMY+HBMLP2cjQga+Cnf0qfRquIoa1sWoENY5p5HqIT21
aXIpe/8AGYGAPpaK08d+UdRF2i9PeydZMQ1dPhjqzKeGC+Ku65bqGjRkasTp
FKs9lhxkcspNAs5tG5hg5AVuOjnArTyQatliVldI+SqONbbGSlUsatIqPaH4
fF9ztCi9C3SgLWZVtgjWnbGLs2R/ugsdHi9RIZlQ055kggyN0BWWXWa//SSB
o0n3Q7l4GcfWt3BDo0oL575/nQ8E9+idFMOpauuq2+OUuuBjc0caMTLnrFyD
ch5k3sSDm82kOWbzN96JBG7D3ZqmJOmTp/OKCHTLwaJCQwlgnOHQ3wsCIbgf
BBRXk1QfdjGPfJrJaenJ1kn85Z2jn4Lwi72Ilwwg/UrlTA1XfGvCKYBYAsJJ
WCbLr1vA+NMiaT3xP/31o1HfRS1yDG8Q5p3iaw/67UM/lRIPd+eiBOMMfptx
xFG55b7AFJXSuFLZACPyEuKk5SjaqfRmmqYH/z1LB2EUbbVZaWeiQLTNmdaA
JfJU49X3mZK9zm9zXQBnbUZxQPj5toNlO8Bpc44vjFjJ6E6QFq+7ZykTGakJ
Cnn4A4NNXW/K5LWmgVIe1KcyvFy8CtbvHV6fPzycHQ+qZZl54vz91aSutDyC
CkEm9bBrA2eakLFQj6MMH6EZipvrmTSR2kdU0hf63jF2o115xA3D6nHck+os
nI06138oVtcwxqpOv/tHesylMWOTIKEhZn7tFimrJn1Urge9GODhcIDH3n+r
kaKPUeJRcJx7LOZlfgQkSPFPu6hquayBvDqZrt/AM1+S4Tpdd+0FIU/D/pgd
uJM8Q1Ma1QejCKnyr9nzKrtHlRWZSRkZSu03LosIUxWlW8c90XwVnwI8jkJ9
qgAVk+DBza6IPWi5zYZsWQ0l3HeGy7L+xhak3y/dtgg0ZUpZpm8d2XpIId6T
79mzDtaHywu+SKs4vmGOLqGAa8v5F8QlplgFYZdU+mb3CAPCfSwQTN+tFF9O
EhGuH8OE4b3ArrUp+rAYHFOTcMa1a2hkqEJe6yy3LiroO218y88UdFF3zLCA
Ot3D5tfwtm8MuZJUgcG0UxK1G7kRGk8csEfaQBmDdJigbvmPW8zPVmaXxsqK
zpN5QOO4C1Bk3CHf9Ytv+JBuocVp23hCrIxXeweR4iEA9/4rdjcRYbHty38d
ex0zFfsquK0yBWyCxX3SFdkqdjV5biISWULQFlZ7JGOrVBUwcDbOou5BBIjk
HDgMYOtmLZJ+obhIz6Yr2tL9vTd618Kl4/GKKUR7OEIBiIb2440yMikTWwsb
lyVGzJMSFZpos6o6hJZdtaJxHvsZUDADiY72U2iTMrqqzzITKXl93hPHB0Sv
Jelok8XyoJDGFW/sjg+7DrqV6ouIt6xyDRGwfqutGz645T5/1KIJiGYrr1g9
vwgXjNYdzR2wgO1sPkoyo2QdCQOfd8Z7lvMPmnCtwNN4q2WkuL0jTU4cijbb
IgrDBk9PJxiol11atKU58ayt+iU4wdf6kj6awyjWNhBMtDfYvYQqSiSVy7zj
77wY/bF/IzbqM+l5CHJceRpWKE6pqF+7T8AFNnGrj61BtrL3BL/e/h/Cc3UH
69LRVRdch+vvHUiw+2GY2XTkDvFcV/LntrOfN3r544H/mCe4ArN7RvcT+NhW
W7T0B1e7XqC9Q3vnpqAG3yXI2TM3xc0tnopDlLUOO20LYIQVFmaAy3rFrycd
tCTyxikRg/A8e4J+7lMBNPWyPoGu+Qz566CC1y/5lw85QW+0lXWc9LB/QJ5Y
XMyY2q2VZO8LOgsPDjKr4RmCpxVbq+5c+fwjcpKOwIadJiX8mRi0TT7jUCOs
MQCIRmJmXKRvif6cLKRTdr5SrKPegmvG9cKkrvYTfOoucpEt2QxPnwKQcY+6
VWEBD1ag1eO90nQp5eeT6Zwud3Z0BWnJhZ6+Wp0OgUM9/6WAe+4bX3RYr6fz
KenV1zCTV3LPAkCmdC7dfHuNfU49S4rUv/XBxvGbKFK16GwVftKT71CRFdo+
ijgAMKEmg1lzCjTgKjQ2TJ2uMCHQYEIsXIxyjZqPASb+bifEJDyEyprFx7C5
DJI7LHVtj/3WDeSADaih8OK8bXn9iYZAEHci3D9s4XZ+OgJziOr0iKlUxt1U
DrznVnvaDZ1PqTxscPIY2JnsnxbptMY9vxLmOygd8kaMX6VA1ti/ndFFx2gm
Shzw3OvA10dZHByah1iz5tx10sxXCuhxPJYlhZSAnnECwhX9nfbS9A9nHClS
gW2Sruua3/1lQZVn1nLxTqLLtFqXWsgrgCLaHsW71453V2xUVQrCO5dvAQPQ
Zcv15G/Jv0TuY0xAdWX53pityyiP8HqZtopFisDKEoeFY7/u6vOTa5FU+t1m
HSfsOV+YVnvDtjhnkHpkWKvNtAzbQRYUnNQsoDNbTgyyHfeEWPz6VkCG/N6O
RIJDe2SRQhIDX+dDnhD7I8EbF0U3DAyMcK94GFq/mGB1pxvkrp/KwbVAYISg
Q3q4WcUrO/7f/FJzkwH2L3VBSzUMe9b8795Y1ptdvTHj0Vr7e4BosV1VZjdL
s4u1dsNcGcA1eC6giVsg+351v5pSlXlZi6Z/PszvF4YeM6d5QL4a/PUxfPfY
C2Yp9DL6KoymOCufYVMnC4eEc46Mf/nJUj8ANgL1mUdPDTDKNgBFM09UDD3V
koeJjHMdWwC93Ui0d9hGVj0bzvPQ6un7n8sJnernCLouTlTSMf2DU5CNMvB/
P6EbOZP1XH9+w1YdNywQgdmy+9Z68Edj5qST4XrP+p9IAa2Lca3tO2qA/+8C
CPxUl/ez5hfD3r8soB9pXSWLUFjPr2DfaOY1gdLXARw+Tf9o5KmYbjjJWoZU
M3ckthyEy4+NFdPYHhP0nFC9vwTibGn15wTzPEi2Xrw9QJMDD8AL8qLyxWjB
duf+1ekSAC3IJyHSN95/xNx44W8XVWp6uBexKnhYaZFVW4zn73izXB89HIGw
2MO6WiyIEZBo77/uA/WGTOJesrEZ/ly4pC+xCRXsMzQKL/0DN2CcaCBBhv+r
C0TzYJc7LYfJmiwEYIomtbZ9z5dTOTcM+DMTPkSJCIaWCMzSw5X8tzWolOeb
1wvOfb4fyqf9NR4D4G6WMjfGwHZTm9GifXsZPakxI7DvxmhyXIea0e22pLk+
fX2yD9DPTdcauxmRyqEKaBumDbHiOjpjmyAMZWhpn2PVVVCndh1qEG9Mj+IV
hwT8H1ai+jzXBZ7JZV5BaGljbZ0iSPT6Qouy9PVdKW638XbUl09w9L1D+J/t
163h7tW0N3hAUVfyqsYOe8QF87jEj2LfPsQtnk/aERIfUhp4ATNHFnMr/yMQ
OxxNVewihoS+46ZB3VWhWqt7hBVOD6D3vCn7DXoIEmhv7mIGWgwD7nIURsvm
UaecXGGB8whW3ct1p3sGwInY5gcBrPLA8nmRMMnnpIafmy/258YmyFSB2vTK
+SnsFaW42o+35GkqoBcHT8MVl18szkBcqGP3Ij985PymzIKqLswv7B15prgf
FhRAmHKNOk5MBmnoDRkxrnW8Cpa7epLmiy36wBNcFvZs7LoqaRJ4s37FLjCJ
lS6NZVnZJ33ntdd3adFZXw3GRe/+8yo9RTCAkNRfcw/uBP5FB0jIdEgBZTTp
qkA6yh5mU9kY+kO3Nz5cNYGn+wcZja3uDONPuW+xFX2EzLA911d6pGniXvt+
mVDK2aaJSfB9CqR/79GLmB+m0oX5Hh2CTiHYIjqs4k8GjD1YquGO2um8H/Gf
aLoCOtz/i9d2KlA/JNWDP8H1dUU17RwmPmuyCMu6nTH61TfP7mCoY/u3zsih
homQXdayrnJ/6oFE0lFtgDYuNoBenO4Q0vYi0Y0J5l74grLMQjG4XahUO8jS
hqfvZsZ5yuJ/R5Dk/8qCZYAuRvGztX4ZovNSUXC422YBGTXTO6ILkM8HV7uf
SUplFzK8FXqjaYUOLPiSZ6GdqhypWsslBhBHFYzxhHDJN+FcL64G7YjUXeuO
E8q/+XS7D+Qhv9G/DDAdTl8rFuja+F1y9z0kvOAVuo3cxPzqRExzpxmqNYkA
8ezgHPvxu2OLuqj8WS6hhMG6fL0X8ymAXii7PDHgfluUaVCbl+q8sH8nP45w
cyVFljnGABvdIQvLKzFm6/IajTde76EqTak/slPxxlYCGoQJbryz1ew78xIx
P3lZCAD/ChEld/546c7RqyT9XHD34CB6EgBIZBDLy77JQtsnmr9nzRGh8eGC
ABwKU0NptKnbIiV8LZbOfNa1uRAwjWaSem+8mRD5eCal62D1nKN9al2BJeLX
qiuH72LJNv4bo5xkOwuOKiVxGjwzx6U03qWyVWcPWst2GOzSEXoigwOOl9Nh
gN/10FIy35OJOlcdAyxZSoqpzs4hk392v/4wrhBqnw0BcH5r31jCtbIvgfnn
Xn5M2dkb6JMr7okM41ybzZgYlHVhIcaL9QGfrBWTRKMN2JQp1IbMArcwr99n
cIj8b8WXb2xbJjnNvRhUbp1yV/hn02zRtccGPOP6nrhXl6Ib3hZ2vpKAQWaZ
fchr7B5dQupChZgSR9BejI6MsbA1xMFzoP2I3Ird26KvuEEewRIP5tLBxqr1
VC7yL/zZcYdm4XchvZabIUVO1gjc1266yhJ45EMrAZ9mFUuroJThDu9JBtAb
3zAWls3js1OX0JdvuEwmfB29IREFH3vs+r8koXrF0NI9/G3z3Ht0CbpRetGD
mHqnTa6u5eJJ4GxVv5HQXOqdjf32i5fETezG+LW6y+MGogahh6WmBHT/sWUe
pLjSchZNOlpgpTNZ+Rv56Mq09zlqgi12ZYwIocC4gVxe0RfhQQDB/AGKhmGY
RwkST/ZsPYsdcTleGNUPN/yq15CdaA47EKN68nZgLbhMduJwkymq5hAvlpUb
Felv9dzmM9C14ouOrx5+XUiiW5mLqOXgF0H+72PamHl5kHH9+pC702UTzIrg
9zz/4kfZwz5gGQy3Vvq5iWyTE+93BeHRp+6S6/Kjl9dyFiihiZd7HLQlOLJk
YpVfoG8AckndF0D3itoByrjKxqMQUisaAHMARdBgnbOZjxmbSqFir7OD6HIr
Y24fCu6IrVbEclRFlP745zeG4CER79ZIuA4Z0EXo0Pa9Y85joX6ENI8cBwhI
yotZ3HohzQ3mJCJPHGypMYgF8ti9zQ9wQE2oJp11001KOdYzihLo2WWtg8hA
l45ddXuqHSj95fxTA+2jeNm1UakN5YAWSWrJbFazaaHqMZkaRxvtiKjzNe1e
TKZT4FCMtJvhxpAl2IlY0nWmrDztrZrQgJeZXjbInm08lS0/DAYmIfVjINTR
F+hasZt4g2QKzww/MMiu5vUM4VsggYSWAV/F99qCqwizBMw0a8HKHbJdzCb0
E0jBj9hvlpMbFrG/bwrVBEEIeZNXtpjpijBmn0uJ3qzKgRORYE+UOnOq8P/n
dgzAtJ+wrRPtnVxgX6AxxrdDHEPDbW9GszSGSN14DfNkSFzkWwh66VkYN+7d
gxaPHIvRA2ei9prtBwufU4oxnXevLCZdMUzAvVELYk0gGjTLlEpQpe7oU/2h
jPwQkMc01kWuZB678mkvk7wzIiTuJzsyRGUFLRhwvj7vt81KJqjD3+dCx0Ai
xaFzB6PEyU3Vjnh5Qv1b3Enb/hz4mcAsesAIr2n7sSkmCsHhqw/HS1I6RPfs
zWM/Lsi7lWtyaemhbr6XVuVIwwTA2IBT9RXH6BLKYn/qvD7y7oD8ibnnvL3P
o0ofJS3v4nvMK/y2E8nFoVKsOQtdalMdsrsp5ZfE1+gxuq16O60759m91nvV
VH3CR933uU1b2AMyXl2cwf7ERpczWkfSbqOSTAPJr3iVZ33uIIG+gX5NVVWK
tAZTIUJcoMvO8HZT/XhFzbo1zn4NxI4rOdq1+3t+iRBjvQ59qkMJLWCtuHm1
xkrCwqpqKqgTRdRKr48pAX3VsJL0kvdnRVuqPK7k3kj+loczZ1X8P1618Xg4
vM7wqoPS6cs0bbiIqI+9KtWe5x+A0kD+U197j134a3cWz0uOqW9maqvncxos
F/guGbVuqvPW3QNM8oyl1F1FV6xw9m4Z2VKJDzyvC3pm6cs3qxo/TLE4dRJH
DUyrGa6aLNBOVVetEGKeVv1Z9S/kL9SfzHQivvAH/gH1tzwWbVz7V6gVNMdY
Dn/cqH5F1NJguA+igf/AofrB+9Gnv7YWeS99DTnGDl3LDo0iyuR7EZMA7oFJ
babccdV5shUEfAuFsUHVRtEcEgy5kGOijV2xeeBkcuVg0kg2SopDTdWEwqud
HcsubcLZR0891tkOkdYDl09h0p2S1BjtQm5sDDOqD03e49kEpJB//Al9+mCz
vxxLAqymeL+dFe4wFWrPhQsfyPSOGF266zmf5iM7pv8xbIW+7LTzgYixQEAY
d7TSKtLbE9GrEeRoQwBx/B8uzYfUMyyVp8woi3qACaxzXQ4dEtqZvxkml3zq
+qUgi6nhK9HZPX35KJO7ToXI4JprUuXeBeZRrHayOUBXFfu2I8peY2+78YdF
22mlOnbJ6dEWtIczW8+9fTEL4hDXvGYvv5dJUIH7HmDnxuLVO4s5N+Mn6ETf
UAhRMmfS13FqJ8quOOxhxrc//g5czRexI7yImQwWtXRGt6yDcIMPTrmNTCEZ
3/ZK2qXCH3lQb+UMQ3LTs7GhTXufbA9F22ScznMR+Rrqs5gHkd/ouo3NXSXV
ss4sfOhdi9HbSH7PRlXfn/5LYqpHjoVfL2gE1UljEXatXKt5ZP1TZH8QOk7f
jMk8MczyI/3G+U3RbiXID3SMPE63PaBzQQemObbRTygLp4TN6mSWAY84yLLQ
P3v39dwSPA1OR2uu05uZeCs7x/6lCePwu9tVKfdzriJHKiS9ghb0burRU2dB
jTnfMW870WPAyoC9KRdpK5GhxmPebz7FeJ7cFIUDaMV5/+HLhZ2hRgKW/T19
h6cqtxZIdU+nmQI0cBto80diOLkR9U9zzkZCn+jn0GFaUsJpknMhSiFMIDf7
MLQbzlMTNqsCDOM70qRI1NO0D5hzqeIvymRGbZWwOD0yL8dpbTf7Cdmjeynx
hcc0cL0UTly6gQexdR6ehzCci4GKzdTnokoRwNbKLFZEYAWr8L6z5c3+Mc58
9jOLwpo6MPHIOaAPNi1cXPjJ8mb+/XgnmNCX6aviWFvCQt0C78hkHS5l8uSa
8somLW/Yj3khu20ancu+xKldet7NxL1W/CQZAv9Isd7fLZrvU4Bqfl5eIdGg
L9XtB217wMjSMgW3Wkcq/0PEcFN14SmHi2t1FguuR/q8XD1pRDYRdtnk4P/J
5u26WjgtByhyKNP0h7VTB8wkg3ObARiwLEsr13cTNTVjIPOH1eJyTRLFS7wN
2VbLyfPtsOOIeJWRjmZ0ScGDVWUApXIMTf87IpVaHtGb1V0mhuOKlkoKhm3k
qyiQUnIRlYRUROIxJeEKHoK+USWNdMa5uAqVt9OwAEZTq5a32z83dwuA/KkQ
Sudnt4rIP3N3Sh8nkyKC6gtjDcFq/GMLpxFK0Z2PoBgFdJllpQ00j+mIc1Fb
zSqXOYe+pMAmz3qfIgekO7F9aoOZmo5kJIKx97K0+FrKKwbo/V1+nJiNKQ5H
Lc4RdRvVklN+nEjtIfW1d1s0pRhfd/xpQP/8BHzUceWhv65mvq2NAxajqDy/
uQkpgy+3r1RDJZiV8WWKPrN2cYkBMOjPinizSOuKrBp9p5warymiqE0zfP+p
5Ei0DQwMhb2SJAvsRSkGZXZPd5NYb3lYOHrHtHzuWzkpje2qfdU1d+Ec4Jvq
iMiX84HwlwhmcNLVWCFAOyOn8ps/prrImGMoxxusiQZ9mS6vY4TnIuDt+7XQ
nJRZ7+Tr5gzHG/4lMhgYuchliN3+C/NYDJg7zbePVLHlqb+IFOXY9qje7noF
IgMehiAhzBAcVnYluvKGkDVvzzbHz64O6z3nMVNIKsyWoygBDVFXKgyyFMuK
QMtz0VNw9VJX/+QPHmz5YfVLk6MNqhYKkVHZvlGCfrz5PWp3CAC3awDKEk6/
jjvC4YtQNnBwmL0BhAS7/XeXduX30kjuJTUDA/V9J7usyffcYGVEHSIFQBkl
IdLYAjspn5kkGWmrZmVJ5dDbi7BrZv8wNmv2jKR5EjvqaleXsbJ8hXIbb15j
aTDEh84xdt/FnsX5zGMHL3Cburq45G0vWsmpHj6cP2qtWuBHOHGmhvhRO7Q2
0z7dIPs3Vur311PhmeJPg2BxAHnC1xV0DNhrKTCYr52XgwnctvbVbq3iMx0h
SikuRnDwoE21bXjeO6ZfJDf32M0QT8qmPmXKLyym4qIBjiEgrlhAqg1ZR6w/
zkg0md2PZY0eHYo5SsVXd3PjGsdM9xySk9o+sXesA+jI545ULev7+pMGdgEp
tR4X4b3SPSt+EYOOwIl8jDtudnxDPd+dh7xQ5YmPFxbtEJLRto8LGozAnpId
r9AslnmrluUIGTKxU0+qiYx0az7EqDXSKv8vvnRwGlvFzS9N19TnHW7Hbtma
kgHOvKLbs/zWLUEOnxHyvtL6u9G6CG5cxdrQpGezuFIphgBlwTziFzgG0z/g
oEY2p6ROkVFsSM0l7mPRmU5ZPrkBo4+t8JNAbfZEwpjGoVLTiX4wP1h0Ttaa
0io+8NXlWeJxdfYrDIyta3T2NhRo5Tv2JqJr/8UbkpBqSLD1REXC91ZwxjvY
5laRjbWvcYomoU70RJAQOj+axHAfXgqVMvOwRIOwANmaPgtQugw298MowsPV
S3HVp0c23ZN83Sf+8cO+rROENHQy/yRvHhxygs4yyLEnDoGBtJL2Y5CWqJ1w
OAaTuWciJuo7TryNimx/V2tM9wn2rBs9oV3X6Vu9lmf5z8cLMtBaAV1UbTTU
b7j+hPzK4V5V9zurdwiajzbDCroVVShvZoRmXzZTLhilAgi8enn4u0R/UY1l
YAQD2JgrI96xv4Eh7LFFJA2d5hsilQHPQD0jbyZ7UcszsTNhZJC5aUb34Ia+
xd5mj5RJsZt6biFka5vBMmL/pKsA46lrghOX4CxgAoxtd6H9j8tCzaHVMWQ2
sRo3dYxQda6r8anCFNTxH3FaTcf5kn4+xDP8dzKPDmvqxnJ7GO/ayL68ay58
S0C9yZD6g4LuPvBXFxEZCkaCOwu0UrLjw6NNnMQe3qWOm4gOUFQ9rKW0UDm/
GqmndgZq0RZByfFJZ4kUeOmJw7RMdKQ+pG6nVsEO9kZK0CjuYyxH0Zm2YMRU
EBXzJ+OtCxhOrPruLXCh2tiqwmhCcJTzWHZnKILIlzA2vMne0W1g38b4SejL
bektNp8PI57llqMW740laaXsUtT3Ffx4vsm82BzrjzlZChY5w/JmlB6ms5ue
rlV3FpesiaS+EFqzTWwaBiDP+g+WfZutq/rg3qW8cdVwL9jb3jd5zYAampBF
uv33R6KO9F6b+CD1eNanLA5F7bTv1EEBglOZhLr8Pel77MU0bXzYFykVHnEF
G1DhdXm07d999qmQA6E9SEhVZPl5eATKctwgVFl6WTGklXKasznAm5pRGXuh
HCsUNIEgUYEZirMEhFH2d5ijwlb3Yfz6fqQ1KIUL0oz7J7FyGjIwLGSDQhOc
bUDT+l7fKAT72HSqIXcv3Sgi6eLw2wtlMp17jerazuTxMufnoKpKGuZOcgYW
I6XJf0CigwPDTSCmPWv+43gBVUoC2kDV0xSv5Ts/vzenfwxWRzU2n6rd52Mw
sKvyWLOwNxnxSoDq3qaydXpfxRaGdaX0mblnvUSbxuFj1qsFEKaXnZB6FEch
hMmoZvYvrFn2EmDk62UfuueWOuxQH7p59oRDJzCiR+84ujPuM4c32dfaR7f6
IiAcAia+ZxxzfopUS83bE5zK7VjTnqGT/a1rC07woom4lD8o0j/sGVwzfK9B
H95XQWL3IV05Zxvd9q61tg0rmEnBwKiYtY2heBewP3stJvfoGG4AMgmB8ysR
jR6zCi2sUNXXuEF23sFHiAhxYSjzp5iiWKXZVgEOq8WinfUAeXA7xFawMoBZ
I37PRylJgFWgYWdnthGODxNh6CJ1qe9K2cas0tvWC+U+9B8IhDOzpJ2Izubt
CGNg0f3RgWKDEvM2/WaYYtpomq+cPAIg0Kx6CtNO61ZQF+dNlA5ajG0EIxND
Xl0AFLTxfJGKMMP1crlbsM5oFcZ5cm4csujAEdgzmXdZJFYOV+mnwK/HSJlP
sYaWHKUoCFVjnWwHRDR+RuDDvoD1L53OtZIo+bbR4XpK7/XB5eYHyJOApjbI
Oc+uRXZt2akOxsV2dOkI5yJoQbFY50+or7XICZj6QGefJrWTi8GcjO/pXTxW
tcKUVcweEAx0RQIeaKH3T97it2wgQgcfH1yxn8cH1Kq3qMmZftYicg0mkJqq
Z/aIU5Hc0NDjYnZQStnwKTPAO73MGurKwCF3/CS85RqaJDbXK3AoIzsTTMPQ
rMdX4jIV2wBu7GnvCZDQIsHRMKGaG1tK4XRbBaCE78RJ7a+h/Ia62jpup1wQ
cC5A3t5M1ZTdT/Gydk2rJfCGuM5N/VpiSSuFPQhglEervMgoGt98MyRZTLfW
46g1aB2pP6JkBkfCA+TmDRGkQx2ISfq4Io3N3TbK5eZNDi89NEOBP8haoaLg
JaHW9kplmYwEf/5KxzGu450KqyeZrKQ8YbD7CnJEsTg8vYvHpLmvaaaTYa0h
s3pI6m+SjZMO4C5w4IIiDD7mnfU8Ci4s6FusJhf0rmOYx2SWOtcfJWaL0srM
oghFS3rcyZJcYIg5IfcQEr6zdl9YOdFZP0i+C+MkAW2cY2cu0d9iOexnrDld
G52gYI7fkeRzEmGqAuRPMa4ztAa1D/hkVAZkfJefUbaKojDWcNW86tj2iBGe
tQ1PPEdfFH7fcwtukDa7l2+EMUNKeScH0hvLM6dB/eQmiREAuq3izTcoILYm
r3iUV3gurzUJSGODZWpOr7XUwhGtEx9raU7IE++tvZZL1xKuV7U1ka4djaYm
1sO9J5BfuuxVuBO3uMNryDsbEpoFr4b+Jc5/uFrY1SZqOY7zZpP9ENbzw4WG
wPty9xxEyPxyy8vnaF0PZWOScc6dzKssv8CeroWr7DfScgKba9eOZp8dbJGu
sSuQKLL47xtUZhV4gGIYyxiZ3FHlNzX//L8PLXvsTEwsSkLMBiBeRvoQ2cFG
zVJWQpejRl4gnn9qko2TQ2kIx6MyQOT0TJJmvXXng77y62FWmJ8Rkc32tuKt
T/WpkopBl8rnKZkNwMEihQi63FDU2izK1nIY27D+ZImJFDyzoNnmCDH4yEI3
AM/5DsUD5IkqtDCYUcm9Y9sdiKj26eW2Zu9r7FgF6o50xjtli/ZNJx6Q21ES
FjKyAaLFUhH2SeBPk+Ax04k6NUfKTdVl/EnsZysWnQoXF9bCs6eLy0htwKNO
qomVBzj2uXMZ5tSrrSa6NUTSuneJpt0sCOONNrO4x1ymWnBWkX51UBQVnr3O
e2LHf4YKwVMYEk32F0pkaY18MgrOKvrjhayZaD19nEvsLxaOmWVTrjIEgaoN
cFl0qr8aYNz9eTKuOiaKBWQKkm6+EmbUqpNx/G0ZHbI/6by7CdAtQ9/29D6V
WYfGhynIXet/Ld0VOgQTEQSUsZAic377BoO+V/ig2S7X3LI+7jrm2hTpqSKa
RMd/X98g6qP6E9Bz1i4vLb+jZfaq7XesTAj+or7Nus45UciIw0e5xAgRgW6c
X4uz50A6TQ31A+YWd0Srs2mUD45ZMXeofF8fJdxDZFMVeIIkKz5WccMZv3iB
vTRBJXTdQpX6cq9JiPUjTSbr4CHTHlq/yccXtSMh97qvpLUvXHaPyga/jKWE
Lxw6PMFG1nOlKtxfl2/4xBfAnebtKyMUaa4HBoreNxirEgPsuwWb9SGsFTnn
eGJop3OPePL8T7gUWn+BfbSUH3mjwMKma62rxmAY8nz+zbw9IPWuOmGainTU
A31zMIDbG2tQFZm6XuCx6CB2s2SGNljHAPt8+VHbmZYeKoox0G9l8RVuGp6W
fiEpiB9TXbkBLq19g1rDG1E3XdHKd+kAvele8bR1nkphhDXBu6tTlD8dSTol
VIqLmdjXUqnEBBt2eQOMezg9z1ChVTEgrLt/dbbYUpZYLUaKmWVkt55hK8xr
UJH95K9d7RSyFNuFBSUbWLLAxAoLMEF07snPui9yv2OIxEP9ZsgkWUPNt8rV
xxD9sQH+/I7MUzFrVwuOgp1stmrgIldVlC70liVz3AtLP6gB2q4ENE4g5HqR
SL08pIjxuSyGE60v181IximB39VcJ1B5xJpQpHYmOokGjuZmh8nnLFqzviR5
Zm/bQzEdao+Z/l6mhSK+KdJiJNKojrPNcpoNl0ncL9IMUmRxraPieGeuzMt2
0RpuLzx9kMW138oBs/iZmfT+vI+EqL/woCV6zacy93bLaLOFlBb3LIlDHqZ9
zh3f1DDOPgTUgrVUlmchiVRlUy7Ob5kJq51u5R8wGsCCXE/vjlfK7sr4Lwyd
ORuw2iWCM/lfYSjUU6dYBwvoLQPu6xjAVamFo8js6d4VyEw5//9GV6jlDo2/
UzJTkJ1XnUd85rVIFt/CSadxJUm5oUctIyvZ8FrZVv5Kd7i9S5PQIH3ykvby
IvfF7nTIIvx1Uw4HsBY01OmoBKvMujKweDcdT+6dEnLEeGJc55PteBa1tQ+G
dFLRtnvg4AEygjge9NST/VjLgfRS6X9BqZ+PqmwJRynG/krYj/ptm/nzpG6c
sDHf8BLranakWce2FTfj/lYn71NDQNc8R0TlrGbMHfxPceMxmnwSv0kKzSo8
utbns7rW3fDbc3CpuEtr414OvtFBFDcYfNhId980meEUVjcl8c4SsMmLiyir
G9d5F2qSqv/riYnqar3OI/WiewOhnLZs1jLcx4+caZU0+4s/bEB6jT3KzPSs
2KucmVWcjziuiQmbq6AWwRfV3c3gKrSYGPvx3a/ErYWkojLYV6iNPvwPqP6n
TIttQHj1Wqw+hObpmy7eEQZ0XytJpeCqz+83kK6GToO1mi3K5ucmAj7KLwjh
PU4P816jaUlgd+idbboSAd7GWMJUmka4s6tnfhl2SJfdd3RVHbKspTfBHxko
esxUbbP95vvPdV1tNU2EucgFZrgCRaEt0XciYcyCm4nECIM31CHuwiHyHSl6
0EbU2Cq8fWh9D+gt9eY90AfHzUUVVKoMUWyafwMnmWs/8puM7/Shn8MhNJa9
HZ4wyJp6lam0idEzMi91/9TKvugVkH7zDyeCogfTRDU482dsF62fppZcHrqM
/Ayg2TuaJynGEYI2koLuOWmLe5zvJaUJ5eCw6iDneF3AQ/iqkt4bLbuQwKfn
uinUpR2+DOEmwsUDvMmdW5P+nWrSsG9cut8xWcg/iu1V+I9drf8Ws59K5esB
60BgcGwr9UyjSTXa/AAlz4CmUUjf9CrQudsBRQDpJYx+aKzafzUC64w+Jb74
IjAOPaE5CPQyNU+e14WQy3sw2i7VnKqT3O5q/83jcbyo97BKO7yMcEBDtakb
T67P18tWL5KF6ZRlY/lqh9ZmUAlLlTuzj0vQC+BucYE1sD9wp5oMz2drfnGl
U5gZa2zGdK+u8ZRCZlCMZuMzQU2ley5bpTnLFJxk7wCwDl96HOdF9mRUoP7F
c2AE+NnpR24w7lZ75iYxRBS+ZlpL2S0PY3JUWtuxzvuSOXYuA7vvbRWRG8YG
jqDDwbpfr/ZwFgR+XMLSTExVZMboazoQU3h0Pdbj1kCWAFnFZyFRiKBXq9Ez
srGFWjgiLavh5ZXvNw+QDEIbeuhKSQ2mQz2eIL7BLHryl15oco9O+X6sFntI
2OGYaccM7ovBuwOPkJJLWmBeHMxWNvCuciEOfGIoIedcbQDcB+oNxbLMsKS7
915Wx4QAAv5KjEX80un4fEf/5bA0dN4I2pTgKvLUOKB41CBA/zmkm4Z9qj09
rdZNPB4XEhvNpHkXfGoWySijYBBpX6kB5ncc3Otyy0lLrNecK6NeCvbMxDTF
A9tcPP/Vac99uJShYqkZYQCGMCiVu/a2XCcEsqWOXiUQHgG8IQg0G6lyaU+t
0qZYoy5DOWiBgBqfn+pmKOPSU0q3wztghW5zzOgsIlBb6NqjeLAj2EPp1kwJ
8W8eyPTDEjs3Jw1JrtPbe24BU/F7PDqK4MpeDfK7/pKfqCyHzZuL5UUKeVIj
MwCjuWrRGueLH5jNNIwNm/0BvC4FF3zP93WQucTWQ31UTnAAd/rt7zwfed0A
loVqZIYBQmzG2D/s7OEVq+/TE8i5/CnD4dF9LQhcCLqxY0i1k2uM/yO1256l
J1mqppReeKlBfO63+AR+gDlmclyiV8kcE6RN0K4Y3l8FaXfN4nSBYiLJrXPI
aLZxPp0gTFEiA1F8Q/uSRq/Mm4n+nwwaoaLBd8yDZ+w5FqwgtacNxcKLhXlf
WI+Fpix28EMUdNVdpXsMSiKgyucepdzHpyXmTdf19c0Ypzg6AkTIUgMtEu77
oz/l5KxK3JFxJxHxjK31rflBtFm7zt1TFIUp8M4AIo2/n6lvUOubq2xxXeBO
DnAeBL/77aUvgDe8Iry/Yg7uUm42Xp7dHLUR0gSmXuTUICkHhX0UeKTHICLR
eTMHRJtDbRppz+EyWu5PI8DWq18mNLC7vAIvzix7BFsWHHPK38EL3XLh+VxQ
4ZwIHIm2ZDB40+a9WVSKXd5n5fQWxhRp7j9/DmJNjyn1AEImYH7pySoJOKdN
grQWwaPIkYbezticit/hm77km7tEYNpUihzUgOOyvn2n8iV/bnIFwEVngNCt
qJ9mUShnnA49strTiY9YWUxk1rWP1fWg4U2zGBL/JvzDqO1QWWNRa+xIO1eV
aUBTSgMs/dLb7Iwn2atzj9jIOubFUuJmChPIsKJ0KJhkeGkg6pc3afcsm/jE
oUM64mrMpDS7wANSSLI/z9WUcXSwBjZ51SJ7hzxM+NiVgRoSIk5rH2etfBYz
atoh3Vr/3plEtJ6Ts+vImrOlBDRk7QJ6BJdpzXiK6LWbFjv1YSY//bnKU8v6
IEhepkC7u27BjZeabD2fB3Uu/JZrHVSHDjcPpzmOjKKEPcjRay3uwpZ5pnBp
5Wwd5RfO4xCfOt34G13BTJ3DLQjbnCeDyVS9FpAROhnPRnuvMuZhT/9qxnzC
yk3apWa6XsoR5rfvFU/BDHTHJuj27PF7c36Eludf25Fw33eMF3OeF0A4C5qV
AP7/LoKvBhd4Dy+hA8yTomFqyYk/w/6b1sduK3t4H2BlLZdBXkQRm2o6xrDH
hQ71x1hL2ZLzRu8JD/2IEY4az6paRtlDDVV3OAyqotkhYGM4KW3GDZj3Hb7k
YoIHJjPXdh7q/DdguE5io8P3ae/mGihZfPicTAiRdDapimRVEFitfVYH9mWD
aBjDX9J/Rt1feHkvZ5K6M/i9axKAZn0IbU7Hpi8d2M3vzPVW+U7bHlXPkC3D
IZtYqHK6eO/wUp+1KTev86prdZcLifqtynAZn9j6NKVLR8ZcaslpAZ0q0yYb
Cu2aRebCsDsK8pfY1B4PvltYcpXl+k6UOLGsbJpsNJq7NuZhXjaNVpugNeNW
9HsRkragFA/n73InxfUDLelvBXt7ayiFgc4piDtLVBgMbdmCkGIC/c7BuQRf
3eKK6CRY1ThDOGDAbrUoguO92uykYFF5SpSFKVcmULyNMpQS2XzNXqQhwCEe
5DyQzW1nlYBg3pH/QF9OrCGGkVjl3hDxZLIPuwFPHDgjLkW7gV7yFUTkIwys
5Rz932OsBjzpvg+4fWV124mTC+NOlN/xbAotO1l/rBvMtsLq4mt4PdHz1yQX
RrqX7+gYIwcgLmpH8BqSn4HYkevBrAvl8FvlvJ4sO128Kaw8udcJ7Wd/UcAW
fEPfibUB7KHsfKFlX9Qt00QRi8685Omyg6ecLa9Mj6sLD1789undCRkROqyi
tqMMxxRrB4z7YiLNrUV/n7gHYFUIBGmEG5kI1GDnWaxFIb8B1f0qASYI5zVq
DffRAnRIAZnBonGOiyAqBuoC328sPrWAiRquvaxxzSsZ7gxf6q9sSromEyN6
bGXka3vdsyZIjQ12OSThh5Marh9goBDDKla8PcZymZL7SNLfC+HQbup+kR+7
6lI7C0bwxdG44zPLG/SURluGwX3jLh0cBwpmoR09WgQ1avmrr+HpRrdKdswg
wQOE5NmWxRDRtKAblIZBG4CySNy1qBD9/FXAuFPQizXN/qyfXlD0xnnd2NwC
O9GhiZvSlSOwuhPLwrEHv7yUMIwua/q76nYyI8Yg2tvVCDKjrw5nF5mAW+37
GYfgUSwAI3LuIC8pf58eG6zoUAOheG6MDYEPLx3yhpx3wwDwO6rIx++tYiv8
Q9gjjpiLamHK1WJfHFNeai1LY4jn78N3AIH5GWm7y/fcExB2RisyrifraWD5
z5bVNWcHO9QfvjqwimqGC/ydsEFsQnH4g/epz9qNqsAzbD14OmS5MmdaQydt
XHDwWR7I40TFoxhEEwJUuSpO/ccc49blcFGiMXHVutKeIa0++v1pZDcMY7D6
a/oE/lqZ6H5IMYZBX0KvBl5zYXE08LvZ0rqlIT7WTcbRPj1n6wsugOiy+90k
yT7C8ymFAUb1XzigDln7VZhHQ8SCQwoFgCpWW5JDI0+4uB1qD8/sc5dnddEj
5nJ5gbnOfUWmFIiYG9EftlkotcjSD1dAEMS5GR09KOq/OcXPePqtmcVOy6Hj
KOx2xOrW2vzvZIhuDsbtEaS7gjt7ps7tInP77g3LO0HJWRnW2HxGGGpbKoFw
t02HrxoEH8M6BKuAo8euKJqaH5tJRptgJN5XVl9VcKLtVo3iRCUDg8FVlpib
dxajN/zEyVFuYJm/Jpq6zxsA2o697gYCua/Y5xoT9QeYjIivqN6gps6Lj6cS
kct9aQNo/svUQ7NhLM9xl0YJxlPLVZzFtSAj3XnBMtMLdAly9IBm54rmhRIQ
sH7OfBNpZ+VObxBh3DYGRSlLUdvGW514tvkmspYdXGON82ocMzPCwRRqb6bF
0ngKgmjuv5pkV7BDfx8QxKaa0eAGFGa4S/bv//Bbl1rzsLB/2RWWVaeXdNzZ
Be5V4wR/eSZ4pzI202aYfX8pf/3AS0+5d251Uc5gzm9wH4gOn8zAKrjOCpY3
EpGYru+TKL+O/j3aZ/WFVXluYzI8VJ7k6xn15PZDPZgwQ0rj66qsoYHXghRk
XEfRR5sddmGcpr0gRqHxeFkLmy7kxHQS15t0KnwrmQ8PvKz71he+JHppYDyI
Ol9KlAnqC7tN/HzdvGcQh+WbDdVQegJMj9gRIgb+Ls4OWLXYYnfOd7sJ5Pfj
3+PYRnKGXLpAvs5hdauOHC4hXDjYta1m+5NiIEEa4sq9JQlEY02+HC/J68U1
eWkUnjHTrpedHGbpsbBF8qndbVVo0NusfL3v2NUMuGjr2FeBgVu/+P5JTi7F
ecteH4vnoMkmU6T7BwlUvg/HFKopzWPImhz0ebCJwKxVDqLwlXD9/7LWEbqq
bWLOxwzMve+CrdkfPYojn9mUstB+c94CWTAifjFHX8uZT+l6zclaCndoNan0
nsofrg4+U78hzkCkpvtKoBkNR3sBZDk/6gQxw5N4Lu0qASf2PASrl336ACsB
k5bS725EDjsYxShwIUtW+4wOqHjPEhY+f4JaMU5Nm/m0CfPAB5FMQxIO4wqG
xXzsx2SkETVaANJJxBShJcPJ0hS/at+B3VoOGSfcuY1GUCL/nSi6+G2GpZ0c
cjsMxSS2vUJ+0lXjn0B4XHefUQK6Ndgj4t8YCC9hRvHptfACf+E6B/GaclMS
ls8sIrf3Ms984eK7DH1cdyNErQH84wMM8fT5QSDjZaWDkrgSKLtFp9Z5AcGl
FVichCRt0+zBlhWq3p44L0kMgrgNVD/PQJHynsuCWRSC0BQlcVY9ezTqAfWF
SBZMDH4+JaCd5eTCvvS+8YsKNW5swPx3BJ6+vY+6OR8JK1HNBwOAdE/1Tr6Y
Jmdfm+ge4rFmcjI/lgAd3TT3ETizJqb4e/4LMZGs+Zd4TZEMq58U2B9VpCMw
/6m4ISQPmXleu1wm3eggnDPsz+Jr1paVVGI25MQkGfu+8EKuVgfBPGjgUlsI
3sbYLLctqsey/dYU6WCwGdeUqa7B/bLsq56NerlbBSY6iM1dPGDDybcfLLDD
2wZ1I9gP2Q20MVA3prR19W4RZAIOL77lvR5LdnEFyxT6otuWMF9HZ9VyZNzr
dMqIshFqAnRYbR3uL1KuJBrR799ATvWCOM2bmiHFIdGWEvpsoGvl7lnzd/ar
/YhJYdsqmsVuqicALV1QhTifwFcJR6gZQvyuxnQav2447UK3lprjCcmo9Sxi
4wGJBqjUCSaMuzei0UQD1/dTOsHplkQqyEruIvBNiX1oR+ohPEPfYeSU4Vxz
UhUAv7FJtDJQ+0e0f1GMRUQC9Gc1j246AbtgMg4UoYqeRdYLspfenakOtujT
7aVfcgRPXzFx6uRun8oCi7/ityLHu4jCl9YDfAl1ux57ZfUQKGY9HIY93kkq
0OOvnleCJpC2humgzZu72AUvw/ONNN1UQV2wezkQHNqao4u7ZRulP4HlV0Z6
OIa5G1H5Zz9TbMv1Eu8s2ZjsE4qmp90DP5avt0f7e4STuVg7M+u5LJMg9BwU
TTASn28NmWKQxYeVZfii9PmFoPgLVKmmUHTAig1bM+FzG6Ecg7pjjiV7SpOI
2OzjZoN/9U2CPfJ59+b6UR4NXvLId/o86tJnUiUY9DF2QOPC9sCS+nJ4Orxn
UFdagsI84PpGWouG4FbGVMHEkzJ8k7zgiHdeDZ9yMSfbs2HgNLw8wOoMKgD/
JuVihJcHGNhsT2BdfvzXRrC6N3iTB6AZ+TCYyzBr67VKcr/yzrfyb+3YnRak
UrMuOOG9KNLwTCF3kGLdJWOQInWzBRZBKq46JBGrElK0e6EksPHN09qbrBxC
3tauW3jsIlIlGtigUq8JjRMGNzB3RRhjz0VbBo/RUCQI26Z8gtnPc59igpJd
QeKqAT86FRLkafb7vPqnDBWg69/c2Qaww6792B8z/jGbvKs+5ujKtYMKtjka
hnbFjov65rSNksqtXK1p6KTJUJss1GbYLu12xn5k/N806rIalUNPnum0uAZj
M0L2CJkCoSX6VE7tNMKsliW6DPu5yYXfa3eqcms3hcj5Su9hPxeJc/4qc/RO
LAuBcYi/gEhEr65P1Zd+UjE4a9U1JDQ8NmVev+GFYDS+/fNB/BpuYgLn8Dbn
QhcVt0bLwtS+FIinejH+WIsaDIlrONT8TMX/88WgzidxpMsYQnhMJa+1yp8S
NdM4x53PZUFlaqKfMZl8rPzHkWu5qIWmVRKnHuNHhQSLI7+8bqviyDfedABj
N10uWfv7LXQADFUGuacrLZZ/hg3c4OxFNUQGA6Qmx2NrIVwptep8jkB/++FZ
nGt1Fp1NxrI96cBwtDNVlIVN5zkQdBSBlxsbuB+okxTRfUKoAA1h+6OIwvzv
UkU08YIG0CdIVdSLC1et+WUGZ1SrVGuDUUiFHS4JjDUTEYCgBSwmWIPmA9Ke
BlAuHTpMIU5AglSTZVbtr+nUJ/snST4eFXxw5EuHyrZ9Lr4cFGe1L/EA0VLk
8eMdQNWxk5WXrQw41NRQG3xNnj2VXSyb/yrAeuyFwfuw19ISPCMkJyZ8nVkc
67gnAC8a1xEOhZculYg+ROOKC8fjehihZGnH9QgfR+fQkYKjH9e4hOKvX+We
9Wh/fmJHhTtKuUIpjxc4RjE/KV0A8Zc8disWb04GZ2y9uIEzOoOmxw7fy+Gk
zrWjgE7kvlc0A0kKU4eAb2sDd4Ur64dSgvz3wUaOUKdCaoZLLX+3TYETafvR
hoY5s42vwJ9XhdIPTor8c5mXKowcjgdBS1IXIxh9CEmAvrxFDi9migs11gXN
rnizw3uW/SlbTrlKm2PdCwOrTa5fspYespxzLdcoX3d3zDVkO339FsaRgWmd
46eCo+wTLH8wxwMFRFwuCO8R9FZIrrpx8wgpfqMYjjzwJIY2TeaBl6Jvm1Ch
9QYGlZ84tbv6609u0bWeF43xVGmsWAsCZNlKPf9qAq7CoMO9MMLqccJHK+yD
tg8K8h+rO18y3AjmFRud1SXSBln0cuETuLI9h/pa2Jp03XuI2vWuPMB5EY0s
N1sJg27NHcUnalMO48vJBQ6Fw17K2IVoMk7rIsdXnbst5hewVnVgboYeL6e4
3OV+r8HMuY/vZ/Ep8ilKPdu+Pral5dVMqx1gxAdosaUFHX/dguguhu6J9FUu
OP1xXn6v8jStCIUTxeLSez30Kv9cYC5jRuKKrvyt0PfkYxT8LdnY6Nt9OKPh
TwDPUHLbMBzwKk3X1EFGPReKR2YQE033TNDs20BDEthvEKiGVwUIkxClUQ+E
qdS+8bWF0Gms/qj5kCF71izXKP+kn2MPeItL7g56ML2dEqgurV60bKmTZkbf
o0SLt5jPwHb4xQSYvXNJCzUc8QEz3CwrXhtUw7NDHjmjsTMFx4lqi6UPLGqD
RmKbYJeI/Yh6ROAHFbxqKejMRFT3WcjkfcndidlVWEw5n40EtStD490W6d+p
O6tEs1B3bwaugj8dy8+D8DLHHc+FmL1avn3A0yKqLW0rJ/KP0fpbRDXW7lnC
cyH2PZdnI+npr+VWex7/Oq0RPPmKfoE3BM9vXFV5VgQOEtn5iFqan5PRnNkZ
f4jG3vEEyWfZ1clQdoB8pdGWCUS6L9KroACNQfYZiVf4dyvaTq3jlr0UWjoh
85P0O+rDeK2KgAq+Rz7xuIjzZE0BCRw3tkraVkmBLE5MThbm3QV32RWbNaaY
IPCKhJeaehoaLA24ZJdEUWmQly3ZoD0dtSoQZLx/Pf0Z+hu3vNVvKTk77jL2
aFMVL/ZDh2Pgpja0oCFkNp+64/1yrCD5jRwlqGT4XQupZ3GGXkYfSIYM+cqq
iU4sYuu9GjL4wuwuJ3Hm8wU4KZTN4stEU+aSkmGsKmzLAvLejXP3pWZhzXu9
zTJRuNKA0BlU/TxoC5cG9QHDpSVtbykOVL31RulJ0oYdnw4G5xaPY9z8cPoS
4tQNW7w3zgLzuQDRXmitUKD9iqgasimtWXk0VFS8xqDDvR9PvalAnlMFWWmq
y9+Arl+qdIvr1n2hLjaJaJLHTknTAWuEsvU7kVNmgmUoh8OqiK62rT1aU+ig
YjK47sO2VIIqV2GUUFPozLgt7tlGH5HE3t0RCb+h6p2vmXsWCk43GRqSG9JL
6HEAn8eOV70GwCc/7ePPtFsXGSsTxj9y/hg4MDJA2z0xFB+/KC5D8/vEbB+k
SNRKS/szpqKaQUbHW2rBs6xNdfwCSI7TeM8TA2Wxij4PKQNMMxVdBEGsvssK
Jn7zo+ebdjI8nOSDHnX/uM5brpXinXW7E6k0/wFNBW4AOtVaHHg8PwFZPXE5
S8nptiynS10oQS1SSasv4x2bA0T6IQeJPhi2afJ4rs70SKkp1+Bx3pXfuIOM
RCVWA4SeSYgoW70CGe3YTpfjFbhneunt5NnweJ8ZEYOvkD36JJPFUa6PdY/q
5+yuRfbQ1uQJ6YIrALq/LAAPfCFUtdQufSP15XyJrQ1TLyDBUJdmLooH92v/
8VnrnjYcCpu3r2Fw4yVLEejFSXN1Yj9O9yxt3FjHx7IkuTb4kspDBubO74ay
sKCNKgm5XpL6wwzVONBHyj2qkTtmrDpYDBFQnLtsRfYlTHsvHXskGIyNAWM6
/8RjuknrpufLYpBI+n9TexE8ATLDmP6nW/OIcMfFtBEH9dIn8WE8hoPjB0ci
DUmYyA2L8bfC4lcBBP0WbRyR6Rrm6N38eY6dCKRWi4rKvwPcZf1Org4S3DhU
uk+m47Gr1VRdJZTXU9DXZ9gXq5zcs6dTaydIN+RlgRZtjTXc6sCYrtpGz3up
Z5/dIu9dufZ8K3J/djRQRKODtHutsst0oz2mmudg0dd4DeEksj4P7aiDLePe
q0NSZoN+iNA2DA3nGkk6j5BxC15K3GtmN5rH5/wCepG5vfkXFV8+vya2xgPG
TuK90V2m6jRTeLwK2yN7LJr3p0FJ6kTlOXSFfMpxNyoBJYCVNq052dPFNYnw
OGUpH5b6065JX2c5tGanC3vHldKVLC23LHeLWMKp1cjQ3d0bixDHOaEsvJpB
NL/ZG+yMFj+A7AuwTQH7xwpNB1W5kJTJ2z5nRmHVC9V/2l+nYkUi8Il+4pz6
Zy4jYtrCBunO2lovXqNgDhHBzn82HD/p6NPfaE64SHxoxlz4xRGXlx5jkgOL
1b2DtPJO762I9NMbdnc8AUDj+iJphXiwiLlLIB8hSw59sV4htZgEPPlkofFW
+KM2sTY0ofAvYNCxL+XqdRuMkkgB5KCw+QkN+UMPofslagvO/wQpcc4xijl9
j/Z5NHQqM3aC0Tnnjb3mroOVyjTzQcDTX8d5rF8dt/5702iaAzrMmiJrmD1N
E3uOrtS/KD5JYiTxP4H/AHT+1Snf0bDGyp9p8SB0IY5Aj9GTuRd5IyJzJEWH
eaDXU9pasBByk9GtfwyC/SF7Wb0b8LLN0L298VonYXRTgdh3ZpmkW7hm4rvd
dxV/0XbCBq3DmUU24BONy1ovq9AiY5/wMAjh/zU1eisrlCv46ceUoWJUYnj3
5+AuLsg5AKzk7KtrPMAIO4mVGE5S3dM/x7j4ad5M8qnfj1mzrwTUL1fBSz8h
cseUo2cBusD9OG9HbDi7YTzkBxCTC0RPtRb0DcNOON/a0YHzNH04qJijzgya
kNy2Q/E8pEtD3zmVbs5bbiC9kHZNAsGMQZdO10z/fqqJkZnzvzOuyosfhKFT
YWvkmCi3VT9aLMPUxU+Uf2AdX+5Ituo491/Er2OZDUliHM4+fU3OV6q54t5P
W/i9pR9bXB/wBlCphpCmlePP6X6h8WCz9R4coXx+Np/6KONTthfmVO1FLZYR
qkOW1ziIpTi7QSGsCx1cKr/OeorDo3oB7ZbLi3Zcnxcn2kTCW4IO2Un9llNO
9YNkK+l/eK3c3FB8elIjrZT0FeeZz6dJrte5XsKNUyoBpc2vDjBFcoJhhQdx
jJL4P+QolyOuWer7VPoSTHol84wazpXv1m9Gsd7r7lML2qpH3V+StLvJTCWY
+3w4uvvrRXpPsKvVZzizacG7cNgN7paUfCs7Ael6Ix/P28OP3391uvy1f3jv
NyE5x1i2ZfJ4p6z9PUrcUxCBI2+6GJP1DmPgOXBDaLruhRxMgYEH3vG6BvkY
pEtOhUTIxmA4D7uz6NQtKMQVuHwBkI2nsRT3pdVWdRNtS0iTQtnc+z0b23eu
WOu835pP0Z1GtnZTNTn9QxdVjHZLKLY8cuOlIFWsbmFeGsI3xfguPJQxtbrg
rDUu5tvUdLffhMZO8GifU84j2GJger4C5przzK+RDoZdH6zAkVIodtbqNrBq
JHNU7keH2zKrK0hMj30pCLrkAmdgzDF2ir8h+dSrcuqlCaClaI5EGF89+rvi
5NYtyiQ4uve3s+wZiF7L8W5Eia3nkKC0TBtgvdPPysH3rGEU1sTU+2D41q8f
TuKf08t8D7ZjFVut4MP2jLh/w6pGy7kVaaIM9g1I3ScVRdE5sEm8MueYDOQI
sGyQaup1gM4Xr7cIsjsCrOiGCR5XY0Z8kflxJXYc+LBIKTxKzZ3Rqo7NZ1zO
MKdaeZmc+5fxR63cmbRXP7puV4hxl3ubAAKDiso+G8IkQE+SACfWEGXmDxPb
7sNx6s9PohWnCkwdGAx9xz6AL72rUGV1ksgrAuSXqOBEIekeNkAfy68Mj8IQ
4MuNerH6N+jzO+qWejygfSRglxst8Ju+3TEnO1W+zaJduiCRfI54QjUA04MD
UqAVgFzZupuIHYeArCYtErRbieHqNvthS0FbiP2PvgK9MpBuC36foqzWjTdP
hAw5MUQZ6f0KWfuPfPPaycnSlGZy13RNcyGcnRyALVY89oBXuv+Tza20ruZO
JuaTrQsybvBG7nKPWt9SzkqUjmKVATDJMakOu6Azu2Jw3o5yULIMxsOplrc8
eh2mKK9jkVi0Bq65vb85W2n/UMqCTxHFE5eLVxnHRhkppinfsN15IT8Bz/CR
2pWDHmllZZDXGeK31oHSl5ah2JRUKVkjQM979sFh9BZ3Xf58XExmpkXVlV2z
M2TYCaNODsQg9fm8AoCx+rgTd8vGh6aiF6QvitH2lTgAR4M/D/ScYCJFfW22
QnQRty2E4jfuw58J4w1eJ532NTrNxsAuBleejCcTvi0UX19Gb7A/ALtpp/3h
/bDb0vxeJx42VXBgWQUiaKEMJKLOXpS04GJ1GADj6BNGr4VdrVDQlWI5wddx
vOZd0/qtjLG4RxnvKnLfcz0utQm4Y1rxUN89LhaopFf58d+qSlKaVqwJWeHr
yWSObENqFj6PZxvID0gBcqEQ4M24UUDxS64LqRti41KE4jBPKG+rzEeRpiHI
uxTTp9RdLWVN4f6VemshIGTRWe5jUquMNTU5aOe9fQJRoYAAEKGttB9sKI6w
ZE5tiaJVJh/igaa28CSmnnUR528v/qE2qQum1S5P3xKDtma4zF7IC0munT2n
CQs6Ykxucrvw8Hn+NWU4upWiAWzI0o5KwXVK4cl/yyUP1zAaDEewbVs4GrAP
i185ujqhGKhI68jl6R2EzTd4Hhur4YKNdOLA5AhhLs3xLdpZfXv+sUjYIEBN
CnpYUUIf8QFONFcJWh9itlZI6a9vPv2A+VeZPcgVn5vaBjE74lQ+K8Y9ge1/
JC6QsXghQvPXstHjNwv/MUiyLcy+8n4vQr0SWA7V2EZ/OuzR7jTdaryMxf0G
XmhMUYNJ6nm/F5FjnudsILSamHAecXWH0kMoHFtzjzz0LMvFSu7S/tK/A7P4
euLjdDNvoDDY3XeWodAqEXuf4zyDvG4wptB08pgcWryTBPj0NgN+eAli60Mc
DK9eA7j2dFH9r7Q2YKS9kr9d0I8EGh5OoBvZZD4f1hYCcFLCTyN3Oqrs20JJ
GAYGqsXhx0Ujq0rXiTuOO82Nitjun0tizJVm+IDluHa/i6kfRAVosZeN546P
zJ6sv+nGPI77UYf+N8L6oRcGGGExHvFyzTLmZrP4EFQy4D7hSsXKUMDLyVDf
lElIHKoqY3iYHnHetWJ58bwT4/r7Gf1h+OYxHEPEP4KQpy3p1zWpbkqFy6Ia
SMlhCitASeNprTVBGVuO8Q6uCEcONRV8YQlaLugUYKJMIWvxnkrZ06u2+Pqq
6POBpfXXW9TmG3OpsZ9oNEzD8LLUSDwVxTtZMrhWBzXaB4DpgYYMaSKuRysG
iB3I3pN/CRN3tKbjKykWNy7BcIOC5GwklyhcBq2WKOUL0qWgtNKdrGi3YUR7
uMbRTktSMev6HqlMk3ynKn4NosHnlUWwuwJMOwy98O81x3L++W9BPNdIS4hv
582pq0+IeyNrEzSFugSL2MtGGAp5GfyOqDVgUnQTiiKzK5VORwL6jNVjrXB9
Yz7IBtijrHXlQM91w89gsYPxzsDlJwgQhitcMnEQas2PWOhXDrvqaN5Nkg0t
XQ8EvjN/xKVIg2+3CtYra09OHyAkkDnH7+VZmzNuwnDLbXNe4Q9cpR62X+UI
fx7wM+JQ3pUzff/eeQ84ZkWxjCr9Ror+c9latfQpfp5bdMqOEs18u+FBEYFy
ivuMVOHYt3+min1J06SKZMR2N0uv7CBHuYURpVLFHWn7ci2bbKo9qDXe7j3s
emcNtrfFFRjHox70JIrtGUlYcmhvunNvdHJsf6d/nmVs2JhUdirRbxX66lyS
MR1SKh8ZuYfaopwV3XvCrURH43jHH17yA58USd4OuibsW61wxHyUNKjH6Vku
MJRFhnJw/vh3Ryq2c4jfOUlfgUd0hMnwF+SkTIVwpBu169nHG9A5WwSL/nc/
3o4P6ljfO5myFfCE6Y0Rnrs7zZUXzV0SWxZ43GgxQ7b2JRWVEC/mVraBh20Y
vsv3PJT1FWks4tX5RSc2SG+DjTzP7GZItHQ/Ye5NEUA9BKQH8IpdRn3M8isu
LGjT/x/TFB6grqFP231gVsvgQkNfGGa9crdaorLmzlqhD8MaFcYCaauOO0NT
Cs9kbnZMHxdCU9y2QJYOY48gNqKnn9kceyOvnm9IJBsdvLf69HC7OxtagvwL
r+MWaAl+bsEQ23C8hi4tfupJAkodGpLvdmg7XgjbVAt6rry4K4qCPa5Be+mE
NsJNDMukv4Wi9zQpoNz86XOxVKjHE/SN715i72nA2EBEZDdOdZtC+cgInuwa
qBvNilmt+GW7BgG83a3cpdoK1hmxL1JnAxusluQLOX4nuRfCgoQE1Z3eYSmF
WJQx86RZkXn8HZ4HXqs1y+un8hw4ykTv0usQE3Pg010xxTKudJmaTRIwNxA7
O5WC7XgXYRlUvI0m+MqJG2jynU1/vTDE3qNJLI2YkP000LHOGnyVp/6LvI08
iPAqy5OAiu9Q+nexUH50f0Rfxy0E7hKgYOmxEsSaeAXjr03EF4wa7LTV3gGM
uxrU6UbG4bAWnujdePiQMnrAcr0M7N9L+T4/VDgc0/TvupYfb17pVlcqIdql
elYaws8iev+d/HoFxFTFwb8SyXuewYCqmSQ1NrcJAsbmSpVN3cc9ICpNCVxI
M+RfXBYmj9zwCEFM2B972cRW8qBgHYHz0wflycVOHZGSa/lMDR1TAmbJcNXR
uINedXTWYe7NfwNzSiO8yK3503ac6uM4THyELtai35tWJeYqJN0hKEEwQZVy
QUNJJ/rlCZQnYUhcxW3K2FfK/oCWGnv74yaxFFMJaMgoLZfcDBb+TMJ94Hff
+4m3kVEg832E+VDG2PKLuA0TbudqnDWiDFKQbGm9ylET5bs/6GlmRY7cEA9H
OQrsMjVz5GwyX/7E/ZmbiifuiITOGhh/BHHVQ9NSTIqrcB33x/4c+KyDjrB6
ZIJWTH6DZF7IWqmoDMKJvQRYcXhBFLNjuE8NwbOAwIjjyziytaaVogO3wwcd
Aw0cPmQk/5DNAfVnJp6Swr1MR2u/skzb7zsfLNsfedtWd7CDEUQwVcCGjQ71
ksm+0uR+CCvQWq3mMCAeYc8sI4vk5jz7Ssz5QqMfEbm+UcmhXZD1FAqB5IH8
eibI4ZoFxfBdLyHGfBzm3SWiOTqFUFpHPy38CYN6o5GFKS3GfDI3cVAKr/tv
sAMVJTDnl/n0ToIAXlNctb4OAW8V/DUUv4hlUjU1CUVkOviJ9qFxsUaAx6QW
2WMSiQQaemLDADxe/8Z+YQU3ew1+o19ZzUmDRsWtA3SD0ghLhIkyYYFse7yh
mJNilvPDRPHWPfMqUZBny++5nwgE4JICZa5lUyEvSkYmQRWC+XwtQbXzIa4C
2Gqj3uMTKrZxTe4ZD1mcmurm+Nnwn753sSv1ruXkGrcygEjWyueZLYc/5eMN
THXCMm/ZWYFqUun6R4GMVOYw+d8jZ318hLPOLVvz5tqyD6yQYwofJWRXNyYL
GG0hSynZZAF0M0Qp8BrS8vpS/Bcn6dJ8303p+vttp8YI9r6eN/buBPzQka2T
nEOAFa1dkCONQQ6PBsYrjGkv8aFZ6I4/kmGUmSGU8/iT1tmfl+PhYoTEPejg
vvNP5RFpkNHKC3/SnPmC/ZS4pQDVQ4YhTd0ld3vgOkK4YnhwfFDpV9MsG7wF
6FpWAm7BBoK8IuTzfSAYtfdGUNiJD1KU2L8813DFhF3UDqT4a43qyMqdXNeP
oCxWlAiNzBH/2fHeX9J3FXVrkDCUJwgl5mJnJcLhwpKhDRYbzdKuCv7MYMcx
QXmjlk72NsRGd6/sb8kTifDhGUbtLAFs0gzIlYdZTS6T8UoA3iDyBKyilZEK
EHJFWoDxYYXpb4Yq/F98srb8TvAMsWsxB7yveRxW3kv3MNum7kS0bsfslvXh
xJNtnEHNIR1CQwhyUMdD6xhoPnwBBVCCwhe4eUDukXyigL8wvIP05fD1/UGf
aQSolHuzfLa/6eoGd7r6Ywq1y2dIZcx8XM3CV+pmjEciHCcG8YsqNAXx9IJl
K+4dSNQUcSQXj14+9YjIcby4DSdDoOq1uGNOZi6otbJMCMOitkUryTTSHAFG
douX+WHLiLPvU+WhN+lzgf3LP+plvEWr7w6fi9yvgLlG8b9TNFk3pyzbea4Q
kdkinCDCnhYdgJx7PG5wVxgdfgsGdhZaV9eTt5Kmb3Fd/i3RSGL5GXZufCqY
ES8O7JijwFSVuA3j29CUTdiFWsd4BATm1PvodlKyvrmgu2t19Q7SnawyMfRE
FBCL4kDiREGzdx2r6R+oAlGcMfCPMjLN6GhyIxWL7YGvkgHEIfx9BzmLQUVt
NtNMTeLOj1+oyfALNPEcCdiyJdwV7rsrxvQbmtjXHwgEobLwO19wvn1gNq6F
zu5LR1TjGCRiSTCiM/jjLmOnB5aivehr4DrQWFtvDABmaHXFUVWOdgOTELxd
oqfwpyGVh8X0aYPXsNuNwDlooLjoaV+myAolrcWsTvdeHYksjirClbOXwA7h
IUeSubZLBr0I71wAm41JOHvudDfmbqP9pTw+Dlj1u/Ld9RqkyNI+xAtRWKIg
bbkvNBq46tzjvUAwr2e5LfGWkaUIlM/WCooNiM70F/Cwu7Vy+p8+XG61SssL
JCQbmTJ0FuvDbYSLcHfJ+SvDBxn2BxSbDgxGAazboTude34KUyb9Ks4AyS+M
CFwYXzjwb1Ld3qA+EDBNrTG33UIr6iPh6A6JToMUrhcVp10GwDyt8VUZJQgc
Fn05tm9qF3u4lTzjprD+0laoYq+ZNUOaxMm78+eFfpKFA0HtskyZNqfjBynr
bi+TaytUUhFvm/2y0N6ALoASmkw6Ee+Kba4WicrH0R8jMjPzHfOE5NIj+TQY
T+OprE7wehmMukT4mtmVWUWCAwP+BEMu4Kf9dprIUiedh+WcXl3MUb1rcsK9
f0bJT9ueW/Q6YoQgfWoNFDYWlQ+93wrlrHgVpvIzdVMpsfDeiPqZQnnE0ygL
c1ba4jpbh1UslLEtf9Tx0zD7yjZSho2EvJ895EuAzeH70jflPDT88I+D5ate
7joYTr+7fYKREz3XU1BCQ5Ml44seLA12YQYqOGfWsPTsdamw3ftvj6cR7W3Y
3g63ChHDBC8StHezdUEv3Uv0EHxhzwcX31+QnUUJynRJo9heUrl3OFfPWmmJ
ppDnkyVFSQ2Pieb5LV+rVDeuuRqA8d+jF1iaLg6DgDgYJTtZbJwEu6wCEXvM
o8cEDU+lhMWVngy60gXM/zEAVa68fsBVMRPUYI/EVilrpVG/6Mc1YwrXdVMQ
3PH17wAo5rZMhSaXzPyl8mOZ1qlxediJASbhj9tI1ZlPRK+fgY/F/osJvTNp
bweQNI/AQxTrVNPGoQK5Y8356DpxmgKJ/YAF9RECu/KGkCcdXD5+ma+zLnSp
0U/Jmz1CoYUxL+Dz8iD+YY8r8r6CDrGRjnsmRtZjuPrL/sTyynd+61VwEcWr
pEHQQoj5FiQmsKSCJQcyCJMBzHk/pB9KlPGTjGoWr8LSvCXJzDb8jjnl2ynx
MOvTMtv7k5ZXJltVUD18B3bW7vldq8jM9lQ05EMq9AT0nld/qqs4myEmtlBG
cxWie2996L3gCXANzVA54NtxTF/eJdKi+zAQ+/eSTsUAwFIL40pg9tewn+C/
kRscT4tFbEAEeJB51+sCutDTx9FvyPDfw8+wPL0hC1pja2DPymHVkoJZnbTR
jhTzzxU+egwD4PU/L2xFfVF8VJSL50kzJ9e6GP6N4Hq/nwKmpTTBWPtkN8lM
qDgLITIiykKYZ3uGm4e//HJTp9qQ0GSE2dPxvBjCyY6gJl8hdslr9hTf3LYo
dldzBGlscy3ARQ8DTmAztZR0JS14k6Kov4h4ViMBtkIczGclb0u0JTpsdY7L
IZgxfDeLAi0Arf9pA/iCkGqEez+tP5yF2G3luk8OIt+6gPoNggd+hZX2h0ub
HxJM/Fk47x7NldNLeXVs0IwEpNEJHkHVL9pRr5BGTP0WPUdw5clg7pZn1a7O
p+/3ZX0+xMUqve1YPy7wNTbk/rK0qW1xBcD5rbhKEGmm4oKtQ/IpUb7wWmER
Zwuuziq9kFgY0pfh0jXRH3HAz7KjymHIV5oPhSwO3oLDnzeb6vshuvh7qk1M
MNJ93uUH+Y+SxVpz+1VlanjoSJ2WthuCJBAZT5n6Oj7EP5UW1P9ZYcY4thU4
ZxBhIG0Ss8LjmYpTXTdIGoUGpAwXangKBqLxA/GTM2RoKWfyd2pUUrNsnm41
lOrKN9M5s1ZISZ3FX5gQ+gGjmMFJFoM4aYlwkQLkIu4Y6WfFKrwFEypNI0Fb
xZfnTWsuRyyb3prN+OjSKbl8eHWHJTdrrLTUR84kk0XRwWmcK9Lk8WVrjGic
80i2eroq5IADxAkXiEVWGf+LDHR4YxIRMpOKUsLE36LKOizWT2zmOr3jhN8p
JPLIUmWhk3v0ABxht2sxY07m1r/sNgNL/MCaxB3ilagzn+vLaEWNnGmL199v
Q6O8ANbhTGKzzktw3T9shC0GmuOvJHSt96MKJj8MWinhuFlbANI7OKj4NNx7
rcvo47N4W2HfhWbYxrfZECq7BxenF5K7THLG8271gn1EVi+d6z61V/+9SOml
xayG5SazM/WpwXSqcmNp6b7aZ91aZLe1e65uXjceZwMTTGTjn2GJp8sVChyU
mgF+if74JzCiOwUSqQ0pwC7qZB2MEhr9zIV426cL5LHg6Sga7LUPQaOr+brt
kj1gP1l0Oz6R9HKYhgFQR8brvhHMjUXAmhbmDIpr3Kb2QSp1+VEj4+pQQ+nD
UDlORizqLyJBCcQYDJLM7JBv3oPZJoJY/ZM8fGJkYPLgGilbgMknTlN5AGbk
QZSkQ7RjF8rwQpG3pWCTwkkVE6OtC7mac3R0Sp5yAyLZXCPd1dT/hqIvcdz5
RK7snkQA/AVIUiDqgm9ob8Ydgwo5FiqYFo1/F1bSIp4luqE20yyDng1t7a8g
qGzPe29JqogbEaz7SyzSOCmvAQTfAulVAc3NiYqvF5O0tB1mAEQxxNFMa9zn
IZUCkhTbQoCepJ4ewZxIdkRIv9okxhcdsYZ/r6wjdQLUDBqHQtXI8YYhypc3
yqOhAlT/33HMEqouAvd8HbIhOmyshfWmMAI+xlrxWGvElGVORgCo1y7KG+9U
oF0Tq5XK3vCKk2UzWvzLCFzq38IDoj42cu9aL9bIy7gT/RRHuVttu/gQVOL2
OO1OOYcO+HQjNy8mZFXWMCEoUqHwJfsvCSUtgAouTugvycw7Ke2NC6izZS8z
RrCx7bWvWegyKy+Ji7NEWvM4PWnv10Z13x+2QNxZJEBNi3k0PasWuXRfRYCr
TfatJTxtayJOXy8RITHa9ddrJ3Lg9SVp0MWRFmYFJB/VUUFpl8eBoKLNAZWe
rnG32go1mXcI3PeAl5szHWZgZXcmA3X/Ub5saqyWHODt8rggf9jqQnRrKe3Y
AjXWqRSF7+mwYm4NlAQHpWZ2nu3HWeKhNq8QpJiwcdPbUujX8z/0tOac+gAB
pCkdCHEttk1js99zOHBFpLD++xMn5D6b5C0kpPmemt++s2UmX9HBuHdUbM7V
WOArnJ3ODsrmpVpg19tStivqpLV5lw+wmeRzdaAfmnOFr291PB+WHbUbQOlL
SIeyjcUSY9qiGeZjt7aPN5Roq2TV3qj1Lhgmj/zKAOy9ZigDNkDv4t8t4QLZ
oxlta9kj8pOfcqztSQmbsk/Gr6A4hhCVU+vg4C+03SR3VyxSuZj/0qiKZWVK
XPKP+iasDBdWeKaeAGOVKEFc3RI20MWOETa5df2tSr7V51u9jFr4GxSFsS6n
NRJ4N/YpNnMVkEgM8483B5QUVYOQZIwX99+ihU3LcDyimi/voq2ZGgaYXxmd
NgoyjrHPCMPBpPyy56Uh5SHp1WOgYocqQ2vTSYj3NuMWg49BOEM2PZyAuPG8
5iXeA7PBzowAQf3YSS2pH6VFYR8EbTRTabJgueosxAKPEmQbb6BiZEETZUSY
CyvlDsB3W3+oFOaFvLJmkH8xWKovtLzaZ1pIvnpyyNfcFUkX2EL9oWkW/mUb
Mclss6CR64LIs4TID02gEi0Ot7xe+h0zHdOnEsoM6DOCokZgxBZrA5yy4ZyW
anxD/eib8xH2b9eOMilLONgQSboRLYrvStI0/WQQ4+lEmy+BNaUBEO26mxgB
BeZ+/I8wFKp/+4b+94fNVsrVbdOL50hMBqE2ypm54RVhj5d+rT1Uv9wuiUaw
feIzoOClAV2wNTyqyiCcasz46fo0x1pTMf/KKfJ1h79AGiToQ4gmO8OE4lmo
mAS8kE9rqV2SKEGx3oTW4yTiVtyvkh4vCmFQHtKVjsxnK1Jl9p8cWDImN3rF
l4PmBcfts6RX5sT8GhHFegspQa2falxVJYYeBs6IdJUSz9EPayLIpzx4YBSA
51sG9c+rJ7ITTMcxaDm+641vy5ZCffJVw2HC/h36CSxA4sNkNNni09vJXp6A
tsFGcl3UTGPG+WSa6MCycl9MMJb0S7EISa8cYp9bZ6etaqI/CVKfK+1zW6m3
/tu3h7yvD8lLfpPGulHkvPhuB0/Y/KVqD4fjdoJbErn41FJsKmbJXO9sA1DV
2M1FNDf6LHQICPo8YvCftqiVBml5lSZR0f2S7DluVUXall5/QYzbF98XxT1W
Mk9GgM6qplNOqbIZcXAenlWwXBbJMRTf2Nsh/yr7wtPzkpKPcou/vCiIwCht
LdX23fgvCFGxQSOjT0b5y3sbUigrjCNEjFSw/EWBR5N1TLZjU+G/BMDY/dr2
G3xFJDf0r7ZJSc9kb4KeSn22y9Prn1Q3D+OsojeIhWvd+qdphzAMDJtCuHqv
m+bYJ/7K8XNPKxaf7rbXFZ1pl0W4wA8T7gLxTt+yIBYWYZSy1U71XWgckPWa
Px4jwGXrthU7/azbuGiX5cAHrR1b/SoW9+N0ZJg838TKQeTVXKL52mqf+yCa
gXin7E5x+eUXMeAG90T25xVg6UDho2JLds73e6czNuN9o4uUbIojbLTMRkHs
Axoh/lOMaYbqVvZHSaOrBEWPtLoPL5KFkgNtCM0VhLYncXT5iyxwTGf/a9cx
ZUQzOElkXz5Ok956efnwmcd6Yf3b3U23w49ZIvh63Cte4TCiQZwhaFKTHQqt
gV5qLcF4ader55ggTVkLFKnzztil32xXE+9GGfmeZRF4GbJY0Skh6bLlS6T/
xMvbQztVoR40aIQ3EeMm1pkinxTI09ndUEM5c4n0rrrC2oz57gmdcauimZmm
N9Tb0f72vfggmJ5wl8qLokbZr/nK+HIFFouV1XTgIk6U8nzo5vTl1zQJOupI
KYMNINYEZEqAissPFm+1w9LmXRDcxiyVTWBmLPfckqxyGN6I/PPAUtuFzeV0
WYjQahJuu0ZKIrpJFRuy1IieAeJK1Zd/5nvWqYuK6Nkj9kbDd3Q6RVpOl4o+
gXmgZy0xHcIgPEInrIIhBUDYQ8AbN6Ga4pR/qvQiCOk1VyJnjRXCNFO40WjG
0FGhY3UoubZRPrQhY5B3g6AINKUOUl97K2XnByChRS1ANB1Xdein5ueCJVMU
kEwWC/aFcgE+y24jHneO97yiGhKJm254rwbgD9MNzltYwO7tF11Oh8spfyY3
bbwa9ebtBjYCFNArA5PzdW7A/oQ6AGx/oeggu3A8GPQGJneqcHsqROcGpCOI
iuZIlh4WxixsEHX227Amkhe68KrSTNwFCK3gK+O9hu0Xl6QICeGml793G6HH
xR6eSFjE5wQs7x3wXq1baMHhG8xkq/vflbYRpbSt0JCkhZo1G/HSZYC7RnLi
FPCGHxrGqiCKmHUupWgN8fCmZoowW3FJb+kNIwaszUyovH82xm/BU1/ZW8ct
LaDZjkUCPR67twI/YZgpqclheDA0JtetS9ZiP5/F+Azg5sLxmAvR4CEQb++a
JVJHENaPWfpTGHMejrMd4oYm//9rBxwmWaI90lnRKup7jBsaf7NabY9M2K27
VgP7YfcQ32HHU9fdryzuBvw/rcDVFAVfWml/+qcX77f4DMF/W9dp86uxMjbH
o33g8ogxt1cUwAqIdhenbu3oq5wfWI27vTH3PlPanCPaWym9O1p4W8edWpDR
t7//LL+thJoEWSI62mTgPxKbUMEHXJKUIChXpstgQQgpgmPJB0KGGy677zY4
zF7eBazwC6iRa/mUF8HtuAFJYu1T74f8N3HG8/nW8qXNQ4cUlUHW6XWN6fFc
4Rm5eyKXbhlkBxaTyrCElaKoZIAbwfg7aZQm3V0wn3G5gAryvwONbcZCoca7
s+t5YZ9UVDsKdWWRJqXj5ds57/gc6R1o+cHDMWDkYyxTTBRXFaEK3NMxUhDI
CNsj+/v+UJB0k6/E+U7SklQ4v8P4klcOmYi2hw2Qy8QcYhuYn47hGroQD/vn
o0HJHfkOoajcyDpPZmJ5epG+x3ax5DUUiIyDtWF5EHr8TSyzmOqn+ShszZOs
Xnq2dm1VFMlu3ugPwq7W+a0PAPseq3s5y313mrNdDJ5uVqhde5KsZz0lhSZ9
tHdrStml+IAYKwWk9oz5mA6NmaL8amwIt4J5dcmN6rlKSjye0+ES9k17f8o9
JKqCHQk74SRPx0E29OzHnNyGznqJMsXMB5Aufje4BwBJteXal886e927hJ8R
ZuPwwLROqx74Fl1YxAj8jGORwk9Ps662z6mCe8kcL3j7J6zc7w6hTqLKXm1t
6vU67CM7xOYSbA0ZGsHs6jlUv+orizA8nUGqAnixySodKsltEtFTxmKfOMfs
7DiVOjR0yA26MX1xxWbjO2m8xNKkw1P2aV2FUBAL3RA/4ARwZSxsbQP52sRR
LlzSeERrPP3Jn3r1xOeoM6tXl1WINREqbzmFip0vVkRzB/CDBkJh5RLXWRAp
UNRsmVAzpbqRzPi8QN/6ShEvvfJJ/0HHcl9D9wa132iuGWb8LFu1jV3r+ysc
aoSMEEOgN0FG/58WgRD51FJ/Ym9nXqEsv9Km4V/U3lBkgrdvAuMrAnyYmdvb
4jD4QIZbVG2Wl1zi/MszWzkSjQvs7xEv8GoBhQ4Ph5o1XKrpSyeN9TUD3vu6
1AsQKyffneeytsKfax2w+gBthBtsk6xa+xKIkgAM6HtnhsE7TpyH0zvrVAv5
U17+xDl2aDHRRh0tvZccSn2BWJegoHi7a0A5YmztoBpKi9lYQOf3T63FZji1
5vv9SvmjdUY8wavudSkH2SWR8i/WFqctDJRM6mbKwZ0aED3ordYVFKHaJMEL
wmEItf2y3JoPu8put3CXw8rhDpOBr6AGK6CUyoc6MzLqnNPQI0NDL/5uJC59
aIs6n5qg7X5f5sEjyHOLjsh+gPo5f7zn2GRcDBU5jTLQ/5EeO1X/jAURrKSW
z6dz0pq6UeumbW9ArV8eAvkctENUzuOqwm3OEHFGTgAYwlhZ3X8ZfNt2tQ+3
vVn3L/Yxg3aH2dXcb9Gg5SS3DRums4f8VJaYkXKc/HQwIwXmDnYVQbMBb0hj
VgzqR0v/R21GLNIsoTNQ4va7UeAKqp2W8+ZgWW/FCkDmVIKK8GwspFArhs7w
jMqR5XAD6PxmFn/91dWv6xUwfnmLe0jjLEsRNjWcwvSUDicjEdHK1MIPtSmz
twoTwMLWnDKv0mrhkAemBmZnKtKO+Jg4mN3OIL/Pl6LH2ulcObK7/ktOP+Nj
tXGGJ9LC0TzCBDt/HxnUuYJtWYv5pl9yhKadnahPcku+naQjC8jWKqoxSR0y
BtexvQly6syhO/ss2FOHkRT+e6XmtBWLHqPtKuCv1rvACn1SKmzQ9tGzGuf7
Z0rUWLNgvOi6esHQb1QVJyrbTpPl37yNe03lJpzLlyl3mZA/lcJlQImOhZjt
YjLgl2VfNLMfqSaYN0v4X2OuETGmI93Dcc2hfKt0BvxblAw0GsV8m6h2dbV8
trLX6e44V/ZdqEQ+schE1zhIpECmj7gYrD/DNEQwn7wlrLrFsUiHHTZDZsMw
7DDVwBKuYNvMwb9rgufSFD5zmyWzQLuhaIuI/6fJO+pAcJnf7bS7kdO2lqQC
78YXVvW1b/7slcD+d2R7eqTp4iMrcGs4hd6yP0pFaBya9VF1rJyuSil789i5
a1ILtzvjP8EyPCE63VYjLZBY+8ukcW27jqwB80FxXRk9jUBsD776vrQ65JK5
ARe2aXSBT2AL/J3mhsc+6y5p3PzSJ3t7P/NFDPar/K8sVRSr0MnYPGN9/RSO
0DOh8aVEW/CwnTgAJiSaVrlo/EPzJGEB6yJtQWixENG1Qj62bBYsWtpljpal
QeueRWI0glswXMQJBw7BoygfOSnL51IXquU2wUzhYb/1ctVmprnxj9ycaRg0
XgDPHnX+hSHW8Qq7c6kSrqGV1136jxdj1OCoAbwFNlRylXxudY943O1X/Pob
X3zhR3jgXt/4IRj9KbbpOvtkRefJLMkvRncFan/xcWkK6v3gX1UvwsBeVnay
jxedZPA0/k73xsLUMbwFXMf4J3C/oSd9RQtbfzvwBOzhAo4pbVMWT+YLirlt
8aJw0lNfpNPCJtyT3A9XUb6q8iGvJhSJ+C7OqmjdZ6GmasHK55yDN1791tr+
xQUQH0jVb46OTpm+ksaYAbYzpIyj+lSjS3V6dSwbODDPFErAfEzNrn5ldtJ5
KJSOwJTlAwlOO3SQM7niLwYiHhqe1FabQCGfetwh/JX54vOG9MW3B2Ku6mjm
POc9FMUoaT9wOCiSXin04rDjQ+yXonPnQqSAxImeeME+ACtAyzvW2Y4yRucb
ol3CoXmymjLnyFksi0wxF21kwDpQR5ZMzXi+qMziJCLm3TFu8E9b40X4RRjk
CkTGl+tyj+/TOp1KCBoIJm9dWjxpMwZllF2F3vPhBTI+mLc24kGvG/KqeMYS
83V54EhkuNgpqKNN7xqPua7rkI7ocTl5ynBSwpebIFze2uojSEHb8DGp9v1y
k9wHxbxTbBcWxEgIUgjfZozITatzG0kIoVoWHvy2pYOghGohnlWBflNLg9jl
2dwlNzgDmJyo1wDNNUCPwhUaXo1MgcofyOXYC7ixExC+GCGZfSAHA9m6q8gs
4q9JFuI1Er3mVo0V1+EtlP8deQHlh5NNj6bKxXT0ubbE4/DB6t3vDUO8tnNk
mZY/RIwos+zg3env6RD86yBNX+TqyvifGggW2eOWiSEOHEN7/FyTJ28TwJi3
dYhScORhL2yD//AwxsSQ4meufJiP/i67EUdQO188LicmGaRf+cz9Poa1Ql/J
YyMKsl3BPKeFHxhi2EWK6yWpdNJKR/NNMqFWIprAT/1WcbU0WARstRuxK3vk
CcK5TeXJ2hsJtsjFpo32mz2T6nq2376hcOUvxwflQVQSx41BpQv+r2laAlq3
uV7TS87pGuMrmVWKH37RehOeZPuG3lAb0CVlJTHigk2o+1WV7ulW3bn/xjcy
7rSChiEJFjtlKm0yXLebB43wR5edonXf/O34UvBzaV1odsjIVWgszymNb2te
MkJQ9vzprUGtFwXuSbHfC9LAL90AotntD7XwlAv8pxvjVYtM9618uhcmw8ab
FKX80BfRAVIgcHQWt8V4u0jq6vYrAfoFBYpwmPNZBCNDQTD5QT4TAdTJt++F
9v48a9UTxi0lzdA7GaRVgkSjAtVOFPNQsz/W2ttmTNNuRBBn4VErfnceOXGA
TFayPbDisOAxEYLeb97r8QM1MDyv9Zp2V853kbymxxBTEbV92U2JHTADbTCk
RQk+ekQSWBJnjjkIoyrpTJe6Qbeb8uQqO9Ae5SikFnXYzilan22Sbj+sF2K3
Xvyu9w0ozdUos3UQueKskoxztghnPxdxxUaZHMXzTRajYIJv7quammlrynks
XbtH47bVHGA3aEryaXYhzvc6pMkZeYJAubwI3lc0pQdC6Gam+NvrY9wa7R3A
y7SqMTq6DrTe0GPMWcUgv21a1VkZ7bEn80tHmO3BLp3uFnvswf1gy7YHder4
WCdOred2ZLfJIVO4TH/GFmJKpciGup4uqmdr9/rcrZq2N8Az0t93sv8xqkq/
bxTQBkRLTMUOziSAtobJH0vNIKU3l23fTDWq2s2/kT4U/wCJj8reQJwdiJtz
G3M1ctfduj1RZHraCKP3uQJ3DuBcLsnWqiYgQYIkW8RFxl9pZaCzKgwbTzoj
MXLCJGqxnnncoJd2Cwqw5tLfQZlX3wj40IXVMDckK47XD55QmrVk89UgBZKI
VTmdfbEte11RwxKsgu6hKi23uVgKXvVWOJIVAxwou3fdUQ8HItou10z2FcWR
FsTaoUT14LlBFY97391c+2vD69tylJJzdE9Rn8U0Rig3BmMeYirn9jtWNprE
NUf3efWKQmeyevqoUnzhla87CAUcnYYgzvKBVmOo4fkTGLEk9eFvydTkeJtq
9w7LPCBDcMd7nmxEqBAWFsb74eZwTN3IaA0s/ilAOvJEkE/gkFoJZoHXdAa/
DI4nZTnAtkK3LxfBSs7bsJAdUoNPngWGwUAEYSEs2yDC7wpAThGZhsUtMDh5
UP2cOA/gRr9xL3p8qEB21tIyS7dZVfhAZknVlB7dADvbK11rr/n8xCsndNRF
Xv2fiRgc9xbBrfGhce3DGZPax/S4BzKzeoDiPvloh15xxerT2zZzE1AcCaOM
sX4MyBXtFzceVPO3EuyoSGoFnJaFLPAoTxyHbq+MB341xqDqGnx20b26ggtT
8Wj6oBZ1inMbi5teKkuCLVar4XUafo+uIGOkGaJ7GPK8CymAmNhsyeXoL4FV
fE0MK3VtWqncPcdcsMLFpw1SqDLDLdYyQ+dptpC++ey2GqZhemElNyQ3XPeF
PRISiGuNkF4KfdpWbaeDRLCHNY44Cc0Du4W31HTk3kP3q1NvmC0d8DhPFRnl
GjvhegXs81dqV0ZIayoir+0d6SuJZt1J/eCdK0gwTjT5kxvKmO1BN8Y1zBfl
vH5rNevbrKJWbqYz1I2BGg+zqvGXMlO4B+Jrg4FwOFdkkRJe00YfXXO1/t71
TY7qfno/Ro9d5zVHs4uzZ+0sZ7WzxFeESDPMBXUsozQ/4D0MZkFoBxtC42Ks
WyQSMUzKAKWUasTXZ3u2NI/9i0jUe3ssa+W5o28QRnz31WdeFHTca1qcBISZ
YiLW1qWiGXQXvnSYXZZB0YhocAwhQN/z49re8tCuzb4yHavWztOwNFRnFwct
23crhAAVY3W7rXv7NVzsWtE7cxROY8YQl5+57Qoh9Q5lsBQDQz4q0Q64lXO5
HF9XolTEdjVj3cEUmBbWhh7KQ4mbm5kLGbmpCFgIxxLXRnRnObzqx7h+FOzc
vK7Y515MMT1I0rJBQgTWxXJebBOH8FWTb9lf8FSDHt5TLHbY86CuLnC1V26z
Z6zWyLt26ZTv2tXifxsBqeZs4dQ0aA8qsl5D65SJzdMH8MsLOsiHaX0cRF9A
z/mS1BIf68uGJQ+n2CZTV3U6bqa8lz8MPpRPckOeGwWNyBE147IzT3LBraHL
VnHtBXAczaPh1Juay88G7b8jJNH0WkBKK6jjq2jTsx+nZb1gRuw7uo+/0OxI
wQw9dIOuGmWGwTCVTqFsQ6pxTMUp3FzSkTxLv6YB7UbuoE3wal+5tlWq/Qa/
ZcvMvHiQzoEJcmRIE7NeuLF31+LrMF/aaiBMKWEN6glLrEoyFby/qnf9p2TQ
LM/2C6be8MdmlpYA/FZmvwhRT5aMxNrqL8RZc9qWADrM6YNP7GCs8zCk6hma
0KFyUS+ixtF4LiB7q7kgTD0MgbV/MVFSGAWGn+lHkVkFasK1/YaDiIlwhzyF
Tfw69TU7YXB28VIVQ8Tz+yPnYriATb78cmdIr47LWMJlT/fUNvyf2qljs9eU
2EXb9i+STPgzFumeDl7SBOCx+/wdO0myUciIXS7mHDcv5CN3ee5K7s+7jC3U
rmanvXCnsXHk9cWFRqlf51/wn4bsntbeBQn1Pa0mhxfGSDah2PLnleL8au0x
lSq79FvINRTc5ppvEVr+PmzcJPzLO2t7VLPnMfkL78HOucNc45Qai8ytohsO
gQ0TcaDEmbm44Ad/t+NqF2YsJo1subbxsmtAyGlxb6deFLsK75HU3MQgIl5F
4wlCwVGcUnB8Kv4D9w82emyqCdGrksFaolb8oUu5FlZft6t0vmvM/Do0aomR
xhGCYwVog744TKaa5as2EEM1arH42Dx6qmKQ0oCbjGJjIohCBHCggz52BkIa
jjzwUj8fkJgqZX7ZkVJrXQDH9rjxwkifKlYl2+5ILztpgMMLDE3K18m3RoYO
AhVg3NKrVybZ9errHGM/OkozZgVyRcdISJSemCuwaXgyQE5IGsdEFAoBhEx9
JdeIz3XmHbEcnczW1TYHO9YDeIjd9oSl9FELb0JSaHZZPp3hWkUgtPuYKBIA
VH+eEKejbtGFVws0osiXRDrwhoAh5RcESubKmU8ICNURF1pdhb28Wkua0+Pa
n/1UxASKGXwOcMAltGL+jSO3Bgd+659TN4dSHB4t3Hs6NOdPGU7/G0DVSoL+
WjJtPGU158UtRxa8bBGe8lsNdLCrDoXFQyUTGswU2VZawihrOYKSN5a9RDFG
qm566oluMKaeLYvOo1HffaprsXp0qdPxFU3HJlpoKDY0ZLNS0mHt/zVrSv8H
Kt2x6aLdMwAJrfKmYezeGqfLaSXpMo472XAB9DWMhVqR/LzMW1ilrBiCzovp
5+Mku9lAADneouP0rG2ZbN+KFG57DZmSn/7XlQHaXOrlUwkXPQHMwa6YZ7IZ
RHgCKlX/j7dOTEVS2JzZLJRa83uv83wUA3pDfUpQLs2ZCzMXWkXgt2ai6WX2
Y5VVKv6heq8GNHsRqBjwQVATD/iVd8Rz/HKhYze6VU6lep4fMpGd19YAf7bs
Nj4Kboc9RODXPqib6uV0UcHy0U9YaIyHPmrCXQqcWCX/cHs6IXA93mJzNxav
RuBtTzDF7nDxeCoTPzqBn8Eatw7JSQN4LbZXOjyDbopIX16XUm0orp3svabt
WIej840z7FIgsJ3/TsHv/h2hqQ3CJWLDsYnV50FDZ+YnMFpHuBCzG7PhecYY
OF/tdciLhUYshH/tQB2q9o73Cuk6WolTA4SjslcIM2/WirxuXd3SqMnf29ca
bJIynb3YCpOQiLxltSd3yARNEtuGY0Pl6UjDqdTaU7z+gPijjnIEsxunt/ZW
5qZxly5ce8GJUgwUMlNHwyAhJcoR5s3QlYUl1rKrKovLJYhrWrmlYAahiQqR
yRy4sdZ7m8q3yM8rqkl8upmrnPQYYeP6cE5yvyHaBTOr1EgUm+SnG6zGzZou
syQMgxdkthDaJ0qhHNNhJoLtunXqiqZX+sLEma9iyBgUcD/zyXZYQAdxvyKj
iJm1+QTryWGbXBI0cUaQLrOxel6W+ME26EpNTTRwV/SahANXVuqS1GUOj0uD
6TxrRTKoQRMMHLSl+VqW3IKnobDyRUdR8HFBwg9IqkKFbvvm+nmR5zU6U9ZG
f9LQenwMUuUnAdvt5RDYFR346bwHf9tdk/N8yKY66Jzx9OZ3E17glzHZluZ8
rrLj//Dj5d0Z1r7bPnlMUXOBjW+NQt6CEVGycN+OBlAFiAPm0FTtPD6y7qWt
Y9FiJLUa/Jzm2UFYnUk2I0/pzoJ9u9HIHxwxGB4yIjFOAdcoIZTv/WOcFpaj
MpsiHxyCvfPjSC4iuKyfRMRJx3CQtjZZG1BA7lsz3xmWtUhKkL7KkNhC+//A
VFWJRCpyw4+79RO6p3O7D8NSpoQmuaI677JBXRGxU6LbjM07z/HQOjT6rGYV
AWEzSMQxDaCaFWUUz+BEGdpNWBKpml7ph3WP6SlmWvYPmTHEBtNhNUFzKqDw
w0kSZWhHkE/wx0rlSO4IZA1IlcqjBKOBXGkqAs9SuInnCCs4CGbpQXp4ehFj
qYPoCnjVISWWiX/k17izZonbP7x1yp14cRgsPZTTIxzAv4WIFY3UOKCxvSDE
FHU9eM3Nbmdx+dgfz4zfPDszlNb4smAa/kpz3ZhNYGhBeXsJwDwgRoa++Pxk
0I66LTZUyBXY4xd6kNNHlF+1/9S43eE+W1sECac1XR3DZ/qRi/HCWosNFJYM
HPgvV6Ru4VJXN/EueTcE1NRvEMgYinifTTPT3ei0AMngqy1UulY5JxAUkP7Y
KIGz6vFealPnY3zDyL9tmHMkeDVqMGIRfYox2BNfDseWu08knsYoqd89TIaS
V6cAhfswQxSGoidPvKvfhE3dzurwNRtOFp2yiSx857tsY1ZtKV5cIo+5MyGk
0JW6sdr1D81IcrQ7dS6f8Tmp3lFsRwP12YaF3VdhndbYXGFmaLXKe6nu5Uud
lv/II/5aAVrWdUUQUfU22eXMo0GDxHgBU5HHnIJ93nqd+FUtitioNuR9Ehd2
n33JC4Xs9uyiLBB1xTHREAj11Nk8jyuFsO8qcI8k0oMsco3w2DNt3kwDt9MS
QsH9YbJLdIEEXHwkt++FhIJ9AdE2Xh50f9M9w89952ux3cDWZMckPrZ5Cyyv
2rfKJBgcdnSb2SYwdPFHoTAGE30lBjvZKiq/aY82RsxEacWNX48PDZd6nvQQ
KQr5dK95sOTW0mR6aU3qSLp8otBgXfHMK3yY5o6/x9GAI+XqxoR9tvbQMv+G
0vosyDKZ/kQpohdSUNXZUtVwd13acz46iTW12j85nwniCIkZw7XvN4LSFeMq
5Xqs8FAHduxnRNSBbT7BGo41GLqItr4yxwIVjc+V1+JbeWormLcKurWQtEQV
lMIAUzm5LU7mVdPjOjqu6eUUStvRCyEp1WBWBldPJ4Z6YGxMtXyuDd5cgbED
fTIB6ZBZCMWNjYwUxS/AY32LOZ+z6tYw8UCalmlofGQAR4v1hi74htvozxkX
FuOSX7Ioykt/ja5AjaJaDnLM0WDHTgNlKfoV5apq42eRL9eIa4cEHVjaiZj8
sgHPzb43ChXfE2YW9QugmDlyupmraOBre9ZiamOU+BEvg6wFBXGH4/7yW1yc
KpDTaRyc54KlaoBrKzT2j5olyV2Gh0qvXxBS3WuVdSeKkAMWaz5sM/1JFL0f
9qtOdA6X9D9EBN+ZvcrEY/HXPE38ZUWmZzqDtDmDqBxKrF9fAkNL1kQzKHIB
aFRj8IINz3Y881auslnoE/gMAh0+KyCvNPJ9vsLB4OssstOpPpRlB4VGU6SF
9I30gzoJRUp6gYjU8H2N1oBXVbnyR5oWnaOVyH2jg+O5Fnfpa8x3UWM/KlrY
BAxwhkKA4979c1hk02s3C2Eupx1eA35pPWjlS8stTy7qOWxzvQw8U1dkKjOu
9ky5zT/Kkl19xd5+ezQ7KM/bjtFljL0m458HFy/aYBH6LPmHug5RQPtsuS13
b/X0q+AeL6mT/t+wAEvmC2AhmHhIDQ24fCAcZEBQ9S+7wzlsdDnlE2lYxfbr
KftyhbTJ8NQtiabYo3AudSchSM+JieYdfQUYknO2gP3JIUG4pfspVdydvj30
Rus5OlAk4BdFnJk2TLNTCUcgFXnUXbcfFMGzF3qfilgQj70R+aPQuNiXtRFn
IIbH+PaN2AF6ymk0PBN/Qn+KWXAEUoVcZt8YKSlfztc6hLQOH3EVEL98KKLb
YlN87YxN4pZW4bQjJSnG0S2Bo64llovoayr6oxLLUu4Owldc06nGDliD1wlZ
hMU0IwfHZGIgYQ7HtX64w85dqDyjqB0Biku7TFg/qDhqLfAwLcPgLIACP9kq
Oa/Vr317i0sDNg1hEyOkVXdH6wfqoVcbfYkTRtZmKECbzTt49BvLCVqlX1XF
xDmBdEKbiigPaWFPD4u0d93TKrNR5Anrj+YSRg+ObfSQ3s2PRNeZsZQdoB0c
kdHWWPSwsH/BzMIiSvNgrT2hPtyCAwPMAYaJNVR8l7BavQuGUZMfPeXZlM1U
V28QKAviNe9i8wqk9NBagpyw5cFcNuQKTiMhq/sgN8PCV03LjJpLzLG+po82
b6xQw8qUOoBabh3TBJn5NJisq1/Oo9gkxRurFIpkebX2uFQe2/VWOQD5FZIZ
q/NIckEMDx1c/OCPp6CCCmInr+GrUS79njjVm1loHu76DQ0TMNi+WXJaT9hv
xgvACLr/OVdUnEuPwCFGOd5/bKQpKIago/qnYSI2N3LpKCjF6U7pszlc1+2A
dmWcIW9DM8HsJ5+R/81swlX2jaXN+t+/TRpltkAcGJzWAvhBpfIbpD3s7t6J
yzLThkfdZubpJwxo8C4geyxnh4rhefHNsJZTfXU/fKS24Z5A8cDOrlUmSLwo
EnDBP/gBr5aw5M0ghmU5z5D/wcvstVqd/7PY9urMZ1fj3Fb+lWrawL9OIjYE
Hh1Kgel+DhhFwQMbaJFLof/71lEmN2e+T5aBQoxIEPTxQtf4XPwproEnkVkE
dcBELy1T/yKs0bJzCZerwEbfqQF3hOgAKl/L68Ugw7Z/WxbmyqRAEiV2E6Yh
2JQqkmvwAk2PXGYpryy7hERw83+rNtOTrY4YjR0U+vCCaCcPohHFbJTBMDWI
+CDLS7RAdLdBr199Ji50jYwap1vDu8BIk65P0uSrQ7dmOeugNMFHwVMGpsHP
SYLQVH4vHBzvFQkFKFPhHpw3ectTT9/XPw2hdAkww10ktkHrVNavkvwH4uEu
aq2ZSsXOlbw7Lo8NKQfr9i9c3W0U+OBmhN0zbX4gFPiqi3pUkvvuK4dNWFyy
MlHRvjAUSOEmx8zmt2/Tvbt17H4ZYtj/HlhV4tDk66ej2bXJE2p7+u81OvLh
frao+pWAJfTnQFcq67Z0HBnTjZZdII8zzr0vT5JOKgIXuKO1smBGzj8Xumd7
BWu+iTKPvkNRhM/EzQcmdxbEGxN+uBwnPxD+f5kolszQ5uNohjXn1+pmdc88
oAWg9Hhp7YsOQxCDrChqot6T3MWTuwNKzy1304aVSfjsAUQ1x8XgF6K0iNJ4
AyOXvGJ34rBq2NPp6ioyW+ypZMXdIjICuEIJmooBQguTOP2RdcqysYQqFWiY
+jzWNiMEt65wodimaqqpfP3Nmaknt3X4ys83/X4trg1fzdsnWf8HbEXwqcza
t/jL6TrmM+5Vghp29uujCzVkKsOuRPHFx/UAjvTTAwIOFIwg5cOQtWaHqE/w
A+/Y4yTVkhyW+q5QHYKb4N5Q/NiFFIwio/pBQ7r1D1JkjOjB81thctYKJwMb
TodMevlqpEc6w2duK6pz+1P45463Z7yLfTkZjtSqyZ+4ktnVX3z4fh3ucw69
bH2ATfSlvc0ac4yKm1QXlW5Z/vHL3LHC7/dxbV5OSiothU/FxNC4FW10RiMF
RH0vTVYozAHXb2P24ab3oqstpdrhPfwNNJvLktpXWIM8hFJwCdCb7+XRO36b
ji+ka0++gkLMZ5Ofa1shlCIPhiFv14CH1j/KkBieabNgMzMUpGSMRi+vW93P
lqOCWF6C+CGlw7anbI1LcBoXQONL0JKPH/49hG/nkSQgsgDDoJrGuPTGHjV2
/8X34c/2RlPSffwp7OA8GAsh1sLUukX9PRZkx/rr1R02o2CJmhSwkSU6Ml6x
/wrd87Sbhj2TkKdNfzJceHN5F4K1ZSw2N7WYndS8csuWMGCd6EvIt00K1wIM
VHTsvupJ38fNv9RdWlsF2Nmyw+pclTiX79qZKIiWO2L+gTLlSYBPKZ2vdcjP
6AdDt9K/exQ+7omJK4j7BvXOfhcoeig8IQA1/xDIf2OFrNqUG6e4fD2b0ESh
5ZEFn8aTM4L1S8saxcZ/BLxbZhxyni0Mu1R+YhR0eNUvmiJiVhZgZl+S9Kz5
7tntIu85cW3y6larziyghvUFxZlgVSYQxiRGHFfy4G62Je2G0ZJJpHm15LNk
tm0Jr3x/Q/yK/rVINhaBZCaCtMFmVXg5ZNV8BaKGYjc4DUL72E+KfBqUmLDM
nW74MAAjpzucXO9+XS+nEhiBkcajm5WkyFoM9uUd5vw8epBKdjGvXdLUkXSw
ovSVIHg0Db+vjzLlWAmK0m6/Kc4SW+HSqZiudKx9jtuvArK+3Oh2v/N+3t8H
PTEGPHXLdGY6IKNZFg7vNG9VSPlrDCQGt6hDsaufdjhQchqlhr/pLfmOW/jt
alMU1cGW467bg9ib3i8gMaqOx7EIVxCh71UOfqGfgYVUgZASQvcwx5J84cW5
YakFvyiCk8blInBo2/zDAF81bEYu2Fz9o3LWui9nTQZYvr3PR/7zSur6dz6C
m3BhymTRBUaEXHhLhbb7B3FVvWq4w0X5S0Qhxx5FGa2qlA2Eq53YaPGudTtx
pyXGHlLieQ89w0mxsU8I5sQWuWr25DyWA9qcyoKMEc6nnOmBRTDpaybr7wF/
q5le3NbyqTGIGA2lCHpwRsNd4TpjxssXZxjbqAyxaSXOg3O4+TdKgcjycUtU
iavQP3A69OB+NgcMmpLRvDrHxGejTRi8yV1EARAkvSbid0mp3Gxt3BTTR8dD
1nM6ZzGiEqt93Ti5AvIWP8VmDIlPE+Tcm+0MmK78FIMHdWZSKQvEJ46BQTK2
oA07vNH58vBbmX9BYqQuvyrphz5kHEB5NCFmfOcj2du6wFMJdiGSqMAk1JZe
RoKuerDght/ifPjhbEcuZu9PMxNikIY3Jmr5dKet2Kow78UV8xwp8b0T5VlO
E7ofTQ1ViMF8i4SHGAT8X6T7yEq4/SIYqiAFz26AII2j2W3uFZ9rCkaAOC+2
BbjPSX02tZVB24XN5ngpDm8P1cdIzJj48BgVAPjL17CbR9pt64f45mg8y/aM
jJtkm1A8rHeqcxvjykG+MrU8NgzSl1mIfJQ/zLcnddEu5jUuQGXT8TL1toNV
4vbA6YpMnhaGCoVkeNdHKEavc19AKVHrhzL1Ew642M/Jw8IMr6HLM00pkWMV
8lrfi0fPmyTrd9WStVP0ZgpBrrTgYwoc5FfLxRSFKhkOdpI2FEDKsdysJ1SN
U73E+Z5z/FhKnXUVpeTfjqQzERk2B7iaBWY0aGBW2rkQNgHZqIjERnwGWA1P
QSnesRb3Fp2Pw9YfJv31UX3x1VMTxdWPQKjpm3ieZfPKJKwUv2AU3lZEmTHH
MwuUvxy4i7FaQtIKAroNDeenGRjSYSHTJJHLqBjLkpWhIoOlMwxEnD6fIiik
HoiNpy6GhBVO6rhcyp+m5dEHFots4NpALFQedd1povyn0tXXuri2wXJcwgyx
nXIijDLpvsSS+16hlUCagUkLsB5myM7Pj9FX9ros5MT2i8b5SyiS583/ROyX
KO78EEY/ZsrqU8W5NJTjX6Xa9hHDynkEK3GA12b5CaiTjHgcjCBVa5cGEpR+
tVVuQRj+stZSVXmH++cIKapcnIvrduiqOariAL1tr3QFXMjSLA3z/r7w5Kqs
9p9ZsCNUTOL32Yq2evf+QCQU7KHE6K0aES/EWtDIiqq2zldUx4ydg/b+ufTk
nXE1l2rBTKhi881laziDnw2+W07FijuO963O13DzSE6G3Z3cGekLtcMHwIwd
kJ+7RZKX5zQ5VHz2BX68bZhucQr6NjFSKSOp4Sge5+MhO7AJ3Vi7LbhsXXU4
no1g5YHwCAGU9AKtfalQh32+EX3A5OXv13rGloi2ESfDW1e0mlo/RIf7AeLG
mPIiA+UJvLX49QBo0+N4KavOI0/Wlt0EtncB1Pkmp5sL7PHsCQX39x16/Z1u
9YnSo7mCfd7eYTqSM0IoDE43TXsidC2C1SjfjM3JpF7WfZ+10AXE5XmYcwwj
JscwoJQda9FLES+SqAJo8HPE6Wxs0H0BTI7DKvoriVe16VtlyPPwfcvdD/Zp
IfEL5FdMlcCxWAWy/0gIXfhao+ntakuoen9H0i+29S+8JvnwDx3eMfGbOO1V
gRlAoPznky1syPkgaNZSgFkDQHTLXECNyOIDlVgvkdav9uZ4mWVncbTjuRHA
RLEZ5IrOEbYhHb0MFnN1cTzR7BJBpN4NhLRTHTyVkuWjhQizbGtu328yW4Ml
DJ+vHFru3dVxlIF3hHIr/JADb7/30SFSHeT3hB8CtsW5w+3YjDunIza8iWus
8bG23invjIAFscUMiPFbJETp6TEov8iJk6lOz+BqWiaT8nIu12Oy3/RFkxr/
qcUiLN7nUHczYgUeNk3eEYzTDfDAkCQZV2Gut21NfE8xelxriTdmyHwP+3XM
KEuJEod7V1auAAXo7LSOY38NDIg/Zs45JvLdxfRTEYtCJPBhHcPMtQA5uAky
MD7iT6M7oq9B6dx8DuOQMR6F7hV/9cPMowOBBYB8vPZrxKjM5JgwI5FLV3du
Nve1Biju1PcsgC7jPsa5j6eftJYPmFlpN2gZQuPmmDGw/aIlDIVcyRSJEEXz
D+8t/1/fngtrutzoxS1TnESBhrtUKD37E7OU7hbatxRtB8O/jmzdWpp2sZJ4
wk7REcA34lw6F89hwDcYCk0DBhD7KI7ONTOFmq7qClqI1mxtG/Ni9YEEvqUK
GoSLlWbr6sOJzoUkjoy2n2aFX3GdgqardYn0Oqnasm0597+JkVmw3w8+RP7T
IS24eXnblvo36IFc3NUjcjEh8TpjUXWY9jBsyhbNyaQC4VdeZNcQgqRJSdC7
bCw8yPOwbqNW9DbMvENSADuszslM/dri7GDq/miifPaLzSUdnQU53EbwMAY6
Wg8nmL1jFftcYBqLisIsjmZDXVEbAy4dJCfTwzwq2hwFOMJsT2h0GoaCS0C6
0GOl7XyNZqjt1izb6C5sloRbGYRhKsYDg4IaWrEkNaa79HeT4d78k9pxXtGE
ECx8VjZy+2dlhWm9+WLmMJFEDJDk3mjz21U8vmahPAPWwhZ2jld24nKczM8M
Z1+3w9ZkC4w746R4cspcSAzs3fjw1CBI85KXJ71r96wDLlehjrpxNxQwGHEI
pOLgHY9x6rYpcR5lieyrm0x7vG0V1dC5qe9kB+WuesjtBFB+Y5pQiQPWLwaK
arhBF60vGibNn3OIgpEz7sFQvVSrDjVBlIw/FWY2MEuzU1kJDKruY13Db83M
qIpyTp4AIGR4UJ0emdScZG1rzh7eOw+1c1Far11x++npAJZpOP5MccC8Du24
i/Q9I9jQMs1EMN4bLxpC0+BtOhwBPVh2q0AGxBbpOG1U21M3J1QUQk1mCDzR
Pexa82YhrXuW0wrn8DUhEDlaOhnC6brKJf8GChp6fI56ujXy38Zduhj9V8nu
zlyDfZ6sXydO+UjzU3JYg5wY655XhiJ/WXwxb3IFqMm5r53WAf48WQPAbnSj
aYRapPF5FGq/jiRr2jFrVMss6ujRd4YRh3XW1Qf3NtatZ0mKUtkF/kBHsjuC
76IzFz4EgPy6Mm5L2Rdq4QDu+c44bjOdIe3olRMLeKqFziQEhebojAg8DjYZ
Za3SFtTm89yhKkFQltY45r5r8Vc/gvrmVJTcG8f8rSFB8yaSQw/a8nbQgPkG
YcM94myBfHpnDlKVYfMLBrR+RuuYFL1g90pm1EIUrP62MVi1OIA2er05Le3Q
aPTZa7DGIgRLubqVYUmc8/jmTbxDzVfNvuVFjni6MWsEQ5A6oRNkBUS0SGD6
zxTP5qRGUptaaKovx57Oubyn615HOkgh5cYA5Ma+cizoXsDY3R/DEFWU6pHK
d70ex1efNXLJjIL/sLKypUybMF/bvZnkobOMgZPcxZti2r3qw8lsobXuJeRK
AZc51phsKQdVFMQFvTU90PWwDIO0H3Pcug1+d7GHcBQvGjUDsfBGlMU8SfhO
dlr5fyNQFnLL4ZocfKl5zSyvS4VOsA2mPI1UDVblYZLVj6HMaDKjuwRX7wyx
PhsMkXDHuz6Lq5v7aGRss/GcwPNjLBbcZPLeIACGUP9imUQ7C7w1PVYwlYxv
nO5ARSYvDcXqBiV+g+6sEv9jIF5WXyLD+EinRfdUgBWJmcAhAPD+M9qrfdgp
LyTGtDQF9yjCJH6HdpRFTJjPAAddOqCqqT+jKGYDof3Nye1bMD4FC03sjgod
8X6NzceW43bkkZISlawG7ORzansl+qHV5dzHaG3lHtJC+EXEU2poLZfidFe3
MtXav25QGIjMHzBdmdNVVAbgrrsOpdwsiVPYOgRp5/uxinPc0vv44YqGblh/
0e5df1MRzZiJRPiBwZuBJWSEiewwTutzEOM1FCwxEdogf7pFgs6ORKWnl21W
mbZqvb0v8Xq9KkzpbpmH49uhEs6F7xhWU7SGcfI/3lZjaRsLrTA9DGtd2OpM
I+HVazOuhDMk7DPZ1oyNl/pcvanUfk6K0f38aCtrW9mxgP1f0qxh89oxygQE
KD9Mf5z8WLkIc/MSVccJeZ43YgdUqc468E5+DE1WpbPpBhI7RSYT0tkzsnr5
UbFcgE2CjucU9CIq5GLEOqS4i2Sn0SvYDXZsXwKkYfKK9OyQhesVNHZHMo0L
+I0AXbskxrPAlCWPkF0mxtRN5wWZSxc5BpwuZn60sZG4dz0lr/YFLScbESif
wUifu94uCYXF59jCUKn1aNr/ypeF6KDmgDlnMsA2pmDNoMH8k22/6ifG/kUo
3X88vyN/zkvBBPjbDjXhDbwTYcc+o2q5jN3/OLf+OqjxZBJP8Cv1xED3IKpY
PZPgArfldHeGi7IY+CM2OETHexyP+M/Eu2TMx6rWz8CzITiPF4yai6WHC6Mm
6jVIwB1I+DQNGnrGqM0ON4lzYLBKJl7eIzA5N7F1T4MsDh71J+4gBS3sufWO
5YU9ea2aFqWM8sLH20L/h21ojCj/SdCL8j3kbOiZ8tzVWUDZ79TP7HAFIF07
xzEvilF3CHbCXIIE8JLWxTBQk0arlpknXi9bk18TCZPslf9HAJDsz0hRDOek
UbSvI8LKPwozeuIeYar6FaCswkdZGxgdn0KdfIWOWzJV9+mMYTDbuIsaqC+A
OU3UjF+eM/gKej31sp/vu8TFZRqJQs3avnBORX31WNrsiJIJ2IbDqTQoJeic
gtleLlWgC+uIYvCUzHR70O8QvuCcWRb+JEBBFnZWzEQMloU5987tvJlJnHy2
OeEHnX4NIzuMt1uRSS+jr93RmH+HowBXT664L94GP3wckK1jA5W1Aeep1Lbp
Qe9lvenIiemJgxDmc/tb27F7o5KIYrMz3rvs1FwsQDjl4sAFDLfD2hHWaqG/
BoeJ/aCyjVFuFPjfS72UzF/n3RFbbGAaMpL5lE2H5sqtIhvkjOPMvrb7aLz4
VFgJ+3yvulsceJlxmTvwhOjTSnm9aGnZvF1qRYigpZ7SwmXucjNzzvNg7/zl
ZCQmNZ1mpsUQAUlxXbbOj9plqQcNLdjKOke1mYLK/asq54ekYTFQ+HOS/tOO
ENxMqT4AnCrDkMEAugK/RrS1Hfxd/Z4rdaFPG2EzGc1sP+/H9aSNtbQODpgP
Lk3/RO5b9GqHNeimA1PVSfrmPu+SSFWl8CSL2vkhqy66ha468Wynrc/Ej5tU
5J/uHBUlkngg5PhrFjfZVovfsyCGEfOConyKVxXk5B96FiTihaXbsCxNIJTy
84wfDtY5VHdcpoObzHraBe6qwT4IIu1Gmm0BZhIiHvpCdLFwmrzzk8QSLKiG
CVHNtaM3GA20J1YTCssLChSpSWRssm8F50u7fyIZFaIIrPTCzcgB9DJ8M5VE
xubpq7h3lHNyLvuk0+emAOeuat7OnjEihrpgAXkJOr14LgAmHaOY3t4S07M9
f1orsqFKtDQ9oSVQZS7fPaZIhMltkDe83P/n672lOx4ggKV6AlQWJAR1cd+A
8vSpVS3FtNzjnTQRBhZvKyTU4UQP1hz9tSIUvkC0xZiQfoj+1QCmMhAa642R
QDcg7Jg3v2Gx4Hv0UYBSa2vVPh4QHEh6qLbxFCAzDJem0cfLs7i+hPDPVkmD
zz1JjiylO6ng2ZzXky0CYA2JHT+AYHQaxAjyH0qb2yGq6lYPOloP53O7eoqq
ZroxXoRWtuAujxHQkjnDxNHeGvzEi/8Olz6jCDRPCofpQgRPLuuGud9TeLZd
328izxWZ5EXvMXnHIfcg8n/prdevTPOKyYwh+doJGsLGYgeIuLpJfcAFuJKb
4udznkbi51dfVWzWHmWIAorZr9KEHosBdxTTY6aR2Lf2Y6Qy9cBai0387YzP
s6hSu/j7Zq0AJfmVYKmfHgtYj0ZGvvTBPOdpCbq0iv6+PcL58jDV/AwHqclp
MzKvDgVGYBPWKm3SF6c/2KmZOwF4tIATKOguM37a39TS7c6B4mRGeD5xJog4
DxqezgQbYlLEK7Ca3PFohe8qYjSh18nJCekX0KpzhTyU3q4ufWu9xXgPqmoT
zYrN2MJzMFbk1b0m7X1qWqOq0KaYARLVi6DtybnTNbv3D5td3KIduWhxfc12
YlkiliK5LEua+a2r+R6zS3A4ll4nNhBRkFs2Vo/CtzREn9LGqv1Jrk2VezXB
dvCb6353L8gf1fJy7FkI8tiuL5/oz4b3n1BeQefk2AIo50GesrxQOdFGfB+6
L+mjNs0C1XTjdPXrnvdIfBZ6Deq+jMUIztbYtz0uzDsNHdWpbv4hXS2lqMYY
wNH7dF4rOpJSqgPbzLoy1Ir20pAJCi0z5KNC+N+QNUpVbG+V05ve+n5/0/sA
/MNWNFI2H/zvJ6JiyWhB+bbGHkfTtK2T3y+UMFuqOfq1VaI9Noj5e+KFZqJ0
N3+6lmeVi9TuNQ0X2rGMkcdX6F4ovIWJfZw9U+6NAmCBb+rEIVh4H2qrrlZQ
xVVztSCW+7TUyKHokLJLuwXKTu1xMmW+l5+l3sO1zie748UNDEFMaPaWVXHr
ei6SMOSJl7wvdjkEKxQQoWJCxNx0waFA8UzznO7uXto/E5KL0mX//zEusxEH
aLF/zL7qg5VU16yU9yaK8Bcu4AGvvc2dx4qOLpOBfbQKvajax/2WrL25JUYQ
kW5UOAWvJ+LBUI/RMmUrwlNhl1w1fqAra/UYCBsqCbOP+B9GVlleE0k04W29
+11LWhopGgVueRYTUaPuqHLL5I9JhzT06+9OkxtgoSrE//NfopsCEJhGi3af
Kx2pN0HF8+tv2cCmqipeVX94oW0PAFxGeqUi2wkFxd+DcvxxhDZmzElieO4K
jmFD259mw3MzEcSnJnYuDpeAitJSecL92QnARx6CCHFwNNVxoMinBHmgiyqT
JtLPB25oH5offLHEJmzAR/8y+ScZnu7ifQ8aI/Oa8uUkfCBrtOhB0vRWIBGO
/eot809dl8AV+vG+IWlWcyFx3oLU3yot2Np3ygqhspjBzWFl3eHQT7Zajm7G
Hn/KPyqVbfMRuwWYPh/1+89vjQu5kHCXv71yRRwFsu1i8Uy+KCooLnRfcgkw
RB1zaKV11xS46kd+xwGW+GO0lVobJWKmvJsIE7ogKM0WxmJQ/beTlt9Mav+b
r/Oq+2HY53G+KaW6hYJl7EA0GigSRcyBVSWzx3jZqVH+G9Tov1vKySbINd9L
As+dETYE9Tkth1sBRKY4iyutTSvkVCYKjc9Xuw/lwNqJRiwDKG0b61sPxuZp
4SmKs1iJqWKhOWJOBlpW7ScTYxg+iV5LsWeaTneDAHNi6WzHb6M44DkIB9wp
rfqFCZiA0e2m7wQNQ68THECkTwdOC7SFFvdlum4tp1AxENdDI7k7RK9G07jJ
HTdf3Olrc7uCKGsnZSGvWK+WY1JZrsNE9bTHYKr5xmW2D0HWlpCluQcN8Z1s
sMdDYb2gr7+gZry437pUTTQzgG3tFgGM4bZWSf7/I4+dAiDMOGEktXFjHj2N
uH3poUh82YJwrXBdWUb9vTVMiU/fxauC480nwaU/NEvi7jkIh507Kc5A75/0
Q/0/b2ow3GmeZIOMaj1vEZJMX3yFlCVs3uzL3EHqKhA+NmFg8ETCcWLYTDOL
55kbfmKSEdE+nWuulHmHc+4GAAhMsvG3eKA2jydXDziWmfzKerATIlNIza0r
dsKDr7vB4rrjskOvUCnJfN/UYyQ9uRSf1hsk5FUAnJKJrsHppgL3wxd3zxE+
nqWaVR1YQTwCt0c2qGa1c3CKsxKt2Y8pQgUFuOwjCXD6VE1tyih6GLeOJ2jB
EvlyyJrafGntpu0TEvcjMGGDi2ldahm4RXeUxY9UKfCLY0d6r8rV4YY3q/Wv
WJI0lwp52+sgKKom3yi6yKOcZYchHxKnifk34lqqzmcJoFoHoAuYgcZB/YVG
jTfmOLElbRM5uU3/NzPLeBpNgZlvo5JdqjvxJHo9q/byGT9C/RABpdWD6Jxd
rfzPsX/98XTU1J0n4YktTNT8XMTe/KHALyrS5MSNVOSKcpoWmApIUx2+7W16
0C0jNQQxqpKyzCPSw4vxr+MpXDBLDppR3/ztFelVzQ0nc6fVF5qfrKnCn2MM
07SUOL8zQEmBP7CIpfOJv95nAwVjjBdR15GxHaZu1cvnc81BLpW18JeW7znj
tSf0tzrCUrWSILQQpLw2QcQTv5w+6oPbFVb/YXoDzBszWYiaQKASrfpiyGW/
hhiHz7gmxtpDqhV9iyb+5HCj/75F4U27PHtCcxjMnKCoYfL97iCJ9JRDRMWw
vElotwDSBHLkhZYOGLGXmIdcCK/vXv3JBESjqFDjT+W0vv9clH1eAR/Hakjw
ToWhKy2EHUzLX3BFlXV4SOUySeD210vP53m6sEuC+IPsGu1slfZ9FxV28Cdi
n3Eoz3ziAyC8bmgkSx0JT9AFFUmleMMPRaFvH3YuZAqBuWl4Uf30rP2YfiWD
miQE0fkNk9MChD2jwzf7d/jZPhNsGhrujOE0Z41QiN7AdvhWSW8LoafaRGQ+
cIOctDT2vASNy/KwoOW8A1/ULnQ0KtpWdXLRFjh+kWyO7248qAT5hb9pJo+I
ANPAtWKKnM22uTCmbCclte+vY7DdvhOsE9ysDuAmD9Vz52px1frekDKSW1eJ
JTu/G2EvUrwzsXzfS8xe18bXfSpA3QEqyGP8AFTjdO/M25iRiLzitJuE5wYt
JAc34ozpJVlALsTGA/zRbYIz514OMyNprtk/FUOlSlqbqWBzM5SyKlpVUKVh
+SIui8tTsp0tHau+qN7aWT/tU3I11qzU5iNspuwTJ9VfCaONRRjOx/woV/Je
bxSKkjyd8WsduLFdnNAqx98ZBovl8e7N7qHcDeLRwUwC1C5+bxXA0xDphEBJ
IS1Xc4va4AMHIn9z9VLPE6J+s4MQC5W/MOa2vIXrAPitxn7wN2aa7D9H184e
vmuJl8trAiffVk7uWKliiKWUXMl0aKD3liFIgIpziY9De6QAoThoOG1XnC6X
nU1ybTcnQgtTo9V+jdLf/w2teI+bLoKq1B4DjbaTmi+9TFcfGk4FCbZVmVk/
DcXN3tkO8VNrSME489KF0+XcwQQkS3mBe1WltjPKzBAomyo24iElWex7NHEt
Fi9JE24jv9pWVJvIZnsLuXnkKKwibjjO2aUTm3W+0WtQ9WsvSrr0M9Da1BKM
VkbPBG9AXUJLVIkyzImp8DBG3eyv1P5g6pEE19dKbrFSQdm1k3cT85uEC2Yl
gch1t+/uIptdYlcfnlH4QJS8yvjokh01tgDZUrPIZz3ZAEpjQtvfcb1H9PK2
29uGn4fbu1B1nXnExodCMu3E4BQduQ7d7ZeqkXU+QBPt61vzoJVhRGEpS6Bs
1+NPeAhVoUDeMaTe5E4XmpEAMgTQjwVPlWHTwdwdddUDUU8RiqlUO4Wzj09l
PwNfvX4woqRTaycAGsRJHaotpZk/2+SexRLr+q9ib+FfKBjoC6IXTyQkY/Bv
rXqYg24y86XrBOpi6iJU7C3LMfmi3g7YO0dcBXUZXV26nr+4M4jLDyoRrRFY
0jlsS3eUGKFR0xirXQC8BR14twsfK/dWVhJcmZO4Nz6Eg0FlouT1VhbwdgSG
Yhi0FLvTQ6dImAOkuNvXOE5cabr5tuPVIQ9yNRBK9ERNQFQURlTEfpxYUHrS
09+/VOESxu4x/ImV/ZkGxHAx/Tli6RwPpXm4PeLwRWo9EuhhmkNY1RW+fx5F
z+0p8bkJCf3IKjVj13v6jsZbAogecxi7JAW133lOEBjQXwDlP2d60/URqwXv
Pgjc2r1O0FBt2suglvYv8oP5Tec4+oHPbwBlr6kUDqdFwhw+k8YD1JKBSX1o
jQo4kbX4X9D5dvOce7Ea/pLltP1zXJfsVFR+iGliM5aE7AeSWdn2KrSW8gmn
bG3SVstxH8wSa3dTtVENy63b/4PGx5A5Bn10Yt9Ns04Pk7gpcOGd8Hr/K37p
dOIclYqOdD5+jI24OhbE1XKxlwUDYAp2Oz6ojqRNJoJ+xkFK1hHJyG4clJiL
ilwruistDD4hm19rzTMR6h7cFZbODOvGAwLeXRoX9OTi2U2yASRYybyHn1so
dapROpiMwykccHjJFj/HafoVZoDp94kyKSlM069UcSwcyr0QXAOz4wuCSc4Z
pPt14Wc/ZkDiMjQ0OW6sH8H85srltaWW0ZUnLlsxF6CChVDvlBbvu1vpRrT6
KRk8drDgFAucinxqh5hzFmBvusiT8ON+2aMPkSB6EK50O6hq9WvHQC09rRkl
IeV04l3oC5a3CZj1TlnCOQQEghcZJWyVFNW+dqWTQNzy5AIb3zZJx7rSOFCO
l/kwuw0bx+zpk/cgE55bufGXJ3HVLxxdp9QWgZ5LljH5X6wMUiw1dbGPRppT
gM3dMcEpfGioH6Da/BTSbCsn6oWt7xVSJ+bFIVxCpiUk76tG3FFDOflIuEmu
HOFuRqPkFBOJkBpkcmcjpo2mjFBhKYjltt7flHe7YjqM39WxLwgV37WFnL1P
99XjGxBrh98eyO3GFr6nYFWTHQuH3cSa58/Si9lePUvqK9afOgVPKvANO2X2
FfXbOUMg2ejdb8pVVGAlnile2f7sQreNm09ZLo0YwdxSH3vfjDlpJhh8YIA4
hUMHsFnXWoyrxmojGT4+TjN3JRq8l8B9wV4O1YMS6EwG1gzblrrocz2bopzd
shS98dahBH+3DydxwmAm6GJE5q0zlrKoEQBE2C/OktzDxzyln3AiMvsJvPkx
yaJ0OP5gwMJagVL+yaT23LTJsGB95fmZ6y8FI8wXXMFdXF1GirChGJp9hSlU
4hbbmN+4STnqKB0odfuG78kp3eeofxffY7UzhSe2rRcLU59yjdYLW3TPdgTr
fcKdJ1CDMqs+VEPztX1J0bHuteB1/WqmRXnblhgVQ+dD9o7YjFciviY0RcOY
vnPKpyzxROlhTq6xlNCFrsgFNI8Ov0F/IHwTLKHG7/eGLFem+9vba7LT9ZTN
hpEUP+h7JCwi5+vNMZpreyQ/Yhgzy0oWNvtvGVppRb7yawBUrBqEimiB07xc
fPT5vYcCjtU/fwxEGN+214Y0lImyPsmwiZxjQaGcaqlF4+SpOqAo8FS6zFgr
7V1VaG8MUdiR4b6eLiqNaPE5KuWZXAapTklEtwW1fKhw2WUhZjVbxzl6gqHV
fXhbv6McMuza97LVLoTUHF59JEJr3lYwLHLSmgQ3vMqRwWyLvIbBqLQpYHLS
ma9mkVBdQPhzWxsyCDyjrjB+KpJ0QbskCgKkCCAaij1wiInlNpJ25z44CTQw
HNg2a3EFk93bequymH3diujRtshCkg8KlTkl4nufF6DhX6TaBFvBLw/xJ2Od
itXBP/+90chjOXNzRba5848CQAYe9VMYvypXCiAHb5pdVedGYDG01gnrBZYK
Xw+HwtjTrmzzG/BJV7XtSlgZ4+VvYpzbvmJMqKXzlVvqpLOI87iiS2pwRz0D
Leurnagj5B1TCw3NqHA9/bV9EtHns4eIFm4Ot4+moiqr8qaaVK8H7xzO61Az
IoD9bj1OY0+/yepLEVaa0fSGTbWBdjSYQjI/0r3P/R7G7ntf3NjXiHwt5VkP
4fqArQF19GiJ8j/Emm9lAFx5BusTW7zdnPiXXUaWEuKqS6YKI3Cr+IX/uh2Z
1od12jyzlYkLRfIK29nxlFHuiuAXyPS+AQwVwNbBIb+GjY1gxnLZuMuf0UDv
Mn+/ws/qGZVVFbvRJ04UvOhP3FcSHGsHiw/EfQmo38QJDnXs653mDBoESYA9
/gsOfMtslyRX6NyRFJz+5rCW6vxdl2U2IwxR2jc5wuGbTHgMSc6GGnqP+6A4
Al+IUiOZ40KG/i+7NmeNkqzK3XvSGeWC61IWXAUVLV03Xswx4LhWcMip4XvI
ogpYTWdXA+OIthk5weA8486l1/z6QvdsACNVKyrgTYwZKUx6raYbYRNeUhQa
n3WnVyxDVwIypDE2zG/8vy+YKkQrDz+ntDPKAtQAY0RzsvbWU/r4RWXhNMrp
hFAJ5W4UuF61/WM8tpOU/pvtoljDkE6Bjsml07s/XFVnh9Q8SjQ+yerp59G4
h+iyd+JJmhIilumyhBs7D+WCT1IpVWfZ8Z6TEjwQyBM25EDU0LuFSG76Ui6H
cPg9SmrYzAOxyeA5gQCfQGn4PRVSsTJ4thE9wpQNH1juE5IH8Z/gxrREibDz
0QxvLyv0OhU3sm4Iiw65Qe1ZWQFmFxKYM/t+zsV/GYVOfNoJqxPsTIxgyqx3
gN+lG03wOq1CjcHPdnwJWn3FhKDIrEZKcsz7UQdH5IRxI7svALmf6/7nm4HF
4SN1IcdpJpMDmCkglBmBmzkS5Kjm5QgHFm2xcvkOTZ1nQIKmqqiQJc0LopRE
6bOab8do35DNYondSIJecLPPO6+UglL/L+Gkdw9rhlm9ZBHm06ihwiaaeuAk
VISRg4naVEdFqPTbK/dHsSZdaAHEKCIt9thGUmDN1hywmxfujaxy/lc6Kgz8
DgEUKUBNmSpWXBGD9XAQny6cAQJJhXNJ46+AAMrVW05agTwChoQcuLz9byKS
fGGep6UNEuBDZGDASm+f+1QLNV2JnRj1wHye/czEJF6wezG/5qAkS6DUZwJM
hTHwxcP3WwI3EhLN5WmJO/I6SKtHg8N4LUHS8mUg4i2QkBhVTUiCHjZxgSjp
5TERj3TwC0GRpRzg5/8EjFKMey65JeEZ3JWQnGbFwv8ocusSWTKvDUmRyIeO
GX63FR/oEcb0Q/kWNzIllFGaNKNts706Sfgh5R259ND6Ygq11h46h5FmDe4+
zIH9iC5f1su9uyVpgbwA92HXSFRaimgb+H3kMF/i0e5dmOkIrfKYsQhFyWmJ
WVwD8NJAqwYBt1mUjizakXzFlVWzzR6m8fERvMVyJqbvIDkwe//qpMC4+xMF
Xc+ay/8kZv3SgNIMuswDBLuy/fUimDJKzqOsywiZtvvpEW6xoZmJvrpTM7xS
hOr0vsvr7mAE0DPfZwzeNBISFOZydk9/KD9H9AllnTbWcW42BR9482dK2sEO
dWiRdB7WZ4T8+qwF4Mf4GXVLAPb5JkDjfsdcAxBPDlwlRwSb4XxjF2EVMyif
yysxfuo4T1igMiXukWgBiTbPNTvdj7G8yTLV+jYQvu2IVpZUWhG/R0zUw6Yn
A4tTYecP+BJIcV7LD3IbVE5nqRGwSIp5oPsqKkZM4OkHx4/1X/TVy8TxBF0P
njnvso2wc1S+sYb0IAz9W5/TlPD5Qr3pl5X0g+1YXm6F0ocTeejQtWeL6Xl+
A20rp2Sp++WcUGpnGRo6QxUkn8oTzDS7m6CVBabwnGsvhQMTgZynesDW41Z0
cQ871VxR0yq5mgodFXeVUPcZpnI1NjqzqeM+lrRZAaaImbE4DcK5jgZ6BOjS
gq0oxRO2p+dY1OZxtfvhdZwGAPTsBQK/z0G2/Pj6NMkVqgJSp4oi4mt4qs10
rs0rZQmcyLFBSp+qMChZo5NqYxXMt7ByUk56B5DSbw0k8JvyVR4BPEtPuXN9
Izk6EyOH1OK9QEhb4nuV4EJti1coox405m/lUtJUk0KrMpNPi/IEY4e6LLrG
rhdI8VHCF4tFjL9SR9RcB4yZFmeJCYjjdlBTdA9NQhXcd0mwxIVmabsCyzJz
upRGM1tcoPBXHAmn6EgXtwucmxY9XWMR1mWy+Rui+0hp5l/oKEpSv+LwGogM
S60DwHsBaePF20i++3wbOxh0Z4uszIRGJbdknwLehRTsM6fezBpDGzwzW+z7
+Kgtb7Q24zNI1cEiRt6h3UlBaEx6KRiLde3vXgUbV7sQGXcHP4Lm+A/pHqcl
3v4aTOWMOoLxiUeSbDQlsmBavLafjQTFhB/YfqkbAN15v1cIvsPHyYNARjSs
Hi8o16mN4zfpL3X1Pp7YlNj+W1FZUzt4RNq1xnA7frxX8FklLSx+Mw1PuxYA
VrhAgRy5pTPN0tvJFiFYA8Z8zypUtP78idfa+MiCeWOTc4lICzoYRr2ix+Wy
iUwlSCKZFA3rrbaLot5RXDWitChFNUigaCnW6nNJR6lzJJJ65JeL8KSqE/R8
oSi6L2myxVJqLDDb5HN736Rv98eLbWErY553olcAZc6Sw3O8l3QWVeaxhlwF
2XNFNr+CNy7h0P0r1Sn51C58V+67K31gXh1FUU7uAx9FXrpyDCP9kzc0HOuR
kPa4QPcikT5nKKdEAJTbn6MkjIKX7lyjmWvb2qbGfywfApi7ibts8Bsntsab
ne1re2YN+gSNO2CTAmxiWehlDxz25qKPTfAbfnhjETnNjwL3FOjPNtd1eMHx
5lcEtpdriHvBrSsPSSrU+FQh2V8I6JL6wvvogORKkpewZcH3JDRfOOKu8Tdb
JAr5ie7+bDWYszrX4yyNOsLOFPHgC7UHfZ8SLLaLR0SHI/Dszg/NFZcqLLtk
3Q3xhBSdFdENzEACb4fYBDceff6yfuS0UhI0M943z07PO90hcJV6Ftb20t8e
PgXWf6Zh3yI46anl8XTn/D1VhqRMyNxBDT2RnT+z/xLKBHkFXkrTpRWWnLIo
okjVLW4AKmxsj7wtqPNChc9/Jx90W0yXiIn7jba9A5ySRfG21W0SY7xLLy78
Q++8uG60Xn2auckIYdVxHliJzm43Mn2ylJRL4Rscf9CGI4H9Mvfvwnjw9Jq0
EHoY1k3cxrnKR7b5DdxtL61dyRdhpsLG+TkumGksxNOrdEajxexpKv5DUD0F
qwvVF51rdNNwcLTfG5RkhvsaJWU7CSLNryS30W0h5Mr3gU/Fx0uyTO1BTfzs
AOuCX4zSgOLPolGv++kI919RlIvaWY+Ze4jYhWqr9IRpsmkXIzPCMSn6e27i
gfeIfh3qj4Hp6i8mH98kDQwPRr2jJ3gtCrKyOXlHvY4GwUiY3ARI5l297B4E
qDIb9uSncj/l4Vz+/JcerJQHkw8uCDjMunrMViz4qHqte/O519Mk8YyDHnKs
NB/LBZ6OQP91lrDY9oMWFE5viq2tOSpstHgesJuQfZYMNISe/iirdOEwGQXJ
vJK5nI1Pa7QTaHdDZpCfAiOM8P5bZTqhs7VX3inCmmsUN8PXJwJBn7du6Z5v
CqNUBTzAgjGxyfutucMw6LXTwpaiewh9BUQNAeTFShKmWERPhnICVvWkpxqk
w2u7yoxG0YLjQpl6dKhSeCMFmkqJZ2aRzj5Xea/5MskS8POG305f+0v1Wl6d
uBfzUKW5cIsyehkd1OKpIrN5CIY+zzb5SuLp4rXv/gwYDvfM6uo+er0BirsQ
pXZwA7d8LEX8YELphmzhsODjBo8uCZqRtpNJxe76jB0ydWdMudTYG7DMRSsz
Abe4pPjo4dhOX1RVTEaM4Bl9l1kmNbTUDIs2vzGd+s5vr9Klow4EQT2jOCCu
7VWry5bIHAT5Wy+2dpqB4NCRe2IXmUFT10dxZOupzJAqun9E5L0BIEuwPeDg
fhoRa+Oy3rEtTT/rmrZ8br1SQ2Sim0Dd6rz6badmYHFlyRFSNe+FxsVw+/DU
OvwnSFraEvobM/mWdcsyJB6s1uy6SmNUi3mbpR9GQukyyvKNiuY5iUB6wK8W
bE9nUR1sM0CclKZk7KxwhtUZc4aBvCxG5oN8ZdtlT0ee/UxldPcMgrOvl+K8
Dd+DKzp0jvZ2jlYjq/GL5vyRtgMaThyjBV7cWkmRvrsYmssK3u1fEIzA9lJ9
0CbtMjZmov/xXapaNdtPVtLu3QGsdffjmKFSw4/WYzsIbYOuD/3le9rfiKC9
DJUMzNHajMwz5Sswm1nf5VYhR1bOeGwMMZAz9/Q/YDL587FB2Q4yF1bP5MGk
FUk3+IfDfkQoQhIMFB1b/Ny9AOpcUnERaLVCJ1cjE9aLsWASo7C0LwLHUkpR
Nbq29SECo3uxP2qn/yZfIPNEZt0AB8i3Fpf3KBn/CyeonXnmvDKuGs/eEIQd
ecRdIGyIENgfpRxFipz5snHODmv+S9m1C02mxwCJKsjiWAx7bQW1HltrGTv3
minWWVeFz2w/nK8V98v5spbEK2avVG/zLTnrIeHq1j6ApL7q5Hnrjyq8zElI
lUxKDeUXcxI9b7L2NTlfNoSqZlkAkoUuUrfzXsDagJfj8vc2jdPZLRxfZvlX
6qRsbecAG7cO6qboXSTnrdUlOYhU6IoVBiG2VJJWZVRDi2uFmHM1bsSrrD+X
EBfvNUHTD5rdTGcD49yLM6mHsZaLD99s2Z5pDTi3/KSN0JywMHM6upv2DonV
jgqq62kCKPyrjWWHRxEuombRfJZs0lDLtOyXolN7vjlA1fz3zdptIwRKyfFw
80rZ2OHpP8ZZbgwDtEOW+prk/pP6ODVEoR7OOJ0UFmYNXlj4WBXG6T175z7E
dwzIvLvM8aHgh2L9tTCay8/GlRp7pIMpAg5wddtB/HCHjo7okUVwnkQswlby
QylP3aQ2shWdhBjcqZBatjAOrv36w3dZsvgD/u7rdgiLRcbC1fN8kYAUrzo6
BdVoMK4yF7lJNUf5aN20BILdceGFG0JNhMGJWGCPao4JxqMakoYClIy7J+om
m5gktW/Onl0AQL6cCmGXyQdItrcTxtCkZ3YmDGdDh4dL9n8Nz0NhU+NKvaow
lZK54xiWzgLydY+jQG4uRyYvJWe2sBxkdq4/4ynLp4fqKtwW9L0uJ+oue7MT
/SW/SJdNHYaHX8PwNrkuy5aKWPvXsuVu10CWCsXi/ACNNxYiq9pyFxhZDVLU
4zT7v2FUzvr5/9BG0xIwbhAGdKchKgXgoDYbKEK9gGznY4zfQMzaEzTyUYtl
g//Ta/1IrNN3JdUUByp3d3GcfHs3RRXQQBtqHhBqYaaE/ZKRo+sLMhNHl+g2
MqGSxEXAJddjwTCYQUJRWBPNoLV+/1PvOd8O1Kkl9DYED+jhk7cMpo3qsFWB
t7q3hFiXNjBexRqijOddKr2VNrjSLAIp0zigi+vsmiiBG/bkT+8FQ7/g6WUu
FXt8aPTyFJsklq0SPPVK2os4dmV1rZ59y0l8LbzfZJAEyBX2Y/SD+UQYbiEv
tZIdc6/De2p7ayDeYTuHDMSRKu3x32VfKOt1ci40FtkGnltoT5A/LK10ND97
8NJNfllxRrtNNK/01d2P5CvEnuZVWwD8kRJcdwGKKPFfgviOPV+QBeF04H5y
so1BOQMLhv/qhpNpfk0l10onHHdn8FCjLPZM8XK+/xdVlVLUC6FrOsp5P0Cy
0bDzSTXhO9Vg+y5aSXMzBG5hwEGVweq6Za9zELymxmyNqy53hlk+cEC3Ov0M
OHNMcXgbhVSyFsxJQ0H9+14EBIJBEj5TNKEphuLp8yUYad0ddghP4naOvzPC
YuSG9w+htAF9w9WO+teUU+eN34D+PxKwbGZHhOX2rY1qJfk3Vmvmon131jpG
RCjILG2LjwT7ONvbzB+K4iimg03mEWpsY1h3thvx7lvXhOYDRLqX582jPEqg
6+7clBVAE4OFZOIxxs/44En7u/83TDCnjoxsM9bCDHOi4eFXvJo5ZK4M0ZSO
Ae/kuZasD02Ee9FCBXLe4kbGLzXEl5+XN5TC1I7m2Rg0KWpHT9J4CNMiZviU
pK+0EaiwiF772oBEqQ9mrGjaEwFXaNt+BSLLll3f9YJuGJWCcc6Cv1V8A2Lr
JEojufjNtGta8wk7jO/BocW2BL/Jnss+9QU8bPqXE9VtIx/B4ancSfY7CFYI
sy+WJ9nMtXCjtropcLtTgKgQF/OaeMMOFvLU+bi4YFnDzOFiPcKfnaijC547
pRh0efs49ZDOM4nI+KxO6Cn3KwqHT56qQK/m6NFmw3VF/bEfEc5yz73wMZIs
6KOX3e6GmJI3l+xKeJhswaoDXnx8nm5FnMt+Xufhz0UL2JuC3Y4WPSpEud3S
FRGdcyTsG+yzJPCu1q7TG1ujzICQN433IiLRpu0wh8mzLc2Xzt2XYJDiZBHH
J4//JQ+bge9FIoVsBT5KxBdvqN3YTmw1pg6nsOFvuzNloQVGW9fII0g0xT/d
smkQ/IexVxdnXTydKFXSUNLsoiefyRAH/GEwzw1qtXTE4+NNAWBlDOkt/Jgo
m4GXph9Ktur6+s6EjwXWaHrGO70OGFtjHonzWX3U62dI2SgO5Z1Egv5CmPHy
dAqbUstvK/w4iBVWGUjDD8Za9/GWfCFg5BN4OYKDCtO/rTgr0bg1xYXZ1plP
KNKhLHXb09douzE74HlqGMwTbzqOGTNfFVU97HjzHGVcowLDp1WYoONwOD+4
FtpQnEf75rf3xBBjM1BQgZD7z+HDHaJfdM2WO1AA5I+AhxQbXWx8mkg3HFnv
GF7m9i8ovyTtn8iPEUStZLBe+PhfwNscOS4DT2HA6tpeyozA/rFhULUgU9Vv
6lrgjOEWKOb4lImOdSCDSgSWJ0vS6L7cGQQm/qlCdc9lEi1BzdaqPkYCdudO
T24BOELNq6OhVTBwtJ5YvQhJsJh9UcB7nH67MvsPW6G50aMYXLauSBBXFsUN
NAcl4+J1635mbTcBg0gNyBNe5po/qZIYq+O82NCbfJj/jJrN1kl6tEAIei2p
rizgysHhwiBOAwDvYAndRVDC0hGeSOnlcV5gVzUc41Q9vgCCmPi3KPu1fH/Z
fOI6kHlkTYYpQJu9XP1LFVkF9hU5bn1ZkFkBadWNLdbWFMw2CVJgnqOGA375
9oDTgjya7ZK2QcOPNBvOngCl0mFxx2/pLGHZifGJDLeAiq7UNkEicxC4CawS
BE4jirSal0ZmDBOEMLCsE8DWg255n1bg2SW8OaPw/pff3l72ERN711U1Aaw5
5whMCaomLcj/XWavmOFSkg2WGGN96HylrmwNS03t7qTuDefHaGdgy3r+DsE7
R3rNcee9nbsyYO8b0LuZhbW89mpDf7g9kCUNGanv4/zehv1Lz9j7OxUuEX1t
xHJUQjbWkD0W/u0PwmnIeZF47J0eUlmEJeicQqExPVnYLOqpMb5l2yBZ/zlv
XATR97UrWkMNnOOt/rUw3mOSqnUwQZmyCSs0cXJFmspdYrPGip9h3NLARFJr
jJnmWiIqbU5eLOGhHVOomQyTxqMuJHZrGhoruKPuplRmo4XS0n84HJA/KjJp
LhUwFq/2MaB2UQGjZGx6qYohcBw2HMtE9nnyBLYxq6yAMl9kRyxG+QASurr6
sUe9xW5vrL1aDkslAMQJ3Oy/57SJdfZcIgvFE3MaZIT63639eUz+9Uqf5Dpd
zhYXNgh+cDFSlgcNHtYxRhWGMJcqCsFFpdvTbgX1LWpBSuOK2SW/M5ZSXPU2
Hw2fojVjVDNbbVYbmpa8Fthx6cR5XSYU9mtPkozisIdJ7TuMWemVt5NFICRS
RKPTLj9PuNeWBLFkel2IVWqGlIW2tMvmTwLGp09WOrFsFHp+GMl0VJ0SIKnQ
isSVdW4pFhF2LNqkknavixLgWbKxLVJqeL3j4+EJhYbgIyy+6eQUxoutJp37
TgcLyYj8yn9RvzDxFCkCkzU7XUsBr46eBLcdGRE3eoxjlGNRMBbOq6CcMyPs
T83Kds5I0935MeE6WsiU4MxZM2+52PSdtoFRaLTZptn81OdtAbbYhyzPtSK8
My9oW7HyrgJ3F1hC83TkSHxmKGwhf2UFo/UowSMtSYJvDQ9YdeiUY9FW9Iso
D3/4z5VmCuMx+XoEkKh+mz/aQdcyh9T14SaBbbnvljqABvYAphRQgG3Gzir2
s92f73xSINP3rrEn3ssuMiWE0AIZHKjXO21w8wt6hPTl+Er8Hyqy22MKv89S
XAm22g7jU4DWloe5YaTwVhqi4j/RDrSN2tjNdSTpeyHLLHM0bxSKxOMznf9T
EHn1fhH9JHw0CoH7lcdf+AkZP6VD9uDS2r4Mn6YmoVOds5N5RBX9hNjIPT+M
eA9OftG4AGiInnL80F6L7KTkrArAtBOibi7ohCTAmk++sdk4rJDmak4u8y5d
hlandmQv2m6bT7a6PmLVmen6HUkMQMj/xxMGVAkNUxzbfMmqE601HlkxwDas
jTL20TLE+FBRJXq/syFSp4IANFwQ5sDTpkf9hC1tDl4dmzfrXyKaZKI+U9T7
cQlUP7DZ6lbb0Dx13ueHjJsAWPqhUeJbMFyeX0fmAOQKOLwbOOStnyecDrfJ
+ZT3dB1/MxpNabEO9jhhKy2VzS2AeWTXG2+HwR9VU2/DX8F1DQz+sYua6wne
4Zuvf6d53DP5lBiwSvFm7V8ZoV/cu34hOig1ZIG9izybkMKHpo35Sb/5r5qV
M2qalfRPVJjSKjB/YEPbDyxAGIHtPBak8UN6g+IazKHADz1Z4VaLD7LQ7eYi
YyVGOtjU+FFIMKtDOhii533xWJqIABNbxpI3Q+GKwka820ly6u1wQINZiHHG
N6rEhIYPmClcycxi/iwOuhPajOhRRZ/X/glENjEodLfJpM6zSNkr2tdlxegz
Een0IDlhG5lPV4mttayHcXOXq4bcoIxoinnlNFCBNGuw3nFt78tESVSWTog+
QXcstLs5h9EGWky4qdIwdmyu41NZ5oydnoLkIehRX0yGl7qRiHuqRXtFXuY7
spp17MNKkg/eO0IErasDb6BuA1F38RmD2TtzrnnS1NlSHsx+zDMCZlthg5jH
fr7Zv6qcvIABVuOGNwGUm1Mu4LbTwufMcWojmXLTnr9OqGracbcDqcZ3ct7K
ddsyG737w0ntKS09h5mN7ygLvvEXQmz8kTbhE5cXgY8ZNfCBeNf62XMGIlYM
0U1BtxmY3kxy3DDfT+4iuCzufvB9yCQHschIJVCEdNAchNmaeZyzAksfShkM
4cdkYNMz+3hBK5C9jBY0u4pCMFAo9uU+5Weq+RFV9kAJbwW9yTo2v+0KE5la
VGP+86pUKfLsb82x2egxhpLwbjlRaE+o+/WhaR497Y6rzClECDYJtOdSIdJz
80rXjUou1+pEJgtx4EX/Fck0ZJPrxz3ArBZUY/GbcXwM7lrhP2cVRBSJEVMw
VdTTjbzCvg5zgJa2NzVSnJXAh2MFXrf0eFHKUXcoN2fT2MBONRS9qJGyYzNo
Ys/XzPDBm7yhzU0TIXJ0CVIxAH6qrYi5Ugb+6Rd1m0emCIulEqPx4l3mRBMH
6f9jrYRXVgBpSFDgCbeT1HPXcTFab3d1hNDhtVae8EJdxUjqLdtLQgSELrIL
4xMIVANyWAmChQb0Jx32Ld6PbiGnHR6uLGQDcx9dA6ZQGS2MXl2eRB48LfJ8
/oq1L+w4DMf5u1FH142hJxecWT8ettaR/y/A8WI0M4WIEZ5ZMiH3mifeLKtk
6QOMoWrGGg7NchrJNG7UeaMFKtwg2d1iWTWWYh5dx551ycnEnajsQ5vNSs92
IskZSGq/jPExHHUhoqqCFrHFeAvU6+WSLxxgX6NlgzW1e5rRVKe+3aORN7nh
Bxgb1nX2F9DX1ImAzLcqBbNfrQ5MrXz0+OKpU3XJO5QIuaW9HID2h/WznpyW
Hqy1RmzeTSS0bnGwM1CLdj+JinV+8mH8I7wEmnHwb4lRT97+WsLWbh65DgkB
tZUQMHD55vRHxlu2FT65M7xeqL7QKVczB1WVHHWXX4XH1YEep+iA2/tjos+1
9tzoKextTXp4DdnPX/9NXB+JH4edCBOxUb83i60xEYxUtKjg9UnRE8ZVS2gy
nkdFl5wMTqsGIL3FcKi++W2mXhH99XFxM72e2lSRnwiQSK2jFUmYfHmgDCUR
1Exsi5OhSsYfAx2L0VTsHpgIOMwcgQn044BIXLqUNdMzy2fOPad8wk0mck9z
HITqoJKVgPFJnqsNOHHGGzO/Ys33wkS2FJJemeob6HaKx+CRm0gr6Gnj4OhX
fi9lukaeeMXmoXvG8WV1mSKgivj0pWHKP1C84862/wm3M0l13bxqEYm4Ab2I
3/WGWPTNOIzHPiVeqIwysYo80CotVSpAakNrWoRG6gSVd9SBfxYQCZyOi2G2
ybue0PxwWWHt6QUAJXYEF84PWgjJkeoLrhvTArPNyP0g1wbN1YTJKn85hEp8
TiTGAZY6yl9MJMxNnqmjmVLudHtEoUMWo+5ndSyKS9DgHcnAr/OJrnSmPEnY
d5oKr+9/Tafq9Mi55tsbsmMDfd0TCJeoFCmX0s7Hl7mTWEqXnRN2FxCZ2Y88
UuSeNu1M2r3IwDczZZ1zd4WggpYFxehYAtO4QlBVFvQgCrNArbl+hRTIDXBE
fLB34pyTFh/IzSEMRwc0J9wSHr9y+xScknjCX2AZDM6M1K6HVx8QAXIwTII1
knsm8GlJvYp9VtZHw9lsH8afqV5zNG6rzUo/COfYsoGozz6wtCbb9EelLIG9
1zEstX7F0dsz9ej5aUiCHKgKYBolMf0GzDQhfs6skUwBcJOcXsXlOoL9fNuE
pbTB9GeKuh8/Oa3X1JDJChM1+gIgjI+/nsefTh0vAAZfCGvS3JS6ztF8hxWz
ubunKlGbyT+Y05Ubwc5wOqqyF19vLNp+QnIkGbqXi4exxEe7zxdy7AxBL5zR
tiGR+SbUtQSsIAIHpgLwyw4mp3pJK3WJtMr1nxOS0RAPWa2OCVR56d33rxhX
NZVGecJ7czR+mV2rkaPDnBLl0704G4sLt9eWYq0KbglpdndOf2vCu1rieCMK
hfwGcVuqQY/T4WaLg//7JVSKdYQn/kRBf54oMgpS4KP5uXn+CpxFzQfs539R
EAB6l78PeX8CXHtdPubGB8LIIbKOFNRP+mHJJNhCku6VC3QVe7lQZcrhEjND
87kaE9vJ+9Y7J6FMj6ckVZIjKDf1aYi05+ReTCAZGcNt3FyIUAUfnGhEudwI
kexcJLm/ILiYLmGwA4jAX/HNaA3rmVV/7BN8pgNiE+qHaUCzUmvwkKrLpHD+
ldvledNPTsUgxbT1Jhri9aD3k2fY3CvOVr4/PC1nB3zZIVyXPFYeiU7tnBNR
KNW0RZoL9dIhb0n0+Wde7tNpHlPYzNjlen3+SvFNquBusezu/qC2fqIxsMfd
2cXrXRZmEs5Li4FeTlht5OFJvGucU5e8wE+pZ/AuXN0mYl4Rw5LlD4g5NKqB
yHhYcFUaGr1rIpXj32kbgB5WugbhGp4sFOt1FVh8C3Pr38k3ERk1kiQCyscO
lS8NBvUNzJ4fiKQsoyQJH17AQoPik0LaFZpDlfEpaqMyWCdLnp/coq3UIxV8
ZfhpcnidwZ7FQwdMexnpGO4rRrFWBjvS8gu5fEuiVqAgyhWD4UPmRARiQxlE
SBm6Wxx38SRmJZEfHiO5hnnYyVCmEweNE6lwLMFAnYrgrdjtCVyhl7AWwjYV
QGFQsyROse6Q61HnfrgAL2Awvgs104LH+dMiFf38G1z3G7UNTrUAb1fprs3O
UCSYmAiiEdNQPut2zQ24RymwECd77E47eKFy9Acrji9fcgRfpPJ+HDydLgnw
K8WNutsKwXN6kbktgFpjxL2aZmv+2oMxaAYgwITmN+RxEaRRkloqAQmSi+oQ
FJveArkGBMbDQQ7x2v52KEC0Mz1Tjipz7KxCsao6YDIJGim/KFAULW0q7tpU
rhD5/+JAcCBsTizXP6QbNPe5xShaoHE1uLRDEMD/cHQhS9AdzAR5ZvaFR6EQ
5/+/LYlV1jSjXQm94kuk0c4RZAmjUb59wlB/UyYOhS8dfWLV/39fR+oosSN8
VtTIRhB8YB86XtDJT6Lv7go8QTGZCfWLUXKTcwm0dKChEGotJqdOPDI1m1hs
FnSf/+mGBlLoIYJjDiabkSm+Mi6Eb5ujCYle97PcYYuZWNwxso19zSonVpj8
eGKy48f5c4SYUT9F8QFpGgU3w5y5jc7Ew35sapxWwKRr3gr2mrxxNWPNuj8C
hJ3j7DN7wcjoPT+dBv56zEBIjaQmqaSAxkueC/bndethkA3W4NYqbhNNwDGj
fCaqMCBYEeJAVIbjq4i9y79otBeDxH3ciMOtvsMCth6E1sf2Oji97scji1ud
6uykmcl8lqQKhvkPmmXv1RqBPUKd5xqMf5SsptBaJnxBaJIvXTlyQJ6hNX48
3PpHJwuqHEcylO/JAUIdjcs2U6aTHL9rGW8QD0wGUoiFzpkPB0lRDiUCeRuF
MK/rT1VCaHBgMO5SErmMv+5aV4ixG96sLr7s2hQtvHQH42dOrNeuB+ep3OIf
D7hVGvBvyAn7i9dvRxiFKX/lfuyB3RcCJLXF/jyKu+yDKOSnmWQA3CL/31pH
aGuqtAzzX3ICXEVBKCz487hq3dR/XvAaqWECT46OVfanGLl9wFUm+1c/BzCc
y+YH29AtljHTLdlDu4Pnm8PRTY0ObV37OqVyHHCwx82jHqNhA36bKeXj0T5w
vCfj0tMQVUE2l4KIvDGXUT/GyBnPbCtHISPNZ8Hniarn73V+Ah+n1MZMM7EK
M4kl32T/BPv5mDUTYGNnAwoYFVgtHxBA3o1gdLFZvScs+xRmau1TmecnCF09
YKt90SPvLjDQmRvE5FDFxy1FqNWvsacE8Ctd9tQDXRYTuuUiyNPvvY8pYOgO
wd0JmEyMy2RYX0jT+CfqGF8l5Vl212eO8arr3CAPbloqPH+JdFEB9gTvbwNo
ILSMhD4AVg+zefWfV0LJlT6cmEU5ha7E/gC5EdAeW26HKmCOWNtyVUQtBvtW
mRJaGZ5R8FAlsnjTCV4EnN4l2POPupBWpbrUR18plK05PprGfEk4iW3WrW1/
/uldjb/Dj/D0i4IAqN0JSJ+JZjRccTgTRMwaFBWYN2CS2EHpbN9XXkNXzjfF
uI6dEDwKNULXj1kS8VQmOb45ZfwjzxVVl0OjzXxHDitAbmY8pkKlt5KIWZW7
gYtzPNek9VqhSe//CPyq3SNCa1xtWu84i0/ixY1yyeIcYppsxYNFn753aUbX
iBWR6To+yq4fwDDFyQDl2nCwg809wspgIeOsMmCcRiBV0mTULGth07A8KvHF
vML4+7nxzNMao1N5CKFVMAA28uLGR9LvEzTdTJFF1IJV7JFcLl5plzyCOYfV
zR/Lej27aO87nrGS9KxCA09yQ9ZY3hqAPhZhUKKuwvlmOSAGoRPE+t/H5eFM
dA2PjaTtlwCrNC/zbRI08vir+aDsEjqTRR/QN/t+xJga2am1BhtbhIR9Xx9P
MXb/UxhnsoROzy8VvimAAOd/8f/iXp/J0DXkIAb6p6upDz1vrRsM/gT/8nSt
KZw6sMfEwGx2QZSJ5ECn9jGId4imlyznG8xqOqWqo3t7kFN/SIvIvTB6OA+m
ZlHqy1pbJ6MAMF9ErpoYGGQKmBovmb+a/F9tiLCF8cL5Ro0bav7+vClpGmXO
7+2FfPvMBB/2MAQ5VD8s/Tf+qDoUUk0M7sE6/WzMZtV63HpfoR4fpEs8sdmP
MTNqKIO+h1kJn3MaeyxspliABSYHaisEgwDsDmb31kZ5SN2VzxJgG9FOZnwt
0+K0kxdCS3glxhoNdgIoT+gC9uNegDwUrJL9hSlbSmTqAsK1lMeULHmv7ip5
nSQMx+M9JERItO1j5sY6Ue+nH+P4iPJnem+SferrL6FmEQ0P8OLHUHdmZcf4
E9kaSDtIdKQ1QNKwPbYu6lCJjGLw+Nxz+sY/79O2QfBKnL5+7OMJBdlYowc9
geuNCzjcf7w1sO4KvqEl4fCCLFH0xdmHiOo2oOJPzywebW+LSpKuU6KXS8LX
YPj7MeNylWun0HCHoGMvO8UFMd5z4x7yvqMPNKfr3gAWby/nfKZDrFvlPLfk
11y5lOaNUyj6v5uagXgbdinV5dyyn1zPH/FVFLWXHCnWjSFsF2SEC7kgWMMp
cI01Wxexj7UHOIDOsrlMKHNWgH1IqUaHRu6+hu/QeRjxOOMsvDUV5V++7/7Z
/2J0miO+7f96THgWFUA0QL+vRdcCWhvGXJkmHF/dnw8aTn8sTQ+zUxyvOUYv
Eb49oIF66QjRyqLSLzJRM6NAxhOLk6RdS0Tx4GZlU22XSROyFfODhO4CUjsa
AbPKHcSkcGHA0yqj/HbmNySjucsDgwdsc5J1zct6cR7D6K3zcm9S7oJMm9Sw
lpI3MnCNHxGqJIZrxzED1HUfrqZKkgSqYeIq99zmdi2YN4VGqm0Dy9f5vwiB
mbefHRUsnDnmNtiSdrDU74h/bNkY/rz35XShA86vp0s9wYzsK19OCMQtRGaj
qGMIGnbRZMU0wXDZqReVH0oPR6kBApjrbJ/mkzaeffVgacY2LcpO9W+2eCak
7lyI9voOn8II/CLm+nlX8akyxaQYtShw2m+mkRyXLWp0LprpQs5xXMQAqjd2
7bwJjVmYIxb2jrIt7ycnvAp8SlVGWJhgrtSMPEpjkHFnEaXjGbyex6TDGp7H
vGD5e4iuV7fZMI+BRKY2VZbbaa8vjt061WLrb1pvJ+X/cKKKnunP1f4MlTND
ruJo1igcomtzuH89hDZqXthRhpB9kHWCMGcTywq8aYzKO+lzTSGXTGDVheK4
K6XkC3Wv10UWTYaTlommz4ai0AfH3U9UJA21cnie5Q6EaSsANz7/AFG6g8B2
ipB2awKEl2E5SOpmyb/F5rcKmwtbCJGrIUC2uAXTZU2dJk+aEBis4+DeIx5S
S4GBZDlIRViwFWwngeZokttxQ5GLAdamJSW0nLx/K6p0bxm/79xxtUxegYwj
lJdyTcLUqD5rKp5iUwZa6HZ+tjF1jz5RHQ4YJ38KaV7Jj98L0gwtqzyUwH5O
q/iKbdWtaOd8/66b0HBGGlZrOXeYrU9BIYtAoAN44+X7+zWxQX+AsI1W3e6i
h6yWW5LG0/E4azNyVaaZUKIEtBgIIKnCcBT3aF+j0f3MKrEL23Drrgz+mSNY
pknX5BuOKHu7PRTNFxolZLQmAYuWa7J0pN5og+Dd4PXFg10MLbZl89ifSc29
KLePUpGbMi2xfTPO6ulo+Gc7vzfL3TB1fNSWoO5YqkVGJh6jVK4iwz2ofRfB
esJKpM+TSA+gRbDjRboagKxKFeDDW/POYRDadJXaSTtW409zF3u7ZgzhyQMo
KIQG/Tr1Fme4Hu7BRkBu2pXu9gmnjos659aLLHrgEWwTlFa4tTtPrUpVfyyh
TzvySc3fDocqhbXos8LO8tpir19SHpkfaFeNo3Gu8/5yCreGgmC9SFb+Cb7p
ZM6Im++PHEb3gxSr+EeCn888ngaGPgNshxJY1UFh/C0xgTh3BnuMs65pg+Uz
k0bWexkRLzmKRTdXyw9xRKi0VrJ394V4Mu5do9hxb66u44iXpA8uwHrxIRkg
2ZCVOdcma8vlwPZVG3Uy2gIUhzGVim9f0b/6nzafn8qcNJ1CuDWoKUYJNx65
gylKHWEYX+LrxkQ14zbDrZ3/KIegTR6FeBg6e762WznLGWsjwrJ8LLXVdR/+
809YgNZBR6xPfO0KVzh81oOc0qYsm33WMbFWxhDHOap2xhskoozQcALrUZ8C
jrFJA0RpRuhR1HtUhPSh83XtC+42ZLGkZvEnEplSfN4YeEf31Nmf8nzXResf
dS9KBTYJzSUrALYsxL6f40ifcb78FKNn/nTqDDmzASmf512ApVmmKYplJyMf
ksRaxvQ7iJClRfg8oT9p9mUYE+xAsSPTTEMSawnlFeZKu/snFYBL9j6SfZRS
WPU0YywlZASCZW5bgknPSgEDjwvnj43fAD5oqojM91orRodeWpkOHDf32jkR
OiaTsqMo+v+Z7Xq01UCntc7gNPNXNMlb5b3rqrCywVTf4psfhxvt16OB887b
N2nPeVXhQR2drR+dOXVtSmLdtMs29K8hYTg43gcL+p9+Tsv022WsT5+ndYQv
YcknRlVOERg2LURIPrwS9zDsGhJ8rfdbaWWfkEwnEeaUdOTBlKk1hCdqSYmh
KCmwX4Uh32Hulm18eESpSu0gYXxP3T3QzBdaa+MvFkmmgSXNJolAXxs4assu
BjJMNj1lL+nATqfqOCYEdb9qLhrLquBDu5Ty+h7N+iVZpoZrY1odmG4yCIHe
1x5KGbaLrsY85yyDu3pNeGRDSnCKTdDj/DKFf0wjcz2P5KPoRDINW6WcxmLC
rL3sCES/HxcndhJYbbjoc495dUgj6NCBxOOt6s3C+MXwQufCCcERdJ4nzutz
9F9m2OuiA9JXz3aAlrE9bEDT2Y4sbjfs9k9CdpVXU3Ws4c1Snw7smwCQdEdn
jlWsPuO8roCgDJm9trOoIYh96cxFGE8+nf9A3yAb+cW5LIyeKFujxEZ8GCiM
JQkInnKfDtv9am20uBRMdJhnNDS33yS1Jzjlmvu0UzDBPhSkHnBvOZ+3Ou0h
g19G8e0SVFqHZ7DQdTo1KLaKnDqAxP0VhqhFsfzk27964ow0l/IYJBxwKpNW
Glwr5t+QdI4FyZX67TihOYEeXqCrB8OuRhVAvvsqCWZSJn8fSkgI+f57tsCV
KP88gbtVfOKqubq8yr90ohiDrNn7kFdpSnFJeJknTL8Um74wHEJnxG8WsEI0
6m6QrtVyU6CLE7fc7NFwvcSIUEoGZbqeCvdKJfqt07OQQeWt9234uA4gLtJC
97lKcpA4KRAWVcAI7yF//HH8jdpRdAfjXVNhZwNe94BSiABmdoD4rfhUd1wl
ridNmmfw51Urn9zZq3dnD9Xr2Tr9++o3mXpUHYzaHly/SHUv4Zo39DTWLZ7H
2zod3zzQZldzR+JnXF+FUrufb5cBpVEJ9VVr9BgRW4nV1zkiQAGS47OMrlXv
roTACEJF4+DZ0huj9BkigIXrXnnJ+az3QvjDTnPI6poxzvh+zyvDC+FVDhtN
tHCpbvqnbjrg15MhNEVKLV38JY5sWPGAdCiW8DqS7GOieqNIpS/EDYPcmPuC
JJVgWE2BVHSFnGiazseTtaomn+TUfpSKhuQJMGYc6TOxU20AU9PmQxts+7qc
RUYD5cD1LaILlzLCqymNXY8FHauxZST9jfkf+j12CdP+9a5rWvvXcOoayOdn
SzL+KvGs02ECsARLxNEp7Lf9+Vb7ElmDyjZgRDkA78S5Xgm1nzXGOIKNvRb7
FOm/VmjKsGLqJN50oFtHvVThwSRCilgY4n1QxCWOy6OBSi6Sst8HWQTbmLfZ
WSQj9EZweRbkHCLzKTGGWDQFDbnmiva6EKCNMg80qVrjNQ1khINYoW2jn9De
C+a6eMQSBB7z3UTNGyXK0x2iiney6kpW6m0cY3r5Jo9RJj79hwu2KiKU/s0t
xMxBbhsJnYToanfRdOHiP0b7iSa7M04FM04CePpKgM7ueQr88268Ndx6j6bJ
2+idMilgkyjiANP9OMRSdBpMaUsx4eA20fha9Is0az8CAGGg9sybDGo3zvYK
c40wkqgNl0ma/nmjF214Qvb9WEapk52sXjB3CUSpAvipxe2KrUtV7r+Ivmz8
SEBx00T0NzX2HqWHjPiXD4pU9SmeEsCF4V+K449icAChJzfjccfEpc8cYWVV
yAyeRHng7W+DMUGZt0P09yMajv8j9NPw65ykx42b2VVHZQZBVkWr02mW+6G6
1EmBkijBx8Cs3KGtX9Da1gZ2+qjPPfXyQ2IG6FoPTMrNQ8me9bTqd3LEDnP0
/joGgvy7osOpExRcfJLmeq/4dPDtNxzKnoH6OGf8+5lRktOScd5uLB5vJrim
sz2GUN3jhCLcDoNDSiIcb4xAsKiRwOi+Iv/uDw7O6J8xHxVEKEvyLFuR/NHE
Li/QTr5rlVRay36AiBEZyTGkIpFtihLoKBesIvsKdW5RPS+jfmJFy7sXNuT5
7xArhbP1GWmQu4VGCtp2rOoheOcdITozqd+9b1JcCVMIxMcT0QlutmD+Imf9
GK/S/hMazKb22n+Yd9s6NJPWccsTFLyDPLP18U7FY10mtVhqPpsfvmnfPtWs
R+MkHDbJ8EY1uLPxdH/Z+mzTsOZwouR37Bp8fqoztABlfslZHTTdU7edJmE7
qtrRF6AnJ4H6NXybomy9saWKkmMvrEhYoTJRr+5BV0QIu8FvdVsWtMkS2m/E
UZZt7JzWyxQWRKNdk4aITMJwoOkhu91smEb5KoTQt75TZeobMWFj2bu89gSP
8lHZznzHqa5mijkdmso5saLlfdEXoZ+jUpR+pisuK8lfQfPYPLM6H+2IVs/6
Yqyw5U4K1bkD7mGKGIbi4YsTXCrGxLNUq0vu9b0UdMs4v0iBnp5AuL3vJYsH
pc4sxi7ZUDpmB2u7cNqTqfSPC4Oy+LgBiBdWZh1CVPzmsW9NoVg4L1hXu2xL
2sxdY8+q7uZ1nQcjHLYrvGrM0ZisRKpxdhRMRzky1fxs5MUX4E1xAJiUR+QB
FoH8iVoDfNbfvUVSVQ2UV9QbEKO1Ab8oaBW7E7p/mcO/QR/SUsOATaWB+EDp
odg2ZYr2Y//man+BfSdyOyGkXj9jQwZBni+4B+PgdMtyGJLFKVR5LCvZPHom
fGHHCVkNrUE6pEvHkIR/Ea8WDzgxJIFus7R96rC4ow6YYZ+VEeqN8XzB9vuX
E84tcKtwUkcGmN3+lrTOeC/rgg7idrHLjM2cFKYnqHamU+/9Wt/N/Ga9C9X4
Ok/uBnkPBpNxscNP0XaSefJfuC76ne+/Ps0DKh5uF+z1MVRr25YQy+edp6fh
/johKui0DZCr3qroQVYB6S3177y8v9Jb/foJ62F0MvV2uoGpsSRwMBxOdHv2
WR+WA548LLXLXVrY+jBfnpPngvz9VEQzGe8eTzHLaIduGjDfE4/fRnlzyvzY
ELcjWUkRMbZS/lWhiuPAiUlLH9Q7WBR89+bklCY8/UrKWVp3OPbCOe1cB/dU
I+gu4ZOt8ADCFMIznAVUiVBGxGlhvpt3OUn7IrUhEjJ/REo2Vr/J6aFKrg/o
XwRj3hB//9BiDrEgPJh9IWG2ermdw7o83Rt+1hu9A/L9RQ39reC2vYIxo1xB
3ueXc9gRMgKQgEjx21uadPeoLVV2i7+aEyrLv6tR7BMXyZbF90uFDjaaByn7
tfHuSplJVx1ZCFJHTHNGBSynBvTAeaQjOcVLZ1UVdOfWXE9aH9A81IgGLqbb
vUTzwPbOVgDo5sjHWPghsordNZCHt1Rsn14Sh4XLCI5yfcjyJlnCLWTgBRAr
qwphP3tjxSVesunJWuqqdiRALRJjO89xv34ZzgaI/jLYAoqEM+KvbY2au/4J
dXZbdeBrJtLFXC+/1ufDs3khUZE++bukkJ0we2YuYJxgsOqBfI5konu0JN/a
hUbhz41+NSFbL/+xmdWxLMPZveEONeMJFFumuEUg+/nWdWa874r37Jm2bm4n
WnlhhqSdbKB+iT5JoG+5yHzAFaKlean8O+Y0eH5O8DE0diJDA/W5zN6ADvXk
OQ3Lzh4bH8O2UCzjg1jju72iTMTBHuozb+AWk/OzmXIgbVEL01FxxE/2shi6
XtqhoQADT5vrBkk13X4/ivsFRdYwreUbnmj0IK7K37XyH1p4Fbp1FskWtAHX
D0OVJBXmJ2krn/ssCZO552UCMKEIvHAWUnBHb/AOFmxqkGJPvMLgMI7qYPy2
RuCT1iPsvwF4sW69Sz+opECi/S3ymHjSHcLow/6GzAYO3Apyn0SNzPlEZm2K
2PiHwtk9tycl22sDJVyMQ0Poz4TcGA3GAjfe/3TYgd6appPditCj2MunLgMN
igQLI92SV4+w56DNzS6JP6FqKz2/b97h/3NLF0hghBUGTRG8s5dSg7cVL+v4
u9ErFr3fcCRYpxjkW8Akqk1+4JMOFG5GbY9ZLFaW4xhjDW9pCKoXqQHli7J/
vuq/DX8QwES3WEv4nRtN8Q5itra2IjKKt1bi9wCz4wpbO3d2SuPNUKzeZfez
nckB1Vgc6dwGeEN3c1FTtfW4O2bmjhSfwH1ec6j+1XkolhNiHPfb1gICZIq5
6wcvCWwl4Z5vpEDz/atsa3ka1IHFP7des7fKRErjE18DizT+KMzGRdOSX+lm
mBr7hvCM82vjbchHNjt5U6yfTNAZGqscYMjy+wUS0bJ4mswKUORwTV00QqlY
Spgs4DC754voLZGRkD3EnAnCXujrHB8AwS7f1J767zGC8q7EEFGcVAGdoSnN
yMvIr9g+wJ82hypg44Hr+7esS/WXGdCouWjoboaIshsAsrE2E3G+a+T3/KcC
Fv2F9iJoK50jZ8lcPe30+jTNHNEitH+HxFlTS90P1VMgSvfX73Ian7EKW6Gn
yvr1TVbrv5eAXKrwvr78aGhwHPnkdZKS03KMaALYo63R9XgdtMAMXE4SpRpZ
nof/PvbmIFxZnLUxSYZz8I1V5P295C6TTsHV4Vysu6XufUB8ESjx8X5HlsvW
NpE/EacZd/b3xRzqK6P62G5A4fYbw7COnDZ1aHc4zKcEoscMoP5ORQYuQ9Ym
5o4TM80FSyNVzPPLBrEzTRQCdH9Q8eapGjuFeniP7zgu8p6FRcZdoxz/yehf
zfwfdYGoouvlROrR7bZEOVp13f39T4vGz/jP9po7gQASH/e0uXbfo8k9/nJ7
eth3FOCGcizfuRQdXQ3DP0mHqKAHDr4qDY/hdAe3rkJxNK44/hXWVSjgquOv
yRNVJw+1iWmZ9eDPZ9dmlS+hts8WhlOTUV3eeKoY3gZ9r8xZEfeV88TcB4tr
p8BEEyaYPR6lkBnLFjqjqMee4L9Kt8JBZnp6HBgdtWxtE9hUxKQthtGxv9Py
WMrCQ1qU8vXTbLWGcb8i6FMnetTyMGx42H1UpuzIBzEf9iv6BEjxnnrQCwJ3
6QaFooyQaPhjxyFffeECDGyATWvKOFNIr2QKg8Lc3I4+XGESvm3pWidilWuG
JIw6GBtFT3h7m7FZI/S/xq+iqyE8T8HHKXa3z31+GfdYTOnrR1Vd8bme1Zw0
Ti24Ww9EDy0ZbPIULf/Yp+El+jbD6XMUhGo9OuP9WsPmDgcPOtuTb2L20oCs
o3lIYqEJyqcNQ/boIQD/u4qfhSjp+1G0jE6oVFjfUjL9LRpnbpjvHowLkq9K
4fj44EnV0gRv6xAGZ+1PCVxkvYQXwf2H0ROW8q4cP3PDxaFSuYTNDq5QwcNR
Xw4tD/d/8eborsxePddD6UUBtgukmUnfhFU8y2UV2I6TBaN1o8tlS56TVed4
6oRnPLdotmUI/OphpbVQbHHMgQmuSdu/QYnZ1qWNx+dSSKVccUp5ZAOoPKzW
ImDOnrykiCSEsY8lP3LEMCbaiUhhbwEsaZr/hgYiJSbZoqNYnGQ5hRjAW2QP
ocf2/Z+lUlO1MhNEbiN/JsvAicQVKV41dOTaumXfgwntG3z0GcS569kGp+lZ
xy6MwPORptmaTu+rcwvBDXbWorD2ItEuT6+7YRwVZSYzFSS/S0OXh8kAQA4c
cjfN1N6/gqddMb6qEqDP6jmYLuB+JG0+4JogZorUQJn+lJ3l42MuSadG6Luk
hmSZEpwenp8xCbkclVYlouvyNtxmn1u/q+3fOnavPkHDnZBvXttKqK6s1OlK
Ww6CHCxtPlTPkNr8IpUlc9TzTmdOmsgyzjyWtQFTobgmeOKR1bHwMzLcEf6U
g3ExhFST/SQAxc/0fIEVVYOu1VbfSBd+Rix6njbNad5TvBsVPV4JN5IydHKC
DP0QPFjQlNwtvhboYZEwOl/i74A+Evf4D0UlU10ZqSF08kuB3p705gnoK+G/
aFvaMmQcgA42/kbIIAxh+vJfl1ITaaGT5SYqKL8vhTfaPomm/ygrcy7TTPfM
WovJU7Oov2JobTpN+SoTYDsVGo5sfQEQH09JfRkaCFnjUo/WmE4uvpGlNTzV
ECAeT0A20I1zjjwXbEUL9guvJrmjFITIw21DvCGuFQf44wm85ntCZBUNcNof
Kwm0AoZCt4ERwoXSSS0TztkvHzggGtbbeYT9ecvMFVYB2gi4+R5vujF2ORqH
Zl2Ffe32jMAOowe4oBy0VGHZLQDmQR/HEhbErs6nsexCwZt23xHD7VAvVAa+
PlUsDXGSZc9HgjKbIIc7+EtoNaNiUhYyMpMcfNZD0erBPxkWOp/Hn12JMIVj
1w/io8NXMn57qVrpxsmIXVAZTLFWHt7ZDynUz1OOer1HmFNUddLSkAyRhRcZ
dDMmDOaGLvFZ1ug9cR3PEnP9+hYlcyWBvMtIITt638hMAmrlXEictWmgEO7y
eNPwRBWRvABN6BexI33GnMjuSWscDxCUhn7KrkzJBvZdfV9GSGQ6z4Uj8SAz
OCCeZASEwP7LtIRam/w2eAE8SPBuMUdF4gg0rCKgEXv0w15CudJefCRYWzzO
SHzIahhkEo3mIFq+9aP8YDzzek4PP1jEtoiGnXIB4yIolQ2s+7iMD3LB1Q3F
Q2E3/RJTWx74gZS5jnuP7KksTYy4vX5E6AsdW5ODpEUCdCBTqFJgjE27Sf+g
38WyfzVvTafdFT47yPyVeJzVKypwmJ6eG8VskXg3dW6naeAOpreHyjn7+woY
a6+bEbL/bLts3PP/tH0ZdT59zaKphEA14DqSknbxMAD9g7sx3s1te5yzGWT2
OqlwJvjHJY9IzB92FqSy3+l1j9i5Q/9qD36pTCV4KnUp1sfkOmWY3UHmYsTk
e664D1vzE4dNL43Rgv5F6erRN7SDkSKsgS5+Dc4yCt3dt8wCzOkGydi2CxUE
M6CAU2Zgh8zHoc6MhNgN6qF3/XX3tyCLibRAjYBUzOd02JT9Ft9OTtIlnhBl
6nJ1eOvV+NYX5OsmBpfMV3LQFCPbZLAPDr+uip21eRt/BZOPXNzxzLewWmYQ
UJzkPNHW4zGWcBsothhrQPdW1wN/d+wYHlncJju+4RapmWoi4k4Z7M3aiSUA
AAI1/uDv5C+/6vxsAmGqT/OlvU97O+SNGYk47QXnUbSCDCU1BGSszf9yENtI
qzoSRWjk722wjVxbAB38NgLz5ogNNmEo+8l0WoX3ovsm8oNxKbUEnthsRS0s
bQDXjn+t5LprOZAfRPM5tmTYmblsBBAQJlcrAXMlwofGDdk/6oA92nyngHvZ
ss5lNF4/i95GOjQGOsC7XKCec3FM4ZFv40Xxhfh43e0YK4CqvImtQgyKcAyD
ehFSsBQpfrozg5iHAOlP3XxUEMFy3c9tZetwqnRqsBXGOpQIy+D1xTk7Q2yA
0KJNwqjM5sQShhX2/i7aqUSJC3/oOCTL+nuQyS4A+6Z/Vp9cPshefF5bA8OY
NwruWwTFnxHlX5O3bSonaTK6gfk/ZYeAfpvfOT36W2n0wuy/68WTZf8gNOn6
5phZOu/Hhybb40NCGfnvp3TFIgDa8MaQT2KqXZVYbaMTGI++zbN4UFz5NWcW
uiDRDZqlWAPA5XSLhRXZk8jOe32UDby2cLUF1WgxbGccy08PnzERJqn9jzUf
t1cL2T49AeDz2zVFOSNDb8WYfSWy2Xaq7csedidFWe/zvmGWtp/Xfe1pavJs
8Fr/l6T5pfNgnR7cCe4JWbcfC0sEjrYjaF6IjAtt+oUvHtsXUZ9jP6uISXMW
C0XuvxVcidoVauvuaPCnAR4qQaAiZs/FLRFUfoDKIbxdDWe22tKwK5dhpvPO
b8L57FsVg2nIKUFUpvok+06JRKTyPChU9ttePlt8D5qYMavDywnNZiE4BTdr
cznulz9iU4FgpRl+zQ/tdd1asZy1gMf/XSnKnVS1fI6gpIdKo0/BSZ4cDXvj
AjssUPzWRCPOiobPcs8wxjz9CQg9lAKA7uBN0jFFzC7k4t8LxH7DUSXfhHWC
7Qo4JoAy2Epz1r0CE+Dk4GbJMiFiViIlizaxuIcAtgEqal/web6hssQ+lkiZ
gx5kwacReB+Jgin2z3TVc1rI+DmYTjeJHx5U1tdYBdgjKVHD8K55yd5C5p4H
iczyTea6vhFlYZpFgNH1MEzZuuHNkalpIx0BTbgydJOs26NCpOPahpn/1dZ2
knOVSYelJgw8RArT5jMuwyVFsMO1i7SkiZqOpmncoKshBDQS579ZiWWFG7B5
06nLlz1FFYuAr1odO7bqANOBfMZm5T926LqdEAr8WeM1htzgwZii7WU0tpTr
zN2KHTMJv84gZRpxLIHRIcWhdQuxQR0Qclg4GKq6iO8V3Gjt6dJOb6QKCYRf
5QfNEgn1+COZ5ZDIwohDT1tlQQkC18vcPOsgvMQx5KLGxnWKtIhk+p+Yb6k4
/sRZMbEnSNr+cziq/RCAO80mPPASYododw0fDKoQbFDSVVB/t+PyS0ZO8s2m
zruxk+3BeleYc+54CbfjxKgRB9p+79zEw64M3MqeYFG2K2O4IMmcBYxpF9M5
5qwrheh5ILMkNmvrp4udyx0AfU36aOARUbjJ8r6JO3YpkUyAAXKTcXJi2rh3
hjF1LNGXpxtxbuDD8SPDGNl6BTryHqOqYxQlYMtZwPiOtSJ0JFWy6tIpWdAS
O8tkGTwglA0IVg35jE90e9cPOS9Ojg8tQaui+1/JWUnF7Z52CJ+giBknahFH
kcTOFA+ThROhNYMOgma8Gk0za0hG4dOBIbm7WjY1oQEhxazbG+9EeDTm2cRk
uqhJOqYbi2fQgQ42x/8Z7EJMv2JAkKI2wD2opO8VUOOXsAct/ldLGDwd5UVt
KTsqawqFOHu0g1KJ2JlvXDXkuMLPCY/PPy/XOiSIgJ3vPy+UUrYcslpeZMeP
8PF3Fb5tGsq+bR3GcNFfb+OQSDjz+sSlL+WFo4l3AGTkgd7zxYPzGpHbCrsv
WX69mCNC1f9fgMHkFa8fKBzW/aFQB254677Mnjc87wHAQb5pkERHTrEWrkMu
vGjxEP2qxDzYTL+rj1oY30TYavuy2unmZJA0TaHwd6l4namIIt3UTFM6nzFj
F5l4OOrkIktyT7WcMeyh3CJogps9Zy+avtheukNIIz8YVG//2spLvYEF5hOx
FP/oSsXZm1Hw4MMjcLrE2+FCh6Al6WjBegEkjA8gdyOtfbp+M/xE6BzccK0k
6OARyTUCC3XmhmQ2SE7JuYUKp46DKuW0xZo3GeJdPjobwj2F19ExnrNrdIBU
2jePgfHVD3JJjvz4yscQKEj9dpKcS5DsR7amijnSRb9b9nkntf229D3OgS5e
OUtz9H0mD1jebF3/Ii1eSOxoujVEPA3x4753GAl54tHwBa2TC08D/sllfF8j
8ZaXgHj9eneyf300Io0Pkm1NcOR7VVvKwVGSbz1cokT+zQqBkVp36me1ggNf
MIUGhDA5oPh/It7og/i9WFfRClUXyd8CTjvVdHcQVMOpR2GZpJ6Fzf4bnZgR
XNJ7QAhcsYBpr/wly7PxyIe6Dm2Dt86wpa/lgT5sl10t9f1ld8GrC8qtg1it
rnwWC6ZOecRNp421H+96u7BMy4HWOs+NjZ28tl24VUD6B53BtMBCOFc9bkz0
zJnlShb1CWFirL3M19Ag2PrO5UYYwRWAccuOpmVip2booUBT5YyXy9ggrgIt
Y9H5rOEi+Pv2AsGXar5jD++jT4oY75dulPMJZKHTqNkwjJm7OcL2kRKR7wFN
+RizWWIBNQDUgv3+nDgE7hy1H4Nwc2BXk8uUJnfSODVPdFs8sCL02l4Tes/F
ExXiMSV++mzUOtQrNtro8Tq/OjGeI1/MuBlzkxn059ICw2hn6zESGXqW3fbK
s7i53TJKlRcdBr+XogeohJIteD3wQ3+n3M0smkt/1Crw4wycTYxQdmDs2JDW
9gNJl0XdHfhEQTOYM4Do5ELqDpG/gicW/vasRTAncyMnd7cZ5KbZzDCwIDCl
1aXqlbaZIizbX32SxVnqZofMJj6wVV0fdYfNgTxgvtppnneBs3R/Alc2GtJc
XSqwZc8WnkAQx0D8ObOWtKUAKDDCuPYA8Dn+KQQjwdtJMST4zPUhXrA9EyoN
bmxHngTptvzHQL/WlsBFcU65Fg1oh4yUh7sWqIV4IKGHpVkw8EcGXJ+bV6pF
JEVXApldcGkaAZfYyaPJs06YKJtmcModbD11aqo254UG73BUYc5QGLJ+60O/
+krAYjxJavsDmSkPEbf7N0xSX8IdRIb5WMQWy5SZU4u6RDmXCX7mLZVgDHSp
YrAiPOwVycCzNb27QgmJ/7CUX7LoSE5WtjSGKEUtbmDpEDsvkq0lSuAtDuG2
dz59McDcvhUmZZIW7VBIkD6I9SEoH2UxOe6SZMXiw6GXgfsc/iC5wmFMWMkV
gsyWzyzRnCaxi7hx/6nURGHrPWQhPBzYQUIMH1RF63lO219xoK6OyLYdnOvs
85DtmgY4yyW9jDKX1xLmuxMl4D+SMo8B3qwOQKoweNaCVRto4x9ez+pyirFk
PWxg5qcBwp1s6sfPvBGpM5Csfyvy2btv605zxJv40tvKKICfJI1WL4W7LHy2
RoZn6R1ZTFGvEeggNDjtJrQihktsPpiLpFqU6U2hlBSh2ypgv0E/smtv6YzF
rYBpgeg4YYp89CBK7u92kga7xnjscOwIuDuTNvxRzvnC9v6KnmcUP7igc1y3
qH0jT+2MQsWcbNOSLwBXwdQ4V9XIZkDCe0zjy8h/2fm/JFT9jO4YTUMOTHsq
u97aMHW7etn8dcDhwXUIiAGnYrY1mzZ7IoznDRM/f2VsvRystAzvBeolwW85
/2Rg/S+LUAbAhaHJWmxpVtKth8ywim8x1UkOtJeikiMm6vc71n3MQVkHpqzd
wHEHARk63n/TNeelb6WheAoO2KTX2++VHi2xIsg7Y9eADcHt23QgbgpOuc1Z
LiXcpyAL9rfZyjTI8EQv8CuIIfJllLalhF4ru+rlzjsmnB1HFp8Mt7qJG83p
H1Xg8eBiDLzp4nQSflyYGgK/AUgTc1egFXxiQ8sZvk5Dlqvu31+CpLrn3A3m
48MMgIeH9sAK3+lQtpi0EBO744Uu08EbcCCPEWi7s1gIpMjYMD1OUSsilIqF
JdQAZ3tSVaksjLbZujjnmpNontrNDKQDNCDmPtfgSZ4YjH8cfdv154ZTI0aK
0jllbl1Ai3hEws4jgVB1c3umng/r91gvT5Sms0G/SsHhsnwiMVsP98mMy3Lx
0/c6vfM6h+OohHGxl3mm+QYoC/icOVbkxi4enaGtEkNBlRyZTjHvEn7nwkF5
XRCcxmgeliEVoDXMHznizSDZjZx6Y+GADaZrsDFVQ6fgzFOR9smgzYpjWa8g
aaqpWyIi6qpAqQI2JEiadxmsUVcoc2gkM8UB0o7QFoBFHLTDNsPGA9A+Uq1Q
uyxe0AtIeYFYy0SPveGPcLHUU0ie2d+aBsLWiq5OZI2trHcQ0FoYEL6TAT/3
Irs+Nc8SWFBsom9cF+7i4Kh1PLHaPjhPhVBj/b4SdEXYPCBWXtAjjp76ttu5
NlxBkbCyJWVqSDp8QoPUZ0lotkCVvF1xo6g4CNi3HtGIBciX+pgWkPCuxpS+
Yy7c2h6+7bCQdYwbHzZljS9SKrDc/xrkNVOOUzgGs+IVXQgdECDq0Rg5K6Fb
oDnddnOS8A1NV4UUbg6IuK3KUuJtNfuXZnW1NZ50FdyZcVIY8VTJUEyHjsW+
4XSg9kvsHkwB7esN61YgCN6FIvOGLLPStpBpS/p1rhDTZ9QONjYTcibdXjfS
rbs7haxjOwohjuiwHtT6Ol85IZhUgWNkrZLSNn2oogegwPRsuuhvyUrMbMPS
o/yRPvYmFk2p8v1xM4h1vSBc7cyLHv1fgQdtdAPeILdDr55knl/KRiPrVv99
u8MQh//Msa432OGwZM2c8gAK1YiAptpUj3L603wsUfWyXJwelD6e/HiIZTQh
NgrZgO7llnWuW2OPktzxiz3JbO/26hx+BDRgvYALg+XqinGz4OypanV8TSle
twA+w5b0y4ARb6E07IYQCLaKCmDPHt9D1JVIbJwi7eAQTIdKvO+ypajitDYy
0MUskNiVZt/G/aTwwCnqv5muIHbWLUM2bPw3RnY89TiZaGwXjcSHZwCy3jp0
1KUGPwcegaI9ac+0LkX8Ic9+UFHLngX8uYBMpcj6Y5TIjlJtK3JbGLTRM/gi
J5bUhuZgOdmhukn5TKkI6p0yHzqbvlfn+KTdqEv5xKxJxlK0WTXhhyaP9/VW
05p31/VNaxBVCgrq2b9INGVXLhtn1/nRT1lFw6nlPpBOXQemEX2Wv6zBBcS5
7RWqA8yzoXyaHSx+WW7lQbq3j56wP9rUkppfNi0Dh1pyMQF6CA6Kq2t5tHrV
szTECkfcbFxubqFa4f+WVG+JpKoFTLQMgZgi1pHfLBMClItpGypQ/olaNMhd
DeL9sqGUPZM99GUMwGzRPlrH/84Cf9DkpHKzmGc/Q3Is/7QimZPpDZhupNsa
f3htFmFYeZH5xe6KJurkZkR6Ndkl6jJ204gYFVMT9x85O79fOq+gjd76juU/
u6yACLlFeA6mJTa7CSwyTgDfHBmdNixEgNh9rRB9SDyratOt9UR1T4l4BR7I
4spNw6Q5+h4AzVVMS8ulvfLZRISufEW7D+s33fNzgaBUrSgHygtN0GF2LOh2
l3XftPMIdiSMy/r/mii1fxhApeqvPs45+/LU645wgCeCz3YwOG7St0u8e6Vr
0kR3uSUwGykhKmtR6YZ2P1S24Ww2s09N8V1OYc+OmmbCVVbLX0FKAU/aH1rl
HBfja0y/slrGzxaVO6uvAW2OfMFIGu0bTZwjkzyaTg5xeS+PP+YGJfXi6jem
40WCzaF7pjwmiCZm6Nyv2nnJQBMguBoTwvqh5+Fai9Gxderlr1G2vv41Ew7w
ezpPe6G7TlRDvCCfTHb8kolJa5kg+wDyjNWuBQlzglO+ABF1fNF7ofAEMlW1
VS9rq0djkv/mGzQaH0BTHpGPn0Wo0Mg7W7hWpk1hTOGl69/iREJpF14GpoAE
vMOO5oC8vWl+9FYLY4iIUanpPHra4at76fpDFr6/cnuu8b8yTKMBRsY/yI/F
TXMYLr5K1G+TVLZeBelwX+nBgh9AhY6dQDlSHWxHAkvuFCrkyY3ECP+3akBD
qpHkDIks/+aLcUF6oMHYQK8wUhV/GTkxaCbfBIOdOkT7kOKvNW0CXzMg7bZi
Rqaz5Z7vdwSXOENCXj14evezyXj3QMxAtLHxMnZZnXJAPPEawbTbiOHXFC65
PwULne/Do2zLFmvlkDXKRu6gnrs8Ai2KVq5Seg4dOA6GlsfjFnEoqqoHLQIL
CFf8thbqepjXvKOVK25y7BFBia/qZn62Bi96RNqzDZxBw13w1H89Yp00nHuS
UQV85nJCs6iQY/aOx0kiHxZLgB4nxiPm9aDUY1KWKCzLWUs+Uv4tKJYv+20W
NBpi+8ZHL18Nuc+XOo0RVQg9g4jNV2Bpbd8IcVD4n5y7cOblaboTGTHmJews
sOi7zCiDzYwfbUcEryjNioLIz4G57rUNf4eNZbkB8gIlcN+O0N33+USHuBzI
9xnIS6EkWpAGX499gMDjcvMSrLXvBwOMA0OUKTQr1wzfxTKa/9Eqo05D0yFE
VXAOLysAyHWsEPWMckQkKUjY5Q7uajrGZsYnXc62WuTmK9mDUogriM4jv/vt
wFQiET9szl7rV/5xF7osm7SMLXFiVCdb9nJBAQCizM8Wc70jUml1+YHp//fX
m64G/SuRZNtH0bq4d8Bm8TKdu4Tp/jJsng0XHXx47UxgBX7eKc14753ypps3
Ftl3m5zCyS7JFJ0pV4PMvDbP/PZJqrEAun18+T59lb0gu7PASIq1rw5xcT+P
kO56+MeEoo2RYnM52axzn6P+CzVeq6HqhFaIvQdvVYFvzEU0aBy7y4EM1iIL
qdqxMCsi/2AC64wEFu5GIiDQsBmK7PmL7Ey0YCTb7aZljdkO5nNfxIi31eoD
cNq0Z2ozzKJGtD1+acpliViExRgusjwh1OfLmj8y2szFIvfyBIzlRLSJ7pKm
dNk+4HATkpF7O46AHv+TEmntx+kGYIYW1eOVLjX6x4CVnWW+Pjpwgbpk4Oea
rJq5n4fOfrntT1hQGSQN1MOokCI7AW4jlPskyAxo6Xd+eSiph9fL8aZgdQxD
jxrZVFLQjPBIsGU7YZCgTMEcUjwmj6pSbFiCUntibvW4CRGCdpEwWy+WNRTQ
mEKCzJBEMZ0uUKgwPsnHJV0+QCWJOz/X9YPint6VdoSbFl4vQ433Gti+tr8G
b7HhwK29Pt/XbdUpLPM30CKkB2QcuTZlSc57xXDha8Zy0YF/yAvIn6eFP1Qf
H8782GCAe9lYY/AYehyUH/zbSJDInVmE45K95uV197zxpyzVIHuuIqjeYPHV
2RQnTqIJxkdNQ+uvXmhfimI5ioDDGUgvkW3Uhw7h0fe2B4+cEHL28aOFBwdk
oMEeKdZbnJ5AZowOyMCrW2Xv95uaPvgsWuOxG+oXK8BJDlQ5ZT4q/QZPFSor
OHrGn7/APTMV2xi0X7v7uh0flwwN2e4FExegXF/EtJYxL86XfM83Fy1vIT2x
Aoafci0DUXcUkdV7muiXzF8687HFbKvpixAPbcE4UivsUAyQKVGjyJc1ccPt
JcbPgtJyZ+Yj2qMfga69vx6h88VPdw6W4FrK8ABDgTuru8JwEjrCoI8pOD2F
m6MZhYPBu2yHk74PIkzMP9AGyWrQdceSoZoYqc1OrgMOrYsr44bFskkPu/Fm
xxxUOehXOHd/AKzgct1CjeXBms+EuI43/tjW1EOORxA/TawpYOsgOhXmiiN9
mllOGPFnzIBbEFhC5w78wUGPzpK95MtvI52Zw8d/MiRTfBFhwI/h7ePshXIo
b2qipZLSGxlrfiYX8/qeTEXAHbIcpicl1fQewPJEVYV9LIVzbznxCUuJOhmK
3GNDSm3iRLyXiQrknuHTsrJm9k6Uy+bHBiJEeePKOmf1kYAlqYbwzbIXeCXk
u+YoL6YKYCFUUBOO5NeD6W1/qLCJwsNG8O289/Fl6x2Ev/LAegavisYyclFX
VY8NwYUp/grwHx/h74jEO0d8zyN8USk4sLJhUgFFQUOeJQ7N2E+m9EkhU6ga
jmpfFeHssxN1FORAy486Bjo71YX6au4xA0bgKkrYXgBUvcE0JCkaMncbku8z
i0XrSD1RZC4T+MzK74n6vegTiR3W6X9eJaEYYOklbW/IcER/XpUHlpv+UaQG
MPc1sksZzE7jkWXeRMHmes9NAeuJJs1O7hXNkWvdCHodh+u40ct9+HRVFpYY
1lVwuSgUR5Md1VfFzNYVz9+2vy8QGXCP4YDXJBpfZftHJBJ99Pvf5n75/hqq
Ocjf+q/4zYxE0Ok/KnWpP2+kWVDTB+F1fzLZsBGt4zGqC9DqmURoTJmoUjPz
CHfHnyHJC/ljO+Yi1CnvYD84UWC4766lyjkVuQ4eGHMN7ZtYIJaleuJgWeL1
nnyTSH2eYx8FJglIH93hQ6WGfkMPcc7S3Rh+BQA0yeW7wBRmiXmj8GO9gMd0
UxP2bjpmZy1Z/HVHmzFRChLJmgl4vqoC+sn0Ch17jLHYfGabKcUnK3Og4IYG
/votQQYcX0dhmjdSf7deaGXgnywh1ND57ksl8C+aeBt6fjgVvMMdt2/iJTDk
SEi5+qLOy1GMGaNC9kYmu98xnAusveklZ5ex8LGfA58X2jMHxH/KN9y3YHhP
LdUagm3uIlLmXsVGb+P26jW028NCUU8Y0Nc3x2ZqkpElelXiXs0iUWg0CYEo
LwR3Evxc13HJgGh4mubfxi8YWPMdpVKEO+dJXPwMDUUtrG114N5NH9enqZNU
TEUb4maQHtE9HdfT3x/0VRJkETwN7/BnzS/TRj3zwyZxYM8qd8/k79T1tdI6
YGdxF3vHzJMZ6oqUtkL9fvgQFu9yAoxh20jj2MBD0CyaAhUvQenM9DTeLaFB
ImANn7XsKq056rEPLPyvKjRfx9tfc/3ujwvLACJj081CVrFvl5TuBBz2+3Bo
IQn5jF+BlPmLvA5Ah8yibOtLAHy8e/QQH8Uxj0EbzR1KCMzaJmo+o8z1QeoC
sZ7j6b6Dj39vRWW40ZWMZ1GXJE3KEdiRJ/K8hXcs8eRie4lRhA1yUPbi3V/t
xQY99dV5n6rEFeovHznuLBWr17npBA+zUSgsLZMWl/onIoacYpCkOkAWW1DH
2tf696en8WkiuerXV3+Z0pJF/tTx23rfyWwbHLC/wtU82JnGWiaX2OnOnSIi
tnYxLZPClxm1WcRXQBgq9BCYrIJlAw9Dl+FcKwlDH5Fck83iNn/ZWZioasYC
roKqiuj4ZW4QfLAjJv/W/69ua0/jX/RHWhr5pB99nm7BmUZYt9EeW8SLCrXy
5rBLV8NGf3KNRsScv2coyOLiPM5oXxbu1KVjUAEzlg3qNfbb5bhojzYWubiN
hjso6/XUpu+HuUUrPPRbEQZp3OlHIf358MUsqCj7QR0J962uCtZEYbWhoJKr
fGLLvOvOOOAgUerJIAPqMfL1NCUn5aEQbcdZoDwBy8Dc2ok9llL+V9KQf+Mp
6Ild6TRxSY8D30SFhXBTLpDDgRUHnbWl+QHk+rvhFdG+SdROuI+Q0702DCdB
cNfiLphoOrQCcnK4ZpxTGgVMOfahYc37kpWZ9rozTjmH20TViUUc5dyywnVQ
/dmrk1DlbyKLbi6swsCUtDpfpwaVKjYHQ6PN7vOAH9LYmlAW02TOW0Pjf1sR
QsdUMGzLar4pF4Tgi8SagEBbf+yTyM8RgMRzCHD3G/C9Dw0jHIma0FajzW7M
BmzOsGGW+WZzre06AaRfICaZgEKzUxNGQDwgpTIryBzvMQ1PshmPen7pB91r
uPoP7ahX3ZjSTwwplt0qn8m7Q2UebOJ5Smz+DovZzV04al6CpXDv2GxEeGja
cJk/ne8Z9zID+NFhj6PfLZTuBe/HsqpRKslJ/TB4P3uUJF4Wc67xdZv+audW
THZvZK67JH94yJYFJRyS92ekfy0J+Z90CESz6K/qDcQf/RqYPjHfT5HT4xxU
2RkoBUtagESJAMtDonrthTQakTEy+V8DA8jqBERH2I1MK2EGnerJjzmE+3OI
dYyZAJdYUYICvCRw6o2Dz56z/0fD5kgP4p9NPTtXfQ+aEJvmXzcfLJOZkvja
ZbGDUNYIOS514CR7QneGj9INqVYQqqmRZomGkjhWFndHB6k3cElFc+JTKfoq
Ih5YbSlzG83xQjfhsPP3PsYW3s9PMJQrXtey0ERvvdSGe4MM57SfFcIdCtGa
FJoMUa1fTHzhoGbSnu4uMyICZ7EC842Sn+Rf29bBGBCP4vi5Oa3ufPHfcpDO
MUU1NDovehxvma/MKOOLDvjb2yPgD3Gm767nQKkHOUZY0FLeZ+AG4iod4v/d
ju1Dr+MTuF2h/93uI17UWChLDhzER17H3VaK8J4fzHFD3V1X0wGlKYMAs91w
RrL1MOwOsbi17iK5Bd1sFaWSRrz3oQNj65OnGFYKWijFevYDVV0RFI5n6vSu
2CBodBdLzI+zhQbAzgowcN3+Era898tXy0yFvs4qbYfFd7EfWhzMGIlO2lwh
GqQAZQDiAicVObw2WudjQmFAGjQeZS9guaZUirKGWJrn4w1NThLQbwyPPIrU
YkiPPo1qzTiQWzP9fPnYF6P4TEuGAfEvGfQLOMDN3HEbkdMS3l4Axi/41LRD
RSUSITurdcQUpuSKZyhyimIWocbD9j8mst8b4F+NA07nZqf3EWEHDGd6gv32
P7AB789QRvo26/K5LD69CUv70sU/SaLecCF4vpnANndyvTRSN/YgqSAsBkuR
yY6ggCyKDGfTuf32C1kds8D7+MZtlp13m0j+5uGmrvXZiJ2PynA9wy//4fKd
LD+Onu4Xm4TBS4A/6lHCI+CZ8OW8xJLF+Fcom0Ut3dGUC5Llbd8JNnuFTKNF
+KUHTQu8yIcTZnRVJycx0eZeUh6+x8A0QafXn+I174hDs+BZSdXUDJv17RcQ
Y1huVChiVxokMGhd1UhsTSh98J5vN9fzOZ2yivnPBQsgfH+sQn1qDd3T6pDJ
LW/hqWcSz4VOk229J4jU+YSwA+mBuR6zDsF/zi9EQGG9ZXHRGxs8K12hJjCG
rglrNAtRpYFpf4yQ+AWbhjEYAScp6BX+my0e8qsw1vLpqayBVSEgbBp/kyBs
W4AIlhAAGTBockC61wpG0nD92VJyyYBreG2JWbZOwgPYRPE7ifGIH8uTPdHW
oMuWTbKidIK6Sq7HTfDtr7f9WuTm4DbmWEKS5o6PsOFwrIjgE1IKROt9CFan
XAOK3svo+7w62rYA76z1c0KiEy2FwnxDB3/4FF/g/hlOFO+PC/t3KEeQGjTZ
rSSTbmNkfgWPr3H1LYTHhimRZWErdbNRx6QQKvfPYQZp5YPiyM3CXW3sOhd4
62W+21KgABrWnWN1vyQYYGCoE/3B4bWpfQ7/lFspRU/uCeypBv3M4cqGFYsK
zWnmqFXHkg+2OelhK3l4nMUcrzNGLeUkfFycX1smgsnM+vRKOfseyV2ulpa5
XAOYFHM9EQwobzFIyaNVOIC4A/PGMMwd8koz0wcHHzLDFKMTRIbLcgh35uTM
tc4zRzk0APqzx1hUOfGEYoB1EYoPS/RmWqK1omwS0sI2a3iXl4Qxy3UIQgLs
nfCOPEd6xkXTsoHWGBKd5mbbHeJA8RMTzuUm0Y1Q1W84WIW78yDxGIS0Xows
vCpB1NZJPoA49CCS+XXZ2NzaHDWgAHKLw9aSCR0gF6MOSS3bfaGdrfmwiKcj
8VDE9fOOFXleGGctapMdNKZunZ18eW7Fmsl8s8hFcY4os5xXXUjpkNuw63xY
GvQJ1wKqhypMTHvpon7iVUB8R+FyklL6LcdxxuwpeNp9+6TA0Z2dIvTqEvuH
ih4Nv29qP1Mc/irhU4lkzdHcwdp77lKF/kmkycY4GK2zE6Uz22tJgZg53B8I
gCbtjT/VnOYPc/fveUuSnkUkmeg3Sk1tyvKnLOLnoYv2OdUZ8YPCmT049EUS
J6KziLbJm6qcaUQSW2URn0/AGVxmVlTGVS7+PclQcHYOU+JOyyG3bB7IQorR
rQ3ROovhTWzlhWsHrixDwNb3yLjeB2nn18Qj2/vDtZxCI8O5Cqc17ykLGzT1
9Bvj8bxL+Hjw/K2O72KvxE1Ozj9JXyi0Sqewm6JVTgJhjciKjzcKOCCvLLLz
nDjWQDwPMaccb9xKDsBtEgEh+RXINoXNIuMUe452sW2VJJjT/5poMH6v0eux
MlzayIGHGOq3l/0eq04IlEhKwoirLPu4Y0eElLh+2rclZMar5aX8BbNMSncr
WSc/Q/7d0Dz2RSPfaoCY/mPReIlrBKGBuTTibJFbxKcbuc7tGsrmZrMH40/K
cgPjFeD3Yf+bWjSt/f9V2GJg/HBT9iY/mE+1d/UlPlEyA+/lG2pupdVT8mF1
vmbeZuXKuTdpifZj3dO8ooDs/wBb5I6yimuvne/iUBCkdg39xELwOYRDzXrb
ElXsia6++kC2XwJJfQWN47wVCwIHyQ9WcM8cKDgYQOj9ggh0Go/66KeBjvsV
teUZpcQuMgBJGlevpso0ocT4sUdPnNupK1OjotE5QrhEcDZXGxIshE70U5Kz
PgYvno3GX1fEGZmvIoBtnJMzwGj9WGeOACC5MNPdcKdsOFiLC4TJdJGzjCkQ
PtWoxg70i59ssxIqRgwE6mlslK0mTb57HCWdfSUEHh69ZEqFAtKs1FhhYZec
+SHvpW4Zewa4N8MQpcdUMM+qJQ2VLtRAPFOFTEAWvf8eRRocCrdSweJS1ZNK
OLVGJZmo0YLhcKIQezMcNrZF+q2zmLzgv5RexfQ81u+bknyq5Mo9znA8/9MR
FKNcauYFU3Y6jwFU3yIFueOdKEYIbfzz6fPpMJkVmy5q5azJkLmOlJoLSsck
35ui3M6V0JCf3zUSK4RqhqmFkuwT+hnrWQXz4UdLu65jUM4/tsxb6kLEtbxY
uRs6r18rOSa02+xcVvRYTIoI9IVdLjYS3dmySN+pJinssxGKvg5caND+57FB
SKvURQO5xiXTCkzdTwa/+9BidSj5R6/6TnSVeUo/vbsS4zCX0OEThFNqlhg5
Pk7BiUrGxflHdgAa8F6DZBgHWaKSPUO5nN0DRSp3seOMlz/WLcW3OAXh53jE
6qM4QxHXsMIiharKkprFrGtdYMDoF2GhHZFZUKo1ie8aT+oBafAL5mR5rcjm
s8ySJ3WGUTeYbSVn22vEko4OL/ZsRyEohKXB4eMbpQolgiyGg6mFwgHrc7Db
CzdqEjx1sWYfBRNE9PSUhVrk0/wCbceN4SVxtauswyLND7YR/YifgSeZm9wk
CXBUK0NxedSB0wKKR6Vjs850v15ARHkz9eLBWFi3yEQMHsA0SUouHpiSgAey
zomRe8m7sXDtpo0vAks5CKQSXiUHa2BbXXuchzdUCRH4X2XvyQFrmKiFrMjH
caq1SPYXQs2o+BFQs7JLQLiM9LVB58NeN87xQXFMUCLZGhkNXyFRj5HRaboO
CacP3Di6uV1L0ivYfNFNJ6bjczD7HYtZjktxkDyKvpaVIe5uLFAj/OfdHAtn
6alDCnsgT1cckPeQMuxNd4DMsH7yuvjabUWivlt95qGVFW/A7gGxZaAZVV1V
tqUenFX8l+MAeTMU1heyTQ45HkzaWCv9FyOwe0XQlSfeByF+Gdtg9PyxbhCT
KXICpQIf48rZFcwn5dnWdG/R4KUXgGuc2pcO6Chg+YKa4f3aYIVV1nZ6qF41
k6hV1Kg5ktKqQcatBSOMr5zmNJl9p/dolN1e7aZtPPZnwq1r16Di6Yu6LB3a
HZQ3acmZRV56bsxpxqX8T8c9NLxYXkLvwK4KrvqkEtSoTnFtbyr2/nmhi+cM
fw5jfpbABm/QYjoj5hrRNQtj/1B9mNwqSxWYD8waSPwaQkXWF9Ssy9g2Y/89
e/KjAhV5i9PyMV0YTqOSmTAymwW5lLdKvcnv8MuzOw9Ow2cHbLVaaLbR8jQr
u5G1NqbRBblWM3Ja5pXZZGWZbnjKoP28hykqldGUMukATgHtTMvIyXhi5HjY
n7rGqbtas6yaWuCFtheKQxmQE3kaCxr25q92eoyyQF4vq73yfilADhAnJi8I
X3663Ob88Ofe28tQvVXW1dn5PWTgCz6HshO05K9voSW4ODFl72aXpQvpUJeK
OnmdpN3W6r5DcCup8/mGlrFCzmSuZj58loImuTkulA/XAVdMkQ3/Vn3vtb8k
gSCGqOmrmz+FKG8F/Onrgc98wGSjtz2QFiPorbT8vhqCjP0UTMxlnxYI6R4S
VgM0zsGzalpptqbPfT/ZHNbcHQjJPrE24WCIWcWVy2mMXBBr22Rp2wTz5zCB
zbp1hjKx3d6RDkCSV3GkMEh1L899mDSEcKcRvF+bSW6+cPuPrTRoGcUknEFC
EJXHldqHE9vsRCEw0Tn6Ah+zQ5feaIy2MeTnQax3Hle45EK4SZJANr0eYChO
ZZSYpzNqTs43U0+8THyq9tUu0pI7gImNMzF3Kurp/sOhsq9Xur+nD0s0WMp/
7mBncD6TeB5WiyN1LQSTHHKqSNbZwe6mmvxreWSwsWHKTfFyH7fMAdW8xS0l
dKrsQXzTXMVgNVkHZu2Pxx1W7kjpHd6LOZbxjnJZ2jL1fXBpAuaLHloTe8tc
pU5RhqeWc2fKNHBgNeAFFhm4L67IlWutR4RXg4N4FP7xE5XxNl78yb7ogS6v
GSEtbVPAFG1Q+ZspV8rGxuJSdmkm+BBX6+Xmfo32mXVpzTLz9JVLLF4/leNV
EEn8LRwngg+zciPOkhmGh9wNyaOcAuSTM0V840rD6wQmzQ0aqc1tkNa1WDgr
i7WrxtVBS9vX1KRBq9Y8ug9OxYxiJ47Ynzb5EIpxAsdxFVHIVohxutCDBeCT
hbPrrUj+0sEqF0NCeQgw3QLnKROmEVk6PR9/LnGdIMYOHV4mndmOCv48YveY
pV4sVX7QM5EUJuIkVwKQ+nI/aiwpSrJlGgSjzKEhwwMiv95fYgOVb/+EPZlO
BvSJ6ATXieHdSYxh6fuanBiwRCDzN2h6OBz887VvLbWCsC/D63Ol9oAmTlWn
1iRipPDZhYCxbDNj2IUxeGrnY0xFEWqSGQUaBHwixNO7u36C6NaU5BLNLXrP
HF0PPy3422YR6EqOCn2moFP2yb3DrQeQLAsYm3B8fEJb0Lr5YTo/heJs+vRn
YIQb97n+2Esvm296MMylNupz9Hk8vcTQIaE/x6fLxIwy8UklMkuqXDlhXj54
BO7WqwYwbVrQcmz7BMRATsi7JGlTd2aXviDeskhb04dRgwwM2OmNvcQCgxr6
vkkvhUbGboZOzBJac2RX5k0PixzBrT9Ou2WehZZviq9Q2XyqnbNmBkKNMmyE
9akZrzUL0/qiF3IzF4YidoIFg5HNs4o4JlQcf1ppALqU57d/RtmCPUHTX5J7
c2V9wGmr8YZ818sSL6Ni7erByahcAABuVlKcYoubrgoYQWYQL0rHUpditFEJ
u2G88mvxk9wFzxw8jjQFReo/UdewQI3j2OsK8Wk1sc+loTjy6U1IHsJZgg4t
yPqy4dpAUTCxumwuzJES1d04Do8AGbE0dkR1/4YheVISCZTQ06Tw54SDUrj7
f1EvaRcuG2S1Set13bbMme5JUZZOlayL9SgTsyJ/rPEsblsYrrK0epDQaM9K
+q1/6HFLuQ8f2cZV6fBqIL5S+96ue7eZocWs+U9P3ixB7xCnKsWCxtErbSUl
mbj1m4NXcKJnkQ1lkqxTdS0nE1Q5lqerBdyBkON5jR8oMMUpamItwvrtiYIj
M3FxkN/0QS3vNqGRfDd+dGUBNu/o+I8HLNTdYI6ZiQE2eSdvi9OLxHBprAyf
BL5NX0wbFE+cUP0ZooAGMDiUekluEXIxAvQSQn9VDx+zbz6Q92F+QQrvQuFH
8bQNa0YN/tiBWd43jjyVxaEX1QjmvtjYgx2V0uJa7acpXwX0QaUfx1HbWVm4
plaChSbLRK5VpsiP93XyvcAca2K+Av+yCfDJvaHDUL/aWvoIHaO8EQhY4n5Y
IwZgpmSauQ7dwVxFI7NAF0gwsbWlx9ZKINRI4S1tOXfbRSQ4X/2vT349+1PA
y69+kA4zPZ7xcKlydfGgoLvgXsl0iuXlJn9/iyRJqvnbDgEcT2agzrIgcJhi
jEUSud5x59t/geN6G0mzueS62JThtE/DIxUiAEz87LQjN8pYT2kb8A21WIZC
DxKtKdyRG3infSeyc07OnidF25LNE2bT32DUzpbr3llNJw6OL756ZnLSY6/W
TYzP7DIkciu8yITaP57B4UGGXmzTHgkYYEfHtVfqholGSFaVo0bsu8C75Py6
JSSEAbU3H04+ef90KtF++5oETcE4otMkIty2L+zslTmRO7o3IYVRs6971znR
hhO+ptuPUedpi9dHKw9JpSQ/0Vf8vyVCjAhbuLH/Wk51DEUi9uaAzV/Cjq6+
nm06NSAMD4Hxng/M44NnlO65EXVeMmQPJhzamvVg+k9c8H5U+c6Iur8wGyBy
tuyn9240NRSxZPFLWCLhxDfpj+yUO0p3++ivdbRrfjXu2sqU/D/QkxYYvfkB
YqsrKJwELEDGJwX0f5aOEIaE0HoVgrd76ABsDW5PqDFcg9twE/Ab5c3kACZi
eE9dQhlaazuW+qPB1P0sRMBed801xPB/99re+vrEsb3jFgzX8AsUpJXdb2Ey
cFpuxO12hePDYk++J3QmyItXOtVA3kbRijxdQinHPZvRnnrbX0EURGLCozWX
hljTNjJrmFUU4sMuZjhbBVkOFsg6AiPJ4hdM1KuYsK6WhKx3tz79N7qUPgWL
PvgRRfh5hitmLF7K9mfWUGAGOcRVUaCQl+kBkeDoRaL887FXDWZZE38yjTo9
gAl6HvoO6ueqFJKY/V0/uM6W8JzAkHZal3x5e7JWHir9RyzNbwf3Fda4IIOE
mvhnDimIDf6TAjOzRxtF0E+/6OjVcLXoVE++ByPypsvv/5ocvo9EQ944aPNu
g9eDXgpgZEPbaqkfxPLovyACYnwiH+y1jJSdna4gincJ58i4olNbST9gG0xx
jlEl/O1Gp+cDK8irC2DYxazjjjz+qzTIQtwNY8lA8GTdDhVP8jgXFnM/kkJM
ZcrpzlPdEuxZuQBqs0i8m7Ocot6Udf3SHkU1ebcb9hpod9AnMjtmHGMC+XDA
/ht9hA7SZo9zaOS5LEflHhTgT9cHqZId3csqVPC8msIWTM2CtIKkeoZyMF4O
KEGIhLuaOcim7xyzVGlmyi8oz5iuvLtAhrwRgY1X5mrK4ZNJ68QTx5ebulMZ
9Czk1dGn90Mn+VIF3HqyZUoMSy2KewF3uOig7lYzYeoRKPM2c9b7eg6b1QUt
tC+UKdwymzYlVO05n6Ao9+ynhxG8sGnu7UjDkKIPbSFZC/UtPcIzWLVKNv5J
+kHp0xcYH304EW1T9dwZBDVKa3w2uUWbsTslzIAtnM4mgc0ARmYkSe7/6rLO
xQejjifMFzPVhVwu1U+ximk+EAbsN3Xfe0T+DwEV0jpx0sXjZ09CfVQ1Gsq7
MmG9kQIvTZmjxihRxSvpvAYhZ5FPunEVc/lzU6gL7vGHAFH8TbcQaQ861Ug9
+HamRySL7dsZ6NNGFN0jHU+NtW/kWDXjPvmb7CzSXVAFIWlcgnUGPXVSS90p
5bDJVmqI2SJMdvrQVQFCMGakWzRO1Gt40dKmrBJ+3lNESf7ashmKrv4ldkuy
YEtcoErEvRevHMohKvZ0xPAqrvgeXO4CJasi0FDAu7o06AQNjfJ3iSQAtdXL
csg8R15xXTTrhnpfjo9Qc0Bbcx1e7zH47ZHJfcFtILsKJQHK3zTs8fMJM2Lo
bTkALhzOdw5viJNR2tmrSN1oUT49zfiHB7KWltZ+6i2vObasC9a6M7mTMUQQ
Pm9GW+KYwDK2vdgdKxJIu41sEdZ8MZqV479TX8SSvyc0GwygX2nKNnG4mzPM
wEhrxGHrt6zTCwF2iIrfEBd7Zg6eqPuJjVZNEKBw0dWftffvgwr5a6mQl9yJ
QOJ4qOd4Hgf0OLFSPcj8/o+YwzIIxZ7Wa4Uy7xK/JXtJbTVSDmdEMvEzK8Cf
aQQ2ORhhgwX5rl0AkalHSd9MuHns3UcE/drd2HZYH3L+aG4Jtbo8cYW8xCxT
YDiUfpG5AlP1IdHEi4N22oW6HcxUVjbw9il9cBV9MWVOjnVwr5id9CNXTNBi
uOKtdaT266ekC9Pa6DeNvZPz7sZKHJiS0fnIlDRK2sjgsA8p01cRD+Z4GITn
Ao03mLo9HxsjrGqoWNaOHPMqJp/yozuEWqHHO6R2aA7bobFn9jFEbf/XgiUI
x8dZ4Mdakn3LgOPdMWoOOH2/8dkAlsy7a5rJYOKgrw7rskDVIOAJJGRsiUnx
7aBlTg4MK3SBqTUc4GhEsRMYp9D1cSzRIceXC+/88+wzzFqk+nTtnwtZ7f54
tLocifZXnYQbFLTnLEwGuEGdM54duzApVTY7Q5zVFDlcg/T8t9xuFmjOvSXO
2zLs1YEKS1AI9fwiDTPiCeydzomFWagBjWvc3j/AHZvu8WIg5CGkKIEfIofP
7Ay8Kblc04PpR1UxlXAT4+a5O/DFXUpsxNY7Dcmgtu0P+gfGR4NlgJUekzn9
AUmk+f/cG+h7nzheNDoumG4EBESJN5acGMZCIEccVWpAdzZjIbNyJxhb3kfO
Yp2zT/a7Fs/tYYa7dmpedsSZVkpMTD/txwtlSt1mS91UczZohgXI1Hi/s5NF
wR0+sbguNPJUaLsapz/6TlCqhx2+nsLr5LXiteCX2ILHQJFQBTK8oZOzPTDj
kC/iTSDLq2L7kdWgUWjK77M3ZNnd2RwK2Hq5JEVAzKNG4C52ynqGpdouiYOg
H7msvO09npmQQZjXvdk36Q4WnNJw3188XeSOPh1MnVjNNVX/N33xn+W9nkVB
J6EcQYf5eJkmW7UPCnOXDhe6MSSz5F52SWVhWtrC0DDJmm74spnBW6k3CQwS
t7e2eCuMRxvddlH0armuyEAYKMj2o7oFasgtLZjrVY1QfrNbaDoSKeCL35Xs
rHGLpIf9X6JreSclb4heU+HbCQay1Z3+BTYtZNnBbEWEYpLc7PVDGPdUu5HZ
p/mn+YPG8bww9WFFFv3J4vc/DWOTtBshbyj5FJR9f0ZcO31+NApNb8ON0NPm
n4woe1y4TVZzN8wHqeYiFKi4HnNKNq9XTLmKC6x/vuxAscRfaRRyE1vaBlDk
SjtpLZWNDxQ/pqSR3dnxI4scYeDoGZNwHj3HrMKrJXtepPtN5u7T6avOg9yp
PULJpYOFA8bmShUrvfsTnv1tH3wdE/i5/TrWEU0BgHF3kvE1K9sTcuTY8JfY
+SVNp2b97P6shnTsH88myiDsO7mM9Um6kb2Xpfb7Y+U3/1W6MYNl52VVZ+Nq
YW2xZjCGUMA/laVNAJzxzGgN6fPOdThpY5k144heBNUduTfndJk+nIhE9poG
wW3T+Zt90DdBN+pCzlfcoZwd73J0nrtlce7FlLLNMKiejOV2t178xC7fjQ6H
XBYnFKFQ6AC76QHPXUOMUi53HhnUzCOdGmC+qBKyo5038R9Bpm61ui0l1v7Y
w2xkLPT9126MjpZe2p0l7kaa9mMj/jec2MPX+y6ucpm3iRlzN78K8QXYb5K1
LFMFQLHjRhLCFNcUbKpPFo0PsaAcB/kpd2rH7WBIDu2/AFT77rYABVtDTfmm
Uu2mbtrRwY0eb2OT5L2M58grFFBU7rFNzF1+ZrcRoDCML+vPjCg7dkSrlh7S
WKRjtKH6t2u7mHxTuiLjqjzUfHxqIxXjYMTSUkCAVZgYCDG2ukNo9/HTEda6
tnVCyHp7S264wqUO0zHsgp/vbXSMfFKoCNM0cY3/SVGpFxHbtzosY0nUbiev
wZ3ZKWGM94S6GcXsIzIKfyOENertIWhAT7nMBgRJd5Pb6iPohxxaqxtYyDVR
44Ag9fGURFlwervS2ordXVdtstDH9H7YxeRIO7KYvI0Qn5HBOGzxFTGNaf20
hbIc096gH7QUrg4NNhmkOrCxbz5ppw/oG3paDog9zPInTWrHEvVSxFg0YMU2
TUJjKtPC/yI3vkFm+GJZiX3M4VkqXnJDOglSBAl24LITz1GFmGMf2ZYYJc5i
Xvikj5qtkh6HdaJ5NBC7k1XHIllNbm9hEKCrz4Z2J94eUlzqFnOM/iieIMBl
lH/RNFe1VuAdk8BBH9OR5PiZQ21ik5OPuu20Zk8L0MogklIcO7mhTvRHbIRK
2uGx+yz9drq8VzSa+6ktu5vZnOqqhRsI0m8+aNDcqXuD8K5Qq8bYd0NYbVMX
+oA7OOg6rw8qsvgdzBhMV2xyDmDplmZS4G9+wGQdttD4QTXIM5TU3ismEx2Q
zo2l9BfzwtbLv+rE/+SA5iiSviHY1sP4SadeMyEeaXbDJuoZTjyLo4vlMM5s
+dmY3LnEJN2wD9l7CNTp/NWMsU416E9gYhpv44SNyvLd2YIs9RwQs0HdV64M
oGL9tbolfWHARTVLIQR62Jd3TQ7vQk63aTcNFMz37ifXls+hpXI4pBmQ35OY
B1benM163l3gaogf9gmsUH/qdb+VsXqVOS05NUc0tTp03548kVF0K6it35+v
cuzu+l/jDqaqnuK2bVjoAMx5RZbn7WYVIEw6iGeMwdydF+xqNz3i7Q2F7wWd
owbrc8uatlCGMErfKhGEOenLg6u9c5i2Ez68A8lMdigS8uhafSoRGbU9Rv5n
wupIAar5ktTrIr/UT4mEBs50ov+8uWEdbnfNt3cTQwfmrENobD2L148TwqI0
qIavg30TQmo+jtqIRloJlqb+tKvmg9YWNIK8YbOnGzTqmPtC5xahc+8tQ/P4
lK24Aim10uiiCQ+eg8c4mJPLIKvuHAoVwD8SZns+GWeBTKftoSE3L5RBe0JC
2e4fpV66jZSkyM20aW4LQ1PXjjCjBxND6oyqchY6gARAurd5f1EdfWlMAc/C
85oZxvKvh++BFzEsrLcIBZEQGgqLroBQgfLPl+AbGyISi6RAhS48ybR2qyjf
j/aCprlBx+9tAFDoTN4kzC1fqeSKI+uvdXhx+h8OuQWnMPSyMClbQzHh0XN0
9AdD9TOeT0SUFlnmRUs05NfYAKCeQN+iL15YIPafhAgFxmGqsfvsu5SpL4B0
clK7f2kl0F8FqqTxNLrz+1JkjrNviFyJZH8thy2/ajiCmBPHAvIoEuXaT/EO
lG+UXh7eXmWfN0vBDTteHuAJ3lmnDecblE9cv6lpXuCupYzv0wD/Gw9NLY0V
erFKd303FbNeC79hg81JePHwtImsEMnRK5DjgkxeMSpy6eF/HYaj/Ch1BP41
wjNjwh6gtYX9LuEvXec3hImp55AZudDObAvPeyZozHVcF9X41fz/Zp+hHWCu
u8dSyguPNmb9L40YvfhTkxOC28qziLT67FRVhcmEbQJbJIO1WlW/KRXf6d21
mt11ZQdLOY3ct03ptR3vxhnMYcR0zIlmVp5aXSAcndvpihNInZJFPvXERLvH
IKiHRYmsZpHFK7lsPtwOcf6Bc17XMz9XEJE1SG1GsiW8JlbcJv+0Wyp2JND5
1VBMlODgOb/utNrcMeot1+TVfBrkzFyX1Vd+sjDsuZhtvrT8l3zShJX64Oej
1WqNQjNdxFZ690i/OSNdnQVTALLHRk41X/x3ghBPHCs5JvjrsVzdXuCHMTdm
8+LeQbccaIUTZeXm5Eq7Sy5XpKRV07x/N1dWVZnhIbzAD1qRCjZ7ZWMhSJ/m
kSKrGRTwLPOxuxCmI8qPZLrtkCpKr/fB4cn3VqQERDYQh2vBUUoLDtglRaVS
pwGq5OEYRTiq1YJxMme3kdfJwf4P9UkymA7qRuu/vRlws4xWg1eOgR+s7Jql
aqOGxouyjGb2ZTNjZQz2L7wdSB6UjcvoIJZLgyVhv2hdFSE11uOXHNiIJmIJ
QW4tPnPsJ4pcYy4YcaY9qQQYzt2lb4bL538xYfeoOklrXuv9AS9uN09wyhN7
Gg+UJRVITQP2TFoQHhMYc813oVNFf0yPLdmjurD+kagF79kMtdhULAQ5htG5
QicZEbQczQaZzMkwyU3ngQ0Fa7AppQmZ5tegs0yEVqv/h9qwuIeSgxJpJ+sI
TLLNfx5oa+GDrZh3WUz9xSM+pV/6og6jyLRJWTx9KLtucB2TbWOqFVrH7lq2
4/HU708sw/dc+QQezFuMGrrs/BsJxkU5lpQnYtnPm6ee8W3lEKlqoQQUGNSY
6Q/bHioyvHUnSQbqK3/ZhpQmHZAihq1qnm09DQERrVsxOFynN2ZPvdDKfbsX
TKn0uWbB+S2ZjR+CE+DUcw9wlz584akTsCrFRr2AgOpK4yEPBgi39JfM92L/
6+o5Z5fnVabbq+OkhK3NTY7ovsobtrhDg9BeArUhRWhxANQku/qLhnveH28T
UUXnhHLznLAwdHLjEoJMatWlc6BLiWrtfkstynkJ3qR4V5EHy28Lp8eDgUqD
qAV0/2lw4Q2aziUjWLSeRl+IwmeCHinH56OGHLc8/aNQ4K3qe3BXW8JDtCQD
YYhovwiGBVh8Y8ZSiM63KD7DmdZ/+L437rw/vziZRaEhcP2WoeuaDSM0zz70
PdeTGH92lRA2FWzYGSlRObTZhIzo71fpyngiY45/9XabkRGIrKFUtyk6pt7q
ni1QHj6CHt/eR+PyXh/LzE0uysq78G07YpqSpl37x/XvOMkP2vil7lxioYri
hqo8sW7xQpCGX0pXNr5vdcat2q9BUo0phEbpnzbmr97cwueQfbqoVOHQRJ9b
gt+tA3mV44OeEpxHeNZOA0iNqrtMDIicrjpEbDyAwvXbrozYMA1+Y7Nubx90
hXc3nwsqx5Hvelm1wfIpQ2zt6rJ6NWoqIn6yN+qKwkB8VkFFjTehOXZBBTuw
mHzYEYdmrv4E9lLmCxvIQUHfJ54LYeWRWVw/jG+vkoMPuSseatoadGCEZK87
ejVt6cT9vQFKh6YfmmFa1DGQuQ8fZd+Cf3xIxALtrosyZ+57MxgZZ96BUD4K
iTkjDJ0H3xhIvS4sAXE3Z9Xq5uHylrVPTH1bg2W8XzKbZaG3/izMVLIvmIiQ
ppong1LRz/q+wZK5EX615+aS6B6FmKaoYg7DPTnekjX2XqO1C03hb5KpikFE
LbIgItRYSdngaL2x9l0fXFj4XC6xxlyojM0qZhHgd8jG2OfN6vpNFdpEoRLT
wrJhjfvFmCYenVSw9adeH9KZnjgdO2YPew+5j5ahgx+mEcSMljgYzO7mH5Uw
qDaqFp0gHV6xrirOcMyQkUFF28KRm/bhDwyF4vA/QqRqDIYPu7qi5EN2dPHK
WGuDAlsuoZo2maMjQlERtIjy5O8rI75LmOWuJz2PDyZm+M9oC8Ojmtgew987
laIV1B0zE1+DaSnr81ThX6ktEBZ3eZjP8xnw9gLs5nLca1JM/0AikAQZb6wd
nzioi0ujuT7bS93oedSez2NocBYsQ+xEntMdE9cCNn/gywilO/0E4Fk10Bbz
4qqFIkOTS3RL5K0Ela5NT4uON0WWEeqzRU4e3WBb9RtrGYgIqvmrksuIiPLZ
BsdnUPn/vLJo7MSGD0ehwFfK5oSIUENq0wSwg4MvAwMcSTdDuVVcVUVO75lO
y9W5mwMbVFCw9E9NdQP4zDxkbv5d4XuBvEMTGD2/+mbJy9YyDNGSKNjoQ+0G
amMkUlnJrmi9R1ZVchh3T663AtdyAc2rrkAgHO1dlVU5SHu/+/TR5CS7C1tr
AC2uTJ00UluIXmab/zmwMcp1BrkYo512ZmP/80cjsKFifMDQpOiF5NzJ/9Y8
4aIng+Frd0538hocELasyvnXlmrlKl3+wkLXxwxV0vCOIVQdVohzUIrH9hZJ
NEHT4oQB44K3GMWag8xKWGcLSK+6BE2EjA8/4gMQg4hVCH7AQsu2P7htxduv
YXt8CaZ6iB5nC+W4F3ereuRv3tHvILYMiKzNyombMnfo2FNDRa77RgT5kDpf
ZuqcdYa2Gk8pcuKX6VdI17sjhj/hvR6UgTJFn+2S5HcHqniCq74woGTlKhnD
y4bP56aeyHiNlR1903HfLsKdB3VwoIOXwfPk0YgxlfZvRoc+oy7tIhnnwhGN
TDDvZhw2CRE9JrVV/sR7OVELNTApJIg39d3sGXXGgDQUp4aq/PQNA4rnmJDl
rlamOQZLEV9gfoT30olF/i0KIfS7MRpmoEwTMJpQxX6QpYitnx7QBscQ54+W
97LvpcJd3vXBqbpUwAPzv6JdVJSnbAORJKncD8RcYIrKJaqUy2URr3IdCwAO
xQCEKlSlftZo82snsIhsVbBmIt+UEZnZf2FtCNdPx0w5wDHaV6vJEQFCBgzo
Ok0zhlCf1TU9D/J1LqsHYx28OZ5sV9qmaec2n7+uG9ueIc7yH9ZUnIlJB72h
38g40uregnVFazUKOMI9xu3jinS/unv57sKIaMXA4KzpG6Q0D3VGGxSvmRUC
SslVL8g1efoBk7DD61kzUrck6xuKKhLz+cOPMT46aYiQi8rIaKVzzihKTcYs
Rg6Dg0CCkH3cM5Op8WwbHtB3FHA1Lxs0dudUi4e8+AIQ48kQh1Q77sOqmTqk
K45AtkyEIgcIByErb0Bv6slG1eoA5XzwuHi8U/QDdZjn48vECr/rSeCqnN4H
kaaeytNUBNRdQlwDAupeqRC6zb4ZxPng8v1wtdhzMk3rAZlTJXO77K7yCoLO
Ju5JTg1/PBRq01D6kZO9bH6dUHj+ggYNYxBA+8K4qx6SkLAORePucVlw5ojD
ahj7jlUdKyZvFhkl5ULYpYzNj2784QCWlAbNG2Y5AR+bSOFW/+OHwY//XVzo
VcfDjVZBg7JA9RunIbVeU2vQNErmIwhO0djxjgNyLfEzu7c95DTbr3zdNDAl
kHN+VJ9BMMHlvW81w9iPFbtlLYHt3xnoLFzOd5fAaSwri2x402ohhaJnTZhr
7ATDD62bRVAHYPbng6dxF0Cxm0rXIwJOj5bWsvv2SOCp8soCS3KKRDiNXEur
aHBgGQucexoxWIMLpP84e1jD3rb4wc3peHfgf4HNx4yXn7D/pfg4DyYTgXyr
0t0YC85C3JegmyKsTSO1xbfQ3IJ+pVrTTzjJmAI9PS98uvkzuRfLjTULn/Q+
Jez6SOLd6a7S1NV6iQgwliCtVkCNoA4G89EnXse8bneMS7ZPuobI0aSslKUQ
VfmkpXi8SzhgYo8rYdDowZWxZoE3jDo4L3HIIkFbQz1DXdXHhO+TEo6Js5Dw
TcWvt8wFZpfcFLfZKVVbiqFhMCwa1NKEhVvcf6Hog2iYLu3wCJAP+S2ig87W
RYjaY50prvzYHuqIOA0dEQJy3gLFawWCnJ7mjBmh+a71Ak6PuZmRu9EdXUVM
8y7pGabALWdaaVkL9Ge1nYVYGOlGI+V3oP8uVAnBwEqEp6caHjd7bDXO6dbh
vHiPzStL/r+WKW4OUjXMIzLa9fPU+FAkENdCxPZKQLdlhrRnTv7CXjEPp/uz
7vjmWAE9iY5C9U09/s+J9qK/YadFoGAvKi7OCcFejqb+bFghagr8tkNgGHVP
gdAaCYId9ge60SDFFDpDNIyvwRa+1XugWT9TF5Y2sEcSXe7y7HB8ntPw8M9g
SHavSJqqLja/RNnbdoCh8lK1ldJl1g3jNpNu1bH61er+XbNHX8kP12Kj27pe
q/ASFOdv9dY7LjTAGwAnuOODxN+yit6ATZQfV2qJiBIUWmqm7EmFs1og+atY
PksYDN5mxwds/h5e2vCfPgKSYz7pUaVJ7G/zq2bVWM6UZfYy+CTI9H4fTzWp
AMwQpEnX9uSxzu9MqRDbqjIT2cpcfZBo3VUhhzIu3+OCwsTMqqvssc9uFViG
WkZcqH8xaagfE0UhrFFjloZ8xLxpd3hWbXk3Lo4z+UeV3OdaTN3q3Dsq090n
OEVZ8THoK6wiHdTTlNpSP6YbrA7kWf25DF2tPxRZXiDTU+k9DZhix+yWP4Wg
xi4/SoN0xe6rqWMLXMViRdx/7R45DIXWevzoZfbv731OJKGfpzw+4DVJrVnN
xQQWNKggwYaFtc50itUL62skDTrOoPdYdC19yt8ulqfn/es1rJUZzAU8NCyW
0YRPl58JE8k8S+NfbZnvNuK/gVPJw4RNVqtGHWf0Wa8wi17J+v5kH+UhxadZ
IURRzEXKaiKWGAJFeFCZSrKTTWm+ppx4hncnUIECYKRZDC3+kRr0A7W/e3lM
UlScD3E/f5kWCmIOg1wWoN+CWdFo69VbCKqEKykTG6Kk7v7k6d6bK3SaJKZX
gW2icp5LTkQ7PUw8NH0ubH7zh3CfZklwA6h1DCZzvBKVCzbNg+yYrVA+ITsB
QEAsWCx9V+H7XfFrwR2lY0grXwkzt48Cq+ghPuntZ+ErOkrR1RdiCCz+REQx
I4fQ4g8CQdEL71gmIC+9OMrUuEDw6Gq0wM8wI1E27R7AG+Wb2IJfnI3JWqT1
5X33/645+h0RbeHg6x4MAwLXbey+nycVCrQbTnpZPbf9IcQ5KDkgDYUb72Zm
OPK1zsZsw0lhZKR4ZyO6lM19KAhMMZN4hvR4nT2W1qVrfuNQkvTEIP2UhLFh
4qlmb2mRlq7iM6QHutsuqFL/YY0hHAny1i5uwuZhkXcIELpUbijvAVkm/MhB
rVJ5rJVObnzCPRH0oMfq++r8wl1GNuqt/aLuNNYk/88i7EzEMrT3bryf9sI6
aDL4jtIRePOOy658BlNIvyUt6udyN6IcDKTPkzgnlCOLXhOk+poajB14vpQ3
QY2IZakXc+5mAB1SeMrLRROdCh2ths6pStWNwrOfCObz/R34T5DYnnaakhA7
PYR+D+CngNAIUPifeAMHJAmpnoFHZhR6D1oalo+4oQIOG4UCbbmY3b5WdjFE
zh39G5s6w5kJdx6yTOv0VFI0N+4bsbX1pWSTn7eOltIdkZVhiVPLumyohe21
cgBEiygIqzlFxQTehaIGfxteYmEvKco+MuWhnd6Cn1qLEEfCFc1fFyc6f8uT
RdRsShIeRq3V/IBf3zAbHsoqVp/gppjjZ06VAxMyWOwvFnl74er6ggQM4hPW
A5/p910Qb/231JmtIYNkdIIIbvY7FWS/lqI95wLftg5iOTU0rD7XcIkSxaq9
h8xkqe+NerQ16dlb36higRnU73UBS89/pMfid2q5vFDAakqEM176X2rTXehH
B7E+O/lNbUtMg4ZsL62iS5B9N6ojJzv/uNs9ei46nceFpM87wtmXe7Uk7WVG
ev0EPEp98meWVRyfghlUBb8XwY9knhU1y55Nkvlun5QlABVPEGC6NrJLVORX
bEcTeq0F5HJqm44DqJmJBmQmy8bPARdFguASacXD9onOdS/SfO5cIWzDcOPb
ubE+zSKUT0HwI4tvSS+4rLIzpPzQC5wQXqb8cErCSBVo9COlUF1pmnyiso1/
tXDy0iuaD6wG6h2MmsSnw/6O4SKojgSyockTJGe45gIjLSDt7KNq6h2w9rEO
xmiyHKxHQpqoEzFhLEEBtIffrJu8DCqDZjdMsBH6nqEFV/LlFpyGip06kt4x
YwJewFJKDmSTcsFeYucmjsJrKy/5V5ogjyoBGcNdst1mUCcVmHpeqKh8vHwR
+vaMtO0Z5+S6I0Al9uWh10lZ5gse566gpoWPywK/pLguoCyAXhQ/4pHffQ7P
Ybf4mT0+VqZ6gOg1feVi0sTDGuhDbMfiABzoq+anwsFIkOXLHkLA1qd937qR
llc/7VSvFRxkdlIA5NYJEEHRWGZ5TppQjmxSNHKSjSI7z//vNtMhB+ehnaYG
vWMKg9D67WbGXCaVDs328lZo/XXDi5RiypoQmA/lMtim/I2FbuSYPPev9/si
Ia/HeaHHKAH0e4HrNijWwXfxhhT9FxBH0f8l0vNdQHGSBpDxo6KVCVaQnIAI
m6jma2faLrfZhyn2Ba8T5H2BzuMUsTK1PIOTtuAUb21Tr7FDhoRixAMCdsgn
q+lv07T8rl+tkA5XFWed74ieQ4nTy7Aypv4GfmY41aj9LRHQ5Fp9o9a7+91/
csvfrz+mRiiyhw2/0CZsiK4MzILzJy8gKNtcAdq5INL27IXS9UOoGzERCHYb
p3vu4JNG2qVrtYflB5+Ct3i2uh+v9nQZMIJQWg9bdh4vg/nPHVqEvfR6kGd/
Q1zdvMasvJ50lck/bkUNE+k/JGDMtA+q16QkECh0xDrMwqGCUdYHytrc/P2i
jR57REpYfQIgdI00abCeQk8o3K/JFAe8ePvR+bmUAztY5APEnemSGji4v7Zv
L5aRVCfwd5HTs/4beW/+Br9yr9X9SS/zflo+gcP7WAUwIRjLUvkB0ePRHmoL
l2LDT5hQgRxLo1p+umqCNVyOO2vA5u1oNs58gJZREkUbG8vCkol1tXfCpIqs
kUNagE/D3J/nd3ywFOr90Ll46nLRtC3Zuvym+Mly3t3QgQBhDGe5sLsRhmyE
mQ7uVkfUukjS2nNgDA1OBIK5iw53dcjyQs4IN/UM6yQS7rzgnvmQ6Mkc40KU
P6OQ2KsO7fX5VQVK9OpVXT2VA4WhRObwLaDbsdNbZfjBYyQhw0DYaD0iaS4d
cOZyCRzTOLd1Zclwuotj7WzBJ/j/ddrRfLa26M8AidAa3h4nd2HnVeENHvzz
CYcUpvPxyRNqGiVmW9WA7FtzoxlPaH+wHPpTXvfa2+nGxI6Yh4Ir/RC0U+za
8HJY11gZkGpP+nwJ7IhvgnLKcFkE76R07KBqTlvxA3PgTIigKYBOiovhLLR6
ues1F12StHwqe0Tig2cZcxnpzy/SHCFN8TRihT2L91XKPYxOQbEN+AQKdvCF
9cHqno7tyizvNLoQyUoWVP/vFDjroGB8y/5xdTsaSolOnoarBN8Xe6z3uEII
BzQYjxHvUO8BeuHm+GbS5vvq4QwBLyT//lC/Cxyctpk5PlO8Id7pp3GolCw4
M2GMzx/Ohf1eT3/5+bUv6ZvI6ocoWfJWILebPB3pHB8YbSK0XujSRDzpTTlg
NC6zcdHXyc69s4u4n3IuwlllF9VoBQxQpUdyY/n3AYflpjB7CKrVxbpFT30F
8zAp9a22xtUArAEFjAyfJnRRI6EHb6uh2z58ZfgHf14Gz3wf3G8+zGHH3rTv
/KCHAGxDTkoKOMIIf3jZM990NCBTqFSetF4Xsg9+yKHEgrdXofuRTg5JI2mW
fJFbgf3Z6uZROulZ+YDgHJeQYaEZ4GAeFzTwLKhfazIaDVNAsF3DjumGNmVA
aI8KWhpfMx4U9jwtBas3UTlVY4jMYd4L3qiud5TBZTMP3WlcT1zjr7r1Wq8R
C11TX42jBiUffMqydafV3AAdKDtYVu0KrlDF8ykJzEc3kl+hfzXxzN3EhGMg
g3t2LEKD2EaS6QvViayqCasBz71R2LxpMLQ+SChodObV1MitPuXIaj1EbMgA
x5GfA2I9m742XqUAcf/LZBIHevgcFo/Ll33J0DKRvgzwoCrUFIoTaLTFP0ND
smErqcTo7Lrsa356Tu3/lhC5fNZ0/R6BNaLAG2gx5b9ZUoslNp3CuFhND+uJ
FqRSa6aDwz0eoFrdYbCsp9g7joonFQSOmDmbV7T8F5S61/+lMaBh+1aN9WG+
NT3udIiJRKTavXG0Iaw2wlxMJHeCIv+K0zk9UpaA30ibf3QKdwxwQbc4ToZe
CDlGru+9nooPqrx+7UvTfkkSMHhu1j4KrKavukTDtHtsxRBHOxcXsoPVHDAm
uINp6wlq5xEVDpvtEX5FI27UTmUTb54sLqtXvqaA4ie2C39eq4Y8vMABV8kb
8YNrRl4eHRjjrgjCyqlpxCoUDmIT611wwb4pvuqmbO1539zXABM2l30mK76k
TsjwWOa135BsIzfwiaeH55yCw63VhXXhCP5NfjaEiBDizHIfFwRnBFkH/YA6
ppAFzyCa7OHeJN0kPMUtuf9UTaapb7rj+MXsQGvljM80Ge6s7UGDkB36femk
nLJz1YwYoCLtLNTmh1pSfkpccHoGr88jzGYYYFHTtH3S9Z446LfRPgbIOtcO
fUzkyBrXsUIRt7z3jCJ98lJecMwoqTe5ULmNqwZE3uT7+CfSYGrRIiEYtVx4
7JLxnUuRXvHTQGeWIj5QP1t7cyf0oaEYS74I5NJg3G69FUVxkpAh224h5IyH
9RAu3kaZRAvhoADeCtWVb9g8eWIALZbNA28gYX8IBTK1mdmb66RpvfV6hx9h
kx+rSjB3w7TM2oGQ7Gctv8uZ9jm8LepkOmeesBDhojHw4klo3LOgTEDKmF7C
cDXAymzHOHhaagx+ApYQ2Mrj/Ll7RmCq2PA8OcrXWWEOaCk27GrpvJxA+nqf
PUHD+05hACLiSpk+u7jCAEvHYth72yyUkKAqiC8IXh9Xj1fKST2jJVYH8W+o
qaXVRP2zs89fRDO+dutS9n4nNw8AdzTEF5APRRO33P4kCidfjeTXysTVWiyE
XDpFsotJ2fGf8jHSmjU5aBG3OSoj3vrvB6nXMQ9e7DivIF0+eT2nXjZVW0LU
sNnU2T3ss4YTg+HYXE6P/hpmdcsJb/MpKgtD3/To3GJ58HPIBBoMuJgPtE/a
W+CunyYWBoezr/4Mu+YZeSHMflBQg9scolTOXS+Wb5L054MDseEkKjt74697
Q6IAS3tvccmkwlQxiCgmmAhpYzcyfxQ75h290PH28jUlFXTUcIQW7v0PM6+J
+oyZjRTWc8DE7lo80eykEj7BjYXPNo8JDJJWQVzCmdURXX9xj1DQsQgaYFeP
oGoPCAKvxNp3FOzsaHTSEqkvhgGVFXXzvbYnvlEe4pgaSgQN+hUQQEfLScpx
nxXNo7EjhBbKSHBh2i/2G1pE8WDa/O/Mf7xyd3DtAIEM+EQwwBbbEFYc/Z5F
GoEhhg3y9JG0tiflbw5zMRnfwPJ9g8vyylDnkWdGawEW4vAl8VXsLx7eHsQM
a/59mzdBZUNAJj92zsrUp9vRJ/6SbNkvILkHcPtM4bJGjBOeWl7SrsV7wGME
6xZ8stQArkG3AznccPts6vQqpNoBkG9Scxw+ciwBFekYm7xFCI3+YgiOAdc+
J8Ht1Q5YSJ4b3S+eMAutZAvUJdM27eh1dw/8Sh9vtn/ckYcLntI8pTr39NDq
psL15mxE9FYF2QHK6+553L4fK0m2sZgDuxhr9ZL6GpiVHYGqPWfymXKFvUH1
soyFcaV/7PuRhvJChLXjFeaVlUgeqEJlZ7+IuOg5T6gycSky78OIuQJK7jev
m8jU2N4U6W0L8PpYVUUF8NiJZ85nN6M1j63D02knLZOJlRJXr/eI1ZpIXHE/
jNXf+gEmpwsMmBGDS9ejnFfbNO7thfCX5Tju254YYiXudRsU4W/00uumpiD4
iX4sksVnjAh1HG7GJoacVuVJfeG7C+z9WEvH/k9ITfuEoZ1Jgep2ZPA8uqAF
EdTWe4uCnpDDHVP17ru1mXM9CB3Hk5ynyh4Ljspxja5zIgztKqAoJ0xFWaFN
BsjwDSlBv3uDxCaLI7kK2qnIudOOYAGM+Bgl5mW26JKymmAut0e8DDDpzuCw
U3imGwFvswVhBE8Ku8XI7doNBdX8hRpKawNkGM4/FR4nxBqdkcepi8WRPpPa
CuSE+IhTpKecmoFbE7n3662eZ6dPG5qqpfKyALYoMOSZEmMZi7Kn98v5ouyx
t3qI29WApkiIPruhdvYeqXQr+krHbr12bwvwDmPnd6/5O6jKYloYrFjv4vSi
JM169SdCwJIAeaj4Qg1vA0wxoeJetyojI9lrPVob95qkPMfSWojVI5Syc3I8
e7aSpgKuoG+AvLeopnrWCkIQi3ieh3j1hPv6HSuMsSSJOyu8zFmCj9G7RL/R
w1v9I8Jh/dc99+/KcnU+40NA8oJ58xarQPT/ywyp0TorImfHkeHnuqI4lSRH
kmPT76zzaPvNLGyIociusPuu9ZWjS6Pm2Yjy+Ohp6gVKyDoErzTVM/763RS3
bp6Ee+RSS3Ua0ZckGnyRnM3/jgrM0Xc7zGZhMbWYmtB+ORrHIEkQLdbclFfg
+cwA6jN0tRkmR1Ar36BOmjrru45u2XUY+gH7lwGfziRgj/YaPZ3dH/4aQzLG
M5NY9d/w1BMC52DnK8sB39VJppl/+QrLD0fP3uQL35d02lWk5mA9tgPjOPhj
vJ3A7uEq+0vP6CxpW7WlEUoCK7yTPcnBW9Le41CGEcxF8Y2gez+HyKJtaess
imaitITyjJgSjPyOPIoVaLgdr95L+nTDhu0I9JFzWOvTwINjdqopFX67mAyL
q4yT0NvY6Bppi6zTo2Ws1S3gdFKt8/NBC4l+0zQj2O9rZkh8ZhbWc2vBYRd0
5yoPDZY5F4D5eiLEFYgOylJPvi0b3DiTVe/BUAHcWOQY6MVjUQPTEeAbhaYk
lYmCi3U/2EjzlRInMjN3w3DHuZjADabfZ4ox6bmJTe3zKXQyy6I2RCOqGieF
3DJXLzqCcqpOM8RtJRygtl3fR+7Ia4q2sNnVjDLbbN26q4dfkxb7i+VPu6CR
8u7/Mg86jzflq3ZQonrvZMTY90k+y+gtGJRDDuDc/zf23uOHYr3gbix3xyxJ
yMxcLraSRL4XiKhApGBe6/g2NBp3XdUPT1G7xd0nY+U2ytB/78w4Ul4XUnXw
80jn5zieTXKTV4YiwLwCLFZNm8lgT3X2a8r46lFDK4w3JxlboeR4AM2Acfyh
rkVOrl79ZxzC3wCSfLlU01FWTBLfoK4RmZFDLFGy16WHIVG2hJk9vXWMIpaC
ofeRuQdqQ9uPfL7SofMwhyBcTlOJ0Ajk05Yu16taYHLUj2Aid8V/VHB+N24S
15mH0EBGwt0moSyg5j4lu1HECuoMvQTweLnxQwwjBWaD4hKNNvlXY3i7Je0j
XvktKLOrxozoNVSVfiweyV+QHc2ylcVcbM1Mxi7bJ07k1mPG/Z1epp36g70e
+XeAtgq5xm61TGQJZeokwVTI2c8K7X1+we3QeLV/iaC43LatC1Da/2s9NHiV
UVwTbwrLXJ2gBAKg0IjYNuWUK3CMxD+LriQGSIuypfOvTlpxKLpGbizBwFNW
WJ9nomUKEQsf1+IbbrII2UiMNqaRxiTHJ9OC8lEmcNS9EpFMbCDWWTH8jhw3
ujqHSAh9BmdfsT3BbBTYBDdElB1zEDFOgo5yA2RVaDUh8QIj4/VtHKPiuosD
wVgd5rAIylxehy2ymGq0AuNE0jAQQmadthWE6fZHBmLu4V7WyOsiZXlH+jag
rrVuaxgrHYoXdP8YNlyacIIEgObKaI0CvU0w5RbTTNvU3yO4I308Ge1YANnM
bpxIggbPa3SmAjnSoGlBefwOWLcrzF7OwStO3xiuvW+xLIYrLGNqbsUrijGg
UDhhW68PUZK+55gRDXhsUUOIJtG0EUYROUikd1GNdx+2KUkx7ii5iIJM0ETc
bPEuxh8JM4wgXsuQWx/jG9q4M4w2ai9T8a/mQziAAO+xcKTzmRCGDNUs6+mU
DHr6M0vUxrADA166Gc/+f/aIXY+lnlHTsANCj9jy/fqivaTI66d8j8eUvyjl
7TdnIK37RynP4nJ43p5FRqSizfvi/x0R02yVNGHVJiUqhpiu33rJvkccP7S8
GAnGQXgWpQEW1tcuh/ZiyR7irIddnd2FPcufY6rid4ECwJl2g/D+eYl+mXoA
1gwUBZPdI6On0yob1wPMdCKWWF8/iY8QunGlIs8WhAZ9d7ZIPZFTk00oTG/m
EEAiJvKFrYTdWZDZzyDOtFImSPuTzCRkYLeftGof6jJzSEDxecit2106kDmn
5D+UTHUZMQYg9f8He0MFSj3a/gjeEUnAiTh/hxDtowMlKmDd2qrW10TVLODl
dxdhMBnjOC+1d8nVQbtlvNjhjkLMn9QGlTl05U96Y3Y1tzDJ9DyTpJMqiTvZ
6yOei3NEgfjNIpD3u6D3pU6FtgByo2B9NdoG2VNfxot1FGKjach1TLOEoe97
dDYYb6tY1b9s5yEf1oi3ZNZEcDIeujNl2oVjlVJtcr2rrVLz278bi3Zn3VXs
PED+BGD4n/lSeuUGOm3gfKfv2oquIGJSQPGUE1QGV+mePexQP642Y5S1yrUQ
Fw9WVaPNbsgzzP13WSQk1kQdsmdS7V8/8/GQ4lM7lbVlPte8bX7r5GwB+Sl/
az2WytZVb5cA8YRTwycX4WCADVhdW04v6th3EAfEMXSf2p4Pv/lPGBMPeDBS
XoUJ8vWyXNznJASLpRlVy5UPyhP4zP0AP94OxJMWLen58PludHjjTSKkKNfV
bjPg0AwRB6cPNlygIukYwR5RjuDE7SZB76Flwg79TvqReoN7hz5GgzcJcx2Z
W56vMXmsm0DpYXX1Nc6bJYTWtRWc5Y5wn43Jh3hyXAPLTV0odyD9Yg1haLzk
2d+SKg9vEgtqRiir39pGFc4nZ3siclwh14wRHAWXFy31709aGfZHR7nyPmsR
sDQ0DDiF4ez0pA7J1YdntPKClO7PLncCjgfOSRBrfzJkaRhx1RQjDIW1oxvG
WxTKChiZp0zuMOSekdklVdkxa1Riw/Nv1f5BHVrgIFO6mlcObEvN7slvOq2c
juRPbNTfOB46LFo95BxF3nUhmuQPggHHrmT4iEn0It8bE8KipYIPOybtrja2
mvbaGNwM+g+nv7zY+VrV41fsf3McAoX6Fpxyt0v2fe9ziDSxKMOnkZnhVdUL
nG3bCfZVF6uA3B1KViI5QmAvygjWRuA8EoxJTbMKaeY2gXHLZEINiaVr9Phz
/s25nHOg0G60mRfEMXDPZte2lwaRFre9x2pRW8FnNdoHMpiYGqY3po9vlL0s
zSSl3UVmIkCDKvsy2DWXJjoEiZnSWh4devULigRCKPwLLiUUwyYSEfYf93Bs
3hd6iyddNZPzdATbDIRRSzuVFpO1495hhrfP0ZuSm/CzprAM/cxs8QM/rwsF
EiOBvoNacQ9JMqATxT2bMsidlFio+trp7LKFxcGeCnr0I9/Asv+BJzdyzVYi
WiJ5p5GHmGOYA0jLwfprauey+RJ2QeuCzH/A5bWLtbpl+df23uvt/ymaQFL/
j8uFBnZdBX0RIgw/NwfTX4nmjFG3pXhLJr9XSmjV6QJIJlBZBnTXlyvhlNw0
ASJCYtMHKX6LFQFODvJ/obRMVFvRLtGkm1QGq7meyRaQREVV0AoZwRJhvBwX
y7mYANhGLF4X5YxCgi6s1TJYe8F+LmnZfd4a1CrO9P4vEfAknK5mfQ2bz+bT
fYHEuh8rRzcExyvszNBQZBjeN3GVA7JQ91Z0fNbDqq95Cjk913ygG3VSh6j7
Mb5yXNVj5NbqK3xjlfLLnTXjpHyJP3/Bj5xXsPreJhWmMI0vhmKiC2XSRkIP
QJEtsrx0IDGi1fG1/Pr+El5XVLI1noMZ6ULVmhlhukhlF0gvUF642M+HKkoG
AsxnQf0A4NuRFZimex6vIRvpYY7P4POkpYrZe6XhOBA6M+sLZ3LIjryVr1qL
9tog7pC0YveuK7Gn7S7Idugoy5bSUUXCzn4akzU0rxR1eui+WCV/Blgr7Rjb
LPtFwNmFDnk3VyOf2Y1WcSrTw/IXhdV1xD6TORTBf9et18QaQGHzjkrEkiOE
wOdq2fW9Z4Y5xgLNyPmf94+mz7PQqIlu+SkvPwmS49RZfvquddDXpq4xcClz
J8uEV0KrlOMS//0JNW3iUFqPgHISRpXExPB1g+iObIyJdfgEdUvDhDMzxYF0
JvkwPYBRqxcbEKMG3KuMBYeYSeD1IwuuPs1mgZB238oYNMBDjgWK00a8n3AN
lQXgBdWhLiL6GonyqYXK7JbclpTs7w4Jq36NydTNkqn9/NGldkptNKGBkMub
9tXJAQkczjKFBwxQ7yXkZIfDRQ6cuD25c+4AoasqFCsRQUQcNhpsAKzWuBfr
0TIb1GJGcFr/T1q4m1nxoG3zxLHXYtcgdOBA5G7lEsYv5kuPXC+xOBg1yMZp
a1HSg2wm1lr8NmDS6wol2BiuIudx4Q2ru7JEyokxIifE7dXjboDF7PhE9tAH
a7p6vtKUJj1J+vpebBrF+j1w5utczHQgDomUXLPIGy7i0orl0dVyPbvwh5ys
fbrWkYhLGyW1ou8iv985Lah0qRLRsp6a72atU72zOXd0Ki+4t7bOymvKIq0A
e/T/iNZ4X0uqSiTq4LieN/bqYf4UgK+m7ZSlQPgVOZPNA48YMROVgQeL4ItU
3j0buvIBq6a1VbnVFrDxsa4ZU1kz1k4eBsVcvM48EXJhwlNuw8ETid7PvdLs
FlhDAw1nfMsmNl9JyQZNgC8PtH+a9+1zPoCMKIhhCUXAM11NmpGE5j9WfTfx
VY5LSSkcnBcY4zeJ7czNwsFSq+R/FL3xzSSvBbEMjJTetAyax6qjOLEt6tO9
kqJI9yeZ+PlghJ1P7Z/NEk/I6j6x+3CgB50YkxDpfBHidvT5YOtGb5HKaxWK
a2UzJ0REBwh6FM3g+pcvfZpXq53MiHko7mE4tY2151AflD2XoMsJT3veZ43z
omL5p6qvsd9NO1UZgnjZW5ERLqeJkei+sr93oaRwTgq2JQIw1ySGStFYiIeL
qcBb4Yzed92Qd5uC3ktHSXHiO/FhLTb9h8bFN7GN32p73JcDfT6npo2xPrXI
YzjXpyksNT66QnNbg5dSptpNqz/3VNtXC7sZz2u9nApPHnLh7/LYbbsp27wv
DAxLS0HXPYiW2c5i6FPl9NoyaHn+bP8fq5JOSgbQoZ2upRWquFhpWwUPZamu
st4ooH0iIMFa2hkBXYNF1aq7F5/xHTzHaVaJL6rL58Sc3FyJuYFXZ4TpVMOI
yiRgV1VrH6eLOEx0O91s6eNRxfn+iQZ6aNnNW5ENQUf2N71uP8OgEcP/0Tqq
xg8ty6+jr0lYBMMDKKKz/Zrd/vPB4RbpZGNi/7Q/2+GqIrp1/ePqdotlpOiY
+WAjMo1MmardBZuHAIWkFgZSaNrGhR3LTXrA5NmO55OWQrTRU8r5PtZiRHUj
8zbJxHYNLKvmD0YbXKM2LfYrWcBjX6zGSWdlPIDhOmGVLbmMWjOXmq1YRRXt
lAX2YyPDAuJa1LODbKsF2DNWXTGb6AVb2/Hb1UnvNeHsKWB27tV6M+leeAUt
ALNlP52KNk3vglI8sHH+bmoXVxy8daGkSS2Pb2pLeN4tIrvJM7ZNz56b6odO
xV+LbQGWUlDksFYPQEV9dPswwrrKoSPKMx/PeBFDVrEYVXZEHcO0upYRoVsa
WtCiWhSQnpr4KBm+78HTLeuBcVVuUJGC3ESV9CbJNDoCSPGpyTfe34QcNKoC
Vu12BLurLc/r7oEy4XOuyCZ5WB0gM2bODhNs8tozcxTf9DSAIdqGmx/hj8xX
1fIUX2eNYRBIf38lK45t5bsItktJhOyAOPpeX41a3Dxosw14TmVxUN2lahHT
G+OA1HKJKMQ0vr3IOkDfJf4KTkO4fg+Un9XrE7bWO3DTg8AdXVeYvyWvnvWY
B/U+HWIGzalcP0glQMpgWtXDTeIjtHdmcN8+dNg42yY7VNgJeFnH5TL7wGQu
Ccys0AqMFprf77ncKe3hcSZQaZ4IH1297Uy8mw7sXdSKbiSLgkZc9q2vVZAW
ZqNidlDAXUdZU/Sddx+uodzCOjqzwGGr6sq2ptn2hBtSw29MTPmcuEp3j5++
hFJO6EzDOfDMv8D3q+TDNQNfqcmLvoygeDhxY6YXaAC0o2UaO4d6jvfeVotw
r4kMkElDBddWIzKme18mH7Pe2MjAGFf1yI5A8/ft79k0ADYFeioxVdh4nC6b
NMcM1enJPW3Y7yjqBIXikbE+6ZOTx1KojFUnvOwQZate6IgZ4Axcu/g7hI96
RO4IeB7XycpN5voSIde5QRYZvkcAAW+xK1LDyvrBPcDySeBTgky3SV8ok82z
z1g5GrT27cQ0YtsPQhBx82rJkA4VA7P/SbFPfpcIX84cPEnkE+hV0XClSCHZ
PAh6V3vIpUk8Of1k9G7+lN5nrl7D2NhZxVePRtv5mlUk/n98GbQ0YpcBfx2K
0+Nt8t9+t/PiD3AIMyRuIc0/XPosS4wtVLbsu4XIKUtAVZAgyC733UVmF6wZ
8Zy2aRlvSfluIuNk7klS0jio2/7fYYIWcHgD0WC8ghlgsWCWDthms7sgJlxG
HlXtwbwD8XZVFERsDlHBzSoNkac1KzzYFmHrStFsEGl/s/D6gpD0H/8/W35V
gILZyNbfUfSvDbIjelTVpt3W2IqX+ZdzfYCUn1rp2hASzPgvYkjt6smZRwcj
rvzMXBOzFKSK+9wy9fL+bjwnHxuGFmtjuX0HNkKO+JTojGDPYMQAl56LCc42
pBpoRaEzXDeSLt2JEuvIgnzgKBVL+/tctGhme96MKIAMyfr9UEukiTp1whZJ
QqybDcrwcY2JgcvaEs0FT27FPwI6QDX/Hc7DPf5c73KVAosxfoZ/QPqFSL3r
HzhSWX4V0XdJ3A64Jo1RtrALdTlgUUvPPdPk3lmcIxDWhPu6g4cCs57o9OUq
xu4nkXwtGeJx6s/ENWkeIJPkvzuuQZzSQvs3bxhF6z6Eqq9tjXYba8O7U/+u
8CsXdU8Si7/6YZ0NMnt6Bhho274y9GznAiHhhL2Dpv9lOnUooYFhxxMUNiTn
VhsFLXoUuP4kQTbEeqo5mCkkEg8bXemEM7rHZkvy9uoa8kdwub65Xy0iC1QH
Vvq7iC/2YcBZCzHENxCvD0YQ/L/hICLR50cyHnM9eNlfOdlao1EGOuyIcJw6
kIX4TFLdIMCnFwOa/AwrctlzVVmen+mJYnIiIGK34aeDHqx1GJ0gMeS7rz0G
T95jhZz1vgX4+l3AY6BZS9hMt3dLkFw+lOLe5Uv92uoVTf1SikdxuFZRZbb2
zRlQUPh4ww+0H2B+V/uTkRFgCGuXNtVrMg/146wpHLSDwSYOBpC1e4MhjdL+
w+vQX4k0BgSANPCEih+QonSgcVdcV9dF9HCbSygtcA2yPxY2LJQjOxekRpIt
ryGgdC7HaItjEgnAoksrzNDF+Y5DTPAekU+dq7vVjwykDq8p0j/Zx/SgC7v4
kXrPyY1jsJDtmRNG91RBV9gVFe9fGbpwXnWHeR2IpWHhgDgQsEkUVo/MTYip
px+oB7RYBVLIrF2zTJlDbbKRK9KzVfLF4v9qEMv1IgOeAHwH8Fut0ER1Qt9g
A2JVjPSUI4le6fCVyhPcwGG5GZ6WbZZb5tv+kqQ0uRSia+7YZTw6XNaU8dDX
lsX1AGMIYCyJaJVu1QixNuyLmsPY0GQBXWgfqhNWkAnZVI+euhKYavgFTIEX
sqtyhIO4IibgDFiaZgqUfCDNg8i9CXFgqyDEEdlbH05zMTAHB34gsopnOudp
S0mfV5LSTECOnIsGjtBs9hd0XyI2Ovf4LpHT9IOb02UpS1C5j3HMpqYgCg2q
NZkAuHo54Tyu5vjRG4tvX6ySPpxoYgQAW/7+pETKSgot3NOzfS01wPP3IZtE
7UDhGMnEiSFsPBqcQd4/lFhwd2aJVTh7ZZmI+tT/quk8ROvulCs5p5dMHvpr
nAwBAHTK3qhFwD0uND/v5wzLF/Tq13czPJJvnQ+eQn6CFu0ZaVNeb9SUizZU
DiN1ILA1sEBk6ypRPCcww7KwxVpeYZrgOUSd1TDfHpnifv5yN1a7Y9Ql5sVd
mXWIlJskgmxqgDoCihSi/+jQbFual0pwad6DeOTQ+2hYXNQMWUMJMjwflQg+
Xmi+x3hPcAtovgpp86neaIoNws7QgdNjcq4E1ICh0mHKxB+T2uKoD8awdlaI
zTgOETkxU4p/pTgnVxl4oz4rM/yunDvNNdZubj9TIngcBGM5dKVruBP1ptjo
5tP0/OudcT14AyFK/ck0W5GhPDmBuLJdmjGrs3reeO1bTV6XgYRzt07pqvFC
QbkMVORSffHNAa6SC56MbDHPJDQ0gEfXFI3rPoS7Bo2UF+pE0QJ9kfnZLACW
pFL5NDqAZWNhSRWnk9AZjMho2plTCZ3fldyDVOzpdWVCMyn3mZDbQzm/uPzG
DGvhPqb4RiOzzMw2OHBehvq9eX//kQkycipVgd2JrHDenxlD71vsNoVfjy4h
EyJbg5i626svEB6mDbrroGo+3ssy+xaUhlLjYrkUp1xFtAX1+W6hcZnzz/0e
fEcTk3A612TDBBHslOtOmdospAScJAO7KtckWp5a7SYNNQHSPnFwgj49+Pm0
4GNW9V0NvIoZXJHh6eYBz3YZ4dd90AWGQar5gywFbu3dp88pF4S+Jj0PzUSH
+QVcx9Wo+znrokVOZxi0USqznVQYOLsHwUOnfezN4cPXvLF8vI2tS5fI9h/i
bOWAoqQnNyHvV7NDZ5n5lNNJZmuo4V+R0bQZQyMnoGHH3JR3xttT47P0h7IS
TgGw/dM5HcxAhJMgeksDg8AvcvBqRbBEMnHy5NE7f6CISzwBJUuD40d0qA5d
VUT+KxK7vKlK3O7ksRI7csIMv7irRzuX9AXGIb5oN8hKhsWGMoAzrg9UD9Ju
IKKQc4iX7jROWMfbIS25dVNLegBfxpLdN/UC9cIDjXQF7cHc8m8Ou0R7cdb0
5R/c9UNTNQ4zPP3iZAvMeyFZPjQt/olcMcf4KvAvdRaZN6NvbgtPOEMWG54r
lrGeWo3CLLF++4w97PD9pf+gd4NKhbX400KIgQABS9P+s/lHwkTGUZdRCkDO
KiXIdt9/ZUsynzusdcXbna7uFCHZOWYlqATJShbK0AsvKc4X9Brre8LZW2AE
5ZoAjVjzhp+1Yk2bx8NGEHLobHQ4UfW6nqDnQsqyo6dUJPTlwMQYh8jdEE59
qygXb9kjH748XFw861lN4/7dmrb59mNGb10wmgWh8aiywFPDZq7DY0yj7gh0
nU3cjOIr2W7Xfl9v8U5sMWP710GIUeG0LxKa2+kZdDyFoZa3BuEBHzdXGsyK
k+QQ1iyhxUg7aqVsPcL3MRAsqASJNIkKRmrm+7c34ja8fMSUFq4suz7KWTk5
etL7YKTIF01JgEPHyidyon/KGisG0ZGm4tyIJnbndkTJAvWoAU6oFhB+XZ9n
GKsRvcdu73+ZJmCbbCHfK9pLTxi+V6nJjXhaPO2gh7W7aISiZTM5QMN9SvXe
VgnuHcDizD3IWu32IjgOylKYNs6hOnB9Li07mucYRlUgtt6l9Q5r+EMUfAxM
vSgJzrgtFAPa2ckKE9GAWwn+KlJGN6YZtnjDj6PLcrvF83067ZoFcRYyFE13
PUr5qXzIPEkeWKklhtjhZ/W9oGsIxVSx2xZauy9aPrb9aVh0Z9h/h3wu57WY
vVnPg3T/H/13D9j7JTWf0NXP6ij7zHAzJzCH/Bf3U/aOzBi1eWo0wPv8lvZn
xiTVSEnkqRglsbnqwDi27zh60aGJN6cdW6razwSS+M95Z8lXZfFQlnkrh7ps
PrK0bRe66Ti6m3I19JniMeqj76+sBYmM6lPTQ8EkYeXaUUKCbtKoDqWEo9/x
Flwk68NxBo3VzHW6HgwWlGChGG2LEJEL0StTQ9p0tNKNhLk2zDN7Yrvywzy6
NfScs/8mpaccgyLZgkOlUW2Em+Ao3eoh49Cclp1NuMSeUOVPTFP9pKJJZOL7
1C+dQiSKv7MkkP0O+7e+7JQyvUj2Hn6058HcxP9yld6oLNuwUwnILtvRej+B
Jbth9/FY/zHIBm7SLz8dj2wtsY58zbTqibQrZnYfAdSY3zRa4Oce+0CXmVXR
djqz5ZxF2j8YomH9Yn40nJozwAYE/F6ADkKNToqR95V5Wb/SUnk6pgknBRxC
DmF9JScNoVWrex4oRnRgK3UNstZRy5+ZS4rvdzJvg4FMURjFwDs4+XIertCz
gPAoTKiCtCCdN7hlmBL0HenRJQI5Etzz6dtZ0nIkmjDCqRhkLIDGeubFSijY
hKfDliHGNT0ta6KKGcA1kwsOxrXWEVwbvEpcPZV7sSVSIAaQ2w2t2ISH2NB5
5RpNe+gD2H7aLkHx5MD3Opb0kPb1zXpsk0GILZOt3AV3cWLejSoy7cuZpOg0
PjUndEnsOZGSAhSUhd66aUgeK0sHMO9wj3bwgC8SEG6XmKO5SUUxp1I4Xy3w
Uit3qOXbX9HkoET6n4lIWIVPU9WHhtNDk0BrC7ySVP+Bf2pFbuAesJfwxjXd
Fe9cPavG7Ii9E8XUeKkRaAAehyKKvkUt4EF/3c67hbxU0O2gKimvE1KzHo50
zhcSqIhL+1wY2P5bZzD7iQPIMmvmh2qnwUIhZASE2upWJT9yf/KcMYWcrjeH
StKufR0NOBA8Mqf5+OcEEuDf9b9DpGlvwfuF1Hz0fZoNs3cAofH0xjdI99IR
XNOexH2mgbJc8XPbPrGdvzD4Jd9aITsq+ZZKNtocW7i43iBdxDzfrUwxXgte
CuccHpWHrM0S0uxU/rTFT56NQ8LvaARFop4PfUHmCze5SK/WCVNJvSMECHJI
AfseWaIEZ1HijJ/6lNouVGsIt6kYDhfpmQ29JUa49zb0bbsiQMVQXTPfFVHz
IoOgqwJS+ehU0MXYDctGtjUmj1agSA8yYSyUpiE9jiWK9soN0fsw7Tsyuvqn
sG1dkRCiFWKOtZ6L54csumURKzAr2lEk9lSUJBzyavbdJtC1kcvXljR8+v2y
47uUBYB9qntYkEyk067YQs4b6s0NeGPdlAsenIxE/ybFRR1HoRhp0sN11gu2
RshwbklMOmuE1t/xcE6Pq3peqXjQprVu/HQnBSwnqbNrTVVlyA7xUPn0bP4s
or0/U/nVNQza/ftdk3KYOTAur8pP/LIw9UOJ+aAerdSG928liTCi30fxsAHc
brANocvUKVXU5rEHLoQ4FifmgcC9KWE1kqpnHlxa3K7zVgCukVuoLfwVm8K0
ZdZpFEIaLaFMa0SAUhg2141rNi8ZYJ0xcafSAg3VXJencx5b9OdI+5Rwpp22
cYSCGOC99KNvhfUFInezZElD2W8evfPSLqOzaDxPZR5X8zUzSEntJwiSRIdE
46Z3zzHH8X7tb6w+v/lyBRm5P6L7auJi8Xj8YeqHluGTZ25XpLcLRsmZFmNU
kDDXZgGs+QfvJ1HBf7Jw7YlOZA3LKnm44QA3xpzOHrwrJA2o3jlGG0iehoPQ
mPYmaVv5h7ZNU5eBz6m/jwkQY8vGY7V897TLpgql3KWXRNsgIFTKKwFZxhVi
f/P12apDijRHcA6+U/6hVgbnIq1tko8BBnRt1owb3KkjG59ipCqFPdphoz4U
fJM7Rx8cSVEyn7JkWjUJGVl7LQM6m4dG8PjfOf2aBbq5ebBTQOssvZuqfV7T
gJghXroRQmSDy2efA06WBh6xtXhO6ddCRSDb+cui47u9ends5L8KSN1BKs8x
49RDemyr+qU611n3YHlX+ENLVwIW62N0plRJaFRUGFfiWDZvqMsZvIXwbp1X
Bu/gwyB2R+lhZPsueFM/knnfupdGZWJxlvu3FwhDmtvy0tvfkBO8FPX0qde6
oQ85XhWm7DOHVROEkr+FkgUgPwCgFiNVHspsCELR8Wl/mXLcxGyS8+83Mzh6
c6DElSrwTT2VZE5NFoCJep461yPL7OIsCw/fVRNKEVlxyXCTb1uiE5b72CBJ
yFfoM/HKU9zBnA0TK3rH/pUZBFMU92N+Le5ewtrpB/P+8x00TaZgZhMkyV9Y
hkXQtt70tIftmu2tIyBLyUHeTMPkEQlRme+NJmU5BCaWJ1Iw5bgtuAMILwj0
mD3phK+Os1ckPGXQOkwh8t7B4FI2HKNCy/GCS8vpnAngAhPd7lyxrXwmgkIG
bq49RFOdXjJGuuXIy698uE8TqI+0WFnkCE+6OiBq6Ejm9kw2IChwpp/ejfml
+H47Pu811O6TZc1hwlWyoC46fHgu9euaGrdSgpLVxko9ULWYPgTYVuPfFkCu
OCPIHqZ7l22yvvJJYisse/fqixKK8t7Oy0y1C8SCnWmsmmCMwAcdEFn8gmqM
gU265sktgDlvIv9kGy0ENLo6KEs9F9Bt9jBDfwCq0FZynJFw4+hzTRIy5a4v
AuG+RpWjmyFyChlIorKNewPEPmCTW0Q0zKUm9/eITQvqbdi+JX89SpGT570S
fHxJ4bmijpMPvMnyzE3wMb5Jk441I+1kn/Ky13m2UIZuyhai3KGCtKTlI3B7
v1zOP6yrLt/ald7lGX9/1cQm+KGe0XjaS7fh/tPgN+hU/8+FUubD2s4ammAw
/T51D/olY56g1k/P0cDtcxSloEbH1t8W+cxmKxVygw6hAHZFU9KfMjXZS+FD
8/w6W7pKg4mDg3mfE7/CpFl2vJv6q2DwbbJexoQcgw17GU7Ebbr7CVcWf2pc
cqZUX+WEnKLij6rV4DlNOOaia8Wi2bK79C6KrgXSXSYjfklQqJPC8fkJI8oQ
CsO9ZUD8ruMw8vLnaSZAps3haklxbVkWNBJe3GTUDZ7Ppmw7z4dNaEDqlD/s
IqRlQj/uFQ5qfeGT2axXPfwl2DdoUVgB3ICMQSRqYI7aponcIraC5gjngMSc
va55cMXbcWHonmSunXNJkzzd9h2FdcXuqwBMTXLz2/P/W+MjaoV6CboxQQ/M
360zVx5ZdHbKEyrHjF0SWMR8v1q1YfiA5hymiU6SOpmj2LuFcUdv+usJ6SBh
2c21AyTyR30+lS9udAlp0DL2thMAu1UmYjPSHAi2Pg+n8OtqV+K11CU1gnpY
f4khNbOfAnjejJbVRowdZijfXMv0sMcbWRdeZCjNH9XNhPuF0qoUVWSKnvzg
8hsKSC8u9sY3r/AhkR55CtLtcHsjxp0gVzf01ESqbsAg0DjtUsM8Uadz+Jf3
oi70Y2+iROt6Z/1EF35SQXnDTNK/zur75RMGuxGj0E0lRlSt2PwkJGF+2swb
AEfimWE+yRsUjSQrrDUGeBKqSX58cXqQbqDlzw/vEcaVwNIcFZQmuzMG2xw1
O+MBrpibBQd4XhbLkX4gacnBrMvLFtOcFKzeMWNqdlbIYC61ELei869mXo8B
Kr9RLQMAbWprBkaCgakG7o2JBeiyF3Dxgj9G5o9uvKuZnn9nmtygEwXVF8Vm
7Ktcs6LMglCEA9OolB+bSKb7stzfaFDmK5fANOhEFqCwuZ7zAKL888hMP9ic
Shw1ahoP47v2pGE97Zr6l/x+moFX6AElrvSFPyIjJCiHgiWTvvNzRIZ9RNxQ
aU8g4EzNYwcNvPVUbtCxd4zvCMSLHZayI1yx1UboyAc/aKcDdEROKDjb+uus
q87IsUdgtXnmucB5r/aXKn0nirEJ0tzpYRtKhSBnPrGnBIqX/xD7R9m8+Z+P
kHegftzTVfZGJ4KSO0d5WYliJdnkfyE7k6P4s9ZguUNulh8SbP74fGv19jTr
UNFjlVa7o3Wfi3w+/ej7RAZpck8b39o4kuTiJGJZ3keN4uNMyb/DS4IXigN1
RXgrCfqRw82Vfdb6SHVXvSvhme9IEH5m56ojbIzGpQF5lrnpE04GVCLSP2Sb
6IC4hFCsp/E/Rxczn/9SCfKOMEqp/mVJdAsX18W7jmLOw8sMM4xq6pgZiHwY
mIcm81I3q1stfu1r8DtgfuTcQgKMcIocvqkQPt7AEp6FxEW9xZp8iOJ4qeS9
XW58sb2eQTFED4C8XHaY+oSWJ9nSmpBRJgJ0zDDBf/g5ORZTXOXbpq99akFc
zl1SAppi8BrYc8AeTAB0oITEmVJqONYhMebzsAgldGRjCL8ScjktSbmzZDcI
FNkvPpJbXnzhYNtBoA+l63IZIEzu/Kg2o/8HZ40bFTcGn98H0Pj0ygKk4Jo4
NCov9MzC/or9sIhFuzGfCzCueNyoA8RgghBIVLRMJxk1j/w8X0YM3PNdl+gO
LPhbaeVgic2ECXwOKgjjmxKlfSff82RoJx4cOqKx3xMTf+HLTHtUZ0SkFLQw
slR/JucKlsZGKRiqmr8q0SHmlu7h3CEVv8uOF0RKP5MBigNbDBE4R4GBNsfL
F6k2khlCvHrPhAGjNVWd5W1FZP5DxWBnm8ABFN9sxErlI6r7U0O5lRLm86gJ
/2taEiS85uF6ORyy+14oRzZDVh9OLdQ6NFrLMZtDA030hmxRg2R+GnPiFZca
TSvBHNhwILfB6JaIDOofQAuDhcq3LJl5axQjZTNP+VsRhA5DLXjpUmhBA/Ll
SGv1EsR3UdWq9eM5jSBCzb22NSIMMMWgQ6CEzCUudx/HR/49EQmyEmx5Pp1Y
XD0sHK6odkKYUnFFmot+E2czUoI7rUMiDDo2O+1cTyZSxwe2dDGOzgy1yyDU
0Agp0mPspESLD+frZxL+kiICpWeovVPGqm6ZjuH+we+NivqVTkcxT7NJoPJ0
1Ei/yFXX7unQ7n17BOF93pblXHrWWTb4t3NepwTExRhNGXZ/A08CUoie1G8v
nN9zxOEV5shpIpUTftCsi5p2+Um8oR95KnNtOizgF0KoTVsislDK0mH+rQmc
eARMQm+9QysZcb0yrMJ4+Ib4qUI9mnskXZ64ZPwtyipv1fvABG18+jIP/kpV
RJSBvyxGsENvgy0jR+w8/o19wpNKGNd5WXOwiZH7qtbXgx5b2KezQwtcFxJe
zlVbidnb+brKRr/cAJeEbBka7NWSs4aPOucpXPB5EB03FEwcWrvksc6T8Fx6
MK9dqcP9B3WOAD048nOXL35WRT6adwTBbv3l9A0rsthCoRrSfrrmpMfoVX1H
1tKvqI+5kHksBPkRYOpyKxXGUXT+v8fXwLY0Php9w76b3pzNc2OUHN0lRywt
Ve+GdYLCp6L725MtYTb6/9OMMUT+xZubZIngalsAjSFQhGMuyeuqpmn0BNTz
xFzS7Eqe+mdCFCZbd30gTSgjurLX8KkTOfreCOOUwmZjQfss32snYbp1mXPc
5sljz5d4uOVQ/LDGyHVrqKlCl7SLYMx+P8HigK2cqUn+F398xOmgmr6+MmVW
7unYqpVTBItFgqdjRTe9CqTjlcIaDVoe+iobMVvJGUI+rTe+CSitaDHSnmg8
WVfkZqij1wfdW3ojt0bagxMq0hHzo8+hscWzlVEh45ceOVS1A5Jn+ylClC8+
6gY/KxRO1eLkSRofor+/jf8axOwaFMjuhY2lonwU2ubPjtYEylslE+C2WFD5
hU+FjXJw8r8+W6MkkrPb948AC0Bbr7fsa8VD5pbYkIoBfrZr9UlB+q1oyLVZ
RRyRVhAKzu4SIrlUAX5WrTwG3yDeaTkyvhi/hGDql/6xlpuFHqnB5VLR8hHu
hAolMxjDL8zcje7m/Dn9LFLxeb6HQ0Q+mHXA620e1ZSJlqkVcxEJJ88H/8KL
ZXqAZ5MkUAtOrpoKThe3VQyaGtsjlyO79CJ3Y0avinr537FKxqvOdyC+/NEd
BI7t5q6Aw8gEY0NZrtCCa584hJC4AS2mAy1a/Xs5gQ1IkyFXg6w6ivBoctNS
JZ6JOWSCdaUiJwIEXQBpQWxt2EaWJIyR795Y3EiMql432H+jq8yI9ChtTqZQ
vl+19yPi34DAVJTGXwoqTdpxr0zL3jGbQb5M+CaLjCEHARHvjp4UeIP9ZaoF
hF9LlkeLj8ugJEkhECG2j8n+D5XSDdCX0X4F2GTXR0YZ+j6KJ9HHdhfCV1f2
0BBqF2qKg1vhHRyV4NeyuL1zM8CkjQ3YDfyTHZQmmBtQrbyaZXSWHL28FtoG
9Am7L7sLMUZA+1EtXE/oA0pvQHbgKE1E041PNVkoHnR6iZglI08oy33GL88o
DVCIRoneYS6UwGzSIQI0rBHlRGzdgOcz/l98E5haJ76MJKPAZFPPrq77hsMQ
MpH+P1fRq31rp90dIcOI6hkURWPYgiZh/ytk4OQ5gStPCGSRq5BPZU4J3FOF
z1WA6P5rmK2Wga8SB0fcA4d54szrmyq598Yyt/O6s0vTEzPe+KaLUk54tOyK
/dDqzek96s8cGTdfidOOvqUfagbSBgEKFQ7O5oUeik7FCDh5vGBDL644I5ap
vljd0Wnhq0mAV4m7XX4TvuGckdgBxYhqkVH2F/so31/nPlditLhYZH8sendV
r6UuXjV6DNVZJ09ceAFpFiYiip+KCK2F9hRDtQw0pYZvdMQ5Uqrw/yAQo8nf
0ST+yWTqiCFjNDnVGer10DUgLVIhC0+UTIK48y2X9CvFa8OizZmwNrDob9dV
t4tGQFrA0IwOjS9tHabGT8OZGNfrgjTuDS0ZZmqbU65oQ8rvr20do3bwnlRO
TeBB7Cb+W7ks63kSuxacPwJSUHAfXtmG+Jx4fUa+ku8Ri/2ma4WSE+68VGdD
a5U49AYltj4GWU99UhWsLgl2N1CXWfq6BZ/Tb9Zg8xh5+LBAD3jL3A3sObDK
990Wm0D33mwsAybTjMsask6SZZvg/0U1kbICGmvgZzPq/d46UdesEd3vm6E2
zTLXFqizz+eJyG/p5oG9Vxo7OOAS836omTli4T/qbcqihK/xnHpR0DrLMLgj
BIefWU+JWNdEzbERoet5Gl7tZcBzsANUsizYJjw52Jgdo9XDDSdS5lECiEey
bAjW7bDZeDf52FXfIy4dNdnqumOcdOcgDazJIt7v0PDCWv5c41ckXAyrxHEI
GFCbVFB+78LUsRWCekFkE4vhEJX3iv+OnMYerf3Ve9kiLCE7prS3k6kwb9ib
dXugu1M75XkLLT1uku0ZPzt1JFvihJcMONJRnUQqQocMROD4xHTmigLmxuI8
DCRVpidJIXtFlo2pNDqHLpIE4WC5X6p2EaA/l13+iTGpyGP3CDydXcR3vkOa
lPhuigJGb0ov7eErDVjMvJ8pwEJrUOVHbFURGfV/6EZg4uXpMDTAo3LhqmFD
Oiee0CIwQZaOTiSFGtqQRmCDg6KgXS3L7OZd/rB/bth/TXgXKG+eGYiTb2Xv
FKwcNtcVtH0hj3fdY36108c6CrtDRQtUm8XOM3mbcxJL96YrjH8tblbt5fLy
hhLzyWXnqoYV0Mjuz+7O/nOVV3SAi1yACqneBMAN0r21xoBn2CRUIqohon4b
7rec+EOQ4RK6iQYNoK02dvpymJ7eN5VjY6kYNPmcM/xL0IZzKU4cMGZtwcRN
BkYId/l0awTBUC6ZJuZr3scWYmyKnwBYl+ohHMr2SBS3yfNaBtuWlGKYJca3
LkMnC67ViA6NBhbS/zyXQny1cnox2nhw6aM6GSbSeRhuFJc9n8tS3ew7d1Ah
Jk+nbo3uHrCqyPoqjj/wtu2KmJyHz/b4wLFROjez8mklW1SsMr4CJ8fFwBu8
cZKwGe0pN2VdZQbQSIO1nZ4C+9leJinCg/ms+e3JWW/mR5eL0fFdS5SsFgvn
087WshWio574HwmkRLnnCaHPrPk0QUfdVJ8AywqTK1hAr6+hX7KR3oBRwYBp
wVQ6G8EuX2XeUgl9LCH49qFUtvLq564nqHBRddC1CqjR0GUr9OmiCw4VbrfM
2QW6LA9pe4oVR5Q88GE09CG3frlJULjt7XJQY80oYTyXoh5FB74DHjmCo9oi
5lCvunp1zTn0PqvlVwX3PCLmtDue/lIB2ACFCqwMoOFX+eYnwIrU46psou2P
3gj1G1sOfDbqBrX7sLA0qpHMuKbRq8xsZOuLWUJmdw0H26gPDpkZBTceLR2l
XMTN93H+utJ51A1LDvMQdsF6336Ux/GW7EYy1UwNCTCYvBbZdxEqty91yXER
SMD0wGyquxoRBKNIL5J1gRBB1+QnA1zAmHpY2Na9yf51upjpGPQMXjI+bnSr
MScpowbtdRdM5j3uHz2lQWXUmuNrYNhi9nfQaFERhTsPxxpROyAclupHvJQl
+QmVp33ZDVS76QEVYKeMFUCj/vBkvdFyL4xlmIV4lUGI0/HU5w6CwRQs0DbV
VIpIgEKkk/gl0L+psGhsd4ekFevxpBddwbDW76mJeV3HZi+GK26xQ0hlAmtf
X0iuq+NxReoQwGFeT4fKFVUFQJbn+9bCsNKtUIkiYnFBd1TycCxSOwU3EQmc
LaXLUGhCPC0KwzVJ0Pqn5fRO1jIYtTTmQmIiUR6tW/PAg9e1YQHlOD42mII3
5rJsKKtgjt0HJk13z3BlcJdSbGHir2o3zi06w93pp52jhN9tqfJ5nVrltGKc
SEqYo75zh/LKPshA5nsJXr8546N8g5VXh/evpsyScY3JbDjGGFYMH0QCLdlr
m5+DiECplwuJ5yGRa3vpBml83uoeQ7+Hd/NefHE5bgqYV2prDklkKs58OtgQ
1EVVrJuZUxXrWgP24gBy2QdPyx7Mm358vwikNF1CnWlczSp4UC6uleLnk3iU
BLe54Gre3hYoO6hvsQLdaRtImpT+zOZOkQ9mYaxvlfqpPDq8mHDFl1aMd3vC
1Xbjkffp+uj1qbeNytexZUyQzD7IVwZ64CHk9pe/AGb7pCATnhPHWgsHO/zj
l4jO3fbc+cyNga72YWp6THG/KDPbwe8FUhg5iTWtUOmqgIeu5Gjzue8p0gna
pWe2BUEhp+r12zvj5g2KvbnbCABnDbSOD/XHfUb4C5rucZ4DdhMNa1SZB0g2
iJnQavKZsw4rVktPk7/KUDBy8ylq/FoVhlUv/HUzRlJHrlAtTtqwOh76uHbx
L+PEP2UyRRr2ywY7PAwJGRimyauXtGkRk+lDjdqqMYhSo5jxx3ySxW4nUBIb
VJlTX518zqdyDtM7+nUM3XyObviWPlRq5lLqlQD9zoV4JRlf4drK7cd6Huws
pwn2Am9hincW7AdPN4Gamdu2Ig2cIEibluBAQzTmYRDOBLS21uu7WU63sMgV
WzhpSQ0X/hZlKkzkLqYN0BaxYzr//QAiC5QgSg5+2JLvM77vBlOxTgflurRN
C4/VTMSSvxMSX9NMIyRoN3QSi2yTXetimd3ZSLHk9b8n66O7aTIZAUYUmZrk
+K6CR4OaGO/CzUu1vfNO0XH55rcX+ZAlglwQfF16P4SIvyMatPeVg7K/8kof
vfD5bRs7Z6X9y5moYcxHdVWeZweiJiM8QCLUk5TiHSJNh6K3hPL+u/H/NSHu
FWiqQ2KefXhLYcLPZpyTOWzz5GIHqaJ7CDpQtEN3GGPn8c/tlaYmnbVqFP8w
HsrnxMJPM7pdNahliKbDiIGSZmJzpCnau4MmpoCF/WzS6m0MRfRNvn7kcisc
0sL4Mwh83la+umk36+k+GfxnWuUp5f5XVkSqD4KbNh+95k6/ATzuDj8sbqas
bzUoIDGMcCVw4VDjGdPrOiOlNDTP30IcsBdGg9oBdSUie13sA71eVOdzvEsc
iIhvhFPIJVtxqDLOEdwRXvnWnJw4UG79QeDD6hNsDL+5N7pR/xW6PckwsKOd
LyLd6AlrqkQgwPXE5pd3d0ErMnzco6eejlxRPn3LGFQOTJRqdnmhbtSVTLve
IgR6aa5WiUeIuq7UMv5LQNwIesb3SaB08xrh/3RRzqek9XZ1HNpHCzn11raJ
aBmu+bqwlYLJl7oY4MEJHGb/F+wKqHRjh/gDp+o9uckS9Lc0zk7G697561f6
4nKH+KjzBxdRcc52lBiQBPGmEmAcinI7iwUzh4BmD3wZW9i3bXELYA7ayq8x
oSHgVvT1UMpykRk6iYwx7mW0zNpPSjmGIOl01tyWAdc+2SyWX/Wf5UbV2FDa
uiiiDxkpvmy0GbYNCepVc0NA47YZsyI+RLIAteVXc2E5STIXj/ZUct7Y3A+q
RIlpJVFfpcEw7JtlAq1mwELLB3/pXMoBoL2dNJP+kTqqejUFym8hvVHamX8T
PKhUBG1wEGj0MrrgW3LMdJkpo8N01s8AcA4lY0NFn1XJ3yU+7UjjEAaB6SBO
OyJ7DoShZBpnPYyeP4B/hXTF36+E5cxD10gNLzPamIy7HMVvfkhbzes39IPV
Um32zcEOHvZse0jYUrKfQOhOGlDQF0L2Pv535uzXCzNYMgS99C9rV/6c4o8W
Mo4c3uoKtK23ed2m0AsGOm2sHSIt1TXaDiueS2ZZ7muyzwrXnj/OjKpa3zsI
p9wdoZkERDVX3s4dUUo6iHxcZlkt0xUNuSFnEANVomkWCcgo+PC8aOBexdgd
J5gDFv/sICx9VNCN9fh8M1XffP1oRCcqy/+UURynTdXkPfbm9m6bcJju9Lis
CiglDCMCkqV2vGxiPnvNSXmeIs8Wpht03uSW2S2wDU3ukynHINxLI51FnayL
kl7Kbx1BBJJAJHSKjnOpK+GIUeiXefF+dwIskr/N1H/zdwkwuBE9mRNLoN0l
lG3LvsBZP8uVW7Fp5zO/7k7RyYuMg1/f7nJrxXp9/7tRIdHAbLODjMKCEXFT
Pmx+LE1Aka3+5ARRu7WFfaIrhGTLZbSe9sLBKABFpnY6EhtgUeh+LlFYm+9w
/3YRLQ8y33Yi7FEMB4I02KzqdaVYhP/u/kZsG6UbH5cYE6F0++LoYNLZyDwj
/IlPyCcSRQm+xVmMMQvatIUbhxSYIK2wX+k6HuzlgqjS7q5UiQLy2iBrPHeA
Y1sceAbaGo1SzwTpj3pXxrfrOy8eq+CKpzKXKKWGUZ1Mdd1lanlOeGSeG4f6
gMKudHOMyr9xwRTXuUhCU/kkQD6wyU7wFgF1N2AGnxEMFwXgimeY2qy+4DRR
gjTMDtNpJWRWPNcPGPNwEuTLo2v9u3SGy0Q6eOQzr9RWpSnVwOCE7VbS1VqF
TGCmUWP+hNfOtFRDe5M5QgdzZgsMxVolbJ/YmjLmAYPdrX5Lc7ZXKcEihdmT
aFF8Kyl++DIzUZCTKtdlxdERife4ScJPjHS8SpHTgT5OOoH0vyEwbZgja3SQ
H6oPboQiirlXwGLGaEO7drtVOmiupIvihrOrT7RT1I28VWY1du8euqsVFRkE
tL8lVujf5hQfSHHwe2i02/6Tc6i/rCcQoA+JpNDSKQtUMvDuL4V0d24hB1t+
uoWYcqC9CxEVsvgl5OTquu2FD5x4vwN6FWr7dYWEwxUgUWmEhEQNn4QzvSm2
Yw/c4GcWQ1pqC6F4j2um/+Y2jtly9Y9OVXPh39UE0XeGbCAhmJCVpRVt1F+n
3m8qSQdAEzYj6NjeVw1TaMN8llX7Zy5YWN7pTo467sq/m0r0gdOhArTF7ojQ
uqis8K36dn6dzgvAqFzrs581l6yrDsWAtVE71iN7WxcrNuVz2DgNc8mUP8k0
RlcH+0Go9CwBGBjHe72KOGnQKsUGITeLSU1tFjzsPQiPRDki3lPry5zS9t3c
890xLqfCPAnzBeQfg4sNaWohcAbI4wwdjhj+Kxx3skQvZ5eb6oQR9ZpjKx7/
076nTOln6RHhDmmOqUffFJsCXdVd2SjCzXndThKZLhRUGJXV2o/0LwIGscIN
NArp0z+vLRja5XXoMkrYR4lncK02uS1UJvqxoXCWbg75e07uWugiKl36I2/u
hWfIVhG2jfy5xAyqmQ26IJWDoQ2hI4RI7VC91xRVP/LBP0N1NT2XuYYsfU9w
E3G3n71gpWxVdq+hpnPF+8huXCdJecqZgKZmpGXLOsCIHwKDRidifPNKhTeC
nfDnXqS4lRggBdyK1qAWtxlRAC0DNfkHMkgS/C2bc2bRTkS4Bk54CV3C/G2M
S+t+RykQsGWef4/SAoJV/bN96x6OI4szOFyL+w4LBaBA9Y9l4uu4E78XYy29
2Pl/SIvVI/i/buAZIteeJgRUg6SXC9eQoaH0yuJgSqhq210Z5DKu/coblq1t
l+mo29U3b1Zgys4QNhlH9EDkcX9HoYFiSo8T+vEIKczF6Z6H9hI7pBj0L05X
M/XyLKOMbshH2/9L0y5uY/gwruAiN06Jr8zZclXPCTu8F5dhlkJ7VeflzjZe
LgZoLa6pOKvszWftgNWY0ri3X/PzOSXT27oV7RffTNyFepR836OkkKP2IsMA
c0k+JNd39ushJBHUTxzDSfg8Fc3svDUryJrikO96+RuRwdML0HJRZmPpziML
fpEMS6Q2WDZKdQZqZnb35yS6ZnY+MO5tzfqWVFM6rtWqoTWEPKBqytd5QrUF
zxDbcXHmNzn2Nfq03H8f1bHaJGfcvwZl6bGAwpjDO9d2UzWJZ/IQ9Yjqa8Es
OJvyZ9Vs+YyZl3rjxhYensdZtKAy9x1eRdnOLsPo7HSYWEPxVQuwS1AiEAhF
jXE8uk4lKthkdrVnZ87TqIXvaHASqQZzXAjzgVKUw0fX8L9nXoGJx5Q3ZY4n
cCkaAK4Lzg0/3HHbk2L/EBSojL0c8Lh8Q4Sed1Y2G2KcivxTWCAK4VITrjwh
1r/MEZmoiyEF3z9R80S7ajRPb2l0dcmgFSj9sIgwBp2P70ldDa2UG36Ohjd+
xSCwwZOjgsdE2cszRNLtVjfDA0vMR6MviSeDeKFXtxt02m6p+DB1T9YvxWMa
Gl4lGSBEEccp4T70/LDEy5v30f2LB9UW/xmLIv0yGO1qu7WPMnuhhLzSQq1k
IqnGY+o1zEZw5nsAEYd2rkRgevFBRJ+j++Af3e4NUVkw794NU7paHsJ2CuYF
WMYYxFYZ/rCACK1MrveMh5/HErRmhTHtvg6lkTRZo5/l1szEpr+QnA/mII2G
HEAUrVKUT1uCg0wC8km4/TFvyTHwPgNh9EZzPBUvWsj68pZaVDqiEuQoyfoF
ZK0bncthD97MqZlX5jQFchyFUoB2ybmJCw8jc6mzxb+iZQlCsXyYHddLIYpU
Mr3vR08+TaajyzttigSPnArdIBRhlDRmdjWOYsLYQH9lq90wz2ZN6OP7jGn3
LBASiw4W39TCpOnVY3xtVsXGNup8xPRE3ECQ8DsntRbuMPlY44Z57PbCzolV
LTW2aDrmZ87X5bKn5+kO1fLk+7WN/JWcTuFmaaP6gPk3vVQZG0JwMPNvbB1m
qReaOArcank43teV3Bc6D2nqknPtz/TSsHl16mjRzed1IF1JY47Wla+F9uWc
2Cjbwd+h8rM29Z5tvo4/BPklqjznJMVGVXWbLZkJhn9o/h7L2E1mI085qEtx
98gttfttiHNOH5tzOD5wtHaZEKRYTsQeiIziD6/z2OO8sEcbn3aLEdQOMvuy
Q5PaIidNvnndtHGP7CigI41fdXi9PU6Av+TjWN7C9CqFrMRxLk5nvOIGTgCO
Cg/iRw2VHHO4UwK/tGQ0Rhvg3i8O0ldlLZM6xY+N1efVp3ZSSnbt9yCFGiS+
6YqhXoITdQhyl3NEYoloMpKmCPkqa4fpwZGoTNQhiLxIh17HDMAyQSSCk2qK
tGq4q5CciLIInN25sFcaBn5cdpc4oXGA7yHm7+Qm5vUOFBy1v/wLAXCrovu1
rVdHKVgwn0tCcs8x1UGuUrQ1vWYgi4MLC/2nWGqWouayJBwoD1VI5rskwe5L
WM+yUmGRaUX9kO8RhaDP9tgAp4xxl7jIbcag8KRuwVH3yLIfis0Zk++x97LA
iQNoLiyqeBvx3JdDSDguTjjJUAoIcxwHzIwLj00gc/TC7mivdf6OWQtVrPiT
W4Mc8NgKIboD7sq/O67otzuaWaPtp12HWR2H1kc6wLS8Hn1BGVe3onRr0ixQ
h0e9nGIiMWyi5zl5dMv/NqdjEdalch83EmWE6QX+u7IaRN2IifJ9tmhAdBIO
1I2FC3+qKkd96wmwi9+98FYwL9PnFUuRdZdbeuCACM7cEMcpORtbv7xVbsfC
xt92vj24lm3YLXiCnBCyjGpMQi+5qDLBM27DT6XTi0o6UaLQdnev++S9emhZ
KW/8pftHeNbvbhEAGDAD6KSSNrRrL/zh78pob9X4UTxiTUwUbew53X1G8LV5
Ra7ex+OmYbIvCxyHEhCS97QYu3GJMYnZhfSUjZO1S8UYRwWPPVyyJnVHkkdX
QAvpYiJrCbbuYX05is+8yptOKjzWWE+dwyy055Lu0xtAanJ5BbHH10Qa/YdA
DxWPsNAL/5f7XUzDMOxlcya6sQH3jAv8d7esjRPbjIaQJyhfIIUEmD9aEyyZ
CA2Wz7pKr6TUJQGfept7In1wvOs5axWxPBdTZcZLXGQRiBlSsUQa5Jyb6deu
rPNR/s7GRDgkntG1/mHJiXxz8ha5FSrigfa8jaY/FgknASdtYLDMNuPG3Jcu
pwfMZRGj3nOZdx5B+YQE4gIirwpbxPNW3yvSGpO+oHyAbClF+cjDNK2aUXW5
Sb4eeEGUuLlmye8XGXKXo1igqnGmaTrzlK7R6OL7XTzMOTn8yJL9qPMwmAHi
n7qPalFg0OoOmyj7powp2e6cG4ZvJof58XYPv3T2Dgt/zDNA17iwRjFfKqXh
XUyp+ZaXQtI39LgYy4IXrMEJa3VNtlFn6BngxEU8PUeaepbuMV1R5POQnvYb
2BGwtdhZJLG+6sKifduQSxBBGZfb1O4uEF//zQQJBxYin+IUk5qujPPyLxnp
Swh/andQVGZSLrZxMstnIsmM1+x1B8Lnc4omutVQAGMP0iPAHd8DARcthcL9
A8SofTdL8UkmVGkHMQRal1wHlajeqsXbSRq/TOIGArh56N0kF/BKE4ChSVIm
51QlPQqkX7O9Ls+MjdeC8Xm8mre8CJIiH+z7pHOTA55BSeSQGEQawcRxJhOz
xk1uWTn7gYa199BTp8SIl7WlhK5cbXSY6KlPiLSlVNOPU7IiyGTiv3TFU1Tu
lPFX5oITTbWxm/UrxYrs4zF6W41YYaxcVAN4GTisG6Y/ln+fIeIARfeoCA6o
fPow7d7ZCITt58BLwBi+MdQSVBa1BFqmxDoNtPqbSEKn4dSiHZaiaT7sCKOE
SrF5clJFwG/yyIWtzdJZebniYPbfcf4hWvYV1620jRO9n8HGiANOaIQeTgNB
C9AhMscTUkgTCAypI0K8Euc5asxLblzl36ia68P5TzWSquvaExqgMjpPO+H+
ex9YBkXARm7WZBiSWN9WGvcmZ+5dpL+3u59gS/k6vaK5Po1f/IUumKZ/shNa
RWCCghZf/0GC9OkQCO86xa18aBO/qpy6zR25TQqmwKp2tFS0SXdj+TQNPX/6
0MksnlUAduLIOmma48CwHBotbxArdSDDySFvROh5usU61ZuQ24SP/szv9Ez2
E9QJ4vxk7puanVg/fnKx+s3KJ4MoJMoMfk5fbhrEAd8OIPx8sOdqyNSd3KAg
PtG4mNZg+r05AytK2aapjNE9dQQjQy3R6RjzxyC8Q+W8abRfPX/gNsAl+Z9V
mr4tvW4d+B2oov/Xw0M2cM/om6AlkVA+piedGILJ8uqR7YWzG7DJgjXj/Xnd
KKNGVFRzNe3P1LU2pLzXTHWPL2SP9nA2VkGMfD9DNOYb2bJaTTqmnuawcouT
57d0FKWNuBS8pzqDokwMi7iYHMHx7KKJA8chhHh7glrVTTThqrRAdLdw1415
eBzwCzQonXgMJWUY4wTAq69hOUMFKf/1LNY/kwsbYlQOvBbzt5aCaqvNU2GZ
vQefy6fChWHuSjOmN8seTM/ABt/ES6HMJZl+vny2C+xwRJjx4g1il3HfHuMK
gsU5p8RVWaGYn4LamW573dl3KPCgunCBrrNSPnA8k2ltdO6AjCHQoWnPtvaz
blJGFTKKD5dbTFbnUeqnfHa2DEF8nSYV0b1+Qbai0ka2QwJMM6RqY9uVNwl5
K7KjtNm/xPvrYVo8O6T0t0NHrUpWPDezTH2HXFVNquWs26g3RDzkirY09T5a
AN9cfQ7GJsSeJfY0m4b2IaiBhCLiJsDS0ZqEoJe37xDlVgDq6R02fs2zvor2
7bAItvYvQiBIbBkllZDkdso6nRMRwN4kNjy8WroNXOU5D97Ig28XDqRonQah
08A+1UgJZdXUGtBBzvRARG//2+4P6Ji3RB6Qnz7Qko9/jeNpdvy+t27HvLsO
xzzk3mqQzO2gYADmKMHOy8uUt5Ynp4Jana86VGGSmF7GMKEES2Lg8PyVb6hm
DtxSo380DfqV6hgvenGz/MnaPpMH+2+PTCmFTPurfHJDF2/p1upbssD+Mztt
mTj/7Ysh7mSae4uVJhew8bKo6zN00V8d6lSJmhGTX8H5LmtR0R9cam2jkBWs
+qPPLj1PWtSlS5kdUGBwt2u9CyTM0RY6F7Z6vRcvnWY7S8D0kUNlbik9Q4FV
Vl9p+yF8VAhpqYwQWJyQsccIFe9Rvm0gbb+FVVqrJAarMD8ZByrAAPAXh8Xw
HvOSlXPHAXjZlbXaSBW+OeHFW/bRTFRs0GufIQ/u9MsdiMWArLNJxAKcPJyY
XWtUtRUm6TgZUOGQ7cGk6LoSCaHbK6ng9lDlJROb55idrMsIzPusMq5Nij6h
o2Lo74yt12Lj7FMExoOnbAKJaLCSvCZ0h3/d6NBjmXoJMY+sOxbLCyH/7tyY
JigoTM3y0TAo6BNpGk3IIZstxHZWzXV8bl3zZ726Vy97KpEn8Hihg8fN1HXq
IfFv0CRPssnsFSCjSP2c+9ix2ddIXjTCVTDv5Qg9QWt46c3+DJlSOTq8nhdV
cZXZcmZtnRqwun0wSmt35Bdz14lPzEwstA9KP6MfJWG7/aVMLDeuOXxeVyfa
s2EvtTYfETu0DSACzdRX5I00Y+Wnc3qH2bemY81SUCXVkdLCVspeRF8WL02t
DJsBsvrQOEIcxdDoTfRbCWTS//PlupKuyUMadHICdlKS5zupsS7BdVZPU7hh
+nKt/OYXal5S1X22Ppt3JSJBnkAOEaP3BWEfERnbJJRrM5RYFWgHPu5LhvTJ
/aCPw0pLeasgSXpMAJo2Lw5btRrAfUMjzZzQIRnXbXflcq7OVoD7R4661aB0
qATtwA2yy8EtLb1/J9JC45F/AhuCDabgeokph79NYj2MLrHYiAkD7mC7oLgs
LwxRN5hzrGl9GSV6f8N3z+Izi+ACO0i3OJjQ9v/+Y+moGyitBZfDKGcfomwU
b6lHo0BnXeZkHDw9ely3rRiHt7V7M7rUqQhKiNnGXqfX+sDkKNd+5YyN++5b
wv/4F61NHongWAMZ5AsAketFlP/TIedf4QRmDL4qHLwReYuRr3U+mal52JHi
w0mcdA0LbOUP5jMGhFzTxyvcM6E88XS6G84X/XqVmx80zEa+lTkSf2mbCLWy
ZkiVo8jrqxZujyZNhRuufYToCvFrBxrMJij2EA/ViQdrVca/yWleC0ObOXz2
XT9Nz9AVyOEH4WGdoxEd0D5OVmuHsiMIZa0qm6BE/UwyMiSBBEzm2X+tgd/b
GfTPrDOCYMcFsyRh1KEI/uMc9DAzkpnrCTuPqM7Sf8TM0qalnjYwWjKksHzc
g9cITxAHpnT2RWxPpsTVWeObeOkzOx3oQ6JyvUF8eQnUDVjazAoRt37O9ivM
vsbyJo5Ox4l/sTu8p4W+UvSLWqTcjMmSxCKwAHEi2D2Vn6UnLvHZhKyoXiMp
esFRlX0NPmoR+b/xMjasZ/UL0Jytwf2J+pfUrRpnamBiGUyoUBn2HKNdlPWd
uCC5QrS4FzJo3rJop3hytyg6hjzed3FZSvYFdNqTx/7hFd0tvRm2U18VLsNM
Vx8LN+QkU1qdFnLhkc4dptxpqrtzNSkLaB1CzUKJAsPcMGl7lVKC32B5ys+f
oN7l6MyMHy1AZaPi3vHRImUSawcRPYL7dMmXyR3ZJbunTeBch3rs9XWP3ifR
kH73SBYJczNgwarfSgXIfIibRn7g7pEAkWQuZMq0Pi6r1ACX/7g5E04GmeKE
e7J+tlj/AZQAK0Kfe3K5S576VhGEy8f7HvG52HeJJgPCN8SLfFxSDjpChZJ5
+bh174F0xNJ4aGnJ6ePWVela/KTjtKW3so62m6LSnpsYqALoZyQb3QTup/Eh
Sw6mehmTyAgFE6IGMDTt25N2gDri7ruQaJivZGuI9bA0ehUJ1fU/bClvg7Pr
EneNd1QTDjhWKsDaSY08QUh/CyKQLq7tdwDa9BHHA/ReAV0e/Togwfo3wuy2
4MmmOQID0xzjmxuVZQDAx/kpvdi7oQR8rg+WvyjRusIkEaErKJpLIlL9OLi1
vwmh500GHJtRnlEdzPHQtyZchQXNUwP0ZiJKeVDa94jBn11TJZ4MnjAc57fA
aIK9QGhgCCZkx++y5q6hitIYRLiscirw6hvVoBZdWm7FkDWZUNOm2SkOHdek
oTbxv6M+o7xuhsCyiwmIam89NNst9pllx/MkLBRKnt35MXjzHTONcxpZV1g5
fizg2iYUJFVDfQqiIeL2GxX2KW0X8CiJuGzCS1O52TasSNhJ9IOWP9x/HU3W
NvfFnwA8sCcfSD4TVtQWxlgmp6TcWxAWVmzf6Z434Bp64p6D0gpz1gbe34yQ
+Cr9AIgCUovqrbyu5PfeSuN7YBet91cnmNMO8iR/Tyop0gPqdNrnVfnmjMml
xH/ZFzJuw1HUu8hUnqduWrE8xnu1Eicm6YUOFjQ25vDCgG9YA84345WetZAO
7MlT5g8XB/b9xc/t/2yvjgx944po5RIVtYfHKckBoWzqGvkD8clVjs2rwYDJ
hRC4Fe3ZXmwuq/ysKhMG5yuz0Y7T0fD3SVTGrmo1O+n3dhNuVn2TOC65r1v0
9UhX6Qv2Nq+U3pskwXEyyrI3rYGAv1hrN7H0iPuNnkMM0MzQtQvsX7XNl6fa
IhfDHrec0pcQfop+zx0v9aN5TsgzYfssthuxHV3s6JzHW02RbD5k+JQVAN9j
rVtIriULOaqybx/ZyNG3kjyw9ni1ApA/geut3v6rtqp4jO+AOMahqAJtwdgA
U8fNweJRDa/9VskRRbYxa/EMCcFo3HyljfIof6xjS0KmeeI7D/c5SbawMfD9
6i0HqaWao9tDZP/3Hs6VQOJ4FrTakm15jBe1k34sBwj2uebiIlQYqEJYWjv2
quD5u98kvl76IBtPuzLdu5Pn7dmAjf5FW6uaT60gx5qQw82t7IarTHP0/5xb
HVDqptuKIossC//QQafCF1KWfagRJ9vw5VkLLjwhmKY78yntEskCgowbO73i
FVVYYmjF3/Nm8k2MGakKxKyhqSasToH4jCGXawm60oiHEUBBQ03LDzYwH4bR
oNg+5IZiCIJPIdhqbiTUOPaBcms6i7L32cG+31L5n5LaxQ1GIDczlaFcpNRH
QgDRZxI2XwbCoQpVcmh77+wOIjE8cAhTGggjC98MTcgqKmtHiqRXOrrt8HMX
Pi8i2E3hysC6dS7Lwkfz5+3K8I0o7/nTLZvYPpDD2DA3rSP2hYVOFwmX+H30
Azffr71pJlDnN2wE14j8EYKSz8Lzc1+DPPb1OslsgtnMnO7gNiQx/jEPhLhE
bhT++NKg3EBHoAq+s9eYmySCVHa4JrgGoziG23wUr6CJXs0z8+3Dru/9vybZ
MPxsjoNQyBE318YLqk2dxDw38P+lcwFKVOD1yWe46pRU125Z7ZtYzmZ1cspE
DDQlwaNPC4jfI4JEyoOUg5ATmjJvotahRz8R0wwTPNMRZOR8rVvbsSd1w9Nr
mnThNUbE7F2sA3v5wE1l6d8I9102nHl/ujU6l9dhVsTyz+tNhA3n9D3NfpQ4
U5f+zHJAaffRJyvZHcn0C+rMocsHEe9mzPABV7XfiHB3yEH0SVGEIYWyBOwb
1volRrEVIsGdzGF3Gf1Cpr0KrzWxkw2WlCjsleHtydJtqW9K+EwQXc9kLJd0
IrdlZcA1EubfMBQsowHiP9COZ5X9OjFegauYiQTH/b/I6/DjmlYSWBboMEvM
LEPzSZkDooeC0m5YyG93uVMiCLHkb3GJLGiE8c6nod6NxV2JjtaqiueuYZhc
fQ6hhBve/3BBtrrov344+/+vn7BvOMTKUOZcqnIr5S1UZVU1ynXUouQzY6jL
OUcdX56TUkDyI0OpY8y5hZOpV7k2xx+GoynDXVe2W06KAZkMLy1aRmf8YYDP
8knedpVqTXc5mOAEUcL/544Qj4ApZAOnthjz8v44HFkca0idhUboLKKmFOB+
tNx27WwRlju5GqLTz7IlNxz64OQqgs4FlwAKgppTClOsXsMpLsmXzTh0CkT8
zdguDN0gWcJJVz4PAsdLS3PLbkNau42zQvpJYjc3IHcLmjs5/tXH8Ip6NE4i
08cuyulhlGV79YY6d6W14Z1AhPaO1IR65JM43rQs1NHY8taLZn729hNIqlDQ
TfFy8BT7ctqJhFy0AqC3ZD4bGnI5nOlZQh8r90pZ2nZoa4SmFDToj61wm21E
bxgXPBlBalBTZvETjE31MbSTT5Vz+hhFOjRC273FqVgTomP3SOcIMizEJtBd
k7LqNO+BK7nTcjiliVvSgyJ4aOeVQA75R3me2KqKxNewmGEWrmdiGPVt996u
uwoy1T78EjmZn6C0AKxiMSaV46armq0D9dKQhP50oP8Y9QcZEMS7YW8G+HSh
WfzYwMs8zIRzu83kbxv5xYunFW3wR0MYCEOxckqMn0LtmsbdZ2MwTd1lrM+d
He1bD2Hh55DWssnboP60cAGLSlBl/7enyZj1DxQGVkUY6LVvLs5odYs44fJ2
AYB5KS55kNkoVOrgCQ0wa+g6+doigTpdpZSrjZSA7+ZSnAbbiGpCriVpVSjz
fguSXohTzBrfoas61uvSP9fRj6hJs8EyLdEqlgha4HRCpKwGA+v1S8/8FH1X
x7GlP1WD2x8HWalzofOrRdW7DYznwjRRE0NzNkNaE1HjIFRBeXw9AkuRhqim
zkYDRvuvAEpRMlkQiD1OGPGdA7qfKfkC0WgaSx9lbZt9GlgXVequmJ/Izth+
zyuibAIIgTHYYj5lI7z4lL21Um2lPwfCBeS+4Ii6GOSRF1lQSYSItHnRr5kR
ZwV0joRmkON7HSYBWz7RkUQYmoFIUpeXktqBStBo/6aCUFYsr9nzRhCe+eZ3
thyyZ5142bH6krvIlvhkfpdEPK8GHCez4tQvc0dBCTOUpykTqYh1SuhPwwtF
PJrg9q3GQd1RWKHuJhaBb/+zsnxm6dcOaxPoePPvgCyYnjrLnzM5NszOeMoh
aTgFUjG/bGNa69CVKtRTDzCNZnaAd3HCj8hXxbc/Dl1+DrUX3ZBOBEXI763D
weA4exmSJdTkCWGMwydI1ulkvo9HSvk+P+DaLp9PGBEaRIYGsc9ZXNX3JYFQ
dJszDnf+Wm5xm3gad+rGZeSBb0qzknH7qGIJ7rUj+ilnHNjidxT0cg7bXb6K
gJlAcUK4FTNnecURhwzTa1IZpsll576Vdpa9cpm3/CgZdioVphc9+vDioQjg
lJHMNBu/A0cAeQwkGHnVL1DiHfatN7FNjnZgpSq8Gpk2PR5iE2hVuZWi7TU0
/Uqse8A0A4h5NhVBdz+w5f/qNA4bifFPPjjmSSAeECM+1Iz2HrMyf6K+AZ3T
VIwjMDkMG6zKhq8ZuMr6zyk2LTw8b86t4g9Ye1a/6pLNxdVSmSTLC5PiQ4HZ
1IKG5RhVtPoIuM4dK1Utl5aVUPnaJC8C8f6g3XTsACcDQXaa+F+N8TogNhaH
YZ9y4GHjuU5lPFj1UTGzCtz99GtnKgX2gNKKB4XjrpB4A4p4Q4BFEVMJraUj
HE9+paVjmrcsGXD64HlM2TR6WwX/scWNyLLo2/T9nMpU9vFt9xbMN86F3COD
36lcGLhOGO5pUmHNiLNVWxZBT1EzStI7tN1di0K/iCQdZU7iQavID8OufeRU
LJTDlbOnf+nG8pUwuPyck/ThZsMFOf9TRatTgwf4+0TmeSh7ENCIPrq6XBQ2
vmAeRKAk5gT8c5Vy7WxY+IXcIcApmwRoriPyylQbd7slqDs7PIijxgTidhtd
XaDT3UbG3S+mHUiCa/ajHFvcgxgh9hQcEJSbO6G7GvGNqFCJgHWREfVLc/io
xHDP4Euqo0/XdttaDfdknid26wtDNxXeO9p6Lu1eJju8KhKlirp79pP884jb
On6V2fd/ubsBdgARcE0MDhOoLHzF55SDs89pIgpr8vLQH8GciaLwLjRrAcNs
4OKC3Fhc1fcLfw33EAiVWUKVAsRgULSpm5QPf3SwG/MQceBT9qsYw+AVwKFt
W3cUcapkPdvKouUoBv+hevIeQ9D8Sx54iZHvbKj2yW8i9Bn3pg0dUsOgz8os
IVv+6kqI4466pyZDPJyGEUCwOMTODw42X9q/eSYLmZXAbvPv9gVEj+tl7Rd5
zoXIeL3om7NE/cjc4BPfNKTS5/RyC0+T5kXEc0cLlyv3bZRy9V7x1D9RJdsM
SjpwPhsVkq4EzxVKfZF5+j7+8bjKa3CX1PYpLcsPYHtThixKhU5/arTAj5eA
sF4dhTRhoUoHyouY+duIiaPel4bbZqy0lBuSW8eyoL++q3JiiPNF+gkwoq4p
gn961vBI+EUziC53kKmyy9aGYhBDMTynCJlozsvFnFp14Lfb8VfDeRYBkRAf
DbI6Gvuz4qYsFqrBxgErbL82h9dUCjdX+zB/iCFVFUvJULbFrdm6qEGkkVpv
f/MtMfEU4PRXVOWFjfhYiU3LfkFxB69jN3Wqujk5JQgX4pGYJKoyTGSerYpg
SMZt/XQxl+PaoAegktf7/MlSK48EF4OjbikE41xiY/MQwiJ2anKljfqEI/vX
PKtT2zzV3YihGknD2blfVWK6CtpFQ1wzckOYtsmc4ZjP2LvWJji3acnt7+oa
W+LLIWqN+1nViOTVrmBEmHEDSweoxb9JOssPP+eNEub0w/ZoddnhFiERuOfV
IEfZf7Ydtj+Muc2jVq/Ck1VU18R0prhJoay88uMxyf5c0p5egWu32AyvXTKB
3kuoOvkjYySRp4mvX4XBpHlsfbpHX8v0YThQ3iDT59M90dBj3oPPj/Jf74J5
+Ni/mvouUeFZXCdEeSs9IEAwDlvXgUZDy/tlsPoPeEmXy7FNux4IUpqleeWX
iNIYBBKwajL//YcFxT249zNhEetPfDMmEGfLJi7Euwgr7zuJMeOGEaC+Q1fV
g1DDVxP34ecNgG4CCIlf+QhVByo2S7+Zyiu/SPC+SiYrFbZbUObI6TCyGAUs
RZqReqKIYKOs6Kz26veCillGKzx4YdOpjjNRpRv6ez/BmZwUbRBmSyFWoqs8
okc4VYDq516Ahk8L+uigfUy1uweAv8+MSY7i4QHT3a2hg0vofnJ6reRsnHjT
8qMJPkO6lNfD1Vy4+jHmlwdIDXjWjYx0BU6u6N3mvgNoBk3SBrSpc8xvCJMq
r3aNlLexcYABltyt/62G0f1l5NOA1hGVeL5us36bcS3FXsF5ZsUXVixLGWtb
EJN69vrt3LU/rnWMVhbMJPFgFG9yYl18oLwT9h2qDn4/irY9P7wLfqnq7hv7
7m/IpUN61v3li+bkEwDdfMQtr9lFrkE3k9cXiLqanituO0NpAES/cBuWdeJ4
eq/XiNK++wdi6ewhA7WDvWGzNFB2sO7Dwe2/UBn8NNfUb7i6JOCnCVKlgCN7
Vy0tFFGrTL35q7IEuR1lNvYl4LQ5SMyHOteE82yhqFFNRCGEkvXTDg4EMz7k
XEDVjfxTmY5+6t7y38XnMMTuxp3kqChnQxeq3muVNZxMC0hOSOLuyayUSAVR
U3PQ5pXocSqegmcVt/Xyoxo7d0d9Y//fELaPraWQJ8QuTOszSzxeEl6dQXs+
QNo9BL4EnB0TnyLzFv6X9nU0YNbcf7x7gUA6k1VuSZ//eEPALXeNIa4TwUJ1
A3auyKDYX8KjbsHvAW1Qm8zrHc3D4vBpB7CkF2tisozyGrXrlzEY7GKDIOH/
dK7fKXznT6xVxE0owsXrYpYJhE/TewhcCbH+dC/cxWE0suxHLZWiDcu0ZTbX
8yeDIdJPXiVnxSbJnfZJMWl2ht8zPS85WrySsvzYq6B/Q5fUf/02PY05uZae
UERYpSynEH6b4l/Lg+e17Nsuzu6w56QV+dsvqdv3XlwH9z/zBh0gNNSA3TTl
Tx93y5GFaDcEeCUS6D99hAiBTGEeTZtlRqIuOyiFwFTolMRGJ5gJTeWIuOII
JRkS6RX8MQIpkoAjyNQdF9cDHLCldenoy4aHZgrioLoYaFVbmygzA2+5/pMK
VM/XcXlnW8x+DyTpDBrv23+OJ6RmWn/ZVhNC6DCLcni1VcsnUYQmk0+3gs24
41Bjy9jA8w8YitOzurvppGprTvIq8iL4NF8dCCDxG+Hm7RNKrrS33oitBgXq
0OsEseWr0bV+10qO+obU1qLu7HRmscX0ez2GbiSqwrYOMPmfb912JyfqwHBV
C53XLL8tEvPWulkxSZzS6lZuBowfoy60A1avHADy1OlMlngYeVK4PzH/91Ok
8R+eCQ9frFO40frUrAMomVxyeAbwJV7auhm71DDeQmnjLXqVSbW3vgv26MRn
4u/eLH/TycAIIQrAcxPU0AFO66EWqivcqqQlejqnS86bHxw+m6+xDPuFxVZz
JtNELs/YRjDSwzIw2jx3Vndd683FKI9mQyIJIiaa4+12WnAKIASJJdxwm5ru
6Mths5kG5kaAovMojXzAg6tXT/32K7Szx4Wq8VM54We0VXL5GJArE8wvbaeL
lHEFVwvMLygFMgpCUAqgzYaSKYTaPfa1EEqX2zHNLkzg8CPg44pT9ccRAMBf
3hsb5jwD69ltDbEoZ5iJ0zHICpNuXmrSCuXgxVDrHL8JbOt+1s7ZLjS5HnBO
8Ly+TVZs+dJbmIGpLcwZTTGTFG8TTi0v2UQ6zJekvWt6po1WOdSabba6t+h6
OYAcWNe7bsbtV2CF5JN4MjBZnsV92DGtXMP2KPZkRCGMtJXEYdF0jn3xRSHJ
9xLregQV1lYqyyf6n4dDvIHFokUZ2INPYuKV6Tk6XyWrXxdFewR0RKTsKtda
NLaWaspDmTySnlTtWPXn2WaMDmszVtVVwjQvpxUOFV3LZSjf4OiANkQkpqNw
Qn/f0ANljoC6PMl/KnijJmXMOEX7luMUajAzbVs2O8AfpUoCz6gQOfHTy3kX
+0w4IUXup2VbrA3/t/i1grN975WJQ//O8YJssTKd/OtZEMBdbpIFvQL3CPs2
Ism/6eIoz2YBGrrScg8T7nIb+aNfFkT9pux7H2qDgowmUrzGSCvL0OBZfVq8
og8xHZ0/Qnn/RaBBmuxyJSQYgEBiHi1V6G2NankPy+PmeLkv4BluOny4L6Ku
7MpzBozrck5T2+mlTcAoQa+nFIOHgDX7OGShACn4DtCPVmViXjpS99LnIgnW
V6KvHR4D6mnHkBGnL/racqu6LefNMzj+Lk5qKkiTM9J6jmNtRdwah9mEW5JL
UJDm0VWBOYBWv/j6g+LQ++4Sbc7d/Mc4qe6LC2ujPplTG7hgoaxpiay5VnEq
+nAKKNXMPJ/mr7HBFDUa3Wz8PtM0wDbhk+wy9GmAeIjx+dEr76K9ykXCVpl9
u7Yot8MPW6imNVn4zm8oAxUES4RYkIbqK9U2WjHK6BN8NU46dV+ltCV9Kd68
ohQQgAfDpMgCMiMr1H7L0FIpoUsrFknR9exj1rBiP/nHprf3LqxOpoPKjMNL
d1hTazHHU2UNsW82S7UINjSgsrQ9EAVEOUGk9i541zA1CKteDYruHlLDaJmH
4wekSmP2Zwxo/4QoX3yg0oSCP6z6UMbKgDbjGUYHsLJxYVsYhmykwHULabLw
uEBq44PnMC7lbwbVRMQK9PMqQByO+EG7SEitrVvon9/t7OKLY0j4UJ6pdo2J
Zf3RuXJQgUM4Kv1+0nNUoR3wtp3tlgOGhsBgG84F/16ZzfhqdiFpFP+aoQ/S
pp1p3Xbvr76K9djAW4VPejyWU98nqgGIJjS7l1B6BMGXEYNiWK3dxk73M+RG
lqe7pJdUd7ik3729QzLM1OqRHTY7purwTFRQWVL2X9XVN0GEsIOUdvKJwFFm
AF8srAruhCCDEfn647F0G+PHGE2bzSIeUqUKymqC56Jn7sNu6IqnPQaJ3sBg
Jb7wVsLp6GpzCuP2+RIPiLiyAAsiPcjc3p85v3jTTWLTmzbkmabWb+lgl7OG
xKFtsRwjLZeJDQYjaAAOEKqyT01VcXQIeIMbJxwYcQYPR3CWdBwiLtsyaBKD
EDFa4afBw6rHOMxEe7h5POVLjRCCAt8/QlNEYYz4NGLX4w9Cp+Z35uuM3R8p
/jiwD/CroTik3yX5AQiguyHhlLfFAQeXqA+2ms6o+EqEN7B3koDpfqbiG0zG
jkqlPEJSIauECvJuEiWRIxROQ1wZam37uSjW3TWa3pMv6FMQ6VIz3Z9xV/Xc
mwYZEs4ydTNZ4MCHYrOM5NY/52BDerldWGUFNti5SOMXfZIUPqkZtVzKLH7U
kBHKRRvnofYhWUn7I1acQc66qonYz+8ne48JSHTGepYTDXbE8grD6Y7rESJf
cEbnUqbVLlNS3lY62o0vRcrzhcXErjwIovH/bRa1Mjl8iIOFAAzzXkzvuj4o
ubbN796tu9whCTUegAxHLl5mzGxmDNqH2lH/utaeKDtS9rdRpWq+WDHbenYV
Z8BJkXVVR0+g3NQ3cUbPOVfqQS/eiWaSGY3cZZ2JAUd/GdGBh0tESBrf8nLP
4oXhcVbHXHDVt/itq9+uXjLeF2BpShCLAGfaszoWOf19r9PtHsDQ6HdvdcI4
yZXdJUK6oI7GE9j/2IMKtiFcxkES+b5EJn6+uwZWxsB8c53GZc5hqxwJbODH
hXGSE+5ipg9Ea8rWjKK7JZRgf2nhsPI87aijYJUNResrbQtJqw0urGmtSW7g
rfVg+DxpMi1K6ia/NNMLHqLN8hVWS70vSNqqfpkgN2c3FPLOuLbKsQoNpfyY
UCLSagm85e+0ptvZ//+ScpjcqBRUrVLrQUcDVRugOulkuKFjD+TLxIiz+32O
au4AGFvjozr+hh05eNULZZX+mbVcwiH/l5nbDpzMKox7PG9BYj9Ncn+ml6bM
5nwzMSZX9AZ3lXQ7oMNarRl53q5T3lCWljeuL1Z8hvC5dNmdXjVyOh27Vtyf
X5TI0ZE2cbRWrEi0qNxll8cQ0ekVyS0gxG4SdBeULBRGe9FdBHF3Z6D149Zh
HzHEHENmmHaHe5ZIdUqT8ZxtDeki7tJxwNb5+zMYtC132+kvN7pY5A6+/Vo8
tgMiqO4f+2kdZDHrMbqfwvBqUiQNonQVbWkXXTcOFQIj9KpFP1/fV0hsdK3h
T55uYuXDLCv6KTiJGQj1v7IjqiRfBCFQaulEhkxnu4LGMW7PmaFn3kyemO3g
njHHE+ma6Nww5zLvdbNfn4TJ+maaTaqOC5g0/P1FuyYGMy0fDs7fbcOBVIBa
0MWlfKQSNCMgDhhWFBpFp7zCVor4xL4RcJLFvJNJzUFCoGsADx8yS/z+9J68
ThHL7Jc1PlZkIfcLw3Rxf5zmpWstRrxTx+pD1Z1UcXAoD70kD65br5H9htxS
xa7vyXwg8McdceHaEWgBz6J8xAfj/zm7PXr1hQmX/mhmPEbv4+jti+Qwn36k
WaAdJStY0ge/YcL0iX7iBactkzqd7zwwTJEAN/tUoeFWQEbWGPKFM7l2nlE8
Kzio8LfTlmSbk7OrsydPpQ835O9ntoFAnAi96fC5ngz53oxX/36EJyzJ2E7P
2di72ZLK5Yf3iehJqHQxrpaxhNiq+ZgA/xSTRxMf3tA73EC41jQTolS0uFIh
A9n9w+Lydx7uigd/MoEVfx8T5V56q+lDgTZjXwtXohepdIreE0q2gf5Oop3H
FjwE37s1BC6F4sfy+dUSPBzCz0XxphmcIxDjDFQJF3qwuaPP0xYpPCwoiJhQ
L9QKEpCtqtJr/jhW2Pyxf2S9UHQXN8qg/p4OSLw/QWvx3C0VJxMrQUYfkWcv
1Ux3weuL2Zy8LxP48nbeD8uNGxYlBD/yikawoQJgXl9EVoNCgI38XE4tl2lB
ozBXoXjpBhCTU99h9l7pt4fQxXaFZwbFa8sipKuyb0EJLdE6/gDPc3nsYHEc
EBGCnFZWHL3DlNW0aT5uC+rvO9BtZbzXjzM5IICfe5WlHRpQha1LFS0FwnKX
0zUzCxc/P6VnXjDLYxKuoo2Ap/dj44VMhaLwGlgZ7SROViu8yDuedw6ymHeQ
hFEuMUxSqlo4MBGmaj8MlEGB9GE+yjIgcnn6ak9xiuQGde330VYjW1fY5ee5
mHxTDgdPjVZu4ibo/ROpQeaWKC/NHWTA3QxAXrnftUSQW90t/LxTMLveK4JX
X5rZF5SXA00XqcM3YXnE2Omwy+cCP9MJ3wiS+3H5yXozFCW8b7jVpmed2UQ6
XDpzNJ9EeIFzz5PxhsVUzVxhOvMkJMGkVEFZxZcQGi0xX0LMBy8bc1s471ai
Xs5W3v2OhzYiQP2HgDqTuLfExm6GD6bubTbkDo5PCOiTUUFSkoOZKTwYj7un
NiOdiUVg+rAD6KrTl5N2wdUDBoeIUTO5clfVnokmOHCATsJ8U0gyKvVWBqAe
3b9XN6+4NIjpY6nXivpKiEhPSGo5nuwkptqL+tdhtMCy2TWBXNSKZF8/cmxv
OGah1VkMPLFqAfxdAflTUi1s1wH0aETJvBZIK4yWngqCCkRtLrBn2szqxfyO
+KO5vhersdlbHfPjEngKwhxU14AZY9RLeq7mmkXt9On1POfFgR/i835RQiA+
Yp8oh+97QE6rkgc9mfYMszHDNan9o9WeWCsrL9BRb/SK7j3F19tMbTuh382+
dwQvRCQmVql25yFOqICturw4ADhEF6G+Qp9LlC1KQ6OQyIOXYAgElUn+51V0
qGdsHIrDzwVx6VVEfptUPczZFH/hjo1ZjaOghyX53WHHMTRh6iX7t2/EPx0U
cOCGP+lxRWCI+ZlD0kpPelkkq9HHcFLOS1NxbctKOHWX9K3Hx+jjYHiZw3bT
gyn0YDANGHL2fSRKUqAXoJASf8oggQ7wrrD+NuVEo9n9mDVQnSwMVC50qWXW
KOS+5HlrChCuIgTUstEYlYhNuRnS2/STRlRrfB9Q5T8l+U3ocqGIWdy83DFK
ccD6yeRG9FdsGl1PXmbG9FUWYxcPfvTxWud3yfoEPmb6M/vcgTeiC51T9/Ig
wtkX4ic7RA16mo5lVGZJK1Xn/wJiw7m8GTYy27aSApWPk+WnCOnwjNFCq7g+
H66JigWAv2/612UD4FD2Z+DWLlU6PxyRkxNd2Vpmke+cGOilOoQuAsc7X/Es
FGmIYweo53uW6rEFF2XHlrDWaSxOxgs+lmG60hrjesJwM7/U71MpWJu8ppm2
iS7ysODbrptmonUVJYCB0/oq4d7kKn9f3tUlM93HsX6sUxOpI1DHTzrFLjTZ
ySJ1G+YyYVLW2TZ+VQI6/vTLh0CDGEdyP/aeEudZtokpoPJlFAsYyR5nqLHV
GuGE3rZS58LmPv02VYucBIlJFEY4gbbNyWm6eseAKQFSpBTaeBWpMJXkSSDI
O5CDXo/vjdqst0kp4kSATUsCpex+4rEsG3jwFTMaszWv8cDbrJ/UGd6TmRYV
Zu4ws2WXmZO9vZSxv1Ro6suPg+Lvr5Hlj5S7TsIokYNLUdKYLMyHo3x3uOwG
q4Tes4iWC1Noy/gbmLc1MV9l2yNS0jOKhbu6dQnf4udTJHtbrNtYYZFrWidG
KF1B9K3aDmDagBJmAp+GalAF8oxRz9C7PrbiQ9ANLAMf6KUvpnSxV0LVD91G
WaOQWVhklTABZBk/D9rEbPh1IEn04vieSFp8xi1SLcCkcJmKhYmn7a/Wn9ab
BjtdMwx3pKD4Vp7/JgE3NRBjd0X+F3AOFk7azpydXen3Pqey2HevdljdBrvU
9zJ05BbNrtEyyaKyDVvn7fdvvnUryqSpdAWf4s/OTw/aCYnMckrwLw0B412+
JZIlnV34nOL7ATi0Ka1FxSxIYX/564UDDS6KXQFl9cf7va63KHfGwwFv4lJf
LKSXEkEzbS7YXlLdyL5yetAPzUYHU51LEtTq390Nt5YjToV6/80apGHkazjk
B8tBXhgZ+s2jgRDTYzRdLZBowmmLyBwxrAQw9A9HORz5TkGKuXgvYgfksnpP
XKwaKHBpihLGBQIiv3i+Q8cuWaVIYzrdtcbogc8ZZuBP228x4iwcEkFEvF1A
mNL+t6TGYTdLIPy44MgGICj5IOdkXFE4Lo7R5qh53oXkmzY3orTzDUt3ESMx
W25MEWVjhmNsGBlKWHVS2obR+q+fflw5VsbtjD/6FGeatzd+aRy1eS0wUSJL
VlTaOwckEq14hNV8zhcsaFXbBf1TEklfb7DG8KccbXzx6oywkjizxAE5UNdm
4J5qyy/P8x3QpFHXxZ4lMDZW5NhIOaTtiedGXWMyKNH+gCohWq3WmSvPJGQU
fhJYdZgx7qCjLo+YhPK3hfzLn2DkE8InNvnPDZM2usv3zCzetkoqIFBOC1Ul
nB/H4XVGqb7GBQcN5q33mk9IOaU+s7mOyZUD9Z9HSA7AjGGvcFcqICWS6FyO
ROlege/BPgnMtEW3+MAeXUlBncD63PPauHvNofJmxYCooV9463TC3baLR1lp
1oV0TiWSQzXXEycoq+H8ATV789SCdDxnQ+jhNZjPdTLqAdVAZspH8UFEe/0i
o/bYrYX3Jnjf//HkBsZwDhq/9bvhbPUB5BrgpglEs238mLJV3zYDB4sLlWe4
poGdKAnz45mCBB8H4sVkBRfDBme4eSIHbv+DSReDJGaiKtG7jGLwkYLr192v
kwuVD9r7f+O0ylqJbjR3qe8aRViAvJ4b0QOx7CcqGh5lJHCD/dmBtFHf5HPk
1lcP4vYsYjywLzePkAgXlLsaDx7B0sz2sExSZHwge2C856NZ7vyPRaDXWzBu
DOaa6fYelX03qOf5GFPrXnr9QtU71rtdvheCAQJqgPvbrj/tRU0UcqTsPvhl
A4gmEChIZqy0cjb+v/GluwUPCgyPUAWWn8o5XDGV68zTbNZmwTpIBNkKN2md
rAoNxiNM+dPTnKMQTwNZW6Fmt0OopxfrFi0qsTsBKuviJAWv+7I7pTjUs004
MCqjk/BRuiSJMerqAoRavjNwd9k7VyNP57gVH8G1feXCpNuuqjhUuGZxQymc
fwFkFlmt415eS7x0HmfBJ9uoyjSfOzNGPspvfIwij33bexa7Ngyf1yOzL3NV
RfTQhgeQhAAeKCKCR4rL8f/jR5Audh1hOf3gd5+rI40eMXN/QTlc4PeTYqgo
Ab9n+MRiypkSizpiA5uPpJ8S5FMqCeCaTQZhbg8dxfC8rdxWTmbPJ5PhoBLF
STI/sJnAHm0A7RsVqyy6oTvRRAb7g9DZxATk6iYJtO2gKpr08XCjAiiyA4Og
NzCe7VRdOB1D5fmXj6v7sr8lTMqm5lLrOkMLRx4MN0URsVRd2+LcndHZXSD2
17k3xxl3m/xsqZ+e6BI2HhIVALmQdhso3DlL7xX5bYeKIFA4fVijQ/NKMye/
+/X1QeuP2ddpdgg+q7E6iwroroRYCsX4pxmcN7qnsMQoC4yqBSGq95eSm7Mo
YmM4PthjBrIMNwCIuHjj8s+CVQNGVEUhFXHswacDvGnRip3dQpFZQ/WJHgNi
4FlHTD8EJkhv8001/rMBRgcBYiuJjXJe1MDC8vdXkwVAVOIwLRTdPSqH/KvY
wKgUWYV3H29Vk3vzxsdjp/j7VL9JY1UzA09fFXkqiPbGWRn6b5Ac3Yu9tOFm
8emJi4SVpAVvxWM+HllSRSTEoDGw9hC4EgWqJiGDYROmwJ2i4+HVhI3c6RoO
Ci6tM9IgroCduTz9E2uGbALrHC0t0d3YgUHP7jUTeEl6vlJYzZ2kOznL3qLa
sKlm9i7S4sVTDg5KugoGoZJmzOBh6u0HaQWNORX8gsU7/5voXXwVpNmjh9L2
OVzu4tNmib3rUsbzHKN5otnCHLFTUeUv+yFzWiRztpaU0Xdhm2tSH5tI3z9v
4wuEqYj5zfEEhYSYM/Js2hoTr3MTwtd45qVXAl1b3Y/C+Jnz4jjAX4lKnNSO
q8Uv1nfKRDnzxX2ywykMWkghQZ/yNCLWn3+sGQR5meWXvBMzIOrNyNbEeIsz
q76bl+4PSllkI6J6BGe/O3oZY1gPWKQWTRHVGN4DTq6uLNJ8WzuE4l7hkdWP
BnyzmUHGkA0zd6bnVIyijDMXQtpeeJzcHvFU5V+1PrDZlP31iBqLimCaSX3P
9mwuq/HukriHiLNIDR2w5uwXEsF8qeuwDU/JTmKW3tDEnMrKn67ffhNGAVOX
qRlCaN1eCfv3WYTgRYBQ44mM51w3CmpkiB/D+MDWcYdslQcY7ZHmdzBnUWOJ
5RxyWTkpqZ+//sdtpk6xQmSSyTHuriO5F27EbWMcFMYM+ZlkC0xKX1Pfv87y
ilYo09sGs4XpQcaKS4wB9f+DLfu24eXzNb6O1PW62Jswcm4WxhWtuUgacqcY
/N31SPA+TpM6QD3mKdPaUxNZLYyQy6pL0zw/OcED5UaGZOcmHHx7MI/kiSDb
aCvGLVtwsoefTO/lWu5f0kjXElZRwjqbR/iI+ZbpBQryCTdK6vayuGkmSIVx
F2Q4aRIExrDXEDKMF2ovEwZWnrdmECK3bi42hIYLYLfbR68hBUTIlXTQDWSD
zEqN/3F8huedMG4QFRe/3tJCKLIAklZGINa44vkuy7GENTDRiie2sIUtD3QH
IjouaLIScPoopqN4YBtwRiETS1PhijqFLvS1jBSpmBGsq1BCBO84BA5znABG
g3RoUytveKfHculwRDZIee28Q3f7ypToSrxjc5AEWxFmjkgFHo8lMLpNrHCV
YgzaQZX0jnY+elj7Kk8CTPwlRiTn9OoP5OdAD1khF9aEgnwXlokBnc2BA9FT
7uZrWr3Ctu7yzNeiNU5pHrv6D5rvcOXDQvY+qHKnOrtJL9iCXOLHqRm11M/4
2DnaPi9hQNIXiKOwKSROoir7RL3fFcY1miF6wfNXhbalb3MiR6HL5/jyquXt
vylvJVMJ3oZ5yvyksJVVwuQxItoGSlSW9WAghr5dnDXj5+byphJaMs3y5yxp
M3E54otyyVQXsCk3oZGzF0owtOCD6mAPQ+Ch538iRRnfRlvTQULR4c2911cj
shcYn9d3E+3QPW63rYl5EvSkS3LKKHamUX/bEmh42hoFeLJ3HrsNuXjRuJiv
yONr3oZo9e9w7qQI5nfSxm1QQE1Oxh4u/XcSxBOjsnvh5Ilgvm6xGqT2nU0H
Ez+BNqfftRkHDTw0fRw+wxXrow1fpFQXsqUM32UPcJ4Z7EeieORQfk6nLaRT
okDSLalAGT+uySrS0NCAxzjIHo6q1i9u/ta32zJzoTIcDN3bt5W3vY3gGOsI
3o31oYBrGL+960hmgbs6N2cgNOY7Z6WE1iZROvPXPt104dtJCm5rcnyZSNBp
xaFAF2aG7ewx/a+xqhdb5+/uSPDKJ/IrHGUvcr63nnHQWiK10nIfvAuOQMrf
zVhb7Z7+OusFOYteMAqc05mXmMDctnLDfeSrH61J0fh06DhQq5jvLWqZ3828
M4JYkOIJAx4FmTWpLEh608+Zga5lTxXXoWhLYehqFExe6JQ5ZrmLA7pDOV3g
6KJi/LxkqfdYKg9HQisP2/IiIl+tQ29ysJOfNRVpBWall3W5orHg1CRXrDjQ
AE1SZsdox/3RzhHx67HMMWtH6GLnS0FPqLRXIvMHS93Nt1Gx/v7YbUX/0l+S
yFWZifExJhwADSgRzKs96hoAqvR9XpDITGW5s2L9Kr1NMJ3XnD6J23IAJ9Eu
7I/kYw9x+L/N8UFyCFCg0oFrFdqbU6oyMlOsMvXyEesxEDpvJILXWP6mkfAB
K0bq4dDbxNmI3c9igpUvFQzUhqWAmDhvzJvpJFdwaOQn/oBj0buH6oYV4JXP
WcPjK1Odd9aaEzYhpJqBksXvBpl5T+d6vDBb6wmGJGM0nDDzOmV2S6tbAaN/
L95pJ0ACVYU7LqigGMQ0MYq2+8US4nQSKLApoT1uVHZD7DRUpbRfgV9v2Ul6
7wEf/7zzy5oT6I7ORxzJgJK3pGvQ6bZs49IU8qZtA7nZdZrVn4elSKNyD/oM
7ozFjQSHF2GIjFMUGDJmj07vPAth43km5OvvuLLh6J6WNneNmHBl1lQTpXCD
V2fewaaIv5ifE7g1ex0YVFKQUUFtKd6AXE/PY4z6ovQdHqaV0Yumwvs9bW4V
RclKno2Hz16UsC+2V/Fs+LnisTlr/t5yOiPOITwLgKBuuDaQpAsL70mFwkjl
FXZjLF++KoQ2QBMznhJcWeDdl86mJduw+IIROK6rbItdSqnvOX/wT+ecdFHM
Zmea2sL4/wx925GS6U7wVqaLHjYV6KYruYK8jUWppCVaS4VKkflqfDfIf+N7
qDZJe02ryUBq7NDCwS5dr7SXu31ttELRpjoajJRwOsq/ZHDFyHc6SclQhge2
AM1DTi9TSjVdvCVeMFw/P1cGtW9/GFjvQ1tHIINR6D4TXr4KeMsvjA5+8B8j
LSMdrtTGlyT2bhRMfyUYLBJBjohNd5Z0zbah01YXZiLDkhWJ3bZ9YNCZC97a
hIF0DcE3WCIM/Fec/8vbUlMZAACyMqpl0BSR2dEoJKJcUQfRq3X+poV279P7
UpdxCgyuNV7t1WSzrDXnhKV0LBUU9oc08q8oI7uCi+He4RWL+m2ojlFnogLu
cyoBdtqMl5UI+app7j/JS3QBU+qdDFaGilDLR7D7vlJabpsY/awTxbDX61L3
6OrfhQpUWBA4FbyYO1QC2dnKTfiP2cQF3nyTJGet0ZcvyopkXv6rc5m0hzUE
p3gv5F6INfXgbACc4O1YXLbeBLdoSo5CIdO12eO1C+MrksNcSVEZhkPhzo9w
R/vEpupqdkooe1lFsDnggHmcy/bqDFyCO/1Y3aGUusMkf7xzsg0wOibhr+zj
RHTff3kJPS+NL9C1gigfUxrPUyeZijQWiRDKdydXB5eGyuB1PSs+wmSoJcwM
UfgAMosTQutn4qpqmXvuWQ/rryyNlYN5+elmGS9o1YGsoxUpGp8HLqw6z8WZ
+6BAcAVllKv6FiF8ZRp2TpWYafnfWBY11fLZtjaIye1kDQvJ/13tQdG60AwU
XLTOQ0eMHbsevqkz1IDYdqDGI+P7rXeYoYDrdFHBMjxCp0Lb8cnRSJrjWsPz
lYOIwSXLc4GRRgpsXJlSHc6M6gmEjDvJkzpcLefChqmHo0jMLL1jLzuJtJZ4
48ih5ScaSzXJvcd1qt8q54BXqMDYWe0vjiHtLL5FbewHFuKbPAoxFo3qnwEQ
WZb4EtyDvfV42xoXNdj25yknQ0xAOBfk/9b7WqVEH8CEArwi8d3XaZMZGmW1
JGvEsafuvM8Mzk30hEnm2VJu6OJs2H0qoZJexYmwhfIuFZvCwSmZoz/Yrtby
ZmGGuVdjqio/7CxlyXpjAYyG+qhncQRLFEf2Zu7FsaQaWPsHPj4H+Yn0mUgs
LJhMAe2/WWqwqXJYFO8LKi/RX5ZWma6kbeViQsdBiATlofbty5nCF8bM7wvP
HSZA3DBep9h9qaOMMvM8ILaV+7ybyeRmL/PdplTEeTR/p08+YTdvW15cOvk1
apK39T+qUTo83hdzQRQ0hzo9U5WdTEWlM66VqeV40MH03odsIlrN6CBJZ8Rj
3rSXDFlJtS2YNjdGoOZSSgD6dKMr30NKWokwtGefMz2USKPrBfNX/2Ca3JPu
iF3fcUtm4FoQM5648fZ2lIAYzrg58gpQnquSssVP1rGdMnQ+n6Jdh9sT8jNg
Ughv4bn9GqE6xyWkSyJbY8ck0v4atyYtCTv+JCqqda9x1eOapu88oGFTxh53
EC55+PkTIBaxFUWoiu9HxUUAoO2NwCUnoR0ZSF/9dOxhMSjQBvM1gffMSdKr
LI3b19dVUcDGJdlfsoaZvXBSeQak8+PxQhM6HW5NgH8ntUwitXq+X+6SoyhB
aO2fL0WiCMOD7no7Kr5gwcnUpjxkJzwV0kfnsAHjXwFQJ0RJHXyF+S07KrOK
sg/qZatKWP9twS3Alf1Z7A6o/yxWTtNQXQu12ogymicdAfAba+6B8WfQLCPG
xzxt4x/tcdX1be6xs8+gCtJJOZ6tmZ5F2kXEF+DR4T10uei2wNxsSNvHitZ9
11yvPup3fEhBPYkNyjccQCivH69jKr4ILQaF9aae5wP/xxlOymJADNqbmTnM
AXo2BntK0oJoz7YsDMydDgXZZBbKU3z1OIN1Gh5VVLGhLUSxt39Tv78RfJbq
rpJebCS4z0RttiluAZRIPnzoBf9W7W0yoWxp8cjpAfIgEd6dHi6zGirFkJmD
pVTX9zEBcVVhzqO5ZvzJQjG1yBehVUAXVEjrYO9IMJ/pxTxUaQ9YCUodBpid
inmJkzcuaxFzKKTR21QxpljKIVwA8C+0gVpAv//HucMEf/bBL91fpre23ZKo
z0EQ5Jzqk5zqfLj5FVvwzF6aBeL5JPAXsHUYjcHdE+u4BTDrmG9JKwJQAQB4
gpiI7luINwV5vyzn5qFHqeMJX1hcF00yhXTm14xaEddISFqvgXM1fAAoPgMe
MUwxUl3uMhuPszA9veTbTO36tlxyx77YfYUZZa2eg3GlNw5AO6StF3zAWlk7
VaN/LGcJ3BS47SDgBUcdOzIZz3BTbxo67k3fpHDJA+GO4MFEJvWYk7Rgk1XV
RBv/2Pg2zLQS8dVx6d7JgveY6FHqoNSdEprH2b5HtmSmkqK52k8B/xw8J0gW
5K5rycKRK3exoHGjs2Dpouhc26OfZ6h5JN3P/q7vqUXyR07Ny9pnKbOQMUK9
JYKj89OIF+XW/6m4XD584jsgV7GssI9icLH6gH1HHipHVO5M3QzklTBZQerz
sO7vPgqnGSUmhL4YI6KJw/fCxK079WINjWw5Q1wwq1CnVZQouJUgd3YJrIT1
3MWufejmej75hu3XN7m577cL/Plo0UtY00vX+01AckEnmFXy2cYKe8SUVq4i
HHigHiTv2qDdHiAD/CmH/dPTwH7rjSsfSKP2UPDmsDqBmVIcsdUU1ctT9Ss7
1nwElhG/i7MDnuNppoq+AtVhR6kaC/2rNhiuIANgZkB+IxQtYtB92zV4rnZG
SxNS+jk7FQhScuA64g3XazvAnM+cAYIvoaCbr4dz57xUgatPxXZlfAp2sYgp
AqGB3mgkcV9m/PIlp00NZ/r3rqPYmSTPNBT2SO8MsAj4OREpieqGYfxJXc39
caaI30/k3thGm06u7mE+Y89icgKFoz7IxW1PwbYy4XpdREbcodcEnpB2Frh2
tQs0OOI7XQl+nIf9mcoWuiyH8H9Aq2/Q2T0bEviS5kZk1AXnu6Mf0yPsvGwi
RxWk3+1mx2TM3HszRJFLSWLv0e//IDUKlgNB5tMGLNFnm4lw6eWx/o08p6O4
H+lj/xJQ6rEsEREe8OsuokmVvQg0bDDYhD+ECgDfQY7NV4fZuztdrfeNm0FT
JdDeQ9XsFMYfjiUF8WCbQEwFnj9UxoWXw4Tl27qxBN8zkgFlpt7B4PT2ZGW+
K+13I2v7bX3oyHDy2MIydslz8sAuAuKBZ30K/wMZ/f0m815VD55GUL3zbDsU
KdSAOTtPt4Ws59WrMHvYkwZPMZr6Wfpys2AgyiTjXP47eLpxtlgJNFcHmYPy
Es3ZZf5MzJZnUt9OZqyDXixwYppZU4UeBViEqlz1WNeSyPuraWgrPq0nPHO7
XHtWdRxWeKluyNpyxyOAFcRb354ZweeIXxNwP4h8xFOrUt40x86oGVTYxEG5
W0oMs327rdfvYUBUdrKDlND2BDMD3deznsOh81x6pdy1Egg9Y7p/Q1MCiXWl
0DZ/jXMe2+dxUkl2Wr117FJrwaiN8d18kxjH7jzjZI+kgvwgWEHh+VZ6GAl8
aJxrCyFGG+XqTVVs++Ki0PHefnoHyTWhjTf+9A4c4a03hXKhGTNYJQV2CfLX
Ftmc4Gw0mQP3g9dX8uIOEjAyGqSI6d7k1kSGqPKu9aWYb3xuEdrR0rHha/dY
mG1PVOfHN+OO1xMKoyX0X9rRzzAvyzzRJYRYcv5CLPLJ6GFM7QCZGcifTvEG
N7gS6oKyiptk3PvHRXGUQkpncF3kz9lmIz7+jt9JN+Nl2uR2KmEQd0fTtEJq
yXH/QfzW1P5BZehgfeBrk8+v6sqGeIWo4doM6/95APVG49KnENYC5PfJjWUp
rGTGDNU92M64wK/OfQgvgnxu1XOCbFdIyFhaN97s9lLYSdrAKzLMUcQ+fRYs
mW3FWzNwQOsfFVmUoBybJLyQ9jzoIbOWF1jrbr/7fMxpWUv7KCsjdr5L+t7i
BHZYuoinMKR4z8WZOUYpZACNLHHDEN418mP6LF3iF3uUFtXOb4mpOmruvCME
Z7ZmMQFY3Elsygr6jLS9572FHqJvkb/WpbE3yhok9ZMCAEgnNtjcVCyRTqE+
QaXfcXMmqHRmjjVboHf6IIhUmA2fb0TdaXH8UtTxh2QOJyqGbBy8N/fqxnt0
wARbbDLbI1OIJheQQe+cBeKig71gyF4Hz4XvMtzuTHHwFbDQZ7/GiRCuKi9n
0TI6gUXz/VJZNk6cdqWXfMs6LBWd6eLnMvVX2MxtNvpBbZgh/Jb7UEffvbjh
B3gcSLg0b54mJ0xwgysMNFk/IObODEGfCpHpNWbrt3b36h6j/F7nUdgKTCs0
05JscO5HudcsflWVDAtLhCNxh5Gk7wz2NtH88m5LzQbCB8WXPIin22KvuJxf
WOyyC1PH2VFtLAULw06h9p0sW/2hxuOAyR3TzwSw/gvVqw7pCzfgBFBwtRic
2gAzECzASDBZCGnFhsCCfbHszOM91p+KOLWywomgoGA/667p/ml/J3a14IUl
uBDEpgCguKIPhAycZ2jScTCrc6N0lOsTI4YvY2RjyRQhO8Mhpe0FjcEckjkk
hIPgT4d+P+QVwel7D1BA9lGRhHWw3VxlpgxJfaSnGxKuzhRhkv58xDg5dCYv
kLc/gGtGjP9vUITXMzz4SHGBnADAJznQCota+OOGohP7AaEDgAyOYkhAcfFe
hhoGQDSOVaJiYjYGuDA/hwgJLv1nHxxMPF2os+KUniFXtCUcWcd2LfHanKG6
/P4WFlrDaVal6qoFdDZbBmWeRnLMemodb1+VoOSgMaQHnvxnQdSrXqbtcNFz
Q6aIByPwera4fG5V21RzuSkO+EZvA9uv/h+OJRkRs9EZlXQEXEYwgFAD4atw
oJHO6N5rNoHPJ7HPM5MGhzi7Mnvh59PIpK9FvTiHsKTzvsKDRhdpvu5e4Yhd
5mqob8vhSti2NuXkvJ694EZKza7KnOCUgdowAMmp5Uj0iad3vbn3o71ZNMJj
1Q5XK3Wfb4z0lgqYd+y6iuiskCY/5Gd6oW3TW7NGHZvRxIycWcGRglSbTrYL
6cZFdesOlnr8Azs7i446ldkJg1LZIyxmKHTIfgrI6iqrl1nSUP2gBwqKiVyZ
Ji6v4djwzjiR9QojEtkaghYaLrluI0VZM91YPPZ2oxIla98efj9C5We0EiDF
If5j88TbgURW7YWbi52df+xm1WQT6pjpRGbHvDvbQ+xclfEd3/Q53KWevxr8
oiBHKQpT5cJoXwBiOy/TbVXxZSVWsF4XrSbHMmR6RZrb8E/SkvbKmz8E46+W
8ObeLqfx481ccQh01gMVfHOEePwOx8yYQ31HPNSX18aLAS2unYa0gBU9Tzgi
wkZbIf4tN1abWbmTiDUB9vTeAlITBiZkbT/ky6mbDsq+1sFCwmQCR9tuvWHR
GQWrhslznWJelegfHqgc2WDt6zVbdBOikPulNtNQ1di96MlfnVA1DSPJHtnI
N16LDfYdW70k1XSShpWoun0JZsQMWjJZUTwXD+2s7ljIQ/XsgrToaDSGyV2t
72egwYC6a0RhjXBVsg+xg/D1nk0qN42MAUShkPv6J1CBBm3/tGJjKRhCtwlz
mHRrBV/mcn/++MaTBrrxbu0+P6oyakA9qevLcBJa1EO5/FuLlnHVSgDjjNGX
XJ2sypJpId3VsgrIX7I678Z+K1vaphHevWRZLhFbtMdFYm8oXkEZMOBm0zkb
3mdKvRYxVtwF7XsaQt3TnxE0yWmsysYg3GOK+t4TE1waP7JoK53XCvwYJBzl
RDh1DkMWgHLmxbDB+21/PSqZpCIWtJ7BwU4eJqCSF2v7OM5yEWacTI+pB1/5
1EcCTmICgHpI6aCXZiByZlmkVyAQDk/f96/CCdkghXVSYwrcFassOb9MJQya
a6eiz5uHciMT4xa+qBZPyE3UZbAV1IelXPg8RXqHTOGfjROWPVWnCdm9wnTt
sjUhPbimcUIYTi9CXcMuNT6X7bspKs9orYa24yUca8W4wrh3GaFevTgb4vWP
4ilf4rOpedQtx1PdYD9H5vm5Xn0xNtInfxetGjKD9nL0pg11jy2NHMpo7yo7
nqhz444lysug393ApPYyI4M1MPRMOvG5+/5qFzdqgfiOa21UURiRV1D4e4Py
FJ9PENTR2VnZv2ILTuuyDxSsl9vaqBI+2/K2HHqJLSfp+LjgjEYT5JYy8aGI
J/SqrbkY+9uwC0HNQEb1ds93mTkylVTS54bgYR7/JipT8I4TL9lXJN0x4v2T
upcrj/SgNGHpUF5wSpcy9HC97PnvrU75AOabyeA6uCVccXhLjLI9lIuqXFox
/CKCT/B0laX2E6a4qY29U9OxwHM66OLs3zA6NndtAcjji4C3NtDcmH6eq+QQ
9d6P91v0gs1qiWDD+98ojdAB2aBERT7hQ5C0pCLlAcYOD8OAEZHy45ChJ6GV
/VZsI0bolBtEE0aMj06z4ldcJrQPh95N+NIEgpXbnWPzCO/aOmFcEeoVjRLV
fq6oRcIBT8Fvmp/walPwCalm/7q8tDCIsSWM5gYwV7CPyA3VYobDTnR20lv7
tLcjEWE6hkCXkDFuSRb0kLapPTAIuJk/oj1JJ/GqXLVQAJGIoMS0Rqq7Ih+G
Vrts3qLeDyIpDgHzARJBJsQc1hMaGi+wBYGYVL/VoetkHfKSyzxeha7aC9BQ
Zx+E6PI876VXv0N+qI75+FVJvqDljoNDKkRTI8At3+GdMufGgA8oxAPSTfZL
Jk/dyR+XN9yIdn6DnHxn34TXnHj3aOF8hSUiSez3ukh6U9Jp20F8ghD46MyX
oFcf0pUAAhHpMWBP+Gy+rBhTAX5MsSG5+904HhuYOT8PMNfPicb50rGk564N
kKyN66HUBb0KwGsBJf55WiMY0+o3cgeBB7NcfBqgf/n2kb0r67qW3TaZI+tL
TyrjULP7aeuyh4DHHksBjhOGd5Vl8z7Fr+26HzBh0QFjuXcVVjCZ2O9FWmPH
dZUiuRdF81GK57nbHei+6qX+POE5U8r8k4v7Cwumha+2ml6M+uHH2GyRcwb1
1Pc7TPetDokjisGqPn+BoDaHl7Eq0Lj1hcUT8D+i7saWbL0c6HFznomA9c3l
2mZlWzvP+URKoRuXIuIS374MrUPtjfTpuBYZFDkYcK3bo8taujXPgVovYg2k
aqd6aIhJ8pSg11Z5in90o52YW8L6aAsxy84QX0kTjS6e/cwElMspam589EaD
phULVWtDOZJ/5g+bur2TYjRYA7qThuw/7H06tlYFAqnpXRsJhv65y3oTEr9R
zf9nCZyNp3/eY9I35CakmiZHptaXmlQxYyOLtLmk9YJaYI8C81ojSN4LR0wO
kCjVKivuUVKDhzsyex1g8QrI62lnMrrlvUaFSZWEUOLG5Fvzd6BDQ2/PKiuZ
WkOuGLDDxWfVgfyn3Ttos0zuBqHLSRAxbaom+9d9qaVXGGX4E3JczDXq1UVC
xxNtqLtf2aqInaKU33uh388aCSg7aZc4cSFylRVkPlH7lMpOOg/Rtuem9QAL
l1+pV75ddA+sz/ibm5OPEIkZb7V/dc5yQIia7HoIHSCD2RER8T3ZT0upTTE5
YH9fVZ27aPx6E/OdLKaU07/oJi2r+cp2kyInDty+vB6z4QRlQPlLHlKugQPO
VJaPO1h2vlqE5+UOuC0cafNSZKJQ0CmTNzajuDRq0ufL6hKdJrqNtEwgxShs
dqi5688kK1j2nWm56lF54KjL2HJqbDxJyMzFFv3wEvAaDGFHuCDUZbt6Pku6
uC6W7gMt9Kv5CPa4n1qxkP58eMAZMoYnSn72kmIxmV61LI7V0osQSDBgPNoT
3DuyVfWwCr6xq2+JMT7AZ18Zf1Gms6rx6wSjZlge6Ev9uwpuRbBJFItu3RjL
5XmHJzxaucNptHaiDg881MkaL5qwceRlZrto7z6K4vvP4Qr1e1rKxLNTCYQd
mqWf6XgHBw/hWQxrKBMySX63T+Q2cgHG5UJ6cqnhfkXzWeN8YrUPOfDTFQM/
nGB/MKXcd8trXE/oI+nHz8I72B9PYEmceXBpbY3Ru5Fj18e8yCfsJDNmbaM+
7eRd6jFPvDBnlfZSKA7UouZtyE8y8lPF2JsUB2iVPZ7PaG/CtVFi6aK5BHll
V+oceOTA9qyl0Q2c/1JYCXRJAYxv3LbnZvqdW7kMiKyRlgz+KzALxoatj4Pn
D7xNy3bstSjqRC9IFWhAUR/cZkE1KFl9aYmPj1dWGcA7W+xUpVBj1yWUfDTZ
kvjEuZXnYhB4wjRlb+KcpIfGRPsjcypMv7tYoqQYq5mM44JiQ0OQgCUHmINy
V6dlQa8AwbwtbJBkCwCHIbtY7j/5nF5uqQWzBLYXWkbftkfqop9p77t6v6Ji
Riyt65cfg469LKKE/Sw7aJS5ocP8ekeJPhns9/nMi5e29pXRWAF0oZ3xxQXD
64QQOfpWVHy7/oNSqOAjvONEfTnOyuWzb+Q4McESzBlKSU6hJZP5K9P9FLqp
MPu+TmaIhCTKb4xaBudt25SIR+aK7WmT1RS0ZJuqduYo48Prq2F4I5MnCGgC
zoX7aD6jKndgObTKdc1zVHbp7zyNzqCJhvei/ND8pGzzByRActjSNf4TPah3
+0IMbRvkT3ZyFzu7FbHY4mKYn/xJoZbGo4vjtZ5h0qGsSaeGUtQ7h/BR2jMj
UpPdtTXRH8L7SZJl8ZU4iGHXIwaKgGwA93qUj/XnShOdk/s9LCwIV1hqikm6
8tX+ZmLdFZcoYdXe5N8YPvRGmIlya5JvGJpHC1czwIQ7kcSE9UouB7uSvrAL
oj4VcK4AmXHVpeJ5LeO3MoGhQKkVBYLL1Krh5G4TsvjPXEh53/mXpOvhXTTh
vD/Ti6ScdFIY+KgFYwpyzyas71y4LGnzVYGViSefzqLmzQGqb7ALIVEI90Re
O14CigA48h2umYQmiY6y1saupM8BFPPsmFNfTOz8M384UPadSD4/PoIgYB8w
HeXFQxFPyb4ami9fVrSWThjoB0xCCiKPdvyqNhiJymF2pClLH2BLNzpx9tto
2a9iMDmFZbBkgjPrtL30mQfQkhYgnzDT8gV6AzjEBUmFoDhCneBHzFA22VCl
jW0bv7Z2IeeEtSlEHjV7ZblPMzTj/MuVYashM1xaVR6hrCoF0/c/HvM2eijk
DHavJDOqJSNi8s6RNEwV3zkao0ZXI2xgplgJw63YDwOUK8Y+CvvEykXHAc79
nW2w1QaQ5TX8IR5IYIBgFlHTAWFfva9Z4zfTXPyFGEt8nJ2fuoHHFKtzJlqi
za4i0RB3ONK0lDXTR/gdNH1N6tcL55NUTRSX0Gzwnc+VOuuZO4kfICxcHKHc
F6ENgdbLgJm0xCjqNbQZDS96M/mvvVRl7D6lTh3eGuWhuLyvwMRVC0e/a4nj
xUVuQK0tzrQzjTb4QY/kza6JRk/Ud2Ov6HJVTPhg9CiKci4EQjVGJghBxPBI
MRH/rDm4MW82xLNELyFGp3rCw49/ry22/qOdw6ti8iPRM75mjoP8thjeXJFT
3mIQHWVO0SE0ExnE8bSSVUGNdnSTm0ATQpj5cgEOiswku2qa+LWNyiDrBvFA
mjSiWNvyB+TIDBFH68yqB4pxxbdCpw/FJyJvjqLmIDUPXxgqbioK7KFkkStr
Sl2UrmXV/hA3L9z2nA6nQSslcAk2dgkRDGaxX5HiJiUskPvjfK5alm4HoRUw
hQOjktcf6GO5WdmI3fTO1UDxdjhUnOiVgYbVjLUq2pdUPqY5fCvs9HZqIXDR
ZyLGb/DbLqPn7o3aGBEzdmtYDUNpRRCiyOseqFxvqJKn6Up4E60PLSLLZjyn
8dwiAvIHbcs3DpMfd3aeO/G3ZfJ/AE1q+ljaaA6f2uLTLoPjEIwFo+trnLrC
aMOkCgeMoLeTXrmsBld5QtllmlJx+54fmzG2YmyCi6wriu/Cp4O3F9+QVrxt
1oWRopzSQs638vP5/nAHP2+Q1BKSyQxF3h+SciyerE/nn6g3bg4Wugz0xA2M
9xPJnms5kJT3A2JdwaSdHjgfM3l9hUcHNYuG6nWto41E8lb0fb7cPVuZvdPg
O17m55M/UHR9cIINufVl1N1IcaL1dYuRxEKit+WAtROip80Y+YzKFW/Al001
6yagMlNk0J7JfZ2R2O6y9S0NGVFCnHUwWwLZqWrjEAjn/cTsgv3igLcq8XFr
Pkyw/BjQWaA+iYiuNmqmU4NL0ateTyl3XSjA6nriRcUQXhNFtBJV7c8k3kMC
PGI94ovXcg+n+9DlepOA9Faqk/E+7OK1VrtY7KYE2i6gnQeKRcE1cgRJZzkD
hYzH+1l1LF3vN2JlknVfhkVNTo3I32euirM4fbMjQj03At4SfuSpTRA7IfIB
WOiba+EAMFgjuBTFvnWSW9MaYMied13DUv34SLCZKqUqsHZENyH8Bdzz5k4j
B1GcLqN388JX2Is5k5VKQzuLfdvCMPuw3SRzOslfLkGs48Kd8KF2mBSdWkFf
ubtBn/VVnoearLeMCrJ9vThPic0N5/dII4AgBRTNshaC6zAior7kh2D9K3Bo
Jk5LWTD8fDBKk7JMUENIz62kqWeX/YbElWZNJyezlyoOHAFvv2JR9Q8W5ev+
+yRJ+zgB4SjaZja95XB6uFlsmgKOQyMA71WO2gYDdA5RlsVGp9F9IkaqLSkT
O/HPMFHcpIaXPMScHR82EYHrL2dCt3zgqABi12gRSyX4dPLP637qlartNCIl
Bxvoh4W07D1RLgsDRBqpCbblTC3xNN2rl11tqjZshp9s3MGjUYpajPK4ECXX
7ZvZDTnAZsQ6U9BiI+JUlInU24raTbf5uYIFwdDT6aX5r7rU4k5meDKpoldL
ib8cu0AO1o1ADD/M7RNvpWS8ofDNaTJ3e66joWZqekybfs7I3V4dczTQr2XR
zTxHOmA2dUB1a/tBQbZxT5q70/XEayLEjdvH8qKLKaNKxPOJlwtJgDkryslJ
fkehJJa6Dn00oS/ZoLN4bD5McHM4BZ9+UIBGEjuDz0pc4/4JRxUwpbq5YOES
gsWeqJQOIhN13xIDfPouB458wJJZ9rnZeIjrbbbl4A2FsmDu1pxx+PWmWoh0
PR8HfHqJpWe8kaHoZ8ruytQ9IkeTokyhTCH8Q32NHvic2ZX0jO+kfwj/jRsS
u9RanBDtSsr8SFupoSiMB/nVwVSIyJMlTF7KjSJ4FP6Ysh6XvkVT/Mkj4Lju
MxFP5W85dY9T/bumc7MgFos9fvia01fmLNd9rwceHXSO9WoxTnGjmI9HTQtm
gD0D8Lrwoq+EYB9XKMM31lGTlOy4qORmWrEqod8WHK6HlqlGSKSeNBESl4eJ
csINKIY6s2CfrXT9G6vVXQr+/GTGbsRVHvl2Dst86TMu8Ah+5hJt0NDo/9OX
tVfGBT+zsVG/twvXS8LSRZLFRH9Qwr9ZdqPlMN1ClQ1kyFNMntgA1/YqV2Zp
DjrlzK54lFmvHXHfE34wryrQf1/W/XX6ijF9MfoBkyEInNRJiGPcmlXbs5x1
v/4ZJSUl1AhJkpKd6Bon7N1BANkcetW08RHdO1t408DdMJwAYg3eZI4tbrAI
fopHRlZnwbNpLrQa6GMTqRhsAyhkHls04Ir5wlBm0iOEt8eLMmuFYmFszwhs
uHkxMpVNagvOI0yIk7C8s4UDGlMukUzPQiWcaMIb/Av2FpxYMNC0vum0VZr4
87mMtscvOnpIPxt9MoGr31Eo+MpwiolyCeIiXniAPI3kTNWrdFnErkvVj/Ah
W43hfuL9+jSdnWR02h/s5gzhW+KE8UP/7BqFspCpA5aDwHYS/ThesunZ1VXy
eAsoU675D4XFuwFENSZa2YabulxRz4282cXsciars0FMZZ8O6EO4jt50Wr+Z
2utUBNO0yPHzmQ5zkI4S3dG47FUozWbOGoW/MaoFYJ7BLUu153W16p87nSKi
O2bK5fwwy7ZEK+i1a2VaHwjfXFFKFqGsqkQDRbuW9GmlTuDckViRhxpKq3JW
65MXe5qamVL7poSMZqg5WkZ5SOVojN7Rmt2ZDFyFKslXvZvqiSTDqTGw+2Qz
cBtghsFAAmGcIldFIJcpO7w9I8fxxpfZ6joJJybENmigoz2IqZPVu09/giwx
9h6B27Z7+nmHRILB02RS4FV+/z8hSDshoiofnTXjc3rPvT2lGLCyr+k6N7ty
IHNi4euJIqSc/wFa4pT/JP2s7oHZ3fjOWohxwmaR3mHfWvI7J0MNpY7Lv2jY
zMQcutBEBJrSIWULO8WPX+Q+9c5AeYPjxALK+Zlm+k+qrG0DPcRzrCWvsuCX
2yWE6dnhtMoIV6FAfcU5qugSon3D5UdUpLbeILWjJeFy8lWaRvPaBwELIVId
wqifgIGCoojbulUZ7w/Jm4ConkwvVIOVeIWdP55AtqIQq716fM35c6xvJ5gb
mUWL5qT/USEgNrsvz67jjWd0DPa56UfkVlZ262+Qt5YuSKbY0h7h991KcHlR
PlgNiu64Rs6gzuSJARVmlT6JkNZ+ASthYF9DHn8rn8eKMJKihLNEmbsFcV7n
Z0WWiPHPnF/AC3x9XLpj6S+7s9XDOf/sqiQr3ugMeJWQh1cDp7BF8N8hvxQo
K3yL6noDuiQlNykmhjZnpzQ9VCh8bQTal+csXvDRtfBc7/b3q9Y9GlC/42eb
O4RpMHaHSVah1OuAz2izlaE2Ik93pv9c8waNrCau+NrhLPzx0MX9/T8xWYmr
XkFBP20LdvkZNp3g7gTFXhWsHKBhs654cLR3b6GuBNxYeNsxuBdapsfbdz3/
PJOyyqhak+lQq6L6izzCw+9ji4pwHCpgeGQaPSs/Sbz/zI0Ev6kUQfPzDChf
cbIiQThF8tAbhc2mDyjLbad5lirqNi/meRO7DBIA+lrK7GpujBpl16XTBgY7
2eiEZUDr6E0UE3Uh98fKl/ITwqRN/uvGIUXhaHk1TVGegEPl54o5ijhcitJC
xIzTziabaei2dSdVtCe0Iv8VmPAg6ERFfr3V907214/wVyxhT4PecAlVYlgs
GedYnBfzPSvFT8MwIaQCEgk6iKPLMaRD2WejFfDb7MDi5cFlFK5/HrKXeyxT
A/vTL53H1pugaWQBjsQhjkJJYltpr0ORRbp53X5DPwF5WjT5fb4ldyw+HhV8
3ANvy5oQcDhsceLhSlXw54ZA7RL5z5S87pJ6NRue1SvQMoCq/d+RvxofuyvD
pma3feK3JST2q+1+iOdfqoZP5yigoiNd3GDr5PTrC1RSyMSqVfafE3oxSJVB
PiLxhkf4cnk/taEqfBD5ChsqP3GhqA8/qtBp7HuQ127RwFOa/9rl2bNKzY8b
ySXg83wNjTHZwFcDrbfRF7a0FQO/5CqdJJ8tMRZS7FwIIZYdzmw713uFU8+8
31Ci7eiQqCmhwulkbRQPBr0O81rICRgJqTHIzYdEzIwPdTw6iQhN+EDyYC32
O+O26q7nt2it4ArIXrF7nuBEGyvw1k5R1CrNx4u5bVkCVtFlsV0rlWeSMeRg
tCdk7FofZYyfySD0Tx8Bddl/B2mY13V969zv69LJUzwiObrrePhnenRNkMW8
mgUuRqRc8ilv1SmLrvMIFd/fNY/kmoJuYjX2tyvbAo0owp6/boe3biW1Beyg
WWQTqxk9BdcXu0/JDxdLH5wV5Yl5is0XzLv4FHSff8ebKQAIMnuFe/JzPIoL
qAB0u9RxG0I5KziLWGfQyafcNyU0hp1J+WLz5XZGHzWZDyftFMgUZ63UbrA2
GCcKTyrtc27dCg1nvNbVbPelX9XMnuUfeBMdWexcE7D1y5tSQNZ/jWn7WbRI
4cCHDPeWy5nsihDdEYbsNo96XfY7UMo1kjjFNKBJMsaA/es+XmWPNrbl73y4
nHQi6jsndPHHQPy3233B8I3E3cTQHeftktKYa9IEVSID3qswh4c6DTV9Xooc
TSAO/1YxZbmUUNUoPiq+YVfVqh8T4OeGbzAaG+NbK1kHmZDSCRhwKADojtSW
lnHz9XatTUGd3jIKrRsbkYYPAFOGlh78NYlwYILI1agp6vfnUAUU5N9J9AkH
+7yLbKFf3kKqDSf/jhdqhGzQUSvVcP0DHBOZfhTb67G+08ZnSrY/oC5TmrUN
1KWj4yJHTfaUt8/oT+ej0iI4EmC+GhGFUhv/LMxYty5oK6VZKDZrCv9E4gv9
qTksbWNQ3Bfy5grAr9/9/eIHpffpMiiDuzv5ak7rx6beyZYBaq9/fjwBm8O9
H9jPuP7XeDmdweyYPCbX4nFag5c2Or6BZ8VwQsIekiDPVfdySpvr/PelYPwV
n6dv0Y3HHKtkC3laGUKXlnPnc8YfKIYd5ivO4dVPizjsKhXXMpYK2oSugG6E
UJbBA0PcXswQtmMOOu9JwZ1pcJhR9sTsKVSfIRZKwmDHFtgb5s6HHHSEEy/R
ZxVIyk6PTD+qBFCQfVYMRI5Imyd83LOlUYDJQBtVy0IrtYuLmHCLfIJ9N53I
ptAiBiWPq7GUAr9TLzMm4LOzfK/bKtvsacm8yAPjlHWjR62wxY/9drcejeaK
w6Lo9ZsEbrdSw0MTo3CfqfJuotCsJPl90H+d6AEIW23qxnY3yDOhV6aj0F5M
RKANKEln3VKKUFrTojdw3dmOxKB8KY0L8uXVbyNoOb4rWM6gaIQZTdjos/Pj
1H2iSuCMmJbkn/mgnuJ24b7VixySVmWjTS68u0Em8/rHuyOC7tceuTc6L4NH
TRj8TmGVJtG8mFNa6wlDxEyPsH5Gaq+tJR1db1xjWJhVLBVHmGenFpvInhyy
iJgvmIVdVsXs4AqFDFxZ95eyT8l2FqCFZtTRsBGEDlVFdHR9jRkKWV4X4PPT
SdmdySlhoyrW0ijRBAvmgIWWTEOG35yqFxwD9Z/it43rLx7W2UTIe69WSOWX
XFVLXK/lKSyVQXyVtxtP6znKNyN3XNUMNpr6L0ffZXXH8lpr69xgxhH2nr+0
cDt/xpIzrL0DetyUNvx6ovK8M8Vf1tIrOrsdNz1paMlt+HdcAsa5cXmFFa1J
rArvzYTkuRxh5J7iGKE14nc0wrIbcUfL3GKlSWpbk+X0GVh8tSNBCS/A2iGo
qJdm9pWboD2I3y1Dw5/asxHkiJQbPQt8XUPyomkX0xE2Vg7+JPjYuWuVyMpu
cXBTx4iyk/xOI+coiFHVtnYTC/ac6rufnlQbPGbxBFvZ11AQyjni96/4qacQ
3ykin2M4gz0eEqJ8uzZx/ieqiNm2w2k2HSHQf+2dY1CzWt8Pvto/v4XAGP6p
lEVrv91T2qULG7jLMAP2eBlWewJwx8X5b9G6qDRi3gabMj/jszI6DqFGGpYx
ZYSD/wRbumEtdSnb2eM/smXNSFHfREsBb2qeS1oN6WqCgbezURp8qkXz/sZ5
bLNJ14vZ/AZKxXTcfw4vGz3pKIF3WqVMQbNzYxbewKj+qbTVnxbylT/27iF/
0Ys+DcjOgV3pCLtSDwaeBEtPMTVwR6pD+sYktkfwCklQHw4obrakl0Is8ur/
n+URBpIytc5EoA6g1rUriZCO8L0wjr0jf7nnXWGyvy9xyOzfeI1s5Tx/UGmN
BtfVQAzqWsmMRvPovjiJI4+8DE1ayVoUsEKfpxsMk+1BFGJTSbWtSrwq1JGH
4J/VmfNuq4OVVsUXBI7makGjhKiMwkuDoGvfjj+t8lpL2Itx7ulFTLbxYGTh
QctVyLr5b+LJb0ZFaf5xbUjlxnsfVy6m6TGq1BMmoLuY2lHKE46xZhCaJKqr
haOFvAp0Iyo8MSGgDumZCCWD8sjd0PUjT9HfE6EOcabT324HhEMDswJ8oyFH
Fv2AMgCsonbIF231CZPUiPzrq6tH1mF5j8UgizxhK0+ufIoF0NBCMM2GpSrN
xe/24Od0lRF0T3hEyiU21gkqkX19JoluCmKkvGsg+XrrxcwqCEsh+8BnC6fx
jVqzr6U16pcx7LfxVUYW+YVrYyV/R6+y3qfbcZ8Xgv0iBGfcB7AeS5AHaMoL
taIzOaF8PIqULO9ZyI7kDLRQosdOR8jyGs/0C8TPhg++uQSjNkdcDeqMP9f5
THGyCtJi4Kl1QLR99JXx1TqPkXKGGK8Za0BwOpLgE33ZV8i1jRpR3ROeUKo/
6ws8cGf3dk+2eEmfTTJVF7d/YFwmTdNGgngs4woNulbFDeGbuyI22zjgfgjK
e2pQQR+3FQFKsCxyapDYA7q8ag4Uz9Huqm5Le8FTDe1JGIbMQmU/pTyUDKXB
bEye4fG/0ID4AZeEWk++5mUftTvipV6u5WlwLg20Zs353MNofWQ3fbT8T9J+
Y5RsRPtoOpMeOqGaxxbDKdT/ddp4t7Y0Z+AtQQcji66nrKvfB9mBFFAnfQT5
lZMgPZy3XkP13jpJ8qs6QNJZ3+dpDEP0ErNc/ET/D1DeMRZc0NKLbLxY0pq4
Ns+Gc/xyq/50dla+3KGLjx1j8J8V94gtdPTpplfcHc0D30AZkj2x2NUTEzpt
8/Ee7rBFGBT59ux8l0TIo+qj2CoPSDOy96Ij4KkjrTg+8/ZmEZCjgPZyEJFB
EeAiLdbk+zcHR5l1T0uJw67cWGqnLEABwJlIAlh7ogbPTWLpMkQF7y8TllnB
7ImTqMWrZ981aWbrzKHUvQ3dFvZ2gqOhwCOHPXvAglY4K8ezfucRU222hB+/
XVhP2Bx5Qerp4r/TaVyrXs7dAPtaLGrKEkPQQkktzH6R25ulHwjkmRZs3Qws
neVAVrALOi8Jlx9vudQ+XTkRS6HLYTlrThRQtpoq4imCYPWcoxY/uVeXGPhJ
73kT4tMmWVFwg2r/uY7nq0zznpNfrFNfYWGw+U5iwsbAUk7VxLAjobSslxPq
rqn1xFlRTpKqknbX8icju3Skn1WN30uNQdHZiqamH60RJSj079MFezqmz9VS
DTPUUDH4+T611zRUdEhV5TZxGv5YLAms1nT52ds/aTbZ1ztHeis47pZq/H1f
gPbMatQE3aiu6fD5Uc12oHbp7MaMP5gNJgozdIj1nPlgentWzw37AATOyGq/
Iu0cwZwj6zZ7pSwVcWU1/qeUEfeJTanvN2B0wQO3BBMMTvG2wj0dJYdjpPjj
5MdUjX6LeOdZYU8WT0RWFANqvJwXbVaax+RdDPZzFJogphVHrBvcYD/Uocwe
18KBaaI9fkRM4tcPs5iFlTd+dmTJJo34uwprTeLp3Z/3omEDBq0ZF5u0npCO
JprLjNUTsovk/dFNoiSzxvts5LcHvjlVRTrjLxx+8iB2TpOW8tbDLVqHvi6O
dAE0IAswWEXEnaQxEbVkpmjcyTVW1mBTYba9wBuczzXu6B72BPqrrQdPHwEp
EOwddgqWa65Jm3edKjIjXCvU7tcNuZrON0Wyw5533196OX27pFzCq1t2NcZ3
CwbpKBh8XZk69EortmE03rGkxFypEl6mi2bATP8t+MjcM3WGI5SitBYRY8Fg
usnaESjjdwDNTNIuA/+4eAfESw8ADfx6lAJmkUe/Z5BM2EiuPnP8i9VGAwrl
5aaF6EUp8jiGC8QS5CD/qzbv6HVqVdH/E5jWiVqBMDL3/dLFGtn6H86PNq4A
E6N3djFkyEcYNZC5E0L+j8tC/8wCe0sDoVHc/+6bjzW8DmJFktngeafnVBOx
gCaC98FuWeWUf9o4F1ZxtTfnNmSAJzqoInp2WbsPz/Q70YL2DTW7vpGkjKSQ
uDkjxdurCdmXwgjK9qRqLL7mj5DD6d3RPLFAKRfKWjCaR0OX9qhpldOGGqCR
RRYzFXEF53ihSuDwCJMsC/4+1ehLre9KLXZugOSvrV2ub0R44W3POLQhBIRV
6zTj7/G8zSY2KO+vxC1xZTBn9NTpldhe8Vp/ix33SgwCSchBxCtQ3uPnXT9s
glRVNks535DxY1hI9SaWu6j9DB/vq5JOto1OvIdNxKEFm/Hfy15Xnzv0xX8i
xW0U9ywvage6DRjyXhXLb79gFIodfyT87zvB1YRG4Ptmu6d50OWTakHqlVcx
AQ3oPPLNWIM2a6bp17+yhCy3PJiqgnp1pCBtXol9jB82recruIxUnFS92rwN
sHWPcmYpE170cPcZ7hOBNEgYI2yE8UeSS+rJI/4wvUIwNDIQ7GhpiECoBbE2
fN9eHZHshDT3F+2R65buqJLCMbjBc6AmpLqX4JBwlIazRCIxHEh0prg3H7Xf
bwIpGZVFd9kH9+OGKHaTvW4oNOWpK/A79eMeFZMGMSogujkGxYvdG3cbG4z8
ozzMJ3AfTUSjSAZytxug6ApUyZ+PUp1mhuMxanp+k1I6EXdt7ULKL5mk+1Yo
53oS3DTPqsjEYh0t1v35S7AVWRBrZhzeq5MuMk6/MJIiSup4gX3VrzXhrJxj
Lauco9+KKi37NKCRLg/rmZqNFjsjXGC9MlzaE3wIJSr2mzozGvgXx3chDDap
Pwon9rM0HKDm4cJcbslK6AGAWfmMTipmPtyE2K7edDhjMO13DmuC+i949dvn
Uht5zELVdWVHQs83wgf9S7jkeVr7oNp1l596+1cMFpUum+VIcpj6CAc7u/YY
pMfQtt3rPoud/43TWqkF6DevGCNQWpRQY0hpqRDXyu6EqdbZv0/Bmz6QRv40
PWaE+HW759dyOvC/VfRmgxR/vpvuAt4lM42vgxhGVUo8lEuWSbzOOU50wxHX
PuvwFp4Bcs5H5WgEWUyd0EwMDxaHmNELMWyxx1mcS2OYLsl7PU6af8pj5JaK
7hDCGBUNz2sbWQ10SsXNZiTQgFEJV1Cri/THWCAvEjUAL6x+hNpWafIH2T6H
GXmlM28VSIyTeuOzHaB6lBsiSmMjk5nKMOlLGQpZ3wY9OtYBrf1jWHU5eMqk
MkuxLfggpAXWVMdo7ob3gncseyT4O/3WbzUUkLKDG+33oJM/bhZBE9uCGr1w
TSdvE137WqpZkmBfEp+JI1JAXA0rQdnb9jpTKiEv0GvwL2uaJjuWDRCXhp4r
B6OmpRtiWYpyIk/yHpUR2852f0L+cXVRnTctE53qLENGOR05IM1EbfnWOnic
Mycw+lyvyHaaa5uxtddq+BxhvrPdt2c/oNYVRVDIBqr0/dk+yb3cnehRTRPA
qmqbzcIgzsqt3iXPztDE90Tjvcdm5eEjkgYzm7wWrDbFmFgsxbvFj6p3ZuAe
f1KF+TTwDl2CPA335duQybskgm3mehb4tg/QhJuB0AVWNGtyLIuTC1TGjkHE
DA6YWbLL8USU/Thq+kXUf8LF5x3/CiKUwBA4rIgTLNp04j/bh30GriSacSIh
tTZrST3DN+TEMNLm1bATNG32whHS18P99ZQXNlPaLIIgLNR9NeprdBYUAchO
YnxgfDrBUr6iCLHsoVRJV+4oq765vR9vtgh529lu0AIJSZ2ZWMTLSaQBO2Hw
fbCVC/Kr6KcrGKAheXPf58BhVwn+hXrRCxM+V/z2p9TaAb35P21Cq4bnt+L7
OypXS3RIAeNBD54C27XuuLc3bCU1W9xAQFk/07qIKgnKQHvL2yk3/2YzVuUw
H5LFcYkUmP4pKiDo7zFOkk17h0lwco661CniR75GbRIsmArQ1S4BJXRh8xO9
rQ88qloMR9NBipPuPTHrVEt1PBIhd3lB5JYwWKQVvKW4PRDYF99FZBScrE/Q
EBy8nB1sNnW1FfY3J8hLSnmp8VBLIvtiA2L6HwDk/0/VJM8M+PqDpQzOFNpN
e43aMPn6/U5kVowDqXMykXnztlpKgigm3e7f47IqIlmEzl2FYbQVQcvBeYog
zJphrrJhqq3go8c4idcy3jsJQ39XZaiqxdX66dfS/MpUbhqDfeJmerqrcycJ
FJigRnoh0emVjRBSbeur60G2WjkWuZqjdjqN0yJrRAhORyKdYSl6L+on3rgl
Q7ZHra7+aGbktmfF++GUQj1ie9d7/SiFD36Urv0vmQsIMGBYjw37Uy/q9/Ud
+3IcyG0B5+ji4cnQattCHXsGL4OPSf7VRyXQL/y+fBRDc8+oq1r0VxssMuxQ
jS93JhVWg3rYQVE50O1wkEpc1ZTD9u7BAXipmNOoqMJKv8OKvVijKJPoWENt
hFEGIr5ZtcDACjhQtYXjDJ29+pecRz7ETh4QaMJpKuhctzLZLqZxHkqqCa1j
XqtoYMf/3Ql6WBwaldSLIgMWulH80rWIII/QiY+zRV8vuD0/29aH6pZPxEBG
uMXmabnDIdkCe3zk6ossKDUQYxkvEpDHI/LpQxXnLv6RZugnGQSHSB1iG53M
5JXXynhNtXUu7w1xr2Xh/JSNVU1kVTtlM3KVu3Pihccsm2d8FhiYX0+NTwjU
IkdKd3wCup/dZa8NDYrrsMfc6hpgysKX5Pi2lGn8UbTT3F/Vp8hnnd9MJmpD
RXUme8ZehgL6TN50QcGVhsR4e8v+vioG+vdJwwdS6q/NgdezEKktxnu7vXMk
q7KVp3tLA5ODUJt4/g/Ia13A89S8kfySmQfPIwALIrHM+e2PuuhE9CBbABm+
TfQUsKEojpqmH960KRA3TGEJX+928T5g7GKUKs8Y3qAzvJW1ocx2WOVBBvTZ
GzwcA9CWoxMVPPSAPkTq8i7TCNOCtvqSJf85ZCewJl3aFVcdf8MmFqj5ZeW9
BjPln/zktfD2VfB+FBRZyomUz5pmjlaYXI99rLuTcdPx5kGRQLnfrrm3IDc6
99bM3mMji+F74VWxbRgCU1DLZcDWWVW2ns0NLpbv1aMx6jk28iHCMDJGqMK7
gdJkP6GbzBLNFGz1iGHbA8v/BUDqDNi6H3tm5ZYnt9VZ32/Nu6eiwkmdhR8v
sNKh1hwT2hbYLaYbi4MaVJdTiPBaDv2LSl9llwTuluE7scxX+3imEGCW8sE+
5IHT41qp67n08jgI79GEe4U0CxyUUyTR4NUbAZvk8oFhyangC9A1oALeRWqN
z8ouPMTan+P/o6ZwgjKT3aXaBXRdgnfqG/pTmJXXY11dOTsNZXfeqLfA4A67
wISUWXMZTuVU8ZNKx6BT3HZRNy5vWgUQmdZeq7o1G6GVdOFKGru4mRcI3v3l
QchS803j82nL9vuai9XjS6n92pEKa5llWpD41gYZnKpdlKpH6Na034NdvVHb
QSuAbFqRC+Hk1Z125xzKh/wtudpdb5yzygvVs22qKb7F3XZG1m0GBBKbJYIG
skX1A1XFOiuAYrivsqOiQGHj2tqkw9iLs45ZC7DGtABghzrwRdfOGEB/RQF9
DR0kcN4hs5O9b4HJDGaSnAA51Xbd2rxj9B7GhCPS62wgiKwb/ac5IgdigzYc
gH+kXhV6YdJmGOAF2xmwYwZ45wGaJLiRdtdLTlJ+7843uiB7Lq7HPbkdLeab
vx4wlyr3aBayYxTbJzYQ64ZNs5mbkw7e3OzktWM0k/Q13AW6kvZrcxFbUle+
t0gGmydkL1yHy1o6mOLzTyfKCYcoum6EgGna/TkfqpK7Ogj3Ms8QPuD0tEFx
9e2t7eop6TcV9pAPCftc6hBzxl1LqgL539R/gcPzHr8EtNU96MmVxKDr4q+p
4X+kESyTM6/rljVj4f8ovZLkEK6dRpmMMio/aYqkb/+C97Qu6nrhXumOXH3s
5b0DgTKmbWGRO+3VSE9+f104vBXwm+Hb2ndb2jZ+GAIvZRtdGWzng/d9ywlF
AWcIyb8ZPRd1Z6j5fMlu85nsxvx5Bp+FN0EXcnwPTcHgMKv0mSYrzdUwRyOo
js+hZZeBgejbknaH4G13nUMTd/axzV+gBCQyqfnrvwxmP3M0Ka2HPleNUD86
0cZ63fnDpOunzyddZG6jbIwQimmX8w7g04Yffu5d2Q/uS/v+0Krgq8JyQKFN
bkPo5DTv5E+6nVCibU+hKQPhPDp4TLl1zuRhshJEAgOCayleR811rb958e0I
RTr2DzTBhjpJBHbCH7EqfX9Qtq73wRXmw3vT25bl989Z4H664orr7MJ9O4QZ
JNUF8AM/Imxg/Trm2egdR1UtEd2FC8ul2kNoCQmadPV1ZZGBV91hkiTEF/YZ
5kpAe635f7czXpwmpbDQGA0/WeWCmBLKKhR8FVmKhxrI6f5MbBusmz2guOym
S5bCeCKrpuOvsnwACLnumn55bAqP6ven27kpTXcJK+xBUWI1vDFoJHMu0Z1L
/QFt0jMSQh87pHGPcVtnDO67iQDKkShf2+m9AZG0rSENxekQmQKHSXy6ccKg
pq8pe7Ypr0XH3AyR7gF39/xWlj/kCjqqnR0HlC8TVt9CrncTKONuSRznqkDR
pLnL39BcZJi8FpBgaSg6/unUlV5s16cFEBfDD3ZCLBKzELehso/98ga0ao/n
fSH68ULVE1TkWOw2mcglHV0U2KrWbk/6VJqe7LzeEljnNa1rbt6RmrDhVBNi
fFszktClGql9xUS3vPHxafNRMBsJC3clPVr6WLbdTkzPeKi846XVDBgn8TNJ
iMZyjg+F09tqFPPaWLcGEOsUHsvjrzpxvayj6HMBNAIupRMFHfRSmJ5Wtqt/
XijYK+C6wpwXW3zh+dpJ+NE+A5pj2VkspC+FJvHbiDJ0Qcc6vjSuHBDwHzjR
hV/EkOqowSZlHJ/55Odz4Hq6ahOQ9+8V2WeH572tqq/Rl9GqZW7MPgT9xfyN
U2XTQmvuxLsk79OiUb9fXjZQp5GbXETJ8qY6Gt9gYP0zclLgr+MDPpWurUyM
YiUfE3JOuXJWKWIqL6YRITPWz3kFT2YnwXD3uzvL5lacwES8X1rZBiX89HcL
jkAWSDcmOOQZdZQYS8/f1E4bPPlevKAMD1nrv+PukepdbLukNqahYWjTUn9z
OhthRpuarKcirtgbunj4tHCpRBazlTKIVM43WJ0IoGG1vUJc35BwABIuZLpM
P7gjjfH8K21jzb2dPQ5sOPVWlmTjMNCqMK+P1Tz6Ao+/7J9Sv0Z3fz+0EIoQ
x+dIbw7Chb1xOJCUSXZ9j7ArzscT6QUTjkgA1wX7YceQLA5yYP6RR6vo3Sng
EVvbVzB1Kakdls2Ko1YtGpeul6FHOVVUaNPmiZhVe6FMFgoKPvLF0rxSqksR
58BXeqtf2ReQlQL7Q7eqQptD39e7L+pc1TbnSUAFxd0AXEMZNiH1kRDerhPa
650USZv2hLoKWLlcvrrSFKQ1M31wlZIYW474G4KhfoPan39HPUCMbVIqgqvy
McZx9qOb74X/cjqJBtfhsCi78DYN6WUzJMMdcIW02M0Es7Hc9rquv+1gzKh4
RvwBFKnFRWYZjv5as5FAv5tfiYcG+b8dCR3gufGXteKweXwq+2WUPopyIzmt
qocOAym/0AzslJWbWmnFGN9U3BrWT/DM3Wbtp+m5GiNM+Rd8HuNWi1nd6yIR
GA3QLa9K3HpPz0eYr8G8Apmv85Kijz70TiD4z3Kv9xy8KrjCxpPM29qYFqSx
AXX/15B9Ogy9k8uTHImMhMJkbY1ievp3gLVJ+0h1p2ZB3I3wiv7kxu6NEYqT
a0lrYbeznK3Wgze0LCjJHjTy3muTPsm9R1rblSXlxp/ktwKbNV016SZW4qkg
QaKfS4Dc+zF8mf0VawRyGeoBlIN+yFX1zug77R0vsnnQPyusnfEIf2WRPbee
/z9S/E/r/iyqAlZ/wpnpvdtNdiIlNZYK9dJzN3gpTqkmbVO8mmPOHP8DDzX7
EwfLzSG6vX9/fzz3RfXS5c66iNpIKx2d+1MWtScvihjbcxESiNTKRH7tZYux
I+StYw+nhJ7gE1AW4tTwMhV8l8ZsSeR4wysHOXMsNRqYPBvNASUqxHnRvWti
EbK2iczLnhVl+LqteG6h09FMYz45+RJ++jZguP72fx1ahhoJy/oKvhOL9HQN
+K1z4VW4bKtjw4MDb0EPjodPVNPcwXwxCBGUp2bP+El2ivPF2mfbLR9qD6bp
iBpYuq2l+9aiJ+ijol4l8nCKvUnLipngldyrnrqmKEX9+bjEdcPDOnKbhv3g
ZV4BsjculT3+43JtC+mRsflMbfIHY9mB4CnxCQ50ER97iurW55K0YsA+0DcT
Glx3PbtsvDffXu2nWCVEDK7PLLMA7BtgcZmQsFRA2Y18rUY/cd+DpCTpwhzr
GELJbXEXRbhatNRKaij+xkND0zZXooxYZcu+GGvV84VY7ujH2+DpDoUlkM1r
aYTS5+ox9bDzdpcyX5AhcM558BqW/N8MpggN+yzJA+/mLvSkkqWLTekCRw3e
S5+HP1qSBFnV21iQFlAiZ2DwIh8kH1RE0uJkqmy0AuQwXvAH9gPU8eiez5t7
D+o6WLqBZPs/xN2CYF9tdp5bUy+DIBIhzCkBWlJrHr+/9BoNHD5KNb/r+Go8
F14XXXPcERJdvcWmYOxCG0QM2QlXL1tDflqE7zckQsqErEdKdZpKHpIqIGge
esdZAEisrrCm5oVRhccdZ+pclBUmUzT3SYUPyBTXiaIHJ1KkTLL+KIRjHWCn
ztWvPwKLRn62Ug/KOXH889wM9EI4vAEXK7a6VUFqrbkPX+kXEqUqRRwRhbVx
5HoFGLEzRC9Eeu4TGI6Vc4Jx94aqS3vYGFslbAVLQxqc3X8EQDWcOS9ABhEa
dq3hJvTDpBz6ROZUsZqKZ/Kvgb6hD6FkYYW+iFmAYEVgtQOgWEbX2MRIorfp
A3IOU6KZnlxfWj66GKGYAHwqZzcUKcVNprI8kl2O6uQ+2vbJXcWmgcb1kVfI
9wMYM5ZK8Gt8r3wQCgwQx6I2FyFy//gqJ37j1a9u0cgugUAF5K3uQhR0acCT
RX2s/uaZ4CxCDeeuPhqnK5r6nEqB6P4wCGaXIZzcgEijl64kOGRDdLmwuayx
2O2mrg1VXfZLM3sBhU3cBUI3FT88zZ53QDsPH1CCFNHZ16o4BzM++Yrphm5D
uueDtQu0jsHU6lQ9UMTEz7hEAPeyINJZQYtwgrfuB4g8ah7f4UuZWppMCk8M
kxq7YPkQI8tXnz2abxGdgCi4fV746b7hNNJeZb6Ze6aPtMQfy+QATgR+CyIq
GBrVf3V2T6pcRzyQtvl2drsaMaWwM+cdTincjmqAYWmx2nerhATDAHGoAJew
3rGe2eotz3/2ZFDYTuj+iTIaE+gi/uydQSOmaSj+/qTffoJbza4zMe9ZMOoV
5zXOg8LZKE4LVoKJirySeUcbhYs8SLBJgiEjcSax01I/aHDzmhHVhvkLVAVQ
x3dsG03xsE0QW3U46boKs5LJAc+F9SOayhAlyWdAZkbmWdTXPfmuRequpeGZ
QyaZs383BwRLJr1bUYwy3oXvnArLVl/zhnpfRd0n1fwrebC3MEik2s0lRjAP
oFBQZHrVRybcd5YbIdoviZ7VKdt/CHzjxfwwjLG+/RfboCjajJlSUcUAPC4p
8zf7puDJ9yPJh5/YWeFjHayPY3qFp+i6Tz+nwBzpNqHlWPvrGspAr/JzKL7J
BRQ+w4VcMPyhmPZ9TK3gntzHTzbrrEpttLRgAaC6YUfJ/3xvZeRLyib3fpRy
QBopnA7hKeuANYdm42k5YzZAsycHrijW0oXUS2JPzaBv92h1vkJm3jBayGvL
bsG4uP3D8tOj9kmcvd1ljnpv/ga3oZePUyw2+51n2kVWamNmOy2ZQlpXK0PX
RrgYuxKPWWCaLZ57YRRqOGT5yMzOG2T6MbibvCPLlms+tVB4mUi8K7JRQuB7
AsmRwRt0CoXITi7lYyYcrjBal9z7p4aYFOSalCztJ2aJJBdLDm+SyKY2+bGV
96f00wB7Dx9PwRExu62tFvX4LpQ8+yDRono7gWKuuYi6efeB3PV/Fn/vddZJ
3mK30xUGTySZXyggr4S6HeakUyKRvyZROma6uRJ1rcP/xZyTEiDOHCHxPFtT
r5hRB1eVpl9srszW835hnKC48jXvoB8c6xf5d0/2rspkAfN4VDHJ4DLFqzK6
wyYIWClLBFXv2l4Z0XwwumaOuu9D0CgM4pA2X8S9gwTO/jP6gre8x0ljeSKh
OPVLF3qPv64zB1j7sIjVuYquLMfJNlpqBEIZGRRf9w7dE7Hmn2h8spY3Ti/D
B83Zq5weeFIUOHvOsaWn5SXkC96JJr9jeGflop9avZHZs7mSDRO5QEIvh5VO
jAr+FpB+EybKhMFYLUB9zhXuB+PzK0jDBzsDsVu8kS90ckwHuIblJraw9ze/
h4EqJW5yExCOQMao3HjTlIPEB1wcwZRDBLQuiTW0sxUBFV6g9mVjlbff6IZ1
shG+Ms6YUwqqbfjAaFExkap3w8qab7fXeLKq6EgnJsJ7S6uqNhCHWzDymrlu
d2AbfJPJs2Z6L/tRqHv/UrJtSdnAxc2UIYlqOh8Up3UQS5VQXlgyB8omzQTu
MZN+3hyR8k+5tmglvCZO7aaYKkx9Cy4+ODG6msbNsgNQSqr1TMAmDeXvp7gy
m5Q9DAlzCARkFyLre0uaDjgfXGRuHt9mr7ReUvN9iM2kgNe0PJ1NhDPWTHUR
PwV5b+r0Llbg8XdvsrMEaWFyvc6lilsksEURNXP4GyEZUDtJ1Su54yeUDyBv
vqLNie9k0n1ybzuWF/IwWNYDGXGIerSotuMIWYav1KLxR0DIsRgjY0OUSprc
WeJB+S9ys+zzD9hW7tJ25d343U7foZj7x8QXgzjHCb27zOgkVaVhMBXDTOAt
9ZVNxnL7Efv3LVVwcTEeAt8W+2b/dcBV81N1iuCZ35LMhE/iU+Zp5Xk+YKF4
aCuQiQm7Whh3nZ0nIcdkXaf038UkvAi0YY6e3Ri8POf1/KAeSmxTUx6dhe2T
KTqm5Y7PRupV37Bl8qWHXYg6SkgLtvVit0Jb1JVEFvQIh/hZQ64Pbt8NBbLV
IdqDzKt7uabQigRawjbADqkf+Y8MJoedKjDTSFQiQhDMoy4r1a2BX1cWki72
CUm7r34ZbeKM6agDZrmNEu+uo23oc+rXQOEvOUci5G4iwybYGlwkTqrmB/VA
U9V9YOqnt+/yBHKZ9XhmeodjZ0+DHYOQHwGZwp+q+YI8S+zMe3yE8q927Rf2
Jr/doQRkDNEZt/0q4a6EyAVSPmiw0wKKaam/sJDZ7FG4Ij132ZadOpT/rkqi
emyX8fRqDXtcCdH7sBel26yT1/56RD6MWZBR3AcbQEglFll68bNiaerbRTPb
wLwrRfhG1YuviGFMI7LkClmWnOahHPw+D/f8RbyaOwMhK5bK6FG12zSU8QbR
a/BY8QjSImn56s7azXC5vQSw0/Isf4/Uzoz6ynp/kFa+m2hHHcwMR9e+jttl
xNZQ+43/cMqlnaSpVXhfy0FN8ZiVri9TnoJ1J01lh7AxnLJfV47Xt+f+ECfD
+jP2KZaiAlqIdehgJna2cfK8qlO+2NBrwh2KnuPiY9AE/v+H9mE2K/iuZcsu
7wcUeiAG+3JBdsftpEQKbYsODGY54u7LpGACS5c8bK4tYTZttFj7WSy194ww
XaJCswjKidIEExQLZCmn23fGlbCsuEeG6DxIRae+PyvC9hXpBIYA5TdqpVJF
/KMgaTjc+mUpWzg1PljqrbIjXjoAjiqvO/ZXbsIKdQb0KQ97ETpqVZ3mTGlo
aoSqaE9qp2q41dLX+iTPag9UrbFEKqrma+CYpy5YLi/7RBX8ZForM5VDGOYm
nFxzvH+tB1CTHhLqGMYp15Eyn5fkqou11CEHSwsngzGxihZUin7W3xBIGN25
w8khBV+JO9GcmeCoIyFKAJLbHcDXZdT8nkaaUSfXM9qqf1La8lxfl09rWYt7
bPVmGayh6IjMVuxQXvLnE3+LfX8XE67ERaQyebKpvywe2lEFBGnfMOdl2osj
dUjg9koUeP1ggQj4RIg7YCDNy3VO9yUR+5WMoyLF1Zdv+La2jOZjxRvHsFoU
Ylx78EqDWZVvtpRNnh5LGGF9eMVLE2ZtNLtHltZ0HPfM7eQi2s2YPNz+W4LO
vRYVTvW/adHqB9e19cJva8I9awKarH7YCoPXms7DMSm9oTHaVlRhB0Knpx/v
rI5HRqpLtjCb3rmoFOCw05uJdEqI37Js5MdM9grr2Y2j8U/Xad1z/4PlJhCT
ZPQkgmbkCeZV3f0m2o3DuihSiAOuejJpl8BhbuOLf5zwyCAGlsScw10tc1uP
vP6hztvPmhH7u6ZRvqCaMDKlieyvU3B0QepPwWrHuWIuE9MnXnixpP1hqvuV
eV8aDGU2aEVJSCGOD2ftluqfLD3PF3R0LyM3IJ5Xpfrog4q4S+iNtDEwRhUv
7zCF5i2IMh1XJEC/3rggiCyulWBQgZ5IZ7q/0ZBPV8VrVbNxucTPSbBAXMql
qP4FliZjr3Le8M9MJpQQFlbWnap7xHCwNrmqYD3cJpEUEit/kiCh8ljMpe7t
RmkJgMGR4hYmD6ZqDz7eNFd3kyKydi+bmOXleGVbd0wzCFIoEvktqMxcOvVK
X3uhaEKzSfd9LVtDCPdBaGMoVPy9MxgVXsjmCpbyKmF5eGn+4XLqcAQ1ipL6
zhk+vds26FNbJ6DtVLP2ZsO0Yp7beb9cXZZMPeq4Lfv58SwYpj1zQYtVBFnn
Np+EPztyTMcvZmjiIQNJxIEyb9E1FFMRdDQdHcB+mfexHDIdy7Wee7km9nEt
P2TrdPzi0l4cjEl5kRL0kMLkww7wBMiSuuCLxiFvO/jPvMQDmxqyovX3zxye
UzIqHg44CWnrCK2QNBJHCl7JehF2f3YdhhyV1Sytwlg7sruF1M8//KtxFa0e
d8yy+nPQSLQkmands8WssNR6eQUR+gtix4nV39IbZ7DUcH2n7z78OvY8b4k6
Gyqc0ZltzMYS5+FU2ra5ZPxiL4IiffYZSKMZSvqSq2ymraA6ZPy8IcYFtCxG
7wpHKpqqids2wEmi188L2l+jszrVlJv0ILhIoGsxNY4BVEaqmAqZGP5PLHx+
Fc5gPJM/KIZM1qzMbeCcszxq0S4fV61Pl07HOuMHR5nF+5ddxfsp9Ede2EXd
l5V3TQoWgeRQnt9999ktqKT0swLy2+Dn+7Z+TQC2Ux5MgVzEhP4bboQyA3NN
mq9qKn3R5WDhQinAdRRfdOdvjocFZH2wu+YkSNbonrGAY5wUs5xywhiqMXVA
RL736hf0B1mJh+GLv5kh7jzmuucvDTaRGIqKwZDnvbJ3vG1vvgrvRn+gxIzq
XiLOpgxbxRvaQNN2gJTW6Mn7bwp/s/yRynB0SZkV7zDYKVhH0R2w1RB+rZtI
ZH8GL+buUJwuXRnEEDTuvHRcaX7fdBjXx5M2Dta8bUszdyMIXQWTmK7x4opa
QZ+8n9HslD/rS4BfIwgNOTc/xg4YXv5/ukETTI8BzCBKcGniCub1MBvhe45Y
ygD7DTLc4+7pGzLWb5o5cPFmLWG4u411w/r4saMNIp9cgRVJ/aKCCDBDgTK9
8TthEvHUYx173h5ByJlJTo2hOsygMeso5VkMefvBP6YlQFsDw4XbuyiaGEQt
0YTgDEYQX4pzx4xPR1pxsPPPxQY+MdgsxHdk2D2feTmjGjZmenjmpxUlGDb4
2Sg9297C/CQfWfoR8xHQSp/esOLZ11kL4uIgSRWOgiaZNtanliW0PElWp9jz
nqm+wjd8Xvio/JqEfL2X1ZbDCFpLuM4MKUO85VM3YkrABeNl33Se27phl6YL
HRTxUOR6aAct+8V73xcRRumftDd58b3yVkL+X7gxKB1jgmmlbkzsVz4RvhD3
TVvkjtYvi2FztSjcKfqsG3Xh9gYz1+tv+KSZB6KK2tT1x18QUro6apO7AeXA
3jU1VrkXkozBApdEkO0wFnjyECCzIS/Iad0uM6jyp0VNf8D4BBNiuZqh/dyd
M+1l7FiTCVwgQDeacYMBeslg5Bpw1Hig2JbY+ORpA6ogBrNwOyq56yszxi+w
QdAVoAOH1fGx4D/vAtqL886so6XeLjDB3xAjH/AVTopcS1gMuW8bq65BFLGJ
SgyN+mivBc1kgY0LI0QZ9UaZ9kXZYHvCKC+F0YKqWkUFOMkjuCYPD5uptEdP
4EaqnOfsQTcc6EIat4jEJRpAbZ03qcV5DxGSOqyqoxuCX1Nfg706G6LkrjUW
sxbLzXyLnYVibKsHMSse7h7Ih18yTQJkTg9A/cdSXWjlTMLhrG1i3IuIxJJM
JoHzUlbdWZhfOo7F5avadvDxp/6PIjzQQUi51jPjQQa2Qi/go9AoqquRooHs
/f7bWXtZEpZqQNykBxaksOa0TGGZTnED9FHeIoKDxznxaguAz9dhEDyP5CkA
Z353d74I5VuhpCWGZYiUpoFgS184xeXe54FoT+iHtr4xDd4rbn9V+T4brjgA
5bk0f8BanpDtk1vegcLFXU+kVcg+PQDFqdzAsI1PDtvnSRSVxLp93jnz647y
NcP/7McWZbzj9LOSBHizILff1OA/4WOEoyHqf1IMJ0ATzrVPNE01kxPL5saI
Ukby9cVL6Q+4JxUHOVLyTiv9/nWpg+wXiqk0bxFfdFDa1Spnj0/SHjra83jE
tUNBT/33zfc14hB8W899i8VbdACHXgyzxV8+WP0W1hCz4mm+RH8xwf/GCe2n
AW32yYEoxKBlpV20V96+V8Z7nwk4sNgoiOzWaHey6o+RpgPsv/jtiM22tawx
e9oTJ7lqAl9mHecJKE9AQhRBjKnOfIIVhK+m225sdlGYKfL6FOO6O7WAcplr
0TGOEm8TTil1Fj7K+JVSF3XOXiotaBSQvkk66CxzxuBdgBQt80TJfYc2b+IN
MyNwBnG18ZSF49Jp5EPUnrT0JLfydQ8aK8Iqg2LQFLrLnPCQH3cptDOjaNaW
yCRBgTSw64VxPm1Dd0i6FydV6XqzbXjVTeaVjZML/ym3KVig5Lfrd18xSgNY
HMsTowwWYzWXRA5/J9pg7sdyePOsvnBqGMqHv0kSYmiDmJNf4iO+NsI1IYD0
nzBGJaXxrfVbhjdSUOMAgoyZgkgqfHBfd8CHtTyec4iuBHQVkEq6cLtwyvhx
cOcpj25Ew5VmpjvvHW6goPvr6LUWYT3EFYL3ak7gy7hxpBCA7/lATRmwcFzp
+dJIJ0wYKZLXxZAOhPlxJzGZ9DVKEShssIfdJhzwNUoue+yVKJ6H2ui/tz+H
HNnuornsAmGV4X7CI50gr7fo+nKngEu4I78+Z2wOzbiSLv0uD/EUSwxZQOlV
xgAqyd563SImJALuT6deqArC0Qg4g6H/DUNpxUS1irGHa2OWGr4RSAPStA75
Yq/RctGBr6SvUNerg8mcE5Tr4pRhmGiwd4s1ymAgz0C/79MUl25jb2OrGEDr
sNE1hdWuYObneza71YmcB7Jbo7+i5Jw/N5A6bNXPxhFTfcgNk8h5pasClwzm
1bu/3cD1FcEVtipfGV2tkyasbmVIXHj2aR3WpJ+Pt/jtXwJoSnPOTLGnPClF
9vLKCbzqYzn6JBQ+JT2UjlfgO86kEdwo1zeTL0XsgJKJiSyupIWInBbPQ5OD
OYPHbXXBOZvUwXZ++P4mIY4gOJdz5h05YRR11ohbS3CfWorTmAI0y7iGNBZN
zg+HNxIb+2+Uys2DDci+IKZVJP6njRuuMnb6xuf7oPYg+rzK6jULqUhR0eJY
IQ+SVEiZ7fOF5snt4hm3lsvuexOkNwQwFXrbQJTrvUkKEPVe0LCILkS1iJ92
RjiVVM/eMM4hi2m5+n/O6uBuZwQp1cLhEg/lZhK1n7jkdOkxSeH/unlNitvy
ecm4LXOWpJeYUrfTLiBsHHnmlU+GwJaNDJYK7C1y6U/VhKMPDwwRW1G9O10m
KlfPomnx7N6h7kpKnWDXit1d5OMryn8Hw2U9W5XVA5YLv0W+/e10Wckwvmbc
tg5nUfgWI0wU41+B7FwjYxxc8wBxnW4EJIpaSqSwYeLnTf40VfCzVe//Aj7J
98YACASyUMF9OaYlVeFalo/GaCwtm5lcyXe6uSkA7NbI4xcUSrwMA02jEpac
EuAgawIV2KnbpRhpIesMBKSzoMRY7ly7+veqfaHCxLhtgxX91O4SeKE5nI5n
zzPAFDbrEvp6pwkGe/LNM6deWvCEPYj4QTsblAPhUhLuasUeYXGzn7xHGZwH
4ZiFULjc2G8cuw9foi96pmYd1lTJCzMISgMi8JVE2DhQ9rRrJjK+SVsb4xhh
B31W4wkuaXVVTPRVV4g74NgVkZRdTkOdCi8BxZtmrOfZRco7aSmAqdCRQVFI
QGxnTdP25rw3jsIzq1X2JGIHjSky2WG54N+3q2GZl2ShKPFeV1sdL1uky93m
R64DUDaG598wiyL6LLRTPBnA0guuM6LpLkcjGmlxUoyLK8tOHfDXzoFy2zmg
hwCFkWbjK0ZkNARP99a2M5xTbM28u2nIh6/UM1sb4qVZj5kHzb835QDbQiZi
xrqjz5iqtkfr/Be+9MnCmnFSM1O023R5gCoh/S2ASHcz3aiNsUq7D5k/jQ/x
jZL7U3O64MV35KpgbsaZVwpYPs+s3U46q+xhEfKQDt9nSdNqu3eZYK9+nlse
8NDOekcjZyPu7wnNQS7N61u3esUpAYPRQY//nfgPmeB5XIYD8+UxgmmuaJjx
d6OJFABsDVhlrPaSm3vBZ5Q2DsuuZIAKVKP1fxH6Ntm/OGyLLhPTO6NpH1sy
2hiwTXgO6XejfoUsRjqrUAV3texE/uj61uyHOjc1ZL9VdYOGMcVujeSMlj51
2v+dx3LSJoGm7vnPL6q9rTEzR083J/TcwjnJrFEsffdhvUSA7tOiWxwuT49z
4JpZ6LB77PT62D9t3zA+KrpZ9vvQ45m6+K2HIA9hfRMMGJ8CqC2xQpzshj/V
9HJn+6BheR5XsBWqqRvTrIKlM+ZpvoQCbE9EbNCtcUl6T3ya5MCap8aON9Ms
bmEA7frWzLABMVqKEAojqWU7/LHnLbYnPaWChLDciYoLhhLyklk9hVAAmo+Z
eKEN5iPJHtTHRSWDmGZtMuPru4E3t+5dax0cYYBKMlqsZHwt8LU1jQ8cnovU
WUePArECsmBsacbbUJJ4PRK+wyI5UJAH84B2DFVeA+aAkER/e3+eLYKz/e1Y
5bjiUCaXbqaLNtuXN29xGhZmZ7YgUjI0vG/OGAI6ggRbU5OueIUBciM81Ft5
Fcipe74NfHW7wN475X7gBwDHXYu1O3FLyQmWhvTB9L3DVrf4IHhykWTKRcAu
N9XyMFM/WA/Jms9lUp+ib1jHAOlLORKkdKXoDM3bFT5FCiWmRKeJhpMzWMta
d8rn5m1HbSTgJvKo46tOIa9F2fRX747UsE6ZAi303qK7Xl9H6VVaFJqBjxnu
cwhlGS3HQUYllyEfMnm8HbWFHlAiVSaGdJiRnbJk+lemd4EMi6mpW9DXaczC
b+JSvTvZ8/4RjLNCtmrmwWdJYBdO716qBKdILHrATX/Pi6DYw6+btXQhJRI7
bOWVBpmeTxQamn4QvR+/k/0PaV7/oVeJ+5ZNGwaw2XBoFM+Q+ltsSa0ZBqdJ
kl7wdjBqIrw3iZnX+6rRxIgmX2613twePT4hjt/1mf8HwL/7udovs7XaXBQC
ZsRWeKH7Gjsff5oBpt5k4h7TUvxRH8DoXLscCBH53CAPsX3G2zZkS1YsR+ZV
alSsOn2zHqDJZ9azyc3oTXhfhpw7IjaL29lO5hW5kVYfYVR2oBu00I/8APkX
dCmfNObjruppHgUDVIkKgKMdBrwR/5mbslN9RCSbAHJ7b1VYlKoNXGi+Dm6s
GxP2DHyZsbWookynX6f3jTDsxp384StxgR4VWlZK5ayG6oDqe9zL40y6m8b3
NWSLwHaAYq154IpbSxxgtB94clLdSOR/155AKX3IeLfv4GsVVZbZXRz2mFlg
kdh4NHS2CSi4Z4/pdliAUb60Ju/cBJmUaxwb6Csud5e4ZJba3+l/pnW5Tmam
8Bt5nw/ghpdK5tK5QZNBAIP+Ap/jBxT3UuxC/ka/I0hxtXcgNvfOJJfir/xv
37EU+JQxa5b28g1UaedZx538nzC7TZ9KK8yckyth+FSrRj+4uMwMVZ2jIKVm
q3fah7Uxy6o0XJjbjYBBlpEuxND6Y+zeorE7ul8ksXH4whJCkCiefiI8IYd8
AXmE0vJi410qWXw5Ll5M6uFcD4HAmfIsNcGVXHOtBo2uvP1FvXXIayrErJ4T
zjwT1Ib2s27DtniO2joA1wfNBgpiNphJqrvnmLrafYqfBkyZxClFatNZEMQi
yUqcKYvAU9TqFtEqAORKJAvkotSOQQjrB6HeLF+cUChXPjqD9duClGdPaoHN
T3JkzxMbTzpaG0A4r2/tQ/ah9CNEYAq7r7DE5IQ38Lz71Xv7lxbqdJzuWQeE
c2S4dcZneDLB8ekBNU6JHipWayXqXdYr+qFLgNB/xKI7qlonbRkc0rugbiBg
pq0DJKhp5k6u/rqeSdwxWZ1XclvZSbhgRRvs5T7LyPQo9u6naUXVDsY4+faD
07OAZ7HI4Gf25J3TBZV01mR6BLl/l0kP4SibQx+EpgLHLUyom61K8xGGvbHj
kGegKbP4wT4ssF6//uE6cqASGaJIt1+5VOWOwUM4AmvoCehWInBlVoyX0bL6
C/2ZUCWogtC82ch4BNfs1LKvM7FK5qIbVvrqQlK+CcCVnV8L3KU7C1w2cZbI
ZyrAyqBM1wJ3kBooJkDQAnSeTNXgO25v3xmP0LA6zjZIkGVz2/6uiBO4uSyf
QnQHS1AKc3Abto8LTcIbi6UjRvK0Q4jKlg+K6d5qxbhe5vR3gCVNMYluIilP
JBEoPgqjIO2c46bH+lFvWYB3rIkEwrBtGDqI0LgHCVj3sY4nHQfoU6N5VD0+
ETobVD/jz7b+AlSSSimOI86nl/tE5Vgb7ed75Sn8iNhMpbd9f/Qc6SpUYrhr
izdgniq26GRGrxBl3gOrLHGJm0HgDHl92Vz65UkZtjJyLNby15AK16zrPTzt
e5piWcDaIxoMwtAlgtjp+r5UnD/OVBlytStoldpp28GPAGwTSzFmaAN3CNYN
lIcczOjwRTgFRWofgrQNd8ml6vyDU5YC+nwVswVsXk1jaJYYJJjL3hiwXJ57
XKR3EPs0yyybYkcNzCYoMNno2KNbgcmV+Am0n0nc3OAGkuosptqPfMVuZSfW
6pjvg51lQNAj6sP9B+UWUBZ2Ty3v1QPBodzDZMX1RaUXjJr1NbQA/KMLAupC
3+Cs08lYx4XN1F1FqyXFTh5ivZNU3j/3zS23BANwmk9M2w4is9/93T9GVqE7
bh4fYuLNIkNE1H3Q0yvFZTadjxpmsspJ3IUKjXdXlLeS/43eZCUwGReOLDY3
ey41ml3UOgn0wZm4fHHrFJyZI0JjXAnRp2Maxmdyf6mhICegVZK+DayekhAJ
Jmpn8kh131h1lXcvNu24ILAv+w7b3OJ1Mc2NnoufOs+3mxlybI3D20tNUqTI
QeCHmijsrK7chDIuvlDM82w03fMRKR5Q3r8jedBeIEnx9K5Azm3fs1gI1ZY0
yTQJ615WLFXAKDweGFf11IjRq03a+pSp7FEZ0CrdGSaCgVGCoAB6GI7986iu
rsLq/TZixN4b68yzEx1m5SWwy3Bfb/BA2S0NSK0ouWIlF6bSDpR9q4DXSoD8
wpH87RgXxkdyLBiSBIR/SBS8+Q1rDKYmS6+kzGfNu2I2vVahmMJldBdU/o/j
TC/DNBm2j1lax9KG9Ag/Xiu587qIDgbBJEI05R+wS82ETLKpKO4N2xKTYZOJ
aXJArJodmawPIAUPgM8wCyj33XAdzHScUZm8TSKHYbAA9wkIDeeGUFE5yTuT
e3Ou6o7+A0zMTo8Ckq49mERhmMVesK7lBIh5ieqLE7Ygf0PKfS0cYeylfHPL
iexysdaSrxv7n5L0LOnNA4rRVSuzd6K/Snk4WkzejV+ubdM+Y8oHIZs7ClnQ
MFrWSxIAr9l604vCfejsvX/SqMjSDkTIWuk82UsVxEmb44TLDl7QKDm0ElBq
d1N5fQPF9JlZpTWlRWPHcIB8lEcBtocAK5N9CuW4Vhz700PKBqZCLzaNmKGL
EOL1b34RSaMwNhmhl1DaWCiqPfAl7nKIxAhj2mRdAedBwPzX3wnHZ6Uj3TPN
LORzo3TWZm5KN2bB1mRxEyNZh/F0zAq4JJLHXiy6SR4p953F2LWFoiaqOugL
izXQHQBFyFX2HJlsOH0xlZlYLvHzsaYVek/tkz7U77+5bUAtVapwDl6B5kIO
wls036uowZWgp1vALyoK2VPVvbUiKcDu4PPIIoA82jR3Pvimh66DLqHAxrvJ
xj/eUtHlLSSl29TVtYsTO5ZjYeiHlZCd4q4EgcKckVrGU4Q2EOJujxwvzovO
vOKGSj5IK92vOV4wWFBsWEXk4wFkgWAhdFagOcSCI8xG1jtPA/LRq/Xi5mC9
taBVW9aNEyoyoWZsE8mSSoNZMrbvLXM6fQpG1eV4WkwZkY0i4baVuJnb358a
8IK6BTjROaQ7gcWZH+2fr6iWuWLVlXsp1eck6KGiyrxRD9LDR/cYCJuLVY2V
r1Lj1h7zu41RDyRuRJEzpzJwZYY+M2Lm/jTpgBTyhDEkB5xmlmzRSGajEAhg
Au+ag0zIHW4OO+N6OsGWuSKPiLj5DBHxO3cp7o75a7p+on20B9Il+KytLiDm
YIhubYgREtgRvnJ72eHWhA731+XwN/TZ5XH4N3u35DzKdedRQ7O0tBKDtyCI
6jQzsaORKc9s3tf3GhQ4sVaxre/InL7v7zDy8dnxWYGqf7jvw4w8EMK1uMk5
rTaMo4XgHGoo0qF+0JZA9jSpxE6zo6QrjUpyytzcQT2OiXF5NnmqF4PSsJHy
abvsxeO4Tr3ywP8jWe3ekEedQZMp6fmFDkFPlwPDSwRlz51G+NMCHoZXEtTK
ePapg/KUPkMcH0OI2j8jJVK0UH1/BxmlwhfzdJTJ0xSy0hR3HOGbbMRrMknN
+eNkY+ezpAT/ZsMZvrW6qRjvDK8JPi6/8WQxJ0ht7aThX0BdJPALSjYFguVZ
kRFBsmNPiTVKcw8JsWeHWW+T0dnJyRQfkfmBDfWRO7aavuDHZjqcqzAspM84
e6biC4Wddmqrvp6KiphrNi6O7jCi68uEGj9DYx8tbs8Baq2OvvAyldJnK4nb
T88kY3rkqg767MVrBFB6zFmS2MXxUGvgWdiwgtdvGuHMBmEIRZ14OE/A6uLy
4LmLWgWiYnAFpO1KZ8jJHe9OhJVM+WnR45MXh5oFWNzmX4vThtUchamRCC1M
HrWOOZqDrYJGSTfL/b/rOrH/E+Vra+A0qHnrxP9E6mmKes3suKRoSCglZH3c
IrSI1OcmY7M03YxCM0lukEokR97HIgMgFM42QsxZoiQNbClGB3r+ljKe+/Gi
/ka/d4Eod7OTTGhmz+sYi/T63MZrAL3S4kSVX8889y6DJ0yCI4iAMGiTwO1+
wHi3GzBy8SJ07DfjQ0rZuYkSjhUSn0IQ6J5Tctl1Gfkja/2e47bZZa4vZarr
BXikbBuZ9mAWIKxWDyqyQF02LzqC/5NusTwPVvujkSdfDeS6xE0MRiGSFlaL
Kx+5uTeln4OqJlbtd1SLsm+1XeXdxb0HB0TX6lwC1Wi6m3Pns+PuEPnKHPZV
cjr3dpY1Jc14AYoba78PkNdymmWVMzIc37ZFr0DE1Bx2jvNM090NuvOzmUaS
9eHYYVXPBMj/VjgBae6aUW9dN5jfBeD2DJscZ3ZGxrH5jLnhok2uIYUNulUq
1TfdgdqFPXsQInwg6ag/QNnnR24QkfSmLpmfySybq9yDV/gZiRROirBFJDTu
IzHeu4on33S8UZP0BlKDvgmPVhsESxkzU6LoPkiJE/JM86qtnzD+hpWM/ZCN
B1iXDMRVK6YJSWLtGtWL0iewniQY4Zvgg9ZKKvSIXmPAXH9TmmttcBrS1vV4
Ak9nZW7O+wrfVIDlpdp+Lk59uPdJ8sP/sndamC/8CVhkdzCeljnlLTQfgaz4
EI/EED2a3ab9lGx2JLKBTGwH8o4G5d0c4tgO3E+OmH/dR64gw73c4wIUquLD
QbGGPt5M6Qt+WEt3/2gx+2RQzoYYAtrWReHCB2R0aL8ZaEWdhSKtq6UmmjhG
2SWXfFm+k4Qfbm6+ciBnjJwTUEzm7UzVs+big+jWNioAKHqr2dmFeDdTfSt8
t6NJvDULu3m6HYl5/B99vgTLR3c3fWGnvhum2140ljrz/ni8uEFAqv/JouTu
JOLOZLLYWPE3bKcErH2lZUMMWy+2lSsmfdHYBosPI59JkbuHUMo2iAD/IzWy
pl2zO4SjCqj23Z1oTT8NPaup+eS3Z1UjczvFXYUKuDciQppEDpMF1FQ4FIY/
fH0c7fWR5DTrphXWzuh0dKvE5NuhIk08IcMbFspTs5PcSqC4xdZKCfrnqooD
PD4NdICfiCbXibFdOWXEBjISnCqo5bjPAZAd9tYf1cMKCjBHlG475Xb3bpF9
aj4AbJ8HtodxVRn7GvEPEQQz3cx5B2b79JWWCk2Jz/g75XACnNhDzMSXCqOb
8E3WLa6DSuRLbrkqR8AJtiE+9rYlARchN5M3AHFEzkY8z4tIzfLEkmQfosnk
pSq271aE0PHK31zqGdp5CBnlUkWEZNF4kDYmHBXuKd/CxniQpk4EqY0/wYRf
8ytpYNdK042UKoqqXsj/YM6+a3vDepjHQ3tuOQIglZP2d2wEGVUdanQuN7yz
uE10wVVUQ3k5G7WvSRnClBjnQlsOCJGV9jdRhuRCT18U6YVde4EVOCO1rEBl
Hz7m895KdQHiMMhT3o8/H98FXu3rIQcdS7OvPKIHG+H6uiPi+PTdD8xXTAFu
wfb+YwMYrFdq/DgTHeS9jU9k1xRMPN48U8kkBDILlnTBUsMRgMBJnZodT/Rr
skAkyIzH0BtyNdIbXEv3A21U0IF5LHAE6urALcdevUHX9EIv36rUDxQvdrkt
7SeCnUv4cJSLxr7BkCJpH8y1hYWkLiq7IUhjc7HbbtnG/RBBh5G5NMaJDYcV
QT+zVVCnJ6Hvmmc+0nxEwfNURqMcsxy5p6lyoStOwUNxnDO920at41km6Tu9
bhbtGgbtoyKWmzc74qVZsW4dZ6KFdRvOPpT1hz6eqpIEMXPhiISiiuZUIoAI
Z0AuEJ97PxeEG7Odq+iVa+gCdMg4dydiT3HjSvVD9hHjLp3hAM8M7pSTL3mQ
IV1wI9X2LlxapAyb3yfVWwRteqIDX4xvRW9UYszGLKUHp74CCPTJ4pv6yojq
bXJsHca3IRhZFUsD2vF8XD7OBCAzKZKe8F44DCpvPibS6Fyrl3jEGst1OPOC
v84VMB1Wr85gOm6MWgH08Ca8chAgrJ40zEI8cxhCiiOyAKGUlm0AwafxLu+K
NFHWbhU66GfZJm1e9bQCTWKSoErbMUSsqGxRJzXX3N24zjMouA37zadSLIKw
m/7nvnDrR+axeX8LD/XKP7fMd6E3D8SYoXorRJ6ve964a9ngzQ98keYUTbX/
ot/oZ8O6d5iAgLu4x5XYXz4tdSSSMcq07ScdOrrt1jOClkbMwUpNoeGkojcw
nyE0AI2xoDP/BNbeVAwWiiwAgVjmpmZWkIZmG+2DMOLf+uQ62rQdekeVm3gc
HTgHs1GWFWYnQ+O/bTzGcTKE8LzPOuGSkNAz8+rT8CrW3y0V4Tsqx0qx7ndF
AC7cG6fKGxvPsY2/JNUdQxWdK1tahn8Ghaw9p1nI++pEx/NKIpPbvJGAvD5U
E2Gi7+/7aHYuaP8bJD84XdFjNJ295GiJayRMf9NwdSafZQPF9uCckeIo4+Oo
F/NsdLSIHotQRVCiltV6JbPOljP2CC/4dHmcOSgdN96UF4s1Y615A5TbeM6p
3TE9A6bT4AK5jyb0biIwsDtDy/ft2nPbdCNmxrl9z/LmtQF62IqJ/QIL1/Id
JG82V5IdMOT9+TTqyHg8XCh3TsrgRA6yxu4ZtVIv7a7x5CUlGayNDtTQ5Twz
8G9tzUnOEJs0K9xWRfqpyUqc4mJe2Xc1zSFBTeCekk6sgYlZWK9W7qsHGT7o
nY9ZhJGADzR+fBCBaUWU38VcpldQrTN80p/RVuVD3Z3o6WHDZUQm+zhLc0YM
364OiZpl+Zsyy+rXYCWUzEIDlESUE+V9WA4/6U2BWAQC+FNaJUvGyxke60MJ
WVbUDBW7RkpJYdN/wK04jBRQ6MOzTr0HK0w/7Z6Qbdmkm+iPwStXpqMjr/pd
GVCv+g4czgVuwTTMg5I+YHzIieluoumDFm+E2cj00Rtmk/+kL0cyPUa8MnCs
ptQ36f69M277nSB/zLsQR5R8dI7fbOX/rHbgRj6PyBkv/X6ayfWqmYiGxOWs
3KF4Pj1P7U7L1tdTymU4XvOr/Jzbve7y7CNgQbI1LD0eWSFE8VIdldiZdpte
RGRkKDZWOOPlWnTbUpRf1HyawdhvFv2+AOXm7IqWyKU0itwoLpHmVQGr4Jpy
626xPSuzmuPBerZxx8rsOtpZdGw8ZLpxQZiCLU5lhFDEPH7LOVDoN6zUZ5an
UxaGk0WsiCtjSnAIpH6AmkTtTV+aDx89lQjfCdbfB9PvQJnXEjAgC6U0wZ/V
uVhBqM3/uF2PQ4SD0aUzvfDeqfKmuePImAsfsL1I6NpajUvCossAb8R7zWBA
SuQVDI52x2OJQjKHk5+W+BzKQMdg5ink5gzBW6zc/1UU/TU9MuiuHFV3mXB/
XTt7bLMI/xryTCROW7brAuks8vZO1VOPGYkI+SojBGKt++dJcCqWjgoIn/4w
txcHi6tAlbYCMaNcTf9/1+4n89rTFZG7hNhhNIFB3SdKTSwLbzMQDpynfoVp
tx0nxjTCdI/ab9LYX97+BZJIc/cEuJBKI8dwqQWEYUO3Ko28U2sdKfOqtOUk
YsOR14oo+0hVxqDM8ow0mj6aLSH77CUl/IH/o/u5jOIvKzH9TWDIbnVYXbBj
9RRwHrjM8sGjpAKMcG3NuPMUT8rSFspqdTkore0JGYvIQWp6V0uRchUwfaNE
TFQLILxVdSlQi7vcHGJHwPhiiPYQ8iFAPU490I2HcabKsSZpn9hubXF7h3JW
GiolSiAUK5vhIpNzMyl9fu4MidKp+RdE/shfnz+O4raUg1X8tsxmxwn6MgOl
HWDeh5vVgxVoT849CiJlytrW3gzknew/DUTonBI/Asl4jad/f3gkx3WOuuPw
0Q8C+IsJe+D8PDmDps7vFzyTFhnN2sUIJEOJBg/5rW4czx+Inc4HAsBq755P
/WpWplA3fX38HHYnEMzkiQHoeecALmsVhaZN3CzGCWefqKiKIIJV7ATlRaeB
SmrqG2umtCopn46Bd/J0O9dptnhU9wmCZFm8xYF2KGtRU37RvgRIZXRXzUbh
1SS0ybBamAuqXFSTSIlL7m/gY3kce770AH7OdRhgx+5rfTc+jtyHS6v2ciy5
pPE9lfV3BRAmyTdrUTWHNSJkx+DU7yTQvV5ZDvgbojvp5vnpxvlKzX7iy4wv
WOxZBOwcIjsqoYubioK2fsGD5ADQpGG7sq/6GexWkz1S3zxIbUjiU9qvcPHQ
ePrNQ+/t+5s5G1b/rImXGWaGBSeVjusMVfgKxQeZnBwXFd04PNGr2N1Go915
qp3IC728z1DpzEqTLMq83ZyJutdWzo/7JfUZAIbA3rtdwT7egnWFlMy2gEPi
FokbVvHTV6OpDQyQFEFnfk2LjFvlm04XHBseBykSpLNZilDDFQIXtWrphyCZ
l0DnJ/N5nwhsNhJvBBzQLYoISqel3LNalVyhgM+EuzeqlMavSZzrYwg7j4Z5
Fyep+tRNeSOE0t+xoT7gWNKGE4V/tVH6Tg7m6ufa8AMSSwMYXTqxJ3qzu5NQ
uC6PUOaKRDVY6C4tLUL2pRiYnp85UUvxTICNYRLNNSwtEMrBfmQTSv7oNPL4
PlTt4BbPLt98v0Je19VkzOx0XuhD78YY1g9aVCRYKcvnMQ29cVtgWb+TPQ09
6oCPBEEyF5cu5AXOGhX5M2ruIiXoNV8HmWUgLK8xtPCPclWuaWtSMAmyWcTr
5gVsuhOfm8Ag4m4RQvPnCkUjbDPV7w130blZTWwu83P3dz9NvcS6TA0S72fh
cZHnCfM9Xy2Jz28BXyDxe8uGs1LxxdskiJMy06Ugt9ZDDWTMLHI+0pgG1alC
GZ66GQVx35F3LJya7Hj2Ts1/kN02Q/2RoQMqT+W/bk7Y8+2DA1pgrStDM03o
RLJJaW0QJM7GerdoBN+4xpyhTrZz+gekP3WQJH5l0rOVanXQ2y1MRMTNqeLy
9zKLzbsiqrn7nNbuxQMxxiDdmTSQ83Dwr7JYj48ECOxvdZ9lhxcnadVxZdK1
QQEGlXLTIkjXKE9jIwGEzGID8JB4+v/TY1vH0V3tUHHqysHeX3AeSri9XqUu
5gkBflFhsobiXIiyfYMTW8CZt7MEHwsUuRnqRkyoFVQSh/qLS+EUv/X2+l+Y
6alK2VjZmOXdKUIzr0INzSc3D8SEUcYfg/znyDKVb7tUsqSU3qwEykaMusYh
5UtFDLTqAPanLKf+a4c5UW8W1XJNtCgLE2youG6NxRz1oT2YqBiiaQPZtGgV
uZr50ATWfe20/mLTPM0BNxlns+tmbHMOjZzpKrhyhBv8+OOc+dwGwHmKH/rz
FkkC1gp6TrgsyENy4Nl8cbCK8IHpleW/DGoSyyIVT1hbae74HJiUlFJA5rYj
m3/aPzC7VeZq6ljUpG/QGYeH5Cl2rrj1UwN9v4onnZZaid3wgfO5YN8iViu8
1WSqBaY2zD8+/3D1KGLHCR0Uyz5CcTkhKFyPayykCpmlKlUIvNjL6WK6MYai
9n1xhmWaYD+XrDmqgOxhZZMjjbOLboL8EbrLgvYLXNq4EX4Kz/IauYtJmt86
OWAUdecsTHYHrPB8rWXqT+jaE+bMvLOr2COUX5s77dGPKIgsLJHEDewyckzl
pGFerqGPVTtn/LfzttfWmW6GMQxrhKsoosimFzECrkHC2cdttfSawYc5FyYK
DmB3AzEPUjmEiIEfuMN/JWDZtdl1EoBZiYJtsv8ve6zU4Xj4WAdfzJwE42Cu
pNZLzao6l2fOWGJM8pdlnIXDRohkv80m62WWiGLOW6p1ZmBiTGO5cExErED/
UNbtMEMGTDsNAEsLazcWru3Ya0D7iTImc5XCzypQqN2AhYPeLH1+hpL5AHHW
ssdXFZEY7qjYdLdepTHmCRBe8simVqEzThQnJstZnrszHXAsxcxdNg9zohia
0xbVzBRsbUSD8eLT8W01mGBORVt+KDjb3S9oxrq05WB2JOKiLnit+arraw6B
c549gp3gT38DQH4SqpSffD7n+5C+3haokp7CQjOwYtmjmqzcTdu+ibzzDz37
O0j4rj+GH2Zs/pUWk6gHDaO64XQBoTqNhggzKcnA9qsGEBgEozsUZIoMTql4
xfTKvqGG/oje1qS5L6XpMsyHf1M6E8ctNZC1AQg8nF9ba6r7MLQk6av55mpi
yUE8RI2AxRllVyuU1+7EGcA0Y5mba4NMAIumIH9L1cVYMnh0GzX7b+RxiVSW
VYCJT0xmtDrZV67Z0mqoGvPpL/4u3ZK/R48fDcP9VfQVC8UsIFgEX4iqyWUH
6ciBn70TG83yZn8wDr1Q0Ppr3SIw48Kx3Zn+zb8SKUAQWdjTsNELaYHDVjmz
T9vg99P2jrfqWSTFIEqcqj4rzHtAbb8wVW9QEUpXhS/tXOnvJ//OQHTnGfY+
2fjqI3pt+6rhlHjhLs+JTW4MgnaaE3rrFFhGdYAxTcCz7NU9qZo+nSuPugYZ
8tJscyyCk1MnCsh1oz9t5MmHwtTWbUjdclmBBL3m0S9WY/+vHB29LEMjzohX
tTdhNx1nm6HmUuvaBVVXCNd32YwpLcn7ZwhnuoJF1bJaQFex36VaPNYPmkDp
n9puh8498qQjxK9zzy8jGA+tP6WKa4jizFvGkXFc6QC74SiehwVqClCo5dIB
/gHCoU83vugJ4RVUI+COlkjOBIeExr8R7PXpQh5nFle0Lz4gAhqpq9unRUL6
VdRmnjWdGlpxHkZYxdeypVsg/Zg0J+obtp6nNnDRjJmI5QfVYnM2uI+QknrD
i0/v7LSp5DKpmPkIhy4Te6Kz2EVaSPS92gKDNPMnIQ6xNsqWS4V0/nleA5oZ
+f/nbboQm0hIRlcHHuZzpma7QBi9bleULroHOMCZLvavcwDnLmt9qLNOkm20
8Z/kAiBPJ/GoQhYP1/vXA7Wsv1mH80Ixo5IhUd98uQCnZfyPWkW1+6vdOXAV
XUyos6bEp6SyUOonTr81IGZWlYGtEST0bYfv3lk8Uyn/3EhHv2AJyiXJuDZD
oyVMtHZeyMnoUJriVEGNm+Gbe809vwbh/mfjLbuuw4JiCE82HNbVGNwBm0UF
suWH4m0T2f0hI6VzaM1BI6mfWZhp+EqRaUwOr6LR+EQoyFrG+dOB/4I+XTKZ
nTLJs3X4g54bzWaKN8/gyVqIEPQDvrNZ9l0SvaNgb+6F2I20mLr+Bxc4azuO
vXAP3V6NoBMuZzl3c5cLUV7GtA6cJUSxIll8VTPdOYyItdSg4wOIdDTj+EvB
SVbudMALMVxL/6wCH7vCBwF21TheyK/ZlLYDKvQMs04e2climB0yOWrY9LU7
fKm9Up4+5SeGW8PAs7yrmZa2NC/IyVSEmZZ+zd4NxegR2RZpIaxX2sToQs3w
s2m6O9np9X8WRcrg6LtZ1DMdsg+xLhu1Uh5oc73QDo/GfpSUfCum/l/ZoH0q
+d/w73lRlnlfayHwD3WWeYfQemrtaO5PI+VlpS00HmGXg7HxdhpPvakuNw1U
i+f0bCfUdQsaQQMiZ1yoVlGx0X0XdWy9RuAjphT7DvpwuRrpfymI6aGK8t9p
xiG0QKcJkiFM1370oOvJogZs7uSVZUyGVaB0ZBC2kIklnV/nJuf/LL0F32vX
Zcav8ZidvfAETCXHZUbxQk1iOodObxdeR6Q91s0zhX1gsGKBZ6BgaHfqPrGT
0b50u0StTMQ5nrtNYubuxXrl24TDbKdpc2uDyw4vQx4vda6iKrtZVcoLWGC6
/9+5iD5Q3gaXz/8S4A8/iXMiSiOY8vs9cSejSlWtp3KoTOi9Kjs9ZLNx02q7
4EcL0YJAh5mTg6cteQpIqgbmONDDMV0+LPn+ZSNnlzSQ9BcoDocwczzjZd4Q
CFw3+jS8HHRjYr4AYscU0Uw9EtFKT2ORSQZRh2uhGf3VJKUmTLP+bn0GIuU/
AFajsWF0KjvxrnYa08ADKvfUbah+XCXkebvXzUkbw3OABFFA7HRTfg8G6wFw
e2uMZomdN8+PBwovvV2WEXShFNPQI3cU1tJMm532XGYjZfYZJkAbCuR10yA0
l7urD5bNuy3OAHYdNz34OUni6+XJzbzL2M62ImyOjDUC18YEIgR6e3nuzR4U
VKzuwEBxF70qkI+VVUFjmE3NA5RKce5q8hkzVO4TQKGHFyD9a/wGBhkqsnwt
aeKqLvt1WAqp6tyw3rIdIvYcfa14jPFXP6TzoSBme7b8j4rBgvhBWr2dDQtV
x8V0qEEh9e3CEct0dDyBWrnejJYPyjU1Evi5r68mFdSdpfLjxa5OIHg+5Ehl
0u7Ea1OBtlScBlGQ5qbgPBnDS8y/zqRLhjjlEwGGzENETVnMGeYgA4JtWBdt
/4it+FslmTz3EgU++TcVbHg+nNrYLnTr19J3KkVYyb0z8F7jNu0GpEpvhr5e
9bxpUB+q0KUf2R9RAN6okuwGfEvOR1Ix/63OzTSG3uFPlewMjEGXqAtUkBjz
IyLyo21lC14qFhHHm/izmglgsv39/yOIEHUt20+0oNUejU+D/M7ZFHocpIuZ
f/BGCZ6ohJXt9iAY28Z+Lk/TQh0e7oREjfbjeemuJIaU72hjwrLizQJJd11C
zG4ST9zFNGLNxOdVrGQKAc2XFnQp1yNAzp/+Nm15NLTcZdvAYL3pWj7ZS1Cn
aG2p+dQlCSboHjqeq6tnJp3S8cbWERG/CKMOZ+/h8wSrvwekym0x18myztkn
W/1xxKJvyn6tgixukOQT+OF5KwIsnUmcC2NZyH+QgKYl9qd4W7xl03Ih4yU9
nX7LALp3GPTchCSjFlyGX+/PODxaKvvp0qZxGMTwxHIbJWO6bCIR7R7v7MKT
efmRaed/O7FuJbh9bgaAk33UThCGccDqasjIolxc7CUkFnBGNE8F6Q3lTjv1
fKX2TdLaGmaGZoBHNMswdA7Hg4qzZ4+XuVWJbCUApKv77HjKukcYk2no0EIc
Krx5uhAP+rB5Z8CZWbj3GA4pV+fnXSzfQ/T2Vp3DYJoXX0O0jxWMNSnU5FIi
7xhBMbbFK1Dan/Sd13SDPYdwJO9Zcccgg+7FOBJIJwxIuD7Vk1EHpjnBpqQA
DHFWnrIoV+4d+ldI6UNmJD6+0b0bubkRw/hiVuuToj0TfLod+nDTZ0XEabhL
gDIXe6oPeaHGwWt7LUKCC6vXgvg24VcpeO/EJNBUI13DC8YEScxSn0epKNNA
EeEJzqbd58fa0lkLx4IG+6YW7PCpiRHe39GPRGovpDtswyr0fZKXBCXxEIFK
hP3j06dOaN9HPmP/bkc/o/1KYVemZUpwcnUdHWn6x1rUp1vumPO8D6NKne2Z
+KwAcmdLbAQnRBel2YE7t3smytLWNKe155jJRMiLpu5lyo/UufjFukTp/Ae9
gx9lJ/ky+xVOnqqZ3uk0akkoc9efTNbK3vJnW8XwbeT+WKJ+Sii4XRnYX3jr
4zQO1u5OBkpEAGJw69bTx2wDnDehVSYfXJdY9DcIhIJ84jyOtyMgaGk70VuF
eJ3tYV2WEzRv2YEExD418w+oLSRkk5KpgNl2S/HtgjpVb3sGJh3jdfA0w8o6
rmt8FQxOEvLOxJCK9ZHKRW5aP4SPy3hy9bGn61RxbVeNnyIC7l6VFFyghbK9
P2WvGP8NOGkl75gqmr4mwYb3w0tXfwPhQRfpxUDcFEJ+dXJD5UTsKCd4RAM0
Ey1z47CSMXMDpe56NuGronM0dlDosPb+rL/Rvp9qiG3q7T0mX4DJuDNivybJ
R4AOBY6AP3B8NyT+MXlyXEqi3xQbQtYXzexH77AgWrP2nbNu99EaammC1arl
LC4+5PXOx1BkZnBpZ3J9Q4PTplfnNWxv7RAzonZw05GJWUJSD6NYFxY7Ca26
ka9gm8h9EsAapnCjPjiN8RGnxr+SEQ57dO4Zkl+gVkr/iDNbm3BB3TiegMgJ
5vZuw3CM/UbWTs2YV9v1mZ8cSco8/Y7wbBco2rh1iu8p1VKvLTEUncN6Olpm
slxtToEnaPjLzA2KOWw8CXYgSnPfZKDAtcLBlB0a0VeLHew7SuaMk+j2Hl3u
zuEucwDfODF7dIBzKubML1k2d4oZfqZXBXp/oH05K4x89vA/LMYdncFb3doA
vJaYvkpBm+YV2kMPKl7iTBRURpgm7SZFAQaz9BhtYZXQT5vQKhlMI7DXLcp/
/pDfmtCgjBHYoc8kGC5CSvTAq9JSLhCKmjrnM4Su6jTHPRcn3QqTsv1C84ab
MR606U3fjHQmccfFya3N+ROirPDS/YtknrhhFXQLjciAmqWkShl8hQkE1K0v
mQ91+zwMFeBDmarwYd5LYmWvsEfE3lKzGjtjx0tiURvLeLRbICFkvi2mRtQ4
UgvzfdzkIlrsS3wI5aHy6PQNGy7ZMuAIw/DC6nhbXH11Sw4Y7KTcT/fetHuz
uAHJvKi364aoqRjqOtFg+SGPVy11aCg9oljKsFNKEAHE59lloK+16Pud6Jq6
Uxvlsv9vMciQxu8NvWH6JKZequQcLSoJSG+eL/jKjldkExCAep3PwxsC8sxM
kulqpozZczb+Ni3zHhTfssjMw7GqVwNnGFx1Zt1UCGKM63EpBmP4282y1M2y
s0Cz5m/3SGihIqyBYjWpVENhsDou7w1tmvpRxK4DPuU25EwO2geUxQWCRK2m
adHGxCYB1r56S9j2JGnlh46y1fkpoJ8ldZ8U8SeRyIjt5m+jNOWclzFmAQvd
B7nLgfU8r9j+2zdeFs61X6ByXy+UDfLAJ2Mm2FCgiBzxcooHOB0hfVgtUFnp
QejtoTfukKYNxW9nJ9ROSuaogWo5ZzWoH3Cz/0qZTa4qvtoG8XXm/GTB0ljw
pi9R/4JFba5cBimY3Om5hWgy7X/zMaPqqs4qcRfgxXeZaTQvT3X1XiphFUBt
FXP8Wft7fG+/lflrDheKCjoBJ4QNyFwYLJkmibS+QecJd01a0lXPpHevjlqy
3HnYaInVO3HfgkzXlxFFAm99mceDYZBNaLGD18s1gj7U8l/P22OyppWrvshk
a5d6c9iKPfyP5DksHBhLHU7Kemu/G2MfxHRstcMEShgAZ9v/ZD8l/NRbLjXD
Jyi1FQqn7eEYH1xXLL02FN3j/261tR2XoDHwIak9gVs5GDZ8ZdaF/P1Y/72y
b0HIMI1jWo3DdY9aBwQ+01qwPfH+qiViQBnia3PNgPpTvjdrtWep0U2nHUyL
A/GT4HosM1HOyU6OsnB8FpmcWECh59l+HDHGT27+BNk+tlc6METSrWCaDQBw
Idwq7UdraRBug9/CWrR9XJrcGTZ/fpaV6VQk7YSJT2XaS2UGaWlfTFF4XY5D
5OMDx8oE3tQPiqUIlm5S0iMnefLGYf2Awt9YwKRjfVQHOLGQ2DWDNqS1vb3s
RjVy0MLgVeQU7D99Df7/G/UnY0/GrQIEtbaIDxVGVG18VDP37e9VC9FG1NKc
4LIEGO2zIJUTUSnmcBrM+E0YNDOUyx7qRs5XzVtm7qyCHidRQd8QtbdW87S4
E9vtnvD2CBcI6gnoCa5m98pErprLt7ZJ7S428xTtAQXsNyqIqSwipZ7p3z5k
O9pc0MkZqMF4E6cVb7q21oZK6OJQwvzKcosCSIfo3HbsLnNyAJ7fgPgWfYxZ
MumOk0LMRFklsGU7znl+unCwGRvkTg8vMSmdfUmJHO6RIhgONzCn3yTcWPC7
OF8cHWv+/Eojer2CMO+rcLOQDLsmqVF4NV1VfNTFZwcGFNNwuFwL4CfXG009
Fn7KX1dkX+O9s0GsLnzkyqoyK5PTPpHCqYgzt4OaUITOBD3x+72/mvhq2+72
4LoJIWv/0OfjiaK2vRGqEGg8nDvKyHl/y7z111AxhLQepULk3AiORZpZT2ya
bD+tMqgVJSLG4NuDoj2XVCk822uUOhi+EInDbFrh6jkZvq5HK7IccW8wfubn
JOLTsHZWov9x0L3NB0pvkaFPCz4+WcNaVOMzEZPijz1NCTTEOjn04TDUw3Xf
meEcc6jKgKtyUqnElNW8SohZbHcuP5XPqRIDO4cDevpPajtg5Yw0jitT3x2r
JQRfX/AfPrwXZOF+YrGmYouY3M4CgFBG63ukxz+ZwsaLjxf9IU7ElRslMwfx
NS2S57WmGT7zj7r8tX64raqA/nw0hPz6fE0KNEb+97/LEril5LuwyFhJ+fxb
9DjnaR4H0uYkkHkIHsrSeuz2BQMmczKlhfMYXIC3NkGBK/xS1XFHzsUA7TSZ
Ztcm41GOZmOSMaW11jP1NuWaIcBGv81QnH8xH+WnCnYG9oom4zU1gnvxLS9L
GUWThr88MircmUL1d+oQLTCrDhTtBJLXVRcRmuPeIbDXxU4tlZT+GMNiiKu8
lHx9Btb4UFIp+XkOOgCUGckBDF57reclc7wCMo9R5fsmjCcxddsBSzZk7/aX
KVZtWLvW1a3tll1XMvzr87w6U19lGOUM5eCAMAKBZxjKk38sqm/+83nVQrdp
b2XcCstr8lNV3ak2P4r1tc4IxLjrEFydqL56WoonKQxn84MbqqRyfwWBQOqm
NbToFpFLXih+Y/TY0dmdS6Jihcqkhfy+Oh4KdyrUcPZayyXs+ANELr8L5eko
sigbqmfhxBW88r70oZerJrGpLs00/NEh9Bx+/RsNDDp35c5rY64IQ+2Hb7hL
rjoLRDkMUpuKZw98jRV2Vty+SRrY4S9BgXAtttv8388X2Cy2rp7m43utuqYW
X5IpDe80xBPcS9sgrVFWmxxb7kL5AHuRLnBqRUmVn0GGEEMt8/lBbecr7Im/
6Vp8olVphvBR4kAGgjIiF2LN87zLWP4m7Cz2wJpASKg3K+4LZaDbtTg2X9wX
ZvR2LeEEArI/YFnR8DCUp0JFhdzPBV2v1+yMBDDXF5u4WO4VN6maDvKlC7LC
MnnlyxwmStsNRFG0WAiynWOAQmGlyjjUQ1h2+43+yP7sfb87rjbW4pfdddyo
rO88Z71LDdWFD8Ury83amYnfRDNLq+g8XQxQx+q6tnY7hi0iRsJvHVJOVkF+
PEVihDNwen6ylTCLGilmqej9HmnbgvuK0bjpu8/g/9+VnHIwhtzo6q5kmCgb
AyfyxUHe+WksQIYH1eDoPjt9kDD7KIsWOXf6d7HS9CNcTyTRXTD59oCzCclK
WdyNosWak4t1ob7pf4DEPBiNiRtlTRc6eDP4GPcRseJd5in6V0420Mx0/mCj
xRX6bg1hJirrNaYJt3LBQWcJhn9Xmi2FS2sk87Cj7wncj4jK9bFNvGhteErs
9Rfi6A+Ap78knDxyNLQNMmd53pgYgpcf+o+7r2SO002czjpfZNgCkVhoLEwq
VoMCIaVx9f9F7mtAkV9nfFwS8lS0SDwUQLGarS5i5sFtWjwfwGZ59vEuWQma
MGE/IseeDPuap4XIlegltLUeibBeUi1xfzH/k83VyPw5hauioHJPd8KmbSrl
0SXrAZ/scfcs6uxuLvYtIr70TSAtB17F09ucZ034gJ1ajAbviewS+CybgI7a
QHmVuG2O32PRZ527wjJaoRyCxZ+bL8C3LFiSzQFYRZxIcATaat3sp4HnoXbH
XXbQf7ipOeT180Qyg2DEszSwXE4JnmoWljrsYLHVbK5jG+4JW8fGuOfQt3gw
W2t5NyP83LlHAYDgOKT/cSZpUNdbJtWjDu+2ar9PJLqA6vACvGkb5WaLNl3Z
xttUAkGKFyBD4xIHK3qVukgztyuQ9fL5t/F6BOjjVw6YxJGFQJYF+/0qsPQl
TjfaWdWSHFrAM7+4s2+oYFCmbByiKiV/xLjd7l0edRLY0HJSZiqSOZGfAOf1
sHSOTEop2z6eSqaHRv96s5PrF21qi1i2wN5crWy2IJH20Yt2Mksy4bgPv/r4
Fy6lxBQnpuHgvp1SDsyYw8tSvMmtNBZQ2TrhSx+qAjOOwabnRUSRF9gFoW+6
Pb6dEz1f1CC9GA4q4OJCB4zoGfHvob9VXZ5QcPCIKZbo1YPgMzBV/A+EZGHk
65qK3+FS04IXLt9KChfvQkCRd3KD6zf/DAs2uV5ztZ5zVmvdIt921bbgL6ha
007WKMAsvgiGWEfQDkK/1sdk7nwKNvMJJFmF7iTF+Ib2iWfT4+viLNscWRgP
60Hjmm2zR27CSHoNyNSCQfK0MCmjL1HxKsj3vGrMCNHWsies/nzUB3RuUCAU
I4fiyoSVf8cTKybzM2FFickVZ414b0Qhxrf677QNZg4x4ru5pUO1jtGr5Qf3
QbqwXd4o81Zl70Us3+nbt5Qv9Zgr1lKYLodwnQXxQrrzhwx2zu59nUiY8fZf
f6W2aNjsI70kHyxVaWPP1YBqekiQyiVWeUQRQBv6pSAOlM66kUsTi6l+HWrs
VtwvXe01QBWG3eHWxy8enocy++4B50OmsNKU8JtY/C4ed4PCF+8/HyokNX0h
3GG7V7gjeSMzdusKLlbIAtAcRcPMMVWO8wn9cCdAtDtmvsm/3kPwYxm3Pf5k
iAipiipjI/TZY9W69Dz2J1c/5tH9MLOVAghqTwRfyQOr328OT26CXGwcYHIq
icqDkdPGAm6gdF6F/6zr9J5313w6Va9bHqtILRxoEb02XzJTyLyQuIT7t7Lh
LtIiGem7oObvOW/49e+Jev3oJbjNw+P1A07xml6Aq8B2kiPbBQ+GRrJd4IfI
g+L9vcBVJIeqOPA7I2F6VTh/gB5erTEq7MK/J4iafMjOG2rcuU+OW/1oubZS
Qri9Yq9iPZdsFsFigbRNtHsj98FpA0aPdQ/kka9GpGVP1P3XIBNHFXq4WVWv
k7na4dOBPP6kydgg8h2Jyslcp/xmQLgloAaI/ttTqE9C5FVRCISVYTkj95Tz
tx0Lx7jUoeXQqll58rKa9VS23Jo6vPfVaK3GmYZ745a7QoVzs+Ny0e8oYKBR
/t093foFUPBNAugNgYx54qU3c+uhpjYkuH18MXPG1ZJri5kZHe2qqOKCifNt
vfgVy8A2h3nxIjmnznFctiOzDiI719oXoEljWzke0MHL0FP3lCp4Ddaokq0B
roeL2ly0SqfbzYNP3a8OJim/JpCpLsiqo9C6oNbDCXtOq+QJQVWK1G1GHHk9
k1gTqBDB4IaNRP7fYieFVHiPG/bjWocBMHaWPDHIR3WW8d1ySAa1V/lfsArA
LKhtpApXItneOPkB90PvEk9N2dSil8UAPBoZz9mJBooEi1lmEKwy+K0tLD9O
YNU46xe9rhiCHjAlvjNrCD2XY7aHkHJ2oWJkOvkpWSrYfmN9QcsFY2mCK83t
5GUjXJJj8xTw9Cdu9UfW3Zf3N8vCSR99fjNbttR9F7dAywL5bhQGvxZRe5lc
s6hNVTjCxmBPhluXWgCKuscrE1I2x9wldcatAcXnoarPe7fKdc0oIR1mISGw
oWw5mj7F88IRxkihZpuwMwiD7B71lkjPusz9fRvpcVJ0zc6iGRU1KLYZO9aa
UxZVKbQkE0yjBU312lQnsGint3MxbmCoW6PbjALjdKOLzNDD6I/YM6DMlb5n
R7sXoxfnLrsvEY5l4iemxQ5LVUS2uY/miP6Fgb4aG0offCXmVnqnYizkuyqs
Bc2FE8ZB/YnReYa0OkGX4dPARbvZ8mpIrvaqjcd0p2bSfRTuUgkCKrRUEwA0
y5ZpU9cOo+3Ce6ZJPmD2fJQB7PnZOT5mhuQ6ToGrSb/UpgQL3FnjoOiEhFMR
/y8Fjlw+1NHt3/nP0qr6U8DWqNuf51PTsxBp2UrcBfjLJIbl2bVU3Qgls3S+
7q78H9laP8KE6/Di3TiwEK5ovBKhhu4QbGGJSeeKCwlCRTpaUQ4UaFNNwQrM
qYjRpTbtaDR2TIDIeb6PaeVL0qke4jogQwSklsQImcReiJThuAtnUd8+hybt
x/Zx1F1kkTvnrnLmTSq4cLhVAH3YyXazt+lDWefKr7akR+L5tYjD3SIMVTDk
gQ4tJd0c7Od9NkX+TSzqIRRedKf9+CnkEWaqCWsws5xE2H0u/bPWIUEhfnsG
Nrkt6B9jbqmHgvWc7Yv2lZO078dlILrQdJ3PHVHiz/iIzFPxGxyo6IkO7aW4
0kThIYxidjKeih/RaW1/I+f0v9mV4ASR3fhpJL/IeJsNUZVayWsinPBSmaQZ
0HC/udJH+2oXDsYaLdC8/8w8wNi+NhBroxruCx4/hkGmyHVEKHZpl45WjrwN
B+iTtDVq5xRn/gd0bI0K8grV160bJo5ggN703T6v5M3JY0BfPIyWI7bGVFLV
NTFOcjbixtZQwsLqEOsZ5k1059GXjbfIATg8ys6dsVuNRpplo0MUnjflu22Q
z02MShhMBvRwdUsFlwbmelqBoZ88vB7SRbR3f2evjefZNVxiizP28lhW4Y2b
f1kW8T+/m3M/TDeMg1uFxLmsU1TBUPuy9Q7snh5JK5wqs7YD8U+X3PA11B52
wkvSQzzHABLnG35WimMXWtDy2tC1ANbBRtzheqIWIUoAGGsbWFcW/KPBp6/K
e/A8yElMYNfJ+y96M249RezgC6liwQzZV8wOO8mEIWmaB3VSUOxOtSN9PbU6
gS/Dxy/xb/HXfhp8QIf5xfI44A/IZOV/s0pNIRvQF3JfCjtmUTX8gSRfUT5S
9VMq/8asjSUkLkadEMhuMfteKNF20VjNQX+DmZ2NIDp99yD0UGUwEwWFdxzK
9I6H3v0ZxRUPu+fMMyir3KgVlDK5RxoRwYNpdPWbnd+4ebGE3gqi4jy/6tkn
r4vgdiGoDR+QfakjIzTCFe9iWEt2TMGtXylWsfme/dU6pa0BfO1/xzwzaVbl
vQlLPQ1UM0M1sS5/qORHpBnQ+40wT6rPnV2cB2cbttuJSf4VaPx9d1hlgzaK
ED/+fszB+7JZUKv+NHTHSCcpxDQmFXXkK+QsCSYGAiIqNL8nE08fzaei+nNr
SfKPVuEGLwk8sV8dlRYoM2IG1vxBa7G7oL2l9qLDsJptQMganMQcYrwNVwj5
mb63Viloa50aqoeduki/JyZYDJXeQ0WCZJ0stEmLvj/Fzdiud1o8Cof/0Zha
UwnaY81lL2+jYgqebPmtPkPeKMgdYjqfvtr3Sj0VD5CPDLPLS1vZcb48SgVN
85XXxy0O0mczVTIkKyd5Ib5enAu6eKoKGV4yWfycTNGDeJOz0DFNeaYrp8I4
qAcP1byn79cgynfH14/QmgUrqYyTXPnJre73i7aP0999s9g7DtElLFYIHmLg
gebDO1EswTIBsjpdXCzW2Yr/qSYFVFs6NKL8rlu5jaaqW9ElUAoZgXGEa/J7
K69V7Wu81FY5bAx05Y/NCsjN9MM5lC5Fl0bIvUptfmCFS01rB2UJxiRJuh5x
F+o+GZyfbW40uRK2Znh8U+53YNoIEReH6/wnwDd6GVbCLBB6FcadGIM9+LW4
qBL+wSZ0afXOei2mhUs0ypUCwYryWfwQ1XEnMSGa270IGuUagCLzyP5bjvI9
fkt30Q+5OEYhjchDX1xgJTPFRF9CWF87A9BjDayifMjH4cHBgdv8Wfl3BBEZ
G/qISNVDW/BwsTskjHdzMBlMP26CzWaTZJVoinMdITs5bcf28W0YOjmXjQ8m
yBnr7GgrdGQjo2VKdD1gFXoZ5N9VSJLU3+FcpxdG+KPSWubNt3qR83EZmR7z
u4FjpOCJeLAEPccaNWnevVWbenAJZcbV6vSf7p0es6RWpIKqZ+zyq6gPQyZi
3tNsTD4GDU0YhpWyrfnPenlQvid85KAjNBy1G5BsLayHzzgOf15qEiLFkEmh
H8mupGJvZen/BFLXyTl3qFhNngyVavUV5LVnUtRaLAVJsB5nmZ3Vpn6ZXDJ2
SiFBJLf+KmRh96ku1k7aPDzPCgFoVrjMKcswmASMmL21DR47lvwY78zeZije
aOtqjsGCuzZGWve3By5479ioSQ5EMS5IxgN20i+YqMYg/zHHzQkGPfJB2Bwq
g7+w3sgab6FcHBhw+UvP02onszD5RwPDB+PtjDAv6oWW8xkfPoKR8+kttoq2
scuEQGqYqIFJTpzqibOoaKu0eGRCa/mtQlmjqui66f4zEkZ1mxo2ZP7viJhW
B3g+VrdmVZeG2lvb7KW4HboeslIV5bpXJr8VgB2sW8A9/aOUJCmg0tGVv5+b
YGE3/Fr9GxKlFYAkGJ50F/lWOh9QlDh2uVR6Rh1+GBo0GfkO2O5JJk5IqpWg
teUjdViJKTXUuRXoNmsCix5gSRfmE2LaJpBu1t4MV+7UYEi12pTZHHzgYc3d
L1HVzvwCjGUGddW7Ny2GkwRxrf563PJJC/pAEzmSe6/6Gc9Q2KyNJOeYbKe2
ZidRoncSmWPMQNreiT1pCGMUeXe504Ep9YY9Yj67/GuuH1drLg/gAL0tUU2a
hbkvL2itxo8YX6RPDvmkPDoR9Ld0vD2bZznYMkYagPujp6B5L86wjUkdcosN
3DPeu4vycKjE7w86VYVlwhWPUjn0cBG/RzPRe5Iug7R0GtELszS6w5efgwal
kA0KqfaIDxZ7zkVfz/RmJb0kl0p9krSi8emUqkdEViaRPnde3gEh2eZP1Kzs
/a0hyeMa4XATmSjW5JLVL+OFnpOlVvh7Gpf6T3AyTCgBxLgsdKphOPub6f0P
1VwzC5jDr5Y/2aUfdCcfpAnaJmaIIw5sh1iqIudxUdMDC9OYBbonxAHRUvVE
lE83mmXeAgV0+tfFO7GFwcQwmrsByNu/jGdFvW4y7BuM+xv0NcFSdubBor5k
Fhapi5QaPBhUOjxd80kOYDk4KAi3jHA/V4n6oPHmQWx80OTRy2ZEDWrWDGny
v37gjBml9AtkxMw52loahF9WeN9CuiUfejAvWhaVUhxZ7s1XtSjtAON3wSiw
43tQM66f5LCkfkN/jRhVmyCGh9igNUo+KaymhLN+iHEf97gB6mi5kfhqZnIt
gVSUeaHQ1ubu+NdtQqkauMyvs+Rw62mCXB6cV1sAricIhItcYEujlUoaM4MV
w2WgCO2GVIL0bo4GYmRa6DRFRWAzY7qwChPW6zlZD+vwmhURAWGjYFECdqwx
W1+VCAXcQ9CWfXi128gvAY771ET5WLK6L+lJbhWNHEQihxQQFO27xuqgHLqe
SImC/DVsWFVmiA2Ao8lKJ9jqnD3Kk+OAy4/GqrnvAuvpoBGxN5c5y7X3jezX
Z4WIU9D/0w78fs2BNlwjz+8bLwg1qdbQg22XOAhKP4H8K6a5G+9h5rJRvaPU
RWbVwDROn03dP8WYmG80gbkk8O5RPwOHKE2tidIlKVDpOWurYO+bSBjiIP8Z
8l5Tch77FQPEztGWVwdXLQ9yMMKOZTTwPF2iAIkSv+zcigSr48eBnteYuCEL
8R6JlTLPwHlksDoziNllrzgrJ09MuTnqmYnmzmyLRf5w1XdYLOrGXKPM/KMZ
6wqAmiBhPmIqdcXe34Q4ANv27ico8OOlto60G3WKB5S+NzjHaH80Hde07UFH
S60YQFzsQ4TwX2pSmuem7OOU5fnbJfxoSZfeCL6yCdxQaL4lKBhUMeTWYxA9
9IScyk01S/iMsXCjEsJhLkLBZeQpE31igOpwbfLJjaiCeHDwPPnjwK68GeBR
xDB20QTvyufHvC2Qjn39c7qFu2nCrKaZ96CTnyXD1Y8Jnxry9fQK891GAA0D
dBdq/s/ZFx8iS8Ve18GaDCijiTvtln215B3P6T0sHa7WXQrjULR5gwPFjx5o
88/GfdEs9lOp47BTBeCfQNF5+9XWooCraRkR/GWuUA/O8h1VzDat39hpuLza
lKzEk/j7G6SrNegainz2dPU7OwL+Y47PegFoaOdpNmtJZDf54hGsDfddyw/m
CsHw2W4unwk9wgHcdR/GQ1o90zEtq9E04iAWQeRsdynzXLTiJZlNkLipl60o
hl3eaFtlF5RDF69YZ2etBDINLflv2fv4hEFzCD8jFw4SlOdDYLCL5D8fowj/
gEng3WqyP/YbVIQu+GPZ5JOB3dXnb8QBTKJWo7lRTixnM6FS604cpN/KJoE1
SDiDUkUmvm+9MAkBkJ625WMzZupwmyqH253iO5MMKl2h/POltqWk439Vnepp
mVLPX/PWBCCWrxBNX7imRaIBfXflLzpKwH+XIVeYh/MP/K1s8bYvD29DLoM+
CY6jttM9ZB04DlQAQyiJhndeZbeTbRqF+LW8lQCzS63XpsxrskRtJzhueUCh
IjMP5DLQGbm5sAA4rlN/pit/2cu9j5RkigVYdivEOsoWK9b0h2oSU5TiV519
BQShW/DAAYv4Eu7qMtppUObqKIJrvFcDTzWPAAVxnXTeIjMOeXDGMWBJgF4f
Yu9Rkv4CE2WLZ+DKnsI4OY8zAUx9hjIR5IqnbHUvqzyjXCmvE5glCi8OhziN
8I2aB+371VpAnK/s2P1+fRJDWQTVdovbdvRa8CBpXqbBoEx5NCLlBGYVwdmH
brRJhAOqbPJN61Q/A39xgrQtaOVIO5rkG75HIsmCDJCbPQq/xOd0PAsdSMkN
lDvjokvRATrk0952cR5ALWBIWsyx1sj2zH6GV5kt/OBU/bJBWjmnsqJIKx5R
tA89mrWdExICfPRgBbeA5U3GfLcrYEvV1xOx6pQfrz0jrg2Vk9mOxHLiZ3M5
4g/qSmGhdDdjV/jgfB5nQP9a3h2XYpa/vpawaPK6CahurWXnYrx03sXWNbnD
qxSBAkk6M9tD18GkxeEHkE0xeCXHjS0dfYDUo1+XQxgvt3tVn5YCCE0t9I3W
IOkVDxoxzSQOxteDjqiAnagv/ekNMUsHtKc8W1q4e1YGrKR/0sa1sUjTEjjT
gF/6RAyn+Z4JcFSMzO9HvljW2+6QbnGUFiD93D7I1BBffWH36LaB3BR+ldlN
EvYF5FKV26Cc9UP7tAKb289iladFb85JKHZpQjj43EvalxiNC3qhNGt+pp6c
g5WLsYgY1QHhjvNf4MUXXq+R1nweE04CO1Jrkdykpb40na6s+VSQ3UwPuHiu
HjC+K8dhTnYzagbwxy2+T7uNOk03GUrs0ghDJn0/k9MEv3j/B9e22sd6/7Sd
EbJIThnIjXcWpsEFGcpc0/Vhu1OqqgeRyZqfNu3aPD6zghZardHPoemDT/KG
roLit9stq1a1z5WAszj41kEIEn6khzZ/qsjKYCf8rjI9C7zkJB3B6IkZaA30
OdLSomH1CVGOO4p63i/DSVIXhHe0X+CrhxQ+8rGnbcKpX3w3aW96C1T1Ooga
EXtP5s+ZzruCMmvc/FOa3w8eXwz9WwD4Wl8UFLoktBKt+jxT3hTcXkpA39Dn
8OXbR6Y6TcVkrsCYbqm8emx15eqvzXxRut8dIFR9u9yS7fwVNeJcKhAMeL4b
DdaVyaGQ9HItKUKgoxqjED65hLhUDOQ+mQOuHKoAr4FcKuEFchOUtEKBmY0C
cHqJGKf31oyJFexY5fQmWKQyH8DmD7ecfBhGN6e3igsgUdBWaji3K+V+jERR
J0MVv0vUkp1nvgv78wRwc/Zh8+acVTm+kPV6HEY1HRKssZ7q1bricPzcPAFv
N3gbN4xKGXuNfKHUWX4kW8rYpqVvshLD4DRWZVcYgWBjOUJ8JhIfSw0Svjau
1Orl27s3ItQi1gVs8HJImyp8rp73n/iOrRQmZY0D7djkQtTqhoRNyTrpuuUE
yAvGt/jySbpSPBrN3+4ofgyoslF0fOqvwYxQndnXGtgiF9hq9thpuyL9p2wb
csLePxt/ZiLRYxXE6KNRABJJfxcCZzRqDApPMYwVzAZ256H2rGbZ2tuw5DCC
oWcVF/CW2O7mseuu0PapkawyWbGAzNHJbkFxRbzJs1NKd9f1Yr3N/5gdx+rN
yMSMTrTIbafsFeWJVWoSAlDVwX/r65kYDbwWkvZtBZW/ZY5Y8ssdRJNijX8x
QY0tDKKXwMD8m7moaH0+lEcLyPNiMhCQx4lqnGOMOUPoQybiqgL6cLQIW+tm
rHNwY2wFvu4Pcx9aGSz+gC5rK8eo0/j15H1WZEregreYcMdskU9otJv6Topk
ZhQNdX0wfA5gyvbJB41Hc1/v1nYMWhizxDbcElClLpT8J7Cq4ot9eaKh6qSH
PXpgXVx3M+taSknB6Yh/6uEL9TQxaDr6TpUs/jG3wbaszGLc56o5MH5DChOD
rjMxuTHaxTfhB7r4TUUntt6jVG5xlB3Mo1KE8cyW5tOmyQXiFXrsDOYQAi6O
B5fr8UwoOw8H1rV4XUEZlvmvxMgnmHIDSFm5xNP+okFFeX1oUFCjn2K2ZwVm
sSx1Szbr7QDdpiPwbeuJVGG3CXz/Cy2up6q9gSXlu/UGd/ITxZMmoj/kVDTE
AZs1/ay2z4GvAN6hQId3H3qsPzJnq+ADvULaFNnpjkJ1fLwWE+6wr1beJnTX
NV6xUj5oFOVR75E3h8jwI51OiHU+Lmx8A1GW9rBmf+IJ73IJm2mNb28qLCCJ
2LcZ14nkJsj7OlggNWV2Eh7pEUj4RCF0V1g8DZ2FpdSFon07zHvQR5GT9ho8
xsueMCJ3oMr//2LablR9GWmXTV3z2CMvD634kaDji5itStnMpNrN9cDb3c+O
xigY/NQKtHW1aaP+GeUJZpWrf3nthl+fHW9g/I7L6j6r7LelgUK31ZRLsTrX
wsZPDkmBDHyQX2d4gjMAOrnkMocethFZsVHwZI1RmDbHlPg/Iur/5DU8GNjy
CjYRnTdXEyaT1Pp207Qp3prRGu4zyLfeYROD0HE79qHHtSK97DXONcA7Xb+z
t1lZd1P4csQj+WAdu7C1ZaKLy7Knk+fDQgBjPWcFRjGsnrzD6rbMuzRqlsKQ
ybaI/bvjDW7ZhRPhCENp3Xjv2+YXqBnb+o8zY1ZnbHX9GscBYRVUuYlV6/MW
yv9LJvv74ew51q6uXAiKhenv4mYswhi/afMBbgeoQh0GekZtgEXBzco8lnu8
CBCgRQe43PW7nY5WFTFKTWl5HaBhX7pc1jlUjepF3wmmZJ4ZI6IU4qp3/LmQ
aymuMZn1UZtvUra3uOvNjMHA8LTB+bfiyaTpT0c9bdOWIhL9LS8Ju5uEct0N
t/sr9mIfIyeucFzMq1EUPaPyMvWU8GS+yHRJhIFQorcNBk+xshvqVocDQCct
/cLVeJoUj/z4772lUOtuRz7RzMHI4sKbQYNiLd5OhOuLBw14HXRr1CcmlbkE
OFr+Q7ysC+5T/vNCnI7JFDSO7Djeo95LzUXdCiHGL/NdEN1wBMtsytWUTdk3
F2VuBxtftBtISsP7BfQ1if/zvUxX4cmT8bJtiECmg3UkJM8lnH0ZhmKLvsK+
TD4sGQw17mWOzerepSqvUWBJyYfM4ZTxz47AHluCk3l8cKCcMBTHWAbyLATg
AGXW3E9B7R2VMymGbah9H3FXRaE+PLhwPu9XXC7qBOAEg/S6tjWR0RQILuqR
JTjfEg3yovMMK1dT+1tfmvrUl/PH8/iGsRfqocM3/AEifRVto5EumZCrcAHm
dpUsjXAYNblGYn8LGQfQ0aL3hBudY4EL0qzljK+dRFfuhrMXjhtUoPTdhPpO
SZvJbLqKWMNZ2qhPBjBsKz/gtJRm+zKRzrH+tQKqwCsrJTaiQWmgwV6twhqJ
+Ez3uqvl5lqiue/BGyxD1nNyjTCeaTTlKze8exC7OP44MV0AeWfuIC44t6Gd
6pnp+MGe7BRX1WVsf3STaVE2y4F81pGmQQa0+OvzbU8JTF/uYwsRvHqoznUG
lgpac/Wh+fqhXtelS2uLBjkG+eLCHbWI1RyOmd2+dScaNlj9Od6jYp77nNLU
3oRIx3mUg1jp2PUgQ5m/ArVUHGoEmPNd0NRhS8TTWLtm4JNHIBHwsCOe0ndP
gejfv605naRy1vxgil/QEtiLiYIVEpKRekj1hQk2P5j7mbPaCDQYbatLHATj
JAfFiMHcI3O3r0umBqIcy/3nipJS/S7b+ecyFPKqXj99QHg89XMnQ2faG1IM
Q2vVzZoG3ArvCru3S9thtMwrRh9BBwcJtLx+dP1D7SKVtJd/xIAIxs+7TPE6
FhJahuhc4YzR3umpABtBHXaGClGyGy7V+v9rCRofhlicWzcWB0gVRHIf040B
9aUwgczCvEDmpceVvaUOCLe34H48O1PXVPSiCfZ33zduZ4LbE2yBiXToiJyd
W1Jp1HdJNzyIODhY0VfSp2KylWNeP11wcS1p9KcwP7C+ddwKjMOqDQpAAQHm
pYKUkQE4MIM5LIrqD3sKw2NhWTkMM3EwqO3mV/kVpxRcNjLaVJNm7V1opeKz
vih/9AQRHFpvx6YiL9TovyH54dKuBfH9bcOk+ZhLoJXrn0VUx0Nkf0uwOc9o
tB9ufNyiX2lIn/0zInYUq5jpTXP4z21DQHGUbBxi382DlX0MznxAw1HNxZ4+
WbJsIW3e2+rhjaxa25JkH9uKoLid21erHn6oPpkz3q8PFuNaOyHzN6c4GTG+
odT4G/TnHCQNUewVrA0lliu5JAc2jK+yD2DO+lM72UtBNQQsr7sIb6RK3DiH
GWq8K3xIekAfryRM1C3+lShbTnV3RG2gJPKvNkfnub0Aa6xHyWI2AVPjSYHI
51EmNHEMp8/d+vknSE+/wdkxxsmeUzjP8W7s2ji/j7Zv2iuM57eFBOEaoUBc
Fe+6BQD4X0q/gmk2BQ8CShwu2WYmPILdOW6By07bhfU/lQSwEGUD4I0qeXbH
0NfeDh+HAYUNqh8SJFO2QNcy9fTv8qk+Rd48aPo4bWg7ITnS8qbR8TX0T+uY
WXTzw99kJ5juzum5UbNcu4Y6KRekO16Q4LJRKRvPWa28w6yH4gquu21O5pV8
Uy9Vs98CiuyJa6JxNUEHXxbNTZf8p9sGp3WiO0nS/agxFs+HlolYiLtSbKw4
LmuHydwh8OrkOCfWeOkc+z9agUD4Ri/n/D+n1X/nq3DfhjZkAhN8kHNFzWXG
j91e0S0L76eXV9NzTxJvHoOYglDmiOaUlNvOjc9NfS/KCGwzm1bLR6y+Ylcw
zVpnjO+lWEaCz6XpSsU0I0l140JnK//hkCN/Z5qhedyHo1B8+QVZWyxMGhCA
yQW6y0XpPr+4QOMxQGDvVRvC2TB6EoSBrgNCdCvMuML8VxlkUzciZ3Vxq+LZ
KyzRKWHkI3wFDLqWr+Ewwmo3P3DIs4liq33EZFvXgrbZQr7dKokAfQHQdXWo
+mcBj5aJzfQ9KkTDUGEGGQPNsPrMuMDMRZJ8cObZvnguejqbGsA9fKxLYUzF
/xCJJ73W7q9IS9yk06OGB3smSkGw7vsDOqe/In3A78TiMbWYOegGzR1CCKeo
7exAmm6dfN5XKOWWrW6+ozcBe6PG6Q3Vf9WG7FxU08/eYtFlXwhABRCPpC63
pfW4m1bTjMVPiGemXFIV2aka93ZN9CJfnG2EAMJrYILKaOhxdS98pEEH2cIe
gz1BFLXs0+XF9Jl9/p9HA3NX4P1OLlAdF3Ac7NAniCwd++n/GtQR/XbPrLVW
J8NBevUsTwmpKGXS/Pk+ecCRw8dBSOS4ZW7mIvK+ifLRiZ/XKxeR7fe/saHD
7K3ZwWnb265SAPyySJKUIS/tk2xI0E8hBJ9j3/Xblig849SqgkhLejMzLzyY
AolT5lqKpY6D/+uqZMsrRDXDZ8Oa7LSbWVfuYETG0Qqqt8sXCpTtDdsN7+/t
3otbb9HtA7oaeOCI3e09MZqNmi53GXXd+a4xH94F1j3ZDeI7RcVWimK6I9ff
1JMpQgi7d5U6XJJhBXzEusXzAFXzFO9G8AXtoS3WmqtP2Cdo8tVLIcK4kVY0
aiUdern9I0OP1PGT96jkj9oDCqMtsSXCH/yOThtNsvFPejTCKbCbTStqKMbK
vZoa7VhN0X0NqLr16UIx3vGztAkQfxLqykXPMAEbt2LnPatIknSJMN7qN67V
FOu7Ksv4JbaVBLcrFbB0ujgv6KQq/6PhNCiWyvObNwwfFD+IPyLaK3/zuvu0
ixC/9iAbGBzB+Ut1iqdvMTkWTztHEJ1nL11DoQlTp5mgo3RtuawEPVqxBzE0
qOPaQxkekFChgPEGHfFy/pHbfuUYwBSZ2QJeziLGhdWyeD6zfjq7g9PHcT+l
kXdpcb1byhKd56VZkd910Z+wXurCB87WympOkFvcxJxqIw/Kq+46WFJ5Hiby
dUEyDYfYRWNCZSB7xvT3W4n2M5bg1FxtYfWZ5aoSkcGTEyTJACrF9k2XnXJS
m0KUwtds1MXuPXhbzhLf19F6chO5rOLVZftyZ8NoSD9LuXqn0DKRKlnhvdnB
6e3eg0Bzw/80LMvo1Ky53/3pizv7N9PgFshgM6YiZRjNTppfpLH6oIvcbY0Y
Wwtjt174eomSmPlZ8GrYz8ZsKpUM1Tf9Sb6xCP7lV/2unYxBy20jcSYGc6x1
oLErCdejb6n4L1IPoDZ5zGsj1qv0lTlI4Wy/J2klsDher4Pci4LOjvgzKmgg
52XhcVZ2Cz74+qGihKyIFdkbmzCcixA0+WRlQSC+u32tK3PMNHVhHG87jrzw
T3syLzkAkvgFGnZwvTT1DLPBvWFmZQ6KAQHPYOD0fMsWbEwHduFMrR94giom
8I4V6/AKdhpNJCDbex7ga+AuIAzeBaGneiubqd9XQz/Otw40kCx5Iu2cu7q6
i+eiK5yS4jV3IPzYHk/RlBQ61G2q1WD+PsBtXpceM19U4KvI4tjduPxHRarj
BzdmONHcZRrxD6h/3LAz+L7ceE6LW4ZJkW2RTmJ3w+vGpfAyYns6FEU/uVXn
JJRp37LJwvIxmKXLJcqFLM37SujnkgaPquNGjn/9n2Gt1KQ6HWo0fxeh3xEu
ZM41YxiA2qjBA9SJAMi2dYdsCideCbegFfzaloEJQ3mL4j4Cs5DCfDfImTFA
BmGdIZhEVu09PfC8TsV9OKHgyNsC9RIttXDCSFRFTWY18dd2slf13R5vb53V
/K8yvhAGQb0NTLPC1ltJ5EqI//AX+FBu4kyTkg2JA41tG0xWMJmmmwdSYm7l
oxzXior3L/xSFFuprH5evrHp+7j36E/+xx2BKxskjLUD7w8zJGuSn8aDRLuo
cTPRGuHX9NttoIFaYNpU4IP73jT1OF6kFpY9Qz2oLm7cPWC5b2c9TPQRdVqj
uXmQOQZj6d25S3wPjWFQDl//C2NxqIdkDADD7yE89JUJapOiCrrxWmiMjCv3
eP+eBBXVxQYLe/wIL4ySssZD8WiIbXkfIx9fMuEayj7qLDTP/mSot1b6Isgk
CcD6ct+sThirnzSONDUjnaFczSc2/pG20nSp/teiBhIqv0OcgixqP5TIt3cq
fKMoX80S23RoiQ0CXqC/K281EqXXgFjbn0OCkcb1zzN49TL4l5UAUvRJinmY
7Xy99lhjHiZwnLyvBbHKM1YBmjIJqbRaXsv3xucwnj9x4QDjofvKNNaUAMop
U7B2Ghhs9xOK5tKXKdE/JR5wuMk75yLSZjwKnykOl9K6+LXUZxAZrMoRqXQX
OFvMEFlwkB/j7gBNS2fj4tEWLS5BAUCqawOPEA12oVTo26MBp6E80yCKQrtS
XLVY96HiVYgOkEg5d6+MIWdjmGxuS631a0UHMzkUL3hvcrUXGTP/4izz5Ngc
GHItbszRH6oO89fkDrNxPc2LuJYO6+bVPH7BPMBkXw1lv21EzDbIw3kZvEpW
nwJynGLJsYCorO85RRQ8tTpxi/Cilr5HdmMXe/Z8RC0EAvQf5Jztx771Ae/G
HHsK0FxMeyhxPhMXtoZncEGR88CJ4vN6Je8jn7NxVCnAQ/xg1JST1vxj1DVJ
HqdyIZNEu6sHBsAzWj8FJ6m3H0Qjz8J/6j0NanBJRkcnailBEwRfhToD79VT
cnohSeTGj7E15c7cqbHW0m/hqPurtwzRnDZVVKV3B/CFKnP/aG0o7aAqLiX+
fdgA2hzWQfo+hn333Xvbc5NyOI8lsLtb9evv7IpcfCQ8YDFRrzrtbRZPtEBf
9tm61rWY4yqdHsOrY07foASnW/qUIKY/D0Hc9sy31m9NtTXOU21foO/cvrf1
TV/f3H7kFTsIcxFTwmGn2CNa2vWihndsL1CmosR+yyRRFMD2KsutcQIMGVsS
igUmza1npZ0pylJfLrx4SO18i+KiE9qps0IcGDWw0AzXSc2WQE6Ixs6nJnBw
2hix6QK7P3bJ91+pProaysouxT0rUJVdNFmwGGqTLUcN1oIZfR8m/nsjaFp3
atL57Cg5NrKzcLdhSGcmMzbsswqPbTAsYPK4EPyDUhmkDPK3lmPyL6EanbQ5
lqLHU7Mw/OHOVvrpkbk8CvD5SpvEpB6/0kGn6ta+SHZEZviXxapt/AqqfkRQ
1dPRPdW9bVdgvEp5QEKwxZIIKV8oZyNGRrQ16RCqNvIY0oOl435rJRSvs7VH
dOtY0Cohn6qVobeWMwtM0JSe06AJH1IlntBau/+hcY0PbEYGe9TtF9NwHTsg
8hSSbgteuKoZc8Nzpp4SwP7QbJ0Bu/du4iDnzIo8dgwSDgjwLPqq9qnzNTd4
oLEqsFlRDRyeatYt8gs+V7VmDgU0BVb/P3n2NafTkoQg5CROU/FuH2gCPUgU
CGAWJxigvmmP6jKUCjYuxWLkZ0eyFu/7g2KlKpoc/RJZ8RcE9TOH7Oe5cyhD
X/BEhv0jiUW4rTDE8S89CbKFi37xqJyftyk1G0Mzc1MA6ZS9+ucnJG7b5Auc
LuNvAQATcT+WjF1k82ueVgKIFhUN7Z6Yu7evq5JO5OJoLWFUHpQoZRJQAzWB
f6GQ2nsO92eRK361cFGVEdYvCoFDUHhbRc8KgFOo1H13oNvOdXO3Ii3yMqkV
LPdiiXhZ24+y1Oh1tpcqJX4EyzvI/MS9FL+bqt5RMUw9bhYDKmc668U0Reb0
bRIiLHWcU6049C9jdN8Y7nNAIWOu+yFTq6path67iCJW2nEU+K8peyy3Y5fq
1ixKB1lajou4p3vMV4nZFa6qjVCS93gXn1FXRl1a1aw1diDSRQLYIaLFvB7Z
lBQMue/6b1P6dFvK4H8lQCHtC8mg3+bgLBLPWbcKu/6mnYwF+kOTwsP7HOV5
Qm4Pwd/UdvwOUvhCSgOIDpKzT+kXqnxpVnip9ELNoVu3UGRTjOkv+Us5DWUr
NP/k0OeknoVeGMuW2GP3VeZf+s7HzWJl48/qrIJu9g/1ec23N2fzmo7JY55O
FvpGfSsRhFhYQIUs4d0MMVU7TZg6CHWLTsX5KdcwPX515CdJKTt8oMhpA9MY
VVsU9596GpUO6Fl432RRPcg4Nz7t76sqx98x6IKOMrsAF3Y7/ulM9yRPBrCB
ve2eBVkLmVyF3ZizwI42P0sK8K/oRwxy9fephaDRZITQlVRkTiH5ffRB/HLt
aRs6/ljhivYRW5WhH3H+33IVJucIYKhP5jEwsCStn1tf3UpESCqTTzlqKAU7
ZHeHMABhw0wUcN3QNTgpGTWc79iPKOyb7+NT9+XoZg/5hPS/3zi1UbBkCZqT
+tf2cwscQhhBvHbS92OGLb0YUuNaNCTmINjAprlJpobeQPYcLEWhnwx1ly9U
O0/6hMZ+CRR17TeOkcPFlbFbLXtaEI1FcIB2agqunEh9mQm6r+H6eat4SaFe
34w8ayz7p6bexcefaY42stmvU+Vbdoj7MFfMm17g3RCYYSLR+J/v2xk3+SgT
H8tb4oMn189zHBNfNJAVV0xVuw2Bww6KEkc2XopdQR7PuLhrqV6cdtZCROlp
NZworVHXSHB092u+xuvD2m5o2/vgiPZavRSKzJXTGM7rRph02PFyOXqYT9pc
35pmB9g/hvWTyAviv0qAJgXVMaU9p18GFDOoHeeUghbjlLBwbd/UXG2UabMh
+puK1wq3raTIptG4SNIz7n+HsXZM3+te3wvahCjewRogJZT2V7u0C06Mfzos
DdMTetTaCAYeLU9GWOtqGemGQ18K4NO54lQGLFj3UbsBdEZrHPslVbSBB0nJ
aQS13ttkbGsyOtJWEBdhvrRwt886ghwK+YGaxv8GlpHPQisKGtN0bn/4PciJ
DdvndW3uwl8Hs5fZrHPigPMtshVvhtahvX3/3n6Cs9jNfS4iznFUP5hhj1bR
Av5nH+z3c54TnJVb4h7RCGMEcnQ6vTgVbCBVaHTU5aq3AMyGYSOkK/+AGfdo
1hcqi/jU01OVwFiGBllSsKhVC4yQcfMBZK1NxnhMk8w8uMVqPax3V5rTdVOH
7RZG7lV3P6EmQs8a64M2s8VZuj6jpVzv6SdNSSpZF/cUa09DL2AfvvcZ0XBc
R8ConRX5JyWGeKu2OhcFgFSlGELZmbWtRe07uyEgANdbOTzqsannz+P5k/Mv
3OwK82Y4q3j4DRzxUYsnYI0B1tjaS7fRPYyzs4ytcI8RQwmM269PHIktpVXC
ofXAz08JjCx+heVm6OnrDAeBPHVwTW+CUX3mQpnQSNNPzt2Lt3Wui8xReZqF
8ngYRr65mUOas7hL5jDeJtlNfWmbFLGET4lDRh53YKl+I3zIrN3W4xLPabeo
jmoEa6HSf5ZDhK9NGk5Wp/egHYY+Z6i1mCwERvb8ltao0R3SHE0yCOVPF0U5
9S/KZVC19/uR48dDGfnN7+4WGVmrtm1nu00WDVAwlUKHgnKR/7k14JnYTZQL
Fh1C5H2b+oohSviaiP2owl9wio4/w/W7FsAZwg1S8+TZmeswPLuo4x+MyDuB
dTh5JH7X6m1hA2C+1ke23Qm5VGa6XYIhNz9HpQA3pkY0DnT10NDrI+ZjU68F
CfKGZVHZK+kmh/csmL1S+kY0vKlcDggkaip7mMpMvlN5fyMhhOrufR7Pc/rC
Y11eGhaTnZjb8p+KlGnOBBw9IGIu+yXdWFVgXelMSJq2k/sjWs0b849VZgMF
VZfCrVQAM16EajZOqeQO1X/JImirknR20iYN0JLpbJ5+IWjNFf+GPN7kberi
y0do2Gczz1EO4fHE4PEt0w8LFbIGF/vaBZQknjFQGmFKxwuyOdRqGQNbQxuh
ttuJ7ezlGBt9et6IoD9IzprI+Uge2B+JWexEi/fat03u9diepu4v6NWihk5h
ZdzG2hWumpGVJutaGUaPHGR4dJ0fv5ZV81Jj7s9AmdyTPU4nneSVlsPAmwRl
4LQ0sg1PrzM9/WcRXWdK6igrXDaPnGlu0rhyz10khsWzjVncZA81LqqCzINN
Euzv30geTzrzJIvcN0lBF7sj4cGrypGajptsE+jHtSGerHeuj97oZzsbaMep
QEgfpjcPbGwR78TRW4eo24bXeuVegzQzA6ikEj76xf3uysBu0EII0C2WhnAA
+c61ZkSB7E/0iQKaJQ2mBt2e6RAkacu8ARDHrjtR2sVbjgrMxAFkWlYRacjr
XoyF6e2k2BbPF7Q6XijyETu8v+nQ6gKxXyXyvxBMwQdCaTvKq3svmECe1m30
ow7INBnjF+fPaPvp5gU4IieLwuaTwZxEEQSjT92FyMePEpyOqTus6KxJISjT
fMxsM0uD6cvD4aRts0iFZtBueOQ/HsMttrS75RFMX2ISfa+sN/abAkmDFzyo
OOd8Ho8nANNR2xjo7vjDT5WAKHeNiWFeTRPyWtWnfG2s+/0uDmTcqiUaNad7
qGvICEfMA2PIOu8/v2l50jx3vbbXKU6HmbfHLyVQCZFXPeC5tnZj1q1ERD9o
rDErQkjB6TZ9SQ5pSFj+UpRb95SYnPdmMZwVhZ0r+2/tUNRCR6BkZuxsttRB
TlT7DQY0Erc9IMd3vbLaeLtgcECIn9slqTu5ga7Uy4eMo7xaN7RAnKwWh5qf
MsFHsYd3BKWU2XiSH5QcuXFXnHx4W61/8vJ3Y05tfrEAdkSrmSOopCBc5ggZ
OreTbF4s7omxxt0B4hjnV0s1nRlZnke5EWODlrZymY8/NfVtNilE4hVpt9Qk
gwt+PscGEFwCoZrpaEUuEUpXL34g31ILN5/dhN/xQXYljUG8BnhPlC1WQfOr
vGysG/BXe0q1mw9YabD8237sxcO86mFFvjIuBtCcTOq/eG4DH6+z6PipaLHA
UUsuvc/PSaX6M/KpOaAuleBpmLDtOqlKsAwk061hiUJxPi+nq3GDvHECcjjT
BRD6VBPs/AkhS2sc5zSt9cdTIXL/wGYcAYHFQEITwcpGf85gQoGwZxGsL2b3
B8F8mK0wLJdYrXzzL4346oig6rrbazH0M+OOZ5fbeRkz8lmpNY6aEPI2gbnE
Hl96c9mrhRaRcjlPoZE0ek2sbH+5h7QlErSgTnCjKTeil+A0oz91s+PAyCN1
giDyQoEc+5QgNkTW0r5PdWbOLIM/1+r2comC6cgdSqnPBIrgfe2CzTZm4s5j
pLsAL7UgCQRbROUmt7R0NOlQD7swwBN6f9KjRwijqjxG1Q9rCD92jRgJdUVb
yE4c0jRHuOfeu95sy43j/FRa/XOLYz0wfdIeS7ZPFdyyN6wgNbN58annr4NC
/h0x8ceP1typXv3/93mOzL3v/ToccutqDMYWljqdDvomKDXLofLp/WA7F1dI
31ZMl+gqWKu32mWWIPHOCfK6e8qttVq1kdUAJwWCEUOmqQCtWKEo2C6HCYa/
khEZTezpNZXvFCpC89J1kOfEAhIifTzAclqwxNuEAr8zlzECOfjv67fLW5GJ
216C1KEGuiNAwtqrvNDdr7sHitIETDcCCeArfdzwX6eE6UZuHJf+ByYLyShd
8s0fNXZhy6Ln0X65u3zSeb3WvpC/erLMmAunw4iBcSbPywfpfTOGkz5ZtTzo
WFmh52oOc0vk0TFw7RKi/oG9uTQ1Etnfvj6InLOZp4E47p227vte8rheNCmH
8FPYnYTe3ohMRAjgpZpEDhFl3VRzZ6LbLL7fk2v4UxMaPJgrj3ltjbPy6uW5
QtIApBq8VPPv1lwEvdpfAd5hI10krn/StjWv6ParjJWVRQ/+WZm5gtFlOwUp
vd4rdGfnZpVUHSHApFVaHEgpoR5pPC9a8pEz6nOBMMB69/Kt/J0uamHtwv/t
1U8ghtALPC16p196AXMm03iwXkMn/rZFnS5ZOXrwTSQhqh51qxxzXeZMKREd
ixunwOPxDrD1tU2vNKveQQ4KYbmfrNJEq1q6r/mu06Q+JhalBgFzwSnsUnzA
5uFA62nVebYZeR//XSDgRV1FsmHlHnCEP2+gPMNJCW884jdZgLQcx8uPneHp
navPoclGBNDVTlPfQU1HgZPbYzT0RVMB95vRZUZn77VZvTJFxTv7w2Q9O83p
IYz/ls9n8uZxifqMMKQObIrZkEoyvi3zUebNuzGKSo+2mmmZ55PIb0e527kb
sNiWkCyLPVNfovKuoHDx7/JmHq8dKmDdU3HB0We6ASgspx2+xp+Y3sntGq5A
I2EjSSkJzbfsAu+NoTsLg6DM8rFKB3oMwIfeVmjxr0iiOG75X32KQ9brYfMN
gttdN3U8NaZNl6yWgQ2g76887b87kG53JpILAaBSVP5Jom3U1y+uHsHQ8VF6
Q1s8eAr0/4fJMMb0v9u7soS9bEr/tq7nt7ByFF1dbNeo8NjIXQzZm/IgCEEU
uu0Xfa16cNnar/beZPakT/FSw3yE/Q6mp9O3wsdqjTYM35VfOJ65bq+ahIRs
rom50a7paZ8jksme44YsqJMiHGZ2CrIA8Ktvbga2wObcY45jFS9ggnlhm/fu
Vg8+4zt70IWm3H8wIHVjeKOvC3e3EB659JbV4XhfIoebZi1KcdXzPZZAhZ4v
fc88OB82SNlNarxCJM6+bitMdrdZyQCPfptDnyaCIFhuGSjSFkUckUe00Jzy
tg27Gl9XNY6tVnVbzkdEwbZaiwvmlwjtlhnYmAPoJ4bMPjJ1Lvs24rNak0N3
QEaFHVLXmVlZmPJz2bXKipoS6Tb0ipTkvrP949F8HqHg+oVDTtA4DNjZAFSU
UDQFvsZLY5PBadRyN9Mur4V24uuq1xMB9KYIjKE5Ac9nqHoFm7a1yANYrPgC
r7m5qz41leSFB8JOHUffFbfRphrSCuc7sGUE+o+d30CyzQeotCBAKKy6xGXQ
uAz06dkedWEOr5VS+GTSKGPMhIHInJtXVdp8vm1jw8L71kvunbm3kDueTsRj
CEXoUrg4YE3elUYwKbxYzPpmgf/zWeOZVtT9FCtz1AxW/PNNHSoNejWRWCTu
7vfD11nQacdWHOOBaeP7ncT/OSdvwXsuKJz/e0cR65gc6Plqps7FhfiKlCdw
4yqopRhEXO/P3WvK2RxZe3wIZbJFgun8YLEHfTBH+ICOP7TSIpdlSqnqcXCu
Ewz3uDwgSLdXcxpu0Sk2vDQtuSFZv9rOSJ4WXx5w/uS5WDTzHikcM5eibgQR
W4+7A5sIIiWtqQlbFUMPl67fiUVr60LcW3HNjdXlX/oQUpBdp1onSNr9kOBJ
Zxihx2Y+nFzM9IpHipsKwwUBr5tm0lEG8FrvalgkUGhTod3KZmEbJWJumPMF
CHtW5d8fUHw+tt/0p1SaSxGV1k7/K+4YnKqscxSBqJqekZ5A5uD6gvUlmkqP
wwMrw30cascqlb7goIriHf586i8B5/JL8L8mM8SoiiK3doOsYawmNK9FIP1Y
QodcYAWc1HdKzoHrGyApk4e7cHrq6tLXXb9bczWtw+P72mZLINjRWFT3cGth
v/SMpE0rA3jL3oC/bd1t3CQ9NcebYTjAzmMQ2jF3+nS+W6IOInHaAjREiGVz
oAVfHJSuWqVYkx/qcEvrkBd1nOJcFa+LcKtBcjZwukpeoZVQUgdKNrmn3H12
XG+TB6keYn+6c2jTN/f3V9YqwlptDuw2l50cNnMt+jjDH4oQ+2e3HCheuGAB
DrJeaNj5kCpR16dDivQ7aYhOjXdwLfUJX4Zjkyxr5Rswk+GU8gEOUb4YsPd1
yrMtJYCa/cX8wWDx6y7ZK6yQ4KwS2Nr0MOs0yxl02GL/jHKVi++Si/1KS4Ev
revHrZqo88S6HQAqm7sPdFWWQ6kTuZbxUOxkuOTkzeTZSP4sZklDGuspAfNw
DFdE6IIeWAE37wXwupwNApb0nh1xyL7iYkHKbhxqvxCTZMcEbvimJXMR+uOq
VxNXO7nZHVmVxfKpjlxImsf4HUFhHBNbXS7tUKHI9Us5vkfDz1G+pZsTPHXa
L5eoqJVkeiGoAbaG753oWjbhpMC8x96Re24bU0+rVhZ/IjQaL07imLWmidjV
RAoinvbJ21m4y0sYIlEou3MIs47OgfJk/QfKNo15ibmoLICpib4r/xNar1Pa
44j3CIBT/d23m4w5eTCePX5NeGAYySxfFrvGaVLpK7Ccyw35wCgPI5H9XklX
t5HjTe1Oxy68Yf9a+VVbAG/iajOXNqtsO03iF2rhSbvD48wrwbA1fIHoBOrV
h3SlKvvBdOm+1dewRLHZPJephwtkskCEoZ2oOZPJgRfqp4lmrULMUV7PshUX
qjiJ9nLaFzM04+jw4h95JlpgjicnBrZzpUYFS1QH5PEJqb7GEAPiI1NyPqNl
MeIxBGsrGhA0w7tVGW4+q2lUNj2sJDjY6I4VEyCvhFea4+haMDXKwl3hk/FH
83sgN0uejx3hWpCusz7HLl4T7BC1+HH+kBdc1cMhtmWZP3t2ujYCxf2nnoUr
ULTuAKEqg8bmm4pv7ncXymOV82slI32wqNBGpgEz99vl6kogtiOUFmm4gxZu
zAJTpiOdY2ZCUwPqzL04VilCZwkzp6kSQKeBcPjz7/5kW+MeOtr6d3pKyjHs
+fMIgcHwM5JUujp8ChIsfQRKkCkmqEtFL00CO6rpcujJLbvT8mQ3795FtG1K
ucxS/ZAOGRs/gJAyYVW6kCVo/Mk/FH9ifsvmEq+nUsySIrqdjgVy+fdn4H+M
2IFiwiWhvurikO20l6l5EEUkcbUGgdhFzH5Hplt0uNFyJLB/q/VWnmx1lhqA
z7ysfCFIQBsobU7w2g8hmPyZlOrl/gjGF4HbRmlbA34DSSV/PCcyDzy1b9D9
NzxDYIIXvImQ77umOeQ6QQksMjKqPN2v4irHwUC1XIlyQtoRI1muRWDFWDzz
QeR3ZMy8YqeGjvfvSnpm3AKW1qtpfcYkF3SxWlv28eINKyMWlEieviPtTyGT
YNBwsBAm/uaaQ7QSb0VzRWZyzIpNt4M8akByN0nRvJxEN3npaOGqF20Ly5U+
FZ9Nxn9vFmHxw2neVwma/wVtyXSfIBjkAZg+GXmpjVf7aWBsf4h0YlJ90YNp
PVnUCemawjmKKFFMINquXePd0XG2quJYy1Jk05PIvDTn6w/5CVpmo2t5cEbd
n1J4sCQMayXGrEjiTkH1FKyNO+TTYfkE3aG4iHYQ9JZujymddx+wi1a1kcR5
XeAG8td0MiqRRqo5JjvcLHWzoYd3rxwwFo94rZPrsAasWcpRL6l/HHGnONq9
ZUoBaopTdZNjbfhzIoS+824Vt/hJ0UXEJjk0O3856c1DNpoQwckOeaYaWEvj
XK0avIct0Xm3i4lBxJ5+j4GA2+z6CiSJi7GpzUTBZwIN5zjkp1RYOQtXQDDp
88tAGnNeO4I9z47KN2HimtkYGSNZnOWD6L1CMJLwOhqGeLzz472H9Xldlnpj
FhGi1ybZpC3InzwZh9ARA+zF5UkMk3mZrPzB+CbEnpHsntghpPOA9P3ARZiL
C+R0Ake7r7JHgaiONl9uF9jsXYfRW63Xyy0va2Elnd3yuNvK1Mnk6GoESBgU
dwnz4J3MsRJOoifRjYXN1oCiIKuQlFg8AKWhFl3zSf4Yq5g0MWfRY7C7XerM
Jz2fJ/2O8t0DUqpLQfZ4PS5SnBJSyoOeeYnfvn10Yn0eDSli2zMIrC92cdh/
DjbKXFjSr8VuNojD9ejgIgQdTikOSZBZSrc0/UOSqV+MaQ3baWYw8ZZFjTqA
1LlaFabb1ovTgu+Z8Q4MTB5uK3D7G8RP5+QTl64KjNv3MWSSUs8k5xfPqPDx
qEfq4phID38ykBr+uGhIcG2VGZ7Dk8lJmMceCKL/tQ+czDXVWXfiY9LsS46N
amUcN5VP4IHjdqkt/q1Mk9o9a4yxZFDW2zjUzLY32YawYKfr0s7xJqvcAd2F
kVxd1wNfm5NDG8OD2yoohlIhZq2vGubLhiomOsKFAluqDC8XDZpoj92AwcaX
ShQ0DIDZSWDux5cSPTDxXVYZUuqemrUzFDr63ISriqloP6xGG4BWwpA50yiP
JFREFWwmZldMSGhVhrFg1xnEF7svekj4AKSuuWaneHt8QnrUI0sq/X/Z6pwp
UujfQ6NTcSXJ1sXaZR26IhRdG+v+CJ8o5HkYtvD+B2Kgj+d3cutUDrUkrJ3z
dxRQymy+OsMjL0vnizUXeUOX3eFSJQF0U8zzG79YfrXx/NU5foadB2kTi/7U
nw+wZVuxFU3P9Mk4gltsYpevLzkZOoLihVHeplBKCG46sY9+yKGZDimtn9Ya
pGwGyfOs8cga8HnVveDZWMtRkA2MKDhUaMMGsOfU/cNtGGGzmcQKwsa2lXAV
43/TtpgL2qZpy62iXc8lg+CxyTBPwt2iVtrdewrWdfTii+36E+NcZ2MyB0Xs
DEKd/FteCunyFtQqF6sQa3fTVp+tMMCYY2RJp+cYwz1V8Ofx/3j0Y7TVLi4i
3rHNEdp3gUf6GhbZA2yH4OaDU2fSL0mRPBGI3PuqIgaMGrIqZk9gIpL3g2L3
ZsSp3HIJp5fvZ6j3qX696jyAlCLoQOR4FJYvNCtl0xXd+izAsQvgxI9RXByu
nRR9sKTikOOe6ijX9dWhWylV/7ZvOWnqEPjUjuK0+0/VSgEufZXtOTvAlLfp
agZ2XsvtTaKQ7vsPeVnSmcbLpnAU+J3cczO0FyqXtrX7pZPbwiVBlY9b4MpF
FrFoUQ/7deW6vQmgxaQrB/rcIFReG8RlVKlyxoUn1V4avc0wi10Cmzd/j2yZ
v7sgL4ewjTJRuzTBBA4+JHKjwVys8i8lmc0pld2ktISbEcUnohEb+bMEXY2S
w8qehd19UWAtyTwsdyfb97RgpcuinauTS83gQGxP1+TJgiO7z/2y5cyfeTYE
Kq6L8291DVTN83GieC6uI6EOvo5N5XwARNvEFMLVcS+GAThUvNd51V82r0CY
SSlIJ4IeALEUAoaMVYVmwQ8qWuRxTx3iBFoqUwmEcU6RHUq1wtBQiQzVWRxn
GQXypDByAAjSh358ascfpuAd7+wuGYviumyijnXSEguKV13ZpONQK7x/fZAp
zGA3+JwPBrTfDUrwBj5lTOXpiE3Fybfnd51QZlDzwjMmk3CAUbcmxgGzxgRn
Ju08jENA2TlAxKjMh9JMWKZ4dBKtWZqYuCKg1qUDTAIKlY95s+THpSITNWx8
NvEy/83L+eXVAbZAUJZ7iPBmhfUmF9r1xpEg+1AH0igRxVquyEkf16VOKdu8
fmw7Jgt2cMdSEjO91TYlO02Yj+tX/m9SVQp77YKsoZpWOZKDTa2HGRpKs13z
r6ksPrHQ1Db22D4cW+s5lUAx650/0xZXLJiAMC3B2bZP4DNdY3AJQ4491ZkG
HebNtu08ZQ0yrttzjzt/OXYbgP+d4OAp09mou6CA0FXC3qiW2Rx8mgTC/Kri
H7z2bg6vKfYH3XAaxaV0pbtYGTQ3KnSMj+bR2d7Zev1La1a9JL/Wy0emH77C
lvFgteOMAFA+pWhxdowfAsKhTfTf0fLe4XWhLeg5jUk6LLk/6NIH0gV4/pVj
psSbfwwTvSHaqlVJc/M8OhgYgdB1Lcs7/uI8wfvmW8YC7z0ntrtRO4APOQZX
kFzG0rAHs6YqqbEVrezF9v+np+FHAlU48TZzs5NLhgBQdWiKehNPZ1nkxJqU
osK95MYjZhxkAibyIcuvczXWC+zTdF+3xqKzYfXFCq8iBU2RpUwEh5Rg++O8
v/awzOAHmVn+zMR1t4WHkd7XTt/6lzRYNLBd5h2RGYBAqnyxa/FRke7on3/z
uTwAb+3ZRfSkd6iaYeDQ7BoWVa/RPRrPbEqrQlwaR8nuB4JdrgueooAsy5mb
gS2OFW9FVPy+GeZG1dndBYmp9bt7AZR9Btj8YCTziaNI8xXf6jnwldSi2mt/
xag6TZlvhEw8dGYtuccYjB44HcE2Ne1TfqAUkOzhDT4N9sHhRs8aO4d3tWb4
WToZTs7HtgkiOGbXycUZ8rYb+0F3Qad7rsqWGlLLDiZeWGF2zKs3mR7qwzHQ
hxtziAHaT3Xh1u88P9NF6JZaq/EmH6VJI/hirfHMqdVWWTNbIL2A3i8WvoPV
zvLBRNbygJbwi1k50UyHUY5Qw8u/d38itAOAMznzoIqPJWj8e0dc6oly7drv
C9m1n6W68HChYYw+fC8o6Bo8lSs9g4yBBLEbtXHxoJ3183SrRHoUVCG+QSan
MbYezlFcpIPlQ86oYh/JbSeqg4ivtpUxnoJtoZZ3A+iCsimBH59zMEo0pFuw
XLoNuMneM5/HOYV3DC8dtlkcyREmL4AxuSF2qgZENkqGVBc8ZKPRx5Icfj2v
xCEDK3PS1Z/nuzotoPtfL3qcr4/+PK5CUEMapgZukpWaqRB4kb0u47UzVPAu
w2hPzNhPF/ggQM29/GdSO5QBaWv+k2lTMjVBgQpxJF5bszkFeDTi3M4RmSFY
I43/t98rgFZe6V17rcUnREu/WYoWBCQa+LMPgwRTuCu5ac+hosOaw1WePz5G
m9c/M+C83jQa+zPw1kefBxxyyGPfjb0yQzgX9z2G01EP2fITHwPtx5MeS8oc
7rniZymubpEdknW3RD2RoU+c52w/fhalTnjtgCac1wsRrpw95VmPOszaU2N3
6RYD1lrp7aptYgJOKRFqeNel6qfoSzOL4AT9VBKpQqb6pGoClhAooR7zxlMp
BdFUHOOWRU3GEYRnSYLXhQnSR5H6ZQ7wbLPnEL1vJNMLh/QG6lufLRH6GvZ3
R/CnihWR2gxyecwZMBD6oNBT4HSKM5V0x3qOLzLplvCqRmNY+SNZHUBVr3Pe
5mceBF+K9OZn9giVc0Z8Qy3azhHHxZk15egAbk5WVEAEp8CHs4TaJFLBNKem
07Dgcr1MK7SerpRwY9ggn/c4NPGfKBG6RRle/XH2iUyEK1fMq6KO/GAvBPmf
v7/emUtMU+bE7nud813ioupPF5O5nJd3kttWe4qjuTLf3iaoLid48taKX7w9
MxHxnr+KQ+EPGr5KUN6eoJKxknx5IpVUiIMzl3Co4fBtvgpUI3xfNjvBJ6fH
UjWgG0B0YFQMAxo1/7X3HRA5Eo8a/RGaw6hhRLara1HlH6NHWgpFq8Itik9/
h3l5aSJnPzd6gzN1oMYlLAksHSGkZub3WAwRYyPSlTbo2TcDyVoES2GxsDly
ari5xOzieXsEu2kv1dgoI0DXj2VNgJVoe0svomkhss2clqankIZQMakFShWT
9jQLm7MPbhDTxEuFnq9/r+sjTSfyuRmgrOeL0gbuLt67mruBtACUBQNLiUYX
JwWeoKktIg7TJxjNMNYn1xXHWA+e7hRyKzWE2JsorDoUXHRZMCCmRbmujFDQ
ihTrK/Rakyb8G7fXvVYvqfOEdK69TIxVJvFcI2P9QZKlc7GOqlfC0oZbvoCi
eDSPVpOwyvUmiEUJUH6gG6l/ecJbX9RW1BTsT/d31MwMvYvm7AkjiHRZWilx
v+994mr/7W8DJO7tODbEhJm1L98ahkFkI4AhZAoNTIc6SGIEZGJctZFA/A5m
T39hDndTPdYIlh4h0z3uRdWYeYCyNx/+GIwY19Cb+/fKPYkUVeDu79Fpcani
M5AdEJ34IyKE1JiDRrDhn/Aode1Lm0NOxBvOaHETKSuxLqnB4WBJqXa2kEJl
CRmW4MfUFAatSjXwzk64FYe1EL6H0Oy0TO2r1Ou86vqzX95P0tx+478M1iY3
dnuL6sV4OYhkq5BpmtXBOANTeSVb13Y6NqEyIA0k9wHB2/Wz9bXkvODTLfKT
fyAcOlkVqiEUYcC2yVrvRibkXHX5oA89dEuy67FAYmj1/kSiYj/gsBgCfhj1
A6V7zt+cw35wm3l8F/KokQHd/HWAYFyUhIFbEG6jV1tnAoqdsJLMlb+rWMiI
7Hi3jqcikB3EaFLCXXd4j/nfWRd7R+kcJjjg32akJAwYeGz+NgF+GcPN/ejA
eEitjByibbFMb+x7e9HM7Me/FDkoo7ndZerAhaHtEC414kwkjypLnjoWe9qe
RXxa8zuJyy98uYxcZdvqeg1GC/2VeX7WruBdjOgw643tBkgPL3ljXb3pWZLo
jGHn9JCACUTCu9U8ny0gq1oyHPCPBfKSdn6FCWZvRMBOjvSEpvzIEogCl19e
yz4Zy5ZBbWGgTf+i9eTXLE+zMqmr+8yJpMZoTRumTLUCRDsvuriZCsjTdBtB
+zmxvy/WQ1qKvO/dvOk+naMMMehm5fBzN1fQTg8bwC1fvCtVw0b7Bpe8xokn
Zncg15m6EKXLeWXAcfs+Mtx2rHS3x4qVDfPEQCyEjLE+g1WLn2U2iCsOuK7M
hhcEtcn0CeuynUa23QCf7J4IriBjEQ+qLG+sA75qITAxfpLEuK4bWUlL7M0V
2QXfe01/99i4JijEQSfiV3DGPMpS9B7DWLe+9yFprW9/Ku0QN23qybxwgzxg
WohCOfDqKaxrrFgpyNwM0ID6sIkCeOPA514CPpqKnUqOR5KBbPDJrb8Wi0v5
gfjMWCq1OpuSfVsBPSeMT617xkJaAt/RDblxOra3AsDFVjdZO4LJzEj08lC6
nUR1Y/X7ixYhpgjMSBW/M5/yhwREIvLbYNKlTT/U1W4G5bsCarEfM5kqmrGh
14GkGDPU6QNGHYimTnrQbbcKO9Fy3sxdVynx7LZdyydTpduTw3uXdA6AO3y3
/Y8VaMsHhOYf0SLJgHWRIwtvM8QDx+4yDiOkVnFgHN1sCOIOvFV9W1ciXjV6
ouhFUGsrWrWirTvax8+ZQrbLLquHOih/t/fkfA+74C/mTVU/DD51zm2eONhy
+d6ixsCGkCO0tg7sUu9MX6M/mTAjLuHj6WQG0ilkevST8nhtwdR/hg4V6cTh
RKwrNLfgZ1z7TbmI3QaIM/sH5OBWwZ4yNx0Y/6sndrel50oNS5fKUaTNfAPH
YFTgR9iDwiQYkBmdimuqLo/S0XHLnVPW/MLQhfY67l0LjvJD1bmTMwgs2SM+
oSgZVbIc3awoOMyaeuGqxefdRivWPAYHppMHRn7/sNmUihsYLpxNyqLEXps/
tcYDe3HWabOWIHG2aWEsR/os+8B41f9YVuysb9C7zKwVYrKVBJRnCvsetm+A
VQ5iN91WaDMB/hZFkfDkx+4j8lpuPIEGMxZ4wqWJVAN0dmFcSFkteabScsG4
tmuNc/B/FtVjKw3x6h40cqgr9EETr+onj90umGl2HvRymUYdEXRWKzRAeEGF
28puLBu5arYQ92ZusTstj4RDgRS9nyjUIXuTLYtW4/pH03yZ6WmPPAqX6VWO
l9cpEyYbl5oy5D+DFGLLzAWUvuW3gogbLO0I3pTBksxArDeqQA5cgz/6CQK+
eECe5ZT06/PuXka3b7No+ua7u489++XtcoUw5RqeH//5TGocsh2EoJLQvpdH
E9CUb26RQtb5Ay1BIqZE5iIpqaUPlhrKVqdLBLa8lifWDq/H7z90yvUglhJ0
smpZSaMdhYaYhlKN/rwUFYUJvw52I0VMk9jI+sSQI+aVUw1lEU6zTYOGbAcK
xUGLrWQt34vEwsSVg8C981RCFVXGBlTFe08Xf+6tB45GSnWz+Xn0j0x3tDEI
t0CfIUFHEOPac5O/7VVfnzBbTYKqdtb56w3RuRWCuxlEbq90AA/wdYBUEEes
u0QYAaXPzqXQEgQ/tAXHPY8c89ItxO0H79l/2rUUiuD+v0d0sAo4Iy/N55mD
ROL9abtJvwMPuzSDWWSDiPjy6I0fJwyGUG/M+Sht0NtGbhxdOEvjIZAdhxm5
SInc0v4x5zj7Aml3EZRFJ21XiVbf8+wEz64Qsk649VxCd+1ONzE5lxWb+Ua4
Ii4O29EMZgHTzMhO4jwAKWWrQ6MyxD6sQciXBTYNghRgk1kjHOWq1yDg3Kv1
76C6P+KWgre7lccwq29kyeZeRd49IuP2g7b6z5AJhtQI8fm1cPb41lzbtFrt
4yNOkIktJzsE/5d5Fr3z+fWY6V0mfW2TNrICM0+kirtiDSQ1Qc5+XsH40Vy5
xksaaoOseXNlcSnHqjo/33ATKnDuR/CYH82HreXo+wsLU2NS2y+abXULeEWX
rErn2HMC9DdwX1tPRy6yv2bRT6IrBVMYwlWeBqJ6NjmvdiqYWd2UGT7jKISW
9C1yH4tHtPrA2J969GEjizATIwuYAb133HvRfpqAu7wfsgOkag39DwB7AuwG
KZizEI8wj1rqaMUZthKfhBjBWEkt4mVPdD4YeDSgkaqvbtz2hYkmuQmhzD6V
Byp3H3vNOZyghyhaXk1aaJbmD7SHh6xTEawOpKHqfvBBVz4EtZwjuxGM1f2w
j10jDAfN6tvhi44N4ucvmLllRXSdwWcqYSmY+ROuNqGWHZqPslU6rGMZg4cT
FRcA2BM1II+ha4R0FuDq8t7XmfcfTzJ9ROu5DM/M13Rc+DeuQv4S6sURzB22
YiSLxMR0BJy9igo25XewUzWK65YT04ZaQe9WKWsBJD7o4QFswNLMUBwNKs1P
IWvAb4hDUQcHFiPtUrBtvngIMX8ArTp/mpOyS4ezmJ+vv+RNHzOJ2eIZU3Tr
7qcd0nLYlHEM//3wuYxfYD8qhhTZgiL8yaSdkvEqN9nZl8MXKvXikHo0oc28
ZDs1pU/zTfyilkwnrQwNYaQW2Q+NiymHOqUsbFkaXgN5Suh58LhfQWBayWQY
4SC7+lZqQl/6jeADfsS5X6TyMtM1Dw9o/R/Q/65+aFnylCGzhMG9GjIhjKE3
nCOreDIFSsEmS28I94N2UKcQQReXDLtXOzcF8mcVZqUQr2jvPleaMLU1tnup
Ujr8+DzE5JmDwI/2KLCvDjYYdgxWcEd/VR6H6a+tAbhHTmRFLL9GrdljbJHd
SqzN5iymIerkRuMW0lW+gOOpjkmP9+Xx+juJBHcNqaF6ab0gBN0SAoUq0bh0
ne3EL7OVriJltk+VNCIQBJZnOXvRJwDtwC2MroTMqKhgo2IJDXR1lrONZlGI
Ay0In20KEGkEwrS9sy+MwNKd5+X8EVUKENURiVUSx/BZs0Q4wac3eUlJhr9i
e8puXhqQ4wJRlmjiaq7pA8zQFpP1Lal6fYKnmrwRDKzPCRNANk/mbBpbUPu9
0HOmf4dFW1lsRF1CtS8Hq3rdNUI8C7yrzTzKWJ02j8LQiGrWreDH0HNcCXjj
uMHlmZaj5Jd2cjw2QcBKNMRbvTPNxdvkFbU36OaC/yGQdPHiWXVwnKkD51u2
hSazNL2swaJMD6kYFR8avz9AnghUzSYntgp+B2LlCymtETg6ycO0TB0/l9Pu
+mm6H/G4Ula/9pCpiDFsbQReQOORjCjZjml72bo51YzyylDOIQIIS1R4KH2n
wEQd+55KfWv1BIetazgA22NmU99tgSDKA+MEp2c2s/LVxBGHY/2wiVMAcA+9
mToMqxCsYhYx3j0SV74XWKXVE/T8a/XK+GZtgU7UhQqZEfuWts61oNu3h2mS
r2oamFpU5AlTArAe9Wq3TMp7Jox0JthROXilTbkAH40PAsBj88kAwq6+0g0Z
Rp+RchA/1Xb8Km7TS6ypxsipbPhwcK/jbZQxaX1rlLi+bOX6gnSSeYkKD3Pr
Zzfu2xdPu5+CKoH+HW/rOEQ2vFiBpLWaSyI661+SU70jOPWPM5RR75sJsqwf
46iobYMk4Rye8HliRA93vSHk/NDUNp2N2mzYmkO5liXQdUeKqirYXjVIBJCp
u5RQBjSIRPhoxxdLweiRjyxUicobSsQ7eYo6XSETfyLNoCifLdav4/y8tCHU
TgG+q2xx4bebxYqhqb2M+Uz/5ekQIb4MS9rM4K7iLqCn/0D1esvc/bL5hn9a
oIwQIZdzKrS4B1Gj0mtNzi6oGQv5zvpJwgaqJmGqyHmiOMpxPuxu8ssPLuFP
Wuelx0tGHe+cCmaLRe0KcxfDuoUTd+2qvkGEtTnn8jazV8+RsQgs0w6iBn8+
4xhWwrVX+HAj5I1SbBBMTIfBEOGK1h6+Ul/XRvaV81Zs7Y75hxLgeTBGuAdc
MqCnWRga/OYN/cmXxkvApGvRMKgpIat55zKPpWsbrE2rRRDy8XbSwCmGNuBN
jBGmq5Pvr7s5tEUDMkeW9vCg6Ulq8IGKF3arUXFbl/FVBKQo3OhLU824IgZn
P8Fwmb4GS3F1RcjenOkFks0CjFGKqaci6tNFk4iPsiU9EbFOVkosbAIeCyAD
Aqjo4VNHv6tDWBMv6B946MlqLzYFs7ys+lWTtJXp5DEzKl0h1ArdrancpWgx
Mxy9loxwOWlhqjVGZK7JI37QGFdn57QhjPhy38NaNesslLxuABAqTm1JDsKl
icsxUrLg98jiEr1Z82ykHaOWUmiRwIm00vEZx8PF6JEbJ61SvlSPqdgcvpta
a286YUvzFDt5PU7vrmJwkFdRIO4mnzrTvsjCU/90J+3HkGTVvCdKe8JXXiSB
DP34VjiuDQSSmCn+997w2avzd1uTCmdNu354G+o7cTqPn5HDj3fPFFedXTG6
qIRx0n5Zo9YVuBLD5d3nsJa2qB8J8j2rUpcbOni/r4j9eXhcx8l7SmfHWudl
v3sS8vm3wE881pFeuusgzw16hqiLbb4bdSbQ3B7kSCVKOxVxWzUKY/1rLg3n
B8QqbfkqeRhX1nf1CcLd7Yv1uHDhlWzriKFVulK0NXsJZ+9S7zKLa0f9mNS7
xvTBriiUvv4ZQuSx6RUrIUYwFUUY13Cr/y3rWNXVEF6/FxTX302dMgz6XSFz
6nU7cn7JD/Bus7e6UULwTGzaWnxdmvAmJYgvmNlN6uFeb/tndme9qugPj9u2
z6PmpxI0ZZ7ED3MvSCxEPV5V5WQ+ZdfHIVEcHJlgcFK8/f8vBliuRmwai/pA
vQnP3y3j1r5oq1G0/cwpszpUcGl4CJDaV5oXHZawBemhNLHFc6V8BAJRwsM3
PkkrsuIxVKnp2X5ouIewPC4TNrAGDrdWGh1wBdb+Mwgw2oZhEuDHe/qbYYCC
2Z6ZhUaUoj9V2wHn57QdjCs6miL30iall0ZBBSiMil6FK/NTVmyvF0CcN1oo
9lirNrq5XAiP8cWacukjZgyvdJkkn6VGHBRrvdraIV7q+LGENy/2HlIKmczI
K4DL5esqgrkKy4xVPsrq383VakGRdITb9Upjgijz1y5jjtcchb0xXmox/Yzk
Aw1EDDA5yaZ0XCHBh9NOpcIMMDjS2ZG4aJDd9P+dmREwi0neKJy3p1znNNJP
x9GHvuASbtgDizQFS3Yi514sPNIrPnAjHe/PVonzIT+vLmOoJQZX5UtEzCpo
gbZDcoSHc8b4MQb0czZGLHeGFrCsvLnP+M2Y9FtWmo/vC3PYO7JGhGsa/BaF
NavF1fgRtdpClTMUPbRpgBOkNr0TRKfg2vHkzZlP3NRCA0+FKVdKaR0IWfai
BqzaqQq5iSVKGZiSDbzbd4Ea7ID9hY0ioXfyFlDFWnZVcq4GC9P9Dh2/FZNs
Sbeu3bE4UVjMwjC1SuSJj1UNszzgjm7EOgg7B6COLCLZn1VPdAZEViXR4lNQ
98W/iTE6OwXDTH2F5eeaj2u1CYF9JRuHy0wlkX3+EohKC/kf26VF0j9HbqBz
XQHBVCqI2t877WMWBnDHHNgrgID4T8AQ3aHM9l4iWSv4iaRMRLqZMJ79gvzU
5JXtKQNRWsedXTla4fGvoC1f042Eh7rAz1H4Nf0hlAiZtkN2WOZxzFjA6wwF
Mo/7l63U9BG9NMG4+yb9vop/qLRRha6E++eBAh3Jn+QqpKrBpOq+CgEvs5gR
3Vlf7mujnH9As1W9LFmu/52URhgFJkNDqcfpIQOrKF1qkDXagbTJLi/lq4R8
m9WM0uNUD4wQepE/BjhTRUC96kjABNb06qKJlZXomWf4SWAOh0GUPxkv43dV
7YlzdXDJ5a/NveLum652Vjr+Nw5e3GMdRAvVjZT0FUEJMFqrtop4zES1wwM5
M7jplR+aOh12lvm5avspzH5J9lGhay8nuNQMUuUftAv7w/JulJ48W4dUsAap
m5WmqCdkna273z1qM6CmTIKb8AtV0El5r4x0KDN1PVYAA0ghxq+XjPc/ua0P
llYCYzcZ5HpXmnwK2wTHcLRLotCwqRtmQUL6v8+27ESV4K3KWaIShQHveYUp
KJhiq0Cuw+xDhHW9ufeG83DcPCz3Z7s830xspytiH6bydx7xQ9ds1T4kKfhl
f5ByJVfaQbLA7TnqSGMVZz4GOJYOK7Chd0FgbzfXuZtlgPuby7blBsI4zye+
4lxDBsxlbXPCYXo4ndvHmS+O7VY8AH2GnBOGCy/5H45MeI3oQ+NMom+rb8Wp
R+xzYNVshKb/0U2sp3BNeC6fFVsNXh2OSbZsCLWpW53E3htlAh7jasLPA4RT
sxSjkUQdNzzVcp+Y6G3PMy9LZVUJTpdSMPHs9APgt263zM4l4ThlNMOOh/ek
Gl/bATFm/BNb6Y3Te4ABD7DuX8AaIo6p5MplYFc92AIWLwDxfw8U18ODsK2t
ds6mJ1kCnJ8EnKjAkwxyA4NmA3V9Fpir982abQwUD7OS/g2kkFoS3Qro3CZL
ZuFEsMh2YUXT2Leg+3vDwxtDsXwxuvX3IHhQiWrZt/LcaH+ilXQNCQ2ZNyNZ
lPJXIOlnGpium+OHCpHjH0xNqV3SRypM5Y+3cIPHogqo98DuWtAZIa0L3rN4
Qyp7o4ktp/O0w4xxbtJsi6NLP5sgnAyOXP14nncbY67x1uv58ShztN8qUjfQ
rZTWlNR1ngx0wK58uymTQ5C3fYLQxv74YF356MoxkEwQ6UA3eBskVaOwBxEa
fog/2Cw6xmEJHgRLJEQVCoS/rdLsfIbdknbWybprgWW8VnTbMhabGcbjL9PP
Drj54z89YcsG/CsidIQOCaDA1ZKx81i4F0hQcO0U30rb1eP5HrG6yyrrUD0E
PEbSp6Em0sf3JD6vIBgjVGmgu/oi3Do7pBWEFP3om6Bcr3f7dLLglHdZtEn9
47YN5zmGlQvtbxFUfioiKYcI3OuOASlOmlNVsFJWAgH4rNDMdGXaBbor4gnh
vP7ZGLE8raWVdbcmUb94G2XYMj1iqwfjD7R46bxpM1U6FDbhCwr6hLTONJ6r
TlKZ3SP0NphpMY1L6IdH6jIGbtYBtSdqtNPKcJVC+3+PGfx6fv8kpusQzcoB
ruill8wmhgjTL3zFRKVPiZ/HdjfBp2PQif+3s3ATTQwKFh6IOl5CG3KxYMKJ
uF2/rTmCjlU30qH3aSyC7GZ+tQ0cRDQPPb9651XMHdY5//yVeKQMcwciRXBu
h9MfgzT6ZX9yjvjQ8Cu/XT/RWyvhs1GXL2vHb3RrRN7FfgbMak5sRbLIChVL
0W5fAGgywQiH3hw6Ixc5bdLoMVDwe6Uw/xtdK8TWBA8TDT9tmyLd1vibfmk6
Tg+sCaGW8Ffcf3JHFcB/z/R5ShTvGrVssCGgZ58eImibHVkTlHVBkpfm0pyJ
sChlyyjdruFTm1G1aFPxNMGc604RaZg8D64RvQIGwdDM3whdnBxnS2zcmRxB
m3KXAolEtvOOIELrnMc7hSytVjAYTCKDllsZaA3ke66Qg6pFwNmrOI4qeqSG
btH7gLKGyA76LB1jfiLTjubKGwXl4KQF+pUhjRteYD9s4Rm7ZjJqJ/ZtEsAL
SGrOiKBLxFA1ylyJvopTGAjhsfWXwOOjM3tnEp/MUjuokVIGb7k1BtyaaE+d
UGMmO/HRgjtrixALFPticPy4hf82nYS1zaXTJM4CFklNOePM1IdlbGN7afDO
YDjjpMc7UgMhdXgwT/p2YZkKmIb5eRm4E9BcuTBQx2eOekyfX/LNUE4JJ2mm
CDpRKK8TP2KiBb58bq5WOLQK5S4ay+lpTEq28F1kfRE2WGFETnj5nDhEBri3
zW6/Hn/AK64S4jdZmM/0N9pELJOUJE6f101Bw9YKLQaqoJjAvh4JCBwDxAQW
7VvvCIhsy4ZQY9eF2HrvRP7yh/Ib/RyBX3DwehsMpGbm0ryRvYXMepbhpxQ9
oab56gmm56/g81BfVcppfxa5RM/F+hbVPOnVJOGhgwzom8YlvjcXQ87ONCCf
CIuHsRxWh4DGr5bDxiI/+ZwvMOGHABAEqRwdSVR1P7DYgS635+Hl4AwvaPTw
R3QbFXNtsS3UXd9PKh2U/BT7uUF226RVyhfp/+SagqnG2GMZGwXnoTxOVRbm
MNavA6Jttl5pnfYoS2yDih9qFyk9fOz6O34iPL+xLbPw8zenq81tFfHgN0f9
L/mEkwHWR3Yb/NEIYsUajfDy8XbD2WmZF2OJyuDLe/YKVV2GrzPbD/dAatw4
Y3OxoCv6CgQxw8wn677zxG3KFCulxIELhLz8yMEydtVG3ozHI2P3BeyBFUyJ
VYvPKCwUsxV38dJFY/sItNRh23fGJoxz7tywkx+WHU53YUchP0oMkdJiF1UC
9nYC39YZYxjLm8JeFG6z4bAWTcaszzi7tojWNyJzLg0lFPSiOUnudh3wZDe8
qXGY3rO7zv9hVGRFWHEyiA3LwpQgrENVq5T3OcNrxJxtPMhv+ZkiF7JXLnP2
TYCXvsod6yRgTeb6b7/iSwBrMkhknXR0qXfgVjE9EkwN/YruoRYcMwhEGZOn
AiVDQ22L0flPq7Y0cMpzNmvfCfbraEWb0tuutLRoBnnBQKnDK175biX+wD5E
/aHFcqm0AkabHxL+Z+cYHi0p9/3aG4Pdc5QIspI8cBcppRgkCNEhRCHcXSRu
DsiP67usttlazsawxovdMSC1TIowFVw6XE9M73Ywtv8FMkubcRGZdVVL14Qb
Tx3Jw+sZFknRBkmDahWqKzJ9+SKqoqrr7131ZOkhKij9y5gJrkPX8DXV8FYU
wCw4yYU1uqOV0l9T4Y+efz9NScpEeqjRNS3JGk+BdV0jWse1hTw4OE+PBHlL
qshYMNiIQiR5jVhs0/cPv3Gh6NCeQW16d7apvekwX2vev/dZCLWCIMbn5FW8
LFD4GsHQq1qTg7VXB6FaXVRbgjZiKMrTBJbmfjsK9Sib3YLCbA6WRL5F13N/
CPqq6IPN0kOCeASdRbu1l7nxuUSzp6Rm6hV45xMEHZSxADUhNV/Q+cNeaUov
FbCTv/rrQ70iYQ6Q2+3il4AWd5h84B9R/5q21r1ws0BbuIH4GBWOB80Osy9V
SZbLyRZmWVHrDNMnz9sjnpYhsncheWN2Yt1JuKEiPzvYJ0gEgYM2KwXB+GWW
QR4eh1cnpr4iYoES2f1sl5p0SQIorsrwdMNhXT4rWlurP6rTBpGQsfXwH+Mv
yVKDYel3Q68qDJaW1U6nlK9qIFjdL3VmxSZkqXOIZW4eHwP/h5Oa+NgN03hI
AI4CFRMQvN0HgbbWZH8B+/zgZKzyjmK6Xyl5ev3XL32V0uTnMZbnqd1gkO4X
7sP1tegi8vYD3FTDYHErJ7WWV//3AtevhaIbOVsuDeLonUFpYKgppHVJ9K2t
Ugih9VF/DUU0iQDaCUjndGVmVgeEidTiNTGJjKCC/O3ZcOZ9nBw1Wl3aaADv
kw/gDdGaIFL+ObBMqNBs8cyvJlHM5RZ4qwQMC+uX8OOOjpgB+cctdoc5YKvb
dZwZHSi0+a7Fk0zOVVZlmsza8rE9P+xU7OBy9nSZ29UhGjkGUJ6ksrMBPwui
BZbMg0fMgTHCw6ZyKDExe/jw1cGD4arYoSZ6Os2Gosij1eyuqWT1Zd7y4sFj
RUS3CBXQOl7ZutTlGUuXVXjFWzP4roreAZoooZkpfmJoiNvEH9j8t9fb25zJ
DzOPJFFv6iOP3Jyc4Iv0wfgnCt6NsrQjB0ocLlOYBDNqTv+xEKPUMAVJChij
JgLcp5R671HfHz94NaSW4CEKyUYiMpZCtEd00arYv0mdCzZL0Xy+O8AduntT
pgtDVlKStm9jzJmO8blWm8Di5C6QqszNpteq8kXE2NZSIrbzApL8AMLUt+Nv
u2PQAdj9YDlZCM2mG0ldwWjIBKw2Kf1tDdQ11lRotPHES6jvELAVyT9Qay85
HcxuB2FITor/zfG5EgE4i/3K89YMTM1f8CRS1T/Yg5rf2HsE241J6U1E2wft
9shK1GGkJE6mMUQPoYr+ynqGDPFY+oGBIO7IiXPj3Qhr1nd6Xf8HImLQCytB
cUG+4nO1h4Le851iNCHo3rMMI7/xAqaZ9mwMIUKCgbphNF+gRJVQVnMF1X/B
NV5b2vpxs2D57e8K5C66Zjgo6/etwSM+d/luSen8jyJugS7WCEl5DciQL6oS
vuxx5hIocCioauX3L1k7jOMyiK23dgU6H9m2zC5/WIZwn6266ZnR6Zs8myC3
W5GaSb7lLb4iGKo/ahV+RjTywukZNHGAmBP6uSlPxPjWDr6NLGr9zO7tEc+n
TkJEW3Bh7GVm3r1vBAhiVfrxgzFGC1j9UYIagX5a3Qoyls72TfZ8/+ACrRtn
pVnSsdlw1eYAk/xlvHv86iOOfhwp8IlZNY3WTvkz9EP1//HtLtLgMGzNg1QZ
1Z3up+J8NT3OlcL4Z6tvV28Bay/iRYUt5kA1T+4Pbeu1drGHYTJ03Mx+NJgM
ABGOsc7hPFH7mOQG7kuys8WfcgmuHZvf0X0A7ilNk3hzNID+JECD5JqfRwxC
L1TXPe7QJ1K3SeleXo3oSTSZ7KwoHOCzNAA7ArzI3zIKeAy3/BdJmDlYOI27
1nOD2lRZs7sSN6303BV/9MqNdo+1rMZ7+QgmqJkN2lBCLytGsRTBhFA876wJ
HhFfEmKHAJYzjbI3EP1xpaaz/rMS1wjlLrsfX2QA5RieY/OtcOJn8JJQugXw
Nv1wCtUXk5zm4A5g89T33bCQ79B6M0IAPmTwE4sw64z4A1R1cpCmhL5vc9QF
EwWILC8zK1d3kvYzAK1ocZF/6TAy9IZrjn6kaieNdnF00EFmOuIXjYhNzcNG
eM0rPkJ2+3oK1ZB9cWQZnGtvRHuiIlce5oVVRM7YYGj/SuVDmD0wWuYSj6np
JMAhviqR4CaIxJN38s5ovl27kfhGG/V72ZX/8xjddK/NJ1HGmIHbI73CR6Gb
EbvW3uHn1avX7GENysFyfQtT6yukTinH9cO7LfulJnil3RXZTNHj/W1+UFo5
fKugH5g4JW4BWcoo3NYO2+YxqF1Yj2QRB9LbO2E8UYOMlbZkYCveNYX7d8Z1
welNfj2PstX0ee4aUj8LA3s4hwNcsZtYYBgPr7MGCTcU8WsUjVc9MeneQaVZ
U95rOvpMfjUSENcUHYQgcyI/mqiQMCd0sBsCe1tmIjmk7pd51kvLkwf0AY3S
III6Uq3xj9Nkp7l55bprlUxxOdZz53TX99XRP+nYIqvvusHnyHNoeBXL4EOe
VNGJszNY/8RxIpXcJVZ7kgDitoUftMD7AS0oGym/WQE3uDrfw00FrAZzhQs/
3qcA5Rc9zL0igXJd0zkjO2Mz34FnPdAU5AZunxQ/DFf2/zHoyC/Z3oWyTF6c
XoAITX3cX6942UCr0jMoUpPwB6lH/Ihask3y5C9oOmayxIUhBgj1v8DsOl7l
68nONi7tb8cjbTKpW4nir1+2hp3VByn29nPY0pqCXTfakNDb59lnMf+MBCbX
DrOixGcB6p44srjK2h1EMzmyNBhv6i2uiB1Zg1bC35g+MKa4/1ootUZYt/6N
pzzdVqQRVAw50KYIEgLRxZYPGBcM8PSy/lBW2Ht/AabbEp4BE032WdKigGCk
Dndq+45zWu2V+lptDddSAp6rQsDH6otBUrekpbxsYJM7ZrZ9Xa76LX7xMYy7
v6jpzmeEFgAoFuCOwSEnMSQQlZv1254POeY0hTzNaJsA3McVx6MbjCJKLy5a
1hog9+h1iuphqvLO20FOBsHfwS2sLoXMdSP+T2YxFtS8qqstq5n2cog7KZXr
TDQZagpLV1ix04ZRT/e3SfHmW0VGsL39oiIKWorLk0K5W76KaHhNOVfddb6B
cVmX9+0wpybC5cJN7ygCshyI1mxY7xIxqOzch1uHvQl2ghRJJvcZBvwSX4Kf
Ba1+gEse20op9pB9c59KreObHy0aMKy66QQAP3sFgaGqYktfmJW3dNRrGCpC
j59NwUp+XTqK/Mc8PXhMlku/dmYRk1yQUF/0NBolNPhCRDDCU32Rdnub9PiP
UloD2+Dco3FoTJxBv3odhlqWSj2Izai4Y7E5NuqLJl5OCcLKWZPNWCXib2l4
PsbUBwK06W+8bO0669zSYF/hVW5KwVfhlyOkqXoEx2+fTpE+xnq03rFzo9km
Fcs/dm8ixySEvu+fmSt3e+XuCaY1WZAaerCp7MQ3GKQHgLM/7AH2Xim/FxSS
J4ZY64xebwIXLqiL5ss34I8G+ZA75Ncfv8EYW/eZhs8IOoSIOC9eQMTam8rb
ZoHpQmPuB5ztNRJk+o1DqAvVSjWWvQSr02FgY7Xaw5ssWymEDHLiPoSaEauw
rya4uzKwlQxuWDZfkkY4GF1GPwfIAlYl+J0xa0wK8oiV/+jArVbHRv/dIWY6
8/UOkWlvZ3p4lcW9nbKNYOBMcMJN62a2S7NOaHBegj6cimkukCwShPL+omri
7Sdy1j9Md3vmx6n/ayZjkYEDqf5/QcdCTGynsVlDeqqOyVwqRSwgSc0qRNNf
vRSryvqHhimICBZWO1bn30o8BeDGPUAu7WaV2cW/dvXjISLhImhafA+jVfp5
Sb4SEJxq2Ey1Gp2viOc+JgI0liuw+RDL+NT2+EUp+HzGPL8kAxoS1m9/3Ywk
gC9e4S63LKbQnL9rCbcFyYPvjF0D0+2LtIPAULJNLTytQ+MV0eYfnGlUVyQA
Nwlov4VoXV+SacrfEa99pzwZwkKwEHSRkUtiSAN6vRHbLLK9sSEikeMkTx/E
GzdV3QOhoRE6HJkDLTeHPsVtfb/UtIoOD9W+Vt1K51VLl19uiauc81AVz6sM
RiJTder8AItcm+zScFkYxQOSoBU2yV8TTCYHqNC+po5qj+GVq+ZiUvAn7Jia
LUgd54G631dfVJu2NRZfaiR+c6SJ4n6l49E53aYy8z8tzx1jGGZFwJ7/OVoY
4EgmKvL6yw21xv58EImrHMCQc9FUJpjcxXNg30FmZMFYsvtX77jOP0guXHrD
LMGO/Ya5509TBfv7Qsk55Ha6FYZ4awPWmm1OG9OLffAmySLK25zr+PAdNEP8
sCrZNEtYJ/2M01abBhyenNMp6lwM/HxtXqiwpzdW7/mJ9WJLURyk51Gj0So0
6pXe+fLeNxRNdMqTdHVXh0KD3iAwHD3/qjxvh0e+K7YiWTMYPH4AU141hukX
KWePZtCdvGToUKgIye6LVicGi2U5H3gEjXYW7y589/sQCFESVY038I0qSFcp
8GNlO35b3uA2TEVSiV6JIMR5VeEHmFwDEm7alNNbL/DLGd9Cmk+5tx2CnRYk
+T1d/+lEIdaDHUoLVJH3EmbN9BnJVuNu8HCH/98QhWTC06oXDR0c85xpYu+8
ZDn0U4/j7ukdtzHHvZMTd2QrPWIuhv8NghhYMmPPoqSH8u5d7iyFFDvlk72a
cFtYXXPcXbCgMWjVdLhvzzM8rs87sL6h8y9PURDS2OX549wgg1RlUasijsms
hFBs7dHXC3/vvNj15+jEgfz2RcsjjDBWaUm8agGBYpD7OsZSb4ALLHKBe9mn
WHZf5XJagt6yYbfK353SMYuR9PF8ozWNYZm0t/dWNj3iA/x0gVhNwD5zQjPe
Z9SoeSG4yL6xfU7whl1Q4d0+7BycK0t1PVYXvHd8wc0OHWvfNub8RwRcLvXI
WmlaKOKxdViGvLiW4JoEFk6FUuYuHEuLUmf1+XEly6DvtN4T7RZooSyhID9b
rxdkjZ2F35Et+sHgUuh+Xh2y6Ro9Wz8MVHpDTp6gNypKfT/H51UAywDKZ3hN
cbOL0L2gpScbC0McugVAA4OKAp/alRrJA85TYYTUHoSzjcWbrW9S6QM1GPcD
t5bR/Wkjl1jwnqBT5MU2rSBZtezjlnQZT0BPWfUap3nJo1u529IH82KWoR97
VTFqcQG1Z/VjqfVixyrnYItEPjk4CKGcGKLGIkMTXna/+5+oSWiIxAIehv/q
Zdpz9tbYqiA+rl9AFXHz5o+LVjcdPKSl4Sk3YhPybU4vl21pJfT1oXiWpudZ
jkH21Ia2cZRk3mWevboS3VYtwYI6FoqPc0ZIpQYNcMHGO3E53qrkhZlVMUHD
KPmSPvE3XmKLUZ/A+t3tN+RQjS18SKAKH6+9TKtP1/Y2DnQ/8KD/t3t5s4oR
CQZf5LXF5elLbWUq9IfrqMEDwXJY/uSLW8mx+aAPeok0ZXkLxbnxzncY0EUN
nkoQIg+RSYOB1algZi2uGyTKdSUnxalAT4UGWTh9r2yU3QlPeknNonLf3qBc
U7V8Chvjnj8SNKnJnmG8XQh1A9cZRt8SxSzHPzWzL1GhRkJwCOsFh3lDi+V7
fE1ljBCwsrS8GmGr8dPfSVn37ztRDA9gzB1Q7Fs0bUuKl3+ZSUWww59/T6Fd
3EU4IaZ3pmacELUFB3sJwm+lsWVkSsUs7ZHAHULMuh11HbIenYYV6QrycYZU
A1G3OxstF2SyMmuBheRYEugDzfftbmsFrG7SuaXkYq6eP+P845Dyne5xyQXT
Dy/BaWDae9Ybk52AxswRDHlkox/zpO7bmJRqo84NHEMRAmhEfditFfqFRymM
T3y8RHfQUDaaEMtuvUXzI88tQ86n5uFzldB6y6pQnGiy+W/X6JWMrUwdtA7k
HRyP1Q/HWb/pDXbZED2SQZFfs+iYD78hsFyE7NRQN0VuY47MEB8I36zmxXop
h/yzISdgwxdca5CAo+Paw9+VmUEWEb0cm2p2gN/5VdLBCKoLz3u6DiQqx0i6
UAZGS8pYTJmKV8E0K5sf//6Ikquwmup7zUjIHLPgG/GOb0Wgwmu1LHyXF59K
Fx42fwTmRqJT/ZmO/mUbx24jqdfRA/h3BLFC1RQsS68W/NRze8vM5nuCoN+L
WnV9/8RG2n28nmWyUYQGcnXZ8f353tmpllwtOl9T2pStVbD9ZHQ5snZckdpL
UyLShce32bfCimGR8rS4iT2SLVU+jLh3bRt4OZPwF8531jT/z6ScMnggukDY
T6cfixxorUsu/ifcX8JVkQRhQH7S6/Lr/qJaq1vZOey90yf1rJ+LvpHDQJSq
CLck6be3PP2VpNkuDxbG3svDYhmcF6rulLwPu5oJ8++eKV5N6PiRB4VXQuzq
TWYHCek6W0vLSzbi5zu/Cz7cuk8fke9TiCdZu+7K0tGZbQ9lwcOwoFEdMoSE
ma0HvRxYG9I7s/kXKn5d1dgzzmasTrGFS9xXzwZwmClMrKzYxjEgy3Yt9tQ3
lpoCjqB23JfNjp3KXCvJID6eDe+Y7aRLNFftOQ2cnjGWXIgYuJMkZKHnJY0I
o6p5FXNXanE8S8pX6b7sJxtZ3+LOLzU7NxXdIlgzM2j4p3uTAPhDaSyi2Hmo
W0myhGx2LSbpeEky8uPFg3ZCOKZC00Ph2KTtycjtMh6GdRyzviBlXaWhAxo5
icmPC2E/Gwkyf+mko6qtigqEXfn8tieniCgEcUPWzkaFI7TQAx4KX/be3XfM
NmGGMMiK8y9eY61TbdgawWIullZ3LxIXmVP7WaC38V6iBaBJD35WaiWcINvl
HxbX0ulOwObUv9Y9VpFDmAs7h9aqxInoRSiEYGP16jQRJHN3DPnWYoyPzHFt
dIKvSH3PskcnEYaann7qHPIXel8A1aqy+mCvPE3tDrDNAjwO96kDasLk+mGO
6rFoi3j+FV12y4eLjLMY7ipiQ8bGaHxdYKk5iutg19mznsmM6O60CcLokHsO
j7zd5kw31n337sKdpN2986KP+pU7vKNZ1t/uasWeXZRf6pageKIE3vXaCjsW
oLhvPNxX15kkiu2kL3sCvvwb8HueHSh12uCP+vhXWRqrbLoy6ZR85zNHs5+x
5bqWzoRYfI/qmR7GRld7nqCDYZp3LztOxhbUhif3Ri0w6r+nYr/2RtSGr5td
hhnNn3Yr0Kgei3cDXkJXXe58PXrgOVdBNnlSIxKu03AgxcnRzPnCGFrbdjRy
Z6v/jGqbRkO774jdQ7KK38ubClN68ekKtLLFE0le9Lx/s5J2E9thCrJPTX63
Do4P8DloPwnJe8uWNKwYC6/+uF7hDAi573MHY1DDf27Is+WcTDILzzidmMRE
VvKSH8bcEmlNis7C9VZBxrjGWOiEAf1pwmRv5xq7bEpG4/2vr2KwN8JiF/U+
JbjDgdWd4bxMSeI8anlS5XM1HWM3Q9XAoWxZgT/o3nyBUlxFLHQxXkMFk3Hz
o81LIVnzTtPzicTGX03YHH3T+CB80i58Rzc92A/GuurrEhMLLy4Ft05ItpPW
tJI3zEiWWb1YYRIDXvqNzsqkR+dd9XF5+dXm2ptma9SXJpf1Yoqn6MdkNjN8
GE7tWVvltQGM3IP11+A1u3tKWMWQVweFQ1U+M/XzSaK1YtFOG52L/u0yHsZo
R13Mcra6WR1LD8rFUXW0nhtUVhTLbbAgOv3U6jfzKvBq3SkCZMa/qNoLjwxZ
LqZkAUVktm6E7xGGE1b5xbI0jC/59w9g9zitU/aL18YLBg59SG7eJZmVUCR3
C9mAZo884ahpIPFt4TjZTpe9OOXYBQSZRmfu29ZLEn6rL4ZnJz2gCMfO7NEG
LWegtR6iCweK3ul65FWUDD9Nd9qmxWCjokcqa/mpD69K/yCMNLEXgE/KZ/Je
4frVu5FoP5HD3Ed70w5jcJCQozpo80SgK+QFbBVxOxRMC4cxLHeo9n10dP+U
pankzLHAlEytdXoHq6ymP6IKIIBLwVw+wUtdtEPKpEFC9s1uZ5zHsGZL4n9I
HshlvhHnqCbv6o297kZ5wjwlLMmbuDzLAYwzaBAQsb9ByBJfVGmWyrZv8fib
b0dPoFxQMfrSzIu9H168ZWEiatmoSQoQFZwaFY9KtyC1nReDbgzowqSjw7qS
vCfK1RqQDCqh4d6wI/oJauQi8vb0c7UCgam/d9RXXxKPTjLefOdKwljHuGa7
a/GNkVSX1Md7aHDPqZRqiDDPXatg2kbFhXJnsLq0/6LRInIx41D3NihvI72c
SusovI8pgsP6sjC404XFu33jSeMg3bkC8R0DQQ7W6bH/rN3f4KPnn+MVm/v6
+8mvhTkG8XyI2M8Lh2RKLlTJnSI1zNxQdDQwyO9YZD9p4v2BARFsMbBzxd2O
buRTupTln+F++BCI2+AN6mVpbrEfUu4R2S+OHwZwK8qIfPsFi7bHgoxZvB2F
Vr/2ebIhFPqkgHZTvA9GWimAnhaaD518j5nhEhBl1UqIG+dcGtxK2B5ELL1q
A7JFXFFCMoDhLPuYum7uPEDTuA1G/+qSlUQ7pB912b8AimhbhSoYWmKPg4Qy
VFjugcXq1aozPa6upuZzED7VUPO/DpAutFSFxq0JVcWULBAPLMJUj5H2i8pj
vxoFyrwmowI16Fbyfijd6lwN0lLFemDDDmEZmfaAzPSLOdaENvmnhhTmvRaQ
GyGQncxbuZxt+0JG3QPLJfRNpcj3QXHR2/N60soDbZDXtP8owz9H0sP0mgdI
VASwgSGBlh6KGMoytpby3+OZbX9hJSAClxAcGOIP2kkmBRPn8ZRjYBWEPWrP
dQdI0+021W+9PBiY1rIlwkHeLpn36sR9GNbY8NsiuI3fk9hrzmEmJo+NcrNz
gmlogyhKvKjC3zwEQU2Wabg6ichj8KztJXeZh5PrxWRx4gXuDb6QbBIZOnNK
Tn28jaj1LAclpryeJzvz1PZFqTSnFj04l/EIpMPMvXJX7S5NsDn8EYfwq0bF
kbrE4QVUdzLe6WfLP9947jD9IsCAmM9vTZDyDvH32VmF6Hz3f5c4/eAW5ouw
tinw5S2jwpDpOiX+IZUwV5mH0TijcAguxx7WEEY7hJ6Xf41AThhGMrKIXhto
9n243y6tuPjrV7PSsnj8u2YWUhEVvcrdxVdRYPG7S0CnTrTOGBkYwerLDmWu
nUUTtxvE2me29iHN2LCNvn3Eg9txu2jS1YSdNP8RQr+FX/a+D/wcU3tN4uTw
oVPYDpQSADK/P71aK7OjCjud0lY/mrrlpEf8OSisBp6HcEdgQJ6gYoQP/vBG
bRGay2s3/JzrF/kdXnZGjHRDkbh2RJ7RsPp6k0tH07qjAvp/QwD3FkSFVK1e
4LmQ6jqdTQDYNSlsYH7nO80hcSM5Byxol+sszLAiU82EchV/cU/PHocULJWm
FOhGKEEZCxBqCyn5TIdFdrLSsjwWEfHcs6/He7+wIvYIR1mLlmV73zNIXjcx
DADwmHsx7xF5PGH6Ao/a6tvFJ6wVPrpVyDornwk09IS244xQeZf1S+Dt8HnO
qJoZDUslfmDKYU9totuf86Hz1vA2r8onnhpRZDt2feIbfH0/leT9CWoAAyob
ye79QYh7/fc3KFjyGwGs3erGHz64cToHWDuvmHYZLPf34l/rAEsr2bQan6yT
MCZJdBzQpPDcXrL4qg+dljdWkXngbmQHPfPM0sIeiXmG27rX+7gxtgq/gGka
eAB08pYekWt+oWysCJuSlGsv+Cu/HEEnMx0hjyEzLCp+kR124altd/mpkq8G
A78ZWyXmc03rvoYuOnORF+nO8ViBqiwgxb5hAhI+dukAf/e48svO/MeozUBt
6QmtxfcT6qyhEGR3JeE2ah2h1Al8Ph0PENRNRQBQaaACddbRykxX6+RzwmSi
rqDWRh5eGgIENrbsi7a/xhjB8RCrj4B2K6Wk708kAH7MoefEq00dqxbiBXnY
Ws12ZZQadydmCWNxBPVrQmJY4TxC2MOv9WaSbGph1Z7PqHXxldddVIcjvr8A
BsMo+0xC6nu0BIbnFmpxvlrfCkZgDVZjXfEA071xdGowOcHi3WVKqBH7TNvY
cVXVqyWuuDb79REduMUFM9R9E5KgXGnpZ3I98zZA7ovMvHJwEvm5la/dXM2w
kr8eNDtx4DyCVtIrTbZI5DDQqlozk4dDtr9uTx0Cnd66CEPeY2GgU6oZbqh3
9O1XVhanLL2uIPwdKymPC2XXjjh/8HvsE+5x1NaAvrOuYTzAjIAs7524PaRb
Rb65EEuBZ+J2p4/gMWBIJxhw4tf0yhi4wkHsZUfQLM7DYG+eOLxfJxEje1SX
/IJ9y7AVXfDGvfD4zosGIRRbPF16ArhBS/iRJJK39LP0eHD6t0XA5SsF7IXx
Ddv81neaPK0FcYoJEin5oUb/+tyggYO5eDg5A3nAdD6F8rTr1XSd9dVIqfbx
n8VzroPeOSfBT+30iF4j7sZxp8FqIwNqKDgj6fPkxFIWeWdQpJDbGs0qpsOj
7suZ6h9NaHNT0BoNtdliRWuwywHCYZJBZPKu1j3yNoY51Mpn8C//+qz5kgjP
IA9bOHqIEggHYiyBTExdHd53BfqWziRNFrySszmOXIru5f6UVgdslfA+X82z
Kfti5ZXNKLCHjV2XReGdHe8DgvwQK9mvNhMyacCUiaPKwHUKjIJPj+Ochk3p
yNV3WqQgPQVO0h+N2wr5uC2M4UzsM/0aT9hxWfDuSpBwDetZ9SuaQI48LZiE
phNWYH5KDtFbjquzkVMbt2Y59KHvUrRnnFGcU3haNbKJhFYwMvTUZIftLRPJ
5SpXOy/9f5nn8QO/KpW5ETbK8VtlB+BpTIAFIk0TVg7gQg9zv03yknwu44Dt
1VRITC+rTBlhC2UUB1BqAsxJrjjxbp3/REIswaqGTCQLmVWh+rbFD3eraWRB
gWmNBHvOQmyjEBSwweDxwn0w/In5/P7S1r7DSq0KUH0D48d90avP7BQrT6To
Uk3lIxKN6tozmaJFm/iYlAWxBHt18FyJJBr9Toc5OUF77VY7kkJS+DjNa2ek
4SrfAYVuxMz+JuY+hTxdPkJ1bxKwbCJzY65TQlIcWNXh8zoDImhY869/iVTW
oFmp2CPu+tIrZro8URzujuVKwOldD62eFD4q3SxW/Ep4A8cCrrL+zISecc6a
6FhnvVvaE2KD7LuX9uz+WJWFO/gGr1u0NQJ8xowERHCreizs/3KHHXQ+pEcl
5eV6f9yOFWN1tXSclBibm+gWE/6k4o9k4Cr+DfKP+T1qJGI3FLcVsfmHpaJC
c6qW8dO6kGRYCs0UylqgBTEPPRuA9LXLTxIDhksvUikjbDHHNExjooja6Ili
Wf+/koE1rmV+97wjSi/u0XLy2dvSjWAxDbwqqnlcMl6UGKnfpdYTBWW7iWtD
/XSX8I/WC3U6rhO6UNWC91flsljDsczVT8cRAsP5yCtP/x0vEGfLe/ydGSpl
fQiN+N5nWqqpdm8knY+og7ytuDgNyY41Re7s/YH1KEl1kkjnAd40HVNV2t/i
CiB/kDGYwWbRMJUOAp66vOMItFKh9lCWnneyta0lqccJMtnl1q4SemZEPDLT
IylZIY5QMuSyxsxIhnXrD/whueGu0PlfZjJ4gTPgvAUlNAZ8BlEJKDs/MjSF
prKMRAso1fzSiLhIUqmn/JztwoTMkR2gUQD29qu4/M078Wwb6WTJGiNrj8nb
vER3zZbxd1ybtbtF9KGbA+4QiGPcPwF02N8F+ZZc9D2Y2AoFWn7JX1j18BMS
5xfZhwhTlPZ0kQDNTH8acfKc9sAGXE6kuu6Qu1hpGO8DRnSx3ATX94ST2fGK
71JZuviYhx5HSh74nIQj21KmsvxFGLCjFI9G2VCt7+4qaBEmM/gD/NfPvFq9
Vgn+LqixCmkFDCPQQIW1p3Y1/vgF9zEPT9VH4HZq6uboAof2vdR5fSYycY8L
5xG9oO78CZpXsXBjnfc0mp9aDLRt87ONE4x6P8trduYHU3qu+8K4oy9jNnrG
mOQF5AWNg3Dc+u+2+rPnbDlM3aL0aweGf2u2JBkH9TELHUCxLuVYDdvxCCgs
cVbnFURxnDHqvAoTMGPOCnLGroK6Rpeptyg930ynItbazjKCZi54df+K8pI+
6kEdWYZh+GFDiGK8GWaLUn2WbkMJQe8K8lgfwzEaIGeuOJlie4EsvHEsuFwZ
pg0oT7JR3wYQW65egColphMf4NBvCJNR9EzMdFeod+3jWKFlrtC1SmdKF0r7
dua1kXV98+fR7FSQ62zf0gWQI63R0iTozw3mQnC2YIg8L7LLgGagpnuKjfZ5
brz0JnJd6P/0u7YrhLfxCaTZgC9itkjeBV3FiVPgfYqxuwflDbl1zuwNhW9C
Pqm5XGO9wVF37JieQBQZsCfw5IB/50iS3NI/vXtSESALO2A59krv/inn75x8
AatusRGJa8M08r9wlnZajnn2HNRTQwblolmhiU1emmg5EyXNqGfDubGpwXpj
c40gs7dxQ2XfygmnW+BSyoKqoBtEFrgCorGPiVqL45ksRAjdkqvLE+dZOCyA
XJv30ePI51C6UISHKG/jjFx4hXzASe4ZXB3iupbgArHNXf+w0POtH0+bEUNn
TAO4alY+R98le5Te8CoARjqDe1MYd791GdSXt8y3K7Z7KogwVcjOmHGw0KCX
N0d3UcPK9F4VlMVEWCvPIzJNcZS/SOtpfKnQ44B7kTsI/BmFJoR1ZxUxhBhJ
AomMVdh57BJxsp7jCdRc1CxrM0tp/y5pENBN6V42MW73m5YgkO3P59dCPq0n
8ZAz/kRa4H4xUgcr2nm2OFiP6XtafmvkI4hypgllHyzGL1id5T0HwOq7HczB
02NRtFKgl5fzBDgYHTVFuD7g+L9dHmmkzTL77G/IOARAJXI+BRWKXXNyCd//
GIvWsDHsYExwhS1DZzoKFyqncepIVEN1AygAlmh191ITilap92g1MNdMDNrO
Y9VRmng45RdAp/NKwXXFS3aYBQKh/xO2sDmSFGxjlZC85XTarSae28msZeE3
nrvZa+iP+kX+fX9Z4EgRxsT0AWZqSjG6D7n9mLuSDBHQJHAUbqY/IdSCbxfy
tyuxeBxcFQN6VUk2ZhmPW0hVF6NsnsvP4DQZZzKdUZke1eJ+MTZqss+kIjCQ
Q870BhtIl36SrH29blRN6aDEtBl8oo2riWTAEMgNrXDFnOAHBhvAObMa4qM8
w0U3ydjRH6rFJF6isjYqtQhd1uGIlbP2oOvZWLvbAaO6ozAELamfkjbZJylj
t2lqhnpthxr/tDJxw3h8GAQN++GXbt1PeoTGbmr6MUeQLA2aHutOIjTJHfJZ
1fma2gJO+zwQ2oLDWJYBqXqmtz9ZxF89YuMPkVIzQkpFCxv5QYavLpzXq4HC
zN53M+ZuBGhrIwU59E3DEq/DKrA0F6ZD7eHBquFe9nt780zxBlDq6/tdojgH
UPMxWrm/3wufuH0xjjKgUkMy1l1xgzdoql3OExhezCW2uRQoIsmDsg/OOAj1
azxObrfluCYRU6BTDIuS6dO83opePeQB4tHS04bPHRD2aQ1sIrCouWftuDrv
55JD4vrDFMhJDNtYnSUTX1XjTbqXxAe3gbcCJHViZBbsqD1KAQgqR43zSZeL
kQcmpvvGmIFA2rXR+ziaWw0+7+TJgMj5RgWnhnHaJVzh8QeVzZpFoYBIBDvx
GYkEf1VBaVTOV3CuBgJ8isU+AxlTTQXwVD5Lklu4mgaKpUc/sY9Z3MHOZ/7N
mv8oTWFwtshHaM2LIF0A8bPHbpQmLCpcflOQFeE4VgL3yF2vsuMwk3zs3cve
w3IBWyHhNk0T/wd8HVkwP1w4gLZSv8w46k0+mjph4YC+EvVKn/yFbSkaZVBM
QCRA/Ss1/42UK3sescql7l4POjYUh4X56rMDFnbkA6KCTLUbjIzcc0Q2Sj6h
ySlHPw2Sd7cFvZD2DwMl74X+czwTtsqlInivoVMQryrISMipU4pntT4wT5pL
NfpwgNjbGI2URkhH4VqgINI6HjtzUfBO5LG+m0YFkaowRe9RjArk6syaIWAr
RZTaZunhDdNuEGaCUxs1yBJgDpda5G3OhBbtF22mJVsps7GuGmm5a6zXrDBG
tv8NMEpGH83rz7rbsjGAfXPzV66JzBptxnn6eijsiqlJ92LNL+EHRMpAoQ0p
vKsEnEU3ktWjjaDO9aGpP6j61nKQMXVwOrBjExMb9XONSgqsl8oAeieaWZfA
Xsjdm1IaPfPCEqWQYkArHNmnxO4dAVP/Pf+erKLjoA/ScjrMKHEE3mzHlYE0
cY9Skm1n5rO6BAe0ED/BrIQguq6VMAEMVJNgfCCyCXJkW8hwYQ9DxHp3mmhl
xxMyPX7bkqiQ8307Dt5IVFzCtMwtGfs5pVRj3YjJeI5YMA27gfA3B0E2KtH9
OXukZl3mNhq87xHJchCB2vRHqPqDstowZ95heWLpxSXjIf/lZdQ5FVppDC26
3xY3Czs17sI9p1A1dVw1JTQI+mSq2fI7GXYiEbEP198pLOSTw/v5MUivFw9w
qR9+py54SfhOzQGYwhOLLwEg1rITLiG1cVkidAKaC4f2ip2ZbpW1nyGALdBP
2Wg2iUxERbMSH3SBclXTN+q8SGtAmK7VSY68CKJYiY8dRkM04i0dPLbZ4iGv
B9H2nWiPlfnMpprj0O9ohnacYOaugYh1G2x/bkggyN953NiWKQbU/d7b4ojA
cJlUqI8s3OUZdMVFPQrhu4hPFwnUavX40zDvMwh3vz829l6leeqmFB+ejxzU
GlRrvN8G6Ms3yBpuJISJdrjU8cy3dQxDz/QYB+C/zaFNf3ueHA9l9wUEjCGo
q61Jfs0moQw2271Awg2KrYs80FTPrJz7q9PM3ev2lHr2oNdHEJsjQ9e7cWsj
D77n/5Yi5F05EOhS4n3TZ56ltrDPqgb1ui1R6ncdhf/eeA5kJVji6LMFssXa
aVKNaf1W9nVroUclIdrycdfuwu4XoAwvLa+L8vQ6tdlcP+jxwpAugHCXXBu7
WSGAa2q7nUp07LzQ4LOL0q4yf5IHC2zcjR+Q2bLpE3gXz/fw2NoTuG3L31Er
v+x+YjIjhEzxhQI+whCHFHmXbLoPvIfzJtdaParLBvs/PhKC7LpL+NxVNPP7
HXahZ2fDeoB8XpPkPkMSMgMP/z9IIWQTG/hfFK7jIiTJC2tTF8L3B8uMuOEj
b24MTAKDB1n9uSNShyQ8NeOivpK3R2fhTdOhihq6Gae6X1liDBYautlnIhjf
6Yh2KBZkmlzTlMxRXlkgcBQ2cZtBoSQEw9yfKKj9V2ZF9fYYiHA0RTC1TQUW
cWG8wO8rdxii209hFPuAEzbk7m/m095g3UVFtIZ3VrL0AA67kxepIB5M/mis
2YNvLljgyNh0PJWVdd2TomFlEDLKwoh7cOfBXaiwO3di+/N5x+8qt4RyzzSA
3kXv1hKiQ/Lsc2XpGgLQjWjtB/WxAW3TmQIvREd2mR6DvHf7T0rxsTxhl+pE
gzcONKWU/2QpUtZzd7dEN3jwDGGTSlal9pw28QPbsr11UVwg94KigPK+Ty1u
ZSJHLcl817NrrVKjLWixUWAAQTxgghmbzEEJPH59xaCZdbnVwWRLFqdhOmbv
A51CdaxIsUcp1vSrRE4lvihghqOOJA4MVgtwry6fzmJXLZsCKZIL60yaBGjd
OJsFYjeVJRaoFmBA5F2YBywiRU75iOTd+xRwwLVZ8cjISfwA86NHFuI6ZBM9
0MdsY0J1cpKaR9F4XfkPk5a5JiPSp6nyiI2m/hCySg3lVfI2gSFUsjUX9Yep
SNVQ5COtSDuamWVNrlYEJOQHdeXWfWIBnzUNr33flYn0lwgakYHUpHpKmpW1
Qtj6ETNO55mu8UePAbJRQ9EzMLJjIsn4uF279M43qI++KFpX/xVV/eevVrXy
71b+mfT3DYCcMd/0ol59t9pd2t16lga3/DMqAyIKS36H0mUfbNQFJVpWmQej
u8EABDTf8wcVju5RdVYbSyNCYqAjcwrL7CDIoFYu/UiKpXjoFjOet2NnQrg9
+PF7gRs/of3BY7MmYWZ2v+d1MPt5aVf1pyiPopWZcAVu8TTdAcTneSHcmcEA
xMExUCxvc2PApYecGJM9jUO6g2umP5HDs20CdqGtAl1dW9mmAuO/p/F2AwHD
gMLqz6bWhD2RCbpGQu7rF5eUo3bvr5IsFohJowo9vWGv5Ayn7RBguoYRNGdM
9ZKORuJalN0sYW8SkhZilWxVTPAN423StvaDcNbMnPWhqxpG2a91zqqwA1ym
Xj5VVmhnTLZMqCQP3eNWWhf1FB3UIdnq0Q0grx/YnIrMdPqeEtEC2qwk5bhQ
9f8SKSdggy7Ju9rogO5SyZErtvZVvzl6F1BKoFwKZcy/Z7fBShsOSrAJQEJ8
tkQqorG9ASL6UNHxaYDzbdpqnTuoEU0IXBSUygh98QdL7FdQ+jb9eGslb6Hv
l8bUVkqM32bV1Ud6mvxsz3rKlDZmL0lO9Jb3uz/+NNz8IQ2fNGwh+be1wTli
wZtLsS0nfVvDdtkFLW61NEFxOY1SvJRRTRFwSqVl/XBH1zUzEAMnLXnyuS6k
JkfIjjpjP/O32LN0B4hQX9SJ90mg1Get8oM5qfNjwjudn1vxtMNX3lxDV5f4
TQMPahvt7NYNZxomU/UlQqAR8UcteY5BZlSqvGNYu3ga8pF1uPvB7VKnAT0M
NH+htDYlN+6f0wQXpgG9kQkdhGMKVhhn9dcxJWuKm3xuaXe0bltOCLD4MIV/
MFRAhva9HmrYuk+4H/z09h9trVuvYg+/A7QvTQD1wc0CEimcslzNWT7h9ko5
XYz9fedP8N0JvJTvnX7yczA1evZ0nL10xlEODKv9UsAHvJEQp6QlPFA4SR09
AUFIelqDacWzTfoPw78o1s+UXyg97yr72fFiffD0fQkrHPn4EZGsUDWbfypz
NwHYbSiCTwf20vLoSpQBcoC2rCOG/ou9mcfyOMIxcT+Uyj/qEgfu9kphDE3T
fokowjO3OB2waC/B2EHg/AFmdLSeo5TowX/loiL3n95eDrvy09JN+4e8Yk7s
XHow3uq6fNrc2poB6WtifCn1yss1XrpJ1SY5i37wrsN5ROA9F1PUl4MxeJ3F
JfNAzkiRU2Qe0GR66eA20DV56i3wnr2zhNUEIwu5TgcnA+KFF0I1fWO/O60K
odb/+L1HgByisubkkPUfQ764fOungOLriMs5p5WbpBeGUPngIACGe+1XZ5hI
/Ds0ssU+ItR3945A1Z1utPujQNZXOjHUtDFYvHLAFb5hX0rcA8ofmIdNm9dL
GoJaTNAVzRT4iHO0U/3J8gCuVlrMkA+y2rZZa5npoyDwJYsp/23/gT5SmAmk
kXJQTkJuRAQ3WVx1wM3x1CJv3sVkx198HFqDTIzz3zm1YXzOdBbJGMH/WShx
7hg5Pzf/c24MHQ0mQ9Nn+YEXIt693h1mvDOOXOzOh9d9rDHbcjtgW86Qkvht
hQ2JXuUsFbyIR5I23E/EjN1WfOlne7XGkdCBnySnoE8EoX1rluVp7qjmt1hL
DqiaT9Ad6JV5ICiPivDxbP1MFtzUsFBHv7X64d0W4+dNAKIrlpQmjDrNnE39
8HkpXaFFOrqMBwbZ9WAmwuxuSGAlZonjwZLdZGCrf7OoTrwhKSmHUZU36ReH
ITq3+lGFGTbVRsAyHzSmswW/RlD7+NwGIpUtRYWVYZateAOn4cmQPF7jaDxE
0ZI1/cGQuTE/oLfdedUBsdTng4J/S9jTcJK2wWUZWMqHBHV7pDvJBEQXEqN4
mj6NUCp+tkvd40m0lw4iG90xipR0uvGe4HEY5nQK92EkgKYUvX9oFZlEi6/q
EFi16+pj/hakV1IghVpr0JGwLLCA3TyuxfPFsdCK1+eajI34sdRv9Gcrum6g
0KuAefC0Kfe1gTUOPSYafLBQH/vvwkziJiCdSZTRQsAliG8jk+wmw7Twrs+u
U1F7k9VV7hJ4pn6A+Xf3IkcAc28N75vxhFNsSIwwDb3sRpTdseQbRhIyLdKz
nd3l2ICRINA5NyTBZH3991GuytiCRLUzLRWrstIRcpDOJFidW9pwmcWLZ95x
ozz1DBYWpnXMP17zMf7kFuM9lmTncn5S3l5EJfV5CASpqFkKK3TWfq5y7frU
NI1zMy1gD/UsTSuj//nAwKIx5xk1uD/mMtKuUByef4aCG3FJMZdMFOEdK3jj
OJ+TV4CGv2PeUBLx7l4N+ZWgZ4OrEYMkcB7Yds0PyWGmCZ0NbUXn9FXKEDZA
Ho9Aff2qoUcLa7JSeDNOXOV5ExRvsXsVpak0mtTetlaiHVhcNCysgM52RXHC
KEOP2KxNdDMt6bfyniGYp145gDKjUkxzNEzMnYuKaeW9y6KDE5+/L/RQfrhM
UC9l3GU2e+Iy8qSlICiNZ10U5zAnZv8W4Mg/Hmybp/PgS2myiFT7MbZVrwtS
ZPnccMPlTi2n5+tk6Ha9UvFrACFgGac0+Qu95REIkCGM8vRmnx1W2ebJnU9O
kSKVJPhO2RK7Ud6aIZONCyguzsIswD7sTXDB3XOVwTUYFPf/d4jpn87QY/xS
4DI5Iynzpf2GkXFHng0Jy/zvvYuR6dIiHpUHuGk1jN4IcDPyvGEcaTZAbemR
bzUo7xioyNiq7CNCMXDs+9o7K0UvZxgR2G6TJJmmpABZonlRUGLgDdpTjLHC
+RWU35m1wmD7aFFAOyABL8j5UWnhAWOYnB24XAGOiCgpugaTUEFHlA++kLrp
PYowcNIZMy+Azwbs3b41hdr2S+RmF5c02nTVe2s+0QIc/p1MYDL9sZ0dml/w
SJ/KoNq1dghAdLFuNLqyIDDWDucafBRbLwqELoHji5aU7Tg1I9v9xgbH0Tvo
G6mFKUJqzxghTvCz7lP3OGh8LlKBCFCiwsjl6zjGDSROz4XITNjHVdoEt0Et
2R4hyokD+hzc/63E+9VIRFrZzsp6PMqMob0iHFmJ6XCEIs/PZ4WACVEkB98D
c+29Lsq3VClALUncAYcF0KZmXwcAFcUOw3I4yUhMH49ra90rQnlkS5T4xxoJ
UO1NI4DPxzJQqRcP4Eb5g8A7ZJ1XTDh03E1+cqDwAl2vsig1cJckuhqOkRHV
krAkBi8huo92vktRtaXoWgpa1TOIHdS7BuOSk+tzr5+eGsFiyqo78omBkIVF
kUDKjQl1u01p/CbbW4nIQzNIwMiW/IMbVssAjooufQ4dk7ptsma2unot1712
cuweOlENrZnAoN5MBp41FiVzLSBkwr6P41BEckE9WNiOI/BElb31CQ2Rpb++
UcwdT3+zjQx/t8CcsvMjo/rtwtyAY7h5/c9wMu/mLv/6hokZMpBnWPzZdy7N
aliLTgQo0QnuERyLDHZ7ISTYcjCICBAEi58pRl9oFIu9tpZal/w03jDc1YA3
8SLbc046I4l2frjTginfcM8XERC4AaNw9pS8UBkHKnBT2xRmKMQmRwNpeFcY
hZflx94WF0MJOfrVdobXWYH6FDE4tna8eabyI47cgmnWkfTf8rF/Ch/YGstT
k0c85MTs9vKtCrrxcujmaw+8j7j223H9X+bnTb+Y6HK7VkFk9Y1Q9qWSuoni
sqZEjMD1ba3Kw1p6nSCx84fU/eibutO54MbfSeYhx++FcrgUmmM5hejF4LW6
HVcfRbSy9HQcTxmBF03iAwBeaFFJVHEHHVOEUq1NFda0mei7Sw6Dq1OA9VIY
qJuGMnahZP3cNth3FNU52yjDutEgJM5+0/RDR566cmNN/1bmshOu9oKbU2kO
mmJSwLwAykjv+1OLyQeQsECikSwlsCR0A5qtiKdzKTWStUzCWxUkgID+vDYs
qzc62Ego5D9fDteKU5rhi8pDhQ6kwAe7dPmq37vslt74xoqD2TYogONR/Fvo
DtCFMSOJKlOQ5XDj4T8AEJ2sYVxrqrQoqgCfgW4Z1827Y07GVyaQ1IOsEkB6
857h9yZJ+P3fAiy3k1KPxRqQt+tvdLheGN6S/P1+EvvgYWHwzzL9cl36oVlX
j1lnBqLmAW5q7OP+ktJO4FgEiAsH8+a61BhoSvdzZpL8Uv1R5ISpkPlpWoWU
Ra0vvxNdFjJnTraVYVN23AmI/1qPCmb28cDEBpWYMyis348cLpyEyOB/wHNK
s0z4m8/3s6l+FZmVowRyGZbrdZ6nRszcsWxBEkfAL94jyqFabzNpX1ApI/S6
B2Sr/QKLEOLOwsUbT7F3oWGh+nN2bskG8ECFI49bGDQsfCrRjvdvHX6GWF65
jr+ZDsAX+/TVp1vBKu/I/5FnPdIs3FI2Hi0Qgxa869n2B7OmZQe7fZNqRask
PSgkS27Ma9S79G+7HZxriw847ErlQTMQgc3qYSyL7cwggo7hCqgFlD1joa4J
Zv48xc9VzLFgwI5jZU9phUT39t1X7FSId71bI+ViEnDyBDCIliywZLAs8yvV
7rdwqPA8e4MVPH5AMHWdIMej8OKz8oOJx1z7IurUIG+608BWjhJzJ8yzoo3G
kMZ3lrnzdI657p31oh94KInqxjjzvFCh+M83qfz6nfg7epH0PVGxZCiCxALA
g41nUBIdzE6iwhAJf5KYoz7afQ/s8EXj2/sYNQy9rKL0hEVqCtH8l/keHuvR
5RuDGd3TG4iQN8e77/nmyjyP2z3iyKcS0mwj71llagz53miNQopsJuFUzhyM
a830sIjfmYBF5PGirtq4ka8Unr+XcBZ+MIss5fiGbBNPi1hvO1m/rvTiRZJz
LTzCTZfbEp8iBxsS3Aw5ltFbUFv78Z8sREiSWmVtKm/sLvBvyA9drLSxse+D
EYKmA2+JcLwt4NmerHZ8uOxZAYPScPx+h9gNmZT0VtDYUZtHMuRKAvii9+fc
PzZtA/dAcESIKIpa5dIChtYALXwClmvNUX7+d/dGY/BwHXQJWyeUSpd41YM3
CL1GspXTdaujnCM2oWBqzSFWt9c2fOyvheJRVZFHpz+hy8Neh0RVGcIGEb/b
t9e660qQoMp7ezrBWijR+3OtTAsaSV6x4K0tuAjDYzLZx60/rdvLGQI/7S9V
GsFjhVOOg39cQigh+SMEVV79HtC3WPqUBTQabtvc2D6tXSuZ8+eSY056sDp2
itngiTtkrKKa9UCfVh9GfVQrvXeKJaoLzEGf5iBMboePvkxblrcT2L+G9cVc
8RE6sklNV4UuyJjAk2CGsPETs8rPJTXBy0Qf82yanC/tJOfLwcMVVFd4CIJA
hCNKZW/7+8sElsVMProqyGe4Pl3kkI5YMDSv/V7EcIr4fc9Pakdd6BTJiR/y
PyEs9mikvCC7ATcfdqq3ONe1yXVec46bbphHtg6il0d10l19g90vtjJXsFfP
7GehWpieUCA4UfD/QH73ZEP1W9KuQyKiOs+C/no8jw0peQS4GPvcTZVCxGfn
Qy7SSn0+fm68L7ZqptiMsDYJAv5UpcDhLeWOjnUbUbugTQzLEkHAoseA5Nfj
FWFFwoDT645hKNlIDqTNl0Ug6Vx8zretH5aQWSltgq8HjsgENDGPbfcTLPIl
o1ElGWMH6h9ZfCzJYEeGv1GN8x9JdXtjb2HmwsFNh2o+ChsodAUznKXgnJZe
O//rE71SM04hXHeSPvZGyPlhsLGdf3qUq/Ln636rXV9bz7omTk8IF2c+eV15
5YaeE2NqSO96zVESZEAikMJRc/aYag/K74HJnISQ+fvycUuVdElNLuDeHPqT
ypCgewfGAszowiHSJtSx69zH3BAb61f79BP9Dqw0yKdrslUTLI3u50tsr7vd
3+37vaVgxYMJUV6ll1CK3oWn5LJitf4oAf8iLbmvuiBdjugm+wzxd4cZA0Ox
Wlvmx4zFQfpFx7M15PBjb2jE5lQFR3nBYe0f9uDBPFT3O6eup4lIi2MDzXzR
8Z5sus231jvLVjqQuNisJtWovHoGiZII/4bs7Rdk5r1jZZ2U6xcQ44FaHn1F
f4KrZJBIeyOXkUpmS+CyB5Il+KfsorzvNnM4Y4g/KoljZPzbmc1mODsjQtlR
A0+sMFxI7AAunv8GjFewNr+SG72OcEv6rLdnRI2SXYXtKPfbfRrri/tRT/cF
avnYmgd/K4CeSMI7gWgaWYyXY2PAYu/pI0e9enPdmkT/8LV7YCRhcG1ljM2S
3mx3EN6ak3Mj/6riqn40ZIAdQ8RUdhiSE3csvngJW8ZeP5Sr6Sq0Ig3o1Y3c
ujkiAs4Q5IgAX7er+XUrgdluFuncMrXSMda39O4GdUmZIjSRDm8pnELWdE5a
tHihMbv6sgWcFvQu2P/eSgzlZJvdwvIgBf25VykK+i6VPhQ5/daewbHRalCX
o4mvX/CNmOPfSAnjxw5VvrHXJvvjCuZWkff6tw3a5g2+ReMx4iurodXyfcoM
3f1vMh8Au2Z1Dpr7I4Xf+vtb5DmkFbNIAre7j0QvVh1MVAB2RCPIoUUU+amj
N6xDO4250+QBS/nNNrrVBtw6Prp7jcX3NMxdaK4YVz0wdL3D28pBJYIjF8wT
0q9qID/t/9uZ7FGZSXPmxihxu+Q7PQCr3SDQ5fIXP+YBWu/FEwHvid9RJ7OU
RPeudqR1ZaYR6Kq8sMgUjJLaowd3oFiiBiHNpNHS3gAvC6UePjyvJoDuVlOj
19yFf2nVxzCe95YanAcjmUt4GotIgP8hly/g7U6B+BGh7yw/l1VNCZxMBM4L
Y3nsfSq/Vopyc0lWXABUtH7bZYSwBUC//VIzZI+JDoxwyeuU4gw4PAT/CVZ5
b1mY5CctavgXR+tCxAbD38CmfbhSfTbZpVbtp6ddA2kXeay1p4vfLarXMXL7
Z9aEKVH2iXJ4v8NpHyD3O4wAI4Vw/E+YdiGXd2k18AaJlvpXYpKcX/RZ/5uj
y153qIUVNqMrFVYE7vdDHkexOj0vw5IHeELKB6KhgxuyDF44+WdGp3s7Jf9e
EYHP5NRLeCS/miDj3ThqOUocF9rs0mYOTSejYJAySoY9+qid+kdacfizk6qe
V9m2rY7zsTzXPgP9XBo8JItHBPZrLJHHGe0hDUzhH9sLBCEqpNNLOM+WmaTH
BTzk5mhMpS92dt3m1pk7ZbD+CmUkK3R4DRjwKfhscTHjhYWRtpUcE9A/xCjm
kh5irjJ3hTL4yKHLCq3d29As8Lc5Zl1dzwE7fDdafoHAEutqM7ySFaxPdKoJ
u2q1OAxyOYsVOfjSKHgtz1jieAiixWzhJ9neDaRs1SIpzlNttzpm5juq6hLe
LRaVgyhhxKz1pjevLOWjMFhEXSejDW/01DFp4awPA3lKCvrCLavrXl7Ws6LL
WepVb7B6hY4OuKzyNzuhuU0si+geChpqNe83TK+8CUVLF2WXjpmZE4zHUnui
eohCnSLCCDhWd0j1yKl7JH1zBvlPu9EJkLgfm/Frexlb93Q6x4Lf7lHkPVhq
y3dHZNpzh4jvQ4TT6g27D1c10gcB2qjqS36aHE+qFpu02T4uNVka/TVCaKl4
icRnGy3iwJEUT6wyEmypVECjA8uHFbkPeAR1yNLPrKQdu+FOIcOVdTxKdOa1
69epL93EUUYevE4rH4JK2bx+FZ+fFXYAInL9xAdZOhfBK7MHHa1srJTvrxhO
KQgxzRBdIGzeLxsJRH5sv8ecHlEqTW1zKn1czmI6nkSyREFAyduVW6tP92W+
A6IILIV+OkkaQWT8PAYE2ET3ZlYU6AuyBTWE3HgAEwDyNmYimhyc60MChk5o
7wDnhKs4p2P6V+FKBAuRm8BD3yKvKh7KRQEhAoX0p058aHO2ybtE/v5loLr2
bLoujzmxZMKwRMLPvW1J1UeorOX2gvf3rwvtLbiOXmTGqlSi4NZvp/nwUcyr
bzDCEz9dzSFxC4/v69nVVyOUDlaTYJxQqZfCt6ALgRe4w2z3DAzAB/ZktHqB
O34m+Vvze1BgOq/PEZ6evr35Q8Oqhgnvuw/vc+/LMgbvmW7sXG07ISFITxFW
AGm9CIk809FLwNkNAHTWkD2RJYxnzrobx4vjtx8hFYmDAwSqCwb04G0cC1Cr
eJUzLMpph8rJ0q+Rnuu2M7LkzJMVn5GC1UeSa3Ybezz2B2XCgOVKdyZ6zIYU
DGEMJCK0XQl92Cm42wPhvR669zF93PiaAgUcLmW8HrOzuwVkiMQSo1CKd08M
J0uI4suzLf2nD5fiQvQZePbYZsSuZQBvTcR02Vl4W0hT+Mk6RSkn8+B0RDHI
ET2jp2A6/UMzRzyjoFglAGW/AYDVntHwBNAOWPict9A3cUm7eRSIRS85pBV1
kdfq+HxUS0ajlTAmOY+sduHVxnd5VU/wk4w54JPg7IwcDmKCqxQ5p66ZQlPD
XR/d55mdWs4ELiwKUNYL94wGTUv7UkATwqGWjyG+zCyDeod5pytPM/bpXN7K
lQfyHU9tyF+YSBsV3MIepG+wzU8Ew9dPozh6+FB/XQj4Tu1xuY/WyyDlRZ2Z
e1CZEaE5ga6639lu9EM2vtGIOY/vdUbsUxQq3qT7XiDOAkp7TMwDnuXBCqKt
pZQtSUtHrb3LaqVhZqoAQNycRDjsmZZ/JNd6r5uE7vyGDG2MHerF3iFhFN01
aBRustAcvLLliL02Xtr8NHa+eUmp4ybKca8jb7XYVhPi6qzG5DzZqr4bxyFg
PUePlrNJtfmaYyGIF9l/ZLca22/12rmq7e3OpeaDbYfz2VF/OvvuOklCtnCq
9CitA/LXvndCnaxuETM48vz/0FEY6vCRQ4E0PrAWPx3bFQInXlLk+Ce+r/gg
qwwrrLkN0vXDLnnjyTYqKI8SNxwtvGXELXy8zh9/CN5wtH6Td3F14YjEwYmh
DEkhnTtxO1BxJhVWs7XIzcr3rr79JmZGssTyQGQL/hNhmub0k9G+n4AjXrGp
o9UOlg5xFiP8pjVCRSERf4r7TeW2ASg/9LxbmGEi90I0iWpW4+NuLCyuKv6x
71dEAIKAaKpqzyOSvMx5Zdm7BRDInI6J9A1TNZrkscWRCAHWyDTHBIC4dHi7
gqm1r/Rb6hjmQQfPvswoyaeK5iV2QhJjbT7iH12U24mRaZmFfRnr0cWdY4Zp
slRNNBl9xm/x6p49rNGFBRtRTz7e9SA+bwHHvCY13dh4wmLIeRJS31UrOPa9
iv9PXln9+fUKzVYGuNfLHhuRDYG8JcrWjd4ii4RSJEhT6DpVyUd5GstcNDDN
aPp4GJo6EkijDzHqmSY3u8CmxCjwaBIIhCdKs+TkWDvOZgGDzTY75uscPigh
yAktcmTB0XDAOLzgTxzz6jdN4Vcll49SwjOZvnQN4vP3IGnq7sD6vxkEjqjO
FsRxDsSWdMkAP6u39WcPUwMVED8pk42WIjClsCVtlHVn/k4HhDzwxlSSVixf
wcRhr0kOxBbLm1X4pNCF7FW85K1gOJ7K4Z/w1JfQZvUmqZwg+2bGAS239lh7
Li5ZY/E3b1nI2gkf0So5t6pfcuNFF/CkB9nvBsTTqxX2WZTdZPR+osdEuhFe
B3uR0RMz2D/g+KnGBfKF085jC6WpUkMWer4sChumAJbjw8Qlw4JIpXfrfcLk
Y6KPWLiIMenUE+uHT/0TWgMZlwcEjjYQ+BQ9pXSnV5WVr5q/cx1djdnpyoQb
FPrIswdb8pUE811dfEQIzWHP05QkXEeCDrSBB529lHEKMHPEOezA2Vi/X8TG
GxKhQW2n/QZqZPDJybe44BlE6dSn5N5gWYFoyrf7AXCiTuxQJOkMGm95eNLE
/ejw+QREs0z8thZN0kVZ23LJqkDqsxutw8XnIvFUUwS5OugQH7T7JHwkedyv
bXjZqKPVfknBYjQD3cRqcFZCLhePfKEYnGFTmm4KfJvhtR9vv9a6J64aA1sB
CEGowTJ4O3fp1WkvRPERYZPMKP/5NnrCkmvzRAXOLTpJvFxtKoq4Z7Sl3O9w
y468fS9K6uqrPagZwIRnrSRsuYU7jD7hbBlXDAG4Xd2nUVkgbd9nIA4Tlj+6
mS3KRYNVsZE1R2DUAw/mVk5Kt+YScPvq5M/FXvvbwai1oB2MUxxgpjItft2O
QRWnPA1kH0umgjMA5tqugCnGbduM1khz5CBDqsqqX6i+z7grkV3gXSe7ump5
Q5uQtBvXdp34E4otSLMUuSWzpaVHDJH1k/j9Q/e8sy+/N7sunySbJkHpnaYA
xL/yjH9O2TKcq3AwYlCRNPlg1kmW9LAFAZEsiJBGAcva+SdA7Sm/vW6YBLoy
x2w2zxuaFZB0ZxkTXMoFhex+RHDXSTXUvo/Yvqfc3vfQhWjGT+DXAS3g2oru
FFmDLiYzM0p3Npfq7cIXqmIJKl7bQ1SY4JxQwtDTzI5fDRrGdpj5gByIpC6H
u4+Icl9MaD2pcm/9+AIAG0qxL6Wu98NKVCJSTJoQKV3pefJEIH1BbN1AMr3L
9oqXWfhme5nUhGb+4ZlXiE/+e7P/oded52URgY+VbHDi/TEboGdzcBXlfc8V
vjJcaLscvToEQ05gY5ElVU+nBMVHmxxT/KoagPfXQf/olK909HjDW91bSXcP
ld1App+fRb9lefSzhzhsJmjXPwLNTw0NnyLRg+/eo+1LsaS8wVcrhKI1uIZT
ctDo3RFH9UYuMlR67tq2PemQMux4v1BDebSo4mXyRSUlldBuEtSK2jLoQrWL
yv4VNhUc/v2uPg4fdf+H3meMFulT57fiwwqes3jUgR5yemf9ODlWA7b9abZV
wMq5AXp1Wf/eKTFft91DN560sbcKzZeQcJYEoqkakZ0S+q2+baRmtkuBUPUK
YeLVlvdp5TMwU3LbaiUE1VrRJNOODEabXTBAuoZX1FkMHA4UIuq6HN1nvMG2
aHB3WClHt+6l3l9Lh4IJpgU/Msy/tGthGxJd/AyWqT+prR5+v7sXbANLfAOd
spaa7V4siwiTPlN+V8NAdQsScjai1nVrDCnusKG+nqI9g8B1j2G9joide8sP
tRQWHPDkl88ScTwwqo8dI+8OSQYvOatFo4oKdwpCjNLKgffO34fQi7rqrrPs
xmkeghL8n4U42JcSbipeQZJX23TcVc6/JF8M3sI5Er+MybX+LcOEQvcVri0/
lJZ4zWuejVEhWwQaB7quJwV7RQuIFoWLXVUySh6ajQRgCxOsGJ5cqlPD1rKW
rS3hp3MmduSyxsvgWJGhCuVii58p6FOHXWBhuNax8aE8EHgkd7t1OYnHaKEq
5tuKFedG5MUWctbhY9dhz0/5abihHdTV2UBgG+iAxJq3yyRSyv2PgFTjGweY
A1bBpGNFCC0GIH71rQYpo00eD8mgw9/R0BciIikURFtDxkjkpF13uvl4gfCV
Nb8g3cySkgUgeNEWLl7PHk9Axg17YhW0jVlhJSqw4FkxP6gazDHL3hrLnG1z
Ws5M80+u5Ekkiz4455Jhr7vwby1TFfd8KgPi6Tzgb2gQ5AfVzn8gLGEo93tc
0x+YQFzYm5yEtVT6oVYPIrMYilqp2b0/ebH4arp7X2GdKP9mnilgJCkM1Bf1
RkSXrm0YtXi0qkZVdyOljAQ7mMxsZpVxjVnIeJnbmcf1XqDk9kHCoG3G7gom
rjJRQHYg4r1jqD5SQafVNfmlfAb0Mk1E36VPAR+XHjcEt69VESSp0PGsD2Cy
XjILtJYqC8qEADqGrojWHo+mW59fsLF1ieGuZzQ2QRxRnFqIj2SZV8aZUHfq
BAFCJFvP2YoK48RrK4bo/nLrEjntBoTiSE4xEDoeV44AdzI1yHihGhr/t/GR
IrRHDoJ0BBikeQkxSWGy7TQd7FvTM35o+XeVtp5dtSguCyHh1snkvD0hD5JQ
/MEOF5WegWoD9Y3sNGPoadh09y0Yp2zNQnP271+jy3xZMejN610l4PY+odxn
2w7JB8aGh0T6IBB0aDrqPifUPITBPyuFBYZFJXiZMem8v6lIaD6qXbRil/7P
Ok9gBXe8gfsKlc+jH6jOIOAhZDtrqWXWZrb1Nf2ac/x5g85QlAHXEcOnV92v
UbV3/PdF8mGHNJqS+IITcxBBMsxU9xX8GdS1I2Zjm/8g64uhAQfdgtxU5Mz3
HuiBbT2h/u4Ksfp8VaRAn8wPd2hUuxx0epW3aXYKvuHgFa28/HptzGQY8p2O
3NDvJTYnq4V77NrNT92j2H809xRw1cDrCoOd5/6Oox7EjHs02guRYZjzK3J6
3WjiMVbqOmt7Vel3f/fgwmWsihkMCJPg+NAF40iywW/96pN6KiEBuvi+dkbG
4VMi0smi87icOT4e3IEPq5elrDxi6dujduJzOznDrwYzMnofcxRvjTeVQbtn
SEXDfVwRbCprjozKr8VV3QnNOa4dvKi6LJ4/okLZwZUSc+Zqs71E2/6htE52
BcpluM2WPPtSI1JUYq0Ncl6PTmVPoPibdJbSiCKrMZEbp6sVIsTLg3RgkuYz
pSq1gi0zt/QClC655SXHjZgMuvGcMYSUWKRbhpNEeiG52MQy+GgupnOud8ti
svA02S6KaQU7gR8kdh64y2kgQLTK/fEVfrL2u4UzM8aevmiPSRAB82hn2kBe
DC0XM6H6ZaUbLXo4flIXhSiwALXgCQjag6Hz9DCByy3cjALPs9PXPjqy07LD
16QszmaOjIe8Ka58//p46DoAAc2GQNQSGr7hhfkMgY/zWhfy1tDvuxaLz0Cu
45DAQ54swqFAxsCxOUpuEKiIgNcLqmq283oyou2+v8hDusLPk8bC/Vy4eLAO
jkfAAPe7CkT8mlmjk1vePNK6Gc115WaFd8iwa2NNWR3BT8au1X9fTkVsxVY4
K41unIttoFwCd4uiMj8a5IuxhVIabiDYDwu+KUuGrNMvDQKBotA8I3n6bChm
0IK+PzvU3k2O0Ek8A2bODioyX/DcR27WP/WtbR8pnjkA+yAPZThsekG75k/M
nNrMrp29bX1gyjRtmQtGEgP/A1a+WxizIzunln+II75+9yiH7eLTd+pgl8Gx
lLnSbUKGZFA89FYFVZSW+/vtOvhF+YJ1sbt2zard8EBZxkj49uQYkCr3kJOG
q6sTn9OFTgP7KQlqeb0LyjjN3nbg8ZeBaTXT+YyFkW+yPGDL0g/ySlksq9zr
iDKsjf4eb9tWkBZ0VZ3OSc9Hb1eZFxKNlO21uw4pnwe0PyxPdZh4erq4NOWd
wse9HuKszc88/KdjS14ymqcGEAcnJox4fdaqgB+Oe2PVd3JNF7onKIOR9hFk
5dost9echcroHla9Sfy6ho5y/pX6a5+nAHXnv0cocOo5KLecuWbKnX3vpHAv
hPehNU++b1SqlAVn9Z0PKg/rHJvXtjIWXjSgnfzygRAkQQmoxRKW9C7YkVzT
9mgIAKvctDlm9y+mO6DOabiwceoSniOcqnDUwuIzdn6EtX0dNtKnUyLdj9Au
VudiHg5slAFnJXVD/oArpNZZ8rUQJY6UYhFvHtE/MvWIkYfx6tCdPPR0ILV5
SjdtkI4Gw2pMw3LBIGFUJnSGWIQ30RGlmbxFpnrE9f18g0dkjIQGHKOY6pDp
MnpOkCPuBqaXBtlKjv+IhoSIgSZDqlc5eeGwHxHQpOSX0JHyzH4pKN7LQsr/
Wm1gqXAUpcMXk4eBckXIkE0vfS7oDiBBMvkndpEcOtDxHmho2QAYUgrDA92n
HkRMwYNpv4KSe7rflpDIrbbDsNjyf0GrsPzIcvZl/gFn7sjB7jwPUGmz0AgV
o3gT8RY1bM1x2w9AwFHoWydvebJ9gmerx81ER4+lWk1qu+7pR/uMGP7oV4XA
XoVw3SlwHSuSy4ddCndJOhLtoTh2Ko2R2oKcrwF7veX+IJG+5sbFUG/4XFHZ
ScIHEaROzvBEZq2zFsH0UilS5oveDKAG72Olbhd5z9Fgnw8ag8ea1DBASBxc
r9j78uifAzU9cnJBJEylDrsL28M3JJvcuzxzhGqql1XfXfalfLSm6mRXpnzm
iF811Q53CSklieKj3J3pqz7bp+RCsif7vcWbOUgs1wJfeEkqp5xjGwuIb6Sg
1Md5/h22t+Xsb4iVo9EoA9yah6UUBrqGFezk+JJfwl2lRGLYq0UrFonjEa4o
MwLdhTMrP19TA7k+2ds8OIGalorSN6cvwnTlKBoQm7zFu52hz33dm041RRlU
RSURAWa5U42s4RpXF20TXzDZ/uvROkZwrLH2DcYxtzogdfLvDsy2sCa2u1HN
nHMeJ/IGu3e+EOJKwTBU9vXh3+qOrLinDVZoKyYEdO3AzSdSdKsLMHB6icFH
MkNgxSj6du9pRWvNrHzB5ISp5AwGtO1tggXJ1Fa6SV9ofI6Y3A+fW3IWtcBZ
uZW+Ioqu/3rw/z8OdbJ4/EiWeRm5ygACdOwoico9W1tX6GLVBmoj4YPOh1mC
lYyxC2fewuDzpIuhqEpPjIm2ya6yZMUqHNyJE1dB0siotauz8sJM5vdxZks1
stUJI7npmm1U4P+tuoduJNhgCNwcrdlXhCUyZIfDW+cBUfo2ukeYn4qSwt8m
Fwh+GrCF9cwTRtq08q/CzfNMwoHHP2D2HcatLIEndISXQyqo9rDKxHA6Lmg3
BWBobrGAukQmVkBuleE6b9JThlDSw0BH4KD5PIys4rOZtDYFwzKAfn8wrmLp
ea/msqan/0kSvAw0KDMeeGj1Pn7m1zamwfJkijTnAeN9kqtnEROSaVBZKZPY
ih1kkxN/6+yoimR+LzEEnxXzum1q49PcWLOx7/7DGWbQxTbTphISOgRM3KXz
Jp2TAN6uchSz3hmIdPckXMi2Gptw06GG8ZpJxKGpYNEHkcIo7KBmwT1Pcfwh
oe6R+WSwln1s/77TFCDiFnqE3snh1j7rtYnv78Mr10xwyNDElhhrzzuDviHL
ttuCXlMKJlR6IhXtTl8QCo4GqrSgIVgnyx0tVWlEPWP6awQ//RdHIdaf6ZLW
bRNo8UFbG2B3UtH+ZHIoIAwzPwpX5tJtepW7gq01Y7EEU3kTj+iTrVOQJtdq
zWmgr6aHUburuUawLLaWoS2WqRCrALxZOL4Y5vg/cIptzlCgescCzV9jOatv
tl/vUlfyHf9ZrLIpWo52UWobrWmhqGzJG3RfA7VzF0olK92yWuHQkWql1O14
2fFqDQulF5uNcYU7EfjDnRgxXgmq7z4V4OfL2Q+BGY26pyBHtYgImtoe36Z2
ZkwA6BC1Xt5Yz8nk5xhu81WWTAVtFVEza8uDL84fMk3VDNS/xgEuDxtx4R62
sQpY4cPf7PBSu4mPWNEdAoDRbl0Gc9wMDh9wNaTHwMEwbvGSFS+QkjTGhHot
6Aan0hT292VE9raKb6DHhnv5I0MsjPR3OV2TOC+lJaYCQkY9iefBIqwg3HJb
xKItPEsJuKn5Y2pQH0ZTWMR2aeuIDSACIGE5fI9p3kWnS+YAEK/umsBjqOKG
h1Qb5PChfOh7vDmMm0kdb8SKIzsWi7othBm0Vmftd/au1r7gJ/tmEnTHKUMT
S1nrhd+/ctW0N16uCs2Uw2tlkxw0XkhstUefBCIfwVCgXQRDpVfTcqaA5Jf4
WwCy2DO+BMZA5ZEhBJSQX94FMNhn/9XhTm4Vlts+wfTjap0CbXSE+brbUFPA
LERu+P1SZ02sP0K1fBw889fZUx4MI9KfvIxaGo0U5cW5KKYCiGuPlsRCHxNu
0MAfM8Ho7cX03UBl0bUhPLXCZRl+o5h0PaasqzBPoIC258eiAs05nH8nPEH+
YpOCEiRtiHm9t/y7Tud48FECe/A3/bPeHdn75Fvj9epnPImplC+67J6xKyPC
HdAzG5Pgw+65U7pOtjryl/LvxsQabg0XPK4zlxU97nfMxMQAqy86VtpOzTy1
sJiZy7Txwemc4tLGTB0dZLo8aqSBKgDAfI8apI7Vy/zk42moumTN4QkFNuBI
F2VOMZkh2Qen0E1SS8xiS2je9Fsec8s+bYa4igez2apjs7l8TK51v9BmAzWN
cuz24TesNDCh+QP8tJa+7bHrI9lkLKnk0DZfWVzCVmtkxuDD+8OMahlZUZG2
KyL8sBJSp+FTNhYF72Tib1BUyEfQhVelZzvi8vMhzDPjoZYfUI1i6GdsbLeB
pAq4nm7Fwvppvt/LdbUgyLw7+qtzzCMc3mDM+sj9ZbDYs7mk2ODx4zVDGuTS
d1dAOdkl14Cnsq2MFQiNSuMLCq3FIr2laI3QhjkvjuKR8lYlASS4y0LwI95E
N6Fdk9MfX24iWi4aVPe2TME+xeEfGSekjBeQ8ifOsUW2X7NyTYpwoRbjunBu
WyvpPDwcR0rcHpNXj0DJfulGMDz2iARx+B5IgmaqDsfIpGpKSp/COBZXXX7f
8n7BuaGS3AsqqlD/nGWGPLb15k1L+dcQ2ilmjuHpBNKrs9C69lZmx0D3HwcZ
/E5RCztJRwk/KYJGnnki/ytzVBGeArFxgEbzBWUqdgTjkfDPpUnZVb12GTka
4UTVd7BQZdYCb6gVM1y4akzIsw1bb4l4KsNaDJyiX/LSu5gs42kAO+0cauhN
AnERiDfe2NtypB/p9tiYVEXUzO7lnT/py/jdD3pUAPJQOxMX74fpg6MVcGMW
+/zLohgiX8xd0ugM6bNPDDN+4m+bARtWzwahrsUZbrLUwpZeMSLE9UC3jq6T
jKSHq0SJsMKVwODnrJHvf6DI21y4rH4SONLNHhA9onwp8NSI4ZR93ZCkUvrd
+23553dAXu6JGZxTH/o8LOadIL7iXEP/SkpxKH42hJ3GrJn+eF66lQpm4fxC
gypgiBZtghhMEZHFPrMez7Zwf0nASxLjsCsHUD8SModoIZtYU/hQBwOYorNl
902uBRJhDPo5ScjOiWIo7+wLexUXzBsvYxOIG7iw9yRc8vpDSsb+0OkuEzlS
iklYAFYPEt2aFuWpzGO7XgokgJrlP5y2FvKRSjVhqKG1QrXat0rlloQfblQ6
BSlZjbkGHQ/lE8MN+21gUGB0mjNuuv71KmFaKHiViu1UgWFUaCE9kBo/yvgo
V7HKipKzRFInjUJNJmDkZrMgXLvURAEm0EhqGzBnjhyw4XH8y+62x7zV0IB5
8V5S4qIadwli2iHi3jTZ6NvNIzks7fZ2drvjRKzMBAKEBnLIo8FQlkIk6E3/
i8dhWVLM6tTh9BCx5Dr4cXChY+/GlY/DnBSc9x/Q8Knf3DGyjAbhFvTuzJWA
yZ/aUtiCX2MW8/CAntTXweqIWH6WlYtZ6Z5Cs2CebVoVNmer/txLsk1LcZaK
JXnXCmWmW/BlE1ip4gjA3E0okzgkfxwf/ag3zYnCpQEysvbGhyFSLH7G2gXP
1gxEd7Ev5yKC/FIMilvHrGgOwWV52K4NKLCwrXHXOvSugRseddKN425xIoVP
kLBlel+Kqx+W/Y0LNk5ImT+cZXul4C/tdaqhmd+hU/IFVbole0/3aaDadqdr
EJQBydZoqTujuTrIiTqMwKIDJKL6LfoSUnk4lZJ1FE6BisYQhgZUni3+g0xf
Hxs9u+ATCMkCqfXKTebyG7UYKD6ef3giGoSlWvFajXAW5A3pPhud1qGMQD7U
sfKMHA87AbdkiWEOhN7RMXPmqyXh9ZgF8J4oqGpVbKa3EBz9cC+0AG/1gQzp
pvMmjZWQ8pxSLlg4uv3KHwHUtgGGZYyvmUuf/pW9Vc8SshsZgEmlmu09hXNs
h8ebZUMDM3EEjjdhvUXmXPLopob2MktHM3KWuAeNXv0iZGsMD6a2cs3L4k30
k1jV9Ck4NP26ghWdWxlZSNYPyG1h6cU999MtNQQCYUk7aHyd5K9sR5G2OgQM
+7nYITu2keynXG08tRzhw+8PBoFvnBYGVspcIuE+p4oJ8z6dZKzL3nORwvbe
CgSr6VsY2GSymrTd4EeCP/UJHTQ1DHiXh4xpkYMfoS4+2rv0IcJv7Ch1+9j7
2SxQpwpqLVs1eC0S1VfEA47cxLcTsm6pNdKMegkEj1dj4bJScr9avqncev8N
wUtbEF2G6ZWFyHFDexTuJCwGbIV6pQWIYouLiPI7C1nwXFG/3lwI5mbXjr9S
rqRVcM8WPv+WMdDcSSXZgXSvpL5Z4BMR6jQncouJ9v5qEF8O51M+QkbojOpU
/TwSWYf7kCZ0VCKgDuMiqFdtKXDXkNqU0u5GJ9dugyHNrk7tCpUAZFIUJSu+
NSCpm/j3gDctJxsl3CpQVXV2o6kUP/h4kG7nh25dCrUuagLi+CnumN03caVo
j9F53/ne7+TQF+ZP3M0hU4DM5iVWtg5N+Bb7L4WUE2MEkU5aOmXRIhrHuoSi
UX5gOQKylrL+xVeM+FH5zPA6e4J/DqbOwPDzw37XxupJaRTzmn4XueNqsCZX
HtuTrrd9K76VWAWAg2b96n6NH6RHbb9g0py/rp+j1I6FEvSZopWyeswgqCEt
+vxOLIUYHEYHh7q8W370eZsGpKqnKZALE3tE/B5tFX59R4vPf7ygaa5VT3Yb
kjnpLVhF+MnVrGm31qWIPqgvSdQN0B0HwkXMxSzDF5LXAJ4uHvne9EFRml/T
L39skPgmvHtGgUM2sLNoIR4vA0rTGPqUBIim8xYKozjMYP2u9Ve0eWtEV7/n
Acq0Z276FU35h4KlS92VIUmskiOwR45qNZmcQXT1bmnoRGcxSYc8aOBEATYO
ecUZSwU8UNr5Qxbs2Ivijc5BRQG1+HBLJAsOE4RH2Vz2LuaXUEHn3bwL1AOP
j06Q5Fi0C0ZuiVQ0oiaoerpFjYMaL8W0GdNgvic4vKjkK1o6MPz8EkGIqHim
fgpsi8JqZ5HFrMIh+fd/M1iKR/3EZB2//3esJrWsUFxCmuAc+H95QuqMcf0G
sGHM6aJVJJw5TCoJ32I8wdBrE5qryBUdwCLv+vaevickOQEcmKNKaFUt5EZX
aBuDTfOdalGlm7iZYeg/x35Cma8KpTb4eG6fg+lLI/x49EXlRsbFLLK+kdk+
xTDcVG3ll+E0TnAW4+1YM5bwjYMxVFO0jhJAVlKcDYM/k/PHyAcTEi0YPj5/
ZEditvcJAXG9a2FrVcTnWso1qSOMcAxXvmDGFkj1Ar23kyWUbeRCB7VfY40N
7YStpm3M9gCXP7SqLE//Oj4paA+V0Fi6rYgpKRfdMag7Ub2OEj2EcgLWem6m
ypLeN4EjLeF2KvQ7eCH+5MQbcnTZGcqV0e3QKuNfsWXyU2NN8JAM4yPsqAMg
gASSF8CpyNHJ72yDaK8UCWEPnzhTMpIW9qXUaftse1YTBVPnfbtrP3r981sz
kX8Uo9KK0Lfv42P2HDybKj24MeCkRwCguuRMYLlUFwhqG1UThmewQf8CSMHy
+mfejpfiFn9E81s8lwE4kaYjCosp7bUqd0CfKhMXzHlhIUJZg3Bqw/aofZFW
sRsPZ2ZQQuI1+nZZVtylYejpckNwGx0mDfAZb4683RUoNFPwKznf+A+BCISU
H/65CWDb7/vUO/DWJyDHq6TwTBX4WXhWgXyBODd4g8eUCU+uZpXRZ8QKvHw1
UHhNhiinsyTxn2v0YsmzfbKJShqYIkEuWAL9Qie8udOjQFqRsIC3Z1d4z1jw
Ybl8u/3vdyRWre4e4wy1e1mk8piw4Fu1KhXuf2sxRbDVxSgcfR2s1VCjeFIB
94RspGlTEO8vyOGxQL5iG/f66blmggttrsa6FaObyeh1sapFW0MadQktrV7w
ieNmR9RJb0RiBKAsAmEPt1DRVrUBLVSqb0jI4HTKJCbrhpGIaiw3YrFvxhnV
GmuP2AgDrqLjE61TeL/WtKdymDZr2wlPmLeqj62/zGM0Xc46WdPEFNzOR2gF
jCheC+PtqIA9ou2chF5Qsgox3LPyJaGll4g/uc7SUFDkgXLJfD9llOGtgXSc
acOQjq5zkVHf0Xnb/NIYFDs7Rkc8sPIqiTRNwDwEZEyx5GYYwyblfucB/ZVS
peldmvOLoIyZsD8cTEU2mHByweMePGKAg9aNUk3sC4fyTB+53w2h5CJY8HmW
2IgVCH2A1Mml8V7AZqI+FOj8RdLDzmjHEF7B4D30cHOO24ZVwSeVXHrrjy5y
J/FsZ888TXzynDr+sIndi/9L1MCfbS/kIKSw2E8BW3PtBUYAfmlT5DHgUqgI
5UELgC5Ob8m0wtuInE+tAY1Zs1YoQi5+lRBPd+Igof1ZdelWONxbfgVPfCkR
6rfCBHswsBiglZt6VzStnpVTbHrbb8hmqDqNGgOKQa99xg199PP3XqdMTpde
n/k75MQPhZgquZBqAWGB8b6komKUvy/Bq4ME01W642D8ckShxYVlK1BrQ2Wk
CuXBytDnvL7Lw7dZfoLuxfxw6DnicYLMD+Wqyr8bt4C7MV8HMt7JAJYAMhsU
ds+pPX6QRgaSMYVTTZ6iH2rmbNNoSuALwIB/me9oTAY+uU6eKTNP8z/825+b
lGeU1oOAcQXRxbTLHPDltz3FJvYHIAOXpqAi21HFboHJLG+sahwTGQSXtWyw
OJy0SVgGCyS/vkNEQ0uvz83gfxZRdf1YW9zcxI7cHvmDNzGTQC5QSjYQjHe9
qgcyFIarQsLE2QwIPESye5yUhza7/2svx/c1urBSTkTY0NEq6Zh3aqNY5whl
iCLeSObwK9nRU9PAjE/O280q0ZkOD4gjsFcg7dHouI7k1ty6SL9X8E/oGydO
G010SSjke0AZF7yrWzo1TO0tNwZyWg/eW8nc9ngRPgXN/eOcqUJOf8cfkPuk
45pq9gDgcV1ThIwjO9ADGlD06YvsnRqv9ZpUUYm9wrF7OHgQ3h1uvOWhpkmR
owr6JyLTQmDdm5IWUQY5W9omsSAyBiC7hJzYdQZuNXJTR2XHpqm1U+Lf/nFq
pY0x37/xV+cbmCc8OkxyP/8KYkhtSLqcK0raUM4guMX3yld0BhNeieIcaB7a
HaK63lWbb7/xxA5jsvE9B2KBd9glX1lPGN6dV328t9Wel8ZlHF902BCcfGce
ZzldR/lcpkxjrZqMyDeRWic6VtL+JE5+ZcPkZfObw/LgBmGGJVfyLcgGp83k
ztfAOzpXMIiPWgHiexC6PhyTeYc00qJdKsN8TOplPJHJiCkmz0vj3sLXP+Bq
IB0jk+35WOSArQVXZRHPbynvSZ4qhuCA19cqE8ax54APS2Qx69dRZK3XKB43
mpnm4NgKNHHBABv6OJqIgb8BJNxGEuFTo44duBWFqfBJmAVSWkfth1eWX7ZZ
iZ27ez2XKYxF2+h+68fYXUr38El5vPdQzIUXB/5VGvzPkIGznRQ2kZ2WXwBT
uJJLS/vT1tfRDb1g7ETSDDK0MC0cRpJIKcCSxnpH02iej35a9Mwha+T/gTXO
lkSSXvsrdEGZ/Phi/jMCqtOG1jvVm7vcv6f1RP5bPwaSZgUhz0hjU4MT9cdh
KKeIPLSfGIjV2i2/HXC4D220BGELzf8eApSkWUHPARiIib+wDO0V12FEmccO
wc/FwUHrU+DcYgc/Zmw1+I5i0MgjGi84SmCds8dkcOBI9giw4t5sB0Q2HslQ
7HJoOqHBoV4XhNY3gTWSRsdCWswM1+6EFtbcXZ1tVHOfWuBkOJ/ptFDKnGvd
6zQ57RLzcFDhYNJ7xdREFU/vg/O9+Vu73IIYW2gbZZ7hNoeD+j5+R7jVFm5T
zvblglBZSPv5XlpDIsRwE9gZxTOQI2ro6c2zoAo7R0y8VwFlqENms5pI0Tro
/ezRLxnWFchtI8tm1j4AAAdDJWmZORP2Ql31xIzxJtOYFaX6mJdLKqJAugVK
hQU03Db/Z5zNXebf1kKt67eAqKfz7WNPiIVXx5/TNs+ZsegfdxGb2QCBr/nP
hH+pQQ+g3UXRDdXUG6SWpz2eWSGtFzxoWePzVPnG6O8j4RRAx036wjFKW/Jr
AfA/lMrIg5JENTPkQv0cuXael7vPUrCVDSppUVrPbSOsb4ZQCecnY5eO0nsj
Ty+5AOaWlkmmkNJGncpwurZsWG1Q+rnI1vdBFCIVTvPbHYsrtyghtT05FV1T
fTrWJSMsHUtZcpLOzzcAVS4XK8d581XVtZ8x6sIpHBv0CZY1xqNrrj84dK+L
Mo0LIzImw9d+TGP7XtpF0usiAGm34avgkl88DVf6EggikI4tG3I5xd1mln/+
njofp1LkK94LeKuf8z28vJ28TxmOcy9/x1vPFVAdIMpIEoxG1igqS+sH6jgK
piIzPMBk1lfoxHcchffA0CNSMuO2ZtrKFKPYJIYCNj7W0aekTr60Ys8MLuvy
nvSwnBzrfESYefV7Imk4yb7eKz4nY78NOM0jS6oIcubF5iO4qK5cdrPmTgN/
vo9bS9mU54VXExiPeEWY33t0ynxMFXiicmEc38oUukvpPxT8bdCNvJelPG/b
IjZNPovNdtRKahZoLL6GXu0SYhk/6Bkp6AwXt3kb00P5Ncsg/VE/v412tmGw
I7sXhEufNwgovSNk940lXc02MGwOl145Lf0VAtJdDcOKDhyBSnRBP2ydWT7e
6jlWxKklS+12dpBocOBZGXknYa02dSLjzvHi6USKza2mr2icaWo+yV9lteWg
oq2gyOXZxmhCJNeMImYOTOL9KtvE/4cg7wI56BttfwVYj2XX4qfkkbge+a7k
f0UK3yIyEIC8GROfxKgtY/VOjAibqH3G7YtikmAEspe9cHmAWXqCPSNZYvT8
aEccC0MBfEBusnGEwdYZ5FnPNj1OHRGymd4MoSBSpM2HQhqnXIuiWTlKwBFe
ROaLQ45omTXkW8qv1aQkSoIdhKrja3+rCC/8WOc/MK7hO11fKIePtyVlaIRZ
uME9259S5ZMry7GCkafc7VHdxc1wd0GzZDb/aqTUAeaKU0WgAUzTMob3vJqU
+RHs5abFERaoz5Ha6vYHDmcdub8Q8rb5MzE/gMvOLjr4QiMvnjni5TUrtp3D
NezTvzDo6fKHTFIUHK6eUW5hsIXc5ewyoBLoUX99LXKemEkOmvUVPGDr3aGX
uRVhQi8XJbE2HgcT5Z+o9t96hLibqBx6YE6XFfymG6eBqhZy8zNaWQaujEOd
DT2ns3l9c8yRffXEVEh6p9hOl9D0vMK3YR6H0PFubx7lt+pEWD72Ca7E9jGS
B8rHqO1B6CTffuTgVbUBt/tgiZ7b0wBXlEGG/cdizHnzbdohEFlB6OsxYUo1
Yu6vVFMoD82vkYGY0L7R+N2GkaqkwR5utP4CmN5rMCOK3nLaizBvFS/qzTsm
DNmIMIKIg9AFysLeFtDr9cmUguidlNharX5rIkdNYIWe3/B5s0OUOk7Puzt2
WkCqLhhCu4yM7pB9ByZwORmEJ6mUU33QKp5bNUWADXu8tlhqtISlw/8m/Aqo
AOzTflmju8wFmnC2rcIUz4qcfgaUG7YJdmIaWNYP32Xbemc/COjYRAj5z3yO
tKZg9JBhtf3gMQjz9DAEoQFl/6OKQFbD/iNUsldWpI2zIYWpGS0dlo5r/yCE
dkYGiHQcB+KRZ+/KTm5FbO7sRXkXhnco7+oDSbz5wO+rzdBJzJRCp5OVif+u
pZzWbjwSnX7Z1hHvkZ2iLHgic5kRkBmDRVm/lvzVJPMGbc1xGnwPo4J52wbQ
n3+BaVNACIh9TDoO4sjagjmPHyb2sSYNgVkW+UipAGrgoA61+0IRBautRnW4
kxbpBRiKB6jBtP00eWX9uwGrKR7nVk0esTFNGT6Og0vJYo6DmACqHbqyoS4d
xoKO+KtNYYCQKiA/PFzJIKeVtWwq8OGzzPCOATIRKkuaKTR/I2TNDqr/EdlD
vyPgp7/6pJ7vgttdKJY7IyTHCMSn5AhfHT1aElJ4V2DrXKKs6OoDcq/BIz4q
m2uAAjcw6UOACz04NwU4zkOdMhNtgh21BaI5+HuEmOqj7h12puexjen5lFYE
iC5Q5d8t3PU/GQozhAhcT/MhxZ706DHYTDvJ2AJooD8QKXhLAZetNM5ZIRNp
UC3WO0+k3CRspGayGLPz8LkbIMd7kPnomF8h9Z/rX5C/vRA81WDXufV7BwGD
bFU5xbdB46wsl+Z00gRP5UISrxYd+YywEyLDunNt431d0UqCOF2OT4kjiKED
ho0YDebApSpULttLBsBGdxwiRKITCkvooJ10HAhDNcwuv2UfHRKNagu9U66s
69SH0JMZJFpexCEinViX+zmb/9ZQXV4RYHnM+RGGr9hHaJiPOcoPc41jMDRa
tjcupD21S9LHkNPDN77wKi841BrzYbVU2jYDXjXfqmUzKPPhBnGqqMxuH8QJ
g2BKAwd8DohWCwn5Riv6y6gdbek9MwyYdrxh2i4mkdgw2p8oY/AO/0wHE95v
55AsaEfnehZ/73+bXMz/dTKTLIwmWNX0ZuUv/ileVZgMRiuqfg39qUOQKqOI
0EamBuWm5ShD1gQB7py8Ux4LPKHhGjjoPeB726gmzXSg0qCHJ8MdKVeAejhG
ijohOxW24+V1z6Z8YLo0xdRVDV4Vc+zzY+Wg09xQ7MJS8pWJrolwr4zCnJ3r
/oN2ddCa/zohbzdFHDXjj9LnowVy4XoHEkIgsOkMWuGqpoy+RTbSAXHGGevi
EeBjJqK38ejOyMKZZFgRxK9bv2ILcn1FuitaonYs/34R3iQLTpA1AV033w8k
7608Y28eZih4GopRUSjS8p/4o98OMH8NS7AE3RVlwdOkscqhy+ml9jWAZwKD
TpsXkzZR3M3y//u6zuteVxyFXJiTTYDrH7dFnPCCwl+0D8ASw1BbdaGHgLQQ
7CT/V1bMnL+TCA44kTrv4g7LpPwkoki+RR3fl/qfEP7dNqLBn7sdeY4nhqu7
IxHFBwSiT0VixQ/DQfbuHlnnHjeoP6WmKTmUUgDvrnDcoAvEmGkn6NxursVS
ZxuG/W+2l+2M4x/Ru66qgJfDcgKINB+d3ZClj/mPWL/j4LMMOw9STq4rJBWE
RcZPrQLW6rf5819PMoQ5K/5XgshD71XlWuRzcaq8hkhryPjVMKPrNeb7LK1K
pxoy6GDFSI5MeZBhlPOGKJyPg2+FnFRnrmVCnHZ0aR8xlNLFx1mRwO9QWSCB
QUV/pCld3RXtIflSvsE0RXSw0W5qK6MGDgcxRyHcS/JFLIq2r0XjK8ubZvIf
q7d+583R2mHWhPV4/gyFrggCNp0v/dw1fwrsJplvGTIPeomE932IQBqFvuVM
3c4nGYkBAU8sbAE7czAUBUaGcU2VfN0sWUfjkTiN/5msntl+9r07Jl9h0REB
Yf8wzhwvXHbpFBaoigOk7I0p+oyMQ7I92gmS0pekhUMeHEzjLfE8q68/YSBz
I+XbJMEdC3VwRHJHkFMPz801TrrRsQaQZVaLjYDeWJsUiqXaS4OPgeaigTTa
4PpFOtfW7CRVk0AHp0Rh/ZZKYpx53nSn8/5Hf+MuJorVUFIjpkbOabzDAA38
BPUyrzWxcnAJnOYnLbVwO6Z0m10smGdmV1OrxLTxnb74JMnGUz5dxQHAOdOV
+a8ceT10ngqQv2LOBFC5a1ts/3SsJp2IGeYZuyLhgaQuDe2PiOdDbzBO4Ew0
oXsKbqyTFHkamQBPz7EYhcwG/GYcbL75GR25Tp+Jwozp4upc/rmCOJIJM/2N
IeMvkFzubzLLH/wPiH8DoO9zC1a5EvUmhP+KJzYkmgyMbsi4SzVQYTqqIsQq
VKt7T6QXh8H+4coyNrL383lVEhAsgGNT+3wBSLNkdJYt/gkMz9xk8RTE9qy9
FFrCJ7I4kYlWA1neuUXaRJSthnmHdN2CWlVF1xmw8QYAxwJhUNB9SLv8nAUA
nEmwpONKhLQEpmHbChtOM/ibosqPcD9x3paktRh689qhzNt9mnImwyhBVDSb
QCeTB7+0UqsEhQH/G5+0hCEwRnngF8OgIDSuFCHDSGMncBtb7gXj7kIq5O4u
6I5v5mRgGkPWT8MJ+nQeZ/DAugEs9q8nzasgqdn52U+w6LGV04RyJCaclLN+
cReFN2dB+9hPnIJiQFx38mHTI3wDdg/P0+br4O/YXsoY/8KbGruO5jCNOMRj
/zhOmGThbQlF+htjVMzOPZqxj+tZEOz/EZXBG6T8Be7z54zIxaXbr7hCFLIc
e36FU6NPvS+pAhyRpCnxXz5TEgXzIxly8HgwWuSlCy5pRwa64Bsgltl136C5
r6HK+dUBEOW2k7UM3tKWSeR9TkpkafQb2ykJVJehwWrtPlXBkgoZBRO6rLhN
h2cP3mX9JkOluC6m1s2NCdTJJhJWLNnsR7y+/YcbW4Izw2PVIHsumCFPivcL
56nr+E92ib6xR4x3VhssDVvHw53X3iFev3a90BF3y41d31gFyq6yHhmSklO2
MoQgiy3EfXJW29tDbYYgK5PDeXlh6f6lbPMaBIgSx3yAbTtj2BQCVqfWVtDq
xkIedysS+NkxgnVgBh97Ws/WHR1jbDjNODN5WzfyIdNDhYY6OC+B0rEHFqnb
gyU2Rkyfa9pUOXdXiJkS9UlgULPGj1yAY4wmAfF51na3BFh6K4sB0stDersA
shPaGdNQ4zEQbTSSizCEN1pgtF0HeMzKu4L7t15xq1Rwb4iAWw+KrhnxPDlR
W90LGbS+euQzpXmgkg7BXhYXEsTCX6sUGZDrY3KkCIIak4gEi0YXSx12fG28
po7Eqqtxpc9piYrNBYSqzvESVTVMt3L6ARpYaeEz75gq7pW2ae6dM9o/9VNE
FhxyuU9nRJEH7k5tp+V9dak768IQxErRa9E1lUVhKFrXuXTgzbz9RCXSh2LC
VExcD45MEbZgIZQc7WN5RwPRcg6m1qAhuLSsBAfY+1TC4h6xWersLiAW688x
Y0sJWsb5HpgwHBiU2moJpgic8BgqsvxkeyeJre/KWi7KW8b4+NI8YMgAR3ay
pMp/RQH6bYGV3CALHbgR+1XL/HYESiJOAs5c59L0xfBrBY6YqxjKr1CrGpDX
+aF4VzVl5/DaNl94ITS3zn0yGAmUhCDmfQJ56e7XaCk6qgxMhuYHRDmD8e6O
6VpmfEdGKjILPgnKP23oCzfZArI4rgTXyChPYp/PpqeqKUnBf6LLLl26wBb9
TWuTRDoR6yt79i4TQioo3aig3WQpkAawkuAz+KftYA6WIJTIqhTebsU+WmqL
cwbpuBXhhMZWGhPlxQTZTUlUY2PzXLwelGkYUQlX3TfutouYsIBnQW3sOMx1
OixGwNJxA3An4cVpOUvKfddGQFA8eGrx3tEIA2dFikYhmcEgl0E/NXvuZ/7i
6by4MTMy5ejN+Z7QIj9ywD8CGV21l7E/myQEq0e2xv5Dp7RU2CPLVmL2jRGa
mNc/J6MKj5rmpSB0ebsN2Loos9WPkUsU7M+xdc+razsgY1YePR5mJN2h7OED
P4aa4mKdeQuewNnSHzhzO1Ldo2yqG86VebdWVO1flSwYYKtA1SShJokuOukB
CihWHAsQhNb/Lpv6aRlSqIqTa/M9dx6P5Eg9T79zYQvd4zgiogtAu3bWIjnJ
K/oF85asBNRWfBYx0PxDcW0T50EALkuF8jsR6SzsHUqboQA+5jIvsFa4AYMP
eaeyi/ZT/PzNVxE4DvFIXZv+zizP1wREZDIvw2WcClEiEc1wn6BkvZLIlSGQ
4uz67alpvY/gtc22JW5ZPXQ2zZXO3uOMy47lIDpsU11QIQvf5bWc7e8UhouS
kNbV7dI+vqSNyLcO2X4pf8wJDfmV92iy2bWZ90wBhfxV+hwQyb0U0xKTXhuU
its+NOp6hYUFYmyQN0Xxg1+C4gx2s5ophX2oUyYhUQh0INHIpH91YD0HBib4
9CydyA/eqqsy0hV+IlR+Xh0f5qz8ARfJRRQ9wxBELucfzdfDn0d/viDIv2oG
hwk1tZ53uELJ4ybn+G7E3MXr0ZqadoiK9ENVf0gn8AkGC7b4MFndqJZN/4vV
vBxp0YucMS10CbjMtOfdjhKqaLnRi8jQuXn9RjkfuvRXKNOkOwSxN6sFGRdm
n2puQRTUa9u0xzQbGi+0cA8dUca2jhwSxQ4HrlAhRx2m48qmMSAQY/leZnkO
QP2ms+bT8vpnFAeUwadMoeecvVVaLm3svW20axSpWJX+WqpDg33ek17ipzNi
1KAJvHBYshfNVe/ry/I1Qz085Y5ZtCID1dbavIG+AGetnhXjCwKl2dhrbrAL
h6fXEwEBIbyxOzxktPEQ2dKGNxBPRLxX43xaOfZb9jiQbWzLLEZrKMKpnXSU
p8UGacDHj+Rb6KCE/8BA4zykukfiberd+M1g+mnFL0iveKuS6Gyx12lj1EtE
L7DqjCormT2PYKmfEdseA/mgk14U766iQ8/hXky4MlNnSbzX3VJnxDbJNNqk
4Ms/14vsmpCHumm0iWhsJWmQ+B2Sy4eDQDwJarjoNSlFLTw0h27sqBXb1J6D
vyr0lc88SnZ12obPdQVa5t9EJB9Gx6k3enLMlmIZNErscCO8dJeZ4Zy+EnxW
4gbX09cGVCc3Nd+NPmTASGiKK0bQctWU6IYe2Z+wVmXjc7og1khtCFC4Q0E9
zrx9YLAiHq31MvPqDvYdI0K3C3RODYjky6G6PyGTnDFiuRG+5AuilhHa7WbR
pT7Y9La/QOKS3SCoFwetXmLCAcnqDBnVHekV9Szz4v6DZm3x+vk8IQtgmQcD
qESrn+PcsoWsoiXOSQx4iCiL7YkeEMjAAx2Ni7CTVLa71ydx/3DH4gNm9isW
dZ0ezAdC4xuYSkeB8U0lkHNLY/UjfPQ7KQW2OXhPL5h1PJumcgP/BD6bLcNL
WMxrgYWKlHOLqaxIy3+2tl0HmeTpn+YOH+suSbG/FEGo5Gz/JPRk6gnXvpWA
d/v0VWw4uJSMUXpcn7BCPxWvZIb/1FMnn5lBF3NcbClEs0AUb8y7OTLekwE8
Dl6oIWfApqygjfJ671+mVLE1tHMqmCEzJzAk2mts7IrB3kcZSlRnJ61Kh9kS
5sg0PHehrev1qRQ7cID8MztsRP9DdT3Bny2w++UY03nczJUGF0p3E6r2IAwo
bGXWUsKdXH8hy68HvbF94zAWoS+emHe0293vTLLx3tNzgouLIwEjM/4In4C7
lT4tQ+CaxoFCivBmWHENmHMyE+IDYs9j7XYYdFgHNc9RPCmwUMSGwhymLLca
5HNC1yBSm8kFnwh1ZzMl1Z2TpjbF7BiLwfa/XzzynJNWDpAOCnFehosgVikx
grYjgB46FJ+2w2sYGWfSbsjNL/HD6iFYGK9h/DSav5+rVVI9OEsV4NP7TTjH
Zz1QL386QurR2fCPzMF1ytUG1h5t9ZxX3ZG+AmxGKhUbQZ683sd2gK5JOEff
J98wuckV16smxXxPgfIe6frw0fq8yDaymmCDSDc7h30Ghtp1UbrWmAm4xj4g
4dV0k88sffb9eag+YwTzvq5UCwLhKh2SgzhH8Q/CyTYYQcrJ7dSm66Us11kd
QCLjd2QJmO1u+kszPLYHt7qSeRGyQv1Dji9h9qRiEDoNztMj17833gwH8wlU
x0qHA3z5x4TpS+whAHW1Lhz/MePWyCm6jVc6m3bwbroaDV30aD6fP2DXLElu
FXcCXu1ryGschh1aHJ79Uis1Qti1uocjBDiWQAZREF2i8LokfpYgusD4gauP
qM+QSCdpOsIMFNCc78EsD/26kbxUyjlvZeGQfw/DnU4hJiEAc++Me/9RoYyU
vT8Bld1ToxGTtmA77FDRjq1X6tDvrPQ+6CzQ33EbC80mrfaxVgQKQ5nsnODH
apnjWOYGY/GNRUMxh4RLUDCfunJm7X4b3INbtOsoA8JCJ50cep8oLj+Ofb6H
3nXDX2Vk0+QTOltun37YMqCsXCaNmnXZNY9MzKStSyAH94D/pqRajvWAliRG
9PXNcaiwNFTNTJ4I7aMNXMu+dEYNE1vqq1FiwK9fyGvCMQBeqmx8coVNlW31
p6XPa+aIIIoD0aSOKPFZw3lOVLAm53lNbJ14gFOoJVCbxGavil8HEppZhclw
OUr3M5Yk2AHRtEnP8Ug8+b3DyzlgUOxk/nyAIK9wO391klYg4qiLDfa7UDG3
UkRojSAYMNsJvjgVMmvWeGuWId3kuTWlGr7RbS0hUZ/5bzf2Ovq37DzkNMMx
aRwJhW0/1B2B0nt9ArW9uGVXYikC69hiR7s0uCF4veTDVoHxHLY6P7rMgNZb
R8/RgtUL8U82UN0LKRATOXJglO/GpCxYfDvdXUKZFfrE/vc9wVBXSezWymUk
9Sa4FOy7rjqmbC95oWKVkjMryNWZpKvPoy2G99SzUoPo3WaQS1VGJdzgUWl5
vJYx1p1iEuhHon2Fv+8PzBgcDHApOk0MoLDGxmI9J5n17msF2SKQ+1PBH2aQ
jyUYcemqMT34YlEykDz7eK8mpF3RxspMh7Su/UiPovIOzl2zKfOIjrEK9CNX
XVL3LgbsAMv+fqlzeMb7zRP+dxlttfJTt6AYFSOfY3M5USnSSb9S9c1gouw+
Vx53qoiCOx4n6NYPZcdbCIT0JU/ghSf3h9a5Ba30arDt4TSMpk62QGSTVoLc
+WQCeKRe+qsioNldfkiNxGndeeZD85r4lYVg63KsamlH75WsFOuLogP1gmGF
yR0hxW7DyYxS7WTUKlTtp9w7UZkzurwLNuxEfe4keEVmCOWz994BKUOIL8Z3
n3P28aD7iBGbx22keHpuIlwg103PR5FWls4GV6K4jm9KrZ8eZGvlHlQqfmEK
nDbOU0WFN640ygGO+pd95w3k4t0tyZDwKFL39wNWbXy0s85oqF+JSYWSKFzP
3bzfPk3E/bTiyUR2ynuPlBjEBijC+SZu5waRgYSEpGSGv2BqzHpnVDKvR3Gk
9dMzVlfAagvnzzKp7WacaBnrswF6s/sQF3NEwX46kwLB4kpSpPbGgqnuNaMS
cSBkM4Lcf4TUQjYT4u/Ah9+XL59MOUuXCW/XPXwqVQPyWn0K+kCDFUE0/Qr7
OP1UnzmrjUJ2IPB5abwOfdW5sCdpt/qo9mU4XMBbGFj1Bd22VCr8iiO+AS2+
GnvxYhEpiURV+gnYM8OyZo+DSpCkh5C4hZcWCQCjshXfOkaKQCUluMpbCekt
bCQp7WK0hUy3lA+MsE++0HkFvuTG8zICszxKXYUpt6ZMvmrCkJw7lreZfGrN
A1kfmginC3COBFMUvnRfO9dSCEkurEFrvarcgqp5TQerrnU0IU+XeUxxh9+L
WTb3bAuy45rQj3SNR1RbFmO3zKD/OhQ/6Y46VRJoiMJbgInnCbyfyLeifiho
YyJ3UdB4NKUkqCuweUM7MTOxgd9vkTWEyeYQQKFtRt3VpktxpPiKs0ZajLzn
vUmLhho3GMntDbWRBg2k9iw+Aag/HsUtakpbvVDraAbuV8zGFS0V+oIpqDaC
KvJ00gjQMbxIgsdlhLnBMEI2akvv4HEn0JK9WpqsxW2WesL9h7PMHUL7AA+h
QbzCsKWV3OGUkyllPgjJ/1XQ7mByAOMny+OTzoCNoOf59qWDQ4ycdAQSD8/a
VtYcmUF79jKKfKRYXzTdfSJauipjbxzgQoBxLMREZISGWU4vpIz+evYSRGn3
KVPeEu+0p4REr0pSb36CerLPUAqljPI8OVelZuD3GcxoUwoZ6FO4rXV+AaY8
zA14lzzlhTiSRZwInJ8/bDaueYIxPSBDrVGGKN+6/er95fhCaz0naCJceTUC
0loNsRCg/dvbNKgQ204vBOr2PqrACX1NYpj74D4mJzuZ0xI20gLa0AHafhGz
D5sIgbekucm4QinHPxkySeJIrbjXxsmTx+irANRfygXTPuiu0sMvOfmx52Qf
jIk2UC0wZZ860x++nOuYuhsTk7/RtU54brO+0ALt9pCR5V+ylzAuWnMiEYaG
D3yk+yTmDwQsKgDVekXn3tjSeVjTyrT+i1vJ7AqgSoFJ/Jsby/8Vip1tBfCe
HA/2ZaBM/ydYCcErIuBPowUjORjhwkwaIzIXrrbJ3W5XLxoIoos64HqT2DG1
5xduPmHapWKlddOjMN/V3VaKYZANozpV450aULuXtKbCMeQd7HSA1G//UyuX
/2Oas5SL0cHrVHzQVFEtXFwNeSSsXtDrWnll0hNCpXgn5NZmDTx3DQD/01WA
U8WlyUvfxFc6w/9oMLlJX6b5+95X06So7eliOiJljQRqX89dWE2FiJCyq2Ez
0LB5B3kUhOY7Mn0FJRU46OcD30bxFazGTOQxIwRrxK2UQk+6GY7S52gAtbQt
diGK0C6XCDgOIYriZ25aTCsFQuXDC50Glad20QQ00+S6BzfaKa5bNVh+KtFZ
jrypaOybypLdZjg+J5DtW9kCyeNcXroFZ6WN5nE6R8Rp6oTLC2KkqiRDefXx
eEW8ujS16N99RRkqBM/ivqN/KzlGCwSlMABPrVtEqgKYNP6oJj/RLt3yG+ll
9e4CrgSkUB1Zw/OiiWAnExE+8BuLBDe9xY87I7DjFg3XmQm81fpAiKyRle/4
MkdewWaWkIxQwgCa7oBMdSNC2pjMZrnwwuQaWfbuoS1QC1xV9iLoRgtIcjJN
R/z6LYKrR/WW6ChKYI5DcnCe0Xxa8J6l/3l6nuUwf8eLsthCcRMOXeesVcMO
CODJyKubjd99Ohbsu4k2q/kXbRZwbLNWID8gvhgM4BmTEU4ZfK8Sy9mY8KGI
IklmyfxFl2OGvrXHsu3xz9gGPTbMQN+M6D837C3x6HqPzk5mgCoLNo+aXz3M
B8P1oZ5aTBp3HqbIexkF/whbBnRPQEYGlQVFjWZyS4DXuUoB0Y/MCtO68Lj7
4oUp2oMKkq0WQOi7kwM3AzXJ+o5Hi+uTL5l9308LVSfEylJWM811MCde4wTy
v+mYpu5okjwqzw/oRBuwwgrZ60ATH8IRB56qnWXvx6Ce6r1f2ZVp/faXI8R9
qx9rVes/NRJOPjx5vZXHDwSx0nmukYubZq+/E7SqSqBBAG+4kJphvIAnGfO0
qxTGFCn5A9Y2bGe0Fw4HlFQNGdWA52GRDAOrgIw/earOxz/5m5fhWO7ewUeq
6mO/fYG2NZuwrwnRlIJBJS/KWW50Y1BOJA/tWCvRAEAfv1/GW5IIRtBRswjZ
2WGYJb9iOFMpoyb97IHFDJ7s3UESGC9tt3Q8MP+neXtfL3QLecueQnRDCuLY
C3kDEoNYtovZ6gsP6yZC+zLKuujpovqRzzMX5K7+GH0EMJlJRQoaCdiCumgT
imIE41m0qmN/um8X5YW1nXR0MLSyDrDhd94HNWVdbOFf2cEsiisnrxOwB10v
f0f/xeT/Oa3UhiniIjuXrh6G4QE8yp1Hh4RC0hpbmMzFfURCm1dfhQ+ZdyWq
djAjkJQcwyeJbqARdvi2cBzykWjVWGFUomzuIuM4a0B7rwXkV5Mhh4a3na4N
nu19P7ybqLCJfsvk8szpyvCZ/6OS0Wxa/bgmSKKoB3llIwCAUSSzwQPZUWYw
GEKUQb+5FFv1nvaRFJCeRgf1BNfNccSDBtZlN5kkGNL6VebxgGe+OzOs4J+H
wdBGXXKWse1Ip6qBLggw5LS2X/ylllmJqABEVqGRH4/Iz0UCK0BzgABZWlaR
fa3wL2amfXmyLxaTuaLaSa4+BeycZP/Fzpip9vxSf1qp7VExcILtMkee3q0B
G7NWHGC3JcXW42ZDmZaNSHXXohzd5gfvuPrJszoLXcafvvyBX5BJ59WM22Dw
UW2jh6xrzh/QKTU42WyqqrdbN/umLoU+wYS+L1/8Z4+UdOWUoLpMvth8wUFF
pY+U26h+ly+HGGqmotojWsnoDOVPEtqjYhPrL3uqsfZoMFz5bqvYaNgJyRKD
x+ejaD08ipo8bSkWKvcuN1z26VUnLzQPFdsIw7WtAUvjLMLjJZEvxtzkXkRT
fky1Cev1ro8jJBM/1PjRqSD/i6IKz9FrXntdsqp6lwH3hKuMNVKSKKR0rAS/
v/2oZt0aKZzcVYpYrnLVfzbZcnzkxjP4s0ZS5IQKMPBMHU3JVU4OkaBKTtwX
mwY71aeVj3uqgTZrdFtKYqfKhPeplDZgDBAPMt2tEL5SDX0+SRPqlIHKM64r
2trC5b/Py7b+XMLbWq+VaPP9QXICHSzWYvRb1VjSSaEt0R+47o6Mu/AhGSbq
rhzYw2ial/FQowk8tFXDR8yJ8DEdAw+wd7zWhSfcq0SPO7fqRurVlg6Bwnga
pBbHw8ebonEBvX4m0xaX11SU5xtZZ/2mPILT6CTTu6oK6HL7HaNoJk5cu9hd
4E1hSKHgJJj2pBhwrcmlXo9ugvDnVrk9g6vMVtfSpxJ9fKxJMt7TOYTuH4Iy
b+KEkpjYHusvTj4axTpxvz10Sm3oWyg0JJ7KQIrU7gmgb5dJoaTkWMUvihqd
8yNa0q0mTsqqY9BGXdS6Wd8Bs0ie9ztxUWs90awG4P1ecJ8hhHSo3oWeTNJs
UmA8oK3kVROLg6jxq/397ra1HSC1IYNQfJQsVHw/pJcDOEtgCJA6B1SY4iJb
3RAztkx2dZt6j178ICgPmmLtbt7nyl4RUdQHR7fK1vMq7TZMe11Here4rkWp
BW6kqNRSWyz0y5+E5AsXgjJYviRrEu9+l0qYp63s5qMt3xY0GBvsN1pbwpx0
jqONXXg7LjjsfAguW60JxI0GDENtAJavHVZ+plPEWo7iX02yfT8qQT+vbElU
peDFCLY4NdehHyMB0A6LQhNQc50d7eWrV62VAvslIQfq1R9ihU2BZ4SgCTNj
4ZaHoNSVvQ0SA6dP3d/MDNqz87q7/4Q2WO0yNX40q0ORf0FMCSVNfKavJcO1
0L5PwyNeE9eMOicMFxOw2Qlb7kx5VcC/p8+6CdR3C00D/aMuby3Rh3FmCJ27
855e/YmG3WXSL5n8jSSMLumdEiHsR3IKEXf8tdm8CQiTYBk6gzh63KaDsOBG
NX+T3kxg59CIJ0NXytU8Hgo212WcRtI3mLDT36axw8W7H0PR+nxAnk7NmB/Y
5YYLJszNKuA678YwOdQzfV1g8Vq5vZXNLqH54VF+2Jyx1BeQEa5Dc2/lU+vR
LiwJER83BjxpVONSCU32lRaMXR/JSq9z7KxdQPcO/yWtAfd9QO+WSOqfNjAU
L1yI6BUPt24lq2a+4lbnyL+HIQpSm2/ReGcE3+7gJX2IQHzCkM52Tfw+CyZU
g1DFWl1kF/Xy32u/NfxFTtxucGyVODeKrEZwEo1mRu6qdrWDWY8j3xGXE5Cb
WUEcL147McrXfgJbE4DMiTSt/0XH+ow61Z5gYO+Y8eEj3SMxbbCA5tFxjy21
L17MYQy+ICXCAKXeznLk/zDS0KyMCLO8WowyXnjpLTrrN68DK5Ti6nREje/w
0HVLAmkT/DroqireO54GqRLWhyzfjEQ2Jx2+vXXk1V+Q6F7sn9oFoJprtWaA
9P7DjE4ldq7fOrx4j8+PXNbBGyot9oBh8/bRI7K3VIcyH1Ep80MwDbc14vIp
DcIK5xqRoJGmNX0RWxSt/yGhSLGTmbocsmJf75lnxnwwuBbo53ljntzOzXKK
NTptG8oepcKrCc8/W9pID+7DYkYQbpBY3PLpP+5LkWkT1JyM6qdqRmvJ/UJq
Ujo4V3sC/8EjyLlzBFDiB6eMErx0Q6COVofk+9dvSOPDWxO0nxUn92SeHnBP
ni1Fone4q4I0Wxywv/b2O/oASCMiOXCi/swBnSSJeJrFRNk1gV9GWK/FoOzp
WqkQ0DF8XFIBLUEqeGfmWDSHV3TeaPDFrS64rhtTCK8iES3GYcCJlY8msceV
p71hTrZtGv/sXtQudvT2ymQ+/kNIe05pxQCQFUktOnTn/ntrGUquAaqO6uds
EJ2h1PrViQx5k8OF0BFKzbOSdbhQXBbkWEhJ/6DDjgi5tj0N3+fTr9i+l0z+
4SlyCUnoLZ3z7+Fxrl+UfGl3rmTpoBOQzT7vYzCXPIg9gWlmx0KIGgvgmrZp
08GdMWBgKk5NyAvhWbcQrvgciknuD0+rKjzgf+Jl5iMd+96+rnZFmzIz8pPf
blDNeZjix2rH1eqaEYc0WlOoacb6tTtJTnPBu3xdimoqTK0QxY5UG4hRxti4
/JeaoQ5+1Zlay+5sKCu/9cFxUpmlKlybdWSDFWsoTwNMOXKhB9pdcge2YZPD
ifH+q6q2Fx1ceXf+iBH/sEiAQM56/PCkFaBOEU5CraDDjhCETkdplsfn6ju7
u5XHJYrijWxnz04loe0KLN0Cvlng3jIoLJKbq/jF1eP1qEjKHLYo0ufxg/R3
rSe1QYfunm7ofTAamJeL4PNxAqeXAGbIDfP3OHPiZ+6DI9NIlnqnHzEhYcsn
GFIniiDeNiKU1gZ9dJ6w50uXhoYKVIttiki2zyrcGWQua9JHFesW/bfLZstc
8sh7mEc3824X+R4yh9eSyVq5R3+dSnEoU48uw+tOghHQGABbiOMjAYvtN0we
ENeMDKfCBAzTY9rsHBMClMyHmVkXlRvu8mGlQcLwfXRF0G9LF5mnU03tCt9B
ovecg8t4P72KtcXvdwNQxE5NoCotWwoyjHtVtdmpexTTDjWbdRmnrx4ZWvC1
9PZ6f2z0+8oidl14e9FTCVbdQUWA+w4yF+H4iBsEZrrHuYjNAy6TAIw4cy5k
V9PSUONAnmCFY59vurAClsRTNzVZPeYGAuCIkg2RLBokeEXJQ7DBcbpWuDfY
hyvZbGRgmsoCJJrsTcbdKlwpVHLRU4tZ2eEmT8nOIqiUUoVDfGVcmY4wT6DC
xb2SVm6IswWXj35X8eyEkYYVt8/DBwxgZUcruPqRybuejQZpb4nU9bfr4T/f
bRMwxNITPwzO2mdV48UxDmTe0ZdQgFkueTndxD0lKWO81f6dD9q3gfUnHgB0
UU9/RFr1qG0gam8ct9Mtd4iQpsHtqKmMgomFttnqAsmGsn3XjEXCssMPWdH6
YlT57qoFYbYc+g0gTS45HVlYtSWmiOSd93tCg4CMi2Q8Kl5s6fWRlBhtgHDM
Ol1LvHhnM6OPg24GwwRg5TNJ685O945AA8CVcBPl3Ew3AOuVYFEabzN9Zb+S
5p7bGTWHAfEaO/tcKpcF0MTOwDMdM+GYe4r1WJ2QRgANiIULcDaea9ZXhDwx
qG6HjmEYRdqk0Ss+LqxTN+oRFPZiap1yn2gRB2Ng9/3YdpbW2ZDPREfvJMJv
Us8hvi3R/EpWSgBvClUvRBwHFs/J2/D+XmPO20r+DOD81GvjOJQwryy7EZsY
r3ybufYGYDRHLG29yFzgb6MCNG0yUfim7Ia1SZPVz1FFwJ5vJgTBnyIzak4q
A1et6oix3qXNYb2Y4mr1IwyDRWocmotJ9jhSZN9vyMlATMFauiegyh2xs27L
LGEbRK7oC69N4YXoMYiehoYSWOzmRJZgaXxdYq8HEh7P9le9nrfn0ViHtKAM
ly7SrCeHuMZajhP2YTRsYRB1cZX0/9Vw3iYold/4LRXSS3R2pYV0lDLa5/Vn
wUc+ya9hh7gK1ZWSrtXyq3+KQP8EQ6NLghAAofKZBtZlsANPxvwLkqvycXMY
Y0HlV3JPQPlYuk6j4JntuUz7FW3Fz+AHN30jNICk7O8kgH8k8lMDSIjNWD7q
/go6KpbDzfArO5cQxLBOE8y1UZyMyRVaPEB6xKr/gH3mcLKCwd+ZwdK6GCu1
9AvivGxZdyLNrglr79V07bD/2GlBrkMSlqXQEyR9jwJ3dsfovY0O+3wJ5mGE
VAccMUBdCyWoT3UV5UVyRx7Kq5k2Ckct+hD8xgzivxXdtz8GJenO1HelkI/p
gr3hHYNt+ARF8Eq3MkJNooO4jKbPGpUAviCqmv/13bcXZ+daQUA2TG1myORb
/czSMZWOSfCrDe2493oMS7Qa7MWwocV6KISJE4rYVPLpOZ/XUSlAL07RUab6
kRiWbMcTWAMIB1NhuaNF+bJNlq3eEAPpPJj8NwSR3fgwmgYmE13J9xjLFG3q
EGxZSs8129GglYK6gPEedEJNga8Q5r1oKEJHBezNOBGH2M+gYWwAsJu9zrkU
+DhcuAwXGI7JQZadr8AWAJsTI62+VwPE1CXm3DxjlO4Vqxapk775dgs1j6X1
eMALZE/q9Ce4KdiifGSWDsfJbGJxlF6uEMzdwOWKXKEJeze94aT92WG5teU9
OCDuyS9jTUt3OckRcZOI8Pk5eTcSt0xBAXcRsQ0WPooma5W12rBGX4uN0Egs
SitGLjtAkVIBqmsNAofxVfofn95OJSRs8ermofpJfm7Jblve2T92fJlQCzPV
xXdIM9iUDH03JlWF29M+0RmX6s6SdLsil6ti/W1PIh2S4YfVZDnbpIrOG2xY
jzUwqv35YtCGl+5ywN/kcpnR4/J/V1D+diTwQm0AjtiFXSAWLO+HFHoG1rkj
zS2iACWPG0nqifFCkGuaTtFRE+nJuyGj7OCn6qMMroFz5YeL0fqwNKJg7jsI
5OUSfHXWoZedJacOF8fWvKq4bnPDwXrWsq9s8uQHcgAkr3UKmpN43r53Ffsf
Xp5XBLe9idNlXFiHNXovhjrpvqO/pMa0PzsvnGt658yCZguzdhONxkEkQrMG
3LxG70BTcRn8qvLonMvuwM5JGvdVqe7cz6GBkFVBFNDiAkw7xvZXQnvetnOs
O2ICkgoC58fRj8Wydrh+vZszHxgYoGZM3w0tKdF7ftASPWx6sxsuXvOsEuHc
7HhcDUyLeZdb3xNcvqMPyE+GdcLvxQROPhweZKKfzmNbA3moYpWf65TqX2y1
z6rHPNWLf4wC7Onkqmk1OUBKHgIdGu3Cs1ch9go8Xf9u1jdrQHCCJiCOCWvw
C7mDnDfFuQ7B3QTEfWhqQOJh2UIrqlcapSWBSKXk5V/foef+nofZ+BdGiZ6F
OtrVumCDdZd8Bpg/X9uoZbdt2gO84sQobrFclgfltAFdb/R/dbUEipGRoqmv
RzglOgqvD0nLFaFuQDFUD48g90a5eswZkXIUyD54HpKaBvf1w0LChpNqi7VI
3pa1jQ0aG3P/DDBw8hUOlLiE/JrWwCk7bJkW/lG/JAVg3i4Qh/9+Rq0aGZ7w
jkpeQ1rF/kieJ+CYsax9u+NfXd70isJj2/w/lYCYZwnPMyqHSoaMfnLFmjeb
yoId4nJ445EvTp8SxqxpUPuE5Y2C503HUvwUIrhXJ8+Vo0WwJShknVqqgBvf
+cFeprd4iP+9waGDe2XDLp4vxAlGVGFwo1yRO/cECfOxaOAdsjrsgIsY+c2h
UE1szvpXFS9JiRjXWGLAnbkCTcwFKMLgVk6p4mePVYEk4cIs3I1GsV37YF8l
dZ7sQINjU//lyz+pOcUDcxqGUV1ZCkU/0hcJvgk+bCvCz4AHa9xm4qMryHPU
zvuTj7NfexmK0BfiDazBcVzQ9OuaeX7WICqsFzbYz33PuLEiptg6m8H8vhEY
uAxNaLBzLAL9Pu5j092+4zxe6mvrFq78CPS1EbXauzY548kDoMgXMQpcgtvO
1+8OJkfvV3kim2yPYqwYTiTN89JTp0DznclO8Pk+fe3YioFc8om68kDJ/gts
h1kCf5P3unI2uoyp9x7khAviPEDxjVFOarkgr8c4ed4xSgYotvrsBWNWaX9Q
QfPbrIMqbtcNsXCZi4eKg2MfxCV+He5T43NMcwmcbrTaPwk+DVhWnB/+vXfD
AjE1bn94VUDjVtMPdY3oOG8pemjNEGKSlt0eHTYa/EV7GGy/P2Jd9Jt3hIF6
QKhttpOmXLkROoiXv2nHQLMoD8/7MLWijNWaspZ7HqmFK5SedhlFocA3olpM
eim3leFWvCGPflDmr/gO7PeHz5xWNpLIDC+MRoxSSlGHgr+YOS/NKz/0xlCH
2r6rBAbJlsJH4Mt0w8KU4s9pML8aW97ptC5Xdkb3DxsiqCMIVfuZZj11GkJo
KbG80QUn/eNVZxhR5HfcZNzgV7wKFfW6iXVUIrCvJxKBGaKWPFoKyEkuq45l
83S25rXo4+A6Kp0OhRk/PTQ9225DCoYmOV8Kek3v5RoUgdpS5BU9j1THXH98
xK+7VEAuU32P75D5idMThZsaYQzPbdkkRpdt+qGFSoLpbUkrmbaZCpgx8WML
NxB/HoCQarR6ynhNqLcRzNVqZm2/LVhyRWagKkpWH2+jNSvSFRwIA/3U+S9k
QdwkcPaPizJKFjzIwrJfB9J0rR28OOZeM4RApFY86ApVz9KRYqDOO5+11Fr4
VSTsgfk6JUAxZNq3UmzK0FinDnNi/6/RVU7Pn6LVnG6akC5/zrfCCBVBBlhZ
rNEyYpE+OPK59zE2xatDThNRfAsaHpQCIsXyFt8ZKy/Mx7xhIA7VqY6uK35T
b0k6UktBIyCX6xmEVnyNfcjIC5jDkBtJkB8tWV0MqvCu11NT3uUX1IH4uQPx
Qhj9+gljMJed5v2vU4l4LaTR2+6PY2QVprZ6DE+16Ge6ys8VY2pCOCnMNBst
yS+/YF+vQBZgrwEARJ7sKnDorZuvf16oERscyarSA14KUjAXijYDyQVx+Ae9
+V/uvx3mPgJvHtO3bfNbS4YxO9TzBRJUmuYqnY92ObwTnagl96PycgmspMik
wjzYqE3/XFQ8AwhuPoJ/1LXCmd9SNYyezcNoNX9DsOqDzRZiiUjnmSi1NRb7
i+GWmP1kr8Llwz3mSNNCQ6GckuShLBan4fIz6xXEnCCqZrSBSr6Gc7dxL84K
ggUz0QnpPRfVirZIyHJuhsb2byRb+dJ8xXliqBh6zhO6VRvfQO2OOpwGgm0/
cvHWf8W+0+cabw5khvt3MKVqHSp56nweM5j7AAiw5vHL+s/d+YLWFa6FP9O9
IRHpQDgrKsOYMLEs6TWLMR1n+4q8RuIhfB4Gi/yxtFcauNRPz3pk2EtDEBPI
aGbS6WAkYGF/opxUT7kiRVZlYzGDbMc0V6N7kqFBOthKk8QT9htA/9mfusMr
CxZ12A4kmAbgbjRreWXmX0WMhB9wFMM5tm51qe1EkOOP8TAzXW9riFzWYAV2
QOvL9tXYQ4zPGRZuD81MgAMm1c4NJLXbf7eOrMsE0e7hsnTR3WidVSm8z0nX
uY6EVRrZGSxn0trkf3PjOwpgkJQZJC6RO7rmmABWOjRcs3XxI5JBLPQFd81R
FPwG4IpW8GlunWhXXs4F/iwCnh1m/4pTSoYGg88PIV383aH8LXVnYPF/G8/M
rCC+BaKArtHNnhv7vYrFbyaavfHnksgi3SXwtfyQEljVxF2WtlDRh9Jxd1SP
XeN3b2AWv/r5/S9sbdGcUr+ah6IAwUsAGp/VOZ2JY8B/aYSNCP+l3+csPEu2
7eso37ne7tHLNdVopA19x3jKgGkZfdFSHuqutgiaH8r5S+vVr+g3qJ8TmMk9
qyra9eq0jVoIlZdVAkHxgDcwlPGCUhOIV3nyQ977TAANfw7WOE/pseaT4Cn6
wLasPUXbQRT6uv+VG6gtJ1PdNUsVbuQ3mRr26Ioq6EKW1E2bbgWWLwkqlRr7
Dt5jtTTyLAORe433Q4yp/uV3FPNCMRg2REN1EXh5wCRjf4JGHLpBFT1krScs
uW/Qc2ah0+ZYj3zs5+U/lck4aOtTSD3C5AY33veapEZrFbRBMs2J0YMukdZq
w0/9zhz0MlBwXPLXaWds2+Lg+3qn/cVNpOUgZSnC09AdC31rumJGa3Lz2MT9
UK9TN3KWoagMkZEuzDoryw+zwc6uBCIQzT7i9+01kNO1GRErYZ6zOhoZ1dB0
f9XhCZeQeA1OUK05AqSxcEyRlQi0O/+cZz63sdxKq1pyxa0zLeHQtCmxdSlb
PvrDaEb9mIYFeTurtpNz+JXQXLMhL838fQrEoe6yIMWB+NpCpspNRizr3VcP
tFoXudZxYMy/E1FgRzBUxy831EgvUrqRcYfNzYVyqM1ImkQLClIC2RAs/JaJ
gM2+6cMcVadeDqpYKf8P8C5JNJFZmre20K6FRkNQNtLveaNjHDLEh2oylHio
YmbB+VbgeJs+BFyt6/YOlU6pGl4rzVE0g70vsmPX5PlkBQIPfOajIlIHMo3H
giCEKObVBdg8QWX/fbhFKaj7PX2IENIQO9PqUunL2qsPo/CEaG/NjkyFX0sd
uutwvnJeM2ZI6q6xtoTag//mPQD3wdcI5OYbSLtE5i7RZfQYir6kiaarMPoQ
sz0YFI79EYEt0W0loss3m/f0TyFmpaBLWsdE3pCaf7ijB0Q3km3klTds+fgG
ytDOQVZm1jADWtVvF3dY3j1B/QiqBn9kShGQfiXZl4uMUx/NatwDevlP/z00
XzhROznRGYhGAAAULgE8O9Zf6aDjuEeFEjN+PE1qxTxlmqA9NP7bBRmqhvD4
Ce+CkaQuKOjXrJQz97Ealf2VseUNWPI6z/AWoerqAw/fH/4T9U18dGGhB812
BvPmNiSDq+8b6xGoa2PaC3TYZb+6d0Bt1piWLjUdPL34j9MNTnPJuIVlQz4K
+Y3VHVeDPfuh1Y4T1kt81QcgAIo2/67F1U8/6lSf8u7J5C6oz2SAYKYIm5Iu
OYjarwYGyKD85JVUiT9DkFdgqK+yOyJZ8uGX72KNLiV7QdZZyUmBV59Dtk0r
pYtovd+MXbw6HGx2+oYdxpMkMvuhNZfQ56tzKtN/0QLdFcC393w8AjVV7nS6
ZfVdqUiGBnF0yL2SERA5oATHa9btEaKtDJ6I2BixcQriPZdF9ChqmpVaulSa
vEei9GbA3PaVR93ifvl5hT6v83zldi3X4pQVzqYCG/isVItwRTepFRWq1x4L
LCL7WU00ZBLfOvuJJZKiF63pf236Ur46bMfl8dApbGCeUGY9htAZivUO6csy
gnjxWZFEX3CDviiq3ceEy9DsE99NSeMoC6j4uG8s3h0kf2SsgaiIZgjP/14k
Mp00wm931XtNw/sOkKp2h1r37DNAQjRB7iJxGgPfwaxzZ3nbRPFKQM4NuzXS
X0UIGRjQie7ZAo++llNLo7JKXS0YPCGRdppkI9T7nOfMZKVOpHVny4cphL/n
u2s3samHZ1Mxmwq6xIKjm9ooFvXb4S/5ZoqLUEVPejgt3I81DyY78UIAvqG0
4CW+bxBAsmp6eiOCgCzlUc0mAbc14DQK7C98zDfE1U06bCH824BXQfCl8KYk
Rtl0QlFGTBkgDsq1/hZMcmfDaYmd6umwD/tJW8b6DLc5QdwXqm9CLEPGCr0t
glMxgf+i/wh0agtGjXmCbrkkDasmX52zUHwBGceVZBB+m54UBCZHyHJPBEWr
+1AAtuzR1z8rxMpW9DKIfucDUSjQItu9skLWFxyxJTO5fGj6gFQm2sVQZ3XO
sjxRoBWSWlian67mEtVoLcS4DAJY9YuNZC4pHe6jrXa2MB2TMMA5C0qrfWj6
GBVa16G4K9NFwrx41bsr1e9q9SvIKtMRKozBxUScmRZAJx1TEokvoZ1W9oLo
k8o+4W5F5AARY2qmGTmOeyuNhDehbCL2beR6h2UlR5gvxkWzpI/pfX5kQinM
Ix0R0Opncinwbo135fzLT3V7oO3qPwZvn8shBVwwXRTtBehhQaiSo/+KESus
BIslM4jdE2PgmmBOn9wmgPpoujCLK1HZmIZutMpWSB2lbeOpnkGLDNS7X+St
ek8mrhBKq1EgeVvzJeXbWQCNoVGVdrGetbe/Ut210j0r6niUvHJp1Xg+8X7g
aSH288MaiDkLwvm3ZKnL2UsAJS2oO+8zd6+E18ujPTj6IbKivyXL7yruiEpX
ylizRQaXnYKARrckkElTcDjtU5Jo4ZFIzMXw6kQFYnzPR/tcIXpHXFgwfYBJ
6MWjJguyBQCbGi2nJY+QZAQYUKIfMS59LAlO7LkWn2HQSZi7vOvSaxAZYF4L
mKHcMqNLp8wxY3QZ61eVoNEXokPVQS+Kmhe/BmOKIfECMnVJ7CaBDHqdBckq
NWZvnq2sjwwtKt+3/sLnq6NAH3CU6dlIVtQCPj2UY4pnN7fLMeTn4rCOzBNH
yzlyQN5FF+bNONj71jcC/2SXwABAOoW5KgVUlNRA2xyRtReNKe6wej0MsPxA
29tvwVZN+hpyfjZey/tN3wP5DPZjWMf4Ptt1uRoO7HQbEmcrUZ6SIl3qBx6I
BmT7XW+s7PS83zD1wZnsiZeXCCbJVMeEG5DmgSCBQ8LU9JxniRNroXC2/V83
D98kMr+JpihFOpoWiEtjtOoZoR2RJtN2tQaKyN15ErTB4jr62JEaR31ifqwj
iqfWhSJ4PyuYrgJP/wW98hL+LzNKGsDDVKl7FypSPT8H4oJbwUWjkjIXhqXc
2r24A3nY1L40ATGvTNfRuivnB+RishX+WPheqUS12V8pPYJtcgA7iWiJqspD
fZlMnk6gFJH4eCTmhEri7SAvoeE6bb0JXzdQXqOXunITCJxWalhvQ1RiJK9T
LLcdtBxNw8/12UDIlcMZMlDP9zAgJHZv/8XD5nmA/JQrt/OpKql37fEXf3Fd
gPCz9GbScBSfYHS/kjWZ2RNqSka9gNPzlTli7mGP2Lsgo/OqGLqgfAvU4Y+F
INGQRimQR3Ech+kAEES6Pe6zN2+fhHy6739oik4J4zQ2Lmxk7z/vQ5spGOmd
dnlKPVwaNn1xMh/TsY5arQsb0JC+j+GkCej4+/2yLzyaVb4J2GqTVqUHZrs3
l1SgVUOTjpYHvgSV+JdzAUOywUJBDE4u7PCME3UFyQFPIQnxIAmlJ9T9dT9p
M3gBzNURCLVeKiLh4+lYVMDW9XK+YMwFHMdKlIBDBYMmNnhjY/QolECiLXKI
w4me2AUrnfIxH6sy5L3p1oQLBZ8hKhoFGRtK4/3E0FE1wSErgSNb0gpffgco
+HkdNSlH2bxyMPsdSBg4QXI363moiIAdnwQixYZd8OzU8sKamTEYWKrjA0fl
YHGeXwS2L1NDYlZPvpqnabYheTYW1/tFqHPDfefDTsQANOZToP8VInvpGKu3
OLoQmlHI1daP+MV/Gug3IuCZr9OD1sMI9kCtAuJqnI04t4MhnJo4CoRAxHSH
ttevEQlTRpVnJuU9RUbI3Y3yhOO4Yy1YjE3oE0YfsJYOE/5xGaZ0/ocbAz9w
clfTkf7eKhWgZO1ld82gAPTY1J2qeLUx/VN4I/qvhhroWG2pSIxNSLSm14fq
wu4yBQefoC4XZY1Mp25KRLJ+RX3AvnQw+B9x6Po7q+VV8lL9IMrS/QN4Iair
oFOcXnsoN80ALWk/n/DzF9pK40cpgrFRgW/EfhHPzj1ieMkqQRyeMdZvm5DJ
DLE/L4oiUm6UUCB9yXi5HOk12ETVp1yLOCr/wLfox4/REJ7pZUVUpQni/RwF
+NorgzAVTf0q8PM57F6WAkAcCCcCGhzgUnNy2tMOwXEHBK5+QHRN3Av2amXP
Dt3NqWgZF5qlKp0K5j9YBT5l1lTC1779K8INDk51tAU5wCkn2AiwKg+bP8Po
LM4mCSIhGlMmTE5BNvocaTtNrIj3P1Lkx/L9O/4tTmzaC88BKeXZlNBZ5gq0
P5k1AibD07z8V2PPLAymflCrjCy1EIhlmWQUggTxCI4uZGFGj27RzHlF4T6J
2CtLI6zfQ4F4OJO4YQNYQnu6vIxZDJ+I4/DOIVPDLQg/JgpPQygcrygco3vF
2QSzRrVkv+ukJyNPdvIOAVS4H3lMcKa1X2FBJIbOxdchzCoL88RaVXYgB/91
FXIbhzkwN0grZl7pq+9sMfJY7GdVII2rQSBKqwubEHwQlcP6JZwC7EZVzwIu
+ZYhxY8OWNO/++1Ype/ZojpgYpwSqFXVpH32FBLbNtG1l/w0noFW3LZmy80z
vCsumNp2eeZP/G7A5gN/IT7fpsyiz+3JhgVfaYo2PIzqeLnRmnGdelp+KbV3
QuyAFCrqnkb+Mr7wqA3vZlSzsbY3ZUILB6fwDJTTHUFoQEBhN69JfLG9xHLE
bSo1QawXeSlhdPMy78LOrFCSXLq4X77OS5SyXLT9zSLORe5i35l4KeKrUPRd
8q208gNMCMHyNOzzmjQL45XTuGLKI9/6QSt+pbueSwferbsuwjimgoKPImVw
tBJq7lUAwbmZnJRxHji3zNlMyM8TdjTjBfXGTd5YVkpDJspv2VJnx/yc+aOg
gdpOiepgshlAPcEoo5DYL6h01I2ehzGLFEwNnTq0qZBmHSq7kiZULEUPT1QV
MVUgA6oVabSHdyrtroC1R8lunQlGbtMRQwdOgjmv5d0xPpP6qsKk+RTVod+6
lp643zLPeBPEUNIRCrZsyPh0WisyJWrvPvd8uAE5RH6J2lIxUBJECfND8mxb
Cj9r+uSEAkEDBAK0HDabn+YnDa8ybwWYq0wPM3ifhmIPKotmqdiX4+12dTd4
SbdXQwk1PGpiTufxJBl2Z/Ol6Wind3SSJhut+gXtLGhV4q8cxuhcKgEebBW5
iapX5k6JIuHmDpOsgUQIhF3j6ZXn/VaPJTb3Vc8vg5WgMN4nHlLZIN9reN29
UssxLKYEbWhTD5GGXSSL6cn0CI3rJy3GHWbHxXmGiznMzZGo4y/CEi0F1k9R
J3RFbjGy26e1rXCRdKiSViAzgyYNI7Nv2LBAYcnTkas6Fv6uySrEVHj460nc
AEPqQW6ry6pRulVAwTHkrkP7j37/MwOFadrzS/CAOhHmbRtn/ZTJc+ej8Chz
+u1rlGb0h48N7UpB0EI9/eOyldBfAEL/Bvhx1ETxBQ/NVAxfiLZ+ygl9TFHI
e5g23YggyiGX/wzK3FvirpOg5sWAmvVuElQOa3bZFgB6rrxBXSr7friN5Yh0
QEre4Bf5SNHGAVgEbAmf0UohqZdMeCx7Iri2oyMONDRQFCqQR1elijQA8oTM
iWXQRkONQ9wiinM8/dbFEJVGPc5Re1qtiYprdywmYNDv6bBM+EdJa1xf3MK0
78QnMdOSuidFefjekEXKXPzsOEgmf0MRKO5pYjGGOYx2ndYsATGBxG5bwcPe
Crk3SDDcnMgIztepr6ct8a/1b03k/BGYuALmmLeUmb+CMqOJC4Z8vnXq7tdX
9bW7Kix7DkqK7V6E2xgqvxNk0mbtv7g/QfGg9mDslxnvORSuxeFPu2dGby8L
3duxsRUrDWFNm7FRHANJQ/wLlbBEk469kuLKa7sAzreGXMpbs2UaoryAEaoI
e94FGcqWrlrMuwS7cT3VnyPceh1EjphVJxCg2Ujm2piUvAnIdXcy1TWzEOA2
0org50FhgSazdc+Doxr6Qn/3Xg3pf6aUj+YtaODgS9SG7wcaP/q45v7MiXYG
/p2nfpvMqqFFLWV4hy8rUD3P0n01YjJXrnBuBJnvGCeHkDCDSIOf2cwed/Jc
urPcTfd3dkuqa6tslKSFjXfP/qhlzvcHNLh6I9/Tvv+oPtE9LA3PpnWF5Vbl
5s6H4v6gz993FgBwBz0q/vjSJdJf4frNP0Q1JPG1+m9YDWOlYTGmfRTfAmyw
9oG+Z0yD1J48TLi7zecq1j5OTBmijNYrflpUUbYucyDpPAAijDka4X/uX/yr
13P0SaDGaJrET62nxUnPYNElwmvSOHxD0IZS2hXU5xnHGRMKkUmTnqAe2R6M
rT6gseND4hfOP5/BqKFJgpra5OWXXAOKNKAhAOcL3k/CFV8ENAkHHV0u/EEQ
WxbkHad8JsdHv5myes0vrgGdoZmJl3Wf0Z6Xx+MsQtucsaNNjJtTSGYe/vwt
p+gZ7MUg+kffztOb00RbmEtCk1vh2cfCOcg0ZenaFMKH4rx+L4vl1OlNwlfo
T05T7o0nbbPgERP0max37HqMDdx9HSRwcjHAJw+UVlUvmj7NNmsxO/KDtQcr
D72vPP+hP7k/ox42G+4KxGKzYqkYLpN/e8X+Qw6k0Ox86i01Q3pb/CIp4oF1
5vSMN4oRc6m5xK25vmXI1H/atFAVOotucX9FYXO9G8+Hy7TH4ZGnXpOCidSL
MSZH0utramcNuOjokc3zvbKjiCHcBuIBwdCBzQBrDe8q+RlsvzKbnzOkxPSX
rDJBlRAdgkPycqPOJwjHKTD7vSdftqy4ZdGWtdQ/zzlsLgwkkPqwMb9L+aL7
jNxV0ataKxif6WrsH8sI7cHmtUOp9ORkjPKeno0zHqcTAe+keOH8QheLproR
ZscLZffJd/jH9yaTPySgAVK8gtFBLdDMI3ZhIyHGEw/Z4jsGysjtSiMN3Aw/
GON6F9mWxzC0LUv1v873y+fy9LzpgumKXjHLQCFTyqU2pKjTY1jD7Il4c/eE
cQiNRZWMRM+zmYU/fNImdAslUufd/c1Ibr0veXUjPg6Sg+MQ4O5Oo1fq0Oq8
VEO6xHLmc3Hkgu/v8AtqjO3lKBfPtTluHD2xmwxAP14Iz1IQlVvDsTGpqLBX
oII9ifz3iPhKxTFv5nWa73uPQSMK5evB1XJ1kAdQ0v+pKMzg2QD1BQES6BcD
UEQmaC69SBTyOW1TB5sqwPBst3dRDGUCbD+nLwgEoGz1ZGYxth+TKB4pTWiY
h/7T7t66Y+hUGo762aMH8bH7iMxI3z/XesAgH1vX2PlGBa2btzIPqAuywwAc
AYSIM1LjgH/t3IlVfxK14oEgu+q5GZqikXS0Yk6ikhHesHhqzoQMWA5BOVIj
NFGkxsIRHcZj8Yk/FqvXdZjJ9yPAek8JGUtJN1y3RpFhF+ypHxHHyNZ2uYSs
QIf/nFsqmGhtZvPpx4PqNgNh+eMoTEanWSdsZfU/OImxMj3stwwBAyy3aB4G
t/vryxNt3X4jJWbnCWYKd7KJG+fVB25Ij0zUvPBeVHRKLaxhFp7ktbwb706V
1doSuo1ybIuTNalvRNUtHxBFqacd590zwhrhkH8wzAjzsW7EkkRYqFrJaLw5
HbMIK6Qv7X8AOQGeNSpyI4L2foYmA7Giqaj04FpkP8g5pScw1HNu9gIBLk9Q
XuMuCZAv0mgf5gkByTLXgQ+LDDRS0tdTuRGrKDH9Cx3habuxWoHPucQT57VB
dg8XT3ZTvOwAaaL0t6oeu0eS7huitBPL/Marh55ZHBtTjLl/FzOB7vbbMTT/
9TO5q4IimY3zc4+Ooo9pxiykDS+Bs+HMBi62FdvzcxrnC3lGScHoWHCGF3hN
4Ae4/s/Z6HdygfKr0Vye41f0c0oqTDWyTyp7pYqiLPX3TUeQJnatQg80l4oo
xhRD3DrllzKLwpYwXyDxrHhDvbV0mH7Utny5SGgoihNDkOyYXTbftSaFizoo
sw2xKDCg2r+G33RAdJwAJjN0Z+Bqu6YIUKH0Y9eJ+KI0Gi7CeWj4B5cxSmR1
em1YOvlAgV9ZE9IJqi4BUlCfiXwprGrl5S3t7DxGCu7WHs2rtNgWPREDG82B
qxuMHzsWLCC7nk842Cc0eco8/olSNGrdmN5Uq2SRNwIine/T9N+/8JsCV9KD
lGbcDMvvgg8Zf54kop2YxAP8QULnVP5USzocFxvjZQtSiiSjhQXuZF1jxJ+A
d5aFrtP8YqmN5i3eOe7T6F4gAxcidMsznE35pTdrD2kx4cgSiz+U0vBo7y/O
uyFtPfaBQdqyzx2KrmXVu7YSOKKkMUKMaQsg60I2N8Jr8HOjMek1qS6baOS7
/kiPXh9yy2R0zRyUGOi4h4MSN5cAvHBnXWjbl1BTIqwPuS4UHudbyf2fJPOk
TQkT+k7x/SG1AC85taSQpr3PGb/dUzxX5hM7AiV7le/b381k1UoBWLWwORgM
qkTb4Z7jpXU99skyJF/tagS0MX4HeQLySTO712QbEubz0Kni82y6Mt5U3N/I
CW3dTVcDOKWQM1Is7ShJO7y3I6A2NnIkyTQme9AcftbNYrwR24t4EN5WdFY9
l/qMJgNkWZj2CkROjS2u7KO6su49iyKOT6tO8zruQqFUUjHrnto4iVWJBiVX
hqCPajl6Ux6Htu52XGVZKazv6R+XBcwaVqMxMrbsa3M/N2AumNz8KNMF/o1L
4+l4456WQwPOHwm4XnmwZHR+rq2YWHmEVXGMNF1Chcaj8aMcFZ7OOWaJbfuF
wGuK5bDb+FD3Vqss7CLj3ma71Cyv3kHnLHPu2RAS0tqvRfER2k3kcDKIII06
Cb2sCyMgOYeC0Vu+rioLw7FJ4pJkypPUtW7rwwalTQ4iyoazUHQFeCxKRKro
2JCzYUk/DOtiL3CFX3mCaAZNLxh+YgskVibw6POQr2Sq2lyEig0qBiZjeAWF
XNvIV2QsN4Iz84AZFzs1rdmKDBsG6l/rTn1hDtXHyIXE4AmtKxR4U3g3MOc6
S5sbjwff4ydyPBxJhGzT8b90H+tWgZ5VDvrfZgw/HyrvJv4Otyr2duiPVWAK
L5A/Ie29qjUp/zwsPjuZYdpBKtL4tnGtNW+KM4Ns4sUfKoBQrxTaCPaWoaXV
PDZy8J8XFi75FpwT9oltEtKI7ewb081weq3KsInE/KzPDl1PRJUzDk39FaRZ
dsCqejml9gWrHrNMfIUgtFpFE2/v/BKg6vvpqO4irqrHUCe9wg1JukhU5/+5
U8GHuLpz3LsYZEkIs1NOJHKWSaJQhIWUSJ5tE2mke0qxns+D4hRnNoyv7KGF
tltvo1DLDkjCAVPm9Lb01jZpH7Me3ejhx4he0em/Z2glj0S74CZC6eiUzSM1
TO+849rNvdBBisdlaxOC54brh9xacB+ZdojHa4oysJOYvX8PvxOe9r3e0RJ6
s+NAHUM+8x0suWDwrqMNziruBW9onYpqLcCS0xRaMOy/ZpXzR1JcUaGucK+r
/35hqDUxvqK/oRL8FEUF39mkcbIXyD4cGxTTJ2pl6enl330vKIi+n8Yt9i1V
63uLgK140pJIkzixzug2z+thg7BXek8BF2R8uYpi+IAZXNsotGUPPyQDPGHW
dQvDY9BOMre2W725uSUVsqlcBdATtl5XgxtQrqH2yWpkhyQxkRmhddiMWc9W
GjDBAHzoTO8WFeTa9hD4jOs/hm5cd2vxjPTm3mVAVKdEeIv+pyZG3yA6EQgD
0euRSU2oBv2FkYv/Acayi4rEYXGM6NJ8I3QaESOsqGGdfuxzYyeaMqsjbYSB
H0TgOKGWX4KiudauX+S98tEpU7Ie9spSFTOhOhztaqtQoOtc+XDUQcl5dLX0
DMfZshGnyUsB18ynUxISAA+ECh+sq/nzcvIIe8KA5WcHuiI4CsnKvInOz2O2
XgmZKWDMfPTW9KvugqfVaKMYPvLfOFivs9zdjftDch9BHscdkhvgYLt7G+XD
eo6h8/SqlD+Ok7qgZm39CuUjZ/+CW08mG8QLMW9aSSkPOkUMAaziWumhvA09
3CQexXtgM+hzCv8pKwFfSFpfqhnPQ27EYiOQ7BuCc+zcEmwQvSW03EVavuPq
C9PLXmKC/G3zf51VmiFRWWc8t49F5St38L91/2YC+uVXhKMeYK33jHzNm2DT
+vdBYWvn7fwfKFtNv90i5TI5sDZqWMdYtsNhBGWe1D7XeyvE8sed3ZsxOAAW
XVDHIokGPLWhH2b141VnF+dmzWEHr9tnBPUwTfn8N/rpQ8UrmLtgdXJJtDxs
tfUhK5bbsQT9oVYJg8DPpWXEmpx2XwHQTdwLmNifbQiVilBFx5Co1diGFegb
f7mkG6mx5R+tWhmFQfBB9ZJdPI+tWu47G6Aqch4KxEe+Isr52rRFabMeRtse
FkN7A2WYy46HfbxnyySwIDLKynre5xvanrED4sCbbCpDPd0C1T7Y/ev7UC1q
u2CUb+MJyVAQCiTRgvOOn7yiMf5HS0/MvUPy01YdNgR5YbpCP5qHqM4OeYO4
HqGXUwbeLbfBUfyJLLhQOV7hlbbzcZ9XqGGAa/5F4IBXy26i51sJPGWYXDdr
Ri5b3ii7yCOBRjfi88ijJXWSu7EPX+ZDpU/BHF/k7KgeqfN8+SlDVP3SFWTj
Ffw5JypSSugXIdZndumDOzDQ94RMZ5WkhAc83cNkddngwWEkiD9xJCU4xUCs
Qc2tdLWZlMVbk6PQf3Ia3AusZtTh5gWPKjVP1GUYkOMd9mrW/JG713GSUbVz
r6TCYnPdbYO0tFOHLg+x5Co+RUJkqSojVvaR2m/nSUiUdGtR9aEkDqOpJhZl
jt/LQa5DJyGUhIaxa7vdbkX1AXInc+S6q2zeG3RKgC7nFh8j6sL/I/iIu78m
KzXndbvpWoaP/JnplgV4u5CM5+yypq1x585pVYxW9z//M3/IdQjzPbN4jFoE
IR9UBdDwSHP4eSwVxqcU8T4+cniI+iDbfXZlHNytIu7/uK3OoKS8MmBcBA8y
6BLxbpihi3hKFiQXLtLmt8TtgSwZbDN40M+4aXW3Xd9gz6GVWCkDXRP54Ju6
csd+Oii46WeJ4KCi7L7a3XfgHiYfx1vKDLNuw2A60S8QmaQto19vJgfor3v0
+HI75lHi4JsxXU1GaWjb1Tb02JMmbmYtSZX3jGQRsYfEu2UX0nVwsIrIKpbw
5fr9OsQW720GGZUsxzqyfQGLQdScEtDuh4UddkcgnVM82t/tptjFc44qn12d
DJkJh3xbRRFI6hUl1gl1vZjZwap1/Fn6Hyl7QWqFAuNzFT637LmMqYczRLYE
3N/mQzhhw9uuWQEETUjgP6QAEiSMXyiIleT7kMfxvxTcIa3V+NN+hfs0HtEV
45eswHsJ6pKpMLVgzI0wag9JuSFQWpWFF5pwRn1ee6y6Mes0Il/D0OXI0dNP
6XugHP8Emg2cgip16EGxxrXUKaFA49yz2VlARijSvaC7P2dcye5uMmW9EzQ7
F8w95Dsny5iV0rf91G/O0BhoNSiDNcynYk/bBcnR74QCVkbZlW7WQy4PdfwA
232f2tP2ltpRT/BWSb/fOUsqkNrPyyRVtip54cYV/xHv9JR2vukTiusJ0mLG
XLwz5BLVW4FP/C4K3WgPRAwKhcpL3rDw8Lad3PvlgYvxvBqVd1zOVU7Ycy2V
bTZPjwx1kZRzCGkDvLLIlqy5/gfoyp3Pk0R96EEHzMHR3GH9JccY7/mxyD+g
cb/CLKiTF0D842rC8Y6fxwNcxV5F5wbemh3wdIFPHIo2mSpql5+gQjhc64rZ
+oJh6FkEZfUzmn/ItzINM8k59p3SRwL1HLVAtZ6/Yn9kVa3tZe14UwcjE5Kk
wnb3yOP2V81vaaRAD+OXDqw7RbKyWbLJjpaduopaZjz0cWn6v6Cilv1LpvC5
YAwW2bCOgZm9N1DuWF0vUKgXaZYeGlJsE5TIw5fcWAZ3RoeQiBeN58eDNTTF
dZu5+ZmXF8d6PXhjkgw2DSTlelWfhudV1qS9Ry5V+Ejg+ZgarrgmzwT0giMD
sykQy1fyBrTJUo4dVy7qjevVQOgc+aveUNTzqi0Fu7mTt0LDTK6uDlLMQuzY
auMAOv1te6Cvq63F9DqXeiSN5hBnA2JcX2ug0KkWM+ojL1uRoTNBU13DONAi
liSiJf2FJwCmSiwqCGoGwlBMCjVBd49etkZ/3afYdPZWbo6WGlNx7BnoR2hL
J65n0uCo9ajJffu0etlyCkhXGusoJqjVJkkqT7AA8q1ydlV/Mm5XxlZfR+f3
rSCWCkouHmM3Go2H9Uqju2rzpr2byeyrh8A9qpjq4+mA9qrKSrge29mTq9Nt
Vog/7Crf6Ux5eQzJ70ut3WX1XGq8+0JS9LaUbHxh02aQEbrrGy9kiwqSfbOD
0uRXW2WxdTtuJV1DC5GJIc8hwh0wXeSjjMlvtUk05xVF6DcM6LP39+Ao9f1W
i0voedadt30HL+sZGi+hfSpVznvyImsJD+x8+cpGijyvmrW0VmNBrzdFTDe/
NrViknj4Eet70PW3g1Errw66voCcNRUWmtplQBYQyptvgYPNH5Xuf9iKBQa/
Fn1ZqrjlFzmyPP2E5nTBju8oGdCCNjbDcncjfaVAJXXt0QgYTSw3m8RcmYCr
skYQZwhE89eMEt/CB5GY9hrwXPEIKCs9Du2ZQuslmF+gPcKVPRLnigdGW9jX
Gu5x8/AHE2ruvEsBnSadSk+waMKPfqH4ZDQpFOwXHNLdesPjzZ2lDms39cMN
0Z5y0iONOWxfz0KvkddhwpP+dfnpwZQIe5pu5g249PhVTKtnpeCQNLT6o0hI
QS/Xqx70H5lTGxRpUyLeUFCvY1VgTNJP7CJ0QcMJoXiLIqE9vuAXNI+fm7TU
aE7zARcwid6b15AGtdamRe+urHJz7vxECHwkoOhAj/LynVGOf6fdSsG6AdO1
LS5mY5XN4xXZTOdAqDgI5860lXkChAf0K8eMKB3AzbgSRVhlGuzIoKvM1CI9
9ofEPr9h42XIzh9JaJj9weLxl4+V+ivnRArb3FFoDewBALYbYglO/5ANfOzU
KaW7nTHZlVNuP8hp5eftMi9T6b8OUK7+mP+fEsMfuFdKi5JEoBTBxBpDcjFF
VMiaOXbsbhK+e++DmS0NaFEluxknRd0tN9XL6k6gJzkP3WRlhrE3AlPe6KJL
q9qCxyhCvAnuz+E6MIubYkrfgxC0f6lbwwYmAV+O4q+IrtA3evaZvCObpsO7
sVvuWmGKhKkZVV/NpF9mXqj49GQoPIMBbMYacdDJNoTcKmbskVjpgHTNnG36
T4qulZ4xHZ26rviGDHcrSNyXJD569rQSD4yZ8f+DP7RQ0BW8Zi4K6c071VkD
2bVVicgSCJrXcU/eLom8Wik5QY9gxjiJud/04c4ZETs49T288UYDuoLEGson
z/XwhZURn0hPgrwYEWAuu1E1+v+zbptGHFGclyIzoGDKGFTpDQvJEjlaJlej
rRvMcvgV0vfwUPZ5QmkWAvqgirkgkeRMt3T0K3VV1kRsccREN3iGhwKHTQQD
bfkAFBFMFzJnnUj6qxHZ40bU/Z199pWF6E1ydn3XJxf80NplJyZPlGK/XA+l
+wMha9NatGx4kX0vLXCuqeC2hLgorfgqZ+00pZbKBBaKONUvBa298unAzeBa
ITIOLj5tYAqxyYKnGkQT7oqCyLk+zGgtc0+SFeCD0X7fU3RUAtd3LTZQxqLY
oW+carkhRXkt9vHV5E8dRkPbT2NRwwDqfJhjef5qfiGjeGlD5Ds5FFUD6IQf
Tm+PZ9IlFUXBNmLliXJycBe+Ie3IPs3duNXdcdPY48ImD49K0HnoTTUs9CWK
rJsfwqONvo5/m/nAoPn24dkzRytjZMRBKU5YTbsJ4ZPFiwasQdfrblpmcvBV
AtH329Y//LG/MLTdVH+u6uGLRLloEcTc8VmZCd7qeNPxJj0k8Tjm8kkcoawo
znqAMF+T2kxMXQWHOVGC3OFmxQtrqP5QR6PfRRx2DLACtWgBLySIjTDIb9tA
jsTHXjwvsvxSsElXzsOK1hDy07cuaifmM2z6dlpdOPwygiCJZ0FgW/tP6jI6
i93Zol3Y/TsaVh1PsFaM1Z1YhWbih9rzkauHN4NwFFI3b5CvyVALZ94riJT+
PJ9rWNmlxiD85C1XNvr4iGLuiHaLJyp1/WZR8OItAypyXZeQhVaulKGJ89pb
6nilBw9nflOiwThCu3QhSkv8Di5YO4cwOMm705MoZ9cob/osZkxeqvjpNq7P
C48CMvHbyJyN1sBcvq4scm97CE6QUJjIf8CNrl17F1ZHfM31JcHXFT0EQYFv
o/5jZQ7HIl4JJD98CjMzp26fFa4RbnWbnBHNt198AlX7CtP4ExaRLxAPtcdK
89fa3wwgJ2qxD8KpNlEkMlXCRErd+ARbi9atR0PpcFoMRuXbHd/FwtQo9MNL
XVQK6L+GVBnKZ2lbZon8Ug5+OiPhY23THfzk2aVc4HyIXdnV6YNwE0ELJymV
j40L9CSDwycaq31HizPelg8Xh8bpk9cieq5U6kIsgWyOxrJoqaGZQLVTYD/n
dRzZGI4ESb4VHimZT5pbfkOnCc4/oisrq2WG15yLW4j/vNXQ/55W555i2BFk
xsq13iHcnMDYaFcEW0MQyYagFKrbYbrBdnvNVojC6KT4npqyQ5A/XcFvk0SL
ApmAnyJpuMe/wnZFPmDP2iyBw+3MlXCPW+gZWaB80ucUHTCPYhP5CjJf24nd
ElxWGT9HsKoGq9u/JgsfRdgjySuZWj8sCgA2iFV+2Hdh0FbzffbopU5pSBBy
jU2ipiVkawOUNB9nkLUq+R++gkPrrgP/IXhpeX9hdgv7jQBXC84CrkABibGK
izqzhIZ6L9mb2r1Jq4xQlecFZ2f8WJZHdcUJ/GrKinpULeq4bowI/Lgb/kfn
GcH48SYLDIYmh4F8TkDizZg8Une1lCnhqedr0MRK9wUqH/gXvxCIhzzQdSCV
hFRjtXC8QxNAHYJEqF/7qqW4JHR9hlr5360XqZr8c11uUyFFBrQ1gFUQQa6i
LcGqCfh+iXMI35Q5eet/5P+2DwuzEr4ku7AhszYzrXeerJ9hnArbBpdtrdap
YIl+eE8KZt0QVEbZDrUOuZmdmCi/HOENFZEnRsvIBqGiyFSisNNhgbHiGAAz
cMI2vDZHbjuMr+0jqUjBg0EvuPJi/hZVXvhtA8Q9/ljneA++hiUCzzgt9A6M
qR6RSF6cfuo0h2tUnldjIyWQ6Ts9ep9lnqTit/SJ4lR76QHMf2BBx8syDiPG
/4Ac5wyTP7hUxk3rctQRZ7XV9MoMYO4+LtWfiPpknTocsc41ydESwoic2Obp
xoUxa4h9Uf9GSLLU3ZPw2gz2K9yL0KEQRcO4sliMFx8ZiOojNTh+V09mrQt1
tZh21tJY6IPe4s4sS7ruepke12R23LXfMtLEY9ptR9dZMFNUIvQ6LkKLfz98
PcAEDrAM1YDrlELIzzHqpCDue0QkbX28J6K6pUFHNL/X3QM3e4cT/fcf0GWQ
28w10jslzATbzVMfyUf+gVYHp4gr1G8Em5+0ovbnZqTwJzjFUi5JFMnrT47N
MP7Cr/KuPmHBDVcChY5V9U12xMbZCWCA5Bpj2ya5VO3NH/lE8QM5xaXEfS8m
CWyXSEYk+HVK++Z+MPGsBOMPplRh0U7TUgZwxARYFiRz9KvNWXJjVCmhhgIy
ci5levjj6YAuTyugwHPVyo7iU0Mty2CR6dFF+p+6PrBAWS5l0E5xvDdlnXsm
x0Q2itF1Rbg3agn54EM9h0aQ1J3yyPeO7e8GawbMbVxYd9sRJQaQmcimFUvQ
41H6La5u5mV5aD3pWP7+GasjCiIWZnM9e6M5Rxf5fHdnRxKpww7yNc6jxW0Q
E57bdu9ulf10Si8sqGvAspaT6mP92+GQQaM8Nw2BNSWZK7qPfMjupwpI4NEK
jsyzOrU04RtvDU+eTD0+P2CwYsvG+jQbvfepNHvaiZ9TNbxyGkvNGcFFJMaU
/5AtbVWrdwo2F6qvqnYW5E8GWLYZj2Mmv1wh5mu/irYyLzJAynDT4Zb1nML5
v9dCAI6jipWsDxMu669M1Ox7NwH+tJUhhxsMTokN7ynfJ9GEGWVAv8Ztr0OK
CE373U4mAgO7JBDSiPJoQ/TxZViqZ8fb//QH5szv+QsRpSH5W1yp164cQ5Kn
aTBbZlcIvLTbHefEvMOes6SwnzNzzth22TMf3BtlEHUGtENlyYnM9k600xjg
yRQBHyPUSSuom0cGNLw7S50Yi3/HSts8qkbCn1FaPgRJL7Yt5rWwl9Cy82IN
I22Pgu7OeTM0UbGQt3imBUz9j/AHGfjBjDMaFpLs4hrYVTpekKgUuoSSWgoO
zyXcAPLprpP8syI4m3sE7sH1s2CbTVX2UJi8v/zrmOPlqoF16E1CBfsQbaF0
xvK/FMo9598kUhY9XQXKSln/UipDVubjoMFobI971o33lnNb4UNmn59GZ8LB
vGwzd/m828GMwXNHXNnc3NQOfGF/qbLRufDkWPUr6AA0pAeK+Z500pnCFve/
7G2JwVQ8Oxnw3JJeRQjU6vCEm5ByNYLY7orpozQzmOEZ6AfE78jnDt/7Pg2l
QycrksRZvAxCqcGMrjcLHyItcn7VYTT3ZVY23XuPZ6w6f5a4VF60bJUI0GWm
cLXti56YCHqrBvfm7LZOnw3oaUsAi4sU9pGPxe5nI3SK6G9z75211m5kSADV
UsA0IyPSoKfCpxzxxKfH6Gi38JAQ3jOz6E61ouSnl3airP7hNZ/omUKayrcH
hs5X7H/HlcssWlqnHZ6rFaauTT0adkhGiVvP1Li9zba+SmwjWfMgSUUIUuon
Pnf6fS0hCUMZgVA+fBeZp6dTYN7wLYE6uXhyOy+XcuXbINto/i1ofvbZj+nw
ZBcpxTWlyKRGfch4ICz+I7e+v+IyXLKnYBmz8R3Hsm2gH9URAQrHae17c5XK
nMlZX8NC0CFX9bT3UaHSlXE/Nv613j6RC2nO+GsTsx/I/xSs5Uhm+x1SyP4j
lR5D9eVcYoOCC66qK5YYpH2czFirgdQzP93PlpZTFKLH/dsyOjCabj/8niBn
vqQ3+vLNp0FblX6Ma476N35bjM5Uk0aTDw3pkim9m7IoRlGE3vlMRkj21tvu
PzfoLVAG+MMSOk/ePcrIV8FT6400bKsJ582+XsddtwdpfyLlKD4HyJrOI6oA
cJCCQdRNvQo4ZUer5zXfRxCqoD8VPbMcJ2ezQc5bZPJdLDkDfexsIg2LDccz
ErqPCUOfmCEUNrknA/yPwmtzRrhJtaZLqH1MB3guwJsJGxf0RCBZp7NCOjD+
+eTlMmmh0a/sTKU4l2N4wSB0Z07i8L+CQNJRMzIsP1SQgL4bQuW/EON/7+oe
zFxmfQoX3YUTow/DviZ479/nG9BEN2XN9Cu7NL39JtnsxFU64LoZoBXH/FAm
yVGZR4t/SdYFx36LHEizvjRlBLNdTT4FEsYmYCuXJmZ6KbmwG6yZmF9YrIV1
sWgAIPQDfokFAGUorswaKvnpRwnJQb/He97TmPX4tTxka5mSyT2dsFgTMgD0
i++u3b+++e/pReKdyGNoE7ZO06hrcSVHdNj0Lf2mFkSdwEl1ZV0lPJIUu3t7
wPBH68vXcnFl0+qPOKs1Zi3oclDX79N+eP/2TGNJgSIDLcmHDm8AQz+H2RrV
XD0D7YTqK/2d8LYIDy+vg3ZOA2cq04j7oTGLxiAckjHY5NnhPFWvu3TYLN0T
vqjwWM1mdBEHWkcSg51qfdSg0mSY/r7Kusrd2x6euD/2gUtKgenpsx2fLpMY
9/6Ilul5Zl3g7YtL+Teuvz1/dM3WDHH4YXcVkB6+JwlAjciVjdA4dE4SGHw9
MDAOCJ+tpmWGALoFx/YGNRnd92NHSsGGlKL/b+PEVmORcNEJuabpmWU+8F6z
q+LIyft8MPu8iUutoqWZL4a+LS8eqgzpAJNO9HVJymVB5YNGklE/eYEL/3GK
Z3b2uEHRQTcCeYhua4oH30QE6cLOk52PBP+nxPeeyc2GZnVKa6AE+jLDc54M
50DEjW635EbUg9MoKtdpnMeB1LGZXpsOFJrzC6TcB7qafsBoot75GZMKBx9B
enFYc3ggSwW+SFOd7ib/VhbiIAH0Xa/xT21IsJ9vjkMqXfgSlS7Vq/FM//la
zJ5/OXe12DJv2/eXAzqPBtwdUD2KSLkNSNwTdw7cDDxI0fTViBNnNxZpPwyf
wu6GAv5HmJ2BKjH4WLy6Y7o9C5LYrM4A49/2l1EzxtAi5wK3nTGJnETA0cr5
o0eehSvM5CALtHbjUJheGOLf7SzDrOPBcIHcGrtOZk+0ODBDJ9cAaQ7LaGuM
QkZ2MWI2QOQKGj4+Y/F+2KIIDETUe8lJapfh7d3/jDkZJhZoEcmhHLw+SKLP
ZSRYFPVkYSg1D7L9sc5R8CCY0iaM+hYS3ElGQPF8gUyhHQQeiImKJm3FCqpt
5kjN20+zqM7fx5eEawGr0bp8sxfP70D7FFHBr4kKc4sYkxBOhP91uaGoccLz
9eMd+kD2YTXMg2nVXRnlJKAgC69hqRG1MHvMKj0GGD2amQsgdddkFnL0fG2w
534CuFIYP4cPbJ9vwagRyjAUXCTJ4fm6lmhKzFu24uE6hufSXdGyxQh4/oG2
ny+wTANCyVtXJcNJx9EgzzAnItwKkuJKgbc3xb4CXOzJ35pt8sJkcWsmOm5g
Z88exbJSRVpTMi7ZZueryVI85Fmcb9bN6REoOJgLBsfCadpA+Y6QmzqJN3s7
l9WmMaLcxA5wia/PeBv9VPYEMUWdbySyEBPPn/MFofOC8Xh4TbKwzINHFRZV
x+tGtPuj+joCRXOBAt6SVP35W72f8KhLdGlx16pfuiFPIJRdjAmbO/PEE3Ad
ujKnecixN8K2cNv646QiL6mKiikVs6CmgG79fEM0Ou3eJwzRMXXuHxtj72Cs
m+LgyjFx68iQ1U/yjEwf5b5piymUOUEGPTjA954sMJZl/F0R4ROb9Nu3Y1ut
2X/z/NcGd/39PzRE3YDGWqDzfzm/F5OWCLrgsdyOwQe/Uhga8BGy+SYIa2mw
D/Hp4Iq3QpB1pNHaSERRHxXFU/vItn9TZwh2hHXfLGfS2KCSXYuji5wCfHw8
AKysvd4rjF/3CINRKqTmHFvRiol2JoXWxqlL/AgLTdPBUnONbqO38K3yQHbD
GXpgzFD0U11Vp0CaklJpBR8N4WfMlA2Hh6/MtSOW7evnU08Bxs2OZRvtDtr3
0KMyMfVP03V4Sifgxu8kXRdcf6vZNpafC8cPmwzFTqX3EcdrTgaFs1UMB3lj
JRlCF2WOEB6/EKedkLeTg+wv1CcvJQLVcWObE2k8pUAZjTHwkY7alhBBqCZb
Q1PJrOabqwAhp+d50RwzLdTnbHSq+iMdQNQfKABK+OapFLY9+OdLDwGLTyh8
2wlW5/CdPqsX48PoF7pvDS312WOGyJlXlKDArZxUC/u04NOdfH6p0ndyY4pr
Za9k/uSSPNFvnK4CmCJpDHFF1qxJYNS3Y24rmbb3rVnKs3PBYmlyNQU/2R1a
gx81SH9xQhkk7rjzp1QI75is00xM6kfhlshA56PsEd/oOHmmmncCVaL9a6XQ
792T4i5m7uLUrYRhpOvW+MSbEWgs3ggfj3YY+60Zi6ih4gJUvgoWdfBQQTxM
V0ZWp3noO81+hQ1zNf8xpJvDaqoq+iNDJpCKwh1zKT5fTHD7JwLBtQanIB9Q
a3mrTnjn+5KovyZlW2rTt+5SmsNTG0bQrv0yVVEnQ5+6cjTLokkdvNfsXP7f
dfUs0TTmqV70Yi/Rxmr/iIvJ4gMHeKpj1MPCicMSOyYkwTygDwQwkPwwv5+l
OasFCeu4zisMhBSkKV4P7CpXikwV4dNaBRE2lSjC7M69Q6Us6JdDLKB6pvh9
9xqv7KTtUZcNVYAFWOdOpCse4FddciAHVRkJZj2q1JdJRh+yK6cZ4EYOUrBj
tvxqixhy4fdb/Czjx8zmX1kyCTtvtclLhs8BNwab5+V6R3PFEPHLculpX9zE
8yciggwHrv+1thVyhMPPHD+JEl3gslwVGOppM7dWaODtEjTkApSMETaTLK4h
18nJaMpivUuI14okeS0h632onRztbqmR6adlunj4Oxc5Sd4upCZqtIgdCWEv
291h9SOEGwpXyk0vaCeirn8h/nAoEuvXxtkGg2ODu9Cxrv3fojmwcAvf1FtY
qOPXKToy/pRDChJY0OhXjxTCSLgFSA20Ehm8L9qGaDtPU6MMPMY3jGenl1w4
yXLQWS5BqGPWs6JoJt0P1+oBgjYOu9Fyb17D+C+WVp1pdWUs3mjHTwl34doh
Dd/i8zfeKPOzFWZJy1+WLvCfh+x7Uc+acycXbaL7zROEyFZJsbp8vFq+fP3w
9g5+qQy5/PrY9HXL2WQiYgMPJCn3rL+VJJktPzXVXn6iZ+spQwrOv8c0AjDh
KRFgpQsg9CAmFE9H1/ikcT3upQUrGfRl0/MiNYPZULd/50rj0v/Q7pJLD6Xc
NX5SMZhT4KxABXYP/bkllnk9AXKqQLom371n3WEJbbQ3d/nA2eFDuSA4MS3n
Mgc76GbA09ODxe+X52aWdfud46Sh3Sn5DAXzNQhbFzpL6OwU3gIfJUprt14J
Ef0oG9DlGoZEiVLqBLfVZqdxoFkF7MJwOENmdYvwMutDObyAUZE5bFYxCLRE
3xTCtmjJpuynI9WBnVqv/h//xYFjRTIMsuU+9Oe1KttoAnzJrU/DC+t2Kzaj
yo7QKdcF8cCyeCGCVjsSMQYAn6vZX7/Lawbx84iXrCPVhSc/MLprUyzHYLAV
f9ZxRJCGHNVpmdW8qT3pc5SDlenEiQ5LCuIRzGoOhSvPp8xNCUa6rFG/Fo2p
LoxGjBi5MjokmpeNjTO3lY+gHTDFbvOO3i/qX0TfPbjGA/zP8QznQEpX/sn8
puf5+Ei13urLHkHM0PNZExk+cvTHVykm0uMxPnDgy15eSnlgbPMz+bSYUeOT
Vgffvt9xatbCTN9if7uWClZNdE2NgSofNYuv2Cip118DXLeGSdd4HYA4TfJp
v9SDuUHdRSDuRGf0C9M+bSWb2CTZMByZlDAJ7mdY358lE4vpvUeWPWZYQG7s
dAwzMFEpOCNZQc41F2uXdojCeez6jj2pmR+CZJ7tNkUm4GVw2EF8fL+yxCiq
jgF0TmqtSFU98deHUrfemMDclC6i714n7Iez+EPx6kgRopPI8+wcrWKEjaog
PGMZVEzpEVTRwOZhh7Jv16qY2kzCDulEslJbO+SgoLiBWmmdrJWThz0WfVqP
79pKHd+Ahlv4u4qOpU3DLfxAmlryBpgARWwBT3BLMoYBDQspfSvj6Wj0qWk8
GG4jvrn1d39REyPPCN7ABE8gWXkbWJ7/27lC3cum108ir/OcavcQvNodIuYf
7y84M5MlrG/lfM+dJ6GwwEuzbK9pzYlNnq3mmFry+Mdg3dnHjbrfqwTpI0xO
2tEpIHfX79I5kXVBB31Z0UPLSe640YLf+hqcJlAjEZxd2h65ohOy9DY4SFWG
GDy1UU2iI5cAz82ocqhdgq47uXgMV7mf/NbWVovDl0x7j0mADr8WrBEgLO/B
2qLmoy7LMkXCRONgu3n9RJAbkl5CR0rD2j9JZF33qqNbC+XTtE0g2S2HJu24
7lRp3dEympS3uHwlsuXO3iBDeKyCzLpDs4HpvFatxSL4Rfa4E1UVt5nP7WXz
iOWbpUVhf/3uKmWZyuxamzoTERYr41TWjiyQMp97qPtKNfnkk5PDTyLATeKc
QUvUngfGNi+Uuvjj9/lU9uUsX0mq93KYg2aAx/AQEUdC1IvmQE5JwngomSOo
UDBQwBxqufCMZm7T1/o6S1bF18foWvOVsogy5claJnO0oEOud5SNKrumYIf+
r4ovzG4VAws+1YwoKGppXzicL87nr5k2kJUD288Mn3/YKrW4SLQ9mwEhYrpO
FK1l0Gfov+fHyhuvw4cSHyL3vzX4c+DTfKgpKIbw3TyQASkPjqEXyqUrAY7S
mLz77s0mlWjLjrrHaYFwjFNkaqEym4pjhKZBZzWQ4l7ounwRxlhD+yWF+Qju
6ziSMM60wZPeGpKf/1dNvKgQC9sKErzSbHDtGEqThv5YDgTuMOWLeUi2oErS
KVv6Q3SDw7tfMGLFnIR79KzVdE+OJ1ZtjNcOMThlEi3PbG7UuGBprjiFEKUm
HdL/TkbujeHvWz+tb8BaPIzLZxOMN/+QJBDScpHHc0dvE/XRMDtWKFvnY0RW
aZCtl2l2adZWge19XM3ySDvA6FkuJqlzzEnIPZZ9xDLa9jhggumlvuZ2eyJU
ZLjP39fnKeB35fa4vORjQiAxFNlOO9INggker/FwFtdBvWVljmAbsML587+C
DcRWHY635m/WJIHT5pTaDtWSMFHlEcBw+isNZABHcIUZ8TxtpFy+/xDZYRYl
bGXMI1TEeh8+OOmk276UGrU5HE72O4XJwFBhPgTJ14tgDWwDAfh/OVeD5utu
uXW2iI9+nQDpxk4gsV6AROxgD6CfPR+30YDxtW6KQh0au1JxvXd7HU36yqtF
esmr7f58fXIaEUNVLC6jFV4eb2dU6hpdhl7URYWePBASdRx9lUb2i42Zv/49
IW26n/OzMAiKXmmneCj6OSlzaRqT+EhIEbHEmWgC01CuGjgvK1wQIy+MrhuR
qOegdLokYEQVJKLakJW+70YY8KiwcGkIngM7LLDLAbp51xrOhpaijsWSn0ip
pqCEKiPBom0PtE+i2G49kV/W2P5XxvImXZlfHYZBqU8QSqu0BvZuRaS69eOI
Kiorm/dwV85stRBWEV3SCJhPSKQ7rmVyCCxieAPvo+3nf/buZ0g8Nk7MASVl
xV7YXYDdUSYdUrTPdaRCflQPZNPi7G1Kn9TRt4Q8BjXEEV2nrmOTmfbw9TkD
y6CfmY9TK4VjZab9qQnNgc3by/qD8NvWE93OT84xyBeU5eSxhzqoLIhAnpPS
iUniq+jagmc5WYgNFQPpYMNrxBTNo0y4Ff/VdFWFbNtzTUDo3ZPva9I508db
Ju/86xOwUFB0xJO7RW9bcAA9NmKgTte7yNYGJwH6uij08GFViE2xjgFOXw+B
99M0NfukWJjfd/kDEBc7ppUCyDIHfGAclbPA+XQsBMWRmia3FD/V7YUgGWlG
G6/3KpaaELKovrtrQZ2QONxUXXB+QXx3L3kcuK0bgLsVSd7OIlfam0lyL+S3
70nK6UO0L+rHOuLw0iq33VAX1SM6T2SCDMvuNK13LY5QwrL5v4lEVCeisvRD
J7/3LzTbERCtTUTcNA9sZ3XOV/MQR89S6I1Rv5BoFxTB8hAYtRp2WXqjfGq2
n4gZQ2Z0QriLU7TI7PwNIe1uplSSmQSg6DtRhSvugCN2NW4ZDz0cGNSDdwNS
Ad0kgETUYu0vrGlDBUignP9n8re+qv1bhQfDhPrIZd+o0LbxgVfvzfgRR7zk
MLkAXqwzOAz/0e+vE8UGPhsycXnxnxUB1PlmXI1jd8K2ma4KiOCpv4ZJ8J3S
dugaB+BROsD48UhwKXbfbbqKJYXeb12jJq9ZKguQl7/HYJW59oYv3XZH+Kdt
kxLkF2yd35P3ZC0aVlf9b6q7NhCElJSDouzYdQUvylyA5T0bdyPQADO84wDK
EeVPCjEd9K9vX7VWU78Bz2pH4wIgvH5GGQU7VtkeWVgUYXcCogM/h8/vzSOI
Z1oGcCTM5I6MqxVMB9hqmy5vB0FZAg6vwVPYcX6i5HmksdG7uIh1bG+EeuHF
2v9ggczQ6+mkjkMWVVcSff2EtdUtn2YsxEvWbLTRlyMpQKadWfLiz7EwF/1n
7QJkl6n+gNJg+Jmriky1VbmeuggaTfM1BtYDg6dEmkqTjdHF6XlBK3QKU2Th
8pVJQOhC7AFA7SRLKCXz79XP6Ah6ZyKCD+qn9Wm7dY+qlBc67JbAznuDiPlv
bC1hblOEZpyvQVH7W1hNq+n797u5zX1u3qhKyF9shVTd6mrmXM7fcyVdMG/N
A4/h7s5LEP4qnvaa7AU56e0vtkGjoQj/4naOVtqjYWX7Lv9FPYVrisA7x91/
SzOKS/c0ozcfjK0GDE0JmUiFW1nNh1eRGm9u+ocfoEahUXxYCq4tIkZpK3CA
rLlmVSefn+mVaV1WGEwg7aQwDFXvKiWEa3hDrqg+nNPFu5rbQeOFJNcuqm75
Oj1OGhM5OWRDeZuBjkZxPtto5eeyrZtF7wWb6HefrKqIXYomiAFc5PJQuRrM
YAFsX+U0T7cnDR32yMq71BYKqQY0gd9uHLw0ibtZHeCc/MsgFhkOTAOcJR2J
IYJfL9pzB3F01xpL2DgzlUawK3RJafLMSJ7yIa0F2jYqUyz4a4BeDuxLA6U0
XSt0ocE5fFw/qttmUPiClhLW75q6IRM7vHTna1PnH989wJ7RcGOfzIpFULtH
lVJhHG95kkSFZx5aznjxRmHEwufOKdNkymVucI2aHh4kkwmD1V8ZALHAsLjA
7hhQ7TKWe+Zc9Is37iydFxqktOl1+aITe0F1pFr+Cl0WTJtg2l+04iNEgQuZ
dpc1fCzEL6n9pXSvl4yNLS/yBkfAGoo5z6V0mNwgwam1DWAsTBgdrcMqEFXW
TLm7xpZkNO4jfyqirrZ5T4DdhIFfZbEb8bpC5JvQs7KOqXy0Akc01Tr01Zeq
JDFVVgeJeCwpRs35jGm5zAbwiMDnj8wOI6Plyg8Hl9Uhn0WoaBI1+eWucSYB
/jFZZyesQmVsjk/jhT8yN3VdKc9slxISA6zFN8qZQ87ejJEAfz7ChqXFMYT+
VP0iUm4Sl7mnPriVUVrXvDOTcW9IQfHvQgXWM0d8+L0SAWRTr2QGJaSioGhq
mGxjLReMJTBOIvfoSWh7SqJ5KXp2xYDrvNytKBJeMVP7bO98lPdjo0zwNEjQ
2sutOlP+QMbPlwHRwdM8s8gW95DxWatxHbP2kX3rxDx72sUKQeGAVPfQrZ8E
Ab5Lc7I/7lTMbM4pRaVNzCek0sHlKvcB/eFkWzYItOHlzICuWeCRQfWBUwoQ
Rl8B/OqWIwu6xMlewM9EFIfQ+OC4LsyBnBvaQ4kez3z3BpiTcu09QLczBS9o
uZTSn+ZHvjmuE4zp+1iA3/onrXokqSel2e/J69DuStraqyuluY6M4TjCHVDo
CcIPqs+aNMFA94n7dwqIk/hsXIjJhffpFz+odtxRSMVYnw8pDDVBnDLL4hzI
LzcXZ6w9EI0fODGyzhLdDZ4AiLs0E+FUc8lhWt5+SCmoPVKzdV8mnRYEYu3l
RVHdMxU5hn2WCGMWb1Q9LmHKcyB1wjMPejDYQq24xMjAZz7IQD1HP3uhfI0+
h+BURqZF54SEuyYXtl1Ilfg0KeqnepUEY3l+mg156Fbfy5H9Oy6MRPSGc4FL
63Z9btaD3no+7pQrDCqE/Evh842NCb0aNSL34kZqnj4CgrGtSFqfJqGuh5sb
1BIC2nSRudAXA/aIDdSiAI49fO6Dzbgac3ZbdP15jVuwUCG7pKvdSDTxqd+9
BQNfzZ9E0wTu2FZUrRvd2ytYD7uvXijW3TZK2jVGQOLlkA7G+NuL2ofI7xzs
j1tAe9WABgl/llj8Gxc0bU5EnfK18YWsfgxaOoLgMHFh/ItHFPWaaZxz5aC/
ovk1FWBEvJXMKbS/m57uh3Tdlqd7DJZQmpMRR6k3NceWq+EkDxgdYVQ/gSUb
fsGwu4BkkicTX2gdAg+qfbMazK2VjTCrj4mlaQO9Qt+hEPPk2VtOcZLxh+bk
p+dODDyBzfsuonj64aqMXliFvbvTqDqYIUrT6LZl2iR/v03SgMxu1BWrbTRn
NZGl/t110NHaTYUzV3FdUB9Dj8rO/CAaKsRvJn/Me/GWN/xGqBP3Bc2SuGPQ
oaXNgO8Wphn2QBsTFPL09empaV7BbfV4CvQWFX/Oc1wSlEzDxcs4jFgDdoKw
hl/v1yd/PiTfuK7Ht98I42LZLZuhpbMyXhVQxNrwEWZk8JA/qYGs2otPKdwM
WDIdcbK7bdFCyLUDOSaY95Kjsnng+h5pfjNMKvPPIinJ13p73ebEBlbrlrig
KE+95J3uSBnT/a7VMdQelhqpv5n6WvYArZesIEG+HArbMHrdqCK3oa4RFCZT
f8gf7Huc5J/OPqRN4PpyVqBKXn8Wl6Nr4Bp3k2Vrhb4aZW9CrvdnWS+EH2yP
p1F4Go7Z4vUozs9tXmLOIAC+UUavMkjh8gHS3WdfXZ/qHkjYxi9f19NP8K0Q
XvklFk1wzFMlYYNfbIlEYqrIeRB+6cbq5XvrFHLJApKAGqxh7XJBwFYCsM/q
prjHoOpgK5/pxeUId4hyMncDe2KlzL3mnE75rcTiStkI+hgpTe38cFkge7zo
qe+887QwK+65K8vJpjTKlOyrsdpwREe+nJscnTAp7LmamAfHDH/SGjyQ3eBO
l5L3igMLyZI6NudTPwPE/id42J9+xCgbfotyp1G9afTwJp635IHzI9aLdNuz
rIZ0jbno4RMqLGPNbcu16KfEKmFIa+RkvYbOvNLclvO6UYG1AKZxSeovkyya
/L/ugWwicS0uFHFBzAhpHp6OCkp6Xi9S5Y2HkPYq/4+dzWPnnu7MwIwrQYSG
xK4afOgboKloooVgJ3DpFzv+pZ0RcYuVRq/HE0EOZc/DsmikUMGG2xRU938h
44HFZGjB604psbIa2AXT+vRp3FydAQ9wsNbOvU1SUD0UDjDxV8yjO1wZIrfh
pDcA18YrPGlJ+vVnep6ijerZSr95AtedhskELCVKsUuGOz8S6+pJLkqQwaxp
z2Pw1wY9bP68X/k00F/Kl6IIqyfuGnDbNZw4qCFGJs4Lh2nYU9JGXm0z4zN4
pvfFg+H6yDf7Vkc4/pen3xJFkq9vESSRhi2n1cej3fsospiUbXkWRO/TDLQJ
MuduBGuYl5tqpStnocwWIe57SC3R5cTHFWZMF3U+Bg9P+X7hzq9Miza6rbkv
8zox5nwSRuqAnW85YbcEzCaLoFGGY49wUTsxUwdeuqEga/vSG4v6ViWHHaqe
KpXIf6Ec5uzW80yzolttGSsu8J7ELrgB6VoElr2ID3LdIvoDk4o2rqCE2tZf
0s8ZoFXra6E7qsw1181oQmjLbWed8aJ2zJVkx3yVxQn7k9EgE970wYysFbdm
3wueSwI76Xr89w+bjktFagBtaupW2yCwIsAD2yoJRJvnB0Y9WqvYOxjSYZZa
FoXbC1Adj+U+3cH3bpigsobLz6KH1f0vMKGrsOCiALia0U3rf0Zz2NmVdjPg
sX2ZU4XI30MVaEewyh0mhknP0WNh7rC0OEA2WoJ59aLRaJiXuI5Wb2RwXt0p
Zl+UUi8L/EYKJxS0sRqAFO1+h1xB9EAIhpLMUKy1dQZsq68MRDGSIfObV7UM
5x/hShWunl9IDc48tkzf1sLkzG8LN5R9chfbYgDxAbwMK+9ozPGzQnjJRod7
Bzau0bDgQwEvClJ42rroydbO+XPNdAIJOnaqzjwR24tc6sWA4v8Qe+Ims09w
hRn30UuBzmRmbGHYB0BbMdyKwPxo7FBNVrZAHa/pOmIgQF5xqu9kxIcumTKU
buBRUGE8Xjq6dfaglcXnUFT5uWfJx2X5mKB8mcwKSVgQgch2xxNmZCWjz6qg
+qb4+Q3Vo9et0dHCdqKvH44MXtiVNspP0mmyM6rWzYRDh/sype9ULwvSDG+b
CnSW7tL8W70CJmTCJNmL83ITSZfzoJ2/KXAcnDpYRMTmPlhggvYpJCrKeFbE
QEa1qt1Z3HxAJeegpkut98e1WRrOsXIIq08Y1GQFZjphApdlWkqURC1z3eEs
RgNw+4BZ2dMRwlQEAy3VMwDupawMt2zDGCdwXd03qGCQcEnuKg4+AK8B8vqP
BN6fZuaTrnp0KHXcQyycO2hyY+wLLq4dm7s6H8zDSKg+SYqekC6o9ousRVEi
/GfTj9Gy8cqsfrey4l0kdzuJnlk93p8+HDf55iwqAcX6BdeUGzqmoSz9YrZO
QRhNmh9yNVCtMGg3+r1IHGqF2mKyT+aLUtO0fK8Qqk7C18nPEuGr7ViyklAn
aSL2dyTgV79o62bjZMWHY8Y41Hmr5Q228PeBirwWtlqCTGSgZ8VfPugk/EyA
cR0tw5fJDXhrXryiBqaOiy/I2TQ9feuhy3O8iuFRByZVRM5OqAflIWG3T7hf
Xy4CKvdT7LsyAcqdtzOC3mE70qSqsgkUpjMzM7+PBCd+yGvRQNh5HuPg1gDL
wmBTMj6ivcaDoQZxvbYoHdywX4WgtQSGITJGYw2so2XGB9IrgePopR+CnHqX
wd5r8YgjVkl316b6l9BRdC9598dlXzwYFPK0kECrgEc5N+QERhb8fogJfyWf
Y885rNInFiEYYGXkawde8lrA+11HfTGrbsKC/GMKY6fHYYZRZISwcV1zmJaM
QYkdgTnit4fhQOME2wsGCO7vcGRJvlBG31l9YaazQF63VWjFtUOCg/Th888l
D1FOxQok5drV0LnBsZ56MOmXG8CGCFxUCpCR3BA74QU0am1TaTPnDKoDCJ7k
rHQzjPUEQsLn6JrJdlQO2jZPwbl6tNiN2Azbmql2GYCP57ym4SWHlqPhY7CH
oCBz7Qaq3xhhqGHwGIgiDmVRKQ7HA3mn4cDxsYMaRiqHJ9w3y3gb5HN/8Dlp
AuoHJjCPbcjwxo1EGVW0yF3WAxysEMSmWl1iQfeoqAAlEP5G4H9duecZnJuj
5ez5pQ44d2mClAFg+bh+n3o55Y3VMx86q/OkCopN6nMCGxSg5mtmgOJOyJ5y
y9Z0dglPrHXn3Vlr112SU1RhvLtPSAqVSyGSamsQmxvnugYXRUsLZluKhvnq
VntrKyjntfkONzLfEhHh6PEXLCVywjWIffY2evX0kfI2yZNRwlj9L04+IBOS
0sWJa1VHRJCvRdJHdMeIWktfOtJPVbnIqpzZFK6xnCH3SmaAiTM0SXu+zw18
Px1TETtnK1s80YXl1MI2IuMtzvcEIVNPz/MFqIZhFzQC1Cz9Yq9UcVaRSGRH
vprm7Ge3LGn2pLNfHiq6PAh5D3G48pizTUXmmpKEMq2Urkldu9ZPpuWBYIeZ
Kn4ntPnpECxFk0iBpDaVqnVgvws3j6rvrO+Iba7K9C/2h/9tiRmHBC3rT/aq
u8tWM/NYMOQKtmD8tfNs8Zs8R0a9WbNBqEtcG2/bdjkaEXaE5hXVftZPfsd9
cR7PZTXpku8bVfS7kbckhQ4mR6tBGEBAa4ttivSXLN6aJKkk3Wpo91Dn3p9g
aqBUPOwb4mW+L08idKLHCX4Zosasvi7I0KBm0Ho+C7f9viqkajFuPZUpNJaA
OpigM8pZWEj4JaNIOmHDhezM7a1e9BS+H/yvLug1B0tD4eeVz4TNWSoPPEAO
T5m3IA3wPM4UB0EdjKjPm9QdlurKm2FgJH1bMq1ORGU/KnTe/Hn9yPTZNLHP
nIjb8d1Mv+U5rKVAjJPypcVfEIf3Z2BpY2kOMuHN73CvXYCQXBS++o8tV2t5
PbOSe/PeKRFpRmTJH0uNaDY4iVzYLnhTxrahs2R42TmaVC4NeHhDMLtSC9OV
VoNIUPhjlE2F/Ocau0ldzOntW+ac8DjCNY7FwRyAMGG5LBm0CAfwkkGQL8ax
xj12ASsNl4RphoLagyzUQYceTfyJySrY8PgXd1LmU3S3CTAnDACjdunejRRP
73gsi9tPLv3f+wtFq59Ue0vDksb6LsAOEYIAxODbn34y/+CO4gCjjgJl0gir
hzmCFbI3BVvLtyshtQoXedhlT9rcwicZN/bZkPOWRYMELlF0HKGOKqS+PGNt
Gr7Jf20GUH0neyU0/a7ppQthdpxcU0wIlvDlQqaVB8VrGVuUVBKP5fh/YQYv
5QiVlUVjG3DaZDJiP4y9c9zsQnBy4geHCPjaCvJAh/LrZxHM8sm7Ki45jNRp
2mf47GtLgr8LDk5+e6xpAoqNerizT5urClUNUl6XwT+d/AqerslCcCREJO0G
bNnj6dYWGZALvIOwfGWvOvqvixLQHabUxtYSHA7vLHWKfqlDC1EtJw7xnfVh
1bsvAmmTEghm/Wd23NvqT4kGfQqQq1Ck2whlC9bXmmjGijFyT8sws2G4O6Pc
9L95zMQCgCyciTYNJBPY3p5frVs7ZfgFvEqPTaybWY+tV+CQzcc8RC+dWbX4
Bg6JBHs4j4P348lWG8aa+t56ydij0uaCVV0Xap7P4JolTfHnz0U1G+ldMvSz
jFDL1IhFIiHhJ6dIp/lw6GHImywkCiJ8EowLlHJfdFd/+FjFDpu8IYr9U1v9
sH52gE4kC3mq/9gmwj7AGEgFuR4Wb5y7+EQdq5Ksqxor7XD8JX9k4p0LAKHf
/4lyldb6EP2OrnHEUsVsBP/ofo9ra/vuUBk7+otr08lSS2YsEyN4Lbywsn+T
26CTZG5XUaL3BM/8wFniNctA1GXDvL4/4MfL31g0R0hq1ljKavSDGyNMRkl3
7We6vMay2taQg87ijGktmlltrydvF9glNzv+0bb/6NF5lsefGSE7f2SdwBfa
GzJZS26RIdkbg8gby2THuOQE4JirB1c40S3DaVuxl37u9fl8EqmWgJ/Kpwjb
SKWd0pNprkp+1dBXOkBbrvBeQrwie9S7abQyyqWpqUZeE0yTdUzQ7oXLfQoT
PhYwd4wtHX8bwVXtkNXYn7ybO8zNKcwBeHb99zFmjrGY/qwi3emu52kuoq2P
978wio//1VCstQWCSgGlpQaAZMU70G+W9eg21DGoqPEYpnSgz9jRWAGMbVPT
ycYOouuVHoCYjcpUKKih6Na5YiNuawVlB8UEXSv0igpYumUb/i/ircJcLBF5
D3RCVqLsd6i/xA7dc5WHwLqLAczjRk01bb7OQHMvVmHsgMKgEuZOP5inB5C7
8PXRrdclaGnc3M8N+xbWpLu3fDJA0WzvGQyjTtgYi5PtSI0tGTT2fzxCi7Wm
2kNDn3CzoL4BqcnYBDHfKdeEkI+/N4wIMSDnXzsbLjM+i6KonEJlL6Sq9NvN
MJ4w4MOWXo9QCSXau1uPyj6rxlOeXUs5CKIziS8wd7byuZSszmtm820t7QBw
xHRibDSkZgIrn5MU3NWi5/3mjCFBMB/SDu6SUE6VDfLF7OF/SXbwSiYNWmFn
FFY0KgQeVc/531KWU3Rm0zY4sCnAhMQf7fmvwPhCg9jPsvB/ufs2KqNEbMNw
GtqDqtW7lxHFgUkph94wz0Wqsg3jfNEbVkxoyltcP22vtupoGHhl4uFGAQLM
wXPsVbzDkEf1/MpeZSHwQHP5B4uzY8quo6SUtofAMK/OE5eqRnPxHstyKQEz
JyRFOlnq+SDaB8wwZ8v7DR6Jz9UdiyzggGsWrT/wMLXtKEQD6PCBOV6yE+0G
V35nefcvvJwK2bzJp3GVIQLqpWKt0eJaFe4Uc8hKlGaGE5DKgaGiwP06OvdN
gXznUXPvBi2HdO3FCUXtMAH7D+688FPPSHiA+u9WM/Tz4P2paWRg73rUthin
mVgEwCI2PgT8ZQixaZLeHdPV41Ah8oPXfzMgerV2WQfPeKoIOnLt70SEDU8o
wsflikNKRNRDoZGbA6lSlJT+yjTBEdTBbt6JQjNZETE3EcAWxMQa0KiCnriZ
mkbdFg66eP/oq/0yPWT2v96fxCbPxYhxbZ9fjCeUyb1i84pIbLQGK4FIQwFH
XTK+UTYinSrPSFge5Fsb7kvQY3ydD8J99MhZOmJjpa6SNs/c4IWsmL/albDQ
2uD9XLZ4K7Gr1N46MSaiMVYZY8UQ2mE2qdy8q4Z6zneic6tOExnlGNTjgsfn
0zzng03lrHCtfD/UNNTdXNeurrpYE7pjirwGIzpNOzDFGQp4UufHHkYnSsrq
LmKJkJDHesew+1doq/zU3c2BmqIFzhH2MbGkeSWcluHUo6bAG6B1Ve0/PIKK
nfBSRaY8mhsjytpWOXJuu7jcgHQTbn39DkT6T4n72b2lsxalAmUeL+3ARHm0
2X9B3+EnojDM7x0UmXjSBwaKxYOHAWRNUxrgLzyaAGvPq/PppYHQaW/Kw+hL
2xHzAefGA4bvLQyr2HWX5hqVDzfeYxanlunEjeMzJyLYzb4nCl0t5kv0btX7
sCc3HcVsVZDsc0a7k5Nmd4cZr0wVQgaFsU89Izt6w9Tg21LofC8QaWa0/3H3
2+5zWKfYcsgS3cptH68oDVUaofWaeBast0ibaIYKlbz8HmJ3Mxdz3ZMeRzOs
lkyC5xxnyahKvyHokHDxdIh/OW+SP0O++2LHvgBUIyHVA50rukZvfr/amEd8
IqutjQRJDn7x+RFX5LCsveAiVy7KS9bGpqI1eZxjpH/ioQkiZ+dtUGhy6zrf
hNwTDud+RysifX6yXJTUCQQiB5SeY80tfeDbsP4Orf3zJsgoyj5WLP4Eoa+U
TsBczLijQUx7DZIP/FTLMtRileiPo8hXgiSqEw4sl9sbXPUxp40DlzRwpUoF
Yl7Z3ZoICgqhMEVGtXlDG6YfygEXU8bg+TLsz9OuMZpzZ0D/5iGDfdfWeMin
RlCguUFm5QDtqKdk4WemME4zuVUznUVaIuUuksGOZQ/poGkbKP/kN4uWxT5t
sF45mIqZMPbAxAQvEbX44HKKieQlGgYfPKDWHLamXYUBBWpJYNsm3nXh+CkZ
VQ189rExZdirxAtvxi4Si0EJp9nF4iuADyg81bSCa/dOdCBESn2pFkLQS1h9
fIqYGqFSixQUen51Rq4fp+nsq8CxLEUIBKBGiw4Q0QSjszxo0HDy6HMGAFMw
cmUKBU7/kkjgTF78WBNSdwiwzJBPiHdnjZTxVjp/4bsiIiQfjgAPddo1m7Bh
piZYPoVS5q3WAJPQjyfFI5v1MQcWku9Pm2tKfJj+7+7QeWHjhTQgJGhlWrSb
yyzCZHfPPspkBs9A3fYswA/w2Hj8JUy+UYY/hfr3g9hqcEBDz/RiTWJVJrhT
wzcz6urXgSqp/KnZ4zlQWhyPuBkqU/nzL1CMw3IkEQpYq/JUYW185tpu2VY0
DnD8ZmsTJEJhqk4kDQ9CLDYdmFDAg/c3dGQp98OaqKYXMeTT+n+yRhZDqduS
WwJm7ma2vuIWpYT3FmGRcKjfoWt6GLviWl5uxGgsFWZZAy5TfPbo/huM6ssX
jrRuHuoJkYJtj4ouraBZhPTqLaa4ujFMBxTbw3RR8f1wYOOzeLCPjaJUfhQ0
nc4ACGs+258IV/PpfV1NRnugeYKv8ojCxGPOJjDZniSzCxBu66hrLzW9M7IN
WedE80ikarXmilk5MHIynv6izmfbmCNAAtidVKddNOOL5JbWqX0Mlig6vQC7
EPnkJD0LgzsxoBZx7lBLyR3P99UivSKoIExpsvRGgLwP7u0tAVRPEggmemfp
bPBU0W/wc1J7KiOF/SA6CH/KoC9wJmwJltIIg0g4O1Wy7gRGTurhK2dh9LL1
UQYNSsHeuo1VfbopB1G3Zc4KgA18GGoCMG0dNgylHTOsRtmhoC+878T82jv3
fZ21MG3pHkIsMU2ttkLuyBbcTzrNOfeZLLdsZQ4COR+B7eFM+MhbTKfrjzmp
cUxd1zH7knEXxfdDDpA82D1q+HT/QlmlxtXJut+xEI4no+MI7sdRp35hvulk
xaD1pOqP0t0LL9Z1q6C0DHGw7fC5BkiD207O5FKzvVFfa6BeQPKLGpgras3e
lmz9UAjwkjI4gHRJJeAi2zhcGwKFdttwMADNlbU0jTy+yb8DHKMQ73SjdcaL
Y2PM/jMTInMPmigKj0js7geB4CqPlRa32eMG1seMo+NRJIIRWq+hSQ4LvAyk
h6CFa+S+83jdMP2zuFFuEvD4IFCYZ6V1e63R5A5lSbS9/mkUExQFFeZMJVIG
1xavWIuo35f9ojFEClnhjqgrKxsikcMIgZtlZLNz/5s2d2DzclBoG7uJaOom
XbbdwVai1BIL0uLrz6GC88JUOzqgH8/I40n1KpgtL/MLTKib2tgazU7RHrm7
7eTzaJeadQrWn4yZcwy9dUfMAL0obphX9NEAl8nLprixrmv29nacVrFmf647
jXFzopxCCW3vfGh7kBO7cW+h+FCvZgPcEOv19ZIoOlrTgZND2cxu8cfTMa47
2gG9idZR136130CybPFSZkrwn/UJqbaGOMZvryZg3gM3Z6LXmRzkTGh24sJG
SAGnJZ1CFIiYo6zb+tHgOMobqXpEpiMcGRjFb6oBb/Us2WwNHDJwCBld+9Ob
G0VMCrm2Tk+O1bZg3AiAhckhLq26jiEtUiHqJUXaF205iGpkpKAQqw9SceaX
ByAZaR4iQLKCp5oRjDtG6SSS9+fyo3Sa2gFX4n6Qx4Fm3AG2O/tOQR3iaY0o
4CMBn8tu/MmjZiawD6XmCJXelBqc2lmFnlxbGXem8cVqzTEUD+Y01/z9BvT/
l6TlRvkBBq3ugmGanr96nis3clKjXchOE/5U1da4YbIoWLkkr7AyZ52XdLv/
v2bqspbwI8fOuZBeRaXPRLO8x1IXyav5TTEK7+L1rfCpUsQ1dFp1XRcustoJ
LBo7vvHsiFVxP3LB66P6+H4VhEezXIwDZpFYJEhDbfHF1o9ed00vYIvg485R
3c8gb2ystq06hEWX9KQYcnaAwHDDmx4u/FyouAH3uq/Co6EtDtErmaCpnzE1
sredFX8a22qTtKf/xf3o7cBjue9O2ZUWDXEN1duHULTsTKr0D0c5DPXpvb60
aMYjaaV011XYyBuvMfyvMOeTYnzV3Xky4kZIDN63la6dp5z0nedwYhuXt+nV
TcjLFHH7CUPBtTi+NVdra5vCCbB5j413/nge2NDbP428fAGjWaZBiKrmBZN1
k6Ng1Sr0nOQzya2+rkt5QDlB08ccZbQhCQjLAWjdb4FD9Ayvd31LFYOyNwCx
El6wlpVNVWa9hPIEQ2J4eK7TO7c+knQYYQBD7IV2KHRy0MIjYUWcC8ZjQcJi
ROb2UW30iEMDAp4H/A8U4lsftgS12q/JADWTAouElghWJv7Cdy/zBoYM9TZa
a+OWp+4gTkio/vTsgKg/XWeh0DxfgvRtYprxBE9lx7Fspzsb1Zn841mtaqLZ
rc913ASz6gPBG7m69XCD2qINgKBXT1YzIOXEb3105V6OEmUYugZYXmAtPDBM
XKxz7RaQRKV303QNEdlTUGZqqP8quEf3mxkMRU6iRaQKWGH9Ns8Cj9YeApLS
ED8g3m5sMlKyC4qO2m/fsllmXCwgJfMCMokh1KejKiqfVkGs5su9L5NGxcgJ
2bclrbcxNnF6m0NxHWgL6c0F6etBe7X6lYHkt/b2FY3htbMDYxSNn2tY/MDg
vp6zjCVMEpyv2mcUk/YNamMlZlV7CNRzWr2QbZnbpMcQkkhsHjMuXrSoEHO5
54dJ+U17fj1PvvHLUozYzMSBR7xfQ/PNkt+f7NjG6f2+WN6OwVQF6n8vqiaT
tNunixhq7bs6MVuENXTsd1JCsseM69LHzHQZ7+BqhMRiHf3n96KC2xlOSdu1
93RCnquCfj3sdTuHmgNhIVigBcnOrGoEO7jQZyGRyNR/BQ4SVfqXdM0P5pTC
8H0B7ZUKE/ARdTLNUUo6mAv4NzWK1KtEhUBdznj6/+ntTHY1go+uvn1yAKMv
WZXBXf++2zNahjObGQto3Ly8Y5+BU+G258OAlPbbsJ1ynGuZPaXUJe5i36xn
9zzJUnkeHtMnGKfPzYPicKpu+0b8cHuJTzdImw9rckIo+gqZe43ESDpNNyPE
aZGslNBM4KJyHZ0V5BFu1CEz6MiqQI6X4iibhPVyIA2/mRv8++fuTwqYYGdN
bnJp+FmybLuAKV39ZNXX7VFaPsIkP5yv++oSbJVD6MAAhPHarWVbMuxw1NqV
ICppcuxgHPTIh0B2uZaY/TbC5veYcQrUDrZq3OTT5JJK5hYzZxdxz2gDyIkj
0NO56oh3dKVZj30bSksSl9HG+hAKjJEJEwVq+ocV1vXfOL12JFaLMGueqwGB
V1tVr385Q1M4uGVpxPIuMrUduVmYkT141VWlFiV9FOqjZf7YNBfXsubAGkAY
a6Lp9EA9xdQKP6xCoyoXZVmmVZDQvqdey/kLGr7FcK/3+EGC+UYFYFJdYTGb
cvCHK5eq5lTpGsR8xMEyuwgVkz9ij2lzWWgATnmFuv5Xg7O/xHLNjS3d0Yfo
wRoCpjNqtqGplqNGdMTs/qyo4T7KoqSN2/FanjkOCMr2sKJMsruvawa2hrIb
jTJPjkawKJsqcj/DyHWDCMox0tCnZz8G3od9kcIKYS0cWsBEaZB4a9p5tL83
hv1DiV1LOUYy3+W7YfGzdCrFHDaanj1d7u1bfaUZXTYwptVo7ATMMQmtfS/P
sOQAYgqHZk6H0MI4XsDmIkd7MccyapkgiqcXjrqdCl0lowrP4F/5mtz+m3Lf
5IpQJnQG2cB9GPVeE92PUN3Px/c5EbHu6rAmuBNMXelaFcXfuyNsUJSjQOus
6Gc2THQlEkyyI5gqB6VgQOVtW289vCMQYrYDZE8ULujaUepBCkfdqTe1nY7K
7vLXp3xYycxgtTrE8xwIg2HabTtVYrcLic8svdP7iJtlycuqtyXm40gqk/JK
iOafmvHSQKpqzJIF+1M1PsARLJyrCTw5lBhEniI3RfAAjMEz4roiREq/FpZl
ohO8uZp+w8D8/6Lc+Y+E6XhxeGfPndTqDrQL1DV7HN1WQLI4ePrff/4jGjyX
T7jXJ5nVHh7Bm2DLo6Rm/7Uu5YZuuDy/bbYleXnjEhlLQCEK4Tkomskocx3O
xwhJ4HH7ZQCnwY8+h95ZmY3w0BoE2NBduIFbyYD2wqk80TaOMKrbNEvuPG0o
yosdR95wriD7S905P7DdKlzXP1nz/ncqARTVuxP7F0Azke8VX7sgpB2/qqo8
tA5Rd602ihzr60Yh9YfQtsZRNn4eLIDGoti4wR48CeG6xSdEHwcW09YUAyJj
NsW2BV8gsHzryQ5uVQA9xOhBzBE+S9WmRiCxYZGj5jpxBcDJfbaHojb43Dyx
1uM/gozJHFVutenOQ8VxR/oaSHEAAKPa4hq94sL0H79FG1RdqcGit8cd5LRj
35SMSfgiwnyRLpIULT9D7GXdgoR6koTqAWqLj2JluHKUEgF60WIURhhCNGC6
IVtalQtazl8lYp+zALGqLJmUi2kGm8ErNyz+WlWDs5FgEVN7BroyOMQEw3k9
R+cPgdzj/cbSj9R77nsKdtQrjThm0NNHAOGcG9zuvKOVxK7jZUPnIxLyfvne
srcxUU1DhSsdTKQu+SaBw7K93+6J0MiodQgB4DNkOQ+ZE0jkpWFGU1653exI
IKh5LsS9rPGH0fWL/Sc819AxTwSN1MOmRUYvUI+jPyFfZAB+KmxX65mDamL8
fBVCjFRtla/6+LfBn2P85zbGNeGqgEMkw84OC0vTjhW6ZH/PI8EmoYihS8Bf
AxpDCuox23S6W9+OtTeEGHuZw09cQ1FFQ/TG4l8nXmRamxYt2Y3FGC5Gdj63
IP+tjvg0M7knSlyFI3Qqevn5aad7/+JvIZTKE1djbtSRP/cTaZa9s/KnV0Pj
+L53NDCiQj1VpXdn9QBsPRq1wlrjrQObINoL1IR4kDY17Wh3aCE7l3RJC84l
Y6+a/0vfjQ4lN24jnVJVUUjBHbf0rrFGqwpkdKpheIqkO07XiiHlq48FZ+Ro
hLfzI5EEHXN6MIGNBEfGAbxstgT6T0GfuBuE+koqBZNEQtPPehFjVbPQXyAM
JDmRqPeD0BrFaIHAiICvpcDJ0AJlK6HxjjdojcBmqUSUhEFx1eFRuWEXu7DQ
MOQlbnrhrLCdqkN+7VSlrvcbSk6I7J6vJi1YTzOeTrdliiu+Zbw0Ez59sgUe
xbVXQ12zRsx6gPIZQJva5JctK30CVNbDMD2LVom/paZmGmghsZSiNcQkJwRM
qJlqe09sFURV0WwQQwaKgeOfMCqLsCvLShfmttdYYbaY9Wb12irJWpZG07SY
CnNnl/aQ0G4E+YKcwqYf80YLr/JhPhuk2neVTAS8zinEsWDmI3591u2vZRuW
T5lqx9v9migCpEBepBL7quXnViRwR4O4eK44g3x8tHwPFiwJDZmzz68MmrfP
9jmlGzyGY4y+J4/C6dHfDwZNrYAkDyP+T5BYHJ0IZfSTLfVIizTxWYgrFjLq
9L/Zg4R2ddpWDAEAfVOp6mkjKqRnCaX8yH3KpeNo5itOE44ZogoP2n6R7l+y
L+vI2az7JcJ7PpcSZPQinfw+ccwIRwXFBerDlin4RyBMitwZALgK7YlaHIoC
ST66CyAtf8O4tWURhZml/TBpyqcKjER+nFg6/ObFtJKvTD3JleWZaNkjY2wY
+U6PlcVFrj54iKrEFLGiErdvYfyTRJhPdnVwqtOOoDAPpV70qXbihySeco1G
92CXZNpBsixpJa+eN0qXVHUDBmCBC3nNriS0YxVGemvPTMSjYpqbcsjUda44
nmvxrxAiWnWdRPrlEAD9wVoP229I5ojDwxNvOCsHfFhsfccbOW/Et+3cF1QZ
s/YiusNTZSWOud2g+sus6tcgcExQeaDpN0UERP4TA+Ru5cc7koLk9pYthjF0
oIApAwfxUr82Iemo4hTy/sJVUSF6zCfFgPoW+uU9lwf+5bUmTsH92j/3Fgbo
xWoGiKPaugsCfiMvRHK9BsU3YhkMR3AXaZDY8k+gIRDly/opKmfUyVru9UTN
GZEDrqNaVvgZ226rkuQIXzdc3gU8Lrjk9DhOsZCIqkwCdFKMu1gPhpQkCS1/
C7hWAJYK96H2Xl+kpOWRI47hpcCPWC1aY71WDxj0EadOY6jeyZakjIkcWKUB
HD8h5XtyMKaU6KohmnThud1ZKzrcEDumyuFzFlt3I1oi6/cqZOSdc7qa7TDG
hAJXqfUdF2XXtrP8+gtxGPfHp+lnNW0HVFkF/yGZ8wf9beqtp5/G0PdsFh39
AB6j/s2Qf04GyoRb0YYxLynwP5NzzPyjixTfiJdVeXwKdfLY+IKHlfYhbht9
ZrYG8csqH7FP1lTbaWpDfXAgs36izKAddSiihs7p0oKsszZqjV/c627snzs+
VX91kSCZX/hFx/4e/aJQrgHzKVeysopTGjAeQHpe6xSMItP5edUWCvoiJ/Ps
POEdwGb7iqy3t6ZVXC5Vb1CA01DO9aXTXiQPghyXx/3rzgpxK1aM1seyQvTN
B5k712f6rkoaS+yEviu7dr0JtoM2fkBDEXeiWRbGGWxwx6+mRMspebRpqyG6
k9Zyg8aUDuYjC1J0zwn4ZCUtY8+dWX43hqPCv2e5rWHUdsyvlwCbk1jL+Pl2
SYrRQ8snudWG8T2TPjbqExVRHpZkMenJQhi+8bqRXhQNcYq/+WIeUeEmc8m1
AYsQ8ej+vtAqWk/fqHsqG8E5ZYwRmFBZYAeOpKlgCPMJqXJT//Nmbe7f4iaN
Xft/emKMZyQM8SGao9LStCvjVbcZd4oTw1p197tAK8PQeh51KkiLyuLk1vNm
3g9dTeWGohwTat+/GbotV0k0nGhxNc0z4dVXmptGv9kmDJ9yuZVDIQOvlEuN
Km0vhTknRL+tmHdoJIOqP+OfGc/gYE7xDrdlnKm0g2EDSW+bRu5sVBmgtBmY
je+hXqc3W6YvQ28QNVRUWPUnKOsqEevKtC3nV74otJyKtHNVHuyp45OhxewC
DVx1DB615AdhCz3O2LvxigF4omIphiqFPSTjdvuoQp02MBCA9t8dIzT8268l
lbKX/ugRTYjgEHVpC5LRxbWRMeH4Z0UYMX+ZkMq+TCtTkyzG1/vP8QGDjJkU
P06ce5GZPBh93X1Ai2C45yFm60vbCVZMIo9pofW1r2AN+NwFvI+I8y9CITrQ
k5u/Jp7M7EIQQNxktvp1+4TXudaCt6X90yqMNnQ5m0awPRpCknXPRNDeKSF1
09UjyQ8eEWqAwfL9/mrcrMOYotIGMbylQ8UMnhKjEL7A9C/gPSh1jvPpPPt9
3QUZejmxuD42tJboMLz82YdHG457uxT4e55DXsPWEY5j+R3quwYCTOMvhWTU
hQdGuR9q2Fg9Yet1VuSI98xaQkY8CUTZTgOdsnVRk7iSiUebjQ4/OzuBwf7H
aimjJ/yf2qTc5olv9Hjb1f0iR6uPHSaWpFtPLWs+qX+8CIsB/o0i62qo4Tgw
MP6rDFcU3sTW5vJzd/52w8Cmx85yn1QCDtLdaRWjjLwykcWD+UZcFfLAuP7A
Mo0jhHwBGoYOhWsyCNCHP3kAyCvcysTRS0tgHb1/9AvQFeQeA/hhY0yhnmDg
Tkasv4Z7dEqB5CeyB5gTLCUDLmFzGRSb4y1sHDzqaFdImqehL9UXV+EsNDra
ADhutfQLCNmDzn48omSa+fdr426ssQudOSC4+oA1QIDfbAIoi+jCavzjaY2x
2oxRkbjFRbfWEHMgRdZ9BqIF9Te1/IkUJ4x8neYzCC0Wxj0DEFRcLz5Qn7i6
KAKJ38hmo1v/JVofDbrq7jv7HCfLU1fUMJoQyoxlD8ZSXmCRRuf+/baNKl7g
Lk8iFslWDq1Wpgj7JZ35R8meXakaGZsHZEpZlEA27/kzOygvo+OfMCLnayT0
ANyKxpdqTsU4qB4pT0GZ/Utjer/JjjhY5ha98ebNEJsuvv0kMcFP7XSNsO7+
udEGBKbFQ3/DYJs4crAePIWzJJaH+wW1P3s6dfC7gD1w2zIH5cpAOU2JMrPo
7lIVVG3WZPXAdt+ep0bCg2OzvNRL4muReSQ84QS3U40TPTMFh7Mlo0475MYU
NKyCx7PRejGLBOz9wcBkRRm1a2vFuvAu4nXY7UJli1Azzv5OPH+EEFTgmp5I
L6SRRKWQLlbIaZs+jHnAERJLh7GzuOYH554tIVB02kLcQ7S3xDXznCgfZquw
c+Q/2sYGb4TGEkP1EXcz2McnNRmfKyZhjwDWwUiY15iQS2s90Yka1HvKfrEn
3s59dZ8D1ycwIXnzCuYChqQpyyzwobbHShn20nT7yWCkmdGy1vpBhTDwJQyr
Q42x9HYQyiV4FF2XdljECLP/5E2bNeYzBaEqp/9CJH6lcEm50f2CMGCwIc+r
Llbhprs2ESscOeAo9fyuZa2Q01994BTa6RJaS0tmhLmswPnhYhter9/sC3C8
htOnWJsITXYH/nscSCmuoZFWmfIPlbUpVMtPgwp7qgDZyQMwDmfzmoN/+f+x
QqelLC1/u9SAVcE4yUyyJneypS4LY4hUYPXErhVTqLjPBQdaLy5bKKxW3oFW
HrzMhExSKNGE17bV6llapptDFwElFE+gdFBH5d8Q8nnyuKS/JGXjkLobx7Un
NoEgwRAHTDQUePFOz+3j1a7d3/1+EirNxCZ9LSw2ZYtz8aWmI8uvlh0j9iQz
tpjQIFnmx3vVaP7qivUUKjCayfK00byPxEwQM5DlvXj6UxBcmUdq+6iC0Kfk
Smo1W654u3peXFtgrKCZsqepTK623Xw0zBQVf49DWgxIQ1govBUuOypaLszg
6DYGFsb+8CfDctZb030c6lUxzQ41vezKgk9gnMEYC8hbvgjreRjWNOytLYzC
MQ2KPuo7NfZScT8Cq79WW+VPzZOFYLLFytyEYtADo1SrpoOQL3qQ6oxTLkTb
97SxOdnnBMprNmxYWPdy0nKu/KaNdecjrntUstWstuH6EuL1eljVXVcNrSjK
vUkDD99vuSYLg3e8rntsJy4v3d9ZG5yuhgDPw0nzyVCvZI6zIq6x9n+kQ+3U
Xw2MPxwHc/1re0VeWwkXK0YHBOHivBlmZ9mzYs/8LoNwiRwDR3vMUslYSddV
10G2+w/syzRbcYpV9+lexyJnm7HUEMW8CwfVdFcvGjSF80GxFqsdc/rLf6OX
ByQdUjbGxO/AqbNXI16sfi2uzfc67pzTZMty2mnYQvbbtlTW7PLecRDuEENd
dge9+dFxhPbCWyOzimMiuoQHGRmbULX6hBe+uLYucUGYQH6V9ROaw+gVRvjf
zV8E1moAKob15muzHcIWLAAdQsmlCKZoTcF2SeczNnqj2ysLqqOsURuS/Jla
GAwYHx46iBb0aJXI3tjC31SpZhrGDK1R4kRt5E5S3x29+uFWoxbXcTEUbevk
WfPrSHM+61o2PFTDveoN8zw4JdzWLdfUAKHTdMUTNyRfPO34Y8Nic+vh0eUq
8LFUyBVS3RtPBe1Pj5t3lohlK1Ruc1ZVUIjYHxQkzVULJQ3D4gUWBkeFzSXN
wYSpE1tQMUzRJ3ZOfkcOK7CIV0Vz6MsVTbm9LAAfFjzJLhpmWqztFKYZpvMg
xLouc3R6AxqB2XKoaeU7o2x2ZNIJjGVMFhOfFVNqqRLEYwLec0VIDpdY7R5q
h2XXIbM4JVxNUNKZ2iHJKFRJqLgl3g/jxWIFq6KEGtApmHpj0FqQz3fW6h6O
Osy3xHdWXfKdAYoSYPhwlDZeQ3YLbAMDi7cBE5SVAk/akaYVX/+ZyGdEt9gm
/JKiSSNd39S2hLkFSilXJtfKtSSEmTfJPc7AJgbwgFMC8OglgiEulYZKYdRy
v+oN6XPpQ6DNHDWxY6sJzaJo5P5x0k5XtV7qfq92oFLBdBaGSdtYUYmhu+ie
6lxcQ7h1bzu/gpeAjER7Jt6cN9uyE3mKUr1lMig+gyKqdiLvqcOENOZ13h5f
MonP9XQAOmELP3ONjaLi0ICtCYWxftILItLxse8KFvzrQ4Y9QkgkvSG7HZaM
tkgnb/M2kfor24D7YtKNyuHqQ0yAftnGyp9+lYGLDFnX0zmNFy8wAUHIbzWY
F+XXx0F4zHSc3y8EMDDKJE/qdaMpDIl10j03C14BapGcZpKGswfYgifRdV0b
UGboMHGG//Vrrec86ogJAw0ocl30nd45GJ8CBuWAJ2I/SUDJjHtocao86eNV
RYmvhA8Hb6dDNdgMVep1/DlK3wqRv4cTs6ju6yI5/BdaCL84zWANYxB4VD8K
aGt3vWTmrL180IF9cR6j4YOC8MMMuTmR9ePjd3NZXK2jMrU73l8y6fpfMkd4
pSrhut6i64iXydxdLaY/wE+yE0FYs78XMwEdUrGxRcV0z677xzNUtqVo0lrt
PJ86iaytZEK0W4GJLJ0FGMyXnrXDCQJqfoSvviiIqyUGdcbhXLvjF+7D9uhA
siXRGgZU95UxHyiy3VFz+eMdaBQLX8VVH6prTZoWcLrcZR+Q5zo+UKuFviLf
peAwbeZfMYi2W7kt7Hfp7Y4juQgbvjmRAqydUg2qvaMoAfB1ZbSSHmOxErnk
ABREFLnVYVFSmK8JoUBpSCZ1BWyGjToosYw/I1Dn6n0wA6QYp0rLY8KAB1IN
utMYoE+EhgY9f7eWjVpgz2U5wdzt/Q9PYXVO+ObFoeoDNJ7+k31n1sR4jEZt
mgCz1hBRbnameRovCsfbljTJ9Ym0OR/G28UdHyOS3085Ed8s/rhmLOi9LFlX
BZtG3NHtBf5jiM6H7o2uL3ekmLPvAOc+BwMflU15AFz9hxHXbhlM5BKzBEG/
3VYipOiw54qYOzxQ1CVptMgpXi6E53TBG1lXZ2iupPHvjg+R536QNtW+Rcgi
fKUliCqcuCKifPtYNA/UD9pts+ZVhMOE5DXqEcJW+SRc5IFa56peT3IeY1kk
dUPc29+0m1LgTEMPvMFUzMnSnaG2US+YqeFr2kdMA8gKub85nrEH9nWPw0rM
1j5KRPEKGkyOvP5TjB2ONlWUztB8TvwURZk4h3GcqQcXk/a6PkpC6nSoIT7a
3fc2A9xN5dpAPz427GXeFXWLvMaNAnK4avD9K3XS2AFK2ne83A9i9Ioijoq5
AgvdFE6+8q/xY31WmMdP9renUDH1x7HC4KmqqZq0JmOv8cA/9iTq7QcBparR
Au4L4u6Pb8IPA8TmPKgT3OIZ7qIW+fY2f3N5HmSbkqaNJBW6sN9+dgojgO3u
ReNo6/xBDO5mR8BqmYhVDtHKVibsP7488+uxkSOUcVRYci5LwjmvVr77PrZw
CHC+GbWOFeSDI0JGNoTEmnfqd0rLUghDOqp0176X5+cjrO5je8O80fm8fA5i
Szn13WZvpV9gIwoeZXTVHf4L6BAWUSYTSXbOUgp7igFrULXZSX8wyCYiDs5t
RD09nvEFVIRTrY6g/3egWqKMsssf4CFPYUu2lu/bfBmaJU97HB6G52m0LqGs
GX5pEphvwvGHsqaIAlxIQ34LyoPMw4F9pr0d0PtKjJkcCzJl9xcJsgTgRQyv
fOiXeabfhF2f1fY7Et9HI7laHIRB/TfmqdJM6ld84k/aFb0CRu0Y0FR+lxMk
oYw0lGUivKPs5MC4MphwCrgplCS+ZyqmG2P9hlB6Hw1S+zalOjUKcEW6sxyO
OqzZHgfepDzH1q3GUKkoQjhjfpFpgxtVUi82u5ZrlioaffS4/omK+4ij1ycs
XpwO9oKA2ko4PeTPxk2PERD+adU/xmOtkBdJdfCTw7GfOgy5mZiMMmJN+YnL
Jrx0j87wbQj2ADXlMx4gkknHwZlEqTslAdDJS4gFh72FyptT1BvnojAn/cjR
W48VcVNzB9kYz1Wuo05pceJ6Eq5WVKsRgc70DbS8ewLdFR/uPQhlMoos/CNN
hXvvs/DfLfGZS7nVZGbyr3RjaTR/rj2ctS667Zx7ouLPGeA1TZ3x0WM+aWdV
yE8IkS/2kYhimli9umVetHuURw50ZXel3w635d+6E/Kk6aof1PDJzUsISq8a
BL71Klz6CcoJFp0S995HEA7A2WESeEBfrMq/qevgrd9XNaqKlG/+dNYWb5n2
OcKeOHH1FJ5GOnEVpmD9JRyf9dgK8bJv7naBN2xO7xmj0p349VjuxF2jXa/u
hV7LtXlD2rhIUui/k1JBCwypaXdmdzjcKvRVA+MlCRfNg13afDMfrPDOZlJ7
FrLHFd+/aomB9PD3bt57bApfoohBClekRuCYeIjJuetTH6Eeut97t/JLT1Oj
28PEN+nE0Y2RXfFSSUOsKNilulUvmNz2JEwHtgK+oWT5yCcwVOEMJ2/Tg3PJ
cjDSVwGvaliFhVe2m8fRXkT3sy18sCS0mY2119L3+pXkFbmHL5a7euUniaxa
HvJbQsoeM+ZChA02ZurCrYO51kwDyPnCa9vtT4oKm8eT0dJuB2uz0D90IcYU
PQ2MRm4ekxUqyfgl1g19zO+Y7HtV2AxKxrl7axSpcU+ITsTtc/T+oV6G4dwC
vjBWPGNKY2HyXXpMrpgEbEmc9SwshiUSHEeoR3hRtSX6dEMuuqlAQMXzKTEn
f/2rCb99WcqpiuYDBi6GU62c0AMrV83kOSNm9XBwsycz8TYA/pLFHN5/Cd9g
YPKvBZx8OBUN663EEEOqFDplxU9tMVifkZw1PtLd2L3g7cemOF4sqi8P7UT3
PFd9LZKOvHenh7ho80MtLS0O3aJnWhj2T0Tj9uogINo77z0ciEZEHtOUA1pE
cdamvk4V1e0awJCQI29qW2AQOPVI/0ilxAeyAuyMHnHr4FDM1F3Fvs1F7Odr
uWmkXjeQb4bSczhE1TcZxyC7FPSUoLRWfviXLQ0t9p280ukFtfMafDSWVTgJ
9R8iHff22EraQypfDxF8LiVfsVhsyFE1GgJPfoXlL8TKTsqfzEMotTGan4YW
83/FiFWoJolqTRN5aQHpFQR5OzHBuQUidcSrz88CviiqbM++lis+lcrDfHnm
ahAfVPC2MCYaktGydZxvrpiry50LWUjbsKW7z8XMvHUwF+6UJ1KrYYpVzYLW
GQ9q5XAwgajREBbk3322jSlO2SruVFsQWLqZOQe4PzW7lS6MmIo53RO+7zCw
wGuQCbBAT5LO0wVR5Dgrg+22JrdZvKuVhOYCVbEjQAg9LPt7yB+fELgBXrCr
yqjyjaHbE//XdHDjQeK5CswhPr4va6SFTb4Thq7pRtWm/uHBMGqzB24UmkJE
4vyaS85O1Osxl+i10KG85snYxg06nkIH08/LJQsPJmdgm2VzW0oE5Zkn9XiS
GFBW34M/W+Wz9FjuUXPF5KXpBiSxxvSY/ytB15S7qtOPOeqWviQfE2a0rFGB
HoXSUJ1q2t16wEFK2yNtYobJWICkSGJgtXzlkxVU3gW3u0fbASsr+sFt7/Bg
P1HyS6Y6a22Q+KJgE3UE3NUsh6l6oyNk2wydWfexeg5qe8KTda1haj8E73n2
oTwOWqMuYWJDQ+Eo9Sk7bsO984iFx6XR4p54mI7ehp6hrA3cCeB9n2EjptBE
RxyHkyaZvJO0FO19AtUowhYUlgO/co6GhKLCrJTbh96GNsStRaR0XnuvVBLW
XMbFAtaf8Q35LWZ4RzNKjp/3w2AvYCnSk+4lMzvWMQLPlsHpkJDaTCysKO5q
Usr13rzxEV+UOyd9UdLvUFhBAhOGxgnP9lRYhgtnkjsmfubDDmTyLE0I3WaZ
QeGe6xKdH0z3ZhXTZcU3nACbvK8j51bqVyWNTt5mAiIx8FeBKYqPooyjwAwa
J50IyLRwyxYa5v/oXJ5miiIFYN0cgz3kJsQ/qcf82AMYKQomXfbOpkTKJrv8
nj/GOi+4Z+PEI/ys7+SXXcb4i+m5kvwEDIiiO19yQzZ5Vr3+MjwPGqNyMuTt
SU/HXkKC5/n8IPFKeSMqY36bQu1Rqe3Ue0CvyiXvXTYz32RBDjMgeEjUBJtt
pmxZsSS4gx8nC9KPUh++U0AMmTRyd2/OzdEvxIORB3r6FWK0X9Xe0gXpOz+V
uMw2LkvM2SLJkfn4t8ZehiCLv0iRrFA5F/Cu6vznoLMtXW8LyBbNbnz7YwMs
Ci4liH5bF+/2t31F/M30kZ5f5j6Dp4deRxiP5oKS2jEkNvgNZTfopwsvpIKt
bdVSEJBluZgdv/rhFt9SVoiMnt0SP5FEA8y6ugeC8g6KmOc8oMRCZwGudc/k
HRdUGty3QBrBTulUE2zO4twxW3BZ5oQYFhIrrqnPnVskQkA4ERyCwMSyEz2d
cKiwtiMw79iEwp63xRpgQvKSMaiw8PhbKq77tJgq9m1E1PCyfnMjtLHKrkZ4
qTQlozhQrkzNhDSNPOtxSwA9na7GAQKLBX9pLl0jRAi4GsX/A0cRqThpfbpF
yVAHVnCswUdL/NcpoRceAWReBGJ/BoVTzvtouUkYkfs7P0Jmws0ClLUQrS/p
TbKwj84EaotlSlkpwIk2TlowdOOXN8iblDt4f9xZR1AACW8G36R0x7Tdxs1p
eD6He65hchi53osDHAOu8H826FWNonF4Aqax6cv7xCW9L3F4I1xLmCattcnh
4njNjAS1nfUKkS77/g3LN0PWR7ljQ0h0kQnngeyAiKxJSJRAKg1YTihADKb9
RZckxukz8nwyglkJGWctaH/PlYtXVOEKKiERX3DOumk3Zt4BIjnreTDRkOwM
rrLD+Dw6lV4O4hEmBEzjOgM80v52n0OGY6kYD1OuFNs6zrJNjrZnJd/GIxyS
wpyU32SCfTrAdw1NiyUefnf3dWXL+9zLk08S80jzXU3t+hAD56Uazlic7Lxj
dmuBWvV5pxRfpQUDHrpoZmpD415OsvTh4/AqePs4Azxc/AQxDBDMoWhd1dzI
eTLrLiPiCirjdMovizMpsh9g76yhMh5udJ93aXDouoNhJdlawHIqFUyxkp+r
jVCG2v75i4jc+oLb9zhcb0kti4jQwuXWgFo8mnuZu+Wh6WkSAT0ikmsEFC/O
4ZXMkmi8pvGesBKe+sNOrk+pA8DFpyouwWbwnCZnos1kil5ndLul8H5E3hg3
BdJtUhuguavxdBSHoeX4Tw6Qm+1GfqHW8UTnyDbZSUS7imJq3k2DxtAB4XrM
jYn0n6Ld3fPaiRQMroPNAhYVgEKCXm6j/c8G92G6H4+oNhxMf70Zs4egnEo+
yCwyz0DFq58mtcp8QeBiiFaNWe/VRyaEdOm7OkWi5WNcwe9QTuRZc00LPvga
Cb0ZiIx5usl2lX4rmMoA1D0bXl57VSbX3LfqnmVQYwb1Up/HXvkO028Lydi+
j9fFRbp9uQjXhD43ucU+18C1yEmFssOvvwazsQJLKU1D9EgNWMOxeXEa6Q/P
sHAuSRMbCkjIFERmei/dyLbhBEsIA6MYOfx4DtjPSEyTzfGg9GOvdv0Kikad
PzEs2y0+PRk+ff3O80SvaxXtXNV+aJWHeX7MQmSBbFdruPMYtnCqE3Ee6k4i
dgvFI0mtNkp5FmJsBHkjjkdnEoVDCI8Kx+9iwcUj4r5gOjrHW0gyh8Cu2vEc
ekZBIiJmTPPNnvJAWAQgVjCaXm8IPfWu5nQIj6VF76A4Z1sfofAi5FfMSJxm
vIu6oJ410XrVu/nhNVK0EWTZX+378NOmrcp7Lhw10BIjU3ue7SvGV5eaGWX2
4CLFosCC/ZCas3fCaRlaoAIRZO7Z6NlBP/zbQofwbBQYdEoX6L1WnVep3dBY
erqBJPTpyW5eBWokECYsEFvv7oLmUvCv/tuevunF5FYtxEPXTTSqMrf5/OIj
n350G90nQCaiNX2R3UD38vbYWRjvgauHbcqP15NARI/2wbbBlgeGjDIM5zKW
1o54+brk6QD59fqpiwtwmdiRyqjpy9/bcWq3/vEuU6gnBsZvSSmvzOeDMUtx
OzCHDz5u0EgAhBD8JKNcASCh5J+hwv7nGpavZrREZBNW2hzN8CuTruR1HChz
4wJgR46r7RbWa9CuF/qcXoodO4l/QNGTLYq0yIdQ6CsLPEL2Zhd2+xEJ6iTa
3yoQtBlysQZGfc/DT5wz4NssXUTJDIPsrHMwFCrpUfqpCHCKZMmFPMFyh2Gs
mY5l8wsB7c6LG8rbBblcZn+ySz5KkHWoIQb6wptGwEQWESNuYK5fJQMDNuuC
Uj2e0YEUM4WkD7vRt8wgsROpFfCEzGK+cbsVDfffEViEhtShbLwzspWOK3mn
t+LclsY7x7g4xMhdMAT4vLmAzmO5Bep2M9mIxadya1x8yCi5S72BxS1SHpV+
PwplbA6Sr8v2hMX2vJrRsludw2vl6y7WLarrPYPd2HaHMZQAAF3+/qWS4E5x
4KnjLtsV+LPhAfZLmjELeDcbMyHFjD3SOuwUJMwaQ01B3FPNyiLjfwIGJZGv
pYsf+gR2TI09Nr9O1VHztYyjQS7rEq5JerAtDldvSK2sGFrAXNGFiKH+XaW5
3Y53vumxUKXVhv71mH3Hw3VzzKnEjLcIuGjSR4KtavkToCzOiomaVM1CMCM4
uiy+rnlKGvOdWl6qrGBcUYVor1CDrde1+fylE2FY3epsEPD+zChBLfj8iOzh
XyWRloyMERexFIs0DK/+yxuagpfdIcVwI9cZ0BRnzcRXhlKR96OGEDUhTSUz
03V5T8Co6q6SYrDN0gUUMJOx2pM1vmsq5IqTlWbtYBwrXbCAE2vK9F2pQ5KO
qeWx0FZiiJZlulUV0fNrt5MdCwUnYa80y5EGlvvKgAQepLvDgeJNue9/Nbmc
JudnMlw/ZvhUUCzcRJCCp9SUfzQK8XRGfkx4/+vS3saLAfZS5EHoY1zuwTwR
NeHczNX28NN7ISNbVfr2mXR0qEJEUfpZQT31PBEoBoIITr5tYr4OfNKdDstP
7wT4IKZqkUvbvpdrn/u/Xc6IF59nnIxtxdP2K/7d+BDQQVc5PGYdyiDR5Cdb
39jQ4NN17SbGfDfiJt9bARaBk1/6NukBUX4+9oExyC1Ysa67RuKTfEtKRKE8
ghte+2avFyYbI501zh0DGVX5d8my8251dhmEhGecDfX+F3AVXiIl+KubQLwF
+4OUkiqEHkTfIHnJ8bcvaQsSRBylHeLGRhTn9BUB2BLlMGapzNHRQnyyQzot
n3I/Z1J27l2ojzzPKt6sPkfc++TRm67yKF/+oypxvTuq6TE53deaFHhmAoGG
ODrGkomQ78TjxzyIXOBfQR+2+kR/HdgimGd4KBFjw889NB83zgd9kTjSuQSs
OrvsCn35GUc1buRl+I+sxablCJtp1COnqD7viQ6HZpj55uLCc9fV/gelDIah
N+8stXXoVswriX9oZceZeFucF7OUOM5Od5n1nw3km/iBjWYqoI9kao5kfZ8Y
k6HZ/708Ke2YmnQSUo5ddbB/3/Jl2SuP3XCHXUefdCqRV7r8qPvuJ39U1TUX
zpK/BG34muY5wJ9XK46RvpSqu1Fwc0nfelFNtiJLc8zGwurDvNBj6r/93EaA
1KjOFf5EerWGZHQQMvYwRm78JjiiH+yoSIGvZEZBuc6M+ZRNksEqX7DuOVa7
oXJovqj9k4d2N5GiI2eBr+T2UH4HbsoNN1G+CbMJzOFVa5N/QJdI3nmudwZn
BxPnQqcAckJs3oSaMHQXnxTzslMF/Pw1F/i8vh9uxnQFQTYGLUSo6xoM0QqQ
s7dOW/aYhOib6GLPVYUEhgII6c9Gx9j7i1D8UMXv46UIfc+Nv7jf0isLtTPr
ZXOxu17rJyTeasdUCVRT7eoQgCHW1STaofSpvgFZExu7T8kvdj/vHck8Ps9l
ZZHSFwCvuQ6dxnkLFjjiHAJwx2OEe+V5gsnBX32oDRYr2Zk6BTmCWvreART7
MJD6b1XLQ3lNxUt6cKzHsdoM1NnWKjLJKc2eOKuz0JmWlOke7oZN+g9KMiCY
8FUFl+LzxIXwJ1QWsfDs4OCNiEgrQeMCud1IOfz6m3r4Zq3G7Fpy89Uc3eX8
KFPe2MZmwLwVEOhkeIbcW37rcb/mllPNTJ1rG08pUMDi3T9GEJPWlJgV1pYX
Uz1v285tCBFru6GT2LiyI3G6yc6VdNVBsvnidiTelBHzBVR1PDk93zs4h5PQ
1SStEF8XAZfE1/Bz7ThVKj64bE9pvmFm90jVTZHAF1b2DLG+QivzzasDLdXZ
96U7t9wmQXkKdkxLTSFPLdc/6W8p4hHVF9vRi/dNlq3NR0ImSfz86dz4h3TX
jBqbVOWXBMk70waLY84ltFBipXDPUTr2S1tSlMM+ICeWxnZLIJRUz4YdCEON
j9D8mBKlZ9P+gLrxNfWn7vwrhQmD1cfkA+DvH1XgiF/A2S9hy28rd6xT4l4/
dzb5YnesRuK3F7cBkeMf/+I0wTkWlz/Hfsm1qgn3QRbGzgfkXncQaS6tedgV
5vXg85cDRwfMcpfApFV1SHHOuCo3lXN3TAqAzvMPX8mfVioiZM3QV7bMFLSB
YHAvLPGTYXnzEIosr9N6XOkI0cXIeJAPh5WOjQQvMsfwXvjSOU0O3JHbWtlM
H3Dj7jIgirHyShPeiipMHVgms8MmJgmnxXBxF9SdN2YRFtGr7MzS94jlwlwJ
dy4Twf5kuLQgDagAg2G+Ydfwp5owVwnMwQzOpqarVp1TlBNdD9lTidHs6pJg
z5gochUUgg+cY1Mjku45B3sDsFf7BSIvUlXMyapPB4+3/PhZDaLgElH9MoYQ
ukEcV+v6H/cAzwO9TFX7NZi9Am7ysnjsHxxteLNoPMaNAEQvpmV/h8vZajIC
HATQI5WQu4T+Bfw09P6aejsDSNRiwpXYMlx6VOZG2PSI7hBJBi8H7RDZZlqo
8lho1eXg/IIj0jpZ4dmt/gttgOgEc97pwrerKzXej7HHEjmGDFKhC5QNVibs
1G2srkwBFIxUxzxNTZt0U7990Z7i/f/bZoEz4PFrTizvldo1T2M6y7o6dHcZ
bLVm7G+GbVTxDrYLRkNtExor2rewLvoOSyJdjL+AFGXeFKAWJsZxfBkybqfY
f/tf2K/dBEUu1a+zdpmY9I02S+6vhJncczPV4gylELebi09muFtgZCkfw9oO
PkgCGuFLruhvCYED2+KBJhiEnzxpYyf3Zp24BIaqSfbM95JURCwflhQIt5pU
2d6V9pqNOhIu62+MTT7Ez5RpizS3x6NSLQ45MtzWxqSrzH9SczPCN+xG2Bl1
pFlYzTiGQnQ/ROcWEvldha4Y/7IHrxxuieomOhoo5axA44FsHfLeT2BbKU8s
3/zL6d5FxjdbiF24ZlP02utCCZA+QWY5ciip1oTW6314tYddrKil0cnkmxOz
8S2m6jtzx5yn/Z9QfpubldLd7n6WSyPrGOSvupgzt98Fk7VCGc3dZ17laaUb
xDMDc8MPcSCiLPuTDymOFYlDwD9ISKt6yrXOKs55RPvtt1hF0d1KY/PjNSnI
5yGLQW5oIBr9XNZJp+xfMCEI8No1mLFAfrylMwyMmuS3AnHVSEV7WN/RAVen
AaF5y+ENWzuyGHFrwpWuTj59RHbPYpDRW8ZGaAc0T/yB5+oDng3F/7k8LTja
cJDL0O0iGYPBJZoLDBSl1nKBmryFIJHt2rYJwEbW0iBmDxmwsI7DePWJ0shB
sovIZo9nQ9NprVyrcLGtAmRzWMFige+R9RTn5JG9TOhMfWC+QV8S3CfWiWoN
XIZZyeiJbzvD+c2AzNlmf07Zxhk3ex+c7oaqshX4OQ2Z2p6gKPk5QlfcwZKh
8NU9XryQfsT5Cmy0gy5Q/wLX1gHxjecyHTHmJeJ++YnXbxKowzYMXRaELzhi
dOX5hi+ukYg+X3kw2OgyVee5NYpnx4xkSgzeCA1XdW8q0/Wv/zbnjQLc313K
oiXYSR3xDY/F9jI8nbOe2cXzW5EoPw2Kq+sRtomwvJn9oMNtEfHVZyvxwd6O
LAE0YdnAKuFtAAOF3vyw86uZNYKTBSqUH/AmRqUxHlZ3DdOwcFG5Tnki8E5a
jRDvKnb2a9sI+F/MBG0azYtt4rNoSYXirUb6O7KCdk3gus+ZVQ7CuN7APkXz
+3pFp1fJpkvxNYaWAldYSrmH8bV4wbHwlMUHN21wpuDBoUy4LGJin5phuNqN
yAiLvsj9yQwsFEvdQkYkMHZSShcYD8HGb2f0WqX2xiyoNAnYyoXITTkGtMTP
XGuiUW+rAor5iCvqdtyn+YzLmCYSApr5P8tyCbgXlS0+l5pa7O0pFT2TwqXV
VxT0/Bye/qvzXsqUJb0hvK3qenqCBPawXi/Ln23YIAmcyVXkbXBxFg4GnX2s
VB8788Pdj/CF1TRg5fYCyIlgPjGuO908jtcTIogmbuhnu/dXW8IuSfEJxEBI
vRUXOBM3mWYlLiVF2Lu0EytNxjE8yjVHKsDBrZ3FyUaUTjK87Bto9sHHZesX
PF7tdNRxrM/P1GjA1xkGYFvrXA78htVNTbzOYXF2waJ3wPxBQKg9j9ttevpX
OIPZl1AKKrt2m6d27zlqQSNLseiKIabZRqSIcjillSo+R+RnkCgpyVyqXe1J
cWQUzkND/mrvp0RepRUVSsVGvz/msRp9OvHucwU11JLVtN+KeIFcLm4dH05J
Ky6FQopjVopg/gRkFlIHd1wRwx008SgYwrbb2/TjrD9vU2Uc4CAf0iXQ2hPX
DsPlPKEBxfBMH+sOTNEIh8oB1kD1Dd3FgMb8MBZKgZaNlaYKgcjhMpdWtPbf
OUDfap258njy1EehPEjScZ+y/G4i0ZEK5OeTmi4MU4FRzmts07wNRe7tZClK
NuIN+AkB3rNmJQo58T5KW1afEdUPWmwZOXl7oKDW+hD8IfcTxoCXfZXOi9XN
gBQ3T91MpGjb3uYWtn9Mgbw09GFs/Zffvfvk2bB0dRM5FHsNTrM0nlzNdqCz
d9dvCQ8e21V63vVTAigSm0zi6ylZp8XgPqdoKHbwKIfDjzALYWEuUsU3b/MD
LRSNK4xtfIvuzx2yx68VVidzjTCsNGlFTZ1flhUaP7aQqJjtQ82LnGvWkV5N
ct8wkRc7dQJq8ixBzroxgzpK+fkv0J8a3sCy6/TNHpCp3pecta2v6E960+lJ
qLhXQkRgvlyALmLTgdLKkQ27tfHpkkd2wwOEi5/s/j1q5CbmyhodniQloiBH
iBxUZGYFEp2YXG9N8GsGLLqQcwv4HSKC+iSjiOUuAmP+kKPF3CxjcLAH/4pt
7Y5Trth1s4XN72sjyHnMIDGarK/Vu8KtaoF4YE+b7ilhwDwhUnlhqlThs25b
43dLil2xi8nSlZ9x8kmAKMASfEqPWIPaiwlP3roVJRx/Ev68nlhIfB9yhx4j
ow3sHX9Oan90m9QfKJbRyPRlM8zGCV7ldpijtx+RIpLYqRhSPFekpnwJjpGd
WBCbkkyv9h1dxcV8geyPqZrYJ83vHrldzM6/IeoAAUBMPsXBaMjNb5sYgj8q
gQrgaCdAMQPeP4P93DvAnzpCdBIEVhT2ZjuF+w3HjlynvVLlREjP9DJWs0ET
sn7vHq2sxniogvimYgYRBGnVkqU9PFFgoDwHhSGcRtGjtBck9ZDFENpCRjq6
vEaNAwvskU81LP9oSGpt7Upt6YMHhmf5+EiRsB6pucFUcowl3CSiiwWgcPv3
M1jqryX+ZRZyyuZD02ts1l787Lq/dXNkgrEsBAuNOLvm2pWg/8lCj6fBBI3O
8olar+pK3Ib7Gmd7qG+pNVbDItPC2cDBoJ11GjkD10FPCzeI1k9VDoJLw2Fe
pJR9qQG6OfaJbv7ETGE9JQE8+7wpPjSVvF9nvr6xaboQi4R4NsoUo6lvFvU2
f7PVJdAdBk5BbSK7MMMeYlO3s6hsqZh2pfBj0RbNeTUVaOb9ep9tzapJX1FR
+FHM0WWnEvxB9tl0dK3o2gQ0t3cjdOUn2xlGzdAECyzffEVXX80ASRHsZkpo
LcPoEVt537CuE3bjL9yFOEIHySRzmWxdR3J+QEcDSXz+AYEEok4nhVjmBk7m
gzJmlHRoIpKEvQ1CZPLJsX7LZo7RKliBfr7QZt3DfFPNUOAjw0QA3uUJ/5V/
lseANXzmtzFIT4p4WalNZCS6EgbuLlJpDvkAT9HqKPcw5An8iVPgYz5Zv1Jh
df7pRkpm4O0xsGdoZwcs92Jb4HMBiUB2BqsVz7P2xUEf7V2Eo3dYU8U+g2ap
M3LCDtZbj92JqLKBB+a1xB99HqrqjwGxxPY8BFfAe2aMOWwlv4HW+9bMaK6o
6BF+NCYyK3KIlEkTSXCbUmZrsXGr4fv1wpRffviDEHKp0ngg4FXVAHngiQI9
ZqFDAAti4MgCcOAy+A0P1iKlgOlNOM+1pvEexPaivorNMjmwrmuiPOtaYwBF
d1OAlqIPtn77TY8ENgGHmgJQU2deo8PmXsyifkEqUaHtQAy5SMKCk6jJe471
7RlGM4LJfRCl3j0Qp+svPMlaWoLUzm4fkTb4LuiofAX2MaE/lSzQrWvgdyQU
gxw38ZNXo4MLkoW1SJrliy37paLPAZXcF1heC5vCZxSC0jHMRa26CB/qyLfW
9Ut/aMYLPuFJMi3xmZdJYysTerqcNfXPslATgM0YDZuGODJ7i2agOJ1S6Wq5
eSFT+MH7ZVIB9yLGAl16frQ1EMsPwuWMUzBioAWOmOJwymxnR0r/W+7zfea0
+3691M0o8WzyjV6rSoiL9t5fwgqdT3Y6avnySlmsQ8dJrdDakhgjnrG+CQUu
/sjx4U5vxiagGDL6QDfR+9EDpeRwii09BTzkDPUIePhlOPq7aDXJoXrhzr8C
8Xg+vPLbRzpwWqkbOD61nBLsaaFwJe2jrfO56WSSmuluLI1CVROaAfXlxCJp
TLTCvk+PmxCQlNM99UqIAcut2JfDOMB366NH06O1fhPlBjfmFjW6wAfNn9iI
dyt+wdjc2AZPHjrUEfCf+tBefFnRYNwUTN5i502x0LDc4qSn6wgqRpMNylDe
L5bVqp9ef4YOT7+iPQ7SHaCy1/Fk0Xn9X00wiZDqZLL6yv86hZvEjMuDe1Eo
++64Sf1M9fcp+qT2BHdmMP59ZpF8NtVTX8jOaWQRFqR5xIiBbUpQEiytTbFA
DkGTJ3KBl394tNmm+I55uilwkzhf9f/vcTaCDNVn2ZNOjMevx4o+/Avsj/5h
z3zQXvkMg5f+ysiBTH+ST5XpySLVclDBThyBtzlkFatHIzrIn/si/sF+/IFv
d3YzZA4t2uexXM8q/+bYx7X9Dd2aB4MJ/AHJe9MEYQWloUZVx0fAmxozsqfN
XOtONw1m45b1iPwRepY8ZWE5HlGmwS132nSDTmHxXGscARdAJfWLSYsrXgNx
rcxBGxZmcXSelO01fupdc4oT1ddGkFcb9aUvivIdeszzlkjHjTXYDO+H2Ftl
jjaoF9ePQ1QoklqqeJE5ahp3w7VHtK6gmQowdJr/7ni3UuFsVP0sGjbyIalg
hzgaTR/ckef+BTatoYskmanWZBWLkTQhrf//bJuFBU69L93NNJWLX/hNi8iR
rNhlRVmYqKCB2B4BBrBPg9PHocKOBgUWWvT1Iz+P/ExJ/eLElkZU7ygD2arc
Fk8uPh4R4n6CnjqqmNsPh+apBqotdVWlrm8JANZU3aj7fEM8QNpHtqvwxdjV
OiUDkz2ym3kI2mL7BBR3b1o0fj5BYxXuNVqxnKd3tHnTQDeL4LP26bzce3Yi
1TBugEeqKv3NDvobIVu+FRbKcmV7PHPH26d27qY6C4KSX1GnIYKzSBAu4j++
CPwSZ3t7NevaVN3l2FzQdmfwCRQTGZIa1fTNzaH4hYX/uka1e7+tkP4DgHml
LP+ulzt019zzqPGUkHXmkvWnRj0sC9j5oplgXq9nOiehOIkKnssVO58ca/1K
9+xQ6cHhoeDvnNaDCLE5OrK4fYUI+0vd1/ysAmr6eZshJXF/IF3NCJ85csi/
HjzB1bEZgt6zWL86cTvIAEAoGmXyoZqAVkqfXgd+BYDLP2CaF4q1bfPGr6y5
1tg95brY+jwMyqC7jxdfAj9CiWem/kua8TfRIASl39S60ScjTRtc4K1/JhzA
e29bALWDRWxpWqhYowV1+ESkBJUiKkJcLdH1sMlkiHbxWRs4SfS5EdiDSZ5h
s1+LlVF1mgdyYbXs6rHyXH3foFJCyGN64FTjTrkSQR6hI21cfPoDclWZZl//
GHO4TEvef02ZXiunTqUG1cA/K5kg+kZ/0btx8IoCEIfotTKC2Ted0PaEG81j
PF4k5pAhgcwVNAJKl6iyTfhXdIAFuj/+hw7Y2szVw+Rf6l/1nQvNInWhaosB
TVwVI2MdRKFVQ/aogQeCsiBMiQPXJlQoSzBS9hyiLtzYviNXFIQkpTFnaC1T
/qREMsNag4XLZQfvitHawHA6AKFhuMUm0VGIjq9rZtI/7IhZRnGh0AxrvCn7
9ewgYGyOxUon8qpfaWImLjLXUjjhcMepNANfA52gQlxnNswXAvmAiK6N+Yp6
jxGqQ6YFaMIm1kDKzJ/KaekZ4uPyGSMev3/YL7bp2ihgm4IY1TNWBK2e/Wc/
uMDDNkF8AtxTj3mTTJHpEVB6B1ZhLfnkLtHENSEXWVFZwxSqFIyQsp8MT9PM
wzr21BDFpUHEyyo7xh60F9sXL9pBVGZqBhqNXtV/WKDS6yQogS+8VrSBv58O
l7iurEk8fU4pH8qiI+yzZLHWNZ4TP9UQAI0QFlWNojv/wf4tdStW41SzrH5S
UQaYcEsUJLSKZ6e3+ym5vrE383pUHFEdq2QAxe4WrOiKwdEAieOlMrg+pBsp
rb+97ClmroO+zlVuB9jHB5pbedaVnbY7tViaaiJlMYmQzML8K0MVTihG0Eqc
t/TWVZpjp1JJ3SpwlYSfrYyIBenTcevZEvni61Afry6TpeRwQEuU0pI3ktDO
S6FSl1uHElaTbfTcd71XljNhSMH0B+CGs48R63YTS1mf/AZpxUzSEoQzMH6/
SloAZTMKSXcUFlrfmgR+2bslxX1mn4UtVzm7V6ojUdKXg5aEeT6xJHh3XwDz
IHVKUa4PCV5Vat9RFpoy87eku7Kqs3O9pq2oVX1eF7vOn2A6jPJcbL8BkCTJ
AqQpJCr5T5dG7YhRR38Xnh4W7xTax7NOH9Fwa7uzg2R99o2uIWt+n5ZQWhKk
vDq7Us06USxns9ovfkL6s5HnK6uEWf6td0AVo+XqiD+6a29wXOewnDCj04g7
HS59R3ayQw2weaA1leBMrKnpIiTVsuKcpRraL+TA2UIAN0sGIz014UxMYKKh
Jqxkjb9hyuMr/NJ2PB/Safc1JDSuaunKP26eBUucNMNXWjyfMmxP4nAAR4nc
54vHPElsgvtXYkwY8ec41d6kNJ286TEGy4gS0q3Xn6lICeMsQ7Kuf2wETDVc
N+Ewww5DmSaXxjBabXCx+xckCPGlzSlGVlvB06TElc+JfBdmhsOn+zvGJb/f
oo8PtJVQTj+k0eEF+hfL4jd/HLRgoNZdR6pxQzXvlBopmvTAbY39P0n/JU7J
aJR5/dDk9E6N+zC5G0aop+/+0nia349OzkfWHdp4nh1gqFogYu2IQCWFHY7t
dVeL4R3EAl6JwYdQsaIDLYnKfdyWX3FVo5JOJcEgQy3UzOwrIj+jyk24Fie/
pjw+3rBDZALdq3nvBzBxJshM45cIat4iBB9IkS5xxd9WoPRfv0xhhUwynQJE
6dA5e6xo0eD8pEghJjGcqLvSVAPxsPrxcnVtC5pX+eJhHwhBIRyt0EEd/HwF
59qrgQjrlcbRcdRujo+r721xTrEXcU9kMKDUHg/amdI/Jogf7dmYpvk7wZ0F
k0+f+6XPb1hwOvi2I/HTzvcefb5h+yId0yme+inxZprgzGmyLlahKqXdDZyB
Bry6VRbqgwYQfpJOylJnKyMiJR/uQnTk5P9y1MJ6rtLLVbPqsXcQ3J9j7ORa
d4eYw7q+7KdhSL/arIhseQAStxwMJpK69nFCdBbX2vDMlqZWPF249ovdbOTO
zMHfwK1KTa7Nz2YVbETdWYKN8sVYvMCwJeXrsmP73AvOCneJuUQUR7xTfDN9
J1RltUmGXpJ/YSkisRAJgtJTpzqQ9h4xbVOc3bC4ynZaaulUuFH3PHC5+pPO
jHhCE05UWIg065oZ3PeIZ5MHururM3h2Z8cXpcXH/XUupDvUTFP5fJs+fZFO
+N1q7d96LQtsze+eh09ZPnCfZgua4yyXWoNUiyY0eNzGlXgR62X+WQa5xWK7
tTxzZgD9m6I2Oghz+IDU8esS5SR2t+CKumrApD6IYdeELJB4HDwwqn6AuRPh
D0j9V+/UnByHeY1mCXcVAutasN518uFUwJgEolBZCjMv4T4BH8jDPGWYzATF
IQujLfvk9kaAUsuSIeJcU5PgGYx1aTcMbcuJuk3TzyIubGy/db4kTMm7NkUX
qmsLdUS+L0+5ACsS1hR6jcdEvekhGRNH/hX5x9ioZQZ64M4AUSTs7zoIzLwZ
ojhVJWLmxDZEoFZLlBNbGAakPDV67WcqJfuwX3qZ9Ucas1BDCV8pploJpyQ6
X4NFQUFgC1B1MPIHEwvyYRZ9MQhENlSYrgqKTt7xTs4VxknFnIrSnWVs9O/+
JLX9CQd+43AoR5ZCUdm8S8pwCQPjJMENMBlNuknSmd+muCe0RrN6InlQKRGy
Yo0BEYO6S78+oeRl3iEnp7r6C/GjcQviT/L/gRWm5CI5zhtKTigcpYusBDIo
92Y6SSGMMZRui53mhp7wM/HeFpq6FIlGgCu0zXyFSQtSFuuD5EWDJbwi6KKa
b6HgUBXAinQLHleqLxaJbtL9e7e1S08EZsmcVzEatY3tZ4CknuIdrvptAhUH
U6dB4cxsH79/9FjBRJ/wdFWXkIXZb1nJYw4dkz9J7x9WNiMn55noPxYL9Qxz
6uATVTqzlR1CkdApqgFj02rOLuwi/1R/j/eYG+hTW1kBxVYC25odLy/e8HNE
kSHUE30PBLhkaL898MfG9ZOMEf1rWfdDPs3+4vRJIVrarUPUN4arfuN2UqHz
37e4vhWoJ+zsZvF8S6VykYhYQeVMLmekw57dxwsFeUbynD7fFRQbxqUWL8Iq
NE14siVvGba+AmSeV3Yc6DYdFMqYW6134eb3qz8omarNAJ+dW09Av4sgyLOB
zeBY6tjX9Atu6FaKhdwWEsxoK875LHRrop5be3czql93hMkwScP5Da+YXR3h
+6206mW0cj4PeAsWzKk8WH+PYm2iacJdfj06cPJ8unpYJnROfppVzKvVrO28
HSnVkpYAEO3UPlMLq5iIsaXewo7qDpVIOx6Gty7KKQZ9X6Rdby2adk3G3baG
FfbPSUQ5EIYC/KOWk1PxhB+xD9fEkI0o3EiCv034gnuRAkZtwZnv2b0QcUVi
0TavxF6BobLEeMqc2IkF5ERho4wUEHv4KGRHb25/JdFOPPUXG31pCfNP+DHp
7NLKXvDpfiofJ4DzMxBufzOlb7k139ugLeWVMysAKqL/IQb5QylbHplOI8mJ
M4zDNhX+skLA7KHM/KunbGdHu1ehrPGPEG51V/bOMilIm1rzwiBlIx8XnuXY
iGyv2ZLhD3mqJ27fSTSgYk0yHTFk6/I3+iUWxnZfU8F/gnyXHWouftrFwj4x
WWW6bJty5oNVrlbS/0b+FlRpMPtk8o9lw83eNGvD1I4NBtbfiW20USwAdaJP
/9WY96kyfrhDyIj7hvvV8icgjj8HEWs++uuMtWxHWa3FWqG051A7W4MIsFu+
sXydyijj3KzPqh/3Lmj20VMmzX+t7u2yPImiKyuozA6wodrQlBlvBa81ifcs
eNBbeRHD+gG4OPEplwReAPpyztP0Kl1s/Tm6U39tjhLgwq2BnLJOQiGcX1E+
mVPobHK1Q12N/140+Kz5u4xnc4CZBbcw/BNQ+xS7PLPgEF2vSNFf0xz329Wb
YMw8j2JGBUoJSSKeyUa//X4Npxb8WAsFxgrAHgAc5moPGZNr4y27UWMQ7aYd
yX28Hgttfx+aeAJY3qWopg4/FP5leZoCbm8aly6kIAcOmBu4esaBWovtE0oS
CcEoEATQjNdvgLcMKTzKIh9i8Poyh0muRw36WpM2TBstSuRm2UvIlBoGzyu9
igAkP/UDov5LHHx/pQnyBLmOG8MpIyGCBQePRs23Mhtekog/4uLnFlGPyIU0
ftMRDQaOfHtNlYVEDuzS5KjwBhYRJOG+yXLrJDsrT/rZncB94Ya/qPyRYvI2
taDu2KKir5tI6Cb8jSn4XjTi7Eke85j/2kCJwF6LC8aZOvU4EveHQE5P8Nue
s8lkcGQ8iX6s3esROv/P5R2LpIEN6SXIt+fit4e3OsSEv+qB9J7bbLE0LO3y
M2StmMYEA1TpExxtKKn5BoUoff31D7GC6Xx+zaKKV7WqrzA6qHb9ATbQDkza
pJhvJX5JIn0MGmrY2GP0ZEOxtqF7VvfYlHnIZ/Dc93CHOtMOuqo/qbWA/4Sb
Jhu654XjYe3MsfZvt3bDcvUGhNrYxnhYN0FG85Shbiby2XKwcqo3KG+ka+av
RtrnH1sZVIphYEyfyKtRhnTXqkkrbuWyDIq2GBYrF4YujvVCEzm7STg7c/hR
SyaH5ya0pTN/YgkZ2dg/FVHdszaxoA3p1q5yqodQ56JUE47a2vSwkUdiHVUc
UUN3xPY1NIjOsb1oyxXONTVx9UJSIxMxVSH91aOrfPtQIs9u6MamOPbkrZv2
hyG8QyhBNioSWMWZcJ2bE3CsSEDn2fhNQYw3lA6cy2T/+HfuT6FT4rLiQOlb
M5inmgAiTB9G5qNt/pkHjczSltTQ84WPhVOgN64nEaGgwetx6srf4XnYCulL
AeHcA9yUxiUfkL6ShC8n1TYkH+ToL0k8SwCKdjmQ+Ceoo8a2l/eOa5iUgiLI
moGzBPA8ZzwX12JwROYgHsrv3GyKhlaLpjMt01PVKQgm0FF6RYzcgWqxtlZp
/o+7b1/HC1/lPT2bcQjdG2lI+9hLPA+pfEed4udvpQfGk4T3GBGsl1epLViq
rRQZeGpWkHdohCItZaa30WHT9vJbBgt3sGf1dptmgPGxaDwsZRQ3zyZH9y2W
9UPKV0TaLY9K6G7t+Ij8xGhiu+YwhB6j0vI4EAQAzGctv/1SQG6TZJ7dpnZQ
7gX9H5WgH1d+miaGjebrw+W+d5VQTClWha6DV8pEgxWT8cAoCLDYEhVkkbgN
4N44zOGdVxgTbA8gLS9uubMmQJ4gLFhncfgwYntVx4F6mmpNyXNx4JSoqNlE
bYYzh9zp1KEe8a7LZnAHb6aqWhZlweC3iQSpJjzklufuj3ICLNZIwLsREZNc
zg0F4Hayv0Lq9vwt129pQump7UUEzT3KhN/IO0iBtSQLP8Ve47oHB4n3O69l
tqBbHVpnLi+6b7pVQFgl23PIT6V6Ru7G2Kw0ynKCDSlLbweZyykJLjWtV5/C
hXYQhS8MHbpQVPsvpxhr6B5z+DIqXH2487aWHr0pTONBIGz+Y5Jr2Wu3pi93
L0U2KA+rRAJX1PhEEZ0RbE5fYYDmBzdTPY4SoD00R3APsZjDSylROIeSLA2l
x8OlA8pxAHfeQJBbix4Df9QiSFcTjU94hoSIoVJkp7jI+snXUwIAPNutHj2d
UfsN9EosXgJQR0ocLsAqH9+NQJTufumxom65mIIPPowEPw4/0c6v3YLUyfBq
Uz7MeVOsQ9cXtCGclvFSp/Seaay5+70bg+7GEPF7IC07ziT1eeMwXy8YDJjq
vHLNdujiMe/Uer+naHQ2+bcHbPk7g0CKKBuh9gRCyFd0aAW49/wezEvfVE43
OXjQCPU/YdHrVFLfI+175gEv/kQE9XI1KQo1mAB0QhBM1HRIesVyEZ1Y2APF
nF87lDNTolUsNflYFq9VEx79gxB0JoCto864VeMd9p+AM3fJoB/5pPxSKykc
V0/0BJF1GYK51FKXrIfgEeqGjrc4D20K1LCVJ/EiiPZJfHQa6FdqjcrF3L9W
5ZiQf2vvz0w+ZApuqQXS9Pm6m1z1DC2K0qsnF3syHvNnMOU0EfofY1s49Dui
9zsiboTT04s1ohJU60A5P7JCzRRhwQqGy4evviKgXfs0adXfEkle3/bts8mP
6AlhrtBZigZS+hjNx80HyB2kSsdzKbli5WqfJ97Fz/qPJOFj3z5guJxyQNTV
Rb0joNjx7+1j+kFVUasxXnNZx+xW9NfIRNYYippkR0CXqVL1pvhbMrpdZvPn
fd0FeS+hgHgNYgFy8rJxUyyhztQAUnA/Ejv3f7WUFPm60O8wkZw6T0+psx5j
OJhm8aH2t9lrYtks/zcCPSqcfQgBOo/isr3+CCYPcWFv4kgUQh0otgUK6I+M
y9PbbZpWP85IeQmkVU9cRLaIZaHBcucGl1Jh2bSIu2Kh/nhrkPCqW4XdolnY
C5nKlSwZzQSkzuNZkc5yzKeO1Ni0cmOJ0zrCnpkt4ETZLtqEmP7tUYKggOCw
y5A+bi9T7/HBPh/Qx+36uQvzTL15E8MOPeUBuWQ/t5e+4A5LXYA/UCBIYMFC
P/uF/oDGU2P013+rELDh8Vv+WcNONNFpLQXHMz9GlsulCXLpoBRbEfLw9s+q
w4PlJvP6wgIIIu6g7IgSWWQL5BkFHzQL3l+mCuifwvp+a2Ztt3Qoel3LEIMv
4JfXVTdxke6ZEA9kzCOD3KNzS1V9NW5Rk9exeN4KAaEYAGK8xJT09g4+q2zp
oDoswWkN5L4x9XFLKvceMbayQd54PRiT2w6BxuoZfPteRbfyXHRLez10GA0B
sFPukaActJMZU6Tbk8TDNC6kdJN/R3KjaKgagYXLt2FG+GR8Lg2X95/1jKJv
vFIjK7CAUJuYs6LL7nSHinqfjGiYazCKpOeZaGdoA+ehnIjbHGPxJ8Qg6IJk
On713h6jzKLDlEvDM+hO+2HiMH07rOi3bzKyZpIsa5Sx0hd2C8Dd/oWmxYs2
HMVpChr0tyMafuS2+PrZkTEIEpZ4FHkZhEhHLqd+DEox5G1hw6h6aJQmurqV
XWog5ylTyEsb5Npge8xXyqbQN0FXSyx8qfRD5+Wh9FVftg0Gyyk5yL9H4uhr
OtxpsIR7rROs3YteD2gsLVZz0+PDXmtkrCl415rHmSnJwpG12AXvpf2P+ZPR
rRqxrGKR0zfPQK7DLMwTSZZVCn+JExX6WCihRrXWUnlVOb0SOLPymbbxl6/F
7ApiEbGfyYUjMuOdvW4Mm4yxeB/EIcKa6tZgF2NcnBw/NYmQ9p421QSqBPnK
RFxb1M6/x0qyiRDODzJazrJZMjBOrp7/LwEMLAWKO3Ih/vPIdv2Bb63HdUoV
pFEoZxujGhBYm+ANNtAt1M2sIftb3bx8I5FMFCPCS0utPxkSmcNIDzCi/fuJ
Pdzx+6XYZga2Y7qrx4gS6ZYQRbE1rO7oJwslaH0s6djT89L+J7dgnfdJLT8x
ewUr87lH/pbWtSGFpURHpfR7I9IjwX84lodEXB5bjNqxzqUc4qAnnhW2Di1o
Ii9sVflY7HDiGMWK6pWXcs7XpeaEp9NCtOcE8cm3Qf8qVtLLsPs9BqNiWDtA
Vcl+NWv9OWeWK3riOU7si15qL2zT7pQjF1j0WhN9iuy3psYvcFPYx+lQ2eF8
aa3zrk+GtWD1ervJerkn7tRaC4ll1CdWpMAjsaDHqZXlc9xOp+sbl4sPDlKa
8lY/T8iu3Go2heGihrhrkT0CoPIWUvjsfkEviFpbrSx6NkX/dqtatJO+9X+s
CFE9gf89rJtINHVYeft9FL4cKKsVhetwzmXHzqCVOsltZbAv+Xw3T2gTn/l1
Up+f/ugcX4ZltOxBl2vyEwnGX9G4kZclbh//RrYC15iOHLEkHqPoBYivj2wK
tv3cFTP7vm9ME3qR7lCfRyhPGoXc+dQxtH/FumM6M0pb7CeruFu8nllSa7Ba
0Vgl5S0uVUUjfRXuRnERc5CllFxC7TL+4UNV2PtU/LjyhPQjcxK2jZADtQdS
VFNcXt0EVUC4S8rG89Jq7E1UqiGRi4sZzRlvYSyq+IXwgAeIPx06ZfFC2wtU
TWgVn7EQBQleceEh+Xxz/GY/p9IGis4wJulJ0POJN2hmBk85Ez/b9UPl8kit
aHP6AQXVMiPs/atSJ1+E1+NSaxEZwdxuL00VhG58T49cdISQtcBf9cuET+KW
aeyUKh2MAm2DYNXvXdF3wwMD+QshsL0333T4vsBtjKUfYKt8oLhblScMH7wZ
RFKNTjKK6RToUgjyKrxBH+kSrbMBZKg7rfQ/mFWqdDepz+4TZy97viZn7+dv
xaplNEuHv3a+d5H3C4PCyrT7s4rXEfs/iG8FAv1aV5TWiKdbl2VwVkrN/d8/
rhKaZrPuiZrhPH6zce08uKL9TAeMgMFob9FeMDRq/SZvA8khDUFoWJHsS37c
jmYWW7t6T/AMqWb+FqQd68g2RFUh8G9GVy+Ekw/f+4Tb6FHtu6Kt0bilHLzk
3/zUC0TAXJ536xIM7xJMnJn1Q6tZf/eIX8hNEFNswY8u3/U2ZgLX+Ya/5c+p
HwZSenS8dFQtP8wfVpieaOt72Cm2lOZBdyKNhaN/FJLfaVtVvsgsWnXJs0qU
8BT0XVwONjzMc03dS6VsLAffHMGF1EVgSUEfEd8CauQTBZIfSHwPnQG8Vl42
A85fmFRqE1+Kl0xio48GTCxkQSE8nmIknATKJtE8baeyRkFtgy18+8+jY0Vk
67FCaDuMEGoOoiBiQazXrdxHJ3Jx8mW3jdbctBVZp5QBHdYHBPkhc0AqbkkX
FnW1lPi7LWj5OUkQh7CrlHjw2vuSDp138cEV3jyHuuJv7cEWBJIjtGbM3ou/
RXcUFrWmEZIyAOrGUap0SvyF+0L6hn6jTqTHSg0iEuSZ2tk5htJ5cOF/EKcX
jw9YmIKt6kAJ3HLgx41p/ogLsnc3i06Sf2ZYfV/dPNagUB5wzy/bp3GtqISs
kl1yWIjXaB4EEBFEFTJkEV3qAcM6jaqjS+rTZbK7IXR/+xQboQA6EJSvSRqn
/ryKFX5wMmuvRvTl6CkhIAiuDdFq2gnD0clqv4RxyfkBO+UZeYH2fCgig4q5
8g39eSU/EQ5Pl+TfbmhmEjypC1ZwiJE+1+CAiumkUlue3qMtWyp71xTgIebA
dcC774oTLs5iU+UmOEUsUD8le+ChjzLSGjVUr+wRctm5eUshBzwW34olyc9C
USmWc3ILdJDz+/YV5TbNl9nMNMmUu+2KqWiz+DnWQwPS3cpTEbx8AgSLyLSJ
VMzL5Oo5h6NmTPeG+0yCQpLOJNXSIOU76uNheetuyazrMpShuHYSQDXRe9QU
5jIWXhzxcYhtgtVRSxgx/5j8/aQ/oItCIX16Ilva9aiPrBQRvfobM4k9ZxhO
0+ndQBKR1rTNr8uUtMyAwLfK/UBVPWVZyRHXNAyN6z7zvzbYpBR1xfxOjXKt
k0o97AGHcJv1KNTCWiMb4UV7iUfxvi0JoUTLADdybyDLfMBzvHkjaQfP2Pm2
/S7mS//evJvIWbece5t3MlumRBoYJ/y4Biw1Ii+nk6+J1F0OfvnA5R+5ROKp
NrbBVWHpfPomEZDqPF82J+cTQUet8LlV6/U9mAOnRCsR88amMXQ8OEVHyCPc
AAoIXKO1e5ljL8uGUoVq0Rz92YQrcrtxRVSNrzYS07rK9ygRbI0NeWuGvkN3
UE5L8eFp5w8jh5Ol4OrWIfLFyXiJPX5HwY1aPS+GivYsk8Ugp/+h2fNEY1GB
WCqxRerEJsvrd1D+fEgN9ZJsY1QT7vI4YG/dihO0PVhpggCoKhv6iXynWmva
LjKrq2XcG4pbuGlLSrOX+o6aYOlDN+SMYU8GOR3VFrsroSDx3Cg8IomdqYS/
b1j5qHwoi8YxDRq+/VlVNgdz7WpGvPUrwrEdJLvoCtRkRlxZaV/gxFI902LK
Pod2FdOK5C453mH8Cd7oR/9UUqWBg79KbgLhgmmjoaFvVhYzXdRc8PD/UuTf
g9InHc2OPyy2hYdsbCtQkaLqgi5gYwVFGz5h2GO4Kq2RZd3oUYxJrmuO8RlF
ZEmotVKMR7oFN+9aufSUPgqlxy4o8YMMDuQykApBqZFW9tmevGO7jvRguRGI
LTntGUHXEEeRaEwCT5dTj1BVFlgSKbXfzaJpNKz8/kdXHFcQAh6D3ljgvoqV
yTzlpjNrcbjlnFc8nK9SW49kxlUtAoUnlupFvyRoYjZv03oeIBntFT7DcO9/
WJhtZxK/EXYV3G/UODeaaN1C7KWgHPp82u5YA5TkZnm1vuUt70+ccHlFvyVJ
Vhdzf3cQWj8HV7XOaf39i6HMzqNxxLLB7sP13FryjZs9EOWAaPdK+nnqQ/tW
GaJDa0JXe16TQqkwa9ae0p6dd9ZdVJz1UagLdm6Oz5w+0nVIv8odDf9hBcTH
HOF0Ngk4epEB/TumFaVRF7Kga1IzmoTYwGjFV8E9e+kSBKKgZBADdsqf3Tgt
rlKVvzJTXkj2KktZd1xqqaBtNgO2HqS+76dn2sQ1nzsvh2gfPKtFrag31mja
RtFrsss9cArJvxgk3SnhrrICPqCoaiyJgL6V5j2gbGHGc/6DOBAnJEMo5Ko5
uj2a45AXGiGgFF8IFF7uRm8ZEuRz6Fin2IOpArt0CvuKk5+IF7eEG5ruXquB
ff8FtwEGcoxV1IQF9msbm9YeDnKJ51J/JGhiSCRX+YhIk/xOs5r90tqLfzSB
rWldoFzswYxk+mZ+tnW0m6PMprdn0Lsx3DYVaFEGobyMia1jSqnFQNJyNc6G
AABq0zHNBsRTqcoVljzctCBYRsomgTFWMBWHdskWOkVlBTlQq4W8dGzjIefZ
gWTqot49Wy/c2Y6v6oYIkIFajWnAp/7KDnchOj09/2pPuY7ZMLCzJrq1SntR
QF4MODNKPUHJ2bJHM8gozJMGSmnsGd51NW+eWhHA9XEOCIO+/VoDUNbudoAa
08BmU99VaxF0RQlXBNVoYYagNNEq3LchS1MDNXTSstoteUUY/ObPHzoJS/FO
j/675HbOn0fRPhxDct7w9sEYQe4esgIsNLOwD9czrFIeODNntlF3PHn0FsfL
v0cjnH4jhLwWiBCK2BPRUnQZuC1ff4TLaJ489Doi3+qq0R866CiYvco8boZ8
95B/FPLku8dmuo+QcYBj9uq4F8+ws81ezP4XdZ4t6UHLzF7WGTwZqX+dqrcv
qKav8xUXYgam7dAIyHWebaX8SXI7foITvhJU7bQ85ldjsEGvmFXAJWOc2fLt
hrlNNZ+jE3hqWWlV0FSv0PFGzenZOCvv+ASXRJdi4kWAGKJ3Fc+Hh04lvbtg
RIJ8X45axjWKXEaDyhSIwSKx1Yw329Wjcl4u0R2bxlpq/mi8wqcVIbiCLQRK
rGmchDfG3lYzi6V2s/5d+65H3GCHqXK89XaSJy4SGR+mSNpFu9u66kocQgSu
wx14klmxADBXrXIBuNR6uIJumlepSQTZ9Zl++022xJQh7cPxJdtoqTbWY+9S
DDGuL5zdukdoenoLywzQ3jt/GCL3XB+d5nM77BZ7OWXRWDxtVQcXf9bx8AsF
Un8RM5KhmRjot1q4jmR93apvetmzzteYGA38BQDKHN/VCNd1T1dZ2Jxkj/eB
MYpJAj/XbwlLcs+0Yt5qgOaBkXICEJH6XD14DGNWxcYMXYgYEpR6n+4TVrNr
LJMzaV0t7fjfK563ltTBh5jgi2LYXmZ3ILBxaNBEGd8VRKm6jt5V9T8yY0Nn
FN5SoT9sR0PUwU1x/1rn43wTV868kFXgLQgu7UiC9/b0RqoROPGcII4bwWkn
Jr/Dc8irYep+rGlWHo/IlKVRLa0DG02ZHwR7xSuqPccznJPaENAVa0+LkySK
VvET2AjlKgSDzs34LSTe7B8pxf+EBKfcKTm6OC1Cx4SxQrvVsSTWs7U7T7pv
nnsPq5U2ws1Ck/fuKsw2SwyWplO6xSgyPHZEAu3EppkfxvQ5is/vUiES/nuk
ykITREembKV5aCQucFo4/TSCLE8fWeuCECXx3Cj9oE3he6dRAm+Irwuvnirl
+H7K+RfRAgOXop3fyv+L9WUDIcR1C78hTH3wyWNVTAaUMch4HVP+E0fRW5in
702vpOA+Vq0H2FSVsOmKC//9dMIxErpP+oDy5JD7p9a52/slp5pIY+NrXca6
o0yJ4TFtz1tA+QAUyyAYd34zzvVNgZ1vL7ko2ruiEFf5liJnJKrUk4vb6Ooh
Wtr51UmAWmpyIVrSOKonWGwG9JIWFikBJKd+uXJpcRU3rniphDTVSJv9EA0T
/H7Vv7oIL1EU6b0IqcA+ZTpT3itie9FLGhP/epVKv5xZ7ZZfqJuVcmLVjWws
anc0Mf9yN0a3iRYFTyT/53XABeofPp69/HR6DTsuVnbEV+lxcMuQNoDS67S3
v+GSOtOmuMB62xSaXRvwUo4BToPnYJQ6o3PseEcaJ2TrW93cffh7b0WhbqOx
t1TRty2cIrvSith9DRUGvWHsDFO7hXyoOKTDdIkLICmlhyF9qdHTEeuYnNWY
7TotFWpTQS1onK8Dx3ugTCvfzVl9rMoW0g/ltEv03zY0ausml6QVnNLNP6e9
5zhm054bx2kAezfUIMVT+vrO/OsT/a2aYA6bV8uvmrZv2UuK9439gdoxMo52
QAPkmvlKRTmUDZ1mRkTpmL4VM8r/Fe1OtMHkgsdK6TDjHTd8d/w4ZgyR5MHk
HulRWuktUGm+5KKeaBdXbLRDjDea8+RmcYfsYYQ28NsVn5n6W3lr2kuOYnbe
2b1xOiqow43tC06NegfAjxq7DJiyolwyQ9MxRmwHKICK/e2cYRp04LA0VkSr
87OZWszViWHvyW9qi8dY9fdKR4AzB0cj7SZ1BSE0NtlMe0PIzaxOqZIn6Tcn
rFyAGDrhiBT25m3izGx4cFVmV3ZkD1vFE30hhiOGHyCNSbtU7U655y0gGYpg
Mj8zU2Vh7YI6giNVUHATvXEWSn2tiCE5TMV/vdR46LappwljaCRmKw1SEMY1
kmTyHqKsIjjsudzSlAM1MTviKjhmFNCmKRB7OiRIButFVoKOO1wK2y8fDME3
M2YVXqq/3Q4QrFrY1Ny+rrEllNVyOKASJoilMdh3C2jLEJ+dKo2V1S0t9rWB
QtKnJviEIqitByfjlXstBttsBr9KyaLMBmXa9U+A8Jn11jux9acWpWMghmbp
dXl67igpGpVv+oU2DM6m8EazeTgzMN+HyFbw4ALNnW/1IJ62Odu5SQZNEy4a
6KzgG3zmhtCYarbIH3kNHAO3AsOg4Ynh3d6J8btR2jtqoYLk2J6YJp1JaQS5
kfC/zg7L4WQForOrCZAIovd7mPxeIyWYS+KQEwtyCeWhMMkcpXCaqikujYNN
zYIotUoVYjIGzKvOZz4yJzq+rwSkif1WhftcOL84IfGZzDOuqUQpTkUUcQ62
2A3uD/2O8L5wRIAKcgiI2gR2VT6nwlgADzEKEgxJWWl1NU7jTnT5BCbOxXSO
G/miqw/cCWNZIvlznN1Sjb+RH4Hf3Yel1UhQnMaS0HbHAJF/4odqvdeV8gVA
gDZn3sFYq76DmZR1fkGAvqdv5wCkj2VXvYVFAIFwCrdpButDlKQyZ2vQ8ypP
fAFbcVGzgNOjTWi3fE00dwNDbObhZb6PeLb5Xr+/+7KdJaoxhBGPNyDEx9mw
bJHqtHYEy1iONxPSS20uWnxCGvfBm6d0auRtpB3GAf/RJBvhjv7DwrGpViSx
G5Icxlp2NOR5bGfqiy80x/IIljZP7Vdnln4Zyq1AyVM/X/Ql7RkvKxsb/j+Z
HRr7+iAhGB6qrGty487B8XRcuCquVcSUQsGT+oJ7XqM5AbcAvEo2FwaMmqba
wNPKrhClZn5qGqrKuu4UkmgDqL24Y4D5GtfFg4Q8oeZCgqGJpHfAX9/Jj9vm
sIMGtCw+YOxRt5hZXdzr2snGP/i8g6BR+f1XGXZ3MHC2e44wK/t/7/ufBnLo
z2LkdxyaUH8FMR6kgMD2CsM+i8BrqIOSi45C0Rl7NT3RcdUUfUM+qHPodiSP
dLT+fXBncu+UKvsAFktGyf9P7AxRHCnBoM4D1MwxN4uiCU69sz3D8fvja9Lh
UO7CVCGmGO4UOthCH5PJ6lpZzslmwvw1vQAIvMM6mM5ipp0mB/PcEj7KxHpm
vZDYcwnT4O5CYAceyONMdNkJsCF5VtWSDw4BX+OIdSlNnjFN9CTOvzGRdaA1
FEdCTwdd6IV3YHXGU12xDyt8TqUIUI003kJgq4O97I/ZjhouBTmUIc47pn40
WRQT9ttdkgW4/w8ZLZbg7icDVCvd9BK770vLwDzqN0trVIJtQMAsytkWovA1
S8P2+45c9M+Np58+Mba3TeX6cyO5G7OTTO5+i3rtSAs6ScVWXeH8oovigzcI
8DIC+GlXwL3ZEBLZceASNoViqDlMxlI0GGdgXUCPum7QqIYm8b33txTIcRZK
YAW1hg2mt7vRz06W8bvV9GSRU49ItbAgZSKu2lgACakrObMijHpppYK0+cWU
JRGVyRwtyvzI2S1+jkxQgxEAn2uMlVl5MGDoqO4zBSfubLQ7gEhpg8plB9mH
ywRDq3sHD7fEIZSa1zW9JZVJpsuyN8B59aBG6EPl0OlYiMwXCrugjluGD7w6
vg0CPcWpvByaM+D+KuB9IuUPYkd1PnrGl9xSUveEY+wXGgiPGwEl33iaQGWY
5yPH1+EZUAOzZjaizRzsqwWKHbbHczEdumiMVYti7sPyyXujT33OZWkaTZf5
VWeGQrHuBNm8U4hdxJ9+dajxPP/Kt/9I7otM7acDx+q5MbQMUzVrDEzvOAHg
wAj150B4QWGTlRTtpY97MsyB/GfxIW/BYdf/gP1HuRR136SAEcaTVX5hfms+
kQyrSaiepL/T9hHXY6QFt8Ld9DjAuK2loDDtBbbxTkls4qjrfYXsejIHrHHC
GXOAHFCsGbXfchiLjWSsvj0bcmLusTvkyv/Xlcs/3w3NOe/yjQnl+J9Jrp/S
+G/awzioS5oC+TgHWg7Om3G0BXZixu6h8yk1cJquE0JQqG2mbzEnbqdcw11D
cAsopF3b7W31u3iKB7jJ/4NxyfHlRKxqFvWEPKMiEjWF8dNNLd1aT9DpYhNI
bEZWmFBxjQ8x/iBfBhUmUpuSzsIT3UkF2V8uyFDXzH0zL67GmXAriJIe0+lw
HrZCrPR/U08eMrgu1bsn7kys8XTgveELzhETFWHO5+l7tKEPC9K7KbCapbYS
aiT7VOzRlUomhqY9qdCCPNI42X8qXIRy6kRZYMpZTQxZmPURLINtJRX0Ma62
1YdNa8wEkRN5AkXQGud+iJy6kzly0n0izj1QmbabGdc9gWiVsZVblBkFGrf+
EfBaNZQH4zlq+hg05Xsb8YWywO4API8J+wX0RXtXR1UJX/diFnNdOzpgTQav
YmJup+ZLaTeJMPRHeVQxADf8ySL0Gc+P48VEy3vH7IJbpPvh6NkzkWE/n7yj
PgRcetxYCyJ0orvmA1WmfjeBXeRRqKXhw99eyh++UyrREf5XWb688ltmfShP
g3xmQk6+f9b6w3kqtjxymLAWlsmrOlRdUwf5CQsTMzwkh5TAVB2DnIXJvDJj
QVrxytmNasOq4gzU+lZUghs3gBZYyRxvLMy++jtvUxvsv8dTijUumeF+ciNf
PMsxrroB7WrIAIbTImQlJZ7P6QryLPH7w9f0EpUr21AKv4YlcNMU19TOfXSN
RMfTW1jyN8dBYnKidQWSaFjjyyDIYlsLDefuhRT/pB/gAaLF49PNZ1k4wlIZ
u+El4LlYgsBU2vsCA/Xs3WEgLhM8r00wyM5IL603x9vK3jVdo9fqjvbr3FRe
YCEeGF4gKAm4rugy4H6KedOkizQU89K1/ZJKyVKuPcJ8BEiwuvWqwuutLbtw
hbQGJWqZaCGT2/d7ze3oIjVNeYRyTMJu76QGjnuMFv4GkRfKYfw2B21G8MCt
o607JogMA14GJTyrsiQVKRYi+nsXj3ilpZ4pE6atiCQZY1O2oZdkY0WnWg9U
t/xITIj7yFyG/E8gh0Sr3ISR7Jh339n2TzkQoliw3xSWTVeXPqXhuBHVXjnc
+FmDcNU77D5iC/RaNxabsremkUDxtAIKnx/ex61nCAH9a0sVtGHp7c6df6jZ
bnnwPXOX5utzeJmavDaCdOi6GgRRIjnMM/5myv4exJfGz76w2IOvS6IeCq4o
i/Nkcq9RhT5XW7KcuKrhFQ4HXwv5O84BauBa704I4VRAVt5Ma7wp1mnLxioq
qOfUtb3GK/PIrlDTbMynu0vJWwfjiJNTW91SvZGl+olicHjOhtGLlQ0dtyrz
wUyorkqDdUGvL2JqOI3COJSnIMD1AOYqlkM/L/s8yMu5Mv8QO8jItaEXOhEP
7ARCBmJcBBMWbYVHItWMWv4u/265KR//Ll6K+Tn2mpsp1LCxeUzAMzbCCBha
aF0nwSFy9kLp87oG4XlgsqlZ4hf2+2Wj75G0yvww71vcKEBe95KXtaXXYU5D
8wGU/rubiLpHK6mSGLzyTLj6cCoi7hMLtE79MAu/7A/xd7XlaPPfpBj90zJG
tfROOhRCFmacSK0YKKW88TM/IlG3FUB8KKXWnMqBI3w/QdiKX9+4xFKtmHd9
HcxtUjSHvK792vK38cI9042IzJgKnpViaBoto6rCIsqy/c5Qby4vCXJpPetK
9edtfTzopxaXSrOycH9XJEMxu2hcNOHHF5xAADYcPyVJ/op7o0iGU08rykbT
Qy8LRQFGg0UFV6/O5+ykxunUdmjCbN2czhmp2rTDhqw2Qp1FlmgZzKeq/fm/
TgFltBD38EpseVQaV/+sarSja1AVHtH5qVRLeiUO4h8g3Rlp3epqdDmsFiHR
uJVAOLUtecA/m/zg66MAyDRLWqkngrmORRqsfAvIBadoZB8w9+dwosal5j09
fYgfUbGCRBnKyB9IjfAkuGNGFnRKZxeUqSGvzZVw+zGHjhZv612AqrJ123cA
QBOn6T8sjQhSSehqcceugVRQ+SnGSHjidNhniE3w1YiJo9gg2P4PsrXrLMPb
08oS6UgYrcbwqfGqIenyy7EnralNkvkLWTK3o7EsKPIxqMCBPQ8ggwp6SZoJ
nFCTDMvsZ6OWEigzWPfgP4xG8FGmpq8oLrzkAwVUG6mhUnBPiZAdP2q0CxPx
urLJR5YEKVOOy11OO4G6Kez7h1bsi5iua3yIs6BB88MqfyFcpUpet6ffmzzJ
yV0Nwv73fBiTpgU2wWdzyt0GuQJRHUY0PHN9VsWpoc5KybNltazfb++rpemA
bC7Uh+6jpCJEKQj2dIjgeqs23NwAoUHD5sOk6WqLiYaCj4FAjUcmeSEj/r8v
jW7L1tXWwamae5IfpSnTfL3pxtsVfxPejvexSSM9WZzI3kroRwsjENR/91ai
NA29F3V0gkYMFOGCZ2kSXrR54eHVIlqOGtr3mIcpV2jL1dz1gzd72waMuqvk
jp8/G4wBLgb/E+VCNWyDrvLzgIt6JmRRgHVH7Q7lZ4zfFfkiBKXUVuD8e//h
S5mv7Xumx6KxtJDlK8SBKUYnjUTozAl/ncrIYjC7hLV1G+6NN3Cpeu4FjVaW
c+nY9JYL4zp8SBVpc+oOUJPBqkKcBw5vsHqU0C3YPivG5iwrIq0749HzgCcJ
nCb4DHb/qeIJ5KBV9zQl08tvTMNDx42xOVVEgPtXtG8ruE20EIHa+HLEwo97
wWXkUPnsiooNvHKR/qgv2+fnrjRO/Q/hTvv2AysBhlNUZYbDJZpoBxf3+NXI
t6V8/W/cBLxfBwKv45/q8Bu5f17iOm2/WiZyVtQZKRpBxzSia6WRoo08ZWF2
pw2uWtXixxQQphiH3VHK7J23G5C5yPdiJEkaLQyF0UhBYD8Gm3s0Io5iIu8O
a4gyakP32scXNPVkDsHnG+AA/rI+4c0lylE9cJSEGeYimGD9tQCr/WfAp7Tj
FZytrtOGUHdxRxTXUjVNxRwllU80G5kSVo6fRz7hMdsgJUARr/P2NMoCmTF3
Xdws5QE64s8i/MvhOsdoExP5wR3IfOZvd7RcZr/FJglKZ292DRac/PueSS9W
gxdcy99uNne18PbH6WUGSTeIl4aQ2ZKLR4XSOw/lgZOXeVNIQqjYABRk0xZI
vmmyz7zpEeXx57Clyt+m7w5wTkncJT9ad/FAuIQ+HGKK4WWn0o2DoJWk7uoW
GLFrrx+bcHocanI59FjDOa9HpsV8saE8GjZVA0hWgLX+SAqhGxetAxAZnMLD
3iHqBuPvI8PgNDz8lT5fvpqjUJpFSPlE2zGlFl8lu3nqZcCJlmcsG0+Xim3J
aRjMxzYm05OAZfubo0IFaugkt2sJec4RxFeIwn8kX1UR+11dJC5/ZsZvj/LU
zZqZFM9ue08GcN+Nf3tEm9BvJateivJAISoO627u3uoRYO8vNz6yuzWjBtju
Mad6Ei0qjyzKqPDpiWufgGWqS23IdHbpkzmYAwKS17Isz3F80nfbU9wrntYS
wxx5zLf4r56ugCd3ZutxS4mySfuQOfDcxNIMg97tEfgFGbajROh91oF6SXZ2
9herldGgPapKFGzHvK7IFIF1tX9FJ2ah80n3JjEXPyykiAwwwH/1iJPiUc4W
1l4rfk3ZlWfB2F4BSbMKIgd9nMqo0ss4h4a1Wa3LMYeMsfjAm48doQqt2Hlf
GbF18h6rzcf6evWbCciYDrpXiEN3r1jL6aKLAVYLFqntUsijK+djHlulqLJT
V2poqYWuS0NxB+kLCLMbXFWIJWLgRYR5rcZdKaj8sG+jH57T9fSTW+d/rywA
vQscScHi02AO/pPH5mKuwJYr0l/4VU6rfJoJ2i0vrLrLzP0pX8Oiq3SoWBBY
X9QTeNUIhyLNpd1cvSSDi53+qCKSZeiX2bjkBX6nxxpKLk+ZyGHtO7P4Ae9G
rPy2l8xsWQO8uNBFeXYvnI7UkSghJ9IoillEMYBAo7P8m6XbThSNmtQMEhSg
ylBE3HRbbh8sFAkiLOav8IS451bX76Ip8ZvYGzctAb84MdzxPstTU0Ekyx+9
zmfoi7SqxkJwq9JTlV392BNTDfAcYHH84LJDM26XBnnmZd7MnOnX36yhYkZE
HRRWmjlxaW0yDlrBHQisfEhPpo+hoXDfKfyAFGoMqNMEL6lq4IB1PcP26XjD
rTPJaorqzLvhN5HI10vaBH6j70mxBpem0QkcPcj5N4i0k30skFobP4QtZgWp
Q1yuqOM+pWfablgLKdndMq+UsADQ8ljWk2jHaGr9WdRxC5mSNtC6QYfnIXqP
1XRd2hFlU+mj3CCGQmYEmj4ecpZkrN8tbfhAKwAsO1Jygop3oXWh0TV98yfl
6+D2w/cJQbF6tiTc5Vhp/RWl+92GDNRqBKSejzi0lgi3jAr/A3AP+Qghv3Ex
DJnt1Hl/dRXBJ2atwwLQDTDANXMjcimQL8KKCk8m9vCvlabKOhWAXc4zyo4S
CYl+bmQedkdAma9KX6mYps+mF8D846jxyFBM8ebms6Grt/4e4ciMG8UwM37L
iQGBJGR1wEwwQJ2c5sBGtnGnW49x9By9qjJ84Po5t4QTnSrJJMRzom8MCgu5
f9C9Lee+kJgaGZ7fCx9rrg/hlIoTSB1o1yFQ35AUXGGNHE4Mec2UpQkHvbXD
ijQfkjjchEC0hH/xhHAGaUORpvHEYBz7cWLkmKVmVv3qmL6a0jgpvmzAnPmG
agsim4oRJuOsHgPw6TnIbzh7B32jAAMvmnvFe4c+/rVJRdHvBwzOc0+WPTdh
ejrLWhcNpYXWKiogZsv3awYDH5XxhAJvjXxO++3xfYRpjB0LBZIwcMg0fHRh
1aAn5EXfxQ7/Q6n6f7/bnQJNWhNPSuw1g0Ef5yUF2i9BgNml6L/x7gQnnlb3
RlyWsmNduQE9ufMZbEmGhm8WUyl5u32UIOL2yIMP3DcvRXaSkM5yv/rjcbjM
rEMGLnrnT70kMxMeL3Q2gXWHEfjkk0qq6VQ+kssv/vCslszkrJNF4n7p2rPE
NNB8ORLKhvWOFgRa6tqHnxDcv5GTL3c284aCW7OiejbMBP81ndIll/rrxw0o
S27xb5jbREWqxpHGH63n+sV2uT6KxSnSzLmKscmsJOKSIVxZzFdL/70fH26G
pI+Ij0RIe2F5jFKiZQ394zgOwDYS1j5PHonGAK0zPScN8khvhT9Rd1rMYNwz
5IJzByzKoBntA3WFqBvC16umF2POLkFw5RKLoVKkN2N2ssRSUF7lPs3vubHt
XXYDBBwRo9b9a63u0fzu1g1TWEnR8mHEGFbc6bVOT/G0SRrYO3ytRvr/vJRV
rboSe1hNIPnyuaokh1MJSRgjZxFN0Knu+AbTs43bNTBxowpl9L+pB/A24kyz
wujNA6EkLo5jfzXUzCXh5e02UVbMl3Du1FjuHFWLeIZ5XKQTE+a8xETVt8gr
tw5hXOgYhcQ+pPabhnTTGvsAiWaEEnn4Uh3IC+/NrcZvIHplBneGgvCMPboG
VY2iungos1g1pEf4fGgakP910+2FnBqOvRTnUSzlmqPTKHTtst0vkqnX3WNt
vy9QdGhE4M/Dphc074tMfyTJn6NmHEA26dUF+9xGo2qb7IILjgLViKBK4oot
uLWQcFw/TRiIoQGpKd+Qfh42SNtQvNqhYKrLCU5aGUMep9OXum3uO0THqYiK
amSv0Ur7KXV3kmNXLU7uvjeThWswYkCtKOgwQjvwYedfE+LiiCNLtPWH07Xi
GjkPFpRDB9oREydYPGAs/0Cxm7UqL9Yn4x0zcJQYZugXJwLijEPrabrDf5KO
HALBOv+NP8vG9pCjDlcQY0EBDoxQhV6rrckicHDtcNKv7tcuBXLVxZTzLU7a
H2oX6dNFszzJyKk7hA+i+1PTROwlgRDD0Ki8/uqnRTmKi3Gu2x644qA7KVp/
xPWod/ZGGssTyPUhHNpxbQPcqZ/x3jKtjHhBS5OBFK8ihW17tEXnDE0OCdl5
3XxtWbabN7HMZKFG+b0VNy2UXYQwzYA6z2zkzqbaAPyBk7C7/EJ6c3D0cerk
HsUx+6L/v2SoDEu///Qb9APRN2mVNU9HKFlu+EapOzBQLn+mDzin3CzpoUGH
BacHGGhLMAHPSotcWBxSzuVmSp/Cq9jtUTUH0QgsXwqYxrkb2lLZFSzIrGBH
IA6NnN4vfvnbpr6LI1NL7jxnlxEcteHmsGw83V6tRTyA9gcDdyuSwLrc6KbV
hjIhHswF/1vkadI2K+wGHRBYKlCMyafQDrvJ0fA5m8v0zi6jPYl2TSxxlPN9
8CQLIN+fL/Ys2R8w/aRrYI4fI/WAf+lMstzal78GvMtwowhZIediohjs4Pep
FRC2iNE7N1fNXrq5yq4haFADToPE8PwIVM2CRkZv61ffgxsERA/SbRZ7Y3ie
nXBuOEvCyOKmcGBZdbEXcekAdJusDyzxHA9O+KKKsFfGckItPyDPIp10fa/0
GTJZT9rhJpL+Thg4mX6pEIOf7P6lmHGVOuA6EXZECNvAj7HNrnNG9jY+oLht
dMOkeqwl8GBT3m7ihz1qByjFWNskQdBio+PLcVPkMSfjEVE82OIA8a0YJkXr
H9foOPNycdmWhk1/17g6L8qZrqgLRPlKdHttodjOeg3JBIKdvZ2AwLgdK6LJ
NVx3zUiEoN++aZ5K5Fio/csFr12n4YDmioUJ5PZYr5zfptG94jQi8JijL5tk
QE1AC2cJRDlnIuBCf3GNaP3cATTpQSdhC8bW5646hXwRh5xckiz63by7obaX
Mw0coRZW9HNCBbdZ9IP5mOseaA6WrWj2Vl4PA7EgBefPDNYBbLLkIVqMZoI4
WVKcrrzYNPxQ5ApTQGVPxOwqqET2qT0oHDL3OVrsI2xeHGzqMLayUgQQGN+l
3oL329Pzy30ickUxY7umE9PwTxQfXE6akyGNq6zsGzL0OvfUoAR+hGsnFVks
361w7jjbDrWgxFQjixVW1NL0B2sdbkUURylc+TxF0C8hkdzzSxcoKRs/+1ye
FIHbWVUnVpFWe2qSkaQaMcb9hDuZ029HCxDIIcTgc+ERMPBOqjEGbgIsRHFM
LLKNcNcF7aI4Z2VuW+FJXVxl+YnAk2fbQUNRmn7gfvoQ9HViX5g11qE2OfkH
NtdodXXbnoIvYF+64lYNauVTqYGFLZW9RY+eY5+DFfA7w0WMEZ1GJMoefs/G
vSrZZFcB+lf9juphuSjvh7nLdBpEh+B79gtxa90Pdg23iAB+fIKbmlJdElxJ
vb9RHXuLTm3No64uYpBm+INFIwafbacQLZmrSSvGUwajkpyAbF2VTtShh092
HA6bLiUvFwG61LdgGFUDQ7r+JbqK72KJLLnW7xY4wnOZ8NfhEoCvIhTNLrSv
BfIMIXVW2VpfK7OHY4gT7v90/3hzOhw9qZaG6rOhLc6x+5XOZoReFUHyM2fX
0cpQ9+9yDfe9JR9n5riFKYyuvPiHAkt59wYEv7TqoFXbOxqjxpLuZYyyUiaw
ewTYE8MS/ApKiN0yCecu2RJVneh6piDfj5J5wE0f5Vg8FIKqyhd5h4cPeets
2IlbuTeD7WzmNkgKlOr+8OxGAbZXtifGFgMwH0UOBrgIsbbAHJBfk6VgZKX/
FPJgM2wZKutACQWTDXyGBRAe4BW6w0jp2kTrTxwlDuVNhTOHnBw+YV1d9skg
St2y2YkCfkiPu4TWjzlGKtHH6jYJdjZWIoxDZXteehAENkGI0Lb7XVw3zYgG
k7MHBaSr7LLSBGxLrbPbRNfODMqPVfpcJeVCPcPrdDdQghKlZemI+YPxKsvL
wP7EjCnIZcFplb6KOLZn2N3iGFvc7zlVpM1Li4uNP2z61+W5VhQN33YjkFpQ
bJJ69CibMW5MswKc6vr30dG2NwXrdrTCOKEZE6OFjiY6t62bwcdr2Y1GWD8E
tFP2DVC3ZunfP1cOeucccm4PKZJ4mPytYl2phWfnCwrEA16j0mKR2gd9eo3y
idh7X39ru8EQLaJ2/FxyUm6hsE07rCvCIc+tEwMeYueS7SCepNXaku+XsFke
qnE108xLfz2JwwGxz44WA/H+BZiHHpyrKlAtNnAM7Qoc98+uB4X7/0OglZLt
m/KEgeKc7qlgyoG1NBnJmsOlE6XY0PAaRQRDhVR85W4j0gB14re2NsXMHTZi
yHTHQqh/0RFBqvDj+H6Sboek/DM6lHhMlHD5V7eBNnmVTQfW36mV+OoKFC9C
auaa/Wf67B0oa5Nag9tjw7MgsMG/6oA8LYPOxJPZ+l1OFB9tBUa7qRS/34pQ
KEujY1iBJw3WhGFTuTVy7dIzgAG0ugYmdcFZWb5Y3xRNK9Hu8fF3FUVJTqAj
8QnpdmnUwgKzAO+Qj/2uexhlen4HxHTSWHOGWcvsDP02m3QviJPFZDbnbIrC
Fc+xeUhLrvgZa1Nfvx1EUTRhmzulf/bKQOcjQ3xpyobOaWd3bQ60Qx/buH3n
IdODW98QaFi36ZE1XkRqRyOgUutsHcIkLTFXg8OhnhwPvVgz6USicpRKvg0X
wMvwyesyp7jtd14u4hpgx978BdY9gHrz0XZpYPqDNpI42qH6n0LIy4Xme4L4
p/Yj8TLql2vX/5oVvnv2Vz5yanEHOt5x0oorpcuvLA1lBXqH/V33skLYZK6s
guptpST4ICjRCZ8dLeORExnlq/cZK9YtU8sOTsh9okKQLeYgpzcudfrIDLDm
trpsPG0Npkg7CS3rJFTg7PSvEomgX8Pqj9p8asXCTIyTqfju6aY6WiIJycAS
huKJweZz0YSyjsSCEWPLYSDpJnO4Xe9Xj/1wvZ4UYjqPGquB1zs4ungerRwA
xbD8zOsmtsFTqyyWaqX5LdBM3pO0UAGShvAsG53+Ahm8sivAiuxJC8IgXLuZ
vd8Rd+dCymQbrrLZ23+Fp7Wa31Nkuy6dBc1pyhIl9bOXSV+ITSb0UyYYAqJ8
yj3wBrGTVuUd57JXdxT12MxQ8dspHEP0+fJ/TcyEv+oZzNNj//jehgkl5SR5
K76BUYp4U1wwwLRuD8q5pEsS+8mdPZguMCKftRCND+ZgVVV0G8ZElEGXCvEB
/TKImFrNy5juQXQi9vtSwzVYmi2qnHMEh9758E1JHRrz9DsdVixxgTBsVvjc
pMDjxCdunA+LqiPz/pBWJmN5NP0oScMIb70+893IygndNEuykXH239HtFQM1
GJPODD1quizGv2lpT6WUf+v6QiUDS8ZgnwHWtBUp+HigpAiLQ+ARrrA0cv8t
JT5MbH4en10fBaGsa0dAqY3qKBYmOOcA+CojkwCcae4nMFDaEQRmGkXCKHZk
ZAvsueAJNoej82N/hZJSD8PKrzgEdsN8Mqm5oIMZ6iYJj2Tq6J4kr3/klyMF
/pekk0Jn3DQ8Yvm6FgvI8eGrbaLlXxoJhI6wGG02tSADi1V5Jkg58A7A2ptO
2LyjIXnvE+NTQw8sVdPGy7hvmreS15J/rQmhexHkpIWtY/9FGFKhaMCApRpO
bvKreu5UT1SPXTfWNEwqkUIab8bE/gtBIRw3Ur7wuGv6ANLj0nTixDKvG5bg
8NnFFIQ92giGnG1ACK/eyVNTMaHgHCIDhRi2Y8LiADgr5qMJeC+HRozN7oLc
u1VQP0G+7aHPTa2ITCJynYWS9ZIxgTZzAT0oqwDx0u28oDbzMITNrDaHAGv/
ObVyZaoVeBgZZtft8L60BY4pi+y0xv+iPWQJ9/ApviSCZZCHAMg6OI7lRMJE
5YbSj6wqjQCEBvAw7h6e/8BbuzHjYPswXGizc4xHItGClzInZb3wMhUfKKT1
PjG1xR0wu6pheeMV8lstM0ebp7zftYQTbpNen1J8hOzzhNZeJY+9x7rEmocb
ugHKTb6eq6zaTlDeAJ93WbTW6nXyywAj3f3hUfOmWLGRSGsVewUzcPE82VVl
CXF0TU+x4p2AE87gwh192nWfHYoYnqmBYd1Bzn/Knr6bFs+7a/MAHbXRXaCQ
8FMALfHvTQphCqDZ+yMd2Ru8ZUJTPwLHle2HiFW2QvPLiwkw1V3MBp+Qr4nX
I0vmGbz+DCNPqraSfi3s5/btJloq1ZKdCVmr8xFbwLYjtsXQyt0Ocx5XgNVv
1hmM68cAQliQ3g7oAgffQM3hVvJ90E+/tNhGSUrUMxpf+GHtL9xpQudBhgUe
G8qPkSJdBndqUxuxJUSwDp0P5I00oejBGpGltkwCNVtYAbA5tXG+3O9xq2sS
s9ONI52HvvPdFbo34Ar7lkN7pRYWNTEXijLverFZd4cW13EAQThV7UoNZCQJ
LhIO7cQLl3Bamolcm95La9zKTVR1fcWwEcgk6EYnZoF8KEwZrrODxatmjvWo
ojWXx3q1xeHRS6KSi6UuE7GOO3MQhlizUmtSdBZ8IcPAs5B/sIviQtijaKhg
Q+HxFtQzmmASx7zN60003ocZLuDZh4OhDuriKsi2rjzAruBbfTIPFQLqp/LU
Av47wb2vfBRb7N7emo2Subh5yW8bCdZx/fAA9XB0AhdrcGWz215H6G3/t1Th
1ZP/yqWO3LmOkBtBPhtwjcuHBmC3e1or5225m8zOLNx4tMRAk42uYLYaxb2u
exwD+jgGH8fHhROFLTYhyTMy538vCLlFCPYTuRvJ8QXmUMBKWEuBVBM3TPXH
4V1yfGsiS/VK7CzbQR3slYp8IWDQeyK/B/HnB/6j3w6yxhe7pOd/1ZuAj7qW
vfjbYOaK/LgbnmDI4SsokZXeXBt3qSl8f9TklU1QLpCnY5AeNCoQOzkphnhy
0sTdJ1CgWFlmwgqVPdLVjyfzQUmaqsqIPIb4GsLdVv+x26r0naddeVHaMoum
Myyakj8w666Jde5UpRUBdnZyAGpIQUgHqtDdXNlBSNgk3TFDYYO0US8JRUKu
BYRFlgzyK3g8m/nVrJ0ZN2rVNyOJAAm22+iw40pbLydYFTp/I8FA+pZR1wlD
AKPNJaAShZ9dWtsu53QQRh8XulWORwB7W7rhMbTK64/jzRh9tAIqfr6QKEUn
KPfj4Icy4LFwZsyw30uy3afXt0QWuVNe5TWmBN3J5VTmWsvRoyrlSy16cKwC
3KFtM5tXYmtDRSF0TuOXWhBDcHuP0tjZFN8+D3rLsVMrQJXz8pKJ/sOox7A9
ebgp85GK2VxVc2JP0ZssinJhinljyIq+Adl6AsJscPqaOBsbgwLuikbr7cMN
FNZ4T4qcW2C0xUGeZOYkmkt/NbimnZgoNN6rg7XMhnj/XNH1sPuOzRiTNr4B
fShhyJTC4Os/Y3/U+9HirGrtJ4hRArP8aiWipV5RqQ2eOTyK2+VTBHVLL3fY
gZ7HZryJrT1GZtNy8phHtO7SueKExAMR2Bo82Tv0BVyCNFlhLlscCRto3RQk
67Saxw8YZes4ADMAFxnNMW5jZV2tqH8kt7JgANe60PfExoExAMopD7pnGpt1
Z7OiBe3TLuiqcMEgcjKqIffmfMda+BUrQO2evY4deiJAO4uZRxgSE5IN/E19
v4cQ0oswYxUhhrBsAW4avO042IGBjGkt1SXPdE8B7z/4TVemK7HWvTRlVNut
eNMVLW7oKn7I1FxxqDCuNXmtwbIQLjOeHHyeW67v3W/nRfThigZP2zSURas1
3MXQU68MS4uFd/5IpYaH4ydXyuaRR9bEHWtjDsBlqkMueCm5R2GHy/ZgQXQD
HmIKaghtdPfxDCzOkmLAkBO1wSiH+2QmFsZwWagafKLuux3w7zm13HaS+3R0
ik6mQsGcokNJIb4ixFHd415BBgv9ICU7yiCddFlLYrUXJCQ2U3bxLNueY7kg
8mCbPY/HS5p3FfFeei0txAtgOQaYrb8Qfu+VNi6T6ExOf/xf43tNYYb+kPEY
+9guA2l+biuxXHl8NgYWvuICoH6hGKRoGgF3YaK+Mu1YpFV3JtP5WdM73x9Y
k8zOqXQuNkDJibDzDNDmtdmitXbhul8wHvJFeweHvv9CoosoWHMLvt8DXshV
+tCY3+7nYir3sllK5HMn0ncZ7lFltwT3euXIHEYiHae7l/dKRUXDcIRXuqxL
n3d/GZaym95DvEt2gHeFbAHwQdHrfWln0UOuf2zkwcrX40cFvYB8X/75f6Xv
GdeFE7nVbE2y4N2qZYSrJY5ZF4gXX5zQV8eDXpH5ppZiZ9GQuhIHXT4sCpUj
5L2Xn/yhUr4Le/xbAtNu8XsVRkM6Kq4GDpVE2IkmoKUEiPH83TTXJNw53zEe
FEGWS55kkeLJMkBddmTas1ODWoQG4CbYr+r9OEdIsA1l6lnvx5Iww/7WMcYD
9X8yVpmetyJhUZaxQlsN0XcUIKtpHhx/jSUdxwW8o1B9fL4ELhUJiFY3JkZF
aYVSsims0k+X9/jafzXnpl8Vh3foOd8xClzP5oApyt2hfzjm53JC+eo5FiWu
QpC93KICu0XmkBXI9Xw8cwlYpTHrdV9WafxIHXw3nLZXRlv7Uu8lTPxl6Lyy
lGHq0L+wUgTsWZcvaw9/bkuuiUX+Opz+hvaGyHR1lE4w0L+N+wo/X3JxJp5A
UYL03aVZ3q3HLsGLsOEB1jlRDJrgUTvTL+04Gst5jHZzZbIBQyDrMZaj7QOA
T4Pko+a8SpMZSVaP+RUmKdrCDw3KoUpLVJwymKsL+Ltfj3bhlwu0RvxEpuLK
hIHwk+OiD+A04Pd+/C3QCBUMhkT62JciJbwE2hJxLWbMI3K6xkr1PNUcN3wh
yZChhPXE0ZIzHYh6ij/Sc9KOEvhgDn5nd1Uj5pQ+64weRVwvAniCRTdCmVtx
/DLUKVNngP5LtupvXg4N0hcJpQtgInZFln3OsgNB7ViXumM/XlDrpyOt9YSL
Cjkz1U7/q/KQUxpKAkaCmeaoQdMtKINeKThNHHreJo22TVg7AZEP0XgZLhJF
JZKyImZTStzS0OF0v3GHKWayP8GN1/cLqnnpX4W1GF+je0PWCKuLiaRCaQSx
MZsja7bdBRRnn7piZydCEmPAPaSHMOWbO2ittrTNXzBnUUTw2gRqdQVNL46R
N+Up+0Jgn2E5ZSxpJe43rbHG3lEEIEm4t4TxVpvbpF+umgUa9OUT5e9iwLg/
CPNpY0zb1dgs94yNlAOKp05gCiktzxTHlZEoGksLi6O8oe+QMwAneu42H5Ex
MmbUxEwrpzz16s4yQg9OA8PmkrvrE82Ferjshz8kZb5D+pt4un3c9k4+Pf4d
/EvkOvFzkUtaLfVkAeyjk2WGWOvfTy3Llt1rPOixRcqIc3xNbUkmAJguKjSr
HiIv1+nEoSN0le9X8z2oAlvZGqHZ/OcYfG3I1nL/kNClu/+RTpeuxdZVMxMc
PfMrOHrw2Ay1xdHTXP+efzpI6x2qMS7o0Kg6yONngKNHM7An50vosSRS6Q9S
s3fVyM539pK3+Zos/MrYxqSN+SebLJRvPNpW1jwwmbO1o0qm5CUvysbRV4Hn
+eSjzgMV6XqHr+rXzyek69OoMsOTm/g2jNy6U/0OLg1H9eyGhQrDRvP2db7t
hLVqCCOds26XvRfHXn73T5NfCqQ6wmJXIKDyC6F6W8HmfrqABxqGXXvf+FVj
7WSVx9J672N/lX6TRaagWueio9tsAYWAizs77Z2amiOM95Gi5ArmX8SFHDXk
Y9Ud/mfADvH8z5DJ/B4sA3SpSM2bShcMWTYj06TuG0FlgjSqVYKJCm75OInK
8WJ1zu4Zqb1db0gm1AKFmFOhGOSo797RN7XuVJsJHYQk8sF7NDCRjChs45XR
PjReaq6Zn5tXEv34QR113r1Sjp2Rn0iOTgAqqi0L4Yp+qjsNzTzSbOVjbVtM
Sx/ylM4+ZUO8FFV53Qc84jOfXX37mj/ihq3fBv6esHh7SW9CfrU3ppgV+eDp
Mz92ggwN2WylS3ZfPtkpHGPLRse4LVdRcMeFe3Dfrpv6ZcqTgf4nKTcl0xoI
oaOCRf57AeBPHtWsYFOixODlh7b6h0taY2pW12wGS4LNSoKgISYyEcpDY6+7
gwx6t6AcwCzutd98lOMdk1Sih/V6fQ4Ww0/qzYRwpkvabtMh14E6o0qtiulC
Bq+Eidq8Wwk9FhRqZo/9hwbh6eCtdVbIVaY8EIroBIXlLas/iBI+g1Mc0jm0
fYMMELj+uUYy7Q2Q3BoD/iPpySSleEm1+FWFgrSupJx3IxaHyHhGpRwXzi6K
Fa1+DaX9jAj4zgZahQHv41sU74OkBcaKlCFOH1yCYZMSWUdQ2Lq0Y8ktbeBp
Qn7ejtxR5+jhPhZIIulvkxJHtHQ57/2SLLekRmpxGcFOgfoGCRIohJOYuAvS
pKNjqb6BoNlPlrHcGZ4TZ+8f13bC8GWy/D1QnfA0HMrEZctjI+B+FZxLkN/E
Ot1I0TGCBB4jKH2dGNPuJjcm71rZ7hNlHzdB5c99MnUBUFigQz3NtomiyQBZ
v41YpAakg78WVkVTVTsQpjFVpxhZfRdu1cdO8R5TOqVflmArjGpJo7l5h+Tt
aNEOYaitkqTZ+RL1Mn+6v73Uju6wYhDufcnvTLAZ/KB6IlxmqjsKaC9qY1Sj
EWCpRpmxZp2cnG6LexF+n2X5rlyQ2Qhqttz6CvSL32YkM/2vQhL5rQiM8rSl
rVoD+rTc95BM6H/omqQV39mI3jZmz+VXLlrR4ced68paXmNT8bFmSluNgyjA
kFNlCIO6CPvbJAKKshejpA890lz+gLbKSNLWKrdcw3G8kgTWKA/V8ovxjGW1
OCKVgCa5O1+iCXAx7pJMpJc7n8Px+dL3DxAoERox2YSKpxpVGfvW0CZGca6b
1jd1diCsyg1FsymOC6I2yCzr/A+jflAJPvIXTbrYvB/djmrGFNbHBTFgYcYw
oKYppjOYPSn2AM+fTPKWrOX+o9Oq5ITJnv9DGFNaABG06u/11vet0GZW7Qb/
K5t0oF9auyh1Td5viBO4TFNeuYbaX20ueYc4+/JXB60a01NUVuwlBaV9xH5z
k8qEJ7StYUFAKALQSPi/PyLY7onkqIOO23Q6ikICVKEPP88pFFiPnMu1PpS+
NFk4jKPo2rUNPF7JLtMTgMGM2MT8FOpS96icGocvg0sIMvgccAI4HO6Ei9Ti
9oAz8Ol9x7wcU++lJ1YYRjfImwvHumh1Y4ZVFTxRFkXqGmfqTovHYz8tlmra
68E11uOQ486j/TaJUrLCmhAsHftcXREetl5CPOwe0Qqk/YEWJjhuKOIeHiFV
dY7iiM7wM6+RZvRyYWmGZ5Se17wJuCBMP04AnIPTgffYrrJBDNmLqxTqj46T
vwqac5DcdqR0ii+9l7QX8qaA3YhS0qZWWQAYjRYjlBSSbg+KRrJkVmHQDjAS
jbC6KnJLd5BwlZ35trtMnc74NJ1t+t2WEA9BzJ6SW4iqls2RJ7AzBPunL4L3
OkAk5mB+WuhD8FWVJawK+THTm5qinxfWHjgKhzNzUfYXmafQyo5EeUnRSijt
htgXLZBhWAhOlm240/cNMp13yoZQHD1wCWc7NMK+f9yEUQWYXfWFN0b2rR3o
ECknrNPDdXuot5d8ASQmayKMNAAUvxQi2powoxdy7leb5bNmYgXM7yMBO/E2
b5fU1+s1k4odPD8hwxMLsvvRb+KIUeXGBs6iERwb1B3eD381iY+1aT4K4GON
uz/e+o9h9LPDCNRoueyt0vnJJLT1cTV4m47oSMFQf08BeWpG+qmjhAN18wMf
HSgY+gLEvcXJ6xcmEdDfD5Lp8RADfhAVELjUXswOTM+p/b4a9GO4PQc1cQUM
oVIR1xpCpwqwsCfGvqZxRnncmZtPSHi049grLnHQ7EBW16bxlp9beT8TjX3J
+B4zjlG7wV9jcaQX5cz8zC0RTP4PwvSxvbbPCfZ/C3VEFWblQ2B3NzG7HRJB
KN5IrP1zUGY73lUU6J2Jb9KRXl5ahf0XI33CZigixltRRotw+Ccg9Pfi9zMZ
htWr/h8ANMtJYMpe0iN9Z7iSHWL1BW/9tVg1bBSTDNixKLQ3PGAbigmyjcWI
qnu/4t1n7nw3OooKzzF9lSzqb6TxxtvI52I57lGdZudzCI54rrMSUG4OH663
VObkTxqTVgqbMAfBu4GdYdjFBBgpGJE8/n3/l7iuEwt/+jkH4rfo/RM1YLRk
g5Ezz3we7SI4nuh2HBS6JwcG/KjdxzNqesVutOVe1HAjYCvcHWP4LvsxeiRh
poxFwnL0x7OgexwBqosjtgmc1c06eg9JVf60WCrAegBL7SAazQCaOv3AxEeN
xtdkOiGngz/0fZhIeuwKM8mR24r3D4CmcnRmMPEhMYPruNSqSWrWglNuOP8f
b4T+GV/h32l6cuLB/iuj5a6nFG+ZlAfyyDbLweAYpbIAqmqAzBglSspF3hrb
brmOqDq9Renb13WhVVG1g2/CDbIBfia0koKs5852F++7OOsXOe5rcaUUZML7
8qUeJSQbPRDvXuW3oQs76KqEIYdPUpWUEu0UVh2ITPEApx2/9o2AX3TdiXHo
PQYweE2qhxsMV4ndJJZQSe4NvdA6oqHceKIrMkk6Wo1aBNAVG/mPdTdD3GnA
zAISXuopZjxT5la1f9QsTCB3XIY5jKw09NAQShafKXYC01ZToaGyco3oX284
VkhdNZyAYsSVfavUIRHwk/g9wPJG8CjFxk3f0P+uw0UMRYT3ALTSBz9DuLWD
PTPxiyFwiiPY+41r1+Q7cfsA8eIBPT04L8tEjNr4LaW3yrB5wYhz7/3dWf+U
7/Ilv1YSycfrUh7KBFpJjrhDyhGenfrUDLUKht/5iWhxDl7coQBm74gdzlyG
XyrFFRomkMzdMydGEb0Uq+uePps84OK3mhHOWnbWCfW7wXeAYQGbrXtOA/Gk
1Ww3dP+hQvO0kfenUTowLWrmros5H26880ppPCX39ffnhcTEE6xo7IKfaD//
CVhuomrz9PoshWJgWTYH2df5UEEWFpOXANd9xL/NRocc4ejqebDxVQEUeoMN
1G3wxHjwxnVXgNZlqo+bXPcMxfWzCStG13Gt5XYnKSUYLKE9UI+4RHlzCd4D
FAahgJnNZF6Ln5qTrqoqZ7kE0D/GnI7r693i2IWzP9FF1vhs/kdGh4pzfAcG
UZmpQZ+Bm3i71qoeFSeL7rHTQGEABRwhX3O5qv+g/DaARdmrMfdnf9FyOvwp
va4to3VSbu41MzRxbnRZW+jfpeGR65wz6FQtREqSVRc42rsm1IRZhMgJADEB
M4o+pJzS1/SJtHxLdOoXwMfieaePbNube2gVxc9V5efSvNeklIgIcAvngazb
rLmh/94a86aPRE5oEgXnHGoTvIyAJ0NblVu+M/Qo40YYRC+Wwzg6JUwpsBsi
iF8B0R23e0dO1RN26enk7lBRG0wtFFZtrF3m9EAcmUlebMzGBaIDSjbAu7S6
+2FVgf2jTS+ro6I9GA4ntlr71EAYYfj9BbpeNQc8NCNKPK1LhXKK0prfkxMq
4V2H54EHra/+TgzntFzWvj1RHU6rx1xGkGFduZpHAmr4tkTxkgn+zdQYb5ej
tUrKBPuoyZ8d8x6zszOETlYGQQGCHOUvzWeWhl8VXhX9FnD9qfVKek71TEDx
zD0eNinWkvTTpEHKWInygSed2SZ3f0oEjPaWxfas8BymfWLbKQmLV+aL4JgG
Df8zOVqRrc2f4EcEjfds64qIVUwob2Yj+28IOP12fKtcYbnjB8DOTSx9OPyK
wIPdpiYVRT9OfE2E36P4dSKo7LmoiEHD5tHxfVdJB5EgITElGYevlZYXUPwL
CVC9320a+WXJpOhwtGLHcc8+ljE8VKPSQMTcey4iFYZ6i386vmO3CvyAPf5o
LKn/dw7ceFnlU9joAxmXS6aWbBVnMNTV7EI+BBZ6gE2t2HJR5im62iAUOdDM
xonKQ5EhnhAl/VnoWpoUaF2NGPcPWR1AgLKArhXg9HhGk2YejfazDHY/kAmm
vtPnSz5YSztE77GxSx5+i7+EDaKbRoRmwZgCZgty44qqwPQ3WsKlC3lBtAFg
uv4SIpGEz/r72SEcLWqOnpx+otMxJfKQWVNICBwd5SKhYrWfGNdKB+gvjy0Q
Fg1rREEcxTAVbbheRABFopfQa5CJf2EExXHBmDzb8DadFFfZBUZLL7Nsqhgo
4kRKApKMkAWL2AdnrWciQXeA2dKpvq0S1Ymvh8tde7WVrbjW7L6/ncFtUwIq
lqNufo432lzDKAJTtZVlkn7jS/pNch3OHch/GrfUmQGZr3/YMZQN8zJomGkN
Z86NOg+n5cc5kqUSpYauZB8+voVIcEqdFuoNHOC+QpeXDtwyuh59RZ1KBJMw
45UmYtjP/hF6M6A79eZlsWw5XwHL0lcWTo7Jqoepy+UcFnF4oxzAdID7Mb6A
Yrbz4ppRoVbXm1gGbzd36tvAlchEvPzIdVQyMWyLqGPYrwXKl5iZz1gAp24I
CTninMRGEzhE5ul9h3sXt+iuFxbhywnf+UF95olNf1bq6Z6AzQsK3ALlXsS2
kSwGAqv5UH50KWB2E8efsvRBv7P8U+AMeqQ9bhJ8moxEMOx7qjA/iU/hgGYz
OMTIiFmiDvwLeaPoJnBsGC1HgEJIC5uwjTDMd0df89Qmu/1iraB5cy2xUwZD
WNmaVrkIeJHoU/KsdKc/KBEJrXMcx/WQUSytSSGZVi8i0CSyuCFgelvOOT0K
CviPzXkf8XiZjhCb5QerBNQqlM+U3dU6FksoSbn2L3ZB0qXtulUVbykWeTix
/CTtm06UJy+e9JwX24wF8i+alQguQcH7gZYmkadMBTvhuNBwwBtuI2O0yPh4
PIMtRPAjPs4RXuisHM3OBv6Ngqznxe7oEueSEZFy9cyeMVnHwgqnyiZWCMC+
WCVhXkkdA0b9xRS1uFh1xKO7cm3I8iOqBpWFdwfTj5dv38qdRXeUhZElw1fl
P3YOf3k4+Qh21DyEn880UZBhyM1f4BpE9/xKQvSSuJmEKbYFb05mnLCjqxc9
5q56Nru9XErG8Ye0vdawYCjTN87sXsyLsQ4jEyAJCHkEfhHUWkIoIZy4Ha+k
3rOU3TpTMgvas95Jrh5Mf8cbpCMaVPk7TEk8a4BH6gOx5GqTcfktK9CXgOO4
Yl3MN23OqY0hmSHgLPnUjrHhsddENwGctJkLk+VO6etAJJ81w2giBwTbqdje
d4/3DkkBVN9Ej4dHxgHVw5XEQs5NPMWCqyEhAbeB+jl7FSz0miak4h+3OUNI
AF+6tBoy3IuPzKNFwRmz3oEIhEpRwZHjMFotR9Y8Lrh63ogvkcNsUorxxipm
XrxZpVd7D61d1Ympwb4L6i0LyEXjTyQmKNQ4fnVrOuz3Cb9lsU/MeCfo+zvC
HOPf3wAlEJ6L3TrX6ndUUF9rUXKC95BNcztDVEshlQvQFEoDSLR/Vrg9dWov
zTpjJOsCa+nl0sxag+U/WdjUuSUvqa2OcEBVgVcW/HFlBN0JTHhrSH0v+AE+
2BOZB4SoVAMwKLTmrwOrbEiJ6eh26YqZLyNnwAo5XpBpgPhzPcCumo3RnWHw
2Itum+ko0jFBibwH0zdoEYswa3YDqR3sbTFp9vZ+cA9UAuGN4FlsyPv8oWgD
Cst3szOmfSPJyYNfTOXo5l6StCpxmhwzUs5zSbKkN8AiTHTI/7R1YuMhBZHX
hUQqsrv8cadfS083kv28GMG3pXSFfzI4gdMu7+mU9Ab+EO5lUSIZXAEQvcJ2
rVCpc/gp+N1pgJ6UDTsrMxtpPVbJY5Hrr2dWtRPu3QDRb0fiXi/NaoeU+mlT
L5jE9Pd25OhFgZ0qquMnzZaQ9jirbh2XjjjlMG8CGvu6W64EbtZCJ28bMlQV
HZR7x3E0eQ3aM3udJO9zHFvn/LIuDHbXqaAVrHF3i39EJMs6CxF8PxAav+F/
Vul8oBwZh7F+RxjfTg6cjjlNjPFi1Z1jY2h8slUm9cD40GEMyAQegTEwSaeC
mwQ/IMcfCnbxUzEKslXs6GPXyhILg9VLZ8mJsURA5YL4Uoe3J1I+XJaboWle
Tzx7AuJQLyBPWYkZu1IGvN1KZsuJ9cGTK+FNpOYRyNQELs7oOcCqmtZDMQQH
ehYJ2i4wPqvrM9UeWQmYfguCqWNORv1tVKgjTFryR73eFUob4kXVp9ZgPS4n
lET1ScT5XhMjHEFEQyayXIGborzkXBXvdC8dhRaCKMezZgiFXJ49MibufDRT
hS2T0P3KkCRJ40+U1L7IqEJEMHFTSaIYx0lP7Dh3ycjGkPvu+n6F199ou4Pq
LkdGvmtJLQ3fyKdJw3KBOYI7X01CtU4WlGKqIIdDJOFnz9esIF52U+aXLzpP
efgshH2gFoDCubbYx7QYN4GRiBmaNTH17P/xjw80jcGD97z5Ah+KQV9Ha/W5
0p00p6FKM75yfRUBtH3SljvQkfR0IIDsiPl+nqAtJiUuZ8S4S3CZ4bibrA8I
FL3odKybLYfVaPd3aF1nXPIkxPWe4+cD0MqYoLunwIhDgtG4IjOxVw4wnbz0
CJvs/0rIaA9NqD+T/SpcjZdnJMXogEMgLc60w/C/T/E7mSZwAbpGdTyRGdbw
R28uFGihEc/gFr2BrCH1kWT9oHSQrY/tbwrAvUAP/qLndyyYLxmAvRFZ+IgC
XLNv15jjeP7LWAfLCiqhM76pSu0gPG6szjPv/8nH2rGYItLFWHyTneGifq98
d9xN/51kDHiQYOnYyZimV3O/VQYowKw8VNDFeL4p0lzkm5bZekPupvyiSyVz
X+03VaWx8RNV/uZ4qfpwyaeMtCJZVRW6buhgVE4LAb5vi2mMMw/SUPwACWgO
C/8rI3Tn1jhv7e0O+01GpoYbWBhW410LAW4P1t5SjlWnDmRXhOW6s2ql8jQQ
kOV6e4ZmWGmcWQZScXiYUuYCHu5UPSrZTfBqY8xVPy9eIQ6jhStSiAXAwp8u
hmZfTsEJlW9ORHiXeLwm1Zu0v1EogbNV7wk15AL65hamwH/b2iSwxTJeFW36
MDiU3KplxrZSx+817I6ycobmdcVM/AdQIeHlXVZGEevKFGuokjj7PUW80dSI
pE+YTv8ehNMulLLaLLV9QSviswHQZ88rVvIIziyuAsnvvm00VAr+Oz8kenJe
AVC2kk/LTwFbPPPa3ZEwU156n4Is9KosEOQK/s8QqLsUgPj9HTs6m7r8Iare
craq6EuRNOoPchm3iAMkBxHvWj1tzF8S8Qog35C23WSZx7QUFgZpPTdfy/hZ
/Yb8d0eU6ZRIw1iNmcEIxPrDBu1nI5qEg2FPaE1ogwCjxIcE0NsdE+Gbqojv
5rwENjoqQK3pwY10WRSqbbUHum9T08Hhpto+0aQNl4qKTmX5nIjVXBmu9+XW
vMyCfRHBolI4V29Z/m6F7xyujinA/JtETEKc9HvgdnaYXhlRtFF/8VgE6jXM
35KlRMna1blBxIIGPPAqeUE4BpJfX+D+KDSen950bvKDl/xChZaWo2rK0MVb
lg90vLzs/A2PblQCVMXm4bOLpPmWlV1nrg0v6oct9UeBwZG3HtgQ1kWURZ4u
uoMzytEwNMrC9+xRm0RHPHs3nowexc87WRTzkRZ7/7V6j8JxrDFhyHuH5MAp
uG6txJTTA/F1CQmYY/EDHlribS3dzqekKYyYFX7yrnrU/W5XE03P7p5GcBzd
T0gUeWitbnFm1oxgIxWD41xlxPIzoXCqNXzAt12VOAwGHU6AF9dTTxs96pFY
c4uQOQtdh9faKWk6nDPawfiCzcmbddhaMmo7ESn27PbfaHI6/vDMDP9yvNdi
cKus7cmkqs0lT1oXThD8eDoI8+Wl/3WtOeq31TMc/sp3UWquyjMoQXKKt7E1
jvGkwr6Y+YsJTrMig6VgcNj8kCIzkiNqXUOHV2w28lRA61Xur10+HZOw3xLB
OG/DYQ5DcQtZvcFxxOZX72e7WTI6wOutmNnicljd53xpJT1/sNgAgbAGsalV
6FL2ZsBeLbU6MOFxOccvYatpPrLGH8KkHhtVydzRKutIiCqp8ZCXkSn4rYSI
yF+kmk76pwJSE58kpTOuo2+SZhRMbOc+Lj/xwhU/tXwurTr1iiFvHlZTt14r
EF18Wxtt1sjIwIaOPwaN7GQletfvMF1pfg+onaCM10rHH5XL0u62HMsd7LzA
TyXm6MluGL7nEBYYEYWkFtize5dzllvttHSUfJczYeFph3xxvv3td1OYWqd7
sl5GpaWKrVy5pdfDy3CtGomfOkKvDNwRNT1QoctcwA7UAu3cWDxdANbpI81W
+ALAA7ti7XHwURy3mdBJZDqr9goTHyBty/feTJTFxNF1kIL9Lop6Tk130z5C
oft0uYV18bKk8KQ+lWGCNgswEk/bzUF6u2DEMFWNGcGOH3xltai1wXgD8jyx
LJ6af1fiETjZjK10BnMDWnuVdIA4ByWm8qrcNeO2FguCo8kiabIcReoa/7Io
3r6Wy3G6JQBl37uWDyyFolQPYto3nVuPtKIMpJepAZH/NfhSeRmdgX5OENbS
fjdUiZy6zY8CigbLAhW6MMx1vml2kt0d0neXpvM3RFKn2rpncZrfZ/jpE2RL
Cp7cnGum1W1tK7MA8hRzYJBWB91qLWn0DjnFXub16IlfvgyUc/KWHW9ccoUn
AAQ5A3MZm9+4C6zlQFkRZWuLnu79KQ32ZW4YqeSo6p0hjgNcRyyHXjehPuRC
PhJQziUg+LkrVScKcvUAEtkPBD0V9XOZs87EXEP/e2w3esvuLuXKBX6DTQyF
kWh9Ul4LJQ/lvXiGmzyYZMqK9yrN1U8zcYHYVOsOAD7aYJHiWuK2E6QlIzJT
tC6JnnwVLwWN104il3eqjeeT+zm+XZmuQxd0LRzKygBkNDyzuLsHsq+Z73h0
2/ZCPwTs+O9/cM4HTpXLyspkr/yxWJrIBfMIFVKkNTO6hEoMGFkB60eQAEuq
m/1gQhN5WmN3GkAH1P+HJQcOx7UYk07JJjLcKQOQa0QE43HNglCjdFhBrBrE
eighikGZzFhpFYMphHjRjhD47SgTSkVbcjiKUu7TTRdp9OX5KQg+4SFh+NRG
ErN0WCG0puJhSNew3OhjxTAFDj/OiiacJczDY0lypxvDQX2HrxektdG9Uzue
UClkJ3Gy0t93JVqGSIWBqYmzLKScxAeI/K1vnE0XSnGgX3822C2nTxnjz/KD
E69sO5JUwtVFLptrWFNQ2BrnxVDngqvsPHgqMESX2wt2n5IjJWceSdC6xQxD
eKqhDcN38DPpgg+s2cVR4AxGeOW8yNzaIrwYR6CEWWNpb+Z3ApLiDnyl2Oyd
khm901l+2g9vnMjdDjft1rZrr+tpS82yEr3LjyIYNKzbtes2mmE85fPig9Mw
VXKd8V9aB0esGCBRvgeNu5q168wESHsNNRhrpQVCGU8DKRPWXqX2bF0+PpAS
JMl/xjNiYskepCtR4yQtaWunBGj8AbtVoC6RrWjJGMe5NsCkUnic8Y7c+ehC
WfMxwtZ6EvZmZCV1N5jpM57nmRHGSnlV6UGDagISKmQUdgjl2FIL0drbMrAi
CNFnR7DGnFBkdPNgPLwMli7cUhvIxrgoOPcdIFTd54iGVf2kQT0J4w/gEgax
UQwL6U4HX8yjp3wjifyyp0X0ySAaVroMpB8aEKfmjwJ8fxyMmYeFkV8Fs3n4
MUQIfkCJcWyDM9Lpg9LJaGIrcfwoeUYAMO2+D5BlbML9zy1AOHiE0vkPNHiX
h1/H31VwbATkKmLtndo/vO3+Xh2x8BxHYcJU5cSv5/N9ZLus59QvcH+Vyxjp
DbAoNsG4UjI4PM3xWYAZ5DR6LbWxb6K6QWSijeBmuNd5QHd2dzWCCKLA1rJF
hEIM1Xe2xblcdJkM9vhWWWHkkfxW3tQRkOyjGeGohnARLq81KG+Oz7D/Uh1q
MBw8orkLM67ZxNoL+iKYr2bSX5m5UKdCXpTzYX6+KEyp2ZmYqDjk6ANy24sS
3g0AgL7jY0TDedYLo5JpNNFaKheGrkAfDaZ/rqQSKLGvgabucyfB7uqembyb
W5Gzt7Uun4l3YDRB69rbJnCOWoIrdFWeDmtriPM3zajb4YGz7KIBgE+Q4mqO
Z50dschK1h2pHffC0292+QkAch8kkhFdIZLE65k15smyi5vrgGnvRrdhat9q
GF5gSsbRtoOdQDPNUsyJT4VIt91tPvS6tdZp3xOnCgHOlPiuekD5CO/QAVrs
oub5Z/ISNOEUgLZkt5NhJQT6hdHObd2px7X2ccU/T/pCi0cXaGl3GBiUcKR4
PGOeijhKFL0DwnwpquV9uj5a9QAhTrvO0jGa+mddY/lMR98psDnggSoDA3zP
tGbA1MYYuLQSvhxfOKjGcmgeVvPLtmFAHaVHmye3GnOTMvPQD1ENivSEx6xA
aVW2e0QuHpegq6c+O+Uv9n8ibmT8QQcBaGq8B+8t/3W+rMSjmVJ3hbwIesJl
c9zJX0SznY8xZvvgFgOKYSlp/anykXf8WAiQTkB/j9PsYzo7yGS44tPmWV/1
l2Gk9I4NooVAuAxZiNm+tQ2ESX2N77JJW/8tYnVtsC+q28chHLB6Va3ZphFv
zvBVnB8+kUwtxWYsO3Rci+QUwtPQxtjzRksLC+8H9k0eNw3lXTHXs1wj+01r
F0zLw+WShuLvf+3rC+dKUGp6ydxxYG7cnHo3LufNfGVb2MS157/27WA2ImF+
XFanrxmuH92Dwd/1ZdSXQPHu2UF0oq9Sbj4S54gDGbpBeq4oTB8eS1l2ua95
897OVsL85KDDK3yG94VNt9HJigpMbYSsuQNtGFxQ5NTpgmcLLdMcAWrizpJm
YhNK4I1YJC6cuC1UCULm0XjMH4n4uGkUsd7Jh5LXnTEFYl6QgfEqDk27OBwu
6mcqJhPeFjOvH7f8pmFPUQzmTUNGU3dwQf2S4Zsnsc66OJ9FCJagXOwVWV1k
ccPo8Uskr+0WM+6r9OIACrfT1PJ+86nwi3hzYxxYJmo90o/7iG+QsDbERcfg
UzVYqup8HWBIiyBub7pISWssrxYK1mu1GX38Nh8vKgdWNJ1Ir3eW7xmcCxyr
LGzHSSe09ssc6fR58sJ6/aXatYZsV8bK0eWqJf7SFvhp72TSDiKE0SqtY3lh
xdHxzPQCovaAm0xRspCA9fZf7MzvFzlf1UrmbsEzJed7W6u6AfBl8h4cLfGC
M1O22jfgdIHtQnALg44GKnvsn3oj7vOQcFleiOjSImuA6DUBKXV7tZ99u17n
KNebuWUkNPnfy27k0oHWXZCPeXzPIaWQ5y6uAZCgAcXv9dWmOSFRXHK/Nfbd
lsU/WdTs62AOt008j/+gR4UeRyEA/rnnL11HTJfJh708yCPJxbIB93TwWRtc
weaur7JVp6JbujmXBfnVt0KKgJTqtbR1BoniPYsZqhQ/uTbXC6oYF0K0mViC
AokH0eyh+zxbWXqZ2cqcQuamHCSsupuHDFRE80RgoOanN50VD2FAUT38n/QG
wdzdxfM681mAngcukZL1B6WAP/ivupUciTl1pUIg3GSx5cMPxj5GgMCVlQP+
C19YDdie/PnQ8vfTRlhDEubDnVarK3Gga3qxYFzAy39vXiEhfbRw7rzbhqMo
mP1xkimololTZ6L5r6DqfMbkR6e3tCB+EWu+0yEBAc+QHAUbik21cqoc/sGU
TxipyRgNclq2VsSGdX+RtrNK24gaoXpN/eVElw/FKm3sIIk+N8fdl7yUZ+Ri
b2Mnu84AGYQED3V44wF9awybn9lNhCep9AMEb1/yCvsE7vhN7sgheuDFTvbJ
Ax51Qs/3H9MLs2Cx95Sa1syDGmYHTuRu3PT1yX6Ifoimzy60CFAc1qyUyILB
SzOjCGWLIz3f22j1mBEvs46qripl6tB6mNuLyPv1Sg940d42UInz7O8RLC0W
qWRR/nn5nJ2uJJYD8Uh/e7CwjI+3X8rTO7FGvXHneLQLAgWiP/pTY76RHuqz
JEzIzOs3xKMarwkpGynsN94GEi5D79y+7s7C6ct++oJqJ2+Crel8ZGbbFwVF
EYZHZ/eLO4Op1mxGGix5mUEycJC2k21dketO1T937saqhDIf4772O6BYzl/E
vYDjkesImRwEhtCahitXN0cQKEk3Tz/a8uxq7b2HhpEJG6HBAhfWQLwfPavm
kPAoYrL7HWoTssyHfTe8nlsnhoGd5vXPjIP/lyjskq843Sxr59J9x8E5/2wn
77CO/45wcmvATM8R7B2Ryk/e97SYGTMtoSqjj5qxVm23EmJ/ibBXXtIkr199
pXscqXyte3GnYAvwTIRJnVfb92slCs6l9YfAVprdZ+SWcdMTxW99ilGWkQQ4
w3DVMOHKoX+boOwy2gZBBgJ74961b0Lqz+opApIlRqJBO1M5RBK+4ToZvQQQ
fnpUgphbMyBDUT8CCaonkBh/DQQJuajoyK5vePGpQyIGrP2sQQJqpAx9xScp
PCUYnfX0fymXXeRt1udatK2kbet09VbxieYRI/KhjpV2xjTe/7uNFbhEJdIP
iT7aQ5c9C32Y+ohIxZXVb/6bp896YQyIlpJjykO6oRNo871libLk/EZO9dBU
gP3f3HH0tVlGEWZPwCZmWskIwWssleM6RteyFqm9AoY1ui7mn2+3LQh9UWZ2
3JGmjn6PxdVd1f8DrtmopDw6m7o85L1dwbVQy+gvCMPValk4MvhF3s1mPfES
QlWZyl5EW48UtyS0mjVEpL7K4pKRhllI9G8WsxSPnGo7EKYBLOJl5/CLqgnY
IFh+Bb/CCtVMmD3g8zizOpk29vPFptbT47Ic6unIPRWXTsgj5oHPILMf3nPt
vyPpFwMbOGh3qrgRjly4HfTkT0f4sjz/Vvl1NG4brNjdHnMqhoux8FwIkr9P
hElPd0U8W1M59pHjpTc4Rc/MtIh8jW2yBq64dfQvvNyKgzA6y7UxlHzaWy1B
uLeD9H2kVx4Q2N6tQFyKzltIfZzTrqlUskMRGsGMKD4+vLUsrQKqxml88OoX
t3CUY8Jzcgos6Y/R+OU/LWLajIjLC79xTtv8+wzyg/3bRmWTb0TNHpIKYh30
EHWzmI8yzHX9dTTzdatU80BBb/6YmYnwh7jHK4qdINFlWOHDoRj0VJryhzuo
WDwt6xfIHn/WozHs35p2ghOfqB9TOjoCuEo/ELlXy7K1t8+SYEhZCCz0caNc
s1UNH+PiN+9JsTbZZ52fAjM7cZshbwPx9STMSWj9drdJOCprIsa+gr9+FuD5
T3yX7lTy87agECNANc7t/4gkGmepL7d4ykhLam0IqTwfqwbqMFzJEJr6kgYN
XgmZURr5RKZM4znHBYD3ewqQAygsc/pzz8Z9et6l/I+5VjjMNlb0nM26DAGb
x/8L+yalIk/9AYLuFwZ3k9M4Sw1ZxdapatMxNx7cpuIYIEBMdAG+/QO8B5DD
d0JY55TZ5yuII8AJkA5xfWL5y4ohKD44FLvtjMQJEo+mMgP/BQQcGmctK8Dz
jhicD1Yzk4dhTXbjoWnj0xOoSg/53yALMRIqG5xkFCY09wY6O8p6c4FUeBRa
lBClqUZMg+024S/oChKXxwrbWrcST5tbsyMHp3JTh6Lw8yHgrvhmCG3/CtSZ
LXxQTZLyupP6tyxG0q98o46S8X/4yEv3nG0ZnO/aKmwSKuxH2SnXMFMIH+QK
feUD0/4sgEu6OD9xZcsErzSbYeuxtIcsBdvptMrbUIKczVKqbqLR91EO/yZI
a+pWJy2rfZoSJnxv3ZEnSQgUowx8oRqNX87fIBClSxZ5ZToWwsNbkVRlsyPn
6r8F2XhuqMF0XeLWsKoRAVsmjyr9BzKIQoCwtLCzEgZBbpM8XFXBYFimxZQj
+ToVpc3VO3fGVYDb/XAz0HABSHxXXERCCDEhBqKImaG/U1gS9P4jYtFE+JH8
lU/VQ2cflXhfJReRJCNQKeof0EKN8nPFW341cAC/DFQPaOS9yC+6X8aL6HFy
0cDN18zs3g8GBypuLmH3TPb94RrW7jup/et9qikOCyGBu2s/4GgQ/8nbcMdv
+sbe8tG6mYeLBUElqVz43uL6svMSfRVy0+slfc+9Jg7T75pXjacQOBpozsLK
n0G80zrvO5M13eOfbGZ6JWCNnXTUkFHp4N2AAyH57E9t+cePFgtSLc9WSOHL
tZINiofD8XHlpnskrck59ivYJA5eu8E0KvdVMYe4CXFF1D0wqj1pQvwmqrrV
L2bVfqSqjbvcWZHu5FrUQ6SUo98B39bVjz92QnLG2IfQg+1aP7KJTOI+DcoC
atC/j1DtViio+eDAb6F6pLP/+6OkGgU4vltSIeKRydDjd8Sxn13IXTyepzQV
ivrPI7cXhYARN+H9sAintvckItgMw9n195cp5MYJP/nTCda35JIr4ngjk5xY
0/aHczGz/cfiENy9uka9W0lBuEgB6Rdl0msLKjGGTg95yKGDxklCnyuYPovm
c/HjIYuqw5CW30LKAT0QlbZpni8hyJ4by6CZNzWvVFrSCLpMkTE1YuYVw/r4
nwkgUrk99VF4JuKy2/DVFSp8dP3lNK2arJ8IIYKHqmjObnBy1rmRmdU9C54r
QMzAZexfQTHXRYMnNFpAQGuBjHgRdNhd6KK0myt18KL4aTMY/ARYGuIipV28
hEM8vF85CznKGxhC6XKddGv/q3dT1Pu8uAOOKOu+s2lDhQTXHvAyABz9ZL/S
HpPkhmBR9K8s69/mgd7aE/BpZ/GVjgaeZu1q+jAki8QlELwVNgLyqaiR9bKb
nGPckm+pme/1LCjvAmFxU28r1TPw5A/2UzSXz83hOxlSks3njNzhMSrCwIYH
dlVNfYrbmYeorTifTzttB349jXykizeNagVdRjKPgDJVPpDlorKzLkCQPSVI
Q/zh8I3JbFc7bAae2plmzOcL5SMVy4+MnwduhjM+zAq8/3dWm0jdt71afyFd
qvAc17Hji4Z7/ZonVt93yrD7rldrC4ti6FY4o48K1+7WtWdrNQYJT3zNmZdA
teuJaS85B8sIkxZh60+tOtuY+UzZtryrAQLW1Zg4vtZoDAGUGsMLM25j9sJE
8hzgSQil7s/FOq/LF5gWfBcV5HgDBD0XItU1mRFSfNx8zwap16XPndaWL6Dt
w3GOdnPaaJbkjbM49kIRUPX9ZIkxwiTsCXKNgCBntWchTrsjDFejKuRQAQ6x
bhmhU7nR5EG+iGr1GUTtbsBDGwusrC78BIn84sMr9xIwVEdhh+WCtC3UmxOh
3u3IV44mh82z8FP51wikvXkfm49x7IyWmIHWh6d3Wt3xq2Wq2XtV7xTxvsBI
Btc+Vf0lzvqD9b4vuKPAyU3o57mHVvQAvhinkf5aIysMvI9wWbKyJduRSgWX
VjuOtwqNIPSjRf/zdhPACwMlWY1X0nopg5kODwQ9YxYmnDzBBB2XLaZ3NgQD
HPuOCnc6cTHyD0FN8XMz6vUsGqkVyWH+YD8n7E7PBPOMNCM1EocvXCAhGQRg
T8gDvmDVKODZg1FlAGj3vVW0qNzsPB62rtwebrBldNTPMNUXHj1P6VTQhojI
UEj/q7J0rINg/eeTZU8b6Gr6lxOGjgPo791Yc935Wd7QeDTvfwmQbdbKVGa+
67HqTR3D4lXPpIR07dwOjnKuVqZDT7l0IKX8t63OJwDbE1Qmh5qtHj9XhlLD
vkLoByKiftXT9h5nQX1CKJq+dhMpMfzkO5Lkv/Hyd4g5u0XcZh3r0jrpFiqM
BgJaw6wWumAOEKhS7Kv6KCRaToOE9m1zCw2ywnfPtpp/thIKtLCzylV0fS+O
bk0d96eX9XFfGbNWaPjZvGYpUualTACS5pRaejR7C+grhMziMGFdTfCz0Zu2
nLSQRT7o2Fn2z6IxIy+2DSIRLhe0a6dwVv7PilUDmIiyG4pYUcg7Fog7d5kC
h2ek0ykL7CBC9bIBLX8qwAqNtxNU7EVpS23I4qr/5wQmxtolDMG8H4gDpE8I
bF/ekOUhkZ/A6YhVrSW9+ao0IzU6z9x0oI9TXQXybm9+/eKmHbXYvPoeOLng
o2md6vd2jpnlho1rfS+tps0DB46GZitoPcyBsE1LKRO26KbMg1hgUUEnsj0H
bPelJc9pPn/TQ8S2zww1D9Eld3nq4+IXHvY24BM57Qnlk1jHhf8+po3ENPDv
cI9OEqLdCN2Q4wI87ilAVAhXps9nWrrANAUdc71LG2oB7YO8pLKwVOmnkLRm
uBfa9uNHtUivIclJKyYforE/9gV8HGTKj1/YGfXq1d5r5n/pEiXXpxQR70kA
u+IWzzNmh8lqldh6Z8i57sQ/yXxPzkLbLIacbIScAQpFtjm2nrYkzVV8cNgJ
EJiisghspfQkChDSjxmsQ+rH4a8FHvji+aKiu7wniaiZtF6Gt519Tzh3m95R
FR/t+BnCLUXGT/Q1YbCemIOJXDeny2GCAsKIgbv+bhEKqfTSQxyIPgAdfRkN
NMwGUAhYbUI1dKZSoRKVeWkwH2qbMSUOCxqioCmks/ntPl6gYCLVG1nGOkPo
6Lzw4oJNAS7ui6wNGmMdOv6wi+wXlgCo1AT4zAKtr/Tlwl/YA8pe4jnKVCLY
1uhljaYVso/wHlFtVMGihqFkh3jRAZCFc1RvkSVSYtGgxL8nwSiL6SB4z2l6
wcYh2cJ1G/X+vpIBU34OWEiBarzzTdnIN8Zedz19X35OCnXYHPP4rIkBIAzQ
RkHFttM/a/1Yg9cMHBhZu+IPecWjzGCxrfq59fZNhw11NcGEEtk+b3jXSKq2
0m0m0HT+syXFZu8hee4F1RYQMFTClg5BLFxzx7JwLc++dXfX7WzojM3Xbcrz
HyOwg1B2aeHHYB6R6swfgZcz5n5+M1H1Cyzg+pIqf3FuPcBpi8hQERUt48/b
wS1OQvI2UdaCQY1go6NyyCfyFAZf+ShMad+ShVA4fNoGpp7zbhZzJeW6nMUh
wJ2QsTF72E3OgNAaCi886bTgn2+YdtbDxOqGExKOswOEy1yPybc1DT/YdSJB
6FLnF+CeREYaNin5tpzBfFOpVudyJjXfvNoGV6iEV0UPMaizo4yAJswzbsYy
T3X7QqXKgqHziX/xJ/2iLkUhAk1OkFS1QmA0YoMHSgZrBRf72NI5+LiwlnmP
m1ZrGXIf2n662+YCqMT0urZyVC3MyqOtXGYcPhGKuWzHOtKuRSIAOPKw9bWE
ZzotIZQr5uJx/U1RdRN7DSp8R/OZGxKoHDI81g+JvBE8+bH3dNzk0QCbB5HX
ZOHMW9OJAiF+gmrT5vwSNvyxoTsHqrxHOe8QMUIeHKfJY5N/hGTU+pqVdtXL
jNlVmxRek8kN1UhJu98CPTflksgC8UKPgBZ2hr/oEB2I8tN3YZruhY/aLfMh
fvJB2xr0/NtX2EAFACF61oriK9qvJqSTQTHIbbDUkWN50Rh3JogBgmzDNAwo
uTayKM599NEDhhvwCPb0iNcLTX7ycoaOTPbg87ttKziyPEHKZ6FCxkYcRMeD
J7bVbS3b64lmkZeAlcT3tZF/uhDfm2OS4tEF2xaLOn+x8Qtev4i9Sr+pPN64
Yh42seI/j5RSsTZacrBaC2h0lE4rJSZMzIGJvWMIkjyQ374S3YUODyZFMew5
95SyfsNIYwVZrhQ5TQLci3C6snqC8qjprbgcLPSTOvdA9oIor+2vI95ZbrvK
UTcmXu9kGW3jojP7b6Zeri+WW/qxJJEgthFnvOTfn8AavCK8SuK5nw8hc3Xi
zfqboai1rUILEaOzyS4sRhOpYOrS0tIsf6b7ymT750mAMyjANvsd/6b93pPk
Z+2qyCSJ2JCrBoIqCxo+bxA0yRYybbbvujHz1wVzTyZYmiWm3SCTXk1ICcJA
zGgy4bRJysiyy6JGPcI0zXl9DIx0h9p3xwsY46Z1verCgJJIzcVbS4q4ZaP3
mpid06iAvQiiUq9WkiO5Xj0Twrlqx5wInEU7fBKDb3Kfka7nrJ4o9rNgbdkF
owOdWNpwXCIwsInkV1CcbbXGn1J1XFNWZiSpDIgbwOBxQdAJeUq+Wqz48yQc
fjk1RE69CnZHkjiLbAJzXAN0FqtjEBdcUA/v0Uy5AgHrnI2u7EVKTs1nQpmv
KA8NxZhdCa9+oh/NwLauzvmKFbi8v9d2t39uvXtf0wpMqzJLm/H8APGBQWwT
LckzquJrPU5yMhY4FSvLki5hGXAR56mEiBdFv/9xoFVqHeoA5fMFU9SP4fz1
tv4ic5vWnovqIJiw9U9Dt54LfE7vSJ9rf6TV2YclTAuhSweZ/pDmOylR1TEd
Wwwz5UKcZ34vy1R+HHi3q2KQVB1nuQN+IA59JuKcasrqHUOu+Uu1GKXzUFoY
EG53sLgi0q6NHXJq0Wdmmx66OGz6Ed3KVxKeyMdIjRfHQWpwKKFqNJLzPrF1
m9CQMR2rxetGVjOzy/1zOpRXrVFPfyIZzY92oZWDZAIehK2cAHb+0Z9oCE7k
sxdraM7a+rv/jOr2R8V8qJliTMcirgXX564MsUXmISmTsDz4w+Orji46YL4T
+uP0/AmZ4qD9lbRBtUt6Z0h9awRHqYkO/EpC7Vqh05bImCPGlsQB/0U5XBUV
qJCXYg602KN3wHUvm6JhresMIZepbnMMZftJUqjlkamSP7wJa6HJtfQ4Gysz
JflPfbJycWYK8xE2r5RzB7JUONuHo4nzNMdyNeEfunzcEp7Msvq1gVWFyw2l
1DfHMQ4qLy9chBMwV8XZrNasDHtsb9Gm3mtG+tD8PGCrKu7JH1DhvhFce574
koaRZSegpbaE0GBtpJGY5nGS1juCyyio4jD1DXWkHFenUszs5Tu8yOoWMe8Z
1QHE1eS5y0GquJ1pCaqROkdPzBB5VzRus7aiWAH9tUouRtLzqIdnPDfDU73u
suOnOIdHJgoEWpjIJb/Yx5C6ixoGIOMyFVORHJOOkqADlFgcLJPeHOrS15Yz
EruJkrEfn5HxU/HwP01LITbP9O5fUzPZ01jmsAtz53erqHa3Eem3EWxnIZT4
IuofTLNov3dmQTytFUzd43wt966kF1vW9mfCcPDGnXCEkCSt2UrqB2MVS5Hc
uEksT/FuZvu6aSt7mxoJaxD20jKFYL1a9PSTo8FRuWltOt+aiVuiFEIJl7hm
gtBuQKk1gFMh33BNIo96nk7g67ZobOMCblsGiHoV6cTtQR6xj9zqrh0dtK5G
+PTmY6JTggwHh9koXD7B+DFRdI2i7CFXA+3SeTu8cdCL5YpZAv7ZKA3GrsSc
xLBD3QFNT+Onb467jbclLvlf7Rw2j/ebHoqSEYQb1r0cu28WW0gxE1zbaKGL
yWwFHM36uWVeVhEeS18weVUr6ze4iCBC5N7lwauND1hNh+5LhAW7gL7fUeQE
FO8XHvnhUbylO1cHOVifSXZtnuKPTj5bAAySEh/piFQfyaEjbjwmbVM2tdd2
Uz6hS4FvQBMwIejdJ3idK4u6g8bMOVAXSWwUOLw7dQvW7ErDS4nXJB3f40F/
lVz/b1ag4fva8ZwiwQIApCuJR24h2LqE5uQGD6UW7IXSmvEsR35BWifv3wh0
bo+o0cEZxmve0BNzeACBd9p+50RLKxyf9kDVk0pqNl7kk7JzF7yOu/+iLkjn
3JBH2UXWYx7XCw5y5fsCkueAByAxpLmAW+RUPSjZ4V1PlT3FB8JygRIwWtdF
9Gdot0I+GkDtXcXUe4Om73d+xzc40Yd1xFwCCwGfRRioYwLM0tTK0tOMybNh
QrmwHdT3EXsCPpDg3vHMNQt4mbShU9nBl9iAPqVXGTC7Hh6OUuca33mIRyrI
eA1R7GKJ/HVCqJmC0uAvg9cgqrZQ88EyMrQxVGuYaAUe/WhNWRm99nmNbl5C
8FX9BVrYZ5XwkEs2QbcHd4rMHg7tbgWbZui8A6F7qmgAjhmDWsPur3aCTYdK
SwEfSEPtxlK68Lk6axNKo658bo+nGjGCtvoCCHk2tfoErqRtOP7iKoPXd90r
oPjJ8Z2C9UlsWP/TmJ261UCkKXj7pFWDaNTqrsVsRwpgy9ejUwlQSKi9CWHt
41lAPq33j4uGanATKcxUQ1ffVFeRaYKWefc3o0dcgLgoIeuhs612F1IoY8VX
AbEPnN/CcO/y5uStfb/rM+K1ECz0sMC8NhsYZ2Ivkz+Pb3lDEEZDcit8qRQo
n+PPU2bXzpWVM/g6geyNy4tMajK622DJ7sVCFScd1e9hyy8aMgwk3eF/rHaa
gaZ2BPDdLqltVXt5CYjTjerqGUryvaFeEEDyW4o8crmLX1MFd8ROrB2nPqvG
s2KRBx6dZRjkQKkrAM71u/u1vfvdL2EXLIcBv0sYp1bUBx4dOs0pws1meUPh
hmJtiVzwX/XK4ls0I3LJPguK0BZ3vIz1bK5fOxXHlKWTykHngrtf/OddUbNL
bhlzJQjtlb+1XsxtS9KAzcuTB/6Ksc1N/5rDmXIw1ZvrA3TCtYHuw22uYCsf
X9/iuRTVLbzme7YBJDZLlc6k64G60aoaD9C1WT52Zl8djK2CO7yoWX2Ea1Aj
LISjC7hUfeZEeXSHMyeqYehqTzMFUjdRAmJiikz+SiPNcIDHGFk632b/mnI1
tjxYrxgckOZXkFYWOWmOmOPxAu4vD//v9pBweteEY3U9F1IcgaYrRFe584zL
hAkKLbSACxmIbdGvxjE7JzrOYmA9OnSd/5COa/QFRaQdSFqbwjjX0qB7EDCb
jqvJWyL/VkbGdKxf+JzAUzRzVpHwf5S6t9nZMdaIiouBD48N4SDE6c4d+rTu
Fu73nbi9fq+HruYcmVY5bHlgWHxkz9gw8OsZbkXElGHIeyEu8wfLC8AcK3Kg
TiamB0UC2v1zkQhvBXfNoPpUfswGnH93UFTG4vouuimBhmp1hfWV8slGjeJ3
Dfpins2bbEDMhYLya+KJfUs7napmDyKuDMcwNT5BBJy11uUKcFRE84ZKyz5K
szO63wz9aSGKwcojwE4AgDEhMcQJgMk1Q4KU9sEhIQGnfYxysaH8lCLECX/V
DlXsZugLRiOGrQRICY1mIm0tLxk6ivzXT+HS5M0bnmMza8oAr9yq5F+L6QcL
4DgVUEfa+CEHZ5yVsx/CowW7i7FIlK/rwqlxRjTg3fHbAQBkGAXxMH8lG2Jh
Q4ROXfsLgXj6n3xezS1UNPyPj2BR8yOH1EWU7CDG3VqXlL4QDs+BkmJi/v3M
KHZLA4/mwjV9UdwOgzrCZ0iIJZJyhULUM5YEM1EnYBe2OvaJNpTohNmXGMDS
EW2UnhWdlCOPWj3gftQ2GPlPR4mgkq+jMCnK6yIT1siaI+Yy48t5qUSzbdRx
VTwgDDIDH8JKY/p2x5WDkZfW5iax0ZAADxKZ7AseghGM2kdJH1kO+VEJwg5l
LifBRbW+b9MQghwwegfg5p8gCKNyLAbnaZHE6t7aeBJzQXIBqfn2G/lceJB4
w0pNrQI0gsmljZsxBU+hEyrEgTsNISGM6Fp3w/i7Uu1h3g9l6Uarc9JKGyYc
A3dpwhzFw/vfKwcFujvU1u3mz5YWi39txb9JkBL+q5aNp5ZQATS77Y5nzsQW
IFnvy6EwrXPgJqLszS8O5ffXs0hGnbwZWSQZ1dS2S1HEkrUcpbjYsfReYQjs
HJpxFzNnUBi3gkEKVE1fI//GhwiLFy8N9LN0LXIDa62bccRiaBNVZ0CP1FLi
SSgPxwPUwl1YK5JBfThj6HMcjHHus4uhCIWsvU1MJWg5RPDgv1IZjjBSQaN6
37xi2YD1EWRE+auaQ48VwwLrtFXH6TIp4mQJVkyEcfpt3kRMMAjep1lm0elb
w5RT4V7X8KSEHWw1oPeVPWbWvmgcqPYgGGj2WNMYFthSG3qrO9/JiB3kXWgv
SOrxWRACXSSxWIArLVLyAg6YTvQfzbMV2EjKFCU0gOg7Qg43pujQr5uI5wGt
sY0qDvx9IXUPKffvWwNA9yvzvl1kd6IfYht1W8uV2BpuDfwJxm55C4kopDWA
dPVMayJWtuihc8TgRsjecMFb/jKKpP4oFWeIFgq/cQ+JmjB2fMIWeAg6jG6D
u7YSyqj7/53yMYICbLn1Rs3Y5UDZ8KAIJllooFJK7ZqdQ72JHD+Yy8vPWQfq
S4uIyt/cH+wMhoHRrqAmDxtsclLNcHezzdrD6A/8UG1af/ch28p3oPWNHcwW
GHo1xXct20BmQN9pct/q21xvSfeIz21VEkm13qgZdDZ1mAv+0ooUy/A6qsVx
ppuE3xmjMrju02QVscjCzpnJjWml4i3KRpi6oNnJlmGYUDkDkcHQ5SpibKEO
1WS+fZynxqWCoECFxypDUnUFZ4TYh1lvXdf2ZbF35LPMX4cssZ19g92P17OL
y2ZkCYC4ESL4048pgOnBbnHsWcnVyO7HReolKDOSObnzfM3yFYB8SGK8YCyg
bOeBSGfviPxONw/hgD85XB/6RRrjUwiKq5IOBnvtgK+qnZLzA4EBOFjO1WIF
OpyDAUZc4ObVI466iP0zClMRqZTlMCVr5wuGqHvXxFHhYYY9M3LRmwEWorYo
XFZPxd7NPQdZQQt4YaPPIRFRJCpSA8BGoROozzN3B+HHSfoFJgrlbuPBSGRq
6cJSH032i2dj3cJJudL2W95OXaqqdy4zgpCKYplWymu7m/VayNQsV/k118/p
zxNU+yWiRA1+4RrOJb3Iw6TJDtmQzpgL+mG9AAlNJ/zHeOICBnsgGY2clkvz
4yIlHKJ8h5IUPiBCSPry8FCK1w/R8l+Rm5wCg7e9XMxz3F/PjvcTjEAle0pU
tTbkC8IqTACJ+GxoWKakWsL8SNgVdw5hkb80ZAt/LJWogKVxQU3Yh4UMBi5t
jq2aQ8rmtp+BSBDdmBbYIEyTd9eUP4e76INmg38YsQJVpc4+su7GYHwNn5oz
GgUqaZMvHVNZxEykHO6GtIvk7VD0x2T4v1eucw+E4xk+novG/PS/bauPFrjR
ZLtkHSqxlDn1JmS0FBrEWcGRjZQ9AWojRMaO8r9c+V05H5oqRXpw9e9WevHm
XvPHhajrWbtI/KUgiE+u6zcSccPRRzbx/Fi8gM99fIvufh0VKLHxezAahpWI
3zneBgVIMg+dzMxKLAFvn71sEK0YW0l2cYtRjtfOK5b/9dWSrDz4fu2kVvjJ
TAMtLPKwHfeZHX2tbeEJ/uxpZIZC+ar+y8AP8mI9m3cGfO8NBknRtHdsUxt5
jOXGxcdsLa/2z4t46LcvsjeKZRlwCJjm//aKOYu45/8Vk4sNqzCQFf54/8Dk
pAxmLzMz7BaX5BJ+EoRITjOmmaRKj5/ovsjzxLAYZVxF+dgtrUdv3ZDTgC8Q
K1RkqANTbR2cwZNM239apw3yghngouFghZi9hx5aqJK8vTG+mfI4alpD2/nj
RWiZzjuHysCBiFztxE7CIWfmUgIwhag37ABU+rDMer60YAuM/zfEZtvMhqEl
C6vfYfIm/EdIkl290U67IYnlOVvEZ7hj2ApERC7zeI1e3b8d0xxejUqC2UON
nlQ95u6jR/9cullZbz5NO5M3309F6xQnJilIEc9v2Qesh6I/IxWQ4y1ulWyT
ek7xi+riAWmWeP4VREbUHGqNxmjNwwnQMqjmmlvdCo+FHB0RycRCUdo8v0o9
TTfHugdZ7cxlX5HQ4LVG0LQxQkg2wfu/g1r2Fs5Y5mEHAKhD6OP/36HdUU/P
2bFvLXV9SzwISiYGs+comAP5mliK96eWhtQUNcoCYbwNCjrkHT7lFprHX95Q
FRRy7KkMyO5zChXCrL/28o0jk/9GSu8q34V2bV6EoiqP8LijC4insbkBXGEG
x0RyC0Vnn7ly+p4I7+D2cd8wl+4owpD3DJBIehZrnSaYZwhHR4XW2Jan3e4A
BMIAsFS4RiavUx3MIIASFnLhYu93rURjZr52sg4hHnhx01dXcBQSd9KhW1Rx
PP4XlhrmZfq3dtT/+P0Ud2wAEKTtoqrNwCCLPmwAVu7az9KTMJKCZ7BcXhuK
KtamyF32RqNLgktsdhAha5Qlw13I/wF/mIFk1KZTxG2QH6bkh+8mZpBD0/T/
xNFcpFoo4ShOWfj6Y5rsHaIz3wTrQAeXdt8mIX8DZG7ncU5XAthhl/usNMU5
3up9EJ778RbNsWVTD04pYi+RGX6zcGiDLDLtlkTuY+Jc7Od/8aDE5cU3rzJA
GSk3rE5sNik0RrTAag5AChQWmPaV9gTgkkVHAghoDhldEmbxm43tS3DxR5p4
waEO33ktFJj6nJUxZBbdiTgjfL1Zf4yyY5bGtN1kcywrrbr9I2m8AjXT2Zal
nimm0enaLofie/V4KxX4TkqW0049rlYn5HyaTfWuIfyEZmzEhPHlOln49kpe
IEBU7BVks42b4VPV+eaE4KSJj+9dp7WHAh7sf0EQTHKgpsGb5fUgbBgStOnR
18IUVwsLxzhDn7lxOv7r/w6BEB3UWjRoNmJgEEFIlpBjaO9Cb2Aw+TlP4j1o
f3VaHvP87LAN6mm8umUzKgprQEMflU32DBP1btkj33tvqfn2XCLUTkpR76gj
5YIBhx6+dDSADW2qFYJbwlehH2SZn089g0D5HGG9Gzf3tU5T8dz7Lfh8zVv6
7Nt8tdpyyM+ZFzai+NbANRU6N2y6c3k0Kp2BJF7u0HtuLkr5GFf/BB1oGIAQ
6TsyOWgIVBUHv3vI7aFWhIsz8IIHx3+OVQz2kYiuMfJCrRHDnYinMNr+Yb4f
m0aAs96pkiLZtKv4NW4+NlwLfTVfig5788IRYAkUuRFA/KlEqDG3HZnmO0L2
hxwgumT3OPX7tUNl08emJHpBGtS6uVYvH3jFB1r1Fj5qFvdTmWL/r93mH05V
WJNJy0Ad/tfCT+OCfEBRzU8uepaCShkNPYEHS5xyMtQP597+XkMGwYT2/M7l
S1FRwUcAAxN6o7pOlm46rjMOPqpIXj3cFz5VHvWj53qOkg2sGPwkpVUtJw4z
wKX45UO6yUKNjUlcZgq/1edL0SDZ64iCaq3qGvtpddd2LD8wGVSb+ulI6ODe
myZ1Oej7Wt3jwEgGJQ3618I+60VgjKshhC5u0k43Mjpf/RXvCbpKRHOHC5GA
U+LTTM1PT2KuozSgeEz8Alr6Dy/b93px4f7HdJacTaJEuZ1JknFZsF79CnRp
tYOdOQE1mAhOd5aug4jFs78tvI6mgMVbPqh6k2tWd5ulGSrXQHynYm6jWc9L
mkNJMF+6PLDy9CkPUvi5LtmRyDBt3a5fX7qHEhP8aGnAZD55cFsSgN/byVzX
XQuup6AaiPB+2QWBEDqfmljPPIl+2XdFPnziAFwrpKwH9x+pZsHPxszp6dse
jQRgEeMxIyaNaIezBJnGtqpiYF8NMXylW+JEZ/tI1kISyZbzb7R+Jw64yZ8z
3QlUARssyfiZtujpf6gdl3hczhCnxmi+TxpAaejOpAzQ55oImCGkgqTfnJm8
y0eSwonuX8DR55lbt8Yu1qEoaRXidDbCi1ZZxr/KVE7CHoH+FCSBsc1MT03t
cMmV+gQK1cLclOQ8/0QYdXA4nbmPdFnZSluDNGCo5YbReppBI1ov8B/rNAyd
PancDxx7fYW+uelKqgc1ZyxpIFHjJFocmHkTVf9QF7XR/vcv+cLj8HM6NOpk
pRAbrb+9oVQwoFtf3g8feuN2Jfhu8+7se3URh4a9MTAoDDZAG9O9WE4HaESx
8HpF9kST5S1Wj8drxUwJySvN+EkjfsghSSSoSkyytZLy0Or1DTP7wG1hRA2j
YdyNjso9xaM+KEWj1f6s+ZYgFLq9jI8LGEhTAiiiEvx4bBMKkp52NRaYQqu6
8YhtVjlifDu7ERsebFSjnUvs08pl7cG22rd6IB46Qb7UNceXzi7lZkL10p29
7XGidQfuws9VGYX1mW8Rg89tmzq9qUkO9jka9n66mvFZAjOUvpv3p0JTWCV8
kuhGtX+OmD19Duiu90FIKT6Hw14lhOFMNg/MHxImMmZZ40MVVlTRpXxK+kOd
H+9GqghTzIsjYfY+sl3Me6G1HZWMajzdBinMX8Mpahp6QTPEPi/JEUz6GlfL
IGMuoDyvrl/MXNMDYQcjJ97HV/HszggUlv8oVT7e8zMqMCiZZUUBmZPjXvah
tp3d/xvMeG92kbckl5Vy5XaUA+cz36j7gO+jtciW7zNHnh5fkLQ2htDsJ+mN
E7PrPTf9IfhIESHwMeVEW3bgTmyjFM/9GVGvOVHZTi3fGGS69wgwfpTgTZvk
rFGbtS9tsPo6ygMtvhZ6/nXvNcxCT3FJi+XjqSJregI3Fee23B1OQhr82Nwk
VMGhopNPmfkUZiBbtO5SBPmup3UG/53bUqZ+Iya8Ks1xex04Vm7YozRdEiBs
RiDF4pXWiCqbp4ckSIXOO/M9QPZDHgEemMj3uywEf9RUj8lJlH5OXlDdg2is
Lrwu+I+PmxWHMlQdtEIPFXDk/moN76t/relY5xAhr/iwbbO7Ysh7w0kqN7io
Qi1LhPVnevgWcEm6G4QKk2VIFvC2whJLx6pZMDdQo9GZEJCKqzVH9O3eqhLy
nYK0LkA+ybRTa8C4JO0eSttSGluCUKU3KkSCvPVCSBWu8Q9MF5Ee/jlUlymZ
GSRlpKM16yx/hm+nq7MkuCFTE+gO3p5OYBabHD0lhuOrTJ2TQokAuKUKbcdZ
+q7Tzx/5paJElfoVZCCqvsNwbjJue9RdnZXtWG51MyIu/DKR5WT2OTs4FCv2
8WfMzQTO4jv4Zuj4+bg3BCaAqfQwsZxcxAyJ2L9uEjRWVFqTTq4rdRCvzMnj
2c6gKj5uNOXxi4QMIQWnCSXpEAZ13Bk9KTSS/1rjcPC/10CNk/dSbpWeKN8k
56vWevA3EA+dDDeDJanoYbRXNFvvLKZtqhauhyXsF2G22IkP6KKp+MjCEzjq
/svMAAKRBUQkHC1Ocxs+S/yg7wYXjObGtfZUVpI1qIMf51ttIkebvpcB9OBh
cvyd+4H/BAjnK1EY/oHaSg+fAAsPIUFU16VFody8/pPPcArbzJMrKLI1tiE0
kGGmb2a7IwstT5qKZHtQfKo5wVMje6NbWC+pvbONr4ArOZzBbsMtKZJ+fTq0
KxBRdbou3knTvhC6uq0AVdJUV9/b3cdt7yTUZnajPg/Cc6KvnG4St6zB1a41
DyTy7ndTvZWOAjbnuASm3kUU467T4oMUkM2TCxWr3Rei/lyHxC9iGlHMAgqk
kmynSHLSMkrJHvhyQTNjmHbUcplo3vHbQ/vDDHClFeNXR7GPo3eRxjzyPRZB
NrGX+bHCwpmQ45CkpMA8gYYzeryfxeO2G9XyXjpPIbJmPofgy7sn6gvU7yWS
p1w2qIjjtXMQ1gqTK4Gv9ou/Y2cVCTv++0Rvj9SjbSjP6IIdhCCp4RBPAyba
fcqMtn0r6O8OObjuL2jIGJ2rfEv/YGrFVab0wJ66CjZ5De6+UJSFlNh8DYCc
eOKDquv4cBMZ3SFKzFHAljRqqdRDYoKcr5w1GPVRcLW66MUwmV7Cv7UgYbS3
19EpKiceiaQHsxmsIRlyS2dYhf4QqpwMKCOiYuSYS5fbvfXJ4YxCFk0wLxgR
Nz8f9Sp2tMrb4Ump7yAnNC8sc2ZKLllumn/ZIY6uQm14lgA2le8Qv+mmZaiC
XRY+8hn1zVZ3fS6P4vi1MV9985u2S7fsZg72e+Ilqfi2pOrggu9nOmOW92nS
Qb22EL1m9SCnIc2G0a2AQ53ZjIW57skVwOlECU5O6GAMDcG/2b/5NI+aAoDH
83UT+2OnKX1dksi+gYbrJhitcjE4FdZ8N6si4vq6nwdTmrDKx0ji92aJMuVx
6+z9uzGYHNnntyLBYHzUnXCaSVMB+Avf/z+4QV6nDrfIXepIrIbDFL2ASVsF
fbi5DQyNU6VnRLZSaOX7I+b9HHi3VPZWEElFWJQh86il0uJCkMgYBHwglaY+
u0HPKiludDOl+o920B1F4FDvmHOwdwtY4pZJ6nrdMBlCndNCGP6qMqjbTJJD
PKW2snz8REzUpZdI4ElqKA+tVGpjTKe4Riauc4A/foIfI8+V+YLVQVi0dz3V
kbr6h6uNATJZ2CzMAyMx+NVYP0WJEQBO+IiOvSWg9Qj9WIZiiBp6GwRTElhL
rI7g2Bm1pEx5q0GGL58xs4cFdRS6wxeyBDdPdyURoi8Q5uRNK3MrrgZbbGzI
3P9oEeQ2MRHOU+QHkMEwA455375Q3HheUl3fdg38LJnSaaDF1g/3vYOaF9cK
ZIN7NtctsoPRLkvger08xFcNCiMdGRvWpszCrEKa53mudbTv/TwofiX/HnME
LkBItXp6Oj4dUcfqPASFqMvgvbKEWijERQr+jql7Kcc4qy584f8RFKau2X+H
KGIhkwbr3sLG0uvmC+/7gvkVwli8w1r0+Rk/8FV/kh+hQ6Sor7MYyE3EJw9U
TWfBXAMmR7esAKrNSOEl6aMiGO1k9Svo8nNJcHcDTnlZDUErOtcMdkuH11OZ
XUQzD6YWvHj67hiNosnxOu5iZoVhsfo4z58PbdWsKdJneA036Z1WpvW6iCYj
Wh3uLenXuYFYuxBS1rzAFsoejmrDKz+JwikhfaNIqi/Yt/nGUhrLtAP45J9i
jMYsMsm2JjMmuz4WnYIL/WfdxlwAMczswSbPJNwCQLHfxQYCf3ZveUcE2Zhc
dWdnub5wQr2DGJNLqQbkIAreAh2etmXRPNFiOWkY/mtBNMnpRI9vc1NB8BK4
VpqIHq5M7fa4kS0CkvcZBjXm9uN0dAI8EL3QBubVUXPzpuBjKauG2zW2F4TW
J8bE9YvQZWUszrY0dlg0ta6fynWGHe49OOT/YDkaLkMLZyE2fbEXVhpbiUXD
MVSC2+WfLdOY8p2/9Nuk4zusikQJbVzNTenkfNtfOoaE3hzaypn8r7K8fZAA
JrpCwgCFGd+RzOw57h69ww3ITFXRJ3d90wEMIBkCsrP2UJ2TCAp3XYmnvPdl
dYwdOsaGD1jNpDGyVv5TVA7Rysij8SqOI2uMzbeSmvB3CjXQ85Qwoo+R8zW+
gfp94f0rNq95OkTE7Mc9BQa/gQF70VPUzKIFn4/bCtX9ueXnp0+T2bj2wGmU
khPl8UyVCDoCdr23qkqLjFjWiN5EA8ohdNENqAs0wJ/ZDxFhxOLoexksgLtr
/J8vj3Dy7O8jRXVxvTSnt+lQ8plKbjrjZDOdNnVk1MxvWYD3iSHY1lQMJgpZ
/G0oVZ8FcS5IPdnu9DpZ2B8areXmKV08KzG0hmBQzl4F6ysdULKBT/b9TJsJ
i7XXjXYBg5wVNNIhJWjcqhzBXCZ+EttNhmpMXKhQps4W1BV5A7PPZT7btaFd
+MtWeQQpcooCvHsDnWHb8wMlWvBmrhmOvG7PrNUAPJ5BjbRZ67MNQwGgHpZv
pJltLivS3kAkVjgn6fcRCoSCZPdqhvjlaYj2h/d9bUbTHq/1RS6hwireFYLc
JHDIkBRFZxl6Qxzp7k3JoaJW5SEwhJjqIXOwHL6BUnsgEVLkhO0V6cvIBSLS
k/CVNBIMC558V85H/3oXIu2acAeHSAvV9Mom2ONmsskpbTa2DS13qfDxVGJv
Kkhf+P3ODFdz9+YI0sZ+Lft4+C+bEIg1BTbWrI9fmGHaJNEprknCFYuITDtT
4D/nFLmW/7wofzg0X28soL/HEGQ7envvSe7mFi4Dwe5O1vSVv8xA8jKnX5RP
hY/cg9IT+3l6w0ZYXc2jQJb0j0JkOLHrgPOukyzEnxeh0I0aYJ1K1TFacetf
MPaHBpVcWNvX5oAMkPLfdslI9bRvLHUcuZ+eChnLbDzRTsCuPcb5/LkeRsfR
+Fb2WP51HQ0p8GkcZZTZhp7UsAxcN0gUdR3fLnEoK1owha1zPcOsJ6o0xPv+
/6/gYHuAsXeuHlZHVCLXFp+WBJGJhXVQ9XelihNjjASnZtAoqF7k7m9k75To
1UPITSSeiS0gmq/wxoOulE6D6bHoBnlzhFBTmGVlFSbRQq3etMwr7kryBXYD
CWTLRFhAtEXBzP4sMmYlkrXhWKF6AiGrTjSg/2lK3oWIxWgp/L8paJz73lXF
WreKmuCMoYJAHwyPBFbWzM4n3qBvFTpdAS0yUgHDLQssOTGTzx13c67SHGLs
Mor7rS34t8B96rFCvYxvnKLlhPzsv00VLyLNSa5++bIDSMA6Cm6yNYbYivBJ
NdpcnQB7KIZbUfTfuhMhczqFTGNXnqqnCCA2Mih0Q8P+8wZnwwLvesfSBZR/
1n4ix5cBssVfOwJxaHsohxcddGPoRqq77t3+9XChunbnCpGDUGi77hvEjxVK
mbUvQQEDYpF6jdc9YrbR+UIUxcVmrWMahwEW+M6VNhMgxxev4c1ketCyNo/e
idtedQe3nwqp7y20fe1wRTPD5u1LoDaUI9vz+ypmh7q6aN1fQBBPdjFs0zAT
m34bnYC7ws8BD98QjHjeK2IY0edrOaH9Pd+SsdLZFsWVT/mzOnzusEaMztu3
lsuB0X6JVPzzjVzAenf9Fn4ZnjPadTFl/x5RNJSoFmF0TWheoHyCbggMVy2K
dKdqryAxdYHCvNnCIOW8SRGYmyZIimbdbzzJUwGpeeQy0gA7jAVVl/NjBu4D
PX50KlBKVTxQshQeytxkxqzMLTOWHMlWjCwa3vlGKyfbbjSq0cEy1I0Xuue1
ew5Aqdw+csvRgtN1REATcfPHILh+kG/dmWWOSSuST+IKKpg3MRmLD9EnrbFs
Fx4W7HxW8aZwiTypW5yLKThV/F46N0HdKt8ewfxWTGtppHKXbuF/RtUr9odU
PFLsAtoKeKFRscC1jOVt5K/dyI4yGPXCjjBaVT9oYhDrZ62gvjfFrJqtxdPh
P8q/6G55gL3X/yVk2PMLhpfl7FA+XyUcScV7lnt5GYWvnbistn+u1W/i/37w
mLv/cRAFc7Qr8PkDFNfddtdZRPpkpXitHpV/c7rXarKvVysf0rwkh/S6cNru
/GEkFDDBmv1BeNCndYW3NwDfpW/HGZ6ijX63ZL2JgqVxW3yYzqim8nKbTljY
myymSW57BV2gdq46H3rNQ9BeguKcbNLaFqC72DsDjYbFV4eBBVtNHjfAqqui
l/9YnYq+QxVji4gn7bjKkiQRDcpenBRNlMI5Wpz7csR8QXHUwyKBTQs4o4/V
Z6Gh+vw1T1jlC9EV5WtSC/BolcDNdshZdxNs3YL8CE4Nmv3/6JU4QiriQs5E
bl5GziQxgMKD14ZB9Dscyh9rpjgurbhMbcKVKkXisFPNUNoKZDNo9gljAS8W
z2c/EWRySET01GsQrR8lvC2O3d8mbP5VEpVmllDX2OK28x+27ZmVjO1BG5Rd
S/tR8qmS28WMfJHmurVhbJbb2QQlSGzVYV5fyj5HQNNuX0lJj1ECsGvidQfH
EzYZs09tp6HPIA1jrDeeI2/rFyFLUJL9axfD4EqcTNVHEYiQny7rAOP9DDbk
q1E41piPL/Aav9tqyVBjKWTnJNihYZ5eM3DGno9pPxqFhSei6fHsQ7hxPruy
rLQ4eG2iuhTE/8Jcy8pv0BP4J3Y3LLqR2bAvLyybDwD4Ce94utkZHSxBAilP
A81wLfsfN7X6xKrJs11sN6uy3SrC7nv6LlusGcjTLbvosiwUKDDEah2rEK/F
XoxQNh9cRWx+tqS1oubYHDorqfI4X5I4IXl8sh4eZlNRRw8szaq++UE/cl3I
OuVqN72E5bBA5zqqADMV67S1+UMPHxq56Z6CRIOk8QQNY/UzIUIgzmTOls0x
x3FshDGHXiMFNK9+SzqJScuJx/ccbIKJ04hCLL2E46G6frtDk7NQAmhC0RWQ
9t0EE9WsTHKY8th4TLq7swYiEZJiVsaCPTpn7E6X+mU1PFX5TtunLbWFC5kH
eg7heaczqSGSjxNUyoUKlCtfn3ZTMWHHr3Saqzg1UNUYhc9I4fHeXe99obXa
Q6gnvtMoEAnZ8pDcKgc+uH1PBE33kN4vDz02SLTj4+Pi0vGMx1b6VAgTMu6H
ZfSv0aJq9+q53XQq++UkXoxSwYREnUBXSmWGROrZnCBRswURU+hi0uMzJNZ4
M+jRNrRlmW0+HhD9i5ki/OSQV+gdd2pT09eWW03g8PppXDD862unhHZUs365
Io2ODe0BQ0ie23E1mGWXM5TlNudrbHH7Loh+1MaYhIgwIDjEkcgS5BCL1S/W
rLWGgn1GNQRXm/TavXaGbfwXLYPe/9725LVuhC9Ck2K+/KOqe3XNL/XqMWnb
Ah/3Q290Tw32Ljrwre1cbcHvArMXho60IHfAx4ZdJP2ZR6n+1jsKvGla7HxN
TP9f4UgBhFaYSo3WXxCtf8TnyoprZLEctl9o6iOjPGk55kcymoGTBA5jfH9a
v58LdGpHc9kgl9LMrE2Nzo+Wyv47BGqnQ/1Ox8FiSO0TdAvGneMqqmK5enR4
rmFG5oBjje5LLtsIJhiS/RLvp7mF/iNSa/kIERs4wx5YIB8oU0P07E++g5N5
tiWDsjhyGATkmhg9BXIYLYvi+4A8lBxgh5xyDG+wQUMTvIyv8zQSbS3MnL2s
zvtqH4lKtaegRzf0AzEgIdGlya4hJdZElxKsjkzpZUA5mvuVluU8ZjloM8it
6DbIeibn0sPO/8IfUgAwCtgtVbrXpRiIPw+KrbUB4mWXBVB0nY11Bi29bJCz
Pu+5yL9ey788CU00CauUyLGBQhRoSMBZdVRTExnuuxBkHsWsgpkb2KFQc5Wd
D2HsygO1xS5syNPdnoyCN8XhiEkgkotXpN4fKyUhvqBTpeR7oauHveoTa0g0
jXJqqcTa5yirockfZ8GtVBv7sWVILIB0lE7kJ89+WmJ8v9dlZvJ92aFVakz7
WQmXrtzuAiRhNRx1pTWvJ6Y8qyVeRKd5BSwn3uEFEQwX8l6R2f6v+QhQyrt5
6Z4tDb15vRcUwbmSc5YyG3Sw0iZTxbE1G3QFwlQ62yDqhnHTtu7O7WPMmZyw
WCTn3xeRA41fMHxKsO81GZwJe+qkcfwvR5AKKKVH5d0V19OY2t2/vjjvdgn7
Gi/7Swi4BSyYMD5F2O6MZlpM6KH5NWSYWMJFydp438Gb0ECNaq6vPgtS2x9u
C/mQs6Um6L9DhAR7gM1B1H6wyQ+chArwlYrYMBdsezvSt071dnTs9XTMxB+G
dngqLOeymJP6n5V7moHCv90aEQIksgio4sgXa4zhzZv/xL9odMPbTGrXE/vC
qDMmfUuttcBhcFAvEzTM68vOYEBovKa+brcDxA+lxjN9tGaj7nfMihl8/zk+
VQysdKbxCQKpK4dc6lMUQKE3K8W2AM63mi7OgplfGQ8c85gy31tPsGyW0dmE
goLxDh0n+AcUEWdW/FHGp8tbFcWqiibv0j+I2DwRBnxA6t4GO8W3K8dlJ4d3
iBaYLrndRInHKXtN2W2AxTO8glgnuBG3tQBuive9PdH11QCCkgWK6TcjTaDF
9Z/6e18ztcnrkzdAENYBuC14mbEUJdoZGxCgQLEtOjx1cH+MtUyOD3QaQWPa
h7CFXtXFKBrEM/bFrA+IdEipwEqEmnepNANvrpShfJSEArXxzso67PgXRCJ1
TWuAuZYUrAaFYCeny+WddcEoTgXDVHlM4wd+EP30iOvP3BpssBivdBw480ek
gpXjhrxzHGSP1wY4yGgXp7ZdX6BOA8AJ/7a0Mq3xFtKFL909xUuECpDOShol
ZJILLdrVsMrB6Z/fs19xsp5WSEbJNrYjleXFubBSQq7I2vJOjYMRhDk+Jv8d
xC0e331Fh4l/7FOm5t7E1WFXceETD0fiizP3amxZohH7lUYtGr94OO8k4zTC
FB5uFakIb82XCv+kKlJJkduBOKLbbu90AP5PBNb8HCfP9hy+hHMf8lGjMlOq
OVBpayVZeKKWp77cIdL/GO6m3uBMijtvEasGhwPCf22XzKOoYVMbgFSgPxlW
WnUASShSujZqg/QqIN3LKT52qYrt8r5HAMLD4n5iUNpJ7CwT6YMaGTvzNoy9
CiOQfASYfwztV1h6UTE7sgO5xgF8+22lUeZzUoXrtjl7QxUZu71cIKqjdp0e
hns/bx0d0mwZ66rkvP0B2pXwEhaPaH8/Q7CkEvFmJ/BF/aFkW5SQdSj+dTXQ
fkXGq5K5472jsVf+0kjw9M9d5Ir4xtO0OJvF0LhRwk3rkJ3oosLdIwQbpjLx
vmk+L8FgKhOcShziBsH/AsFpqQwgP+IOvDn3jBfHuhR0x8pHFlaTSj8qqliT
1UsozZAiv9lsFEDWN4putYAjyRjnj9qZrAwBRMNNvYKaaytqdTAxCWBeO5A3
g8vOvyB2bRia9CvCHXhfk7haEzLy8LaiF/P6Y4DjMro3y0f33iqZPKX3vcaI
r+4ERivDv2it6iNY8fss/3HPDpqvj4KDd7Ho94REwYVeZqXb+doSUjgOB5Pq
WSzkoMerfjbdbKs7kq8OD7c6Wpeh79nXdWsfSit+WCKy7gwDGx56s+gAXtxP
cDESuIHFyW3p1c8tAiZ6+y/0gaeaQ+Oq0Y4TyHzxTBvH9Q26a2DYjSpLerMe
fy3j7srFLFre5GHtpxmIdp5x+muCbs5ThC+rFh1vbUzppVaK2RfphnIMvAHu
hFhbctC1JkllR4NZ37YpZd+73VK+KxnPnHAVRtK5gGRN8Z/ncjcXMmH0meMS
isA9sfm2ho+mhjObnBD3C7S8BCQdI+3/Cm36vQRhNA+DV9ycoVYkh8MMy7yk
bW70yl5b392cvItu0qHzJdeGyhBEihcsS+1Edq1R4B1/nYCsJxR+2DoiHLJb
hs4Zl2rJENqah6CSEzYwco6ORh0p8jH+7Y+UHqFFb7sMJqAzbogp59aX6Osk
uU/L0TFVFhAdlnFZMb3WoJKvi+HZ/bb7Ba8ku65po/8XUTzL2F89M/gcK3g9
aG9vFDqfIKzcQimxu26e/eFbBY2VQn1ATNvDozqoLUgVfnZAUQ1qRkM94foX
RBfpXdFqiW58OQWQ3BZSkriBG2VQi8zmkNZqeXwd5iP51X6bWAARx15fHbaY
Cfrg7lpIukynbbKwJvTMby97jMGk3byLu9hdjHMrPXX91Tab9/VVadZ9YGv0
q88rvPDqMpvNNihwsX1A4/GWKF0IVhWvcLYgcv0pii42RxxzjzSmi3z0EmM3
iVLNSFWFxn70/KLSj3RRr1jAl4C2U0r4uUjEJjV3xTv1cifpr0ndCZZXwudW
tYxCCIW2ELXVHY94bIF+YtGjyUS1J1MghOcCpIUv4W4se9nIfoCSv89AzzuC
caElaQn1iu8ZlWWkbB10LT0ixtGfd5dt8HzcpfFI6+/e9k4t5Be+9b0xQU2+
kCEDuSuJVIDxj9lnnGYGYAcQz7zQ3qRhMf+LhU4Vv/8yEy4b5uu0nMSdEmEi
iK4L36i24yHzM8RPJxiv70fSJZ3ISrPazZs8pEw19A66pYNvgth+De/zImzf
s4zqrz8NCmWbNagzvkSYA1fyLrRqNol120iMYO9nphw3FmHozjUdsXm2APTM
q9S0XNO35P1pGRgmI+ZbkbljR4b3exxx00+WwjRGA6+yDT8zbxLrrX9n/ytM
yr+eucP8O6kH0fDf7umslrPyUVwHld+Ks9ljnf/kjOj/s6crgRDs3+68ADwf
B7kO2VHWulAIaEq/B1BiixHbazt2+cZE6BTjULvY5VxOO8ibfVPa+cXyYPNv
QTzCd9JN5xneWw/1m+cPSIIR/3Wr2MYBQkfRTvTvXlK6yREdv4qvWgH2V/tR
iXmi9T/9yJjdoaolkAJWTJb7jq5gvsnSWo2wjV+sYOEQveAWO0goQta8O/7X
ubz6cutOkCOMCh2mL1/cwteUJQ03hGivs+OaJxofBTN7M6HM6NpA5H/hmFs8
lqdxTP+MD2UHFmBtLji0RsmcI/id4TFai8aj3V6cs7CHRa495hIdchcNFi85
GJsWc3CpiICHaapYNUJOuaZAj2iSYd5BByIn35uzXHMPc3gBqQx7g6baKuJq
TnDPEu2WlnX/3RgCEAaVwLOtplz7RPO9jE/7+4WmVJjmv5/Da3JBd6CJ3Tce
C8dQO6hy0pVI6UOSvbiv6cE7PRMp0n1EmpQtGrTDdDX652aQrpThY4HL2HRb
hPsMUWUPOdtfdOStmVKRiwKExhJHuADbqtmH/4qW88uCX5p3IjdZYEv20o8o
ybAxx8Xe5YY/93VqQp9uPYxESGDbQTfxa++zUhYzbgUt0HEyurZ390EqLLeX
gqxV5Xew7DNPmEqp51ljH+ndiDq6Rv4HmoY3kdYQ+DJ8dojRBLq1bNthp4yX
DV9QDcF3NUoWG7ubCuzm2HE+hI+g5iUh/DKcXkSB4ESDqd+EOGHlnIaZAfxH
e7OKzoNc6Nzz3J2cVB4FJvFPp6Q0vKxJo+aghJheRm4gM2recf33fszRe1xX
PvWWWL5ON8egAUviQQ2tce7uBca/P2p50u3ea8P0bsllM1wpCLxC+01JXr2F
fpFtgCe4uEOKfO6seEtg1Sw3vKHs6G8wO4sEqyoaE2uWYnMS/7+ZOJtNpw5C
I2rbQ2NCzz7DUa/IgCg0NHeMRY49jqL4ndLE/HVaUzivlXvHC4LZRmkM/pXW
XJNvejbCgtVuRq9ENPmBwoEDCNauaaOiSLJpOSzVurlRVzp+FeTe/z3idGSO
0WyUlA4mhIM44CHck3whS3o/adhDnnQE/0MS4j+TQNVqNTVDLuTn/VQDxZuw
NoevBkfUkrnbWSRY9ahKiKgg/bbsIBiyO3vttTayEY9TR6uckbkum58U1sjc
BdJaivgp0uReMrJhEiTu9VLeEYtovw1eHKmR6//zvIVEJ2cyxzmB2ax4e2/w
kP/NXBBr48vXL8CduYmAWGFk386M8PD44STg3UYsOr7FGdDHxBFeI+5hcej6
OAI2Sdfkpo5XmZU02V3H3oejf7cNOG+Vgg243J88hqIf0xC56pYExrcyn4XV
+ipgPULQvLlaxLFkHXhohQZGhuHSD4MdtqRytfaFxnUO94wb/ZEnvYow9LhX
+llAviSaipYGkknbz6hKQl12MNzqHgNZDRQXD/8kVANzXF7ZyGzNyt2irZg4
VoXmY+rr1LyWxGh9ihYBiw6QOfig6zHqjpe/vktGq2+cJ8CJcUQaOlHpDecH
lFA8oMCdz9W+Dn2y/G8k9PVtxCdqnb8bZw4yG5aWmV3+IC8ywHhS4P5nWdb1
xn7Xtpcvipo3qyRQ8HJ568yNLcjgstvnO9czplWhkicdZ+kxdEfgivLFd1l6
c04ITqdHffvLyIZkUIv3nt2qsv+9g5EHRJ5RVAUCiCylNNLRO+zhXJOFd3P4
tO7+vi/vBaXT9B2oBpdnsMmK/34NHgVGBB6i8ujx7V+Qe5NBBAasp/l2arTM
3pBBKwQzCHjQNhXVWFupKPNQttC+VWI+PNLzbtcr1ysVyBxTrameg6AMDtgx
R0K16iMV1EDYdFCYFoiA685v7yuZscyADgvWlsebBgS+ZS/SDafe6438ozUy
KPJY4AxWsCy6WGOIKf/gxcWb4w+uI8vnhcxyuFpMGcX4mVOEnpQWoxrqNg1a
ZBFAV4gVbpEZsR3pdTsAEicpLrHneKPTU/PhtxPAJnR+lBFRCmilapJn58dC
HyQNhGX714ywerV4imUd7Tv3UUR/lwnEUoslXUpeyKk/eO4AJDvvHt2Q0zwo
C9SHY317ku7HO1MoMOW6EZaLkJJwiB909ar76364ivfdDWy+w1Jnz5O6sqKm
mMNERNtIy79INRwSC+gS2wFcPpCyxovVcDeyMxfNhMRKtDDDoJznc4mrmF7Z
N17ETOxjExbapCM+7+YnB4x3SfkU0oWYtMKr88982tff/DqgfepVgrHDZ7Xh
oJn78fp8/9XSpQ10GuerDTLVqXcHxXl24m/ag5jCbQpJoRKFZgbWeoCIlMHX
46x8lbtx/e8oldPiH/YI25i/0roApzozOv6GUEciuPCbqVT/yP4to+4fztY3
QU+ODiHnTSeEJ/5vSZyFLcMAYjvc/IFq+nUGM9/tzCjPd70QPmFB9EVG6ldU
HRv0yP19TM2gP/92+miyffYhTVSwNuANmynkwc/ViswRElTF66O047RtxYqp
yuKBv7asTe3S/1hC9V3BEekgGNm5bReTLASMzStOaCHepEBPfdJvlN5PdLSU
fURapoOuZ5MsfsHVl6Pd3N65lWXbAwGS6jW9ufiYBrgqGabaS/SzWMt7T5xM
rvqWNH2uX8VIQI9IL7NN4v6Wz6lTg4xTsqSnqYq++YXh6mSgdF13C6xqP4u1
dIYPAWGnEB8p4HQlfhjrvMoKpdoBkfXUTXFKme3IPPNrxc+LUSgg/FE89mxO
uxVdcT4B4YBn27b1YpnHkfmQVjz+3768iMYYaUuAhTIGF9SwTeXSEI4pRdAN
5YW+PIDqgzpfV0XxxJvLjOmTS8nMtO89IZ04zuYo4ycVveH1GP7je9Uk8RQJ
uCBxYCareuQGMqvvEOW4icuKUdJvmjpyDD1ohpDaWnqRq+exofwTHhJzDecb
qg4lASD/f+X97zcKLQmSI1akA3dqHoRdguvN0cO7CusbAQd5KTAgEMBZ7ctn
6TZe9q96paj99GDna3vyPObFF5FjMwb9tiT6pBOdPpY1u491sjRIyBfJwEi7
QGx9teRNwQhmd3G4pIVuxNF9PE2MoRQ30IfiM4paJTl1/ck79MJZt84V0TLP
Jr+2/+g63J4nLRhTuSaP7tTlby5BQ9gXvyERPMTHhLTOgWmUWq188Bgb7dkP
KHLnMtJwisQIzBmQ3fxSfqzlAl5NqyVnowaE5Nb/Qvx0y9nM7T0hUWeSOn8/
Vj2vSqhMJUYxm3P7A1vNQmffrun4fcpditPoqNfvIQ85VfUpeIZ7QsKY4vHR
Bvfp0N0nlGpZfMW/DVJjB/RNuABawxV6S9f5WBMJQ278KNhW0jMafYSayCuE
W4ItW6aVBdN3dynQHJwg0YiIkcgmm1PN5vqa5q7UL34Am6wrNl0GC+F24WcX
nWSdPhAX9kr7V8qz1lPcG4SF7Waf0Fjso8IPofNqRHR700WcRBz5aE4ruqPo
XfoMGZn6djggBmzZohAb5sC1TXARVTgUoduUwzhNAvz77TIublxxmlUBoShO
ndEWxdpXGkXs5Y59y1KiY5tFRYjfj0HwiN9LBIJVBtHNkJpnuVpEeiP/ahCl
f4qaXmU//65VUZEAkGRkHpzl5xojakHEISCSmi6TB5Yfds0H3QIfSCqkURqB
hZFVVH4BbRzbCGaNBVwVsdyV5EcvuhBf3cMp7aqO8i7J9lpCohaAqnaMRghR
uOTVn8k87q4+HVgdCco247L0mI+LpDvSxlf08R22DA5Hb0E+3aOR+VVF5Jgq
AoxQGNDVHHCQCdjik02+pu6yqE6ibhiZrC1g0oPrdwzPMPM3y0FzEyu5CSTn
Yu1V6OYYOw3iOgIcxZCY6PaV4EQkB/k7klu0uc/Gei9vEe6UI0/IuTptfpM2
224U9V/FTHjvd/BU/CDU+hOifi/QOOaD5534yqlFAlOeVewosIWaElg7HhnO
whcLAie5uO9mu8cVjYGNhaOvqsluvlbq4AWKlakywa8IUhZjk9pelAWIrJbw
Z9loMWPneVCAOy+H8zDQw+lbSGPUzFQ4hd7Z10I3Dj2YZyrkaQbsy7ud/fTq
7FqTcpqHbTIOFfODPZqFYnQwXhAdCea3Bwcwy1XzgyurGYL3ibB4JvHweSio
azV58epqdOiBObwHznFh2JUfd5uthkhOajGwq3k2LwFr9zg0bC2PrxzloCUG
SonMGQTN7p5BFvK4dKXCHmBICCJIkpgOIr+rv0rGF04AOwL5yohBg1EON8AX
MwyXkrMe74cIxKnaaLEoaq/32gtOVaosVFyqvCLooHFnF/LWHB3GYxTuRvN4
eApTmg8VRty1P8CqB0ipUE/0fpHy2AUGfmQSsMvkygLYEDCplDE5YbsGqXSU
8jGzfkhGrhdOnZFP86dcCvjzhDlRgobFUU7g4XbPlAWYJV5gzu09BgRZE+A5
mk/5FwRsjMu+fFqyJcp2LZvMm8fkRPVtDn+Z7UTAXd515L6hgHn1AyOdjvZn
fw9X1IkYg69HYZGWCwKouzphMH9zfHKzj1DTt/eK0jA3It/xiQQDYU6bzVsc
XeFBPRIHGOAs1fFRIj+1oJxDIazstfJ7IxtCetYlvC4znmkSiy5E490p5nJ+
Y9Wa+uXCG2DHAiU0imcMSJ5HmC3BYsGysghtn+GpuNeO0UiFqhH1wBKRd+Gn
2sSRQ0FM2DMgD+FHIAfP35SnwRO6eFiJK5VU3tgWmtUqGm/g6kQFkJxvmE3K
vQoGfvSzzOZO5XLemLjdBwPRP1s+P0H+2fnFff4fFHQ9WvHLFlxqSzQ2jxD2
eHLLv18Xx/srcOXAhEZszwPcEB351SRY9wHgGuo02gy0P2tco+IXcCULRagn
goMNFOSQZSRg3LLjpdiH0X91l2YXSnVnBPTkT+TxakxasEewRyImwvwcxUVm
yMD5HTGSElj+x2JDXwknhpPJ1sm+94okkpLgIAL9SEQfbqsWMG0DKZBa6IMs
qMSq3SdrPwJ/dloKJRl1Vg217XPha/momO0MXyMIWBg2Q0B2leGVUTZJB8yB
/Szh9YS3OjG5aQUl2NC0AocXlCvn5QffeUN2KyqIFbuwDalAAKBIZttH0Wt6
F95OMiKcV5kh/z3Mxb306xGwhH2cM2bVW5hMBVUsJ3bk20y9vlWZv28Xm8Uw
nJR0iqshQgZWLyrM50wtKJbZKF7NoJRIVEOH2W2tlH4auRVv1lV1d9Nuf2M5
l7tvD9+GQIoVSOOfksquq5ekKoYcTwyImJ8oRzaJlWkT1dGk02vt1pF3qSQ1
7oNAKb7mxlQSyjSnX/tymiilrFkllfTrpnc+zZqJuqkY4JlkD0Td1gEdrR4J
XQoxI9ytIkMftz0r0a/zBxgO4w+AoEoAcJv4WJkGdMeeOmhce2YLALAj6433
5Y0+4jBUswGCsrquVFRpXS/r/tdfPJaV/PtdCB/3EFFnKksZ2j+CctLTKlPk
NZOlnJAbwzkwa2Efj1VzddT2elGKJwJMUrSufG4zJZGt5oylMOxi9PZwWsmU
hIlhbxYWMsed4YwhUsNb+Cq1DrlejWAE3V/RFOebn5RXfeZy8OdgqZ0cJ0ZR
PpOvMRfDkQ5y51OEqgWzJbzRX/KVQKoy5QISHM9m2+GPFs1CLLlotsfE1wgc
gxdW2KfXzGU5Sl+H8qtbLhd8RIrUA2pCbS6n94dPGlAzio9QwUYB6J+7kuoX
mdNi5s4yOehkqg5NiIniiygpS5URnQRCgmnyb1YdQpOUgXeWFJCl355nDPc/
Jt4b8XlTIxDsrc2smzE79i61SZQD+cCWFPK6Tkz7A1mPnqW8H/MGS+1urUDR
L3Amf/RMHPr85xdYvuEZQGoCzO4EvMdR45ml+1JqW2DnXtG9tr9ByALbhY1r
4UVs/4wiLfh9EDqgEpGHkKYocJH3ShNMG+m1Vj8mgfHR5XQh6EN98p9gTm3u
BVRujoTtgfNEw8ZM/YcFC4rNJMTeDs/HLizHTJA3EgDgSh9a3luQ/Hl7JTxd
24s5WsMcabXISx+obrZReOGUp9V8jl7dA2S9fST2rWm7hrAyx5zbx5XqxD5v
B2vk9k/5lDgmVcMs4tNHJaikB51n5FQgqyxbOR9ISPfmn4RlWMYD2K9E2/HJ
kkv3eAN8n5nEU7VNlV2Sn1lv7y5duZzy3awfBzsV2d4Dm9dUOO3hAStJMk+M
zgry2g20LR0OuoxezCFvHxDR+Y9H/RA+PFtBcyH1WH9+WxWr6H8xEr8kXCjM
lZXax7mOTbOtgp0LSq4ljrHSSkQA+1YgkxlBLsecwhWEo8H4SF9Pk2z8ZF1v
0ztzzoOkGeduY0w2VCefSPR26wzvtVUHBCPqrdl7v95p2pYa79EuZWK2SP35
HFh2kVXNodgV0XPGbFz9oDLZf1HhBZ3sJcGA8cfiwoZl30IXWqP1VANukpjK
PeygH7PxtITqujRosb+3t1t6onA1G+u1LGg4gK7ZYKkJDl2GlOvSJGiD70ai
hAQ4x8+dph10MsZKMzv2UnSlT4ubrIC+z4dsKdMnxzQxTAqEbd+dX+izQ0JV
5Y12R6IMWSzBHvcv0hCz6lPi9T8wiVWwktNpRaKrIcw+Y7LrdTVBbIe4UMUi
0Rav+eWFsP2t7Yy9X6+n5nlwJkhXzx9j1TISWU+uNYCUvP4pDzas1lEP1SRh
7DB5U91i7hVKPfjx5kCG8vR+/G1NcyryxKYVNKLoO39FcjkUR0Aep3Aflcip
5Vmb9Irxt1eX/lH+dyrHMq9dylH6CFgkLvqaqS3BK+poCrYuM+X9gNT0tH+C
jmaYFMCLeZ/QhJhnNt7PFRrkKzxhHGxMdoyyN4sAcGihjn1fYYEXu0HAJNZf
otxuqEQUrxwR2/QKogx3ZV4cmkhEfLBOKIOKuhoJcFs1GZv0YplIW9NtUHhu
zQv3kDB8fXzCnMbb9Wr8FCsoCADWFQvddjRFEL1QIPYAN8Q1GA4AWyAJmF+0
JRFroYVlIRLa1+iMGVAgPUvI4cv6til6HjYpPyLKUjBBiFgyNSny7mtaq/5I
QHwcRvjL7jG+KQrXrOKs6sFBYsRMg0wL7Y1B8cFmi5VszXklE89uKTVxXmXi
NaorXgVOOM5hfMc4NT2tKwgkU0O4nTJBEKO5YP/BSd7JTFKh8IFYxgutlCIg
Ljb0tETUMZHjdd0FUKHaeQRpmnDj7l9Lv1Xp7LlaRPM71smxZO026NHOCkuk
OqzuRNVqd5+lTJJHmjkLYf4jG/pyI0aVCoFf8mOuRi9CakPXimfc5O0iEiNu
IrHnlOGJ+8YlZ8QwHfaNyqz8G8iC18ugxVZ4TnkoTPfTbYDE7YUemoe5O3Kg
lnPrr2qit0m+wE812nQ/qWQRNgtXo0HKj66nr0ljQECjKBIhYdnjewP+8ZtF
fWDEEyo7lJGqA22ro1wINRsiZjcByu+kEawf4gOLZgZFa1waCfS1XiYQchIG
GPB99U0gmMKWQq5hW6Ng4HME7wVMdNrktqtKJDta02qzhozHtKzB8w+MrGRs
eK7lBp59IrHfzImYL98OZza6xI1qpj6DOGPXr0hBINVER8ZnEHqceq458e20
TTX7DUfuLgQfa2GcOIj0gWIwzw3j9OhShVWIPlpqHnJNgDa54gWLiUkLJWFJ
tAWuuRrgoJP1yaddtCLXb511O5TE0fXY4JkYhNpCxAzJcLkp1ptBtBVu2w8k
2rINkooXo+ZDH7d0Jytz4GtT6gSy8I1E5gllhz9BF/6VFDWwLxgzo2/2th8B
Yk0SIPueN7KhuiK9DWtnDc1nb847hNHDnmWTm+seg3tV0xklDT3vojHYo8S7
zviqkgHsrwv0NKtr8DLwZUmGQHkLBBUjBmWTGjuAyyckKnaPP5zH0mrTa5hA
RuxZ+yQ2xpwJz6bt5m0Sdhf7C//GcnV913ChT5JX0k1ow+shEy5Yzpv8NEo5
BPIlPWUDP2K1NjcNFJTOYQcVWVPSdRzU13JDMBtVfxBDYYyTZ8HDOeKP1VEr
vhAZlIebLxvzCc8mTidFFXsAiqNbOfz9YaaZbnC+XgnHr7nN+FGFSFajPgYQ
vMhBH+UK7WYpK4fMbf8Am/Uw5kaT+5Rdrht5LoaZO/IflPwn9ktfoM/uA9f7
DwLeHCq6Ks/YqRO76eBC+HrnZIfGz/rIK/3k3V8qntc8VbG12YOHVB8EeMMy
TrVyUeKQLEnxvO5U+1CaTE/wao/TnU8RPEYhKmG5uTcsfQmNGGlmtMrspovX
G3EO0GLz89IntaV3rjT1CA92aZxDCdMJQY+PD/V450o3XQmadzaaV3IYaQHF
whNNGpNUjReDSGLPECdU7KPMEa0rWk+21aNoeHiXGpCePB2OrrsdlJu+4Fry
mzEIK8l2Pe9R/H+aHyUkvXl+BnI6DJdBpqCgRYH0hSTaK45/4Nj/gXPTxiEQ
R81frLaE5VOD1OfzOHw+kzYomEv6kd2s8dKmER6nczgseduf8ISAJkdWbWvj
m0u24Mwp3SPlpzPUzDT8hdqZNPorET6Pbk6wSaVYOIxPyoxKDjW1JZdrWo75
cTxWwOCeQaxB6GDk7HP9KmSm6wl0W6u4ErMcAv/ZkAZBpYeg1ymbebf1iAwu
8hLy4eFa+VeBrP9AF6H8rISdZ11FmUgnY7KcfmRZA+kob+j0xrKJc1BQOLVS
DifHNS2QfU15hxCRu8Gu+9B2+6HaDhdscWm82Pv18ZL8wlY9NeTzkgq++m7I
j//ULo3vOBWpMVfLeN3YwDADPNFcsicL4gzA7lpbgNw4b6RpY2hRgbF+/9vp
ujQ82R0meQJNYGv355gWsFqAnmFnbnNpBvnE4vTxDFcqfQsbdz7UfjOoqsnt
cvnBWBblbDaG2wevveDyIUgJ4sBXF3RMzEAFPbSU6SS/Deu1ypQwkFLUvoHJ
XG102PzH6BxflY18ZtLPj+mt0/gM6d4Ww6kWyz6bsJ564L5aL1D/W0tvUpq1
Tx9Rku0gsVyJb/9pIywSVwEsAk77BYiwj25EqGbXVfStbIupcAnL87w7bAg/
dGXo0k9q4j9BckSblV9kRSUHAKs7Ag1UKRNsG8OtQYcrITTbufOxfXfbmvaS
64QUFG5nSlNTPs9bG42fB5PJnA4Q6yrJ72cZHkgC6hIWphGMXK6S2o0PDEzS
J7zMjSi58/5bVU1c6LvaHquzgI+PtNAVAorCfoQZQGfuwaonMKB3lDoM45tk
ztP94E46hHB5MicQcM78Jwexv43qcr8sLaHcJKWX7YX1WwKkLwOthQmmgY1F
sbctdR6KSJToCFZrHRYP5G/2O5uyEv2a/0tVSLMAJHxlx9n0awdTyMUMyt5m
zMw/P3zeEsVdmLHyuzj4KLB8DmJvNgkaSlJfSptRLV/ErzXqxhT/rzfdxlUz
0NmaB+N+Qds/q8oL4yHs5lAvvudOHqEcTFeR3XP16q08HDNg9bWAj8m1vkTI
9eVmlFdjq48BddOUPlp4Q5eCMD0aDJozjdfQVnDOJNBOfxlBiAgtCDlVIKEs
GU3ZfN0DhEgIJWz3mrIiCZ+jjRiE6RGiJsuWgchx/OwZiurXig9RMHEafxPN
/OQgfNylebH733Pz0J3+FvT7E6USdqQoCUW3tXTqcy9CPauXbch6ODpg6D8P
U0nX2zrExasARhPZV2K8luRzgQj0yQyVhZS1kcnUbhsGfqhQdaf44f/aVGOt
8+ITjrEWwc52ePBYnEkG/89+m9hkygJOyWF8/9/AMoL3IAwqfRdZlF+tCTrp
+A71Gthe4UfzXtT3uMH/ll+dz1zOVw/kajTRf5fFuurvEw+274jd7XnhfQpZ
5K7wn+MzqygLDffFMORHdcIkXDx7zs9pCOj6LmCFFIGCc+Xuu1wZflgBMJXu
U3U9mh1+SXbGEzT8rjYvMM8Ar0O/m5BSq0PJUi0u7+kAxkOcrAF/Ys3FsGBp
dSKkzC8Cbf+SLtoYpX7KAmE1v6gEJILBsHwDbBy+T3GNIjGQ96+vORt+g/Ci
o8E6snJqh4xq/6kuoONjrXlKC+KRTZ7ckPHSqm8X48TXf6bfeE3fgNEUOzMD
K32N2XmXD0HODxaR8qNh4bdq+Ii9RlwDVcqK3kZABSXn/EydMfHZxs1z0pMj
35s8TAcKzGKbFnRugs3n7ZPZxFypVW17JsYTEiwJai9xp2JkG4FAKO34hfhm
lp0b1RVy54CnYODrPds2lGdb8CWMJkgPrQ5DnetL6PJVx51DbBC7fUZqaaQl
dhsrgb0SSQcnh//6PRgOS5DXsemcwZNTIsXiU1IiIIgJ/VA22pZC6RPH0uLq
aAdaIQ/5eWz8ud4STIzD1d1VY2desqSg5mch+hzPTCIsXvClC1P13ilgsgrb
dSZgH4bLcqdHssfmBvKYAnz6d5jCjdd8ASM3hukhXtZMhdXYfqq/sWYAg0da
3UkRIZi0ju1dupWEJ9kMBwPEcJYHZz9PC/dedcont27xa0QVVIHYE+y6U/PH
eOjhO8dzUHo7I2EuZHOLrLP1sBzF4PUYVYNC+yQ5Hm4ZP7XTBXGqJqiqac+3
sZZoqcfYzqFGJqcBqsJsOD5xSiZ7KkF9h36YiOnD7j2o2DhG/nE4ckkr3TiC
fFshcMgoqMs6ZZaIHs9ugQP4yAkfDfvNNjfz68ZnWVso94haWEg73CHi+pzu
WM7GQBpwu+S6QvZgsGyj58DOLs4bT+07mKXAStgHzo0vZkuzdR4wCSA70i6q
yKCOoeLzMQhsT05dVaMHn2Bpnirk1/1OdsBhPNWjkM4SNNQDNQLvqT8n6f0n
lux5DMMKmUjPVl1vUlkVJ6eRKaOsMaiVcNPCJF6p3e8xqk483lg5RPqDiiR9
XSFtDTbqJ5vSzzhaOYKA8wwBkKNgknHs9RvFTGM5fcwy169o9VwUL0W3pJwL
IUamUMTe/w8fQd/7ZmpqALKYaZmlelq/Hp85j5Vu237365yV/FS5OuL+1BvP
gASLrU/cqP5Bt/WP0LxDiL4AV6EE/vPkCaAwdc81d44fKswS0+OkvbPeZLuf
Tthhb2VAij/fgRbRKSuNxgK6jlVG7wr7jh/SYC0F9HKx+gcBkKwEFmqRcJzZ
8LwprAjX9B9Jtpatm0+j2WYnlDZFkz5rH0jzfKbsPEmcTAlw10+tkO9i6lBl
BrwBBfmoz1RJrMXfD+5vtEREE0p8SP0eq2cIrsDxiRcFuXWDLo3HrWij/onW
ZlgJZniHhUDVNF96AyFSFp8pKjbcm5DPD+2PZrOyAPbK8uMhqm+DbaK5pJu9
3+OvaOeLuHq0Y4Xl26LGIQiGNanbcWUed9kz0WPPaaqbZjrrbRFLU8RfamBH
NgV5Gv8wVQxMpKusFkDXhnO6H5vDrmTIB/y4pUUJZHP4FAWeUlncUfVgfqVg
FCjp1ucVo8e8J7xcDmUl/NYhZje14RZVDVZ/Zi8pwxqcrQNhk1kefN2Tmaj0
mBRHkCqGSAusAJ0ESJbCo3l8oYJE+dgscQyzyj4p0y1kdk3yT+VOZ54T/zwn
pDo4rrlPvuUCQLqIO6iN7PDjVdhXroeD/2G8jA/HZKka3lEN7eSlAXGYF5xV
at0Kh27ghPhBS9D56Vh/YU2q9j9ner7m5+oDnzB95K218wCfs+S+0GLMiiD3
BQ1JmUziDYmLSvcJKg/gdFJKt9NKz0ixE9U0gpM4w0bW/JZnhrk/Q4DmXIlg
08TGsyARJJxzGjV4T0qtRm2IRnEL1iGbeR2d/csJ0Cq8UwLNk/XsKCEM9EwJ
Pwo3vYwwL3ruy0mPhgCn176BCZbvE4j4JK/Wy67P5La60lzySkb4hzxbVRuZ
bHBanf4Ok4wnrDPXMcvRYuaiOV+L6XBWTpcS78LeeWm+sFyyfWpPvhHJYA7+
WRxCaUmgJMh9f7qnyki7UfH9urmrB32lhfm07gGHVsBppVnmTvCxhMkDMreQ
diCc2w065tkJTIRXEEENmVpQKxRRI54Ul+00l6tB9BMa7KLT938C+2OU6f1/
uqb792NbV7XkTjDVwrV8zIyC8H/XSQsAoPPTiT8jlvf26dMFTVjPBfk1Bckw
Mcml4LQt8QBFD9A10tI2COb8tgwMt2g3roIG/D4mwiszVKgTpaZav/HLdCnQ
RLW4JwZnY9xXie9xJjRXR+SFOk4iKzdl2S7TW1mH79IYHkUahthfSkvrTBME
jue5sUIRYe1f+dZvQu9fblN3kQKzhaBmXCDZKvh/vKjvHwcC1mwK3GgZshtE
VDUScQYvet8UO2/lBSBIxAH+dw8NnVabkItUHeZglGdTSivvQJzjOYSKVeSl
5itTmpB34u3WD+yytqIldIe9odYHCfjBCWh0M2KmvkFnD6JhQtAVDuDjMYXp
EkBDzo1uxb7L+kIKZ7u7nt+vDqo0jpSf1yWRybHY//dQd8TxSByUeTEzUJBC
ivbPAvstLzWYBxgwTqcGwz4H7UQi8TdRFA0sv0D0YZ5LLZ1k40jXC5Y/TMG2
ihLF+Emaf3yDbiuckgYf1s/ypdFhFTNxhB8SJePA/xlbDAWrVp5xDDOxsBHz
N2ydlLqDyu66YHoI6Fh7y0FLmppnTHPB21CY8ZXNcD+Atxq7+FNW0EH+3399
xBvR8i4v7jZdlRIuOxvUXSUJDKvBJD4wdlRp9apelOg9xbjJe2DNkDp4VrIi
K/wBTv8Hm1BBS7SgRKTAHrZgshBcxPZF3Soib5NGJFGGKmD+3AjQfZpdsFw8
kRQhZLaxbWQK5kkwA0WEko0XOBDkSBOIEO3lliCKugjSvNf5AGmxvz3xWBB2
0CDUeaTCffFhN6R6ez0t6UkHb+NE11mapc5i8TgAbQUhY8kWZv4dDtc6tRji
1f96tsdYW7+OGkriMoQ3qPhAwEo0nmmPhCiX/MUQsKN5sTF3B7pUd2SqaBw1
SM9A3g88e+lKje+mbbH8saKPviYujZSgfV+QMT2yNmG3oQ4kqPc2FyiiefP9
7x2XKDjL3i/aGO5Ws7SFtFOD+ClSKINrr+0YMX6lSP8hNAs+kH5Tn+3wGjko
bP8HG6ofZTICw09J/+SnRYzoo/lwKzUSJbOLZEDFGOGVOFX/FIBHZcLDZlQF
5Y/QFkX4RE6XMczilHgVFG7ILPMpzE5Gmz3dkZm8NRFhW169T/QtFanLHqCy
h0sYZ0a8mpV6KRLG3DFbqbxdV87DZqoXcslz2ODFOYEA8O95UOJ3tTgnmOU+
bgIncN/lm2kIH/tcxR/8B3NdTIEc/QKpEYpToCaEVI5zt7Q3jiHQOH5t7Hej
5ZQYBhgxR0NVvezOQ3yW4adHQFMmEkdhAp+iAF97mTVQgl/C4WK4Q4AvHqAr
fDWXHJzAEr9kit8wqOInGS9+q6vGBNvRIcR7bbLSAlJwcMj/DcTJ8KL9WudE
t2ync/Zg07b7jENW/gNeiwBDrUV9E+HAFkHH1yTNSiNz74oFZVIlardZSBUV
nrOI5+DeG+KOW8D5yyFKESVftIGeVhCTDDjT9yEfylVjX+4TfSpe257E5c4p
Zicn/Ep1Aj6+9OIxa7IuOmEDDsgSBk/31+NRaLqzrjngaALzxtXpvvmqx4Uc
4oaIH8Bbaz0FAK9lx8Ym6wTrksdJl3ZO+hNUO5+twGZMdPx5z76W3u5C9vqI
+jKwt4PSRIdUgl4FqVq1DRTZRSOnUKajKj44XJcpF/6rsoZfvq0qnjWW5kut
ttDgtIzXrhQllW4XOyKmwKf6OzAIaVhY+76eJZXqi//EYJ0zNwEHWdLkBjz8
jCuvfXDVq9iOTObb5opu0Uim4x3vbGT/1k7ivRQPXbbMMF2dTz2sMrIZobDT
UH8dRWYAJztDoYtqWUgXtiNbBtXcunQo4eDb45GTUvS7nfeGmSH2XidnMNuM
+Le2og060VNSc6RV2KuXF/AF1PL4cecLs8C8IWi1+Jhi5rntxqsWOwr+EZuR
EYa7JkEJfD9RSflZs4+p7gqgG/M3gVO+HDJEvQbzRx4Bqm7T+KnL9fKDgf1o
i9GQ6T3HP8O/b/x9bl8QopeNUQDc0eIWANwETAdgOYwwC7r+LBPHAR3NK/hq
DprxurrT9J2m1RhHy1T2SDKDslf0v8sy0WeYtCwuOODRBCQDJbB3e01KtTGt
c1VB+s1UqVkgiGtWez04tuieKS9jXCDGiFfDxIzEOXxvSDJ9EsQZOM7gkAZX
E3PLbZRjoRm/VXOU+U2LPt/EmN63wWwGONNm1MaaMAxQu8qqrFQKVIHHEEEo
AVcPQrAbsOFy7zsrxCrDi6ti7cmkAuniltNg5HranotXIEgR087NOLQu4d8I
ZK8CgBEUEhv5OGrA1ivWB1QYeNxWgVnUb5i2hoptAjrcPvyMT6twdEkfjlKA
1JqHF7wrNo7DYgO2losUY+wxUPVSeOh12maNCVMQPJ6KswsQ7AtGVFp9lxRF
5+P8UJGCU8xzFZtVqPTAW86VGUx4ClaiuR/8zGxnhcC+NLL8aKaKKEvnDHZP
hqjNBMZJ6PjKAkHxEou45bTtJUVmEy9RZD/3Z1PZOyflHZAKml+bfyzboYUl
UyZcgBxLNyjuwNoJRDUBvWEOzVwVJOywwXg9/EIGX/zL+LqG4zI6g4uW6HEZ
0myXlPYy5NnUzzhYLEbCyXN3ulYVsZVPzg7soZnfD0skmdem66W9C2/i0Os+
iTh2cux679OxY7j733XZKtj90N/wElzYrNtzSTqdxXcit9b4Hh9AOgnInHvy
w/e+wzXpFt96X5qRru3pUtT0Gc4w6j2zLXp5zcQRNL9EeX4TjsGZzo4ZJ0qh
ZMO14F7EkRNk5+7509EJABWzR4EosHrTRK5e/hRo5iNKE/9Kwd5stfFwTrHv
eSdavlYLmbDdoo24lM8OT6CxYy9PPE6pzDfEQM/3Sg/zx9WdWbm+nXh2B9ce
AcIQcc1qliqYshlVpX9ABE/kRJFww17cHCz2S2QCpLzoUn3s04PCXAUEF1og
2vCgGVRKxtkMao7jIsn7GLAophi3VmsposNPV0UkDs8vgxGwFB+N6KF4m3wp
y0cJY1xwCz4DH1ro56mOe9BI4f1BoXAw10eFt77fwqq3ik/5Jhles/WO+kmj
LD1gcOc6rFO6fOk0mEbMEV5U9D/0L0pNh9T9E9rMvvV/sGwMnJTgAIi3wc8H
WFomXvMQC1NqSA+bpAHJy8trljTm8XS/WCGPAGwe+3TDwHF0wVWrlovrNxUv
04ZVwsNJNejyw4aO5WOTj7UsMtsINUZ6ekaxiNwmysQSI+TB9MuFMfkp53mM
Dq9HJX+ZozqCMc+VE39EJEEoWZFy8DBgLIzPK//JbWfsz6Zog4afx8IG9jzr
R3uqkOOoTYZDRVDAMq91B84wpulxk6/cs49HnU5sNGBRNqtxY5icVpoXuWq2
vY+VBegkH2JVRkjLsqNiVHYgyeg21WmABPXVUYxbgE2MN2Y6IPkchf9XNX2q
48uANDgWA6mCt/X0QUbZjTjPgHIjk7GbW+U8dHVZjQRxTE/9d2gpue7NutNf
IAtMOr9bj4mGhZhq9cjqoqlKHM3mIU0ufVuiQ/1Y0uir86oXCC8j0iwKEkLy
/NSLKOfQmREO1nOGnogqgiCSSqO7si4ye1vATQ+zgsz0GCxK9W1mrG8Lhp2O
wy0S8fl3IvqZ31qPSeSjONmv5LmZUAFskdF5bWDfof0AkKArN7g1qFj64p/B
STi2CHNbZHc0/1lgQ3lPpw+G3Yq4ZD9uRET0TatyWzVFayGrsQ0aEqkpgt3H
Yh0R3/NF4a0UBrSzKFi5N6SB/oZivLakTFzDEe6y0BCiKz479aHp49BHsI8g
zbFF/dfJFxKov7NPoFxtdPyn7wLYDvGliMIDQhQRQLHKVyYvZmnfGyH//5sm
d6CK0c2xp8euHqIdNB9B9YO5JpnS9SPh2v9sO/tCVnkiYT3KdjYWVJqqDNvI
h1+7qJkGLzthiPO/g2dY6qvLbbrW77+E8mKHV2K8m45oycolm64F5HxH9z8N
lB87iDU9Ud/SGO4vanIdvQmfkEH7oepWIXK1ugRCdtDtQISTKK93kOhCt3xL
wEsAUhShmbB/GnkzDTA5Vu136ACEvEp7ypNc6gcVV1vahQyXcQUe0LLpHroC
jfpqxbjDD/dFX5zgg0gyuNT9H+JexAbfUChI5Ytq8xTyvfwCcD+09p5wLxKu
5Qjk7vPRp6rBaVZBscT7/eCu1khrYjAYOATmtoBA9doVh6/u2fX0vJs46fT8
jHTgWvJB4g+alC+A9yvK0//dyFdryksQs4RPGPrE8vtkgV6rgeP5+YnEhSCk
xIVrnznJ5xfCOj4xmCUYJQZ9c38V9QDqdTnnbq5NZgmBaJgdoyMbdxb2XHR3
u30JsM+3Pwu2yFKfZdVMKCa85LSb+TblaY1XfV1Q25R6lWKNRn/zMki8qCIX
PB1WRM6Z3lgkY5zGOwk+kLnPNIXISacRF1YZjMoaMmoIQKdqfIW911Vne9Mh
1qr228kiRajU5gIU6L+a5EAmJ4eiaNGFvsHLr0VQWF8iPbYjIPIirFDKfeuB
mshUGjqDLsos3eJOd8OiOM8R6+8EQnreRQwoNmLvg4GkRPc+mI7vvmv7BxOX
fGrZGQIP4mh/bus6EOnrp44iwJnHoJ9wydc8SfEfh2xfxdplAOhhVQjYtF37
MmpuJPmOY3m2BSXw66JoSyx8RhVuoAgc7eBSRyU9Xi8JuYOE6ndYZ2bNMMVL
J9b8OcKTU1AD7Vxyeybi5dhqSf4NXVqU3l/GvilxJR24ZS4qIxrQCAd5MtS/
V7bKaI0ty7G/WNFbxLbaaDKz9zyBjpdhFmeoBrWGJIlXsZNhqPHfoI7q9D4K
22Bg6yAoOhZIkT3NU+oUD4qtoPJeyYdZ7BhO2nDz51eUk6OQupZkbHuqgoei
CByNHVi5z8ArwN9WJkwdpp88KXNF79OxItptgBVVqhCiFZ2HzV7NW4tZ3aX7
9DxXxwc8W6Dh468MRieSR+bm8ffPxGM0bxzyH8hhqlk3G0Xdwkjt9CiJNUdc
SuTYVR14IjH4INdwjRB7Sg4QHkXENMedUZmeV0wOTbWg3gectXdADo5ulD40
V5q+Kxp0A64yPXCsq5Zcjmsrjgfdk1RgOoDfruW8UbxLDiLHzc/IGcg12Vwh
spRzmP8DkDKpAP+lmXDOJHklglm+Ug5ehxpUca+59tsDPpmsyfTjbQw6tRd4
/yEO+nHF8dCCxYBjGraBLH8oscWQAfrOlEvO3GHQGfmIOrkJzRobCOxkpjM4
iT1sICZ5DwlpflaV17FeCK5uL6KhPpVGpr8lGOS8BMOMv5Rh176moNYT+rpT
AGmpGzqeimjKjwD43IBePaX/penwb5O8lu5c03sJIeDuw4EBz10uQuQTjlHx
aDgLBKZIqvXouyPyc0q8ojXW0lSxUMZ9tb3JPsEYZi54XZXBpe5f3TruV/as
FSVKI4Lv7MzddkQsEQqoIIA+kk6rNUHQhC3AlS6lzcfnabAlDlYKuKb4n3bZ
0tueULJpffXJ2f/dztk9TbeQl7sZ5dBizX9SRDW6Y77mD+PNkhGnBI66QBMC
Z845BCsccP59+2a4KwG+hRnOjORH3xfVG5tl1UtM+KENNshjqnL67sL3/0tx
2KeZY+MJZ5Gxx2340Bgyrt90DGKRgxg0c2meiACqmoGpLxqpqGQB6CAEZ6V8
Zucj/+Tg/oSFKbo1DM72uGpi6q7q8IyemOEVI6NA95+vntaycR/UGobqr5hE
+3kb9HX0i2HRusXg8etbdUkQyigx6AV45XmM2Uia9+FU4/I3OCwX4W0zzHp2
CNEuyk1P3kFfz4kD20jQuaA2qzMUcM4ubi0HtY4tNmpS9dxY56K/4mmoCQpu
n+znP7Mynfkp2KI6ZZ/Miog45QH9OpOHaWnRADhCaER9SkYHOcBbJwPlkm2J
gt0GBnHOCYcBrF0E8ofuDv5tABQSdKLjP+BUDZBItOsUbCv6XdstiVg42Au/
8Vv47y9ivQ5wELpNX3pC266d/00hxk8WlLZiGRbZX2wn4jY9VlDq6fLg6C0h
cs3hbI3PtiUS8FLcFwTgw7TeKBMZYWVu7aTNKnSKOzT8Qkyz6/6okKP8lgm6
5UCIEosYjZ26Q81eVYKHdW3rYdY8DOXq+TaD9kkbiU1Pms6V9LfNNHEUCvtW
cICV92H5HUYUzPXxchny+3N0faFjLcKsA4sc6oPjCcTpCVy61KtE9ZtUVEBT
K21YrYFDV+ZcQX9mNKZvGKC7HcIw1iyqPoSjVEIb+CJFwb5f+b8VellyqxgX
9I3k4L1aVFUx6McOkmXQeEvZl3DhKRJjNM6vw+EQxbJ5hXQU941VAFDyftzZ
oSVRbLN0dUNTIs38UfqLuN3T2O7CHE/E6sZNT0tNno4vCIKgdx8L7Arx0d1K
ipvEVl3YxnZIo86TqXMMoS0DV47aLNCtm2qE+T0s8QB7WGwLNqKkxZ1xG8pU
kz1c+iAvUR10QzuuqP+aLlU4fDnMYxBaFEmA2JvgRRsyIBlpjZOgKGoqS0cA
9XZVgf64cVpYPFsSeYOY18UUdSndHFOs1VhLtVxajkD2Gaq5Ru5XzKYRODxy
JyUlI6H0YoP9jPcs5uYs2/fTR1+7qQBwhEa1JqO9tz3aW108kxCFsQokSzR6
usRTgRme8/yyY9LldMSaqI7R+S1wZXvwpVoT4rYYcJ2jEPi5SOd/wW/Giilx
rit9CfKeP20/XSqtUCuT+YJYvAriigJxW4noAtSa+6ZQJg1/ajMmXZ4vvFu4
GWy0zTS+SeUPOBDrOE2+w079FVM5QslqY1qIvbtIygJjMVAA+i1MkvDPlBR/
yKRhxUcvtFbgjlfl3kvzQDCEtmNKPnBfoaLv00USdGpNXEww3nqgI7KGXqIi
F2JKxHMdHGVCgDPhLgWFy21ot2eZdgzcdIDkyIG4DHaYuzEUgq8UDnYmSYoS
zfBcjnLXtO4C90nHPZS4oknBika3nLF7svjFRm9HuRcpn17MGcyOJRLufXEa
ZjzinK2Q1UQ98jSGka+b5Le81oFLL8bGYrf6in2ajT37GcEsl41950MuaOfH
aZH9oVY6pcOiksEbOS4dzLXWG/Tm+qvmIFX3oLT6Lzs8GccZJScLvJweuVP5
3zx/PDBxZSH7w18i8XW7bnTGaFHo1776ow2HNBh2yRejy8NPoEDbiCy6Bjsv
X2IwdWvOQnGlqBysZhSAxyx/HJUR1gekIkoSR1x55rsRBII5SVtE65vY2/JF
ZPbbrQyaD4zp4iMnUSGy+9pSyQJZ08S9YzNTJOXc/3+yGkdayun8dHNczfu7
8aZ/XOVZTPlvpRtrBj3zq0+eLgh+hrcvOdpMv2aTfLVzQe97GEbgVd0CtSm/
HeDKi3QNcFAZZ8D3iEbbzeODABTwR/tDieVF9BQOCZWg3i2TBPEfZqf1jZe9
/Mksu7hDpUfFNovmqdBYmwi5CBr3SoiWeTytY/JNLT/qFGVlxxUQV8gcLnGM
CsfjlE2KYIWGJeAnFXfNJpKSeNn8x/4YDrbX/tx6WY88Sp3gKyey5hK4JEwU
6ODL3/Ww/rV1oh62s/XBr4WapxM9OpWce2vvOJd1ITplzbe36AZX+l1rwG4U
CKhdkZ9Xkt134OXSTFX4eNvFxQ0aYHpeYsduzOwbpEyqT1Tjm9QYZEmvooi4
Qv5s429iAhvvs6o8kCaXehfztGV27v6IckvBDoUnaFGJJrTqsIQpIjEFeSF/
thDSoErC2PFWxuCbpQnNBJZ9rvwY1QOl7t15MQfAkYfj4pejGU3HTtxR5GuD
NUUq7hat7mO7V9rASDiqWVdF8rg6dDRIy9+313esAiF7NUtv91zw1zROmBbq
vHbDLlV7Y/w/wUUj2wkWc1EFyfBNwgvdqvM6+8y1QaHDgmSq6A1XLN7Ksx/h
zqMBd0JlWFbrjbUSbmGMs71142mx+dd0lcAIl2WfKDWzNKxse5wRKqDeZZ63
xGzwlzGqrOVifO+04VFDsxJJ8dZqsr84bsQ6ZOLw3m1sfvYYr+Ky4ekU9wFD
MuYotvymDVzGV0hxuU8bXolGnuHw3QwSzKAxFZSoZWqEHvOw6NFX+P8yxCJX
oSZzduuYLmsB5ZKPoGNge3CviqVt7X/vfVa1DJbZWbHz70R1HK720/2z3GuX
xeYS4O6GCxBcbS7jMxG9ZPcseL8FX6eUAoezq9EYJk1klHV9E3puPXn06NNB
haAzJ1bAN9i/qdQKO6dyb+RY8dRc9CyrmqkbrSdvCBXlPyBsWfeJz2eSHAc3
F1ob6UU0P1hOwTEhE3wQh7KYwiQqpBYNIaRyuB+ilhepNVCBX90MREmsMYa/
3ikySHnv7+CoDzsQAj22MhS8N0fcBE3qdRcQn7fbAJp6jVrhSJA2gepvakwN
y0PNWQXiYut8sDKXlwk1Qv1d7w6SMGQxsRT+NrVCwAO/V0LdqatxihuzdLY6
jfEi7s4FuVBTpbtX8wdIMagnv/LDQXQnJ0yQHQZXAvX6u+w2sx/LDDAgWXwW
Q8axuCa5MiJy2VnpevJ2qVRgdWFhUrXdlPaIpzqwbd05zUAmIaZqQNKi3rQa
HlSU4uPCybJ87NSljZpgviW8X1wwB2p2GCCxzE/+XUj3WUC3BmzhCrkHX9F7
huOZraGGwrhZFb/9j8U6vqlL/h8giGE8AXeb6YAIMmseawFFoorH4QwWyZyW
HZ5uAW53f6eMkMJ0bUKeXH/cUWu+B8Z+8w0eDvzCZAyhlQSSXLxxQXUtzToq
0abUcSpcxG06jggsEoFPnAy74t1hknVRi4ykq4p6flxydTbIVK6SltAjURX+
Xzm1myFfCE9jdLKyLB6AQ2R3FRsVOQGRm3I9JcEl4aFk+8HY2mT5FEBOPdIP
Ri86LYDKThLaVXEZ/v8Np0X/Ber9D5X2TAIY4tiYQL4MZtSXyUEk+bv5jP9D
+FBbbzKWgLwQAtwM4faIxTm9a1GsqOta3pd19+dDBkhPP7KOW/ZE0ayW/0Hk
LV0EkUoZkqDRZZWNGR6+k0e6UzwdCVsdYRKvUPCkl/5+iF0d69T0snYjrOqv
OMNpJ1l3YFu3W933CqSJQUGq9kfPzTnrWZobL/axzqZSpa7LxVkKFfgwMb7h
PFLo1UZ3NZhzeqIAhkePL5ttVp8dzWpUN6l0NnCJdETSJCPYWQx0IJ1INY+i
cVf263bb/wqniKEZmrs6gbhTHWfRdh4xFbU6yvkw0vlclPXnHc9TdDZ/eXQy
I3IGXc/Xghmak2AkGCJBJ1k8xo625VYBBEbaSOkPm63m7yW77d1wTDg2aOfZ
TFMJ4Ndhnc7iJ2IO4L5n7zxWVS+31Bj4B7uiQV59BSnmt2aLN7E5ESMRIyK8
NiAJxmcQkB7OmF4lVqXXyHwEFrxllcaZm3PSJWPHXx7CPNXJSmBdsAiPsNKK
pO2OEBVt/xglVtFXBk+rfxGqj6fiNMQrv7OpVP6zBc3Efman1J+PdUWWm4FH
0VSeDzblP2Z1Y8h2j2nWxvKD96FtqnINaoLffYOB13kkAqLdSTxzPWkedKEa
ta9wC6fkracXR2mv52OfZ/L8BXiQHyyPERZpSnLnzdRBtxNc2nwh9fkpRsxr
GELfSMBU9sdRep7ygnqxtzWBV6ZxvBvWz4osrGNLYhdQ5FTfL+mxhL9YJS1m
LSMmemP7fLA471jjfF4WZMYk73EYeaDAdfO8p0VqUp+D0QniuWb3XXkNgJZj
uLnftCqCttTpDC724C78Dm52fp1BKFeLjgG6pf4nrzVCWiKJMyU+IUyIMgXu
Dl3DEIVDUOasqaoYZ5YHe95BQMqmlIGzKByDEheYWdj7EhGYl95cQ5YsmexQ
qOVcXOzP05VytCrCD/13d+ia8fKzAWt9upP2Nmc34l5JZX0S+mt6ZcxEoIq8
j4A4KKvbrhxNkqZTj+T8YoQUJLGqwZ5+2DgLsm4vrZYmOjBdRCGdeTETFYgM
fp751edfXIYu85mguPBmOGMRtCnr8IgXGR/U2a5sZYL1DSnzfdPriyc75SUp
yWgF4RefTxytxSaj/b+gABU9z4u2Ptr7XG07hhdawqUzhDsDiZar0GUW7RCL
ADV6mRXVw1SSxwE+kT9nhD8KCL1kyDyEEl26iKA6lhx9MBcdQ0kxUrwW3/FU
eAnIL9iVk8ciICWOohb0DQCn1nolY7uBsYMv33eeWX24x82oB9/E+b/poj3a
DZyPwHZwh83htt+/o2htdB7X2apgyAIQ6tzBci7YNa9/Eywimf6o3ldIvWPb
oNDoehk1To3ypXkb7Wcp81c/NCYDdtU0S2iAhJvICMIXMG7x/hoMGCxHp4Nn
GyNvDH3SRqQ+UTK20oazw5uSxkynm6koBbvpuet3GS997hShfYWDt5wd3l37
tOFFNGSIKO2uldRoHAzX02Nqcf7Z+lodZSq7GS4jQ1ULmR4PKQeT9AUrRCZ3
HD+a2BtChWlO1Ic15HS+lW+IvRqn6fm36L24RIYQkJqewHV1mzCxKuqMBQrd
8KSi+5y3rjEEsv+1jA23Se5W2MJc+MpwabQ1aRS1k4naHbuAXw3JzJKHi+Jq
33p0poeF0Ohv3M7M5LC3VCE0kGc8I9aqOUvgjEiXHaJeSOwLQyrf3Q0ZZU1M
1r2nOP9B4LflgMC58qeiefAux2TXfOtEKgVJtty3nQyycu68rlEZTDs3GmBK
jJriTcD5mTAaW0o0MVPlu+da7UjMceXHKQR62Qw81c1XSlz6U30pmPiDlG4s
zNR9for0JoRacDk3B4hIUt5wfEwyh/vUdR7O0YEPTX11qx7nxkY0DHqBWiNP
C2DNephRoWrcOTsdWql/XS6N0DRRiLGFrJQ1mg3A0WT1eJ+Dsgs0S13NCgGH
QTcRxvMPqllr/bLTLZS3PPVif8wdJGwBlq8lWZijanVGRFxv79fZ5xkU3VWN
+E/SdrN7lsSnFV15/RPqZtF8dyh5WdGdE+M6dUtt/7SBcZNH4xpAh1IwxFVj
Rc3mni1sIsSETwOviOYB6sjETiUNOEJS7ER5Gl26YTSEpkfeO+j6wpPsi3hH
hnmspQyW/Xbf88LOsOEIctqo0fyD79b7kFUpRATsBhR5P4RZN31K50Q/8OK3
KutKIy0d/Vdaoh0rBlMDbkNOBrEaRPNKRzqknAf4DVXseSje+PNLVv/z70AO
j7B7mt7P3F0GNANbkf571HziejOGoUArLYXnhHtV6oF3+4LBF9P0pm+sUFwI
nDLixaGC1kWvx+JDprAfHxGbj/WIwclBSZmEi1/Lvi12KEwZiZU1TnDwJJIN
UPD/PJEspyVv91j1C9LoAWB2tx4xJMVtympvTRV1H5+bwQyQmCcL7D8diazX
weOY25B6ajvoTyZDTRopaIgVoWSjeHBdCdM4OQ5x5X9VBfwb5fkKyp8vrIp1
qQif/7IaXxBUrp8zCbA+XPpLJl9H+5ieBkc+NgJ1SFTYRQC3+XkokV/XPntN
RLYtJ8ghSNqqp90T0TYRiE0fo2zY76i+/jZkgQhsJrjRZhbD9rzLvRJ/ApZ9
gKWZG+x30FIM9y3bLp7wZyM7ei8Qd04GPOG/FAF+W3bNQ2+nMt7cHqhgFXw3
ab2VFR/j1a9AUjVtqocgxl32vkyP8bYW9U5HM11yUQHKhTrSuJnGA1Jq8QNd
uwq/3Z6GKm4ozBIicl87G5VX3vYRdtzwI9R79f2HMF1aploWNDoERXmEneXC
wF3aeVR0WKjnTYjEbSYGI3amm8XMDKcLt2Q0ZGcxR5vMX462b5XnMJj9+0g8
BHjcd4zau2se4rY+dH4jzUUEAliuwtWSBVQUCSEbz1ZGge+29izxFpOwk4Qm
C5Hj0fB3GlfdEwvrO27b87HgdPU0x2/qVeYiTPcqdaVXPbAE9uCRLB1WyRzs
d5y/DIUI667Ky0/g5SHsbmjpw72lar+sGxYLmjsm1AVrkwMSrsjnCjwIgPOX
yOS1kIZU1XRztd9xH00+P+MhyuLhDPBUO/PwDcfBdDLxjDItm7UzZwMdb/YC
eqBRbzV+azG20hjQL8saf/A/PNmKBM4XFIT0g3lSDRPJOt3OjI2/sp4pmkI9
6PamyU3MQNvRHaFrDsbD5wehuna19p22Lg9qQEkTL6m7BeYb6pQB+utFJ0iU
QPAq4iZu7W5TAw7na+kAuYbmWiF8ZMVUi9y3Ebjy4SGUAlruK/YOaNb6LtIY
3TyPX7G6geaCsU0F2Y79lrv8/on36z4VntBXldCiyGMsokITO9rZnkfzP8L3
R0gZT9V8G0bBmPcUYJ1lohITuBsAVOZwiMPpYFcjUAh+if0j8ECFQe+wH0Ly
QEgjxIscU7nBSIGk/Ps7jQdEsGbPmER4RsumfBRAFUGFRsPdgzLvCWvBMjn8
Ae3aAiSe0g2fACP+c+QDMD9ycHfSJMhS8SgS+TRJT+ye+xipDwSaYtymO85H
yuPbyFmJarps1XW1gRJPWz/MVdXAhR0RJRvWNh+KkCracpBSKtTheEgoCOy3
0Muof/sl/ZI5V+fj1csjQXcv14SD6LNlJbn+I6YX6G/WGfxkSS3Bn3xU+6ji
nlPr1CDg7BxMeRvxmsYzbd6mzibKrdN9Q9NUjGO4gzJ3CcRIbSOBcrAFLtOX
SQY8Ac4EtoEm+7gRUjFyj5mpJwbpjOrI6rqiewbqO8mwNtYbz7UcHyXOlWwg
zZ3wCoAPMai/tvl/cJ1qUFf9ZyX+FC4YJ0+sA9AN16AVupPgt4r3uwBaAPRd
6ml3kPsC263Iuwu4n2TNk7YrlXpyOneAht0O1E4u3xHHtjCY2KTpoWEddcZ9
Wo316+GGMTpeAPUxdpVY9ttGska7fTnrEDjfSVWYO6eTN3OtFMt8GkhuVuxH
1deiw8jmZ86WOzKrgqWCgOveyI3XUp/swWk7BAc8shaU8vl5I6le9s7+hIbC
lTs/lU0Qwxhamm4069ExvNzAYSlS0Tf7B1a2/uJIEGsuHqLaFpqZvTk5gf0U
SSjlaQiUrR38iRIM7gJZY8gzgDmcxhhlgG5JFVEHYS0MR9tg3TQbdl2m2MoU
x8AxhDEXneaXnftoRKruQul7pL7c/6SJcZe8cWc+Pf443ADTNrMWbuhe/6La
7vWOMCcX68sIOv0NHdzaRElP0+ps7mf5mxCeFZr7cTGReyU44VmKGsOuMawn
y3Yu+nTUbz5Fw+4aYyguEylAE0fjTXw4HivHs7Vy4vAAQ6OsqnsfXHcKMsn/
R7k1q6z60ywLR9woeMH5TUaxcEGzVYGKBE2TzhhYMb/AbeHMy3WjsxRzw++A
sagkQ+mpa1h1opY6DvHBtJo/QSA1cyQuPhwwv/loeSPWsq2M+CFLczC3DlFa
23DPErR8rY1F3E/wb1TlmudiIALlQrQyIF3gNo6YR1Tr+OntGRprIkICJLDz
2bzm0Jj/Y3H5qoKLvujmiigqwTybXJSaHvG9HXXdouNyYLCOB6oAhCFZc6tq
vi+RsRw6lVaWAV06+g3mStDUgMEv+70UMgPAONXEztrs6EeYq3q5+JmyilkF
1uk1LIYcCYWW6dHnVUH6S6/mwsYN3QuphKvR+GGSi/O9uWDYmHkBwRyELSjg
mrBarTi/Hco3PWr7xCqVCjIV+JMBeG54rFlREAa0MyekZvbQl0GDGIusOSjI
itYwfJZxBt1kpD7NNJK4tCjTopXfAK/t9iDHbAja2LRFPyQ57uXrTNtZtTFp
+n9dVCxOzGhYEsRxijpoJRKCCpxXLH9ZeKtzUHPF7ZysNTJPWVUKp/IMtPCH
yuFLzhCRcRO4PhRpzIAtHvEXI0E4Rjwnual8JtY8mXFeHzveICDOHv0QENQl
oCyep3LqAJ5ZZfD5dlPgYuMonRGDwsEkUwFQdy/UQ5uk0L7U0nx4BH2MwWCz
nmzL3NvJnEM2pjooL2VhHT9bdyVbQla0TUgqlVqjM9nHpou6AjrzDNS94FwG
KRlXIrww7+A99jmCz61WucWWXtAR+cidQttA0TxQ76cSkGu3i1izW4m4HrGN
6DD96+4NYKHUr10cJKj62KETr6FiLWOb/UP7Di6xjXvZc1J9NOrCl9jv9Gap
ECDMK1Ucc+ePge5ydApDglnVVs2IzQcD+YP8PpMfv4sxMOlxw3ScAA2vwUVk
NXi1cQjaEZtG4GJbOBg4wX6JLE9ltlXrEAY6kkEPHi2VQYhntf5tm7QA5idI
rHR+eA1BEKJT01clVs/ibUZm00EDn+lzJYhQuR7kN2cAcPv5sUXDU9/1Rdln
F+p8uN9NGLaqYqeMeBweR4wr8eA3lmDnBxPD6JwTaxTYR9palCBNs/+nBl9b
SP00xJsiL5Y8kN+6F9XBButTAOvpW2G0rH0gm84yXPL5sHA6ZMQa/JVolGVC
HaEWu/hMwZ13Eb7YeKALTC4I6JMKKkM9Bv7rPY1qz74mRomq17U13PoNgWgh
bj5ach31oQ8tA1HV/qNWGPKFKteTaE81KsgzR5MziUc8e/MCixtFvj2kBszY
g/RJ0ZPTWWycSL+t1dAEYa8bWZht+sT9EoBgghcNxk/oIkYN9brlfQhbmDk7
haiIRaYJ0AnGY4Jm1sH8LfXiVZoMS3ZsOwJSLxSS8LxWJc7kpZzBe7M70o5p
sqOaKG8PYdJwW1zCw2dtker0XY7YSauzFE9mTftL+gVDnZKy9lN04774ToFt
unfjhI/8DK3las4goJIO47NvMkMPgkrSt6jONdl29+v6k96jN3hGjkIrt/pL
/9MXXsRfwngky4Zsewn813Pdg2ED4bl2n+ggvxeZ/cDJaKIKCXCBy55D5jMZ
jGTlnu7oQqSnM6pSsHsJc4b1C4kL2yZUZXOhyHkYvwdRh0VTW2I/i3bFiXte
fpTNeHdZ6wFWbBwLr0c7EOLhSlH1ojrqqXyAFxXIX0b/jRiiszZctN5vAdZ+
wnmum5JqHO0JY6HnuRJCjeS4fnnxLwIsBekNMLbyTIU3YU0Y3skayyn5HAPF
n1+pX2t0xWT3BRx7y9f7yZ7nxZrqQb9E6wbYz/9BNfpPQM6m/WSLOG70N68+
UptK8Us4r/5BOZDgAqBOS80U1+Jdj5Kr0cZPFHd1hrf5zzQa1ASYvegdqO7J
up/ZNx8/Jvu5xF7NKecW2zK4lQVtTQqh/s83ZOaH2NNmaLb8YdbXRCAXmW7B
BnNH6eJ8nAMQhznQTcCoeUrR++t/mqIR5oY0L23UcOkU6MSy8bhnN4OEmvRH
oliiMp66XpORFuznTnjhQacGr8QJ2fm/Wf3es7BRJvBV88wZm9kKqhPi5iOu
HnQiB8c8tE7k8m+SBAXesr5XdphlW7LNBZsTKdcl/aqZ1o2SvIGCuaRR2RWf
EoPhHlwR58P6O6m0EhdJhvBVIjh3pTppN1vjYkm53fKoW6uKMQW/MqdDsz1e
WUjOdZYLHJkyJlK9mLinFDvJfL9lbEisZ9Zohfml9tswIne1/lIeC417ljmD
VYziOAVYXe1W4HeXIDa5j4xNNhdLZCUc35axBWqkn8SuuyihEFivbdPDEEBg
dUzFsRr3PW/8jree8JbzVfTlxqwXwbpf/qMrwxiehvgRBnSMergPrBIfecqo
4y3sfS5VwxVWVjHmcs/c+nzad51MzlUb4BO7vQOIsIFR2QIvS39A5iVFI8pI
reSOBc4XCWTMK2PBxHCXUo/km3fx0HrD4mqXFUwo9YgPrUTDPzBT5Bp5092Y
NzhizvIr+iAAsy1K/rax4gnGztGI/uoqA0c5FrYgzFrZ2TtlZ0Q2D+Mpi2CK
AeK04o96HSBw3+XbG1KtO/7feHapm/H4yLRZ6NP0BRtCOFsDUyfdr/hmb5Im
6bPetCzDYhsuhlj677zj2lQxVkGCDUYGb2QwCCBfRNgUKvjJESMhMNBkEqcK
jrMgnrwl3b3V1iPXgnZ8g1MFd3UUxEysu/CL976WSJujlhluM+422pBc9Duw
M1jmPGSIByvu7lP8sZiGTY0FIMa+lQkQprI3AB4F3zSHVfpnh8up7ps8sGKx
BH/sSzlxg1On8T6pi57bvKsllMR0l6NJ1NzQfFh6xz3+QCfnSiX6elj74k3Q
dzGBrfufhcoJlldUJOZHQiCdgm00UKtlA8TvTDWb/+oYq/HML1yvSjW/EC2c
ds1ulw/KFFXs1NDMFn8bjDNNhiP4dYdAxoOGmWfGj51Im9tjVV+Jfy3pMbF6
eVbdWVYkEzRfA5NYRiJNDhxgT8wTu9EGj1MLY2Sb0yF9RR0l4lW+Kgk1I3G1
2hn5pEB1EYzB8gKpTxLoJl8mEVdEOhjQDXaqhwZIxzHzFFFoQFfU9F8slVKe
UOc4W3XXLimQCidvLfCXof2S1HMNRzeNBaDPipxQLhY2sPi9IIwquQvUwxpg
9NkF7W8qiK5v44pFDenttKvTL23l2RuN2HBuWvwbQAgEJiVlYodZTVePFkh0
88VJCsqSOg7OBfyzk3A4gASLHK95fPDa/zSEWYyehsQ7sbHWvavubynHR+VL
ODYlxD4e1mXvx1kCU5X66VWuPC3h2OclJQ9v9VVBP489v7Jxdwc1rTOBTknl
2jDZk0qsb/IfNMPi3m/OO8E6tmRvmDIdVepq4Yhkbquy/RPm3/BOsHl1AKJE
zHs7xyRZsNTMH4H8IPIiqBk4p1y0UwIKz8qUfvHTQW4flfhZQzzaY/QH33wi
p33BgmeNwIeJCauY2EFq43yW7Ds9dHbj3q39iL+bFMNe+U3vP9xy3+7s5nRw
upot+bGr1QFW36LAzU8BnevLMGi99Yx2TNfuC8XFoLciydpuWAnyq99nXuaL
/viKRxwceDnCRhMDhJ1AsdeWph9hUDwQLPWvYEJCOwByKzgD0JD7v585OqTd
2b/McbZpK1ZObfbU1rm+mWapxG1Hw8A8LW1+DzF9xZAsnRZ7bdehw/x1dU62
gwZ/MOaqw7+ANNB3zA440t2pOpdXyLRtpseZh0P5DOOFT1qRKNTGRmzxFhw+
HGaPXp49Xq9jBCqSKMnI1CxcbjpH7/gJ5Vf8/tqdETZ2WWf0oD/w5L8xN+lG
AVhrNc/boWnmccsP8YIIrJNaJXBesANEXwsI5/Y9ZZ43JjCHLFcHihFtofU9
EisnCxfsT5w5YzZMf4julG9HqFqYpsTSCesYrhPXpln1oNu3Mu05YOjo4bAK
heGzE36CQmbiGA2CmhUqXVjtqjKLLP45eqxk3pxzO1wNzLASa5tiOXcy2cDB
1EHz8MpzKEDEUsYucp+9XJGqvTEYKtP3f/SL+gDHBA0agijo8wjAb31Pgge+
Th/6cyocLnYTFDjSHwBfw95zNnBmf4iPuYt2kRcAj91Wf4I7mBinv/BGZHXX
Cjhh+pLx3iiHHtM71jpJw9H/6JwvLDrWVEqmgQKl1A8qIB6dMMXmsUk4gzgo
m2c52hL1zlyysWxqMmnSJXWq1uEipEh6lnzdeS/VaarCDs8x0P2wdR39RkMX
K1jZuYAFrLEu3JY+QcXkFGadcCusRAQQruxut9VrNZnplDU+Hfsk8rdhLA4n
zoziPiimaQLSaTZ7bF18CCjaWe4i/htrJe56JQ3VF1aedMnfakTN1x8ZN2K2
aAkXjaSYExV1K1Z+NfueV5CgHCXLzMannXjGcNuwRcJ/ZzxvUzXygB1jddqi
T4lrY/6lH9tc5pINitHVeUuq3vq5fQbjHYgn65jPejf34uJKIIAnVlPFZ2yl
DgM5QZWqsuK+SNnLzTmu5EMC8vZnl+vAdlqkihT3hRDpam9dMx48npQqvgbd
5GXBe/e2S1WP0jDG8vmHyRG6ejt+rP3nc1LknodJkn8fZTmPzb8bVrnlIXOn
q/CPiS1wrZ8qTLPbZXNJOP6XJDfMdW2DTm6rF4tuWx25qNkPl+htHOdZNRD+
DhPMiA+dgzwzNn9ZRkZL3EvXFc5G9p0FJtlQrtcUZyYnXyOwmikUf27vsFq+
I9knwgUgU4jXjQ4/YbtIlNE96vJOt19KKWCSeoqfc2cqrqc2BW2JaW1ZVOY0
bqcifPbsQD7IiAmm8dvKDQ4SmlOunQ+NAqFUpgqzTOkY3nSRqurUUl/XBhkk
uvUUe99cNLWEcMRxi1oONSTI4pSUPoGvQlPtDYLaS6xAIYVjAtXk/82UOyk/
OiOy87GHPx22SScL4g4TkeDbvKRD+5RAdhIR6ZTEPenC0FNzOZO8G9SEBJnd
B9sWdNzf4WwT5BgfhOWN6TMQEpCl+CBb8PXU1oWE+31g0/TyTHCWTyej/Qam
C9T0Oh7FvKebjigq6+0MxL4QtghiVkePV9T1tabOJ0Pjw150EGx0RvNZSwfd
geG0EP5ZcIxcLdJR3cuO2OpHesX3aRv1vcYEDBdvWt6N4c5vk7MzPzmKSCVO
fhw11TaFr2bq3U7N7Bw5y5l2pSdHNV51e5/ntUc0VRdQPl2TXx5v/iDn/zhU
0qusW5z56pwS6q1xQ1QvFXMeeDZ4h0tbgEYq3CXUFHuRvTwwoWoqSWdy6Dsl
xRzIjKiA+O1uB1vRDO9IiINwsqAHtAAqw/YvKph7LpREI1EEmJqLurOrIYIn
W62HlF/n59JXF9r6gRydXJn0v8ZOfl4vIcUICkdSLSqefQtdskvQFbxdcIXR
0teZg6CMjTU35baNGf7ywLAEbaK3VoVGEL+wuPK0tL+Jjeg67gD5bxH+6yV9
ZgvWaVegU5MK/ReOiFh/l5rKPtfz/pQLCXy5p0zchpahGPbHCBK4vNH0gqqZ
V9EfkXEuvORPW9B8IGP59cVIXH8S00LK2Gjsc08YrK69VeDiD3NunWyyIPcq
7WQjXyZCZa9xk5XuqEvPhCpW796MTkHcTJdysDGzSxrATD11QkaY532gyzDn
+dmCIt2/ziY9O4K8WVja39yt2B28duZMWuZpxiGxCoDs8DwG0MQj4Vo5xYWD
y9GG31uM9pnSZM/iGfYKrsG0owXG5VO5ISwwVSeJYsya0R3aw1oUDJ6pcA5t
qQC1qn/LBF3aukfzdSF2dhwTUqTVp92hdhZV4v/Hnzb4qoY6lDzWapDNaUrC
TZ59A01mLjtAIO0QG/npyDQK7SZP4ZzYLQxVKYQAani/XtLo4wan2kO1Ugxt
adqnpwsYPwKWA+RSKwZwmeNigC6jYYtPIjlSYzgRKp0Apd3T8UUq/q/7qjD3
BV4R1EBf8xdPXxI2TE4MAX6kLxTAATTmxhBWAAXE7AI52az8KGeubaq/bKRi
K7LFP4YOqOk/gxLo+oSwfxqQz9yJdx+RxKEPXGtQRhsuOqP5Ic84wMfb7mMt
RH68NA4p+xuBvNIjjLl95LWv+CfIcrKS80xHx6pCWgke9VqwzzYF4ONdUSK9
oT5xZqU8cXmPQkLrEDvetV36m2tvwDxPQL/uZd85W+BnDwJdKQSgLdgzGaBC
C5ZFP0fy/xQn+8G1kCWIVjtOBZKEZ3KdmKzUdbHwh3q1EavQ4ka1M/OglPrg
xYp/gouf8PtDMrH1XsJ13NlIBn/xiMx4JnES/qI4tPYMS04OB3cLaTzhkwuc
VGL9qp0uvoSbd7wEvx9DAu/CVHift1kXSLnbLAcZuO97UwpyRc1nxspzIeTA
ltS7La3Hoqyn2jn2zVwKQb+NrZbtiG+KfPq+Mi1baZPvqiyKEPHR0m7vKhLj
O33+vuk+sXDaFWzeCyNeJKeeCFzqPFlqi4RDQOyMz9EJS6oaBKHVqMOZ/rZO
JI1PiUgmbOCkRWK+cL8PLGUySLOmy5eLNVu2Bw2OrI/0h5tv2LFTGjPxD6aw
G6ASjeR1PlLHaDA+iCPPI9MJs4izG3WhhgC/5iQc+UU3TT6YrI1WTFtNqc3i
oRvG377pxXHwsWTZVgqha9W7HGrPMbGIXEYyza+u02o3p/HW2o5QOJ9xx5YR
/pWgxUNBjc99bhmCNAF2U+2AScUTZ2d5qWF6egeEm4ioObiNbvMyBqFUIcwI
kqveh0LgMtiqpJLKNLR87CJhUGtL3sq+xETHPyKna0I8o2a0eB978gh2w+gp
iMQmzTeTHlCV8PEvpyH50DWoiR1GjTWGKsiiHo4y66JzeyASOx5TjZHjWTRl
8AridLWJxjFF02npkrapb6+9vlLzlrWXKaXjIsF2uS6cvGjiIky7jRquBAZL
CHPUfbrMJd0NYEQExVNTEviNBcVZoUCtPOeaL841x4OWw2/MFHpMoroCCTL7
C3jCN5aWFPrxwaR5wMYxmEQFCh6UL4k+9hhN6z3L55Stq6ikP0OimMGBrggh
HJJ+MpCiuWk405HyStdldbmgXXOkiX+APxKGBWlf//SqQd4NwbLcnfblWhaD
xBn7AKrAQYnPqfzTeDWk7ZaiLCZT+avjP4nz3YOJghXyLiYZreo/NgOyKw3w
Osuavcau0gIPtH9ldDpzt2kexTAjp+geuMHpxk3HE1Ijm1p2jnWqCtjBxg7k
A/MPZ02d5I7X0xCpzAdpB9mBkH/FRwKolAsbK0wegD31lEXogaiBBgHJRJR9
qLAIfdd6OCoIwS6Fi2ilJ7qSAYB/eYTGTRpZ+1CWAqjR5tZbgWTX3PL3q0wj
T4AfjLyDWdyrwSTtkwoFnm9ApSphWCUJ3y+TugvXcMHw/u9n/BNzqXMgKgfQ
mkwZYFBUiqfrhtktMI6MmlxWUPeHNuCkkIDStupYf9HhlXF7NVJvYBP9WnY5
ejdqdBTuOhTGsc19QTtNsWiqFoswY1iMfhaFGeq3Vjd71arcW3eSTl777XV8
jXvoqEPMZaIPInWQtKCGhO6JlL6/NBF6DGf9Jb4XMEUgIuo9QCN3GkOJlq0O
mzg0/k+oLltUxt42wRJRH3VUSsrDj5qNhRfUiTpie5UdbiJgIb3iFxH+y0Mw
bAm+yMpvy/R4xkJ/juSce6JE29TCTrN0jgUQvRD4GbgeKrMpS0o/9sBTjVzs
4La0FqRUN37D4hvRlBiMJpF4D9NSpP4ISVsuNT3acFpoz1NABb48sAwMWXbG
BeYCiGHlEih948JmsRITEZmTMv3pA4gpThhBIoj7DMkt5mBk3Cs28kim+m4W
2neTd3az33y2iWpjFferLxaT3Ng3iMiCj01PtvRm5bX3FwdLN7bfxW/gqoV3
LSJZ70pnuuFUqTRxgScKmOk6Nux2w8JIGHW3oJqYRQeJMmykp6HA/OUiM2eN
Y1dpwmnniGIDjBHhnRb10BZlVJx0N3ToJfAYVslnXiQnWFOG4vL943ZLAyFb
cWZDkeAdZR0Y9LdcNMXtlnB1qJ9Pe+LNe2xaJfnXbVHbx8i7+pNn2p+vPxBp
GkGQpEphBS+9BgHM0jG9I2RO0fZKU7UzAE6ZqHySRD1yMvdS7G+wuI17rn3B
kUH1gbWuqTisX0cpjHAhz6l+1FcX5fxl41zzcPUgbR3IFES887vCSks1TIII
YpizDaBmDDvm7Hi5XIUDzsejOkbSpID0x40c1ALRsDniMQKmQ4sR1YkzYPph
UOykiYgonwJJR7gZNXI4zQfhUODmnT+bxRcORxnYe/h+eAsTtyXQfmwK4Q/7
kSoNG4Nxh1WL3CNmmutVQPIMDNk0kj98ZnSJhm5UWkbmlEkNUlpuW+shVmMc
tZuOPbet3O8dEGz1laxpY+/JftTp47Ut5cMcYgQaoxy5xlm8dQyWxN6EVaOn
sLhjueaGWYkywg1iZ0T5uWfgE/XrAXh6NPbKGlNZSLElKqfIQ5NIbHOcy8QW
j/bboCANXiZy4BL0RzAlI3d1Zaypjrp6135BcBjNaJXiF8fVhffuqWnsByub
MAxh2zkLWoUnTtD8R2R+BLLyCNx47MyTdqXznR5tq8gIxOxalW+/UeWY5ox9
N1FgYc94W8zKqG7chfuPogR+q/abHOYxozWj+jIT49SMyYEniUVEVE7B1HsS
yWQy5NyQH/BeBmq+wUGKl4wsG41kxVmIquHbZpKGqG37TVqonyVPBWXfTG/7
WfUts4gWh3Q/ofTYWfYo5xJKL0QPyvrGoopE0e4XOZEQEGRP1+/fn739jm2+
aqajquAngTwYiqnffTQlIlFB7Sl/7wWqal+t2nr3WlWwUSjeUvuLEhhffGbx
9lwzAL+JXUElIXnCVY8mdpMzXWptN1MbrmYUwFEh5LB9IN51vA735hC/yzMf
fUiuEfhr1ueWJsM0vVF4A2z1uCX2OdWitsY2Iyp5K7CTexgTM5mWvpJm0rd9
2FPQLub12uZdVcUot5/HpghbRkbRocQ6+2Bmp0LazI8y76XqFRHNIumjXfZy
wt2n4btt/uUu4QXNwxZVr9Fcwee7Htf3km8nn+zNDeoBT0mFyD/rLAXmyfhg
Y94bvg6w9HM900t3ncylTMWTSZDev9h1BkE/04uT7eun80VL/LhNK1rjObGf
r3sy2gnec92gKgT2peXHafDEMN/Rf06G4ALZEq4pIVGVGbM4XKGBhPfhPNC8
q7sOSz/MSww6qFQzGcTEXfQLGJIr75/tn/+Q4c24SEpThnTlSiB9N3YyGbKa
mSKklNoFkg+P9OCFUkTsi3ikty6vYkborAf0cO9A4sHUxICzORHyDEsWFA1e
JdxC6RMPQwK/HXfhr4GtnQLtn5JzHhDtVG7wJoMXhUYQkIYgr3NW8dyI2KPS
lOzMKWjcIi+32hFo+qPGx3pZbAfy9SCmuuwTC33ZR7zOiyO1Eujv2FNrq+Jm
7SbW9MQAjBrsI0UcWhuPuzAXp6bozqtBPkmOUbQeWc4HrdoeuVxW+rVSpQz3
kbcWRHV/GQdMLqlwCm1ynq5amLQV9qhtm4lBeUszjsvt73PJuKEeQ9d2MN8O
1VargE6rHXDFN8vpW3bSnDKYIpb9kPAxTrOzDALH16JY4olS6rryF3V6FaGr
BSBOpMm4/xUtkc1N0ZkRY9dH5n2fTmGDd+PVwI7pxSFCYOFGYwEt0MaFMgiK
iwZJ/+HIZjoIZu2q4XZeNK3yWCBik4qXYkfEzx3yHYSefDL6gc3m0gwU8Bfe
Q+4Kwwb6sFesBmP8hLhrLmzSJYk3EPmFeknvLcju3zy4A6XWV8JQvXhmzf9i
bjVqmQmpb7fZg6NvQEslk7reJ73/zrj5edS8mATooXiTBmHYOf/xuePzUpzQ
lIbUAajai1rp2rxipwmYP5S4Srn79N5VmDGnSvJSg2CV99XTE9rLIE3N3LxQ
x0GWFodNuzk0bfvY8JyOa9ndd8ILktGt6CZbQ5H/gDi2ZB8dW/efOq+x6ITY
a0GvKI+qBpID9UMmfqoCMsBjtR8qeXuXG41xzyzYgImBeS4YbX/EL7KKiR8c
1NvW8oZLMLfWGXRgxwkYQE877kUpbacHEo4UG+ixonLJjUKIbeA/umRXzWfR
rbO7iugl/2ryR5clK+OCbsr7XGL/oIvEwUSGgPP7DQYYVAgqvb7iVKzWST8h
yfTPC6CgEUyEiJPLO6aY6wOW1NXFt7xte12OQx4lb+lE+py5YGmxG962ZUiW
vceF4vmxQmxDHbj5eOSdZrCtInGnvgNZ9OgSZheICOiTXttHNSnRGzFfLUvk
SAV3yJGcsjtk6jqjzraW4j5V37yI78iKcTEBxUQQ5Avyt2xn7JUaRxvs1RM0
ide5tMARasrZ+zQL7T1UJpQSPVhmoefuM3ktG1++P+wU+u6mOgeEz395qwp3
N8joQM7tFU9bJZmD/Hw3NSV5JVVV5TRm+YaAG2x4kch82EgkSdkP2WSgGGS6
s9Dr/hrmvD1jhcUGBUHCsDQIpZhD+xnJiLOKiRzYPhkNjoNdNpwvkysfar+3
bgy5SmZjUAVFvk1U/3N1YfbUohgxBSoaTYQF5tYe8y1fKGs+pLjjrydwgY77
L6Aue1VvCencmIEOa9IKR/Ocf8C+QCx8VyLgs7QBhHH41b1jfZrrlmEjILEf
QR8/jTaDavB9Q4KUxow/yB7MDpX/Uu7k5Nkb0dHNZ6is+t23QL/os1OxqYIt
NTwqyoY3qccWw6K5lkoHvalGopJiz8lcB3VIX9IE01feWsGmxxV8JH2jA7a3
IxiRCL12ry8exQHCUbLXhQFqNI6pheL1TS1/imEibEEbPW6/JHHPJnwskYpS
XnFVXXfPyUmJiC6pFEH551KP62z9AfXSaJTVPHaWYb8NBFJExHDIbD6PIrrl
flogfBZKsgJEk/sDDfYhpUcRSVVMr0jRoH60UiSvR04ykAavU5G5TZsUD2q4
z2FzMBJFQtXm+U23KQhM2n01Z1WE4gIkXJlyeoLr/jfG8c9jmxyWz7Dbo3ls
5EOoa3d8edk5FRSINfgVVVwP77j4I79JX53/yL9F7EVB0Q7fniVDjECzWh01
SuFteq77QXjVfUEsggKU8+wLYPrRDDgb5Ms/SJDRZkKNDh90jULrQ3hPXB4w
AlsblwC4S+NWUKMvGWqlhnmdFa+Cb7nQ0GaDhIjeqNlkmVRnZ51qb+oc4h9N
6IFfR9HZcTClC6rFy2HkSw7nqCJ7iZmFh+8srGWsIMDA5tmeKnz+tyYSLjQW
kmpyTHKQIkwbQKIUfnyozng1veyQszFBMm7GlfT8uEE36T3TheiJJmoTd6eP
nlaLQYfUJWtgdKGhVSvfn6Ii20gMK+76Nksi6Q2ZMjQCYn816qvrRZjeEeQL
26ZPcnprJFQaG2YXxWswEtRe7J8AMERuihuomwoGKMUnMpqd+STE9qzNvgxE
MARNHpWtmvCRmoqQpgG8lgfaTNaUjeLNITIDFe6bwziZWp8PQJlKIDRetkcp
HIur25wW2pYwbMYjdgS2yFAj/q8lLI2pA99HNugmA7XMMdbRrXynIMiltaSr
Pt9btnUGaohT/VwRrQfFH60FMu53z8nprm3OH+WII0flszLHZoY673A6BMdp
H07g3TThdyziPO7DDvtut3UmrQyzEDpcAMPO8KQG+xG9tr2lRZAFrDc/91KO
+OkfvdtBbEbsE9h+FBQFU0ESugMzft4GBPLhgQaFo4SSYDM1KAQKpY/IlWuj
/ozG4vqhe8lnv9MXjwfjQfq14M+/r0yKszMAzndJ4GuNjFPLKI55wDBzqWTx
TMDRLdGjAfuGUpe9IalazzKojJ2mSDK5KkzoayFhYBhCGeeE5FMR3PVhns5k
629HAILTBElXIaItXFA55oJwWmXdBrEpDprzld2Mf1OcMaA0U1aYRlUxZ1ZI
AyZlfzQRwmZ7XHJgcgt4nb/UezU1waOjRM5sniCGYQQ+r1ynRk9uzgEEVm5h
afCSD3yTnKiJVEsUpdS1qMMc08pApv+19/sbG4X8KWs2dKC0PrTCZTim+HL7
ekq9GnIyp/sAnq3QtEMTGYfQiyuU1tes7RpK4cXGbtSbX5H6W6IeF/X5xYPP
tw9ukfwQIfUlvZiT0HOvAbfOBPbFpvWYg6A10kajP/2bIzZcXuKc2rTDJx10
bTgrTgjD3svI3UURRZxkgMlgbo1UDoLyAHoycLYffRzSeITIJzJpg2MkSHly
pq9Dxorq1ux6NQzPUW2rYZwrfT0cH6Dj1VbaTYI43ofM2NIrrG+EwabLHF7z
KWTeDQhGM7FPEarWdnMa7A6o9LAylGBYTKwG4DJuezXSCHqGAnePkqsEP+Q0
TTqxwJRrn6gb3O7WzfwcHBgNpdWdSM5aGyavjWtiyr3h6/nH6TKLWk1SxJvw
275O2luv6IRfY9eojHx4ohWRIKKmvtcy4qjr80ZGDoolqdGf+gMdXJieN0CU
FHP/VhjMWgy0h07TAZPpS734kzuICo30pzmXOi0n/pQFLMprFKCT6vLDCN3o
BkbuNriSQtdpBbvUBLCUV1DnFjcYsJp9EmQAz4OLXbTn97FK6ZVJdEFkWrmH
oy7pAnE9+iH1hBzPSPfVEe572TGahCkV6QvJk8uE1tFOZ68+QJ96h177hw0z
zau6z8dEus3fozxcWbNYiGqaA6enEmw8wUhQ/1Z5puL08j60oRxpnRpOHc62
lmG+Sysko6j2e+dDMmDR4LDMcIQFqaxJsxRC8UY/Bv4xNpH4njfy/wS5DXeb
aQXrOokPz4+Yxcpn6tg6kf7TMAx6AMzxfUDEac/U9/jP3b1gNn/+ysr0aPDC
ce1vFy96Tr7oqlcuEYmeeBAITGQWQ+oAvTdDKy6YYgP8U7jSo02HVxIfwhoK
SW40gmh2lVe6R5PjN5GhM5COfPOhzU0vCMkOKfk+yk0cCU2FR+0JZuWOBiYz
K0q54tu7gZLkeNvBW5RpCt8WpqbeKTy1uEyFUQSmf6gLMklBmaRroyO8nYDK
uot00BWOj53z5eY4qRCcezElIn46gH7wQ9hkF7nAtmKJ+66RK6Ex43btRwMS
M9fbFe5i4zTUduh5k4lNuR8gO7mKG16ouagI6B84zkt/S/+IxAYyfbwAhjVl
P/8j9UaAlz4A2lh/GujQP1Rm0J4QKVV2xEFWgrGWQggzvDrLIMmBasONbTj+
L99RS+TVMbc3tTLdgz2QCcDuZ8NnVTTgSOLqhyaMg0RfphkiDhHRXxW+r0Hh
y3Npxdq72jH7k+x3DYsXhA58fkkk1wShb96riqCHBEEYPnxit+0bVemVdtc0
t4YQ74D6Vr/el1bxwMpQMgRTmWPnZfnttqYDJSHH1ElaupzIeMgPgsKqLThG
fHTqgAUjPtHNar6J6GgzQ16yavMyK3rlogz6jSO/RGPF+dJrCF5LOWYC/aj2
axTPJIbdHtJjjGSjZQ2baFIt9KTM/2ZapEbZqK/Daze2mTJzucBsyWLXmOlm
v9qIDDW7GF0sK39FJXfh4Q+EVzH9w3/HBAEAtoSfCsGnLMUJlsaMTHRdyr8/
mNpeA7yNGVAMGoVL9cT5q4NKOHsT5psBCYZNbm6vy+b/NKhgGKAilNna67ks
h21Ksdbz/GHYztvXeoRqT7nGyUN6la/8DkAmHgNWiZX9ysUaZnZ8RrZ/f4dK
Am9BTYQqaCNqMs3EVihGwe2zNub0YtB+QIcMHkyUWvu9Fk7g6toPNhvKzFRk
yHglvBhgyQgvN8hr3Eia8iL8KGO1Qrk8Ktm6xQEiYJNJ0KUFzL6V5PjBtO5+
EnOezZw0paGsl2/J9R9AO0tHu10QNc0nZoowbqPnG1GHrv0zke/6eQj3sRv3
Tzz8/Qu9dkWCxPQET6rw85mgUkFY+athYiw3U++kCam/IH/alcTbjDHbFwxJ
7xrA1QZl1lAahgaFrnlwkHSPe5Yyc0PH+xTnljoY29xG81uGFfjlrW4cIgRT
uuAnqOp2/oI0fCBr0e4RiYvba4jhVJrIdpLNF6Upgo4v3oM+0wd22EPZ5nae
XIIQdMmGSqOpybmnXeXPw1935PtZ/+Q1QX/KbZJTmtihGDcEGPaYn6NiPUQi
sJe8/dM1wKMzsaXdNByMJuw9jjBgSpikPxAJdTpolxOT3fbAIOwApBTC3/5Q
yte+ZBpKnCE/hu8OPkvFadbGD+BmdfbedBbkAn3eI7Ijcd4sTX7QFgWp9Mnl
rxhV1jhM1JnruJ5uh1Xc8hZ9+y+3XHFh0ajtyybJp0eOpGoNXBni+SbemVey
RYmb7Hxju07rxU1Ky82GAWCIhZ9s4FB9sURdpn4fuK741UjIE1Gw6HHiA+18
AGbT6N7m9li/Li4cu0WUXx06+oN0qhzmlAZ9onWmw505AdPGlRoN3X5um17Z
bku5NhP76CcIjmhquRy0wpP2q/hTFS0DBem0MkqoHiyMFuXLlcYsQUoUfsR3
msOIXhgwnGYSO7jKji3lFifSHeNxcsPAxSyKuaqU14Mr4inaGUtUQVka6vRJ
IRX1dXr1CZcz8/MioMfrOOBau7yE4tDaiq0ik/o384lmWIBkM91pAEnvC6EA
shenLWEVL5WMqddD7oF0b8ckKjreilon018WeQeYCQ8F/zhMs0NbPem8fHIf
tXWJGxzDA7DxvoRmBo8atzzhnM79UfQSHcucDZRlZfD5g92r6cUdhbRi4K9d
Yrg4JzEzTaQfKjpv2j8F5MPILQqVcvsAdtHzNrNUVE4wMCvSHzn+esfllYTR
do75TmllpwNMoaFG2vlm29FrUlNAeIODx1pDW+5UUHCQh3XGZ+n4ds5ELDwb
ohi4QRhgo/Kmk5oPjkVgYMb5/fMmOkAOubuHaCFsFyNQE9QoYzMTBYUnWXlT
Rn9R5v2zVG5RadeaeQ35mU3oxvG5imhwVrboEBB/ueVawbuTtcLdc6oNmMsz
2nOZs4e5UL/j+u8wqTT5zjpgzNV+aPqph+TDKSDrVHfGSROHvtec10sP+DsI
6NBnbV2iXmQNDYsSqjfb7lk0aW8X/PlEToirzben7TufCtk5DWdtWDhjnczP
D3R63WKMC5QcCgitvACSMmd+X83i2E6fCJFKz1pzfM+bgoTV8WaNCoOthA4U
2GVw7i7QjuVgmPJ9LoQbQtLE8ldurEKziRbKQ3isxkVv0wujtz9E/DOMgHT4
4ZrKPqJMJ8Z8HTfhdEGbvOVtpWmHdeG3fc/4ZVeiUjFjJFOiwWVh7yZoyI8x
0qRSOT7fnj8Zpme0FQ2DER4KHYy0CNPm/5h4zLrPVCaCwiIah32wnfrpvj9m
ceCObiZyrw5O3oyBQfUOnoKmbl0QzsVIWsLhG/gDZxJ3a+ijdwfQHoXwQ+aW
ijvPwKzMO9FqUlvqFEjAluvtawKbm6ncXFTmfsefkGVnoseBAQELGQTkh4so
B2TwIhfZyNSoYG35eOzhoUj2XYzCkW+hp5HHhxonpo127BKoa5C7mlbkmvz7
lhIGLjmfgDUIGh5AvrtbtuvBPr9Hm+Kix8SA7m0mL0dthRgSUtfjXr60uOcv
ZEX4LVh0zcfvAfjrymEEaNGD8W4XD1gOwXfwb8fXDZiFFXOORQ1DucEmVDW8
YpUABQcBsaHjJdmxmlcqQkzF4zWeFiDxxix2vrisCX3le0+Gu5S9ADL0vrIN
mYxICZBBwb6eVoJkfwF0oKufjOo2qjLG9Byd/uH7IHIVtFKqjnEDZxrfSkzX
3ob6FYEON6ZtucBbDuYItmG1Dl1huCU6xCCS9IRy7MeJwuSRvKl8CW1dEdh7
FrrSA1HPePxGo5zWc/cZhjRld4kvo4AKX/jmx3AwKJRbPeItS97jW8FASN2c
x6YS39gvD2vtAluX5qqKRXiQUHP1Z9s4G42OwCQKxl2JdQegQbgL3GIoPONM
Y+EaTuKt+Eh36B+Ov+d1op0uT6hlmwiEOwTuz8JYnUaG6XdXzz3S8EpZKuHY
iLn/z2XzFjgD1WmgYN7BYVP1EGXDA41ghyPNx/a+nzitFmwPpUKUY3KqspvD
0/unTMgl6sOhFGZmRvGNTku8OFlR7OZTiDS0mhIbuqJd3Kj+3RQmNWa26bSJ
8Rqlozu04rDwA8MwshckP858GG+zfz0GKPO/GOaMhVY8RVd2VIMJoIUO5hRb
o2DCOIf2IY1GLgEDThaZJDTppdeMmlsbtTxrJOvqlThv/iSOGfEVe6SXm31k
jzneJn33hxSDmd7xdwQcRLaJKqoNJG3BxmjDkt0k0WDLxY5kVJqOeelg/TWP
+oEZX+HOAYOnwUOcP0xWDNM/1HlrrIwM23jbc2SYeKvZsubXaDfteSrQtMNh
gAyweh8fMLIAUJACCKlYXPjYbJzpgvS4t6u+6fhnzmiJ9kWVZF43vNV5HfEW
19e1kgTLoDQEDyHy5idCvl74Qf5ZQ2BwmKHhqBWZ4hRDhNhY7G+hMoliEQv2
2WK0jQ+sO8YdMvAMEnVljQsTYKV5QavP5RzVoahVTw8hlGQu3Yq4u0iSTnDd
8TYTvYG8Ef/WZf0NlSLfFQzepv+QVqOp3/RAtKHEtifcJ3ontC+zL+VWRUMB
EVgki3xd+FFUh/gj7htA1zaxyc1S+O0Q69Zp0beIKb/m1Wot+FMxwn79RING
y8HFDDkCb0r6s3bQuFv2QBlJoXy/MrvgRYMWMgvNQznrZioYjXQQz8HbSclq
bukiDZC6J9S6B4g0pLwm3o8zKkRzVrY0wuFm/Do6oS8SW4nxbjL0laRltXXj
QRl/CjexSR9vReRQPOqh4fAp2JROwL1cpTUy0qTwKiww10hgGkgRY+6bgeau
IZpASbrIWc3vpVtInDMQA1Eu8XqIgdGIlU6k4cNrWwK1Kh4AlGgJ9tuHFDpa
F/puKaaXbE9qSGcvSBO+nNHwrsScWs74E2xJ51/uewX1Pv6HX809A6q14LUU
PxfEgZxutQ30qK8ldT1DWjzDKEtmZ87LdWnyKNeqAlC4kLFrc4v18kwsf5rZ
6ehzLtGE7KUlcQzkhZBgrNQD4gSDiHPAU9Xnxid7SBGbB14eAq47pnKSh0e0
Q+07TtmuB6FBqdoDr249B37BfCsQuAbYJkojE98Ofrbr6e0fXOfQsDhtXTWn
chLWis25n80ZqQhpRiXhMS81HfRrxGAd5lSaE3yLObq/7QyC0e9f2e3HuLke
IzQ+EjZ7AZ7GU6si5LpXlfXGF65dAfiUkOd3IwJAEn2SfePv4kTZIA10S1kJ
OFFjd3ohuxCcgaSxu7mID0ox1WRhZggSU60EafugLfPmlf0w8rGLVoZY/ex9
f+VIMIFmCIlQHufULqTnmtNyHLykzbOHHy6bzcOAXiDsIEu3Zpc1hyyqLj+L
48LbrJM+SDq7H9IkcYWSuPc/afAJCYw/3RaL66P/aj9U7vvGWOKw8ScfS5By
dzLi7AycIJq5geeVGQq0wAJXU75b6ZaQK73uzQ/IW6R07KiqcdYNZHbV72T/
ZX4C/Q/fejr5T7LnUQNQOCLiDFqiRhklebhyIJA90w7XIzckNXt1MPUETFFw
Wsc2JSdU2r/KWnrGUglUdxDnEvX0BxOUJgxfYleNfTpKzG2TLPIHlEIZmvEp
KIW4nQG4SWemcg1GLSweF/tmPVn7QZStXug6a2Aq8EXCwtE9JbRjMUd4App3
J2i1xfT7a7A6QRmINu+PLpYbexsDKYD4msBMsEvPzIZRYS+EpCmkKUvvZZ1u
jc7YsaPkP5M9JyEZXSkSUhgZUO7/Xay4LahRQ1v04d/g4g/hVzCWQ6jKXzcD
myGoGtLLGrax8G/9SCSfraUvzlYEZRuOGuTk5IlVturBdEN1mlooNLlr9cqO
NZ+n/8b6wiXrX/pnmpakjfaYWyuk1hZjfmlV5tk3M5s0j56aBKS1Ys4Co1qw
8BLRqMmIBVScdhkg8gwqfynIvcu2SreDHxpMg7fQoIiMZoSM76oGogb5mFnH
6C0uD5kyhuMKrjuhS2PrBJjIXuyMNCLJqALk6SxORl1Z7S7/LAFhwu1VMeUU
6fjJ/KgmSR6WSZsHCSe0RHnT8xExdAueQ9DEJohLB63rDcZvNlsbfjAwPGYr
mpXCo6IqIjz36ZC6LeflIFPx5osS4LIzX+4mZ7Peo2n/dmnq5wm3uiTMPfgB
cKGFFQy8khiDcu79sH+tTPzWYyXGi4CeQRsHL8gC9zvm1dleNWPGYNqVKUcr
sZeM12jbMC+7Hlvgwok5IW1TIY2FJBxVJEQVvqGRh3pU9RSnqBTGthBkzuWd
L4M9ytk0H0UvQypKYBcPc1Thgoo93nDR7k04QJqgd2rpuSvpYEAkIy9Q183l
sFOwrDl6yzxq7HFq0HCkldzUnG/xHHcuaWICSVFLgg8ipClvCJLTHaX/R3vp
5ukjYax5Uc7ejQuU4MCE0eQ9y/9VuywpSO+IqubY1UBHSBHqDIH3MGRSWA1W
PS5S18Mr1qJK7DZA/7WSGCtL3QAguDtcQoUhe22yheUMtLmGamuRvnGGbXJk
1S/LcLev1reuQRItSb1zMfNO89X/kPQ3ZOnEfQfte0Ni+8FVjdjnM5BWIkEP
d6vzETJFoWDEdP7q64LY8haGEfM/tl2hanT6hW/yZE7by/G3yDwAoLtjYd5k
eLLiAO2teF+oclCerooVLQar4cBdiPQvSuUj4egzRo259rGLkzuftvNwVdNX
2Adh2yh04PEvYEKUTCM1ej/2oMfQoWt9tvW2WyR5BjmelM85Bo13WhFG10IM
vb2IJ+2MuYXKLkDsME5go006a6fqxFq0JYAZKVPWYCbtBd3NiTAKBEjNHi50
KQ3/JcUVy8n82ihzu9cF4u+eqvgXX5COvvXcWXPWL/UUIh5nP+Z+ytMESgzM
8VnoPnAIzV0ZdNyN9KzSf/QEdvSht5nwAY2lYpiOlZ13gRiSTTDDIDEj4VC5
y+Sd8jp+SOa7vfpF3b+RFDXdj1P2jIgbhBbK4V9g8zsgWbbopxXZkFH2cddp
13kZxRYEpJgeQi6E4X5tr0ZANTSaefGMnlPPjOzR8edYxiJ7huZBWkZPuOdU
CMl7UB0AGPQ0QQIw+ofDfyon8tKK9lKUwIDB0S+/H6lgs9XAOWapLfVcyRip
Cqgr7sTF3qkW2s3rX5tAkHsVSiUdM7WhvYIkDdVuiLDGLc8+Bv/cfZHPjTGy
JuSOH1KW7lCRpipYxwciJXWR51IExULwsx9qa7eSCCiQdiiG7ugg2wsJIV8X
e9+PQnh2lCXNmkD9VOwJioILb5mdRz0blaR91yolbx4FtCaOtRwlqOkHt8ix
DrEEZaYA74laS76VVY3GVoxIZPCZD5NXNaUvSy8TfaGy5pBJKsozIIphLor+
ncOxs573Wl6Js1CKtvyJjPPdvDJfdHcqu6W79dUnvp9fJwN4PxrXySTJS90N
Xpv6ywww4eHxZaAQFqUNscGILahyUgte7gNm9nbs9WDClWQKMfbh/qqjxoQN
/PoO0QgDELs314+Svtv7YA2sM4TNfQsJQQORUaKfP6zzAaA7WJZd77O3OBPZ
xEzS280GO05kr9GGosVbmbR67qOM/CPmBvwmWSax32gP7VwzdDmIau1inBvK
hWWmOgk9c7z+uZ4B4Rf5lEQ4s42ufVRb9aFvgivTrqgruPmxx45VNRHYSHxs
3CnmGaDcnEoR6tQgNc2XEVicbTPPi9rpedBY+jEKyWm9b0PIvFhmKdCkztFV
Q4dez3kpfYyGRI/B7y/aBg4uVuxbvXHhJmBpMD+ax6s26MDfWCsXOc5kKFOq
BBTOGSUypjRmC8y7IjkZ9X0gS1I41RbCXf+jJxkRTikA83cvjZW9D2eN1/mV
YsaIZ25JNSmwB57mIuidY54o/F+Dc3KShJoNPBkbPwjKFrlnNpVSqYcBaArp
hz6btOIuzg0ytdoBziSrJk4rP72PJVuEt4kiVT70smCl9HRiASnr9Vr2DGPV
qRcRGO5kCnk0j+61Y7vkOISvF8qAIokkrbgMcdD6//ZNA5LaxpvZcrY4BVLg
BTb8MkxbZbQityHeXlDcG5dgZtoTtyEno9q0NofUiUa6BtmaEdrZox3b3ALv
Lm8+PjROD7plrRmKRkkvYQNNvgID6PMTi2HFjweFhezFIP58cb3WA3qezw8g
96UOatmOP1QE9YB2rb4UCf8FLkYSOg1FhofzHe2Z/iFxlhi7oX+UeXrxZfUe
nbG15Y871ABBWpa4RDgD2mMp2H45DIDLteh2vgzrW0UParM/sEMaZf+bOO6S
qzVdz8VhAsi69xlpB8o99PDU972MwLWeXmxmDogXk4jtWZ0roQYasgVX1vxk
6L2m3MSEF+/IKACDaNKcX2M3Q9cEs96mkXjLHHPaByZjC2mZww1BlRq574HG
vGiG2noKN0nNQGl/5e3Y6qpOdblpZ3+3gm3LSPhqcLT4rDdlgg5XbmjlzDCP
mPJrL218saaa+d9qR4c14W4m/Ku0zpWxAQDRK6NgYZtwK11oL3WYOV95Kykz
uuVNOjrVSD2osZ1O3Sw9sPXzzjvZjexrpVJnc0eUlO8geWtVBKUpr93BRLi0
mfgjngVOIQTbI5a94tbuc7YhCRov1SeV4bOxMPbiCCrVZcARVtlgPxHY133A
QdujJ6TTDQgb7HVAbDR1nZGB0BxRjkRLdamvDIn7KTfT9n6sFSSrkoi188BG
8vJXqwb1udjCfbA775ACxJY2QFgZfv+VwrbsxC+iyGLHcNwinKs2iCSWntJK
42JvUsemjemW/8mjjcWQKkrrW2kMBvD2XM7Gul7gWaM9GpGbgjw6J9+sALRL
MX1AeycACS2Qvrgua6GZYPhCqLmy7qjEt2kTfJP2vKGy6dEa7409MxGaLN1N
YOIn+xUZsrveukfsG1Uti4u1msy0JMpNPbAqF5b6DRabyCVx6Wjtqaw3STEk
WmSdFpkGOk59azjtoRkpw/10nfRU7xEQF7CYfPGpc2Y9myoZweKOJmF33ggN
p9q6r37uJ5wicI79YKBwcm76ye1FPZ6F9hrDFLJjO/QPaHQ+Lvdk8K0rBktS
c8RSwYArIVb5sek37hqBXmxnb60Nf7hITP+X93S0Mp8aXtK+ktSC51oxGNtm
ShplZ/FMbSWx9yxnbbhaTMXwAi5WoiQtvOIY5Yayvz8H6poWn3RVItP1lnAs
kHhxo2ZyfqwJpJfQBZWME7bgVswBU0fJqUmBJcEeCijr6cHj3DZjwTinSEJv
brGIRUX89yifoaHY1VkRf3jxL4mwIfkrJquQiytBsttn75VsAh2VCxkGasn8
maZt5lWuZvZ2vqJJh/M1dXz57DJrzhawV7zliJ3emhdisPY4VcQ4Y4tXoywE
NP871b+1m8Z3EIQy3LXpT/X7f447Q2C7uxbVOxq2K3QtXUi3MmXiN7vYZGGj
tbhBtaFYiBFELGLr3Uff8avBUy+pjKsjOONOoxz9HSck7WAL+f+x4Hyb79TG
XJsq6nLw1dG/s8vTD9b/hZ+gAYkLvgl8mrUmb1h8XwV9wNCH0R0WmsJIbPxC
eO2mnSd2U9GhOXItby1z2BXZnv+K3xAMyMe1C3Ev27okIdCFBMOT3e2BPwxu
WhlhMpE+EDlyynRMdV0FibGB8PyrHMG7x4SnAKyLvrLNYnto3c8W4Igegx7p
DOUngZz14zrDVEGb4d4RyB8CHjomd9VGOLoC5hS5PY7E7pyNfldBLEmw73S1
Ouf6dRgMB86m4i9ZULAj0d4XDjXD/JAORIp7xUpyXow52sUbKQtBKybQVFzO
TH1E6lQGJKBsbzC5eSlhxbeZmRF5dzHVyL2/rGiQJawpEei/VkDaoIgUWKq7
PFWJGhjLQgpYMyna2LDAldSGEYhUrP6IjGp7k7Yn7aAznwy8nP+TxNzNqgbf
o1gpz5DrbAzsd+ld6y0RLbwk44zmo9Qlk9RRn+L8KdqlvW8zI/9AV379PQbp
nnNQ8zZ+9WNOM0ulyCOdTpD11ZzmWJXjDn4CWrSkzcnDuN1TaE3N6HE7E4X7
yN07LgX83h9DdFiOYah7RzfhSyZ855GuO2+BMIMR2G7yGErjmGZMgo/7g2Jw
pKzKOiViCBWFGTjGo1uQ31lOMotHY13DVJFYfsnQrxbbQmgoLpT7RTG7E1J6
ghbPFn9QWA9jAcNDikMYrjn9nGC7ipXSnZSlaP9B10bEufnUw3/Gw8zI61M6
TLAf6QjppM3itFHMGtRNRvxI5xwen4WbEUVfQVE0rK7MpnUczVuwUwLK6HEh
SK7PPw39oQNfhF6atLqkq86a746/ZZDAPSt1ZHoOqE0bvalVhFBTUCbPmx2c
WYL8HilGuj2SB4AGpULdHxjSVEvanyIOmBYFjIERbq3OeKc2ZXcQCqICdl2W
1JFZSBmxa81zcWugol/AacP5aFKhgt6EOgUhkzrCJJKhy+Gouy2NRmGbW2fI
qM2706e/vE9zr2KVK+ZsE8AzTL2dMiul6sNrL3MbttkVhXPcJXXE++zVSoYU
FscMyeCUYcnr6blxpBBWLpXYjo5xjskgIPN7mZkVtuC6x4SLx2lcw+7m6XIQ
sV7+8Boljz6cTr3D00b3Qg9FuS3CV6koPV5e9BYr+B0uomcvu7y1E3bgsvSE
65vkOXMNgb+EyfrVTvTQfKAqGSX8cohgfkQfl8QO+deQ6xL8RuRrVBZhKtjY
FTMP7ZT8M/MneC8ZoWmkh08w33ZDC6H/nXTBjv8fQy4ZXEZ1e/T+dMXfHdSk
aCd82o/upbedu3Z/pGtqca5HT+nFe6cLEXWizndQcLGEbzBjS11EGnjnNyY2
Ke8i0NV3fFRPetlmo4kgutPM7JTP4eFq64qRbirUwFGngpZpEaDrQJvwwe0U
aHTevC0nHOu5S14mw+ocLV/WpSFPWV+6OAOxXhx9r31Y981yKA/nhbrV7vht
tmK1ESyNS4ZOqeQ4DO2IfOvhH3+mkfQneu06pfWAZRQc1cs2ECPsfr/EL9Be
NIaW/b8NJh3r+PBLn4t2EYuLt1Tr7XMsFfO1nSJKsF8YCZoC+bgKy7R/eQeF
pRjojiqvVpk9eN+2EOgB/1tGnp5WmCiu+wJeD5IKdO8+g8lH1pmTf8Qiq+Ao
qXM/PDGbjEJ+j187K0Zbcsq75Nvo8wmxer1iVNmuIiq3osFUSoxFf7T6x89I
sWvQDIzBMausCQLAFk8GRua/w0T3qUyvSKGwUShfan+apHkJv9VFz7QVzljF
Fe4h1Y3X23cHkIWRb4g5sFjELc5AYsJvUcGIiDL1ZtNiyQUPQqz30HmNIdpX
w2V2AAg8PgDN114Zc+aNu6KzIQjPoLs8X9bB3jnFl/oHaW75z/Wsxvll1F3+
0ttYugJyri0BFhzsDlWfUiiu8g03/TsmV/daDwj+J123sl4hkIrppLIlmWUg
xaosuDZJS+aBHqMlqHJ9dRKQdzwGyQ/Pl4bm6a21n6bA6JfyIJd9jJ6yb8bj
sCQ1h9/VV0i8/8tv49VZDrP291UHwrN6ZJndKVNwRC+QKZtMGnCAaHbUPoiT
20v+sIa+8DKtNk7xIIlBSLQj/PZZOpBx5smPrq1ehI0mYC2iuSpiUhmcTld3
N8/5dULk+V9A/WT0SyMw7dkNsMT6rMgr3yrgeko7lgiJU2DiPQS0qQl0yrrZ
n0zO0nYD0SLfZLV+iMThoWzecCakB02gnu/pf0ILN4jmXvSO66sxU9Tvgeae
T9/ZCjYw7m97XlSHYyHLLCA8QTqGMzYz8yMW0o5Ezx+tWH9yc38xbyZ8WNUO
DhiQL5MsFV0TdtGc7zVcQOphmHKU05Aty4AdHvxjks0GhXFKCNEvuGBojQQH
8zReEJ6A8ihSUANHDTh3sPCOYUDsEJYmCeMbAk3kdVpGpo8NRx9Kr/PM2/IK
rOmxWHB31eVEmFDgF/srCpcQSCf2sBgBaXaWYZCxizDW0Xjli32lu9mTWHOE
JIWQ/b0TETvH1q6MFRwwL+jDzptjAOX0nY59Ukebd/S18gOX2TLzxtMiMuoz
6Cyh5hGqZfwdO2Y05Bf3LDdR7HU4aHWJgoGp7qbRc6SFij2tvR+20JPBOHm+
Oemax4OyIAzUOnTmB/PRSdzwdVlL0Qg0P8R1KQOF4RFOY4t98HK70oQ4vAmq
VYRpxwSu7PAUW3obpbmiWdwCotAqrApaqTbg53oAWoBIPMZh84DFR8E2+bui
bCNp+8FwdNJ98iIBujTglyg0jaXuwmE1qTKY0SoVaO+X5Ims216/pR6TdaYG
duBasev8eYiDkdYjk4D/9ewN/Xl71LZXr3QFel5pOanmLeJwReaJo5i0SXq/
g/t+4B7eObduSkQoGek3uH+didk2DmP8I9JZ0JMD7NTocMLeZ4P+NgjC/dI/
/tZtIRFEhEbmKpPPb/RKQPrdVKq0waiJrteb+WdsHriElhKl9PrAMH2nNK2J
V1roRmd5rYwUBtPklljVNp5QbvqFoi4Gy1zf4iYl0D3jcdXKxebCMrJVfxp/
8RxOUM72FrA9IW1SbcHmwRy0qkfAuElB1lO1PGu0oXhQwHon+38fN8tz8R6y
QTRgqSGLXl++qlRAmuls3WkFERu3ynTj/M9ad2CNA/AjHmTinjXLS3NRejKB
KLHoPwm9kzIXHTTTdZ+RXvQIprFU6cmP25MRpa8VW+Sw0nWj4LHfzH2+3+eP
RIFgRRBwzpsijO+QCs62s8GjCuDVc965C0PzEkdublHSVUDG0GBCZD18uawP
LUMNjDRmvMC8ux0kLkYBGoxVuerXilkCLDhXgPImvgMVVWKPf0v5SlJWVvPF
iIAxO60JbWa23N3W1rr+oyArctRAj/bFXxJGEFYqto4FxJr6wTyFGu4MG/RO
APLILlS1olFZwOsiVIK/tJN8mKSOyJt//uAl6I2Am5UlX1WDygAloipc90Yi
1THBmXZ6paLY/lAavVaTRyZ6ieMo5C01eSY+hyZENyV9IFHZe7q9ot3YDKAF
cbPwXr8/QwkCzy1JAVmnPfGSLOgdyzQhQG1XgK/QywFOdfhH8PYN+h8F+vIW
tRVgGmJlKvKX2wltTkskDq4nJr5e+LLbFUq//2Ncl6Fej8TxApG02hLL0U/A
4e07K5MuzyADVqpmBI6aZbrHo7fTpCieoj1LvS+I3+qlpfajCmiEHOQLB7iY
/eNqqux33+JtKow924WfbHg8tGsImTwl/dc3Rktg0dCuLoVxcRRs8OUtwv0A
BpVUN3ULN2ZpOovlPzguEbkANfgNin7SrUWm3f2BzuKirPHIl+XNkDedGaFn
R6OsxQDKu1S0ik/vHe5t+8yzY4yv6QFQnSgsbVBEvDC1EMmKxBr6C/QWA0ZY
q2nFrPu2IXLFWfs1PKqopH3nTyhEmHt70BihOas8ONQEaHUX39FXzxc77DiR
RtUU3AVX+8BNSkQlRDN4ksAbW43IWuV8fRjcFfT2kxfYIrJb4DDNHYEVVbnj
atzku37EJKeFZHNwWpyjr5yyGh8CSi9GUI/Dr3LKmZLPfg5Nu+BsmSYokTWQ
Gm1z4evqOIRdW1PqNpfI8blvxjGs+i8mEORPDc8PMicTJfL++/itP74EzNVE
wvGnkpgkZje/4fouzbp2poaMyGMv6JisCtjSvKKuKHlQ/qjZGY328Llqdy44
GA5gPYtTWR1EYvUq64D3eNJrQCcbCDEf8eaMIsJmjBWYBqE32TWly+woQ4HY
6yZzt5bR0Jv4PaY5rLfBa6qUgBFlhJfEVFzv6VfWlzdVUqjiWHhdNyEbjnW5
UjHAviOeJPIjv0Z+VRMnjVjE7G3HfdjeQr33Mom6tcgdHFi/bXspbvhzN/5y
gIMfcDBRbfuw59vNJFEkVCFdG5cj/xfDkAYm7IyNeVVfzds7+5x/X56vuRRF
hBrQvLH1m/nuBDYn06SpBJqI8aPeVbOzzbPuh9aw+CQ5NA9vStj5GLsO9bYH
di5fvGUvfUY4VTbiSWVX0Us0a50R/0JZ9auD0J9lWXoYwNtXV3xGbRXvyVq4
UPK+Exj2txBmV9VCn90C9Ok4HPnQrLnS0RoDkflBdGOlPjhYzh3aL4peuhES
MXWwMIEXolrUfQaGkufwCmQ4iv7RJ1ewlCK0bbkuKmBzPW5LFvaf9NqKOZ5g
q5FSW2XEfmrGzqgqFAlUBTMw2g/XwX7r80C4qUYmTIGJnKHxYdlpd//WoEWg
7j3OBmUM89JbnKvvnTLjy5EWkY2y4WNLjwbXWt8gOtLPmpCCc6+4aFo112ib
Dyt24vCtSuQ4I7mQYkGSknyTD3jxwqEwohH+3AXqN16CxZCvTWfS5H0SEtmC
0QROr1+h0inJTmfGSfgKWQfLOKAn9rJ4x9fETGRI18/ksHbDy4LArYD6HXUx
0jYt06dOSa7+3aej38vZRLmYmZnabPpPfKrMoiISUUDrcEboXHia5aK0qDVz
yhx6lE3luX8/agu7x6KG+YktwofkfT5LMPqZmg/vDFENU3LWYchQyeyGK6Kp
4zNFO0vY6WTX3kh3ElrJywDse8MVbocoLFLevOMT49QY08fX3Zp65GAeBVeS
nxRlWYvWPZk05IrTGNi7oogPBJfT0JVcQZPl7nkKiRfcOnHi4wVvjI7Wkwcp
ydZduhWaGwFgvADxLkJu3PFisd6RPwm6deYko4T0E3MwFBrwkTPTYLN/Zkmq
HIrPXoZPYPllclWvm2RYnIKriuV7S3oPxL9vvF7aI0y1hjFn46EOIcHd+Vmu
V+N1DfRBh4pLIDKiidDaEBtJ2TxMlfxN8803+8AOMP5YyE3Cho6eC1OPZtkw
qL3NgbSJobgwsOKX83O98jmIyIC2iFvV7WZtX5Q8OJpXQxRQSerS59VzIJ/n
O6caUNQ6E7czQ6p2Z9G6pINBVRgGoKHNfoR5uxcVlvQlIwen25S8+jrK88XB
BxbISRgmp8OsisO7dgwzv+KICebvMIY21lxepVy1aIq53HYkYnCd5/AsTugs
Bb9Dp6HGkdsnZUsmpAI+Xyz2xm485xt+ywTqNdl9zc1q3oWmandDQyXKh7St
BZohifwzfMzpncpC2/SXur1SyAOzepwDP6kVkqdimTDjmWLhCW+4bx+2b6Xo
Zj4Uo/PwLn8aSZ6aYXOgnvkJrYmZ3yJCHVqSgAm1/544626Bd3LF1t/FjTJu
iUd8E+F6Cn4tPtmIKvdEwrsUSx3kocjdiRZuOfiCrbBHpxt1WmkYsbVpwT/B
orm6SdQXR7hmDSg1+95Q83POgmmpbT5Koz6A1mkfV8WPpueW0vCy5AeZn8ZD
R4N4eIpJPh8rb5LXqYelZzzG9G2Yvx1ZAzUrLqJYZgtfd3B+oYHAE6NGTnAy
m3TvyOM0XZAB0yzpkGiY5Hk0A+PKWApZcaISUR3RY2LIX5ZYMVrIfWMw6q5X
51I2/SDT6TQANw0h/iUwxov3+M007Nk1xsy+OA8yhjNUK4wSMgmj3tqERXYk
XqXfHLw9wgInqNPiUGars/gGigWjiju1BR5jeDi+RRdNC2zubwY3KXIuET9G
DGx/tCJIu4kFMtN4OPqMxPoqCn3GlU1+LGEiE4u+CpN0+vYLAQyqA9ID3C9r
jtc1AsfBCwqugoKZ3SHSZfN4RKQOIMgf0nDm5VKFoBeNq9fmYJK6Qsqgl8Fd
qQH0HEJ06FSh6PMBmm70KIVln+IPF1RcZtpP2a6amdJsX2QtXsNZtyn2TDZY
nUUtrgRFghq3/geHUFxBaPwiauraGIGV+t8lwws9YFM+hq5Lq48iPbfVk9Sl
7zgLOWZSnPeKaZ7Rm9PXtiK2WLuqEeWlgOFwdPo2JK66OxPwHJwUg/5kXQBi
fUdTyp1YrKnzSGo3528U93AfGgbBsZ7jbPKi/afgdLVarfnWD/vvaQxnS1OT
gIpnt6uD42SxFcI9o08bfjrX7/KYP9JcyoA9meBvh5ReTl722aDtsAffcRzT
xpclKCX0+5LgGtYB6Oc3nVV+lU7dVEzipo73j+o5O4o/WTA+rdpoZWliiLXG
J07f0fEVTDWiVT6AEseeSqfonUWFwiyFxNcDhvn4I0bg+/FZ4rwTxqJabhqX
vCvlID73dPmBIr41kKmShtAlxhco5miZLx7Nh34XoTUKqpX83wlvdwVyPzJv
AEHm10ERmDSP06PQik+IORT4l1LaUW6/hVej5wj1lhYXHFjh9bCiLeiPb9cW
97MXe/tpnnh01NWlvvVM2K/obeh4IF7v2QqIvjgQJ16bD/rLhYlsbQmn3nST
bfF/MT3EXeYkexjOx/e582uIMoHPY23fBqNI2UTsOywG1H78WluVkM0FTiGA
vTbHPckNYgkY6EKLgZqNo6eDWfJ3tKVEUdNC7IJfRXU1z0h8ZKZIfVsgNEJY
0Pfcq+Cy3dgAQSu2NgDZNDqU9MM3k4erhbA9JCw1OtWmYlLh4TQJOrzGeGZ/
LPEYyrHRbUnVxSymqL7HdSjwGDDQlHLpc9Wslz+KP3xiLYWPzzxncPJ3jMxm
vjcKyyLeKxFKJoYVfHPMgYeiYzqdh6ljRIp87FmFqiFNkv7LpCc2GWNJmT/b
SSEENQYEJ8BYMuGfmb+YelzdAz00eWXsN6Yp+eGlssVl6GmUvMzBg5RLNJaY
5gVaHsl8HyQE2KA2Q2SPJIZ29jtnuwUJNx5g2M5baTtcPm0qCVsceo+DlKOb
rE4H9zB8mMqd4SVOTKHfdArIENxvt5e7SaMq7qkV5Lu02AnE1kqvGblT3UR9
LV6CRZJ8XYDO39OoPZNESVeQRpjRZms/KDbVil/wbgCmRIkEnqME0XXE50L/
oWJBPF/k/CIf+p2PVfSNM2jdl46NiQZ2qBftT57Ba3HABtBliUtYGTf74d9d
e1Sj1yrgKQ2HUPMIscn2ZgDec9ekMt+kcOOV1sxM7n7wgtJ1lXP7jImdqWuj
UU6VfG60CFxosuCWRHqtQyfwRdkjqOGNpQjCo6EMSmj4v1UD7LKudGLR8pti
eXYZaliPjqC0PyimuE2HQ+2LA1Wm1AiMISyvZkkyH7bzZp5QClMCbi8c4Q0h
udc/EgGCyyCu/HUqqTnM38jqwGx/nce0VhNyopdCHAZjArQ/mxiovwVJyRzf
5k7arS281pL9R5DU9n+15knEI6IxDgxrpW0kizSBWcwaivQ9fyDZ+NBqX4VR
6G7reFCOid6p1cAFuyHG5ciJVjHMSHu0LzaR8YIm80S7U1i7oTdTQ0R70lKY
fvIowAn5x3MvRNNJmCpEOZm7V85WfZ0ek3v7rujBiZw6IJP2nCfsx/phMka2
a7/FrS5Ug8jNIuBAQJJKiHXNMA8X0poj3nsdhcRKQN3HY9aWpmpMGbEnpBYH
r8d9gJck0XyES78dbGMWN0ETZgQt0/Rcj7GUrfQbQ7rd3eh4k8q69XjcnNNL
gsRhS/AOoqE+xDhOUMMmMR6uzBC/DTW/JNnVgI0f6TgDAOUxaocjpQvAM2/f
y7EbcchaVKSPc88BJbntvBTj0yHBLK2+PKCRbC4C9dPT4CmeaEEu65bdQyXV
sgHLt7O/QsbWuL6op2beWr12snauYpmrOmy0MrYHXu1Sgdj/bzSj1OLxCuZT
Z3Vl4rCppWCdHL4EtBMOYTkDJBfH1Ai1bFRiWmGMvOjaUHMD1V5+SivY2Wyu
6AeHas1+1D3IijzQn02zDkz2aE1VF1jOGfx3SX4Ct8jWygh1Mq7fAz/xJLe1
+bRlb1NvK7MlKZr36KISmwzr3HNmG9gTtvN+sHlpBGaiLNd60epkgS7uXO4/
NwDWwlpyZQwEDQQd/sH0or3qfq73NZYpokLZtDwTHw0ACQjTQafoq42wy1M7
JMquSBBzTg9kNjd1dAL7O0sxnRjtGLZK13kOtu9azSHGTT0BFryJql9wY0oV
4HeJyh27MgKAcDsWXwGFyYtmBpJ6GaPdYGiFPbclkRgfnZbjDNpUy3HYA/Ns
++95lX02wPj4iYcWt5K0SCmjkRJ7x+yBby/DIW64OPsAvTcV019457+b+PlF
7ZQhERc/79BXr92L3GvXF3GqxwDGdSZFGUO1vQEvLrP3VpVGVLqnxcOX65Cf
7L7/hdWMSB38J93Pr3yofwcsM4YxmCDpfX0QP13OjwRyLL93fgAmZYLQBDTD
a/fxzas94PHGvHMqrP6/KnFc4rbK9e0d/nDvcyOD5dEPUeZmv0vJehtv2QM+
q9/WlSi5SVgfcnu+UFdpyrFOOXt58/j5iI6hFYwJmfNV9/QQpuizsfUgoj1H
OhY1ADAKyJAtuBGGGt/0C5wzBjorDWnDBsQBal+4IW2uqHS4QOYLEdUxXPWk
YBoxCefJkK4kWV97HJZIY03sFbPsHqi9jNU3jR1PE8vtTaMgj56IpNUQ0ya/
GCJDJ918rB1/Tp/GssDDUd3KuEP+FBT3mAIgMLQ1RnFAtNEouyDqyELO0mHx
3vkBOlqMcSc0flnM4A8ummrft/7tpROUa9+1d9rjmq1Kb2NOX2emvjcy3fZJ
TsfPa/YPgieygVt8IJLUMuMafxvUdFA1VJx1eZIBcoblY0KUgfsttrz4bUpZ
EUyzzBQMw8O1P1g7jb23Z5R5d8NXclOC2OQlPAmN+FId5QB09/amxYz3tVsY
3nOilWMccXQLKtj+uvxHbgXlVOyy4kHO4Aq2Lcx8yD4KVBvHV3rP6J3o7dj4
JpOBqwpXMl0jkSaeq8sPMzq1Q3zV7+j49nRKFs+PYW54jkdzh+Gx+mLVcmvr
oPrjj6fbhdZ/Rj2Ued4hxE+cu+TX1R+OHqW0TtlDBEdEbQI1IyBYXj0w6rcO
1u4V5zM7/ERhEfe2NQhP6vzmfQmTPOCHsQo1J1ERTK6jii/kd39/QqdwFM5p
5RLUnUkH0T4zpTdkMm0HyX8F2gHZD9ImxmpKCGp1wDrN8FAfVWl/QxOZw9LK
9p7bzrP/yZuDDkVBUAQJRRGBQmRNi4EK7OOtbaFAR/Y8/v+OZka/8K2LOd3j
AWD37J2kvmWCE6D6Fsw6iv93ilu7MIPdhQrsImuQtzaAupAEKDrnkBzBN2uh
42AaPoU+bI0oklrOxJQiX4w0DHKP5s7C4a6uQAgHux4mpALBiwS4MCtURg08
72tDyB0SeDJCPSXpfVrSSy9RfKRvSBotbZUMG60vRmE3r+6hF8iPJCA3mIUx
lGvirvQ+jCFq+fLQ+rHWLOGq4LGYTywu4pJE2XEt98mrGIN6vT1Ra7eMtuiL
lvJcVBKkiYbgj8LWjs8BzC1T58HS7XWfct4TTyhoqkgEtqlq2Krd4Eooe7I7
f/9IlpfagjdyJ6NImRPqNqQNfpZqT7Nlmy8w7suIj6bt2IwE45fMK/51+fNz
I68YgXaMtb6EptAaSYJo7Z5tFV1SVpLtd2MRqsYjKrDjUuysqVftNhIMFxpN
vKOXM6GAWK4EMSoZTpKD+MUV21BXlgbbse8UVKOSEUvAECS86L+3q8/qgxmI
Sjo/ROI17D+DcM9YuYcj1iWlHiWN+wUvcIBDE6CdZeCjSgBgxZELfL6xV29U
1e9/6Vjl9X1VkAd5ppZ8zOupfmS8lHriyf/ACZFJcuS9uqCJtVYLmuifsScJ
D+vvak8KrZ5QbW7evw9Tn3eG6YOJDNeqzgaFi7iCPkN3KDvsoPKt4qaYz9lo
T8d3AYh9MSJbeZGD5pQUtG8MJPwZFWrpi+MWd9v0VoZ7IjVTkYdudUnI2Vlr
ZYr42F3wWz0y1cONnGib6PjhCLpHvGHd0urm3NESj6mr+NOxyU8eiHvyFfpY
RHUNF46n+NAS/AG37WX/NDZ5nSEk0xYlQN8JgFqkCS0IOmfYeWU0Kg5umu1r
SGK4iIsuuNbFUvyEukqnQncTv3vpO1qLxvlFm/Y3jRAcwvTEyv2cei8HVZbZ
qCmIwuEh+mOLVp0JCmbBqcxvQFiiuxtCjvPZKOh8NmLRmrO7NST+7i4Q3c/U
z551RDTj9f92fKe6ZZyUFlnlR3qO7Cnk8SWIdyvK16tzKt0J/xw9IlzXAJ70
l9bZZv+rJWxQB0eOAJgkZRlCRlcoj8IoL1TTMliTe91c4BbXisXb3dWm9d0/
WAbzIRvCnhH+wOmBAtDisSAFCSmqYTrbQXuK8MVa/3OZFHobKMEGOvDBvgZW
uNr9YYjvFS5NuEiMZFmY40tSJlpKGiQ6z8SFAVH4n8zNE1zlhY9l2MPrf/I9
t5apYv3UNON9JKFrLS0+q9r8YNf+EawwwE1D0/8veJYtHurHqZrL3SFqtA9y
ztEcf/e3vcRaFlZbNmD2QutOqgAN7kE3fC2cypuInPDMdugZcVR99ufHMI4x
xNDo1bm51UFpbK2yPsvAcyAbl1cRh52JpAkkTgbmU4CdwyZTeJCFUECi9Iik
UqaLpZYPN0/3MVnuYWTjAigQ7zPu3i0Of+2U5B0Bq2pc1RpQW+UKbc5gNyhk
GWcIxHaZ9P9W3xcxRM7BqjDCEi5MzYMc5ndoxR8PB8EK4eSZ33G73JmAzXza
6tDNIltGzLyWhamyK0QZmVgme187G8qZLeWqd77Fy69V6PPgUt6R3m6S65vP
scr7smOq+M48i5NUQGYUr07xJQoTB5goXaBHzESaYey8ZYWJteaGjDfUwn3Q
arfo+ToBwMmh1/55/LvZf3zMl48AghHvKWdrpbSiKvafRjDxcH9kK8DDMUEU
M1r8k65wbNUgWbpNq7Z4p3dx5v1XW097RWR9Wh8pUvn4flq5eEiyKPQtdcIf
uF/KoUXLN8+nWAqr9uWw9FBn9842f0tmBdEKxHwyG/XnLSViiZNKWBXnm2SV
XW3v6ZeELRDOT4Ge3q9rfce1Okw3RAqaBcfGPgt6XlTE70PlMMerHNUvBCQn
Kp499MjTI9QqLYYaZAuasuTpxG7UwjpD/I5AMch4+5EWlh1CoonPYEeG5wTe
c9TQR4XrIJ/jrSQgRC2OI8ObLGRmNUn//yGSaLFe6G71PPA6LIhBw+qOIsxr
MtSymwSXh8xstEx1U/umpXiwDhR/FYZs0O9GammLeGIcRd52WdbZ5FD8MOvB
uy/1pzlNgv8bRx12TLGsTlwGv2GwJuCuXO5nlXoN8OsnbDz0/pjECALW4LV4
cCat+giwWWIy1UPAWCuCrmTfqXTiTg1KzmHfdebR/eb129c1uHtCyFURpJXK
jv12+GCm0D3ovG2/ipvpIZlaB6axaOPem5zTpRir/sgpTMqZ0lQSYBPj5n5h
2IsS9bM+E0XKQ/ozokEKMtJxDsNC3m/9T1hBLOgSxm4+n5xbuRuus4neK7VY
afpL8QptJfi8+YrrYCJIRsX1otgAm21HQmT2v4OPsR68fEnoxo+SjqQpM0jO
8soPXRwTdPmLZyC/+ICTeMyo0Vpoh9yi/4DEcluSCzM6x1Vot2z1G0dYO1B6
dRdQ5eu4wSs1i9a1YpJCS2Q31KBCJsrI65I6pSAELmTn8nZABxtZ+1/sqPTB
AGj22PHTt4h2im2hjoeumbh9r2hP/sVsfWC1L0HH3RUkgmH/5BQxbCxYIjF2
z51F/6ML1wXPm+H0A4malBMSfYpLmV22Lvqn8lPgNonfuVI9IBcUnJ8it2H1
Jb1mFtDrSNZ0a+aYw/Ur3+DIuXNrI4k54BoouWEmOMrosHShmLZHKImqfYWG
x0ujS1+EkV7II9QN6FA30x5Fez6HZkmgJ1fI5AcaoVeyM7Y/8WwLz5ytTb2s
uMQ9jp0J5yWjISp9mOkE6AQhXwq68chGRU3FwdcgLWMrJ42xrMZDiVgN27zg
nl8IYqSnFy0et9X3yKSCVyQj5mzvOTEoHwjKcHuvORyppaNvRuXe8vs0Tr8w
HhJRRbn/3Y5er3D0BGRkxTnp3QgdTdd3jPOF8foLyECnVxfiAJRQWZ6RsB58
sY5HPbtmsX49m3w5rFxxCBM2WZsZWN8xcvlzPhb+NczpZuhO5KZwQKecJ5P8
iDSZDfuqpdyULYejrmtjDpzA2j6tmboRgfC/ceGsdLFKmSZqGHLJ34Epcolg
f8OrUVfDCwdyxS8+ND1ZPswRYvdiKS4EX0PNChi3c1qwGwpImbrJek5N82nz
vVbAFOz1o09XyG8+e0D9Nz+ldjH9HtmyrKz6S6s0opoEVaeCJXaus7b+0tUr
k1nkQX3VO9tiZahi11JElMokwQ86ZdcoBkH5Yt5C9UMKh6RNxJB8y+/0Lwt/
cSkv+BTaGHfH+AB7jRfPFRF/lh7J4ZQk93cFLW5fDB5yARMONtrgUlwhrLAN
aW/9WU7ZHk8vgoqflP7k4FabSuL0n3jzXBJMVldUV7/u5dP0G1LFPASylVfs
T0SfQLJ8+8t1zTmH42xE5ykX5krTfrfTqdTqLvoTFrUlVJWSMWh5xxCGn8ka
EtasKcZRYKCbfxXN6FPcUi+uGSQt+fvW7mG/Vs4cejCpLPEi6m0wC+k37ksS
vHVIzfY44QEtGb/RziyfCdB+2RYVWtt0keUulol/uVjAMEFZ8N4kC7xDWtSB
/WiFIFQ9LMYW4fWJbd/M9suYeDJP2wiadH79d2ebPiQib8b3h1PH2XhB7nRi
+zgTcziOBwZVp17C/hHjGajlrQR/5uK/x3I7lvecPuGAEX1xxD06M2xCICyL
jTardfPSUvyYv7FiVmzryEkVrArHoM+HcOfXOr6dYbsHI8TCIk10786PHH/y
RrUL452CwnesQG3oQNlL+p9j7+cTvSXFL0FOmW0RkVsoYVPBOhoNWUCI/W9L
O5FtEMBtCa4P/hVxO2t+3QugWmWHH1hI3UPi3+JdGwYAJUeB5jKB5LEPSf+e
5wX9WTBzJ34eERZZSouWy8lfs47y+1R2Lc+gToCFn2lowKkcx3hx/UV7EqQ8
5nmLzY9Yz8g/mG/oG1kKEZL6Tta2W15d9qKlnbeHyrkrN6T6iQa4rBZPaN7c
/SzyCF42D5tQQbj5LcnRlWjlacNW7xJgN1P8QX/CnBs/ogVQQLgviIe1w41b
S7p7Wy5FljYAVSyR88eUz3f/Yq1gfZXLaW6dl+tgb9zJrwnRd0vBVC5hUjO2
yUWP1wtM9L6IK9v6hSlXWwulHBpQq4Fh/QaWkfAAf6cbRaUkAJgFSzC2d5VX
AQeUdVWNXN24xwaR/HNzEdx3TzgGLcn8rmWeXjT+G+eRL/2kqz1sBOMbIM8Y
GqzIndMGBOXFRBi23gFnUWG087nbqjHQ1OVX7hB/qevzawlj7J4IvMKo8w6h
tMPuBCXMjkMwJg/Wz/xkrZkgSGAEDWc7o/FvEndJr/oHtG9TovyM1/XiXGXM
nabWDGu4lEf+V5sCp3fy2Pe8o8hhSVxnSCu3ZxI2Bq0xwDt23Jx2Y0tiuzbn
2qg+xrlhdRYeo9X7E+dtfA/DWBKINk3ZJNNjXbE8sU+A1/j+QCLTVt0OLU/W
2nd76yBkd1kHTyKSdMTwTYqyqhDkARCMkrct/aclQN6Og4RQBFZ4SJ1Be1MB
CpFwl9adB7/a3EygXfCHSa1czwFLZ2U4XiJ9UyyBvNiROauXWSlsUiui+jGo
EOgBOOGdCVKFlChIwHjjxlG9BYE9qs5WhM2u/0asr7npOy4alRmuedouektm
L7N0IY/f40wa2REBsUTDG1t+v5AlwRR006WPPIyYKqX42jiM0lAoZAKMw/WG
XkTJA+Apd+SDl8InbeZP++ojCnf1EYb9rXgEEx4d9lsVS3gDwcZIHGqLa5E2
TflKXZeQnbLeEgmvk2WQIzJPLZrzPsSRPH8Q/0opsdYuesfYqAg65rDtigzo
J72xfdAFA6KQnRg1zPKBfh1gvF/10Giff/WkewSK5OHKartfMeR6d3OLYs3l
IAv5zyGhVw8L7/C5Hz7O5YNK/xwf2fheB8ANgiVyNP45h6OriahqvdtD5aR2
cE2XrQr1wKScbMyVziCKUZ89/OFWpRcvbu/IAgIjmhuEmJ2uxDO9lw+6H1Rx
SnNHREsqlqxYZpj/AvKDHzU8pK5QtUFvIC7mAJI8Wlbhchx6yhcArga6FN8S
cx9X+Eq8zzfUGS0iWH7SVZQftw0WPKyW9BZNvPWy4uIfGwo4TY3p3A7dMsK7
vot+4G5dr96xvpl6Rkas/hTDDFcWCpIwpdE2E1+UYizxD1+jJCBoWPDfOdpu
maEy9aQBHb8guL0nrKyXE5u8ZB/MXh7ntQ3M0Du24kvxr1XgpPUfugaTWlZ/
5kXEukEMZivZcXxNvFrG2MzCnyEDYMSFG1i/TcNa7RaN3kt6edIoBe5P5lye
lVQV2s1CSKhM+m51Xf4TeYDmG5MOoY5BrOyiJjfPOTOdaQnawhb4eH+qNl27
VnDND/F3kflZMK6KBCFuGhLB4pG1+jfpAzNE6OFUBGo0CsvgTQa4SLuek9ZE
i3MY8v71gEe9RvqluUfEuT6BJP3aUxWHOkUg7cq8syCyZXEgsPw6Qowtn0Al
a8ywQUAWqD5nSyTe8/qr1sK3PgIS33OBnyAkFW/z03a+FjBOFoyg7bjEkKXz
VojQ8TlLRusMq/SnX4zM13XvaVmdFFAomw/k1gUcAvBeILeg1JJp//uMpJNZ
E5Mqdfy9+p5BCDRhGCNS+0D+g7iDvSdymMyLShRYVa9wjs4eP84/c7OZPNL6
+EaADY+uIwCwhJwWDo/Iz5BkFMdQxKAnkEoWaBXk05elQpy+CVcx4hLSSpLr
cuRNAQs6UQTl7A33ZggSZ4SpN8jKYLKsJCDI6YO1WGpUxIYH4HMDrBxHF6eH
Pjh7l13e0YRFj6hohDsSw35Zouzt0wXrRUPVM+YREZ7LI3Pud7v/QUZPcS5A
slvsQW1zYJZuM+yjX9e0um/gO0cZcpWWO+jvLPL0c5E/6woDGs8aZAXV+c3/
cv3h1XElzqq6HljYe1pSO9sz+VEV6Do/k1A4B/j7ERO494s2GUxErEOHerrl
P5NRo3t/VIWfPAEqnkDpizuGyq0oqPYVI4SpWoAYRnL/PjZSJWKJTDNBOCiT
ePMG8OWU6fAAv/2spubTOHIavH7hWqALeEBvEsghepil1TXidcbQ6LfjC2nM
c630nsI1HhVfKENK95c7Dg9NY33m3RWfnqr+T4fS8Eo8YRio2BAYfc6PdgGD
24E+z6hfwzBjiGIgehw+sBQUtgRSgEP92BtdDMr7U1rEHIG9DHTMfqlA4/mW
dxZebfJ7W/14NVnmV0acWiHqLnJQiXqueGqUjCnve48hjDJopX2zDUVetVWE
XLItymKqQa5vC4mYf+u4yo76vTJM2GxvXlC9tR6C255sKgEfpbWgWUq+7Lc1
VCGzS0m2Y8kD67ehnsu0kGX30LLOP3S9KuWhR2SCw9WkzveEo9KAJsuopNHf
Zx/AlU824b1Q3ChLm/UCWT7QzjI4nF5R/IPSzCVKuFqeqooCfa32kpTCxjq8
ZzhXmC/F/9QO4J8gjmqRLj9U4MznXwcCYwwUuHBzOeKLVgaaIQKIIKI1AhC6
yDtp05Rh/EEi0qzMndbEAK4YzgRWzzzAeU+OxrbeJDdmoPPKZ9a0oKWfy/sf
LKa5rgyZjt83i/bwydwJOO6jitdrY023iK+ReYK55stpv6bhW+GkqpjvfZAS
PRTFo99EpsKlA4kXynRFzBBWHwfDk8CiF38SYhmtjDQg3dubCgBDsIpzbWsC
AnkLdggVqvysSzesWyn+6ytg8U9vYogo/NvYM863dsDXBkODdWJJrNeHnU7R
I9qQybmlP69ma3bv9vlbFMVdhIE9kvlrRohkr6WOil8htqKlldz52r4iMzL4
MNbmm9RAwRdiz0/9MKI47UDPsZqcNE3AvYW2e5Da9sR77wEPgYNZkdHvp53H
YIdbVM8ZogxxyOw7wA/SEVqiPp0ha95BiIvAex45c2PdhcpWV8HvUUnwx56B
y71NsEe4+vNiE7e1Q7M6cDmAptfobet5J60kLuILMQ8Yo+gGmYV7c9U1enWv
2hPpssqln35S8TQD3oNeH7phBT0j9SGMWcjVgA4/hz2y+mc7lNxLbuN48x74
NVd/XgGqiRtXKCRZe57dpKH4Od71/EIFMABg3YmPRm1QLzABaM+Oyh1NoC9Z
gEaOH3Z7Qai/vCwHMcgb9fvJj66VRMISV9Bnukx3zex84xpwN2w6HFsLlEh8
oUsgTeJ/jG45zrdlD4eLDVbp/ZaF7pM0Z4k4RLFN5PEO95uH2eqN9rmtROyR
eH5jZOjqwPSB/kzNGz7H1rIVS/aqUVXFDC8IBJ9oElvqmSp0mZbUAHz4pa4X
VxVVLpu73f6AoOOh4bStgCQrvOfo3VLeVMsBClFMurRxHNxX8XHIuA5u5nnl
t535MCPBehd8ZO2zFEowSaCldsAjjUqaf2upx37WBowzsF7bkBcqmh5V/FrH
0G/j8K4hJKz3WawkI1iucuSw9xQTRCOYDPOrS3SM3A6jo09k/vqFb0SPwQKH
FsOuw3INDAFA7NPFnMAafebYybUnkQ1H9mr6gd29lIIG3aWpNsUjNYs8DDUM
MsBw+pifAyKEv5Q2TauWq/yJVMzuAwGf0zrhExzNPZlcnfUuTdSv1Rcv400N
0u83lmUyY3BAF8nfxY/oPWQmlKimyiCv+OycYXD26gg7RMsf1+7mVOlj2nMB
ve9sOSrpY6jhdwA9E231JTAVbNcObcFh2JWG6YKV1K1D4W6b7nWhGQwoZvEP
jya6miGR7v3hb51C+eHPjqraLzV3tlfJXV3+7qju3RPX/uyC0kwyZSatm4sd
l/CsA6vyJVfbKzS/PQTH8IsZpQCf3cok7XqQsrjrXzHevP6m3tVVT+sj/bW2
Tv6G4o89CkLLhvOckUBqqCt3BPiv8222lkE7aAGOe5EpSmRdCLGS4yeSasAY
n/dWkMl+/+fiajhiicGtTbnt5RkqTy1yZVkp5wXHynYu/jti4SnRSmupSQhZ
MYQBL/M/JRe2JexOmCBsXofioPE0pthqGrTRykPnKSJGxB8Enm0HAvRk8D6d
yZkkHfccEOiM1UoUyhypl6xpQBS56IgOvsU1ZVmoRITowpjSORRQyU/Et3e3
hcu7sW6OlGzlVkBwopeiXDasX1ocyHIGkjPkkVkF6IcBmtJ/ZK2aGOdPrky0
0jpWCg+OsQyUhrYOofIs0PmkOX3YEoyYMwBaMLXs5cL+4rMN4DuZ5Jlya1+I
ERZ7Uw+anicCHKdk8g+nw+99JIHRPVSsKzr2ylEXdcLZtY1O5GN6sUNufVJy
ec0wYmZkjnfJ14vrmYf8UdUjLPEq5bn+2tgAIUs46ZDbTzBrqtB6EmkX//FJ
nX3beusVLbFYyWS1mUMQUNLVCUFtiwYvTuY/9KJcpedwz6e+de2wg6K0K8Mn
smpA+FqKj7ox8CV8kcyjo3X2safYyJx72k/5SwRcs5JfHwn2uF3j/uCjx1/N
CozuPeUUbLtoVlV0P37JK9Y+DzsCXXxKgVford5XDS7763MK5zv0uKDeYT5R
1RaGV3J75H/U19ctM0TTdhIKsALaYYcX07mVSPir73qDTZcuY9NmoASCNmFs
bl4DVA4GVMc3j8n8GgS+MzHjxB9KcH9bZNjxrDddCOCAqis1ThC0a3+P41pn
GJLVwcSHxsTO6sg4nfIya2fQeXK935D0admVQ6dxe+QgHoafgBZqr3t2rieL
b4WAl2f/nAx2h6L2K/wTzMkcs+RAc09xlGG8RYmHZgrVmURNmlsGk8SkvKpb
WwbwPLQ+iL7Si1O0Xb+bJ3lLDdGwnNzKAuZbFzb5UgE9aFOUYNGg8s75WLCM
njNG9lxW2bHEJQ/vcl5SNM5MB0cju9hQ9V/ZD5Z89GVZ6tgLrA5pgNTVUGV5
V4GEhScSiaNpY8VNpRT4VHmf4vLUci49tUCDVStnnJrK5M8J4zQOVUTGREUd
DUliZGd/wgfN3wpdCrhUW0lMF+VbZZg9KAE+OoLKBFGipGdIyzmxBAjDS2uU
vsFmTYFh16BwN6fGxhSE3vZf5QyAV8jTZOGMmj3nRZnv0ALNQjAeD8X/YfFF
s4FEyYsRnnM0+wwNmpSsZb95sDrwnZqjCK0hdUp+B+a8uQ+/Q0HJTH39lwal
yfTg1NmmAQIQJCRV56//Htyc2/vinmu7vlZOojll8aAydRJGumfrcSgDyk9Q
eCaCAQ/Fzg6X/kycP3yJioQ3yrPYJ2GycTscoxLTh2iG9rxjIeuWBtdd07jK
HqAPNR3eMhcERYo995EhWSRwsr/LTrrI3c0ab8qa3hnZ4zhRGgE47XiMLYAV
rt3A1+OQYa8yu5NxNQ0PCK2Ag32hfHP1wwoWEEWaM05o9b9IJe3Q7oVtV5BV
RineGcty7NL/1G8ggusV2gm12UfFOiLlD1a2GJu/iDslAwFuaBtB3Auw9W5Y
zrUWWY6O7q458+w09OhQUgXUYi5MAYOOoSBZ/GrSLxzuNFhwaeX3XVbmLjGb
GldvVfUIUjLnEN8JU6krIqlgLbTwYKT97I6NGzOMM91k/C8uInOHKl+3ZtDj
VIA9XWkJftqvXvRnc2sEFGPI6FEEYb/r1yhgmQOcN0LRNECdH/7rRvRPF1jj
Xw3XLJ3EyjFCvsTRz08KnUVd9o5xfFVnps1a+O1Jn9DH0z97wGNuHa4t6riq
pEvpMxv1Hm59K2fuQngRzyUabkvfmVMGXE619bDURahtfzFl9ziyBQTJAJSL
IAdNgB+L39uhJF0w7J52SEVVO6Zmm7dtiPzvktaLpCC6QjXUglmCJU20MmZH
9DpHIujBcqTjPHeCix2HtSWyt+KHiHzQ7CmF2C274yS0klch5SbQ7NRCb8bj
8sdjnU2foNfG/GJOxMpK2pnjcWeETml9cSqXW2PEon+VmM0xa7JNlMHAYqly
GDh3mabxKK2jQG/y+nQgxktcC5D7EULF7CUdDUk38wMlArgEO6/FDe99N7Ev
lvXj+qBehMzy5iLySS02OqQgl1rZRHGj2VVKN8q7tiLQdrJ9SY1YI2H6BERn
F3y25z9VAdC9FbcouOuLi1WAirY5YqnjSfZbgJqLKfF+T9mpGbOh9uz3Tqdd
5DGQdY+NwENcrtIrqT2HgDD4b2XoIcn5P//SYzvG32UgXvFPFW7GmPiq18Xy
Qe1lFca7taoFp5rvdfk2KFg1RahTGAs067kvkkKuAoxzpJIjZIONLgnPX230
yAxV5rm2DVBtOj+tfP5iYSj7gaRSeE53aDM/+VR+QZteKvrOA3CmhKhXxhCe
nNiYa0UHY4BkYk386nfCW8qjfwtxJILI3CuOl/pcCUn4+orxfHYzYg5vbTx/
iap3AP7NYDp0iI6orwdENlxfjzagSBF0BSZg1gkEMx4l0QOjIlRc3AECMMfE
P1ok7rgCGjL6Z0zVjyThcDmxYwiIkfdqsWNDDNmtFg8bzbdZQZFd50GJ9Opn
o46v/sLD4VTF3FDYSdUBuLpzGCSa6FZpVqc5Ef9+4+BMyqQG285O3RlHj5OU
SiULXbVUv3ORvXHUfP93g4MLvjcIj4wU+zQpB9H3HYczeeUDMp3UuA8JzCB0
rh9NJIu17bAfgy1DKus42Cv/uXAUM3nVJjheh6toViA+JMFI/gZ7CDag+MWH
nEjhMQLEYd6bULwf2a0R1Vp0iVqYHtR1DowpX0VJ51P+q07f+sRP6GkdMlxc
0CmbbO0NmK5G5DNcE5QSfjrgK5N28lyn6lcqC7XFAXEJElZEGhFPHOjrQNoM
/fPaI6Ls4vxUOoo0XYkubEW07UINuKAf6TrYSCmWScRXvntpectXPqeLx77y
wndrk9ROWXMPZDD93jaVkTG8Nsgcbex4m83XuiPJK40BBl2xbiTgU1YNQGkd
Btf1Q02kVsMZvxwtbT3FuqQGMB3EDsndd3g9xKuLtYhRwCy6E1LYPFCy5yY7
S2ojwlvaUyraxccugvtolumk6ecfb1SLfeiFOFc0typIVCv23MfSc3yjLMZE
r2q9Lqg56cK2u4hLnVfrGuPuniQs41KHJ+4WjHZMRd5hrB9QDImpSMNSJvWp
iDmBF1IsuaNrlkFp43yCByIyDLvxWJ/cIJYlVRhttL+KYdbg16uqDn6cLj6C
srerSMm48au8lPkTjD2aT6wlo57ifSOLOb0pf5XO9Z2D3veMsj38at//1xHb
msgBByazzLoSF1MnKlJxol0TZtzKagEJ5QXDzsdofk6R7UJGn3hxn7xqSl3+
nWrj0MSojRQ8KQXnvcJqlQNfvUgI87e1+1Z6Kvdk4w8rnIymsbRQInOze0UB
FB9TakgyyP2e6E2vjRcmWrg6QW5QkKvWaMuUUbnR7CpFQ8JUWqNhS0h7gTZd
FfnblGIEREvMo+bN2gksNOxDvs+1pqiCUOSlrsLB34aelu9lsRB4tTvDeqpc
2v5qeGPmSLFMgjZuSMQlHWbOEJpgo+THWoI/yBGOfwOJquKp3y6MzDii5CSD
KFkJoTJaPTxXOajzIA6EyFbkHaGOvVQIxlpVUegcxe9uG1OudODo4FO1YYgZ
dB9oLa2hzpZJw9+/y5zzkdnwpTpiInrzmvN6KJHizBDKe5KY0GRqaVH8C9V2
Sqk31BY7M7Fqd5pmy6Br5tObQPm5F8H97IPd0uBAbnOaxuPuFYs3eIMjTSU+
Nr7smU7NbkXnXdfjkUzxa5exR5+i9bDOnFxifJbVCi9it/u/nTEnwa2E8zK8
jGzHeH4c6AfgFra2fIMSoUWD3F7gC+Xkji14tajLHo48oMcvRjSI24cgtx7J
f98OltxJORbYtt7RLj/HfO63/IqXjHL0K6wpHhg3Ql6KmvKeIjcka6278y1b
g3CVRRZBuvigzEndZ5fBtdgs1f+TUPfjCvwBn2sizhq3boP45E8NlX9BUqNU
AeHBoxdfzJM3R+MTwrZXN2zqSNHxaD23y5Jl5h1e7+WQFC+Q+kiFZA7snbO2
r7DA/6zVuVVBEGPRSPTo/FAFC+T+kjzs4k1qWEr2yj17EeMdE3rFzPB938OK
SOXiGoegKV8KwSMLB95HXKKr7p4BgV3D914qMb9MWGEzJwdgRMmZF7wPsxdo
eT5x7ezFlEchLOYVIx0vESDGsVKWMh7xlnMipV7u3T58q+8Lu1aiPbh9B1U6
7R1Ob9U45967CYom+K9Osakux+EGfqaVnwQnZICToGgI7ZkNkmRgl0TrgvLK
+66aQE3FoYFJ+pjqze/NWWJwWgU+Wd2nHYTlS3unwazBeiGvVzGDySl1cNgF
ayafq3Ldh2wpzG98ggUP+zBrO+IsxAbwD9Be6CHltkeF7epHXlch+mWZpC7K
LWK3jzf3NrDPTjhWrYx/rLe+niFedSgv/gHbNNe3HWJMaVfNMmPEg8j9jD0A
mMGp7SHoMTzIIJ3ds/by0JYT+CGea43mpuci1GFqKSqWUT+nG96SHcJSpaWo
k8xjaYbEOwnKtUGGuAZOgUaVyY+qk6ewzd0Jrmw4pZvB99J4H/2SVaDMces/
07w9DsZvW9XBY4vgQdFPB7ES7Xpao6IjF4m2ZwDMyBJvLUeX0ef1Fh3HntTM
NUnaodnVsnfqRIElOileI+U51zY07+y+i4UbOak5ac+YKuT6/yJ/RvxoqX0Z
CAxsD5gtXZBpSAkM4ktGTsY6uHIb1pyH+TxEGA8P4qARlZGCPHAwY8SxGivQ
tHvAvrN09yJcw9J8nDqwo3fewD3FR9z5GeE1wDWFssRMPRkUaATAXHUkg7q6
FQBm693r7R02zakTwcrFdPpaKAEsBHuSJJOsCfc77Ug1WUTVQ4xsaPwv5FGU
al5IlLn2plBjsayP2OJkBx/YQmfZ2DlMMwGU43wrut0UCL9ActZG7r8xHo3U
u1rV9CRh8PXz9J95fNPBpu6Cju82SPrSo4DnqFCFffvgusxjPf22fU8DlAuG
mLKpy1zqvpOXf4Sbf1ovkGG8f2ffsbelGFSJm+1FEv7a3NK5R04/i7ak8jUo
l/gFWU9f8qmByEYgivGLNEt8RH12TL5GbYt5RowiQdJSNMXoH4EA8tNic5Jz
z9t+bBZBYHRwHhPnt+oz6tHbsCATQLUR451L/JarT/EAkVpztuXx9xcw1wjH
2wJvjpRcAXr+PTrTg6LEX0onjp69njQWSV4XdgzBiqUOLY5us9RH23W2tOhg
oFWDFxpFXoZMjO4Inz+4pGO6qwLMmC1Xnze9piVWKbBaMsR48yfoTJrQRHTz
GnxsmDVeXCvWjsODbHl7esPscrO4oEGR6ts5C7SJjR+cl4aD/4nzKBphqrQ8
JvpANQ8WuVsOJj52E9JhqQAE0epHeTDKxtSItUiNerZhd8KotmZiakxugZ49
VBfjOO2VDUJCCaob+3/fIjHOZmw2GVXuEM0o0v+OIP68JSvv/dt6OTdp4Krh
5S/QoSb+LjQomZEiryBeOBkw3avvPNTgrYQbF38b67KbDzYkW6T2hmsvbJ5t
nAOy+OcfXexsRXeyiDW/Q/qv4m8zfADv/SPH+r/y2qebyys78UMVTe1Hy3ZE
Nfbok6y2Hfn3wGRibcFfSfWr3MctF1Pw7aLbCot7rG1MKM7okWtdvPhAjFTB
bJWghDvZnBB06hpBs2o/wpqPk3O95ShNtwK134/BsQihi88B+BTX+3TaYwnZ
jPyB13olK5Xd6j2hya+PddAUoRehc+rHveIvOqBe1vnEB8QVpjmhtd6NzNSI
DGBC4acdazA7VORXq00VrhApiTCV6M8UNbZ8/pmRmg3bRkJy588uKpjbG8So
eUv+He6FFM68AnZyPmPlGVzSYhAmf76j9tlY/OepLRDEJFM6SnNHbo4lTORe
m7kh3RwuGPojJiLJ0GCbb6acCXuSoRrCqWjoepn1SxRtzzwq0lzP3xdsmkyo
xGUjzwljpsi47msppPaD/L9lIT/HCdl6SMcqX665nhOv0nH7F4k+5ub+LNWD
c8b/nUZw9AbhQEv32w34UWHoolro5Z5tYfNIl0T6djid6pPdBhs1f9oaLdv1
wwYyFXe7DKJTUWfA5JdM2VXBhk4T3I2s+f/B3hatwAbDQFBRpgkODz7SlxhI
twZSd5EAGKNCVu+0LzsNuPKjcxVa4LXLuhHaPw/v3CfTg9Hzg87AJrJDwYe9
2c1EbarC8Ma1QmSI9UANxwkwIDxEfV4vwmZ3hPrNg5XJemli/lOVVV/rFo4k
IPR6cNuTdrC1Pj+Lc25b844DH8w6z1NKIuPfd+FdzDeEGGkjVZqhhQFlmLel
4MUZKHHXSbLF/gmia6/DuUxPvDTqmpZmPhEC9nYM3doviFeQ8ZLYa7odHJBq
P2FhYtsfq0Fko0cbv1aLsJLF790tFSdLKNqB38jNaueHhmgpJiAE9ovzldEJ
UYy5n7lAqBYxDG3nnJ1Oi932nloEJaUqPO2Ykc6wfHXV8MXkrg5oatWJdDNP
2P1vvQKQ4plEGYNA/GdT4KFJRSPXszLfRciDcFSmWQ1tcyzcHYP27Z9RDSiX
xYp5+MLAH2pZMuKKjaqxposVkC8n+rtu8yDHiemxxPstCAWqUEBNs6/eBosf
XHQkwGKX+MAO8sI5XtDYqkRd1Amxr6sRTTYNQffrl+/05Zxz6Gf7im6A++xB
tPi3vzDJskZ+T6XBWX9D8+CM0MvxE8z4jmpbUyfcro2O3xhGgGAAgIvmuf1e
81O6KrnQs2Z8fQ4XxbVgVCpv5QImdFF1Xs8OSg5iUIMOwlOKM/oDoEzrkMWB
sYuIMRbkA7hVfVftSxNuLsxKmolaj4wrxYnEYca+a9blQpo5UPBS8FWIK5jW
gAsyQAHUN1gF7Z597WRll23cZTJJqLP/aaoklTlO3YQDHBDb8vx4dLl0DKXV
tcQOami20aUfsTfpQJDBYSidK7htQITtosEnfLEKiQxILFCJkZP5raREJFUE
XpWSxC6bLLEBsmqkbpWHtFbfmoClDIgiZis099C0fn2n6W0t4/qZotL+tWY0
58o5IbaD3/9B2NpnzxokrHl4RN2VcwR8tdgWpz1ebyU5jNKYS4RiRaffaggf
ojKYr27sWHcVC3y0nquqG/pj4XMvrlYbZJA7y1QDFn+FcwduxgmkdLz4fvOE
gq8nzmRXn4yxU47iHhjz5kqI0qoyDpx2QSc9EOQOCQpdDgHCzvQevrlqa3mn
wV4sbi2j2RZObrYTjaZSbZ9uN8tARZSCP25h6z3wA4BY0uTqgrCn2oLKo9G2
5NqMHdfwZaTPsjCGOdOjb2lPJHvRLAgh0r65RMat9LEFOT58hZ5EDXe7LPdb
d4Zo/DWRVafuLvnoVvqcSJvmb+tQ/xXqX+S7yMaPfLklJua/RBT6IS5b51gw
SLUozOkeCrtL2zrMHMDsZzA5xm+4gr6snU6yDqULOMme6WbrtXsdObVIdXfj
t3q0ql8x9J6naeuv0NOK0C4j0kHGc5zV/0Rk99fMw3hChrhVVnQeIfHcquGT
2rXhBahl4jkF6r0DEeFb1VWJ61N2w8v9UyPJ+nQ6aW8NKTQCkRB51nBnDaJ1
RpZr1rVXho6rFrU7fxuM1YBIJ3hP9P9p86pDzZPNyY1ucIksIGmsIBqi494i
ynP0suBpXatqJsdPpJQ2/E2noBQKQLEFs6ZX3p0OVgOzSj/uqume2cVF+mvc
jOIryakd7rd8wEcH74Hkjc24MiFWW2ZJEBf/4XeJlAdH91ktw9kIO165iTCL
y4BkeAVCZjozwNuUDSFpkusnI+r3gsw7QcGRxeQ50y6PDP3MyG1RXOF4UF4U
wNR0P+7fx25OzLYhm36EYD+LgJxPBRb7+EoXUaZ2DCnXwDiFyTXeGOZuYtf8
M4PmmeV/lOgUcL/zBUk3GMRZK/dblq+8KxdDvb/dr90Qz+Na7NBwNC+++hHb
6VNV23WEDrEUjRlAxgbwGT0/QruTADW/MiWAkDM/a0z8u+Nu6ya5ghhbvsdp
HL2aNOOE19FAfPJbw1fr0jgGFWhj3tWTsysXP0s8AAQRzOKIXFFnuwCbgo87
m58wqh7dPGJJ0mI+RaSWc+yosUP0iybcgF+8eUmaA8ljwGkFELhN640A+CXs
G9zZOLBQXa4a1Lhmzecv4C9MLCSeCk/fOuaiaAS/rYdaU/IfL4kno8r7IM7M
sbJmkg3FCe/KDobNDD4/PlUNDvzPzAN54+hXD78EeU9CIbqtNEgBcv/SQmWr
n8LG63DDbBrHshnCLLGgJM/cVff6UWJG84wdSBHbgWLYTIT0yZVjH2Tdhky6
WLNafK2ETQcwVmhVkQ6V3Qu7VKVJUT36mRNHf36hvApm40AbYRJIENhLIvVF
YD/le3UVtXYs09qp7VzgSDzB0BhUvWUFKKuKv75AUq9Hf58xb4mBe1nRBAKK
lKQ64AyrctF0rB86RT75vdHlFZCDuNKDXLr1EbYhkJVZH8te5M66GbxAZE4y
gINQHo5QiPuVJUBop0TRfC73SpxMEOc+z1qMIVhWRnRz1THICN5JcGHEyPu5
U79vKwq4LOHGC24pLc4RjrZXiFpqKsQ/IfF4dkNZFuMvT6B8SiEztKYjlOQ5
0wE44HyrL0iMi8LgE6RM+kK2TDZQF41Dl5I6LQ1E+/kivqaGrHvaquX8faoH
DRP+8o0P5T3GAB21t1IrPHG+Gd9MP2PcU+r2FgtGXnnZxSGbPqzOqHkTLdx6
2dZykUDpy+fyO4V6mWTyZCJhVWxw4l9CcMP53EqsD8Z9MCt5G1NpEXK7y9hk
uBgSzYajUOY50KMJH4MQyne/CNRs8GP0pjRZZ9XTUCGKvGxzLWWTcvuSZ0Ml
j5LbZzn56xCfqhr5KpT/ScJlnoMDyk1ny2qMvVtFwlvDsxeJa4pQzq+bMKcf
P55R0Xpf87YQuO/gqxuTYpuA2EWKe4wz5XzihwJjOHQ+D+LwxEoLrpg3rno5
hptXpUwdi80BUKxm4dS8Y7Lk7W9q3Nkoc6WPfKa19+aPIcFL4dTEOAmsWQff
QB2Bqn3ytisjoYOtAr0PvUt4WrqgimNbaWDqogD+pyg287tgeczfjxUdICjD
YbVOaKrXlp3EWG8ab5b3Kff8+oR3u7OVeelb2atYhPKCPtdvTV3H6+ARt8BD
YmcuZakV5V33rX7v5ty7T6tq+lUwlWRkVa7XtIi5d2Y1z0vSKUODtzlZUktP
tgI83p+XVty9f+0NR4iCOqOs8pyZni2qhXe2NX56m4C4crfIpoZW8XMnUhN7
wKNHQbqSF0G+ZJrIEjnt9cT2kZXa6N71cFrYph76QQnU6O4rcA6Mwmxo8o29
VofRvvzPS9m5bmHsVGOwDisHqLawHTbjstAoHQ7Rm0wWnPY6qwIM2Ao0FkaD
31EWhfVYoeXOrT/qw9L22xjc0J3cX4DEg3vyaINci49SshWuNcZoMRkYnRRz
zbMzBhmrymR1wG2zJePOnsBUAtDWPbQkY0oh/1cGNYqnlZHIhBeREZl2ZBoL
y5//iVaQjroKo+NhBIhhD2aYjDrIckIAdsDkYKOrLMiVyUobXLkOuBht9edM
9HkiwIwDOGeSefW75+AOiZdcRFLJAlwfJ3UTtYM+P0a44aa2wABJ0jYyp3X0
1N1a1eVljgUH8QaeMx39IlzyNEjLMgiQen2MK7JFPKMnSMqcS3Lfen61C0xH
myK/KIJGu9Q20h0s6uhGpHExSWXQFkrcWPZoTQyhbjNNVqHPO8Vx0HYraxnk
uU7hzqPEIsa0/63WqlyAnACWa0VEEIb2dyiUgk1B+wtAvclCkqzYLGOLGpxK
TBUYrNq10wToQxNMYhSmiBnb+v8tnFVESWcVLowNcNU4NGszvC6eRPXrXW8B
stsN1b2Hv3FVKoYa6wbRxM1HflZ/rinPn6m83x9gJ2yWi5ClnuiZ9yG6HM6r
MSsHmg1R6r8SuMbuqKE6RSlVI+xdqDtmq1+cT8Hd/43kQUUcEsYapJfxFOhb
lqW9T0OWd7nNvnFa8F/PAehWrT+b/2dFS5C8jENZ8jaVazT8vFB/BZy+8QzI
+iIXNtNieKYDUhVPr1ltQ3p4KTXcJoUxCrqmK4JhizZvQeRCfocsIuZZW8Ee
PRKxO/slU4Za8U0NL2EnNG12UV9Gl0nFBuYf36Prh7aGC8UA2daQ4uF8Ki+T
eNJsexGu0pvkHUDJlpDbx8Mq6IXtTKFNNzzXyoDrWjYdY2PD35qKdcDsofD0
0R1APRUYuuzBCkBoBqSYhS9bHSGRqaq9WMox3i3m7SqHRmnFkP87ffkC6rYa
y2KqPhlVeH+2AxqIEhMgvUaZEax/XKJ5HOvY3/1/Vjnl7JkY9zCT75jUMoOH
Chk3Si0xejdwEOeWOsXxJyvA4GF3A/ZqmSskHrw5Hv2nEEuCjXjCDmtHsjGf
z/nWF36PSfxayeVsPgjyMHQzyMGxAGUeqKqOUMyjWIN/fm4btebE3VZh6bhR
IeZ3eIrfhoUXU9+eTYFULt9ORKdTvjEAk9eRnhPFCNykZU05Cj2Z/rq7esBW
V+CeIXC5zPfncJU1cgrlClRyQTRYyaUV82/IB/tEtsd8q9Chqc9VDRf8NxsB
W0W8zvaQ/NljLg+Hs0Lk9B6sD1/bJgsP4Gg/7tCLyFB3oYmnbsc5azx4O9ra
8raTv48dkZkeLxZZkbzdWU1WVZRb71WfcT5tllXk2UcjSIQUNIVDzxE6m/v8
3zaDGKmW4CzKLkAtMutyrHlrfAYG4ef0hx7JLyMa7tqUZyHNE3e7S3qUFyUs
RS5zFoE+nwWtdTsexbC4unMTSaQcdpR+6Ckix4UZIje0C9kFmUBLJD9tPpYl
+MWmZSiU5M3sgkni+idVx6PhFBywAHkummVVcDsCYOHZXrqBuI8+jvDXgoBY
MgiEerSpcB6iWV0Ombfv8QVET2KhW9EDB328EHwIc9IuR0zhvrhzpg8ls7Uz
+VCCtf0Iu9rPeAcN1dk7CtYI+7ZqCyDQVgrqtnp9CzPI/UnesVuRQeMA5HsU
pXCA00n6uwkZe6VuHMDdvsSBp2i+SH+xHd0OfOHUxIt2cJ+Ah4I8OusZGJ5V
pwsyl2hxqUm6KCF5Ieps9IQOI6r1LYgwqtQNztaFKFh1bwq4Dqt1rk1xXFcO
jgsFhqnZkv+M4h02ZG8cHNSrNTh3vufUrBw/E5bYtRxsAtReJcr5kfPu1654
YJTcM2TfAh9NI80S3dYrD8ytwdtcHMmqVjDdgyww/ZpAVZgJD5/kEkBsVvsQ
UoUfaCuIpQ2N01jUwVsZ8CiMgGAlTRU3FbwQdstC9HLfDOAjVFmalqYOkgMp
fQouAPdwoyKrAwAazJTItcQ0F0EEw7PgS9LSQUlVS2PXZyNMPV24fAPUsnnf
LvGNAXtfkbb4DwQiDYAeoJ0sVPqHPFmp6uFU25VsntL5vgH6Jv31wYcn9Ga2
iVlfR8WON+hWMZozWZIv4jaMmAbByvQ/u3oCZCvr2+c+d9SrpyXRucZ6lsd/
eh8D3ydKUWUutyGKweBH/4yu8XYbg8vw7CFPJmJ34B0JfxA1GDcEgB4t8I5w
feBcpgug/12s/Pu+WIkcAsURDOGODeH1Xh47pkFDo9j1UvO3laSdSzouGnVx
kp8RuW3Le4ur94Ji1YD9IpS+kYCX4ZfI8WuibLpEoqSoiin0itPbZfDWVVpI
qIUpjFmzFBuhT5sFiYqAYPrKlqGUFuSh7a6gQhahQ317xR59MxGdRBEOwZsw
0xdMwftNciYurfhPn316n+o+olG7IR1KVACrBoj2hmKPYA+vusPnkYQKkp8C
wvEtWDX3k3LcKovp+0Lg3fJdhskjulFodt3dUgED0U+5G5fhKJfMcdL1NOxW
xAEaXQQdnsT5BeykEoqf8b+qn7c04quDhKX89FtHcrxDWI53QoHaiF8RNpsW
7uP25zo8/m1rXPBHr+LumDyOFvkgpqtpJwY8YByrm8QYTHOzwXmgwzVBcjzF
4uo2Hxarhftx6OrV4hJbzTwcN6JlUE3FRkQKKeuJ8jNffQ2bRFqFFAvb9UT+
ANrTqPjUM1iBPjT4pGyUTt/JQuF7biY+fcudL9FwYoNQEGcF0LmseKTL44rz
uutDBVucnsQ6asCtTWsfeKJ2HJ/Q0sQjFoB3Ikfs7LNa9d9qT3pzxotT3CWd
bztHKDs+UMSUte/dVzb+O2ag5dxx13XYpOrlaPVGf32KmplinDGBHPeUtgpP
Pk51MSMv5i5UKcD8FSqgCtwwo/6j8GjpXskCIrYtgkmW8AR6FYAscexHK9Qn
e8eWvezJ6DGWRedqt2wbTLEL4VMU6rpmhb2JuX0FgemwlumShLkQAVYl2X7v
szoc2MNcBC4DXAFEdy4M55HUOKMiiFISsdD3wbwtWmXxIafPs0bIF1/2xt94
+mvkGoH4/+NS9t+xHrXL/vyyymXMTeB5Z/A8cYhYiTS6mjHiuUucZHtvAkhx
wiPgbXq3kIo1cdeR1G0z3LITrw0t/xG/B/CSzMFXF1iz6YSxodm1T/y3k0k9
XlZlIUnIJv664Mk4LjcaUpfmOWLp1iESuEQZQ9MsEZZMQH2VKwjXhvz7umfS
/c98uNuuITbWsOxCPU3ZcSmyNIBY9M3AZAPgg40C/JyUoWOGCFT3B3aM27B8
8SKGml6mWRtyvVd7SKWNJGg9dvbZUJZ6YSGDlIwgey18wxndQqAgSYvtMh3k
RysddECPX4ad0hBC59wjaVlIDkFRN5ybF7IFJFQ/OBeFvKTnp5DPY3o3fja/
950nQaXqZlLoVs0Gl9+eEYYh1HyvNSotv0Fc3tfEOFj6qtKb8O2BAlFYKCUy
m59Ake7aNLZ31aCY5lAWpERV99nDOOaZTzK8aifzwR8NLg5EvSfBYZ+6DIRP
1tdAv9RiM/WE43VxLbQuhkUm0TCtVlRB4fxn1YDm8dlOeV9zU79kjZwP318z
0runCCTpC7Nje4/PBerxbGWC6Tcj7kJR5AkvWD1uw1jIGeHJLUXl4SMHv7g2
ubbHdkdIknAtNZqYlT1/lTNYxZOUYVfED+6JYgF5QRBUJNP9ZmSHAOhnqE11
u4OzdPbFkzzLDnnpcwVUBiSP8JuEv2BHDL/pmlivUyufoGEYkoXNOAfnzini
co3UyebMwG+VjPcQZdUXgiC/Nuz37Xsn4Pc1YeRCxd3dddU+FqS03EAmN3SY
xXgp4QIrTMRpSD/qcn3VXLAQXipS1LEWvq+wNXkGReuuSmiW2p3Swa0YE+4e
Ux1QxeFy08dwNwVXp+F4Bo0ZI36XIbuJyHn4pSF1CXIyF3+MRmO+EZiihT/z
vCTIxkIPIKb7Rc7k+isePSqVskna78ziPA9rcROezlwktSdkxuyi/GhUXKxQ
tu7sSOG5JMFk/v9h3nhgjP0Zi3pSsRhN8XgYZLNwCtzER1rABGaoCVmh2OL1
tmQW87H7nHfihxtdVMyHxpH8fOxe5i3BvpdM1lWA21ljZVllpojmXFzb3kPs
V4kSjM2JcVSjdhp7tHgbIYbzuupjZRVlvJUBiH2anjhKy8XUKE7pDRgTG7Sj
9BndNyISD7pZtPFFgMw1VW2i0w8Cx/evrF7Pkiy4Djx80ef5Ubux3ze3QmPZ
OE0/Lspt4mj9QfNBFiuBC/eND3qgIX6Y4rzZ/peQamxT82k7VdDQ+hd4XaUV
SqEXa4dUCF4kDKKqE6HY32HcOvKFgYIFPuXOnSXVljuiLahboBSop2Ci9wzN
udlHzDKgf/ZdLx4aVcmxzJvGyEnu1XZdOZOc7G3W8Gfw4mJTRenTb4rHKsGp
77xP+Hh4qOQwk/W9CH9X4SVcgNAG8/UvLdCiIuCrwHRICDkGqeECHJwEXNKr
X/srV5RP+FfVB96XYezNkjZdTE+yXwMUY9CCGO6gYScf2gsrQIh9FfTkMvWL
BrJUEbRS7HDkWKebPqQaGlO4mvcmL8eMyqlFXOTZFtXISq4x7IOZvExTBD2t
yV7pMunsfgU1ookLVpyz1ituCIHK7sz2AOax8ZRsmVOX6cdU7BekiRJSxBEq
4yquHllDQ5cVtFyMjxoBwCYk3TlsBZFkFz1dURfxSK2RLCO10n/KyQZMjzKQ
r0vLCIGNJsFyt/Uxng56AT0P/4pYF49EXdyvX5r8kEHF9yLgKJXT0x/QAHhX
ICR+RwZF8RG2sAe6R3hTb2q1oXJS5vyZio58xuc8AnDo0uHdBbkFG0ZmQRMz
t/Bm1vh3CbeLLZrLV6GYyhf5ajcJGjGI0W4R7M+9PFfxRYuouSeOQZcdF3CB
8E9PBtym3tMuk2FuCtXOZIezJCXrePWobAhXtcdUR+XWCOttTPGFE2nDp4jZ
1WDBJ1G0NaNQGdaZT87z1kJ0c9IrHlBJQqI3YxlOP4L4+RBeGRC8UhH/k8Uo
psM76yo7VeN56uvgrBX08LMl2uBxJgnEu1MkjxN0vWixxFkT7XD4s/2VZFkK
qeYavNfUNcQPBQCIckJqQQJbhTWUXvu7GZ2aHcC+Ud/DFN1fYSUrugz2m4g9
szmMHGR5ZAWDZxMqhUZGx7UBLIsanmhG8IYrJAwgzH8MSQXma7IEOsvkLaDj
qdv4/13eInbP5ySuEtdDW7BYDL63RzDMcZGpZIs1FGCCfMC6uIRg190W5U3K
O+3TElo+xYLPOKjZKo83DEpUIcMHU+IHy1QucKc9RDUub7Op2l7y6S7/ONp1
ymbzglqWVet2KeRaf2cdoHjKFCxKisqTMJhxzta3sw4duivKy7PX+oKTL5Lb
nYiIJp934cq1p9jqYKfTIZHgz9YqErAWdUI7dayUS0YjKxMCpMq5mqqiEL7Z
o8LXenPKc0niLrkhb9o0rZmik91Rgf/czsWT31SJTVfBN/Y7fzNcln3rdU6q
/PgSyHK5fAi8C7oS4crV8xLqknFol0jH7ang6NictZUL0wGb2hTPpGvuW2wx
TIVDS4BgNvQQaQuzSB+Rfv+lNg2BcqkiaakI5cIqgQoM8mPtP8qYCbLA/9KD
fD3Q+lnQZJfYl4mQOD/VVSMnKb9xKARxr7cXqCxXmgsssWhAHT5IHMZ3X/up
J82W6Gi/C9ozjmQV5GOshhyi5jEPRn3MZeWYeP+yCbkx6ADNajv7V/NJdvLv
996zOojb4D5Vj+zHOvOTS/dqmGru+WutZtfCMRxLhOZf72ItjNldpVX7hMFh
rDPzj5jOI5jaE6XTfgRU/MwYqs0pVVyEXf1MHKEWcCdsKzMLnjd9hXv5JdWT
NNUBWjq2XPr64QgdWa/pc4+BXmbKZXZfhiP1cpq0dBBWIIXDxnAoJp2QnvsQ
+4T2vk/ul6pIFdBAwoREnl/gaMv6LQ3xHVWJRt+le7sgovGZSQ4+NqqnLtQe
ooF7j2ZyVQNjO5d5gj5Xc777wql8qWqgQdlZVRZS8bDSgG22japbgRMawJLT
jEjQK/VQygJnbXvIVXq8pIr7ACXi3gbi+3b5opQgpBjhrG1WBhgWAV1p65t0
VY8pqAzRpKDedRQ8K/GlN50oVOSGsfBFbFfZcJ1/ZaGrVF77IyUh8fWF8l6M
KMWVDjpdw9lTRWe1Do/sOkQMS1BYUilpDcOvDaapNc7s/hy/So7GUDNaxuCx
ag3vnqEaZMTmdjHRFbIswp6v9zx8KUz58UQXrWPQNfpep7m5xsLBW6fnCTxa
5g+p5Yei3eZ99/tltAz6IH1m2LNq3T4HS6r2bYr2sMEu14ikSLrAPl3ZSiRf
tghX2Y8ivOmHseW0f9YYbJPCYgyJ6qh087ABvL5U+RxfqNYxQMVzQ9o0omBh
s+BP3wjhEIErTRFQ6i+TnX3p+Z6Xx4nj0NeO/nrAC0GxOwUfI1/u6tFbh1MR
igkt73bT6lZpkSURm84YydHweCKTPYeSrzg1hW89oKHP9N1afz4bGqs9snPE
Xf1TSPG3uFhiFF7062TJdd7nmKsmy+4FfF4a6oPNwfephde4Ct3EmR6Rr957
Z7i1ci3A9VSPPwvmH5UU6YM/br7uj11+aiUgILNTEO4B1ZEh+RfGD8VYWwMH
0OOI1APkTEY1BYmMtii0nME3pnTx2hrri2jHqfQE2LZdDILITXYtmLMKVe8v
JO0RYdqCdjQdGXpIg5lceWY7Gsb/cPcbiFSm58cWM1kjM0MzmyOlaHjaNvAZ
g9IUTjN8uzBWQY6FRE1Cu9GVGjDRPMXP/oh7in3Kid01aKjZJiJX/by6zU7m
9WqR01+DW8vbPBfTiFbwxuwqwxOEyGcJkPrFY3ufi/wHuoKlsDhDgjtLN7aW
5qVkGr5rTG2ZN7QDIaHSZutJrn78wv3VTb3/JJ2Nr5+u/7a/oTtlaONe/9/C
Fx855M/jrvUUef1UUfrFyZxSimovBVLdJSijOk7aA8y0R6zUrnopl8ZqROeG
eAYF9VLGJvxSQaINUnDqn7XoXyMY8Mg/5j3Mzv1MkyefWovxm6qXhXmW/hK8
eythCOCBcNrMfEoDyoJqBe2umUQ+/NcRUXzf6f032PsyNpsOA0q2cH4sVR6S
1SF0ToDF+64h5qhRUSn3Zcg3N7vbPDqgnUvWSKlo2VH6fSHCasaI80l1UIoT
wKE669fxNageJnyuieIFZy+U9QGvYRI5mOEH1P1AHWcCN4EDvXXRiTypnKbp
msNxWl8CkWdeyaV7tN8lQsYou5pzTb2Y7fhcJPNQ0Fn832U1NkVQESIBT2Nm
O5NjOKErArNIz2bGnHQPyt37SOcfoyEnQ75+A4TBZZUM1kodVg4MMPRMiqqv
pOjUjZBVHmH36gdGbiQPa6ozXXLZp/wlKB5PtrajIiuvo1G/ieXe85dj8+It
9x9WsxcDBfOb5zSx5ZGI08tp4iFPqJtGRct35gmn77pwjaGzLmHRWOJjmLml
euXLqwqKQOKt/VQe+S95qK5A5AKBz154PeReYWadxxz3UlYGi0gG9t9YcoXB
agef4ej7stUvHnyfHPyGMT3weOxGosI7l5mgxZ7Eab/7UB5nn3yLIaGjkzJo
TxL60ioWh3HmrAk8sfwqNOfS6XISjvjcQtrmJoYIjqJZbUpaaRVo+VcxNyxF
XeITxSVJ4CoXnxRExe4yP/HPIaFjrvRdwXVw8yMIYab2VmKavIBa9birVVpt
e4EeyAmix7X7MYyju7KgtO9OevLbvE015zwWj5zFWpOga3SiKH5EYBb5MqS+
Hx4SGPrMl1TEzSg4euVLl+fRGw8fbLdoIfVDNj9NIBflrU+xXn6/KuylbUMr
yLorrlEaYKl9PNZ6OKhMDXmPUd7eYwSrrJeGICKmsqH450EXAXiTVWJdpwjQ
ZKR0qBO1IHYyQ6boAV7vLme/M6EEuCLvEQ4qP9eCINQLExGzTlDGfANV1nlv
zFJMCTRS8QWFpCYX0yMaY3pCfTbvAWY0PJocCTHSmwwXTNUXp7r5Du1Q+qSp
tAW7K1ts674qXb4mnvsl8nKhzDWXdMXoqVtu3iY3HVyA5JAvvYguWU1ETTfb
GbhoWEPiRpaYMRY4tJgcACLl1FGQ+n+X5YgXS0hR2omBhIx5CMGlFlOHJdGi
95AHz4sd2easjljFmyqgbGhCNQDegjiSFEaOiK3p79K4ZRzaM3PItMr7nQh0
BvGV8a1YBq1Sudn7tH9GpxRKrGHuxZ0CGmZb5j/+IaaoFKyyq3480tzmfW2L
uUmjaNRWZl6e0zywwX6MMQavvleMEp+nlC1JOnsAn+p2HhQpN7r7IzdURZly
V14rzIwmGPPoEWUFvCNMharD4e8ulPuWolBXlr6tUhLpcadWnHwcWn9ulGGj
mfmsNHV6qTc7FE7eRADFtEziq37prjg5fW2WfJBSlfgzIOI/z4HNQHrCL6S9
7AuUoSLVZZ2xZ4UEqMR1U14X9OfC7y0eBR3h1yqHSsw3UONHBmWwQ0Samhao
4MM+gI6spPZTIJ6/vtg38BagzNUD5BpYpskBnQmTsLEzFt6lThzg44YQegI/
BuxjcfNwYLtQGyfZHNNtgK/wbM5acNot7hKW4SG1boTZqzmDsWIRfvJcBuAe
wu9TH/v57C+qQ911nwd6qlMvRhv71dXSk413Ov/eYhOnQKhhba/C6/FXZXJV
n2zZxevXDJlAxuGHSLMj6mmaHZ0fix9TDHy5+flvYKtuUDC8wp6WbPLw3v9u
VndpR9au6IvMDneC1tjk9LlDnLyElODLNF1qvuWfhvrWZGD1LlgyQMm1vLaC
i/BIRRkVtn+vTu+GoO6+8Nv+gp7DhisFiL8ViVcelcYKCxMcu1JYjhEpezBS
06IwjYsjjRUE5mRYEuRRd8CxtGRfVsvp5AHb2A44OQtMkhPb0KP2cLp2ejz1
GdRadAufBSHjdifmAQUHsLin6Dz2M64YnDnSw8R+c0XGDjF7kt65n+43iMDS
spka82mq3Kj47RxMC2r7+QYt1jNdLfFQohxJHPj84ew4JK7vtdgHnn942oq4
n8C27bmgZncqs3TnO5HHtx6DVd/vlvzj2FlsCFnyGxcn/7TdVTkyrNt5vv9Q
bai7WQKykCprmjl621TKy67aFE3awEm2XpuzPKwYezsDYvS//3hNzUW6uyU5
H7wUZBVUwq1PeV+49/pDFJJycwmMKWTrwn70cJG+MigVG3AvAaoI+vxwiqNy
ZPXu0phbTi2wVy6ahOoDYiJrZJT3VPQNO3i6/ilvUNRuD8nR6NM5qXUuzMF6
6g7o9t1efW/CZxreUHSW5RGK+m3oX34WLcqqq+yaYT07W3yIb8tlpnM0lOOQ
FrVNaXpFETfgG34oc49RT1AX9F0dmntS0rYYO0pwiyyX/is8pzQPrZ4SYkIb
k/VM/DGONduTdmW8mCAb3YKVQiPSBfmBLB5DIpBwi+5V6zgDK1nkHtqWMDpw
oF1tAixT3oNNrU92OS3Hb2xO0P1tM1pKc0kmwqJl8X0ekBQb8JeqzUvZ0Lp+
cDSfRk5SRY1ibzh1bkZ17UZi9wzdz59wFsmPvOu3rr5+9HRRev2w3ynPaeIB
mKIZ6C9wwFPpy5usdlk0rDjLF5jZKVetCaLQOlPv1ZvelbB/G0HxWs/VhKwe
CF+0VMKyDDvHD5oD6RLl0Svn6DvZqSGNboxtxXvIZ0Grhl29USDXph6NU+YW
/CDniPVyVkoxr3otYcxr9AWD+9C+wj7N1tXYvRrZ6O30FbRdy0AUUbJ4WjVW
4PwlY6/rrPPz1bbZWwRfQQ0VA1I1Wrl62FWufYxlrpIcgZS2uIs24+OuqoNS
iVSrdikJ+skDU682QH1PNdGZtVpOJvpq2oUj/VLMlyPKZjvAFOid1QRXf6iM
qKlF3ZPMqLye3RBybxTXqu8L7qr/FjcXjppnk0ROmUZi6PUzV8z7/c3/jWWl
tOksEtG3NhAD3+vIhnDr/yJX963V86D0wK07eaILi78nhgXo2iSdoRgga6qx
CHF1c4DF/HLN0KR67bdOE7PppeDXvWV7seWdaSTRa8GksRLHaQ4l5bpJO3bs
OF8zFnIg+K6P5BJgk1G/GzLDYFzqrUXD/5NWKf/EbMREtiBsrllJ3yt0w6R2
BcU6dunTBfl8i7exCYIfyZfvz7fwjZ6Mp4cFWdEdOR1NgY2h+3gOh46ou1ks
EtWn08Gb2Ds30SEDBX1rSGW32eJFJ6b+o+V/1lxRD6D/9GCvbht/chNm6DD6
8Q7KVAHuK4hLcTf39mY1+umeBG1iNKNx7PPSikLz3UdivNbdU1azNaPnVUAn
75eCklKwXPHh0lqGxuLvzZKlXiKcj5rN6X5P2gBuUoetNwiPsvwKFTN3sk3N
sHe18WMC/HkA/9++zrCyIdtRYSNCHhExR2wMB2yz2v75Fx0SG/jUWXeaC2IO
QOGzB4NZIxCh9wZ/JEGBGL/4SeI2S/GRgwIQdv4NSL1gCurthzbYM7TCHfI1
ZB58lfC2em1HgyWXPwhP3+rEoDs5+2yv5qYNbj388rL97HJpu+5VHLnTJfXI
TbClEG8V1SSXMRRIXL5fB6cNITwa5W7DT3XqVBdaGgKDITpvgTlcmoksf06w
BNBu48dgy4sqWycg9DgRzuNnqEe+Jiwv1FRnSr2MaqXuneEc4DfzcsP3ztZf
Wg3MlMwBap8VXubSGnN5rYYGSm81muR+w1Pq+xOjzr0gTPaJjVEru6HhrJD5
uP7GCA0BlmSmvtqnbaZ6EQrxlzTNLxGa9/qJQ6Z+uCYviCbzQgKFjI6m8YlY
G4lhWdihbI7otEveyUYGqLuFmZSC3/qp3cjGwABFaBvsAUiX0TRKjGvQ3Xtm
OF3WQJ5sOlyRnINexZJV6nUkxYWV6Qi+LtjQZEsUUtpwLMogVvk81RnGPIrj
GTmObYPbHGXtG2GxfvrvpjUmbr4ePInlS/T1ZQhNLEhbs0iMggY2NFMjE2Vg
OMpHta/2tWyYRccUBPBIwDYjKPBOwKBUTvPlhRXN0uDbhNelqcRK3ZZ44My4
xQBscoBpNUrzcz1F0V5ahxKBXhpPk0bY28jWaSx9UJqN2trjiL8BC2GSbjiT
iBs4V553YT2wEqq+sDvHcbFViY67Gq95ml21ZjV6kbs6tdidrxwrqWhDgffN
o8P84Y8aIrUcF+07fN5gTO9pwuukE+9JwNol8irPemPSDLc3TdQz2QAfbLSb
KfFGUzXhvdPu4LRtP5r0r5LZU/S95oMNq01mo9jCEFwLlWOI1wi6Kqeq37DB
3kDLDvMo3pLTf9G4jW3urIFmJ91lfuFBItEMh5j1QFDmZjtjeS+ZQJCiX1hz
smm3T4goScjZ6EnJbPw04MxVT0QkLyMgnxyDSHD1VCzZCevicLEeJuYFqX1S
gV0jANleLvB/Be+HsJCKOKBJ2pchH8WIKEZTyzcGiyDv77J30ESAXftV1BWd
ra+LRPV1am6sixJwBvMklnju2BgwDHkyT6V3/Qy+ftPgDEGGmigHlD9wDVRl
j9LNVRderCZZzbBrZjA8JFPc8twukh0jbVs00bWPlwHyqNklSrNcsCnxYPOq
kv3KCmMc0qKBirR9jLcTLjcMVhWrTT3y/x5rV5EAbmCbsIw8Z7h3UBJJv6pz
fZHknbbqHmDYKJyIIJFCqnaCPJnwjok9oT0+eBPUWp8XL9Mu/c9lUesZj8Z2
JJ+VYMRWaHhb3SkWJknbJQwYOw+FtJtIcVcjCYpZEL/GRMXoxEl82eXvGqmf
Zze8gBPYwzk+3zjIJj0HSTrOKpL9NnwUxUbY1ND7b5M+l8ufwICaf1oyB/9U
bvPljOoVfmdtyYK42uR/uz+nvmFMOzft2dnOdKdq9Glnyt0uXmw48h3tuhlQ
KvCZ5ojR6NovCpjoQDbONYvGeq8eHjFikuQyOfyUN5pomtGAQUwuhraHn75a
9ru6zLFKAWd2pMqklNnd+n9/S5704uaZw/E/Gbt+czV0o9XwLOt7W4oPHyIN
StgRX/czgACpCEAyOm8UrQCmcOHcj2ZvkhmM/YDpX2RaAsojDALAng/W+s6v
fjkraZGuoLrZgHGs2ewHPlY2X+/CsIRsRMM553Th6EuzTbJZmPLDktH9M7iL
WJWQqCrLP9v9IHG7j09DAFo1OyYHT2DI2e9Zj3HSovTUwf0aLF7TFPZn5+VJ
5lj+x04eqgEZxGQzf0zZ5sNF6O76kPuizVyujIJuOdw5xwh9WL/pYuz/Uy3h
OlWHef1V35hEthisxeAnjQ1oSPJh7m5SK8tgJv4kzXlWYSEsQLwMSDWJHz9b
XNlJlsKJguJDMoJ20I0lOxxZZNr1p690u9L0WB1dfv3zJZM774Qa1CgIukAn
8aOzq4hW51VDNHaW73JV72J9D3chBkzAygd5STk6pNsmJf+wELC6Kp15e9m2
88n+4rVkxd/mc3+MKZn97n37PpZlnI7wv8H4mT2zkYRDPc6hutY224HhzTJa
sCtC04rvpv4qQSdkSoYkiwVawZ1m8oF8AcUTkMe2F6zrkMnhhixBvDMN++A1
FJbHtXIXMJI2l1MBLVGYkP/BAgu49ytYDyMubYmI1rXDTffH6S/+PCj2Ogrx
A5jxBbSqHc++IR9sKtddgHIX5bIk8cuu+x3+L6oOGs5HBzWFSWM+E6NdkQTh
Tur7dw4RSu9tYxaifYlMuPj6gkl4pys+WnvYJG9YbipEDIFo62hCPV4uujwC
oOCPtLqjp+zJtv+rCslk/X7CRBwi5403dPF92tSb1/aJiHahEWiTN5BaWocS
nj02PFBj8qaM1DTZ7SaBkTpL6OGz+DZ4tmI1f1kBiOu8FiGml6lGdnIEBhu/
h2zncDPhGdF8YGtvcSGSJJVEyhIBii/Fe0aTmNBrqk59RnEcldK5HknFs8a2
ABHrTQkFFTdKsfE7h7lMOf3ZZVnRfpBEvydjPJrOZMw7y2qbPjhMOzs0DXFk
c5/NGki8cpkbFX/NcmR8u6XZ82wSgmJK4tBGx9MpzuQMdYbhlAPs7VuJfwp5
JoThE1th1nE0yCG17vmRcz+bdJY9CH/6mcfUjOyP52TrB+diEChjyWKzhTZ8
8lKtDEShrxu3SsFIx6dMsNMs5XIIRy4aplg8gcHjNQBNBCtV735aIGEKWzgT
6WFdylh6trRxkKVu6xCAL6dpwH8KZp2fyspiyvorQIA+egOXyWni9m5jYtDp
MeeYr4GHLH5YGPHzAuJxm+DipS4LnDRtHueLu7eodKhkw9Ko0DeRxhJNwCOZ
afmLfAbkm8ZzE1KH98tS7TJE4JB2f/+3pLG1nBrW1rpqnL7uYbDhUoTRrpki
aLioWoxM41E4yEQOlwL6Ru5QmlCfChrm/AKwlFIOXvbOj3wGBsAcWD4OJ3vn
OFCZ3BKHG3PHPrvvp7uwI1EfF2KxDQdJ45qr7RvoIn+mxDtpau+kLoPSyDNC
LfrsWMYaO07RYoQd4vO5Lt6ouxmm9627WwV7PTV2V58ZCpmu4gn5X8rXR8uV
QzepWU1tcJbocY4sZfjRnMzNYjOYqAOfmXmIt+Pq7ENdT3nbe5HLFD6+UImf
8YKxeZ7enPuSYHnOq/nSUGwAuRgosTrhmHkcfLbndp4G7SuXR2c+VhaMC41S
WCuy+2loc9P4bxRQAyDQQdfhae1ZAXMLgLb/0T4RfBGvC2EAX1MgY1x4+9mU
PQzQzvEHM6BUacY5jEiaSVpMuCqSTbftWKp+y9Q7RLe/0QzCygD08dkekJP8
Q6uOKUqroInL0RFUkroOc5rf3TEeWRyDdt2kkq7CrLWvaoAHQ24YomHAzgwb
xA+POUvMHwW0j+NLBKrEgrEOL07toHWi6IcC2XadMnGyVGnQ9IPfInRakZAD
dCg6nmzrSV7l+/N0TCB71IT2uGEkgp0VHjZbCWhHZA39jv4i2ZtWgBD5M2/g
WAfYYuOc0JddPDEob8GKn7Zbmh0y4zTLwgAXFgTY9ULhdUvHeCjUS9/ZWeXh
oqQePSnt2ccsVDhn+byjpE1bkpCyby6dsmVE4ytySrL6LKDpHoe7+GKicQie
1x2z9r4K9qYzkbLw271mRNeAg/R5jBdLdROXQFI+pU0Kp9mHP2HFF43oT+R7
AJ5CDovfJQZNC9lEjsQ8HImHW1+kTGmzQY9nalHABRdnnBN6BqW+9Svwmzpg
qowyT6uqNs1hmPujB5qHvAcw0zf3f3imoz3qctbFPUkp07AjTsuqVDHYp0cr
k+PVX/HRKYKWabX+Kmr8JlT/mdLHy6b8SgPVVjnCSZTL7cdP4bfGbCrcssI2
0poe2bmP/mcFAeB/Am3TLdPhYlx6KHCweCdQih2AdXgfQn5OJXWwj+1hc9vx
25cf+zHGn7mc6XSa0yo5/T8uYpwHvyIKZt0YOmE1SaXsmoNTbaap1GvjxdPn
37k7rPMtegQVZIHgUo+pg+JG4dtrGiwHGFgnknamOXNvEIJO1x5+hrzq4vX0
nrqc/s7lIkbkctogApYEWWhzV1zEkI0GRBoH/uQdhWq4PaYrl/KNFJK+4UOZ
dPPpsrAFfGN1wsKy01zIj97rbq6YCuOM403Cfl2EpipHNkhnGVQaz5j+pUGg
vEePKfhlOySeMhNUdsfg/R38xvLHyOwnDOyywxm7gm05lE6v4N1eAyUdarpO
Us647hd+tsmgyu2l72Qq4KXAFoIG7pYem0s7tNg6ugUn3b8u63TsZ039z/aC
ZiNdPDtoeAGtJs8Sl3NvW1woo1awspDYIlCGROMixPcH+21eILapUEAwWhHV
/l40ezM+HyxDqakoKeyCNg7xRVc79Tdu4OZogav8Xgmr0G3L3wmmuU5yIUMl
ud0StFbtnpLdO61Tw3cqq23isIabEXJ+jblHmJH63BkbXRsyw0yCSRVTAmlZ
KmS7qS6kysyDevYsE71T1mZFDF1BRKarnptixtSow+VO0BV/v+f7yDLmAtjl
FkVZsatgV3WCArkxINCn7tc8Icn7ukjT1zYyTpjvl9uj8+BQjujexgyw/dD+
TS1X+GWpQFWHybU5BpvGz9IxtDs855qf87W7rh6huqBaYXBVZv37aXKqqmP9
kOhpsptbd5H0905BNX7hiygHI+bZ4l0Q/FLMLzP+ab5CxwFEoP24U0BKECAe
vv31NCAPAsV5AlB6jBzRUoWLY0hRsMW+CqprGJiyjyz0dgvb7920u1GfGGH0
aNGnxlDBDIfFtumFzu6GjFQ2OSr3Mp0uXWK9tx29EH123hlcfCa5Rb7T5f8P
oZMqGh6/jxWnHEG4d3ZQs88HJzdtLQEsAcHtjR5W+c6KRcRvLQmaXpxJmbUG
k0yRVShUSqaMIL2uvW4u2+TekNJ4ebS/TT2ddoCPFxUX55m1c7f0U/E4HZkQ
SnrmwqBrAEFxOZPpPLG8PWceMArSsN+wSMwhD4cV47tOAau3DaVkLs1PpyB8
TFRao/1hdO60VeBXB70bb7U9+2eGX8wtHkBy0sAjxiH60uoc3Nd2DB3lQtV/
tgkvP83Zwu4DSdaoboBpi8wcCk3bZDtruTme5rQ3I2V0R6h9oyuNLrITmkug
mZwZtQvlUqhaPj9kS6SdFxpFYadD/CY/hAH/RI/+1psk8S1/bqlBl3lpcssL
agobO5rBzXQTJcGlYSXtIAcXt9KUuo86yqj+1WgSd/hanIPyVz5vgS+qnmOF
dI0yLpWiHeemZ6hDY5ZOhw7LuicErSmGJtHOCp8xkgkFNUbzrXvBEmNGfNMu
IK0vNMW9EWsf+PiBQA7n9L7KWafTmbctms3AwGSm0hHexcABrUvvoAa3bWIi
nLLZ3UnNvF2QiwK87Zs1npiW4amCxFlLLx4JsBQw6LXYVhG2OfNa92uF0V3S
N3T5ZYdgRk+Zw2gYRm9HBzMjWUulFF5Kk/FLvitR4AlXuwIfBpvlu+cXqG8p
V009zTxuWvFQ+qqL+82MtNTmtyLclxXKPRUl1riod44eqD0EVBaaUlgfWkJj
SGcBO2eT2iL/jAAFC/jWHTZukRuOkxn6rSrafQ+4SbFMMtoW5btaeNQKD0d3
7nAZAPjDVdm53XmC/IoVMabHjtYesstrYR16KgkbDDAmLzboBDLn5X/NwccJ
2RPNRonTp2fULwKeY2XX6ghm8+FHPzMZ71IfpN+IkLNe7BSSvy5+r77JYS5z
XpO3fDPlwujfuMvC/v/KBjPOzJ7Mpa6coRQKV+MGPwyeRPLK28lHaXiL+eIr
D+sMG8K8KD2S1pCtEDP+NZQ6aNsuCoRI006YwHadG4crnZQVXjh7/hioWMoK
YUA4yPIE3j97ZaqC1i1CcE55gQyuPeJSDjI03yZnc2ZsR0DIxpdP57WvplX/
uijLDG7Y3T/jO+z0hEqjFBptBFsX8eiwGaFQj+MVbaiQszrLjsrA6TdIyGgg
oeiWG+N5E3PqEyUma/xUsDi4xw2L7krvBEkgcSsWKKxDyYFefJEYkPcymBmV
w3FKYihIeAFe4aJTh3Nc16ng3fllKeGp99Mrx88XtKn/UDjsTCilBF4MB7xN
U1Lis4y7TQ+d+p6Vuiu2/cYVJEU655NuF1Jmy0+BxiWbwM9LoPlVPH+fMnn4
OsziBgVdcEkKqV0Stk8l//0veWBFs5Ly9fRuGQrhrXxSqOcAUCUoB9NUijN0
yrb6uYOS3ZMl2MlnjOien8JbRqDr/4Jnj+dIZP/JcHB5CaKpIh/3TWOeaq0G
Q1644jQuu0yvGvahjIOiXULEf1Dtn+CQtgInr3MDI9VHn/TPjIE9pG3NFMQo
u9k8sa7LKyHR+2OZvgHlW8B6xr4Oo8YJW4eVTYUfG8VrChWHFC66Xf80b8vG
TSakuL0Ji+bw/++V6tEyDUpV02OygCRAgZZmVt0bvMq96TEx1raGp/T/ObCj
s0iz/Ci0VAEqS5C7QHuYEZSkUN3I/D3gUgrDD/0/KttM69IERGACMylKuvXb
cIeXpc8qB6r4t7c+8ZfOYN8VLRiJvMKHRM4R7Kw0SjlgLlCPlIsLmRHqZzFy
5UfQaoh3pYKHin1mQryXWvdrfFsNcCzpSgZ8Z+4z7Lcwt/lBGkPUy39JMo/E
a6/pIwwdakP8nPB2zTJ0nhP3bia2akAk3AcM6wgQMzTH8Dbu8lTw2SvEg6Ho
sbhuV83ehq1RM+LzzoM2amnHYWUIHsUPtlzp3YH5mYI+4GE2VOSIVFBbWOvQ
VtwkVXoW1htM41ayPeV3LF7gdCTU6dmVYOZycFQ3XETFg2yZMQBktCiAXIGh
wABfCTgl1Sx9DVUDsRLGvVS1+96SkaEE2WqCt+P4/1hRbBklJ76hSmCfOypf
hxtnwlABwlsUz2x3ygvvi7fVi0MmaXjgPsnTeUKjanzgMmaC/GEVZ48HjSMe
QKxWHR7wBLrG3bi0hCwm9rVo3c4egORc94QmzBD3QfwR8mYtrvojPyjKT2+8
DRoDZRFO+PKpjHq0gvXxZe7JfEjyUoUjCu99gx+nSVW4d64JJO7H8krq5GfO
wlreIKFL7pZ4ZC/2koqJpQaAoBfXQM47AQqElrFZY1lqH0/EyYm6NVdGVORj
sAadJha28MDn8Arubo8p4VYn+IBduXTB11HxRghT/DCwtQ4FUnBD4ZqV77Px
eLOouSylVh+/kBjUEAL8B4tKxuLPgRpIrHnOoGmA4++Kwnnz8/osapznzsJL
UI3HW1WKdZmyZMakWlGdklKmpPZMSw4INNS6EZEdF+pBuZpeleVjdjZOP8SO
EXkCP8GMGWZhiPYl8hbFkiumCcqVqDbk9coN9q2ts5WyMu0FB6OlqXXEc0zn
thEwAcCNEEegG+Q17EP6GNHoUDBcoQu3vGW/K71vq25QWvstOKe7sDg2UTBt
RDZQI8I7Hdoy8EaDEs3C8vzGoBcZAzhBV+AiTs/zNyDpwzpsIRu3VUoBOuPL
Jk+KQhiqcX5mF4oG0/f1O4tdc6BTC1NAicRmh4pbqcN4D7oVQ6Hl7AMOdfjj
FHUldSyzWWcU0W3RgoENpAzBwOTtp/G/FZNBs7aXpglAnx0OfIFciq494XJR
VBlgB+9BzQfrpU2+nhGQp1+scsYtT70HTdEW0JQa2qLX4JL1rbUN0MQKL4Fb
U6nACQJ5dBJ4kNwdfjAEpVcHddVsucoj1GeAkoLZZcFzGBvOVHFbA4isLFlR
mhOn5J2SZmiwI3OwTDzFYgSOoxNq473SmIKSCVjUAXkAnhE3QxLvDMcO4pMI
J0DaB62W95942lf7gbFOzE1lhSk1D0PTXWY/XxqGgYDSFoeWLJsEcekNSZIV
Kem4R0BO/k28EuoaI2myB/XvEYzzUG73WUUUilspIHQmfPd/011N8/rDOyAP
GZdr5Mdx8lL1IamcimNO1VC448Q/5+ZVpYDl8k7NgUtn6S5WDZqzRa4iG7sc
j4dymu/oxDaz1yqKW3lfho1m6CMaPGNWx9jcvTjrdjKlq4W8+brubAcA4mqi
SDEsL0DiNhlG3zxydYb37sRElkEP9hCJPVB0DCFQLCi+jnO0StSEGboCoPdy
ko15yGaPSl9vrR66RdfObZgOyvLCmzH+9n5sqa1HhsH/BAbZbhrsG9o5+MT8
76FWfDURxRZ4rod+86zgZYBAzjEJGvgJ7NdQeMsT088WCrAUoZaKszrupe6b
JNKFAC9CJWSK501fKmSQ1ZCp+HwwM181ovv1iLy3MMQz/8tSSDHz/hYOO77a
ar0wCyibZxBDFIfJe/bQKqX2X4+l9aO90Ek2ZxBrC/E3unnL2iLeB/gaGs3B
jHR65ZS6wVXqjFIU28L3O2ePMEVqS/11F53jsmDdMMN+skTnm1G/wBUwH+2P
hvNdRAsKwU/dwzmpVTpXfib8msuYfImm/f4a1NZdSoE4pDzwOnDUM/zRcqPO
4sGTnc456Ww4n5ytX0/ie3ts0Xt8VBdjz3GE81liZSu6y/ooLn88Q8vMG+xw
94FR0GTK9EbUBRXV3hoLu3DH4Yr3lsZA+LpZXx3Si8kFz7PqkpGNEuiYKnIq
Qnb5inUsxKOUSMOumz0PNfGA4kBRMSPvN5CbPTFYOa3vSl5SAZOfhjCECTgB
jJ/Yl6M8m7wjDluQR2N+7WDa4wnCZwPbGifxd9ziP3c723sjXdg6vOBziN/d
m94iLb+ODzXgODl0Jiu/YWNM1Za+/9DMLKO7eymxA60RfHJB7D+ETcZJC0aR
ei1LICXnF2r6TwvxzCzcAXMYMCD6SnN+maKLc3MxI0VNCaHzsonFrj5ghJhf
31jI45/9+ijKbmQvwpPlzIXRLq10iSwv5fqsZ3R87QeokbhgGM1C5dRE7fHZ
eQNXghpfEZ73tsXLNdO4RgNlfaXD7nqm39sXvkJYK8WpzCPIiJU0XMuc7Juc
9fjVe9yefe1UOHmK8fNh1cIeXI4IJUzlgAGpis850jqxNIZ0fSFJVq5SlF/5
8F1XyJF16fxZCT6gQT9/XFzRKe6KrN06nZEoxii78qA7QYfVYODYHJDyabAI
4f7W3DOe6JzgV+h8gmNZSHEP1ZufolAzpn8I/apjTjlix6kld3N/XBXDm9Sj
SiGZ8cud9rCQv17k3E3hEeGkU+sPRcTzWvJMT7EJYAmGS0jufJTBSJoFSxI/
ghaDYX1bcx0ub2fAQBPxvcCmaQdpo2/2fuzvHl2bP4oEFnXuJ5yuD+CVmwpR
u9WmNTBVWnKBzYCr0QZpVsZq21rJxdrOQ+mILIguEbkckV7VQtmQJjg9LYcj
npf3/7iAHmYegMLEAvX1h7g1lDydNwsTdH+UQG/KLkpm4I8x8CmSY1hYenau
10XU82yaithj0qiJfGy530qHC0Ixh04UI7BZiokQHvCPsgnktLTd6HAT66JP
qmZXiYFv4v4gwo13MNmCT0tHsBUCSONSJZrijX7VhpklZASEq6hbR5ZRtP5e
uJb1NZPbq8W1VYhNl6Pwic+H4k8EfwVBH1Z7RvjtkAxKj/etvFu8cM1E/Q3g
gdr5OX+iE3bZzQ5OH3sh2QBo3MrUBOOf3l0Vsr+CY30dLiECg1A6ubJhwsxb
mQT8uO/mZ9lgSHsqiK5zSjEZVlDPawT8G15UxM7oEtaUzlslnFlJLyg4EK8k
FyY8E+S5OPscBj4JQjbxdeCcNbZOkh/qJyubxnjzoybDbVMywCaMt5MNO1eH
TkHvfpxLaWEofWbd9bGYUvO/tWKUs07jnckassPuZ4rWl5nquvNSR0LsPsc9
XN0SHXUiRjGwIV2aMhbRKk8uzDpnZgHZgHfLTl1CQwYA24A+RhpL5vuKSAxu
QpB5OHGfRnbRuC1gOHfKE5xtXbsUpewGehCl0/WU72eQLjLbI4YJxpfQn3rf
lhukVv+uzEKAifzOaF+DEofmi4k8o6TjOGK3V6vPp0+IE7FjNW61bu2Wp2fa
ICT2nhI0mU42KlJBxdd9c1m8dC1fziQsAxBQnPumWj0i54+sXxL5zppj0ONG
NiIrNtf3pl6fHbRnhqnV8FwJDlkywipJmVnYbw6eGjcp3zwnJunL/3erTY4B
HKBodZUcjCjwIq5DYgEhB2tDB6q3dRESfFvwPEmgFL2aphCkRH5eY/o9Fplp
O6MuwqOLBFmK2tPEsQwVTIbx52dLX2eYyO15pj1XsrLM7O9m7o55Bs5kcrNl
Fva7hgOiTGpAvxPWHZJzVw1K3UJaZCwL0LeJK35if9rp5D2VnV8/PbB17G7w
/cEKeHlpYN/O7AtmbmbSS3xDu+j/sFv9/+SrK3rOoAbRcmDzgL3rsn8jn3S3
n0jJXcSb6dXgQ//tGjJClQqnyIgmNdaSmFNpirsZLb0Bgob50sjthlMTVzt1
6rd/gDx1xK5IxdI8A38RnumEZO+zBOQ2/Rr/EX9TmQo8rHCSGA1UW9YyKyiB
GLCFmT4D4vjK2JsZwZsT2LXPMh4ffIG2bDx7tuHVdtUaTxqZGYe1ElrvJIIs
HcSwr55JNN/NVyFT4Zn7drQfhnqUmgZo/DP8rdx5iZ0PcfZ4D3AcxvhxG57p
WwX8jWm3ah+OTvMuZMVsXd7G1ISUM+i65Ts2QUvHz0eCbPMoFdPqYAyKlXms
hnXG1er7um0PAZdKp1AegCQdaYfeL6F5mr9zyRcYl0HrFZEjKObqEF3zDOLo
0ND0R/pKhbdsQ8IFACW7zy0S4luEjduRIs+Lv3MftXNAjevcj1gRIXWLvTO9
ZcAJkiTxKxopoifGe5vljslBFm1CskSpBpHkGXeux8SYEm9E+BSKWk0mOAeg
1CH9lEOvKZj3BozW8e32MTOS5OpqTa6CcgkPUFbpJTWIvwKZTyYkkSZXgtdS
GmZ8JWwq4gNMBdnNHYxqH//NcoGVBUUEgOeEb3M33oN8d2/Vk08CjaK+mO7f
SHfcemNjY3IQGz6seg0iL4ZuZXazlUToyGQ5nG1mzVyuYFQ3Pi9WOpgtLB0B
sXIsgnT1SY4ObOmdS4X2vi74rpvpSKOVK7w+NWj3rDCQFxuaTK9ocYTsiV29
hZzRXoIfIRcQFKdA/10ggrT6NHWOlN/QWY1kEqWXMFKx2kDlLDEVIirEGSBa
7p/5fIHEKAe+SVpTeG/JpD2ilKgwdMIpURW/OlrtX2I7HxXFQFDfOX3NJ7jj
l9ZQI9V2hX6C9REqoTKeC3XSpn928WCPUp/w3GrAjcLl/h1aC7LOSGW8HZaO
UvA5MWyslq4jjZynDqu7ygW/DVRHdk4yyULCxiULTt3vvm0crtLtZEr9E/3p
1ARhvjhxbWYbFoWxg0HRIyyjsK7MdhVjV6MBqMWwA1TBo+7ZLrXgUwL99xVu
5uoPtCXR8n3mR5/hLqFfD3YQ6zJJ+wprNB/oe2NM2EjkDleUMnHPM02ZefjO
ya9xp+l+ZemCdpaTwcg1rRVm/adY7RXPGxT3bzzV+0kyanWtwg9EA0inDe5d
GZUHEYBWkx0vbTHMRN2XwmPz4HjT06colgWkpYGi6et/nJg7Pry15fUwQB6m
LfJuqUyFlDfN5pHhHPIDWNsY7od4UI0F4gfs+CXewsNaSSQjYjN5NGz8Zh0j
YEqoRVf46+W3ZtGieHL3uiviAhtPLsfQZ/SMQT38c1plkU0rkSZG51KKL6/+
6ytEW3kTCnMPz7ASexLLZ7SnHs0bG/KhplKjduylRqZC3/+zXHrXcxqQX9pj
BtuKQ58UtU6v7DUjzF1kNPFwbshJzAKUMRlWjrF0Qv6y2qnUEQKYLTHONUbn
9rYEdBzW2WCMuwpShaDUhT8QuH5aERvfagB5nmrQ04YcZjNP3kiEvfbkrgL6
Rk56GUaM1+BtbtiTVDYo5n+ZQ3lTFxLXUt0GThJ2adzHfs5wXp6T7Rdqd+D+
/UovMof5YvqEGlETmiNbzPN36NQ9KVvR1r3AXHdOcPo3YK9LzmXpBVfNDySl
FNjvidw+4Bwn11iki/46LxUN3+LrjbZbZ/IajWTDSl9e44SDvWke3xXgIRvw
xXKlEPml91Jy37tNZ/o5EzBo9Umt602lhe1CePlzukaYluBEnZYGXANxd4+U
qOPerzKjFTjV3PcYYw4fzQhTmrvMA+tpebZnFeD6mFGNxIcvVnAL4hxct27B
DVzftfayFvK22qn+9l2JZ4KqSn0E+lJyovB33Wnjyuz9q/dcCS9whliB32pu
ASc8nsv+6hGa+MJ9B0oD0hojmkArwJ0/HnP7y73j/TM3PCYsFtBBfGsQfWy6
HCxpVKdfiFbXQ6wMiQcxIT5342xq3ZaGbPXhpaa758FNxe0+YqTsLKrgSEfj
+Zm1lViIxyz/fAqh09g7jOw7XbM0uAR1uPUz9v3EjcHn0siXSdo4O0IF0lcY
tTY9os43P7tYCa0kV2bHWhoail1CEd5N3DPVECrTzT55TyzfJhP3V27H/BAO
J6ldOENCffr/Lv7VHK838AxaDd1DOh15L791vhMjvdIwRm+tr16j83VY61CJ
8dLZCq9woC/m1fHViu/SOf47HZSkeI089qw4rIIW1OONMeZyD5Rqo/ORsFHI
+jmEpruedxnvzExTi4TEV8VXYbys97K9Yy9Bdr4pu3ZXmrtFlxr3COVMwQuy
BONzclTu0kVzH8FrQ9oAqc6oQTHlsnClR6gShSWNtJAXRSVLt2+z3IN12TZ8
hQAta9YjxFzK8SL9mu3rC5t8B14rBRy/KHM/Lm7d65lKpI+YhVquf4Q5d8P1
FvRnL2CL5+yydjBW8S3b1kJZyzvvZsUg+8mMGIOKWf/J3SJogYVeAmDiDbFC
/rFoMjl+ZUuw0aG8tNJ1w3I6pDnUs70I2Y4b/3cFefj+SbSRldFhtNAqb61f
l3CXd8FYvG+1Lum6j7+vO7Bz+I2HK2xFzx8FJmc29IoaqBucGYZ+qCVY5Lv2
oZQOnuuISX9wWV3ff/tzVYEZA/F6TrFe5pMrdgg7Cktao/v5NxfeCLxFANZ0
g90O65K/ZpfhVxQNJZz20EXxYVrja/xyHO1fNiFiY4zoyKy5fDsg2VYIW7OO
DRt1bKMg9n6DNk04Wz49ON9v8PBdM3iFS37uYsTnBndR8F+yNnMuGSWHFp2N
nGmsjL70GI5tcYINWhKM35+gaWMO4wv78nC6CAZYVtlcougYx91cPoCnj/QG
sv4/kvLd57RGtIEpd9KvZ6YcCnTzZHqBVGAzRAXvPWZVZ1DUp4Kd5o3TPvpM
uinuIF7KA8yxM5JSxDrRaJXxunWRNeyBY0ispv4e2hYQasD57hfbfZ7SBJHC
waUEnY7wG8TU5IXWwD3Bwa90fX4YZdvPjgysEvrEoialXExvD9qyQmpe+8Jr
iYzyJTwiuQ8jCHQPYSe33/robZSQZMusiXFqFzX1NVFX/lqYQGoBHh6NCEzT
WYs5jbWuv6cttdJn6bDcTNjNmRJ8wiFANvn7Awkas8Ax3fp4BuJsaqRC3k8t
05MJzy9khnkYsSshJhJ0dWcKMvjHvDwUzAHFR7RTc01uauGf4boVX2ypwo1d
91h8mBrorsKceaUMtuwisDVNKckMuA+EKJDL+wDWz8UR/mfvdht4OHu123C9
Xp523V0xm8udmk2+JF6obmqfYjzQAil/akVUbNBEbNTlVCYnEaPygB7OhL8R
vGg2AK3HIyRHYAS/805RlBGrM5fQhg3hnlvwaDgc4iGr1AB89wteDDOsdIVd
o8sRD9lVVMY+UrO4vEAkHjPyhFq2NTerFtcB+qBcs0mSK2UMHXoFXLF41yEa
Su6+71vDjLD+yCALQU3dkTIPQcxNT2IA0TfARj41nr4gJnW8jlHCehe1vL79
EYS+1w32J4Hjt8wTZmGGO/mF6t46OI0lv2POr/l+IMl3AaiVJwpMjVxS3HbE
oqLcWiV4rkWZ/GbRviWcloyWXQsAhRssXFzEPvB2hg5GCXnqDnPk2r2zkSQP
0arVtSM1PHl3KB/Ex9sD1OCkA6+uqCFvcZ4l5c1llHzSi2BUjex125U1QQyM
plIGGHRWANC1x3lpafRcRf1ijCz6PdqGdmvj9qKHX67DWvBN4HvMUPDZE+WG
ZE0Y5cKA05SsI5mnJlR+33/sDlgV03e5+Ym5tCwqq1APuGvoYk73qn5vGc9a
CXCE7NvolXb+vo4vQUS0nIx/WdRgk4TUpGcZ5iT5pnoDJiRM5Et+v79apYx9
8liP+fNtMCZukgbdmbbDkG0/qanSxDELQnlNzredcnBQNi5rU4uzxQOUHf3h
uoQdxkczYRbF6jlpqbl0gQC/QII4x5gwj4CspfN9lANuP+0uLdqiSAKP5PdZ
oFWa5W1IelidAnJr27vScAGRKZH7DDSQukkLcQs/p3qB4nxvBXUM/Hso36ZQ
Lw1cR3QG3tLIa8D3i7lo780KUDSoUepP4FW/9wPP9J5wXL3VsYY548yI74z/
t+raYqjYRSjzbY7AB9ER/I1+Yfb1q5xLiuPo4TncY1G4DJNBFOduYFvhiZ/D
xKhjMGxqJOcX6SH+rk2VrB+WDvf+kzGOfLYBSw/stCtzSRBTP2xi1DCUbuB5
X+/7rj9RkOAuqMNOIybcCUWt2hqEJUHr3/m1V/hh8j5YTFeYJ0lPrgKB4mlv
0PgXMpPmu++WfZXiJ06iOb9bJs3Iv5/+iZt6sWJSZ+Z3ZiKGC0zsQtq185dW
6Znj+UM1ZI8R3P6TXFlRziCHfAHlgThWfDyZHjTNZ1bF0xvStP0BefExxtvW
NmitARqUcbTFIMyc8vpy09J4JshxeBWCTDebAeIw7XQIF37SjYX4wCGvqSyH
C6QCD6DeSyyLMi+PZoJ6xq3lqUdNuPmQAoqbdn05p2d8KdpId+nK64RkkW91
y6fiV1ZL8+Hh6LdLio/Fg9hzePGiahuM41diu6bfXG6YzAHb3mdUf/Mn3nGZ
jPMmA5Hd+McTym0TGC75l7nH8Am5O0WJFW8V2PySvFonH6xaVchsCh7KsYVt
pig0rva5Jq8hcnWXUsYvcvNJYqnsznLn+MY+79xI8ou/4RkrNf3BmG9u6kW+
DdVvZk8+ai97z8yT+LXl5jCKzdO56rr1/v4+/nT0K9uvqOWJKfiu0Giml8tk
YKgyV/xPkl54lTFLBvU3do07BNYEuDpwUhu0YBdNhkJOY+1AdL2hWP8tTT9e
qQSHvzzz56S0mTawXJftBMl0ARCfmbDuaHD8CPCVo78Jyx/HtC0zvac0sr58
W+U0NktivBwheXaLHv9XRUZ/TT0s+AFwwhR7b7f+YdQ8EOvqtK5IoPg+bL0R
nWn6fwpzV1GgXjd+3DZ0qyaoDwaXpcRDEy2qQhQ2gyMVpRRFbm1pMF4BJHib
ULw4iEK2Un9ifx9GsAsNAv8M2XTS4ZhD6u0TtWhxzyM+IutTmFLUkUZXrBVK
yXuoEH0W6eR3b5ww0fnCeeQ5dQ5kXJoiJAm6sEz4a/r3Ns6AuDqq/cHfHnDM
Anmw/lSc11PK3c9HIkojvjbDb5QLMSyRkHkrmlGj6RIFIJBXfJntYZLOJepS
kBPy2xCZOp9BYtX2vG06FOLvRQAYCR6Z3PgWn4wqC95wsv8y64meYQ5QO0Vr
Z4tQ3ffF2lwsZnwL91bPvxMDUZRKbcOO7eRW6STOqA9joy2eNJELhuRzdhnQ
+lQG7oS1/07X7XK4HW1iUfwaIHiAmrUD68oFJaar9rBW+DAKr1Fc/26P37RR
io/pqgUnxkLlddLjMeUV4NwryBzB9YnC7FxnTw4vUVzb8Llpgkj8VJRBHhiV
+HwSUw8Fk8AvzHmlpIpP9GClgHdSPMGPal/3d1T4wsrGnsBOj8MTPYzKqdbg
wmM9JmAQIe6hO28yUIALXQIqrBzBnfnYAHzeSsaC6yhVlPJmun7liu5Iy+n4
2JrQCfIa58mQoB46gq6fbLyAOkGX3y1gMZCbCrYvQDFzCVZb5HaS3Pu/wXHK
IdbUhPDBd14L8pPLBD7CThrP4bgaBaLLTWJmo6f6tTZKfINSe4CQdR36eZO2
Eyz6MgTJult6wnl4Exp7Q9KYODoFx4PP3vmqd0tg9rfIUFGtBrKxuUdXn5s5
m5tHzMl9Rjt8tCTCjRX2WwieQbxD0LQ0z73tvA+dch4sBM4zPStmWO7qIisz
p4D+ybNgyCHDoz4ht+aK6wyRAvoBvMYuQXw/arqmgX0LR8v8vdpaYP/qMMYk
OgQtrCC1ZYXTaqmnp1hDTClPfrQ3IUykODIdY4nzwlMI1SghBPtVsYMhUBK5
G/vH7qslRXjR5pw6/Py4szTuOeBahBWrPxv+wdqFjVWRtgKBK3wPxx/eDPMR
yK9BqtKwygxkOVjiw8ribJogjjMaZdy+qEwOL2uzrO6XqN0n9cBK9TxC9tMr
N4YQG5zoDiVKv1ACS8CvLmy122XXbDhnT2imJOgfbV7RQnbIy2o+YUb1JYSH
DRfezC7uUxgpoh7Jwon/OFjjXS0a60vUXNQbwH9mJAbCGvZEbSH8uLGGSsU6
zMBZ7JXNGxD4UjDkEggz/20X6y6ariiVruk2TE1a/kozWRHLaxrqX95PaSJ2
6v6/r5Vnan1bfsY5+KfzYBet6ga8MxDnXRavwh/Dcl9bk6V1n+1h43eEOiaV
rG6GvviHFtkZe3G0TFF4kncNB5rxI3VGb4XfyrZCWLyzk5aOfGufqOp+Zgrq
KTf2uA1QXetkpwkDNtsW5YP+aKDiPcEgMetCxLukDgm7HaoHiBst9STEOfCM
VTBiDBD+fHW5FH+6RWjzr9JYAhIPlYGSvnjGBvbdYbwzuQv3cy5Mgv6P2BUr
tBqDsos/DdfAUeMSbAZ8cB13jmX9V4MT+r8xq8/eZLO1P0yq9U94f3oz56b/
oFS4zxpQt4i7hoZ1K8XHXeN7giGQTW2mAkQ9Qv3AIxyp3dq+7k+eMfd3eSiU
7vbHEBpl+aQ4f90/JFW7C6GY1lfPH26T8W2F5erj9R0fXi7VMa5JyZvts+q+
HATQWH1S54A2KW2QVawsxgnIcTstK2j6vULzVCp6t5JcbwnnICLHXyGgmXIY
eTpy06L07Y7JbgIhby/Ojwk+XdDPVrZ/6SBn9Jf52mvvvuxMYCqHYhh+54oZ
Uz3YHnqPGeiiulPsitVaV1tid7XAyFQNm8OiJSLHzJwIK1QFgqu+zk6rgR6t
gIx3JzirpayEzwoWB4yJRde9L2WIJYs7LILvQ0Mc5qWPgdlLZM2ZyOZeDNVW
GrU6+/TqJ808uJobePUk2+D7cM8HbeGvYndt2yFF4KXYUzSDYLZNxBlSZYf0
luFSC6Oy6s0FB7vBY5BX5bL/EPNFV/tPm/XZe9R7jGQC0LxXFf/zLVTsh3n6
LSZXKPqkiLyeozbIk0Hie6SGocAITX1Dq4qW2aKsgaWYXtRByet/aNNyIQUw
iDMB9Yz6C+I3BYJobF0oEOpeczkyANd70oOsG8H0sMyYqVQWx7GTqBhNHmOy
qdfVcdnKnSgDW4ihBiPAlYoSW2NaidtgxXDwtDX4COAOUCPb1ujwufc7SG0S
O4bjZlOBRgGE379XfL45svug3UcjV1uiAsgtvg5NDy/GBb+QkhI+OXMY7P1y
P2uedVTyfXVtdabzlauuCI6T8mzx8YWP2vk9fhw70K9eZjCs1GqPhoPbnIXz
qcvxNS2jH77GRCRM9QfO1FSR3AFlaQuQryblen5EXqVxQwp2sobcqPciQ1HT
r5qOcvKsiEaggmMYhLRDNCZJ8LGkfcykY0+yuTTPjEmdCOGtRvIe+Hp0jkMj
0GZXpPauaiReH+uGycXw5fc8ugbj109ufdH5FdfuIrgXmN6iL8FHKqXL2xYp
HHtr0ZgRDVJcec+6WQSp0VYb5I7TGDYgBt6tweO7ugJWSvd4xAKWM1DJmSns
+3/h+oLBt4lPFsl+/vJARMi8dFOuNpZ3V9poG+dNkQ2/pVqk+i46EEH5WPq7
gv3w8FSOoMRXdjLoJhMtT8yTUwPJvIC8qBhMGysTsEF4u0JeJmJUraf8D3nF
avSvx0ze8dY2Ttpj7g4RG6NlVZKC1jtqr4GYr7JQr5W5K6IxNoRpNgCemMbX
uQh/ud/HVnFROvTdFxGqB2BcqtzS0ZwQb4ayRobbOxn8Qrhw4WRB77U9YyXC
HjcWQQTK11env9AebcN2nFALhAjsGcGSVSqbBkspAqSoNvHdCFDQ7CNdEVeT
FHjGobaMf6scBg+CR7OC3b3LsJFHr9B1hRJi6+WbwWWbyHkvF2b6bJx9r3eK
tb4vXi1kFj/we7xebAwhj5607g+4pvojPwnVU2E+xTVBbRTaXWLo+R1pmyys
miiheE42EhpFmpLI3ic9d1Oq5EmX5H4tmqUabS644pQuvfZAZuE8jurI/i9g
5h0fPVeudnNl5DnUImAg1RHXSOaQu2EPzsSiuhKBnY5bubEeMzluqFrFd9cx
YrwEEh92M63k1FI0q/blX9A4w2205vUsp0H7fry/wcMEoJYEsgvnFF68BQnK
LK6V7h26ck6vY2Ik7ZWmVMFDIjr9GBMNGwbRm5R3RoqMd36b34ZTXL0CWp7r
i5AiqTBKRu7kuFJBCdU8neXLv+ksAghP4Og8U7bezAHUmvjQdIxhBG3djo4a
VzrBHQ9owD1i6Y6Wszja2ZPCPCpsqORO23fSLWqiBJYJMq+EseGABF0AUWR+
lQb2+2SCtQoM00yheKHPfAIXmKiY6LCXNF+5aeqho5xw8ajG1llBZ8oS28Ej
/GdM2hBueqd5FvDfRyeyNwKJt2/9Usc1oL0I7mJnKud25vjUCMID/W04KSfL
EFkFNGP0XaRpkS8mvt0IVWMSqfocXUF8BCwOCnOTJRTBokjR086VSRB6nuUD
kXJAeLXPgokRETdGM7VyPsR5kJhkS8PDiuamxOZJvRL9uSiDKyNtoDY5ByZs
sZEwC41w1xyGJKYcpOTkwfa+X5AYlgYzHtvfNODjuUzDfqr5c7oG2+WL58Ei
WUfIjQ1QdJWPzqbh78JTa7Brchk48jJCmABguswq0haRXOeMlKUFu865qGGu
vKvVGut50s2uAHEb8fEiyWI9t7EGg6N9Hu74IXNggq1Z/I9xjES+DbEbcbrz
DmGYtpuYNB4T0VhEUB8/46X99lJcSuH7Us6sWt5sBNwWtAahIewedK2mb1eU
P6a8JrSXsW1y71NV1N2kH8gWYpWpp2ayUshJjn0hJEVwml079kj7iIenFvIc
pgOqR3n7dfpTGEO9nX0u5TzqcY8lt44Hkvk9BHy8P61EkI8WmaSnMBZGuKYA
RtT7dXiP90ubHNNWHvR7b4EBt/LWVJtDi9Y1IPeG5LCQZb+ZayR35NcXu/dP
6SEsf22SfejUCZcqEDUt8Extr9Tyg9jhDbEyelnGwutos+K/LO3N9CDlEnZf
lJF2vMuTNmJJsMfu9BLYmFvD9ApegstRHEWMZMXGhYnpcCrzZqzc5ew1Xda5
ypXlaxHE6vQ6CTPa/xt/aw0g5Oxe6xdaPQY2Eh8zdzvTcs4fM9GGtdNAI3dr
fLybuxG2vlmK8lApmyPkL1v4+yd5P1PJIQ6cfiQOPIrVse74KGBDJKmwhUNv
4Oe29fjEeV2TiLkU1zXnFHEWEX2SwiHBqLu5MUQtwoT4l55757VNlOAqS28D
yxDTceg+74ULbD2u67aj4rApxlQ74f33iawmzMHfIqWYkr9tmufVNL7LBgSA
QR5+TEmqSi1fG4ymHaKu8XWB9Tg/WEsyYPcazZIKznF2e6qLjR9LfIKpU0WX
pw8WyuCa+ZsayQ730VbaAtS5baFwMnGSDbIpvvu4+GAM8YMGnKI3vV76JeZb
x/MeQCEMxOXOSJYNdLdcU2GJRotfSOJ67jGXwbUgtvmbHSgCRYTvMQld8RDU
eOftJneT0WHGri7gChqfNd65goF/91enOCnB6wPP1JtfpJ2+obY5v99cNfB/
2G8YpVp8wx4EflVKsUBiLgLrHUn/NePuFPHema0F4V0G2+CpTrGSVbtgoxKT
qD4VeIhq6FPMk+b/dKORXjEoPJSbLf2KL2ni1t2Mt5X9Cl7EauYEMntY2cH9
O5niBAVPpO20XVCC+g7SVQ4JTgpu/WFRhg8X7am7PFi/LO5pihHzzieeOZeT
y1LDZyT6VSdDYksFjkh/uEDFeK4uQWUnj+BEbDe1nuj8OTLAQtw7GhJ0gDqD
KN1mVgKuc2t1z0GWPFUe30zpXBeYKHYbTEoZCkwq+l9exDIl8KSA+wSCYWV2
nupTkGJ9sz1+qG8FfHB2lhDtOubzO5zvo/Hk3USdoZgiHINlvrg8sj+ATOn5
d50sJhCg2qPjIXQ1MCNieRvKN9C9hzew0fAnyugParQuuWSthzp1Pje/dOgq
12CIPQIzq+GhyFtWbiSuIACgud9urQ6UB5nXjCtElLvZgvg+1mYx34xTPgFm
Xc/MpGxoWg7S1bsfxgkHBueVgS8Bmvi5H59QagP8PtTmU/Jo8VM4+AM57hL3
li5dqwEi9v0NGEfDhq8nqQNEWMpUP+80EKqXw6C0bPxc+vD1PF6zfPiv5jbK
qpX4EpurCy6+ehTFLClUQq0C14xpgh20IH/bJhItWMeh+aw7SPwc4RbjZK8B
RFKBP4Cnd2DQOLYNh5lLUqGpzS702Xx7lJwqFNv1777gMeuzDXLrPMLITX1M
9Vx143PMNIfBpY0ebRQHq6WLn6Fk3BT5ZwWYM+Joe+OXfuI9LZ/O3n5VVH2F
Or+L7vPaL1obLuWWEbHBFajwlW5lB/EBodYYwxYdnhx/rnG9Y0MhvLmREWMG
Uv2Q3dyIlkXkbz2ha6bnCAoNmNbh0QUrnb43jATFMlJOFTxRrLhRa05dITlF
FuZHzgYlR+dEvi/on6xgw02LBYDjNMolydcnd9xCo8KmE9OAeSqzfq23gifp
nhvHi81/MTeoWp93efzkJaGzagyvh9n4FjKedCTD+KVIK+mCYhddcdZ92Q6M
5px8VYLlFSuYroefr+OHMWQewP0iN39BFfw0cYo72qgBmiAzzCT8W07jEweS
POXGgp/3dIoHoF4KIPK8mdAhnPo9DilX5om2fPo3CEF8vv0Ak5svWJP0n7hj
A6LMnvpQLDFStrIaNYubE6JHPXZ+pVGZpk1MZC9M/IQ4oTpXQP4E1mwcSvNT
oItLUZR2T/O/gQKquNvTObNvmwCVb00XQ3uUSJ3qtu+vrVTzuNLJ2pmpBdpH
jq5CisqLqKtZw3GsysSLDZdwZkRrigXTjHhAb1D5gytn8uyAzTi+FiEi8fF9
AFet+PxisM1QSFSAbOPfhd2Ewn5SIGx6hSNUVES4BNJdJpj4A9xV8oOKnbWp
BbAGgQHpYrcbodFc+aCjvzklIu3udiOyYIK9PN62+hFl9N/WflWcCXHTppRa
HZ8NCuYFCZytI5BRpSH5Wwdzeo98zMPXxgY8+qzLF+QjhaKYCvDNYAD4Nkmh
fssNNRizgUeZfAtMjK+SNvoovGbPN8pxvQ7eZPC6RoNvtiPqXWcQc+Ox9r81
KjIxStmUJ3+lSRr8eV+efN5ZanPr6DccMINy7Wljc7yD2nfY3wwTbnRgKBzf
BV0fsWZwQcW89UQ/QUJ40TXGwmXtPorwdCmWGLRy2N0sxx7VbmD6K45G9/lG
3l/IBMFR0rzJkt5MLsLdbzf4YD7kOxS5kibC1m6sKVtufWQnkRIKjqJ1yKvq
NgpdxExZljnXmZyUjufifdWYeNfTLAhEdGugDc/s72G+vb8bQlXq5nPjZnbS
7xobnvttV2m2/6pIEsKWyf6emE2EyT5Jg93nwgM0eEKLzVgnb6zhJui1eMM7
QC/ouOBazLVMB4baTqVy9D2rbAiOz0ezORwezCtrUCQWGSlbCLEA7mevuEEG
QxqIUVOW8qjygKGqLAly5j1txRnY5bJhoqx5suT44epcv1H3fGNC4JCUnXtI
NhpC7GDmdwNmiJnmEAY+O1Be+FV4CimEnCu+4Xo5nfylz6io8M2uk9AF0SMW
OBj4ksguWL/eiZUKTQtBXjAsvJXJh/KuO+ikmAWIwPcZPt2/woi7pQg4a2QC
AyujjbOPxlg1PXlxOXpI1LoXWtf30w9XMgwFoX4GZlkpb6FcIxXL1NGxc/GA
tGFp0ouXz6SHlZx/bxdG8A2rrUmBYtWayp+aGXuhXY110C3UIGg3JbL96vKf
Krl/ZHtnJ6CGoy3eRY1NvA6lVIXyiSwn1KJkQ3kau5gfFAUwE603izo9gulk
0NMC7GF/NpZR5fnXusqNOifQbO18z2/10oHO8jKPW34poVayLsa4UVKbRfOc
v7GcwyaUoBBdNJusImlz49UsxVxrev3aoPDKiJwiUMWxDly6Ny3Ukobb6FJ0
nfu28JNK5CA9flwTjpdOHXC/9QYnEzWqygK72otsdGYsOw3D/xuNHGjfyJFG
eRRVglIz+mFWQAIWQomCaASyKxFhDj07TfdO7FxPHp2+T9t7R0Ve0U22DwT+
ELtsA116lonYkEEIl6J5ltES7YinZVYcaQYyugI4aXiI2uss4fvYQoyRRPT4
6SSoy3AOmTxc2UG8S7cOXEJ/4zFmkGnQYf50oQDDA75zcG3kBMNLlPE5Q+hv
MNAy0/9/BL7vJLLaG3DZPyhGj8ljCZHTHGylhLmJsY2zmYeBXhCQcoapoUuK
Sk7w6hUmFzer7UPcHV6V17y3Y7dKXwLpgp3wKcQMkedjGyDQoTbQifw4+Z2j
mjRYsctJOvXmTlS6x6ktJmUGItrq8ysCDfZFCvkP9SMF9nnyI9nZNXTbVSGn
2iP0hpOVOvxjdYBIHWhjF1ODWdmxPfIdoBIed16QtO1hrpgxx/mmUOQcOWbE
KbWp03DATI5MfW1US91F4/+jjY2+UW7yRh5WzpzCgbIZ4a1Uh9ORm0/0EBny
JYt+smWbGy7CJCAut3ajFRACD4TXj/WqBXUHYuYgHaG1lRQOnSTYDUqGEqYS
iPsnb0Jb394rbhFer2NMfVvaN/HUSazOYva9Xt6v8JGP5SL7d+lO1eryAWgs
fcsU0kr4Jgem/P98Fn640zH0C9xSrTi5EXSbS2nsrwEZI/8hDHo3+iup45w9
NLPd6XNjOzGQdicruyD8976xRTMbmzT4that5xCC1U7kJ8fbyRNXsKRWIpUB
fErnLqHEVHqAY2yEnbgtnXAy8Icifr3NA368z55OHuewjHoT/cVmub6I7x14
+15nx1jxztyQifs4it4B85emN+8KXOiF3IwtMZ6AH4lcmEhHcRJL+bCtWW6H
dWafiyDV/TPrwkd+9PV8S+HpC1xC8Oyo1bQPqr4WFrg0gV12u+z/Y8LqBeOt
g47/Fb/mddU7S1PTiqWApHFok/SF3Bze7nBx7BaFTSxHLv5ABs/OoOvvVDtu
aeNfo4fAH1G/C6efOHvaolkexycd2mi40mr/A7b4Vnnvftm2oJd15rDDg/wx
yv9sDlX9gNnVBTuH43PYASF5uZor6OjVNfk9IAt+vGOukZl+CiafzPUMyL4Z
zXQm4MOiLOgarvLu4alGO/6eHl7i+vd82eQoa7OR/JRkFaNimh3G7zJBKUBK
UeFB0mR6K2CP3vHvPoZgaX8vbzYwm+pODm3ApPU1EeD+/bqtM0ljUQ1TMcIu
K1FL0tFzombfhV5qHYIj1j4JYaK2ndOsARx1/u+kpmMU3bXdK6Kggv97KVr5
l+7NCihTaBU+bP+0SM011cStgnROMGDgLBdeq5ywITstyk48AOA1fY+tr9Ow
HiiN1VAPJoOPqD6T4EzCchkAcywuC/QsIfLbL1wFCMZVM8tbe14apqaMOCOu
bEolfYt0lb33qj2hKKA7OLBf+3qm+bdWQCsC6akMncDulKx9UtXt9yjmP/IW
4CkplSrrqXi6aoKmi48QZyAzDM3JgkP2FezLm//Ck7QsqDLMaiGpvY33I38A
FG7KsF/O9zSaqBMkIyEDqDUgjAKh0yfJkIzxPFi3VRQfNxv515t/vZ623xgc
sfDgijJQIPq2cYyVXkGYadN+YvFbkn8QFUZZKq7LpegY2isQbrW3iam45lz+
/KNqeldJM8aDnFjpOSZ31HP+mf5/D+F/Zw6PKDnYC3ppviwtd762LhDf8I04
pB2CQsz24Z99B46HE5lHPzbJ9bTVwvL8RAW3jXJ/QAGViRQhOJ67/d91xGHS
G7d7TOfG9NyzarAqGgIvvWLQ4m/S5+2TjXX8fmQLupdRT9ZQE64+2R6ExD9E
SlquXVO6+k8NKjRsbno/v5kytVTQh+5HfEhjh8vVoAUXnd54sCHtf9D92v1q
3mUgWawe8I6YoAziUHsl4BaHBjRVVwpxEJDIJu+C5sr25xUGaksh+IasK6JQ
sUK973NRMAgjZoSbqnKIi9IIdURTxAvmnBxxoJeGSw6Ipxz9kY+kI4QDxbKh
svAJ/vQaxlZu0296UrucVCz/ZX1T5zVdNWS+Wt0RXVkT1XfJNTJwUQxpncQZ
0HuPIknGyhCsDEZfgETNgiuk2EkvPC1p2hxgz+gTN7CkuTClPmHSBk5le3XD
v19r4jDxp20aCBzNWb4zWSaamD9MKUzS/3cqRBITk1857QtLJQQQCRqC1Qxo
9U9UUm4yq22i7kyX5kOv8gdyNjOYOCp4n6H10eJr2Ymrm+oXeAO/gWH12Yek
ASY9SVTnBrEPnjhocWl94xXgsgj+W0Mz/L0fxMBAxK1onJ8vTA2d+erX9xLW
tyPMmGL0Lk8COR/DlifAe8ZoWrt79guLQfKILITNiIdGCZTPOasV04kyT85t
H9c6B5awDWwGQlUV1MgMoFiD01J71TisZArxLeiX+ychjdcFnVQf3CHPHNtE
wTdrbuerWwqVSh/1Tixb8lrJBX4FucZNTB92wj5xKZrdgL/kJsDJbGhjy/IK
PRPjFAMZzCOiJd6rTliUAAcNjmwV/nQyDje7c/DtORL4hmYiYTJw7qN7aZwt
onfCOuFwzA9myemBD1jsY6EjxGCCAwwHlHe6XAb8mzkS1ubqQahGzraBFEew
SNpuMHuerTj1ZO4pghEQffdaGRw9zB9TndVMLZNR04PhNMtyXTVUAI8yhH6B
1GoehVQP7cOOUNKVXwuM8Sps75dOBRxyAL6AuH/o2oePerWyXtPaK/Uejmtd
c48FgoFF4grcQKxkCG0Xa/epJYr/jI3Q6LDUQ0G0k1AWmj3cX3OASG3t52B5
6vIEeYiLg5gi+bHhQCLil+U6YFDxESduEApDM3ZB9Eb1P4IEHie9sAPDuw3h
CGcofPxZnV33BeLSZoZ9D9lLp8GMLUpxAjKuIeq2amx8wV18YYhO4/p/2KeA
pVRcZ6LsuROzFOxktlyPkEovPo/Hqr+jzKima6k3EeBZKT5ZFdqkxwctbolB
3Wqtwyik+qPw/wBT3GEaLlZlYg9+NKlntMAW9XtsBJKJqCQlQZCDus43IRMy
I79A0UJhd2TzRYPJ6S9ybXT05LJbjhPYE0np/EPl7AkGFGogucaL81AW34Gl
MDby9+Bye+bxMWmj57namr5gmgaP6IiE7Lrfneq/UlNFMQEjaM/8GgVPTsrS
hhTCWj6YHR9M96Jfzw5o528QqKyBlvAWaGwmT0SZ8wWfPOtUtb7pVAMB1TRg
VZZyKxSlCgNlqO5jOpVogSX/wTY6a5O7K853NhSDAyHAg1bP8Lg5QndrMGeb
N16gUtSEUM/AY7H67upvC4rJ+J6ZbFsTEj16eEBNyHaesQP6++HL7SO7PYKr
bbl9ZaWK8fXSXK5SbpO28d5P9wQvviLlap5s0d0QoGDydk2oBEh9HuC8k7hg
esYs/nEQuQSRzrnm1Dud0yNHsyi7H0cQT8pzN/+CTmTuutxCOn2L2jk48bdA
Ws7xKR+TAlENwjJDcll/CYL5ev7f3IZiKYpR2TcbtuZAW6eTRfdQtSg4PGxW
zcv3DEwEMzb0S1bzD+T+HC4kYhpTMjk+PjfGXApnhKN7lPC+Hn+o2exlIPgy
Rm0ngfkZARs4FGCdenLLp4L44f/UhdrroCWkEnqC23bUezZCuKfhoLeE6/vH
gWE/x10w+oByPKwll4xKTexN6ZRAAPt63cCTU0uQ7ImsyVuZfB8nmV0cqj3s
5Nm/CU9z8VYObAdGHiilTgHi5HDRls5ky/gmzFUTZ8zESg+xW8KJXXMfVZ0P
UGdffKCVuDFTLjjzU2Lpl8BUg9OKvEnhvR3htYId0XJyIlIe1PE7axtnR4Zl
zTSxRa2Lo57TANgsxLxPzhhagsXbz3ECa8lYfobhzFCSOCbUYJW7yIHSz5be
bJYLkpF8ip6rdBimPsuSvl+YEb8jMdGmBh/obbdEjvo255Xp8vpeb9UgeEhx
LnzbBxWTWOUr+CmDNLKCPfxQqP9vNHqL/PFU8anrBbL0Vnl5VG9EUlQZcXLp
xu/kmQZCBFAedk8gKtHDC/ofqg4A8aXtofFRSxegktYPD02DsnnMxwaHlY0Q
1B62uzAM2f29apMMK4ESwn0x4sCWn7CQWPcHsiVX8YMvmbwl3n1iT5KRf7NF
T06+S74pYq0kb3HK5LZuO3SX7uxhKWn/6iMmYv+EXLayJmz1GToWj2PifVrC
wG/BaVe441XdEivxuiI3Kto5i60wYh1HS5A4XzAFV2oythuUuZNLhnhKGHm6
hNI/uIBnzbsJKiF8TrnLIym+ToWeYPRAV7qDxwxovpi3y82WYwzsRIwpvTCT
sb0mYoL07CIYSFtyTkPDxmY7zjtAEFwqHeZqMd9QK8r6qaKI9LqLXWrnhBP5
FvoxUfrMHlfhu5E529fUYhdQUslnZRBNzA4Xu3i9W0HbTGxUxyutn+Cs+iMW
vYH7i2MO1rPe3qSHD58lQgVomqeGgHoxWKe2DvhSR2cWim9ODspkPCerYpOY
8S58yPTnQbJsAkLCt3GEgkeTm7xKusw4MwKJcy4sfualxEcA150yn6TiuE30
7hghiuznuaaEyK1lsIjhJYAOtPmpjg9tvkn523+rYlqOFCT3xrnpyKa/XOip
64M668w5NsW3i7P7ZL9djmV0SBoNWPELG47noyvlFU5pAi9rtrDtIIFvkZYv
d57N4RJeV8DbuuOGpoKcWdYCrEyI/tJYQH2MNkaMTbXIaG4oQuyHB9fZs4+X
Gf75o12pMUcLymKniZrDKS5WAGiug11yAB9ZtM//S70lxR95k4gtM4odRG3v
xkEr9qVm3hIGksTjAvi32SrywZPfHHTiWyP1dOunVK/PIyGTBrha9QSP2ale
+9rQ5pTWYgeUuygeChLFDG1huTXImlMxLmyeUsctUS6w8fIpsCQ/sUcB3ajR
wu+nFlXSr3ojqIEpCPdYaqvtHPddVjCzxcyKqCBcDaTTFgL2hmwuOhMlz0x9
5d2DelA/H2dJF7Hi5+esp1yZJ/lHTyFnFO6NSPbzvJgKePRg121xOOK2Yooy
p5JAye6k8cVRiaENcihT3nO7i16dC0vGaJq7VsKmKwJ8UpmLu60if2dg3rpO
W0AZ1w6QGPPWVR72Usd7++ZeMbOQgK93xvmK05CTA/4IZlCx45EeFnGDBvJF
PIaB9nvnyTrAyl5ZUDHQCHkHsU8oN5l8gsEqR6z/Ggrr/s/7JcnFbRXqyYPa
ZY7gOZuML5eQT6h41kQqZyxJqQFtsnAdqkcsdJPyXKZTG3OjmP5wflF2UP/u
2qhd/QRO80VOm0SDo66sRxNCjQNzh5AtWXqJ9+xEgkD35aRsgHKrrPpJ4ltd
KoQqsBn2Rf27XCXVNC2UwdBCnNnEGIIyXqTxHaEEaNszsPVfNNl0oll1SR3a
Jhb3vDwF9rWPd+dPL2a5wgTrgRNCv1d9FCuGO0iUzcWdaklz+38zm6RrCJ1p
5bA3DKYFJSmcepQm/V2bmGjM8vjNEAnSOr89rVL+Caus3CY2/mnhH6wiUl8W
JuEY/ahhZV5JSiE6C9YTjKlCUbX06MtWRw+NWwCfkvZoN/IeToKL99dPnhTP
yXtCAkyWH361AwfMZNq12A8H71ndBlhqbn6v7tWRZfTvMncc7JTEn6WEWcid
A/cpmK3/ZhaqzENU7uHoByPZaebJoMgmAodNyUvLm3A3zhbajjRy64cduU+4
NMRGTVl1dCjVASROJfbaSCcL6tPlRKPIiep7wfXLYLscX16f9g1hePOM9iws
sTkFQ2aFCzjplvWY0lPILW6OsjK8GBSdpZwb73i8MvhwFWFovTDqMHNLUwIv
w5JOF51mrA66n70wvEnLR8bmYJbP+UnrW+R5C7a7Um81pub/tOsutq8U3F/m
lFUYhFnK6/zdUUbbjCtha+pLOk0a2yx0equpSsWrHJV9aJje5cZ9/xWuK/kw
gv1aAxZl5AR2mDJf9DWfqwGjgyeMa73V6gynThA6MXsRN010Rlh1YHzcvVT5
Nx6FFUg6I9CJmxzphHT6fIk56R9UFEProHKAPq+rIUJ3uHJiDUri9AwipY/9
syA6kzzwnvlpVtRDPQQiDfGFksLUMngLYMnQnb+UpHbgGNR5Ejw+BQY3KFJN
4+V3LxOoO/ABC3litpC2Hd/4UfHmom5jqOEX5AhWaDJHsaNwMnfqJ3BMkzHJ
HRZ9ii3xMra51++1fWuMj7qre5xKw3ysE+NO/m55Lh/AKcUwF1cd5ou09BRW
IaZLGeyxUf5BImb8giabB2H2Ks66cPf5UbZmU/KG0jCAzeYQVCYmXAwOuSiP
2x4pbMpX8xt0WmX0jxE4a0LABtrOla9XWIR5QinsfvX5uLLztENbBYRT18jJ
za5kvZgowBCNsG2uHgs9kz4eUvpfSo8PhK/x0yE0uUY0iAWGBwN65qx3o7L7
pv1OGgd0aa1NdFCJr54i9saQnQiVsnEMbe1xRmPc46ndK/EBHydc/bo6Xk7w
OAvJlqH7UlTEvY24kDZQCkNXtOxVDFg8oGbjwSsPtUNLVxmpMKh6aCucktxA
1a/a+CjdntlHNbOkvU+ogxoR1R+41NuYm4PGwCZ1gVdfv5tdkQOQYF38e0Gq
+BFn/iKv3RL4y4qvrjj82fkvAsleA9WrFQ4T3QcLheW3J8BLcm5XB0fGUSbx
OoBc3soMbkZAkhsdEww325vYo0CngiyybZ7S63MLK/R5FvwGimk6STirbZDl
joyBeu75GsX/s5bJksDtC16BO7VUZCxMzRPjrtDWelcFeGT6Kmwh/L5GRHwR
osj3dsk5xU39Xzz0oTslqLrBzwABlRH0WpT0AXWdb/MV122sWjY0aQVBiQlL
9PhDSdxUXVw57EWHp9wIPHUUGdqclTmefaus444cdG3actiVdjBLTqVVm58l
FR4s49i11dZLhnOQXxAPRvnbV2dCZhVW9aaEee6IvjX1TgMfln1SsycOkKTQ
l+LgAnHiiKS0kMwO0x2R9Kc+jtQil7UzRBFWTmTGK/prqKSLDWDO/W++t5MP
6qIJ2miPkeFEAmevdU6zrCggC/HBWV6huzo5UD9Addb6bbvbOkPxuVbOv889
kkYV2a9tXg5TrWBqxnFW9vwA/YTT6CE0ftdXaXhh+Ij4uJPKH/O7ypyNtPJy
PUF7X4BbcxKvy/pbfgZ1MxgIDA4xv6WBXZWL7UvwSIx3govhXi9+wLPJMe6Y
SFvFnPwyLNUkeClzfkpeN3eMSMAf4ZCkuabshcTtpDTXbKpJVUXgru0FJsKP
ZuQb6iQ1mY+/y1WEuxCBTUFcDmVSQv9e8ARGR6dCZzsq/0TF4d7nHUTzcabq
KR5i+XD9ULbXtzlNVPn5ZHzRj96PNqz8egwVfLD2v5ci+4aZOtK5bfIVRPdv
stvni0z+26X0G2CRvwxFVLZXbWILHAJypQO3hFizQMmNTyq/t3M6VRiifB7I
+w0zZNJjl2Py/VDgksLKHep5CEj/+0PBWEzyKVj1BpluhEcKgM0KTXR5Nf2+
fysssVwJ2LajFt0GhJCuMLk3PWrix3+U8UdOXurZe+qvK/f6TZhiIjvKm2ZO
e1EfQNISSUiowu0uQ4LHEx3HtojALHz3PGcROTTxVq5InR02nDJgMhsiBIWZ
rX9pCCNsnuvWzQX8/r5SGQlIIso4tuDrc53ksN8XzfdHOzh8VVsYQqOyC2s/
ID432GOgRmAmadwf2E7oDEkKP/K6j89l0qQ+v+IBr0rVI0kJWWiFNnkKAQkQ
aoQ6zFZO7c/da+KwWlu3JZxvmmz5NV2mlcJlL6+f0cVrxmf9lLBa/H6fFsFG
PKn/02AECgViA4SU+6ob/rJ8ayQyv4yS01pFaVGnn2gZSjSuVEeODwQoMjBi
MUH793aVoJ8qYUr2h8GafmDrFBcaqrJejjJB8u0oTKvGN1L32kBOlLb+PU1e
TaKZfsRQKjYNz9osHaWRSOeRhhxNtHGJhx/lbnLDo9Z+328nAMYV9E5sIyYa
kMh9B8tu4tyBvYPvtf0XHW2Tbgr3E/uYQsIEOpuiA6CFA1EYuYfB+N6tqema
UEvqxKzvxbZJ+mwCvbkxzNlGOzviWMnaJg6yWnuITBefW8EK1kOYUMSK1MWy
eAu1RdW679wxwnShJfYiM0aMwf3b+ciq3ZJtTVtm3EMZ7czVKmzP7Ap69zNk
FiJbj6kNDtj4ywaZKet7XrGkb0KMypB4cX8KFZ4z9Re2WFxqX9BdD7rQAVac
b11xzKe5oH7yJCvoEuXoAfzJfiteVSN3YU0fWjMnvqQrEul8C6FgxjhvVaiZ
18k5vss/22ZMLe3ikSj1Wki1AOwfMbkIYmkl4RRzBwcGeuvncd+c43jZBGSK
bVsrczsAnkVGjdO86pAgoTIQcVysyNy9wA4MxS1Zy/KmWD6XtXccsITVUo2Z
IEBi3I/w0DEGnwIcOTNftVXVw6VCxxXojox0BOnAjyaDsUSIJyKYQu/lVZnw
4l4cSufnPteuIxUKfFyctsVteNDBQdHfgfUa4KTK8NCDWiRRqEiu0yZq0mZd
KTqiNKe5jyqMzNMYH6aA58TBHzv1QTlXw683ujSefYqLcL0AkG3LCPwU9au9
8LgfZqV/0LiRwM+EJgmIj71XpDotIhaNOdWo8OuPFad+e8LIZ5/oVxafgd3m
t+leCzCyADquzroEb4Qock6I/VX6+XscUxBgMNaVsXNDi6Ko1ZKd37Zx/gVu
Lnn2fl8XsQP5KKN5dUItXQIiZb45W5MD1F4dqk3Cqrk9kvD4pyob2Jd7Rshz
sxtRYW+9sdtkXonypWXeGd9P02UbXvXKSAN23A5QfwPCcElffRX7inptDzFF
UqiTMiqcVzBcfHiN5TBQYHYBBhZeICNe+pswvyqR9Bu4tC900PPdHBJ0AvUI
RWfNwXYcyaP/USWt64sIp4PBlMosf1NZMvJsCgwRr1BdpgGPYwRtAYf/pU4q
TeQKhwft7fP3BM1VsojSzKMaZZYYXsyP+N6F4y+/2aIbqrKH/hZUtnToGlks
/H62HgjQMwIiMywF6Tb1Tjo1o0iM4hd3l1htW0FLfp5B/L1zeY0a30D+jOaj
FbT7xBuB9EAPUcLk8+0dcucA5oGAIcEYrmT5X1ddnXTbW7kT6AY/0JJTRBF7
ct6+sIiezz5wpMqv8CCmfvKSkMLCii0JzpnEBuzm7K6yiKPYL8Avqt4xfZEk
kk5/9bFAWVS1YhnSz0AGWH2mB3GC362sMpuu6XUBSolEIlr6bl0v1+DIyc6Q
+m8DhaLdkaQPlRwoF0WCLVWzgxuE562mpx0yOyIV+SD66B60c0QUUAFF5ZGH
RC1yt6VHo06Q4HDuei9QGVW+srYWPldeNQvW4o1yxy9+Wu0ZBPY5i+QXZUjJ
QCyt/9CfNls0qqSL3uJkidlFTDR0unZ3F0sDmozY/6TxSvw3adQLm0iEOyxn
NLCnx3nODxyHBgn+T5lkZDrUN3Aprp1xVh5nAZalIwuz4h2Gww9vxXblucHe
ptWHcKzqOhZg2R9kXPZPgNw50Ri6zHq9yX3csxuEEzjIhCjnnGU+Xl3/hSei
iA3aBe94qsmhcfEDXpRAWaJh1NI+/YHp+/AaVOH3at84NYg6uzmj0eyvJOgY
Gpu4494xRrPDfx6TO6RP5HCQG26VSMzTXqYV1gD1qFJk+CQgSpFcA2ny25ah
L5BC88mV2S3F9YbbmzXLZ2VCqL/OHh9OK6dDbw2eoeZL5+3CHTu1I2r/hf8u
rb79rjJEyTvSPxr3inuAxihM8ef7cgqstraSDfCtUp24bznW7uweFlV8alok
eCnaSpEzOEy1eArZ4VCR8YMbym18v6iixwvLRy8k0QLqISaPRpV24WbXUsNT
tAWhjkZVj3asm0jK9RZFKu2oA5bZ5iwwI6oJYRQQvyjYkwcCZLpnrgYTarw+
zBhpA42Mrk99/hmL4qNB5Bofy+3oZVfJ5tNrnpPESaJHYiQTGgOsWf4AmTXH
Y4htYDH8NTgz5lKS37jBEmPPWi/7uXt6KtoBmkuEffsiIqvZ4dlqX5tFkWbi
Nmb1pWMo7wTyIAGZJEQ9y4x241PMWxqEpsOosLgTBKJ4lWp0/wnoHI1gBNvI
cDQilb6IPly26BE94aaVm0L27LscUm6cpiWAoT4b2SUvL8WACnuN4rC2hvFs
x9dxmvO7gzUkU6KeObZ30A7evhsd4uF+gvDAS94Hb+cSThXaNmScVntTkUsp
e+lQMIxBpX3xvrckIlBE9f4rbp1AoxviTwuPf3XwT6u7+k9FfKAeVHUUx4pV
BzVFUFu4pmni6qn3XeSYvcL+Ct/0XRgwK15i6q1EA/ZP+2n4Y0CvtzdVJJdd
r+yYCYtUCZfu3cw5VV8698rVLiIOe3r49JnfzPLmFhmnEKajDk6231gNCI4z
q/gpdpnoTTYlOj3JfP7W6NUcjtvefiOPC1DBhLbXv1lREm+HTkmeX8zdG6CM
BGW9ya9V+HcNuKWxhmgTrOBMlRolqVvCH9a5wHJDKlWqiXURAxGQMQ/6QD30
oZ60yi1KrUxam/Gvan6gIm+4+6YDOftSnUw3T9nYqdH1P+y1rfg2cTBoPUsI
oureZXN99QPmiq/k7BZoGImdQEontSySQ9sIRm7CJlnybBlAqtLLbDD3ozpf
KitsNGjYGuvFzt50UkHjYUip/PFLabAKjLESBxw7Nb+hSjO0SbPttovG75WE
3BI9PfFB3SadJDJN5ZXbzufpk5NT373eY/t5wVdWjU1leOEziDemsYBbcXKC
5jw5EUKaX1RjawJp2wdNLmH/mW58Nhgq18TxspzK0G1POsDES22ECV9PC8rn
fUxguTtts3Yau9R4s6lqq+8eQh45n89M2pHruHE25QIxu90Mqf1P6s0VZxPq
F8hRp+9STIoJFhtLPR4n12b4/s3dV8fk0Kt7DQ0ZiAmxrvEwVrcrPe3bh3S5
W5E5iZbXcrOJUHC7hkYuesOjiuqSzvMG9aIuGg6xXv7Gbdd+MQDDG/GhJ+fh
p1SGlz8nPKkE6vlgwYfMO11irvBjrNqFLSIexyzEYxcLCEBFjtXyl01H2Yyf
Yu8XkILp2x7AS3CaVsyhB1RQ7Oya9zivzvD2nRffmGKz1YSxgHM81oDaCj4B
uPxMHQpOok1WfXsO1lPYOasD4C9PXU4sB6OV0m5VcJSwQWxTe0bWdXXLB/FV
Ec2Ql8GzHZ+uFBwwo5MgA7NMr8NZdQiIA1ALvzl/UKFjOCkHc2cgxZbfWeDJ
uK/am6L7tO6GZ5arlPemMKUie1flgz9tkYrGNrvUIOYRe+XiOEvRksgsPRQi
97LePEmJX7V3vN901lGvxD7SPEuDvplpjfz+WfZ+oqUZjULAbdHxiwbR0XH8
7iSywICOrr5XRgLQKvRKQ3RKVLLgg+VVxvdPKzmpdDV0a4zf3ZTF8YceYmz7
g5bA1zciQII6GFwLnLDbQmsWCVrcLJKlHUaBvbXS4bs0ledVh0RzyKkTzIrH
hpNxnAIRXbV2KKHR1mrzYxKEAbA68E0Z3CdC0LX4pHRL9WxwZ0Pf+sAMnq8z
VW5x5yp7XYO88jWwZwLiFSoMJ2vfImt1c414CM0QHowSizb0NXW+knsMwLq2
dHKgqLrMdbR3H3Ucz1Cf21l5q7v3nPlxcsmGNudvsxbZQZtEZT/jvuBU59aO
bhXVlGlpEo++zYH7PvAh46ck1wevzddV6mbJCmaJr3dQo0hg4Pzr5HcattAF
kUH/8NmuCZ27xSLzV9u8hX9ZabNH0FSTzlsBnlBoZiSlEopN10hb8MOQv1G1
dhpfMiWFnXRLWpoW3bi3Knv+/+8QarCAHZ1Xn+B7oeMqDHQYqxMZ/6xSWUoG
2///P53TKem9g5qhp8KhufdnlkEMQL8CtXtFIw2XjIjBOl4zpkC9bbvXi8Hs
l3M6W6u941ibCV+V9Pi07Zvn3GtC/pI9HIv4w9/sMfpcWDuYP2I55wroiGWf
OIk0nle8sNlRtKK0wD9uxeiszTx2AXcFQokom69EIaeRNU0DUaL0WwQ4tcwS
I8CdUQ9OEfGFDvBU8+cjiOhsSwXca/iCZP/A83Mga0B0Dub1jRLxeS0vLOAV
uZuBvUHEl637SOauLA5rPSXI56Z3iJsBAs7H1kx0qRyhNfDZiQo6V8uA97ix
R4AYD5JwA/RyRC+NLWvPNKxExL/PRK+83sidHOqLJ1l9osGaD+KqeZRA3qld
H1puOG1ngTgqJ9MgtllcxfpcgZNsl03Kg+sNfVR5H0MOuFoNiwRU1tXFVIhx
QJ4BRAnwIQqvTOxu/6g+4RoYLSqxop0T/qvL6MnLTXes+LRp79JmkTfQ0qpS
9F8ajWRFvKdvOovPC68ngBrkRz1YtO3PZHlNN0rR4O83B4RqgSC34M3CieZJ
76E05O2rHz9jNzd9b5U/zHF1DL01xEQnLQItoilJjIF+kHgBTDJ7AVhhBLIQ
gL/bi9vL9qO8TUiSdQ25uf+uXdyyOqaK55WcvLdZ1aURWcIDLIwFxaUoNVPc
6ZpBs0e+Fb8lpLVX6XeA1jgG0R0n8tO5pGZ2e4crKqCD9uIu2xx00Ek7LhWf
CoRdUz5FYCRybBCWbi+5H80SodQZg6no07qcc2HUP7gQpPJGhECx4dev8OZp
+Vesp4ENxEdhYcJ93kTdNOkHzEIn4SP5JtEKV2GMM8/KHCO1MnKoMPGRd47L
OKL2F5Sxlx55oA5mJ7dKWuvoLp24AaC7bwRulxQJ/fqd4qPOlymLZqklD7YF
63Rd4+HkKXjrDcnU6EUTb3k0X7ovJaxm657tcPelq++rMzntP5oAIykuHy4o
1euHjVtJnoDKaVLmvb+x/1sYJkXb4NaCjXUsJbCWcLXI5XNUWX67fbv+HxZA
LaN1hSaq75QfsBobgws28mvr2cpR5RoSP+DP4pD0ehMRQ8Rz04/gyKhkvaJ0
69K5E5+Gnr3NVCWGanaOvZDqEFGUfp8gYwY8HMxrAZxDDBFysF84mPMSQ/5Z
l4Ai1kKSBwUAF0onmgF1t2WQ5X7/fQCDWaX2PU9s3mZvYxo+YuoFt1IVLSkZ
z+uEk3FtW+X78kp/PSatS8W+vq0fxBj8Lhee0uDM22xUsfSfZ2JeQDN3hD/B
GNyn+aLfIu9cPwyvsgsH3EYJi7mk/QBXAEicE09loRNG3xAho/HLgOvLWU5k
1fzrzxDJDhrC2R9DM/Jc8Hxvphk3CupeV+EM4/BITDprfe84rPxr1UuTj76d
Qm8xDwcJJVcKmSclpWf16rc26VlgJgYiQfU2n9iO/GbL9vDDgMNmMnk7WDTr
ghjBsr0+4k9fRmL20zDcTqDg+jVDJxJ1gU4yf6BeoN3TybZuxC/e6p34eQQN
RZ8pE24EosMpL4JTx9WotTkgWYT7o1qeA8R73HIFAEF6HQ2rI+uRPaSPfXx2
a7xQloZ7zBMukhXCtFv+oemWqnVbMCqMeoVZVAiJD0h8NPz2Vjl44hR+zpz7
AWuYviL+NHWmaatOjztPA1EFmC3s0Qcr0pzzgtu1nUhnlry3vv3ypJwxK3xJ
M5ivdgalDCYkq0YD4ItFjfIF41VNcYUw4TwVLLSoLBXdr0bQQpHemU0rWDGz
9VMVveDltKQAW59yvucnN/xMDQWTwnpuKI4QOARnGshWvHZDcuATNrYWqj9h
fmO/SVKUqj/bG0c40lkJyulI9FfxZj3sJf8Dvxie0GlZptKvgdJvaXVNXuA5
hth9G67ZMhao7qWT1svHHLogPs2Zg3+bOyQG4MAdc7+6WxA6TrcHU1HaMHiy
QViymkSXvFiMIRo6TNhwZPNE57RYOcw6lbLWdWUzMPGawuJ6RbF8YXJB/sPs
3PxjABxNhAEbn2/QhOgUPHfqwdrww+dbRZsDhz2AQTxIliVkBP3pD24RZG2P
tBM7HSoltsNqGHiFLxteLT/fju7bUYNqySkjNXY1pafpzgSVNQzCda4nXly/
tBXA9aIcMQfzMpq+rbx0ZDxeCw6C/Trgbg3iX3UpEdq9lyegdEeWXBkYOEpp
2s8vNE88U0yBNroGYl7bWHS6MIfqIg8JGhwPpJ3bSDocdqN8j/bGBlB+a0gV
yuIFeCLD4oUguVZJwxidP+gTqCgDUvsr+KGxwhDtoCf6kIQb+aSigL+NK7Wp
Pg0xJqtQJDXCalG3ohZhh7/zuBuTVmabwhvJwtlowp0oDLP+hs32tsDSPTz6
cdYQDqGssTloW9rq62SjNXtKu0Cxb7fTUN1+DztG154MJabPXYxzCWKQYFRp
xCS9Mf6seZp1flxswdFkruYVHGgPR8dRYYo4GYwZx1wgLZMrsv+Fp6Rq+fCQ
0424NwozND41egJ3QWT0p6ASlDWWPH7W5CbZZZU+VCcXSb3yrORIUxglgWLF
EkA5PF7xD02ucWtc+s/fjn2AMnKJSpJ3tNZZyoPiiRxjyhEEbv03dMdciM3f
2DCFSi5BbagKeOIkVd89V2zQ48cFkBPJ/5oGI+un71squuNaHZlqmhgbYBQX
rSnpgT+A3FZom/6oGrz88wDZ3SRTnVubSHtIpGMEL0sHv/oQmqoghzALcK1D
+vezOxOmBY0UVT3/5DpK48kJ9BGx1HbDoo9pQDIMtcoXagul0WDrcbDYQV+w
1UWVXtb4FE43c3OIpn7Sx0nuxX7pz/n9yVSD/w5jSEtg1iOQHR/QVLIIdjZw
bgiGhiNgpqq97pwkR56orHYY+fn2JTeNhb5GyALNOHYO4/XM8atMna6humkM
wqotU4dBqyTctu53w234mXHh5tWkv13Uww5kNkhEpwVyYavb9oC1ECf6qUeb
pnxbmKXFUeHGAnAUkQXz0bxuRjeEa3uOpchRBkfpsJUg66halcEp5t8rtdti
Y4YciG8s/eWiejiGrTBF2fg6TmosE6oGSoFk8oIW9T/Bok/Pk1uGCa6w+9AD
yIOm3+YTROzX9B7I6lkFIRScHdJ7TR0m/8MZen9k+9hftRCRPNVjaFnJn8Gy
Lj5BME2Gk7JWZXb3ZwFIMb8rPCJfD+AIbQrM+0AclP1d4FJSRNt51GC+SlWY
d7XEwBdzkRPzQi/1J6jFPKIKwiSqX+0jkcUY6Oa7faRQj6eZer2GHKtzKPOK
YRtJ+q18tww78hfQTLHIZIQ8T+HYyZmpmiigkHa+ldskI8oX7eYPbpdQILQ8
Bt8l8DNjJn4AvZiVZ42bQ/NoYVzpDML/38dan1G4R7fVLc1r7h5a1fXSjRun
A5TabRHoCw2XDX8R3w8OC2qvPlKbATpjsJNUPuCz4t4N+LwXpT3Mvu5Egetr
wuH3tUVZp5WSJscxItzeVQw8+wlRZq34jPQ6mOegbaK2pJzRJymyQOb6Vpio
Vljc5Etk7fyBPTnwGpIqy2Xo4OUsankjkZE644nbazBcGjpH7f23CVepcUnE
CpJkiU7Xn7XlOZ069VUxNzf6cGEMxRpxC9KmRiCEptdFghBRkZJRx9gLq31F
s3BivJ61zARKux29jztvikNl7ChGNlGEe/NGUQdqFVvyKB+rc3RreyfvtVTB
zPtScjzWn4RPRa+1uYAO52UP9dAu8AsHMmEK8pIadGWLNbi7N5BZ9EmnYMPu
eoIQTymr8ISYhmptxOCu8nGLeQZx3pI4SH9PDvir8Im4zUzctMa/Mi8FT8EB
K/JW8KW9lb41yOlOfCtWNNpcRp0E8BzN+5h4MwgugcSAh83lPliFfWna5RGl
0iS1jjWFhrrx04EXmYJlTZDVq0nmGhHhkdl1nE0bga321aQJZZaPBEI5a8IZ
gG3LmEcg0nI6+hzmHlQ+JN1ViQCbea6vtWRadP6usJNAQhSxZ2onF1H4sxm7
QpzMetB3/IV+egnvouPtUMDJiiGLid221JETzdULYcTEQOyBqpPOo7+pvnGM
IN4w5/moPs2Up73P4ce649/G11f/rdJUmeMPmN9fmK+iAHF/hN0OKgF90/Xp
tgmR1pouuuZAS1ucELo7El2hAqA4jOlsc/MVozyIfm6Cs2lkSQSS+v5webfB
Hnc54ruowTN1N2Zf/kF30RKVnWyRYWRDzSiGVw0lq06vKwjhhWy0DY29uW7U
DZK9FUYbK+5zY0kZJ9BZmWUyfGaWwAPIwdf0Ku2P1f/89buztyBoi5sRBXRY
pJOs+437Qkm2KBQChWzgvFClS+WEOTf0bFvrrUMCUvsGW89Z+b52nCBwZawc
Ov+dS05+VFnVm810pnA1pXDEdqPkZobAnmt39n+HR9OvmlFm75esTdPhH5xR
7VhBFOwtYKjPjq8sP0pXbvPym4dCPHpoCBfDGXluyrxTfBfQjilEPejozWdX
Ow5kYM4+fgFPyZF0iQ04F9bjgO9HT1GlHNBx4Rpc830XyW/RQ9I9xV8uzOzJ
Dd6pfyUWRR7lN1KKvsrse9bZ5lwrYynau3XPiEAk6dbHtqbrT9VJbktS52gH
oF4ng8D01miOezgrGmiUHtZ3tppSZBFPuBlyNaPoI3K6jUgmbyE9MYSCbVSt
B4Etg5H6Z6toZoxE03nDLChPeRQ1W/CM5EUPlfZsI1KbUWJ/L8lhiB6srpyi
/dkvyryOTWJuSKCpaPv1CR/JOm80YxUbj1UjfsZJwy3El/+BYn57OrKA0qPI
Sah9sLT/1OlExTHC/K3d89lRWmMzxXoTQKohz2MN6INQocDWQHd/0RgFieQb
CuwkdVN1SARM18MmTpscYgebBT0jbUmIMxiOkME4Tz4m6IokP9bzpFyjVzcV
J3ay22CmFc8JMujtpKnJL6upbADRA5Npsiaw7+UOdbrRXdvFxHdB1HSN6GEz
mOFfvhASo6GpMpP0DwKIVdlB4bOZGpKxgRHaRmrpVsu6in8m3bqljkRqSb66
CxXIW8/TaRbQ9LamOB/JBZQgOtx66f8e3mLY9EoyNePnoI7fZYc/X8sjHn+5
QKbuuMpPXBVYEnEoJoxbPJ09hOILEeEEpvwF486OR/zVMuDJ1NRL2+h5sIYA
HX0XUN5XcPs3Xw2YIZnKlghbeQZn/OtyE+rRh92ZIWs5K14cJo1qyP7q9jFE
PAO3Mrf6Q6Ond5YIThbR3br5o2KCsHmFeHCX7e/i5K3V4jBxrI/f+V5lMwpx
VKNj1TRbB9fEpiCB2nacWwoNt1Z5eIyFB0htFOTVgrNroIkVGmQuEhROTcXO
hHVX0q0WS2OLN8wbqo1geEEveddrj3FtGiyN0sxL4c5OPfD/2b5lbu/cVEOl
fd/TNkF7Y7nbC0KN33VpdWPTJHojjCn/q1EogUOtas/X0lAlIsqUJtBGbYkT
FfEK4VKzuI6WgxgBRVPkn9rE2uY6P3sfu+/TB9XtaFlDHWmglHQHnCQ5as2h
TEr4xQ3IdXhvosYsy6GPX0ZUu+J6j99iO/xpvp6mfo2pvVpetrsL1tGn8wiv
rwjjkUfXWFU/SdI2omuexJ9sm3ny/3rzqi90v5iSn5AF+7WVltYOp3OzYlut
PLUbO6KmZglbDu2RYUDxuw0gx6z6oAimvCPsfvGeAzzgxGIeyeco0xzf/KoG
8dsJU3YwaS7T8H9r/iwCXQxr923Nzw55IXtviez6/IMALjIIwsESqrQCBw1q
LSF+a1dP20KRJqu8hxunQ4FCYzCPlGawUsraj30iH2AragJpoeleZJ6Zm94J
t2/N+BzMl4HXFf1Po3/GOu6xFkhd4OSY6dazTs3/bQjmf+sqdGItmB2okmDC
XowtPp4RPHDJIBnGkSorKo+ux3t28R7n3Gl4huC7rgduCkvywvhC8LadML43
KAuGW5k5IfzSBEDzm/QX56I6eD2ElJte+qNeXyTaamF7+opkhOesKZNDyGlP
obYIOOLgAJmu1PRH8mJY8FffTE4a4ATn0cDz6QkXIFg8z0/OJJp6I9DM3TXA
EcYwOm5bFMK+wdK+50xEP0uY3EP0v4eWFOMrbgAz9+eOGS65TBNhxJz9Vk9L
ppUEDAV9HxFYA0M9PRyy7QfVNc9j+W4pPdIKfPYQK3FpFBcSjClJtfYFMVx8
XsqdlFVntfZEW8Ph/cFgcoNZtQ+bujlJ2irqGPmzP+gcxK0+ZQjIOZokQSC2
D7CL3ktfI4vLo1rur6AW+sKvKG77pzDHv6MBO9db0JybIy8xxsJZFPltSdUI
wfJf1LTec/2IBITObv231ZxjQYGkIOkWN5b0HmQAZfvU7aWWk+F6vUsKibsu
kbC3dUONf+OMdONTEo0fWCCF+VTRNVugXgn43RWBJz4gw7XPjs7Pu98hpPyn
cM9wCWIj1w/YNtJiCxytL/WrPevdh2+V/TIl7rV8WRVPxaf5wNzgZdehTnQ0
JoOnMBRY7qq6yZ6pdjlsU6yX6r9t2YnDQWdUFz/Pc6D+2NyUjeL6M5uexquT
i5KLytK1aLp0CDQ7sTxuVIfvpEEXVexuGAkSawHuocvO9YLoEbq1HNAcOLUF
vO3ab9w1qzxsv1IzoJXE8KXaRWXzYRnSV7TdPfHhd3OzVogNOM30uViMQTSc
cHpu+tP9J6aFISfUNIsByiWf2lL1S46USMyLC+rI9dXWPhg4EgwNqO8MWJv3
XO1wq8QDIj6zbdI+JhQKBmghJZ7yB0bfHE1jqZdn5ql2ZjI1wXQX9IakRDDV
+bEhpWZkJX5JjVspRDauzjWJ0NyeN4FF6fhAdTqAizkaqVjYKTxT+GA+rH+R
BX+hGlhsfbGyExOAIe0xCiR1hPDzGbYZsmreANPn1qY/GJBcBHSXPgsMKzh8
kQuo1tiZqki3HEXAl+q++Y199BClN+lDEsT4CB6El9zC9HZo3NuxBpVc06tX
K0+Nc6SUVbsrundkcB2T5zh727/PducxXQoOIrMQp3xuw764NQcjXfZnKEQQ
vwXosXEaFk4R+aUIFt0OR7NSxmLyMNcveealInUJITntAkuIsqv3qktIIfRz
s/i0HgxNHHgaFqojMlegRLYeW0Ffl5L8uR31U9ahv/eSMLSvSyq7uQv5cAtJ
08rE1v1wTB03Kflhmhgu9uUzAesaErjHNbL3Smc3gtdqbeju8RFwGymM4tdH
BnykGHWDBTzcvDKNy9SzRzWV7S/T2f+dDLwp7vXOWbGXwWwPZxUbdQCAlWF4
/ioNetTX12og6X5UlKiE6KYgL7WiXGrcK0dtcPiGdUj7JgTl1SgYtO+CaxCw
C9Q45K7tdEraZGS1uVcI8IZJA1K9LDLC2vnESIHW0natLLzRJ6zLez2cMzQ8
OkS5Da3pDL5kSDoiuIjk+ARpkM7z7VtURFI5+riNLbJvwc4F9z0YSY+gHVIx
RLzppX4BZeDQENLMRJ4gFfx+wre8VIR94R13nstB5lfVI4J7JymtyLzj9TKH
n02Xril7dIP/qnPuhY0eR4cZLLmfPKabVDqAZ7l6jiOyLYFxiwjqlhrIlv2h
1HVrRQE4gTjFONmSbe5bG1zwnZ0fRt0CotAqvIzMqEwELowOJ/YVzeAyza6J
Xtio/GG4M8+I4UiMJc8QKTfFZM1r4Vmj/jmypQFoLSnaOB4OJIKunlhxRfeC
leUzzZfhfvkU4hUYY/GWwWoATBvMJkThFqbewPK7TougG4j4AiAibIppfCAW
AhoXIgy+9/wtGULj5dl9GRrk3jfATdh01/TlxlIim0M3zgEmGoppiZwzlqCA
LQPMj5UOf/E13i+gVhUTA03LJTDxdko/CVUuxX+DfIyP8n2g9napGrcrMjr+
4FFVzO/VxErB4yJszMVP9VBz3w8F1BsXoJ+fuLSobbNXuutenIsG0ojtDu/w
MRMoFS1+q2yxQyo1HfUJpUwUTM6+KDIi3BXvJImJscSbUh4YWe934vMs7WZ0
MO06ggDz6IALhHTuN3jF61OKjAaYhggr91B5sjvdZXhrS+3uon4H+/zykBzi
KssNQlXBoILl41QCBR4ce9ir4y/xU0qGmgS13RgGOgESnDeelSicdI+ZqbQK
P0DZGL83RB3Sd0xXYpwjPXvGIUWpgzyTFJTK9zZM4BCjlIjKsulzRMUvo0Sp
Gho0q+kbqIn87ngFLIlaV/7Rtk9qL/bxOmi0HYSVA4p8YLzPdfBixfdzMk6u
Z+zSJK1DWR/K7AVejqCfhPIlkgi1JiTmra6Ty/M4tXsL3LfZ6LhH+DItkxzn
XtqFDYCCXIFnU7c8DjFSfhjXPEoTA+xzhjVFIqgwTnNHuU8kWhIJ7Gi3lQBI
cltXzPhePpgrIuWChyF4qmnBU+j8s5IfxMbYuKM6Usz3kWo3qjG+JAEiRUTf
a9arRglztimkHzaQsuZmUta7+Zv313aWhY0Z2KEhQ6+O/d/I6dCCrIA3vT0T
wWFCUR9yFvWsFXL5lKAvI1Xx/WGt2GVeWoshlaACMOAaXdOLPoDHfl8Oauc2
hr/3jNr0RyqxufIvFG77XkX51u8b7j7DMHwJhmI/njmeXddsHK08XT3Dtigg
cy2elK1XfsL431Y/41rfUDAiyqQCE0OToXacAEe8TZuQEQ5I+l+Alir6scY+
Y2z0LMojcJkiZjM5Ila4NEBC9DO/MuCdKV9DAke5itznMDobYGPr/PwSzv4M
/AusNo1hhAsc1V9YXAd8aMjK5rBXzisXtuv7APYvLWcFckXznTNIOdpAtunM
qbJjPpKLf2uGgk0NfZxFhXLsli+QJqvPRFQUaesftWXMTc1svQRYdWSnVgHp
FD5OZ8sqECnbE80KFaqGmaenIVtN1XiHbJ7B583y+70i4xPAlxZQkqZvv3n/
2w7tYyzi+kooAz9OFnOe5rKQ8wfdaT9XT2dKufHkhe2Y3RQ2h6dfB9/XRhYw
N/ymf2sRpGpj4bCxE8RIzISN8nfq9Oc/Fm7V7I13zgYVAmTMPudTFvb+kc/+
+95cBJDeA6l7WltA9vm/R7p0KuOQ17ki6tUxEA+LUNjil4AmZdSZWenyQOcO
VSmilWaln6ZgYlzTLjEiBxgPgdi0ixjIGzFWdx33MON/DJ7I/3UDU3OFzpnL
KRyZcEguoNdkwQzIhH0qfZbV3RfgEafXe0QgvnsoJXeKCOIsusBIiOU3EEP0
54wYYRpkgt/wZRrQ8caAd46/Rn3W++BFT7KoTN4zQd/uUb06qGFKz5sFKJIT
WlZWuE3YF8DMeefpIIXo9afEy3svsAA073WuRrTr9OjNUrSA8j6LuNF3t+wh
bJ9BRxMKOpTjtujML+4waf2tKOmPwS/ssFljuhmoAY3rNEC/7821qlCtjt7L
EkxHEBSBLWFuUNzsL0B9FMrgLu8fZpiSn6GrJNrMxbMQyVy9C9edkPvAoxVT
BD5F90TT02vQWPhqQO81O3zG0k+D/jExkwz24aFnROPx4Ilqdg5LRE9oQLLm
Y3m7K0YFAu8qT1rQvAHdTwQ7AWnJrSbxDIDmto6V3Pa7bfTVhwZGn4hihgzW
jXuwIicEE3gn0IuRMb8CdbF9Q468gy0gFm9jHiPWQg2wQEWP7swuS77tXzVA
abECAHUCv1vcQl/RUIrbUCM3k8ND+GgHgft1lveHCJC+F3BQ8Xa/+3VhtAqH
qQvB28L65ztm0vgfe5scYz+GqkcrNrTTMeLUCBRx9hneCIPC53j6tGg4U3oM
eHLzZjn1wiDYQrSmMD5qc7AyJgLza8KaoLVl+x8KbotW1+QPqvMzm7eyr3a7
2bH5HHbiATWMcv6EPoo78OSWFi3H4Jn2d3r85QOMt+y3HBp+oqKVSu4xqqL0
61WA0hR4d5m3NuoPu2JjTynMONCpX+r1g9TmMvlchPlUkk7yO0yuiUPGk2e+
MNRr5m+uBgAdKiI15eZw2kP2Ylq4YrboMafMAixLIUR34KQP1X3LZKuUYsp5
vXDiCPwTNv2dYPkBD7DceMYw3Et4ANpLLzJW+V+GYuNCt5Ivb47uEBqDrbmd
dn1TTCWwdVRAQAKQKJKoiwfX2t6R+x+OY6/cF4BLKA7BT3U/a1Em8wKeH187
enQbeR5KWtAttGIT79z1CO/E2AMT3lSk447aqkkfyHvo2eQRbQ6jox1Yz+33
Nn3h+qPmhMEr9YLF+8Uw/SKBYWYITbEhPuBNkFvl7UTTW2H/hQt08Vw3Jt9x
uVN/H+MTOLXS/MYVTU6O8ExEisPg++fVbLE7HIr4YpJrXDWE9FRSKbdDvfJQ
P84bSJHoD3WUtdPeATPfxz/klunN4Ulixw+un0WcI07HlA2YjDiG1VibBUZr
LSZiP1ccjYD1nMKJSmkJ1POD8lxSqHg0jc6NJgoLu346AhmZcVeG2Nlax5zk
20E2j8wWV2QkYEnoCojUbtWtcB2oIGHcej4i6PcFxd6Oeku/k4WIbYikRW+s
LFOS3VNj+rTQLfXtyJWtm2AkBZU3X1g0STOEVy1iVw0vW17Aom1qFaxiyDOy
IjdC+JKX7O2ueKppvYoKieEJgvyW/GQA6H9ZXDhULr/FKJA931HyjKXqWMH/
Xux+cxULLLFDFaEydeaYxOTS9f3SV3m8ipIq6gP+t9j/a+r0u6PjQkA5s5uh
mcp0D5TVo+cB4j5xyCD2alsjo4Vdx3TNo4qqxmPJhmjKA2zlkEgVX3utcuo/
YaPl2H6hSszicaEWSfqJwZXdfVcmisP5uGUeOa7C4He/3J2dU28c6sAxz8BO
NgX9NJsLRJMuEw+A3FCDCxOHAMLSHnxPTNg4su6PH3xW2gbMTjxzXYgYH9g6
tI1jfmE67npK8K5y4W0JFf36zhGj9jupXNKm+fEFG093y+0Z6vEsHdzMpPbR
JSLicO9aH/wK61GS0Sl1ttn0G58gN0HBXl+jgd8dTEkrbkdr/G+W5yS9M0TK
+Mjxf3qJLuStlTcrgg2m6SgHK4Q1jNabRyrYzzLLDicWmDKkD2VSnxI84uGE
bmKt7lvXpSbOLUFfU73HMB5By17dYKMDQKWGsk5wd/axn4ugyq4YA8W3JeT3
NYDoj22Nv3lP7k/FvDDrrmKLejqfH0xR8OmJfASTSEOgZu9TRserGG4mlsmV
onZryJV9RtJjIPNYOiZGB67BstSJaDGK3tmkY5mvKelyjCm4NoMtpk3IY2w3
zs938Ymo1yLOT3EyyS72vOe6tbN5MxFhz8ankryJ83I4+D43CFGJEA+PD/MI
/ZztyyTE2FdNQ8qHa4NFNUayq51mS4ZFme621iyEAk/jA9Z7oXQrUIiFq4IO
KhnbLKge+5I9ESjw++IyLU6W2rtc91vcEDFCAF+yhpCumKlOjCplP/hTw9f3
64Hsa6uEm+oUXOdKQrxV8YC2reThMO/eB8OEUaqtnVE4CJHSZw4SHb/hjIRP
//Gmvne0sZYCHFsf0KKWnUy6uBok9azhYeeVlZLIQXF2k/ibBStCF+hxtAnV
B/u0UFuv1ZJM31j1ey0tkCCOvlEEXzZhl8w/uewmxihb2o3GoP9ZmOXzVMgZ
FpIfLPtSw5/RUNMI1mhmqtGcmHA4AR/cz3UmBuNtbZ9YB8/aaSjB6F0+3iLj
iqoaRhajrVNBggPgBVF+l6v7xyRUj64KhRyXi46uAdZ6XndQHc1cvGfKa38v
gu/f73vkZ0k8Nxd2rdQjVizw27oFuhhvSQ3X6QomnLfP6K4sWEgKyJDHAy6y
jNcfYwl/X2RsiO52Al+18NAgf45wqOJCjiU+QUkWx7Sqf8FIwSMvDZ+K6OiG
tZLtYTNX2UANvW6d+xsJNB4gLZjxYstW6Vzvj6eQod9lHEMEJfKT7a3d3v8z
8lm2POgZyLUV0N9+6XtS4VupUhtkTMGUSY59HXNXvSoZ3faqtQ/p8GKGQ+zn
EZ7es4gvM8P4PGtjtCaA805UB3jnXtt2A2MVWLkqLAQu0/feTwwY7dNFLrIX
IxzLj2bSPB/qbi3IXjW/Ubb/YA3yPJqUcnjWy33TctzEUC84XWkMT05qe8sW
PrEEyCiGIuO/lGTj7+sDoVyZ9hw+pBkHg7kjjUjdSFRu+hjl6F2iGADkdCSQ
QWKOJDsx02QS7g0FvuWFSXnYVYV+d8PcECkj1TC7Q7YyRs15gRTm47lbnMAO
Y8c79sdSBYIbuBQwSfGz4ohjx8aw3AUTUIhHRy0EFh5Z9qd4/Mf3Q+MGJlLJ
K4iFb/IB6R/klT/doiX8y/5vYI1AnRvUvbBthqTikkqSl48zocuTuL51ChWg
Ig3CoNBg+Llbnb9/HMxjp7erZub0UDI41bCcixlZ9awQbE+USf1J2Kgz0VtG
Jk3JTGa2ENBhLA98Z+NsMyF/x3tYRx6Qa7+PIbFA+kB6BkaHwsH7smoSYIVE
XOSQm+tOCxLbX4yxvY5JP7ysP+TE3xHORH5DlASFenSikQxrkLnAZF1uc1mD
JU+7G2S1wG0SWee5eq+OLTFaP8yxjR6pb/7OEhWVd2lU2DpiiOSGfPRTiuFI
r5FtjIVM0qzo6Dp1Jjz+8ICGDPH3Uq9nr18cUXoIX+OpMKDc6RcENHQDS3ZA
9KdhSzMVoHPAefuAhBLHfAmWHSiFjHrLOmHUdPE3sN/u9BhMVRZtYgq1TCco
JYzrJjrIltITgVOHUDogaz+16uWxJJbLW97NSUjh50gaC4jfYt4/fFu3JPDV
aIl6qEtmQ4p4VzZUkoernbQVBnlBKPypgRqgwvWxaf+AYjs/Q8q0Ykua4XwZ
yFttJ5nwiHxkxkDvI77AzzIsUuFQgtEZ/VlnXEQoyJdNqdfZM0pASEDkBQLl
zwQ2MAFTmndiXflnM0Nqx3Ff2FxJFGaPObaSFGm6VWrYZ5REWnrWpv2zb9ix
niQuoojyVt1NYk1T5UMafLuw7cMSgV3kjpurr0QHY36EFhWUMHOuuuDGvyoB
35GUZs6UPlmB0UrglJbjlo4YTNUzoML4FSQz9x4gdN5xoyGq3QEzwNgreWEE
bN2vqKr3MUN6k9uJEiHWmLART/2yoFp1JT4e6+3G7/61a76D0QmDhS7zsh1N
QIspqf6EY0u+ga//nd9HsZSKBB6ruIWj0bFbR3gdtQrm8qd0WfvwEnBfpAoD
c5GPf+jVHdgEPls7JmizReAhrgXi/EmqbRKasIVvbBdwxMyWDUO0jK+0IlC8
yTuB5u0nz/AH6TcjcBIsNvvbbyGy6yhLkBumTfBZRbPPbjp5g62rTOv/gbCz
61YN4mnTJX2SHJtSqeZZz6PjosEu4gxPFQKsTHV5pzBV2DXo09dm84l4MoTM
/lSJwNY/sp3laeKIvJPdGFOm3Dpv7RktpeBLoYnymZwDd6Sc4OxbQExdeOMX
tXPENVr2QxSWdowMSbjeRagg+GIru+LV9yGFffVkn0tC2M9uS8QwyPTwvmy+
1Vu5rxQk+Fxh/ddNXt9oBRnU3Pw9OoDe+QD/oNK2nnyeR4Fppe71tY1mgP+V
97v2OjkVna+67iGVB3oam22iOYafLB1Eub0/nShYbFsWEdDUGjlsfAf+nGFI
lF4sGRJutvnRnfLVVPbzliIWFoh+05Z9X4laTnUn75lAIae5ic/zM9emziZm
V5sspYvJMBM/3NwFtjrQ5AB1ShJoNNLwv6vuzLUQfd2vmN+b3RYLEE2LHpQH
qVbcPHytsR2XEuRkRZlj7uyykYaNjKOwe/1cOJv7rjuSYqECMY81bUk/lgAh
B8/wjmJTIu99HEvaiCMFsdryTT9xwO6aoLfERPVoKNPaqdAH5Cj9GzTU1Y8L
ix6hObrjQmYE4G7lAxaJQaaVujAEcrANWdDidjEKCI6FI4EUil2bAAPHGsoR
1op743ozHDXL+ED5WpIVOmotWcxrka6enyaTfHDkPrifFSRaJK5nYUwAbuyy
0Ys6YHn7vs87EDAUyIGLBU2rjEQ2CWlVApmSuYGAntVQfjVIUTm9cMCMnCqC
onfLL/l2tBMi4xgALuMh5ajwkFM44q4anSebx1nvopTYhH+hVuYutCClxtk6
LINSnpmlZtx61mbilOfWjqpGrFWUTXAHSFXPJx3+t+tqW8CLWgfkFK6FNdTu
lhX4aMhTiJQXRK/fbfoVH3dGuTSQyEwzFoUTAa5/lDcfupk5zVGfF15UDK84
vEeGr4rxBbkNMprbC/dMVVa8tYhtCP3lYJWDDvHGdzfR2dwYSHtofHJmQhsa
D0ZcMJsRn96Iq/aC+MLmFTHMLL12ujKSSVQG4slLNbqQx5B9AnLsln+/Tpej
ff400Sbzm7mHPXAlN33BiFwdoSwzAl1AXILGTHNf8vbq5b67x2YSfkJSodrY
qNX6nb08xEyJS0NgUteV+X5XKByB1rFbDtfpXG6Wew7400KxlCZ/xNJnBs1R
IJAJvtMEHzltnwFCzXUZOlBHL9n/Mef5oQf2xbhIyzNPxn39emQoUOwIhZUa
j+z3O4bSfpHMmxWU3z8tZMjV0REfKYSoJIazUemOnmu4mXhnS7msYrwXxh7X
SxvDkU9MBLHcjsiQbDn6oJDsFnccxU61JS6AxCYJMfkH4EYk0p6rWNrM6mE3
E9IbXCv3jl9ZnHQV3+VbPVKnX/C+zgBd4nrGbYi1kCm8r84OgNryyY8F6raL
lbhnu9SKzCEgL01U2XtIWphqs7lGWxOUd9i6QkTzLDdj6wZ8TBjbIDzsfSD1
50SgJqnaU3vQDpHDhnOmO2XFkUsR62Y3loB/CbO+I3gomnDusU/NVWGPqUwY
ITFgT3oRXIGEVUxbEOmKbtVgpStn1NLl1TQazYht9BWsoS+D88hr4LtU2uRh
NkCEvlnbRFCT7B4Fmt/sK00uQaWdev88i9g9HODx9xoa9ioxmkD3sfTim/Bp
Aq0AM4ktzlmJA7edY3WVvC0jfMYSPD/mzf+JOUo/Xak2/xjl2uLdd+vRCTJi
YJOB5Tgq1uiT1ZVdn/PeKTDCJbODdOSJ1WCPW4uLmZ0CPKbJQvrpjH+o2eO6
YbMCcd1RKxgGuUCCpiZ1ebATB5C8iaebFMBppD7D1NBlMlmg1sZ5yC5/SHPh
V1FMKq7DFXBtyPS1NqS375BAVuyE5++hghtlY36tuttvUXKQIQklvRj46Lqi
vCWsl0MNvNIBn0c0Np8wb7dSSG3NsfXUOsSs6kNLPsb0PORRDHQFkDbSkPG3
OduLRs1priLud7NYOrMiXao8l2+w2P4YXaNgYbeaaYw9++4RiuIZU1+7Seym
KTimWx4Ft2oxb/hrssE3X05fuR+YOdbQowgEiNHoyRfk+FTHwDGoDhzjv/7z
VfLnbQ0ZKMwwKmo0eeF6tC9BwfgWSYdsd4aG/w+rhHoo+xf333+o2LuobgfE
RUGq0wDs53aguFlYCBlGVbDhDWrEYi3C98yPYarHUIguQb/7giGrmW2xE/o6
27vuoDJrMeoVD03vRiY1x9WGTn7u6fcSELWULoJhPFkXb9fP+2Tj5rUemEyX
ZNUe+WaNxV4jpzxoLM4eQoWZN9BlQ0O7lRvDQ0yTPRK6dg6JUn19BSTa5fRo
TFiZxdZxoV+y1H7OeNQKbqFUh5MVuQN8TPOicJyXw8ZDUgY/Y+GfefWlRRSp
DoulIsdOVs9rbFkVHS1kUq0hJpNU8Qqmj8l562qdHFXRCRgD31DfYzKTjMHS
VGPm0FQDAtPh8FWi5WATZ/0DbsU09j7M9yGU1Z44N3OPlbGA6VCluZWxXoon
+d5h9QyIi1/orfjUw/wGKuJGZJ1/NnrZ/1WFhwfpyFYcWmVufXdL6kf/BGRH
VXFHVQsKBuEFuPeIS6hCUiuc4Urx2eZM+/e29/kOtkbSyN32Modz0SWz0leK
mHKi2/4nNuxfPE6u96Po44MXsk82IcA726l6b2gvxVRshE8OX5cUDEH7+kSN
2zsv8tGM+7vuyWmmFIfHa6GZ4a3TSnELMunbMT91kR34QyQ3Te9U++RaL+sf
sIzAnp8CZ9iskOEODE45NMJikc6fi+vFX8VrLiAtCs3aX/OZPFpoezNykDZ6
77WugRPH1r+fZHDd7L7q9L/05vTPbrxxO2zTnGmc2WZiXJ0xSv0KRQimJe6m
tMC//pGXGuUDdpBIliXQvrBIiRWH00/1wxo5ZWdfB3HdOL2ym4OrK4omv7n8
JcDgpBtfFaZk5A94++eNtZSl/bsRuCyi7HkuTAA/Q/lU2fs/5PE95nHR32Wf
9ZNdeVSK1EvaYeHelajIQyILH2EJ4MRa/HqLXCOEIeaJ3xjunvZZ+GAOfUuE
MLEnjtV0Uzf0Xmzg/Glo9dQ67gLvHQCxez0EToLzljJb19CbXG46hxHnWlyh
N53HvGYuq6bO5Hn9jz9GSs2+yGjOdkYxzJXMuCkT4Nsp94CaKyl3JJLgF/Kn
B81pxl+3iAIiihVHpr8fdRnVKo+9y4lm6tKOCgoK4nRQRIvplimI8c71CwEO
1fnHVDoeI5+RvMUNEDotMttUtAQftX+y9ep4QWZX0dEsbi17aq7f+PwJXKzX
NaHTLBH1GyhbaskZcerlo9oR72Eas9ZRhG0JiC8MGhSk4VGiI1SXOJkgV+3M
wI90aqFQGLkb2iRxGznX2QVB+gU2D8JqGJ2rTPRPDXua9DoN6vfx4r3BSMyu
ooRk8Zrab17DlsHW4u9Hx4J2+fnIxAiNBbcox9uJCygUtE6cA/Xj6uhiLNtf
/JZ1oKpchR6Go+Z5+8RJRTYniFKunZkS3GAPmCEMZKm0rje+dM3CnP2qhvba
KuD+VKoLH+wViPTo3gQT7Fqdl6u0OY0buGiXRBEeloW/IejhlCdPA4fssuQV
ebqOR6nQQF04DFngYGHffBNjCCvqTBx2cylVtBex9HHO5/QOIC2vtb7zzlXW
TtmExYPtdhyrf884Mc/htQKp1wSRV7sJG4bi7stIjedGC1XmWf9hoyBEoSFK
r1lSMw/qHGj5qpY3gt5owIIv5Ze9wFlG41GyBiNgg+JFt05M8JET2vXdiVtl
PyhhIg2Wode+uOMbFHIA0MLwY08/cMnz+U1m5AZAVYgyAlwEqgbC5UJ8fuPc
4Xt1szwlNPbkYjKav999ivCWSzneHHCb5Sb3qaF0lU61KmGKlfHnLoaDBjnP
HIs0euQmBs7dy7MPwJb64t6/C28p/DQEQ9mpTeAt+GvqV860xYLCODkYVjUR
VsSbdqzhTgJcoqOuqmOojqtoB4QyRWsdqmkRsSNcSM3hs+8YC+Kf2rI3VQki
3M9fZEmo4bJlgDaw5c3/XglM97L1ngj/oYgaZ4cDVd/rIEyfOkVwCnvfgWn9
UHxykeeukMLESZUdBhfJLOTLztAKL14ACDnhdMHTbvUwXEEih/NNuMhgN2pH
VGVozDLL3zudD+H4ZKW/2/p5TROEC3PRTL0VnXrb4EBY5RLejDX0iarC2rdv
POkFu14Rqhj/0qhMYak425JNGyaaluVyK9+iT2vWihrv58lQOZOAAcqmHk09
MWSFBrTa/Rf4B8Hx3wLhpofigtWoufu5pw8cp/E3+mFglM8y/RidpkHl18vI
O+k+bptJPzNNs28L1VnWwlyRZnh7c7zHzRFoRylIOwoud5OlpFJ6Btt2cGA7
lKxQDbDnpes7ZUCo4/MFFRTPLuCh7mrawrJfxQGjnINdwmfYGdgM2AO66VVa
aJod4hxdZkL1WbD4piGsVKiuxRXqc3DC1tqN5hdPnrmCbruFizph2f9KdcqI
Oy3o1hP3UG82DqAQeRXIxm6gF6BicFXnQjZzOV62NjwIsdd+OQFpE9UfqD3Q
0jydZMXzknJUrvXPN2rIRkwvxzIC2+2E90ZwKmxM3cmS3AAWMjiRD0LwG/yy
rFZOU0SYs/BektJ6WM91rYlqgsGx5MLs8kA93Nka6tACnX0Hkd2qB+CFmQba
4l0o/0l9XG0MlnsQMYMyvaXi/ksT84qgTCjdqdHdLRez932CWN5KtTKgmIs0
gGWJvXphAKSH/ytJibaOJwMaxn9mVFT7rb+rDUfbfZPMVwFBHA78AxcXMzjn
e1tmqR3zP8oGe/l5aej58poXwDY2b0u5yg7JxaVkdl8o5wHiWnvMSZL81Xew
BLy8Tz9cm+tATgMSsVF3eGZaWXKzTIg45GFWWE05uUFi+IRJXYeDDI9p3h4I
fZHl0B4wEZTF04lZ0u46DA/RumLXrYacZ1HrPD2aWylkhvoL32pygc5x9b7m
X2FvtYpGe0Zj3L2v6Ax05uymI5BeUjTApzyNcMOGTE5eWTskyFZGh5zCIXHY
mYfybIJbvqmYYRdEZtVHpYBGreqzfysc4OkNuuh2LwGZrW7he2PTOV7LPApn
sOZ4LzMeTXBKz0dydAGCyKbsKA6AjTxIEIRYYxcPe0Eu7q59xFOEATnlw9cV
o6Fc4rwz84n74a4H4Z4Rqx+XkRF2AiWTbDYl3hEKaRjhiqOCLrlctG71KOfT
4Pmrc4FMBlR089HyKsKQwwKWAOWGhsR6lc8BAsyIcxITaDD3klNRiNPM8FVy
4aWdhpJbmhIJvVCtn6PFxn6adeXcOsnTaRdAAtjijul9zWRrgfQy9l3h3eQc
caIrYe17wmU1FZH0bozWryMbbLuSLLQaXbdSaU11HEvYGnnAU/M+8mK82H16
oVii5SgHbk3q1l1pDLRyRo2yi4jUjzjDD0fWDB+csi1QtD7Z4X1205afPtOD
qno38Cx5Rmlj2vdfMpIngcniAzXcXVPM/HLj6Nr3HX28w+ZLQhfLmy8lJVC/
U/IlhrN3YcfScoZGa3cR2GMDEh22eLXkT6J1poAVxQVNU6EatTBv+mHBb/mx
d8tbvWSkDfiakoMyC7CCmvN3MMmb1y9NRMf0bItliBeknmiVp3hyAYDRv9IE
h5+FRNvDOTmu6AfwsRYPRPpEdiCuIP7iO0P5RC0go6lIgS152zFG4kHL17RF
kHw3cnUSxVTp0Z0iClJv+7NDXxlngNAx1H7lruy/r4dhVY2iNPReIe+EO35b
/l2wPzXgIlpducQ9mhaZHMi71S0oU0CVzmphzTGcg1rMBK3OfJvw04dC9SoS
iYkktkHzhFS4qOZne/qAQfu0dedZ4MEUTKAK7Z/y/SXMVnoTqNLwtxqj1QmP
jHxekUFnJwsFR+CwN2BAN1hro277nJlygY9c0U6nkiFnuSSGJEtzmYSgu94u
dmdFx9GNk1SJqzltf435x+jXpoiVBbbG+E4r7l5OUPqx80ulxWdoyEkUoyH7
5OMRqeq4DdTlPgXbW329mqW2plznnyWR9nRSziEv4AxM1eGvGwPciQZWZm88
2KD9IE5ZdTwBMjui4+WqLKrZOz8yWhtMk7wNzjnXLxL0PHJVgjLk7GLeluf1
VEcpN8wvdiDUYwB0PvyNaEGrzVZ9W82MTDic1DGIGaR6jecgrblLjY1EGtcB
YSbI0pfc56BF1soFmnQw+9Vc7Zi3NB7fR5fDdXKJ3C37bNz1YD8tgke5VHky
0YNM/KnqRKPCSUioZxHSKExkjzApi93eLf5O2W53j44WrObfeNPslqejDVOu
WVFYnyernvl2oQwQLT9qhvTE84ioZkSX6ObQ8qKVMjE4b4X06xCC5G1aqJ0N
3MPNvDlgg4ErK7raZ6JfYtBC+gvmDK2f8xCgCZPCKnOkI6SKrzfwfBCShUNk
VjEvjBKcNdthBB6dI/Bn4DfFm9v8JzF88kES+rdT+o9BOt3Gnx7/J+dXVX/D
6uT+hLUBaaSJR3yWzW1jm5Ikmk1vM5qr7IzT8c4S6HjXHH7qNAdwuhbW8nPt
2SlE3vHjXWA4ZPs+bJAYjRlm7HXgurzK6SiheAlWzYYR43KSSQDlNR00zknZ
B3l6PxjjstO0cb3t7+GfA3r0Au3RZDG6WpBjOK8KFrIz48EBUgjkoIJfC2xw
+c+1TB4I6as0xgAvqhzbs2WikNkScf+RaJGKoY20LoVi5hxRrItTTS3+Tffk
fzAydxGPPj3SHp14ZUXihANora4pTKIMXfiM9c1nyTmPpG/UEkNwW9DqgdIs
GIkv6Ky2r+ifz5GH/bKkkwF3Ngp4QrnI9RC3/7j23TfLt6ZhrVE2Bwg5CuLy
n0GOdEt9Yt3wlsCY95cN9AAKl2bz07utFYaSozy786E0p5T0Qqih732PCCJs
zyC8lfJ9zULQugTFov0gm/Ye7Pt7Yq4b6YO4dwM0rBo2nX9gvGbBZ1jgx9bB
u8x+p+tSjlTspZ57nVJZoqP7j0wLkVrZ85I2SfGIYYKQSYMBoGSAawTNcFFh
hKkaCr1jZiFEnOjkVCsV6Aaa77iw+lq7UooYcxbRyQ2KLENgjNLwmsDOXMgh
16TiNdhyhPH6OSZK8D+Wsi7Q/KlKLgjSuDHS3tnF6bcOgg6mPiReWWYkR0WZ
z7p/CgRx2Mxsqq7Q5nlMwmUWFKjsNCGiO+UwVQbTAfpwa4ydNa3qKgY2IZaC
nLByoMrQMZe9Gs3Eam+Ebt5/HL2+pekumTJrH2PXTz/7uN9kTyH3yF0ZIabS
uDJvTSr4B5GMcPGd0Eynw3G+r0UDMlVbocki9NDh501PUZIsHqBL+wH2/3er
aCotxouo/V23kWZBfr2UcPn4DbOUrx+yDWVbKz8iO97LnGX7j40/ZRsdR5kK
M3DdC/Z5wpcIldP6jf85N5D50p8HnFw7D7CJPphPcGA0w+4O7YIt/rtnIGbt
O2RxtaEMXDGPv6pUAMb8cgGUuAmIbDR3LWtA4ZqRdSGEf5c6+KL70ebs0jNj
8O5vBMVU2N+frgFCa9KFuGHn4KhFIoPC0C34vNAqmanzyvuzgxug1GDLwn2/
wjgMD3v1tgj7NNq+rhMjg50NekVsTegdpNsKKKHHtZ9FyGCjYQJiV7sKbP62
zGApT5a0+NEGZdWme0vtEMh47oWcErRllP3gueiOKO31fevgbx6fNA93PMaO
TXX9njPxSYGOmlaclzV8pTN6IuMS1PtZmY47Z0P+gcNkT8kuhR/5709hVr/6
CBu4DgFD7CthS6NVhSQYfycooana6IAhmx0RrDTqYxUqp6uf0bitdJEOJ5wn
NPu2cpIQNeczXW0mkuP6/QlhQBIJ1C2VLIQBUrwUXhVctUc7W18YEQwizzbe
bsGZY5JrK103h4ooQN67xHQqvSRhQWeU59S9zLKQaUVXDTTf/h17vT1NQfs1
Ocq7deL787hJ2L5akBYTiMzLNQaA9e8ieysGTUp2oDp6UVLgUmDjBGD6sJVz
N9gl9D8qFOhu/ZHE6o9+IywWjJ0m8SCKo3fjbq6/Tzm0gIyPAK2nh+jqP1j1
5TrC7oqlwLdVNmAHYtjKxUcGj+NlC0ZJ3K8KVsBBpaHYM2CmrVc6N2F+5i4K
Q7//W35a1MM5LdiKNonbdZOtw5l2OiWZ7HfGWASrpBq8OsZhADZKLd581ymo
5vu5Pa8zFOPytuUuL/ahlhsgaVnbpjwmZVjH5udR3dKbVRWG5O+ZvP/QKgO+
W1psK/VvK3l1X16/zvm7Q/AzbYrMqHBRTbdfHykMVp2INRk1YiWBWDggavwu
xTB/kitODiSq42FKGft/ROBlKe4y5dBlw9VaOLtOSVFOsJUv0NVVZNSPve66
/2b1l1+oaAbvuAGSi/w4U+tgzBvq/YTnAolRqS7zOAV9m5NeTwbztA1zsuT9
i9VqBWk7cKMyBHnfUQ8oqgkZWyPE5qNdkrxJLdmmLEWwI9VmjTxJMCJ6bGbJ
itkQteR9LdpKy5jGL1c63hN2KTlVIb0UoxBZIc4ZIlUjL7Mxn7qmszZ2A84o
KGW9yVCFXmceGrY8hbnXODgisyZhzrHrdmUVRUPh/N+s8LqssPfAk6R3OKaN
r/+Re58AcZ0oVy7+Np3Seu2XYAMFczEMR7dtNgDHwGX9hnAzHm7gdRp1qubr
NwvRdk8CnTgPAh6U3KmnZuafd+j/RiPkW48THNIR6J6ZP02Req7FtZ5RHyV0
UMkuD2GZd5ch3NjSwfZzQIzYIFOzXoZGDmc7/6IRJJq3O6n3ipggzR/fDzVn
YiUVdnRFUUPwRWpddgwQClaRQjHCwSS1MTdqxhQxkBQsMrVtr/Dh8wpNexYK
beJE7OATj1Lrci/kecmDK0fDGPW8666T63Pr9RBLOFm4mBcJ0ZlCyQ4D1QX+
IgFtszCAybb4S4jtNInUOfbHemn6LV63tP2eGksGSTia6RsFNn7WQKvsMj8J
WbsEObvwbHj36eqtBzJYp5U2WEjnHmmU71wMPxafVdpJq2DyggYxwzgtQjjX
G1PdLo8G9gJwK61PDxbGm5BLaZI1GMubRlXec8QNEdF7VF4Kl98IuY7e5Yo7
VwjRkykjLY/Y7iFmgUCXU5ju/Lispl+cuE++0AGHjkxh82w0c6XVznryyCrd
9t+Wv/3VzMaDzL6nP8SdUe17woc7TApv1wkaj3l/bVwJfeQw7qXxKVsOXQtt
hUCesG7rU4R5d7MSbz8YMazGlnBPRbP1NKNUFMqHG3H/EoCNrcvvdpz7QVPk
hN1Mm1p2JgK9WI2vNHUEYQMBSjpTNBQobW9mceQhF2tkmAdFO1ysKiPOepa7
xZTfeVGBMkniL9xHRpAUA+5myLUDavqzaJOdDjbwkB3y8TCqovXg6tTDM6/W
RS5M/+n3D1GpD51lItFteriYF74H7Y6nxQaiDE089Nv++8YV/3v4CIqj05nm
RodifgOeIeCS5GdSa9UDiEt0FiFWkMC0vmZuO132cyR8YHHVxaVzAFlbdtio
DpMFkzFgvauB9TzifrDIE0/dixsrVLICmhlRccrGirSScvGEgNo0cvbojU8l
CXHzHVaXu8jehGhSCi1QMYesDYFR67utk+oObALXS2hGDmvxWoHpF074Toc+
4iy2/KAQ905BYVezpwaEBCkqLXXhxRjWgHi/Lx2ouY78gl7XBxeEaGyS0t6o
vKnL+WRO464Qnpr8Sd+qJcNTh1HkgwpU41uiko1L3ogEE+8Xcka+mhKsWAsy
8tEJGQ+59AK+4F2LXeIZdlsPXAjmu9A9TJTk2SELEz80LV5JKzacKJMTiKeO
2sXZsQOinAHJ1Z09ZonM+HS5TwGhIZxpJC9Jf8M/xwrrAGzxoFq/BX/9xelw
kr8Eb+QDWgs60pGcidX4YlT7ksT0N/EeOdrmZ+n9RftlTPBoEP76mI4zcgJ7
n3ZQ+c+FnGFG3N4E3emkkppE4fN6VBieRjCz9XXIQbrzbm5/5zUH/vcoTTRy
0ytZBGlXz1laVbzd5VwUwMLG+FfQ2TxJYe3svUYakW/rHaplV9DL51/8tF+w
o1949R+57WQ9Bi8QVHhkmpqNyPRDD2w+WI8KhgBlcbCRI8MW0/pVKjkHoRoj
VmsFWPPszFh0vUWMgwV2gyMmeBCZ4ZKH6nMJsnTOou/RifbCGKofvQDe75mU
lPO61p/5t7gdDWLtjOW/qI9iGMtjFlz2In5AD/j1my6SL2SCnUVGIjy33rXD
cdrsRS1CqBr1YMgysaMcpSvGS3H0KHLGSa/GvykyEYChSXAD7l4UtZERoxyp
0VXGXh1xOqQn2E2PhO4MESnr7AW5CKH+9ecQ8znszTX8AlrttszhQ8eGKslO
2ksKEU7fJXnWPnACC2dDdsRPdxBwS6Rkw5oZZv0NG7wVZlrTd3OF5mmiE6zI
OCD6DkN3hJPW4qne5gHiCYGHyND9WrHyxP+xgJKFOeveqzvsl2bdhl9gMprx
v9AadtJXPtZxnlju+bZTIrhNhuhlvlyTjOVPV+X7tXwGvkUGAM7ZeAAuhX4j
rLjuXX8cLsxbAUphSZTA/CTHeUg3NI2cfNNNqfI4gUegMtg8aDAR00hSXPcG
/ADoTZPEr+YERVwvpTKUdSmFcmgm77HZh2EN5hjsoBBVxhvsBTIM2APAftJs
2kjQinEQj1OK9fc9fXPvoiXAzXisV948M8TwF6lpye9XKHDeTx6OjbXC/nxq
uFubSM7Ab3ZvEAbf/Nj5NoS3c1K7B+3LrSi+yeA2vb5SDAYkcJSxOwUftjDj
BJOY4KIe2EQTMTe9B1c4lUdt1Y6rpLMpXHN5hiPOuHRkeRPfcQuRO5V8DP6S
DgiuO7Ze534YhJHpPz9KBqtVkf1epQSw/ZJJJWUL0Whic+1ra27F1r3dRyRr
Tev9yJfiUe0GRuGLeg3VsnNoaKmtGMI36KPaysrdHFP1O8hko8cXUstA6EKl
9BNwQxwVlb7h0srq8tl4Er4ON/+0gQcjaqB6l37f5MfAFeePG0TpFtXwwdXq
q+zZ1jygDlUZcRwv7/XZXg47AYV7QNoX3P1oAID6umDY/iPb29JAztm2Ytyt
7/mHZXaPK7zj8o8F9Fu5TR05fa9zn+SLndUUlGbz/yJR7bZVWIoyxsl5+3C1
sJfU5YDYwJFbgCZxOXVjD9t+W93N+xdST3Z1oRefo2Hqnog7ND6qBO63fD5o
2iuIJyjr6F2lziByms6cZQbAehJczd+W6WZJiTaipExK+wo7M95aB9n2sc9/
XYB1qfhERUH2JWnvf0mL4Wh8e3v/fj6WVENz47M+/GA/q9mKg0J1tuja5soS
ao3893ID0vUAd+ccqS10VgqVuwr6+qsYo/TnvTyMorb0e8Pmt63Q09BorTbn
BFMDHwaCjRc9hZ7bLU6toXH8b4pgciwLUAsSufxlkSnV/c2K6OFrJwkwNzWJ
aNnTD4uPRGv+IAZ80b3VeWMR1yb2sRe9Xf+AQ93ELkruG3G1yoYTcI5fRXuZ
EPeBgh0ST2sqEszZdf3Hx4ex8udePwNhcgHWjTxk6mkCQORqAYSMkwbWFgOb
7g3/TJ/kuwe1IxZQTxPC4zNiBRd7APTDbP55ETr5/b/nJvDehY5fbmwfo2B4
kPnZK0LInjIcp6euOyTh6qr+NKgzo1egpuwjytnCPq8sjwdXtymxh98FRXxU
EmjbjRNbWRA5XXcB13UA/7FhrcjgSQju/4MmvE4cV92SWxsDPgo1Um0SIVco
K2UpPcwMD7jVywg6Vg3Jq5MofreFP+uxw8XP/4i2tx9v25+IQRcOvpkcG6iJ
7honYYSlW3bRmSI7bPtG6FrMw/ubAmbkHZkEUAK3r5X+UTibrKPaSnlPaDQ3
XmGDDZs05WG4bOCCt9nX9tGK3Z8VQ2deuoeuoP0CPcVGxUp3XU2AcOslRhcr
m1ActtGwgQmn9DtSlGqOrB1lJXwY/S/s0qWq5M5SpMdNQEU6Lm/czikdABB/
rDep8vdVehZ0949dZjTOsjQ33NYLM8xf4/208VGLb2nU/vlc7R4N1AKR+LKV
k+nHlQA3Yn7HkT05aaP3kvf1RkmA/+FdOmsrFVY78hnJOQKNIxODPQIpISDk
k8MyC6tunoalfDsNQjwBlJixKhharNC0si7Sc/mazL03ktuOsSModucIf5RP
H7BAGezUZTKnuVTGIBv4QJ3O5bSrWO99OCkPqOogjWC/ZfUD487k93C5Sn3J
oWkc9V796qtq7/nTAXtNQTQO4kKMAKkW8/XBLhBrlq7dQVrdZav6C2RLyI6R
kHloxtxf+bjq/t9PSJtvyk6MvaKoXH09msBIzmkqRmJZdGsLP9ncMDmI61Il
13K7OvuKGbu3SUGKAhgLfdw3bwnpuFpyyeuzHR4wfiKCeBzo4vDJeUfc8JgD
aISvFvLtE0CCAxlw497eEdp4QT/+7LV3YBJjH7jQkATMWyHAkwcjDafWpVCH
6xSWQ+dtKOvYUKJqPXL+DUgfgrkVbBd/nP7GKV/ihBu5mRl/LxF5iJT8EYJ5
RyXZvB559/PCotpAw++DD3+t/er0wC4CqKfg1N11hXOpdc8x+OiJUSFzKIQN
rLWYTp/IrurEKUM5fMuSBaADcZIIHMYF7J6iT3fqWDch/5Rv8qUR82mIc3Dt
03ykfpR3Qqh1RAQ0mSUvy3yhNYRNn2YFiAeOxicpCA4pX8+aMPrJkMsuoq0B
xLkWaLmTN5DLrCxbORyH2c9O9MwUA9p3+hMbIPRrOH0NCXya3em4Oq5no3Dm
l8SaoTWgrc4bAUMWMDbiKWd4+iwEHKQXRi0FDg5fR2RFzAj91IlTr5V4usgP
L/I/FtwG9GbV6pGbz4aqQjaO8Qla18g4aAyfKJhU7R9tr0DM5bT4yXQP+ipz
/muRPhuXJXw0k6KENJTN5n7huZHthNY8Q/9c6iFh9f5LTvHGhT9jmpNFq+xR
CXviScpSa6xaNr/AR6kdxIKulG0r0ecYZrA6t+C42J9c+N78sRbwXRKz2ksS
ifKmtb9uKXlizLAnSfAijHZ3zR30EuQuZjvR1iFqRxA5IfbdUqo6HHs9Iq8q
s+5K0GSrfWCKtwEN+f/Gp91WaRP5V1IIGjwM7we7Mi/MbTOcihf13wohzJVw
anIAs7N0BVQNWkNkyTr+sDAUXBWag65h+yb4Gb35X414TKZ3s4R6XLrWPwJN
MjykazCrOrobHXH4/tj8CLhUuw1uVs/XEKtLdtKwA5B86HfiYutpTDxExv73
B6cPnHaj0Jb5dle+/u60U/rFbn0XRhI0a7kdoyeID2Zi858xuEn1vfzDqIQN
mJwRWtrNrNfXNzQWhYTt/3q4c7Gx+ea7M8J1C73jfnZX0OnYwHIwu8zM/Gy9
yUT2vQFDpE07SlW67PtVvruxN9DkvGtWjVDUHLjsnMP5z2SNIs3fHdv7RiOA
bQHnrPYj8Hvb74y41wYSthCY8Ru7rEoYNH/BKGdykfwIkZ0kyrt2ntKPXVOt
ZShHAvR7v3afwOA/MYjybBBJbaPbbCShsWR0GrzRyhEoKBGqIORWT9Fg2ww+
2l2FbzdTR1mRTHB9VXn8eMnd3DR8ZArydzQ3T5B3UFWK+oMfsjYqUPvbN0Rf
LKyLCNno4B/fJzeGjixtY2J8IHV5sSF/4tXzxPGR4HzsIqVlR0UFnNhMblxw
7vs851pvEWG3eJPmBvx4Vy/d1eu+tnk1wHeBGlbxlVyixQ3uO8I5TOjQa/kG
KswIN6s5DpoZMhdpwVzskEbLeIQMQqv83e8Dn+78rKMNzlJ/jtXylgUVwG5S
8I9I09U2kKkNxILYvZa1cSNacqbeqXQsl9ySOV2H/Pof26YiuKfaBUsmzwjz
EZZdQZ/qVHVwzbMIk+VYfNbBYS9DtyJP+NzNHFFAq+w+X2UZbwkJMBtxkVoU
rIGxVr9Fb7ZsWDlAHDF8D9j1dRBczH4FZon5JZClOX+eyH5B9sZVPTYwXIf/
QVytYyOLMixwEhJBvtGnAifDsESeE/8SRwxpi+yc2x7zjHs1kwxkzbPkbbwT
L0IJe8Stnc8CwneY8lctycBZvfyLGiCqKv/Q0yjXi+3eMT5CH+ZjQI0U3QnV
YA3i0tgR7cHiWwNLnxc0cJjebMLoiQi/w+MDX+QoE6Wy/aNMseP/cbCMWh8w
v7VW6nK3Beg3wCBbh3nIcP9Q4yI8c/9GzrtffBszVg1OeVb5uJzkAvi7l4JE
Z+xskoEDqkWG2WiZPNqElKsHiyCXvUQozHi/MsbXioz2bJf9dZyz3n6wmxwt
BkW3yjfV0NkO1LTYydI9YPMWSAnN0NnQKuarydseVi2+KZ76iqXhQNZTMGZW
wHT6BnHZYSjQ0jLnesqrRnX/Eq4h54PX56v0wV04cjrWwhM1uNpmguCHUk4s
LALT0waG3lFp7srZTf3pLAfp/j5UlPjS+mk3JJXNBOrrxmkMW2rdyOO2jbRp
eXRsPa7J1thIJhB1hG/kDM7xQ0juGuCKIcHT+X05H42WNabd6XJtJ+/sw5vP
lVIHGs1IztXJZCRDqf33bdj61kdwngq3R8OcHP7Y4ixhRSuclDGYTG/Y74Jz
270UspqWAal3UVhkolcnufTRtS1mqEkdm/DxLn1MT+1Esx5fCy7stHw+gf71
vmrbFVsmRERnakXMTBQq+BmYJlDJbPcIxDS2NkuBft0tZ1wWGco/s1R6VPTT
wtHRiVKXzc/1NNTqLtWX7/zfUbaJJYc7+MaI964Lsua6ROKKHqE9RXfnHfMn
2VkH7ez9uc6x7Ym8Ntbk9L8UaihQ2TnW9qnaEmlm88M+7Nn6/k5J8uh/at/x
uNMxj5PLJNhWo2INTiiPmW5xeXTvXSZO/wNhSjV9LvLf1CU3r8lLkHxgTDPY
MlPXYvOD0M7gTG/fNd2OTCTfNu/uDpE9PJjUDNlUVC7gU3XXGRuoe30fE+RP
nnFMbmgM72XIz3MjnRLK7HICwvVGUkW6WFYwrsTEx+di9hmiYYxs8UfjU8yx
8DbhZONpbb3uWyrzmsYw8vkLHvw8d9GbBJK0n0zzQYM9I0IswAC2LMpJbAxS
df0vOPiggTEYLj7qpn23H/AWDI1+/HNE2SsrlWLEv+3v5PFBe1DlHgNDncbz
y5TA805e1LH5d/Pj2RgoEiImsGVxYn2X5JIpe3KfH0Vk33bNxpHT2ZOGlKW1
nm2wuq/eSq6wbNrdUdOhXiHMJUqFDmR2zZTEIl6og9KCv9+zJGBNY015e3E5
bAvTx7EoL078+PWpxI01md5s7Z/ejT3io2EQqcFpcZfGtUG9hhp5/IUn8At8
olHDzQnRkqytUKHn2OAP1d3ws3Wl4BbMTFAHTcHFc078NXwR4r3WMf88PD0l
fO1KeW1feovDZoR3yK/6iKsgekt3UeQQ7ujFXFAr9ldkukt7czFhVbhCwM9j
f50eWSDgCIaMqcs5pZpsNuKISGQoHCoTrv6V18tQIEcUG1swivn6fv/ANJKo
Ldu/TZVDcLv+tuiNKIMw577OSDm91pxwK9rpEgfWF2P7r7vfSeboJM+EtgGL
Zgg6crf1OSZr4/kteoYM6kO1b27Ew/y9zR5F7N8qMIFzLDpp0/P7pOzjqXXU
uUAN6g+MC985S08/srgCB5cgEzj05TYvUq+9hzuHFo494TFdkKC9dJpN33S9
KNZctgRCL1A1+hHDiYR7Knu6kVBMnoa4TDFKjVVlGOv+9nlPe0VT4z3yhc2m
ftIfTDsD+CUK+HS25OH8MFgGxo4wNgBchfUKVF0/4aoD2qiTgFTDZemDwgLH
LMiI/VCagz68EwDdEusmE8bEgXSH2LfOtXkqyvcJ8PlOqgdjdn/VZePStYr9
funkmtCT7tbjdJqTZoHRryfb21y4WMtIy1fkYSxH7ipy/3CbYwCxVnWQyRhN
njP054hElWMkML+OL7ZciWIJ0PgBvO1Zws8uLHdgaFh/rl+CzSFH/brlUKKb
9HUCFjuYMRRStNDXq5a/+ZtYWYxSGT+RsTR28iJL0v45aulXhxv88JKjpLZ1
ab0uZ8SusAE/dOwv1bytiz21RSIltTccyEEB0Grj4BEiZ3qO6YxmTHbQewrH
FLQFNlmY+SEm3p2r+hapw3Vz3rJnFnstaLJeVAOk2DDW3b3N7B0sfOYQU3iu
JoFnLXatD5hlNxzb2pUUpK+v9E+/G4mYlzM4EAiUqyeU7onEKpKV41JR9HWF
eoN2piHKI6cEU91AOvR8qYj2HVsItPE4QIqdNArO3oLghLmtMQEddxDZnz3c
eZFq4ow5DxGkYFygRdD4aDTqXTPzHlfbYp9mj5XdOTyYfXbp/VHdtL100H7e
uKkSNsfDDA/Cy78wXVMm/2h1YkB29GyXhtqR+mIUDpMuEmMZV2qiJvYU1bF7
Kfd4BOpktsB4twM8WZXXg/1gwUD9qP/4Z2uwCOaC2SVJyNd6otNzX6xBZILF
3R/RB5zr+mTnTjtKWpTHCQwW714FyOiXQbZRrDCLmqwPCFmA0rMDgbhxIymH
C4c3YBEgTyQEocvT1HFkmItT1q95D1vyYz4v7HCABZNauoK2vlWg5PwrZgG7
YoLjM+loOsHEq5YKceLd+Epj0KxHmZ4cBvtVbbKk3cMCQ+nBBkDAZprLwTL7
l49s42nPmTglEyH5UdJ9/kPn7gngluC+FHDHFUNH8Bt7bBwaQk9LcNXdsc30
eFzGLytHi5WS327TgAeq6PxW6GsfVRzvxCiKMBvNHMxFnCyBpzaFXxGEgni6
E3MAqK6wK7fZzW4W5YFGOZRmUgirLVAyhjrfTnXiFihuxhG29GxLxrEP5jEU
AlCAw+UB7CQiolVl7mA81ND3mrnaQPQv378dt7YhUBl3o8qSt0mMd8Hzg9ZI
IAgSSsFHzFv9qNc63yIqzpH8fuq6PvdR7zhaX4Mjl+81NzYP3g8SGgUyE6P1
qm7nfpzYAjpi3NnC4MwQe09qSojxIX1y7BGdclx/I01R6Mgzu+D08G1boDi7
PCMsIOtbVf5mBPF1rdZIN18TRzEA7pejTGgSDPhg4puxWIrUP242m8sPESkw
8ofBrqFmtDP4jc9CXcTPYfuZcemCMh4lQ3qhbaw42XoRk/Kcfn58CLP3rcF/
2+zhzx6yq/eGx2sAGdQsdmW1dAdnNfIUHK1BEe7SQkUvVOdnUftqJ+N1OrxH
EXjExl6H1obGgE8Q+dG8eO+M/VdZFP2qCpoSmsnR0nK31Ut1wlZJvbPsvTox
ItYCdICumWARvwhpnyhffQlcTqIRWAxj8hnK3ve4bnOgoaTn35X9YR5HIBuL
zHgfjKrPsmkCBg+RVmzzfoA2N6funpJSZMBSVRwoGj7oZZjUaVGWbs2jfhet
Ws+JkwBHv9r2ADi6aSUHklYXDlOlb72kP/VDf7hr8+WiiEqgCOF2EQ909gTv
p9umKykq3jDEttTf6cpKdxMrkto3g1PyaGCO3yTtTk4JZiCxosskJ8nRQe+W
RSkM0sdr1+F+aDW/1PekrGdGQoK+WSFqKYevchuXHA2/n4dRHSGV67YZ+f0u
Cro8oMNA5Gppvg+mAD5VirnjGpK6bBoS0FuxzRai5WtQvNYw1RyhpUJkfnd5
qH+HhWJKQtQikPOcKrGnq6WUeT00XYHA/tAGntdliIRIKyVc3k7XAvb7Ar6Z
r5nh3SPsojGfrfhhtK/bHNzYX70/TdeTsKHWb0AOoPu2wFNskruaiQaZevcn
lvNVIiyJtqpX8JWy+jVxjivU5FhSVbV3L9p/8HX6UEXtbwxHVD7MxJjeQcj7
nydItwC89jCrdNI2qTL33oCxhw8YZAPOl3fabSL8YQ29bhcpqkP25FtrHxbi
ICFldftedN7mKNbHbaWrcwWHYS18vd6bdmsFt56X8tR/e5Y2t3i9+kyDsltQ
v2nEoteQel+x54EmOi1Y66rNy7cQBHWfMzQWeABDL8VkzRBJWmA7AwTvR3pm
vBBRw2A9B30tu5HhdCvTKA/2EY11ks33uRowDqdkJeK016xIC8mFGNTjqlbm
IiX+NgZ0FecVbMskMuKlFbPoxUUIGoj0hUfQlHfBllbrm2YrcaTotfj6L/4t
OBkj3CXtXinjONDlQDcH18r8vXJ9SVGzbgbOU7tc/PO6p0kvnDSfxsWh3yoC
B2fxM1rytd54xw3YcOcyXJ6uD8lsxHJkb4g+eAArVBeTmq6M9zkhUac8v687
qRAaG6NvDYzAYGwZoWpRD1ZQcQR4MSGc2X10nbEyXMO3FLuYxBfNEu4RAXdT
WLFxGypLq57AlOsHD5FplD/wh8c6yuYyDgyQpviAxGYA2zg0tBiY5kgNDudc
vnZdrmvwMMBgUZymW/Vp2TYT6TxZiewCQHzB+m773PKuV+kvqHlUvYzyTFlL
kFyAt4VzwPRh/ziTXrbEyYNbQjmqu55PYL0Y4sxpsGO2R+NICbqQA62krZGV
cJWaocP/rxCwGht3OYG2HTHCOV/fhW4LMoAAW2TLcKhgxq//KW3ynJqp7f9s
j4xzBeS7BZB5avwGFpYs7ceeo4IPH50d6CBQle3hT3qwhXmZb4W9Yfq2K4we
fE/QZZyECoEFbL0lQbDjad8/Wo9cjxdKIKRUk2SCyWIT3lW9Hk2X5oRWnYUs
rH0w/6U0H2B3W5vagmaRr/Jpto715g6tzfcxSogYYJYTh7yqrDiKW5Hw7QQG
yNCLSUVbcj6WVKLt/8zh+2kKx0TIjoeeF81di9K0S4fA85/fDDlg0mKbZ5rB
b1btGhibaRiSATjOjCwFigNHAyDXuqialGHFMKO1gYH4v+v2yo0AKKPNowNd
gxFsUkgWcINn5B87ir/qXSAERNRu08P5eRzTqQNn0AT8N25pmCl3Z78KUS7E
zwB8crbOsdv6y4O3rvQzyl4KJwqABNdW99jTNLpfqASTLuIpQW+6B+n4Ep2r
WHEndDYfOOsys1MA1n0AX8U+VLZ+a97PAeGmH9HjNnn2wkvmAJa1WvXcrLwE
oSdHSJDxgH5LtEAcIJWYdUHwQkrHI70+1AaviyoDqLzM4SVn075dv7Mtrc9f
dLjA9are1Y/RrWGLupGJrI47o4OCJGDvGOM6UtTn+S0qroomhCdq+sIUJi5v
vLyC6VhnAu1WbRRxwakgB6KZT4s4D1e5tsvmhvjpc8IEwkPe0UvXjO7cLcpL
VJAVpYMS25EbxreU1fs+4gALi+8Q6D0VolrzWSywHHm1Jg9N+6jGh0OI21mC
CwAo8ucGS1e/NMyOD3Z6T1uBNjTSV9ANFmw8liVtjGq9r7OhLNy3p4yhiYXB
eV7FvHkBplaHMO3obkxBT9E0Y7zMHmHUav/OFUhoBL22tjo8+9jR6vSLqCyA
mpPwx3BI7wzUcD8d7pOQQiQ64LN+XnTqqg8cXaaYBf36wku4ax6gJdcEBmYs
88xH/0tIutrXc2IeJAHfG4GFzXOn0F8FOCkzyUrHk19I+REw5JSsuvOfByS7
cWF45l7NrshgtdI25XW4Wym0qk1At+0M9VVNwawQJ7p/ax1/Zo+ITKAAwzrl
0ePIBs+i6vJdlN8Bx4AK+aQYhZCn5OwxPpa8O0u6ihtiCddYPGZ1GTonwt7U
Duc8BKqpe0s3gBS8kfNFrlJ+rhMsqbOQEaAvkhtdVt5so1+RbR8teeJhP7Eg
DCL7t5LDey0qYRztHKPU86T78XwyJBGqnLBE1IdisPku34kEmHrOiYZiZsFU
LVIoj0jf3/cjV2mVOs7pROA72OYlRYkRb1ApLxEUQTuR5AyEdwntHi7Nmp27
wJ5sJbYa7Qa1MLXNfk0XIiTXFJRY+XvXOpsMf0KqRtExam4cOYwHzbI9GebO
7iQo9mjcwGFYc1eaEYX5q+wZsld5I5AwJQhZCqCd5SrnpjbIwyKMFJAIAUiD
eMYKaF5VL16dlWyhjyFNHJReJeC2vgjuBYvZzDrJfZ9npX0ehC2B+1t+qeno
JW2Rz2fs63FmNqYqTu/6nXOP0X3pk89tTbSGGT24aJh4Lb/RUMLOAY20R9l9
IqEVSvM5/+MQP8MWA5trBXGnDVKypUdmIjaOqhZsmpJZdLVNVWBcc4EvIWux
YVrEn5YYj7NwS/7YlDwZkpIe2OHjuV1F5XmMKKQ89owGw6KVRNlvkN2qWgjV
KH39LfZ0cNEoc28vfhvgEDoNWTGaHKsMmjHMOYnTSACjfguNwnRK32wiS6nP
vpjm2pi4027o8Z4NDQhp9ERZuoZfWe0QqWYizW/c1nj1HYxR5I3TY34p8tez
pFP/cFCEERSCAe49ssV8fJs1ECTbAqkxAuW/aCznjdwGkbKLOB5OsU+OPufy
tYfoWYYOGEY1bYU//vmp38fzoh2auTMy4zhVmM7+EP470MpAQlAtZoMgHPyD
ucTgPjRDc869nX8iDIJCGJQWOYoOxBZqY/pebnEsVSnsIv3+EFzpUkwTEv6C
k9tE2gdsjW57gH+w7HvV87nv839EnjLoRQULVymjIZJ0FUo7FbXq0X55aJ5Y
eXbOUCnQuaaK51q7Ji1yhz489JfXtJ4NXBiay47e4l5QVF6gmCa7yDYAA/P4
fo+GcPV0Jk2bS0vKBXtuYhUAfVq1sUWxZI9kjz/5lefQ0zLRc+2ThlPz9Wkt
eubRhA8gah577Ry2P9NyjqRMs5pgFfRAujRmdxV9F7B8/mgZtVhGZmD7IwDp
P+8kuO0SI2BPUgZiUhAIPelB1ve3mDL+Ts04JhVT7eWrsdiBDSSvoYS7+U53
aYmmOEhFoaCm28x5o88VsbNFIHHMvWWggoBMCO2C6MkJfNNiqJEkQGsgenz/
Ry+VClvWedFE/zy48kFoLFuO+f3aXlAxTju5DE9vkwVDpYe5JZL0eqQgG+rh
7lgYreW1+F+X3Mzw4L7HuROIfD0TaXYcGOYBzO3kjAfK8LhXISVVge+nWLvQ
iLhQyiERMQjX9yRqFXieO64kYWqe/0yUD8ix08TpadCd86d+U2n4Sq9PGRqj
0TPEUcpRmWR2ZXF1F5EDj5fJuXv1nMMUsWUXd0fMLNKkMCJGLwKg+j0l2f7s
19bn/1ZxztlDF+O7WSblX/Ws3FFraAF/78Qe8kg3rzTT+48bLIDZgvVESjFP
GA10ut/r5uLdisrT98OxHNH/KtOQ38+bhOmMqrBoWyIb/uwq6+kmhhqzoGPF
nuaEe7EslP86EMGVPQ1d6V0842wllMl20aS5eu9U0NvcyuCiiEiO5e1sK0u5
98OlAC6q9FX1iserZmqb5O+blHU9eyl8fLX+GYZtsNvV+NJMDhLAG7ylYiWr
2d1ifVOGlHTasirMeKbGsXbDmHfJtIp9jZoAeLHXlFLhL6D9Bt6Tw+8/kjVh
FzqJdLhkVElraCi6bpBdsH2EgHrWIoIJkBIIkX2nM3vstSwFL0Re8Sqa6NlM
9hGt1JLjzdDTrCAyp+hq7RD4I+avpj1zR5z4MvkjZ2cmbfD2W4ofjzDCZYCQ
gg/jr1Rjdkvgaj5KzMTZdjIVt3PCm2jnEwOA1huPllxfeE8IMBXZrsXMsEOl
tuj/E1rnSHb0O2CCPIq1a3WGyWEnNXYccHqGeNkDFP9Cq8TceT/YMEfZsxlV
SUis5ml4Xn71fdKUlHL0TOX4pjdxbIR7q57SAeD6Fw/okBhLXKzxa3mi9tk9
RzUMZqN+wWKE6d6FWd/5cm3ZLJVFCYi14xzmzuMTrEFt3Wa9xJ3Ij0hsp7J+
Cb5MwM8zNJFlUpNQNpAKhjx9NudKmkmTFmxgD2zHLp0mW1ifuzw1pNWdNKbd
fJVU9+xf9ntULtKy5uDOqkp1jSkjX2YEgmUDae42Ibt85YCaV8iid9Y/dvJL
4X0nAtFE9aKsaGY5yw2vMFH9d2S8CfKq0W3ll849FDJ9YLPRvu0K54lBdGgH
4IwGQPqPdBNbHOc9IaTjrAruYcQAXPCft4MLRKnKJT4EpefGzEO+nf96S1On
YfuhIBewUkcHwVdKsbKEKdJS1Z+9ACGhS9N4aW0lhUUvdSl5GUQFfcQw5Mjm
/HHJ0PRMsbm4XF4g9pj9uV4dxHGIyEyrvFeCrOGrgZmtGjXfmy2V5gJ0VWAG
/OIAQ6fj7KHu6YI7at7M74n2uoNAN+ozMwdm796acmcsbm3LVS9gQo3EVVrf
Njb2qqSj3xrdhmc79T7n/7nYkqX1R531BwtCX5evLNsxW8fo4mrG13W57X/9
Qjli/UDoQYxrElN1I8lwhvLBK3aPSM7njRFCw2z9k2IPqqHSjyEmxWyY9HvR
A1JWarv1dBTLz60CNSs1c07vfWQFmWOvXTRJzD3qjgij254fVVwYp8Qw7EwN
anpqmcvv6zlel2xBpH97LfgGB7hJLQ24CjNwQtGegWGnn4s7+LyTnQFkqv3x
ws231vBIcmaNgwotVGqeef5N4GmCX1vr3Sp4egecv9BZ0IYKmqYoH7yO9sIn
hKC2/tQ+eP3QmSjrAYzaFWQoSNhyzj63bDfIMc8LaZs64qnJZ78bdGB6vrmX
RNCfwY1BZEBe66cdCEr3VG/8g7M+Ycx1L7F19H/s7ohqZH7uV0QAtd8AwRJH
gfghZPZrHf4995bgKfLI7diTmjNI8iYAO1EViL2atw/Zw0HuPa96mIpADapS
kEcxV8+NZ14eHO7dS0P8xyl31Z3t1KBhnxRAkVILPbQpiu0ijxCO+ZNMZGme
HcG3Rwo6Ah9q7TpKyk15Yl1IgUb1sa4+NDkpXfvhhzLJ6wDXEBoU1yrGbzwo
i/xJu576g1pAjGlXqW3w+iBRq2IFhUqyZTlSDgyqtp1ro4r4VmEc1s1dH6GM
TcPlIJqInddgFdMInHhXqAwKxGyiPKSaqUBiYnqpHmDQid71ROq2j7KjfBFU
5yHliE4iuOft8RBg8ToPhEk/TzRfh/npwQNVrd4rh8gXvOYFak5iNT99GaXb
21JVFXqsVIZ43fCaw/gRgOy6M9so5t/wP9NO83AmVDT8xvoO/HXm1gx22G8y
b6OXuXKTvXyz/IGxxT8Bu6uFy34WWquqHA/geggeDVlEwthBHK8MrTSuJ0fq
fSrKPJQLAZOlyIz1yD/DyewFDF8HyMFz5VFJkPZprCtFOYxAX5C5BipCq5eo
xDZERkxPVObAy/qHgefvWv9TFuQNkilzP2pN48Um20PgyR2KPzjjp8vR/yGN
LSOPl+7qb/xIshSo4C9oqg5WNSzUAjkPjgaUUHjIEpXKKvBlQrwx9RRbzIdc
/chUF3JmJxeV3K/4kT6/1Jmn7fwdlz4uFcBzKusGF+/heqv3bjO1pXEwF0eY
wvyL8xnA8AyXmlW3WNv2sgTkvDgNaCdL25cOrspNxsuj/TFZmMmwSrcPh2qA
MY+EyvalnmOStS3zEnRwkjG1MUv7lQFtboWYyIktM2ZXshX3zx8MblYN1uFm
27aPz+fsT5cCqIEBQ2x38lNWGgaYIawntTdUYlGFStOo6/2H6d3vuYOeK9CB
ZKB6Ob/pryjzYxPKChy1NATUtEXDLfasl7NOHPQ8Ylo3xRXi4T5hP0TnnW2l
wYSQEJFV8o1iVxeGM6gjMd2eFvo03iL9V0y1iwJMMbwA7ATw9e6S6n/cxbDz
atXCuyfEx2qrQKY/tFIDTvG6AQkzyqvxZMPGl7h8Q6yf2xMfWjZt3yWs+M5d
t/CzLO0bBpfBDGX6gU5uzmDMeNEY+3BJ2YBHtIcY1ND6YdJ403S7ZFrTYdTR
DAk8jJl42sHCus11p1eViqGEyB2dqClIDCl86V6IcuA3AJafS+lG1WpLlYNv
963mG7L97cyTUWmvt/4Wwn+xD85r+9zZNH32umLDvtwtmXgdXRqknlgOAnv9
BfTe/8hoHdj1E31cnAi5TL6FZbWDgmHA3Y/tyV5Jk/Gyqmaznn2m5UodtvGU
F3EPPfi2fZtiComDkbjIv1/cvsA9DMQ+P9htK3DcEmhNU7a8TwkomLy66+9G
gWruZ/9NAuL0Fkrig/OSaGhLgiqwjYFBGVkwZBQuCj9mBEaOs+6Z9W9oksgO
FEE3nm2IJ4bqjakHqPPozMl+B+PIN6x5xGs3JGufFFzffektBDDtKqSje6zv
8ozVWEJG7smEfrMm8E8hTMcp3h1IDMBoqRLsLh53WWqy6Ij2hA/nA8S9qfiH
1dU0znYAezZZGXD/1koufkWe7Lj3yWLCtEVBs8hvMUtD63Lu/Ayw8XQvJus7
T1nCTyoNUAnpARdveG1utUy5A7uIJTvpFs7Gw3n87MI4LvM0VEsOYKD+BaY7
eUjlQFrJwi/7ojT13lGcger2ETnW1wCq2KfLfKjS1ayrhMU7Hur10OOFoLYE
WJurK2pbQzvQij7+/GJnProIaZstfE+96KZTjMlH+tReRTp71SLTvHapX53t
cw4wQdi3NI+a5jDcL5J3V0w0vUrU2n4988/8Qk96+S1veIsiLYzB2z3TIwY/
vMrjSL7LuIUK9Od24oh2dhqSsRXLGwkEefWrojqiNnZ1mLfAkUnlF8i0xlNs
gKVo04oLKXq4Y5KAMiF7H/iOc7bMm+Z8vGIOu1Jc+C7G4UJiLXDAJkLPsrfx
CMPsLZ8ujD5yUx3kBO4LpvEmTlnhxlyqLwYMzsM2prbOzY5CiB/KBcQlk7DB
8mgfO8p6feU0rsWpHNZeAEcMvC90ds3t0x+FSeiVmPb+jSPHk8GoElUAMear
nW41Vbg18Cm+V2ake+t8RuBGZMdF/cT5eQRv/0htZKt2fVecQ4UBHm3Nfqpq
CcT5AxmADb+E2xD9T0ev2iuk1vl8IUJAsJESS0dpVo6+MFeBxRt1uqon/bFk
OYAevkY8Ad/ppFSck58c+QireRNhJxC7RJBaFZgitU3GERifuWH1ctWWZBer
/r0peByz4UTg29uP8/HSR1+gHGohkcv4gS2H5bdpnIaeS+i4YfixpyNEPGHs
Or+IfjB9wapFHccv0MIm88hxdc9whwwKhFXaB+3G6EetI4IlPDENBzsmYkQI
5VMzOMEl7frvdY+SIlapa/5G9G8u5nsRLpJ6wvL5kfppyR4FCcjEwRG8/91g
c0kHCyEUaQa4UjSgmhbt2jrYgZl4fc9X/EsRijqhBOzQjl2mWuAAD6Ghw71K
QdG7tqUNf5ZqNS8QbPNSOO0QB/Ck/uDKxG8W8F3gC6QoC8ZS9PGh32ssipb6
SFsAsC0UoJGlUYuh6RBla8Yz85PYMU6PjqN/HFhzSVfxe5vhjOfIH2vi3KMx
o9SxeEvD51r5BdxCMTlpp5kLg33Ga9ZrUExeq7vgW0k7ZKTFZnzPkctTDa1T
u1weXNncWjllvCQ14f1nUJLL8wzXAcdvaU+2Xb9KhbBY1rcNcC1O24OJiW1I
x6WOgJIuQHfZR23uxxdgwpgYYp8wkbZNPABsJL+Pv6tAD82nuc5Dob9WWnFN
n8vi4hZC1/1FtZkMNWAGcZTcvuU0JkDOaaL+ZTeg5/ImelA63Cey9G+awZq9
tHNf5tqqoFpFfLAWrHvbczAsgXi/SZNnVQoO5+w7OSu/5ofendZxSWs8pnhp
hFyZXX+ejpQ3iNWYLrXZ7S6wZVH4C1vt8/Kv7c17xDxPAtxVDqBTJvTPrTrj
7+3TJAHBR4ovMH2bH1mp2j92aOJxx9oH8pt3WNvfHQaW4kv3M4D6NMS2wNAb
W8ZicHaQtpCb8MA+KW1qPRGDNlpr0III6tf5NqVxqYOI99BTouglLK77iKiN
rRnXTD1Go2Ixo7BrS+EevPtISv2QSboE3LwbaKFg0TF4MUldHToCJmcILPPP
Zz3DRVAkzY6f78m8z4kXMi4LBU9Tu/YFsi7Ko3IO2nkpYOBP/6wgmiVvS1uy
EhDoKn/QtHm3yASwDZqkAY6RWUpkbxjNWsFTN3ho1EFcElPHbfDembyFpdNH
PePUzQfQYRVaTfnKcGqkCQRTQx+i9hb/Q8HmN4vmrgCO10XRhiRM8JSNivBw
L887MlcjznoGwjZ6TAx3NBfoqKbg3XnmIdgEovDMiUdsZkz0VOX+Y+wSCvJ5
Er9JJDTY1ZDi6ZFBN3io9aVsCZzn5oMtCOdkjOtF92rIVFFbbWGk1yCOYnLD
oKOXE/xyEiIHvCtq8Zc0GoIpZQnYn2SOjk8XTPnMiPjUkGYe7nVKL1RC9jJ3
cRHzH5BGJrrye16Qj1Sm3gin81jTenHnur9GUQt6WzKVggzRn40qfmkoBzYq
c4jR+B8Vfx2lewtEglzn/i+yCNhBSrMmCp2NQDo+wp8C9gWFeLyNw99//cEl
76j4gb08EyQl6SnbYny8Y7KPiy9hhHnwK20t/E+HxFNKxUhgwJijiK73BTJR
z7vXtaesi7Sc6WCUl7YG2GiZRRvE0QeV/LukLoe7IJl/5M/Fupj5gOFDgguI
ncZlCt1SAaSK7NCCJ4ev1GKhSQoLGnrKveznsEGHaVO134wQCj+WwOH8hcfG
+mmnXr9QM+1QfZBoOFRKtZnEZ8Sgxcw4JtgZvWFi0ob7jnUt9qTHpVmSwYry
la13TxGcojE4kEIYlbLiGGRLQlCrLMAtpgIETSeL3Xa4kCKR/s7d/Osq8QFj
6CY7EjnGgXfoeB6jC78XsPF3N21obJGML9k7IU2LeMPXs3XbXSdIkXYWMnEW
6GWrw+UOL2YxGyO+zFCYYLRGsrUT8ImHQE890+y9pzer7J0zJUxVJJUulqfm
TZCETggqj7q+oR2ja/VKbbucVSrEFKmPf92QkKNDj6lyXclTJydUtUYLTKbG
jidPhwVpKJJDEHhV2sD7uZg0R6HEYOytdOgXlwT1Qj0Xc6mL8Qk2bDN3uHeh
U2+NQklXPLga3m5ICIZ2/fORESrgbS4vqGWmt9GAxNsdSvntf2Hs+nFQJBGk
kTgPGYa/1076nyzfAONz1y36B9nUJP7165/vB4LJilEsyPRl4abU3bnq8gbQ
e+5gFSpQfJWhcCRBeZplA8y/bNji7qWlZaqcxZ7pfN7YjDtRmJ56p+fCAj5Z
ke8GR2dBI+qtPylKqT/MEXwswQPc2FTYs2Col2WdcT52hqbxGZShFWbLHYcv
FjWx7MpuhFCQFymKH04iDO+I3SbyDqHSuY65K3P7TGFS83I/g5/+7I7Nd7W+
Wx0kaPq++Y4Jjwnv0b4HMcx55tC46lXNeNIw2+dDd6BqPyN197Dcnkq6jrM2
XKSlLtz8yMqW2Da03RdUiN0fiZloBB+0dorAU4ESPvMG9IXWs2QMEvU/3g3Q
V4s9dBH6Mlo4BJrosXGhf7Mi9thDLBC3H+RtJEpoIopdUeMHgjJmNJxxfXlU
bc08vGwoWGxwuKXyEiXEbpMg/mPx/YLWkykozyluD8J1np0nuzquRBxqmn1A
B9mUnmjm7nrFYbPg0mgtF0uXJJxO7EwsCTgBhaC/77Y1ft7Z57qmn1qLhkxn
dl94gyb2SNZuDkqC44BAqUcKo5qz5tslh5C+dTNBPVbnOJQIEsOv9namaOpT
Exm/NQa3qlpUlJ6LzlyXM+9EXcLWMTVXgFDV0jO93qsqF2q9PNHcXQDezKNb
i634sCAkykyLE/sOFBKl1gWlYdU1Xk8uq0f04yUlmnRqJlHdid5AaHeoZfMM
UjuvITGSHTiK4TztFVwWqO51Swke/bul6IQnWN7wOzyOeymPqinZ/BfVRxNK
qLQCVgZ5gVCGX/g10VpKh2T3b+uAQWNvKqWXf9WQt87cJsqgppWgCZW+DLJm
sDckRjmdsFBsriL0QZOk7VJa2gDNdAL7ZfLiQxqEVBDu2kGPyXsUWAcfr+6r
RKdm0ytvVflACYhGkDqlp0jqA41+P8P19WPbwoA7ajTlf86EXSGECZZPfB34
N6Fb8nIOnouBlTYY+vkJxBfOk04SZ82Zlsk5QnLefzGJBsCGpRps7keyElW8
EVCGUNyWzVlvfTRm0itvYWGYL9KXtvJFBkU3fzJvnrNm4b2ElAwbs8YA0hzi
k/WEgJBJcD34J1L4CPnJgF4yi+eflUZeWDqSRNplJswc6qdRlMy7yz+FOZEm
9oAtQbVR2m7BPPKDd3j+iAkb2bEsJwZ9R25ztSTa3nHvOJ32e2L7lD/rpcXF
sjHUVtC5u16bvPRZ9YYv5yQHr/oTMLVzTVHomf+XEjB8NX/5QBrMm/bt8lbK
y3F0KBpFcQZB8b4mhpiccqcq1D40HTglMHUhScfVhGjDs6om2S4boNVu8NOP
JEF061QkhZd56qmoqz2U0qTyHgDQp1QxW2u3N1lIorU6g/tPb0a3sNsLa4GQ
6UESOydpD3AgF/P4nExVkNsz78O5hQbexBZtP4KDxkDgg0ZM33oijD/N/Ukv
HL6wmAqjP7UVsUZGZGH54UBIrgvNVt6VrhTo323l9kJhYgvU/C+VDBHFGO8f
14nY0N/sPbli6beYTHq4xEP/nCgECaN7KAIsKMYoW56C6LE4r/2GIUZljF6o
UvOcEYwXPWFcioSEco7fse35mcz2CY7DW5ac4QmkQCt0Y/kGnu3J3Gl5ffXI
LEKqXLoEP3BRQWdaEop9BpwFq7TbihiUgx+i2G5I0JJJVEkl5lwWxHN7c9Xq
4zjXPAnmWg2V73eTjUGggKtI0Xi1qbD+Udtso4KV0NYu6v2rO5bMXK+XLx2J
T3v6MpkQ2xWlEZd0d3wsMjN9rdSSs9M7/RDLsC7V+Sjxg8h0NNM2yqWNS5vD
c+D9+H7m0LNLcTR9+DyDKIUb7M96To1I5rrgUF2OpHxCFzCDjvcQfy8Gqq9A
XXFFPlGCKSYrXr+xeDfE9l8x4EkQouhp0lKBtjytO4bHG8RZIlm6In5+gxig
Iv6dzc0o6tt2PRH6exknacNgeTGeSacOqenA6cNBlBwru026x/Af1WXrSvCf
AGS89tUVhYyRHKoVwHj58lhwx4EM3wpRXHDk0d4JdPXBt/g/kSAFNycjl7Rw
aKetF6RCwQZlnHCBGydTAc1MjCKUAa+aZs0cs3GLkykv8v6MCmeyBJkcdg8W
kFmg3e5ENelrXF8reCAKZepx0AgXxuOTVV0fWj3JRAHGlJNDLEGhyO1p5L5A
a8HSaDXPFQjZ7YKBbza3yn1m3CgoTFM/A52mIJXYE4lu4LFlyyU/0sXA0GMu
wRhQ3FPpSaaAxIRO5TbrNa6KrAsAo9wYB5H3o+snzJ/mtg6k9Yd9XZ+bMZKY
kYVYJC7KF0vaoMXQGMhwjsSPCbh9SJR1JVQBONUT9MHkyxuzEET27qfVuy+K
pKh5Nb6vWi8AVu7gCx9xIEU0L52jI7Nm7ScZeRI38PhvFlukA3HRSHTgavH3
FZQodYa/BZDDVzeHmnc0CNbyVDwnTEDO6+71RqG5e1qv2z8gA7C7Z7sYOftK
uupkKY4/4ReF8DapJR+3VW9rzV9b5xMbuvxIHrftgM6yrpmE0HnF3BBhYvBy
b9K0AOI1nsUnq3L6FkiiWSh5+dg6KzJdBGO62dV5e3ArrPnvdEXkepYpv4Pi
TyGACSGe6wYSaabknBb+uPtKscF42eY32G86Mev1EcriDk29LQ68bNXkixbA
8x+z2VUn0IouUtUNjGU1RbgCvIrrHvn4RHqhqQLP/mdlL2XlV4L0g+csKjj3
c8Tnc/IEAnsMEHiKjJenK/gzYgg3dKRskUvQpbPVAqgC0Tre8UZeEEXixqFB
A1VIF6+60MESCImqaCkiPBHVryb4pdgu8yHi1FqH6STiU3Bo6azQfFG7E02N
+vzDdcrM+GkVrY6k+IfCLoozmO0f26+rLFvs72Tz630YrOVbHzatR4XqIekY
zy94W2A3I6/zGPXhGZsHK+UgtACuMcadWpkq1Fp+XuZxVecvAGpqyuy/ylrC
cFPb8brnx/CdjXzso8O6Ik0/r+s9jS77IfMWETYGbMhlyrUEuDgzubv4ppj2
J53ZDekGuh3rPp4+08M9adtZXM6mKTA09/tASkXER6Z9sZuGHdJe4U41XRu3
+vW5F7qgPUg089qcspxsv6bs8y5tuE8dy/u1Fc2SjOVGzvAMIiMeTzAmihjG
tjfzL5vZaoXehTd5T0YDLUp47E5FGUYqNZ8v9uAFfoExLZ23ORZB8e1iycVR
LqAbxdjI2RzNUIr/ipV6hPmJ/QE9jFsolOqoDXsqTzN3KM9esiB4oFNLVTDP
GZ1wohalq21Ea3Ge3QS/l+43V340fPtnjzJ/dyl/UdtjLpI9lqjPbcQ+r0JB
ZTi7udwbI7llkeO1uvjLKtSVeM9Y8PcljPohRAAsVe4YIeFYQj43viZP4kt2
/vj6p6CXMh4qWRvKnQPTydHV/kI0ciM9cg1u+UJJFLyAkO4cMLwkYzlj7aO6
EU7N+I/dYGlG2u7JgkYB3pZFoPNb5SYaYO9dUlnz/pZwOMQPlceToGqsgHvp
kESmBQiZv/MUKZxlgPudMqsSQHrbT3LhesX4iEzJs8JPBvXvjdp3IIPT85Xh
houVWbeHv6VyfYwkH8yHHaEqeYNJz3drjVCS4DKlb0hO+JTag4C+FL1tjV6l
aQTOw+fs3fLGfCA6t7822w28P88N8UXh9NS4gvaXNcjsR+E9CnHMY+nSqj1A
zkxQtUaS021zhAVWr9W9NHBIHA4Jkj6MyRpqdpx6e6mvcAitgvcnfWbSTlDF
Ss03qMx+QqZEwlvcnvaCMcR34WbEbNX9hqd/wcrT+KGmJ/Iiy37Z7TJ8kWsw
yEgk8M3qAPwOncGcEMJ/AH/gZ0aqDdCLcvDt7+f2aAwUDlxDoSBxO4/OH9wO
j2QXmSwVUkRnbRWcUIbGx1I34HObeQcjeq1e+YqL7f/WQ/IOpCyiaFMcp+L1
F3HvJW7gHzdyPq752sYJfNBbsAA4JNPgjgJUlZ6q3+rw68ti5xd+39HLcrOx
JZ9tUlFVBrvsHY0KLM6PwgRpjMRJD0feS5ujnA6CrrckDFQhCqhB2jgCd7Lk
IuZuim1umzyLCmJVbHYrT9eg9wVId42vo3W7PaA1fhcBiQRbB+Q2FuTE3NVp
ziOLa5Ha2E9Uqva4vSGd9V2jNTAwim9298UrICCx1uL7YS9KHeLkFswUweSj
0/Dvc5Ba/zxXQkBCDotkc4s7vPDKedAIsn94buEpUHRk1KtLycKtZcQMxcAt
JBXH3dGQjITJqJpQhQJrqPocgi7az8geBOzDWM2zBliJjNPM2LngM63e+swm
yKSg+BizHHpOlateUNtv8fFg9sQfZQlV5aVOOsbUH1KG2w7brvFwlofnA8if
A3sXTI0zNOvTBVCq96Y8+3lV/LG260GSz8/3KWsRtGz7adapiHIW9NQ6iTCA
iAc8KSLWk7/MV7atohU8XnHbDHHzR29PTROTVZ9Iu+e5rzPGN1ijlna6ct6u
cFnwwCz4rRTXeFku/lIqmxx/4xA5RfsnhJBifNBp7AZJ5zLNFYpM5lKIbORV
xXVd4qDH3fD5PPkUTswkNbHnSVtG5BpYrEzgr3HhkSUliuYxSNe95jnHIn/Y
3FHPh+abB4Z5wsY32wROOtcijYG/4SgO4B45hHaUNQhK0i5OCxL6xk7cFkmO
cmETrkvJUPL4UNurRSOR2X4YNyNaAiToN4cHQvAsBpC0Wm6l/k4+gXVJLLUc
3kNZ0aBDm7LPH3rurMr2Nwstkz4eYmMXc5n4ToBvhLZL7f2+a4cyjo1keRe5
D2FxHDiY0aTKe8W4JbAuyegRzavDgomQl3n23Hcqt4VN0+m3PuGU5mdrrT4K
nWm3JTYC5izoDrQCLLqm1YW3yPnMB3v0xEil1ui+SuvKkDpO+4O3IwtfeJQ+
3gVxQ/XKAmGHzd9Aj6/dBWWZ04Hy/YTOXmB2egtAGS2SJCEJIf2A28qLXrTt
AWQvja2PXCYewFV48OsLbb0CWxx9cZTLSVvNr7qfQaDbk8kHOQCx+pzVmLmY
hTPGVXyaPaVKSCZgYjtyRKvh+t66dTNlS7eJU3XFFErjneMEx5tnUTy4iqLu
IAqdtpcbPu9xOsepVBV0PrE3E5Jr7hg0aV/OPNbr+OlNsPM3+iOcAKpAITAy
UDtTOkQvF0pL5qVATwcN2qMFXZW4EiZTpilfXvA1gFTXDEBqEEJxAFZMRx2q
zzWZox+5lyW1UbMlTsodH2Txy8T8xEimuk2F6ADboT3RyERObBXYCa9FtzQy
X4MiymXJtYVpceeVRl+MFtd0Y2A9a8wGizcy5300IGV7nNv18Zkv6ip//i2K
4gop9JdN8VKgUnQSiPrPqsamgCd2oB1KRuyiFZUqUD/hQBw0ZnJxRnrOBDNs
c2FYfC9SsgZAsK8//4M4KiJ4q34/DgRg+ppbr+XV85PnIuCDLvFy9R8n/NS/
4TG6esrS4FeobKw2qgEhOtt9U7hBMczL2R35y4vv+WeDP9Q79S0v+2rcPQaz
IkjBqhuaJot7zZal6hkc2Z2OGeWSGBejSe2Q8/kik51l/TfQ0fBnFmfDOBiO
yosP2/rT9PpqSFBH7brqMY1HLnPXF9dcrvA7HB75QXklpgQ2ZifImXSwSxw8
jk3ET4ACD+rGJn4Ux4BFPENw09ffxLr+p2VFEI+Inw6EWWm2z/DN7Vb0+xxv
L8J1gVfFVTDWDR5dNJRgQ5+QyV4b1+SgcVfWN2h77vOxcf+iXjg+myRnivDY
n9AFg0QS9KX+M3QlQDaiHmdsvX3mGyfwwk2659RZUWCfBfoY0qGMeRK6n40g
NnnoCCWyNyRB1cTeiMwzb3qXQEcOSoQvmcF0j9mrP2XxfrpY+lT+8XnsuJ3X
Ljem9yq00Cp4gdiuQcJA80zeYDFAE0mvd9HT8OufwVJPUau3jTniqsF3lCC1
bRtD8nlALj356+XtavDJ8PpFmpRbCebnFpQKZnK2QBg6QEZDhp8nOjDgJ5wN
8ZvSRVq5sHgjV8yYZhPRundjlUggEaa1gq+8Nt8cWmPCuRGc1WY5fcOg7J6P
8Xr/1WRbK8jlGjxl9M/hs2Iuqqcjq8+jo0Fwr98Zz021NCW3C8lN7liayr8g
YoE8XZrEWXxullXUs0Cp7Dj71Xf4gzQDkHWhRnQrk/cK2zqqdfkAxwJTbl1n
CjvJZGxxfZRF2VRNVmtxDyVHyOBmbUqucDurFSkikeJgpvAr1HNsFdG9tqdm
5PiNY2VeZtGVS9VQknuC+VjeKIU6M62kZp23JcOVcfTI8s/tQuUhAjRkZyh3
yyAJ/CiDN/9OZyeLvN89fV9YrtOCd9EV9ricUyUxMNEHtfoUUT3uDgRNwgFx
VuWs4+rSh5AMKhOybLlcBMLxfTCQm8e7gxxjd0wUmXRyHgyUYJsSVT9rlTxD
kge8PP+wH0e8d1P8X/fqAvrTQZv0ubr/6P6JWvIOLsCZR9akoZhBBGamjNUU
zZ1iF+erwgUdT6DSXw1POj1XDqDyG/EYBjsTprPLEbnDMT7FuHKgeYlqKK4B
FSkhkXRKNp+K6q7qNetFhFJsekaPesgbaWkv8qvJNzi6KXFiWivjv8iodq4M
DM7PD7OX1+ZyH8QhDBnY/YEcrsNWm4hC8w7KRjXq3Rmt26YlYxVOhmZS1l6r
SSHLrasH1rvVCzLNWE9KVEUrr3TJ6BokDE01SoUrgXj5rSAw9WgMJcy9or9u
JxJ4BFTM0SZ2K6Nt0ROu2LxFkw7UTre0auw9ClH5N2gjTDW41qAU4cVHgzw5
xAEWc1OhdJm0dWQEnJlClLIrvLIGeaJOoKKU/9RzXs9YVeVruhwpjkTyDwv2
Jxmk7kVYPHBTdNb0IpCkRNzl2rugyViefR950LnGv6BC+6Bhx8xjGnj9qM4t
9MqU2OSCktDk+OPQ3egE9rWnXgxA08S3DTXuC6DGVFe+JRhhbF/yRED/qHvF
s9WlCAv5kEh91oAZDByOr1cCLTL5C7KGh/RX0Qot7QZL5xOcoAQF92rbD14H
bYTDigT37UDjFhJLTWlXDanBMTyz5GSm0/pqERvrMxUNlPuBlvKfOAfuuvZn
3eqyBat+nsRb4wm0g3b0eiqOrQp/LUlqB2wsWQwxAnaKg7j88HVjeeP2ezTV
bLFe+YP3JfmoyEj/Nz5YI8PIxeZA4q6XSVPmCKquEeVDgSCSl/69IcfTs3/Q
WLDTGpQeAmPqv+QKVJ2Cqkd2AUxgN6ge5Ge+mPv3wN7GDDJsEubd0Snxx1TG
kuaDLnAOR/Qom48tDAc0BOoRBlfLmKfbjk9F5BkS8qnV1QRiHa7x0FFPQlAA
UM6CpgC9CaKk8DivmbsO07KHj1prW5JCzNli2hrz6HTEYr3uttApkC+YFhn2
uCtbVotfMrCsplwyY8T9Y4IEiCrXqjm8A8So17YhsyjWc7N187qCGSnzbZOE
tC7vAaKPXEO4og7YsKNYV2/N6Tp3ExuZVm7gycKMYLfVbLjfaI7hDK5Cu09x
p6eB46Z8KF9I7LoMwV5nzZqxPWeAj6e4MHOyS4fBFe8zyh1GHm1Q1z4tRLGq
LbxDGcDjIHiIKxRlDeRJAvvGhLVrfA5C+oc0CTkE+S6nTLtC4t7PWdcQyV9N
ZScg6aQiBpjG1OQuv9FiLg5tBjoeCMqaNYdGpzBHQq4QJXTFN2VfNl7XO4tS
F6kxS8cVX9AA2xK9NwiGO2ZAAEeJ2/lgwxTCyyoWUWpp/qSulZpxJB8Ia0tn
Rk0cqZQf0ErHmSob75oirT8UtxzmtsTWtjf3aWazloMnzitZ0+s1gMmPnj3R
mcmmifZtEbdMWt5xwd1l33k2T7E1cSCzK8C5W1NzGWftIz3adXxMH0czrWao
z+aZseE8xSIEkpg8E2M/pcj+hjArgW0+hcp8fUUVZBHXc9IynrshwAxa4gMH
mfCh16mRPEtH5IVtgmCKXOTFeZzxQmyxL1OuUImRKqPm6BcN8lEXrDudqToF
l3hpGnlTSiJhYbO814i45hJ2dq+SQfof3Y6dLdXKPB0fQXX8woKHWuWHj+Mp
ZKpzUoVec8242Ncu9H03Y+7hz2OZGbxX76Xo4k005DDALrC/syQxmTRB8THm
kXrZQxjw7q33ebNQZLuirvR+L95K1eS/1QqQyvu9NxN8gDdqSItHqawelroD
iBsdsgYCrBq2gO697kwWve8MJu89OlmyJYTp9g1TFn3OlSJEu99SyAS9mggB
tSLThCWMHVfoYjzXbXONyL3CdOc81luIyvVtguSRB0tZ2HYT706RiGY/RD1E
EU6nRiZ+rO9HprLzzJEXv106T9HrOgJ1dyHXYcFOSNILpeHnHNPMQwb9S3BA
4mP9qwg7lg/DynXIW7x3OJR6FX1ekocQsZ6jfl7wRBVcTqvCqsVuDWHdjWiA
BRMcRjxkP1jefTRyyLyTNe31OzzFhP2OM6DPhj5rk6oDHDxxF8ccuM/R2Mc3
PIjsj9hOQRZcSGRUhTbUgmAtam0IUm17t+jsPAxq1LO1e+AaaZ/yxjBPX7yo
q0JTwdG98lP2WWvIMakRerkRJzYCPxPQH48g3qDiyArxA2ipR717x03+4neI
NYMY+UR4JbjzDiCPw2TYRkivkIscqVmDliA5tkb08A/fT5FVWAZlsmN4LP0K
rvDY39qlkv03xTFYqHNbZB1v+iO34HMWXA/yDtlhdvjJn0l7ubjLySuct/2l
xgxIrraGEfQ6VEqNcHXKBV0FIcXfd9l2ec8rEfy3XBnmVndw4DyuwQ8/in/d
s6wz06fAL3HBgk06K57cSIwLtFB1se9c112Q+IG1R4fxX8O/45aM7IiPzzqC
8+nrSLUiUQnKR8aBNb8Uq356zM69TnK2c9gp+WIBHgf67E/F7MQTbHSWoYqA
IGWUsUvmRjUDsU9qtMndboZE5W1/WP60BckhGeNSS5XunPbLAkVQGpWZzpHp
Bz7WXVornRrDBWu93sfpFbR8UVD8vxUhq507DRycCeBOtK/me8RNvH/OLZpb
5SLMQPY2O9fQl3uzv+cAq5+f8tlPouaZ6tlnzgGb8GbHL8gEdxzns2E8UrRA
fkRbzf/wGtRpbbYs4ji7RXcbIRahcMz2d+RQHrZKkz1rZxLrso/9rsseGwNk
/uSIqDVD/EpgAPgT3RjgKT5W2ney/W4sW9wjqwf8CgCPIbPWOucTdg/x9zTa
L8reWwV8J2AEZMqFybuVfUDMpnHPQSftAfDSjWVPZlhmEEpKszkyaBsXiuZo
Ss7wRSaWEJeaST3TrSUqLEVydB80flMsp8MVmmMB6P8h4XvCMlrmAJLQeYDZ
q2MYV39cKdS5iOau+mG93/mVZq5RSIwjs62jqDxbqvww4iqYWGr+iJ4tNUIh
a2GxjNgEyequjnN0jjiraeaNJLbFiZ9RV0+Sc9YcvOkvYYce0GxICuUiJmSj
ZfY/8AfHw03qc+qvR26nOaFWh2kRg4ThTT6cgZh7Fniip8NyMfLYfH2w3fQ5
nLhZ3oTwVrrjWK1redJE8Kpj9/bL5UnLJGJyhzovUHSry1Hw0G6e7vWpi1CK
RHSs1DTe0LtWWB2Sy52+jvZdVD7fS3i1v6gzRTOeMRUCHKnpuEQ8QtoHEU7f
tJ3Ucl/x34X0xYuVkKWnzTHzKymJ4dzAVLYm1vITUNAHGzKHuhD0aOppJGpH
p+miNJiHa7B68D7PbWxqxwHRK8uth82R3kmzmPXaLYEkM7NlR4jOwIELqlMx
9XwagLYwXy9d2Ap6t4XTkum/j3U/ROktfYkZSK1gEShQ+FPHl3cNDhV9iS7V
PkH2kGBA6mYrsjcbMrJ/BYMUEG41u9IZ8Pgu6vtA0qUy5GS0SPNgs+HKpEgg
H+5FfIcKuC36sDxDl/SMPSmK6G2mUyq/2A0kvaBWsxEzrkhCpeanP/jtjCUD
QePQVren3/IvWFW0bcX+ffak0AcByvlyvr0c/6w7cFeBgF839fnBSt0rcReC
T+henH8qusRSWgRodlmNMKkJ08cWmDWw96MJyTf3OP+plGy93HY6cC/I4l2J
cgQA4U07Qn9aJRfAvBD5YqwxkQJQgG0mvxVWXsMzXO8zPRwit77XERZDXHAm
O0u6+ann7K9Naq54mL0/Af3uimdUz1V09mBg4ncDoo8duXGoLlxp5CWqhBuw
m4rYOK0vesv1XEXORgCcWPYZufdYW2qUxJrq+OKXh5piKmJcau0npkuBhtHk
2ZzHD9QWdC94cfDAabclXIVSh0OVyskF25JZBE75uRJWVM9MhemG1v8cPBj8
9Z938YVVIdpqDFX4Io+RkU6ZIscr5KXn51usz1c9c/zKSAyjaQnhRJrtb9IK
Ps7Pk77IEfke2AVHJBxqYE8gi7lN1NECrJO7rh6coP0qa6CNPFQTDaUL0nF0
fYukZ/Q9KoTWzHYXDzCTi2mm5iE6LRALyHAaPo4AhGSrJcYLBWD8k4ne1vON
Gi6rVZThQ0MT9uXfZNH9G3WtAfdbouyExUIF46ZxoVNdlfB6DKUQ11AjpbGH
0Z8B2UbDY6ZQe7KSUOZNliuh/RqZPpJtBvwvLOqExgRQtZMuWpvZY214nF7j
NF0nlvpMJ5dV1d9YL/viy223Mj9+xnAbm+IcnT+qj/p66tPmtaH4XncMbN66
B1lVPDZyJrAJaywhzKZESBswXtCI9ASSp1T4KdLCx8VzJBVn4c8yPhSlSLfA
bil9Ib8/LtmjbmlyGxZDcUr7UdfdpJcOK/GsLVOSe6Z6WUSFIcKEDVcRhSvT
DZXe3ZNAqTPwEVthgqduYR4xhaOu/HvO7E3ZGQ+bo5/S1BLzvULGwOJjRz11
HbuuysZU9XW5N14/MkFm/tzQtN2VHuDXI6VlPYCPx1w+t6tr+sLkHNMeAlKK
BQO/GmK3oQz8olZU8jLLZqRMf1+5xi339CZCggsA0AJ0aCj0I22Sm1+QC1/f
3HVjy1Mh1UHNySEQkPrX7XGxH2VfVmZWapLzdvBkeVJOx1nrlo6Zh9ftXG6G
RT5TP52JR0yc9UKBORxlPpsWiVIgQuF7oJFDn8bsk7+TRguTD27NKxWXduSM
6Vq7SrOlwtMQMNaERXVx1H7aKR3AWYTThMRTD/aIFrylNy09t2LuJbGuQ4eD
1SjHwH+bsr93V3IAIZGFzgbbBNFPkgcPkzLXSU/aFc6xqFQVP/C6yIWq1rMS
cfJ9euxDBC/ho9e6XkAeKJgKzBdguTCdwwcu13VXwJSf1qHX01oyRXN6rl73
0Bejk31AFIEbKFguv9lwEInWc2EJRjyPebLKprsDBGJEmmAjQv0Tu5DxiLUc
eDib8OD9fYRt32Xr+k1VVe5GRTsYbArOcgwWwSpAoBU9UZAGKpPCuS0imOBr
Pnf7ZuchLcGCl7kHLQ5YhmR84dZHNG40qFgJAXgzYT6aVlKW02f09CtB1kIr
JYjlSPBKyfxt7PyVQGCBWVA0QiCJ7eWPW4hWkCRbycaa5A/pfddE2jEY7ZuV
aeEO3CO6huWqv80PXPB8h6fQBzduP9ZDF7gfs4yp+AP8zY5yqd0VutjC92XB
aGZB922xW11VHYZhcXnksm9Kv9mrsHVRnZU6cAbPfreQFZLq7Fs7nNYq0reh
wQaKcNUIXpIOWvNYLqOA51NurWNwjGiJ61DbUf61VzreZTopenyRFJ8V3XMb
GIXyxfu5RH52LAVoWfQ0zadZrvP4oT76K5q0lNzCC3dKiOLsb3Vv663zsGI6
4Sx9zV+Bft+/8E2WVfdb8smLM6AeL6thXwlbAKVKDtXXUQiQra67RcCbpQG+
9XR6zXleuBo/NVlNj/zqJyXCTadENSc025zvAAaC/4iRr8rZyNtbbNPzzvXr
fAFY+s656o9SNGBc1xMJ96Xic9gjKEsOZCRup8BAzQSOanWV5l798Owi2e7/
jRPsDSyREKdpC1IPYLHDKIyCWoEGk/JPevoAABXq0NkYgYWKmohPaxGgr4BJ
LpunQiNNrQStmNi0qkKrPVT4EZtq1wwh+W8eEcMvtJ4GEvzXPDp7re/NYOTJ
8Z0MJ7y620eJFUNeX0vhDwC1SssVY91BcYBiwaEa/IKs5QQjsfXLJAjInpFb
vEHKjnCbNTuHwvo3jH32rQs4MFmY0DYgD3arV0EvBcwwC16Q+yxs9Xr/6Qwb
k2aRXy5kW7SzHmUJ13dkQ95pDoccYdvOCVRLJ45U9PTmZecpeQL7PZA1UwVl
F+vDt4AtxpR1AHh5uw/j0o5SDrGQyPtvVPs6F0DpchHPHSO3RGrWzURSOG7r
ci34lVCLZesvmM7k+NRWRaWrVU9wT825iL3rWNKFHrd0Jw7mCM7wgpb1kec7
666eWdm/4QhJODtlis34AH/gLB3DP0Gbw5tVMlSeoklw7E2rKuO2fmLiFrb3
7KpQLu5/VnCK0mEiFHHHVez316cm9HBVZ3RnRztIjVEEUao/cOvDbXvnvoX5
TgqmiLY5BiSp1sXf34e0X02ef5Ek7/C7yAjjhlZQZm0JHXbZYRVe/SBynUDK
9dxUl4dLqCT8esVkzm/2QcQzBueLM9DUh46t756MxgwkMUD35n/k1Z5JNfUB
9ic08GjuI+NbmCmsXhbNRK35A9m1Q6HQx3bBm8BwK4eVTDzpvHWMutL9YQcY
E+CUS3i/ylF8l39avAaIfIuA0gD5JLAixyG9mF73uIQYg1L0pNirZt5QUeiz
RKDMHfc/YfTq2JIOTpDTbY8Km0u2yR0WCZjFeQ1DRomMi0TBTet4GgnY3Mp8
xK2iGV7szFL68p+RqweN8Yaz2VZcTKCS2ON1vWiWdi1KZZlXdsKeQNR8tEcN
1jiiYpaA2SSZdPk7As4yszQpjtope2gtdNpZBBh995tdDzWR3B+O11Nr7sOU
T4QDwGvNE8J9Vftr2u6zIOI4/oxo2RCiTFOYaSBgidzVq7xhs1CCM8n5G1T8
V2qXrEpy5DtGp94vbqrAyp8TOlAufd97P2J3Jbb+0pgSS+gpEyMkt5iVNIAO
TdQH5NBSfRygrrNFtA8JGVp+WXlrcEbr3SDMHEwcyd+OrbelNrKhUx+jKNWY
G0hjtAdJs/Z9DdN/Aa2MZVg6YjBvsexI5f2noOjosugu1LfV/wadqt4oIJs9
rBs4CAKvav72e0WRKh8qBvdecfuzQW92YiqqNo1duGY7CZ7X26D9KvDkarw2
hFk0+GybsClgmjZJMA236vA8UkgE/eCl8+I7UQrhuwT8p8rr2UInxGoaBWWx
0Z9Z1Tz6GHR+FzgolTnHkWPxmw3hVkewDF8+wcmoC+DNedtVMAIIJjVi37BJ
JEF2F4y+unwUBbh0tJCJ4MY6lPHgee9GZOd/icKmW9hUAWcO+aaj+HHLm0yz
aIPWhZo9vKuRg4kQMGo47Osl01oaQY99qXYRmYbMd2MnYau4x4pq4R7s7IA2
qXpxg296yg4w6YNE9DZFeeafqAKXqU/P2au14+tGs28l03ViZDPpztPQPRqp
I8JqR71DJICFqBavyTVfSsMIuILfb09rOLgGaeIeHJBla2QGq9+9gshNz8ow
GoUyEO4WYvaM1Il9nTkKpe/TRG20LUM1Va/Yf4YElXfDKoz3ntTQEd1amdj4
yF/4ue0rPLPzqIxMJ6dQdRW8e/+qFLfiskrupQf9pqf6/RayLbAZrGHfOvNa
4FznA5/hpfYgL23OHGSHqOh+8O6uAMMeZb7pwhvvBZtOJdit9X1AVXvosl4Y
YtZ0GcAtmRsMKkAeGMK+6qmU+gDaufQ/aOw0eVJ3zekgJRO83cvYvofCTZ9a
WEjSqJNlb1uTZpHaG6qpCKcsT93BL+3Nweatbq2CsKcBt26XvsqUKOaqlxvK
3iGcF0af+kHBJCg5aZlE5qbpauPn24bd4unV5U0jhox4XX0XRDpk3MElGpMk
krTX/QIjSPnP+7PhYdIHxDlCVcqhG1/cO4KoirF4wFUt445TCtuUOMOSR8R0
9SuJ65slRhB9MwH7QNroMabPr/wGMfjynSAqUa/CQdV1OAHpgB2you57mP2m
akIS4L6fE7HJlmzsLrVBsmFH+wqyMpRijXFldylrxNXDH2UE/jkplyzG9+yv
GdhEIKiEw6V10Ei6392w6CURv19xW/Bd3Az0zoTZyldOo/zzb+DepP/lNE5X
QETGemu49YpF8XIPxtZ37ClUP9oWRzAQj8fAhKEqdpAGDupYmd4R89lOIcvn
+kc2stdp5wT/Diqhr3l2yMCtI/erN8D4I/6DVDsENi0qmjoeh/4AMkN69gvp
LNK9xoS9dGOd8I62uOv1TbbH1WV4ChvYoCEDYZPjbyBQ1jzSYagWdlP0r2L5
fsL+CICWMF83C4shLShmFCjmmdXj1rJa3rftiu5ZQD3IIBlHcCmZPgAMO8Tw
sibuxEC6wfeKP9nqDolzHshwm+TEZvprlkBbkYINYOvBuDRGK93qhJrYVNip
pvEthKqQXDxns3646/9kVOFc1rbbnFKYIqcCtHHSMaW2ll9fe8xTbTmx6ik5
Xpgx8TT+awJ1c69flMsWqPd/whKCsDITeuzUJ98zr0SkVwg+g3mmSAfqArjd
PcllD5JmETMaUQr5RgjOkhTzG2L+lqxtkMshXvBOYozso8YEE1WiOe4mYOa7
mx90RpdfurZYAVLNmK6/jxMp6yw0RM2qtyAT5hexGb+mFnFJpK9aREHlSLMb
EnPJr2et8bNH3bzuWghKI/55JSBiXv6vMdAaRHoSGkrFWxrhlbzdLmimC7oE
HhtJ130KbK05qpH99/LWOhCxXkRLFNHt3NybcfbzucZenCypDviXh3ulm2S2
B8OVnjyX24ed7aLrGa4ZfffUF+mm8tg8ZFqP9/eVPst+XZnXJxj1ouWSAZZ7
eLndHlfozufrT3xUUWymM2o+gLQIZlOjrLUv3CIFSfQvPDXlxwgBHWSk0HXc
4F7B5cz8plqDsReZg3dksh8CONTV/AjEktJLukGMTgLZ1nLA37PdqI3Mtzt8
plBsBwM1NlmWvT9IjWFKHtHQXEuTTCqAXbvYGzcG4gaEzTZWhWoL0T2R0JJD
GJkmWhyrdicSDQdBHg11BCi06LLA5DXhaxQgu7MNMI6rH6oBdjOhG2B6bb/+
PuDWrRqM7SN5lKmIushRLztQ3QOMv/fSt8OSAqW4sEhzZR/U0d+Nd04zQshJ
BtVHbZz9pVGhHvYR4wNr5xvEGaXy4ZuFySePwlmI1L2UqjtNRbDN4gA0jYJE
Zhftj4cwmkjkWe0+Rp9y0izYNpkJ0oS3/kkN0wvwK3x1IZ6DkRCqSl5GwCr6
xlJwHNX6dhMRB0pFbxiOWN9rwmu04sbX3z+xf6s63xov8qT0KBX/X2Gi+Ruy
qaFkhD0huTEt/fYEnoY9lfFzLZVloca18D+8eJPDN/y1bC/ZmWg80VSW7GXZ
qx21zkQio3k+aEUvkGXRBGaUXLBttCPM0Ee0UUvFvxghHUfpj3hNlebCV4j+
wjowfUICJN2ZQn4K+vE49rcbduLOsv4fTCoeAJIF+9ojRvvcyfhqVHWpKQCE
j1titq5uOIxtUTzCZIiFajQ7JqfBAxwCtkdtDqDs8jzh0A7zRyO5bZTIm+Qi
RZIeEiGarukIXgZajfQULjhTxHAvk7kS58IbELLwlH5p9gb2Myi3GcuRfICC
9FfB8JqDXF4RmPV9Gfy3CfOdnEp7Ujme5w0ZN+DIMW67TQnx/c8Pm9If1a9t
NtIWp0FQx0hVMbzv0BpIqY/fVgdYoQgsiLcdUkWcmO6XPEsGm8XEfd0sMhU9
M7N/VvLgnUjlgwFVdOZlKYgpCLyDZ9AEVCzp2um/dzoUAi17S071m2b5y/nG
3V2Ma3u5ZVhIhTMbHaqTaGmzPzT61LDrlknJv90Q5DRdGb77548E42q49tNd
Bq8CzOqkOaDelZG2G7IeAmsYlxK02E2XDrZ6M6wyiXKQ+EZ/5DfVyVJCcudp
rCtxJbIpsN4+bWdW4gh+TrVvb3A1a+OMshwMnpksIVeBK8P9JXNTTujvnV/B
HZUF6Hgqw2XWCOvYsnWxu1pZw61pJUsnsot4om6lj2YSoLtQIA8dFeiy+hOr
W3tKuUQinBgwzgDC/AenqxwJK/bwUAc41k/l48mosRA/fA06Fg4tYSjifaUi
Rxhj16bvuzCe9lZo4Ydbl/1i4LbsMvlBcw+HqvodUhugfIW2wVm7H7VV+KFF
b6cm3TamohjeGTjJhK8TMtz7ABsGiFBHMnmI3R4yPi7zUAzISo1zyKK2/MGm
1UIwEzIZD1y2Mx1f7NDxnqsRNqzAEk/XpxJkenNcYaka4GHToon/dCY/6CD1
VhcAQnPxGk6G4ZS8EcuannNDAxhE1rwuoFwEU64WqkELXaaFmoTGfpxqqtCi
zkpCbkqQtk4E6+aP25cm2EiEp3e7drGRkcco8A5GUWZFesZf49U7fyRSoZx9
OnQQp+faOllHJ1tvWycBWMEDhy1J7dSi1nnl71jDsE4iMk09PePommC5yVXS
JcNpxPZAhYIucURNRp0UGeUoyCwKRG57V8C50JF/feA5YJEqAXsutRF3/zE6
MkOBPicqGujWvo2jodOdkbFBY5+VIbuhmjAKqbEQHUPrwIRWBCEcUOjotsdt
Mf4ixDBMp0lANtQTsIDSvnm7VsMNq2vKdkhl59yUiStSnmu4VhOUN25BfxH6
PfmnpiYHiR9oU/p/inOf0boS193l563086grQTpNk023ivXzKhN1VLzFv+36
joBEL23f3sBhHcyZK6CTBXwXutEeTmDsHMmrfBgcn6NL1tQiazkSwb/jj+FO
MqRTdVdNB8+uE9/tMI7hHEOJLuKMD4871gDUs47uF8Pw+DNLRj/HdHHMyqW5
qV7uRdo5okPjlp+rNLIuh3Y1zZWcmZ+RxhbtjUbaVioz9VSaD8fN82wlMirq
qAN7gFWgaMyV/w/WRnAg+NOi3ZhL4Y6cUs3mb/z3Q5JtpNahp5NE+khNlPaf
JnbqPmRkLjy25hKqXQDob2TovDHkUFMmKfwIe3P+4zdl+p/VTYG/frwnsYXz
oUeWeWe785cXO7Dm6yKyTd0Ku4SwwNJWkejs+PxsUGOhja6MT3h0ngiLxzEx
e9xdwJ2i21xG+e+3rnQujLSl6SY8UsG2XJoIExI/B+DnfliySEMZl5kF0sON
rC69DSPbqSFF1ccjJhE3M+7Si6+XOkTd6BEcG66rxDLiHtJ5XrRMXjPZJCPy
M4asciycHS3yqJT/Wgs8hDa5Kza2wGJK44O/OjWQzOxNNP2cLsMXCVJxMKc6
Te7GnAaukG3Om7kO+Bh+9yO5/G0E3Yh8lZg70CJRlRjBKhbdN10mwiHx6dE4
5xA919KOpDLle01aK+X6DQH8mdJ/EEX5tG1o/9Ub2ba8/ShbnFD5dMfIFjOu
gKN+p5/NIV3qHxQrx3WaXWfpYMxwISjRFkVHapsBUEgStJIu8KcghpDDnyf1
9EzwFOODgqabm1bkF9Qm5rp89cMLZM8IeCc0L4BADN3AH/bVt6vUgsLNhVs+
xFIAKpF5qz6h1Zgm13WjT27NlwqENFjOi2MjSzmMFpYqylv7SRcyZgt1oizv
pJqa+ZY4xDXSj9qy7Ts0nzXzwRgLPfsVp3Ld0NBVr/Tq5Ae/xKEA3nVkihDw
xl8JLekSbVi9nhvbM+idqoVJpYe1P+uv0+EyuC5e6Q+p3ThZJs3wYLqYYad0
ahN/wPyLKZAHDNDyeqDBuekl681Imzn45hyASBbSSRAs5XhlS7nDwXmsy5gn
vcEcE9EfjAaq7TmBF/HYXnGFcB9YiRsf6YuBK8F4denGbK3fprrky+vHS7xM
65ktrZmesUSrT8lekWBDuzsvxIOAsPNDUpPywwpEekc/yYqcMv8lcTvqykHo
XwDzctnf7s3RWgUrfFhoRYdr1P9hDewORVQftmzSqOIyCGTpfO1NmxOZYRHD
4BWcC3B0dXmLp/eeW9ZDaSeI9TLAjN8Zb8IcvagxO25l9GFz/ZSn8ol4xZtb
zW0hI0e9BDBGJ1yOlYbpiefUQ5QOPCeCM4mtaAVT0zGpddpAZmnmsihad6Cr
TsGJh09BjbV7I4AEpBACM6ZaPpE5Bd78i5o99GyhDwCVbCvgROwGm0Q8fzrO
zEkjdr8EjUZOlze+wZspZNKoRhwnb3mun5QOPm5oU1D2K+nsJeFsggQWWzhA
rMIhCd0/Yics3ZXWYz5ZWvIJZMtSbLn2paIVnGn9S8JNsUWdnOC/423oVD0I
aPdwK+6tS6wLDxA4isBZU99IxYrAoOF6HRh2PoBwSVnvSKrDaF5IASKFC+rs
AipVHpaOFZAU3PZLLr3tMOSSNo6lsa83uyjj0i4Cdum6o5/1Neny0J6W2tzg
XOxf6zjOOWNsbf5t0qfDAciKYFaEsWi6znZwNXRFMbuDqA5CPOzKy+ynL1Hz
wKWxhX2vMVQ9+a0dQU5wlsCCZIHk+JhkqR7RvZM+I36ZPMvHTvsamGGScqW3
nSonpdOMnSNpOscP0dftJa9cYySjuFIRZvylqA9xsndg88h96YBIALnRVkTo
zkdzgQchNmv42XzER0sGOGOUXcHbC5k6yT7aFSwA9hgimEKNz+V5/ADaWD/5
say8t4/FmxME3vBeXchszHo7OkrocLw9IPnNFX9CBAcVcmgrmjttTMvRKFpq
cYAp68W3hn1KgrsHHgtK+emDQesp0C/zpqPh8b85sP22lGqOudsDUnjQlMl8
WPRMyKcbbGod5TBQUQA4bNxCSUlreyHctH00WtrdOCSMEYp6zahIY/55rfVs
13WuLz5z5OtU0QpXe8xoF5HvfDqxOgr3Ly9MSxFZ9Y0NEVqGiNWESNw38Mll
yfK85E7zfTf+YCUOoQyuMqBhKl3ZQkVvr2ec4PskM5U0i7EeYvZ8q5UWc6z8
rIisjtQSc3Ts6nj1MZaFFE0xC+SkLO6bgzMltqgCpyoOIkQhIJZoTGfPliXk
Gi/YwxVgiWwKroasw+Zyp5y6VkvHB4C0no/194c9MTytFhV5SMhykb/cHC3j
fbmgQCq4pgj4p/lsu7/zdF8FI3CsZfH5lUqMPyMKHp5+b1KB0QOQ02IcG0jY
FJ76Ri2M02DcQbeiM92B5CRFuU91kjd9BLwZDnalWKFh6PE9o8+tH5w0Yylr
fl6Wc2uwnGPV96332h5cF1rXotpfz2yfEuI2pRdN3EoA1vQwetsdaosyIylh
pyRTvGJxbQeUq3TGkaFeeL5m7B8S5BW7+WkOsYqolfH5wGLGH44vPmZWL+j7
dYsp+OQUqhX3Q0W8FLuk7Z3avEIYFNOlnQQqR9KnvjT5NasQG6bzEFmONbak
gL4Ps6OgXaGUxi5gh7XfaGEoel6Mp/qTYRIb7uDuCHchonMsKxLpw0OhMWXD
eo7qJ4UhUT9COuwD7w1RdwBEfCb7uMkdH06CxpdYc4zY7wlOi+tyMdjvoWK9
YxQpoy9j1Q+eaqJPA/JciKLn1A/SRr1dWFCzO4Uyqyx7eSGpwEVxB6BbGLNq
/s8YSI+hlV+j55QelOx7EY2D005+xNSZKWfU6QFz8+GCxVgm8Ty0jLSmL5h5
+hA0dFm46+hnrBpUBdyG1yeHouXWG06oNeQNBsSMhNBYL3VH1wdmbgaBVpTO
MHa7nkkfmL6Zyi4r+UnaYtHE6ScV2j0ePmOzL2vMUF+wT6k1oYSfV8i3qQ23
/QY1lMI3lDYqzfw+Qd1Zpp7wL9P2rAg8Sa6ncAGjmwiXxPgG9JKPJMgnubxi
mqZdQTYDf5Y80bKK2WmqV5AbYRKMPwgl9duLxVKkYo6zxMOcEjW4VC+xqKPf
36zi+Z0ICkOZggUD+HMqlYTVUA4mP6ucyToej8A6HIVBXGDrH/MCWMM+WpT8
7DCa97J3iazKFOcAJYHObJwqlV95SfwYrA5305Z25StGKYH9Cw2PoolYcFUP
sAGIIIipWrXZ4DMd4imkHDhukcMgLz3cIMyM6VWOyM94CJTZnjx5f2G+CMpp
6/8Uz6X1zEdwVI60xR5U3PHVL//ASXiwVTvJOtWZGq54fnrfIAmHlqRAJK4K
EijA99RmV7HVCVi9lDcoON6Nk6FPJ3LG2zi+63SPfb1ZwqOuzo4K3SFHwsjf
3SvQBRpphks0QrpRhX3czmdJyyLAv4INnpKV9x5eHXiC9QQz6QwLlBsY9r3P
YpEDRdHTsdoyUQ+NXPIMgsNSrkZSvqvCeNKW8YFmYftoOYHU+nuZvdlifxgx
sBGB+wX9gUYZ/39MfzuEwbGMy6IHF2zM+43kKUFxANMm0Up5o83uM6m5BAcz
V6tao/WMbwaKzHPRjPBZ5J6DfRaM7uGlYj1NkjkdcKvWh5coq92impufQVlX
hNB+O2dZJ9QceVjKWFqGCbOwk8rf3cQk3nY+lB3BYKHvm2H56GuEFji7l5Hq
9eGNRD+1s23zAPmUxdlJ1d0xD7utyjPjnbolC9oLLDEaKbcC0aEc5NE53upi
ikBzSC5kRDMHB3cxL45sJPmzdYnaiJI+2psxo5GUL+KANQaPAcXpz4Mx0D14
mZs9xQjxzSbyybBEKbRjipnIkmABZd+n3KNcSF0S+F8ITYO6ZGX33PqrKelQ
fzVz5c5daMaH9dMwhQk0nKgxbZ6yTnI0Rm5RbqqzlFndtJrlbA6ca/owCLMx
Sry96gfHDXGAcUhGKLLEwAZEAXH2R6+XivmbAi+pBuZWtS+pUxzoQZSuwtfl
kI2c1tYOZXVjWBzcmJLc/bs50aF41dm+3rE/MO4GkDHwGetMwo/PPiniVyoL
EPjrTn/bJiThtJC1BhTxRaH13A4Azhy7w4ApMoEBkVah7m1VsTu0aJYbo0hC
NzdAGkdx3U8FnFQsud227IiWhbxoP8UUlIPEe1TZ7X41SyDwFcwIj6JOafaf
IDlEvMJKr2Pd0nIgXm4qwN1Eii3jlUI9pkPPmnAVf0xIIdiK7dhRMV43lfbv
jtaQOW4E89PFIXYd4q/yjr92+vXev8EuSYfW30oZVbbvjA2KRgVxahZJOYHc
xha0jCcwFRNUNE8I3Hr7DljCLpj4KcLmbuuEcATMTvDyM2bbw+Sa++dOpYcz
MXOwG99r3WRN6+3HlKjhZ2fZsEVmZVrbK9F1+UBdCEwOaqdtqMRFCsLSQOc2
w8GzqIg3glcfllPc4yiAoToeKwwX7SM6oWicgdQL4QLxcAF9pLlNfEiGEEAl
Xi/tqyVOsKM/nQnL1j75qJxK6VvteRnTe7QFgeMsRIxqA7Sg8DNViB3C8BHa
eXjfbI9hpABd/xPm+QRwcl1bGt8JAN8iIaIzhZV1cuzSXseTvn08K0i/P8sT
Clu/mGmmDTWCWVnVjx9kTWL96Ud9E16q7NZd9/W8uV375t0KaQr+5d2gH/1g
gIkEJHmjeRWMxAB3IW0X4a0Fk7oVF7OnQZSvmI2TPQJ4Jx1LWPUYtkbEQSJV
On1Iw7XiYTjQGKHaRcKGS82Ay3SKibtfyYbJkLzGopa9lPhU13PawshJEaAp
BYuoHDorGfese2zPgTsJp2R7i7VJC3gCFbAXIa34ud7lIrEAN2gcaU6KwMgH
vvm/Am0S9IpRnxq9fqOVHq1c/2lnIS08sA2klo8/V9Rmm9B0Fhp0kptYejIj
+xpZnk5k0wZrfBrMTT+nWqhVLRm45ixTrklTPgn9TcuQAiLD1LF5IU8XUu6U
jr9voxeTE9jqedg0Xrjr8po6xQrxUUb8facRlbZqioJDQu+20gLYXadXOLJP
BdCeoxXHje57ZRAAYHCiGbyH7ssJKrNOmrtOART+hENoy6qu97QV3OraxfBu
GLivDVOVMVUyVXDZrOmU1j4LS2ZnpkALuuFsOVZF46Na02FM0PUV6xaTC4hV
pgNVTT6nvRwMi9YWgfwBGmeAkVrjt6DMMp9Lg+8/txpLdnH0QnNSuvkAoPtG
0cjqPbhy0KNoUJZrKd9cj+ho187MuJbPpd8zpt5sWH2EGz7CByzz2UW5B/lu
T/8oBj/gV2/4r1moCgkv5DipNL0q5r2t21+Ho+Lrlf8wjGA5u6UupcoLQujt
0PAHT0IzlEp/QOAfsSwJQOudcoDhh3ceoi2Ie7/aRHb7ucaDkUJ285JQgD2H
//x/lpkqVGYtWqdq9/CN5yBRvD6xw6+1S+s8In/gWNlfbkRpSeYiUQ30aA4N
M/QG8GSwUvpvnaXfw+xXfj9kam3BSvebtXrTpRy9UJf1lnQLTkCl/kbVJ0co
UKWdVNaGkRJCXZyrOKG5gYCSMOOdkeG6v5pWFol4UhwwAc3wgPqA5uBocMMK
miNR0L5FWbSC7AKIBY0CnO5XCrJgyZy7ueCMID0Uujz2dx2MCmuGRj6JdZNM
gsbPsoN/c2Ttsq2Taf7n1yfeK0aCCYpPjoW4MQw47AonUxpe1cfVTtPt9qYF
4Ld1zQyEJqG6UAxDpL2XEbQr20K7HvMPOxMlRa+UMIiOFVechT83RSlMOTO1
ID55Wclnp0bdZ4wOvzoTcEGonChfTnGpC0MWa8CgmDkKPo2PxR/YQJgGRNnV
hnmWjk6+SGXGWDxiYqF7On1Q5zQcSzYHEDV7tIQMZPGw+E7iBR+z9DZ408bN
4jF834tLp9ffjcaDQjnYULdQst9sH95KhJ0WWls24v1+YsJUzqSfY9tMWx2z
JgXaHGLcvEvL9Hj+jmB3zktxV1YlvmvCQ0Vyb8JbGOshxqqWG6RPSdHXCXAY
apSxkXP/JBzg31Gy+lW1l4JT9OSEDgP8Viy2U2LBT5FooT7WgkXpmOIrN7RZ
UKDc258i1A4Ux5La+sMLLi1kZFoKAVhlz479a5IexCC+rPEIMk7nmYfHpIKb
IjtjqXAWY/kZ/u9cMmGMuCyZQiuPxXNxHzM0cl9Ia3940gaUN1KsW8AHRJmr
XHoJkVihCCkCfJ0RzyC+TpMkNqXfEq3DrNwllaotk+PJ7ORRby+U9r1JsnjX
dZFDXfqJ+sr02uDopdKXzt+LlSMZ/TeEZgeBWtc0hAWoAOdV6+j703PYHOjd
Tk9wt5dR13LU+3EcYZdI/X0qzsJPnnYmVVFvNa+gIsAiM6mKgOQY0xcyYK5i
76QE1OAqsudTon+x5d1ORJ3T6cZ9uO82j1y4a98gA7HaVoFNWhB9uc3BVXQE
L0xVAAH9RCr0qPwLM48kI3RDdQ+4LfYPlsbqPD9hsbMJgfxZmxAyahKtr6xr
09tLF40DR0SrLJg15ovM0D5H5Bpw676BhRUYdCjsIiAKQJHVHQHS+bouVo7f
ng1Ba9jxfI1salgPKWOmaxrfWjNYnp07zoSoivNjp5wQHi+Bz5rlmRWckStH
fbxuNtaPEhjE+MU5WraGVtVnfCP5M9o3+w23v4xc3PJD9VzgymlVgVHnHCXk
v1c+jULFqO07JCBfm9NBK1SOg+RTuIuONnKEbxvpoM8t+yu0g4FeDl/qB9+6
NwHfY4ByySl9AWcVUMgVqR+vbDAif+uKIa/ac1NffKREfbL3aZ3cHVSp/VnV
8Yxng/L7DEmNwFfe0DfYlC9mQGkF2yqvT+2tIetux4IozlSpcOXMKIXh/zcH
k4z/XqjFEOlap6zWejObX6j1qMlBpk9jDm8C3DPBQb9LcLyetXNNhfY7ukXY
o1iK8J6+vL6WZzh6TNh5ixk2P1kSJEsyaIIyyYzoBcex1DMZ2Zq/ffcO5JzV
sKkdmM6nF2ouXXwFoQrv7J+vHL8ku/3KkjSWVmqQj58ZMW9YuDvrqrEdvjqa
pPr8D/gOLupSsaZzpY0L0E/txXh1PZ9Kizknk9U1uE3Dk8s+vXKdwURKglaD
vLkN9uPluU0oyQV554RNcvddC327PJvZ7xZSQgspWkijpDRbuAr9Bz9Y1k36
TSmWWvSAIzOriXKzIKBbjAEKFJpkwGDk5EjDqQjgMBdY21Fw1I5aaBqrXODq
owVIWl/RHnjFj2p4Cj2W1R9ojqhs9yWsNzLcqzXNmOrqwaDgXAjIUwyltadr
uhgDGfbQ7Y2ka1rRGH3q03c4+LQY2zyuyPWbLIBs3WefSVNa00lBIycSb8MG
wm5TzpC24dsaQflFIak9citnQk1lGavaMQQ/Fi71UZ4vTCi9n5WPwEuMhIUp
UYcSdELbcq3VdufC7VfliS5kndQtPgV9WRMgOlANARjvRRY/uICezDD1o6Pd
YGGESVbSBci9LM1vLGqCSrMbHL6oaXMUFvOHBhDRo83Ec4/bfLXQYbCX1G3t
mGk8qrLjkWfmZ1SyktlgF/LnXefEy3XXG0HLfXWX9xSZ9fVPA5bEJsoIdcJ6
Ad93g1RHC8koUPwVFnKKwdRCr6xiQ8O6eT98qGPz1OzF7Y2N7WYKXg7uJHUl
2p3YvcOKLn30UBB41+wMak2xaiotyov6zZMiWU+gi/qXtk/w6l4gERNv3N0h
T2oGsd0zrA55bWDdT2Dg84crSXKojVUMrVGfGS4tnjeiwb5/o/Hw+2o0JCpS
J9/ndhaIjxdQt4gCcrM/5XGKtjmWrO3Bfw2olwOy9BR+nLoHOeupGWWvpAzD
4r5NRAkqoyONKPssaoicQjyzFuLtIaTXAAWavxOrw3VWT3a6uSJxStNC3cP9
QU/b993zkAw7qsLmFRiuzur4sed6fXvIEdEzjfEBuu1cXtzv0COUanI3V4rX
Y1FTI4YQTwFsQ9aXws2VqK0qBis7EssSE/80wiMwmX2mHCLoJ63MqmlsUddd
djY7RClCbZHimu1smo8owSI6Ctez+kZLNSvsurA8lCDH33G9q4mqxf1ODYL/
K9subI6OfsFdRjY1CjhA8peVXleiPIFrs7NlJIhd1XU6We6kFyJQyTD7MRsY
PYGDEZkIEsqVqK/wCt4vi4Xb87iW8ccHuRXYdToyx3c8UTUeFw46mpEcGfhu
57eg5F4y4CVtGN26rnJIAGNETdEaId/2G92W7p8Og1aDgxU4YJZQ18y88rsY
aAksjjB9cMcErZuPBCGhyi/6fXFAFn2aSRPCr/pqIGyWilSAHpDmOUGmtlG7
5d5bMwD3wlA7p15s3Q2svf/d020m2j0IHOS/ieK/L66Ovcgn/Qo04q4Bw+Ei
4TedJ5mVQpASVfbgmqDRN8ySOXpl2cQCmCE5DLIvpY84YJWkYs7CWbRKL4RQ
Agaq2GaF2F2PG7IcpSG1FGWcqQymrg9Rsvg8oJOBDvWGy808oT1FwXEmbL+5
+3YwBjuecAifwJxkaBL3mKRs6lXb4pIudUG+3J7BzmaSDm7yzm4Z2gfEDOMg
GruLxsfExqA3h7WI7ap9Pbd4msCx+g/cCnDdjeMe+JXVEt4WIdeWixi7pmOJ
49HMITQCuHR7mY7vsTmDracAlRtqs0QbWHucQ2mzAmIwuETzYCoraNp1UjLF
iinrqmedSQZXEOVAtuVd5C8JfnicNCO4Fd1dk5QeLMBpr6OuD+9zKh1YntE1
W3psATMe8dJp14+cZd+6QriLvGUMN1RphOAsVvxegwtL91vgCywL23aHOYpL
i8ZY3WKjxzFmwpywXpAWQYDlFMfbTmpXlP2A9f7RWw8zNcS0Stvc44mt3ra7
H9WRs8/lN7yfbS0MCDSKROvfMRpyJ01moyFCug7Z1l2ytniOVAEXVjeqqFrq
nEs/XpaSjLjjSAkV6l7gVC6Ob/jNQkSrlVWaWoO2YAK27PZGLLuGjcVuS8OP
o7waiA1K5slfSD5W3DT5sEQl46QhOa2AcMAvTSyZrwBZDF403sKVzLkIBEQX
9sIx98y8VO/lKQuex9XNlSSCSGt2WYs8BmPCq+Y9wBQsxjl69fjI/I6ymNPS
bvN9Tt8hSGwkIfUDIjQD/ekGRWmli6dXepMS80BD2AMWV5O0TFVpjiCDREyO
Hq1MB3+Kp6MgXKrj4cb95STOGDIBvUzIRButcDT9cYPAWOplMkic9hsOd75G
azfycmxZ0+L0m+JksS6NNXLc7U9M1pWiNxrBJf427iMTPHmubMZNSSGgkQdE
RcAcbiIQrhjX3PWPMnMTLkcb57G2k2w74kFk5eqXU0eeRar0TWHf9+nae2W+
uLlKspQGAVAwUFnDTcN3wck7yUga5OGw+lxLxPjGPmF/+qhy7a/dD1pN5QeV
G5E47q+bNRoTrcnt87AnX3Ji3ARfm7OhzD08kDFzS+uiw60MP1gdzwYS1yR0
Ep+oe40Bww2NoIHlCzNbxVNWoTNMesf5nRGzKYe1rxZbQGNf2QDXYHBSfMzM
6ZPaXtllVi9ZKjGJi2ry6i2Snz5eW2cDtY4ZhZm6tAt9csbZlYwLZt05c7Ie
QK0wExfGaHymQL8KgMzcx5N+xJhVMrM5pk371NAJbEFqhr4xziBAKI1nXiGj
A11FwISLhS/qkn3Mz9jGXR5zBaCIMjS6CMX0k/TgamEd13mtp54IWRJA5KaR
uacW0em2rRxFXtESw1H8Ze7CQEU0MMfSGYUae0ILnXdqni+LCU/3aV7Rzb4R
VlgKne58p5iydDjdqnJJPzTetwFWzhur9r7RLO2FAryr7xZ9yM0rwv1bY0DT
Sre6NivGysL9hJRJuDxZyP2AfBbXxju9ALkmOmyw0kOG5sDl0pPYUWE+0Y94
xkyJeZ0njY8rfrrhOHw1aF2JUP4/ENJHqnGp29nSlxuKsEAtUg/dtACOL+kC
tWChVgYBNKVHgyF1lMh4JlWaeYYsqFkAmM9/HgJngjnHzsNEIb0FDqretYGo
gXLvWXyo63IReYhJCQsjscJhgzlM9o+24bhI6H6pxmz75mY0RGMCUDP0mF/o
YJi9eGheh9c9569T7OcLg1pChSCgP0K0ub9FQ2TpR2XIvPL/QpjuXbww77oX
+0eCyGhSeeXCV5s/Oe3qWB0kS/JqR2UKl254onYw1z0I1BS70lJJrTCqs1qq
Qj0qC3bC9dV9miUp02sO+8oRd/JiCrkZ9829QCqPzE56MyoSFY9SIymt9cxD
0rxlEbzovnUbAQKMiijeTlN2N6B57hK3WQOYzrPzAz8VF2vIz0+inEip0537
vEJTbfF7BlhHQqVcRbfMf49HaBzURdhNIawXAxdejfIgpftBQ+h17jA1lxmF
XPNOY82Y02WbIXKGmbooAKMjy9V1lHqiHtOZgqf5BhpQOSwRzrauI2WvOcVm
Q2kZginekuqXau00IGjOO/6isZd62RjSu9VuRrXa69gJ5LZTbXO2hGz1vD0n
F73BIk5AUKNEXzMRqoMy3D9UK09iJIH87l90zBq2SqDSQ6lTT+oBVy9h09Lo
QQz7g7xjbtyQpFnh0bnzude2bLgvBN24ZJe9kykCQbjp1UgG7VQTSs7F7PKa
F+Dik49xY3Xir/J/e/rcKG8vTTE+326ohPFfwOcRIBD0AJg3nfVtsoh70EHY
aWsYmBAOIFL6b+MLlArK3QakDGfKT3Vjur1JPDlbz9Tx7lNM/cm3tJFMmYo2
ByTRU8RL66RdsBt90wrsltnQHrbR4q25jSdVILjApkAdNsL/bC17UqA8o6an
KxcvqLboG/ZZJXUT38ZfFZw5CaR6/Hw/vdn2AhxKPonMr6gJUsKKCuAbwLK3
w9/JVnKBgt7di7Tx+GOvX57IBSZn3yhIUXdjvtvIj6XrNHW0NYnLH54zfB5u
3h/aJhXdfPhtPuLAhHedzrraqYEszWBLXe9sCZ2lZ5Jrb+1haMFaOBK/y/8K
pVCAT+BAYRohqYgFpdtPnWjXl5OgDJQK3p53mCWjnyEP1d2v0MI1Thk+1hsZ
WvZt2OA9pZB9B11Ndf/WlU9GJTSrMSoy+cbg88bchlFOsuCP5WcISBOacB0w
AMWuepfI5fm1capGlE2hVi9fWh6zr2xh7bGkIBhzJvRCGX69MCT6CMe5QdTg
9ckog5Dkn7ojZuJbjvrRtKTQ17CGYl4U3fVb4GfMcyYWYDOZkfK9a3yth70k
Gc3SIryIUOfcKHtgz0GZ3ucvkgdXLP99eV75F+gKRusBKqTJ48nVB781qzLv
P8eP+PeyePwoWM+Sy2ACCy6rWVH+/IcKkhl49R295w+DKnR+QUrCPkYEU2a4
D1dPnyDNVsSednFzIw75B8nUPxALFGhAPm+3HQFc3ILcoBgYO19o9bpsi0DG
wqjuiBq7XYXKRRSolii+i7Z0DuOdDH/HdMxAI0Z/jIV4pa8Pl/38D961knBa
wABX8aOwv2+PIpPkohB5UiTenZ7VBDGTjifvRkQ1+PA7e5G3wE2CIsQIJYeW
sfCnWFnSUYA0b+4Y3aYrF8YP0dgw27+aYLHvcv0b+J7V035M3m83ObK17ZKs
FxnzrVLwXsDVzG+mCBx0qUFNZBsJ9LUCAz8h9CRZAZ4PuavR5NrxkwsOHbuM
Nw8DBaFHC1ES6qGzOjAr5mR930PkXaKX4CV7nySh+OQ8QuYk6P7vCoHddKFF
7dx6lBVSPn4pCP/8dTHMUADoCM3HLMS+kLqYI75qTs7TwFQsmcwTwKCxP82W
7VJ1SYA61YhdeVK9g+RUN08t7LRtxmzXjZkzoyzsr52IGuA4N2KM31AA5Glp
YwhVx13woh8rovEZ/cCcbyTIL6OnbqPEDDUKOn3KRiyMzMDN5tV676CrPPa2
OXCRVReEwrovb8fML5PtbkBgtQ4ATPKN8FsmNWEMknDyQGKQR6I1gTb77VVF
mg9vlsOHjG2/STg1cdjYPVF7cWua4bj8bhoPVndI0bg9xARJlsysjld/umGE
ZrdiNtwZHV7dy7l8vbUk5G8kuISTv55YNMXuVsPVhN8+Wxty+G6jJEzk31l2
LRt6BRYBDTYaaLkDLmvMMcMuavY+s+eQHab8oo1S5+GqbcswU/W9GAV7sZyJ
/C8wfmKqPumGM8+9FguwIhmeyMIBuV5HJ/QWqtXxPTOQQ2o+TYH3WkQkdVFJ
T9qbqE0AjOaLzCStfivJ/0Gl8Yt4jIS/vvFuLq1u8XZcnspa5M4FOt+Rw73X
kanN3z5OFd87V94IxSPPFvKWRyqcdSPiLy7bmfMvBK/ho8SvOIsN9yU/TS70
xIKK9oZ6R0UeQ0oUzn/9k5vZP/vcIkHKvCaNsmb7EA9uWpd6wZ/dIfN8Gcwk
hzgQTbQ5/Q4BTrI+J0/z2iZSxdCUbW3UOOYuhDCzwX7O7DoFEyRny68qGJ7K
2zaFNqpX2Bh+BmkqCVdTXQ5ulzbD6nEIb/11IPbZVQV2jkfV/ZI+nAaI6LTT
ZYOajuiLaSDPZGGP9d59X6blj4Wt251jWHuwubN3yq9iIs0NDujxvUBXU/pC
PTqtYQFjkkpbnQesSAYG+cKEgwWaFqqsGWNhgKd1e206Qf97b48rn4tcLyyA
OOGUAonAWUAwbotKm7ZIEUV+p3AIDkSc/bSj01tPNanzfMiMZDzP8JlHJreP
lw2yvkutXcRl6XFbWFcHCh43xD08AYfoz6bhZM63vU8pM82pAzbby2NplyIr
XchwA/YHzTgp3YdfI/uyH+4+7/XMWIL5jJalH/PPtwRPn7xbdchpzaTr8mmj
2IA5Kw58Cv0ZZBKXSLZuh72HHYqMqlYMHY66nPSoj9x2E5RIEdk2/YXLyx15
Hq9U9CJRDA27pYzzOxnpyiVAp38beuBvi1eOhsaJRpXPEcuae5lCOXlJlv/c
VGpSnfsicK6S+aoEi+G7bxs+wOHj28ddGvYVLkQtDV8rgFOaZBIi31ZVGMVj
rys87xNZeokgjbeicPOYrrBN6CcbHQsD1NBV/g9esHJqBwseAr5RpWRkrp56
/0vwK7EtyoYRvWdBfPznF2qwmVaZ4LIueBRtngs4TxpuHEi7R8u0D/skg1WY
9WLvNGw+SUSHANzZjkgZkqP8rVgjqINyal1S3KfVtzpY7fHJiM0r9CzlPaAY
nQwnf6leKaMrn1cZFotC/tiKbyeWv50WPXm83QCo5C67IAWV9sYOCrEmnuKa
CMT5Qg8fM00qo84m67N9qA3cVWRvcyVCgaudhSr3pIGnRnooZaY7B4SDrola
tpwST8ohm3QIweTE3iX0jwHkecoTrsOUG5gbD0rd/6lTi4KFjLiQWglFZfy7
PTs+it4AjmvIxslRc5w/LFdjstNAhADaK8j5Rt8JDl5mrnSbDlu0rOqfPEhp
WwwJ1aO07gQpqBsQkC43mK14ji05Sh95vAW1yIZq3WT63jQ7XOyzx6fdSt/8
Du6M9PghF/KZZl6811dTe8qdM3K6NNDzSbEI98TKZSqK7ZwCB7EcIeXn2xNG
uJT5zJKpjygbzU6MFzwkFCWv2tDNk5zL/9FWgJ90SPKxVL/aCCk5zOTW2PmF
VlOVQIxxRL9C8EAtefGLf5fjcOHNrM8ysQtQ+BL7G/y99TnAc7OoDQSYS9yf
QwmFSq/0dB2nBLGH2NYx+P8S2Pirl88zEHHIZ2kORbTh6IHrfMxQsMnetVc0
UvZsrPOF4mSAQm4UA6VPi93u1ktgxFXOD+4W1+O0U//Nwv0FmBB2fSVkMv0T
8TllnjWPaUgrg5va92l3qWWxGxGS7YOYucDF1SIcRpynlnPT0s8Qk7DhuTze
8a5V9u0qBnd6cq1DcqUsb1SfBzO05DD9XtXsWBnCmp6XWcTmzhYS0VRvOw0u
aGmd+kM/vqPtkL07jUFn2Tv1zLvllCBYJ1b+g4VsZj5BPNDt/1wMFLF3eNgW
Ybw3rbp0pQpcGu3+MuPChmUCXSQtDRz+lDF+gWzUBbnmm1I9QNaa22dxKjVu
+kh2JwpJhWUMjH8ra9mtRvlC8RMIlQaG+3XrviH4I1KwyXbCY0Yyd7HHXxLk
13kGpouKavK66Lr5A5XmIutbzhAr0w3G59RUIWMXeR0FzgepYUjGKXPY3l3A
sZFdfRJSWhh10ZN/8lb7ruakSTq5c6AG/8NhqDdvSXIwTvz0zjveEeKSFa2K
ZUddJuXYLZci7ezpO/TshFb+P5qn4cBTKdZ5oSjTv9cyC9pTLC2gMUlGJTZR
fpbBmRmd+UCtWxo8e9RK/hEaj9odbxkOtrCbn5lLeMUgZuzTncZGFOOSSnwt
ItGnlwi5hbbB/vXlMWfQCDvppogauQQkXU04PWKF67j1MRq5hTmg0HP1/mNJ
gU5kK9g2qSz0j7L8QGJK0nLUbT68QBJzRvK57vEqAfjv20HaUDM+V0tyjUMB
r0dymybJX353ARZYD4hijpdBriA8pdAiZzhXWKmVYkzil2kooFLfKMkcP9HU
jVGmHeVz2k0uhnLykl+p2ACWGF4b9XeOfVuxOf+QF8JEyv6PWaiwXxK5M73a
q241BVUEcS7yCIk5DNoBAifoMzKeBrV+oxKCbrwGmRblbbxforQWclHZxrE7
SpDGwdcZQ6CJjotXvwrRJzt2u70+BwmNxP74btVovUnkxzgSEMgrYAZH4NO4
yFdtpW94YkwoNQKhVEhFe5e5xTBIR7lPTRy25ZSroeEqqYai0acZwztRjLsJ
qJza3yhNIrpgucY8wWhtOgwr8f/aO2SN+bKRs2mQYXhRueEcl0OJ2jFQojli
eXaOJDtFYj1crVaE7l3jF3r7k/6LbPbi733K1mqmj6mgk/gH3BSouf2BAAbl
djXZJ/+hBT70NIexzB0wYFRPExrauPpxLlcP6cyxOwQZPept90wgaKt9Ual6
yZpvt3V6QlyH70ylZlQXj6ht/+mAEOzh996Cv6GCpQQe2ZTJbY8zK/EYXTaV
FrQ7eH1E9p//kvCimK+jtnP3BR1G+5NJQRWy3nV+TCa26WjxGjhXLboAxB33
PFiLz4RRKGUEBwZqBVaCq0xSjP+JXo/Z1Gsqo9xo8X6k8IDEH94y91SeYDri
uS1dS2NougqltV0vOKhVIPST9dAd4iXGP7t3TSN6Kleph8J5Rc0Ew3R422ji
iJa2KtaPwJYxvxkUSkzsOpdCIB0ptH1PhayHMlRvhoVp7/ZwU1kdcaWB9cc9
ROIsj59wY5KsJOkzL5ZJwUaXzCJcHnMQ88ZdvnCx0XyjjFEXuthUDquyn5ez
bsvO3bGlNOc+RQm5kvko2o7UVj+R9/snUeu+CWuQ/Y6KAIJNWqdI/4B1+lkU
6Jauck//Mvtkcxgog6hUNijr81e0fX0JD5jsLIFP8X0/GGslETYucm/pYf7T
h+ILO+AHha4xW/gzXZ7fCUHVxya4NRa8KMZQQJsOeFHvvCsUPW83bJGEUgMo
GCj91EErXGt3XtFGZcKLs8TFo0dUQ1XatLW3stFVrtZkB9TpAlnZLk6WmzCh
zHZ2ksTOhHVtGSxLO52gZ3dNZ3Sx66XtXwu8uhIzMB/4gVyI0KN1GG6bRJvN
v0KoVq5SU5InWGX/xpG9BT2j56LfYcwFM7D1uuYQydjMJFPmtBM9UH5ObMQG
4WYKaQcH04fr/PKcCmjTY57Wq9FqzDK5ESwUKAPVx2pe+7ca4JvTbineGRox
JXYPnx0EF+NSOahe07u/c9YQdal+FT+g0fbVjISHRv+1OrcPUG/JagZBmbNX
0udi8WYtMqgb2cwsqdW2+Er5CucHFqY6tl+oRN7CnPQaDpf9kO0JI7Zc36St
HlvCQQ9dHQI0Lr+7pSDQIYTBnCpmXTm4CjI91BQ+r417dqwxy33XVBxohW8k
8i0fS/j5lk1Igcd6ZkKf59pimL2uVDTkZtL4wNnoaM5c5q7lTd7Vtn0GA3LZ
2Ht9p4d2VfSZkm8jNjF/zNOAvvba2ivQLlAqX0b2QY8GGpCgACrtUSHJEf8D
bLoGf9KZC4BTWazxXHk5yio3xRCGt6zjZhGWHyrfj/fYOQyDv6r0qcg9vHyr
paNHFlT6ulZ6jbRBbYhW6uJDUnlrywlxL/ceGSdeDsZv12b34/VkZ3yck+73
HYmP3mSrETvYubwvHpFIBsWUfrp200W5iL40Z1HgT7iK9JSsnR6g3R7dat5J
v4db8bRYb1kq6bBRv017sGdS6qNbs3aU4XYwd6Zh/8eTPIMVi9tps8taQShd
Hh8R3qZxcFa06oOKG8Ubv6jaaqB/O9y+eOQWGoid4yPukFgbPC8LZFbNOjK9
/2cm+/pgNtu6ocdisNzCpoh6yZB39Os/53R0xVjkHgom9fdQI5efJRpkvJ2K
tr3VBLFZXuOvgkzA1FQYkzqKMkuZW0Jmb+W8taQRKAdjGYut+iOY2Kl6e/yj
Y5qFc8CNKj7R1cUh37HvhOWaRyzfqhYS7nr7qXS+CbmXewStlcoCD0oxpVEv
puJCd1zEALBLQoYkqNvgNNyObHHlAlo13cv2KQQoLQlWnuEDlxy+vl1XXXI/
pHmniwbGyEPEw2urkWjCBPRvICW5AM8BdksU7/jd+QFWbkWEK7cXj087l11a
eP5HNiwOyMBwKXdBeOmnuFe8lwgem12Ai94Z6kApkhcQMg8mgRD8wdea/DrC
9YZmZs1s//mCBEYfNFAq60RZrw0/4fM5XWaRwMsAYgRTJEXcSU8qBdESkOhT
ygAxeji8y6hflA9ZAW7oSqtgc7EtWG3jgt/TBv6C1AyM363TgoBtMfzcdl/l
oPAYltV1NtDR232hMZPThNW2Bt0GxsQBl3n5gr7DzoBdvsec8q4C2NsQEeUC
3CQiWBziBLJEUVG5SDf11Ktgu/OVNDIZaWUSqYToWwr8i4b3b7MLHxGx0m1E
HFwtwdKVN+faTKnylB9M56Lmq9eJePp+gpkdqRjYsgzLlKTDV06T2shKCEte
1wrCqnOyYWeGHfg9zFXJJdEwi+J0u5qEOHdcxeTBBGhKTc6jSbgqBNgspSyL
cy9TxLtdRrV5jLsFfqBvlazwSTlP8udzlLKB4OPd/4LPkvHWyf25WmAj/oTR
09jTji2xDtSPUVifcW24bDyPQQye6wMI+nNVTrQbk1pK6Zq8QEPlFZQBqbxU
m2qsu9VipjDZY5dBtpmgh1oRdnzzkVQ59q7ykI+ipmWO5BwqJ5bL5Zhr5KuC
8z2JvACE83LyZQ29W1OvQBWarmbYQ4k092keEwff2qK2uev+roDsumMI+ubP
gJ2RgmELXDVb514P6qvl3xW39neFWYL3n4/zj+H4lDeK784jJq2oqzog8wii
VgvZtlRWjo6R1UIGPWQ3UDSBa+gQAIb00y8xj8TymJ4L3YMM3yn94SqTS0OG
H+M1esosFPk+DMAsFPaE+IHOIlV9PmTSUnTOWqvwvvkEEHyU2VKsbB8aGMps
va8sbEDtZpmSGcdKesPn+2o5dvuebJVgp9LjHygfWlVzBtvBl0ZGewwpHfna
WTt+8QxrO/ylpEde3YqsTNENLB977zMJq4dnMfliIUG6yEhD3zSPBbPPrIYC
2C3aWV3k6110O1ZkYIvZSnnJaMw/Esq9Oi75pvDkE7OWIZbpZUGhYa51IsXT
zRUgPmsx8WwHp04YB8RutmoxuqGNEHwpHCyNXd8/0fW6sQcJjUQKW860OIY8
ava9vegapHM8c/rHXwF2Gg9Jb0BtxLxtM/wNPPLob+iouBQqK8n0tfXu4Xnn
3Ktgsso9X37Uupcvg4p6uA5kbVFhoy+XS6dj/llDgetbw6Io/MWWbw+LD42s
hnr24MoMww2J0rMVTIt5OoIlc8t92OavN8BCWvCnQ8MIYEh+iGdpOVa8lZVH
6vlCegRTCjSQ+C3/fL0jlABKNZNfIgepR/2SRydPDgb4JtWKeWve1K/GNva6
wfVC0uafwYHBgwEy47/xXur1A68KSgJU4clZPpyZY5W1Ih1s+x63hq2raOpM
hv4dAA0C/2z+xfo+yHcvh9LxggZVYku1ogzsNww5aLEWqJWbFSvPz2PP+CUi
U/w0A5QYCX8MIdOcBj/Xny8QXvJR/YZMOwGGxyLOAFqPwgGiiIW0eS2QBwC6
o55UzFyfXsrqKGMCTjZa7YJq3L7PCr0QZwzvyQdfnjVYDx0xHY+Pokwl5ATS
YTSbQqXp9YgDLCA3qar5U1r08Nxo5DHgGj1tG3ON36rmbORFXCCh/c7Ot83u
tKLzDln+TXdmKyW36zzVqb/AwctCkp4mfyZA0BfE1WBQy3o1l/qauM4vjIfv
Rwj14TuPuOHgIGOpNq+a5WgZn87oUv+/w8twFqU9UA/aav8bnofht62X/3Zl
EATjhSX/TwOod1zCTZJdBnMIs0qagiLwzp2q8inRCzmxBr5ic26Ozjl5gfoF
RlUJOk5g3Ojbtf6swnw+FDb9of4d4UeZCi1LKc+TBW6EfWOzrjpkniPdr24W
JaZtlhc/HSWtqZIgb+vaecGBYKSXdStvseilErk1yWaNGu53LrNISay0o30M
go3Of/4pigCX0NzzGE6wa2hGb3az95MKoOIO7NqmTGbaPBbntrW4kV2Jh8yI
mMeqTE5TvlX66J3CIvh2iBg6AkB2Md4XdULAPfLa0Bvqc1ge7g+3Mj6Chbm5
dGKTAlFPH9xvD6cHLnhJrl2UoosVGd+mLZmhaYjgX56ECesA+CwxqUGfdb1r
x+UJ0uFSAJ9ZjAo8qANDVIginGnutMv0z9cg4yhg5ZZkB5cs0rg6mmaOX5it
qSdcIRs2v3XHx/MdWZvjIVpiHKiS0EBzX+8GnayBynybkkQcOPm/SQdDjPs7
yVwj6JnzhbP8UPubAiUt5NK+7purVcVCV8mdZ5V4wtwDMbTalWRT4LUMhIiJ
zpyt7YrpjW2olJ1LM4d3oLjNfMIcWe8scfDln3djHjRj905NkOls7H3wtc94
T3K8isSbUOywv98qcsA839Ri2GfdSsTOglr49GGGCEbvAJJWYJWzlJeAK/Aq
1jGt/tTNIU8kGmQkFXDuVojPviJz0qNamJdHLbSRWhOiiStgy8pdD2WiRdry
0GnBNaY0/oawPEIJgyreFr6Jy165n/51krelA2IS5lzWT0Bwo3D0CSgWMd3W
kU5SpBpZgc6lrqrxoP+vRSC9esrKKX+X3RAW7yipRjfdxWqrbhFaTKmWPKaZ
7Jbcuz8Oy+vNr3EsrgaRmS1JKnKp0O4VnK5UozS6fJdDyHJS5hNz/5Bt1Jk6
0NoMehPrXdypBK4zO0GiigNYTaxQ50uFl/dqNtuP9xYzSmd612n6DlX2VjAL
deZQf6KUlLr3WzD5vlRd+3nCBNmUdsS5QkxgTNtFmoUQBgeJ9DJFyunk1HWq
H4HoFwKJXBxO0wOTvfvlwsHPugXeQHwi/fi3jT8M0zQ1JDygdMpwK0P+X2L8
gMt81NWVcrr3dWkFhwEL8s/jaT4qv5U7zakjGRIz/Z2dSPv8mlmMQGAUvQ7X
SApge4OKR8FTrkjDhXPKsYPoEuN2RVbBOFK6HScUszCiStQnib20gz/z5gGa
m6bj/wF3tXcAwD31dn/GBgGUlduTTJW9pMgivoROufIG9lKu8SMURPhznesC
kh0bGdTO+wmS6DXGaIw682FH69B5+7uuX2L4ZuGEJJvED8tifdv/zEgB6Md6
BBM7KwzcT1c/4g2fTfiXxCWSD+MSVqU15s1j76k36qr7buYwsKHmPZAUkw/4
NHqSpx3s8x0V2rwbK5qd/+VMNT1gWeXQAWfp4rn1cV2jZ3pQdFl7Ydj/Bbak
cdtvitOvp3wbHzJx7c9lZ5S8wFwWfwNYeXcjgAJYWVi2fEAmk5d728jruOfK
UZ0z/f9kqqtsB9HnBvMF2H3MfH1qhW8bOLxgLQMu1tiYwbS1ldNbw/bYaQ4i
8/gvfneOzPjoNAYC95EWydfK60GtoESzn83tJG/3wRxwUw7QawWN4Xh40eGh
lYdM0vuGEQ28l93wrWRCDddTSW3GRqUIbAB0bSG3hNkPLJV5jrXgTApQNkS9
xW0Fesn+HiVdw9k0dJsg07QC0WCYF2np+1wEDCibqyfnUH6V1XHNgtQUkMJn
/nNJ9LRv0ATnKs6U84p94p2KB0y0WfOGmgEQI5OSKbzmruYzbS5SBlSStmKr
dwdvm/J0m+gc8EGlxvX7fFt60ZETr3dT/nP6ziqPZTvRnaw0ntKsw+8N6VOA
cdgLn8FVQfLJ2SHMalxFYO3blkgocngSbAHZBHITw8KCv+G6noO2GjNIAcCW
wYAwRWz+GJWP20fj3yuEeZeYYJ7B8KZOyPbofLDAbROBh39pAhFSMN3BXT1h
nS7uWd7bDnNdtwBDIn9WVu12X7rxOzr0znC+FPAgIVn1zVK42tK7jCFq1JI/
4rcrw6lSWAXE04X59ebVee2ktrPjPBDdeToQdW9+zj+9/hyL0cvaSyWAq80a
v5NpwUDCsacrawnlvBsFeyRE3tCllG3TewHdz/86EaB2vVHJK8OmmF/pzsMw
sdkE1rmjSP7jmRQ168zRkkTJuIduQ7HK5z233C/vluazYs6WTlxcZPQGyxry
uj41oirCBAsz4ryZvhfnEiN/NMMPqpDFGY6JZystKhb8u4W7cmc/gTIFSJdK
LIECy+hCRW7YTprn88LHrA4hKOrrC0huezAZkulb9Wd4Kolcq/BaPkbVik+X
liv10vySFbRzrjptnHjzPbeN7PSENjDrjpL0cP2X6RP5x52J3xp/T+3aFQJB
HEeQsbKlsalnZeyNub16JjxJDrnJWSAGxcicSyMac+k82RCxu2CtZv4d9Czb
reDYlrUI9TXtOFIWTRMNzJL+g5jpJ0yW9yN0NtLeRDxX8kXfEUcViMx7skB8
puqHi0RpFgGJ4LAi6dadr2MYmmRR3lNeAnzi8mmmQNBEXRnS5BgQ3Q/gq1A4
166M0CLDx1FNxL3jmp0LLaqAiVZ6k4Al19peObiF1p1yovueputT9nC2qynm
OFh+gnEG1vR6pG2+Jrm+SPwPgTo/Aguv5XKKfFMpeAgqIEU/6JdQvkk9clB9
yBdMqoV64dNlT/oINpfmLD8H5S/FL2brwRRgiJdqa5DuLKzDswwFwtHrZThj
yFENRiNdKRvXAlhvyP8mY2LapgSm6n9oumAumUbZDe0b7SCdEPoVQh0y+kPL
K68WgCW5GPE/DwMj5o0jLy99c6wFxfQk6Re4urQEEBQBQDNaF5gOQmxCaelD
W5ZNjPom/QVsOvET/LRPCJpkI0S3PukROuGNaNbi8viCB5hT67pNxOT0xweR
IBF1uM1dyVmly07S6pIuQPap4AofNX/vQBeXJTYXeA8xjekvSUGkbT0NONlw
P9e5LpGYtKHikrh7NLwwluGquLossiSQs6kgAJ5DD/nc3Xch8UbjY315o2TZ
bb5l97LMPOCeR1TW/+XGrWOZNR7SEhT/mlxQ3TW+jQ6KENxQwgN6qHqUX34p
lwC+nzrV1D1WQN8qlIKnNz/5zFtRfE9XwUYjg8ycnolygVKEmaju5W5Ce4xN
azdsGlKaxBOYL+eFnOqJfVdj1FWjj4piRh1y6nWJXu8VcRviuC3fMyVgmDXP
G6uSj5F5IZhK7Nxhcs5Wp9IQ3c+6AqM2r8/EeIC16blv4zuafIxF3Yapudrw
kIkM+kfsugtU2palibQp2awGTfU2W6wjgLdMZmrgMwLK44Cdw4OC0yaoHENv
uwey/QsZkxcYJPOxyUFEPTqGy+oEQckTGYFgjBgZQMalFPfXBoqolNI8XUyy
3Dj/bNUCitz+VRm2MhgtvuZK+/12haI2QUJZrxu2D28zIO000yrxrwti9841
HsQlV/J8fqms2AKoPOYggQDw/azC4t3+yapypBVLFeABQGCsHcA/kc9LWHi6
sJ5t9wQ8hzijQfQXNVDbas8JFvgr7DEkrP7Xo2gaS8W+RBJ35Qc0w3mtASlk
1DvmRIjRRxIF49R7YR5MYROO2ce7DV4tTIs8QmcXZnx1MqClVKj+9Uy1O/zg
dwTEFULddQrKuWEgF1a658spS+L+d+afwHzPqqT9lTQ1ErqfQVeZRkFCpg6A
FfGVNi9n2o8Xm5rG3FggmrGZqDnz7CFErE/d01XOM6iN1Rle5uqLNdaMOC1O
RgPr2tNqOigsjV/EwhLj12vEyXULbL7wWv41wIBaxMeEsa4seMKxpIslSKQF
Hvkwox+D+F3I4laWrYFuEih4C7nA2/OaxBBVyINh8mV1CZx/jnEsmtD6lEN/
8MNPgUVPcEs253bGCgavIWUK4OyFoeHtlqWFjCIckrO6ke68eDRVhmiA8d4q
DlQgym5+hq0wmAUV6B2iHomvRFZSZf3j9z3bLC8k9t4BotWh8Q+GynEAWNGx
v8BhUiV4FuLFxF3TpUmqUv8AoydQUW+iDXVUfdN5+WeMr7tTWEOX1z9eBA/f
pgByIJu0+teWuM4GHTdPsb7HpQz9gRwmai6t48AATGzQHHdkhCeHNUlNYs0x
zuAWTgBTFRwES4mJCLgslGf9ajM1OrDsbSbpTkDZPK7OqYq36eCyjA6jSvnX
+wMlQdNpTpnvgiovY5PRfjQDCnhpIuI5ei7s+J6AfXjOtJcf8Jr3E1IVhFLo
ZxoKwEU242Y3OxvvA28UINIMXp3GDlVJJLpzD54jvutSUxeqqGipCDd46Epn
2xIqYFnQ48q2Tnha5sX7nVOdxKraqXq2FBvEJBl03dE6BVTxl+XIMuf/cdAa
k+gIFARS8J6imsJqk6iq8KOFC0y9VKEN2r4sPTW3jUiTakW71DgI1BZot7Bb
EJc8qxZfmphtkSV5UOiOj6ogQBooHKSwAq3kFJwNqr4o3+W3RosGXvdMxhvE
PrkIA2ndgWhlP7LbvlVJqJCX1a/FO1hPk1x7MhZlAmVvaRGlIoAOE04GgXNP
PuX4FNamxy43qcxAtZerj2tXBuSePNNS4NI1LmYhXurih5Lyjd+eKMNt8VGc
WYi0vz1xY7Pv5B7zV2CXQRVqmBwEuaa9RzYhZndnq5fIbHagC+e5QfRDeu8O
oaox3uNwUa8rPdplEe5iB/srRkrzDLmtWSPXgpu5CAx2V0mY3GtedRS0sicu
yXpxB4DI4VU7IdcSci8gSfUKazUi+zrjEY3hKA64E+W0iLIJLkidQF+pC4jy
+TVQF4zdIFqL1Vc+gK/T7DIGodbHFxWUbRf8615pLrEvQM8A3IBWIisxpc4+
Mv19M0xcZBmaHXf8pNRvrmVO8+2wgj6qsrKqG+0ORmiJOM1jMw9KMHXVUlfU
eyHWDoQjh5XmH5QoH+2HonDYStzLQESFB1PA5ZA87wANuh5R6kqBF0udQHf8
v6RRh5H7UwoYINlmjly8rKdpUpr7v8ag9F7QHfn6hxpGI5X5KoKn431UHEQI
Os2GQJeGpP1wSx1KAFbSZ6/Abgr7vuf06HdBoTJ9f6yDPH3XMTkuQDX+Bfsp
+3+TSw/UDGm7w/aL9KkCpt1HSmArCP1aucLQTvVX7iDsjgvui2ks9+FsWgyg
b/sTojB61tpruwi2Ozd2R09Hywf6T+yjsR2IfTskvXWiry5DMtVd4HhHicTb
6KMGubhjLHFW8ak8GvDKaA/TjE+cdn+Fe1DyG0t6Ene1ebVfMm1s87KSckdE
tWFjLOP16Kf1i9g+trTscDiLiwjzalNwRz4+ji99IJEjYkCNGA1ILJsC/q6L
pFedL0QmlSQ4kw2AKR6d+D/b8WKvXSMyyi8r4ezcf9qXkX2Wz0midYLirfLd
z30/u3ijOk/qWWhrGF3nX+/Txo1iCKng3Nz0sGbwuPPsHkUZ4izBbY9XFL+i
bVc4SXzPKuoBQVQALPKzntQ6xHBH7I0LeYxHlS8Oe5Cm/H18bcKqehhZP/V+
xP1MxqXwxXGo2EQWD1I4QAj9qGyBvUk9awM19iKLoUnz12UbNlE9a+Y4XQIK
vdWQJXFn4R1l9g1PJiOwjXjH2qfXlHGMg1PUeyskXmJ1e3w9xc6PpFQjc23n
dcpms9739Milp5X8kMFbUukuZHptxIfUqjrF9FZTTzBxCJUxeDcirNRTr8Iu
kXVPlmjxUdBlb6jedHddtVjrQbEIUGPWRpDCXpww+3A42QXPA24lDEUmktUe
MlRJ5NcxVawH2fqpfGOMVORp4kYErLRJuNHwcsHrAG1DaQYeC+Wpm84oMAOD
8pQ2DudsOjRJo7rUpywLAoJ7D3nG290/IOBmAd3gb6nec6++B82NCdj6sE/0
Da0wZ1cDZfsU6xtv8kV0qH0tpjcdp5UHzBKr9Oax4DYQvnEFmcMl/cPa79qV
gcTZUqIkfKhCJZ0yV7GVcN2/Mygm0lNiqPPfWojUZ2oaBFHovFZtU7ZTkpRr
jidNWg3iOrUjO9fk8D0eUB0hQwWKPxXPvUN5rk3Iawx0o6z9dhbH34OUEcmD
yvwAMfJOii64pGRvmcDALNhIGKf2HLTeTJKu9xdDLiatF3lJvhF++vaEUOJr
SIfkDdwfaNZKv2eusYsn1rtU1dLke3R0gk7dIWfv7w66a90ZHrrFVddPVyGS
rF0x3LVRh5l6SKcMBP3grvCmtFiPlxLwCqxFFQ1EaHbY29P4cOtlZQ9Sk50Y
/svJBLXP0Er7FNVOKda7KqRugzROj/tNRwFlivRkqUn5d5N0jN5tZhvg0xI/
vettelklerv2E/maB3xFHMbgjXRP0svIrSZILfQbRaUVBQ9tQRrLTSdWW9xs
yPupMUqW8gelruRPZh2X1Q7vIjbLHmIAfn2uf0CsBdjuz9wl5guThd3VUd1P
tjy2sOdiqyna3nowJeT77qOa9n526lDjSL1ys+paX09fPlc1q3LO0EPxXsKq
iRQDICN8Fj6npTCE+sYoeZs4K9wYHRq9NghoEOayJd9w8zIcso6Bi/+HI/fh
n/tj+NFIBOF4owhaDA4MF4SPk/x8xedKyZtZ53YKBXiYKYwFfR6y7bcF9RYx
5jcKqjeRYlLkNzrA8bOz+D8IlVONFAe/QaJf+aTUiyAo+DvHzdB4JZBBOfXB
OcAAhvm2Kj36rtgv8yJc3NaRGHq2/7KWNQfOiWLk8cON/NTN0FkptpWY5iFV
g+HToY9cge10KqaxpQZALzF/crie3kP74x2XEs5ik+Whqg82SVCQYsVCnUJK
E2PKPqwSaDZldzJkc6zQXBAiaV6Cupw7ADnOB7kINCNwqEd60EjSBCxO4ZOH
dF3IiIkMWLA9vexLGu7FhijcBWt7a6LYX8c7VH+nf73rMO+5p7NjD7JGSXym
YFVQKsKjt2nKzT7qDAa9g4+FYTbOwL/wu2xLdhGKJAbeiOGsMM7AqjiWTwv5
enPKj5ov3iw54RJ+2ZpDFlT8uJu17HNHZRegmZ0P84mn2IZR9FrHj9/vb20h
eIOQxXD0B3pJ0NnhM/kMv8mkVh/BHuKh080PV/d9dG6QGYyOu+G2QliEHLtn
aag1oc44lUKMKNQojRpx/xasZWEZy1h3kENuUYEow4Y6S6CbfCskmiEtNMWZ
XueNJaOHnVlCP9JnP22t0A1R6Ht5IRk7xvCiFJPXoksFW886kNtveiEmGdCX
n41lpv0bELcdBKiutXZnHwSZ2ebf+esMZeqfBMkdDxqF+B1f/ehZ7r+0hf0e
YlP9IwVOXGBnqfZqWTbBKjrJRkkvMB/e1q0PW7l0IilNxBpVxtnPEb6rQAcl
F6toUW05tH+X4oyabmzIHoleDRLBUoQv2uXzgStIhqd5T87hn5+5Mge5VTVq
/0H2GHtcoJxeA3N0qeeyLTjd6BuST9sjkYLFlpoCQ1EJkAFPoPe73CRNww3B
R3rRiRgNNQ4vLqtwTluulLvRndZUwGmX9kgbPEEKYsQ0uFy/1zyMQooyY8Yi
AxtGWlLYmZGCBVCLGWri9H2PU2sSQ7aF6Ok43yUATJqvq1EUxMMrSAJcyxuu
fZLOvunWW7ceuIt0VqbONmJmpIgDkb3VR6GgVZJVQs/H/L6pGO/eKoHV4a5/
aNRkflE3sBXlEzFblvZNMjIxu5d1TGmtiGrOROLw7mhqn1eKasT4LQWCQHPY
i7nGNOIKaNMlcL60hm9CONIO9ZrAp4xScGt+bNnydK8IuLWmh2FpvBQ/ZIRQ
Qm1DEuaUbIehhfT29H6AcI7ueG+BNAyFaRp3iZw23A4DnVbl25Y6rgbKeHVG
UUKfVDC8njbPY0LOfmJOdND1hI4rWkA5LpQLFUf7pxmimez/J84X+9JCA2J+
I+fhkT/AX/FY1mnqSiMYKIVVGKXDG62GXikLXroWfM1buHINmTjlTVtB8+Q1
JtcabluM47ceGdq8Nq8QCAfKfsydodXpTPCRrhUVMB21KSO8+VIufh0ozZhp
dmI6ZVAxi3rS7shI3PByEgkGItDihbg3OtIkatSzCyPa42yy45xet2Xw2P8O
W7Jj/QCf3/aZ3jOaha5x+Vb061r/ZMeUlbwlVnLgpfNOZpI/XfIzLJg2n7Y/
X3uCmnPdh4QZFRC53ecyA2hGDFhyyO58dsgCxDPLlXiDt0vjrbd9zEbaLvs8
bMtLMkj8AYdNBO1GllRPkMIXoQaKlPKrgfDYnP5e908Pg+7OmukESveCV2Qw
vzvCqGEM3ailVkJ4tKOD1TqqshpZrfHcnQV7Br0W99JmPOdt51UfYA4xPUC7
rtHQCw4dGLT4fQd4nkWq02e245BU9dAWjYuWgNUwBnu2lz/TIvlvdnN75L4c
wpxnKYoE7TEMiViMNPlbwgJjTOTfVrfpORV541nbEd7j8rTZnf7Cb7IBfO66
YFlST0JSF83mkidj5IE2JvJG57dgKcC4JRNsLvdhlgPDQ0h06zvHo2HwRfdx
2dT+wVNjf/vVXpWfA7PVqNxODyRSvkL53+CCFeMub1dCY/Sj3ErOK8u0WYaE
HHC1V+1HR6yCsap2qlP4tt/vGbYWECqfeRpuQDhAzgrjryuSjJrrdtR4TMM9
9d9GUF0xZhcWzZQbYB3IaIbx80+piteN4C6OEr5DHRlVtMUhag1hx7nThsuN
KIHjRZ1MYLKkJLvyGxwEED38vW7SysFYS9EJ2IR4tvgGKGyrzFUe8nSll26I
Cq05wQvHdF68EecvUCoLnLya3nKokVsikso1uYatlSr2Wy/VdWNauU+Z+0e0
oLYKLtIHYGhTFU7bUvPD51UkDsiRS7P+L3XRMp8UmsG2uyybR/kP88EkZI9M
5TNiN3h6pCfJTMTKfF8qtc08N0uIlDTwPPUhSvyUt0kJKRxREbZvn6Lki2md
kVStXbUopynGys3iKdQ5yqV6Ybxp1W6Oltf95r8IOGZPQBCW991fFDiKcJTF
vABh6uD/RF6erDf/A2jjDS+5h4kcquI87QiNnuU3zVosPd5GeDmLNU0qjawu
aGUmwHYsBaBDcz/2dZ/sR2w3oQzTOT9eSjYjT71UEfsJtjm9aaQhHOd8PLO4
SinuCirsdn9gBVnXkUIGH8jSqefwjQnDFWY2JD5IgsOXzop2HucgWwrAuVy6
coiBrG2fD5bHRNC1w9XnS2jizFpjzYx0CQ87kNqYKbgrNtMnC5hQ9bXY8AWL
X2bmIPoLtnljVTLB3dWX7pnbTxmjbNBsHEg0S4eLCLeHsviwuByK/JF5pipG
0IVcRSrGbobrN/DgpAlHMExIYWCzq7uVoemCL+3DrB3rlpXxq90vD064mZhf
JQJYUr0oKIxsnANkLPBnZjYyuJx1PihHyLfYFXxAKJQADrQHSnhAQ/4prTJH
jL9HU1Ap/hNRQih83Sr7OB0RzqYk/a/zhA7RW99oJd8xeZ3g2CKa90YWU707
HJvS4FZTRJCrR8RI6YcGlYePMRlrWb56S8QcV2bIoMjWUHKUUCxN2w5dQ7RD
Bniq8naO5g/IPrYe+njZ3Hd8VkF1ypBSd+3qF0GVRoXvi2Gcy6g1Ucr06f0T
oCtQU2n9lf4UpWgXvMr7+WTlFjsaGGUDhnehpc1HT5rZZ03qP0/owb7VdKd3
lWeC/pIoLxgcQQZHLgcKJki+cX/uOmLwgtqWpoyZUlaUgyeAh3yoDKOrJqml
lRixV0Sy+vbTIdQ0yidOkWPkcpCqBC12mBvJYrzinfrcEmdo2jWFAX2b82hI
CtO3WEURi5+ZWJ1oETSUwDD+3bKfXvOh4ORJ1GYxjmeTGa62H+RImWJsDGTy
/li2OqlMF3Eejkdo528eTuCHQJo9BFBEvJmnAbd09vly0gnKw7ASFZFQD9x6
XHS2+FGf70nEzDb1espO9XdLmCPHNm9tEheXnwcg3G+KVASKkaY1oWMr0Fgi
5nCpe+TbDCFdVjJ7hHZTs/Zwk7t7D8wb2efI++r13xdYCEDWNpsSOufLKFZG
wPb5K9Mooitg6eAdB8MO40ALZOXDF0739tNy43lwOlaZsxICm1RnYz0YMGIm
m1R5+1aAldUwcPBGpBQuElkEz4zOAxIZWIEGrEX7ptXsfOUZdOCm4H9xjl1o
ku/hdYm4apfGJfOHpATuFie9BQopmNVhKJEPi/1HSH2t9D5Y65DW0IAgBxNv
RERYSq+kexOgqnzFt5PoaI5NKiLanRLFYomAAWfDstWWIHqE1sdmPBkDgb7r
21w1Zs4nfqQB8CaGnN0FupEqfZzs3kdFBUAVK3v1/ZlBCqRyJNvMSBG79sbK
PGtd6MlPN+loWCZhKoNQt+pBzslRecmcD6JDUclhnegHCCaO5mE+vwvzMPaO
FkrLmJ23ME+SMJar0NRmDraJAK9qQ2+Olm4VQtddc4azsJpKi/qF7DyRCUr9
doxswiDT5unk2Z90Bto/4OczWakpj9Vvq3ZY/A/kj5t2Ks1oY0Gk0xw3Noga
/1pnW0gvg2x6pRcT9OAYxlm6R+0+htK9H1pxTX9CLmsFOJA08cj98gFExH36
PVe2Rs4uQDnEc+/ncvTrtZUNj02F8rJItdZuZL8DXNq+xLais59okq4W41/z
fiZYF/hW0fSHPmjaZO5MRVgi7V+xbaD/XP+e8hqZrBgdBKBetPgZviE6KZ86
O9Zj02WdJkCsk9G/cI0K+nDeIbkdTf4Uwecn85eDUZVxK8WHIQycewXB6psR
Y+7zqvOtf1PPrzAmx+9Y8rk/kO4k5MGJVMKrlDqkrPe/pNyhKqrYcPxr6f5z
TLAOTV4Kkw1Wd6TVE/aqewVDkdoBZBDXudNxZMP8mH5PIQ5WDztv1btO0wYj
12kJYwxgak0KXfAnHU4F+CR0k0YDZEoXpzsltRdzSN4xDbbJYKw9EbbsktVv
uLNCFq+dU+p8a5ar672rVbhING9U6CcJ/Ml+Ttc4flxQCuoPR8GvvhELofsv
cJm/32a1QgQkz16CQTtfw+32o+XRUNix8gkPLJEn2ZY0OdfePonRXMwFZZqU
J+rFcfsJ0b3Wr2u9hf3mWPkVcWXlvnLYuZA9Hlm5+aXjuolWAoT4ARXZgaWE
ffaxOBVusfzU288ahzVssGV7vhzbDOQCkjk0EPzTYl3rbI6zusT994qRyS7t
coWmhZrnnX1+7axUDkSV7cBTJS9TuYPUciQAhWfMZ+CdyhbU1P5tcaSlirg+
nPch0pgUszGPYSkmJ6C2AGxZz5UkwNpu9qdDeyGDq/gm3gmfuORnt/nQhURI
oZ/hEqWiW66dsfDe5/dxht9cwN/HMxA/+uU61+3LjS8/MSXmy4SY19q3//cj
hAxEahJot6DAx0pej72hMTJa6R5HvT5K+FmylUrWFcHTvqGIVQm0pfADgtcU
HPnRiGlq2nOvGihfavkA0Xj0g1wS1pogaUg5opRC4NZkJRBrdek9cs2KviMz
YxzycCXtA4sUoiheqNUggcy40oGFcWkV3dTN7qGaeJHmu2ND8NSm7skh1CEi
yKf83LFXaH0RhYeUIFk48btdFrxpjL86BgvbDTkuh3La8bwVjj0KoIpFcgPG
YLSJ3ybws3+2F0zRJ4dRMVGOEBeux8zGr5lKzMbhFyZHEDPTKLfShcE9AbAg
EtCnjbh1qbl0TyBzUTAFqbURR/qsoin3GI8fHC9JC9tAyxiWTM5NlyyTDtoT
b3br1H41d3M0uDb3q/1eGD6YfIxtmGQrMxbA3CLLG7fnXvMofsq2SbDmGzFA
TmUrBvxRkZX6XTrxiGI3PTd3KjR3LgYsCmBlNjOvrLYeZa0caxtLrNPV5dRp
eGLLnN4MlPvoXGWlPPF9ljz+36CU22UX/YlW+GJvLVEZgFvi5eh4SuOyBdTc
khccyfZQ52t2EOoUyNtnuKyBfMKuC/dNQx5q1DUa86jWqrj+Zg14AlkoDj/n
VfYdYjl01q7/Fx+IPAAdZAUjCFURMwmlv5K1K9WBjGrptjStSOs3P+CmEPqU
YfOh4p1JMz4BgfIsPQlHlq6nvZzQe329IAx8vy+kLDsDxWdkqsxLgJprR0r5
f3L1VC7CUcCicV1jUXtGvH/PyM7NR2393egL0UDj71kA5JSZlmlSAn6euBzH
2lUaI+dbsIxos36u2zdWuJspuNbCy4v68NHO2m3fkpcPsI9Cp0OonXkbw0PJ
f3+lg/ehbVSSds9X7dbEXrvQc/P59oJiQLMQi9v5Uq/2krFOVgute9HGgxaR
m2sc5oTI2H6UKJODJotS9eKJZkQmAjayAGy+XQPJ/RRNuWABCcZsrbWvwJgw
PEEstYw7xvwZQGzkllIueZ+SKMab+K0EmAf9WrF3jX5d8xRs+S0s5xN9Q24f
rUrV9S4wtzV4XVoURF1kkvo6H0bSOrjedTn32wyg9GMmKFceO3kDTn1GELUf
s4tgDthn709R4unW1+c29atp25m3ypQ+azPHFeG4r3YfHeWPWXznijSvDCLj
9HMmPSn6p9HwrPt9fRGzCP/tAeaUpNiTGODv6bI8h4HLp1QNQ0z+d5WDPRd3
zflk4Vwkqo8sLIksM7X0lcZ/wk76MjgPNirYyrUHslsn49wSin+ZZo7k80lk
tp5zn+Bgiyc3m0HiDgcxi1vDAWRgDiGMvZvm18eF0M7Tl2CkJfbcq2lmvs48
CwzDVjTFE2eIENHbfhsgSPF2AOK0CzdNQs4kEVE33n5xhYoRk8z8ZKosbK4p
0T5Pdh+iDjXbFA96qu7QALLgusILhE47EPlQhlYQUHuLj9S979rldaZBDqxP
d96AKrBDZSoyCYv4zMsO+iIwK5lbavQSIUaVpnSVuf65FYKwRqIgk5Jb5EKN
WcPiEHdyIa30U7Lt4DGDL70Rchy0OmPrEpTS2IcfWNdL73GMe9pb4XfRLB5J
7C5P4yt5HqkSPAmxUYsr3nDSJ+fEXuQtbKanToaO0xoFANKR1xYXyo8N5I6U
6bJypD8HSlZ0jcH23bodkWr+FyzcHNQxW6tGBOzAvYhzu7/14F0t68LlfGsQ
xwqPlAuzzmCgBwGheFEXdY7eoidTjarA9wwFojjOo9AQjjpRAvQ3E7GkfE9L
IDowGbEqIDOgGOrM0RwbIdkxMacc0kqGMVDNUt6IX3yAffskgcznt8v7LoBn
4ZdDKpu+FA22UBu/AB3x/8Ko6ICu+pnerDASBpdfgv3L1nvE1VIyQfYfCBre
GMK2Hty6S8P72wHz8ZquvQrY5jCUIPKoShGUbLFX/Cft2qCr7dz0I2sj9bAm
Xcq9NhuWs8pZ/fD60EToSmWlS4SYsKx82zZQ7PBRfdXMqflMunFOoH2L/NQE
KZZKFEeNxy99ED1oRAQQvOBPOi+zhyhx+3nYN03DtcyLi0ZA7+iDud/AwbZD
0XxY+3BHEIfHfdTG0X/Xh3xdkpW+Uzt7jJ4AKE9LRR2hXu8C/Ji9GXhEGxn5
5p+NI8ogLtsfbFfuGUD2aLHN1oEkQTESlaIKAN+Rvf9+SD4J1ZVuzK0b516k
ZwL5SLDkvwP4g0fOUNi09IDX3TaWdR8CrN0yHB+5EuWfvHaLYVnWdm4HmjY4
v9MvEgH9WViVZtT2FFW1+WgzFJCiLk3Te7+FiWiu+Z5KSbKIgtJ2YP15ZGK2
+vDxKDBIV+lHeaNxYpv/b0VAE4jrAF0dbixrLGkA/5UtDHUs7M+Rk3Mvetik
DWtjyF50CbE/RT4a+wVdLuEIbm6ZdzBP/VyPbYtbrGLaQ3mL07lV8iyR/T5Z
n56uWe02RRUKb2DkjtCKI3jI13mxAMhJ9zSSjG0QzmA14RsDrnF4m9g033dr
bLJnSd1CnIlGHE4GpQsAHZfewZcQqn34jncz/WpavwlBLhbryypdnmTTU+ov
Xp25qovrCmAWaGILNZvfeIbwg8nxvC6892FPALaFVN1xZtGqgf0taN4Lp317
MN8+S95C5RiTKOxe2pDYVqazW+AwPgLW0cmGhcKqqWoo8Q2/DugzXlhHGPLT
HmXBkJFniDdcj0wa0Og2xvwqES5WJO3oU+QVQW2Jc55EAsfJUee6tQZeElIt
M4iWo0cDLYiih5U06lbcP/98WoathHIqmc+MTPYET/jhnTxo1Cm1lHCE2LRv
npyampmI4irSycggAjBwIgNYjRBDu2G4StKK5uhrl1BSCfTbbOzeFI4wX8pS
UbfA47B2MqRO0Ysv8SXM4bNgdbtybNDqWztHCBc/z07LjpRrx8Qp7WQgrcek
H1fLqfZYgxBdBaqe5nBfXtW7N2cBIty1+M1qnCC3nnrSTkaLXjiUO5OS569n
qjla89lmQeor0gsgT0U64AStBZi6DAHa+AeAXBaMOnEuiWbmZTx6pCxDzBYn
Y8UvxnWiHAWkR+we8LVOdedANYCvQWPxeatQitvh21IW+xJV8l+dT5AeOtPu
StQ+ytC747ou2IBkvhlGA2aFkMId2co8NB737d3ECBURRUJDT6hO+WXY7kTa
Il/Sj4HuFiZEFU4O6fWwmstwZiEsohVk7HV6L1CJOubEA8ok22QazrKd2ch0
6SUzYpvOhzKVHLI0s2QhQiAC6Lzoiw28I6lj3+VCQmvLT/YkkSoDssrWpCYl
q8wzydTLeaqBuV2uOSuWUwrZNYBx0flJjmawyDrvm24jLtj8x/gNI9Q/RvCK
bcm6t8AbVOBGFhK8i+MRBC2D0D7n5L5pGXkw2P8b0afT4EmE+o96cy8Uif8t
2hXBv3Ooj4DDSAShiNNODu0ur/KfM8z0PS8gG1+qJgsXHnAuUd9x/j1CSu9l
X3JwTefnxVUS7f9EMt4mvANrQFHkD7yw6tZQ/SAvfpl8EPgXo66/rRKm2Nmc
ZfAGNPMMne21O1OYSdP8fESthu0U0R4FgLUhpo1LsPI3XB3ChTy1VYZTlwPF
8emWgNZSDfSOQ7PSm1ByiJD06mgjBPUh8dTwwUX85F1gNqj0wA6Vham68aaF
qCj7xhqFw5fea4UL29PZfI8K2zdZutNnLzrH53852glyWR1zLDCHyOPWhPMN
prYL2cnDsNjfvoKJOnaBejl3Nukqr3SC/AF1ulvfumbUTR7bXbPJ3rCNzBxz
SzcvT3bbmra9c8orQWX7RtHwPBcPrwYEgMM3qbzRX+N83ctIW/1RP4rdW7FF
GBbWGgSpn/+HBqj7JDlipM1tjUtFUhkm96n5R733sgWXBZCP1eHML5RECe8k
UYpualKf6QovJh6cVBthl1rrabr5BQkEU4toaMiCyTFsoek1DEedc5Q0kNvC
SLQPiPZ6NyorTaePWdMP+N9PcHKjru7vLoPl2So7zKUcgySeh9L6KkJoWlgk
FaosFP2Z7amdlGq1G5Hvssv9sRlfcjWhFfVWLeUbfeH6tkahpLvTCmfjZyds
x1amKIy03uFz2TeuE0xPIZ0HzS/MIxtCg2ZOsUqYvxlY9xjaw3tOz79oG3uu
s6/DBkehhdcpQ2AtWiT2tiWVzp2qXBgrgP9+9ZnUbgSMgrVl2iN5WA787L5j
QobbvdJ0p4r3wnqS5WeGd5Yxear5tlZdgtB2tVDr0foxwVkzrzIHP3OE1erB
Tt28iQU24UgomAu/Oq88aFQ5KY+oFAOBHM4IwwePJXCzkK/TYhHTCjlAtACr
3BleVs1bvsr08ZPUJYeM53QC+sYMgpJkw5HQa0yEMHInQRR01INfSdyrlEzT
np+Y8o34RaAfF9JA+fcqgWVenCwAXDQ/NlT7ZTFxmDfhyXpGBSG6VqSm2Mvg
rMRML4ZNq/HCUq8e4DV1375FXlTjMV9pekrMqVnXT7f5rzGV3ceEjw5VBXt6
bXroGP5q653I1OXIa5aobZcR36R0+u7RUOFIXqJiH9XFsfjboAg7sFtXq77G
CjMDZyVWxjA6msDrkLlDc12Wo3CYrQXO0uFMpZd/H9NPBEnotacli2D6MDZm
rPafddW3QWctvjfmJbP/Yeq6859dlHqXlYlUCGzOBjfaEaGM+IkjgO3jXa3Y
mdvjl1al37nVNPKr4iXUBWcHAamg9tj2EhpqJttgQPAkQxhsJHYcPEI3zDSg
mkvEYQ2TcRAzhrBlzEjTcNBLm7JjIwS3OwyVuunNP2Gv0H1VK2gpCD2zI8C0
C99KxWhEGbCSkeilYcsddgBg+j6jSG6Mh5YWXJOc+BO/nqdr6YCMl0KO56Ny
z4ImfHsi0GONgZQG/JqjV89U7B7ycWCH/uNswW0NYwN14cNm0O9+BWj7Oyav
tT5aT5iA9Gatp1yefO0GEvLmit7cpgv/PSJDmPiEvb9P/9Z5Sn8YMuf6UB/5
dgxcvByy/6BUvowCv1gFsYEsgdmvhL/Jud6XPFmq+jKi4c5Gdx25lAusm7vv
c7sLcCGJWI+KOrJZwWDdLe5tMCXIKg57GwJg8qXle3JGxKBPRo+wDdC01CsC
tB0JaCQ82FIjK94jwNPZan99D/5UnJcQEYMusQtwlgva9wTRk2GsPr/gloZA
V1kX5fKnt93o/OT2PmB1jbMysPq+tJKAGvZc6Q+M0llAQN8h8/7nRo6Dv4NR
AGA/RxDZ+dqG5bKtcjl2CdQeJHQnWSrq07azRq7jxsIOORT59Mejb3SQ2dY1
WL60LGhCcIqsWzjOYWgHnC2bo1rvuqtFKx5cwpWpPPA0dc/O4zCp1edQlZno
cUDTW4oyf2x53NxAVbCZdw73E8lIhI1Iak5if4C7S/UEjlDYyuxm8pEqGURm
sF/8tVQQnfpJMAXL3eA5ZEHgigPmfmqXr64Cjm24p4ya9MuSrJZreBYJrpWd
GIclXE00dsYJ+Z2aZFuGyL8R0u47xhRHXpCoo88RN5DwZhEa6OGxsUyHrbzN
mMX9XJWftaybzxMIj8I1LJryMNW8hKmYBCeB4JEf05UnwitJJlHYarAtLtBS
z3VFLhEOyH1r3L0qkWegX522MyshUgawuRX1kTaTUON7K5veA35u9a6eieFX
9Mltgdb8G1aWprZCBDdjcr1jepNy1jH6Bg6ym/yv3k7uK1tn4h5ZU7JtLU9S
c9AKnjTQH0MNIz4TwQoBRNhQUN2gThVnFf1ruDHyS/rl8Q0DITwvosD+JVZo
fsVdBPEeCsng+UA8kxpCN1YPlaMNmuyTXiQa9iDTJf5WgdHngH7hJzhaBsID
qylwBxSoS5Jk5qMLK6kjCe6UZXtT60VM7okF7DFNoDSI6TBF6xhl3/daGzgN
XFFVtafJnogOgN+2Xt4I5zICsHoC50BMkrHhx8QLoXiKkG9Xn/QD+yCbKGCc
sbuJ6FQ97XR7VYREfIeDzirZrOJbJZmOx604fzW8NaP6It61yEwtgAsgUtap
qOTvhWRz9owqHxH4XxAHC1nTUZv82IjdV9rEb/TKR6md0cFSPkIj5B4lV9En
OLrKCAowKaiKiVt4sgA/FIwCHSMdEjihciqcLvIBr26c/7iQSz7Vh10mvmb2
lJ/D4muCltbMKxYl6qaLEvTJwv7i5ZcuCymvBiUGGkeiD1wOW0yKQuOendyd
nDnLsbgvsI6JWt1gfhtoDXlwc649Agdzxv2KYc7JztDG99XCImBIJGvuY4zK
qpZD+OUHUcQ088Brz1dXubYpAZATj0eIFuCCC+xi3UgDfsaGtzwWw78rJWmx
i33dVakdmPE7uSl1nXhNYzAv2qfMWKm9I+bPv12/ayHFcQyT/2aHSxHFvpW6
gSYgpxzXyyuAYCebbt5/WIe5eikH9DLOhfyxlsQh+KpUNvZoJZ/oRpLmUdtr
tVw3ut33siEpUnvBEimGzYRRKjY+aQlqAPA8cCqySmxGR97MnJLquVggPxw0
xVwEpOzaszhqajx6c4q+8pUAA6kl4gopvpKQRFInO5vuPG0ZJVQW+7qJqSx/
+ltkmF2eBegEvmLveICmI3SOxkULkVMreDKeMqKQGOFX3RxN7whmVPZIbXhN
YT7EchtfL3sMJNQw/Cy4q7Wfgz9fkZJnzUnWWNvzWGFo9/2pjFq1i8cKyHUM
nHeNf0B8WapKWUtDKNaQtXUTbNx5ATvSZrBAmc0N4ocP8OnmFu6skhXXGNIC
bro4Vj5HDVMWujtTNz/4zj5vVmSoVn30i6tIg4qQYnwrLyHY0VkZyeLVuhXn
dC4Ejqk/2/MDFY17y22aAhVXnFVGPk3rn1wJVO2r1oeP/1cgr7EyK9FjQcCm
QOo3QnVNEXm0L5QlUjZHpzq7/kv7Mn3uNNKR2CLqAZ1KLR3LbuXKEaHekPbU
y4jpNRDhnaJsal6Q/jYo7GOwhgB2NhyG4rS6lv8AJ2TU7Q5MjnrYhJ70cBjD
ogAhNVB1Bo87WBsEHAxuxXU4JWXkoDDtVA8C8dHXvMduV4KgRLobxJXDPuBF
ahavRHhj8LACDCte6gvbXJINS+SJXX0zSWvrn0AyNqtdvlBq6vQQy1EbJH5M
hzJLYtrLLfzOK0HjzNFp715X5Z+Tyu/FYckOr8FGr4rod/uYd6vipr5rCUVv
POHfBr7QP3kTZELH0/c3/GF7q77B/ndOth2b83G809qOxswVbLB+tTc4tM94
2/DhwlJF9Ue/9Wg5U7A1zGX00y4SXeBylntxpUaVmEp8ZHviwVHRGCieayGA
MAC8j4mo7dTaMsNJbU/Mw3WTGJ5I6ZowJY4DRRSEuYDTIZk0teZQP1k1GAN4
BGkvqfrDPqOSZCUNKqh3vw2X7VLJ2M1QURDNZdxIg9+9XPSE13yVQHN6+tnv
syXevPbFJpeTmJ70tUd0tv+TJGS+Z76YH4MFtpNzcZF359drK8p3BXa5CvXD
Z+/lF8tEgneRbBTvgaHYcvE0E5rMWIdR3hVGjdQCwQCWzA2GPxOobW9AQ4hc
drJck4Prav9OcO1wHcR4nR1nHF/Kx+D/CXRJYtQ2MJTHH0VEjtcFnxor8pNM
BtynKDdW3sMKio3WFvBn2d7OmuysFMtN5Pr7oo2Gw/K0W8IoTFNUKIvcemvV
wQ+gsxibWK5tDiNlhtJgqml8OiQNueEL0/WcbW0aQB9CD6+PADoL2P1OZry9
K2+0Ia6JugQRhTNZ4/Oh06S81xzJ5z5NXXZqZUTuytOCaxMsSAlwTwntQ+K9
FXPzQHDrmQxrWTj1qJbXl8sfC0E57Jo9mMYn5vAc/6QU8VNBhnHrni5nn4R7
ZmQUaBxsweul8VGHWHtDexAnxJN2D1yUVHvrUSOFUWZbnD3VIFjD7yMxpqbZ
wtxx2jbQCgeD1YBLkx3r619VGnLqHs0k2H5TB/U+Eut4xUfULGfcfDzbT1b2
iWwBxxyxNvj4EDG9WRdEumOidvoc0hd+pU6/DDb9wkZVJ7qp+ktwTvsnFsMp
MM0bpgn4RiPFmKBNNdMJq1XI4ZiI+H1e8dOzhQAKz+cejWKqrtk+Ot6/1eE3
jC5V+txZTo1elfWgxvbYucde6lsePMHj3jC7tfiDqVcvqvppBoH+twZXpaI8
cNCtWGd+7xy1cIO332KyqVUfVUOmg4xbW64sWuhH7kOazjk1YmjB+1tYLDjv
MkaaT17HmzTnT0utUqX/QQums+NMeqJp2TmJEHzqPWP7LY5VxEGqu3NFNVyE
yjHkcjlYna+s+7D/EMA4P4f+OPZUnLUuDM/HRkWzVyAyGgZKx/syUO3yXNO+
1sknVYrWIV9itOSHvsh9tMzRzR7K6N/HMQMF6Q7+9C61KJ2O4NblHY6w4+ql
XIJ44EFWz1wrZPj05d7w6FOQuGutIPGbD166eyPrleGFmzSrsFS0PdsE50Rx
00AtoDG7lLbBmoO0Jx+Zw3KjEY1YGZyCUwhsHXosPdE8qLYlyNFzMbEnGwCp
2oo+uvjZgCQhcehuonNu8PQ5r09hdfKLCZKq90AtzTiwRNhwuVKfMgNJx9U1
/qvbsMErvW6yowlnXjC4C69FfWHJBXIX3XQHD64k1fzAf6cAl7kh6Tbl2utv
fGCMUJM3yQmuT5c2q205/9tbpPQjM4aiEnqx8jEj94ZSD9Egqfov+lWPqZeH
858KM8StjuiS4Eb/HMMqGwvG3mW7JK7mGeqJL0vO5nPvYnMUHf9gjZAZNYz5
Rx5UTrFpP+++zM27jtNvHsvNShWGrA0u6PNUajv9aLq0bRGbYyKntRtQ55tF
4XD55DnM1TFiAk3IXlPuQYaB43c2XJ33meljdPSFz9Qa/Wu9MZQxPCFVKbTX
gKGkI9HlXJLDJeHZJejrXgrqY+aC0POZQM3xXn2QmlNHvXAdJTGeXfZ6AoLH
5bIwtVHBrfSgcvIUK2QOMikmFBBfElPp8yf9bkVvZvxQrsWP4TtGTtt9ysZ/
pMHkIIN0PUDA3Hoj5t9gBRud6VV+VFBDl0B8omrnL4ueTUtvEoWSryOe85vm
ceC/2rSPPsah3bPH1nw1MhjNYjS3Cs2IJFw/mBd/2LmBvdRKyB0rN6DwMzc9
zu+QJFjVcKk9KDN2hKXiOM86d+ywwSx9qK73qGbkN2NFyIIWr4l+I2Jw1EE9
3KWy1uQRTZTxbs3vdcujdwNu3pDED/vABnndK7qbfuhbroilpUzOxcr7XlCA
3GxP0cgeO9X9qTnDKH4yLeOV08WR0H2l0ciiNPYT2HiYYzVuSbF9UNNSBmqH
ewNq9CgLM6LP6lHebCp1vLGQS8UwcBr4GcbZ/QM9pszyVybBUlDyPOCch9Dt
QiywQXpCmsAsV6zMF1z/oxyE1/+Cvk2n/iKx3aJrsKPLO6Sopc6iPS4N6xOx
7vl5uh/SDbvRm/PdxV1UraFNRpP+DjldOvSIxYaJLss6th8dTdfUKHXXBxRS
rp8eBjwtFB4AeLrZLE/nuSeAXv2vTJMNwkrDd77Q5qo+o5I0lGNrsywZvVxd
tl1pg7M1YTPdPuiceBumB1LNRrSXnJoZobde2pQOCvUB3b6l6jYb9aUrKftj
x+4HBrh2Qg4yjcsi/fUKshVPtgi92SzT8R7qh5XZcUGvkNwxLKs1uRqMSoeh
6SHvQ7Es5xxa0eGDW/xQMZn8Yzo41+48Pep0kYl7TsvctZ6seskoKzI+uxgm
Okr+hte9USkmcRj5gmE7wL+PIwXdcTYdkvFAGBeHvN7DO0Ya4QRPXvLcXda5
2Qd6Kz2YNKjt4fwAHpm8GFE2Ot1RAvjkwHxcnxETIil4GNOFWHPgyeJMjDzW
HwmCaB2PpbCxbGCRdkuLjyZVf07BrTYSamXXfmkdTz6S61AuOYIzWG1Yi61/
GGctJW0NwK5GDSwwwFix9hYQHtlhQERQop+u2S+kti+MPw/jIiiQzHkCdUmG
e2RbJzl4DjaiatjsVt++KFrZMOPxV14Hkf6aN1YFwcSJ/lwQa1zS7B2GDyea
OGZNmB1vb+EisEc0glUlOKeJm4ewRfT7iBSmBNvw3LJBDWirG+pEDxG9rEJz
ef7ae9XDle8Ydgx/HHcRzMtYcEAH7PRwJzH4ikgs9+3BeKvuRrZnQXoiLZhs
JVFvxULSyS4JVgKHsl0vpOTy/cQcB/mSMT6YkrTVrdd12DE7QAqjld/D+/qw
VnYWNCBTcz+gmOalPRXrNPexIv6tBLVfdLfWUdDco152BZw9DYrQ7Q96tVDX
Zdd4eShY+paJozYiNikjOerLXoIk2VHI5xRNG6TAjTx266y5TpuE2674pHKD
h5f13ec/e3Hhkyb8w7wtFLiwp8VQIQf/GgOnSKEF7onMc7r2P1lo4AhzNcVM
cuF/ODspAgWh9vRLrJ0ZNOBDwfWpoaQwIO67zdaup2cl870heVYlzzoBBXJd
lIBcx7+bJF8fMPnmZKKDJEUBqPAHfVOpolRkQ931N27T0xWR+7yZ3qbX0HlR
TeCw2DF/NjxZFOTK8cAM3BCmYFFSx3O0A147obecVT03qeKn3n/rMYpYWdtj
mJ9IRIU06MXLikQk3rtjle4ToR7mdi191Ie8U09HRi3GoKKMno/BwsmDAp2T
UtCWzSTQ4G9LhoNTxtMNsSThxM1JPJzkMzKCCpcOft5ZFCiV5sg9qsxKARh7
IZuzIPUxH6Zprx3Z03qGLAuNuhoS1GXJeqfeerECFjjgaktPwmKMEZI4Cei1
nh5uLJhTrdHlwAsEyi0+oeYiz3xd6dWW3N/wmEZ+TtUtFogtZ6nWFLfYUM/s
kSN0+D2bg5Q/uIzHxkWtbXSh2KzRhXViNU/AG7tJtIdq22QQHmUrjhJdg60M
OdiXje6CU39zUmSOZFR8efni9jww/o9k1dd5v33wH7kk2xQxCFJrXxIWp5JI
JVq/CNiZ1QCvV4nA3ZpVHl5fBOzLq6LZC3FeABMjSlifL7v/W2RIz5qwRHYc
4lw54tpLY3DojeKqvKo7bKfRqnqh7Bfa5g2+N0bkauSR99pSAnN2u6rgJ2Oy
KyPlHE5wXq9X0A2NCDkJfXV4WoOwANR4GVW7ZIF4OPkwUahF6P/ewBmbJ1bz
tj8Am2WShSoUinW7sQgTsf2Y0Ojh8HIWRKxy8JWG3zfQCvhWoohJ9UwIHeiv
aaETjq0lkuguVDxwsjUUo/1E4gS6fCAE34GZwogpRYEOr4wkdces3cyETlRf
hPeo9ZRd3TxyzghhRtp66hfPVg51TF50BBvZZdGusV5e8rAQQ0KXhFb/v7xO
NRgFkY541bNKGOnoNy2aMwLGkfR8EtmnVOsx852Z033I9xwoyxPV3hh2U/Y7
qP8P7bupes50cDY1zwv0PwWmkBn+FLkaZpwh7Iaey65lwijIWnhqSO65d9Ov
ow5X755rRgjJTSBTGnK5aoeztN4A4R5hwqdydPVnyZx7+h9Jr7pW8tGQHliI
MUkaFLabxYZgTuvjZOGXBfqLbGZWUzGTgLeIayaPuv0VsOpBN/emDiHbTyGD
5h4sLW9jDjCpd8cJikqOG3PtrzfC9RtEu3biuDVvlY0dbwoJo7KNcKnVY+Kt
bZ+xu4D4eZiKQ+5mvywPIrv8G1VsjYk23Ijv1NRqyEoe26js5BGv7MaumjFk
/JekOmn8hnTa7buWjDgbeWnziyQ4bTM4uScyFSU933H8kpw6vU5t2J/JGaPe
81LqkCy8u15t9WjzZ8rnqfaqP/bq0td5xDTyzafdV+mHxzgzZTfdivCWN3zN
N2fq8b0FDx/hDvq7Kjx+tlsfDNA7zqRUYHL2ETRux7RjvIIcuD3qoVJs4oTk
OvbBoAUIdx+sBiD/mtGJ8qivTOashV9X+UvYiWUwP6yG4TqXXit0KyM909rQ
72l2Wtai3H7HmHSoARLMyrtFh0dv2EWuzwQ6B7Bu39ftFlp9TWO+5mG+8+dW
RfbzM9Lng598h9GZJBD6EnZsb7g2SbPnIgm5YXVdrtlGs8jRaFClomwhKpNU
K47epA6W4tMwj/b2f6q5nCrlKi72X9ge0EoBJsAJIxtOLQdbhnXSTFIW08V/
0sBo59tCsGQolZ60cDiwMXQcsvhLTjYjHOiGrqLZ5zhunozeYuAS9lz8l0X3
YHPZ4ZfM8h+o7fVbTfYFuaJg0oANNxpc55SmUVA0eUYzNyJ8c4tKM4yieVSA
5YIh8oeaOSPBdirNH5gjaVVzM1617pEp22ZCh6R6AMHsUGngxaMRLZH/H/kI
pDMry276GkVo/4bAVR4OsigBx+u0R4S4MWbEaxSwH1vF0+vuQe05TLbefUbJ
aeKjnk8v/KxMy48fnPuxvr/bTzJ77o6+CDcEn7Wvy9Vp4fJld4JpDaUsZ3Ob
wxGbou60y56tkFD3EwtR5YBZ7FOgMvA1fN4psNu2F4g5721IyU1a5iVOzTQ4
9jWJ28ptr5Ibw4Aojkok3cBTxlDpOqKB88zfDcKkIEggLxElNfdmCzpYQO+X
RmjJfAbGp8WolxHGEr4GohQDLkYwPsJYw0YgY266IpivwIv0x0lR95mr9dOJ
3IsofSvWCQqwlB40Cb7aW2hYc9yaYfbzICSWGPCA6iTZWpt1U1eSr7DoFwJN
Wi7T56JLaPSCXz6mGBf3k0wz58+pHkoAM30/I9QEg9UQZo/F830nhoKXxlkW
I4Xa4vL51Mmpkx8sQe6DAMMhptxBDbdByM6RHnnBTPITw3Y9mdSIXB9S5vaM
BF1599uzkReYdhWKoIvlR93SxPHfiRpcyBmUBoFz1NpRTIbZF+gXJXQyuf8H
qCPJdImsLCftXhbbFzug0A49gJtSG3qD9GFHy7F8SDhZdoCkDqAErm3RnJ4C
iA6qeCa9lfHtrjC7J2llsWcvtQwoGU4lm5yl6FwU/yWE1BPZFwrHr7a26qZf
UWMTEr6cfic1wcK3THiKyuMkdtXmc8hlSilh0gdNlKi8mCwc0LrQWX5INmhz
8fvQlc55GQ5WbSrZcznucDI47h2ZYQDau9LAEzGxObk+QeuLm0fC/d2Y/avh
1jHdwDx6LrXU5oiUG72YoItnG5OLqjSArF4QNieVCIZmGTydgcs893Pe98d/
ahiGNqZpCd6L47qlNo0ofcThHWJor/B1oJ7gNwpfO2fChlrTw6QgKpPf2n3D
GZpVVePJZbMXcWD0INvVG0knDNDsLZAdH+oFaKFa4GeVH0GS0IOh58PQ8BS8
grvE/GAtexVxzQnxnpUFObixkAHQNHesZxTkES+x8FnquxIZLDocO5YONz8K
iDnFOIkhhzChb8R6nw6ltxCfUscIGYmTiFEDqKU7kCeS2JPRUPTIrMKqr6eq
iu68op9eSSy7Ipd9lKhYpBw6Ixbu1i8kTayD3dfciksCsqAhVU5xD4wzRLFy
9ZvsbzKqWWVXsbZzmR8ecqKWMh4nEd+KimpYs6vPjGNJbfi8cx/IezDAFeNf
8GdQS8zN7yOOcXiVz0Ym6XQE5PsWwI9A/9gC39ZoFj3Ifx73gXqNKlVUFVYy
/5tcwXaST/DKlfzNUqpXZTq5VZaqPTGrTZSCiRi5tbDG/T4eeoekK8TUxpfU
PgVyTp7expIY4Y2TZ6Hi0OHY3bNeUc8TUtgvHit1TcwA672zluU36TPmZ1GK
zlnnP0BMbon62Yfy9jrlzMPXbv8wO3P5N88eP/i6WhbZ8cqq00ecVCmlyJEw
nWUzTa9SUVQ8kbyQ1nq1vBZNgeTo8r7xbsGJ5gDgOjVSybcSHxRdA1t1mAX2
oYNVGVKiQk562KtSYktBxkYWgkc7lMxKgU2B3/8vtxdsm2Y+sdIZkDcVb4SA
ilwVN+EBoETYYgZR25djATh3mMVhFLhbmiewrxRmN50St44V9VpaMVVwjDLv
HT8IiZpmW+RkjLtmnupzK7SylSRG+esQ/wgIiSSmIotupvHJ1QH49YRgPIax
udkO0GoEyuioQdbHS9rwIWBKdYl8SRNQMwTT/OR7l7k/A3MYLPlsFohVlijz
tm9LQ9fB72jbvZZ6RnnSmkweiLoWvojEPbudWwMJXnhe7LwMsxO/aGbkrKzq
xzPpxmPjSL/Hx/DAaT6aMuRyTDavpxf+DhckWDTZUPu5dzCeGawmyNw2njwP
oVBpXNNAgiKdUN0dnmLk/jbP2FEL9+c+Hj//6u3UCdOYkcuIe6tpV/HPe6SP
lAY2I283rQOxJbRG88aIAQfwTMIuqh4/72PCmv+FlmAy0D0c9SVzAGcYgNY1
5jFLcB719x8uub3xC/43+VXgkPZe23sK9F6HuKKXAoyG+4KIF7Se2nyjgiMy
nvvu+OwpgVKqzQIi7IyIggMvHJExuN2MCnigx5TDEraxmuzrcuFgd/A2DwD4
K7xVupgdkQR/gTn96Tmqc3BrjeLrvvOErl64hitLaTE59IX7rBbztd5Cx3B8
MHjM+TRcWuoulxMuEjeqJPxw8EelkxDp58fmUGvIGyTqBKGFW9/ixZohqi4I
v7vas9tjfwvK9b3/j8QaGOeDZcBnnmQiF5Nzf+XRwKfRADoIxq/ofrvBFj7H
ftevURJkMNXdG6vtKL0ayCG3fcYCwaFGs7Wc6u+6z85WxzPvOrt/CJTv3yuH
l3riYaIxH/heTwtaUPsV8RgSaraV6GOGX8uckfJmteJmt9hhoqlG2EbicL8R
HV1T25djjLygG/OydwpRCI5cHQECpL+cJzcYH6AFAjADsdOofOHNzNoKiTYR
Ci6ER/Vlwad/vxceSdG170BiGWrrohWi3bru1qMmLyVJjrqiBT0uUE03xQBJ
SvdLjXSuzJHEkvX4bp2n4f5i4Qnwjfwloki+xQyWjUqd/Ci/3LddE557vY/q
S+DAPZ51IaiB+dGNChcxHbA1t/rqy7/2lMUvSmAh1W0GqNAQ8G5nKF8xcBjE
WAPaJi7A9JglBQxadvhO6jNpQzmsNQqjq4tfEVU1G0W+aibxm4jV9KOex+ND
i+sHRD7bb/xETKlqJ7opGcv/cyGzSGQFwV7Xm/LGtvv125c4jAm3ok4+abuf
/dIa2BZwVOYzLyorMaHiQZqfQWCJ56kcdNQrDEZlkd9ojgekaJ10abNZMhXp
lalaCR2GrXMzOFlxj3I/STrLIIpOf3L9NVjMLtKd6mKgFYlflDx8Uos/8Y5Q
SS/hKCKSPhEJBOt72pJQZuGliVjgqnU6oq9KnCVznRjD2yEF6h/LMsdeZ5AF
sw0fbN06XOZr142ud2jO+XjSoZ7dh8qY/aa6KIVmrRjJswGj8ZLscHWH9h7d
tNFczXsZaZcKClXyuad3XBbu7Ui4qzlxeEVwB/xsV5FDcp1RGQJasiwo909q
3QdJeyW8rUpL9tR8mnsxv5hJCLo3zUW40PAsyv/HrsRV290CDrVhsVNH5l62
1khzmi0s91LhJd8qNUo8HlLSXK+R3uUxOvchAaJy+5l9Gxm3GPW4N3JJ5fWY
H4dcgM2Hr4r8AFP2s7aVmM0vKV1A5TZ7KzdWxCTtc22bHisKw7uXDTCErV0n
zILBBEveU2FpKafmIEGgMY0MgPmaQprORGkb7BkVetN+40ih6NbCKf1bKfwh
nPMwtLHugj7AhBzF8EGXY4vQ+n/BfWkdwFBa8/+fQ/Uar2knRcphboCHrDwu
zAB5Bd/AG2bxifI4/u3iPFJb/C/oGefN5w5QaHX+Wq/zD9eOw6HsYPg1S2HH
mNq5S9QphiDx0WoEa0tTFUPdZtof7oznAcpVoAEUnY0ZXSAsG8+NtHYS+zmZ
qj3ZpP8jhqA+2MhT6LOKxw7qQvISpZZuIFSPvQxCzg1z4HRCsFqD+Ugjl5SH
yiknws1b22snchCDPo2Pu3TqXprwFYJgoI5bUuw/w7K6NBgGG73vtKDFXWPI
kFxGgumxi+ZQsqlzUdVdJBA0RRlP6d4wKgocNLuFpwZ0N3Cm6Y5GVUWey2Re
vzUU7vviZRzyxzmuQlmTpYI6hFNR3d3I/vkWAickpbknfb87POB8CggTC6TJ
o1d8sIyi1TFLF9XuQQ554rkvzLy8y6Toux1S2kZbOoIIeDF5Z+Eo99977OwY
UMA3T2oEYKyIq9a/x11kBsbwzX6/vCieG+/gcM4hmnIbu3jBU1z2EYgyORdI
DIFyS9pNzqQhOoK2szqTNDTx4DEvAJjFySbZQA+Z9dsC5CMc2+2kYV2Aw24P
B83lLu6g4lxwcB50m3i5zdUlhgwBNMRH0M4x47vurf9R+QpZJlJdb4guDh5B
C4MMQW5TH8szls8GucsQugGX8f4x9WOnncJCQlbF8e/DQFBEDwUJM/82OjS7
Vwi+bbbMXLgYKJcFnHeYZ1+vwXFesvoXEXTiO2iNdgDMXlXiK5RQ0r6Tw/2/
P67BRfjWVaZja7VVP3AmXlu/yr2doER20rMgMrIaJR9pm/RDutimggrpowti
yCB5RWPxlVSKqQm48z+3HvDaqr/wyNZvH1ec2ySW1BnpAiCqTuvCmR30xi4q
oVDBZyEhvR3GmmUeeXdVLOM5Laxd8Lcuuwkb6ISnciVJ56m5SHUuWeCHVZRV
HT1VEz8xjbtNjtU5JtoXkPnngnvxRk5yqiRzVHMOoV1vIR4++023YC15Vtyx
38njT4o74TiSLn+u+xy32j5XRtGm6zod+cGzNs7u4B55wzBdbwhJccyzq6x0
YGJNNMvrQnbSmYOrXU0nFnD6VsJDTn6fe4CB5FJEqCyEGEVDjXTtxRGixSe5
gpWrdZZCt047qH2RwNE6CGfxeCaBGFYH6PAjjZo24SWSrXeorK20cextOD4e
Oi9wAz9wCaw+yaezAi3bsrG1I9I2cEhXhNcEEaeBpDdG6hM6Y7hvLBDnaxI3
NzeRs+z7PKlr59nLSbCv4ubsei/iBcZAu5tIX0ygY+f+qIf1L9Jf0Ggfeims
SlvZScDoCGJhC9Yy+ECBIMgk2+sXKhyx47VMbVMetSp4QGkSfL5LZEWhpf4m
pnyr4Mvy5QxSjLMaL6QtSf+m/JSn58SAFQ0xrH9I5AiC3iWjnrmmugixOvAa
fIijeprunjOBzochI1AU+jrUs1mH1f0rGSuVt43NOPjL9v3T3/rnLv/IiC23
gJy3ZUw3kFio+sx8eN8Cc8kYqnutCFnQi2QYBFenaO9I0EcEvOyuO8gT9XYY
K6fnf14jphmevtTn09dYO4AkCLc1OYzcy4RUP+iXakLcRSXdC9IWnFFQqrjE
CkUu773220RctlfRGkxX5L/8HMlsGSmr8c9Gm8sW3zADQdvZBcRLDJnuAtCD
Nqv+hh7+FXpHg6TQDNspEM/uaXcDPSHX0mgYhwoE2Ao2jhmSCwgUQP1g3/Y6
aJLOwInAcXp4NFRprOnLPytNqlK+zjKspJpsWwSM6K/lN2fMLgDFMWlyB0RB
CR6y8wFako2iUCUSbgioHN2Zu7s3kPuLdUoRyWioDn6ne0evozDiswPG0vm/
xVTJv/S0Dcb/Hah2TOoBX5Heg6uGkCJVZRk0HxUngfo+jg4S7f4juppvC6rt
9E4FmbM35m9N7omCVMgO85FEyQIdz2NAMtU2zlpZ9iAnUREMi9iT3zABdx34
M+FfTZMt0OQtre0CtA487LyEdg0LLQgQsVMjffQ905iTIVth3saBV0OJA6Ns
QrIThnZzhWOpOKQNbfxtFhyVpRBW2uigBbWSI8YnCUZ+qdwW4fcuwX+fyPBT
K75XWUUnIcNlA4V/z1rKl6+LRnCrBpqIhozoQQJ3mMqtA6bAqsO+QrJ9ddDL
nGWsbmBZmOEDOE2baVYQHAwCEXTvPFncCI7NU9aWNt29XGM0264H3ebbdJoI
MvA7QV/t4YOFXd5FPYmCi8opMiPKIR/KnO+pUHZNm4rgoy7k72tlDFZKhOJu
npEvm22RkBbJC+nYn7AzuG4xKhFtYe0KRG7kK23y2FsYuJ9f9SSTu+YeEgPq
Y7/0CzgeEiyLERGM7PBo8dOx1g10Yd1kj+3m8mhnFSeBwTQC3KjIwiytgCpd
dFKsbRnus17CwluHwuksaTJjljm6BTG2pdjfsuJr/sITXL1lXtbiy+1zXcq2
jmhHavXN1rMyImtEfBNC1oCIqUyVLm8QsJA3n40BldfAcqjZNwRk565sNNmX
lzJYTF/B6nPzSLlB8PeaBJFtwD9DtVOqVqerYl/8xsskxrjkRvsfyvIwLpYl
TXklYLybfPd7oJx3gBiI9Q5nd6onuzQsSyeitImyyI5K8mqhAMbQss92QP6r
NFRKBEa0uNU2bGMmTc9oyJ8h/lqiTgjrx9FCK0tjgwddufQWCMldPgMBtTOt
lr+zHh3K9beo+jALv/OHDqUS7I+FmB924LRoEva2O87/s+SuvrmKr5kqe2c6
bQR1e9kigAcpKUEoZDjaS5myl5ReFvgPADFh4bmUXA30/GLFjFNwZPXwCk0x
tAG9RDGw9OV6Zg3Qnw7g7J9ScNCSAk2/pcbzS6Yq/Ub4HjsoDlfIKR/yFH08
rr4JXrd/lW7PuXTR4s+k6Ts0URw7Ib7PMR3jeGwVVcH1pmFyAmMChakZC994
g2r85raABXfo2sxLIf9UD+E1yUfIAkdIs1itTN8bsXMbNZ4v5CkXqQdGKZTQ
8kWpUD8bKvZsoNFx+8woR48/LfaIKDHXjqQPVkDtZEFzaljXAixxoz3UgVZ0
YWexRZv/RNYlke16DPBfW0oicL1bnML61votAcvA0G22LZziFVIiB9JgdG8Z
aq2C4d/RT76HTElYrSERo/sy2/hCR9EAtBMs2uoGtHlOaoUmBhTCZmazCzbd
EbJ8aOOzbVkYvZxCGXwqyv+9VBUvQHAUdZ/zVgffI4DprP9Rk0qM0AeDy7bu
Pkx7jRrpaOA111UXhuTmoC3epvZ54glRH8n0vJqb7ncQufqvnyY+MoNtqVkx
59WpOB7mokc4DvcNzu8HTBSj4b73KdV5NTju5D2yC9QK7ZfttVIxkg0auznz
A5/gGLmSeh0d+YpTc5+d7f6KUuHOGM/DTtCWLQIXagY/4oP7WRAIX6oHnyC6
xM7kxWWTOvNq9oHNuh4sRa/deiNhivLjDO7AncsPf2EPX4VHlDaIdsOrSKMm
8xxynrcXoCcl6/IvyokX0uSXBT9LS/K3vt9Xt15fZMD9XFPP4b4+4o9jmphZ
wU1kjWpjUiMYjW7syFdMrx4j2hmzszjLyeCETbB1atOSJVN0B8BuB/BcBl1c
cpaISe5uUDqyZ3p36aaVO9EtmTDBjr3LpofdXWlCc2O3AvSmKVVD4AFctKeU
eworKhMUOc1YEVN4ptLlEx6P9V7mYuk8PIGYKSg+x+0TOj1nUP4v/0EdbNWM
oqv2ZZLtwvWE4ftMUu5nQWNdwwGCxYw7Omc4+A65w1XPz8dgZsmqnXP3a0uE
GO7zW6UoKkZlOAqjqDsKwTMGO6iw4hJi9Nihd1dRwfICEvpyd8LZNC1KgQGK
qNNX9MKe/1nkphnMy7rn3f+oAQ7PLmY+SCfFAgtkGW/ZXJ5SGkpH32SHzStu
/ianBH0UIv2bEiYfx2/hQBTY4+DutwV+wNJ2A2vETFli67WLdQA7fp+D13Fr
iUokURYDmkleDBPGr0J0Z/lVtyMTxQsyyCubrwxdNgPcWqV7PpLwEEEUKqqw
o+FalPG2XR50GAQ3wiOobzgRFx/65uv7HWu0E3Sg8U4qGB2qyvu9MFrKhPJV
uwQPxodJJqpG/nIn+roiIkcAMbAt1tL4bR+pbUrfFtI5PEnhRbNxH3gMu0uh
d9DYoXh5MNVsllWp3klPmr2OinBfpocb2EkaQJyrO0W6qZ05gIwwQOhzjbkJ
i2NdbuIbg+miqNkkgqRv2fxdJzRogw7MtBEjGONwzTYmCUeIOSlBHejn42gF
uGeRHefJGpPlBZIx6cU3O//xNEokpPk380IG7QNit7q5jI9r/CwrAJ4vzT7Z
cs885jr9FuqW/8qBbE/nokAsoyWk6cHW3LlpeBWoMHfriFUGG4biE7z6mJAN
90oKuKttzSa5mP9AV77+O6wV5Tec+rXaLS4p4gLrbkUuJB4+m6NbMTTvLjnq
bGCwmrrhlNc/bpry8NDGG2P7uRGGLORY5VxCe+ahhoQZzjfyls6F5wpK1Rqd
BikGK+hiJy5jrdeZWB4n1bSNt9JnuMYh8qpGTW5ugaCXAPhlzrgVK7a+WAYE
oCwQO8eaMqwwoczsHgGO03k6NtoRUIIuoJTs+PF5txzIsYhBP57LbXnBPFyk
JjFQmfyia5z6JgMZWi2HMJNguoo4n6sqIeWmG+rEOjVSzU2UCTo8vGfP3wKm
/4TuakZaYV4SFETrRVwbvTaeE0QoBZOSSqMskIOVfXRMomjEMMo4NihOK83e
X/qpCobhZK/P7rmtm3GyvhpJXOy1cb9UwuuVtAsstn7O59akN64ykpqQjsvn
m7OhNWpK7370ANINouNulUnLiq3qsVvRHINm/ya6DZTutWl2ViSsIIRbZXsG
GQJm5QSXyR7TNGB3Qt8GRK2fbgKzvykm+Bz+l4za0fkEEshvtBfZySRUmY43
6fYk1tOLs2MsBhOF0A3DBUTpx+7hsN7H74gyAmHToHdZeXMmERCPWQ+7BfGe
IhyBPUBSOOphc42flp0/2mIFQjQwfqSITOM6abFhhAfsCE5UI2Vi8WdxFifl
8e0cDN/cRtm4QbunSWzJu2tBa3+x8hMegjmcvqz2pfvGdu53tAdZ0ZeBimIm
/VQK9qyONHbCOTGNJ+3X1D2KRIqn70RuhB0AX4oFhc2o0epmFK+0ud/v7Kw1
6MAMScsrm91APpZA7ZlH/a268bFCSe1V1clZW63Dp2JrV6vW/Ja/5fUDyVri
jTv2WJxbBA4/KbTKezMvZjNDUMDxlcNE5BvjPPavKM7J3Kulr3fiOlCwk9Yt
1SDtnmHeZK8XSbuOpMEuFl4qWr8UGPu0/G8kwczfF/Geznegp/oK/XfKGjHh
Nnu0ywPI1sg2JI4sjfyderOnasr1rob4Tgy4t7ybFcLYsPMEZAeG3FU31GAN
LxbHuFbF2rlA0qRBruF5/UtwQt90K2Pa+XK32kldpf9zRJtz/JjAA35V8dGC
QVXhA0hDhMf63rxw9mlLJEeEOPtNbyITjBVNQBIXlU9Q0ftGgeKHffXsm/P6
v2n5ImvbHtfpf5Ajc585E8Y7ZLIq1frDy1tjLskBRkHSIcAdFSw2wxIMawlU
6vKma0KM0fEMsZJsoQ+WOdtME0Ygv/a5mdE/FnEoCHP6S3Sdar0U2rSQTfz+
IYlYo8YXiVqE1qXorEx24NlK4LLFVTMi918BFGn5tkD+FZGxSJVMnXeGI6Ew
ol/5hEgo6ib7fmXnjgbrOlQjnsPPnC1KS/69GnkZ1G3rbq8yaT3a20oLoAzv
gLfJhYQSycp2aMv3TvjF3bSDSE14jALb23QMlbOiXSSw0/DPW2cLeqe1h6u5
X8ZD5Fa3QJH8VrijwubBArUa3ZHNHcL4RaBcY5X4yEuEKHsnrpPUPHEv5Pli
OWOrkQlqkBbBIqpVch/2L8ebQh9Tj/X6bVY9wd2Y5BV6gniebtcJeHloy2IO
TVsvBss4BGKRhGwmHL7i4WoXDjXnrHDZ2qzRw4d0OnJZom5GvO8wD7lXUYdc
Z0oLerCaAPitiG5UwdvkihezmTnCSKT3YYS28ftNVu5R8BJgEbFpkpQH7Vx6
4x+l4Edbl5Lid126RC0WGCMMy707UKmTWSTj+b+hE+BRXi0Id34NHCWu0q7V
I2mOF27r+/dca84u3eUFi8nDZvDthHagPlA1p+dWLj6rAo/1SrP0yuCfuQ3e
qsIVaCmtKf9wTYdEIYxd7CPi40/CD1vr1B7nlHqIQAVZU79Zhl9TZnY+eIId
V/yrorSSGsEWzWa12D8OMCB+ILfdI8BPNf7ZGIfyJUWHYCXSZ9KslS1RGTBv
Fc/+xWHT1K1xW40y0zVEt8c1gQRzww1Oi3T0YK3A+kk+rDblvifdRkfL2NaG
amYqsxeqRLikr/DCl1f7F072S1znrmdk7yetwZDAhhx5cD54ECr2RebaxUMF
owti6b+ihMpjxwqEhgrC04MTES0jyD0t1jRjs0QmlinXkeBUjM9A3jeRELtv
i34VUQvGYtV7R7ozEeENtz2iVsGvu9/FhomChS0vCYF1j+lomyoCdJqH+wm2
+xKx5N377oKMq70bPaPYnw6sn7atvVdbCiUxrzeJ2YLvSosQ4ZegxxP21YZQ
TqdHmg906NkPIDWfQ0tz6kuVPIW+6hHk2AS+imsxDE9o3CEv8Enx4je/YuGs
Ha+hUfo8DZwrdykL9fmeFxLhHpCvuvh8Kq7vgh84bJsRxyY1RNGT8dcVVGOQ
Qw6D6Qy02ESVOVuehFNyqxfQreH9QjR2aBHKFFVOioMNbsseLuD2IwiYNm5S
pXC8/VeLKPSUzQvKm7hGu8mJl/e6d2F3DbnCEW8fZ38Kl0jjF3S0NWUgwqE3
2i1b5KM7eGajxcnBJhKNvdMk4fkSEchMwZ9IORQJTHbkPtE3h1i8w91k1q4Z
JZd+PpHHXQ9aMnR7PjAkVZD/HbkRgNIPjr96oRB+dEcmE9e2IQbeWjCMClvv
b0T8ocEBfr3mtyY/hWAQ0CoaZSBVcQeeOJyBlrILY12C12f4GMHMgPks+Gv4
ziQ3cBEYrOwLRjZ8APA/wv+cNG8nITQrjRAkbWSCf1JNL+jlUAxUoEGeby0L
+kGE3EyHShpQ3w56VvwuHX/ImZPsFnnQze3RXvRbyUSi6TKA6h8CEm3NG000
S4L4RwLw4qtM5zlgAabFb7qq3ZmzWaJmwIVimD2bur3a5JCOeRuook80xYXz
2yMOXr/lpE5BcNKv5Tzkjvm08ZqbsaA95pdd0O+0Lf339dpoLpDy8sFVCWtA
jMm9UaFwJ3Gb2rTGD5SEG0W/fZ8Vqh/J2Pq5et2yRfuRye8/bd4pz9wwUpYW
Hm5splBOIoqmxT35Od+my006Q71nxzxoX3KteskCQl5+S2RaRYar6Ben+DC6
dPQzUQ8n0tQd0wG1ngU3IqubihHdwFIH5oDbczAy77RdQLWYk1YtzrZkzGye
JBBt47lnQmR7tGP0jLGovBMfpX2Ddk7CNi4tyLNKe8tJccggHQZtAultdvWb
etn+BoMNMEksZBSJMh2G5jKEpI7sANVaK41HKhdQ4SVkoy0vuZ1QzK5LMsDu
H7RNvmEsky7wbVM3x7yTxEQs6/hGUVCIxx9yMDK4JTITCqkjYjsnrO2GRLl/
/aD27mDpFBKgv8xOZgPju8nhDn3lCO4cqzfSYcwZYkXBGE10ZEcUbdGvZJbD
K6zEk4rRvTV0ivjfN+dblPNjSsWCmjJaBwKf+lsdXhb41FBDRTIdOBgZGMM9
B3l32VOlL0RI1W62hwIZzniQVNPBQVvu55gPjZAdr58u3tI6S87uxa/Hl5dm
dWHwPDBeflml/A+Ib9jQOkdQYn+aAK3c0M2HiHAr1ebXXUGrsZLmXYRTmFk3
KRUZt2e67OterYK2G8Dh4bmXKXM/Xg+FIITEwUm8F89OTYWG3XP+1x/h53nW
8kYm/w5f42ce8sSkFNXeeM1O048Pc/DXJS9fNrGVJ4hvIgvdLKAUyG5Kdvyo
NC2eNJi/HRaaKPlpwNuqvclGG3Tur4Csb8Px/V0QBlJE4OcK4BchROk9japB
1zkfHH3envmoRvv3kzE2gHtXD1l8ySpvxsTChTEBdnp4NwjaUkCNDHwBxVZ8
NVOs+/BP3w+VokwStMkOR+swp0Cal6dtYKkxe08wSGfMFH4HjSDHFfEM32w/
OldLWdrPLEPwhCwP/22hvI5j9HBgnxjRixZ5MMMCCEsoJFjibGu+Ui4DF2+j
DoIDzE6lbYfb+cybxb9LUhUfTEQiuTa7iTdEs4mCOdfwHkZFvMrflDpEr7mp
gO6VbqSGzX/M9siI/gpxQ0oLihAalbNv7+knXyh1J35DoHchlB0hIR0zK0vQ
UfNBtLxMdfE2kpAelgq5/ZbWcf6HRSR6SMUD2PzXsdstyyv1d8P8Uhr6WOqN
AdRHGaZJ4Z43k1AfnL9QgWUGlysZiUkSTeIbYeQwRWYmBDyhifS0QF1oamTr
WhivSIYb9V9RLStruUZ5ogt5FbTEE4ehiOUUDlAI/iqaLATNW1UWeHOjIVnb
PgLBSG31Dxg0Xz6fOXAljsKRRE2727qV2kg3/Z+V5vALU4nMeYE2GPyQgZlq
Aol9MRFYiu5VreMdx2/dC3XsZQY9DARkR8OL0kAAr3ocRYmXZgwWIfalSPd0
MJug7tcbDlBTTMDBYSJHVA4PGCAEUy5GWV4P6S88KglVg4pWSgfHGdEXTFl7
clwwLWzJScjmi+EWSX7KQ8zfgK7s8DU7HGG/Jz1iRe4gLtOPkd8mMpFC+7kG
O41u0fwzfXyX+9558FV/36H8b8tr6dFKxpMsWw2IPfk5G20ZiXB2ExDy6q38
Cyhl2pOFSyCBgILVtkZ5CdeUS7iUpO5U4RFgh7HGZGanIUqlP2VmGDtBXRxn
DZNl2e+tcLEgouLjWhdjw8ioQvn/q46qq4996O5ekBjgiW/LaIYv2VQjSTJW
YenW0dHQx22njOz1vVE8P59uy0b0fC4TStCtNKWkjG8mhwX46AbaW0ZYb5Ul
DgxUxWeIJYKSQpZysXkvYfBM5h54QO/geVLVG5AyQIMSqcz1ORo7ad5dhF6r
azqVnJLq3a0jEDch2iWEVIui9i1E14eHNGSwnQs34CcHIDfLaT2DJZVZ5ozU
+xNC9/skwK7G0XQaJC1niZm4Io4HfpkDXzq9JthUcfxXVG2lnO6Jlsd8OFIn
mDeLCWkWqsl0xOlv1MxrUo298G5gurS5ll2zC096pHOdqgQmZLPF4iFy9Bxw
tdnIvTODA9Q5Jtn45JuKJ1ZO0MEWeHp76a69Nct2TXc52C7MXqhr9H3/22RF
JmVfEEkAjykYLtDhB0SVhmYn8y3tIko90WtzCPls8GMWVxCZOb8IkF3cA85Y
98jxN4r1sj8FWxWHNywqXf649dIdOQEOUTWryTdQYQiGRvg+xIdqxowMZp9k
17t/z90BKr4hdjjJRznsYdEV/kMy9JCvo5s+ke2NFEcjX5FODhYiurSoMteC
WOszwvbEyAkxwIcSYidHOYngdSNyp32wqn6gvdZU7P65dBqrg3zKIH2e7pa/
puLDKNwLrtmveCqoQnqy/uGP6nTtv8nZzGWj3qEcFglPKoh2FBbdY1T19wJ3
DccqECt23WjX9Ei/s6397hyt29//ky2LQIESAKqU3no3p6w6yeaUQzF56g9R
q0Zw8cgwj/psnqCQGZQ+xf0A8e8TcpmD9SUSO5WyUxCrPn5zCs0I9HssKlJO
6UZMF/tvA4RU2jZMp8lYm8Gi0z8vvyESpP+mrrHyecQ1ngxH6RPufJU1eNwa
cdeab/ha/GhEuAlOUQ5DEt+ZVH2Q2Hu8wkgLtzBqj44GYMsIjCPaywKjoWso
3RDGg9wl+Ub/Mp/XLT1JoyOdnVh4iOFNLEhpFcTiZFuR8IaTuh98NrfGxNUb
qlzAjumhnqvukz7YKeXfoq810aRMlv9ZwLgPKaMLU17lcrOYsE66rA9+IFyS
ShVzRnmQh9Gcy13TVD5md3eg5d1jHlKyF5F6fkwpwyXTfjxrqymOCL5/wkzc
G80VThGw6YuH/gNc/CeHwZS9gwDDeRFuYBTT5ZCEDiUiMjGanKUyIA99cpex
tyvSVBWVz+Rq5j1CnTSHS+qdvsKzyO96VrHhgjHP/ytT7QKHlSxU0VGqblL7
TVUzdyAMDpE0DIYEIdkGzrDLYzTQa+CSTCXePDLprDG+j+WBiWL/u8t9+C+E
YKcRXkEcsTDYF/dVZR88zzcJWqu4T2LSVy7SXTIRMyqT12sz++ygBqOxaP31
Z4PKzadb62dPfPSuZdYDphL+OsWrlESruztMqZFl8qkb19M7d1CP0iM6K4TG
spNbjVcSFAaw621L39p7Y06/nQX/DCOmaGLlOfhYMzizDedtjaySC92atXuf
xSovIVg7IWlJdqzd2NCd9CzKlGI4XVXmCPw38I4g87818AoI9jg0+5HXYEmR
kY4+TYcDWhf8w/UcrCP4KcVwte7KSius30Dg4jzU2NxC7J4onaXN2TOhBmUj
mC0vUvJhe/mxG+fhXF+GhF/UM3NKSzvTshwue/Of81OkWdSWKmtNr2Et35Rq
TF8RN1QT3Fz/1IEPP8X/TrOhVsjh/1Tgs3WXK0+aaDRY8q8E/H2d4dA+KRHx
yHxpGpyW6Px8BTVLIdSciNi3JWJeoV52hMAhLlYbJBFrKOc+gQn3rmjMEZ/j
qd2gQhw8Ptg2TmaGrqMX3mIwTBSfCg9YkPkAUw8Lk1I3cn+6n7h41CLBnvNZ
G3wvmpWzZ6de72VD2CVR45Ws/njtYcvAcjZ79MK4e6uTWby2l1pCO1Ud9Xto
7tB5lYYmPEVRjcJQ8KqtQ96VucNDe6PiABI48EDAhOWPr2O9QQLM5PUEsVfw
GB20SzVaFL1pUU8PXIsueE1Hh3tzD3Ns58Bssa0rKKZar8yfexlm0psIeYfq
pT060AusXY7CsyZendyTBznULbJ9y5UGYoYAdmroMkFSWoD3UcTx1ZyBbLKe
utelKIhqLLaW10HCOi6RRG8ah8wKIfJKVz5+EwDnfsligVacEbtKHBOsRrVU
RwNMrAVnM1Bx2ca3uIMq0RRTeebwuPr/f8/3cRbrgBEqT/7EwfYmUu1OBQ6Q
+jaAbB18bM+fR8Fvfg1LuNuW3LcDGi+Sgp+SOsO971ZYDWirxRRL07mmu/7M
snx0lt1jrchGG6r8L7fFz0YpTx5XcbDUpyu/8piYIxaM0pmSNCaSPrJWTa3K
qYi8NwXjoOixgywllgy4m8F9yNFyJ8eBGUbKuEsN2y+uhUUHS/uWfybX6KPX
ZhHSNDIs15rOBGTT45hdHP0EviAAV/WCbpAgz72Y5E6FNLM6GnDOEdOYrMy2
6IYdbx4gcMoUY6rnb9CPTVBPXTOHNpXTRARRC1MxGUa9d7dzo9WGWg4RIrAP
kzDHrNm2NJ8HZwWlFHGNirgAzpyO+4qImxCEmV8F7lJvs3Q1V+MBmVdhipys
Q82o5pG51gpJCAdQOwjxQLHJ0dg7Ln4dVg/R1n4IDnN5fzf6vjsl8iRCxfyH
qS4QsUJi5YSrQhsrKiTsYAEYNc+YEo2FstCwSf+SlrWowljT4oTjucGxCyI/
nMArZ3nnn4tVt3QcrE5d23j+9HiO69bBYVkTTPUlSnyBHRpviCl0wF3PQloe
fJLUYZry/xy+yJCRs5d411poIeJFpy26VP24VFV9yAboIPt4ztxoouF/zHr6
O0dFT3Z8co7RvjXX6T2rmTwqo9z0QVVFAMZSPzvAHauJTOPuLM399YHXYgcy
4CSVU6mDOP1Ep1/FNj7OKd/ycYi23XoLuwFxrnRAaX43tQRJ/Moe/yW6oa+N
f3aOjIr1oFsORBLtws8ccQPmxck9W0i/J2EJX+nJ1X7E/qLdwgHJqPy8wXUE
2836ID3l8RyAN9h/dYlnM3YGVXBzn6APzEE1J9d23yJXF9n6pttszDuuI2I+
DJ1+U2R5O/gbnvV0Um4EJnp5n5BcDGjSD/GsUtEtV/O+1PvclhU49Ih0DRB8
A7pZFwgwi7K/ZPfdFlysDtm6CHf84En2J9CMm8IDCB4HU8431VC/uKflmvd8
9ChRCnZT8EdR2QkPjZBVOVxFbxM0vjtGAVr+YYFroDsg23/dL1tAu00PTKfI
kaTKGzidbglEczs+N8GhRxw4BKWWPK+o1R6U5a3T3JdB8FZeO58B1B5/qWN6
Z5VjHPEYkZ3B68qXz2dFG1pTEMgsjq/chjF0W89rX74vWmpdILnYTwJo5Pgr
4HO3OGECgbxtXFjsxqy6fTreS6rjWUnU3Qsx9EMOw8VhwSzV6Hr557XnDiVs
VjqN1TNu5h10bG0iiHf2H4mauSnkRQ4LoqC3det+ToozTNjLdK5cjMHK/VKk
gWFzRj6i5AxKZeSLuOLoRVLIXP4SSCYH6d2ZNKqix6LCMbPz87AK6KXNYOJh
SVXwn/1wW0I5zaVPWoFkK5O4/8rqMN9t3Ykns4RvFFE02gl643N0ni/4k0VE
LYp+G7jT6phhvPpOw2yJLKlH9Wf6h484Zf+/aOfVFMsqSeunKMyZvdJ2jVtK
mcdyupZ92Fz+AokoSOy+CDe51srauUKQL7JtIm+Oc/Ty7JPmSLob6XVeugqq
UUOXviRsYF4ktMY3XcI9r64oiBYFuABMq64XfjVmSzvvGRb6BVA+Gp+0EJXV
ghF6ucq4wVYkTGotFygNBt3gmbLXHMEv9IBlnWoPwcwnvTyKcRsS9cA/DvGW
w7HPn2bbttG1rqOde0YNE8/ud4O0zR12Au6CFF195NLZ3/MGp7Oq9CBWmN1D
KkUBSzYYMbH4Stix8sHKXC5y2uIIDT4qxqabtt5MbmxGyidFdmqIZ96BCFWc
N6jM/AOtTMmkOT/H+pgMNVSDqdnzYLs0cdq5lcfmLeAQDR57bqTe7VMzkCf3
v/TpJAws0qqbt9+bXWxy984fpZvpy+72Adfmf02+eYbU347akb7vrzhZ0EeB
7lMmxdGdqq4tNqtrolViMqfsYQD9en4TeTWfEC7Unz3wBDaCDgYMkCm3nXL/
kc1VeJOueLe5+RRlnbBDtf3jcMjs2Ww4SRQ5Uftq7mTcofl9qaLN0+tVHpPr
FHmzlX6T4E9J/j0Vgl42vbtEH+zRvKRW2lDzYjb5jVKw3z00OAraSjy38Gcp
tQfsrmaY8cj8gF7p6Lq3P16JC309rJ7TrhjTr8X89JGe05deDSfFyPVSk9EW
zp/cGs+P3/pCNNhPxmxsKym6w95rLongf54T3UVRvxBKx0SCo6OlvMi2Ktb4
6B9rizFyKAaghX362/eaf4PVGLQgfQ4pthfnVSyPHlJLxxMFGAsD0RqktOeY
/+uEuC4pakLwIpTH988yDDwm2CCSBgFJGrrTJ82g851hU0hnLLypRlX85YxD
SvKSVIc8CFEGKEb2IfhtCTwMSsEllHApiMPvJKQUGnE48XSXKKbgB0HbZ/iN
imzOOZQYZRtbJ9nizPzHaXEEAM4BiNPEd7y7OM7XKqJr/JtFcBNE7xKuRMRJ
4QrSJcSW+4oIQ/1JjJyIJ7ny0/Y2FAxIU0sofKy8Ez4lgtVrcHpYH1xomF6C
5H6w/KUlrg6V+md2VnjEmAbJ9DFytaMBnQovYas0u8Rlw4Hcqfgr42/V3OOg
wO9hOkTxFqZldrYS7hFDk0nZoPZZdZGGfqOw5mo94+abHlMKMzUTloUcyROW
FOr5wBn8P0J/nzxOl5UOq9X5P+dTl+bk7aTfkWW4/FcVHPfUaB+itPUgw/mz
BXKeTv+uqXY4NIfaesfa1pJRZDoHP+TDhw9zZfp3DoFrssCTdcdUNKN+m3ML
XOUbg1E0ZQHhit5ca61PGX5ooHanXYMSbr+rOUoosg/VgKvtVaXtT1n0ODSy
ImhBARYvAjlCQUfYm+YyPt+vv3/8TrLCHYE+Jh4zEG8vPDIeyyMUl0QfafgO
bQPqFgHb5Cb7IH3+32qwgYVf/aFvIxwJZFu3O1yAE/PQnquFV+VpCRQENq5w
1bBOglufyER+OWNLVFW//tkXB8XfZ3N+uhty5aknIr14HJv9ihkiuWDEruDS
wWhW4PzHKY8tOK7nfjqV+ckWJnKQ7r2q7P87wQgHbkvn4RIqEzPpOJrrybK/
gs7cfPAyIPOnQxRK0hh9C2ACjxe4ENFOR+RvkT1zzmZhBgvNYF/dgUPHDYSJ
mMUU1DpW3OXWdPKJ9BpsoNp6fxXGzuKPMgHUmtXdCrl/Z2agN9EdpQ49nAHq
hSVH1rC/iVgFgv3x6/oDeVPJh9eiDY0SQ048mjd8Gad7BtIAy+wXbSR951jL
Ps8dIy/ZNmMTxsNTdNQWb+RDoOd284lDS026+H59hnEdC+FNTwhsp/Vf+OG3
CWYj8Nc+00EwEEmydzA8Cc6IjXVJDgJZoYysa0A3H7dh5b5f1XmYAPwucp1c
bJWlUL+G/tLarUOV8jUrN3NCrI9H/V4TcPiE9AnhJ3RGYjiuzUWi3VluNrBn
GMmF+v3rbAnllJc36aIUIjbXFXtMLY095QCQt8wKHNvISPDpZI/0Me6Dq3Um
fDLiasP6TQ3rS7R20mmM3XXrGpLuLd0fpEqhObU0aRCd08dVyUX0vxNoihMA
fxDKYC4Prb/WoOeIssyYZNrwXhcgPmyxmqMIgI54ScQdoXq4VnYIpOMkzLVT
KYNFOLjsnILtFD4W8OAvEuS3D8HGbpSgPOfhijw/u/hqZETc9lb+SgsHWBel
6qWx4NCkBX9ljECsn4LWJInwPVA7GPV5n/5fC4v0j0O2+gOUn4nvyY1BoLFx
dExb64S4JxdxRnGd61Ds7U/4jBwbVvBY5FOSsz7kTXi45EhjgS6oIE77Dvfa
xELMMg9ZQi/CcjjiP12/1C0k3tRrQP+2RUFGwTxzjI3F/jiXLEmgh/iTbBSA
pBVCpnHY6T+Une9T4g1Eq/j+KWTRfk0MePtcZsc0+suOuGoHLZ4+YK2NmPN3
TUUfPpryQWP4p32o1TOFqho0AprqFfqq8zI89J5RXhxcHCpV4LxDcYV+cQYm
HYUa5x3qFm4i1ajc7o1osY4TRIq/WUOjQXoLtgr4L7cYPlylgwYVf+9l5yx9
xpdkIs0xmIWX0HzAbI5Z2UV9ItNaPuAtyTn5FyZkYcZ2xDj9NZn6GPo3PRZz
SrBP2OSVX6Ieor6L+GojaaHCPttjzWiq4pAvURMkADfIPQ+2qG3SEoxM+9/g
nXeTxc1iU+19gVYwbBMO+0VKHEjtAkgHZNZ+wkYEhb06E2AeyGqff0eiVcH8
Fx0paWd/9QbWiKH2NruvaIzgLFKHYxEaEsXyCFK3hmEn78Aky2ILxLRQuEXt
pps7wxTYh5bQTYpLKNf1y7TvUDWtjxHyg44OJ4/+t6/k6NT1sCiVlsxY6pB5
L71T8xgH9JrXcnGmzaRwDwsf+Bv3/M9vMx3COdVwyx3CGyTqtlBvnWYbFf55
HSCCm7+Via6pCVNMOFyYVK4b6OPrh2wVJRhqbfCkQBHZ6AQiJBuF7mgim1U4
PA2AFPlnUvk1nD+XfbtFviEZz0vmqY7u8EQaiGdI+655Q4pPLKrb1ne8HQfZ
hNX1Qety4ARrqOfnDGKx5nSHnYD6VuBwfxW/nBA/07Ujxkbjb5WX1przRJd9
sO2AFOcXdjEXS+qf7/C+4A/M+yEE5LWiaFYTMjenuk47qUaFIFpFcrrSP4b1
NSnXX8485G8lywU7WeTqLtUf+4V/+5cXvb0KdfTmUK6umu8gVGvjyV2OzHCR
FMKdxNSQmUCfEsFvF7WvhhgieFoHGsZk9383yuyKXYwgRudtAiDr8oD/xsun
aKUpNpGlb49O/aURAJopIbw9Nm6BrAH3MlZ/ChHyp7Nm44/t+454ZSKnDDL3
oQDoHBuDcblQypsqtBr3YOgKT2y9DzgvEmYb+uTYIeVguo83BTOUM4MF3S3N
z0TAfEWO3+VNwhuyVBcxv+gg3nOFdWRXicE8E7Akek+NWdIuMa5/B7Wd1QG1
BFfuY0Ior+LLvhYoKCfYDjGL6VSSe/t+ZDsEG6HkLHKYozsqFwqyFeQuDo9z
nF2kJHAbhKO7Lw6Uvmlc/Q/l9RZwm6yG0zzlsjAAVOwLws6La+SSX2owdLcr
2xzqSaD45EVvRr7+EuEhYHL0+9i1sLDbOEIf3ZM90HN3JUu+dHDhGZDzL20G
SnxzpEh366oeCNSluMv78dv4WM+ABQU8yz/nEET5a89Xpf4YRbAQD3sR/a7V
bP8Ks4xXWQDIb8QmeJqwWOexUFZZ2ZvWPD3/eCRN9C31eQkHw5D6tcZrizWH
8qJ+dKDKjwi6tCkp29vxfqlyVfx0+YBAHGoWBhTG0HOjWiKA2yfLwnIr1J12
gfrbYaQKpSSR9UZNxJyHtwR/lC+3hIcDRJpQg8yNyM8ozA2mJzjE08P/tVez
BECc1RKz0Yd23icpvnxoNzkT/gNEFTiP22QNdpXX+nCRvS3xc+V/Bhz2lFcF
T5Ms1UXQahRn0RAbREHsB5T5uCYy1Stwg6ikE7CJx5ZsiWOA5rj3WxjanqZl
i2kXXrPFWTvfEtrmi5IM0SXIEc3PFq2uJJCiliuVBxRgSXu/OzsC+h14Cbbd
ScX/L+m/HeeVPgW0+NBH1jVF7iu+kCoVzf4ySXjMgvn55GEnP3d2KV+OEp13
C8KPV8Zm/s3PYsrir56VCSxihy2COORdPH6/Mf+NOt6r2DPzseulk4BVtqYe
FFTuVAi/TqfDivhAEh7JcEidgDNKzlAsoI1o/QASvOyCvC04EFIMKdLaYBQu
YLAtW3osk4aShKrtx6ExfihauHc/0f/QMA7MkFJ2jCfSjqbXwj7SntNEcZom
hiuXrxdXOTErfHJPSpXq7lKYw6zifGCJe0dGsqHGxhDxcyKQgeTVZjxPtjAv
pVkGnhsmXb4xYBXyFO0AB53iaTqmPv0vRBujTEB2LOzKKxmYy5FBBT3J2v9d
nCogQEwa3Z+kPGDHlCcHAZP/Km+48hlZbTcKhe9FTNyEz+90sOOLPfqNUB3f
bLeyGWFRik5PY3BI9LkR4cf1yOl2nYFF7j4k9UfoGxJkrkqy/HOfTboO8Hip
rkRLCc0OFPfQRAamN49ScqteknxUV1kIt46IUJjg2vcoMYoHOVr9E8RzsNwQ
a8tPaPbmGbaQPS1Peg/ormFZki/Y2ZsTn8GGfVQYz+sN5ZnoaR9vtTbOYxNT
BpMyThaZqy0njK3dCGNPBR3JoGAh6POX4BDYhLsYADCPc3+HwdIK/u6TouLR
dLGtuktbZrUr5udEl01uMB7ViaT8ktHV4DawIGKudQJ4NkH0dW8GbmOQzZLn
iKXEswcZx8BD2ChtGGkspTzJKlFYxffUUaXnXkkJPfvyhKu//vggYtgt6x3f
RaltjbSMiQRsNjh+Iq4aoev7rq7CjL3VTHM6mWeIq66nqFH4BumSuYdlywSE
7WpoO9z2sEO+BJggxJcj+Dx0FUymu1TmBaA/8YK+ZVN7Hu/MkC2DSrjawO5O
aJFl2BtRwJDXZZG5eAsUcooU6y/Q/QGBniIJISXvCG+Lg+nqmjB0Ys463vb1
k6N/wNjMOmHBs85JtWOS8JOWWe8We1X2hj6Uld6T9zKd9clIoQikFlWoSL1v
eAeQGiyp/vrOJ11D+9Z09aK16Iz2azMUy67DwL3AVgdyZlr3nSRItjNtl+HS
R72Emlf8EztDGqUQY6ysiOB/pqXLiGs8x3VkKh2dImobcPkqjF1AU0dzstKM
KEXFWMHgR9TDxobfSYRNjXgZKaws3c61IqBzOh9ytJXlOxAD8H1u1EHUe6td
NiiOkNMFpuZ/NSSUkackW7BqWZoZl2MWUqSH37LrUVgPdSQpbE2X5MNTy3NK
vsCMQepe25Jw50yIcbdTwbk2F4lVL+tuEZ5I3X5qi0ivH0MUqjRpIR0cvwsc
TWJLsv3KrJFmKkqZZPsBGzyyGabhTMz3Y2HnB2Kw4zspbyaLpun3ixJWijcv
mmSfeopf9UvLDeQIcImVdFFQUaWX/RpYa4LOOOKy0LWpbjo3sdIdbPnUdm7X
ZAZ4z4K/0IUdvJislCuR+X6GzZK++3LduHhMuzZGmf0or3RzWD3VVz+fASQW
XxXLXkf3VtKy8Sn5aF1jUCImowOfnUDvDyK4nqauguups0n7jhzPdgQzr5DC
fm422DBmNtquVybaI9fJBn/oVtDPvRvf3g9AFAPhBtDxETgNseD6FEtiEKoO
hbvKrojQ6c/3ejBiZQl/XXDWQdsDvQdb99vLpRqqmZ/FaNMcxExUO1hScCyq
O/ijKo2AeVOdiUpHJTm0slUfHNMN+hHo/QcWULAqZAZ+zdnZpBnCdMJgAbqk
BTsgP6yeiI/GzcpeT3bOqcTsoziQjMj3+Dv7bbUCd1MmoJwFfunSDxYFxosB
4FIxDCZwRNcmAMZTtA7/cakGqg/kOnrD2Kjfns56BqwW2pKvLuv7amRdjEja
ALPkxGQ+25p4F+hEcVTJ/jZrZ9LWpOyooLpnUVvVa1oWr0yuAVWGn8WfYRhW
o799D5cWMCWHIIF+B/MWwRP8NfKNiUQ6vhbvTO/XCYIe2P94+JqWL3vLB6gQ
v1+GDTJLwRznUHni+nA0VE1eMxEGJCMeO++myf8Key20+WyZzfwzn22pAQYF
zs8tP1iiunXXXBmj7ruLM4EbYTFB489DOjM0Os17PpQ+M1n3TjigiHVWBl9k
H+OpFS87roERWlaLMLWZTYCVC74SZkWHSVfLT6l6UAw4fiOAWzNWVcWfS3xw
tE8f9Kusf5IA3J88YyVjLJ2NEPmwP0y11HvyitGURuCBj0EsbSjUA4weT1mx
ENG6NmlX2PBT7QnpRwwHeO2LdkGC67LRdpeyQsRshWtWS89n+qp8W18wO12p
sP69i0je3ndU5r/1o20zNOU+soJurfcaYtVo3ciRCf8N/4arfGBFSyrMmqN3
n8Q8jfecZK6usWOAchpf8WiPSMOBzJszQlXzLUwa0AtVkxrv1U9g9sxGt99N
6jQkYxUUdpm/y4nBb/DLMs17FZTLQXm8j+NRcrZuSE5C35IRIrY4XVoj8kJy
lWLPmwB89n8rpxXXAAKvWjlgSjPpyXcYJ1IeOulul2ZNjMXZa4FU+C17hVKo
/YjjKun80AM69UYZppOKlqMFp1kRWSEa3YPgCe8MlchPPQc/aMunbunuCpWR
QOOZzvVzbX7JtcFcZv6ipEDxErJXdrvT4mef9n7kq5T3ZXYn3CksMz4ydU+9
+H2DjK/yOlbWlJO1uHCPtY+p8PteqqtAtLlRTFOX7EKuzo35NLey/lqFVdDi
QEtFdrt0EAi81ZHUaqush/12bKqo2MHWcxN+Aj9Dy1BR0/H9xfCHx6IlzeMN
ROyQwf6dSIhiYjTUYqOqVOPjv88khvfBWIGPkPzRDn32TqjZT2DZGq+CVFjZ
/cgKYWm/TFU7cZCzQN5DLqszWrqXbVCMXy6F6BLoiPM2/SBRSgLSbspyl62j
30GKq+oCYDKCAUePaGqqzeOjC4PwfJUL5nl1urztGX55OF+dScG7s2tQQ2mP
fTAE+SCeEBfeC7frw/5yYmnjap9qArtZO4K8C0QkJN1xloCjvr2n59AggELM
uDwCon602RDftLPYTtjiLdeQ1kEYC2S0bPQyQttftKvtmn2mwH0ZHhFwW3Ko
HwveGOKUsvfrWmP9Py8fpooT3R/b/SflX9Xe1E8gbxfheSQ3tVuZ6M+ryE32
hBkRRci05UgNCXDq/GtbBvzuAo65TQRR/K+fjSktsWqaNPA/i08tZbm1cC+k
4zXTc0W92Fch1cezfd8KGyNRGsWTXuECpRhVUfcFfW7Bs6MjvttUkNxjiv2v
wNVAyCs+GDZhfx84UjMTb2GWcDcwCBqmyXXKqB+DZjg8Yt434nRHWXZsKN/+
zILCd7vYbwG8CD4n7L0l4R2GvMWbvZIrxLJlTAQJ13lFyltdwuNf0uCq2Uix
is5i8iFDW12QEZ/2OYMAl19aMpO8izzRuikwdNkgk/dfIHTIPRp2GcU/egb5
zm+Iz81O6zRRmpggdoKrERJVyz/tQelFdjkof2nNDhq5dc48cQvKfb50Q2eJ
22qxX+vyQ9MuEoebPB7KmfA1DIiDKuni2768VswcWOxEQA1ECC2dKlwXW+1y
lc26ixn+KSo2p6xgru+SZdbolS5P75aGmAmgoJqyOH/vyuJB5hU+1vREUvDM
hYXmEkT8KeHOJQFonjt2mMWvyniLm3QUy6OqZHriyDx2C6CXS3VkQa+an78B
3W6cb+yKxZyrcZLJvE6M5A+emWhKhozeF9+pJW33eNGnw3sQD1una3z43S5j
jEshcSHMIKaBlQmORWwNrP7JwqpPXiqhVooiHkOn5o5GkI0jCKYPH8K3eCSx
iZfo6u1YX9gD/ARdF+PwqQExaxyzw8kOGp6xo7KJdB2d2nsg0fr4J1nIEdPt
ZoajgfyhI/9RJ5xh2WTxOmox3Qkz24oczMoaLtf6lqFkKOf2aUWG8bHENUrc
ivLE5IT9x5fFF3+JtxCucZ+9bhQj8uyN0UmyepvRH/LJZ2TWid84NBiqdkIp
z8wRkjKhzq+kIf+neEaymH0Uy4PbZEadepP4R8XYJcSC1UM76Cmu3tBwJgHR
ldzIxLF+8fApthZN/wrPgca8Hr02YFKI30zzGx91QtO+5fUWN4wKjmfHzjTg
kxpHkL9vQSwrduqmOSHDnRhphv3hNi7AFiIBCxmadv1fnbYG4n/jAJuHTBeW
ywfERW1+J5isqYFa6Nk2jKvQy0tfa3KdjLApahlNyJK/WEMwCx1lyw07d4Tl
eYtQXTtQq3pyLlpr27ntimShg/qSRPTxfI9owlJUFB2Tu3U/wdNwjB39C9CX
eVXa1qK/gYAI6cr5WgJ5WKLqhQU0Q2zHrJeve3Wlq++J1MetpMNt8EWRgXKC
mzzDFtDOepaM4xFKtacfbkRopuSp7+kHA76vLMu8Z8LGFk0F48iy8dUoxNQC
el1RWFOSVmYG7Ep8LJAD8ZN5TVQFlwb3C2JEnT99GJHoGDrouhJTx8vOOqay
MwRW99EmzqVi/v6AjBYLKyA9x3zf+fZb33i50UHs9rGmXOlMhpBzDd6gstii
RfQ42gSylH2lQAub8lXQiH0kgAaYk76zsh3cx7OkSI4evGy3NRdTl4xNpAil
gTjbRUjdOWu04/vTRgVq09Kmzt9dOeF6AE1UJjqOfDZSgLyvKBunBC7q5Xir
mi+OC3qJU66XTJUEAKNidRxTAWBPULCbC1fDSBXj6DB4bwK7jt1972NyRw63
umA4/YYjTJPeEJthfJYVNcR04NPjnLMMTAn9IqaeFYfQVZWiL33ikjnDoEeV
pgOaxpCY5QYVq7hEx8CBR/hItNs5TPuOoKEMVcBti8Al6x3UUelK8Dt0oPxj
8uXtljsyCqR7KogZQK68u02I/+y5Zq2Cj+ETntJGJuFBW+yIpTSOhlnHARaY
Vs59j/7e0YkONe4Lbk7E9ymX4a3eDm+aD3pWOTwXIkKAa7JVXzvc3a0iqPSN
1vnwgZwCyu6PUQwzTF0QwkuEfF/L9xK7Tns1jwdzLePvMnKgiWVxAPOXiMqe
jSN3ftD81GhKZiE5nY4Rdz2+K1hC+4JKevk910mcgVONOGPZl5MCdGBPg8m1
xqdO5LcxNZPPaVDJNbzB4iahPpeCR/MV/c3Rhvc3TXFPpfY3iqVTWAhefv+c
gpgPPiys3PQ9Uc2o6JFOZzDGk0U7nwAY/YQCal+z/XuG7DWtSb4dvKJJ9x1Q
EwCPCJOGaGWVnraTiiwd1jPXgcPuClFrCjaV/WQ8CK/0hIOyBreANPw9Q9Bg
YoY3HDXzPrX/85renIGpS78sYSH1hvFO6OQuFYgjrJYoBb3nP/y9wB5ZUszd
JcNPtXgKGEIRiXSaf25Q/B2nOAxsg8EgwRZ7YJWqBCMZnAMB3Cvgv+ySiKdw
FapjQH+MiQOOjvMhjJ95dQ6R5MTXtzB2yt54sUanBoP2iD4uCEe6bEmpz8mi
JM6l8AD0bD1jjX+MLCQYsfAp/Yh+cMHrG0Wy+YvP3D4o7XC/TdJpnwofNGT0
pYEezpuf83/4kqlAYfvvYTOk3ec4fVxvJQ8dmeyWaI6HULDuxgkFc6+BIW87
SVZRF3RMvCQBS+0ypES72zaLeqFvvE+LN5+zTuJ4Efq1bkAkDyWK28zT1v5N
HqR3vBB+qXl7SN/UDIjwqzQOewxQowwvXIcuoAzcc0P7SrDp+XouI0tfEPsU
mg0iRRXmrNmYSFSfum75WPi2FQZWVc1RoLOejWcJKTySJEZWrDL7S2O/qr2I
z9RVmQ4LUG0HWtPzI6tmodDd39JI1pthOXEfv+dATxbq2MpHLZum1Mx1mx+N
fdTSsokG5fGPj86x2MC4TWu/9+S+xT2fn8Z+J76phrVh8dXpMekbtstSblf4
1yfNr9l2GI+2E8Q3Ia89AMRg+zo/zwyDhIR+I1NdwbAN7b0mQWMRbCWal8fJ
D5SJHK1vEp0w/MG5nSsBSNyCvsm2PjSAHUlsFyT8Ksun4b98BfaMpz3u4WzE
0rQK3CnbddjakRZ6SlBLlv9vkuLMTnAobSbP6k8yObhgRkBkRZRnoSp9UXx4
Kd7ZZHRhDIZxjabjLGhZ1GMsOMWVubczLPprbzuoCoawPBdMSqQ6WsnUZJwF
rGaR8MwjvpZf523HoIc7cwq3iQPMB0jteCaHdYyBZkhIdJ9wlmF/GlFPd7ko
fSs5qSp+bWlbTR3RHolE/AW0ZRI4HRPn4Rw4sh3aStxJXoNGwerK2Qe3S0bl
l02QyXgw/5Q55MWy/BErvxUgtOtvhRhTh0xLvNVkoADumJ3aGrohHn1WAp+W
dQefc6zn8GkDaSHMdFWOju7Evvctv2ndy69gmQam4f3xjGjvgZAqWwTWYxl1
Z4hLLSPeHsK3r9HDtHUb873VcrVwLnxml7XOvlb150A5Ev75060f+19Q/i/l
+eTL3FcsWRYs38TVxGW6oi4EQt9z5mi6aD1W9lHw5LUJze+ubrN8qLURSskM
ahuzV7o/dAbdt6kPFcc+rRgiezAhZnkNBiFB8R5Cvsfkn3Gb5Jejg9LsL1Zt
A6aTToxbMYb4njgZ6GSHTKT9xCoqCbQlky9svDxepGNnx+12FJC8ZXzDreZc
FM0jXl5w89LmO7fiEm7YQjfW2sdE+ZRgX3Sc8HqCEoOPI4BgLD7LDVYTc8v/
jYUtwme5iHva2ekFR10RwbtYQW476J4C3qgM+w0W84j+r+uKPHCil0PbHzXN
4ZWHVRlHHlrSX/0kMwnsimA1Yjk8O0+9n9r38XIWKuckp3sxUKAAJ9iRtjjg
FtujLgN18FsLaGWaNhYIBFWgIdYgXqL+9fHBKTt7TqCyjhsVUad2ZnQcWn8D
504OPgT+wrvPFjTmZ3elc93V9OLXvqOzZMwCb7v2s41i/PHQEtmJWeCp5Xm+
7M8bv6eHyhbN6ejZygY36E2RL1tXvGOMAZhSrqb1FqEwyJdGpqhnw3Vb3K54
0CY7LY23boym9DEiUUbYU7mQfcEHXLiNbAr4SljKnDkdh7pGkLDCiA1tlGuI
zySbZHCUyJgwyNCPn524cyI2pzYEAnj7C73CbSiK8IJCc8+ocfxhBjbJdJpu
YdHb6ZUDPbM79+Xzuxtf/EMJBR0t5bDCSdpCN25NmM25Mr6MYO5hxZOEVpAo
RKjIIe8NxigxhMNc+ph5BZGQYffhmzL1JqFSqtwCujZw1ZbgW4Wr0lOUJSg/
nXRlsHlQbAfBWEqoUfRXeaC5BXuWm1mzYvHBh+XEeNCdhxVr76ejWXFcqKcF
DZ18ymiFpAUcrH1vZFKAZDIzQvtLoB/TI93RUEgobzOW/yhQSBHIEn5OOT3C
iScpaJj7zowZwt+JXyv3m00QbEtOYlstXqqc5wNr6g4pGtO+OlsYxbrcMGSq
i2HJJahqaRoAGvDPkCCne4Ep3nn5ERqPCoUkRweNhWzlUj+q/VwG2z3Y5LNP
+L4AogcA70Ag4+Di5eWviaac/vfGyNpvo9WsPg5vzd9/PlUvuEQ7VZdRmD+n
FaIyNCJGjOLiXiOjjFv3uGlDhumK+J/kFKEB8hVmcfz/LTztyU4JvhuLh+XV
PQ+dgCYtLeRzp4vOyG+UfRxw32qhrFTGF9v9vbVmmp5ZQhnPY1MLwfZbXcI9
imykIMyz5dhhU5NratxmJ7gkzLiZHF5hQfKinctkAhEC7w9DGnsatsd+J0SM
siHuU/lRZ1S6bfU0YrEtAwrMmAYeFrKeXlUV5NpTb7J4taD7+kOtNisNGqi2
XiOOnuLrAvXOKApCS1uyO6J3j1rq0Fopqu8+wuiRlr3qMCzQOId7h8ZPoXqE
D7cuDnIF4d49PY7aptcSHExxOnrHauTEDljspwS+HO40pdh9B0CxfrTy2iL9
bja0CsxsWsEZYP4g2ykk9iZeUVg4cwPfGqsMw8RU+R7fGlXF+0xtMIIT7T9O
lxM02JqzHFCHsfIhqVY0tj1WcCSdO+q+lvQy4t/VjSPDk5PwLjKtO4R82KeW
INBQw3ows+etf8JT7CEC3l1kWQtAA3qB1vaeirVckiHflnlfiAqbsZQIFiZ2
+AMXuobDJFV+jnlZb9i6C1EtbUQfiCV7rGpOzo8QjQPCFljx3CF/R3OY8j6T
7kT71KHf5Nb8prTyYLNJtMrkqexlyD+MAUpA60dki/J0RVHOe+CqYLgqYksz
59mESTtREYsrfrZMafLDIXkqQijDAkjEAaUUYsNdMeZRTWqoo6GLrmoHPSb8
86U5jgmKHhmVQphCMV1E3AwdRkrkrpvLRzl7UGsKjKGC1Xt/TJtxU//dch85
L/YWckofLvJfY5WVkdkixWOa0Lx4mersDqCSTiwrUsueykEy+qZYcs9GEFuA
3dx16glO5qnoadEFX9RtEjzGtNO9VqGZZtT5kBwU5XwfG9/7PMiin9HBKBi9
FYNX6Wp8hB8Dv8r9BIQHOT51aAWKsR5kkmmVwCnvNCadwrYIBIVreYpEOBld
eezFUqfo66fhrMf6leITuzYPpRD2Q4QzNttxakZy8X+raMnIRvIAREZ7tUHk
IhnV56mFwXX0/XVTmrtX8nj24EPyEnBnuwaSMlgPEH/aEP8NlNt81uTQgm6w
v4ShF2k/QcMP8h8j0YCdpf6sXG+YioaG1UfzIaY81zOZQhSOYSfnH8SNhtOX
IifFr1jWiypxrGNDgCxiVpeLPV9i2H007SHUk3VzPcQwEX1Uxi1OTnMf63kx
2JJNMLiI3GT9zpwgvTDw9eSqUIN8MteIdvhZeO44uwe3DOjSdC06PI9zBNSW
mGpMXJUvA66HD5Pa/vnOxFZQY1AE/JQ9I+8/XPL+AqQRrBHB80sFFps1AQZM
0mq2pXOxhGNoo/5YHY+BN4WvLEbGbIKN7zojlzNv5dT2hoh3CzziA/rcH26x
22nDLh+SNnpurwzvCfWJLyN1Xs1TBx70ZrmWAYApfIBWe8id/a9OBLMLV1Js
A8bRA0HxfxF+9MBWA3QrWytfNO/axg4PnhUSOtmXdVVyTsyGbJPIls5lLuGb
FpOTut6SHmduD4VX2qHp/rQz45HRRcb8bwZ0/UFy188Na2HXtheO6Qt2db/c
B+aGpGREKspH8DhSVHjQS7E4kTHp2mXilIsqrpgbAVn7resBzz6HwUkxsy+f
oOb9vGtP9MhowASSP0eE+koFmt+EfecjzuknI3b704zaybs6OUVIJ22JddoQ
EEbYIEBX61vLLNJHQLHeWaDxPVxKCuM2zzxrzlrv1J/wukSiYzLsVZaq00/w
P6hSlOJVl1oq0o1IonL9fZYip4C4JuvWPDvAS5RQL0QKzkS/fWzUPzdBqYYk
rdBLXj9xsYZRq3/nzPbPJFHIBKLG8BGBQOYop4bchWAQdVRr5adAVwwhwMuc
6jnbNs79yCincSHvtAQVMA3tbE2UYklHwqJ/J814BOoZOi+Jn6gOwuvQdb1p
VxsO4lIsburuS4ActJJt0oYq7G9Ce2DcnqqBry+kOtTRXbvj0ZU1JEhumQcU
fCsVmksss5qwTx3sgEZ/Y71pmmQfIduRMZnhzYp8CKFudrcgEZsp24T5LO9b
nHVFwAAmNl/O+T3TqkjXVPRja0NJ09730pAtUPNXiJTVdFhVyC1s+i9ZSy4H
qJsdXEIt8zU12sHGPlJhLexz+UAhMwGXjK2RKjJjeSGlr0Uu0sY6u6WRzmap
xPU4+kEMLXp5VS24vYVSbX1LTYBlGqu4wbFZgUzC6KLF7RRxvE6CDYDFIUpa
ZHIZ7RETCAt63HgzxHxP/gfstsN3ZsJ0E8TRSgNgWIqxCuyudBmpLdbvY8L9
sKh9vtKuD2D16pOpXRxiPaaQfgL50CYkUPWROrXBTM9M58tq9czwXmKnGmGi
k3E9O8O5/B56eExL3qOZ6PLm3zjTjvBQKv+Ev7CFAnCrt+SSjykP6So13BeX
qJUikpyhM3Zi7rG5mOPwtBPGJV4qpmYwbsAPC5xuZrDTM+Ydg45Ox7av9W9U
8+7wKBkoOkV7yI1GWLs8lEQQ6mlqncZgSE2fhU1LByGuSYu/5kiC7mAkgfnx
73VbSHcdY6Nw2ipPp6DB3A1ocit26/HNB1/oDQp5P6h1YOJYqRy2lYZS9MSd
h1cDvrZHjuX/ZYr5hQOZVidiL0fUCs75qw3WS4M9UrkI+IAU3nWiw0SHg6oa
OOfb5R+4kEvn0Ef6AxjLrzw99qHYnKSNJTk1hNtgo+MFN008Tw+hUVgGm2Mo
gWLg89vS+2x31RuKMAXVQUsa9Q2a2VNZNwgJvFRaUPZgj6lV08HEpJ3Q/Y6W
vmsCC5mm9RJcdBkZYdJ6GWPMEwg5whQJKQ7nNYmZqUKfk8Ie3Mow4RPre4RN
ClSnq4ik6c59MOrv+NFCXrykDe2opVyOI+FfmO8vpHVd95vNgZguBL4/lt/a
3od//6XhFCKEDDtWXTxiftZpmyGZYqgu469pydq2wLb40+3hbtk0W3gLnU+q
pn8Ge1Wo9RBLHjEd+vQipzf4s2R+shulVI/JTfGWyAlfqABL6/0yUjP2OZ0l
/JsudhXRTCl28+uqhtboeNRT5wwuVG1NvSy5JLvu3EEz04QKIT0vDUSsYS2H
vUW+yug+Ykcte8kEyWAtKrNGojDnhIMXbbX9ovcT0WJDbxk7fzS2fYEl7XL9
7q0QDWPjvCIpJo1B/DlI5MjRRb5jX6FZqiH4Br4usLS9DeD2gnN0e/5y3bJD
sVsWMjCHenMGeAovrbDDuJycBUu74xoA0bdbvziYaE9gFnG8VI2v+ICzi1cA
oEwZZnPgQx/GAO7EJjFs/VBgU6mwdEMtbVP9B9xiAzzNYBNQh3r6OUnCDcaX
/pxYsDsZehaEJnsOqqvnlCTGckrhyGpwJ+Hs8t2IJ6KBNCQFyCvBGuHVha4t
SFIKa4IMJ3vnX+e8BL+ZgQXsbSnLltihI0/sZ1Y3zxvKbCu5R0uLT8PNSbk8
biGhgVpBj32b1wiIgoc1gEQl6F4Ob+5wyAWL/7aeNEYWYk5ihkfTlMzYdQd/
jhLN6L1kELRkP3SzkFeSydHW8saJ1690uWX2o+/L65pbR0VGwqvZ7eD9UR2a
L82fbusH5RDvSgZ/56YGjhfJ6rQdO6RsHqcfeMNsDFoXpFdTtpW46m3SQ/kx
8xHz1jUYp9/ryIriX01s1XL26hZlu5i2goNOZCHz9ripztxuDLuytY4uAsAe
0jdVkcw0nAlcjHfGLk5pNwR/Om6vIGkaxPRJnQa7ZDlmxH2QieCQzkpdk7+u
kvU1ta/wtwHTBY1euzMU0go+9mszoJ/HpOFrsF3sbTD85Fje1MGpKkQvX7ed
tiJUiDm2NBuAwV6dDtqLwSzfGUKti6W4tVqgj+MNUswAAjSw6XCa284ZZDPg
FHd5WKu+75eKtX/KjT2j6iFM4Ig/F9oGRkkup20y/XbBWpyS8xerOaO8Aqyw
cN27UxOW2feOu1DYHBFxB623SH+Ha/jcr2gYzaJG4/s84VUbGkh2SlznO0SD
aURVpyybj+KKEjENo88LCcF++DcCVNMh9W1OKBdB4pTNZASReSH0kI3v16mi
QZFBWMKbWONSdy/tGOhXfqn1hLGuci65hZ+78X41U7eDnIqW68MzfO2luT8w
owIDWGIEzrXyhSu3RVz4721bYc29rFaGIBeA4n22eHYcUieWSAzusRvI70Fu
yLDP/7lsZJgdMx6Gn0e9JdAEtwyJZtc85vo6P3V8795WMt/fFlQAn987YfgJ
hZGFpN1Zn8xzfAEB4g32O5xchBfrXACGE4ZsO32wvD+arUesBnJCUfsLrQ1/
XetC3ayPBpx1/SvUzlB/v2oRr30DJMihpJW1TKpWWWOmJBZGt4oclMas/R7m
vRLXj4X6w6Xw9Ov/R5s3tlfb7LsFO7rTeaP74h8Ti7n4NDiYIfe6zv/3t+Qc
p93PhTgdF4NY1A0RZ6HJHDBoMARNuGZkSsOp3ZlLtHDVR6Kqk3lYpj4gp7MT
J6LyrWX4rhA1omoyco9M4nwnrzvlqbsE5zOJWXGIMxABv6Ef11W3XI+In+JB
Hxx6c18HgoiSMTLz7Db718SISe3CSqZlxB90Wc4Q5z1BTBgNXj8aVMErj4h1
JdMJJ9nLmL0uVduYEwqxI4Q97B/rEbvc5WNKzR4Lml60H+tvygIf7K6cuZjW
0/PIrthZYcxZk19P0n/NlM/HKb44Il+4PVq9xtr+pu27lzP7XESoTWN57Klo
EYy+YRBlBpLgQe27GEcAxMiVE4tEut8VDXn+N/tSjyc7wIgSrgIJjQTdi4F4
JgarSXYaosMxoVpYX0L1eNjTZrUz4kEfSiC34/mPd0O5genidK7aeBbtZ1F1
ny5lvDTis9Dh7zX0V2bpA8JpiOiVQWoJgBd9w7j6ZcQ+matETNWbwOpQlH3q
BHUEhAlaIEKdXNfGfcrd5mx9xMEjJw15eNuNBuaDJXuMzfkTINrqSYI+38WC
DfR3F2KafJYukn/np+BH+fco8TgGN7N4/ndKBXOJIHdf/hPMYaFE2whq9e1l
KuIeVDmgIMjg7p7H0TkRa6WPsHOnut7WNem9kzYWvaNn1NrJzaptsK1jothM
yWolUykXmNWU4+di05ObEO+jioUY5MWBMrdaTeyoVUMDza+jzZAb2BW4ZTtz
q4eDarCPcmt/uuEX2pJ4LkKVauHYzaNyUqPabim0FhL/bq9DczCKCojyDVg7
KYjt9fRO/BlZOQf1LHHI4L6kRBLr9ECV1uMOlfSNIj8T2NB6zLz67/+Rjv8u
IYVJ2vrsVYRU+jNv+tUINUGBOxhXBAoeXWPpgKfIEmpAlOeSOmnxPlPhSfb2
N/2Lhwteon4UVB06Zx6dccu2Y1+syUrsnoL7MQPOpLtGxCIz2bsLG5rkmB2u
6wMHk9VGeMetwM7KO0g6WnhzQnAX7wOT88nYVKiEo7olJu/JTI2OaxANQ5Xy
eOXks2PlZRiuHuZZX8VwwRuXW64uuGqOJ76m38DNVbKYRVhXFeyE2z2ePj1p
i0hE+eW273VXW1Ldpcy0Swa8WrvTNNRYf3OJ/rKCb7zdZaLUx686bQGolOFx
ZzI4MhSq7eIMkGcKA1zupjuaRhfsB0dg6Cf3GcTHlUOFctFZlMMUyq7i0L9B
JvUtN2u98Z3r7ww+xZG05Xg3lwHVqgRjaZZuHYV2WphXXWky7UX/UIsK226P
xG/Yllsq45mwmfX9YoPVbaH5+gSTU10Ou5U8WkmIqv6ozHCOw4XgUMnhq+fQ
2x7C2jqWX3CXhMWSKaVS2l9SUhxGB2m9E+Gk3l4KGU3evFtTTXharXgaVPxm
DA/UqsaK/iCzLtxp5GwLHCOFD6mPPVfOpoULCD+Z5ObIHz0pzSTWopq1mfmd
oqdXbBOWfABT2X4gft++ELHBMVyizxpKZMkolMaYNRIb0ahu8Cf1xDdvDJCo
de1SdYAvNnzhwb+r1cwXoV2sZH+26pnlyQsB9JwbndiicyXV8HjuH1Kef0ah
y+hMx9Vm2nPh9fqCd9jAnWLEFdW4UBFjH8okeHrJRHa0fjd7zrS2B91162Ff
7/BUmC17/HLxEWRF7VyaDzm4AtjL/UQRaxA5BvCrlccGac98Yo5yPEjoklC5
1io06EotA5HivI7QqPTcyl3fP+3xCWW/Xb4UF6DHJL+gc9v7208xFuSrQ36h
mNx3/7w4U+pI0OuprIk9CAWdkR+S6y0qDWIOPYhNQbFyt4tBd874/QV5YW+k
VOOZ1SYguFrrWAG5w0zd64bLdZp3QqzIMw6oE44MmM0pMr4uGN4lZ0z8NizQ
ekWMXhLA0Y+H0gQdR3zLt7KmXqu7GaQuoTXWK9A7B3psl6JNv8fE5dshGtYm
pfWk+VXlHRV9buKQfqlV4EbAyR3O60WN4rj8Y186fgPRpEH/Fp4fwBXpqQFc
qrPSMUD1suZwWW7iPM7XxnK7z08jpjiq4cpn1b7QZzy1g6Vqs94GKl+1LI1l
88iP7MZ6icH9RIM+4del/WrTpwu9UmF1wBILXVD+mK0/S4Lm6bl5Rwshcw8/
sVj2BB/pzOIxAuikBwNtuZkD2oahGPKyLeqqQuYxAVmdJolgbuXbLLzAMqgo
x1LLE76ZIBC5dYj53S0wcT76Q56OqZ2Kxk4yWjULyFa0gssj7kX3e6qBQDjH
IEcwdaAA9tas7Oc/tQ+oyQZMUAzjuxb/TRLeRK46mhkbhHH9krKeL2HO620a
JlKOXtlSgBzxWekpND/BVb01wFQWNF8RK2e2k9l5gHDMoABKtCwLWKKwB+dT
2/j5+TlXmxv5rshcarqrq44ycdkYc2w07z9LGOyA8eywDcQ4fZwOzuLD+WD+
n+NuRQaEs1SoYS5hNB5AaW4rfsvjzvTQ1ZWKapY1UW7BBw8G6ipg4fk64Zmi
fIpSD++vlu6EUWZ6MtBqysuzkpQA/PJCfNE8VXF9qFz8FeJW5Lu9vb3+/s/L
Yn0rHhBg816MX2Y7X0Vq6Yd/E5YCBy0ezAMcXhKNeqmEbcferc7voKwKkhv9
fDn2/KidAOhBZedqvIg4y8HD+vVijNdE8VKL6xLNdSyucWwNDuXUyV/5ixJZ
HkH8kqSIw+zpHhiAL2YIpfLZIokJgUO6xI1PqvUz60BBoj1IVHIMYCREDToH
ONYZDcS7/SiP6uur1FU2cE9VHwwkhOPFMFXaCmjY7uDHNOOZzT2PYVkkEIuK
WmXNxdNo1muyXsrWZOdOwPFDSp+tWK7dzXqloJxJTKEWrFDBuLMz6FQsvnBo
yzBHvJh3ub+ss+DAxr6unD4Yue5tRrTgm6vwlukID3hT3xE20+YVW4oNkcPz
PCVXuk8m7Wv0fFgdWe0DrP5zCq1ad4qw+nD2ONz9jW1UHBykCqZNMfHFjUbT
Ml1rvhKrlLnw+x6r90wHmssj8kaidxwocTlGFt1ZPlF4xACOqBHmoTkK9S6y
9OA7OR/yuFT5+f9Ra0SuTzDS6tCKM89jejKHI2vwrL65GsZBfrlcg3XWmjoH
cztng2hydns8JueBJT/IquUXO1nkNhmOF9MnQL/hq1Qc/j2HC/fD8AebEzIR
7WGfvo/ZdXrETvKeIpRnIGzzU7E+022M4xQngvzic+NNDKCksP3pkYvOg+bB
1VY2KVzqFol6AMpbH7vwe3ixHikFLvmv8wv6ffTiYT4NPC2OEd6J/Z6nfPGA
9mBdroMuWnW/gOb13x638NMrKOJrG91PG7yVFDfIvzFABybHDHUFvNHuereP
P8pToQj5+ttU6s8/bHPUQ70e25eXJLEbz3R5OjwsRs/hEPv0F4mc6qa7XNxJ
nunoA11JFVd5/dcJUvrdSnYEEEi+Vdpu9M5j+p8DMyR1F7FDDbXhkJXOQoOx
Ab7/nTj0RLLZm40x11RYQqL5DLSKY39kxw/TSPoc0NnDb+5ereO5KMpfjnsJ
h4nkxWOHAGa/8y6aeHMkW0H2sVeFOnoUO4p2db/Z7ZRYwgO5imdBY4sRyKjz
p/KVQfVFqCzpcIIVXdMc3z1pWwVgSYtdjYC+3vBYI5iHAHx0EiPfyd/82QWT
SMDNEU6BcpdTg6ULiSbQ93VaZy6waZNBOziOScO5WHyW/gF3xaPWcUCClRJ8
2yMwJHGp9zxaFxKIn68/bBEGeN/ZSsNZjMrMOxabBsZ1cc5QEs2AldZf5hOi
bI6d3d5VE/t1DFQ/fQeuhyguWJO1lxN0Oii+Kc4VQ7JmKHBONWTt0rruPr6F
hA1n6RSANCE/GRZtebfuI2Bvmi5AI0JOt2Dd5AFi84095DDeQA6/B3ZEvr6E
GCtfT+aPZ1EnKtcKo+N/8ZhveE2M8tgY92kbG2I5oIeoJHRLsqv7VVXvcCb/
BlIQfFWJ6GkWb+vx4Kvp8yG/Bkw0pyhv25IZrP8RyXdmtMmwCQLIeC3Ufpq5
OxO5t5g0K88OpT6DAjObGxuKu/A4LQRlj5i2Lw7kqVi3qPSqccXjueLksF1M
8rZQ3lg90Rs0WqzkIQgRBuRyBW4DpcHwfDyuEfab8y3JDV/1WKjykZciXKgk
Ct8xFWMTR1rypbLeHG5o1GOUxNy+JoIZjlu70ex/nrr6/tdtteqnwCM4O0wP
KOnJ7/4mw5lZBCMIgj/HSNQDsBwRBTXljqUWxsUWkm4/kvHF5K7y2svxaOx8
4IDvCjSveJrOfOToEIRzdEVbtuF6FJXTcauM8LVZ9KqzY5l+0SwOKOMpzlbS
oIDDY8VX/sza7pm4PkHgBXCj7gH/1Srr1EYjfeL8rNmKLfxRMqRRSC473Znl
cmWCA9QfNL1vQ3jPr+cM6WUMmHTwIiT2Sgnf5nqvtLgR5A70d0eA+7f3YbGg
FDe7WPGGoVnVAnB4FMZmEwYBJUcewDJX9EI/6Uejdkw2Tk5nF+7npfhwU5iQ
y+jxmk5eVLaVK43CnHti7cJLJ2fOUnkymggwIN5hxO9X00HOChFIJXs1bEsp
oDc8/EjeY5gyHdWNhsbvF+frK9OQSSKUWXP5GG2jOL+xWaS7gu3i0levx0Dn
ORiqSVAXq2uZYRi1d4PXe/XHF6U1m0qgv7fm3hPBHC3hq6dVJlxqc5veRaCH
ABwIBOqRfhNFs0gfoF2/oqsz0DDd3fZyjjOgTRvontaTAov7Sd/WJ1pzioP6
cosDMAmBIBTAFbjyTbrKoF7tYJskHoU6JTjKBopg7NHBbx2DsjoFj87AIRCo
WtqMWGxyETS+K4fzyyu/tAeMDetdY9Fyon0k3oni0+xyXr+u+heovoGG/TQm
zk9uQbLfczTbtqoeDYrUTxp4gd4IzNpFcIGcJpBD8In4JzKeD5nzN/J8oB0c
uFQynphkqDPERuJAmcM5g/TvL4UTOAPDBlX+Ygw13/pUe8mc2c6NRgh/uNbC
VsrSfA9FGPpMu3NXFaIURZ8W5RxhDSayZ6uo+ZZG5XfZLrfAaYf5noXeVua1
sik1cZDkfceP6Nbi0MGncZnNCNmME4mOp56X8cZwDHfgdHDGUpRyIXU1L16W
yb+wam554yfddBKFQtQBCfbLlaYiDQvTugaspw5eL/6MCBeZOve1dyiSNxSq
KRgzj9yo3SIs6j+pjM93CziwLjYlaoSsxI8rQAU1M1RXs+F6YVCkCylT9d1P
iVgMWq/gQJkmbRePHRo+J26uai+zP0jzE15hLXIUtOb0kjjhokY1zkQyg6Hw
A7LtU+WoEI2SEeNzN3RiAk0GJhkVhXjRZyjbiapCsjKD/xJAxcRweB5wbYFr
fmsYqfHvp3ESMtGLMLilemQVhjnbaiRjzFroDPkyxiBF88GE2RxRIC70Zrqi
IsUpwoP172XIGfot7yXPWjUePL/ZxtwbfwVHEyrDkLgWw6vg9j1c0sa3Pifl
gCemNAR3igxwLDNOru4ahTPFujd1whQE6T171GVXLM3QaMVXGYrUHEncJ/FQ
8UvgR47ShORhVobzC6/+2NPv6HVqybkpaUIv4wReZp5nqUCKrLSVlieju+q/
tQUKmfDfovTu75USU4ONOwiKdZ1NJnDKRyHoFnWN98kjADUV3fHRXOMJuG40
a3TUSUmgOhilk8A6hYbLBCymFzbqInZXAIoU5yggvSGwX2w2OMRWE+Tq0epW
kIpDafaMMtcycCCOib7ynMqRsVzvBrdIhiQ6sudRYbrFljKleoZhMHPFrlIa
SbSMmN+qZM2all8sUL+YKlxEHn56ZZ1M8lW43ZtM0EaTCm3GzUZdcP8nxa9r
mHnI654kCcP6mytUlxJwkf8AApLf1RyfgKZVBwjJBx/JW7pmjCOgDWZCKoa9
5wRbhlatMi55h+XowiecEyPgYuSMAXZVvRiDczd0eFiUcVICJj40lOHmlYiC
JaxBFK+QafwB3p7+4Xqa6b0TgoHkKFld6lf1w2PRtjaxApzj+Qdq8QG6311E
ug3Pq4On08ota890akiSN6aZNgLuwh22TdIL/xTGK0mhBPFTlYPvYkJjadFD
yW/O2KLdHGewq5myEyADJ9RfIt+uXmkFafL6581URJNofVIv5JbejsAVJxQN
ApHeD/EdBmq18tO8t9D9KykwPlsliQ9Ky6pXPCucOnDSlCCyriFFJzBNgPom
gBRbkyYlqsXgVMYsgQf7DjqAXnhQnNH5websGzbo1QcxVYXyjyeFeysbCt5e
ibdEfdGJjYLHTN3/n35kBKQ28TE/XuMk9EAJYDJ81/6yjlH/76uuSToKPEOc
PZLfBZ6oAFaTipX0Ut/6kRxPtw7pjyLQ/B4M+p69Z2MYcLJin8jnWMb1LBrE
R515SvzbP9RsZRRv9AnFWdnXlXzEbzAoj9fOJ6o00pZQohSW9btdZ9LXqIqO
x00oSFKNzavSG7Q3PRR0EUNOLlvqRezQbQ8o0tFDGr6+fYM6pMqLMLCG/DMa
8I274ZjxAKeqz0IqJQFenZL4iaTQmV2/Cf+7OTsgPM5zMhIiMD1JGj91cJr6
58OumFD2+fgNl9dIYQxPGJ4rqNwLPofH7opHP6U4Lo72gd5utgvMN8nnt9VB
M/vjp/K9QzFqM5xXTnwMil9h2GMU19rQFbcxSL6PZ01RqqGpi43yU9la0tgA
g/258WqN5Y7qo1aQDfZdINkRFTX06ZdqZrB9Mrbc5XWZiQqjjAVQ015tcpnP
qBtEYM5QIM1W2TzqtB4w5fhW+PboT9k2G3k0kDRjDQoo81G+wTdWS688g5ew
wo3uN7JzCpzcLGg4wnJMh06XvmILuT87mLYi5SIM9Q0hy8JDXI/JOFpA5b4D
/JgLc2raMxQMJ1FDBu/cnoQliPAjh9dDuAcuVwVXQAKVWZTOEPhnA0WHcA3X
c0AGKrsR4PzhQi1NyUarLWLI07ObIVqKwK2mJkN3YJhgdDmGWEllnw0fX45k
QvMYtwSJK5xOFS8Q79gFUh3Ir1OwrMtbJALz0BA4q5RxbBIC64B5fYGQG4am
p4YYnNxKc26c1vEz9+04/c2UhvUSybgWZmorYKwoFHwJsmmYxohbY86CnObD
Ql3hF5BUiXfRHNWAAGuS6vbjME92xEbpRJgiGiMRkA4DXdnto7gb92H2+kTz
OAvjAwMtkG1rqe/5VkWEx4rDJczlN1ZbOymRTA+wR5hL2UVnYwYNXngzXXZS
sKDiJGWtzly2CbCUox+08wCNvtlrQnVy2dQ7p7Q2xeRqAk4ECgGiMfnQmF8s
dbLMCQiUsgsiYudeLEnxVGU/otfF5BtCAeOPJpHvW+Dtoga3DcYOewjM01FL
TgOWSOoLb+L6Ppc5Pj85suNXgX/rMjTvaRxQGyxlq61UyAqn3wnQqRPNZAlb
DqGyv/6TsLjfFTjpOeu8+HR03/G0LelishDyjwjb+teBLCIc6rJeT3roXsFC
xiY3q9g8TO0hQT5ZVJCDUSNl6IKoxSrGbRWy4O8BVnWDZcFbTy5Rjd++Navn
aWclZm7st76UH1HhI21fzR1RDsrHKMgHFoRzRJSGWhmYVojOqucsv/sJ6bJR
BUd857P2aekk/hnCVK8ZTro776gjsTPot8FYuKdpBSMyExRbGji7odmFnsRL
n/1gru/GIsAWYxrfOiU1v/qcpCan8LGxO/VUA3AZdscSy7Jyj4Xwj2WE6qqA
svkQ/pXyXgyZb96X8frtgNDAISpl9ztdTv6ofvP5+8yP/PJwkUDrcL2qIg+A
T7hCEENBh8EO0HxXA/0KxEj/8qJJKWB0vKXBCIbXnDqL4Mw0HR21uovySKhV
ZdoNNeN3wL4xvbHIKRRyIxNW574ULXfJCBOLN3ZHoRwoC6dY+XJ9ovt02YWB
2ZmKdIOKbywFWFKkRhmoiY8NFa9OeDY4lsITE5PYXTw5tlSZGBt7fV/oqUDi
oKghKH+JJzFVZS/mi2q4eEONffJMHpC2QWiXnFbESPZ8AIsjzOstpNyhGvKA
+t1dPMCOHjRAsGDp0CHBJg2ZsjdWC5A3E44bq+xXgXRnJc+5LyBHG1+crxaj
K35SCItM+Bi/eEZok1a2/mYaNqo+yKuW9z56xxCccmNEQuTQ44MhT/90plo6
2Q5F8rhGDSxlinuLA48iGFqPcgBq3E85XiSP3KilRP7U+u0xbW8ADMO+Erld
5Z1yo0nNwbGrRdjplCA2zY4EqqyAwmB9zcVNKdqtcA0jbyvaMFceW4ELBwjB
Ckan31jnb4Q0B9a72DT1twHRLRGF2psckX5dxV2wwPiaqBi4rqF8iuOyk8Ba
ptmr5WUeQzNPOCZNu49+InhHsZBOq2hqJlTzn0uRahvf0aSguArnF1oRRiS9
aqcJ98/COpwr4nQXs6NE4FeFWlJVoeEqegvPimzmbGRh0F0UE3EwzBTfBG6+
2NsT9pcmIiHR4ydIJyt4yWzFzZ2/YguI2513O9vL5j8KHXKXm8dHVRKM6kZG
zZPdLifsrpGb6PFACiZSZxq17bHtekbi3ZL2bWHf1NAJEIHiRy+O7DsJ61ZI
1pDpdZrK5fiYBGcQ5xeGH8BAQGyqb3JhX3bPHMOD0gpJNUrm6XYTk/trwru5
CzeKj4NiUnxzvE56PkXslqt+GGct2mXalOzDtlx/nAQtuC445Fa6HyJKXa3o
UXLgqSnAoj3O01IV08ADhB6Dt226I5QgNXuFuHolKDv24k5a11VM1A3d4lDC
PnqnMhz6rMydWJehFYcr80w+S8GEF4HrfWMSxAZfbK4Z57G5r3/A3hS68Chf
MCKUeOi48cEXoS58SqIE/7GDz60v8eHXcXXWN9m2DHwyYfG0yVDDBjjPDhX1
xyn5PxfV0ePR4Jq9e+Q6pYYlQXw+mEwGadPJaufaERX+6ePCe7JRwNieNC9J
nbnvXYwmKayjP2/c24YAZ/FVOtKpKdTBhDPHV1ajtPudsytuF3Srz9Q+lwI9
E5qpVktu3xaNt6n+PWhbepGVY6L6yHMbqhpE3ghSCcWbwaDgNMSnsxJs3eS9
I1zHHFo6KOruOAWD/ZExdlgm05KaVfvAOF4GI1ob1QvexfyUAoDPKZ+1DdXa
cWGZxxA7YXB2oq2TxEaAtSaKDwRpNtcmkO6KaNdorgFHO1qDe/YSzJIrFB6F
0xvhUZ9zkP/7wVJRceadk7pr7yXPbz9nRzGaZH94WXyEt1zWr/R6+dYa4iJx
+yRjci1o2J0cL/O6J4JLotA3tEmKwFOueHk40JwRDU0H3bLTxNVlp8Yer3iV
G9oQhFhWvc7H+R/0IIsT35GeRQggfWLjwXs1QWqoM1C2+0/7R8SIo7lzEEkl
1g8xvcPk4ci7BmCmTdNIW1kfZEYvjrz54cR9yw7du4VhKab6cM1cQp8F3jYH
tXYlbsUf93/uFyrJ+tXmDw8b8/QsQPmL0n9Rnnvu5T0toWgVFdxEYqH1a/fn
TyxnL07MpR0PvtWhgrcTcTCUCJ3r4IGmTTKENZfIxrMCmMurwT+Iw2XE42Pf
htVu67Dc4KqiPM1pb90y3eTlZuJvlRWD9BCH46/gRUQ9VqmQrOVeSuxQNehE
9WR3UC4wE1j/gm9L13b0RlToI1lvCqAflKOG2NZNM1TAZSDp74n0PneEpidR
4h+x5gJRaD84768+9dg+2OkUbqW4aZi2lltPEPFI4SUoL9sh8TRsXSDEP0Rx
2QPdOYJL1MlHSpiyHsOS8icaNnmND++jGMCjX2pJ3ES8Vxxbd+Izp9Pk6Vzs
FA5z9NPplIdafJhZilw9eXXro4e6caNH5D0mLde8//pweoV4leEt6BwCnmJl
mEfXX3UXykKO0lrEoXZVP7jhUs0Gr73j6dRrFte9ahuS2fjpIRCmo9skH07L
QpMWGzDq/ogj3daORDHdSqVlNsCnjkevxjLP94TBLO0cqHlNIod9EcJeriFH
cHuUUrvIAmxvz9xmJAmTv3zAssGaC4DN56QDcKWwALcR0g8xA6/c+kT7zctz
8IvufYFqORkPrtv3X51dbPzZvn56sMstq2lJ1feSFv4L2UDpxD+Bg7DqlpZS
wFCFtTTcFMCYfd28E18CoI9Hpttp0btDjaDCM6N0ov9Y6eaeqTkCV3+a3BdS
YjR+vYpIpGUe2K3t8yUrUcXYdhfXugGOOjeaKEUv0pvSWPi0IyyhKeOflmEJ
bDKKLXjEcXq1xMnIlPrnJFnas5IFSEzrhyVLDaUD9Lo0B4nCnZsaFuwvYIkY
DbZBm3tdkjeTus51Gwx6Iq9m/r95t0YQ9NzvhxpHgTB+WPacKsWwR14iM5lI
Ktb/xAMJd0t0CZAZw0oBXDnbcNZngoe1cIP4kWM2xMEl1nJ8q48laW79wkJl
wKjGscYsra3haqHBE+OuAsBnXA8pKcOHObOFU6WvK+wh5HDVBDVS82XOBW6V
D2L5zH2ZQLvkUda5TScmarzWY016JFV5orMZP8/Si5xF8h2tKrru6rwFwIcs
RquJHYzxNj5odUqK61+w0DPIZpl3trjpN3AbEQ+CsD+Y/+Kz8IUe8oyPfS2n
6gDYWf1LRQQ3JI6YMFgC+FjISmn+V6a+ku2Q9BV6mgp+Z7O+CF+9BYNXDM+k
YwwlqeRPKR4hH8HhXIUtTyHJIWdyoQ7AQhIX/74p/yynMq+ZryUpB7LZpiM9
IO+n13PTFpdSCsOjx4FW2/AnxAK/2dZTPoyMdddt9EbfQOk+nuY+pdIXKotw
cVe5q9EQyPCpSlnacWlOddUH5K6Xr55vu3GaqLHPaLloJFqG0R6kXxmBtYpr
xHSoDzBOqYQ9JiHY9E5Ov6XXt5nXK1Ku9MyVWso+RA0/hWi/TawM6RFrvunj
OTLO+iiJh/leODazfn2FP/aLZdGx2J3TDCnHnA8FfCJzHsqaEFrQqyI0GaJZ
CNV7sN88b+zDJRNmQqCOCUcsbqgIeP4ONYLbv772+gi8+6lQBnvjLd/S0AtV
r0/mNYR0HW/zq6WyHVCKPF9ad/tgkx2odq1yXpUsry/w5s6Cz1dJR0na0UU6
qPQQ/LMn1GFE5zUYsQSIAINa/sMsabdt8Z5LGz4UoHLlSMNKLWif09++EOJE
NFU/qSB/D/zNQ8WkdwV0h/M39s/HtWmEV0DKID5UaSrZuP0o3wJq8rbWX62s
m/1sZibB8ROp3pQjOIZCXM/IrVERRYYHjkxSeMdexItRd9sDjWFn8geXSRck
HBv0Vt++bMqJWrZwW+QJWT5mgUEwqHdKNYxO0DXutrBVhKlnMv5A1iTtS+o4
o2wAx13qxv0jSvkadjN5+37ocLNJfFc828JChNFBGtoXxzP1qxC6C0tDZKgH
azVNTXvZ2xOh6AO8ehZa++0tkBhHlaSZAUzAHjxePpKp5VgrGXBJrOE92N1O
TxKSRO6K52cxF/+kaTjnM5nz7DrXbiN7Jc0R49y/6RighseavjEEGmWX8Zf5
qBK+1yVYhUlOMVa8N2KzKO6yOWmAK1dUVgKQyuPpqL1iyMZl+eBOZBHfe0Zy
qSkSq8x6K4GhW3aUM52V3PdwnrogYLaDs2EPj5K4YTI2OBj+1GpkRN568lBc
Rq661Zqkvj2wLcdH0TkZlEXkDN6K/QenM0pmXwKxlOvjETOZs2LN9x3O8qu8
dxaGmCERhaDHa/FCvO735u949Jno5PY8/MPywqHNqLwDJqPqWtU/M1KqCFTt
1ezhMWoSfEPqTfcwGNgjeDV6OKril3smMdQD80bZ+r7n/1Vb1dojSSAavH4C
x1oCzBgpAOuuD78kEc3qoiOEIYjebIX4HU/VOA0PL5pNFmXftVZmz8O+3mIo
PcXTa6Fm8vlZUdu3TnOqWGbRzTCRTPKWPusuQBdlXqRsNwun23UzvKiYosts
K5qmaPUVTAfk9w23MwZenbYfY0lqygZCXm5W0E3idw7q48xAWXU8t+4+noSt
ouHd09h5dPJlxcB0SSO1FWFQMnaQpa6VTl9iBFL0a2d0sJvZToBdkH0cPrlx
ZaGWN0letcGsla2TL32SD97q31rgeRbW9PDVGFa0naNIfB+sqaMPSTs0kS+Q
nZM7p94rfjjkvLpjYGgkCgfQkrPP0olqm+hwm1uOI4zoJbheSaUv7c5saZeI
PlH9ysQZR4J8w21et7EF+lzHYG7ZbyKo1E2fIukHTqhwY3hWUHzuNpxjtZgn
LZ6sa0Lc2zEWv32ArfeAVc9gjUssOjMcbDYpuO/mhUsytyz6Nkh0SdI3FFJO
S1YuMX2zI0iXRL0bC1lFYTniR22ochWQ2eVkToamwHsukKNdezHBisCqRcfS
PFIq2k5tVzsYkieaU8J7+Lx3RHekfm7e1+KGxGNJqTMkgzPFdrzKuBbZNYEL
+hfqj9NQF+Fevf6npjdHHWOCTRjYQXgqQ4EciPcE3a13O+8dFypBmo2NIKu2
DnM89zyRM0gD2cQfshbFObD3V97uYdvjzRis5Drf2hS+OtOPicxYhTy1uRjs
GsrQAET7+9S/BH2NFcNezTbBdVwr9Kx2AgDBPU1hOK/Ed01lhyAGMJiDYhvn
qGgEeHZX/9tsvF18iWA3QjNL83x/BqAhFBjVQxPRkjpgXo3arNWvafziT9zu
zglSgwkD51Ihb+2v1Qt2+9MKp6BukZJsexs86y26DpMemKBDgko4eXnGYx71
4vnOitMM+eeeNXrW1+d0DJ6NmZ9+ISm3j0PtuGdOQr1me+FQbpaAYRh0T6ps
3A+dp/GG3LZWRP7xFGSUtLBB33mXSYYy7j4KIGMdCe+rbuFv0qgfaojAs/6t
iefarlIT92DVBhiDDIJwbkMkh12i49BHw96Xt6YOLtvsZsLo6djUTg2zY64m
KRUBc7Gmqupwwi9TFnH11A2A/5gOkZRSkqKaNmLTQeOeoGcBP7UzQBLqN2x9
cJwSF95o1swQzXjSUTvTP9dLCeIeOZ0RM+Q7aBmPFps3atfa1JmZRp36ccyc
Wm89K2Yel7wk75Mj/86LAdsQ8yEEOd1W1ysDcWULtxkY/Sr07tE01n4o9M0Z
avSt9WTOQVZwYaIvj69+nuLPYmG3gnw/0Nbg+0vH09BUIkvFD0mOCBhZfkSW
TFfG9r/qLSnipYKsb2Z49VujfW7vfWeVq1CPaLClP2LDhaZZdIQu113WS+93
2d1s2Wji/K+BlDejZ9zOkeB8fmMlIbRfZ8iy0Ee7sAXw9SLUlc6pGdTzzpeJ
2zahIbYEPk/qsjLgSbXvADyN6zqpzt6/XJVeM3s2/yXWU/JX7Nqvuze7/9z8
BxahQnnIwP3qXe0Bx+6BJHekCleK7jCY3eymWEmrEX6je4eas6/Eb1WD6mbR
EaSio/IwDGejFtdD6ZbejaY8KIFobpiqPN9BfXkn1XxtTAp5dbd9kq0UUhzN
OsJojf6FhUV4gD9nKNwRsMkMMkkekxqUn+JsCHaH7Z+iK1g0Fgo2RPSlQ01n
hIQGoMpUh3XwkgfkUCeq47Gr4151nL8FwimtNxEwaPORpNnjhMzGMBNqUnBT
ju7mZlTsdx0/R30rPRFOtruSd2Xvm4Yr01ydiAjYTnBlB1VyDaOrOggb0iqg
B4eeHRv7gcvOXydA2DJcylJx/76nhoJPaDYzraOq1GvyPAdCjcSbKACd3gfk
4H/a//Z1mjlwqm15EBVm5iNNcwmaczgVNtspuc0A0VpjuLKgTU1H/r68Uzj5
lB0lu1BsECK0ivZipIj6SmqVhphQ+rawmcD4W+NKv2zlOElNdk/lMW/VdQNU
kR4g9qq5gFzHtHl0wQOwN/tdocVemsc7eXOdRzA2RasOMbSeb84EIJFJqMsM
ACi6kiA2rwIo+HW9x1X/rYQwSDxM6I6P/W3LhqXkgqpfpyKHGUtVaV9yB9XD
riNcj0ke5Jbwk94Ls/UZa1AHR7zfeHmRGCp+kkyZJbTs/YL6Ei/GQ3RiDK8T
UwpQzs3japWkARWwcaC0OxuNbWmT82MQhWC//jc2NLdvrzjztzVFljpGmr4D
ArVXfn81xWDlELH1ySysSKNHBZcWvnT2W4joCGGV6VZx6NiZyUXZjezfG5Ga
61c/IWUpZp5nhpN0+wQZfq3kmmAHoB5nZOXUTzbSBqKR1VDm/22h2BdVXzES
jIBQYqFepjXFVYYNMdp/s/prFiUZuZtuQCZ1Va6k/Js3oYX9DYiqL+e/L51u
9UPkMhSwkfMtcIwsYop0FYeYGcc+vrOEq6+eydkJX0GMtZnsPArjYN0H/7Uv
0hXLLOHulwLzK7DMh4o1VMWEbt1omoIT8LG03gEgGVff9gH+svc9DUCUbfwe
y0BKrC95PSLa9rPyDwOsc034lhavK2SLuXz8XUvaW7o+tH//ZrSaA7c2ZOqt
+VtfRFchWmTgTIVHwAWo0kuJsBacQ1WfSyoCkMxJ46aJjSQeYyZRGMcb+SxH
Dv1DwUs+sU8Q+CAFXCwZGw9SI5PO8SRzZg9K7XxV4fR6xsmD9Rl/ppdbXjG8
WPqjDwi2eN9qK4U2yjSjJ/cVAvl6WAq7UgNmo5w4r3B2sKsOwnkOL6EpchVh
5nVgMn6/t8S6Qv2XVkgdFp9GzXIU3ecXSyz7LqLSH+AgtVd1scI2rLhwpInF
uxw/UvorS1gnOf6/XWgApTrsNUDClnqUPFS7KyzSYJGJbjlOvJcJv61gYuwU
S8wwJJ08f1IHuoQrch8pdcsXTxQbrIoNjFaLf7dTwu7G/niEaiHYn6tBAjfS
Tb2HIfNl6VM7BrjDwhMne82jEkSNQJJejskldl4IbL6b/8KBVjlHF5Nyrlvs
abyLYwy7KneJNbT3PtbC7h3i5YtxPQ6KUkVkK7Ye+eaOjb8gBQKl6uPFHHk/
+HiKZbhZKeVi8xiDtDgUtQ3udGi/3ef8IgJ/bENLUJjMiiisAehUcqV7Hg6I
FMnLIStCPtQKY70dCqn+UMj/2rlm9lEKHKDqEkYmGdotQvKQhJwtrGehUY2r
VKg6odEnAaChuDcTbmt6fCU+l03xKXcxjchXUlaEOWm5CgNaeDRQUnG+K7Px
MQx1B8httRra7CAu6dMVqpyYlJkqs7ZVYzyrbnDEuN7U7dQdbMlhB+9QPJkX
Gqn/7UgiOweXvWWsW9GrVxyhvv3+/T34Wi2NvEpkhMHSqA61yNfJIhpphdL+
qWfh+jJO8GgkJDOeqPi+6YuT4k2Q4peyuBG/orjcMPqvqMYGUxM1TYQRKO4V
wagTNFtZled60g2sUSy4Isf/WQk4WDP5TdHAFypkaL7l41fC0aJok35CdaUk
H4GXz4VY3cIYQo5hTRD82wTSbWhOgcsneWn/RYSLliGp8PC3VDF6Otf5tvMi
kzEykXFg+6eO3sJq5GZZdosIFCwRsqwCLHp2H5iguxWSLON8nds/MGFpLag0
p1e4EvlHcGpmlgLp18xHSxeHrf6CeQpsr8Ir/55GHp/G6qNuwfaPcphs/4F0
+ENlKupLMF3RSM+5MyPiZiDbO+nSMBWS2Wh11M73wbnqH6b6h7Wswo84gRXl
1Av+IClMGzFjjwWDjuuj+DxeOcb3ATdevbOp0edkQBiT38FNC3JAL7vu0ImP
bJjSzon0kTMYWtAtZ7VyjH35rPhV51dx3+xYfvdtTHGRfD5nXl+oauNhtD60
vlVtTQVMF2UnEMAob0MX8rMZ6Hxo95YNNb5f0txTZfk3uMVVaxACR8weUvSH
UcuU8VsWevTvNzqDntWGl9w3ybZNjNkhnR8d8TEWW5U0owSqELNAQHc+n9Pr
MOpJ6g13eXAPKHu6spG8UbzHMSm8HYAOIEKjOExw9saJ9mceazmcNVOp6buj
DKTa4NNPV0MhDsTImmpbCEag0xzUbMUedyH4ECZazElZ9IbhZca4PCrphNvb
I32z+U8MG91sllaNWE+JKnKPvXMuU10jARIg+Zvu1XQbw5AYF6b7l8Oqvq3p
i5gFrTFrZ/Zw3a2UrPtglAcyMYAn0u/FMVWEPJzDdlr+x4lptKnAB+VsWb4m
PmmWJjXWeVQ96+6caARaxZQrZRIyMYzjpdzT+wdgSsAiDJTaALOsB+F9FQ3g
EzElcl3XeZ8vgmLYtYrEIGcmWuSGoiJbBxUCl1CUu9GDmWNGwoVlv8q2Tpbz
+NjMS1ahlCdaA9ROmEiz9pd2U1lDB1j+3XdNrExLx/y5evtamVd/L9/CwGQY
9M1Xct49WxZxm7mqwmCW9ZsYS4OCdWkgVSXvEBHpy1J8zbf7U2ybyPZqKPTJ
xCIKP5edTq6GuYZv3RS5x5kqTon6aDGpusH3A4/fe5xn0qmsU18OlOfcE293
AEKDk/E2il+lR4SN4KzJ0lU/HZh/Q++yMuNi0WIJE7ToE1Cpq/OQcCi9nPNW
WOKAijlC6VmqqC/rvWQRUwp/CwcNlwOe8R/83RcmrXGJZ7aWB0h/Seq9glJY
k0RdnkSc3SVK/vnMtD7dT8xbSY0LWckSCZJt1NT8eqQR6qc/YRfpR2BY1C8X
JcyiUWkzPRFN8tnGiT8DjCUn4KY4BBJmFeq5ISFWTbB+ukVHI9ZVb836yQVE
WGNBcmwp/2A2j8pnmYk3hvKTuHSPIXjgZ+0a1oeghu8b12DnfoJrXgg1XsGS
MI9fh6n7D3nN/whP+JTUWCbqLvWAb+BnYzur5R/u4AhYtqvfM689yKg/J2tH
LJbiT8k3kWU95hwg2PYLYWr/ZbCgtfPYy23XVxsjpWqJkspyU4Z8J+fClGs7
ZeoeH0NCkeIGAIdGn6qKCDcrSZBKiZMqixFFsUMpDIYgAhgvvOfiNik9QQ52
y9gMlTZpZ61f6e/HUf70/5q2aUMTiIJnRg/9SlvmV6fufRAluM+GFlAdOgcr
KQyjp+SVNmEEevmk4X4vPYmq2ksoTu/2OsNirMv7Y8nMEaynS0xJzjM7AZA/
N+ZtUUsMkMjeI8HxyRSqx14eKJ76hzHxjUzI37NbCGYo9LpGRyHc5ERfndEq
DkhAKgLhIsD3NFdX2fafz0yjoDWkLzMGm5ZVnVcubQrePkKPTa7EVjzgyb5X
BW+PWcVccNNjeYJJLqpDsu0GBYPqtOr7O0+IeWkTx9RCdCd4nc/xE/3ya6wQ
+yVC1IuDaY/z43ULAlC2zksU0SpAcjp5d+YFr6nLB9LX3vNTSXRrCIEXgscq
h1IjDGFXOR9Rp+QSafkPcEoRSanuEyEWE1fv1JAEm6BoMSWeoEf/hM8m8otk
8hQVKbwfxrNAzzfKyds0vYnZoqBAqw1w821cUlpOzl5Ql3KLLYa6Sck8og+Q
hUdx81qIOn79YOvkIhH/Hpmr8YNv02gE3FX4UkIvv0NqER7NqDCikfeIyhHB
jyDbeh0KVf53IDHoKnIbrCvffS8ezu6dLvfoh+bh0dCzpwEFOk3bNgpY9ivd
AWWEEuAHwu21LcXDue9JYrxwJW42XVByshCCoyO2IKgBFKQfUz0VHK3i7QRm
5iVbDYfgUcVwSth+uBVv1Ov/ruGZR28g7J5bBr5aWU3xzwDn332A3lr7vMT3
jwlz1EQ+gjIZvZ+9TIkKfSDBW5mU3a4wyaaWDWv+Bb1OxgbMdDETbXuDrf/C
Dm6udKuBvwFv2YM3r6LX3lgo+2ZhmQ5adgQH+uo3NPDeQv/EMuZt8+VvnOko
IQr6VHndHvWiF2O9tU0H5JnIRWi2+HU+0YZrmMqVJbyyHBp6HF4dR+duRAvV
MZTngPp0gVI7xStlICxpn4CNfhfKHk8/vkNM856vD3qFLTr8ivKrlIWFJHSa
TAwvPhYVnjZa3RJHBaY3G7yPVgIvpbGQIoElxkE3t7KRYJokwq/WCjT0H4T4
9CefGYfCAQDTeUBFimIGg3Pudr+Ovu9EqCxhBfICq0OSSOvt9jWBXxgL3hnu
S3X1G0ZQ9Uxs1anGc36ujcAplKWrCmLJ9eiwCBNOGSiByVFSxlL3s4a6XhDM
rfXh8gu4CwC9LotQOD5RMVi2so+SioJBzgFrTnjxoTUEocaXY7taMrTkwyVc
eZK8XPVPRkGznZKIne7jrYJ7ylR9gDrhgKN3+hR+LXW9Ubv3hcv3J2SJcv8M
NaNsnFcocflJ6ieePJ7Q96aj4fsRq2J/FnjyUtktKfaJ62FvujjM0Ft2iM5d
njkN2YloQE3GK2LNNqOEdU4KE17phCBtV5ifPgerrPLyLrQ66HB/TmyHRWVs
4O1Xdcc7ZsZWvc+etV72WRIwxt7R8xmXS0nH8EwJJdHKk3L+zj13DZ7K++kV
ka3NfrICXxKr7YBkC3t6fMdy9I6KGVa+oz3GlXI+yfAKD5TxhoB/gbtLh/Tv
0e09tuCDRZ4TUS942z+6OAOvAG2++VxJaIs6W1BDS4lEljSXgJ7T7y3ou2jv
sOzGTHRz0lQRfrSbzvjEG2b2ETAldrsEopmZfyI1jDq7N8SR5YjA84gH0Pnd
Wm1IM6JP/qeLLDy/yoRERhgWqPkYZ3bvm5ycuxLGQP6iFSHgvD4bZRGEl5vg
dL2yEu1dwJiOLWAmPQylOJPB7wEwVCIECzQG+UBfW8uy+K70NIbFk5Dw2QBp
Sy0tUzQujTUtDyV3hPs+q0QrZAPEZsTI1Jcpnb/S+hlBZqzDu2Jw4sqnfeJu
ObzVr1ZR7Nc4j2HIDP7TA4Zqo1EqpkhIhDDm7jOFIfdnEKhoKG5kuXpvytK8
jO+JsiOOHcD/Cdg/4b+ee4PE6Srf/TUmL9r4IUTruHonfnpjxL1uYLUEMgD8
+f/XIdsakMW2Eenuu56SjKNYtrAizK4IXYymsS+BKNU1PvYOHju3voRWhwfU
wpx9iKvSyFhXGP7WtBFkAKI3j01LorkbL28VRF2LVowajrNzNJIzB/IIkWiD
ANoOOe3El9peCEUityM1vl+DqYENqajkETzTTcs85eSbHJCSaFVxhW/iTm5T
gOUPtNwSGdCD/2Kj/zfDV4+8RlxHIfEXb4RQoY1N8QjTJu7VRiRuQQwxucTJ
6xP61/qb9YWzu2Tt2JISmb4t7uFq5eGb5l3a0wJqqqVV53/ZpFIKxpO2m2bR
IuWHp8+SrnV09Gss5EmZ2X2JWIE5VNLLvVUCOUoD8Vd3wlL6+6xMB2PE6+kW
0+d3pbTEKxC+6IgmAMnTdNQQFWrOXpmm8Ph+wefVHoeAahzMMs8iUIH5/wBa
SgqgF+BnUX7CP7xn5WYymse+XUzuCXy5sm2dTcUSkgDl80exQhF0MwowBZNX
5H1ZwLnUvXbLvmwtxWbdw5Hi3cF1DBFpxEzs8DSBCuKWYDgTVEP5CTrl3b+d
8xS8evaVoWbgJ2ohaMIFS6H2E1Yj3q9/2oPLHg6Znf4aHV+yiTf4BkoOpSZJ
gKr8xQApfhf+AaGuQhX466ZrEX5nfxTHawAUzWaI2370LwjgyG7wMGbBqf2E
SS2MS1ltaf/WnA08cmCAFBuLJ51K3zjkyG+ZRBcQfiJVv6aonNuYSirWLABH
ThtZ0UoQctlXG/RDsRY0+ztwtWn/gmTiUSH7MVIleW97qh7YCibopL1v1PD4
NsGynuzZgVI1eFumrJ+PyJImeoUzYHHazr1zPjW5ra5UL/PKSyb6xmppp66B
2bYLCUicUhs1mPSldD6Q7wl0sj/r1zv9qnoKcUvrgvEzRU/4bVgCIWZPpmjW
ICo4VITPq8FphQMdf874B2/HbuKO/V5bVLX/l5TOlcPuP8UnB+r/t3QD3cWU
Wn4pbg+uIyXk/JhzwEcFpCZn4Z6GKbnrX2tVJN65oy/oq7/aHOx+10rkEHqV
mS31HlZT7IJLcTSSIXrVka44w7YNB4rJRutYNITNL6qJD2pqX333lGDXyeQs
R6/6X4gQRaziw7Rd9fdu8tMyIfv9sUTJytoePZJvlJVg5dXRhC0W/yfuL8oe
JjDpPNua1ZDn/yCxsI1cFKrN2rGmL+eKbM1QkQts4iTwFr6PNpn0xFbi1hFq
vTgQURJDoKE2s7huJg4IUx955EB3VOiDGroHuSTn7uQnfPAcI+mrWr7Vj4QX
ABHmGBn/oZEeGOdyt+QKsmAfCVEpS6iRiEsQIsn4X/g3TRnL9xhJTYENcldy
CZAuO0mPpiltpc1oaU0rTpJ04NlIbpnYlRvBM2wc8bHADTc1E3ZPC+THVxE0
+RDXSiHvPfKCbE5icX/B+88FkIygT8DWFXuV6sFvD3slfJ1yWBEjJpCfpdiy
MWfNLCEZeabeNtErVqqJPbSQag87NeSg5DaB3Yn1TK80chIWmfO/nAFJFDUS
MbjsiNpQiZFHyzyLIZ2IAjar9JP+9EqIqgY2TINzBZIWBlHhGXMVQoj5tATb
sf/oMvEE2F9c4oaMVNkVZXbTdrMIs8+kZMezW4AU5cwzR46P4tdpBqfutJP4
LhEXfl4LU4MbaDfadHAU6pFa17g/s9537V1BVA9jI0q1qmylwMqfUk8KbYhP
jFHwOkz+1Mqa51POzcYzkYV7A9i+bBTHz31orJ6sRdRjD49GIcuH4vZXB02F
v/fbbmBvwU2WB58wnQKA80Fa8kNUsfxQdNlIMPtna6y4Zedow1p7xiqlMPuI
RQ86M4rstj3c0I5iVTKHuuNds3HzO654R0zCemEoChpKurKKDgiLPBwNwilJ
qn2zEzrF/Q1lXNuWGx8VZ6qav8FM69BPqz+VYgzKDhyNxca11siV5DXB6R7n
OEXjwv8c+v8WZQur8Kihi+fUsVzx4S9DsTAjmVg7de8IKAvw9rtlJRmxVM9f
cjzvkpdakNTS8F7xyq/7hK+AQwcTfIsN7MnWqgV6Qmh2XEqWBZzKSwG8WD+5
yx30aYOgGHqsbLOoFPQa5rhUwywSHtha3Eedsh8/CvG4te3zcInnqy0va+69
6vm2oyj0XurYwmvMBljU7zolBhjiq6yH9JAA5CrBfAm/1b3kWsyr1JDt615N
RNNwH4JbdfF3uOPA2FZTxhNZVt6YvzgzyeNImw8F9AC+RJLy8y6J8xQuIfGA
qP+vE1ynVQsMIctUtYo0FcFu5jEzMvUBmgoOMUMeRD8OWMysXfYhcwleKuTu
PwfmqNfgWLBB8MVsuP7uDqXtfL+sZdrLVY0OJMnRewZXAQ0P8XXn9ra0mPnR
EVNpfLGA+wcAHy7OUSht6moIlLuAXgKu0m6AjZasgg7UQRXfRLWhrK82lKEv
qhwFYRxa0GOsBuN5ElfZh0DMaI3JDx5nO26WH4PQ/20Q2qSUfet0BAacQVdO
jb2UBVN3CHsEQQIjk4GSk5APiYmIVf25mxws9WQEPusLxuNxswFcdCZdan0K
QdMLDPVvnpCSDCxjgr/QaW8YVZNMs63OtPrNjhMz27ex/awiRxB44CGmOz7N
tD2MzbUeQ2F1pcKSq7F+YvO60lsUibkKLcX02xOY13hEJm+drJjT76zP9ugV
L/VXZuTeNgezagpUlsoavbQ1Qw6oV4zQcZ2fgt8LyvZusSaFMjiqeM2GajA5
ytpAxqKWhteX1ZPzWrsMvgTztn3BLv0yWdb8XhvLkeG+GzKs+jIPfrfUZ53i
JK6tLcnbc9lVu4HCIiPNdp8kYnt0ExzkhgrVbCo7XPqFa+Kb4Q6AYXKtobzA
YK0YLirE7U0Kx3OKIDxiGEEV7YWV6CTA+MlyiLzeA8xw7+hwFxBgplWM09g3
MRuB7YCxWHfqvskqfm/zyC1xrVfQZNcWK7j2hFR1BSDeTrx/p3zKwKJiWqnd
G1/I45W0Di13a1e4VeCRL3j23MTE/Y7F+e7+kESBbJgqeu8LnUIppTkcaT2X
Ji/gy5lRv1asSX+6co732+8HSGeVz6lbKytlyfp0d00F2R1Y4qnthMocQO57
EPHXXxUG1WGYnO9eRcf9LJk2nRMSpQj8sfry43ZFiA5snV8uWAiy7nulnR+K
YBUWxnzJztsw/yB3BiUpUZoTCFRRTc51Tsos+HJ5asZFbZuJL3cjn6vXxZYB
CECZF2d7XXTw9Rzbr/hCwloHqHsbHCFhLdeXAJVXyASloBRgJ2vMXZC0kGxs
THl22Gkx0aPCqpP7np1rCl5flu9BttXvjlH/mD2zco9SMrvj3QtpgR59VujA
u/rtfAk0h4FPegGXECCx/8vPyo9IqZFBxabyH7ElWHR2u71EY3Q4NjcHrSvR
OrV4Pnb15ykTCVYg2yfoW/IZHQNWSRCnomj/u+2yNNiE6yeU4flPXsTRXhI4
azU8PxLgRWmlOM2/FLBW1lALetYoqs3+QzdtWgMgLHCMuwHiPmYHqn1jXf78
FKTBKWnhphbPGn+QUTmrL1WYJ62N/xt0nR4t6fyesgihlWDj98jGPKxC9L7z
jPi44IW8vbpwBR72d0XrDaHx7aoZSNLDxJaJ1wzMQEXiGfFxOKhGk7Rhc1d6
LZTutkeJnOtOazFnbWlxfiVDF+M7HPxkFEv11LdYQdSNruWE5dQxf4tGHsFh
I2eG7o6q2bshiIjmH/3dqgrLCL91azd8xY0gu5g6yfEUUz03wSMGjefaeT3i
pqq19CL+VEdq3LaRu+heipa8A2E/OBk74/KJhIO+2LmouaMlj4KLPmogJbkK
Fce8oGAVZ06WG8phJdwF4OR87k41GpEGrO2iIB7vn6TyqKh6MrVLXDIus75n
VVlgv1OT7l3nzVeXWxEN34ggazKi58b76lYeZvK9STEVYvEseELxtMoqlcBz
6fjckVtRP5Thy0eYAdhVEY/y/6Zk7W9NpckDM8PSFZAp7dReytl3IJiPbxsE
hVWYLZj5LIFU95OzO4CK3JgsNrOzrHgflTnb5csFj9fSQO8qyqZ1KxywURaw
VONKQP7dFn6GIgGQnTNb0is/jNU1EYnj29sfMcLaQo5udysuV2fOTRWNYH7m
B0Ij9tKCBTP85lRtlUXaudIy6+HLAd3aVButchPZI9pDjGqzbRefoBy0M6JZ
ubpd1jy+MqZUmwwqGakaD0jLO4kMPLILz7fHFQrSCWkn7brEoVUFwb2RrgyI
QG9b9BZkcc2nlIsm7Smpl7nJuB+E1JLfRqLbPT5wdrxqZaSGv7VrccBDXUPG
gXhCa+y6bc62cvnrrXs1z0OBK1JWLcR6lFhkxu3/le1FAip0B2HKWbLZaAjB
lyjB63yxxJ8b/7sqFquTOoz24tjXT+chz453Ooz7DOEZjVHcafp4+RYSRljR
rjTi1gRxcZXD6u9TiKPq56zCKZLWKlPjOsSE3XqpSCe4QUsg99HD4B5Ddp3y
iP/XyO93M1OlJ5Vx/NEtnBj6SLxkjgJDuuEShxo8tpWB90dW5LxHd4a1A3Rh
dSPj9BG4zCmQFCbWdpABNhsd0ezkRc2OF1gJ0b1oM1KApJ0NP1igsEsVuBI9
Di5V+FnwrqkZJK1CIrno/wzRHEf24gpCXQZ6fmEdKRdQfcFvOJsqq6dpn4Tx
vTu/OP1KGBZ+KVMq3/v+Bjpx5sVIcAEno5GHaj/NzYiR+ss2KGnbvWAgnkFM
apCgFNXqQsgKt7MX5svv6WyzQGJye1hb/W9bMWeYN3NXcsbdmi+61OosH89h
rtH1uP9wAlpFckf3hkVJYzF7GESGPKnDPtJsHXl/BmC5354H2bIz16579x0W
RgJ63ETwMjhcPP4FHZpLinmMSbSl7nNQ9zYVt7eyWSKEvXX2US1J3JjLKhQe
vLGLp19qlfPAdwCYlvj1oJ8LJHIVgKmTfDLxMcqE2vGdZkaRMHLYdcJax8NA
AU3zm0K6gFch1uL3UITAp00GrrZy697eBcG4hWhd9VNQ8zeUVloTkQbvwkni
CTcFWe0Y8M9pde2bwWhCOWzwt3akWrbLpoQeFZZaxmw/Iwix9JHmqjq6LTv7
4sui6g8oiyA8QIoZPQgl1NBsCzwauJaT3tcdDZMiK6JDgOhgAfuc4ytJDErE
mMEVErgWIZQWH5CcjXfr/r2FPMeegnY+TOREOogQuDVJJ5VUUE856mMpMYP8
yRGU2Y+M/N3GyuNYSKf6STAp34xFDiXrFCebMBANFEXUtsr0JkYzWsy8sGPl
LMRWZrwDGBVHJo0NRVkBuDnlkvDgWZyH5bqDIe6qvWd7Jvfkym1pZKlZJh91
AalyTDqy1SrpneeVaWq1heuQP18I4aS8Ss/gnXNpy/q7c0WGfZkZaRGJMjyv
m/ZtJm8jxuchEpGIG6jfdVaPpx0zMZA8zMYoDEXTKykU2ibvlABMX9Xo3EVM
yT2Uj4PX45vUQ0jRXkKdqwwXqU7R4b/YAAxit/6YNB1zRTzK0Ljyff6agvIt
lg6djCEi7ciZhh3BnUTXCPgrzgfPGR4/OW0saFF6MP9d0raJfQtnz3A4mkHa
TQCBYyxRVXlCyj6xVHhcG8EnCZgI3Y40pIIMupLj2KKO5jzBz0GKisWgxmJ3
rNa05S2MkV8KK+Awuro5VJJonQbKJOC/6PjWamFddo0bE81w740CslZodqkI
iX0izcNGx+vZWKREAFuKlT1zJTZEpD88cDpJDsy/uc8GEzBGrOhOVqZolkNC
aCCaU1gebfqzeyMspcRwi7XD16Pt+9mX7/QfnJ5j7tqTw0ZpUXLVI4fxAEck
q8reXoLyHIwjI0+gxK49SRo3yK0Gide7QipvrSd2rR6WaAxaastn2Fc/LJgu
kp5ilMm59dl8Kt6ZwYCmyj8k2plkAif5M7wfeCk0t5YRmTmH2nyZ2TUpTOTD
6a6r3lUNxSeZvkCsqs/Q87/tGDeqGbOZ8ajCyl0n09oovQV5Nj1vD1GBWmQm
8klmos7Z/hTTpPx1OfdueE8b9ct26LifjUvmQM9AS10xsFeg2F/sAcy3i/DO
lFKNQ3cht6IalSwkYDTfL40wkWhFYm0Hg3IbCBGj4sEpAYXnS/KaGK/gyTX0
t8arEHGXsZocnamYqE4U77TlrmtXrzY5lQU6HZ50VJTT4SyUa4i1VDSu6DBK
vTcxhglP5nuOTWTvg/BX2jWT/lpW8p5RwzFhf38WmalKRQahqUGa6Vy3OIZs
iVbDKYaatVcm2gixLBycm4E7bBx8ScHVUdjsnZJM6TN62tKivUGI7BlZdLcz
L3KTzA0HQjDjLl1OB+2iOJvi7nDSxV+gvQ4EPl2fghxfY3eCeb0UtaygmB9S
2L0oXDvycbzlEmgSmGEI1A/nb2SWAPagulBFm5S/NZMz9c0oW4esrHj24ZHX
vc7II+t2pryx02gdYzKw58liuvgRqGYkZ3VT6vVCM+Ilww/w/n0zKHkyMoKj
Zj3deNhZcz2ozcAvNgbi8y4xQudcE73xhTRn4kV8vH9Z406+TGvhDWaogcKb
WnpnubOztRTomGgHsJgja8wEYvz37tH5hey8ahf9KadvQToSjYQYMhKi1B//
GgN4+57Fo5e/eX8mMzd9SaVKxZwiP1I+CVPSoTMX36UJ76YJ+VNYfojCyPmx
ex0tyEsXPpb+1AmON2G4Kf7/JXRgzz56eWxcinDiJuh+mIqurbTkl/HxMkrj
cojKThgqRig0DEXybXvTX+lSStvE531TAYbjbGgKDIU2tOL3b6pDp97ZgloO
SWIgb6Rr1WsNLxakR7j0uj+XwyFJHM98wv4xmc5aWvmkaII3yWFIp5Z8bC5e
ttBZDIjwL2+bd23xQsxLMlkM7QAycQcgSw9a1caeCnOvcGPNGTeumM8T0cu8
HXBL1J+2tLP4Y4cXsKZ7Og9hjgFMao9qt4xw9Ztd3YcenkhhLjuoBEnVBOU8
mnRenIMacboqUF05TIUEMfDjLar/ybJoBJ99euex9mr+EicRkmorX2uw7gzS
DisM6agqBg5s6wgpnx0ACWVuH0nJJS56e1PoPq/qU5yMBURax2YPi8wX1oUM
SdMn0TiojmNab9cnQnOLr4kJwJkmYMBDiAamqhDpjLYjCH3LAZkYAvEimbtE
+c248itZ4jumE+jVcxIxQGabFiwg4fmGFInLMUF9KbYRTdYGahOq5uswNV1+
50B0E9p2rYt6gBO8ZmmOtjCRMuPtU/hkYBPnM3bGm/U4lG9G80NooopD1BCU
Z5GF7ItRQhX/emT5oqHwfIJ0kMyINvRaqceaU/93NiTDQQbmLeK5zLHOIIpL
kHWJmK7GmRHDT7rjoee3bqKCvbTxIrHt8xOqIFfJxm4xxXpRNGW/y6fVSGWZ
C8c3cRK6ibhdlGegj1cMAh5DvvYiCuPPZzf9mgiQVUf2LmqSM8H0dwnScOEy
j/Mzv2O/baPTH8x59HA7W1DfH04J7xZVnuZC2+/Rz8HEN/04j88sDD1+oaCX
oh513bEyrVtzK3r5feNE9to9n+yokLWiadhJ4aOmq100OvDvEUfpHRf3eif4
d/nSlLDL53Osf64/623pvX5bZxTfCUhIt9h0z4IBn+aiZGrJL7Au0Np6iwDa
7mCsNH6QBgw9c7+BKepi6YLQFOEkbemVehNocwCrk64+N13H4AlB5cGsrHtk
fzVPPd8FtdKRZZkzsNEsANpw63wjCW7dsLwmLV2mvRF1Cn2YuRh9dI+qCEmM
cH/mzDpiIjk/FIC+4Cm0wIau+i97xwBWNcaLOL+VqUwlHqG84Z64Mvu2OFfQ
GFr8DhVA0JsofNDtAQpxJedQ7eC8es0keJI3//Nf2Zlf1RoSL6/IGn1Faht/
VroGtWefAjdLXTsv5x5MmhhpFqqMZBEVUgCKXklsREpBgICQQoCFWfxCqrX4
8EpIIldqfNfKYICima2xh9trf04SvA5oVB1x5/BNcG91ZidoMHQklcb8simn
QK/bkxyBuT0XporOvaE4AsGNPWEKzxwfHxWdPJTJAzmtOx+YlDsBli31CgdJ
N7/5HNJew/Ca7itJj3JL19GgeyTKM9ZWneb/O9K6hpIc/2kh43eVYxTWhMZX
uxkrpTlTx7gpXetZyYQ6TbKXAX/NpqIfcLE6Z1vXe08jaBV3R2JWchIvp9RO
7p3XRC67lsGmcUQSrwaagpv0XlB6ZBpxzZbS0RXHVXmDX4xEfbzxMJDnGJa4
ZYQTUtYokZKKIVq1EEj2/hsjRGkRJeZhaE8bZOKrSKqWW4wsWfv0impbnJsP
GCuuGg41ElJ2fW5TXVzrMjtv59txOPD+qowyhhr+iv6Szz67NqdG7utFiq3+
Tab6iHJTrcjwQCXoTZFQksj0HNMN24x63DzUKcLGufC8bY/BhpsUjtKJZ4uT
4KaG+oipBPtrWd94kZGIGcnNPuvSQhnbTmeLRqK3ZXai9JnThKOrL6mzumMH
gXOTK2Ueo7KSNnOaanrYpZzV81Pt9ZOqShO7Bev8dnIkxTUWHNJbJ5g1R6X5
OFe9oTjJCOJRhww1YKEes1rU2AOc53j5tb+ZGJtJtl8x8ZqXJdREB+xHNKEX
h1vuW3rbkGaUjtmqFPNg3VZZEVt1zEKgUftHPnzfO9Dv5YyLKlKKa5N3Q1r3
5+3e40MzyIcXbP5xVluQcfoXDLShude1CUesVYYKFlPN45vca5O8RKGrWDMe
8ZvzTfGYS4Cs42qV7kZDer6Z6EfRoeP1OH7WwQDNU/LbJeS7Ubtup9coGexz
kDZmFm4nAF0+CWu9truh2LkobkOJICptuOfImo5SKNDVEn6lfik1/HcIrZCE
pXInsOHjqKUhvmVeYkZIZ1wZKj7t2I1f7w2CpZQWImlth2sj8GIVWF1CF+cg
o68mq95U/hVb0Zl/E1Ltsh3ra8mtUm2VInBuR259Z6xDs0jgsLRMQVsEWfQg
liVgdmxr4WudbDO/0RXA2rZDPHTZX2Ic+g+kh9FsXgPSREvbyYQ0WZLa+wPQ
UdvPn9G1oFfbjSsqIJAjWdhYAnG7ItGw62s/mYmuCpRHhSRk8hYOY+KjbwLH
aclQJsm18lpdFKDN3////K2qmWMJBiglk5/ebqjAvRC79nAg8A1JigNeQTWM
J5yNzTmO3vNuk/f5Tv/DxHlwSLblT9QucwytgsG4RFUEo4JG6v8mu/Hi0oNu
CGiczJ1eUStS3DlM9rs1Oo6NLT9Nmc7O+f6ttILyTEwKveSVBtPAYyiAfE39
LAlXG3+EuirgPtZRdBGb1AayOqo8YUW//j1a3CQJVXSs70mYJ6upeeNdYDRX
/+ZmMAGoW3ZDnP0ODCqQnicObHxjJDGzqPaGZkZTtf6mwgCWBG4HzPCO8msp
IrhWkflRM5uk936fcsmN7o1/oAJocwS2IEluSTQJLa5mg8lvCasFZAJ0HVRB
tJb/eoyhrqHR+AKVk5D5RnHJ25puy/+Ldpgv6kO9kWko8j6s9wzJLaqUrOwb
DCHKLx5fApU1IwoTNHFSYrqG2CKp28foX2krpaBk917xpYMRaY+YE1iVmmRk
EK6DFDGb2c7ONOowZGG9EYIcSt3rMI7CXWjbSgdCaCeplbiqRI3NIvJ83kat
Sjuk6xngDXB/XuQCRwKoCgyadIKtfJWYPKFnTW7t9xjdXpwQo4I5I2+vbslp
sUZg57/G0XukxmOHuabLTVwD1Bi6sJL+HKhd1UfVCPCWV5SgXB6daUGs0GZa
taXVdSbPOdv/YeJ+lx8H8dE4rvTPGQhtyAoJiCkgH+0QjFKNHAw/wjrXN+XT
7GOHVxrqnTKD+LxJmJQXaNnmrMMAtUnFT1Ew9OX5bzOh6l5F4pwK/3nzqJjF
gKMMpw6TNGYNni2W/m3wICir10ejykj/Cq5H0roAVkoB6T8ktDU6B9Y9GtBm
ixzn3pXMTFieypQhZEBN5CXYWAtMWYPYGaN0CI8P1XnQR4JnNTfB9ps1xWTo
Azbmv7XcZ4kvvPApz6QKY49DOmFaI0Efxu2IgqducCi8bGr/sQarD7LNOs9V
ILjenmgfP+85v0BSNEy5CWyKqSNZLEd5Mz7E1PtJOyCJvZ5zQ+ZrH7bFI5Lb
E6Cj+cdHunDRqsUWY9YPglcgRjHFPh5GyFv+ZeVaCUjgMID74IvpOgoxs2dz
WoaxJ4JUbq8BSa3bnGAHlJL3z1xb82DHAG0QdwfZIh2M9pMr7edC3AGjCych
FWMOJEBhR5wVmZW8prPc/zMmEI2y1qYIEfudbcDi0TbfHrtchL4lZUcKX3nj
EYcqVyywdaDFll8DblNmxWpJJAlnh0IL+hSBSKgTvdJzDT5/7BRReQetdWP7
PD2u6QkqkxbQAT4HpoknlpdkUMR0D9jTJWD+8GWeCxOJ6x62gt14tfUw0cd6
9stGPemlaxeY58BMRCqxDac+nafL07/6NSOfLwXVX2rA/AjqUabImG4RxVed
O54rqu/k7osgEd9JSllyRK5BE/7+XR+ye7pUVy5JXB3QpEX2TRaEBt2pPq/Z
MoqNvCwowSxv95iYEL3MR5YGWKThlLVcoxxIaRAP5qxz0unu1alLmmgS1510
SsaFpWZV701ldtKWLFq+x/hFA4qlSxNI4Zc68qvft4OnzfLX2VJRVp/nZtFQ
68n6ocvcZBiwvb7AWE7ryevpeLd8kovM9XQ9mQFuV65IkZ3Q7cZq/GJVGy4g
++6Qu0UnyM7ckUBEHyW3QVJok5y/5FV7zQtrLFqoHNvbsyFmCPwqCsdZsHGS
/FayrCTlG5bzyUJ/hS1B8M4MrHFGJFBjrugEvWnyBhtqsKkvgihr28tNJoBx
9apwAC+zBG+tESGJ4jnsSWWDYj20rtMXgeEjQNw8O0KCkkInT9ZzFg60bRXD
8oZbGjS7BZj/u+l8GT6m00fcWdy9yUqa7inZTJDmQH2rexp6gJeyYq8KmDbU
iQo/FCD+KHTSEcxAvQHXczHSoeMYcUDAJ2zq8/XfFG+1EJiFrmaI9/OJ4l2c
JlT0Zl3IJILmPw0rpadFAQqYusB0rJ7+UoCRR0bCmCKWRnrhLEdxe933moHY
DrykxW71LGpsp7YsrhkYbnfiYAYqIIgi1DFMq4KzNlIed9gVWRdGNGekY0Ru
KQO6b5hWbEi48b8Dpdal155ywaJIsoeeWFwzzr8krgTdSuVuEZMgb1AZggaw
8SV9YO6p9ITcr2vGYYjeCGNujD3oGKNrXa/Hnw2px36PcwRHeolKGg8ukRIA
UpPebnG1XQ9Be2UpjhyoE0X8gZc2WTJdBXX4lFy4qiwGW8HZ3+rWi5t9Qk0N
+lBqIDSZOTXPvKIBorQuS1gwbMHoMhJC/EGadwBt7oQGIFayaCtgKAdttn7O
+9q6QGq/BVfIId2EpsKGRlAwgNPiQfzm0wmE0YmPPdSu/CpER9qO5If1Dc/C
0imEWezQu4oYWXzTVAOPyZ0J3THdPEH7wj8PjGhWAotOxzpWUA1CDCROz2sY
r5vHkP8Lr3ljGCHV663GiYFGSRKJE05/XA50/4A4HNXpVZKJLu4RT433H2sf
98x5LJTIuaFqEAuuqPj0ZzkWqPUjfXh57fWYPuNrXCShaWcsgjwO684jTExL
/FEExd2SAtpJVR/2B/5gI4ApqTdmMlQQiwFvirhkWyijg5vq/EgT2tyKrT8f
9u7PtwONnqrzl9qa5B0m20IIHTzhDpv9de1gQJWZAO3co03JJQDKUS9nv54C
y1A4FWaojz8MEJf9534wRM2boytovpXdC8Kv/KJEZKrhq0DXQrLJXmQHUo9n
WHEEl2Jj8T9Vl1569aIh2B8lT5qomkltnOwj6fOHrP3JTcwaBo49d06hdm5b
crbdEfTbtv9wdk1b4DVe1u88EHKaA2zMUOiW+cVPHCS16bBsI6XSrotAiUWW
BObpW59IddwOtWAXODO1rEZwuKpsI6IWlothVomdMMWuaqZw+wmpn1FfPOJM
E891Ykfqijtjw6itglFlkrSGFGaXXbi4Qx1uO22rBn58sc62hzenZKyFonDH
uf7EUdDfZh1kuddqnb2zZM3pGXCCASuV2D5usMPfxi7vnYR3VzxP76OyS+Rp
6ZWKwI6Yywkq8dQGsOmQE+yU+tm5ZHg3OxwjZDIJiYhch2IVYPeDwRcw9BqS
qB06fzY+7Q/ak3OBeiC3HoZIKx10Wwx1iOIvZyAXs4h1SyrXkRoLdJzbR4ML
nf3DXAwQF4gFNaPtRPowvjJBUKbDXj/fCbzPbYvmV4d6opTg1lXNbmSnBNxA
AE6fmhe4aCw0sl8lKrViSnRXcyI8MUxBG13c5IxnyeOtJQEW7i1ILSwBy+B7
LSp68efCbi9II0jIdUZcOv4e1nxsUQMr+6AYyyS6Q4XesRsY7i2YgHaH1gPp
XQKxRmJOCnSaXQ2ZYrsvw/X/2wIibKWSDEQifzC1bDlby1ry0o0vCZN/MGIC
8th9GmYokmYccRe1bCh27LUo8C51xMopmcnT3urX9QHwrGpcHSddJh/0eXaW
sOTC1bhRNqbcamViI7tb8DpN2IX0WPhQyeSjO+W/DiNIXYAvwGIvRfaLUX0v
m4AON27ma0wOTUxU3dgjh0u4og3Xajf0RbLgZBeBuOyeOFuHPwAfzSY/XyEX
gm+pTl06awJDDVsdM++/+NtDKKnmrl+XyXWVSGghk4PUb64VCPGcxAjff3aI
cuZKqOPfaSYV6Fff+O9wuNxRwXWKaMCnT7IRUnBd7QF7QG3XrC7ljrd83dNq
x75GWulOUrB4+1m/67Jba/TL1g3/Em1pYVWwV5u607Ki5ELS/7MmkpvsgMwY
oMRL5Rka4NdMmUZ/fDI59N30hd28Yx8zmmICYFh5rDRkjaC0E8jOHJCK5T0y
7JhXFGKudZlGIttSkERYIjtFV3jeL5/JSMOP6HTbeYQFkwClvLlSEauPYjLV
8+gsSErTR1mfWR3f1kmr2fWHbjOKD/AOBFjM3ayTSlwsyYUErH4EN5Dl2NiE
xYxXzpls9JBcoc6Jj2SqrNjodaJ3M4s7IaW6/sLDGo1J2XoEUKIhSsBjMqvi
b2vK7dFQCc0Bkq7BVuDGZ/8Tt/MHK5w/pEIwh5XbrUonGxcKB3GwBMkENc1g
zwCC3ksDWK3yosbF+KeMeHgZpOBaBHnivgF+E8GACAfETiDH2OA0HR1JhlJj
zDZmtN5uE2mxAMZhDGXfyUZf2Yz3j8QdHxzBN0CZBISqOXzJAKtwLpGL2htn
RWkIMKuOTYHad7wcbPKMusYUSIyoR6qZTMvGPY75fklEGNW5QDzU1YjkeEE3
nXT7uCilCiAnq+pGv1m2XecdecnoPphkzs88exzqqB172wjTM3NN5VdFrMAR
5guhDislS8PM7aIdTsteF6OJbGs4uDjaZyNH7J9uQut7M9QTFf3087KmeXnE
3Hs5U0+rwZSDi0GlfecCWwFJegestNkqboKKXsBmoqNdXuOuMAd/cbOzghrb
jSIcDiT+TiTQx0Y7wGUXteRHyMpwdZpXTBWoGjm4bWpCzIlhdSWk+W4raLy6
H4q12E800l4zKLf0aJGPnSdSsmsyYJ+bX2hG/gmGN1h+HXrDlIvVaii5K+l0
14LP/IOl9vcAo3aeQndVYzAGyr6pWebQCli+bDlz0kVk6PdMGQ9OSBJgrwPR
6ZST0UrynE7a/7ga0528qmqy3+Mmkw4pcfaApMjEZM63mzIbpB+R4Cz4GbGW
AMx41Z5/4jsE23wpu3dRn0fF/5hpwaOKo3m5jVjmxQeRpIdxA5QBexerLckd
Atnb9OtAjDeWOaqlxEuTDYw8sqf2CpaXAqun8vY8bLuZmCy6MaiP3kbsE0Ip
w53JGpB5+gN6b4UIN3gkNwh3fAsrL0cJNxCif2iSTsx9xuzB5U0yUuZSyefs
a56glwmIY5vUaLOnsrXNIuarLZBTx5H7VEYPTSkUvG5NHLGH7JEB2+I6Zts5
KmdGqfcuLEZYW4NTpU/Xi6oSs2EBu3gDGNIqnM8s9InpPhTATp0c0l06upKc
3/aB4j5AN2QJ98w9TyPoZIVGstTR5AgGU8M1RWvC3A7H0VydpnuTGgXrDXhI
LkQl10M8REpq2MyfHjbZGtpeTB8JkmeL71W95jgzyIzcYOQdAv/ee/zWMpOt
h3mWN/8nzApVe1mP14YLMzNHJHc1pDc5qgCYLwwiWHB4hBMv/Fa+lz31YrHg
kl/EGGVHsRLwzanpGmLgkJ1iDCKNZKsaWgFmgZxQZBm1TG9cugsaPJ3/P/Nm
t2QXD7BVd2qbwjFV1/7ZOEmw52jA5dUOf0JrqEbfp63ocZaVZUVO1jrWMP4h
6+17IcZacFEBS6jGwEtpR+TK/wJLI+rBJnz+QIncZc6Rk/wpOL6+nzPkVYl+
3Wd9rlLLZjUUCgOx2COo5fRxk8MiB5Zr9q3D0UTlOKkmfxvjkLw4vSQg8CLD
/AwDU+Ott/6dKocHVd6cXWz29NFX/5fsUAsttyTXIXNduRmf04uHajHUjTxg
8ONlhgEvAYn9vpJ1ckNfNy5qu5dWrLajEg1Er4rJFzUdA7P0+jZpO7n+8GjS
feO82Y1PsTg5zS70BW7mwaDkq0mJTuD1kaT0R266iS2ymbfDYkM6Gj8VKnA4
V92LpKi39OIQfRS/+Dkaa7UDlwOubaNUorE1N9pcLNgefdRhKkB5ckqtC0RS
mpTBWOAY0ZGlZFsDmG93MVDQHNbplNYhWMRQ4L9raQV4wHBO3A9oplGA/aJ8
W816BGqHgfagrkXnWj1W9ndACH8z1cigZ/DUhjekax3XcjOu0H6LQiB2NO9l
XbpNbYjWptZK08uuj3DrQXzUnCqEQm86njOkfkZmT12FtQ6faaSVJ/tgXXEh
6Q9Ehc1ZuHSwboewaiBn+K6dz4ClPhFxUqCWogqxbFFxDf5lojZGhyW3H8Ro
puXtw+0B3Y1ZzH3l0/fAkzln4z63IqeYgY2LaKGRj9Ew6TkT83R1ObXVwjmr
m7XVVsOb4Cqy+tG239GtqupRaZlJWKMce4xphXwc3tYmnv9LcSE8rLRdXWML
FihJLf1FxMXHwi9czay0dwy50aiidLbBf/lgURN/Cch2SJnHV5s/ra5koQjO
BuNIVAz5eQE1HLE8UBapaTk0HJBSVZLSudidWDO5WDeOIUnXNkqoWUDufoTq
+zmrwaQZvlQ7vgNojf2Kx6CcTIZG1RCpFOks60C/PqeFVCzNIS7Oj43Ot8Pv
hZCwH/uV74xDN3+FO9nAhpmJzKqov/UHF/oY4EttThgsfukXf9COCRFBQzHE
+OFYev2U2CttndZYpgGMJrt2zy2qTotoMvSXgU5CYd0NFDm70C4X15GJxOn8
mCSxVed7jB5xm8hI7bDQT5Ji4uM5um99jZTmOUpLtAZcDittn2d0+CUBVkEd
o79rA9bNYjJoMpKGfVrhK97BnOwk0diDgOilKm17rrMbFZ0aA4CRSpc6W6zS
5tRIX+ESLcRPcfkf3jgKWuCEfWh0tS/gmv4bbWCsKGOikYM19NlzsdTFp15Y
Ty5GcPNpi7QXmhNBDvtLOo47ET93YN9gN4hwluhnyZy8btPEaKPICq408KMp
g9FatVukn+IQEEUICcSkuPPZzO8mYjLD7zF06b/DaFlPekPf5cS1KGWrvWCH
2DsJ4ag8733J6hSsCBtkfX9113IvZLyaBBDy148N2VEO6AJ07e6+Jq9R5Rk+
xJtJF/B6SYey1onuGPCH9mrzymM+j5LcAXJ9x0lwteZGuKRHjVpUu8ZKV8Qx
WJSVA4Dfa/yCQR1kEF6Lt0sAw0O8Z66hi6zk5jI+cUUDrWu7RDjA8U4HuJow
n69NkYZPtN/7przKj715fc1Bwae9th3+WrW5E5phORiNbJ/Lgxe8TOhfJlY2
ZqsW/6gyB1iT1A4E4nL4M6o9TofnU9DyFo5+UgQ4ETw0ymHrzEB8sM1b2upH
PncsPuzocLKBxG9ydo+r8XrUnuyw5idz/xPgxMsNsn7CGj7kV4XcdiGodeLo
Qnq3cUcgf8bk5f/X9aIa0Zw9FcuGn+AOJup4EwoEWJ+5ovdj61FcJn/UTtdr
ohD/2enbXZB0KeUtzEFpyh49bqgqWHexDjJBj48UWV8QfNtNF+9u2EMoUWbX
qNwFFHqQdh57XZFc/sok2OIJcW3Na0Y91NsDyzf+uOVMPv0BHPdmG43Teu+g
oZxLsib9i3XD/72g/WPgQRy02Jc0pJQcD7LO16eOBGJdyLzkEI/ZfnksNQl8
nh2w43Tk5zI5KcAc+3IdPNtyteRQLH5ebEXxMPgKI8r/tm0u3JsjZL0muYGu
CPdQvSZ8sQg8H44mIQ8DQChLXiDYtd1/b1PEoJIhSnczHKwHJVjgRzItJdN5
aD9wUmocklM01LZvpLElf4j5132bajaIxDcjli1UgV/6pVS87D7NuRqZ19/h
dJnYZFBNNsNrDncNADVneCEN2LxXhocM8HhJoSUJGJiUqHV3NCQtAz7IxGDc
PT+S2hWgq0CkusPadPrcA/B0zAGw/4uzRbQRgcovrrF9S/C975QalcNcgXZ9
blGlepd97eFGViBM3vZfVrbeM9fH4WGJ6W3kve/e+Wkql2dgJTQGiTkPRS//
u4/a2UVGPyUE0Iffy0pPnxzvqMc4t/pLVeVQ7kBlYmAstu5L5WRccLDDzmWk
wEGgymKZqx74GqmMDina7slvQ1A2kkkzz7hNOReDoSKxi9R3onHwE2FO8gJy
EOAfjS84HU98q1sD6zDzxqp6Vg6x9TvnKfTkTLU/AmygSVjMTINnARqYegZR
7eBQ8h0UtfKa+hy/vGbJTzbDVZ5jwzJZKlC4jC5dZHYBxxs0sSlwjaeu7U3q
JO4AUJJHxkVsxqVHvVp1LUyk7UC/C3Yo42KO2awfnQqEdoQjhufUNBOCgZua
kaN3hYReBlYKGVA6BsL0yPgK9gAf4iI07A2gvWp8O0ckn/8F7v7n5aDV23bT
Vo7iyB1VAWaWsQLHyBeI8zmESFVg862K5TiROlPBGLkWBgLANRL3esZOs0FZ
XY30vAsIWm7/aXKJU7DzqNUx72BeyDH9WKBbq+wresvM+Gnp/b4fTyYZ7T0U
OpwFwQbuFpMtklMJgqLeEhy30MYfhYBQnaQt+tQ4HKmXAvQ/yO0X4x3x47sA
1w/UaEgzqt799WxYHEvIFiMqzlDzfQ7ohumsoWskS+OogA6KQGAAIAmxUJZO
a1S4ZvSwgYfKOBHYDX9fj4hF8/MrFsbWDnIP+pj9IC5RWV/J+fZWJIEPGWKx
qSkBBJ0S0sQGMzff1Cv38YYWqzvy7DgZXJUFUfYliVlwrp178Oz8eB5uvkJL
5A2bJOK5exdXe2FcxCByG1VeX6aBW7qfjSsKNb58hHpo1fyBvWHUkUuKeZKp
8qVXebf40PlMTjZb69YrMq++TDFtJBRPgEkgRGkZwqtrLdm0atg0+fHNW1BN
yEzTIg8M9fqc/iBgu1brkbs4xVNJd3KANxnGJGfOUeTObNm9QAyz8vtm+E/t
RRKNo45/279oOEb1tkFzXr/noVdnAmyklaFnhIDW78UVaqNDM7A7Z1GthYsp
jv/QEDzrzzKN3t1TfDU6Z4R49/wsnGXEmBvvJsNeGKWyl3QvIZgd/or3pYtQ
aJOT+YeC0f6s+XtEf9/bG3ZGCt38wFFkkhZRZV0a9UXp9TA2NUzuvLyz3Nue
KvOH9eT8Tg1fY8lSfryA4uetUNhwgYM6W4Q1LGw+0HSYxHaV9uzydSmwyJoR
N/gBd0f3isPbxXcB7ORiTIzBCJUB20PAk6WkuxD6DqmEPXSO2nQ0XXBEnZw3
vSTaZ2jyr7krYzsY/2QOtSEiyBbpBqpjDclDI59yhRcAxBcYaaUY8i180Fnn
mzPHSp65mLWq7tv/ULkm6YMx1xyktz2kOSCVfpy13Fp3zDM6OKgsczBHJr+j
/REsstzfGdJfJWmA3pHq7/Qh5srvTMwUPorU2adHkKdnrb9dTiteC5t02NW5
fCElxrqgp39KzzNIdRDpyUrSopwWk4APDfIct5EJLVkTgquNaNR5AFlAyuLG
00DfDNzKV9vw3hwI6SIlDo9NVWFORCsTZH3ZPcfuykaC96zrvDx8x16gS87/
Q2p9VLqxxU2xZJ/JxODzCbUnNWol4nO8lJT1Zb+o6Smc4DVWDDtlbREykCqY
e+1Y2OnwOAqVccbJBA7YxtApQomM9mtAbNivwziQvaRx9iwbVGN1GBfeKxRJ
8Mxpth2TDHFL4ZEKVa/FTziwIy4s3Qr+Q/sxwD/RoK58PwHzMYjWA+LNVxXw
ci/+nK8qsMLzcB2oRAgGvAeBI4gpQYf0FCapPWmASGmq9TT9gb6Jjh8/ZRHQ
hq73NjQ+OXMmgw1P/h/gkSMxjuurwM334AKOPXOX16e8zaD/aa1a0zM79tY2
O5rNeTj2CJRs9wWQikIpKJ0Tra9NMPv0uJBkDqW51V/aUmWBvff1Y9YzB5+K
Sm7oConu5EK+vUl5PRmVGyHI9PpWA/9jrnkaqC9XEpB5OwfHcYqQarGP/0IY
74nDQO1ICakadJDB5ASl1KUEu8ve+xHMEjiAJYwhf2FPRa6n6n7XPy9RceN8
/1cJq+Wnmua/4hQ1NtihsI0BypPskCly7w2Ke/tKqUnM10PG0WSluMFIuCml
UwL1gPakuMjEvxlWcU0bhM93AwzxSayIeX6smeYNPJtJsH4ay9edi8OcDNaV
pJaMCF9Ez3pmKkDGPKER7mpDIMrerdoLbCwS9In32qwtneuBtWZyLgNRhqHn
TPvORLa0UhoOjpPxIKQAIaq38uVZWtoAFCo4qmgFi+ATbBHS/kVmRO4tBION
v1V5kXXewSZb8lxcCzR7S6w6Yq57U7lnjMeWfic1oOV+oimTGcnMoyOeeG83
nJ9woRuquTrddEa74dEOPCqArp7bcTr2/ABE3iy9TeQGUWhddgpjsapsk0Um
MfuyfSsy50oQQgDzyvAQ+nPWA1d3NbXmnt/BHVwZWPnsBEIE+oq3mizlR6ky
sRqy7Srz8L71ME6TCNJpW9WUWzm+02nhCP5GocOubzxLhgEl1wEhE6Nvkdbb
6DxJBKJslYOZQM5FD3U7Qa/Gv1denu4C9JZVeiDNfr6C0Q3FnoxQKElWucCK
NxZ7D2xKJD9YLCH+oWUjj2NPjvRDsP4wkwwUC2KjG+pmG5GaLxuVi77wPLhB
fLAg9So5GHt479oYO7v+Q7bYDKKtaw1Zrclb7FjkFF+tOWadi/wZ6JXgbrgE
WDRU4scmuR7lnlYC24MPdpX+hi62/RJ1kd4oB6bkC8dSbp+J+nZNiid+UPFX
mVkEwp/oo3YLnLEV2LiaVcI+M7TdA26zop89J/ia1hosf7ouoRVUeTfzTTY2
tfPjJlPVZnw4GKmC+2E96wDP/l/NlGeSlTVO+clBqfRJ3rvmjpLan8FJLHzs
8zKAYak6wlB7mRLFKzM9aqB8zCy2PXNLajCU0DQm4dw+PzdHLY3mXmv0HXQx
zhcVOfS/4ij8gOQiJpUJAYDM0lWqNatiQuuBJngO/K6Lr7MntlvJy3OHWtID
LPWrdNMInKIbCn9P4cupTI8y3IisdjkI2OiG58mpvUa9wgQqNzP/Jp8Vun7O
VmEvlD3/FzcsmvUGXOZda4H3+Hc6Mnmrj3J6K+NvNm9LSOOLtR/nFIePoFLR
aOF+DllkMY84+c9y6jv5ff1x4qFfhbKbv0XmJqLZNRKplqQNaj2p9ug/gx7B
se8ohT9aM4WJNI0Iy6bL5z2xN12OqpNPJjcq2cuHaN2mU27mCX806OxYLkWG
T7/vD73niC1p3ALlocqddQ03Kknxce1mjqi37dV3Qpe+Rno7vubLrBiMpM9b
i3KrvqmgtRo8IRifmS+6lnp7IbeN54e8/FqXcEkIhvn2vp/3XtjW4qxjIGaT
/tdF5to1ghBaDE4O5PExsx2ZBoQN4WRqHQQ585grLKqZSFn2YIkoi1riK2Q4
qRfxhn+BtLIi78qPdyQnAPf9mOBaXtTYpwnukw8yDEIAzzEHnGpm6pPCEbc4
9xTHNsHh6Iffj9UIblZ7K6DJ99CMd0onmG3LzyaIg25/KRe3bzUEU6y9RyIc
cxTyPYYEuK6m8OIhKlO7E6+zelm6FcgUk6tvV8n64I4q2gRdpaCHz+r2jLZr
7rOidfqgHYCs5j4zPkaAf6pmKcPsK7l84L/tLit+vJFKaearAEf7t8J6z8Hg
LGgJ9r4TjOEs1JwiDC7WjyKELP7d+Ag/Ut3Xgg9aOKm4l8a1wfPGqxBTG9nF
aWCqJ6LXWsCEAVUB7aOXy5cYBp7FuhLouVu/cELXO6RmFJAH/fc5g7TxpVgw
u1ftxrVLvMEnATgdgof+DjaX8nd/e5EzvPU83e9l95DxZqmWxV+WUMK/BEOE
BniYE9zmMXqTQdfuZOcSHRkHRwT5BTjpWALSiMAeW6X0LEwhF3H70o09FPcc
89mIWoJ/6bmJJo9LHvC/eAxaZzzMKi2V0BqXbz0ex6/aSKlsM+B56njSb6am
FD5Y6au0ty85XFheI8eFPFbvWmvIp/7bc1grdgP+k6vYf1ydZ4n4BfaAaPpf
sc6aQaajIHEFxN6Uykn/1136xRiYqrOUrvwFtHgAlFuvb+soTMj3C+qZlp4f
jhKtCLRXHFbQvdSdMZO2QzvaV0zryECfobjP1woPwpu+F7o6TGoNYASkeg6M
IFOaytCnh3LWM8FY8RM4mNADbAj7PpvTjqLYHG3kWTcVdN7KYdlGpX8p2k25
0Bmf0SXKILpD3WI/znFCw+Kdr/WvdEwnRvJVy0nxPu1NylyM6LwvBjb1n24+
yRa3kd2aEDClBF7P+RGE69YV7Y/ZFYir0N08QQRtX651/AI/okV6eNqABC6u
jU+Lgo/A7gOGkN1y1YygO0A7t9nFMWVBJa25PqXr2al4qOu1OKflT06YOJPV
CWWhyUeXceERzr8JXHvs6IZBRmFQfqXbd9xEROeCFneRzDNJdXKp1pIXzMiP
n/LXQzW/6I7R8gx8WHRS24vUmd0xXeTNwwxghgr/Y0ZP4hu07/Yj++994xYp
gRuVMO0ihQuew4t0yHMbUePuIIXBLk+g9ZPemtM9ppAKvTw3bDMxjtSlixdp
Upx9aonMelNy+6K9cdH+mnuHi9jRPblCjF+ha8+BhLe4AUxt6pCmS1mYVx+V
ge7vWPJy59gEi20ECWA7xYZegPm4KJoRE5B3amEmMfHGDbbVwpnspeBIrZdk
WMsfy+IGn686D9oP0dAefM+N+6Z3ehp6e1B8VJlYZIdsAHJ3hzpdheZXOUE3
mR5+sj5CJIDEhSwBdjuxP4if9tEhyKncJnr5oBqkncQ8CO1LmpagZnG/S8eU
aDU99OQ2LhYQ7ksOYMT526O+lZv9OrgsEUvdx7viRPCdrTxt3t2Y5IOAfY0m
fOwl+toJ5cAQrTCll6qgj13qwlSlvRyTfGXTAzhqN9YowBZLAMIU++Y9NaI5
/tVRPkc5DJMBWy7E4VR4hHiRwEb4rchelNb5rZ5TW7U+NVheiQnqRu15klpz
uUG2zGhI+SCMI5HCu/VXJFDa74DGF2Q4d5lXqeNCHAIXRqmITmKr0PFCThAX
GMynpMMhCdDH9+bo772EGuCHXrXhuHxuVhETtPEOTlHqT9+3rHHCLvVGykpC
trJ17BbgCq06lDc8aemuqr0YHfWs2bDu5bxKrfUpA8fk5I214zigNdCMll90
1uOHoJShZsEmJQEig0ek4t/w4pqQAZpWQj54I22NJpaboe3KPgmJRrmyLyQx
x2+QYC0P0OISv3Bwnk6qPeDd9jCDTAKMmnTxKtAVUf4U+sRNb/ja2hzLerO+
iKtHJR4K+Ezud3qE+2tkwgcszMiey86NAQyioM2CxU+dinvaC3bdFpAt/2Pw
kpixp3lTVUFAqLqGOz4mgAL/xVUsa28sjibbDgAqOH60lKbr4kL05gBbUce2
bhREJIT9sRAAmqwOiUL4KxCcEALg1xsM4kkalerQrxO3d2NEPqXtk/PhrV/B
ZIQeK2AcjAUDV8JpY85sY+IMqqRjJeKEHEQ0t0VoIjKqFPIcmh9Bh/b4R1S8
Co7/RKytswZTHlE9FjFBvRWZ+faKuLr/omcQUkU8XrkwWXjQo/AFpN8vslTS
Da7KP8QFroJmJx9esgYPVW701esft8Hxll/sTbL8gbe2/Eyf3Whgp5Y7ZO7r
fuamsF7uP/kUPAx0rKNoY6tr2Rfk+hoCIUJXh+7jw5J4SGYhVGS+VdGsH66+
FsQokoktx/86LHYqh4NEVDHFMBhmvMK56ZoiP2QZtGVUPu9DgwYVLuNg31Q5
xiBbTzcFcyeldPAHu0MMSq1xQbGvW/1xEvhFC7zOyCClFVHy8iA6+n2PrtOt
m8oOY2T+q1SPHkmAsX98lwk9AqMMMWxA2JImdRpYfHe+DKKs7/emtBAS4TjX
B9uMlB9IXonew42HjnIA6itK/F0RIumrNDxyBSdOacpP9jkDJvzmCPGsBFmI
nYAlplr5h8ukeZXP9n0YOQ7u4vXLE6L9zR2JUDm5Dso+q+88JqcptP113GSx
UkGMZCfKW2AbAV1M25Hsby9Zt7lVYeDLantKENZSmLE0xpSzIQ11VB5jZRNJ
aVjlwktf9mOeyOTqNSLkb3pjRv6n3UVymgnTimOF3qUVN7v6u0od/S/D9iwi
aVEO3e9UGxMnYA554icltw1J4BbR4jbXujhU4pAEeHnXPha2zI8yVdfyS9Ki
IcpeCuhR2D0NhrBNA/pGjhTtjK+5E002wjHd5vDBZ4X8uvOm8QfgheDrb4/9
iyGFf5/TVq0ubblHLWjvwM96I1D9yvsVOnkCC/QUHsMVVlPACuQ7cd9wfMIA
u+zd9vpm35jmf+FBfemhuEQCykcbwIjMu/gXjf6vdl+QpqANm+ca3adHExmo
3utCi6CliVJlonQV/IrqyDlJneUwqZlZ2J8ct3jMEsQR1BGDIO8twG5lMq8T
lWDSk7/9XO27rLWpakaAywVWjNNDJ0LRC1BSimhue1AcDjFSqt0lotL70VwH
gpGYGAMLxLnmkA0mpWzSjNNmh08c4cjjO2pXB9GnqHB9Hr7brxs3Y+dqVRTw
mhpJQ2dLNQJ9SdthAh3Yj1sdjK6ai5TKbFO7Uqy5CKZ7SZlRnIVPWbk12+nn
ly7GJ/i8V/+DtkkO0lLha5pAmojkp/T+SLtNU9hl5KntUMQDQpgwKz9EKAiB
wNjzSG4QxUxYgUwIRzbDXOgnyVdWqor55/6lJAGqtQIYXz2pkmmRytFAOOC1
awlDmw1yW0jfzX8vYAX0zeqDRGs6MUXpJ3za4FI3nm3L/y1urwQZoM3w5N83
zyDPtjgt/WMJ5zpvAGa00c6oqdXQ5U9a3YZLfPFCvo6P+4zPwKc1qU85mVsN
xd2nNnhVP3w+njdYLLfFvCfAzXxPfbu7/+VySV4xQoLl+whi6oSbyiO50dTU
BLhvy6fidJjtsRJ9P9DSPpM9YvK8aLcndHKMX0jF0XQMI8+T73vDJilVAwTm
UD1CdGhzsGxtIJ/JmCaJz6AKmSFsv45HiYK0UaFknAI1L+cMJNeOB9BiKQWE
4S5lq8wGmbBa2NMlha1HHw+6dX4PXKHy42yZ/DK4hR+5WUlh8eEAJng9awIg
UI7arFrDw5dynfOQ/nT+xk4JkJHMexfntmQYbS91cj6jafx0IuTfG3pVFBzu
lXCp3KQS0QPbfP8FWlihIrL0U23YrSoB/IcP/DKgaH5aLDhdXT0qBJO16B19
isDFRyTZAHdjBOKCGDtzf15ihGxh0SlFfQLsEwTApykxH2AXe93IUlPKQo21
E/l1up4fjhfxa+VK9zm44ehsCCbseZ6D63mRJuErTMJimFAMhnCc8ZFpp1Vn
nA9VEKAWqLiU7v/6HzMCh/crzkbW45O6okSdRQyg+Wn6K+LUFIgkmUbLp8gP
kmezvrrRWMnd/trAxHARmcZQCTc4nvLfusVNiutsZChltz+OW9ipvMnhE2g3
BWWszN1dLHCQFijs9tP/DgKqA3RFbK4G3BMSO4RZVfV9u08LL18d4k8eAi10
UJwA4rFDZEGVr6bqzDz0rco/fca2TzpO3X/dH9+Hq9IF4heJyaORN2JLdOJy
W0flTLmsjlLOvYAPEIJfcl06kJrxxWWl7HwyP1pfiemTqlcgkBUS2KjIf/Ew
56QbDjWiBMWneIEWRstShtaePYshTaEQrscW2K6HcGNiU/QAo38eMCu5a5kX
RqK/QOW+nN9GG+3lZmHiFtlxG1PFFRPpI1aPXSMdHGn7LmDhZ7ajjmj38frK
fzr+z0Lgu1gDNpXdex2zwECaiWOzMUvjPkXrE1qLp4DPLm7HJFjukrC034JS
18yuKFSr7jnurS78w0Rsrc9viB1wgRKTMnpyDuJ8WGgQn1c3KPneK/N3C/nf
mb03nHG6aJWEw4h0goANARJe6ZZ2UHKzMfnBFlCICzC2pqnybDYcVKKpKUuB
k8Eb1YIaw4mg4IceonDzspsX7mgU9hJfeXRjxZxWuL8GK+dnsoD2tnBymYWi
ETptmWB2kVR6tTzupVIEQ1m9dqtdDXjvB+vnOJALlRe+lP+W20ACk52cX+ri
3xf8cMABcRbwTcmh60RuRc+W6bzQKHSvArigHOTdopDYTi2BwqMHoLM8UuA7
TAvrb/xbxTYud1SkMHBTqvIPOB7sS72yH5bTlFJgj8DgnPuFLgaEdl9sKb6I
C0JSZ+Gb1Klgp4yaRFBgFwjRVd8g6mYBACfpfVjkXtoHJBHlOo8Wo+2Cowye
CoiUJakDNyKgPTKVtvS1Lo8VTSoGdpI2JIShuwzTiZjvx/YGzs/wYqnCex1p
H/Y1YXg2v9MguIUe2SPS4f+4bRa0HBtA/5meTV93ETR8zHlL3QlEBk/fhtaX
m9dvDDG+rZB69gwv4JvlF4OWwIc0wKgr+h3dHlSXsmIDqvFUJMjpb2dIEDd6
GyvW7KVQCH2qhvQnme8MOohJi2TQ+mvRs9JGLQBEiCjB2mjppquFtBRz+NtQ
/rRr/zQqqTFDawFJPDJnPgcIFoXy/A9JcgVxYoTR9zqjQ9kJTdpTHJMLllDS
GhGtmEGuoszdoVIshHO7cunt4LYmlwLC7xAZZLwE661NivZ6lwOQnvBPWpHb
mX+V5ootobrXcEs3PbagcyPlyXCi5GwwYRY8Si4p1ywfqoSILdOawOzQLihK
o+lUApMYSXZvylbG9VOe1GLMtnOz5nAC9UioPeorXwFYVWc9RFlJsxzkiqeW
/mnPkUgxb3lO7sBDFnXqRTAMHyJyBIvafnFbv3+5Zblxm2+bUHq1QdidFTWy
QUP+u2TIxioN4AJC870nooN2Ful6zTfB4QMmO1XpCnJCYk85ogyfhdwsy1v6
3sr3ysgnDUx0bVEm0jnKn1cf4/zpSqdKmSjHWp3iirggKEUBUHgYTTOK48y5
YLXmin+dhdtkGXtwQyyTFc/WagT/0yubhEj6Sd6ijeILANVJ9p3jP2UN5kUS
LOmBVjEw+4cx/6UdnoqkqVfjPYa0eQYr5LXjP7z0mqqVhdjURGT4IGOQ29dg
NI1A5Q8wUsgjO/kaTZE4BoDfvhkZ6Uuoln7SIPCgeBLuQgysWr487dd8u5ZX
1Ycw8yt5tOCg24fJI+0JQm3nZIOYfKk2jCs4+Sn5BmoeRX3BV2vOyHWogdu5
F15/5xDXY+eDHc8vHZKq1+jcqNO80tyHxt70ltjrX/FgnAns02LCykbjHjCt
yUtSwenRH4a716tz4Eks+aj1D3/qOR6IoK/9MsfQTD1MREJL+lVXc/COmYGc
VHXOf4v1ZDvdK2PAEeKWw6CgLipzTmEdkcSFhnY31v4ppM3A/7bT1Fg52hIy
WMEhqi3G+UgsCPbgg3D0hg6EmsqWSB3LzZPBsDW5q7ZZXXNpnntkrB/NAs4+
eVIH/Erjz9NNjBnofJU1Ah/HzLfYP29GEonmpthLPA1WhgPq35owvmNp3x5s
tpHN+w4swBJhRFheRwr9sHdCGjOjlYRBs3iyGlGmls2RNLeYHeqvRCchvBoE
Nu3RbqDrYIpda4HdAu/mHeu7yyM42NGf5HahJveN3LE2HqyllelLBEho+WQk
75EF33Aotnsl06XD+Zk+3ULBgj53Hx/zBn/WAE2QZSGA0U+G7g0ywVdneUGy
ekJkTRDKMLHpjuc+y1EsBu73qftlE/HkVc09GKgPO05h1r2A/mMV/z22oRHH
deasjWXZosrN8o8JI0Vz7vkFASBk3YqUYg97ikv4GL5rMvQ1tMIrh5k/CwPW
+DGHb+X4r5rGmdOmSthkfxgaxM3KhsRPF7J2T2w0m1pSHai+p9Ca66YgDzaI
OmSh9w6ZZc/YpLEdBdrjzozHCad/GyN/sm8bEWIu+umSP27nX1w1jrzMuhlB
DlFIg25GV8OsAyvQLkef0Vf8kk6ELSdESdET6mNkR9sz6mPSXTeJqufZ3mDk
BpH7XioByOZeNf31VOG5/lbP5OcFhfBGdLBbmqHDrTTRIASDzu0MLYHJXqft
PTu/lsQ3aKQKFzlMUNAspDRD//WjIPN8UBiUYDpinGPHwsEgTzSJ2ThGMLSI
p2rKaMUEc92CMVxJHg/3dFoTBOpvCP7UZe2sOJ93fKIS1u3YrRX+wf7MyH7P
u8pVbLeJTuXVoLltteFSPz2xRcu4gSPxas73WxEGP+Mh6omhFejOZRMqaitI
b55ld20U1zRkGSR7v9Zr92ZBX35T+taPRoXuEB0TTcvJcQrZzEE+mjhE8OrE
INf46BUuQ11bBx3Kjv/qbERRZKslGVrVRMmMNjhyRvWbyzMoYMFCQ5knaj3t
2zWgE0NaEFoCGvSQQ8/oCrRQkq+4WliAcjYafZXf31XjYrnLK0RVWrIMz5A+
ZIgTIDLjI91dCio1qjHCcpl/PlrjxhWNDQK2xIjmP2/I+nooORpVWE75Q1b2
TlN9p4vUkmXhkV80ppsjOOW4R0LiFYeRPqSIPgO1906fk62lg8ZgYqmtx4PJ
a1kewezdMJmMNRTOXz4c1Ij/Jfh1cBKdrIWltm/YXx0W8tyUBZldToxEJIYA
dsce7fDLDoKA0SEiysN0R7kaTYC7DIjBWFiAvXkWuzpI2R7j4CHLUoqJUqYt
gNn65dqMk8jlxgWDUGmkeLkW79Yuh7gZsyiKhxPwB2cwgIRikG7PKja7vebl
zOeaaSRM9Ztq+fQyk+z9lpVF38mQ10PESoeyu5T9qbIFeQGOxQrZNKvZN5o/
d0StLPVdBU0OwVUgUQKDKCrIQzdxpP3Jzx8KjM/ERR4PFxxVLi1Ga7n9U9sw
iT+j8k9rYKP5iaaFP6zO+m+9JWfalbD+vxA6fWBAJRGonX1yrqb22PYj09Gf
P33oFoYoIlqX9Nc9qhQNHWBAE+WaNweby+xz6Bl9Xg2yQb1Aj3Iw7I/33pLN
EYenxsU91Ml8L4KnNgswB+EiZTS3/DGa4rJVw4d6Ey3/1HCy7cUHg+Ga1zMS
p2+m6e1NELvPKUqVHNh/R+zdXRj+7u5sL7NHn5bh/yrFee5OIUr3yV+bIAq7
hA3UE5FV5mRApa4MdOyk5XCxq0bMAd/fq/oWaCnt9IqRrz4B66cocOi5Gw9y
EABq1WeqxW8YeM/w0vQo8qD3+SJnGMNwEHrIA8QvcHIMQq6vBxLJARCIeuiD
ikMpBRKDTAPsWMYtwt4aluCOsOXNSajeyrqVwE1JeQA2pz4dtsZhxQjshzKh
JLjepIhzqXqfaVa4lJxfLnW95CYZfZPsWttvsgyAownTDpEDpT9N0w55zA+a
DggmNEwJtYOz4newONokHVDqkklaebcMd+hEkvD/Y6/YJo8u2eXSrOE4ucpF
Vz2NjOpRcMbKN0AcaLjg31NJ4FCOkVDsvowUw8kSc5Cv0i8JQa8cxO+0zGqc
lXKeKq6JwMdkYfIdzkg/px4j7ocEculY57rNMpwNNm55Ib6PgjGgqSpSzAOj
1IYXQEPjo8TqcUU+vnzzpAdSAZlPlDhZJqVN4xrVN2tCScCxDKRR9qqlj3rW
3aChYbVtsYWhNU6N9jNfcZZ2i6N1Cq7JMnbIOQhYlw5odxh1/CBJqQN+i1bl
+OTvoArHROEkLpYb0lVvz5dwEVb8fkHUnqpfwoWhcTjzBDMijtiDWbK0QEAc
UBHuU6uP4CfLjnjImybfj0kUEiedIfZw47U1oRrJTD0huc0pLrU3M4zBQGEH
zAoDdwi0KosEFR2sCC2XpWcCUrF1+m8XDTiz7v7so8IVYOJXy1JBgkLx7puT
qlDq/Fx9QSSqIyrFnFv0yHLhNLy/3w4X9X/giAW2OU6etvnXJHiu6fShirxQ
Z+G/8MiD4IsbZOSBTLocZQCKeevSaki++0eUXuezgIRODU9P+KwxZ9jjmzZG
abNwKshtE17MZuCWNkFywf7/lctrg5M/Hs5TloYrnT+xOHW0K/xppObu2oIW
cS0uFSADPLTXiZJ8zV7Kp42cPbtKfRM2Wm+MFlv1eueafYRHwlvS2m+3l0is
BP4uEbDbOIwFP5BFZjHaBgbmCWihEdCwPyqyGV2+ncu0FyAPZnqRWNUaFtGc
eLTOWMmcVrnk4M4yygbYJUqGFHup4VI437i9J6URVC/SnKMMqXHXtK71iCCt
BoQwrXeI006uCVmo78okr7pzIQ+RF7EkzhAfd+dYNGoPnhHLXH/+I8Cw846O
HeiPvdVel6+ciNuFgcmJ5nzn9eb20mWArVLymp92BU4pbl+KM+ji/z45f6di
IF968uLGi89tl+ysHT8afI4Tf3b/O/WqjKXM13F0eb4hCDNTem/HINoImlR9
/ILFVBXIUr4+mwGc28fSDmcOCI9JWUfUm0BPxAKlz4tTX7FMFx0lmW2fc0CA
WoWlIRG9Icklzy1KOZMJRbe0Z5EW4g7g7g8jzFjy2l+Tb6ktmo460Ri0YXby
Fc2/PbwxRSB9VhA0NJuZMjy4uwDMw1Lb6ctc/pv/cDw09dV4RME8TcrT8jh7
7u4tXw6t3oOI1EvAfJdCNAflpGEYKrZ0NKbTIlLY1Mnff6KCu/lUPOM7TXd4
zgtR1MuCAZUWztNeJDooWdHift/7LYwB/Tzb3DXpSRy9JkTDmyRI+hfAfFbC
ZKPM1wRxN2G1M940pQwoEJqn7OVIP/1COhApZqOWJ+o0I4nxW+THMowyYT6Z
v8+9IZFRBDkSsrcGnKOB6QOwLAzIUOJS6LtAv2uClnkCFl4mXmKmZQHULqpC
YSQhU4CgGEDYzkU5RSp7V0jaMcoOflm8ZgatjtWBTSlPhpkB4krIAtCLJMs5
Jul33srzeMT/R81xnZq1ET3BAOXUz4fFg+It4BxwhcWn2IZpgiPCDXs8ZfB4
t5YcCoX0Z7VAJrZjDKORUpJwLqNlofVbTrqevJvrwzygj31fAaEtenTV+Pw6
K/amEbYJHMDPRXnN/w9zHhQXdKuAQ2CrfeJ3ZVRICTgTQUE4Ifs0F0jzfSYr
oBlAZvYVRICzeWDyFS4iouvTg4YtltHOyB4YRgi/DTEmUq2qzm3X/Up24sYw
z3KV9b0/3IczAKwf0wQJviiE5T97vmCxEVjLdYYO+snHhWZHzcKeGkUOorFo
yZ13H2W5QS5MlCHUKFPaRP+ZoXIT7A2rKhqd8ytmTfKOQ6e06rUQfswEnYfT
a1F0ZzVWuuLIFsRr8quQ3obgFBGc+k+YWvmAhL/ng7pm7hQOfGuu/ZA0Qx2e
YErH1II2hjkCuIclot83NkiUUSD0rO0s2BqIUGRVmQR00oAAKmE3W+QVqlJc
0skci4kFuDnDijQ72/EA0v4oXPCKJ2wBFfcahPDO8Fs/0f//QxyKQzyoiiUS
FJ78pB4uxOTocr4mDGBvxTKjOmqXQrZwASKu+ubfUtd1rYLaT/8qXbtivjnb
25ZwyGgfWUT+s3VnVmkJHgMHx/QaNo0TUt7CjRz+xriRR6gG1aySMZTZXwp5
YhB4ypIoi8VX7DygTe65t1guEla11Hdc0eZ45FhwhOvV6iiTG0aB7BTH9a2X
QdSpDVO80j2WP+O2Yq8kUBXo/PudmVfkp1MsFK1amzVIwVZk1uIOYLK+kHtw
cbFPC7OKn5irWRLVESk5e56pctZc0d+yksVx27/HEbCNuRqEK9QRzw7S9VCM
sjBUfI/AVN0o/su8Y1cSR/Pgx34Rlf9yZZSZCEqihl5wme9XWfn3UfHR9EqC
ELEiOixJmLgVq8pb1BL1iVHcVtUo54uYF8grXjMeBAQ8F8rCeuvdyRhAs6oj
r1XK9EYyAoowGyPfV3+a1MiMQ1Gdw3yy54VlU2bdZh4Dyn2e7iSBn3mwMZKH
vz9/pecyLn+MIWAb9D36KY42v0ks06lvYqWXjd5x2+mXTlkco+qmD92idc4E
tjEIkIq2+V6ryB6XRPJcS6LY4pe6mSu/HhUIRnIxGJ4cXTrnIL3caXKK+Ai4
Pu3OxWXyFptur5hQMHlnBTFCOt3DnyOcA7Xu+sxQ/SKeO5OOm3Ky2UcM+iC/
KSdeMxHzcpvF+gLYFlg7cWe1h+ZX8FSS6A7Wfg1FqYmBLX39Lp7k6y+59iVN
kvty0rvqm1g5eZwyFhLI62IdLsbj9wk/oll360kmD2XKCzFH1qjlGnArIhRE
6gsnSt26DCfQLD+k+QiYyQH5Pw1Fjb4M4CniDz3GHAfqZw0IVZX/tsHMhZbv
866G49uEI9ms80IQqrKYgMg0BKPMRHV+vAbp0lrK+sW/Z10LjFoN8FDN+q1l
fVoV8lbpsXbOIChaVe4ODxmMFnZdmMYzkVmNoBfRfwKuUq43amlNzlSwF/p2
+kLyZDD/UPIz330RAjNeRz+tP4YjE7vo9bGu6K2eJNi5Addx3qCxlDm3mNWJ
JP6QeKOd/dEyesZROAUdzvrVegbFwFg3R2jg1PHNgbtYmnoSH9q7xulABJd0
3jXB3kicTDRHHfCY0UEafeGPBgL7EKRuwMpCTg+/M5V56n0kON53WqVF800d
SDjcnqeORE7yZo3NM2wsrdxm87L4yN5TbOs/CS1n3qzCohHylc9cYHDdehpc
gJsclBDjFro69Z5OzT9WIOlCpkwswJnRNEwk7xqLZ3k4qfMU2ulaSDick/8M
UW4Q2KTewD4SIGe9r4GJwPlTZ3MEhcjFSmNHNZQiMIqK7JBh4RsM9C3GVvr+
4TXaSXhjQ0BjVztWz5aVSp4t6VTwXNFMwOS7220Jn392tamrY42mG5nos6p6
nijyEFd+EEonDEVARfVtj9GB3XmZuw64Uy9Z8fJMWoZ/hHNO5ibIWITfmRWB
dVdtdbcWLRFmzUXry+GCbt/4my0+E3Boy+/34cUXirlKD3wV9PnuzkIoKyXe
pUA+6gfyd45iB/fLYAY26Yo8MVNMMKOuKvigw7yIoleRh2XVDWF2suPjtfJv
OgTwWII07DnhMQKbsuJ5wjjsMkV+K2bgnsuJblZzG6LaAlkhCsrmYltaaYjK
edpYVx+EExRSJOZ3vPUaneUUPpQDZvf/Bh/yGt1CGJ3ZfmTqsjZPFtyOfhrT
BGyDZ2im/HSkTGC/uZEJxEwsMKP9zYEvfiVO6P+R4jkfT6x+vOfjsMqXPs3X
txgSas1aeuUuAFeQjzTafpwc1ppwRYyAHCj/KUu7hpBxpg1OuBcfajPoCueO
HLzTerw9mI9stJ6QL2FA7sPTVGt5zkjIdBtAzTq+2bbDK+GtEd8yRkKlGn0h
pXD1DQHdDV8x0dt5QYGXhinhWKMN8c8S6GDvFXuBG4ZE0BXk0Z1BXMllROio
Zmf5YnPFy1ROmZUu1ptlmDYYu3xB6b7XeouO5SoOd2jRqR3lim9AVeg70X0w
iVhevYgfNqMdPUY22kTWSFYQpXNyzvfBMJyHxQFPT5m/R48unZxiAIhOa2ZE
B4jsyhPWFo/90NsoeTjn9+bPa7lSOKnfcxYhuv74ZFMpGR9AGwVj1rSqXMz/
jdK330MnMP6LOVMfXcEcPYLlcpeNCxnCzZwnwjdFEGzTVEky7ZDA/2W66iHM
8fx/tPw/fq5QaJx7soFJFmSuYIT7tpGGNMTTqH3w1vkC2V7F+BrjwWGbhNsA
6CI6Ftkae/ErMFVVK/V5EY/z67gcp0FBLwSaSwngmmOFrXjxzkHLL+Xmlz1L
8K9Nn1sYkKxiJcImSVcedvS4IuHH3dtdGpX8FP8H5AVotamJ2wEUGuscGB7u
s1wYXZ7w3/FBkZ90MJAzZAunu6AzcLzYhbd9eTnXOHLC9Zz0AQB37dR2X38K
K8d48iV5khhpIifMWVKJSectY/3iHA/52EDtSKY6GeAtFYeXiYlsUASsys1B
YEHlbEKKf2OaVTtrPUZV0Bgl7LvM7OHpbf7qbytbI5VYzO2u6cEZy2zHCpEq
d2M3bHjHK4k1w/hi3E71y1K58TEgef/NeNlvQPqQhx1/G+5DsSOzhLm4Xc6v
PHK2MtPMf31TztIiRG9lcf3NHZc5VbfX52+nZkQgn8U8+uDcmy0gkpHgxRjV
JRAzCVPLLXuoG9yqyX+ti34VMg+CjVNissK5KxAYZWAjj065vkimk/DqdtdF
9WGD0FpnmIvJbUTVV5PduMI5/4uCBGymhjzpQu3Hx4FnqUnLxPcT8ndiUOnK
cihwTYR7qsIVXMc9yq+DwDFi6YLtzdJbGIAY9Ag30theEN7U18HDjFArCDNP
HPz7YN+iGXIbg2oSpncReTkw3dKC4FshWt++rvAdkpDE4H/J2FiLHvvDnu+7
Z/uuvPiuFkBZqQVgU3Ys6rI9XrJtb24XbeepQo6W/Hspbxw1/NVM+cQyz4LC
bNQiLqoiDek1luIebBDbzGF/0OjCecNsPBMjl+pXbbp/mJ5r29N1C58/OWaz
pt6aeRxpLRVl2089u9bLf9U/s2J7fy5mRvzMZCNVqA840QU2Wt1FrhMZq/qa
tVqUAjUxY9iKmpdnYHErZAGOx7RAQGRSrG2G2N2qCcgCfRCHVlB974Q7aUEL
AOfmnMDtX/x5aowMO9rRtF/1xXSxmC4SF5a0uyTMm85Ry7jnnAFC6rwougmN
7LMDcwriDBRU7pvrl8t8155E+R2tkWjZFCFm4Rw1hRD+KJHv3+jzSTxUQdUf
wmZN+zL0W03k72NQ0FYn42JUhY2cdrHyVuX50d7ZiIdgCuI9bHQCSCL5DHpi
GjR6f1Xt9HCh01JNEWhV39wofzFvXmb4Xmo3mEYZ31oAVMaRlEXPKgy95ttT
FVtjfjO75XqvG6x4lDo3FuV8i+148/XEbeK4eP6tiS18peXh2iZmBjVTh9zC
Jqq2gjslg2VQ3hLf2QbUN1DxYoJCM83wIBGUOsYjkChI2Y7INfvAmZOiIVh0
eQsEXhomVRMYYxlx4TWBKbz8KbCO+Mv/OBRDhT14zImLxXRJV6lZIX1JIDq3
rYxaSmRnWOYq5xnsi7GEZBGVq80tTrY2jVdZS9d5CWUGOv8ruECVtCKY8R1W
xVlP2aGeCHxYdbJ8w8W3sJB++5tnhpawpvRXI3KefcKFLwUnlULakSEieuBL
b3jF21QvBUXxDwK6l/XXIVpJq/IA2W4/1vaUnPxlm5NykUz5jK2Dyb32nJtH
D0c5H2jbRjVWay9h6DQlfsiKYBim/MNRYu7gtO5JBXzmtqn3WB24CQyWGiQA
f/+Ojl0SD30++9D0Pw7B3QLKk6fcFODmBikoswZqwXAMDvStZt5JfGpRDb0X
MJUpOHAFW93+YPbEflLFoDaq53wu5R/ct1ywTz608O1RztrNhhUwiVz3kJLF
LCeT5O6/LPI/x7bEO0b93zOnVC7/xVFyvz4rmvKTz2bu70Zi9e/N40+UycHs
gJIGQUDHkoxjNitogeD+A3sb94yhXCCdTbqxVjcCGBGwSRnga1Q20qaWEjBv
izxKRu9nVh//1SzrRY3cQejym2cElcAONz0Qp+mYvIwzjXcG8tt/VGvSUiww
b2uTdchlLXug6K8zhqiISADiRWLbUAElgJhNRUw+El53F86+3R66fsOdetjA
SQYEVKl54EfqBf7UTfIgt0LACKjudML3sUpJUQO3dsud/OA3/YjgVxm3IGWW
CAYxgnG758wutbaeirdboEjuZEeXJv2et1gVAnoAIpRm+/EqKvgEYzXrIK2R
ROcA2Nsz9vGph5sr9+a1HrdGys5sfRkVIV3VB4n5wXA/0UGojkN+VNL4kXYu
QRKV/u5Szq4CfKNZ3/eq+8e8PM19sOrvqPkp+oNEjvC35B3RGmpCcSL8oFZk
oEKSqjVlQFxTBZTs2Yo+tvXQ2nNnc/ZXlI+Q9yK+yJktA7YJCOMS9AtMXHOu
DDfgLF1d+6J4YVnnJ8Yhefu7qcd3V1I83Z9wV4uxGQGe4btsOBBb2p5kXerP
g5mwx+lo0IxXhTs1zLZXVDag7YFExO0yOeH0EsJqEzlsw01M2LPsz6iSetFy
BHFCfxPdHWirMm1aUUNCRRjm74utso7k1qCBXiiI5uuMG3SNjrnK8FCdhnlS
FW1fCHbKlpV0JX9gp8ck/AXIilaCAnaKTveXhs1Ohw/2Cwni6lWXqs0UJPuI
W1vRhtG1/nSPK1/0bXplYYELVhvpzQWsOtTK0GAeT+lb2GTqcNz9UTXybTd0
+8xCS2v3LBMUW4z8iSiEBDeFFcfgmx+pK7K6TDth0yxtsMcZNtIeltLxo4Tu
tLmaeDW9qWsuU3dylO4412l6C0n6XE4H2NZ1l53SZQA9URcRYdUQxaAy5xwR
yAG9h1/bBFs7GRAicPA3UTou9CwmrRB+87xX5pADN/05V4IsOhzrhwOhPD1d
1C3275IMzCPmNRwfECOtsRyOwj0/QQw3OGMQSglp10dSfbVFQFG+1RWED4oC
8LzmcMDYWLqWFfm52WWlAtf26nnpnZZcRMqqOp9OLGy3whNdoSjl8g1xgINQ
DZDco1HRyUYevqZi7ztF+eMq7XOOKx5iL1j6+x8OpGI/4a2uXSo8ptA8Djzd
sN2qaUGBD4qVRGWejVQXk1e9puIt8oyG7n2bNmJO3vocZZManOU6DhOce6kj
COe1zCpMbQbLStxXbA7kLUti74CTEE1jdMIGM8RH0uhk7pFRjmqOvn+KSaP0
4MWkrkusrFxwKkLzkT1XfG7WsPZbFmuGIv98YuWm74ZgGTDDlkxEH3226Rq9
8jHdm2EC/9Pet3KRw/MLPYzbCwjqmsyBxgNW8EjSSHxWTSTwYRXlqJxSi9xk
ys2mQK853fG94d/v8IMiWWwP/8uRblFh8m0X2tszYppT3oWTXxUXG4GFWM4B
kfXP94zYYwU99A+uIUGi8OdAdRD2VCt9wwrx6GGSb8BC5XhU1XleU05DHkZa
7IWSPsAG1j8ufAKyuS3BqYi211qRW/JPlAMJ++947iA1Vre4S8ty9+YC/Zm/
uO05sxx4z7yFE1eJOLK6HN/kJTf5eqSU0BiPXRz8nGMdpNs9PPaMNe7KI6iL
Lj88KG0VKIeDw6T6sCKR/2xHCWMjNTedLSKtbMUEQfd5ey0OjuyDiVvPfZNb
gcSP9LaqVIedSfsFN4pU7iGUCaeBwpusEYRYAG+zdzTpuTYrzM2mlG9OMKgk
HH2Ev5bdriuwweKH86Ti89GYIY6VHc1tVhRIV/XVw4ex77qbxzHcnz5yUrmw
+CQk4OvT7GjK6e2XkMOtMzvKtGpk4ZeIOMNJyyl21/LBfnvyYyEu4qNJZB7K
VaQ3rxH5F6ds00C7jI4aK4lBRBCM/5TR3aMy68pXGHR3j1Qs7dmeAnFxkquR
Y6ZuUBirkmqz3IlrpF24ZOp8M1ErGB6Jrsh5khXp+xXACCtKiATb0GuD1jGL
hoKDgJJB9h+TFeebkrNIxl3/3skrcx5d6qZ23LtqdeLFf/dRDpjvZRkGn0OZ
bWyphdeZSx7+DWwz4h9gMqodzVQuAuVtdXAjw+V39w+c8nLBv7bP4rnEX+Sq
Ia9vH4TcKiX9/GiYJgVLIHnNDbFDzTW+x7ZyTcfBnC08xxj+uobTOe1gKg2m
7O/r3fE9JzPoORhdeshygS29S/pfpYJJYAXpKf9NCr2NvvWNaUOvGVZrMf9J
qHxCORr7ZVtRBdqv6mRPytD2kSBcs+Z/3OisRoj2+qwixhpuhfPlPY6zd3Vv
zejPgpzepflZXNFhzZ+FoZCKZkAaMYA6uA5XpmOzBZa+nS32IDxxdD8ZPVYG
NcZNOpFwXwdNVvVNvFC0OBxYtvw6hkBlEL4eAukvY8LKwWMWUZgirgGQIbr5
AP3Rp+yDm25MknVNRrGTup2w+55AfaFH/ou5ckRvuuSP96AQ0MZWJSwOgo1K
eCqmBXz/Xcz9HGyCsY2xF70V4B+BoqoXZaW/q/+hAM4LqgFXdoBlSQteVPQY
CzakE/wrHrpnpGdjXriht4dkXHrcrORcm4xigkdFcSZr5TU1ZjCehLbyNoa0
rZebFjlPxq0Fv5YjWr3vB0rZj3TBucLQhvCKS5KGg9mjIlcWk9x7mxK7nmR1
O/d5MQSv5TYegTJeKjc/AaxbyuGQvcGgZXYt22x72PTZEs6s7Td52EguZAKF
Zhr1vqVZmaX9qyeyPWS3OOX9DqXeepguPkIFT5dxT+yomYZXBUOQ3MSknqii
qKcT6LBpQO86KMhaXjzw2OjY98GWovRzrWnVqWeBXePMhM52PCwV1sAO7nKJ
qgYEQ7jYAqOYWw3ijh/Xbx4/5xsF+h/TMHUZ1kVVTbRsetrnX/Lr/ZVXvzf0
nwj2RWTJAO3bobJjUXZCMVlmYHqsmAQ50MLDoveFPOO5460uX1E2HjWzuiQV
L/Q+pkY9O7fxXE5Iu5ngoKOUxSXLv/CHNmKqINvPyQcK96+xg7tXSTBz+iVx
X7LfXnp2qRJSlQGUDD26ouvNO6Jv28WnTFfUno2a8bnycFqubowZ6oIBq6Ya
TPf1aGz+LTZMqAMZG9OSi0qsAWbb3VF/ETSMPADe4Fz7UOEIxolKR9tMvjag
auUkXlMcqTe7HHFgSswEYJ15vnp5cCXyhNebO9fCMYX/HMCHjlpWMf176lKQ
3FgRpzHT4/RNJxvJWACeuvklJ8hbKnmC7AA3MzKRaQhxs2Ios5uaFX6LoEGv
4RJY0jU/SZcXBEq+HTrRcVpTNfKAr7kfydRtkP3zZHGvG1RGtzxfvI58nhQy
w6WmBPZPm7qf1BfZCXFbukYZACcKgSNLIROJhTQS50J0/LmYObImwRutoa1H
6+vVVEJM+fULYo99CDngxodx9U4jU9edRAiinkv4eunVZejyCXDGNOaN9woG
BYvrN5hwum0ytk7IVUx4DzVCxf2G5b7RdTIqsuGQprGxZRxd65H93zE6vEu2
ZbGaeF/smUBZ/yOMog2i3IAMD0tZzL73TVEOxSOk+UeMNxjizpHKeDsP288l
cZWHIRB+GNZfiA4hhJNmnIzAehk34iNGAlCs/yCUGnhZrmvoYKTGYB9G5qzH
ln328xznv92j5dDCc/slvmizbeZuGsXSigi41E/hLpfesvrd1xf9mdDw8fy5
IIQs16oPlLw5o4yIGDLK+rT+QAleKb038yGE1TmSY4e6jfHheouoe9IfAIi1
xrIQy9qa4W81Kzmy1bsmzly7dBQpGCjfGJfarPJAIPiNLb2ytHShjRjKb75V
hNxl4E4J9zc+TVoEflGlKHi7PdMRUzviGP8cuRYX7rksYnU5P3TETUet1m1d
REEgyt0EFNnVZBMNwAAn3apYv2JeSGlxhBdupYzprn9Blc/vxbvameJ5PhNE
pZY9+AIbfqRLcnndyq37ivtXgWMELNAt/Oh/cxcMypdHgqE+1o74GFDv6fCl
193qzmqrVSQlUlK/FGiJ/ZUUv6RGqFXZthDJqLTAAs7Be3y9yZP3dhlEYDRI
wpM+XFFPgJ45ttrDkUglr9SpL0+lkMNIIHfur3KaGP+dON0RF+jhvtQM70vQ
gAXlnXyWEA4Oy636KCY12B29lkOLhpgJKFqmQf07uh/Vqgf2AQOi0HGGH7Dr
+0/lLQeue3G3NM3mEUaHOZTv7GIjrdyeYW6VWF4ZXAJsRFbgdgyWdcJp9U5R
CPaNnY6H0lSwWRrZM9+XXVufxyVRr425uYbn+tA/BEMS1SGDOSKDWQKPXVeD
PV444c6Dg3I4vqYKEFNczdgEfvzHjUtsEg5UqVBNU0iNUOazdkxzocyb/OCD
mdJXjweZmvfxzIzR8toAKluY4QaHQL8Jh84+GF/h7ZTyf+dd3Z96+dir271c
QAJ8A8e8b8LZaEDN9yLc4H3HCGdFKTVwk3BC5O7da3F04kNaINpCE5/PGVMI
IGNf8Da9ToCW9TmG7d1Isufp8IUlFOndP+Xsx7j3E5H9wXWoLP6j0rslUd0E
YK8N+FLuHaspT/9bbt2Mlnr+bCr8HEbbj9l8Sed43Ls43FoZYolkqeTbNk80
FvcHfwDyrHOWQSN2UbbHVDHh8dlsUgbRwD2AelI5XuwfGz+4lIlrvHosUhJ1
7LISWHFgXcR5U5WjZEu5k+KlpQ9DHXFirMZfsoR9BN91g6WKMhescMRQ28xi
rg9bs8jwhXcM5g/fn3/Zf2bJJxpt0GJ7hr5q0shtuOXfqbmgQ29GZWnykQVR
V2Q8Wv0c4sz7ORsZDXMU+VqROagtV6B7iIJVQDP2nE4sIKiwP/iPlA1ntgSr
X5dzeHMB26fGhF/79Qlxkt3c7u3KTabeynCYGOjHI3BiTOTYfWrQ2DBdoy6O
d3SaFbyvwHNKIsDE9xMD4MGRiFTGLaL5ySrAM7XPMWI+S102GepsuBcu1+/3
ukhJFeoDrkb5j5sgKv61P2yoz7pjv1e+rPQ5cXZPQHb2vR/I9JxRrNyt16Rz
UfSk5wp//L50TCnqh4XieKV6QyJZg3nFfMy54peEdGbI+T1dEU1o3M8UYguo
jkLn1X08CXOwZg+bG7mKw9SUWbtm86sGW1fFMSkj36/Ay/H6oqXDSRjsJMg7
K0XNLHC/sba1XSqneWa8/bk57NX/QZ6edf8UASDi7i3WCT6htEgqEUsXBUYX
k5PmAf+ZFm589YDD6Gd3xj9aQhBf0+giz/LRiUSdmik0eCda5Tft08qD+d/Q
GM+/UQ//nszdUz6fqgV6kH4RcZkQ6UUeihtfcyIps6ThoZPVDfDGGYv5mV0d
ZLJeJItaMWv9e1DQBeFfFb8t4MgkYVIAJAb4i6BrtrlAFlEwT3poVutLQrAY
xIsC5qJoVbD9GZCk8iPbxxcihTWx7Zba+SqQN3eyucqLEQ/Tx4P7HyQ0vlT5
M1kJqzc+VUQkpy+5gH22eGhZ6wIoa5v7jUSjRtZLKHw5g7pIY6THgaVq6pNy
z32cSyUCdQ5Lk6GgmmBM58p+Oc7QQzos/8IX4W8XCD3bK1tuEc2cFChl8FiX
F+Kv0c6bkSuHJWPI5CHthj6+yYiUgijDdH6dP+pbQijjzSLkEfLYBAbuH8WC
Lxy+nJgjboufO8tWMeYD41A+n+fP0Sq+uFsBRgBr9VDV799Gu9OXRkXfB+Di
XayvaNjKRr+WL11P9WiCu2CBNioCiTOM9F1OSBcuDDNGYrD7vIKYHzGranaP
aH9vkG3PTexcboZuLSBT4vjLjCCi1LfSs6Ig3KwapmqXyzOGeXJnrYnzKVhR
ZyHTqRcISX6uofq03j5Va+IsHQAOQVSRBJjVCD1CMfGDc9wlrY96zOf/vksy
OJoTd+CqJw9oWhRQo9Y7jCmJGRoBwbFBTT6zAuw0zxlPpAzqgnsTuZkvQNtg
8zLq9REMVGwTA9OZnSHLCk9fJin/F9p8gCxtTBRD9yWM1Dkeoiwfw9L5/BqH
Vz/mfYy6KhYuSo9UH0R5voJz2l9eTTzCf+tmU4aecHh6LnIFqUdNQLG32bPZ
FgHgBBJPc5f9XW1hVm3YTasyjh8lv+VnnrNl+hA9Z5Q+58JlBtJ+pBs8rndm
8MlXZAFtmzkPpjBqlzpcuy0kqRSxRmJaXM1w4Ab17kYJhTQjX4ipdWEfgJQ8
Q2o6abjOin1Vd/++Tv2Y8cBemI1TyFEBzXYqO76YZAnPrHTLFUmWoPScTIFB
Yz01DcnECnpi2gpDFGwSS+diZFOgCssM0Q8VI49s3zWgdiNUq3wqs10Akzq/
n8UMmJKKSoTjfDB6AZdmlIccTcpNEY733A+jCiWdB3IWxi9vT3WSHKsFcTq6
dMgs5yX8IRmNPUxK3oVLxULWl0dUANKZi6zSkb+BVmgq1lKIogvFAHWtroiJ
dRYySb6rkJD1lo1napdI/GNUBN9gCRt2ylsAAm8PYJaP9D2Jx+5V3z4p56wi
BYSvt9x7kC+EB9rfMNTMbZGAe2QBD6KX0LlmRKmilUneugvbhVOR2qCsfgqZ
1J8YiDfJxa7xfeT3b6doEZKqX7rkLxGjbkX3DvtvpV5PIXcfMdrTUFY4rFEg
4XkMdxfQPQtVcP1ZLCXqFBD8ORiGsernhiResACPEg4qBProq93Mg8pECUEb
LzvO6NyPDd4klkaSpavYMTR8Cab0gPkER4P3cOT8qK/2D159trfVqSkK6IzO
wVGSIbJcL3aULHGidDBKCTfTM4g7ksvfEt/W1b5rywseovVOTNGmj/i3BLe/
LmN48V1hZ6yvmfxuJFGSBQB0rDiAeFe7CHJW/nsXxEmJA9/xDDWe5FprEaMD
JVzmR/XgDgUGVn1jTjP6AiZb6rZy1F05CT1aGCqlzExuiP7lNETNDjAeeYxF
39qp1e1avZpihPvl8P8MDRRY/HTBUp/bQpzpf1sl2ZxG03hphr6OZUknb5Mr
VqV4k/SimRsHWy+FQDN8lWLVuOY+auL75khvYKs8Q72LHFl9/1k52gsnY5Qb
n6SFrPtZPJifgSjoMQM5yKvD3nDlV4gC9jkB4oMag7iJH4zR0EcpZ5Y8COaz
2Rjdgb7GwP6UqQ+df1+BrvYydNyKb3gb8sTvQOf7WjEkoNRzTW3PX2Q9dgXu
+uB6lsKGmuisUyI3kq7BUYbXTeXF+z+4KuAFImcpoF4BvAb+uiE3vEeTPQOB
DcZ3GU2TolAcY2XjKrlk8vLAt1g1FB8k3gM4YMHeRQV5sH/BcAEY5ejVgr7P
7ewuQVD4fukKRn+MYavumhFK6lVgmpiquaQ/TR/A/3gDUj0+Af4oiDQavzza
yodgbuGzoR5qoUMhJdUoIxTs7dCN6/m/1sx09GdVuZkbSDFZ0VvRtbDjluO4
F4iTMp19p/MOne+gFmQA+iOJLsninmuy3B9ioMU019r6YCEyRTX5fZ+mOj8n
5KV8ReqvrR4qFZsJnudOieJrGljtyAifixodtSqMmjJs6DR8e/yqEh0Vc8Z3
1DNHDlhQn4Cv1lQ0kRAmRvD9ks30M/2RlXw9Fyv+pZDlvRom7PohROc1OlCw
yKXFTl0AZmxf2pMLKNxnH89qsp1YouXM6+6tjltsFICKf1v7PTEdJmw/wcUg
PX2XuA7GWG6agc/iJ5YVjc/wl4vlZ8zR/kupvONjShzmPTgz1/hEVpl2ksmx
d9zBT1etD7rewDDOJT/ScVRCtcAzL84yzrVLwlgIvc3VkKhT3CVVjdK8J/WX
wdTQImLWUDG2uVu6xwUu+CZk3SoMSNvdJBXBY26MCB0mkv2XihGErgxD3WRg
HKb/H4U9i0UvfPkc0NjBpEjKvhxT9PO1MM1b+37Thx51ifJmeE4LiPE3+q3B
HHJs9ENrSTkhl5AeBcO7B8PfVZ54PHJ8Qwo9XkGxqqjnTX0P2xKshbxtbubC
rx9HTy5qzvSY2kCT/ewy/BBkaK27enRKs6ht7B53g7exo+vIeDtJ6DCsqSmK
Jl/AlxTeYfwA+1llJo/751vZSsHkdjFGmbibeXlg04YYGynVyHmtxVhqByp8
JjmztfhtJ1C26hV/Dzx7/Bjw6tLsy2GlhR5jtnnZZJcbOYjekMkWmJ52s8To
mg0jelM5bRHg7dSA+mRKIxkCPQ9ib+PCwSbvJB23EkSWCyI0OldXeyiZge9/
x2HqPz16F//5MeFO8LpMAmmz9K4OBI4qXNN34xrVMBDxuc1gO19BAAaiV4b2
ZldFfqf0I9ECK5uKpggMSE0Chi3d6heIS+8XnLlDEgSThc22xtoT4iy95ZUC
RdaFy/hoQ9+4Pzid/qbVzv9yhqnI3U5lUxLflwBaLJ/YaF2I8ToVNZZYhhYu
i3dG7F3SH8pwD/N8EBtN79ZxByL4uHWhsba7blznsD8NXyxmpE1FIYKqHHXf
L41VVoGstPWB28yTvFWbwga1bQ2BhvIaXZ0SEYg3v/U3ZQBe7fafEEVUzIpo
H7G3bniqHV9+5on5MglZD0CtQf2cSnTqVWbsZ9jl9CG4Qb8jnwN17igjnmZk
4Vi2y2kWk21hpL6GoD2fGEbSJR5Q+Te/YpB45KRW8R/xCkSg7TwWAMYsaDPX
+TsOduMAma0neyB21Hx99qI4UffaBQ+5T7rvz2Bg8V664Xr98KHIMcFlW3B2
SxAUg3yvOiutxsB6TNleoo5LtPn80GycezM0EWX5FpGMEyEwt7OtIylqxurN
8MOoTbUYcVgGGJ3EtJaLcLtkRlKzL97yqXY9IO4mV0ol+iGwrxXiNYLtmB3A
dh5/HMhM8H3r2xtQmjnHWSv7YIgoKLJ41hN+Kj5rFgRToKZETwDZ1ZVwvhB6
TKXVUf/YfDkxzpE+4cFBsUL3WbBLMMsDWwS1leic4Qj6fLpGkzkVSkKgUPOs
YCp+hpSjHLQwhvWBmqzPEnavxag8mtQxTII7px6sE9cNnSsLpcZDMfLfyN/i
2n966BzVjlctZb6HI/O3MPsWQ/1LAOBQ5wqp9bEs6Am6uTIP+QXF1ydUToAl
YFCJL0KTisUxZeKatJR5jR+40Ae9IEDfwYI8IbLVq5mMhsDagSr2yKeS/yi5
lz+Y3QhV5qgysqCGq+v7geRs1KQV3zm4sY5pNprAUC6IvSZGj6t4L40k54Iy
B3Uu4T2hFwiFpMnnkiDn0P4sdLpiktzCaKq9MHua6ZVPgXCZRSzzsrTubl1A
KcI5gEXkyDcBkLvGhMYEaFjoXmojP78AFwO7qGBhRxPwARkyP9337IyNlVtB
4HuTQjKe+erL+7wMCkOpo/hhd9FdlyRK159zJwoVpBzZu6xLgy7XezTxH4gB
jhhc2WPTjWT6VJqZByzXrg6XGFJ8zsbWak9PaXx1u8tH/kwUIzbbipkUvh+Q
Z4AyaQ9jup9RLlV+jixC0WTin2RNef+sR+NaKLy2SKIp2Cn4/9vKxs0+cwnn
uJBoHByep9bSEwBGVzXCDBwX7Bk0i947d0BvUpcVCVlN91K8nqZ1c2Llo/TW
EEpR/fkbRz/hVhFLWqr/WX8DGvgqP4K/MhVUsyqF1vYVHJsocbT8zbldXfWd
oOfQVeaD2nwEvEgvGs3M/0VH+JBik+9erLtdtUlQa1QYiw6eTMmG1y7H7fIC
76WSVWtlLmwTR5dtkq1S3tR5yiiY6jnT4pacgOF/Qscu2jkI/IG0eEpk+iQA
BCnMzabcOxGEEXFl9mNBVhTy4WUAERzf3frjpx8fKedcg2uZMvEl/U8HuS1g
FyEKgqDrHhIhZGWo8hbXYNNeVKJ0xdWOP0XIh9D0AV44Ue7ccVuD/DopEeyS
z0aneA9dQ48Q+NGqkRTtN6uKaWzH2zAwPeX8OalRichlrIDgrbZWKbuHIadi
RS0QVRNyxBVsE6JnyyvGMvrIfmSDWnfHGQjVDKKLN5FlAf4aQDbRZmGq/qME
kRAZdv+uVaqY4u3JXm1bausEoGeWCfBEOcGcIsPhzab0VtzcRgUJReDh1DP/
BQOFrxbA5UwiefNaYrX7ceHZQJes/4lr0oGxhgDxVCE1U4K+3YbrRJy2K/o6
N9NvucyInpVtqsB51U0kqYdfNygloRv5hCPbg1RAE6SAAmRTlqMStygczWj/
qGQV7H4zcvC+daKwXhd0ceY/QQFbwnT7y2bYo4VfG1MLQwYRBB9IZVOandbb
ajOY155hqlBxKxFsAQmG/XAxABYBj88PnhKYJaEkv5/MyoBP83wpYJ2WTvh9
O2N0ZMpU2m1xWHoIPsVyk6fqOetTn1BWbikk4xRUumE62Hr6FK2phK0L/cFK
hyfBcYX9KPjz8nLvb7YuFI0wta1BBRwklILCMH5tcNZew37mDqJ2qR8q/dpq
74mFtlYvTbESA0CoT0mqUeeg8DU1SL+EpbOOl5wyaassrMjOtTwUhHZS9EYC
yc/E0cSQ4BO+xmE66HJgh9oBy/FTVY1qYa+wJzgn8wAysbfk/aoKViQwRX2H
zGukHzhYVDl5QoKGyGtwXw+Bofe5m9Wy3c55nqheRele0eonMBv+m5nPY1QW
4hyr/Lx2xJfl53+w2CfGDfjQ8dSvxvMFjiriBDUBT5bvbnirlPyU8PAH3eZB
7yUwUEAN7Ce68qzfSAMMvfoCFfnY5x7itOwYbyhWdVCcdIG5vOZVL2g7UTH7
DD2Br0b0p0lDp58X9TNXqyaFGZdvEW5hn5H42+88ZqQ0B2l64TfOuGm3JlRh
t4OiYShJ2N/TLquGviYrmZ65qXlnvgv52GZN4oBZveLj0nhEyLzr00uNXEyA
IcX+LTQ/YF/W1tMVlTeDSSPxeaP/Cd5K7qn3jgIo0ck4aAipfpNN+MgmHU8S
fy7sCBNd8yIBUiyjbVuEmuPBFEwA6+m2rte/2/k+kA5KTa48/u8pf6GJv6bf
tyhSBSEsPEDXZbJjLor/XSkELYP1v2LiHfUMTvGNYkC1FuELb5X3NPe3QF3e
/dQYUivw7xinATSYe+a3iCFGrqNkC1qYpgEsIM3+0rg8dIUKCh/FL/IkiRwQ
XMCzl91It9vftV/pHbHgtN1SkcRdK4tydl0aTbEbd60pVYolsN1N63M0gigm
8KrLmHJDtonbjgWrA+IuHCXClUi0oNcYIXIPCIiFBdKFXr7m8huNLEnFh3w5
UbMRRA1JmdGnPQ8+8KyrARe466iD065hjVCD+U5/RvON/OFfADFb3m/NOyt+
XIyXo85YI9yZiCAm26tZvzp7lqcq9Mk+8cYAUJXHDcn3BBqiKBGmj1KvLDki
FetYqaMOfE2tBLtDQzx4hk5j3wLJM/qC9gH6Dezjg3EMHbh4E00624adn4uc
yCR389TciBFBCQoeR0lvbxxJTtYWOHpS85UJr9JGKHMjrXPzPRpJ+7JBxijS
r+g4QUX8kDkjAMqM4zN5Ge+0nNFLdbc3HH8tv21M0N/CCiM2KFzylf34DuUF
DvSaXY4G0UG+boATN9VP9ZAmoBaSuYFnXxakJLX8HqvZfwIEfhTuxQ9qBKe0
F48LbO7o9Wix9+yDIUTEC/Yurpl1tpci4sf2XioL/28A2ZVeRAfYgyePc4mg
U8LjcY+jtdvaxMQ4Jh8JEWUPB9g0ou0fw14ew+jrM1Fo9b1+0gid9XBUyKZK
OUpCJUqSg3+ucGJ/QCuCeogEBJ2ZUNQyclHi3IrnLMXq/MFy9ryiGEM7RSsi
BBZPmn5viCwWdCt+lJyvyGnWUyKK6lSLZckzje+9HWhmkuL4jmU9ntp7zsra
F7+lBLkZduGHPx5lnojOs8Paki7nMSCeNiK0oBzM3tCd2OXWotL6Labn2ro+
9UIQcoV1pcUdVWR9mX7gm5GD8eXK1badz5j4MT7NybrMLRa0hwu6UH0dwO4C
0POVnKRNYwfBaKgZZPsm0mDWTL1f9iN/w4R/3Ctt2txx78SwHrsL4YjKDnnh
hK2WABXjOVTKiYKIbTDgEBvIkG8hnrIkqW7D4SI4walxG/Hrc195Uq9AQ0A/
SLRFc7JmH5YhHPM3/MbvpRmf4wb4a1lnIqMGvfeZhzJRuqOPZptJDOpPjsGf
C95xBaLr0uuzuOqABCvQUNW8lnztp2lwN9JLAkBu2fdWbqK1Fe9sjiaD6WeU
Q3C+4c/KPXJHMmOY226NdCXmzfqDbnKnhvtOu02oJFTf2e/Q1yNNEZj1O+Vj
P6MU4d1MpSX+37YRqTqwPnW/SanvB+pSEYsNyFsSZ/bAJ3pRHZISLEk9Uqr9
WFQXvyMY+Dft44siPx0iXem4EF64ycEqFCWt7OMAU8/KuvDo5IX9jQAJClEr
lpu4NYR+MsYxA65RiVfOjIsbKHjlwFq/fsUUzz3SxO0TtVkUh+6LOlUxVtUq
KNECbB21FS4CpKEg6oxXQUNSTXKd0Tpik9VSRREf6ansET09aiM9IP5ttkeD
/EotGxqn25XuJ4qL4r5TthQVg1qdjgRRLQ8WUmtqWmrmjr3ni4/A58xlIoE4
fVAmRfdBNgvqcjxvOZPuxH7xttiglEn318P05tmFX2u5K5LzXryGB2XYJJgl
I4v3mUobAnLzAMKfl0kq2pD9NubFb4s82dSeQC4d9jhVtFLv/dX7ZB+vjGSk
Q+ro7dA6ZE8WfyXE/n4AB2dk5jt6PUrK9pu/4i1XMZ27JlsdYbAQN09hg5bk
2p3ciTlxFsqcDAwt4U7fhgS+UvJQRTiGhhORrb/p+kVqfezB3GZULek8u2mx
33i1oaJ9fDDe/T1htl9CGEA01EiLQpMFaFd+e9EzA/Bav5BhdKn6N50Yrq9v
YVC9A3X4Q7xezTfKzNg41y1RiWnI1cGMfcvfLQy3fTF69JdsqHNiSV6PFJ+w
OD0G+kXUkDOrVCQa6EjCFmXII2ougXzpojA/BAbmjtObsEN31g79Xb137gu6
10ip8PL+8A6aGjMa/7xMx4bDTq0Rrphb8GC3dWdTRS32j/zPNfwq+sZr9hWD
GMeYMbFtcekJs8MnnEQvvbOSYYQfz8jBXvIUYNF+4G9oskcBF1Fo8J2+x3d3
e6dAvEWL0orSGo04wJyxZebogPs8/3ELyFwR6QVWl3JZdGjyJjCFdJER9F1F
RJCtqYmJqEjHNelBTSKqs/akSHvLneolNd+unvifeKn8WJ1yv6CA4yhjuBOz
vmAw68uR5ZUG9X3i/vRaOCZEqAL4xGZZTe8noYQyZH/VIO/ckMKUOfoThI6s
oLqPKBp99ydJ7B8e6BFxS5XiurWkeRjkaoK9xkvhy7u5QVFB+J/kYHS9HIxW
xeSfuPxFXQd1rh0s5s9Erjs/nUMRlfSjHnbOfde41Qluu/L6Ga1rkBzzLqRK
veLC5hpIzCLj3oh0sK6fcLpGQyO8m7O8lwUubWJ4TVYMNiET3SwMajU1eoKG
Xmv99NYU+BwWBWVgU+MABBdAy9X+IXIwmFMvk5TlzdY7yL0zREsFxRasdSIj
zwjt5Ix8tBnTHvmnHNyX7OZfsb3eB7i2MfwCPRStGwYkB6AQkTuZdKqFzk+e
VilP87MUIixHQ5JPwT+yyn+eI/3lR6ZyMXMK98hNVXkhxDPLKeDQC3CepqKu
35nxPEGtVMGME+dQRz1PaV1ujLHVYSQzJwUviO99BTG2QqoEmi/TZWhbmwLs
YTeiItBhpaudhUbhq7D3pvZuOFy82taVq+92ZPdeAJkZu9f5g7xIFpuZI2H8
Vc8hQeWqNa936uXGNtHCBk1sS0M9Y78sMTIZRZHamXNqBrVlcRKOVmyT3Jq2
e3fj4PzzX1zWBexdR6XMf4aIrXd9kIfsUaZ7ry6XpaktHrPtAgF+lipawcHP
ygfT5t2IJTL7LmVgf17zbTyDNniIcUoekxKFT248pTR7bZfYsSGNxYqAoG2M
QOD5C1WcpFJvBjCbcwjjfwPXloCOfFVMwny/wuZnPE5EtF0ueUtEFOkqMuBZ
sD1lG2AMYbd+nCRLhlu/mnUo0853YuP1Bkc3PC1yeACRnWvgW3kE+to56mvr
eZn/CF803AsybUjNsnw5y0ETlwpPMMjmiI3p8ndvAP4PnJ4lOKyzSIfG5LEJ
zBODPK34Id77w9OArY+1OgKARLjysOqHZrZvQyf9eAB3U54vZIPqMECswVUj
dLU0nnY3KjNkGxlHQerBky6nqfRC/SELFf9s0cgnLJGtivfKfbteV8N8XyDB
HOfYEseEzXrt/117btkLj1XqZEsdbLv2D+UyY/KnV6ZG6w062NWzEur8ndJP
OZLkLFbVo/D1njyj9IbFVCJ2B5/uFUoNrP+LSKw5nSdARPhfZ1kJNOmwqk5l
VDSbbGZvWLM37lxWt0Vc6AEoc7tmQ5cquRHmHy+ja88Y1tkp5TanFfkbb8xq
EyhLsIeR/5OqjG7JYY5quFju+MIr5pModBwRAGSHjIrHEPJymz6MQt9gRK5t
cuP/KSyb0WxauLXMlAJcmnt/N1R5Gn2TQltr03b/B602vyZZgbgB/Dxc0KmD
glOP8YD/4yRmD0lq/5yG4n83n9j+Q0IrTRNh3BePorOiY1Ne7WSW+k8SliSZ
8Zjd67bsTqQem4P7kskd/esbYZH525b9ULZLWzPqMWqEmFevqqh9JnAHt0AF
XNtfCOi998dl2dK5j9HiwPNXXZlz7gKyr55YGc7TIyhhOhXXsNaromrOagOq
7SYEUOeQbZ1bec8rBAjSdy+kq7b6YIWhMRqtViq2Biwh/l3M+X75HHHxAGNc
Jdw5DjKw6Sp6qZlmiMglj5jRlg7a7Jppp+aU9fgCUYDqRgYKSVSVSIbmtHYD
i2D6U/y54GOtIYSF9C6fqEMXLt1WJ7pS1gQwuWkOThQBU6a0AEJ4WumS9qAD
wHVT0T+yqNRcEPGDuSpEhAOQFwWwt+QaGhg9ebxOYkBgBshPRFHl0KC+ESdX
THM+al9GUsWIF4xyyb11bby18JpOelqW+wl3bNmO8KAFLmWTMIT8PKBmX8T5
2FOiCJ/II7M2CJIgI2OLZeqG6yxT3Sv2j3lZoHcdU10hhUqAL/L1p8u+WIrQ
HadAFLri+1c9+rriI1WoVlH7PEdSxT7YKOpYVvFVDgXK5mmrt37lXvUXkqtx
Ee5gvf1s5hidF8y1slbladu+LJGxQLpTm340tgJqUz2+zKvyhWWF8u1+pxem
kWhYRUMPr5H2MQL7CHrgCWYNMNZpMIldNEnHFnSDAJVGQLKYyTqHU15NFxPi
LpeZ0lXizSFUA48UU4h5RTn/TKEY5KKh5dNqUe9A5c9q1f/7uI8rZdErNpcx
svd4LhtZ2a1xfHGuSAd6onvPk6ZV4DrC9s4IqRzrNrexFClyTshitGRZGWWa
TjIYIUQ3G2Ged0ogtWux6If3JWr+jPQ0qDj6vpY131kh8GTD10JWXxUSlI5W
OaPoNZ+kxzEAXj6ohEBMV91Mi02UMIM473VEVVFkKD9+xbRFYeCMBeNGSTuC
UMM+tJmLQLv7spzadu7CRVnUqVPldusspYEukHJQD6RtYnFHQh2RYfSo7hsD
5fKIpFaIDGMrZgSrXCzH0Ce/TPfP3OoFWPRQoO76Qu2WgivR33OoqZ8QstTz
O22mRvtoeminJ7APfIKkPUGPpSrtdLA2pQF3MbNRcsieZgjt+wLHfU3bZmTq
aVp2IM2El1e+1rQw/KOdmhAcF+8Vfu47cP5YVHizeFi9Msti6BH6zu6/1Pza
C6ig8SNaXJZFAry822qJNxM+XIuTnVon9HXlIvPrPrxyWPwzA2NHJtNe1BSe
qA5SZFVJe97suzdbnGKHEtQtHcJDWXd59yGg5IMLP89yMVtojA1e8wGF75KS
SDPlCQHeF/Sn60OFN5pjaHGKaKf7h/WIPVGlcE20eDdIonLWDemwvanQPimU
HprUuPCWJLTOBmlNeZEBZqzOzE7mK9bjQvP9txFpQTxZKD4AFXMs7BLLrWJD
m1GW8jKiZOm/ASuMszuzV8txw9kbo10KA5XS72EFQ/1efo6tfHEDO98IPLg1
yw6yP6SB4g/lwk9yQPiSV+Urbxpwo3ojqy/KNpcIUBuuYVqv0J5h8cLzUBap
K15pUt2wwE4Wx4E/sejBlVoewuAFgZTnOHkAWywvOw+rDL3Vv9AraGO7Z2Ak
Ly973vUsdO81QsLm8Hz9qKf7qMxRAgpu8SlED00RmpelVdJi+ediznBWUQH0
Wn5lLyTMnUh1qr2m/+63hLpMldtkW0LE0Q6PKZwZ/X6cZ+rfx3fgyrm3oWWC
eZrEYShR48mMfqdqK/yulrUz4FzZG1/hoziuHUFvzvvx30E4BOSy7/NlR4U8
GnvvpLV3snAh3VBJyMTWomOeODNTVZnNHOCT/wVLPFQ5x7B4L1+BkN04E7zl
F7pWVfUxcXDHmnNJ7gCTxKl6P3D7647DsGvmvQ+L0kzwNek0Qae14Iza5wLZ
BHgpt5loLvbp9Pl4n+Oq6M/59oAf1ZtltMmX5Gjui6pEhaKBdZzxIzxt+abn
kzjVXvFxpuLS05YWx4GvlzyRSDXvqeWVRLSL7LbiQyDDJ63goVs3yd/LOoqP
U/0fCeKK8pOuFff2mNYQMxXRpMQmwEqDkkqWv0sg2K4/oD859xi2ld3vrx1X
f1H5ZkuxKsSuTXTzWQJo/IQ6MfiWi6cEgLEO9NmJeP1+V3802qq5KMN7TzWY
xgaKpQw8EgQlbMY1UdDuR9/WNa9IZnKW2DQm4YP5fxq7ZtiCrnWm58Cdl4/a
zYDHx2uHErZ/yn+T4w4ULU05deT3z/oE+t7aIJueBocIg6iGNojFkQkhReWO
eIlc1yHZO6tTz/gj2YifEf8Ll7xxkrbH/rMsH/teqr9kR/qbUTCxDd6aAjeU
rlHD+BGcuysrz6MKKPUA9DQW/ASMHflDkyifxWHkm0aIJMNxobCggjKFgpza
gEZhbx9rtJJq0FnsIXPg9lxNyC+PLDsyTsdULZfSrHeQ0TpFMu3+hOo2m+9s
Q5hZ7fhS18jUYPzlqx7BcmCUgPCAZ/mbV6n43jnoiYJZRQyUYcj3zTEBJoAZ
Xo1zqaAiZP59C6FmYy6hdFWlwLrDYXBKTfXP2mjEdBZ3KMkmnV0irHYWIsvf
ynErDrPS4jQ2pqbFedhBUhBn4ZIvWrad3WdTcUrfuuuW3ehq0FZUywQVrjyp
efFzonspOGlAG0hfSzdi1Ogml33SJKjwXfgH8ssAaPlNPDRl/8XtwiJVrZfD
xhAbb1qkhfXT1t5H6Zh17fdJzvCHR5LWcjz4ZNWgNccwpONc4A2JpI6CM60k
rjSxiCcG89odiMikPGccnAz370n+C7WIutegGfDrxnw2dCDCnfPARQL29u17
pdfaNIFq0Nowi35mY7xparo7lnX9qRaRGeML4O85w+VT3B/WFmmyGwnbfCuW
jEgl6inkeNHsimM380HKD/JmQPzLdiyF7GjO2GlfNuatiXoAqFT+6PqblMlT
Xuu+FWzMUyfYQlfod06pzWMWC/XJ1kZBi/B8FozDPRlG7e+6/UOUlEH7be9s
9Dzs9JklYwaAkvzSsvou/kKmw8kuA//aqAjfSZKhWjIT7lptCxPFasmvDP7Z
P5JKfX56L1vk8jCi3+TNJvSbDbE9TOhnni+SdSrwiWz/fNWFNFT63U+Z233g
xWnuPtXDD3J0C2wwJmRJTEvSLbBuVGC1uayhBF5ebhTpPkGx6wJW5Sp62rrw
IQurwp0d2mrRwAW58JoY7XQ96lY1WqAaxIsJMaEw7dUrNPbgu/nAjvttxJ5s
S+IiIHNc92unMtY3DEWUyOqPb9U1sYlydnu93f0lb/wsPEqJ84eNGH0YLCw+
pfRgtA28hu1hoMgP3nQ3CEK16G1t7PrsL//Efm/jYeN8R0RzSv1k9at4ELYf
2u5eKgAxrzWgkl6rXjnVC/7rPCeHSivyw4+oGOZUjrEaMAtqT7vxRl2arl5g
y4G1HajXWXCMozj6boosLKAN4rfzEswQwrzOcHOD7jBD8c6hjx67KcrKKbP2
KcwswmUYH0lK7WW76dQXV8Xjc1C6O+V36T5dHbhekHYPXGof2OmPS1TcXoe+
vQroyM9odHWHy+FIJAuRnsNYDpDWScLtvBpCgSVCUuJBR/L95y3aoQwlz1uw
OFJzqBRS8P9T8nKsbUS46JuXsV8HXxBDO0RhZWvmdo7Vj+NNmrAbkR+gXl1W
7RN/kG31gz5PXnAyzE+N0gDQpDSHyydMYmbRgGh4ceTPgkh3GYTvyoJOLGjy
MnkJrgr9btTfD8iKdsiSlaw8Hsdwkuw6uVQvhoZ00rbC7nR484VGvin7z27D
TQbF46S0+uqPsGMc4Rcdzfxlg1SUhMriiPwUwWMbxpVqv4hUusHLe6fRV3EU
zwj89ZdPtkcXONmY06+sx60/sVxGu1dlpVAmSrfdITGhmTR3pI96msXUdWVs
EcNcebdRV8Oo/8tMYc77ftUFf2h+zHL9G2VjhQq3kvTAhFA6xyKnw6bYjY2g
A3HDgrlfGkXuNOx4mnhiP8aYdeF0yv5DJMJNq6lzamAnA8jwAtBFUWHtFCF2
LYz+jvNzEPD1gqv/9OxjLYCVf/0joU3DkXe62QGwXcQ9ZTCLCaDe4CL6mKov
5GjOu0uIKUl91WUpEWMhkcS9AzShuHo5INDxXIyvp4UUjecycCv3ARuLRgkC
QxtyNGchejmbmXrvfSIjquBghW1uxzpBvFh3y8N96skvARTu7ZKTT/gYzAPE
yWaQY8Tf8GlkBj7150FadZR92alPHL6AQTbMcUOyN9GbfvJJQ5RR6eU8+B0+
aoQQyUqfGLuXIlGE6wU1gJGXySqyfML10fcux90XM5AKwGLHL98NLn10/TwH
jb6cDP7p17RWIQZKv73ghnVWpI5aHrwlhAI211iOYVS9j7HMPN4hrKifSKRl
wJjxl0hqmznX4HlBavqf3kM1JGu2ekgOxs9NYBURy0brLeCtTbcmQPy0Bqv8
gAO7TAfykw+Mx79UW7tB0zwoOEyV+QhqcGOBKYqqhDaGpKajdDs/6wbYvHSJ
KacAiNlvSU4NP6Dmqtn36qHICA8nce4NfQLxvmdUGbCMR1s7zWrSeT73hf/J
fgIMUIqveumTyCuVa5NCnOSijH52h1yGNqBNXJ3tdp4D7YZAYEKESLrlj8Ut
BT5Q5vICYdmar1DnMogibR6GCSHdYGSfKea8xIQAJwZFGXVTuzqJn5wb+50P
qDTimI/lJ5A/BOsK7PWqzlJLTe+7Ew9pEFKvCqM0eto4L81M0clQbCMIdUTn
iVW+K1LuoAb1bJF9sy8Bxz3qaZ1o5QgwYkL07u/reVwBJsPrvliQ0zci4vfT
wmRNX6QS3tnkZTo9mmGuPg+sNdZY81CQxTZLmEtUTyO/gVvrRVbusChvO6pQ
7PUBxxshCbyxjrMXZbpPdgh+8Msab5GRruIQcH2RTmrcX7MOvIAXMVTJgEfs
yJBPK0mvFnIjj0h+yV5CLlyEdYx3QYvh/dBxc0t8gG21SWLXecIFjZ03s+nQ
/gq4DW3eOq1aa+GGCVECxqyGg+TQiN4S+qSs9U+RjVa+MOGwtBlY001Nrq/M
GEd3xXPI2LNz0t9WzTVKujYrGvEH6vtFMCfE+2LKRHM00oFckn0r8dIWuwcb
SeVkpGyo3k9if+NHe93fyFGROQwbNIL+y1LjopXaf/QOFbvenfz5UJxeXAK8
aw7kTf8F0hIx0Jw2zKE4duCtncfDnafnRmlwFiJmmhefeXdBNiGFJZT7xiZf
WXGwUCtfHEBHNjFrg1cCDpC3y00FuozmqYvY+/+tTKnjZCfewiDQ+tblKESA
ffq2x78PrlXbR1lhIwHJUrbzyEJxGaefWy2Q/k1wZh3lnUX0dEVtawFxomG0
yNSk4A8TInBl2JljCetqpIszAC0rPMOvyR4Shom/RKIHU+/1ariRDlm1Ew/O
OK0qKrH9ER2yEzAAx77hIOIHzBj4qys4Gv05te7z8fI8Uy6IwLk7sPK1wMnD
/3Gpb53SLMs+SMOKUkQvErYytFgGudN6afm8hemn6K6puSTyGd5H2PX0UV1+
pZgAaNrcMQIoB+Gxjw2mSOkRX2GtVo/FE9mWkXZWEctLBCwamakDMTvaJ3qQ
ZaM74aqkuNsPcjdvXs+9eOUjioXQW0ZRz1o+y2IlUI8U0Uxy/8uhHnmppp6v
iNKZsULKdjzwnZCSijerb0ab03OSY8xvCv91jhTbXGjuIxjiZ3iFt1pA3WP4
7g6UDk7d9uSwcFVUl3CxMEH3XErrq3mfM8UokWPEb0VYZhlS1Pmr2f1xUMjK
v3owmbMy91qGsYHIoMW2q31R0EmEORNwxMmPYtXf/0jjsgobt3z9/jRgYyYE
JFlcLQGjefPP+PdYLkpzA7sL4AZvJ6n0iS7K+b+B5AZ5voEeoo1g7zReX/zO
RxHNaHGRR8+D/D1ckQfXqVop6DNWmMwjO2Y5x70L8cLaBfAbn/5RxGQEH2Jz
b5ZUVMEjqt1GO91naJFnAUrFlhDgColiPLKsTxf1PMPokUnwFBsRCxdaXcrO
adgHTjX+RRIZ9dXPQf+IR9lkH3bu/2nUIZyF29JzspCIDdrdfP1Lcri0Dg/j
r6yBlGAM/p7mhqf0rT6pskVfRDxNzTwTd2ToBCZef2BgWpxZcr72y0kcrfXq
AdXgdfykcVbISnQbz9hA+hw9gouHQ0tzpVIF/HkG4GajRWKVhtt6IEMlUECl
dhxpSCHqaKK/tQlBwSwGO/mYV0JjZ/ybK36uHZBx7LSVrY4rJl7KEBeWK4TJ
7VTVRB0otDezn4lQ7GMLHVJwL+Hu1PAiyYTzm7I49BJ9PCc9a+69dKASSwuR
c20T2GhxZVjc0z01paiTiPO+SqoEcs7CYuZGxN4t63fjpvGjMdoMcErBh/rY
9em9UsyAxLiPe47cpRBM4Q53nquDDRBsGC3sOyRgKv7fEXuZAKrYkLujBBjW
4aVKA4ydoLWDSL/SeoHunImSumCgyANFl8hZ2Fx6b0j9KQ3LiZ0dCr00B6Og
jybgKxy619LYfahfD0tRMKVPXKiZAQJHolyDrwt6Nwi5mJ3rtWS0/2MsdqbV
DTKqXWfjVIRL6+xiseEf2ar3wFVVm9JsxyTfNEh/akcDZiXgvrQSpLQdqbCM
nVXY8WDLlNwYaN/EqpAqA0vGkkJ4kO4sKGKJUO63tUQiyij5z+UKsNiyUDgL
CTtMQZlfF/+0UQaGLHcNKX0/slJK4yk/ONetl7FNzTzyzDatGAGZMB+ZlwJA
z9WnJHbuTQsvFCwy9wxzC76ZlUcS+DR94Ijh3wvgI4u24K15lW7dlBSVfOlU
s5b+DvPAhvrehj7xfcSZFpBrjYtFHfcJ9i/WQxSvOTqaE2L8skIagm4Vnx2P
rN8d1AWfsGa3a9g58IGvXC5zTMqFZi+cTGuumcN67mwt+a6cxEyroDhXHtE5
RNVntLJA5pQZYugvKUNfGOCNtVbEUIFaoKgOThO7HOiozNFS0POLGOiRw3b2
3y2G84pdX/3e7ssJG6/873lhiAnv/TVVgEap2Cyt16peU5LfgZjr1YTXxdz8
hpYZSfAP8TXFMIeqRpFR+vh2yJ4LqXFlAzJrUWr+5SxYbreb57ZZmlzp4sjZ
ALK+We6X2jVOFjNwy0yzKOWbVdlJ52qQ+LZQ8ZY+BJbBw2fECgIW0vz6z6YF
nOkmIxoPoKujadcIkOim8o6bU5VsrGHGhxc/bXD5Y13pCqcSqjVU396H3BHR
1awnYt8uaYVnMddTl0hc0Y2gQPeEQ/8XrXMJwW4b5oFvf9WqMvExNQ3k95rY
VtmLMPPmHxHSBuC8V754djG3LsmhYZHRRIDrS9pzBkANOaEGZw4DOSMunn3A
PT2Le/ImR7QzaKNv9QCm9sbL7Uex1CLbNWML0G92e3yvRjeq3/PN9kfmkQX1
2sIG89vCvTCQzpODQ7mdiNMvWP1SRmM1P/wPvqGrRryft9w6mvOQDMjKsAiP
O1McbslLHrtLkyOZT4WK2wuaTnIfsj4bdLZXQq0YJdGpEq/z2K96D2RhCBOQ
u5V0Gg8r9eiaABgAsXQIti4irFWeg7CZNktIeHBbN1etn/ObyGSREcq+hoRM
94hU51+7X9y9+7mV9Jwng0TbIpU2LG2gxXjLkYRlYI7NHQL/pNmNsEYekD34
KSuheKcNmr1nlam0V0jJAHPtjeKzukoE6sRjKvH97vJUbquNvRgmnoXwuhz0
lYbtlm4jFHX/L9zqXzba3U01Hn/O73Qm6fQ88L33dYl3BP/JljDyeIN7p2go
nf/QyI9emMfjRk0jBSXVNlKDpE6m0Z8Scd5Ej3A3AGHRNhtnJZdZ+0uCx9Lw
nNXUHexxDsAHvfkQyjuyhC+5nY5ga0FKP0SQq+UNbZ20sGGqu8ZGrL4mgiHo
a+HmkbxwbU5NyELH23iTeZMDkGVtOwmjFhyMZaIZUw5+YkJVW5JyB3R7eyNi
aqq00CbTNsfDZeK1JKCHwC+KR9DxPFFvqn2hM1ZEnRXUWKwh2yk8lFyq7Tvl
mg9kfgqWx/wvi4OHD9aD9y4GbUOcohqF9k4SKssbqKybcyr1Z60DxS2A+z/Z
I5L2M9u02uBwNg8NMnpAETjQ/SquBacFVGIYpyXufhqdweQOMnRLp6N+8XVB
GNoZEFtgu2g2Hm0RjKjF63He1+NaCVSAjNAbk0oVKmlhug2Gdn/pRQgUHUj6
GmSO342aFOwsXZ6B/WzaI46NyzRnw34c1hCZudWg91egtTzgKt8jNH1yInbJ
ZPIsRClg7GMIMfCFLEjOcAZEZDouvsY1BgvkCi/l5rq/L1YGalC3yzp3lv+0
NIwr/upJNspxwZ4WA6DZAjQqRYx1znARclmBBTCmZMvgsEGIlGkL1c3zCwZ0
w0MFeF0d8td84U52Bp+5inr+4Fju+aV3xcz/NfRNTkb+fpZnpMnZU9NRfVKF
qCtXb8zrp/+MHi8afYGjoRQ0bFCVj7ZYpDr/GTcyXf5aoziBeMuNKraYs5Lj
ziUC4AyWG4wIeK5r/h6MSKdmTEEvyPNtUmd8pfElU2NHiwoPvlzEYIvzHnq/
f3HCzNbQNq6Pt/MzFgrfVWGrjdz0XN29B6LuXEAFszBdpPyy9/6n215zUqV2
G0fT0X/PZUs/rpm97WBIuhLrJzQ+NT9HbyGsMg+ONAIuPFHqP/zHoQ8ImeqC
uwnQAqCkONcDB5WEPl/PXJMX7GT7gd8EuGqXBrv/iK2NvTcUXUk4YtOYrv7F
PhL04ShjeyQwTWBgPc39Dnp1scoy7X2uctjl7C9hb73VEmQfifX2vIcWU80x
zRl0fD9FOD2tAjlIWqgS4kWwxT3U9pcCJSh17DCPvSVYmAtrlwiz7NHtkTyp
gPcuXlqIv/RANFtp/XDaBEvIuZWj44Re1+GelzQCykY28O6acpSleH2qKepe
Hcz5mGaLoibjavf1vzy7akuWwZS0xyNyV4GM+3u9Q8chawmG0Gwa3Vz7T6qm
GSHOzuqjlQiVORJaCdTrIVzsv7Emyh9zLRhhXMzakJqi6DsxB0x+h6GuiT98
v+6qhEIUisuZHqVxvdjl5LcBhx4/7/cBC2V0GbFfdGa8/kfWsDQQiY0B/JoD
xDj/4Il0VUI9Xw5WwqV2Cb2oPI/2FdUuIkpgpTxDOehBSEXR2jyyTkvrGMKd
dJRR9lyi0ycs98cNQ2dQ1JSgBLztXjxxECdJFu8yhmIDqN9H0NlPGRaKW4tY
9esbz6XGCISgXoDUdDBxPhd8HvZI5R1H5Y8HSoS7NGJiUkzaU+PeAk5Pn6vw
KZ/s8DR74k0TiphHQm5ELKuk+nrLBV1lkwGO1enbiiX1lo7bp29nZaRyzaqd
wPClL0KRJ04at/TWd7Ci+vzjJG7Dat32+unvwPWj2+7GUfjEBLzSzNJ0K6is
t5+2sorm2EoklPVuU7lRoaLXl6UM+3N4sg46chXziixWbMAFpt4EIdVMDC1i
gZG5R0dwaNdpUxrLTt37XBUGG1XEHQiPfjwBU3s+awEmUHR5qPHmo27ySSLr
sv+ClEKv8j5hayy+i1IS58j+VP6DFcSmPUx0k5CLGfVYrdgYzqvBDywdRo2V
P7RlBnyORc0L6lyldYVcnaZwOP24s1cfzDIgrJLFiaChtgpDoIjFW5m3g2If
SbmxyBwwJeYhT5r5noWzEhj/tFsBgxZe9WTihOWonX9ESulUgsCNnVmrf7T+
uKM+enEkwUiadaSa2TeqLMIUwktLr0LW54+c2FzwRZor3vLhRQQR9bTpxVPF
Mi+CILb4GyzdbBa708cUXHen2IgQ1m9SlMdsdy5fEXyGJ+JLYN8Qe6HWAAxS
8TpOve5dYQJ+OGIq/18TNg0qfk4Oe1WBs4CAwYaNQZdEJs/TyxmL48fgqjPH
53UJ6zsOnCu2q+gyFeM9INz1XBoS21xzPltyVMQSJj0BpoAhz41c6EOnzpKL
5Ba0cw9KtOZbP8cLwK8lmZhoMpaIKvMVkltnpkMq/Nqbf+yZRiB/XIPD9J5B
PW2ZR/kdhW3eZXjjxs6ZUhkmv2dLEQmSgVt50P+w4vvomqw2VLRM9lUQPphQ
CTyPE3FbM5MD3VVuL/kq36Eo8fn5m8ET/rGPwM+ff9mI1XP1OJgCtAvr4u/k
vVbUEaoeSuunJW8hobuGxvb4pbIlZ+/M+RS/wlRGJREx6kL3K1MNS6HNOI3F
6EYrCpv38MGZ361H/49KokszEbG1jfXTiTm9tGtC+HvRlsYd7pQvb1ziGEPL
SxUF37lwHA1b9kwdNQ4KzJ8YBooX/RTnaFcmD5Y3rbOc3y+UuHx68U+7vsM4
w360xFqqRBxfzjgzYKMbfkKp/PpDczim6LkzLHQW6YnEN5d4f3bf3WepYNA8
3ftMw++xHdGMBscqVQVzgapnFkiHVJgXkk2jdNXCYkJ6jjyevcsHEjCvu1ov
U7j1vszlt6vGQQs7HGAHk7leI/4IW4C142uRwLY5fPl0gWQCWn/f0xQE4qL1
lmU3p42TAo5VIU6dVEZKp0An5rExqtDV9nReyBv2sT3iyb3O4adzfKQmzEm0
U7T19J8uboM6n36Tuq4SpAkWY56jL0xskS2fKPyJsFOen9IHUVDC+YHPUqG6
TstAFNDDmOUwVSqFxZUrwpe9RZIQcxI1ROTHjdJfQ4IW432czWEuSpb5Z628
0urXXFfx7OpUSWScOoyIE+eWOCdKSd3YKzeTw1KeLx2IOXOO+1BbXJa5plHv
VvLnvXgxpTDTSsszCc9pbDhqO7KsbhS98K6Lf5rkhSDELVJA9nmB1OE1NT0w
bMR63OfJz2M5ZtxF49fakis6EU5tWJRcVnnHyipWhU7DqHFJe/bbz5bD9/qn
pcTM/fyOT8wZ1hu52xjEUuylOCDL6WAKpfaMkOMBXKOoVaTxFgMT/m+DPDhg
FVEN1zCsDW6DwC3qYXZ4fj+QMLSpTE6JeClPeSZdn5PH4eKbJ6P50r8hmVIa
LCYANv8DKIM74BUsZaHFEG0GMMX+DeytdfvAjAH+Xr4PG66nq62J4NYDtqKd
9A+EGJzOJ14i9MCz5UOcCdy+WbYdgXsHQ5RPIrcMqgeZI3UowiE51A2UhTkf
vNtV7sjR049F4KaGzWwnQo7KFr6Y9yk4TyOsNGXI0BS6/ThNnqO6JKJgJWmG
Cy3dqK9Ct9SYQHVGom8Y3ftMhxoR/lSum6cdwlOkdTbF0+60nIYc3TzVYxvp
uRTc9+jdS0+HHW05UqAnK9rwkd714lXrp8MXsvgLUN9hcS2TKp1UTKULCVhK
f5CYSSHkuZdid5bxcYmFN/mbKcdSrk/kx7METrQg+oqntXpHNYo1y5AYc9yU
O1e68rw/Px8+CgmMeEzyBtFxZR8HqylhaFZARH4N3FsfI8NAbi0xUZ18p0oU
uzoBP0LqQqY6NPj74hQRGFZGJoZgcWOxyqRXRD/+uK9Dpr+Z+5hQ1kx7bnBD
0M+9JNfzH8ygXuJBaAFLU5YfmYk7Biw/do7MoTwjUaNVEirtIcO3THPoqnQj
+7dIf+p9uIUZXFTnjlE2lHzOVwgTNeMZr/Bh+c8suz46jhNf5Lpfws4A4hZt
c+Bwv8yLo32nZksN7PQ2ttdjUpL6T+KyOibdMYv3TEhmDFMyEUKFju9OU6K0
DCLlEOUs1hHGLnxxgfax7vwmsc7NYx2B3L291yHqhCzsB4RSw2ervIQWc3yD
tXUm6HxTciC+mvIAIaE12rL5vm0sXiOqFCWnTo2ejbSr3MFg9rwZyLidj5gm
RI0atsoNi8+dkZXTaJ6uH3YkyFw2Gfx3t+bDtjaqhf2e7ZCG+UlKACRdUmB5
sot0vQhmmQmR72mxyAVQz9482AdNZ9Fcy0wbeqyCoaPSiSfgfuMGUewkxx91
8RtCK5sdW83FqfzsIHHKiX7iBrSYavSDFMWBzwmqNTxwIpSdnmk32TsqS3ET
HycmEsl2YnnssW0bNhv+kSKrKoLT4OjNB6M8MuwGUEgezWk2Us3GXz0US2ya
jcr7nUVywxkG3uhTpeBjes3Dcn+8N58RkrIHUNca/Ok6NoTca/1feXaBycRm
Dce7qssmWqufa8xeknMF3gqnj+4uo6AHNH2JkBXZaKKjuRkPE4GRVpR9rxlO
uP9gvLzAUKLFW/Kepxbg4oWJqpXhN3Ad9JQHtQeMkxkO5zati1SfoC8H1CeH
W7u+uv6IVZbjGrXtbUrIL0RHoWWNJdiV8npd6gz534JWzT1E7IDxjIRiPBxi
zxS4fS5rm0LkOfwfaj+Np/JITn5t0y6MCOpbK5p4q10NtQXK9x3mK82Rfn3+
9c4LCB/aFEJB7Ri2kDgopAgP2LeXJTN2E5Z9fOwOzrjHzjHwgE3zKcqJU6q7
iJAnsv/YZbs2PIo6FJAhYo6bCh9eDDL0zLMMAoBaf0CdNo2FqvTavsSLdWur
qqy7zfMWtLtS+2hv5uVnzDn+oR/zC7SBRiR/sB3fdpUC5JScR64P1gvPiOQT
VjhCvszLgXWghz1VRGHqPdU3Ar3Vzs9hfqOpnrOsllmX0IKmPCE/aOD4EeX0
79obP58Q8j+5q8kSN6OmCPCyY/lp4DncIXGDLl0K0arHv+s3toQYpWzPfPpW
S2OwlKaRJEWvSHK/6xiHTGKU1ofHX3IvMA6cq8O+8PAa+m/sIfyNFA+VSFoM
dueVbHFRDDMPo4X9edorboEpcCsKrLkB05k68YaD13FijphDtTGpeID9wR1D
7EQGkZul9mbxnoV5ABXdhVNG2HAvTTUd1ehDvq/Zjk9ZnQKx4NZj0TtAyXAr
kWndGQftxn3BdnL90AAVuwgTtA5+pJGUEcV/4gAabe8cqgf3i3MGBvxN8KxD
cu2p/EglgaZyQ+Q9/Q0cLBOTzQiG99R97B1cNVx89dXTJjaMRttXWewmS9il
6MlK1NhRQtSaOSuy7kHzVLiSs1Xg0KybdG6MDfFb4VHkZSbsFoFjUdm9tgdw
18JL/10iwuSl+MGJ52AAwsopsgLHOjEmEWoCnVxBpwrzYoIjWig87Us2qAyb
xjhQ6m6sZNgodgFmkH3EfYVxDUrbvn3+RzWNsj1FFdJFGLSvHyUeAEIMvRqr
dGwOAS2eP6os2Ubrf/rBwMJdkxOAMh6wd/WhHFVPGEfkeG/7puyT8M/bOb1j
ffSCru/JkNFoPRCXeKrCMyD8yN/XpjoIwNqaRPAyofUrw9PMmC2Ar+qA27hK
ILd66koPXJs0ShC/9wLLTBDg7W4qboqa3MTa2nGZ4ySixm5xK51+XB8g57Gh
iPSrteTADuPQZVcz8+V8o6MczTb68yGLmCzgT9GrRMZPQpuP7oxFwDCgnekT
DoVBSMavwxoF1fIgr9qOmtVA6+OnLt/67d+mq+sm3XVCaiAzpD1ndgpnRKeN
jM7Tqt23hUI0G1atbzQTPJLLANTnbAggry2aFSYhMaCUT97sz0Z4YLQDwJ0i
0CLd9g/jtVo9n2iNG+oKhIwMMumSG+f9hR5HaDjl00Pu0ieG7czYaNtzLiy7
uecEnwev7fTJtPjDtCEw++oyF/TPEd8rCM5hKbbOtXqaky5u6zTRPokeOf1W
nMVe0koPv1UtiJdYkHHBU79WOueanzWu/65XLQaEhz/h8R114daf8CDIb2pd
lk47dYX1/tIJUtuAuy5xIldZO84voqWCu0NnMV792Q6rtinXoGE3niB89e2D
EzocqerK06d2cHXr+kjkQTQq+gBeVZSwir6ibE6P31Pm9Qzn0r4Cgp8EJ5T5
lznCsriLGTKGeJ2JERZG9ag2PPt55NiwW4zc/gavwX82Q4/Kg/t1lrJPIG3P
qMC16rwXrQCW59xZgPNzEQxpXi3CIRNJwY9jfAKvkaubpy9NgDnS0gdbllFu
HE06ru9PrGPAe+77Qm15YIEYt88NoBv+gJcwpcP587Fx/EaHjYgG7tYYLVUw
ubJrUhbswlBMJRT/0rcXOkWT75ScMPxnoSpc5ADJT68woZ28qklQajXtDdaO
9fvSstYw5T+RdEkh/BIaS7pLMvTl64YOPXVb8VEYNvwrI3ITi1OueOSyV5rL
u5G/qtfvKU0k7PUO3DDf8LqF/1cFX8zMZcdZz2ZWoy1IZJHsAoG3wj5MA27e
uulvpUouLQrtg9OHrbpGuCQB0cVnvbuwrWhglAroNHWslxu0JeRPHT2yLTpW
di6jBhQM6YKmK3/oJzPClYb9i2JCjnpYQovrgN2TJ8tJ9/MSVbuyTT/FDdK3
lkU5G8CVcjkD+hi88CJOYsV4aZMvSXLx17MCr/4t6GTEu/0hGysqOC/9TugH
gcq8iHLgm8o0H+Em4d/puy7jQaltkmT+Wow+edvRaqP0bAzQoTyta0++MU02
5CZcllu7nqJ322AUTsmYgi7Lx0XwcJXm+6/Z1NQCp/KmAzn1otF3r4aCDAxP
9K1WJ13vNMYrJtz+ETzDqFSx+z65TXL6BATGOCqaQPyKDrJZFT0I/PRVHRpf
YO7DRRd2N1mcFOP3xP+RK8bqLF4wOZ6ouewKZFWUHf+64peUHAckVLq3Ih7F
6eCNO6x4Zo/QJYOaz6lT6jianip6o52ihdzT2GmL9u4wUtsERHZA7mqhadG6
bhk3MgYgQRlI1F3x4GCNkIHeyv5VUxPI2mx3zfZGAXd4U3e04Ubwgx2wYimT
L2L/FRp/dUNbAfdV5EQebUoZQv4UXydy9+VCvOpC5Ph5LAReRMyj1nUDfEvQ
rjvwcrsShCPfLsaH8sk4OPxEXVfTpwK2456CP/vRRWOy/SywZOkTWaU9w2sj
hZo30OlLCOcYbVc8nJHypA7jtsS9d3CIjW4vKzPCem+b7aCVZZ0U4+M3Yo8G
rKeXBerdibDFj5MIGq8JBbOFKPoDPfdHqAfVxB48q/7SkWEcXpdtTwWd3bhX
KUy065ytIIsH4Mf2rOAMZLW1QaJnYdh2hbQrQemOkkccJ3JGew9Veoz00vQh
o07wo2MdzbhS2fOehgrz3mPTwjgnk+TwP09XckCNA+UqDqLepMXIMyNuoZb8
zsKQpfnIZm4JyDPzLdQrjWexJqFBo/rDvP5OdlmT9bJLg0QvAvxUPFTyyO8q
jxYqP1vYFq+Gh//xQAFkUpeECjWSPkY8C/qnosXbWtdLwn9y8c3dRAcImNe+
Nn4CYZ4NE1eCe5Da2mhexJmw9OLqrutGiEh+B4SmRU/wT6hAGVATEiYrCHg2
9KFYd2VHiRmeCV2JoiFWyFzs1jIdNR5Cg72YlQRMUcQp7W+JNS37MQ9aw7N0
QlngbdsPO3OrH5x6qAvvhRVgDDjSueJa6gXATfcFVIc7kZHv4Gl8ri1VRAW/
S3+gkGHRTFLT9LjVKjX/6FC4zn6+J3oQ1pbw1o2r2+U4zIpmHff9VS4JRItn
lDlITXAvfyQNx6u8iwoWJKRp9Q6Q/PJr71qKXi2oZhaUdINRSCQwMKIlU8f+
XNxDgTYfqXuJqDU/6jEP8OmaqYTMH8KYpeCCx+j7DQRId08bmrSYhAOAShpX
W1XfyzKqb6mXSrr69oigP/urE7r9KNpCjdgSaH5syP3CUGgiNok95I5yqAkI
xk/7RcSIRa9686/+aqm2G1QzhlFQGAzBrneWjZ5h+cdETQV1yCT4V9J9z+Tv
0MSSk6ajdQV/v7yDr0NxjufywtsY7NUUSpc0WhzxGQJV1lVxlke1Kr38xmdv
XL7aXc3Wfgf8M5tCQ5XqbK9DSa/+p3obVkQZEAy3oP//QsH1uX+36xUq7Yzn
6RUD1gAPZ+zVfYI0yZl7SBVoaypYsitoM8w7AVzn0g+2IHIYFAwUIQHUmPWs
buqikPQ1vqLbgIcDeVQ0bO+gjpZ/3FSaSHjSYlbVqdE+0y6Lrxw7e1e6tpLE
4D3waXuPVh4vujWtYNlChFFFCXup5pXpHpWZ5lky9KChtKl49Ka769TXMDdI
8D3vhJW13YMMnAhyJEuT4mn5ayCBNGYGpH7wD7zaOG6fjh7we4exrp6sAxGR
zZg4Lx6V323BcTpOTr+5zCjym+SXrL5/p7p0EaT9dxx9W6PO881SIOgdO+dR
pFZ6EeFIVJn5GOit5sv1jp1CPb+pHuZB8M2DmXMcgLeu8cfomNqnZ8Jhq9/D
zt3NXNe8pOWV6qI4ynptkpR5xyC3OJgD0N5JqEO6wSqLDNR0wxjKcFPKBQva
FSd2ZXChaefBAPPrq8HUOdsPaUsUCa5JDKVVFZczodzuUNjlJJJSaPikiZfB
GrkX/gfc71HPqxZkm25LodZlxQ+5K7fKkyEBIHFG6ctaT5g/bgD+5Aznjxeu
BwV3jZQvEwqGIC1qix1e23m/tCQbyW53VM/xewJJIIvcreXLhfiv9Sfv8VKU
vwSL2OQlPKq0HsRQ4u+eXc3DejG+yNgGSmV5yt32FWTJ+jtkArNDRIOgT+dK
DlKKXf1LZmDfUmnRjBWyg2DCdDeQxEKg4/PQnfubrPa/Va7dyMZXP0MBvmIT
oD1F7FhncTKMrGv1LV5l2RYHSJtsIMGfcKAHvNGO93SWmBRsTdvgBdP8ojoZ
xwMuzydtmy1nrfGqciBThNiRuVgJ8IoR9NE00O4PRHZbpTLmDUyLedlzlaCd
T9TFIB5feSVVR0wmsOI0lr3QRa77t2F5FrUxfVzw5H3rmdTJTua/5rOffQKE
xp93MbUMFv1j7TInvaQ62lirjLZYM8rKnFH0HcyTKdiqGfnQfiCNnlvdjEhj
TSvOXSp+Ol+3c+8rI3o+TbGCNIfXtLHGuQWUEqKqhZ19lWG1QM3wka9FcW75
6auVC+gk1BMnvMKkIY7YXklgXXntsjGQ34KaBt238W8lV4Vg31sdqKJ5aZqU
3AZwBVEFbpx4TUrcAtlPqDvlgJV5T6DSHnyUUxxINIZLHLH+l4MeaakwPquO
aJNXiZdlZYHq24SSOmXYP5WnK3J6u1DjX/+OYDQaK1i/cGOuVwHBo6J4hgiL
mVslX7oNjwClzzqu7AaME3dIjFXkwyo7BDniExxZ0jPZHN1VBr/ziEPsra0e
GIl28WAS+2kb+7VBv/+gptgutjG1a6X36eNCzayBybNy0ZIxVPeevBfkRk0T
+zXKtrDSsI2xzBA8WwcD37ke/qzCXG+1G2VLQWGX47ZXHLNKIMZ70pXKtA5t
U4A1X9mQNxPjUFbDPges1WITzszDcPKSJZPRJ/0GUm075DqP+eHcxrOstJfy
8N/CJELUqhh7m57tuRcKkgarQNiB4GAPwj1BX7AbRzsrDspU5PPCGqEBrQZk
mmoqtY0R+hW2PAl2EZqP7CGy4qZ3oY6ObbFoDMto6JHfUApSdF7UPRYaM4sP
B+rjj2d73Uuv7YPcX5CpxKO/feA4exoD+TrJPCHYn3fsftDvJthJRM4p6C4f
HM1xk4RFE9gW0+4Kqf4P6sbFBbBUcOshMRU0J61kfzbY88QACH9fAZl0Mcz0
8zkkYQlcUAkN+pRHpAIhX36dQluNiLyCt1ykJDIVj7DiP7IIktXjabZ66Dgp
cq6lLzF/7ihdljk67t/dODeG8caZQkG563xZeaPO7YHD1Q5Cyc3Ld4v/fdNi
K5/QNoUlsktlwKQEbbwq9d/JeFsfK5MROoZ9azLtI5KWePojZ9fyvXUcaZga
7OIIm/19h6pjoM9VB0MgjyheTJFM2IbfRm9Alcdz5E06hTaFCi/f89mXNuUT
eAUwmKdD9nTZ7P1BNY4Q5to3nqppg2QqL2DLHnSxGeZwdCwneIZkiCHu1CXR
MppGnk0FHAL+S0SQajKsUQak757udwkzx0nHZY9nOTs/ZmmnBoPF7zS7YdDk
MyO6gIwQP8269Kew0ayeDYOKwUtlg7QPaI5qRYb0nqeiRzrJWn2SUzzzJ6fE
J740FdfEYA8D3vT3zuj5glXEbbQF2h9a83OOM5HqWBXRpNraNa7ytlSn0Vxt
CPImuayITp32xOWfPG1PjXfCzpCrfcaoLx6xqyEpmQNmUCLyLwLbW4Zzas7O
KGi57VXYFBkfAFAbWobcYDzdMOiBGhM152kbSTGWT3trKPk7xwNhd1LdmdmB
2tePerlFtTy4A3GdQZUskLTCRx6Ep7AiaCRSUb0DRVwVt1q3O/WXLu2VX/Uq
FZpDyMY/8boiTRFfIPle60gNiwc8N8jP7mt2tW0e33zJCMaq/3YhrrGE5/p0
Jc23dYGYJiO/Y9u6ZIj195SeB3oZbu3f+V0IB0XMifRauHN3odyqnA6xqVQL
lg5bQNnXFa/mfRIBknbs9GIMRfImfX+J7QtRDmioECqDp6zWI+BQXy6rL+hW
B0727r+7f3SSRzTSDZzAyMWuHGL7zPhNWfqEgO6bX1W22DZImGO+1l5TUVSz
gKVfMyMg0ksYCnRBryItnTn6JWxuMix+eMduQcXkO8GcfVn08c2DBqH/j4Xt
u4BdeZl3/KVmH9QoUlrNtctqos4NeQ3IBoWS+EZNevkVzC5qciPwHqtBkRjZ
PDAPkRqCKjT78Sk6AvpSu9Y0zgQvz8E6A0d4Ov2jFpeY25HuYqS4ZL+Hmqfh
RwH9sp+OA0AoKK6BoTzIyJjKaiqlzUAGhAb0eK5oTDUfLdu1MkzyHnKj5f1T
wFeHYnn4MyfbHe7XKn+WnxKCVAzn8FnvReCZloF8NfeRoFfxg3QpnyOldPyG
wDyU5xxMhqlVFt67Kk62JpHdPJO8cpPwV1HPbHWA1Fe0gDD+8vzjK4J+5rCY
BczAJPs2ibH9/tflJfKyp7mmiWhisQnD2XO1QiQwZQOBfS3fy109j+jfM3XX
M7ihqKj8RxWMT9Lrwj2zpWrNv4DeU0WbC4MNR1NhTzt7TWURIgXEdpW9MnXH
Ie2xdIVT6NvvZP7XMFZoNWNviS2jMQTzjdT/xA9tt7p5MfqXUxgp/8uQXjou
MEGeHB/nWLR+Iy/QuzFUks09D7sRRo7MZAF2dPmoGfW9JqJHXls5dnUCDGh7
n9JA46BcjoJZlCFSEM7MthdrgvQ3hjxyZD9ZFzDop8MBzPlOp8ulyhwOXIDJ
M0lSKEgEtLs7QIbUFCvKQjNchJr4MRlXKJJU2n64LQgiG83oilschB5rDIzB
Kwvvb9tTnBAj2Se7dXJq/17ri/HmbphQOS24Yn87pvrK7+3H1NVm3HFYIumn
SEU0RS80oQD9bP+JopLDSb7IHp/14TL4zv9P2d8Fm0TuBbg0bCDSyE6deEYz
Yi04fkIksF+P93227YD+MrU1A9W2UPXtvrraNeW73+Vks7WhoFEKl7vsMaBd
AR0QefJnOJ9ERvu0WTjFI7Z0q2B2gYIGeOuaqw2PtCENrCOJvBCR3+aKnwsB
NNFXGKpuOZuyMqbl5zul75m+RftdwogwPTb5KBTAwSLWR8QgsmZkRKIkl9uS
5nMbCMKMz7EzsFkNy32gMTvLWE58WY9J1r3ghv1FSNGHFNent71O0L/hkAL+
VezG0VqXjMuJ4I/niYX1W2CzdQExqU+m3ClAqqNz+53CQcWZRSFSUet1ebXZ
y3Y0t5dZvNdQSUjaHTjU8tPveyKoWfXLCS6psEQ5dX2z/gsLk+8RU1k+UCeS
0G+6QmmmnHZbG4tYMo2qQRM2Q4A28bvuno/adM3XVLk2njCJ73avOQ2ZLDvL
FPBMwnu0RAh7ItyC+ADTxc2A2BVLJv/Kk5pg9jhK7pLjuT8idXN/abeiTy+U
PW/AZNZcCQkkqHY9sF/DFClJm0BxsmAXF/rmThnh/pwBqdQ1BmLUhkifTKyz
vgQ0UUWbMk6kF6TvWcek2BevQpzWOWIRgZDnLmtcEGf91DuiMzl2SmvK0ctv
VqPsA7U4CoAeG2gr4ne7QnCUIG7rPQ7KbOSBZtWpHNairtkrJ6ZzB4lSiheU
HA3dyC9/3yZuNVzciM606IQPb+OWyJPe73qAOOqMHRtCQIZ5REf7Uefn2lmX
skoFpYy3uNzIgMMMU2Rhqq0nYLLevBBUReKP1xLaw2C3vSjlka3mhbeV+gGl
fMyxPTX92SITlQpxE32eYubFYyM5cx8GyNLQYOjzClRjQyOMt+4pnbYxgFP2
DRTKAfbSoVS6JWt9ZYXtQ8xT3vrFH0BRmsQB9y4wRRFsI9eNQYskBb6GI/1j
QoWlf+nkv8aBI0QvekqXrFWqvfNsusc0F7ODsYLI+4tcxfBsqFaowctpkXM3
8VLpdGbMncpR58khKFmkwBMByDKLlgsCCXuCwugLAkhVxqG5VeMMQFCsKEM2
OnFbUxQDQ6Lt6mHb+JUmuAEtP2rzCE6bXQnREREWvs+tRMEQZMw9JlSeOTAq
eLRHqZLpHwe40MlXcKBj7WrF3gAPa5K95jTHDrXZh4b61iqSWkYt9DsOk6/E
3jaam2YpAdsK7isgCWR7Z9W82KVRebQOs7oPsKeW/RZt99dwAaShux61HnRq
Baq8XsLQmpJJOOIxOdwXEzGRYB1cZzb18xbGRWbnNAWGlZDGE7kkOda+UMfS
pzaGb7Bt6mry9BNykjVxH9sn3U4TPKPPKunrS1TfT3HGKiVTlEWR7Fy2iqmD
X7xz18vRhysCfJwfh9iXdz9Kh1pvBOuw1FKrDRqgTdbHlOL7jTyBQLLsrJ/8
pBd3+e/YF+THKf9sGzHi+O+2j7VFkmfnMY0K44nYPSm9cb5LgOXmOHO0bvRU
pFz15QdFd+A1G6Nk+XQ5IdqLpq+OQ3m1QxLrKDMbpUas3sjFJR/bAUWUoOjo
MRVb643i9f1KyQ2PFmHCG1TDfYhajh2EDRlr+BR/YrUPTtVDzrlF/gpXijaF
mXJDt/LKKZQSzsFkQdaidGWQZDjM9i8aesNgvpU2cXrfPUBgDC76ndY45mOG
m5R6y/82U/M2Q+Tz3mMvOxjNJydsXr3ME79Z+UNEy2lPLLezjVyXa6519Fjh
9Q7I0H6hOpWUsWdFPPY4T/q4ZNSoNxN37EU7CmXf+mM7gPRbP/aMh4FniOUp
Wlg82IdqHv8Dj4gAgBm3NM61ERLsgJ4phATBkPhLR3ZsXbSTf/5/FnjN0woE
awColywLzMLfWq4ODWtofkoA851mXGTTz70jByrBjB23g2f/VLTJcmugAyE/
cYCiLsxjmJZbAmJT+Xb2Xaqx0sdRrBfKbcxzV+2umKSrhIp0vDhQrFdPA0eo
ArN0925QP2tE2bipbnP1eM6cAGL5lMyhfmK/bSx3WwQc8NDbl+R9LBiBYpUd
Ckn3Dl73itxNJePaw/3h/X35/nupEHxyKJjy24vvC9mMVCfmzMqV+8BobVvL
iOnsQ4eLckmEPnE6HQYXLKp1QkDJSsG074kb1Ow5XeaUMM0viSmn353pycyU
fjAqonqApCVGt38aHAqbpB8kdftJBD1LaKWYwfj6Ozjd2w5tpB7IWEV+PSGC
DjxR8GW578nFq1PantZPvUM/3rSuzBicfYTfaR2LL0s3tc4ceABY/MDxYx+B
7ml9JHUxp4gq9Z2cKaXBHKIaZHJylySnR9aPjcn4S6snPuM4UoHpcuqps0gO
2reeR2qyvEH6ILepqWf5JMJo98+YNMMqh6KpxdXHAddtdO18TaU5v9jWUKfA
KYznqYO6z4C7PCyxu10DJO9M5DzijaabXPl1skHZX5DVOmMrSfNMYN8iYuLx
5p+YC8chBHn3uqYl7lV8wAhAe5e+EX/awrhcSSes9UW1IHhu0oI4yY8PaIJC
cWITLOKgPqUDcMc1XDiPW/xECI3LKgXkFB+mfQvNjzgrXA1RG6YmcemEjLQ/
0ENKEJ5W33xipRR6ogJk1s/O9nDIcjQ/D1d4slpH42GPlvKnyXMS/w4iTjds
EjDwhMc6vukTlgld0SW0q5rvjMnUIImKq0Cq6jD3KENmDesNmgWtSfzfO2z5
/dCoWUoSE2pveGFDadwJhpc1pyRRacckkCpkk4UnhOTnoe0dJ/gk7gPNz44q
bvdPkQ5CjEk8zuroeTdDnvMTfuhoO64/TmgK1Lp8ZyXh106qjN1cd65mB3oH
dFz+QQMmYQ5k0DqZrLaubrUY5eKL4xD83WRVtX/FFVNw7IousSJI2tx3vcWT
GM5tcL6jAlecbPePQ1HPdhBXHKzNT4+s3+0yEjfv2GhMc7UpU92ZxRjm+5KT
KLzQ9Pk0fs3xMb72FS/NQ7C6ywuM8PzsMr4KgEJ5dhrmz+Ekl+AuN6B3SV7r
FLNQP1mrROJO17dwE1Esd7J9WiTdi8wcK5cVy0iDx0yaOZOujyZX7bZZsy9O
k7eCj+y/5xxjtfPebbEM5axS3ilYWs37f0vnkVubcxG1ML0CEn2wXr9C/34e
xrp3yVx+aNY6v4H8KJbEuPxuGM2l/uH0RVEoV/9ik9gcO2X4fJuMD3fJFI7g
vkG01G8W3cymsM9aXES48h8pLU6uLzQrpY/4NDQjPUi9Iz/al7fR9mTciNu4
Jho8xe/WQUH1s8YHg5qrSfMeSvtXwk3okVyawfvWY9G/s1+TPu5EVTTluyW7
8En8PUZmjI4KfFTPPL+mG46JBflVsY4McNtTpVYHqNq32DptZl72NbkvBQn+
cp3MVZ0XSBtc3c7TzFAm560jBYU/SZxuayhJsAS6Y01xlvCpuixpuuiTcjsi
lQyivAguXkcrIUctrFvcrlf9bg+OsmbKDuI4P8mZsrKdJK3ze+OANYBDBRJJ
5xHiOFrEuYXirLElLOi0C0mPDBee16sQie5K9FDk+XLf6DTc5Y3ovE5B1kQy
U21LJfK6XR30bTKXTyrv6RtGBDLP+oiIE0/35C18GZuaA+WKPspvwSdXzvCr
8ZqQ5RodsBarjewdF5+qDyW0hhMr8DOuSCPsWbsXqEuFRR6kReCLYzs7pshH
pr122FsBughXGtz/V5rGSqae3Q7VwMUutKv4Oh7YnB4RcRzmjGDY2ClTLd83
uxSL41oDczbZNLopcBKvGF5bBQtQHzwpwvQmIruuuRKDO/vEWZmUNHbRWFVN
wWvC00iOz/6gb0zMuDrCNXnV3gBAfAUtEHvLszlvR754GVR2YzDac9pcjNR3
1Z7MZRZE3b1+pOZPUXyBzRDULeeefMThylA2Y2XbXliGnWgD3chUcVQYdwq7
vNd3BXcOGmfkC+2dqzcQlY1gBkZ5LxjgRryYAud5TNchy2O/LpF7PE3qh9eE
OG8Pl38eZz5R8i1jP9jPHBdVZTziLA27AZYIyiF3xu8aONyty7vdRyMYPqtA
14lLxuOPiELkDZGpyP+8iT+wCfwPtXlwCy+EyQs1AltPjigTPE0OaybW2vRU
+6Tmx6kuHbPsAZWJYYWR8eA4pkQQqohCC8PlrzIqHqx9GVPrLwkrJjIW4FVg
8Z3Gm+K0ZRBZhH5OFyEGJvtRNLFWqugUaljRKBun7qj9sXSovl3GqRbOJoum
mkQyBI/xyUi91w0ODZpUfmTMetp1FMWhCg1QTZP//NwzrtrXPfCTNS4+WTM/
z/dF68eoOq6aOoGEYbRDVM4MMH30kfblygdaEmf/+RqU/aLTHBUH3q7MZTMm
itO0eLJrQU993OP9CVCrBu/W8Hc7yz5Z2bXJpxky3JxvRVtNNfwqFCmDExYO
EiIU9tMlEmo77lGN45fGQ3SG8vVoJv1FddAY0MZg2dBjd6LnVSoxf5YhNHJj
9DpiCS9E4ygbwhiriwZIAmBXMe8h1V+TBJEZtwNHAw2SF4mcx+fXe6foiCQC
V+0ol0/QhBU8KsMXZ+VlmvlB0bibjHC30DU1WfitkNYljG2ZuaBGKzZqRhsT
uCQJGCCF32fOyVfcaViQ5ca8WdMiibrTbR1o3O5jVsLQqo6kGNBtFSjJgwsa
A/vHHe/osS5av87o+UHsumZXk5/vVwFoI79eg1W1dT5QUQw6UhQJ5XIZQ6F5
DrYSCz+9MbtjvDySBXMGW9S2oX/y1b/gIzT2LcLvJiEcK5oz73X8B/eLiTJx
P6MsRsc8Jpu0dQliInFyWqpeA1TAyzPtGJILjyVGY0eTzENgJhKo4yqtpZwu
HaEFZyrTCm3ARYf6LcDAmDM6P+bn2khKkeVd5Gox+jAkFn15Pg8p9nRCutYw
viS1T39dNaEAvoCAc0yvEknZGy2bdPNwHhVObWdmpFfNJovSoFs8QVQ1aJrV
W4y7RYyJBb+plht8AMJX0JY7vr6kH1axk6QMqwqgvkOpoCSDM8o7ZSpGpTuA
4yUMWq07t8/5uOnJtnVzwJ7Wn+H+wWNdUiRFImTiKyWZAIi+LYdMOt9ysOva
OXryFLxMbp5f+Obu+OtgIccN7E60CpYh6fnt64rjz1/SGJJ8+1S7BjJxKwbi
25qwqaZl7Yw5ck/pZ9fbo/a26zl4vjomH8r1yPnKy9BMjUsF+51wzM2nRFaq
8mPNGCzrnN8oa+GkAuKQvAGDTgigrInwDIg4xbcbyENwcsyVNRYzg537Wr53
Yqf+qlfR9Er55nLOPWjDs5vmmsedwgzwrmE6fLUdLzkvKqM+kTS/ulLZ5Sfb
dU956CjS+gDth1NtbmfKB2vaG4UIvbIWtzzCd4D3s2lSLvi4H6eGrnufH4/j
LtublD5XtEWkl0/x65+TWFXSFkyG3wz5I4BAO0hfv1GJd3AbSWm8e8rcCFxv
p+NCxa7SQoLjkp0FkfVuboOVqRdX4R8ocDK8RbBKwV1u5lU6kQ7jLXBO6nsP
bDqznQVaofvwJmiQNzSNc9f2mEHav2g1kvJXgBi1qM6KdAJRO6LswAgEHjIx
OIzfCUU7PsWJ4/8HUXt+SVpRHdu0vsUX9jMswDZ//BjE59EFc6xUD7aeCCrm
ms/ND0xJMaairIFvsa1gMSS0O4N/jUnpHuqujJ2eUA3SGpFaO7gZON/AGm/2
cNV4/SJvDoh2eUGLSFRus0AnPTEj15LqD+CZNqdVhmsl92MQGjQGxaEp6RI0
CGTM7EoIhPQ1YcOoP1yY60vKK+6qKWJJekQEu2vW4qayG1NH0sV2EbHMKuP8
2QoX0yQYaPWlwZBS/apfI+yWNWSR8CpQkrGvJ0NDOkhApWsSWxlpFpV+bKNX
hmpYBkBetzWgQGPp+ZIC3LUvZ5YDx9FPOp5pHNyVlHe8W2EsUTIAASJ4Nwfj
hOpoVQrOqqGskWgR5KEItm4pvCBvAlReSQelnwKCZ5P4vao8oxtCYw0fxA7X
mogREfBOEGzpDS5mke2DguyLhboKZck7xSl/vZu2Atgndq0pw9ArqTJv+osT
M9SQ0SPZaMaycLVB9NoMfO4A/gnlgi+E/pinNvczpn4l1h/XwVqqIhBt9Yvx
/x7Z5pc7uk5PcAI3T7qPXMk7mMq7sfYRDnwJGfOjS38nrgK3zX+hBxfHfHLh
YqxLj6JtTwLCiHAgt0jj8i/JBe0vIaUG35/HQ31jxg0s891lrc71FbB0XlvB
PLRfkIt2DCjj6l07p+nRslBtMfwH/ygpAkBMv7b21xoL3f3x9Tt+OqOQspY8
8V3d9CD/JjTZJTeFvhAeBtBa+Kj8l6KwOf5afEzgSg6Wg/dQQiJVU7jPBwl/
k94Nw7FNT+EL6X1MgmYi4QEzLnL4WPisO8YbLGo/ihkp07YL91h/wlJF8Qks
kDR0dWwfmJMl9gVmpnUYnevZnmzxmn6SQCqgVQkbYRaliUzHsrVmVLARQzb8
U4KKJ/bz0vi11IiQgqUGSbnzKktfvhgIoxSz4OEaqEvoi0cJoJ2Towcz6COB
JnRA+FxxmPzIWc+A8C/nCFURDG/A2EnNKCrRB/KlqfSOIYEjD7kS+zCtCL+P
dU+vxu1iZRFu4z9gZSU/oqhVkhOQXOj6miOhqQQb6WwqkAh1rwrsjl4BeQCh
Vl2i/26n+PeQDHpOn1dMhBQN/dRA5edXJWj8pbxCCQczGRV9UraVi891RD+t
4B5aTQA4bCoy9GxrDoWmQt+52JI2jooScXzo2KVWSNMZNZh3+DppTM8+QBFG
zp91N46ziWvmKkFBGMW/3Ruw6AZgA+n8+gXgUsCJvR1Dx7K0qslCch+9rDzq
ZfDASdviHSRSb1oJt8j6DrV0u3shbsisd++BdhcRx0n5Eji2f4lgsB1fxpan
8ReoEeg1UtrGgMX7a9jQVujopC1qg0RZl8i/Ys7ZrQiA/Yx3esUV+5yZxfP9
bDSbsWJz5ai8UoTY7RWUr/ytbBLJgqAZITcNpudRrkmK1t+dRAGVyAeY4Gwc
V6LF7TE4VOUgj6zwKWVTpYi7lSRspi+SXT+L4QZH66/WuWOncxOZHhlGBmdR
gC98NhEdh6p4VMg/aqvPSkJlGyCmR1M+cYGnmg46ySIng1VTHwmCsGnRlYEK
/qbHREt2lrXvfutcQVAsy9i1h/yPpJRwEef2brod73hFW/vrmCKLcIcvzBmN
mTIK68Wtp1Qb1Vwx9wJQAhDZp9cMlLym3AYsQERfF+hnfHytdjyt6UjjTVSL
eKhUeydmbYXA0AN84UtyULKjtGBvhOsdnaywalK4cEKbi0+Dbn95QKvREnqp
vuvNvAu2dPjRhxdJJ5AGILKmCiQerX0daYbpezmPl9674re0pMezcIurUcvd
D4JPR2RkE9DedR/9xdhC9A2PXd1zpDFvHAWDwNZbRThiMQKOBdxFLZUvca41
MOM+96+JjQu9/UHbrnXUcjOM1RtUPcrZH2Gcb5+zHr5eeB4pWrHAxoaBuun4
txJ9sjQt/3B+HOhMi7385bfWQYyaZc2tVEP3nJ1xxgzOxSzy4742rTDxbbWK
c8rDr2JjWsM7ObUWR9FOTvUOKn3CY+dz5oD/SC4guXy+l1kfvlS5z4LD3GNZ
LEj3e3oWTSnWsi3nlc5ROwK1bujlDV2L1tx73T7xUOosUmLprLjSyKykZs2i
Vv+vhi3N1pteIslAAzELQkHgCg0WRIL6+NDLTl6R/p/cusNChYSQMGzzO9tW
QsysjNkU4xHz/xSswdOOpW0rogmDYGbZiYZsLjJax6aNJtkRK6BjxPrniWCA
08cbIJrFQrrB4cokNez3D5whZJ42f1xwQlGZ66p/kP22+NoM20L6g75aiiuQ
R8ltbviVb04xO/CJlQ8D3lgtFHUg7ysuOgSyOtKAt7ToZniREaANWaXCO4o2
z9jf0y3J1PLQjs5cn3gGPL/5mpasfo+8Jd+FE0r5DCRO9jDHKOXr/xO/vna5
TfkJ59gPlTYzD5lQZC1jsh0ppmKiazI/NDlobHgBYdhadfVCwLZWVimI7Yga
kLXEjtS5EnRL0JBN7eMra79xWGeAH1zgkTzpd1eXlTpHJVFD7LwkWZWq/zKg
Dl8GBV7+Ga1uUPZ/VzLJEfsdZ+dnKp1PeJJPCflrTCQzFBK8/nCi0cCNe8VS
6Ag2+S3Sj2sKZktIkbueQ0Ymg9I1a8MeGkIw9YDFgQ96wAq0pmN8vVD/0TWv
sUMGDKBi4GwHc9HozYPENqoERz5nlLd/lS2fhGxFfAIIJL+83CS+DYOAQOiW
z4cwDhsmK0f/dHysxEdEHO/K2t9YIkQOyQCXHNCYUxODzePLm/dxrMkespi1
LnFfT2WXKHeKEHxo9m+FzrM7Bi96G3foN8NYqjkC2C+/KhNQEGBMhhuMxvUY
2q1BMKk+M75Y7ybcdiY34oLsgn/xQHD5/dU83G0sZaX4m42Mi/D63olhDDq8
hVws6fjzG7V3QC3vrKfvAbVDhyL/Y7FZyMy+UyQPN1jB93VwoErVCX/GYLCE
Z4UZdFuinn97dXsoD9891TaAEasEWCA2hDWS7NLhw2P2/wvBhWmn8MNfwArH
MU2bSqO1pV/oNLLAxsvokyj4TFgDuWRY0MaJex4kWY+IgRwU1UrFyL3ms5I6
FpjRS7NZMpX5zC4XPq98GelfriqM5JoqzJFO5qGV+uK94I1W6dNnpSjNU6zI
6iTx24186Y5APPYRyj8p/0r+YZCCWJ6OEcO21lMDRjjj617Y6uCP7EQa0rAq
MWCus6ocMkyB6Kh70O223CPCrYaumb5pzYgZZKB2K4P4j5U/rMclv2u7dqWM
ax814Z+k2A2NZUOS31d8luL3lD9v4v0KUofLixvpoXsJtnKlb6yGkUfyKB3h
TAFoDeTfPWHbRqJT3dPRTha1GdUQ/Ar5nHf9hGRIxMu7CYVHuBImRPcEPkA5
CtB8IbMuhbgZgUFcGz6mlqpGn1jGmSuy6OfJVv04mnt35KJ2SCOYAdKZQArI
R9BNLz1ViqH+xjFmjYoS7ogAB0hJanwFdos1x/6aDPjXHfcLYeiEcs9R4PNd
WbYVRoQrl9squGJ04Aob4bXiC4oZ4KDARzn71HMENWjEXapkSZHaHH+Owsl7
iE1X0jVTZFZHV3EzIQUbar2/KN6VogNobydfOmWio9sZNGPeTZbwfdbLwmTk
n2Z4RkV9rteNie3T5nMassgEjsZqyMyHgVGZy52G1hxdZwvMGHonQaUeshP1
42Yb8EOzFWvE1q0rdmkpEd08/zqLrEX/2bd+AqRcuKIcgy4EwTeF2ZqAWreu
zFYJtI2KUrQuNFVHNGVlMJoQM5CKHl4VPeMGlVYhxlwQyqQKDm7RrUEggEVu
iUEU9VcU2BvAj/oTL7lhKek40B8tgUfTt+AQ/IFCB3lUB1X7thQT38nUz88/
Okx9/9jZHbjVTVJAPq/8eu+GSR2DSYDvLGr4K31Cyy/8jAxKjhP8YXB1vDyL
FCom6B/X/RMjx8n199AGH4Ci+Bo8R10i+TH/zy32hybIVpXUJziQbCU50eYC
nEtYM78qayO5/TaE/OOy49DU/uxfU3bKtQxCjNGL5+VS254gtAzvDfkdR5oY
o32ZfPYQZrbrtqJ/86ZxP/SpuT7mk/K/ZIaEmC8lEbY56Ub7Cdv7pGd13T/F
+icHGITbAw9G56NeOMMbZ+0s07pVUdpvTOkA0m1kp+2Nn6Vm6u2nKJrIQEvK
Kb7JSlP6BU+CdL5HfOIKY+M52anzP2sNF7wHFoSzShI1ZWFeb4Mwefd6dp3M
Id58rFC9w6sQZxqab0vlcz/x3bVOE2hacQS8OMXyy09GokN1A0l8Sc/+SwAo
5Y5bIkEBJsxZEWZ4cV16CTafw8Mm28ZmfsRxnYP9gcRzKX/Gvsnav9I5YHUd
82WptklQsNUWK703itgT72KhRMP9edscGBoDVk9JFx2VSyHSexPcVrmc2qN5
JLdCDs8kjJ30nIGKF1mQy4EsEMj96U/FjvOe86oJAcT2eyAtoqZIgFaq5HuU
2dZtrRJ9rAgvMtqP1RmxRmZX4bPC4lFIr+kF28SsJNgS4kpoSEYCIuGl+7v5
HPLMMML0rMV57gbKLgIuHSPC6K2jObpXwk4Beie5yK7kME994tj+YYSir/ER
FPPqSttbFZKdDfLQ1lDIIRhS0hlMZnPiAuINsxb7wDVb7DbjCfEKNE452M4D
EWwozesyJDcyaAf4uTb9eRJTFBj+0QACp6wltelVZQTrluah5KzWdR6FjriK
UOmqH7oK16ux2y5w4OdYJ0iwRAcQunAtdNkk5wXCaR5iqFDx1d0pwe5TovbZ
aOjmZH7n0OtdPHCWlwubveME/DVbbj7KBmjtyGFvAAa3bzVyOZbaUTaYYn3g
X5OhTJMG40ZJ6KJLKi1OyDrKuLObvg2BARXWDjebERFFKV4K9zFbPKFqNyZQ
GH+Kf6iXz/hJwYFzz/DlHDp8WfGBZE516j3Gw2QQiFWaYEdojTZpE+1DFiYl
v02kXUP8wOnDuHfHf5Mfwszdngzqs82Ss+12GFCXURVNYFfq6EgShxFmdAKf
RSanYMGwe417UGzVl7RWqCu2FyzdeygyM+FOFhw96SSGCiLx2+p5TYSx916K
znNXrfJ+KGk2oSiZvFOmPnlr7a9ghuD+hAD2bSn4RcD5AiMBQitjkzYfkDp5
/REtEWpLScckl9TYrJ4Tglhr+exepjSVYDlmiS6/rh4JKrvTTOJ0vRJaRItX
Vs+JC0JLkuh+ODpp8KxEXLlUpKrWwGOx3ECZlujfQ2f2J0l1/2gbFI5xrrlM
PvNeJiX3FV03i1IUxUwULl1jh0Faeplxx8/eC0rhzBv/VoCSFOpQptoOI44L
eqGQbMiCEdUQWbeTT26aa8hgJyWQGhYG/OubBRWHDIrHGniCPDjuD7U3n5Yq
QaOt0on4VSo/X86D78wn0ugRU8gmGHwcDBT1AAUHofMJ1WAlg78vnKY3iupu
0FpmJJVinr/LNZDRnPir+UnQFWAvbZHkxhOclhudm16Wx72wM/sIcQTjTolf
bOqCu+hkH4e+t972dTQMp4xsX+uu3LNcdWM+8r4XZJz1s5AaxNYf7HV0YRd+
AncBWyay+cdihMsrkSVXqTvCaea4KrcYSTFED6Y3xHU1NJQREFsFvJSXtDjm
LchlvAtUboaChGc6yzzBVEUnwj80sH2L8YFEFDFd/2vccsm8a5tA8qREQMu1
54CI/htqI5eOB/owZLJYWNVZnso2yAhTuk2mDd8V7S5atOO5I3O5nZ8jV2r9
3bZ/AK7UYzwKVDTbhspx0X1xf3uPFYuzny7U5S0Ss3waNW0Ei65W+YeZfrD5
ES8R3CrDVmH0A0/poNeAwyoHAaj4Ifxi5Xp1/Z9OXuXGnUd6CC0BRX6YgfbU
G3dX3Ctt1LpYYofc4dH6grejNAI2twnMjhG23HUwE7Db09NoiK+5M0qvWu2e
5vkYMjwUhUF9yG8JrPYNyGL/Wd6iO+tgv6awhxmOkjPOWbkGDilCjRkghp/N
WIVkeoX9NeyeWlCmlPdy+L6/hL3m8SgrFZ91npcUcd6Bw6R3HFAycoeQ1gzX
uu9PhZeBCqqXKQ2WK1xY0ZVoK9DL48mGDy0VyjLykmziyTgkTcua6iPrFq+5
6f8XUf24ZRpdPW2tuUR7PAJxGOf43zT5oi2tUn6fsjxoNiX+DxYm9O9x/jbW
KBIDU2mNKOldQWuqw0j/xuxfMGUBevcm/z291OgeiGB18VU+Jb9n55uZBre9
NvLlH61c6Vn5jdN9mqSB6XLEDgcFZGrnLxAfHYnYbIszwdmwOp/AmYAd+GX6
0h7z9kx9U/xZlSVzZ803ItuPQsXrVngyonCUDiGADCQkzleMTDFcf7xDw0UU
N63ta7Sp9ez+2VqHZdkOM+k49iR6fIWFOBAy+XmiPmiu6AyfFZqTsZ/iN5cJ
xInHsASFCLbMAYHZn9iHqWU7Ue5KXDMQG/j2f4Fwcy+2BrrM/AfjIIkqEqu6
TtE+T+cYT/9LphB5tX+Dc00fpRc+4ZivCWCAWKE3evgms2/HKgAPFROWJ4eM
IpAckuSL2SxBKP/tqFvQvB65Q/OANgylf0LQqjTMQq0rKS6vupny1+D+KUVl
t31io3DJ58htSOIbmQAdx5EItnQcNHjtcg2Ypwl1t6EiCNfGdFk8D/eGAbSS
w7L8NN3+nj3CNOQgMM9IMc0967UNsekfXnSiGEN3/EaXAbX3sqLz+aKqQRt1
AZ6RFc3xG8maBtTj7gGdkV6UDTOuBqfEagufQew2E3jr4JMkyeLzrnpBIVBe
mB9ifoNkRauI84AtxfLreicgmp+Khc3n72z3TMw/6OqQ5XDRXAbuvCttsyXa
2R5SF8E6XIQoair5jv0utZZui4fGLn2zuyjapeExkizgiAr32Jh6r4Q0LchF
ehE6fAaUR/UJEy+2jQQN+U5y6mIYjXSP7xmUzLRah5WeV6Dl+BiBhP2Z9zH8
DU1yProETa/NITOyUC22KkM56K8Db/uqxVg2G6ZAve8kSPyX/4C6AwdK1nWw
rsAd6nHum+G5XhXolVzOHzUWVzkdLnfzjn46TCl7pvH8xx+DaRnJju02m5Qg
nWxB+Lbccpwoj9tgyfhSlinDg5FiqzvTGw4hZwKLNy8VFFn+fG2h6bOsnWco
B5ubGXbwxG4PxoIXwWnElZiCYCDM/5KgqI3Qo3XbeyhaS56tkDgaaU8ThncG
821kD9GeBIQq1Ofd90jqaP5ldzaOvrvltIeng3vyzXDzXzUmQZd9ohknTjbX
3ybq3PmyNaMnUAzypL7QdVNrhTKnWjaKc2MqoSUzPkvykAZj/5TljTUI+QCn
V7JqGe3AFeRzolyUU98CG8pEoqvpuh6CMJWSdII1fEdrOVafOLLySOWSnPGE
Wr0U2i2vp352XIN4kocQIJuJ5zdCZ3TcOE3+AKQPybRpNnwJbUEbL1Ev4kmr
7U06nsSkiEuwcMoMj1ryGQeAQe5adnOvshJv3x/OdZimYF6H4dqju6Z8wdQ/
fbOser1bxjxvdweUukEsAu/LhfYd2Go6L26MnrgW3fmSaOYdhjFXgpvQixZJ
g1hmAr9q8PO6QDobk6uP/ULXc4lUy3cZOqqeSxyLX7HurnwK+AfaqniTtz7M
UZd/t95yp2M6ieeBejhJR2/2XYtH1KNky3WBpuVze1SpNpfirRQI5TlvQb8M
y1pGpVwki7P7tErbEQnX+fnLsN5FaqTU8JFuXe6zGXOElPiJy4DLJU4j/BxE
R99fThvGfeSiOrNvnPCP6CqEHTWQQmqX7NH2Kb0Dml2O865ijNx/zD9emAis
TMipeEh+ZY4l1bkryyw9+/OpJeDxK2TcyVu6i/WV3inld/6wFYtPgnZgMwLt
RF44ggBlh+FLzvcu6NwsHBcGb4wUXrIzOL8LFeea6X2IhxhS/sCde4p1Vr10
k0K1EYAuR9Bztz5QcLn4St9aN27Ynan/Pgk/0q1pDO5LTZwl/ifK3oKTXwyu
eiI1XU2iQBjIOiJUyGnR5KTEDSjOB9O7hc0BPbbfmnHeD3Q3Iqi31HztNY6S
sVIdOkuNa6/wsDug2hxfndVFDDzmQ5ODtR0PQyJ6m16ID6iJVNZn9P+mZSuq
3lemwLal3Tut2j1d3eaUWS/xdxwy7FuTaJp/P+GlD+ChiGgr7tFhDE1voSFm
JN7A5XvZAhkeLZjR6VdWgyTUAb/Ky/SeCa8LccJbZ1HnkiSo8OAglOvyippF
ZcLaY0oJFKtvMrzjTRLa5rUfeoB1v9PB8HP+Z5PrXwUctS55qDb/TPExxtHg
JOgZhynE5xj6kOM02NS6SuqmancXSM+HFsNAs4oyv60GkEoiRYHnDFMEYXhB
RQSM0DZIkfT/ev2gHNz7/kxAo6NYtc5DJMsKP9b8V97iMQocr+6BfCTXb/Vk
sswPivfX+cHilUgGM0ubW6Rq/r/trDlqH1T8b4tU0OnA4gzOmCE7csg69x1V
n8JsmiGIlxX7lRxzx2EH13WLpAENP3aU/u/L48SvIWI+QEMHR4GbNUV2vcH8
LuhX6EKhCCZXX/pqtDjI5Mm0TTUhk2S+ro2wv4cCnR28kBTp0PL6+NhaI+/D
oKfvRjClrIE+jRgb99S+XwZDWAdbXMOTVRNJXS2CpnGYn9Z2SDHW9JvvLRCn
o45GLY894MfEw4A6QzVDOQkHXpzs99yvMhLLfBptbLs/nwLRpVU7MEGekxUP
+nLx/lduKrEOOT3tsSS/VOt37SU0stkIFIm+Gzlw26j3f9VxRcfAqCzE9PM0
qHcn7wV4QP5yvhZbcnm0mL1XG3yzFJwjW8yIa+KtRTxNYW79+jbRkbjcZVBB
0I1XUa22lOSE+w/DSJFZZLHeZF+zLpsgPoZBKgUvU+zb3jI+fwacAMFUK8Qj
ksyMPklzl2ChxqJO76tfiFsFNEF0JrC1OvFezOexH1HRq7o+PBZg8ne0I7Cu
2gBjJ0BKkhUglp7eAtwdtPFuW+8AmcrXflXzlBmSNcJk9USlvOCoJUPK0jAZ
UA0U7Rn0/gGzbp0GYugjHrQycDeMSm9KYkw9J2FTLNmSVwrTOm/t/CGlZFeU
TN/m773awgQW+ppiB73JsVzrCFLyex2aeMaEsEvctQSEUmZk3BlLaRsK8Sm8
JZ7U9e5hCw7NMy1clTdwq04bC7izQ+3LK3bP7pR3A/QuPQ+JqHC/rCiKMib0
4PrLS/ZxNphKdzzGKp6VK7MjRtNaMJs91MnlaCn6Odq1Izetb33Iy2gV9R8r
yxHAFoLyXVs0NQmH24VRp52R1mF2UPETKTc4FbLq4yoKiEvXroPpgxFIKF+2
1OOirKw5szdnGbxo99l5RF+3Es3U/wfUKpB7LS0O7wE9mOc7DYVGvKza5TjA
pZmn/nbZodgE7Z+8wcoFaFSYzEg5AADxH4Icy0z8d8BLkOIWAbus+E99aiFF
+TyCg7D2nZ0IBunLBOw4qCpB6DvE3e8L92YXefFcqLrzv7ftq9NH0jqXVmPU
e7eIoneYo+AFjabOnXzvvr0DA5IP5+dpRTU8rYEjzf+9kFOtdgwbrse5nBhM
QJBM/t74/tXcY6pfFUa4ZrNucQ4twIJDB5fnZyGeHSffU5hf7LSUuMlBr5V4
ALuQz7Zkwf3xCKeYcs0FH5L3fI7citFo0kjpDv4B1A/MCNnluQUTpCwoGXwn
OmKcaI/JNy5iJ8rATN+cRMmnTRN5lfHfW/rtqcs57xGYmsJXCKIMPJOAp5p5
yikQA8OtIZw9UP/j+ERUus6vWic5hE3Up0/1RmTnG8DkmbwmmS3jvqVUZ4+O
G8vKclexYCtTRGcTmMPGuSmCF1VoAOox8MULHEqqsFX79B0e8s7Xnymh3reF
eM6JMjll+7N1gtmmz6roLwfPylxVIDcNh28XPWYBsDciRUrO++nWDcVzM7tV
DgYUDzx1ESE8P/h1oci3rNuxI6Uye+PdsKwWUHfRXiRsUneA5CG/f6yXkCcN
CKgU9vjoKlkVrBpf6uJpk6MfgZkD34B4gY/yW7O9DoMuanliEoNgDCYhxpTV
pBy0FNxGMj9sBMZsCrUSMTx2bkG9Ph4KpCoDB8+goPPnfT6CfJSXoKEoKsLZ
8tBz3wRIHTdeSovmsFIIFXwaeVKrTyedzDdHL12nTPbBnGOIAQMlvU4YhdiW
0mNnqEuNrhMUEUnCK8LHhRGaxVcIEGbus4KJt2kZqIHR6P83M5hCjfa3CFKk
7LWMw4nFtBR9oP7O0H29uSG0mf2XMcQdf//B5EMUwBMat3m9gF33n1+KdnXy
/nqLfYPznmsKPqT778Jm6cgXY9SxMIM7dy8PWWaLFqY3OZmOt5Yu5e/W1CU9
n3qvJ1yHArZ9CCEi+7z0l91oXOp1KAl6OWCKBxAd2scxc80BkWd074ZtokMy
CY2zL2ebkdODtJYXRtKZX3DFnBIPKBEdImhkvV/zVA7jPv+PZ2/xeLmMjqtM
nrtsmI9niH9ENmwBd/W9t9QrLDuHI5/WpgsG7wxOl4M9Kov2riJKjUpo34oh
FuU3GUaScSFv/VoAR+3IptR7Jh4C+DqZLGYvTK9FwJjYxbZXJCfCj3nePzk0
ODCYdRKuRRI8XIJ2BSG5qOyNtqH8mvSCFmLesLSOP2PuJKKCXvBTleyw5WZr
BhgewrcRJs95G8sZpW5L7qTZsyGDCNs/9bzqDHg+AK5Gy1kbLXwXCb0b8QCP
Zdfe8k/CUclFF5ICQ5q6eHijfZmuNyGgJ/ALZ9jUvQv3GC2uUbK/YLTSS1Yb
ekmDnYCrv7B4S5YQwINnqJw73+X3wFpJbRVhw6WbVaHXC1wcCLbvwa3OrT87
/Q0txuL0NrjQzWPupXkjko91AQMvQBy/XDfc8Q+UjmrKOl8RVMIrYt3v7gov
E4VaHaY0eriGXZsswEBke6kMueACN7/wejnEpieTXu7KgRi+B44CQjKKtAXP
dGwWkEzuuRSanvr0a0mbCuxuQXoZVQ4mqYW3jwCoM6VLJISuOBF712KHX9XQ
RsF60B42uUiGl+SBPgUZWoNktNOi07cbxKRE1QvkPMIcjJalkYU4pnnij+3P
T7JbVC5wjwuOkrhkEHiRGK6b0bZQd4k7GnkHcCOSiYUmEnVuL+ExjeFpmbwa
IU38nHt35Mwe7FcDzEu4HqzrErFOu40WQK+oHw63AnUalcK0RmIqdccfiyMU
c0d+smuYMJLubt+IXMPpajKIj1YOPtcFjEFpjVqaRuWgWKkntD67FAnGQEgY
z37/reTKWu5l+22RCo913T4ZSlWWq3KZo09q2GMWwv9BfxTJxu2N9kJBRt/3
nVWyK8UWcZ2rrO2kQE/e9RfvnUau6pdAm287K8IOuZLEeZsA5fhGk0T1Cvo2
jjzGAdfXXpWIei1sZhp6CDvbTqsIsVgvtaZfJCjetjwAbIzEw2X1Nc2aHPSd
mtS261KweV1WIf99FOCJegvs5X/lEU5Mpmg7AJF3J/DVopT95fHolDXqn9Nm
qNwPbLGW9oR0vn0jgaXV7E+sQwmwZDtCR3bHlLir0aNWvBoY7jS9lF7NXcjW
JMDTass54tkoYUiQEROlo+9e++g1SIDgoQhCLt4wggPoAVAuR4ty7Xh6QIfu
t91+4ak0UK+TMcfyREzsc5r/m5dzaOy19f0VbL/7l9N+5y2Ma8I5qsj4fMnq
I/YxG/zSokUc6SSEDDiUr0L5zozFtqrZ9H6hzjRpv425f+unVt7hG3ZOug7s
xaCwTonpQhVVxnBaMyqY1Axoo0xpiyfrD1uEVuiGpRAmV7R88KwFiHHlN8CN
ypZOm7OWJG+FSt0NTRKlUU5e0VOe04IxH8Ymw7X+mo4R1/vxjSJpCd08qY6m
U9wjGm0go/PSvaKR/6vFQBC+momyyQEVCA4YvBGNgcq6s11ji5zmlOWjq2k8
wks5htWmVyAdJP/58x4sezsoH2F/NaUdl7a9Ckt7mndVjvJDj9A4RczupvRN
pxCa/GvtOcAHVZuTUCQREBzu8jC6ajb2Cj6zMYo1ONQva30QMEfKjPzOmZ+0
KuJuUqePcn6/p9DlZoZvmye8ZBPThfS9cD39tTAMc1IM3SCIb5f3lGLtgxGl
A3zJUq7Ym1g5zAQ37R6qPCXT6Nu1G+fPgMf2l7dzI5+keqMKOJiObH1fU//B
L5nQNM3aoxIA9KL/HSfwZp0eV/4iDbN7WsSaFxRINhOITtMExUHvSYk3Mnd3
QNQE20kW7mm3wCPC5LJJdYXQl6YEwnb2jCPKShVImsq9/+djjgHf0uSVvlK3
xZW/teY3AqkYOLJE5onDA5nUASS7Aqkt/4UV3rqmnbgG67oMZkPWqyO/ZNFu
O7IqN3tj5e8Gk8B8hU8HiTT6imKEq2dGMGPuY+d76a46a2yCYvSC8YQvrDaI
x3zAHxR3Lbk+5BlmY0R/iOaHCI9yTzTWqtRnWNuVZ9+V6xAwXieFhHHBrX1u
WSHVoJEBs1Fk++QceI0ZDrcl1JeEOmKXXclT/35EfmZER8CnD7TGTk66bzqL
aOOYRD6oUqoQuHv78vvFI1u3sBdufS/tBnlpl+n8+ShIGFkC0sAvFkQ4xQFm
OfMS49I51buDgYpvIupUM7IBlXu8ib/dl5lkCRFsh+xSsiIqjOwpHnsUs7JU
Fbk3ZmOecHMsrhDEDjURINzoMakln2NecWoB7wUrBn1USlezN5D09LMEy+gJ
5mlXuipz/MPIFJecNB7K/SvNoph0OmnSM0HN3ge37Zmc1vn08T1D4H+OoYvc
hjXBeLJOjS5NIGW9qmQ6vxTsTnLm7ORrGM6nRWjnjVirfn/jhP8yVT1ZaCyM
5ECwbUEbMQJByQPRqig5zMXDI1RCFwOff2JUAlVZXQHfQKESKUCqBU+/Swz4
251FfSn85dJQsPfnWcMp+whOMY9atgbKHNkfKHP5rdXWq1FEvh2jqGlfc7S0
J8vy/lZn5lyALuYGQPraXYzJJhulof7nr+1a5JwDy3jhSBKJQzzrjpO+n1fe
UlgHdIr9V1uHH4na0u9KAGyQh5BKYbSSF7rJiZpOyWOuc/zJLXGtlO+SzIh/
oWlDbm2RFzrBFQfUPHwfHUssK1wr8wHs44BaG9uFisB4PwFy8Kz2+rT6lnhM
mrqm9p9slJdFkf5sZujoSigmwzH3HUMSBnnqDGeBM/uRTgursG/L8+K23hpI
Vw2rmhfYoxgxPe7Skvt9eenxCZfEbJSoRTJOrKptxQ0A99SzNHtrCvkrabVN
9PULR8rqoQM+fUaJTx43gOglqdZNmn86TbdMmDKxWmMxPppfAUnjoFHkgpBA
KLwaInq6GSkpMmQIlFS0nPG8GzI5K16AiBCuvHDM6vICxymsp6wPeFZL8Tv+
dp1WsripbaUsW2gSemUfR7zBkzK2kwozE+7x6KCM70s9j/+Ep3zHVRkPQ4ro
S2SGuFESfs1DnuiN3eYCBb1iYcixqZEHI1L/yZWVtrknWxLUkkHOChQCjaAC
GqAHeOqhLccmi8bD61ZVBQa9XYaojzeitOBW5+bAXNhGEqLIKk4vfOhhCSVA
5TsgT++lMMhyCLVPwkPnzXCfbrezSp03peypQuy8+zPBGn7+RjXp/+RGbg7l
X0C7GopuSIq35WsoohFURcERtkMuWSGwV3gWWXP9rxDroBUaFg4d8uMxQBRc
YlAlzfKUJhee2tw+EjI8YgGjO4jfhWl4qQG6fe1DKS4gtVe+RFxLEHCoqPG2
7iK8plet16ln6SaCNRW/6+YtnuksIQnIB1S/sURbfcVYp3f7IXvYN0VMIXDl
CxX2+RLjPKzwWHjaAw/7F1u/pMAQs3O1seGYBACqO94TSyOHJVZ/zfEIIXTq
89WvFLHVcwfswsIMMsamZtO+MFORCq1kQ831qTFsEO6IgS1z3YmHCbHyzYaG
41CsyoFVA/nHP9JhS/u1/i2Tftz0GvOSsejyO6LCClAAJvdhTEXj/Erz+zD2
9H7no+WE8gx84d2J06WfDUUnedyevcnYkKDf2+ohTqxd4AxBY5U0q6HbZLfl
FLSwHxoELrCijaSTl/L1FbmPifk/CPKf3UM0DemOLmmIdMhli5CL0Dos9I7q
ZzHitDIjuwZnTQYRtM8rMozC3JnhfwVQc2E2gd5X7MXVk9oWh2gl4gF2xIa8
L8/JPbavCXzbQwLIeMSHFTm5s114XaWU/XVBJZF/XE+AuTb/eytfbrqDCN4L
8AyoZblJa3PGTAv5tejINqkc+7O8AdqM0EsYLgVld+iP3DLtNEhx/cXe/6x6
5uDd6V5y/djrRcsJI8BA/G4SL33pAkoKCsoaPbsU8IpVvhdr/RpKyp4IB8pT
tJwe/JyQgNko/VlFFsAxOZCAcK0SRsWlSDmwDY27ciHrA2PPEj4tUx3AX2Ue
rQ4vTKsza+eQ9Q/X0HHORZLSg4sGOJFsxpcSBJCk5pwIwyJ/4w1kL8izBZlG
LlH8ZugtN8U5znjS5zIkfMMVMAYgGHoJ1kIY/mQtouO0vkovQxNUeI/BvzUI
wmYMfFKTRzjTyGkHfXZ/2bGiCZPP+XF1bZTuVZKxqGyo+K1gyyTMzNN+Ezvw
unObC2Z2c7uCmqyEqRHTyKdFe9EpwiCxkCn4p7uHBTaZe57xuN1CjfLANXJx
OF3ME6s+AGdjRPMmLvE00NKdmXJ9OC93YlxlX/Nd6pkezE2rFgXYpM6/9SdW
Tn6KfFRdYakz+bR7vnelD+o3ZBt8qkZDZXo/YRhmEk+V/WYqOH4nSz6PiQ6F
63t/7wOyjWrIpN0lgCDAklp7PBnU2NmsXyB0rRokWfA+3nGWTgZdhMBz5yUP
u26Q1uE111ybM7GtujzczrzRhV+V0A1sjFA3ZD1oQ6Bk5f2qadsHR2nEuk8X
4xbtVjWobhcjNh2ub1jeJgqxNlhmmnOQPd4iP8XRnN45JRferTUZRttrsiG3
oNY7m/VDWAzFpGcs9pImOLmC4KDrHol0UO4/hAWoSBUN3zn2utL0gIp1v3Yf
4QCRua6cDWyvVAYEgs7nFiQGfpWsRAc/RS9UGlwLtAloN0h9oGe6+90oCS8+
0TnBLRWui45LHQ1oFwLPxsoJ+qPzaT0VGUQ/rEtgs0K/5icU3av/9G205OK8
RbcW48HDVHjUseKcwli0nTBXuKcHZlP4RrAtomug5goZgutPctkJlMI5IKbu
G8Fo6YjAtbxjCtBUZ/ekhCrL1nuPGlmY++WPRR4/FXIAgmwihohsl4mNf9cq
2COoIT9gEz57YX4taSILDCNflkhwMZgv3BzjXzZMy21kjB65LxH+s+qSOSnV
vUBDXWK0HlRgSRAP7yX0Qyu2nFzJFDML75Rc+QLUXglzNPsAlifygqZxm4xt
WQ5Xz0buwlNqMzmGOkSQ7Q39FDXVDwZOfViZ7nzFmpWykmqX6Dv8ADHspFgr
y2Ri5PsSzc62txdTrm5O249XK1H2diz+puVqBYGlwEz/C+sv3gQAVwdMmvtk
bv3wy30ob1iJuB/uON6gV5/siYdVN5Gcqecmjlgk+8tNU7yYDFMQtbrv9hQe
4Em2B+WjYbqxaDJBU00W5FzVHcffnNM90FR32FWPj5I7ridY/g2zP5vAN2rv
UC/+QE0J6L1ZmvhY1n3JJrcsUrEAp6bHfmdRbhN9XIGtSYly6brHgY3x11UX
BLRlFHDBADRjvicrnNZdnIf2gYrYbI5KimMP75g5+T0xkbxfBe2j0S6OTBUo
/ad1uByl3zJ0axBwfDBQsz0vjuzf8oQ1rWLpzxjMrgX0cGzQhdPWB5CMFFQF
yE1MloK+QVBvh+Rk1XVqQcy0NnVmI3HJTsyJLzpeY7HkgXqSSgW6m27sWnX1
5EaAneAHBe7BZSDm+9PwW9WiCKG24ixGSwQiq2oEydjQZQR5rwS0YlW457Oo
SJd8GIMQu9aa7pfOt5nmO1zCfp4A6FJbhjwMG0mQqkn761ESM8CtYeCDdfIE
V8yHKvpMPvTCa1h9sG37DAAd3IJyWxj7l4Rpyr6ngCSG1ORUYnjO76XZwMtZ
ZusCuvwfjXOWTbp5F1AiIaA5VZohGA31c/1TQlNxPN9cf8c+vzApgkKnaYsH
JAmHOZsktnE5c/1EgKo/lFtJCfzoZG5ntpGnaB8E+4BPFbjiegviSaqU3NEC
S9uio/Stu0mwTSBWFw87aJORZrmwol1YBqNdn+N6iwuUPqYQu7yFtrg6qV/5
uU84j2uTZgrEAWcBH+/QpsJE8XWnTzyYeQxQI68SnRIw3hO4dGOF65ROsCaA
nkm9KPdtbj7HsGIzxdo+TmilohwpUJmXKQtH0fttVpe6OE19OaXYPncDNdiT
jZbVdvk3tHcvsg5pHrlXaIGbEPRE9vBJ0AfWtlgHl8LqnoWvuG5iPuV52JmH
47hkZQWj7UHG3UQBOoYxHlt2TnSDrDI1MTxzuK68lL/G7djnBf1tKeEP+Ia7
4RXy8cetDI1KMLfn+xMOa9c2fKrg1P/RKuqpj1OL4/L7xUzRcD6U3atoB8ee
Xx2nKved3vYK2NQKvF7bZV7yV/vU9XOxiZmmyxFGkwc31HbwDoqqzXakGucw
HtZ8J2x19p/zxvBXDl4aPdkLAb4FFvjZwHqPBjFOErgo0ihtpqFMSbSi6hVI
ZUiptHoiBlV2K0taibRC8d4uG85iyfS5PCisrAlyc1dEQvUZOmhxuUVmx2v9
o+vFE7iCMTvpbQ6lP24Bx5IotZjCgRWWxnNVTrDLwNpYKtlAElhTYxl3bED/
7ZUKHgv8TfBCki3OC4aqT8ZCC95uw65wbmZGlCMVGvagy9+2fgYRJ9aS6f8f
79pSjO26umJ8XaxVnwJf3zWV+L138jD8RzgV06/KtfbKn2Rmpv1Z3jPoKuCH
Tvd/PBqnu1NfiWCoTAyFrjNtUWMTGzHFO3yCOpeqrROA1VzhSYFwk/28eS8r
/0ZGpFdrDcX1WYTmtvggMSzRk3hLg7QeVMIp0BWb1KMSUWcVm9n48Xh1SG6n
iCAtOO4k6v1gSuQbHfXUBi6CW1Tr9+vkRm4NvnrBzpdo/EgUsobGB6wnkM3B
BdAh7bEHagZJJC/uiS5LFcZbohflLJb1XjnAiGOsv4p6qCGItOCo3vb8x0wn
gh90qxcV+KD2pXwGbQPUhYFTl+qM9WLkknIvS35lOJNFpE1dVrPXzEVYh/Qz
lcVVNBQza93h1SKaBcxwV/BYqPvC87JulBpertIzpV4KM1mZY+HWm0FpY4v4
J+Hr42KZjxlvBlkpY9FKkktkbc0Z58bzs88YKpC4eqwqdssPcJmtkM6ek+jr
lk84kgbkcsqIZVSLLnEEEnXR1vqG8XwHkPMYP/WusNaKEE/2Sv9djEi1uJ2I
3pr1Y+xYTIXDERUVtx3MKBCduDbo0Y+zoO8dMBcnrxu1ou+wiZx2gXDl33OS
hCByN2wedpSGu2FRrRtRKJa2ibGv2qMhjcBFE1PFl3vqlr628FfIiMu8SDZQ
6Yt1hZaGENscPSlz5Hc992Jfo8LpLpcMeEaQFjmPs2LpIR/ZyAGNlyH5dLwU
S+T7nP1yuxyQfemz1GKHqBPwTA3yYjKJJ0b4ASVj23iUV6ewfXupd55rL3rp
nnL0csxNNKA/CNsbM2niaB9VV0HSZMShSEWg5DOExKDxc+Qn5+2H22q6HiKR
/U5q2Y3v43UrA+MrofYsW8nEc0mzxbfBZPxN7CSC12yNpLtAdkItSUd5xEhi
kubLRKgU728eSaLMNEnjEGDxyWNlXGZrDyc/Yu9G9WzEwFS6OaiRGlruqOSr
q80wAOzHMx+NwHPY3CKeCltFVpbK0+72ukv4zCm/zU9zIGrUT09yeKBgXZpS
Cea/pC/hFfEt5DUiqwSzWll9KQ7Tu1Xh5mpcTbZGsFJ27wxls2EeDeR2dQuO
KZpLRS5zz3qb5HMQaRJK1oh61dwg+6TPEG/wueYa7brLn3EWZ4E6MTPIqga9
iDt2hIIIJZXJzBCxp16Vqe3FGlA92tSgTwdWvm6sgiFi8LuhoFAXKMlt41H/
WbyOE4XzJympvBjAH3itEGII8QQtDdy/QuNkGBoch/cB/KK2L7VtDZJyGOnh
Cxks8ta1JUiGgBbo76g+t7sdPhkSlHcBfn6AjHR+YwB2OfULzA1tHxsBtBvo
TxATbAAcMZShnNtamu9FvDQh21Fd5xdiiUneNgFZKG2op7eJz9Znp6oOOH1T
ENqlFutFVwEaqvtCR71n9gIo4S8GIoTHcctwgj5T+hLOqJIkEqSz0hOcptKr
ZptttNN02eGIX7EtkNpKpiEWtB0t0TdLMyja1v0NWpIzlZchOScQ3Vdyk+qr
L4D5I0CYyQCV2pPoEEZ3r13JGd5vah0HxxvkTdiqUqB50YWpPF/PxN3Mowyo
L/iwI5florcKPFNe9/U5DqU4VNU6eUh80f8GoYB/0KCRLtND/jnjmVaMFEho
8dOVS+QefWbVGgBiE8CC3//K3zrRonGlkh2K0qcqbBl+4RH+69Y3uocOfVr2
2jmDlo8tk+BJrtZEC96jWQI3NsVn87OX5d1IU38bDEtcSZhkeOU7N0P471mx
pvNlYSyOtS/NN2tHBmWTpN+ChZuV9OQt/9GLWv3EKkm5tWL3IeDKT1iPOEz7
K9lIoJd+sNEgcPOKSphObxf3xjMxYdGVlQPwKe5dYF29oQhyvM2gTps/q4zE
ehisto/hvs4PCv/gX65VEncYxrn2Con7JtKeUJubXt5WSzpxBoCOOJ17OgyB
CQS4LfMs4azLDcCpBoR+iq6VmTViZIuZBM8yCpkxNNfCFUaZyKyM3fAyjfN8
Pl63RMJCBNJhkfwM1CgBmyMr0MM6o2x81ocABXZXXYfcfIbhoPyml+RGfBQe
j44KCUWbn0qFWvXi880uhrBnKOk5dOhg2966RHnGQian9iV/Ug5zjC0zjgxX
ogplccAq51QtgyQCCoNR8aNR65tN6Yn6lyXN75NeF0xvXcnFgsbQFe7CHCTu
dB+Sbjv+tqmGscOoYznMAbRB7tnOO/KJlxPnVKg/4Sp2e5gNWEgKsOgdSagd
u0+g2K6d7wsEO5JHAcD380Ki3umF2YuHyTEYTdimz4cKn2hG36BbMx/jkpUc
QTMnI6I7CMq4TOSOpcWd+ZeR92p3JVk7crDFAcbRBFxvGDJnEJ3szuK4Bmux
3ZYqVwK717RdpDfogRkV1g6QFJquPYvVb9/k/sOWLnZz48CDk7vYjhfyMpW4
g+9+AVKz6qRevYwFrmpK6+YO1bMH+Zps6yBD9R5JHTVnvRMxjX5gJVQhjj5K
3XqlJ2eosUYh8zDOHaFzqXfnI3YLSyogDE5Epi5vtQ5Tdgu7DfDDXhHkqnWK
lin1HONe9xLTivYUiVoQ347Ctmwn9Wj5WDsOe8GHX1ufZRmyFm0+8Dr+tedF
5ncaKEQ3LwN1wSJOgXpeKeR8je6u+8uOMNiEtuwq5tvbyTEeSguQgsj7umCk
S9f5PKGnm5eNQtJv2VqeoOj5Tdoug87ly5athc7AujT2h0yeR9R5q0/y9FTI
RmOLF1zS0vLxUktdw6+2xZYD/WYsphBUzaEqn0egNz2ZpUn0GnYBL+SrhqYR
YQ6Be2TMbIpwpl3Z8kTBid6N9qvxOmSr2JVadBv2WRX+HX0j42lNWc9/yXc1
xjyJ22cMv7T1kyil2kymbQBJAehUv5Z5oQs23M3kSG2U72RJPtvkRX612A95
1NimGrzxSP+EyS89c9n91g1O7DtiyciT1QL4RXRv5f61mjRdltBR1dOWb+j1
M/wrMHprJ5fhrbASUhLCPH35WShudo+Jd54woZjOdd5vBPQhepyTZ6qQsPVC
qWYQ2KH+jLQlAAWhL94DKGqXdf5rtEciEHWDGuFXY0GzWuJcFxJNib1GUeBd
zDuiU3/3qE5epFHis28yILDxaiHe07p33/qSs5VePcI40j1QJVBsafEb1cc8
i6a8tEuCUMA/PgBrjuElt7ehF3evjHzNuMTw3YQgMG37t+gHneUimHG2Z1tQ
yAorA7I8wJYCgzyBrlUP0g/f5tWSsKeVjbap34TDINI+oiDkPOWzVKO9X6Iw
S1VcCp7iVg2LbAna3cFCqEb5NX863JnzUQ5sUI+Auy7c7J/6jlnMA1dvQw7Z
LHvyfuwOF8bUh85WkRWYTP6WAHT4PeR3t1y4t7Ee0lSzx8+OcFUkW44eL/Lc
5aELwwuYky8YkAYoBzmDwzR3fEIjbuYX1pr19pe7TVptlxgTM+/t8nLcekbF
5SpD1nMkYas9QT+hnUqhQHBNW87fzVBuGtyQQzE4FnUG3OGAWoChnmbhrfgq
+pvtvEQK5IKw2jXm4DU1sIYsqGnafiU1l8AHqPU/BlCf99ajtJU9pplglGCt
1zhSYsSNroQ3AmNdlMlHOih1o2Ds6Akn4lbMfXGjprmp05u7s/JEXSVoKVxN
KkBQ0fKCpVCUIwFaqPuT07YawR+/uDKu0RvPl7dbBFxIolUSlXTocKLoE6WC
gZFaz75qp1Id+ot1zSMQI5Pq0L+wNGp5gnf2ZOsn7gGPtlxo9C8HpGuq0lzu
AgjXWlLl5xtLUpkZEf0K1JrNiX10eEiTJoTdpZXSDuKud/lsVsRM8UR1VE2e
8OTLGLEd2aumZGqKa4Mklnceohtx6F5HAElj7HsU1OXYuqlaZJ0G4X7p1XpK
P7BjT0G674VSV/+WQ/Jh0TK9Wf9F4FvuZaJtzm7cvDgyqLI/Y8yy/BBY6/RK
JfYIcF9NW1BEbE+EoFmFW1sQyof/vDBB7E0Q+wyVuYs5BBzGe7IqdMEDkCRj
btvm44x+rfk/5UffZleutCichUAfN/yeo7EE3Xiazb7MRN9bvdABiGfk1RmE
0WW/lMeaA02hHUJEyM5615G7FCJpWVrf2ABScTy9ar6/taUS2jg/xOdbybzC
qDOAp8AH/Ja0OkMu/aJ0yKydGWrj+OTH3+NDCDGC2aF1tC9rENGn9OU54bTI
XRtDqHsMcP67eXZXejp7sre4sA8n9qXkgenHli+NZKPsgwkOaN3O5hQ9CrvC
0XoPbJ6B79glPQmGkSjzUJ4vdLad7igu/pivRU/90VCrQ4PjBwST24T2gXNk
RJX9QqD2teBo047uVNcbxgdbjqt+rD+OaI2Urjg2jEEAlZKBARbzKKjs0Mc2
NFWY7dEnvUwNd11lSqEE2EZ0O4nzwEsnymOtm205bZArYN84JYCLvsgVjgKE
xM72CWCkeklHWOqDwqklkbBHTct3nTSdDyygND8ihUz4kN/LE1B5tgFL2+Cn
OdECYi+L+L0XzbhaKrJ2mfp339pTizWYnFxqCQfnZmNRa24fcCXgx2lQ8zWM
MJ+RH2cx+ERYwfPwUm4ygesGGC0HOUtaog+dHgst+qGog3Ix9DzbcDk99VQO
DIUFpv8JosaQ4/q6rNt7FJMJDKOvLWvwPGzd2ZMG3E/JPhOABzyUIilvVLQh
tJ4xKAoMuH4T5QQqGwf4REwcO5fw6TloyX2v/ljj3mxw1XcSepdUOTPGmyV6
tcnYBq1NhIO9nvHvaJiJeGPFwLENPCoaI22LxPkA1h2DuXCjRTQfgRnwD1MJ
LvJK0vH9OySTZMWfBJ0y9Jn0SKVr6ibjbTKsU+u73Qh6afouIelXF7zKDIqA
XiCEnYBa9qGxQ4usjpW+89tgfcjvPcTNst+8RrVYtdRKmg7y5tpNNaVJ2LpJ
RazaHOcmPIxZN2M+zCMrRp1Hoxqu6n6VRBs8A5oE/mdAMfu/lJSlzaQcELAp
yjZihdWAKWfxIF+zSsQVT9LZ++uPeO71rX4KEdD7jZjvojRQEMMEjqbvqaLZ
fdOZHmNXmSZ3KrAbBSL/Ps+JTJe36Fhxv3u+RjFPcemKDSXEu4yBzjGqLfyV
iX6qaUEYOaoC1G2PIbIk6skcRTdX6dS1KwWbsf6KjHArR/KPY/24ND+P39Es
8Fl8fB7wHE2HREPIyzDe8eaRcmpLw/RnqCHzXPsfAR+/4t2j4tOS5ZPzTN+1
DvKTTDjdKelCWdEtT8hZ5Jw8TniFoIbyClZSomr2ADkjr+O38naov7j51218
x8pUAgdoPZH+eA0kgsKJbIiPlZXwRE5ozQyNT3n7xkLjfsY9C+SLJ3aXO8hu
DjthYlR7MfmWTS5J/PiKsNm+FWo23Ff/6mLYW8SwPRZ+Mj0i+SxTOB8P2YGR
BBUp8TmxBcWKt7i5ucOCrkK5OiTnN5wZFtmEb18Z3iJ3NL4jp1ycwu/AQaQo
FdY3hPLWwg3vWdcgJ0nKmEXO6HNrfbVhS0YW/1e2nIk4Z+9pqeE7jmlUqqlk
Awowp+zS59gBJNmwo8S8saPJRbLKfizmYz6CUIsb8yv4R2pNIDOAmGyAptI6
RDVvR5Yg7Bs8TTPoRT7gsnCOV9aCDg/iHcHD0x1BYOOSzXJYGvubzU9QdmRS
SsuigsKK5mTarboNWcvMtqcm4HFkG+N3POWiP3R5fy1g0OV96q31NJTgAB3X
u7fJtcH5KCz7XEbxtcXpwjtG+Bn+jAwg4prYzL6QZEAiT5QRbkKkKpuRC8m6
plZVmIJHuHHZXIODLo3YREjXQG6JMySbPd4CAd1pkzt6mZEm51Q9t/4MoZGF
QSx5Mh4JvY7NjdkMk3bdeCywnzMdEcMWI1UQ7T4uGZhvXxI6io0BN6NJfR6t
WAD75bCGs2F2hHTa8MoMbyLFsddod+1GBvEownjNh6am/gO6tR8PhebEeW++
v06UHGeOsJBChzf27ObgRJjlNamGtS3tGCANmx82JyQV410zXR8be2GmTZYk
7tG1nul95dOv6P13s58yBZu4ISDhCaMQJBrQa9gGxVKmGt7gXVtcgGUnH96+
3UF++qQ3U15uWMOMBIBwscoieWO/UfHObHLsdziLiQyI9snUx5OZ1P0/Ns26
7wm9BDbziRPS5i/rIIsvbhaLRw2dXQkNmrJCImQpc/Yjl+ouFaE7QLhxRwKc
dzC7MPNdUBahkOSjxu5SF3AwaGO+vjHgsKaGlV1WRkwpY9UlhpaKtXB0nXcW
vdNRcFW00c2JE6u11rvSw5z3lwrj+DuStGHgbi3GW3uUUMJ4sXJk5Utjpa+O
ZqReB1UuffDhZdqmA+4zBwc7+FSlu6GDEXglV1QQdJEBitQwoc+icGptxCBz
ELtUuC20K8d3cLuKpBmvBdj6/9dhnmFoHudMbAfT+VKjpUkgCyde5RJgME24
GDZVTeJ/xaUA8BzW1tn8XUExYMq+COE2FSYxB9BwFp0G0PGQXz+8e5GkRo8n
URgRfX9/4uWTHKdzrsPhRaK2pPT+3Ka0d9Y8h/IWZT/9bLOag1Q7mN1RB0pw
dSFpd/geWntbkegL89/HRqeAVP+4bZ5NH4J6ej+LIcT2vFkAvfIiZGhYbiVY
jMjZc/DDZ29GWYI/FhfBeAmPO8CharfHzjbmv6P91U2vNGCqZgsfL0+MFXU4
Ttvy5ymbO08qZ/zVKQs8u1jyWpfcW7wQvjVR0vLAusSkWhPrNm+eMTYmjmkF
MDT/PDBbZ4dyFtyiXLY3tqU3Gr2mJJY44HNLOOnGzBc3nDGQT1CVRkuKDhNg
gOKviAX9gljSX0OeM7pMNnPD6F7tsveIawBmzLjTMfeHmp61Boup4ppqWsSx
xTW8AaZYe+HtMPB8KJ9cT9TXrCxaoZIxSZ53X3CCiPYIMAdd4cJ7TCc47MEP
SYwR+iqSOgjlqKv+hwSkZvk+jZ72ySGaIIuXjyymbYpzXsHpvFOeV7FoTjju
wKMZTnoq0LG9hovK4T6awNoLrX8vlE+QKx+MchliUQAm2T8tOOCu0XBXMEPs
ImVIq4LQNqYIDMcflHRf1VZjvbhexDwpNdhHmlol2XghVl39ghIHm2f6vxxy
KY+kmSIuZhLaabsPeSdGFIne+C8lZjZW5k/cYotMuAEDkM+Mdpu67OjGpp99
zM8Ihsm8GgqeJpIQOa7+Uum9HZXSzKZYunUHbKgb4W8eLcB2qyxb2dGwh/dG
2WkCtcjwtX7nLCkqlbTplPi6kq+ZQIFiBRKkmwuxP2YgYOevfpDsExmSRKJu
Ahv1aFGIMdbHWdCwxS2GnnQqj4IBqy2R/CrZ8Y1UQ/D3xam3n6GjAzcYtVmm
JkTGKbN3/SXMVKs6cdcwfvb8vi3MYu4epHgYehLQij5A7kugHRPJKgnkalXY
4izMoQ6MNbrToTNf/z/+eEZMvhFr4gxhvbhMIOOfXlGO4YhXhWOiHuEJYuqs
un6Vz2WUbGd49wQVlGZEfdkEOhhPlGl0B9eTGxnY33m1D9e/xYi2NJx4pQPX
xDS+405ewv61tyBvEJQl7WFsn1oVUQOqrGHNHM1+XAZjYMW5oqmnAEfSThCI
UkgDsoFgr+LLHpJgqZVtxfPl1S0g1rwDEFcEED2D/g4Zl7CWkbye5+DTWA80
2WUJTzGd74uix8p/Iqo650J93FyFTLBSH3pkAI8ZffdUlf4LNVJi969kVPn3
zp/vGA1j8AYCv7Yz20H9330Cj75Nw9i2Olmm5sHwz4DPYnpptCO2ppe4xmUQ
t1zzPCYsDqEERELU4rZaDnWl7qKR4TZ0V+BqBgIw6BM9E2glN+fKZhv06Xmd
SmADQ9DTSU4MKQj4JzsLP4tI4fS6MkipjIDD3+4lWSnpjQg4GKxpiA2rL/V1
D1DG9YDoCfw68aa3199K4HpKk3b5IVwty2pqvjQ/I6cUpkfZyVtWGYS54MgW
ERB0UJTosVuz0E90qbfW1bk3Gh0iu1qXQftJBmxeCUProu0HChbLQqNFOrbX
i3s0km91blAw9Mb9FG+6ibw/Rfqqa8MK3Du2TREVOU6KjjGc5ssNHm3aZ33X
sHUaJ0ocfLX1Sd/Kac/wPTz8HIsvjUsrwqeTviWJTQPIDdtUvkgMrnKqOtGV
yYQzmjk8q+8Dt6yWQrcgFnDQ9ehjQ9l7ivheoubcN+xw5xD1eqW3MFftCf8n
dIotC48i3WoNuZ7obejRtoE71YWJbuUv1bM8i+P0IPUGHBnSA1UMnfPrwq9l
1FKXoOSypPJZ/DD70wNeBU71n/+4MfHyMUDtzhnn5c5BehALu6fn+eI6zQNv
6EWT6a00jO/AvAKPzyFZkPUaEr3GpYtRzybtURLcWe2jV3Jv6RZHKPUm1z0A
4gsc8oHLkgn56dtS+JeZ5rHrzqu524nztXDk0ahTItrjq+TXfli2aHNMcZGN
wasOi1MnIOJWdhSgc3cN5R7QYnkidAgM75Q9umvQaxeiqQ3/rsc5Mu/kcREr
ql0/M4LcI34oTN7PNnug+N7cr2ktvGSvmWPewjXTkp6Kxd9CDYPMKBIAZdGp
TACmrePGaqaiajc29cHb45Lt98722A0eEfj4i39QyTGN7RXZRMCL6oUQ3vEq
vIqTvLZM0xHOqXd57S0nj+Ngll9ls8c4b5hRR9Otcvcqqq2arZ7spyJdiKrN
WJJ8eguocKynfwQBKlo6VOBJBFmiGRZuy3pgrsRsG6cA3sRQ0urSv7pMzOGD
Gvf5wu1Xg+JJfKOh8p2pV7I/tYHILMTxK63vvZGEdhdoeytw0zkgZHhLTIqz
JDccS6Awpx5WoqQVkBNfZO5e8iDbmRS2UtFQtkn1bkZNLUael9hGoO9dAGAS
PfvymlbmsC6DkXlMCVR+5eEeuDY+g9tsR5t/TczBlHXxjwIYp2ooSAwtljUR
zRgYU2FC6+hYNlzsA1Hs7zYt5xfdeXDrLdUglS9MMi8QAMmVTgNQrwb5iCvk
6bm9fsvAIpFcK47PFnyqvqP5hwr5dkYI4VoPGSa4df3lf8a9kLifgQ+5riCD
5fBKwrQhaM2j+9w+J4AIhJxWpdCsgCHlLRn/mcVDv8i4XQ5yQ/5hTYQ8k/fc
Sk5GUrEaeeinEp7+DNXGvJBrjRu9HuGz+QzRL8TVDhnAanLdcBLoSx4NgMFn
4KRVuKRh9k1yMz/cgG/d3PnFP7jLkEjQfrJHbPx3VDw9UVuIVgYma5NE2o+A
iPuKV7zZHtdptHcL+PIK8njsf/ELwYTkHl2eWdL9/f1h8iBf8sOJs9e1qD/z
9zhlwxvQ+6M5MxDv8JruATjwo+s/Epot2fWAvGzydq9odROQo9yijGbkxZcn
snppvan3r+VGSVbASBne0fh89uc6mWYlDcD9IfeQl6iBvcMXhsBTmxL9qgb6
JeuH/kE5nOIE10tRnOBPadTsMwjUhaMWIlttBYpR3+TXoHHstAoLgzk8pGat
7vFu58+WON0OZxdBJfivvnps1wWhrX93VpG079iFkwfX9Ougwlwb1lbW19JO
xPc3NhwvANQvhsQPpQGo3bGpYuk6P+chy8OiThmVKhXSNOH1mVkxq8TIh2T/
1Y3b4bEIpEkv+nKv9TKJhHwppEPD6PVJdD67tUo3ydHX5Z6Ph0FR0LBGTA27
DL0r2dc7gVHJbEzSLYKT1X8sMTHUlPJn+AB9nAOZ/zXFK2+++pS8dHj0rAIH
UY0pvvr4bRr04BMeOyXKrAhHNTDFwoxjG+Nq8fvajQlnDWkajRjO8i7r2Qm0
U5nS3Tqe7qWmD9mIIwNZrq4WSl626rnlRwNQQt7BRXTafVWypm2WeIUNyecV
HtPs4WewfApFLsDhcap3e7V0HiN+V5MInwVNeljbltGl6wb2ovwOh8+OsqTL
Sbe7dFQZH+FWb1yhXpkuNcvAuTo44vYlyst9BP08AbKop7fnTQV8MD4r2JCd
e+iks5RpPQokwKazU97wcF83jfvM4Qk/HEERSEkdTxlaXwK46D0B8MDu8DRO
Km8I4ZyXi+bNgulfpHrV9MUuykmq4HmGk7iCWyrQ+9fiJcUH+j+6V/VSiaBB
ITmj+zqjQd279bAl3j5FhzoheilwQwC5GyPrv6/KAoXRjXKdOBvmKKTs6mb/
Fop8yjYDLe7HLdqkhAmEYt1lBDR2FRRN8EbnvRl2RtP+X9hQ+fgtIwdZYkPr
26tBNEiA0ahBdqbwSjjFjZ2ohZlK1yFd5S+9F+v4hhpomQuqD/8+9XX0UcYo
h1Xr/7DStdG07Tsip2GKpnz9t9fWo52O9LC67u8pbuvGB7fyJm1qnK4Mf1Ik
BZJo0DVUVBUAocRyacwU5NGiGYXUAte/6gy7gmuj5d/vLm9LAAnGfMN7er9P
fWYFFA7KkKkTuD94CuvOP5TW6j5yElEpafEO9DNvEVHPsrzb/RPZxB8EpHyt
zv7Ihh+2mY0gZ4E9/YFyKla1etwBl9Cf+ebdPgAEcgq1BO5E9m/saXaEH+xf
WI8oSbgbb96k1qAtidr1UExYHBmXtudCS3LxMW/mmYOyrfAcTMkdzRfWQbQA
No0Utd6SsdP/jwKV/xArvhg0zPUcJqEe8riBHKk+wN44oDfCK1umIAALOuF1
Dq36SvqyWNl97MYPh+wySDOI41P7c9lpU94vBPGK6QNfJyIrwMxQvUXcXstf
1POXqTb8wBAyZloDtRpzkACwagFnDrfzTCGBCHDkT9LrlOE7JbxL02FJ3t6+
RLXSnod4nsaj40cz00LBYgATnuvLlQIsAN3F+bcsn8Lc+rffDB18aphO+8yP
vAiPj02u8dFnjDpTUeY7YjJCvSOZurcJeiPTxs4lLMh1pxCzvslrQCgmyGAz
VjO9IWlaUCQIy1aWK54pmmyX3COqxajVW/vKES0E25gkatxWJa2Gr/Dr7w5I
pEh7W+/4wKfCV2FOK1oD1pgBXF3IwshvkPZbZraSGHS0lWRG18QZD/vFfMwc
pmEfLYxd6DOl56WblFxcql0PntuwX1ch8cfoNLn13OeZOuP6+luQCne/R/8E
JaxAmuADAg7SKpJ4PUh9qGrjzH7Z3ICdPy2v4wkUqX1Ea/OUeHiKaRde03O0
z8QVnGDPlU7jMIQ/LHCAsma2YeMM6VRChFIsT0WVVVvbOVQaSFmG6QHO9NZ8
+Ao1CISBDOc8K3sgSz8Vgv9SaEyY+4ADbpnyuINDo1plL+WoLi224oAEu2X/
z6XDqMSnsjdWg9BWmFs+yBUnTLTajEQgxwHdZ6cqYdBIWC+d2+D5Ft22fzXK
/CrwmG0Jk3HdtZovrzTkoAlfDkFdRAu9TiP1FDn+DKUGRsJu4ZqvA4g9FjCN
QHcl97zWBICWd/HBm5P4562ZtYImTj1hcIq87FFwMsW5ccXLIOGMnyz6MvsU
cdQVPrEDU32BhclAl4u2sEDw1FdlfgVPpMQ72xZwAnQJ8d30k2wRtAj0Rczs
B0oiOyfAz2V0iT8L0W/hooDBFaQTAQAPpLzCG6jHgMxLGSH0yExzOfEiu7r/
g6fz47pgbs9aer6ta5+gWo3poxxd6P3fqTztudGE+nfDRA03jRr48oGiSSAr
zXKZwB0PGNwJQx3Kj3/fB+wT/27CucotF2KqY5X0nCzgSmxyDmKl36ANciip
aVhh3gof9GpzNDmy0dSA1TNyQ78tEebO1n58TYwIDXg432RBgRHVkFZFkyDX
ca0vCl7p7G9sHECvy+lNGQfV5IBc24o8uAg/sl/VF8b+OkDNirAl6u7cv+8v
zj8n5ofaNPoewS1G28PkGwiIrxsLqA5pytr5W8wUw6t9508BkxwepgjbwVMH
/tjvE/Sa6ncMDJ3hKGA+3p5pvwWnFe+JoOMa75+aPV/y4K2fVNsU6SfuB6Tt
Wg6Yn55y/HWVwCeaq8XKzPwCK7JLZv5K99WTwOiDhpBs+XiBgBiOQggCemes
sWs9ZvNNv8A9dunSIDDU1RR7D/LEliakGkgCyoGhS7ptNq0kgTb3lwCZJKgO
+CFW8zI+iq5Sb1gj0Fiq79Z+r2yUHie3AYCDqn3ZMaA0IScp/BHIUlum+lW2
MkORVzUpHrCXeq/47jPXh9675zPTCxtSqxeGydtvLNyVnHF9Ow/XoQHPV+hy
sMR4I8l1ObA6ce3xz+lpk0GNP9zZXLMssT/i1q6tvK2V6xeOjfLOGZxwEFmZ
CYjkIoUiyWNq7OkrbIu3czpi6l9JroS5C/TVWrki3Qg97LP8OEFXEVEBgrCs
IUHLWbLq+OZw+3K/l5n1ahVu5O4r0p5VI0+kVOL8sA9kIjUMYcJDzLClkkn/
ToBk3QrCf//wvAAW5QuecRLVupgSIvNh6RKQMGBtVF6EVs9hfxELrVdAVrH4
NoXXPmXmnv9vu8kqzsDEjRASRqHllw6COW7/u1YzFsd2icMaJBy0BoZznij5
OeU3+Y+RWRrVVLu4JJi3XcAOm0f9IMVVO0LR+cZz8PGs782EeL0Nlr4IImqt
qNEIlJ6AbLiXpV6uGA+Uac8quKQFrvcjaw0gFbTfzK552Ku0lfMeIFzL6lr3
1e5CbskWdyL0+klma4eXpR5EhQmeBtFOm/KSdY/zRFbKIqTSWzQ5fN3qmLtP
wUGYR6pvFPnzJHGb1noYNUSq1qiTmBS5lTr/6l26VOBWNZmD83pn6AqEBUw8
sCkD5j5LMEv9vJk6IDP3aOytWTnPinmh5IwDmdj41mE+qmyCKB9Pllyk2US2
iwU/LXjG9ecs8oKyNMzH/JJIzyFtrZEqEqN6DotUj29TNAx+uarRIhO9YfwU
n71hNVhn0mAlOM2Mrs8CCSMeRDg21ccDi7fLK8f9lp2H2GAto8OX/Y+/T6pQ
cr5sfJlA3YgnvKn/2+RR3okhLc8lI8vPpbrGewaAxzZoV+yNWBQPE7qUGoiI
rc2uLlOf1u0GHwVoUHkm1vspYGuXaH4ZiwcjizPcrEK2btPmV+yWeNUoV4oo
6Gmdl53Wl2Yg0EoYWln0XTy6CY4epycoe4qMODqdlJCIlghKXZJxNt5Yz1VV
iSP5MW6jwfDgHUSy0VYveCrC9iWxKNCOQpMQ8kSvugHsN+0LcUdlaatwDSCS
YTyrDKDjhfpaYMyBi0VHQSGXhirwKobQ5MfnMw/akTuNt6YhEkpzgKuouEV+
fGfs2Bf8WIj5mbK1W75hM6gH+xSLWgWlzEKAe9oN1AsTnuM7JE/Oo4nCf07h
AO2YXX0Ox62Zn4Es4BJCpRPrrfKkv6Vr1dJS8ltjoCculpWuscwy1NME159j
O7J2McMLn3bmSpEjgx3u6bDjBTCirPnBQldmZ2kfiHG5zaMA/Yf9/ccCShI/
mxv92BYHpqF4C9pxrb953T/tBh9MAHB/mao6Nr6utnyADntQbQeYALRoT0pR
EtBWmf9Vx4CCo/6O2mJaH3GUMNLXuOHV1mNZwfsfFCToAx15lZomAnckn+IK
VJ193Oy+/xQTOo57deZZffuE774Ay1BCOGLxDuZm3GfAOi/RqlSKOeLE3Aik
wYvaEJYx6epIZP843Zhgkvq5fDiq/CyW4OBlPpSy59Y+FVuV4evYqRhHm0NK
fZBBRTCzIMcANUwxpkWEGxuup1S+8Yn0FyXTcifbsgiDJCMA/dgAbdWTWopL
w4VO0HeC0AOI73jcMyLafMlePfTYwcWA5a6cwS0WGW1I4slnViHCUpkW32Z4
8qb2KQAZW4Sa9v/tS3+iawEtGeytOk+9R5vqESyXPVqT2yJ+XQUur+lk87EG
6ig/f5fxxt0XkgIfm+gJsqNhQc8rqzUekA27TTnDz8zPbGd7G9iSGWyZlYc4
6y1y4KEaNNBALWWe3dWAHHk3/Ynkv7zwSUhuSGQfHHxUd1NJOv0JaB4f2Bgr
MsZ96jNEhmdQmAnhD2Y/OAmOFaFTdTvRX9e3zePmUhTEtomIDmjQzDx3WX9i
2FMe1jlesLkm0/Ft3fXhaCigsNcJrF4cKVR0/Jl6/KqJlVL0ma/gJa+ud5/B
7+1fEvUPjsmsuHwKjZuK2qREvo02IXf4SbI1WZn4Dl/P57LqZCd7zgbWqkf3
u/xp1M+MXOrC2MwZGEld1XGhjF1lU9gKLIGjPQ3bxwm3NZK3Mfn/hUIi3D3J
lwwxvc/QERkvACAhBanIf5FoYy6UzOp+xjwQ+DLCyS3398a035rYqf7jyNdk
qXkDkSpEIipPkS7H4Q1pRmgjedB++fVaFwxOc1qFO2B/JxX7OYD2gcfIzuHd
KqfI7y8RFutUFN1M6UeNd4G+H0AkKhAMHBohgrSmkwXssDfwNIzFsVFJZWIu
LG4q/fq44chvkWidjStxWLCOw0RPP6MtNxSJ7KB9ESVZ6NL7O+Xfpn1Z7SH/
i5uP1TP9YO3D1eB4uOAZiBhQDjGh++rsF7290MD53q6p0rBYc1rtkKygLY/5
nkIZwI83O9pDlLQR8xM5sM1bVG6VcOE8p5JCt5vHq8Vnj5D65uyEIH0osv3W
nc/9+3exCjNPQK4kR2zCffyD6iYLVcLQAeoIMq92jLCFRKkL5QWttyY/fl/A
rKtYV6kQ3imyiKz8j905wvSS+Xn0c3iq1OwlMp5hwrdrIiAY2QyMKN9FoGnU
+jr+B+JuhZbpU4U3HWlmDyWu0KkC/323HkLkn891KANpFyU5L2BNGOXfaoRe
qWtF8Ml/xkefBiEvDXa0zfJ3QSSDf3By5r5X0xm7rOax+IUvzBl7M9Uov317
qR7lkv7T4K9D2ay0PM5YsLsIAa8sDGgwcRpWQg0YiRyqDw4FgZozDyjf0qAl
csZKJ6trnvXrTzs4TxId6w053aXDJVMsuv7ul5ma6vwCPp2rdNIMkWK2Eq/7
K5Gfv1yCTUtoNxMh0D5Oe8Vsf7yxkr80cNqE0NZqKlNnucHzOYtDkaJ84XS7
yn3JczaJ8kBtL/ffMLCrbm/1IEJrJcRilsc6i3JZyxgOSmSmt6+07yDKGXRb
s2i2BTQh6+axp3TI9oZGtjfwmDnFEG0fsvYX+8jCTNsX3xMCvpv+MqQvO1aO
jPlL1JN5KV3qhxgVD+v8UhyNYDFWNQVbIG2Ce16YfAuqYcSiDcKycFOtdtfh
soxGBn4LwAdhSZCjVsQ5+ri9fHIgrYLbBfzL8r78gy8CoeO78alypOTNk2jB
1ZAiWvHAUAHJJ6e3dllBAIzjDu/rcLOkDJcSi6JSLHIRgMk/H5HZF904Ka/c
jsdyZzaN0WhoQyjDhnyW9hR4HhMHfm7hKONJeqdNG0tW72LXANOPPuv3TDAp
aUp7Zu1QuM6n9iIn+oN5lC3jTiQM6MbuETbAGM9Hj0sjzg/Ga9MGTixQaEI1
M4oB9iBbA17gOhOc03tn7OyyxWtIu1wrhMydZgn6+Nf2Pm9KmC6LchRJUDQq
+YE/fTrp+qJI1twJA4lW/rqRrmoIQU8juUVybh602wQEwLVAITiItneln3AP
QYnaaKWaTU9roPp5xGO+i0H8BGw0GIXWXXa9I1GJ6MEL4owXWUT5dhRA8cuF
gVeGsYKY41ZvXvNTuQpVcTdrwJUd06i26R6/iv9BE9cxdSK24tqRy3mrUNhz
4uxeB1A2cZt7T/nBxxbi/ML0+Ry/Xwk3JOHZ6ocrTu4h7L+5+DDw5Lm6XWSt
6FMmTg62AMEDCiKJALkv3Eh7eX9ERfTppDQQmnzf1eJfYZiYmU65K9Lj2dfV
L+ZQW0A6WmehPM8TolVxHGzJ79CNDmzQvUQ/95NHwAiPd4TJIPwPtRKzaehp
HHUW/KRFjZ/+xNJs1IRAvF6jHQGqyCFLGW6I4Da5SZEQUwnZ3WqGivdJomAV
mzsEGyw1fiIzqA/0hex3dhQkrRBQaZLQBpsf/1/DU2A7Qda5Bvur/UQe8QFR
O6P5KBjZMnbc6DatPBXxugJ6J22LiczrIiI4yHRPiD69XvUBo5WtyJ07VZO8
dIP/m+7ZMPI1LyvDLHgNEHHLvPAryf1jRw00sQOnz2Snty4e2gOeS9gXvSlF
Gn8wxDshyze2ZJ7CLd+eiueVc8bH5U4Igq+iHwBzkEZPaZreY696aXTNXvjg
Ob7+BxiBawRXnmJZ4oaLXrFGa6rSPYk237+8YTUAR33xagY8tT1ZsNZZhCX3
DeXoRHikEs7Tw3Lo/5JY/89X/hkF4ldmbys2M8s2MZfZwT/Ms1Z4JpwN6jfO
kygkBr36mX7Tk4A75eZH5AeE4R+VFvs2K6hBecc10kTgeIYb24ipyZCf8hHd
5JiOb3mfvKpA7bLKXCRxNQp/fXEmXEmUJmOkrVLkJUUeV8Pzy8fU2sFXSBcv
6qXHqGLcCbsQ1u1T8LJcI8v1h6Gxwl/caYYVILNok+PPL3duV5qXXj1WwNAr
tON7cYVzeSP/m22SEpgqyWOvXvI+rEuasF/pa1RtylVDZztxQWkyB5OGHX8J
b4GqKKN+/P6+8e31W1KTrZFHkH6FPTFGPD3KZ2afy5k0J/roUesVc+jxyUsb
08BjS84xWqd/r5Owxa7u2/HJqxskRWn/UsWa9KpLBFGHlyYwfEU9wu1Pxg5m
UoFCgJzDXJSGOT1geEhxQUCXCaEmgx68OnCgCIhq5rdYWeT1O2hna+jrqARO
PFnDEXTAEwd2LQwhS6A+YjLOzLMbw6AM6/jqswLqojBjVYtUtOxGSOA/Sqpq
iCkVMp5u9/ccYIvIVHjDjrqisZ5wdA2AQcZuEMWiNJmzhfA2t1BpXmlSPal4
PZWcgunP1noBfiCTqy4LjpdkUa6ItXEKJSxMVjDDTAZ6vkFrJBpWg1ng/9tL
yZDAiFW4cMddP2S0CQuMm/0hY4reXMqFBDgKnVH0yN1DSulei4tJY6AG+M70
1Skts9LqtmGAkgt0zdpYmZmt8gVqkAw11aZORC9Cqs93HPp7pc7SA1n72mu7
jRisviwyClbzCFt4XTw9a0tP4fLAAyxVwPimlNDKhlo77p8Db2jWbTN7aqqo
G34m17i+eZZBx5JlIFd553zgJk13hNTokMrk5H+rFcVZ6evNkDV3upkvmcX/
jFaVhnM8iLGvCSXhQAcZkI6BXGVFhC0RXt2UBykXoYquyyauCIa3irExRmhY
05jlr9CJmYBxfYYvTgg319TLws93A6RcHHKM0u/02MKFNcSn6Jql8zCK4mnY
XFhtiYUqrvKM1KLmteCl1THEydsFeMxKGjwYcdmi62hqcahgpBvoXNwp47QB
RvDGqkcclQfw3bhCPFT84/2R/U4540NAzmWN9G5oNJJhGFZRZ/O8b9dGIbGo
WbYKpM3gxL6aDngMrNocHS2+j7MZpBBhdB/kBUkydZsNHXuLl3mt5U2sZna3
67RSJaiDW7uzlXpaLI8AIhY2YgBxevpUf/GZ+OGMKxhwU271VjVQrNZnnpOk
HYNVTb3CtEtAR79JRkBsz92a5mmQJ8D+hgWHlRog6iySmxXMGtbUZ++OB6yf
PCeJeDfA2kMAlYQ3DIeu+5Fs6PycjuOTrmrYi+4XmozdcEwMDcVYV2Ui7t5d
dHXsp6Ty2/upfvvEAdjAZt9orQ2XRXqpsy+T6FU8EorIq/kD7uV/vSIO4Kcp
KdgRyHUPFbLnYGrDm+o/eVwk3PpRcr9xb4stnapPboxZABD6VuwrkuhTc6MF
Uo+JhUh8Cwg0DxwxkaKL9b05UUuiyvt0HMhWs3uP7fk+e1npT4dwviBQ2zJd
dWjzOrvfYbZ8M9UAi3G1iRbIjJlBT9D3FS1F0l+aByAdhZo1hZYhfGVkSYrz
k3yH5/patwYia1/RX/rvTy7FdAhjpcoNgIGSvbIYN1KbvNORMpiPMPSwgm9J
cxdLtIgzmDPDZTkJTPrHRt5pCX1mG+C54ffp9WeYNeST5Sr21wLg3vJczQmD
g9Ym5R+AEsBO2NDMPpsHbr7bshstvJgva+LZnThJRdozBRhzZb0EftzNal2I
XmNCvgFQ6gMDhR4b14ZTH5c7V7VTPkIEkDazl1EGSsFSBAnAyWL7klDjGJAl
c1TXUEYEjhkLGadM3qssYg8emK/TmBijn2yj2zjdNKI8mqKrjtUwEaHhasf8
1pphGOmzxSASxQki48Sq4CUH2RFY+/6Vs8mtwZTozK0UfZW/xc7ao69z7bYT
/h/Krs6AcNri9GJUqjs3xCRypeBQSvKERDdcXIxtz2y7h0TEcKncZQRI6py8
NbBSlWcPKHvKTgx/aDsVHdgyJ+h2+BQv8nsYPNm2kn9XYjooXBxGZ8qJmztt
RwArXeZgMl6f4/1ZGy31gQVtdjdeXMNtaZBBuyUWlJ8SeTI5vO153Iw02S1c
+ZUCGEK3BkqNxyLN/0DBYTr1FsrNWNxMLshJQas152mWY86k0s+46m0sGKXg
mvvUo/heZdnRKUzpB6xtP8bcisHl/KulikpFRjtFJKZDP0dRUG5rCLP0324b
5+wEvkrvlQYg6MgLFnIH2OdqyXHbuGxMZ8DPAbaIkYzm/Qjfk7FTb0oEpXrR
fN8lhEWYNdPyJylSPY/jDTVZZXw9vytsSt993n+wm5ISAqyR34BdJ+WZfu5Q
2S6ik+fw4xxf7wWWUn9+FWXBp9AtF+5Hm/1PvaMt0oQME3Yudg6nKDyHqFpp
idTewFSqu35Ux7Cb8Jh9aq0JQcKStDYZdBkpb2RLcMLTJ6rfF8Ldt6pirvkF
NkPgHl8XsRvKH7VUz+toBRCs9b1nE6f7cvyX+P/EN8mM8wpFXWEIICNQp7te
lRKEpd1UMeYVhZm3XHQiSKo+hVExzfyKdiZRB0/cv7h0Zhv1pQTXxMUSXgn/
ktdw4uhfa8tLxM6cYee2bJiaq4JEtXVmLl3qtkUn/aemDE1nWZeffkFdkk8e
ECsNeCNiuku1+0EBQRl+DKj75hc0S3BjiBfTwUfjQYtKi5hnSzsNzcoedPog
xKT9EEjMtXrZxH7SJuEZz+J+7K81ePYdfEBL7QXTLlOGSu29ez41r/kguFtk
cx5+xNW0qHvApOxVLqW8UYZ+tl87qrsZE0pOMqVUZ3vlDW1wFvpJrGzlhraE
CxH3RK2nn5YGuJ7K5COmnFlu3pSP8jscLtKFavR0f0YojVFNk+SMZ9ZR7rW+
IjEl5T9W2SeqnLT/cx0Lhi4qzbALiGB+1ZwkctA5dsDUl/kjNlV4zfVfbY7A
pGlHubbS5jDJbU0Pnm3cVT3Xa6dVEReAX2pve+zs44pEmku59xNA8QHZs8io
zCU0IEGnwCi88yxnUW5ABNWyzCK33de0YgSG57CCNTd4mhJvSw7jMz2LQUP2
q0K4pFtraqmipNU86NiOi2WxHNsVUutUMXmjkkX2Ccd0GYuSjm9OE5OU3zvb
1Qje9opjELIh7uQoOmSjvQlA4qjySqORfK9DnY5Cik15kcHE/mhB0YMxJjCu
E5HlV5GWq2RTX2qSZsAuDJGMeFnznGfPPK2cP8Ry4JWSrQ9GEqv90aOM/6ZH
sATQcQli5tUYP/GnDMI4uJU1hLa+wJAx+j1JaAXoFODTnOZygH1VTibTnz5v
WgAVX9KyuwGGaltHdT7Sz4B2yzSXCjbO7HI5vg8nDfGLPc+9HPV4IXEMbWQ4
qudgT2NSVo9kAJZ6qI7XVLQCH0Tzi641VUxarb2UlKTpa1E6eZW3V2ESgBfq
zxbAvXDsCYKs8OqvF6MN9bI/ixFLO3ok7CGIXox1Ca0wGaw6gy0rTnvwZbFC
qyHRebwBw8Uec/C3YAw5xwMI/HoKqe9CfCOL7NVqPKHfCry+9p+LbadeLa61
P4HJXf9TEgcVDWhKjGX3nnVYHNkIihxNPjjcu4Dd2vD/mgFM105xJ/5RMw9G
zbLooAu68OLkGaZK7MWowccM8uoMiP/PFbBG9KM6xoqiAtltp2r+doq921LR
vEqr75g6A+jAoT1UdedqaFO7s+ODsiPg/1YkvYwETKepFf1TM3VTHeIpZcnQ
FosZnX5tXbKLW0dbKAP8cxeuHWJROkBAsM8UbetgscNFKe8TKL86znptYnH0
QtKegdGpX2j75gAcR7ThPioL4UPF5s0bXWEuVJ0x4EJV+b89XTX6M7HJRONW
n7E0GIdltoNm7Q2BiVXpi1ugTi/4ZRW0vcrhU/Jnyr09qqYRiS9o9wB9BEY3
lScMJdObfgTwx7WtXy8ytG0qjf/GOVksnZjkTWxQxqdLyqAzliBb6itwSaQ+
QK8quG7g1eJgvjMf0mY9dgZtRkAH58/FFTlSxz6/UL2oWwRPWF7YU7BQiYw1
LI5M4Vb0sOkkcX4BracvPGgpoj0bfvAPgsB4n2cbALBOL7Px0KjYtHQAJOfu
FbnzqCCzFpSiiJmPfyIde7ZyWoaE80rQiep1uDYc66Jjjej7qcRG+QNVL5xt
qMRXM6hyD8M9f+BRCg9mLy2uj0jMeenv5fvNeAjk3oDZGVtlCQkNfmAAOQn6
FqhquX5MsyF22Y6FRPIevtxI34D1q2Oc32m0PNYEFGXU6T9HNnOyHWyqiemt
YV+DqRKPQsUHZ11SN3wp3IzzIIrKuDuKkEiZow6mdAx15RcHxRYQwLf7/01H
9q+IZ87uf2TsmPu3WOr389HhQZ23aXa18S/ISHXAiyTYA69FXkxUZemQrUlF
JP3eOD2XQuE7G0Nmb6QE4WRy/Rl8TuiZuWByICZdDp51uSVTVH/JFQdwUX0A
5o2kSgtGjRjRUzWEreAL7/bBtHwqjEf0orcq1dIEttWjLQQAUhrzcC6grI7h
J7ljrnBRcdtpDZ+TpkSlOIaxndd19LVgqLkgKQ/6IAwlu73Yk5Ym9ryRJ4gZ
UaolAiX01EK+wejzuHGRcy/vUM3LS4pm0X1TGhrRVgziJP2bZdNL/NaUsC5r
9XixDY51F1qsnUrImsX1HCzYsJmPAgCzqYbi9vaKJJZDCUM4J3z0srvrJr5p
tREji6fAQG0XsT55B0gNfkIh2ypiJRlor/vx6sJulqObx4E3zsaFbWFsyN0q
um/uqx/MBeklbGdxYB/oktxGkweyO7xhr2+9eY35OToUrEUiGRxn6kRLpVg8
3lOuOAwUAoGro1FE5FHW38kQdO2NuZUeYWAgQpVL9e2Zaa89nsBigxGeovIy
cTQeJaQrKr7XSNVOt0//5DA/k9PQN8Pa09q2PRkjjMXBWC9G4FcCToWktASx
6RLhqk8hNUtaUZiadOMJDKy650zN3j4vTUT+4HrJtIQFmivH/lKHrSDu5lve
dpMyQtmYX7Hu3ysVX6+bDmL1fKbsRQzCL1YlQaO59nmkk5nv0DQBn1X6xv2v
YT+IMh7M60fPDwgF3YKQvIF1z6wM+Ni8os7dpb7aMu1Wn6AS9Y8pPZ/1JKVb
6kDiwyjSEcLDlI/+GpIT+u+sFw5LTeWfNv4XZIrSRVuMFh91w3VV36x+5o+i
F37tUcEt+nXz1u9ueUUuC/lJDw/f7xbz+POP6Q6HF2QV2fmQz5MINUneXUqL
nn+baF1aGOFUVNX6R6TPo3naoOKLMMcvkFwXIOzQf44HAH36b39POf7mYhzs
CTNGQ/v4tlreRyZih8wJXOV706NtqnCrVV1oscdPZ4NlELeuqGvIiejbIPt3
vpXYoAUhmtcrLiUbq7OSZ3rsLqa0aRB77tLcW8JCZcJNtCwiGeZvlxDYTDKT
jMk6mf9OVB3pu3MSPDis5L/iHXlJE9BU7GfepryTc56UDvCywFxMq0yS+BX0
3sxKaHxSTCEZlXH+pSOHB2xLWRpX3WOQkGtbHB2rAl2Hd/7T43fvy46N0vo3
DPA+SQCjnup01oppLpt7dBsNiym8wgsx6/C4k2AlikS3FyU5A8NLA/eFsjU8
d7Nl3ALe8C3HdHqHSzU3fETPge2840kHhSzfOO/A3vCfkDDEoV0+ZdkJoIn7
F27LB5eJKSFV5hD7H2eQLjwvWH46BUMkfEEHwAgoASe6ik3j8C+XYW8aV85l
JalxgkIXNwkcfO/RW3gOL96znRpz7WIV8J6OJ6CCRqqMCh86GiPI434VZWd0
Zp85/7SEl7eSrpDzbSQ95j89CXjA9mMJ8O25ifh59Pi4CB7Xf0bt+hLjpkKu
Qb3+DAoUOl/XdiTfr+ek6B7jNl4FaJK6E3AvOfWpQ0UQ9FpANoYc4hKY29+A
H2ROEMXes6sTUSn8mBieurAO6PGxqdqAQVk4XLk6gLKxG/nBYq78+Sq7owcC
o5sEhsGW5Sp3F+cGXfuR3W8BdfffVE2CbdNykUfWNaJnLnIvk+0nabtzH/QV
LG6l8nyRiSPaz1Zkp/AZexrbOuzpyKz2VEpC8qogvSLzyM8P7iebqi40npLy
GkBRGOPjh/34bitpCXJi3/m+LMbPV/TM3RD5MtYBHzBHeO7Cok/Nrs6B9nTp
Vs0xLr6LYobF/KMZqdKH/adUp8JAsweUSxsgw/bk9xM+1fwrNfk9w+pixpWv
FYjqLnbxp7UXwChDEyHdEEpCxk0V38aso87/f92MnmnkdLMrdBiDPrwR4K1A
9jmLBygwOPeMPrYY7o51dJkqtpxW3AxB2g1VVjF+9y68VmNfBrhMkX++Q0VF
x6RODGyVUvyWiSVdJTZ21a6bShgkVH/UyvURALzeJnoXcqWQLOdO99tp4TOb
WBkCrO0YVcoEuQ/HC2OT+3xvr+MAYpQgnfm3ICHTaN868xaRRRxS4WojEIap
SMaPdNisPwFkOV96EafGT+uqgbrkXkJ3qXqZRHNb90cXlNxqCHX1cQI31z9M
rrWv+qYYihjWVtP7kLcCO1pGCBHk6rumcJ+QKjku7cLeMRh0TQnWrV93x28z
4Kdak2omHoT0vujTgp/4lrcz0CAIKMaQYtglLVZv7tF9731xyg/aNc1SUkH+
TQoXGndSi+tlG+egTFLuuhXTkcsV/Z3MTwY7Ij7+7cqarEqC8IB2SDQZtyxG
g+pta5Ai+zJH5DS558gCt7/Vuz7tjqT2eSz1fe6vDBJOiCdWpdNpR9OeZGwi
0O8nUvpxu/y3JyiIG+gsbzjzdNSeFZK2tYtmdI3fBjCRaaQV/JjC/AVlQKAk
To0abkjRrvl2qrr81XzECN45Mztjyv8iDdGY349SmQb9K3UwoyxhVEKxOa5S
n7NZOzSg0L/kgQZYgcjm6VmPa/TY4qJ588mduQ6WaQ/I8EQNyeKgYFyLWZ4Z
v/v2h53L+mEYps36rZfFdbw56W4Z4TO+8E3OFJorV3YVn0tqEF0pINzsgQ6L
S6M1eNg1yZYaaUVQ4VbrAIBSBwd1wTYWn01GRBjYDXPTmAVAjmbog0fo6sGv
YsptUp4GbYFJDDA7Ye/oAcrwQ+dE1SVXD/L3FheFb4XJcgLkprH6EZJTFupV
oENJP9GBUslqTpD8cA7W2nz6NyKx1wt4sjs5OZ5enjdcFuwlr9XV87d77C0f
TXM5y+XAEN8tn3gKpN2ohjE+sfbi87XZSUgfmgpSXEpMn0iINwChvG/64FnD
OaIgOYopuCVWPvtq6phxCJftKXw3EA7tGr0Z4NcnZqs9FdB9RsO2QhjfK+aA
SefsEqEiNr8Vd/MSBTrf/iEQ0vBCFAl/DRm0OsFCt46tSMKxwHxtaz6rPPim
Ab7WGTxddSV/nwilG1avKdMStx0TIgJOXKC6UiFWDLYj0LQDOqXN+kBwbSgu
+M7HwjJS36B1Ra3X8FJRpR/sd6r4J5szE27W2KsG3OKu2OxwH30s7hWMFfiD
MpuDjNW2PhlLcGmrWVWta+27gNKOPw6fk9VjQ9WeAvXg6g1h5uq5/p9qGwQY
1kR7j2rU7n28pslf6X6zJ1G7RRjEMwtDlmMx3JZM0pKh5HRJOOvJnEF/+2v9
DBw0rYe6H+nofO6bxQ+bR6otU9gBke9XNtuxHTfeYf+YSuX0HV25a6tRgVaL
sAC2PMbi031FKaBt0umLNYxOc/qcwoVnOenSsG41dCMy57KQgtJGMJot1Hap
+ORX2eS+0x/58UZNBd1RZEL6KtoWDYYSrsG0MviBA8ouAZW/tcTUeTviFSZP
9uRUpa429runm4P/0MTLyxdHWrvhaZSpbW0sBcku9FTesq/EV8D0wi5str9U
9iPZixvHj+w++uX6e6m6hsvhyFm1fyZjUWPg4GtUeesZQDUv4Ko48sJFEU90
EiYCB5UO/ZbCAdQsYNm9VtQspBnlvJripJqnXdkp8IrqBqG1z+WbCUwMFwPt
BPJEj8eUMIC4FyeOLAgwDlwov0HJMrUzSs/w+Yw7zEcQJeLQQr319s7fi32A
2PTbtMdkxwyS8lyo3wspRYzE7G/+fxdZVDauJEJHvgFZs4jpPmGR+SMglmUN
Mc8sz8zvvGAfmkiq39DCalehUTTsox6tKQ2QFCKmq/KC9QMEzHIF2xZ/7N67
vTDcjWIV2DKuZDYkbG6CRptJDT5K0+sJqYeZkB3d6MQ0XqZPTC+Wbnr4HR//
xzDCgymugX9lM+p6pAVPLvgd0qzT4B16Yf8ZgWwJ4FKqEqV7iCfCheXfGmPn
k2S5PbUhvMQWCMttPO/xXUbhKPNBV7DBEnhzCo+/kmSnmYJ+t6uBymkvJmVN
oPWi2uQp3Q49ZxJ9laTEr9rR+iEz6qM5/A5uY8SJKWafhjllI/Y8Y3QfU2Dp
mdDMQVtf5U3BKwqOEuU6ExCTdr+h6oUB4AHxXL9yr373RlqEOlaiOe1o5QVx
BFGm1NXZ6XRbGOESVSB60v8tGOxiZ2WKZilbo9FoDzSfzQe0RBXjCwWi8n/9
aoKrI7uNlnORFPCuwjEj3DtSAQ6EGBCQDqEH1H7uSCFjzVphi1DMKI1GprB1
F1Uo6p4VNswQb9qx23Y3Pl8F19eaGiVsG/HUiWPpm7P0CF+IwiBzp0uYZdgg
nOM9T01zFHDQU7iTP6oN+LUAz/Cu5sWawCpa3om0wZHdSNtFqRQhDUlVGKpY
hPvtTOspWfsjLCB6SuhZCmRk/hzVZSilq6J5A4qZEJq0Wc28dsV+LyOu7DGh
5YFTBhzE/o8nApux21fsjuFZpTpC6FStpu2RgTbrnQScuN6x7Gxtlh7pXkHK
n82Ldrppa8POphaezEyhLKaCXuvWwjpCfBw2oVfyZbqpbbGeIqsfXSU9g20r
iIfN1EVtk8q6p0htc3ff7B9KVN3jQnCWqe42g6omwHFBapzSDwVXClzT8cn9
vXhW8SWqxSN97vi6vJWQszR4NiT8HXt5QzvtS6U4pXBtkQiob454nbOs3El3
u4w6V7KcaHFBkzWd5ARUqx/Hbxx8F0KbLCXJ3ECvR4Pd7L0OT49UOr8LIsB2
MdQZX14sL7Ig4GRj83btyqLWIfZzZxxr41dHFtZhZUjdIc4gX0a2jzgxnmhL
72W9bUqK9gtv9jcYWcT+rmiYelkqfvET+u1uLIdXHBSNrlrjD7sfOkxEfNWP
o/bMJjch1CTfL2TBy5YuOvDZvDozDeAF9t9/1Z6EuYvZOfT/aX4E1bpIWTqm
QVPdaiPUYcexLgX6RuoeuGk6Fe5Fmv774GEtawr/YGeq9Nt8aFataPvv24zK
GXUMnfMYPUElXxoe6mlZFLdI5yhiM26yvYPR4w+eOeeZyYCiXTOrrQbu6Nuw
AMlgih60yrOG8jd7pV4J/7iGwd7b6YVmvAdGr+yBsLX1Y4cvjK+5uYoBS6LU
1tAgYf3sElNsRHdJpMXVStMCf5FAof5QG4NDciC92o1XCYwKAJDxSaEGCrDO
VNQLeahfrTRyzhupHN4/Gbc0ZMkZdImj7o6p+lm8yWgnGZ9/8xPiVPYdC5ix
DaepTJJhwRcGeWq8jXP69JWC9id+C3ioXs8ChHBMgBShaIO/Ie8B1MoUOUff
x8CnnRcwSHzZt2lv1MCzDKOgp9MDRT6OsNpU5fF7pnJ4nIIotVu8RlRzwZLo
GOYHaHbmRnr29VkI4BuBM9aHR/BL21nrXHuaArts7r0WlV+YxL0F+3VAoBV7
vwSU2pxSdcdAXCOMtVTKCiw36cDo6gcWncyy0d8WIYxIp24Bvk/0jnEK1JFz
nV21YEzYAq5ivfPY7+oseyvbF7GkWjDNlEWfY66VZ1l/FGs8iLR1oalG0b9q
lHrEO+UD/PMxMENzFtbsiWyJmLa2rwIG0I0jMM+Jrf41mDOkmuEFytFDjmfW
I3R7x2IPDIVA24jElqgjn1YRrE1OnCfbPXhEPwPlXlDpaiXAif+0mDoTYBsV
rVdUeeSJNBMrvgZJJwpoJJVMstXOenYJadqbr5/Nt73nKsTZpLx4T+LxpZO8
c2mRnGbRZNPr0GTI3CH1h+gKr3vfFQ7aqkNznvu6sAM8+8l8c9v04Lr/vOtH
hN3KvUQfAZKrAw5O89KZiznOmWfWGDQvL8XPEwD49lEQ3as6yg2t6kVw9gX0
Ix3jvz1vCinrkzSOEP9bQe6MDyqPSqJPwV52xn7nUt83jnZvfFvTc04gwHBz
Yndl5135HbclJJC/BPcWrxn/JeR9yiG37MUKM1Dbq30w+XrmMkZmtlavVQIZ
12/p/bbvZ0eqxCWibY0oz3GCMEuAODSliEeQF6In19EwqRC8J8jR8dP3Pl/6
zRWdNQ+OZdjK6D1SROJOL3V2czUQSkMXx5GJpmc829oLQsshUuAmqEOzYbdY
fJB+ug3n6SCMYbLCIqjaQ2ag/QMZk4tk4hCqIou4T1yKcfTqk7pKdJW9Bq0x
DFSZmnOkavSdJRRr2OMXpZqhgTyQCJRMfYWWY/Q4rpp9NZOlygK/EPWlTY0G
c37E+2TegUxBFwm5TDLd4GBdGFmvANNJlSU5mBcEU24k2BwRLE1yFJvVc/Qp
MMv1fwsiI6Rj47qrC566ZtWrPrmIKF9xblZPQPE2fdtS+XQTgdm4XopX484s
aA7tg/uHWp9TQrFKe6cq+yMjvxWNHXyBKXWEqqu/DAFLiPBeaZsQyZvFeNgR
L63+fx42KYjYEouZOyB447aB+cDOE4fbhmT5JoEdyN0z1tYBCVpKGyyPtDFG
KYkgOH90zuOLQhB/cBPmZZZhFmvsKt/ZD93guptwAA2atlIZ56jHpT+N6Es5
aDZb9WRnZhkdf5uNRslTqWODaPbEHCcqxKRb0ZCi5pmlNmXsbu/3nZKKyvZG
pvCGnwWHTL7qut6o8oM0O/+IoTHaBLFBwgbZC6yEoM8NrOALvHcSWOcVPrv9
sRRyjX10YrwYA00Q+JjFSN13uKdwAG37LtSM61HuzpT24oaXWBIRqIPHIgRH
rIupP2t9gGCHGNF9WFH1TNhWLiofR1ewB6rf1mJy6dlTHZ+SAVYvLpjHfuGB
xJm5uoI9PxNrHdtOwu4D+grBVVr7GOVoYKwfMlZelvimfrPygsWdxzO0eUSd
X++2LgvjbEwFkgpsF9Pc9H3D8qL7aGtMQzFEwkSpTlK+r4c3fWv4K1bjN3C/
suQU8WW/3BjNdp6GRODHjzgl9oH23zkE4tINeWrYGm6uP28xf4Ulv6sEvlCI
yVO4Dlnj2RprVI00J6wYlo8XRxCgqgk9tMTOflp7PY7y0UZxMsauo28cmLKy
ZP0t/DAcnNPeg/Nx1i9avTAdRp9pjHPUZVG3sPt3x2LeWvNw8McHew71MEIg
fcXzhn7EVi3FKwEQxAUu9yuW+kDacmoThimLI/ctqJn/z00BApMMdFGpFct6
+Uw153gYuBSTt5hspGSw6eXfXAIPCieeSnMkL+LchLuTpYbI2IldlBfb1CFh
kX+49yH00AQWbNyfwc+KcTa4o83uXnDXbLAyIPmPUwOjzY31IsZZFlMLvazv
J1v1Wy6qgVxKFFUi4qLLahsdrgejqS3beeyqxjnfc0XQyA40S4AOljTEEnao
SsKSx5Oo8mzZQ7D2HBlXy9YEiedHmqtnBJVV6tfisiYMS7ZHOZeoD1ho6TN7
vQZiEaV3fJvsAk5avve7bJ41VTIuFDqe2o3I3A99Bzu9kaen5bqKMFfPzn92
TmO8QCmVkqNFBnx+c/9OrL/ZnO5L9Mta4rmryTKU8PhFVJXdB7b748pr7w8e
2pF0SRnOsoUSMn6z67qpmmayN5CFEmbVkGVeeejPJ0tUNH0luR337c6Qg8P1
POvneZs7GxTxeC0KepciCUipkM2uluqQKh1A7ma1XV4qElaO+yJ1qe5tjkcM
5ccWBstYP4zuP5bHCKIG8NaKRH9/nHODiW+ifceaX1wUBD4Z8dKfWVeD48pG
zPl+ClPX2MFl/F1V5ZVQx0DLqyUXbATZduJuhLNWgRRntxyGqucLVD878C/9
5Nu2ydT66PTyQlzpp0OWAbLjGw3TUexR6abZo5EsqIhQzKy11tT3Nu73pb4o
NkCJpCVJRDL+X7cRS6GkCgBCMeVl2unbQpdZOgBJyExO6WLn39UuccKr0Rrl
kvcDESMwpdhMjzgqJUfZozZ0rr34Lvgnl/qxCsW3ESkr23trpZgIyCcyHsbn
G5RtyCcwQ71sN5pjntIyGIMfjmS3oP16Bihb8ay5QKZpKcaMoSMeOErKjeUR
oviS+j45NDqhaIMnfQ5ocZ6Pb2fqL3WGw7lpe+RBxT46rT+5q9vwN7RLfwOl
3UzSvscHotGXnX7JDYsimoHrhE/LCAQl3+c1HL432WlFGujsk9yhiKZl0k4r
SnwQRQiKhQ8/pgKDbCldDX4SrMnqV5OAUE9OGJf/rSCeV7skxyYKVDvDBUt1
C30WGOG1s23hK8/j37erQOPcXVrq3CuEbSVG/hXFUETFKkg6YOejA3C9l+d0
YeJvVEFvdGVdr0VnQVsYT3emE3+IMXjTyw2UOIYZvhekZxUbyIKaqSvgu+xK
FUUke5o3dpecKdJ0gd1h6j8/yE5j3D0grTOrDmcd/8xa1Ns7OwfN4fjLNmgP
LCapnEHdAfB9fgWXcy+IfrRBzAR5lT2KVzcqmm6sEaFjhsUyUyM3sYljy65m
JrA0o1bTd1LgwpVBmh2lsrMRhu5rYZZghqXdiH1uIBMHdTs+dUJ6DymkMgr6
56TXrkuG/41yEWn1H8b1xSMUeNXpXf+ZB7DgUIaUqCP8B13XeLc8OBKsxuem
qMo+oK1XgwjCzPvmppcT0GgOTy0lHEt+BGKd4uNekfo+vCSa7Vg3TzHRIQIo
FuU8ZPXjSNoo/xVLtxCKImB9/jq5lcmhU9zvK54rA9iDXnvmg2J8piEOzmnc
KZDdS2EA47XusjqvTrACqXNhbWqVCT3kj4Uz5LMflK+eXTwv4cYc5EvDw3Rq
sfzmfh9oK0T60oOda0re1djXpAnjvJAoL6G7f+Zzms76oUiJaqJKQLooUTpn
G1VPZ7k9iMt287YNZrqDWXJdd2N8a0GsDact/CWqrzlSG0cA9o1yo7QqAGbU
FdbIt0hGMGPiXmxY6vIMJAby5yM2lEygEq9QR8CZoGXsFm9JT9lzMyYQaEEE
0+u574Fi/U7kA9qXzdUvugTTEZ5G2fW/BIbyDQYF0DOht7jdy4MCmd6uMcnq
dknDNpR6qPcwEx81VVzB92BIzRnQfFMd+Z/mcrstrp467Y2lFyPumBgiDb++
v2BAjXAfEAKdvZJJoS7e37YTjD0YQxmZNgQD3p1kTN0/ai79DNfM3X2FLoWw
o1u5OClO3fTtTFZ8IO+LEB0qak7QBF0+8vwKVcCog6sb5WKw9wbARJLwKzzC
jUHuzx0Rn5SjWQXZxUt6GrmpTahIBhxaObe+uFNJnwWF6OGzQb0wFHo83aRj
3CJftQYZp6WRE/7YFzI6VbAy1sMnk9Zv/KT5lk0QFJBcVd+gHZj5GpNUkl3/
ilWLhzd9ASUcvp5/eqra8Rzbu8flzV9xVE+BRNIiP1beDDLFwDzgdcL38lzg
vmxQFngZ7L0cdT9RY4pcphYqa1nj2qwemNCkuBJEh9BhSNdtj00qvcAWDbk9
7intNuzogSG2eDs1b8B/RlzjK0CeSbphh0YaXQGBrw0jyi7FPCsXdaHXpN6q
24bY71xHqJcFYDlvWdyGRVwyORq/1y1f8JtvixcL4zhX4PgL6HizWcEv3Byu
hhxCFUxmnjSykF9Lgo5xfEQyUlFlKRxNnWyZZaC7HpHL+oeO6uqJuzv6yAWd
PK3CAHs2xQX83HkVmM3o5woFvTfZWL1HhQlKUeiHbfJWqUNKMYMIuZi+7k4G
69vihm2lkm3Rxp8MLn47crobt8nawVVJ7EgQSKCCrfzF1SOXTw64YaQ0Qv43
ywgLMwstOPy1aAlzFMmLkvEKcZiv4bl5PSseb3Ab8ugZOi/DzebSDw0jSZUu
/PHUoiGAEjvD2/pENg7tMaLbL/In2EaJIdTBYo6cb4OVc01qx5wQt4CBl/pv
aPwEVoKxQGDEBjpZYODAfmCIH68QM52iHFGAEG0Uu72W7nqEgNxoicJOpVYB
qrcoU+bvHrRMMZJ/JNEzR3gs5/7G264/9HsLLfbDF78JJ1fBqJgbZI0m0ygP
WJrNfxslGIWIATl7Qd+08mVSvonpfxUq37FHBk3vlLwvbbEZW0tscxfogJ/j
n1sqZFs4OMG99ibYLx/WAqg4FY7Kv0oMOVX6w1cFaA1qPam9vd1RDMpoJ7e0
uztTwvoHbqaciSmlalMRpmIKluOx62f+0W9bZHFXxAnk1+y/E9ghiT0YCk4m
p8+815Gq0ypaQJuGCRtjn8hGxc2+cTEvJcMSUGIlZbUWSQzGIH0bv28xYLR6
YllXU3fXIH36qGoesq87RuIbQiCKvwU9CzihvXQqcW2niVzU6+mWlVtSn4h9
BwLWl4eu5gMpd+iBeu5nc16hCw1O+yQ6GotDa/ZavsoCHIgracYfBVEl3gkm
CPvaIiuz7cvL0F/+xtYFEhAZPTAEtxV4UNznHG/fa3fEPZ+1ToBf4YsFT4ZA
6NRL7zxU+8Snr2QSMXXmAgChChBQ8jILkYclD1/GqyCTkpjnmgmAnr3jVlAq
EGCVOh4vqzNSRb3dtqqg9LT9los+eOKpGwGCDh5jmLvPTvYPCx0hAO6Q+jJo
DZ8UdWA1QC/FeOUPd3T282U5lYbGH/7lE8y387epZVR9iALq8FDwJU9/ThVA
Nqvvpwpo00RXEC6oGXXpAGWy6o00NJ7hHPr3+vopSfRa2z+XDFsLozqiVpXw
689LRCBBzC98hdV+qpwFijAwab7n+PSvoSan3XIYporLbGS6HzhShrAgoY1C
jQ539v5fEAgDfl8VauhW0IENrLu4S4G1dRnplBjU2IQZEAVFBgSc7IPsJ/Up
Y+0/abGMWS72MVuqcLPL0u60tCGZxAmhT2/GgPVMsHgDsngrwKUH2vwa/GaH
6+9M/aLNKAWwf3afGFUnwcuN2jJfL6KNKOD8yeXNtDCvOZqmI6I7HWrysner
NEsp181Iu3dMpZQD1auf7EBMMWdfd/PDv/UOJOYibABQOXsUw6lSaKmVgC7T
v/IwX1epJm+KH7DCBPU2Bg+J8DxU0sDjqvBgSEVfik79UEYfIDsciVfRI2H7
hqAwCNktvreUWeoLHlRC4pCMoHOWvF36UZsZc+9RY0P61plJiCBZVHXUZlsf
6mIcu3cXwcUQOavm3xWJ3J1hfCNyC3uxd1QNXk8pHQK2rJD6S8UyvpzndqCo
8lhUe5t5dXg6t7v1w7Bhhmy8ItYBm/kiYic7JNIqfkurCOXYSW4jkZ2fSX5V
TbvjUotDureB9n9GsxTNda3eb2xnQ4tEk9PbPcMuspE36bWorvzRXGuFgndV
sZYPfOIiTzdKZXgWW/L6kslkryz7TdJiBhiA/XZqIZVtucfvjmGnxGCIDdhE
Yhk2gSOXV88/YBSeGwsGYoNSOreVGjr9zUUti/qbeuZT9EURrL9xZxcgpAz7
1bTXJ3zeEV64gh6MBiy2ds/WGFhzadKod3Y71N2eEO4DdTk8La+Ut6AbbXW1
jJ7remLWpupZR8p4TGSnkKSmEutiAVxhEV/8cQjAzuFyZFbsK7d2gD5kMj2o
xZPIatplcDGpspnDmoertyxQBZIcgl85yx8rdvexXr/JleIXQi7JRpWwoyJp
LzTWphEe53Q7D49dQTuFe7DupFJP9qrqtkYFL/k9Ohx2onIMHMsUFt/MVIiI
5IKNo5CHLDUOLhByYFRMkjODqQ8e6SJVLxuS+NmoB06KZ+gCHjgEfQK7UDCw
fsY+56Y+dCiwAHEcgAKB9t7Ia18xmc18oF9Joqs5dsVt1vha2BdtQPBXSkKe
BnR/G9EeT2LxnSpXAJ3rBzTNQrC9dMYFEgA4wYFs0utflE0QcUNt3EMsE0Oo
58JF2K9ftr6xN2aFf5lHK6q9GiekN+AR2ZlnR+A/xekldCAL/0d8UomBwYrN
3rXLLqDpgAPFjdmGT2ybmcrdCO/ZMEnMZj84cH3mOZUpv87LQfpgI57Tggt7
rcm950wIc5X0zSPiXQsp9acYSbhURYrZNoVzdcUUjmSSBbLPfq5B4M1NMCAb
2dlnOYtKLOH+neV1tpA9gO3LdZSA15EmF2URNx3+hP4gWMtzOSyJR5HJahOd
UIkC94NFcQrC7lkBt+Qo3WJjbj3vufJ6iTl1QB7Q8l3YTcNiGwpRhe3mNyAj
u2f11SvHnZH7cXxKYwvKxjIuLfh9GtI2BnbsrJXhyzIs8ts4/2QF61F5uJNr
BvxaJWT9ejRR1v/R7WEeiGi1vuAZKUzQYE3nZcEiEAKeISsnTjA0ZPi68kAI
N/2tc9pDgJH8vri11qvly6qLWAxySXm0kzOh3JzQtzisrSxkVl4d1Y7U4Ek8
R+VtNoT++fgtBRdMw50Dz3e6IhDTJ/voHO2X3/tiwDd4MG43RfUARO2b0m8a
Wy6qr7O1gH38Y9cf3/FhguyaJM3p0GxVV4QLjlIwvHBqPicLULT8spb+/909
OL+4TCPdiwY6rqeZnz0MuiMGpjnJZ1MnqiKPkMSuB18pTPwd7bOdg0wVrGYV
sDoIq2tav3lS8KvreQGrjzF4GkCUjYhJQyVAvbK1Eh8mJ+2R3T1y2VHGJ/jg
umAeSnUbRrlScoVlr2VqFzXH+HYShONeKmgIx1EBqIdnmVrL0xjY6bmv1yo2
hO55REKow/k2eH35fHW1RxsX2HtlsWpEvSeRU/NL5nynY8G4kffXxa5KmgDa
8sCD0ieAYKXUB69kYMGJjpowmaL3hUtsRSx+4RHkJuzWyQoQDQumpBZr0+rg
+4GWKnfg96M5AYDCZX0eaEBTKGAmR6YdJnjyqno0tskQFASKNz4XsRvKNbu7
sToBEGygsKDQG3pVXbDUOeme2eUChOuhmqSfa+89gckVZ1Ai99msbSX2Kl0A
O8KvrQ1icr5e1PAPnKm6nMop5XNTAgVHR8xfj/XOFcCclHcFUzlRqh74hU92
hePpkaxQ8+oZPrMMCTI/r+ajMxdZzUCO0KCDk32+8WBIf17JjGloXytHFRdu
7ukQl7oJiBrawavec3aHBhD/R9RuGeQv/f66H9Fpdw77Olm+ntvKuicRgKrZ
uSdxOPukUQkywv1sTwRg986oKGDMh+wiPnywimZfogpawiHV/YfkgLOOY495
l+57TJidekNJIbicnZvcgJXrYdc1B6QYsGYfZBWEYjf+6lqxt4tNawMDe4v3
si8ch0+TiM8PoQOyzNDAqWWQ854jttWM36udXTMFOOM13Gp6UsIV73Ew7S0x
Y9AZg/tT3OojKqTlWRcLMEY0ooIAHbhA8TDl1kWaJRJC1VuZJZkBWjvr5lwQ
mxonYMHDqhmtnsCPPN5VIOuBs9S8KOBwl+ngmXwAhB62MM6J0pLfjE3QA/Z0
dG/gq4SovsB2OSXXk3MHPA+bipAieUHx/PhNPdxIQRehD/PoL2rePPddWNAD
sVWmt9QrQdRoTVTHRBUcK364UfAawtu402h3ulAf60KLd5BL1J8IbT8iWro+
Ggulpi0duAlUfrLZTkiV8kukF2vjV1m1hHiRiBjSlTyODcXtpPJwpbTXWivT
UOEdqDdJW33fQO2wQorwhFCKcG9NIZpgZ1a1l/0kVFmoWCED1BZA5wQROoOg
MCrk+zhzibHyxmmqU38KILDbddPTbdHrw+cnsEGo5UVfZek34E0Xvn5WySXy
CWB+274ocJO3B/5e+OZrbQAeQq7aTnpvYJgrZik9qGUGKlhoFcJTCbd/dq7F
AuWBDBKJ/lWGl8pxQVQ+BfxZX5VkbSrvdzcgHRyfmMghrSUF8A3Iw0gAaOfy
woCbMsPMCdBp70vxmcc0qoBChY3RJm50E1HI/mowJRRh0XWL4C3Fz9AnkwvK
oWG2hdT+lAbcy1TgEarm7wx1xOmK/nB/jneiwF0KEHv1sFMyHeJPaboLIsT1
N5SNAWlUV003P0e9q5iZk9h3prqJf/vBvRHd5YQNj4RVD5u+v7pJOheQuiOg
tNa+rHgQ5LS6JQLFwIduYxl6IZCNsANo3MQGI8y6URqYTSW6GX4HEd7yuDZR
jdORzlPQTUYm4X1q1iNRkYQF9rU516ltrmIY8pVnuM+5LQluAxelCq1hC2mA
rtxA6aioTESDye2sZhBDi67hHMboTrtE8GnV+Dqn81RkiSEgNuyyMF6uJTkJ
pnQ9Ehhj5S9jmmmemv1aRHLsCri6s6c3t5RNWB5JMZ497z88AHJ44po6Pqs9
I6mvM1LBH23zGGYSyL3/t2M/bCyqvWNKhhQU+JaQsuM+SBmRHYbUu7a9bPUc
A1vXLq32wb6LkyBLSE8i8X6zjCxuOYxTruYcn6A39vkT/NCLv7g8vqC39w5o
qFmSE4SpyIKjiNmVrfYwXcSdN8MtAQjxpizfpmky4yBi7Zbd5E2cZ5b8nypE
2CKX8/hgiFXCBB/ogDg2gsdufl62/nm2G84R3+VK60xVnJU+vGbLYUPqDdE/
zBE0xk4HgiY3tngddPaLDz7Yq5gGpJlnw4s6zgQIU+M53jKTNMubK/UYga+t
70e9Y9JKT6myg3FogVEGNMQq2kxFz0pAmcff/UUTCQuC0II44NZRmOhhdD3W
WOM1XszZMqREggC1fdWs09iqgOB6QYIe/XeSdTW8ye8R/25YM1cy8np+T0KD
W2LANiOhaekMEqSDrnVOhopqO1tt+J5RFD3Ll/Fepm3Yi5+06QUehERkvciN
wjzMelIXVuFo84oYRPUUH5KfWCbcvqbAaT3JiDsIGn4Hi3VgWUqOLcCXgPnr
HDAeOtqtmpU2OJ5Q/se9OOpCWx/Kl2Nrg/BmCfgPfWvTtwMedXzGQPxt9d21
30vdOj9D5sq5vOXl1XlMzv6SIf5nfBZznW1abSZMYtFD2GqvTmnE0A8GWb8+
97Z+ECw3pDVA0DT3y/jZuE63yjY6Au8/dXMinOl9uLn7QZGosuFoZNZdR16c
gP5NKrEHNnCkWI6YJZUVPziZ5Cr6PK2wHXpluCfZ4rxSHY8PZTrXt25NlB8x
W7NNEMoyfWIoWLLLRlmRMEJgHD6akUL2+/e7zitJ4u+nuQ/Ma9ieyR1RuGtm
chdCGbvHHO+hkcOfP9uGe+fdSfpQsTg6nsY9hLt0HWZ9jViFopGM9iyhEbNj
wvxbNEuav/IkUYQRYmKZeCBPQT50/uwOcOEQXDe7QreH1pt0Rq48Vzv6qIpb
btDDGQzenfodC6Qc/sSbIvJh+V3k0F8mmgIBxu5J/d39KKCJESdlxnQtJGQf
F8P9zZeeFmmjgTWE2LXDzW7Vg47tLZGxP7/4H0dCDsReNY3bR4yWluIcmUvs
SbWrMHEhnDlRE9Itf23TT0IgkK+/5WNTal+EHhY5XrAg3nIugxP4VYSnVG5P
HKlTyu2EPT+iMUapEvmqxm4pYGEBCBTFBqtlwUquXyrNdTuRfuGf7F4jq/NH
2KyVC0RT1UOqUMZQTdNcpEbfK3SsBAhkOM6gv2lu+9Nzt4NtWu+UkX1SXE65
n6f4iXQ6p14+k4KPWukbNxrqWDIHBfPUgnd5f0dwDlyH3ChaNLHtEmsR//qm
8xedNpICmDhn2oczAsUSmO8hPFc0sJBamLuLSG2YF2sei+R7gl4z8SRmNKbq
b9a9HekKXD66jEa6eWH6pugGisROsl9Nd50UyMjKXSQ9e3yeM4wRFRnem1H5
N4YprVTnpj3wFN4AXo6V2T6O5IlGe9dPdJel3xlP3NCK4W3p0kmFvhBLbDp/
TJuYnZLMmFgPlckMLWw6LUcywwwq2tNqMmWbd51Xzzw+46uPXmj9FrLC+mrj
oYFg6RaXBH3VIzdwlqKRYuUMQuj4Kt29a+tVRtuwEib6PfNT3tPmbFPVdwXK
Bvn7qPndHQ4B9+rlDMD/JOIQBNWhBIxRGrQdbMbGUtxYWfPG8ksolWyeRR6F
hk/Q+oE61htE4MHbZapDPhMh3FhkWxuJ+0lwhoyOTWK7T/Q0Atwf6J0LCJCI
O7auDsHslapq/nPjaKc6hGthG2P/c6X4NDLMMjozJfBlaXrp+OIMuSNTateF
+fWtdrSQiZtf4+lKalW/k4bsh+iV+NVAEz92n3MF95ascEr5X/Yd6+376JSe
qmt16fBJs0mcMZZv6zw7mn29vt6xiIioPKOMlISUdwRokwg6MsqLCSyV81cU
yUHX3NAGSemZ1A8l/JbWIWpO4FeT9flhEvpilH2JXJMufu0QiXzrxHhAb4fO
OWEk4A9iXgMVN76S2DVNn60nON+WsZQf4eClFYaep8DvvQ/DNNDCNPLFqOSt
DxMfAEQPngtAkyfoSmBZf9pXrxr/BDDeNAokNbFEJXKYyZrBo1qYETQxkDFe
hrO9rJa3h05vQoGv5YOoKzqrRA4FDqg854v6WsPJPTQTtNYHnYG/CFKemqqu
ag3gIdUrgPq6Rq4WsxSAbP0JJDo/HDD+3g7jxEhL8GuSEh8StiFk+5UQoh14
KkuaGQw9ZbOE3n3E6MrgYe07IO6JjqhoXfMlFYdFvxlRyheOX4NP2STkBSFk
gySL0ZzBCkX/BwQdLFEEUKV4qi8PuIyPC7T+Cn6v5VWVSzeVChKMxI8gxuj3
xjmu4f8g2l+XOomLVscXpdBHqCeioYvagcZO57CAPVBlFtdyYzZcxfbsAmq4
Ur7sH4A8oTuzalnIcxfXY3sXNvvkK1wA8z7FmkMh1+E3HSEZ/Z/Z4V22xjuA
fhtrUCv8cyxo9sq2/xDlupn++MPQpowdruJ7wNA2X05uA7u53lcriqdJW61i
+TjFRqO+tZEw4wJXof+YSI/eIS8BQDsyxqTdIOrkSvLFYXuywtJFjGVmvz5w
h/vOu5MHNXfmW8PyZaavvfBGfywERBi+gZUZf8D3hgZkwWmXWGgA77Kv+l8z
x6syXTKRcY3J4o12G1p3IQnvQHCL0+bOPcxqiCByZ05RMIFGzGWXli6A9iHc
jZteXQpfMhKgwlD12IMWDc+UKevrrmKuI4HV2L6OZ8KqUf6IyWqUuhHS9wW0
ANCM8Cuxre2aV3fpFO9rIvrQNCceYjg5yyGHcMMfjP5YsA1Km9ZhwjIbrCgz
1YbbX3WmUt+0OJaAmYZVPWVxwchfECcFfoSbLBM2eJMr/uV4TLP92zgw2UDY
FdKJmoVThm8kFvIWh+oIhxTQ9b5FyfvKuqH1sc4bnDCBJ/05oJQ8zol23hkR
S/5IavqbkUQTbPXs+s9cthwQIKtZFefUmdTVJcPZb8hs3v+Wx8G0UY9mZUrx
3CMqx4R0mdIC3SQzEyBPIkCa0/mqGISdPIi69gYaLEmExRmSpsnvE1zyG4uF
1pVi2AC8bEByN74ZYBwqtBhQAfEf47NJBsQukY74MIxxrsaR01e7vX18SVgb
skp7HLouIoAsCCE+MUzlmfTwY8znyiix49/KeAx0rKWjriGecO42lrM9iVL4
rgajH+qdTQULvK3MkHZZjQvzgMmaPxRl0gVWO2WxhtEQF9SkR74jf/EBdqxI
l7WZe5AWoR3vBUBPvQo0a0bsf9JD0rsJYAXHooTpIO9tmNCLA4UJJVDwImB3
hL40Awl+CpoZ0O94oahW66EeCe4bazb5VwCiDph7nUPds7ZeKxY3+dL+xtNt
wLF3Dhj1ZxiJb691Nq/opj+coK4jMLYD9OnbM41nTQ5NJuF1i9je1wuu5+yK
gJ0FmCVlP0t+LUYU3s5shKACk/dA17zLGlrLPMEX1dWWIMvtVjEPaQA10+KB
stDKDpHI04Wim0ueJoVsyTyyuF7U4UkbDvU4S/qY8Wy19Dp1HWfxlcgf3n34
5cI/sgBRXoRY9d51Y15nEUOPqVcDQPlsjX2JX/i+gShBfJlD3efppnkDNPJC
uduAoiG7qLcGlwfCDc/vZl0pmkogLtC5Aj1YiDvPcuK0ZIGOCOZnxxd3yYjp
RLzzz/N+nI/SUHmadrXLERLZGq5VxQmNSCqaAjsK4XgxhsbJZthlQr6+fo2b
DARR44w5LyCip1Ur2em7ZTmzItVyQsJsBSloBG9u10r6VFMB64aZ12tBat4Y
jVlpUG78t2FwG+T9IfTR1rVWq/fZSE0XkmpVOIr9sdZ/tY1DkT9SD4ue1JVj
x4qYulMqrdKKSUQoTH0WEnZVy83u/eNUEu16LrgtIfT6Z2ASAD8sG0He1+lH
/tvwy86VHP8i5HDzPd2b86pgI9M77EpgriRBM+8/ytt3R/hwqNE6jod2qBRS
zyByAixpCGnXeCD71J1J7d8OPkt5yBsse3mSF0jfqhZCu3cMu0dcgNRt3AvE
JyLbfdAwdSEUe7sN9EgnQUnBMblKARUgq6MvKgBdxU0jOMbCc1AJW8/UYS3D
pw1ZGVvqSc8PYHmWBJCda6mjF/EH7UFkesBELDqUEX1hKaNi4YZKcV5fu46o
d8EPq8t08U77suywPWhKrtnorpAzbKwl/Lc0DwU+SRgEFtcQA3uHIFRkmpYe
yT4qf0SAMvlTFGbf1Qb2eemDpMfCfzsSyR1d0fiAN7zzZ+2eDq7StT3kgb0J
98DG0GOFuCWrt9eWOd4PCMZQAuhXKZogMysEyfJIhoOR1hLpQo6o8hcbpJmN
z4u8lbuKAqqLSsAbBJpNfj8kNR8+8Fkc1RVWCnYK+6snzcJRb+pi/d8ctuOA
apJ7CkpBOD90NS8pubZzUm/dgiqqRs4ELrcuXo3WcrNTVv+QRH/AByuxFX1G
HpF4DjTvmDLMzNAVFISLfYT0paiUXdqkZtmJJB1To280+PTwASLjSJzobpGj
Q33RyPYULNqGSARcSJMf+yX3Rb6goOBY1zHPJuDhL1g5S8y8HIb5mDXGnMAf
8PTlU2m48RLbQWuc/Be+v9xKNIJeVCZRfb8lFZt2O1rjqFJa5jAz/2fWDrn0
i8p5gIU+K5HfQHXdxW+pS4EF6UbPQcV8EPGJPWLvMve5TeV1sQhhd80AesQc
4bjhVU0WJa5Resr1vgwT+A8PlYQY7qg3xauGAQ2TwEzQOvvPuYueaHlUuNlN
qVWT4YgHiEyoCrvJyoTiuPOGNEuC3Ix3Pzf3qjLdC0rAMF7H0vomY7RqVs2F
q2H59xHlNwyJ0urw6idheImqsiRzLsC8eU66UX+v4sX1B5Atj9sB6vY72X36
OLFJYOqV/6XIDLenxM7t+EoFAoUoRq4q5JgcLpDcwgB7ENQX1IxEkBEantYC
aLnQ91I2PCKXnRLxNQEbLbXdnw86a1fZvo8YXENFqkrn+37GMTepVSl9oO+x
hB7CAf3zv9X978gIqP6i1LR8qWAdqaWPu0fNvXRW31CwZzMQvpgMqd/5WmWC
Bmg7ySnLCjMl4eZ8T/xRxemWUYFNZXfBYu9RQChtarqd1frvxmDla2/QyrIv
n3EmnYAVnJeiBDMGxs2RoLMBFt+wfGOq8yj/9Gsevkh3PjUZdVmeu2Vq3Bv9
1S2zyXgE4vxHy00S04Bu4z1zz9U2Pwi9znIFbnBSIYiXLAhm70QkIvpuSxcG
7foZzmjvYCO1DlQMLmO7SUvSXa/b3KFoRzvPeY14e3iAXFqQXx0c8Eor+qIT
nGCTTqOaJQups5M1ulrdx1OCwsi+jFxrlf33xtphI3qUmYqQJZ7753n99k1W
/f8wy2ITuloywgwOs0u4dhOQwvxKGCZhyW/gyxb5KWKcMhblEnGoCQ3dFjd4
/2WlmTCTjIK7JIUIEW2XGoM5qUQhlVVAz6nE/bM0jjr+Y5GLBF0Z/ULIVl7R
Tmc9i2vio4+M3bgyRjY4AUJDv8q83HDaJwmOzoOwQhaWiJOXSNKPyG9Tkzu3
gQY3Mqkh6MmnOJ58gt4zdEKxXfmkNaf4hMqTLS3/vU2iS7Hi9J4NYQmCsdd/
/+TY3lNWQGARb8y2de0MQ4npFtYEYCRxxxT7XRkaHlUOa+Y6hXY9MagN1iZx
eFGr93YILAOscBzaKHVIMhmoBBsWQP7Yb8APFM+4kND4OjznLxvn5u7wQ3eb
cTlsDsGpUCu149h3X4EdnbT4StTBz1Pi/GvG0on8/+9KcUMg5xqqqMCcCBGE
ll1nKYCvognDtDCLkFzVZX8RdEPqeiwlxEN3T6/BJaOM8JIXEZlRDj1FrU/9
F0OHGmEZW6ltRF86cgu/sFQgXXB8tVDp8f/ZKDtjAoNpIu9gizf/E8GFuj6A
/XtuXbfx90tt7eG/pQPnCCWSKFa+tpmCtmHwpshkk3mTrX63VsUtKqtIU8II
280aK9cf7gMVlCPxjHkn5OLBY+ELu9jmr+NBX28BQafDoI/qjqe2aQN7FMso
YI7K+0rZV8CGMOxyVEa62mdRohIHUWQ8QtdrNdcsTOzB5/Xhr1aOuIn/Ej9p
cOsXvv3wrk1SXVSWc8DEyRrbeUImKU+cpd8124EepUU7gB0XV0ucXlBTWyVd
ZG54kL1Qk/cOT+lQuK93vBKTtazHcBGv1M9lQ9ZI045NRCvb1pxQ4cU8Ofz0
F+JqUlLWftnmKdWrlMtACSX9fZO0zbQNzaImu04uBUeBNNgDoqp9RbfNDhe3
oaaTdCdr4piW77sbBhZvosg1UG82GDyg8RzWX3y1Pm0diqeOTvQ8iW1K4ndF
Xbu08XrnLT2C8wrXBKgh83XjIorBYDwdKnNh8tI6hDUDwedeJBwn7itv6t3B
sMdGnT0cFJpUitSXJTs0XwyPOJFf8P2xe7OSEEsFPHYu9LyRcYM1zQxhTf7x
XEKV+/x4t1o2yH/JC+0fCxGfTy/Mq1GS5Yef2mucZtewu+itCDsPi2HPopk1
rIzc1qGHNbNoEn1aCiTiYAt5HVkU09Dsp/7uRzs9yw5QGb0jyMOgLlXgPY91
lhBIRztq1IvEvW7oX7HwtHA/pITGY02iBlC4Z/NglZtM2AETlULOtJrlMihh
8cog3y0V1d/UMaZj6XlU7dYN1XA6HvscAuhRwCOC2VPAzfrk5xAtQr8yRlf7
s3UIUtj2tzmlqtNJW4nYuW5MRcUqag2PXMg3k8YQIN8E3Es6Hwg4ZP51fWyu
3zN/KmegdWQdacGvofRJSrLmkPL8CuOKqV0aK+k0EEvB7+fTX05GpKafuMRx
SDD+0iJ4DWlw5LQF/1r1RB3P+hyXQvlsWjXXrOHAmQFHYnave3VBOz/foAKm
0MHDcnjlNzVG0l8M526q/LMc8nWG15u+JpdYpoL0WktV4NKjzb4K+Hl5140l
3yLqyZhlDWjCuwrP4yCkEzDdcUhSKjRyF9zUPQ6QWlf79zGCTpxY8GTvXvSm
hbjoyZJO+ByGXt1IYrGQtrTmXpxN+nxQlhTJFqoZ1JShu7c4TSQAK8+U6v8g
S4VX3OREaL7LMcSxe2xEG0mD0cHUrB2onVMjzYeKXBoBIk99+YalLpTMFy8f
rkdD4Ifwf7iCZ6ksPvOynBvDv7wveNBcCCk+Lc6oNbwztANEbG90UyAGnEBL
Py6ISqvG0eJmNvn35qKQmRfZewMsSUuNO2Jzk6SxZpRdwtSqBsj+G1NefASn
NVjSdFUNat/VqjV/bGbovaDN5268yqAPpR+QGUoO4mkrnV+G+qcawAhJoq8u
mIrW2sQyXE3AmSg74slKs0REkOszQbaikZkuIoGgVkFlxCbbLrYgSPe9aoj5
I3UxuM1w7d86ST5m+fj/jspw6tKV6kraBp9YZBX9xEIdAJsoKtwqLtYcUPLU
/bYYY9kbI8mLPyd8oUxoep03NQMlKBA1OltTmCghhY3UF9jOW4PhNYiPjJwl
gvM/h3eA6Gghq5R3wuhhN+Vx+MX4QoyeewnOKzw0tjMFZ7EimPmDZiNNpeVD
V7xPJywBtbYp9n+EF6QqYkobzfZWBJ80QceIcSw2P8iWXSFf/3DQ6FLIFcGS
mxXEyILZq8uB+1RzNrP+Hp/nsmWCKbXEbCxzTV9abwudXTg9nw/uxkJ6It70
JPogF0vbpvYn8Hq1tko2ldPleQwBNw7rJiv4obU1Nw2unL+PLFOQgUfvpBGo
PbF42T9F3FIGi+Q7/FURgLEngnqjQQTtuqKpfoxQ+dn7+1+AVU7PNYD1VwKb
vyyfW4/wXGGaPrznq4JMhJPdLuOhO6Z+HbsaftwCRipAJOWXEhU3OTDOOWhC
0HF1r6RjsVLYFrILWUAyHa6+KUKAaWAGunY4vzMeVX6F4khJ8JItHhV+xglf
4dnlHrsh7dqLK5IqtHXkT45fr8fy6wv+Bxh3N0gUkj8Rb06hy0gmu54ZQLp0
G59dnGM1izg95tbggPY+2Rx+k9exvy0QZCQo4a2T8AqRZmOwGvYnt4Bt97HQ
I5V7Yvptd105iGLTdDH/72X4liwv7FFNMDtBDWpgtnNV9sr4g6R0B3vNuhjb
CPYxAlkrZM3YH/Ex33+6TS5AjPcy+Jn7QoYxtmSOzOJenIYR+kM7DuIQn3Zx
r/U60ywc7SAHosDxn9uccEursYrQ8E/nw10LZ1O1dGyaL4UYfnZu4s4U6bGS
dqnnzDppkIGhq3QAxkxTkI95LdgkeC0JcFtVK0EcaUVX+KfSWDb3ZdHuhhYc
2GtWTnhgl7bJzACK5HPe0RqP8xJAEf/Z+If1HoJF+gWyBJzZyGzM1HS81/sp
UO3ea9hFSPoMwjt5dqG/ik/FqZZek0e7zskd59YBdLpSUY5HIVNzSyS+OaH1
TDE2RZ2P7JMsuKc6WELZanFyv3hs31Q1rUzEEN51tKAl0T5ujZUEI2cSiSUF
nIKUVeKCGHczlXGyK/aeKsRhrOwu0vsIMNJ7uT/5z14G7digqd15uqmViu4s
dmTYULiAwMvHEGQFbSPTogDAYuFM6O7WsvRaY/PVttWAnsp+7vxyF7BbXdvH
ANFnqVUrz4WRRGIlBSrfkFzGmEmlD/7HeiAwuQlIizSYFxVf+n7644qPKgmb
NsNSiCUqQdTyghe7vo3O5+QM0CgYpblTUYBl/wGM8Zj19ZdvDmyrIZQXy5RW
HBhlwnHPULOwX7bwHPnRIlMqRjYmfnpJRJyVSkpnDOS6/EYqDpx13SFXNAh4
1uedDNcKmlYfmQZVtPHc1E1BlUzN21ckdQHu/b1MD1HSp5++yX/NT5steJ2i
gkScnI5N9Tc1+SukhgfRS7Gk0p48iIn9BnJfcVel64gHbhquFG4bWusAIHcq
uSBPvjCX7Qtq7xJM3dhE1g2UtpM4vAHV5F7MMhCCMz+HDuWW1eIsqcyZOZM4
aLtyixN2z+6xCMX2ia/hgor8lWfDIj0d9L+G9C7hbqvkpH+dMO+3PmUwrgVn
+uuLa17p/jv/wbJgggLu4k51T5Ahk8Y2/xixXaqcwi//YDFNpYxCw278aIi1
HEYY2OhQHQIeCxSUkv9pasv/sX7EMbpiBtIIbCrBKqVm6cuT3kYUOe9rCrqE
a+u3E1TdeP+seIjRQdcg2rvTEkWINB0CAIyVEjEIu2dSdti0t1MQ5Cima6FN
0hC+eUVVkutQe6lLusoSE3/y7ZqvqKKStTWDO0LddE6i13MvZOg5xrG0vcDQ
/WPK8mgJq2yboX7zkp6/N/Tcz1CH/Pj/CZxTojxhUlACzQgqkuVN2T4XN+pZ
Phfd78IEQLBBaUbRdr2yrZagolYsV/npZ7DNTJlt+p0V8vhTu1VXyUN0lSb1
yZwB6KpwYDJk4t8S7yXGk/pgANxOZcmuP4YBPcIAuePY7uUgEAW338fWhGpx
OqJELDgWrzy6S0JDg1k8f8G9AGrFMrvjE+Ygon5i9GRCjsoojwOa+QjBi4vK
FigcZKYnUSVVjOMyVaBikXjqjrT9g7onctkkCrh2Xdd7LCozvGh5cxYy5Q1d
UhDeO2X4PP/IVaFHy0j+J8RPvkGyQSjDd74d6Sf68CG1zBGZd006ZSFGVQkB
QmRGtYTs5u61yB9k9TmfYJmZyHqvrox+59W3d2IauMkNdyrgWnaM78bOfNp6
CJ0CdglUyVdj0gi/ZSd+WwDwLJcxPFyElTxB/NN0ScD5Tj1DEHhWWKeWKyQw
q4wJZoFS3HfrihtmEJYFu0b4BBBSIvRxYVisThhQuMIqrc2FwG/4hKWM2VzL
UWD7sbdvLu+8Ierv3RVGOHjHprZW+JHhh6papmXC4LS+SsKCh1+B70IrK8q0
3a3eO8xl5XVRxo48vfHqJQu7+XYsGAnZ7rD//nDzT6qITsBN1xXZxeBa4RmB
NDgBdoindmrLRNn7J44FMPcYX/MOPVZl0zzZKc9wYlRNqmFdARtfqRUqZj2g
CdvpXcGQGLVmfyMwlOlyjOq/UvL2j2e+JR5ApMXJwgx6AUaWdkPgGJ5tIAk6
R1fAzasBmT+oysqMPLJf4f2MWP1EtbiT29UU/YTLH53nk7aH8bhl3J/JEtOJ
mqXTpROMM73QFmEh9W72U8yhRuaxY9Vy7xKjK4SASOf/g4p60hbb/AcrRjNf
Yih6ISLYQZV+9P+InIOLXprgENVw9l/bAawIalYkin1RVQcG/Kd4F+NDGqyf
rnc0ilYHr8O4sNzgapTPyu4m2/NdVqk5bOfJWDcww6EjNI0w9yJzlovAfmVB
qafE1DBVEx2x3gNhWMqa9FPcduULhSiKQP4lNtsfd2PuU5u9wo0v1m6AfWeX
HBo+kz2s+EHuGC4NIAwDTimy+gZONY/6g/NHaZmFjT/j7gij+7KCnomd7RNF
mYGYSn8q2WbXW1VvMQDPmszIlrIB1sgNLi1GTVNN+N4c29YiwvtC235hNwdO
pSbu6iFi/HKHo1Q13HGtnauUAsuQaF7F2W6MYaJrfXZzy+rUotdQt5Zvy7qs
1RtyeXZG42Wd1VlI7s9kZuZ8+LyyTVysSc7lI5cKFWUevwLU0cZ7bUz7ae6M
B4tPLD4yK/w6T3KZNSy08X+4Lk6ntCPa73vs6poqJe9wPool1nH/JbMvn+bw
Ojx+S0aXK3LGbkruf9EnEa3C91mkRiC06cHsZ6+fdHCLenvZHmrQuGm+EBsb
OUwJjHBxLOAT1XNbvmhpc1JrcY8wJHKwmhXJsDtlperNb2C47e2XlMvCwB2E
jwmtjFnDdwVq0f+REKkeVBhRNXb86Th2y7TV81JpXPU55IAqBWikiU0XZ7A/
/RH1a7karscpKyxzjwMVsm0frWHJ38JGExoxh9RjuppMwtpj7b7HWx9b5uek
XcOSlq2E3vJgV9XQSEKbgUtOkefD+UgId0u+YWUoQG8KG3/X7e4/jfNmhJL5
duoO6JtSSQr4Cz4BZeE2viM+7IjfC0jvMvOIEAeiEdlqw+Jp2mQc2PjUI1P9
hmYwkhL5a3Qfxtbb7taWinPgnfhsVj99gAwH9BIRe4CabPnhYvTuncIF+Kzt
9HydB7I6JXU5BVOruXb3LZgEQphyAIA9NTn1OHrSQVFDloSCqRhieAi+vLhQ
zXh4e23MXIypO33N3oZP+YePxBWjnc79UGGs/tq3B9tu3nGCOVkxSsV+Lj4D
2JwrIY+5SX7pMaUQJIBWtyEBWrc++Cjo7Vg+g4xtAYj6g4nLYIGb3khzwlTr
Afihv2/3UEG7DVAVByGMaE/ImTSlBVJhY2wEFD4/z8ROVhcZdDHVOqmhb2SC
q8A/N7cEl3BB7StU6kAUW+m/TbtP+MBXIzVcf0wIGyBp/dAggmVCu+RF/GCv
Kmb2CKYKzh7OmyZoCrsAUvrusWkTKhkEWjqKT630m6qP/ThKjFnCL5mnRUn9
NZP73BDLdiZfC9+O8MItBrMbo1xezCtCCRFnOMza/BXhO1exxpY9iYKcUb88
NqxJ4i25+u/v5RTibdUBMLxxuWk++j3GvUWa9DY/P8VtkvpvtwkL3OKP3+sR
FiaiTFPHaZW6BHiAQdom3bCHpAL4N77ZIpiEeSC0dGil8LxCFGCwpy8jMjq9
Bhz3c3Vig8OTscQRw5t9kOpBSACOzZQKX0oGJ1dxSdKYXyeOcTij+G37yFqa
fJV+VDiMH1LGNDMmK4ShOJkSFWiM6M0ejLaITEM6jQAez0GKbE8q7ygMRANs
hRLZYefBda/lSYXJigPWzSQ/SBU6IhL+BQsOi3xofYW1KKE7Jk9UqWLVq3hx
cQ+dO2y6ijXpkY3cACcSUOU+dzbUPyUMPMLsk9YR0GGQNcjbLVcVa0MeosiP
oIQ+Tc4LkveVrPEGQTpSr5AVR3eDA0XJjsPcunC2Aqd7KVxzS4D25qVTPtgh
HXUJjcSnCoRK4aWRNQjEXiWNVZg3WUKwGyuY1pTIu4NpH6Yx2DXQ1qqW3pMI
DceFyYF7rfL2F/aIAiLdkbOa1JrZmgiV/swZqlB1JnXttGtOmShYJG0z/jvT
qyW8ZTpbEUjZooqaWTjRqTA33WP7ICb50JQqZCjoIk6oEG4evLyuxitpbe+x
a8+sYiB74hnwBgKffVMro9RT85XsU381KKr/Drj3PVwQMXyVqk8A1iinyvjg
5U3nOjPndFCu06sqiRpIwGYTVRq1wuqcSEeW24y4FVwGooe9fsrwCCU6rAMS
mxUL7TOlEY09fjYkXv8Hao/DqaAoaKyq9t6W2oAKTGRRKVRcIZDwudPGPIGk
T+M1FD2fr9luHRDkyA3mqyr6PjL3tFqCdHcrcd5t66N4WVrfN/ToohEH6Qc8
8uu2b/WR7ofwe5ytXvsCg11kIYDi+m3aQuKUSPVSUeiTS7jy2KyDavYgfqcF
HVNTcXR3z1vs7K0vaQfnA5QRLlvXWxAKpooppKgAmri0hFyX+2kQkRq0jV5X
ZOqLMC0A+LgWx9IZurr4hORHTUATk2qNtx33jkZcAcKN1RK6cId6m6JOr++1
Htm/h8ALvU0WJKhEB+nJrieIYiyUTUnPLlpc5xai32EzMdRgaPf592cIoNHP
me7SulkA7unQg4RVR9l6eaL7kLEZmYQa7u08YXZXIkZr77LdNDddCCLdo+0H
4iXNi4IBTb14x8qRbD9fyzoEPudvLYy/my74u+jtP/1vxBPeHF7kQ7xpzHHn
XGtZ4ZRL2EzkDWHpTav3R9rOS5LvCGezTBov7nYzq9P3yx4gd+4FhBtYccvT
pzCtKQrn2IJGjz5WNpAnQCuPpAzApPHQthGU9VeXLvyPLarTcEVNkIZYb/nb
bwOBg+RZzF952eYXl10UiZ9eXzMT0MSVpy6vnNgDV2wDLkdGT+A4oDnLDKWT
Wyk5Nr1RfHxcLCssO7lBdmcvAKM5VPc7sXidzh7oNdYZ7tCH/kcpQo9dH1xf
qmDhJt22b2VZ6eqQfT2ptwIONo5Jxz6rfaMY0acvu9YATjPnxF3upza8c/SO
JPunO0YxTuM1voCHtc+b+gW937BtI7Qpi6GGoD7H5hwkl6/ZpwnOckRzcAlM
B1Jv6hNPTj/tLpmYiiutpBUBhEKhp88RpMn8JFRFHqTz4eaIE9Z2vlPaiYp0
87vpTSvftpFMM3NhV6hrKSD/8+Z0d/T52D599pveLEBn6hextn5hrx5p52wT
+nHZi7nk+omM/diktuPc5M/ndUheiigvHma7QBlSCZ80Yv5K43yC/Ab8gxUi
00p+wNLjf+o+D6EGpL5oLXRX0v6TiixjltxZap1CwNNkY6HhEsvuMZG9sDST
Wnpl3wLSgs36DvfG0Fj0wNALHtzQq7c8BxjQU/bBCwXzh55WAOxldY5R6j27
BNcgVRJLmwXffAUfsOWQ+5B+gnAxf8iegk1RG+GOxSVYmpE7Gf8LO/+HeQzE
u849uaIJEyU8+FGRWUu4zZyEfIvNAcFj43vQNzmDvvzc1MnoZG0ikfvoIit3
AnJS0hAgBBHkxoPQgqjBBeYJzPDsbDuM/C1Oo0OnsLhPj70jVfIkP04MpGXz
G0+jJttiNJ+V6K+APWTTafETX/37MX9MEW+Ua2EXfSzBlwn/sKNcf4G5iw19
FzAzR30jNExD3cGnhtzk1YjjEd1gXDnOIofYNJP4jbEeA8Cc6Q33qDziEMd7
3YVVU0xEn75Q57qXM29sXII09lqq66cVQrLg24WbgoiVlmHzv4hBcRt2RfuU
it9o74xL6rgMnVueg+jXZv1WUFLQpbtFJ8PADt0r7ROizrmM5vhM7HfWFuuN
L45q3ZxUTh2QDLXLEsUzLkgNmqNyvoYWOtt9b9b04nn+uWOuKklRwXvLpGqJ
UQuxBnZ4po6/l4KZPfg80zP9jv1R4+JYpUb/L3DRiLzYOIjS7iF77PnrBmIi
CdKSBhJk5m2poXCqPkkYB4qvtbcLnpKWthTOVElFSSPm89eYN3dUr8mM4ncy
wrSJEY7/+ydCVfusPcsIEZF796BXKJdaYMnrHJRYwsY7XdK4gk1UO4D/5+L4
ySTsTNofnhPKxkldarwchFxTsNTxqdrKJSWMsW9vVzIDRkvLnq2WraeQnq+l
bUPA+Hz+saUCR2gslK7RTUODiDyjnIpcv9uZqC3rNmfxwCeiCzrBCpt1afbI
yLn+CVqZ1Gl5EWOPbxN/cddCtfLyWxot4RqJXKtaayx3at7dUUxV/zKvVf07
cvVCyk/ftnUhi7iEa0fMRDSS4G/wUc29CnyfBuwhE7IkGjmiaKUQ7Q57wPSV
EmWgRg+075B9XF70/BLv4HoY9tbgPer+/HQL+gbk7ZD/suO7du1qNqFV1kj+
uRiPBAfbZDD/Lq0daO/ars/7EReLBhGxI9IFKuk+Z9tiW8p8ZjjaZt807AtQ
RI9644qc7+Z5Qhk8z7LOrejyViXKbOd90/sXjApLulF18Lmh3X/tYjt5Oh40
4afnlvLJsw/c42upq6AngaCyq9yjXzVyy04v8vn3+tvqyS6xFJp3hPerIhU4
vosFNEOw0gMeBL+6/aAc9CL7V48NXNRY1ccTVwSAPnM+UG6bFt4zzIR3bYRz
aym59Ph/86h8yB9DtxORxTDXy46Hg9bTlCSG0CwfY4cKmMpKEg5L2Wbl9pmY
qv7nW8BiL45zinttmYabFncwcWAWJt1hbhCNvajE6MYSobpxeIZftfm+hqhA
msyAF2J2lIRU0vwy8PwsP+w+a+lt1oXMJHFcqS0DxsY9MJJHeXZfBxrfmfvs
QQTcVx3DDWeHRC7qWWo17Bwoqj6lZs6dcpbEnotLBD9rFB2Y3I2XFcppNzY3
sdUHjnJjg3xmEl+pnRdOts2OaXilxoi6iFp4VZT165baSuz5ZtE6mZjsNTNE
fVaqSFhHDtXVif7RQaLxB9Rr4a23ebXd5QvHocgl6r4rIEh2qDiEBXJ1zVPw
dUGMubRKGeI7Y8/X0uUrDZqPFaTQGHE4HYC2gzmWRYGnwgxxjpGxTPvDvk6P
2LY2z605kp4/kB7rZ5H75oD63dRBX75Myc3B5DptZpvxQ49g5Vrwwt663fGl
f8DDtGJVaoszCffGdBYuFCYNE3EYC/keNkIyh7+Fn1alNrjw0Hz8b5jxvZPn
iwHPPG73Lq8O6C4WFdF5TH1tOmoGNxDKWOufMLq6eCVgdIs5+X1AfB0TAUeE
bzA8uLD8mPtoXDUzhx3k2mc5UddZzXyrJvIJh/17Tf4vV/rfn6SYB7078ydO
1DOLpJhfK0MYYJWZvDqi7DnBRRUM8ZujOWNvcRVg/conyVRfVa9rq4fUw2Dm
TEYv0huzD8magNEShY0vHXEUNODAVtqlXuIITsD0UmTPHzsXkLZEppIi012c
75IGORsqc9oXE6QIYRqoFD8LBuRqrGVUgvDeEgJWvMRKCExHVPv48zjry4Qh
GPPUttop/QqSMnYd7Ki6qOKa6weZ+y2RahEHPxBgxTYTTFe1StzNAc2GZFpE
laVSSoyy9dAaUX8dTzWhzqCrQ2Eof0SWo0PS7Gs6+wbFsGDJXA/4D341KdkM
CZNgDf02rCiavgKcTVz9ZsOgIO7ISFjwMmV1iAtRcMK0dj3pdeRvgFHYGGX4
5lKeIpSbewC1kV9pTu5YuFhp4O/Ld7Y3++uBMlUyUHYhf0TXZCnlKWxZvEhM
l0ghRSN+94IX/fS1u839zzo0omgshRtF+z/AAtngCeXUf8SgUBjT/oB5chop
v+CiULxf0wlBklj2V7omkP+HiHzDH2lmWCYiGBMnbucZZH2i5/aD2S9M/5sQ
39PPj/OODud17/YgWcP3atnr/K89h3OlSQlhDNt8fY9G+WVNBZQ+wSizEzo2
VVso92ZyLKTH0ZoTBlkqZpq/kG8sclj+qPCHj8k/BMzDosp5CASOKbVNW0Sw
LIFXowcf1kfUXTX7K8cYWsi8s03t7lY0DTIS1bhFPptj+lSrzfv2h4COE5rJ
jd0zEumkMpeBSPxpCBleeE8MtsFEkVfxZO3OOCPoLhsLa0C9gjWeMCtM+sGl
UFQeAff1OjlrqLP8Ach3VOEWZ0NLaCawX/QjZjch+0qL3cNzv6RR//LPZcRD
+Awe3LdJ6K1HpFzCOWm5nETjq25yyipbpb99BtpOpGK/95Xg6MX92fgRRn3G
QSQl90BEobHPEFaNqYwxm8nZ2Wmdvs1ER3y84J4uREi9RAFkNPB/oakI/PEQ
BPMvucYLoGIamlE8udRF2mqihn8NnhJ1jqaaD+wuVwnH/ISEVZ9TPb7r9ci4
TonLtDGkZmHiZtluPKrpsuW5e1w8Q1tyAo9obfCFGBTYdAu0UrZ7W2Ci7FUk
9l82tV696kfGDOqfaBWFTXeowWyNzBU8Y3s5yIhoUNaYTc4beSdeNU7hf3B3
7jB3xhu3O7UIcVHipTpPpTGAWJTkpveHwK5le1aM1zWCoANqXW/LMwTBYLCO
T/FR37xsn9CcEdk/LxblM2veNjuqhv6lIQzWXEZy/ZVVZEdoB99e7zV3pCTs
p7VeojoXDuDOz5l0t+coUNVTrNdgL+IBT8QGAc/z7UQskO/1GWnDYNcLJeet
NgFq2e87CfLNguRBmHHxD2fwX6akBzOIoQaehtnH4laUFpMrd81ajGkmQN8m
EjTKbsCGMFK4CYUY924jxBA45rxXboO/4jVl+Kj9gzEc/3TqvMAiPLTuJ33D
DHSkJx4Z/CiNwPrmWMETR0LA1MYh+iPuv96YjQnCdwUHKv7xjC1IWMQe7h+7
wHzIUpHl7YbHaAr8rIP5XWxgA4bKhPbgtgOg45D3SfhczAnq7AUe/D0Utovk
XkfKFNSm0hBwW94RhVmwm6k9geag+qSBSvH5klZZAnfKghtn6fm2TVTNZ1b8
NgHBbSrPRfuLUrU48F0Z9u72EzJ/7fnnipRZatyMcLfD+UMM2Ew7VnCQyiJo
J8+5jNGkEtyzMnqdNu5MpXESfGc/DYMYCYJuvMlXbwCeW2Jwu0SnMzNpiv1c
mI4pAlvdZj2kEIyFmUnfWQaaEWEElmGWlgZ8yTM3oVeORfl0pOyPaK9nUwxt
dVeLx5Sq0kotsGwCW09U5jB7TwSw5g538o5aMCKFhF2pww2Qk0aQoa11EdOX
OYh32MFTTioGLJEVEk+zneSAqOC29bDf2PsUEj4mt4qyeyoyfP+UzCAF7XtF
TPlWgUy9bxCSQkrS0o84seglWILXXxY9K5WYI4uoEpEB4IqEDnkfpzdXdDKw
Yu9bhLXbL51uOaqkJ2DoDiqLGzHh/2hnaUhUpHS2vE1rlP00A+EKW5sNX8VD
TupysSAsEqV6C003KKB8gQwpah+lwutIVIz9LnHgb0cl1cSXyPPMqrtS4GzK
LgDSrUGDHz7EUCCyySpbivIgY704Orp8evGBeAOq3+Wd0UxKjF4b93Zraz5j
tIGvo32joYjQN4aaKHnaVJNJ/RjwssiY7FMDrYzlbbCcNc91EYAvd9zXb8lR
oBOwooa17eeQDNLnEhiHcRdbDxnRPD23x72107C2iKNhDyVSBWudL44Hgs4s
AGjq7L3v7KP9iXOOrlelyB+cyKF3ZTicvX7V27ueG2kiMLn/3blPStmhiaJt
C8NvH7Cbax1IM4ZPAebfx+WC/P0A64X70apiZRKYGbhCh5R3yPAD+XekL0eN
97DzIw8kso1fFLNugtfFX0PV+DIlz8FnPhkHoe7Lah0rIGi6usft5y58XpFs
Gfoz7ZdsIM8K4Br85H81U0Ugm5qtFDoU95b29v/ue80WgoCvWFy/Esynp3gd
MPGKmFtJbbZbLYkbjf3D9NNwZliE5Vk3fhRbNfJdHv0w1M/FM46iepi7izdy
OSDZBKxTbrKuIcyVCdfh3v3/cNhWJfC/fZ6MjzwIm73FHi4eVq/JQfKlRe+q
/PXVlXcHq3Zd4HxkSBEKvE+c7aq65tYBiu1J0xoIZ8I9tnkqWq9/njUbEUih
3ky+rvgXoNplrvgklNEtdlp5qUlsUHYadjLhEs8gL6xO5zG+B0dmTqyAJzG1
ZIOW0Fpu9eNYzwri+k1+Dnl3MepPEkD6SQdpgqkRR+b72Hj4XpqYXWqpYcvZ
RCtRehv7oSqCays1tnt5VBsO+m68Xed9o+75PCyVvlHe2vkZ1Z0Mvj7AqQTk
wwtGnFjpACHEgelVt1RZyzdjEAjdYnH1xmY4tH4CSQ1URkF01I40BeU8nWir
DFk0pAwrfoXlmSFXvk42o47ExwrBgj/dZDD379S2ulHzxrEJD4GKOKg5Rzt7
Vns2jsWH7dyakkOoOC2L4RJSOFnEcqtJobBJ0ZVSTC50++O867p/Yf/Sq7Rl
9jZvJJa0D3jFl80y5+lVccYvR3AYvsyoU9OwF1rcmaXKYMlZy8kM4CTV+vCZ
nYgVQLgydgQ5QgiUPDnRPBbNHswAI+zsJF23YAD6T9dfi2XwXVFMJy6fqp8K
BVj98pB8dQI2O1k4saN014Z/NNZRSWiH0NMEp74aOUgIi56Z7C1DppHub0Dj
n+cm28z+hIrXiG29Q0+P0TnjihLzPN5kuhYQmXcO5sVxtaMkjstmX46ggedN
X+onYNmo0rddw4QWXCfh4CMoqkrpymr36M7dzmYIulqgTeBVAqHPQWcImXjg
ZEjlj5Yy67ZBy+aoAI8kCc25/QSED3O3KxsTP/1UzcQdhg7W7v5v9XA02euI
xCsdeBr+bxmH8KX521Plsly1K7kKO+PdzKWX/mmvx6/27J+dCvQc6B4n4GhY
7HI5RyB6aXIp2cSeghZkdh6wKiCIS9I8/ujzwDKXjBUcxtXbK/yKbDSIyYXw
jFYrWOzWQhJUQTcbmKjGG5uVKL3ribc4NbA/jf5FYsgVm7yFyFCUmyzFCsZA
LWojMeFs39iz5ptc5/rXb2iLnVu4WlGlIMMd0g8975lAUvkmA2ZLqy2dUYKm
rqOJ9KYtpnvJ38DFBHZ2Ytz9lix9GlSKRmq/ACSO/JBwbinoeQbgsIZHVXHG
c7GkuJaxmlWacjpKg6l8+aViqDmFRmdYOEgWpx1R3y4+sgXd/Yzg1UlCyV2T
1Xh3pdK27gHt76Ink53aEYQs/JgDQS2qjIsTQj1X5IVhIPxqvCp7PPQJaBFx
1Fw7DlHQORYV4T/apOoQ12HPQAtm8vA3JTT7pnWosUfdbKUXVF58GXZAxuED
Cyzj01gmMph2KAT1ThfqC3y95Z2q1Qs3CMM9kHHu5ZbrRqKkXWuFBNNkOegC
Dhn9XEyLLmO1DxjFpkUX1mJe/GdnOvklFCPhzRXokri06RUlGtIFqSI+SLQs
+KNIg0+whcSkluYPcqAODD9T8MXgqzycyBxEJmp4CT38IP9+wOXZfBEQH/K7
r4Mug0Y1cZteD2CQWFPT09KEEFrrYBYfykeV5EgzsvP1KhCzjFP83K+Bk1/y
HXfj2IR16oipuA32xDBkF7lueuXCq2A4fk093NOYv4ML/qT85QqbuKI1A9+U
4ShMwYbgSZq0I5CMPRyY5rm7eLkBsGKkwLYDGex8S3KxYUFXtgdH6eN4V3cc
zscAi0NpEgcd94E+n8Y9BmPPNOwu7OoRKrwH2d/g3IZf05yqjiIfXTTRuqWk
PaIqtwz7WMXilrWWt1mM1oh8YD0mt0BH4zV5+ENYfEsFOnmYy3jW9htodNRQ
ORK1G7fKSUGG3AKx/C1Q7LcpQHYn3holcqpMg6h5QW7dv0v5Y9v0iEHlX67e
uBXH68rCZ9nV07vaDCWcQzjVGSXdCslrq4oLNlcs6NVtIMulU16Op2bjfumF
LcBHbL50TFcP4KXG9A8GCP5nwbawXgTjQPHtskFpyXV57lmJkzmIcy+ibLKv
GOzQymUdF60BGm8FAx1a+R7jsXKzTgI7DGXH6K/pRliEBzAtvHbO1uNgklCT
6GH9ybarT9pswXoHAGJIlI73iNYZjiQ8v3K9TjJ3VDRmLd8XwyO2GNwvOgDH
bVesnHoDzct5xc7G+n8f79Vkh6BCfCrT4uY9yhI8XwxvDRcRgvWwldYf4gnz
d9pWTvNfR6fXJPQS+A/Ca6VC13nzbDtehulVuA9RNhL/iJnR8EvlhbaTqyKk
Zt303yzeiQfvMu3jTn5TD0YnCLKEYREcHUSAQpWdIm7MMOM+Kr2TAT/7uPFN
5BeXgCG9PAvwWs+gZ4WHy74PFznkSTB+T5Jc7v5+bq+fOXGZ68Q7T4N3RQD4
oBg3exSq3oxXKjBcRyudK1KgWIFtu/vJ91AN3vXEvMsoRV2fvZL7Vq0jSsOx
k7z6HF3l7kfpmtBFwmO/weWMHqrYOdQhUHHrynq0iyph6nsOrLn4EXw6Zt2X
mMiIoc9IHe6sAspJtmJkiHbUKLdbo/WI3yh41yMXeJhu+YO+S/N+VVCVezym
PBxvN2unPoxhI6ZEYZCqsCr2hDI6/Ngf13b87UOfF4mUHiZ613/H5jM0zywJ
A6AXRq9TV0EIGbQqFrdoMwjLKC8Sf8Rahq4emhSrcgupsD3nFTbg/twiTSbw
EP/73/R7x3Ot7lgrkNVh5FBNDEvV8Msgxa/xND6L77TKSqY0UAcuhbIXmBLR
UHoz69IAlmuzYEFvlyzJPxbOkaB1PCQUnUbJrc/L5QSgMzjOiXHXppSEMTVE
oSxB5rVqPrDUB09vtY51ubXMG3gHf0mX9x2dbPzWbZwzqxZqXTQGqgteR88H
RUDSEquyti+U03ilsPKnPa4hE2owN2WuUvWrZaOaTvy4yrKwgBjaEF2pSKJG
wW7y4fIPn8HYUMGFcv7bFzVoRT0lylyh/HSm1CQ7oOpMGux3sD2lEsJCf9ru
eVNxOuXOrlKF7p6GrOR8IbD7Bq0TwHIWdQ+v5L+WSZ83b2Vr/k3kjs7HmM16
jiDFIoOdTvXH3jXuHS61KfZp14rRdMTBLF0IBq/0IsFHUf0dj/KQXxnSoYPu
YFf+eX5zvO+s9eiK7YChvSpXBrupTjgLXcHb8mmokcokqiLRllTwee/i5dhZ
VQ3yfXBiauwbgWN/RxIwZjl2ksXpWgFTvhtOvjYsZ3isq9yIh3E5ZHEFJGeI
heDhUTptscPTQpKpezvJJ6VND+7WtJOrwDsUNc4xSzavEdH09F5YIm8dsKpm
ij/ENZfnBOEqUyG2gI0Zj8y59+Y7uLFiBBCz+xMB5PM3B6agGWBfczArg2I4
vQX6aUZHte0hwL2htepH58XFGIWd/jLz3kzRKsfuREIO21b+UyFFaZ6olSyD
8QBiBtbnGTqWxD7U4rTV17FFAZ+hDTt7DP3Lqr1CYVo05V3jicZMWWCbU3G/
y8+XpqBta0ihqbw9bfRrP/eXMmVw8SUuQJfDsKR2D5Eri8M1rhELL+v92IX+
xaNAZIpwV7PexfJ+UL+HAS8SEJ2vttpOMLTDKSkiQM4W/hvFEEpsra1kVKQU
Ack2S81uqyHYjoUJtjMtfu907eCPNk9qtO7VPgGMvfOp2WT8yIyFySDFKMAd
c8sLW4oOtwgePc1uPn/47tWnEKYrsVqPHeAw8568z8oFBMWHgy7IPd0uPBy8
8+kQUCbUVr0EEFtb74Nml5zwHQaYmPa2NyLc10zPYnQzpnkaQU2WyHki5B8W
0267O/a702MOcJS9LwvTzpRQZ4qNXLGnlSzziLmBKsAOsnoxJAqV6lorSyGk
CdZsy77g8wPnG6klP0SeTsnxS4HqWU75lcX84R3Yc6RO4ohOqH7io0SaP/bk
nksReUjBEEiScwePnGNgwsONqnilePTXqopAIUpaYolvome434QuHvs0BRad
lQTiadn36eOJY7G7fiGZPDJWabtGnspvJM+HEvCklo3ZyALL/KpNmOnTy94a
SXn2+64xbEyb3SGgI/3QXpYhxy8/sZw0qsZdrIEmkUou07as5/Zg6vrwXFs8
lciVL30jJTYer4QqQKRQsoh7beVfYhtrulIEds8v1eM8lwcHx5vhxAbMtPt5
D7CmE+ZVAiJoStaoho1E/FTNR7ajINwUZ4yz0eZTS2ycVTvpuVmB7sQ+hIzC
eLHi4BbWYFewnxBuFrrE3UegGf53LpGsBMHsS9jMeb21nWLMOebzb64A3RPw
BZY6eX+wbSPwYyQ+ZoSBIRDKt6MHse7C1PYdfRq57Mvfpi4rIUzu9xN2RgAB
Tx4zcJXUhtCBlspQOAq09r6WAYVK5ffkqTBNLXFGjEQWS9j9lLyKGpRIuql8
Yrm2criIg+Oa2TxWh9990WAwb8LVD6wbBvCm9FtXQ9DqGQVoVmZdN9/NBewQ
QhlclQJuFRvil++0zpU9NsUp0AEb4DMhRUsnQSrteUVo99XnO8PFsBLSk4mQ
ZFSsQypnS5lnKOKFIQNanX9XtPRhPWFSJXdpHOviYOeIq1csmytQEtpqmr+a
V8y41epMOiGzLRyLcLH2d7jJKnmUMQl4KX4OPmWo+f3sCSGeSrLmhuxh4/6D
8AnBlrPYw9UDl5lKtom8L8gSskH6YvAWaWtwk0JFgbhnHNM2LhTpr5MygbB9
F4mViU3eRzKaP6E9Ak9SYKBqQtxhLvppK9CyPg5E2f+6XNO4hhXTulIUKh5Q
+ZPHERefYesUdZoOry9r54xUgrZ12SRdk7Kb5I/djjHJz3A5MsKy/p7qdt7y
05XquwkEFo7DIP1us5fsbbTrb6RmjtnMh3J3SWS0ILsfShvL/HFeef1CsD9D
C9ee5lR8Tf5EQy7M1LPj2jUM+wawMjGVtsuYqiC7aIHvLtjRYwxTtpJL8d0W
fMz+Bhfk821IjmCwIkRhVYuBG4wvAzl0RZLEa5ZVTI9jaCZOeN9IiL3JC6Ji
+5GnjoiN00cMnLsSs5FwpfMSHk/3CN+qKQ0j/2UmboznuPHqjqg+IQ62pMhR
YfM8nGxI4O2kSwJjhcYbTrstL4u0QsbV1uJ3I+E7cfV58IlEFiX2wJ7gLvA4
aRL7dO9z1y0U4xiv43nuYg0JtvGD1RO+dmOwfgJM7DQoJiEhjKoEoMee629t
BWzNpVxPHH0Tp5iyJNXgQRwF7qJDD6FUV/HvYuRL/c8iga81tgmgilnLae7H
lLrsPzm4pntmWFZ8T2fD1XOT3G588zlKVfbtHc8VEkMJ+QdEY6IeRmz1z7LI
zfCfTO/hKliujwOcWg7HCsHOQqinw8Q2IYRnGNKOxMkoF/WmnNLzVn+xBXQk
ykN7UKdX36Fn01HH7jwvgdsN1AYmQzTo4NDg3XmE5LtSZ7LFYNRhToWbnKvg
+mbJsPARjpKK0Z5CeXLvUdZbGsmH3CEM30MVDjEWWEhsLJ6Dp7vm5ptw6qUF
1itENW5QIqDwgKRWjo6GrM6z8jbM9+HZrJ+YqyeuQSwWdjIHpCs/Nn3HE6em
XJOCg4bBCdGHIm5QW4cOg8RvqbSrtGyxnrQeI3gwIonY2fjz0DnfU8PS+oBi
8o6DKgA8FhDSN/PnEHJV0NF61crzGM1bY3X9WQcbXn3XmKaZE6wELgg0RBUf
hTN7iiHKmisl+pSXy6TK+TC6uJBsZwPdHOTKzphpPX1qCKa/6A3BGaB5UGjS
rgK2BIHaEdQCqP+yiYpw63osMhF2Osn+0t6CK+RMhChIIJGapAZafZe2BugS
JSMBpFpp2kGxs0xOcgn4K6LiL+4Ol+Gpm4GEBrNZ0R27In8bb6bHnUPPUEGE
0qLkWP1fZgJdYwazYd0KM1b9aQXzaBd+PD8PfBbdiSsR1AyJgGRbPw9u9Qop
Xc/RQfnMU7FqXUeG2MjNF1AQ0UBIHisG+fOWzfpep07B5JPkNkY3nojEKKdL
RZHO48yvDLOu41QiWbWz8k+uEmZEcz818Od75uu+hhTLEc0ss80WXOn7Bv/M
1hM4+ooKfGOg/yN1G714jXnJvyog0/7DnoYz/sHvOukVKrxchaQTz1vkFuj5
cClHs+YZEeHXtJdI0t01CzXBIwEwQYZ7OEYuCA4W2OpLWVO2MOMgLKEUvPTu
7SCuUh1L4ekL7MpJTE11AeBRc+d37O2lxeJvHYktMoqMFFzDVpzGn5bF5GaZ
0JknNwJHV/tMf6BbA3XVPrJDoX2G7UEpkABfkV3lKDMQYLnZp/s/FS7T5IY7
loOZtyc2ZgFESxATWudzoaISakoCWfyedsMBmgqmpvcpKxFMjLOz5Z/nR922
ONYmoUTJp0C/oesJbr7B6ZxYMwpz9sqo3Md7FmpLsj3SQ9pXmnU0VZwfuEW8
3MxnQglygqtsPBbKtVUZRK15zaAeFEFf9wSpePPAU69rRvq1d9TTdiEtVF23
ehKzh5WSLuWTgf3KviMC4KQulYHAhmJrF9p7CuojvBDfu7KyiXXHrXSASsI2
wYnt34OKmM3o5+LkuSrThQT+ozPf46PB8P0thEnpWRvuyezbb4E6fREvvRqs
DJ5mUHKdwWBcMpnuwKOe/l2ROf13UWdD17+6CvMzbp0bMj6DDal3/fOXEoc0
iSNBpt4gUQ2mFy4mfUgLUP36a+Nh8Y/Ec3ELP0yxlN2k089T6XhfLhPt+thj
jz0GJgcvSpDaXiyIvHPORs+1krVgmuJq7mvk9sv9ROkLwrii4gOldX3uj/aw
ZkF9iF2LyftTcOBr6g9KQfgvR7hhJg7Qk0LJW+nlx/c6rOatOZfmxQKcimFG
p3UIVRo79HxNvyOMXGox1f9JjWjxp9BeuHkiehH7mU4wZQeOTC3kbjOWxDZE
7TUzdEykz14QSLb01r0J5dnQudytepMA7eSxSncO5cOnd0kXAbJwSZgp8AmK
EvR2gqeUaxXQR5D9396mOXEjVB0Jo6yhJQcYjMyZ3HBfolRUymz1j078Ro29
sGSzsH9ydV6eULPkKfOfMGA+b6wQ229CMnz5FPwf6+vZYDc48pMJURdFwaAV
oI/uX08PtuFtztSMOy3Ua/XVFWzqMwiAMd5iiqMg69brd4Qj2uSzjZIMpQQp
VBufpxqTgcsy5DRyraCU7ljf2grDuc5X1H8zGHrsdR1947Ht81wJ2ebD6jQQ
WsDN/v6xf/FQsMc80eTePDRu9IJ9uvUGnkBklvIHhm53ZxMSVApdrpS3LKzX
vKPi+fe/a1wBqN8zDvEyoRjdBDx3GF3sFV4cG8os3YmM25dsdI5U/pWh9sm2
cc3RKew9q4ozJiqpjUdfN+3gTrKnCQy4R5xtyjXxWcKC/XHGNa1VLWNdPkFo
spq5EpnUSWkaieiAA5eOLAhxxQecK1yBgXHj54her9sDHmG9uwiU1xfIbpEd
hw1SNjT38OOXcOeZV3IsYozj3l2oug9dq+FKT5t3BoZyTAjf10yTDHxeIAOU
GtJ2JgRMA1ZLN3Z2fk5a29n9GCFun6PPOyuQUjPI6c0qCeds9pZ113VZMLN9
IyJ5rOY4dq1Qxdptbhqr+TTXRwSSZEPEmQ9FFtK4dZArrOMVxUuE1Ubz1GLR
rYMKNl7x5xiBAsAvS0849fMkWQCLEyM82WRuKPia6rUeawB5yqfIn3PehcTi
9VWjX8zSyjNQFq6xx7vae8d6A1+b23dzTPKa/QIbVzWzuhrDsPmHdIcu/j/H
QVWZ1CLcyaOamV7WEGQC2+s7XxcYn/xQrhLAUjaDeGWOkFWrOhqFTatJ20LG
thjGIAQLnnqZESvHFxNOuWVT7pRQDy21MnKv0DyNfJkgQMO+NzmH6infYLqi
rAXrYW2tKcHe0+J+sUf82DtcSlLHDJQlSqQeVJYkC8JsYmrpLi+L6rnrgF7b
kyfLWhgXe9dqISIKHDP3XS03Hq6Pg8PdFh6HUeaRWzbnRNp4SaokhcOoM9Jt
yk7HbK/mo6JtzLSKK2vbpaTWpiVy7J6nah7HhsrB6JANp8Fg4Edyi9Fce6cz
DEiKDvXGtBhXdlmnZ87raTer5S20CZbpRPQIX3ra8iCTBWT4bf3sg5LlS9N2
UGCS/9fhLdD5R0hw0OtjTzwQtgo7VEtBaGKpxr3QTTc1j3X80zpCPcC+0ytN
lTIyhLVjkhpj5PFBN+090L6Arsp3jOs7jKWcs/1gs2B0sUOqrcHOblPUYKmY
JqTlZX0wITvg6UHtItrGMFd7sV+hFlMzbE8i0FHZOFk5Xw9KirV4Fbu2gJk1
ISHa+m6WAhPTq56yTXONMvdsHThzTqR0tpUVu2XnISMJZ3eVkkeIZmGelSuk
opjhOX0o69fm73sgN63NQgIPJZ5Fq8SfNJFEdrCNtpfwR8zGDwacSgSnAEg3
5yc7T/s44Mk2++FgSoaLrFf12KEwOROTDvf8Q9QFPJ4oeZvFK+Y+efoRR/gw
yaFLkLfnYKJG3+LiYLmMJSGevwotgpug7WVSnLyFwi47P4mUmVKAoS7R9uiD
wIMLQw+Xofc3XrWjXjMiOKNXy6gU+uNS02JJNKtFHnOPzDuI+j5/OiMg2xAi
fEPNchCOJ70wZ9WQb5J/0vZhi/g2yNnt9ujXspH1O6Z7QUmzthLBC4CJkq0Y
fi1NrcUX3SsByWRUmL55I0hOG6PF9NMKPB8axFWKrKbW0DXeWyH2EwhSyb5j
N22uahsL20pfMK5Hhv4Kkpw/cnf+4y3ePVB40Dj+CTIkLH5nrLuMHcQIhU5A
kQyogEG+ctvp9wWY4grBEe0WslFsp9Xgtt1qQyINF5VNDsCF1ivMeobu63bN
iOdfJdzq1gCVpd7klkpwqzZoMd2k9tyyzYQh19VaZEVXrMDZFsuVopIrAsqe
dwAE33X27LnmYVNm2t1mSG9Lchs+UEm/EDGX/+4xS7oBF/MwPHPttaMVCmaj
eSZixzx3Gu3xoP1vgJPaWxvYi0X1c91eLC0JxZqTWAD5YzaLZYqMyTI/X2eI
i96JfLWf8bYnb0iH8jjrm/D4degsIYeO1MfXZXODNAGRx1GPvCfugNJCgUB5
hlc0wQliDyKsmGFpQn9aeEWowoTsn03aXqatB146cWk9QLi3tYkTtW8Atpj7
j9xLR+K2MbVHfr+6ahYGEN+QtyzyoniFUGr6G8sAEevsSVcvsUXWHx7RefLo
Nr/2fXH//9TSpGbKoaGjBNyqA/qY0IdvVf2AfHvYdTjx0KRB5L7SX09ApT0N
FjRurKh0cUPV5Bc/9pSa27w/EDU77BWZiV4N3SHlq+GtcxIUbbkZHFlKmeQw
H308S7irAbFa33BTnm6JjAlDLFodUCtGFnP4hWRGo4ugFs6q7/kEMQVDJre4
WBaem9hhorfr+ljEHlk+K3dnTX7ctEMIgCl+RIrxMyowPjkJbbVGybxf1nj0
OFfn5FC7RpoteE8ZD5W55Lscw+KbWnqSs6BA1HgRGVi4PP//yn4X3tq/MjwA
UT0fMJZCgvO0yUZrXzCZ12Bm09g5qnZwXeDJOqrRne953zLwQtnIT0k6Bf2q
hpyj3bZRUUA/ay8MncPkQ9aoqsUr63rS123qSvbvWkyXCKi+KN70FiOhtv6W
sFengEOs1a9EbqWcprpn04CTIpwq+4F3XsnFOQj/TeAICBpfkivz1r5tKb3C
Fv1GgnC8rKAfFFzTIY/BJG6o/Q5nRDcqcj77z8O1q84PuN7sls5Q7ToDRlPe
wGQiLcJ+Ij8K8z2eEsOJNaiIaVMZey5t/6dC9CyeglyL44b6ZLEUKR6hG6Np
fQbLpLiFtdRkoh1H1QxcJ1IKbHgPGbC3pkgWTl+4rJoPjqS2Eu+2RQ0g/KS6
rkdbK8CeXl0XGzQvzlZEG+PDtX31v1L50kbEHH4qMwyQwTd+7Wd13ecEeigz
QPET3PiQC4dkCNelGD29vH3IBRZxcdvNOcybaiMXUkr6+MSwd+k50ZhONUkp
/8sCHwfEZlXp2WtiglAge09dLs+sFaTmFyD0/aqV7mETD93BHHurrZSjaW7/
coQOFnwB9NFSdZN9lGVtjqEJhqix+NExQjgoJ2tkg78T4eDtFTS+cFpPRvtn
1V6LKaWCjyLbxpovHTikIhKiJtKDJkNiYGTuCeKwRkbFQJ5/0DqOx76g+xdn
tciI59yge04W+iKhWSqzIEUeyJgQ9+WccRoovMJUO/IzROiW4ShfXoxNmOYK
r3EfhbbJqmiviHgV0y/jAbBclyO1et/FMFJaKQyDCJNik3aay0XFqLpR+IgW
KRkWxM4pXpLqn1ZEQ5gtwfrcpWWQ69mGiACzzxPISpYFUnThJruKov/AUAwg
yGVS1bu8AZ15GWN1Gk65xomeFqjWsr12YJHYI3gwxVUgAp+oGiFzIkBZ4pnt
mhexfCMMQrKo3kc8D0RFm/4Zc4SL+XSF9pOmdGefPTnpOYsa3PkVKTnFbnLd
qUNj0poUAe7NqO/D4dtEhrNVSe7OScoxwyDUU08dbs8+ycbYp8kH2E8ZGp8+
Qs84Kkib9S8SkAaSEs0u7vcmuvrDHbSJyfm6Akifm6258tx1vlA4Kp/BqNk0
gpJIrUvdB2eztB7SeXW4kiPf5sNxVSEcrs0oOSaPGfGaLib/iXf1QcnRMs69
eE05uz2CnrucNfN/uqwxhUDw0DOG+yY1K5//Z69W/947sZYE01d9wjr4ae8p
aY61EV5ZLwRwRKRT4RW0L6/9VQ6Zavh9NXrmcsZXGIEpG/ast1MMVocZYK7T
lcnuMurdA9rDPS+ieZ1buFkfh3DrzR3YQNtLjrxOOtprrTozTtqEc3c9cmEN
OVeBx6XX5YJw/a/unDRloLC2zRdBsAN3j2GEvy+YLxN4ONM6pAk/RPkRc9tN
mIZYryL+2xRecgxwbaeKdyPDS+5/9a9EObzGOhXuoo70mTTg11e/r+S6TkCR
3DER36K3S5pLDxdVSnAcoOAp/IPqpsK5RslAyBDohvLfvI+/oySgjrp6Z7HE
bbVhNHauaMXWmrdeXWUS8TvTlMVdFixOuoE6GNeYOtV8yImKv5q+jgzO+EAH
ywaS3h2Shkrf/YVz4Nwxt8OxvnJgdzo+LKX6mMXh31rY4lPHnQpaKNSWr992
YYk4Mz2YGXecwN33pSFWEMrPs55kJUdj4aNtIxyRf5gZRKurnA+AQkspgoj4
2J25AncwIf9oT6Ehizcbmzk2wwk25ewiNpPcNM+c7q9DPCh3fqehCxh2pVtr
rY+ZykXHerjDV9FjJCN5ajywk2qQEzwwWd4XbFKSm7KW0d5wFcQNkTVOwZgD
9xmXyrL5PCvNUQH+xAOMwt+f9pjUSo0YPLztIc7BF+QZbMledhyXbz/Buttv
ohisyJ/7TRplOHQbQC/cc9dbfU2EyB+0QZ6jsYcsGO2gaEM/UwYObVRVQTqV
0ejuS0TKxuAgiMDai6yNrR/F/WDsBsUFgE/XmWMv1nLLioK5Tg1EcD31JjQf
58+ROLcpDBaInWp/aftXa3AaW7obDXd5ftywXM0aQA1Yr9eg5KNrSaoHCkE6
wZV87M9Tm/MvqZNFohNXOXmD/wdgzT/srT33tmEgov5giVmB7A5hEWc1OIxW
0HyyZC7Xbta2mkGUHYHlQXbcbTK0AYG6gyRguc6LVtqVmm+LO+UgZpgv6OSJ
+x+FmD3++zprmxC2KbrdHp1IMx942nR087T2m2XUtNxHJJ76dukZTGKzF1Mi
zn1H0vylqih3CHQsIQ96U2QpNbqUegXgywFZeJ4IvWnWJoVQXY5En40DGLD2
QXi4rimPuaZSQIyeWMyJ4BYpDmhF/ToOLXAdd6vrtOI8MVrtuXgITX3GiYVr
69MZD3duVHTdOZp8xYhKtBDWyFxzsgdL/72c2JbCuDhwEbhgU7ouTngkqZXc
/Uqli9Juzvfu9tAm+uWiw5upeLPTbRjFotmlDWkuRcym3BuUtRBgtQ2qSoIK
Xvbx/QhaXIIsIddLyu6264sAMOg8r4GEUeLFTOV+/EtXRgpknMPWA35ELHlC
wTRp8HZBjnWvAm5xKSV1kZ6pud5StT0XExxAXKHXT/54JNICVw3qyEc/mcH1
wu45pkdBGufui5UdOUKrXCMZG8160xA7I76YSwPdPe98OhOwi2OzJqkekhIO
EkQe7JKO8u45Nlii2qV0rkt4lRKcmb3kPVNSUEbckFyQbmPgtPabCAPleUH2
nC6UHWSVr4OK4j7Haew/j+U94Jf0zodgc0EH2HUXoYHiXWLyRY984F5WJmE1
aH/rxC+YvAG5I+riLatBfyd4KHFp9iRPAr1UOfLVqg0tjW8cib6+ufiPrfsn
TY2ux9zNKI96oDjSsuPZYbRBrpimHE1Yz/PrSAee9h/B9KnWCHUgi/4b3/+C
s8ZpV2ohN2d61sDVyCfbHsL+I/HAvW2dTj2W9Ctvm9zC2jN1Vg6XlWF3aVHN
5B4nasztA0ByDVh9ChFan+GE43ZzAu+4z6FzH2zkN81toM7Ok45exKackyH4
bVdus5yOtkhdl+67Xc+9gnrYzm9/SITDLWtjASAYLiRr1B7k3+K2zZzAvVPr
Uq273YfGzILkMgfkVs5PHbcF4ImzAPssk9Zrcauxergv0190l/hPSxe7ahYn
0b9SzbZ/VjbhtLfru4Ks3wcGjkgkGarVJvebqRj6l/FMOFl1BzhaXIUVVnwW
fjHzEV4Mp+iKVwxCtLoNbT6Qgszm44i+6A4y/31K6DQ6zgkoATNw3G2ntlpc
06KJGPYHQaBbosbrRR6U4TDLVpC9ce00Gj689E1GW/M2E+1DbZnjqBn/WB9l
bQNg0vDYrfl+qxXgDL0SNfCeKosxP+xKB+ekZPP/V/49HQ01y5MVCOyCTd0F
gxIxDOkkOv+Mj0N9yTb312I05V/ARzD10jBMwkv4Zi6v6rI8NEGkEYfroVfe
CTOVxfq5zJ8jHbaaz5FwVRDir65sHRDUtT+2QxwwziSdUeN5FMlt/AOhTR9j
HBiNnpvlSMegoaSMYQ9gqbSIUKBYxrACMXQ6iTyQUGgHZWQ5ppQMmfSLC+6u
UfNG4BD9XgbL1dDup4OTUYlEwdsWbdo3WFGhD887Rs17MX0fLN/raLxbZdTb
VwkJDg07wecLumvNphjYKPS2bmHhGbtMkeVxK2VUDDg/gbcz7vE5A0i1Zquc
WpOBKI7I+nqWcGAsrKlmXHGkHEpqVNg1bQKZEZIkRFy9kqNZ08VKIayupRys
JCa5RYEUpyCF6//x6jISja4gbihsRvNsRSyzOrrQ0fCISsfyZPO9Z2B4yj/i
0HTZqKRJRKFLIXYKGUk5U3YhW1ouccBGU6loauKON0CPQy3RMi/k7G2C1NxF
/iXkmTZeLehVtkFrbUOyRugoeA1Jvkfi3Ko9pUZKnE6pWflv4WQ7RI7CTKrw
zrMzO32W3NZtetw8LhfTDBRCyjvxYqEO22Tx1jFtYr1QbksA6t2UlHgoWOoF
PQTqfYmm2WVpLQ7/pl0SenQ8zLeSUFMMOIHNpiyEAQow4mVB+DjhXJpgyHRR
4qGZ4imicrQlP70BqLnXPjH1/9/LdnY2C696eDnmP+L3boIp0SgUMBbvH/yC
ZOLnnkSei05iecA1Uc5gqFOIuvkATVukRjQVd4//Zlkys9I1jiRM7AzeyrMK
ZHkbJzDjMmdbX+2Spv1niF7Bz8LOjqk0VkeOrlDQEUY6TSYzViQoZHhNYAfw
Rpxtail0UzIir4afQv+9D0d61KT9Q1I99XuFle4ooakLYxT/5iMnm4F2qYvq
Vf7ANcfoEbF46hAsrhJvKnnQb2SQcGLf2Gz9E/CxeYLVa4ZzzvxiI6HYFkbp
DU+EVknWBxx3lr5CkBexq20f6iJHlGzYaImERouT3BdZfyLHPidokXIIf8HW
ydZewF8bOKdZ9LpyO0aQyAAwIrACDtrLJ878qH6aSqMfsVtmF0nQG4RfSOwy
R0G+6retIY7MBeMXK2Da167d7I77V6efsgSpDbZsp2MdCF5YYP6Qq6riO50A
OuNPZVHRR89V7guPmCSLBqJLR9fQj07pFOFBbovAe5UV15xi0jZbaBogQ/jM
oWfT448soD8GUJlWx0lLX1EruSQ2f9desLNyUJA0u2W5xoHzwuPFL0oZUOPr
P7kRqtkNT/BHAbb5inCJnaRGimVZR3Yxg4hjo8FQz8czpL9NTxWu6j1w7gDq
aHbA8fZ3qLy3Cwbkwgz77EA8KwBGLeSxkIyArZ5uZdEs9Jk6VY1AbYO+8Qf6
Rr18TPqrgrkxf9VssU+Wg6HIgUi7hToIJU1Y+uqt3ti70Jg8Hv69ooief5W+
ne+6sobDDauYdtCYEZjNW/9DRsJ2j/KxwQzdczB3I1h3EhnFdYJ+FzKO8tig
jugNrT+km4478AnCcsr5mE74LA2nYtn+pM3V+SepeRYXNBvKk5OMGct/kAJr
ed8o5hjWn4xTjOBecRQVsA9YdowH1m4WKxe3v7cEikWKr22F9ye/Uvb0L0bT
60J/B465s2rIBQcbA3QLsoVVw8UWy7zv0OAv8FlzxR4NpusfvZ7CiWSQ/U5a
r1zFc5XNHuCobU3FClthsMP90HHDPHFv81hyYuMecP2w2/TxVY9WPmCd+fDu
69QWe9pD1VRIA7iR1KDrYXAf5cQNVW3LQ0k55Tw+04kOtgPrhPL1BcazyuN0
dcoPjQq6696Orb6k+EPa64cYbNwH7BXttobvfITPMk9OF/hX7bQ//oKJ8kdQ
aEHGSP50fXSWVnF0YqpWHgdtwdXQ7rEMataHz2v76KLqe0Gi8JXYqQU4+7Vt
9Uei2Y0GtKMyRh/SUk6/rU9L3UPczC4+V8j1QYJ7k7akjT9dNS4bjzcAvouo
B+gl511wVdgHpchxDxbSMpAVDad56TzXklRdhg1P1Eoy7YJo4HmFd1X12eNj
Y9Vc9MgSORichtJH4x7WMuDqhHSCYM7mxVNPwV2Lfc4enTVnlJyvB7I4zgTW
9W/BSJxvVAFHDJJj4CPq/K+6/HQOYe9fG1BcUiTYPECjWk+Iyl8XwjtBoaY0
x+pR9JMMhA3h0oZ+tcV4OhwGoLoYKfR9o3x8QmdRvCSQHAPzlmslnoL7rDEF
bRJcXfEbuNKCtaedOCDhP9jdntPZNRrASzKHNbTJ1XJIvTrbp563gvspJIaT
qY89m2W8wgvNxx+Vi2IvoHIa+DTV4ZwcsKThMNcusSBWXsuR0yivMNYR56q2
jl9HKJTu3vc06gVGQPKv/09E4YI25jB6FkZSIcvGkS/egCffyEh6uibPMk0k
L9m6bADkHO92XHL9MxxTwlsBm35b+YR9ssaTKHvdy/dVRNa7TNLxVZSznoOk
3cLFmSzH68XqlGgWxTZheIuxPwNrmvgxaiKH5OpomfRVkB0ANbOukY7V76Mw
AbIYt0Z/bgqHq628xUMt4hpyvc8c7CoaeX8Ij5FFB8gHUz6XEUw10o83wLAL
IQ0RXAra+sDhajiDhaZrjw0krIUwzxMHCORMU/e9gexwK2MAiDsg7LCiOdOJ
DvAftMNd5JWMxHnAfuscYQs5rrRpdnHRmpPJvnxnMUIQgu+/mExodXtUf/kk
Y+tCPbp5/q0UzphjbkR3xcUUus0KDkPiy00B81/eJ/V+W83QeXgD7/Uy/LVW
/iSIck1oP9qN3YtOuGBqEoIeI+SICFbQ0UK7zTx5zykGYxMrFywoTSbxpj4d
hRQdOuoPb6t5HgkLrh63/cw4zHbrtKaCq8u6ogY1m5LsHg3nbY6RB2dCII3t
CnzFwXKcmdh6jbwzaKwFx++lzYNKvGubG9TbLRSMUwxrX29WnnMj8gtYj3Mg
2jF7Ijqn0T8IsAC2OqSh3YSHErLAygyVx0KGRRl8v/WzK0tp/oJOvRg3kmNz
2hMwKS7fkdjfINDiI9FbpUj7qmczNWzqbk10qmhd+P0OcAmdze/7lLTWe1DP
Mc3GSB2TlNMihT5y0OAqLpu+t2PYCZawVAQF4rpfD0tpNw9XUa3So7fHWiUT
w8ycRAaXwvaxe5TQUV7fX/MK5jrniKLTUxfIn6dHmy9iRl01z3aDqgimXgKp
LBiPYA6xyBIrFNJEgsGHoo+ezJUzQ/RbyTCgtz9Of551GBHCWF+KJRco/bzr
JRbw4tVtTYpHSIVIbVAtxL7XWyVI15tthWZeBRv6h5U0k6oI71mbYMDutviF
36u1orqYigLi+VaTYWRMfLz2RnQFW69kGm8NYIzbSWlOwH2Jh3zZvhid/xFj
MRHBwsCHSm4ZWL8ZaDD1dv/4xeQkHGbG4QP8a2X0d6kD5ts3gvZvVJ80yBdU
JZUdeoA+fdz+AiopEitY7TJLkEoWRgqH65tf2gIHT7AIpftbGT5fiza2V7Ns
0604Nm4FATyj+zj/kXzD/pNVgU16eP8KQ4CoTaxPWwuEe113EBS/C31vV4z/
KzWd6iI7kywTlM9xZgc8qGvq2OLYj+3Gxv7dHCPP0f2yjpycT2/mEdhXQHtv
2uiHIn4H4zzH+VADOml8ux4/st18UUc3XcAiV2n2X9bvKiaW+Z9/GwetYX60
ov+dKYhzgq7ndAWU+y4FXwowwtClii4XwePVPwfKPElQUPnuUdQqnrEnxg/W
+dOFaVL1nIOciYhrvyU/A371HimaARUhTC2bn4a2r2pRvGsfMm02B379Am33
E+hzKO/A9iMtox2KZ2eAFQux2NsaxrDCEwCiG3Be9j+QNJoz002QJQWV/5sO
NfT2WiDYkW72mpisFIxjq2U7I1h62iGkEMVerdXJLmIQEVCu/Wmerxr/QzcY
kjpYkxJbu5HVJ24IO1K781JWFwRzQBf2rv1DMmS1CMJjoEIRyj6G2HmlaiWB
zoyINPso1sJ6aH+B32qSEBemqMhF60i6zEiKChACeSi/rmY3UmH7+LT4OPsw
KG0M8u/4y270C2DLgpsz/FDhW6G+ucknG1lW1RRhrkR+Whfvqhp0i2pg+P1d
WSv9DvIXNZ5HUCPYu2ta5LWggp9gm9+wJ8qrFe+Lj/DOhjBERaHIOjaD++K7
VGYy9VkysWt4Zd32eGyp9xRfQ+LB4de5dIiaz+RsTEsnbfx4fN0zDzUwIIEP
nmyGx/mlvA90xV1AElQwmb1YHwBU2Gi/Er4rqqpdYsI6XmJD1XzgA/bhPzfx
x/l21ylTYGTAauETA73x/NUIQwpLrCKf37HJiOIKR0qYLNbeiV/yQEu7MqNR
Tw5u/5DTKtM0ERLCXn1pKBGoRIMuhACsWfnETUQ3BRPSCTRtTJZnBZQ9HcPr
abMysZaXsnBMpXzeOTicKpH3oISMS3pyQWuIrlFRQMuwCzmEWXzmLUcQIRR+
GelDigWTShV6Uxklaz+MPih1AL1VBoU8A8yNuPlKDHmeMbzfojXtZBlmHry0
UhZZkYHfSGKeExIeCWhS4XkLN2p+zIPmsb0n3PjDm2Ji0CbY3kIn05X2EHmH
m2qylVbBGCr2MRLZ1B6BQo2aTbcV0gF4tPqnZQrrwM268ZtBM4HJVbUyzo0q
PWLqPrc059ColEkyT04aj1GxG8amsxi0fpgHSKaMOnEnMPjBGJKH3KaQrei6
DCUpNUC3ssvjwaE/FBmiOPaS/B2lpljfnBgrFy4PEm7jNo+LqRZdpIgtQWFC
O5K9tVvrPlRm4sbMnJxru1D/9oYXB1w/t676yw1aWlZc4wwrYz+KPi9X1/8d
438jwXdnU1FSMTgv90yyNo7y6mI4OtiEja2LSlnGKlDX0F01WuHkjCnP76+r
zC5bMCt1yfW9MReqVkuDnL4dU/YHeIbz0Pzd0y6POZHkPXqVhcO911Fzy5wm
WZJkUJqF88uWbz8ZVvPvkr+HMXJVVgAGdExY1msHe4lrOS0Q8+waEFOw5ZL1
o9ZHkDGX58pDCbxkXC84Cp6wTvcB04Eua0OLBLwfOYm/9kzikjpaaeRnQsi5
FJe4TFwax7+w95q90oQNIRlzJ14eDf36+jeSTgqqQ08FPinlhn75Gp9UiToy
vdpJr5U8SU3cKXJ32O5a0R09BnPMcjyLP70vHBouRgVrCR4kxLMNd8lk6hnR
IyXebJSRqxrVMV9nzaRT5Tm/lgdWeqJ7a0hwo4YQvTdciR81fwcN5EbWHIfa
/2GIEnAhgTdflyFYIXDh8bioZRiCQCTy1eTpTE6KGBkznce/sa+fr/jjvrGY
3P3M24Iu+hbHh8rmV28BtOpB3yTGD5LuY24L2K15gO0wbvbfIMq8XPcEHiKz
WB73ZaWvU4G+DplfXQvy8oU//Oz7nFPFaO7zAz1j/SqnpAWcFZldOUFuzuzz
Ql3UBUeV8vjjC4tQqZbi0EjzZuXifBW8lH57qFIJ4buq9qT9dWZBWVMF8afw
Y44sA602lsB/n6vLg0ZhGtnSLZ+IU9AF8ICXeoB8gAIl7MGSBwyGdCypNy/O
0XVYNumRCa5DX43CoRYtQwxlZBYnPA8R2fXyHSFBY8IArKmMwBKUKbjDN1PY
06j72DpTmvKoz6IRFZJ8NvRNZZ4FJgz8U4cw+DTvoFG7p2xgrsBrqXelp71V
kPFlKldPkrwz/sSn153xkdtcEsNljH52r6BKNt+EZ+SXO0NIeLwp8g/Z76wT
Wf7LOM7xC2JpEXIoHJ8S8M17D42ujOuhuXny4Bi9pITKuTCXvLYtq3ubxzUH
x3Hn4++VGDw8uinbJGg9+2hTL5o5Pakc6sFhC8mACbBf5HWvGy+XRYf8+Z5m
wBMY/kCd0MH7XWrMHD2AtA0XUwNKHl//B4UbLt0tf+Jwz27+Sj3QNQ/mnlNe
MjuGoj6zOE3Gn2QMdrd+eD+b+UwM6jqyr2Np4dyPk1HC6+fkG2d1Hy8gXr5q
WqV08eoSqMKsmw0TeLGUJrRtUch5R4DbiGra7Zh3d3+rMO+CHvjNdDgrYvGO
UA5w9yHXu4rRmYW7dcl578q4vqDF8NClPpyfxOSF8eXfJ51p5tXLj/AsD21D
8pSPeCJMosN1RxRWKfBIAXB6Lh1Qi7DhsgPuXBErlpHL/Cnr1nritrFKo2eb
QaaUtZpEs3Eqzx4hoYlJikXc4pPtAXMWkfbG+rMOT9bF2a2DZr0l83U0QZjl
iPHF7N+SLAhvcYDroFe8jwdsqBKtMbI/0ii6p1rGc1GbbVhgqablNXIkwiJ+
wduCGiWWK5VqcvlNz5tYFdwQ6N+EFVD45N+l7yJ+wqCT8B3bp2s9CyQdfj8n
g7LiUhOsc4Oi8eBgBb8BLtks3fRS0M29soPq+KZunjbCfymKZxtLi1aT4+ZB
WKxepjLh3txegROjsN1jxlYfPvLDk8lj3dJ5DrvhNdFLsesjraKy57hnkeIY
5rBZgm8uw+8kc1sfqJqUp3JF6GwjuEDzFts4sd9k4r/W5LsdVDkY+OPceLkZ
xz58Lf1Ib/PcOF70nUb6bf2v06Xk2JY2otCOLXC4VYKjmwhAfFfvb1xxn92H
m5hX28iAtsal35Gz0QuXKBMi3PfqQ/lKPe+lVwWdXw/SttVFBZcI18Ava4ev
rn5cF5u7uXHbEMAnJkJ0MNl81jZfzYTwnHR57VEJjnzucDJYsvr+qZhUdlPJ
iLiC3yYcn4zrz0mY5vxTxQPu4Aa8fb0ygBrRPxGRfg5orLIoABmG6AuiE6lq
uvJAVDoPVixvB59Mb186Ie7VR2+oVQjI6b9d9N0cQH5a7GlTyXLGhZ5TLNz7
h9Gr+Jcy9sUrpOc+W4fbYkDD8f+laWssBHWD+59EZTfsGc30J+6nPDfqh96S
+VJXaXWhXCL+uOFYUMbWDjQFozHAyiN/CRQAHJFPVSQLq3D00fgD9zX9LEB9
5gPjnh1no6xOhlrAQ4DQgyIli8F18VNJ/WtM9AuEF6DF+++o7H5ZiLK40Znu
plB8uC6nr3IOG//hHuS1cYtL5SDA7kpKmvQ/ejb+q1rOTHLHxj9JDfac/gfk
qAUgKwTjAHgdiJ064nK7LC+a1QLbelwcWAFADaHy5oNOCwGU1oELmBGNSnUb
tPyA+qkYRXIfoZY17xO6vwkGNYj8iu0dXuM3hg5gTTIVMr2zGcD+8hZ+fNDB
TQSmjGCMCT8aBY5el/gutlblYcVxTIV60e7KEYMvp1MjVo+wIR9o0BYV1xa5
MrOh1MtTKjeOrZF/MqNoNl2MZPcgVIBvnH6h/rAMz4zwPtlQsPxZg7H4dy5n
Iuo0goRUOxLTzntg2Mal60gl0AgyPP6XSxBnTLRcvrpVX9+wFU06B/Vgi8x/
6vb/ZO0RlLxBqsM3DQ1/UvOLr/dDZ6qPmc9eYhdUK6nKJURU6rP4jd3tHQYH
4dxs4PXvLZ1GNJ7bemX3238ePeorQpyr8RACacBiXoENdWfh7o4UqHXp36JV
qE/xAPLHh4NsKmKn0HjljQis1uJqRmo6sDpzt4NmFjoK1ModRHAIVNDgEMlG
Ca0GV1cTBDy5PqHh4MqAdzUNaUQ3fdNcko4gyOfXgQeGGjI+mJCJWaAXxhwz
xoowfLFMwQX/egehYzm9iI2+Ax0aI2Evdq3Sp3TSQONnWEpWhVmKxyk3CY+1
XcdjNEMkIDOOVlK0RuX9mUcPhZrQKWOAzSXk05lgQP1ipTKSa/24QeuUeOu+
Sv5NjbcnoRg5telwN58YvL/+l/PQ2yGrYkQrDY32JQsAM71tBPkqZpQjAaWC
32Kg2ft9RSt/SEixWhT0jyfB6A7eafYbVDsFpV3F9wBBAfewdz7+lFj4PQNr
+yloKrwbjEpzXqryCYTNOAOhpSzVsgs+7yiKmRIcKv2kzFHb9Oq3FZycsB+r
oyXzG3E/wVgBTQp26XdzdKRKl3PkqgFLJs9ErQytQ4THak1RCsfPkkM2shrG
OiFvz+bjgwlQhOrV+Gt95vl1foFNAk9apSz7yIhqHrz/kUkEG6Qo1YhckZBp
itg+3udQyOq56WKoij1N9brsaWpB7oPqsU1BDkcsumqd1ws9uYBN5NrslFxj
jyv2QprcbT4TWnq6xG1SedsrOkBB3ieWNnvxS/bfDVx9r4iaJ84wkN7u/J70
bjGHxTQ9aXuQSX/mBq+2dbI4YleEus+RoPhX9sWIzvlZWFsBDIwsaMecTMd0
vvcwhVKtPNQYDQqxIIrqVxf1W+/7c7mOWv9zTDR9k7xWfKvKBPfvhhFDYc4J
Zj9wILAAEC/VAJ9mms+/0xXAe3ftU95ICrybhf+zjlpdQZEK2ma83DzUfe4V
Rb7ScvJa2s++HGmAztAQOBF6hkjBN5rDwJ8SnIQuFePWiJqhz3NkTFomK+R6
vJeFSjewkOhIKCnz9z09ouGoq9Zh/e+QoS48nul59HwahKAsbI7nP0fqwjJw
xCMHo7ZuCHZznVRaxzcV9pCaJoPVM/kjhkUfVwVbzHGE2SxljJsCWynovA39
cWKc5Wc2QmCn0yZ5W6UDdAXGnirgAiwA/u4IwPlPEUdac2TcD2zWCO3ZbjOC
KR1+O6dhyhfPzh06IfRF+7pJlW9gaUzamVvzC1ds/xqMf1yhB1/6SxYIO51b
B7XEDZizSGTVteGCtvxokkNaCrmf7phatDH0MAh22p4Pkf7+pys8CODXexkW
FHrMZQutJEzL+GllxUdGRiLixdqf9wAlV01t1GbEdn3ueUGGn+BPEnWZdyMs
T7nOwAT+qIbqT3hWPoxTB2lGb7OjjgCMQy1e/TntGEeJCfVANtbK2yItyd6F
PUi1dioLetKWMH+YcfJXi6HqoVQCT+nXBs4LrJTZYZltdBnEY1TrZuaCcF02
jQAYrybLdylRsmbgrkt8+Kq7koIwMd6TOfqz/aZ9NWOpU0HuoWiB6PKJneFf
DdybOYHzEQ7LTM8vCp0eCmBP6mqas00VRuOKdKnk7pp3Wsytk2Qws62WJe4/
fKgKNMDGo2mJtGV5l332r7cTHzeeyWn69btyqsRE8WmIMzpDvzPyXaHRIgei
d0UVlH2VqRdsvKqcHEAvbAw2Mtk+TNObYp1679AFNYctoyKAaUPNTsUB3Tmw
WqKUZGIczTChy3P8rIeYS81zXe+MbisqhUbiXLXCcpMsthFKs2jZQiDxsuRL
kLih3Fw/2AecqXProY0ILFqAg7kJNlg/b88Ge9LCquEjzqxeyMmi67f51eEE
80d/GiLxZ0v8AB/X7r3L8/ooQxY2b8vvIdLcXVtWL1PF6kpw9STkN7IWSjZY
kMuLxX+7qsECYYjAVasVs9AkaoXEf2rcCrHXeZmnmhZI3CRvvycIJG0qjRxZ
zF546aLgJQ4/0267J9aQ3wrrE5Xu+v5pAcAAm/Ey1iQvKCnYqSnNB2LiyyKa
D0QznCjoPTB7y1W2gosuPHv4zNYTUNZUY/JehLMDGhqW6C7ZZu86ehL9T9fK
lqClqbScJztgtdMRJESf0tdFrn5db+HSvlWBZ7vGjoz2lvziG6ZxzR9+7tfv
zEjO5HnWf8OTdsZZdyQrG6dXexJcgEfVQzEkkw1iM1VanBBf9nNIdvpX4tk4
8aM2Yu8scyWKGqH885iWqn3Tf/AoAJM01+nrnjU5KXPazAWxpNT7+Ls43qtz
MbolQlwwYauUTJizTRKk4D6FvXgYjE9VOxaGJS4Zf76XcHk5ZfGc+RxSAUPt
hoNaUda2016YypvfqAyfrulrnmZcaphtjcsnz3a7+D6xvYhgJsYOE4bol5R/
kAUzKYSUZ4gYbHCjtBEwbIuPVFwyiPn6MS5d+WEONPTO9y/iZbCoIR/WyLb0
bQPl0gdD+K/v0bMUfZEFznjB6N0nkT7EjAwjVPEvDxGRNWLKhBxx7wbDaLA7
IrTgb6GCRjHPHMocEND/+9tncjzkHqux3HKnG+wp04qlctlaHn18PWaa/rH/
V/GcHpO5cYfisKuS/2nP2AmA7/ysCUhPqQr0JdLBgGHPLFfjbA4ORz2AUoMs
1O0JyjNWFPJLyHUZDPS8UqAtTX9zTfofpbOey+FkdpGp7uJcxH5fcrRO8jAU
8ojYwO18Tbqv/lyncTGF0WGns4+17VewkDtYqM23qqIN1wIfMvhdBegKxhSf
wWShQxZ+G4t4CKRNf4RMAs7mxdKzdnT1f8Oc0zfNeYS1SoIrMmQ+seJfr6gp
uVCEpwpE7p6VKP4fcGzMSQWjawjpb/GPEouiE9/xjmkQk9fmePYeILRiBCn4
XmRnxwzcIaLY2LrYsE+dRPAE9Eh1L6/y0Sxy3Ckhq4L8iF6pG4Y31mBaggAs
YknOdlbfCZfJG3jgGMR3W0cJzj/IW0eARCsYBpPIV7t0I3PDUrZB3bza50Ea
xtcsj3AuvdEImVPZQzHxY3dGgo4zRRuyDAPruAEr3GqzmTwmmc4jB41STuic
RN6UpRI0Gd7dKaVs9hnXY3krhmJTGWMF2Q8/O2/sLG0xN0LjMqL09gW9dKpy
1Eg0rykJRFaxGzy5JA/IAdlgD0pJDVBp+/ojLpqqPF3UN6vVqwTXDCUxdESK
ydP+w+Q9EbpW7CwiRXQsRghE/LPD7W+aeII8j27bxiOa8sSW6N0nYOOWaLvJ
a5f1v1XnB/17FxUpz7b6ks6aaYjscfj9rC6IwqY/mhSElO7AyCagjTslk3eP
Orfam4KlNSN8aDTq+1D1KnR6WUN+oaLAlY+piP+BZESGf3VXsbJBsvwgQcnl
k3M/9QtX+2Z8yKv9FmJjeQmAlHO4gfYpb2I7qvTYls9ixmof3JGoWyaVSexe
7TDRaBAovOvdTo+hksosDeeXJIh6tvCLIZlGp1A/Js3IPE/ubjuyou8rQ9CZ
n9yq1pLVpbVa7bZNXRPvRwcjRqCt/sgwA2dNC+gQVRV/hixO7uik+rll9Rjn
UFqiLO8jBK10Ba8kBF2FyZ+zcnMV0Jr0nVhgVQzSS6n519kyBv0sPndi8qdf
U1VsGYYJceUkUbRZlMO8x2xwxaOFVovJxE9miiNu5hYbjm10jeqJMQIkXO6E
fxkc7pR7TcDVaSSLY87HjLlXq8B/86IMSSvPQr1vQRoL94z4yEfrcqeL/LlZ
unsaDCCIYL1zCjdYpY+4liOR/G+agm1rQGKkk0vUZAkTjcBz1d03A1DObUkq
pAz5JuyBTDt/FmmEJ5cC0K/QyxSCGq7mPiFl6XDTPtizsH4LOde3/BGijbJS
Vo/Nb+IgLXP20ujEu9ftFx2hFLDm5mMqxbZiSwxM4Q18mYbt14FoYnmQQEkq
XN2ImH4jessoJz9yP2cqPTDxLFaAgrg1B/ZYBpUYQxJ31ucXtedoGXX0JGIw
yxnMLyKSDl9LuuzlQfnDBxbPPkSJA6AjiLZdxpqqGqfzj0NI4oyn3HUk09To
4pvAnCZuE+74SRXAELNGLimA0cfAOvWKsEIhtr8WbAHSKzYQZ9Xx0/vnB3cd
+FPl47n5yA4TFp/H55dYEWrvyQZ00sqKcAiSYxpmZW9RTChyasixLYBFi4KN
k7ckwLjxLvKKouyOy6e2G0OX4s32IqxUzU6GGixhgW9oMDIyM/jZf5bR5fZr
n/Ve1aH/ZY9S4o9CR2DdGbaDHejGnMx7Q4mt2VbQFQdGYzn0BxKtBdFgeM2f
HaLGjdYyY9suNXfWFUsncfEc8b8Y43qUHLN4bPm2dcLwkjzgK/cbyulGYRD+
OyvXaCYMthFhyWMkTivYmF1bblv98A4B/DFcHGL6k+qoGJhLQK/U7jt2Nk4B
pezHRww3Y8sttsgwucqiVkjGMuPL+vHzMtVAlvrU5aqRLRjR8YFca/xUPGVg
cRput3lpOnkyWnUvAyQGBJeaPuBMhsh62vonF6nTB1dt1hJMjDXYhdoLs7kw
xZh2iN+oGHlhx1xtqGXUVPMFAngkmJfD2gczL05MUbYjGcVFP8dHtBu5GX27
v+b+pmljsFK/1vvea10t/kOdXT07cCp7A5Zi9uteemYYnaI3Qa6o8uOa/7H/
qSxuJdfujlt5Opa5EW6mHoEIq8J6Gq2rP5e3lbgJr+A8S/C9xCpmQl3wKiGB
vpq/fmZFPgddkdETDv3fwDCIPcx4k4zIEw4QBGUy3iq7/TXxBfc2xgr+hd0l
qloZ9sPhUVnpCpJVbR8H3Ssqk1gPuv5HDNnvqxNt/HR24QTBb9sIjpVsZccX
TJ5tqsNRTmwl0/ymZ6URKU7ygnx7CXNUszph+PpstkTJhM6jfVDsnH8qv/pw
tqSmwh/+BMbiHwIcjCPoCVOFEGLJug2Tk4qh4IAYFn45OpFiKEnhDbJi06np
m+A2ycdrHybtCufOiQI0zqwAvMZmQ9AwJIO7C8ZWme1uc/37bsZR6nkyCMWR
vakpqLctMWvuyxX56/TyVoI5wcNBMbivgqmzDygJ5MnKfRD2RSWdlB8bLEnp
epkJHAw63ZozKln+gumJE+CNFhc0T5SI6HkBTPoUW4koKmS1VTEau1x0iPR6
XHC3E5CpUFCoj0izjrdGF+3tScuXPGXmKyMVZ9mPH5RwRlbN1paJSI8Aljtk
GZTdZ85fty87wTmiDvmvJcFhTLOCykH+VepQR6CdhPstbKpaaXottNXxC6+0
wFQ8aJ0kolZZ9UKyC7xt2HFV2xvNMT0vW4CqtAqhHE9NezKfzGDLWgBb3ftT
DwwYJtMC7LW1v/Y/lYvC9QwqhezKbDxZIfqbggDcJquSi/z4rM/yZgtoyfWC
w5trRUd04oWYoWwQwJzUjmrLBoX+x1s+XwpHc2tMUEfyiVwWb+wssvixotbg
Yw/xDo+QVL/rFgsYJ8zNbi6P34RsxuExUUFsrxOtNPzWFpYAYXlqac7n5H/c
vWBXgfL/jLrZzNwfrZwfQUUzHgR1DjyCU18d9kv7qwpaPz6QwBoMoxjSxNCT
8cU4ODFpLr5AVJpUdrtGfoq0RTwCieM5P+YHMS/HlowN9r6tGLdeL7WE2tJ2
6xYVnGLcwjfd56B0bKqg7JurVFGz1Vn05l5cNLfAe6upJuQuRd5xVOHDUNUV
VSW7OUFOl13hxI9TwJKd4Fz6u71hzU2CCROwpbCQAxTKi3KztYYerlx/fD/2
5gXznVRw9veB0yMTO3ydjbN196pAzqoyxK7zabG8Q1+eMErw58IMn6EOYw6d
hxiaAo00qi2dDP2wuGMvr/8/noh1ORI3uo9OQkxtlKNk0K3vd6j1kL0NyuWp
eOKgZ77h4UVkpfCQ+8zBOFpcz11B7zfdudWZM4ogv7n8BvzodAaNOlYJ00dv
AIHgMCTtKGk9HWgY9vakAbZ+zb1y+WY7ErOARYyoAvLMEbT+SCAYNGWCfCoo
p8C89IEZVb272CfSXxnVj3pnLVgCObG+SA5A9oq502twBbfdfEDUKx5+KII7
QxNGn+yVvLK5I0Zm0Z5QWt02nsKIKJbW5++iwywt3hyHqKh19WJlY/mH75rF
DTVnaWZg+tO91qtRKF+r6o7yDY03QCDcmBD2uRUWtzPYLq0cwhZPinlLFo8h
IxNNHMRqBu7VwBXHKdiKMGS/PUv+uscbmnNjpRjecEyglN/ooIQGR3LybrLy
gfLjluZF7kULg11En6W0knxoXl6ozpcyJDt8u2YhyF8kHEm60YQ3GHiNv6Q/
4u1krNJG8KX47e+/hBRuP8VdxOq4IxplLlJkJDJUhE96ZGGVOnO9PCP3WNNb
pPgyCovDA2W1jEvFnr0vA5FlGfd+d/Uw1sdNcItVn68Am4hMZoHADRid23YZ
eIaeXsQDOqwWArYZ7VLmCT/xkQ29m/OkBuBJxZ0WhTJZld5FqJ6365uLWsWC
vboAzjZ4jb86ksrnr5iQOnv8Pim7iXE87EaoXp/4S3touunYUguwokTTMtQk
TrBpy3Ju4DtG7bxVUARPnK7KWOy3rW0VMlPxvH6DRYh1v5yFMhb+yjtlXQGv
8qzSdxZ/WbMoZ4Sc5Ub1lY6dAE3JHSrrRRp7CNLwl56IHllnr3Jj5EOAb3Jo
GKjpDE+Ay40GJCgcWyIlsxC97vIBneUD0dgFu0fpuXkeOTSeibeduibE1EpV
cnUL3FLQfwbAZx8gektFxOppOZ+12mJbRO4Uy1ATulgSBxycNbfJKrLamZPj
qeopSSNoasCQh09OqYumnHo1nPls3uh/agGMsgxU4AWAxf3qOo6ic0txK4x4
MdemIvZ2cwy2aN0aoH9WxD72wzgky2Is76RGdqe8uTgDkFVrngx5areH84K6
3RZmrXhvMlDu0Ai4+DKT2YadkbzqWGKZVhB7n9Py6V1GdM1JDjstTNln+atc
4teSIGkabrUKLVrkScBTH2L3hh7eqq0rRn26fdtl6H5Cy6PCsqbSn5iWl7Po
J+oq450ZLkrWO8W+mcdk1WDzQ5Qro2cDCz1NWUPFPe0HOi5+1RDT4HjHhAFX
CWmo9UwbGVXpbYFPoHECzq0B7jJ9N4LRcy36KpfkpY9BSVbUGl0vgRj/ttKk
LWX9tcC57W4UBh1TFf5EYFGPHCKnrrKymMqaQcDqGcibQwZnUKdDpCrPw0Tc
xdv4O7vhBr9SEDQuoeWcP/pzDAKxA3i332NxsjGLZlGFrntCk2/FTs22FsA/
kiIH4gOK8TsUAp6RT2nOuDkq9I5Xx66VPLHS4t8ROnLAJSJr84nqrLPC3ERW
LsYXBHF8soA2U6Mn6UgMeyuyUqUr774/4acgMvbmOH9qPiNyQYAw+HayVPLj
MCl+Ws2MOJAK+o5QcpiGeEFwOZr/56ymUj73Ug3CpbAcTH150uIFV1MXBkFu
AEndEaF2bYxFCkRHWIeXe0P08Ckd9Y5Q7pE7VXVFF+s8nqPot4s0H9HW1lt1
w6nwIDSFkialRdOu3WGm8GjKFiV36HYag40RKQA3uUN3lF6Tig7g3zaaca4x
Zdv2xlVFnW67pRZ8CWHA9N1GdYsyKns5JN+2V3E1jb+kMhYkMS0SVMcTgWSc
B8PK9FtHWkGlW1QtKbVoxz9aDKP5h3Vl2HmCRK0gjWc31uTRcE8rhhfRT5JJ
WLe4cHvQP+A3UT6r+FgIuwpv7bSi8y6nq4ZoM1sJvLG3DgHt7K8Ck8OTo3k1
HhCkE1IVRtS3H/FbDKUGS2wcj+krI0o2+0l/6ktBPCA7Ms3QH1PpHElnb948
hOLE17nDL846Pf98b4n/lTEbFyKuc/uCgOPkTnN4BPy4frR/vsbycK5gqNBp
g9VzaRWPE7V1E5+ipszwba8wQYYnCPCPxdKxO9KQ1CbU/GVW0NAh78Uh2/Vv
mTOzOe87SVdaFZHCmIb3qzpeXZoWOrqsJ3/ulMHUKfB2oXjMaXh2GvrhUbO/
HAvsPgflzYTzOJc1o+uvbibBDqmbnhfIF3wClTy3ozdhlOfmBHQnEgjjTz/+
MDmV849O4DhozYaXMP3BNsi2vLrWTYYx4ho+uqHmbTF287nPEnHjDw7mimbN
zPkDDSh7oaRlZnyNe2pXUcmT6Dm6uGG7lqYTM+uUmaoRo8nArOEgPRxVkWad
yo6lLVlVClT9XWoVFXdAocAq/lZ1EEk7kv0UsucOwKEqk5ZmqDZl6/GQVc40
Zjf51WPJDOU8wKV4ayDrfzaSsLisii9JULxP1ymRP0qBKrGVmkTtgGmJ7Fow
uN0Zf6QB30NBeH+LwSdYkupm68KAE9JA4q/CJM3RTd/16j87dhZegxtrvSde
+fDzL/2BXOjX81jTH/HDwSzr4+IN7xKOjrgMUgPhhgMgEERaU8AnwiflNT2i
SliZ9GC6a1MZv8/3H2NSrYIf75oIQGY/ldBu9EwC/8cQBaIV4pt1mg77qWXN
J8oXm76RhCWKBUGWwUx+WjYE89SGUDkYdCOSG0wG1VxnKCQTk2nd2WSs8z4w
YhtRBtVQGUJcFfrXDylvBp4klr6zpU4Qg6pI3sU1ahIRIdV7W7WUmWC4WeC6
QX66F7/kXbi4WYeCtoV8CnuGEdPC2RWn/fj0WzcxCJ40AhPVVAj9LZW1urvY
f+3ovaKDsIt2vcZfxhW2Q91RuywO6eQv+/M0+eCqd7r6lgYHdkecj5h+uNB6
uEU0UvsU4IVrUgMpw5iSSbQL4TpWOrb8AplIOt+LXeNwHjWO6Sp2i+LaNh2h
v4ZMdul0tj2KfXyM4c1h/reXJwOvtPgfhkEN8mVZZQEqtYNc930dVzMm2CFW
yR5Xk1yo74KinaX4P+4ICcGjEfd2azqirHLBPAuNpfgPsv2W+G6DVGGvcFGP
ataEeRGMxODNGwp0dui0isR9drrql+7ZCiGkUGplbJ8s7NjZrEm9EBadvUtW
09QL52ClUMiDvM16e3yS2ifhl8X2/XPJgNTPfGCAeQI/g69WyDiUDDD/htMK
Fbpz4ESmjmBPLvQTk92qqtw55wolea27rZFoEsIxCpq6D1+DkA6JQ8OzMETC
INF8hPJ2PSxiPC10kNZj/q01AJ/QugtXQ1TTLvt7kPYYT8n9h8LF22tjebGC
IFuGuRLeTeXXfptrTe74nUXW8SNyU9rLY8hnSEMcabJCiS0cUPY42Ju98eTf
Yb0j0mdCPEa0Cs+2B0jbSsqSnb5GOMTMV7VYy86GWdcRT123rVrxh9GFAxow
ACmf9+UUdLp6TTpNDasecDeOKgmKdO40eZq6dnBkUzxBrAVDtVpxvIqAoZrU
uL6XW0WVEglJjkeJI4BYMGez39tS3ey+MTZ+EvyF7iy8wJAtS/rybY6s/T83
gC1bZn9PiBKhMFRa3edBgwWEz6XC220JLHaYxVMVozXYCYJZIuRHVUaEfY6o
fUZmiZ4vQI7S5G5AmbhwXrJrjzDalx0FsDAyYxzhxUELkEwz2amIgQFyJ6he
uJy+bh2XFzN0oxY1HbkVfCJyEUGFZ0qWXkZHnXs2GVWcukzfgMb/HtupdxCF
jgpW/+EOKGp4U0mzFd1H3/cqrei7/ZQRdRfn5+fopvqXvEPzVSRm1lsl+IAs
aomv9aJtmeYUwHyv6tiWuJKdy6c6V8GGB7iS8KmZL4ptC7dSbhLbRCwOm1kE
KtmRmQBntp7Mg8QN4phtVTve/xDwuqPMaMpaz6g5EiKAkMCm7WiE+4Pa/4gD
1dq88HA36AI1frN8cT5Uzv/cLVANgZdfNxZ0tINn30fDpH33MtD8OTWAMQxa
hRraFMBywYpBvizfkl/Hg2Udp3baEiw08GaTh+CRM/N0flUeDidZzRExAnmp
bHfH2vjA8J4RXsfU8QC5obyhqmBQZ5gQ+iZ5L+0r5CIx30olsUVzHuQebdIg
0Hz67LZ/rnss5Mw83shZ6Q9xblpgti8dJzWJKAomj92fWmpEgBsQlN3R1O0c
Zx9PnEGvyQ6c8nhtqtMGXWwlh318TXypwXJRgRMIUoAV8VwltCt/JKB0nfRt
9y67Pt7h+bQZoKBojOohRDspC+zKDHigL1446nFCGv5r+x90An4jw3panR8h
TICAiFh/1WKYyDepchEvhe69si+2ZIHMBobwSPtSm8LkI1eIaLqxKgkaTmcf
Yk9GscsxRWwOaTy8m+T1RrtXTS4/PmkTIIzeEubdkXRYk8UhQFaXGWnbD3t7
NCznPNn00RDUwdokhbbwaxABzo7KPjf1u/8W38hrQTdR7CssbkNBo89GoItB
DkB+pvhfq6cJg8eum38WOStNL73HV4mAmzWTGkrtnSSYO0dfyzccOaNlIMMk
dYqm1o/pX+GQJ23laiDdNp5PcT9PN2uP5yakq0eK3ECCOp7DRKpwwYZvwuXs
9Ukm2EyPL/fkSmptEUsdY3/QAB7tA71omHl138HmxTZHFnnblSw8GmQ6vzAp
ZSw0I1ft7B3CqCHmkH88doz5nEe220WLhJOffdZziDd5BDBrrzGt78EIZY4g
ehtNjnAUQbO3ErDRLyOZLVg7gRzpCVH9PJSC1JXKqMjpyQ275u+hMFFyKLI4
GLuMqemxk+GTxkHLzB6IobXNQrkv3L57bB7CMpCnrMyfnDhq0U0ySVug3kRZ
MvMPwIi2Q0KHp1S26hzGEKrkYZYi1rdhbDTLKJrB4aUb9RG0klmHRPpf6o/X
q0VPOgLD9VSJ4b5u9uYT0G5DavNPqOBBEJMcthY/AR4bUY8ks0+eeRAtuA53
4IisC11PSkesOKQbG4p44pIk+RZLptVtP7gIsUxVBKbuEjpLag6a9mhSAYzW
U4mjBw2ENJMZb8p9sAFlOCrCbxYGS66czyPZ7hVi6kU2hRU8aJ1c/shVQqiP
TJDbECTas+gLUueWfygDw8hULY65OVTN7fRTz+wBOS/JCVBuPdXxqdtzHo/E
aWlYrPO8sbb8xdxAc9KcKQ0+4AZZP3lRImCWaqp/DFHZ/VSb6UYfbSYAIIAm
7pSpeayw8yrgi7DOYvTTdDkelmGosGODkgAOHum1BoMHk9gF+8lkZ6KyeG7x
TIy1hltbwUd3PI/B1uq90wPi0uYCBQ2Rq7W0cSzd0mzl89LFIBOaDi6n/9QO
v/g4P7fqMnAiCxyqyfGDQ/OhrSqghZf+GWQ+xDMZ3IlXR0g3iAonRuvYx7cU
0m8cAppb9Zbf2o7xuq8MPABaz1yrJG3+UAdGDeuUsQliNVXGo1oYc2cbisXU
P7VvEzVmwq9okwnsJ6J++mtfxYBmbLJbMm/kq8XZcsK+WtWq7rGCbkL6kGzT
kb6RI/z/WTi/8DN65MJUAFBNdy7RSr2ct8FxAmTfn9rfCu8SnAUifYXahFc8
RN/TxdMpL/hJHiXue6cembYEgP7ntIXVATs22O0RjIgc4HHrF2a5ehFqwry8
+A/JTqh4yYrj1jSk7y7IEXlKJLOIM4MjgMlQizjYVHkqCQ19sF0XX1+v3zFM
P7zNWhKlu/0nEtnpP8V2wQEBqIl3nbclo3sBoT8PWXkKXvk0YjNILrFGVDf2
MrR4CrT+MmeJ61kkLsE+Zkw5QHjrzT3dV43ljRiUHZSlsaV1WlGfhyda4oM9
FugoW6bMXC7L9o32VVH0vQnUx1uEVKTQlJvnD9FbbcaVdGWUDgmisDlK85zV
sDZ+zh+Dz/3Kf4hflBdnP+rLfkORonD2Eu5pwabHoSe/0NUMKS7YXoQnhYDG
lhDeoG0nB99aFi37NGsHXP+RyXSVWdDj7UX4oQWFhUpS3qPSLaZun0W2VcBk
pa8Np/DcJ2LdXl/+cGbOugJQiaYVGWyCS1HJ2uzsyCiqR+brX2x/iIprMQiT
/+Lvl9ptdGsKZPefjfxhXi+C7+2GMjQ6khymJuQBjGDqtT4xpRN78TZHbzyI
1s35AKix/3ZGD75Seb/g2psjMzTutYvxXA2ZjyJ3IRGs5utIrz60xM7bATev
ThV/2PvbrdQ+mUkhl/UngJRhQHO/wYOmxOnoPvEyeydHiDVrfkozajQu2s3k
cGPFLak2EJ5xLYrgXLXnBAJgCSUfDs/dB0Ng1BKvvrGN5B+Io3LgNx+2jG+C
Nhz9avBdlQ+9yeVXN4yo13kqOCc0s8gTKIR/Cdrb9fSnxIjpry6IMJakrdgY
2AmSvA6AAh1vc5QlFDltVpLRpZQKJXYWbhlH0b7N/RZlP+jP+Dl/Nr+J60nz
rAltIliG793ywzINUEzcFhv/w/scS9TJPQcSq6pWevPQKq4Mb+Bp+J6rEcyh
WwdpKf5GF3ePQuUx4jho7N34j8O81ABCMnDzhHSYvKGfzhvlGzx4hpC3TUbq
Xc5mZZo6+R+uhzCNDOhlDQCa5l+fpGrbOPsLFT37jb46oa0u5N1jLA6tAW+C
w0s3IGrATP5h6Olys6DCtnZdpgDzKkWyfzkN47DKP2EVnRgqJo1KVLj5eIhR
uRyrcrLEJSRkfj1G59kynCLWP+sdc35J12W6OzsdqRTfW77iScpDM6LlvXDW
hgpRiZWMtkUuW5B6oS0Bla8WZd4OrVPhZ7y1gBzKAcxUGfs7XjXclufgK/Cu
cSikVJ9EEqPrObjxldKBZzN9g42VZ+ABm00dpRtl9aNTNe09SaZMM6VhMR9r
k3fnlHdh31ublnktPmqjwgc5UZRUDTJ8QMU3AdqN8VP7O2qNC4AYwQ6Orv94
7dXTOrLJ4htTdh5ac8BdRFDIqbj8gkyLCC2mqJqdru66RPI2Qi3YIkTj+yte
VWMgaWTbxF1E4qI4zxMuHhwJTGf42zH8Kfx6m8EnbfMy5YByHYh/0JTABLCi
6xcGEFBT93uPd18H87EhPHPSmXKc6fQloqZZjt1bc2qaUSAFXNb0eaFBUTh6
3wv1GZj7u7n3u5aZrnff/hElY6ySSY8iZr5t9RMcHxO0eVfoS/seQc3MqH2I
de8oCkipz/fKcwWW4A5ezHX8o5OhDAGE+h6pbwT+nKr5RqflLAIhufEu2B0c
64R7QBZWvUi65yL2JXTmLXRUYv1iSPMQ4+dKhYex6gSs9V2FAVl0l9/ndZ+z
E8fCsXl/UT8UiDYaedwyPXdThrDWVHPk31nqo5Kkwd4qTpXY5Pmb0GoNNUsY
qHFnhNKL88PAs7pqVQ2+QhL6XfOQzFaYXdMd79Es2BzWKlg9ikiT0XCuzGi3
V1yABFSTxWehpw2n78UaSHR8cVXBWkv3dwcKitK0cctkE9cNn1/XGQuNQrZ2
3E6FUjvS2nd+EIe1yUuAyeZh09L+HX3q40UHa2oue7Lj4ujzmVFizt2br424
3vRGFjv2H7zh+AV5RX3uKjyft3d0PZvnF11IhiKfcp0dHvpKsBPS6vqs3vmP
v6xSFlQxETBXs4RCYzTeMZPG5YLg0Yh7Z3rjLbjHbXU9CMT2wyUiehXHvQic
rpwMqgvepjOwlBQC13Gwoey2K1ak2/CXPGExOD8HyT6y/5dcNucjwPpqX+gZ
jhDkhehZhiYNXBdA6xNioBE2PC4j3vMoy/LW8GyZ1UIgikRO9W6hPvevN0C6
cVKromWriMYxBN0T5dO4IkYFBJ0Y9mJSA0XwlXg8mn8UKRUrJcAGLqaKNztX
G6zdiUGQUn698WcJ2VGMHRv7Qk9Y7T+ms+e1B9ou6+grJvvRkoW7RGu8rxGu
OuSuRMA0fV5OedpYlPvf7kgz5Z1634YluC5QqfK592olk3KgTBLstQgRyVnM
6NodFdPEVSxBmKC/dK7YGHSXyQYrm2DWsgmJrniB2P+wYQHLRvMQMAqAD1rW
kkCjlFB3Q31WYfnqnDa3KaZGgtwtifjtwmwVtC2axq/iRNsoSLvtR0JVhzPt
Qm/zhBK3rYhPdXx4LmVCgzFkBdkfBj8iOSMhm2vPZzq//t1GKAu/dxyJUhBU
5866FsQ+1lQQYn2a8HeJeMff5hHCrPL1xkgjXnniDSuh9eNW/7PaKw9s+H9K
NXSqR1TemIjTyLS7s1w7F2SChIxTsTBskGp/7NaTMQCDU2W+jkR0kU0vWIAG
vKt5PAWFMeXlWzP3rNhZMiYmJnXNUWCDDZUfg+ONdU03m84+QxjDjX1YWxNL
OpD96L1j+k4qhrGmuuZx1ft35mZIOsqiQ2xvL/6p2zXN4saXDBFD52dq7B4A
tmEVQTzeVU4cZpS3ws1gbe+CpTEsvAbD/7Lg8QlykJT3JaqV7/zodq4JpoGE
//IVwv/6je+/m/GZX2XYs+p5hhMD7MlSmvWiEq9kQZYL5sZVM10rYtYhtzaB
p75rhzdwtYWyftUdbVrZ2AlP/QzpQ7VSOwrHIz6mP9dMO7P80KkeYai9e65M
Z41eLn21Gzarey5GYrpjam2QIvX7r/oalz2SCWBggcy58JRWEa6BFVNpO9bH
3PT0ILd00TFFuFUxyQ8U/MM5w/RysfV0+sXZ8SYm+QE5DysmxH2cy5z67yjv
+V6+2VDR94mVBOk9RdrqWA6pVacd1KfzrAHB4uvHRGmxEpQqyHcqIjJlZA/u
XzO/I43BcZjiM0eg7py3Ih9AxRy5Z5LLbuylGprpsEn+f8aBBf6434M61aeo
ocjdHckeY156CbnV9Gg7s/+Gx+1ZvAg7Qe9FWIbaGrKEDT1V/nfkec/1/tFv
wMixmLtMicd2co/lYuNA/d6/3p2bGkg5cST1SMvfG+FgoAyEapsoJnZXRBL3
yYdzk2aPJJV7/04tlUeTN/wJ7d2fAvAp8QdwZeH4XfPA0bK9aKvlnPelvL7q
q0cQCCg07Qao1SeMYPIRKraHbWfWbqdcrP9skSAWv7sS+5PTkDXy8Ekli0mE
1Bq0AXyTTODpECyhH6heRf6Kh+V1bmHgYJzMEKz5FWtzE85fIrzj7WpMSit/
Dh45rLi57oDmTBUH3lk6uvqUsV5nO3jrq7ykefWWESL+cJxSc+0bRr3BMAH4
CHuaHYSeonf89Wkjmn6Qpgre9Vhi1YWfpTeFHm4oZJ/k73RNVZZD3ZHke2XH
oPyVTdDti3G4//jj5BMV3dNE5Io/2mfpOGnlBfDOi64Gamgm94MBn6WGQPOH
1L/CtE3qrs3udp/4rw9l1jM63WgyYINxPgQ5f6lDc7869zya8V0Hf+nphtZq
PeVgpXvzP72bRnf/0cZVyAPySDc/lzg8etHJoYqcnaagbr+Pk9lyeXSdlLza
/EIg/ztuoKDFkrdyZcKd5svsDyepQ0vH3f5TY/hU5rWPqxSQGcO9DmItX/Vm
xQVT/501qt8DiC2n8HKvT+YIZCiPFC0smk4pFwVvKG1lkz+x9LUJadzRQwuK
XYDkqXyLjpXC0tfuoUdxAzo2RSyQtp2usM6LsmxFiOQm/wh1bUpPkY4zPFvb
5fxQ7q3FHJDjuVVl/z3+2bMnAjm0H8hIBJyfu0ssUm9zxm2NKSUGGiTVriXU
a2kC+Emvcz79DgtqST26lljevjn+wKibPJgVhemYKRqGgrtw8TBt8H8u0Mo9
ivyLO8N41TklcaO3N2r/zAVO5+BOYyxEUDKOpPOB6WyofWIE4UxKYcyJrCte
1LdVoT7pLJ4DiexZE+1oDBpGPeh23RjWqzjBVXmbqft29WU6pPYA1TI3qBm3
iKpky9oVAvagBkGOP5lDr0r1/m+qQzO+4WX7Se5tM/DTo5riihm8lkNBHKW7
YK6LPCU3xIIpa2vDQ7DeE+uqdhhoHsUccrMlJeNwIXmA1UhlN0hHlDud+zZq
e5tRbJC3t/mHUMGHyrkoqYvd3hrO/f1bdx+mihO89VYIh36mHQlA45yonVkZ
WrgDDxiLUiICTqzE+98+FHJFA2T1+ZJtBW96v1sa9d/+bp5EVhdeWXLSqBIp
NFKqxZ1sK7ooOxRaC/r5N/jNiAC9VdKsUPgJfBRaJffkfOkHAXCmmzYiYydI
pqrKM+YR5/YQw/moLeHKK48UTtLhMjeG0xaODVah+MVYHb0fzmmrxV/kn/lw
flLMaOLZuC1VtN4JCu9gQd8RZrTMlDxfCtjW9IMStwoeYrhUVgsysWfGOyvj
JgiJd31QsvA+jIcFJaJVwiByv3EezEaOg8UwpFtGLReSS96cg1OULnkdzsoW
czg2BdnTmq03Xy0dO4RsNmv7dMOXgNL7ugNJJgR2JbmW/SrhI3b/1Jam2AR6
+OR3ybw+IcHTFjab7npjps29S+8bze9AHdVF37UED8SaX4JQct0pmyP1Zr7k
Own0qwqLUJcfG0Ot95+VpoCOxsOsTmLluQnW0+XFkYqqBAgSYA5FR0uXxdzV
5rv//LfbId0HdUnwHM4fVC5VCGp2BJrajzcQzqMyTNo3lgSjvseWucNTNW2E
s3o3OE7stUxneObw9PTdVfqnClwDM9a3RZmKTrV8WTVNeJRoXTmw6IiHR1J6
u0RKeb03CEmxoF7f5Hi3ptmIWo9n1ctWMcSdD7oOWnDMft+79KRk2eY2JIo6
WFKcaVhNjwY08RIZhdQTVX6TIM5Q2gOnaAoqobcVs/4WgGzgE8AbtRGscQCd
hknoSFmSmmy5H+jmOpeO9BiYCuuLjyXE/eqN9wNx2RgeWOGwpp/QZvZcSCNI
lwvam47+aSKl/xFMVpP9ndmSMk3U+arzY2otjwlxcbapalpbMYhF8CfKe2nr
sjCtirLERxA1B9bNxAywL+gFWOxlhyv6jP6+2apaUpb6mpNouZyaXqNw8T12
cZtorZYR4phSzTcWaJtnePNI0Ua56ODTUoK9hAGtMbTTAtGDa4GiP40Xi4WQ
L1Nah6I+jaEdrcfc7+hlh45dBRTo9qVm6Me0HeW902ak3upCOfGTTQs7WSGN
gq6BecH+c6WHdjyLwAfDxjXq0aVxMZg6Itj+gs1oga+2YcgsPtV48IWU/dKD
Ih3UG4jFmOarLMA3Ze2jDQ7amhTNqtwJJ7TvxKZ7sLlGMJAjIHSzOeroTV3C
BR57q1ibcx2AvXHE0BKTlYUpdHU/GGmTlsgi77OtGCgH+PPNRSWBFk0O8Z/p
RYtvHfLFWgoEuOx3gDtJa4WjqzvwPzJAf4JQsb5ESLbto8OGM7umfxiD4AJv
auIZsBdn/8EfnzgapLkqUhhQm8l65J50iY25m7Fjr2s5InIwpbJWKZMy/uua
RJMap2evxmwPL0CqcWRRzO+vOfk6sxAfpA+TrVl7Ow8/ts5Ah7PPEDSQ+77F
2JdKnrrMOO6IqlytP1gwka+2q7c7wjK7qOiGgUXpenyl+X/MiwPTxg8hgOqR
CC76wfZO3ng/plBdmGezFmCY99SDkw7Tysa46ni60jtRa130/wWIJ9v//ti/
LpsoIis3IrMGe1BRy7TDnZ8U3i2s0V1uHv2pv4P+dMhQgwvmhIYeakurwDl0
m4FpKtot8PxaktCYayd99fuVeT+Dr8zOny7gwS8L8TfOVOzcjoYYf9lQ4W/3
63kyxyv5wgSZxk811MTWGNp3ivGqm+tEjjSZuY5pw4dtqWxGUeh0MnZFlDHd
RlKRodwyMHUDIXHYaf3LNytmxv7eSxRXnJcuF5Exih5F4YSNkCNINUq7SwqI
IwKJB/Qkn43G9+g+oiK5kg8YA76yxwpnWOM0xHHCbBGhcnD9BJ4OvKzeBk7j
ASziRss4lr4kIMp8VWPyz7koCjVjrV5loA19E6vvvGHi1NWzgjcUG0Q/cQ1e
yhT8X95OoxnWso2p5Mrq4Kwx7aQ/Bji0JaSTT2wBrhO9r+G8e8yWHq6GgBXl
8eEGUMo0zclLtQUZKqdbXHHE8GFw+wmU9ErftqDEF/lSHH5lQZuYz3waYJuo
vyANB1ddO5vdj17xcytWPjGfNMi0q+Q4OHV+GMh0k94WaQNBNGP7ryTgWW5Y
yS9BPWhCLcrxad/kEjYuhbwS30nBGN8G/oi+UE+bFeqTm5ssC6pdbwJ88NAM
mN5OuGvviWzoCpEjfU7n/ucjaeUZLLlNFnL1gbHcbUvPq4VtaJsp/5OPMjXX
SOFqgi1gAFi+XM6WzhDYcot8kj0fK5kAB+1wDDueXjibT8c1AB2K1ZjQ9iVI
mOmP0X4iF1O+H+xbOe5cghkajqIa+XseB8OZcd4Zm9P49IBBZhhXiU1h/wAe
fLKX7ejVjdWvn4gBelfzbaXdlAAKtyDv+GJoJnV6El50O1vs1c44M4gLmURM
oJyd8YAKlGCXLl8d8xfXansbymBq41UALTVUfesr+url/0YHRvvib+VtrtpO
LbllvgBfUtjp99rwaPb965H6MN4EzOcYWLhyS87RllDnckp+y5NPcOwWkuqn
JBC13RErRc2PVccCT2Hbb7dPlQ9xQ1y8ki2ui4sffb7ELWN6VAjnWTba3H+N
E6DTCyNYEl2s1eG+pIdVxtqIytsj+uV4ossVFHyyTE0d6puf/3khZXu3bREs
/nUwuywuyyhrv+l0pCJ6s9WHST82m6/0ERrFgBNa6j0UqYmbVRUCOy3FAUAv
qXDepR9n14fI04rPyu5PFJ62PUaLAipLT9/dM4p4tJkqI4OuGaTbaCErbvEH
4v/Brm0TkpRD5FIo9iKuI2GiL6EPdxD+UqGqVv4q0z6+1GFPMRT+luXn+Qgl
kitKOXgpiErSLlZeTpaijC8F4Oz48HmeVV2nGGIdzJmi6tM17yvNDJIYI01G
zDbVuoKD5oKBASoPqkkW9O49+tq99SrSgaMAOBIz4lscCX46nhIz0NZ+fknB
Sm1AQjW0t+JPsf0hKb/iCpFeb2MM9ce+theD0aEi03qOik0c3PptXPP8tNjb
qIjKDHbOs6VU3w9iLnJLMU5SpDmRbrz4mICZUPPjixYqDpQbcdisJwf3VnA/
Njjg5S2PKhJIelmQD2mjNOB+ksDe+/adO93tV/ROGAQ6QEubsLw1UlcGAAmQ
Xk1SyODzJY+Ycns/ciefk/yrZprl3O4ha7/6Qx4HwOo0bbhCp8P8lLjcZj3E
WgAK9dZPM7yIouQ1UA1fMlwYy23xpgpRDQUKd/Yf7CcIpDfCmxzpIvlKUVRO
dSbzHMCxNfPqe6sALmABdst1CSwpLdCf+AAWwH80ivXTONJlK1UzZlfhcvUn
0mAn3fd3+XnCgGehqTOCc9Z9B0yUXYp8pZj13R0b6MfqkUNOykfDfvgqpc2E
L7trBU/0/wibT64is1K8yY5WcNpM7UeXMjwebmaYAX7Hy3obBlsMJu72sfV6
7n/lW3LmMbaAC6u2jOr8+wnwqO/y5wXDOv+nxdyOd7VId5gKcUVpOc08ZUC3
YArC6q3k5sTy0bgVlvbxx2HmQEHhiDhRfija7o+MTeNjQ7t8KPWtlMRAp4qX
r5iVPjInAf1xECmQ91vi9obc1vMQHq9kESQDko124aiK7w0qetifYqY0TgNG
eq0CxARF/qWuRx1r7XFrbmFLmXrKUuC5xj83Rah3PhCHswLMZB/5cKMdUs50
2TQ0JloAaRx/smCOY3/pGyfHEbDrJZjk13gC67Y1a9OhuwDWeQMJrUzmwGGG
EiAXMy7R3vHeCaxbJ1cCqXSb8lO3xnoJtezJ6UZTaGtbUAiVjeV+3hTFaOIt
dBgb6ccMrP8Zfe8ey+FSMdN/BTwVhRboxZ2ownJ9QAsj8Z8AicpCe6zytowm
suBYTqM/K5GKXwJvkJNwWnNGpM7aM5DRvG06KBApQlmJWWfld09SCmlHx2ty
CBwxGMkzqAY/77Mb4zKCDLHagUklsbja7QaDV6Zm7aN34sSLaiv8JA+UYFiI
HjzhMcXB1Q6P4LP4KGmV+U+dPPQb+lRELznVvk4lPO1HitbfaOmC6AqKsbR9
j0h4MI/InV1TvsB93J+kqosbrqKJIegqk685iFOhlq4a8iVv9/ENQvfOhAEs
POnv66pUlUFlXFqtw7eXpgz6P31f/o9afLBbQSt/x189xqMPW/QJZw+QJTdN
G6FJdlTy7MlI0lF4vYCRHzRr3hx0OAHSr2PRrd5xAHpXZkmJMWv9N7Zgx2ZT
NUQH1Aix8htVQy8JN+fhURmtFrQ2ARbC0WZBJx6n5hZSP+fEYRT8veMyQsrK
HKPOQeWDSJuvp4FAQ7yVRi3X0dxfYF8TPM7KrvAIMAy7vipMwtIbPAu7I0yj
bsuiQ39ScgSKSPk6v9GgaMuxPymPKQMm+jEwNbuIALOxvF4nyFbzvk/F1crk
Lj+ey9isYWWxJM/sWRDRWw/LrSMafCMkOPt6bgyc9jCIUwyBQs4CtAY04TRu
27Ms3RIuOQ5hqwHogLEC3O3m0oNz9FrcmFVRHXMaJVaXQO+Q3FeGJKyWlx7/
4WeIb/MK/cNIm95yTCSZngfWZPPL0XSHUapRKmMZQju6Oq6L129azCe0bTXj
h1Wf5MalM2ZGU+lalJXWxCwRVCagm5VR60A9y0+XuHHsCxl2r3qkbwmNnk2w
f71Jt2XIy2h8J9mx7UoSge5uhYziKcDEOqIyx9726P/ycTiIgCCqCITihjMB
8P3rE3Z9/ywux+TKyqSvAUCnBldAIiofVfpHO1+vdK7DFMZq1e+h5x6kH5pc
OpwO8pUwjuKtUjWobOXXbYdRt5GtcVqSOLakij2omBAw2qEb0l+alxBwrJA3
kpmuvtbrh5d3i83WFQZskNYm/cyf74qiX+kS9LlZ9Ehd++vp6YFgeg+NENnz
zgY/E2+7QFirfwKnhLzBORi/2xOp/2RKd7by8/9nfFdTnHCruXqL2Qilb9nX
oLNLw+jnPzgBkXWbzfeYAAU7pRsHGV1sIFi3iGBlld7lZobhHPJaJdi1BFTt
ydUa3bfqS6iF2Zd+WCScYATPxBrlOPBpy42FUC2uIEm4IPCxPtzbHoohEc0m
ZjG7Vyfgn4IFFc7DPEeFQP7NZScuE/Uf1znDEJxOX5/0epHxUCi0D0So/HlR
sreMSY/mz7QchKQng7HfdxMlLH6CCYVYJxHOft2EYgG3C0OpAGCYtvTWXMM6
JHP2cf9cl5/EEgTwxAqhkl4m/YI7yu41lKTsUyY9gv5jqVxpXi8fRdHPg8Tz
INCTjcxPUt0O5zaWtpIR9kBzdI5EQG4Lt43KXF/gyWoP7THM3LfElUqQ4Y8y
tdjlljUSO/bYvtrdLr6xl1xLotR6yyw7VK4F4w5mn7Fm8L/bQrzGzKTyrAeG
0Fd0H9UE6CGYCYndjJcdDVKXDRFRUdbPZqvRFyce0BcPYpHHIAa7ZHmO5l2b
OTX63MiCGbUDz8cqrpoobpk/fwTgW6o1I0xEA1nYPCmMuuDM1OTwjxrbCMSE
zwAK9H8UrJEyBymFyGd4fnjgQWBtQp2qu6W4TiJ9viqZOJW/GYPchQd4KMR4
Sz5B6We0dcQkabReuubMIvNZ8SBprn8BCVdmfe+F2BOEsErNNhpUkkZW1HzO
Gz8NmTVRVY0nRTChVJVVCxXK1TRUqDyDHbgUGB5DKNykdpGtxLiN46KUhrv/
B++bryA3kBg9JOCl1qllBpBQEEwFB875sdtPkKNtUeCDCNC6m0TNBV6dcYMk
vEQw+4+5i4pvYaSRFOkKhTYf2uEYJ2YKFLOTzNAjCFwPmu51dmYuc8dr+sag
qNzsFzlm+1kRYHjkgmPcdQEn36nA4s4r4J8ayHGBbdAG6k1jo3g2z+c+rpxX
IlPpyQYYKDAL/YsDdOfeqy5OfRwJk+qC3YVPaYf8OvubPUPhotl5Y+GeriZv
Gm/IO3BwD7X8aDS3HQWRaak+uG7rQWpVd3u0/SGWToQu/N4kWLfy/JN4dKA4
Yof6gnLZ8W19sw4oVZPMLfEzCNW7KWu2mQjbTvZVg4Xoj9CTg4oI6Vskb27e
wpCsqvW2wewg2BDt5B75wGMYgywjZISa+y3gAYjD2w5HwEhtOsjrMtwDOx7A
BqQUT4psLFgT5DA00lMS+zwBt+DNvgdHga2Icgwic3rYJ3u7pfn1cz+33Sy6
6DUwu1wPRj5qmP5NR8Sy66rHJY3qQKX+CldEMa7D/McTcSp9KUAFmYr0Q5Mt
Vdhm6Dm0yzzkNMNmlSSGucjMEstm59vxeKibuK70bfxSxPye0t1v8wovDRDL
od60qNir3/JW81g4XhmtWLUBLox4NGz07ho82GYCG328Vq78UsYZ952vwCVK
hHOo+kY946vtX0y5O3ub2929u74cmvr5DZsQn6i+dfJAeD7/8+LBDR2EFyro
fNXduTSdE0xSuuFOIjZILsMwzD5g6/Cxvs+o+oVqORVvLPFY7ryeG6wE/o0k
ueO7IgHTvwmowZ5M+KLhHk0Rck1zFKlR8nPpBfxqliyZ77YbghxLWcxGx66C
sIbOujI4KQMz1IQLLjQbdNjP4KLHwFQ0sSTcAn3NQf4F8PL1T/pRJ8bI4jfw
nn+muaTW8SnhkWv0nCsIaq2HCraOLFV50jng5LlWGF53w+tLujDNW4OzKTEp
dXk7mO786xr7DLaYr56R+76+Qndr4a/j3WnyJzwELRew4pes7w5lEkBOQ8br
PD7lfK96fCAYuH9digHo5VO2QU5CjDXZT++CLoqg9QlW2KcfJg/iQsRKUrEv
eiz7mGnFO90NPjwK4rnq+6Q30X3YDWrKYKl9XFsLDkLxnJhr4wNYUvZ9Y6kG
xKSv6ZtV8Yck4vcxiKUVQEFpKsVRmo/TG+fHhGjj4snEgdbQSTl9HsrPHUSI
AoK/WAtk+2wJjYO17LSrW47Ey1jYSGxWkTFscd7bOxym38XbHpAQL7WZ8b09
QbVT9pERIwhHGTjVtwQPhCrOm4DNIflznwWwrPzve/qsfoVTU25JqDzhbtwj
xgKrfw81ojy/ITMeXAlA9hWDbL8qpKNxjoKMWRT4BtpKA6alTazdA9Ql4M4w
4mbjuSO5m6O1bhmWpZZPWu+crqb1iUeUR6FXmwEsXkiGDBYjKD1B32GcKA9c
eAvaqglQmWV8qxvXgddX5PlJRB96fE4NmYbezyD9fBUcjqJ9gE9tpk7Q+HAy
vE7bNQkTWKtjzoduz5uMnqYN8HgE+ZcYKyS+h4IGqGFcUhDFAV5saJf88t4B
vjX3TJ/w3sdehPCehHkdE+6XvdHF3Vugsc1zxX852Cw5CgMFJsytr63r6F6A
h9++Kq6YHTpIiWRXzYCiKv7QEO3tiZm5/8OGGiIt/VcC8Cx4TJq6AP3Yj6XE
GqqrR2L9hYwdPwuV1pZtCO2vUco9zszGjhJCKLoB6BuSL0KdGJgcPX/5tKK+
DrI0ns5mMnN3hE3qkppp3AW1CqII5RZ7r+ThbilDSj6eSkgIr9NFXIKIwJlY
1RmQxspYwC74VKdlZqrTbiIYKFqvFDFDPTlwk35cIsEi71ke2tfWtVWI/fFD
1Q0hCY6vTa8jD+29Ki2aHA6b4a34Q46qOrrS2pFR7ijsrkWUBmKK/0vRoWlP
Ji6IAqMit/hsGfK+0otW4/PvBXcZZuQPPE7vxxM7FGL3EBUoPfEQTetnDiVm
Hd4uB4vO/0mqL7hP3gC2QGtPf0XJK7G3/Licq1WM6Oex5XAml7w6js/ZNi2y
Lw8n9JhztTy4BQGval8jHZWJYPnupExVg3YoQ2GkpZ5LTrfyIIpBxLP6QXxq
NV5C6lXS3dP5W7ZItxFEhlLCPSYp35Fo5WIfzAc2SJb1/3NV/GQtqI6V5qvk
QEWT0pnmA6a5wQSa2NVeVESrn+n/kkqtArAXQdqyUwWkHRWRIAog7O5DRxgs
YERXXbsUHCxzeZb/nSVM/EzZD/pBgp3DjCbohWdbhHcZnI5dB4QfcufIV7gI
yOS93g+Rmo1/bGJ2xBDLiQpTflBXensJ8HNushnHL9xbmq1yJ4wvDGBtRimx
H6nh/9mU4gKTWTpOHBZ4P8Y25oNeHccFNjT5/gCNtkV8V+1Jyjcw4uJgpiYs
FxqjgTR6OrQgwjGI2XI5nt5YZ4ZWOxlbJmAzerozbpYB9M+dxSD6kMID1rWx
ji/p330twQZynq78cQlBeXl7CD7Jo/xgoE5Pq4DgXOO114Sz+Q3dLGgpxZqS
r/vJypwsWmzrkAvKy+QRx+KbtMjnqGDT7M80J2JzWszJJq8rxOj1aMuw3W2s
lLuaOsehmext9olXn668BLetOtmGgmbRUV3XBwOZs4FEuJFEzWaiyWjnfA0G
2C7XQJy2rUYYwsw8D6zDIH3afskFdmi20pM2BiV3r8EWHC+OzfXviDTmZLhp
dJszUDUMZN5PZprbzWGX4hgI8GRmvpGRlxB5TDzYz/suG4uaTZwowKi5bXtU
8PFYs8YCRqbn4KWQ7l5xrmSvlS92GPHG2PDQoTvLp9UujmHhUqLN8gkPogKE
BId7Ho4nzVu1UTq12PJKXeLaHhcOys8GBz6T0Ewa3NjFeiA/P79mMzvY2OzG
p2QxR2J9q3oX683ycIHb96+JBs88xz0R8P5Cg9+a8wXfGaX/irSvmn51XoyQ
wHqQW6XzQs6bkBPzn5huKLkfDmch3d6tDlZTfshReItELfQOFQDj7ZWvp4EA
jlybGjjFn05HZjPcMakfecOgyqk4DpAnpSG4PhI4JHp6MNSzPeGz8hc4uqil
WE9a6+nIFrXuHe6CqGmxzMzRnZTYgDCkm5kUpe44vN68NCXeY20gCukm6hMK
01nU4YgskAQLS3Ze6dT6ssrITtOGT+P56rPG6EyjY/zwybQ3N8H/Md2HhEm7
39JV+D4Yd66VWoZH2SmF4NTgLz4dUl6i3kMUMjXFCbIKoS0jYAiuKxcurg4b
DyQfxPBjJXkd4pFk3UbFTvKLUqN6eee/urLwhp4FMDKbGaBws2lsNE1ffm4c
puKiEMe4Qg32aou+G4sZKyXhPog5SE+cmUoJqzVRITJgtJsAaEoNa2BINQak
JeLmGx4/TWSZ/5fiJdIBbizEBFtjXHqNQMqxZrrrOXMZ0w6YyGP9Z8B3RGto
VG6kFB9iDcLpOupJuAFh2z59mHJkG0c+z7Vwxlm39K0YfEWN3x0uM/9xUSoQ
bg/5imXX9nB4mtIhVp2CV4Pmt9tEwPPnfQyWB7x/9GrSEds+6IVllwSRAFGG
3sKbjpNasAlqdytnNV7KxpDUhGnrBbsirS7xBbd+BaG/hgJscSkXlz020PAt
oGalAM2spZKgyacMYPqG0YgBk9QfkwD5tfFallH3lVdZfOLA+czu/YQbDSS7
9uEA+CgxkDsYxKrAe2it+Ngri2QjNA8jGIwsqhjJAg4XdkY2S7hLUuC+H79a
cY69ILTeopiifQiVbtn2aIHs+QSTIaVEZ+WUoy41Ct4V78K2T8d568HY5k/T
1W/FDoJ7EYVdvlBvYqJSiws5pstleiAVMPTA+D22Dwvea1kBuXgIpMT5Tjp7
kHMSn1MgK4iiuT4+ldqyVEZyHH7JtJFIQ8BywG4LlQaJCLRoK3hkHLN7kYIS
OZashmlr+w6wJDA36M5b47oA+QyStFpVfhbv7zwYOMcJJ/HoV7bnt1N8Nq2t
R4ttbdV3ua5Ti/omrF7b3qN9owQxekrbWbwyH3lkaalVZEUO4SCF8Xn8XZXk
tvWoUcchfshzTtAZRfKQPkaIynrxDoGdE3fx11b7Mz1wteM3f3fTTSg82v7y
W15Kgr6IhOFIfwe7w0Qz2rGPv13EyqJbYn13q7PpQWyxwgP/wSoz7zLx8xae
heYXRCBTUGy6vYVquWkNT+VjueKQQYJPeuDt0ODF3nqSvW4QlBzTx8IfWLAG
1olWVN1Nq1XvHiSDhS1fKuJ6XSDp374mS80AKDx6xwOkHnTOtLqirPWil225
cAvcfiNVI1HRA9ZhgAkvj3nGwvyVedsNRGGpsxDdQ8lDMBQWb0aHUbnPLjZW
AEon1n4hdeHpKtM1ko4xU9tDP3O7pIK+/q2C7gXxGHk5xCO2nnAmyhhCbatF
x7N1JEJbhANxTfhl1e1ZAfv/nhomhFkl991NLz/ml6FYsqaygH671R8KBX8e
byVfNXnjxFwGceebFVZ1/EKE6mJFBBNf00BzvCrYU3jtDLGouU2/uvVcBHaE
cUNZpvqCkbRohgjtGJqbsNVLlLesCWo1od8QFomCG7g0rs5SXm0Ex0iu/XhL
73TrZSeJfugA8vwsq2AF+fzsdP4n4OH7R4HvWKgwBDLo97cqDCWZ/qJob/Y4
+un6G1v5AN6ivWnQVlIR2WD/HcB0zrBO7UlHz3TjQEuVACDO5f2we2+XhHGy
mjBRGBM2eZG+/gC43eX1MgPg88m/SVXFJlccD4n/NsMjzMEkt4lI/WwYYEUm
dS/dGpC3pee2j647ABZswjmCC6R7B85yCA1JlU9UPuB4otiiAMdD5d9L+mXC
qtB4H5Ni7akDwe1QAfklGGDHrYrZP0SIZT035PCPoDCBMfDH40FvxhSEHP1n
itpwFziKL6yRdzl3ij6m57U9EXmv60QFP6MNC2U7d+JLVnlZBFFtpajFWVlB
jdpg/+B/2bLmtvluKSg3vUnJcGbF5rw5NxBR0ukBYb21WzMGGpwfscRuTQoL
cEKSSJgnP8nP35JD6wMnxGs3Tt8bJ6EaL3HWeGnfUs8+0wh+W5ow2Mf8PIeA
V/qdouqh0PZ8Q7ZfJIO7gDMB+uFUiEEMA+wAmsPaqV6PplccD7iUQYNkEvEb
IGrIvoRmOVg+OLv7wyGW2OqzCm6kj0wU5tZLz5g/o+Urx/BIZG+4KErnbC4a
9zN8P15LRr/1w/+VIRkf0A+H4Fi/msTeoht/rYG8s9prZ2j17LcMqYk31adV
9VGQZH3+Db3v5BOyjPcviupMoS//O6nCuxuTRaLSf7TrcjHdF1dmfV2uGZuJ
flFqvDA7NW2tVgrjOKZb0/JNbvjtyFPiAdaRfJmyZ6oQfRsuX/viYsJGk1Ll
lr1PZ0nlGxituhBStXb6UJslYmk05plV8o42nqee3PEbsbyMy+G/n/o0YTVK
ThP57Ca3KeWFQvuNStaSXJiSww8VW1LYIQ+St2xw/sm6b3qC1l8X0t62aOja
RaAJVuuHk/bEg8ere/8NSHJE/1mNADZ4KigjlxNZtlyiDJ721tfywKHRvWtS
3i3rQDEz7e48Rw42b+Tjotev41jgxJ7wC4tT0Z81RekYRIZAy9BisPZ0q7i8
v/9UYwR/HbNhu6y6JUBuKCCfUeEsLM9m1eoNaGqzTS6prVuqZRqupp3KhaOS
J0fwBEwBqjrKu9bnd7dlddmlXuTCOMmILSPh9Up9I+S59AOO+ny3t3rCAEJv
JF7PuH0IqrisDAhQRW7pcOHGVLEaudOkY8Ln1ZKtCP4TLXt+Jl1rfqxEQ4Iz
ZgxSxXJDWpYvGpraV6EHSeNdfLYqkyT3CzXNt5/SHab0FrcPJqkTUxR7nbv0
3aUkh43VRyCg4o7UiAKWJDN58+1LWBfrFKNqI1FSo6oM9YxMhT+HOLY2gkPu
LJ7KbRXZ/tLByYMsgHbOky25xZJf8Zv20jM4HC3fMFHtB2OT0vH8BdQqbP3J
YKrx9iZJp8SyriBLJsAm39TlFR3vJPgqda1cmzZoDeybjzsYRxUU9lU+/N2E
wTCWExLWnhPo2GCBG19B1esjRAtqCVn9+Rz5X8Zxxo5oIGFLAbfhoTEofZ3u
cR6AOmuYjIOthG03hemfB16J6UCVEXIf5S6Fo0q70llJhIulCzm1Qosv34Fd
f8IB6fef6CvW9VELZfX65Ex+7AdiAwxC4ZN+LxiNAKGgA7g/7BPHBZxedzpt
pPMtgerO6BOOJJYB1yJKt5Wdy3BlzOboQdjkSHUh0elh/fHENn4oGdBYM16f
WAnnw+PBQdjox3h789iBtyxoSjQvfCzj3c8NrfAeC77rrE04Tgt7GIlqUKI2
oGsn0kvfpNSpr4hPUosLd6FQ/AzE2o42d0Z7A33XHUYdhRz0PeYB8fwA42UG
hru0z5D+aHLgi8YpT1euaMlDrhQwu0DSyoCIUP1Dzz0ZSVf2qXCUPHv41QoQ
NnHYV78h2g2orErwkHANEzV9bdkGHNCn3H/hNbdYcCeGd8VxO19wORLQ3B6d
TRQQNelX919pHp8tHdheZgL45TKZoep08pR/XGsu8smSaGIGEMiTAuXKNq0c
L2/g5GHmHiBKb8ZK7H4EI5kvJXEj2N9TZKaSkgNL+aY6d9eVMlwVsI7GdDgm
oZJ08Xpq50CFP3mMnFouIjtGSGtazQyWkSulYX5V5c6kVK1rrbaCkAQXhny6
9q8SnswI0fqyPEVZETNNrJIrWC2zqc618ZfTpRH1PxntqjfGjkvvgPzCBz2s
UO8JUKEGf+nIsVZukbRs0Wm13nKiS8SMELuIzGjG4/6nVDp/ZG8mtlsM4slS
RMUCjAJmD+D02wbPufwDPKOK6oonbC1cAC6Z/Dyy5XGL+KrXPTz+xxwYL3kG
xzcRH+Znq2bOTRpf1EpIJo1HWKFlh9Wwh6hzVN12jTJ9mI/zgBl2Oo8obsli
r0aU/fHywTLr3Y3SfKJmNhrfAbxarWZgZceuS+Qw18hcW0NJY8UcnomlFFks
QQgLuKOm9cIqPsa5Lh2nFUjzI1TUfF25V+i0oza5wkkUIq5oF/fRDjgOr1yE
bOGAzFwizuLlwcV/jEY+9/Ko/TWKxbasn/8ZoDg8s27b50sv3+1RFXzmXtAp
bfMk0hrB9oNt1GPTkbr5rs5dSNtK0QnoqFaQ5eHA5Ma+ERCFYWTwVPixO/PH
qvVvZOV/2amplZZC5Nofo0FSY6UWSZDuexrIPa0oGiwtDcP80XcmYfnJWkdS
pvP6jW2SZKMlPJ6tshyOEHD3/ooTLyoNQIAKsk5Is7t6X6cilLmWCYSqedb/
JINa/P/SrrHo4ikq1o/8lUJcPJ2Jecjtu7l1saoB+zU6IPI9srpGjiVNVG51
SHdkarskEQzJJp+AiWrgghNrYNfZTbxpheMIQf7JJFQionE3aDPG7GBjTN5+
CcyqbGtxsRRF+V6w6dpnJEV46F5skCS6s2Ned9pnI1rArgEtXCnu6LZZqHp9
QxI1sgKAAi0aj4mUQQHUTCNfTF+ObAjyHFzVbmm2UTK6ZvFXKXHpQP5pFOPT
mkzJRJ2eQcagbtN9hMnt8UWO1jhk9GTSwW0qbdhjNqJ4OLRoX+KcOE61RNh/
xvECusLUlFfIkYAQXkb+Dc6K9MJ6ut5HFlt8YWYuSfejRpVsYoNKOFU2NYPp
uNyyhObAZzzncAb1BVvyh7kU5suM2HyX8g2i+Xnqt+mvVyHro9YaK0PpNcJC
xecv8SvNO8grpwyqBl2euACRE9tc5Ea3bisrCTX7YCrPqC3P2TA0MSgYA4ma
oJFHrQiAjFGjzSqNhHJ7l/ZwfA2YEKtSYuhH4ME8oNg0CUQUn7Qr53z2LF2/
fTR9ZaE0CEDMcPjJAwnAC/MXDbYouY71W89gEDFqJcAWM/a11+rsJYStKXyM
za0mGGpLF7E1sIf+33sT0f38M6276tOEM1uoiQsKkFdXmirKVPQT7B9EccKw
Yfx3heYm5aAy2kfXtfh70PP0+uve+L7oWcfgXUFnGII7jNaaNjF674I1m1v2
6F1Rhhy1Xrp6bFqsuStUEDDxvMDy3eGB1GMEJNn/9HBxOsTVLVqs3nILjvV/
xNiwfIuAs766OuSK5GDlainPiY06r0FgfDg22J2MrFTH8sZ4Q4eT5JmPtJbK
oJhJGpPFbj/VUvsVw+UxcG1BCaJCKmo4dDHtStvicv23d4QSIE8S3/yoyQip
vVLf7ZmEsD8phknRk/CiXIR2IzzPaKPHa08aqbEY8c0PKGowobsFf+pRglB8
v2jqZ2tOFwsHRf3OfmF8EM5okg8Z2+q/AfruJpBfhYsu7K1ysr3pBUl30y84
JePqXCKSoaKsl8DC6DsEa27pZLxvFS39ayRUJWleREu1eQtu0TVJQGJoynqG
7vj6C+BrzUYvGs1MhQr11XZ7F2PIQOQ5A9Cn0/baJ5HK0sx8sgUrYP3fIHAO
iEBomIkty+90XQn5pbUANmPXyLPkkYhTbY45K+aCqaa+U+9AS0nOXwrG1fBV
d6dvK4H9GbA81aIwhbft4t5LrRIPfJK8PYn8wTEyELPNbzgAjrXcLGaMfgQR
kaW5q1XBPiyxRY34qshb1Wq47zBGqPovoTb4kEEAbLsAmUso1fT/esoBBIJr
BKIiVlPbDRFatmchWvlSQbQtcBFCaEBzd4eb0wg4rG3gpkrdgjE8ZXL9Esjf
sSvohCfMw/71MFafwQtj11lIcszpp2WiKhVbW4YWQU/fgWyj0NSymnM1DOFT
bcfjNHWYXRGcVHC7Y5cEfbI7DPMQdgIGhxSRALctKIsie1tbLbmeIR5zb1OK
l4g9sB1WRKwHYCAsDcd+OLDYkiChW6omaqSub2IE1hQDZI0f/Nibdf60zBHh
jH2sMaE0wnoARZXBZiTnz8yBzNLLMXKltZbcIXcTlTjUzPTi0aElVwmcm20p
X/JlUBP3unii9Ktu4MBjVfunxQEoIJGLdaqjCgOdzH7XTFvnXWYBPAxTNGoQ
0JlDpismUjRTtIaqqvxBauwscAazKy1ORWsp1D/T04o9gmAGL/7mdWUiBPAZ
X7EehMRZKMWXj2U21yAN3IJ/jvKOz6Y3J0elOveBE/wsmPNXbRcpZpLDqHes
Vt3PKIRXOA92depQA9kPUWu38sWc3+CO61mFYCRuVjngqfe07sHbwKeftd5S
Qfgi4MnYD9LYjj63EeBeeHzPRz8eBIz+jmvwYzkUg6++UslI2ckUAdiB8r23
03/nUx10MOWTCGGi13gZ9hyPLUiOENhGndZaJD1OFeYjW1b1BOvJ7F01xOHN
Mq8WWiJQqDyfT4NN0CnFPbdKENLN1agfdUFIjVrF/5jlEfU17HGz/N/JmPG4
fPAZkUQD4QoA1A5peJOXBcYgxyeUSO0b7EIvwvOwVcb0/KrL8oeZg2ovrExt
Uuomt8v1rJlvk55eW0fcXuRPIgYwyUPvkfxrhoqwcwHQeHiOhg48+YDUXmyF
2JgP8JV9QaDtSTo/PT2ySszgnPe94rV14XZNNAuwmSwCBOg1ibody9lmnuJh
zN5ZtLRpNYTC5i3bC5cNDj3FjOxeOD2dUOipattEx+zr5944lNNCTFZ3poQc
3Ge2Qhe69J0mLdLgbz+vdWHHpNQwdLHcg3pjv3DfvT22TAUcmyPLWsL1Wo0V
AR3JIDVovSS67hLl9uPbY3E4+lWLLcN9m0w13X4fBWSfmTSDKDNnQmg88nD/
71uDr3qg61JgTkS0EairBDQLaaCH8EZWgohz+LKjSsiFG2OSi1qu5EiigOam
Ef6vzAXFWMhx5+iZ8XbBcCafyk6Crk6NA+y/9AGFN3BRUvkCWSHMJ8MQDOUF
q/5t7+xKb9RBAL7rDHmsqzFMaXXfJgi9yC2OVTpUdoyZ59QNIgpqfbiDGd/I
lHZbPFSINEU16LV03DEsT4EEqHvo2ByAbZLVtrMT+GX6herccKPO2i8rglbT
uhxSvVsUSfAkUtSRCceswwwjB1XrO3cgCcPPWtsQyHpNpCz5SH2pv2FmdeY2
gZSvgtK7qntUNF/MmfMx0iKK/XCNedktHndVYj35lUyIBt44tC/jn0l+SRWP
i4AyCl/70oTVhENRrrV2rqIeC9lRgPxZJQKYSH/rHYcMMdMfJ7C5WAmhHloB
4M00vxQaehBIckcb0ssY7cS2YANZttnwtnJkmfZT4RZZKuW8VnMJo4Tt6AhN
40dW26CXL9ZbdOWkdmjDwAwMZ4ENfrMvHwAOljReMuwOei0SahjUpeHOfcQE
sImSRVIkETDwHFJ++v8NOVf9PzL3ZwdlaKXkji/9Gw/gBbt+jtGnDrTmnZWu
DmNjYm+nuSV7zx484AfGnHHht1myvwvcGE5gCn4S0GFgVPlM4Suf4uNrJpPM
IYuDC6SntSkHFXbEcUWaWlFZuC9+P7fO6q/3Pk9JgLOxT7MwjeB3VPQ3lIML
45NGMFTEDhnL9AsZJy5eFfCbTscFJukCnazymoWtj55GPDjNNXwdcmKz8bVC
mCMPQTuXRaKCyS+6LuKMfPDej7K6LmezmGCEVQG7o3ch82RATDJ1oT8iFWov
18Ct3vdlsrZRZezvnuE2sDM/sWxR8Y49zl9ya4uRWm486neTWmGcwqf1G9Nr
CqK2aR9Tj6R+yVuhQHlFD4aGs0eDLu3LKI/6zyC1uyYQQAc/CXTz8QuaXKGg
K5iGqLrMA+iqELK+GHpJs0nZRF3AOhLPToJA1kQv6+0ejvBy02oVtvHff5Ky
gSwzOhQtU507lMEIO2G8Rtggpn1wYGdFRLMu1NDShynqZ757TnwnJbufP30T
HBmw6jj2UsUnTKDekn02B/Ogj3nnRDoeU9clyg/n4r6TBIRXLcHcJjX3F1Q/
D7fLEjnXBJMRXdcFZh9Px0moLkFa1XlFZNrs/NPqRKi5OQk2s/eoAW6TNX7Q
QKfnMs40qfcTloENQYiwBMMxyt96T7rEEiSctv2Mgdkev5rREfpe23TmAnOh
gdVjP6QxnL/gYCvchUY0WlBcvgnqQ4G9xzrG/uInOn5FVcDRTpICbMkAbkyB
F0hZFgpCBRdAVy+mT+zanUh/22VGFczf5Wlxw7i4+/0bzRds0aT1ksDswmgF
52E90pAEWc0ToondfEUrdwsz12cg3JOVcS1XORYqjr1d/ogtda1n6T7AcXem
Hal0IY2pIdAJtQqLz/p1tuL9/EDpHyzeb9GK7q3DEH/lgNvo+eLIjT5fl3TR
v+rhL+m41J4i13xmYlLrV6dXfrhxwEkFY7lhclCAa+bXIHVoHXLpSNkaD5o8
DyvjtPtEPNOo4mY8qxlMbhNrTIk+o6tZHwAxM3D3e3Aqm7dTo3JwiAAzWTqM
PA5Na/jm8c9mn2HGNpb9f/0vfiKESyiLFqvfYIOOIAxLDMDKVuIPwAcCLoAO
JuhYdLQUqQiZhT6lA0Ba6RBpYfvG7BFfQ9iCPEr9001qtuRrkaeL6O0L1o68
RO+ugocjfZp3ZZvd1aY3g7TlviaWgRxzcF6mXMC+nJ+xdUuc68zaZRPNiS/q
+t3PuhtCDOrRqYtSOfcUIJARRwiRweYwzq65x0H1wzSDQkXoK+3cUVk8f4m5
3PGwtaJly1HeGV9ghx9MjiwpMhcPGVZ5Ujds509QZdOmgVNO/zoRKNqw68+J
U5gfqTdkviNqdlSGGKswvUlftAt66rYqrBUExkTmUq1LdXQ5xy+OOFR7xmUE
QxlFoUfRCLAPUotCKms/YgE8/Hec6EStxcgf7mJPSBr/wAbJ7WUJyDr5Gwyb
ohGRiugZwES6JbQH8oW3hMpGlnSi4klj9BCdTzNws/96VxYseJd1awsdEtmv
uVAESyPKlVpFdf2tLU4lSuEIr8b8vL2tmln5SqLcsd+JFogaDtdlKKTQH0IU
AkqITAhGtb1JTnN8CtpVH8B5s94Z+RcJXUPT2KWiwjlIzXGfXJ4g0E9Hz4yg
/Dl19vWefTmlf50TK06mDp9AdiCmdXkAqay10GuNxi8Y1wUz0bJWqjacu+yU
SFXqPKa6O8y8THnN6btYg0wbnrWwk1t0UBo32XsyF9ZW2Y+WLHjw3dZEY/mk
vbwtxF9F6uIcDfUDUmbLmEFlyuvTGvLFIZU8wOtU1abqM1Eif3d2GPL9Ehiu
EKGhXB6+qLY76nXKXPJDefB73ehFUlgphtd4TV+sBiIk+0/IdrcFGeKkYxPz
D7xlUP/hn0uBzTNkeEpyQuMQu2Rw0Pe0+7QvZyh/no7LJwzvwaThidnj6pSR
pL1QxIaxMUjbwiS2p1e/XMtu5cjWq8h6dmh1KHLlAtTJYm1Zf/wph0A06fxT
DDQYgcdiqczYAGQ6X2XpC67PxjUzrg3KHQYpezC4CJ3ciypko+sCw4fEPQwp
llixh9BbFpGLs078yeTVY697LtxVaptH74vp46yZVwP2i+HGq/Q8ZlXzmV4B
nBKj5GYxF+bTplQd9dlVasYyGOgy8E98w/6AfV+wilJGJz1vjMLei0B2rjxP
sMf8tNzyhYNDRxwTEIESd/hwprmqpFiVhFS2PbkDVxH96VxzuHqQnyxdaMOj
YgqO96l8qDP+dZ8jya5WReKnYx4sRiE+/u0IsusuA2U+G3Ev2zw+m/gNtVn6
T7CAfxYJP+kVGHiOCaX0ZoHtNYUTJ6B332M5BVaMK638G9Tz9F2Fhr/SLL79
wUG9sYTVDZp0awjdqd8GosCs9K9PqYnZ0Y1njJaZgawiSWeJH4K+kr3dFGvc
hUezvMmTR+aK9kiDyinwyksGqqhLV4p/ykVPcBtytac3k08/4yW1I/6E7SyV
PEGZn9VxxChQBLBippdlu+WoWzKjefT1Dg8kNJXGFvnZ/sJwOoijvyurGHNi
xOmRI4XxVBq/aryiGdybjsT4OI3LipKpfQ++uHT2dj1ST0mDouy4rCeSlFvB
wdMvbCx20zD2Z1NtbLiOEJJoyG30L+pbwbpFU4a6crbLnIRicyM9GVwMKVKp
GTe3WvwpO32ef3jK6YiPyepxNAjYvLTNkVfyexv3iAwojbh+VDNdPSe3vvOF
DJceWNv/KG+wHra5XbajIiDIinfggrUqnky+AASyzWGQUQSKjtutWu6fLlkv
pYs1JYyiiyax9Czno/PA1W8qD5QmvblFg1fmLkS9HIoO4Aq1On4s25qyOXRG
GWK5l4D5i+sSev1M+WrZ/ARsioA0j77ypLCAREJe+JMmE/dglzmraQHET/Tj
37V6G35YbzS3DXAR85ag6l/O0ylUxeugLae6rTpWmbrG/YD7uyVE+gPuI31I
f5jqNtVn0anf6A6F9Xg120ibr74XYiQUZUrHazF0CVhe5CtNhuJ0U682ZEux
7t6c6KddYcWZ4kLMxtSnWx0n6rh/jV9weP5oUqQqKWC4JfAmnbAciZMaPqMP
TPpVb/5cuowJHRb9lFgfsdtBJIImsqtGf6hFE2aviBWbZ/oMtHyJ3NeED4KH
wqge11Vetr27xadQvOCuXx2mL0iewcNrSixFgxiCcSYzFc+bIYclFrufFG0n
HOCaduu27scaCNYPQHg8CXSIFMl8A1iosYIG9AF6KKLC95eJ3SfKaqmQ4TIv
yyXebYyfHdNuUWSNJ7/C2mLoF7hxUDdtrup0uEsp36NJselh0l8hipkiHqIe
y35m4xgpfCCCxSWaGBCIqGuHYvmGu/cDhALuCVyn8W+AMprFJzE8j+sTGxUY
/B6xXLm1rvxVgV4tbHaHq3ItLGwKe/lI5sINroTNI4GixEuXRCQB1H1d8YJ7
lCffPgnwZISPPk5742OqWxueeaWU3fPo29z7ld9Pf7QBev6qzB69XLhoS3XZ
NCW9tnt5Hs2XhFJVIP1rXXxy/oWU1qhL30n5x5SwaLf7wFAKHGpHgxF4aIei
c3jQ+kdW+7UXcl0qwmv7pQbqfiPD2QVzcMiXcuA/a4mWaIDLEnBA30+pP1yf
a2L4YIm0DyFIQKmq6+getMqPvwHM+RXrYHjntSnY9CKfAKCnU1aKidghYI2H
GgRQQJztXuS2W1056+GCeYcX/hA6dnvbnOjSjINpTt9HBeGM0NjFWJ3kY8S9
ntG0lZzcNOThgZf0QBD6NSDYN4JOvRUWIvMOQmoLj6cF0+FaIhqvMopnckfR
XGK+vupGKXUt6kDz9dww7QC77+XKRsWoyBUZNHrHPYJvdofeRACvSwi/8V9Q
KINTGbWN30EqLz7f0iO9fSbanUvp6hIW00oSDAXpye1e92pUt+O7OlM50ft9
2WGkGdPzWMHYzOqhMZ5bGR8J2HXb26teXq/NoCDSzK/LpKHrtjEDDkn2qP+2
4MFUoh3uWXX994DRG9AInKjPwTVT4JdiFCJSiqrK972BwP/B7+K8OpDgUxoz
rj+cbkq48YBMUWascHFxr/v8bl96MCMDa6ZZO5US2ZEu0HoBhRL3zHrtbAAZ
2RGnyma9ephmfSBk5uCijC8t4MPdeKtnEqCycyEJS3P5n+5mGCjFMxBI2Lzs
53iyD01FVPv+RDNTSxJQTVMUvAi9MWN2h1af2d8yscXmWaWijqvBk76weth0
bOw4FiSnVAYzEGlyf4yK1i5JS4Z7ROWcpGwjVylnnIxnSuTjfSOjWJQJHKCQ
WWjICEov9LsPeFdzDUXW2Dzv7thCCw51hpuB9d0OoUlLv9qtbZgnmktr4vdG
m4gsIXM8nZHV3g0ir/6sY/xiO09IuAztapW2OVeExjSFTb9s7VcH4tH2Z2s+
1DGdn9gNw8Tmnboxe1V+hyI7tPt704stsR/RTcL5hN5IV9cUtXf5RJy+1qhS
dwWXFW5e/04g2cHMVUmEi5MtbsqnHVIA+wZdTax1EhIOu1luqrhgJEumwq4W
fit/CwnIlSLCobuRWBBb74Vh8/yzoqSWrYsPyzDgDe/Xp0UOaH2A6c07woQH
jD7E2ujhGE6Y+2KBzJi8MD1IvaLJgdknTX3fslOG/+vqz2x5BEpjjOV+ewj5
qPFcQzY4Q28fc+VEybMZTsjyaHlkbDWPDtUJdZPjKkDuGjTUDNVSZI3X3DFd
8A2h6qzrT7gb9e/Etp6PbAJrgrilkS2mbQ4ljpnRBpLl3MOOc/TLFdE9+leO
pRHeDF0BA17MkSmcqLVu9kfj49/Y1i/FlTJp+ooGAMFZTD6bTZqfHGth4Bqy
dWqr6GLNBX43og5sw+9XvolR9/6BQsWP6wnH0VenW8UZgPxaOCqmZeOrgHAp
VjTApb689pL0n/LDWvbpvzYSfScDRf7ZlomMz94/uqSJbgDyR68YrWLSokDQ
iKeGxUY/0k3c9uHI4PgJszqrkLUPq1QD7xhIgntz/psLGmbvaP3XyAbjE203
nAbwi5UVIyVCn/JPfjdpiMGwo+qocOVZp/Jl4UjKizgQ0MC9M2T9UzUfSxrP
P4P5zvxlve8tlP0IG/di5g1JWABPxRL2gP6POjUgBu/ae7pIwE8mveJ+ofOz
T6iGRtrmtcsVfC6Ya6KzQjXxnS72hY6y22BBUXX+IAm6jkoxzxbHXYQNYKD6
PoBgNeKQoVtCsZSZn4NDN9IqKwFMCue9tHzdtbzCvkbvFsyVZH0aZ70g0UVH
dbL1S+f3wVEtSXFmuSFqRF8BSUoCt6692pSwLobF5xddOWjKwBMwimiw4V8O
a2t+sgCzRCABYQ5xJovJZ+BKbP0ZOxMH9sYxW/Cq3QqTHSQNlPMvdaTumQa8
ig7TDlegWPZmZt1GE3z2Hsj/WfXKHFCvkZ7ZRgxNXp8i97Z1nmeg5IRiNgtg
M3co/m5oNNCO5cx/TQ6guTfs/uqyc7AMqy2Q/jHnRBzz/guxJ2QF4nXaWzNR
a9fQDLtehtXnFqUewX3UkWHZl/YZxbyMWBR5A7Osz327bZAHGGQR4gV8+WxB
YKbxkmMfE5T29Q6wcnrhSOZjsrKy60bk4cSRbcXTmE92AvwP6mPtkHK0mw/8
ZI8RMBYkJnf52AsZMf6DVM3AfY1mEqizv9Pf/NNHxca8UYxP3kwRFmsd9P2K
kJANj2CPRsL6Lscx5WntMoIQRppKCNTYBZU4pajNWGI/AFnQK/mZt4jaBrGk
WAMtZDti+n0xHgvK9EcdFra/4PoDlVVBf8N4qk8ItmRI3XJCJZBr5VaQ1yjq
DCYpJFUK//68NrzxbxWSNcy/s6y4bGl91qt33tUdov5Oh/w9TyKohSdbLccL
N6HskkXcqQPeI2oLEFqKCpu93yawW4JIUVBHy09ZuWhumKrwaEkdL/oroN+Q
dChdDZLYVJuorhl3JMO7WeLa88MQfAwUJ8KI8YXFqaugaRMDnEFs2aeB3ZR/
9FqP4sJSYvZOpvwBuWXNPkblT3rn6qux9/kl/n84Tq7rkfQxJ9nScX1JbdPg
wCOPc61oRF9WNNg/F12Ful5FmaKszaUJHqvJzkMU/k6v71j5WxufCH7ZITO0
yd3EhBOXtb1cfRoSlQRqyDU/UyOwHgQR+HVzRo+m0pybYleo5TGrMEvkLyHJ
w1+oh6IXGUpu+FsUxRN/wcn4V88Fjr7LpNr/0LP1wfrI6RbHEUXwfsmoEyBG
AZVW0nfJrYsGUVFK0s7VTd8Q3iq7NMk8A77DqBJB1l9Kv4qjFJn3Tv0kvwkJ
pwmqZWrX9d30ZHS/hOV/BwQr8s/J5H0e411VALevr5argC5Ad0plXMtB64yr
m/ZAR3s/HgDqxG8ksg/jeMl7gWCXfhpJmbzSsZyOMBqWH8VJ5RqRzUIXaoJI
9iDlrlO2hHehA+oTDNdgw2MPs+s83+L3gbYebljIRggwtjzkY97ICNS86bHp
aXN7jtwCFDnJVPgrHh/lcFFhePCEGCy72LmYZokEeIw8DAxviqfzy6JGLKTB
k7wkAfh6o5y7DmIWSmuB+5v27vNfsVOrEOMovTvAOVUGOJs5h8/QUhyEhwE4
wH7qrAv/S0o/Wu2V0hH1ixSXQgZ+YYo+FCFTaNgZD2ie7DqxpvzG/93EAYva
H0gHZgL7T/BU/bIrFbk9FbjdDHlO5qUqqyYPr8IPqGPenpFX4ldCitP6Gi0o
RBdmwWEqWyHaDbQutsNAw0pafk8CXf4kFRI7f7sWo9Wc57ooKkt2BPLGUXbg
U0kmTxutUroApJKb7Ac6CO+kQ9aceCn7hpDGv3NuUhzTeaxCGNAfsFdU7cLy
hCQbfTrFSL4vfpyrApf7HFbBzkCQxRpm771/pZvlGOWljXaR00wjftozQTH2
JxcMWQMIggVT6jOUwzXsUOGrnQdV6CS2c9FDLoKrf6mZm48XLWy+O1QIskjR
w+dR6LBWVsc0fpxwNl616CeZNNi3NrnU10vKpGtMoRLgC3uXyHZ7/FEzuntF
TmggTD/ZkDIRowrq7CrNRMFdiGCM4FTHtvX3clixlCdQknhNy6O/ol4DiF83
Co861HlSiicRcj0i5IaEDvfQ87IO03v88G14ucPHartEAP15+nnDtQWHRWUZ
mvm+o3s2ppqP/4Y6WXXSaWtA7u1Im/zbw642KcrZGodp798hOFIy+od40P4q
zaCJvAQCwblwAIp3bTJoH5PpY2R+M4dJvehBrks0ncQly+lb2kUUpJAGPpA4
Bg3WptRMVbBq37ei9Thf8qIzFcrNJuD4UV+CTZrz8y6ltPaeSUzH2bVE4pRs
kCVgR7WlCqExSn+LBPrsl1hPKFKHUUY/zwqIsVSXU4vnOgBBv5CCD7ON0Uup
Be/9uLcQMRy6kl6i097P+vqfjFku8aXmgJUBieje+S4sjkz7hbmoUMr+zvLF
issU2nx5QfbpP8UBNJesh1Yb0MXkiZ/bkJmMqxX3171fYmOnGmPibNZQFreI
LFLP/w2HSNSq9Sdx/o0S+BaBln7+nXqbWh5ztktKPxc6WghdMcz1JX3VuRtP
Bd/cdUghlM7sunExX4UOGF+j0j5Th31ykUmpyyzjMeUz9vNgmAkU+0bx7LfR
OeUpw5H7trGhXuiarRZDPsvOeSx82tCuRrNJUgym4jeqaucdnO1vMUcl9Ud2
MuxKGMIBaqJQ+q8+BY21w8aHHM5hfeeXIRpgK3NYOzVlSwWx4rE8Ndb83/h+
SCoYjWcjwbNjckWtCrb5i1DYmbojoOouuzOXerzQYAgUY2265iRvQxDEIAOm
fqIVU93q7r9ZFXybmizV0O/51RFwJ81KWh50yGlcez4U5WF7+aoxZyO0/r7p
uvOvH14BKxtiO8o1j5je1URJMeIcj4VSQks8XWHbgBs5aEIhydPnPAFoRlp5
Wl27X8tx0EaUYg3wjPQZ1C2+jahVIy0ZlvhakVOg04N0J33gfgLq0PrAk2fE
BZvNG4ks64s0LbuqM4s8PHoCbZv8q2ykqgU2ARL0tauq2scP/41s+N2xUssR
zKNwG2NrxyPVpKTr+8yBhBpQPhks37USSaiBAz971cvSSw3sIXKnVDT52RnJ
ygZvzCUULxzNwWFporIZeBK0Ly6N26kHGIF0bW3yX2MKtg16OAT/YOuvBPnT
vkeYT26lYwQgfZw+Nw90twmx0TPRXS56GP7M22NzvBM9Wpe3GNM87Vto9uXA
aKwf3T5gmkMNtYglENhMjuEHV7gSYIQ3JScsAlMhziYmicnTHEzlTXbG6q7N
2ZnjNlhopyuffE5v/DDr7yygeXYHsRWF2N5WzWaT6RalWoDgUcvuXGy8r70T
a+bEpIFXRZXi5LQ/hS3YASQtufhtJD/f+93NTozcJTGJxLup1GjPr9jdQhvG
aw1aJnyISoHwCVMvaoa2/zgrZu/MQkoHc/L20CkgCg00rdK9Plh5fhFzOvtp
/Dk0DCvqIZMc7NafAyyzUlnHQVAB60m0WkeOJv44TCFXKPqucLOGZPZkRstw
p2enYu0bcY3eej6lmez0tOo2QowCwuvkx0Tg1PvC4e+nFPnjsPW1lDN686zd
n41M5UGzd7ItEp9zKY4G1wscdsjCNR4NwLd2sRDOtGICL0ee1xVuhjIL5z/J
zqjh9SRGhPxv6HjOrsscDkdsvtlgJeA9N/Wf+rM6WSpcR8Lszq1yTJ4Yuz40
qClFtnV2TkdU5NOoFwQ+R/euXu0FtuYs7KC0VPnAeVwj1PSwpWDhETWmFJHQ
qt5u3mIeNPhe2kVN/iyP6yuE2enIeFH0u/VmI0bWjTMTDd13ZwyuX4/w2rPC
SGA3gJFAxzqUXBwaW5fxZpbbXP49KhAgvcz9OnrGqZsHZrk8VUzk2TpTlc1w
yvYtKLqjiZGJh3Tewso9t81KFjN5DjhJGMnYYK2xrQ3kIIsPz+T3UrO6/EXB
bfSh1GYxsQYrPfjkPWKVvH0kU45ZpfRMcos5NtmIj3k5WHzwYzG5WvhWgnn+
NYfPUFDKtvcB5k8QrzSuko9OOka8FbRVJe6+ekMwDt+cZTg7s9WXb9f5vQDT
IkCTjN30jlxE68X3mE9CDm72vUnQsqG4iALzaNGg3DmpegbwrY0npGc6Uopb
t4Kr46LNChL6OTfO5GMqAL/ENw3zLRxtTSoOYEvButCskUqbNEaO+vk5/Tue
WwnZQb+y0bhvMcCohou5BzDIfOWdgbfxLG2zwwS3kC22t2FsISP5eI1o/WET
XEJ50TcW+ev/K62SSZZG58aYNUZnFWqAiBG8DCHqsqdk344v3Z1n+47QRfmM
jBAaaJluAdjgcGUA3JQdKeMUzEtPGmeHNp+UjLpyVUfSU692F/8OzPDBRpjO
uwLAAmH5e8jv6jdI28MfL3ko1C6N/bSJX5ZarJcVwoEuqVkkb97WFwbHbpd0
eajM4KDYATIv3d2Zf+5FLEmdwQiP+ALlH1KOIJGhTgFw1ZQFt1hEP6fnKr+x
AZON4cwc9GEQzAPf9BhT+ChooLA2QSPIYSbTmYO5ZhA7I7bGeNI+0SCek8Kx
DAuVTYViiXaaBtCKs9jpMt3nhfyRfju+ea5Fp+kb04zxy70sHEi+QcPo3gjz
dOgv/2ilKXJS9uZ3OY3W+ek89Qpb+Gs6wfhDC5kGNiYqclmKZiCjDTD0xB4N
HxdfM8ExcPT3lFjPOI0jTnf4VtupRT4xEyIaSNyUeZFQo6+10nrl5OwBW5S2
4TDzg6X92TSTYTeFulE8tCJDw6Wu6i9bZq9qZeqt6h4UF0pghT/LmOvYUsuD
4YbyZYq2egzh3gm8wPpXTRvjXHHAd3YnK8GP8rubG0f3Odnx3/DIApAUVVkN
vzoJItW52OMYSD1MobOlcbl0u8tUjfLIm5fl6RYH6dufzKxxn4jJUiVIebRh
obqm7IBPkn6SdYN2GXfE6RkAod4SyAZUB6yY3GIFP8PBbG7zBrNXDydKXt5Z
elU3B5Wkvmi5XCSyMf9nwFAsoGYIUjzlAx21P0Sazuv7eRlUafJ8Q/EIeDl8
CXWhp1SdXIrCgqw1kmY5L0OWmCEYmIw2vVlFXWopubwMvdeGWHCFNWaui4/t
fhtuABRDrtkK3ppMBnxuIPI6SXXfkfv0tqKFXNwmurJ1T8F5Iu5sk/KMhr+n
7/4s0ktLA9/Nfi3zAJmGuUm4hXxOMhXvVQCxOicimKP4rfREz7Wltgek7yCC
FozSa7ZX1OoadsC5NpoCTUg0/a4N6XE2/YMbwnzBAqYa2PNkvi8sPyFAq3Xz
KTS3yn38Cpyr0dzyf3tVzf5+sJwxM/uctejbm3wNZovZrYIcSaxYDgDDrGxX
09HG5QJldMyP95P9zZzrOy0sV363RmVtcHq7pUSQqv3e5pQo8rrJi1u7tz2H
9RpCfUP2Cs8zzIbmBYRawf/y65uP04qB5VSiUsy5EzzYcm5Ru7WxLkPs0Jem
xERinij08W1swO5te+dqej3HdskBK6yJWD4Qvz6d9k/WSv4Oemx0p7p1P5Su
iqS6o8L8vjRx8/4L5pP9Fa4aK5uUNlJei/GCpsKd7xowV2c/LK/PKicgQdnU
6qVDjGw4XNIhmneIoLS+eK4Nm5gaQusJEHitrKJAPIj4s8ouX+vwiHDxSeZA
EnHe2NpuLZm6F9C0kw4vHNW26pUdOSiO2/lsxDvGuv1jyIKTBO3i9HKw9rfE
b7YD8qsMXePpU1FMJSQaYH4KiRpzJbKV7AJrdD6Lgw3bU6+QK+A16LAT4P2O
Eu6eCqtNnx+CAf1vx/6zM3tNmuUfd+ThUjVvs+Iuv+caTv0QXXQ3qukn1UOL
DcCPECAdl/e6pnRDAWZyzBjl2Ozcv1ARfYe92G3o/MS7MHtCOSb/BRJGaz9P
iJtl+fUb/SGNyAbXHd1AcKUPWoWGxXexPPKPSPozan2JkiDyp2WiO0J1V7SC
Xca5G7Vr/WvRM/tZr8SKji/wNCIMNiPtL40QaHvcEXZ56iGoshjymmnsga1K
72tPg03RB9AjijNQb3jIzcFz8At0dOZ0QwOlpB7Jy7IaPZx/mu1WOm2WQIt2
4dm/Ob1aKEtQ4RJrJDqTucY7EZhV2jUv941G0vUChwWSfniC3FzwnI8UgLoM
M3kHIIcHaW8XZZiQ429e36DrEutzSTeuRlSV9fvkj0lVKYwIcM1lt7yNZxIF
JE+VqjmNdBhRTTAuJGjIvC0kaSBlCa2E7+UkkKI7rcGDYQOZllJuSv3db384
QEIqX+oBR+E/KUTW0XlNPQdFKp0JJMOyM+aq+YqEkJzL+Mp2DWgeKO35Legn
lN5yUd7uuz77X+1SKciOVIfa3nBOjhT/UmhfMIzS8HdRpqd1A1Fh/gB0rILg
EeyQ/gzY0ZHB+57qSWiv1Uk3HiFYRIujAAr1Fmr4HdJSFzRCoxg/udUhBLmU
yKIlcIEMDGGPdbke2WbsFOBYtOY3bPEkADG5rXDR5zuqQnigoDc+VOvA/EKi
3HKsYGAR3sDwxst7YfGwM9/Seu7tnGbSvp4CTCfvbs65VGM1jJefiItR03Hq
Te8jjE91/ObwE0hmn+8PctsKOyLUdmMVEj1W9NRHGplHGm71OIDchNEH+g+d
M72Te25XRbmsdRPRZ5U6wjOZmXCFA4Ql5khrR1n+JqZtvP5YNHUd/v0eWh75
gJp1MqOw0GEI5n1VyrHdOB+u6yjgqO62yXNp/hlr4HlGQrsxDuMamk9ZMC0j
Mig4TE5ADLtR0Z2FpWYN3Ol2AkNoxsJNxlU+gqfXaZ3VzFeEk4HrxEAz4aKQ
xoWpmED8Q51Rs086QI5CS9+SaDVAlvRb03XdDr3fxNrpwypGZ6pYhEVWHBe9
+YYSyTSY0AVDCf0vUmCzDdff0YHC+PL18a8VgDccJgMMJACn9rCJkW+oM99B
fX3EhXBhrRQh/ghvxyFHWzLO2geVls6kPWoOxf6/uHejcBp/sfjEKAZFgKgs
/95i/WdfbWjBpAyQOEf3wS97tMheDGZnx4e8LzJJJqlxFuFtduoiuM3QLWq2
m8xARmsDnIL0STwYDHTnwaeYQ2Dq3xFxgZ3qJnxFUxMFHXClixnlMw7p6GFe
l2KsBa7s95GJPPNOG0Y43NXOf9AN1zybQofk+cqBMsvGqeUgosS3CdJZbsU3
foKqMG0Es+YGRzDbvLWK0tBVPipOr9eQCJrXSIP5VrtVqIQrGQgwl6ib+lW3
/fJN+uyVBO251hcMG4Ewb7GC+phkU2yNoxg/L1PBYVrRBSROl8NqKoKrxnYq
WexkMi2tV0a84R1u5I4v8ZMV1v9Dcu9YbqH82ThJH9Z3gC32tDQhqxuWPvga
8hQLcha5YUJZQ1JHpXPRCYmG3g32rm2GDLQLOoZjWJwHJTl5rnPjplE1qota
L03psY5eOLBj/0LeFyMQ+q/SwNo2OK2GTaR7nhcZJ64C3JlOd+mHve4XHK0v
IPxfMncG6jo/aTJKZDGiUtdc/GobB0Lcs2sK5+Qofac2gbYh+hK1vFVAKLT0
u2+fSSvKkSQU/ez4kdDalrNriwv2M5Iu0szs770CgEgE5ECw8tkJh/1PxuQ9
iFVgPsh4EIbbzSVWlJL3DK/pN7YhS9XdU0c+FFAcwHomOBg1T//axpSym561
ImfDYicmjlDMdNNlLDOilvk9OTdCJ0qCWsi6dS4tHthlxVp9JR8tvZUfzTQ3
/IwgDm2DvTiuHVMMHtjz1Pzh05ohmQrq1kXdo63hF8a2FZhWb0KZm406MpQ3
/mmdS6Iz1hDHZKT+ainlkmr1tvduSoqdqVZCQHlOgMSaIZOPNjmgUGhp5mjn
ihd/LyGBz6EEOASoWmlTa4OFMIGQb5/34RVXI+4hdP7MGz2fFpJ8DgsZIH1l
EoZ5Yga1pH9WZRQcERh7o0fT7Ar6/j+UH9RL30iMuHVmmP7yDQ/YiMli9fJY
agOBOgj0zFgE+nYL0T5WIf1ZoNYCx5K59spS3dH0W0RtpjM4D3cSR601jYgP
4kE3CSTgTuNrpc4tO18fOTgSPtFzs3zfn2zAIQq2UZU2+SNPXmykeSjOzgdY
qi2NsxYeo3cBmQaUOKD7hsmQ8PZFdHpU8loh8FtP+LXY7IzquW43oAj3BX14
hdVawasL4CKHch5haDAABVuK0XFyWZNBjQOunlimqFVqEjfZOqA2H+EeSRl9
k7eMObrHitjiInEYkVxs/RsdEpO7Blqx58DIrY0Xi25n/7zlmgG/zX1/Eyq4
q1W6wJix131fSGRiy+kfZg0CJXn/bMunLHlurnnsnsJi0+UEFi/zle9zMQpw
F/hmlmrgnbMZKBsp+JbMPfIgK+7IoK60Tw/PbMqNzJH2CL/CN4MNUr9hoBkw
qZEMvqNq+6XhUctGCbSMHu9Y8A3nT3pKEk6XfAThLNsWQuidDdfxojY0y36W
gfuWp1lRMafyB+mjPZCrbr8zRwy2ZhnMxoFoLhG7KG5s+HgfxNCY6RUmu3fA
AruZefHBgoEkYiSzCcvI0kgwTWoFzEYV7GlwXhXDB90tvVS94ijRcyIf/3rz
CfqIy+y8f9CTDYmSGwVV/EmR/tRCyIm4UgPQ7mNB9DIDj9BkjgcI1/cE63jN
PC87djqR846/SMtMEmMC3sKifFWMYe5f9y/tmMgQmGl3cO0uwGKhWhdNakfV
ZzAimxhqKEgYjl9ZJuYxr2Osc1G2AVC9e+MYO3ptqvXse9c9HProQg0UKpxE
VisaZZYKzKrlRNf5nXLG1wAkKo9HZBz73yH3TpO49EPrmWWR1ByQNdQwrWdJ
jmlq51WGjlxp8VOcGaybGhmZ/UdzSCn160NGSIGOA8IiRZmBQQ5Zpe8/9tbJ
v0Is1MnLCMGLxvdji7NE/1nE94lpiEP6MabDa7F9JNR4+6B5YnLtNVdv8Nnm
YEbjJg90+kB43HM/ypQmG4zLbNmf1oxrydxpQsYgy5z6KHKA8JKYoWOX6SZY
TCJfX/ONjhrCDp+0a+WlxEfQq+vPtSZJ7V3NrSpTSuEUwTZB/e5olIzvvHxw
qUPhVtEZ4RY7vtzAL7wDyg4vtiMwqAbiYs4HD4LE8BXqbLsy4WZm+eUpAB7B
9eBtw9aVfipESG9oNhG6V/Gndy+4eU3kmX++/4UB+K/CDk17XO8xYzpiXsiT
5nqqzAriwLQc2HzaZat82rd8UIKwEVBQEGjaqkJtn9F249GpExQPeAxqB9iG
72j2FfusiIAZQ056IlpxksUZDi/lDC73sC0JP905KJyACj6Phaqxb53Ul96u
fxfTGJLTam9JwKjwua5Y8faVZlhe88jXcED7zdP+/Jx3ebypyv8K308NXDSN
4BPDkuwUY6sqCIwHl7SCB203nFUpKN8vhOAHgxBNzdampdYJX10s3CMVsdft
mQ02p5OdFUSMTVTzgBsxUF8Beg7mjtj17CMJAEznL2O77HvWZudLXww7/4zo
o9AeY4ZO1EYix+tZZ0l4gE//5IZSYHPD3ecU8n6H2iNsllNJz4g8wnmdLt0E
aHtk9nujpu18Lh/RY2ZINNqCCWrAplCv60BG2kT5JaCBekfOLd3IBo+nC8DM
+uFx7CnV9TvmJXbS658+kf9MoL4fXtWg4x96s6q1EjCK+5G2CG8nLpzCoQmz
YYmz5kVlMlp0///ESzwANQy8NqF3BEkFN5qLGhJ1J841qZmGfbYmxwN+BnmZ
fmj6d7KWWu4ohMh2fJBZlc3eK2tMC3en0AANMjUfUwzfT7x4fJvjW4KMGzuQ
Hl406ss80RH7An45DS8ZQe2uQ9KYLe0vG/mX8/lAxSS6zVZKRPwahpkBEVDO
1Kod6tXJj/oiZ+e0hR2WFd2ARyzQiaH18PK8znGiYs7NdZkyEmwsz3UBrHio
UFsPgbnhB/109nYzS89CV3mGq+8HTTHqAkN/e5LV7qjvmVDzgJo5N7RYXTqL
3R4JSrd2n1lESEyOIUgsqn5EjzevOCAakLnrhhdBavbRtcgmbQ6uL/WDxK2Y
8j6fCyuoPGP57CdbTzz5NF9zA85VWU6TWPMXfvOU4SvAcRLPAX6OeDHsWlOd
34uyI2JQdH2kKW9RwxRHTOkdzhUZx6ZqzwFle2dSz3Taq2Co2qu6TCSXv0+R
gJWAK95BNvcfQ+rW9AuNZei4Gs0CFNKTYknoPIWi32FSwrTqJq8ODP/Cq7i4
cGttf/sMCyADE+l3lohuNKDTIDUwC8TFmhDVZBYryr0oC4Vjwje0j0u6MfYU
QWgo2wgledtfQGKW3jXsAkTMzI8A3X2WA1d5QYjWIzgR9FiC0XPJxQ4xFPcD
bb6EYewBhbrVMV6bAIerrh1gTt0VTOeT6qcZ2y/2J4OmBrGy3ze4FSISXn6U
4SxEjzXTeNT+4KzCTUFKBi1PxqLsUvIi0h7cI8QRofA2W9hVjUXNTzkOu80D
f9geB19RN5Qr3EKwYuq/3rXaaFQcpF7vmAbdRwqyCCCAmvfBf6UDUeR6Id7j
s8ZL6m4o/jo47X2gZq7mfxLPM1kUfZzrR5E5zCwTmOa12yxFevrUkahR/TkS
LgsAtqZYHOwugqu2+lrr7mHTNQuZYmL5Fr5pyL1OJnzysnVIxWjA4TwLnHcg
Ppot+hD7hxWWOMjH/rIqZOCmU4BOm7+dz3kKLP0geUE3B4WYCCv7ThbIw8J8
3zAZNNulRdOBiT9WO8nqU6oK6fG/2xh/ftFiImrteslg7OohMjHB0UvBzYsJ
9973JzeYmF9Of1IHXepXhvHHLKXj9g8/WmTe+FjVbQ2maIFq5vTxinoQDcj4
ifckCIu/ksO4k/xDC3i3YRHAF2fMU96l7UFoLC8gECMKl8LP/BGXHyNejaGk
QoTXMGmbiJ6DG4c0FW8wiaUkJxdoFjsXRw7EMwx8aXkxTogaeyzBuMlbfnyK
vu4M4gASoBwG+8IuGeBXz242MwaBUmwhauNGGFB0lX8BuWDADN16IAu+gKlb
0oPV1Lbsxmu0Yli69HPSsDZ9YF5TqpgztiCl8GHamHDN9lqBD8Cj9bbq/WDb
eeXfHmUqLXBk2hWITNu5kZHMA/qmhsG0hXsmc9uRe90pKENA6jJgMdHvDUz+
mjKWg/36K/vA0JoT9QO8BY5U+fIN6I1gkwAo3DTxrISlYpyRvEdfGtpfyLlR
+grA5jaJhdg/Yu1tYptRJspvqrXGKyc5jADHo0QAI7BkVOgfuVjMAVtMW19y
nFV4Mwg8dCBT2UoC/d2bAHkrJ4IZsEXwRu1ql6FWghjpmGYfw56IRn4duAZf
nGbuM6/OzacuuiFFG6GOCPbymxUMV6AAAJB1BlWfzDrOOua89cPTyff1UNAF
LjnufUVQad8qdpl+BcIYOPLTzQJRmdschtIhY/idaPFH7seVcWOx05mdi/lG
cwVBb05b+VEtvOzZIjtHB0woxZN3WyrSKKvZST6+abx6Tf9QydHXyynyUvCE
AY843OC6JXPpGTF4wcnq6RZZHIKlpLoLEpBs8+Q2kzsVbEHMrpIKB2orzV9v
UV9DxgTpnCJmMNpWBpIxn1kWPeVEf8DhrOCtTSC4S3eEm9NQcVAlBu+8eNYa
rkgJZYZ6XNiTRrG0B5pgUn4lQwgHaCiAhs+dvSjthOWwoblVDcICAxhtvJcv
mu/HxAe+PSgNN0adiMFl8+MAbzOP5dXUgrUYDJN0eUYKelk1ACsJSqnahb2U
z8Bqt/zBwCMS2TlMjq6t3i54yMP6gvTcRwjgIB6Ux33ejwveQnFWjDanlHhQ
dvz6ml7sAJx4oto8aQwd+W4S6muObxCEYM6KW0MSO9FJxwjlp9fz1fSLVvSm
kDLETlZ2Jtfhk18jzQ13ITjxTjXGb9eb4i6YB4C4UOpP3aZ4OWDldZpR3P9s
w+pSbRGrrqNjqAPSQ17X75tFTwkT5wa5J3Fjv2NDSbet+ZH0GVIiQ89X9VHl
ruZmzjCahPdZzho77J7LgVURbKRQTWjRy145OpKSD2iwv4oCdBOqcFtP/aSC
TN/RN31r2S4bJQKac41GwovvhXHTJLaFtIMzI9AY/Was866DbtgFWO7tfw6Y
tilwngKBduwmTw0P2OUhZlzrtrd8/j8PKsPn+anRJsq4hNwcDgiKLnuiszb9
/bJSuZoecA3H9Ke15SwS+0lR1Rx7PUzqzGTXg4/TvPVrxInI8FrU+W5+cCnn
lVpDEc0gxisfG3F3mfbRt47XZw1T4lAAiLbWjI2FsJQCsMOE0aNzM5zIYPQ+
BEn33eGcGBJQm8IjpkSsP/JilbR0xba8O3xQJKt6G59qOGH+J4+DytONx19A
gH2CpWAopx12lzCkNq+vYKv3uzLMQfqPG9kFw1sI+XMohtcCVGeVaqqdMTwX
iuPaZWN0HG3eRJd57ZpRJN+/y4Z0lJCM7IyCTQ8NygUQmcLAZXuwtIwYWqYy
RMFgSfhV5IR4V4hP5ALCM+FXNyxReu/bMgsbTEjxyKbapF/2xEBS+n/xkFf8
r3ZjHEB0BtKJR7u1w/SGQlHJvX4DKkHNXwmsFebh1Ggp6G5UAoZLxbp07PWM
F8tplU2OAX+NerQswrV5JUpQm05jJls02RQtnzRZSzrX0cHlg9J+MfddVY2I
DRGUawbtEZgRZwlze3pcOUlER72IO9vPjiI9Q/cpVvN8a4+u6SGdvKPrGOvi
itXZBuHU64ftE3+rN70ZLGzO36hGvTkWI0H+rVGHMDWhNV9cxUIatUgtntdv
W5hu2lPvicjIDA9ChKOVzHLmST5x6lzJbAh7HLO0ctg9SxJdV2z+OD5vrDNd
ZJe6xRyXCiyc/syjW5D3JuACjwE0SVbU7r1Lx8uVpDsU/oNDbM84G2w16Kur
pYZaMXTia+oi/OInK0c60OlZWcjY9IrIwyjGrdfT0XTNAr8LIW6yiJtbr/Sg
thacZF7PTF5wuDHZxF3Rkdr4GYXOukWjQTu4qlI5M2DwkTGC2BXjsYJIX11/
R8nwBh5FLn2arShg5Tdngpla28RsuFdVFra5qkqh81LUVZTkDgAetVbCHCjz
1Zkv679PhcysxXYZXSouBprdazlBtUCtpvYV+tC891vv4l4JjGdScsiHG9wS
LhPbCBBpKHxnBLmCof/6YDDuVmKnDww2Hqb/OiskTSEmfUl/wlfLjR6YBHEB
zsDS/HnkRTWZ96ga+jjoHdtMEKGd7b8oSTirI6ewMTImja/uEluPTr7Udjdi
sa+RIbG/bJYXhuJzyrMUONIcECJfTs6+2WEv32NTep0r5yFCY7ewQQylxL/f
YyK63uNohe41/wQLHJKAEJRge07hWqWNmKwu4r5d9k5VGP3JjNhS23H8tGFN
1Jy+4b2HXT7BMCqlR2QFgL+gdp9sjbR/NZC/noGEw5JfdAloE3/eysXX4LEi
KxF9Emy3CREvWcNDCQUCDQaguPl01U0EM09nevU+DaSC3G0I/inbrL0f2YkM
sakLuujDJmVZdpOxKJ0xTEsglmS1i94a6wB3/klA+HOj+6FDeHRPmVmRadZs
7/e0hEVjYD49UKRGSVxfn4fwHQHVMGK2MYVjw+6EjKbF4VVkdLE09ykXIJj/
z46VLddTQW2xEGECeTOfy3KPZD14iAx1thU0nVTx7phzYxkDucDMY94wUMFR
9Nr5LwiA7OnBZA4PSkUJpH+VvtkHKmk/oj+RvdDcD3WsLhZ4aSuucN4jEGQd
ecBKMU/HoNN8Frozshg/oUzultExB0ozlxzkuEVr+KoZSu5srxKqXXQl4+cG
rYSc3RFdaQSFNYmRLEdJJjPARV20z9aHFN8O0Y8CWXPK1GqAe6/gg8ZXEDDk
bHT7Ai0IHdO6fI2LE3AY3ID/JgMs4ubivH5KbRtR+E7CsgrmLyKspJfzUsPT
eZfhvweQ1zcz8VAjDbsk0yVapANPg1+cc09xipaNKfya7E92QR0VrFo9kvd+
Qsn5dSwheHOHyO5VQ57ztN4oHJ6wiCqQ+STB9pVnhZ+z03dsC44x7VkXeaCD
NeUSiRgrbYdCu++X2sVrrh/vu/Al3Z14EANyUVWJcDHkymfem9943CYXOapS
mYANJcXQ7QHsm/YSlspwkeBVY6Zr23jR6kCMnDGGDoaqum1IQcGrVXJPUjlM
EWmkYcTRtGnN09Zwoyas7q77aqtE7+v3jv2PuQNKEoV2P1KF7dc+9vfVGOf4
2amsIPAwBn9syetSFCtNyT2L29fUyTdu6pWRswLUUG0tlwRVlBNoZJHMmn3d
EvkIctJvAx0azZSktFqAN7cL0e9gc3sisnwWT3cZ5nLBrZDjoT9xVKBukKQa
dvlCZePxnZnmQIilgUq2NbJ72hWyLRZejuRe4auem7nMtkOuKzcqjIHKTImY
1E53Zxg5l0ddPy6fteSctjML7Mtbme2d+PkeWV8rpArky/jyq6tDeMdCszC1
QyYvfJyMif6rzIx8bX81TvXdw6YeNSIQcA/rc1lsKToJfFPORahqf+m8g7e8
ZnrJXR4EmkncSO+pjglZz1dpO2Y2YUmFg/aDsDFoVM7r1AmYU5MLXkc01O+L
M3PGCGjl06Nbn+Kz9SqqM0vI39Wf4ql+TmB3/SRN/JD4kljypDPfOEDbnGja
r53aK76Te8zYvcFx/X0D5HgIFn0sXQjJ+tRplDgQy5zAdk58LxV2tkXaz9Oh
ZrNLheAMHh4IsjRrauhDxfVeCdv4kwhRR4CguVUW6DjB+OcSymDmwTDE6Q6v
udyF6ncygGrTdhw6Siqzp0tFGSRpmIsa7XsAMRQQ9udETVE1RK0zRJ1GqZub
tRnxGZk8HB138ZsM9a/ZkIQejsP0xadP+sMeTS9pRMzoohBFh5q9mwIE1HyN
+G/Tu6iaiogrlQFXporRlkp6Ki60yj1Kao55APCIo2sc87mlNSC6tFEfoMMn
0dxQ+2anYC9/hr67Xt04ACczEvLk9BnrVnwkzS2uQH+ZRuLeeIljTM/6dXXv
7ImEfieGbMadBvhfKIuni7CCI4ULQ/7a2z8AXHC29jyXzu4nuQ6nUnavuEy0
Khg8wkDATup08CuAz0S/2CL8FxR5/aZnaXRbxkKlQM8ZfN6alZ+eVG1CQxq7
Ogp3dehqB0yzGEHCJ4gROtp1/WX7TOLYTHw/jjn8MLqjdW5pePl4DVLzEeKY
JLosc1I1OrPn9WeCOM6JPl61RGCeT2vbZN3HcZSpNVQSr4Y5SS/Y9dYtqCsm
GYV3JYQY3zk+2Hg74haY2N4OYm37sODgFFg3+HvS2Y00oc2tNsUOJECYcZMP
mAWy4fGOdUJIAVOeVzqMaG98yKmwr5nRdOaqz2UHvrIFDTtrGLBvlaoAetBR
3kgH6BPTQ/KgxjgX3olBcNlIVz1Qo/lUTt5RVo+Chu+oIe3jnEdV/O/Kry9Z
gvSB4wAMHfWvH/UMMMzivhkRRCfBzhTz8tapzA4faP8FMd2iTPvuo4o8JLnA
mBh003pnNDb9E+AI1YtHOEHB4IGBXnbaWZBo/Okbkce9PVE+yMSuywqhkunE
SyWEgwFLLgSsAITNERJX95sH4OK5QYeIs1b3UkWuBU22MmGTMrNza025uccU
VX2oUSBVsLSTcHCwkbM4/elSDOei2pPbT7wJeHEnuQ/+Sphswoc6i23hEqZh
QpzyCID5/XrbcGMIGP8qzYnwIkxWDLj6ArkXvDZkfAYhzohJQcv92HKhIU6L
IKQbOmE8xqHaYK7hMn4o5t72+yS4XLH1IJ1O1WQaL4RRMkyQ54m5ga1nQurk
8sDw9Si9WpvxQJSHFDK99+tFdngAp+Wj2erKSUBWh8/CxtK8Sy7bFxSCgyHS
nKNrDqw1pPHphmn8K8tBkJKVsbpYPr9voMC+xeg3rVCD6ac/TMBykNTrz8JY
y0gXUtzCocKq6sQAnfPbrfXnvvCFJ2sYCYdTSDgIuNDDzlFec0bKlKQbqXfn
v3LbjAA/oolWQTsL9fZ26sJnFYFOY5MELO/Bx1RmapiwoIE7Lj25akgsgQCQ
h9pXxBsxvFotO02TyFxLbDvxh5t5Kvjlndi5WdRoZiZ9YSW10dtFX6wMxAsF
OizRzKjepy0MDQM0l2c+p3fwwYXm8OCh+N7RKFg/f44cQK+9B8L16L4+skVg
1aMw4w5YYPJpBJSuG2SQ12XmrfjyeDJryEmx259TalEDb38xI96UP/Y5Xyaj
W1jZKRltNUztN6+7VYRtZs9M9XWADnIbBYFR9dUAFYxDI8DCNfPidqzBNUIv
FNmlVMuEdE5+tV5ZcS30LdwzAmsLmvgI0CmbaO3FXAATm41lIpuKPNClAfA7
FfhGgpGgZHyERrb3+FOBFjJShTwIMfackEmwMtNYS4nPQQkm4fZ8Y4Sl09e1
kf2AUYIW2xRyT7JeJfyzVEpE4rSYbqaYqH5DIOuWwhyHF+CMw2e5VBGfVhf6
KHqih594YdPy++hxz6IPmN5umL3hjAhBWJ72J6g/rmLlJWP1AMCkDU/emlW1
fJjDzMpiiOmSziBmSQqvQTP2BYo7wliX2qYXJOpIaV0I7w2ltkaBd+J9zDui
eDOYk1KyDcRJurLIvd3oQSTTNwhaMAucMe6xEHQln5viimhpn0Ho2kvq+r/9
fF5p8jkbLX19WcmoWnn1CvEAhJavkhMMljyB5LlyBq+BteLEy90XjRiTXmpj
PtqeuEzmjymsgXRpeQv38CTur+bua2wKt1WczGeyqdPYwLEXgP90KXfTmf7e
WFVfdcIB3jjCys8vhe3WvwFRlClp0xoZavNOfWrT2gOe3XIRw8ADgLccEpQW
8YvwW9JTwNdudoMqVSnEZSbPWKofrGwu+YZ9RyGIJNrpoEHSFVZO0i1O+2Mm
GNytuqAsQ5yCBr4D4QckBD44I42BX1oypZAAhztno1TAELF0h3H4Fcad89J1
qz5UuEf8/N72VCFGpoX6NOGr8iTFtCT8u/pKxrUyfrrrUfuMZfB08cRjVLZU
G8HOC8ZvLlxCe764gCrf3yzv+DuG7i68fLECSLe8FeezL7g9y2+dTNYBalgT
DPLK7QoK5CyfKIRUqGu5MDYkRUojzK2uS3GsQRL9dRQ+d5CkyHpeStu90Qh5
jd5stlfLS3zQ8v1ZY9DUV32830NyAY5SU0mmc39iWC/iwBNIJXwzpC4Ms3Dn
mPTU7u+uxqvIwZo6nCftmVpZDaIdNlVK0YRpJhfgqwwYi3HNbHTgiJ0BC5el
x3f1sjS8WV5myy34jKAXmZAt1f6wSdhoxgVEx+4XTqDfH3iCnNHGbb77dnws
d58xhYg3NLclFnearTw9s3n7dgqIafqYY7RBarFWelK4YEK85NmGBp/RKEgl
PMX6+RCSqQsQ3kvsX98B14F2Zp832bDCVL76YM5DG0JVMWGJKOBsgpoAxpSs
UIJwdTMe7TA93bLIWFMf2+q7WcNNY26fZDHLutMbFGOuXsRKsMj1ihtmYAAP
xaiGas95pg4zkHBxvxIswMErMXKKDkrBXT90p3CcXZcJXGevYG6dAOwVIlif
J8hd1HLjWy7dxtsPZViFhHE8s1E2WOlGPBJDWHIal3M8kVuBVoe2IEB6A+Nd
UU54ej7OpptOOyFSNChTvMsMBouXOToSCzuTvxSjCn56jVjbRFI7fMc3TZjQ
hZQaajz3cQLjU0Zs5umamB91KmGq/AVJZWrAtxr5WNk64q2Cxb6fP1hFVQhb
JOBFmCk8MwQd984N5IW+5Nvg2EWmpYQLdHse2z8qT3meQouptucKYWCWXvbB
+lcbax6yNLomXTFIfmx5B0+ljE2LT+lK7GP0TaJRHhlrf+kcTC43GcwR6rKL
MHips5ikS5lta6NN4PsHGceYpoeJXpstdhjKkz+tnk+4ArG6oyR7PjYtjeoC
li9heE3lQx2yRQLqq1S137mKO+9j4kihgVGIW1bXDTvpaZ4qX0iIs5ey6qZe
6KsfV8irCPazvqzU1AwTR+4cWkLCQNRT+WfS4zoq34NM5lkpXAxG2R4qzfJG
6XpMga2TdFosivDzMUwj9pL/N1XdhOmbqhId0zhgkEwcG1NtNLttWVZnP/H3
LsLjmZG6V1xEqS5hAGUz/+068FP20fXGXzrUgJu/vCkEbbsQSmH1zZREi20U
L6VNHmjgH6XdshlIEZSWk+BAenj7x/eHfefZ+sVmgcgSsjT7NVMPEyKyU0Tz
EivaaoEpXckA34O/wRBBqPdwQkW0FBp9vB7iYcU1Nmb7vrdI0at0AHA1C5kP
EAhockCMxLrmDyc+EjlSL6uQlKBt5CMt4qLkfH0kFeOoi4oJzapN5ZwOqUFk
VPlGd0bwfbu01/uOLve+zXISUxggfa0xfZiWo5cVFW7p2tnxapDjuEB3VJf1
bFucWgVRilGjx4dPMqWZG20GjrMak9jytYFwPPUzVuhfYyaAu/vERoLPT53c
23FL7h4PxqitEL0Ie7GP01WAyEjhI6Gr2FDdJYCPaWZKZu5DcOUDefjI0Rp8
vIPwYFuN1PwLqhhhI3zHXqXMylegjutuFszTnOruOOap9KUT8By3j+eU1DGr
XfOWHmynuMBSzVOyQeoEsCOYHTalPrAye1bJisLtzqMmd16F3uGaNqi9U4Oj
yy0dUuFKZbhnUTA/y6Yq0Hy3PerhHOIFIIhSOyRnugkJuV4f4606GOTBC/yi
e2zuSH4yB7EjDyNwyMurEEHZUySYzRi8Mm+YfWmE4oKOWKxBHL3Gu1p+i/X9
QCQ+3wmgvfC3hUIBigMjYvp5Q8NsOsdqVV+UhUKJ7pmkC1pw00jek2EDXer+
QjO/sX0vxTaz88/X0wr484F1+uI51JYlnPSshVCvFfuWefNUD3MEqx1n81z4
1Ht5C9oCegCvVrOlo7IVpgX5dBulq7IVGdcXKGfcTKN9tcdzpPQyB0pMzam6
bDwTftil4aZjtX0NYbVnPTBUOZCG2t7PxfRD3T0y3kMW3Kq2u+jQrf+FxxE+
UiPpOm/Ky0ZqwF4JTcAu4xEvyNuWNddykz41mKpbi1NEeTwXt8u7ZXHu1Dxs
SaqR5RrCX4qUuoWFi28JnCNiYvjVI7QGtVcXujSZES6mhf1/q3Fi6DzvJMEI
CuFdeASeY1EUrp4UIV0vPMvUHv+G+UTeV8jiVinNV9TK/we7gAOAHdzD2IBx
WJJE/V3EfOE7IjkKhbqf3OHc0RMaVM4yRS71Mybnoqs0M38dCleFst05XQ2n
o9a+mXbCF6E6ztOrc2r9OXxj7+IlLjfIWifJh3vrGNGeAkp9xOWgXrJEdWkt
/4wAFGG3PS9dzlFTFczLFa70Nsa/ejt58AWXYm11h5tmqF2TJZDajya4NnOI
xS2Y5/Ihq4lp0AXfH086Eks9Bfm907Kwtz8UaU0iPycAs0CDP0FiIYbOiINA
x1SS6+GdTW5ju2kklo6AlSif8pyMsy919awt2h4vR5mCB3ny787GkGL0qU3w
d39Tfsz5UZJpPHTUUK757AzNTVsyzTpKnAG135ay7tHJ3ermcyc9lG2DDSb2
relZcLC+KHL/NBselwUpQOU0UYlwPVCMJ6Anhyp8+njGpzPxATFaql5D7DXN
8RsynI3sxFXRkEbHXoxUy3WkK5H7AqofN+aOSx7KuS46wChJA+Z0z8NwnUHr
7T9vM07r1u0tFWiO82iy+h31tssYJ1tnXPlymPLfcXRa+n0oQ+qa/1JP/CK+
XPSJma1/Tn3DOSwWY4ky/9OtO4xhyILxZk3R3zsEbfpr+R0O7aJxVEJuOQQz
cksVTPEzTuPdyNTDRbhSnczwSwfrzpcdkRyQ4f2SCHIhVVBwHGYBOos7ACVq
PJ8YybAUVbioK+REbUKwL+07NMYP7PC7tfRjnHqo6yBsbvzGmw2kCyo9in+A
PYyUALWXQ9OLev4gbfmpxSptKhIa+HkeF6bHYscVKFpC9c0SqLklUeKx3DCI
8jpjPRlmNsfUr14B9bRot6BXEM1KBS6v0AVG3Kx/9KvUK93xKMqxW04nTCda
ZaiIO0zUTX46PkZe3QKk2YhmpcVUNcXJmd1ZEIqGu3EFiDGZDDdXmljiPbpF
S/hsa84DL0jiLxvU8P9fYEeyZI0Et9k+Jgpo27zLoam0vh4iy/6b7sRgq4jE
6z/NR3xHzUUdae6mWZNLKnakcA1cvE6Vb7xcJaiiSTNv1sztZTl1bZQksw39
skLdJYzXHAvO+bkLTWnwfNLoYyb+z85L6mXJvRm+MCAx72RZsEPTcAe3SIlr
U3k88rzbec5ii+zq2DiNVyCk2bhgPWc6k3583wPt3YP5zloSjVGSV5b4AaAC
CJ4Rxtb32cMVxh0lkvlpeo6HR4iD8ZLBX2GwG6V4Lmo59ufBuf7ly0El3/JU
hLxwHIYnFe9cdRNOf2O4SN+rrPD7VYaUFKCdHBvcldiGfcMcUjHE+RZS2k5U
aH6eqKQOPIAyWbsmkxrgmgzyuoQMZTulXpZmz7cCPp2eq1EP3cl/WL/bW7iU
/Wd/tCjnQ3woSoQTMQm1SdBcrJ8WOKS7ld2lUy4YbTbHJoYoaMhfjMI/n9gb
psNcHwSx5+um3aiqG1K0B0mer0LcOIv3CKGLQwX5ybdMzPpplJgQ0EnvNCdE
JPne9zfchKCgiC/3R49c25pBZIsWz0iDrZtliFC6oI3uMDJZkd7e+J2/sZ2F
+p/Knyjx/bPFqcPa3aR3TX+mmMVfedhBAXdkD6l9x4EWl3sxSbH3GsEM1mky
pPJ4TSzXhZ4gOBqgHhZNSD9NDbokxw1etuypJZgQUwEIbu7ElPyWrZ78AE/7
Hhi6cCJpkYHcQZ0ORGPHqvyygv15bL4s1EeX1buQvlKB79Y1/qCkYlHE7/hO
aBR/bBVSjFHlXm72rq4McoSlqtW52WVoSTVRITSSBO4DQKzlPrsRXcQWna+i
zppcxkiFQPfpjzK7q+kOHTd2FY1cpQQ8vCsyQJ7eQYHMVVj26FrjZMsudZSc
g92YZ3t7e10MOE/SeBJ1fTHN5oAbPbLGCjVYPPrbHz5dwdmADfgrhhB7sMDV
YEWhsNQ4SDGZVcU3FsmLKimZW65PxXDgC3W5gFVOS6PE5hO9dZm/AwryGl/y
8QSA+XeuwV0vOLmmbX3v95S5mW5BlG9HiyfcLS138fuRc8BlmT4JLCa/p1Xn
HVtL4OpUojQsdrqMoj7NQhLVOl4/iIKB7/9BU6hw6+yvU0VRLCpa1V2S3eda
H4m97S5RGhASrOu8vPLxWWD4Ehf9hN22gldaIwZ2Awx2P9K+gQvJUYcaFkoU
jr2QOSeeN36zmKlojwPHtAM/wl4XDcG8WZMya1pOiUVaMdKVbNK5qH5XsfSC
qUMqzA6CNcgyAfVazfhhWxipkrjvTYL5lwrE05l7w0RN8h5iB2ELoF3tiWSh
BYQcQ6h/dMFcWtzSPHMgg/fqiAGBf4wKuRYti2SY49tdt64gyibx6xY/CuM/
REJ7FuHmMQUnOpV2HtWY68bNSmSUKSW//I0a77V591mSXfFPt/iADwMpZ7kO
H+yUhBX7pAkxaytupZVzNqeXBNuKi1JqUFTZG5tTnH0FZJarXJdyiY9PLsmL
HWDX2g4jagUI27IJ9fMvwtenJ3QYkl/teKjmBoK+5sTxIgXGnHimOnE0lABq
d2cdb89mCXcmkSH06rz/fcwKFYSsZ1lQIvAuwVt28MB/M0Vsw+mniDdl3E3t
lBOjq5FwBNSC76xc2Eq2xcR/DNkkWz+sLj0H5o9WIemKqcNFOH0PRg8dWlCJ
EFQgx6MPIOFRDUbfj1xZf4lDZc53wPNHCuq8w5Zp53DceVjeT/EeuR1oGwJ7
2WMmhU0eRSXHh0O9vV5uKf/Z4OhUH8yXJnEVWNRWb2PsTVe3yP7kxMO6Jisa
CH6rNhr2sQAi0iqG4W5RVK5gsq0r57fLU2lXZu0p1CVl1TntDUY838VQqcIi
FjYCRGehnWB2E1MIT1P1mUj2idQJyYDeYmkZN4bdFCjikS53lW46QyohKkxq
ByXa2fqQSQyNBIs1b7u0NHs8G2ivyVx2pjr6GYeiphkjWIitODVeDnzojRAh
7ud5z9rkVNKT5wyX1zUoMBYBUcXU1+AtYa1tghHK9rejNGThsO8iqfEaPfA0
aT2vo2b+pvOLF/RjYObcNteLodUvEoYESUgZzcwq8MpubvrvBJp6AnrIgt7m
EKQaKG+yJl1s4lZde7c+x9S0AgcFakkgOfQHprawECxBs3bKHgvTvK3TYK92
B8514FaEQFUtYsYIKzBUcbgD28FycpPbbawHgY8a8zZqOsav6sgZq5YNlI39
qmKWh3RtAZFUcCXMPaawAfZ3yEF275ZLd+pvGdz9/CzqperO/nv+JxkHV9Ow
CHrtnlSvq50h6tngQ0wfFjTwEdbeYqICjp4HcilKQQ72RQlWyS3YCRz54vrR
AE3/HBonlbL2Hjtq5yX2/jqqF8m0eaFtToRTx+Oet8/gXRImyXY+5JbDKmsw
kXNn1Kl2YpIp4ytnloqprI10Sz59eOS4Mkj3g+IICCFUe/b5CuqoRaQw4uew
2fPNpXclP762t92CcVcf3IZYkF3RMPGXvIcUocMNl1qTE1Ur7newx+X3CT08
hj/KzF1nemlD+ZEL0yvYrr8V8lebIZK+O80HxD/EVw2hhKM+eU2gKvnl1g5o
gYb5TeeHPDMZiQ/ewNMgdxi30JapZMGYBDl8gQriDugTA4q8aDXXhWm5K1sx
m8A+i44gECOkZwW8ZS79fgAHnGnHiOUgABwaEV9temzoCJnMcElHe5ktto+9
L9Tod+qpc+g08UbqcNmxokUhK9bhvmn+jRzzoIGK4RkeBRQWV2MqTCC+SPci
GGveLIcSM85Yp1SImLnnmG2dh2g8+lNwPQdtIXX0bXQHeEAyHkvZ/YPzN+dP
w3OY+BeGoWd+T6g0I6mu8OXY6tbQCcwQMl1wgN4TLn4EZWKT9ME9VeomSG3D
cq4dMR9xp2LVRcyU+esxJ6wFlGclVXaEhqWsqv2uICMPrhDdOoVnzsSUhUN8
jflbHrRs2Xwk3gkjItx+q/28/s30P7c5ux8LYjMqS+S6rbCw0x0cSaSO3UiW
ravNevE0s9qieLd8aIGkN8/2HNC9C6MLGakCx8cQqBxhrjI9ghqzy1Q6EoZ9
56B5PL5HbpTMGy4KLrdkAqjV94TzasqMsMFheXVKLkUX+kACi/u914TDL6Rc
iebJYtwkZiIF0JxqeepWOQSO9eOr4gwJ4A70momHDGpno10+ZFlqS3xgEoh8
W3+vbVDjcT+od/PRLNmaJ3e88snYHVwUDPmcrrDruTuDb0eZQtdWEFq5PFVP
sWwtgzodDrv3RkJ6sjDeOZp4zelhaTFrW4/OclMfEHm+Fdk53kR5yOVwzjgW
sj7G3H72lUUdsYBcVcY8OFI/AmDOvGM8tOPmccW+pBFC4TMd+mSpI93yPW4x
zePczQoLw67iUppEFXa+tChND8D6hJBXu6bl3dj/1kG/Ij6VWiYpAeyTCFEm
UyBFo2VTdVZavKWCS5Tz6m9rMhIV68FFhnsZhIQGegjwjcQHvwoB/17XLApb
t56dGJ4vCEADrbHYFG20BEFYC/zEIhj75iZxYygOKB4fn9tmWVxGZvGZuQ0q
FahTEr7DZeLY3zb5DZWjN96m9Cisk3lDIrrms7Y8tRTmMniWiOtKdh3cmrkA
OrEcxcng5usgHLN/QdFopKaZeLYTS/PLNi3p2bNS7M1i/fAG57g7LJKRQr3s
UzFJvpquBxwbB4252Uy0CIVpXafQ2B4XmVwq9Sfwy8JFqlEG7ZczVlM129He
gkVrpooxPZTDSY5TTjuCY73ctGPdYm2qumjZz7Si0WplNBTo8/Y3BI1HBmkd
QmlbOToelaihIDqJcL9LYSD7nOz90+0mI0tVE0lsxu3CbKtOxbNcgwKDZBxX
iGNs5fuZ8PARVrPWhuo1dH8fL9NccPxJd9m5FWHD+ilcdb1j4fo1Fte3jZE3
YXGbJetakd/CyqFntMqwB2AJOi5wp2xnQp36ABlxhfLLgbQRBPjmVxkRGusG
dOqbfGN+UiNJULmxzcbYopJ2Zy/wTSPlHHdOC5N9VN1NjHcISdLiCCx7aICS
yiE54yboMM8lt2RRRyplmQXSzeYHd0dfxNCFKn2fCqdtPXUxxpfa+p2ySb8P
xttM2a7sdJdRMA+f+8fMbDMSidDRUM+COPsnnEV+i5vn1Wk1KFrmXchXonH1
Zz2Smk1gWF3EFCSNq9F7NNPb/5WKoceEGoddIr3S0IoS4VW9wj+8i72GXKSO
dE42TCbN9NFHM4yPtVyVyfp4qzmNexRutw/y7zW9uh+Ssnx1E87s4kS/9tjr
ffR8IvMvk1nZHLokSZx9ixg9omPCXVZUufcXMz3c2kUxOUXZh1VoaikIWssh
BGtMTRMzFUY2DpVfuKb8D663CgkXmpPhXLLAh8+L7Qe9xomOcBVBX9K8zeR2
Fe239PRC1MvdRwsplabLCvSPYG3G3z+H1MMbd11NoxaMUvtnPtCgAz9wtagg
5JsTZ2OoVpI8CznB9IJqVGc7IrXaoVoea8Gb/QoxpWQDdh1K+emGLwlwu8ym
7KUFkJBrhB+j7nXkSoEAaLAQ8WpqpUqOoBASVRxh3ZwsaKOIS/UkxYLfEhrH
QOr5ydhiY9r/THuAootQZaEPAGwLUQrta/mkqhW2IMSrN9OXctiC/ZGNJTW5
gZZXsYMHwWvR0X+s52lNhhqhVmNCiwqZ/3b7w6LCnx9xwFHUl9+DnwtDWvxj
8RgtAJq3TtmXaIJubAXBPvv2q5NEGiV42uEUTuQ8wgWEq6VNv8HqTROyos6b
fzRNcOhqS0PbKwqeg8r6sB7bqiJ/GSFzbWjkHxZlqw+zN4oYskYc7+vMAvfH
9Tp0qveMfbjoEHqcGKFfl2Yz0BnRvrwv0VgQX9HulrsmedlY7MQv5/TH/8s0
KmB8E5ROvGeCkY5qJajNaRgbJZbMIEPkKiOf4DesnClftic0z6OJZUYg3Lbi
YyIGh9b279EMa5uOXVE1CY5dXF6pvU5MPmK2LvVjbSUekLIAkbZy5+B4SSES
zmSg0m+DzLw5cal5UuVqlHdTftpNOCW6meq/jPF1q3O/A1wAl/xLqJX9ZEXw
KtLm8DOIluYIABGbgLxIgNY+uxo+siBEmty4VDDetmtUNNvrXgxHCIqDO/5I
MQ3vMMgGzv7mxngvFK1vmHV2NWNps2/ums4FT6LxH8F76BdSw09mmK3CC+bc
/Gci2RtvbnORfbostxYGMGzqa+0D/RBb5lhAug6v1kxvuOB6dyRwOrXjpnqa
YPYNuBU95r4ARVHEDJGlsS0J3lXt9/cTMYICgQ8FrDnOSUQoCsSkgDcq7NNv
y3T0sYlyu2aZtzQADdMDFBez/TxhvlIoZKmgO+wlpLHCJKEDyCJ6AuoOpszO
utnwJBltVuR4Xj2TmQvUY0Kc+VVZfKnUgjUeC/YCwqXCLxDa9bxDvnBmucoy
nOOrUQjZAgo8d+J8mOLgqNb4dlEsqZOR1aEUYm/yy9R7UMt2xDQZ9iRcBy7Z
tF33HfcFsIzvAwzcnYLAuyeDTUNuGbYN44Iu5B1e4OUqr80ETrdVHrK9uv5p
nxlUDo/ollQXNYZjyUeEQx2bodjHK3/2OkuIF0KbenFRAusYBfsYPi85OKSb
/DNQJmIY92M7tvHbsxKd3FniP6hCsvyEZlkxuDhuYDd5bW/PAeCfUcKnmYsx
ck+1Q6qCaqk5dmCLTr4Vk7sZ5EJ3QmYqlcEWFFSaJG+wahuYdURQe6C88hJM
+OvfzqKnv+KsQQoBsm1y2Xbu5lLPUwyG/fwAqoisR6fUS+fjK+JOjpkcUjkB
zq2F8AQItN5St4K44h5J3j3Wd7JSmWle9sfMyz+faknZfZ+8ENW1Wk0tm41f
2r/CkiVds684G89zyKhfGtJBK1ei9aM6IbqWkWAcDnhsTb4ZfG5NzmMijK+c
hvwA8BJoFIEH2DXbEkwk4W+eO14PVw3it6Nxne++WTBs2IM+KEcPJq1deaGB
T2nXLQEazJdtVhb1D1tmrOFmYhIEc+fWHEPTVd//96C3ebCzPCRB0N8Q+vB/
OfiIK34mzHszENvJT1U8D1pfaU1co8/WAELG2xJRwII5CMfYrByRVo8TlcVx
gj3ZmravJttg9qJa5w4HaLn7TzAidIYRuckAj6U4VdhLHti8gupg04a2DGwe
ExNeyfg5nBVXfZvlS4AKUjuvpdp4v8ux1STVsaqhveOdmHhBmMhqfoBPfilZ
72zkiiPbiX8A4lOZ+vL2NgnQn0Z1nP/wDZ3WukYKZrsq06/DHTFuvxqWgu25
SJ0yPkpZyzX0TLmmBzNRQQVJJgSFnowidssm73fL2eCOtJJdf9PZoTcwfUgy
HxWAlRmrb1wp7BoyKDpv4lGzTEpXVfpf0YlcpOnvkVViX16GWE53Bd6KIm6I
UwTo9/c1DQvao24kKFYSAj3XYuZhimeJNUfFQc3ezbLuhezUDwtaBiDW1fwc
QWTMg30o74BvPuQA/hmpnm6dxap4PK1CsF0iSKP6I88+V7edBsYSCoIFGUNQ
Wd2HPBsplmd8Lg8LA9fCjucGiVyw/L51WyY8P/sm7fccPwMDYucV7JJhadZR
OmMNNUOkNIOW8JLe/b+aNQEtoma07ADLl3FNB14MvtM5ivcQj6rbqQhHAa27
8DF5yL3ddPeFOeoJUvUCY4BxVPkZeJzFppAvGTcCguEOueruwc2SoAMjOEkX
DeWz1GU0bQo7v45Ua0Gmxd291NuWWzvG6fxnG2I0VHYT4ewmUxn8A9UZZJYF
VKgpVN08TKZaN4LeO+LlRs8B8DW26VbGKlyw4YLGbVvWB118Zm5lTIkzRNLv
s3cQBMDGXm+de629DMPPNeNqGiEqz5EplhlLBuvrelAFZMTBAbRrqD1unxJn
5uvB1ol0j2LG06I7Aw/7h0x5m8chSJi50KmKIpg0occ/w+r7ChrBxt++bv6V
dNQWw1en234RBMzabnMzDHrb0jJXN6W5sQQgASl2ftKjlFggFek4Mi8m16gk
+FND8dfqvZvwTKlSF8C6pDL3AwDPJ6Q887HNT84ZUBHr+sFM2Jd2Gns3tchD
j7r1YoOFrkejExpV/yTIKHS2Rg/cHQ2VVb83idH7BUiGG5IJkta3Rrm8LXdc
kxa+5c7FfPeqFZY5GMNsS1p+fDoKJUWen+vmmd2TT84sDjpoATMa84eVw0US
cOaLkSN2ZoqiP5pxoOB3/Ss+bXXz5iRd3Rbgt7NbPw8dr8JT48YeuFwcq2zF
zCw1oIQW+NjWhCJlUGGdnu51wU9q8KYiWSHrocTWEW2rC9aeIvHDigXXkCjK
wCek78lV+3RxaaXcVmPupG2CYIuCHVEvdNa+c+QajVpxWUms8S6bECFu1RCK
obeLChUbznRCwoRED144SX3o05qEQJUCJAISpFN0wZWfg7eIRA30ke9YfWK1
IOSWqmAQfIlBY6zBk9JwcnwQoTgw7a7Uod0J8HdhP4/ALeSh8btaAFAKF1Q6
o2elF5HhsrqUKa3oYD/vte3sE9ZmP8S7X0/QCcUTg4wms9s+4I+Vyeh5TVkw
fvfpV5oXfh3NbvKppBpahNbDpA+54poptQ6DTcvKHreEO5Ofo7t3mAhB9Ig6
qSnLeyIIwwT4VAUtEMcGXY6Fx+HogjScTvZmGNn5njy9WIxVVc+235PnNf/V
Yk43fehYysyJwsHzUbHaTlnh9vCwouC6GqgogzlJkHehnxFyv2ogUDOHh7Ij
AQbbNyFxw2sARZBaMCA0JgiXge5kJoo/CHf5yaMqfa9ChzdQEKjXA4yBZfVS
Y5ugrSq7VWCS3FPtL+qNWhFgTUGZif9rBk6qqfgcmr+p7bkkVqKjXVXKQrAg
sKJNtKswC1HUQwwjEU37ntMalzBDzGTfzi2LyALeOohOpUghvLg4Y6qcsdgl
9J7Z7JJb1P3f4PUtFDXZnFW/2u7h4svLQ9rccpaGrnQOrCDxCwO+6ucTp2lJ
0/umpNXcgIxHtpsjkN1ZGs5EyWjeTt+dEVdyJbKNde/Rj3l6042VIOvdrDOO
rbiN8cnSZ1/8cu1W8iDpehQ4WN+l8fnd3UQoCRHywrCE4Gw4LIQ1j9rL951B
rJcjT45nTs8/neYKGaWI4wgM5GVwN8h60ZyEEkTbJbWlb8LzI8TySsmwlp03
we+iPQYdWY7SwpXJZGPCO7dA0jEUM3MfhznWnMd3cIw1BVnAHMOGgJADNGvn
11HoPQXt1puj+McYi4yCxKY1iTgd//crfHllmp/cnNQQn7C3LzIYGluWE8uP
fcl4sWjuq7jVZRxYOE0KFcEV2z2+eZKESdQ2IgGiyR6zQksTS56uKiLWLm1G
9LQYqRl2yEDkVaGwMJptceLC4AIIfTUaN85cPiXOWTnzgXsOMnqyo2ptmG4y
5A+zkReRo44qa4baHLNrVgAWoyVy8UY83hncfOjrFzrrz0TyO+0ZQM7Td2/m
/ydRP/Y6ZNvE9CUVPx0Ele/AcK9A89UIy6w+HHJUmRcMi8Wbs33Tr/cDdmvq
evFcA++uIVHlf7bvZwmCZ7AaZX/3bnYfluuQuiY2udkYj0X8p+5wLu4vfuhd
JpVsdXDW7vDeEJFQfyBNDAojib7qhGmC6zQjrEQ/hH9HRk8EyOcZKhCTmHGI
6UZCMZ7aSi6yYXTYzok0HZpgJO4spHfa3KQe8Nh7Js1TQOoVN4WlwRDbIGjv
LwsfJOsOaZaOOE6tudg5eH6DDFqSy7VgEqS7cl5sEXoEvRh2iOxERlv/+co4
SCUeQDskiyp/UwElQN4Hrfs52kB4Qq8476q5b3EvX4i9oH/C0eCYVyFyOmOi
48dha2NCDjYkYrQgQmcABK98zFHgi5WXn58/CrRiW3ha5YMCn3QO0WQhlo58
sUZUOnKvPiqb2mmD0KSBDzhdGUI/bru6bnlpXG+2+fE1nT3zRCbrynQRVyXy
ZGMyy7dlzVbV9+YxrGHRdXDJKLIlFHBgGZ+5jnmaBDXBE2sepZjC0bu1SCBp
veJVV4vFKVDlInw+EXnFDYT2RpCaEmy/tzcom/ePL7+DwnGJJJ4KMQjwCRZw
Sz9ik3JuoAMvVnJGPrhN/iHkG2rRPeYrl0xiEAoXbrAo0sAok+TiVpHkG6zJ
1OPb/YPP4iaKmIz2642i+37dlKf7URnVcUBpYMP1P+RoFzpX/KHCTmlL/U1D
Q0l9vy6JQcY27Dzl88REFqH9cIWUL4HwS/VGyAsCxYGMzYCOUwT3GBNM02jz
ET2AtLSPTXu5G/KuVdczKmgQ8DJ/l2Ijl1JjDXLj6GwGuEWJVeizkJ2arz2g
BIqs8Rm3q/334rWQ8RrN+4syd7MTm3IersgsryxpVYhTSIx/2D5IfBp1agnp
jkCHWrt+Jg5HvCBDHlxasakWsPcLYPRiMds1dHtf1flv2/AaM9dKWOLwXDlP
5nFKAUbqc5OeN4YQ5A01JQqVAziqcKUlOT02eVUNBAssZgolkX3sKRu2GtzO
kAVYDKR7ZWMFC+fDDzuwfRj275e3cR6oKWkYUckXkuTdb+2oNLQa4tIYLZGx
fv5n0eGsJlR+OuyM8lLrfJauCdX6gQtrHnU9CP0a/NQlV6SuVAqobcKQ0IHd
syNAs/Rev0jFAarSpB08KM7gPFHhHv8c6pe0NNEhWc4JyHio+7TPo5Jn6ACl
NBN3RvRHMa2AFmifXviULElkbPe7BN7CYSb+eByx1kHsUxBxyNzmdHB0V8KG
+o4xV9QUMQbbnHnF/Oek1Da5SWbhYpE3LI0QBs0BuGDZs4xH4PP5Y4ldU7Xl
psAfAPEmJGm8lmSWvuZtscSMYpDYNrGCdfGpbh5EayQfZLWaw6M5rnzOSWMX
EfrevnSFA+InninNSbtccUv+LeBwrP2MiPccw6oRmGws+uSp+xiZS79gKzsb
qE1CNzINaxc11SSplfiMbC6qnrBTsdrNw7NFAxHhkWECZAoyy9WHVYUqRTql
7q5ooegV7vzH3aaMDMEWSar07kdUFVytQ2469jLo+mw+7Hl4tBIBoagdWoBM
FlBS4A96GJE/Ke112vxmsJZhifFNXrfMUIHRsLy89NAwoSXGUNk7WQYOHiAX
YIs9MvohQZJIp5KwGGPfuchQ3l2k7DyxUA5Rdt66veGUxyZH5M4yFZQ6cyY/
tZxCf6lkQViraxIw4EwGD5y795j64GeEu34BNYIP6mxMXAplkSlUJcRqLL9e
M4SR74r6t9jr812XpiVySUn80unq3dsNpvhHvxjNdochscg9HnYLnCTkO/ZV
LzzbifepsBpyYS/gATokuikUl6v6KaZ9114MeZiRFAH9OPuInB5JLQv+132q
VNtYzgunvlPblYs4F8pfeKYqPKw6koejIZdMYHZLqAMtnV5A+k2KqQXXr+Jz
uQ4MJedBeHo5WWCCYABlO/JfG1qufjO7Mb+BbWMoKEd69WJ9wCcyjSUm1G3n
p7ZZib3ES8xQ11E0m0w1QgM1y3E46u492urDZwQyJWag6d9TByXcsnORYyHx
RZ07g/bR80Ml1dwGbgLjKfTCsyuwRulqMVscAPL6DImcJrCpuQaVwMmYr79L
zLhjTCALALRhVmE0M1GZyJwAx13wyDBzSRVPknMic7nUep24voRJ9F4dvSTU
NmWHrgvS3GQ8xz5ZXM36DzwkD9kwfYw4MSuypPf2pdWAHHVvKQuRfpzzPMeA
/X0Przbv9UMY4F1xExii2Md35EpsPlgfVXI+r2coo7IUWSO9JgRx8bLqwpvO
RqyAUOKGz/4p1C/H7yYUgdItizL6HXwtjN41KCybH5NlECs5WLWNZJ7bm6BR
biVc5vZatCgiZxnhj0jPtUdvZlkv3J4aAT5v0iU6pQfO0hPt4SgYLvoiKnRp
kqvl9C3WnDyBwMezy6cDAwjs6kqo5xtjGWLtNnUqNlBtYXCKk+kTLIOsO+XP
QKrfze05cQ7DOiYq8gpq/8kDKpqpfPZcCoD1/XFsyTI4Y/3thjBOoIc7KJMX
zqL4JJi7sCaXB+FDpXo4EUwkoITuQfvsv/hfjkv9Ro6+7+3dYLU95eYyyLdc
QLqhk7P3az2rB8aCTTAEFstJcZYK2sqeGFfgi99/3lgZj0IdbA6zxR3M9PgX
wpU78dCCipjlU7R+Y8dAefsoR/e0UCkgknni0cKp65YPY8JAapyO992JlygE
/HSN+1BtmDu96MYw8YRgcgd1iLFmyWzzH7LTfwdaQTxCX2IzloqpvjYw0l3h
e4zi1iLmYiv3ys1YzrAQnVmfzJaFEbY762Ktole5ztTijarWtNXN8T3X6hpp
Lb4Z523VZ+s4PgEP5gkcyTuutER+4Kd/PXt0j9eO2d9qPgsNnFav46kLkHb4
7x8GYloAGdlVaiUHF2Jypj2GaTkMt1hIjrZl8gb0a8yjpa/E28bHqaargz5T
j7muxinKqF26FAEzRhDkd6X8gRxPaeJKW4S0RVUUuSic7iMRxyHocDDSrJX9
WPv/YjdDm6JWtoDSmClwfe59fr9aRjq9tqi2aS0mYasxZtdPqAkrpFXQ/C6R
WKTWh+C9lT2AQUyR7SBNVjbcNmjxCc7sdNLSffzH12HaSGOAzY6h/lTsd0fC
qB+Llfq2XSHiFTU6JF51ljVy8Viyl/bhc2RHwfkTb155mmdK6hZXJ15WvhlL
QqqXPVrNW4dhJGrxHkddORLhASLJXz3QxCUjH68wSjBPpIkG+z/RJT/oZhQr
VcltBUfv5wAzMcz+eiQrnjWvZzB9gVOfOeOYwbZG6eF8pv8Yh9RQJfk83IhS
mc37PL3QMj4B+hoEa100ADYILpJ2IfuZGjAkVa+V43cs97qNeSJldvZ1EX3o
Z5Ieajs4DORhPDDiqX/pd3NvzDoMq9TdDBSxUPsPZIxj5pya18gdzBCgOhqv
aZJQpzLbVqv/7GFIQWHFYk2uUkaeI/NcwvGaraTCmg+2aHA1b12yEDkZj619
osm66fVmwyTglhtKoNs6BxaIRnjGB+dnpTu1h/+WBRZiJ05oe2P/VE3nZnC2
XDCJcKdkWjMJ+9lAOOKUKJCgfGS0QzLqqBRUQR2xqo0alJo9F0vk2pD5kJad
3zDJ/q63++Gs8jNq6yUBitGl7P/ZcodzaFnf/t2pl+f1Zl7ex29zctVdP8oE
U8klnlNxupu6eQdF8YIuWJ6Ksp/5+lk/2c05NVv8v83YQoT33Ea3kJ6AvOMn
pG8zTuH5ko8xj1dhUh2vC9xuOa+rsgmPTTjRIVsCH3yH+EbZ61LO6VCLeWpD
D/Rhl+8nlDY3Vt1RHH5Qwoolr3mr5JQgi0qBHkic3oSDehL0q4ZBODNiDPy5
nqVVqJmhtEpCxZ52Fybarkf9qqCb0EZFsfW2hvlXvyoZqspgKW+Zu6e/shdJ
Cb+JL7DDNckh2tt/prrlv+lqICXQ5d2XKPKrcmIf+cG+RVukja/IK+0TtOy6
u3dARFnH2jhZuiL4Y4ItOkzcgrex5JDudpb8HTqAcf6EaPlIdawOOsC/vdTR
SwG6f0okisk6pMO/EPyd8g1NR8WBgMIQlXf9Oy+deipF/aVmgkN9UJaKyRDP
JzAp9zr84KB1uCl6S0N//AGaCKuv53ZuySVE6VTgiv59ELMyoWcQcacx7tNU
FyCc11Z4SUmZ1oUstLvKlovNs65OS4GFIHpo0WAh+9wxoOCHD3lmq96kESpT
BQ3H5BlgvURGVOjRCfaT4DoJui5YDRoJx2HOOIx+EyrWZQveyYQsicQ1PRyC
CCRR4MDA9kliza6XfTUpVqaxu7EyqXXZkMzEkutDwZFmnvtrAMJJWJPgAdpS
IIzkFv2e2coM3vTmoqChiZVESNQapNE2iGOqKReRHCBrP1kW8poUJVuAHVyn
Lt/EFwMNUgJ5EsNy8j6nCOWId0ir24lj5idP4moZgxPQvagsI69xWv2RNeDQ
Ucwaf23VT37/gcfGBQykipP1P7jCUBwnMYNAL/jtzlJFPHyeXUYF7c9z3BV5
WR7+MKp/RR1gKI/kAByXEeG5NaDmuPqSCyVKhMiO0IqJgSzWD50ITZ1wcVlS
rojHhHmTanC88b4cx5VK7ImQX9PdpI0bmJsa5vJRQuMvwJI1C1rs5gH4su/t
KkB3jdNe9xuna/aPOHIp5Il8R3jpGJjP5gI7/J2OzburggQWvzBv0L7wUTlM
cqn4ANqNg40aMnBvVYXZI+GKspBNq9c/kyz79ycAUz3xvEvAwULDD73edWFm
QKKHsjFEXnGU731DwWF94T86VGJP8UW+Hu8augee9/BRr40QooPKeXxWB0tF
oFEAXQcrSnkThBpHAWce1cJE3rcKLdBf/F82Xr5aOHyO0KAUXzw8SkdtlK6k
YrTujNOneN9kcxJk4H2pmvnLFXaiqxr+0x60GgvXkpR9EBCzFe0zUkZpnJVA
2F55ST/KIGod5Suy8lzE3K6snJSN5uKYfhAOkmJ9B48lsJYstqs7Ea3/gXpn
Mhu191U5IqOCwYpfBkwIgsFThH7aDk3oDPWnygpyfVUzUw/adUi3LzNbpgaf
pxAVjVBWeLl6A1bf88eoXbQLrYF5rGHVqc5FTpGCEDVprvMHXMhWcwqe6r35
pocfRLb6TWOgPVqnCZCnQ8WUAz+w5P1kIGRkzIz/g0h4G3vmwVPHh6G+Q3f5
/fyLtYi9lXrB8crkzA3zGfkQgfAW9CG6ckvZb9r0swqQ3mkSVNAOmC9+GDeJ
Ih39njxH2nvBrnEpHtDbir7t8wzuqEIPFQdU43pN258fNSPQdH2jV7hpbNAK
Tr/J4guqG8yuwqT1MooAqNmpURarqi7+FnXl/499FEb5Y9vQLMVNyNvP0enA
E6sMmxkIl/fZNhWrM5y5xgnQrtTNHTRhXr+g62UIP/qp5IhXBMKpIKfwP4Bk
cZxNTz8N5d/xli4Shla3ho0w4Pta11KlpT4ss//QRSFK8ih8n5T5ZoXqfAIr
vEDvOqo+KnYUeqizUbixmw53HFQD3nFo0M6j9ZuyNhSzu3cJny9LaPiz8wBD
uni+/402F5TYIBlzEXyIm6D3+y7DOPHMQB8U/km/AvYboCI/Nj6oega9soAb
CiBpiEI9WHduZpitPt6ej+cmSwuMDjWLh/jbfaOvpCtt1jE1VAbZ03w1YFkT
XlPdmJdgRCreQ5ULyXle1r8n4bRUtNRpYqAhKbSgbyMMdPH1rZzoaq7T9nWl
LjVR4FFLs1zTac+jLr+JOscSQpmA1fEoff86HSxGfPI9vV3kFBPDJigbN7iM
rIL/gVsk3uaW2Gz1qIx4SicTnIW0qo3QGogPkf30JMAeoIVLuToz/F8tiEZc
pt3WDlnWM8yf/ANSvHcvwRPU2wKn3eubEDuBArbD9AIYjtajid2Ud+5hTLmI
1C5DMG3YDWarc2Kwzoqx3ch9Hkwv72Z24TKC01yYrGKT/+juNMdJpGEw3r7b
Sis/LkLw3yHsOvDuyiHIIaMQ8HXk0VfSPG4irfXefoao49w4ZEfxQbfS0vdG
eyrSv0gD7jFl8pYStUncMDfwQL8GKx71Eo/cbSucDoFtMOgTU0QIDXxULAZx
mxcInvXuxavveg1ANj+zS51976vHXstY6DrQ7olX+vW2hP23fKByJIQKGtvz
KIhlI7V0jTBy6Xx3f2TcNMdH5dDRNhUG6fI7xeNs9jlCFnZ7CF9AtFyOww0O
FdWkb1SrEESmWVV6xFYErnfgtu7rtz3glmFQL+Y+MwpEkonu4LXzt8zYqmYk
8zPQyQk2nwKb0KxTWk1gDPAzqqIILpV3qVU4FvB4e1hBqX/S8CPhvnfHs0BS
afK39liacj1bCHjEkv2lzfsibGTf2NsiJILxXoiZEAGVygBwYTJd4JUGFn40
AammPYLKfrnHR1pwk4dETuSXIyuyYPxguCxAaolEA+UmYBJE/zc+SrUgZOv6
YGivQ8CvwBcMJXNMw+qyhI6Yo7gAJzlj6O7NID8+LhxhuGyEavx/PyB085PW
jd0QtznP/ds153c+UTHq0Rm/iM3yNr0xSmJqWiUIGPJscir7V3vGyBfyZETp
YS6Dbkj/A3fCTlZVCCoiyGZ/H7kGKA6ylmkpJ9FWKdTgjY8gRT1jHf3+Nebq
G7txezVNzmXozqQ3u8HyGsvgM7kwHHDt3SHbVGjm1VjjqdhdA7LHYPh7OPU8
i3l5kFSCRPETaESzYbhjYQTqLuUY8B7I0n5MPg0rTTVHbARtNyaeHMYMYxzD
sXNQcxOfH37mmDibYk35057QpvwjlidQMrYfX8m9jAQJm1gKEVA7NkpkfgMc
Tk2iWa06qervxrz1REHixZsA8WWIs1Gik27bTbE9XWECw8MJD5+NHIkL5N6q
HNGm260CvQ9CCkeM2bbsH6cW5VsPUYjny3dC/Yxco3RliKE6toOz4uGFD8Dk
GoJ0iAWq+BdIABM0PJAEi6G2MpiIcwdAkKaDivRIhBL0b0QYWWshlvZvtc5J
Bb1N+a/OVNnEHZROG38oHoUi46SWuVFSMHZvlIFuEuNS7dppIQHOQR8axU/K
3pnO6QU9+S4tMCFKmW2xJlaYwWo1ZPzdQW5ZpsBfEDlKMiRbFEqkez1JaV/1
UhDXQVr5yXRmk1MlH9h7s16k8O58kdMIYZffmTPM6HlvSQqCgJVwotJrffL2
ASRfjQRWUWyGTEpA5SLYhw2SnxW72dRSZoRBXCFsQkWpRDVdxabpitqeHJMx
LXdYXixZPCkjBye+tu3EO+ZMz3Hdl7MTpu5a+v9NYSrrHnjJXmRz82CLdDHH
isJxdFoYiLS2+0bvTWPdAM03Um3/js+nVXEkR2bAjk/QqKl2bdsE3eMuNvRt
foPTqSdPteH7wTbivocKPnOo3POU/RLJHfTOdNrLsQYtB6n4+Eo2JmOEOLcd
OYpcKzrr0FYuU+FnIiCRPFjAS09Z2a617liGAFWF3BPsdVx+OfpgdCIa4wWs
uzp9yHujfjgd4xxvQvTQmsDggPJuPIg5lqcfuDA6MYPTx+vX5hKxeEl0gDAJ
//1sWpe/yzdv4kO7FzYgnAgaNt5c9kfgvUyDRPQh5yJATbeiuQhoNFWwgict
MHY7fLM6rE1Ihsh6KdU6LdO/+Q3Abh9+Xg52Nkilt904YiI8a2T8gs/17dxK
MnSaye0fh68THhzMxIf55IwG4IF2MSbdkxNOnO4z5sStLYBJDJHfWgEurMZO
HfCM991hBMJyzRmD01TzyYJmOfI9WeCPUuELNajerSqbkrQXsg2LWQIGLGeS
5JLFUxcWNwWHRNJh8gBVFZ/5Eg2pJHP0kGrbtnWFQRwHUBew7wANkCeQ7a5c
86oALKk3+Jbg6dXMQucnxBYZ/9f4YT7yDfUcWS2gv90LiSZgQsy1WRPa8hGv
EVpIDz0TeD+J4/nBfhpeuvNrb3alwzL5/Gnbb36fHqSCT3Pm8p4nYBQG90Rn
+bLR2sNS4lcc3UcsngPGnqZfmRJ0Zup3OvZQhFOXd1rXm+5W7WGh0wuxbn+P
aiaF+wAvUSovhhTAqG8wUZZCsrGRczjJW2/SC+j78pTqtt8JkRo8aEHpBqzE
pEX1lbV/zp3XDjLOB5LQ7Wq6Z4CmvlYKcXSxMSEVheP6f1kEMUZfPqN7cKO3
VxQpvOO1QlqXjpkNOplj1HvaZBH5cIotJgveUOTRlT6l6TmaCRtGoUm2C7My
5ynOO9q4rcuPPsHsuBdmJ5E38YE+q94dCh8a7NAXMKyxfPkPByT2uWlx7mVw
uK3ER8KxBNG6Av4NM6UI4O1eQEBrMDwabEttknW8LVlXjnA0EIAmZnMiwYi2
Wexa3qSFog0Xq//pSe+XPPCps3WtDtruY+23oWtBltdJbZNlBVQjnkklvz7S
FNWxqcET2PjG7/DSMx6xy/+281ez8uSNvKZpWonVVCMMX2YJd8IGZwbElwsC
KGNCp4pHVZdPRKi3Q1hNIrOm3izFnLjkfd3X4XkamHc2xkAc9ZxvqyFFQHVu
JHd3AGg/RkmTEqiA0Goya4VUoHmcA0YiJpASAjL+i7wOHv2rYCYFv5Zq+0/Z
sN+swxP2mKTKwCl6PWVeSlEm8NdTUVwMiAfjtPqrHgQ4lR9+0P8bmkqP57O+
K77C/XWy4Pr7lUTpeGusWiWPWIJqecSYSyhJU2Un2MPrwR3BEnVfBLY49H4s
rbsdIdaG+7Il/m24k163TXJfHLthIzi1AeVm3sdsD9r9RUr+6GU+pdwNRuzZ
SU+MukXH0HN4MvW6vsnTYdUwPJsFxJur9HjutfM5Wtdm1Q8+PLdGBTe3eT0T
Ktnz5skQg6hG6AKjxcUAoCBtwVHTuv5zbXZyD3tSK//+Qr9yBqqYB8fFrOv9
LkiT2envD+7obln78QoFdGSVajHWeTBnzgGNRwW/LzPfFi5v5jcbc8KWZIRp
hsWMUtIt+Ac2GEhINruvlS95ZkcVsz2aJ8pFYUeZwQ8lVMx603s+vMM65Ut3
BcdmXRb+W5CPEtpog87ib+vUfPDn16J9O5gbV6GNoZ/BGOxBsFOpL4JQU/j7
VeKU0pJDWRr4eOdF05vtJhI6/7QY9ePZ5mtH2oNm8jXlztFSKlv7rKnDabB3
NvNeqcUa1b9zMxhN6/xqXDwKPdTFqzx8v+7SKZb1AKFjNi3qeyFjL62jgaif
tUq1qKj0AGAU0+WlsmwJUHIvXb8qd2gSCtQaGZ0D+wBVMVEF+sWb99DpKRkk
9HOYJYD/r8XmrEa7TfnKr6eug3BGaAUa6uKTwgjnbC2WOFnYc/FTAg9VAc8n
x1jleRHx84q2uYRdzJBNHKb2d/D4lwzi7TAupAbm92hsV+wYOBHohG3fop/q
5LxzbJkP8hw5qvwo5eD6Z99I7QzGIIxmXvBtp7B9540+4Due6PWvKduE7mwi
amxupaLRmC0P1KGj/CPF0BVH9ej/9SdnxLDBG1kH43WfFMVqjQeOF0EyOawT
X6M8g5vbYq+akpTS2roqGQm0JsO8AK9YvAbNn5F5iTth02D7puaKibI1itWo
BWzvBP8/QHolNtGv8I2GDniSfpdQwwHzbWx1eEG6u/RSMOjQgWSXwqhntiHi
3FKdrvPc3UfJG4q/sOUMYRHgtAxjePhWV0pZPb/mK78POEf2FXzr3L+eSYoi
MzamqtbIUpWaAxD7dDjbnhck+H1IZj8BBdpeAa7zSTAasr14J0N8tJmcFBbg
TrbqqxpO+IwwaflrzVGhkmk/d4tlJKnTbQE+jSUmojcyvy3z4Gu0Ym4QsPIy
T0iM1Un4RJx5rWNB8tfaqR9eunhYZJw4g+goKxN0K941Psv+STmq545uTnX7
SX91MUvV5gZcRrsi2agehMiPC1t83ybmahRaz9jra+KTSYgKkiczcv76mMBn
1Yi5R06oI6PKC8mvTw3l+jRLjMWZsxYIXroy+7PZOnviqRLkhH5Y6yDHEYKl
eBh9TRthMywuuTeKPRsFR5OsnMq5kYT75GTREH3aAN++Hhkz7bbW7pkXNF8O
e7hGXUZ+X9/hU2xBpk7r2e5Ryr7ktt9KFfHcQNz+Q8epRdC4SkaR5eYOA2LY
lpyj+UMldXJ5j5XZy+ROBtFAf3YlMR1WsxNE7zyc3HDE55LEgRHtezHSoDS9
fWh1mE/tklQnOBFZJtTRr6XblIE1vCz2YZVnOwBOKPWxPPq3yVm6vayG/h1J
b2DM3RCqzG7IfENp+VzWeJM8p1ApaE2XewckqA3W++6vUMI7MT0IYpOjNQ24
7L4dpSxTn+MOChtJiVtKOrZXWr2PJOSiGsIzwUpesMsP1u8ALj1LmNDYPkTR
zYQw5ICnHAo/mDlFua52M9Jj89V0VcEW2DerqFKkCU97fBf7m8/SG7zHLFUi
ej3L1QQdNf6rUvUS/kFKKb09MfGjFWd2t6ExvpPTVpb9lG5DIWzZyTKd4xiY
H/UwIndi7whohiSKuvbW+SOQ+AneQN6bIQpt46wK1QvdXb8/jZuHnPlIyyCN
F6JfuadiRBizKWDBbZA5Z32XS4l+BpYCE6NurtQQ9DH9kbf08ArahK5WhCuS
4SAVPvznl5og7uRKFJIAJyDj8gIzFKI3Q+yl0WjoG+FIweqbCVgHKLmDGdJQ
tkcH3xTTBt9I5792SdinidQPFX58ahQ8+0mkj/dE8H7/eNT3JCdspQodxbUG
jzOiPLtNv4sECn9f44qTY/kEzJMh5bqYWtzmiJTDBpzomy7DSGueLXNSG3C+
qLSzfBzuEBIWzF3529qs2a7sOlgdlXEWaFAfxQyFnKLon1pfAIlKVU3s+I6a
YsBELS2k7RfzV0xOo0LrdPheFbplQdrYubposEg0/MslGBL9aEsNLLMQSlyC
8mtfsrNaKt85ImKG0brDex9ejLw009lNqPy1LD1mvg3bE4Bc2Z2nzrTwMR8y
9+WMXPfI2JI+G2cTQf+2RqNGXFXOseOGlJg/1i1czZqb7uBTHWDSQ/ddFYB4
rX4pJEDg+kYvJFIsduZOf+Raiog3E9Kl7kuS4+Pq88ZIZ+cdeqaMiiTjdJPQ
nVGPKafO7i3xyzc95GNpHWK8FT/vioA4KnsT6WQ4IQe894KSXBgKaOQ0b+Hm
L5f3BCKzEn+95HwwRMKlB1eczBlVD5PLBEzMhR+06kW6SQko4MVUebc9ESuF
0IWBhnXXhP2+4nk6XM2kU8Mgg37z7Z2FRUJ25/vQket+QFL+xm7RbmtB/gYC
/QGNPTztfSpxrMiE18zrNUTQgV3f6z8ZPkfcSjoZhqMDJyiIW6g++yHC3pPM
lSncEMJ1sExbXdgKcS/Zg+8S7dH5AkAnTfg5WutflGNRmCRuLVFKFG/r3LXx
QazGCg35HrBk/0srdtQ2wkLAlA/XxBKEsphLgJdfaHz7cNCSvG+BsyBpC1V5
BG4thuROwelb17WS2EhGglCRnaxKtLjbWKJBM4z7gqayIoQ3690UExsUNPu0
51M8pnuN9aKIGeEkxx+FcHzvkUX0hiKhqEquN9kU0mgrOResHTsruGCtX7V+
ieZmKVXZhpjRNbnzU1mgSkuAyoRtB687Z6U1nMBlbV/tJqPX5w8mFgrwsP29
Pc95tcDoGHiZsfFTONHSrHINaKbxe+zq0s2XC5EINcuSQ+qavF5u8BK0unAJ
+bRHU9yXYH452FA1Fwjp2U15ruLJVCktViLhHUs064uhApY3U1F1bmXJATUG
G8mSM7vDlVY9nXIw9Luk8s3XupN1mUWtHl8aRbZF6zEuM3ZJszAxcQp9Nwky
uob4Fk7V+4LotbwWm8ghJuK9CMjgnPJmVJ6s6Fm8qS2Ml6c0wRiqMrlS8NPr
3xa7d7xwE6mz/vYArRebkH+Bw5PcFGo/uVB4Qgs+AATshDDIqqr5bajEHA6g
RSDYcCySXkJWOYqX07zmki3juc2GXJzx743IiA8FOBTdMcMSnYAK3VTkSQlI
wuCHjoBGysYkGSnqBe9SFHqGF/QldNnIJxKpqmn4E1O8XcZHfthnWzoV9yk1
f7RvCWpmgktcbN67BKC7mAvvhfHgQL3jBLDw4OXBB86fMIm4HqnBX6yh18M5
AFoyP4R4vF2MsgJv2f/rg5TEdNYkvohmTFOOkRYFvXSHzGRxpw595tvll8Ir
wS/Wcs3TSDNpeywCnGH23QBk58mKw6D8QcVuqA3i68pL+luZT5dYMvbRzXHr
a1DRgwpLt4TwQuP4lISK30mFUm7hLQv3cmc/ZZ3454GvWtJmCPdwX1dazLef
ls0bHCNxpMa/JJ/iAHr9GnE+4JrWJgHB7Q2Jm4t29EVVWGNNgydK9qa0Y3Ww
AM22XRi/FpiUNiSSOj+0HYygLYDW8ytcWV0CB9JCQGFNTczxkxyxKTORAZtC
PlHLfy3CYXvungGnD2j/jGfpPOxlCDRdg+LPQxbhq2OcLbdT2bQorH7zPkzE
DnI0BGZOUjba7z3BAFh0tBRzkfwqYhL26lRD51dQawxw0lmgAJSmtWPXSft5
5lXitDdRZZlAEG2PKma6PSgSRop76dlaqViadynoM9cPHyxMpdCI7505ztVy
zdT/ZMmYoP2OiaCTs646fRn+vADUrgp6z7RwYa0W2vMwb13JyWSIhQoZSgkV
V+eP2m1t8hja8nW4wJ6ePcnzjoW45yPXT9oJtKc1GCOx29kVCPTYRwlZjzuc
YPenO/lkGcgkOwztDUO75jDj7bCclkz47afiBmwD72vKt86fqeE7w6op+Eup
FEQM1ASDRSr04giEyZv3gjQbqa4Y1DBnYIyVrqryPb8VVXX4F0Hu6E/r4yJ2
VsC/2CMkgmYHMfC/COmDbdK2RDGg7sa9omStweIUhm+CzvIVl26JCzstG3Iz
IFd72bO3TXSpi5paIjPBG5uE7iR3ik0FhrYwTW34Z6r/UrIow99JMvT7q8gx
rHQXGUk3hCr7ThfLaItWCFXOf/luWnlbDaOyQNiKS16YhVpznQGT2/j0d7IJ
K18aCRabGf5oYG2vW3f9hyswe7EGxMxSglPHvuk5anm2TBqeqpUScvey+aH4
+DxTzEVB5mIkzDF/NQWmTUAFXP6p4wk+iE84WnXuJzqg9JEOT60E36iU9Oqq
QgBgk3ylWQttzr3FjQEVyqU7kFmH5s8/pHXN43MXi5WT5nBD9ZV5jtzaiLk2
a25vI6OKtmJK/mSuTTQtOqA/Fcxyqa7Hpu0zjlSUcb0cgl9Y290m4yR/TI1q
i2ENF5ol/J8fwt0sbOcv5REiS735nby+1GrxP838DoKilsrARzM4KkP5pWRp
OUWx2Ex/35Xg1UlEga4wmqM/ZJXBMpRUY9py6ljGa/wHqa6OCCfDm1NFNvon
w+9Ix0uZ1FXRGHdeqmbHK9n9HNSJ37Niel/BbC8PaSUYj9FvwTmRwLWpQpuT
iW9v89sI1y/r5hMT/85ORop8G4uKYsm/xy1/afaV7YNqHbLlFPC7oCCRM8lA
Ibs4KKpw+eNVf+c1SEj2P6ycSOPXZynFlWsOCxip29T+0soASmjp9x9aAJnG
rLscJEqKiU6pDJjCe+yqAOFffOJqnfqfA2mOJML91R7pbUuM6OOF+8U6bM7Q
wg5siFL+bPrJ/XVLo5RAA6kL/PWODciPMsaCH357kjiAnfuibo44RBW9RKHS
oBx/2SHsEbPTK3wzy73ZOpc/AtviI/wZ/hybasLhnfU58F7cSgJH6/kT/+sK
n2DiFX8xd99kEsB0PDag0YkfHgDz1VKZwgFetxP4W4cDJ2RkkR7wRSR6Bdba
2vrAw1F4XVvqWakwfzksZsoaneRi2CGcCQoVKbzFVn5jR6sl/j431c+1B+m7
S6PgcHrOImOPG7eiZ76+MC0vCqxNrZqcrVx3iiXzXaR94fmAhCXmwiBcuUc2
YWQpqpTqRH3H2tJL6KEqZzGzLp6xwjCHBHjrzslGIIbxSsdevgHDOP8O2AYi
eUKS+R2eI1WIZbadfSQaQYHSNdoUrvj+BQGckEt/2Jj+tSxleMhWy8xApr5Y
V6zfYx+BkQRh+Q+1a9oY3j6I1IKkA+fWOxkxvJyeQ0q6Ac9/vFKCcjUtHpOr
PZjlrDpKD/Z+O5stpj+o7786Exh5zzUuoCt5Yl0fe26z3Z/T/cLrF3tZDPWd
qvlqA73q3VDKk0SayBHmKAzPTr5q0Ko8F2V47LpFyzuey0mWr9RQAHyG13jq
t0b2qEJptoJXyKgfFh4kI/j45/i5PPJX9MofdbiANLT62PwmjL81+j/d1jwq
z9QAKuqvQNRAIZMKu8+zZeIvol1I4aJ0GszWpzi/Qrc0dUip5fCBpXYTPUAh
CJPMXI4mXAU04knH37ErThp+DBli0EAI9NEF2tohChvj9d+eNzSl8AKMRuJp
2CYsGr+J6QmC8LffwBHfnsvGgoorrApVPFwHPlNwBdr1V96DCAJLv7DouVLe
U1s+wVPQyDzBj5xgMklG5Yb2Tb9XYxEG4SUAp3Ep5mmZYfbUOQ0QbjztsDM0
jaw1ffL5KoXIWIMGYbHXFGWnisb6L9fHqGinCZvlgDYjuxclOQ1hE2A1Z+lx
p1B9d0vdFT+V0z+o44ROzafOuevR2/cMZXR/6exD0QOLqsBsHGJDTbyMtVXL
djS9p43qUZyWJ9C3VOylsMymjrAskE2ndkObv88FtO/vtWOYby5psvwYOt36
BJCxHYVbQe/idVNT1AnPGO92ao5SSVjoNdoZywnZbc3OptDmDVofPGIZVKhg
hkBn+0+oJmYPXNMLYJGG515J7bw6nsRrlnIeHbSHAgOh29ZpZ0KEVX3cs4Kf
O/Vlg6xZQcJm8cYTUdty3M11a6L/hiKIFMyGioT1zLGfVPMf4uOR7oJimHfj
Cp9ut706UVJxlxVYLyWiloW2B80zYP92akp74R9HGGLXA9VJ8daiZihvFliN
BmsjmpG1w6Lbr5M8GZ/4XKJmKF/60niltaAkThw0ioRU09JWb+J6Q9fWZdib
mMZFV8q7YzyEo5rIEGAjX3lVIdDS79/x0lCqJvdfObaoRJvp13Cf2lMJ6GlA
nGeiQ4khf1ycZGm4SLbEdmfgDN6+UiYQQJBx/46fuBHoMCCIvgeOjElwXiCU
W8bt+nlFmEmQanMee1dSMhZJgFqrCpBhpQ/RyO/Ecq5k/SpReG7In/Acrkwh
ElQ7iX0oCq4/Ejr6tEg64sxUDK1ecUsNVWKHDF0XzFq1pYFIfoRKYAZaqQyF
kEzw7kL8UhITXMF5oFzQeCYmjASxvksrXG0rZFHiTCygGYjOcw1bbr6cqQpA
LJZBn7IhzNCuRYGifu41LsAC+LXVoKWlmMEtz7UvzQ5RvXsE7BLWrJgEyT5e
uaC18WZhCjmt5QHAg+IoskiL+q5pps0HV9aDiXKlHN6MT/25m6Fa/ZDOXk3L
g8xNtMjniSsAgeKT0VoKO2PAJ34Jr02nq2zMJKAcZPWBUAtHrmf6XQSVze8V
TU94SRGH+hp67VJpXKQFvQ3uthIvWt3kNE73m8xRk2NcHwtO/IAA6o7YOYYF
9gBcv/OGePiReokLdyovIPnzbE+zH5FujCa7K6lR/DACacJK8pvUUVFUEubl
4pgmJmrVjvnSQ9gS4HmlQEHdXWgWAUV0mXeKpyDAvd8LHtJWOPj9lHbZVgBK
fpQxq8rSbFNcfwV3jwkj+J84bHWUeLDe1FsrzAZCiC+240/1QdUiRWMXJHsb
Uw3IoDs84WEULdZw8rD9pgXuv378ax+Bt/2DlWiOj+fEjeNYtrstmA9GVJSv
FGtCF1n8AZWrwccDPZR+2gbgV4tKFF+2e+LFrSGoVOQDAGzMimFCJTXBIxJl
dm186/w1XjUerIZpIyVltEmCe9wi+ZoBYkUFlOFNgGHV5489njwsPa/drFit
CzAPPkLjiuP2edp/TKwhp9QkHmX9yDE5Ejk6zBQZlpbA5358mHLNESNaVdxZ
T8GsSw9K6S0Y93NG8qL7m0JIm7naEfcpiWElXU2snlUsJBBd+RwAzmd9I/yT
kSCexPvU5UkQ5j6KgfMU0GV8uz9dHqHIKDq7ptXwzjiOIrfmz57SOYmi3CFt
tQDUbkKda4lLSIZfOubj3TMutsnXQ4fHn6EM5hf+PSl3/w3z8Jrs4AVWUGAC
hM2cNuS5exshB29risKXosg/JnTlBBt0j6NK/H9c3hDrfpoxcOyAyMlpYrGU
dkf5rz/K3juP+wQ8STg7kkbavyn/sZHltZ9Nmk9c/iaXlYGOPQKNUHMB1+48
9GJP1gKCym2ZJV3pmHrVgojhJju9FQga9oUbAbSMoUKSRM0wzUoQ8msZSWq5
Ojq7/DZZxD1m+/fexNH7oO3zMWIfg2MILhztwT6Lpwn9+S1oOmiJYuK6lDI/
mQGdCeU9dAnqj2dM95nZ9jeWgcKtFr4jL/B1c3IWhyYoRzwirV8Vh4lumRVX
BRVoEEzyh49qrTMqD27DG8uWQmzkm98AMVMlzrQHaUDpDbeIMSXhFodEDq1c
KNqQJVDf3p0m8H/6hfhyzYtrygvzuIzYtECkcwbDM8ezK3coIqLNLej4CGiZ
DWTJy58o7W/TdER5CS7ejW8VW8AgictNRVoOKD+jTVZhb1gA9i4gtPKSU8rZ
IEkLm7gUeQe132s0qKB8GmLQ9q63NQJeee6hUpkpyTHM0cMb7bOfvQzjXUER
jHJ5gEI/LXaKWgJhp0yTKfXYiaI18qzAxyt5tl162nqS0jcDIn38Um9B3id/
7YCgsCxJ85TZ4Re9VQbSgV4c/y93lfgxbL9YEdbyIMzvxWf+xxwpPHy7ov+t
mg7lOKAECyvtIoWyONc80D/dlWrhKWZlEUl2YxQJuvAG4Vo1oyigzUM8bjow
lLMnrJJEMDU0s6j2VMSSYj3VPRiP7vy9xBhrbeJC2GFj2CR16L38SfKy0vMt
zb1aFnpTG56SOiqXVR5PP8eCKxKlsrfvrmTWT4yZHwqIC2Y3VNzzyk3OHXGJ
fO/92ejDyMCcXjoZb2w7WJSJiqPoufnp+yI9OGqqNT+CFP9llquhG+pgyDTR
jvSqldBpQfQF3eYC7QFQZgn9Rn7aWDp4w5a/abNpEG0EAXR30v2aJTjSPfMi
pwyjH7fUBf1+3duzoT8AQ+DTyccDSiEXm6paS66o18KEoo4ikFXiafsPaG1r
/hz+kdXiEBhy2kXM3damDhQNmGc3BDcUDfd0VFeGyZriN+ZX0ta5d6QG9xPc
5WvXSqp3Dg/IQIKrcwFPqrG4dtn76uNhWy/+GIx+zuV9g6FQnLV36Z0Bkn8d
JlZ/5NlX0BC0atudcwwHwaMKi/HD2MCzU9JwxP5Xqw0mGEM7hvVseFtDTwcN
GXPUgsQCLrRG8SHWxDHoSNpCSRDlZzGYicnNFA0HExtCOf289uNPR6wHP9UO
1FkN45cvMgjw4ceE0fXB59Y6UNoF3ERk6w04wvyRTSE2wMA8oXOUtLc7X3+L
eyqRy0HbDdeUOXL++6sFjRAEfnz69Z3cNlR0fEY+iMGNHY42G4d+VOiLuLav
XfnqC3RA92WxHSHuWERGkj9QZjqUuRUOgQ3qnfJRkMAQi5vJO8WH7rXdH21Y
wXfX6bRpMOqD5aF0PRu5Q0l1mG4QVRHkOsWT602YL8/6wa0b901cAPQiFyjW
8D7cj1RyXriCxCAubZExoa/FtgZraSY9kz6XURhyt896ZUIlM81jNDJqph8X
osPfhXCgoEN/cuurJ09v42kgrsCOj6gpi/O2B5OSIettC6vtX4uJjE0FfvSZ
Qu7Xg2VsKkcFcwVq863agrR6XWV/Keiuu73ljLwJnUhZhgKls3FXAYc4MVG4
gC4nVP4opAzchwpf/IRo4fnuXIa80u1C60dal6cjrh8XiwwKQDM8ULeYRkfo
73gCKPCy3Nh48Ze8gCSA3x0khcRg8V7VqoUo9uXy4/Cooi5e7qEloTqoomgv
5oK2jVkqWYAk4bTgWbJhJ+I5/iZIshxKbTTwbPQ+2/qq1IkWqRp4y0MrjwO0
eeQ/aQodn7ij5gkz6twsiFuTc4m0X95ITS9gAx55S+PEhMBe//jH4fffBXVF
7Sgmj2rx004oj/nWSxbxGagdJx7Ey3WJPgzSwyTVifllU1vBBifrjdj/7HA4
7D4cvYbFsSLZVVasQqNshsut/EaW1uN0K6Pewp67YB4ihIvusMxedSUEVHbN
SMvN9mbTaORpZE26PpaU3V05fsabiVkLIRKn/JrK883DAIlAf1khzo5lgQFz
GSHp0BDP7zPbgCvQomIYw/rwWedcsL54lyaEjx4DHeqOA/3Iq8HJmpXLdOPN
FMEycRk/sqoMDBwk4dJs/CB8kGyvla5V0hPSlosAGD2litbsbcHC1oEvzGbq
niM59bYZJ7vPlO/GbWAlwz1GKVnCtPf5sGxP7to9CLNkIUqnomJTe1umPzFd
yFEdv7equDycYEhrGRns+iCRpe8qW2ReconsKI1PlwcI+LPnIDwdO2lZ1Auy
xkGQH/OoJU6Puxp20JQya8SyH/q5cVQyxgnavueNqZR+yKcs4iHK0Z3FvkdV
3/AEtMnW4NAdY4X5Aj0UyTr1Ok0ep1LJW8KnLME179ft/hS/YvZetiSL2r5l
+jJV+cj4julyftYDVxnWl6LNSoQIIenExaD9Y4wGDBpiJ+BWMYP7nvJAX7Jz
uwwMfh/l+jM7xrKbM18sWSZECIXHQhRn6jDWy0GZmzn+aTBQ/52Q3pPbuvvs
/T9DzYhCaTbQBYjjo4XBr7p1NDdYZ16SmffvlnvPhVSYiXvEY83M0f082XIl
IyKIvVZXQHSl/WvSjEwrPmGV6+r6blVC6QCcAzV/OstMrI5zzoPoxnPRyZTJ
jbXUzlS+EuM2BDbnKdDo0juE+/SNWkvkUaOlU3OqPbt2XbWLfBTwL5dJzfGD
iwrKq2lDmxYlsPSg6bkE/x+i3FybO0Sa+CPo4uiYFrBK+vt77QN/WA7vsJ30
yWNOpIt0fvhRYApihQosakzoLBuwFuUe+WBqp8N+QxYLEEWiVqG4hf/u7xra
5jlipX3ZGzF7izSL/dywY0oM0n5NkDQTioVoSvivqUFCz0Yu2qG4C+ImQsqk
7CdwzSLlWeJupS3d/eg+f9beBlYhfKcKakzb67VM/XhnBElU4beiYNsA6lmd
ES8S0xfiOR/NEDr29+5C0HnsbBika72Wl1s85/NEhCiXEliR8oevnShGFK1E
L1A9CAAFlKn+SMEq4rtp1C3P82Pau5wVrDtnbUp/D5kUymOFAdOJ/OOGGfvl
jIe7SKxSid5eKPTNtCZ8PfiX8axdPM+QcYZ0/kru/OXGrZs72pG0lSNh2ePZ
m9a4tLzIpERXjFMxyTEw8IEmHRI16svoxiGuWeox4qMusrzF+Rv7tM+bw/Ie
hzYJqsbfXrBw5uSEQMvLrLiA3smog2BanpRf9Rq/V41vzDZqLHT6b/6Klj4Y
cjwLkfVyUJ6I4uHaG3H74C9L9PIHyu2djEVHfj9rfUjRQ0eYz/08m/ik2SK5
V4YyuA2freitBp3gK9y3Z+cZyV5Sg55lQ7PKkx7ZwaOOmh06D0xsuZ34Q/uA
bA3FnMPLQYf1vKC0h9OJb12k/rMx40CDbXRYSP5b9yX67xS5APBrJfrVk2IO
yoFjr+iAB9sRus3PuRVXcpLFhSMEFu8+wy7WoEkR7cau3oUQdW6CVFq3FgSr
MAFwKt3Mt83j/cM21dtcDYX+/z8QxQtkqj+LPlHQ4mha0FBRQQF/3DeCOxuH
vM9GEqCRSYVKEc97gT6JisNeM+HOF6IZhhbl85ULIsr8c1kBIRZ6wRXwfuKo
vD+0eUuIOkYW6G6M5THMiXAh9iyxLmHk6zOquy5UDfQ54Idz0Zv80Q2adU8S
sEFaXe8P++AV78AHPKPyAwNYxQJNWTL0pCR/4QdpSVL/c0d0AlucdDIMpLVU
BIaAtS4wDpc332NdHam4fklswo4vpJNcvpQOeyIgksLK2fw9lNlEeG6Ii7DD
ApVxFam89I4MbG4PZGtee4Jtlz0bgQKjUrVPIgrwd1es8iOP4VyUOxNqjKD1
70B0h9UXaKA1s3M2RqzSFyjLGVT5ljLnTxuiBAs+WlGxjfy1IErg7ZFPHV8E
thobnIt2aBn9hISi10SLM7pGPKFkjuJy2VlMGnu8iT3GOpHoi9hCYegiDe95
l/nDCIAG1dZs0lfKjdZxquk5H91fp04XdnLFLZqHdx5beAVzIRM+gsJhLg+c
g09siZWKMmsLU5MSqr9pbPjGQNgtJqejnRINPQ1ufOP77Lbk85NV33K4x+y0
tNuB5j9Rkw1c5BpesnTQJ4ASxmXv5XgFfFEASZ4yfQWMK2rS5h8QUw4hIHq8
0AUdOKCs7l8J+SfC8nvRLayNltzFaVBFpNiuNXTsRzAiMSfghGv4P/2XXYuv
+kY3U6L02PW6xj9FcTKdTVIWrGVEh+LkXNl1q8x1BEBvUrV6gRA02/hMPLl3
47o6VUVkfLjkjPfvLWvyzKy4ZZKZu2T7nFchl5XyfYNkUmgLOK6cMwAjpkcO
x3D77ijev2xztuenQz8SPJBNWYgJG9ko9NsOllrzSgqeozoL8DfTd81OM54I
nj8a+DTKQOReuux5Tru0lyTY2sY3xjSd2J3WX5WqmXPRfHPLUanlkE+EgJwk
IO3u9g1tbd+1NLHVa23vdQBHQXwOvLEpZCSFy6PT5m/Fq7epp25BBD8wCPKt
lAnMNLzuyU8sZuMfVun9ylulFvEVOofXDea7b1tvLwIR3hj1Ayb8rtJmINgC
ZUBgFGcsrYdO12G9zQNft5npeYOUsf/hbpSOA/qCGOW40vjX5AV+3Q8shU3x
qUIP4ew8H0ND34qmHQIDmZB4RWeB1MCfA7inatuDOyVWIluFf+ebexsauX1c
+28bzzaAqnOz72wns8FakwyTqFVASFMO0XyIDijXc5KcMLGzwt1rik4qFPvz
nKsTcaMc5FJ0bd8Ci8nyciT4x5aaPHGaE9JN0VwVQrB9BGciERdjWqJuCKy+
+qaaKQ2n6mpM033C0qHbYRzIkOvrZsCI0Qp4zFFBEwcN4J+2S+LhjT3Mhklz
5ohlvcVYLMLyqShpp3cuta+dfREYqUAjKCd79eP3S/gdZg58DwIYnIxM2xXs
KmZC56Kqu4PaXynYCAkToUam75XCwGOX2UMsEPS2cJJQ3fwfcRWaFv7KhqN+
GOvxLsWSE8jUqFsyuoMNbfyREw1MGITSe4eXZ5iIX3x+NyQ6yHaagfF/gIXF
DOHFEq+RybM4eXaLw6xC0WI0fpeqDze1jqRaKKp4j0r87fNRAD5bFZvfgDqr
+1227h5dNYqOnhn6DlFtjW0DaPBRfrEYBt/bjVBdlKQpZDKodlfT2lKLSuvF
X1+yc1ECQVllZKlr5G6NrIBn0nN6NUTUL6eMXBOKeXZ1EoJCC/p3naLce4Qk
xE98wNzPEQ6WVny4fSOSH70MoPAk0vmFx8fzmHJZHdJbMewSY1lcYs5DrXUA
Wc0z4bWJjeeBAypyKTUIahf1E7BDwHg7KbVfbX3RvRgneKnXvAyrUdmXMUsX
0A3GvHSTgdGcJ1jZPWzlJtuqf2Zzv5KO9AvGKVSo3JKy2jlX5GoNE0dvA/c+
s6BUHiCqi1fES9QQWylaje6/fg0p5OYcVFjHt+p8224cMm5TtnU7Ri2Kiblc
S5Eqp+o8KCn/iCp+F3NIL8HVn7o/NdniqiRwxFP/RopsBj9B7kNraRAeQi/t
ljtpamTIwBZQ6Lzu0xtYr9r3c3pRdkYpUDI41ZhzKTSTIGTBt1vyc0wXK3Jl
pCZVGd/zRSvUOV4sZYR0+MQVdHUfNQ/r/xuCTBlXjb2QrwBpCcLqAmDmry/G
XNqozOqfOMlq1XM9BxiIUmeSX/Vdpa+CtphJffIDgFlk6eFICXdWF3U4kEkp
WJnpPXNi568+TLYiCoQlca4cq22gS7KVtPsjX8OelvMgQAiY44RsFjk8Jde3
6Ciq88StNOFUhFEETI0BWVz8qn5h9AhgXMmE1Q/Kdke/rtfAJFVYfeNJ4qme
Y2xxTy6AofiLiAUSecDDLaGh93P/iQGfZt+lQb6vX6BK7kV5Zlv4yDsRQY41
3bWJ7Kft3rvFxZijMUxe6v7sffOnppUny6PCgS8RuHpoif/lj+Thhm04Uxa3
HMrqgTLaANd8ewUloTRLJFA+XKX7343G1wWqJJh6KQLmpDni6/Rowh1HQqUB
XOoSH0nWuQcAWK/j6g7XtKfRcUvxgL3SUgMsC52QY2Zv4YZfKWCtTQ8FopAu
rkFl+i22CoBrkbowD36S4XaDxGyyL+Foz4d3+d7OrWX2UT0YMKAACOHFkHVj
X5qQ/TGch/+71UmM0VnqahczrPanKkg+Tq6qrrZvJ1sMbxmpxiEFPBXgryFL
swhSWp8PD71+kmF5Iy6UGXd9vHA12uh9pjan7H49mQE3+CjVNcVMIwUF1lLI
ARmqog36LMUBovAIiDVNYloTScw4VzV3VCchKrH9fVI7xf6DfcIERRVBFSP2
0MRQNHuNv/N0goAybwTevca+aw1xUDoxJJsxRTm8eV7l9QQWH86ziVFVhDL6
6HjhxxM/sWmjwtNerFgm87a62qvJbofFKXT+YdvQknU1ftphb67IzSLXH6oI
iwlXyjZVKusv7k37OLLifr+9OoHmzRf2LUDJS/JoA2K006z0NL/fduMR5aPt
0YfGjzjuXbxrZDiwxsK3Yhosyt8Kr/FpuClzdQsGhlPbHgVfV2GT/jB+Ivlm
sUDcdlao0WkDpJnTrM3G9MhkJnbM4RakkMiM/BggywFiIVzJBNT9Q4cvC/Ax
KyyzbiYmvR/3CNLW2Xu2UW2dqJmdKW5D2dDEfwKyzlDVGtGPbBJFXwD+y6ro
vwV7cfrp5h3akfKubOvVGJa8g9Ar+yl8D4ftK6phR+i+qq1g6ckXD6e5NBli
Nmp72mUj+vSs9nr6DBHSTh90VBJRTh0I9j5TxmPlg6vMlhJnrW3mJfbMmYVr
uPNJufOFwEIZLK0sqH8AIlvzbGzDv2hguyYwfrp+1Ln6tlqIRs01eGQUdM9J
LC1QrW3DKhuBRFDIJhGvcP4iUwLKbCsfcynY3T2SFnxT03qHYn4yoKv3yBJm
EoaSqlC/Va7Mj70ac+znnUT8yFKqRRFhuOFkYvDes30SUEOcV/KeKyCAJpmi
VvzuCNqQzWpq22U0X4hhc4KaTV3sumFQYGiAM2XzPFNMh5Mrs+HVwQcnf0bD
6Cz6OcZoBxsvc6nx69EEttrB2YZJKey6rxEZLp8oO+FPIhTpnZrSFVTSe4PN
y+eLQYCI1r/ogJ/bgRuqYL0gSYq96+BZlPN7aGuaLRmGQEdRxobUnyEn7C3g
rca+yigNNBDOteoAKSNqFTTRNlHEXuZdMJKuUjya+CsMuney4wOp7NDUxG7Y
CK4v1QxAiMyJ+AOzTcgrgb/vSEzjOijvIa9djD3B1uhFcUTtFsQYgeCSCwvS
qZU4GzFtUdwFPwzGI1p95M5LkkE9B6LB2oKO32H96i8NdWpeFFPUY7+MapM+
Vz5m3EWXOZqZHN4Z2wwOrDHzoWxDbi7eFM1eddGCRRjQXzjX3XTtc4au6icE
+gmwnT+QdQkLR/RHlj8W9XJiSkKnXHxU8Hvaqw3Z5Z3aZRcj42oW4d6hmqSK
SP2QGxRCau3RFyhCxey4DvA42HfPx4g2vr9JQmStroJcSSeMAobI0BUCLr4D
1n1P8bhxculmgaqnyaSyoM1hk1AwKAERhWHcN3AQ7G9wzjhtRN6Y3mzr8zKs
/574XkM+cJaxdq/0GNkd7BTvCCI1s1ZDwvs59d+pWTqnGWIMrzJ/JowFDXbx
fyp12Hv0dFMsNpFesHVaRGhtRXUFfyr9WzzqERL2plMoAK9ME85Hvmfe+COY
scY8r3sv6mk3uD7yJE8ZkpRa2bbmUVOnodpp3P0mNKzQ3ZLCpqu9XVc/g+QR
gvlTmHfmD0HjLxaBv3jY2PfRwG8GTwgefrYivg6sDz/+Py1Jwjw0+f4whIbn
BKJ/aduPgS/tPEQdVYPTxi1p0UwDl6BfsuwZSkVBSWAmk6w/IqaIgfHaRASU
4o/nKlFQjQ0xU/F4XTvbpFPvnBmSf+CQBP7BU6CPKdwmAZXhChbMoTxq9Cgs
DBoAfNuXcfhhaiO5RuJK6z5+UgYLWC4kBm4YdbUqKNihXVVHsPDXk7Vi/pi/
DtRLnVLeIpOI+Ef8khnfClYROLZqF5HtmEQdNT/9pqRjpERwBAQO9dzWHuWp
dxewnDm6CV5KXmZ2pRgOmfjLqwK6tSSBFa12s85Fuk+qQvyrpdsUNHzjMkSv
BcAzP2GUZES5HH91rzOr+qcuktwT/Fq4lUjm7X0d6OI7+0roIJV4/+nJ/4v2
nEXrNpDqMGU0HZKaeRIFN1TvN1pTDqbhXpGiyW6yJK2ON+oCbNEI+TOmuFau
+fJGY+r+LCivNqoJabKHaBntFWYl1ulQyjdMP6CnORPIqyPirey5BUp5aVTu
4uLCfV1yNUJJD0VRxgpYqmGne8rxvPfrTEaU0XnIcMH4JQpyCwuPSo5deNO9
QmbDKTQiha71y3dKT/KJExWJDmUlDFYTP1on3M7gP0oECdxJR6dubtubXB4h
unc4RVWCYNT5FjxZXUYHtYUqS9wQjc2x2F8yrWlNI+4oRvdSKI3mamDMR4wf
XpXHL9+0MG4GJwnGHHQDU0Z2kG32dTl6uWGkVyJYdeIxqx3n0tcL5wFa241G
pZTe73AfyDJP3wdxicFjRNMNvOtPHmTn/LVsHgkno6Wpa2EOebt/wen/wfZP
b2unmwnmZeg6Kdtz0s3VPQkWHhdQq2CaAONnRP6CgmL8TmhsmfEKs8Gkd6Bj
WOOqLs2AN3hKtFQ59GKLSWd2dJSmDLGfpogwAb6xqCOJcndAvu2YyqF+psks
e5db7nxKR3fO/nOaIlfVbzWlz4MDW05rwmjqBaHnidvUL5Pc5SiiNEKjm/Cc
CkfLejd0p/TM4u3WsVrKq+zpfocuANomig4li5UMiSZ8y5gde2K2ZHPZWeAy
y4xEHcrwJXLokScS4OtyTPeJfQ85S0jEbKZe9feI/S2eotYWO8thvi61Kesz
hW2LSrhbPscPIOPIUanBQxHYNISuNfG0551Locd9DNrgm4LOW9eAfCrTJYgI
R9kvPs4NjyTyfX/PrAgb4u5NspUzydCbTQFCBDKKE4ebQ8sr7g3RH/KJNQPX
5be1wE4+nZ94oTNryapwM7EoHUkGb6xaiVI5jD1ga+V0clG3kdQ0CwMfRiEQ
Vn2TQhHfv8yeoG/7y3LnsQGO4EcfM0n9iXaZahm39dwGu8jOqfKRqPbK43Gw
x04jOmf9TDmysRXPdOahHXsfFHMFaVi0g8itN0OMdUSTBiqtuMtEEQ051Fpc
ffMougsB8PhD0MFPCs1WX4T29JZYri9EEdXgcU3Zcse5efPJBIu8rcwf7kc1
Mkwl5ejClg7kEV/03m1dnSMJw5i1h0R4Hz9zDTMQZF/l90o/nZXnCiV+uBq8
WrcZaehyqMbfrcQBOX5dDQiL5bDkLUbX7/pTm2AKwRZ05bstl4WvDSMTokWe
ylEF4209cyYncUwukEYV9EkHwqPa6WgUzGMAZr8t8apOvc3QKX4K8S6My83d
cfq47VJO6Bp+fwbHjqD198c7m3zCj66V0va2AK/9Oiu+IiPL24ycFPkIyVEm
JhQrEq+QcvFt7nnYRy4aeWYxqljxUU6L9+lOmfT1h4YM3G4/wQkz+8yONjXz
ffKxFLoWdYhPgEPfxS25ZM1RTgNj1WUOvVupyjvxD4qmJYHQ7Yp/VfQVsWaW
IWAlQvexIV1X/SSqTgm2usMYlWdlOf3OccZ7euP56WkcvlHft70YM7kvwbXd
eEnGyGpKgDfA5pOF0YWgssiTffB1rpbtT94yEqMKGHUKbR7SkG8Ccv82G61m
HgUBggpnvHKXvSfO70F9yXOX7WFdGMz8ptZlwWtNyWLyd3DmEs1WGaG6gb6T
VOgQk0CjVRm/12MDQroi+VDU2TzOcZoYao4r8UZNe2nyfmHDMCeIx0nxaVVq
0OQ+qTNH5+BvEBBNwGJ5e3r4Y/paRwAtPvUbM8IcvRY+Wcm5yZPSUdfcPm+B
I2KqbDoCY2sIsPfO9iAUxT5Jk2glmINIF4N9LD1OuR9EaDOSlFdJQLLbJ01M
VEko9t66JyG03/BLGS0TJxDmM9Gc49aF06lWHqOSpHHKjBiPgzgzgfVrYTcR
J+0h5nYSCl/eB1PIK8KtLehsmxMGrtuyEcIOhenN8FbKwywdPS0AEgBNekIp
tI9BrHMdrCPgu79AIFwPuIwf/p/PuGrAjDGqmvN9ijqx+DVLw+aaUZc3L8iF
WcmLHfIHFGQN4+rJ/qiXr+h5pwXXWEftxYyose1TfS2/imyGqrdOG4GZ8Fhq
iH62AbTgR09R9KoBsV/SKXwE37WmbQFMiH+FvFAvpgLB2bCzioMpUM33i5zR
RoHXKkYdah5SP049kq+mAVYgmhKQMnGARudgj5GcFb5USPXpgqgJHgm+jmnr
Mfy3aq7twR/TGOIPSa0b+jz6bv8DuNeBlwUSYpnjhab08GC9GOMPIYMvpTH2
ayh0SxjcvMlQCMovm9R280jD69InBXQuoTvURFPidDluoUj7+dofJWYEWf2T
dJodIKI+YKdWftZFQtfZM/yecCdGM3kwkfOYijOq3xfDXHKrvqkNN+NpNT4d
j/QSUrsyCEksl1tKHcWfLHdXZGw0ECjVg8f0X+ybsdcBh7qyNiq/m0GrpaT1
MWwIL9b78aSlYSkS/y0WsuZz6IzVF35fvQSXPpCZBKquFpiJG/nmRWuG7MwU
nHXjhIjiyHOCfW9z+8tkp2yC9JbEuPjgpbRDc4em0OlDILSCCyhkYB8YL7SB
oLIksXUtofp5cgClod5CmHE2eK//rua2KvlbojIyRgGCliAvy4Xdy8DyKtdF
2Rd4McT6QnZoxxr4qYYF54dwGrPRDZvDoAzinxBWy09anGglchss+Qc61mB3
N7BVNse20F5Of6fKdex+XHAfZxUu7Pf4F/NEbPwa7J7AkxS4wEGprOyUVijT
2ept3EJchT66IF1Yf1gTc1HjJFENIljcv8XX7joWvqObSL1TV4zBzLOvabcR
At9mj95JcxG/VEZcpwmhYaXPQJzC+VdHS3sgAQdh0iVidrx55q+uqr6bipNI
apZ9gBV81ZQKCKMuv4K6xFXMtK0a9MLxHABldc46IKvrsWGjMVe7IeQjieoT
p1+CbRwVDpen2WeU/rAfM6QLf8ARVI7sJfOEsC90VV2t5W6m8rqvs9G+E+wi
nNOCGf7FxDMY7eGlCUfI2HHeJgQFHnfyZB/SFHi+ygna15NISaWOrnB168i0
ghbxRnIYQiiKBULe9lMo0AzzscxMf7qPMLS53XIngcrATMszwQbhH56Rc+Fr
CYJNHXc3Yjm69m4N2tJtaa5ltl1KDfiIz8pPzLHGI/LtMg7D8EfrbY9z+xaV
MRotk20yDz9mGblP11xeQWJRQXkTOxTQbPNL9arZtGMCQ+trzKbIr8DvdhDW
QK9boyi1xoBQZTxfY2SZLY84SvyPx5swY8mLcwVSOEmR8P0w7d3Cak+65zPF
Q4Hemfox9V/Jt/+D5WfAcwX5zTOBiL/uCfcxLXljo6qhqxDO8UpnGl3s4sJN
q09SCsoLpPVbxyUb8/sadGakYAjVigyclqahAsAgc1eQKzgA2lF7qPH4Y0fi
uTMwq+8UK3YtdrQj+d51/ilv3KtV1ZhHpvdnlYPGSny2XIbT17yAn1CuuNCv
lrWW7FGPGcC46MM9Xjqe7O/UBAhWfri0X+5CQdLG8YwTT3fqYbOxkSuhCeLE
6KyTFQjqE5FisHavby5cPzhEvjPEiMhnbDPTSm/uedYCGb1RBMifKA6wkXHZ
iEQymQx2sDVdlU/UBK6tgQiEN1DKMcYYX1ZzrRP9UAYF+piohzoUbFOgG9FC
pRkZvhcLw0ojifJALK+z76T6V/1A5iQCrDHH5+ibuO/wwM+0wUYVvfljx7uG
0oGZ+swX27gxwmGEjkgJZZAZGRVxTXeNk92igLKom2SHihXygvAJwEKp2v1b
8D2JkcYApwP8GdD5eVYZ7KPBv/McHtGcEXUL7iLCe7o9ZdezOMcTcVkXfkpk
bbEOdwckZz+EHxiNWJyLExHYtBUh0fVZ8OwPj/CVvvOMY/A5yu+HEVIN43A9
PGb3g/j1pG7MAc/XOIJejN7ki4cdXLrSmdfVR13C40cCgg0+KuWn6pULhv6t
eNj8uVH1uh4rjDmiNs4zojdqeYPpugUoXDP/JzIdzzazWQXqWP4IoZI+RCjk
17z6qT6aw79klb3id0IrL671l42nMz1GbjaE/l7o3NfeMoWVvfwzAx+5LZVW
1DPFfRHuJIoou7DXlOPjmrDjnoiSr/92Gd2/tT5ezHqYGNRH/m0fS/v/+q6p
+n8gpozhtMRuPlSO47FzQ/Eok7eErwejC8GABxfRfHif1dyX//z65XTNqBvj
EcHaAO97ToRqNSEGWe7Iffk36/TGJL+mv5ru727Jg23TPwkCqXqLE0JVurrI
t/K4HHAeE7bzVIIDHd4YlMX3ndiAhzRy/j1nk/hWWDuOogMu9P+M3yeCk1cG
edfdK4oIMAWr4+LhwI07VdrJKMlkGj2PAq17cS/3Uu/Pb1Z30HXDBr3XB0qQ
zFQhnwihOsnawt1EpLYzY/DFKdR3TfKT1eIuNjv/0NwBKXm0hr66wAkP1dc9
Fav6HVqd1O2XnUxWaD1ZxlC2HOjFOATvF4PiVxO+Ht5w28RiLzY4PhlTAVhu
lxQGuddrTNULoqbZ0SXrZgQwoW/fMMRUprc6xDfeQtsHNU3Tv2e8URUjeU76
W1ID2rwiIGjRylWvouQ6ILGjIf1SgKIC+Lb6/5B8jvdVtlvX0Gln3bEy5Yjl
GMRfI/ZnmIbyI0W5DiESt8x9/otsUuXk259MoCwIClNu++Hhuga7umt710qO
7eti1jpHdm1BaSwuztC7RtuQVRbhHIH2HZfNKNWEXCdfVuoWRM219+SeR/9C
ZBl44DdRqjj1sdcaxwhHPtOe3CUUzm4FjXMkOqwjJMRvGKXzqOaIzKhrdTCR
o1AHzJC+o6wgKWeUTx2gbyw/r0TUJS2Jrd9zcLrNbxMiuuBz1z+YoeWDPPHs
TO7NWTXiol1REP3eVLwcZ1zVzUkPLt27sJd8nF4rwUH0KUNet+laxwNr2B0e
D+E+Wt5JSutCVWiMiVEOBXuF2+jskQ3VLUoxZ4/AhvPj6l53Y0L/KPg+iouP
WLCopc25h7BUsHPY8ktdGlS2jgSycD+AoUcf3HyMANrmsmRtmlCZFODc+SCB
0c3uQXSy9R3u4/PdofzHAmbSyyswKPfk0aXPq2qs1fK0r+wqTyx+6HRlMF0h
0krnFYqepAsbwfyK45ED8X1Ev1EYduPa+NwYbUbIwsmKrp39q4kky5qKFGpx
ZmBhDd52raUJnm9of5P1ldUGbNXJzcA/d7aJkTfB2d01dYHOwBa0Pm3FJpLN
WtpI7n+qPZJJFhVg0Otdvh6Nb+Yrp02Acdg+zgrlqN7+x4eOhgUulqU/p7cB
SM3xxKGu/0mtWv12K4ZpLB5T//ht8S91TLUNBaUgN5TKYxQM5tARgSwdFEFS
w0Y6i0jR94h6FLwNYzL5kDHmOUGbIuqECFl56nv4sB52GC4b1MJbOmh0Oy8f
vO1za09LQz+ZBUbC4XN5eSFE44a0Ed6rq/nbhPhU/4fnG4mzMUtBnrhbB7Dr
Ws9uJuIAOg3K5VfgeV16ImsFBay6y/ECxqxjje7KV7MleLNgJHOufWFxCnil
mzgce47uA7+d0lN7hMSy7aY6GnAI4fYPgc8WT0KWgw6VznMtLmIw0duRTTVH
3d6AdCuDW6F4PReFcyZoN4LTT6qOwKAq+WPt93QxcO1atOWIcqGVOg0Z+64w
JLC5Ohn7M9k9xekIrvMPKScC0RndoeM3EToo848KbobftxxQsXoV7O/RvpHM
SdQ/WVDqxhPO1a75gP2+nStm0fwh//XuDMATBfM9u9Umdudx8QqLsYz6YUcV
vfTzoe1Pkj8b9vfsV45CYO7L6HZHkzDI7ztIAMwYdusNcmNxZMxNhlX005Zc
7SXiyDgxhHxxJ/JvjeeDSUiEhasIOP7qIKtakfpbjIlsx85nHN+Ii3bRqsYf
I2oi9hpgkY4JWYn+tNvyZeSPrhGkImWfqyzWnn8ctuf0ic6oggreyyW44M3H
v2h9s07SzLRioLTcfqRVpH/C+dygsZ47E/hgICDpeXlxdtsmOyfeDsRKF8Qx
NSFNX75XgcKcbv2bJTG4+RAYs9cMm1MsgBMIWDWU2ebqPiteiV4RUig4Wp6K
wy3sV4OvSoWmJ4ChYmCJnUXEKk96Mq1hB07VVedQhHPw9iXzDfSoxOUiXbwa
UcCt+HGpfBtyxbiM/4YE2spFxJOs8N1j9Xx9TFFdyUVOohIS8mX0vykiIhmc
hVizlht4jJFFAvpOGLNJYOj+F+2uwA57KPocNO4CYP1eX3M+l6IiomVXXCBD
2tAmDtTFBsNMSvrmFwrjpUEqya0CgARyvDLT41EklotdeysXP23jFJ7SBCLs
V5lUK20JplPePLbeNF3cYkBQLwWPG56CrxBnX+Pi+pRDzRV1B0LuQwk0L4rK
gvrUP/f884nRxCxS0e2KRotGeec2Agu1sNtzbK0cEjovJmiK7Bk+H916AIud
Dh02O8NGcHZ1xQwDAbXFeRgfioBiWV04l91ZwUq5rPwqv1wr/l1J9d2knFdP
p6uH6Gb9r8WIb10T0A5sR7t1cdLuMuqsm2uvD4946CxOcdRo4yQncaFnxW2a
Ko7mcR6RFuYuwxL8xw3EssKdfKkoWdGM7ZBjt+drcS9DnTHUmIcbQqK1/2G9
q4wtwEHs5Rrj8OzRhpDwzRkoCYz0oe8FhstxXdI5oLFFsgIck5rLJutiB31l
lf0sSLJRT34VzJ1+fqqWSaRV6kc7e4CvzIGXE7FYw0ZbvHyYrgbnpnLuimii
DgQdIvLLEnXwjp+661mkZTwWHdny4Jql31ps8YjI0YLaC4ow7E2ELgc9wDLe
9tD2q6O2E0eajtKIe22MgtTBve9Cp0PeHLiXfSVLNykFFBek5OtCfQVIkWsK
iNGJNXJp01xobP0o3QTl7h4wUGw3QIUGZi8rebwhpwB76RtCNhvvwPWwF0O5
iabkRjUtuPMaw5h2mOxCT4NQle/hbSh+IUeOSqOE4mWZGPhLYt4h/bC80FSi
WYEk1pWstZMj6Ms2h4WqjLoycqFxNL6HvY6iW0I4OpOs5jwqz2iG7PYCLHCd
+qKgr+F+Y4EJZlGfSnenjH9An9w4jLUOFyDbj+yE9mUfS7nYGr+qknX3Hyrg
25u/AjfGH/Iy4iWfy19tV+/pY5V58UV/UXu2J90bbwfTaqe4V2wd+ZIKPIse
8Q7ru4XfDvmNifv3/pTAG9yz6IYChw3O1f87nc+ce7SYMkZqg2sOlqFaozg1
JVRS30gya1soW8FHmqd8ATiY1WGC/5aRqtP9oGiPq4e5daG+0m6s1grAeR9E
7nAzPaB0k+vn0D5zizsn5f89KMTuf4MQ5DZYFAXtHmmPGvAnhL3692VwZuVK
aH+FxW1B7fThOIdVZpwCB9EKJp6JYxqR9Iv74UOXHjKvlYi0FcbMQG7KmPex
TK7B5nTKH+CIR1cQMXbwmJzQ143Mu6QD5claLpT+bqt1Ry/B3h4yBYS8m0FU
1CLu+jJl4b/C4a4ef/U83UmeI/AthbIVyYfKXUFkOzS66FBtnjcNMVDPgeFr
04GwRBm40+p6GmzorXHEdIWK4aCAzdJ5/heLPrFD1GGSUN/C8KZO1IlVmmsp
/bOUy3BmuCoMd+6TikRtiVAqAS7FrEQ6gMF7wi8hVml6lOugNlPtFvIGI2vR
BJqEmhWvlNQPbJoQ6Wa4wxUW3A7VRdB5B/CbtkY3o6CMqNZhfRzjltvlyWXO
TxOKq1M8ScSWESde+Brsqfu1emzY8/xEsOMD0qjNXk+F6ymv7X6wKeCNi9lc
unHpDgD7l1hLNL2qpjEJtS18Gxygygp+aroZm/vwcSB5ldNzZuU+xEAPnMRl
WG2ojrX/3YfJmjxB55ypgbiEWMQfraNrD+Y2UddWCK3eM7RGbbI4JvLTamKy
g9E0NI8BddjiCm1DBjwaushOGrCJNPUwQqd4mIkXEZJ6g3iqZYkrRIUuJUBY
gTHidT8EzPChlyiBVRharKmEZKt25miAS585PC3MECTaMWua7VMRh5E/CO5k
RFcxiP2bkz6gwrL+bFq05k4DAEafUl/IXekoFWVyzOgu5hC26PHmK8Se6XXq
yQgfwNi1RlAiett/0fqIWtv0/LjSBLH4oDGQfIHghCnvFIfU7/BXtBv1KqY0
9RwB1xDx5KBNQfsqBnKwYAxTm1q+1ryqjg06YgcOisUXy78ye3P2uT5JwqJZ
IIQzeGmCCW0egJFx/X1mbkYodFS3z9dD49ZNLPNwL2cyZPtqQR82q5+O+ckC
Gga4MYSp1IWTfQ7r2lljSip9WwSdM9OtBpHKimZSaHhi0TQETuTjmxWmPz6s
yLW54qzeYT83W6cld2R2Wp6081WoDP72M7sv4a0ZKZej5j4qiqbxRur3C+oq
hjPJoqcrgGw49349IAAABwDBgyJdX4vfE+oDknGHADpcY2SE/Fg4qo912Yid
gB4WlsNBHiVxjXVHp4kWttoSbgNjOyPIKvqcNDxbgkp8vn07HdE40x2XpW5v
MMmJQDiotVEWcDtgE43oaUHSL5Ayn+0abeZKHMPBca7gqzKW6DDBL1lzis9I
q5299SMV6epsg3Rx1uKrIzABb8KPsWepYjMnXGQ9RXLDeKQDCrOUGcfD0PHJ
KSETByYAfjbOp8E34MLUPKOKGN2wxEhTyID3Sj7gdqYviHyzqPJSV8+rZqf0
jpxqiEyddkde0FaMBcE6Lc4BkzsLN5yGdpn3r9fjX/JOPPVJcDDnqh6R9UlX
Hgzb1fwf8rReodDouvTg8kOkYKBjdtJOKKIa60kLCtZnc1H9EEMxHpHFnLx+
WSq9GVwbtwz4HwpZQyJX81s6EgF4gBBQgiIdf6XL6Z59QWpedGl0dc9oBnmd
d1AhpP8Eu502omfh6nssGobPbJtca4TabJHorcfkDgtGz9ScvLLt4dlAigcc
p0UZn6rrXQ586Xrlns+lNqclOJE5Eylqe9GXZck5fODawVb71UW23q8G04tT
Yl4L9UJEpnxcAtOTK+hDnHfw8Os7xmB3vr37ZMtmknQ6Kq8TIBca3Qsmp2VC
8nEfQwn0m39aRFJ2Ey6Q4fNpV/1R+S9+uN2cuk5nfaFvRaarQFlCYbnXgvsF
LJxnxDTv26jft/UN1MdRSBMBWEwa7F5ZfMfx34RE1QE9ND+2qM2DsPl8bwI4
iTUole/dBvx8GmYrE9NXW3rn8e1/LBXDQ7LeUsT8AUyKPK9Szd1YhWmZz4rN
74n5pOZg0vZ+2D1JOCTbg8mxOhi4Vmvnw5Q3dcDO8V0IUvMG1Oh82VUNrHfO
eb1AdwL4CnI1cPMfdW06j7O6JuFrLtVa3AoUGYCZAGLRiNwGl1jrbPvTVQWb
bEAClVXshjmFdkxrv7jTrIF2AxSM6cHX2Ck2xkl15YUKRd+slrekQEVhhWlq
rZhQb43V3ISUMTUTAO2tc9zgNenKRxgR8LI6at1lyEn2qGwX8nzx/lhxBUDN
T+Ef+Wlz8u2SP+I0jI0sJTA2J+RnKYTOfOkIKppHJIjg49c6ZVIkvSuEpGyR
KDLCmhZ4iULFBLQ6Nqgo1hNGt1SrJrXcWWNqMTe95jdgVzWhuI2GDutFbWsP
sW0hkYltAEDBRW4No7px6H3Iov2RT8qfTzYpe1d6BCNV1sUPYfKfQKYR/1Jr
JwR7jusFEp1xwcZVug3GEYT/hSoyvA7M8Ycv2x8+hR62+d89rhRLO6yXz7s1
A4DW3FBhAYGOWfH3bHPbZre+7qMiX1NRxoTWTwwehyncl4isEFfGi11RmLMD
B0sRsMv9hbh6l4hYgWjOd32TzBGZ/fF1mtsmPqHtgk6hLXEE4DaQ7LVIZFyQ
T+Ft9qWTJHfh77z+UZp7C8AIvrkdffMRdgT5pGthjztGYsSW6TDCmkxL0hVJ
iYBe4qzsnAaN77ppjxNpHd3v6gpwCbRgPDLSVcSjFJNOzTpYhh46PiEfSYHr
e+3c0aVQtd72PH/mM1+1HDkiSL6hbaCvJ7PuhuhBowgmxLKU0dlxcwi9Bb2A
T36L3a/WvUcTE2SrItGWr4HTT4UwnjhC3hbOX0I0JemweHQQiUwz8BX2IEKd
LK+rWsodemDwibYYSecrFKMoEJXDxbsNyo7dKvpQqmAHXo6Slbhx/hOPjgJT
qQE=

`pragma protect end_protected
