`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
ClN29tNILxpWfk27Q9ttAlmDAmgyJpZ1edUGzJEWiEqrpAY6einr0JQC+MBSKTmh
9olXTYfsr8DiyvobjiWAgjzc7fGahJX0VdNdDX2L5nQJ0dvDWHb3PDKhYsSeQ+XR
+y7afSQKFo4zEcr8c0kVOvXi9UOT3J8LaVrluiughDM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4160), data_block
rfSiaDnm+KA8KWq0Ky+5mh268Y5CarkPSXx2gx6PN26nT3eoc/0ucp4lPIaUS49u
oevgcOhrI5zCooZEuSRSwwq18ujOVttO2xBkS7CT6Z4xw9eu13IDHsHYXJr/0ckH
2oufXoqzNwT8/OXNahCtSTM84iaBEf/ZwoILxUhiFzCIuHtFhU+C9P017P8rB3jg
TDjC1nVuFdWw4sndgvAu0bA8FLm9M1N1ML0/lJtdCxvEqsRpABWsSyuowhN4GBaf
gCWUKPGdV7/7twhe1O1uzzr/D40fX7VLaKk8rTRtqtVwhML0YIRST7fKKuRdpZ0X
/tQ1rS3ipQ820AGVqEWV3DwWH8I+/c4NckS7E/K50ytBo7gz2Xl/E5H0zvxD38zG
01le85yW08+W4vxoKPkQFDhqwRRi0BpNQKB5mo58UO2ngMHQSf4nJmKv8q2XsHN6
ANYZzlPi8WpOMIcIuJPmrsb8Nahvxk1HNJIjYvEDBEd4bFDOP4dD9SqME/4vWcML
FFClx+IRx8w3nScc9LGpK3tFNCsCTB+pp8GA7Yi6beDlF+NFunTjQy2YIBIqPuUU
pIJq9kvgaGZFPq1kG9blnKitCQpiw+6OVnJuU+jihJvQ7DjVUbHYaljIOeWoyNJX
trRc+wqqMqAUoZoixyRCzniCHMXvnT3lmCaqOjlwXOVNiQS7uB6jT64er896KY7T
ozPUGRJDhVDskGSL/vjrq/GuK3VUtdsVmiCSkIfpWCaajo2ySIn2rH5WaQ9LAbwl
9QiK8+CanPSzaS4yP2dR+tVRIkigafG0sdPZC3cJ6mCagbJP+jEiDxz4Wr9p80bY
AxrLXym0ysHskoF9YL2HeSyXXunW9xcALsH9x/8lYcK+iSu8rjFI/StK64fcfT15
WnhRnFcX8wnGGeFBb47oqUgWpkrBFCPMTsMTUVX7KHUd0HhBv+5IoJ0ttIxmteKr
EklHabU0MX0f2KlOVk1bA8DE2dhuSSr7Vy5sfGscs3VIpwqitHS1WuxY8Piq/3Tc
8xP0z3xT9KIzHmKfzS6fvnLBgcERb8atIQlyZ2CcYUPFCq8JYTIb12z/kVdlPdTl
onMyFIOZGyk1aQV+qOZPbPIUuRr93sSkhV03vacm6CrkKGVB2a9gitHiRqphENGq
SSDxpLCqZgME+AQmzLEaM5ohwscMOPdmR7W8b2Wzd8OgVGKAmIjX0Qi6mG4vvS5h
AHK2dpeYgc57wOKf5rL3Z5gi17W656UTaAVJtDSLqsmzI0+t0XlclEUyVgkLkJ1s
xhrezouIAfpWoAXqhSIelC8Gq0SlExwtPBhi1f24lDQ+SyJsUFzRax+T1KM5nEwk
b3yaXtO4WTeAUo9BfNWkV1LzgOG0NibRjqlnAsUwesJCNv9+X4svW9BL6Q3XX6uM
WDbWo0Q3Fd+8Tc1+zlHlER7/YDHFYO81uioVKsJnXPsRMji84xm7V0rdNIwoUCKX
aJoYZWwVE/aiSci3MeKi8+RrmxQ9w7e/wTZUk+Dlb28jU3yXIEioysrFSmO2cINL
XBUv5ls8esMKl02QXBdzmMG7mDe9gK9PzP0n0t8Kua7NyQK7GYvA/IENbAIzAtPj
Q9qgvl4N2tVeXBD4UZzdGfLlsWwM9aWtutDOLGtcZ3fC2rQF0R6Eof7hDXvuxs3j
5ttJndEHKk3gy2KhtPUfUnZ9p65YEQQXbkuVdj64erovOeuFpKWT6onYz70A+5Ne
aebCCyvER4eJWO3PcX6Q2Vxd3gXySH665qzwYWslxypsyFtFR2Xwk83IR8deqKMR
d6H3I8lE/D5KzATxkSxdAkOytw89fzPq3GQeMM82GCPRJ0F67T0K/dbFlNaoNhix
dkxEwhpmgamscd1kWp/hNLsYRVUiuu0Sgy9pdehVe1ayRGuO+MRhLTNX4veBSlVU
r3S88z/nTFC+nTQz+ZRokEMVs8Tmfe2+bru9144nPXaKasVqLLTmIoLnil8+mJb0
bl3tXfs+ZgL5sH5dWsVSyHwtLyGRuJltDJDXnIadIGfwlwCMz8iAblPBdNe5RWc+
0NPSNAVwNwiZz6Ri33jZZ5X1yIuSOmHWibRG/tDOvm1X0IJ3NS+metalGDM0v0L+
lQ/Tc87wvdrEO5CgbCVKCb3CvSaSi1rseuGxGmnQ5m8LnoWwaqoHKEdTmNXt88V6
p8mWn9ISzumrMpgF142BsOm8od/7tO9gLtxLyx5I9ldm4Lru0KWcCygg83QWPRMW
OM23SC/zp/S3XMi+HakSq0dSjFsUHyimAJwaUAtXHHrbPWmNhbCzgBgelb2oTw98
uirD+BerSRcfXPUbFtlwtAb+J4QuJTMIn0iYMDI6go9dr28vA6Osfd2rF3ihySpB
VTAnhjl3ACOiynsOVcUP0QlHuFWksyWKfYbL0QQBBRHmucaXCXQ/bI0IWvxO7LJf
A/WoYr2x+zAqBYAq1xWlCYzPsT3hRbFtHqJpff6lrfPEGcmrJEjTOpY1i2XAqWzB
sGVsM+e38Oyhad9trJJQ/u4lxpjUKaw+NJDjGnsliJ0jYFx0sIC+DbdB/3VBaAgC
zA/xUWcFYWNkllJcN+D5/DZKYgyYa4zpFTMT1mjBFVzx7X9J+OOgEW/TYMP04TgD
7znMcLQBlV/2z+5KbpPXLxNV0dOAoCS7CzZ4AgOMAt/ZqbLdgkMoFFB1psyvw4wf
waJk8Qg/jN6HMUaPnP8Yu0hhGg1mrBUWJsgO/P3Padtb3ZJZYUXI6Tg1E4I1KHVX
qFpJT8VglUfHraW1Q/IhlnXOUpzGXBW9QelNjL/VH1ADay/HD96lsCByBhBo2MY6
Mh75XPufQD73TMfQNdQMLlcgQTAGd0gMEVNO41oXqtPP9/VisPglTOYG6nff4q2w
1ePt3kFaCrZICvP+BFEUOXMjObxo+5Ep3wR3N3trViAzaSKFilTkOC2sJAmZAqZx
jI/D/qrBMirljBOw0I6wNm9NsT68hFJJ+3P+HrVUBKZeRwpZj+yVgL0utzRaMrUx
EusOlM82fR8sAUGFSFkTnluWzidlnHrMij1U9mNyGnJIdOKTifpggiVT5CgJ3aVB
In8Vw0LQ16/8VGQDzb9Urgdsd44d5od3lJutkhBNJzxJ/HGcpWDu4fh/BM7LTpH6
afqeYIFy+sKHaC+RKxP5c2h4F86rs74btiis/pOHNOkuZdhOVhXfMCL8uaK802KD
QPRN6EawkOnQ9uvUe6qcviwaHb79sHhwZJYgu+V5Z+O/A7zu5qP81SHTaQzLdBb9
92zmn+ZYDchqF4cfTHswz7RsqoF5yFOsu8MVR0V0BeQG/T1nWkTj5j8LrI9yx2hr
cn+wOy9fmVBxLSneNq8LleX1zY7BvbOvaocrGkmIMpejPl+NjOOwaO5N7HnoRxS+
P23UDdzRk+qnWq03JfCYOa7JwVSXoFCesH4NuJzCWWjXj3SFRjyG7plexE7gsOGd
OTtKREonamUlw1qUjCnKHau+sitd5/UeuxDJIg7tdi7I19TZSByidPNib+3jdbFh
Y5iemEx3gdtAWcQBL2CeneTngIZdumdYwaUctdmcU5+ioHw0OUiZEYwli+U5Kl/F
kKZFuKfQhvKY/b5ALqY2wb56tdSQEc9Sup+9p5n8a5ma16wBKYzmPuvTAMwsQtDu
5hhyXZhWwdxgZXrcf+SmTfLFU9djYwsuN7Z81hLfc5x+0jswtoqz4Uoj9FIKnS7U
4yGIdndYm87boUWpPSSU9u+/43EFkNHuuKalRBGbNug5gM/JufZy5x+55aL75bJH
pPWZJwuQz8JxbW5w6zD9n4AvBvuy5dvhPaNP9ZN3n++L9n7josraMzNlv4K7+lt/
A6mBrxnsUhEyAfF1pkAPwgwcgZwjYJ6FBNv/79+Kz9o7GKJ4Ekrh1M0JWpI0GJic
Wkix1BlUqyjAy6zlQcQbDJPHUDR+YZXjTDJlz9VqzG+icPCv4VB2hUF16DvzFL/1
IwtvAxZxTK08F2Q++iGkQWKjGXTe2ct+sGLAvJs7u1vCpR15UWQNQESoyWBKKqQH
0zgH0TboV5tJq6ypYLKojbp390KKkTBSFWwcCOHfxohWcuDAXKSEO+EvzTdRH2jT
QjwXNOAv1tpxmvHe13P/7UL2ymJqUSAg2+19jbLzuCW+gDE+sE965eHP5sO+nuCx
jUBP+QquFmgzVZrtfI9yIGunmh/JfB5/yRwF0V4BU3BW6vPta2jvOgqlhN9lq6WK
GyyOt/3svWoA2cqQcOrlOIkp2jWAjMwAb3cAFY6Fc/3WnzeMfbJWiUf34GyfYb5c
CagxNIF+M9My3I39HalQIe/AajFxpYoro5/gF11WyoGGWm0CvqTWkqsXvo6WpNs0
E4rhjiNTwc9tUFTX/Mld9FRPDL2cQov6biPvu/VKhMg9rgukFhJbXmn6p+VR54VH
P7vVBLeJcA/DAGhTCRc4xr3kw4NPpT7v+yPVnjMzcGsV7R7N0PRHndQNEcYC+XWp
TvOmMAIO4lUP0/Vp5GeKKN1Ctk34O/6fNBzFMZcMYmO8yJ1rr5Wq/U6tJM36q5IA
9xME1+NkJYWnmbcDackuzI90qOZMt9bdLwsvFpTeyDcttI/tfo8wgxrUzzl2uZEJ
PfGAjOCBAjCBsocKKjd9GxRPQGzwe2h7yVqaX8xIMySal4X6ulgmEuEBZsyuFqr4
Ymcylmlh+vDV+0hI86zwuR1FYRXyB4hjFOLTK1aXu132Kl4YVAusifycKsk+aEGC
FpCuc1exbacc2jsc2pHBYAXZ/nBB2MQyYi0tePE0CMJLfbxN8Y6LfMogT8PtQFr4
9bVA+I5a42477igjMd5fLXYR2Q+N7xZGnUkgN2711d3kX6lGLY+GQMDqUc+BMReu
JL8Y40+3QiXhd6js9LeYZvlQ5w2exX6Hnh8p4iJFHkhvqvUxPYut6tkH1vq9rU+L
iZq7ESOQtilrvwPgFEBMLtv+b09UQdyt9sXIXc3TnaAcUr5q8yCafMuQTJWznuzm
eWjOx9qSmJMKdv+PoeXZQGMGUbNLp67yBeCj/LC342fgKPzUEnP01GdoBs9zyd0u
Au8nSxQSWrcq49zBqrWiNv8nVDX4Xj1PGqqvBwCwtfYTQ/8g0zT1w1Lh8QZK4zxa
KrMNjSoFmsY4zr2XMdZmzHhg5VRJfD58PZrHOyRoZskd4+D4VEjj8VWNKg0Cj1qh
bKeSLfbJQ80kA7eCdUH4BXfkFtcQbJrejvWFO09d80hbrpCh5DCts4pRQIFK7BeS
3GciU2nfW5fKpRqB7cvV/nP/eXbQVBzgwSLYh7HhMitBmuPn8+QV5DyFHQGSmf7V
vp4HWNhOj2Ns/xiN0oTcUg/F3p9IENg1bceVhb7xIVHX79F1K2OOCiqp+mx5qUxf
bZvtNkydtqAl4VeGjDlrFxS27aUY6xXqe6kEXkM4av5yCjS0UJi3JfZtk2Q7qPdF
70QV+CqPsKJrwCNe16UHWPs6AHDwBl8A+6FKqlFe4v6xNT1Lgm08buu2yMGvxkPJ
EqljFoLrLBJ+Uh7jL7VEEopQYYlCynkm4oaQyUnDUlU=
`pragma protect end_protected
