// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jhvtq6GXnwN/A4elYnYA12V4Tq6bvgIlUu1Yrbf/s5Ocjr2HSRj606cv10Be
1bcD/e4legfEkim4H3XNORGdRlJQZxT82+q2WnuYhDOwwrXnAPDBF5f8ZLhB
MBDQUsI9xb050uXnduE1UQ53a/7KkTtCvkoCEMzTfRngpYZjl3yDYD4BkMx/
8PmqSaJNJe/5d7SZZk8g02rHZ9oGg+QfzYIqnP7UZcNFqsuFNJv5DrmQuOLy
vSLsS2zTN8eR6Q8FRo8WiENucRtLqagP9ancOYh35iwu3d0vJfCZlaG7vOY1
n8oRSxwZPiqDr2VYU3qARQT8Uk8hLRe/69mZmoMR8Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KIEGlJbirn/Q0hf6o7Lat5RWzgcY0cinxx9OUHagnNpANRAAShgj1yVJFwin
k916Lh3Lx0eQnuAz5mw2sBQWiqblwgUTet7IsqPdJuPDU+280rnzlZWGAvfS
uL5Dv7c0r2zJogIl/XGeD9sTh1cXQ/P1ITp652OXn/Q4zmUYbScRz0+xggxV
M5+JeCNLxblzyLfQ6ZsHr/9N8aYnB5UQTE0TNZHTFNeijCDj247C2TWX/MmW
gdeQSFtp5JMJZZDb1rzRXZaeoDWHsX+Z3zU1BX82BkXQQtYemL1MR9U1RQcX
UydIlW436Ik4Z5PPz5SETsM4PCBAADr+RKJdBhSXHQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AH4Ch5bB33duPjVAUduyfryA90mR67cyATkwWzxTYPa1mARvwK9tANHaFZVV
fAhishW9EbalBeYDq8nE5Ma+QCdC5Ieqp6xD0Ng+s9JZ0wtbWoyBEDuzJvCP
Wv1vQflDsRVlW/bVi5+C75TgARSThbfVuOrd50gZZxCo2iw/9KDk4pFfCgVJ
9XUD3qxIlcpX4k4DfidNVqmNYTTF1L2lfW/fbyCr3EaweNG6GRngQsSHFu13
KeMaTXkHv+ld5LyUVc+vPkkm5YxKZCqZO9Knk0AsIBg35+t24tSU8BbrVusQ
0tBHAb4HNxVY6PpbB7umdzqy3cZQy33mgTDQrp45SQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q3ki1uW6OIXTGacC/7lWTwuI5b9hJDd46tcWWmPLTtQm6J8uC7CidCGt41xA
BJ6A/P/6ZLpUFvNX5YKh/Hb5/a7dtspJ5vzfRmVveS9nCe1q9QGKDgOrwn55
3Cr1RD6dWL28/Q8fxZwlxnAQvwYM3JRzACBk+oNwTrjf0uuXen8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xGqBmCdumlpS04oan29hbDBd1v8loNe6BKdvuOZ2Q5nFY3FXV6tGMRCfuIEp
8Ukj2xlxVoQXKcB73JaZ4tqquzCA2hIbCIRgIGMqHiUudX2tWsSsQstRbDR0
IdNPUAinn7gBp9g7YfTqsmbiIYTEwFZTNXSqYd3zFLgrk/QMajEABPZsvwx/
czqHTKNrIa8YN2wAv5CEpTsBNpWzY48od6rKNMajk/9Fd8y29VAI5x0DL+zR
trWAtSnXr5UmjtFaca6lsEDzYQnqsoNP5XBiv05zqNp3DIzjyj8+0FZnjvCc
KPP7xMWZQKfP932E9sav38HH+9i44eztUccZl7UHI33gqDlrZ8eHRzEkmotk
x6XTLbdt/gv4OSZMYJqB1Btc532h9Y5Gcp2si4x4whFso2uGZ047OKddHK39
xYLiI6+MqlQ9pl9px6L2t1IvqITZegf9YyqK9cAox8wQEb0sXonzsVWkkn0l
CA5SdPMBD8VahnZ1xKtGKeK9kRVNGfS2


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NnRr976TSU7y9yCmzpZRtjF9lUzy+Oc+TJuiZmn9nv1AYM/TfMDQTxHnhrqa
IOse0KryljZq00gf84T58iZXOVJlMc/SotVxj4wRTt40hGNqNO/7N0fisUrG
5/oN7eyIxezzT6aQmcX33GRujZ4V0Of4UIPd5tOLCD9Vxnpzzeo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jrZWbw121WFInoPj5BVBmXSINDfKGpuPxbmUqyGlOvjTXnLaigyxOkV+l58j
eoQebhhlcPKsuBatpFbO7Nu1n4wWukiCnnkEIZWQCEfhdAmAhrYP7KcgAzNy
6wtz1hMSCNH6t8AmxrtqxhCdq3kAeBDUBQIVoxBSeoZaddns8tU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3296)
`pragma protect data_block
CvRTt5+J4n72bk6ReCK7+sYZnz6jY3amTEurK3t4daweXshdgdV7zX7nR1Ey
hQ+eUxr5TJ2yQFNGqYyWC233vqvzrs+gpU51t+BJNf+mQOKyN6rA/radV38H
R0nM2z3x9VWkHSRqFxeNZTTtSYaLZDHpc2TudeaLI5XP/ThtK73ZWsxcXbzj
KXoeCNICEIVbhvfy9CQmL0AGonpTYPikAF0xIQZug0diSnS2jceYaVgWpHJZ
2nh42Vm8I9722rYoDuzelW8We10oa3WCL3w87/mQJZXC+oDnl7oQOQEQy4ot
pxoXVgnAMo4aQb5ybhHRang00q1RO0Im/ARQphSTF6O2KJ2NnYN4GQ7a0fkK
CLQRuohzC5RZyBPINahka4eFD1CiVPPHlY53HtCuVKueycu8bhXJ/lqXqAlN
8gL4xcDn7078oHCitsXDhx4HsZQJnPG4KTOWz/99R8dY8zYIq+3d5Vw8Yfz4
EfXqLu9oE3yoY0yDcp9pq9Rpv2AFvrLGrXTGuX/WqNQrfd5HNvo0jd6/IYyg
WzdE+YvcPlH1B9p9ZtUkV197GEKXy8wHgbV9WDDwcTEU0fzv/whzQavzuLlq
SVLJQIbP7Jj7Sr2Bqxg+bCpYX0tRczxp8aQGKp2Md5Xv9ZmYD2D/Ry3hL3ye
KkWKcZviVJiIyPSqS7yEUklAxds7EtlZkZqmv/LpEcZxPZV7lOcl7K4h0Dpc
zwFpZvGp3AfVoT30g3QXlxvCMVx/r5HJcMXY4GbTj3pzn2S4ocZ7OxiE8Cpt
egtBIMgFg8t3a9GnHziD4z7qUMSg81BK2NWdhJuJHyMFpDpQiwlSphzi4Z8c
qWEPyhF/t1VQlSeGPw4QGG40hS/W8SAvSc5OqSPKpetOCzMUJWTSXI5nP3gY
OphjUWEi/jBohEblTY1qHDaSF7sdGvYJOiBqnA9L5QnLMC+dMwiXzmDh0G5m
BYSKpTWDpsfg2dNtTm8lMjTmie4y9ggK9wCHJUUy83k1UfuYguJAfdCTdWgB
Xuw5EOw00XKaMHkJ9Cl1XYWCgs4HdxbuLQfEoBaFCAMhqxr4IvQdKMn+r5Ul
16dbWhy40Yo4P05rCLTOua4D7BQ05a5BFSmrQ/Hto6DoDNB6Nc5WbfamWB7u
KSocC1y7X3HD4qyEoYfKF639oH1eGwO17PKXa7hJ77ZG0b47FkJkb1bzCTvd
L2v0QWolD9it9pYGL/4H2S75JydbtLKeFNCPu7fyMUnV4XD0uWJFMQ35OnJu
AkVmdoL0upTVZ2i9i6Ak4+W8diJdP3BSYkiZwKhDmDj9PCBQ5FPCIvUGcp2j
ed4k22/7sSXQWeWlgzrJeyGlP6Zmg8qtfvqepEG43hNfZowm6eUpCh3XasvM
/5JQi2tneZtoS/RRKna5UDnPwrIoKq+DkPskKZmixie0sxoONlP5w0eI0rtQ
qj+36jA0/9XvhwIscpRIbX2/BHUxQIgMWiUbiOLsVpc6wV/EvfZIb6IgPdXa
WyHjS4gdkgYL+371lU1VXClT/P202HdE5agp+GvH0v8bGc68QIHmNUZjxP+V
l1rNhbi3zTgOOS3eRnGsCXXizQCd1hnuIYpm3CQpi0lt3hs4/TzU+aIkdZmy
MQqJQzmxWb8KKDg0hL5Hm6DqNKhZkFEMLEvSZlUCarbcQHXNlogCUnxqlPah
GEezotk5q9tBPjLK2/POpXAY9sZREzZzZFNsD4Qi899nUSR1Axw8uSsZARcB
ncoHFYTF844NsG4MlIlknpTmrvKax+0+Xh9X76z4SutJsXYyfZqNJV/S8+zq
yQ7KoXamnhR7YmlR8quy9P8u0Ml+mija55iL2/RKoDp2RRT60Qe/cOXxPURA
FG3E/LxKcKjHv1y7ePQ8Xh3xpvuCRjh8uf0kJoJQP/5ZTCXrKki0MTBxpL3b
xB7+Xe14xG9VWDs9ypjA/FEH3GmHmVXveiRiCzDe8LQLI1ouTGq/L4VK61f0
qGEIly26ZUKpZe2E9eK3JGk150OYN9NXI0hoiVRWcbit1U8K8b5azuANevTb
4PIUTlp7P4eSLERGXTc428aLxF50iur/0Lsb/fAOi1RXTOD5gQZrw1N8uR4x
ZEm1xbOIDR9ODki+V2LDEWCs+25kDYfZzZHaQ5baEKVat18xhZ/znhaSs3s0
jMq+ZKf5d4aq7WzlT6wnUZ+/BNqyW4pzEK3UIJxo36unhllkheuQ2HtYN86K
OQHPTJatVbG8uP18CYaLqcAnF3fbr3/ZyIHqvL/s8W9B2DjtbZnjQAJexbNx
/G84cnXA6WF2m00awk5aAQ7W9SVFMocXNtsZ2y0SLJFVaT5k/tXt5rDCflbU
0+1cgRjKAY8owAkVTN+qc02OIYBdKdZSvb+uWVLKN3uUT9f15htHwGl9nwF6
pCHXcJj5QKcOLxP9R27lXeaLWLAK+z4b08T0IkLXu7rU9ToxbroHvSYwgp6L
E4TDH0ljOb2SHi28Di4Ghv4/K2UCu2xyjE/8DtSpkT1lzFb40jUJtk9ltaBd
4mJ3KC8nKbGovvDHcTPTQaqopmY9mRi676u3X7FYEhefHPHw4TiuqoSJNh86
J9bqPT7ci0cT3Cq+0BEov4XVSRx6M3ZcYZ4P1DOMoS18SY7s5u5c04ptz4jN
zSXf/2E2epAGmAqVnnqehRU6pWj2/XIK+56XCuiM2q47PaoD2650eZsWZxmZ
PzLUT4x6TqtSKD7Jrkc/5+3ppfdVINETLIWftodruLyXtloGNv9dY83Ra9Wv
C5x51qUmMLBkUQVUPtBaFPkm5D08EE6zq+BhXJJs+v+VpBtYb5a5TKEe3mvJ
q6jIhu+RbIfaNy1On/TYiY+QEF7eE1mbwwu6KhYulZFK+udM88njRwfj7rFp
suqNWt8EN4x+mFABmtrUFjVt38XpQwBkfckKyIzVrHk5M3Vijw/JuN6WSmDG
6Z2+yksYfux7VUrNBWbcZ4AXm7xYfIsSV57YHdHOqJwT9meG/Tp4y6jzzXiY
SNRzSTI8TApEAZRyQaYycgqkxJRTs6pSkpu8WwHXEOVV8YO6qBTbZtT6AV3p
AseSPU+4+vChu7LQcNK+QxY8PA7Kh+8Zh0OkjfKmJypIzX6lF9k2/ybHjDfF
dyM5f7v/h7j+XxwyvzCMz2rPROf/t66NGxHjCdvlcnD+pLOFOXoTqwe5esJU
vWrTMkA60rpRGGQS4bkbwyP8tRTXHTnWeV5Nfn8/DyCeNbI9TTYpWwJ+rQsD
tLC+7Qxwx5CVemPlGOwGXd5VpE7jStZfAlF2R1nGvqSKDWQcEtiNHROY2tSL
GJ6GD8+aXVAhaiGuORNQ5e5t1A7tglkxR7xli5nl6cPOMKWukK5cHhLgjRZG
bhPPLl+7l5P1EYuEIJfTgalV0POX53KYfbF2gQ7uqxcgV71PmhAHhjWK1XIc
Vz8OFFknbTgLUjgTMF1Q+zEhGsu2JKz39d+Ip5cMXi50NJSlnaNEn9qoBJLs
y15iJGdi916qnzbNUx16Ar2QQqcqFifb97UZiGsXfOMUCGrdl9bzXzWPKwDD
WDSh+75FrTBnWThxeV1ZcNXO+whuVAzU/nlBhSPgOP21VTTcGTpTggaS8pGZ
cUXPWA0DVYyOOF37mmuvluYbOkL4tm0vMnObxd3wnnlx/gfyck5gk2ledmVf
loqcsUZdHPqZlZEiXwN8uQQvM7wpMTVUC7kDeNxJCUH5YdVqXJ75EMlsHHBm
UKGA/GbvTjGfYs6Wy1xq9dEDjSr3Yi2H7P8Tv7UPpnO44j3agKR1yqRVFY7l
g5+B/bsCawIiJp6AVQBLrPiXI9Ts2nkMnLiFbmwmvHwV415brX2ICU3iVc8M
1kh6o+mftWlohMQYo8iFX59l2IhGDP75RgVTGUQ9MZL18tmCUGSaeOuf4EPA
L7HOOOCDCyU2IffGewAgsxHUwkPqKrRmWEH0WjP3shHZL5SlAyJMos99T2zG
1Urpb5haKcxYzZkTTSanYclCxCHS/zUuduz0j72ecvrAJvjg6PdclRwiS9uJ
HG5AAEOKKAut+f5Z/0o3KoaAfnxV9YGcKXMyVPA9J70yptpTpyd14M8OTl5q
XQwTbuXGZzXCIaj7kP3VDxPOp0twQhQfcC2EDh+BOsbFS58z4O7fzmycZnWJ
cXa/YKDeB3bz7SLo3ltWMDjsjeDmVZTDhn6piCcvjcbWfXjOjPaAh9tr8wKd
cHdqHTv1kfNg/COKyEjhV0GOO9heTF9Xz4KISn6LDMNhqAe7FAGz5WUEOhAE
lQtARe2cOpAma/73FSktgeRRdRA8cfD/SJKMS1vxSmvm2W689NIr+y94b2RH
aMK69HpQVg/2KnKqD+qy4t7jKjo/5qIonr1YK65hLoWXVXnYhGUTcIDyfKq5
YAY+pR1ZHB5ksqU=

`pragma protect end_protected
