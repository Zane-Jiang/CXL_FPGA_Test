// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8yFzNEidueoTrkaFMRkOM4yrfXyb7/D6xe8pDGjQw183s9wA5AcgC0TFnSMV1PfH
o/liFcI8ZsYvjn+BzHRJA8e4IsyR9osn9ASIN2w13z37Qz7+gKiutEK94V026/Xk
hntA4gcZcUirwNIvKxJ6y6UJ5t1uKvKKWfSH+Bgzu1KwAtLNLaFs2Q==
//pragma protect end_key_block
//pragma protect digest_block
3q+KoVsFDe7ACIaZp+ldP5JgJW8=
//pragma protect end_digest_block
//pragma protect data_block
XtPn5HsnLQYnV4J5+UkzLnkGY2h6B1uQ9aBNSQ7o552BaoDLoKLm5HXxCoLMjrVt
hFsJQI8T/oet+YEN8TrIwOYQ0JMGmuaA4fISsBasTLC+L5dpJ3CFzxFdowr3TTo8
E7dKL4p5KQH8MZoOH1V3BDjJBVNjqXIWLvpFY+VTBVeK7mokj2ymJxgTpEP7uSyn
m9dI8c6iqLHTHnGMIUHG0Ai6oRiuC/bbjW/1iafC7aayA9dXcUzBU/1H+o20a9/z
FwbKeu6+lD/2YMjq69oVTXIab+WSb5jQgbLJ6g0aIP4K83bH0Hm3XanzWVEy3PGN
9VldAHYKxRerhsvcw+NhKJobhD/7Q/lcZoriucePZ4A5rvctdIQwzVCJCjRhue3t
UHpP5BOMy9sOOX4TGO3x3EUkBI1WyEjRWMWhWSEFQUv5/Pe3uFcopnA0lKZjGGTc
FU2Rkr/auPSTOXVXkx3bGLKyJIZ3HPgNhzWVOb8LOJy5LLHkzJarruW03SbOQ2Rh
xqsfvdgc5PokZipLec9kEbSAVjmO1HxxQl9UrYKrwnmPiLvganjf+Suq2Yq59qcv
H6qzIt6wkKo8uktYxerAcVeSTGuoqLDnLMz2CatLlZxwm3f1bi4U+xhU366tc2vC
afbTTbUEPUAVZFyiV0dua7nhmxkQtbDh8zmh8kxS63FphP9Rz3MS8vwpdja/LfzL
OtuUz79a9sLG1pHTyntj5O9TXQWBDN11uipPqjKUgUZu0EwhbljdcUVWkgHuaoxg
/Wr9OGdBe8HwjL6y83LdDeyORhvt9Q8RupxO8YQIrxgtMdWUUEkPW+8AMMaZkpAV
X3upz2+AHv6Q1eJynhz7jPdGuZh4BxhV0Ucb9CMmtKhLQCxegJQdPsRKR5isThvq
JmBPL/fcWofh8VWOWhMSibFpcEajn0DJSJcdhBXrTqqpj9E2G9hLZobhmHzHYyiI
KoQBlTYs83uZxIT6tHonFKrwGXPwyak8j+FKUXmL+ldBnTMYxFkS6UafbmXPKMCa
SStur2O92hFT/xBc01/1JpKThfwmSCB/W/FgOf/YYsngi7Tua++WpiBR+D34k2oN
OpGj0Q3HiQPARL3mzSAjtU0pZk+iUgwakmSG8EWVF1dWHLTeXB+dXTsRR5WY3XL7
1/rOcH3N714hlT7FKP2mRcuXYkXbEfQAD9P6PZ8v0vgCkHU2UZbA31IIP7x4ELki
WkBeYreGrMq67dqr1UEiblp2gEFra8Ue4fNi2kRCXuFI6jRRz3fKUGfIj8wpv/nf
Ged40JrWvS2q88AUyO2fd6KcEEJC0XpJJjK/wMXiNnWqoE973w8kfqeF41/sLJF7
EznjbSH2cp5QpkGuD1vtbZMKfxOaNMtTAohQaKDyuAi6ihvnilyTO0UuWUx5G70q
COw3cv2UuYoQN0cp9FSR6fw1zI/V8jkAmrC76n25aqtt6fPigoyzX4MX5/ik3pzh
k6gpmkhUaDS0NMgqlwTD+TApFAGsSFE87xSpEcdUXay64MgnB/r3NmHZq5DOLK4f
gY9y70Y8Mpj25K3sdmWSk8PLXeTKHtgtEuxhbdczG/fq0DNGb0+ARkdrz7WosMlI
Hb+jr/ES5n4IL02e+LGLeQBFFRObHFoGK1XYt88/U8TYjHI2GnLX+SBDSaB8j2ir
+afWvj2y2yHqolKBsHmltIEKzrkrbfP4q3+taX6YxIGMMiCJRNMyiRqbErcamI8c
qszs15KcmCVZmEHGrbYAE6is+eXnc3RF2sbcQCg2+04LfTh2Q4fSpgyEUAkeTzpN
AOZXwLC7RkFgJFWYUsn8N5UeYctKqBUEgt8cuhvVvF35919ZkQtJz4ExRiYznPNV
+FxI5Ihp+6vtRmGWf6oAq1oU4Wbv7pUd0OzEH3+12AZBkIJjoyYc1Ua8tGfg9d6J
G1+dGY9IbSu6u3O0FArCIHLiPkwfZsui0/ez1FIv/ma/5d8VwUR5/3zqrFuSc79O
Bh7xlG6Wdc8tUkt9wY69fz642TZqfX4GQ4UIHci139ZyGahGC5HTRskS/J5LmLVg
nYfQp71b7G3UpJcLNlvQEkmIXPI/Z1WK23H/Sysg375f5ab8HXLrAJr9DzkTHU41
MUBEO5RIjr4pkxtqW523FTv2ODou94jCUKDpjE1ToJK7DxN7hURArZMKxQQpnQ4Y
ahH2tz5OFKpXmroZh/oI385BHgKKAgJHokzix2pklDjWizxDm61yxAllufe1dHRX
/hjy/DWsDE8rr/6ErWj1igdabMCdOibA4ANloQXo+hP9c+I9jqA1fsMkB/oJOwvX
e54fVqE9ULUUPJ2eiyIU+ZJ+GXCmbsnOz1dfIcxUx0pkL2YUXAOCt40q/psr7aDg
tqRnKOJqJyXvUj6INaoSM1v1CrUp8VZbMzNZBWQL/dpmYKmD9Ge80mlKXqeZ5nLQ
CdvhBUtsfKe1JN4O5Y6rYnxa+J0+KTpo85fXn9FiukNiC+QKqpB35q/dR2vg9ecT
JoqK0DCGWqGkTbtJaxlyElit4RLcfi9x3aqswhszoT+BHOu56gdV6LQZQXzK7GpU
Oz71TrER0gII8HYU4Karj71mNskh2uOjZv2MZ6AUNweKI/6Gdn0MUXJ2zNvaNlPF
wQ0dfcpDrrsHG/2QFTcITKVyx7Wyg+4RJY7IqZLvShFL9KsTFkDnM523aqbnk1OB
8jO+u1M4dK659FvzQK2hGx2X7HDeie24IAwYtGe/BrSUSRnmzXgvMdfC351wvCuj
nAgOyzGYc2yDXkotB7xhdpsp7hpbnGv9TuYX/gtt2me1zwPqwprzQAZPFUzzjLfU
y2gIHVeyRa7bnwGsN57xoarNJFFBZmsbt+/SCAJfUuXGzw1p6LGHLSIt5b3da2ur
U6QJrqSUPN3nZsnaBaFW5CX3GZdY7iZ2jpgeo7AmXeJtJ/QpJxVEUgYq/N+xA/Fi
/WDy+VbbgPyTyWfIC+RXwf/ZHiC9iUx/2kHdcIxIC+cS1NJ2FIotfazxuLM123n1
gE09P49s/IwTB1JlvCYNloRPQPgJdNCkqqLDThSb5bonl/X/h+HYFDmXsl7q2Vw8
SvOoQZKBuKrLTpTlLl2u9MXSu4txmA8MLP9FbGKg213Z65DPNi8Z1PgXEz+GCFc/
ZseGsl6ckjrAF3Z4x/P+taJcq346wlLaEnM54kRDKSxiA/cblsI6WibmA88lKNlm
7oXdGotdk2TWF6sDWYJGJRPVVQKP0fUj0TkyYjJ45G9S7sFkfAPfIC0uagfkNkqY
hsCwLD94lpMHlvvNfp3/HmUn2FubLjIe/Od8R3Kn7Dk84gKjKojQcbfILHsPcPwT
xE0D/12vUtRHviZwEv/7dtmKOTlN2ot5Is7CILEBUelnpd2AWh3Cng6euUPj9bGE
LMsYRaiU/AZvCUBd9Ofp/tB83bLq8OQKNr6/fQ5nY61rHp5CL3qH5kI+n8/VI+yU
POXLW+3dnbS0Un4Imy3txEsh7ZQWzcEGadyMkQsspijc3RDQsKDpzr+uTqToJF2X
SeqABYSy0gWiDOAkDIi/Mb0XvfEcGwiEEwPIN+FPnsjf5Kisx2cNMKKxnsWN68Li
OtdErLuKayb4kVQ/MntbjBTOx3zK2Nt2c3tedcx+/8bq18ekq8DtxGpBE+F+ITTN
+wKxA7vP8MQAWSycqF16t9yJ+o/x8xGrupOFqeUjUVRqyHmDLQQiq/9R29yJAeHp
aL7zUsdz/hNvfSZsOFe9hmKczYcRfNbz+9Z1sHzE4fmAaHuqJVObfwfIIsejMWW3
ega1qNFp5hgVFWMiojvNOMaz2lXPyEtVEbWCiMkAOKgTI1qjCBRd0jPXv3IhJPo4
OIb0xMrDKzEFK2MDXaeDlqf9siKVFVREEsVfGq2fLv5T5e96bBfGyz81b909GGky
afeVJ30ARHrcvEpAydkCiHy8IBAWo678SpeScSJzqmze+EkwGY02zh12t7DugPSE
9dJax06WqkO1A+FgtZhypCDSIUfazbDDGBymqnudOZgUFU+YQeRJSsSElVCH/NQ1
e2RVvtW3y/a39wKD2TOCh4bh4frxkdShvFHZM9NXflNO9K1Ov+/jmoGhBXkcUveg
ZRVChVnjt51rzlNUQ4L/Na/ApjY+xXfkN7aKIq9pPAOEVRz2pUMJnGE2vssFsoc5
Mf9pYX7yMehy58veCSfoTCqoG6/4QnSQfwLEWVjHIWYm8yyNEjVnRErsRvrywdDU
ES4E8RKrJ0JNz4PfbqQDf7gd1o0hZuL4jP5cUyu5khIq/9ILiVEsHRtG7u0bGQv4
K2uhmQPdOr5gABkGA57PIhyhlzEm5WaQ2tgATZriW1mGRev1975LJFjowQluP40c
/IDva3mNHYVuyhlWZLNadphfZ70pIjNYZwqsnAGm2MZ0yKaIF7jxWbSeoU07V/5N
x8SSWT4buD4r1oa3TrBkL+TEkjMQvH5B5gHsSkMf7+fYlTsuE1DzDHLE7tpw3Kfa
pB95WtoSaRvmg7D6aGadaGntp0mOn0LHFWXM8ixJ3S6izh46xcQXkC6Hv2pkHduC
D2MVxUFQfOdt8+uL2zDR/TTP0bU0S9Qfkuo9gWAdCrXfsPbGbawNDp4G+cm8l2/0
OErNZ0sEBgFk0H+ibjhGXCMFhF1JsZnRf2VjZx6FyCuMD1YuyNkPr+LOnqeiWrdM
zknJP/TLYUtWKV5PyPP1VmCpxwwMU/25q4sMYLvayO4F16BzNGzL8bf6XUOfCeOV
FboThCvprl6gZzDFPF8zTCvqiLFlgXKEoJNwz1onilm5qWxMMBLHBEG+ZZMXyo2+
SxFsTVnJPMolnWbzK57sOZUphHGaVXFryvNmoOQUZaRGXpWrkRuzwoqsGPzrQ0Mq
fmvhVOXoSeYyZ7uuTx3Gzs+FD/eOzsXtpceIRhkJaH4Y3N8cybmA8AEZmJhnMRBp
qSWbcUKD8wDfNn7/AU05ujZanWesn9mlLS+bK7cJcSd05IpvrImzxzkkqNkVqxzD
/X6ED6w9jgiz++RC9UddxA4SbbvIKr3j0f4nEs69gEOt0IYeCWEiKJ4YjpaGbiUJ
fxBZlwjC9mEJwfLaTVTqAIiBiPx3ZhXnizlgh26KECeuFHB5HZU4FlQf/cfdMbZp
ho50lyKNJs8YD3saLmR16B52DH8RZV4sToGoC1/K2qdAaxt4E/7CV+2tq9qC7MNg
QmmcaNEHl4cyMW/N9NC70JtR0C8bkSNxmfEwvGOXVgQup5yuqa91pn220Gb8/hGJ
iAlyT+KaipdgEMT0a+q4TG57xaCP+ncmqlC9KIm78mshTeJLXhpiNIuvRe2Vn3eO
3aHxsvKF5bQWAPurfRSoxWJVtH6iIRJzk7U+1rcCa81xjRn4OZ0s0p1WrCOXPje6
BZ6JuJhjIswqBUPIF7VHXswOM9wUH3+FXuQdWszYpt2+8Q9lFyi+mJUqOVZpuY0D
jxJjQydBvZBkcahF/Q9Y1hbCMyIVE9T9TF9LaGvOdJ9++7k+alKqVHHWDxb9dYx+
ZjPxlU6xFnblo+r1WPr349kXhYXwTSV1OBDouOuqectLHR/vq/phlepWsp1nFGkc
XNKxOJJHtFuchSaWSe0C3VsWg36RBEEaM0L8oNW6+JwKAMtbnqf3PGFTKp/4kAjS
Xle9L6srRXMaw8/YVnuqshghaLAjCAfW6G4QQbR6ZBVf064a20atkrhfiIumuLsV
IvRDvZoTjQNEwuF/zImhhUjuQCi/se/a5O3N2o5HX4d4QOFi1TFjryqL9t5pmcE7
W78QZmx0WL2OiVtyxlwnP+2bp7uV3sUZzfGxxbt2YeU8XVxAzJZX9BrB0GXHuvty
HuCVvQ3Nv3LKCGuIxACsAKUKok+G0FoT1wTsGytj0O/Q7Y9JMkDoqEhEIcVnUo0N
AW8u5BImLwhX3buyGfF/U98wMESRT+lYPP37/4GiB8+Yt0pwMeWDko5iZv0TM1D+
txAAxPw29ffNFCA9y9+6BSyXcPbHnhAKN/hdhsUL5+V1XUa20+X5pv2do1EQ8lnr
ES1NmozrpV8SF04u55Gf5t/+aWUG2Ff58n0dTpJRvvjoFNoHL7YPa+PrS0GgVMx1
ZX5723UoNwtldsVDxLaNSJBnRI6XLKflWzsiUOPPDThlvpVY+KR5rpY1lWX6aJlM
mAQmNK6bJm8wxraB7Vi+Wuwj4WQLhHC0CSGqcklNaUFAtF5E4RLYn0PmlHaZ9S/t
wKwmiOAXalCTwJ7v3+yNVDKroo/TF6n/iM+FwH5a7V9Jr5sblYx88naZ+PB31eMd
21x6+lyqE2d4FUlRfBQjfR1dpjGYiEcErRYL0HDFRWfniSDi0LFS/hMlD4sL+Ehi
R3P0qBSbyaDzGjFkaWZcDormZPjKZcJYpmWH5A1DYgMw9Jn8083BScZuG34Snlts
NQf4XtkynxYURU2re5D1lH7fxC8vZiJmpx+aQ9vC0rauzwJIiF8RxEurvQc+47uV
E39tjE7K1taTqz1M1K20vT6SDf0n8CaZbV57TNZyrCjlo9o32fmsIc4WSVgHnCH5
RxanDaRsWdKOEpKsaoo71RMlPbFHkEuaDERD11geC7FQUPqGHnOnxnWNW5JVCrQr
zgpQ0EyL+hzUs1dzKoYSIB8/c6vfxxP5g/h0QS3VDTVy3nYl7GTuGEptqvstMlbj
0BWMlmpF69WU2ULcdIOaFUEWosEu96xsNn3zjjC1MsHgFPHfOcejbovVoa7YAxga
tTMB2lu2/l5hKOeb23TVnv1kczsXOVqKNRIiy/GqNJUbuOmlhLUaQmJNX2fOqduH
1OKt5/T7yhtanQUPthHazCkUQO1eC9nlHsqfv1D9qNYUpcGYyiqBWvKGFsDL11Xa
SSxArwOQu5sMwGU8LlG6V+EgaGsQMNr9eJ9jhWbSGfb9gcKzPtZvxpBDh+KyBmkn
xPjTrVdNFyhKJAbPzTSWDBGSEopreEmXuYZC4vre9NMBOR+eY3/r4jNwiN6opM/o
t0d0eWjlDOl02u14E6T5UQM3N/9P+xBb0UEbz83pX2KfnDhSm397KvTtJPcPzaDo
d5yWGuYtNj1LR+iNmSLey7xWRHHP5yxD68CD/tapiWQkyw4VICcDIjEwZVd6LpMD
b5n/9NFnOHS5PweoMoCF2DaWLkzWZzUqFgk6C6frkWOWq97L9HqrEo5MINyP+Zod
EavefjTEOlQB6wikbpyD5enHkJM76lc4EqKMe+r3y57UHfrQipMn9RTUHnx4ct63
RloyDr81hNZtrWrbPCwfriukJ8pCmrt68ea80bbMHqCFYzw2fEfkqmUyIEbhbx+I
RH3LkF3IwDyBjSRqn0DsnnKhT09geeiMeBbKORIhOnyn7++DPM5aALSPoo+1EcBs
rfTntKWn0M6ngch7FtEhYO6Sw6a0+yGrNZ+VUd1na8Q58sy5FjX4+gtj+zyIMjfA
aRehauE9nz2F8lq1kMOUVwVUQjsyc4GbsQBLn09rwdsWTU+R/Cue4lq/wykNeQjT
Ff7mE/FcOlM23AAm5lYVwMNu/mettxKC4KIrRtA60F6Jcp1ofiDLxQ6xdx/NuiYq
HIvmiaA0+hbtysifGNuc8FcAEiEXEK6UnYuJjUYAUzs6bW6GkPFJuRxfe37VABRb
+DNn6xUs9ht9fugG7+KN/ZXWPAk9GWtXHxwVagRbiMjzVa8jA6G+UhiK0edoSiKX
iOHUpYVFZEVrqlLLieFlE6d8c1p68TOYJ0UU/NcGzT/GXwt+UGrPbdUlu3rahOLX
T2m5B/9Z6+MZ31DcPZHZMdnvAbYFzdQpH0+z8PKL59Pjw/ckRXJjk2FhMyPzs4LR
BkTxfmYbOzpzYRgF/E+jXDOfwmgn8zVhD/knjG1UAMbdxvVM0sGY0gjG7JA6FH53
fSgg63JD5FWhApkwNhijoQ+3v5nIlREWWWLmAfobjMCYPWzVLHfKyEoMi9Fa9IKN
OWqdrEzqMA0TMDDDuTlx0bmkNjDwP/q3wzgc879sNlBSX8HVVK8Ttl7T6+VSVuEn
webKagZeoUEMW0DUbBpXojcl6za7xIh+H2Q5Jzt5PlRQFSbbZpQ8hXuSwJCPA9fZ
Hg1TpTFLqJnPtBzbTuqWWavgS2OXBGsKerJI0SW/ppMhmdrCuEo07vpWuhLxYXdj
q6weBhOqw1ZYoYxnnM6Cpg5AnXU1JO8pQuh0V7J/2Cq9t9AuhW2aS0s5unUssX8Y
RnkqOBq3Y6mB90UvnrntFp2+ze8p08dmS4Kw0DIpqDAemTnJIzKMrFU8veZZkclm
QGkO6pU0hJ+1nDgLAX3G/i65Yan1Mdz9Xqydo944jATLv7Qe7QMhE/Rc3R5Jdt1H
D57QYV/3+NWP6QX61chSHoAQXHHX8UN+wQfcLamcp/HbVpKPJQ42FRA6LczQCYSj
No1aZGziqR/CgWQKP5yPllJPaRO7qbJJVaARu+JRFJRrsQJbEiOsPgwNV0lUosVv
/SXRvl0pCzDO03257X/SYN8a7flzljxxNYrOslXgKVZMqYY3HoHl6HOcE1HixL/G
xHDJDn3rueHrVsCzn8DXaG5rgwYu+N2VbRm4VF9n4iQgP5ueXB8DeVgyujGXGD1E
B+IHKZksxcNhZhOa7DUgGdwJg2oA6YpmcR8oL9Li1KCCxg6XuzWYRInm0ofmJkMI
iTvSJ/bit1vSz7AS7XRzoFPAHslIYiqQpDQ1GI9eli9OCnclCLKiLEdz4Tk3EPpV
wMIbEhQSa9Dfmf3QfQTqyVOGnRF252KMSnqaI4dSytjA2Kq7bq+aHd6gm8G0o00A
ptZ13xm6im2zz1f4vjwhP4RdD+rOZzbj0BkaztcuB281BSVDc4YXBgeWHwb4oYeg
HXBf68SlZTKEbUYk6xpHKLV9KiDorqNhhlvbcqKTXGpAAjK7EeH0LoNAz9QXM7bH
hcuJUq4B9Tzw1aUDRxv+93PVX1uGgjOV7Ta1R7VJy+o3LivhpBeTH+zJtkWrbmHB
b9Vi23a0fKgnAIKSGoLc37/BnmbD0HsaDkr51ryRNQMM9IweBCghBrjL7lwAcrCo
2YRIhJ+EUQpmNib7COfoRaIaMTnXoZmU//M9MDroQd2VQREw30RPymaCxAyTt36Z
Zvt5Kw4sPM0wYjHIMuHa7oCGBY/drrzqgp9yYFDMN+pH+ADwyfXq2hP4GXeUXL/c
DeU+7e92DusvzW/bxapCT8kocftranhPbVsjKTl0RiwhIUkWSLEUvvfI1S7dhz7F
NKIKvCB/LGUFzl6hktDHkPP6eAdfuOiI1aoG2kgNSx2wMjteTAuiHsvUbRHA7OR8
ylwC6on5/IJ4HMxlzoj6Ajgdpi6MCgDCl4Z42KKmq5RGBe22b0Dl4mWLxxL1YbAR
JICVuGm5544T+ykVna/lMtLCKEPt1DIt8e+WElm6MnIMq340wZZexWGCu6bzsP7B
f8X+ufNWoyOGiz6P6mx3KCs+Vr+zcTL56G37ShoPU12pq8lvKeR8XTKhW1xEMFw8
oS1rUAVNj8p2HMHTS1GDyHAyLgq79qaAReIvsbbY/VrsJBQUD6F2XX65s3bY7m45
+kdAdQKUGV1Y0vUjHXpZyVF9J0uUB1a1sIKxYMAsWt0+weVXZ/uU4F+PCoO/W2l5
Yywv+H5TYQkPHCp3+J1rvAZLrNJikYTy+TBagYQVBDVO2BmBEew3YnzjV/4tpgFw
M+F7bwxHNrHv4AnR+O+/uE0RnEOx+rmcQcDU5K2azb0kNXtWY/4rrVt+vvmIifbF
D1dY1ZxEYn78mfn56ypbUwcEoMeZPJvkQNX89K62HZ7PFfwUQHappH2/U0jdi51N
01o8S/7v1wblSUqpe7fHiCVZVVW7YDbJ4Ea8XMZtHw2/MgXhC/PChY9NNzB6A1TG
X0LpRVmJ/zFQf/6KsKW/cJRQgp6sQt8OhgX/oB9eHdLJLW4a+HdV5D8mAObv9zva
ZIsGwMtZGVGvCfASY3ea1BJo37aBajnhaH7yaapAaN0ce4bU6nv+d8a67vfllaxN
8JCGJaBWfbyMDLkPom5W81GpXUZUlDJP/95KW4Am4oaXo3fTUgW5uUvBcE2iurQc
yPxxbdJOoHxcrN8ATb95UNDNccj+ikrC4HBb8X4w6DGIwiDmdjqXdwcRpjwMuooK
QPOV81nWyFJ+EOKNW9qcPMfqw7QW/i4T5oUgb7HCBNfSu/7ivuGoiGA2VeuC18S5
hgCRCad6K5QYOolAblBpJ6l3a+iN6RR2WW4VHCF3qeD2JYAURJwB2HGXDr1h5hFr
D+4/CSYzpulF1XfVHebBWIgYImmtTvaoA6k0DkJ3sGcPjSbjU1Q7y2spEUXWqoJ7
KNCVPz6rw1VX0qm75bRrNoqjBik4gnQaINz5z6oKrfyNrulqxSUKfrXFpH5giV9f
5cql0DqoUT4WNV3FNT8UoDzCQ8caSwf6qO3Lf/XzStCQXKjnmqgUwf1iFjyVHM+7
haRJHBbxyr1+ddBF8/y9zDHBQQJfdLQGOB1M1vSHmx3mT5bxLRq92QEzG0NjCcOK
qeU3LyyMmv93uWWos8IqlPjydCDX65dQAjKCZKOBYu072UHB1mIB2GooyzjKXpLs
4WSJ+I/R8j0BvSodqL/hElgVZCXz2pySSE7S1wctJ9TxOZHgmItZa6T+pXKTxsDs
Yig52L4d9GdCWeQyi1+cI0PCGQ2btLEh2EVgdPhOhGkt7bltJPSxnSrh5HVasFNm
dBIKR03tzwNVyJyKMnYfc5UjcWrhDXkQVn8QQGZpM0xzX0XmksXNN2KaR6EZeES3
d+dupKEyCVWW8zo7cKpxbEb9NOa1TdgypO9kEwVDF0i8M83YBeSrdEFnmxqhlMmy
fAW8NLFRIxsuZ9HhzjIVJeSXqs36Ca2ZAxgyhkxUyMdXnzergRm9GQlogMv5GfnT
cs6FPfssch14cY1R3h5lN0TAeUHqGGn4tOaBGlpksOdPgp6c3Q+xb3leaRtwzX6C
V1nas3T5v/WHa/BQGsU8sJgM0M/GAXAGK3M2iiIciVPNrFM4KPj/ttNpgUR6U7cn
/FcLn7hmE+UNP5YZGytFdcAEwGrT5FRBbcO7abjy1yqyMqhegjI/qh/PTeZlaTIX
Y2tZUVVY3YposRQnxnmxYr+U9+ruC6agKJ9GO8fZzmJFHX+OmZ2iboHvHX1uXlAk
09y6+V8cGTRgKctgC/d8VdIlSrMrWooppFS5hr9LiYEFluUoeDC8rKlvhg//a8UG
4sjMQXBYgAaEnIWzEvHcWbWg2aWfQm3XQ3BOmof1cEqXzFS82pTe1rtSOOtJdPyK
goWFnW22Y4C7r3gSEFPvSqC+e0DEjOrXZAzJpJNirwyX/DmT62G/yYOm8SQuDze+
5eauSACJvLXoefEeOaFirGq5TPddzJTUe6xBqTbgPVVU3y7wxqws7rmDoPk3DZi5
N7GYnc9r9J1Q8npmg2vvZRk/Z2aLfTTmYqqr2OIBswrIlJNTI9LflM9UhjF4N9qv
BaXHZ+xcsmTlzN0BFZdlQdGg8+2IlYCWatELqZPjHhzxkaTGWf86d948LUbh77ff
LG9LAkI8Wsn9bLh9nty5NjP6NpUYgcFc9kCTnLuqo476zCO/CdXlDaZeq0T3VLrS
uKB1YNnuoXhvtr2R1ElfHJ1rt8d83v8Y/d4W+BcEGu7IV+c3PtVoz4dCsaO+DujU

//pragma protect end_data_block
//pragma protect digest_block
gZSRnRR7lFlrRI+eN0GztLTkZto=
//pragma protect end_digest_block
//pragma protect end_protected
