// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
UU+MDLwAz41g46ugBLM+FJ+XIzpTbHRYTJVwnTPkUKakhm/dmdc4rpIef/eykWf2
VprkgwqhqipLlh5txKO81LWxUHoyYTn8c2vn767DVb5+X6PWE63e+WbC2fqkgEZA
YKSHp6kopElEB+p1boqMcFI5ioLtVFS1ifY6LrcQr3Y=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 99808 )
`pragma protect data_block
g09Wg7bR9RbvOGYqlCaGOEzJo/34SL67b9svC3fsv58BLGd+pxOvh+oYeCwuYWdj
CqI+Qn7LikbVzo1RgRekQcn4iqeEiIet0qkmSKimNCL2DuQfjP0f4pKGl3fbfEVd
pEn/idebLpATBAwgiePARRGGcGo3QzdhIsYlFjqjOBhQutfkcFSB6y7+MDZqxYA3
J46uZK1QCtDHYR/xzV/+ZNDYswhV3EDNW+iiTWJpU+4wl7Q0oHyFIl4YbzjrjmJL
MW1e0mNvCnEvwxnreKUzwctSpDRsoYNPuy0EOzLoerjEFLDYXJDb5H++HAVj96tu
mAuiLGEJPCA0IP21nx9G4rN8nIuBqIRTUu3MN7uMwhsk+/QCcTERapv/tGL3fwMX
lyCnLEspNv8HwJLCjELfb8Ivf0JbMPrcPO1UU5dja4VVDZiJPYDUXZfk3BFww414
0LLI1lWGJnvLtwUphUGtqlmPnmXXm6expudTJhFawcEsEudIBNl08PPhh35xMWaH
hEtuxqHXIxJLwjwNh8aiCO7Xw5Z3MLK9Gn894iIPqodXPeqjSy9VFCyFNY+M5R54
9KbJ9ZgEQaTM4sW3oV7OHh9yPL1pv07OfBOGmzPzu9R9hi0IICfJW4t+fxLfT+jh
WV/TQkQI+BRP4MUidPT2BHS+1wAGC5b++yk7PL3sn5O0qI9HoAJGnn98KLjouqpZ
01zDvDwUq9xQSjRN9xTvFKpiC2b+hI6jCX/45sFdzF9laYCyTNQn0m0s6Uc5/yXS
rLIZNyvcLuzptgG6GyKDkMtUtP1I37OgpWAjXab6U77Hht7T3PAscCYPsaApyx60
TayFIHBTi538g41mIIzmtxt/6maUqtM9YpnIg0DaROYkQam27OIJWNy6+KRtKqSy
0puUWgKeWth+YNtFldH2EKJZdskx646s6xR0XCOX/kXonFvGUqyKHhMAGFQMMNuL
dybI+NLQeVnsmgg/HdWBwfVWT9VqyX7xhESACvZNrSQprabA22geJ9fBGQBDtleP
qJ+Ii0er88A3FiNm4DVFwkmLmnKGT20uV4+Zv7Bycxe/VXNLwGD+MdLh4i+YPD7g
MMQ2rDQYPI43G1UUvoI+wXftjG46DnuynmLiaCF2fyeknCMxbkvvMzbo/0zuvp1t
dW/NkGJ0wdM4hcpyNQ7b3dQsDzCYb4AfflGsO4ws25lb4kFW5cJTPaojNp06H+7U
lJcgeRMoKdsbDMtpzLXT/LN9fCfdwkHfR3X4u5GPkUzpnNaDXEPtNTcDG2/5YCFR
/JsjZJDkAygoy+NXxMoxEqu1WJhe60Be12fUhHMfHtSABKBETRvjjZ7/Qiw62u3i
Jl1FQZuewA2zkaVnFOCseNpFOVqJciJZrhCmezeqUAIf0U8VqlcMMkNlFdgKfZs1
ikG59BYeFZjSIXpbBl0Fxm58Fjjk+DzwwkOcGUrz36AXV/geYQRXxnmzlRM9sgbP
p6CxokIqzQg9zRrrNvpkBJN8ZMrvqgyzomc6ZaQd2vdr1616a7RJEbSn58lDV2tI
wsauqHDMSYlX2QRiJB+ej9siewmANtqzmLP1KUngHiqMTr7NIsEy3FxpaE/ZtV6k
F94airTAV7HFFlbTb3V8zf5G4mvM97cSY58qiDDr3+cGGKAtNGo4CoQajEN5Jx67
K6RUVexlnWa1ch1S+tpwL7TlvxthMptgZDwWP1sZ1V+Ecn0nZN0BN8gCgs6CJMg5
VWZWDKYG/zsMcNpd4ii9XEWXXpxhXkRrQ65Rf2NSa3AEaflClJCadfHAhemZwdrd
Clwa99Xd0kRooaa8sxZQcyhlJtq1PIXD4Nmo3j6TuvrgxopccTJQXG2hLl3tgA9a
+EqokBNbzZ1tZ9z9wQbbl7nBKHVYvgzLf7qpDq1HM1T/FySEpX41MNxIosFY2NeF
GR7gblDXBQe7Dij2bOzDR0iFtJTiOkQwPhIK2BBbpagacSohYWiXdkK7yz3yDxt8
1vaG4ohxh/u7kqpyM7nUizWgjFmQFUplZSADrNVMjTx/rFLQfoVfHsZ1eH5f3zyG
kTzaWGkNn9m5GPF0YjcaE3agsVC28gnA4mwHJIngTu+ADlLuT2s6AE/gKDuLze8T
WppsZDqa7V6W9bggdwVX5CrAFdpQv/98Mlzg+O5MSFi2nFd+qxu7ffa4o7pV0ujI
E4yjrylLzw8BZ3Dnwyz9Eej5bMTGdwTlhoC5YE5/8nNvuGM2sIXtPa3rCQ5OOMD0
9Et1CVCdIQoCHlp1xAmm7arPuZ0DLzdXb335t+hdoDm7oiwIfAQVwBJdfInhp9Er
dzFGPFuOYVrOWK4OdgEvtY0f5K1gkt2racz+sDxQK2HC9j4XsoRBcCptIxafBlWC
xlnfZmXALiYpFqVtpEdm0T1KYwhSl4Y9YOcXS54qiOzdAO6Kd5FOxPhCYgbPnus1
JnaBUCJO8qmc1m780QAc58fuoFO6m+UpoPMbYIOAG2h14XAJ8kTqTRyIw+IJ7NQx
TnPpQtSh0equDVLkL+UrqXP4ZEmn8w9T2eck5hVWKb+wPIejzt3KpedL/bnGlyvd
0SIYkN+hKq7Y3GBPQCa2DCHgCOZsFWOM5tmGBhljp1GGfrf1KVd3PeWL/wcO50Zf
13n2XeHI5xr3iV6Iwj9Vyjlw+mfrIFJY+AQr7DCL5YPXzMD3xed9KEO5IPKvarO0
CAorfuINqDxfGwqcJ2fcgN4+qhNfKoZ4PAAGETx2fdBtiM5Ta6dXeYnHK5j2k5Rb
eReC+m0PCgvtA2TqngFpJ8E7h7eTSJSME8dyem7NmFbieYNPOzdQq4S52VqgSSKf
6KDNjO4nxLVYbp2+nAjWM/VwgPuqOaYhLHsFZzlLA5iEMgasNlo0qxwtTfvukfu8
pXhCkYdgNrqRxwkEfbeyCnAvk+3ZcGJl8l0KUXCD0NkQGLnIcTPZeSbwfA9B5l2N
W341yw/PD++O9sxYAf+CK+0C99Kkw8PnZ67WvG2fUV69L6cZ0m47nza2yL3xe3ez
o8lyNcLb6sQq3TAXKxkAx/slHpHm4nWmwcNAcGzLc6PjTQ8q8yD17Fzb95cXKTgH
zIfe2cMtEiUEpXYgCYUqxUuFA72uJ+REQuCiQf3KUKVYygigIWpDVbkJNUt/ac6N
9Val+IQKW6KpFWO0cEPv+1sF6TxvFHyuhO9mggydOPo9o1wr+0/9RBRYSLrJQKV4
XzjUPe+LrdoZdmhyKTdigSYiCFkLWpXhAAF2Qb21tL2T69xcPJhB55EVDyHbb8U0
k1uGYLNc30l9M2fxz91dOg5rpTOZEP5zxgVSwjRxBd2c03Bh4Cvl+eotiZNwRlFA
CcSu9WNsaR2oCHi0KpnDxACvSB7m+caVrcHIKlvUB7Lfva+IYt9RTgbMf54ecAyf
4gaJAk0RCqrGMH3xi+xOQN+ayEBexdX5/pcjoiQucKAuVe/qcTJhP007yU3Uenkc
Obd/SjHQePEgOLLOLxwjJb2cZ1v8JHDAZkB319OBnj3j+/tl9naz1azZroowzGPA
esi9YtytFfwFUDB6C/jUcXsVLRgpAdbXxv+7Cn3ReT3MV853Qui1BoYfWePhWlrq
CFf3NkVssw8hBAxB0oH+YxpTKkUEKoP/bYYVZdQZ/gh+B277Z9i/vXh8z+9YI7g7
rcXw+TrWCJZIfC2SOcGlncBbaSzbv78H2nyhxeA/xVUocNQW/7bBR4nFwUlgtJgK
4sXjPBnHroTuU5FdvaIe1QmYk/7qYiEeaPJe/u56wMspKwOr/ObNhBYDqyKY+yRj
Kh3v9AEtKBfFXYFYfH7Vjd2qNkVHwcR5B9WjgKgMMYwPc+bsu2ED3SRU4K61v7Lr
EHFT+CnyHEMj/KwJVQaa1kIcjWhndtvjsCgL5rGbTluXyY/mi1MYz/hn8dZMyfet
YlmsaLuiw7+JR576KJa80tMstrnk8x4CU4RIoqZ+REG3O8tnoPgXhxasNsm0qWzT
3jNBi+ZBnJMvgpiyvPcE3ZBDzOs59GsUTf5vrlT9jUQWgCM55OGYIcF7izPliDAp
kwobFunlwtTL8B38ZLvigos1qWm8z8SJKl/4k7XdM+KxtXBmvzk0ROMbv7YYhlj9
UgNohVwdia0v+qKB4GRb1/AgvJPWUpeor2DhlqO9KUNBqYNFBrkTswcU9hIyraH8
SVInvsmmFk8Z6d8u+b4Viuqk7vL4kCp/a6WLpRv2iTNOL/NMWlYsFu/E6mzYycmZ
KCN7VbCcc69R5xGY/a4wUNnob7DpIzEjxUXYdl4hwY7ZFUV3t/EHFax9BzUD5mEU
cLnkMiuJOM7jGCK4TWYPQ/JBTbFWnVGP/UCAVaK+p+1KN5RWy0BuncLi/AA8tx/F
/XEtq6auVxujnhyDjZOsYV7x8VadTekSlauLW1puggUXDFt74Ul8cjHm2ASyjqkM
vW8rIgNpLECCA0fhO9x4WIRWSAGjAJPNulMj3wRjhptzNfdGXRl9cHj+UNgqB67/
QKKWqxQZ7rGwA3vq5MmcDPtEf4UsF7EhNlOivnT7lg0W4GLWJkSVJauFGRBubqF9
nQypTDxbHzW3pEAn+fH3D953O22Mc91+v9tXp3iH59mM2frKIABy3e/PRsMjV5MT
EfeQtIgKMJaE4RBY3LrXdBGUo2L++eZfMCsKNUPquQUZ+g/FMpBuYAcIVWizuqgV
Wj15Ud9mPj6sE9CV/PzH6QKE8w7/irJF9TkzsVIRLq4oVQh/jTxdEjBUWS0/1ITj
fqRK/YNaziV0ED2XTUNJSwYtEaksWsDRgtsWXGeMGce7pNe78R2QMMQNxnwL/AJ8
LWx0qxv60b+zhSrnkKZFQmM82UePt7E7PKeusIQD+VwZ7n3PyrMaSUnr9yGtR10A
p/0LyItkVMPwLh9xB07J/6iX/m8k540w2mM+8mzHFAZyImOJofjpRIecsg7IZgVe
8p/+ENiI6TCuSrZYUg+Dhlqa5QStnurPFp/fusrfixIeqJGJO8imcwu+2afVphY6
t6rCgmwIKOwgbH/xriJ+kM7BQZiy5+3P25fTfo/9hn9gpPicVjVvLjU/iBZBFke8
aAc3tjIKpRMaTMike+3NOvm4VHjA6tK6CqrF3WS87LtiXA/llIvzbeS1cAko722X
D44SA+Ki+BYCD6SItSSQFRLXWdbYogaDOzK3MWVgMacv6LwucmMsCZhjXr4Z5D13
4PZo4j71H6WlyZL7aozB/wxCPklNPOw1VeRwCmd4Io1ZJFskDS0M2crNKwer0QK/
/Gu1HP3vKkTaOsC15daDoLjzZbsgkmND2kEs0rIl6bNP+zZslZ4HTaxSZL9Q7RCP
HLolk3chG4zSbhxVAHy8Bo443xp+v9y+KIH6zM+YSPzZG5/hah2wzpVbeLhtzc48
dVSPlJ9YyEs7TWTD7Nq0539NaC98T2vl3djAtKduqeMu81m4oJOLT4P0DATh998r
XKhX3YdG3p2TIYCvyb4kbqUaANdTPAJUUh4OGJL0Ozh9fjXOHtdZ9QalI4eWrzpY
D2cQQdffCG34hhPfLtRqQrJYbQg2qY1FzMo3e7Smns6jTK1650VH/k/o7fjcn/U2
4sjyC6kNvM5Pz0Ro1cOpGM0OpMtjDnlZi/XBVRDKaPKzpw8XwZrVS3ldbesOB49a
6DyTzglHTw7Fmtahvxgokb6asmAtlVDScX5s6OEb4iefvXq2vyhX+E039Cklbuvd
4zYXfJngHvDBs1eqpYo9y5123SA2qMfoot6NYr9bia5lOEaCSu6T2+woxBdHg4ik
tCrQciIThpSwxMxiuSco+Utyz7Az8DvTtdhOa+BqGZpisiOMzNlZNWmglP1rvJ8y
BBbLaZz96a2IlkUFnokpsMaPTs3NwDGTTySe0Te6LXLsrD1N2m9OZlA30v+WQXE1
n9yzop85QG/PB6HnZnBMsAS5qiYqaz95Dl4Xng9FoYyFQ1z1xJSxsKFSivWuS/p/
F5wzISRpLf50B+5LUfn4cve3DZRC5hYQqDsjnjgfvRzjYjfD0m7Mf3Jp/MuktzHK
mGdL9n+GSVcvXQ6yEv06m5gq3wyr83eqf9GErMWfYjYKvcdTJhJ7qJhyePt5hU0w
ebtyrVLioS4fwZeFwRo9hIQTN5e/hSZgtYYIrCLjc80NHigpEbQRZBwMIb6PlMJw
5J4MALgHDLhYNh3mrkqjQ9qvVicqgS8YTfyW93Yi1ySeQUW0BNcCmN/VJxzkpnT0
qMOXVCua4bN6+cAoS7g4j3kzE9ahEDslBXu15GeNEHO8YWyb9IpgTIDEDo2dDTQ6
bo7Q5iZ42y1tQhaWGVXCXWycCSYqVUo0s3EvNtEA8DBN11etREM5NQIPhXjKymyV
1wSZuF0BV7yemCI4C3uotOFAeahb1pg2UUHbjukUAfFDEk4OSySP4Dv9a5Z9nQBd
VcxlI7FQrqsvSoBfyNGywUN6rGWqzcRdHbrcuQqxKy+c1fXsfAJBf1LV1yUTA1KI
8ZvAr5bBxwrszFYVgPM578WH/GTY2HWkieKE2FfPDrZ2F/VksV1uTSiPyUL7aVNx
rWlVWCQMlwvQMwzy8uLcxn64nBftwzS/bBLqfUCNd8FNCPX0UtiyJTIA6mVkDy42
m4IEeMkmb3pzFewHLyLWo69LhVLZfmf26uMR7z0pCLpGU91Jq6Ya0xCxkJctB16s
eiv+M6DIhKC6yVaYjwRPRsh9kxThq+KPGNXdimaD0Mo7Gt4OJZTgYlC12MQAxkCS
qzahL7hHUS06iB/FG9aIlejsHy/7V4e9Xya6ePqJiu3HbO1ELc/diXqiJguYJ0ws
eU28quQ2FAmitEBntMWIeQhOrBKSCIMdot2WE7n7UtdqhczS7kjAs6CW4wdV0Md8
PCZTzQCrYlP5nrmCVbyUVgjounM0vfjHks3XnoSB2bcRyvAFSKYj/uYoNOeOD2Dx
VRPmaWzXLCncQI0w94hgsCn+C+Y2U3YZ8/M1+RYHZIa8Qk58UfZSTKfk2GgGqrBr
KD4Q0SHiO2N311ymIahuA9PWUpASQ+66IbyZr+in/7ixepYvnZAtOnS4AjRUQGfL
qmta5RsDrfVZiw64ex0o+QVbGHWRhP3MyV36TDPSBNewiN5UBSf9+Cp5aDzgL8MG
UQ9xnS4d5Xd6zh3eSG3TdPEwLqukf2kvytZec/Gzg0kn7IGJIlu9MstJVXx+S/2c
arOD2AVsdNjhDg/1M5RUb39qlsHvBYAiW1ABLSV3o3cLTzK28EwuqGT+7EJbY4ro
RlIbRYmfz/rTNG8Rgsg908tLC5vEwCA0j5OSw+3jU4P3SzHbQl6gH1LZyGIkArW6
Hel1ti33pzerzsZHe4BOlti7z9UdxG/Y1CxK4dgqaJeyfuEE/7AzLI08wDH9hutz
K0GMU2PhB4BSHD7qQrucrON8f1fuVt3a+09Mny3RYCRw0PITyDTWbytLCTT1bzQF
Fp6tNubDLYZWVASwLAAxntOo3UBwCUYVKFNJ+HftwpmVmLlo3AvkTIJLsB33j/+y
2ra9KU2cA1f6EzY7cy2L5n4gCEZoewcGCsPOFvmdfXolz+Rzo2Dn1A9Zh7Gp+y6+
j0VQYlmcuWpsley51SCNY/IfArd8AFdzqGi8flzfHQTWj7KdvssOWZC1/heUY/x0
0wc0wOJoSy23iY2tl576irklTDwjVGaksXQI/KTkqxdAR59esKpaKQXQ1cKq7YQG
svUPDpK9nHOXoWlGLGAAKkwoqahMnbpphXqFC/Q2vN50LXiAOUdR4F10NifPlS7n
cjp0WC2Smi5mnhjHkCHj04v7icAOn4cdy6KB3Li2jbkvmSM/rxkZST9SfLDVa0Bf
21Qt0cgattDZyAo2O9O+AK1jlH/tVsOHgJNscKPiBFacVUtPTOPaRCHxUnHc2ZqP
YNkVFLNvobO/nYlT5pDGtmCgcpGfuOf1FOJShzbvYVOhVIBnrIXAXUYAz8qe4Y9/
DKlOivUlIQ/opWyll1xrGfku2G8MYQnWk02OwiIcaKHIz8v6HsWQ1Hp027bXFSXK
n7n8iNNPTU5OwgbWmKQPZnvQIoyFE8FRstYHzVwnAM/TKPdsVzKRi93cXlpMrZww
lDKAzfKKQl4m9hC8a5UDp6RhQZG2LqhxlTz6m+D7TcAxK7rz8+uTnuG3vXMqsd5A
Pzic+GshF2CmIHR9tyDpUmHON06duE3f6trQZa/pg+Rm3u8yuTr/BGIJssDm060I
q4QuceyAItv8QHDBAvgDKBn+7BkldHGxsmUf6J8zcTmHa3W8Fc9qE0d4ORdmnWXB
nwAWmWmF+SCmPnS6mi2OBW7bDNjPKgH0hgg+/e5bZr/yRfm78M19qPTot9Wt/R2/
aXdvWkeL6i/odUbUA4BxdRQ6LNyCox4NaXCHk8yVfKJvUlL34uRiZ0yyXZzKtMhx
ALJfoycX/rFB7mmQqOECqi4+jIuHWP5FziqnYAxxY5T7JRy1+HQPcXLYxvMpMoc4
1DCnu2BCVeMoxnIDeSflbAf82Ar87p9B067DdnPrgnfIe63BftI+vfdo/sumb2l4
5+q7YzHo97zV+0A2/TWqyPs/xKbnkG2x2dtio2XaVgD40IifhDOaCUMt9KQUFlaH
NMVTFFx8q7/K7+YdO+U2gcEvk3YdxzVfI/S+fVvKRAZavJo2140NCFNqrHlIOCf3
BYefe6PuuOnhgTTqyD/kSBaJ//BnLqutuszZMoz+e1NSYd7pNGgxo0ZoFNxsNhTk
tkl+cd7NPaY/f7/MB69P1ZSsQBGY8dY7PaeBELHxPQmn2ar2N8R67ZfmqF+APTli
DKvUZWltSpW01KiUsXrq6MxoXWEG41EiqPj4PYsEsJJ3N6NAJ3SDQ39+7ZuT7CtB
bL4dry8f1Uc/VQrmCSVP9ALOHTvimOlOHF7oZH35wqbEtnpunaq9gEwgs+PKbyyb
zdjos5CYojec0G/OVgbWi1UYeLIJTlmsYawAsJapvS2klH/RuHTv/BCL+gC/GxnB
Nvpas0zsaYjmqo/dEYLGmvjGkhOifg0rGg4yXjg+wi0/ASZg03JFqnja7bCsi54B
/7G0M3ww/AXknwZFWuW2UmDPilqxNWC1TUsfn5T3murMcoi1NljCBfz2yUS9uCdR
zkq2Cw/wzWpmYZc8lt2Mb+H28N5mH3kmPCK69QfxDj5aYqw8SLhzUCE3LFKBC98K
fKysL5rVOPsEpgQvxGIaKWCJ43VmtdEaDvpCdoUx7UkP3+hVW275odHn3dhkkSd2
UNBjFp3AMYT6TG3G1M1vKyb+smBGUJJnJsSfFJUk1Wa8pWhKIAfJFHLq8TgjZdSq
73vwvxLY6w9k9XTKVCaabW00gdbDlb+Vewx28c25QBoUjmjaMh7xThxWv92C2l8H
lQ740fYxSytD/Za+VTZHtg9Oa30OHq6uae9bYs3CEhHC7EdfXPeBZwPkFRo6gV1z
rcBxEUa35hkeFbXEfQQBy7qDeSNFsFKN/2a+r50oJddclgWvY6eJeQcwDYc9fc+F
8XcUmJ2CvIAi4jD0oEi5ajn9O7gv8BHqAKpP5XjYiiccqjHUSE9n4nfb18IlAuHl
pFBlB83C5/m9zyfHUk1OhOQcGceYbmWycHglaaI/di+xJuoym7/3T2+cK3Kwu1N5
gLUWg/cWevVeJHSTwMMxb8cEdgCsRiV4QjEDG8WjrqF1/D2FqqR5UxZ/QDghfrqm
II7CgoA6fytD83vuL+WO+X8/PXs2qPXI8zPIWM6Vr+/tJpjZHb26Y143kD0PmhsO
7DEHVxpnwTrtFiJXRoeAN84oPTBMSHiVkCMF78cucwRifjgZtcqkVdp/rFHScRfR
Y3aNRCAJ1Ul9E4sq8JqGQFFScvZKEzOTKcSw6RwkqqwzjK1W9SgqCFMx03fVFIlT
i9TNbqv9F4PhT9hMqQw8QRyMLgpBvOf5iU0bAR1ne6YSAQvZVty3Z2ylronKSesF
X4nz6SY0cH1jMlt998sAA2+O2/3nVGVMZDLRSMH28PPG6ix2O2VDcCjRWrYgbCQH
wsxJjRVazlRIjznReCr0uJVDCIg1SlLTcx3GsYmVAuVTWCRHcrnQ/5Ktf+5dKAFQ
J/rrIWwLPz4hQM/zkWyIYICvHDLmpec7uLaTxA7r7lwjZ2tmuQdT6W6BBcNAba17
5Xe1ScCQpqN3RwroYVcHUbcTpGZhbkRqb+oQ5tAj5Sr5RugGYiBfJ4B/LbONVLgh
wQ7oFepNg7dJr0p6wIIHNcoxulQqMEwYsWWJiwHVgOPbmP9iK1D6+v7xtl2ac/r/
IHKC/vYLlEcl8qI/rCq6kNaySwLGS3dyHHsB/SsP4IVR2AyP6HdXHth1bnjs9SHX
eAubyci1VMCBQwGrqt/2o2e/hsQi51sjsRtG2kYGGWsd+IWM29HSCn8UJafojYlX
A7Z8fXvG6OeHgREasey5PwxPvcWrBp8ozRLJI4+czif+Rmges0vufXtRJsaUeoTK
mosP9wN4NO5T5T8W2ChJ4lie3O8jrA11gaMoMe3GU8/J8Gd+ah1H2Mmm0cuK3HSG
lwo2ea9y7k6A1RxdCpTuk9Wu6z9MQQYBXKTqKU0a0q1LCDczQH3lM9Bjqoq3Yvjv
fRhnbW3pomhXKzm077PKe4nc+vLtibmSXZVnhcKNhu+YIz7iH39KQQgHH0Ac088b
pu7UAsdne+5ciRfmBtWYdbzs56BTlrqtYeWP6EiJZLJJrR4sPAFf9/bSstdpKlVl
0skbqhYAuD9JAMDCnMRdbFe0vQ2KbGTIxsitMekqqAZmpOdCbM1iKo2YFitj/Ojk
4QYvuGt0wUdH2XHVKDfEUfN3i9DXg9iq6vPgzfk1MJmmmc6JC4TRDVLBd8gWrQrP
XF5/CmyM353Jm0+zvYhVXkNAvLQSbnk7KzWxVJbHYf92GHSmR4b1sJo0oHjnV29Y
bbpDHXmkcECx1IUEYzxEzrtP7hqTBeGQsmFAtFPKzpoq2DOH8s60WqvEnoRBberC
2ivklGSmFHgOJ5iJPE+OalXoy5ER/pYjlvWWGQzif9/FZPyuG4+Xwii7SyK/GUCy
NGXNk8a5ixwmf78DP3vYKMrzszdJpGUsSQNRo/WoThmYfWYWsxCiCh/NvRlFTPGb
+A/mydyAhrtMnCL9CG1QLSlCNlehNmx2VgRRtbjaLOYZu3/xvhe8sanUyHo5DEge
WRGJDqjCxWrnR676EoJm0sjWMSMKBORpEo+CRLyrbMrwswMaBjHFAEBurLwzu7jS
f+JkhknjYii+G928ncNk8rMJTreDlWGTbtG4jLw6d1Cz+24s+yfGAfOprsq7DJOo
AWiZaQap88nX9OT95HBUcqGLcuWwhuRRupjJ8Wiz//1YD3MRvVEiqnSfJplR6K0Q
VTYemQX4Dx9pyP1rS+z7Znm0XYO+tm4QaqzOFG+aFMlZQwKqZutRe5qqs1gjeh+t
P4QF4NxB7ja5YOeSqTYyf0Tt5b799yZYgkhDeR545ZYm1yCmpLUiWFk7KYvrisjP
iCpR88SYsJ8eW9o3R/p10n4RfE35ER8S9JmufY9WJCACH/eCiYDcz2+HZvlECnYR
/OcqP03nY3IxRw5WrmJQ8YMPKnG2HvT3LeZXkTDTayoJ2z9/MfkOWJtVRoF+mv84
em2iFOIiJtWkVTrmM/PEN9N36Ajk+wyeiCPQCOWyZLQfbaKcOrlrHOn9zrvSfzII
TVJQ9jFWUZHihH/GKA0uKn3iUpO2L9dg+TDUeHadILJHT8or+i/GELGwQ64sWkD0
FGL6SCgIAQC976/cG/ew3g4KJ3+v14CHEsLjVC9VaJjzDX5Ve4M1ipGfxnsyimyc
EtNgGLOyjKCLYAPnbMyFPSRStIKOXPx8bncq0NKZ9VCdBXxvqCwrxl2QJdnhW+tj
afzgOyZ4D17ukCcLA51dysSevFiIy69HQ4Ap1pCpTH0rew/siSSt7D9OIn4MGy+0
CopryW/bMTaceZIgRh8INu0RvmGkM54N7lo3lyhVrRIsyDIzbHikNGjNTAgX0czB
oKRD5pT57OcoNkb/iO6szCYPuE4XxDt67iXtdCO4FLqS0MAz2tfV7V12ddsxooz/
VMXkAxcbrTDHbo8ce4/UkKhOpVrYeGRZNaea58LIypXNuPxPPH6NeIN3Lo1FtQa6
mMIr5iswkLxOkJTA7Lqg0wlctAccJVHeGFol3PZ2SdWE9w11DI7JDwtdyEpv0ICG
st05TIPE09nH5lloIYG7INWgcsKfalfN7qA7n6uJXSvRsYscfn0N27EhSG1ot6B+
ZBrVSFsp1BqTl2SbrbZlRrZK2AGZf6BDKWyv2RuD8/v8+xi7S6cxXMS3Tc/dAVfN
ed9S/DLAgK8kpsrV2k8Oc6TGVWqets4ktx2j6XFsPfqQo4CtaSPsVNLb0TxSayvR
rPYMLQqN2fzBFnxUEu2LwlaxgicdOZVIuUbh5/LlQJCsO/Vx+xe6EqK+0RAqRUtN
JUj6E1Mr2tUzWt2bBOfP6kgQxnZsOsBfHGwPbZvlcQv2LCD85PjqSiWFLQjKPexD
wNSQoKgLUjFISiqAJWHasIdWYZljs2zicQyu7izUpITMre0zC4HwbKsdd322uPGW
oKswgxcaeBKgT+q4ncnXPvRsKSAsgcBl20RzX6axu+HSw/XcrOGOidM/2vCKUsHg
sD+eUYZe35fP/QOhC9TWJrnuPFFYZP7YT3LOPjNu7ZvJqUsGSeMlwkLHLvR2wdqF
etTtFM6esgPF9GGrV+hmS0t7X4dLqSEDFOyAZCuKP/N7hMiGFznr5/Pvppa9S2gd
ipY72SIcwBaOSgS/9MnyJBATyz052NTqY80Zktvo0s5ZI6usAMN77w8jc6HkrXyA
Aq5UAIKBNP5jNmeYXb00WWUoykPf30IUZRW2W3CzPzL3+qZCDwz0UBhYZGG6Lxr8
g/nCrE1puZSm+3H50R/aTSQtflDTuab5fMf7p6q0QMWqEW4IgaSwG3KC3Qc+0zhn
trOIRtN7i8qtSq+zNzF1K8K+Nkxytu8rVfk5n5w3kWY+v5CD8dyt0n38AW4Hbta/
iqMxergM4h1d+8jYfWaAaXeg06RiENTLrqw4vJ9zR3Oi5RiOY+WFqve3MhYlYqQ4
oM7fwwUqM8r8Qsk8ByQLyYGeNIi8buPyGOySm5EIPPuJMsqO9SzxJZEbeiBGjXoh
m6FARMgFhwY92FHdtBVxitNdy3R3xx66lp87ubn3gL02pIQztBwrqotgW6saf/8c
XFtMXfjg1YTjzbRu8YxlPpS+FSJVj+VM7yNy8aqMv8Q0dyoiuU/aVxYOVCv6yZQ4
H4DHmxQ6R9p/zxGzUel4VfItX6E6zb4G5mamzT7zMte0bQPOMyWfUHq2LTJIfZPF
nYswL0+OKCRLptns2xud3+IdvJ0kgX0twfo7oR7xuXb0INbekhq6zXBzGRufSRzX
s1dVR8yhofLTGfTRwUFrKAFAhGP4aHHlrvSk9EFibt7kMucEids6IZvjytGY0uTu
ugonWBAir49CyopI4sS688YHyoDI56DbHYbWtW3934GP13wVRVeeX9RqsKxPIgBs
37cDSetg8ziAwzLx6aAznba0rTsTXuL4Qi++JpRx/XfElcKHJn8JY+PtcvjSxyPn
9Fk2UwZnTnqb9/0GnvIAKRltSUOsPw0IEIO9rMor+dWron5i6uhE4WR6ET6JruZa
9gk0JxK1u2UodErx+MnWqRM8QOfjgnkM/+zQcOGbiyoU+mCiZxPgwq4TgwxqKANc
AZQcWdfTfBnXZsMmroZyreWLPp2yLYvKW/8PHXyUgMST+zAnvFtF0KPFm6fVBD81
Ao/QvMSloiRXKLfaOdf5qHjFU/PbTZGKqwLHuEDOGM8bPP6jBztwXEl1O2nJSLVc
wcsTX8mO3bo55T/AVLNRXcY3nu6ZNwIDuCnofd/EK9RcOVDJM9LII8O6Xj/kH6Vu
k07Ja3VNSx/XV8A4Yx38kvZisV+1ijPj/JINz8oRhCUNKP4l97KwsNisT6anfhgz
tOatmYTBX5twevfJB85QSocXRtKpGVlXEz+L+iiMDm7UZx85ppsi5UgTmIe4/sw8
UvICgAVsVFUbzigoJDTmHC/3K74YlB//QxxT6vL/UKoygQptIntfaRL1wVwpx7TL
ckzjeLyXUI81UE+CaLwalZ0+6SauxExeDzRl28ZPf5OGQRx4rqIPCtZAUdF5ZlJM
3S6eL6cl8zOvIKIVBuM7CDWKhpJV9aEOJhPTzLVxDN/HN2T7GRWKYkxJEskMrkoa
8GiAH64n6MDL77/+7mByygm17jJ+6hWs/noEg5UUsRai+Iet9/oE8e5JwvtIb6NS
stQDumP5DfGQQ3tfdfBzdeLimJXJ4ubEPVnEpWG7rA3i8dX6jea6lrb46NnPJRV5
0zqnzYNxW3fmhze+oR+7/znDHC5zNPXWgOUCvHRvqcGKC7P4EzsO4+V22TuXKB2i
GUdgI9zVc8xqppOT+qoHD3c1IiLf4+C82pD/Jxosnr5qeUwXF/+yuJcYKC0gxd6W
PjG6aRMs0WoRzzO2FA/qSRwiwEMN/rgiLASKMkt9LyZ3MLL2DU2mHgCEfUY+gaAs
QJynvhex5fjEJ56J/nvxzE+dQuG/e1ijOgKfvKdyXtJpYcDTUgIwAfvTOAlM5NXV
zRbB4xFgwapYOzCVYEKe3FRZ358FcIz2Xhy6qzgkAcY1nHi6lnFjGUJhbQXhpc4+
qyO54FHTf4b2yAwyO3hJ7Git+Gb0grEvvCZgRQv70htXn5uMra3DsysKfgtWSIWj
CV6XReRhTw1d8FnBTJHqedsTXFmml/olF4hTNSg8j7+gfvhyx54DhaweZZdv5FYs
DtQQy8BmXyrhUIcaL5F24n2x4G7m09XB8Ny5o/DckHDFtMgsFjr5YEoZeAZ4f7QR
AQ9HcDMAN0U6qtXlmQpO7LqUXfMYmPlz0isYJPsu+cMR/vi+165b7QmDZyNLlRoh
VdLSn9evZ5sn6/gEZT/EAIF5oLnBlvyg7B4BdpIOLSo8BYfGeXyukTBtxSyoFS/e
neRlDAfKlNTAShe5UxJFC5LJJtwSRNXTyrnejLFm7Qtnx+NbOuA7u1Ju31HnNcKD
ZIJrRVEqrUj43gs1DrBSOUgayl8UNsFuWuzxbbcBtjgAHcynL2Suo7o2gmuM9L9w
/mOfNgBqRiSqB9mws9nMtXF1KLDfDzH20IPnyEJv6e9+k6wKrPLEJdmunhx1wve1
ur9nlDh5IfE4eQhBEvaDaZvAglCypR4PbfWHnuF0XAtJuBiU8fQK6AvpE6r+SBNv
KenSRHDacjUYZcv8faw7NS1YHf0/eQuxsf3GW8j7E2I8GsZhx74Iok/tJK9JDSjG
zYI/c7XWXO70eY68C4YWJJXmXp08WlS5hWR8UgKPQuwUo30I7QT73O95buMB4ZOQ
vGpgUy00z92Ci//nmfRMXHABnK1G9dfHkg+CGO3m/FO1Nse5hWBOr217Ya/j3tPN
wXpOYH69CGiQa5s/doUu0khtSmSCQfwEF508t2AsrsuHLqsoUC23WbqCpN1l0BMH
1Lg2yZoSdasyjl8vOt/V/JsN64CxEUpLMF4ydyxIwtkAie+mMvcYfjqQkq+5J0o9
RMGfkZfIqsjZ3nwUprWmvTH75K+73TeSq/e4RB0sUw2bNB2BGO+NciDmj8lPwlMS
XGXuTitDlWZKLVdrQJHaim939ySyXYBx/FtV+lVc+Axf9u5c2KAHMxwWeRjLrJcj
Ekc2s7e/zus9QhruFIT1kQoTXg92mCPkw1qC5SqYi3zrfpOSWe8wGHPVwgyuOvN1
sQyNggZtLUgzhlaGjqq7TI+M49qUQJyodcMYNJ2rlonbDjlh1qdIVg0KMjx6bEIX
LNmZNUJK0pAUZwTjPWiOai28y766sqi00kL1aWBzqSt151u2AnBD53xPMe2sWvep
Lqq5bVWMujfnZtHLh/T6IbX8wUrXHyNmKuKtMmGNgry3EPtTNU1NgZawiCZiYVWO
T4PS/1aA/Y2047yBuDq5/cnhq+DrOgGusSxYvZcRo5uoFwncQhWcRGP6DautBwqB
7kgaJIlepopAUQHA0oNCktqOc/bqDxXiODvKQfRK6RMbfXocOXh5miKbH2elWPkF
cxizlg3uiYCCrY7Qe9lbvOkVjO4+BI5Wjy3IbNJpCqFkgxiScvZnjZlC5qqEJH/V
gcBqBhiOF2NECvxqKLTh/IU3OjOG6d7hsEcSH+8JQm2LmgmMSUFLI3uK7RZX7TPZ
gVJMbWJz7kxaNC8h63jVAg6PokgNo9aXCZMSkwSK0wTlMtZeN0XjZXh2fD2WyCzg
t/rEsbFRFkLvugXD4Cfw+y5hP7jicseIUFTtMirejSjBQA7x+5oGGDRBsq8zNtXh
o32DjrryLzzfIe2pGDAOHgUqIAxUWV0gQwur1uSucl5UahQPxz89ZHXnbZaIALdZ
cOR2hK/d/MZCrE5UP722JFGXCfungEwfJ+u7p+w4t4HgEUQCQi1Hv6j4TUK1HocP
e8xq4RFj8GKhxlk5NWkV0CX4GqGWJKzZ9Cj4YwrVl7YYv6FgFvxddvECsTbWK1aw
SUewrLIS/faEihQexsTIQUT6LIOgRH4w7lqy8Ui2SqdquH8qldq6YwOrykDAhvGw
8U3ShoIJVsKE/aASU9fgvrFl4m519RKQS8QmWIbBov9/gNRKV58Iock9mDRJh008
qPwf4AYdaMvsFR5fFuVqmjYGnoiFyoXB2sEXwCHTyE02bNM8lBKnZZPYV9M4ivP7
roL884ddJK5QJX5dYlMGeAZAF+MU3Ojg9zBDclw2XAUPYA0wLByd4beGiO0DQmoV
QCNf5svfJfdr0dhi7VN28bpZelPa9I+NND5rp8pVaY8LC+PM9+1jGoSpCvQ8xtrW
vVCRqjEuwzKXCflj6vnidMqdNbcT7xaM0HajvKUaTd9NJJOjQryUhPYsOoZl1b2D
XeTVPZmpBOrHBhMtWxRoaqjgW1xufq1OvstoJMkrybAYqVR65EO0fNEATAXrkizK
Nu70E1555F90fKd5/5+omzuF3KK/bwdYwSmfa2QG7M2oNh6cLz/nbXsLsN/CV5cv
qiCAuoH+BWizqgSNdHWHDzxcU8rH+JLEWROW3LGUc9za3vaiBng6vEX/DlGkAQvZ
18SU1rpG8nouFGzxBB2R686ckf7z+64G4LpDA4ESeFr8RiA473QCuOCIXYcXOAlQ
qJcBrrBLDWTzNoyo0uck4JTnSQSnFedFIzXMsWGKbIbhw9M8TCeMedbh8sB3ABrX
fqmAkddRfiFW/TXgkE2sZ1MdDB9AQzlMtsKSmS5nX87ehEnbyUIkP4ptZTo5ZXaS
y4TiUMH7MsEtFfI7zeOus8QKY7MF9yPGJ+6ighh0Q/S7f3BMgTiaRbdRvmRK8hK3
Q1B1mMKT7eHev+TNZJcpBK24Sq2q5opJUhI9WmQTUpQoP/9anXQvL3eyy8e+H+g5
31ocQYoyjpYv+9wk5UAaTUYBAf1l6jhCOvwwxRvu3ITtbhAO8mTNLd2RSCIMjJp1
iX8aoqXJCYuIIvInLswYIiPWvC9aUklAFQSjPkodyBmy+F+JvhPlgvnoPTD/HrDI
ZL4MbX7XCYRZB7DS4hgI4oLmXdA72WKvaY27tdDe+y8PvEcTXYrHOdfI2/7lAdqD
bWr3YzENxOddXcqYfsohHLa8bt+fKg1NBMjGaPoG70KBOwK2IgyW91Ro9tsPKfxC
xkSRFd11K2hKmffStimtM28l4Hqw9clL9r7dowvFwnSypPID/wD5niagxmPB2hFv
UwXtmviNEuor8kd34NO35IC7AabuIlMzSF2t79H4Jo3lhgr1cW7vgEcXbuaN9dhZ
b/VyCV2a/UzR28KaHNs5EjZlnbUNzesYpib2qhJNRjviTY/jD+zpH4tjfSxE4LMn
ARHrJMxWpwponobS/xUX2DxbHxqdf/1Akg2E0qZ9BysceobiINO6LHaZwiiZiVjX
ahUJE9NjWX/LtjjoTcRmVoNegIhpPHrR1NRmnEz3rzwpBq+zZQg2qKpGsajN4qDM
qqW/bwNzQFKE5AhlW65xsd4fvrWH3dQ9VgbS9+DPda8AwbErv6rUMck9mZQLxNwm
+RQCs9xrWEaCywA+bYpmCLwbyhUDUP8DhH3fvRMQVTb5PkZZyst/VWyPPF9G+qip
Me87MAjZQCyrbuLBia+9ln4JYq1ZRdg0OWFrBqNE6MlM82rYjq/FATSYA/FVg2D7
d7PYI0tWdRDQ6OX1TFp3rqgiqZ5ZD+dh+rlcSF9gbCTXEHh9ZrY9rshLL8Hp53cN
esMdhKLvA+O36XeC8id8bCKE4QgdOuJJDqJkg3C7FRpeayVFIOVj7o90p++tkQuS
ISQeXpJGwGVIBu8qHd3l1Gr1xYj8E76JLY2Ijn0x9SLLxM4CEY/rs1JMO1T099Nd
dlYCHWUCuFNMD4OzmI+Ze1djbnPAUoNY7/qkaJgsmzX1aJSmkLCeq1srQEN1hYJt
Ma4Tkl95iowkPwJRKVHgMhh5WvReJA+jU+rB8rThA4XphHKDaUEgY6X1YDASkQLY
hKeDUMKs3kpUm0yJoH07tTH0UsAZnTCdluqQMgvcJ4exOWInFPgG+fk1MMjpmrHP
Ws7+tTy11gL5lRBu6ps3sF4zNxkm7TX16DOO1E/HfKjKeyjjwjgpcgzEeHnNdy1s
DmK1K5U3kpb1pl/FuVOl4XQ32P8eLpIZqSdpv+9Zuhv3iuC80eBEuUTBKfAXA6IP
nHdx4FCe11HXuYo6Bmbz1jhGkmZylCtPYyMqkCs+MKEuDAmK/nK9Yj/1oaZvOYng
QYElmrlhC8h5T0GZTmpP6sdNivD78HNvJx6wBNxtPAWT52MlWsje1SkhYDR9sFy+
Vgc3pjf14bkMhYcfyTfuEm2DfMoys0mNbbw4YpLzKFo3ystvN3B+5uip6sUhrezU
NzLUEp+LWUVF4e1NOJh13qFbTdUS8GZCEADABvAFjm3sQISEJd0V+bOMFWeiIcPm
v4jbeL220iGbbd92aYYWga+pnWEIfhsOb2H4w9MYUk5v0/woguS/u/7OfB9PWoqJ
3ca2jmYvDgo906j959E1g0PxMQiGygg5O9r84ikj6+7c9KDTmYPESnYccXZz4rbr
wBTVjapIcGsbc9Ud+RX+a8O/Cqd4TqNmxbALsdTkQE3E1EDaru6npIoEg3vZ4rd7
vFhtRJvxpAiwRd3I0ASw4Vlw7xRvU3GOfrr/+jDnDZeTY20joXY7lg0R67D+qKZ4
amj6MXippwaKL1Qi2wbLJqgBxCTK4e591kFazm5yiE46nHaINu55XPXV2NORVdRw
dfHa4lHS1ttPoL9eE01ieAG7Yy6gPpD2bh+PoDPhx03QRf5tYAY3XHufzHWQA3Wl
w0i6dp9SYiIHYJfcNQcxo66Njbc9/u072kZO1yL6jXHjmnPCtKfNa9gpkZpSkCaH
r1sj5/6XG2rMe3RaY8VfIuQnEgnca3vzXKZNkotPfViepK1kLGiPjI1ZKU9Jpqt9
Jm6LJnNM2qolglLGu7gb7ZVSrnSebZDbLKTktZL4mWQz3jqqJm7Dn7SI7yCI9hsp
+o4xa901CY+C+mW8XbFGvy9LfKzdlZYq6fbyvzIGsUE7b7zQRNut7wwnqhqDD3Wm
H2G7moISxDMRlAf6U2cclQRaxIDj7utkUDWpk6IHtBtK6cYZPnS503DPsF1gxec4
Zmaxbj2DZe955WTRynnZYYZeuGmbEraGGdrQ58AILUmlrQtbjhU72WiNZpe5TtQr
g76ycYYq4vLmZjZ5fITm2e5Xak1ls7VsXgQNEVXFWJcSkABrNQyTq4n/pDxj+rrj
n9krNFKrIpFOh1axCCdpah6+T8ov7e/nBZrUHoI/fqOjyYSbBA7+Tfvm3xU1qMzI
NYHSgaxPPGEt8NkIwVTFwt9hV0kIwlXJ6x7qYXwwOvNz3BpdiJez28ToltaHqHMW
KD/PoVdVRvNLe839vAgp0htQMfXgPYK5n9V80+U2pR5sCDrIQZowbVIB6zoOl3jw
c/HGxD9LfLiWcntNv7Sx/EnD1BCyQaTHlatrFAXdXwB8OFSmEszTQJqisU17D2HK
Q2GIW7FxsedrM8UYJtwXJTG3hOs3KLy7VJ3cV5o+3oH2Jm4u+v+2LQMLgr/dfQZ7
Az8un1YFk1ArJJZ8aVe+M6Q9LaS40hR+8JbkTiHrsCMTJWKQJ4ojk7H4eQWe4ktW
ws8EE6G2a5GW1PQXZa9HP+oZf1MzB3Mn21afhjEGNHu3erPF4acSETpMaoCMA1Ce
tlgKciRiMJRYWpE5sCkhOoxBtRpT2KXFetjpKJ1RmTdCOruVUGYBDiGa57Vqb6HY
irQiaZDlLoknsnJAy+bfCEAJogFmHyBgdgqY7a0mZLJ+W1E6qHG8r8f6/8/4uIZq
xKhBFQvLGtZmXthsTUYN+asr/mLcvetxeNKC9lJngUN/DwHq2Ud/4slfF9wD5Pfz
1Ga0OXeAY7Y+bIoxKK/Id7HV1+NbaksTItj+5TO4JQnPVr9Lygokv9ZKbOYZtgrr
WNld5njP6uE0DrDxhfDkX27LK5g35pyscwC5KUhxMhJLPLxipgtw9k7ICVTOkoUH
B9mSD+HvqxDw9aQGD82ofzZbr94o8puSFa6RsFalaBbHhpvFNAsIi9uizBDP1GRT
UTRh/vXMbCsuGknUCP6qBUfIiTX37QQ3qg8umwZ6mZMPi6em0E2l97nON5zttFLz
ei0qkrTKzF3hK00iJM2sxFIzAzDZ89YeN+hiEPeqt9l67kAbGgUGkCpjhl0B0FUu
a9uO2RwrxifP2huOwjBd85xrO9LXHknJmaNbYasaZKWgPZV/9MyBkuDp6ITn+B99
RXpqyUdtdybgLb85lT2lFCQWFpYrK7vdgdCTZxS42X06CW9se2cmeRcV3IilFBRg
LPlmifI1ZOn7e/fWHl5jMnaDbEna3zJBxMzs8OW9QZVX9FVJgQWa3apg2cYsen7f
PIOpHLi8kHaVYXCnaED6ThuoXjBBa+Awpfyf5hrKkDtN6518NeOfA0udyRo2ks+R
aVSSvI+GhHF/zUunBWHOUaeFx2I/Z9rNGN0ggdl/xgYGvy7Yh1M96eW6+X7H1K/P
TpZ92opsQI0pdnomEEWLy4+8J42C0A/tPa3tGbI92HuT6fMVUL6hDCEGQmBHSh9F
UW3D5qnwJH5CdgLNxEQakG5Wq6ZS1UabuamKOiUsBfSeXtxirlg2Ls5KmAXecWAT
Yeo8ST7y1wC+VEHWMBPq9KAyqSu56T7T3au1tGgCumMJ1TIYjxn6ZyxDPz0QZlQD
nfMcszQhg+z5DepcWmnh1V4sZPLkv04va3JMiE8YXuMdXB+GJJJwibL8DsUqs/My
T7VazzjJF8TU1BeMY+2RmsQX2yd9AoN0XhREh78ih4ZzWfvXFQULrTfr7HNp1BJn
ukmMwLLLt0uqymfr0xtnRUfX+l3WJSvnraknlMDaU6ndxtYj3fxPU6t8prxmiNGf
lHvnTWQJHuxvsKTp+pCPxFT0Qo+rIHw9iQQuJCmYolJiyiVnJqOxMw64HsxlYgec
rzGaDYAmfP0/a1okhD2K7f+neUJiu6lp/tRnuHHLiHDvk1FcjcvNwU7q4hHucM4q
GgRF4cn7BaA1UIt8Dr32OYwnDH8gAU2aBVQE6uWJPnjJQIRjHYH7nZx3vjGqlN9i
YpFO30IZr9hjh3SlMYIFteTfK0wfzWINDnGn84MDULLIWJJ1ITbIE4Ot9BnKgHbg
KXkrM/RuTfKmtOrrbuEHhRHv2urAr3pqc5pIZWolMZzGcyCBHY9+50Div92O441e
eZ7f4Og2WGUNJYTFKKUdDQmelg66DW5HcaR0/XMYaCPpW0ghmM1nkUa7E82YQsO3
Kf6ndh6C9wIq8m2h8D7Ibe3pDQD8TGz9WMYs8R60pS5YjnZ0GtspqIzMGS8M/woD
rSopDFr/kx88Pb4xuEj6834fGnPXFT4USDHIIKC8ZJnu1QFy89yHPVnoZdVEIcVs
QAhCkybtHT6cgxGYTcFwB8LdkVyRf9s5yGysGt/eSqsppXWaxSywz5rn0kECyd6c
aBb7i07lpIhUREbpA+Nd3mXhEhL6QHVHEG/D8dcViLA9mH422Fa1/2FL30mh+Cu9
ImLBAgt20XJ7+ol1pVEnRXZ71NisUDkF9wIZWrZnRns5pkdmEJCaIcdX7q7bcpGx
IwiFsmYz95Yn8yxiO+TulIeuP0ML3ZmbrRpXNq58wCcRBaJVUYZdMAjOAkqBD2n2
G8ZLsROMxDZFpwsg3fzb+g2LBdNYn4WrVWd10+2Q7QSzatbW+MJh8qWKV3SHnpX4
u2clWSn0x2SxMZDirHFEpP7aaoo8v+SnTvWOaR9J4yAyFtlsBQ+StMM16XpXe9Sn
DMRTkeAEMSUpKeyJ8GWxx9UY75kUSrBvgj8iHtu+LjEoUjVMTyvfNldOjaf0HDjS
B25fjgU0kYenWgDfXXebO0H7lZW/sRAxztaI+4zmAzJYkFrtpITSvy2jFfXmyxbZ
XtWisAh8An6CZCAREIqeKSGD9/M5rUtbO9AETpnL6kH+w8rHTc308tZP7NSX+vrA
p/g4YTiKq+H8cS0qzM2HaYIeoRhbwMsHb76gnCovgvA9TcrN42qjjX1hHD3KcCC8
S0xwrRLIiu2cCBLN7N+tV/XCGYSck3NPVkKK2Cur0gCdNF5JJvMYdg9WNH4DJvzu
1HfmHbD9/nr1TNYd7v0r9CyUqw9dcN2aTE0jcShaZnGxM4/sOmd/XYSodZNOu4pw
WKnAYcZo0fPOC5VDdOJSMh5aaqv4X1O3fUBLpDeIIRVvWLSnTFvo9oGxAvb8ZW7A
nlAjSzWivHN9KivpeGhduKEwmXjUbKGkrboOE/SVbQypsNcUa0ebMN66GXObeXeQ
p/TSVAyeK18hb/Zg6IdI/OWcHoZdDAVzKIAI7PQQ4+rhnedtQk+i5qxjB1mDU/s+
3CfWcIVGXg0wVGBCVupi5ZcqxX9+OLx/paRswsz8mAX9GzNd1e5y5zjpH28XfbrT
21bnmNqWq6fyyBsLWDEYtvHh7LT8zhrkVJ2L9USkCxGyn6+9cCWoWwY2lo0Y0af1
ERKAL+4Ui3LSCqshd/raAf3x1W8Crh+jqt0NhR9+NPbNQvCxL6UIdAaBWBjrfsbK
8qoZbR/LklJHvyZA3XUvyt3X5uq0R1RmDFUyb/tqr1qYdrehyGe3JGJtN6fDXI7v
G/I41fdqPxTrYNO3jmrBW1PmWzs7Mkx4rWSL7rd9JNjVOpiW9dqRQxiDaZTQxYNp
BGcXuhIKQ6Frini7A9y7ha+ELjgWMJnkp07yx98n15jjM6Vpu04UuWylMWB9SmWZ
856Wc0WqbX4tUhss+TOJ3P1xwGfqC/YLYr8a7DMBQHvJk57lukAYkO/spWnroolY
K9uaLTHWpSMKPvxOwv4tnBmWiQE8nCuPU+9RpAsvJcnNB9bbItDsE2xJ3BTKEd7A
8O6XkCSmGOresIWkDvufckCloWo4EFG2ga9edEyAhznQzj8xuAoKLGXXV7ipod8a
/OBrf8ES+fuwWWVLW/uhguxSRaivjrcRy8Yh7cPMNT4VouWMBaLFLH4tw3l3cfLo
I0Yn0whn95s76ibznB5ge/mVz+YFMRXndjBI5rlVhCFkkhELv6XLQwPeNPwZdx0D
uWegSIbr0ZQlqRa2LcHKcEDxt5L/i7qq7JvpJ/Qb/zId/4d48h64tq/j0WRFalXc
euTn4QeJPW36DW/WafHORZQbSoSWDmYauzxxigr9s8KqEdtilpJpacEBQ+K44oPB
mquUsW16/RjqJ12MRnSU+ijthpeTm7lOyG10EbzDK8yYUw0//YBykzdOk2ddczEi
jiFlM7w6DcpmobVGM4P1ZpqJm9pYmEdEDbaubtD2vp6oi+Z+ovTgglV1jjgVFbeQ
J5UbvPmdKEH9TbjEPgErbnmIVPcXO79RFXidhOzPp2GOh+1oTEMVBZr4z9yic/5B
rNqNalXhV1K2NxD+h/AIZrL/bODl4WtraOAylDAtjhXtOFkbeOch4qGKrIuYuMNk
PMjoVDcJTwGexXSu3gdLEGIGYvaO8R7bFBCF485w+1goWj1GKjx2RYllRgjalZBV
lUQKdugl90EHJztf5v6NrVWSh7AjjhfDwRjaRy5igJpBiIk4pGJ+GfbJ6bs+qzri
u8cnTNEi16cMjDMBE66ObgTZlEU4+XxpmsWNzAsdbZWtLPiDCUE0m7BGn8Biylya
um9hN/3+mx88e8d1JOIBYJurkXXaFUGFpqddevMKmso4P7QGlhRWn41x1ZW6qcLp
41qHNUd+zfWLa233zXpwn2ibKVpsXla7p0tUxqeJmiBsdlk46kOXeCUnYpLilFMx
nwRFyIp3AQ75ASQG8K0pedmiDvCrUw8bzZTktKPIF5bwla8YvYvpjjJQieApcQNr
pbJDxq7gLgB002iNkxTLjwqPB/EoL+ZZGsU9ytMn4Q+IsGwADVEqs7fbRoScDSKL
qUySui17auVM9ecK2UB78R97vdqfTKYwyX1U/BlOZ0XAS/+9ie09g+YF3Mjt2uLU
v2m37a4naV2I14JleUsDGEEJR56Izme0lwg6huLqrEQJ25jJskfRyB2BhySjlbP5
xAaYWK7cxUtEbGbwtfH7uGehLvaC57PTM2GeZl159Jt9bNNmMwaI+6l5IlXnM+64
/6dXnn+WatYyJgVbsxj9EsREUYKO7CDu7G61XNl/i4UAoJqcyzszGWdrn7HeWP6L
Qen2BBuZ98MIBWmBgRK0KlVMb74zIHNyNFjiZR+wkiT8ehORzI7ACFPAkS4av7on
2+NgfcjjUkeSukK7EaDEoDQ3zQZ2dqEJI6xHoTSTsJy9xqWK6ZOmZ2wI1dFnMAtc
uQRDz+vhpCnOaNtHnaSOyOf3bJXp2O0nbo7FWlYbPvQsomuK4SK3+eRnwDDKnPGe
hsQkzxrKVD28Pe5gV+jvgNWy9Z64l6FixKwDYmq6VuzYkS4m7ly3K5nhwRzYUAhN
yuCKuY45HWSe6/ExrMk7Fc8Yyn3QxVXdPht0+AOtCt/6t7yOetS+tsJoym1/FWzD
YwZdSosHqlNVchV7f+gowdFqswo27zQ0pM3YbFygYwpLONTlFQTSzbJ0CpdSlgKN
J1vicUIg37je/TUX1AJTashThqJG9Q9cOetxrWoqM60tpVPyQdCzxz3N0l+tWLjB
qbtdq9SU/4Z33IU3HcDqzxqc1Zd5PhKxwNayy2ca2hHJdF+ehd08rXrY/w/r8XZy
akfJIcAj2C4uWENcJkjXJzwUrcR10WWowQDL3iuaYs+t9o0CnRlvHWXflFDuxSfI
oOeUdjWxORtYMUWupk0lhUjpeJHnaKKJsWa9tL+yYKc2cu/EU0UQf2gf6TxxDH8o
zslH82vBRpmGO25oGAuiERB/fDRabWhgI7NNB44RHLVWH5CcKYoCb1fzWkeg7+fr
sDfK1RcP9nB5p8B8eQHrMqfOvy1nm7byR/wpi7OB1ocStpqCJHYXgjIdMhwCTFjA
8JdlZJfJj3A/KegAEtifuwywg/1RE83QvG5iIRuh/HthS+69sRup6YTHN8+irThB
qNoKmWAmbPPyWBsrRWoIlUXDxqlR67E/SrUcKEVGWMjYDTcHK8sHuY52p8vWZXQf
duQB1L8JyxHVz3wxMfACn1pPTctxshPKr0dUkX1LGfmM039qKbBsyw+KOCrIAIhL
PWjo2c9QHRv4fJvNFwb3CzjFqTokzbu9cXtDOyDIpz6DpuEclyRFCfe7wvx/og3O
roy3qrnmFKjdNFowf1cpl1NwhMtrjypOx24P6aEHysY14ROc4326tGBAhbbJJ2Gk
XKuRfATXsju01IoLybMHQaPNuEbQQOeKY1xxShXgKDtaoecLFGOC5EnHoh7iAoxc
NXM75XaqA8UTSSGjS4UTFj7d0Au2GixmN3jJVEs7oYQrKF56WmJ+p1CF4GrfcCEF
YCMBc5qZnVkWA/m91ZrrSWjelr5FJ1by/BZOt1EwBPi8hvSvVwPXaFCGFopWvq8/
IGIlIrMEeFkFqJJ0aPvf0m+l2CVaqWiOxj9I/hZP49NYinBKSAOSsVpJk2ArLkDu
NBXSXLa5vds1NTwE26hI2tFcT3hYgdj/4CxgabLZiIPQZORf5rAeIl40yE96R8an
2GtHEoC14Pcd4l+/Y73tG3SFjmRPHX2Hd190sJNaLUWpGYKPko1UMNx5kepthpEE
m8Yjpd6v8g/pqfeUmkEKf3cAZe2chLXO2JxcGc869TZbagWmu61y991Ehp4n9xM4
OsmezRa5JrzG9mIZGAlI3RGkPGC6jUnA/OY9q0peY5A9vmrVT7uP2awnR3qp/OkA
o/fzOXODysezCfwANWm6nAOStlE9NFoJge3gF0rL3gjdorRQr88HvhAlx1CJSvOw
s7RRCHvxhc8mk3Bj6abmmCjZPvUOkIhtaBFCURWG8rSkG0aMkOwxArdj7m0EJlAs
agS4ZelyxB/MAD91F0jQj5ythef3+QVCY/lcez32QIRcsEolr0LV28yst9ttJO8F
R+x08G/EquqTCalEXCht+2BQlyBmrK6et6oSjW5LPiUUSUp/6+5lTF3IwB3X8SpL
XmSmuO1YnC5xxUiegnVEdOojDr4wcd1+tMMnpGlJqti6Ew9Jch4WxcSF2AogqW9K
nzAEwlFxHI5xvZRD4Fj2X5ZXR1EW8d7Zw8qBfo4Z1qROlAokzpjAZuIHoEeF3YOr
Ryj4PHM7RogNpHLZifsJa1UQgFKqfOAwJNSxgkrpE8V9/voZmso/CbzswZ8631yR
tWfeWtEzJUx9pHNReHfcemyUTtraNKWdOqqTigE6ILR+zaYf5Q4IxdEbn8sxVht2
rlSoMpLBCDIlDp/Mz8/5AYn/6sOoBTQOupZQf797VcqAwrRJKRh6AVPUg+wXVuAB
TMJSt9y//oRc0D4KnZXdPcekJ8114VpBvMbmKBhJBSZiWJed25IkEtaSRUfZDguF
4pq6FPdiOkfd6Rom5MfyjXijjTLHrTdvpqDIuHztXmwc/CyMcSwHVz28O4xCkxZt
Dy7XKCT8OTrDHP6pKVZZ41mRXac99h16ApXOb+5TMiLB9KTvNUzk/KvHCsf8DYHm
AJkkwgrFfpni4mhPkaelyD5Q8p7z8uFwRx+bHPUHDWL89s1XWryLQo85PYv9wDQu
a/yQd4sLVSIXT2eZP4WbxKyS0S8FKhmTe5Jvgy3QyHSzrQoLrLuiQuCEx3/JMiS9
Hgn7E5wZVjcVso39Tvy6wqV9ocafwiM3M7qUJaB9GQaqDxrMs/OWLA37mzQWgL6f
Yf5rXOfwNt4aTJwn3Mpl4J+1Jt3gG7nnHjJcYuYLYEdaquM2lOWFFnWfYwyrFMA2
VPpZPfJA0PFE87D/NNNAM36q8moZihyJwvU2xSslWOZXGWEF2DT3s6pDp/52o7cX
ul8qflVpwuPapQ2J7XsYtnUk6c8Hk7fkXq1deyDivmouVqpM4U2l92UzN3JmkRlp
diI6GKqxRg8hLlXlGEs8SqqolYv6GoRztnb/j/CarCysoHd7gKDJhwtfiniJ0DXY
aKv+EmKEnzVKy/DUA0NXrm9AQ/Tu2YcPHwXB7IXmpaXUaP8p5/ct0Cb8r0AnJ7aV
kDNmNdGEOkZpxVCI8o4M3worldpzzFzfTnh9b0A38jaiH86Xxg4ua2whmIofiIfv
mh+08N4uDMPbqPWw3JDg0zr6V1c41vuEN3sGUJ34psw4WTBVCAmzYv5y1HMQzo7D
sgXmD7qhfAkRpu7gibjXXHx9CXJ15bBO2keMj6xQx6UEv6myrqutiXKM/q2LhfZs
nnYM0Wpb1G1XbHJWq23ss2j8p3xTxKjKKrMZox0Nn3Rpa8D2cNjKRgT2u2G7NObN
o9Q6e542QvUIJiIbrub1g9p+g2f35n+00L27bTZu6wbvVKX3xLx86v2PAIiPzgIT
IjBXNP+xnQudSJHjr6znV7xVj15N2IU/roYfR4toxyrAIDqc7+rAfrQikzbgmsvs
OhB/srHKAQr4JNkr4/2Dn7HarWJwNu9SuAES+NNmB7UR1/p82KGQwsMg0avxuprU
7INakyn8oetILSfho2ZLQAKy62dgkSNDgYdyfCn96xQqZJbsZ/sPpUex8rMwBX7/
7n1aJesUgBtPzQTu4Y0XT1WCztV+f4CrJOOAPlizOyhshdlyUwZzPmbCyWbGsFYT
Fh9EXtO7BaJ/sCqVT72JDD7KeJ52Bj1pVcikQAGpJGZvZiA/o2jk3r9qJtZGUoeS
bxvxQha/TeEKvei6VQBaCKjTUOJqb88kmgQiKAT0C1kirT9wOwIkfFgE91+y75We
q1p5AQRqF+0AaEFsUSVY422nQmukaYVc2gCF0/wruLJba1qWrqMQscHainaRklH/
MnoqBHk33Q/2As51mvhg2S+6bwcQnWGQImWjeEY3EB/dmAtU/l2uFZewUvhHMwEr
OQwlv+Uqzoewmmcy5LdBzg7MKi+nL2W3bKGQSzwUa3Et9Y2V/2OT1G3Ca6iIh+4r
tcoXvLPXjNyLxFQF8tQIWhYIVRnTnZyRtcYAFbfuyYVjatFsTLvL49kxR+yuEcL7
0ptous8SNoqrHLlLFmx3WuOIuWugOzJYqTA5P/ElV156h7qKk7DqYYC6YETEVUIF
Vnx7NRqcnpUFbl4gix7fzodbLlMdqLqkT6utkPvibwdLIS/6lwtMRHkU1g3BAGh7
rO72OGko8kti2TMvVsdAcoemEpBTK/w4ovck6nL/zkcSx0ml1NEOie5PZHTZMLeC
7ur2Uex8+ToLVlD6ANfIwpxyttmFULEHk4URr4neR09Z/MejhB6bdTWE8aiad3NB
zmi84B8eJpxLKQMlpX57JKuHJ1vzze1LPHa2NdtIzFRRL6PYkYUEVdPze4mFH/q1
1zsDxdLam+DWiCgVM/vVEY9i8uivpurhcf6bR+j0M/mKg94Mdpja/o9McoQucjIN
95Y1vdxl2OgPzfOvX13bG54oHB8YYOFf+L+D+y3LZXg4011Ii2ZDPIVUaY1SjT4k
BJ+ueEQTkexCTCyTMnisLifkU7sbWaOzsVocZT+60DFH/zRDXseDO/bGIYTvz5Rr
3P24GanMTnNmBNy5Qz/zhbfiVbT3mF+ySnau1PE74l5t+xs98MzOS3S/KeP9yUW/
U6B/hdqS9kwoOWgH2b/Viltp3QLkVDRgby78VQS3xzr4pP2wDSI9pJzFZpjsiIuj
Jm5les57raQEx2ecQHv9K7dU8tTG2HKhToU4qdtP2HxPi4IBHOtzSLhBVFzE0kN2
rVZlphia9ZEAbrP7yDy38nG/oWFzda/1cdwwhh2TfAlp1ZIfUoa8fDP9ZKHk6+AW
bnEJ7amN/deS05s6p4pNMVfAOt6J6e4RXYlZybD1ih50LZ7yyLUdfJ3GVRdoosaA
jP7EoUfxbEYJajaxC6SK8RD5dvAhA2YDZ+gsMemGB7hf7nhEw913hGhwnQz295P+
5FBC8CWFwHQ8KFkwAeEqtW2Lku8GJVK8yRmA4s06Hdy0lpm1lvdL8Ls7nG+1GeBn
Y5qOh+IR9YU23pgoajjpRI7vfhDvGsnZ3RGuA3SET70kmcermV1h1oXh3vexxywb
tsNmv5CQFwYQmKKlkwgtMaANDhYFVlkTCvEPgWimzi/97maNLu3mIq66QpUzsY29
mOOLMbdkxq/CSgnrHoPjH/wJwxhrq/KQ32rNKQ98khAGUvEZONwy6iehdmrIdJs0
ynWUd4Sq8xwJaPLQMqZJaunrWK+4bzE7zeCHBJTSP1q1qvW/CE+l44nvlJU4feNL
OrlDzVFswcA50BL7Bef8A1fiAVnMXrGZgs+ywdlIe6iomw2x9qI75CW4LAwmO+aI
S70n/cZl3LCAGWmFLaMEsRCTQSc7bQXtaRnxWcx8Tpj7fr0mvf8bzIH9ecYRGknr
BPjydP2kJw7t8f8DgBlJT+VoVbNj01ovSD+4Zz5elvYpiLdLg55Xm6U56w67GKMG
GQEeuTKWgyKq2HL3OCR4BUvJOYWRcmVbgzUtXj1A4gmOT5V+QAh6YpSvZyE0S1i/
bjX4Lpn7bN273SG5NY19Ehgkepf8fGx9hFbVWeBaTp++xzr53gs4Cj9wGJWYhXnx
eK/7+i7s/60JB1Vc4VunZnTbkhGl+6fR6/ZWrKefdSb0sl2ZnUHCgwDoI/zGg7a6
khN3jovHclLq4CGIIvMPncRdf2jNCpcqnq7yL6pUxQign4gU2tb3I7bFDiI5sawX
004trJnAfVWslqSBQyh+vydOa3HQHdwPfMyI8yeJSNxcV3TJAptPqp/nPFIgGS7W
lcby9pj9nsCvI8ZYsb9fZm23S/sESx1N3cVBclefMoaD6I09+YnHosIRqa0ScxGY
Z8C8s5HYlTm8EcPRJ7neV3AYJwFwcupqs3fLrYE5Fp2Wcft5Giq3akgtAhIiLNkl
Cu5+aM0BDcBAE7o1lyKR1d0N1iCMjco1jQQ+zVvhZidWyQan1j/tGlDKrVQ2WY1V
YbjpX/WRNghGU4K0Xo/16gW2+N1JVptyhKpv2LGH2C4Vq845OLkhgNVkIhRWljjL
uH+1TazRJ9pT57Q8FpSBA4nkr+aDy/FsbyMmRw3Dt/XqAxrSnPdq8BMi2DIYQ6VU
gCFH+g3c5fBoAB+M3JOJow2lluV4VpgZ4G661ItXmiFxfvd9tUSSHvWuuPGOgxpK
cKkJSmSi8LYWoCUYqwOljDnZPe5rZHOuLDCbZAlP+sn9cCwrT8iEdkUW6fdh54wx
U1bJGURWbkb9rlLn6Wfw8z1QEI4QzUPjOynYXk2Y8L0upQEcOT6oDe5dTb/+jSWd
nakKl9WnqxRO8WbosetoRTknaPiUCkQnxuN6qC+5FmbcAu54uELZ9Rm6El3wkz5g
8IV8zCTfGFExV5u4ZwEYHg5s6AdUNIsZ2s24AYC/OhCt3tVA9Wl9hapW5n4kBrgh
uLw0azV8yUWZxw81xsZasNjaJj7jziTKOGsyc14Nl1HIl1eY+KauOroGx98lU6S7
PgXArovZbW4eYjqA0DAASMWEmUmKcYytHOsz/cnT4OFRj52sy67IEWDvp2fXbuJE
b/ytrcG/NZasI9MdqtyOVf1C4gC+hayDUAV/rVw/44AeZ+K5b8KxqQ5N13waQGA5
+Uofozd/1Rqtmx/7/P99Mu2Q5oENIfFVH8Bo6UlrNOqDuWYrghU4ujbBk8Ff6X1l
SfWr1bTDMn22WemTnm2PiTISWCjxm0ufKxkHXzF1DrKKyvorcd6VF72BjA9nMR+J
lEjNaHuEWc0qTGKJFJJTcQenvn594tfNNeq4HVhfWgOYSrtpmd5NCoHQ3Z9oeNyN
gop5Hf9tvREP+kMCXGo+KbIn1zhi55HFDbAF4nsVyqj3UPWj12EvWSxFr3AL0z+8
aqZgjcMnFrvLR2nHark9t23UQqPlIckaT6tGBPR+h9m8yzXA4u3WBjN0fj7Ed54s
8gVxnA8ZZsOZ8gsG3pyKwlV0C7dDlZn9Qc20d7uVzSbF+DIm/R//0C6WbFhcArhD
lYwF5nItqZqx32X0h0fxWPYBSbemFiofBBRT/HUfGfyJXEjbdCI2cP0+FcLSQ7hK
7MLz0K1Ki/jENyAvakKQUTrsrSDyCGpX9UUnuAQbI27a2MTBCmXZnBTI4hl+nQpC
93zuRPPqjZZZiZzXErtxdRtenjI0BycQ6GJvjLeVBJv5eQHBCKkDznfrms3Bqb1t
0clw3xpaQomJWwzCKHsxrWanx5UXoxpacZfEpo7Ib6LF+Foq4waukXDh2b5GnAtx
jBQds4KQPuw/ou+avqhh8x63wfddiscE8nkI2+pvtZAwuAYiH4CX8f/P1rU4kUKq
OsOYI2sbEMXfw5qLSpJf0z0uUVA4OqvVlvOy7V/6SvcIZDfzBff4o2m/3GQNOnGq
8OYzp/8NYTaUCaXjW4JUADP1y3iU5HdiK9TCbCRJHjmqvDbc52NwhoBgfOJYDKrm
S/CFXOB+DOn12joqmFLzD//7obTe813pAk8sjN1xt5/ObG3WoGY7FmNzOZKqE53z
jT00wKUg8hppm6CZm5qfmvJv7CctywJEjLv9L9LpAx1B367RF/z7EMM3/r/OdoMy
RL6dzEwJwZH0Ak9HYaGdE3q1f3MXsMtw0oNNCOVC8Oc+7sDeuPYITVmkUKHOLHfx
E8Bh9dJaxyrjMRUlDvv8Q9ztk0ACg6Nb6EyJS5qd9qQAYLZdz+O1sdd/KKXMU+KY
aUkB/CAda5HWhvrsW751Q935uyeCOjwb4rjonK5YXnrljDF/kS8LLUqqx8OyQ7sO
cWgykXifNIKzNvsyBZGG/+Y/ts1OxH2lUZDKD3IgB7fP9aLqxN2mwwZskcIMiKUU
Fv9DyBer7LZsM+8pr0PvT6A/xy8ymupTYBakLC3ZypXJ+9nU/EuAe7lDQPzc8Uiw
WnJvXxIJYBNHiqPkW7KREHPAYyioPAtVucOFVX4BC4z5bQh/PDlKikpCHygI5j+0
XZ9jDQ2gAaTAZ+x7D6QT1x7fi+80eSfeSTuG7Vo4AIdjLARFTW7VK0BVe4GzrfL3
v+43HAeIMbdEWzY45Tmb48tS/1V5WdJrcyfE4xBCLBWiDvYC+4wunFffFNbsed9r
ayG6H+xImLeyU9IOadsfjvkGmBqroFjWlqT5atYQnT/KWHvt38lomNJ8I9rytuZ9
QqHTZU/zROdfbdjjbNrJcOdGdP0zcd0TnR8ddgJsmFgqtds5ZqyEkkyKITtinedB
BHCxZCzGKP2bvlnxirksrvRbDqcJMvlVbtwma9XQmetizioVkWbfHrUy5IJPbb6F
iGXkGqiHrLB+kQVN08ysTBis13G+asLTpIiHlM+uyiSDrMMJkXl3xM7q7DJN3/x2
JcK7psC0drWLrjk/eoula9ju8Ym4xgLQ3mfMWr/0rarygVYrtm7A/18WTMeazp1a
/XauC7vLFZLVagZmgQHthl0qLa3fRQ+32mvkaFhmC2jfKWs3e7hYTrkZTL27dEwK
8oThX1Flwm3QmH/h6XHo+wPHY8KhemfzI+xoWIrLsmwx8KUR2J6BhjbT0VZlbyv/
fyk0DlQKdvISevHGA1SxPO3I76ULhZUJ6CyeXl8qR2caQiZhLkXEkOuu9DOl9c+g
b7gLBN0EyA59xjhxbgAd5hTv8qmA2cdSvuLU0FhU+hUsmtQEuTRtJQ8IslHUA6pA
L+U/5jXB4HxbwaW5pD8tFUoH94FxPW4JqV/6RUV7NI95HKWUZhUkBo9ZpzY690DK
SFPDScUUB5u86dRVrAw2a4oI7wu3WO++jwSd9vmzA0JCGmidhAVNo2un/cYto13r
THe5j+HQvw2qERvkJJWoMTfEfd45eSrEYSsr5kyHtqiFkf7YVegrlTAadwhlAQHU
cHE2ujzSF1Zyfggx4fjGtSxz1G26m+XBVkTkNHm4JoN22emtlKj3NYu8andVt186
G4MH7Fm6hu7X5E3u2Fc0XKsZR+zH2yI76/v6i7bJPdGOJ9JWrmNfYJbK/U87H4Uw
Lk5lfKWMciNttGh8rMDEJwY3t6/I88TbIkDiP+PQPTB3LchJEI4EehuSiSjOt71V
7uQK02Nf4ngbldb7D5PJARS/hw3UL7NTduWn75ZqMyFz8p0SWDiFawUt7+34ULRH
b96iLveuqeH6jxNcVezHpDVi/+Vk7h43xfkKF0dMv5n2sie58ZUCBtQk+USkL+ah
g5Vv/KQJ50/vQcyaLPPiDf5JhsyuBGbtLCUeQc8N09KLJP6CW0UI88Ul0m6T77xu
4jZ3LgzYqkoFDP6W0hMznrvT51LjIFPZY18117XaRzxLDQDSSltrzgQ6Tzk10yMI
W7NR4UFKCG1mxYSutvi5qM6B+Ghkusa10cLYa8KRz6AtY5Lt+EXT2KvhFdiuwJMP
6j4GIVGD2kWkUX0C3kZhSo/JtFKnzke+Q/qE7T9YYUBDN1VLdEguw6lRC3ExUYoC
MywGaUMRixHdIxY5diXVCu8JT1oyA0Y9TNCX6/frTLKQTugutAzdITIrRAgsmbKI
2riXtK+w7+RgwgoOiSn7FNxaMZGc+K6fUWB5MmH6pqIbCMDAqGX+5lRKw3NRd3Zt
WbmHsIssZz9OgAmdz0xk8vTwhO/dEzSV6PQOR/bZIM7dKSjdcn6E7nenpllPX7eM
zA2d52yC2Z+HRcii7q3xuVhMftr0iSebb537nCtCPYTpg/8Efr6/RcvCWK0CjFiB
/WobDUPbMyeqloNXqAfCufFV+HoVdaVf8YcEEpM1JR9mSx6ke4HjEobD9XTcAyfe
YWERYyyyT9XWWf5hsnu1/iOBKuxUJRdu+cr+VzqbVRvhjzBxJH7FvjJ51LkxCgvK
2d31cTt2sVccUOKh51iDayTzN8KjC2/Q9NBe3062msRoSZNYwWS5zCA4RwcQEolm
ZBTSjhFyyCNZq6OyJ6tlCYhVEfU/DKDo77uKoc127QEVfe5uExvUiIxHoAURwUzX
T57UA9iNFmLZvtxG57CPfhjZ31KWm4gKPsMkP0S7oXuWSp2k1dnu2djgMNfwiC7g
vAvfgrR/fyaKjulJkbMBMKIqUlJh1f8NvKUb2XXCTeHfVgmTciA4P+94NGpzGd/F
PNg0doMZgCjaebpH2lLHZcn5RjZuOJb7zlVaJ/eqHeVebK2IOVUHYpJA5TnyGAmn
fRwax3FO5ei2rgOEXZ5HvaxpZwaj75X60jWqIqelWrqwjob1CYfVYc8gh4e5F/1r
TfoH3ahA36F3/rQfPst2CAuutARrO5DnjIZW39HX4hOe6N0XltN2FQ4vincslLc3
VVBe6QUu9WDBPo44P2nvwWEvbyMEi1/TzNK9qw5ZKuIFgSKiydBFbh5D7EQ7lAHT
rxqrvXAqFTJBiHrYr9qevejePRTOFu8I7F0NzP1cvebjDCYQOasVVTAPm5QFOw9I
siEDRlovSylxIW8xQFzg7DF/zrE5rokXjsiUesgc9viM3aTmRHoRghvQjVz0Thpc
nbbB9Juh+UpiyqTuyjxysu+aG4j/eFzjeBYBDEASGW/UW/06WhR4h1deF9dVAv7q
9N32BXkP7dADf8qMDwLy6vWBOB8Fqz4AU7MKfJiRN9eZmLf6fjMtkt0LSFgRuDYL
nGfTBz8UV+BwrBO/W02RewFvh8Ah8ZR3mBDyJNd0YAzE/ZTlvUbVNvsJ+v1rxrHU
6kljeHFvo2SGTiff/vTv1eya1E4spDG+4aBAfYJKy81nQrfu68nzzvhx2Ygs9QcB
eIy1xWQ06rfDyA2/bxFQLhi8IfWFYQLoZI1LAJGKUNYKTe44Z7MPasQ7VGPdrn9n
8Epgobs9Ja5MWZbdIL7hfVyDGaf5PEbje5yQ5+Ts8xgsrhthVNlNg9Zd85Ymc7U6
yZN4VxVwNV/69hN/eIe/+XuBKcfNXd2PQT1CmgDAqNLAFrXek2u7yg7rjG4N00HC
Gxsxzpeb06SQQIixW6M1ns1pT8lhaNCKoPpCv28E8zz3F8S9zs0Qfi9Asyv/cf6U
YuvoHAVb7dTHSQTyaSViE3HHVTnd6zrhbZEqmqWXEn0VkT2QTApw9X8ay4iGe7Mb
kLIPkXzj18gftL/T39gQLsnejYtRtKnGXWJZ0ocWb+tuv6bnCdJ9aDlqbsOGCFqF
kK3gSr9p3x6d+tTZ0MopUPEC5rx4TMOOm1JA991Dy3U72+OHbyzHJluLR8GXHZyD
kmSNoA+O6sNrEeFd1W1bR85BqLi8yA1SXw3L1ZxxvTGUzqDjMDuSKDQ0wbT9hekG
0AWnzrD0jnlIzcfXlArQLsonF2L5+lsDT6qBP3iC16ZYWiJISfP5G0V2cF7qGAmk
YT77YmCMwGI55rbbUfp7vNg5hSeDe362lS4idgr9Dyu2XSq69Az7bLsFkKNFiZ6N
A+hKGHefkF3KdS3Po0KYWapHjlMC+pZPSw5Ul08eIVpxkkDCsGzuyCptw/b+xPH0
um3g8nYTxz//lC4cpfRL7HLQYN0Q9NA5C4AOLy834EzXtqXi9GtjPggsNvZw/R8i
vIpGOQ0c1NX7t1/+iH558fiNypRBC4+tbObiTA76TevNuLJVAuoMFnLcOfJC0bsm
BpPA+nYWQu9SZRqOMBkC6zFlWXTPJJzxEEkmUGJ2Cy7MgsnOP1G+5O7T3Pr1dOyb
KU0IH6vPOxvFc8fUUytX+F8kDOMkb7RPEAk5wPoID7zcS3wX9LXbeYCR8UgZwCVz
Yh2OCSPOubkpkjS4rp48gAwkcWyR1JJA4zqUvYSnlF39sHczCoPxTt22pIjQVTxP
wPmIEaLaPBCy0ah4A9zM2vYV6j32BI5eUUlOgUbgLYbl6hry6lHGXjWcQvpZ6iNo
Xt/0QmI6ygYcqs8OREMBLu9/U81wvsDVwo3oJZ/s1Y7h+ujdpsYOltw2qEzACMav
mBiweFmNU/9TO4zHpgUuIC13zAA0JdghbWwpFbRr8ct0abDRU2stycnrTw1qrmT3
R4LxGzZXRGba2P1Ux0xq2lgkpIIrYLQgo4RijzYQABD5cG4448M3yzJUv/rSJ8Lw
UNq22AlLGd7jkHePEWl/fM9Iw/D7QFq+6uTC7WHTbFovCB+SguE826fXbpknisjo
hUtTarUva0QIV1lC0NrL6VFIWEC6SUQNDdCqu3juVkYDivwiAGkQtqOf+XPbF+uz
OMkzZ8BsTWlci7fLx3w86iXTOvgTZLfJeSdsFIk4m+iupxthed62lCHG3KdS7Bn/
4bHcR+Y0vnE1RR4zmxvMc57JNWkRUVDPR053PAUha7NnVAOOm+bLEbbN0rI69gDv
ky5pd31inanDhNmtxdY2tylWUX5HqYlUdZbp2vo+szw88vz4wzkvQy5eyfKmXHwC
aZWpl0suZUhjU/myvVV5nM2NGP5CSmrMhtuggoENL532UT503WxqUYky8NThRGTv
yJ2E/xWndXFwg23QPVsMY0WrQp6x5Y2ibfR3xf5lrBiDZjw9pk4/g29CVMG9ELXx
EvR7hUZCvoYnam4tEGUp8f8GtpfxE/CzxFU33lnSE4zTKQvGoceX0cxW0wjKeEhG
cPLnSlP9/m2cP+qn18t34Bq3gYN7D9cYOBkUpZIGDukEJA3y3QO4Tffg442wjxG9
2jU/0WMTV0V6715EM+Gt9QzntPj8gnHeh/gt85dSiyxZbfXjESbOlwZzYg/ttaku
GDhGIfloeXWwiYTywpJYtP/2qSvsAvlSbFvj0ZAFFYRuh4SB4x2na9P2CLC57xxE
OnYvpk9B6xeKXjMVkHSPXrVYobm29tpMGEKGNXQSqX7Q9h1c11g6VsySl2aRUCjf
jf7D3kNtfU7yzI1MvXse1GEv4kZXsfW0yyBKgQipAMxRNwVI3V5gbckaskkmQd5t
gTCV3kkC1Cz/lPcqTPyEMqS10jCzEya1y687cXxHswYrqspxL4zzCscrOGyb+bGo
ZBhnlN1tQ/kamaV8tdP/wel5Nlf+yebf2/wcXlfV9BufPDt5zR+ABq5RGexl1nUN
bVhvFmYB8G5nH3yPi+L21FHK8pknXaPc/WdgOTboIt3OzfghBAlq3D4yuapjh5To
ecnDIxcsZ+yTyZEo3ZCUr2RtgGSHHkZzn0RmDqjw19cXEuLzMelg/uKVUNrz0dyi
rpYG6GmtW8Sl/XsRkJcjeQH+buJdVkU71dDDpwYd5JhO+TXPJUX5oJsPO59S7cF4
sw+AAXom/Vc1EBR9UAoh+gBdjAv+PfvpR71M9Zk3ektijoSXdWon8e8eGl90Y/qI
DBY1/NXVIyQE3nAVBKFTSJE1sYEkFSwQTBbPDgeWoYf5YyR1pFcCgSHhuSZ0Qvh2
82D/QjFJcm18RwpP/K6qgON9Trnh/b6rDXJbjtTADqqc2Z/9OzzDjvj4sI9+qOv6
Tq6i2Y+Nw5LfTEZRnqORlX1iPCyfXmaE6c67DsrHS4iXWKyJGu3vuOz5mV7aH72x
aZNpjDgwqP8GZUuNNd7VRXUSBd+wf19k+0cLiIKkSskOHFcikq4GDkseXIdVXytc
n4A7IfksDGi+kh4P+ADTn7lRxfGab5iiGhQh9brBnVj+yndp+KXmxznrBu4vuBgM
TIobvN1jxtBe9WuJ401WJFGW4VUUGUYQoHURVOWZax0ScTtPWvciRoKvN99iBhRu
H9ExP2RVhv8+O105890lILpGX/23BcTBlaO9IofMFCjN3ZazqgXNBsEwLOQS6whl
XLFCi+z8+o6Cozb/UsOGtJIiub4rjWYmOcG1mdWv+rlmnvF121V1BjnJo+7xdF+u
I6lhE3xI07i3P3jW2+28Wg2NTm7sY0aZQAwUxGDN12YeIDuwzxqAzidVzakp+LU3
qLSz0v2sXj3zsxNxAtWe7WUYnRaUllTTXr/028rg1yWCkWttDF3R7CIsha5uhWJY
3M+tOcZ32GtxfLJqmHL0iLN/pNAzc9qsRaGr3wUc6hBYEJo9dtPPsbSiAR89pZdR
K3TypKKxJ1gVfuTbB+ITDdErGXcnCFNucAp/O2d08ji9mvPLHlEEhkf65w8taWG/
/iDJgq8JSGz1Y+b1kzgbrDq9KdNtFoMg/rO29sz0XQVjV28Veti+nwxJ+Jr7cxUM
0VPB3VR7MdHzK3AGS/+PG1F/QmPbCguNcb5pP9yIWD2r5qumalnt1cDFrqWPd64H
Se/Kg12Nkm2KFqmnCchHc++Pzo6o48Jh17BmCMexUycevb22bd4m6TLttc/ViANc
k9eKYZwiVATAmoa8uYL+ULFmppCyljjq94t9giQPhoh1QwMZ4lWpGqcN/eM0Ms1s
oeAR4TvrjS357qEwX6EKKKZnUPDWJeMGSsUS09KDpNjRdAKf8VowsDXLip4Q2IVN
4Iyvw4sf0a8pXSU9RDLdxe8gmglWgkkUxlRAiV6rXx7AXNaBpnYjQxEpbPWxtbxM
ts8FP86LE35HRloo1/ckuCtNUDfsYPdyTuVedO5vvRnfGDYqipfB2SCZNStrQIhc
yOLErddIpvtMLJYOQmArbQhr+uygS6ZUWcqB5Kb+c+BEitH8NWWiADx4FBaLdQsi
dHAoQHX5ha5zylT1Use//K9EmhwA05MKN2e0sUuAxQ/hlq9BFxiF4819Rvq9uBxs
2uZEFjd+YB+C+U6SVX3iFKfrGoimg+3qjW/POfunMeZ4vM87ydJo0JB8G9az7EJQ
JQVXBhaRJElDdcfmlXM8qM1hVJlNXGWKxRJI/KxbXJkHT/XI+OLjez6QY+WYEzXZ
Evf/XY5lJhFzROqyXnEG0YoIg5/wB8SKSBSyPUxdRA4J2a8zbM/NtMjENYRH84v+
W22GNAeeUssdnM0o+4OUsfXfvGhhsQkmmKGnfQvOSqX+pK26bl7YklfG/9yLP7n2
HtIhdzKSd6tytzExIPAMV7g9Fk+ZrwFRvsxuMuR2hS2vpUK4iIJLp/ThJMqHSdpG
EElpUMeviR6WD3JXGrciV0xAF+sQ3DeIzUN/tetMSYpilsopdoZb1G5ckbRA/l+m
L9ZdhzSjVI0mDgGa4pZ0CU8AkEv8XPvATpcIbaZnGwS6z8epan3K17y7RuEA/mkV
ASFV4gQVvNCVIKC8U+M3dZ1W6qgoSUhxNsMkF2DKr0ROvWE7XHg7QY3liebn8Axr
M1g69732m83S0gz4Ov1LZ9jen4GYvUL2yVh3scdjdy7Y34c66C0z75gyf7ake/Qq
sEOxG43UmrbVjkPlLxwgz7qM2CvPYC3u54zt9zLAMq68H70Y9LfMAJJTUElzJN9p
IgRwLo1cKgqdXxV2sexw96YugpvfW2zufvJNe9lpkdGhRLmO5gRT6qAvikJ33j+Z
9Fvk11rOAyA4byOTZxvwYZF50vU9HHS30rmxpZ/ls81fEwC7XH19H43IOYt1p5yv
0s6yj4Uq6nroCjMJxgvVGjezwgfu5PLe6FoXt64eE6jXW6CbnBonO/U65nhqD8Es
OO5uxcXcaeS173idOG/z2nPQJd8Gb9rmxuhp5ATW6DQC96OW/JbCKIjv5iF4wq5b
hKAz/ADrqvKkLqfPjU0tTS10blcemYjDkLZxfLQPeWEwyiFpow8U3GlIXKoLV8az
V4jJH7BLND85BaYZ2M9uwlD4fxVUtDFBpZcppJsc2zk1CBjxay6SLtUILAfv73Za
BX0CC4kC5w3s3L9rMQE2/T4jBGMh1VdCfECXVNMpjETc8bwtDQZhj8cAGPx9mo6e
UV0OwyHxoRQb3FTMfeCOGJCkC8fXeoVNEqbCDCHPfZg2h6ZwhTS+Rx/BF1UDAtwX
Pdu2XhoNn8wJY9T9Su8j6hyUGho7Vpc6i6/N1aWkiAHnNBYJIMevTb2w+FqxPl/O
/ZDc81ZWpwPqw1wP3r+anubfItj+CWckpaPNF1kVfVsGLPqDXN4EhiXwzxHHN6pr
NOCs/8r+Fl1sgsyGPu9Kuw7qzyxpze2HCK7N6kOBD3asa1k66ePMEb0O5FyGd1gN
yy3SBvqavduFTNLBL8hUhCT11D7KIz01KotEuK7PLpVoXcrIG2GeMgadSrlM40b2
9SYZ0EdkBWcnWRkVebDJGAsMRHrxeuNYEm6JgeKYN7Em+PhC51UL1cc5NRk/wICK
pxZIqvhinhqTcS3mFQTpoxfJoTAaw2lqsHtiKrcjOiubaw194l5fHVYLQPhUqvrG
IwUL5TprRDm8MJhvwjha+RdalOWds78rW+EML9klmHu0RbQJhByg+q9xIfFCm+Bm
9zQc1hnufBEFZglnB3Eiv0P4ZWpB7f9GEoaRFRAcFA16UkBU4l2z2G86dQKVKizk
nAPoRB82uGAvGJCv5CSmIBQsoX4emVefqvnN6L9/QRI4HkuJOBkC3LZlwZfiOwrw
uRb1cBAPEYNS6b6wXy6unNxTtqPifIqy0I0Tr1y5fDuFFO0/GUBYADvt0eFmN2Gx
76i+1gfg40YcO7xDCT98qGXljm9pyGxCClsW1Ez+GhAdX/1z3sOPIa3T803Mdo8a
IuZltqy3eYyygewn6A7Q3XHJiSrzgb/Xa2vJf25oQkqudBsrW7iPN63rcj3VzbCp
eWkdzVhhL9uffcEhxDnA9WXmyNV6EFtJVJhXH/nq5MPIarvEHwIPVjNT395dNlXE
Zbf3mXyqr1cI55uCkGmzFRWe/LYcKh4MnVdF23kCaiVmU36TpUyMLlvfylUQDXVQ
Hpghxr2QoVCGb16Z9FCzHR3/QO0P+Yd22bTS4+Vl8baMspmgHb/H+GMvJQ9ozr+3
U0e/hhvuUvGvFSAJjCSfy/pB3+Own4iPuB7X68usLKxF/ZCed04lPnHRRLg6DDCr
zIp0E0IXuv5pvsRBhwRR8MFZgGb4L4RDuzThnWhup+o7H95qHMfGuEOSHLxxaA+Q
d4U89ZMSwFwvldK1kOFDnBSTiIh2U/PRwKL4or85NyAm9D4AFaWa7tpWMdX67see
6MMhbT5rwQyWOco2C5xVLLothpyyKlj6VhqMxnG26JQ7LbANwt34qygdMXyTsaTj
PbUWpF23BmgpjbT1BUueBgQqWdrYLWnBug1GVFs1x/Js2aBaBsXF0bZDbucElNSo
8wwSvnDIt1k9cxtjv15v77U1WfxERJcRcJj16KCRGjkiSPeRWek5JEm0Eqgq0XuW
0JEy3Bst/b1DZifxw7OMCSBtShP65XcsOdihXIbnsc0B5gKfDc2ApaSAjDT0lAsx
rkZYGzoUyXrcC2O0Xv6G8bmd8y3SGnXy/tAb1kEdZMoBFqBukv8Rl2nD+5eQUmvG
7xpddAFpCKaiA+LIF1SOJ0DFbsKkArD6zHcw9R19PbyNf5z4AGKe11ywBg/0wx5S
qeM3K85TWmiHyLg8WIWAiBZPMP0WKor7UkCI+V1axzTTmEwVTQa3cLY54vMSTl8Z
LL8EY2X494Ugjn/azKjiyIY8kX3eVOd07hfCHtNI9S3/E7MdOk9t1u+89h2ed59r
zEgULnQUAhh4vXkmFVdVbVo9sns23oLSPa/JP8kbAYivLN0cfvKGTvZBzuLBLudi
sgT8cyeFMziu6K2823+4M4dIfwGJOiNzuymdS+s80xr+PRwrLPiMTOi8a6I0ZmFH
8ub2F/PeGJOZ/A1WNwKZA9L83c2CBam9scOzpMvFu10skxij49hi4mkF1+7fWZB4
VusniLenMe7OzwoAxFgoIXN0E7mikG4nDdvok8GsYspIGXwSsjKMHW7Qf9MwgcDy
PwyGUYvexoeVmXaG7pIakImjnvukKlF8tEXdZzuMViOrq7KsZPGdZfpRsiqW6GnG
Iyuj9mG42RujAvLnjCbVEMf1Q/cL9WDT4e1YthHjpXHu7R3rNVP0zIFHqjfQhAUN
E2DwTFmyIGgTqdEpi7WiEW15tLRibjDq4s3x/BlLhZ5exThiL5kfdv9PkK4wdCWt
QdZFn4KGG0TwDvdaa2L/IC5hxbvooZ465psBG80XZYVJSWkosg5BIQaKCMr5Eawt
UfYV0I800LumIZ6NHcV5WHIs7wiVWXAE9uHhf6BpB9GQ5oa+jr58q3EtS+SqhhNr
L9cDEeqrA5IZm/cBSFMLgDh3Et9xfmQtXERvgkqR40i3VlqHW7VsaPg2qrl8zVlu
9I2HbETnC/mjU0fBPTNbwG0uXWsvgXIxIGYgnDy9Qt8u7gtkhhG2/LVLd+hGp/q2
xovok+nROi9wssQb+1v2NNyuFs2FIYoIn14I7+xjZ18UTLM1AbKgeUYZYLA4N1Dl
FNu5WwAjtnYsB8OMh5ZMbd9wCqOJrAj3ansyKhFRydFc/gv1iLfTx2/Azc8tc6bX
EqqLd6j/LkdZ7fS+Wss3goRRoW1QAYWkitxOv+d0jqpEKNob20VAh8kYLWdIjhmC
G/NAHs1Px7UJ0h4dpXbxDATUyBMWQbJ2Og8t0HkAu7CwO7JayqE0ps1ISDzhr9VN
J+5XmP1HjsoFfLuCiebkZzKRXoGv6xM6Ua6dtBagTNHtjrqScExIRRu3D+jDj7Hb
IvYl+30nJFnYV10v8/OJfkrH1Z8LbYRUx7iR0bDPyO5xCPkW1lc4oCU4yHTW4KSN
LMhbutmGOVO8YYwWrrKZ6nY38CA8QAp2ZpDWWA6puwtiAlP9BEakhtqasjXWAt0V
zVrXu7cf1pYAW8GLQZBf1nmFxrXcr32+zik3Fdjile+c6T9DUMhHh40JSFukuz6m
vwDbB2ie+AjtBM1boJgS9xm4bMIXpR1ZkGaHD8aQy6V3V2hvvr95MgBhLgFsCMBm
c4nn24/JonHyHHhbpxBK1XU7KqWkSajQ6ATFqwEtaMzLOvC3HtbJ13K9tbhwNX0i
7TcZgqg1JrQjeQU+SfX0CbqGJeCNfzX/hswbhC+AkAcrbmlxmph6drA6XuwMtx3w
rocGF5SOfWqPKGt1QsHwGzloA+07MHU2AeKQW5bVW7CWdfQh9h6rBvwgO4tC9fVl
6BeQ0HVTjjfEQP0u6AUbj8+FvesAr3SQ9E8IoidJJWixDsvtoDk97l8kat2rVLnA
kCHL4lgC2MfTt85+gsqrTRU9mncpxiCA+TrfsAHB9kuejPYdUQlSbWFnSJ1mPkQs
vPV0p19g2JiExV5rwFZMFWXwI55GNwxZt3miQt0p4176q3f40lyo79vy0g7cB6gO
1z3j9Iik4Z0NhDKRG37ILw9TYYN4Tf1WiObYorQqlohI50A9xnwPySAtEtI2PYsI
756WO1x8cxrIbNuyfD0yTBUYuMoJIj2BZfoAm9fcGqUwUIfNHSJr0ini1AxLi8ca
bv0Akxb4SokcAJwbYtHCYhHxT894a+YfZzSKKErHG38vqz/Ghjo9IgodIQ87LbUj
aWX8KYzEy1SQh5eASYAUSdv5BrtA49mkIsjJkynmpSpXCNdgsgdPt4ZGvQI9VZey
qDHn9iBlK/St5qEvciTqdSkOMEuuZE09wfbQq9eYZnN8AfKxpZNh4xsiA0ibR9Xb
N9Yev3zg0P5Amy9TLeanrrKE8h/EEbOhRtSRffKz1/ZIplB3LeO0dLVC/CBM4LJb
STszxE99Pw0NGPSyGtL4S3HfCJLMPzk8o7GIbhdvSwAqgRW4by6dhDdI+XQ74BGe
mCv8fLEo+eKOxDaIPhoSSLiFy704MTZtV07v1TeJZ3Xyk0N8j2ucW8Sk9Z85syKT
H02womWWabmqd8aLvXjCLTfe2YC0aYqcevsE7a5pOTmPOs8NwSwE2iBDtkyRwYPd
Vxge9ypoKT+9CoJxKzDOtHITbbccG05nLX1td7mup/2A7ajhMxgnXvGUrtUn6j89
v0eeSmM5pJbLIrG0RW6+1jjjSt4Z3U/p38O/YA8Rkvk17g36M1+qt8of/sBz85un
ZaHQF181hLUiBwaaPecqrbX7i56Yt+n22zqFSTPhBdEwpyRuyHfxXv6P1h4eTVSk
CUlBccvPvkspHeN41b3xoKCLBS98kwZfG/gD6OfLoDnh465HElwKiv1PLweVD37Z
mM8KT1onbMARjFqgSSHVCrGLhAhbWLtnUnH9xX84JzSAD4RVOQukefCBi4wk3/LC
LeKo73xGkx0VTgi1X6VNyzP608Jh6jaXKc+rV3JU3SfqEB32VYPLReEOUdkyMUi5
vvSnHDYfLxriEwNWWllyI7sZyCTw4X4qkm+KIx6jKNQNESXsUpl2CDtvzgilo/DN
tnuBhD3ZVQPhi58okcWg1SMf/UESE5dCJPHwFW5XPkzr1i8b/pp6CrmJV+dz3Q3d
YT0kdyvHsF2SYzFaGkTdJEyfCscpbmXrSePqYG6Yk7vEwEZZ0OUVcBoFS0UtqOJm
pHkw9gxo1rYt9HmW/BD53ykCSuFWQHaGAxNIeBg5LzcqT9HzssC4ijQPNM+QJFuk
UVlg6FE06fdqMUCiY1dXUyG5QBc4/V/PPXkCno9mXZB0QOhBWpIEis0fp3Tgngs0
qoeqV9UCKQWPOP6XLg/ss6UpcH/sNNqd+MEyKTMoXnuTKWQAOmklyI8nvmw0nkzQ
SgK2yfs8cTxGLXbKDF2Hw7JkvxaBbxvHvwDLxd9ZcBX9wplpOaJAgs1/RDF8ffie
r2Fl2q4fWzDn5s/Frnx2JGqJD5wpULACkSDX7kBdjdIXEZT8lof9lb7qBE7ALcPN
oC4wPDX2XxcmVio+kYYjtH8OAw4ILNj6bgtbAIO70rap2/hJpGiBImALcUBd6E9g
cEmwoi4IYNMy1UFLXJGp5Yc7CHKhX1+Y3tGpzoRklhp3d7sQ8z9VN3p4iJIQuOoB
cpHhE0IMK5qGsaULeiOey1yvndmuTEOibSnEGl95g3ioZq8wkSlKoZBHIQgMINUo
x5eNwjOmqa57+hEens2/e5STXJRK5me4q6WrmU+UUSoh0hIJGyQb0z4rHjweAC51
7QeIkC3zrl6llvMf0Xc32go55Pai8/I92V100N6S4+x3FhM9OWbTlsLuw9prt8qQ
TiE6PqnN6j42YDzUSoPoOdbOB0y4QXj82oCfgsCi1b6y/xSO9ZuBlfexCmtCYFH8
CLVA9RufJkAvz1fbTp9dgq8oT0k0V6LRCAgW8pxTpgvrxXC/gujaY1TnjHTOshgr
jt4eLmTwkjvXpJssLP2gWfwPBLkArG3/PwQZ6yizc4N8lDFDFv7xMZBaHkd9I2CN
81AVCh8ixVQ+0aj2VSZ2Ou+iqWfT48u+CwfQBmNrYOm4P6vSzgoeJATTQi8sftr0
CShylzeC9iP8ZSdIHyxRwHbJgxxtCOSU/FEM15XXINxdkdy2toMo4Gy02olMKU1r
BCcM/Q/PiudtqpIjrlv3EHCCmyh/tytFRC7w4/P0lE8Vdp6AiTR6YAThtxTFtk1j
I8RNrX4TkMLwZlBjHjEegevYfatOoPVKNvr1lbD7j4X26s29qViJrqTno9Anpuzi
ZXQrfLIwzlVXNrdru4XhehCTCEOVmYZVE4jwW8X4hL1Hi3kIedH29J79z7krWUIW
4qYnlTS3LSDhvcpK5ZNv1+dmlgBeKrAVWTc1cMY+OCT6YH4RcdrfYAGYwuvNq0Jc
zDYvmLN3Ra/60tGxD31vzZJqwHt8OKuetZiExaYMgryOa2yuOX31NPxGJgJZVS4P
uDONo6mdpv2g9+rgBQCeEkgrv6nQBNEPaMKjktvIwgErSgTGsjJGGjVdZ3ONRKx9
fMNXv3QVPiqnNHwfDqfyw6zaWcptJv/E6G28wtWyA3X4PM+MBseYvft3gCHG2zLi
86yUIyA3y1pw0I3uv/exn5vUEZOh0lGgwftMcA13Kj5oG2aPbjH+cQ+HBf3xyTqQ
QN3do1K3t5fKYytZ3RVc8XRxqdy+tatna4nR5tFYEjkMpevbJ6T4kh18lQFMgw6W
4tRT2Kf8KjW55aB+1x+tYHema4+qbWtSUcLutH9v5Midxk1Q6JBT8QY6dYGdgveT
aMEtULPhf7c6w8C9O6xxEFv/NJ0ECDCCiJtdHPAyXrIfeIz4DiAFQVjQiH9vWvdg
EZD+nkH2Nr/M6ldql3a1Ozy7WN4H++Itag4X6HTdhdwlE5WeU+DuktKzIPF2f4GW
iqaRd8az9Tx8v81zAbxdVVPvKl8u/fmt2rEIalTDY+Gpf1Liaprsxo7apBhXz/pR
vnp1bOEvKs6BTxdmA5i4m32ZjJ5SiudZ+DXixYaOZhoCSrc4w3fBsUQOlZLEz7pO
oGBCIxl3tl23xNwKxlvwYa/9PgziXXvDcPOI3hI+v/q/Q00ZV4sC9OoueZdAsClE
UVZEKAdq1pqK4iKMBs+pu+ty60ibzUU6pEFwvvAQbf9CblP4yJz52r1S4ztwMZIy
bYPyLYQaJyf5pOh0D/F1OiX+5p5P2yux3v12y/gx/Bl+5rvtbR3YvvyFLXDb6Tz4
CwJtsnlzXGjv+8OiGzZdhv/3rE2TJ7PLSyh4YHHnsWwpxOiJ/XQm3bM0MVNeLsz3
6k/uY3BZNhwG0NFvsPJO0ENBKnjbcIvrR1UGpgR57SMdT5+XKjeQi5ACLxDjZ3XM
a8panHOytZIi160kE1VnkBpOhVW6KfRJD54vDZu5xkNqTFacJQqNgGvKDzRBvUCw
+/GxOAeNzAl61scfMt22IJUo5/GwFkJCadK4Kd9qmxhUgRliP/AfmrJmyOr0ie8b
+40oPOtckdNJ+L1Sp+6PkW2c2knLd3OZa78f8NF4c3jRSINAcxidWV2mzCXTxhVZ
ridmTK0gLcK/5N3jES9yUdHXDjaJg7hnPpxAbYT+CZxooI/ocr3Syy0Dt4v4ZWt4
SxhDrsknTa/VB8hXje/0KSfTa3orT6tLE6/cwGnQpif93bRN5fGAMtVcULzoOhAq
ZZbjklk3Cib+kqyU9mw8uf7fyJ2hx9XqwFdkDp32evB+WWzXNBC3J5j3fcfQgUWa
0mC33H47HcvEheLvnh17rccnN614Zh5D2h4ykho5AFp8nrkUTi9WiAsEQv3J5bw4
6lWMl9u70xRtM4pnw18rdthGqVL67ByPIIcsmGnEpoUfDOkDz8leiIk2++84taGV
i8lWqVbz2xr6tFGKVPcKgDVHlN26uBXxrYgFzy7jPXTlO+o0ULus1KNLszVeD0kx
0Re0kIHL5GD5jLF9RYCLvw1mB4oHKKn3ivi7p+9MubyZNbGQVoDq0FhNA9KoH0Yu
h8opiGRozEhC9xumsDiQrrC9X736ht5huXkWDw0hXzQn6gCWaSm03JHQt2WnN4+R
/cVvzqPiUN0ouaRLWqp+ZVckFqBD9PkzJXwEJmb2dNcUflfiOHJmBEBjgnAzTTmR
XF7ZYHKNo4j/7WdDX0vl06bVnuK7dZo2gNtyFO0tDnr4n8Tb+n03fRWNewoV0b6v
/n8N470fwx3YEaHSNgmH7Q/xkQRxq5J3v0+mRW+eu0IqVhfLinWRAfZPvO/WW1cU
GT3Oie6dEYxjanMNNwXsgRCa46JWnFm1wpnT7i5sZB/JNbBEfIz2sZg54/bbVMjj
yvpsU/gOfWGb8qzhXkXT2jW0d8QTzCraJuAbAo05huRUiFrikZcVwcLtHZzCCzIi
fc98igsYrKMcmr4xtaKxq7pH/B8yKAd2aYeAG3OC3ohsbCfJZTrmKyrAYds7vgKg
Y+TISBnbTS+0G9Vn4V0hdz/yieu3EFZmf5q9XfOalqFf3e/9NY1pNqvqPg0P1fqj
WVuEKuwd/YRFYIS6GnvN3zemEoEpYYVNEtzweKozjNC/MZf9Hv9kz/74Wa1xbn2M
M/SpOXDm34oWSrYEt51oup02Hz5oq818cnsOU48xLo9tqy1fsP7OLsocpUtYl7fM
1szFGtCEqwcy/+y3cANVimWRWbeey+AzwqOiecpdgmi7MaVpatWQX6Tw0Rgkzr/p
Mr3Mn9yPIUJ/slkCHlIfML+mupQuXHqxE0cdP2UOKLG6Hqmv+C9fdnV30haB/rr8
SW1WwMDRoFlNmEw2uQhjA4uovu5sS5O61UIMffjqJxgL0RWaR1u3QZjBsMYr0sL0
Z62iTj4LuCk8hqrgZjACbEjjumrUIWeZ5Gv1jqNzshTRHthvvsgeDUk7WdEdAFN0
NGrP4LR3veshQv70ZFvGUh682Xr3nBfZU0QL23YKfUXg4k9WvTHvyg7GY93p/UkR
U3WXkpiKdtq7cHsegF8kbQnCpurGsCEDehnpVLJ5Yh+4xDISqJpJL+tTn3Y/hp4r
qyNrznOQ9V/kSDN90mfbdX2/2Ddp8AVNFrR6+1FgiA4O4l8tj3MoOdn1lfCJ3xay
RdxlAw64iCpf/B21rE23DXgc7RVvMbtNPn5TXfNf8Ie7SKcx1q06L0m8T5ijPRQ9
GG1rBvn4UV5EC7K0tHt33Q1CZvDT99lyMAjjMIY38WBsxyMbqKHaz92YRLAKtWtl
QcLT1MnhXEAzLvn723wEyfpeOtU/IBITANBNTDGbQjllnVhoAeiOi+5Ft8yEtRqe
yMh3amWniucD/tjFSveDQMVPFjhldJWROf2vZMJJ+23fvESya+bSYq+dD1EWeZq4
ByIp+yAVxUxZ5DJeukd9RY6l0DKN07uptAHRzaeJTRPfwLB8qII6IYVrACNOUbaG
d2jY1QwMNmmHNqpUIl+sSNAINvQh9e+j7Y1euvuxdkBvY3kjLF1Tgn59RdKJdiT2
L7jKA8JmV5+7QbyXlNaci+Fl5BoR7pL5Dd1hJPiq/LBTHKuW4sREChg3UPCMDuwv
0uksQr8O8D75CT+9fQOcDGAzBDV5PKV54eJqL7EUF/jFL/D5lQIU/kYGKH2LE25L
56XBO47hrWNvpFZUfPeOEI6sPyO9pfKRNVCrUVRXRZCBaqGVU5Aeipevp0V4NLQg
7twhtHKlGgu0kLsg612NRcz9wBNXMFvQwS2KIlkwA4xF227d3W/vfoU8IMLUHm+d
B+05wu8/4+NlaSk2q+gnQpHFVxyQHAEO57rgC0K7q5sIDiTcCXFA29UC9163ppRo
uHTqBigKIecSlceGgDpy7+M2P8RSx9mH7witkxVecu2sBYgjentxjUR3wWsWq5fa
A+qwXFsXs84PrBvGHO9d85V95qXbnUc+wmGzPxv85K1jYT+4wo8JGGbqPoaWQJwP
dVaXV2tuWu0rBQiBy3BRM60M5vpmSLol7NsSewz3EedAN9CTxZZH0CtvWDErwv+b
gOsxlX3YZSTOUexB8wyxmOlpxyqDs/GtBetQgQOFm74xN8CbnZWe58iHrYGhcjzy
14uhaGGHaLkzFJPAMk/931nQGqe7WtNCu5OM0Cq/GmVRiug4AgK44HsloZ8pxmdp
Zba3l0Fzo6Q743un8Xvr4sRmTW4OrDlpGs/rHT2Y20N/EpeYe14IbHWpk2jQP7AX
T5+Nw06YuO78MYNPK69haWuk35W7lqoUuhWzcCWUEoqMu5qRZZtS8ogAzXK74klM
TFKYE8bdKwLoQ2B9KpdocGA3E2iyurA31BgjtFqGnixEDLm+pyiBjM/a/G1Jj6dR
riH7l9RAFsHPx/+LpalGH97lE2gFY4rOgRaMGY75W2qOBAFI27Ji/4mUowMJGbnF
EfGcDWl95nCa+pCPqUE+83aFTkuKu298NS9Sl8RkP8rnNeUSGFLDbacNtXPbcSOX
D1J7yGROvk9eYCCj8aFhPF/Jqd+pI75hD+PaUzzXkO8TkiIpPffR32EVUX6wB4eD
erhkSxQK7vdMbRSWMRVleyzCY8QO+FZCNitkmAhT8k7LLycc2dxGAAitD0fQXuzN
lFpBtP3h2YPL6rpmHoxfG7atC+rnfVatTqn8OMeVk2Dz6k3lVOD9K2PngafVCOSV
KryfWVphVKXLeQB/+78Rvh8mhGnziWsC8vfFlL2+Z1DRlu1nkMum0RGk1iBvpkT+
Zg52sXpWzNNJF+lc4BWtnQaoJlYM1xPdzfAFDCA6Mi7DBS935reSmd5rCUblHGkj
WUf6MU19CSjlvJnspCKhd0zh1rLPrgjPBaxBxBIzcM7GvFianYR2knTRl4X/KAyU
wO9mvgR9ItfmiXq+k+QDxgElhXWugiizkI08qXSBRWvPrmBnI3EsOQBdO2D5sAzg
MOGtRh8yrO6DS6hA4CRhk64IH+1HN7s2Wu9/SnDrJsv8X9IBGdP8cGjQi865hrW0
Vuj48Mnp5F4ImgJg6eH/Eq0cm4JjyHHtkSKILYhg4176hjP3fIisZ9h0zLAGAZ07
aYX3VHtgbSxLvIIHZFHt0hlwoarRxXyHC/HvSM4M9exoL2iWRXKTatzreOqr0AoB
fZmV8bOGiueZ5kRL5EQsEfLzcPgwPmpQEWtxc+4srdOavacdVrdQ45znwtW9Yvzv
RQbX12WDshsN/C7Ff+iQxgUYlK0aIlMdHX3+QLxuJ5fk+d4PdFAtyInPCpR3cLKV
chHUOJZ8SIhgRXJ3wm9Xe0spVXk8XvNvuxsEkxPOXftJYaZBoBAvkpCQpNSDAssH
A5rnF1Q09J+L+eT3XDAlYmJ190N6nSCeVtKpDgwOl66mfchTqDZbu1sXqw9r3e7L
dG3oe+HZUPWwY9VMlWrVCQw6EoTGfxi9e0efrtEVomF13FZtwrq8kUocJeyfYG0m
EScivnYtK8wnehiE9GzChOp2O3xsiMbRRPKDyclReTXSNi1fmBzJPao3hkGYDM5l
QGjad23Sxsx1IIIlb3v6OFF0hALdcsMKRFXFUyFeAZ7OHT4ebgJcokks8XQCLeas
WwClb/FMo6EYhWh6Xs0wV47X5xPdG7iZJIWbUKwgUBtfu1MV1GcoIfKQDe4kWrap
APZVIxwP7SBWjE9G54s8kMb4sevPO/1jhThkwvcW4ZHPtIwBybYVpFoZJTjaSCPm
KAF21t6cLhbm/rxAvAopUWHgYXmmnTApVKn7fJPFyuBfDzmEYuaphm/iaeiNZSf4
ouhD3UiMrU45ZWiJ3PqYrTpF0jvvWBRRGwon2Gg2/Vek42zxSBRopEdDCe4s5WgD
BtcoSXG9jJD3lEgG7zsBKMVDRODrCJ9VCkPXtYb791S3ZQY+fgE7oey9NqTTkm02
ONOueZKPvCjkWXPG0uAEomx27iBrvFS2aoj2L7pcDIiwkc2D2ZKFv11N6kitZcnq
1PjdD3olCLzMiKDEv72q27NC0EDoVMUe5nxDtLG+Q64Yrku6Dqu6y85qFt9LDwdn
GZvv3+hil6KnFn15T5Y7GX28E0U/8PUQfVQ3QfQUQVu7jlp+tPtjEl5JJkfte7EG
5oNZzWyxu16k5lT84CXzfBSdAZBRw59eaD4qdi/FyEDvEYtpKRByEVisUrh92SOK
gxkIIUAJKXYZ/HTl6G3Syx7GsYeMRh77q/1Wc4NRVFstVo1JUSFQ8Yw7Blz/cBSY
sPUWIuWZuiHAGGwYK1yrUwEiHq4vIBwl49iTZFndAbOS57hvNyQD3DhXfRVcszhz
qDQi7rFzdZggwJ09A3Su1UD8Nau0bhtF//D82qBnoUalLhGGlkagMyIyIafuupSy
zBobkFA8nu+n+LfTEftPOnMGfL/IvX6AHlDSFvOSex/z4cASLl/5WJIA9x2gH6SX
4dvM94sFf8trQPKRh9xe6qxQOxr+IchTxLAb7PSbjd73K2+OnU+v2oCpeaygJ3jD
2PF7/kOlB/j9ZNH6NqqP+LADMj1UwTf+zjMa5S3dPgcWjuNTOHqKta5zbLG5H/Kl
do4mNLAeFwVglNUB8z6pAO806iuvMnHQmf7wHBcddGVnLTl6vNRq7aeMuDkmmi4h
dPs93QfLfpu1raCmisk7J+Pgf2Ozr4hLyw//K7xpR2PHF+K2ZDfS1sGASOT0nhKO
U+t44jtFsSPrnTN567MWacExbBu05sx5P2S7yq8WPMaqDqeLrfrsWPa2cNggIUwr
UkTBqhDdAzCSMwVUo7fMI8XlxH+0OqtL4wBXMZCf3o4DKo8XBEaalSXlSWBh+oiF
m2WsVgxqm9MaPcTxt5gS6cZJEipMyjM+MwcilzQShgjOwkHS/9/aKZP8q8W2J0iH
WpOnqi1/kcF6u/rzJqUzStp2EwoDZuEmD/OEYms3XVE9OM7zjrSPxnJN19bnhiR9
2OHHZACLb8zk405oBU/r0QySQmY7bLih1ldloW42DG0NdS7eGNuPgUBkeOOJOaBR
rfQPh7j30osk1GqRkF+hJJO00ccnY1sIYZvrr4Td9sHY85apSifirXYSH4qjw2EM
3iPeWEgEUHjdvW4wPbuYSmQA/f47zIaIDgcfJohHYjlKXfF3ymDbq8OVdoe4kkOs
2tilekGdUq0R9k1f2il00OerfkI9hUvTU6zsCVhI5ZVbc6wg+El2fSztlkxNROXC
smvhW1qsNuZ11iymEaE9XS5uxkPktpQqlpNSMqExdPl5t59F4TREs9uWf72XTuQz
6Gd5LiK4K9L2hz/vycTj9nae/L6Otm5WXyWggVXEyGXAC/EECDKov/hfPc49wdh0
7cop4OQrb1UljlY+/ps0U9YZCAaPZ3oKbx8IEdNFVMlNCCYrnhQQUsnWTMR5ZzEo
IYWwK2z5Xg7NyMubB+MmHYDW8wcMT8o2LOyMzxCiMXxRj6ojaO1p6WmbyZL5HeFh
1sxopScjXVELc+6lotoFghhGFm9Ba4QCg9FA+USpK130dlkvBWFzSEJ81rH89aT8
MRfhyLFem8blADZwbQ9qSIZ+KR8kpJaGctvYn6TyEpHhj4WAi4IPpvrZgJ6QF4ft
hv0cbKKeUPhQC2Z+m9cP0lKJOfioJNGYYKQ0hJD/KIKmi4NcSIvGVpUG2dnwKNAB
P7lFRg9BBFy0Hvv0Y6o00Pklek+TPk62gyfwtVDsp9ykahGDtZBAdeJJa3bDquQ5
PVV5TS23RYuyLi9FLAwojnoljiKvkVPcxjA8Dr+/53USrljGAUAKvR+PCxAB7h/j
fiYmzSxS1oO6IY+3gpJ4ATEiBpDqSrYB29zvOPLJe+J3zrKRpfQo0sNY9oUyYM4d
gaB4j9SooTFPejNAwSjBAKKxA7C1jv1/2wswb+uKgtQWnj5qOzSe3om9OJCXLHcz
MLAdWjYk7MWZfsRwwzh6vdeO+sPS3EEjvPPPjmaT/tcw6skjOPg9j0ps9Cn/o5BO
MCygOiCony/VNssF9n15J6GntUij7RSdFCEV5DXpZHqt1wEnUOxD18jbP2wKGDlt
vLz0wTLbhrm93wuvFJcZ0P68gj9QWhBrJyoVhH3LmUmBN4dsf402/gQ8WRnrCB25
ykDL1dOile0Qn1fleWBlD8QqmzY0yFRD9Qo39L06dHe8YkLhhsWK3EWLmU0TgDXe
W2rPsvdn+ad9wEx9sUeINXIJRWowjGQoOIX5V0v3AeIx2tbx8r5DrQePk4CHJkjV
oFlrKDdlVCRiPxm1pR5wOiw6RsmdhE6DN39zXcTCOKrK0ISKnXuxHBMUiAlGjYYQ
vrvgsMfsidhLhTyR7Zh4779gbWsODiwWZ9ccgqyFGXx/X3Dv26s9JzoN1XH4jEr+
C6mluZ9TUHqWeSh6bL0wUfPzVlsz3ZAwVz+0ghn9N4Zk8BBsUQyl0sn0jFC0hOPr
QAq+AljXYNM1CJl8XfuUVsBPubmAZ4nu2SYTeoSmDWf8U6jSKDKA1NFAcKCf1TfO
QyPT19ihpLIQceu9ZTditSyx/x8vIkyvzGLoh7v8aZS6nM7kIqH8XDqDyMRH+4zs
ay4v+NW1tT7+KVa3YzJhwU/uiIOjmlPdGk2ZnjfqQdmJSJrcOdwp7NZ5inQXkhHi
rRwAMeljeQoqqGe+h7rP3nTn4zXhv3V24/X5pbyMwJzTqNEDPZ7b4Edivw/qhW74
Vi1sGIapo8ub0cHKZ1nXOb6YABbqa0Lq1tIIDui3D07/b9RkpTQOVFly8v5Rmm81
PAlgESu6Eka6ZEtLbInKyE5hFHwZffNu3L/A5jl30YEaJT3N19+jhH2TtM6Y3T3M
HlZfi2fn1PBLmhT2DQ6A5Fi9N7uNCzCtYu/+2xN1JjcFK/jMYk11ZXnUKp4FsPXX
l9ni3dwEVLdw2tbC6rV+rcCieUzaWVaQfbK556+oo1pQfCtzNeBbva+HayOV+Nck
L9aEPsHdF1Cg5RpaxGPo7uIjuacykIFIAGncF1dUv6hz3o8tphcfTe+rCAYJP7K6
yLRS97f5LJemuYOEefOo3PCAF7m5+Jac1woUzlvuGtNpJ4UOLGymy1ngJcl+e5Yr
d24lgjnyPcb6WDhXufuc/hN+4ydWiwoxi2IqsP9LAUa53da++xEh3R20JmRdEGSN
slJaaqesSF11ZmSuHoE7ppORf8VuMZvbMGwpR/CYxRHp/gHjr8edi0/1jug/s1R8
/7pk01yiWf3pqjSzKnbN2rtA8k2Gf3cdIMnivpQcXhAP7uWyGWAbKbjR5KP63NZZ
ximCDT1dahh5pTFLAWvxDI3zy5C4TSCl04wmz45S+paK4vg7Nk80pitdJpLi+bCi
vrUXzuNxJKWuzudzemOVvtgfl3uPConrttF7q1V2nr9Z2beMfWTzKlD2Mfr1Lj5e
fbeOV/g8v3WtGv8O9ew+ixoSCOLp4/LEYIz6Lm9f55rMj8ugaIzps/wvgpGaR7Cg
rauZtCIp0N+aYi6kqjb0XIMujKCiHuV7iBxQUqhmVmZCWB3jgqz3z/MXMz99qiH1
YjXCTGJtohsqlcgH3rwXlLFGhckskn3gZ5AL2xr0YJfDnxEXTCgqCq35u6pi4zKo
a5KDEyLhkmjlf9w2OE3hamxANMjIRhg4TIIvY3yxTsyJWSNUzmP0jzlBrNdVzH6a
uaPWTogayU3QSs/E/C9t+qqM8SAshkf3v9m26YF3hfCVyIJkri/RKSmWtUPBDUsF
ytYh8TThWyhREtPl/vp00+qUasAj7nX6OBooInQwUHp58JDj3JI7JOLMHvt/Z52t
q7zGYJynL/POExo8RiisrqrUOOlNp5l0/bmpV0pwviK1ScoUw0S2hAXHbT2INBb7
PwL3f2Y5g/pdTRVqCkpZaxXamn2TsjIF5N9XLUJmUVPdUOLJaa+fpL4eOxk5F9Pg
7d+Q9Q9zQEBCXqYvZbf/pg3N26ONPiKqZ42r9bblW/D1rAjq9t2MDN1nGT2Capv7
0sT8UK0JNrpMeC9LpxJcf42JTdD4din9t4TRiKnIQD97qr6rxEBPNJ9b8CtN39iJ
iMjTol98/+j82fpYv8p/9Oi3OzaknLgwl/Ante4NtW/zJ80FDDVWkWPBgPtiZypu
Ltv6xIOsgKNXNgMNYYZu3U7+b/aAM1V9uCml/VhwyEFyxwbL7g9YWCFizbnPQrXt
3FJy6a/hxspdc7rDXDA088EQNEk5fqXoZKZVOr2jUbxskKROY1ubOltU2mm/L6S/
Lqc80G4/BGgs0IoY3Y0ZDPHAZeNPnCo/ets8a6mQaNSV45JgPi2fPPVjF2uDHRa9
NjTpVnh1HIE2H2BopAuGN5K0/par2bvojGk/qeGtNfgkPi9zqDNvJF8PVMAhCDbq
JqY8fVPuUGr2kCdmQNDsBuRkqPG5y6JEnNhEpN/g5WiJz/Ey2Q3/2Hx2Ph4KgoLu
HxXU6aFfE2XTDJmz1Qo1Tb4fsYasS0iQrS2TuR1DQc3PkrVSH/YoV701EGiePoCB
WF3p2pmQluiN81BVJvdQc4kYok336TSWHRpA9cqvvWPolksTPXGj/u0dlZm1SdnY
Xgw6R9HqJEnTXhipYp/9Ibm2S10vR5WEXCMy7YgXT4xSU+YUZfDlkbOAhRsqMPNz
RbRl8t0Q4KksLQrWhre5j8zaApL8chIh9GeHNU754InQmHV178OAgx4kR14A/cmk
ZIVd/C3igFbuIC/7Mcs3ThAXddGII7VSa1etOgW3Zyr2pGZ5sbwlWJdy+ljWu4LR
3YighntosZPJQBH0NdMf3s2ooHQQnkjInin6lgI4mS8RKjN+HAw8HWjJ4aYsX4CV
JyNboEtcQS0GMbXjLSeipwJoKOOVwpjn1TIqmMvMvL0c3tM6JiYR12H08OnsQCjm
eqg3p3Bm3RK/kSrz6ceOcv+2MvDCfbmRspYgdDvjtzjJrw/Qcqc1T7cK7HBJI9Lc
FmxMUErAwqsDI7DiUGw9Kqe8kS1zmKoIGoJX3wAIMEF3iPGXB6OOueiXLZWbH1p1
qc6cjogcZ9YU/OMzYAtwJSDIB34J3NU9Mr+tSR7lWvHiBb0ZuJMibpaWuElYRObX
Y4SWjDwRk7Ib0Zi9j+0mjPN9arP3JCjXv8/o459y0boGlTbcmo3mGpCq6CJbS7M/
sE+SOJHio5JihD53bGdR5SJta0Zye5rRJw66nsNybjMDC+N62G5PHj1H0YOJQtZx
yECaGQB1yRwZ+w6pRAs+t8cI1ktmaWKsOj1GN5wU5FOyFK9zCp7rXNn1k8Jbi922
miFw4D5iCY2sq6s3Oh4D8IEw+X/hulJlWZHCm0Yt5iflae73wUuup83L91fYCRRR
K1lh/pG/7btMyXx9Li2bmNVYfSxUTQslePbrh1X4WyeCn0j4ML0TqJ66MbE8gC2C
v/luikBFKix+ffj5ucAEzLW1xHLetPy01EGwyFITlicjYdNv3uN1ih8py8PTt8Dj
KwUPJqnLRlt+LTEuPpEIw8r2tufkEhK1b/Faskt2fWfCPMjrEmQXcEeXPstUACsa
BRey6vKWCCWgJDUbyDtN727quZkG4WrTCZAqgGl7o6mIJ3u2OelAnVJVgaJDM1Mc
RwFBAYrpfB5iTt9lkOrKMG2sXe0j1kbfT6rxDXBOERM4hpSkfZYQN0giCwe73DFH
xMW3s+KC6NeeNubKG6MtcznJ36w6gvRNDtRx4IsG46WSctKUatC4O+uAI0RwPpB5
dy2W0TbCyN6GN832/C/6gQ7QVf7+D/cv//bc+PhQwC4/iXoWFxhG6GIVZxfzuRE3
EFWyQLydU5uUwB5+eKMC/x4S/XiDZSANdY4aO5Q7c18smArjHB1VGxykmqt/keJu
yNaLsGsMxY9N205WCaKqK+jnHlgvVwma7EnhuNcEiJ+VJyIfuaV+GBH+3i/Je+04
/tqZyjAd8IsbdRcnfDb6GUfQiLUpJUxSOun5TbdO4sq+HTu1mkbDknZ8I8VjP1TC
ZaymPQfGoPVWVwrKR3GWUz0GlkRpntIZi6A4NQ6v+XAOUV1EOdUdSZ7UO2LwVYlK
eZTzbAAg9pb7qhuJsgos0D6BvqiwUu+ZClrXdrM9WYcTDDjy8U0z96KpFlG1tu7E
HV/rKNhMZ/ES9VFWPVZDaFthJ1nkwMripVG27S4vj8NbnKQzOPXgI7xBniOpjFk4
aJHhofPOvIVsbO/pZ17c1e67MDj6mVLBzktrBV7DJ9mHb+KKAFhFyesOrZVgaBiP
8oTfx3C1Vz8y47O9eY/z8/Xpra0tshi9WVOgU/IaZeBMQw02VrbsytM3n7W0rZyV
/7VzSpsg4JWMvLGcxEi2XNgMqDJKGM95tA51JLJw6arvif11Lfp44SIFysmZb87A
rp6yknrWnxbqO6o/fxvzZIBCzCo55h6V6Kg2uZLkzm2h2I38UPuCkjwee3q8gjhD
gvo6LKarkgvERDnnOpm3rVdyNhnx0crDUuNFBIRZDE/5Y/k790SafpnTZjLqWVxP
wJB7EDPE2mezhHBR+nHLv+lGeP6O/y908b5rPuUkCphbuuIvmU1xKkXthCGxBhnm
1hmi6WMbfCZusy8WMi7o+xCcN4EL/q7Shzvvp/0GVn60Ty4XYpCUydL9mVPCJe00
76m691rFdfud02zHm5r3QM8DlMuObyow6S+bA4OX7khPQTRXV9OT3KZtVAVAs3Xl
uk9mnh3UvQIaeIa8BdGIwjBfdyfNlZRfiZ+G7HUxw4xkap4cMaS+/3CJHmFlc8DK
Lt+3t6gHz3roLy14ngpdIEmJN457iWQRxWSQo58zGTUwVWs2n834bxZumHBr3Xdn
bgd5XM99YhDpCOWjStCsnyPGz7UBZOhQXBr5nifMntuaNCSH4e+qjyw7fpLpbVXk
VYu+cNJzNSVcI608+y8XmixP8JX5YE54JTJLT0WwQCVYILcZ4V3N7ChGUZ32brXD
ofIn1LganEMXJezyz3572TrhIE+iR2X3p3IJmzna1XaRVISZVUdLkpzONH1VyOpw
4BIx8UzJeAB9cAURoNFnKDxVWFkIu/nhlJlWCAYjJr/q4we7bTwFC6Q+ug/vcRCv
4VAjUGBBkCdxP1ZiVvN0xSA+Cl11AbHUuTceANQUM4FgmE7+CEa8wYE80OBnPgJq
LMr3iXh7aX8kERniLbUiiioTAHs5whgFogceEiX98cqbYNoEnopCS4McR/R0RFJO
wQsI7CMTE4dBllCu3X6eXuh0eZ6E/MzbCQNZJZlYdrBsR96cGopQw3hEOq7UJ+1J
vmobKNJY3oqNhMluayW0usG6567o5CD1C4CXG+jzPdcoRXOO053IUWFBV5gyaQyO
Wi7SIOzkM0ZRcuNo10MbJgp6VsldtKUO2n2CJyAyEWQOrOgjmQmkUwuyp7k/eXu4
jDb/O9Sqij7EL0Uwo5kPrjjA/YHF+Ag4krXriUcnlz0hOYdSYt6F2okqhDTnlwrJ
zf//LdhdOMA9lf9WRZTHoezRJIdgFRujPCAcF0cHJ1LG/zLHrJpB360SOUEq7YI/
5NJh5KQJe0Y19GL2UFgHZfhiJKUz3lC4Bo7XNr4Vz4VA20NliKiokamOIIE9g198
mttGdy8sx7jumNW31gMZKjk0i3IZJtVdgNpnVvnh0EedDMhKsr7EBW8CASvAlgYq
OhtKQc5hclg6w43zZAx6cPd2lXWgN96Xha4dLwacxDtt6co+aVtoNNqaV2U7hkAR
vdx0v2Ceb6jW5/JcwKo2M0kC3NLpqGTM+qcoLHXtx408P5yg2Ux32T8BuHoCLIe7
rwz1PXcOghm90Sv9N93HlLaKkK5IT/CNeDZlisriznz8ze3ICthOKi6Wwbn4fW4o
qTjatQO465UtBI89UM6bnSx4ZHi1OdRW2gfIh8fq4slONtQ4JHDj+xO27u2aGotG
rlnVS5G6V9YC753p3Db4kpc01Aoc7eDYWyyVI+NJFn1+BVkqgQttvUwmd3c/kamO
qyxrsR8g2qXt/tfIbbc9yEaCWmh79FegIHgAj01a5BTTD3fQANgTZTL2fizQ4C/U
cNWt06KLovGDzHYPjhc+iePAtnj2BIBcFZ42r0da5WtOdd4h33p+inZLhyR8FZQZ
K9Qz4axyITga/mfQqzfczmCk1utooioXLHA+UPyXNBTCmfKrrA2WMYQXF1GjqJxz
/763XdD/gcMWNeTM5skcrdq1E85z9lzG2SrjNUESp66LN74eoArtijYB/QBVzSdN
+ig22ZbKrIwKpGOBW1w95SoIBcgfd8SWbsiwO1p1SyRrljda4PBhJOuwNCnzZR7B
vUV/p9CjzReOcgoTAlQUMBYCNS4FWKsWfsghP3eXSclqJ9lIJfpu1pDzUcva6ZGV
057mzzRnexaSqzrBmhAFra+dDX2sCmx9/kBOoasxt14QBWbKx3noySD3cAUUHDi0
wSOcWZlSMEG7zjyNC5EUWXOmGbB8YDUIdYGh0ZdfmWKp/BHW8ujLMQQdQB31qotj
TxxQW28l5eYmZzU9zkFSxsogQAc+jO/uTvX8uM3hQQxSTOQxZ3NlY/D4oFfdeIcB
uu18Nh9thqdelmuRvgv7dGTNEIRL2a2u2uIZRNYhXHZLwk+CiGhMbgBgqvhfyAUV
LHdp2mwUVJfXCPCgJ4tiPOXcccRSJWcZURUzne/0JC+RIahBQu2P5/W+/P/Rnvvz
zIdzs3yEQU9y9oXc69xAkI7Is/AA8vWP0a0JfeWfY2xYQgdoVJT/vVdqRypW4eLw
8lqB7oosN+E41PYgo1ww+dwCmvIJcR/lIF8ef+U3xytAbNmvayYdFMbwUXdSAxxr
Hx8g9LgtX+1xxPCJJgXl0u2QfIIruxVv2mFPLcg5znM/mV2XeDfHQujNk+H0L0XJ
sSB8w8aV4ys39aJZ2OuFTirNRxDsikFyucCedG2kEiWc3m3GgeBSQfQklrfr7TJy
Vby4cS3xTqopkHKnc/JGvU/p/zn7BDUKPFuxfMXYnntNgbTv0UsTs46SYYJ8DJDn
SpY8IjlZPMbsXwOo91Pm38NzLpNJfnAZLhbCz0DDZPzNk71Z/f7Q9Ue8SVQlkgFB
X2B43jQFzxGguSxxEiu1KB8+ZXyI08GvD3wPL4Me5/uyWm4uV/zSuESqSKS5WyMB
u17fA6eu0NVJx+NuZpigKmw8xdOdInvXyXoR5JecoAfJ/rrojmd41Z599R8ZgDOw
eqMbOprweTWQJc61ts/HX5p+wvpAjqq2r50zjuBeq1wPqgw7VpX5/q3KsWHVfeMT
aSmN7QWfLE3VkgHYZc3sHd4ik2b/1NpbvxqIOeoNtFpU01a5WloKteLB4fCKH7Dl
c2uDmkTczCtw2JTshKBdHG/d/Kf8n19/OQzJkGTpD2c7Fl2v8wnW4v25k3wEP3yx
pCvAH13vVC8R0thn04Ll3Ufqv4COgqcc2F1l6nwwhIPIXcyEZx8lCnSG/Nh8HaZ0
9wkoLqDCJDZ7irYS7zL3Coa/jdGBqd8V+hXFQx5leXqvsea9nSFkxA0K33pabgTZ
SnfhFnoWGLTkClKjqi0VO85VXPBxV5I7+lOWp6U9ah9RhX+o7mCFR9qp6ie8C5mH
E4NV4AI9Pi63hnCWSatA8RoQfYgqXZ+hEJzdema5WBk8knimFg53/1OTulS8HW+s
hsTFoO+IAayrMVz6on7SkNVXwai6SJhkFXwBUFS9gwH5yukunMU6scjPA7SMOf+M
YORjxJ/ZM5GdjAjUvtFk8zwAkwSUCQwN5meIbTGBwU4BvnOaBEvAw21Dw9zebxLW
8tO1pdjdw8tTd6G3afg5YAPcvMqKmUKi6VSmdZBB1pYHytqAII9lmhdhZT8heSDI
kmeqOETEuttbKhv1IY0nwsyBAbFfaNr8oTPzpA778rahJitilfgcqmAKP7+7rPjw
6nCkEkDqFWmFrdEsx7/ON8Q7WyA+DK26ISjP8bGKDzkZMLciDqC2ljGjRzsxaL03
vswvYra8TNkBog3NBIchvVyYq+pEK9+52yO8J4kMBIgGMMp+26ZTHGzZTBFsxaAC
mvzEthSAPUz1RhNbwEF5A/bH8144GH61ht2T0yEevLSdrRDLQRUvoQk64e9xOTJn
Za1imT1Q2Frpxb6aes1LEaFY6CtXgqKb8HA67kIjxxBtYzg/R719fi+CXom02OZ6
H6uG6VwgwYf1zFZbZgdmixpBoSeGXNQryybcAxJsrsKa7cBzATGe3gc1Xmn8+DfS
OM8etwKE3rLtTKCkszCmVe1Ju21A4hMkPlHVJZHEwCrxBbuLkXHRFDdJY9A8Ggyk
sE+EllBF50Jr0+yoVqVEK1S1VGfTYco5KJ4bAi+3brc3XAuzrEoT71w2wOFscbZ9
RnusW3Qt1AtanpCdZN5OrBz9CScvVdR7ZhAxS9heTT+k8Y57uBMJvoOb47oi3/mA
BUF+JnSSFBwvFq43ItsnBP4VfinQsgdSbIfTqv6KYeWtx5uBIQiLhvhBzYHKKfdK
qoLaq1YVTGtdH3xoUy2anFhhOL3lH5vc2ZPzxdOYRydtCS7aRyqLzIYLQC+FGgYh
XWnwv25PCx9g6RzM2DDqaPufjElvnmoZefxzsgkqDRa6T7HL4aAl/rUhmxF9L3xP
HxNWJ0V0fjH5u5dffdXVw11yXpSyWRg4oilBeHnsMcRlKwoXTWOBXDob9pyUGsFR
0XAVNW03YCdJYDYytvef+vhp5KTuYYYeZT/+/d1kGQfVI4v9GrlZsbO8hZEXkeIE
w45bNncI+vFQ4x2XR1tjPZdrjNf05SF4afoGB8pHrLYrVg8D698lCobjuXyKUchU
qgTC+kVPtggwml5K+RXrI45ey9e0gsE0hjsJKW/DaHqysXIMwUYLsmVWkHX7uMH5
urC91mPEs2GCzudDfAkEcnplevmWbAfBFk+y5FXhZwiHVimXGhrLyclRj/sqzWFQ
mVaRaSXCwXeQ3ztEPWJ2cS9nM8coOj5uXdc3UaeiSLhsnbW7UOzsgvt8DDCAswxc
M7O4vY98hEEnK51F1b+Zwaa4ztqCqx4xlX7mfrVrwwe69zmu28dtxAmWCKq8WP7z
lbaDCui4zzX8BlXGXgOIzco5NCPW8vKZ2XsYmAHXDY0e6oxujU7BkGM6rhw6tY8n
YbI1smDFQb6Aef7yg8Uw4TkHRoosq7AnjlPj/cZVSLkrFsmdd5Yl3QRd3MwVIebC
uq1H4MgCmoes4NRC1YaNVFjXLnfxPMN+XjK65rB+7s0Fh+18TKIs82Sou7DNUWEf
MHn1YFfoFwy+38nTEo4sE6Dw67gyetp5g9LZAaD/QUHCD4SA8YiaWTGTuPBKJ/Tw
6LqNzjARPQdcy5VgWugMhZaymdKKOzQiAvJ08Spk57nUtoOodqffZDACI9avTOlt
tcDpyXbEj254bJfcxOcjXoYnVRK5/rhQUlFPGP8agwWX0vYQy4xRF2ddewZyQvDV
a7HJkveHjODhw3nhxfmH6h/ly9M7IGFpmdzmWXuJWkVu+M0XPC4UUmQTXvocuB5W
PC1R3WPwvve70CCeb7zJ2pN45qld/3u0qfQFCEXhyOdXJnrG/a7Jpy9m7K6sI1ul
6+ZneqiL3FwzQ1out7ky4tgdt79RozANMcwhVpy66dYcsFAU1xXZF6M0Gyx8diNu
d0Zg/4JwBGTmE7fFFl3das7s66e2dRsFmSy8nwfhhLO4W+Aj8c4KVS6sf/3hiJt7
fnfJbJMpT6chJvnFanTtP7awakqSfUw7laSF4P1Eo5O/+bEk5xSp0KbsC7U+KRbN
o8gkkARzdMLVWLtPh4auMpcG1ck1hIu2JaCLjqPLP9OcCUVZPMXlWRTAtHyk9xbJ
CcTe8hU/eyQ9v1cbM5FzOf4QWcR7i2AdbYbzRu+CMvdTExWv74cFJ6xe9h5tcvBs
e5rtxx0Txx3SMbSMRA2pyznbRU4zfmLRfWS8HCyz0PAKluMK+rcZJCKa0FBr2UvW
+8TT1OYfnRLdyvoMgjDClsUDvdDyD7rQ+To7POlJhoPn7Sf2VyaEpXgO4JsnriCX
8YFTTcUoh7mUIAcrfrFYSLSMhwGlRfhHvzbMzXCvUi8EPjYM2RJ0Qy1PwEenJt0h
z6B++pmAO9u+Pllurb9ouD3UqOfbE27j2QhiMvun9flFBp9FGqDn77cX7vbwW3L/
rm3GzBSCehvbDeU42deSXhSXbEPq9Vr7ROFLZvM77kcI6wGvFwGgaZocTO+4vcLM
dp0ikyv4iemp5TJvGi+7G6Qbky+qhVd4cfohBr64r4vfklVqsS2UE+NbOws2W42V
ha2KL8sxmKAdHDVB4+8f6lFqMlEAzBdTPA3a2FhT83HS2cHR1ZmW4gez4rBYRqru
kvy0lq4E19IoXECmH6a6jkUES9u2zr6QZP9pn3iyUL8E2tobNrbytl68Em/CjYPp
035YaljLxSB6Rm6uswItyMGuW9QRugYI9EKGOEkP2csmqq7ob9+1EhqouXL+8UqH
KB7qUKCpgQTTya4PbD5jgj56h20uVd6pubxWDVIboyYbtbuqZtpeRjKnYgepRCja
fpoHkLe99cVv5dirBJ0xWyHK+zX7Xb55hwK4v/bt8HUQQ6sKI3TpPC+y4Y1aWj0t
5OdHw1EmGSTJ2O1sKznSl5ibBYWPEetypuoxE1m5b1WtmdLaXO3iWa9aDtjSMcQw
Obpe809jln1MNfb0z8SLOtlppxfHpWzNUcgNsS0la9h2gyEVKdzJYxLAJ93LLPrG
hqDGBRGHd3Kmw/vn88DxcjFoY/NjZSM2vc52+Cd7NFzjFfEUkNiRTPMSF4nhMUwC
M5GQXUwCbKxI66aK7BkD5Dh4zht7r141mzA7700q4tI49pebHEs9nTW2fsU2jQhq
pil/NSxTXbti+LFWaarWiE3NK0tFRq/BlKkiePLXOYO0DEbI2tQPK3/TN1xXqIzB
GHX25ARp4hx/fxe1QRDi2hw48ZvpZ0Rh2q75SOUugQgVWYcgLeMPbchKlNf3Seq1
JZqqubV+8KV1E9i44w90PCw7BSxrgZ5WHYBxwJBcgd/pnHEeoGkAxiYLjnpLWGpB
KcoZKG2hcEKgJMudRq2sQkugJpLnDk8QL7mKoeg2Gj/5l8M1jR3+AdyKg4r2z9Ce
Soc/xyEAZ9ggTMcZGbZglvE6zhiNAnIZ1+xN7qf3hWG7PFU1e6qNE2yecM4kAlCY
6R8AU/hj/3pkpOKBTlAAJIIvj01JYBKp0Qvotvqh6S69x/106iQgASemvBMa86s/
jjmAhUQnZtbl5GSHTCZlgebPC6FRA2b3nKkN5fDv1erIA6nV2+GRMX9Tv0wpDRi5
upXB4CC8No01aSVMpGCAzU4jd97PzfSxjkk8Ah9m7oaetLzr9JKBblAk4EzSP0dh
yFBpsno2GZKSJtNy8kNDyOObMT39vqm0O1x27xtF6pZGtKEQw5UjBgnFFKL5hDTh
YTOYLDpLtENg/je3m9ILRodV2f/GuXA9CIwgtqk5RHXh4ebMl+f/HzNgUKMk0K3j
rbaROOAdZ83U06lepIS2kXB4mGvyw8yWFL7BWwoaMyt7foPYaa7hfchxfh9k7fZg
S7O3JDkXAbbjGP5/0chuxNZTY9mIbBneXDeITTl/Fk/FyccuwwR6QBGvCZQzd+mK
DlF3+fhaoJNTDXhmI9tCkJVRKJTlIRH0XZR1aTogjGOzSzbd8+IzCZLLgYKeEpS2
CaPWLyRv0U8p+xzTKLAYCVxHjYKVWNSLuCQXtGgxPbd/vmB+wNWbXaZ5M56adutq
HLLoKkhctHvhGgjue5f6gyH7yXO8u5EwZ5Jgdfn9FdJ1uJoUuj7cU4S6GJW1U1o1
rhD0YbI0KxMW0WJp1/tuiYYjuAcqebUEzBjxRvq2ZC4RRLcvr6Sibdki/hxn1jFv
+vQD/H5AevdCkOWAjPAWQzYlF0hnRfLuT6UW2POYop35jesomOxnToGzMpflay1P
L9dxKWRwzIv2LH4W8lH9N1l5NZzNVLW2nvmeV2i0ogkthOKKq0sXNlvm/ommeDdM
+z1sjqg0kdhY6Gh9tx8Kx0+CMuJyqSbkyeyfvmXCBk/9NqgyV7n458XzmxrY8LEW
45HoZVyWYzDE/HVby6zwIQ/MpNZZTp36Ls9a9FPEebeSTy7bvLjcpM7UBHC7hlHF
zG7sEKyYLyRmCWEJ9qEzm7aamTQz+/H1o2IDEyKZu+dlHDJ4h/fAMug20jBy8T8z
ZSh7gzQeyCyy+erQhj0JI0NSpwnPDepYIO/gOW6/YIaSTTRsrxM2TCTJfMz6flcj
nELTNgCm7Ido28HqcNZGEmTklePG29NkJ1gw/qi2Vd1lbtOoElYFXzL14InmzecV
4Ae/rBSKWEEoy/YiZAKkPaVCmTGhDCokgOpV5CxA+itGs6i/t7Ss3HluCiw23Ty1
7g9BsjyjwL5vlTNq6RY3pFLD/ZM11/0cAaZceiUxZ2ZGX983PBcnX3LCI5XZ4MM6
9OHUpGrlBP/0MuB4K9m95I4TwLoKf4/2I0aMUp4ADd+DRcZgu7f0Itohnj+/OIZn
26tRJYisXETCcMJ0oS3GRPVz2LYB7qPJfepB09JaBzlKh1r5PGfCF+skmkYqmsx8
xrIqAVbbg0bK8aPXMi7fRRnt2LgXio6Su+fQ53S83fNmd8I1gsmvoISS5qV1R/Nx
51iS4AOnG98qBZt3BdMdfqpU+UREqvCYNaw/6Gj+DbTE5e+Bwwgrrh+xJm8vN92H
oTZkWZc8daefR1q/ArKGPUYMK84cL4RLnADybvZOXbB37D28DFcckQLGxxL76C9/
G7vTF5CG6CUgNL/HVmn2CvwXdBX5SfjV+QviA6vwwOOp6/zqhgF5z9nrhoR4ULlM
LuFUpmkQsjzozE4D1N5rJpLQFVS/Nlv7e7qPlt/Uqnnt6CgfdHb06E1p636CgR76
qfjVEILNg9wWxE/oeIMQMnAlzGlYRtP6PPIPxSXGfXVHibYq/KgR9NV5r0yXWA4r
3wO+97U+my0vRSRlfJHekXJqBHjvv9CE26yuP04XJZ3LL81ZrLKPK7W8JaRpyl5a
FOelBLShATFosuC4i/H6dfSWUWnAVqTqeWqHCBk/NJdvtLD3yjDLyk7HMwaUp+lE
dum3JNJTt1a/EtMh9sBA+/+D+Ma2jlD5iXj0Orv5HNm9FstGtkyrhl41DVMQia0H
fEfkadi/CMDewXDR7It8GCffTg4CEd/TMroGjVtcl+mMcQ4pY2YLAIO0lrWsGm4O
JpBUjRpVu4YMGTvkxj0TSj0euQ/GASgi8nLfhl7QmFBgBCXiT6aROVUi5UJUVdQu
Tb9B1oHYofiPALzEp/7z2d54Ac6jIpH2UEYBRtyibxkpjkJ8QLagxr/yOkwi4X+p
bWL+GnP9Nt/9G92IzoQmT7Ewd3/+M1uwEPvUyaOxGlbw4Mx0eq2n9AG4ChHRURlV
Zd0x7EOZjgN9YG0ISjL7tJPNWKh6kA+WvPyMClGDXyBQylqBWrfNQG4hONAfnuST
KKDubK/Ez3Ndwvp9CWBBDq48+gOvCuVjywg7Xf67UA5GL+I/nTRAOQs3qgUB2M8l
a4D8nZtO58eB39v0eVKC08dQVNhdg2ek2OcgL2WcMq67wg/08GNieQXzUjiWzAQx
HIs1kJukF4MGFRiyMJKGWnZ1psKo2D3A1kqADt70SlDhesQrmZXeFomDw1T5rSYY
TTftYHOMAAMtzgB4YEx/zAOV519Yv0dVQMjPc6MHxzXhXjcu9zPJPfOlbA9muORP
obK+b+j4vh665Eqkvpubus9ERwpHwz7QAUcbFq2y545md/KNPLtbZSJtTf/Hei/J
T52hYQcsMgYeToMl4FjW6tfmT/FtOivu6Jzsz57ghuLwr2EmistVMyUpuEk2P4Kc
dlDM1jgSewdIaC93QQS2dBOXcTPo+05JAs/Vr6A05/TodM2EyNtluGAgvizLxzsx
KH+orPDUblZPDpVHkBygLAtYSNvrtBp5jivi9L6M004kc6foH52h0g9a0Bz6FURp
XLgKg/Lvs6yFvLGw1ysCzLxrmvuYxAZyrEzxL6tG2uniXncTqyHPX0wlFYWRGkgq
UQ7Nv/4D0loINjJo/wikL/NL74I9V7r0DFUgGUeZrbq9Pt4aU9YQRCgxcckmA8De
R8sfGjNmDq2l+jJS2gCA4UTPfcHiRj9d4KsRyPBba0vH6r25xby4t7lxy0ZrO6ic
mgxzKG//HcBFeIuyI5BAm5q9b4GQkeXAHAXuumGaN76l/OTD02q4OMEmYrlyw6wO
sjiSzFLqY0bLGMd/TvjBpeanqSMPZTDjgpGQK10ulcrV/J6g1DMInxi/8//B8gn3
+LnT7shJ1xavH/nBBCC9oUXkxhM9pGuHVr/CMVAwXbOYoRX6mCUX7TrEgRgNXGpG
KKn0PedzZkfYF3RscuuUHrAw+XmYIIeT1ivg2m/ewYXiLb2D/+t2GMVjGlNznLGQ
um+tCus2UTKo/BSqBdrjAbBI01cSiaq+L/0NpOhqRScgxcLTo7arfwCDrhIX4VfI
49nWJT+VQVin1hasdkOBY7tzR3g72Xti8T4jjQ+uXjiREp8DMQb6sr8WVSzx/BAO
mOVvxRg2zL+qRV3MglqZUABJQx1RM74R5/fZc4Ga6HcRTMlF267iQVoRJMooXXQf
WM3wGV+Y1p90PUJYXDj3gNt7vgpUL+J0OWCS+yjF3uZV/OMj2tfAgn4CTZ4YuDP6
Onk0VUey8RlQvDBk5iaP7fMQ/iis+PI1iHGCc/G1X/+cnMxbrpRO4tNzO3J4gOE1
t5Z6wTVkff3YUDPSBn9uWYiQKVLMSg8oIHkIqTVe0rSWb7utgy5BH6TNcxvt0AfO
1tI58C1fsLy1OsAK8G/2jyv/vY9uKVMmlskT3CDcpJowLo9+An99sUkKSPV79rMR
EWFLJzp/+43ZQc4XMS1VwHCP25Jr3OICebecgDEeu4oXbVeGZQTPq4jMaikqCkcd
9tQEDHfS/QkkJZ+e9m7CviUGZ4NEJ1i6grIpwFIXUkCX354+4kAUqwVLG4t5AkMs
wz9R23UYH561POD23ORpLtYa/Xkr85/3Wh3iTljB05itxaFVlzcQlmqtWLIStxSn
xHvwXMODyoxLhvRLN7qfdanqQq2n5E7pt6qN7TtvHMpN3B3XAkOC/qmiRORGSFUR
HdFDpxEvjFQmTTgBnVV0Pk2rzWJZ0xKkz5UXN6nd84OXdasw67l+vV628HXfwjRi
+kwmEGEtwC0f6/AzPrHVK7x3cgeliozBgmjdrP4wi3wSoI5LFsW8+EPh6hXpOya/
fown/IuIZBbc+RNFF6blyRaG4/mO+Nqr5U26kFKMDIjvJfiZMYSTxDDs/TZMG42i
JyLvJUI5S8ryOMDG1qrbRnSHS4Otg1tUyGZiLWNH1vKNp0ypPk9S0IMD+ERbCqnA
zHHfdU1grP/IwaeluD0/7vDhmMcNs67gizZXyFG120oeKIGnrN0vgaMTJn1cttU4
mGKK8i9b/ZOYyIGcRHTDxuD4Tu6iozCFIpbP/5X+SFDzKM7dJ3vsrFM0Kj8O08Oz
FYie01STZQeBRJH3ZRvdRAA8k85dpOoByhi+U03qkyNV47c51WpusvQ8tysVL6zZ
jim5jk33LnCBQTfeG96OKCS1cM32LtqAr+au5WrcYYqzjzHv13oCwIeMsIxvNc0t
ZU5cc/CessxFJUqAruu2CdaWht0+CZFj7tVKE0FhUZdH3aJrc/u37aV4HIgJS0Ud
1T5zpgMPIZg+6z43X6r+zxjfMfjylXNBHDQaBQ0qRxjyGFElxZo8719RCb6JBGl8
KgnnR59W0MUoCP0MZOfi0llYyT03zzisNXHrXd7Cx2NyUB/1SCG+tzCEMW9LYs+d
fSdPanyLO1x6Xf85RnGoX1chWBwG3JF4Wc2dY3DGNMUH6HnnRayL10e3B0V1EqrX
XSrf2/GcRxonzN2Zg2Pc2iZ5VO0fmphmcU3I9FSR+SaAmTxW31BXBrvgE6AIJxLG
ji7a9FyMaEaOy6ZOIxrU/4dGblHJYlIOcf/JdR04h/YH/poXDWEO4/YbmMp6H/ea
DEzAeCYx78jA5v1P/PYbsxXRCUKgxW4Dak7HVtPfwrwy/i8fh3KiufDfHTQyP57/
ux5yXIfCU+Xc89ZysDwepse2nRXUBHyrAQrQa8ONtRB5++wAnkiIZOZnIkM67UvK
vha2peeYXfWAzfAimea1k57OIQ3OY+NWZEgBCwe7/LnJQ2A00TU2Zjagz95mQFky
BgfxsMirTU1K2339fAFlMRWJRCAQ2MTzKKcMQAlAsCR5rB3gFJ9GuSGPKLQ20hy9
P9M+sE1FgmWI96FuLjUyVGjYChBMnovLK/An0cQG9ecYoGjwtC29to94HP5t9ZnF
P9PK2RillY9s7xCfuwXKYDchrWCiBqnrn6/6+QH+krNr8KeW3cJ7HQQVkuU0W1Lx
DssCzWnb3zbkYPeJUBdl+Iy1gcIWZPDJiPqFG04Dszg9+ch5YdH2ZkMWl4CYJ7yi
+Fcu5jicy6v9Ph/bIAFu9FrgkkVGU4Bs/ncGMaUwBikguCc37s9+pL/uOr94SabK
Xg2ug0GJsg7lTmID+V3fQJMTTm7Q5ahflI2IE1ABUbPfQ5nYd5ti2WQzUxaTffUf
n9OcX5U631mVrh5brAXkmW0P53VE0FVZ0uBenshJzlCVc591CU3PpOCzLXOTOAou
VXtxt4Y4GCwiGbAQ5JJRtmGLSZWHThNJj8M0zNUJsgdPdGM5kqoaZDBJGnA3Y2cB
V1dRRrVPZ3eXfvCqQcSJOnz6JH10psolscVOEYwczpF7B5PmdOQCLW0SGAQ3/JAr
igdyOinMY86y9QasratpOrG6JQyhS0AfjqBo2UZnZlzAglLsUVkwRpAqtA+lvJ7a
ewtiE85gZ/HVE7Hyrj3iuS+JAQUtdq4swy4V4/wj16A0ENjAOXJV334+74LdlRmC
zDx92GrOOEYhOWfox1kQxabCLVxlzqUaxNVg+iuKS6M7bMYU6yHwf7a40gHmrglG
I2pWymf5O7SffowBwC/zZHzDKWlM2vxw9G6i+tZ5y3c6nDtWpFVLstMoOx9YSqZr
ctPhbJGmvLqVcP2tp43skhlusmSfyFdXY0muw0vVCCFzSE481Z9FlCfDzOz5wUG9
pJAO4nZYcOpVeDm0YVeZvE2ixFNP3WEIjHxh9QzVmG+1OICfDu1dawwV+qWuRtyp
MdxQGN5Mea+3Kxj3N4BqqLukD6A8jQNhpiWy8UVgwpT45dD5S1eJOg5nYw+afddC
MLCRkMieXtTcdCW/U8hTqEpTGbpIpkJK91WyLbjyWT8+P8PFWW+NyUrN2FZwBj6z
CK18p3UKYHwsBR98WSwnebDJ+iA+RVvGR8COqLbp4nIRK0p8khfwQtu1uc2OZsh5
u6tcEfts34aczamnKOSa1gB7b+JTTgOEwmKSmwY6nuctfSmcFBRB51DR6aTlb8+0
+fuZcbBMETZ2BFCYHb9ALtC6S/JqyseWCg2+hb+2Qc+dP2ZbCy+82T3iwg4S9z1R
WG98HfbqtoIwMi23tryRybGW7Emz8oC+68icjoylpP2c9q/tNWWcpTHi9Fi1SqEC
pwCT0HdassFv/DgESYDx5e1JHDID6bKuV29tLIaGHKhziUBnTJ42a6a+QvKR0rmC
0E1DE3r9y44M1zvpI3nLXXSxJJC3+cySfvN1quWPjj1L+O9zYuLYZvRDaKV+WKlN
n3UdLKOWJIuTYgOIPxQdOktWOqp8Ulk0WClPQwOy1uXbsvv+VMH5Oi9vTd7P8HS/
dQ+3ZVHHmwq6scbipZPSNtlAOUm1siy+LNFzSXGK8Bo7DZpGk3jN9Jd5YNb5w6wH
+6UdLYeq+6ii9crDB1JJFGEvSc1WIlZlkhJ7ccYB0yRZYx2rWxj73fuRewMus3w6
BsGq/QNaMWY3nNgAVerCdWD4xpnv+hFOUpmc40F9H20twDLFTUVeqw/ec2/3K66P
Vd+Y1o7him7YCXAyTm0mp5pAIP+vUQ4MFcINjkn3sirkdyXeE3S3DiDca/kgiXyo
xb38nWoV6fs/ig+b0aLrRHgw1Xc2UgxXf7X2AcINI/vDDIj/2/6ELGFOChPUq2ZW
QxKBG7CoMFD6gLBIG0PrGDVKUeAy9lrPZ65MIpdOCHfIMA/EvIi2O/QhviR0zZsH
GTE1eAB+48kkYKaLXyOO4FR6mNW77w9oQRpQtbyJrfWu9bZvnFIVgmnGWXpLWwwL
NFM9X0LiVMXYr5/EaOwUvxRKIsyZ1NoEh1yvg42/8lc9rejG0KwfqTifZYNPLJN/
XY/gl00dqJIQvezy5s3mdK/xo3dmtIeEZA5vOd+daDLoaKxKUza4fvaxkDxpGrRA
jTicIzmJQsJ06OTXv6QdIwsiWR8eG393tBgqo4SvlCpl/VHRkQvoihveW4NLTESm
bkeXSRiMtN2lYl5k9FFBRfnEey5gjtopWdktGupRyPKts90rCnc1DwmkAXYttG89
QE/o1OxoGArcSB2YZUpQj93fO+cdVnqI3JN5LbvPIaJNTT/jfeQJ0soTIT4nyo/z
j3ilTY31g6Cz+HW3OdXYgAiMQTAgybMIcg8uCVa+5Pf8TXsB/jNIeU6nyAC7honU
ryeE0b76TqTbB20wVqhmTD8Axgq3YBuBzcCOsVDzosrIK/60r5qmD1QSSA0baIQ1
US4ZrEnUNOp/MQjELSlIjb24fY+7ujZ5y69QZHbX0jRlKaXRjK1Z7xMH0vRw3CDq
bifrXDgl/nCYKeLLBo0peu2uYxHkbuZiWDnZPOQ/AVuzsRE1dqm9IIzptuduMlqa
lZgHDqjaFhXO285PPOzYKK68BLzklbsjLLkfHpYztNOWaAiAGi07du90S6aMX5hs
8/rlqCZb8p6jIQdsZeNhlyK6Ogh8coBFlEVSoftmTG4g58L7rkfdxYL/OodYGXCw
T4pkqwiV0CZ2CeeI1cSMjX3CCwkKsJfoZrFtnE2lBHOOivk+tzj7zsKtmU1FnWbO
8vbKws+tr/SelFkfBer3bqgQFKXKmVLaskeY0zKYLpaGeh5bkIG9+YuvPN4yRsoN
1QSSrKPXa4rmLJlNNbfO0seK41szHBG0IBLuFSQjJztncBDKlwPC6XUekLIsUiY9
k7K8RVY4U2DdrC6fIJbdAVMfwZrYIpkSDo43TPoguBWcpFDWzBUc8wCy09o2g+3Z
GL2aUoWGAl9MuVpkx0hpu/FLKUa5FwRxQ1DiAdQvA/q6rb2x1owOkOl00i9blbJY
TaDZRljOQgdp16vPM2pfDFIRTs3cP0LX6LDAcWBbsC6RqGOcReQrx+ZSNJr3wylY
/yJK3EARPHtTyoxpjCb6xDCCLP+klji9H87zwgG+WgT7h9KJwEfbqwTtzIYeRP72
FhxdUP7LptEqD7JHZd3SZ2CcTDAehd01b3Tzp48aXxOfn++yzegDgIkV5NRiFR3x
4PytqkVeDe33EFdhbEVLuNTFOPI1grX8IVflfH6hzNp9Q0jgC5qPkJviE8thD750
7lyA9wtDFtOjqvOEZ8srrLTN8WkcQDN2T7r7jnzXySpAUBXGUIqCNDkaaRLHOWfN
O5/LQ6M+5aaMcf1l8Xb5ZSqtOWg/RZjCQCwSZt2D+BAv8AfghtES+8xWPchQmLxU
ryrk2g9FPkWOEY00ZGTJLoUMkN7pMPlK45OwkGjG23RBDHDF0C31eeAnJjTx9hmj
KKWkr3h2+nugyd6aKvJVVzBBbol+X8Rz0D/FjbAYhNB6aECdmrpNVWBw+cvztV+2
2SVK4A+oxtan605tLKcK7L8qVuRpfv3BpHwsKV/jI7NyV0p7x/+vgXp/lV4YUxUE
zDegy6ewDe9LgYVGhFpP9UficQqbCUfx5X8W0tgwiDXDW4hO+ZFTCAxOyQHbQqx9
NUunoKpa9B15eVB5BzhAREslv9U7N/tpnXwuRP5+lFCe4pTE+y4Q0d2MX/9wgYES
Re1XEJSQYDfoQsiw/cugz6S/koHqGxoXMWAtXx8qzXW3O6ttHMqu/xNZnomwJhyH
mYA8Qz/eHay2JxRLW9lyHVEWPVw0j3Gz2YofbMSnMN0QTJFS/Mu6Swh8EKC7L4aY
n33JRZWQeYRkcP+F3XldXZz+snPhriGUwHkftoHk3kH5/j48f9EF28Qiy5omd6Zl
8CthFAR0ma4E0ESOSi/CuNxLHo4mvpwMnuUisaz0SVhP24H6+C0oHw4Zaoty+zCk
5RP3YV174p/l1E+okMvynTjntvG0qRlmkuQZpLJuCq0HiPmhxccVzBvvLk/nmijD
u11R9pDlTD2u+iylBcPJoPJKVtiLydFow+MxveUHJeMrjb3U7Md5kJwAtrX1m5gh
g02yL1Ps2jOEgDXj+7HjL+h0vHjQOtMtpb2Fo0P2D/r6ktI0sxCigyg3tuZmBvRd
heNGvv1zMvnxrrlc26FYWLyj+oU/ml526Cc61IUSZgL2gPB9ejfq5IWFfjD2OWHb
p/70DbPZUhaENjbrlq6zNUUCnNbND2RBNO4auBAI8PPXc8m+Qhr8qUQVKNFJEF1+
FTUa7C17hhZxnWOJ0loYrZXdjI9RxbgtLx+cajw0Zp4J9ADlUWNWfhjbVZ41SAE2
g9quV4E+2gYK7XTFCMS4BDToetrJbD/AOn0nmrMl99QzOVQvpc45l4gVhZ7vvWbb
Pszpx0HbzN4K3/Ij12RXJSsoAzcZD2MseMU+wRmwDxlDUBWLmzBNXzKf9fX9Html
LZo9ZylvRKgntKznSG9/W2wyKloPsNxIvKU6HoxZ47Xq4bQGwtm/zu+pdw4lV9z2
MOlHm+lHs7NmSHM3Xw8JqYQnBw0viFTuKw9su8CMPM0R52MyHSspnJvvxN0mP4K6
0a9kwplblion2V5WBnIZhJOQXlm6BSkivBk20FohO/95MhZk36I7xejlezElX6UM
6SQxvhiADt1PVYh1xwNJuVe5/0CR0hF5PC/RIyYwSkCpa01a7ttzGn+ApnOXIGEk
wUzdHSTyzO+bFGmmIPRaSPLTNZpXxlp1ehxdjTA3d+lgG9xPUXHqf5b/s+vnQm4F
kPyF5e2nv3QPPUuc3MLtcZ3xJ1qAjOb4Zn8ItTM0z0go43wFwBqaeFPvLscIY9ET
ZVrDe8sGgw2f6X1tbLSHZ8MKzeZbxuIZIad2DZIKcWeZfVbRKqw/G9pvZ6VAX18y
01VPxr/R9u7WGQZ/ETs9c31NYi7y5Co9G2Q9AWWx/t71NQDK6JpZp5LFNMUQ21BR
2pDT/U4BdRaqn3FLKoRUOCcx9GqzhuNN61Qxq7Q929RdrdFPgEUhrxoqmnlOIVoN
9Pq1ONgaQDzon3oJvtnhPE7IdpfMmUxjIdduOEK8Y5PAHusT7Mbh1f6G9yBkaRIT
SCpwR5XMWhP8pnmKlsO3gAGAb69YyV7REu/QKfUkFDgR5umFK568SSYKvYtRIt9X
9Zjnh6aZedRIPSanSBB/u1nHo1qOYEPXgO8OziMZ7o0CufuShaHj2Rfvfn3CDvOA
WVq5Z5h+8i5oIJe9n1IJLKpcxiMo0MV7Ne8an9YcCv4hRF/vs7UATDSuV2K2hGoP
6c6w7VvsppR3yLntIi5nTKNc1qrlEehD9KNwug/ue+RC4ISIku3vCVkIZFfPf94h
KFGGqWyZHUkGiaYqvr0SExXNXbfelpgIDAS3HhzLnXZbYlKctKAfupR9UFWiYHzU
37U1h8MuCjbmULS+dfDlBZu4fK2sFarvciaMIZUbWF5f54OcKm6+A13/qnulF4xB
Dis3jv70kVv+Rp7V4IYMmHwIaaF/41ofgeK0BKSOFBru9wQK3j930bBpPwHoR6hS
hc2Vxxfp3CpGmLSN1+908mRhHUVTt67C35jj4JGH6cq4fdn3RucW5O5eJUXfvDmr
3RyO/DaixiJ2wA5f4ADsXqDFEgKqb4q04hJ8tJSS8pON5QmAPcli1DAmAKU0Bttc
ZZGBqp4/ZkbR0FLYE5xE9oUtaY2oDI90N15xhm4kbjID5neTwDOKSVwYIjI4BnYH
r0fdH3w06lKSClFhqr+iOADEkxrNR6jR5zDYiVUK3ZKTBblcsjlR2VtwE3bSWOQ1
RsE4MGWsYYSAjikQX/IjfRg5GggFar404BUjQ0shNdJxoTHYWTn7eZ0t87C7JP/Y
k3AcYuwlHn/e6S7PsoeBBsK1MQPGWQoV6BM8/wpzdUajlSZxbwVjf3e0dRtudF73
FNVhp/t70CMEQpeQWXl7OoWgb4l/iJ4wHc/7vfJH0LVFmekUIZxMecfMHYGVhVFE
TsIHN2n7rkrHYhteoz0ntfa4s54d/5l2KqDiuSvrBsm9ZgAscx2/ihjfnirEJ4+L
14pRUy0iXMOTgLAC0X9yvBVnuKOpj3jdk+BYdS7/F73a3rNR68XBhw4x+JGwt4JW
9tBwqUaDDXG/XhuF4LysSwfPMbtO5PbQK5j8B4gct7sQzs+XnQbosYkgmgS5TW3a
TPcobsdH/7nWT+KKhLOKS0mKvhPjS6tAIz0J4ujgSpOprBNTer+16A2VI07H2/xn
JgHu3rst7rITAptF4Va41u/TmMI8VX23+TWux7GhLcnhDGokBRAVWsPEeTXmunPH
4TaB+RZbLi1rFJkeR0GyzkO0SQvtRYR6QGPmiDSyMNonfTvFQp8OyBCS01Jkk8ql
alzaZbe6DgiaykXSByxWrVCu6JKIP8zX++oK49DfjLRRMxmJZEW9WK0n7cGjVleg
KUYAxPGxh4+3G4C/KDB9gaJ4VMRZVzbKhdaYgryr4L5lwi6M05dXeXbDiJ2uOvRQ
V7DYcqkj+yKyeyphFh4kQ8KeJdtje41jA/nct8nZHYkK9/uVV2WgFHCs13Q0pbJk
Ew/9pCxH0YzoCvpOz0o8o+0HXDFpCzJP98lq2vNWtp8xRvmj0XO/7zNOCOnF+R6l
oZOCCGfY4JtQcBkccgMOCYETk8UanLhJvv2TeWkQV9AzmNAEnG1Uf69Pqp1gyrTT
k6LyFve883rBpmavR90afpYaNaMbScIiL7nwLsvP1Gy4DGa5HLxv+YVS+Zb9098F
oyqdUr6MMWZmW9w343pAgowvtsXUFFx8yBtuc9oi3sc69xz4nKHEJdG9wpNocoJp
mWJhFK9/DC7jk3Qqmitl6+z4eHpYxuCizHOApB6kZOMLlRtb1/3li7wpfBzzBwmZ
UhA0OqnnN9ScsInI+kaFuzkfXEpRpnbqE9TxPQpXJEYCg23vSILX+WqHtszZSHIV
sRYkcrQk9RkIt5yyNYTdZDX+124WCU/P9gxbLSeTVRHItaHOnKz+bhTIZNkfuNRU
aD4sO6es+ogV69oCvJTb5gYUZaJPaq8I01EJz2gTXSoxeNH1cpDDgNOFPYryP26L
ea4DqQO1MGl+lcqvt+Z0g+9wbMss4srkozbFVayL5bDX10kCo5kkIE6wfzF+2EEQ
NK/w5xta5aYu4ihMYVa29AQy/j+ku0bQSZ37Zo8Ax8ieCMidZCLdFjO/R4Xh+Rg+
foys+0wQYRJOu0W89O/YGaFfnoZDlJilly+2mPKrVMcE1xU6mNSQh5jEmii3pUD9
1B+MWbk3j4yqrLUHD3nLQy/Z1Iu+kTbqc3WnoXr997866G1NcKWRf4J6K+4RRfb4
e5HgzDJXGVkUHtmHS60YAENXu1knED71kFzXrvoskebmvEqhteDU65hPE/+Lbp0N
MB+4QHlk+SjSXiKODHH5vk4y8uKjvfWFXw9Ipb3bbIpo+kAcq/WkrdIcE9Q/IBj2
CG70GXFntJd5bs/RdHdjmVEd4ohO5t6qxzC6k8rEM2OgRh3tfuwKYM4BYvYNxlx3
SZAMnDLeyf/EIL1WhT1VYAZOCLB6qtytNNxySD+sXtn0C3SB2nEBH6V0ums6qhBQ
ki14o/rke6Z4WTE0xOmZr/TKsjQA/uQ2umg8EddJZyF4RUwQ4uqmsGJRERQ0ylEj
/xB+8SmSaoWHB9z5utTCvIRMx1ZJBViCfui96aYJ3XIvzInyI7cR08HU2bUMOTr6
nfRfS0z6APAJvciJeiBEr3k3Y4jc5eynXE7bVp15Lml0OotBAludj5AKVQt95IbJ
YkPHKjQXVgUZofyNtkJRANAr+GmFghp5IKs3SCMjLfDrPJ/1OrxUcx4RrQ1RJCVN
JWEq0Ay+mueAu/7oRn6rTLfBiipcWbDEWujF3XlOhKvs3V2v+IbEW8VxquZKUPiw
huCqOCK/Fr5Qqbwg0genCv0zhvKu4mfKklOKDmlrmywfNc3MgjQfY2j25BkUCZHL
6RXLXObRCCRdIJSe4Vk4SvpcY6v6UjbC0CAdKXr4qB0xl9sxMlA9M0A5GGv56sJ5
2LwcDpixFEYNCQyQzh+tqHOtQ63lnDegQ55lX/tTh67w/ag49Gypyt1V7XX/mknJ
7zimEs2dLQ2vNUb+M04vXwKW3tlgirK6k4uxISROSH5oAN/0H6P6frUcLohxXsiu
BvTBhXFZ6zp6wIQLbPp1BEibhCE22n9aMz0/342oXsRhY9Je5Dh3KDtzrtCua/0h
arVye5itJj5SUvJGbeQSitoHXV0JRkbkKRYh2pdt6ro11Ke0WYy65tgDvVXtk7ju
0mDO4TJ5w+jtDZG28QiWoiXt6d8I5yUcdGyCz6xxRWlXq1pU7bFvPhHsNwRCSzKr
UZ7/jdikwf35bF8HAFNr5eDM3mhUCr7tTac+eIOi4r7p/gOqzvU4Wlwj26LCHdTu
DE5SBx53IqEWxtmQOxOjbR8ons9Y6NtWDWT78jepeEMRbeivUH3Da2RcB0IV5OKv
PKotpx/yp4iyPI+LKXiBN3afeHWOr/wGRgrggZaugOhGFMQ73A1fCnReEKXTMom2
ihtEC5iCMvVGmxQt5GIazUOKPvC1KASqWClRFQIUnpqItOZWDH40raUQzyy+VMDP
vsLWEM+fiRH3iSwj1C7CoyRs/Y0ZdmOq1r0c3MDoeBp1EJVzfxYyR7kgirHZgksy
tASCEBY+YTiqGBKW+goL2fi50ugdRnlba4UJdxabBSWUWTOzgLWNGRTCTr2x+TUm
m5KqgF3FPfONh39GVMlSK5k7tRPK9t3jG1KhFTuHMaLxkq+PvHRcBwZJC9RyBa3V
5oaDIk5UALf9SQQ1hWwyZ8F7y5eNBOuMjfNo5IUloXbFXc1hS2uJY4lohWSjnm06
ArRmdK1jLtRXZQZzN9PyMnalX7f7m7r9ND4g5sJuO1bkAHfPIk49iQHBzPHMUfgf
evTPAdr8eEulNY+THO5iOeQIpnoiutdkp9VbMXf0zCismCQTUUgjF7H+zkP5MuPg
WTYjixs2EDLflSdXLFwa68hYnZvb3K51+sogYgiDD8oriWtk5Hv1BvYuETmdAg+I
w/TFoevEQx4TbO8KbVRPEn8WmQ6fVx2hReAQ6TgbGwqQvoXyGpLwtewothYp/CZ/
Tt5+LvQyf9RDox8YqfjZ1FwAyrSdEvTXW11dW+4dyyeGpWa4giWvYTYb5nqKqM4r
OfpfEuktYOvJdVohTOL3LLjBtMz6b4VVtabsmf/HtPCLHJGulmuXOuMTn4FrLVrN
ETpLecqvmrQvJYOfLZ8uDH2vxnw7nL3m4eOl2iZ/UkFWLLE8SA79kusais59JfLi
81BYuCjKr4AtQRnSMzpOLEnYEbBCNrzDcNhPF5tpmjCTQu0eSipqIOpBGAFKfiZB
E43JrPAkxdNDu6NbIb2wKLldSaBACIMe/+Qpczt00LurCcq1BKjcfGFy1Lx4G0Oc
67MyQa4aooiMwFg5HEflQrJU48jPpE+MH7QSsRZvKUdD/c5yxpkrnKo8t953jvja
eScAIFY8v3g8ZCCrG1ulLlWMeIuw1OGXDBWve6Hiqk4JCaoBdV613DjGE41Uv/ev
xhd4+zLpR0judg4iIq+ecTYgdl0Qs8RiSv9hMEbAq5RJnNvbsYKJjtd8eXSyaVML
Si/3RJ6RxwbEsmh4fjSYhW4KFN6tGZHtCn8QLLivMi7y/+Mbor0IwNwac/I6tGYY
qEJsiPn1vbSJ2vVPYV4shb084AMC1MiAmx+02limSypn6d2PtRK0TTven9dtuNfX
4763BKZ7GEdULtFnmNyFX+9jiRNXSQsqqbUkYtdevRaqBKlTIrvnrzFgmdj9s+pY
wJS9EvrA/ahzn2eEc4iUfyyelluqA4/Q5MCMD5OlMmT7Efo18o5X8YwDmFHIr27M
tckewyQyXTQPJ188ngXePiIbwfzOzZSUWFYjZwCTOa0p6hv0qac5WuPLzdhYMjFh
HmXEFSri0fl4psFHtfIpiRlU9sK9MNf6x+kqAGMO/ydV6t5aolbLrpyveyL6b+OH
mmiy9LdBOjnK9+HsfSrncOBQJlNCRkfRaRpWfqmTMgdtAGk+JTNyfH9iQKQ+k3UD
rTWnr8tsKeo92M+vonoFzzfyXQlfJQEcHQafF32jpj2e4Y4ogDxQ6o35BxcNb4De
DdERTK0OjUapdyrXWoCoP+MHcwQflY1PGtUCtSHBZZdXer4EHNs1ONrW4mt3M1YR
jBzh3QY5kyIvSp16K3NrgQswaBiY4Fici7bxkIddqyi56xPuv2JgJraQHGm75Re5
J/l8HDFz+PunjWyoqSbuRtn9IhFov8obNfbz4DNxfWpxlus2GWuRaWt3HKv+tSyL
cEJG0mi1HKki3akurdATtqkx/2PL0u/N0Qb7b1jS1BLsmsQ00WCNrJK/1zV+nHQn
Yn1OPLxhDu9JcFkew/goAhn0jeykFFaQBBgoRAKRva9CJiY5abZhpDEiauByRlg3
qhohyaweCbjOHdVmFEonV24BxBC7D8WknEYth68qVCdae499EF3MsZrPyBP3/mUW
sDqSvLOYO6ICzhccOhbyuVbPmb/kbfV7x61C4gT3rtaGQiOfIAPC0AxGp8nbwjdc
GvS/IxeRMYEkgK8PRz05fAi4/vho/OUY2OgSOIM1fcY3564arRzFNUbjEBGio/GH
I0nQeEXGcir31SArcgvJP52+SgTJLgv8le64G01jBMV1KQMHVq2sw0YWOe20Us43
D4RQ9E1rIHGFiB4tymwgBt++xwYOrWP8YB8NGN3zY0A1Xo3hvpFZBAzTL5qR2/Hf
PYx846h5e9JM5wC3xT1IScw12/EJzZKBRkn9LdRPW22NQ8KHy3lsRAZFAmUDkj2U
5dVladUeX7z+I8iURzrk1UUUWhz3G+jvE07nAtWqSTHC1O2Jv2VjAxx9YGRCkAv3
EPRvmrBh6o9uyJ7fT3s3K7xFRg+oQJFUt7NqMSCdQqwGJiwy4XyhoeC6HYQIVAOl
4NboDjF/iNv8M1DUO8HKLz3Yxn+Mc+jNeAV3C9E/5oiv0/90PKLLErYTTdUSMR+d
e0vHdt6C8ENXnoBhCToipP1M8TY979B4vFtflnFEv0dZ9F+LEl8/dT35nE3SM6gQ
sDxU1fZ9s/TNvLZtVW5xupqWsb7cQRmfla+/HgPUWBiuaA5Jy93YTbsMG3ZMEth7
ev4a6JFIY0BWdFh0bnmgj0XpFEBq45qAUzOypdp+h+tOop9lfloWIYpe5vjZeUbV
96dN/Q4PrCQPNCjzgB8bTBJQTdU7PA9dNHXEaNjVbIuWRkPZDLoT/i0S6srtWWUr
kcUl5Hb6tcs4O4ZZofrJaHmXxg+n0oUuf9szavw9TlHHfHlfXvtDb4GOQv8U6Jxa
fTcKDwibvYUObeoy0utHEOo8umVgwAgbhE+v4kpLKhhodAO39fHM25r730fMpGiK
uZcZ5fm3GA0k5iuq0jx5SlpD3y/xzuMh1g0e1VED5ZtVezc9+nbRWJBfozTTPoqb
1N+ieZFE6WBxzR6v9oTPLpOQSdOQzvFrCKAOm8ZImdSp7AIGnURuVlJWeIZsSX0V
Fx9h1pyrcSiL4D5I+l2lPRWphvGrf8ZSEGIkYz7MAHbzuupksBpVbGNpCafg+X4M
jhO6RbD8aW5jidBtJFQBTTn3TAIG1uEswM+5CvcTkohKL34UW9dEIsibxFP+GkXG
NZq7jPS/Oivd5K0L+5R/UAZAD3fpVhh62O1akO1YdF2Wz+pi8m0ione7IHYz08fq
I+0nt2NjJEwuPjXb4U4DbYTevuVXBVJP+iHPenHPl4cnyVYebJG/O/R8LXtAnVtG
2wP2wAG3tvXnubgkdSWwLoud2oh/9dkBiO+qLw13rl9cfwTbb+yKI0ov1maH59Ad
fUIboCpjLKNINUegy4B6jkFyC8GqcxoEMqWuT9Q4auAQ1Z5XO2gytmLcTtzerL0K
oFkJtcK3QxXvioc9YdxntrBHCyn3iDRwv1TJiUaXJd8AEv/29/ExY23Gs4GDenvX
T36JllfTGnbhndgi5/7NhEHFC0lJZEY31qTMVPUsrsTtmISwRQbiLEFCWhyWlAnX
4smyzIdryF6YrC8xqp7MJjkV/zLef/AlXULn2jezWU/hYOoJnd1PPyDBtxaJpUd4
4799a5sMLzS+eTeHP2thE4sP/MybB9AVr6jCSjW5UMhrYh+MxRnYQ3IaotlW9dhh
Gu0r3NOM6p5YELSWDt8czoPH/BTjkn92BHERf6Z7xNrO9xbo9dqMiQ8nqIcayn94
WgjzachDJsBPQlrF8uYcnaAYRcSYRkDXK3NZl0CnZjfJq0xphs2Li4UHPz5MwFUJ
TsGk1f8JANnq5UNego1JGCRYhAr9u+Ku2Q19ysoPrPPv0TPwaTMDHeeQWUhjZ5Ur
aDRvRHpfnEW0ivnPygp04mDi3bmiR1Xya1k6W4FJqUTsqoz9KgTF/EAc2cMMVNlZ
eJlFP/nIn5G8ZIAkcpwpO02BRdIsoLkuuBNdAwfKlWgktiOJTCrHYr/QigIxg2Th
9/+7/c9mAUUgh12NCe7uKJPyLoI3re2EIZXdE1foIVNG1Sl/NHxRa6Ck7R5BuGBF
lh8dyfMP8lAfjeQ525qF5gU7/ocnSHE/QjV6PgND4IhUD6vujyj9V+Yj56I6Pvfo
FDPUXl2UzrUwb2IdxciLOFAM/ZC92Dd7Wf3OOviZDp4YaBHX1KYJV88A5322lxs3
WHSwxbKVxDpXeG53CDkT2rHPiBL+K6tJu9cDN9ktAsPKieLygLPprv6y7bTgx0M1
ewLzwYCf1lv4iCmjHjAa0RrOldpanUHCzHrC8pG7ARQ9Fs5AEAhnXidWwvFgasXq
CDdrW905q3JBCCc36ZUq99KV8zpWclvNw1i2b2t13qNlHSqcb7wIf6k05XQtkOPm
lsngoW/l9+CV5gZARwYMdedvath9tIhg7Al/2qvRmaF+EEJM3SBJCaBiWIwJpvKA
BPIUIvZl6ssBzVK++n58ALZde/yDOCtYlmAKe1cgLHu5lGblXQS8AjLdRtMwQKve
SWo2xN2vmzGPUhoj7r5xpreJCpFipaJcnb6DDoW3Wk741rN6gxEc4586dy6ILYPk
Aj0+FYln73XfqL9m0phVhC6nG1kap66t6rILhH6eH2gtvtAeNo0CEqsEjMwNZIQP
7xwo04koO6456K6b3erIrc+sczdoSFJWKzMTukmd/hgNR7QjeVgnJaCKYR370bAW
lGU5pd3tq99KL/IczA+/7suyitY8GZWqN/S4+fe5AFU86xiudthUBRBsongsJJpz
8Lk4RLSBz0xeJ6HbaoNikO62keqAHkV4fDCIuo44gTD93Duf8FM829zwM+3elfZu
9uMt9XDaocN2R80S8PWCJbegbo+dpvzP4/OU/KoHvYtIvV0rzBvU/GDNxEG6v5Bk
XMIqowCXgeDtpApsrbTxyXiWo4CLydKWG4HT37GfsZ5yNL08qooTijkDGHbvR7JT
B3k+C7QmdQK1ztcmkwY1wwhYjGdg7FdJfTihkfWBSPreP2k1QSHaXvtFAaqfU6xw
kmTjre2/d6za3KeAau4FmnJ93mgCeWCg5zedzppgJ/P75wPs5bfymfaTblJQOamX
gfhn1m15KBSEvPAsaS0ihVwcAXtPixAOBFvzHoJtCdmua5pQrfpqWyOYSDvXaJSs
S8evIMBgu/tuYXT8x7J39bkJdyTdoojrwFfT9Knx/gt+qNMXagwtW08Ub9ufgaCm
rtFAOW5BKZJuD+NrkYOd+N/P3EU9WawG5C1ZitK4122Yd0xFw6GbaXsLqtRvCkD6
PMCbfPm7xWlAmpvHe/fouY/Tb1OrWZPJLIz/C1mNdiQBkWZYcp8yYtnJbGvhrfpT
g/oxsSz/4MPECzW3p1cSGd1B4/BNk0CtWKn69lyJUz9vE5NjHnONNu1N4kc1bHVx
ASCH2uw6WYiBTfpc/T2OjRcGnxrgeadmAqZ7Sp2FlgnPmvqLcqbpg84a6PjkyZXu
QduBZ2l2AOMKNVUbbKTIdoFQ7APZnVajI6urott4SFY10F5Ocf3dQsiKu5ZqMswp
WdTVu9QlK5kOhiZvDoq66uH4Z4w51LYKza0DYb3zY/63el/oQFJgo6z8MCjiiAQd
hBbHbJxqZEvL5wA1HDg1c8UmC5e4zaXcPo4vx9k3c3UPYegQuBwfq/seKnT/3xTJ
x/NmuunuiLMKKFZG0+bngA0HNe1MnB2i9BPgw0DUWcvM290F7NbxeJjrIs0qH60X
ybZiMDy2rJZHAve1RDn3DPJYuhaVskvfRs9nLofpYso4ndz/qdlRXNO1P1znHl0J
FzYCn/5t1lHGbgeJy07DiKy+a2jnb0qEj18JbTykIBkaHrkl7kFPLkrVZ6976EoI
0MFSIaHXE7tmkc6hM68cAfI5vy9JJ+85evau+V0Uy7pqBOZpi1dgWzg5YAwUFBN7
fDPlkKIWvJcYTfqHcg0B5PM6/ELCH8nairwTy47lr/f++SDpTrkSbkHom0btftxx
gOZN/29iwAEyLYTQP5nF8rUNJb33HoQxkIdrLEkpC7hXu377y0zyn1yxBGp1mjZN
XjnUc//UAFXr0PwXn9YIPR8xQCQK0N7JDB+WPdhFWs1/Q4PinmNXYQVvBcqQQk2y
c7PrQKbmvGJ/8aFmi3XAtZxne346wERBC8N9NiP6GYYHa86vEBeOKQGA9h9zsOwA
TMWpNFFqAY1sfXR03mhyhLLgAyE6XiQK5i1x0aS3CXJIRqD0RNtRT35lVhgMhw02
8O78qcgyPl7xIn7EYnGK/DQrjnCYzG6S8yeMLM3DUKh2j2sZ4YV0uuE3HhxSG3Ti
T8yHXuXmeZHOhAmfunuDp4sOLwPeK4FJebhaSo3g+obfpS0jk4A881GTPFM/TxRx
CCUqWYDpwaXf41pHvliAOq7ydcmJMNkYZ3pjggqAyZR+8tUZyn8k5nrtPhezqLzb
dE6ZQwDdw0mFCtxzUgwNc1gDMTN6eA2/kdNcnuKNVA51ld66Uu+YnxqMK1z4R1Wa
K8gb7ZSDZKYod9RDKzFWGwaOQyD7yzfIc54S+XDfFRM3HZOqUZVV0hcR0EV268E0
/dkHm56LfxXKnBQxy/4ZGi1G8XOR6y3LcSYENHSvHh7JX1X981P2e4EhhIAPY7AQ
1xVpmYRRvYSbP5Y0dSj6xvPuJHjrxU2gT1Q+qhEJ1qGofLj/mrH3KfZb1NAvuRZJ
v3drQ5/ObBECCJl6O6UgvUoBxjajDrXxG45r2NxN2KK+80fpBJ4rXks8RXy7oiHk
qtwd/5n6SJggnkOcgOG2kpPQoDtHsOfXXUoJ6KmcexkFGUrTinv1jpqP5BGcHUjS
rZfcQblhehzei2XpHSHdT3K7nRDF6OjIxd8Ual2BPbWs91VyYG1XW+34pS8tOdny
4YHBdoHrLRwq1OpwiD4+kIrtECY3yOK7vcmijZFse1+EMG8Qh5B0vFpajdGudCfa
24kbug5V4B62NKgrqKHHBw56m1uvBM61oqU8XlzQgKqOsMT5FPosSbLKASAAC/fa
+JZY658cd6OA8mv31FQ2Za6km+NBY4OOk7qvE4BtyjJMtRO34CJ+AfGssfPWKVu5
IbOiiqPY9EVBG24tlvcOFdXcvd3rN/1HRr/BzP9bH8WLxiuY5heIRvyoh563zv0P
sJ066WT6vqNfoXvnqL/uflXzLYcvi7kBhAmO/0HQImYOVMMhAZTQOd3qq6PF6FOr
5od2Q1ewlpPFCMSh/YZVUslDv2CCKFfipuVCEqswEaFWVmmEmFIUCCK81U0kYpqF
cRqAio8xr2EC1GNxHE+jQppW5qnm5A433Njc8T/Tr8lf27AZfNl8rpdWXxWwH5JU
Jm9i0xVcIOQKtqpHw6Nl85rdg4dLf8ERFglFrp2Spkm/3Yg4WKorJD9exi+DpfLA
zxrWZ/wgZ78NoRVlcW6PYN6FZnwdlEeGkWL7TfrbplNMRMhWhQOHJwt4ACrdkAuS
e5C44Sqd0M+UP75PMMoB1N1EyM1Wf7T7B1AH5FkIqYkGRayIidZDqBidcwJL1NKs
9kIw1voaPhHBJJHmpiafobFoUITxi+pe765vMke5fJscI7YO9MPDRS5JPJdc6L6O
pT/GWLoFNIRNNmFDKx8ZCFSSFD9WEh2k7ZlIA4CA5ajvoYUfmUqgy6u2AKyXDX96
NnPpPeby6rYgxURjdR9Ne1Wi0GXpY6VaGOYLKGYLmzq1mVDFMKGCsT84EZ+r1xUR
IAKfgSbtVRiCwkSKtl40Z6Zl+efm+M9NWFAYTB9YKzvFnBRTigVHeWo42PIX3Mlv
d8VZaS+OoRb0VhzvXQLbAVPrr9+UlM/P92MgZ2LoDxAwxkakwcf7J+BZiZh/yGjm
TnedDoGeEUM0K1tH42jsuaL0QcvjEsBMI+Jm5/KyNP+9gXvtsxy2s15MCYGCexW4
gRUgfYKz/QAWENJ/LyjcrxrnJz7RVSmcmYPQesfhYGYo7jYQE9L4J/gZU/4tV/ea
SvwUYjqDaPYDKlefyZQKldnYO0jpUIZyT5uRbPS1Kz/0RRlmdI+MR+8FTiBp8Xq5
rdzn5uq/uQC5MtV9OyelUafhuNQYjxi40nABNJsEKplIjDQqjvnPzpAmsV7vPTkp
qJdCc8xke8q7UyVgAnry5f3MNeH8cG10iEvy55WJSh83WFc4+jld2a6apEAJQnFK
RB6ZKReE+SHvNfxrNf5aUv7QLRpBGKrCQ8MkJczokI9BU+k7SzD/4frvpTVf5w5+
zR+IGTWj64vITl500S3+wd5wUkzA0ILFYBIYbVPM/eAZRaqTT4DIZKcsPBJNDlK6
cDp+cD6wOt8htZ3Cf4RD6BMWxk/6LiXcKAKN/w6o2RnFfvAebrIlR/OeXNJBkyEJ
CmAxJpf2uBymcZrhDjANan/6IGbM2DvhUs+Dzbt3d9RVy6W9A4hJxahZl0Q43+zN
NMRUNtd5fCNv8azx5mTeZQkLuvhj5z8v+5i+pOlZJkLUtRD171L5xEPJVTxB9Axx
SGhpoNqvz6dGo/IdJds3vwet2y0QbOTUvfwe+aDQ9UFMTlbhLuKC20a1eoitbwH3
fdxjOGGtPrg6vNuBew2cwcXATJTVDM0u05SeEtbcx82NsZbwL7rbq/QQmGI5VZZ3
27JorkqydlFoGXOzTtLhGXjZ25bWbVP/acdRExdKSZhg9VU/m/foCLML+ja79iUC
nmxyWOE8YM0XjsTqER+48mnOSuSDtwTULwo5zS9riUeZs5Zsl0n9cmzA+i3juety
3M4BYnf+dEsqEIOs/fLHLrrWenzpvzrZUvBdGw4y20n9Abp3C7L/VpHnmE/+PY4t
u5nHXqcSfvOJeG0JRaRs14knxG8aqfAQLY/tf6LsX017QAzlPcVqHEUS3BYuIQUM
y7rp5ZhdU88aIDaWspEV0oPL/pu8WmDYU23FJXWYjrQZfygLz/EB2Dd+DBx6XmQX
7/M7R6Wm6jhZreWwtHnT9/c4qO6NFLRVcNhlsnz++ysVN+W9ITfci9RoNuXTs6IK
KPoZDyJPB1Zb7z178RC0birL0mOn7IFHGTL14qRA6MdnhJGiwCll24TqNoa9bw3V
Ligsr5gpfA/Ob0oTBlZwJmPi1i4YcoKavzfTvsNJzBzBJkhp752ely55hK33k5pL
ylzj3SrcCZXyq2hu0RT6myYNoj3yrmJahudkWa47WbT4EwYoHLeTDDk1MAVHOb9C
l288koKTlehcB/q4yuY04PkfJkKwZOY0JgclMIo39WMxkNIJA1emzlJ59xjHuAVH
JzUBKdYxbUVNFEsEo7fARPy+Ty6sULMGqvnJ1Obv+6woIfNCpTlD4taWL0wP7tEH
SCmxpXfpFym3pOsx9BCOe+LqjbFtn2JCv9bVKZs3HFcePHdhbVWc6TFpC0VXk5Ia
ZD0jsgR9m/oLf2bYon7hWTKNEof49sfcPjLVSsX0nGsJrmZSa1JpbgeLBdkqlnxv
E/H2jfPAVyl07sw2A9t7yiAE6SHl5aNPyLrdqTSB4X31wbwR8OSAHFxcqz4glait
wSNGNP4DDoLK8nm1doGMcthbh9DDqxXYWcAWZD4otdWm3h+A7pKbACff/ADxyJg8
ebuuxnqT5f8u9sVl0nyrmGMbvgi2zxxWjqTOXznwtcQjtFchMnx+Entv+Tts5yf6
y4SbcDsYJwW+yGpgKwnwb+UlZ9wauoTU52pc0DnmZwgyFlDMoPTsXV53zl+mu2Uw
v/wazdX6HOmUtTo33iccHWhJhm24L1t1522uLj53JFjyOCrqG+iHuJsXchLFucP6
Q2qnlB4zBHzdPhM9Xc4291iNhkpGRgOiCuk3UglCxCa9bEpMx2jarjABmlKgbDxR
EJMXYB3gWOhbILd+yd/3CKgIQCZaKMj5VN5BkCjAJKyvnO+YSRh0OP/4B/nJ42gW
5Obg/RoKVIrNgZ2p/QAjUxzCFsU23jeRkjPpK1Z2v2ipmbHZYP7pgD+aK+UX9eq8
FozTORhZ2whE1G+r6WfBhRBF0SPoLD3q8lRn5A9+Uln4aMFVmPMfR7qoItf+YH3u
RdwHXCkNWv7Pzy7jfrmS88CJceOUxapt9aysOUW0wr5gEjnTszqccah3Yw5XD3UK
ygj6AMJdJSQU2ddXSf087jHYvYDlm5A0PtArac7+BsvGv6qxoqVclOpDGp+adiec
QLSMeHhUzT8dy7jNJmgvcb0yf0WOlEJuwZdujTncf1Lv/7cQoCrTwpUhdidvwPEa
26xqfv6FknJ1WmurHFwgJffSYE+5+USrG5cipTlpeWC833FD7RyiPu/cGOOlhDQm
3xSlD1bpH2712vY0nBu/IGPfx1DQr1yMlWBxX4kGCfn6nzDVrPgtlCAOzBNH1aLa
sJqGYhfMctgaU0/0ryssxdyTNBm1UAk23t5+jaPRj6IMCvuK3omtrxjWE20Oa0y8
lhaJOa2MTiYoezkvdbqusFLJk21uRI2+fM5UQeavT9hb4MDq0TMsicY1J6GDRYEm
T/oq0tHHtrcoQ1BSxCB9ddBaMZfpXl7XkqsNv6bAJ1ne7eyfKQvPWTwvYHhpbku1
f6I1Ji07sQXM81HdWNyCpsy3SogphLgU33kZNH7ddM3oP1jncvk/RKtNaX+hcn27
wlIMB4yaLZgGWoBbZo7ZbWjMVQuTX4S6JzJEdm6wJZ71j6QG2DOFnhWXEya12SiU
4NXML8lUgQJjPEcDYvy+Ec+MGw3CW3t1FPyX/sh59jL74/0MRVD59LPzwKcoCpNz
wTXbDwe8M4pvJEPjKqpBpk4ibW+l/boqyTjCvksjPTscdVjT+iSHmJuHBQtAvQtw
iHO1SLLj0ASH1XcdYExfgZwxjnzjv1MbOzYgfOX2KUAqEj+Hk5AqH7UhL60K/P+J
DwcyHnkn9ydSPU6prqEhK/vnQXnzO+FowE+eHaFoKgQ0VnfHtT80xcor8mV8nYSW
JZ81InuC4IQCS4hzrKTsSI/y12gLjo40TdFDR6gHDYvLyj0mEHnsGUJyW3kjt7QF
JQQ0igCHHPy81CvcHu6j5DdDRPTh7WF9xBxquI0UYEJEbHXgL0iOrxiwIFiHzqTe
LHya8xEBsScAufeL2nv+uK9o4r1DqmYPPmbELVW4QEzT7nbWcb9RixERIG2LozeG
MvsdPrHXmN2/xyU91CtaoC8CvmvMaRjXUZhmTuJqpVxg9JzJHxE+Vz4lqoKf2rqV
ykR8/QzaFX2U7zeM6M2svyXFtdHrAsaxlG7BazmX6M3U9+UN84UCtyrFRSwbuy74
XEppLDO5+1482RqvwSeIivDb/ak2ypfQDK4a55kEX9QsnmYCWHGC150ZTPD+t4G6
/wVFAQkjbbxmWHRk7n8jR1X0C2o1zX3pmlaVjR98X7UkSLqgSDq7FEfxQJkPVMym
+Z0r3s7IUn+/zm4sof4bB7kyuUoziKnFxzDAcbVsCfptZtXpfpfJ08pkw+QmLRFY
OX9L1Xskuy+Iyp2Qypk17kfTkNtxxqxQ21h+5xEXOj53ZOfzqUilExsLJLEuZsIf
ukoF/ZKR2kQqE7PNe+pFGpG2wzhT0HQy3ZO1trV85gR/j4aRI4NBkvTYU/4Hz+D4
P/VPbtekSzhZ6QG/KFn/F1IG1h2G0adt/t/WNf1d0uwBD4KuHsoACrRJhFqvK7HP
nLo4kUGDaXTSBa8fugFqLOs7mA2ih9cbGQ9TFEtzg0ElX5AAocWoFX6m7eXetSVO
srj3QzefHbuLtqSkkolYQzMu12C50BgcBzqR3hwELBjMwUmqF1rJlBQrg7UB7G62
Luo2XuS6n81A5n6FdRUEEI+ekQeu+K6EtJwqUqQByyw6A7uhWsWZhBRLYkb7Agm3
iv+loc5AbNIsru1faVWrsTUyUsODhgKl+PYDqFJFdXpjTi3oA8gVp/1jMEdUoIDm
Bfw+5VHEkh2lm4yasEXpHH+z7JUrVuq5DdWdON9qHj86kBH6GnSD7Hq3d02AhwOi
/NuX1t4D+dkJx2kSAuslCvnhT9GwR6FZuPxE/Yan4NuSyEvsVUO86NmypIBo5on+
JD3OzSCxEthBhzx7nWKZhL2qmHNCyJULsUObbIYOArcngxOTIVdzbNmHEO9dgv6Q
pNMQLqBHM9B97MxnDkYf6f+J/Drhr5ox7XOjzZp9JQf6guHaGx8PdmqWBIWqQVrz
tGT/kploZL05vB+D8kZetN9aU8Knlit7GCeO2styoGgZTJ19dxysI7o56jryWlp9
P1yNMCmY5BwYkCSrZtWpu7KAThtiVhVI4Qrh9wS5Nkmkld9LGwYwm8UDhnAVzaT9
cymGGBGrZcAG2Yp95iEIbTO2ZvWWmhwOlZkuPthokgRGCSjRKqvsd4gKdjuX4jbV
auIHOv5tDlytxRAP6Fla5jaoD31s8JYr1gAjBXLJBB0IJhSM6s9DvOVPUenQHbBi
aFfHVXVN9DaCprqnM8/+X5Wakd376WjfC3fp0XFzmUwmtOfBcTF0JPqG1bHnmuQR
0GuchF5vHtuK8qbOg6pc4V9Gvwlr5jEbqxX/ZsL/plSkm0oIlR49T2Kg31WW0mjB
NBj4xlDLib/Lz29PVA/8nhduf7hFoiU+1ofIlu8Q9YrWIXZ0whZYu/Osr/3D+TYY
phQzquvXhT/7yagHshOyC2Qx0GEQAQopVtFmsQr5L5ER5QFKnFvZ+ZCIIoKZJwIW
gfZhH+wnl/6J9gevIYTl4WneCi01hSaQOYBRoveAYE2a5RlDKjwMpe09535SsNLw
+JEz3lSGHk0RSndLkw8ZQSe/nVldMAhYjlrq154XEbj0TmB6qnF0f8IyLlGzIH+p
jQp0cU7osi3auwcTtWZWYn7C5mpSlV/L/Att0R8a5lZFAoZ1V9g96YBBM7grVHJz
/k7x+8uAMd/Iql6cuOIIEsplSZnVrnu0NAVouTmDp6p/8L0DAbQ1QtkL1B8lGlND
KkpP6kB/RVJQ0ORmXCQxDXhvJ1t/Xh7FEMRMQv5XV5z8AEhotl+bLh7ha6GMtGLk
9bNQD+VHdqZlcC70W+LvGCq3xHKYHa9swi6df1K/yA8gpypPTjmUzrVOpbXFzjto
LhAsl6yFybR6w1p9vcT+5/1W+dD2a4DkZ8m9i7ScbIEjiZw3QRl1Wv23sbYN2Zhu
4hxMZSr7hjGSioOAhLOxNIjN1T6iaVgvm19MY0J7TAtcjHSXextKlYUJ9znzhs53
4Nfq3C+SmyMnlT859ArYvsqL6FsR+zhAjCohAmgtUqMXM/BtL3EM97xRvwYCnmx0
fEFD643UNq8bRcaMcB0nNWGU3/TBlQNTMPFhHCIcjJd4koh6cPVjBh5lHaV4hx2z
pjlNwvVAStXtyMYcEHx+y5Cd+6O/pRk2PgYXTowuL4FDcTWITqVYP5BcxuKNKfUP
LuXnRWv9g02N6pDsj/h87S/pc+MYpvJ5EOxReKnC2wJsBgBn1QVaucYx+5qlLXX3
bPEpni3ickz0zc4S07zr176oWWzDf+n1bUZnsFtkaPoGV++okxH6kRF7LpAeRzG3
Qd562I2o9ZWAdnYTHdiDPYaaAO9Mrrp+KaJAnb8hcaSbnc1DOJ7iVsve6HZ6qRpo
u+ovPwXczYUWFUKoHUV+bMG2mZK+P/TzJSxAXZyTfboOQwljMH7cDcpmU7JbT2vJ
wJBAvJa213Xy0jpatv2gV5svwLeYHUO/pscbHfMp1AdvFyhoZqKdzorEqmiLoSAD
iEFqysa+dDqNCV2nxXBsrSQqS054OSxC/AU8jSCXCXfNvxuyW6YbBqda9VqWXf2d
ZmAFh0Htkq9wL6haH8Qf4F/1NlSJlgIXb4StaFj9eqTbQaCzLUDp3Hau4ZOWf4xJ
0KveFcCCtDbmctGVMRLerEjGRRcGMpgZhz6LlV3qXyk36rxYkpTxHvP612NZ1MSv
st9iZshWuELP482HoBq7QcA/Aoib8m+7D/Ff4QQxCMSbuNX15qk8c9GwrralPEhm
mTzTQdS6TcCsK44j59FJaCf03JnU+FNVvwMX2AsUHmlMGneUpYbRpl2adIWDWbW/
PBVmVA5PjJtfVb0kCHC9E+xGh5sxQOaFvviAggOzVc7CjHew7GIAyY0X85dspFe3
PKhzs0RqGtA+MqHm/TUYQypWv8DNqYl5VQVBPb4I1c4WIwpnc5D5PhRuPzl3lKMz
3wfC/v7mvK5eGc9Mrg70cKdrRI1bIHyLjt1gpj4V73blX+Gvz75MZAPik4RKTpDS
HEMvMz9gUTNMZ0C6jMEM7NeSeMwVbXDru9REu7kTVRE6FAd3HAPOIJ9db1hWxMj0
v1PsE3GJ60fbNjS8wWZkTbpadZeOp5aDfkjYe71L3Um5cChOYr2mgMPeD1o/joeG
c6/dd//Catj2+6GC8M84CpALKr6IhEaY1HmM1xk8Vbp9os0fbz34Uaq5dmn74bXc
3nAwNOmKM0b2Ad+pw3FgqmOD/r6aJXCRcznMGZHx056OUPOvqfut2Mf9Epz/jHlq
QQt8+TXXvPQCBYHC7fb4D+BnCGpHRF7RVJjQSW/kjwODqsNH81doGrbgrpIlZZ8V
pDqIewWZ5mIlyRJ052+YunGAd9Tr9yGzjpdHy6Z5nhogMZTxbhh43ViK032d1uPN
viaXOqcritRZuNJsXd2Dayf0PJEPclys4Xl1zuK4UktTNTm7fss6pOTumpHYO39C
LijHk7efS0tHnbcZssDOnAO5MEzsf6/B34Z3fL4oBQd/23528XfcD60UtHF6E2Vj
LoIGMTkcgV55hiPDe7njQVzRzn/IugwFsIYqYAS51GjbWSNffueAp9+Dc8+5igcN
NPG2KCABIbOO9WwUJajWDREyphhQM2IJt+nbXBv3SkGeixUrZPXonH31VED3N51b
ml2o+6H66geYv8U5bb4zqxRv4E33p1VAyCd6dOfG7FL/8kuytiCkMO0liYskbYlb
IrcS8jp3GKqbXZ0iXo5pzmi42nPVbE7Znk9iSkTDP/VaCjPyY1ScaFyWHea5A+PZ
bOniMgtXzUsdWiULIZUU9bbsITQsqnHZMVEDIPBQIZ6yisjp05clGPvO6FKJ8coZ
G60jLt4kdev5eKKUsRE0qIgXE1fd9cFU+WuimesvrVYn9J0XWhqguuG1PpTEjYDz
0tZQCqTbDWbpn0vvXGUh3TynXV0J5agR7huTg1ZJIPlAnGyxKCoeephdKga4tTXH
MsmU3nCmRJup9haCJuLEPIf7l9tDy8+6dPRtderDTbwTc3uCGCMwrwmE+HfHI0dB
d4CqIfgic3/5LE8MkK9m1meOugA5q7EA6Ng1IFjZOcllPZ+RJtsEn0euYnIN1auz
/qQek0xYLfNPWZPL8g1aQLXEePddnZI9VfohbRHyVk0RwGP61WfPz3crtGfFmnXZ
eSMqHTP3Rg1un5StoDiESUewGVMxMia+10JHuI4VUaz437Of9gEVUha0sxvijXNM
Q72Yvnpw9sVOafHZFPuwYXqVW+MGGoYzPbF9CyDpaCTV0L2koc4HHpZuOrk57U3z
LucBebCjqYQHYBKUStA8s2p4rYgsrzpZ3vJsAKw38f+VPx64Jwpk6Jj+RNESQX5i
4/ty+hrPOYeJ/NZmfxIU5bkTww9e0Dn6C71CpcnMEC23mjv0/KyP9RNwj8vHxela
SK/0U9PpcHcSQ8TCaXY/bVia8+zpIDTU6hZvdZl0JHOiPcs42v2MPRJgWXvj0S8k
8P2EfFJGsHpQ+iW6MspdDxn/SHd1E1UbbJzr1COkAWRlFRpqVpuG4c65nPMJYgbO
l7c2SRmBPlEHIFkLxfevIrmEpnUKjIbZMIPQJShtU9LKmKMyZzekJWB6J1MXlNvg
kitau+ww7GbvT56fE9dOWWAD/79XMQLlPyc0M/TFZpeAdYpi0NgQWt8xv0+WK0x/
r+pxthe2vcfwi8qEJenLGsnETpI8EinXGXcWtPVFwZDCRA14fvzJe75aokUtIL0L
WlY/rNc6yx2wIujT9fY5ufiRwApv05FIXgGiNbgyZIdcZm9K21nPzmHz2sIIQC+h
nsArom+Lodm8+TgOg+odSO0weXfZDaFILzvICjZ9JDqkNrBy02NZu31HFQN75Tdx
UQBQxTBSirbmZXhF0p/Sh+y+JMB7u5kIiSac9IuRK5TL9W9xAPDzxpTHnQIUxegP
rqbfNWInj2jL1m+kPDP6QckDN3H3sebtx9CB1MJayqT3Px6CmCvSDzp36+1IWIJS
YSa2cP4LdJI+KlYhKabTSbRhK/0wftjn46rLWOhebFY1yyxJTZw/y/0OO1dsJsV5
y6ISJiRMkeFMcpOJxKtcoCeV0DkCe2C+Hj2r65Ij4MKnCw+ohdyWMAP8LRNvSb5g
XsvN7C91iiT0pUu343GN/Af9Iech13Uk5DBhE6wrGvEqlY7f1oAno2QR6PWQ+bPE
Ly4ew4aEP8R9p7jBLs5lOklpE+kRmu5kNoKutycXMMKY1abNaNZ7su3Bx23LHzGL
IlcYqJbQLzDzBPc2JcnWdjLU9W9+SvFDJPwsIlLWg1gykePLugmt9YiTlto+aPBx
DkWJ/sfDhii8m2YXgHWnwXceoJQB4yTHBcCzSamZ9ShwNZqS/0GJp2at5JWe9y1m
veMKsJEFM55Y7NznYFonm+YfbJRP0rbbG1gsJu2BzevHh1VF5vI4WZ4YJvn0rcHQ
ixPx5t80WyrkjKIAE1dAy9ucuQNqsQFogVTQiN1cmBOa0NiJTufeC0DBh7/k+h06
G4a2r3+z6BayxgGyZ7YHx3bW3gFmwzvs8aYJnmHIKO1Jvv/45D7mDXcVvz2IjxKg
c/wNG61Hko64fqiVAmG+G401oaljqjjUPuPExbPFv1za95Sywpb5aAakAbP1HuVc
2OPeEQWk57jky5B1ht1tcU1Z5bMNQ20jTdu5hsNwDMw9bmIbAhpovwlqsruv6ZKH
+COzTlZRqabiQcmCVKXAfp8j8rdZ1whl02AAJLIGimHogQdrJE9emahmswqTzKno
zUn2w07Lfy92NyyTebtitnsN5COS+Mft/uWv3JUPhvp8Kic5cF/DZgIE72sono3Y
n8O6g7/d6UqZzfVFZ2KTV+9qLq7XgWwDokuSeLJvdBm43cmoWz8wXcdOAYUXHcw0
MFBNArjDNMh4IOT4wb9fQfQbqMpkD+nAkLl36PCrj/O9wclDpi7GyjMn/oQi5Thp
1hBEv+LslW4+7j+6tGf4y7otq2/KWmEwdT+udWX64CLmNaYOESK6M6sMFRYxgOku
xSM1gypi0g6w9bUKpTBA16/YbcEXuKn5T/ua0wXK+rnAmeW+ShAyV1uv7kjtU69H
00aiyI3iBGwiOnU8l4/Mq/1yLGm7fyNFieuPPhRvw0fUYFF4NtuGTW0DQPeN6dbw
ArEGIXI4NGk/gSwW3LHCycbpmOlwPCfm63TKWpR1hBEfkBE97hLxFeBdVMc/zreG
/0bQKwUJO3oTeJvWZGe/+cTYpcv4OLGmWLSXrN635F6se9iql6TEF7u9YYjC54mg
uWfBluzWL9Vd44UtioqSD0YqrRAffOihc53x2KLyyRSu8BR5vCcOhKLfFrkZfKj+
parHWM/X3akzYLyAS05wE0M80bfUBfMgrXMKTUtpMA9ag5XLbLFOUaxTt3EoVG0V
kSfNUi4A/KxYnxAMEci7OzC1d7HE0bjtA21QLY9AGNKJXcgT6yuzJtf7zxzFxbKd
OgZHuqc976kjRd8SZNvF8+7HfGBIXyluohuKeHmMCkyLB6yM4SslVbJAxMBRtdeb
UjSjmcV2QmjsCOEUye77h8ggvgYoHMfW2fWaovoRruZoZ2Onx7HyVCDkfz8RJgNu
ikXGXlK0sOkeHoP5dxjtpHArd35ZQ/1pu23ord1GpM/J1Ulj1b57BqwPoKQ7T4wM
N07/iEsIwGNMUsliV7SJ85peSO8m7/X9nCVBICGWfIqmwybUb93mFt4A9vVwvL0y
BH99bH7cJF5SzN5lZXgE526d/hvmPWlL0+dmP2+RHYc2txWrdig1YeRGiFCmI+rm
LRjxk6Izk2j9Lb/0Y3mNtthGMrmxiiLiZN3D/A5ZpzY6xYRUHAaMG8BW42RWIGrD
zuRhsny/FqRIE69OQSbn8e4cGZTIkd5HeW9hG9s/GGj4SCu4OWe9Up0F3y9ojCgD
4v9SiWtDmYlzazQe/3p0HFdamZDM8xc1U9SQQTONxyE64l++QT4Nn+p3uan2669p
Pm9sPxGEQJ8FasfFbEsLns8Yf9AH73tT/i8mYvS6zrTybivigrHDHLLhNX5Nh7du
zxlKxehM5JcZW9rkXYfWNsMmL8/inPYLAaPgV2wLtB3xkEK23v4G8NTcqH7uUQXP
G+ySegAs7vXl58vm+kKfOuK6istNiD4Ct7VfXr+dFgo27udAQ8rCRQWmzT+OXoy8
wVgf5wAQPiP19Ih6HSQo8xSt7FIxkKDfv9IVnBfXeBwBL3vKBaoIuBGL+hoxNShR
QDlbJVXoD1ksfdWDJtXcUFxws71JgrQEPfuaKV6VUXUK0j/8dqBXLSFrPVzcZI/V
tP84uyZ0u+itEX8bb0ESgaa+mCU39hDxAENYNcJ6v8afyKTCbMJWoPHisCA3XaF5
MLCpJPpLEEnb5xmJ8WuZiPccM/Ow/cGlovHWcjSbLcD4PU2mVMkcqJGbSWMH+TdC
2ajcB3B+4NAliJlP5VvhoTph5cTkNg3AP6B8H/kmcNZcbkzTMBGN/yCo+iwWhG8q
oEVslfm0tvGJZ/LdmroFWAG7xo+oiia2Kl0FEOEflGD/8I6fnWcQPBRRsiqHVr58
blUoJ+u+UP+Qi4DhP+UnvSKwtGReP9aE2k9JEJgvxYjhFT4RR9V0wryj7X3tY5kH
rHm+i7umvvfK5oFmXrG+Tp0D+dNwWJC311ll3zglfeYpOc427JNEfMccxgl2OUsG
smkEb9rgq9Fwuc6/8HUbAHNiEgEVpcFnTFuVTbwJqrey/ciN16yg6L/CQFYZzOSr
iG5gi4IGBxBy7/jy6GQPGf4Om5vUeTltmkksOoioe+cNbFwiF5a0GjFY24Ltja0h
5OPKGlVi+LUtKn0dtcPURzSEyqGM2VaVoP6ALbb1SyzLndXvi5O5jUAwGBEIE+VO
hUni+rOQL+VPJWPkslIXEaAWJwoI4FdnkLz0w0Jm7FGEfm8u9/FrXKn8L1raBKsO
POUuZxWEFNpO6+7vfuwdxATSpuoEu4K1n2o1n7PPHqp9tyM9gjKLPPRKBJBeG3bU
qWKh6XmkcQ+hAjJi57f9K9q/R4KQXkt0PwIPS6yk5viq9tPiZg7aJ4awzAHp3OJg
/rO1wMVk9VA0By5JuXr7n9fyFWSYXu9PUsc098YOoIsp3sGlATs2jHbPD+A/kVK5
IGQLjrvIStwfCOSxna/oXWI6LAGyVG4jlmC/3uX5lP1D4AgPVYAXAVy8JQlFKPt9
V1PSUPwYp0qe4FtFbiPzo5f4ICYoRllyhbMG6kVk9nfjkDitCH7EdZobS7EicV46
YxW3Tyy5Wipt4/z1QlhXpYYiSmYCbdbY4Q04wnbiKVdSmqagy2hHPa4mRSznWpWH
DuVLAFT/jmkwtp5ZB/NwrdqjjKtg5HJQ5xb79QDlYuNRbYMHGvg+/mZv1+8ZPCPv
ufn4KaMplNd3rYdGGzkW9v3d57gONzeSRsbAC1qmIisTN81V6/EqDK6MZlFGZglH
ik4hYvqoJUjqhso1SMd4y6E1TkZy4a8qYdw4q7EsYaCgbKckY4/nvrN9UwPmeefk
BLUkzys9aRdZApanwRu152JzHrmAVxUF3vVEkXNl6LxEmvIQSLPiQ0Dg1S+LG60N
xHdPwN+3EvVpFv4zRB3GnCmPUmMFkDnwx4E4PKZ/Jv86uRrSBNNb8gZzAx9pAdfO
a3pcwNP+qLDMspfm4MmpacLYKvv5hhqxg5DKu9FNjgddxGLykO8mRHHifoyPl77J
2icrK6yPgE1XR/bwKqyGrOcVurhLU/3f1euyBV8rSAhfUwRtyHrqi3+DNvH7C2Xm
WG1F44cssmdNXJe3f89P+M6hfGXNHEMEUd9CoH00xR0c3z6HoWT6WzBrN4CATnSK
vf9BpTepuKkEEz2JhTOF9hVMYPPvzu8fukDtwVNYxRhusXGIj9Ly2lHpx0KFdwME
+4Ix7fFdBRecsUeYPx00sCHh8jXOwSTUQGxc8FHN/nRO9+65F5+Ex/zvoTLUhkTg
K+nrxM1BMA6r56MIA6uC31GYwAYMZZrvSjK2MOmJUI7C8WY/KzGCKUi5+TcHxZFz
TtX9Ew+VdTkFdgARZM38nMPuN5mYkQnWmeIT6fLrC0adn/HXCTW5lK7UZAC/ZgBb
YUrx5evjPIGufBNbuXNn/d7O7hKA+uQ7wOp7bJ1+gyDHwHCGakUZ6NMkDYHpWf3m
iHwWREddAL8Y/ZdXDXG8EYyFqZn2PMuVepfyBHfCaeLIXvqCBAu9SQSWip4yH5XE
hmHPY3D90YcXYrIwkURRmWE37KLcqsOizhpo1cISsi7SG4pVfFEGQ5CRmGax0A7M
7AcPb8STvg2+ljucqsEITvzQknmBSS468xm5mfJ4jKsbcMkiq3BHlL81DW7pfy28
2EFQhlkJ59ugew4dx0YF64FbDVoOjerFo3vYqLKAcUy9LkzaHfLEEyPB8XfCJCq1
xo/lwcXHaAqAzynDY46EI4bxEGeVvdeOdx14gvuLKOg3yrK7y9j184/jwqgfsPQX
93Knm8dKrXsCYSobuz09vz6Y6msPW8sKyrhDL8q+2edom6R8tbHhDRXvvXHkqDtp
1MusNaYkh8uCCJQiCWVNbf2XWO0JNww6o4yofPFNig+yy6nAPVxnNXNmdGJgY9AJ
MZq8ItQiEsHxRTN6y+YoQQkL5yGMcD+Tsq/YcYDWvvfQAYl/1xR6Vo2Vos0l/bZH
RvQbVzklmHuIiQppCaiIb3OcSIl/cUzoTaHJxl+kUE4qd4qUa5aAtN6DM1rXmmW7
h1JtpD8Dob6NlMzeKvywksUCFo0VpW7iXGG5nfW3IjftNJ1T2IpnXnTz51oI6E7L
Zvcq/asPa+TzSGo/gr/O5+toOkiQXTgYx2YxHa61HIgkTPI0SDwgeCt6dRvM9r+y
3RA/QiI8n3Pfs9ZykGXmzxJITk8OPmIgWdHlssk7IiMYtS3YFebz3ONZGyAmjuHH
YW7pBR0Zt2I9HW2EFezc5KrScfgW56OK99NckoSsdgdH+LelA+uBEXJsqeBIRv0H
a4dUaleDyHEB3X0qup0JGOm7J1qsvT2sHrbiZ9See3NiEGPbRJ/o5c0E+xwJ/GlL
1MqnRs/qSTU803RH9eeVcjYFe47ALHHvlcAnPIa21PYEUss9uGpgxIF7Ii+QefUC
i2q3FgxqEAavt8SoQdzmckp0j2+0gLkA4SUINQYa6fyNSIMgMFbxsGkQXYVdryOA
6zbcjKVZP6+Qhr8u2Oobz6DFXuuxItGBxDWkI1/0r7q4/U+QcoY8LD3oDNbJbxqx
t4fzJOsW16jZs7z4Y5mYFbG4bjGu6KwxtqYu76WuC7pbbAFtELcdJmta/FRI6tak
JgI8YmAn3bEhbMgcYj/reWn7frQ+USTaDmOSnpxKtNdN4yT1za9CgHl8d3c2iGEF
McENCsywvZHg96SIvNW8QVIonzTQRbkOgzrLFP15CPO6M5kcsbh7vCFXlmAD+hAR
qFLiGnR2JDOoJw1z6TEKh3EXLrUasfl0QLtnSJReRKzQFF83ovnq41mzf2S6Wh3H
MHev8mv/PuiUgnYGvgxoXPvWWD0XdwmoMrmgyvm4zHHg+0pz+fX8n4uuMnzeQOs9
nVr7+3Ejw2H+NWZAemHLgU547jLiI4S5SDu9PelUreh1vfa3fPdV6jLncxbletee
kAEzmch0B/R+UxcdUGOt4DC9XhnFvvGglmB6s/CLhWh5av3NkSzffq0mVYS7EgXz
l16TSBoiPnF0Ps8WfjalVwJbgRIuOU66/evOtjugRzmeHkLjLWwNdds0kmLb+xPx
Y9PJeI41+wOKJs5LybQEkZki1PbbEh1IT0L2hNZJoznuOwG0KX/mpiseg/GtCqSt
GlOGDp6Z4rxQScbDVcbR/N/1Bhi68ShTVFPoCTpKbfbupDMfy9EszQ/GS/5T90ss
TAR4kRxfmes6p2AUtfJELJIfmwOSgkpqdN4+H8nOlhh4B6q8IdkWWAn/IzrrnJIS
KvVQl8GRjEzLFQKewmvOcck61zgNv4l3Uc0HZa6T/OQ3geDQ5Fur8yufRjST+khM
DQyBUPqwha98kwkq4F7FmHa5Dw0jBsdzLEdye80EPlIlu2CoeEdQy+lYDFWJjgaS
cvQaZNkGtHmSeldrQuvobCorcE+XkUuLH/7/dtLhw1PnAWLsDyHEXEhTINAADahn
pX5PJUTlEWD64y2Qxw2aKY3NyJNNVHyp7I6grmGrbBDC8IXyTsv74wKBomUUougD
K/HfFjp7kgZrMgmYB+IpHBsjhBRDxYUNA4AAV4PZDdUynml9hi8+WTyRWgTmRiie
zXMn3oyWXUvENLOZL8wat6ZXF5tbl60ctMPAqFU0BVI/1eAfnQ9B0XLBPCi5WFZb
UrrzU87LHf/CitQqezlSliwpfFo3yvM0tm4ENcggdxpDN66+/W9ZioEQhIpZtOcv
cGH/M0rN4wMe9DlvkRbgjNendd7mFZJl6z1UbAIcw2Nq1BO+vnbSjlqJ2aPkvXYw
5oBuUWV2CQi0Vy3Lnuh8vO8EQ3AmbXvoXi2DKR0oUn49TZYd2lh6DdvCSOmcwAxo
42IqZEls54HAjgPYzhdef6+zQTqXawIItDYrIL8bEYaykoewE+vlH5aZmTMjC8zm
CZk+ENS2lZGnb+ZoBSMSziD2MLPAB5V/7hVxiliJJ7TrFdqDYPQuo+NeDlZqlMhp
CnlmTl/Q9W1oyBXwMCCzmS/foovgi0DID9HCHd4hcIumEAu3LpQAZYN+6lV/OROM
UN9dDtgW+FX3rb+YUx2pFfS/whUqFeb3/I/6uZ78yvsXbJtLLUF19w65+ug13QmV
170xqKkkLtMAJjD55rxuDFB5V7cXVpflFByAfythKTAs/+oroHrb6AekT8ABtGIR
FgzMVexkJAbXVwWqonsUHjJf8T9+Q7uV+yw3IUPOUiiClETMBVI5o2AbwtHkAxgL
bI56YnocjuPuTb9Km4P2b1PyaPzYV570Ar7LtB2IWBXKojZ/bDpBIzPoATrIaOAL
aG1V49NqpfjD4dYt2HzrV5/Xma6AUlQoOjDzw/F78b0Hk1BOBbklKFTm2I+Q2G+P
nVojyCUOvtANVbbdZNGBhxJQznKmGhYDPBsEz6w/nWGaMNOxneDVsCS77EUWvcxs
hh2g4SDL5aqPB1/CAs5Gk7qsNGN+GC9AX/iIh+zaGHWMBHFTK8zK/ciPKyFbfQik
QCM01NFUFbjRn+TK4KHFqUDO2Lraxv9SmNcpXc7NDCDuvz0QN6pz7Nq7BxNB+rJZ
h8MnyiSjETUhmid3sWLbTfOHkO1IYd1B1EuKjij/UNbVRB7B0r1e79AOWYOY07a6
9yWbcQrL9YMgufvFNtueLNITWNsJCC3MQCZ/+hj9xnWfum27PPutsMY9PgPilXUJ
DyPfP8wlz1idX6mCixKHgwELbD/FJ8Br64aK6WoPOhYP1DAnxxjDrQKf29q4dVPc
UcmajiBxLxyF7anbqS42W5SJpaJNMFNIKo6FfuQZ6QHdF1HUMGhvdbR3q/wI6jK+
VtOYVqvOKl/496yitl3OGCst9dbjGdLDaqhHbMLoZRw1CIFwVWoVnK2YmY4yGGiI
mXWqXV1wzijijzAW4uQc29sQLMdLTLUvj4vbQwGwWhtUWkg9T2FalYFN26iVpivu
xx+SXc3fslePjahUYf+WWdW210Dx1b5JRpDRiDkG3wNllpgv51BB8M4bzrNFwBfu
KsxCmfIrn6GNJ8d+2DS3t848qr7PTg7V4wcoZP8YEZQN6CREJv5Ey33Ai2vhJHW5
+5YIUW/fiHCKcS8yYYVfu51MLcL4GpYCbfga/7gfpnGyU+LaLRFCbCc0KT4E7+Ly
FDXalLl9f8zn6P1kuIDa1l2rI8ffYkLMb+uRp6X9KiF4lHg5fiZSiMlyN9FDC4Jo
olhWhAd51kDjun9KAnJaEOy8RwtFGQnStIjkigCMiMmjRUmWdfowTrv+Ho5HH85D
hKteIyIeS5uApx/28KQ7NE8dYQ3Y/S3a38S7j3WmEufORSq42pB7pO1LZheds/zu
b8bFyQrO0dc61ZzzNsA46BxXEYCptK7cj/BNRTyD2CLbj8xiUxLEAbU5wcXCQgeq
BkPuhDT1EczrzA0ARL4sNTMaMRZsD8gYigW45yycVItQamp2IG0WzUz+wfOeacrC
aUo6FDdCKoCQvRyB4hl3MOau/zPpGYGD7coHYGYA5WRxXnjLOmhpNoS8FOqnuzs4
G8oFR9kpNBL+5fPwWBdVbGQSaWS4irQzr5+4zem3URznrbJkyxyID4D2kFdlqsVo
08Ji0vqh/U7AkwKrkSSBLW9WigSUP0Ga6qrs/snCCYehC+bnAj5CE7/oFTeDvydF
3c3pyLN5kTyK61TfCRVnkBK/abe5Awat1jy+nudbHx08bTiHqTdOaTc7Gz5XXq0F
+kIbU6mPjh7lPUEhpbxzvjO8M4VFfsnsDZzm6l5UP0TDcX4r6m4WUq3ap+PUerbZ
HbKO/MrdDnvH81YYRsMm/TRmoWoHqFC7DdBWpBcw+36ECUPUT12xgfuMyoM8NybY
Ain8qRyIIpwAaqwfWX1cy/3wr+GhkF0sR//o3ZU9xHwExoNTpEF2ol6828Kp+TYb
C2eVBTvqhR8GQbqWPGlIQv7q5z8jL2nZauLAj7uHAUUc+Im5H/JNQEFAAHsz3BR5
oEKP1e5Zk+iVEh0tYfmR/MAM3obVgP1MyWrXV9GAT6XOzlhrhm/p2wS4/a7WPS5Y
S2uqUgMtmwbKgxr6518u82PkSFN1qNswlWLegTouWGvomjBHvhdnoASrHlbOmVdp
/0oWM51+AvBFL3ZqlhJksg9ziIW/5n1qj0QDf3o/OAGw8zCsN+HgEreDweNcgi9i
X9u0kkM24JClc9+jWzSlDsPcEokWCkO5B4PC0s1Zge+ThtPlcK+WYBnBZhwOKAYu
ts3qPk9pk8B848U5g18QCnmR1QfU8iRFcunTOWDimhylnZw3yu4sxjnopjAR05xX
+NlVoj5x0q62apPnbBQwp3qrYlf6UqJz9ieNP2ESYulhQlDWueObY5f8FRghxbdt
fOzpeqVtFRJHH6TQ9VDBgspqyDOKfWUrxlgoaNpgVxC5PNTzz39duVvx428APNzm
X1asl3y9EMzHCw0Xm0NXN8MuGRSFf8BpKMJLK9cy8rR+WQtAeak8CE9C5CHad4ne
xdp1NSDBYe1WgOjsZuxSeihHAKHMs0iWd+hH/OLcMNF6AuP24xUO1oFM8eOLHT7c
oeqsMAe+eEq9xqsBK/ENLHigRC0hxqsdoxQajnAyTcFpDssnQI4kDpSzA5I5+yDF
oVgpjFxO+fLhNyIRmzvXCkiprim9Q4PemukUc67MtchhoI9u2fCcexRil+wu53qV
xvcjUErVnTV56Qd39wATCm9ancz74C+WC4oQHewa4jLOgQC9l2ywIoOzRVoD1jde
7SvUovir3lAqQG5WpM5pDuJEiLjfgL4oYR85nGKsBY5vwSOFiVESRnOo19X6cVDn
flC+vybjIeesFVUCZJ5mH/I8a5HJe9zUf6IF6JSWyaz13aZQNjfcRs9SGK6rMqHe
DyC87jsesBCaoBBri03Vk0oR02jptAn1CSGhr3QetJ0CG73nxmz2cGfiXqoKEG4w
cN8ubFLU2YqpN/HTgCzQ9IkYei/olcMa4fJGTfxN7DCMtmNCmILiAhutaUNzv521
H4h31tFgb/MHxMzz3UYQdBhY2zVC9c964M55vHbU/Lx05MGJdHPWZwQ61wviFF63
Y+uTXDTpw8qmyJBjTfs4zW0wVu3XgHogRAriBIgyDrlDgyFnuAlpQ3FCtC3LLxGj
5IF2iFxIA0HUxITtxkQwWczK5gqUE8z1aB9b2VaDY7lbO+6Kes//P2QX5Hh4HwDu
Wy7OOdfygzigrsB2ZFJg6cCQ9i57K14tSz447Y5Ahm9h11vDbNBo01EnqIqhvH6O
e0aePsD0sH4oWy84qg0qtLMPNDOyzU34nk/W5WSEbikaqmxM6LrTVb/ZWM6loT2y
/TjgKU2OQ7Rfx2jnB3o17lANPdg1sRHg1nZW6yzlBGLvlNNAL+L3MlxpamdwrM3t
8OirQ/wK+Sp5mkLyJVxHj21kuCTMeZqRL/lSh3ClqI4CTKWyaM0FlrXcHGD4eDpz
C44omfHHj22MAdBkyQKskUNwHwRXIjeehrgnWpBu4HZC+V39i/WwBaX1EaCStvhK
5LOK/T/8GYvbDy4cfrxrY9HUnQ5AUjALZstKejlBsUtTBdbWBeEXHPhaqnl6mKvl
LQkfRZ60Miuc5B8ZT6B92/4vunwgHbG+z5u7/iBdzM6xN9+sSSO4k5jMVbpyyIOK
ecOiTLHjF26s2hJ22+iJ6sccOCMuyhyIHAzMSUpea0kdgR3iletIQ0lce397C4k8
balj6yPMM4GkZNf4uhhOTaGtKaTp7xXI6qidBc2sOsobALYGjHY82w7SNvypwI//
k8kBPPVraAlakRAYDvVUuhcAT98b84Qp3onbmegxoSJzVXAIQMaye+QEOCAp2uv0
z4+nPJ0sx41OLmZY8TfT/zazxZo47Cje+rPuhWptwSM0HPYl6+sB2qq7iqMCX8k0
hKRG4LvBiHK6E9bFzcboOcPcXMMRzFKrFU00mZKYpp9er9m9fLrGQrOZyP6PabPM
UQuebsy3v6POqkffl+TjvtWC4oEkCE5Qd/pH1K0V+i4Ma2LIUhs1HnJjat85d7iy
8DZxrrdb/AqvMcz2G5LSq8jBed0ECTswb6euPsz6IQMXfhzI62c+q+vjmVJGOgsF
RZe5ivD+IQeZiB4P+vEgOerua6+PcMPbd9iiZTkvgqGMKfu/WU0Lgx/7BsziGEq8
9PMlACtu5HJwqaZcbrQW/SZurSTQDdOiKiW/6lDUfeBEj7cQ1dvXIgWqzZGOVNoM
T3c3wlWXFEOqa1Qeir8Dk+XH73xAeC0UtDNe6MzKdw16O5M3zQt8AVSUlp0Yv3Sp
jYRI26PDH4NBV2GTuj0FqAzByzktpP2lf08Ok9mXq7FyRHGlzupiR5l/kn/RTcPu
zqP3zB1zSpx0QYTZHql1Jv2WTW17qwWDFI/kTo4tmW1rPnJ3tTyp1SU6+9K5Tcv0
IpntxVs8lbZWnC2yIlSepkr3QYORAD+4F3G6ZS6VQ5hSg7/ZmjrGgdsxXNu2s5bg
43f/PqQZSa9MrrJwBQVlkKIoaIAULf4FKY5n4bP+6X+osAZmk74WlQw7Axy4rFIf
dlGxO8xqrz4MAk1WogSoWvobZuHjKZTcgbWILMk/Mebz6TXZQCJC2oZldX4hCivw
1ZCK8NeIckA1iWoCL38NhcnMKKBvz6rypJ0OSFhFfTaWdTAKWWr0KxuYMNRh9Dmv
G1RZwxViuZpEVMW1bd45gEi9wqFPu+iBbPIRWfaeONMrzNgGcHs1HOWsYtX11LKu
bDzMr8uvaEFUj4OEPkXTl+9ruLlqjY5JKISJ8jlarIadvHDd3yhQ7Hx+05rho5tI
riCK+tVUlS29iNrud3n1wZgzerPyL0pXZpZASXRbTjvV6WXXBcIZdF0f2oNWje0A
s9NaClxuodfXsIDuNBSWeNMr+fYQ+9aNuGEnm0Hix7DrEGDIo03pf6Q6M54V/QAi
80GTWi8oT/KLCIt0v6qX1gNsNGSCam3unBpDaPS4MXCcHObbshE5cE6k6SILneRg
Xd+2uim4VrGrW7up5NQ9uOPa3h8X9k0qBbXZzoyxFxnujBz+cgNkqJLk2BxyCdZF
SS9vjoyELBBmGC3zNGweMdoO2N2JLgkc5sR5+EJVYu79FE8moeMM9BJTADW9cS1r
2l5yZfsJXqCqAIZgUXPU/kiMJ/4LwTh3gcaOlrAoLBoSrZQsusiWMCHxmStPbBn7
yDncqMOWBPKF8oRwp1nPNspCPqh1b7/FlDAEr1RBWCLKb7YNZq20KVeYHsFdHFQb
UgPbgfxQNVDkp//ZBAN6HLDaEosVKdX0oKUG7SMhWaADr57DXskUCvyxVm/0wUVl
9SSf+sAxA3XAlUmZwBzESmt3uQqYpmFoUMh7HKxdUnMAkf3nPWs7nxQRlfgVa/7k
W9O2S05OM9jomCtRhrEQy4l7YkFb1CQUAtRl4fUzTBgu/FhuyKN/tDgC9Y0bfmi3
YdeYoqOOhc9e8oTYS3vgqoX9AmIszz4AT7yKe0S5oKXEG/jUlCpAb2wMWZJbwIyL
EwTkt2MUDKbYPWgZpZzy3SsPv9VBZ2MUypmtlJQug25xOe384Lk6CL7urhUtWdPL
xmL2Xe4VpH1JthMCXJIeOO6zUaKHFhjIkjFuWr00nSi0AVwKkuPpNle8AaxXZYe4
oZXGemiXdssDYw8hfHIZuzy7503TP+CHARf5L546jwzsU82hNEZ7KlC5ooUq6hdm
7aChUxSLUZeTnZJAjz/INZh39gOzez5c261yGVCwpzsLXUetR/VqCSSky8hXZ6ok
/DPrHtZXVCothOM+n7KeQvIUzpAUvZ8HimeoZ0oU5PIsGxe03pDs8tTDZHHoYgv6
Gl0zCx3C2MO+oEUwOkuNvguVADMzu0uljlt15rwBpqnddibWsK23bI4qDSNMUoue
VFj+7WIaukk1Q96xiM6JP+9MeRRcKlFiVs4HwxIPnqeDUnWZvY/q77bTa+6g9EDM
vQJWKUsKnF6wb9N50mwUZo+AWIvqkEgc1AqtL1WxwSsvrT8cx/iib2ZzBe6Nm0fw
4wiI0mnBbffNhadVPZ60KEs8F7Yxpit3qBwZHz5qP8bVYj9SjJfAegpzbxAL08A3
DWEC2R3IibQUSD4VUfJfnVURguzI+Izq1lB80HA27no6QCE77ZRpThfPKPbQElRM
CX1TzbfhonfGlOzUokJavKIz3AFZDiajon5EmQe9bKirLlLVWLbEwHlmVtNztOSM
5Fbmr4FyXg6JvwOwTt+1RbQukB2pwbKj8PjAvTl23lNRQF8akCj55QBLe8ep4iDy
l0V/riBUvBVJCfHkUmNRtK5uG7QDDlFxkPamg7Ijpn44ZUvhTwR6KZAZRQ/5AghM
t+S0peg9UEC5DPIxE4n9iWnHNXbyqMI/ZcZJfbc13P+JR/w81jwxRjp2THzD48sz
EC8kM3P8OO+BZL8PdkuzoWMd2Jlmc4S4X78seMWiXemN5m4PhklrBupJEUjrykjt
Dp5w4TEaECbYHwb4mvYNpR4V47oKGDADqOOizHOVFOuEaMzMtEjtbsOJ67ypyJwt
MLT7NCiyBnBYqXUZ2qdoqzWTCuJM5r3S3BCuVu7OupBJy3W9+x4EAMuOeC4nuIjZ
zdiHtY6qeh13muFGhyL0C4oVJxmjl5R+H9ffhwLTNX0MWk//F8XwTCGgJ8dvqp55
gnGARYltxSh4Xta49UDJh58VyqWihMa1GjJmcd5L6T1t3vG7KmX85fwJ7cAQyvIp
nsL05ckyV0ZxLxN2MDX8qFby+ODzzXWofPx1ya2i5QVJaz+ddwKjFxMaCgzxIaHo
BRNZF3sMc7Y+TT7uwwYdx2wEC4Y++1V/h6ERIIvML9FI9bIbxNRlNtVwAJZ6osGY
Lb2fvtdmJfPMVmi79SNh1z9XkJHNZvdKm/2NCjoyd4M8DV0RZQIc+3eB2NpBapAD
Si1lPK4HL6UfJttYxfsaPSilUwYNMX7YBrCHnp0FKafPuy3I3nBgF3XRCsClpB/e
3SuuADpWW/qAwv79nmHx1caumClBeBWYqZ2Lok7xQGIFjOvJJOr0UwDyOsCk99yx
y94ywIflzifigLcvAY6MG1MNiZHsD9OmhLE+gRIuuJhwh7n5pLVy514pBHZ6PGi8
/NdimQmuNsDkq6Opie3smO85AgVYas729J7XC25ht5xDiJFSbaUq9ZtQSfUk9YOa
8AWMEBDcVT9qWfo/eG+EXzHYpWPfYbMpEqLgiRpiXYLJF1fiDCnLfb3kHtXILnPF
oErkih/GyJJH8DhkBafMHQgyYvgbhV6mshgVBTqYdDgYVpoDOKDXAeFKhgOJDYUA
ZCRDCKDqNy+i7xff7KRyKEWaIsRcpG2aEK2ilSwz/L8QC8pq0AoBlwEDDCAWblDS
09AEuuqPFW9gz1+PLqyBJk7T5FXP87pda+B4xeIJFpz+NsrFMjxq9w4FX8ddDPJw
rhLH3OQcECa63hiWK2ve5rS6FkMQJrwAqVnmyz3xbhTkX6UsALd1TTGLglpr05Yi
1kwLkvzbFogu6ONohDDt1DTnNvQ1PmP8Rhfkfi/UH71WDZ5wMMU1UJf2pnigvEOR
VGGsZBGjCEyFF8AE/kaFLB6+xVakfPJQ3tC0LwJCrI4Q2i4t3qJlLIo8CK+DYBeV
rZGhDnyrb5zreXFU2dL7yafve8NJHtKjqJYYhTMa550mgxArw2tWA8NKmPKm7UXf
55eILxo1Yn9IzKn80erIoFqPOmY9TQcT8GySHriTOVsvUC4kusMmBYnpqO5rezFQ
H+YDlgUi7xx/Dihy790rDI7NbzamKAo7RO3JoGIBEQHNzpFr29gdVjl5O3zdUVbK
jJDsoNBGpm6TRI1ms5tyrHvwT1gJl3W400rrBSEXJQe0/I8UGVTjZ0alFnqi1bYG
R14lGBAPYSBGUEBgIBcddqyexzskWNTBrooZTWNgZlYGUIwkVsQVnEd/xAd3bPfy
p+l5e8WwHLcpi/DKW5uGDzRj7xMbR4bKnkE3jeYg6/Q3qRrP37x9CQvedLUBGYdF
daHg5nWQn4be4E/65idtcRN45C3RNmz0iVgH8Q8b1Bk+BBFI2UL4pd84lKfBMXAQ
SeL2WTf6QRP35aQFLyaCsB7RWdZlX+WiBOZ43cIDt9wh6f3XPd+Ur37ZAZYIQxyd
TYavbHBgprLP0vUyGN0ye1W6Hex+dUatXRsKYJfdF3hcrSEyOwhTlYC9rIL8bAni
OBYKuxStVWi/ON+By0YV3NqKz62hm6ohNjpuv+2fymr74zNY6MMwIkuI+h2ILq7z
bkSgMzozB/ykEfk6ZJRu7pV6QCcXXO+gKq1AKDUN8R2J0I0OXcy9JPTwrD19v3Ur
X/YmYKncmcuPGk3LAynkBXTjfW5KTe0oBTkRHFWpf2Pcpd+C8hUmspm7Yp+LWZbA
G62fnEu3ErHVJWHztMwsMB58h61//KfLYbbGEaXrg4ji0JCPcWW9A34Y7xld1rB5
O0vGPK10D+BQwgYGi0Cl3Ag+KESZ9RIF1MwgSUvV5uoWyMPZ2E2oPmEsaXoz389k
qeStfqc3sJIneIMQ4nFtFum0sLCYeT19Xfws5nP7M94wg4bvWY8pZHIHK+7s9ZlC
yPitWq+SnA20B1PbMR+5BThNsJKD88r0jh0tzHAb3L/2Ljs35jo+AqYHKybyRT+m
+Sj2vz9Q34o78xtPdVO5yuuQ4EwwK67JpZUc2EwYR3iTAeKv0vxLHciatdAiJxHo
sJA5K0HR56RtmFKntE0teblxlz3llTVtADGHM/sii4jj3EcOo2jdSuPrMQKXW/a/
ky/uTA/SJvS7xrJIL8fm6SWJIrQk1nvJ1s48abuE+q9xD8f+0w+8xggDmS2qJAWi
j4R3/DOIjU5MM6V1i5tFDZRifvTuwCqM0coIEzfFargtrWn2ubIs8i5eSu1zXFXi
5VHhIX5GbuRku801ncQrfgOAoUhIhlQzYhs4o9rQm3r3AdzfPmQ4Q6wqIcTGlTVI
27GtyUyrpuqy0hRmONSwS030pdftG1d+kWFouhWrj8Sk16UEqgxJWu0MNlX+ciS9
u3hvqkvizFzmX3mES4O48gDZNT15YLf2Pv2KEfOjXjSt0CbADvay48XqgDDgdJUc
WqcYPVwzfGISC4MRJcMhPNBuR1LViWwUShdC2mWRjcW23gRdBH9dMSivpH0Ao0RU
I96du7Zglmpk8mOtUrxYQQqyVWVv67knqHKyPgDFK7r8Fb9izvCaAI561UBhJVWB
dVTxj4H83zwAEYD+F3nU9Ly8AMAQTp/hzVVyRLXql8IZmr8AJat9EztpaCovWqqN
88rvNNTv08aSzH4ehgr/1LCPHUbg3d9eqPKUdPKus1K8ZSR7frfHw9a3jHqIziB5
zqfLxWdyXlaHUL3krDI6fNpBVqmDT6MIj2bB9Kvm/rHUtRWtdxj0D1U2L6dnbIEe
MPxzkXKo8xumy7HVsbSWvJcWO2G4pLrbzTvHJxdmq5jx8DD78Lw5Gj8OnPUM/eCe
fdVKkXPAUbSLxzDqrnKws06vSFZRDCiY9F/s6oFiMlaPL7SbRpqxMvCsLYQ18wP4
1to6yimLrew8/MR5F9PgfXStPIEeOcsGDXo3FPBJxSzScCWeM+T4nEvLGvfU2MxF
QzESrFL9vw92COz2xjw/3otifpzTIrawy0H0PtXVAfN2mbWGMFLgOPnN5tCnC8/I
j5JJc7gIaqf3RTqF2CjGSXWPgOu9B94jn7VaHKzO8Ixn93oRECkog5zexKkKiQNJ
zEQ85WLjEqOQUhQNhFV5CnvDIyuPxwcQKi9YYLeRHQzb5fPqZbVafbBtncuodvli
/P8SCYY38WahlpJfbCsC/xMXzZGYL3ak627h+9fOFjhO8R4RUO4GNyOLjZ6rXt5y
tR/J4vMdOCZipQm04Uf4HlpQfIPYdALTO/SA2utvSuoW3VI1U6Oz3Ba5ylC1ZrJE
BzE8W2io84jZz7YefypuxpN59tGan4QqxlBuEwE6eCSTr10u6HGbDJD86zshziVi
fnQGQW29QpCS89fOYOC/LjxOhtIXHVquByyXpEXQRXhNzPtxthXyfYTTvOBEffhJ
4RIixZXdgHXRgA14T0H3Hu6JDQ4THvecm519uvZHUbsYlrWw7ih1h1D5FJ3grk32
hoORZaZ7E5iLS43lukiY+yn6r3G9NCdZepF6/2Jqkbe7W177Tl3+I3kFHq46hkA5
tGdpuUTbIK0AGxAnJ7F7snofG33RF2ByrZ4OPLBd+A6+BB/LygFAcJbeL3jevNtR
RgR6dtjExYb4VE9vPBCCHegzaBggxPF8L4JaB3TavHidGnluGhRlVeE5Snos4NA1
w0OUBM84k2equmDXCJDu84IgdjDWOWvdqizB6bOIY/xHtCdKwuJQzomU10RFjTt1
ZPkXDjooLGz0Ya+tOEArwI70CeV5lJkoLD78kGqlQCleu6jCErcHQZqRuZsBGSi4
bL8PDf2lyWSEpZHNdvT8iirORSgSGsAjabfQp3yku5HbtIOEZBqha/HiT+Mpo2rM
AyEDvt0BpooqoT1LF/28ISskHpDTU8WlYOUadz5ArmrVCP9PJSP6NZexJqWMUb05
SmmcbCEFzVeoWlzJdzUwS+AFskeKVFGxqFNlyEDroMAkdPV9TpdzfpQxdzlYapEi
mXXePD+wjgfnwxS0/VNnHCjSZgL16Mpyd+hU+rtW7vPJUktCwhP+ghYtfddPCiuT
MDF5qoUwRR4SNP3qqHvy2GIvd0uRDFXBgtfsNdEOLv4YAefJYgPswr5kgFPi2IPT
mq7QSR9yCo1U3SL+MDNCcH2+3hsALtYjuj/b9uhu3jvk9rSk5RpTLf/cEOyl9lCm
BPULuyKrsKbFJszEFueWKyg6xDuqqavS67Nl4/MwlWn+IGkbI/mKMshPYGfH2FXy
dolqdLh8KImL6ouJEcL4Mip7m8utdoIGP96cAQ5jaoyxKR8nc39JRYKLUwSHeMip
e1CXIXmoxTeh9qO0hVPNNNBWVH9B2NwBMo/K5tuux03lNYn3L90274sLyvearH/w
j9yanrz00DS/jrapDTJ8Qc7hHchmhSOMZIsIYp0SgOBanTWQxgx+SVCh9AeK8H5X
vXH9YEdw+wp9sq2OfEpVP3Ok1j3dR6naonoedPYx4oyZntI9ElLDliQLAvPIszf2
7FswcvPyK+ODn+0JPi9ZvwAHcbYUSQfZqZbgH1YD+5+zzstvF0Vp96eO1yvCc7N1
h9DNKS8AGM16S2wWODAO+iVXPAgb5qlbpdkYyx/Z0bCVx/GEPkP77Eb8zVUiCxeg
tgTzSJJjs2jJgyf5CC6VY+51JFmkWjUxRuDq58VxMTtIg0qv4zGfgAfW+dJdXT5Z
wBr9mMdC6Ihc3Vu4qE+rw40BJQXY4+FSJIdFnw350wV9APPQ70unE8N4DFwkjAZ7
2yND4JBOmn33YSAjToI+6zYU5qhbxCup9as37PJp9LgeTUdBGZ7S6OTXuIudCpXN
ZMLZMNjWbxLQN6sCYoAFcXBxQrDX9FtpM420Sye32lM10/RBl9914r0CjyF64lsK
w/2/IFf/8Z33djhT7vlXAeGCjOqOXbzxTikw9TuvQKLpgmSrpmeF8RmwRvz95lRb
Xs1FrydO3y6EFeK3tNxBbGXRSDK97BO6D7fOTE9XG3YXwyd2DT6AEJK2kAbonxYg
5d2G7ztZrtHwPckS3QJUlGescRAA9ELBxJeo/H8oj9oYWY7x6a854EKj8HngwdbS
iGQQAyJ9fIpRCYT4OGlzxcmCz7H4Kb6Ns9gmoY7tSClgExyIGieIpWv9mt0Pa0xL
HjPfYVsIgcsxbx2tfeLPHMVMbXDL7eY1jmhlok5Ga6ytYv2F3NEYinvKLQNM5T+L
pErPAJZFrsKQkRXn/glr5KHWmiqHYrj+3XmQzg4p9R+lb/+raA7FGAG57qwOyZLq
0ki64vqowMZJk7POLgeFv++iNT5ERDMvVEePSwDWbaW8S7EFQakwfuLH/a3D1XwE
ktDA2NddJkwj5skhsS3EeAAkaJ87UuyT+FjrGAzdv6CPIUFdS5NsBB69GeQ6ZAll
eruGyb7Rp2qnUD6JRz+57fNeJkS+mQupghGzU3rUADbGIozZ/VqaU9vepfTYVtXZ
d4KPeC3EFgHnCZak+tz51VKNkdKTyL6CSX1PddXaSt/BC40DcxE14tpv5RTiebhc
fQw3VWz4DWd2sq9mZKJ0/nN/w87MQt0xzDhbdbe6uCpaFjIlBUxlolalEVUf+z9+
vdf3/6yXeA0VsUnxzBggf5KBZziNz0A1ZQMfKweMi7ZLKAeqaCiyLC4przhGPRET
5GcKce5xKiCkchVap//pJUP6LawkNJ59ngrprauaDqOvsIv58n+gLP2jXF3ctHSf
/i+ecG8cXgpg995dTkLUiG0wTY7eyDmi6bTyu7ucE8BYTn0Dok00PuLFScAFO201
GxEcPhNsC1lVkPirK0IshnMt1x0ywQw3dY8GQL0wb2qWb3Ge6SGTMJOkmGz1GQcZ
QSvBhiWZ1YuvXN5ioYlxhn0xBPdVYyixbExqYteOq+yZ1LzRwV2jUc3gwN7NLQio
30kOj7Jo6+JnUJmRieeQHMLP4C+y7ysPwTCbdR0C/ORxZ2h2Dx8ODxhMimkLdgru
SwFXZOXIeEph+EeFjhj0gZpmbW3SrgpPvuTd7yF387V6JyxW34mGpOhhxDcTB8HU
e8qrH7meLn54AM6AyUl1r6hT1eOTR2aTTTq8BBC50kDYmePq0mQVIqlQJ6bOHhIH
LkBcuQoxzlYxab5aoCoC/F+uRUIlTwaRsdZzrowWCLxdX8wEhJ+PR2QK1LRYx7ee
tSgUmZi7KwjltpVdSNlXkoKFlT4xQK9NWAaKHMPDaR2SkAIvrSHtZavGyz3BmNMc
ULMsOZ1FhQErqyNzptCYSEbQB2yaXmxTXruLSkHcJ8GY0E5T7480TVILQQHF2dbA
iURamR8FX79kzVrTEHGI5ViNkGVlMEQPrjvNtPfa8XHOi+ZXdHDnZlOT5CoaEKbC
QFyQm8Dh8TRI6DOxhvkyHeU1JGvpZewGikFfC2VBfd7/k8DIrENi5mOc42d0Pixk
e0Mlh6t972snApn4PuVDOS2OMI5EQ+FTZk+yQ2LQDDa1fQfAn2cU79WzQOLiu10N
Zvf+v0W6oBW5za5Wp8/ti/VIlQH+k5zA+68Jbb0CJyph0FqCKyFezNAvobkAGFH4
f6cRgDfghpxpw3vNSp+k3ehqyTDaDRLlblFtLqGJIHKWJvbMmzYSWbPg/VOxKKi2
wQKsZCOlijIxBz6byOOkcaRnnNLAlCAIIUBkBVn2PZWvWB7Pb/SjcPKll6wcl8xz
gtaHcjKnNdLnhpyxN33NdDgeq1vSdKzEEMwsJwuEIv9ppDe8ECxFL6Z8g3AdjvsL
4mAevTvOTKWyevxH68DSewCVxLbeQNKs5qqzoIca7IDb1iTV5mnI99B+Dm1FbAb0
i4gBNkH0RFJvupj4OQKelLVaixoKzHfYkUZqDrj1hh0BVYz9EmCEu+vnj4DKnzOD
rz3KeFDkRh3/w17f9+I8bEYUjcymgz6a53HVixl4gyqpmrkzi2tuPv9US/C92nVg
nZ1V+3sG4bWK2XQVW4yLtcrz3iUFuFbshCvYrUyxbQUOs0GrCICDjcUOFflxx+Su
l50iGEgqB861AX6FlWCSO4ggQghZ75lyXmAIPt2acRqaUPqpuBO5TbZknuj/r4X+
SXj+B9+CWlN7A3/KM8a1vqTiRPeDZIpLNoanY/YEb5aA0JF7tXkYAtIZkueY4lkJ
hbDT06oRxCKhc5U2N7u4zkB+Im3wDXREGG2AwrSkMYfaC3olk7svVmGZsLewdRYc
gZ27YBG1FTHnUbOfMlv2KBRJnqOHNfcPc0FQQvMGh8iwFwVLeulvG6ZJUw+LR1y3
LD4FjGMlxRsxVup43H8fQRVHoA90OpJqeqraLCjYnTy6pgEaQYG5BW9AfvUfrchA
rWq03tMS7Hp1thbPVyf8mins+4Z2KAk2pNBk6VJi8/xqGKS/e4f3qR6p7Eglalx+
mPDlAUsQ1+uh7up5f6WFIta2rJvgGe2HoGbVsenAosPS9olNdeWqiYYipBLFeyjS
UleeDEhBJpfJ+rCMavpwcn9td+avVfJPbpqW7hJAXTxprIL1hrugja0d5bX1/DOX
FLesxBD8+Q6++fuVD+vmWSxm/yUVha6qJh7YmILopX/uofrMqLaLkcDcYaLhSUrj
XzxrkJby34J61sPJCUBFK5odcam973QyDf1zGg7f0JaU86XoW5EfSWnOr4t2X0WT
TA8BbuN2KyDjoEeIWff98PC0KS2+PwX2Unks9ZHXK+xoYgH5twUz8P0u6YMlUcim
j4x+qLS6swdpv0FjtngOm/7zS3agnW0+aDMQplfE7l9tllj8uXLzsnfzECXiUlPl
U7cD8m3ecz4MUDKecV6vk+WWJ7EYkP3lGjGt9mf8eWR18AyjI2NvwuqpcmYRZlWw
aKuHvZatrPAldbnQXCdIdY3ff2NhbpTZBBv9kH546hgz23q8IFFHyp9/oUfCnmBS
mWGG7ZFXd+1JReGl5QzcfFjmoaSGNG7+xEkiHDiGWIG6hMYd1l8QqXH++DbmDL/f
7oA3WebjAqMBj5aua8CcDJfeU7hwc6MqqOeiKT5odnApmA56CbFBUbGU4s2aqfxz
DhoaS74IBlQu9P53bc9LLHcvIzN3pSSCXN2rVVfQxMhKJntN2OvcghMjnle4AHfB
w8XKjqnXvcFTs2ML170bNtBGME1SonBDLTO5DFXCzEp+TJacVHpJVZDSTecxDUR4
4x2a90nK2E6UlxnYkKiqvo7eNFmiCtgDsT2TWUeFGPsQcrzXPIL+KbNgmI1Xzk2j
EGJ3JQqhSH/urSwnajl4OqfHlfrvtXj6pdPsuIByy+q1TI5eJEwAWyKqH4Ka/QhQ
ZOU6A4Voh+uFDnfphEP5QqXnuVFxfxTzR4J/aLxU1IfrUy5Z9XzzudDEKYFklgDN
t2tNB8r9CR48qIqJ14xIj0XXgoap3iYYAQNnJHwDstrkbgHCFFm3qsvuM8IActnm
JJRYV801EY4x0AYe54nWsq1umyrIv77W04Ok/LIAdqwhWN+d9yP1+I5L2GX+Bmbw
OFDf/jR2rw/sAIWAgq7pFvxJtrlHzXPq4hgzc5DRwnbSR/nDTaKsgJmrp0lZlBsL
zVyTxHedlv6aOA+N8D+h5MNkQLBuH+BByGhpYYM6oZNyvi0rlxi0E488VHcCq5j8
LPJqIcAIMOOXG05i+dV+N/Lf1qYA9L5szujWhWLVuBYLyO+6hRBLzXf9X2q+kA9R
ZEBuG6uZzqYMK2wXdO/9KNHNrDr3Q60rfNgJARTzCPmIl3zlDRbwG/UJNgix2I+p
BrH3ppK+9t/MwqfcgUz8W2tEaV4KbatMu+OntTW3XuQlHmT8MDEq7arNVq6xL33A
9Fa7t2RIlVnJkbE4wloO478TFRMjgKr7nh5stlb+dggM6G7LXTzRz9qTIRB/pxvH
shNfigzgErYd2ayug7crosfc0JrSyDt5e4eGb3fK3Msx8MogXhFmc90kk6DJuexf
jsqnspSlQ4nbPQKB1HSnX/HlmU0TAfpxAlJ44u+5JlpdemZR5NqKl2Lv1QqdTith
XFPl015utGCfGHctl239PFLBinIUsPe0oaru+RCkMtdKuWFzOMxbkHdI7ZXsNXK8
692bZmp+m5A9KLAvUbjcrSc1sc58WXptsBZ1QIr6VXMJOFTCdBJFOmuyKTmbHklH
RUFsC0kxemUvfnvIbzmVX+SQeEUN03l5uu31PnSWDH+8CaoVhkHG/e/czYMHXSRw
/xyFPBr6nl7FB94FI4NPPlZDDQPQAHFt8ZPi0f/u11RNT+N62l51krbT/+/wozjW
M8O6dN2NKmWoR1L/W3SpNhSUcW3RlA74Emb7fABHCcO2ZmYRV4PkY+lGbubkQ8Rf
m9QDinQPB97cJ6Pedlu37OBlMvpqb3h9/dNx7ke5fcP8meaKcWAQrWayiLNuX+sX
FxpDwIXuaVQ3vVvkM8dl7xAuSX/RCPwgGxl1A09npiklxIaKv1LELY3zMYgsjQ2/
FefwPZ/lKuRwYoncE9uoNseEoOG4A3H+n9nC35etGuQt9T16TiH+uF31sJsrQG/+
91qM35TdZPfw0CAoSagHoidY+U/lLINds9U2ymuog8Q/NjTsgxNO6/gFRdAHSlE9
rTRrfrIP/rAfrPMUUnxnIGq532Sc8Ki4SB+ATv1/Tc1nuxz9goirFALQefBRPcm2
jkCWg+kmE9FWdWAB8TwQQ8OH34XAr8nL9mcLTsuC177nP6EW75ttJebnVDqPeoX4
t2ChTF9AWaSCIOEoK951P6zM00/hyyBQqqTdYDhgPH/2VDs+klBDgm2r5O+LcVPG
VBOX4dLm9ppxM4rPqx/UN+NdCIYhJ8Y6vjlckn7rqcGGaJr7sMjefzORqBR3+/DJ
Hvsn6hrELU8RRS4ZwHRIx1uYDKJgaIW8HwDqFnj2TFgYfXqcneINFmChlcUgAfKc
EvOo0y0zOK8DipyjxSTljbM3L4Djf+48zi2RrI2P7+8KNHkrd2xcQNf2pwJg5ovk
Bn31xaU3jvuCDfwogXPHrtaL7WSJHRXlqtQIuH9zE70KdB44fGLrOIiSDiZ7wcwj
74jrRnVhYHais6obkeEixdI4N6ifKmUiLvstfuWOqyNRwNVjtyfPPusZZv58ndyx
Vzr58CXSLwYT1R9fmF1/3p8JG/ZIGlaPtXbH52igg4gXgAjTlrDuJWKK0prH57W1
JhZkstYYFf+34vNT0odjZC2pqR5VPrMOpCSqiSkRHNSmIJbuSq/3R5cLwdCpXNQr
DySVdcpyWUUy6L9xtQOnofoGneHN2YCu13ckSKWCMpg8YOWHNKelU/sFOGbOS2C2
0VQ6coK4cJoUeYE5E9eps5z0avI6e3ACH+5YG9xm5+jc/9FAXKMMss1zg4TAffEh
NvHNSCIDSl5soryMRd/i0N42YGjwX8n0RDWkwRN05H7szKpPbmXicvHtEKhNg73t
N18gbtotbsywF2tTBZeKZlBQtGodPyyM+ftBvE+X2zsF4RUSRbxe7HlLVEHa+nJW
IjxHFYmXbuiO/EMKst94LBSJXROKhUZNosk2T7GJaTa79om7DnQrTLpvvlDOJWos
JwQRjbYGAwESnUY8GICs+cdP9oVfKB6doaeCKzVyS68pDlB1t9g5ttR2vyFznzKW
zDKDzBo3X6eEE7iSY2MR63/6nsp6qn+AMU3pPTN/Vuk0SqXXIc0zvg6epE8EEYx/
UMeNiKwNYcYK88TeSGQACGOYflZLEAF8+sBHvb8Xsu03Y7Uvr2fm0vudBz+mgGot
VgQ9BcyNUg0prK3c1V6YM/vgMZAs6/Wi4Q5uJ6h4BEyYiuMAG+/TROm4aNrWttiE
H+0kQxT13+wFA5BJ4m4uphWa66idsJgYY3hcNr23jE/lu2hTgf83l59xVNs5fyDw
DcXHZKATmmNYhvjL9qxAzwdnJKWFizshy62UX52c6AhIK/SdhqcnnY6s73a+xuoJ
H4/U4WSavSEZBSBX7eCXWG/YnDNU4J0wOKlI7vPN1j4MgRfvwvI4oiUY15HSRPFf
fbMwyyITpQXcwzwVm3kR29gdk75r4A2qV33Nu+15rUoyOyR1tXFlhWuJ9C8P59cU
ObVU01bj6uWGmTiPY15UB/FZ9XqjAuhKycLJfx94FfKDfeL1WBy+kAiBmXmpcUtM
NtWqLyIdSnZQaGJ11/jhNHooWnb53IFxGbZgPZKNE4onkfRpuAAdB7f9h2j8pEkZ
EWc6kBkv39HckvRek0T/yEACaIlCQd3fkHWrqZ/boleUd1E2uwR+EM9UBgoYJzSQ
YdoXWiqWA85Np988uzYFIDuXowlKJ5XBlx3ITKx2nSkJZqPn8hFw7oOzHdwwxbKR
g7SJ2SM+AYooBIoeegUDpHbyGGPp1PNc7LLJ6wKgNOam5iSylq04qFt+ZOm+IkYc
ClSpVWyzRcSyy+wy1oq4zapOLCdy6LJapOtrHOZ6RLd/G4KXClELuAFTJJeXGjJj
Q2p6mnJKdki7toAqe+zt7x++Lh9ZgCHgkdDEC+WVOMfwxNB33/k1rMywJVXelMty
yTDzSxS8y6QMdgIxxkY2ZT4iyoHomOTbN9Rw+IDhG05wa+BB6WAXIUzTCQJgss2N
wWiUHl/Ca6q3zzUJlvbfgCGKeiJEasiXlC57FP7f90UGjqxas5/UNvQUbvN2+o/n
r2GXv4Xkb2KJlGpMTUpgYYDUtA+HnBm+qduADtfad7JAydmzjVmLL/7z/tEaXWHv
JW0XQQpaG6MwpLnXM2qr4Hvdfd/WyXRvYOq5hCD/kPTIDv8cIvmvjple7IpCW0UK
bZvBrAdnNyb20bdTpyaUtxzf6r89oJDeIDcGywHzBoplxCDoGOz+gvieniSdB/xh
k3tpBs0jnDiD2VS6CcgFY52DMo63m+Hka5qKw4yauGcDf/8WAy7v8zJNCApmxqY/
Qm1z69pM8ymimuj/Ii0VwTfh9b3PbMWetGtVEQDh2IxAjJoy34tBYTYOV2OeXndf
yO597AFTFto98/W4B9xMctsRjgaUZMdcr5DcKbG+O5qEQMGsMf9AWqg3zOVvMgyA
Q5uS+/MhHZLDpXh/PkjnkKGEm7ejO7zPQL9xkOWVcx92/LGJePoGEHqlVpkvoebp
9FCg6r9ehjqENAA49xnV254oBHryDJ/TXOTFdaHXluIauasDvRLKGkAf4VGzSsmv
jNyg9+H+fADV6GR5yatGQgPJyqlCRjMWR/Ws204yFfYmjYIg5XFKGE4EoCq4dCzv
5nIaMsXSp9avVvZ56SuToLVuKDBBBUwAYm9hJFBOETT/RwxXlRNvIUKu8y+4sgY4
2glyDbSFwv4jXN7iijjCDrjVIgtdi+IEpYsn7I6sTS18d21lk/h8DbmwRSG2pLHO
oNM4+kErheu0U6rEDBBg466nWAJd5INAlGedntbOYkxYVULD4FNl2N8uN69H9cj5
KjkNKoPFhZbMsjPekrCIY8Vjx1/wDsThwSWdzwl5tmu0GM63zoVmG9LCorMlpAZT
DgTjGSG+VkihHWr+xuVFLrr+SNxSqKFNoO6yqkEZ9Jr+h2KSkVXIqJ+Ce1K7arqt
p21CYkdq1lgWLdlusKlI/V/tlap0lVABl66wl/tvHYCx0YAnzcKDfzckIyXcHHYL
4dkRAWyjn97sNdNIPPNF/QCvFdYVkHUMeczTYMnF1q1j8aZQvl/BjqSB/VR659BZ
XRUsFJNoD5nEUQNMSXBFaUpr8mmX7owQZxouDmF5S+jH01suQi+40RBdlcSAjs/F
hGCti2M/xLWdgtX7HfKI4wX7noTm8bgKQmNm29shnNSSTB6YNttCvqXr6kS8NweO
7Grt/HvVyeqT9aO2d0lQHxmuMB1GfrVOyqWDI9vxg/vxk2rCaGWBSfBD+CYf9/aB
AmVmIsw18YKDTkuznzN3V8pCkMSN+56w6LyDcoyC2kuxCWSAUtVAGsGnP2MGRBaM
pctLZ+BNcr2qV52HA1wGCLRUdDmcpRx7f1+p8F1AfkPalNPYSIenw83KbtKateT+
AfFx6FSxdwxI7ZzVVyDiduh/D9ocmGJnFcX6IZj0nqoLRmliSogM64Nkgu6skw2H
DcFeRrJgRytmRzypgvVvfuyyymsd4eqDBrUFzGw5VZzJH4hHS9dNm0Lu97siOODw
1ZoyJi8eF6Z2SFRX7kSl3J3vUDpzM180eATPh07VM07OjN/Hprht1K9Fpld6qLOn
PZSGex8cOCbgNLfywKy1QLynluj3F2uCEZrfG8OY3/bYLdEU+kw/CY1dXUMknHZY
bOMCTNrp/Gu1qMI1dZQoB7CKLWEaQyOIA9hbCRDYpq4/2sr5k6haop6lSFi8rCCZ
EZQf8ZiSW7oCLRGc7zsqvUeua11SNCXofpHFFPV/wt7gVhgHsb0TnrbzPVK0CZg0
bNOy7ml5zbVCbop3Glfahte8DOULYAaeSZ6TW4ECOKwiS9J3Ers30DXa5Apgi/u9
TN5F20E3he7Fk6Lp5EJZq6jeZ+s8tReXoPT1JVjAGol6DE0G+mEz54TPEN5xBjmy
QC6fW0TlrHMMhvOpeZDEkWDhVhdUKXp4JIraXZMF2cyIanZdfhKXDrl8kZcSa+I4
UCUi6Q83BTM9+EUkTsgdaJflQqFwJ0Wu1J5yVV2wsSNfPvu/ewHL/E+V78yfKwfv
pPArEIIcRMl0yNwJ7TP7yMDaJFS4Bk6uGs4eb0uiMET5DVNJvQr/WgYe3tK92Jie
l5AjHRAMch6e1QbQtDdbubItKiZ64RMJ5ipaMz2DkSjxbDouQ/zlwhDc+U5uW7F5
/FL0F4BOQ1adMpxUVGqlNk2aeYLkQxZmLmoVVPI+/OX6thWbiRxD6rSzMTMbZfjc
na4t4+zs4niaA85NJD7U3iY6GwQfvb0zs6h48WmijBwMpG1C3pm72I+6vlVKzs7i
B9+4kQsAmPbdA6Zx8eugZm1P6ADmQABVZuzahYfx1GmNUWUFeCYAtKMshuscToz9
tnGgdndU2OK8t8jO+8I0mG6aCJ3AJ2GnoXXlzH/SSGEgTaJ5/WQ6z+jWcrgFeslT
7SD19DmF5J9jK02F84xvAxx0HpHmFbdmSXCMMLtAyCjZ9fkVG41CXS4qQ7N31eEm
Mf/NivLUgZps8YA6o+edfI0gedm2Ub9gFI+PwPGy4eDxumiNsKJvg4KytqUtm8T2
D2oEr8i2js6lq+9fOnaw3BUafIYNco4IHgs9LS29562pjpTGXodQItWdeG0HjSD8
TbzrGC7cVkRZQj5iclAG2YoTCmGKhJf05Cm3nw30+LSHK7o6OqpSagxUj8skqSO3
nnAyGx9IRlMZkMUgSXancD01CNRIS5IjxxlBHrAoRQPOZgGKsgnj3CitJSUXTOI3
PNt5KfiVLIQu/KbxGIp2yP6XfjZy12/3Nie+2Ub1VDo2J1qTNl66RWdt4VwEk9jz
J3tafS4XPLNId8D6SMlDsLo4q1qn22Nc4du9iJ6RAb4itjTL+ue59GMaGWiiRMTU
R5Fuk5O+cb0Ss3xsLBJlkTcP+QjPvLgR2L3vrUVVQ2DyyUmegdVqH2Z5bOy1ouP7
AlG2fvif2UJtVHPUUFudgN6pFQLs8DtPdD5vDKo9PEq68f1gLdkBefeq/ubkB/hz
dZNXpJbsxqSEcozGZbMnbvbT+D6Dt91CDr5W2h22oUxrW+Zl8u+zQYcfalHgMp7c
vJUSFz4K7/GCjL1CdLB1nCwofr7qhB87+wsAb+Xd3962JBFrxvxw9K3eETSS4fbG
/08uv8wBPTg0CBay0uS8EGxWTJkKWsR0iuYi9/9QObFq3Gb0toTuJjnB0THs0A+d
bUVVw8llSo3mRCc2olWJDl2nkw66xq0iddVcFwTqqVDFXhre+aSSmmkxkG5FWz+Z
f7IDatqAu5IbN7KKYoBVEmHyHwOsx/meR8Oo9ouxj39RefSRMREbi/Vvk3YMYzL4
SsRRaopgXrVq+zOyj9lB2n9v2JONmzN/n+8Gqq9mQtmjp2uWviyZtRPIbPVjNYIY
vv4kg23rnBIQEidoWchx//TaNyUH24dFtp9F54rlTvDX4wXDNCeIf4t0Bq3nA4Ew
X9iaDf/BM6EPLYcf8ShOUZjzRDBMGm5PbcFJmnYo+OFKAIuRiNpacUCKO2BnZsjX
lGn8ux8f9LhoQOWbrPwwfv1ApxgMuVJPKZGlRTA581ZzS6UowUtcu0qZj2dgvZ6s
DKa09rmJkZjCX7vY+exk6rMi3iedrGlahliQHR4e/KuFyADds6G11WB79YUYYRST
w+/N7vHjpro1ruuHn1iNtn27KCYDICpTAebMJQE2ijT2IMQV8KMnC+ToJnXaIpIN
cXx+1NvVRaGskEgJVjUFvo9DC3sbqS+dzcI9d5faAgeGitzduTKNn81QK68rFL4q
5UGtDxwak7BZJgdlCeKBx9qw0XDwu0mlDlh8PRd/gsyenIzc60bATyhLlGGPSvYs
Cme9mr0V2Wvfe/lsacPngjtA3cwUFhTUNsUbl7V3s1ypsBpbgnjFkkL25J/cVnWr
E1wZsO22DSF5KqJdeHRa8aA1FcziTp5l4oLxNiUwYGl0GW0krO9TOZdqDdxMfax0
tX6kBXnkeGOcKDA4EjIs0UdU7MYT3lLMk1vK4ql1jkuXdQ5lW5t45viwJA8r6kns
uVSungn50XrP8PyVwnU62YuoiglGVxnMP9ihEmRzq1qVZ2ix1jFEs/XmRk+9OkT6
2bOWf9+AiKcKxO7+UKUZ2c8I0PLlKm66AZtemPrrEdchQgVIzcUB8bEv6lEXHHQi
MW/g3ImnA7yCVRvgErfj+pz2vDWkmClC1BJyzslBDoisKxItv1pgMxaxXBt3LXXl
HdfkjNePj6rvv0AyvWj+LpR6bvvcu5exQQ9gfV0+hsQUboF3LWFj8dnbtgy/nCI3
YwtHX+SLFVt2R3kem6Uj4cAuSMhZlmZd4WKN/Uz+Eb+BCBmhN0cVbokloqVOo3RQ
1i5eER2v54lr5Vyav6a7Zg5WUgCU7hQ6ackEqjHf1dz0jhYkdq224GLwS1QO4RP9
uAyToDUUKkZNdRp7BXFXLNUl63B7RTWEm2tinTpCSzk3h5eZgAOStxnklsRvLRZk
+jFz4FsDZWC/jeJ/NC565qQir+oJmlmJ13Oxm+0NgrBEpt8X05X1erJsCBcZk+E6
Z/8LBrvoNXY5LkaMHi9XNsfMQyLmvKV9Dw3LfpzgtevQvMZyxPcry3VNwaGYj+HY
vQWyisUeypldDzPU4WbnUslcNOyr5hPI+GHnaGc2Qjzzp5RHMdB96uCPc30mNnq2
WvNjfgW6UfAd1lGhtOCoyn8Nzydlgk8HvOsbNXdT/o55rf1WgyHLnlVQGBOUM+HG
4rmqUZPLy2kgZKXIOHQ52Lz6IiTluslwZCLK5aAXdqSJF4SH+wZfkSZ7vloZo2Ix
W6K2mRCxF4QCdlwMfPbO8pWoG0yfDMM6+RSagqLJISY5kRgX8XDl6U7tWjrW0uB7
+PdQ6/WJQTObTT/BrlgA0mhSYrhD/t+RWaeRjjFhgJOThkjDzO9Zi4d2yQzTd6KS
KmPSQQZ6OWsTCG9Ts0+aYIkRd0zB1m2XjPwqqcwm+VeXAcLYPx6S+Rrm+FPrrApN
iLTSQwQQR4gVlOEYggQY3YjLILv1l913GUv0vrJTrzjmhMsVlFQm7X4ELq3Mst3S
U/grVstLxnoiyZeXRAML2oz40QpzS9wekX4N5UwBBQxlqCe//9u6mT9FvoJuo7Ab
qJLxml/KPs8BzrrSivSO0dafmq9cEALMg7MgBMY+B8v0FjrNWZ6ZHRc0sRHb2YNF
OahYTgghfLFC4u2ang7dGBPFi3Fm+QKzrm8qSLeKW2xrhGCrDLscehTbkKSZ6PUV
QoOz7Hye0BglOqoylBEFnnAyRWRmwn6vw05MLys/SlRClZvxrQHYwAyPnkS9SSwb
L6mvAgYJvrAJocHYnks/5s1KIA/DfBqNyd/eLmsBocNMA8WYFCC+hnDoiJBgcUv1
uOxpskfPn22SNQLRktZGkp56NdEqBBH+3ZyxfsZFkAbAR5kK1JDcuEtvRQ34pyCg
EejO34FwgAYArYGpV8RRC3ammNWVJLtIR6cvp90AmM35/AZIFeN71ubwDHfd9Vwu
YZE5orbPGzfx0h40K+8fca7HkBu/IODcXAd+TqiVWYj36NyESH/xsZcnsxGDnhtF
pbgBP1XJhlWjY47zD/mKK5K/sOAzElyVdRTZ4VL9+d2HrnQCxK+TJ98KFl5uBsPP
EWfpHYDYZtael19UCHSrCyVMELp9e8HyBT3uqTMfw5NDiIvKVUz+HmOdxdd+lbP8
tZqOhQM0/WnXYQEeoNrCaxVaJ7KGar/N8Ri3C4b789fVPgwmusgCcord8i2elo6c
mtdIfWTDME9sZvkyGlzSrPO/h4sSlUZVsUIZzouFUKgW0wSHiMFCku/4bCoQLfML
FmJOODR8xyyYCXQ7PaQAnhBthPzIicXZvhCeBERSar24Mp8naOyAz7oMXKVkiQ7S
7w15czHSlEJFgyVV/iGL8IdBCgtsF1aSuoIu79EJm1eNQ3GK5Aa7mTkPkX71X2Z/
UoZxYAbsnHznrZZbebYV+I3uHt4Zrd+n57aJ8cwGt9llQIKVkiLkAP4HwYG8GMxR
/yu2DzIcK6aP3hNfcEL+cJK2BrQDCqmV0Hd3JLa85gkrfYgVWU3HI8ZRdVeXTeRw
oWLKfjXr8s9nS7pFqC5sTGEarOw4PWo6zGumrm70gkN6z7BEX7mg2p09Xr4eLMHm
TTSxCB4gCdcfCAp1uGmcIp3RiEl6mdrO0vQmizJEEp0a/ViO7iDvp+HRV/oXqlLh
DvhfoEwU8Fy5ynmrYD+fZmXd3wKDEnDuuJZr5kGMCtRvm2E90PILYt4C2ARAHEBk
D3pRAXBqz90HLFkZdyPpQJ+B4+ctESi32GRhG+H2Kykhsm6uOrnUv0IYSdQSwQ+0
oedkI7qdRHIoEVlUQZCENLLqpwv3cSvqIMEDfp0G76yySaPzSHc4QUvTmrXWriu0
R51i/beKRYbHqwc04JbzhDguQVKHlOZZmw13cb32toQnpzsi1fAlfh6xw1/fInX3
mpVQ2PVQ6OGXYcm/qVdIZXW1tWBvmCNsEOB5AAz+sGe//6MO1ZZhtSMo3IXRrnaK
6AW/+NBpUh3FJTIO1bYjPeiuYvNp11f8Q8VhGdeX/s8xHgUyqlWSfWUFfUwhhdiL
LicqvC3DlHE1QaRyGCjRMt7NRNhDlg+lbMcMmgixf67GLpY8RrIFQwM2dQTOTcV+
270oWVNVkJG3XYnsk3O7xWqR6CpXMpyMesqvmtHo2VXTyeD8Mpq1Ffrgmkz4tFzO
DoKNQFac1Ue+zhpN5mBgTpZEAyH6X45V1J2MGYKJ16zJ9NfFqsL6BWueZVYOuGBo
vQqRu75zqptys0p2NMxwBZYNHtGKAPgzuSFN6G59q5Qz/Vr7tqQeLX6+TgLEBWBZ
3y7RwiMm1CQ3EWAs76anKl9fJ7Y2O972D7qZ0J35WeOn6ew3bEmeQcXSUVz247hE
avx27mwH+FCssnpH9Rrgnz7lMrwvERRFOg1LI+hnf+923l0eB2TL40Xx7yPbT5pP
ldpn1Cg7uVyqwvOj32sJ98T5LHSTXc2GXrJDYjnsGfp54Kp+ahQMtuwrOshschaG
JXAKzRdrBRxFnplitE10+AoQWDIWNimmrGRDGrt45hJQNKR+4sG6iISceI/DWzpi
ibXpR/hsKOuonx/W8/d2YxYv9iLb3SWqtmkmm0t5azecf6+8um7RZFz+SKDCqsP5
HC0mA4yPgnY17B68zdS5fWtOWK20gDeXf1j4Akh17b5b8QONmGp1D+ixtJC5ZLaJ
VU4wZcuuYvyFeKirbbJ6Plj/PeeMb5Sf+vW3kHLny5U2nhSLYA8Z8ZTq2Kmp1aIP
EAWHSDv6Tp7GUr6iGOFEdGA63WyLNGKQ8Oom71THMf2PPePEsbw28nWZ3nQATl0D
X31exU6gmMNEUHhRzW0iemigp8xWHsxLihR6TrutO2pPW0AfqEg9B6bHnii8NEgl
U6KJWdaeLdDBsTDzB1ko7GjpPIZJZU+WbdcRLTKHnf/ejvX3sDos9PP2zJFLjjNY
1ZsvrIkaMnyjSZt0yf71Sg85zeSFks5uxgXcYD8wQDBqBdJ5ZVd/Dvwi7wTGG70k
N5mXLUfirkvtKE5d8DaDignn+dxtpeYHF3D6wmVSNbuArsNOnetMN8I6Z26eoXTg
XSZG39nbe/DmGyRKCp07P1KvEgy6stbtgV+Ruk1zy1IDloTJ0UifZDeXj4+G0hvc
G0PCrLZMCJZuwMBzJ3FtjCqyrLOOdgbJYHOF91hrQ+ddeRkTso+Mm6h+/AstK0Xw
EUcGK8K2XJKz69n/qW7MJYsHVBLPt6CzxPPyCRC6hPt8JjZ9b4Yd3NdRrxYwd/8o
H8xWssIEZyuFjmdEUtQAZr6TI4ErgcMnhrbVqPE38FZU+n9yzF299CAoKrIB0eK2
9c0dKfBnYKx87lsUDcWrrndDeNrFSLcnUhBaoKqhxNksINfqmxINOAjNoz7ZbGHk
176Ii6AoH+5WLe684SXBqu7uD+erVSkqmNaSjyO49JyJWYMVx3SNL+2dUZ2hsxhA
jaVds8xVpzZFjiDtOKCMxHq6bstlnyNb7OXQn7bncoRXFg9VcgVZmM35vOrWGMzb
fKD2mJogmJV3uP07hFgPgAYbgW0wh0KJSbf0vIRuTGsEHJ3En2Q/avD018HvEmHe
d5e7wHJc9X6HxCD3NM92cbeYdT4TVNAokGUEcmHyYFFkAdW9YS7dOvDYzTGb/cW3
90hE9BrucORCa5sN8m/V68KZHcfgtXttd2lDF5c4zLbSAdCh/MfOIQZrpPUahbuW
9NWDCSzwr/vv9UBxHCNwsTXMfa/9tKFVuEh+NcBW6uZSCDL0QQDqimzNNUAKcx2Y
QtvmfRPXhNzmoDlW31GULZwG6bTDr4JGX3CLNJuDApG1KeQoPEpLRfZD1prY4FfJ
y8oJ9bjs2WZGzTBmfl0T8lMsD+t9Fq1/6UvS0kbW7AuGd5pBrkT5Pjc6ZnVbGCJs
yC5ujfqs/0PvI63qERVrocEK/j6eHa4VoO6Q7xfaw3VMmsn8buB/T68zWZAaYv3o
1pChVyOgnc8UIymaEySOING9Jftd4rj12yPYVIfA2RujCZ1j3uHqTwQdD9qvTsTE
Bxh2y44Mrih4Aa89L/R2naHO3/RfJbhy91c44s4lxfP29uIXaJTfNpsI9nR5QCGX
1rbKe8A7oroebD0RsHAcw6Ubdyp82zLlXe+/C3UUnsjxZ01a2tMZSpqhgQ9gA5BL
sRu0ZaQjLQy16K+JED/5fyAkQtKwk9JQ4SG/OpbvKqNKxwy38SkOSp+j4/ddGGN0
auPtufZGZKCH8QGdDnVMHM50y9MyrhRln+QahD8e8wkz2DpoIAp6xD6wnfNUkYwu
Iurhl7rWVURO7dsa20eSDf78PpF2QVsQuuRy2l1Dk+MEO4EDotsVcYDTPazCHUYD
He+2vgNa/eQgBYipfV3MfwW/FoV8fiRlSmU1E4ft1Kl+JZeNvRu2j6I8sHTkNWre
mpM0/epKcXhmiB74c4Byx+zZxToQEpstaZ1CYAaBjvCjl3Mk0GevDMuMDv+RiNjj
bptAE1+TaBk5+MvhVa210f9+XqMX+dMtFYYT2/Ox2E7hnGhV+YlSe7Px5MRPhIwa
tiBs06JiCROlJpCx6GkMh11HzLeRoUSuHr7hilBiSmlyPH+ZKmaiA+PC+8uCXVgj
i8HaEEBjgRUjAdETMlK32Us2JGFtdYsK8Sbgqp3ijPE3Hnv5dZD38E3nJ7DwrQll
XKo1Z3pq1Mn6yf7nbpbcPYdEY13/OvpBJBjpunFdYQ7ycoQlznpX0VPPlJVb1OCg
WIUe4R7bNTOkr8GJbNbFstxW17jQWb8EWf/NcHqCOQWV1xayNAmAWaLhUIFmeehv
+4hKYpSjaYRNidx6X/gX6b4kmc9NaLuxDCxFF4N+JeGCqvlWlva0yOUWRM5+8+Gb
xtpwTRszIfv41MtNtH+15m1xGgZXJuUH9T40B8M+bIReSSxhrlvNK+GR3u3zu/sR
6FNqwvgJ6oEDY5WPiMPxSYBQpoJ0qSX3QpsBFPXMNBKTdtDikACukcqf88yD+isi
MLLjXBJR/L2nuNrDD1iYceUVnr1puMrcnD0h0KOzNujxm55ourW3uSbt8h1LQZPy
SeyBNkd0szcHdyGgEhr1RgbCAhWDHC0D6vRU5OIi/w8yZifqZl6F+S2YwNUrxiHJ
V6gDKV8zZpfDxZa+qdVBrTBNTxGRfEazyeneLKD2zqLxrWDOTq7z7qMcZ4iWfyxO
AorFvh1llh2nDWu/jSPklm9YHC33nskT6Tos2BDrEqKQSkhVCKgB+OwcLE3HThNB
yEsNnRE00o8J6bT7AABInwVcDDNxYjLdBm4IXkWC6aMaT0xNcZ46NnczYirhvFOS
gBbT28D4KROaRaNV3wobiaeGooGvSORjFqCFaqx+CxQA7G9WwqT7BcTLLHSSuklw
0V8PKemTLjCSU2HrllmvyFXCQz81QGTuzvT7g4FXLsJa3JNrH8adZ9noA5Rj8wUz
oeSPYYhzpJ9JCUlY5EX59i617WPToeArLPwQ1f9Q3fWYFDz0vKzt+74f3fMUyLol
UdnjvrHExx6emI3EQRCyr+EpQ3llRZua5g9skxs3c6sKEpvJZVk6xzDjHzEOxLjO
j54HHUdaLXrIzntKOykOy9YRTbr/5VXQvIv9/x7Vo6YFlS0+d+B3yvlh/VJ5EkI2
9uvP759AMO4LafoELGPswARWsyJ7loqze74hZzUbpCJ2KgtbYXnsK7I8snkNEr+2
8E3PQ3+AdGN6xqZOYeWxsn81XQmW9s2nqLGDQQA+XWyGBIj0GgaRrGKIF8LT//gz
0QX8q9h1zlgXaFwe2tpvRWuOo5e6eTLoFbI6XEFV3Px/T7NoxrEKDNQoaChS0Emc
jC5AOlux7X0GgwTqoKD/lY3XRiWgA0jHP6avZmbBNlqjmqOEl0zvwc2LUSEh6T76
Yvt+xR/s4pEeuv8Ht4nO8WJWvIahXR/z7Dar2tf/cX8czYy4U3hhrFqzrfjy/M0n
Hjbpa51ALhg9LwAdZlNMnODf+70/XLCsiRXuomzj3mk+kkPbYzQiTQ2gVi16ots+
r0DEnSQbHvodSjwVp8BQIWRorZLss0Y3Lzd0aIkQ21f+QkyfYwQAMzYVd/M490Tc
YjGrsHTeUAWWIR2jsR2aaANoyl4bf4M6mupEvUTTgQxN1VrwS2tmGxvST2O6q/eI
W50CNYyqxjKNGWDycO1ZVV3li76LIc9WdsXjfnYXXzVSMR00WDrda/cEp7XtVCzJ
q8S+f9WEWWHKUugDbPcnqsqb3852S92opTVYDQt76Y7FtbnSvmTjOFa0xdDf/A/Y
D+bwMUusDMbWR1gPHtoNnWs1RLks+FWvht7KbgzekAJ7yvNFjT0KZA5de9Sxzhen
3VlqGHwcCKDZu3yazZazzRojPIiUhnwWZB1bw33pJCAH9ro6oDP4qbj01nmYfSKJ
o7oFlsHIkoBfvwRjVKY/ars5Ya6dF54xwN69o3pxmA7Ew+b82VJHQ3OSL/wc+E0/
CQht0ohw6DuatZfcSYuJ5dmvEFheh7DV3j4CcP0j6mvfoJJRhnht2ytODpPRVCZe
qkJPQLcMPkB8RMYUONgGSjktT7evbH8s7H0qd30khUh/S5Hvd5iu0wJiMSreMKy/
sNGmFemO7Np2HP7FJiZHl2TAXhbUqdePRADrKxIL7B7+jjCWYHGk3Ns1/ft6B3jq
DD/5Ohzud7NdmPZRJzKr09SmIaEhczjNU/PMrMXO2Vm+ExrfTpxxO2hHfSdaRF4x
u24oBq+TUhZbLJyTSUM669vVBCfziQ3l1xRma5gqB7DtVGcCGnikniAIzCt024O6
yyi5zEpE6dpVFoyedcS6occS04DWSdxQQRb6olHzc4qWTsbXQtxhyAc4fAhKFclM
1AMcTH+TrnpoTx8UNO51G5N/dsy3FEbSEPKTta+9PgANFI0hrl5k1Jqit3Y9rQej
FubPyRP8roe9moxofSfMs4IGS7CuKhK6BET5LjyLg9aop/6psgBq7KH6HkzqhhNF
P7fRNzDRK8b90WikiGnjBI42m0rAfp0d0zWJPidCUx0agP/+0dlCASCFjnuJH9qf
VnYkJKX3cwtmLbwxDxcs5q2cQLTbmDl35MDG/H7zWFtzxruD/m0nJ7akYODa3KHm
aILae9geUC9EP4v1sQr5Wy0jb8Lsk+DizotY50xPTOaM3/QeftvRM/ME0MOmy0f3
qSpr9/i3/lLT81VP58qbv/pzOp53Yh2AA9bEULtHvAne/oaT9tl/Qa15Cr/qCC0k
W/AL6IH2xZAmhcTf44d9fTZ8f1QlVnPvejRaviALyRc1d837qgtZFoIIFi0dxtfw
9kVEjwEPjCixSqnyDIBqTt/kiOw6RWXtZxx63TYLJ9r5ZadvROlgWk+F7NrUUdGL
rLzYhr8443FdxvofH9LX3ICCknVmnaIWKzRD7v1HTHvp6N6S+zZcRFLtZAQsrUBZ
Cwa4pJEGhDT+JXXHkSbpW1JB7US6+/Z40d8mx/vhbytkrofsytxThu5BYGJDphMY
Xn47seZgq58EVFgJMxn1iX8bV+eR0cVAmu0wzBZA45QLgZ+yS31jtgPCQa0Ao4Rw
ZaFmBbMJMzZMj9ymY2MR+qaeJNEnmW2IqdG7Wh9bYen0AePVo14b37UzuPVuroaa
Gvtfs3uLGni3fKCHmy6Pr5uVB3sABzAhWKE7tyPneK9GHbWZMCqK5lUS1ODpu+S6
fBuz8kVUEQJEyudGjDiX5LujbYECL/nb+4tOGJLzTyCYjcuqyEV7AR1yQlKbvXCU
zofnfi+Kc72ewOzTEugKGPuaUfTFNiyvD0Cv+nkEmPbqbcxB/rOWdyM67PyRAMIV
ai/FsWoh7mBp+UXzS+UU0vjHzbzthlkfX+4pBS1Pi929iryuGz6xpoUXkxiKq7SW
6sITePaCOn95WFpQSnD3yJ/9bdMuPJDdEIRnDwAlc7pEq9n7GiwHP63bHx/en921
Ep6xR20lMRRfC1z+ZamLNYFqlKU5NIKy9mQwoJDVT7ta2o5FvB6dRcl/nN6JgTeR
uAVGX6xgwUirhgcvsaG/Hl1xcJnPLLJ3KZqKg1u6kqKeXN9h3U/DHNK0y1h3SkfE
kfRVmP+PqXR3i4XnVykbHZixd8Gh3zWg9O5yj+H+oJ0CYl5/boIeronDXnwFmCnd
Hgut8CuXQji+zZde1iATn2O7mKb81GEVA7ih+tDAQ+ULvd8LWR4kQUZBlk6OwXtM
vTKWOKYwp3b9eUUf8SdvQ/xy6pJqS9jUv3fJRiuBlUg3kjfC8POqBZxkUs5gqZn1
lmVpD2Gd8TbS1Asp7D38bZ/D+oM+HwrRaLwMOmUwzhQdZHUTZi9MHgn0wADYL1JQ
POSs3Yz8G56sxrm8ZX2SZWEdLMqHYRVh9nPZTgxi2dWGUqfBRIenccHB0i9o5ZeK
eaPucbQAKQDg9arEr6mLh8oU4n9u0SqVuYKDCbr9FisBNuXn4Rk9Swp8XoX56QWi
Pya99ntzX6jYIU904Ld5lIQQocn9YZSwMvWdd46HKeFdFQSutbMehV8TwD1goLwc
w6LecrhZUt32farK8/q9Z1TIe8SsVmZYU3yhM4IR1biScKphTQqHUArsYhsAYtSa
OXHtCOxnx68I9BHZZdI+gQjumtmQhIblD2BdwtKjlpcdQX9w3AXnI2Cy/aXg7PZ3
wYTS0SyVumxbvaNAlnpFgGlFHC0J04H9pE35bEDzRXEMwDKe8lT6nxP/oE9F84bU
fUyxgYpKxrCmvOHoTxV0lK84HvfYJkDz9M53Xb+HZf+r9pCCLIX3Cz8GDqXqqpCi
i5BGZIOa3k4Gd+p1rmuKPDkFlfIpdCZXc2laYSoO4aJYh9C4xfzpDHc7aDZyaaI5
xTh/pl34G+Hu921x4c4ZDKzp4a9hJcqZwhFrtu2rV+pmfkbX2zb6Nbmqxzt/4sT6
RZX/6juMhCJ1/AifweRELJ1cFBOVzROp0kMjcno/Ifvf75l90poNFTI3/4rrYNcu
ci47xQt+TOadRvsSOoXqYk3XSz/hIyNWIzQJ+WYeM7tRsVCQ+ZR3S4m1QQI8IANK
WiKyc3+jh5heDpO5hDJ5sWkKajjapJnF8F1/UAL6X76isJrCMjdKf5lSPf03FOyf
uOxim/4Bg/OoYXH2ioZt+elpzNC5LilHZLUDOOfdl9S9Wig4HO1ig4qG0fgChs7e
zTQXpWsWXVWK8uQQuvGIGWjuxMgXqz0IadqVhX0qtrneP3QcDfeAaBECCfT63f66
rqcocTvugvvPcnM6HpRJY3uXfzK4aPMKBo9one1C+qtjGzOSLnqqMtiK3lytKib1
0zcaIZo6m0ZaWdCCW3uXHQjQtuvm342vyBd6hw5XJq4w4fyBDBZZ24now93bOAaH
Rr2dYK3AK7vGqRRa0ZZyycAEfY6dhHxysvLOfu2AcDLLsh23/t7UHAcl3v1IAC7k
yhKQKAWHvcSJ/vSAoT85Kw==

`pragma protect end_protected
