// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
F+8OeSl0x30S1rwaK4wEC9Dm52zkfi7ru665U5LWuD0hJ+ock+qtL0lcO13ipRS+
FNOGdjD8E1rg/n2gs8HfXhvgfIGMhxB/WbKGT66ASoGhJuDrP38D3MSt9nYwEwSP
ynPQJz/aXkrClq5XFoIRLluxK6fCR+hGVVSBJKZc9nU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1152 )
`pragma protect data_block
9FNNEcFsXtXoQ4QcdowK0nCGw+wHIefcY9jGJ7etgu+OGA7DDo2OcvS4r/U4b/6a
VtXxlGgBfdSwkhoir9KkQVtlj/jWepkDLEkAXAU/VdyGpnH/7pLy2c5l/u1rH1MU
Qv5TNtZe6eOArD9PaDzU4X8rjK7fWW/JS6dU0PKiR8T/hyjShrL4RphhzIR5Ocef
b6nPshOCaLTJgDAfo+5/CTK06v4CHzEPUHm+ICVs3l1UuNX3FI3pe4Og3ihNmppA
fLLgNwAyOt6b/pngIbTl8XmxM6f9TyBTUnvhXlfqdphvcR+jqVBs53bMVIXTBUqN
/wl56PsCI+TIc+C1YUb0gKdMiZYt8VvsG8+Fud8EwGrfx144bm3baPQmcRIL+s6P
S4M8l9aqXt+BAvRCye16HMMGgBIOXjfsZMeUbJPfI+Uwr7ceQwBEYNUzcztalPSA
myzUEllaanMQ3kE1bSdi7jGmfsraXhV1hP5CJfe/Mln0tHqhf+FfaBnfHL8m+o06
eSbm7PjE6oxKc1VZvUVClXIBvlI9fAclg4JhoVcvSolftcX623Kce0Fysz3/NgAy
gPku9HSRPNOJg7VJBCwofjjV4jjUXVFaDw/2Gggi7vqG04eC4hJnwYeV7+uALZPm
xH8nkbM9P0Wng+eypGNZ/xRqoOuDWxZ6Z2AHRLvU+yA2I71fcnHDG+glTjb+gOEG
ndLCgS7Dx94wBW5TZIeCLt27sHIXcubtbPbuaVHqM2PemQo1S5mguXn9Gxi4XXZF
830CDhjFrJb8PNEZTkSpqu4axibMgmgqmv6tv+w7mZWQGNSm9zp015SYFhW52SBN
1i0fWrDFcyEmQh0lEOn7q4Dy9XKYwYuWHpcI++27+rQ2aI06Oub/HsBx91edHoAC
eGaON+9dC86XzUgNcDifrQuT+4hQ/1Bbauhi25RZju+z957al99xoBhy56aVMFZL
lqjnmHYHvc/CirOHmiGHkcqB7T/aIFiCUEORhMdJ4mklcvKXn0KaRggtJzDZVfkB
2G1kGtko7sVKXm5P98k9lNyYRu8wzgWlnqLN7GPS9UCr//FdLaqLMHIXqCtIN2/F
dUYV7MTaRtciWTzweUms0gH1aJLk42IQh7KFIyJUspB83tNH++9mPjvnLVy/ah3c
u8ZVNVYzWyP4oShYtp/gnDYlQVMiBBijfjzHzh93uCWR1Wd3cRtWdzAHD+/Ckzj6
h+1PHEQH8xuI64PWcitB6w3MmZhXpbEdw54p43SmNghnPVaZm/ny6jNc1rJrseh+
Sz5BvT1j3MWQI0V83D8DMR1t+p+/uPmDpkYd6QXTB557bvDPmJFdgH5e+kwG+UyO
M6K+ZqiHs5+8ByxzqAC8E0KX0EQ0XPV+pfTMafBqJLlXe1whw5rgCPDepqwyTJ9F
cCL6DFz3KN5O9321618KZI801Ypy4wuyknETbLZKERaQ10A9nautqqXWOSXAkdy8
Pi07Yb2reoAqTyy4o65sDLtYgYlW58VfTKtpoj+NWQqnucJHXHoDojE6QYhR1TO+

`pragma protect end_protected
