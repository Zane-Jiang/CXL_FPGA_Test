// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
m22fSlDHjASRpuS8kIhfi71K9A1LVwFwkjM2nG5VoDs23v90axtKrSBr/vAoPmDi
ECLvSHwkalBv5VvijjDsM9IKI0V8mm5Xh0tMoqhl7146niBqTh3qHj9WhIciiRTq
kC5cmvYNlh+zDDtE0VIPGRk0dY4P4xvyDoSbRMcnltH4KSRjjIzKUA==
//pragma protect end_key_block
//pragma protect digest_block
c76Jcsb21kA9sVNIGkn6bgOgQ2o=
//pragma protect end_digest_block
//pragma protect data_block
c2C+FlKv/gviSG+uOCGAonaO5zerWXXD9kydpANyTjoRWWy16Rzx8f9WVv+T4Oam
kgT7BuVTGWU/7Z/yDq8+wFwR/e0zaFA/oY72ff1ssKeeoTxTmL8uf2JNh4JpN7R/
bo9IpctY5A0SEjyqqhc+klRMMTFf28SooH5sVL+vDsZ/duuvtvYq9BWkoj+GyEcu
lq+5ndlXPgprl+Ph3JDTMTmPeA+SlbhAJbtoIFU4wenA76zjd3cbpcpR1+28oXjx
Nk5WbjvgcWJdWBt7ujS5ArFzbKfO+Td9m4T7R+b+GGavCz+x+ADBpbQDZ5wkdy+u
6M1pOoUFihIQc/+K9K7hsPSUkU2VvKAlxCh327vbkcYTAfm/C5uPxg4voenKqnt8
7utqayAjXjvtJ4ayRY9KxPBgPxAXXM+MQ2UhxeVnNKiMydtSh21PqxXhMJP23FN4
xPXWcYjz7U+c9MWOoInYRAsGAqTm+MYWZLnc3WbIfE67Cskm6ZLrSiAH6Pwtcq2r
hBUJvARakxtL2CGicnEfImQHupfol0CfW4FlPGHTa5ufbLyR3Xw7K1HbR2S7rfIH
OiBkYdlDvZhE0XMYsCF+Ue1RnOMNwLleyVH8CCGoPYXrugXkYDQsIYt39KWR6jx7
gF3l55Ki1m4UPtq0hPYhzwL1ihTofYKWHdXPmMGoxzJ/mWs0rhVZlmzWzWG5kFjH
cVzhVrb+l9XxH9qKV8iOznETt5UesgGQ0v3DjIms/7TE5gKVH9DNKesbWuYB/tSk
Q5o7FVELre3vNneskBo/lMkAb/eF4hdM6Q2TBqrQ7ReylBv2XknLDMbyvG0rGx29
p6n85jQrfklubQkwXsk75xWgn5qpH7M0Wgc/aC3s2A7lf6y/FePkh08yGho0DmzR
6ZufjSp1mWJsNTvBNsuhA3M4RJaZwERWVU2FfQ/0Rp5UijBg2D3B401TwdpEUrLV
jM+kiy1cOMn5yKbE0UlHi2HxIiTkOT3DH3mlc9Kk0z0jGXZV4KqsEPsXgIg1ik6C
9uBbx9mLstDuQyEQnusl1HiyptFwlYVr5TV8/1ML4TTvyhPO7OcFWGvXGplCGEK+
hopnIeNHDlzBUmPCOefVBqbUrAvvarsINO9232lQmPPm1DWDj4+umcFxzu+Eqliw
EtnTZi4N4oAQZ1+9OCLOh7eLiNnWAaAgGZ663U60Viy700zHQxc8dHnpQyBWwrXN
s7b0boT2HUtzlBJZtNTwwe0v0mkgjOjtZ7/TpgXjxP7Ahi81gfOz67PuteYID027
Yfb+ndSCQkGnjqyTrxmQq1xhjVSE6kf+2SOjwu6C3b9p+UYdG7aHObj4AFGIqIDT
+/7X3s04D81Npf+BvuqdDGvAaysFOjiuinOsPvO0v9o/P9E6ZsP4U05dssuqp/oc
28VEPu/kFmIlo3brjhAYB90japbKD4XHn2tKj2qi68DHFPBNd8z2fKsCg+MRbLKG
BSf8YTt+8SqQLlJgOHn5wMx192rbdG8peWYjWdfnBAcpbASk5J2k/Mc1Z47RPmQw
sV3meTGBjI+NvY2v0ZscQlkKCjumYJXOEZeXlpl2vFtzh3CoDmLKJSnyDS5U5HbG
kdCjQT+H0dGyghW/8yFOY5jryQhMBLNd9JpW4tAnTudD3xpSECkrRwd79WRhDm25
Cvnuzn7m4+m2VGPu4Je56JOhXlixG2PPh99/aNwLozRvY/r07mepm2aWc8//FFvV
f8rko1RBGIG8zHS51N3YYjtU97jM/2Wy6x+Dl2izcbvFEKQCLtczJbV9IwBNUM/P
kQgupjaDzjTlEmj/KSCUDPXe1phL/iU/fIP719DY3dvaVr8UvN10YY7+5SxJ/4hI
gUdrrG8TfK+nryY/Y5/ZmKv/8WqWOMgqSSJGb9cJLIcIWbrjVHrzhniN3S89eMcu
HaO0/ppMcVwdt2GzmEJ56O9bNaTYv2KsF9ovgSPu9C8+/17HPMfeSWTRxUN/+jY6
YuBx37iaGHY4mch2fH1ODkwc2aKF6kYCxLCQ25/PAzsxPWvIyiOOKVlgyNVCn7tL
WR/2uuY0rnRbaQxoJ1Kf/ZEnlapK4o1pNPm2CB4H5AlZVQ7e/mW9eMPHHjvTdb8M
lfXucx7ST2+TCYyU40DBnpjMPatM6dlTOnLEW81HRFS1RHJMgbZ6+Vhx6xFiBLd1
ZjFlXJAAAUhLGxnfdMvY1982ZCKwerKtd7kuCR7Xyq8POJ6RqYxBq27gso85KjHm
ro07TdduxddB7VcX02YNoMSETI5toCJ6dyMDctgUQPn/UCwBgoK9FV0JYIEoGXdI
jm7CFra6YD8F3YWwG28eoJl2y9WY5yGupYPrNN7GcTUNgIIkuW0AwRFYiQa0ipVf
02KZcgUaUYgjIHJJCzdZA97z6mrhShN5FMF4xfTcndMiiZzGC8l/g4DysBIDWim1
0bfmIJ6lZdF8K8iuRCUCBlXDnHJhxIbcBePn1tnrvngfVbHLWP8dyOpBO6P4Il9v
H60NoiJj+4D6T+9CjuPp8hfAcV7NQ9wjUBh80Ldh6GcMw57CwuzCpmLwKV+/HOI6
lZE8w9zWCl4elGRkysnXgpouRtDcXmfVuRK6yL9imBEx98V3SzckTjCJnSeyNRxq
+5w+IIHmGpoDnii8hqcrJpk8SGlybTFLe2SCoNc+tJE4RNJqn41ygjdtBEp1tac5
EXHteRhhMz/RAtKoR+wQaG0IXaj9TooT26eGNUAyTvqJorG5uem8vBEN+6fBatmk
kvcC/Seso8ZwsqFB4QuZV07WYukuoId4r9gs71s+dBauo6OJKbP1vHIqJCT+Zto8
iFFxgMHu7YSyZ4kdprD5jTZR7icEHMfcbZIsfBC7pwQZzdFn7aEPEpeMiw2HTSSt
TJEWY9JWMWkZJHokhaZKJjkEfwoaP85a4EA+57MiRqdTfyg4W7VCz5fsk2uGbElM
Pdvhyr2TONTts/PLKfd+cXYcl+X0iWjYUMYCgP/heoBBjclvm9cRDH9wbA6IRt8T
VejGCUQ4gqtt+Dj3mdopvX5VCu2LHRg9Z+H5Q29ln5ygTnVe1O9qUD2TzxfrMhCN
b+2ryf8VGRzIAwDkmdIX66SDRgGkED02d9EgzUsmw/3a9KlWFfu5RgG5xyrYU/FN
ocVNrall+OHgR6uZa1fteCOvzqXP9YY6LHa/a0cywPnmId84zm87cpInD0NsOvnV
2eogUW5Ua9I4WZTd38tnlBKS++rkkDdSOMnkP0A/BMQ+byYykoFetRif6HJa+gqM
viJl163Tt3CNiwW4ySHV10u0SHN7fmXsXlxHpU1NQ7eLGvVptao8udRcTqbKADJs
rQF3cbP6QSvWHX2ETTkbck3BRz90Kzd+7aQ47y1tF3YG4olTcnHPswzJsU0o1Smr
RKBTXTSqbnbyIxAZuU5mIyJYGB7VKxqzVrGeW8X3THaRuShr/X3iJxluYXhz99ht
/NI19o7bmUmLS3ybQZWkD4pBTE25dcGIqA/Q/xOQbhLhLuoUhg5VLj916v3AIZ90
w00CI3GlEK9VwcOPTpRTQvkwzY5sK9ZOIc9KfVoV6PPptHX48bci84iz0ZO6XoKF
DVagW/swwFKiZHmFVebddwY2qjeOhsi9PtT++wo2LHIc6l08KAKl8JRjJTQw0RqS
Cy5TuOOLIfOkopbF9rkqnrKyaCyLrIglv5ZCy/kI1IjavTwvrqtbUDbOFVlhSjxT
HGY18vvzv19rPunevE/mfT2rDONek04s4wEg5Oly2kET/+0d+vtkVcx3kRax9hdi
abKLiqnJnGiVf0GFZZfJsUG5+7xm+ssEqpN5CJ4W+qlC1McGkqx0CnIsZo90Ie/z
dICRj2BZDKvlt376nFcNxPeBr8N0oivubOH7yBFmCf/CU01Y+i39GuXd5j+qTogz
kGMuCzMKwwXabhSSD/sEfd6OhMhaprldAojn+vp1e0IwRoecJeoPvd8YjYmT67wD
xLeUN/wTm5E555xJUIfctHTM/cVq7J9sEGCAUc0CdCkxNjenTHXM9KsD6bv3tqmf
fxXfZTg7MVNubksVKQqQkprt6UD9/D1Xpf0Bl3RHicvKoP1qNLQwnJ7kfSK7aENP
TnnjN0IJBwSCW+mcamK9H8nNBBh6ffgQlmAPp/b/iWEvTwXRF7HFD31Luw3xfYEi
3d1+Xpo8qPGTQ/fYjM8/HlfcDW2UsJAcJ2ggBEQxc2BkEn2UArc4ce9PPwjJqmvq
oqXz/IpNvUEYn/rANisOinFBMih9PCIWe5qZjidfeVbx2exgvOpK+2R9x7+EDpdo
GrXO1qylXVFbzReJGWTrF3SxB/gt1ze5JjVeVhLJUc7vY6v4GC1+WP3Fl6peUKrD
62WocAqaOUigFb8Su/kMo/Cap1uHLsMRaaTPGMF+J0o1hUvK0QrNpsZWZSobEvCl
pDESg3UgYRf2MtqaPmISOBn5qiuTxrcS1gr9XZog83GIeHkP/r+J+meIavvs1cFd
ShUM0TQ6vRiWa/gjg6dxjGCchwLkOBI7rf0LOxQyOSwZb5DdT8Xa1LhZLiRf9gQy
/tGXeWywGet8j2nhGu4zcsso2RA3sReG4IJ1PrjIx+LDZuKpe6Vh6AcDl+b45Vfq
ATf2+cM5rA6Yr7AbWcxTrq2M/Mwkge5l3oKDysYZsv2CmNBuGdubDIFu9ID36Sv0
OuBDjPM+h93kn55mmYCDpJ5Gz2dm54zjRgCQ21uZFnA4y146isl7uvHDMBY8kqre
BC4NYlWXfjgWJkdr+3s7BA0tc6Xsi5oQjlhJQ188jYYlpM2zCRnw+4P5MF9StiaN
JmiGzBLMLQv/847r6OgQwBEY/x/hmnWq95jSvnmxmwsw6JaXXWmojYV6eeqJbrp9
rfIGBnGwiWBlx7SSv8EuJJn29+JO0Ka0Tq87JETUEdsLjUe8Yalet6zKnNmm8ZSR
t10Gezd5a+MGcjlgh+EiIGXguka4P4ox2MJdK32jXyTq0Ei/4AWC13MYU0tYdfAI
bQ6CqS67Imq+90FIqThS/wqvX//kk0dlfdjCNqv5wZvgDfzy1I6pT1HkCsF4nmhE
UzElhn+hSOSuWTP1lTmRL96OKWq5utr4H2OmYJdJcghHMmCrhygi39I2tH8DaXsk
MfeJ8sRQTULhsKQCF8gJe+pn15Rn8HXNgztmu0iCb8krBIBW1JWrogvsf8arw/pZ
ii5U2/3vnan0x5rgyQzc5wje41cCp8gYkKA6pcZV0F9qTmFul6rSMjGp62SA6j1a
0a3prnyXFr9nX8GGoT6xNUpV8tQRQf/Xv2cq27FKsyCsj3G5HL0+c49Qjj76M3YB
cdJgiUC49eg3LE9/z2dbpyVxtBssaytbrvxmNOUUFqztQXoPGoL2JkciE0cH4vYD
iwMadzJOS1EUutinkvCepPgKlwvmhDPgpl2oT9xOIWl/o9jHo2fHas04p98Lc+UK
r4IDwh85PVbtrpb0bfFG2nidBIw8qKNvSyR62L2J0nh5EEnnNZJcR13a7VVExG4O
bhCt4Rah9l1a7CXvvNw0k0CEu7brkOPjf2fLhIBPUt3madxf4S9DVaOrndZJ78tM
wLYC9O2qmg6oueGxU1E80oJb252S5N00udgrw7R+1Y8ROAfR91KHNvQ1xLCHzlgD
Ur/7Q6hX8Zq6gba5MCfaeYEaIfjpae2mjPYBYseYTk2OlD1EjvZhIxIXMDU+gtSn
6QySELLjF+m+LlPu7NBYTQ==
//pragma protect end_data_block
//pragma protect digest_block
5d01er7AMo0c5Ou1KMGvYBqE07g=
//pragma protect end_digest_block
//pragma protect end_protected
