// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
FCuk3CWsy15buTNlgfbkofCwHzFo0goPlcZFu+r4cp7qtqZpw1qjJS4kJGAGAHZzL0OGvo5Wezv4
yw3McxYwfGrMjQxAArFh4mS0a7TkGztyKeV1WaIaX9Qr28KUXzBscAl+G1uOkL4rHkXDmTvfEgsW
CjDZ1OpkbzbWlh6B+eM4V8VXYlBxD0nlWl+TXV9NsxAVdkzu1/gkKuij9vZ2NNt8R2TMrNE2MUCF
Lm9s+xtHwyNSs3Yk/O8SfM/kyijrNJRqGdbBeLNVhmJEyzCjT+ULOC56su1s652ch9G4dzTcCVr5
mhpstnDLG7ObfwG5Ua+cpDHYV8hAfc7K1urYBg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14832)
6ohYqge12nizelkFa8iyjD3dxvETFfTcVSWTek71MTB4cjyZ2VNp9ehDcicXR8U7VREstkzcynaY
YC+h2WZH4H76/cxBLVg0T+8pkK+EyCUrL8rjgJWK/8y+MD0mwT9L/riG8luHgj8z7DAwPsxUmxCb
MkVkI2w5jioUB9phY1KuKvRHP1u9nURojg1NbJCpYUsA6I5g4CBy/IaEtGMxHq3foU0sGaSRY0S0
TBrnOGG1g9dY81+zAvNzxW9o/rHl5oeqNhYPZq3pPoxyD1CRTOhFx0TbTOfTiNbidgha2r2BzzWN
NUlgNVaPFFn9naWwFpmX0kLYYdqxjtpZvjnyrI2CMVDXEfsEijaKDaGqMttZKoU2IFvSSPcTd/H9
eEfDgw4voLUAr7cfBX5N6tMySnD1tgErJHq+/O+oOKQcPKjXUTtyFAVWcxdNBThhoIEXmxNNzrmJ
ugfDD++ODQ1dR4upRNHyQXykWCYQEqtSTt17LkKgSak/1hO4YJi3taQkaRbKLsl3RQavWhdKokeS
r5zU4rv4Ibp5GS+7mAOMd7fzdCpANqUZxsqUS4ylXF97DBQOXJtfcJ6aumOPh0cgI/afU39j8T53
gFPm6dUCVf0rkOchV5a2aCMFqIPL4YL5p1fYNsjuZhjl5BiADpEy6W/ja+LKpVQc3GCzPEIeIq9S
2uESMh30vV/NkTzqQ5e7dwH1/Y/2V5SF4dSA6E3FSCQUm1dddtO6ocDAa4AoEN5KCDz1Ds6H25hD
4vsRH0WTKAUdFPQgRP7/tRkCU2UhUnSYX4vQqNw5jxfMg7P4pJ8BFeqgTYUuIQ9z53unPwxgflaq
EqZZPYj0Q9hLPWMhLrDT8wdkscy16wQR8/iBtXbSq52VXs9vYSccJql8GpgjZeqPOdgHmPwr+c0h
3isNKq8im2nMTEq0uk/c1fCKxYlQJnLGjiVMyRrnY22v0oAYPr2eXsFUXUzyk1ReZkYF2fdOBmzy
/uNquZ65xjaUH/mxuGkFaNk9CCyNbSfO5TuCF7gEqlT4m1upbfaaLF3jHd3O9+8oOr/HO468TWl4
akkJ7yO+yd65WrU05LUnI3HkFGF0Z/IEYJzQCfVEUXy+XWh2/3p7zbEQRrfx13i0uKR1krRaxiz0
WXfhyntYMYR/LXO6BDNyBZYVz9YrlcnaOjV5PpPebr/+GYU+CIw7U4KFvwSTyVxi/WVfIYtaLEpe
rhk7Wk4sWx4+YZDMEStllc6kKxs1yrgP4lCEbENsF9D97zXzkAz/qeCHHyjwQWGEkOJQE+oHim99
ww2+wUQa4gpKNKle2mK3+2iuM0FV0Llrt0hdUndTwpLeWbqyHIWabStFiUlWRVOIItWOcnruVQjz
gY3bykUtR+FFpScvxeOaGxABGWA5+gxYKXWEcKP348KTCSBqjJjhIf015gB3iLUFb3Gxg+elYJP7
4EnNP4DCOPTkrV9FWnDCjCfGAdzeyW74znHgAimkrPtRJ40z1yExpTXCU2uSTwRwY4KXM71LuEMs
UOJHyn19hhU0cqr1C4bcreK3dQMguJSokeTRMl9wXzniwTCj3DnLZ//3qRCRmrMcyb6souyMSpC/
FjmCzrW4HGMSr7EMq6fem1fhQeLO7UqdY1557lAOJS6MMWLfxCFT9AQVBR0+62DI0DbEOWrhyURQ
jPPh0rTN3+rw+9Bmn03tGHcELlbG3sWWwDabMQUxo4sXX+sJ48n00+F28FIxzL1VgH5Dfodlmg6a
fTNsZ55wCYA2b1eP0yMpnA1ywIBm91l5D0kEDgFaOgaEVxmstSi1NcDzwQgT89GKGEPbKhECm78h
Vqz4/QPgLBTLf5HPLBArsjZhGMunfkSahJIA3snEKVqKxAK92ovtZLZSShqBF4hr4HdQ/zvsOtxw
vwZ8ocvVk9yxVO+InQ5MpAWEi3ilw5TN80x5k4uAzc0itwQdrJ7Jr/9KEc8qA/SykhwxoJKty0R2
Xp3Smtfv8zlEyAhZ/BOOPoc/1r7F/h2NiRTZc7/rJ9FIs2ZoXURaRrK8XBuEg9Mi4Q1EXDQGf1Lz
0eHUO4l2+fvPOcQTW5GZE7WHYIuYso2Ugt6gGm1jerb2UiQbbrHw3BBFLdkL4g8OOg5lqvg514gj
iRXD/Jfra5lWOprU3tV6s3Gv1/H4aXhVUdxTs7X0TZzTspkNEcusXFAz9fPmJS3h86Qg2ODYkgvs
otKOideJbubzFH8AveWX4mt+mSDz1k5psJOj4drgy3bo0VckgexlY1dfesr7yKFFVEhi505QeNEA
K7Pc7RgDWsonSPbrZ5XfdokikfjUc6ewv28PMsL3ipKQpD3kmhtA/kSlIR0HsNumzm6EKYQSEW4s
0Mmjx1G26JQkC6WJJcUWeFAVa2kSzAp6kPB8w+bDPk7kB4xsH52dWCUB/n6fahke2V8kaoCu93C+
dN1+tIds/+H7lzh8SvSnkOloWZsmprw3UGNrf+BfmMu756iSlfB7G6zTrxyRieebTWcfhzB1Etoa
azqmfJSkO1KwxkifLYu5Y3h5nKtqd+Vpyj8cZYvxC8bbObfXSULgWY1XBBj7DyN0hrhMv+Vjy7Nk
azvMmQHdg7zfkzQBH3H2yhXnjboS3FiC0iJQ+pvvypd5cllDb5rIG8RkDyQwHT5uOpaUoK8p7bLr
VxJU1y2YExsONFNtyFFEDeanmu9vizXKuR5gStVj7skEXbEbhqopnJbrJmqcpg/6DUvu90CwSZf7
Zr9TFxycjkktjdK1wdksv+er89Jj4uqnd/JpXBLUHDkXXC1A5BEDvGb3sbFwtOp1qdVBLYd2qWGj
MJHnuw5dpguh86ZN/p8s6wDO/cwXoDnETEOu2SQ9TC9//Acc7n58wEjyhLgS9Vx99p0TUIbQuc5M
/NG3eRNshGaCCquJtOSqWEhAx60K9dwd0KKzazdU2Bhrdn9/2LsEg3gRifIPKeTpcpkXV+9/baD6
YShq00Oorlhwi3l3qDmT8zEJkwIHiphH7xSz0V/lSceDFrZk4Nxe7y76WX6KFeA2Fwgw6eePo/Zs
IKyyThDVPtyhHGF/1Wq23wG52jO+W4qyplmAD/3K0VnvUL/DhooUGbjBt9c644MTQnAFeP5+ZOoj
U6Hv5f3Wl6VCb0iUCmu0wiiDuD2Zi9lOSELZj91aypnoW79QIjWfcW3+xkqvGMS8/wZS4Vz7dnju
Y6F00Ty2O7y5e6Usc2Ze7vrYQse1AHkg1ZUBVj7AUhPdJWW2KeWMxzBG0YJQ4a8YeF3U5WZ3S6+/
mo31r6Jp+4LHfjlr0VhiVTHBH3DmZ1sgTzd7rjVjtFcrbx3RMD/uDKh3V0DPrgYfJzfjZ3NQnp3s
IRpyVUnppWQy6HK5knHmoi3xGLy35QkvwyAXM2Ee9Z0ReHDj2zj1XPHg8yuBcVu9x85stQi9x/U0
PibwqO2ite1TlOMewSD6XD3GOQn9KQ+V3VPtXjkybHJkzdcWwxW0xJEPLceg5X+3TwjMk26FX0U1
ZtZxVhNxIek09xihVqobUxGmRheMAg8/GvjK8J2+Zco84bdZ+H4T0w9yIRwhewnM6J7FeWjHzUrY
Y2MO/94+ST1nQzk0Gq+C4CzYvp9Ll5A7VrS3vzypSb/LbuJN65UlmuyboWmctXEKFI0DZJZksjkL
xzZuwwpPtn1S67QNcHSl2onkH+d/LpsLe2knpT0TZVL85by31V9weS0ve08HYBs462FKneoebqI8
c+noBsHMXAzHykSz6H6Q1BeMbhwhn2a3d+r9h94DijICS5iuykw2Whrg8VihAZaeh4op7fkcnW2x
og9hehUBc95wq5HyXMOEJzAwNc90fYG4g9cf+kgBK0xfNMfM90UeAJmHzt4VPQfr2HRiQSMMtlDE
vj2dwT1bjVfbt4oy8YMttvkuN9C0gKZSfyE2kzx5S2vX4cJUH1vZo6OA2vYaz/b5IsSn48qwJALl
jHuHOXpjeSgaXJ3JvJoLjj0bWMjZuEEWxasL0/RikC7XJ+pHMgkMAuKvLUF4HUtNA+++R2qkgEhU
b3kLr6GfUYMZjxsuUwJZ17X431mP0sBctDIEDUxr8Gb9icmM9EweI9KQ5J+fCP7WYbHJytUwmHgQ
pPVhERvnS8xMxMu/QNWbwRXYFGUnev7HE/vGhj/HLikqhHy1ffzS2RuTLZ3GZTIqlyfRQEQKKYgB
XIbkXzkvwnOtFmEbqvgQQylTKRmIymWVGTO5ilNDcfVKbU28Amr5QKadd0Dcq2EoIVeOPV1gL1of
LzzORQq9CvL8y7LLI629aFqyeRKV6KQ8SF0U/QasHXD9V0XpbXSYkO816VbgONmFlCydAQnWMYAA
xogiwYwCELhaBUUrpz3v1IF4xV5He5TnjsVl8KAr/yWZF3bc4ewgsw0fybO3MRJI11CwqOma8o3y
wVFZbqvFdFCdpv7jPeFphVV99n3OS04Xq4QRfTsCIA2lVZruhRSCx698pVJyX5sWOXXzTNq3D/+1
D7pjYpBwL7C+LEzuopBsfBkjq6LhXGVUm56SG28mh5Y8pUMNV6WsnIshxZye1lJUdNC8BXokte+R
ldDaJOYAAUCWCvACcnJjzu4ofTTGd1SnfAODyyRulbieituBI61/a4NHyxdCTCjnFDDmJL5eaV5K
Eh0LgDWBXldqKwvKGlqFedcfwMIE5+L+XR8u56SdSalewIq6RkyKSmLnHDDlHphgjo2A6F6TBKW9
+haN8Ro4D7J9bsBidCuz44f3Yv0hyabweSn6bF1mz9zISR98GMLGZ/RqsuQOGJIzYQoXIWpYtk4o
YJhF2JaP9kTIN0wQV6Z1Q1gz+q2dgJMiaLnOS2qOr4HMKrL5QPg6o0/EOOAsDSMiFxSTOE71TA2q
NsX/kUeVdMCXH1W5j9WxDPWdMWddobZMkFsn/hllShKhR8I7FdmCxq1BUhXkJKfB4Jzl7X28or04
2P6xGnNnPsuCpzMtOJ+xnFut7xkCXn7p711IT2R02DcC1PJp++ovltnt8r/w6HpWe05y+6E/EXDO
/sP9Yqk+SFaezcNY+QKIP8pMEhiwXBPvPgJqn5sjKfQRqCzSwOL72spxRnpYyrncR8v+SGMd1AyT
ztPtPLBX82/824FGqDLf/EBnxB0zeKCZuY9KbAM0eqitnj0q6dTBQftjGj+c9GlV0Pnutj506dPi
eUwaTlJVGkNDX1kjS3bg0MI+jf12sBfPuA9Qw174IBVgfTjgkcKUu04yUtbSVKmfgbBTPAW3LN3z
R0DqiuYKulMgxzp4A3EOirSi+8k6jH1LEiixszd2XLJmkdw+msTEpQvIDx/eZ9KGjYzNl2dD7MPm
fzUYPeD9BiYA8YoZsP3fVfUVik4G53id/xeu9yd7Xh0OVDm9Pyl+zOJ8ouTLkFwTsndm4xeybQ4Q
SYD9m+Pk0mLjXX0sMDzYJjIAdypjKKmCHEMfd5DAy9/tL4sjjQ1YVkM8Po9peAZ32zxupT3//Stt
VgdpJgxXT+tbx77NwpFWwClDK4OzyKta43sfm/gd6ZbKWhKSg+lf0NUmUyR50LcQBfKhDhHBDIyP
KDP1DpcIsbx2y82L0wlh5uX/WITm75YXci/99kwgC001JIVk2iC3XVplX+eqTMjHI6yPY5Pa+InG
1lgHSa2fxd9H9A0FiJ0SSl3N017ZrPfZ0Tn7Ooei7fMSj0ndeUsWSz+eXUuVk0L43a1Kx6x5o/Kf
fiI7Dyqw9j9hWhEaJslqUR81yqP4BA4o5Dkvtm6CL9PlpD6DoBrhLIOV78nZg6ix44O0nmakB52c
j2cdiN9MUJxiphb6n89twRznRsp+28MhnJTQzO1aLzzv2air2WwQClD7Rx+xvVxvvYJ3d6Tmz10r
xeBhQfgdPngJxEED5j2cF31M+oyvVSf9P9JUpr+Ns7tZAbLVEqxJFYMmj16wgLYmVs+qqiEn+BV+
Zfwew41nIx49X8oEb2jgJxmILrZGEUEmK43p/ZvbrhuHNkfxgmzlzsewhA9KQsBiKx8sngsb8JJR
PJ2hSP0rfgNIg+SxmQlvQujgn9r9a2tCS4VKv1V+Tl88aaMNtfBtcZzft1KglRHwlkgHL/gSHgu8
OfcMgURy8lG1VlUzo/Ryv42ArS66fwfg4GsZlsvBtIc1aVyc+uJyfYb8vKeEAXO4LzkBpKOWyG4E
3zZL/to3hb7ro7oNdgKgxjWW0k7QMRJaiqKpEscUWjdOEooryV+NpPNf2HkcchnkswwwnugEd2CO
jo6t3YolqW/rEAKU9b3LMEvxFKg0vOGglH1vRayPASSodjU2qnN7T+YELF1MdjlUerBGxv0JUOUq
Rys0HADH82N/LpdkS2DwtVUXJVCwUJIl/ydtWYquPaqiBuqs+ouhhBILLqPJaS4DKhiOfqwisuPZ
IGwhGbBhcZ/OfUyQWwOpaV0CTfcboERGxvuVqSlEKsbZ19bdYso5ClnbC/vdSfNcbSC4ATWJmuCa
i6C2Z+Hu29Orxx3zA9b63nvQd14gLmmE9wv2h5fpgO/7nSxBkN6JgmilBhf7LdOowOrF+7a207/A
6GWamD78h0LaAyXuTwaBkkogA+l9JHW7cg3VdMfJti3qLmqsVA9UwiF/YWKPt7KxPVyEEyGQxudr
HSJI/GI1AuLle0K8qZ1rBhsTvEkl0eMNhsS4/3R3LPQOVPaiTJ+T2akIzfQ3aGxskbNrY7GDzepb
c+gOfA/5lHR6F5WTylrARC9s8dN3Mog/UFaZDzQLkQtyejnBHfk45KACxi+iJFg6SKL8rbuOZSPJ
ksa2GuMcv0Rt8lEYTKPJPMGcESjSYw7DxqyU0+6ps+ZJSfSkgjfGdyvtrkIgeUm4Ml202nIouyCx
sr+Nk6CKqoOjoHXWnDpU0PmwuoP58OzVTMuQHTP0TXkaqxPi7qMdlBbQEZTtfi+NUCMc4vK+fwjb
niaNyGhXt4O98L496e/0Y/DtKY0HgbLdKdXctCmlZpIH+X6T2/DO5WyGAmKHJ3+8Bf3sLcySb+Ke
d6pUKSG9N7/4QZL6NPRYqnrH3n2qBT+qzz+UOJnW4nHw2Z/CBcagKXBO0iUEgvWDHccI8H6JpEBA
/WSSvxhYuVdARcfsNKzSzRBQxat83yGN4DqUwGfiyI3YO27m5wUIYEMzyB7P9h8m/xgJlEJ1H1nQ
YM0/uYp+2eOcpRZfNwa79jRC7mcnJ7829JENWwO6S4CUnsGhc8EjWHhHseKgCtm1jBYkTWXgjn3R
CGs5YVxqYCWqAJHqgojHtGgZy0CjEiqJRR+WYqqk12QOPf+L9zYlsZh/cs99MctldD+cj/HP48j7
ZDZJSRpzlZcnttSGrZ6/PcYDVX3dsVJoz78d7Jt/xao2E/YkxJ1ktI1McQQRkXCc1ThKOaP/WKVM
O902IEvPs4wTOlhIknXvAGg8FuE5DPaXNBjPdhw/NpiKlPrZreDUvWPwKcHyEgld2T0WVFR7BjZs
jcRwmsXneixwm4O5FUFPgV7dkOr9OD6HOVEVC9/hT1PTTGX+f8NeBdWn3xLH3e2COuj/ThdXFifR
036h/6dfba+vnDaHdU1jjYfhGe6ImHlwQoFAS0TqGjXhSnKmrAycu53ZYDO8kE9lc0xKy5Map66V
YcjVopl3O3SEm9tHLeLvUiZZY21MOwr0gNvsOOI9JlGQgGj4FtbZBbRNqdzaJBfQaecxAkt9X+EQ
j5tRDOe5bbE3C5uf7N6KolzFIhC2ZcOuLq0VIEvreaNMlYn0mA7riWsj9oUCzITcY2eTvOb3aQiM
KQYRfn9ip5X9S7Npv82eufSR03RJ/SZdkYMeOhBb/lZDKSEzQwqmB0CowiuIg/qFARnVDnpjjB1Y
16XhwawRPJXHDjAblkOQZgRtvSpJWFS2FJHOAwHLb7O3UnrKqcWebuTUM3q2aANPUk/BxtddSIb/
ucwsj9PgisFHJeHtCxKD1yFmEyumfkUD+ENpAnr82vTJNT7WjR5xV7BEjHJJ/YrycUg1+CIrgNhk
i39vBRQN4r6qewQUha5lsUJknEf+m/dTjBIGYZkWN8Rof2zuxbRvWKR/b7TtcXFhNELuUaKvX5fn
f4IWqpIQQ7HX/rTkgDYMCUbbhbzXpxogUD/ymCm2ZKs2TpO5PJfa1onZNRLNw40GTuz//7wQOa+0
N7HQ04mK4NX6EBIdv6L/syNvQeBG7ygfuoiNICo66P3vFgXBZp7xTi02PcKgsLeAbqdgrMxx+FIY
bijRIxJBI43PRk7SLqMOeuiRxTPa8HThDbwMQuTd2hXqIjwP8rjqWrknndxrU1rhJHUJsKvXyI+P
krfe8ZWLbrqmLvO+3/WJ5iPiJuqIhUN0mNMqK2y16EEWVNCgU2ehVVhjs3pUdpPNzfQCbRdzl79p
MZe9nwuaG3Uf8vMdC920ysyqWNbavTY/NAc8lo9g8TOgJEcMRMyNt14Mk7NYSRzUDoEiD5A0YNhx
mwYmrxrIJJdhana0RXIm9RAs5XjHaR9OX9VbjoxddduO6CIdgwkC57ExIR+Khu4m5MvthhB963rZ
JaVuEIatCJQuGGvKJGnE5MNlMqxKAupsheBtevaOvsUHTNmBkzjHhkvU4pdDBoW0XuUGyHzEkEDC
CXE2wvgGcRReYn4JobHTxaz23NBEFeGGk6Z0XTgzYVrtM0iTItPwbgz7Fs9yGtvVg4LJ+ZRe3kyN
SZURLpc7cKpTsZa/q7aG7XERrsmND8nN/kU9wYz//ng8uKPOWNtxUDbMtPzuEfvnWlgQ9uMbhAeZ
xQkK9irKkKaK7IxEmy3IMTO13EIgHUfbpj/T1NFpO9Eez+l6XPLzJxotqxWta/FWYl0hhjN3HUUX
oaNermoiL7Y8qrOsDVUQ0EvgUKH2tvGvAbmaIZsyiltpir4Y6eYuNRYfie9Wxw0w877+FGE2KzVx
yg7WucfUKXrnpvWgS2Qp/V8HvaL8hG43keEVwbiXw/vwsCKqDyXm2Gq1HQaA7DDmX7LqUDL88hx+
xjUXbaE7VwSnQAzeC+aMzxl+U7Pk7VepYEADQHRaWvovzeWJggiRhQYf/wExrlxGOHZr4zACYoOL
k+E3MQn0Px7YFlqOenV7aV/WUZlaWv1V9gnq7CCWcnsEc5Ykgr/kbwzTnSc/CFLATRUSQsfJCgI2
Ge1X7VeTAvK20OIb4FJe952NRgcWcf3ztQoSRSwhZZExH3gg/9m4qvOhrQPveiTfWVgTjUHc0m9F
+F9LcYuFL9Z2T/Htbq63jh4qEA7JBQCudiKLVrX102WKyGxiUVQhqlSlSjmR6Sr4dAxJDTWqPL5P
+vEjDr7vEw9bmA8Zz4c1ozGD771tcuEKBEUlulzgN09Xzq/ws/quvzsVNMHwv9qh+bv+R98bngPg
MHd5MNvtN//iKkPoYpksTSN2tqC3cVTtuYombMg1M9huxv4pRPrhgSHDEwF3H1Eqq/5s2bY5ORMX
dfp3jCaY9U4knbSUjh26x/hGKesfqLkzqYdypjQlg0BrRTUJEtOe3UI2HEYvDBnn75SCPmN66zqF
JgV3l4qCoE1HnA1KPs3erqATVJoykMvlPZj/LTHNPjRrXgqL2u811qBYR9Qoq6E58dFRlUM72lIP
Gtf5nF6oJ7ew2coDMTZEPZ+GIu9lq3WtNZj4bO4liNsv9BfHIyYqCqFJROcbire2iaN1Ay2GSnrT
kxeSttuDdxkrck6k8x4B+gITFzTQiRx3eeTjznC8Uv1GhaA5XeWMHvyco8n7QtrhA+Yt3mgtYtkJ
5lPY+nt0N5zSN5X5Xow1iv4osmlTU+azY4SfkvpyCiHCMIEyLdQtI1UQKFtf2ofCoE9InqRb1Jvs
4CPHNknYIpnNZV0e3wTx2+ruXmiIrxwPaRd/QoKoOM1f9DGSUKi08zCkq/R8WAF93X5taDvwF2/g
TzNiwbNj3Dyz0JQnCPM7p1Uigcscl+nYTMLKKjeCUhwoHZMW7u6bYtnRVSCUBKcGO/rQx1c/7Qdz
7rXncWTCL+x7Iw3bG9mydNpuiBeXojE4gGhU4qEV76IO/XduDNDxmQfHi12YDlTwOc0NIEzq6ndK
AGytK62B8s9L0NJBr9LMytBMfp5YiIJCXqzdGvVyN4I8vysji4bNMuDjpFanpbbRFc6+BKU+mxR8
kRoIvmbTLtWuPzga0RceR5e3Wd09fqxtTFv5yqjGp0NeFyXFus0B+ue3wUwQgbBG4JHynNpTeYM7
7IMmDAtVUIgnPJV8tTcpqSRSCxc6OWEQ1OSVikxtwNEnRWcnxqyzxtDLl1HT6lVeSaXaT5GmsclT
gvKROMtorLwg9DGv0xStnoPXEdl+KQXoyaOpexgvi7WEaLbTmADBK2Wee7nHkKUmxPW9DpHWjAyP
dWUzmYYN9/YgZ0+Hyugzg+7P2KvcAzNZVmH8MoZRzC9mX7/c4y1emZWuCBqeUKE9h7e3RIQbRWQH
ZaVT2XKX8ChjPG1RsgG2zaWzf/rtD/CxR9AP3LXl5NPYlHnrwW2ooWGet5fMVlDE5sNkU9C45A8M
fBri0wRT+oEeaF+e7SlNHKX9ZF+aS6u+0IvpJGYufbWdTyCBoDKfdiOlolkI2zAsCzdEnEsdmL6S
zuyqeETQhO/2SfClEo9Pp6qZUiXvXHuVSOCLwcKyEEfeWrf/pmQsBK5tMf4wahi/imSWkZDmd/xm
7QRMbB9ywogkYHDONHCY9hbSMAf3Z2L3aL3oogod+OOEvQu+4QOYXgkwRMyyoxR8I1zg8KaSH1HQ
XcvzjRBOsm5AhH6/zWw2p6ZIorsRNXDwCarrrmoeO9nhEFUsLfF33tjPCedzKOCniWWYig3ZPTSN
avN2c1+PZsTWS+aFdlgNUAULcdgEMB50+UBKkry1UmWi+0e74ksu0Uu5lc3h0DbMJR9WruTciLf3
NvfJAM42BwwkpkvoYmE1F8LzfUY2a3maKXVKsIIXC3t3Cu8934E9uTLC6lMm6fGc9LF3mxmva0nf
+DYeprGc8txtl+sLg+Qf1qTe9EBUT10ilU2jjOCuy1gRnn5cotnnCJKSw2l6142rNrUMWqTlQd9n
asGf7ccaPrQmPuIIuITiFqDxQq0F9ysUKW2oAj8eDnShE+wkpUBYhYqt6KLoHoI4L2T7sdsfLFec
CH1CT9Ebu50eueTP43+rH/r+tK3Q/EknLzz9kx8wLTqg9jVS0NPXtOLb4XOLCbpoof5AANuLOcFM
zYubXa4fyrSvZh+aofgXNq5a3Oc//vx0NBkrnCofLcFF8Bct+LXyXoF8fl17HzFFwWo64g4U7sHy
RcSZdHGUP3jnMEDQuwjyStA7W35Q0vCxYVey5pvGwWyJI8QTJ5DaijfvzxFrlnKxoAOFc7DmZASI
PClEeoElCPXK36K1fFSApuCFypSkaMI98EsOD7Yz4tAPOCTAm+USyhdwYcW4Scu97/kEHxXQZKxZ
lVVZU7/LicZvHVrU9wh53E3q4juyN1KPzahCwJ6HYFQaQFJPZTVCnbB4StKcO7CuCLkxt35c1jRJ
2tDzAsJCRJuFiPOyfyUP3XQGyixmKCM+Wk9/Xnd9nyfxtqzhJvYbwLLPENCNoymLBXD/rH5QYbtP
a3mv+2Jm/wPSj9ecCL8kWkeHlsxT05mZ+C7eziHEt/dGBa7kPEjWD9mATfbB3TZhclIt1zgO4XcF
fJXVmF9rOKV2oZTc6mz/CkGXWkiLFr3IFxCkSRI/dtVCZ274IMAlTuuxB9xxZHZm585Lc7UwGOoq
M3kxWGTusVSRJVz224qkfUsaEGbK5QG5G0shqYapWnTmv5+d9rmGOh9H/etmm4/6EIimNIlkb05U
LIXP35YsJP5h6BkEwVRj1Y2uYwTX+OTu8SJFQvZpsCsVb3wYH00VB9ENGi+ZlQ6J2SEqtJT8REB9
s5srhLn2oZlO+ogvjCzqBMX0XbaV+yD1WU9oiESwvYt0IpC6qj40MNIAVOUlpIUpODtqE31EpmEy
Bf1f1y/s396dsVPMUvwV5wganrI44V+UUhGHX3aiDhCfkoPmfy1F3m3MhDc+fZlNn0Kgi+48sKSN
k+SFBkrqk+qlQN4B0kpo5wWMkmPoLPjs1//q9VKWzOaZpn0EcP4onaE5zjR1dWr2HBPh+sFt7nP9
BXyTTdTslz1kG9/LZTlczXB9i5ANPpA9cfljHhbf0+rALY+OfE2eX1KVsIEs2m8+jshaN4UFbLIj
3wnq7zakIi2xX9uPuMe9hjYsJFGnTnIg3DAMa0o1B5oK6Yd/CWJ5q4y0kRB4KqsoOH12FsLNNq/u
hSEJHlJknCUIQrY75Og6jMziQ8zijv22g/fYG+iffqbbb5BpX/JgRoVzSfF3cTnIhdTm624WVMTO
RVqHoR5N1E/dd6Hq4QGXkUZ04rbD9aUC4ZDY57BoUOjXu854ACU54OqV7Aw4u3HNUjMznJP6cvwq
qU/LnJk0T22hKAw2ZCevNHgtCeTyComxblJBZlrVVRIBWUKPBhs2PU9NM2n5MubD6r2I+zU/rkRE
Cii4dEHTxyhB8oPV6Vb3qvlxFWCJ9BE9W8TJlEyV8XAyqM1G79ErBCqDNRm//JabkmHfI22ebm1o
1wyGfGvM+g0CwaBEp1dQippVUk1KfzwJvlpS+KIc1259ZIvnFd5UJQY9jbmEBNGktfM21FhAAsM8
cSRfP7B0YwpFs5Jj6sKVb6dhfF6o+cHk+kAgZkIzwYi/uiwp1WI7RfEceoTcm9EtLH1sb6JHjXDV
qhypTMTfu+pBN/4eai3UrXkW/C5+Mq3kqBnI7aL734s7g18LnhbsNYQBJivaU0KDzXCzXAK8ZDpz
zv5X0xrL88zAm6ydB+3MzinpzQ/QvEKtw7lsNBsiPGxKuuB7FWnwKEI/80hx8xJfkkEWA6bOiCft
zZASBjygGe6gjjwJJiJ+zPvZra1J+2FYYFrwwUfFwqOWMdF5b+KtcuPV7HMLUtraNz4WXn2X55kg
s+ieHw82lntSGbqAQWji5/S/z/VyNKiQpxbJbMcIjnMhxiYNKrg2AiKuyyk1DHXZIZkE9QXIR/RM
bat01Hpqzwxl9vlLRsGUAAQu9kBDRP1H1uzGJO8I7S4nFnI2+R07sEOLD8Up1mP/ibV3BcreIDRv
2mW3aFxggcrh0AGYVdd5FA05BfEyxc5p0z06WsvvEJofN/VivrRKXjvYs2dL1SlnfSDN57GDD7RO
OEJFrMPLe9sz0g9JyEAhojgHhsRH/zX0ioJXR3HgFHsBEbnZdeMUjMx52Ww7uFIKScbV1S+ykhyk
hlsZu8Qm4K8l0XflT/nUMtcJtmHdAuTsrUZyjTQD5IetsD/s7ejBymlbjcGou23mQ+WVeeqEdn8n
2UeX3aeDDWvyEtZ/8sp4tqTIv9AzJOtw2PmPpUZWZ/qIZ7oS+WrDN0Exw9BZjnyCStChSR2m4kwh
4QwcBdag5HcWF6JYBnv9lrINjafwamp2xgGbLd9MbfiPpqrKlP3aRpWOHcb9LL5rKQT/DZUgxVbl
ATW8lYQ/DUwlvXVwCghRWtaAZ2Sfrw/ct0o51rydvdQ3rvsLjC9oCgJZ4ShwGkEuCFn3NuMZnLGx
E30R/dMkMsojS98Go8fUjUAc4goZPPuytcPV6MiPh9mcygxTuGaVLLmTvmlQCZxPGCOTE9eEj29C
XaSIS7VviyCp5sqPI7k4p92tBcFe5D5v4Bwpp9vQH7M2wgQYn2rA1KZsx2BNW7/KqNQcNrsHWkg9
LCMtvK9TQ8UMgvxvxw7wkqeO4El2qP7ShK36uyZTp7zHCRDoWUzNExk7aMP27qJ53rRc+R2qN1ND
fxElWhu7QIE3oE5p0i1H6RxhMg2nxxYa0VahWUrc9kzOwh323KWQz58g7WVBVNL2kJWmgl63QKK3
D7OmaCh0PpIhBKWieFvk9q5gXufrv0+sdOo+juCtB5Zs2c1ff05vZb4bDEKJdDY6dVTn/bsopcxM
PGbFSfjDv/MEiJH+gwCUxTxhDeum7VJXPgtTrFni9sTiho3ga2Gpw+cVu0njQuZLV4KiBH3l0e5o
rjPFaDFjc2d4by83syFXAKTjntoJn0hPLH28mFatLELePWRRz5mP/hhcS06yf68lhvJ1pKilWqsd
nmvEB2+SOe2kyfCkbohbv2RfksWVNqzUSyYuZwxSettVN4Kdz7rVwg+vYmXyKCC1w2SBsW4+JKsM
otCNlWLj4Gz1jBjobW30FNT98jCGqmL/2vlEcnOobGPBL2fUiAOSxsqbd4pribv639mZKCsdMHzF
0eX4j1RrD5nvbCHCsbcW9v4rLv1paEi7k9nPipDiDbXJDMlAzlGKY94EOhpetrD8bOcs30RZeQgR
i2iRzyQzA0RSty5sK9aKQbTNCnTQLoUCpP+jRUagfph3EcXxHeiZj59Y9EaKLJjTb0PrJJtKhmjH
P1CYRQhnDX0dhcfAHx8XoCEGMarYkf7woN0cFDcQCj4k+bZSvetRIoPyvbJf2lMMoOYvpTafOv3B
Q5WqIpS+QP5uipwa+KyPcdXbxO1lG4Eh+oJzjN1WCtPeS0sK3G30QvKjBchr2IgscAKS1QFEQv+w
GiIH9LH4VHON3bPQoFcQ90PTFswJ3SEoG/3memSa3tuZkStzSIsKp+yuDVursE6A5fR4uuE1czAa
D+VsBWTHUeGqs09cAj/6ZpVP5EBCv9jXB367zx/ziGcb+GN+rckGmxfOssxJdJDluqPLcJgwWgy0
jjzm4QL16W9Oy0J8CpYV9q5Srl9+fPqF7AeLECC21ruXB38GwwqJAdXxlQF/iuMrmc9Iegcy1kFW
/32IvEkak7WSJMms2M2oLDHGMh4NtjwpFHj8VpPVm7OYEG1L+B+SuDHRpXEm2fh+xMY6nzRTBjBI
N1JMJMJjPDj/uExrf7eauKsPKRg+CDDxziRybZCLu09q8K94IYMAdncSrhJ6W3lK1xofFL52cU2E
NarOJ30uaRVXZ5A6VEMzLqEKpOp9+7i21+okLfyo3ZsLdQOclTuswZTW3J2lgmfinCPuvXhY2yZW
Qa41Tb5oOcyUQX14ZyT/bnpb31gSocaKU2w+CWNyJMJvZqy0t0XjhmrB3JxDBp1r6wnt+H9HorkA
txywHrPXnrGgzAnntbkl3YT/YxFm2zEsSWwdYvYfmWBzHM8g7XbxtbTDAhlwYIIofCTLlpVj6dXq
N2P2davLAzFKOMlSQTG5ZZLhixaMkf2nCn3pE0bovauOal6jp3/F/LDr1sydk0irU049a14qbXrL
exTK0ckm9qfK+VFj/sLKi1DsR0ixJyduSx8Euv99VKrrZgJEpJNNWuZLkjTVRH1zURiea0pfJORS
vqhF3jCBmvRyTKZ4mg95naqknK9xQgqtn2/VzV4WB8/r5ras2yxP1hdhwKUrZGbZ11DZoqdfo4rp
GhinIVgnnS4KwAyI3WchNkGZKfGcQB3Dv+mqm4Jsv6364tNoI60TNtMs+cloyGBKnvPga8ghQc9N
ZdowolMxnEXd/cyPX50RrI7RKzI29G8e6PP3nGKhBrFeVZgMtwahJ8FlPaSM3uyk4hRQ3/wtJatC
fzKSjRvIrbiiZSNQN/feO6qLcRxGsJNdozPzkB32F6hIkQR3AJCnCbWyX4O98BPiXbQqQGihLQ+q
UvNK2nM8l8Mj9UbzsSys/e19nXgx1qniNACOglLaDUMeeCxanbknqdUvbvjZ9R5db3JAQdGto24Y
SlQGQqWFVy9CRFn9cTquIsSs/qrQVrJ+XEwB/bo55pZ27jYIbvIjmVV+aO5MgOwtI3AUrNwGsx/H
ZyiXxcXsf2eE4+9bsAvIvABLIXJ9vimp79jWrng5D/XPHwHgs8xQzxaADGw8xqPVk5/p/Xajs4vk
oaVQLDuE0vTGjze/zt7ykw5FlkJoxShD5+Fr5T65CzWIYbmo7tHOynymCajnNfVm2maQUzYpFB41
TVbLyDrnJeBwtVPQ52457hCPlNbbBvUGUd2N4Efq9+5oODrVVOIpM0IeYV+O/jDDGotZ436RJFlN
FWw/nOHddbaVoHP1KpNE//8tzFFo1S+JIPSU+7DeA+eMCOMy2rbmgkQs4HZ0bG8xhn2FRqRk5+d5
A/AFyIEA57UnzroE+MTo1rEnnBJhyhZuoBnlWT2EZmxPgHFl66RPH9veY6qmHt+s8MRqISNPaiYb
BCfka//Im8qGaMYfuIlgXacGMPy5fd/SWPPd3rvoBhEQRRlteOPuYgpqFfIyo+iT1yFyW/sWNuiD
qooDPyzKgNFjgCVzkI1H7Td5ECv/KCTsH60MOnCNG6wH2oL9dvI7R7exD96dB91rOnh8CTqDXrF0
32kg3MFpAWNzx1bErnUoDo9M+BoWOYttAKLL35qvMPJA7z7naCG+o2zKZREI7dMgxICzVLbfJMjc
CHJcYEuiyoOg9gatwllCRu/6H191m6LvEt714NBIPmM0zIQj6D5iTJz12ay+pA+V9tR/iByKAv0j
YAIDxjrfdORdm+QpB9pjlPY/53HJ2uQg1UANyAMX5dTMfeLrCH19oOCngyxoSma2dI8wa3Pp3ISt
Z2HmAmUtmrnhN1WZwY1oE9r0Ds+EYvNEmOzru5rWM3ZeDio1mvOaHK8OJeDx5eESJoLFpUV0BhCX
EEa/7F+45qNe1dHrZS0l4FMzmXOnulxX5JCSV3GlYmQD3Pishv3SYjobuOKHU5Pw9acazf/vbM6w
n0bWMSX7OpINGBMfjr3z7amvwPX0GHuzwD/X8thdxyT7S0ZQUb/ISwojAp5mJ7Ggw/3XENw7J6vk
aJnOhxm+VzTEh4WNYT6yAFup9LM2CWIUeqcksxoeK+rvvahEwDDtTVjEf5Wg54IXIj+f/dJe+aW2
Mi5UiqAiZ8fWLalWg2N5rmHYf02lgG3r5Fcj25xZG5hVKf/Etp3j9Q0lpZRF/MsxFxA9j67m2erj
VggaOO/rd2AzdDJU17aYtQlmogD4b1xBM+5rxQAklx5Br/GRxPbKB8xf6cim3NANiRXcamF/XHla
wAFFKGryEek3/E3xAVADq6DC4BY5Gfn01eBGv4PyCyEtlfeTty8t9eORV1/Zl7vJFynjTHuWpynM
Y58MFZX5DBNS2oeLPZXA2REgEu8u89SPOmGwFBi8Kqhfkp4GGMJvw48ePmwuEY4kwMioxYhPj3Ti
KSOyPS14VUKM+qOji/lny1iL8weey6ul3pzECzeeTcmpQlrDe3SzKlhALphaU0Mp3ym5ZQQKGQvg
9gQsgYsJz4md2FRpBlVNHSt8xNbFwiTM5fDxu++kkHGCbEUyUnwJ4BcsJbsjZB/Ddz6USZzj9duz
ZvErtdPBdpgHo15wZWFfqkLe1Tfk3Hktmvz0mWPOoK7jwg3OhYV7pkPmSyA30FzHKQfL+Ka3GbXa
feZ9bJ6EuN+MjcUUubzNzftMct/cAfmkjjG2nWP3bLJbmztrgG3LTonp6VNaDPfYYG1rr8dcVVO5
PubMGeGtpL2J97SleoNYIIn1Cc/hl8Mmm9SY+SaFTW/OMXTMJJbBL0AZdyLrA1JBHRsG58wA7mdI
t6gXUy/bkYYFCi+9qR05k//DS63KFzhc/ph7ajvI7I1B84Tyr2ndyU7WlG5H0OV4QNloWtzvqwo7
fQXDJ6sQKCbscjosNExX7hkGPfPEHZM/YT5uOBlaXSrb6I2ugttX29L7TTxu89UVUtz1sFaFiZRI
AmuNEZIeV3LbnYb4245TKThRfDhXETaAaeVbPmuOrBnmeMf1DekBjVCM2qMPJuNj65d/4qL5/QdM
8eGMwUl37fWEenbcxDShQ0zcbvow7lSiUpEMt5jcXAsQDEsC8FTvL7Yp5Nume/aPUudqtRSF5lUd
o99f49wthcfXfLEH7alB2/OO4D/SuBfB6aDBJ+6EyVZg0tyTG95Je8fAll2RCtDu5YbJIZcTIRop
doJ9yokXefQnoBnyuGAm7+zOf+xk40uJ8McjKqbUFieurf9VP3aXzmhPrBesnBR4GVK+p0Uhb5VQ
2bJrSqK5treN+64Mssy2LVY0+aDv02XGfeWZeYB7ESUSBlVMMyQRSqLi5K9pQPWbAdvft0SPYWkI
6MBub9+9owe/9FBNzq/k7CSr2Nockxt8+/ckvgRTOcBxjvklY5/2GTQSt9yRw9ZQzJKfSQXb9xf8
wyKV8I5zp3dkV3s11W9W+ANLM3lNOpagRKt4BAsBKkYO1ibCcruhjllKgkZukF+lH50gPGG124Az
AX/oz4Xo3PZF5ieRwSASBT4U3E7qgO8QPw5Ga2W6yu+joPBRaVf+mH5tkucDNncMHkHi7f0smgmL
bXRcEUXXKuPRLlh0yLM9xx16WITEMtbSp0P32xx0Tp4PlQzXoIsQyQDDiJj1wVPlHSj+p1ytGGz5
e+3Q9EyCz0dYe2TSWhjkJ/1HpPLY2jLd3eVGMVW/sPoa2PW9HHB9oEbIn/twhU9lMtXMLvSQVZXY
IXCLszZpaWuTs+xxCiIbELW4JRoIAz5hMEyTuAnbsogX16gxBIia4xz39rUbCHMBlcWCrRKVa5Ho
cElfdivjIxRiIb2m4VyYR7CoCnjdnofmynq0/f+/c3fOuFkCBM1I8ESOwyw2uXVeAjO2YkCkt50b
pNJYeqlYiRG6EE8T11c9o97G9tvoW9PXEYEejQftb2BtX9H7JfuECPfOhvZj5TkBIJSYB+YCLdcH
Y+SybLBbHA74g3IIOGfLJw8CpW9j0KR7BA2927fjV5LxZj2ODVdg3NwSq4T8YphZgW6Qcczhax7n
aodf+6YbXS5JvqQeC/VFIhPSwGai+UY8+Tx+TOsoJdVX9W5C1yREO8+4aHJhRfL5kJ+1JCNNFuN3
aKLG4U2qloUEVBjh08Chi1ol2h/0k7p/Tu4u+zsKn18X3NaF8Q4bI56jtyE+tBwbNxAFAra+gy9n
kDOwsm71/FL19lBGWfrNDiKe3SdE66U3BOqY5KhfJ4UVwxUicAEnfOk5KJlxucselI8FdKfTv0ZQ
SuRIb4Vc2s0rYsVs3MDWW9k3vpjoO0eZJPKMwrC/fb62pnLyQRHtYLwgA7ERyE1zVi5thtBJQJi4
iYxwVVBSpEiYAt72nJ7/BKlLecfGRDfUntF3VWM5/ZNBDZuTqS3x1qigYMNZP+EVZltsxHld3vTq
HSmwQ0djLwlV5hc5R8sCesdBytJneVyYFMZLuQyFDOkIvwgtTDWaQEO0lA5/fND6X1dXS3NyvHPP
QCObsFl0vlZR0uW76jPWCFFNtGhmrgaGEfe5mdqhGePj/EGXAM5pXkhsdo9onyJF1ayz3s4Jp9N6
sXi4M1fxRUaIC7gaWwQy1LVdGVp7D9eMjc+u44SzSgEgojMMzJBBJw93xgmV2/NS4RRxXDItbXeL
q7Fp/V491GVS9NS1PEuHyJSOSCeYPEqerNffWS6YARfHs+frG1FPddFk6CBgrKcgO2gOGQ4ocj8G
QSghe85nqCc4iNVSwJhRuzPhypwhUcr/u/EHOO2qYMKmzceNwTvHoNR9gFlI8oqA8cZq47gPY5c4
3fDFs1sndb7SBIECr0OShLxpfWGXp/6RMNGNxBOzk0FRQARLf3L0LpvqDqzN6vbvsw6p3H3jw7JR
tJ2sa4L1fULYDE4E06D1X4y/0/ebiPdI8ti99ubKz9YClWYR874HIMwDZ0DLS1s4vOVTUszLirON
PcyJOBkNQTXgi/H2mNgbbBpBZrgQ7gHtBadnSbmA2FMbjeFCXG3WcKV5yt4I9JyXpnHCWpIRTTjh
C/eVxu7GX8jfdRQbJ3AOjojpzcbLkN/2W8VJ2cvuip4aN/eT+sQYUKue6yrQiKQc1J0e8iLFqBks
8fcKr2D25FAdFuSZ
`pragma protect end_protected
