// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
svs0WVl4ekhZHdHaVt229U378Psyff3etB1IP89V9jEmmNrGEnBOdr/UaPI5TgQmJAlO5xqsSbEy
AY0u9fdcAPJm/jko3aNSDad1/I0GK+zAu8Qdzw+khD3dzgRiFNdxMQ/fFEadkZ88ZwWQduJDgGeW
5Q23ZYBb4aAKVRc9iR5W0TCsV1vUu3fGGhIXdz0gPpxSsqhoVfG82V/e3SAuAIyCfbTopSy45zmx
ji/YYd+R3hN+oIWQP2nJStGmRyYIf1nMitrCAh45xIf09weodoF5SrwfsQRCBmSsV76JSkQd8MkE
bLAtMfHf/sJxG7YT+mKEQMtjDLwUjUwQxocekA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6688)
drpgNr0d5auMjdOQUDDi6kk7zVRjKQq7l/ekINFhOUVh6szu8Wegaa0YkDC1B+tObHNbXNPXKtgc
/Zo/6ZA6VVpQ5BXpk23ROrvCRxM5e77Lf8PvCrqogT7cJ41biYjgV/pEW4j2W2Fi+QkUw7kcNES/
xXu68SVU1sCLFPAeqINvK1Msd2nRr3RThqidSPTk4ni7l8DF+VpbYsP4kMRBjtGPIr2v/9VJO44L
9dKnvinyWcuC4udxlbjqF+tvICIsxIrJJp1Y6A65stFzoGdwS2WgTICih9DGFkKnPL/Pt9co9fwu
NBxQGnIakYAG/A7NviUvh2noWJ9yh1bpi7dcl+p8h56WRpCJtSb5GcFKY3r2HS0MBMrW07ln+NNw
8EmhBlabmXyTgbSEX+BANE0MQbfMoPCO41UBuvkAICWL5LFbGgzhpibzLFgEZLnrQjLmih6jDDW7
4qVCHr/Ba8hh2SrLdgqCT8nXy1QnhqVzSTvrGucSbKpOO+YIOD2tptAJJZtEyqLAJbmvydmvgmVV
n7DQqEjjbmwHV9Ra1jvt47MIGKKkObHI5YShnnpghrMFAdTBLRsKJJRtrtmCPnxai6jXaZ3rE9NT
skTRB2TZtKFKFtjO6muBz16rwhPpUbUDPg6I7a1IdpuVxC7qf4cbWExksLidR6YzVM3Wrn8CupFg
Tu/6fGm86JdCzXu1rjeUng04OBj0rT4wE/mNXYuqjnD9vgAv/z9fQF2rLlAhWNlcGIyCInw/NWqb
j7Gu7AuWzTtpS6c272dszSrPCkZ+BbrrcKkvWTpm5TFkVSn59USKQqTh81woUZL1nvFBYAPdmnK4
ncW/L6LGg8/7EZVz++B66EEdOB1Y0qqrjm8Ha8isIpPKRq0CWzdMtCwzKOB2oDnwlcTAA6V8qsqO
L/LRCZXGb8vVf79iFYuvxVYnTfE7My6lEHk8U/8Mk+BkXVd6dWcA9fDqBjyQ6dzcDAj0CLVi8Of9
YkTpqhZ1RXr0QksAy76aOHyUws8mP5crIvGgI6/PQ4zVUeVQeZb2tfK75kfUNFyUQXSjVopRACSc
nGWN4eUAHfFaX541YNKP5sJeYe78d930bm/JHFFrNtW9u1Ac4QGYsp2QYI+5Wf8tKIxW18XhzguA
yomqbqcBaT4oRT1Ks405XQdLpdqCv/6tO2KohvP1iEAO17XAfooJciEigtV2m0AUzFHLbYqrEYvR
eHcSaf5CKYuZidH22rX2Y6tToivu79uawMAUaHrDsv0nt3RNRkglZCB4Shl3jtLET76JDtaPi8S/
VOp4xam02GAgm5Fv5tRJ9bs1SYivBggCcQbV7+W8UnxcY72pduOofvPtwqfdUF5IgomfVChos4cE
bIyOx6uarVo/sbd5YtDY4AZtbzlba79h7HzqppuUJG6MomTnOZgIb2P0LWUax1gDTwHYhEwQEELN
uzwwebcAbant3o6DcvJ+e2auK/jPQz6maPIXHAtJ5TcWUWF2z4TFJ8fHQtX80QpITKImdqklzQSV
OPfpKas5fP+Lw+ZVBdY059mg9H7elkGgyXMW0JH8K9aOtMR4Vin7YZOZhBd4B9+90IuJ1axL/z7J
Y78t7JPG5Qjq/u1yjqgbEgC27EkFLuUP6YRYmizzhb+VczDuBKFm/BQEE2TWEXh3qVqKMsSKztbf
6ilaDXRYSwwdY2nTCVKe/s/unGHKvoXVBAyj9bl23wvVPjcGpcjn4luXo9Bww0/TkZh6+3sTNrKr
isuPEO4DoDFEoFsWZb7ZccV2bRFdVEAJSpoL0ho3n7Wzp/pOIZRCrIoNpZEK1gu97alVDXbpT9M6
ULXKy6ml/TO1XIPKU2e2Q53qUYu21m2SagGaE+iozhZOFLg1+JA/CdLEBf2UbfBff5Nqe+tgAyoz
SKvMTvLVSaXV7XYpi1Q6czNZsYcT3vkqrpnNraQcajjcue2e4kQjdGhiNUJtEp8Xlc5ER3BaMSTp
ulluqOrO6hUKaAobFn38+5nTS9q13Gq3udJXlo0XmMdWovjGa23xtT1jeObZC1y4VDCMl3Ttsflu
vvUaIjCn83jCwS/q9Lzu5xq5a3yHQ6HBIgTJrfuZY7/duKKzKvFOPt4wuZItON/ADXpE6VRcpALJ
bbY9DnWj0SJ9zuCFYszN41EBXfes3y0vzwWqWMYLPA46FRaVFPoR5ZN/MsnVVlz06++XQaNHJueU
9r6rrPB4gPkZMMlWd6mIlL5GI5hErsTQJw02MTbWCJBxXNaJ/f8vCDeth48eHsFArtEMjCoFlpvk
01dywu/rz6WicqFnkV65NxlL8WN5L+ULwPVjpkZzKSAZsn3whEShR0vV+0ocCd2aaYkgOXRP4MI9
jXlZnsl2asXTtSFi25g3PFmnm3jSdldEXsp1IWCmpfWQbZjPZ9rcDR6rZggDZbJjVeKaQAjZY02G
yB3jeIkCjp3/QXnIPu1hADIRHCwJkLqbrsj5qDiR3xIPfE7y5hNKWGoE+AV6WsRKfYOg3r3YQXaf
Iz7wzcOVQhPlUyThF9Me/MOIlMEs48d99UYCvynerLI1CNohdJoK5BHGNDk1bpz5tWl2h/r7zYnb
gmUNJWHH6E/7RkZABpQ6+/557r7JWj1fUPHJRzYrFZsc/I9Ymu5Z7RU5++m4ea08MbHZCbQ8JOb7
dJVRXzrqHOuhULq8DHIuUk4Z/AwnM6T3ZzprexOTkKaLS6sI2vpQn+QMnvWC1NAm5LYSrQUekVEq
Vdaiw6mphNv098B16jG3Mub0WuvCiUak/aqHa3vz1VP+EXo6FHcvRq0uumq/6lX2PyFnoRPLulFI
6HnW1HMLoksD3AwynXegNNcMiY+5EhKa1y+OKmTHwAyYBXowUWX25WVdwBVsHJ5VxBM4EGDwNRER
NN1jRYz8qSn4tnYyOD2w520D7R6xlJN82iQNtgI0yujl6m0u2JqxIy6Yp9qjwH3mmEN8USejL9Ep
R52DHdCzHtJlLLAabZkGxTvpMrz/l7uGG4JgmZ4L/tKoiTueEVsgKPJjB+krmXx0uoFX0ySn7a7+
nufCDzYIhCygPF97JIp7b2hzjigzNsJLiU6Jz6QVKcEHLTmB4TVK1+iu63AwMnJwJ7YHZi1CF7zK
xLjQWKbnQoO491ERoLPrBLL3qK0ysmfcvMi1jZtaQ6vUVDyu7QEXuq9QVDBlV/TnUEnlnhAUqJBp
vAC4VYN2BMyDsTBedbBU2tI8yTcpN4pwz3keyE9LNSQjj4Ox8+hNWsRhLXIq3u/99JK4niHW+Is1
UfUIdF2lBDVb5+9HFHGd/0hWIusG+Td24WMNBJrhZLtKplcd5q6/3ws9zaI1Q4cNPDGrCcI961lI
Y13Op/boynLHSMiJ55Rg5rXtnR5yKW1PlkArj2r8RPnVmWxraD4o+0IO8qyeoxY5wre4inazsG8Q
G3LdPxs8bWdjim5z08mWubQJC9/0j5GA1wwYahyuufAyyzVFIYoBwtFcJ5KR1oqUtfb9gu64po4l
1ghkmX6GanN3jp7o0QWqdcPFAVhmYbV+7niAGHOfgDra9MmMscPyMYvfczsv8zusIEz2uwuCJwxx
QYex8VKXASxPCmTpURDj5NUWiGSXkxXHELsH39HhQIpyAPLQj+ul5B5KhV6Y4LWfMknV3uKcUf7E
W6mVy9o5xT17u2mcyAAP5zxIuL7BFM0eww3g2X5H5/O/g8D/edr80E1qoVtchWe9hn4nGda7By79
lCeiyEjftZWIvXAG+LX9rjryGakfk3BqqCUXt50jWJvCgzddf4jNDtnVqTHhPWI+xUDzchU39jp8
ZIbEsA9djH42ZgH5mkr4OZ3/OEP0vXgVJ5odJRT3yIDZYRH5687SlRUMwBBoMLadmGdh9B4JVtq+
jcmd/gR7kAWXGSz0BJrTABVysVbDriDG9piXL9dOAXtl5hTg/oHtBv6HI5V7DZ7ofsIdSA8yEXIu
hnPMvqSwbrkWpTnBhXztudYlrOlIM9UZ6t8xoUcw/iIIX/9H9qtpO6t+zs1pSaSoqse2qakngbUt
FdgSPagvtQ5Idl7yFbMUN8eA7dtq3OD7q3P/Pscc/OjnXP5C8Sta1Idf0tt2YTK10C2/anwb+p3A
qigfjkNDLAIKQpOMs3x/TwFLf5dSNq/6cn1hQoxDFSAANYGA+rgU2Cf+/cIiQmUmfdUKYJCA8ubW
aQ5BUwRps1anBq5ZKFyDYYh6J/64UoZmsixtJfyBI4FLMsQh8lJLMONw6XUWKgAqorN1y7BFXt7y
bXSt/UHiL4dChh9Cungspza4We7RsdxKBKt8//7No4bVXyg8/B1se5Nj5UsRluvgV8KC7EfcY4Ho
iyugiuP2FlwG/7+zx+GSEvRzJEyACvaVOBm99J/j06h/aM82utvNyNhUar7cUaFuF9YHZ8RFFBlw
aW6LFj3EZIy+iGos55Ib2nQvHSq8f55dVqCM/m0gaktPYTtifyYmPgm8j23s/DeaDmXS0OKT33uj
LxU3HyoJpQZ3ttbDBvvVmxSGWBqsudHidJRApQgDpBQwsraS/I/Wyp0PWF8SA6MlLnr0AvFetkLT
1EPiRJj3lOyY2JGz4zvAM73cRt5mGIr2jtpz2wJmUgy4DYqLC6NMrSapCXKg2vzd32uqAm4eiEll
yzS9Bq6FBy/fivKozQwCpsAmuucpcAq3gvAc44PJLURgHsu2yMS53sdndDLkIxbNq5DyMHpJSaIh
NKDK6wCthgT8E7XI4pDXtXzp+U1SwOQOdJ7V4j3M2zRhErfKdU0lgTBqEqC3lQR5rNrgk+0p1zsM
WZo/liv4WbbzszcRJev72UPGFIfoYOWv/5dBdPZkw+sBYtz0D3xA6sItyB7DX+Y6f5oLIGcNcbD/
h8NXVi1HC9v1ECsIQ2xjlBKMkz/1B97Nk1DUVS6V1VWUHSabwvEARr3ZouNYKxxuvl+lZBKDqrMb
lLMlzWKA6vsVBh1tx+TSCppwL4rZNLL1I2sXNtA/nwqCKVLxgah+87m+ksh4o5hnE4TU9mnHNt0o
xu2np9tkfoPRZeKfzdnlkT61g8uEmb4ASpNJezcNsGu4Zv8j7NS8t+PDv74lb6+t5e4MALkVzaUx
TZQrUPFRHNCSj55QB0EFdcbyFLOR0rfG1lptl16qy6gmjyqflj/GS0CwJdVE2ZZZCKPwJv/eYZkf
PCVbKqxN4RAFis7tsL68xIAZlZoq+10DNTAuFDz59nXUHOf1Qd/F4Mu1gwbzqZHsf2Tisee5vVdO
QP4YyYqERgdqtkdBj3IWTFO1NSpvEWLs1EnViot8SC/Kl6dXnk7oLImAH1vKjG+/8czrcd7Jhyoz
Dfd0QQtMQIDZDCEhPTvgCT+JwvOI1przkLuHYy/mN5Vqvm9xPBEL5flg89Ak9JsaYpfibQwcC4CV
ulR1eKdaUauurFgEfJdmmNdyCW840qw530vQ57E/DdwE1cxiAoB/vGipfPkHAl9dC/hJTZV5nUFv
voZzQB7nzCkUNWzTs2SF/DNtBQXDOoWSyxeJ6hXgzRJw94Tc0NtcelZQ7FA99wB2qUE2ZIPHpKca
I54X7ZOa5arpAg6TpBZKmJo0Zi5vO3BDlxcggunfxf4Y5cCsTM0KzFY1OV8z4AKhUBXDkMUBurbv
4v28F4RMCkQDIcBiD2ZawwZmbKqnMKgz7RieK39257V7bQZQiu21TqhtIkMeWmR/c2qNM3K7ABOa
hG4nVdFkab4nbdd0LmUQEPWgfQao8slbpfu6NqjK9XEkhXJfVMrDromFIebkZljtyAmgbmp5jMu4
7c0AvEp6GhhlGn+BXWk+t2sjljgV2hHEAMIDZ7k0jibuCKle1sX/8+vlq5riR4TyFuLus3CKrE8z
cSy2PbApBw6FMYNwtqlRPa89xrF2vEcl7YWcvt3Uopo3Zk6fIHYOUNDeZfiTPN5y4ptvU/8lthoK
f/S3ZWQXFxqyL6Tw3BlkLfOj3eGva0VtQBRSoaWWfEdud+O3nzBwCsoLs0OMRASHBuYKTdcv6f/n
1gaZCCNqgE2QQkcLw1naeYxH5BTRnElc9oGxBpHd/CToBS9WTbr8SXllpxfjDhHqvyWgkasGZG/i
1z8LXGtbOuPtrj5xLc2PCc/MhOHXivjcFmtrSjmVnys/82ub4rM1oa6fMRUtGZPnoXyJty1FCjzO
2nYONr0e6wW7qFNK6QmOlSwRFZpZpP+lAqZkvW9S6AiOV1XvM+tbhf2RxXx9fCXVqepJ5jw2L7gY
VtKH/foeiZqaCjM39faKZDPBfylbDnXHISkw3RiswKqMbjDxyxGo7FPEvdn50tRYldW5JG+Zc/io
1Tsrc3LkuapmuGktjNbNiSvWZdTSzv3Fu7dnr38zHUHpFlC4j72BKuopq8ZpvLXlgWQfbROloJqg
NXnRlGW8c1/7Cu05H8rAT7IKrrwWRD+FpMsaQy7uOeG77s8WVzWKySdvwJgJ5j4CHxjqk/Yn2VPp
bakT+erkADRhhBtrxP4EIy9piCmo1ekjEuDNMQ9Jdu2rRMhLL/WSTmP0sjf97IH7UxCQ8UysxNyX
cBuMk6/4joimF42q4neNyuHnoD8l8X7MctAsMZdzpWaEk1EfdTO1IWeUjKGFEMsF5MJugyPtMNDi
IOwoPiJGvga45nry0F9jQ/tIGRxi5WRnXvW84suO/7rc2JIhbE0fx67UGKZ8C7XauQctLJwnVTbI
OaVLV2PmO20tFzwKF9HugIexIrPElLtV94nVAcKJ9a7UNMPJCCzVLYBZZ12JEVzkvOeT85xYF4h3
Xu8M8GB2Uc2RdewXSf/SRqrCVcHqZKUszs1bdPutDMJqKoi7eajIrT+YLAfo/5H2Yx+t2Fk2AEFh
9kB8lpexufsDYxwpEbx+E7g59uh8KTxnliyDWKdijcXiPM/jmtl+rbqKpzYC7t1sOrG78wWdi2kV
MrfjVhGCdyVLMdwQQ6cl4AS3ATffwkcSM+KPHUCLOFAgmaUgh4QxEC9wBsV+UYo9SLhwuEf2rNJV
Ua6wF9X9g2wOfxYHrQF3Dq9DkYK2fYiX2WPgCIYHE5Sux4yl3cU1hgvMt4aZFvxXRFAAiUd0bBA9
kCJtZ3Zo19GRpmpjB8HjMaTtDFB+3889UBstITxOL3agltTrBPwjfoCtKzqWOU1vzSZyuCswEuOm
E0STLVSqhKzChU1fw5uzLzr2EU7PdSDh08JFgciLsRSk/2fMGEmVdssZNnKuCq5cFc8x5AQ+Lzrm
ZafIEgFrYzoxq/INXwv5ALso7AXh681MfqafgacaDcA1ud+Zm5zZkIS1rf8U9uu/mB8N+HNgl91D
xqGWixuzIWr1GmuIaBHS8Vw5H0erKJtpY8g4udG5rDAlUpwoSiIut3US6gU7uBp52v1k2DfnsXpK
lfwjI0GFii+ViU1IttVBp0X2GvQX/4E1zGdFZAj/iXwPuOFoX74Jzwmy2afBboOYlAaJ8+1Dvq54
tcPJZwAcUsqrX4P6kwji5blB6LEf52GCy5Je26Dyv68+Y3wh3TNp8bpun0JVJp7raruFnqnhByKb
th7LRBuzRzbh569xJyHkHoSy+9TNJgqN3UDJj1WNhoKr8EduAvGWLA70r5/UGiGAbJtr9uEJxqNM
ZeM/pDBFVfq1Uz5lJZML7Is3JKla4fURDjwi25IQTjZvMtB81NY+4x2Zr+O1llq94VnOK7iXDC+x
xRGdtOtD8oEtGhTBEolYbwGZl35fKtl2C8Pl95goJDZvyvbJxw0gGTGVl/T/Ody2HTNk5fhwE8q/
lqQBw1yXDJNIyXcdQ5MR6VUtdIH/yVfkP8BvW/JqCrSLwXGvCJD0/W40mRb/9LDMvYgHa29bS6oq
5JsOB2uY0AwTLp7Jr/CkZrhRVKZMMn+G/mSxv/ut2R2IedbFIkmfRDhpQwCwVvI6YVso5l5lXd8w
iVUyAOEvPmoZQ+4DY93fPCbAR14682O6cyTm8fecClXHouJx6xZHuDbrnkxVdd3EZ6Xxcg/Q40FP
94hythrHNOkXT5tISPrM5XGeh4pNt1aDO+wyxng5blz2pDe/IT0PabZKUZXcO9K1XpV22UWpWVSW
OxchX/CHv67N3S5ukh3uDPvso4mV+SD8wXNow4rPTVK3SZ4U/hVDTCf4KF4fN7JejI6U7tmejEDD
X2sG/PGkpFdTw9WzY9OMYsMUNBMyfNpfUK2PuTPwho3eRSUBlSxiQ0ySGlIdByLCpz94a4fb6icD
5ab1p7DuAhzzgzlWNvw+4k17Gy4WnbWRHbMMyhCGv7m7igjcQRVcozG6V7CsQneOlvbrFf8DKw2F
rXqOBbTAr73CoU1T90zIznXF80SVC6wT0I1tHH36cevcekHy4h33xIAQXwa8VXT5gbixsoolOldo
/TYpMwQYcOiY621I3sNFA28UY14eLamHDqLDf+1tXRW2Ahv3DejIEYXsFC/hylPi9088R1sw2F9U
ZCzce1dJxgMp0TWRzwQwdWtKFwciBAtq3MxJ9LDdh48CCOWammNv8oYcEqdFNC6JZoGtQDR1wGiv
cFnPEkRMFb+MbAzwI5jDuWGLio3OKn/VDDPNNBlJh5I811i77EGQBMKxDxqn3maOn353xRfnKFpn
9QAPyDyPb+h5z7tLRg6n5cKYcDeEtTpYjC7Ex+34PF47hNZzECJ/ooCTS4OInqeqDKOFWs2nvj64
D/u4mvoz0B1amY5MwpaDw69Zlr6fEUYi1mea1Z9kiSEXC+Y9QZyNldBQRV4G3LKouBAGXwieAntc
kGUBp6n5NUIZvS03PBTMe1SG9MIGBzI55Wuw5oqvp+Ap1xuNgJylk1FQrD1fe6epmgN0fzXXKzGc
FDu7j7+eQwyaPvvRbnG/s6clbvnpUapUvgun6cDPiXFEkgkvjlKiMOKILZpb7fWcxdttLctFPXRs
HrveSUSrzyEvyAvY6zTZbqr9ZA==
`pragma protect end_protected
