// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
NPoq5ivm3fbQYtNKtPrU7G3A6aPj5kjFN/o2Bo1Zb8uhMa9ZROq+0AFL+jFdH0Qi
LfpdckztYBTPQD4x2hmbhzigzaedfq+AuosFQ6fsm76Q1EktvcpXRZJl5u3rtY4s
6sJ2hTriKIl5gEi7jJKZOR9Q/yjLlkajAI5UKvV92dMREc6IDjwMFA==
//pragma protect end_key_block
//pragma protect digest_block
DP/9RRvZsPYcDYKstmRwxfo4Q+Q=
//pragma protect end_digest_block
//pragma protect data_block
TaueU/mExUd8nJRXh/bZe1NZl9bnN+bXinswRPVGzrE8WNpzpt+239zGfXwOPU77
fWQhPVR0rE7mEnboJrZEh6hQ1O9OLRWQpafZaV82xxykPt0ND9CQZYz5ROe08e1n
9YSsnvm0mCIt1ksQOFpqPllVVuWu3LCMLa9mX151IXITCOpc+KtbK3sOEI8E1YCw
PbKEXCBqC0IpKxrhBlur8tNAnAE5hiB1KeH3rcBaY5A7AKq8q+IkkGhDvYM7dPL4
pIl/m0cG72+eyppQcJi78kgkJDcqn5dknh0I0g0uK/xFUy0xQ4Ze9PKXafuieM+W
4KD2ADSopnLfM6GNYrZjfTsjooTsg0PFmM/DRFoNNHrrpjl7KRvbwTVXaqgpLqNH
zKeT0KnwP6+b1erHnaLPjTyB2xHxrt/zK+B3JGKtSaR4nbduNW88We4POp5XoWMW
M7p3iaLFstEge3TzwSW003/7Tz+Dc2w4SSIAmB+dEhh6q3v2IHEqBhhVerhd4Ka2
/rwhTZojI8yIEURfO46Vlh7nHHD28ELq3idyY4PpNRB6xkpuE4Ako/NWUMrjS+V6
5gtgd4/WZNvjZ0deU+B9bDUdWQAhlM5kjYevzPU54VwYxCt4FfY1Mgqihf70fn0v
CKXrgWNcRnFUNU1wqAjkhNpJMuCDYO/2c16XXiXQ32Blsi5oF+IlHAd/g0b3hH2W
oTTm2L12EZxc2jG2I0L410TaYn2f9jFLtTp508DDjcLRZdENHticfzWFz45d2aJB
gOqEFN1KwFtbKlVnLoutvmme+SP6BNlCXwiJAOk9GT4khrJi5kAMXCzZD90Kodzl
/s4kxyGI3qqrmci0f/3KunqjTbVZFs4gNDUqCgc4g/n2rx7tR2wMX7Y+0DJialhW
GgASj3wzI1kVbrciipQAQaHQ8Ia5gII6k5s7+9jSTr+Hl8ZQg1BxAM1FfnkKZiRJ
XA2b/YwimY1tNwGoONBs/MRn8wRqm632JH8cKXcjJ3eEFL7KoLVPxSZawlZ80Cem
7SNuHjxB/ClAEsP4a7T5UHNQGMyBPhv2YgBYaVOlzUC2/12P5FtsushQaO3T3asb
vxgNjOmEj396Y9XNEjmNkEvW+ItIgl4AIKBQl+kvOqWUl7Nvv/MeNMY4eGLj0aje
k/2ZfCMAHGbGECIK+vJrrJCnZyHRjWnVcdZmayeLStqb15YcIGPuDV+9XTJNFawl
VuZnr8ExHP+tJZ6WgHLSd7fpNWuRG41C19k/HVmXtkC5GULRJVE7uVRQ6GJB3Jf7
dG/z5NyRx34tuuIV7LAUDI2ZbeBXO7EJY8tsCbRFLJ+b2DVHuWryqLMAQldcmFvT
vaZ2ybSheJh4uHoqsDJjBxE/VyQH56LyzzsJuv4EYfc5FHKu3gWzqEfE/LGJZL0G
VemfEVLRDQKsULYQN/8+UWme0n1zSkvC/URf4VR7HZHZMdao8af7crd924695k6Z
Nxs//JKg49rsMn6Q8R/G00jRqCZI8lxWQIfcDP3P3g+s2ePMhc4lF6Qd0vgRjTI5
k2ROF6fhQBWNbZKB0tTUEDKrHh+XwuKz0TrrU4M4CW3tnHrGyAvE4+reWLS5kraI
FNq1RZKEp/Vg9y94Ru7l2Hwyg7qXV5z79XirSytztht1ttwjCIMbqtyNxIXE0HDr
iD/fpQFA5PiMkWgQMAOaJwMTy4KhJg79qRsDHNRYQ3Rwk7moNluSXg/gH1v4sLF4
X++ADq8rJERGcEFpGq6TcHgF/W3FfH6GF8AUMovDqHTYXxeEULlseE2dWd080RHd
2hAaQtgOTClNmFirnQjYQucEVeb0nOv7HoC802ymarj0TUZsIZ/hN10jkaeiF8pF
HSqYpBEnyypYvz1kYX/YAIxr368d22m50kGBYFV5KqC4iP/K62uakramn3Ng+63O
D4Y/sycALKeROL624xQhFFLb0ZbtR2IjvLRajttdnaBFAV2pCoVWxYwlgN4WoVBv
Rzofp6lfykBnwOqQ86bGIUXr5UPJ+BKxvCU/vmMrwmQ1hBk6ENO4d50Qg9uEFGQ/
eLj260PDfVPgUV4aTZ187HMobCzVqoe0t0lqfrhOtiFu6pNIqWfglqlttWYdz1hP
CmYpEbfRXduG2SxB7CDgr5j35ixFzTzB+XgLVHwjJZ0wiku0GrxPVSNanxppJEcI
ejX47X20ZOM6szzsNWGvRc6te5gMT62qi0zX9Alf1bw3BBzRgre50pJNTy7/0wRc
Q+jo8ZJ09Gce3/yjcF0bI1GGzdAS4X9sjKCFmjTtWjhK7M8UNoWoJRi45Lb3Bu6p
HtRUilKzt3RS/lnG1AlpMoVQXp8O1kVBHtw7y8J1kUIVc1cPkI0mm9bURyaeXxns
uiKAsWJmNmWqnvUHT1Rwvocka/+5YhDc/jB1UO9uSpL17EYnKr6EqrcMVnuhPntT
vnJOZZx9qw/Nf6OAPw8PGI5L6B+9iSfOhVZJxQGpVF1Ad6W7PcLI9f9cOXzLK2GY
IrrtjyC43HR3bG87TFfp7pCnH7Un5sDalERMF4ZdMq1B1LXn1HDy5JPadug9E8D3
1ouzXZChmvZ66hzx+bZAB4lwbMJ5wT6PDCOLip1Cl1l+o9Dx5EATO11CcX7RlpDP
G66RKR2jlLZCmxTO5cdgpR5ojTSU5PvOcBcIX/vJ4eKOBRT8e1ROh+3sHgsiry/u
+1S2o4qjMU/LwCpczo4USkdGebV86u0UJwGVx0aLp6c/RU2Ol/77d/KWsMonpxPh
wYHgLbs21beTiqNkVJMBrHfbuykw2yOq5zo3jD0lPe67jtbNiub3h9UgoUGXiGzd
J43yJKhjRJX+7Cbp1sG4RIqSOM00wKdM23gFjrkFBTVE/R5im3Lv/u5tpjXkYRtc
xRauAne7IoEiqtqmBibiZXUaZj0wsC1MEvplic5dPv54KYdSFZnmBe1uJD5ECLz3
oB4Ayr/HR62Iuw7qLYWrDQ1o08uRzvRq2Y+XFtiSIPkFhBQHNoxG9STfO2io6Vaj
Aa4XSI7Kn1bILJNkdVccsacd5uoKO9lpX4CvuZVdf+RnOr6kkdTyVN5xz3F01eRK
y4iuowOR2GDnw8vWSohsFibCIVT+noUDW3EX/vCzlVK2u1qaaqXsZcaezp/NyjPX
xSl09Dg/kCu0RJnVe4QdAXNa708MU0aKHMuXJMFy9CGqBgOHPONkKZlRwpfH+gdu
PU/xnT2NZ39RBe/gCZjg2fQLPRR9gO7KHjywjEQQEc9NO14eMpylQK+YjOqdoZrj
KG/6FE+LWcuxYqtfitvimGV/xBwPQ04gZx2v/Wm2xdSYyfJYfZKAkGXYhcORNU8y
6vm4RlqZ3qesc2n95azy4q2rt8k/7ZoIbTbFPrOVZmhYdDpkDdnZodeQ0Li8Efqd
TN3XHmyTsmdI/f8qvqprCG2llX8vJ2bR++x2lhuAigTF7ssYi340VVvM0Kn0klX5
Vrec1Lm61E8IPtkw6y/Z3jPzJ4dm/xxirEIrCYU8KJ5JQ4V2XrOWeP03+wNg4z2l
PMuUZszsxD08ualsNo6vicgh4C6oLqS7EXZa3rdy2WlIFys+qBVf9EA9p5RAkrIi
uMuX4n+hpGEhRQgDlxEs4SYb7hVOEMF/lt6fXGoid3ReVyzP4ImK39M6l8xEbhFS
c0nVva9Rhooc5uBI6fW28wn2x5Sa63LqZvLOTP/0KgrduvxOyH6oJuOizdhP580q
OEPCtzL6Aj0i95NHWJl3tGU/j/Sd19bqN/oxr1Q3kBs0xBnrFvbOd0vCSg1TGW+r
YNrTjgQNWp7bwy4uJc2yl1feJUEi0yjP52ta0gCnaik6AQ0BD3t2pILOst8Y5OgU
QvITkjB19z6GIALxvVdnRhZKSAPYGo74WoCSig8NVZ2RmqC2purfFFEBo7OGpTUw
9BG6GkiWOCw28Jgltk/MNoaWBLi4CyG3U26H09sJg9aNOsawiG/j2x0n1ropCN/S
moV6HZ5+JSFTv/2GwNdZKrI84TuQvq5MvIBZX0M8tTSfKmuCyj4nJw0LTPHc0F5t
KOA5UDJP/CUKNd9BxFZvFmOeT/j5ckNcbspzpMV8mOm4aAQQ1CSFZyeotnoIQ24X
D+58+Qm5CuWdptqDbSG+JMDqL+7mpK/IWmQBGqg24B5QkQ9TBSo6IRMVLDjOhJDo
4g5UsHUEs4Ic7TF+BuS0GrmESkPuKHE4VWG3+XY+36i3k/BaiyHh9DDraTe7yF18
D770xO3/IgnWQLXKh5vJVWzmp884Is4hzIwMxNWZifAxcvG9lQn2Nnb3hXowe44B
spmbfMMQcUXssZYMiJGNHIXgaS3gbTqXBIJhJj685Kj0BF4c48cMXlR2EDz5yuB8
CNP0P+voaJZMMDdoC4FdlvzCU/fMt3fioxAnKXjYTXeR7KivA3//RymY/Y1h6Lh3
MoaAn/8JDDR1heSmxY7ZOt4oyb/B3ib+Dx8EGo73mccdErFh4h+fslt+pPLV8/OO
MiyAtmPeuAKC4y356JxGhnhJjj8W8/UF9tXoF13/EOhPzNRIDfey4em8RPaIAx+T
/DzUjekFo+aTXnWtXRQ2KwxVdqb6aMlqKg033sQICysRlaFeD4lqTwPggTPQm4p2
N5Iqyyk00OTk3ugzi87fLHDF4IpbZzFCNp0bGw2cgIv/ce8Oo8tqkAI9RuXYuMph
k1l7FEL5k9aYr+262r0lW+WZHlFkJDfmR5k6MX71eM1f8wiNXsDpY17/+ShA0Ugl
H0VuPQsDyNCV7hv/hhhc0WWsmm8w5gqiWn4SQaFFOGg+bEFjOs10vXM8RtWpB+F0
5olf24wcbMOQRhrBDNjbo7nWShMEFBqRK3iDk5tI7XDrtyFZ50ZjdW5T4pPWxQ85
g8DneabfkWr103QgVENx+5PrOtZmJ5KJmXAlzA+olNQXgkChywMRrqqmMV9uPnCg
bETj9qf/G4/CKpt9099FcRL+eZvv5kBVLdc4UEoKcPk+HyhtcKVdaAmHlt/vKA4Y
kWIyn/LLpBdQ1lezvd4NPgPfo5/ozn49BC7s8DK7G8QydDwuPo3/i50jxepsw+8u
w3i9Li/bJSBXBSIZHjugIfdX7JdJzkBjL+8FpAQs/ywVRHomJpXO/FuCHYDn3Qzm
NYfLxYDweV1B7i/HJA1bps8SD5IVBuSqHG5g/QsHibkKNxLICDfAWZ5rg4gMuCno
2rJI3wg9GmOGNHRzgBexFEremRSPU8gwHso7aRh11rDdUizyuUN5xMKtjfMUK2y3
YBN1gP7CYaNwQbapyXQRZ9SXhvg2kBqi3vCNnXQuAFppP+EfH3/sZCn0Aa5TYljd
lkIEJq+vSiaInpb5ClfXYACEEMRrj7xnJeXcfwhaYujlRLY0i8eyxU8po2C+6azt
L0FXIDrRyeQEatelpBkC8ZtqxKom+H7DFb/z2u/gAUKjOUd9HU5T5uhNtEkcQ0qd
eTUyqoj9zCfqR8Lgss2ytqrLN8HMLsCiXzGJAhkvvjZnA+364NVqNKntoNxgohO1
Mfq8VOpVNEg/gC1CMxhXof4w4EZqwTXnee1Vy7T6PSxB8a8wYiOcAwYEACBX5WPw
qNivoJ7pWi6nJ+yP+PCU+Xu3hIOXyn8aqBB39yAUj2L47NGM+/bdmCDZFSnYprqM
8pF/GXwznVItiUDvqb31b02I1cpEpi/nrVlaLqDVW7FtlBnvJiRt6WEeYPcxfxNX
LifymcYOV9pZT97lx9gyk3J3VPfY3MtZbiT47/w/Arnyy+8ids8IjDRUPjCjcBm3
CmUw2vaqv6VD5V6I437hpRJEKJPPKXy608X0KkYyyZiLjq6SnTE/+uTUy3rVqokC
sZaNIupTJvB/ICXxsp57zm3VtVBKrkjMrr51kxRsSl4gSqaOFpplvk7+4DE0esCO
AbY6QwpgEmQ0aiJ7mYYAaSG5YJFsrNdhjUYAqEj3+7ApaoA66Ia3YFpJIJxavFuS
o9q53HNVcW7CKe2rXD39gO1JL+JsuUQBTLH9H4WjqKO+MCjgE5RLOt58Z9c056Y/
l5n6m7/S2cWcF2MTBDFhYx2mV0C98JsHQnOsXJ3qPmevi7nJdip3eXCDk7N4oI3z
pL6UOEzm1zdMl349KYjykD6fL+6HX7yHK5i4/wBhKq1oR2GJqz30af7jtUL+b+wW
XtDyAchYT3AnT0TvHKBf4Rfe7OK40IMXTWofg3y58JnAP1Sw2l9ZYEnlONQBSY2H
Cii3ssZd2k+X7yZGaNV2sw0mQ2KKX4odrP0fcPedwkclHxKBEkqnQcScM/FfxFoo
c3zoFg3WECjNqZq7kP6cYO7EYvNPhaqft+zAycOjozI4ngcRYVeMlwlq7ydn39Lf
TmrWQ0GVlGnDgYTPZp9NzPsZ0Y8+0lBkX+qLwq115ZeP0FULqJIgD/aXcosHVDW+
eGk2pBkQ2oJRlWcSk4auq/f11kg2SxZ1H2nrasdSB6FxA1JJ8rf25UkEYI8BMEVw
j1lIs+AO8/mfiToHueSs0ssoWQigKDxvegFQqVsOFk24MRIf7h7t0YGDSznx0UQm
HqMqT8DPJmfl2zd9CxRkFJo3puE4L/4wo+BYd5dNF5fgt/ymM1P5STTSRAGr6wyp
0eq5jhWfzV1wAG3is3ihclJlXctt456uh/0Bs3Q98WwcDGFhDn3orukH/2x1M9w7
7hZGHxNlah3smzAhXItsbQjK0B0dJs7Bbu+3KH9+KBR1Iol4tmbx6yivx5rNYkUl
sKZOeo63oZuwUsQimQEyFYXavc05wnI0jXIJP7gUKJLZyWHUWpqgoLL1dy+WBoQV
60RwDWOJYsLNUJ9KN2co3FG5fqKQ0vY2iUVZr+qKuA0/BcpDDAK2Yas3gPpSpueW
foJAh/Ac5l5F+oRUQWewzY8cobatmg/ePybcCqYlwOB6hq0oOGhK81+UIo0UE7A9
9jQfF5MztHVSp8m1Y8MCIOdNA2+F4+/egpjkFKHDZZxSHdMJF3n8SSqvyFcdks2f
MjwQabt4Vy+UGDaAhla39D6YrbpDr1q612qPbKYVaYrzHKNZfCzRdH7k0UpPGRX+
LY9GiXtjgo6sB8UFnFNgl1UvBZ4m2JZG1Z1LTr5+xzEZsKIljuN0uMUG+fVJ+z9c
pasImfwT1dUPf8EBvPgO7Z6sE0xLvAUXxp2wjw+LgLXFlyZoi9ccfLbNBG3mmiXw
nBXUw/58CT5FzKJ8Ijo4tRwZ8l9qZAxM7p0FsiIwijHCmieErF9p8z01XFM2XgRx
VzKSLe03ZPoRimbYGiv/wOXbfnUlV7krF149Yx2IMc9KUVTqL7c1LPjRmPFU4Tzm
iQ9RSdoPWkxSym3gWpgYa6jBZzGFGUs3jJX+e7MGQA5w+B0RDrU8/eOOqO9LSdaI
hhMQfSLuJHPFkGCB/Z+b2RnQc5+8UBFXvFsDtDvArZI/QA+MkXlYVje6h8Wc9Y9c
I+SjFAnNzOLYTlpGdsqIm3FbjWcxaThMEAhd9+ZmmSQB48p8aj7wq1GGsscOZnq6
nuU4y/3u1rCslwdksd2TvY0SDd+vNt8Ua9jJ+B5vGCHkNdXlI5gBn7/7MHLNxIe+
L6pBzPb7AxZt8hoFU02Tr0FACPhX5SB/dtuXys7oC/8SrWM/fEv4ijnkemKPqVCc
lRclG/X1uwUMyH9NZphBw40vVfBrayEhLGaL1RIHmwRONTPzMMU0xUN81HlgqO3a
wS4B3aQzhA899jb/918eO1BnnSJfP86Y3FKzI10YZZxyx10XHUPdph7dwbh1LpKY
BzffQ8OaAEiWVYt3+ufk0oodORsIZKIDZ3EPNNfew03f6dCXxZVBxYFCUIqqFkxD
iUGb+d8Wtp4mnTqTWIwaY/AksObuECTlAO2pyBaVw5u17+i+52UnZB4cd1wA2owc
UWbSS2zOuAvZDfb9o6LgXGmQFnT03KFMalAjY3HWlUXgL6xJrp93HGql2MngQCz2
2zW/mt92RDAWOAg18McuvSlfUz01CXcFNjzoPUCL0T9FOQPLEa5LYCMEpudxCaRS
qf2TYbhq2ypF38J0HmvuDju/R/5PEBDpqMp+F3Tf9vvdXqpmhKkzaxJCQ3LE89OX
eswndIaGrGTLSRQEkd/sa/EQr1nY9gIqjEOvouNCCWgWwTMYZEqS821X09t+kGp9
pQJnWDBD7+6LLkKI9CTufpGQ9+Qr+NOzPB+ZZBqz+ThqNYh4RzAnAJYImn1PBzjJ
OB27bbGB446zVo8xqBTqxVCNoghStmWyDRgvtN9USX1DcVyiwIWdezSXvuZsbIlL
3XgcMRtShPiwh1cbfKQRxFnPiqm8a1NGQO0Mic5enNW93FadyZNuYU6dsquW4Jgd
CUA5//PpvsHkRXLs+hYUGEUcYcUho5JUI5D1u35lWmndaq4BNw0jIvXu9FTDkye5
u0KSdWwUNs2W4UcyluEBB+JzBFzaal92w9DnyRkD/W4hS1hJKpUNw+o8R7A99s5E
hMZ1nfKZ8CsAr1V7Kz4HiFyPjuoJZQVJRP3wyFeqrqWopV1RScyO/emtBwfR5q8x
zfYMancGUuYb9f/nKtPNPcvPHSqGasy4dQZhFJyWXdwOJEywDgugRo7zBqhrOnI1
pW7Y75TsdOcxxeAyf1dW3PbB+G7wqIk6euoeKcN6n2v54ytI7C6H3OaW/n8QxC6d
JrkCOFIDVpQRPV0sh9j0lL2q/Ld+U2W2V8VLSL3/Y58JAGLMP3JhiO7it0LC4WKW
PCLezHpZwjbKVBjbZogGy2GyiZZgcMgdGtmbsasBvXyM08PzXw0WQG+qXqGW0/CI
MkvjwvUWIfC9T4WLveeH3yvj1h21jcOQOMjwRTbVRN/N28tMA9dMtwHuY3I3L2Mq
klw1VJVC0VWrZjsoYieav0QDhj0kL+aJ8eEJpHClvPLNL8cJf5IF8ToDDDpjIILh
71UoQwm7fE9JAYfofGGW6b1Mse+PlnPKukwHBfMKls71b9Aee8cP2I5ex9n69bfl
Jibfj1tJGm1Exb/wy3maWySWpOT61d9hKj/j5j3U+FuLo+/Lu8TdjqCmz1TWDmTd
zBfxmj5X1JLhdTC9RVAYtESQrdUZM6GMdpzx8Xo4NV0uvnxaX5aG8qpx8+4ezl0j
AJfIjiz4EEkeFBw/DGjoUUe7r2Y0ADVcYaAy8rbSX6j4sDFRQXGG0UqwW+uRbXpF
MB1L9KM31IgDXClDNUJVVVI5HDfYKoRINzYyrNUiVDYLJkn2l5sevN4slUHosimF
3crtsemttInQ2NgcBdpIrNiLut90q71XbyvI2xDwKVwSKtdFN0+6B3MeDRJRe6H8
ujELp1b1no55+40+ADB1ybyS8sMjqzbVRX09fRc0Z+Kd2dW3WXB5Zcw8xIDq5jHQ
d/jpMiLWQuToRRKwbPmDHz7eFDz4BCakQGyVu7mu76kfn+8IlaS2J4/YEFmCKB/B
WcpLqk4f6jYWjK9cFWyIRJV1OnnAdzIBhXMjPDoxpPs1RJVs2BgFm/IMpHZaNtu5
0PMcAPQ/oQNGeeGRdthna3gYjxEUo7qWEeu+Y2tqCsmlPcpKdVUW5c0ADbCLeoMU
Y6swTnfII76U5ZL7Pb/mc7L3YLsPKtjtsM3yc965Hwf2bg9L/2MMUl11g3FEaIPD
mxM8Q2RJbXy5yAhVfdL5h3fO9XJBPd3k+3czMa/Kicn46WUfe9tzr9hcbsInUh3h
sb4Mth5K/O6sGYbNIpW71zwN8BQcChks1YmwwR1VZNG3j/8Fe8w4fhG9ZzarU04F
ZYTCFmQotGkbCh58Pinzu8f7CnpeBXjZUmtrCrD3m1B9pBeERvX/AC+p+Hdqap3+
OE6SWcHyl4dlEC9qTtYgyjNhZrxUmgfB6M+dV56ckLZFgmKqytOyCqpY56YXXDG7
lZgXnHSwAYRt7COrloQa9rNBpSD9zJOEmOukpTatL+t88fvzhCT3Ocdcvr00qQgC
IyPJMjIOHFVm/2zMW+ZnN3K1dj5+6GHu2emOoDg+74VCvtAxu9fGGfb0WRTfVwq4
1DvUclpolaEInqa28ceOcePbsDfMjdlLGT5IICzeq3xYxt/4WmNP4CTl38tjR5gi
KmW0YWXhC6wDWT70B2Tf933jC1zA2hcrA+pfChm6IxnYqcnCE/rKPqhltpFxUCUm
lnC9JjM9g2esAh2AHPFnvJ4LRk6TQe+/RDNIpjMTC26rcuCgizrl0mbkwErsRzl5
4e3eyZqrIle9Zpracll29mpHCP9Z26vtp660YhdF9htmfsP1NYFavtrlhFmUb7ZA
otU5Q+gcqrBLQtHIDPdwhFRMBmKgdQxDzLaUKCl8aFdBWR5S2RTouNFbz2mwCQan
8mwxPoQVMoEiHA63kK4NBAP7oYVQboxHWqMMSMcJRkNdw+94kn7oQzav9LcgjkYs
7KscLeMoIeO55KLn7m2mU96w3FxefynddwM9x9W4yj1tqd78TU2+16rjRClpic0p
OTdKpgWQ245vzj1j5t0Hk/mZkGwAfcC/bgCreTe+CwVtkFAnLTpiet44eAH6OWwv
YOzT/brzatgAyBlUG7xhHrD9UDpZOG9/J7tgrmNHEbKKTRfjFpt/ni4pTvB1nycS
+IG0PWagVd42OgNe/tkoElc9buQ8WKJHdOV072mMAliLtFMJqUKbqIRhcrda1kAI
oG6WgkCs3h3jAfeoPWaP3LtEbnyyQYVJs/nIKB4nX9QDIjf9d5hv9prHn4CC5li9
kkrSkUC06/nK4H8iYbDEdM3RsXZdgD+eB9WYL/kZKX4UuXwK/mvuXj5SMYpbENbk
X7Qtg9q1msgYs4voRYRCrqFp36ob71rI65MyJydquUBYwTJ+3Rdcf1DHvbzNiCOt
A7Q+AfEjb/VVit43haLbny8/4laZPDzl1ZF8Kwu2koYIsG0gCkD4y5Mt7/O2binL
In9cwRNLphlWICkDhmDdQZv+XOZKfE1C8JMrUFDbKrxM9/nTi+qtN4q+Ij6cb4N5
L3SMfCKvm2q0IjHiHG+Y1DugiAv1f6pkpZ8Np0olkpJTKWKBf+OStRt4AJtdSm/h
Cf5eMU5KBxBwFWhyrClyycU61nCK8QNniHsc3UObKoKJKP0qgWolsITlt8lAgjby
/Artni0d4ObIlWpKmS+k6cIYtanQYaUxj4AIeUqoH9nx8nQa+CF7uuEz+w6zS/ue
GMvlxWd0MRPw1aRGetN7jKMpf6JsXAmIH4qTDBbuFRMpDkBHf3fx4+sOjuRuXVbz
zeKQUUX0kHMgX4GDvhFYQaNe+eGS7QjbsodjM6mWMONL3Jof4zgu/lElE0w7Zebo
f382+q6Iz+0Jbyw04nks1b+TsVaAS+dODpJZ5jV99fGamGw5pqwij/6Uj8oSRaay
kTiFO0t0tPAeBkNkYlfzx3EJOy+0p85Mg0FfwkPl+PGi8ja5iwhmHW6/zpz8teOg
/sSBdVF3xPY25r6RkQwzg2mYfQ0fFVtXI0JnpJuH73B3/QDWr3vXvTxNjqOC0eq8
na9kVT4/EJ+Cax18ad5dsBTW+I61lkwEJoFkPodANwi2esZ3iKYIT2hpqdreT6k7
/uoKLK0BnvbIWSXM3MkOUlQx984by8dgwSglwN9ghC1CD9GYIv2uJwe1imsKQI+y
oWbDar4VNrOMYRPvCSCYQro5wvvHXksVAgqn9LKT3s4c11Jq9ZWBC1SsnYs0s5qb
LiNW+VGEFPEWz83NNOgb9T/O5m5yFjCaXMs7zHg4or7rdQIIgqFAUvdobwKgKzvK
8oz42O1+XYzMNx+5yatDsLt5krIbejFGOUHl9MkiQ5NoPcSxqry65cGUyjsiJVWA
XibInVE7c0IR89nbZi8eRI6H8lADe/kMhsqzyPi8A2Ug0WuDxyZFUXKfH8Ozfteq
TeEi0v/0YjTyuUbodRPZAdK+gJ8a96hrx35YyYiGTHMXjmEor7VPW3A05pI7K9y9
DCSsSdL4pH4epo8wgp+GepH4MATCCwBdujnOmFdamZqRGWXql9KRg2bEpvg8AA0t
y1irQ7FxYPG6cL2coyh4bhX6sqelsnMq3hw6dBj/lz7/a3YdyELVSoHr2ExN2cE8
dmFH8oxbOQ4G2jAulYkgDiMGy29RV5+aZGIzGm9h9JeVbnA460bCmTFxnz+f7KJs
FFRLVpsN/d+Uq6HWNg8nQT273mkiDStXkJ4+YpG6vdPGYv1GTu56S1Mgw8UuQhdB
Q1ee8W6z9jtcqPXPLx7kH73Gs+G1gGERhNNh2KDtveyy+2R77xzS3epSpGExe21K
uKWqHT2cdhrRmvXl6LvfGd5/6K1zqRN85+XC6c+xwzj2NNOgHztZJFraNMCYJkhd
OrXK8JZD1P/YbZhLk0AxVPrpdvX72ewErqmhbBuzjR09C2M6R3LaL7I5ceXuG6l+
HcXh0O+UX8efNfBMnoSQ15KJstr7Ojc0F9U1LvY9pNpd0B9OJAP0dFoNKuQBlGzO
ewb0h1GXVNYJPWlLqjtZOGaTVci28ZJi0+22sb/ZL+oGFv43UpKcLcYXPIJlUT0R
3zCIznw1vDceaCGDDYBYwpGlOG3RvAo5CHYKEmtZLwZ0DOmJpbUNYcIZad1n7Q4l
czFiF7wElqT++/SWGI32YbdRJnJeM54IOWsK4Z9AtioIouOuteC0nUJ+3R5suVGW
rPjT52P3h3Bzc8mDdMbKr4Q6FlS8xLiQV7FJYgx4Q4EJpJQfgDnxT4kc4rGtajZ4
p9RkcMbq1EV72kjuJpzQwN8mJF0/zY1gCEZRPtgnDGRA35GLRKNnGseYFCvJVVGH
QCqyN7P6JUby8jt376NGhnD1pD2MwEel2tXAApL/o0xPq3+KpQV6GAZf/kKmDhOU
MAqW5GBS6DBpAVQmoJPh6K82toOxCpC78dgYz5ZT2TJoSfRmMiOIy/qDKuTTK6AU
ntxTMjqu8wVvEWDeBKBPe9RBFa2NRIhiPGgjN7siHxstg0fKb84wdRzXn5/wjRzf
MFi0WSU8zNc/yAT1cNhtOIBDVGePSQbSgJKtVWPud+KaXTHE5cfjAwy/wwmG2H2j
XA8uqBebx2p7oaInbFeRKscVi2TuZcaPtOV+rUfyHTJKdFLYnrjIwfnCtYNPjVn6
Q+LRkFU7KVSUpZd+rxiIO9c7K5QgPzVsfZ+3wg+OffGUuPgFw7bCwLP1TvdlRYXx
Rgh9Z+eguYHrrOx7HqGvGVOPnKxocxmwsoURYPF6QVtFepCsqqzreEMPaFkSU/uZ
TBHzdfRHcs/M30HMhJQ1/84J2ec0XK92gx+LfLGaiTcgyzGoRDxvlxevXNWh8VvH
n01Cvm9cHRgZRX23xgcRD0W/TpGM7bM593vYXcqTn0KZ/OKOOOUUEmpU9XT1QtP5
s0Q/M2HWBFuy+38VkN6Ev/Nqd6pzEAAcWw0mOlUJ0wQE/BtHOBhs73cQBhrA/WUc
ZpVP6n+uHyjhrdOnvkxfWJMGq4cgCbpCYROgAjgbTCSgJMnCEt65xT+fNWMwLN5N
czKaMu4/dULKAJbiPk63YgXOnVz4OGbmq039o+L+YyPkU3+FcJEeNBGCLgfo8v3n
WX+LwsNT/txfviN0/o6ag5ACmR7vkr5E+Qc5EOl3JZngAjRRds9kXRbXT9EMTHQO
1TIDVv1DKwH2Dx+FcLvWmaXNJ13+Y8Mu/CxXwPzaa5TB5aFactJmKIReEnNxnTHB
bYGCyp6KmTYk2PUrvokLjbGTbwFl9s+mDx1LgZj6PUIuSryQFN+aAhj9XjGhCHNK
R2j1cOpo5B/maNupGphhH/8e8GG3Fbxr2Bb7E8j9yFarakpOvkdA1wxr5BGLtDgi
wHGzYm84nPyhyXe3lkhgL6muMa5sFQ/Ohierxfp54ELPRu3ajDZ7G/xZhEPfy633
jUhAUqtVH46nDj4nCB1NqRvHKUg/m4vGxEeD+/909kA3JyiXV4KuyJGf34uJr9gx
4IISLqgRybf1DRHiZ60zApk92L8p8crrkjaLeeEcrrTVyu1Es/GM7szWo5iVHZnc
Uqj7MSBBr0dF887eryHuyS1kEhcPbIWxmb3YGFKx6ComdR+Je7tfdJfMHr+72ryk
raFCgJvTMw/mDGRSGWEjXPaDeSbmjyYq8hcQIes6vGdZcz+Tjfq+69II1H1iRAyz
e2URAtxOxLOy3lcdpxCuZtyI5zEmC/ht78ir4Ko0IIweoFHyueG9kXnF5R0CA8+p
MeH56UsMkVCZroCmvK4bYxGa3mgCgX2AN4Eb2HJGRWHXbz4Ox4ZAUrvxlVxUPJcM
GHjqsGSHyEtXxcLJJ5tLB7ThElzN3LJINeauXy373ScxIsnTDj/6mnS4JAKRhPWC
xXOafGM8UUaCN1fYPy2HpBgLSb02/eVKe39BBUdQjjPUxjqa+M8+WmYn7Os7nGub
PCq6c080pSEQkS4I5gsZWcDArMIrDDyuVIZ4nfGgEG9ETcOpqcGze49GkkxaLcx+
MSgSxoB9lsdcdnZaClgtegb+K751PaGh6+ak/2RQ2PU96n6DonVBhGAiK54jdAtB
0e2zqZGn0ishAEyjyn2pivw6t3ZeT8L3idt2JY4WIFEZ3ZQuuY4wst/Kygdw9Mad
Dm4998gnpAwkPtkBoJ+OHAcN2tiudea3T71DtypBCLwY/ICMNd/oyx5oRzWWMdp+
lgLQKhyPiPQjnIFOFIcRU+aarl/r0FNt1yGapBI/PjUeK/T6mpB5LB+gbIVrUWK/
0kE/CTL0qtrTqdTpTmuWV4X0JvVfq1ua1jQqSLHI5tXSI9yM96Iz77OD1cELRC3Y
BgLFKZ3feA1why0o9NT8Oo25zSa273ULMUD7mmEHzO+J3GcbiGjq4xjeZfr4vlfF
S7ebng7eawGKjQfCmHh29cnC+PB42rCjEiYAvytNP8EO/NmJcFG533MLT6UIZWwF
7H9iYA/cLoxlakHzWh1/Zz/HU9pIlkRXHs4AxtjlbkaiPrpnHXhmGYpfljtwX/q2
5NOwqMK62PhbkuKhM5SY9AXyaJZyopaxPpNuccMUfdf3NFpWwpIhksXyqH/OEZRj
VNd+gNPXtcVNvQuASybl/U5IQPnFVfr4jZDIknaoRZyRyXQNy8XpTlWGXfs6MWN6
lKFdLB1noL0pWQq56c9xGpBpt5cd663tHml2eGGvOB0zWr36Hk+bFqPMQJ/2WVC1
5uWfCYjYakJpbryZF7JoET2KOkzyfee8Q0cjl4HyBU7QdOJbM0IE5x3JEGfhSp8/
mW+g2OzWWB5PEaoLy5kFd/aNXmegQ7rGenVlEsYDQhxHOkTsDXkJw2QUpqXooKk6
NS190twZ+l+KkoM1QBfyy1qsgaOb9kmpqDDcF8g7wkoQKYCrAdhqxp9nqKKcSSAN
3M3rwHSF+MSdDp1tXzUeP8skpML6xjW/7SP+dlPqBwdKq6xfOSQHBjiFI6zPO4OK
0Oq3lbRIdBJPKtmPDiu8mp6men4EiC83K7W+fhfWSe1qVjBpiXr9DuEJ6CkzYhXm
cZDK+kaoPHCa+YpY6avjBrvO7YVMyTpaLpxb1TS/HeEr/mDIQwCscJd3DuNn703f
5U0pu9gzyTb7WzbXTspbsls5K5Ka3XNu4SoXv1kJWkDblQ73t0N9ac0ewZ68VAgN
R7pe6n+M6i0X8fh5zwG9Y6n6y1wY3Xmmhx1wbuwzmaT9ownzdLrZo79KZhkdY5Ej
u5V62c0VEgX/lZ2Vt2/siW66TJxZBfEdZ89hJjdQwxkWScNpMp3gaN0Y+stHst52
fnKVZDvCIrIEM/5cb2JhEaG9TqeaN6iF3bZPVLLwTvlmf+MWbsaDZKxmB0Yc8nhZ
n9EvDB9+RkcPb6LZ1sg+xznCBPkYUPN/0jhdVREAmQ+ozar6dWs4q93vvgPUHw9F
FpcGUkCB1z7iymTvRmr2QYyoWfhsL6bYrosC+vUKNGG6PlFd51BX+lE0Un2vHGFF
mkyEXA0CSoZdzMGz+eeDPTndToQTxgBxvDe07RZ0gNZW3oFYpbTjs/KVwNbHbROU
mtztpeLEmP0t3mkZxIjH3KKm6rB6fhnkb9pgdmXxIOKKDcUaE8UB0S7Uq+gyHvno
LaxKO1S+efQAgsDpdEiqrNnzdbzgWoJinkEoexQhajbe4Lrfwo04y4d1PuFoi514
bMmUllKEgG+GO5SnTLFmR2si5hKjudTklrWQN2srxP2WptZ1+Ub/dd5CHkl8ITfR
wP+3xWAzU/B2/NOx2AUJVTYSJXvFkqlJyNFGpQXbw+NXRMRV2KvqX8UFiLAEnmcj
kztEUyMnrRX18I+qrusIJsmV8tBlsx03+LCYcU3hvNmFKT01/s51eBYTyHVzWt82
d48kFJ/XEJ+YClxhh1cLw8TVzIw7hd6KFEHQs619XfHhvqu67PG/jYt+Bmb1woZ0
8S5gxHtViZzVYPhAwDMg2uFwAvS/4c2FwAH6u0ruSZrPcfUbJ7TGAMAqsCL+f1xr
2XwrEC089ipRbH1yqo6xPPk0YB+hrgf0L87CNh6mC7t52Sl8gT/9D4xmdqXKH5bR
XS0FfXwfiK+uf3Hjrf2Dd+TjQMYNch9VMGGBRhMuSbcw8rXCTOm0VWiIV4l2mEaA
6msnqAGLXASH6ZxQuyKnWq7u9YnY4CX4EHRS5dDzHHJeqaFmao5JG85/HaG3Ls3F
rg5dF101T9ZaTYDuNuGKb/E7/2dmocE/ChmFTmfdelWgWipAjkuUFciIUoCj1E3/
x/xhJLIpuFVwcav/l1sL01gyf9TcjBIIiak6j6MNIZ//4aklI2LAOjza6lfPYFwE
oGT2jy0Q/2IbxwZ7sprVSXYhLnqDGGVsqohvc63Mvy54m31ANBMYsHf1rZ1JQKAb
KvM8h3fPMZqtnCXsCk9qgrA9NKChmzMb98QrTfDDR6HpKpi2RArPnEFWjLDN2i3Y
555l0tdUoa/3rcNw0vfvZcMFoRHN6mYy+vcmxTOEij6mrTAxnIfb8TFRuYBI5Ine
8XbQbu0fngKxrgkQJTMoC29NALOpugzc93N843X4yWEjKob3lqKxMmbj7mPNEnO+
JPKu/8gUkSzmuLDNAi+Vk6lfuedHWb2yh7VLax5LD9CS2LtkQh/DjAa+h3vYUnkM
vsukAlNZlVA9J2A5B/+INnmifBmpZX5ZYJLladdaVaxTnDDjY2GHO48MEtVHM7Ih
N3CsgLAG8WSD5vbZ+oX7a1dROTc711nL+QqmVz+2S0oqlzwGbA7IgyWJbVPNRNMv
WL/4q5hD4CK3W4wY8bzowhdyCzyeurUgFq6+98f1wz8ngO9il+tqn6dCIwbyh8mV
ZwBGRsmqbAMG0oBmhqyLYo/EZwNvMj04uL3avfjNtifllmawiUeQsXIlFgWrS+wo
q9yOrtGW2uD0X1CjJZLZshG/S+3UhvrTy5cNAyUUjpqf2FOZB0NdQPCSMrCNhEfu
vIZV53gFHftmIppOrdenOE7C6E51ME3RXvSlYY+uPnUfKoDn2FLyoyv9p6fYowpa
cSRugq3bTwYVm/Qu14Kr0HJ56ckhtJzNxyVeSZeNvcRZE/uloeKyI/x/btvwFN8Q
Yh4sT42f2dRzYCR67Rx+OvooHaY2shQoCc2arHq5vUrUYhyk6V1FJ6hs+hdgWPFr
28LmZDADALLUOIjhxF1fi5hR6Ff+oaQjO2cFEX3pjXP2QCV+r1+ugDPr0WE75Tzg
Lhb+po5ktpGp+EZnhyuqHS+ddAtxcPYji/RS9S6vHYglVyONmmD+F+V7v04zkGS4
FmsbRHVPvqAvop4yRpPuhCCwM6nLhm9/mai7KiCTCeDd3cNwjrWh+4V6FrC8o9fz
J0pkAd4slL6FgXOsJ1UGVEWUm7QAEf6CcIQCrqLoFRcylwj/wITdAHzKyR6EXRAg
rspxcV/+qcWsPUWnPXCmGt5i4HOeLnYtwS64WUKdt0SHpvFZbg96Gw5XpsvmG9Gu
fcfkvzeunFz/imMbDlRcp+AqMVGnxHNVMq7wgoEkMVWTGMg+NPir/O9GJxjSgZBx
mmpO1yT5unog6N1B85IQvsGRHmpkjNpi/j3cHknA70H14W5vBR5GIf69zZCggr32
GPENkAO7187lYqZwFiyNVQeBhqkOyWy2ACTlYf9NNPy2pidvgod7d8l3IA518KDg
lvVjHeH5OK0Ydlbgxdzp7Aayogh8RaQvYRXcxBy6ISEsrMoD9DpZNLmbkyBf+nOt
Nd/B89SpL0LRhckpiwcgTNj4Eh9UyECvdirxym9+i9SSFr4H8FNLrx4y14JsS18c
4YTxdSUhS/pPQMVoH70TShCqL7KyjksiNpM+KAfAi09AVMUshp0aRfmyUWED1Mnr
qDbR6gELV1Sn9hIOCjwgIYGnCuA8hHw7aqnBmHdljdHtDI3htjUnkxq4Eae5tWHl
AAdDwuLgbIKsJtToyE3XUSw0IAgntJBN5ZFfaJxES0FNFI4N87rpIwIomcXrGKDm
VumP5ZaMDHn1Kh3heHCfFk7G4qZB7UXyelGQL+JmcK5xiY+uC5lKYkK16xsNfEAl
oadCZeDPcr+ReaiwNrzJa4TI95zUT1CPhc6XhVIaAlxOJJTc9A97YxbZk6aJD67A
d4xJT70kmruz/Jgsa4ZGRMutFhqtItHWqooTvPL2vZJlNGcRs81EWZhSvTSJOc2D
ZdfJCh/lr3QYfpcezcpbvVc/q4DXOA8J3ul6ilerkAwyI+bZkYi374LdVnnugGbV
7vLXf1M73W0e715MiPynUPIxdAbJbmo+v2o1KS8nl/BkVFXvIVyPvXIN+rpK6dy/
zUi8TKfVwwS1g8fp5g5V1SBOZ4BS4uwaWoksNlakL2DbXq6mnkTdvO9Dtb83mouQ
oD3wV5gnmdmElkqcXnQLaP+C3LdoV5yVZ0JYNWQNe1AF9pKfhcuorN7TMHGz9D6v
eFMAiqiwbGCPmd0WnYE4bH7zvlLhVym5lD6u/epIjMcICh1dd/eI7TR59CZdc4I1
lnWoGn8lzmNjYQBhjJCmYJgQNHcpsLBwBoT3Z5qgo1tNgR4KC+ZOoO3YvNad5t2Q
qRknxUdefgpcfIz++TGHbZzCuu1aKynA1uiKlePu28r2N5V1l0fSd4suMTIAqp9o
pwYDd+Ix00fBgGPb8CAMIC6TCpsSja4oiYLLHGDWfubCuPNlKwYXOhdqeT/N30v+
yP181SbI6U5fMUvdKMlAscHWdamgyYMJe+ZWi4toMGg5Mlbn8N2P8t7D0MDSTvaj
J/5ZyiLq/xvouWEuvD1cX24hzgenxACJCtVGqvbW9ZGfp8BiflVJxAEruHHZGgks
xcm+YsvBTczzTktPutzMV2M0208ksjVSclmquTmbHKtdF9wKwRHLr+vfiSnsiNt9
fkFIKpfzSTlHNkZM3twJhkK/sjI98YHWLDm/pVnm//14QivepcXGBMXDKYApE8FI
21HJ0ERpVqlcdD4tP5bnNfWk6jzHLDRrf+mEzrKh3mhGzD5eUubvwhMJHxa0HhIE
JLvwe2cnBGURWH6GDJZFEhsPdizF5iz6JOQ8+xIM8ulxf+NS47h9Fq8LsgA7HgIv
i+q1evNhZ8/oNd5/JgOnL0MVXECye1PkD+DCrIW/NxWH7kvyboSVpcmMm4fpJhmt
BZmhJGLMY7IabKN3G9YSVNs9uNbMaF0B8T/+yVQCT8QtC1jxEiunHZj8Pz6OVELt
FHAYHgZuj/Gx+JaYLgZ+D0l8/DcAyqQ7It3s9PazQCXZBFukFKMNcdgOdhEkNWTp
Kqj8Lex3/wzw3VvWiVGKXVmva/GmE926qsxFS1p5WhESyOoDi6MnI7PFmu4Q6Dgy
zjCFLf302siMs6DPaIyMxjYLWjVix0sOII3RxPjC8ya0upnsxyGqD/tu+j3RH5h5
GoVmkn+vVlHVjds5ShKtUQzySL4kruo8UmXH76KCOBxPZtq1YsLq24prhDvo3SM4
LFQtW2/68fO1n+a9u0BG0xjnwgavrp4vKb0zPaHPZUtZOGeVUL6i1GMvjIv8UHS6
6+nqm2hpqcHnjKk6hm/r/wSWd+BG0OwXcHUuABdH0K58EsiuiSC8WcfdjLgu5Err
CuSdIOL7cQqdTv5jcJUgZLZ3NsC0S9cJFA351Zb0VQ69dx4KgokyNZf0fPgTF2CE
EOyBFzvOfzEPgQYGazNygfvHLbHdtuUvXJ/8jzITgFqfNw+joR1ntpzG3EbLNq/T
9OBdN9QRpmCLffbfGaggaqmu6IkjatLpl4mtxlOMVrkEJWHY+hcK7sOqo2ulRVIi
5Fz8OZHIqf/sZWVvKsdTV4ZumQFaY3yuXC+LeaDdOy0ZKDb2ZJ1zZ+WoNJ3SPorv
VLCz8lxgdBF9JDqG4WZ2+LUaG/yAUUibAyN+aqrkqQM2iSvz+kTWwmIOmzggG5bN
wi4Z6auDOaA2kEoA1Bw3cqgZpWk9gkY6BJwbgtHI2Tt4q4/rmt9ELKdQeDiSR65q
Fep235L6ylvhYWiG7vfoOxjgc0MVLg7HbwW2AMJODTBkRQhY2pTBhdL+gi3zVH/R
fADFsZwCvFXIlv21Z2u9Chc+aLmOeYAgh51xCxXR8yUoHgXgXHCxomDZva5z06cQ
/g4akldDRXjbhrgGnwMLNRBG1/KQZjf7h1nTCMBkpmfgW/W3Qo4Yhp94rIPO/KxL
CoWPabg2+6tRLEEi9TTkvLU+TuEbvjUNuf0JMaXgJK5kedORVRBoGg8LMxItKrZT
FyQsr8eANGt2+6wz1kjY1X5A0fHTES/3qZ1+Np5s1QLrJoNpQ4HoEHr5wCn0Cjqv
aEgl68JWx5GRm9AINTuxqrgHSzcmHIPHZ3/4utXO704IwySyp5QXZ+VtWOtBNVvL
RsND5Wb6u0PPveNDuIRObHQORbThnajOetKvrjGtd964LbcaUrQcGNdiZLls9G3S
UuWJ4pADyg4P+XsIqsu1nTx2djSqp3xPjgDFwNcJdkE/QWqVbyZiDDhcpSuLtRn2
o2EVqRFAtH2HeYQALpcWxpaPKURoua56m+XHFMj+VOvAzJeu76azNScSX0AnDYF+
6Kcfkmppu/7Gv9TmTIhS0XlAFcKsPDSi84+K96ZXWiQGiqDsLQ9RW36j8AxKQJyP
mwWgi7PpAR0SeHJA5zv413QndRtBcfPW1afrF2DILuiMwBJQd5rwf8CgTQFWfvm7
E2sZOzwrXRzQFAhYAPIUw0gbg28DKe1b+SomX1M+3SeXPq4QQ8H4WftjpkCUPvyc
dSXW6K9EHOlPTa1cTO1c7k5beQuuK77w0eZWdTtSyP63E2IqLu+3paVi5LrhALqR
a3iq/Grlg9WRYEh9ATemjMlL/FDtGv6fnkHt/dJA8/BsJQ4fIgJUlXNZFF+jRokB
6usWn69bp5bILT0f4xQXRiTCF+Ep8VarU/XnZPNLAmKeERFhZpuYIJtRSXK15fF/
PGD7xdbF7SktTw6LHPUe7n6r3DtwCoYMdzTYZiv0wcPtX+VPmyKfKnComWQQ/4+O
ghyRfNnPm1/AVb9+7zcN6r9rAlOpt44vi+ZO3lsYMAVbVNgkrXZR5Pu4l11NkFGM
2hn7pKZhQ1EUBpkYWPTBNkxB5bl7MngYUh3+X+oqMXxISG50580ygBdX/vXI9g3y
Taf11eOljdVDc7ebIJA2HrsOBH5OMasogxVS7JRe0QZnLmXSXd59RHVfP896RGwt
1HstA9enZoG8iYW2EzhPh5r/l+r3pxjG9HTvaxWyVf3eEalP1QSMtU01ykq992DB
wtkJreT4HIFd4aNdFeRg8QLBlngsA+dU61AhXJ8f6Ed6z7YFjWfcqa2822JlhS7e
LGsg5TV7lPBp2GFL7rUIPsP1jUD5cZNemsqiDtUD5bLOLWz53QNusWVke3Fr6jne
0wiIMJDSp20HTmd3SUVDlX8MOfdTRzWulH7kgrIMFGorAoXXa102FdCpQI/lpOTA
yFM2sfZX3yu3CiZzF5fSQZ3uOaQgsqfyQy2pET7xMtqvI9UAaRsFdfFBzbpPsK5p
l5PFFEg6vVsMQgb8cXM7Y7DfvBecL/cikS0qCqVDATeVb4eu6iGj79mL0+uReQed
s7T7QXRTtp0XHvTU4gcQmAhVyPKtnRLdPCq1LuVIx0dlflm9L0qCjMZNLzr1txSx
z00OGP7OoT46hjAHRoFEGBE2qsJWJc046ioTMC75f9WxjBo0G4vbzX5Icpnp2bbs
P0GteEttkmsUQvGeFtmwadoOn6F5RY6BrCAEl8ZHUkValZZu95dmKy3YIOkLh/4l
CSMgmiCKqdaQP2acuO6v9I+O322bViKQOtYDZpAbR9UYLWQ4YPGzkxNulTnEVVMy
b9VDZcLDRKUbKnRcq8b4VIa7vgAtZspqeuRw/1LARZgpmeGVh2MulfHlxiGboKGd
uQC1fWHGD7ajK7mBOelg9WMzSoQ10poWqZ6gBQATyWGFTfKRH12bRLA7XUS+EEud
kM+P6B+wSakJq6WBNnc/nFMFNHuiPsMIskbS2kQkWHl4C32247QP9ExYGGMNuX7M
x3/braftf2cbXOo2XUTwkpOB0PQm4M5J4A+WJoV4aJ1oxTidQFjeIP7xTgbKnOdv
icxRuszdo00AZCimka1I/W0wGt7n4lnM9t6jL0pCwLjQB3YC38GeNH4M7xsZgqBV
wmc6aXLr55s5cFAnkBy5y+m4h0Msqa9E5JIjv58adA/PP+2q+sPcfZQOioh+dDFN
lZ+SUEZ+guKFl/nViW9urpQn6xiDKyfuqnQbhwQh8aVZL3Mvm8c3KauEZ6dIT8vQ
XTK7RsitQifvBP+wkS9SiDKcHnv5xtObM9QkFQzgXLYnAzvUiEJrwTimbU+ZVrm5
AnJhlNYAwzNzU/rHiNMtPf9qivd0xZpTjovcSlJLUt2XtWP2JZQrDj3tCRnlQ8NP
K1RnXOlkYu/49ZEWnKXgGrJ/ELwXw107Isg26VhZGYgwZAsCeWhKpPcJu/83Gadp
8iWEiwM+SpVu+nWSi1xEUI8FcID7c36T6cdsQkZRzH+c2dXm+pPHJ9wTWYhS68bx
2/+5OotdOTUs8cT0PX1E1BY2PtKkPlLx7e5GDNwij9xk+YRtip4rmc5+cuEa44c1
I9KxpIQSEYh3MC4sjwfZYmztJ+O11hwjPaxS8OjYmhUJ+JR3EfJF/mU8S63nyjcM
hJO84rhOewjI+hK/2cc12COBkWxJLdQxR/tuzV/BmlifBqKK+rrZGwGLp0UiuOju
Q/USGCBC1zZUCUAzkGb1Opd81JCPKDJFwBf0zP2FbtoB5Sw6QpAlOg7RuG5MuRl9
cpgT/zlwy3vgJl6OkZbWae8loXyaQ5bUnVRFMWLB2jcDEJCztMY4ol6ufJZXoeaf
vgzwx5jR15YL2BBdotRy/Luam4QHVeC0bxYHSivwdNPAb0zGZHsS71XFVhrP3X55
fpvgVs2zrIr0uIV+VTDULlKzoLMz87QtEfgK8ihx1rGOpY4f51rgDJ03P46WnaCE
nmhk+GuPLHIuN7OLZ8wPXrSdHVLkPlGfTUnXFlkIfyQCfi5NoBGQubwIHy8uP+QO
7lTr/xiffYx+DZvDeC9wd1MsSCIEzwvFBL1ZijiyiNZ7P9ULmGMOfVanJhs5gxOl
hpO26KvKaalQvSp+cwQgXzqHMVK6qQ2bSsBEaEekrX45j4x1MrrwiJZy+kX/iITK
PfNfMc6+TBenwX/5L7nCS5QmBBFY4I9ru9OMGLapRE9pYy9KbhhJgLUhc+S+84Pu
cMQHKaHOaZsgUtmRIBOS2iGhQw0+GWlDJ+Bo/sNWR6iwvrYUhtCmdy9xYID0I66N
GJFjPVmJsDs8hnSJ7XsYPQH7n48Gxu+HafDi3UG1kbn2f9zGqS68ReEa1Iux321N
huOxmkrlPk8xG4I62DU6nU5OGxTY9arfFYVorkqydiBxLzKUeg5uUUkNnA8N7Fpq
GnOUjsC4SbyXsneYiihIwHhVM9IhYPBEjERdQ85EB4PD1PSvCTcbi424tUqAJHw1
Db1VSq1rZHy4Ji7leRz5Q4AyxbEW6+uiBj8kta+jss7PYkwoQXXDXK6/xZGNdOPq
5bS3meNfTM54hwKnA6rZ/CXrd0ws/LMEUMkvlvtdrVqkQoOeU18WCoejxfUvAqD4
2rz1VJhP+vmIgCZlyxbakNEqk4jDjRiuYkUz3v3I8LJQLCWjULsAjCOO+d3/8bc2
4V5qTRb83Lc+YB4xJWjX7128K9D7m8Vh0spZNvQe8D/ADZfz4xZjihrJbzGibz24
aW7lyk3EXgHQyG49rSODva7wwDppvHHv97qeYRG43kzwlp9bFmpgeORTG9QK8o0y
rmVGJjJl6CpCdGcUNeLb99rAphzEeIxP9yQHAUhmDUsoEV0MaAjuCpWoQpUL+2FY
V6dmV+BjD3DX5xDy/C3VmbxDW9KIpZAbySsV02RWaKTO16iGbxnnJfRIvNvT3FeD
8HLPaIpq+Cc4gkyFTYd4CjgoQBRKtn9Ou7nYdNdkNu5bWhoBecI2oOx+ohumiCq1
+olcyypijV8vL4nsAzQoPViB9FC9jBtKwTBBxX+nlY/FkRqNHJ6FMx1DafdnpnT8
T0Z6AFYWOD+OHHExCD1zUhFM54V2Lrf5Cph0b4c03UMwG32jAPgK3NSQ5hJBGSb9
rcL1ZbwJmuYBwgHiKNjNXvrCq/Rfqq2SkSdTatO/o6Ozha37fFhXQdDBEuXObSHX
KjamZVQdzK+hmO49GV4oKVDRV0iiH7pAmsLrP4ljroXHzt1W5jbXQ9XbjI9zT7iZ
gDEMMJ0s9NuDXLi0d9a9nyzQvXu51bOHpA9ObAaZ5rCtWlB+8RGoZrNr7D/5TAP6
19HTHe8bw8uvmCEkdTG2m6C3DmKAHkMjz/3RCKNk4X7xC/ZwMePVoWXDzGx2S78A
8InAOcaMzckVtYoRK6+3D3KU+oerRnpmMkIDJKbCVYEjTZz0v6oVQKLsw6eM7UBv
/ufCphpcSiG1//2gtYRXFVfMWfL5cj/02BzQWMTWxcgOzqAeBxV8GEtGMAeMcts/
BYfdddprmw46F5JFHYFJ6OSPV3jkH2DYlQ2ZpME5N7BlKMiG4/ujTML2q/n6G4sj
3G5HlfQLsCuUtutGJQ/TynKWF2ecGfMRePGRShe4InopWnGs1CI3LfaobWHbmkRl
rAneHLKiiH2IE7vvukwR5njtAHnIjavUjolPWBS9HJ8k7h83GG4PfNA5jJzW91RU
gOFbWDpUdu8AhwSV2tkk2BGTf8TEBSfNJoHhGfrQIE5U2Jq1TO0IsW3vC7SdEoAP
WzzXyZCpJC77wyjx7v0BkJcD9N+unKE0fyek6toh5DPaTX91kW7oIFoFw3Zet037
Qk1sJvm9wmWRPrSuqa29x7G93eeCmy+09OHyo1jzGItBe8H+tAMxo2FPKkI561Jp
lxiW1MeaUY6ElhOP8WwDvcwQkoA94VfEjiqv9c37qe1GZkCY3t0OW0OjyVewqshl
CE2w7V8Hptk7y7C8GQvSI5pNdXTyb7q5hvxI6Fl/kXh8MrDtBCtg1cBknmP65ehr
KUGutG5RpyN+LedkX/fkrGAfOtBEiNK24vHjXYahBG5rKRdTIOKpZwglU3gw8bM7
5IwAMhFPvZhL5x4H/Zjrr/wkA2RixqU8qF9PrxpxnJr5eveOe/Z/QW8SlH3+1C6A
uu7Hm9luTbBo097SlrSuN16jKv5W3h1ms+wTMiQ/6F3ApqsrzYWWrJhO+DCwX334
DobGGjSH6xMhF+qi1+u/6dTqmsRaUGXCGxW8DOIjhWRDABCbMGPsBzuF7vMWHqZ+
tm4sfB6rsJ5AfgjRX8Tbu7Ii/W9NE35tb6M7yNZ4G51+QIS6x0BCSrZqfRDyklb9
IUe/AlLZILjOcZGGdW+J/+RirK/8xL5Yii/a5sfa2njdcFQTDop/GrqQWaDWc1bY
AdzcFKtYzd9D5LyhzCZ4fRoNtwl84sDvKySB/fj8jnFydtMeU5Jug/Q7BrT03Uw+
UBmSYvTe47+C7h7C6al0Tq6HlKuQY1Gvt5WQZVJOB0fW9NIUjy8InliWw+jRV08R
1HBGf/MYUG5tZ053ByQdiZgXAX4FBYvKh3F7m9RCGelazqZz6ejxZNEZCEYqhM9v
GJVBE2ie4eq9eR7KDd7GhERCY/vqCuGobOUiQGwvHH3HJmhIBgHmm6mKtP0rYcS8
cxm3AIE5evMoBbIJFTkk/0ia5fFZmDdAfrBJ1tOgDb3tedkwZtEKRpxRuUSb4X19
TdBl8/euQIUJHCq2fUNNLKGY6udtXQZ4UnIYN4/DB1fd1Zt1SJ5dgsx5dnSok3eF
akdPLesmYQjKWRL1AwYhR35AHdELqx/O2XBqGoEcrti4wOavMOey82MD7K/g/4Ez
s6+SX+SR1xuDAXnMXQcvOCYKtvQmHFa4z070wX2ErTG33JFs5kYla/zyPXGLSd1r
tVqSvV6jDCWEFL4rn3XZMUYSRitEANup7122nZaj0aZypO74qXfTssiYEw3FZ6VE
JsfPB9Q1cao6rpcdN7yF+4mLmomXtYsNJyRRJecGyZZhr0snqk8Tw2zsdD09YS0I
dkGSGuHt8mMDXQXPTOjSp/hxGF7r8MPza4K96tVMnad7JRl2TeLM68z7zrhkZX5C
chhSWaof7PSCkucL00NFljUxpuQRvR8EDlt0dMDc/m1cK0S3TBbN5SZEJ7Kg6Rye
ibkUbxNT7E+WM9Gj48VL0Uw7j32ywtY2EOj5jAs40vOzHbvC9kHjtHlYw0nnaokR
Lq3o5GmKuZ9jgRanY0rcrrNSQFK1Lguh3JJlMshZdmU71iAwuts/KqM+hQQGsQwl
BC5YnkB7zXEt90rxQ6AiDwDw40H+4PtZ0Zzfyf9K7Oe1pYKUbg6A2FhRsT4zjpMN
EOAy9nVSfpCtwbw71UaB6ZofUNBP5DgR7G38P3gtuEZxQoEEnNFANWalV4cDTkPo
GcoYMsTuW9fwfukBD6YHxwZMzMRBb9QhUYI/tzFvKbKJC9QaSrEJOz0ynLInXRmL
Vqd7pSIqua0/CzSPKMJbzMXZmgszmqBq7rYe+P5owCeyyfLhw7jrKC/MYJx+/4Xs
L1/IDrbuZqkEILjX7oPd5qnERum+ekdLQL4uEX6W03P+xsyjTfppxZ+/jct+ByUO
+g1jlSwqWc5VdUw/hTf6uqlQyZ8R2duvl7G9bjqk0wdkq+gdC8yoFRHuYu0ibK/p
EqFJZkPWXIku5wI50GOBizSSaii1WZ90gTQunCzXB9semXnvFtUL/KWVq3HxvFxF
Jg7iLCGX1wRbCm0RFZmEYxsrchfnwvR33llbiZIR9zYuA/Y+ymKneASW8IsLyEGc
AaKOCLT5JQBaR4yEqkuabex5O9br48I9i7vbsqC1V/40Xu1lRzgeRm7sEjnIbxvv
qLRN0roB4Cd0Sin1T3kxjeBI8MiuHktN1mVZoyQKOVnbPPLU1JKIP4WlKgSxpvXq
s4g/s40SZjjxNcwZZ7mLtmQoPDstGM3KtIyIdIAvVI3PQXDtwLBfvzuboH9xXpGC
uoMHPkGyQUZxHO7t3/5QefftSHI9yXpTrbqjJ2LUVdJE6W1NAjFx0Gai5a7vhlru
w8f85VPR7RqE3YqsXNdDdBLN+mH0KVBXfz9zLF+CBrmpfPc9dOxkr5w5ratEpq4y
r4PHnj+Maw6F62Ow2TSxX614p/OFnnpUzA3qPyGUce2bUZVcafvOTKi1l9VFUE4v
t5EN34vgFCGqyukjXmw+r1dRAHsqJBpi1d7HLbehx6OHJWl1+HPXQjaPnaQsx+np
lSOb3t7A7BGY21jSYc5DCXdZjA+CIdFPvQDXLNRYFttoUrmfWV0/0AU0L4y9Fh2m
u9P+W9EvTSM6PsorOOFZJ57nuZedYuewJzkAHWdzQ5/qiGbadRCosFXccC7xGU9T
p8/sPxG5lBdU5Ecj20B1ZfY5Dp8+PT7+weL1OS493FBtLpr/vgRU3kzo0vRXf10g
0kxREcso+qaCQDz5UcWGFphUkrRiFoQJh7WireoO73WytdRxR75dm+gHae7HsEWV
whZurJI+cpcDn+xTxrmN1PDI9Ll+tyFcdkpahh48B/3Xk80i76NVe5S+RKnKdFPF
LIbT/fYeHA5iFANtlfb/u5JTF0E7IbDprWFrDp22xq7lWWJFbq7LNzbMgNQXR6Ye
7klJaEA/erubv1awe8ahIT08zmATlaW3rKO7uioDMS3ffWkjhz6Pkk1SUa0p+huG
FhtDMRp3qjd+3ALaYXu3vlm3+brgSCOAVF6rHPVatMKFY7icvk8ptJBK8jVbBs0u
86R6YTDl3LxHBZvKopQHhJ4+/M6ZY6NfROJFwZ86sTPTBx5A+kbXE5Y4O+7G2sK1
I9U+v9oDxNY7dIACME2BvaeTWc4jeLm6SqgZKij6pYDTpECRR8b8bLmb+DMWzVLD
zZ/ZzkAEY4fu3MtFcfXtmyDjCbUE3RfbmmvfENm8lwli/TT+G1WxecdXcxjB6tl1
pUYFERJe3cmCmPfNwQ1teaF7afhg6ThNXl8YZLqX6uUZZj/ityGk9HIq7Op4teL8
5FunE/UE30N4qTqFs2HKTKtk0cRJPGAOcchKctmU7EaIuWb0NiwZTJBjTPejrrH3
pU2FO8+RMcfYuhtb82Qx6bEtkP7YrIv9SpMBmXbBhG3VmI2s2vcWM7SqByHXgWb6
aAXkqzl/aVP2y6qqTe8Pr3qHwrKDDeMF1repoeg5UjGmk5BHMc6xWhEH/3mjY1MX
7QdSIwQW3IqFxr6fZGmXVJNmRp3SxAc/SV/Jv156RW30Aff8Y4VHMizx/+AyRA9i
rx89OQ6/PR9wO2oVMoWAhx2FEfYK7JMse6Q5yjUEZgQlNsod7dlVcPOIQQtq9Dck
oFbrpdc+5BhGVfeOVTS2BRJC289NAg+piEtWyNQA/dZUKQ7Sxqt/iMoV5dh4Q/hj
3rJ0EknpZE/ljOGIyvzVqpGwpXo0LRoifPw1rWurNgunhN+x/7dQjZMNxTn3cVUt
4l3Ri0R65eYyDmG7V1Xtxfk2mLNN1bHszVmCJCKUlN5jnilBeszKbuaA6ZU5YCtU
cIetnPKKhoCsocFYnibL19biMc8gd9G6v047Zsk81rmA51PbAdxyoh4jxSEM0bz4
e0AF477nEBcU1VEwjsEdns49fDg+QSCMplOviZyNjkiVaMH2RlnxQ8WeGTszRYlS
IrcbP7wSqi044TC/i8/eUALlva/5RWIttNg9LownnDbkpgX52QVCPl1BFJDdlBg7
Lk7G5PA5+U5jkHoHxbBA0Fi+NzwOUti5YzC4iY4S0EOn3P60HS62JbVWHMN6CUV6
myFj4Y0Knq3SOR9iV7Cl0t+jJMz9l5jyHYkcVFVAAdNh6UksNLhCmZrbSsWeLwYn
tXF3/GbgY5pIs8sc8tRgfTHD5w03eMXy/f55cVdvQiAWkuUc+k1aycKxtLLOYU6v
bihAZNGz3J7UL5tBL/6VcJQcLAMkqv1ssoaLkxtqZYyWXRqc99AX5dy1lYjgrriZ
r0NAU28EJZepTw5Poaa1RrtPsm5wtTtoxVSU3R6b0pJK5cTtrICiB5h478+xSkKN
n8z2oTLSVDxE6TZsBkMjQapPUykoRQYte+G51Dsvx7H+tU25c+PvzK6WHMA7TDWQ
OUrp/xGzpG+N/sT079rkJfcUnfI8lzJMSLFTFZiZ+f9sdv2DS5k2c4D2xb+OqW7P
BENDR+xsUA+/dIRlwKRWuAQTY3UjUS/CSRvxTR4hgw3lh0bTdJqyyRQeg5jSf5Vo
9T0tkWJBVzLWTwVVX0FdGLoZ2T4Bz13YN4BZdChvnMH3W/CqIwztykbMoaQV0Bxe
JDf3E2AvYIgwr/Q1IeMsQ0GHbpHA/RhREtiybZLFg2mn+OUkK70xi+GshtS1E6Qs
UENhgmiSaXA2pvLNXS1iuHBNk/IEJulIBP82+RV2oAwELHvi2JNAhywWhR0HMMYN
HU3UpUN7ZxtuQV8l+Ou5s6OIwz2RCg64/s43A63zAcSn317g9hQnh+JbFk3uYaY7
ZKR8U5BqFG7gUO7Sq6k9zwb7eldqMUQ3My9y2JJmsMQKZRxm9VG/cFfukK+AftIq
UouBCXa4BD7MhCBwcq8Q7WXomQ70sY8hRP1Tk5hUCxOPqOUHcJoZl5oI/V6Vv+38
DRimmfrjCX+6McowTL8/ofX+p5LsSdy/wiHo2u9A+cmzm1Y6lomfZsO6DglKnEmo
0K4AeXo7j7WT32YAHzWKCBFs2gcwaFaPEwH1q9p4sqR4J/ONcbh6C3cuxT5tfzfj
YOG/0xyAN6arjnHHdwKNqCEGNbf65YVmmpGpesq9XkcDzC0Yc6WRl6wInxwT4ioe
QTVPpskiclwRtuybf0mOoaCX+MyPhXfIYIBF2CHyD9cvX9ClcuCOEmf1S3+Zv+iy
BNe+b0di4kvm11GUxf8KdOWGMVPojisUR/m4fM34qE51zIK8H6LWVlHs7pHHxF/9
PJiJ7rC4PZJn1BWdW/jpr4bZl+2+BMkjqFrY/fH8XzscHUnPDPYDWdiIxl49b0Rz
2ezrgwPbYebdh36c+4toLiMe11EmVPsY5zZ1/grmK/tmCcm/2Qki3LmM4sQuSysV
70Xfodya43+5qxuB+Z5agiUVuD7Q3qJFxndtX9Br5aZ9YR2HPNpT98ikg0ihxNFm
5ehAVzxuD1oR8/xoi57spsYgJdt6uvpZlprB6tLV3LvxCk8Td9QbQLItgUrpHStO
3fzSdxLux6L5Ct2P2fOOLe09mL7L0On+1B5rA2lLVsom7aM1qa/+OkgIv4jh/iUK
NkmSmQ1iRAdg7oKuS1ksuuGs4CtvoeSlggLPHIFIRhqK1YAqYA9ohKcqQ5GyFMzg
owa1Ueo4m17GuI3MsC1jgO1L7T3OCmgytxB5A39RWd/yDl7jUZhujo1AShKf0BSs
7ltFE/r1yhRYLJVC+0Z1ILa1AwPM2v0oz5F9zmLVvlIB/0XeMs48x7TCpefNpcq9
oqkgab4ZwkgOIub3ap4kSJ3rnb3khWfNGvPOdUREBv47/msggzuot98YMq3TsSW0
2MpZfF3UpYOKMf5JRczG/prsRrY8GUJ6aqLhCf4fBXqCbIIW4/cnf0XlWyOLU0JX
y/psaoFoPkjQQegt0YjgEOdZgccL0E+owlObh67LbK+VOPlhqLehcRVxVajwF90D
xtykmpF4OgFjxxuUBMZrp7sAOzemOSit6HBk58lKUeF1baxGsT1+FpMPHeiySvG1
oSdo0spZNtkS9yArcXO3A+AcJPfNml+LpfdBKAMLVmbQxlV3vv3dtsJf4IY9hiV3
gSqPHGSoPI4DlRnxuHAUlnfy4Ah2TILxdNXGfajkbhuyP6a6UXI7fxDGKxM/Gl4X
rgFuc+RojM3D0Z3PX7DrLHVnFyzsBhUYtvH+RZpVJU+0NGowj8blh6H6+J+nVQVr
ljf7RoUY3Qw46IzGB5MOz3lCjdhoGsPwu+QH6GEC7NdoMnSHRYA+Noka/JB4crUM
QPBuSIEF2qfrjCypsapluIcqP/Ndw0JW3+WyPCqpXngAnpdHMGqvYrvweLy3VK1J
z4V1tn6JTxrJEjSWdo9yIs9rCHSWXXbTjjHDtLEk7lSKPal3ihikKxeizidcmExc
9DjyH1z6ho3cwyh9oOPHJFIzX4ctBWvYrMTX8p6bpngRQbNgnf+VF39tHlmq+wkn
VCwYhvY/1O4HUZxuqLeCPkNQnnF8ksoz+QEM/Y212pQYqMfRUUsmqDPFRYfw/RMf
RptqOlqsNBoUm9BkWzfH6jdqYJ7cjhP1A9Kil1iu9F8m4ANr9iGDHoAwQwuv6VZx
H73mQUqC2o3ruQTMWuP1F5PMZ89me2zm4PR/8fZMtUHN1wxg9HKZnyZgHBD27EKW
kH7fzw8VG3gYLuRKhh6OHI6mhlojK9aYvc7oHteiWDbrnqm3NAzz6gBE8FTmumXp
x+tBPRgVHevg+IaeNT5Xp3r+biDcGSApvh5Gxlgc5s4Cxz7zJK4f2cAK6rZQUldK
C7ehDqvk3R4GHT5qDWtGF5YhIAHJrbfUj1yWG679FJGmufrjGyM+d6++/gsMoTuw
r19hT6XcCSkHPr3M2L2XRVubSYx0Cnow5FW6yHbwtytpsYCmLBISe8Hurs/CTeyT
LKgeZ46WZ3d6Yg4xmZA9z+BAjX1sSqkQ61DHWp7OnGW/GhO1eXF99Z7ZI5ZfDBMB
qF9YhlXLi2LigjCbP79dqlx4Y/vo7U25FZJIOeMJzzrwVzDrN61INbeXs4gymFMj
sGCLcsDsHEHxM/7p255jX9yk35Zaar3A+yLk/iur1+tv7/0+uvjHJvUqhfdhH3rc
62Slsu46aHG5srkcXEicvz/htsrYp8C8Icu5R5//M7KnORSM1Hp8JxhEj2TgNCcr
/ClFz830LzMOrNI8RQP0jEAl5zG6j/wsHbCa/PMglUJQqCjpOCYztXao2jb5pso4
DlRL24AJpvDWgqL9h8JYfpCAuDTg5pNESULWc/gUVHchOGRxtbmue9mE7UCQy1Rt
isYIHnlUR2xJnvVQzrFO44i01eH6IfiSR1isDjBj1LYChdwkeQYAZM2p1Q5xjoxN
hBBJw+leLxR2qRi7fwBU701k7cekUM2GqoQPcQFXklYwy9oPEPG+pPsTcg+Lwpxq
bbSO3qjWALVHuPAsJPSdJzjb9rXPo/Fb9JjTxkze4islCXJxzmDxtZgGZHIwWfjf
iP8gTKLu3jZ+8f62dc8vkqAgB8OB24cqFigCG0MwOvTH2yoB+UNoumggEkTY9Oow
3BlUzHtNUCEOM2qC2OsXQGsiSCJm3VGWgETGA1nYyw+Gqwk0/yp3lGZuYnIHWeJF
SlBafopSxpsJ9hJjAy3KMbuPeVUxj4u705Vr5eP+kfshzyQ2aoO51wsHvoEiTxhJ
8Z5N6+ChcUgoEYe7xvOUUiD0PlKh1lgcLdP2oAudyhfPRjj4Ad0S5QsIXHH0AZxG
uCyX0gYTXPNuzYkYlT/XG0K1Xht+tt9rm0QDwmNIo3L/SxRSopJRx9BxJ7BVLvuL
p/gCHqdgxLoyMKU84pIoBc+UX2+y6Dd5c/TszluQRXhmzeVLBq0qqLR2GhbJv8Dc
IexdkrPZ+T3K46+MzXkhFZZMPzzqzRYAHq2OA2a2FisVZBnXwND3l6cTYO6KPFtu
0uqOIA5E5SWRIcyIbReAGOtjEBFOVZkjjwgJlD1T+W/k5IzvxeSKNSXiGh15b9cv
0ZibxkxiJN7Q5YTVgAGp/MCqKqrpRN13S2RB4fMiXlAqbb2EbniWkSBpw7F3sYOj
GTCaou+TuaVrd+ODyGCKGmLf3fxPHXQaYo6vpSYxxtkp9mYCz3K/g5aFD2evEIPa
POHYzyxazDReuPv0dJwjmBEvCQkcTvwobaeo4k8up0ktWPJRBJ9+Lo5ioe/aB2b1
Ihq/6SyI3fOLDCrcnDgvPsgOXoybQ1NDzxo+Gus2dlzMaFx5rw7Ynx5imJ+D1DT9
hmmQkMCmPSwdnhoQp1u1eMqPaP8L/dQuA51yO8MIef29+VYFRkvfCBtcLkq71dZl
uRHKvxs7STFAy3NJTklOSuLM1IF02TpcCEm5MIbK2H4ZlQVJwJ89RiQWvrpa3TpF
iIp2gqnxM91m2WE5ELKleCqCarxtc7AvxF7kesHlafUCB4HH5B1nErsOJzFWrjdo
y/IFk5hBj9yqNQLq96Mm4jTAgNhhW83zcxstEQ2OTKMjwA7B35qfplss3c2BDMbp
wYrB4eo8rqiaj1ijWinnzo8Yco+2HVQRTj6Y0LW+hVGXxRpVeyoE84efeW9Ts+rK
KJZvgTYiwmjqCXDWNFrGu6wCjOc9rqdP15ygEs7ony1z6uCLl4PWP06WTh2Cix1u
OAunaIMRfzviVwlcTBox7aBCNw2M5RxvAU6L1fnINOX67LNUUXqhsg8Mp/HC4RFP
84/w6i4DrvJI/EOYJAAkdWur4+5hetwEr06Svs6WSaHdbvK4WBGXEC9skWTtQ07d
sqzOS1CkE2qDMFQuq079/3d4uqkeRSX/CNvYefV4eryPMLaxPXTZ6horiUL6RfBK
RCimP0D2TyqN1x5y38FbSBE1vh7DlBaMWVa0e6JTjevGuNmFRklkWKm0gSEfndJg
DPW1zybDoMfN1JgXDeBSUz9LETp4BtUb3Pad/ydNiiIu3MtaBVVN1gYN5QK2ZRO/
1US6VtMt3+cD6578G6rI1gIJRB0bSORFFR0ulJ18ZJ51ymT3YkpTgJ5SVpAq+Z6B
2KCkxoj77NJsTZ3Ro+O1swLiBYSFt4k4ih8IGgoK72bPmPLd7FdOVreYZB1of+9u
QQDi1P/vREslcseJVBIvB1rXdiZh51LnlhGxCRbqNCm1bjp+xtsU8M8OoiD7Y1gt
YhiUEdKJwfiDqDg5A/ek4KJ2rYqrrLgTbS0C+aKS5iki1XLvHQzoNHhGMbdw9pB0
yYiYqXmxLKNV/UCDWJaHG3rMOlCxxaZIIAeqnTSV+3xqXE6DDkA/KG9rqAqUtt3g
5JxGPIPbNSyDvR63hE6OEMvWjTLzak9htoGmv3cF6FFpsoXfOy5sU9n/ca8quAFy
ksay6Nxd+7yXeZMCiS5x/ef3vMrp24EuJuM6KSUUsgzd0da6WUiexfWhwj+jqd4M
cuWSJ/vpnfWjUZh6f6VDZYlAY0QjZ8cjFLYnaYK2JwjpIazYJt0y55+uGD8A1noa
RIfgu3U9sfzzEdo0qJt8JIpx0azP46Z56R8oEdyLqfjPaaqVE1Oopf5WVB/CutKo
WXSRKymFjD/qybLoKLTp1UNZPv96QE14I1B5lL8sQomFvBUddFh7tBzgVLwhPGoW
ci/UdjS2gYa3UPm2Pl74Wfme5M16UrYhY5JiVCl1SJo782Ri8lZYwMSSRyq4cLKC
bhJ1R26w0XKwvVKQMPz7y+/ctNBtpWvo3K4UP4qRAHMbemL3CNgeWGnZrIlDlR0B
5+GDYO/vv0hS2b02uQh54ALfOP6OV86MHGJQ0Epr06UMKHmYwZEX3kVG+2lazfTN
QFJE6MZ4tpfzw11P+ovejKgdfyxrahFm4yNurqLw2pslc4kIjtPqirGpddI/iH89
8Xy3etL58qrr/SeoEg1Hhq8YlrXVpoaRKOdqqsKSPV36Idnv0PFaBXDEN6qAuM7j
LXjk4y9v8YvnjGWQ3Srfnh0M1OCXEQMddX0uP0Uz1XNlglpdl1vpRcKna93pQyd0
9wHOJDwadH32VTUODQobfK+/piSn5QI4MpAVvnG1Y0oiW+hxCvm5ZHb5XlLGWe8K
Lfe4mE0q1fvHGgf4XS/JT+3pFEyZJ44x55G50SSGClieeJmqMiJBGLkxswX1pPVj
h9Mk03mlEwo/R0+VYNJ7ldJWlSFvxnOsg5h6aht/N1jcErfaI8Uas5YA0bpupW7p
IeUfZ/kyRmCXpD7sZ9NFw3kBUEzhdJg7XKHIsuB1J89CogAI6Ysqs65+tmSK0mY7
U+S/r+dfRKrOqZvhUDlzTIdp1ykciIAKAe/EuSGH4Ow8ow4vxwRSTdp0Kg5arrfw
1m+zB9Nb6zRI6qyRNBTBB2+O1S6GKEHhwG64mY8mz6whhw1dMb7jfCVpl+sviWi1
OdvvHOgNnh9MEM/hYfza+ec1FutVzUzLR8K4bpYWREr1hrixWLqDGQ3ttE2s95UN
BIL/1r6ORksmR9PLUdDU/m4C+jWBwRT4djLt5hh1fdWMj/w08lQmRh5LBZiwhmVf
t5kLPFAduMf9i+0Z11WrHiRJ1EZlA03+py68I2wTdsadUXA8LuQyOs21JPGx+8Ob
bKJQCU0WUkUyr9vhd2eeAwKLNCk3023n9U6FfO2Y/d5oRH6mFVLngeW3rZSNo0t8
toXQN0gIXIe97vd7MrM/DWQjRw8hbaq9uBefhWkmTX2powHdO8ZAzsYSVQo8eNP1
q45EwxQh5QFU28/RpFgpi4w1dSi6tr3Jmru2Sser1FeXM2WkaGTsG06klXcyuKVZ
zGshGl9qx2Yy0kXL39DkFZzEma+H7JNtYPMX/LCb5VwnG4r187xcQCc89iwP0CVQ
1xG/jLd7HrYRlprCkxEyoM14c+Gs2lx8afCc9rYkFR7vkwxM02ZptbK+IYjArP5a
zKHmjQmLiFsf/Y1H4FrG6S20AG/rV7huTk6kvVsgyAz8ktyR5Uq/0IS1MGdePcIt
u7jpr6Cy7kV8eP5DNrrYR4zqwOCsn29KnMxnMYO7zL9f8kIBf/+785fGx0AZtBRj
AwfsHnkqN9NrnM+5eHjz7gJ/buxQ7a0HaPkge/bgFSzIovT8jgiq40mRt0CQdrDL
4tt4roI1us1EjkImmOvGsCAl3cZtmME6ZR9v6Xja7LubTNrEN6QEcvZ98IbLHeNS
yfxsWEbH6RqOZQKzgEpiNJ9yu8yn1dnPLIz7gpX2/P+v59WPG7ZeTdb5btWQ/vG6
Gz3WuwAMIKl3HuRnQUvxyFrU88gngezTc+g0G3SY+0lzmgIFKomS8XUDvxfjwP13
KRtYZ1z3iXx0aH2itHxlRwDicUsKj/YfWhMGwJKQBDrmRvITl33dK53+BxV56n24
IKlMV4D8f3ojToNUpe4e0T3ZrSOJkP9zqfkdh+U3YtGLEBsNCvlEsCF34Kb13bmo
v3xiEyrciH7+6SOdgtvn6CAhUI3oaIMGlDx+x8qPmcB5r2G7YEmVE9RjSiPCMpO+
2dm+a/LgKr5HCkaEQyoKnEQDtH1qFd6GDhTZRKCxeRshUUO+Yt9iUJ9Xw4UFOmV2
08en7I9JWWBhKw2RqtrFGSiJSyPsBFZWehWBIok7YvZRG53i1cqU9YsZz04H9mrc
Na1n6k8bWnXnZVpvmxnIET2RtURrHqLZybPD2ey9JXwZJueqkwFXFj4Y6s5Z03s/
6FR8Uw+iP+XuEiKsUiZbk+dlhIs+9y9wxmN02OMjyMA4MZk9ft/vlzm0rHm0mgsD
lTNpCHgaxIJ/7Vq7s9Ka3Ju1SoCCq3fj1k7RKgJcvgXDDoHFWvSKs9+46GgHTsqK
A+nUloIkgmkVSsaOQETpPgDbfc9RcHfmjtsmMdMJNdsg9XXS39VOJn0Q8sRRewl/
PoiFDJIgZtxb5Dwk8nptE72Ies5l6aNp1SNzLMAAvmoZzKhI1HxBt8MnSwpQzN02
nPoKt8fFPdjJ7VD0YT5A0I2eqMuXf5Hi972BHZagjNrSmuKRjaCiYDKM+hTCwUpg
UUb+aR4nglczEqWX1j5dh5gU4MfkPl7HSIArQe/ya3iZgBDZH4KApEnY4/wYmPhv
K2AzuMIfqht1fFrGcNCfLgdJ1eQopvXRhAhN8ZIsGN6QsSqiom6KLqd0OuC7SuJw
iY8g7Dyf+xx8Bqe+n+VfYFgPpliq8GtKgI9U6EudvCO/iLy7jKaP4Tmbyd3I6Tqz
zc8rQ0PMlP05ejRBc9XrMow6BxgzZVUXLuOlVAmVxDI3vefQv0NFEHLU/SJuUksZ
1gZyTWdiDW47F8bO0/XiLXET+ICfotsDYKMyM+jD+DeF3yvPt5OCtHUM8nlm2XV/
At0OTaV+PBFHG7Z0ecVv8VQ+Cz9dBOW+RhVo5l7cQORatgevYsH4EQjMbD1THQNz
408XTG6spkwJE2Wy5ErA2Xd+jET4Taa963aLlPc2Sa64PtVUPOOzi921IZDs/DB7
kD3hjAGRGoM6ZjMvoO1bIC7RKpL7GH3Ch9aMs3Ew3naCApOlEXtZuph3fK2hcuSa
M8oKaOpBtHZ667UlfSYQHFK3CbDp5AsVKb7vcOQDQQ8ddEK6SitzRCJvxNDq36mZ
2luf11LhgC+oaqK6zLDrZ20D2HKljahSIGiUzsrK1PaKmzsfABRihO9dK8vCgBPA
6gq+HMe8dBiO//QT7msZ4nmBcvg/Bq5IgpNUhXQggcdNKvwfk7aAr+rJuP3Eyqd2
4EwItx1lSUXNcufx45etABiJQLMTOX+eOgedPwmJ9AuyIGleVsFCR3upDOhgicin
QKrsjkJ8DOYldydIhdhOSIyCWmbbWpe2NjPiuJleMZJSBzrC6C6YHL93pVn8MjQK
p9vP3QfjmUTWCug2tdO1J2qrfcm/xyDafYoiT+u2t+u97z3a9+tUNAxg2vb/UWRJ
E6he6PzpPV5I4lcuZZZ2TO6tZ60MeLFmAD2hGowWjZ9R5lAcsglMFrOCTpu9CuOv
xZ2nRsjSrtYfJhcd9BqbqjF6fRCxT9vRsXP7+WWJ+ogAyfk14wLY8Zyo/gYFivxv
GlE/AWZNWFaaQ9QTBWs1Up0FqzcRLxGZhT+Kx0VnkI5znP4nhAtDtnAH8DC5QZb5
Bh24gs0bNTflh3KoSsbHyMmUz9BCaMLP3vBxcR/TrskILzB4Qg270u9fcagj4Mhg
64zYXn4jD8fMuOgxC+6LwP4vG8BU8HgsKScVYhlE6+GTJ6Tsul5wrxMCCribyb/q
aCBJ5SCkBh3cAl/h/3GObeA9Jbf1fH8DoSWfxxzouqWiUFZgIZTPgK8Ujx6SS4OR
KyoDKsfuXZuRK+UsTDwfEnDwb93Ee8ukJhlvxPn0WaNn5alogho8lD9vTP/CdLCB
gvkdS8za73P8H0TRSAoK/TDNB9m1gaZLQolPhFesR5cKU3+bIMlt0yeY/vNxhby3
Wp3g3T2vlhKNjwpfS484elJiFxxFLZ5AhgmWqp/drBZooCsQMP2ZqvlWriDARV05
ee4JfN/F0tCfknlcw25Y02WjUk/9PJbAT8w1n8JFbRbSie32Xrau3Fi9KFGLEu9r
0oootn+M996dntAJdEQW5h5imTvOJzytjcLZ6LjxBITccBj+5yxAY8IUC6kKdth7
dKQu4ovIA/8ZtHjHu2dFmRL3EfO9gQpEM1Tp3U9HOaSDmLhI48BXAxhcIp5br3ty
8GZLJftdZ4jqS5QJcPBma7TP+cRmyg0YTlXeZ1hrM6AtLu7qtlu3ZgCs9UOZOclp
3QzudcwDJM6COigQAmN9oeC+DKa/7ZK0Y4bFElt64T6aH0cHpQQGaqH9zCJWI0T0
UR0CiipwBgbavzWmgETsKkD3oUkqX8JyHI3QX4ongyrw5/Y+9QvrZ0KRqQaE50q7
VXJ2Rf7tQe18PpymyTMPF1QfNZpC45qtekZ94F6cK+aElEQEv7EKKzereqEA10YV
Y6jGbHm7BROOJa+Y6qsUGA5XEA3/6qpL4Nh0R4GVscvC6TxU0kuDRD09Ly6xUt8P
76ltQT1JBhldX/hhkk68lvP+KddPr+JaUkCqvMlqf0AK0oqX04AsqxMgiVHkAtIh
TZCBQ1q5YMd9oXx/FWIKSfTW6aw/LDEjYO2cHCSo3vgn7EtQUcx3ewcDjFrFmjZw
9KGfn9ZRlfZ9/ol5c+2CUthdmN61QJPio4XhiDR40RK9+z+hYhUbiH8nSB+B22tl
LPxRdf9UoSOSkkU+RSz61xMXNSBCLiv6+U+64UoO2aKMnD9G6oo6NbGdiNKHWMx+
eVKpngwIXWttlmE5cTbtOtJAufWb/JZ0MCMrUpfJeArgoThHme8LQtgcek/JNK0G
nO8p+yMitdu/Ks03itaW4osDiJW3M5h17OlwUxrAmBUxSmzzzs21NnH+Sw/GX7Sj
vcDTo7bshK5sU8frhVxB/4Ulj9/7En84ECYBf8frs3C3KecWeOtWdFTCGGZZibAz
ytCe3/C4xHZ6kREuGPHQ/C6CDYPraqKZ8fpuBmY0Ne7ILtBdz8Qm9AXPMcJMI1t7
qitR0FV8zsmx0X6L9LRLj35TK2tUBJw+0ff1QXPFRXDlJQF4EBkkaA5op+ldRrAA
pvSPjYPHr7oc6NJxvbxgI61wJGIrWkWJ8sCVR1xy2MS/P4VCt2IYunNQFVxeIn+Q
jnz8XujNnNORvaRT2WhQF+o6YGXHGQEWPxeno2rLv2DK07rVIfXj79vwxuEDOPHH
9Tza/hgZhPM2qeAjkVOOj32oOsoLsy9YRpISEuEaKj2WKumUWLHVjjt7zk4oD7hV
rnhrNZuiGYQnelXkeVlqm0j2uq5KvVx012H0IWQH77+Px577kB+NcJbb/oyDoD14
0O1Rcl0ee7+6EfZxQGUHUkhprcjahZN+v7ir4SwwvjwWul578yYiIpE/hnitQkZQ
lZCS6GGqyrr3MjPCIBwqceYUo3ymVpDP6MjMlAu9XoLxjLohX1lz+9IeMhqXjv5c
NW6cI18S/PLeqgM0lrWdXYytj/8XVkW6pEF/vQetVcn4qIS+/J482cbjAFSBfKKA
o/cTuOS1uhBMUVLlB281qp8/2dvuU2Jm5zqrzvRJQSqcjtc2aMi3g817XZAbJnCJ
nGLGOTqsbg97jBIEjb3xEe9LcWRDbpFCbSHThIqVg9ITBjaCjT6bZZBdpzuPb+IC
LqzadNWrDDcMRN0f5JqB9/LY6SPO3TGPrtFri0qF7WLvAryZH3FFGEZ8vlfzqRyk
S4jxioRZkNCqvJIe5DJGEOQx65GwKpKl6IuaG17e+c3VwV7BUi3MkogAA85dkoAj
5AwshOoLALukqTfkNCiYPUTgWb1P32MmNYgy52rsW6n4/V4Sw9+/ae/ehZ8+lNpS
ETpYHpK2sqV8LJ+hroaO8xzH6uU7+LSPE9nCeUsoMkpdCVpEj+pJTqcSEw5w5dDV
eyk0wInpOZnnU57hW4zElr3gEowA7foePhQV1d9gerjAxTf2XtMc0gXIUojbJLr5
YWrru+Zryo8j3UtN3gx6KKy/+e5Hja7RQ83UxNSwtsK3xi8/9yg8B91HDLuh4tCU
Q1gp6Lwl9qq+tkbKL7oEHSlCjzmxl8sPZ1ZIk6timZssgHnvMr6yuYc2Kf4e58xC
pEmRjyHniyyoNp9p6L0kwSAc8WcxHLRqo0LaRaA8aNNi7vKVehwj8YuBv0L+jQMF
ugSvzh+ZQ+8VfZI4WJpFXvkyQzpSAr/4zZ75FdzAzgQcjcpxdB8RYXObl5siS/nZ
LCklTEyNwGbYlv/XFkB5hhNiKtiuJUlDloPKsLKaOQBYQntiClTaYo8s5titwr4s
zyFwqbVu0zmxbxH6bZSTR9kgu6orQUA5Fdo0WKRD81+gkMwsJv2OpPxBZeBhWsxR
aKd4yEzhffSoOM0C7NpuErgAqHaMmJvlYlx4ihW4jm0W9SuDOCFiL57pHTL3bH8O
p58hEmxo5eU6KeSNHdPT+wAohqLIIXJ6atwyeSiVdsk8fjU/5PMIiyKHXIEN5oKV
Sw/hlggSaVmGlMA0dZzurJt09/1IeS30EM2RIaoYoePxuLVH6mxPWDsk9kBmsdGI
OiYVkGg0NG+9Dd0z/ajUVGGHcjpCVOsAKRJHTzCS9W+XLtU56M9sNHzZrn0ueynm
Hrz25XGBAKhq2+Gd+kGYexNcHzHRgpNaMH8Ixp1rATFeon/EJL6Oj/g9llRCH/8R
VD07H0cfuIk4y8LPWromS7gFEZKmsaLZseyxEbK4+S6JGg7/fkFR70pfdTojYh4j
XcHNILgYzNKr1LFmmmJK+YXrZ50UY4ZAOTfUlH9xNoBL025R6Fx0R4J2AMts1VPM
wazcPvFaleEKhTrxa18Hp0NWYwZiG8sfPKZQI2zH0G1ZwgxTU9PEymzUWdl3naR/
7zM3AlqKA04xVcxEN0vQ40TQjp9NJHAmh1sadcsfbJlmUaqymuxGVgxCe1neBwDa
DmYZIM16JA85VRFCSkrMmakU6TmwFP+YwfairW/ppnIMBPxzenRrnxtBfo9Wce3x
wcPTPZ+gvJrXZhTF+vkdjRqgnIZ2PaM4enbkrl10bPJ2y1LOLby+0Okrr3UPDRe/
O52LVP8AaPXvZf7EBFc/Hj2HL0D9OMlLy0JHc97qgL5/WW4u6VkJCEW6CkGYSQUl
7BTzScvR0W6OmCEKNe1ByMrTo9wHf5CvJpnbeWCpeKMBHfwbmbHb7gv4gP3q5VGU
8HqezmoteycZLFJfxbGWGcZtBOtcTUuy3GmhWZkMKuWS9Qyyk+nJvSPoc4shnPWL
Eo20VAl6t3gaVYEOTh/Qt1UStTvkRsnZN1yWpO4h8uYTlyeC1N53LOhcwLIHijPc
aPh7Uk1r6cGbckWVi828vCpdBimjVo95189BxeTGOvXJxfe4WFs7dNhku4f6jl9c
FRZ33naG3NN/cOflreFV8jlh5PmQKI1VEQ+OeUNStywfrCDUEa8KkEfRAO044UsQ
8ly54GhiF2tLf5aJpn+1D8K8zLpFMgJenrwp8naHydO2woFc0UAATdeNTQ33QLUq
N7E68foefxNx20qk9EpM5bk8k2pxynmB3gkj7qIF9RF9SAJkk3NYTn6vGKBVACzM
ZPi+lMcp+NN8fRQAZOaC7S2V3hbNTG+6RZKH8h19xNsdpR8uY5Y4owM39zdMp1Hy
MQQ+2wAfx2VEWxecfL/D6EkFA6Y/dR5Z6eZ6pvKLV90lOxUcfNEem3+Y02x5yX9k
Yj2i+yKh12YcE+f/1er6OvklKSZpE/xhNJ51kFJndBCRsxqdrKT/hTCnvNs/KhCa
dF9WjzUeLhdBrF0GUr93NFEzFJAFyFCIhWlvX5WJoc1kEOwRlfilZEGAME8rHouO
9+tk0CfaUS/UVhV4BdNXFlKoe2Xe7e2+ZR2L1YcbWcoZ8WsN3m84StUAfgbAhE6N
lqJahPpDFzY6yx6rL7RmXtZud8IkzXtIcBK5+6VAFBkNQlGO/tFo48v0Qy9VkvB1
Fw4LQWg0oGvsVqaeLd68f7ZS99HV1RRjsPcPydbIkDjadzWv2Hnb8BycRVShmlE1
GbAERg3fr7FH0ZD1eoOKGDURk7Yat99GGuoV+7//wAsxQxkc2JPbNo6adzNvqFBG
ZTmNuWR5fASIM2kOGN4Kagn8+/vML5R2pbVAePnplaLlmxrHXYo8htX5ZcqBE1tN
jelNngIpI5F/4Jasa9uCV+PP4rXbYgM7AvNhtMY/bCA9ObE7KzViX8Vb/fWKfLJ4
WAPaLToLfSmqp9EwETqBqFPdOxGj1EiS55/YvzR/2p1oqm5TDo/7f3OQIKiHzaMC
+SeUpVCFw1/fUpwQT/tNgQODVgeGQv05htia6jHWO+GKPCV9K8SRyVm/s9DudF+u
k/IsLNRFgAd/2jJcHZPKeIqZHvgARdhTyHVQwzw19BnDz03OhJLuL3ta0ur8JpAf
+G7h8+Yi/5JhRoTrmhpijWBVZzivgk4XK3G62EkAHRiyPo7JU/QAWWnzm8gD+9jR
MeuA9mkSIAFUOZqBzCH1OIqyTAaEOkNRuW1GFs/b7KUNMVyrnt0nKvS2gg+MnAfN
xnKWXzXwUqLelvHx4X70yJJ7UqJHrN/+Ogj0iQLN00geF3fgFC+pCqdtrfi5La1m
x4fF5Kmmc+Vhl0/v8Lj+HyTg6EPhK0cbpYRLkGm2kHUQEj9gPcCwxO3P8K9n+J9F
GRYUM/2AhyCI43sLFnkc2YB/s0vP4UdDP+aHKCnijaHH6ZOm0XfhQJYSMsow81d7
L4xa7uo/ysEvXjIHVb6E7jFya+PZMmwWsrFCY2oX7anwm55c1noI5mH4tdItxTfh
HTrYl2EDXSLLo1FO/+OODstMquY2ZhEXPHZ50yVnSp02mnF0zC5CJoK2o634ticG
bxJhpuU5LpFRtOP1T09TEnpne6PFwnIWzVnJy0vJYDdJcHoL3PF0dMv1o4LA0PSq
ieEwLuNGGNnILBJZnxoIxclQmOfyQ4NBU7+bM3s8eQq6KykuYYl9a2orpHT5evtf
qzfPmxeYkxY6wBQzUSdxwS3Ls1Z4A6jV3Qz7VFCv1d9uBS5a/5moTHltBFyA2fN6
+asUbQp9PvzZGilsVSD+GCFy/njxkJX40S8lMQa4I2FNTAb6YT2aO1wWi5f6sZt5
U6YtqYE+3nxyst7s5gDn1tppvGpu//TxlmCn8AwvXwwBw5jOYdaNqJwHQU4K0SWR
7VJpyPfFy1TVVym+cocbZgu00oQkRMnH7MMQLCFDrVNjw21IOAQL3xz/UL50FlPv
lxBF+Xl76WrMI/QUigge6q+Xkvtg2zDcmEixe8RTheaM5hqNhh9OakiQsr+0VcOc
Zqn+stjq8fKEwLXvmHS8j/nH7xOuQeUuASBq3zEB2iQie4VdEyDXIrc9keHgZX3G
69LoY514XmqO3djGF0Bg5r10UsH2qehP62cn7q1fKmPW2VwiP+TA053dRXKsYBWw
rdEUtQopTR4CmvJToybYl1k+k6ki++m0jXspwqkr0fTCjYit4hAQt8ndU+hfynUr
krzmMPWoz/hBMoyG/JvGEayvWBSHFt+f9vfthmqAchnQyCKmfDW06425rzRGbpOd
3lK5+/w2vhHel+7/pC+drbKswd/zHyW7TwvWN1H2rHB7hPY8hMc99rASjhdJ1ehy
g2ictqIMJtW5hywYLhl4jPHt/ZHkUbNhzSWGdb/dOPy/YUXsfv6HqsSM82fCPPC3
u43eo0BiVV5ZfpfHjgkEr+l+2AgukJthHIl4C/qGEe8OpSOzp0INEjlDrHzfDb3V
tVAy6ev8BLLOqvRQR3CR9ubfSNeoBfEMhy8KxMzHXaIut8v/x45V0WX9Qj8eX1jX
YYj+oHirJ+NGKby5eeHDW4vR64z01t0uOGScU0C1W1rv1XNnrTFIqVRkmYL1ihr5
6GKcjtv2bR4MmKP4vK88hiVaqZSmKYZxuxg8tiaNAxsfJZ70uZF6mzM/jFtyHHwR
qm9taRGZ275IseoZxw0eDUiThRNmgzXr4vMfXm0xL14pJ6kCtoXP1pxIN+p4QiUm
HQMiEz9efqtFvoRkQhx0qaFj3ihl9cSGw5pjiVtARmq+jbzwEhqaTnG+3acftaKx
YnWar6NY76G85LRyOckf3MFvPca8GSNqj0NX3SIfMdojgD97RjVU+1vKVWHXXgF9
xmlqihZJXXIoffBg84tjHMe3hZmmSBQnhmaeCx9NmiQXAK4IEDoZ84elwvE+dAmc
rMUjntu0Xzb9SMLdWT8A9Xu0NcCGALSgudU5tj1gJEqz/eVU+xYmGiBzsBNLiCks
uuE2t8V21jFW3FACPi1OLP/5s1Tm8e2VKpBD7bsOTMXGEOmUHV89ozUsb/nqCx+u
s0WI6tum6y32vx/iUQ+DTyQoOOpxlfbhhe+VYir480DIBUEXxZSow3uX60Tr6+FO
7LhEmxSVoeRBgx4RvoMJg7d+lj2DwN9pLhyd6qnOO2+VcthuC8FN3eC6PCere6ML
w01fFX8kWDulWDvT1TwaqaT385mhGbFcIoelXhf6gtg0TqDqexoWqQxIEpg5EpnZ
HppfXwR2ln9Y96xESFp0Qpx3NJcmyZzIeI2/iRCOE2MOmIzsGMYZPSDNJhX0/BB+
RJnij8H1jdyQ34JTgOP8ibMIAECpcKWsQkbYY/0qm5dEBeRuH8jylcfDcWcdg2oS
iEnmV3+GM3knWmRVV1tmXvNDQua7ymrinI3zaRxDMPaoFdUoVuRGgxBbzfK7Apom
mrYMfdSA5y/ho//NlUa24u9utQA45bZHrBEM5o1WtPWy93UA5AsdUbEI7KGIdRvI
UTnDVoIoAR8XzhMOV+hzN9rIbYhT7T+6u8D+AriPLEBZxJlQdauyy7bZ+jTXJvis
2fpE5vMHOruN9hpdazPT+UcX1qZRRZo8MjFVaRGgFcRWW4ee0IOydYJK3tFa49mb
G0RR6COwlLJ+4nD2jMOhG3W59Xml9CwFYlvZJVDd31S4kDu6pbI3/t/UbdVTme2f
ukzJ+jzWoYohKoV0L2jzOzTyIkPe9T9JMsOB5crPXv9eNMDSy+V7R2XPUSkKBkYi
zRJ0AyZQ2YPi+nnl+s3Nywsw9TXk/U/E0Rh/HHs6gwDy2TnaYuf8u1d65mDRfgle
+oFSPw+RVzmnpBdSrPJ0ghDKvvC0bvG1fhNKL/EIwUiDyP2zx0r35BiuuG9UkJjb
xr5+AMI5PdvlCENngX3+z7Y94NvvWKIB+Btsn9uRFXJHe3a+b1iyGMPsyIjm8O6v
5agGaQrNIsVme1OMv9sLJzO1jOCZik+nzOu6UyDEOHrBCDjV16Y9W4Y6jrH3OC+u
3HAIcyfmbVfnW9U1MTCsnO3dJ+bmQ7D982Bqi6Lgmp6ISw2sFJQ2mUYAuCIgUuBp
Zaiwp0Z+sb8CD7+iIdhnGrD32StOKQWq3njrRxYyghNr3dppgdz6fp7S6kcWri3P
ElEFqpvHIbm/Ekbwxd2na+lAb771/rl6gWELqNnvJz5r9nFHaNohS4Oxe/FoC2D8
KT2Qc4UXB97JJjn0xRpJhXcD0yHYCR2dc4zF5hQUVV4JKpJYc3XX0O9lWG8eM2/L
6ggTH1BNufMOXW/s10sInZptqzUnHTPFrQphkiHoGZRKwg7BRhingw5YQsLkgaRD
SL7kHdTiugahffxuFepFtaObF1sKldJtHurmANqdZpVjkPgkYE9lxHE6bWyHZGsx
dYxxp//TVH+nuWAgFZ2PMypJ1R8Ffustoyj0m/LL6ZravMRBdH6x9gUrq4/2fooJ
76UAkjT4JP6a61znEsyDYkR6XEY7LV6lub3Dp1GsphPWaUyahOdQUKu86oKiMi2D
JmMlIj+U4tqSb1p8/2wwfR24jry3yPuzd8UBmP01iViGQ8flC2zm+IAdelrLN9RZ
Hf+cX1psdbzarkggBBrrgyP6/ZQqVcJ+O43I3Tx9ebZ226YSfSNRZ07UfX82J+uP
4v78TT3+zm9xEznF5jtIdHq8eFY25rCi4FDnb1+8WRK//RxGp1Z0VVNHNWiY9FBp
HditB5Ua8nmPqEkrzmGeb+Fiw94bUSsRbZifuuvFyctnIfZrYvsX1ta2bowml7on
0evErNFb5YJBF13wjjEvJMfg/aKFK/FFDlbgVRccIDSLZD/f8r2fCwqcLFt+Cpp4
4ijs0N5j8hscZ4hstGpVVspQlUp81Rmy7esVmocqcFBO1TbBBs3weuZ87yvffl89
C+WYICqeLZVHbsykixCFz42wLpv1MhHe1iwXtBoU7/fQ+eGo4v/j1G53J15izSv6
2iu1N0oVxTF/QdBHEXusOYvw90WCG0Any3xDLepaSPdndfmgSOBYx+SmS/CywC0j
z7/nguPYlQLv+IGxM1kgcimfoIhtRZ8A7gUprGLAHIHzJlog9yX28cQC/isUtXGc
MjJkawi3e/Yn/4VTxiw/iQGjZWvxG7Sol9dappjCvsJuA80ArWHn2w6tXvkXQrwv
Wukt9GiTayJbeRRcxzS7H4hdL/rOQ88Gg4PVey1xzpqVbWyQbeXIkgEg1fvDcLq3
IXh0SubHgrDNM1DD4JWwsea9g/uW5FLoELDd9OY9xjljGMdv2Y+4URVdVjAna+lk
IYccoP3TKZeW/amkQ6JMPSCy+dd+0XZiuowiopIufBfxktlT2RLlok3ab1qiIJc2
3CtAjPyBPyiMmfg/x2UrnkNm35U1UIA5YMrgDEACmkJ5wsxj9XDi2W8Y0Wb4FFRA
eXVot4Z0TxNe1TIbBPBxoEYidc5dDdCpmFvNFEob2FRUCjbQMaXHVqDHTSg+t9EA
z2GPmpDeLZm10aBTlddS7ntkwJvpEw/FBvqxJd/nQ68dwkQALWrnIbnTIeF8kMg+
LH+CrYkFUOzF5JElLC0ADLCOysOipvCPtZo9tz4LS51IUX2G2ZXup9TprbGaK27S
LfRsfU2D5nyhH/1cTnv/Sbibaf/k8aH+6tbINiLpbOCqFIXWZPYl7QLOr13rHKpV
Du38plwmslBr1ZCwYsBX/U/nGgJIObW15UgQYGsauqTQ0pBKeVGaOBzen7MmG0zL
o9dV6LxXr7Kzsw+jyseCXB0WPll4Poi1aoOoCGfiuNiBFAhWpKugM+j8WbPdCi/u
kgQDFRh5riYd6o6YXDyUUl7XR9TAVVaQMvCpw5mUqD+63FS6hcz6jGY8c+/5X1xW
+JgEf2qXn/EgUns32o4ia6A4Vo6ghN1+0fZ5q3r5J1XUczN5F8AIU7yis4hmsPPJ
74P7bV34kcSj3rzwq9yA80vfKdI3rGQ/i453xfneZWX6KBEGgRSZsnwBVcASoIt2
eBSPclutIKde8LrrbBuzGebZsf/zZ+yqj8QVTZgwtZhOqUr2bBqb06AgSqAAlI+S
Sj1snOzlMSjk6m/Hiw/PkSHEaYdDElB9Fv+iQbstvf4a8PGk0CavrdeBUea5UFOT
ar4Ttt7kOoCYzHr1qjZcUdWmTA7GOtfQmvC+kyPmhEWrc9DcQYkk1KhpKm2u96id
cZJxHWyM7FCWcYEPMBtafrOfM5AlxAqCBMuHR8zwI4ivje4hIC1fWV7w2pKKqCgG
5pKgQPhnXo0CRitleCUxsLakoxuD+E6f8Ek7LemRbPPFVpRCt1Vp8SlEkRME9/rg
dEgvb45Z8Q3IE1XTQUcDHi7qGLDKz2C5+1l3bra7OT6LUocVYwYNsugXjKpLDB8O
+VZM+NgBsRXs12aO3YDkdcZPFV8mwPfOSXNMakBltTasP71sd8gpSCocc8CfzpZC
W1GynvSjkvTG5vwMpZ5xUT2fnfrUtuUqp1klbWin4arRPcGJHa7UXjx8cE/U73eq
VUrKFlzmCiViBGLZEDDFTN7deSGzvSlEP2XVoKGXAhrEM8l/3DmWVisOTEJwUltI
dvuNwX7jFScQ38/g1IyDYd2tDCP5JlyGsN/Y1Lu7IgQ6sPwrOuunnfYaEB+Ro6Gm
01gdKuJJx9Fc8luh7+zdtRTMZLTK6TqtXVcJb8id0VHrnSlSgqUcbIltoy8Yg2tO
IDobcjEf6X7AvHr39jMKopH2HTgeeVfICpABc7duP6BwNds97pkHjGQH4qdJqfOx
4oVtjq6zuEP+ma+Ye3WhGyES1TSkPeGEfQpE0VdxDufS4ohVnEW2f35OLpBTYa+7
wLSv8YsU/FLUjle+csNSlttFmKKYGk0Xahbbnk4//fMCeGTKdy4hm62ke0PL8G/3
wrdi0cXVASpmG2FxK3KSHgB1H5VohETQGp+9lg7ZRYEOJgO8/+4ZVlRYtDdPgy72
qehp6Z/Hzr4Chre31eoIq83ob980N7aYv4QD27sSIGr7x2GetdCFC2Jr0mXYyZWd
tgIWNLOtlngee4t6+eMhff3AE5pZqCeITUSBZ/86coSfT4yzYdqgb8gU1++XiUtv
C6qOMiSWj0XgRuIPXt/RIkswZLwXhydIKFfgkzEkQ0mVwOHN/fzA7+2XOK9+H2KR
+Lt/BqSVM/ZC1GzxpI9OC/gZJhz7VIaGNmGlQ0o2/pzP02qntm42RUyGrUZP11p8
T6CWJEIOog+lB1/lrZlEXnxb2+NjNR4cwv9vEXhqkvqufEuZtgksQCE+bnPvVI9Y
flMLC9LrcKZMf68pJXKWgEinfFckhC/P1eFyqKA0rrM9TMY1AY/6LXO/Ag6PzYr6
Z6U4ygHFxpAHPVNUmdSOapkD+216dvoX2Sp0n4DB2YsMVXsd0AeYPBI4zmD2plIo
S9Yx4s7KV7DkVSqsS+pU9o/K1pZ9psKUToQdGNr23sNzyeWt2Pm5f9G7ZVzjoP9S
9TQJDIZUWqNHpJXp09aMpLFLtn96XF8xzvJ8LG4hq3F5T4lUE17p8jEsrHGcAMli
q0WXA0jtq+I78b3RBtX2Ge7Sd5qqxBnrMJaAVOiJ8F81dc6sgVPkefbgZjClcNPN
JZ7S23jpdPPHozX7x6cpPoPL1qSZwndNd/XyC4fbFa/Wx4SCXlnoKWSMuo20FPIe
GRya95Uet8PVOMqF543AENpOXqckeH/0lknE6qEiKY6rygMlmUtqLcZuUKnect6g
DHR2eoBlxBKNKkSZjDgc8vMY0gQCrK/dci5cLub4idj5ShfPFK2LEXd6og06U77T
8AFQv2TiMIyhVmjUK9uQAbU6iX0Twxn1dAGIgytoi/QGVDJccJIs9TyRyuFi37gt
c2GxSiKahsRitRgv9mi/Oo78eK9plxjaVwQ+8Vk6hryWPFqcx3CSgxZJyXH+SoH6
ya62qAzIBrRRc3oNc61IHUzNjvEph8qDZDflk6KdS3bj/1zq7Nhq25cSLXpaHyzu
1jnX1H1f/Gm9Dfckzgm2oAazIQ2nBllLK8K23+pw2jy73D5r3NzNALtamJFUOLj3
z0VKHTGgGvT0ImWLB6/Ggwu87d0Y73yIojznoewLdUiMctdnSr/8cVBPp+O36Xod
6qTuioeb3QB2TCiuIC23BfnRNBOcPuDEs7Y1JHjF4ssUfu/ZmMDejcl22MhRXZbA
XWABL/FI1Cxqu6ltYe59BVoff1NGNBJISNgl16nIz1TsmqYFwbrlIAG7dtXWe1oN
PP+XQZ7THC7McCAaPrNWpikjnGwVMQ1xttPw4Dtv11Royf17xKCzxHZR2evrYFhd
3aEysxtOiNCOPLSxxYI/fkT9WIedADf6Rx9u7os1X04PYvInQxO9/z02plkZqARR
z7HFPf8tpUvbfilhrerStlYbecz+bEGF4V3QfCpB1JGofJR/+gzWWwrpJyJxTDWa
9d4WmHYv2Nu5LVJnDGN/ggz7DatEg1q5TWQ+bjsIEc3YU1c9rrJaQv0z1tkHIh/g
cCO0hL2nGMJxY2FY3iTmX9zIet+2e3bH3Fu7MTsnd5RnLa/y5urYc9x4okNqony7
LtYefLWMwRZNFfI+HxFa7YNZdAD1D9+Ch31ir5x7A2k4l+b6KUowslnzpoi9HO9U
7sl7oSk+WRbQmiwzw2krOjvWJxtRK+6cXe3rUfmCkRyzFPfJlBPufcLU9CPrlOoy
f1YgCVLaCRKiVvsD5ylGzuPVYzHtUvA5d3jinVxCWX/Bv1fvFxgaEkmokCctpn+y
nwRuEso252yl+gFKCrPrA3tiGihOkknrImtiJecnEr85tBEHY29wd1XU1pft1xqz
K0RRFpEzP6ymrJYwHPnkpSVco6TH6BOHqLVWYseVn9x5orODktNznT0DeX9JNhJu
Zy5cNwVkSLO6A2b1KSBZKdvz0GzQm96jpVjYSQN2v78jCpZm6W8pYsw/IqkB6m8m
FfSX8INWtWMl/r1BOwt6SjZDVjzbeaztXdFEkF6V8On1GMIe3DR/eLi3oWrHbLqA
Mr1UxoRLh/Gg+TEINQHrab9UiJuuKC37YU5mIpvppf0OgbSuTS0OhSGKNFrW6Em3
+gOvjjNXOBt/CxhofFO0e0pl/DcHrnDtumO8aKXlmnynMOiA9MkSG3hqPMLf1gDw
tYkl+KaZ1ye1gzz7DkbAy0Of3pQq0GPLtYxMNk9M0RXjkWizszlL1yPyh6MbAujx
T+XZ6Lg+n+DNXVIyBUbE4y+09/FVJ5eh3cQoihCGxwVvK9PTPny7z4zQheRQ3PWq
/k5NeB6ho7f8m6s+Q0NbxcHj+lbuVnGJlEqt4zqIOWgk5nJ/7K2uZ78wYt0QyclZ
VfeKNlAC+8kI75s4Q2/gcnHA8C0x7OhlmMb8Vu6Xvif/LOaoCHpFW4KMjPQrS8SR
5eI7aZ0G8nAvhj1uqjqLnudOkvzN1K6oB/lELXVgcSYflb3WTlajxy3n3SC0vxr9
Lfyc5RL4Edx8xUYL+cS1JAXnyBRRM051nxHohAUEDZOwht7MyRWF5COe2vilZcWo
QFq1GpuXYbbvVuaGJM+pvnCIjKMAWLb/cz/5+atPwNYDHQoRrjGr/Yq9Tic7zvjz
D1obHdLfJ+LdtwHNohQQf2YFK+KgVWWTB9Oe802kovY9T9QpqEYNFCdg69vJT/8E
dZnIrfHqPs2MTvHsweYY7j8cV4wVEYai4CF/Pm0l6awoxvSlS3gZmJF2DqJiTsvp
PrXaedFEXCud0HMenyqr2t01Ow/Syo9e3kMijwuXZw2DyIhrxm/gMRSp8xj/0Gq9
bib+zjE9aU9SG9yATNKRgQoXCD2nShm/dcq3Do5I7AfGNXbsM+NO5zrSReN3qUBt
kB8v+5tP/jW6jZqID3IC9Kcl+qRqzDUGYWjVRcPO9ZJFWT/eKcD/aZjlpo/77h8D
iBsvM6odX9/R+lv6oWfbNnRGvLxU3zi65zq1XYa0QGQAOwLv2ujYq18bzTJdnw8T
L+DgL7Q7U2KSEfGCVIvnFmz7ARhcqC8wVq/nqFgF1dkW1l6aL7iDi17k5mvinX2A
7Rj0fH6X0f/1cUASeV9LEG8Pt39Xbz31LdzTjuE/fG3bT+XVQ0j5kswFMj3jjZqA
AJQ9dzlloMYCgMSY30WKKHl5w/gf8bbiJIGauiwz8UeeUV/Wq6k1nnz97s6jRTo/
H30UCPDcs9g10dlWNpYbC5+Ix9Y1U8Pl0wXLaE+oRCx83fwE75Ciro0JKJ8+vZbZ
M79jVJJlmYgk+k+J+WUgFDhEinodZT+FTK9rHOyfAICbLZmzkRoFsyL5/kNjurY7
VP4NMWbgw2SuQ2lljaqgYyzA6GkLNClpURlQ184bdelhZvc0PShhHfc4UW1qtHre
vfPQtZ9tv5MX73/ymIomYlbQ6WcrD8yeQbRGV7tIQPsykU2aY8rgbsAIg1meURVp
5RFWP+ZSb7D1j7bGV10WCNY55mnWGz45H7gSXz0jverS9ZdDc+hsueQDnLxlGulL
lWvXgF2VAkuJBVUn0RQuundBNJue29DFnf/ifDakXWKABDwOOMaQM6QrIBWi2JwI
Q2zyDWx2JjR1UAKyQguKbIMYHC3xTjgSGWGbHqgV4oi9Idg8Xuad2U2q91kYJlr+
S+vULUWlZ9GAAILtULhzgXraBj5haJXdyqrJXTdYinq5ehD3JBr6BAwLLlUN+wLR
upzUhwj/JvaBgMNEDIpOP74+OIJrn7/8VbwRiLDoovtENjSIlTAzVCyx/zYjbn+y
I/RaaXnyrbvyys5vBzXrB+cdV43CTWrYVzDbrXyK3ENM+H1TsuBAUG/Gl+VGYYo8
qQzk77H1Fhaj/x2PXc8cMN7faY1e21LkzIGANDdl81OE79y7aQeXgi4elhFmkqBk
Y0lqTHQc37esbZ6tmc9VVTl+KEyudq7gDJRaHR07xSdc337Rl+qBvhRFZh20fiJt
t16LDCx7U6KevqevsxvaZh55vs5BM0PrxglfFcxy8cRJsNhsiF2PAqpYf+KWHeO7
kdXMzSaL8FAnPYz3GxsaOFNuEtbaoUlabEVZoIxHAc2xdtXhZtnbsz1CC3JR6XPm
y8EVSOGmkASEiHiPSKqBVM0O+JcAVZ1koQHmymfdlZ9/oaXzWXGzxw8sO/k42Z8V
2SEVrc5D96Id+LSRanulUCAkR1NkkIsr/+ehif8+jRCz7ZIzfTEI1JxagVRtmeFM
nu/m7yDOmX9eW3Uau1myU/FpXYXyvrvV4rlU/btxxUeq5rPugUm9KayxzIIdwNsw
+7tnEWcrX1hxRG9bMUfbg616fnrbIOGHExTnjrworQ3kXZzx5h+aAbXzese0c04S
gap7KixR6FMU8BV689anEU8nOrqtXWVnznfGxKUmUQLQz8LsKHhQFB/16FSf6cP4
nxULdXIRfbnxIJPXl+Pivuwoy0PJhO1JSlRQbAYx1bi6EcOz9i6nOCh+oVmeB+QE
t/5XgBED9ke7IDMpuBDAhzcOISOM3VaxHsdpwtkPqjf7tHB9pLetcFPbMINjrcyf
+DVbbCa6Pkltbk8iCmh3x5DzrjjCegteIFUm4C/RBLIJMceblsHObKVE3BkPf2qw
RtVBf1wwjUUvrA844Pl11KuQhBKOIHE7lUQ92hnl+p5aqmCqzzD0v7kdpzPLoxUz
1o45KQPXAsGB1ekkFYVs4xD82dX82o472o1jvVKJBSQmqQnwp2EIFRiRDDKlCY3B
q/F3EXlAfTA66SevWVCA7y4vna+fT33cTeu3ooMGNwTREXAsOXkyvQSIlHwZrUa7
xmlrvVmhBqgyFN/uCFgSLZZ1lWfySsoWC2L1DNnHLjz5+4l//O80vGNwT83bCUJS
REPBXRD6W/sY/kmzcvOgOzDqYJn0e/LJxVOdAbY+q1V+Zg26TMQs+m4b0y2Z2dXo
wCVdlju4fGNxaj+2zOqiT4Dy9FxEJv+j6jjV5strIeRNYdpj89R5aGAqqiPRN6g7
bWucRiaAJq5sVT4OBpVcIPfCsM+hxtCJRagfiJywZbpKEmiGk4YS0LySSfxGi+Wr
0su7IpIi6I4ktsuP9rmVIVsxyMFszJIXGTUdCWnO71RTJ8W9Ryq4MwYcNXk7bDMg
SWFBVJynDsqBh6YTByvGqFVjDiLWQzwGom/8P33TRZnLqf3V+pf24RCsz+ZpjLxv
iXE4vyYk2BbvTcAywfWxT2B2lE8XXnIQTAPsD2Xburbf5RjupM2lLTm7cD8zJdjY
DcIn0a9MZ4DjtmNsWyOdPiPGAP1QFp0naA4V8bbGMHoR030B4hIgPic/iAr3uTjU
kN2i6PaBXOZKtqLB2iXQb4BtOc9M/2EBEdcgqfR58O+1uM6LDXIFPUGQXsVQXVCI
wMyA+RicuFf3lIHfClhkq0bZ/SguklzCgpIlT/CI2ji6Vj4MZ2Cwibp2Q9G17NL+
6T9e9H/kf478Uy79EiLOljPP9bU6LbzjEDcKWWT9nJ8MjE7JQuheUzoG1SFJXvDX
y4t82x+WqtD2sGDSnB6W+jYLT7CuqSOsne2I1SkXtk4gL9+NHxawpwkEXspixsza
rnCz7Ec6EkrJr+aKeD8/nc6U50szEhO0yK5qpjfuhJnCbLIiZAAmuAZStc9/k8Fw
iHtAJSo8k32+Jd3P6nVqbA2Bsl5E17qQVU9ZnEorU8UJrAZ2Z8BK9HHG9Htj+oZc
loDnZFsp9YZU6+7FauA9qu8VZtgwj000Nt00Z0AMXrxJvpB4yak6JUZ90uhxxue1
8yTIyNCk5ATbe2b3BNEAUtTQfJCNw1LIqwERezxx7XPkOg2jCVNq8ZwX3esLfmbp
RRvQcCP8G3fzjKoE6+WoeqsUwmop1FV25G9+tkE+tfr8V6WfV7hqXKywrsPGc11P
Pbn4CX/oGis++mNZuoJK9a/BAdLvintZbDHY6hOIv/TDPFdU1MuWhvlQZZL7GUpe
RLEmrgnNjgWeCpDK/RdptQeWV6kmua4uJ7pAjJX4IsZLMtvo22qG7ZjLSEuvhHzK
yadh149Y2GzAV8NjAbdM3RD4BBYRBsIehWwC2TVRMD9QIQWKUUy8fJ6NHztWyy+S
P6/HItJIOYqrGPzdrSSpPcvRlhUoxsaJVQuFFWLWLoibSpROCheVwfaYqxYBbDA9
HndW22qiJndHALKjEf0CjL8So6dOa/pfHhET3m6CL1Gl/fgSFrefn/LaQBEe1GaZ
Zf/uaH/4TmrjvQflUb9Vu2+1pY+Sgp3UqK+a4u1jprCnelT3ALRX7IfJjI+ryFs0
filLKU9fACPlt16nBefpHNk5YZ9mSGaXlf2VHLj71eqzqU8NNEaMC9mBSMVa0AUd
6McXU0cvMKMsWvN3e8rhdoiWveS8WKIM1j9R2Mwtgcfwt24kCPGm/0h3v4pIgnXO
ky8aHX2Q1canrikY7LPdwTHYcOXfb9bgl33IzgXYUVcYCHJbT+5rQmOJ5hMPrcJb
CeUiZ92BnPSePKFPHz7adt3jGiqvBvmAiC3Rte8HBcljkWf7L4nElXQ8pFvvDcoZ
/sbeKlD/MdLwHAKi0VlLflTsm6R9copv6vtK7VH/gr1wAUwRNIF7XPbw4+kU85in
c086uL8hdVh1a4S2avZRb8mQJuUaYwIsaSisaK59ocfN036fa9V3vmvQzdqskLWY
33Z9EF3GiSzLwZOmAWtyGf4ww8k5xlA6jSxdptgQrUDTnQ/FMQApSsTIZWeYg0ph
z8U+hg3o40sriVrlITHqJ7T5WxJipXTFDcaaFcClxlONs+Hc8bZYna+pIsZUjWrL
qGk4YarnWw7xYNmGIOnqRggi/c1f4TSind+wuA00Y0C0QH3S2nORDcatMgwiFGxn
p8O5ybr1RskL02GYlrmzFYa1ld6xld3+x+KkYDoXDkIeT4FYPejdkokPPNp4NJ+2
ATcafbunDD9D5CkOA5cP/JC4RpmZM2yAzGikMt6I0rInKg2Wx5OwGb3wIrKukX1G
cgpvhu08So2d40URFracJ3eznn8rAMrvuPu54rnyhlOMdc6bF+7kULbqOhKm1o8Q
utugwO3G5JNRvAp5lBJBYAIPHjeCk3V55PuoIqub9Wdv+hX3BpUtvcbXo7KPHQUP
M1T3aPjd+6IG0gKGsPJ+ZkxKlVmhrOnVop4pYi5V+t4wzFHYtYCl4JWXA+cimknX
6Pui2RRIaHgfv3DCVSg6iI2E7lWBj8Fa6lKzIPaK6AOiUf/NAPJynz/fagCkQUIR
xKZEAYc3QmbjDKP/FsrDXh4JUZHo27Ag1jYPbwlx2CyAe8BGzFRZfKqNY3iNqIJa
zbzfeCJmRoh24JHnKJgqBnnF79le4BWZGKI8tl+kQTW9PnSBlUCP6TqAe0Kaa+PT
+8E+sKm/RXUrIASf8GlGgObb2Kzvh3tsgYBL1Ha1Eeu0mXv3+dL5dWrQO2Nn21pX
UvEysbg3vY19mT4XIEvZhrdeXxjm5YVvNYohcgIodVgRnr99cmGkGkFvfwMXPlTp
OzfY8f/3fX055nKVMTv3I80hIbj0fnhACWePMcNmo5j/VdZumVXKlSQLN4TpAGjU
xdQmv+7+uxFu2W/txJf2L0H+sfXsq02Byi2sgYYatx/DjurwZ3pQCYAWBjNV0Ujg
lZZzlOt6BJHzU3Mr/CORBgI1jrpV+/8Q8gee7yioAU44fHK3J4hTK/gQq8YhdbLb
BIXALluUBO9FRDy9IWxiVO2emrCX7AxqPr9zeqZcOZdFKsfX4YUIEj3K9nTNrZZY
Rc2bqLYg8Jkr/tSc9FUePXVRp3i6LhfmArNsE8lTzC4eYNRbG3WWTiNIPODGujrb
nZIMurai7k1w3KzhhmgJiyaFdLbnLi65tWU5EI/Wmi/e0VH+fD0rPvCuoer8Srkg
Pg9F3O5RthRPuo+i9BHlKqEnD/YmawHkHW2XObLgVdFEa+88q7lutvguHA57TPlB
WLBIZr3Vfdnr5ZQ6kpjHt62PuWS0fV6RK62Mm7kgH7Ph+FjDFIn3IQAetfTo+lcW
WbFzUrkmAMVyN0NDT03ojwpN7s3Q7mahlaC61ZVLzMKQjTnQXIqFALqjjKDEA2of
j/c9+x6z2SQV0kspMKaNH/nq9BhP0Bw/j5MURSyWr5z32sQJHLL2phD/WGX25SPr
mJo/Ebb2z6s1B6nElQcZZW61aNhcNxZ5HTvw88FEgNoXpxfXcBsgRMtuCMG6EzMP
VvOnk19LhVChZLZCq/ffAdPD95worjVNMddm1Hjjp3of8UWt33CeA2BvcvFO6+rH
nlsxx4tjlio3ovsVFDkvT1WdoXq+kPJnQIcVo4Wj0ScW2QnzAAF0rv6+L0t99WA5
Wd0qPlF34scCEvvBiE8FL5FVhCvylE6feVaynewqp1xoSaHNE9wJDs7bWmA1o/i8
SLJwzZNZjsnzUurXCTaOkzQ1Zkv+MXGngZq7H4lPOGr4ecC7Y2+NYWxSvExZ3j8i
+VI8oSeyGS6Iy8ZUz557nohWhRAMUQNoWFqAshCyylNvrlRb/oGvgMnvUJjbxCBb
Pgc65V7qhjqZsqeXyfVZrE0IhrHF82Ln9FWmm727rXuwN3RU/9wvOJ0+zcvUAJex
JK2LVw/UyYy0+7uGEP8zIfv6agnw11FtGGxLs8R8on68JWdb+wpSWnPl+f68qbKQ
cPnjE4I9pDAHScs4TEEhG4OcwqkS0Fan7XDYcD+hgyUca2BiNOqyXRVbjfWLxfa+
lTezNTG5YsO4/vTzeg/weainDgGz6xyMsWWnk15lIQP3vuJXpJ22rYEVPU6X0tOP
JAzS9twmGG/YrEHNYkLc+sexjK/f1eJ98zPj2yIQzbrkNvxlCVClRDkaY7vdc+NJ
NySQteEPdIVpfslly0DPjKRVZffVRG/+HzF7F8gRervrykY9OhW+xcAqKUOZaREP
JU/TnwUZC2j+WBKZHPnEfDdk5TJRpSZON4uykn1gAFvxPDgDWo+AkbDxOUBGqzsl
5lIEgC2Ct9qY1nB5ul+k81XL2QoZY4q9b8RYQp6SkmH1VINyIicl9aa85UKw67rR
gKFEE1WA32WugXzfHE5FIZhOQX9dhnPbV/Y887gvNe+JCTku8/yDaY1DabdxsKgk
WypJfgLAKsPOZnnVeMN6EokKl6IM1c4MAzqPOnHuTLkCdugK2De0/RqgZpUDfzx3
/Try8QPUQmwXs5Fkbvix9eOMPHhLrJHQmH8xrr0U01UlPysSw9djwXFbym/kICtq
wnl6mZH46ll8BrnCEpr7td2b3q75lide6XWbfHHOJvmuNAHd0Mepmnfrjy0D3Ywk
kbdAPfas9M8hC9wRxEBi8RrUN1NV/85HCrgoxQ5NoP2rBp1CNzXuy4i3qGXnFunY
QCYDqOxxLGwtPzHJSR3uRjxonJhNpVwKGw611h+BGqNWD/XWCE6/inCEMW1lCgiA
XJJm614de3W1HwXV3Rz0MtcqCLLXkBV/J650teb+sS/M/KcYeJMyGsnTOTSmh+TL
LrYzXcLVgi2LvH4IApQnUuxej7Zjoem+JEvwyXwRdPE+YtH8GsWgKIS/uVo+s04P
PBD67VBGtVf9ETRjf3bEPHXHzPHzOAnTwp2I38dAZKmhS+1qh/fTBPAtPoxpWhT6
KfZfcOQhdqLVNDCiHExHhAug1V+OYAt4+6CscRs7PCeA5TOkVPaPx9ovgM5CjlaB
btU4nPhliKxR/umctNDoO/t8LB3EVqIYyxsGM6Ck9e2MXKJR62Or/OIQzyw65o1z
tR39wVKaR8HocQ5mNyJXa4/oWTuJweK8UrbdMPLwqMwpFcpll15+SXl4yAYfNZ+g
3vW5QKS00wquQnR4+qYPXxuOOexOeXYWrE7DRy//4eMcYzjMqqgbogSam+XyKeRs
49N1Vm/J+E3UWZ+4O72V6PO9QPQXuvcSRKznr8kq2Be8mvfd9p3dFKMqcCxfqU8X
0BWJcI0Pt1F51mJEDzho5GJW1HmWq3UvEOb93Dt1Ojmnty5qwR7r//IDint+3LN2
jubyI+kISYy7mT7vz/o7VXwcm/do8KwCCizxGgUCvTz3jhVdi7AKai9wZrxf5MCh
lkg6qGPrHar7OtiNuG5Tf/r45/bhyAFs/BnImYGBj+8sTBJGu6BdAiH8U9FWvGyW
lldyvxtymlbsv/GaFSSTwe59/oXlv6FNyAalh8LGbb3VJ4fuL8tqROq/nllg7Edt
v4dfknGMyqTS1KUBOJw4+6m9SrdZCxqUseOKThg3GsB3iJl+klzfhT1TKVU5B4nL
yY+VbDSvcScymhQP00wMQF4e14Exp+n2Alnx6pcBaSjSnNlb/ryg2zdFjEgnXUrT
LYDktTZLDopwfLdfNy/6bls1mRXGN0ZRE/QrjQr4ESG8PFEh2w/9JxVRLuiAMJpY
72Utlif0qUBWjxQ94KjDjVFbK/13+i/5pTuXcaxp7YHRjWpEENTT9J0YffRd2BKz
EMKPbFv1YdEpfcRuc8tmvtBIJo8a0vq28qUT59g/SqPH/XBzvIYUYWl4unPYDrhf
GWJIMvtrQjeaiPXLVMwKrLDtdP/D0I9QLkwiO6IjIwzGFA5P/5QBtQ5xtwBeS23u
piZpao0UYqTfrlxgxB311i1OrrdCMa40Nq8XXl5sljV/xxIOIJAg6DCY1PD3GuDP
EK51NvCLIQSQs+STJ377Wfecg/HUgUcfZlx7+TUoWiNgF/QgtcFtoY/TKkcB2kVV
8ELxGf0w2Thtr8OC5p+fAQ0vfdAZ7SKiDxcKX/Hy8mvXoHfg4OxLovw2moBjevaq
ZmRKMLABd6KxyojZg3DhQurpXhwQ6KDpQK2Sb0qhAHTaKfJbL7mtocaRXkecgW9v
oF8Um+d8qTe4WFjuNaGotnVvpg9iexeW2QHJ5cDnHof8DMASDXHj9FjHj7slbFZs
g2SZnWKaD6h7PwQIDhTdyKnHMqMKFhbwd9mnRb+iAFAqoJ31jILPLk8CCmOg29PO
xYFQfl5qQGBK9dfKm1XDCj+OyvIyjklmv/n4pkylAmxWOIGkKsr6W2BT6t1hN/4m
YrvjcwSknHueO/K5JgrOlVdMdBqHOtN9M1nGH3yyIWVZ7bjtrr3PI0FYYT+ovomv
GlXOOaQ451DRfTE0Uh7PH89hyho/NtMwWBW5uILbqqeIMM08W3E5xE7YoSNcpKiu
8t32fSx50uG/9/T3TNIjlawy6DIrEDnpuJ5qVZbXvzLT/IQ8C95IxqIfFp9Y/ZMv
RZyQyytTb4AzE2bK93Z7X1dzEzE9KMGSL+sHH2iK8NtCejThg/tGxVIsHGJz8QTi
TSZron7cdLT1EfwPd3qx2nhs08zDHUC+XJ9GP/OkDIKZP18Tt0Q67SHApiL+Diu7
oNwlQSmokX7MVa9hxFx+rT0tmbX5KyX6UoQ/552pUItj7srZATxh5csXcOg+yS6Z
l+sAiMd23FRnUPmGV95FHKH8Qjm5QjD7s8WyN3zOuyIAPerosMPaDfeh9ieJOzYn
cLov6//DAct4f2fQJL8C3daSkCBbywhoygYmBxmH6/ihbRvbi2ElhoFV0y8OdOzU
DaEQ+2eTy1icGXd6J6Drpx1QpVSLG9R26jl4Zft4WrqvQg6qbQmJV1z2+1my0F/6
yeorsf6W4qZSm885uA49ygOwrgCk9DLVdHnelKtmC+Oa9Mfr9l6B0St75qmJhL0x
vOWyJq64hxYC7W7WvdnqlD8N/VE3gab9bZuw0Y7vj8eE1+0LllSwxhrIy8YfolcM
I976heboNpzNhwHH+QHymG6+7CEzyq9pFG1HMfPtD4PBW6e2lt12fkWLNOtJfqcC
bxItvU27w63riYDfCGrc5t78pm23gmh1b5R8z1b5aQtHibHPU9e6J6JQ4XMsFO5D
R0LUfweahct8RLBrwHMmmFAh3e3eDE5dGfAiZg+hJgaNs9yBWo6pNtmkwxyunHJU
2qoLD7KI7F7MLP7BlxE5JksXmifS/SXoicdOGTbsNXCr3/P2SoPZvoDGv9L1m/Kg
fKnZmUxTVTcmd6DnvzWPRnb1eYOoG0bJwQ/p3lgrk6/RrWgUwPom4fjTc64uqKED
ItyAU6gIcySc/WpDuuZ5+8IVy0z5rzdYbCSA375bAg+NSGUwF7LhZWbexbM8i7Cd
LzXOB0OmhCdrhSMr3I+VJ94UUKQUIQgH6YojGVok1dhaYdcDJsHiCqq12/767gvW
OVHDdQxsein7jUALm/yqS2y9GQJKyEGBfQEsVpNpMMVLdu0+Bk11KY5KU2hClD+A
Z/7QhiDIekR9iKnL+OMLBuIaJ7yfJozjthUCBgWSI6bm4m/UmYT6grbp0khRZrR/
6kcemm+rS0KrExfY53gHz2/NKViCwaSz5WE5KWJG7IiLC6bcI4+qh3lnMN9YL5kE
31Pgq7X8gJkKajUrowqCEJr3bJBpTTHVteU+pznJnYkAstvTNMfa+81wRWs/3mjf
RVlFBwudJ7uDtP+Zsp2q3DysaFoZKbOX7LPI8vrFowriRwimc1H+/c4kHC7GLmVA
wiHmWHktFk0E/4TP+6TPK6T8sFp7TYWljVRCMNibVcH9/C2ux5OZGg8yltzokL+a
ZHtlYb0qdW6/sKMlrJxyqEDszsYwNqyM5tluRLuxL2THzlApsbpKQKQ3com3hgBk
ZP+mrNFKXJMWYVawpF0stAQNq8EluWag8QrJzS3uX/hO1+xdeMpHJXGmHpmehsvh
pur2NMP19phUgJX0NB2niWnNduWMSFEyIBpZim2v3vXTDejWA4LEVJpefATFsBH7
63VlqlM4uDZCKF1s1kSyoHJwzYqfRQA9UC3UZrLbAcMQEEumA2WCqo5Nrqa0xaMQ
/lngpKv8/7xcQ1auoQixrt+MLzykj+EZWE+Qz65VZ9x0VXXgb6C1n5H6Yv3AK5/D
7Dx5KXM+Tsee05A4rEUm5quq1+mHCzvjyuFChyTRuoFhrcfjIZSKT3vCyAltwUCX
RLJ7UMRtRfbqFrMznCWSRQb2EEdS8tgCbzt49dvZog9CwtXxSwhBi+v9TlmYqAeZ
BppvPFztTns52WCVomXdxHiDNIIJSDmwr2pQ0Jq1W2oa3JlqvH90/aDDb4pXrxlE
RZNhnAh0MwuUMc5lQ4rxESp9yvEaCn3j70LDvOKPB+r9jaqSkl3Bj5HRyG+WGSEu
eoTaya6peyGIILA1/J5IOLmfNjm4iSzGtr6YHsvE31cgrUb7hYtWAKQu461NCwz8
5J3raONM+fnGiYzPLB4ZvINdBpJRO9njl4UGEdGqmPsBZlfZL6cfbQPd1eBZDcu6
aoO4f60osqfYb+dx2OUq9Ow6NCqe9HNgBIQFe77X0F786/GqNhbjt8m0pm/aUHLx
uI8CX8NUksr+VZ5MbNVQOPoNHM8NN+j7P70ubGwKkrkz0bAnAvse/cj3rbFwvIfF
eZflkTdSFl+9PRrCRY2YDuyRpJbc1G62dxZ/Uw32mKQzy4UqbqGA3izFCZsLlV3z
6tkUJ+AS8X03M/Gvn2g8mMOVMadW/+8ep4OCiMQ4Anxi3UCdRsFd921YxQ6XyHMA
QcgFPDd/Wifzu47/+IO30V70ixw1OC9KfocXHg0ndyFg1F5dWaZqwVoGwWhx0cYi
h4LDuCySj3vdSQE9j973hAtigkEKKUwXciIxnKtSkUHIn4eLWEgXI+XBOijEjL3u
GotkOjAeuDnnTa8yOeq8lxrf5GBOxTa42lOpQ1xwzwjUc0KYdAdNbtybfaNZ9QAv
/yIWbvSsAaCeMKC3eDw8HRs9l1U0QdAiEV6w0mu1yFXaLCL3cCKDrYZhdx2039zQ
7mA8HdW78yjl+0zXYgEQNu6s3MAH4WYOsSU9cZPKUQzCU0vo2VEwrReqXPQU6KgF
/u52QyRERtZDSUTvL7je5P1os79UKib+LzFtvJHnxblbKJHwW4x6erOGxpnKOzlE
ilQ7PzysrC6nNixRMF9zCwYnfBajXSJ1TmUxVlT23EAvq0FS/AuRzdYo+h6u8n98
b7Hq5vvC31ouoi4ik3kcKHiEIr/P+u0IJg+vNeUTux0jQhlM6/iWXQcAR0ar7W9c
veIw8o3hkRXCFXGgL1DaKp1/ABgRxEDz1XA5/9yJUtnZWgVvWB77N5WBzUPzxyBE
71Jqw+nqZ5iczbbFqjRTTnwTGLkEcPNM4eNhfM8GzawDQh0yJbIW2WZeFG6Ckqc1
R/rSPmkPP4vum8tv/sIjfucbvEhlu/vEaicWOpdaeT9FN91tSDpaJaSP9b3mUorO
wWwfVM47uN50ROXLYzcaUWVLhHQGuJMrIiwtsQ03ncMqQ9YaBD/TYfzXB7WdQldf
2if15hZz/Bmh0LBe3RVFBRvNs2HdAUSc0XJs8wi+N3rPhLTe+cHaQIij9mLd9VPH
0uDjotrhY75kMiJYRnafSI4p+AmRO0MCXiawBIwfw2Ug29lPcl0i6o3CiRjPajaH
Ax8APEL0bc/Df3ZhA9/pRJMcIcjle+H2HdxhUJ746ELf+oNe9T0ZN561OmgtAPW+
deJVtL05EdOdSCtdTzwUAG+gBzGVD7eft1hdaO1CaZxAaIRLK9nwvDhdQFyTnKV4
9+vFZ0SPD7sRBFuRO2YF0dbN4R64IdZoY7JiBl+nAd1tNiJUGnvcdnVEsmhgZMVs
EQbf8qEQHjOIFUEiXzuilup+92HCOtcPJk8FDMIQBCuEatjZoQx1C8/kH4UveqzP
yg78CfZBA0q5hkSx5WttsZ30JOg1c+TNGiJbwkwN++AaMIzM4v26tv5gjlogkayO
o6704HKPBxndv0mLq1cX/yW9xbAQyv1u0DyVHYlYk7Fo8bOXyp2iAxRgrZvwIJZm
Ah4F1MlRxU/XACPTiaDXVBw+Q07wgZ/gMo9LHNFXZPQg5LZtLEYoJeHBexr0U0LT
3TqAAuOl5e85xLQyK4mUk+MHBPk2WlTq046o4oCSJfWWswMk8rMWS7+JaU7VRogq
w6DarOfRHadqDtCLPt4Q9s4KHsdERZtATI6dNRiUb9ezxYqyIFprRdvYJLQZFdnY
ntw3qs4jNOeKr9wif6rURIfqqSQMNe5VGvNbRklq19cmAGwjwSwJkUc+EDjODpsA
txpCdFDwUisnlh5SQH3TNhouGOQDz3vSkihYp3/HUDUGZ1zyuTFXKjARs80wP4TE
mnkFxHjeK8UAva6eCX3KPzsjWU5XXNTAD7Do0u5FccbKOIA0lxxgF2EIm/aRz/A/
XeTl7+hSCSqvRip/7OWt8Qp7DANVZsYKuGj1rv3FZbygfKZq37bZ/9CRMofSpAIK
e6EbAsNvAefVKRutV/9BHskoghmj/pIDLdj5BiJY6tkPdm/ty/3BlcLdRR7oFzsE
NxQEeQYtxFkrJopr0If8SUAmpf077XJWAktCu8A2QpY08DVJIBHj5On7yH0JV/f8
mQsJYOfhM02Le83K0+ll+es0rfAvKxZp4d2KJovfrwVPV0cfZfpIUb5pCiowBejY
4IHNb07ve2xYkU3foA2XG1MEGu0WAvZxWGo5ju97MpExZNoxMdOZNXsiwFzX5gaU
EhgYKDGPL86XQsifzqzjlEt8OzBHtezE4cJICIjMNuFQ8f1H6n44j6bdisu9zvRk
9h8tc1sPRMtNn1Yc/lk+zFRp+7uJXBc06rYO1s9X25GpWqZ9Ez8M3c9f303dDq6Y
ryqXktvTCEIDlmcFndSL/Dftqu4QTEejygd+ARqTHln4rbYqdXTlAYiqFCghZe1x
lT2k3Y79yv5hzKsCWGXVyLzpG1jUaMoxj9Orkg5dOCxl1OClKuHZMEQTbGYyg1nb
kO9M//1diwsdz3tG2tlrHQkZAArBcvJY7kgG9JtLTGPpA+l/hPxkrKCep5RuXUqP
U4BN/NdIW/Y1+m/GQlwaodKwX1jYvKObdbayNaHtt8FHL5+wWqM+8CmGX26+WggS
O0zdsElXJPJva3fEI5zaPjE7w5wtx0oDAR18qUvdto3h/8SWrcOZnrvyAPWfm3IJ
8nG+OiSSFRaQd5un3Ketev3WYxl1Bmlv0mFlgBcJenv4TfsJcWwyzb63V5YhpCIu
bF048GsYWVagrICBs83Tdh9Uj0TCgYsWc7fnWx1dmVDI6mhoxSonOw+E8GjYpl/e
0XFqD384g+7fT/T0CnZqxLHLj6rIMOTeTPKp3YCEdFvliVY+VQjXAodAaFA9bkfZ
2aZ0/1UCxBfqu881U9/OL0MyLoF+C93HdWe2f48d9nQbiRHKKnnOhAYAkwB5mXK6
PKzc6x/LkGh3sfDXOBPpCkjG51Q8JIkob2/YMk+2oxm1Vp8yyL9Sp2gTTGuuSgpd
9nIcJf1UBMfr60bMyF2LzMK6gYlMZV528EpZQexa/+flr8I/PUpd+P89uOywLAE0
sbCzzeB9Pqjg6Sy+eK2PEvobpwPQejuvMBb4K6V5v+0XdNIMJx++PicgtD+PkGmk
3HUrEPSZVEzHUdAzKDOIf3ZGM67d0b0i5miBt52UtEDGViDT7ymkMn7tu6h5PbKW
sTHt3d/YXQdcZQWC8SAOB9uC4DZ8yMYk2KthIe8IKE2+Zypi00azPqX7+P6WHy4E
z2tEDJ5BWExj4BSMMKrEp4WunT+Nr9LMLEW4NymKWi1S2CE5MV1VadPoNJztgCqf
IsEDnXR/ZVXExo0j9DyXtA2gDjcCwqp1Y22wH6eIoF6u8zANhTuRyTsJnlG2etGK
mMdAZaMsSTPzG61ZdhONESgmw0sGLM+9CRVvMxtGpplACbgmUuaSwdNpe6BkilxY
IIqfxz+/wh/2oZ8ZumHQl/6bFG6Ior3ufa0gyxqe5pOq/LHjoIhqKHOGfh16X7Nl
cSK2xUb2T+GYbRUlZ4Obyl7ra+ND4MT5PM0/gvqb0QbpdB3M9Rv52kJWJANPujr9
M/CXIY5Vh0vK87eGH/rVtNKl60LHi37lUjKUs3SvtsH4gPMMhBjyFybBqia8IMc5
cn9yYFWr16Wo5wZeCvsDAONOTF8J8uBeQIsRvrVyhE3UwtAYEJKqRR0kSqWT76y7
c20GoyV5zS2U/PO+4r3WR7N5zPJWRuwBZXWJdsnmbwtfrWnlLIF4jg59/5mauAK4
uDRPOUgjr0tREXm4P3R3O9hmfsjlyERI14RvP5P6iZ75bKm9CKPdtFvPK1/3DFy5
mTFgLIpEe76l2GedE0RD/vfTTP5BLzwEinJSicHIrUkQBVGLHFY/MrZnt+q/vXhL
4HK4LSzDAODICvnmPJo3cogFDszigI6bHgUr8UcvgAlnY64ZoK7HpAUZK9FpiU3k
4Bm6ELgi3UhunhyQOQQi9RGVt6HDOQwk2gbSIN/oz8o16rnHiLszUA2XzXoUbI5l
ykDcKKQpee7pvBxFE12HeINMLm9IlbZ0U7LmEadI01zb3wrjxAbZhUyjpJY68pCR
NvB10gvAaQqqFaQ5KfFYlAWvIGTHOut9uIs+DJJDPz+uRDJh7U1VfmyZ4Rni+zWI
Mqxy9t4gIp6p7Ck6yfrCOiTyF+B0QYYjX0r3Plj0Al9HQTD1ZOsA/bax6RS29/I+
D4FuKqxI6O9kOSRIzss0ds4PMVDJPBYOt5LSS0ie8lc+FbNc/TQPrlT2TLAU2gQ1
dNAK8vkVeCeF/62UPOqSFTFe7tWFLNB/AgzVF9fU9gAQ9kMB+9s+owwGwGIl7jvt
d7aqlBCcRf72E5zZCvO5UgmZLvXYxbvaq3WvJfEMF1QySv+HUIKQ3z5PDlQKOOqc
9JULEAy45lEN6pBVkZeJOaXrl5cYPMY6+yxaEemQXihDXY94GClm1d2RHTNykrV6
7KLCm19GYUzOibOViISKv3Iq4M2Miew0YNNTcndxJcbM/YEaNfZm/q32hwhkCY+x
xXNWbZMts4KU7C6ddId1XvCbd+FLpNeIhxyd+k285UN0jv5c/+C7NMu0NavvYMMa
busfwcg70+pHpGKS1mweeAhB+H4FzWiwazWIuqLnFVbsJX5vwXNUD+wjTQgTHQI6
XNL/TF5ms/h7GIAHr/be2cDZc1i6Ni3i8n3O20Ds8TWVPjhGX0ndBs36b2EuSQ68
jP+qWStN46igZpVzFqjboKZTm0IRfKYRMDBme6ClS/t0O26uz9i0l6h6yu2fpLIL
Nf10ScB+kc7ZxpRfX8yaa+aeObvDNhi3rVjSXPTzJh+CTlsMNSB5TWBpuxsbqW9X
FhLVw1GtoiFX0ykpwlvXmVVmA8oG7NuOAch/L1BFLWa/Usv4mEMsSywDsiUkEW0S
CrKHdv6vJyPxByg9yRRMN3EIfdM7R0RvtRNZ5cQVIcr91isA6OVI7odAUo77QwuN
FpW1gXdUPlCW59OnTHQcwHzcgaePXPF29XEiMPQSazvE2ORPhOodZucoOEEtKMjc
So3MWqgp9UCuZzRIiaQ2V69NnpwGmseoElPF3IO5X1YZav5wEoBHDLMwApbs2WPq
VUCEroSzLaUi8nnNmcPxJ0BXyeda/baP9yPLgOaxfwkTiUGGj15pFiTNCmNXej00
/Y4gtOFOQdQ4+abb5IpsslVNXrzpzZNPSjwqe2gQcO5PSeai0JIdDh73Fm1hVNF5
XM7dzgFXEhtgyO0ABSsZpx1BouzIwJ+TQ+kbybrYMxViSWxuci8RdVsCoxr1Wro9
aQZj5iQ8K4jDifPMyk5q6zrs7DLumkBrY7tXfo5gZPI8oEk3rrAcA+Q3S0R5w2D9
n8Wb4Q1CZLjxiHzr/0nVACtYbBMTsfCegJfwMXHca+TblxM+vSNJUkhwWP0PpmSB
Twa4PJhi6nBhlvml0dseq8V0cwS8AwWWHkzqPpd5iZC5bAKw4adtWybMaIRd3O8p
y7vZTi1qVZU0cirhUYvZYraX0upIuCvd5qeFwuSaHcEP9CbPKfb2qx35hCfqzNyb
hBVjqrJwU+mtdiVtAFe3EvN0+hyKc+3KW02i5CK1W7vhoLmHAmlbKDpBHOAKrZXk
UYvSZ2Ds5YKRue60MtUrANQPI7TjsRW5sSbj12XH2StouZLBW12BDdbwJjp+PYnX
O86HOkcWqUjA+m/AYpjjMMLcX5K2ANMo8WtCKwCD9beDPOG2fXJI5rvyyHRX/dcz
On4dFXgHurS4w+H6/GSSSfqFWYvavWjQ4oS5UsdRRwKFcNDzb/LHWSn8g+EKGhsk
MIRKc/RtKH/IUS1yJwQbvl/AZHVhYdEQj75S8FQ23Kzl4e9FpfptCUBSfmcmr7Py
o9jkQQjni8gz0FabI7GLcNvVVWXK+PfwYgHL1MqZVLYDYpY/DRp4P9BdpxGzREWs
DUPH0/U5Sp0FR+TfBAM2Mlrx1NWHBjdgq+QHfHQ6bpwxa1tS2iaIXPHnDpoeOGH8
9Ucxx5DrKJ3Z2Tl08zx+hHo52Dn751jiRpICKoh3e//i3cDO+IIFdQhP5dRvAu2c
Db/9CDLt/XR02/yCwW/hJ0enBoE7qhCwrGbhva4Zp5Ej8tVA9hh277MohOmuM6+i
Rh02YGTbtSXZd2ZNhFMZ0KiGmKikG+d/LGyU7c8ERvUrd2VSIAj231Js9N/Ni8M9
HCKU52girvHZc4jYW9r98CT2gbi3dt7F37nVC7sGUuON4JrCU+1A6DxQ0k01WHC1
tNCDCeXPJr+orGQLvY+bhdUSrjeLOHtKpQWoZkhOcyNIxSzST85PmNWtvSB8s3uq
K+OHO0ob5JLH+y09ZPRqQPia3l8IPA/gQ2MoPhQ/RSLhdpHSEF36kLiwQB35DWND
r+t7BdjgTjXW/ifGu9NqPGFMxLzlGW5+NEnauE23559cUzKdUWKLpmI1PE09dFTM
KD3JtuzaMrOE8jaUcYKWGvbF/fR1GULc5ECu7on4xOAwzp7mSB9RF0k28vIa1zDg
0tQNyNYVd9eAohVuro/9QYjqQr1AkdfHL0bJfrLjUFIAFV9aUGjG0y3Bu7RfCcap
PSywkCkA/gwSyyYMClFOzPbgg7TGbtnr9r/RpXs6G9gskzOT48cNQLZHPYYGllBK
oz9wJTr2yn/QjaI8ZFbqVmzldMWK6lN7CtmlnHJfkkkAgn9Rip75ZaDqdBjJCC69
zdsMCgGVil2XBjr16ZG8qFq0Sjp+BXEIkVucqenzgj5cdmMHS+337FSwBioZbbWp
nxt4quTgovq65ZWrlRlQXm5i7mKlAHfOr6o8LSL+ivyKyqYQv0KF+dIicUoDICxs
ZLYWxohHepIOyJQYOxx6iYIb9BXyzARGqpn80fLFc7yM11h1N0ib4Lu0tkj1Ylrq
SLNnkvAmRLjX54F1xQh/w3UakqVxX72Z+mI344cPm9V0XZlqqHT7knHHIeaXpWIq
/gpxsQGFpEl5gvxB3EWmQI//w8bfPET0JklJyfRsL71tX4KBCpmot+jrL5A0lUAT
R2WclbwZWo3SIgdXES7s5edgn9EEAqUB7RWOx6GZQRLVJyjlatgpWVWX013q5Cay
HRULDgaqbSkL7OfBMeCfPj3eNPNDfN/DIb1/ETbJ31clfOiuaJcB9Ghfm38sYMBU
m44DV5KaQVCekPWOqqW2HYq1b7FefzP2DJ3N8qsJf6v8U41y4po2pgQ6o4ovhyF5
Esqm6Ccu9kigADTRY40Ik3D7dpLQrnUbfzynBNzog6YljElcDGOyZZbUPNANKLit
4xSITMlmIOCKmOIyAXfN7hJgEu50/tQIwuWT0dpJjvJbFVqmLqqTnaNCvOroBWIL
UZY2OhEt2QHrRu07K2sk4e+80rjzJpxFI83lejHNfAioFfM1tA+vc/ml5Iu1gnSW
Of5AcbN8WeeAKiG+jqqJ1hDIv9MuukrA5eOBaUMu2X93lDNehT3r1FBJyGQI8lsi
iw7MMH3kInv4/rEOQJ3aGcnmz6sK8I4PpU35MsaY9adRy5kDbNiSv9ckG7Fd6f9D
SdEsanQOJA79LephR5LNglMXAGGZyvDUyxLVsqCnHCodXNig1HnDZrVIfLUULVPX
w1elRSj83yObMN9OuCm45TdCNGniTyeBj7Kg3Li3NnLGYdc+YFzgHSoc8HH1yaCR
QK9AV0tdgluXz+Pcam6udvQV4taUvQvk5iSn9IMsMVWKcoVFpQws/HlP4fdFIGO1
lMvFha9njbq2brbALxaVL6qhSlcmD7ezDcDupcYU8YWWgzqGdXMDTaM66wMluFVp
BGA2N2PQTqVtHEWDuAuZgXb/UsJcYY/c0oQ1VnmcsaUurSOAGovcBotS7wijOZVY
9E2wKsdNnURv4mtsmpC2HcXHCeh1x34uPt0KE8fRpM2BXWL9WCNf8pe3YC3ImP4d
BMJuX7tGkVgElUUPFEtMC8lH4MtwhaQI3e0+Qxo2eEuIBBKx1HfmP/L3pisd0zpy
24rP7tgeoFoq+kOT/JFqMUFzBjf9cIQeF2Xq6Q4hRClzo7QQYwh+E3B06omJLitq
fHg1c2R78HYEB0LlcylDgL7KL+gog1yVtYI7e0vUvm3x8Swpo9hswLhtW5sczD6j
/qzDjwJ/IVYI9xbKVDiPHDjjv7NOslH+lD0ee6Kg0oq9yYlRL7zlzz4KqFcm840s
0C655/LQElTNAeKEXU8MwOCDfFnVlInllAmieIpb47oEfqDfHZPoytq5L5OphpVa
zD6lC9gDAbYbLIFBxbAggpOjSKyBwJL1Q4tO0nYGmtHrwjZuNC7VncLyqSm+IU5H
eJpRx4D9YZ/zXEC2vm7RKrBJF5y5O/ifMSK5sbGBad9EXrE/J3n5J5Z2t8gDVu3S
z0OwU6FVilTJulLrb1/OreEChg5sHN49gafa07Hqd/ws3x7q5hodqsTzNnAk6AHZ
01r37xLoX1OVCVwISsqwAd3c1duHNBATW1h2/gmtXX1/tdmDkwS2pq5HWX6D+SSI
mpSbCe5TbjU33owdPagoBTEtYpocBZSxPuqMlR0UcCSidnDjSbZ9iLyfvtlrZmq5
mpfqj0NlYvpXRdmVkADZflZx5EqH8ZuPihE18AMTQK5VdY8oNIkMGLzFjOkmMa63
PLoki/mm4acEPCQsBQ2Ih5P1fY1Pl8EZYue7NL4BbQdGClMrfPAF1TLmmASp83aB
OHtP9Mv5hYuYeCah0fxjw1gxAd39HpsLOTVEY6GPQZnApEpP7eM6oEQqvD4T/cPo
XRlBQJFj/X4xFiNpx/SVzYaBGilPDNdkcjn1o7c7srnrgeVEkfpbv4aWfCnvKB4q
ayeP+IuXJy+1mPL+f5LPQafX9+l10el4JnYmPt2AGZkMYDYNnVD4vxRmoOrsJyRA
8rzYkpH84pav5rbUFlZAPNPlINUsXGxcoriLSMkmDk9/0CLc3ZPJ3CRSL+7ywZK0
D+YDv+Dfd9BYVwOvdheG7NmHudjH3QfEr7hQ082viPElrrYiXbXvZnKPKghz808X
tz2xZ1nVW2avbZWHPPy7Ao0FUCq/o3nUn8HZnHiyXSji+umocoliFzPaQmefkA1J
HPzjVXk7BGfbJ6EgyK0M+aTZnWfkf7VZi78p+0g8Qdm3IJ2W6KzcU4/5daTFsrEt
z+vWGVkB1o3aRyIeInZI4pKq0kK/B+ISJsA36BjLefkqrT4etv0K5kFFIpITlk/p
NIW1V9MtDoNsJA8N8+kmgE8jYzp0DT6j+UDtpiCH+O6KUCHaWo9hHhJ/XX1h5nlY
G67h2V5rv0+ZgZC27yIr1mCbBTXJZxDbXVxdShRnJ1QySL4AqFT4AbzsaIbLCKs3
9ozZfBqhyVQAzsQoqCpGJDZ7jaq7bIrOZczhyYQgTirqPx8sSMw6dHx/A9ZrOfnA
1nK3GFrflxzsR9WuG1PQNd9y5enT6SCRf1j+eg8javpdH5rIfAPzdSNMDda577/k
WtR2WNrzCcvvlcQvedR2E6F0HSW2ZXl3lqHuCnq7w9TMbmnEOH3s8hjhQG9Z35oU
U+Yj8aycdkXvwse0G0Bauxf8Po0RBzfBcqdz9DlsLpazmYbs23wpWf/OiY/UEqr2
cn0AVY/aCQBjtjAsfFHv462k2hyag5Mt9s+jeJ4nRRsXMYnBKfegmaiVPZbJ6E+x
B9KlvLdcwBXRH3kIjLnOeh7/1JB5cQty06I0vvwjsh7Xm3C6Ly+Ipw/xWwP0qBTC
G3Z9K2pBD24Cqku1rTOBfMCmccR0dtO+wDxukGuNBWck46/HlUOGixwCiowZQVPb
avtXJtpirbJNt6LufeGvDi0bjt2dOxhgaZKn25k+S8Uq9/fMCEzaxxDaQEpeNPGC
4qcbN0lOiZiIJVFVe1tx38gR0e5q9gNsDTVkfLyt1EkKNkhgXFlO9CSWGDXxlvV5
cQt8tT2Pb4Rn4h6f203z5yYLG3ZB2Rkk1JGI7L9lA49yCRUAFAKK0nr+XeWbhF5V
RyJ0IujuwnzO0ZGigXBA0NZMK46F4YUSaykAXfWTfB/e/ev7va46cSR/AdEITq/0
I9aSoG7xHMXXBL59BQccrImnrS8vpKAiOXaMgBESGbhb3+ft/BEYu9R1TvkccCt/
TjiVI+8aVUVCWkwEEHiNfreDwylAyNhoTOahIbeAoS4HuLrw7tVqgk/WfBasOOU9
iDAToGZadDS4Db+hUrUzSgTXRGbfc3Q3vIprdaXt785w43tidOWuxsB+UyYZMKN/
nJ2I39zRy2P4l3P/w/xjNfMrnkjDS/NYuWIm8wqa4ahtwZ98qtnZuE9HwTXAKZ4C
SAOhIgWc/Sy2/69MD8IrrtQpDxh0UQN53/397Hut6vZXBRZwJr7U6yydqMoI89tH
EeibA1doA85tIcbeMLyZbQRVgbDAAU6I/EbxY5Y1ZR2kE2AhJEiXb81RHZQVbcxh
TSh8W7m2cB6LpDtvV51QuYYOORZ+q6bMELZthoPT6VMdYBM9b7M0hXHeuFPbyZ9J
f82w8cgDvuikojM/5hVWHn5kKN9v0F4qwhpv/3bvr3ZpZejCG3oxv3jTiZEwIViH
lJX2QqR9Y5CCTijicS//7qorPD1PEEoX9QBGQgPSEZS8PeB4aPoMm3oI5MCOy9xx
U/4sTkqP7/ZaHVLSa+nBWn/b6D5RBfTmy8sv4bmwEBBOQ2VnRIKv6zFp6L+ym77Q
DqtRhqIHUwhut1tRrZB88AZkM+XAV2jYSNi1z8gDfF668vjmf6fRedNT3y1ACLB3
3hMKbrj1Nn3TGl6zfKt3CtmChwm+SOD9jNLGhDsS8JzdikpzK5oMIFlxsdZi1Di3
z+XTvY2JB+6PSBPklRb3AnC8OmlaKE0dr8Ax/7cXmowqEOEtow1ji8LuV04Opf+v
M0ooI77ttXljWUD7DQJOuSz7drDKhpOKtA91BUglbb7zDrZooEo5N/QxhL9t8yNv
DLp//vG/qh40P7fhbfF/mCJ82ACk3CusrUhcmlCCiglKmA40c2W0NiMfwuS170rK
Mg2a05VWn9HS3YYEZw94DzuRrxWKcLUkCAP6fGFTlKDRabp6nBC4dvz1r172hy4J
UKSDDTtW6Jj+to+yNfTbYf0GS7MoqAp6QXJ8MOjMqyaig26URgXsOuiacsNowiUV
itMz+cw//pwZFTKtMJSZUdWGsHdxNdx8yQEyTE0yBv/6W2/LMs1iX3k2XHi4Nx9G
xNfskb5bfchkad8cY8Bj8FXdElzVNB83/ztyKyW88/dFPsQ7JCRtDY4t4/9wPinV
uSrUECkL1shNNptf21a9DTfu6Cmb/i8wUoR0CcvojclOaRtPjtJpYoPzMSAbmT4x
NoDxnkJgI6d279hDJXKhxB+1TyseYCYsXq3AkHVx4XxksPUuNvgjSddNBPPRfMlp
HD+aWFgao/gex4ghMSiHREkV4k/dEHI9PeIGo5HrXiM2p1BLO0aakOHJSCTcZ4ZV
omHwZQjycJ5j7lJqb4lUBO5rWy6e1C3tPV/J2USvDpRaFy1VA7zyXocDfUF7zuDD
cT9ubGemwG4SsIyokpF+Q/nSJlaKYPYeIgvf+GNXgzbgwots04A0Q03qvjZaM2Eb
yVf6fjHVUhfEsL9im2mR5C/LKE04r3BylK38iMxkjtmHpgkG6mIXvz+Osc+r0Pvd
8Jowt1NZMmSdeLReQQ3C4xKFtMXMnAnbq9qRkilIHen/ZoeHkqDJR0kXI9xQDkxx
582/Q84+bqFoYbM9EfFOdRNSQUy7HD0c2HvP+4xywvZ95XleuyXaViirHDkkxcvg
s0Fhdr07nTBAacbvhN/Wn8Z3qc+gQgXRRt4lEyB+/wLKzydvlpgd+Sb2VLOoV56v
2weaf2oHP4QUcM3KhyboyPQ01PP0VG+WndVhm+pPzeIw370ndyaARcRmoKKEeYlt
eyGO4TUUKrkGwcwkT3IIf8HMEjKLUu0K+LM9lAnsgldWIIjzspd8XXYxYykLN/eF
Hr8zJvOTkXL4CXc7liF0mQkyyKWF4mIZ8KqV9OEfqDv2+fxniBSKPY/E93oe3XnJ
RnbF5SOZI0PB8+lJcvcePIpNbxCku4DrVhjmDIrQwd9VieDxxqYsc76KM34gFyii
ziIX1uaHhI+ArRW5uLLDSwBEQsst/31QD1pb7Giowv+CGOxaOthhBaGd7D+fUzwQ
uVUdRZQ4W79GueozVE1hlnjKpVbUQTinTI4oGCi0UvzH24HWHfBajUus9+aUakTU
ciP29wO1ql6bWlcR7U5yzwQoMZwsycPTOiAcfqab6RwjOjQAZmHo3sufpwXWJ0Tr
SltLA0Cq80wGIwElJsFuVpNPR0KNAIFQyKW0ECroyZXJQyGt5Hpa01gQxrAqeI3t
KSITqn2sB/KHFDugfztwRDDysK4YWqIYfmqhTfQmXCk0dzKKTpSrvzhiCJlw88Io
khjyG85KzRPkWX+yPGTVaZ/Bp/E8aWGO7GU8DhFmmRQm3q7B8zl39mBfjoMCG5Ld
pe7qvID2/rDqlkjktQRrNDt7pobRqVYkcL/fDyLs3Ekiy/+kLS6pwsYeZMdAJ0vD
CxY9NUJbFRLA0cGgmhrtToD/PLfywd4obCOKHFthka5fBAMhWwV0VUTrBv9xDgnR
s5SaO5IQm7EN6CH9fhq9it0IEi3wAiWLhPz43hEAX2u3y4v13iC9YkSBvVQuTNzf
rUCarBaxY1I4KQZszRndfMXtRGrEk5rTDCVyAQQ0klVxbjJMoIv3dP3fhsDPs9Ms
v1m+kWtMFjmntC97tEzbuhJ9LzcYv9RuI41FiBqz+l9WYw4DqegPQ2pG/axMnVv9
dSuHEo+bVGbzlCAuoQq1m5rgwnmQycpsTeHjv7jpWPIQbcN/l5Lfou8j9UFVvWen
ZLIk5yG4vtRivOJo9qnO8u5nfLTCqJ3P44wYlY6NbRq91BXA9u7OYMyzfL4iygyX
PhiNX1j3e3S8aUBx46sHRYZwFENK4SeeMig5sHUeHD5+35ypzDMv9KUa8BFq0CBx
aZ7QoG4AjC7gyzyk14gjVLHb6BMNMUw46UwewRwnC8XwpvYA9y5XLTEyKsqxilgF
Tu9/F0r+LT13Xu7ruYlreh68vYnaPWSuD49PTvmHCpHF7gMHBO1obV+DFLqzVB+g
3XC0tA12WBf0mdBIxzX3wWeO4xRfSI6GMFAlAak0en5VDBzGYGQVNFlwgzYBD2Ao
ZCOIrZjhp6hyCMHQjyqAsYy6OOHQNsZEcTBFnJY/9Q+bNTDG17SDvpUmllcx8oDx
+GnDhhMnUZwqnb6DC0NdQv02Se5N2sJte96vdabyF4IvxCr1dPFTyDNPaPjQNBRq
48GPXw8xtQany88466TIYDKm3jRv+3ZLRkt3X9id1hqkBdtycdRTWtdmBCk7S+4w
T2YiWlZbUFOHi46kqQmU94xFZGiVK1v1xbD5yp7pdS7cD3PH4yHB/jLOHszquv2M
A1Fb34FPxu1wahoKZO2qwSD6nCyX0eLHWRmnJo3nWBEu0O+RIFQsZRnTPu+GgvNN
TaIWOuCdmqXSYPcsdYPZPR+51w9xcGTOQf1+X2Mnwj3lGP/LCGGMtHJEZHqnRdOX
Nm+DLvnvi8RIteVldDckWAj4fLKC8E4PgvpqRCANDwAxhhj7/+NvGEmQLcuurZW0
9ipZYG9PTILufJGLunK2YBohUfG1MHE40iMNgCs9qzK8REVzID2SeVsZCjbMQ9gY
8FfNoJXb1AREYpShfuV1YsgufUoq1TkTZpX8VZrj+USJ9jnzAaV18/2sNI2iGgPf
D4etlMqsZ3/pyJsabxFtS+kjyj7Kk1hvOQk0nsNGsSOpAPkKOkh9P0KrWZwEGV76
gqxXa04U2G2i5prd9ObvAE7ngf0aUQvW+3tbSyss26UO54AryWDsG+gvevnZLszB
mAwuY7qpIhVhnR+Uh2X7wx33r2VcurjjLeDsJxziiKR0jY5bcCBaSy6E7X10i3yQ
FWVOY8uZgkf76LO0CHGOuDdF4jGukuERyzPKZ7Jy13Vdek6aDbA2sxoUR9Ba+Nym
7rOhkgLYzrUDIovwfPyns80Y/lhxOYaa/G3Z/fCBcG3AiQ3M5XVNuGS7P7J0KvGC
QUravS/gM5LPD1VhvyLTdRObrJAdzanLSB+sYGiyKSJcw/aYSjb94Uek095A1lMX
tFGV50c5YfjgGeaoqvimwb2HtR+K2zo8/h5+xgqWiHVg1yYrlF6yeBJJuqb0xprL
lr5rt8cruiwwZ/NfV8rWJeHEkcUlsOp7tt+Lt8QpUsBVIVxZiPCWyOSDtY1zah67
ibcEdf9Oj3rYxB63E2J9rE5p3UVsseVZ93xkk2ob0HoARuZGU8j0jcxPU0eSbOFX
Sn+dnRBE69Te/xwjaI0SaAMFmLigHxnKr9j83iNGz+ZU881oQTvEJClMPn9s+xi6
n8WeMpkbv+bhW5+ihRhtYRCwk5j3/CW5sgqHsCOuIHwN+AUe7DEwePPMKT8dA3E4
FRmHPfc3J6bQdVUtcnBGy8f1q2m0VZU8D9VpBhErSqZLCx48DDKo0x9eDV0JIHVr
ITtyFKJgbR3d0CVxv/DRHOdvHNNyaPWiKK3E5kO2IUmP5LwwhRLTtP092oNOoW9p
48FHaqh5xhnE8kvJIS+584BhlKxNXe0VtRzW7eRaA9yZPLVi0lyNoV8a/8WMtu0O
yzsHrU2UP5Htsw1LfU0RL/M5o0KlRjkSMAbannVI69CiGX+AX4EL7hIWVGcz95do
VQq6fusnmmQ8eUoCWSKmO01UieDs7FuF9/LAfPpF5pTOUr3QTDi61yjU7L4+kPdn
uGBkR+1ba+y+nNXhT5b9OZxj3bKq5nxVSIB3EPkdHjx17BbAgtICyJUEhBi+FSxH
IYrBV+m08+/RxNVTaxX67IaP2KLltw3tIdh7SPeOLCMbh1QEpRcFG/tnYDg0K8Jw
u3PTir0eSRugt7Cs0QyK7EiWvkIv/lKlXNdogzTflh2IEvMJq1G2KE/3qZaglMuY
WgkhQqA0UlzaB6VfR21v11DGJVfj1fGryaI+KPORxsYeFC3XNmvOPExOTTjG88fG
lp3mr1IR3bQEln0TZzpr7CwR8YNFrRFpNEtIKt0BkczJUoVlakMrsI3tXnwjAYvN
xppna5pM32zaCKxN+cDr6Groi1PwWUGfVr4r4nglSO+G578DFJfAfrgzuZ8flDai
mUekuntoA54Jw2dZ6fd1BskSnTZ5HRUTZXxlV/4vdCTJgvHbiWvDQ6/lsg/IQXOh
jAkloe6RTkjRobV8oXcj7uG2IOOVn/tGfI62+yUSoQKBDE+VblkBjNo3i/JOTF7d
VDy6C9mjx4sxc4AonqIe+ZlfKmHja+cmunlaBBzxT7Lv57+wlTLvBPc7Jdnp4v9O
MFqetBQOCx/iTCdUks1qn5E22WhBmYSPrMPU2h0q2R0sc2ziriYoXNsFzUwn4X3Q
hXpkE2oGEc3SzQkVlX938Iq6ZL/pd2tZbbtdb3+gGgVsxtXExyvdNUBbtfcoyS61
WDHbws/zHQ0kbcxgR1/DsQj8TloOmmtf7jtTMdlN03nSKFb1w/I31Tt8KIVcQN2B
lwNiD9xcDI87q+9JxQsUjLaT7ezBQxM4eKHHBSH7sxjmjxojVOJlKSu5hDBLDFsr
lJ0BzeurMAVjEtvzB9DA4ZctvBKxdV1ybdY63mPlwbkWGFvIKMAk7I1dBTexUL8h
j7aX4ci/gzSCVzuyft8nxx4NreBpWS2vJ35weLl+8YoeOr12G8/pFSID+JZqze4Q
r7SC2OkDYJj/icsvuAgMerUytrLjl0Mkm+EjNFLfcq8d3Px31W9Mp5nFfQcRfruX
CAuZqpj9V9VSfAsDJBGa54OMzGZr/OHiN17E1x7dLRgFmuYm+XthC444nS1WORbH
/H46Kpu+LGuPlVk5Hs1D9UwcYpBNXHZpGK2duRzfs08RfDnPWpfJiTcEgh73Agyr
Tdc5Wl066ZpuCvtVG+TUNForQJ2/nOAyg1pC4wUm+yhf9vi4zu1K/c+JIoFDbf9V
UzyjDdu6LsVJqTYRSSEpfpW+JaZAX2NFUo3d7l52XiWRqO03dlI2NHAaHWKhf/c1
KPw2I0SrWGmQBSyf/d0jWEfzzlDYT0ZQ50JzKA8/MnRMODgLto4iNpthLRQ0v20j
V/DQuLa3l/vhej8EoyDNPYatyyeawtxEVZyuNUifw2+lZ/yUiGe48AqdpDRG7iqA
8Jhy72a4tEeCNMqIm1pRPRAn1S+p+Rhj9Xl/93xN2InfmbMgdH4kh0RTgSW4pVTk
ji00uIBo5vPcuSLejhfvJwr+Nx9fn4Ew7J3m2cG1ZGnFXu3uzE6nypUe7tfwniYW
vYaMctrew3Bc5HxHfRpYJvx3ueNo79sp5c4aF3eFPVeeh0iafswGx8Tpbd8n7AB9
DOPbLCsRBEvcEOgCxVNy6Rbobov/9sWMto9nCSu0PYKrVeR3UX21b5c84Plgsn2N
AVKeGwyF5ywj2b24r6OpMVT5TVNiaSbFQbDY9T+rMe4RCleA0eXLZrQT4iKAc81i
d0i8aIcEfdJCCsrCya+IxGQ6azUV/+AhdCiL2y3N28pEwvpucCLtZn259jNGnRJR
yjc4qDG6sDxZIybMCbwr8HMHQFOnvKRXjy8OtAx1SGoGvjegsFMAGCBfKiVcvxGc
f6p1aY8IeNMUq7pa9dols1gcNPzW/68tl3dwpfxW0BT1NZyxxb+2Btc3qCYd3nFW
dPTGY//PKo6Zkjfjj8eNB2q4UBb6NeOHO+6iavK43xjYI2gY8gh6uXb9GihXzlB6
S+K6hWsisYmu99UDMj8tAaPYyD1kOfhNOWHJJGdOflhEcJjSUD1YcvvjeyB3im2y
WcTQECa67fV9qL8zfpESMGq3hiekWBX2tzNYEZX9BfIwmu51tZYQ4kyv95K5z932
Ys26rYDpTECQDqYmFJ6m2NNr4UxsToODMvC7WMvzPCWUL2gOjLi8XA5iWK+Hl5sO
XoP4rekTX0TVKK5TH/zIPcFKpL+hOodTtLDVqSYpxCsZwNhSb19GUPC6WwmsFj5J
GGFYI6Vuyzo3do2GxumHvBpZ9v4BilqUZe3Fhy9MjByv1tPh9+hBCUiM6CWJRGya
6KzuzROn3odt96147LWdlR8fn6x8WVIhs/g3ZCDziKDUsi5lrjqcqZTgPD2LSEOA
XS930d+gWP0MKGTYy29weH6h7stGak6Ik9LjP2IqDn9aZKssY9D8db8FsOp/L0Kn
GDM+yXZFTHQkX22pWXTYGqa8mhmYX1xW7LGcpPmsd/PZziGoYuk4A3HuaVXJ66ie
c4A4fQMySMb9MZDb/IGytxODs3rq3Ebq8zVuaxYA+4XjKA/T+EB7sjQTX4LWP4wN
fDEjdxAnkUbj/qvEzUddpsV04j5pvZkuxAgyLaUPZqsBHRl7mwpFnP7Ml0gqKDTP
P09nqyfzM0wfov9DKxa4F1cg9PQQl62YY2qOVYJNiyPB8ayXjLDPrHbzQacOlb7N
HFpRrJA557XTSR7SjsuapjvzZ4HV7mLjsn9JUxlSrNPHdzutMviHvNEfyqO5wAxo
/8y4XdBGoPYhg/neA/3DnimizBAAJdpub27zY25QebwCcmZYDAcBb2dJwNOUEKW8
N48gFh6c+6t3YXht7wJtoUv0vzhg3d7usT06i3p+JDbh+0JNlzFp7l0vREM3liRR
DZkZl8sqcNV5xRu5p14cNLVLUnMfA5NyF/UaXRnn92JW6+Frf+dJMqX1gmCLpMP+
YkWn/cScwGSwt9plxzoM/XmyJ4AxD8UdyMAh/Y7uqMqG9I4DhxA+EbcL+tQnhaaZ
Ea9XNY9s1CLPwRhyDSOKJsWWTvwkMf6KUqaEHJJsiVctG0wiNta5wlt3IwZsOi9l
Ve28xeTVcQhKu9MXf3WYCPy5uqSZ53qek0qh4ZI2qFOcCULiSduX7GaBZGgXfXDz
RPqzpkKgqWwiDSzekB+5IWx8yEFoZzbMiSRKxUuCcXbHYgH88Gm5xwrWoU3Q6iUK
Le5zwCWKbrvKx3WUWb9TkzR89yckU9Z6oRSHRkJHoA4=
//pragma protect end_data_block
//pragma protect digest_block
4Y72X9pR2cPFdUiijXtHetEwaEs=
//pragma protect end_digest_block
//pragma protect end_protected
