// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eBfVKXDUIBLOvM0KNYVR/RpBqJUvzajOoGhW1nZuKgLeYoDyHeP87iL/mdi5
dJuk/bDtTA0peeDsUMIs2NseR4PRItQ22RayeHab8taCpVGJYTvtBS8CA+se
KSwxYZZlp9MwskJ6mp3+F9oFhUwxXWBggDmPdak2XmLEjPBDA2XS1yqBkErU
0/MI+Cj+yS7DGs/MoixW8nk7m42l/CNmWZgbyqmFe1w02QX6/WkZSARbKth8
XnCbVHR4PIzKXh4ZXpxjGi0T2P1hZ1dSJrxqfc+Jr/8/XidRO/8oxiEftRn+
DCM708RU4Hw4Y3vc8ECiY02TzF2Gm5+njUWfYnAexQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mRxfUrpvdVuWYBpmYjtZKbNGHlliHFTdnnsSWSd7hNCUVPsP6AED8qQ7r6C3
BUWJHavmERb0ALtBbtvpfy57FNv/LUEV9NXK2SK6XMOKE+VsTxuKZ0pmMO4X
vVl7Ia6VVWzT8VGlRMGejcl921hGffbZLxq5okSs3HetUyjVCJiNqHILHdWK
FsVRFS8KfBq5RL4xM7WtLXfI/I6AncDoXeHVueq+HXPd6dHbtaiyfD58VARe
C/f23noPEyAL5GWG/3waD7BpgpSNQ4bmRhoxiQegiAckB4H2870dOmsc4eGl
kKmtGH19bN4Hhs/hfD7LWy0Xv7IEqiZUoOWb50Cyqw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O06wR1fQl2VH1v/HxnWYdJ2NoBWS0U0xMYWmcoOqDncLIF4FUqbkZ4Y2RToB
4PA5GmDwuXFdwAuQqFERQLbzQNRjUiC10vFo5fjD7L+Q2O9w/NlpCelWZVAm
R+Jmw6E1juuhlcOWNQDJ9SqgIxBc8N/GMjWk2pZyOiipXgF1ogQmx4SdiC0z
c35Q0JLE+HRIb7vwLpKQPl2bp0qOZ8qyjSE6TX4q7BIHVc6Umu6lUbphJOJ6
hkvDwtHMLdAZWYU5Mzk75wiRFXB2cJgLLUubNpxLQay4OIa+lQY3IVjvWKUs
4fIAu3GyTeY1YHBY7XogehhWSRxRhzo/AAE3C/3aiQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QZXjdUifD/l9BtHGaFnBt9qZvxALU95udaXHnZSfF+431fNSSkdfLt1dmTv6
q0id7r2o2i0C1066ULeNoLWamMFGimxI71JAKA7PHYS6ot8Mnbq1q5Z6Txzs
wVWHTh1RrWpo/5nh5IkerP9SCsTZEy7W+L5XuO69EaChh4HKMKY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PFby5FO+X/t4OWQ41p4eNbfZOgSeCzl5FVKjRdpQvCuN1jRotzHUjc1Otfmx
wZsU2S5bFKb3ZniggbsyrVJA5D3paPrE3NQI7+PjmMypUAvaRPGguefAltNT
4RLSnDM0Sfr6mF16y9+KSnMUYZHwEN+nJy0p4J84MfP/tXE4l4lqcToREYjz
vmG2w0oPzqJtEDcRdpqkl2ZH3l2cJ5nC+FyxhO9S7egXju1A6Zt3zFIooZz0
LhKwMEofGTNWH53jwlzFik97mNaYsLjXXkTINm3pRpRgh8jO14EnIZHvCV9t
sSH0eMzqj8CALnrh6yrPYP+eFgI4LWW1ptdLzye6My8CJh2Bg06lIU7SxKW1
z/fwrKsVuaNuelw2wYJanLJd9SeWkthF7OGSmlVoNCGB2bOA7ua7ieJF07Bp
7lWuB0IzqML+WusDo9SGQoQ782FRnF2djgb0KFKkcSnasXK89BejpLIHes0A
5LDqKyugZCgON8pAgeMrGCvnPKTArooH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cvZtiSnY3TKn4Oooetci8jOOMBgpZ8UphpZ23bF66tGpCYY3EC7m0m6ws3Fl
L3d2pgiXvO4atXn9hivgYpE0yfSCyjSZmaeOOTkmbQ6pHkkl9f/Rt5cZSDgF
2GzRMy3+Gokq5XuW+8mBaiYfEpD4LB5tTNz7tJRXFjR9LGmKMaE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p1UdMSo8cpoGVC3QzcDj4rn3M88uSEx08Q809XR6qQYgd+WUrU+dCLFNxqM2
FYob8hqbxwOJV563O8r+tWk7gIBZaq79oZ1xswCpf7TSqRB/bdsd1rBuhg6+
7kmWqwOEjvZ5up8CcpdJucWX1aPjOucB5Xz29sfml9roRrtrIUA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10784)
`pragma protect data_block
U7DYyjrP9PbaWXcXf3qqj1GY88x3RW0YhudGTFjISArj2JQEdHxYEjfega76
QyuLn+TIJE1642GRIyFl8azIZpxZKLzRTCT6Ztr3XxYruFp9OSK3AKz/3w+L
SXWruqYZhnphiIruhG6/ygOHXAIseQIQU5kapu2Tc8rEVtO/ojq03yy2dbK9
n9pdMXhv6ow2t8Gwa38vog+QQdc8NvdZFvES5Jo/dYCWte6S7scTsIf9PJ9c
+yW0/yOZODgb2qd1zhTWls9O+TLtWBQWW+X3akiu1+TJ20ykozEYIfQN1UeN
vNyBtmM/aEy+ga+zHnzzafMHioO9VvkT4yidov3gtzFxaaj5VbLwYtif+vx9
O5PXbbzV9kVhs6yXBhN0QkOH/U+YY2flZRa3EYVNm9kKLFqLO2xLGBKElKzL
RQEteyuD01+p30gsT+ovBqqnoXKCpDwyLax0VSYQapJwDzVnl0VXAgxbviZ2
Sg0OHXf7VtIvl06I+rfKf8SWPaYwrt5vBQcWSQfPaK2h0SZZSgDwWolwRE+e
XRxcHOsUMDQwfugEplQUkQZ10s1j1G1IqhjBo8FQmRIh/J7uf5yQJ6aI7vV/
vsqTvq1TeFIfQm7wPuWfFd62yRCD8ReOBk0xkoSIsruRoQlxplPqPVgtlREX
kE+GMuxTnGoxmFIpoavWwz3x7AFavuipYcp3FKUhT33p7b4vvu727j5JT+8Q
7N54ndvpuMkp44p4IToXo+kvbIeb8s00T5AK/SLKYvDBE50rZLyfp2DsNr90
zE8nfgJsuaR6VCqpsj3HxevZbaLYCUugOb3texoFqFzpCoWu1fGDBLM2ICRw
uLjpg/HWvDPsMkW3psCzdQsQ1uuNoXlNt8fvCFjrAsEfGoNBTEMjuKipMZ6w
e3CvUaYhrtKJ7Ie6b3wX0k6N0xextYnpJeqHYPvDPvux4bbR4uVUgZ8bPWWo
bdCSnVHBeYrf7+MRhSQTJunegMq7wnV2rSxhbcaV+Q4PdWeyEwF8QBZZoYOP
inYeld98zB3YnzkG3fiPh3dQARTve/DFeSJV8BunJiXfJPLm7S3l0D6PaTPz
cKial0m8+G4xv9fBQB6DKcv+dOEAwKHCYpD7WjftpqBzpeh8XBlWQQJNYnCS
PWFrAAfbXaQ8QmEy4FQ1rIBAc4BFtN5fgHHl3JFt8ij2P6iztA5WoC5UvB5+
jEXD9smepECVhJ5DbM2bVEUVqYckxOtpOse7WtSd9bGJ3e/6Pg9js2VZSXWQ
sE3yVkap+XpAvBV07HhhFqDTqbL/fCVdEpKx3yWxdpO736NySBUpr19urCx9
kDgLtHneQ5SChRoQ00f1C5idEr4BOT6kgz1zr/oOFeyJBcg/PagDsWal6nDk
JDsu4LQ9BA/ctaRHRdMCE3ZBYafPOijxsi3t35fjLqtmtI5sLJHbn8Eca3DB
yoouiKTRF3kokBSjRzk8zVxCoVeeLgOMYkj4r2qVzosjhfPvaTzdgk4lv0aw
90Sm42CKv7RfV8dDL2QsL0UmQQEhel1qN9OS8bPWs98bxNvlXc0O9MTrSusP
ieiNCUl0A9L5DVt6ssolHFTCA1xCyRqwCIpKzsIJzoNVru87aCl4BZuSYaWy
6h4EVQyWIKjkxB310tNRG9qXfedA804s32RIeqGDZ6c/2jRfPx7mpArsoM3I
TWeU1XCGYBAR9W9IXmsVWEMAkhvX2i54GSnBb/Nq9E/KKB5jbG88L0eYXsxe
wRLcNRWmThcHg/9p5BbNmpGSiCabyhcoZgVkQBi8iws5SHcqaAkLJ7LXI5Lo
A5ZhHWxqpNQofqge2WHT2P6gXK3UnbIZGznZ23dGjoBmy/1XgrgjZKxRUdkJ
5TvRmqEIUX83qdEnWTLriPP10uVlRzAoFzU1tvYGfaNKDhhl3cAQ8g/pNLBC
VD96d7D21KeDVE203SOjUw402z2PtrlOzTkHsGlLcMRIECSHlWlhXhIPo3v+
g7XpK+vggAzJwr69OPV3b26+ALFopvxQAzv75M8p06MOa3/hmflOwxnn71H8
maJclJ03huQAjsz7iFFflFLpyNvVm+GwE4SjG7Ks5ptozFJx9JMJi2IdMd90
nOOZ7XaY5gFc35ACNW0wwAXpIl3HFLJWZZxRTaLCzNxlpu/V+clKet8vcOa6
MRad179YRxWZxVR0DIH5aS7hnRFXhfBkopuBrZKThBx8USnuv3AHrExkOd13
QxoUkDo0diu1Gz74ct8ERS97HiErLV1VPKanF850cw0R+u1LjwMyZbQLCT74
Lj/cKPB4R2gI3Xqrd6nggOcIfGdC/RAZR+lhRNYBCh8/ZijyIL1a5rBmdQpc
RPDvTIxsbss7UpkuC8JEUSslQlZh0Biwzm7hFcD2X4kRBGac7rKwOGrJR7S4
cZlIoZcj9YBgKyXGiEPh0aZhwcl3kHq+GnA6qpjh8spUYnEHFuesRGANpFR5
UUsqWg9+G5oJiuIUM5jtBMtzaq5BaWnYOgoiUouNQjgtpawdBBpYXqL6RWDU
dmo7rRBhXotYy/NnWU+40ibGav15ERRdXF9WxfepnV9zmDd/RcHu8Xw8i4Q5
d7BzBmosCZQqdnFol5RItsU8A7AaNaJ/4Z306e84eR4PTdnBu9PiDJLEvE2y
yt6z06o0lfllu7zmNK0Gm/DF2a76kfyE+dENhj5Ocmb3qoJlAiCUyWUfg8ko
eQFx8N+udsKcNOEZ6eq1kJv8lAHZsNztA72SVU/JbCFEnZvPkSlSbs/AZOeH
aNx0a/m7Vn4A/a9Uj2fOz0p1cEDMuaRO17eJ4TJ/zlYzEEJgLk5OUJxEH3NY
/F5enRumXaAobErUGeTHI0pg3MWWq5fpQWGrgWDY52sIYCNHjBunZ/uV5CMk
gzLKtpz8CVK2rb9u1fAF/ULtaRd8g2rPJ87oW9wB7RqMyJm+f0kip6xNzDhf
tsWCToYG9i3p1ZqujN9YhY7MVunOqX8g0o805z19/qdNxjdlwfT6yMcGb0Zh
pbjbPSQ1pEhNHWqCZ4he3fRssdyw3THY3yNCAE7YNuDcg6ezQXvlE55XRBVi
1oJFltpUz3sKHzlXPqRzgGsHl4Ec3UZxxg4DsJHqcm1s7Cg/FPeIkqR2lqR0
5ZIkHjQ1WT/z0pGloqAvLw+CK24j3kunVsgXiyyfxvAk9MyBJzBIQT+a8ohN
OvDjTU9Qu0iAhXyTg1zQXuwaL2LQLI0m3p0WsYxZ6EcK3C+oT+0ok294yxp6
W1+lPsMuxzIsyxGz9/eHXWMyMWgpGCa+Qs83NG0yQynv2CmlNsFAC439GGyg
wNjeeIpBgUSoGm8/epK4ZqrXamOUfGRYJR4VUVjmG40/96WHIj0AJ8vZES/g
Hk7bdKqOmDmUkAG1BGqjcADYZrqqXlonzkCo/fUg4OjtKdCmM4gRBC5iRpSO
uJ1Eb0GfGA5zW8W5fE2GeSNCIraRKQt3C5vWO2484Uoy2FNee+gRIx/jqk5w
1tidz35AIRz5xv0XpZlRY91iSW/Z5s58IHBIXMTrH2pI+6HhcXMTF8Tkaphx
X+UDnipCP4NdKY/3tRkGDAObIEDMaPMSerrnU7aVw6her3ZUu9s8mt/u5MXU
3y121xiGAVo0p/zaH8UmERvItqIs3zOm96ljt7OvJh0Ci2+ZP5dkoeFr3Vzi
4aq7vOGz/4QSAoMmffaJIttkpsatJnceI9gbCLWbx02HhP/zbhz3ZDBwO6rq
LblsVp/JCvDy+OlrItUIwQkbJE7VPYQmM5ukKJItkZ23vEEj8XoH9cIh7t0n
Ljmly4HRy8LldenONU2NSA5YgAmFeBpLtrqUO45iXRHOoypgykLZRFcCBQEV
wG5KBAKNOTnq4P/JNQTF8VxE0ITR9RaBwv4xWeQZV8xtXM/6P9f0Li4NysMD
VqIDiod0cCSwTWGtlc6Gz//0fG+gfbS4LZCdqLoeMrJvoHEzyJIZ/G6Tepw+
0xXeNTLWh05iVNC6nW3DFj232/j8esh3qN9/v8WUMJMt4HvY2pPIWSHoL8km
5sCykudZ9pBd3mFCnskZYMPxZ0dxPb5AK9m0WEEKYxA7WGUNTZ2j1ZR752Uo
cuwKtKDBF6Z8Hgau6TSS7LCr6hq5zx9gMvcnIuMEooacoUSwone7mmsGU4rB
qzO6knGhXadJQKOgrD5wVfkYEuyQthJ+m/pC3aP+v2h9YJzufHHspSE55bU6
AqxufVc6YsQXid9smx5bkFICp0eRVyir1B4RP45l3a+vh/Rl9mXlUMJiFlOj
vIxaIjP32s3zUwUah6Y2Tb4k+casFluXOgUnHLz67DIPGEkyWr4Qz+l77w1G
Uq0q+BYKRAFJf4HYqvRuq6COSv6Egi/qvqwUCrVbRvJuNBg6xso+M1XYLcEk
17VCtpiSsjjESJaC6kJrq4WXbwOh672fAJwJirDqcKYXG0+84Iita45cO3hF
TYiW7WVQa3SQsjJeS/HFhmn7jfJ6dlmWSUchtSSXMXbu7u/W2CnuAe29SUl7
3MosyoD7ObEomF+pEv3e4voGRr8GLCvCHGIGdkQLxd42YLDXF57EMXTnmxtC
VWhvEavYI/97cQ7/ZgqvFRDZm7GQTWduYQoFJkoopW8nDRRdtZZ4YwoQgTgt
t6AxnpL+gqZXNtiR4sYBhvVUuDT6ArYFapSJahg79rq9M+zdwt5cMwsR+vwE
NCs34fyc4D8y26/W3wcGyxydO+o/AgyxVQngY1pyxklwn80qyyv/4KQrN1hT
n4LZFgZdS1t9CrWobkXFw0IMOmniiNYo/Q46ZFeNw6s4cDepGX3oixAhdotp
L4/emT974sucKz+QNylVExRmdmKRIdxy9YibiiIiP36+NB9lKt0L6wx0+fC4
DzUUO4dbjNPuFI9V9guHFYkS98sJFd94VpcO/jY7RdF7M63xRO3rrrlTUot6
tXcUPIJMOkoPKp8n/CnZ1E5OUJXU8/fZvKuIi/w33s8vQg7qe7tLweZKkLWJ
I8htDWrvaISwjBa62VrvO7hJN9jHYd+/wUbcuoeMdIZqhvul34w5F4WfsHjQ
Pt8hEZ8Le/XWlLHljgYJvhacLN6/bdFjPzpR0CkrDGeYQRQ+kp7SbmZJdcVx
bfF/Grp+wlFribQtngv5GKYAdFwU4Fg6ut1v4+PTKrqAJs7sn/0pkq9MSJnU
t1RC4giAxBRwYtA3/VLOork7VQR2gNjgnjEb9giZGN834CM59kxQMs2cKVXD
6acD3qp3AVhvH3SiTRxvQuVU67Omaput4wiZhKCFPBnx6U7f+UMONSZyuflG
ARAjKCvTFUsP2ZjeRqMB+1+dUDlx084ubOVjpeU2fsW3gC/m6iPeGBa4sSQs
387GdliVL6mxwfhmbImVM3KdPkQITwO9SbVzEUUIqgsOhx1YwV9vxYqX/BX8
/8NkeVUkqB/JWmNmYVqdgdIi79/F33woTKoUVfXwEk6ffKeJ34d57cdd6/Yv
eif560SXYySSwasR+erxAwO+HQlqzz2AQJ2MbI2yAnzmuVoA7JuK8+9Vb6TS
gVt0BV1NJH/U4Lzk1gDP1Zs1ZHc0iF0ABh+5csQ2PTZoHEz3EHzIkjiO4Rhw
/fTSPGsEYbiH9+HE3Sl60+TjMygKe9EPPGXs/nk+OMd8ZlhsFUCzk03dkzei
t5IDoEa8HUtbbLApj0FYzjUZpCpJqLShP6LvT/PO3UW07gVwgCQeTFu74VoH
RHZkXUgnfHYt76WW37aA3bG6pCiV2qBZowP25/SMSOGpLXLxlW3SQ59H1EF7
YtxjIACpj0GXDk9o08Lq/yBuUfLmS+4tJzTatBywRU0yI2ouhDUaPOo5mZl5
/wMnnhj2Kg4Y5x25S1NRUOjdxsp3v8KKOyVkrM/dz1DsMHReMwklj9AJ1H6v
by/EGShjnoxOf/vVEz7Yi8Y1OOcakcVaKQ8Y/zEJdA0urlNmyc82umZj/404
dxt+jK8A5WZCrA7dAcyAj/tDYS/SeShGrb9lEuYFZqpRhNZP4xbkIpWPruIw
RbXMeiEpbHKJDnnYaAw5TNq1n92jF18bse/mWi4NrxC4DGqST1NrEj5wj1zC
fjWytNPV4MDA+t9MsRsuK/3ZnTMyV8nuo3pM/AnHjTzUw+/ZM6jwse3342I0
Y+s4ofpEE7VQrP/FmCD46LxLsdNhGteIwRPNB3ykWy8ZzOTi1P5K9AfZqPYB
hY3gn4tD9BQU62ltO4Cl2PGUct7Br14nTELcqgsMSOuW27Decpy/ihhaJ9UJ
/9WrQNf62GqfAeBpj6fqI+LnZsKYry4BR6DLNZ2BYvFimqgXYAeVEYVUA4DW
+zQalR4x9Gpa+hoL6qjQzRunX5smlAZARBJGueZvow6oSX4aoYo+UoIKrF4R
29NjzEhq3qWEtVdX8NUexeGKVul8SZMWMythXB6QNB/LMoITGxAZ6bROsDyj
xumyNR92wnu1Xd1qUXUA4cSr2qe0MkgVdhRtFxDlOddzLlox/tasJXPaOsNi
CQbz4vPmUUzFuDmOEY54yybB5iUNtG80aJFN6EeK1Q/77ChJHVyeNjbZ/+zN
HIpf0phc2qu2bL7WjtnHnDx+vgPv7eowg+7/dP5sT7CDPCCZsU9uBf0kpzNO
+lxYEwutmJ+Q6aPCZn91JVmlfnaIU+kiQcWuZif5tCXShk9uJX402fC/7v7X
WShGVHHTx93vmm6I/jNt6LayMZtbiv6tNLFKTx/RadTZFp+2bKY/YbLIq4Te
6aVxcSWglqjp7jIK54lBFDkqUQadsMasF6u2ceTiNVsyixXdzecG7W5HbRl1
6V3AdGvEFjy9O54dSekqIcCCzsOKsHokU0fCaX3EdBaSmf36F4VmsM3joQPV
CHhyPmqFOXI4wlO8xaKMWKJYJXOa6knzlw87vgM4eDEeT+bIK07D3ba9cHI8
OiJhBoFWzHFfl8zmvL8Q/T2WVFyl9Vd5x6R0VTj3eHJW5ahy2D2sdYP2PD9q
3Ag5MeLzcR1A2pcG7KiHGJeFHD5pOB/glJt7e1PEBNO7Sia0QMeMRH9YNdJp
/VGTnfeRPvsDBb8AW8uerCopjgmd89NxAs+dd1Lu58dEWfCSfeEqtUZeZ+rY
066h5FpQ/jEzrFOb9HedFqZHmHCnZ47LfViVaV6vsTRMZzzDke9hImEUpEjC
KpvBnWATX8tH4nLj/4Wp8qqBqRtmOuAIUikRIytsROdHx97TzodSM5G9LL4q
Dq/BcIbINUevDhYHY3j4CZu7CjW6D+3CYjlHEUxGamIqOcYBSU93fCN1hWA3
8bu20PFDLdmJgxXEK4zIA3STN7fjGmmHpzO+sh4PvAo/pBfrIX7nJL/4a3DM
1I1dxfTBBEdC5tlkv2jg5+qbSkzyaHmkUehMl7m2QVSS0/LqRM6Lo51Cjbkv
TAFDqAxmRy+swMKCoaAMJigtN9OPr1/k1jj6coFYU05F5Rg5YC51AWZnGfJ4
/Q8qOyMuK4wAsDETbflFtLijbvhFjSpvz6Yz6Ra9RWvV4ubLUw+kkraC5fDr
dDSBr95tTawtkH/8mS1aoHoo2tBgYfQ93ABwd+z1n4bFsxqZZORiVfrNGBur
4+2tcQ0dpau50tAIsV+Mf1i0C5b9CAdsdfxLhMWAuJkd6ESYS38CTKw5J/kf
XJ2N6ysVvzOuxucrbWgaEblGBPclwdTUUmoZwWDo+tPbHD4aaxDbfodUKx1/
1R2ZI9jm04v6+oBgVK2KjzOARTcpWGwfUjgP5Qpe6HGz5+cBry7/FN4wYOVo
bKIwYVFTiQYrCAk+oftZW+rlb05YdYCIsHnGvQhcZs/XJGDB59y5Q5mgC40m
cK7cJK+PDYtxbtx8TeAYyQayONiMy+07WVY8vlSLX+MDwERd3TfpRrkLglyV
W3oBC8hAfMuCdbbYufgKJU0VE4TTz4XPmokdskayu2DvutAJdIBZUMwied9t
dNiznqrNUKenvC7CiHqjaHRzj33oWqpjCfB016K93lFsROpKmzv3PvUbPtn+
1qCov95bvEvLkFzqO4yXqy2qHxGKu9KNlPaK1ob2+pWFSQShLHV5U6WB7HHF
7s9lyLbj3ufbyzN+pjOuSr7aSReaae232LSzBaURbfYK02aUiIEF1Df4Uh+d
CUFh0cj2esejoFPQHGyLM0BwO6NRcJuaKlIj0kOUO4sV11duuVlw/A2VFh1r
SnumV1rXNgaaB4vrBIoEfK7Ag9klqXt7pTj572Ex5zbPHPSvLnfRbzfeHl0t
B4YyECvbzIxOwD5dy0lZhNGa5k6wszpq7uydIKxakqIlj+Q3+GRdykedIQnk
1MkhMR1mdzFtiz5NGIgu3yrh/rj9kcMHGuOXWiJnv+p41wtnXHySNeRZwabC
VpPLdYkzcKMZ/J8ZG5Sxr29DsjxHRUUMIgCAr6CSCxxEEXrMsEUib9YtaSDH
0YP557HMmFkBUwoN6evj4GneNDEFcwrC4lbH8tursMkvkKLTBwZh/ODQ0URr
GxtGxWipmhdfxzZeFQ2IxUEuQIf8typ1r23ES5tHtSwXQCjBmbMGc+hC70t2
szf24P5LHTL6BkbnZhLxcc9fjD+6ofKNmtjBLke8pV0XwRXwhgk9lI+v06F7
XbYwYuaKA9ahHqnvKb6XYtKqhktkylv99uOYW6Ny3ZumhnfuHmgmOiGuglpi
yYvFxiHia23EmH2CQXEasmvJR6kPtqDj1Nl0Lqmxlt16mEncq4oZV36MjRaC
vDBqRDCOq2OLBhv2sesQl3m4XzvMuxozwnK5Yp5QIOnz3T8ZK1lusIoG+mma
a/wQTdaccrjQ3nbhwHwyTwXt3/aQKjLokGbz4mLBJHMqECFZGa/h/TI0AdkJ
KhkP8rqY+ErEUqGOAbE3rPdySRVX2lggP4A5BzGxJccqAMROe4LagoEpoPme
rhW++Y1oyV99vDe96LCNP3ZkTJXVx2g5RJJkHJzWIHWMu8JYFh4qBo34cUpt
Gth/Zt5IeyQZIECPEJlv8CGxPevfO46w4IozFTJEEjTZ/JGdoOS82eHkNsWZ
pR7PsoWLrgoGFgXNqMuZOGopEj/hjAnDg6gOBwWlAFHN1k2SjrcwfLhuSQzi
s+EuoGQLrrYdFAX8JYFkFuoEUFCUgrA5RgR271R5lk7YjXn1oHYZ87159ElT
5cMWy5LZsdHzgWTo+65WhA8WetSaHQy6QOUDFnt1DvMVvdXUxJnhG4zoRwPP
JKHGFDrF3PFlUYJ2SSBQSOJHpibXR1awLBr+u+psAMUc0MYMGdmDQN6IHJ7P
TWFeN+8+vSFP03z8yR2bRIF30m1dcX3HLMLMVi8giLo3hntF1+3Xu/H4jkp0
Q1beBMBw2+P6lrL3jd++AwAkYRCounMMPFsA+au8BBofjbZxJ5k6I5NTYLNU
sjOGLbn8+GCFcapYTnpjKJwV3r14LYkj7g8ZiKBWNm02PMg93RxDTflg7ycS
DCbnSaEF9S7OEzI4tu0Z5VGHmzuLALgMGseSodXpOvhus3wYtCR9TAQ5mDCr
2eXOJHuB9p0ZfBd0vNv+wwY82DOImc6WJQdqHBEJvr6Yqaq9fGRkM/yL+VvQ
OsBk/up/j452+rWs0zNrhDKizbz0wCbtBnNTNroCf47dPfX/ppDJONic+5vO
pKxnjN8F+v1E/g9RHpfD3u+rTiYxA440/WuLgWNtULYE8pwTqLAbpGo5TEgK
SbMjYX8rMAj2DAgZtYRcZcZMGGe5+lOqF4V85ARqHvtbCr7urFLkmsGLMQf8
OGMjIjz2MYYUUk9xgIDyexiXM4enZh9DSDQvG/oXqFecJE4P7obMwHHj0dbo
ZJCDl2AmnGJcz601TrDhvR9dTkthbZdO+MEn4Dhxhgf3bvyGYUKf9SnBYRXL
Q08tc1ilyPe1SqDzpDXv3ai+xUFRGCBO98tRxuWTSGXg2paLQhV4VPs8tRhs
snFCAY/mT7wLUIoNs6PKnDV+8Cey9q8Jl/RRLk9JYbcvLXyTF/ioo8fYkH4b
V6aOsEjNNu/+NWi98XC4sMOrsrmWaGqQ+g9SCKhNvGI60Kx3spHs6NRvljQO
qqklZrOz/RnI16XWbKD+pGoas1RJP2YAfoB0tULh3xNxDCazmvmC2cXttgN7
q9o+zo1gVA64dLi31A9M5vmo8s8UmNZRxvicp2h4FfxrcBKEb8HznZgf6xwE
UH/iVMzQXp5hLvzqgMTUW5sdASA+htE1usyFUbpeXGEMuJhcX1jvgNBkOEYY
mzwMGFkUReEoRr828RmKIN7223737H11plsZaS5ee7GitxiqOShlhglVrRUA
NYRiVjAO/oGbjH4n6l1qyT3XuaO1aznBIVy+cEWe+qs+aRzF0vSwA1NPHMAl
g8q9doZ4qnuIP1GNs5oQmbOwj+lXXWS2aS4oeyZH2cWTm+iF7l6X3F02NDl7
XRvaIVYphdEKlXTUHOj6rvmFV8kxpI4IV6x6a5cqS5GXlGQaFoefZZUqHvkS
yfN5iMDHonhIJHAFGAJ5+qTlqqS6MLm+oHH4nHr/11YxPYhvGwXs63rN9wbJ
V3b9uypFAX5iIQzTT3VCvris451y0LdRNPH0ueeyv26h8R9bM2j02YE3CfZI
oH+7k4RWfAPPbsgdSb7GI3E7jOPk3llt5t5JqCW6XRt0h//Z5hQmkXETTweB
jfnUEG65SWsoCB6xdhMpXwzweuzb0oOlUpWjxXeaZAHjBOVEWWgvMhlaxzOt
AZqBZkTJin02zabhjJAp4PwBhfkxZLQwoiq7PPJ3n/QLXk/TlG7nbYKW+jYE
3qIt/a0awMuegpyXiUPdikpt+ad22DZx6VWBqVMPki/VlUvMyeSKyjW22ndH
NSvy4XDZjPNe0l1sp6KirQ9GkBKFxLzYpemTH46YLYaczJBhQ3XOW5cA30Ni
tgvXatrjCXy1cBxDnYzjQOxliNMkFoSHAb4vesrz4O0gToStv9G9spBP8WlL
j6yGqU1eiwIR0B+OYjI+1a4BdZgpU+Yx9O9OTNoTgjsWfS2CSBSodqspuvLg
N+YZ9Tkmk36jc/BlKfQgN2JEjwx/8Mn8uHvm/FijZ82vt9ZfBl/OP6Ob+lcF
ame8cWPVifwTcGDPsvXLYwUhz14KhBUufF3wXoCUSIHN9I0wTJCDHqUtMDHA
Y6SHEaFOW7E22RQX5ekeGJr36qejp9pQL+W0Y0A3cWEMByLclBEUr+wvZ1lN
qWUPDHKsYyUa6okLEvsa/5td9RYOHlxaQF+hitjMwhke9WDs8K8M2OBhisYV
xcm59PPyjAcqmJfcxZI3Z4woxZ6kifcoec17DQdUa+io29/ZyzW92UGemDI4
aajW+zQk6sx2GPP2iHKVAmWhKSa+3RY/UZbEju3lzJZDKSi4f9EacbxzJmjx
ErrEgazmC2GhrIhOdmVEzoos+FaXwJpJy9SOZdAanytmSQKOybzZiXg6WBAG
dPWsFg9+7hRjqbPXlIJ5pjjec6DV+URx0LmHOaf+WJEt3BXNxe7vLlXnUTNj
9k25QU+E2EQDyK/SsahZL8BGlT4b9PUfUC7YmchlC1ld9D4NwdvfvWU8AGhS
l+JnhPSuvNsgsTi+i1hpvBbFQ2mLxaipE+VS85ASohmLtaFzEL2gqN0kJvrp
cF9sBy9i4Qzx76SfSSWEv0zJBx7Nq1aCDrLis679DvPdH2egPvP865pl+aw8
3E7jwrjhVKAI65RzYSrVD9FgK4mFuIXLRNb6Zsr4Qn74/cX59GjK0drcLSxc
aXfSijKj+IbIriADwLqqaFllESECDN8Qt409paCeEdKUi0NPIgddLCjF70vy
G6uTCRF1HnuNjbINk/sxcUP/SbutOo+a6sHflCKDfjJQskWp1fen6g2zzdGc
J+zuiHSteOdfUbDN38DNYF3KpJVgTRvt1E4CTSnNi94QLfPM4RuiN0i5+DYd
IBQqMTvKGw3oD+C3i8WKJ5aEK/DQR/XIEdXVkv15EUg4dKQV08b0n3K7C7Im
Yji68CwzmXN+JPwpO7guRojZ5kzcJIzL8JMQoH/G4bBxNJJy+sJVktHNZArY
YLK/V2NLg34nqEas9awTVFXdkg2KjlycijEvB+GH4afTLJsaQFOM2kkSDGN1
JgbQqksRNH8FD65k3p21jhLzA0Apkp8vfxu/4aWfFXX+fI6p2Y9Gp9dV4R9X
pGRPo0qDJcJtBk6JysRGfqnbTGen1OtQC6RlKbDbpidm9Ri8KNd5VPzO5ton
hU5d9gc1UXtBxUez0Fo3J2eQUSZd+4cTTKDVcuenh4Xoex1c7MEozNuHAM59
Zsei1u4AaPiE7sprLMRG9Fol45Kyf1QDAyjQGNK706FLn3C0c8Po4fdfkjmb
np01V4UGg3ZqLmZ7OzwsqeIcK13z3kf2dPDxTMwEYOKohDZe0+IJNJP3Pd+w
EqWn62rUgAxwSMNi5Uo84Yb2Z2Qh5bMN6pYHZ0wD4lAXKLHwGhyF0qSfAcbM
VKe5ysqOwd4lrbnImrTx+16IVTo++2gzK3raQX0f21gbAUsD/BbBDPjJs3zU
bLcRVQc75AEaQ0Ldf7Z/ROUHUEWYyV8gaC4iogojzP5m9f8nPyxw3mR0nNPu
rt6egXJMtyiibJ8Gke1rGV27Kuqpg8yEINcfoqgOfpwsUU0YJqhK7ADn60ql
p2/0aH1gnajQCjpIKaxp0HlOdkgmGXIR0VCci9/0DjERduqZc5YWxkhnjkxM
c349G8P1/zUyXwvv3WU/74TKAXoI5ilwCaD59iOaHMQ9Pm05J5M8pry6EeWw
RXQ2C/RajmGyzBraro1OuTh9xifOfUidGkbIIgZsOHhJceVRtEEf9TcP4GHW
txgHIZnxzJlMeUL36LwZKyX6hVM/scQcck1HoA6bswYbvQeH0ZWJLzbyoxyg
Kr8SKtNC+B2SscjpF2ljFZ8hfGMT/K89o0ayJ6pUbmdbwzsM/ZeOtapo3GUm
CfxiGQggpgysoAMuEktzbvzLmJsPIILgN3FIWlAmDKaoLcVxxGWVj2L6xmI5
+tRoe1kNjpGJQBRIuM5zkDkLsuqSM8Njs8K1t2iHHyfAS/bAiNG7vzn4+Jex
xEh5WQYU4jKT91Fb1TNqvlmqKD2I1jAokwD5jnrU/wdwxENdKm3yEyaXiEIQ
6KSYSdCGjUQng5yvuQl3zFclQFjHfu7KpOCyN8nI3LaSbvYLm2sjdLuSiUiq
SVijfM7W9xQEGq7Xhm7OsFRrobFU5Lr001o6qxyGyhamg80K303E36ISAy58
o0UXWGYwzondw2AdWbwJjfihBvknH29vYnxy2gG6Xx/Ax5Mt+ku3hj1BZ/0v
AO6PIREg5irccS7Spd7np9eJX767CqZWrP6yKNFxUzCacJ/EYgVDfQXpYIuM
FrmJnRgyuaSitK9nqlYqM+5l/wM5uM2XNkGhTw5a+gf1eB7OPZF4RiBMOqls
MbYqebmSpqWsADNjOP/ZKNcpd91CQc9URtZ29S2kYLOwapA7AYAItjO8cw9F
w6wQUZM/TwAwwuXxpGv+EzLQFMm5cu7y+gcBfzP2XV2ifnFN1Fi4xNDl34mk
dJtCQVFGTR8y9MUL4q4JcMhY+3jOeVb9qaLvyxtWZYaXpvEvFuOjY21x1NcO
G7IUpuuibfopNW/SBXXiHkvyrnU0RFF77yaYdNwe29lCtH0UxEcnc0U4d2gr
aTwrTJ7RtzLLLe4MtfL2S2oiC3UDo+Rtg6ypYBxxFIe0hMdZnntdgL+6bh5E
Wrke3WtlzNacP+RNCc1X0NMzF7Ha+i2qYjzYqHjIUIq2PuRKzHhgyGR7FBBO
VJ80IjH+k0LT3I/YgG5c7GKj/WiiJDDsn0FCZ9ay/hO7RwSo4YtzXaIOdO+J
4wZAkM2xJSeK5ek5SKwwEAFiyTP5OY/s3d+FSOl1HHbqNlgfxFpz8YjXnOGH
3qLQstmd+wLv0H8/1GunBEglGkCYSfFLrZa29OJu8mP3E/OonWzneylKrC70
wgn5VO8QacdieNq3Clpb/9+A0Zy/DKaHvCkX/m5FWjsVUN+5AoBwMrF25Vo1
0+7gjy8keXAd5gO+J0NUzdQSUOiLe1kdaIZ6KEgOIK6cLIdnk8AgJYiJuBgx
E8deTZdCtZbW4Zk1eF/tx77xzjck4bIDJevwCV7DsPuQiO7TMSU22KxweJyp
/HU5UoJ0RtGw1mBY/yXzIHM1eRn1/GPfcDaRsTh1qErJva6+zNMTyoubReqX
yakiHo+Is6F3XQ55kZKEEMrr0sFZMa+GliaPiZ33vGp8JtthUX7KOUAqpnMk
3cT5gQqnOa1N2f7ddRuja++Z1HfOd0IKk8qYFIZaWRTI/ARHWaGxRUfMOYwW
Cd0thKBZCO3W+22+fX7UmK0LCv2+21whVjc21y5TfYNXl/gOW48BSLsGAeAY
NKYw7Fyygu2WVGEiKgOzojaoQ42yZnggvn4p58g=

`pragma protect end_protected
