// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0426h2LHfcNaRiM0t7pvjI+DSqHCQkARyGokQkHcURu1QsSyfERL16JcgRyR
HuBvWZZ2+l55zrLB+Ydh1wO1uLkV91E+BGvc4JgeKCiucNChxUY5IU0Nun98
fShyYP6BtoYJ2zgBv+lsqxaGw8tXeIj3LJR+rFddCRSOTyd8WtNcl3cBw4cL
+dLjCMSk9A5twj4NDcqKSXVA29BnBKghhQdK4nlS0oAoHIlHJn6bCXRtgcdL
SRAO7yIYhLv4PtbmmVgFr+wK8+b7VOXnGHGwIWUNKQqo8JLEMGtNCoTJZLz4
QSOHZwb2C0fWyiO6xVGTPs6iilBhq9yQiXFwZFIUGg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L/BB1bqnNaADjcIwJ/+BPMAZyAjY51mDBfPHXmnw8tfk8+SbXEDEXKcZ66GR
4UZYYXpdd0TbcBsrQ0W1/H1JkT6Fpk7oukrLSqBuyOuG3SBiANnpt47rSuoH
vq2eG6Z8NmJojw6DGDBoh90kl/Vw3QSct9sUnA6oMfcbGKIKimV47GS2ZdCn
OuwxCizos3SR5N248g/tRL0XpdMVSxLAxcnPRPWbvCfPIzLauy46DgNvHnPs
GMyX0B4KYUEk4ew+kOMzADG+OSsT40nDQgJ/r99bikoUc9xmXlGVAtb5aeHK
EeIRsUjb21x14NMmBI98ew9UHU0nwPVgNngdraSzrQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VUJ2E1vTmMe1T7ZHVqLltaDtWQozIOT8ZR68yUOrLDy1gYS2fhk+G3a1Eo0A
H8SfvITEMaGlPmDeAx2YrdGt+LaAWfE+1U1tPOYbXRRXtDqW5TXXzPR8ECxV
k1MDzMUMm0FAZSiHh57A+7k+YDGQO2w3gkbmVPPLsKp+h5Kyqsj+jrRGqFwh
7XnZbQFWubSRa61eOlg21tRW4jb7MuSCpFpf+WfpdkgSFOoXKEF7ziXNiaLX
NhCs9mLGutO6LGbN/YMPzpujxpdG23jAWRqlqCy9OkJ60vTgjFvioazOlZjN
TbWt9/QK5x5/0LIbZHqW1VH9bNEdRgrPZUj9fuSumQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J7MIbuLN2wdrjuEaDjM1xGUJys9vk7oWIBr/wUTT90EPIrmKKcs5e76tgYdp
W0A5+SNL5TwIK2gCkN2FbTjtxbwA4CEFzO/fBgrypagx4T16FuUhsDWxVfiD
kcKcyKh8oIA53kC87+Rkc7CEtzCZT093hS3rypvsdEZUFuQMBKQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tQWv4YH2jrBJbug9cwsPd3WgfEgLlX91JuEcCO3NaJAmPhiHs1Y00iPXFNIZ
cxHl4RqUYVq7fJHjWXwqSeXie0VOOedkVCRygLU84RU2NtDW72o/RC8R6aoX
DRglNWgDz5CMsg/1DDZKByO2Fo8RLomWuXzM1y39b4WPjuB8AYxWCVXSAjPu
LqKxlne9njsFxHCQ9C+MXOpSE2bC3F7nxsNy4QJbt5L4KXsbnxe+PQKcV6gl
MK19N2eqx2CGJyAs7f+avpBYaTEO5JKHWuiclF+vlNpFhW9/fh0Kanz/55HN
/a1Uy+NRSUvS5lzNmldD9PgnKvfnWd0goT0ForTfVUJoNrubemI+85vMYiNv
U6PZasZ9uQcctfm0hyInSReHgc2KW4T4/7OxDvpq19ULsCdsNpvEY0Tmgd+9
r+p6gg+liEzmIi7abbNmz/BfzkLy7zaSCKOoqPAwg+1Lr0/kLIb8JNMMLQOr
5RdQKratvajQglYHX1oHiIAYNJ9Gh4w5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lLeraowQJuR1QGREOCDQ1t0PXl4ScpoHV/bdJqDZW2T9X5gydoWW3dRq4irj
wpU/doiFSfLnmvqUKiuy/q2i4J1Llmp9VVBlGxTbdmVd7+zw9O8ouK5dSmqR
heG5sDhpFm1WCGhlMmqiyxZEVk0j88zEd+ZCA0T3b6MkRrEmwxE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XdNqFQzE6J3OeBuf9SD6R2QAmiHN8w5KihzZmllA+bd+vb0podhnC0vzPGu0
Byo9fCof673vh2VCgrY+yfyFM9FSpLvA+sQ2rsqMMj3g8uJeb4O6qFqEkc//
WcI7cNpjndts+1rt48vw5a52NDVyuxBboixIvBGHpsvJU6a8fSQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
b2gHVzRfOxUz+wYx/DI1VfTPmibJ60srR77TfO/+SkBwYygWRfNXq5vbt4eq
WNn7KV87X3Fk4kEn5csgrf7Y+a/zZCf1rIT/j4UdjQOSuLGy0dcEqaBBkhw5
wXE4Mtdn9AKxopMEKhWS/RypLiiIHKoZ9DQxt1+qOu3Wuwwh8uB9RdW3VtdO
kES9R49/Ob/8Qgc8aYf43U8ERg25oiLMnVOBwzSZ2ASzrrEIedap6sloBimR
uNealkHkhrdXmDbyZ3ZFYoq++33b848ou26+ao6Z7lAGtk27tGwvWtP7a8FT
OizpGH+0E2m8WYs/YlThOjqP0JmD2Q4zdF9xLUcy//ehFDp+tfT1PgX93wXz
KKyBxjgCoGeFrSZcULCpRE9hlktu0kEnxGTSdV88WCmIVeYxFD56ln3PWwt2
WdY4tTaNRZD8F6RmhuH3TIFUv49KfNmwHxpbRl4KOS3k+YdrDbxTXvjfIJQn
DBmHSMyXr5grcJ92UOR7FlpJKQxhVFr6uvPvIL8rFXibbpxlDxbLDBrbXWid
ddiO110IXa0ZO2J4rHZnpvdazJE0ULYO2sL5+c3AiOx5eaDoSeD0TgG1tJVP
2aybdT9mX2HPtr5oAY9xlUFwsNBOWRRh7hWhaf/Nsm9cP2wmsPg/jasmpNg8
vgLcs28LdydTbfru2v9FAdwmj7SoqbeI94mA2DxVhBPqBL0xeuRv7j/kawvI
B3jb/L2uYLYqwXkP6Px/xbMnFu9ar4sqTOBlYYznfd+1iqoNxy1meZTy/Jz8
ORLDpRA+YeR2l99X2JDsxSpiB/pzyNP3oAp6nV5y3VIcRL+bjxFkeT/ter+5
kf3sgrWBBfmwGWosDL8ZF3ycGfonbCnIzaXf3dajt/v5xXlzmCDfvIkjM74i
Kpo2FuS5E3VFo8qQBcLjHmhhXfrcQFyPXGLEgM2v9o8HVCTESiA+KivBNA7j
R30ZiQNk9H0I68t5PWd/UPUNY9G2EqNJehJDCRpKFJ3sOKU4f/oQftk9edLI
Xg95PBOlkICsagW70vt2RqyrLJT71iQb8CRVBbVp30OBK3zFNkKAcATtVz0b
dokclfq2Is0rIlbvr/it6ZVL7ScpR+pUVWy3WRV45XLwRPb0YFXmUARqgLQ8
eTT2tGWsTBq8pI5aXjDQlTvI5CN35uSizOXEVDhsAoUylj1Jjtfi4wMXqMh7
eB1pm0QmiZVD7SCvUENMAA/c9U15iRNxp+Y9+GXU51oIx0EoEreU1foSpBeT
x4LOx6RKBrkKGXb1PlQu7bhMpZ+FZE2pmWnF2lN69JAxyo66GTF9OGl742d+
f9bTyBG1j7/D9UxRsI2bYedzfg4MMnC2wBPO7FP+yhTWKD3eUTM1yX5szJ/5
3JbPXbT8LtQihbMVD8fwZx/Qms4VQPrsUiB3t7/ggA3CLUvB1wdnlKrb340h
YXTRg6yH7oQeB+JNqe0XVhQZPmJCP1S5oX1SLI+HmXd6HWjiK9fKXfKxCn71
FDOMw0Y5cKH/KWsecu8XJl4fonASCo7bOcyVkHQ2GN+BCM0+5aKYSlTKnZ7p
ailw/IppUil4nRjPtwATMy7RKE+GbzYzcOKC0vGI7Kf9gZH1/19pmJqxFcmA
xkrFKzYkZ7R9ekDogpwgQkYxjxkCjVlPz0udWr3hMxIftowtiARbLfE0rKAY
U+fZUIIfTFIg2ybWUbSTMXHgxSY=

`pragma protect end_protected
