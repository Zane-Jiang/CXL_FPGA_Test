// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jdsjP+nbGVYP0Q6Xw+T7KCvzDd4rvL4CLQ28vDJR3vYlnlnsEhhqnjJmfKNb
K0TMj7rePJYHYsD8DRYqmq8UeixzngRKsKdHZNBUyRMQv3JX5ghME5mLzAnR
k+9O2eOBhL4MrnWDGDHzOoMfdx6Fyb6OX/IASCTWpbo4Y0vrPg1XTq/L2cQE
iwsddrl3jQpzOxc9wtODWEUKYzF6AQQ2CTeisISSFj3NCeqh41ms6Tm2NonE
bAlK6FAw3Oh/xF3LFWoMPE0fhCVWIoBouEGMV8BR6mKUSCU1Y3/P5ShEZD6o
nA5X23+ZNwTj8UpxlJ4Mf4mMoOs4+0M4Bwm77PCq7A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U1/oL/bLIdIOcPdwcleCEQQPS6eP2Xmk6dDmK03BZtqcKgl7iCdnrhIfWSaD
SRSTJnv1OfVDpr1lqjJHBvxYvGlhlTfThxKXXlXOKkHRjeCGdXToKDTLFnf8
Onh+uDdHV4eUAeuc2T2HmV/bL9IZNo/VkDi9RIMW59Ej41Xt0tjSwBY7vO6J
HzdkNobtAqWAiS3r0JzowoZzrPtv8jby/7KRl7XiPJ49fWIi+ATteQSVF3c1
se1UQlimRxDnaGIQqT5FyWPScMTLuR6eIjZ/XNXGQNheQWggum/XiGiubiX1
yRnu4qcaOJYclsHoSHYLzttNZeAxThcg/yEh+/qwow==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EIA8Nc6oIM20DUtzc8eiP+LH668cIcDdWCPh3BB6BGwG5rjZ252XWyPy2uek
uCGAFesVkmSdCZAv0RMb25sjuWyu0IItDsALJfbBoCW8KDqBzeow4liCUC4c
8gWkjQ0VGdcJ0gqZpQfVDKbdcZaUK/5Ciz+OA8OuF6CGPjqg3zayu3hmHzBb
olm50IFiFxN3Clv6mMO9eFNhemep844ksqv8s0twkdGSdZPxvkOsNanqmbIs
4NspuQy327QNJ44nM0/UcwlT+lCnJmyAg86sADAnu0Yp+fwWGWqSYemoFVuW
3MgFqoMtOonmHvHFa5yXCIaDiGnDQ53YnCfmIO4N+g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Cf/TyBegmx8La/8cQLgQg5vi1wyknAt993tverE4ksSvw5B5ndw2X1Hsj3fX
H1ZYm4SVRFtNJuydW9ZcoEfiYyKDfR6i1Ca7W96k1zzNo8rsbmqc1B/hhdUb
eZ7XybA57Bsj1+y3zYC0EERTPpRotQdtudL93NzZqOmxSI57IMo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
qlufJ3SeRoryl3m2ji04Q4bw2lnk0TWxX9ZcSJkGOapTu5SdMht3D2IXwsDa
zLLfFkctM2TsI0yG8qq7x4wRCYatwsFN+at12JE2/xxbxfcr4jiC8LX0fIM/
JNM9NbidmMP75MbZxjeMwz+DCng4lVoEag1nreB4ENAg362Sy0pB1zwYezL6
t3dZ/YNqUxQzq0hGZX63iH/Amih+mFpYhUiW7OP5tA6wANYOMDI9xEDfs6EQ
IkaEW/UWfbvsJQzZCcHMVpyyWegqZCzjQJCdJlJpBZlfwJn7/344dpxhfrAl
cAWGqRi6SbcYfh5PkL/yfhrIhelURhT22FuxB73zJGRJSCue1BNntidRn4tw
o5/nZj6AXwDXS8d3IV6Ouu30vMFZWmXUfqDylx5QS7eEq3Ri35ipQj0PTOQJ
VxV5udbfZmwcwAW+uCek/1pQ3WFaC+RRraOpX6rUMvJvf/iiGoPys3g2SE4I
3mvhsEb6P4irJZYj0tVtAwCOehBd+qhr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AZpIo++E7EKYjgJkHAXEomETc41S9QR2BEl2AEmXZ4V29+Q4+hI1H/iXar1y
vcJb6/gFCDuu4/lbjrlIuv4d8ZJogHzeAUKrxa0wP6Y7we1Uf3R1LyCEqGI9
+LFEQsJM6M+yC8CxjUISBAz1ymYzEb1fTFgZPLROKKqPZ4tYgA0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BzTFFXLXLpOH1GOVwX1fowOFOWiOxNKMQkYHztq3XA1OHEcx3pJ9e4MAZVVC
Qs/zJunO4PWxZIpZh987zK+rS7XZWJt9DCWcOk1jfbKLkYnC0TyVOjSSDHoy
IaSBQI8cbmLckjTUfgNh0S7v6iU2PWhcHlnnk74ILxj8KONOmgU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
PrrQplhzHvPcKOTF+asRug+D9sBv86u0yGgPP/PnffcVtXuZMfcJ9lIZfkVh
IZZ/awjRi5oITnJTEJw82Pvt0kM/3ZaCiVXm7vwMk9aHNq7swzvQ74hk5M10
cknO3lEMWcbzR5KR2j6DvFYpdW46oaA/2CMvwNJlgHuC9+Y6BuHHsEReuPeb
Nw87tOzZNLQ5WG0JKJoIGy/kLwgp8pACrb+K2cxOPQWLxFqAMIRacTEieQn8
CnX8rCa0KVHBgTXQI9FAqFX7MPK+TsZ1czobvp+0TokrOruqAqDhCgtSC6rN
lK8KWkAnxDKHvj1GlLIS3Ewy89y4N0MaIQSTdUWQzTM4DYLyFE+Xu+WxbbHl
OsQl9isC/xsIqG2HwpHgNvrU4OZzfKSAfXcmSPVMrt9ssXHvVEGgBpEAzCzI
5JWOUBELpeT8jxIVddv9p7X0bwmrQawBuC2EucAXBrWddsFeN7yftlNBF+sY
Ee7BRVJ0K4qPgWx/xvpIiL0pAYsgoFsQU0baGVh4C+29R68PtqRvvuMefD2T
+9zguLQUW6LMWgerv9hS0qyG9l8uqOegpOCwnYPJmQMOboz8HVbKphWDg3Md
/3KhqzsbCVAPSYnx4f452TPhUly9H6MPSPqoGOoYF6tapymKyuKLIHiF5ohg
gZH3VG+pZJyO/SPaxGrZ6+WLLYGZDoi4R5P6Q8ILTFGDVhdROIPLf4qsDYBf
+0sXmPNeUOTGK2pbCuFkL5tyuUVlpNpK8h4CYWdoMAscMaOrko8FEd8KI3WF
Ihy5q90mmsH0zTEuOHTmFP9LALF6F+7mtyM9cRNEvjC5XbAJp+JA8fBsFGw6
XjC95H3NJUWCLK26FwhOxn/DL1RAhpNUSDtOxX6andWCehV7TyLxtzXl81zU
ymXymC3dRFKw4TL3rAxXZfTfGeZLX94iDVm0H5Ufwbz/zah9Sehfnznv+YBz
dUlx+bFjuUbvXHt33Yg0aBqYZR072PEx9M6DPn+NJNAXpXU6pNhiqWL0NGcs
xfDCD+yhpCmAgJenxcdkfF59z4vq7niwNTJiIU0XIXx+GQ6iIda8EqLLyEt/
jY6O9sljF4jqR7ciM2c/ql95cQ3eW0KKE1WRbeEl5HBCz8dfyqgN9CGX4lfn
OIhy3joqqa3wobCgMlTweRnbg/JcF2hcnGOQoni7KEfMNuLW8xC8b1wB7Hr/
dbYn8MDkZiXKwcxWGB4/QtonrVnSG0od6nzaLGNS+u2NnszQXljIIzVKXEmZ
m85JZlGHMhz/CmaHi25FOONV/YDPVmtfHH9f23oOuY1kyPL+J3OcpC4ZM5yM
v7KOUHRrdsuYWsy/kWSXmXekv67o98HdKHodM6xJbxV4vC8wgyG/DkLaw9d/
up11h5Y=

`pragma protect end_protected
