// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bhvf1NDPmglcu9s9rFE8fgZ78jEz6TQw0Gk8s8mlovGBUIBfDVh/aLn0fOFg
OcBxZEcc1FTXC1BBsMIx8UyF2RFrZg2XkxiAn8ye6lrtckih6iKS059VylvX
2ffjb1lalDu+oWEEqqLcxmT23vd3o/a6tTTu+piJfqT9303R2F2OfPURMLGD
kfL2QTu2xqIe1UyaAlsSaGxIccVUQMzhS+O5L7Z7VDK/vOvb2S4SlZFFAluS
jJe3cgi1zqUgj0YrVe0ok87KkPP/jt54DK0dk0rz7bFXM3RRaWOSbJ2A/lOm
bv6LfQGbWscevwkUDEYuxiM74Qr7XNsetAjkrvUeFg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qvS9mHe0MXN7t6F2Gc6g1r2zJw+YzhY8q9NTBLzQz49GHXWJLGcib5RBkwul
qaZv9cdGRfx8oCxw+7W3gaflnMpqoE2BTnqMbPJP6da4eZtAuj7pYdcMsd6t
L1nrzJSHjq60yjEpYck5r9W+BcvZo91uvmUZPXt3/J71cE8gDpWDlJBL+hte
pvwyN8yz3cDtJRPDGoy/sztadUbC9QflFPuFG/Xp82Auzolc2D8kyJ/IF3cP
xC16n2xEZuulmsJzyETHgfOtkFglbc0o4bAfJz7YcF69QybeHi18WArXSD/B
wnGROw6ND2KwIVOkBWkD8vP/ZLFweduuv8ZJ19VFkw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ibPcH9RK8ihMBA0PTG4dOC8lSoM2SO76FvdzYP3TCpeOxtXeW5ioc/jeZhdO
E0zrtjtfebGLegB2bjSItJqftkyZcbsZBz5sBicnnwbT8N2hhZqVp2GESd1q
4CfTgKQHWgmkkc6ELi/PFD1d4tnBfYK6xhms4mI7lcahv7pnWtnZH8npPuOi
NBq+AzPV0hDZAvOzUJ7VmxegguWVEs+UXVKfFdJpNyKk87bWh9AYAgj2wn1M
G329wbhBycosDzuw0XSPsiV3agz3HHHuahoBp26EFtUBTabGbS1smu88Amc/
1I+bghaveGs4j5QWHJGqepdnma77Yo8Xjw9aY0t3zw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C826eUQCs/Nu2mMudn+Ruihrau/AiyPC9EprrZuETSxqoZfkq5TJ2gQPDzBK
RZJFV74XEXrOUFHgafWe+F5Xgcfktemx0cKSaxciWtqirfj2AKUspTby3TE3
IsODK4OH2/7fB4cSqcf/Z/M9qslXUZaLe9Z3wbHon9WPt9+ZY60=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
RAcuxE5FE5EoDP4EvclNPgJdPvckH2fFdJIgzANSEGZ877sn3uamuKBXopCs
Feb+QibVt85qaRXd5gcMovcmteODJ9OwsZjPZWP5gY4e2Ky41MnPRCgwZSOL
S68WMFIth5mtjC/7A7fey6CgbDzBZ45yXUEqV4L2WABjE03voRp+4cxDGbFK
BtJAT+fWHd8BMSN7AWO8WPbc4eePw8HkE2oqybwSBRPKiaK2e+MOy39prhV1
VSHlvqdHjw4eDfjyosbAIZicZNq5TbRhB0GvJzjUa2Qc6Cb7+rk9rN0uth5n
dPqR9iflAHVDgmyob/v411qwcAzf33bxqzOc92uuHZaHrRgRQCfrFFWcumgp
ZH/0NvV8U233/IlNI0h2YGmxHgCu1KlRL57tZ6TzmPnyhtAECBJGZGuW8+P3
K5pWocS/bzLT3IOJSPINAeJlzJvoTpPYc0dPumlhv6KcdIBZUZ22eiXcIjrN
zQ2Z8mGJZXSx8yJs82o8MhGv+yONSOAM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TWJdyP43uF7CEXxUn6HFBpkJYxGJSzjROKAgaKB0oPjtjZamypb9Ijff3pgL
55NY9YjfBTlUPUYvLyHlMB+voA7Bk8MMUZt80QYhCEUgcK1wfuWbd/oSwRxp
ZP8DeF1/zMRxpxu8kjJszC6oimWNQTNQaiMGbszFK4VE2mmVAXs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G5QpTDGIodVjPiFAUyG0dGc5F4oe/9m5FAIJn3PH+tsop6AHc5qxZ2+hw01v
L55T6HZW8YDFKNxdccS/eX2E+Ts9JBavmNYufkR4/mxvVIEH0jQb9R3/IRc3
O6VDJ59qyMIFGIMPZymjw1XT10BHUBK0pQhB1eKBrsBZsnJV3m0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10016)
`pragma protect data_block
r1874zhVLVNSZ+QG4enzYCsMZ3aKVW8zmQcG5VXrk+9Ig+w3nB6d/bU/lM8u
701+m5W1XUjjreQI47OChadSJ4y1tRe3cisUnrPiYgJ2K00BDIIHepeLdIDh
VcQ/Ivh+pJoQ6k55YcxGO5sviYgB5eTHT3dP+G9QYdZRAm6SoQiRg/XfTbMe
+KfXYsFo7uKARFWC8WTiF65yGY9MgFxdeIXiARsPwjQCk5huqJm4De4aq7Xe
5JJMQfC4mXwUSb7ldUiRn9e/d3IvztoPbuTlY4v8PsgPZrCMphYF9hbPDjJq
0dHnuOT6dBgvqTTRUGWgEtmnnZCbXmAeLIVsZ2GqUhvEh/lOeflWWjYzOVJC
FSI/WQiJHukP7L9UiSycEMfbBDlBjn5mqp2RrFYue+CbWz01HS2zoDZ5XUYL
CZVkXwZDD/YX0LmJRpTSx2GNbNKNmv6VClAMg7oTkH/AyjraXaL94GlnKUqv
J2mdx7CwNVVGPvsCQV20oVVWBg8yqGKHhDnl+99/Ra5iYpgclVqgD4l55BG8
RwkmvTg7y3YQnhswoXWY3B4PWAjmsxwXDorP98+lbOdPmSW1KGWP397flUCa
LKRMb+NIXL0ovYY7a0mLMTdkdoUpoy/ungnRULD3lv9I8AoyMEQQDvaC6nGQ
tZej2gBBO9kA8T5NyWU/rr4FZmzrEhSu7Ux3L3T2nIH/NXqxXPWZ4Z8U0InP
QnPwbu/DBpXGDNGCxir7rl+zv6srTdvB5Qj10jgX9iszOGDiQ28ZjfmHYj1i
Fbu8s7whhaRwt4C+rBKCWXfi/WBCW2/DGxIsKwREIrgQyQZNDb6f/LWMMpNi
xdEsbYshs7vUQag7AfzrRxWxklDvKPnFMB/LbzPMPitp+kIQAXxBRFIDPGcu
eAk0pT0t+/WGdDD+7ToT1IytbuuWLzZwvBS9hHHilBlGP/04kiZL5cs7KSKw
Vn5081qrWLVu4YVrZSXuO7qs5LLbyadf+uzIJoIxZ2LNY/Bnn3q+ErDHT3yB
Xij1E4je6bAQykDxbYlCYXTrcDWfXAYplnpuXxjbPi8vZxxsva81OKWEMGrq
IchN42oKnsC/3gr+bhwIJCkD3IdjWmKJ/3v95FqrxQrIxUv5IGBsPSEEmVYo
HiHherz22QfsFZCfXCXVt2i9j3LoXWoWzxQZoyOdKh6zRhPuv9+5FTzYo0P0
wAjHXGcr1pFqotvLUo+Xi4p78iiXw6j8kcWRbWQZrsEyKFjeiBINnZgKuutP
nx60R4bbpJu6CbJb9EeD47RxvYXRLKvXETZ8Gl25tG4/d+fCyZQ0DQPhTTFw
bZ7TYCi4iSv0lvvTgDBCx/Y9dSgAlUY8JkqV7OkIz0jXKRjR0myESYATbQnr
v9bLvZSfCg/ncLS70nMUxn4ZdeHkfYTxrJk0oya8svingzQBISYB1XJvZYa0
/kepjlrkQIo1dWHmjCQ6foxvmMxDkJzZI9jSHOZPOa7fJ05UT4aVNUqeZNd/
2ya7NPYeVTrpP03HlAxeoATxvdmoJ3gSeZThJjUYwW77CWwXjlAzjQ+afl67
NGQVSrL2ZY9RP86bxsFttHbuWxhlYQxQD/xNKZRfQ/N3argC9MZdlsz5bSmM
oMSP6w/X/KrSr3GXUxVmRfZghavD/XT8OyeSiBkT0Gdm1vh+g8Ke1/ANzKbY
PxQ2uGbXRYWFSsuLaAv91ga+PgMnpfJQDPPaYZzdmVLAUHKXYy5SS9Ncq055
C+Q10g1M2Wy5SGk5hLf1fmaEMgnTg4mQ8bOzJX4elWhD9FVa7lnVtDRYBHFn
ET1n4waM5o84ngxDT73T3autrISqWstLlRi0Ln7H9F8EgAhvDIMZ/xKuHCms
t/jys4CjyVt6i0AFTDqJ6QDwzJrLQX1uZwKdum06EvETnVlVUNMp6WCkC+Ss
DNNw0gmXWfV49GBe1WXCYQgRnRPE43sGS1RzmYMjjcwc4n9mM5rLAbOABjcr
D24mHfETHHqd6PaWAvHpsCCt0/+l/ip+1rOypMAIhV4RnzNIvE3tmutXnhWP
1DDbm1AjPCrbIrKhTJnsSENHKn7JHhPxwDuRQVGDONRCmzAhcACi2z1byH53
byN35MJAoxeagEvHpJoH4tvNh23O30ToFZ3pD8HXSA8946eSAaP2guUQ4ciI
QehbpuSkJYI6o9F23swnvwb6gca78Kxol5DD1HY15lB/hVraZxQJi0r7p43o
rwzUweFnt5MKqMArpHKZ2LpGcwY5kQUEuH6OAJ0QO33ptt5zJjhWf/D8vJmA
IZV4UToJa3tZ3zty3A7jYUgj8ECB3fOKeNURLaMgSuyGfj/b0q4krf1oRQT9
fd5xVHT+95ND2GTecdbnTAI4lFBaTwg8NAst5nx7cx+cyem+j6pwFjOSuTvN
NYkkBaWwNorIxcU06wIUKz+fPAZtG8BRfdXj0ky7Aw3ohZeSv59FW6oE2HY1
nFnNEomNnyoAHzUTindMlBqo4IGFryNg2Li5Uhx2Bu3i0Fcd8X8bNAfnudy8
K29NYuoX/c9oZlBXF87EV8qYl1gPTMBAJZNRx+YXCfZzfL3fG1US9lckxhA/
6Rt/IBFfIfrAAHAfH3e09v00Ft85/FivY/HRpEIxj/50FAVRpcFcdhg80B49
4MUsHq3v5bX4xtsouNJ+PKlAapqWaxratZiZvp0FFx4c0HeiJHLB0C7t0W7X
2SFn8N6FRT5Zsar1E59+503HrkT1CY3wDJHZPsDq/ihto5D6PrJ5Wu+M2G1X
EUP7WmutqnejdoyDNQJH6u3aT5UejMG+lY4RfvAAubCOtGYCw/jBNem2ImQ0
RMYeExI85k3COtfJmcEQ/hiAJX8mjIjY+cTOA2vH18/aeyW1vLfn6ncJDdB3
zJ5mlnoXrZB6MgsG6v25NLoGPfd/IDPLL8acnWbYEBywdiVSTlRvtz1wxgFm
V3gilgqhPyQGr4gDdzlkC1+LaS0kbUl3o49lz4Bm6K81LMESQV5Qp8cObrd1
xU+Bcrr+KVFwdt+pTcI82zPyPl3LNYupt+fvx/ugVfYxfGfOIp4HSWrqqsck
25q31oIrURugDY+gtRVPQ3qZu/dNm9l5FVJxjxpHTaE79DxJMgmN5cpDeNk1
+NeBrZaqgEhUrgwoIruvoejDqcoUiusL8kGs9Ct9vMFwmN8qELNEnw7GdLvr
kdolOdisyF1uJE+jgVTCLGaTMxXCI2X3UA0d1ohZbAtWAkVlHVQgSTYCf/Er
QsEX19wzD0fti4uMXuEkzxJ/IOZLeKBJEmJma2E6BMHGRPtPHv7fRWld1K3L
Vn8K776EySK+Ny+rHvfiWvPFS8vgogXKqIFm2+BWfyLJWv8XhVn9z3r75u1X
3Lq5o72KTMBJ8Lj2UAhZluwHzsOzg2hk5edXRh319iAeXy4N8r/7sJ913Y7x
vjZ9AaRlinQVIZcitKubkWMSadjhl7lDrEwYiPUHI4TsAcrL5KnLTuOd6g2/
4CPPfan7gIrjIIUf1ajMbKI+Y7PS7nH6CaWmfg2LU34gEGSkjk3JjZXvLP7O
KyWHCvJy1OQU/sCxxKBsAOJdsixIOTHqq5CfxVYbNcVrOUhiJXTJrt303GU4
xZfjfWNL5hr01CAId28BXkYsUdMdJqNckj04F/LvAdiM+IrWa7VLPzVX9yRE
hd8JE45Opg4OW6VnzhdJNC5mD5owqdoTVBosuczR9zF9mBKOLWDhIr5t245D
nwjLl0swRmjadhQScJV5G1UJlffkF99Jas2krURX4Agp9x+HOg8xN+FBJUTo
QBTvJ0H3RPM0TrlmKrpULuCykDHqSfuwGnJ8ho36d3F4vOGCMS8uMd6yxdFn
wT4jtPNFmp1Kj7X8c/4CFYg40ETaq54NU0bfuiMIMRlxXPS9F73YqgEtEpxr
VMVzYKfjf5bZTL8zXs2bY+1VnJtHbNSL1mvheBJoKJDudXIL+kIsL9Bp3754
aKQPQ45vg1+hM8MdRjBW6evQXbSnbMQMJA3tLJiF3GHWFgy0UAK4z4LY1G6S
/eJLMvVTZPx8qYpFbSPQvMta3lB3SvLOMXjDbq1PT+yGmgNKTBYIh8BLv9t6
1t6RBXz9LO7naN7oGSdQrxNkw4C2zBqFB+j0+k/zJ/9nIaBdyVNpuvxwHJCT
WrFq4IbzRjn53oQ9sY8Ub//4fjp4ze5X4ciU9FbEhMBa2Pm63dwzTZfKtl3y
HpLr0ga+2AaoSt/Ni0kbF0S0z11YuQ3m+m+bSaahDjUsXVor+uqml5cJbhUA
IKdRx+ncBjkTwLnVL+EACduiB+usKPoUEmd8V5Y7dCNMrzy9SxSQTTIh/s75
aDeyaDbLnLrfonEwMaYx5l/rEJefGiGxR8iGhx6wL8ZODfmL95rGKZEQmsbr
ZbkdHSV+6rQ9w+zsgMyI2Av20mwH7zkmEPqHm7awbap/gHlZoKGlWanNsLNf
tHTm0Yo486sBQhK7BYdXbOMhey4dohZ5IvTdThOLMGpkjpquW8yhXKuduT+8
drIHMWiiz7BCRFdc2BSXdqcoCMedS2oKkt+flLZuipPWgxQM5VrjXDkk5hJb
a5fBMhJPlpiUkjhgi2PlZLKdN86JBT5nkm75soIEzwuWj/doAdzupawyLOWv
cgYQoRd6jd36Lvq3MyiEto2mmXzZ16pmM04V1L5WYxGqOj54I+0mJnEhWkh6
jpoCepUoB+wH5QVI2sZsjajShK9JmjflnKHiAt6jCKSUEG8mjCMDaKN6ilSO
dQyQiaMQSDNwLZYSTVq39o3Ldea3LN0K0r8uA6A+tr17l26zlWhi1U8uPAh7
02qWdNecIbuwm/ADZiz6hXmQGEg6Editngl8DtuSzlWeNgNfJJn1zhUtklO8
9bvVes2X6ktldM0PG6zkTZ2tMPTd870VT3DqfT1sWkhzAd2IZfNs1HiqOew5
EeZEU+Rhvzf4voyH6QlqixqqTCJGgEKhtVUC4sAFyfzYqSYX6Cxeas79bRir
kodMDSZaVFGkcxD78/5iWGn8WKeW2tVEnvHRyu3sX+d4lZU+lWC1+bOo+Wge
cx9r5+CjsON5s8CZvVAZucSP/ROp/Qo4WsU1dtxIXuUURxy8ukC8xE/yviWf
gqXDMAWxXEFdUpLfs8mhKFgXVnv1pzk47wHW880Qh7xNaGE7VU/7Jj8Oqw/R
zzta/56XuiQSnvw/QVcodoBr8MXC9SNYyDlJq94EgjIWOdy5daSM0ZBVnCGl
V6qVcv7P+B3o4xsC0SjtRn03vGg7Aiqr29T5fGUzBYvgVxZ3AdAclJXyQ/sr
wDtmR5bpErSnrRz6OOExjUn6hHpe7f0jS+Maq9acVsrM25jItAkFfKifkDe9
965cYGGgSoovZd0ezJTeCka1pMDMD4iA3VlrVDtmueWdOZvRtGzHrLkdJyFF
/DgeEBJFuHwgKTw5/1MYGSZd979FbG37/XWOz7Xa4A2SnRBBYgwdY3gsm8c+
/rNiwI/54583/yS5sn4cKcMwSMppMojJUyLxynZvuVXwI9IExYoep5o6a/7H
fTUvqtbsESXsA72oaCRKc6DF6m8MzA9zD+E8v6n63b7rteROW7a8KYiaYPew
+hmY71iVXbVIvv5q0xUqTwp5GcKZwMutSUwOpdD/QCh25Qu5ee7lecWHE90B
fqDFWk4GjqeeN8GyPe4d6eyFrsjQRt+WWXefuoIEVuAuBxNvFwK7UIbQ6gFj
tZuIn0wgBJ4E9EPToXst3Kg4gUMqz7wKg2EmqflYdwTNHA8nS6V+hfhQT05F
LFNWJu3q9cF5l6paKZmCyG0Qh4Sior26diHDSuv+9zMsbKyzQ5UIsln3wrVM
2NnBI0kIz6upp7n8gXvkaWuPM/svCNprPfDI0SV/BVQoT4ktZI1dAi7ticY1
DyG+vgRZXhGYK8o3Nmtn5ScpgQQe2XBfXGTCLDzgoNt1WYlaJwJJ68KkB6KT
J6dIl8W6Ge9defQ6OPukOQZm798ZhZxN/JtP7fj56qCdeliENBLC3uyhu+w7
cWh/izZ2QV12kes7/BWZuVx6uNCf6LH+MtRFWsXbzKxPln0ohnRMSRSEEtw7
wHv8gk+MEXGQpkSZATjIKw8FCpzRSyyYkOpc8f/ZtPXXrugnt2/+g2+hzL/o
X5fEXM+Tn9rzpudTqK8wekobjenGu/fvGjoPQxORbVvVFXDbKfAIesdyxjkf
M47mA4xqsk0ypKHRsxybMFEkfSd4uNZkk4F7Hqdznefhjd5FzH94mC3ZuPWJ
bUlBeDxuwo3raI0uqxuU970Aa6kueU+p7xTqRAakbb3Qcy/QFILK3HcHebYy
oeZ27JuL8WAQjd0nmf3ygebm3Y7hFfLNtC9zOax9FDjP2SQ4EU8XTXWjCCn2
Xgsa9LYPNHxZOl0//SYWGIz5sAGkL7fePOULwta/NtoP7KfahdGGbAFINztQ
D67q47VNsE49wDx8qqcr61m58yp2MiS5IrodXCS6qR8OWn3nm6pLgPW5TIwk
wIpUelsJcd1uwsLoRIcjQZgbFZ3kLFGuAeIEJ+7FupE3Uqx6OSffX7iBNqLQ
zX1SAVLs+YLfVKRRa9LIa+pA4ZyYbbI8eqk6Q6zdkrXUDaTulhuR3B7CHsxM
GyceO0Sw/H59jocVkvU+38gVJno/IJnvjZILz5yazZpaQOQeAaXr7CEH2RNt
jP/b4gYGUlMGao9Q8EUHUieCcF2UVgryGqp60grhsrDum2GGy699dhU0ClfZ
14kMEzknQ6uZhFQdBAnKC1lryKPPsssx1gk5OgC3IqsOwtQcWM/Vlv7hMif/
b6ArS0ofcPKyS66UjorCT3MiSEomlQP3ZFOqZP1vnjmFSz+LCTMYs4pMXCou
v0uGVcZHcGHsISkGIDIfq9DAnZwiu39/Q/NB0v1GSFPPLV9VUTm5uWedXxsx
LbJxoaeCUovE++KqLCNnK0hyK4JF0ngXXpGYiVgV4vdD1JkXotaHWh20K9j8
ymtiFIVPd0QUEPd1TdbXpEXHKFmbMI5wKRQaEHpXp7leQh3wP0t9PB9BIc32
bQ+0VRo3sQSWmm/ktesWnlkTGDx8kZFWU7clmVaTcqXaqyPmzJqlMVG1oTyJ
LFl+VyqmTBayrxS0+1OjUCuwczNQISjLdzjECcnZ1YqqurMzbAtXBExiSV4R
FhnOrMPmRVzjKZlCvzoZUzJtr5Nb2cXpX3TgrMyaXX001UMNk00MhYucNhTC
RAoMuyP2G2kYvtAbqw0Hb36RbIUAn9cifs7YnysWMBD56zSW5+wj6aGLbcTq
a3LtB8AHH9cxuuT5u2NA7u3BbRjc0JNtVOeH2iRP+9q31PPOWst33vP/vbFK
pJ+Gu3jr2Vs5nAVye3e5D/gUbprVYnihwR3f7vf4Ysu7ULxSMCDCDBh6KM1Q
dph7l37duKpV9xDu5COyyn+02r3xziJDRVaqjLF2xsfOpB89LLW4seG5yCSO
T+bOZ+LgGP21Yewfp08laaQstGA5Ih4JW9h5bXGsmCXTOEI5ZiY88GrsVT5J
ZdPxgAjQVwmScLpk+bh2e3M/rJRXAO9HksBHZJlH5DcSB/rABMc0RTkdn7wq
czFnUR0KwjRq3xf0Fc98tpIUGAhD19r/XXij6L9YmSvlrPO0cNErxNMjxltI
cH6QwqQBF/IFtr8Mr10X4eEA6lvyAVASY59r5ScXsITSX6J+qRbzVfylHSUJ
CmfhE5y2NuwNw6UoxgXg4GKbl1LhoOvR8n6UULoZrsTeJyOkoUvQv44gik91
tPSmwDWUmLir2U6mKcK4dth0DmyOg6M+WSK0BOE7MlzEwRwUWV7J2cdO7nVw
KGyWnTKCXCH21w6DbpNyvimayIqBbE/96NgxtQOgmTjAIwjGOb0m0x32IibL
Lb0mMpfB3WbWan3ajs6yzfvI1a6tAldR3dkAOlf4LrOzZCXYz6tBVBYDTSK1
6nq24lOxiRGghfFGhsKJTY8jgvJ7+jZuh94RsUW6zoJj7veE4cfQSu1TEU4y
ihj9jHIgSaG7LJa6V4I4QlLL6kL2wfhOa4oBthWz6y8iIrcKqNLEYQXPJTxH
jXdd+a+Bl4sHckHeQQ/8vpFVG1gv0wdEc6vkBAsYPffC6YILv8tmb0nMajNh
/f9Wc/78z7fhNO7xaytJrqp/ms33w9wKg9mysCQUfFo0opZwJGsdk19Lt6c1
FIU7NohX0f3NZZd4njPOLsujR4fcPEiDRdVUeEiFexDnndoyJeztt38jB70p
D3Ed70JCQha7qooipEFH571/j3jD+5YJ3c0ojWbCvaBcEOT3rJGhzteWYC6f
b0FIQA1v60Vi40SwUjUUNvtc9dVN3LS3/hxJ9YDuVakKGmDm53grLnNrjfP6
2pl9s5GDGCF+DAhN7k3zSwNXw+d2EJDszgNZFws0ykCNY+n8m6NfDADtb1Ev
fBY8nnMWXpl7WCkZ4VM9uF/l7riC8lgkE9LgEeVGn/3+A3VbH4yYCrzD3JCX
UWuKwnaZ3r6MXywAL2/YkLyLP/g9BiPsQkgzCNxSSCX+N/rAkkPlR33bG73C
7fDGBCIRsjzsn6CeAATnp+iF84ngc5uJAMiSesl1+P7fSH5poj36BcRBkrKP
WMCXcqihCSCfAMUCNB8hmlVZNNb4dR53pU3Q6UpEvACl3eDLj4kN1ucWapDN
Aj+5gURctVBxlBqv3klTDHepGzqY008h5tcWkC5YA7aT0iJdRczHfORyhXxB
4WjiuiMWl8L+rvX54JVlCrCqKTzcSBjjx5Rx4t3GEJbUmCaMX/KdyqwpoXNF
izc4IY2sScLyQGHKuOC9+JA/X23IstwVt+TQSEVxoz4x6Gow+rM4eDzo+V9L
f6KRLJv8KnsxUHnEuwyNIQm6XA5ROUn+UEPD7uX3TqDEoXockuI/hvo1b4iv
0fF8lPdf1DyP6256AYp02rGLYSqzCwSgoNV8bJpCEJEsnq6g8NYVzNPGtOPt
pKIziz57+hrVdxHDQoLjlZN4DMcWG6x9sRbaIz55ntPI8El0o0h0Q288TDxn
RjS35+c5I2GDB4Sb4XAskRN3vN48YENHtBPmWtvHYUmhnelW1xVB2OZWNXwt
iBvgh6JRcdtzyryTKQfhlbE+48/rFQQtlE1LLNn2SBI5cBAZ1CMVgWHyM2SJ
OQaVCcCwmuWxRlvqnaPhBG5a0qzIeSktFkOUeRoZZsZBFOI9afwO1E/PWkHU
JrxT2MFhPcxyvEJXWAmbYgG6CtIg1peYHn36Sp4yyAsgZ0QNrbKrh4hU+WyW
mP42gF9RgWgZna+MDGI/VtHUtO9je6IR0W0h06vnwnx9tr8c9y4XCvl3Mwvv
xt6hf02VI4bkmzHoiN028iZp03/U5b30YCKkNGVZMvgSXBlI1+c8DLqKcj9Y
XPVcj7Y8bsdJ//7XKsd58LR9Hb5xWPoCUwHiGxmv7ohndEdyAMoDb5upikiC
lKWcEz93Lz8ErBKar4opxVA8D7Ws4D12O2ZwxFKVEM1PSFCZxYl/gS4m4IIA
dxbrZKjeF7Nwuzo4u5Gf3ztHGeBTjzJffFzcpHGcdWG21/N8GMuxV+G6q1Fy
niCIr1dJcXllZnz5ykaSp+dXOAnI6OxO5nJpZZtHKrbMvGuVewRh/2AzYbIU
m3xDZirC63mMBMT9tuhILpr9UXVOv/0wJUTI81FVZUBjJQn3c05l0Py9t4Wi
q9gu2wdWPJKgqmoGi1yKBRlyYTQTZ/yDc4TrucYuq72X5YFFYfEdfzgIpcZK
2y3HDK/Rvx8iW9YZ91W4bLESuGlOxH9s43veSziFLOlS2lYwwN91jF2RDQQa
CZk4TrxERdoVmNYJRORIG2oeH5zs/8Kpn04UUAcFCvOaGfuS4Hr9Sv4XKsxo
2jgxE5iwc1l7578R5Av73z+qMyoDWCAlreVqL420BCVWFdXUFUZ+o82JRx4F
+pvBbgwEA8Ikn5AQSimmgcDsXxsIGs6yPyP68XHL9mZzrOWErOJ8MsGd/tZJ
JFQoP+CdK0yPc7uKLo1Esf+hZi+D3pgq4jWuCc3b7qVX/yzzCXSnuVmQ7+7p
H777pCc7NZBU1MJC3mHDdj+hNks+s0Qcq0TEpvk824xAHm4916Us9mRcdj69
PsWgYieCzgHBJ8plkpQnT+gyb4q/nfciPJSimz8TfQISfviyHI5223o9FeDM
SvPSLmEQITR3fsfFCmhsPdXh+3DpD9Gpm0xETEfBCbFIx4IBU/7oI0ngm3cl
5J80AvKZC/FGJKcQ5Vawv7Av7A7ZHb2CWJxSR1CSsoV75zHVSBkRE94QCSRf
5NCYMmlCl4oU1PpVWidfGxepTc+F8ZkN9rf+XTQk+89o9Ln5+6bkx0V4X9WM
RKj2EWfILnjhEM8w15cwXSN0A/Nf8YnTcKpKRwj7+rg1iKZqUKFh5ASgYlI2
5eAUc6OhaS953qp1/yf27C17qm1WFqLplPvUPBiMMizdyqIkrVlpcicU0HUa
OnsEU3h+NSFP3XnJ4cP925fVgkBPxL0WxJLYKg1+kimLOteMVFK/JYf0ETUW
QO1HDL2+bsvBpzlj39aPTeia/34QSyoTeQD1U7xctmYs0I3ex+XoiqUZJPac
iaOVqcweAdfZyHdk5pB3+nbCDQoFssCJxKP+DW6GNOkZJIc+nH8SwG/sNyUe
DS0toee5lrzS+q35rDWZRL3TLF7V+aT2Bk+mB0eHcmXHVJjLQRm2Cz8wqZhG
Z/0gbmjf2oyDok1tiG20cj7wzklSWVPXuEa20TyiS16KeUfxmKqn5Zfr1fG1
sONS5+WvACTpkfyowLWUpgyPwauq2od65YvtNkwmU3O/4ZqFTH9LBmg7UpYs
qITk+NCku7e38IXVJRiR3XdH0IXicy/bhaLwVe4miBWb9BBbVru684nS2VL+
1ow2VM88k79YvQvZyKOgO7a6k4N10v8lIifQiR62pn2ykyjX6U+OtbTu9Q77
t9TOzh2vdmu9zSbKGMTxr9RKP16HRdH/5eSFdCjbf3Qco+upoiDiaMz8AFac
AAqSIKM4woK/Tr7TKN0UNBBkUbKAbzJZtJVU3b2/6plPMwKs6Z9lmiCHsSSQ
pRhAlH+XDPaxpck9LSLUj8JnI+3fauTZXrfvalQBn3DIjkYEoBcVD/QcwTvG
Wzf03wAmAF2R6+k4o9N6WX1rsypyTOze4tzo/iVXTUoOcyQffU54N2xVGjY5
xv2mF21Gw8PZSO7NV/5rKAHv1hZaHAmuTisbmjND1XZwF1gOaWVLg1QqPIWh
h+bJwBPqu4FBFSnonQ9G7m4iofPYup9XiLwTP7n7xCTSXbPmesTqQWgSXjmo
h59J/NbT3IQxKlcSRQlrrwegFnpbO/zEpZe7cV/OhsntLeKunCMvvRW2ihXx
89e+kQOQtVtcuuDzhPGEsGoTPColApz7y7Dt6JpVwA1A4iv52PxEXyGTk3MR
fpB6eS66zFsuo/JZumbDVkLyrSZAyHS0lICDoXBzZJljsc64x0TgxpJeWvWm
SAQehePEj/mBPdBBSM8VZus46ZCyGXaHHvlZl7aBn3zWJZrkUBoRfEotHK7X
DIY8Uqre0il2B0T9WvNSHQIxTNqJau4D/jMIPLk8HssZC1V++HVrnRdNKitU
DglTkNh6qi3VceJFxMJqKW/EySvyq4LJjyOPmhMZFc5bVuSL8OFazTxgQuKo
4Ymnxl7F9vD3/sfP4ObABXEaP+hvCF7RLZ29H86i8DGhK08zYlNf9CIlblB0
x2vpHkgITZberE5Xgna+2lM2EqvUHGKpeI3Hn8/Zh5cjAmTkXVIGe4EjPkV+
lKLKAO+kWxBxXT0/O3lobFmwkd1rpZpHQG8YBgCZGsdI3r78+KZkIfwrtlF+
sANCUuMiA3x/Qlz/ZxV/tdA/HYTfArKgso5/W+JmKzphBBqA7QVnNSkCi26j
XwaQKuXuJBxb33KEJ4ZzkE7DHopLyF8bsEI1VjZin7FP6h2vJaqR7Jh4lbS8
ML6sxDOyeNJLZDd5cWziFkT3Bx05kCHNhRODqtUUiqAguaG2cc9ZK7jdLgN0
XPF/wEvNRnD35vS67hFrD4C3Yy6c/VFSPxmP/tpL4HhkgCyzaRgoek9keBjq
eZBxYIShWZTdJxDy5XvQhGe2eC+aj5aa+YTAWE48qUmQ69HEjX8uAfCtgTV6
ENOcHEi7EcpRT2c8VRAZr0g95zRjKognDC8EnrjPSRAbrBvOx1wu911y1SrE
QRYonUq0N7zzW9akoLPbPAQGBWKu9V439l1VCe1nssSUj1km54VQNiYzE5gh
+jTlAp7iS6YLzSdU4wOhIZKSMxcipS/3N1gQb4ZmAyfAxy4yAJ9UC4/dBQMk
mSFtKOQJHDRlu1CLqBKk5EngrDy9mmm5hOZWyF7/G+rL2RSjjmg/bR2YLLil
AHeWEOToeMcKELhYL7CqPNDpxxqffkaMP0R/0NyJP5dv0nF8fP+HRNaZWhie
+Svt2YPjJLAz7vRA3V6yZnwiQlWUFB1HBzII1i5J2z8gCQ4E3YbZHUg6DVhJ
F3emCJfipYgQzWbLLRFXJJK1xQyubU4ZPbqNg/S2xEta6+YPXNiBV2ZYc1Ib
Wb29WCXM9H2CDZlgPGrGGhw6UCcrGCYUZYA2Hps+dI8nEMfKjFRDEjMFHIqi
Bxlk1EB6VbTTxO1CHx1s5EaYixvxUqdu4LaBPwQstSGGPvXKZt9yU00iHhLD
WjMmxD8ovAfOgs4Yj7iya1ux0s5kZrn6FW5lT/5yNw8YGfHBD78qnbxRv8wz
9t0joy3LS70ZUTttbBYOqnm/6bp3i5QzKTclTvn5uyTdE3SOgeW4G1+9KxUR
RUNGyk1QC5iZE/u0mRdFpcMjHBrpr9pC9gMIbDsI+93oT09K45NoWV5gVoKm
kzJ6zhROBfai3TwzjoGOn+vhFgaMD0NWpWwE8Wb/+WFyO/BUW3iSkK+GOCTT
Tx940e87xj6IiQCF3cMao0UW8Xi9bTgQhShk9qwft/Xpk1gBjJt4xC0hotWe
ORIpfDHYTiZ9Y3l7Bb2KxFgF3X+mtdJw7mzK2gKi5Swm8M1Kff4H12gWJ6l2
GJ3rjlaTHKgQ89omCZCOM/bmnLLxu3BgVf6VspeBdtFf87lnFFDMkClTAMd+
tULIF+3wTrAxZRwT6i+Pu6rVIJstdqd1ng65LRYL1kVa1r8kIFBxGtFjSFWE
Buyl/iQtd4+Rucs4JO9vGRGTtnt/09MVXl9QPvlDv757L+2CIl5K3YpQRuTV
DvHbYJ7MTsV0XOJITKuoWQLSeF5XFILRpVCsZ0Ia6vMaPq1UV5yJQ8m+2dxN
Hr923F/02cu8GrJ1svmsLYPDcrZHsTUTPI2Sw54iqA2ry3FFoT7VLTCBtj5z
szdss39peCKz55d0DvgVMTkFXjqWbJvSylQ=

`pragma protect end_protected
