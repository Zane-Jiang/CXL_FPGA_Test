// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
rY+hFmXNsdz+7kU2u0/sHYabi3uBIVjt5gtlnh1AAmiGEtWvDcCSe9xIrzNtF34o
ZV110DBreDa/rywE1QZALCW4YnTZwXmZlB9yZr8c1dA43PHKTr6hFGt6rNazbTY+
UzC4+3roG2x5LW9csdcYjxnjARVO6eMttfR0T8zYfhk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 14528 )
`pragma protect data_block
KbrNVWteI+CfK6F4PC8kA5HQSLZSkUjx8gUlm68rfRMEJ9YLjExV4NDkuEaO2dO9
ySOlREpFq2PBCIyRCWXtk6X3CG0kDeWZTYnTLGQ22U30OFPXwmJYvPO8ndPai1Hy
Rezz5ztZCA4/FmEhpEMDsHCTAeCYQGDW+RIDyRj1oFVlLIzrFLCpvc81o18eK2fP
adulsK/UBydwEEZVqThIvs6f9bdVUhAXVGG2boOQW+RfCc/w/fRgCcbkyHK25oVD
LionVx3ckWMNRKPRzV1V02MduWjLLt/Aml8Gh3yzm4QmjUVLcj32k0om1+GlVeBv
VY+nyTtllxCuOJJn5UOicnXP+F/mvPlS8/W4DcWK8crAjuJH2DY2j1zkpI+9REKE
2VRMDbW54xVSRvdYVW6HCpIeR+mDrha7u+VXWkAUa8GrgH3qT8xet4wtVXQHtVRK
O+2GSl9w9ZqNw1nqOZNw4esnrjv8Fye/l/azC9q6rtTPCbm4XQtamuNq01DLfG9a
g+jHUCaAJ8Vl1vGu/JYVx6u6TeEF6eP2VAVe3KUyrMAGCJ9CCNc6aHTJWNkfxSJa
4VrjxComYVdfsdXsuReDR8kg34kp+KP5K393U7w3MBAVNpsrVGgw3IwC0oOGlbXB
u3pRh69wGwxahf3ywqMghE3ns0eia5qxGt9b78DkrAlTrRit7sqq5l2BzGcjvSni
P2uOpzGxqMN1ig2ygQE1C3Qc9AtuwlXaF1ppY/BBvrwH6Z0wTK9lG2SRUnSoSQHy
u8I8P1Zabt0YTjC77PZ8mNpoQRPvInlE7hxiFvO1BBM6B3WsIQYE5f4bIPF1oDTD
eliqYpZOB+J/tab3qb5sy3v73Fms3ZBaJ8bp/roVTvxfZ+bNbeZwkzmjwNz8GdbC
2EeZq+TnsJTtixYs3Baby4mAo+DEnFt6x9aZQwEFlfEiiRVZF3NLqzfi0QEttuHr
4qa42OjYFLHImBQRD1oqmJ9Q4Kdbr/09CCPbWtn8H5+QfKWF0vZDmAaosm8wcX1V
IY6LYATAQmsLMTY2py7IdifWzdrX1oIyasiYLG2O3w+1STiR0mpG/hFgYawMos1L
4TYZd+x258ASrc/ohHNjmKrUKceVMBygIEAA2AjmIxBGw3f1RLAl4aNlH/HZurjZ
fLJ/GT4iXztF4dlb0eivCt8NqqKVdQvckL4ugTFZWgdrKjI7ZpnDBCwGEZyuvBsl
fRAqoaWmsIfK269VuMdo7R9j/kP60jnUqXoBJ9WX4MBPJ3l9GM8tv1qaa3EUKVh/
aygnNyPm8TVfeur6PBoBYcNGDf4FACiFm/JFRaihkhB2igCmvRkV/LKIhIFKrq+b
iCmMpEzwZgTu2jziGL1M5KJ9+e35Xi/h3XPmNbyMQhynruoZCQnCRAk8Waee6k8a
nSyfpThjlHfPvqJjcyWlJBVkf1k36Wnhdlygvv2x5A+3N7AMKaVLP2PrzYHkW5AA
6taLSSFJ+PDDVFRHvgFkMIAy10NozxWtlNA9rNufp2XURCltt/y8T8ymDLlD4meF
nTMVoMyebpS9gOphFGOh1d4JIlmGa/ipx2O3KwBzJKgri6EzkRK49Enn6+C6JcZP
1yzePZEF+1MsZ47m9M0LmUodRjyuKBHOc6nh0/ZIxmcmDastOrKyAMdt/3ThTaGN
jqxgy2Rd7DhObPNW40pEGVcyE6c/W6G0Cgc/PrWiF61vlE0LRX/YaUjeTfE8iVPq
G1lC1PUaffF3s87Lkw4RO+1iW5QzEDjUnD0Tfpro4q4r/XC58bWq3uvpoe3IF8jQ
VIiAeLJy0kJFvwyM2av3quuPn6PkuE8bDKzdB7py6ZpexzmZ6bTwRdIFod17DvGX
+kPIK6S4LHQ9BKDjgaebTMYUwzPdbsLHjuHWF5/jZOTaeByMwfQ6SUmBz71f7kPj
4co1Uk2DbzR6DBlukKj2aVuMMZy02KSbb69cW0+fxG8i7s4X1b5B5y4BmGMVCxGH
cFsgNn4w2zmm8BaPqJ20ujwjXdVSEK4NDf72EoxdV+CquQtIZ8W6yZOp4ambWA+M
ZixCIWRJcEcwm5KJEAMj3cugQPreIpr3Xbyw2pcu/POzwBciiCK2+BeBgBWCdP9y
UcV5XWK0cXLIeCpPqQEc0N3ye1U6w/91oUn2iEr5EIJ6TfYPQKf0feE2cisEo/df
MrF5ibEt2NPsuscq4VTjN9P8SP5ku08GHY4HO8I3hkLcVztDktLQy5lAVDc5QWgo
H/89OwKXuhrzH1dyYjwPW6+DRaJ4bD4/Idt/RS+t1NwZUKI9qmRUMmamMyw80oIi
4dYia2r/VgLYLb6nNo6c7dhzNaRIisMz4gWcMjAVPhlLxGBkVDIqr97TtYPJT1CC
FcjBNQzqDy69mo2Cqy4WIJKjlypvrPot3kAsEc0guIUgIjWJs2Uv6nLe1JcasU01
ORaJEAyGcem3QUwjxNX9U6Dq8emXHjqkWhGm4dBq0+yQCrs+cYqmUlxSPa5Pdh3A
xa+qC/pEnJUAtjl1Z6w+ktdT0EQw/ox7cZzq89qm+Ombb0SYUkhIJt/pWZYWKr8h
cxIwb5uqScmDRsFpBiYfA/hx3NALhfNs9zsS3h/3tyga4RqRjCMX4wQggF3HLynl
bNWe2d+N/oOpVR5789mLQRbUWJmx6cl/ZyaCub6pOFQi8jwZ572fODNJmz4pe+UE
vtHrzThdVqlW3pB2TNMJbCRyvdyrEOIlmgkFk+EOCSE10CBhxuInYDjqFQWY38rb
ajeorfH514jLjL3LjxYH0h4eJ6DUXazi4Sg2FigyZkdBvSlpA1qduL20mj+LeTV7
4xKH6Go+C+iKFjayQ9g5ma/RHAEIAFNA9YIHMIA5dYg8yGC8LycmufwJap7NNWun
bZbtI7LZzTJgjKCTZ0B+yb3kcnB2XuLcjrXY8aRNSKsVMn/iVj1XuZiq934EWVJ2
q4fWhup579YKzt60LJ1sZWztIHSAog/778G+JGcha3ISEHGnMGvJhbexJvkpSabm
RCt4Lig5Cg72hFMuC+1qtOtOE3Ngtqqnk+m37igu0+VUJeWgMuAEYru92f4z1u/t
wszKmCoZZIRYrZ9qsGNdc68qkseXoo085usvyp2Vo35PZkqXxufREAVgQCuZdlfM
rWHgHLd3MrQzDXIlImah39Uk2NNLrKX8K8FnMIRm4yfAZtQK0EV3jB/9j8NKqOS6
8bj/FHm6wgttzI8QMUVmWnhXMcyXPbnANek9IHxJHAXvpReBY5nx9d241IBpkxMx
Ubt2tx8XHoxQANOMGR3s8h0VWEPsZO3Qm4/+boVq8KCLe9uisJJ7C1aKE3yO2RF7
NmmJqy75lz8NkJ4cK1BilyoKq68DUsoyyyQJMqgGemAmC0Bg8XD7Nv4DPRUXqKBB
lRENRDUEpn8gWN1V/+rk0fH5WoaO/FVOFo9YcuK7MnxJYCLsKHD3rBRNmlWnc4OE
3ilnmDsTuW51p0Kb5riaKsyyMn0vNu6hkNDg8UjiIxrzVOu4UZmgfHLp7nZg1h82
kwG4rkHijGqdZetp5YUayCRnhp24yKZXZw3Rx74lXJIK8/SKuuxIUOnixIbx4p6r
V0m8Z3kexWMcQ9ro6XWGQF7HLm/vCydSyEgf+SBIBLe69rrs0PV1i2iIHpz1ETZ3
L7zuDCqRJb+Xzp60wPTtOjuvxOF8fxNeuwipzJG9xguu1BtDgjT7f0Yhh8UsZZac
Q9ipF2EJ8rzCk6myWId1xZPOsjjISOqH0fPHOMouVTZOiU/K0kgf21XZh8lWwhxI
sH+i2kcx/zsFx9LaAPIlVq+zaR1uIAWN34cADUmZIqX6wbYScnC6g2JgPQP08Us4
/qMF6ML3xj7THRIA+QVf+byJB6PBWsvd9/l47NAm3GkcCxG0Km5c9CcattNs4QGD
26v8hDfdcUEGnDCxo4wbvoDEo1/5j4UFP2cpoOW1Y9xMKZvMtE2VFDs+WEQqB6NK
Lv/HwMwv3N9s6wfVZdnU6fLX1dCGgcSXFjBCaYD6nBp1hhXicYkG4Q4lWhDxPpj3
Ewp2Kg7+KPnxxdJOCBfiByuggZG349ky5jkifF46Bbd51/oar8BX4wIKvphqET3x
untsM7mVQmGSSEAd7HvJx93vzPQkztmKKHLWnrY83IP6FV9aB7XyveNljsSXOdYZ
ItmDcrU7v3bJEFAP3wi6zxxKenca54hhvgCEycpO6yE/QHm3Bj8Oh3ViMlXE7rSX
fktt6ToOaail+Ib+vLMyjCn8oTVRPX7k+ZIyDUSqlzzaBd5bsIUVXhMmHXjj/cma
ws8iziAKUzVu7Gv/VeYmz3atAoFwhjfrpzUG/wUBBvmG5Jrvd1HIdDq11b+Yz2CL
KKetFnaivfp5ev2dOXIjQF2ouHy0kwgVNNJW3uu6oVBpXqHCzIlEgO/JFv94V238
cF7kDjDxHRyLTxeVQ4gkSnR8bPedwENvDni6/Izec3Qihavu/0/8fqzGs4etoSDP
y8L+DEWioaEgkZI+TE1uaO+AqQyyzkmm2g1et2spl1EZ0g1EJjZwtzcTpOxmFyzf
586x2Bhs8LxygFbY/OtPSvwcJR5plaXW7mnY7biOvAGW5gIZXrHa9rxKWG7xFMhe
xjT1twjpMZfcvjy4Hjpjc3/d22ip4KRdDlkRYBeS7DwrBt9aJpaAmVqrHhtzvqpi
cj+l20/RycA6/dQu1AXYjpDdaLcMTDnZDegbxPngBldmUNxM49aDeobcZVgmpCbp
0McBt1lWwS89XkkgPcZI+IobeUr80sHcTbFexSN/CpVFYJQHhh4IRIn9HB8++Ich
24Gv8s5TI0wsq24YYhkXvGwyLbOiLayks3wjrCy2oRFS1x8zTWpHPFEc/OCVL5Yk
+KhhoDfYtWXIPaFBZwxZ5isCCuBZkJ3CRYy4moCSoQq+320OeSGTqKeFSFXRJQ3V
H9O+ZmbFUaK5AOpe+KMKGhi/mG6rldFZ4/wIvwr85T+TJC81QXmOdpDpAcZjoVIf
xdmuJX0+kWRgir8xl50t0KCFi9Cc5HVvFtxZvclIgP0SkoY84Gduo8Jc4WZn8mWZ
BFYTnJ0nwhXQs+rAqrIVqJxIL4CtlxXzsC/IxMiLCEWAbTBjAfI0RD8T34AuBh4s
ExYtm2rlKgSrUn6+2w1n0H27f9g/P7D6dkt5vnaIwbnQe+LzXRrvz52oxmH7IqQJ
rukIiQqzwwNkjnyFQkK2B24ZSLLRQZLCRrKT4GqGJJ7Nscqx82QzPiDk6mubvbd5
SdZIqwjIaLMMcspitur+WtiL1CRSMJiQ41NYvvBtLxxsKPt3LSWE294X6JCBTjC7
Q/rnQ2L8puXV+LhqE9xLJgZO4ASIoVzt8GDyMmOvxwndDiBIkcl2CX87msFWFj+/
+k27x4WiVc3lF6kg52SHi1T6OK2HoBDYs3lrxKJblgBoHMEJRCR9HYyaw8RWL8VP
jvMcJebMujUHY0wRaBKioRraYXOuZ46eedGkJO1tVyIHQfUBy1QR0oH/498kVi1q
IUCXMccgXlWVyYMuZLGp5K9yGIHemLlxIt+ckVf9SZdrYfvZuCqXlyZUh+QzLfx9
vB9kIRaXE1h5r9rimZeZmxTzDqQ5Izilu9VseGJrhySjAmAbI+OclkfMoxvOesbD
h7LEyg9OL7JtSAhWUoZQX6OnASAcF9ICrDF2SaWGitiDzjhnnMfKKXkP1Z2dufd+
nNY2wOrjFRtyBSn/NJtegUBrPEgQiIEZgfeUlBdkbfNoET2wT1WVmX1MgFDHulcN
esE1A5+jBwdw14JhPZAIhli+6G97g/8da1Bq/HMp3SjMlShKjsf9s+c0BoBHCU62
E274BDfyRMZ1m5lGtZ/dpjO+tTwHap7CWRRFs//BzSZcJb9pA+GJ/apYxb7GIflj
vFzM9iam4IluDCSYTlJIlbHCfYshx+0azzfUDBEzgErwZzTaFx/g6xduWGjmpfcC
xcpedCOPUpHE83nfNF7UuKDAkRpAPprd/4XENhWAxhteNBkVih4yQ9FsaPXYIQB7
X8x/xS91CoGeG2nztJg9tntiWEglgqva7hacleEQa2lSmZ5wKFYEeY9Ya6mUiVky
XEpbimCF79AniTqwayqAflEpECP85l0PIrO/MyGH6n9FNTzmANbV/bPFM5n5g997
P63uQuDQ6texmsqZyYIy8NVE2f1Glp4s//yp4MHDDV8/KXqUnWLhgJtoUQTYgVt+
AxOUjF9jK5Bss/3KhbQA7AVEYsI+cTIWhbVX9NhpMOBblNVnfFDCX/fwaUfGd1Sc
1oskcR7GdYjXii7YlpKVxmXJ/eEGQ7ZcPiEXzBYbFpJPlXTu6TF367/j5VawWFtA
a3DjQG4s+EAJpIZwrEwFTls0TbGkfgsYIjpJdT5gJbZ5x6QZXEYlHq7UvC97a6Ki
if8GII1ShpUQpZBdyYbC6gy5Osq+h7PuEoxdkV2SulE7wY4uL6BuZ2s8jVK7YxjB
E0EAkt1vjenJ2HEor9nUXJiL3KqFoFQfqCZ2yoyy79sGO91XhCZTJFn7q7cRgnsH
iSAygnD+CsOo69oqbK8XcTLVFUNr2eRicya+5QJeRrHJb0loflM+7768U5pXqKnu
8wxYXCUaUi+OnuC+fO96FEpLtF/7feLozZBw1e/mgTSoNXDc7/xNZnejOyz+96VH
VGot8d/vlCJwzZl7z4wQ7A7OkIMpnL9htWJhdWYf0q5/8LsGdH4e9QSUbbwWrWoQ
pmDpxBDcF6T2j9DfUsYa9+iVoGe3t6ixsjn/0ZzXousmdCY+11HvfBstV+1hdFYp
y+ipOPvgNBDIpSND5JVMnPq2fm/4iZ/SQX97U49NGe0FHzzE/GVuyemVxs6HkvFw
8qN7VR7taPSvOZhXrl6RyCHFFjvi+Elq7wUofHxCuClzb0FUSyXniV98hQ840YPq
ORBR0Qu2Lxb0INUdLnBmVJZL/I1G/4Wr8THS1YA3DvDgnqpus5q0F58mnUJU/FrK
Bx6rdik0jIfzyGlAY+QCrdHD48djux8R6ASCadC9O9fw2cQtuor200IkIrZ5m3pk
L9G8CllBTnjVzYD2R4flecYB59NGWQpKQsWrPgrKQ4PvtaCKwmvUjVAnhQwiU4JN
5+Tyun81aYcHKU+fv7oCSF4htCJo8Mj+ZryvCGfXNWOqkHskP1EvUwztcrAOoPMi
SoMO0lrGXhJuemS7HJYvCzxFGo3j7lK64y5wiCHhED1ftGY36bPnQjZQREG9MMKC
ua4grqqIU9hyQQDL1YX/CnSL61EmIWdvoyAmK8N07/ZlLqBkdrX1KeteU8WvVEsx
W8jwHJvYegkHdCBIOX7E62L3TvJ0hr8ZhTF6Xfp6im0nmcpI/XZ7fljigYM+cvx3
k+dtGXueaZp6UWOQINVnjc6vK5Sgiru9/xgHvV8M+SCyetoI+S+MBcELoBkkOS/O
vLz+oBQ2VF10D3JbMtUE7Cxtfy5QHlet0oYmioZywcsGWqG8i/qBR0QP04qfonis
mEjSdLN4IoyWeU1eL5jDk1hr9a8nn3ga2VgqgOfc8517dTwEm2o/RZj8u07NzVXM
HkkE7SxTHfREpczQIjUOTkK1ewkdEjHTL3kZLJ6K8vlKiRsvIpjQpi2YgAOyixte
4IaFJY/FFFS0yHiSoLziy863pX2N94ByU/RkTUIQ6+gVu0ek46YVh6dqLeW9ijDB
ZWWeHj9Y6us2+2KIQ03k+KxNjLsU42Rpwf1eAgmgsOau6u4gbJQYp2MrPzMDC/EI
i53vWJsB73G1JNZA8mPzSIGOmBmLoulhDkx9h9IlfiZvLLlybkhipJvg/ek1F5iD
eq0nV5hb6GmQNpJiKTUj9QsDbQZrlM6fRt6oh10wbyMgBoL7nJ/mTxGH/XL7Z8yt
7ryUOP8iu7gbxoqYE4mBo9L4OjTqUqKDZRkTqSVf9vMYiw2dfJQJG3y8AniDtGpZ
zO9VVrtFHidi8bBvYiOtko2NR/6ajOkJCAH3/LUWXOdpCw56SJtDmymQzR4ylbOz
mk+TSUP0qHCdceDa/HvjQSmwVLs9q0qzrFBxq99ktPCMjWU0nXYFs2O5tX465NFg
+SoSWZRSdgDTyrFKTjKzOp0U8CQLPNxsvVQvKvkIYl/ZtW7BjjfhF1u7pOxOCQ0p
AC+WCx141WbgHEwswNqJoa7zpM7FKHoQbTTC6xytgY1F1oUXeDR3ljZXNtKnxoGb
x4S00WTPwHFPqDKa4hNuLfc3B4KTKIUVbKxnQrbNDao9Cebt9X4aDuzFUmJuidTy
MfJhDqDBf+ySF7d+Q18+8088QAEsRWUqyiD74laCxFFMhU/Yu1dhR6k5HSRF/Ns+
PAXXrrG/ePHHWlskFaHR90E8lLOm2DZEthmGL5XRsOfBuk3RcNAI6NgMvIo0OlZB
Yah8b9d3+3IczqGhEqELw8CWtLyE9GRqpA4FJDB0mwIm1JcA2MSbclSmyBTKTf4k
3Z9ynHsWZsk400UFa74Q6jjESLhITPeE9hpPXc9AHV3wSd8b1i07n+uSF8TZ//m9
NBJ/dfUUKcBDyQpOeJN/IeX1LtqV8NXLuhvbugaVQO7sKx2hR8nWL36H2EG1fbL3
QrpychdBDtMIMtJpu0yAMuVnw/5+A2uQFSVWBHI9WaTQ7nD360CsEDQzhkoMCFMx
4Nq5bgjIXBHufNG9IhnAfKr9R4Io4M0sxKtBZ7xjmrksVFlpqpO4frzFfdClzHPl
rLEeyWcY1GZiQX1JYA6C+y5yM2Zr90tFsNcjCN8mCqpNaLYzYB9KUEwSpUm35oLc
pTOb2RT4P3jyX0rlNdhw/+DyZBZOA+kf/KHPUyFmn6S64TtyEUDQia1YHFoY/sAR
Yb2SaRmXOkss7RQ6bxoRTnLWWCR+d9z6Kgdmc7cd/3H621fd9a3WNkBPfWXRjp9v
Bq7BUxqpSISrqSy5UbmKd73SSAer9BG+lhlX7pgX9zrmCi+n4Wtiq7tSVHfS5ueJ
rlDOnhPkMmm3GB2QDLJz0Pu2LvCgi75tZLFOf2l+2AdZffQdejOnwHNCb2UdlRxb
CQ69d+p5rOKvEGTnEz/D3E33aI+Kr+377ISQYjLBg/PlKpZGGnFij+UphLu2FTGp
VyR8JBS4uyboT9ZskYQ2cv10oa/oduOxnl8W+avaSkCxgwT4od5PZdaQFEW9BcY9
CO1RO1iyEaaSt1POK0YrSjydMb1EFQ11BNpsrU+dsnZgfjPAqW8uUq1FtXyh28Mm
Lpzedti2FWlBmAqdROSTeupinS4iLFQt4gEWBFBCIRXrzKr/QRgef1J5Q957+G0T
H69o7YxEqWjfEuKYligjvK0FEyKrgGdSA88JEacae99HNWlArU7lq/OGFvggQQgM
DPouQvVlIzf/2LO1tKUbWLhxC6q9r9rae8kuJD/dGq6VMaauqr8j73AL3sCQgodZ
Hk1aOlh21ikdm9Pa3/WL/dZBcqglsaHgBx/TlrbBm82IYr1RHLN8WteDmb7DpFCn
BDTNNugabBTJHEMFlMoLceYA+dqbIEE7GsbocoPI3qgO2anqGW4Aed1MF6L6xYLh
LPlFDOWfEiW0Nf/7aFM6DDzq75wLpSQQZI6dDh3gH0Ui441TMT8BnH3RQKq80moA
BFUr6h4Buv9THZ6JnVgnr0mNU2+iyJW7MoT+LojHWau5e9foQPf3ziNor8wQA2yw
iWqyQC0gV4KokW+epXIyi58LoIyQmgVL1fkSO1uvHy3+bHb4LKMA2PS9xuqYzzpY
y8o5xVtO/u6KMooNcHlbq+YMnCm0yJ/eV7NifOvTduKFXOv0aG/3TgiQUojMtz5q
vioasSorKcOOA8VAs3zSQP1qXFj/sLs5pdUznF+BPKjCAk9vdKwOZVfwKHRrE7Yi
1wgaIOkOlX5X7oQ7gcjaS5/s7NRjpa7tG5rvrdjOPLh0iIyAd3FxNttbkNL4/yZy
8aNhRZsnHQVRzNPthWyqZbsRumCm+JcDUxPrvhOb3BJG/QEOMh582DIFYw/Ku4Ew
vUDUfVQvAjBNpGoz6E6acJcW4+CiY6f4TFDyGYkHDA7WLkru3kJAdAUa5zh36MuP
dLIg97CUe0QP23+Tu3N6iqQcVerxRnVc7rRxL3VsozTDbYWJMk0OxdjrljhIpZfq
T7IvY17dRAdNLI9LlkKVVUZ48QczmNBqmQAlYQdb5O0axiIxW0S9xaf9jiwvf/Ax
CSMmHLWXZnShRwnDZOEd9o16BDliENQtzyFGaNLty4f9xF8saPXXnYZfC1t9cD9c
ho26Rx/W20cNVKk5yqne6ImaRurJwcnRIYXIj/A0RaDlsrEc/Ef2x2KV7pT2L3Fa
8Uyl9rsUAnHEG8urer6pgKNLf0wRQ4HycSjFk4hbBOOFsbHq4aqCushfNxmR3Vjg
xBvlXdKGYNOJd5NRDQSyIBXKdek3Um/L264ejliRJ5h3IdseASamzmFUF3yGVqud
h4DDi5b3BDJeZ7Fn9wENPUYRoh7zGbOgP+JEQSTeNtjpOPlmzehO+ilG9vb+gnJA
0hR9TJATNA6+HLnyqTozyGvf0HgviRmszMpGmwhRH8505Sb3wsisEU+ACoDJgaAn
KEz4WvJNgl726sybFxVtkVyNLUbbNsKbSY4sJ1s0B29483JWgLM7d7LXEP3ftqkC
5c4BnwoKiA8fnheljqyRDWzfFOTZEyPta70HjCKWoThdF9JKC0S9Cs1FvFs3Nq60
/ly99bW+M6wCJwxSWfzZTC4LZSe0MJoP1DUKGFLVe5v2JRu5VZNXHwwXmi8+6wyh
mtWKPEBckG+o4PBePu7aEYry8ZOvVK88K2GW42h9HZZXapxUtX5cHgvg2TkmarOZ
XD/KScJe5DEteJkMG5VRA4wFNOhqwblc0JeY8SCZw4CDmUOY9DJs2ZaD2VX2lUOt
uR1K1Mvv8/ZhcDP3RE0LwKNgYLGH7RurAfuLcIy6XeP8dsGCy4J2KJbTEl7pyt9E
Jq1EAz+K9L71q0ZSggD1mXOr3UJqUq2fxfcmoO4KExii8r82wKq87YchE/5+BUdH
aEUv4ADaeUIcCPonWwuFOc6js8oaY3qSRVpQdU2KVUtBTGX24eXJwu//JCt3uDhf
3DpNyrsBAEETRfIKsYfA2DEgTCg6yyJ+HnhdAiJuI+8uhHmNRp3gYm3LPxP1QvXT
x52I35GfzW59+zvWQbYHU5ROWw7B+JQuRM3WuZy9it6OuJkEBboAVLHgzuS4LWMq
hFtoza1EGls2/aCd92PbDa9NgLaakOLuXo911I0PnK3yvOTMJBFsA6QKsYkykmYN
3Sj7wW8SxprC66ulee0D+ZPVljfE5Y5tYtGX5reIHENqkU+Lw83sW9wV6gB79KyZ
2l5lyTl6OIlRajup3k9qu0b+QVdHILYvLERGCRlHtMuJDNN85h1B8/du/M0s8Mn2
FSxYa727b1qgJOeC2JGqL4rlcHtZg0sj4DU2r7xnZPTp5D0wyc9exlnTM2Zkzpyu
4WHu3Fup2QiG2dMjI7Gp/LEYTJQ3AGK8MHyrBmL9EyNAQiYVvViglxGZtJGE0P31
Q7rJcgS38U0SqPFDMMbJWYUft8Lrz4q0nfuDOxd079oW7OLpi3vacwGac9kgt4Uv
M53goQNXxRquJx7xLSpFXv+e7+PO088MFhghr+WzEZSPS0QpaSpLCvRQz7kw9TT+
6Ghl86lnmcw3jWrXSDYyvLzEz3Cse+b4Uh1+OwORFF/Pn2Q7H5oeJha6bVjXPx0H
Nzih3sQdsv3crDYijDjSYtjTihSxCyuwR5hsWZqemEnxgKV8V0ouEy5IJsqaX30R
mGAlkL/eeDgqBnqAUdFmuOuCwmE/3Fn/KiWfnPFWj/+k1F7t4oRuSddZqpskV5u+
AinRO/HJOWY/q5IzVrp1YJQG4t2CF7USFz5dUU34ixZoBe82fsZMtddKNq8Ynp+A
tmwyslamGyQ4AQKACwuLuJUmAO/egpslG6S7+ajqd3uY0gxWQbzYROadr0RSXMrm
kejtN7l21KUIoqmSZIaBwGqHDnDvNdBN9ztujQMozz7iu6s/M26ZFPMPh5lLw+r1
ARDqYVOTSzwmb8BRKZTPfVvzHuSscasKxK/exqYnFYOK4uABpFaawWMxxriM9CrJ
GGXDP2d/no/7Wz7GFRpmz1rS/9Udo0ALkohsFLxna7NzA5lAxVjcvVgm6NxPAgz8
KczvXDDB5wQZQO7msoRThS8BiZdTf31RcUxnpLdpXy0QzxS9fslXH4YkiNBDruFN
5ZB319TtPfhDm/EDkWrUIa3xAuRtr6KzUbjXbzweAiVfzxqGab8oiuKuUkzvUQrH
0CZg9rmcxxkk1DCl935DfOuxTF/hnUz6SQudiJHsWfKN4MAFeZcwlGgNAfYghQ3+
RaDPKTQpxtRPJnXeIyShclG/jLqpnDmm0Jtq4vqRDdyoqUeaRRtTa0maQUdhjagP
xkI8YeiV/YeingwbagDUFJoGGf3zQ1gL9Hpg69JX+EoKDlz5d9dj5yfBKmGvdbEP
A4rewsYMyCtcxGstDP+KISe2GpK/5HgSZt04HgCw9eQMKollQ+07HJuBYDE+XApQ
XXdcAfGnjQTNhp3qirXhjR2PHF+hyEK6RLhDWkTy46Q0Czf0NELk6WQipKpsj9ai
akdSO1xxzIXnsfCQ4lPJgEhakDK4FBJ38Ey3dHgIkCrdhb00bMeKAURf5OHZMO3d
EFpdLscKY7otc2hPKtQT1bxcf9QO36d9n5thf/CeIke4SP8Bq63cRrlfCd+d15hJ
IVhd+89mK0GXyhfW7j0nHxtttIcVMQAF521Lwg3dQkieS7k8FeBbVsPqIKW3LZcQ
U6B0Qe5Jd7MEnxvqF1JVE06xadPjofqQ/RNukC4N2V7JwA4GKP9y7cu30CCvTUTt
jfL9ZUoH2F774Dn7PO6ZjTwf69jH9UgX9dSwooXH9W2U0gch8RUFt8hFYAvZSZJX
i3OA3cMAIZvAMJCb9vT0/YlDESDdWa/58cuQV+/vc1UpZAs0K9qd6uilt9sl/USK
xNE63dKCI1Hxu1pm1xgfUPHnNYPUXNIO6vkUHWSTF9lXG6Yt4N9p9LWDWDnjwJ/H
2VBz81ODhw6bMlLu4z8kjduLq5wdTUA3JE1WxbZ3pn/0iy4BvDlzKW3KYEYoLLZ2
R8DHI/Aj4Lsyam3o/63C9oXJmpegbtKMfZJGa7teQAE5eLKooYniMWECLYBtDd60
3OgW1o7KpdVbqrVNOlUM5WpAie8HIiHMAe/0EcyqUQekcvfbqq2zl+Rs08eGR+VX
TCl63JL3jQxlzu4WF4zTKvguiyfPX0yX9OpxFFEw1f2o9JGGwOQe0cSBcPiwmg5P
lmhrAhzsAG2JxGBgWmWZ58KhUnfwhocE5gWbppzVRm4NRNm9mMhunkPVKCb2Cn64
afArBm7dkDaamVYDWR8JdKuFucaRI4LcfiKUPhxt9dEQvZPDt5aUO0CkXYVMgHIE
oB6bdAKVMBXwj7gNujehyWfCxRnh0TQt3QYaXbULc7qdwor90DM2P9dRVLbTT9FF
pbAYS6dAlCuypaO4DtIvGauEd9OqZQNnOARfrur1Lz0NLH79te3t9fC4lwIPAbin
s4egmeGjHg2iA6xyz3cPIiVe87FhP3vp1AI0cl4E/LNNN+pky94X+qcpHNiB74Ez
YDEDVmdw+epT7I16ddVmCsuMslgEM1HvsReg72ySvCzh3KeuRMkvsJdDS4NedYKx
jVvdRaoSUz2pjsQl3QFcT+6Wwz7u2AFl3ONPVQFZkwRgxLV+ylYCxrv325BWAG6x
Vucmr761HzJJ5qjsr07nPOqRShn4cfKn1xkjMnS3k6zlzJ1QLsYwVDUqNFqnIqvk
mWnPa9VQ3qpsC6RlPSCFG4ZOwAMOjlAZkV8DOBhTLLE4+3OhXWwMQnpoprQZMQ3/
vR76uUNNXuy9VpGgoPohgc23bNZdLPyFnQdFE1QLsEDE9E3P1QPtU2ZOBvY+TdWO
qM4urN9Gc3BaOB8/FrbRdNrcux6vzjRcKlFZaXbf5tQaF0PQ3EJVfSBKc6rsUXn8
OTpLKX6AgdxZ8XT9LWMV6zjidGs4Jb5DCkGhp1O9LYhyYTWC4YWjsX755wUaNClg
O7Duarv//FFwAtRuTAVw9w65HHg+xzhi88tY4gpatR6iikWF0AFVCFC98QvGbEvH
5t6+CsSN7bzUiFcJHQJFjIhjd/rV9/oXCTpe0bX3IF+rQ+i3qDc5uDPl/cKHVIzw
2bRCSMA1PjtzjjVNaTiNLNRECWB8pTKWZWMRsR+NDZT3GdLuCQd3LN5k/Qx//4Cg
HTt0Iy1SHSpQZGuX6BXaVUe4eq/h/h7c5l24ijhOUQtvf6yNGYdpzq4saxq0rS+K
unfX9SDaYrzu+YRrQ/VTabdkq6WQhqr9U5iTblqT8Z1qWk8UqMRX0FM2wYI/bzF7
vdBBxEoTORvI9mRophcLyw4pE5+seNpcTJtbmLB1e8990rMQxuKYtM8ORCF2I1HI
UQdlTEhtUZB/yZbFSuV4snSRhCPT+p0WmsWr5x5XWnG/09TOA53dp+YDgKRuvvwT
nYOw+XIXNrywQlfsPVrzysQ+fx8HglFgtNmhNfHQtphJjPfq0ayQgQtJiuvaDyap
1SCYqBNin34xLd5Mij5EoOf6fAgNKSz4z/H7LylgOYU4mjXBxT3JBsvrDFJlQTtz
h9EgPEmfJCIxEo5d5m0gpanNBmuRMEq6siilFSQA+TPBnIEhZkb8+TAru/2A1Nvh
I3K9m9OJb1vQLOTD/2QPHk0jD+EBn/VHOpgId2XbARvX4fE6PgQV0vHwrxpAmanD
/e6T2xl+SlwUVKPtwU0YvYhYXZVAaQSUlIReIdm1H3q7ihRtlHa0r9Zv6TSpeN6o
p8G/VlZgYyOY+w6TSoplL1FuSJv55ePKkQ3pzStW85+qckceJ8WbDZFdI+R4HMjh
LBGvH5ozIZ8DmktXp6Nguv/ltvmyv4o0rYYtORU5dORUz/WsIxDn9q4ZNL080DQ7
X7XTbAWoE/CP6ORiEH0rTTomZxPXHnVxWb/sPcHy55y3f9klp83b9zRdfzNLVeLu
K8G3RWFoPVQksXre8ch98Oay8Q1BmAd7xZnnAevSziRdS1jQ/bYAWhPIEZsXECld
/0NUSkoIGmnXjkRf8DLt0Muwqi6DWXRs9T9pKgDW+iOXjDq+NGd2afRgHIjjX/Bo
jm5z1Ew1n9v6lbU+ccm0CzWJZO05kD1bYUAHxNOIR3oIvttnXUwQvP1OWJQIZs28
ZFqn2PR7lOjo/zSHDb1S8IhBxU1rFrxvfLAsqaoVEf4f9kduF9bdjHvjz4cIJ34D
iytFcNTNR/gnDZM6d6E2IAWIGpozqvIDNL7uF1fCCEewVxn12L1X3DLl0Wfh3OGL
l8VzjylqLtz5DvwPwFSR6aPz+OU3/rh8UILzV2apJyWOqThpnfN3Q8NxBpwMLziL
a90hh92icES/V8mOm65VwXy+NIhhgsq1/V4sxPqNSWv7JaTV1hWpgdjLot5vSdtH
KS8PF4pR9lE2KnPNtfwGHLEzR5KAipJ+lgsVmhqZgJInYS6wi/otxJNUX/e0fP+k
Kv9QJtf/FR0FBWVFjqz/M9HO3aIBcgCvE+5W63HD32uFhtzH26ey/1RG80tCTQps
AMJeyNN1DsT4TKLgCpU01sqUc7tu4S7WY7QXtIK1jAdSPgLfGajR//WvmBYTQK7I
+tpPBl61YQG/dtmF3wMMi+GvRKTj77vKO1XbgnI/kVO/M1UhzxYzeXqswXV7VUtt
lxioziPXm++X/yfN5s9iyrOh1P/ykaj0I/SJ0Fjy1Vtb1vx7a6+ZKbdysSPONQXa
eIWDP2UqKAHm3ziYtnY4Sa91oHjJmLJIboYXL2n6Bgv6T0SlllGsVvpFS0vQzbZH
hTmupCfvZoY6tM7Wkkd31KgRwcgPgvncwD22N1fqJvDR6Spis98VzDnBhCQMet+y
9dZgAfkaFBJt8FJFUCyhMSVtZ+GTn6zBGmFIAVYZiX9RxCM2P3OmN3T1s05oPNs0
KCqECtalaqNfdWYacUheN3AWaaGjDsEivk/9BBcyfIDJHjskO8O9oI/gs2w38Ng1
rhjeo75TOXqhb1rmK/Fm8npm4a2ynCn9qa4wnx9iYzoFFWwhf2btddU8UK7MHWp3
XOhzZPNUnzZ9YA2oiPVxt7vDZ0jMTnyNZ+FSL0WrO88un32V17uyFmDQLpk9SH3+
MazrtNxz/xvffm5wS9I03F6t1oV2RzyGMlUR3qAkeSZ3n90Y2oGkRUoe4MRt/ALY
wL85dOSPskqrHdwnupfFnbYCq5XxVGe2W+gSp5+npZnbXv8kYH4/rYO0DGLlzTEx
LcErP5GSd9INYZMN1iqZ8EbjIvWTZbr4cZ8+VKKHkBr3nBCIqXWB9Jqr1rQuY8X2
h/06hqFW+dgUXD3veeAuZqCzozJ/2gi+tb8oGbB383r5447sM9IxZasL7NT/O7Lx
yCx4I7dTQceiXCJkn3V7utpOPcpR4yNvFLOYcBzId7C4LaSYbWTr29SdH2rKch/i
krEErjDjf6JZ34xPzI+3fzdnuhamtEJZF8ywA/AgonwEz12yn0h6JwbRkFFOsDeO
pRLarRYqB+wstsyzdL6G0C2xt2fp5mnxPM4NeemoG1R06NWH3efHAXyzQeVjwVK+
hrN8uAt+UjgEWhZEL6NhL+BtUG5Cog8CeQWre7pbkZDG7/628pYYxzMTwEp63LFo
Yag4sTgkCYzRIr2tMvR6WpsPNnx26OsClIAra+Z2HtiGM1DuiGais7hkesSjtdS8
FKvfYlKgaRq+bZMLxVMniixlkamiLe3w/3GKqZrCblb4r5FhUj336riYJP7JZRV2
wQdTbYK7JGxOUEHChScYecTyKLJmDilToN34B6hVM4Cw6HiVGAm2oFqfHiXjzbJv
papJE3U09abR7Uz+hgZyM2mHpyZ37xh5z7eH2d3NHYn8d6Y5/cDQBe9UiK3xcfn5
IuU6w6Yy1p/qq0nhZeMy+4LAhsGm2c1Flm6GHDUuPSNfMCaV9fndtdhE7G1Ftzu1
9/bklzvzV0M7yF5H1kkCp3ZifgU6nz3BKgiOdymK8Q3HOTwTxZklm6jj5+8dgSjV
gqCUyZZHVY1WetYZYuUAXMnH0P738X9COEN8J9Y7bGvPTM6MA3Sx3XFhhBGyPfij
wHmLS0wE0rKWXNH+rVfOFYB6IEslXww+qnaVCv3b5q8M5rRHifg6cE6rziHjCHqS
RdJSF+ZXy77l2iU08NyuDzuF+HtgGwW4D8aveUgIfctWMcZCzz5hVZPwWM7v8sBa
93HzYhhzxWqA43wyHCkUaaVjkXE0xUa2Xw9mF4frZzhhOyR30pkisEj2UCOJCXDj
MfCvhntRG7Iw67pF/g0dvnj//yo+ve0EfboUXe6MhGNSDpmyt9GJVbyfWHHumYlb
k+98cOSRZqK/gJsPEGOQ/yFpyKElfLQJ5pL8ydB3nndyPBi+V6s4oN8Fh6R5mypM
bgAbZHhIVJJOekepuYjBi8gIYj01mu9qytl/vFWl4tUU5pzvXOcyuWCgOQO1xAfG
tMKvmFWmw2jHlbeCwvBEc2EhoF9EmXglyzp8UEBNyMzOQZDqHnMBBV6TIINRjw24
ur3TlNc9kmzUTaJBjR7lQvAC0BLNIGzDNzs2gBzneXm9hojDtb7toDX2Ie45ND+z
h7cnXINmQV3A4ZE00l26bPPLqRYOvE2bi1YU7Ra0Z8IaKKgvbCqUL6kCQRhRM0sq
sL1137v2JZiWGdbdfVYX40o+IKtoTJAqonWdijiyFlWodv+Q6I/Zz1KgkqdFTvdd
amUeJgh8Y6ktzC8TwuLHoxqfcJxbw5PXNcnmW2k1DmdZxvbjibvIgd6jFfRR4JBd
BXtrHrpkw2Ln2JAME7zadwgNimYlVBW8tlVEuq2a/rK1SH3tMEjl+5AcIiu6nloF
pjxD/sm95RamMoHbX+fskTb3ZwbcoCs4e+Fdy5MRxhHu0w6FWH9dhxvt6Da4fzbb
lWA1hGR6Bw0bCpJWyt51g8HbCHvX5CfP4BOFjeGgGb4QQruIziyaUjVgMEHhHRjg
lfrEOcN2n5BVuhTJ6HWervFUy0BVpHh0/v1uWZSFNTJ392U40zZKWefQUHrkQrRp
hQOliDocJnFlY+y77asnB4K4s+/2GJ+8IUk25sLjRtIk8h/VkxXUieBYc8bXhDzC
vImxMYJrsNsT9IglnyVxmROve16YjCW+5qXZEwIoP1O7PNZTtiheh4fX325Ip75U
O7BSmPVV4mN2M+mEEDrV63F+wfA+oLnOBVatfKX/dB2GOdmA5Q38ljLX4R1SWtjn
VchEJ5K6kvozz/AIZv9ox/ToJpVBDk5m4Xy4AMxlVbuA6c20gJsQ6/NJOBXt3+X3
XkOUWPcWPgRHUgEyz0D+7W6PnHyHk1L1Yum9mYHWaT/VtYA2J73KGIOGGlr3sP+P
bh34V3gkDkkGn9yXrLWwftRq6cta6vVb+O8+C41Ms5fK+8xVqAALTX9z2EjI9bdc
7J726+5PD3LpR061JInjQiM7vRQrsB+2lBsxOoIS2XNm9DrN+A9Z5wDlI07rTAPK
opRLJ12dWBLn9dAf08BAIQfPh5qhCG+En0k8H1VbFKfdH+cNhBqCQcjqlfLEYaCA
tfu0iotCmPtcWThk1yquDzPP8VnpL5CHbcFjMwXzxbrP9dPkKcCjMcwfG1CpPcjA
QuVxE4gaC3+EcUVGb/JIyP8FUm67wTo3PA5xykPdYhsnfw7jb+m5FyaeAV3e9SPV
JA1bxDlvgQ1CFig/EkyQ0MTqNkVfGd13+4BgPMAPVPb/BgCNCm0t9ldPr1kyKWsN
DgP5hBlQBwFtYwlZOEVr275Cgnczz/e2/z/91cQ6mD6TiAL6ryOoCA7JzzniWFkn
e33bgjy260SkiyWJbSy6mhbwgC0coogweTzdWlRwAS9unztClOjUGdMFs/XrTn2n
DCzo7NfLcm9sBAhy0GfCVIanvVbuiyje1/Gq7pSLgY769TazEtksjwsmsrzMeqn7
3HXkvgi1hlCRpQj/JzUbvzLRVLY96Qh5hPPSZhKMcDPm5WHFtyRZJLjhf6O52SsW
GJotKaAIy82OBNUL7a1GzUbAuH7KRTDOO7h+Igp1ktFEKfFRklwSCDWKPn3E7Ko8
t0GMZkhBB2LmO0Qkmp7x/lnqJAcWRJ/icJVEuypyPHaJX5EMA4Y6vpfSV+jY64d5
7+w3JtazUJH/WQfhOq5X4/VQy96YS2YRPXhx52/YDfEZTL6aIqlu7HgaIs4wN+6U
uxiJMtIYzooamOHvilMVT1VCY54gONISqIkgFMjLuqGbcMAs0kOO4+EcJwkel/sp
E6mwGKw/1IAJ49EqbZ9BC/QH1k0v5Vd4laO4n2pMcTA=

`pragma protect end_protected
