// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m+cfwLv8i/jP1G5a37hXqmYdazwjtsDXcgKq8nIfxOL9cUQTG+0aNRVfYSiV
VSSO7RR7MLzNCgRMCtxiU4lPloIaMCoHI1ed/OEPTXpaeAsvuHdnqvxujhxS
pY3Bh4p9IweySsCMmrhFJDo7Y7r9Ow7hA/UOruTpQKnjJH4/SAuMjE8QgGai
mQPtqjrrHxMFN9RKGG7gr7qn8mrl5RrO9H5on4FuKXuncfoCxubsynMB7oGV
SsukFP7qQ6c5RFFYAOqgnHMokippZOsed78Qv2dqMN3T8/cco8q4g9ouZ+0I
GNj346Ud30CIlUhi4QD2bw1GqHWOftfggCRZZ5mQaQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WgNKJFZGWBIDEplA465UYmYVAtgJjMzZzsCsmXBS5fqMceild1wHNzra9Otu
PbDEkMJGA/nVXhaujB4XGipXV/mdTtZRRsHNFIPkSBvOC6bg/uOXHSDYWwGz
cJg00oBxHudTz2gDJPnkz8N8PUHBOnOvuzKntlTRKAic45XcDcMtKLA8goeV
1CFaga3qnbLFcJIpSHBNRjqH4haJZpVZEZvT+Tj9QYJzLkq70JhnkcFqTw4Q
5olgR07LfbFFFGq9Eqk0KUwxZx1I1gOxoGNdaHXfeyFgif4lYi68mGUZagQi
Jams+PHPaudLtvOukVPSHD/k2oFXaGQo5DXV8pjd0A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JYz9JoYWVwaihpVtBG17jbiTjqRmxWQ0t3163yr5XkXfB/c0TV9i2Svlbat4
2NTELIeSUHOn4s+1rA8ssBIIc6HT6xyHVeNRR/lqQ8daoO4BJiPhnYNDHn3R
SkXuUXsQn27elHbZSvZeyWWFMVhuEg/PDjJZGkTSGwotDO0kTeyCI9zhUsA8
Qh/tctORwBjvKZTmJTLAxNtyYGX/9LvD6hZ7ZHZ3X69882w5zll45LpJOpsX
/eSB7ZXZt6gbd18G0XQH/R/NO//P4myRR4uviYWPHVxGeDN8OZ6ovQTqZgb5
/OPCh9wBWgUPwpCtZxELg0pc9sNIY2p4aAGs+zaYLA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LSXYO5ZLycOw3zJx1LBuN+m9/8swkzYxGHk4PHKK/CdUL66NtzKn6HWnf/lH
7uhZYxAzNLBhZGbfGvu7bE/+enRLwM+DbucEjv4UejWvXbmxqw7LAeXdj4HU
Hg5zYSHpuCBjgJWvugoN6mW3GON5640Gz/32PYX4b549jWjZFH8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
m5R9QM5/BG9vQ2hSpYpK/BictPc8fo6uZ4XxgSdC3EajqP4S9G63tP2f307P
sKYr+o7MFzQH0H14g7Tlu64KaS537MptxyjcdlmXfag9CKIw15w3k0IONnfY
GNKZC0AO5kucrxzwonB31lKRrNukBYL6J54RbZnafI9wf1qn3gwJLDnzbr3O
BjIOMoUZQcz9kfugedJ4F/u9f1r5IpNn1pZ8rUwxzICCUZ+pI+eCoHcsGBFD
0QUCPgNqjmk88tdl3+jN88j2fBA951STA8zsZaRPviRnN2Pzp+T0u3WuLMLP
1zqszMJXBNG1wrTky6Itb2Tu9E6c3B2Zc1zjNcCjENcneoixiNYanw40Yqct
dI8l+LAjP9X7qOusCI9KQeKEeDHLKJdEyfgF19E6H6z5JojBQRKCdrv+DPHi
38qxs4t8cuiNXFtUwL/myy5eYmIKzYAHOI1z0xcncffvkkWkvikfc2RWh4+l
SM01QCfj5Rbml2Y6gXNeQk3BjNbaVGgU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FBQU0RobmUNFthod34kPIADU/BL5Rm2Ap1Ak1sx5yapt9SOEAk8uHe5ZmZiF
GLFFeiuIOaAzEkJDWnIdOaJT/1fQN43RUJQDOE0ztbksqRpXuuvSPHohUpxl
R2ngPcj1PEEran8pwP0jSd9nvoq3DImVYdA0OdWtIjED/Y3AD2U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
V953OrcSLsHQlqjfglOHJlRdAouD6OIqQdnThfUPEpIm3yoOEoM/YmBLmiQU
Be2dZZYL2/q7KGwCIx6/Gjz506krlwQZaVuF+nHaaGx3YFaJLqH525TVQCCp
KgV8lxc/FgIhdM5pP7CfGBKU9vFFh/pQyXwFF4ZVtUNfAF4hX9k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 42320)
`pragma protect data_block
tzmRgjAQSpAS2AJWt4XkVO9KQGJfjvsVlu09911W3mLX3husCKvFETclftj9
aEGpoWn6Un34v1aPCsEPjkwdPeDxMGJsSWfnoeHXbkUEr6rt50vp9mdbK9zH
aY020N7GSgKym7A1lweBSya6Rjt9V66L7gGcDhgBjxuv5zKLcAX67SY+aFQc
wnbG1XxsLBO5JJyNxfJvwGbZtrJeRIngvyFeAy8KFRK6EXyBMMtjFHADAYON
g9FKcgXhT59srFWj07s2Q5sqCuMMhn+xxCAwwq98FS+S7+ywVJbUFGT5Adzq
A1xZF001HLTUc3mAs+tcpR16E/eGswPNS3ICtmAK3nPdnsEWf5Ca/NlgsffV
ClXwgF9QPkFnGWEw+KCZMeKwPQRQIlQRT8/5bLIbUnsLVxRU3sNZsd2stPv3
TCVvg4L82yiZsA9W07Ks0GyvUuSzzwmyvZyKCHXyIKMhAuHC8v7M76MO7DwR
EN9LHhKjeZ96walVa+axkXJKUe6Swc/t+UhsR4N3fK6+wI4lqHvZMSnKjo5A
1dXXzjKRe78jyjFTBuHqaWRP+ro2CSFEdlsgHypD5zynP2bu0J5Dv++UNgGB
KeUAp3fSZZIVjmp8rsh21mpLcUpz0e5lA2HT5Ln8CClyjGLs5TdjfJm0IPcy
cHmEb5Jz72nDUzBZzKmn29RT/zjpTurvwJwClqhAvXrvO5y0VKGuyxmRDRAm
5U9ruJVV2JYDws8Z1KkKMZeQdLE5KBZz6khaxOXmDJdcNLJR3bOrSBQsMXwD
XqsiItYUwgZA2shuU0TCpipGSbUKMQmOf6vxU5iKDYqpy15Zr18B3g0Xk3xd
u6wZ2NLer6Ik2PGh6AhbsCvZjqdbhToT52qfwWEQZ3yjwMFV+uBauWOl6+mg
b3LT2Wmpq6GqOw6fZPnPZC7VyVogD8EABq8g0r5EPj0GpXOSy47mfqyCqjvE
Xkx70xrmLGJXFiiyFp9re+mpEz4xgRgxSlo1skrwFzKxmw2SFL8ttNFBJbw1
mwH9E893miQ/aY6BnjlYfCUvs4o9jbCSRKmr0I91cHz1oM4SNDwX331AR8f1
/S5vFxcyBrq7oPLty3HZhCFybBwsSZ/jA3ZA7XkJKTMjwN6WBK5dGqdTj6st
nEKp3LB56b+8BrDN2Jtj1jaCiVQPnFS8dQ1bfl3JrLjxsLR3LUSa6inKrQ6I
isjoxtUyhYX0G6I1Hd5tJEhqk51M4SsyGy7N0RA5ZQq+/o1RvuLdsxOtIiAw
PLS35Gcf8k6CV7hujGb9ZWSR9o8T0rtzdZLEgwuNSSKL9OivSIqA82mai5A2
PvkllMlACiDhjGQkSo7TeZaptcyGz1BOC0LU1DAKpQBpia5j2o0hOvdVrJRE
+1ChcIy0vXKWHE8wAepeTmZAuvzrqwyl3/1r6rgc78uCjASuvpihBhzAffpm
Wa+QaaFqRB3L5JXEtK8/klOL+x3j4viRgEbcn691tvSkUd9F+M+Tl+igs0k7
BT0cCt4yDs4VeUmZMpOFCaJZSbG1/Aa0u/GXVfXhYXca4ic4ylJmU5/AW30E
BdG8CdpY0QQINuqc/xYPe/Yz7T6CZB+stbx++Y6DTMmZUJ6KCAtQG4evNFS0
mZdMQykJaeAoPY1uojVqZQCLWhj9jYPxXiFyQ2uvQLI9uX5h10MOMX5GCQYa
AjW2lX34Fr6TUSlfM8Z6xOtgWApiEuev33vU0UYeAmt7M8iNVW2NyEETicFe
38fXyPTkzMWYLBr6/RG3UzUfwaRWZCqDDuX/uOXfs1IwbfVvrmIkKW7U7onG
m3jTVsoD1U4ZwTmJQurZ6zRov/+5wOKGJYLpiBPaOGZTe4R6E+1z/xH+z0o3
+0SpmWR9e8a0iFzzvRjX8NXpMFMmo868vB9CBAHSnHPm9qrVzF9G4oh/ZHsR
mjx1nwQEqHNyDd4smf+eZtamdEdd+q+Vcx+EqcwhEmffizysaSTRYyRbEA3G
JUTRV8kSk0cSdIZQT+GuHDL7wtQOikqFkQWVpq08BSwfRkiwc9fLbV/rJys/
iEgwqSwujt27wfci2DgoNLm3kCCTbqIXRzACeJTD6V9Enp2xrM9+yGkG8N2x
Kg9T5yJftIFmlmlyao19J7+mbY3uabqVBSfYPm0DAeqMRnGe1tf9Fmeh6wLa
zxXDHufiCAJua3bYAthB/mfIYTPlkpLXbd0lP7Bwk5+7PnELPGo/kgMPi1ej
oFRZusf3TfENjaXo9VXbA7tS02B3yh+7L7dKV/IkmgY7R5MVybIcT57ua2t5
GnUEIsq+/ePEB1+NbPErCU7BHJdiCbKYwVq6bUN28I3vyWMa6kkPjhadsSDR
qwVzzBFm4Miy0dHvRrW91y080q9bKW0XoBcaomNFosn0Q2h9Vnyhhva/RARm
xdntaTMC2pW/30QogmzG0EMzZ3531cHIy0f8IMvOF3w+dhP5sS/a6Clvg0v9
rAQKxSEaOUzOLqD3MXCydY7qK5tED1WyQnTB/soSDP0LB4ZswjPhw+Ca9V45
kGW/J7HPSLQXa+ohQ00Zy/A2F1qhLpEo8iMArYMbAKkuqDZQnytlL0Mxd5cI
/xc1C0iTt4tPMSi0CIpqRbL/9oL8byNjALhfnZ9j/Al4j8GGEMRtSctaiUOO
36du2EQN662tk4HOfUaX7DB64EJfr6LeNij9MkTVgnCUlee7hP9QjUSxDKBW
RPiMlQbzh/FZwo77EBUUVwPpwZnMpc4F/KZxaUYhM1frRHrWk0IPyPxd3RKx
q5nhM6cezOlR9J0OGmNs+OqvempbKtszNXUJZi28gENEFSEGJSonvu1p6TSb
wWQJhjIbkQpoNr9LKbzM62fqhU/8F2EHbz00gL9ufwOCcnggJQu8d3apZwH/
QMIHsA7HX2scO+CdHr88JP4twWFPPjF/ZO3scWzJ28E1RkoEUHpxP+XnLViG
9gVMz+KM75uwvjNEmsrz8sxDwwGRzT9j35dvQlNfUUeGv7DPlbhbamNOwhTg
TpUQApSnw+pG5tMuIjAMIJW01Q25NFdkIt1E5fFNYE/L9Lq3lg70sDm2d/m+
hVGzEbswN68uD0Rni2MgJCFzCQIVkg0wHlmsCDbl1If1NL8wvU2TVdkgMQKF
sK5VwWdegXrOa2x8yCl0CSDF0j08BtEYEe9F5HaTh3Q9zwIh+63jddinEF0Y
TXOJCILMjnUCSCeRPomvpMWlvucpjw2WKV8F3RgYnpWrbR3g6ydwujvddrU9
d9Z3DDwvPpS6uUQwYuk7gTRJuEAX1dtEaMot1RoAasCgkhUQ6GjKy6iOJbGO
LetMr1jevd+jbgYcpzFtQbukoc4RlCRmZ+43AM+jnl4S+0txQ39YR/L6F9GM
SfWiksVocrrtrhmlybNGjKIR4zPHYoEc6hZ/NdRYEST1WOzpWcckn4KNU+lC
6ZwVRItqg5X1cTwRfgYgghSefqAoSh6R0UpVBZeXsks+SXq9XuzAU935vw3R
GNI2UWBigsuvi0/31i13SkPviZHALRE6FcpR/a0HtP6p3a/fngKa1ETYlTh4
wCkuAerhZmEgKLTbqTEBdz8bYhOdP/TCGEoG0Uc7HTXrkgKP+jIJjxvssn4F
kao2lqV+wMUzWCYAsWbADHQnIe4O33FAqSgVisUwHVqn43xdRpe9l+qcSq7H
Fm/BLtjsYbC/jOBlP8Pkm1Bg6gDtHdlDKiAUnuuxW9OS56E6NjnhHTy4erFL
K2h4WbQS0HIHDy0L12NQUi44DrTHCyZX3FYHBuyuvpW719ZbhSzfcGrRy/Ht
pCmqg9hwR0d3ctIRI/2uDy1CzmhPsvohE6ZJZ0sxM4HRfiGAJYjz8EV8hej1
og91EUISwXciFJhKH5q+tFOr67y2XmjIfZB20p4wa/KjLuXm8Ky2Jaj4L21r
Evs8Y4xcypvKdkFpw5jG/oKoyGbJCKR8+JssCncjh5XjJKWWWwxAERltSzWc
jIbfPnHh/VfjAzTTQW3v/3mbdLFNptnzE21g35Du5Rre80wOrY8utKiESFpW
M1qchPBlPg0FidlVIWinMAjFCiEgoxcIE6wgzD9/tjRn1lXhYDA+gSkFZ4tS
koIC+r3GUGxG8XZvPVf731c9cRtSFwzupxiis1MlK+VkfA99rTeUO7aAq7AI
KQLYKEf2gNTFdW+F/CZuc3JLrHBOtnRG8FKUQIM7scPdLbwpMwKWiFhAwx6o
3hiNc4+/0ljVoU/X5K2Y7rp3EL7U45zKcXE+poL/pqyT4ylD7U2WNLE/DQux
Znv5JHfsOjXjS4s6bdt7XKjj9pdfKvWkY5RIzhAP8Gl4BcmT9X8lhimK3gAg
he10WYz8s53KlHJyLRHFZZgf/Ch+qk2jBArmGf98e/S+vZh2fYHLr65U0MGn
E1W8ikDaTdpqHbQE1fcoVyS0ifl0GwYmKJDZ6rvMkTEZb3YzR83ITbxa1dg8
3ns5cCLUPY9GYaols/hSpiq797KqgStClfmpJTjhDR4OYwZ2MFisvIfdomSN
dBNqdVcVdha9ckOlUTEbewfqt2pQISxB+vmA4zTsYyTnlctPmqgJcrhBfhch
WWOLFsRQ7aq0tW8U7waTOL7k6ngB/Y0auYjxECQzrJWc9MNfG9IOM5XtX7mm
GN6MaGm4qTFeT2ep6mgLe352LmFm21fS14lR28gmx2+uk9jwdzVsa57CSKUP
pxDNlUs2lA3NwGNF4nPlLqx2gEbyngd87EWc/v40oPLEUNgvZwqh9nGpUifA
hj/rDkV3AJkVCFK/1Q4uRAQKbnXTa+KKpgveJ6j1IIBd1JL5HymS10UKKtRM
XH49uCBd2xiBPMcejzQFJNS0xMTky0frasQ67lv1fBN5gXDgDd+oXB8nSGPQ
6xsJXiamP71POyibjTb8qGagh15oy+R0ZYfLXBoE6UrhaWApFxNXP/tumJBy
SaRNveSPGbdU+xN+1o4mCPoiwrWqr5+BZszeKOplwRuNeO9qpCmqPqegGwz8
Sh2NTXHZZD4xcwNhsynPv17IZYcVn2+Md4xz6zWf0vJhE0uqonGkzfNXJvzs
kMm3YiI4GtlEsaoGv/C4YWwGB3isCV73fMluhMDIpDqnf7twCf52bOd03Ooj
2cENnMalATLwbG+/pOOqP2YfiMiezFWL3UOAgKVg7o65fSWLPA9zXboeyw//
iocWBduQMN1aPwDkBexMF9Qx1PKYmRyzsFk7UlT+9U9z8OWMeWfzGI713Kxc
xy2e9uKQzgwEnomLkkaE3868ltk9aAKC6fBKkuVCELsWV20S2YedcPYtLccR
Lntt+GV0sLyq9rp6tZtsofgprkLgxvaggshSSjO/+iE8MX4/RJRIG3F23ZKV
yUgXjsqtvUGg1XJdOpTry1gA6T9mOBfe8CaRoI5/WkPRJESl7sO4BxDoFAPM
dFfUUxmlHdAfqjdVEXgGETwnRvFRKA/jsbiXxLlVt5Rxkgllc7davpsDbcAY
zt19AhvrSJBjWakV/+t2zDUXpO2tutVUQB0a5BsOBQXcTIJNBO57eVnyiDTB
FDY4Iv+5fxzlMbDJ77os+IJsdA3tkDmio4xSDe0tPDZSh5BSoG88BGrOPwLf
sy90Ad3XMGOAqTC6oKKAjies+ICaxg2jlyrQxabPWvYYiIQ9LGdd/QbqOwTw
Dbb7woAnV4i1/WQTfeS4zESaS8xYYX72SxZEBkT1Qx6qgFko9PQp922t1DxS
RjytSyYIgYtNB1QJ0F3+0poOAjwaphTY1cnGB0uylT8AfloboEqTNlXjUx1F
lt5EoB2vHx+8pYMjDzfTd1Igr5K3bwFfQH7anij+YbKb6qX01F/9DN3wvG0f
7ipzvD6v0IDB+mouzjy2+9QxrTtHLtGcXG/biQR4sM9cwnkIC00A+YB1+mWA
naOXqNLB2Jdl6qUAsED1DswpA5OXQYF3jOz27KZSttUYVb8ywBt78f9MsGWh
ZC+TwrnFt3Efk0kqdn6fG10DtO414sVKH9pd6+DuR2G/SwrC7Ygr7OP6X5m4
yny3QbvfN1SDUoJtfqqpu3Zp+LGMWF1vp5a4SqNHcPpmVANCLip3qS7dl8RQ
jeuPcfkzyNClIu4g5/zCU2MP9At/ZIIkJO5Kw2pbdy4CaOHfAg2aHxXQOrH7
VuPW/CKmFN+86HsqilcoEsnaBmsCHC+X1d9gckDoTK17n9leA0LfAjr3I6Uh
6nwB+YjPe4Bn9Ho3VCSe6AgXBklq6qbp5rQaS3QdZzIxGnlf4E8qjs2KUXEa
ZTTs7NEbdRtZkoHSFQNMhM33dBeBrnp9+cQ3QSdKQSpfMoF0dANQTpKjiUFU
0r3lDqyGWBHpqfUyHQ33Uk6NdPvEB2+4RK86M7d5Oj4U3Y5hBqd6jgxVdL0Z
TDXcXOCnyglGgqJotiqTkTyUtyldx3tk/ZoR7wiTW59ZXbu1cT1wBeXACCWu
PE7UU4O0cPMTtdoC/WpwoV+5cnnJKfT5lMb7CjuYiobqhETwjRsU3Yna/g3T
hG/8Iau8BjRR2E14rR293M700yEd/rCNH4lmLhfJkLLvbyjsppv39GH8LujQ
sjnbG7f0bcu8YhMJ1zeVoq64hXeMKErysfGB1MfzbvlYQ7+V87JnLDiOssRx
PPGR1QcoYhKXznGt1LHpWUsSOC6gYj9NbfdnG0BIRY7RHBjOCPLw/wP9Mzb+
EnJvaVV38bXAZfISPkaS9IXzuGf7Ieiq4LX0XQxWwh58sjJp3mMEIRk7/Y1U
/5r3aoIdG7RMZhlvFdPTPJpKEQWYHxyJDz7ZafReAvCRRCOfUQQ+vXr7litS
hJyLU3rcKwDyG5YGAVYLrveTU+Ze6SPzUL1MynC2nHpXsVv2IQWUiSM8jVPs
88BeZTAWvFrmh0evbgCzkozW7aha5TiS8YG1dZXxHgqzn0a7gsDG5TBjlmKJ
n3jZrdoeCErX0CCanf+C5IOGDkaL3Ibpa5Q/VVZQRVfudoE4PqhdrJ5BWBLq
D52/RdIKkSvFX64EgB/VUI6+SO0IKo45piRAboBCyzTofFv66krih53bl1X/
7mttmNS+q9tZzuT4RfHTSWw1ENTFICD56ZdALWQpKK61dFYxXmWT/DHAzIIk
7HbqWab9lnJHNKFT4AcCdZznsrsQkpFeEGFUHG7Zr6Bp9vXSiOs3T3PYbTVe
zsyYc7TpbG71Eh/3kRpfzLHB0SjZYM45bmva5q0ZQm6XbOna4wlg9qE4EB9u
hAppyPxJeeyvcXMo7UPq5hDH0MSm3NFVAjTyYikqD6pctB09uevB0Q0R2+yK
Fc8K4fkS/AW8PhXaUPADe2MNV77Lzg4wWOhphGNM53x6Aa74GL/L4KB9REBo
rLNF1jv/l39WUymAirEk/M4QKL/aDGlNSIFmkvAxaBm/pHpsze9Bd8aNrxPW
WCkcCaUyu43XKVR2a4DKsZ1Ul/L/tem0K2365uSE4KfPPByKC2vXyhbdhK84
VIs9zeeyddV85KCwaJFOoAqb3pmLE803g+7cojtumDKQOj4WACJ2RGCggFaY
r3//rxzASmsW/x/TlNomo6GIgnGggluVxE1v/hroH7qz5WhF5z2qV3aU4YUm
z5cjp6yOWtZ2ixrA6GvwHmAIQSdnijL53nBoa4Ni/0awbx5ZJ10WOmGc9EQ3
WrTKtV1NyYg6xht1tqIfuq3bzk8QlLGWOiVeGkqnSnG2swSxADDDZ6OGvvtS
XVA4hUz69z5lqi20rvFX7YS9IEFPCqyofaaL2BYh++DArdT0nfTT7v+LxYdZ
nzp1kk4TPppFDhyXYoqBG4v0SWCPWF3MMp8FfzyUUzHxzOX7xCUBDlUobN1j
VGQMF+7T9g+hp5FVW+SrDWAM0iPLHwGvrmH/hq3n+Bv2jIHvZeVNOeayiYxv
3x0rNJmqjTfJl7zR/tlhDHYwEP4GjHJ4OTtODSdHeFlA1FnczujiQ9iVIxC0
C5/oFjQpBfCQe28u8dLo2RyvCXjF83pYlQeZpj+G7FvplQgym+fHMH1TLwQt
xxH2MdYqgxgJcpGS3mA3JiPV9zuY+Gp2oWvrULGKTsA8cZruQNqHyUvStZOZ
n4EN5oUcFf2U0G6I+mSOcIP8xT9hLY6VHPsNKkEu889H8QPnqOMCJ4cSzRpG
yAY6IhRXolPl2sQhUSmDXgxox9NqPn98SGLpR/8uDbQ4E9NcrqvrpyFlQXm/
sky/A/biBRkIQyqf/hi/5tX2Sh8PfMUvPcv92W/pHy4aUzhN8Gms9AkfoB2+
KixB2oGRZU6mQqFHxQ1o7sA5aj79K95/vu1Og0xHLzdw8mcgfvow6sj57Pk1
DrJ7fHeIp4JsYpJsM0yLKqohQLZmH21UqqkCcYiPfLyr28I88kbx7QWYWWca
jBEB4rIFMdMYYs1DIqUkoNngwQRn7p7PMayzFV4VbdOkmvsxM2o26ZI34rCw
th/nOH0g6h1d+7+TktwTtIuU7TWbLJ5YXa/FgFlcBrJDQVsZVjt55HGBZUq4
j+quiCilUE4Rnuuy4ddePJoJfO2g4Us0kLE4f2TmBaw6c8L/fj9M+0/zM2bp
jfbTGDlSZhtTOyspC4s6V5O9U/xxkEouVw9htKFNIbo1X9B3MloAyQAsC798
vot8fSG+KTk3VR0Snus5+K+tnX1uggd1n9lLSF8jVCt9U8w8powFXobCcEtE
fTI6gEkZp7jvSyta+kiZ0ajwYm9lUJornxF4WygUK79+6shuNNhtXf5jqFm3
canG18WOirBdY1aDf7sm4NBB6+iGsNJdU9/MsordR/jE4bIycSjUX7kGzcdB
bEv8WyGyWq4gg1aAqkiq7QH/mtu9M76hYkExmawNWeUjPcy0A9xEecDjT/xD
vamiOIEhR2expd9qKMCc7BTVWz+gVYxwaujIN3diwrCMTR2krQebxd2hA2DR
LlGv8hV0NsqBCkKhpU9OxsOoknV1meu3CvUVJYqiZjy+GQ+isMq3G7FQL1T9
++lowMzxYBxoVKPqp+xYpu+D/4vTxj5KPEMjCz3TWu3FIDuvIlAIMQeOgmF/
pi1f9a4KOtcDixysuz+toexOdsboKUn32mJKEuUkK5unrhI7/7YdbxV0mShw
TEfjenL+oMq5wmy0owsfDHmezDpHApig6JcN688/dOpnYUHH1KpJ65p8ltjg
Za17o+qjHHnZy2TezA2xVeOhTU75Q8ZYZrTpMuA12FxC732l2C2M8VskxALg
frDIDmf7YzgJpUsRm8Q2lRYRouSH2xMKKgbrRMWOtwPndcUfs7Bg6qGDcLSA
40QmqYkpnMx9/XW4xF7oNt0H6A+B/Of2r1YFkpL2IVdS8zwxjI4V6/wxf3u0
WbohMmQT4musc2chYvCwUgx8XrHo/A04Myl9kkzkzT+t0UmuprXVXnfr7fA4
mu0N/xyVI2Z/mHVw1YtY+3e9zaqTrE0bSfQrnqMElV3PFwENW0DXhehD/+0Z
/SsV9hhS+r8MW7mVGfCA57PiGEUnOLDBvV5rTORNmCJsiglSF+lsKt/+I6df
lHZEDUsZ6VWzs7NKfkGvHwelkJrJaUJ7NcE3FzAZ90JmaslQOSUFX7Gx2vb4
QSWsalscEsr2Po1f55gTwIOasAxpAoE9hDX4NshYKuA11T4lw+PIU8LeTWHx
ac3Wjer4J+XOizy4DmJqxFjZeC0vg8D8dFq/SBCi0+TdnD5QhMysIk1dPO08
Ypn1zIfwS/9QYOyoVc6UZySTAmBS/ympnFgmt1qsjcfXE6NnCBReeAW54PFB
7XwHCRWyHk0LAReky3nUjHOLi0BZ8VR4AbGN04hRikrhytXakitc2g3TRhdG
OSAM01G+5MKEoLwwhiCSUy1vpn+hLdjxnTq5bST8akLNibFIWbNYsGg0swTo
s5I0P1GwXF0LFGRQa3nPGpg1ieE84yC5w+Ml9Kcp07VbizYRbFt42gGSsU0G
8Kl2B3j1EwmyMBiNdogAaH47/oHi2mpWa4Bq7zt8MFQ3GaFabNi6howrpCb+
mUD/7fVAF631VG0qiKZ3DkYPlid8qUFzUoBQ1mDMhMDh9IPVpvWI4/LfWgDp
+qSRu9Rw8CtEPeAaIqFbSr20venSb87idYXNMY+8dcachbxJ7ojZzx7qJet9
kVze/VELnd/ffuGEMmYx3Hx7jNZtjm6oHNLJ4mrVsENp961wM8kUpalJ1Bp2
xtSljdwwlIy54L9vlDkYYI9Ch9W9IahBAgTK7qb86GnIiCT1Up5Nf5ogwHpO
lA8wj5FBz7XKQmwtWiY7IQEN/sA3oC+LS5NEvnm3siO76pJe9P8VyaRgCvQU
NCroHQnk+uM3oL9/TvjY8iSg2/yF4Ag/JZ3/0Zl1G+huzHdHk7mtZDkIW2xX
HN6NEbWMzwUqM9BgFKWULOaWprWX59NcBYuPaZOXgP6OAwFBcT+VHtf8p5pw
Tgvu24eELYDSgMnwp24oGLR01h18EpSAn5HwcHyRp5tShKvGbdsnSFIkHZEZ
dfLO4MNaAjLtCEAUZ6LJ3i0dN3z4msXRpXr0FROp9+4TpRPlfHEJaNYbItSz
ExAP45HnQNr/ytSU4UiipXejBaUBD3E2YMWcUI1REUtT4KRaTgZSF28rsvkK
CaoxVGQWbA0v62vezY0mDUqAnppWNwrxJfpPP9H69b017nIszv+JQHsR3+6s
uoURYI2QV/MpjQBb9lRkO8pbUwcPnL1eYgQbM/ggwWYfXZo5XDW4p+P9ArIA
Epdn/RICQsZEjQsH9Fd5UFEwaDZvez8VQzorIHLP+cxEqu/mmmLGy3GVz9kA
jd/UrdOnh4+Cv2Eduo9LtdnsnwmuRHYuCIiAsyybf+hEN91PxwGkA+BGdcXp
E6V3d0Ru2VfQZ1OjNMb0OrFe2+82t9AbKeM9yS32Mz6PRIh19s4EUW291AbZ
IFp9BeXtINQOzQvbWHGbIjFy9VjR+CpxePfQxDBk/XC3JCeXdEi8rB5/ruMK
57pkdm8Wdie+kZw5Z994lnLq6iM5sfOmIGAb/K1as8cdpP+t2xrgRome6lxf
6RUwPqyKnyxFT0SyHP638dd5v8dtsrubLumuOL+4I2T7RwB1Yf5s/dv0DRVN
P5PVVJXexU2OOUxgjjx+rOlHdIPFLAwhH3jpPhIQy4kEaIUvtbd9DPHVLgKI
KQJovkT1/ojH2GTqwPhDkK+Zw/9O72KZYhCVZKz8jydLDbkNod9wfpQWPKFW
nvF8Fmrs5Kj+vvAkmiaHqZnjchCyvo5MUbBLoqq/KIq+iJanTR7lGkQ/PFPl
S5unMEOScgPZriH29WnFKg3nA7lGgcdQoil6pU2guy0xwJ9ot3NDLyRvVxH3
v9KzY83pWLd2DlYadEIsXTCQ1HIscAhnWv4l2/fCa9citmySMibB10S0/+Kt
6krzq/PBBrmjeyx5PFU/hDzjXESVyXOnEFTowUk3lssx83etpRqly4G0sKhU
jrFcwIp4hKrFLbj7da6vqngk4voQAFnQqsnXEPD853kO5afcKRU95YnQMwiu
SzQBI+FViZ5qdE4aXAymuBKdZPP315dkkbbRe7Zhzp66Up/Ywz3PQ9FCu+0n
A3n+eEg/knxuw2fWNdqOryU+POmebqfhw44DgsZzBRP7y5j3ZpyrfYNxmAKM
rBRuRrRlhinRK080sB8gxREwX8CS1Ej4Vbi9bubIPJ67hbK9xGOz2ja4P15E
ZQyIUQUFCCpHFBzMGj0MbbeKGXlLjAT33HvzdO5vJPXXu19TR/UtbDBMJzat
QoVddSzmEJ8kqOk6pS7N4+q2CmMIpnVvlkrU3ntgITMSuBu1BqKZ3tA5STXJ
Hhssa42rQz7kWXMF25fWRz3bSLvUWrAxzymjPGJczCLsLBPEI+rUAWfvXZop
uWfjDdLFA23c03gwy+8kSCt+W0o6R3Z7+p9h0tGiai4tdzRb/mCS6GNazNpT
D2z+TbbkxDNsIdhXwfQnQskwlXWKNS8pDjvk9LAxdRhlNZtbsxqncSLpEUwV
V4UaGye2IKmT9uUwHT+YdCFpANb3GaX5Y89D7Tjq/daWhsO1VfYAlWdRnSav
WhHgYYTSk2eHpaft6A5VzE9+h14UdkzhTyJAEnpCYSnUdrPBEK6odjXLYQ7w
gFilY87T0QPnBY8xTcDC3MmftqicrLP9x6XfnoVhVl9n2JW6WHquwjDKIJwT
DD7MS0fVdZxUksUJ7m+S+VqkD3RQDWBkChxQ/00buhiT/AT5nnCly1foBFwZ
l4cDepi6Xr7tbLlJEkB7ufzjO2+j+ScIPrwjtvqp4fjmOIHzyZZunPzSRmsB
SD+FW09DAMIy3w0QtEGZiJKCgVJ7z8lHRUCGli+01K1/ZxRIL4S11BNbDAxz
MiV/LDwZv4LDT8rlM7LufAIg6JG1BfsZJNJT8SuX0ftPGMZHRDIs/D/AeS7I
0BCCLcwukr69RM+tl+rCSqzNCe084s96AJGI3lwugbkWHxmTCd2bdlu6rsXF
YHMbDPJdVqy1mwL9Tz9SAj/GRbFGPZDFmDWR47H2bs+CrIPX6K0ang0SH3gB
DKj8VdpjSl85Hdih7lV2PGLykXUHHgdYvon2wAkQwccUjNQs52mGwww2EyIv
yycUohtyh32UFhfc3ZjzValGcteSiSNgOUrNjp+b2MFfhzfShbq1FSnVhJpu
IGIO5+NEjaQE8YM41Tdlyydy1Nu11IXI8LSJSPZnsYqhc0UO2hn7o5pP8FTK
IBL/fQFf2wMRAX0A92fdohK1JVfWI2sEhCP+UIWgle4Ueaqbwmr2Jn2jZhs0
G7iOdqPzJTjjwAuFqwpeY68t1yfgyN7g68wMJ7z4nUY/kl0lc7aAk4PgNtTf
7/qmfZqW1TLL1p1wHOs+xuyq9JPIpnXl/DdJEuEW9m3CQNEsMofnCrK4W6s/
LOiLRU6H+yQthrQjeot6CeHtPQuZNhq90XuLeLKojCAu/mmSVMtD0MBrFItt
n6UrT6+pVtULLm2tUlNZxqB/I/uxXC2bxN/1VSqvCJETuMFCLxKxwh3YruNI
p2RzogRKO/yG2ovv9I+tqSmg+S2xRtDulaM1uvyxD/72av5Ui1FGmhI847nK
wOW+Rp8pEYxa0oXZ0307hKHmpnUtWZKrOfHmVAr0al4nPs7/L22HKIft7LZj
mHsU7YzcHGeBBmtd3SZHGr6OicsZgd0ieBRMWvc05y5By+PwTlY131gW6SeI
CrK7eAVwxv+iWBDAcR68bigffowNxSNmqj5nvLuioe/nE2ztrBdKDzC8B4Cp
2AOYfgicPJ7Pzcd9MuxQ7u6Mb53TpRgE5eNipTXW9DFpJebxhuHa0Cht/wE7
fS5PP6DI8Zz0cCenNu+R8KJiCcIVfl0V7j+GsEOcSlxKnr3G66AueWVonjqw
aK393rY3H51P63terlTB1SsotTFbMpr9MYnr3J+ZZwtjLn6aetqRxJ6yaAxu
URF/bqvDI5t9hlLisVICkgCB7QRR760P8AKxbmDPZysqU6ukMDMDxwa0+scl
3LHNKOnRLfN75/inGBGTG72/rEKF/x9uzxFI9+KOO6jvkA6oaaG1eFyQvW73
Bz+y2XxFvEZ5NwIRFy+cfugXa2iCg6iR9g7//AXrmfnxiIjAHWvxnYLsvRW1
sQgvBdIO7jZOLRMYB9JB37sUkF637pmK1K0bfVGcWghvo07jgFqXEloMd+Qh
r0o6YSr2ZupNqcLCRiEMdk9ND3L5eazpEou0xC9LpbR2yR1IysDQPqm21AYG
XgxD/1zPQbGRerrMF1VoIp0wXDjRONgLGIShD7NoP7DAZ3jVMsmtULrzCpnm
gYKtlc1Rb18io8Hpy0sd2eEvqDalkYJ7MTjTh+z0XePgSXLXvmcJpcpni7H8
5DhYL+TpG1JIj1aeSECgYirYQvPIo39+sv8bsUW/cXjvNmv8+HM0Bg1sKAjO
Z55lKainomorPUO214GQfmdMdMIEVXlmigykPxSYxEjqqsjr572aevVQvT2B
t1IwfA19NEOorbX3WEKtgtx29LsqG/ef/5QX+pthS55gZybPYMud2+9HckDG
rOrW0FanV+xOvIHb8G5EsWEOenVyBGh8bVDledanF9pWlIh1iKXSGhzPqK53
CYJ2dhP/MzB+eX3iZ0ygvifDzf9coVI6FSwUjtJ/0DPrYCqxNKwLNvROzSix
twZoifjUImEEIAbxhTq/rl94/+6nskw33gTp5RtHm9QyFbwLA6na0z05qC1I
PntRr+TSiwcCWhwUpm7YYjAbZy9J1iCIah8QyazWOf3vM5B/vu+UtLKvRt0h
yGsTal5cwpnDJj6S0+TT1FbsphsLNfhKkZkUgPqtweuPYW/ne+w6p1bfjBGl
hiiGWKI2sz05kfYTQTyv05ZhdmW4iZV9+XXZMckvHv9/l8yw4RzRCHCeHg78
Sak8CFltHmre0cA3/1AyZYu7DDI8P4cqR5wa9fKYRB6OxWtp9hH0xTv+swJx
t9+2zwlB+hAbePaX1h8m9iapauj968FZkd2WZGviy7v//EfEydVjgwoIlrCY
CFBCA+qU2cZUMkI+7nLAqAH3NCSFl3O/LFwMm+NXsWd5tOrTRRf2eBZt7PMC
2wPurTyknRmh9K5Wn5yo88FU2MdmqStfujts/8ezPaB67nArB3DtAxFbeOhy
NfKIhWS+bryjBZVp1uJhBX2ZszNK3dD6CXtmCoENst0oPeBkTtctv9hbg255
bNT5EmJKyLDgmWj1svG8q/8vEQ1p6+KL0g+NEhBh7Gzmt00NL84OHidFZrzh
1vJMq3UZud2b9Fb3hD3Qcv1UuGcxclDrpXtWj/+DJ7+snaOSwPplVu2nNtFx
MlsTcRNi2zL2sRV5oPZIdH5U5WDxhu+xibcKuOVBMHnjlg0XaxO4deU8oETE
ex/EpD1IAutSfcQDsS4T6dvx9CeK6z1qTq2F2xKCA7C8sHVinZZZmNoZLboO
dF61loeawTj/I7YydJhH/28LARA/z8CIpXLzqLhGxO+uMoeyzPHxyQgJw9+A
qXWWkRVbicC/48QvIo4LLkGEzSR2GtvhPWGjDe9DMmp+nbc3fRMUHFT4SQKY
hfzftOWW5BpB4tgRD/0JbeMrvgRnEOFa/wy50imzNk5i+QPQfX+VPv9OtIFM
Ic9UKQ06lgb9wwJVd0zL9vzkEdBucH6Dp0fjk994+pi6WZfl/atCOpt2aADj
2oj77BvzoBZS0EPa8b3Rlc0Fbl8CzWce/MyFkPBfHbBwUu/CdRfSayOjj+Uk
M2ssPTpMtGZuhk49UVlabjelzXaIjeU1748Cp3nTLGjzSwjs5zjvWgbWBrBf
P74TerYUSUZR+65jP0CC0nBzz0OodXckB0zlWTzTxPiNeNZWAKnFP7i1UJXC
IPlkGdb2+5Dc7HdrJyGJmazX8n9l9BBoZQFnsVec2hPhV8wvCIG1USO/Oigr
KZJ/0GX0dv7LnKFard3zdqLMPFzIIMIUzBrdMhQGnWkRgvOpJ6X8nc4oYSlF
8bJFxhikDToTz978acdBA5ooXtyvfSo/kP2MMf1tyPDzdDQSxAu474Rw8oI8
V5XpOVOfGRj93jJGk8X05Ss2INJtrPPSqYRM7tPn0/QMhzx7hhZ4GbyBVYPl
0be82xV5SFrkBYFmaDhTbUZ4alMNh9CyqV/cMGGoabN33hiywaHTsgcZC+NP
iMECPtngTo73dvLazeLDK9vlDYsrEFrwddmUsG9Yhphc1U95WVlKMx5ABi4U
hov2oPznHACwro1/BgnsZF5LoI5NMbZeW/yfeg/cU09y+/KBvDUuC4528oF7
TWxGJZ0VSpe5gmBk+MF1nhkKzdkIQ9D3Tda56L7mWJAf+bRjsmzPWRcEKOoQ
6LipbC/uiuJ2r3J4InBJX5JJ4MMBceDNUJeU47rWkNNgxAPIjOcbMVXf3wSv
WBYh4JFAKOsQFUi0m+pOqMBhLlfe2r3HpX1HuhFORebn+uVr+lVSwvZo6zqr
JXyENOpLYJLtflG8UJYI6EgRE2/5fH0++grHNA5TUDYkKKxEeY0eHPW4EW8p
tYTXWEmTXPPgn9dj+CKkAVXYd99y7Ep7Rm7S5CmLFINqGywAVN7E/IPvC64W
CxaHxfto7vXXzBP8jwZwRZhxC049iGlBIIh2+GI/JRgWhCZ2CpQ4DgIWQ0j4
vGPvf2o6TEayEaX15zM7BcfWv/n1Lud965Fseuo4vpDbzdgeORySNBE+Tlr5
mUZF48UKjQkH/ZkSye+z3cGEazBmZ87O55rQt7DC3GJlwH5+fb7SGdSa8GQv
/5tYbVGZnm6y9ZmMqqPUEOGl0DpSNkPLAvvEhF9NmG6OBdcd3dTdoxCzSJUe
EkixG0j/EX38A/rrXpOwxIhb8ldyNaxlny04/iK64EgYkuSYu630PEoJJqMR
ATdwdAyd5NIriwQjhEWS1BoHBkVxZ60oTWLSASikFCeZiG0oIxNnlLUXqzFS
FVug+c3y4xLKPKSCC0+Ri5JQVh9LIu/NWwK/JzGxljD2MpYG779V7NsHMr+6
iQAP+ut/R3hgSb/A9uAadf1UyJJsPHybd5VLDlm1xay/FkEv0KGT7gfx0E03
kSHQA3+QGqalv0l4nn3152eCGuPHeV1Nle5aJUp/gBjdTHwMHRKfAALh7jsT
EyZWodJ72VC3owrYslWbvYcOlNnIfbBezLv0GLbR6mIr1z/cEabGqjYBDYBb
cPnuRXjwfJz4H/T3xgHaCZwy0nMK/xsnkfnpAsqJ9/TYoiKP8PZBL50frtQa
UTjNoS+tXXPXPkQoxMBlRttjnz9PnuCD4nl9W4ULywmsZjCbSUNDJfjQ7lgV
8jH8iXGQZTBzwwrDgpB6m76+wb7WOkHcEzC0qse8RoeRWUX9ijLrX5tESdxC
YK97f3D6iCY0ysR0oqp2uFX7rbvmWfEZpI7QBIF7z7cYH1pDZ45r02R0s1lQ
+anAasMyVQLVMYIZGhIIeCDttyAFn6+0WJpnkH0uYScMXJXr+TnJiUZwhg4g
8uKXE4s5Fp4zBJL5yfOh5OdZFaVPodyh0tS/rbRLQhad4IvzwYOIqA4ZiNNP
h0jn1MCl3uPLWvsxooDvKkRs4oZRaLSa0zHX4V7jtx4Rk/ehn5MGe3ZiC5MN
Rf69eCQYpscQqYn5CYBt0ppmuV2NVkn14okA+LMKZyYdYvv/jNntWIP/tLci
FyWSlqY1dbRXeN8DMei3IAejwd9Ab+wH1+waN2ogouUAzzbnDTnMp7yQ7Wrq
w07CCwYDq/mJHVrXXd3bLl8q/kgCzYDd7XPenxLJTtpwpJnbSIc5mc0oh6qa
1I3lsMdf0Jppxpe/jTNtwegs7OUgXwt3BlnnD40Cry03d795yILMObsCApT+
l+C+oAn2cq00YgfNRg4JaO9Ek+RWV3JNSwIxxC1L0pszrl5nZZpwr7Ru8ved
131QFvh/qh2Jj+0nwxJ7rtHtaiuSfHfM+qcRAoJ0paNxIjh9ZQDUXCDzJp5G
DHaeJdLZ1Q3OMQMYtxDDit1qdXgm9UCcFJzbevidjtPIX4oecAWz9TRAEoew
nnV75y36EehFWROA3RwGtxhPeIKbRIdZkx6Y0QrJvGR73mm2aa7q3NnKmLXY
1v4MLzZoFvWkZE2rn5GrDO8f82/86fDn1dAoSCAUtA3MHvu4fAC7Z20oQw3X
KxMmhLXTFg+jpyGSdxlu78KxLtvvfHMa3ot3+1qFFOuSdKJD/rSoQ+fLIDCI
fPa/5qGei41mA4vysQpGzlXxQ1uV8Md3JOtJ4Y85MHB6iPMz/cwWIMKLoOl7
K60hZZju6wsjWD4XP9BkXBY33Bs02Oks56gx4DG+uvsn9jg098dAVXbBywD/
9wEtWHnWuSxyAwQ9wqg3IaTrRO0WF8d0CgM2+DmR/8io57kPYAuavg7uOZY4
m5q7Sfw7EpkNparuNalDhhJvWYAn3orsOKLA4a2XpCrYwsjwD1bs6+HeTd9T
73oJDKXImdiDIQkonJeGoBJwq2Cw2dmyGJd3ZZ6LScfUIqT5GNiEAM2fJZGv
pIbaiOlpl3MnaOMs/ogNKUDxPoiZU+mXPC6EusVfJHbtnE10R1VicIw6axYU
jpkfN7Qtjzz0OKZLjjIppfa5k3LK/QN3IlImptXAvIIw+lCbRYg3r1JLnxza
acbTrvEi0DADzIk3/+XbTvzkEzyywR7dBkMfzBiW1K+Uw/nxDC2WKBkvjdPL
q5OcqqhZehu8RSAwgWaQTUYNSfnwJBrbtNS9rN1bqaOzQD/88gDcRTwXcUoV
kHiX3N6Af0XD257xCp8mL50dscxCstDBFQ8tpVYBS+zDgcFJwUf4ijANsAzH
wMpaJJOclohu9VUf0m+pj1osdMk4MHwiM6vQoU3/H5tKMudJwoIzyJvs8Jdr
Q/l1mWSKhaOvDmP/XlVFRh7bgk1lZitCR/erqVThBXc3obI/WSZS1zdlE4Gg
1E1GswrAAmFJei3nN6Kcav/GGLDorqTUMVZrR+QkXw+lYwXUINjCwMzfDtoL
YY2Ev51UJeHUlrf7U1z2vp0w0MsWFDVoynijGlBBletW2W2Sa7sBHfsegEnO
ZupArSS4r8B01qN86xyQ/P+slsDD8P+MI0GG13TGFHIkiSLglZIPvANQHIBl
2IFfnuYD2bOkagO5l7D9EwnWrgVpPDkAZsnO5PAt1yD7W24Wupz4wEop0oIJ
Z15Lc5ZsjVf/I2FNGnXz3misMCQ0xBPqVMa4VGqsZW4TNb6D/E0nf5rLJnYa
CA0J4n6HrnABDPU7rpUeu7sHbb2qD4YO7xjZ1GN4hSaSaafXDEwImcA2gGGW
dj8QoPEYlzPl3qOvcvLVZToU4qznrK4/tpVuezHYjjKUbU9FJFq65lK3CWyj
6aD9OaNUa2I6JUk6HwmiTLQQku6yFUSBFZvcz70/L1GWBWFE6W0DbmklICP3
TRsQFTSXLILwYue8R7A5Cs/krPeFdpBekUTPExkZ6sZSRlALz8xiwMuybV/v
MJOiWr0Zzn0jA2K6xbV/Eq3LnvQh7PenYcVfq/2OTs+LWSgkLxw6ks0AJQrU
O6JRG1pS3OXTYxslp36OrVMlOqws/qHqCudXep1CoE1MauTU7KAipx7fHYez
tQRJVAdvP1VQShhMrKG944mkQvLpi5UO895vsf41Pc3RHcRQ6eSL+SMOdiPB
GXharRFH3PZ2MFIDcj+JOap5ZcoRlNeLodKSYybQlEqKvkuFtChApSSLweS1
NcLayuSvdx60BSuTTEM4jL+CxpHQH5TvLRcwnm+8mjpnWbXwke1uWo3O/qhJ
vgzrJquW5KRLr1t38v2dB9bpuqItXWFwCac37Rzjk+eUbC6msH2UC9TellyC
aefyXC5n/8d6MLbjow0ngL0j8zqDbGOK1Zze9F2KGiZ2bHh96x2mOZ4D3Y1s
Qk5OjgPq9k/zJ3mCrQL7bis0OEaN40k/AY8aS8ddQEBAuo3ymNGO1Z8AhUHT
FN4J3wXbW34gUE6vHqWaYD2udVFelw9BWbX6/vABLirA0Zw/lawOkj/hgfbe
EPi9E5tFk7B7TvOKkEgoXzE6ncPxDBx0rMqAOWgBu4ecGke+zdkmuNNdaQFU
MORJ8YpsnA4FM/fIwsIX3STwygUl48eNq6s9Ib1VgOXqieLJL0MBa26/0jlT
uReDF7pMZTAgJ8Qg7dzOWQNaacg7V0YbpYkGgPELT1LPvX/iwTOi79De/CWo
i6TtEJcEGLYtag9zCidCfM/5IeFvIXnsCdEQz/SeAqYzAqDX5JXVNHrEPc4w
Lwk2gbvEjKmH3pxHT8IgBp5fo7vdtpIEwCpRIyYLmryfsXa4KFMn4Rzbo3nt
zUZRt+ZVjLgudi0NuOEG4gUiNQW8UaOVg+zq6YrErX3UM3m9CeQ3R2NmZHb4
a/xPF+BhtbixGVTYIueuwsejMhvl1XUUiRcD5ycLBfZeC2ziJSCTiIeDyWWg
5b6AnMz/HbNi+z6e3NrRZGV6AkiXmwO1La03gB2xYwxxat0hqYm6yTeuI3Zm
yFV6TzROFZeK6s2iibIyfeNEBgHLDijXPGVJc/IAT0Vp/yYkqIeVvSKFJIt+
BbiBl6acp80+GVQdFctrsMFlutf57gMSD5Tt0cXc6rql1Vxg3z9bi33O8xmN
3hp4EIrk01ynbWov9Eriseri7uNegiUwvkeFiaLagUFohwWNmVDIq0fxP7Gh
RqoQfOqdUf4A2sIM1EGx1i/qiHXIqOq32IKmq5uPgeOOmiEqVr6Pz9BytVpK
bEtHCdyaO+wf6BWde54qwuHQ/rWPZ9R4fEVfewiaDKTJs+LoP8/AHikdnxKo
m6XoAufOrKqe49FPo1pBAFOUp7YViW44uDHesE/BlqBPRh1DbVidau8KpCYQ
GZ3rzf5/NxMB37HRdqxYa/5vL9ni0IlHOzA7BilHRrbKkNN9KLI2LGz109ot
US2rvRBWZ2O1O52OUxLKBxbCRqnb7Phwobb0qU+TbjiAZU+UIaEWfTuj5q97
lxkk1V7qzrCRZafhoDAbCvk26r1OjRppiUadgLRMbUuBKyeoJaznY7o2VuW8
LZ5xgFa+SoTs+Xb1tAEc8l0VRg9xL2n0xmg4UHSofy7D1qBkjoZ/arm/WjdZ
/8nL68A2z9ODFj7hVYs6wvNsgEJ4zvyPDeHxkzo8Yz+Wzh9TDDEWbeGjVIng
NgjeK93kAsKzCfIIm7fHmXgpNye/Ueuw4tOKE5eWNQlvA/e5KSd8Jpdu9tNS
BE4aU7lCW5ZDyZ+V1nH7PB+8jxp8KosKvRl/4MyZLdEJG5PeSe0Xic+vc0Fi
5Ld7GhbBtIPRCqiBeKMDqg2JsDNchZCGjGq0rSfGASVZT/Qw3WodHa9eB1e+
Fj0GmQV8t2gKoawVXqaP3haSmbKtqN94utMfDvWqK8U4yUalRajw6bq7Ml97
RRns8io5kzzC6zudZCJ28zNXD/iyOR/DVRqoadSWntz5wDYLwIE1xzxstmO/
LZ0kg7asqc7+4VdAqvrr3Yx05bTR8abe9lJFwdTQLGhPVseCHYRo/xXwrl+R
wzJkOfz4bQQGfFrSoNO7XZbzTsZAKqYvGW+C0pH3DL9W4Z6nYMrzpb53JB/I
0yhgiTj2GCbyuSz4rr1fdoEPF/vaUr5PJmOB9nEtFZQ0ad5y1V6i1ssAdCUG
B1m7TS1Qu3JFcw1rh0K0w5MI07/uDxIhO6KGwx8VGQpsembi6lVURfTMs3XY
mylja+j8dTn0asFIF1KygIsMkuJLmoOe80t0xJeUCk75MwgcJ16wrNGUsu38
vfQVw0XgCFMMS70GO/wYYSgE76dj2LEkfcwoFV6XMHgUhRcpnsiuCxL2KXiy
5mpzSklFNNXKOFaDoj+E1Mr7OQoizfU3n0gUmHufNMwZEx2MDDTmJh6xqxFo
LinWIWK8In2Hx1rj8Noy47nExA+KoaE3ZkzkD0m/B03fForg9d3ab9YN0hwu
mGseBG8JkUGKteM/15fDPstCogygq0ejN/ebss9HSH2h9I/QUNdBuxaL4IWU
TCbbryTwVrP+2gfmV4vQ4FJSnP8WOSsjJPEej9JYRZqysqMFK/df2rsVITLc
e3oC5ZfcxT+JUlLdFF8UnSwjFroGejBOejBjRsHACTd/A5MOoUQKYNi6C15R
tfzJuf29Zd+kZbqgrIYaUZw1lcpCjRHc0l2DEUVt1IurTadqNsGQaITsiJWJ
w2ul+373YrQ6JgmJuxqwzZG++awPQUQRXZ+lTgtarFOOTz0OYX2yZ9X2ACqN
p1+/DF6xCHXXlILY6GC3qG0NFw9Eu19cISQLOsNdFkYnVG9fumajKjcviqdF
tN/5mrho78s/R2xJph00Zk/EIHyumXF20DHXpXmyiWdFlDBso1Zm4OZ7JLe2
tZfyTnsAmDI7jkD2qRy/8hqjwTdYrKB6ZkH0s8CLVCvpfpXV86EmNzdZlXka
2RHYWoj6k9/PxcFIM2sRhvwhYkwWvd1slBi5LKtQ1ztspSrHQ9h5/2IKMQ3N
utEm34gKEPDLAyBxEkeeBh6u9hkNf/1puUr16f+DZRAtRz+wjyMpavfjkZS5
Elo6fXTlJBGx3ZVh5NUYNv8u3qajqBXL2byKwXwUTd1xpXlESIyY17hUnv8P
c3TDJLN4jmhgN3SU8cvppzX+T0i6JgS0avgSZCdm7QFN5kzonGsf1lDOsYaG
4aA9R32mCk2/O6byvRR9JgnW0ET51DiP9+0vE2JnGYBKeUbZZXesh72fk7MR
JvnSjyP67Go7/w4tYXzUQOG/4owe5WRCFwvNd18/vknXS9LtYXJYAn1vbLxQ
WsxTd0pe8BavYKj+oAFY+m7uP1ayknbc3E81JxEv6qdN9ahi2Ww7GoNmz0sz
Hve9HGGRJM72j+Vjvi7T13Q6unOELiixhpmPzMxCCdFh0/qC03gt39jxpJT4
FYVbLUMypibWMvK+jk10TSizCyq9g3Ia6Qb13NO1/9FTM8UL1Df5lb6YApp/
0xq1kO8e9+AjK+nOOA3tbetEwTaQUpn+SD8cxhyN3X6RD+T/W0ht7dKAI5de
E6X86W/ATveXZjhXna+3I5GsHZv/uz22jQFaXF/cvU/xRhN5/TyAnb7w0bHS
OJDmflpo95FySlcBO6mgY4FYzY42omSxaicw5FWMCB2KCZkJSIbopEUUpZD1
acYzpuTKJ5kBXL5ZwTnjYv8IqQHUd30Plob/CfnoC4hi2Z6GH0FY1Ak8AUnu
aiy1DmBWb9tIP2zcCu7GMiZ/uy7a5aeu69QKO/7JMS5mkpsuuCP/StI1HdTo
7D6n3pJcyN4pIg+RVK23mX5zvIcdCW02y1UFSIzdIvH5Lyc8DQoXNnrQvS1P
BcVsVsk3/QX/l2a/N5LlNQ5rS/3S+ZEMdVtJKu17iJia78vgsWR/SmqhG3Dv
oPMWLmVtHVBFj+7ye6Up8YnKUvPqv0rpAZUfPJ4R31zSu6Y6d4htWukHcWaY
couAgGhxLsCH9ZiI72ih7ZcBntziyMMX6+d0UbFbvKIJN6u8NXMWuHuSQfh6
Hs3um51mJz7RPKMNz/isc8D0YwA3dieaiBXP3uHPGG9Yqf4RMc/JiHs/KXiI
6EOtF8KT4bI+6CQcls3wz0uiAZl16lPr8s6uiZ9DFakCo5WwGGd03rvVNxF9
ZlVkklAPHPHqvcXLLjfy4toVoOBnG2N7NRZrEqzkOXcwEFrEiUcbk5plOnuo
lcTLWp6UYpPzno9xGEb9cAopbyV8GPQs3pqF1AewhxT0r/Pbxl1omeNATlEg
YLwY2/F4hZtUuyBgdxTy7yiBAKnYVpZ+28h9wNpIW+FePoSHoN8FFtBpNDCI
QiKqgd8jaU7Zgre8EQ4+tojfzhQMwhcofD9ch/WQDZnCe9XhHNH1TNhkm36M
R324dHWWeUC6dB6zNwvXa4evGbsuhRdo8Nhp2U0fB5VaehHs3ZwTUAb5QCgA
+uJZEVqQTzKUMmB7DxU5QSMQNMuuTQ8DRSDeoX8by/Q7m2rvN+Z4lhhrS3YR
Yr9mE3afAJI4fN1X2tV8j+U065YpxX49gSPnRC8D6BRQozPdlF2tkD45ow86
7m6+Wl+/XAa86OwjSEpGuLR91tGZ2yKLbM7kF0gqYGTiW85koTyLICxK0K55
uuNujDcIQ8rNCe7Q72mZYuhG2HqW+zwLQoVI524ktxDBYOvndUFK465mt2Ub
hYdvrl8OGmCNW2G2y/lwI9Bnlr0ptO0j8jXg/gxHNNSsOygDYCtFgMOl3tlo
H1bA7yXfTGJTVdV1RG8loqvPxsJPQxicX+O637884SxXqFXB8Pc5spdD62mU
TBx0xL5MkG0fimSXUKhZfe7QqO8YM85UzJ248O+IXp9XbTfAKk1YQ2pwzNs4
EVrP8sJWlEgsDZmSExF+4Cxn+4aH2HjLerxp63Uv/JbxaS9/H5v2FtgKtjos
2ZZJ02YbHem+jBJmkrtSTlFN+F1f0G5SdwpFrnEqD3zRXukDZK956v5Hr5J5
zOYJkRNiAb0FRQkJquHqpHOtTvID6qlUhyWxIHEVtUVPeTJyOvaq67BeguNH
zRxN5h0b8NmJX+r1A/7RM0ZgMRe4mTfd3PHeHpmNeSfp0YfyniwyvdJloKTw
JcfMa+KzB30nUt4W0q1dFM4WzwLhJgM0yNs4G9ujxElGxFSsBuLDhUNTsPcK
0Ou1p8UAmFTnfUrQ53trQ2mht+MGu8gOqNZDOrsA9Z/EeSPkRTf77JR8DbsQ
QOYiRd6YfXi3lKCT7tph1jHxLSKHNpceBRQf2i2x0UtHrAjr3eLMOi2K7RGx
9Jjtefn98Z+oRxVcS7mDG1q9kp9pyjVbjv0LBiCCQ+mGGPWu9me9g26AdPTH
OgXj7QV04RwUmeqQ+8AlQjt7tM5L+JkW8A5z9KriUIFCOTwsC7jxQPi87Tb0
Q5t0T+MaQEhEp+igKNckcbNrW05K9QDXkOMjg8jzn34VDYygOvBfdj2VfTLB
5cDXS0VHZSF6eS9Rwupr1H2/eUA7dyYS+jfwV1rEJGco/0G318iNElsFYZHN
qUgSmReTqUtReGJZW+QH0gAPKQFLMNVEIb87zFPXFeBPZnbwiJnO1u0WA8Xx
GKK3bkUEU/+N/teGDYyVTstaBEUQmqQs3ZtkEaLNWPSYlIHQB5oi3PU/Ttuv
7cJc8ivbEOZLvhRddjrimhe2jq0w+Gcd1/ASmSuQZhZ4nh7LpLpM2UAwNVw3
82cueGAClnO0CHWEZfZOym+VNOY0HSj9DEML2R/pCYSK/JtOqe7I84BFmbAG
El3IX6kC1n73UBpMKhgU1v1B6FD7wqBIxxC9QnIJU3BqNrVruF3NiZP2qhWn
I7Nof95K6IP0lppUjA5XjUyC4jm89WV3AvaVO1tQzczXtbUjiO9sPcVHZ4GW
VNjpk3IEIX7a9JIDUOfp8miA7SRbV1cGokNKikWo/IWETAxZ8gdW+ruKN8UJ
CaCtrGX0CW/47rnzpOGOGzLZsa1Yph4V/GrCq9jW4k5+nlSy8QUZaGn6EAcG
dZMKbdoTReCdPQUx4zcMKkTNzCru4en47ta1UuA37/j+rpBd25e+6riJMm89
vszxmzbHHRPmjxb6/rW4eYoUr/sXVmvVIT9lWy3eCBI6R1Llg7RlPzVjIg3a
NofiVtBwxpEHThqA5OdolfrDrd5p+r6C3X51OWJca8Fv/FmU0dQCHFK2qj97
ytQ5aCqXy5KElu4IPP4NNnL7isSS3gHwdG5IDNYe15xEosqFdse3kcH8+4E7
l/O+FFt0ArnZybGBGvoqUxBIMjU0gniC/SJd4Lhqn3cOaeyi7CpiBBFqEobp
ehqHNHEl9eqrqIVZ57IJZum3PlkenBqU40ZBW+eM/q+jyFpTWMDoSkARuDgT
0pVTsZHMqfUaTxCPIMARgz+ZPUdDRvCfmaNbQqMBAVjOeOudP7Unx2aNorNQ
tClvacpzaSx7M6ViG/L/5FxE6HLoCoeMVb/sulOCwo6SplCNC9Vu9GfZX7ZX
G85POjKKo9o4FfyYgxl3AsmAQfPV4moJsm3b9H5FGeXnp5Q6BuY9EnKlikmu
uoT+GclssnaRHbsKOIsN5eTshU8vU1GKCtmvdZ89nG2A8hsQaC5eUue5D2LA
cfEt9/nQ6QnfvkSFu7xtC6UmkRUQGwaj/ZzpAgz7rJP/f76TolCnUbWCPFS5
lUmdY4XLxkbeskfm4PmqHtpNri3C9oeo7CzujqyFqHrSQUy+IIXU+T8m0rb+
C5gp0jJ7KEnFXd1kmeZEXvsM9bFxPiPalKsQ3N7zEmVCnbnBUNOeo7XzMj3o
YmCKWEftlNjZh7kfL+MUZJvAv3ChIuZySasQuIoy4LTnWZ2odFOpmW2/JxxP
aVEUQGzh4oX5RQjwvvAB2+DYn9J8/jSSbegShMZhtBtuvFVHRSMh6eeBOopM
p+b0m7hYXzYrjAlgx1s2vkAMdGrpDq4CQCFXd9M+qI06KTQiotQtZhbJJAoQ
G2hKTJinae9UJ/83HZiUYxN/1rkjwPXqjpMnljh6xyn7s3W/+EaALJuS5k5E
nOX+5WRHtJzmBYbnDoRWed2meNnNhEo8FcqFywfuVi6RMsYagG3bn/Y2gFza
8imoEyM6LKOV/q/TYnb/FeS5lG7Atiz8xNShva2Nr6UDqfaybqwtMlsjFvRw
iraNQh3IgcohYfO8x/eBsG9FTq4YYY5BsSyUhT+t3t7L4VqGjcpR/0YfPPwI
z4mBpOdaQ/KfixU6x14EFDQGP2jnzykeF7CuoNYbVMzOjIkO/wmKw8wCxCLx
uHLaGmTZbVFlVRYfDx7gjYnj4QSeQtzyYJKAoxchBqaIbtgL4YFZa1x682bp
guHJx98qvZU3ZzpHNCopSXBMi9wUw7SJC2K0RzVuYGUdxJALkF8yqGXnRLyt
tb8e3+UzkrvopkFVFJY9/0ZOfCIHFvscjONqaHyoX8wSbCpMHGb30elhVoAe
4J4C1JIVyYrtANGwsdYUZbuUBHab59Cc4nJowDBbYxBmQA0lyeloDXS6fX98
pNhOEGTb7lg8jfGDaVJ055tMWIYFRM0FzoifaDLf/PYgq7kUqwNViCKraLW9
n1K1OVOEc8o4qp+zYyzwZLNjJDn+hUpkLvB9T5YpOphfDmyzymct8r73aUzo
u/QXxy6+I45MPD/VZ0nvibb+zX3kJYcc9KykIOiXrJkVP2ndF0BGIFHlXTI7
b9A4vAcZw3f2idxGByNOJ9BFG8VE/uTj1oQ5tJ4t2d5gUwXA6Yy02Lldmwvl
lc7i20zJwKFs3tW4cFOuBOD84dGYKnFU2g833UsRE0mr37wu7hFrQIupwLCf
+uNo8SVhDsxxbOmzt4HcCCEQMOVPkfQnL63LfTaipdBIfQBKszuhcxG6ufNt
i4ADQkg6IwyONxMPWG/duKv3SHtavmLKh0WaxIcOthWE4ZIEYLQi/2vnVq91
CAM8Wd6BeRYwq1inShT7UFuZVIrDoZoniiUDi9YCTvK+cEgQOBpwdNWwZllD
qLE/sUTA4vsQt3BVKYvk37mSa1mdiJSvjSjfo5/sn6d4PQR8+AMCmEjNRZof
JTpefDDjFowX5vgg5j2SrVlQMmqMmlANwIqnaTlXQK47tix7xHEEGvt+qNd5
W9B795mAYn7U4p6v3Nq7su6CPChI2ZIq83x4oOA3sXbk3uTpsZJj9r3ERoSy
Pn5kLozvZxfpfukWUANvhobx09ep+Z0PwhrWwEvtTIMH/42p5UkCr8J+WYZ/
Me/37V4n6moHxgo5ZjHZqiIrea1Wput+M152CQ89S0CF5+ECqzdeB+rz6/rv
NXZgvrBL5rlReSd71Y+tZs8+vPvgfG6iIQz83vo0oq1aInw1XsVpPZDCgrT5
m8wtANk7cUixJaTYAt6CPzWgMJ+/DtD6unfalclXjSipuTf3/LtLYq62bV1b
dqPXbGHDNtJZC3Apho6bxahXAWTMVcdJFIHy2eDDXpAnmmE153IOOitcGroK
bGncxkafJBXpTKt7bO/OP+/JHeNIQoe4df6INKtcaUdcaJ4bOdE3U1N2sUmp
csi7/Ku+cH7XiLR3qjkmcqFPBLcm4BFzB731XsxMT1piGTu+mSMih++Hf3wR
AAjMuxT/Udmdg4UA9RMJhTLLGsY19HU1ltieEZgcZSQ00NUvsAMPKMPB76HH
HuCGk5iwQr8xrZ9fKXeQAiGxYnqe7J9Q6L5N62ebqIw5UBFlzGNwOr7+YjtK
y9mpYm9pwbem5dQqgdgYDXLqU/yJ2pUtJi3nU3mK2pqzyyYmnAymWT7Z8kY1
fLY67iGuAq9o7zT07bh66fHavpKpp+b7CZw61YdwLE/Q2h0ME1CzKT6OCPip
y9FYyBw7p4NMg0Xi/rre344FVIPf1T8l+kKA/OY8RO27M8/WKR1cr0Yl3dJp
wmSpIFqj293FtEqlNrA9wVOVvyVdEnSWsyw8SnDp1WNFR/292jhSRySXIWpI
U0LhHI7qzGUrDElOso9wOlRiCV5TVkGNUi495ch0osX2CabmdF7ERu9sEIsE
Ko43RmhLUdVY3g0XAAMRvULGHYrWg4R9oINiMkKYXB58cwYWaH7cMQFGxKFx
G06DR93A9/5HF5gKtQEGywWcKCH1RRgq+JMVt8XIUw/CEzq23pfgRfqNrl6D
s0aeXX7mV4OayuIk4yVLjfvZYwEO6OTP19zmQ2+Ei3SavLhZHiIkyqxoFcmN
kdyKeKAeU8YWHSkg4GPcmQOqjEPm1h1DkN3820OK+UEza2CNNTXxzlU+LixJ
PZPPsUNoYi2kxMtOrLUukjdjedpB3fbuy6Aoz+tKy6mBVv63W7+vQ1go3YwF
FX8pbiTFTPJOCm68d+jxIDzxGlXHJjkZnE4c7MHuHgaSDMxwxXQ2TtYmT8ee
wOXBcTUSiF66pW9d9FBW5U0c9TzkXrjF4VmgPp+jm29vk+/TKLnbmXzWdILG
M06CPTh//s1/VBTJaV628DvxLjD02nqZhTlOWSbAvqkb0i7gQzyQvui+qpXS
eQgAyMz1XrQHk2gCKGwhgq2uw9ibDcSV/6m4poK/Z2RaOaVvVcg6S+5WoJiI
xZLF3whG10bhBDFaFihvFQVWCMQfWHu5oX5SJPUmWt//bMEmEHaU6bZ1msGT
GK4E+OTNjkWc7cNM9lvHYpgN6/02wIOQpRo9z5+6o1xoY8jjqK1APEsb8D0g
iZziO8yuPGYGuL3vyyF9HgHshE4YuzrBPLUVsbQqb2TZRJO5D2prWeZmFN+9
VXzoTg0ten8HkMgWbllJGJXVX9Dc8XjahxRWERGJr7Azn2IoM4H/5Jtnnkm3
8ixyd7ZrzymY2cVXxmeo8QKdLOj1BKXGxNzFIFGz6E76YSfDLQe5izah9R/y
F7RuPClUL50tiV4hbj51IaHR3eSFY4nDbuOuvaOJEovXdscnuZ9cqtEFuUOB
g3JcPOuVRi1n+o39UiWOEcr1BpgqHBC+DwcgK+yENQ9uiFXN/HcjAssdNAIs
JdGPlv8OZt32jkojezmYfo0E6pwbxbkDYEXERsfkajNcW1Nuhkf6Pz3Molf3
ONdtI6FRM6YlJFFCBbve0qU1M+FNJH3veOltXuGCUmzD+zVXBNBGKFzEhSMc
AMgP4My1/E3hhoQlOVVbUSOlCTVUb5GONQcL9WYeMwRly42NxRsN6yiG3F3F
PaaK/V9LiooT9128QIHhrAAQ8tPU8tPkqp+i307eZPpy+THQTQYqIzsU5Azs
LQJi/Kswrm3kQO4a7x8/Y3B9foMfRNPuUzYXa5avPVprgCQLTEjXRrFlA4P9
2Z/RvR4Y4uMdqivXzun9kz2U1nm5p/mFP242l4uvWwZF6lfVKL22fgQ8newt
SRCYq8+/+F9HYke33a8XEV1OvIZtBOTyojwaMxb7VozViZYiCyQ+3Qu3vUrT
GB8EBsEnFSPegTP0UePmDZRxuNL2EFqEfNYvgAtYwnKBiMojkIoSeT68r0Q1
bIT1c13fIm39pRD17zmVuWmO/gcfquYyt8Qtqch9Rt79R8PWWK0JE3Zn8LUp
0KlmZ5NR6TlvEEiNim4MiJCQJWjB6UhYWGJ9DogBPVY7NfvRnCpwEX/rk1+f
72b4w46RjIUbMvaHAdKO0CfNVbNDfftZLogUWLgX20+M1LgvXUkJw9kSLq3Y
fDcKyOVVxmcmUjhp6aO/8574u4zEkN7TPzpf18gNxImE9kIIvmtGPOQrQ4Xt
obdzlZt89mMVhDybz1IQN5zq1r4wL08lud9K/abwaxLONFXbjjxbpbb5nQut
hShn+3YzsDggQE0mYwS6r4L0z4AnyA5H9pN3803YJQOQ3OjYdC0PYzS95GaR
OXuwJcMAL6/q0etXF/WwFNc4VZ6uvI+awoY/cba8vKzJ/geRnGm74R6jIRCV
oT5xGoXGcS8fNegD5k49m893NojiFlAAfumCPyg60g6LCtaBlRh2vLjELBVq
8eJGkbupmxQ0TmqlgO9ir9XtbOse1WKidK8jWKhmZRMdXcl15YkFtI8ypDjd
oVv7rhDDH7LtUVWfdrUGfNyCEogrhtXXW3l6zTjZ3g/VSrk2r1nGMAuq1uLz
sDHqdwfxNI7Q7W70Wkq4w9f4id+x0CiaBFvL563sjA4zXsYb34ZrKFuicpxK
v/Yr6ur8pnSChHjDVRMuETiwYPW5/PeD9kvdTOqZ6F4xd47QpAgHrETnOH9k
0BSjW4H/MzPw51hONBYSjv4sp4sxMbwhgZdIm0lrU5E5yG6TwaFcGyO0WO+5
VgpCun8ElhtlxOPLRK916JyrI5NzJqhDm5lgVW409JsvqjQau0JDst8fqOxe
GznOqTVGnROTyUrJsYjWmF7IOro2T4UF85alNPnKaaV1LguMVRaIaxZXNTK7
XKTkMJ2wgr6tQZ1f4yyTDYBQbbQCM8a9eG9zvo09GrLLWeEy2yd/x7cw5GXu
1ptTLfza5QLKcpFQxgpDlAN9V3CQlg3iycrZ1MQJ1E9g9UfRBXdHKwI0h0E0
H7IdxXvBg+HfK4KsURRIvQGRz3e29Rn/JzDCHLsCj1FhvS+zhh6ePkvNQHIf
u1ZoIWl6BlyX0PSaQF0vrUPROBLExZbeBB2hmxV0yJEep+Oh6vkvHw22sS2x
SeuxDUf6ggR6kLC3xOcnOEYlgwKEMzRJ8GHL6Y6H1Mi43Sl4L0rlklsp43Rn
6diYDPDCEQol7DeEWDdm5gsnbvOYy78KzNnieG/NfCpaAy8mo98oNhgfI1jj
g8GeRLh7nClviaMzO9oExL/5udCvJUaX83xGNXOln1CpFuarYoD+K05cihfT
9nVB7ABMeebcFWAb3UE4LzTwLUADDzvHdTfVZhTYHNuxvHVXfa+EmbbcJuI8
orUOvnz+wN7SnySdSnF67g6u9OsWKTJH8RIUiVEAVoPoFHoWF9XONdQOq8Y8
1e6ZUGZFiYnRNgptslONYAXZZmfXlL59VPUu/WLcAQlfEtuJpj7AH7XZRdhn
MEq0w/gaMXJqM+rNbKHM/0Rte5VbJpCVSOqdphqVKEbU6cjX1JRTWHCEahka
Ilrftl3A02acdrq/9tiP3rKESgZHmubBixl55xCHF4hvSIuB14l2HcqoRBD8
Uwn2vvCJ1j8qWs6LbCIGReQZHnV34Jz63JlWoR2W0jtNLPFp2TAAb0h8WeAu
BH0nT1jG4RvuSk6fw8lXpe817UqhmGL/BTpbbh34xjh+Abr9Ls9C6teT1MZ8
D0Lh1kKLgUjF3zydKbMWZFNEC3thdIuaBZ463iMgQ+QfqG5Zw6IQ33a1C/WP
0xkFVOWLSJIs1om0fVEkM0MMtxnJNUUqNNGCLS2jMiuG14zSAUV/bASdbqIU
26asfSbYackzyEkOHJgd0eYj2zke7gra/DvUdllfwp6RVOKZQl1oUdq3GGvc
9R9VRs5fvmVI5/En4MoCsxpLgSJP4wubOEzC2Ew4L5lRfkoBfyMxlX0sGPGo
29ZKYSvjSRp0Zxs4n40kTuQgbjSNl/MITFWbJupbM18KSxFNu/yZ6qQKPYwc
kXweZBU+ypoL6qXKf/AfANU4Z2aOy2Jj9nVZOxpvWBLljYwdz28pDg7m5Ayf
8l7PhQCs8h6x7srwikG0JkOlKYJP9lqRyUnkF2aoJVNwLyrGz1wUJHTFFW1S
EQLgiW2FYm4lYFHqg2qirhSDcfIGFbtREQoF4MWuIIAY/hVMLyofRxuzFJTl
y9ft/1H0xVt+c9rOFhnY0i0eK1SAr3pKElXphUwOWWEclt4aBXZOnF6p/gja
yefdTtGL7Tbm/blo636LsNgH4mSgdY4BlKE2D3rJ5eLEsEd8M1lX9uu5zeEn
9g4dEUri+z4x7pmiz755M+LzhZ59bbmNtTz4TCJzcoWnJDTK/9dZnWPXGKJ6
tzZAKGM7Fydr0nVgxrzE+MquDHspVdolqgo/wibfAjipWnsejwbUIj5QA+Y7
fIYijiOhTFgsZFePbk0NyV3h1ys3lH5r4Wu9MhnG2eJC6WAkaJqqHh47pCTy
tmWmsWT1RCLehI3pqS5bso8+j10JBi+x5VLSa4vA2JygX0jfy9KiXPKy3s69
499X7FT3XbHhRm+Z03djUbALIlX8jQpNra8HKArve5iqBTWMXiR+4NAenqkt
P8CLHUBvQjhPXPzE22KpkLmYfPwrosNJdLSayp5Xw9eOw13evrtXd9NC8qlJ
SrwMKcXGBKcNzxZLLr4HO2EzywU78e0grlJy8XMfjFbyhUC2LtgERN4Uym73
iZWGCNL1MB5iHcArqon0rBhTF86apwJFOdMcA0ojg9ljodDEiPU5OrEIiwkK
+Kj1AblUA+SFyeAAYqYzm6NYayPp4MTCYyj2Tvk7+BQxHMKM8DSs15tOukcO
FB+yaUV//fci0xgQpZV1kN31Nv22ClQmV4S6aNqggLvAxfqw5m4xFwqtwyBc
qX7dDuK0QPyuha81dYRglVKLdtenrZd6Z7ohlkNujUzahXrdv9uAb3tdtlNq
+/weUBauwzZyUGMNQcBmnmFR1JabbYXa3NHCnX8ajgSCaIDt/4HNg7P/jiir
BZwwiDkb6kxroeuW25DskFUuyTp5Kf8HtbJUce7MtU3pRIDDiXxiXxrwH52i
vBGbKqOsp4GkieWW624OOA6JXxFLWirDuSAAdWiORQBrK1NLWy6uOJtT4f1u
VW+uEx9pL9sOtBNGHDqqN4VjwdyvLSmYsG/P0QrHY0hncPoiVLQPBpqQmVvm
iCjO/f+Si9GLpWwD40NZXPKrN1EiBbdI2GeDeqhYSubJqhPhQGa0DKAw9UIC
Y59WRRL5yA67zHkgENIEGkuAyQFrIWp1UZ2kO5lPyVu7gGsJcWYtWm1URzYE
PXQE0SdQUKxcpQ7WZ2UU0pCaY0ERelMgLBdJBYVft7rZPuhKq3ci1aAPAc/9
BKQwXACk5eC6p24dxqxeiP9B8Hj8bKmhj3n226sL5VeOLBM8rNfqYTCe3l/q
e/x1JclFnevrFsYmBw9/cJs3VFz/ILd2aeXcJ8GUGWrVM9p6Kn1LTtUlyJBg
fdhHz7wfcyZCTABHApiL3kTJfjrImNLJ1RTDe+61O7tig+WZU07RgMyVHefB
ficrIbVDP9xQPJ/9JlyftzZS9DfYzfcbJyTrzOD572B5h+Eq0gNjlC+qnJ1o
z67JomO6KF1mEFF8sKOzRqGj4Q8LwIwTXFjdDXKMuliayC0vtv874aY5Vb45
x/3g3/e4fX+DUuSbfEdG7hFid5/clh5tVocxI4zkhxDT3BVimzUk24MPfzBq
qDv5g+fQpj3Xv5IkJQE72Zx9OforybLjCfd8ZXoQuQ5fxLE9+wk1QKb6HEAL
eq01WnK2H1YL/f9VYyRLfAP7SnCA9SW+gnX1uUr7rlmOnqk8LdqpUjTEBXGG
QwluUXFr4fzC7lrfaE8xGsD+vSdS9URSjLCh1pgDZMviIFBrTmBrOuH3twpO
ILchmg5N0Sspbr9OO+CT/0qTFtlaLp+kODkB3oEc2Tq/YaOovmrF0weH5/05
GfJKvXuNY+hD3Vn7JiKr4ctbYCee/mMmvb03RM1x+Jr7x+0GgV0Azn3UL62l
iScf3NK8XDwnRXJRKIExls6VGFekipYuw0mQ4CWc4eBDODwzr3eOjMB2Z7RF
C9G30Lfwhsv5o7K0lEPdhQclBwuKabsv0oVFx+Nmqc+SFYLVu/leRbAGPJ+o
Tgu+2CgM158BAc77xrDn/owCAa0PbiNU25xMYNXYRItHTpDeI0OQS6nh+rTg
bz8y45YxienAeT6DLfzBF95Gwslp3iCXSSRuVeUrfiHPFl75Q+PWYcA1fcYQ
W1s450brv0U4zjK5IkWE2af53+12L26f6HyVcQ0UXRu/00xTIm6M+Hz7PA/h
ppFV1evGJJu1d/oem1fEfMVm5p9xKmAKVBFxhwb4ltoSl8aA+fn8z0zXuejx
XSMdCa2WUb7NB2QvahCnnZos80cLp5Fy8JwKwjF3DyoIPxhIaVxs3xB9Oe5l
GWVoPVMFWniDjTvrBW3jFANmmKCcEY+ipv35Ru/Y/RrRyGeoMASXtX8rua7Q
dSf98W9JdlLs0x1qbg1Qq2aSh94HiNo/7499ObX8FrbqJMhRwQVVt8fc9sFx
P8irhPqkySjgxtw7Gt2RfW2WXMg/+V6gXs0nWV1Se/913ST3Ttr4Jkr0n1wA
1rdA5YWt5U/DjCMIqbQcJbDz0DPn1wtI1TByWta8iDXYZdV4DAgWXdqAlVVC
hh9DqQvaB5w27ujKQkSIY2ZbsXB+tU4INU6XdLyvDbF3Q+93lKV1368NYPqt
P8+NVohBqReryEHEtaM9ZGcL1OUxqQAjazw8n7GcAXEwwpgAEDbXGiAg/zMV
vHEs+8DSc4/vQg3Bapoxf/b6eSFAjo7GG3LuMHVfA3Cppf/mx58XbuCytz9b
dxhXnNfcZcX4p+WON6s0IsBI0kwMOJEb5dPx7O3d03ex/cdb89isU+ou5Weg
jcHvRQrS8U1ygz1ztwUB6ikBpx7C5vQEhp03CCTZe+JknmoGeREKTXrXJ13C
2zUFKn8V+LUpIBlOcYw7APShyUJyuHBY5oKSitWvPYeKIHTPmd8rL1zLCndR
4rUhZMaNEe20H+xEt0miVDEXaXEp8CMHVlfXigivTvkR/xWPRu4wqCWlpuza
Ghh8lDKBz7z9XGUPytL7iXtj1HxgEmN0JEftYnMVbF/4r4T6DmWLe4OFYk3V
serKGIkTWwZbFVG8YIAJk7jEgK6iPUCsxv9GpmtnNBSoO77zYdE8g39SuHDZ
G/5BvOrNWJq9ZH5vjeiFVeeegBzaRx0i+ZyugA5sA5Bd6w5ThLB7DcJTzmGJ
c+sAPBy5m20pIC3NHA5U92iJ+/FQwsb8BdhWMc/d8UxXonb7TXsyC0Ju3rVr
paAnhL8CSv/NeF/qobkuQBUolOTNNRGoWiBzxuLsa+C0unqj/P+sqoh0ZK7K
oOLAXoFN7D9IBo1+O2tQbYVb4+Wg8XyuUjeDRqObezkhKbs4FDfVSDYikSRn
WdZazJvWgB1hCk0DLBVxRyncZ3RCCgZ9NLDNAp78yjLwS8JNaiTVDyYaRAX3
ad+6AOgqY6cLPJmFk0i2AulF3m5mcbIAtJMjp7fhdMY8Iq1BojkWCH3EbRRD
xKRPl8JZv5qr/0y8nXF4v9Vhfewxq1NqhHS+WbIQ4NluajjQ6YfSb8MTm9e/
RV0BGO66QZnYYBBEOCXKqyIyYFhiQa2LzNSeV+cptZ2brgBtcS1l3Crzlffs
Kyeuj4Ae5O+H7pnjhtw4mAS0tVIW8W5+BkB0A6UovWmAC3BY6bYkDyhXlwri
JiQhZYfK2pNW0sB5rM/c/HTFrAfPvZgSht6lI6BVfiSoUyIQxz9g9b9lLSJj
auJZRQRFrUo+gI1KzK3Gf0Tw9+znoOKQKBy0NnYOfKXenuqrJiXVvIjWpLqT
aRzmqCv8DGR8CuheR66Tw69Ndky1lfdteJBUP42qK2j3ttfWoplAd/IcfuHK
Ox1AW00yqr4B8wM+XxILfnZPCy6gHboTcYX4Ry6DzS6k5xGpc+Mn9Q1u/IdM
82HprYNYDn8TwSma+du8jgSKKYVyZkzt5Vn+f6luHIuoyx9erkYWK9rLFaRT
zmnuKDaTyjaSKfKSuB5NWuiN2db8KIs4V8xHTMHyG7wjWLAUilLXjZ+XfPgJ
ZZX3X9B6dSbjxeRDBm2wyMBE1i3VFzsRkqfbuukJ3D0qZ5lRvo/et6IK+Z0p
U4QJTaEFRBYqaq3iG7A17CXBcYzgmBptE1rB1DwEldmam4BJWRLlsjaZHfzS
tNXCNPKXLqhNnZ2hMGQ8rKXOV4xx3D8FpRZppQnFBeMIsdTap9hO7E8QP8JM
6DuosT5mYRVHkd7Tp4zcpgOhWsF8mPNaSxmap1SRkjpg+3uD4kI/KnHEgv17
6Usxqet/buSOL7coCJsy7vRMIEzOk59nWZKkQki1P7FtJqDh2SbXnMFpY49s
aRl4KPGaXomiZwGOxABhipw6NFcFWespWUDHm/Ppzb2LhGtbJpSKUC2p5Se2
g1yCKgKeBReZRujR/VbDkYu+LP21Z0QDBOWrqZx9KuiZ/DBS9znmkV3HPb1L
0RBMCncD8cvJ49Ol9vQ7YOOMHd4FBNyaMJcdDGWDNRf9lWfE3XsvttSbfpvJ
FhOghb6bhuOBzi/iCmQr1y7erdOX/GalN0J9pkFBCZrPK0eBm6Ctk5Al9Yyz
oS8mCbcmeqIXgxwoV1JbdNkCK6mUKaNSovw1d+I3nzRA/o5MyqhahBlMKU6E
axcVan41oft8br5R4iFvuTAbCnynQb7wdVaJkaNq5N7JMdzewN4PBusZ8CPy
i3eUTjoPkzZJOEZPQklueEVJlaMr5fu8WAiQid+VbiV3rzmx/4pHLCUOxzc0
jO5qVvZ9YZdglEsxwJbUuhp53lcn2qJCIIkDUb/daXBzCSi7TkSS8mG/7Fny
216jSQbxobffOrGd1SoBq0AMC+dcozYxGYLsxdGsIlj61F4UJyNav0dkiXVa
/L1fRhdOQOvwBRqpsuHSqqRw43uHFSauvBk+5sDVFqeg+7zjSqf+lvmG+Mit
W0c9PiiuqSD84d7QnlUXrauxZZA/5fwxUUTDWLZDVAa1h3HyrlLiHbVBtuC6
2hooPjowKTl6w1roW2KFAZPh70gW3yWWml3N+MfptiUN8doLDzUZj2dQ64AJ
o43DXMIjROBk0AuB+HKntU+4tYw/CGpLEl3tqW7jZ9bZafBBdD70lGhlh+2l
P09DfsPH9X1+iCh3b/Krr4Mj96rt7fqy/Li6NwG/4FjXGs61dzvui54fGB2E
uiq1lRei7QAjwRzPv13DHvhEjqx6lJYQrkAhEtJQVJ+4o79qDqwKJT17mv2G
t192pNAgmQwg+62WhuWgYxGuGPnCWtlgqreZTSRTtSO0mAEWu8qulbmsFj1z
0WIgnRyqU2g9dBAITNYTHNwCSRW7R1FzGwioOo4p3jfPxvQ/CZ5pAJKkrgxI
Wk98KVCdgWcKWdYuvzgdsoVaqf8toGXkZLPsr3g36sG63dE7/uq/VIFSJxqT
Xxhq3QZVKAoJp87SE5WuJwhyRFOayeKDEmRb6pxEp4QXEdooBZFmEOh106YH
GXUCBDgWLS2A2BDQJk5F4bcGfAV+P0dEUCFsWdeGKWe/bu2L9vZKZjvDfmf9
hcfOrozwjXgi7zLum3m6AdADgtwZYtqMMnXhWyRLQvwpQ6eNMtJdUPL7IUgy
srjkstpaeQ0twzfWrBmXy3Xz7KOn4Nb8GTZi2L0kaAOas8/cQecPZNYluOAt
LJfVTm1jwuhLdVj6Xk+HNXp5ARDme4Uqxu8SyGtqzbve+juFiu86zPGh+JsI
97pfZ6jrgmsZ2Ockh9PPULaFRQyIuoLXZbL6Vgy7/EpKcY8MCN1SFdeq98Vi
Bwr1gpIHY1S+Q51Z4JQsfLrTCqvszU6cD4FGyf2oD8jONW8ZKtOzo0cmubwk
i/byyV7/0y3KPZ6u3Rex8MNVIZKf880OxrVYPnKaQzSc/aYPyMtMdgdgZB+Q
fmlw2a8qwFbF3HVALckgobgf6SH0zHNc2LN65O30WkdtORgcvwaFOVhc1BRB
j6vxS6bn6yOcVb/8KB0Nwp+qePI+/N02mphPprDSrUzqcc8HjiocwfCm9zh7
qcMb8sG7GzaFl9E57LQEpbMSg9fVCruKrI3IvwchzlKNWWGModHLYhjmvSVX
s5UEbkctQ2by1ljfo85W101QNRSEXm7PFukHjpw2LrKVn3WXiUyBIIF2oL32
SEaf+OLNVAQnR1FmMM49fNricr37T1Ba6JQ4ElKwy+Gt+aEziH7mWXKwawF4
Nv1k+QPeRuDsNdaX4ey3+rN9hPtBpEjGJ0IChl1XrjCjrLeBH9Ih6uhZQowo
Quk1yn+Swd36Bkpb/kzwSQA3gfdFVAf7FwOUYtjnbsPzvCSXvw2N8O9H8dlh
rZAzScAxRDWOlJMh/oi/0ffeiWED3mxqIyNVC2Dn+jWey1oNcB2Hj8PfgQIY
I9Ki3QyD83C/kLwuAdaD3ZU+d93zMXOz4Lfc6Bkr1TKCsZXIpvlp3WN/0/QV
DlIkvJ2zy4ScI6UJ5ZYVH0V07imO2173DM6fra/EYlwF+YfcbxaBOP8ISFWu
1OdVN817huIcVbMLBaChCv1ltSDr6i7Mu0oXOOgExEta3mUX2XbGfSMHLVrC
0DRslLhfQrcda7dlNF59PGecRB8SyhJE15j6yKi8HAnsjxzHVHp3Z8OjgXkY
8ga8bQShZ+It4R2I0yVAGfy6TuoOHBrNDRjpYLiVwu41ssZYMbWtlXCqHSWJ
u+QbqwMEEdcvHJZcTHV9C2BCuNaIYA1IU4bMu5WIdVpDA5CHZKOlchz4MXSH
m5F1wA4ar4kOnBowVqQcVnRpPaJ6rIfgc/u9nULiMnwkxzIz1J+cEIvbLgNy
Mbqp3fJpRShi45K+nY8yP8tU42RYZS4++I2ApBY5PCb7a4peJlef0Y5ShdT+
bVmavfzhX4mfNUyCGuD6OYc1+z1Ip06mR3EN5v9HtkdFPhDdWwxS+3lQgjYj
Y5VmK7put0qedzE5Zacy79tXSXq9dYvIOe+64JNqLGVKpD+sRORb5ryLlxeG
CVrEhXRyP+lhjzRycS0xG1KisTzwyYBWyLzuVYneD8fGjXBQOeXNhd1vxBxP
9Mb23ksJv1Puw00A+5M2ygnbZJthgI9b/A1lL5wPMvKuSAdkrneK1veIPgO4
98rAfjqH/PelaVJBLIkQobc/WLRMhOgVw88scSQ6vYKpNrHr8mM+sfC9IawL
zbphpk3+G0/3Ejj9MZc91z3e69dDLcANyV3l6fE0zY1dR6XzbD8lvz/vsqlp
+fvVQIVx2QhZUInCn2oQm2rvZ2wHqZd0nwha3kordJLVCp09SLygDjIlwKVG
E/ULN3mCT5grfHhBRxi2uiI9iMG5DAIVXgkGl9dfY7nFd2qd46RcK/MWwzFC
ZG77Ngf+NWyBvnqimjNpuoKyrpP3z3F375UeCc/hCdtuZIWCVkMgMKdhB5ok
QvcwBDEk2oPpxwI6CuC9klgOKZGuHFHzhljF/3e2UMEQL8gclpbdfaL3kcOc
U4VHHNjdO7LSM9W7owrT5nuVvJ5rb5gdr0mVScX36Z2J3RFwoxZ0kSGfjFqL
WLJP8xG2GYzjhqwK8AbI21OiBoERcuiV+N0O7aBiVNjlPjJveeeQ98pTAtVe
VlqtXveL7FH9I3YvxD2CWNG53KGboHmD1T+FDGy2lrzFtkWcDbYqipw/ayuz
E3xCiLdGXQPuV5LJAlC83qlCf57Bo3J+s/dMBP68ptOmI2/gvmn1FxjUeCi0
XPG2gmyk/eDNitikP9vKGrNV0Af5snVRf+4nM4GdLRzWhUvqlif1Zx6zDM8Q
cLJkmNkPHNP7NWXmvYtIqZr18miNMTCa/Q1Ca5SYlUX51nJrzpSLoiM6Zl5O
4+8WO/e9UZFPkps/jT2LvcLpEKZEIeBOprLxVHnlsAbo9vUMti7mAR6JWgvj
hZQKzXXtOC4M4wwMBmURFLGadSanL8FcqKKXo2Wxk7u15sGeyoM2E/f1WvW/
vtIW5fGkLs5WgWNEJMPTjjw4NPNO+4fDwgx288HLysLqHWy0PImqamC0scwK
/2KXKqNUl4Ov33AEBuE9po1JlGYpcT9hSsEGsO5CFxKDdf4RiVGiFh0eb63k
zmk9r/KJJotLEojDegRLqJE7BJEInp2rKj8DH8ptzPMAgk4Nr/3yZrv3wjMb
fj8wQQm4I2JOlvWuinzl2X2LAVewHnKLS2bN/S+TSLJ967KGIlsdLC14FjAI
XOwtkfsjfm77m3b4SxB6/K6lXFYPUKyXCZ6E4C1N3w85dPWH6wlsGLBvv5Ma
Rqky2RrKIgUb48NXUgobTMRLHU96qmvO8Ikrw4a2Sr2m3LOs6ilAyfw2yoJ+
37FKu00Jotz7SQ6eqk2h41Bh1Ku748x39HHIxt+kwTv2cvbeyksUFnULOp/r
hYsgUBgSFoqSpPq88DI4qtE40HJbLEMJTd4pbShs4TE4OXDTY4Lx7l+Tpd7p
0tDFTafoupc21ZK8yZN5JwYhk8oz9EzsX3qnlHg+lAUvaV7T+oxHjgRIoflF
KBZffcl7WTyENLUzXN4bGOi1w6dUlaVbDq28SE7keUvYsv3fE+52a8ugwNV9
/QYEBgOcNZV/gwql7qSfNN7ymOJzcZYf64+66IOZcvBNQvGcNofHV2ewyp2s
noYChkEr5oqQOJwHibh8Vz3YnxZLa+p9PmjG4Zhg6GKQ+QRTzUON/gjDK08N
V2TBg2q0/inwk78ZgGECkac8xzZ/1ZjOa1qVd6AzDNz8pPLhlvLY77RgH0Bs
A6cA9gnKs3aJdrZJd9+11V5SG92veun7KToTFJEdMpwszMVJXIHmiiEt+WlM
F03lvaH9Nks5o6HCmmKmmk6HUQV0PYOXrIJ6hcRkFSVxc8NWloYtecfCBud0
cRAYPdNxZc5gbD5YCTLY4F808iM1uySO4IazGqfjZ8PhF7uTM40iraPVTYsF
basdiMNXdtWxT9pQMYQ/6jWdH6mPYbr1+9T3zRz1QeVVKlHdzkSvoSg/NXU0
REP3gPU4DlyiaAITf1tNxP5/eRcVJ+ByR3u0zNw1AsGbakYg9B5dlWRXd/2c
MM3vcBKiSNa6YA9MDLszmyBzkjdD1KTvD1023XbkSt+5BaVpspvapJy7NDOe
ol6BArZbHcbsmW9iMBlSvK8Kl8jYBck/3KHG4tgm4WdvGV8qY57hjJAMTUUH
/QjwwOZ0JGSuXlH8D2SJvRZiwwoDgsWZKH70FVjduiuRX9JY0CzgWTrwQJjL
l8B20NaiYS7HJadW6NrE5LWc8ROkE+SynDYLxB+rMvE19FOV6yVjK0cazDXp
/iCtZLS1U9RN+SsH56iY18bv14sWGZmyeCnUFDc3TEtLeg8qymD3LuI3JuCd
OAsCPVklM/LNwJnGl7i9zQcY0Qj+W/zSk+65BMkc63xriyPUMBVxdgcUKfsD
DqvZPRVRTPFZTNKPoOzMrsRQ3lEkoyybcMvqwzKAZHTXV6hurX+fMco/yK0/
cUyWbPWB0wTCn7VfaBOxcGNC2Y+267W1UWgsYbOWaJI6SV8oU50HrOWOvpxU
4B4oj6VjohF4zXlvHoe1MdgpMOGtqSH+5E5pxBC5/4M/HdEiKUm47wno1MgJ
G7zXLTCT7Kx7DAk6c/ByqIU9+UdgSy4bTVFsB+i70oRpHv4Nzseqhziqm2D1
czkI7+qqAE+qA65aZO1/zIX2HXKpDdqhaabnm2YQCLf/LLVFYgvrDXHmHVFE
CwfVnoTT6j+zN4sr25ahlgDwWrY5W1H7V8mjDBdW4/NmIbcM32/9Sw/AyZw8
drmPcV9qyB8AyiPOFtDKUvxigvbe5IlEBY0cjxZ3QhB9rJl+RFdFACqcAQCx
0x9seUEStPh5imYXzT7y3fduYjFqYnhxgXScbaH4X3zpnZ7XwH9DPwzQnN/a
Gj81clqM4YOjgk8tYDogqbPFHzqbnIQPC9Q14gJYStv2rFBKqOaMadpDjEKn
PA8S3eXEP1yK6PIUviY0F2LX6RNCUlQhTG2CF3xEg8JzUJjln1nlZ83FQVkD
kJfe7i4jW0ebG+wMW6LND5lKIgja6VNLf2aXFDGJ/frZ4nn6wSsWMZoiKCwN
6VVFnK9TV0kBYLFdTHkUuyJzgL/2aMasHAI9M5Ae9tPuC3UlR2L7wtwYKsLs
1cQXNyqaZ20nwmhM5jkz35KOfNZSut4hShSWkaVpXgpQAPOtF+SIies7jtJi
1ijfvdFpSJe/Nj+9BerjDGheN3NFrLs0kSaM08AGO7dbeVqzlV/GdNQbU/LJ
k9b7Ob+EQ5CKZHFiA5e6LKb8bUqB9qyytr+CXkOOX4Xh63Aqt6NlHEdwNgqw
lStpIuOoICI12BK7j0uKfLcJaWeBKrovOfJgI/08KHVj3/IR9WWRpI2RmFno
oUhjN/8+WDh1fbbScEBcZBYl7GG+bhoGyRRXpgRUvop+B62++xhfqGhNOHfs
4STqHaK0eXaIELT3PIPOeAmmVsJ6GiKUGZN0duFdqgb5JG9f8noR4v1VWrrj
9lSH4d5+cSHb1oH9Kzd3s+53pgXMcL8F0FA5iEvLiyy80VQIfiL6T0BXGIng
39GKfkvMCA+Rf7zG3iOrh7kWe5+cm8HCZXYEqDCbTAg5anTHeToZ7zALoyQ+
jzJqoMYvS/fl5c+YtK3+Nu4KcrY8tS0vlRacGbhEKhrSAXT9Pk1Y6JHKVyzh
oe+gtlPR1I/dx3+RFkXcByBDMWEVBlT9yH7I1U50tnpisaXNYG5HbqTQkjkj
hTvI+cxgaB7sRf9n9fhxZGMTo1Soi2iIj2n+KFbJi1nW86Wn4oyrfHXCy0dJ
AEeDcb2pFpEsSlhwwbfgAHmZgVvE+0kUHO5Zobti0E+OLbOnXT47NTYKndpO
C+l58KRHNFh7IwrUPwbhbqeYJRDy2pQttE3XYXQ4m40m8cXJHKcaVGa0ozQx
2kBU2pvII+1UGQS7BiDebjG/4qdhj7MaOk3ucHNNsymW2SkCNPxsQjT2IwqA
qBciwfSDCOhvDrfUhYHvNqsBNdlp6kerE2wPQJxexYfR/vUTbj+gR/7+Jx08
uZtjx8aIeYpLXpXGoR2VLUjurV3RMR3BLT0xt6bc55AgkHx7g7jBJqVw216+
P3Vi8dzC+wDlvGkGd6NYVE1p1uuNscjjbex9KyATV9cLWkusX0gUtVXSo/cY
mFVacDVXt6l9IERf6rOuWLYv4bqZn47jHpu9xYiUE5xFGt60DCR0YKG47gvo
H+4LimznOoSbI7BsHsfgVKRbDcebFxLiKhu/m/JE8PrsKjgV3cIORwk8SfTp
UZgntLCAgPS+iMM3maF5lt419bcKrRPyiZy8utqpdCF8sVznoMJm++qZLWhB
t0YuHgcjj+txb6UAM6pGvWsPQBNJUeYGwhfM/RaiHKvqgjnAhvHAdNJMz9aQ
0MqhmQtKjeomR7M3d/xJoYZ9Npa2wX8os1IaFnYeOT8gMcb3PSO0Nm/1Ga8u
4pshk8ReFQI80LTJZX6571S40bv+aHKNvhvkIOkMlewzzhgt6idAGJDvMd4o
pnhIHr9POzgRRiyJvfdlJ93EZ5sGD7jE2AeXB2Jks9jS8amoaFnXmOhMDLqU
azGrQfODi9KATrQcdQDpgZdoZmj5x/hC4tiId79qsToLf8uB3dO2aytodAjT
OCNcOlciZqiZewwqpodtLrL1HXXhmUBi69btW+cl6ClH2B78b/KlXPw/YHtp
gO/IajfY8DMjyezHdtpc1+UAbqe71pP77YwhaRJFfywCIRmi3yLJIUAYTL6g
1X88Jl4wBKbkahdqwH2cz2UN8ZBUQZQoEXYJuFC0Lcf9lbxuX42I86RjIZiU
ZThvYLvqURZ4bzIHUV5xgY09h4r0cruKva4S2Q2WvAo+ycdS3gmD1wmzdNr3
pU5XX+VJXOi8OqDBUqOf7SPyrolMcPqoR94ZIQIt3ppMQNzwseblO/iDyAor
bLtx4C23uBmcEmG7ZVrm6m3RhNU/7m9LzPDRjb8nmdx6vH5rtcRcvjh2dBVf
ZYiWup+njOgvBQ8JPHE8Ue04m60JaAuFhSXXgz4RCPJXyJ1OqMeGBj57FlIa
AKoEFkGEbSYpYX0joLBqdigjsPqF8sgY9G0ZRR9oRutYeoxjn5loWE1i6SZ+
863k1V0Xtaa9CyG3fBuIfgnfn+y9RuAe9BlSPMrBf2w3WmWNjsarwzKF1912
RMjv+F6JePA3470Nk+KBBGlNAh6L0J23NzDLoHdNk7PQL8EYGEJAcTu+nZOY
DuRIvEK2akjS2rLEIk+9QZK5lGxzx1YQlOGW9Rr+gz9UrqQIGIVn+tx2mSxE
YpvR6to1qb+gaCOvwskz/rvAXjFjhJZpYrGKQ4uKzf3RVE+wJwc0tNwFd+EL
PGxoRGqmsXbLFl1x+e4SwzTnaQ5mNX409YnbQtC8NnwSLeVP27xL+KD4Z+n+
7YcEE/JV2A0uyGdWwHUc5W3JsB9S9RzZL+X+ezsX8hid6+c38yHvYZjCn1wq
K0lwME1gSg6E6aiQQ7ksABa0gGCCH692eihYrT9Lz7nq3mnF+pB8az9Lpgkj
6JJswVikD4Ap4lMCWaJb5IeHUP1CxAPg/EIRrD4vekdZR727AgUjT6Vfc/WP
qJwZAcCS1RyXKSfmtDCu5HeL5BrkXupewbM/ZaTyYqj4AFG+gqhFgoOPt56y
G1h/UAgkzE5I3gaqwEbi82h7Zfc+Pdp81SH5wIKVSYMsWeYu4/iSehHnqHjj
FfUCGjUnxN96Ora9SoYC9p3aQiq03XzSopC+k5b2JMODsr+GML3MPy9sj9kJ
Di1bPCjKp0nslkxDmXkYv7owaacnWQW+1eMVBpoBo1WrXiF0kbrDKyeSqGYO
agakcIliyafVOywP3p62K4d0Eh7qhEWtm7zD/iwlqYlRATj3RkcBno/BbsoY
A+tup3wL/iLFcbzJu0hacipcvrcAq3fjq1iX7hkPrbu77g6KIJZ7svjnlybq
aVfGj66zJM698ILnPnWeU8Gmm0rXt3qWJJQi54ImVL8O/ewZp9vRxfMeGqg2
szp7qmfQrIrs7ehYEZiuiMb97C7KY9R1pt6P60JbSQ9g0Z/58qIh520lsbxh
CbHB59IrsSZnnzwfy2xLX4mszgs5EjONCxBQo2Cx8F+rHMZxtRcNsFnl/xzd
M1qtJ+i74QAivl9OjI28iVQfX5yuILInkVN8MrDVWE+KaQInn4dM0bH4Sl1L
ARdCXhwjOOw9dVLZSIxvx4JBmpqMhJDXm/KYMbMMyeishfenOade2O/sx8rP
aBlxIWILxWT4q1E3aC2co+nZq0lVED41Hk8F8jaQtkB4omU3ZccnuuuOmUW+
DwzPEaTnoiOuHpJ4/cnebnsZuvGFim6NR1vKFIOqPRbZmhChElcZ+5bfEtNi
SLWcJFjPmRYJi3xwFYoKpKKCjTQgzuVEDW5pgH45ymeQd7GnBzoKkX2c75j5
1kn1XxJ5ncVImsP2P5FIz2fKPUbWISOkyqGXA0k6B4fDLXJE7kLAkKk3s9T8
M6zhvbfAxb8KqUZ6G1TRaYHTzXQzO4dnBD2cT0yBnHfB2THBL84h0HUBng0g
yLID2nLJI4+B/lVUxA5z9pNPyKY3IPP+qmPUs8FS80xEOInJuunlthgMNLpy
TAMKdKZxpUh7vasAdhATUUapqodwBS3pyH7a8P1Vj/nZ3wMeDlpSLM13yPZk
Xk/PeI3baH/G52gQhSDt7j7IOpt9jmfiFoROHovCSsTFm6K3UP6gMDO7pQzS
xviGnJ2RBPOZKNhqD+hQA7spNmx4Y4T6qrvNFL1yhKZ8JEemF4fqNdJhMatr
g+XLJNAp6MHLB+UFDzNhzsukLVVTd7wf7hkdOlmrJsOdfmoBiOxA4g9ORq5g
ym7zQIhJvWd0M9qFY59g6+Ck1Dy5OJbX5+4ARB/w29JVF9vN0h68tHWu4QdT
XedT9fwhNcMyxW5lNeW6bcJbG0YZYsrJ4MlM4hp4jU/nhs93bP+xQCDh3UiP
xlQJV31WmFE7jT0NpATXXUfXjwJFXRRNvfHJWyVKg3zpixvZUEq6qSBCX5KH
lF+Rwl2UtMnL2XzW7pb+S4AmbrXKzGOVaDTJV27BzJW9CzPUzYZnPeptgwcB
ofhXwGrOt4DCgi6YaVI0q31BMCo5ResjTOzAYHZe8Pm5TvYcdr8u25UPP6xQ
b7gH44d2w07RjRavchF8BbQ1UCnBVaLoKSTTYt7AfVX3G3gsT3cki7C2jroE
papcNqS7uRNh8j9FrW/ux+0tapxf9+n1kzWj3KLxj98ePgw5vfmHFqHR6Kl8
5XZRsd3ZniT5beWGhXsoRX8XeH9UCgAOL18N0gsYyPtRNwl3e3MSLRm7M3bI
lyq3q1v78f0US/OahUzhfIz7fawW+hUZq4uar3FckUw5OGUjMvrIgJL/8aLA
W+U1mZd31mqnpwAGDRu3p54LX/xfAYlwTZQ0Abcb1knwRQtMgdA6nAg+8reo
Ekk1HI0MKpQFeKjG5T5EXB+wAFFjwBgGwmyCJe+r18tJWN+vvhcCqiGLnEzR
Ojd4VMXBBPZRkGODnfYFVd8sC3xASl5w5lky4e/Fa4xjrRBhFRgB49MOPbBv
jstnP3PA9deJ/bioIEhPqgUA/F6cRXsPOM9cEc4aoNH2gQARaIT1B1e+BsHD
aNd1pq5Lzm2LowmKjjNzOvpMN9njug/2zodu4Mmbnwse7dnodPKV/dHfrzaN
XsgkCPAliS1elMoQNlCkXIB84r0GrtKOvlEaz8s2riF2C9qurIy8FgV6Za0y
bZvsyCtePERnjvDyISCW9EgC3eSlqf/s9UQURu9lS3QohaoYZOCXWvk3BBtf
DEttj04yaJ33WCHlR1KaUu8Zodf+8kW1F3RrE6Fra4SmhZ//DcgGMGO677Qc
kHJq75j6UITnRlHa29v6CS7OcQixc21Jj0F85mvP41F9BQpnNoykyrJ/3N3O
lOHY7mo3mzbJaBtat7FGHLDxSob7RYcMs6s4UX4wFO+Khh8IrNUA/a+opQhk
CzswmePiAf18VWAXg5LCZVIn3x3NhUCt+YxXTh46duhuJETQukhUJDpo7F+s
BEcgHuv0N8tiYW2EomxoNkYn5wf6Piw2GOsf0stMYkXAZzSO76K00sMUKtlo
n2K59Ojntoqg1FM6sCAC6F7I0Z3ubVOs24oqU1ycdvSjictuhZKhDIjhZ5Zr
dkNdA8tGsMoZdMaGAikc2SQvorYPKZkwwT5eiRmCTG/8ny2wb8AB+Nn82lh7
7AkXmfjCYBkhogJ50Hl8/v+vc900uYJTQoKwfv9sTKtlA1m47/Y0pRE5hkaG
boKSeX9j5QNyxCfZzJ7zRVSaqGi1kpWaU2RWT0OYekMMjW+vzWdoT0gHlrPC
I/bKXCAIyKz1BRfxWVbeW6BKnyri7ncaEFTUcqaGKYlqubPRcHmlbprwIMOr
I104YmrLrIL4v+m8Q+LTbJRh40YEzhfldz5VMlI7HfR5mMvol9VcMKkkmKY2
h1TSQwZApHUlCwYcNIolNDk/mL8ghFWi4X9PEPKuyQvt9QweIHCSzL7WK0YH
ooe3KI/cl+NGmTX7cdgrDK2GAQ/SU62kk08gjTBbfJhlSgjL5hrylo/0kw6m
AC15sVODTDJXYFrsWBwudTTK/2Eq3wx+EFOMVaw+1dVLE+WIS0hoMye0zme4
G9HNxseFTT8RwwBLOTqnWqJucPW3huTz8jN+dnZBIctneEoPFLvSDeoMI8Rp
nYzqdNaM/JpGCGscPT0rc4vqMZLJxOVcWvUZHjR5FF2QfBLsJFFB3dAs0h+9
O09tryf35t+JxZ/7AHCZToDuCf3U21P2x6iftUjQQOYluI4fp9jRWDF1FkA8
nbuqsQgS9O0KQ2p4ECJWgD/h8jQdRjS8MniFDrA67E0nLKanu+B0dh8uH5fB
xo3GLtmF7bfj7Vt/Ad+MBMHi4afGxOS+JVlKnpgktPv5Ln6TNXBQwgdYYef6
GqR5chd1WVn/GmWHuiXqgp3KpAENY4Vjtc4+jKS6tuANK/3pujObRMbU8H/5
C101L07oTILqFaYDYHDxwxIdhD6cJHpe1zICyUZQrO6DRprMK2BzvObWxMke
15EJpV7VRG+3UtqJiS+G2QQl/b0D8esyqDScb+4u9OQ4Mb0q+Lf3HqCrun71
EySNnemky/V6sRASx976aoc94HFvV7gQ4NLcbyJH1PvDUdFfv5WzlpCs4Yrm
qjRHtCMcafDLvRBT0T3N+OWXxi5P2JukbA6/shJ8lN/xejWcXsS0L9QHusI5
5w0j7OKLCQppCUYeeafa0gY+AMWL52gjmRyho9rXkSMpElfXg/iYAMnfDnQn
RdFsnvm9ARkfVVNkbfD/wYInGB4LStv5yCa5Lb4C/m6UaTAJh8aXgfrpEnWd
YfhRYzQpVxeU7dZmxyelHhvqwzQmo+Fd2fRgAqghgaB1xX8LUn8O0OtzuzY2
Xaa59P4mJgagTENJOlghXE/taE187UJjwOu61Df8BGjdF3V8TByUILzutHPg
oIsbpizmcyeP4md1WeXsNOKaBFsxpAdXzigzCCRp4OlFVVoL/JaxLnUbwww2
Abb6tvyIHFGct8G1v9Axuzmkoj775KJWIEgnmMZ21P88pNvy5TxlvQtxsdH/
n7WbLcVZ/hKOWh70FeALxYmjTWlQ/LtdoF7yhuhvbgDvxHSeHMXCGmUxa1a5
6WDVMLUBb3irSiFGb11ieyiZ4vbJ96/H8HNFUTlkBhfHaOEaeQWK6n705gyF
aSwJCg10SDL87SeCXSOBPzg1uBuo4KpoSMI+kH6yUHIU8DJUANA0NXKlreHc
OKhvN1LzctfG9Wamrb4MOo3pQGnjZGIwD7tCPszUWCK0PwkgDeNNBPy0DCjw
1rk0j9rakVU+01EnrupxFKcAElYQ6NfhDt0shQpcT2Sazm1bDvfkPAH9j0jp
/4sD48d+wz9Sqb1U2UMExKzzOC0cELSs/P6x1afxomKsPdoYBO8s+tJzi42z
xxdJCMg+jWtuAuF0wcjIrOdxCuEimy89fk9pA4t5JzVi3YgPsKv9ZdCt5WU/
P308x/VbteforsjuAwUjUS7LNaZAEVu0adpO2vAfigOyzr1dZojfGuWlK71b
C9IYXRxbamwkmxE/K/+c2+vS/lLy6EuzGZtl0MaIWWNrwfS8zRvGz6xRpYsR
gX0IIQ1THqjL7dZQ1pBQNLRnpUlAhMPPbuyJgSRnVfLeDbDdALIcMM1NNsVU
hETE8eoRtxxiNqjY6f6jrJG5weEZX2HZjvko40LNWVTeFTc6BfIkQZcSxg4T
VVNhrqqXeZoHK8uFqr8vD39nhkKVu8TVZ3BwbJ/iTuNNjuRCuRAyXExju3Hm
gca4a0hTYSGVDd82Rcgis0YMKQljXO8viPVBB2MjstOPg435BvDS82ofU3ig
XdYxMreBUSXWBlQ9KrYYSkDdUfB4V7YGkiMPKsoyJ23OUNHfKUHvmj03VJJR
PDS82OYEF6Snj4FC0z8u+nhZm04Y2Yss27DE3L6Oq2y5/bEUlNC4mccKxcLD
fOg18rQYjbCPzES9LfS27BlPO3uOgT1tYNBgfkDyG3zEo4d8JEVGNDe5bB97
Kx0yRWjypS6i64gUXtoTr7HxlPxD87IvVdYbA88sfjf/adUg/W//WxRl4UFK
fSbXibdj3oCkD4OkUEIDvkpQ2JRBGlqWi0dBd+5t5Kfvo4EcaPd7FlAZg4PF
6lXoNUNbHUGBYSiE/DGRZt2fk6KidY7ZmjO476HtOoD12Wj8R8fbjNb0x4ti
SoaipKxKxk3ESYzTtYm7GSJqQXiDoMS6MYLnS8y9B0qPUxTJBNvx7yRnj6y0
7biXJgd/ULYv4qa/G4FRXSz3kpu75wx2t3Qj7iJ3r2aP9nA0EQN8IUxXQ9Us
5e32dt/naU4Q4Qz8ECTE10rPOqoHz1WnXjO/nek2xK7XHy3SPBxQ7KKq2v3b
nwFxzJ02XNkHJHgtyAQZwrfVze0TE7rmlLDqtL8tS6yGCW8WE8Rw95twSzBW
Ve6aDtCa5uaTWcyq7LqJBQat9jPMpuYNCAXk9NwRRanQOYAeWUay4OQzSdD0
qtl1ayvsbI5ltC8L0MgLWEvQgnkRDTF2+poiX6wK3jvUC60nZU3Q7UxjAhgK
CV4qPNXm97OpLwoI8UCb/GCREklEfJ79fcEQTJB4vubtXcKU1m1Tzies8K0f
EcM57qgd96NW/tPgbot8mK6Gs97c0R5+4yWWyBrZRLixN3h8zzAHoHYHYJBM
Vg0W69sKY+BGXzkMe1CDGVN03fkZOyPfVbtRA1cXWZA0CDOGVYHlF7tLt86N
610Yxkn4UTj/jIJls1eCag0A9tsMUGaHI7BkkXPQHCzKqvyaDbhc+nBYPAT4
traDFJNQvcnfN8QurUdNarfv0CTM8HtxLBde0nij72F82mPIPKvxR3KFH/L2
aRqNh9EvRd8/fdn2eoEZNdTIVNwoGHFdp/QqnuiMULiz8mIrbaEvu+4JxrYV
gwgSb4HJgP/ETS5QCiZEQaqA9oFiwK8Qa/CPIFCMQSJb15faokNC6zB1/FrY
5Vrnpa0VJeGHzlbkJolYUM9ffvTLvPSWKEGvEFAO1WSl2g/JH/DkGdhSI+v3
5nmCzL0Gd25HFqUtMwZ9hnRebQDGDHimwSBlBBiG3ZUyJfVdLyU59nTJGjXJ
s5lC6rtR0h2WONPtQ+I+Y//LGxv1aagTbvp+IVcu7aojLwrwZtqLTk4zhp1G
gxKlBvLymAFDT70ctjcN/hENHf8iVtGkDaccKzJ7nXkP0h8abeHdimXpzQQ4
Gu2yCEck35IcLPLVXnhCpZyTX1Z3Q6vADJe272cPr8shicCjGdFOLbHUm//v
CHzvm2PDViHVytp2uY9fTJDK7Bvh0KVqkrW027LYOyW1rbQta992lr9MFBZc
UUwN1Ua19VMF6qCg6eGZteKGKTzv0q+8PrExPmU3NJJbyaqJStEYb3/F52Gx
4LachRKJGkXZSewj3GuK3BnNim4aUajBVxyDD354IsfrrNbkrZa/pqwsD174
2miHUfVzX7/ZTmm+h9CQGfkeLyy34NQsBuWQJN4dOdE5jRZPmIUi8YIvYfHM
wwnZbsFu2jeOJl9r4n5cLSXApMlU7uYAlXTik2XqptGEQDZbOtn55iDWRr4l
5HXO90VFp9MEsjIOagw3+g9/qt7bSHfWr1MSh8BbRrE8VhL2wpm9LLp+mg4w
zaLc8+znHoqe2JruM1wTDo7EKQvcB0+8SIOB9RmU7sFhXSY8Nf2CoDXnZqly
2+bnoFnNj4rl0LJZHMW1OjmzcsB9vRYi5clQkdSJsHSaUIvFi/XhuIS9JXyL
Qo+jqjBqrm2+yEOsAcuwcXDplTZuaIdPJP14Rd1Hi9ldxH2aquDM3DJ/tHBH
pB3UF0zmAmFRaPI5OXQ7kE5odMMT5O7vA230oJ3JkflVIeZbhMmjmhw2Blnm
Nj1aMBmd7Lx29dpRy883FiAB63PM0XVhPqRy1B6/oJi32aAgLbeuWkvxCcS/
DlU4+4Xh/zlKpjglie2fpNUozftQKWUn3BaXFfBhuhEbE8BHDI4ecU5/nHGQ
GCLyc9Hea9Pia8G2BMqii8/i/XOIzNuQselbokIkwKI3tql0ValYtPeYuHsN
dAxOaBcrn/w0y3SN0DOuRtQZhfcoJndLiR8zoGrSR/WQ8IVhX/NQW1Oe0yed
vRyWZTu2ydDVn9GMR7TlHaJK8x8pXY1uyEOGG6NsmQ3dZBKz/DhrPoObHKyI
f42IXdr5e6n5UvwWD6xmSTT++32WBhx+DNy00qIZLT9ZZd5ETqZDgiZgU5G4
+2GxpbVlf2np9XkV8KD76dyYzThcfYIxr2+8gy/oSs+IojA21VVdu/Nozcmt
Da/WEEXLIL8qZJZsCet7VqWjENujj8AMmPJNfbgaQlcKhrlQbx74KgnS4imK
ZM0W8fVUgs+xm/esaaDg9VdqRqtWSXNoh5FuLSVIK+HkylivtNi7bFglD7NC
r3kYWLhU1PIhwoIz3t8byh77/lTaPwkMsWa54ooL4u/ChRaDbq/Is1l3q+wV
Q3AgFX0WUvi+ywaAupWuCAdHKCH/aGW2cIGZ9AyTCsOyDkNoLoWi9U8Xkymt
hWijGPUtZ3qSLOAZlAEEq/FMeJkMuvdncXPY0YVhGmHAUv0HdbTZ4aeX9YR5
DtA4WQRFf3aFaWBFy/BpSMEiuHqR/joYzCUD2+ipgCQr0igE2gqr8btxhKl7
7e+2x40VCFWkTFsBQVhMxFiR8NNimYt8TwGmBYT9jlV/6rLNryehZ+ryj3uC
3W7Bn6wdsU3OWlvla5N0yabpdEV+9OAzXUyDuO5QxwWUrFyokbWVhFjn63LO
2jhhTiaH0U3+hGBjvUabLn5dF/3rU8EdgLDDDh9Y1sSbRwQpyGdT74eHiAYk
IRcLry3MC3GiIBsJ8tOKuyCBbYfO0UB1nL9Opks461NzsXXslb2bwHcpat8I
vcZuo7otqkHyE8as3716RtIGVsE/qqso1ikx2OisLOIjEii3SPIVEZzM1rhp
xf6f5zaIuTOvsyVQagjp2ay9kWMxHis9OB7DAqaF8319ac8yLABb7eQgmcJb
HSqjyrnx4Tn++Hru3YArnIV86/Y7OIpFCDDILVfFSvztMcK/yKctQ2xEHLw+
PQy6uOAJapY3PKYbWyzidlXym4ocqyjZtDHqM91/r+Yjuc7fZVND3OpTJ6lB
DCGoGrwkXZTuVkly3yfN05V+DEH5Lx1eT+DubMHvbofT/DbNrbOO/5ax72eJ
lDiHnDeRX1hsWMMtqlcck2sSiFmWYRqueu3uJuyVuaB39GSG2GhX/bfJB9MB
JpKgvysip6qCI4hF8yPbQ8dTYXfgXhfQ8/Ud6y2we3KlxrHzmiANwUp/Ffkh
KqfPb6w5z5/N57T0cay7Ucus7LLeERPk1HgNUSceuuWnHG1dcivjIpk1Qdzq
GSHYrdhJ3cDHnjTHauktES8XDigdtgfj2WDeAO67hvDYypP5C2WK3LnEbNhU
6mHcyuUx+wuh9kn0mdAKmzhiWnS2hBGP3fkWIsKVXJjlKIBvuceTsPCZoBYd
VhfVliYzQ52uui5ei8+RUkHAl/7GaXlegnUOpiZiDrErzGRurg13dzkq5/A9
56NJpbUFb5t70eGqoivcMgS/6VgUhXa+Xqd1TdvRsxYqATzDzlCcMAU2VZ4V
bfsdd/rR1cH9yTcPSYtVP0UUK+OG8tHqQVHIjBRKbeBpl9kGZ1ncR/+yaXlj
e7y4nbRJCizWswxuoLYLG2YbpvCcAg0hNpIAi0jhLTFdZ2QCCBIMJ6DA2TOV
mU6Z2nEARmSRi14n4nN3vphw+/eS1XDCvcn+y+IHYaqNxuxuwUJuPyiHrCl7
NMBOPEeBbfkOU8L+YpT0+OOzSobJ2C5ai6Fqmqi8kXvMkSDc8VPLXSTVKU5t
4VCa/f45sFq5s2V9pAQW67IbqKmg03uSh7JmVFgyNud67DO7VQ4xYQsQuqMP
+fZAgGeICjK+jTVRfq/jhEZ0KrJgcDtEgRC7Yt61CM2YVDft8gA8wO95AO+S
0t0TOxmtU8Qn8uOv1I81xx4CoBYmhMAh6IpVIOJXYyGZh5tnFUZoGH3Gu2PW
pV4jxP+hw1vDZcAz+df8wNNC22Ou/qI+zRw9Bk7J25x1xf/21PwMEcHiGTJ0
o18CUYc0Ki3C7JF0LwbIWIC5W7mfFRoK7w5eMkTHPx/Z6dflQzTz2w2YAbrG
PAMgeJPgvgG1GBLHrLKV/fM7uTJbyhdPP5ZYRgPWiaD7cWYT1S/j50I4bxzs
W28mWSSjcO/R2u1afBDtlbBEKTtPcRJl61z0+0fFJ/p2rY1ML3OTbVLbhnT3
SCl8oDdgHqXEzyg5uaO9RjPPHaraXZJoNt8mAZ09rUj1R4DB0iDN36Bgg8dI
/Z/4TsnVnOn9+Ma3DNszkbyEUyQP/3BJbQJVS78jNFZ7vCyNtVYjvgsgAy1r
kS+qWvPfmBt7rTlH/iKVpSlZykNS+ulJTMjI1jcaDsvf6JVZsCZlMeN5vnAE
EK5RFKbJJTQx7Qs5EmEyP6SPJ8vVtFZUHPLVqrJJJ6TyvN0rJJ7G6h5xrvg7
+ER1n7Dn0Gs1n6riqo5NUqHEM5PuEtDvxB5cqk4ACX8BMQDi/2jiDk0DN0rf
hUkLFZ3DnKjBW2d2mUDi39NlGgbJ8crmniAzuyemmSbbPuvFzxmixWp+Lwbl
0ckhd4qGNCh8eBbFX8JhiLZ5bNjwIkB28HHJzCCRDh0/EifmYD0wpK3iAaeh
ronNbLgR6ahBE7sYn/yaswegGks/dVGIoUp23czm1X8xJdVOmpmDb20x4Zlj
9h5gtOFU9720z3I0/SiyvewftPQtXXiflokcNmkav3OT8j73NktswhkgHu9l
jnmRVGTnY0nqqK4k06yxlqY6Z4+EWZs9tkGVIGLlz05puW3H68i9ZYTAk6U5
cCRn09GzAt2UDHPWRtxIDegk5l4TTxa+MR18tHQKigDSbUXe0VkhQAO+K4Uy
Tx5SrkLAS8UnhmMciLhyBgeYMPIhlOvFI2ypUomEqJZS0jGuivtiJbYELA7o
BtEcb75yu6iMoM/c7zGnKyWVUGnAYA7REB/lx7V6zMFCxUnyeRnUTnb2wQrw
JzrECHrmZayH+TJBR/E0eanuihUHs2GpLoHQBPZQivw8FnWAFSSF6hhbDjbI
bJjEZZy8FxJrdqbBy2P42MNNrmYruVVtbWyLfT6fa9wPrgAP6ErSu8AdBzQ1
uXz2Kqxzd9nQ19+1wAlEKZySww2QouSv26CoEmKgVKnxD2yefWd0YplaCZyB
NX4zbx61vsTRwnumN7in8jl9+jfD3p7A1TbpeBuIFEbFfb1zDBE47y6t3Ars
aY/UPOojd5rgc8qjCt11XVascgoBMDQCfvhlrA/Otpy83uTCREiMy6oD+S81
GUyZ5TRpvoyTGpZaSu3MW0QwjYSPwu+Caxer5fKzrlFsNSNoeY1t2V5aCDDF
xRDsL/Cnvmf2CVoDz0x3P/HhhoGGMG+z7LjbZBs3c5EY2EsKJcIYgOtBjhxC
22nRErgl3q+Vcg3rDzDUyUDDlp4jGqOSzHFQfsKIkgYIVtSGjevTD61gzK5S
QLmL//n961tVbU8giGA7WEOObqkDFlYJz8f01IbRECdpqx9ns+jxQZHDcT+X
2L+Ichpp/Xljp6cAX+n1lf5jWIKnbJ5q/2X2t6FhwsxPiymrmNeWsT84gGgs
yLLon8+PfVvY25TBhVKDCA1g9ClNMXTP/ZYKRzAqguzsVPiQkSW7r1nKkki0
v9TMNsPvlQ9Q9sLfdW5YqoghVK1Lly6N29d4dGHlOt5hOY4odXZBdbw4s/mx
/zp/V9mg1MQ7xrvUC0mMeJq/wO8Oqb3tNtTjnid0viLy4kfiapxGf1rlhCYr
TEnnG1UvYR9HmYMU8AC88jJXdkuqzEg0Si+DaU1HNbwMAVQzsQ66BCuatyWc
GvpIlxYiC3viYWI2ZCkUJgv/HL8TrYTqeZNNY8E4oUT+gx+cEq0jJKXAaayI
NAgzyjM8gDwam6F6fj5C2QNvh1kXrTx6yahVYkcJphTCCSQUCiLw0Scg3gaB
BdjEXctIWvOQVSXbwmQcAU6Dp5Ak6PqVrmA1ls+ExuZ5M0U3AcPpl4mwLKUv
4EQSySi9blS/SLyIho63Tf+AQCX7fR0kaRizUQxB0c3pFTKAmjvS1iyHLsog
LxTbPBZqYjLHeABRGqmn1KGYhI/N6oFT4GziNfbue00e0F6TGSQzpAiqQ53q
ihrHWSSyvZN+MB4eWfqd0/I+RBFTBPcuAOWWRgg+dE9dRzhU/TD0M0Snp/SC
yqeliIvCF+h8PuXReAqA60mkt+bGCHc3DkeTP7XCXg0HGAybeyKaojKlJu6s
D4Qpzqpg/hflLx3ui/f7NnyZAfK7yKJZ0eZcviaf08HfifUMyVh2mSsU0Zj9
WXWcKYbhiZheHmopfN53fy4CVcbqPf+ikyPFv92/xQ/MTZLEQZEnSwcJmUqP
oIyFaqwGd8D50Uez/xbE3wQHuAcQ6+EpX+q6JgsT0OkRavVTwxBp7reSm76k
v5shyNaK1x9CkwvTbFSy97Rd0NsumCtuSJgrwV9sf9qXWKSp12fDZq74b0cd
BTnI8MJ+QgS3Xs5SukrEmIGg6w00JSy3rfPZQXittsbCtEa9rhbpcaLBqrxO
XJcEjLowK8Lp2uqAM/dMfv6Z0Oe/Dy5gy6hEO9QZMeMAqwqfDenbVxAtdBwK
eH/7nK0JMzMFYbVITn6YYXR5cDmuUDVkwAlg02Xx/4ss9uilpyczHQltKVhD
DgDFThtwSvXBk/TxWsBpuWJuAZ+WGw6Ve1WtkuGq1fNfmE+HALrWLRHxQnr3
34x5LiUzbWCEqpYBbP07yVD7FHOSBhpC2uJmgMqmTCAVYzMvy6Sj8ezQJyQp
eQish9s5ggE+QMNWcXvdRAmzkNw3/RlTeqhMfIPhv26bLcp3+4gr6Os/3KYd
cTJ/7ssL4cHq1E7oev50+m243kxIjU2b2Bhi3MNvXI5JQsEN1jay3zmyAZpf
hCCQjIFVuSViu22w6uaH33Z5FDOfTSxMkgYkqwpVa9rBAYm7WHk+kLa9E/uz
semTcgSr2gBVmtNGohHPJ5Zsd3uyZT0BowqwnSOYkntkZuWzc6pTg/BYLMwB
eaehvjZ9p0xTUfIyBIooRilSLMXspWQ5GAKLMsFd1XHgcpwuuqy1J1HeLcdX
vjGeCPnKNXMISQ+wMb5cICPpAIT94Yezhe9rcdg0LNvtMpoiY2g7CCL4vR6F
uqAQhXChWyb++iGg3UF8lvM0cYydr3r60LGIrC3X/6Zr48n//vq279ytT1af
Mr5WIJdl1YSNDTaGFZa/P1aiIjqKdqqRvuyjsGcBnQXNxDLb3r+5HRRiULub
Cw0OGQzd9+/RO4ExP1bizald/v0KSRHA+lLAQCXE9FhMw5BLicVLCmyRragd
vuFewIZU2DBhnWM4b0ldvEW3tJI=

`pragma protect end_protected
