// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
J5v3WChkD2FKsELHT0td8E87IgUxis2oUYLveO/IONSHI5PRLf5LmQ0z+unw7bvN
Clzkjr16LWsf9WlxeJxX3ua904KeL+sn/OF6q310fItKHi/2PoRvc4sMpEqcHO50
M64lPFEc2g5jXydIYMi3FDgocD9riWA7Lo53IVE5B3A=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 50208 )
`pragma protect data_block
rAT491LQEpnfeKrs0/tmzNC9tkQGHx5B8uwfE3JH6nE8FzOCl7KsCbCFB91MVhfL
403Iw5vyNPjOZ8mfJ0EmBmZCeBJP2UzXF/8LWExGWTpSpXF3H/WxIGfAFMrC3pzw
IQAm2EV2J/RA+yrHXF9JTKVbQci1yi45fYVfAOPaGThAu+UIii0a/rNsnewuAeOU
fXmMQK7F2HnGJUNt7ehT4NeqFxjKpBu/9FGUdgTpLO+M+PL+Nn/4m5P32fFlHVwI
sj65eMbVexGNafNTfGcjL8aVaBOL74MFh8mf3u7VCE+ePIabuQgCNHM52v4H1N49
WO22PgPeRR8XwHZN/+3XmXMZVKrcYLEQKZY4UxF3TnbpG6Hzp8loF6/XucRQ5amD
Fka6jy25E+0MDra4yxTvq+kz2to9ncVk8WTTGovbAwTL+ce6MynKQ51h/tHkUPcz
jh9/takesaghwmr2/fCV3yzibcJKY3HP9Ns/Xn3snbo6EdSSHPmA2uouMr7w5p1x
aPS0DVVb8EmwzMyH1yV6DINfVu6nGf+k2MlT95HxipzNnB1t7oEtDaNdW9wTU0Qj
Fj/iqj07z07Jt6SWDz60wp2qivxXbEjhWpAmt1nOP7vHvNcMgXJ5IYZVEKoSDvbU
IVsYlR7i7G+CiSUfbEwQWKQVeygRaxohE9+zg+L++ww3i/EK7XGgrjxnoXcKIx3P
Rz2kCTRiI6CBxVYK0B/3v9Lmp9fhN/U0ybcbhts7KteEltAyHKXakI9+G6TY1Hkr
F+ldh6+uwJL88lkGc9HkhQAFEMkTLcLPjEZUVL8bMsyRzNQklAnqyYIySOK4p5gX
GpwgQzujVbPDqeV74bH8zt1iVCMJ/N6cwaaofTAQsQW8T3SIq/A7seB3K4ar3BlC
vIvJ0w6sBLzR2skg0t+wUjBqf/OyVRQE4JK6mvzpD2qkVisl2ZUgdQurm3nLnk8S
zsPzXubGi2tAFHCiZ8vV59NPPjFtF8eFq+HVdoeRbqfj2SKvlImhYjZA4THVLFQj
yDsgKV2flKBxHBFAktMVGXaHpDB4R3M3s4V0GimQAd5fNsl8Cvg+VGe5h1yQCjL/
rxUKZuQiJ4zbnSdp8JPyArWHUrcKzmPQZJoK+URsjiwEiTu8UAMDVN7wZYD4h6qb
i+iAtD+5l20FZcE4NrqQXD3hK+9US6GcOBvDe8e9plLumqHtIE/gjOja0fsSJIA4
Z3d/TFdQvX9L89ahWqzQalBedcLeabuGq0ZQGGQ91ajnCAuIQAJGALzMys/oyJlt
b+vy5qYoJGhT9dK4tuUa56IrbrvQGNlKq730BuXBF8QERfihkZDu4G8Mz8qKdlxJ
G2vFndMuk/7cRnQLoanq1Sobap/BuVATEC0ZiTYGE5timFFI+YPFGsKz+8je7K9Y
on9ZGnKVlwVMOLfvEmiwys22S1eZeojCuX/sQBSZ3GQCXX2jfra+UzvSSe6eaoFa
c1dX+MhsGa2As6QVNVa12oZcesNAJk2QjAn/Uc/STq2vkVTFL/O2HqT8LAB74Lue
GvZZX16H8tUqDb8TF7ZxEtq9dz1IbaEB5eiSzjE+jd8D+iMJjMEdxzlTBNpWIShS
HNq9CQnT2kDYlM6dQilGn7ZGZyGyam6Jw8gJ71p6uYmtgIlNCKpVqctk2OsDzZHK
3K/yjtQRc59mh7G3Olbi4UnLNsDBnpV87d/Knfow6fcXnJo92re36Q3q4iL3hAnU
94P943EvKeIdTHj+OW1l1dsAhgv7bzviGbYYdNQ19eHTlbeBDvmltBvGFDg8CPCT
mcNWKcUuUwSiABAgiZqrBG8TM2u1yezYX15vZ5vEp7lZK/P9jPhDOKvf6PeAtsuW
GAiF7+rKDdHvPT9E2rQEm8xaOiaAvZuTNTKPLwbZRmkshkuB1zcZJB9a/7Vz9cD4
+ludPjNawTfxCrTP8bAEbzOIaRUJ3dW0kZFEjck2ffTE5AF0mWjp97/InS3EESwd
/y00WPA1ulkbJOrQXErIMqTdr8LcIE3Y3JnniymsakXWSiWgLz2B2GgR0/yobZDh
LIOCeZVrlhVfN+aAezraAUyKyk7kxwRHSA6H7bAzJUAf50ptluaV89QFfG6JXxvR
DaUnrGeGRVTxfYdyCaeiAy+fDkpjRFhgx62HJ0AwXiahh8BNps5Fj9EoEeZWGmqC
bhM9l4o4OUjjwI7pOHn7cBpZXlpHKlqHwRxsemi8GteUULGu3v6UPiVBHnD88Ihl
0DOcly6Ss7tdeyPsIEuozju5VTOd39j7+1CeFqYAEJ6hfZhN0xI1jWSKbZPs3DGe
N8oSifI/aRCGG9WgXMG1VlB8scmG8W9VUAytgd+nrEPPaQI7YBSffaSWaBRJhdWM
9h8fAM55iwjyTWL6Qeoy/YA5sopFbiqLOOo1Ju7FT/zgQHoHHeHhSh0Bhyv4HtIZ
DI4EFZOv7HugcC6O8Cgs35aQuMOYYzD45L+3IJy7Ayd5tj1l0EYPsOxqxNMN5yLL
0CeqaQXkR7rca/eAJkv6+SjbI0Osp+V4a3cigRRU9V5/j9yKsdh+viehoTjztSyR
7KAGTHtVeY5Q4shbn9JcSeKpfCewk0sN/arbD2u2BMMoeXex3eQ3gIaLjS55OYTV
k+ZbIL2X5KioIh0Z2C74KyrTJ200Caa3qrWvHd8bNkONlTzoX7hbNyMpF2ebZVkJ
66z8VLaDGmZy5bifVOoN40XYzKAU40LhADgCGYWR+vvtwf4K2dOz/0m91EJg9iq5
kHk75P3vTNFID16Oca0cpLkb3E7JoAShCg38xJ0k5bdfsuiiSfI0+CLSOc3/Z4JJ
llYskINEccmPbUf97sDTfzbOZwzv2SS4LEvN0qLLv+g5sJ2b0OcrkftUebN1CkEj
Z3yehvZKyfeFNPBZ3gMHa0V1oyRFFl6l2Xw8abJ7Ar8Y1L0nDOsCEZ13W3IVpX3h
U+amCJloIvhpwL3vkxtANAbYv/6flV9UWC7Lg52buQKRzRh42UoAUi7XTtyertYr
rKorbzlO1xKlDBhwjItQLEraAoCY1GCfzO2OLxj4qyZIcoVxyLbEvK36C6tjeqaF
BbyqCgB8Hscq1tZ6x6wItu2bEr4R0rhy7gJO2DRzryxx+h8qo3U/aMqO79wGTjQr
PntWcG32lyzjgxWKqpephmoDCI0NcThiQqf6g6yNZO8pQqH6Rc5O7vv8UWTQ1/xM
MU0fnRCYctrNmCq32sYklE2QZZcRHGz69RpKDFL5J9M3yuphotu1kpw3pxSyw8Z4
8pCUrhcCpymp0/Sqow5rXkBC3SdJj95RsusZKTP89iuraFOCYDQCxrJr6whGvVhn
HK0FHEm4VLHvOZWuRenK5Enr2lbuXuFUXLmJKnHeD7n27xarMlvAEAwmMJboBegn
T0kbrYFE+UAMsh0cC3KC6hmTIjnPpTSP+KP7oAVhkupOSMO4RUp/ZD4gLVlWS9ci
SrqJVq+ZmWV/qqVQT1dezy0GzTawNvt/FMmGanzplBfj4uVkizmeaaFXw2CXccGI
rZnE9dj1A+QqaJShVibbRCkPCjMhWqODOF25VCaNYYuILM4r8S75oJ/ZHqisdfn4
vBKgfXkispoAA8f21gehnlr990hRbwth4pFyiNKkdNsn+r7ul9YnP4I14iDP7ya8
2vYyG2bByRLAEIBZNMrE53GNxKF3pcU+QJ4rBd+Hse7apbDYM8DIUDE+2UU6mMNp
/ahXb9PH0uQC0Q5dpC9IvVHp2MtFy2bnLpT77KOdPgn705zFB31e1ShUmJQX4B8S
3sHPcSRAu0Sal6zuInTaWHN0TvY+YGiIFb9gv3nOTEV24Lig4rh3AzIz5xKPIAgY
QRR8gSGbDxgbHYSWErSuQ8jcnZbTWMEvVtFr9gOgxHnlkQpi+cYreuI5xCeqiluW
ijENNTJpL3hvywCSyZHvg6kJ/rDeyamXmVeg9a2oD6lwJuxIdnlu0JN1bTl7UXaJ
NsEjySiRkk9+O+UVHPVsowns2Lq7RBO8ECg5NyVFx6q4G3pqRllt1qxTlhmBXk4x
HMCdEnKG1Mx7vNnlH/vRI3nHeFLCdwLo93TUpAbUNpqV82FFXOjEXcrkjPJH2Scx
o6z91O/NBIJJRlm8/Et+BadbsY6fAzqLMpxYED7epWqplSrBO9IPHmkUFscfn5BR
dDU7xfF3gKJhOSh+5iAc3ITgizpY8EjPofFczsdd02zRCNox1VIrM2cF32vkhY7Q
/U4lR7PX3eTCNJjnnanmmo9NHohdfMc8bInlGY3KVfpRElJVVY1/4tuCXix1C1wl
tpo+SyqYX2v8e/2DgmQj2eemQoygcr4bYrBHHdNWTkwtgxhGfS+K8Pjj0zy4PnJp
KgN4DokEPrH7TQsnZSE9KuHgpeJYsoDU/cNwAnp9AcpPd1YxFrl0l/hrJqLvYel2
y6uX7zLqY735W9JzPWixOrZxJyyCgpioAzpRjYhDqtM6GrdlCtEXMFZsL3DDgWJ4
ejwQlYkDEuV7vw8vGBrQXtXB5x0WO+X6Qw6cFGWOnfDKsqZ5WEcL7d6AVquQ9eVp
Y6k5AnYJ3J4OMSfPWk9T4hIeMUTEPrusLeSJ+F1ZQxEYwTiAetPaVaLejYhs5uD8
+s7t9vCiC6LtOX/5n2uhe8L2mxEIqofSkXrFHnnlksEARQlHNNB/TwTyNoy7A5uH
2Fid2gxPeDXo6Hb0VuWmGpb+08bg5HuMOQardibzTd3mDZcl6YJceQpyMAljxCps
lcKKYye89WfM1x1lqxu+Z3dRvgPuvm71SwKOpvu6RLU7lsAzojDgIpmXxkU6cwn2
xPzUKt5ESKAT8aywc+YxOpSK0wFgJ5C0MmiMIiXTh1sa2JAPut7tldwYEdfnD8QV
Nw9qAg721yupfno54okWV4GzZyaC3kLQWrJl+UyF/DkxNV0Qv/raEUWAWSk3qAD5
T6SkmvBEIEl5SJC/HIoXHRxA2XGLCJBaDcVrkD0hI8Lc5MLYqvAht3df4hzfHlX2
WdJL4xerVxlMKd/xoYalpboEZHpOMwfCsE23yAhleYXO25DOHVZ+VlRBReYXW2Fv
OBtSGaTO3qiHMbO2guIsiqFKUZutBK6g8XsCSj4F5Hdls1z6zF85DxBFp9S4HkIT
ZSQRFsFP7lxh7ADRh5TViA1zpj7qzGADh6sdP0wEmb7MeN+63rn+d/8r7/uARWqu
zhnEddnvs3H0Rxhgh6c+DMVGNjgLIIhQAuJLdN/H/usM8TjGfAyxU+bbJNbUCv9L
zYmae18EaB7liq/h51wgDKpgoWHeJb3YFjpkDASl7hF56jYZ9u/KxaL7EBURtnhL
0q9lG+1IYIU5TLWHWCkLhWDnefRrO6A+qt7K7SAP85FfNX/bCsdTV4kkimIEYDP/
mRUQ1Gd/UPXDuj5jhVYeylqEZykzUzB8u41pM9NcWWd7jUbiTKX4tmV4nymp2Tg7
c6vrS/GIo9hbwdh/JEbQzJfHy7TjOmMBHYuATeqVu2c73L0WZOh9w3cqAzoUKiX9
K5rgUSs1kUPcTOToauyAUzmEOAd7TYt6ekr1q6jM1xOdzrt/MbNeBPFfV0fWG8hl
tro0aGNDaCAgmL2FZPFlLJoCBlBGAoCT27tOrfHRNuNIr2KfDxyv8Scx+/cy+qRG
TluQrwqRxSF8J2zSzslSCiSVUQZvqAYoMpy1/sG33lNnQaESAcL7VZ9kfjFeI3+7
hTmrnW0lVyrLsev8HbDv0RKFOr2MprUOhiGdjSN8nP8W7aUADQRQfcnxeeNT73jk
Zh0tN2vteR0pRxzY6OPiZdiZo+h/M7Np+b1I6FnEjx9MsglEGYtfPRghkxXdBFcl
L+jSB0UBcDSeQIKymsbc7/HTtuCZ5wv+OoJlg1454jsPu8cA94hsgo1EctX0SFPL
9lw/AhdbZBRVy5eoMggUMtZcIbi5fg/XxST//ZYV9b/9jPz0zBhVr6vXlzLTNOab
xgRkg5wrd4slaIw3yQlG6IbqsPk2EwTuAjcieyugNWWivXZxdvSAkolT7u2vjp7L
QNudoqh6q6qPQshTV1MPciSDQ93ECilc7aS7gdKFQwkYJ5zfFjz9ysBrwb6HtJo4
xno3yhe3HxnFxDXBSV/zZ1gZlrSH/iBmB+UTYruGPkBGYG5h9VIW6fa6PZO+j0ZF
wSqBehVZTv5U8r5CUsbuLI9a20yOj01A57n/Jx2UOJNWaeJFlDIldaBQr5rY55Qc
a3PXCXRM5fu4j0K3NwPT07XdSJ1Y0ksyRt5P4ydm52DbPARmhHXVztYY7XOUK+xz
9PfT+q7pzYDc/Dpr7R3KUJQGx4Xfp5ZY+OlIQG/GtFZFaf7HBMPwMCLvXk9Ki4My
z9bh3gz5k8CUUzZRNWnetLRX00dYIy1SlMVjfK2+ZYkLVrDD27GFZXD3nGpSUE2J
f2UbJVfc5b63pSeV7vBUT0edJrRQ39L+/Nhr/Q8nANweXf5BIxSaMJeUPMK5psSn
gWqtESLUGxr3+qVvVOBKAchEPxN8W57h5K2yGSR9SV9svTBfQzfUmafqgAjD+EG1
M7lyl66EVvTVW/+m9Rck7rkcHj2pXK7ELiVjwgIEYHz2Dm+qdmpSYCDbcHs5/gHy
ioLWi+mHrW1vNfT9hhriuCMjFmy6m8BIXv15rLcC+knu4ucdxCmQi6kaR0htEA2I
vKMmfbzw0rtMejBptK3HSJh4+D++Bldsk87AewqvH0MYFOdfoFVscW3oWLTnlbvc
Up882bffK4d1fwf09lbfhZDwOaF3ygx7fumHL97ShdlasQaBMjzVtdrngq5Q3OQR
Lo0lC0WVb+GeCKVs+ukIL2KOgzvW41X90IxNSvd9bt3K0t8SecYNC7Yw/sX27JQy
fiB0RC8t6QzSzFyvuJd2tM9MX+JzWegi/0TdiZiuST6ibiWnjfauu60rNnkR3KjY
nshz32SqemLQWND3J/nWweXcM3KE9PEylX9tOmbU4zeGwLWkAfALUEg5XW//Fm+j
Cdsf2VYBccy1a4TDMWtGj5SKiiZINMpNoVRoGlIURsatZeAjWPV4DK04sqFFZgvq
GPmvIcl/i2TgWq/YsTIBGaTM5zgmDzs7MdNjhls22ZacGGCUkR/XSUM1BJHACylU
WLIw2W9wk3x87bxX4vXMffg/SWIV2k5lgy1l6fRir8wkZ7aNDqG0pbMtqooxXVyr
T1hIaSqyGuBGC9Hiyvx5FkpVhjyzq90y2LqcZnztLAcUy7bqIUiAEyJRZ0WqvhWQ
8NS8MQWKx5yUaQAnS0khVB9ixlTE7EFagGDIMKOxNkKQ9ZV7mdFOztcbZDzNpg3F
FCj3n3VMfQcm1rWuYNXwGgY3bUFcGkyGds4DpXfWF4PzIlF3wouJgCcuZ5cTX1yU
savdxFtn2SEZvwhOhPoHNqDGgn1UOKCUEVrG16h/IA2lSla9XG6EGtw211CIASda
bksAh6YhOpFA1zO1VijE4lJddSLmGRHnKiTAY/sV15EuTWGv1dd2yBVcNwFc7iwV
bOpJSMCPYHcUs/TpQlg1zBxaY8My4XewJ7rD7ew35phsK49kqawr4E6JxK8bBzR/
n72ncZ1YLdFaywEwEBWJhuFGC0Fn+ECg00qbA5oB0IFyHN6JBN6mztSC5MP8xDs/
/jMFxBLAbCZhHArOcNpZaGOzyBYLQA4+Cpa9LnNKoTirLd0d3aq6FrhPtIOJ9PgB
w7qBwCW3N0LwWSNkM3Fa1SH9AnLsV4mBjIW5mX0vI2wG3QRDtSPlFz4G0HFKohy+
n4w+RiBJ8VyKGGvDvEEfVgTdwQlAAjZN3KFySjUr0hAa6SPG8RbEpMuEpQgMGkJ+
2spvR0Ug5AJLG1XkHJ6ny6uTAZRyjraMR2/NyY/UsRrvGdwPOGjDW4P697yqemCp
TH/eThuSZaRfHeoMtpI3tuBC+ZhBFUpoIxT6cklysA2PhNRY4auYIZXSlGD5so3o
glZFUflPAU6zqN2W7SARrZ/V98+b5uY9Ze0ISXYyOabyVB8iKo73iB7UaFcsQCsh
ZfUJgCm+YuCV3jjWmR0fwvdOBtCp84aAtT8VmOdeaFlVk9F2THjw4AGHfZQS5DBc
ma+Y+QxrMV0SEgsmSksv2M9sJdj86qMlSL5QtsgsIaVEX2sYXOr82p+z9xkLNKDt
yZughznzxQz3lcTFZ7gKdXO5A+9bLaEGaPtqhQ4/BtelORApPIuRjl38UvsWJHW6
1umZr0RG9+TznSUQ4Uexd32k5rj72HSYbmQMF/ldM728wJZoSd5kSilDxxAg4xW9
cXAW25TYhUv36NG0EIyNAFymkLz6+JgGhL3dAjGMvhcUk8oXhNAynnzBak4PC9D5
a42ztFDbL4eKGMVm+Ykhee3+8yeDp87afRjCTQtZmU0NXq/shHg0wnHSBGDgRYia
oxOpvXYmaGLcRTA7VR5nKNXI5+MyeGJFjKTXSx7ppbeyU+gYE1un3s3yEeknAdNY
O8um/NvDSqIG2e0AmIJbIuVlzIolmvXFWQHOf7ppJvijKy11nYoxdxVQUYQu8SEw
DoYcQNkKXTuTso7YP21952iEIOm+1V4gHOqH3lMKg55L9gdymdGvfP5R56SCy9et
8hIC2WktAtWHYfa7DlJvsujxymvlrfIS6E/D1yz6rod51O2C2+UOTA9qYHFotqgM
yVTSurLp+2K6hkAC8HhzecUFraczOKpvvSzYbgM2uP3yYFddOcJdlYJBejSXDtsO
KfrzPBjSjOPzEjIBLBg1Y+J9HD88mVbff8H9uOxyoCkH3qyzRcDp5gKuj0BIkAZF
wy4Cq4wbzxU09okb4nIsvi2mSJV//x0H9nCPa86evKugE9sMG91ztfSqcxBQlp3Z
XzHF7IgE/X+6FH4a9aiRx5esIzOkvKAur4JAJ8tghWWcEk4Hu0ZM2IBgzPqDVmBr
5DtiwRKB4xtEC6Nj+hvQoeHzoke6zaFHtP703msGbkJ0WOTdyhZGy8aaZYKfOCRf
Mna7LKuHx6mgBB3EkIsbzTC7+MYElVZrwQscxgoLmCMfmq7ef+rhEqLhaOwUi85W
bfBn9zZFE2ixTWF12XP2UWJP7DvDQ/9C7bLR2KbqABLXH5nS+wyr72uX/8taJGd4
plTHNX0rmYLn85577F9SiYYZ3g8MJh+GGcp3AI056wajjOBRcbaPbCU/ItjX2mUm
RhKAt7YnkeVPV/gpv9csOm7loAMINLvPuHTV77vVLLdnsOPNvz1MM78KxswTAlHz
fr7T6TM88wp5efnDsiFdsoWsgADVqEHRRJsyQeWfYHuOFV9oFk6ZdtSz7IK0PQ/p
VSAZbddqAHlionGoYjEpM4h/vc8aYGQjSKJtYkueh6+EEe9DSqzvxy+jSK2rkRcW
zj70OT2ZdaeTImdvs5qgHZ1iwcKXryEkapWJ6v3k7nJoXqTc5SyPT06LPiisxnol
qS4jAkd2WKuleSvotDnN3R4+sUniugI716/ZeOe1LwEj4a3erl2n/454oPP3W7ft
02GcLPeRZ/JrmoNDHZWX2DWzohVAaZIpB4W78ve3LNWxbqFGRPUL6cB+d0+8sT6z
bONZNMP++pGXbol7TIW1KDfGTE+f7MJBge+qFzGmtAyAfkgbior4vTLNDF3QjdOJ
+sVmyNnLFX6oLRo4UHtYvDjljB1X3Ka2zCbAtBJhyrq0mo0SreVrbNfNOVkIAEIp
P+oUnYWNsK99Xon7HxVWgjhUlacMly5QIicn+y/aS2dJdT6V7rcZb22BJKGLYN/d
kPdu/gSL5bmXeF5c9Q8mJKxxQ01pQXK39qqz0sZ47RW8aETefac9xmB+7nJHz9+D
HYf6UbtYzCqLmD5AAyB2OpsGyblBSavsZrN9Bby7Ho/SlrKWNG+DcF4Sa+XF9hsO
Ge4QD2dK9yB2+FwIPjiOxcEJcVDFrqJIzl07L5KVkkNrCNIcuZFJUwxiJ/3MVTqY
2hiLKfzo21b8sj8Qa0LcAp0s6DvFx05FdM3aOdDkIFZ0yprnQjqE1uf4zgXaE/2X
5F+BTDmy+60BRGb0lTpYbGH3shQyimv37V5ulB0PW8BL5TSpRt6YV8pHAETCq0LV
R1qh3+7VXVYimfCWmrp+UzUOtHu+sttfTdJtPyyjXiPg1EtVminWAuJw5VN1g5Rk
w07JVCJVuLwvEzm8c+8hRLWGooNEi03tdooWVYwwnNlzga5hx5RxSh6+vKuON++2
4oLHe/OqL/1FHG2pQTy5azOYPDfnzzAAtXPU1W5Iy5jNjB5skZIhXWs5u0eTrSkQ
GeNVSAz7jU+pn5AWwTNxtzIfPA+W6ReM4UGiojVpmYBddvJLNP3FV0z6rK0XCprA
lYHA3SB/OF3qm/uaNoEDjs9w950Id6QIciHIhRsHsRwn132NxmcItmfKNKwefIIW
ksg9XilrLpvTFWfK4MITAfCE5yoe97Bt98Mid9aTmy/z6RhZ0LEvXjM06UdWWU2w
m9mle9xFz8lkBopcfRAn4cxX1ymBLQwz1OiDdfRWJBD8taAu9I1sDydmpFHH0Vmw
gRGYUFRjGg3areFfY+x4A9qikfp/W3DYoYho+8/3lRUbFfHKUyjRm5weoFrNJXjJ
2FnPeLvg7hjfo0kXQ3cp0NZyjbPQA4YRwQp6TEsfzUu/G3EO+UW8FgCzrOlScPTb
vbcdmQZMuZW/CEr6MEZvN00c7W7YcgbWn5V7mAMM795FnG6ztjVCmf1CQ9kpaHmX
Qaog6zV9FsjqQO8QaZ+vMnzSlz4eaIrUifFaThWDuLDJAP0rEm+Vo8QsfS5jMYKI
t9R3IeBqVSqgIt6pspB8HlgK3SLS8mjz1lAIAdweWmmqdOANw1sdaEnIXUxjLp3L
k96Bd9iFboSA8gqWkbJjFEU4vbuqteScnYkmoi4cizfa2fVYJaA1EtgmE9cQmMH3
ay1tebGL21kWSvghYdBgPpIQW0iTv0d3CVdA+BZwEOBPzFKGYkljgnbJfkgMKJ3q
EoWlzvJ5GUjnRgi++QG+3Rq9DWNG2OPoLFKvcoVJPAxwjSeoBVK5axMIQA/Mq8qg
mSz1gwssWfHkFqMTvIQHctBf0khiwpIA4YK6lGk6UUV1meiZEYOG+dcESw71DK5s
fMHCIvODpR6a9kHVceOG+wtHtKChoeUgQ5z3ieMjoxoDCrH0JXgu0eJ00GpmI40V
ZliY0sx2QMdEK8/BmT1TsORwHPa2clO/5kJAL/etZ43LnrM7tJLM0R23W7cA1yvU
BPXQ1cZIRlYyjVp2JOIfr8pQxnNnuNumhhfrbIihuOK+TAjW1eI/y9VHfRQjZxVk
To15l20E7xKQ/0EWllfo+slXgrwGF4a2nu7R+MxfSO2lFseuQJ4lwG79fuUGNSGO
m936Mm1Ktiyqawl4TEmPw/ktrHn2JW8c5VhEC1aDqHlx5+I9AdOdznUL7hLntf0A
EsLpGfutcYzMNijOw1RKTVF96eDzuow3AvTiYVuKBx3nQQs/bTW5ZGiapqUdkaZf
V3+n+nOZ4SR9qFVn8+zQ6OtFhEIBj7YjF9JKKEKYKCNitIvYN1+UTUywiJRdNgLX
UElGvQeV7OqHiMUKaGnQbaIMsle4N8zNJnhll4TwGNaY7EKlWE7Q//Q0QdbXg7xJ
Pm18ceBQLyYeLJqpXn3nWVAkBJObx81zoqwjc8WZRq2/Ec/4/XaNPXMVXXvROoA9
bx6k+iSEc6BHv8fY0VMxsJqvl9tTsSZr3FrdTCp/HYAIXEFOTGohyc1eVzc961Vl
lR399MlAkvzWvBgNqrefmm9bwHxmgfktk1aNh0Gr0P09DkCDUErYA3QlWmBHT4Gi
yN5c3t78+PAkhkkGqq71Jpcyhovy0Hf1+ibxKYwDwKQoItEIhMCOY4EwDK5KqBOA
g3fbf3oLbASL3xK899EUkzm0YNwGiMbZ9RVuw9pFXQrSKWgiRk3P7SEhTezBFozA
2Qew/+s2VxeC2mz84W7iQg9bzigOKFleszNwtXU4F8mH2cA3BdSoQvr3fHClXvbd
xwuqsfhpQXmA8eIIz5rNUjxVAiVTuamJOtIFihexkBuJ72NqaHY4Rj/Z1PfLnZ1d
QrGlNPV7mKlFEzNRP93nT/ToVwKhX6wJt7AMTyiWxkHjYLImvUD7W9xPcB+UI7HN
ZsLYpWYs1C/2/9F3TYq6oDwX1+TrgCtNu2N4M4eveV/XMe6L8eeBb+wia9qtL07w
agTI1IxmXxukTT5FIdm8CBlhWkAbnhgd0a9n6pCgwUM+WDTV11IztAGy2OV5XGj2
Ewqx2F8FFOY1rZNm7e6Xvlsk7vtkSmk2Iy9Xt8H7FjGS5avqRvHECTCtU3+lltz+
5R+XsK7hB/SJsO/qQA9OvATG6ATztJPDfP/lpXrDWWj9KXrQBvrd6Mu14Qf4aL1/
kDl8Sc+c8XMgcZ7TQE2yAS42VjsFKfV52XlAc4GkmXZaR4e+HgbDrjVsrjhW1gkq
ibUAdMrlrgOHwPVjl9B5X7k/4MRX4SbB1ZaMYI7OS440ypXOIHy3DbjJOPof+IwW
eWosApFDbHTiitaAzZJIdy5i6otHMVBL93kp+7I6sqC4I1Zm5nyFD2RhbTU2a1Cc
FpBNdO1BjMGtbGhBoHxcU3+nL5KSYyn2v/x43tx09XBHHpwOnpDO//51BE5qqeBQ
Xo78miy1FKq7+gHD6s3fKC+1oCq2o6m8cCG5mXKssk8uM93Fy0JIafBxihHQVg1U
1ZOp9Xh0QPTMw8OogKPWEiAIJcr+cFkNIBIFLDy4ygxhxvH0Nd5+3F+Ko6wd6EUB
whg5S/J8zwxJ93jDlsWfvlg5EyfdngGqNpB3uz60Xn7UOyjRhQkfUTx+2ObjsnAc
/n5KE5MKgve4BUV4tXzcE5S4KYdt/nqVj72Kk/sMyXOSBsQATEcRhJ+pAbBxab1I
aFQ3jzQkvAHAhibdPM6PrgVaioS+K02BMAudj3JYTv7DxaVg3T9ZP5qeOc7GZ8AX
gF0gCe+E9ZLgGPHElTtyB2FahyoB9P0TIZwcLlaF2/8I7GB/pN41u4QD0+G7THNW
kTjvtD4URIabtkK4R4NZ9wMPWmnVN+i65O2kUe0WSBxYZ5Dmhp3e2fDEYZ/RG78S
fyWtLWtqFRCmlHc8ZtYRomMfgUuWe5W2uqxOGJbfLGwVR2F9OXQ6CTyEIfF+7Obp
WjvijbKoovPw/SSSx26siHEE+UYxOARLZbPydRUObFsM4n54QDsRcmx94AieXw1E
o5FtbTer1Znj2ZaChryGcGl+YHKLsfTf9Zo7vqKxZyUvCYgr4lNLMwOIJWkvWe6l
1AGILNYP67pu2AFWF4ro4gH+s32mlgKeegWMBFT8bSFNZfVcL1LVJds0oNG/jwnY
CzrGM5S5vl6uo0BPxoSl0IK6SJVVrw0YfY+MzUsrcLcdiwmM99PAqpabFTML1NfE
UzRgdVjvH4Gx6xfPUHBJT1HsOdyYyx4eVVnwJVBCrEW2uxox7ok2ycXCLBXOmyJX
qGdGXvekOCbe5uoQIsv+DqeuS1QYnzbKmukfpK4rwLY9FmFZq59qC/2lI8eDB2q7
N8dg+K3XKY91ulmdybn3QBKki40tenGs0LzkvPZPnNtZWA6Rqi8pi08phqXm03G3
7qlhE+I0XK26lKNoAYGJv6VJcnMnHfM/uJBSXQ91ImNFCKKL0eKFY0FuLVAcd3An
cDdF8S/n0YQgOBzLNjkC7H/tlSlrk9Xs8SmyJJq2trFhpYqmHoEJ4mMPoHb5g8LP
k3zlFio2Fqnh3Tfjf7NaYQBmLSTZurs/gMRg4YFNa7uZSU9FTICVDNvnQPpSS83u
10xx+ivJvEUnPZo/Nv2CLF7vFv8jRnlM6KB6PSuO06WnsWtqjfcKIHfnnBmoTCfa
01kN0NLaVjyo8o12W+vfcL3GVgcEVeKl/CYnwM73O947YoX40gwovQZiZvvT/Bmo
Q/lUssjP7eFd47W74kp0MWZSM0FPVDeJIZFU0d7PlU7cFyXsFLZpF/wKiRsFdN5q
UYlM6A2TGjf+Z8bPs2MTuq6Xl8TSY4CBck6Oq8/2RZkDBzP0ngzg2Rsupik4Xazs
yyygrghZk4N335XL8z0QaXAJO7d8Lvu/9ulC+ttxm2t+L/YfxKY7yQjQTCiGpq8E
/BXmueA3OFTiW1xPlmLChVPFrlu5r3tmOOHlCdZMx7zGjHyrEDQlO3s5cTtigLzl
J66M30lMr9E/E4O/7Atipc3A2p4p8u8fbcEwMziNwvzYC1QDb4Lz1tKI5jmkuFqA
M9+eDHMJBOwzzW5mZNXUqWZDtALvPipXtntUxQOIsKzm04wyR9SIHjU2HVRMNSBl
X1DLJzaAcsVCW9uvLMAUgZcAOGZZZX33AJOM2G5yQ5ly4SPlBheotI7vkNzcI0pv
mW7ox5IlxfJ3HW5ybDZ50uej580VSdkqd2Jhi1RDdUDA3bQ+xGanH2Zw8KLqEt0h
D/QkTWlZHRzmS3mVALVDIAGI88rk7JcS6ANDI+Qw+3dtM0vRkzCuOgNzC0SBlOrq
N5AMdONGv/UUI63qtV9PvoNYdst97NPuYzY9KYimN4WzqD2wecBF848rAPDX0ziw
oaSd2C6TL1ytMsEsV8hkvaqzJTul881AE3kzfJdyGF+bbw0eR3lH8HiY0PwcdNiW
kp76AaD35UPGrmtChb3w3bJLfBdGY6jjotNGPdIKaNrp9T74zG3tyIWxzFdyNkW6
Ubts1KM3++vy/5GTyBZMCH6uTHHNbe6XQTSgFgVk4wIUSTK/OiI0EUdj5hCCvvjk
SzhvZT8498LkQU31mfuOc7zNzMxar/KGcX9iQvYNNnqwA0er7y2/GLuYnWEYwSd8
bapHcXBj4impc+zVxT2j86IyhYdcAccdM22HeupdtjnTEDy0oi6TCuWS6byDK9Y/
npu2jVlf5iVApWe/DxKTjjT3ucoRyMzs6t4I4IakSp4UMqGZOf9pAlmStVxOPe3q
LmNkde0TJZ7TZhtLky6ojlV3DU1DEJ0T2yzWcAQtUDn0HseTwISoiBvVToFP5xkc
/G4gFl39UIf/7KdttMl4976cgb7Q77+81E6hhFm7gypWIhaM+/AeB8jNGx+YbpQv
Dkq2jssd6c1MXQMAWDBjYGLcBYnIEQPsjaY9smF3wMLMPafhbfHHjLKa5jd/y2/B
04UcknBESV/U4C0IOYUmVrzRNFHa4W5jV2+z+IufJFlqPMOLZRM/9HqkXxXoP1qE
IyTUR9ddjhjvD0J/5dTTaSENytTXhccJ+vw3JlZGFw6utnjL70NKM12mOF8UnaNJ
YIjv3TnVN+SybNPLbm7AYWqOBPcjlEeBxEDZehKPV80fWXp9AR2aTq01C3eRRro8
uLK0waMXWenOGaDtamgH3mrsNOBaqDrgySV89gKf76ZIEe0+hCa1up2Ivbcvg77N
7U3D1tCb06BOTrhpUjPZj7Ep0aNl8l1KjjoSeEGI5n/fyLa16vR7OCmT8+tYslH9
oCD2ou3h2vqX+3hJiuUL26xq622euDyUnwrkhPSFF1M+YYauMN9t7L+gC65pghiq
WhewkNb4QKiHl3iQyLySYHevh3ZZc8OL/xQKT+bF/wD/zAUtsquzpl8s4dYwOP2h
+6QnRTZ20oh5tHmNcM4tCKp/gAD6C33vipoil+YlEWxOaKFELw+tnFEc8oRD/+cR
Bs4XiwRneRCmbUyANSe+WFWyctnHh0tK4pMdiYi0tzM1Or9D1+InryrS+9HkSgi6
GTo/OKTsp/nNhstdIj0oUf2TQG2t674oTIolkkXyIyID+JdlV+5x9GYoof+GehxN
C9lCIG3BUXp2PXmVv8lfaSgaWoytASEH91byBTZXMB/jFJS2ZItAWpshUazhvnGJ
QWmiSyyPhRMkHB4l5dc94RYO7wTZ7SkLhAFCxmUmF6i2UBmsfLW0H0pOkJJTlY9q
xabrK/b0+mRfw+MN7poNv9DJ2KQcQ9DwTirYllJSxB7QC6eWD6SrOdfY8bmnUh1o
GEEBW++KwTg+BfKXrZPmGak/k0BvPOOxYQTRimyz+NBn3IJCc28pesy768Jrvxx0
vJVvQwm2BxTUfKF8CjFE1+A8aZKx55n0AvoGv+PnY+3FXdxpX3uylDA5b6VFYWf3
ESR23PbBj1cYETOESySq9xHjqT/fGhwzZLbdRgqMEDXRXajcPPZ97O2u3NfEV37A
Y0vdy1xTqu8REKOj/eFPTupJCoMecmV9UM7CJ8fIOX8WDc3ZrgIRVMudrIU7TKfN
PEUVX0trGBjvHMfEgjQOxEh3RXHWz2HYLlpKOZ3leIQj5OO9shEEgkG0NZ/bpVah
87bTV8ri77uI2Av3f1lEdqKIk5LCHW/gYIGJjrYbFQq9kEuBA9k24eh+MlR6l/PM
Nq7DWJY2WJEcqQYKHST8UuRu+UbC//P1dRDxUTRuS73L1Yj8IOWD7te4yeipmg42
Xlsm43XuSroKjG8tp43V+woBIOdcbnBUMVQWZGL2H3XWqzlHk36NkXl31OMN2y1k
qqfevOKnI+9nPKoOrN03//zVzNWhEd7Qs4Uf9CCBLMHoqzfa2luk1ROVJWtS6kSu
iVPDqEpihaD6bZ+HXe0/YBws9qfs/umysiJUVgWbY5cS01A0tEIjl2GMw3PAmJ9P
FKLTOyFfNvEdvG9DE6cbqf4fnz8t9MfT0CNd+FF4odhPo7vjphELd1umOSqRR0bV
qBQUWtrTl9DpIfQKm5Q8+QxevPMwxI3N9BoLpMUTubo30NoHJFRtUJOXLYoL8yKl
ckjQ9HCs4N7QxSDSwMqB2hzeAe4FQsaPk+Ga3eNGfdfMqgmEHJt0FP6VumMkl+gT
X522QEQ20QLxelks55RPxnj6J7rfi1+VJ3zY0fsNV+gc+sMFMudlGDfEipumtoin
1gu1OLxq3ydQk+kcYllqqLnukuMeJsR9mWyb9VfUFUiDnQOqc1+pdeGJV8VI5uio
1SZ6X7WdmPl3D3P6JDyQZJ2JLKmVYSIqM+slAIowkdXIENjXCaYX7CQe8xEFbw6r
9uvjNhthaDJwt7cvq3iJJRJDO+ckE7v9bPluvdN7YjfT0bLqAKpQoWWrPFWrm0As
ffV61jjMkADX7rjbnRyFHSF/JqGR6qwVkCmCGVudvegOcoKrGrhDv0Jth4sNqCAJ
9TX6jo9HL+EocDPSehFskQNqv7G64wrVIqyQI2XuHGxcdZ3Q8gTFcJRIScIfMScx
NLt5cvcc+5GnAbVmXZrcHP54Esk4r107iKih8jm6ScmkzIw/BJEOQJmr6ufmOvao
h4/8L7pHtahGH6qtxlnPyj/Gx9nFBKoCdK58sZofMkaCf9HfSYFZ1R75Lm1+pC1m
8izX7qR02Ousc7Cj9pQGciXusJDkrDaaMMvCSB7wtCsMhf+9zLrpEgTlXQlYiMWG
YATyHwOckiKghW4AdC2+F7DgOaEOnk3E0AZZDZCuqfDi3rlEMFhBLthU9rmMg+jL
A4uY4KDLGcNQHWbvu6ROjs2s32fE3mQZXfcMGgPmsXYuw9MSwlLq8Fk0x6W09HuE
2TU2aZl1DNwFmv5QxEBXz06QOpD+Cj/AYfdgZiHqAzMa9J+2XxQsqh0xxZ4ADNy0
nfXjIbY7XYe6fJSi/k6oFpPDUrKC+G3V0qghPxeWg9R3O0XfAH4S3ahInqGLlmc1
UnWj9ZunQVDpZ3dD8C+y/6XedFvfYSVG15Np+BXaEy9LgLp4fDXrZoGq8aYYCrff
V6G6VLQsOcmE1NDSSX6Dw85IA2xx6UoWqcPqI5SFazCsIWHNk606Y7/0h8v18pSr
pG+Ams47+I15xDIKXa9MHUfXDlDCG73yXCzHYGELiRpRSIC6aVaFUQbLrstjmaUB
6kHoGvEM8OViDoaZaikQr2R0B9durleZKU4AvUzSg4Tobrr2yev+dLZCU04xSnU4
J5eJ+nv61DjYRe+scZK2Eu5YcpEwxToEBd1tl3xUgqUulVAp+Jv63ZSIluSS0A6m
VOQp0FBw2ygluvTfpj+pxcUQhAi8tYhLUF/Cl6LEMli6uOet6gUAZw8yn7ul1VIJ
ImFTUA4Bq7paAAjNrN4gVTpqP8TPqqjRLAdkBc6hvmwN9QD5X5rtAeVOypJEdnSq
fbzfr4WxldwDfYAZ2upxXu4APGp2u5NfeQNrs89WZVWAxvOSO6e+E7Sp+SqXtF37
a7NMX4IDbz4PdntzaWEWjaYYryJiFKTqbdf+AFDcWHwuKHO6IHNTO1NHnNfnS1xo
x6Bqx+GYoFDfMzGR3hdZTdT/npF/b06m3cgEwpApOA7InZRqfaNDHLA8gWDYjCcw
vJQ4PbkgvamY7NmJ21+QyYJjkHLmkwuvbZakbwMbVS0KrdTJlb7GHl3OOeYXQPgu
27y26ik29u/DVY3OWLvJQGNtd8H2Zz1mSl1rJQ9LHVLfCubbkM3PoLUqOPdoAl4E
faHPs5cCl0Z1j532OZydbLuowCAmW1vc8Cjlh8O7r8vjESzm+TN8qqKtViJZDooU
fox3E9BBaAIDezw6VwTOWvSCmj6c0pqngaqp7nsAImhCkFoGI4tFsSHwwXNgD8oo
CcFbzuz0RMteSn0nJ0yF8xwqOXeUTvVAbLAa7m8W7GMKmyTHOlBcGesBvRJhM1J5
5rNrRSiWzOuyVLDb4AHPSfnm5buAbPs690f8fcfVmN4eKKEaHjksQxWL31Fb3Xup
U4sc6mQsk5+pq6txJdFsAqpsAMn/MdSCZ/fQJTILOd7cHXS2Kg1WH0qiAVsi3plm
CQNAtceFR+nRZ9uui8AZC6znRqbm8aOQpcM3L+BGSloCgd++TpO0KYdcke4Wwe4w
7rDVGoh2wy8MOX9wydkXNMV+Vvz07DnmHim/1HvkOOlGG3dSZWpNBO+LlNOpH/p3
rEq4AT/jgo0B3PB2nQOWxRgWcXsJ22E8IB8ttIDu+YQaVANFvRWtW/uxURWZNQyi
6ZiO9JnO0g7ON6QP3raRNFaI9Kgh2JdLjKhqkyv/YOQf4Y51lPVczI1egudGi0rz
2iEs5qGlB0oluqnJfjE0kNYKYAjnwV1nGIBm7rKMF9bR8+V4y9Gj6EBKF1wDhE1E
mjtyzXG9Sr0aU2uvs1sTdCmQBkAwO+2QnqnmFKp17QWmAs/D618Petcl/UO3WysR
G74WHd+yc9IMuwSNxoSpH+jwRBNvo7CzIwHrcGxUkwcGO1gqCpeV6bZmeBPNOtGb
5rchzwLXNNSLirS2DwVpb7hG8cGkyyM8ru/xKnp+tqK4/2XpZz07gXHZ5Vcp/12V
U+avDmt0esImOY3aD8ZknGMu9NQCIIYe34ZjDnPq2X0aAcy9ZUYLIINDSPo2Nuzj
WJPl5ST5guIHuBfmIvW7YRviT0hMnStdnHI/NokjKO57+tBpMZIm+uXa/9tfpTIM
iZARsVxNbZtuNm2BQNud5FIBk+7985LJSIiFUSmPezQkTyknOizrI0o41vXrC/n6
VT33RPmSL9siC5C9Xa7DDUs3OG3IULPPoyTI7NXB5jQInZ+2peVLXPnflyCeLRqY
GUqS27ZCaCneeu4CULvdYTmTIDHq9IO6T1yoQtAQB17jRmJX7GcRKJITANWmjCeD
iJqzHtZyFWxsBb0kzPAqLi2jcjKq361CIosUMvO/FHtXAIljIw1bAJ1N3/MhGeQK
5C39QVa9E61lLWhOJT6wPO6+jmYOoZZHyr5MDvf3w2jMFW2m+Okh7iF7dHCQ2Qv+
HSrZzqELj7xrjQqsTlz6NKuK9HYrt9IKekmqgbttnB6xCyKkJtiILTezF68EUhjn
68x6XGNg/SYSD3EQe9FwRRtdiSKZTncj4wNuTC4/rWRoa3LONchgRVaz7z0Ktai7
woUAwxZYM6yLRjTFQwX8wzAEogaGGJv/SNKXFigUhAqWtbwXbHATo0M47GxL/bzj
0uVmT0CxA3whZF1RVDvxFOpfzo6dNBE2fczdaZKWHj5dieh55cZuDBSmWTWs8clZ
23/YV0Wx7A1pD/bscjqh+VVU9YP7THB6H5k2aXSDoHFGENyHfr0kOsy67EQQiVzn
M338qeqGSPDiEQPxdfy36egSi/JHi6msPkveOu4b2Ij/EMNo+Dxx6yMX19yYq29a
+I8PwVajVlwfEua9JeAxc4eLxQRoKq1a+urJZsbPeuKnSzdHZY6pEld8W2bpXl8d
L99v/fPDSxdn6RQU1jaoI8phF3KVrvLuauWhnE1GiShRktep9Bs88/zWQXQhz3sm
asbuTB/+3UR0twFGCBNANWYPhkZ4Dk50JJt06lvn10hhYCUKspabq+eEmAIsRx2h
zMW+jeql2rGq8f8ich0PHCKbFYSD6lqdRw1c+fejEPjQEnj342+Qll19ONQ241i3
Nxl24SOxbFng5YJyV/8XIHGSgs0wvSc4gv76CCDaU2sEIuP9BWeyZzVh0GCJBb2t
p0F4iN7UIGFXL7zO8jZKwN3K5ToTVHgLdldEWafmmKzp9FLNdABt8UUPB+9KDC29
KgUxrX6u8MOeKC99W/2UxBAh8SUiNQtEdUpUQfOXbo6POEi60Jy1W08O4+EQdEdu
Lr+M+Wv9LGnA+TGTmg/ybHEubgtwdXPVPxtU3WnnDVxpgTgksyU42PXD8bMyXnyz
O1T6YgLBge26zeps6eBolYakjtQFWCUXBd5ohsGtS4xDGMZ+3Hlynicc8sIAmZu2
tAnxc23HFSOlNgvbzBsKqbtwbOQmt/3vAHls5MN+A9Ti0/L4t60hFGGz8Bfu0tHI
UD+NEmSEkaf/j3ets2URY+x9eXVlnbJWEXYGsTNysoDXgbo9kNGUlo4su/tFQ0Qp
VH9keubLi46ukydNcGseT5dAYRNRytWbUre2nCC+JPTILTXU7pNFzya8tNiIb7tS
G+M+L1DFIxv+FT0KKsZuRtR+RmXRT6KrAypcQVnarz7ZUEbm1jx4V+XJ5yBRGsDJ
UVz3QxdbsRotncVib4WVLKdnvuDeE+/Kbwj61V32w4Jtg2gwHRAXIHMHHXhaF9pF
zb6goUeKSLh1DbGmL1iuEiP2c+Kwwvd8VJQGsWJJY8QIhOlJNLcb1NWOrTjgssBC
xusnWJAA42ScIuh8vuCFblyZEDajSO/ZE9j1s7eZUIR/kKc0f82LXOGZTlJJ7lS0
9zNKTDT+jX1cftzQOgIKHzt/fsWFVj03Y08hQu7f5576YGioNjDMl25NPQ/7TWks
RUwPOoFJeEiofgXdNWXxZfJM7+b8furxIt4kvtoaEcRo55hjXgK1pEU65cO1pnOm
cunv2THIh4Lx6dJmKqV4XW+PV1ESMN5avWyXcayMRPqiWKO6aDhRfKGDHN+B9xK+
GISRthwzEjWsqgVJktvXP0WWVBHC/o1rmMGrKworzEG0gDbMjgOC7C8k0wLXHEPB
ACMcYG0MsbaS3I8Zl6nEn8BPSZjquzBCQehjS27+Y+jzGBFjfJ7zRlGAyDf7vSUi
f/9HF7SyCoLtMPhyIcaDVsIXGHuAbkUannUkiadjISwkPIy4usg1c68B3z3SZNl8
AYcuNE6gp8a9GWePzsiYenxsbIxpW7SBD3EbgV37E1gYJQM53LsjqUMazpKs8k54
Lq2zjpK3SPhTOB6NExWgW3h54ybBLlW9uLrjrdThyoBEh1hobNxAxfJSVNrDj0Bs
xpcptZPMsrOlL0MgyxyBrDfJdAC3e+dzRmS/6tt5vju12Zv//C/ZGjEafsz2YQzE
V34Qr4TOi0VZZpDTYz8v1znKbxyg3IfIlus2W5j9HKAmDCOlYnbaQyeXW1LJyM3X
dQibwJbXSkRx6sFbf1+URfvyJtXDd4AqUS4r8tnzcAe/PJpwFB/sTJbNNzAPd+PC
0sNTQbR7VSNBVdvoqWAwTcKzAxQyyOG8LkG5PmBUYidQlP9bL0qIJuGOlUxRxOPJ
QR3TW5Sat+F4ZeMuXBaJ4sCm+bRf/2L2RO8Bie/X/dR3dFaT+fXUiTKnHezdmHyI
F9TxBtWdQDfqF078Ci9Vvq8QcRqyu4AQTv3+18sMDZz39jlcr6HQFyjJT0Bk8QQL
+yvIkznHlfHe0WAwqMlhMcu8k2euqwk7rnAVWiBj11yXqzuMsCYHlOvHaobs4khm
vS/vk40+wGtwGYTmK7EJuVb5sMxP2ptKnmMFyh/knEK0giaypHY/NsBBuJONsOrx
hXu1N3EYmZ3koVjDZlLcwAoVncCtNiP76CtgODjm1gF8XIqIt/i5KHQk0LneFTdP
aobWzbFz58WtDuVIqT4ASigaMZ4erd7D7jUHUxSVEpHfHrsdVCParZvMETeenLTe
vbOfOM4Ah0WkBH86Y1ebuoWgrsHau7VRtolwin3UuMZd5WthJUDWfeSNPI2TOkey
bxdRIuAvil/LHzNlKX1McoB3IhMvZaWQYmwsgUnup1YdE+JbWErPN4/+bdoowksC
0BwVUhYwkKm0dytwsIkI41NersqddNyofrMwFk4md0VyDre+WAEgcpc8JXK7jZz9
8MpRbkeFXxKmYONHogx0X4H9NYxaw62+VsobHMX5M55yd4hMrMFUHQElSaO5DsDI
K/QwlaNBiAlvCNenQND4MLeTjc3KLSaJvBj8oR4xrm4/JCmTQWucKdeZmZo50e7i
FNJM8+veZNXmiJ8Up3hel0AKoJ6unjnObCLe24BkwBToin7RkJPho38Hn5uZYVKW
GSHKnqwudTnlzj+09APOlrPcdFgFnxc8nwtvbwNlumdDuK2WbSchTqEOB6K8EzVm
UrNSedkQcugaKSJnkViBTSd/9t8JPParSnKG8yPhXC1ZrjR+Sf4mmWxqBU8isuTi
hB3vQMf7gnZQ8BPVqs4HrLb/oB804s01PB9z7UgbCneXCL+Kl2hcXZeZF3gO+iJK
LtafQczJ0fEstqCnWgcyE3Xp9IKwfqZTf8mGJ/mmrXkYEeyUtQ9oSDJhIhI/fG5N
APeXPGCpJFXnX1XfjBju2J32VcVzNcZ33+sk2b1JKRdFjg7fu6sZckL+lmxqlOXY
SN7dpugA+vK48jhiMC4PtYBOlGG4AUc6ctjFRS5HiTSnH7B1iNaHOEvE68GzBlwO
9GUHtrkR9olmKwHnXYFEk6ykZJahOo3Q3k7uYlyChXsMAHdOtz+q3iRsAHHd7ZRo
t3HRbqGxd+gFB/Xa0M3ZRHhWPfWYlyDGFHT9vm8iZjUdDXhPzLcSVIBhIuchMFWQ
+ZVPkwDIKNLtviXpOoPKy9WFZQY++c0DRy5hZvIZAJ3/Fm5IW1DaA9/K4TiKQM7S
WOAiVr6f6OeZVZaEPyqK+wdcLOKUWaXccbyK3RCS53GmF7E7CED753DfcMbgqiMU
34bLtWz0sgpQ/AGPjiu3wP4wBt2ZDMBETP3+yXZQOq0GzGkZUQBRy7CnQN/NxKbV
Rg69DdwfzM6IE9YWOlxeGXMNAtYDb7EW4s2TIc+oUOMBrgXB1RhVNB6LWiEwcMeC
s6eS9lJsQRoZMGEl95DTqq+G2WROEs/dFJspC3GSwmuKp1Jc3ECtK6qnaEm89RAk
DJZ/Mf4OI3qyA1nx5O6myWDIWkbgV9VHQIC1IzM8nDSCdNWzJ6cMSWb3ZncPK4zz
RDTMTC6V1pBkY2pt7c8EymXiLPPaw05lkDx9QtgvRZOE6qfiuLrrJ1CpZgrOgEd3
tdzDcWZext1+oo1nIzMCC3araxrPcS+uEhhKR4ZGBrjb9B4g5f9Fbz9BAK3gZsYm
KlE++Bpi5BdVSNnDzr7IVs5YGpRiy4Bho/ltXm6KX6TvOKy0icQZU6FyC6kkIfKD
GDMHg8YDHCb8hufvz9cprz9K7Q1kLo+4ExRkiasG/1SB7UQjLUyxlXtS0RAIW7bF
nX2HkJtxI13/7GLEC9HjtvXfFH6LvJ0CQVs7+LsCjgBx8Ra6XTUwJCxs3kp5E2bH
/LW0R0cjCtZDbi2aM4oROc9rO2LMZ9Of+EXGEWssvn7SOS9qLXEwuID56uba9iwe
1+46PGxrE6+X4TIXZB1tVjFr5FgpzKrdCY1ETpg7wdmGPUdwK/k6rBhrfARTb+2Y
HyJnRE4mTTvh2pTKozrnB30xfSZZPClTyGJaW7VLiYie3KrHAayXIdPCZuh7lIDk
IWHICGKtj135rcoWBqTObhuTbntbtfEkSQryuaz3Km8W2clc8a6tqbj+/vVhrsVh
kuu37oFQX+TYKxU8tWXYmQuKAeS/8f2n5VQNCE4c+LyrbWX9qsdFBOjfROCsEM3x
buF3NWz0cToRMIX4EYyOrFmqylKq5hl/r8tEDQ23Ep+8rFeLfIAa9BHIKb68STBY
naw1o0eiusNNYU+qVbQvMZWZp8Wi+yzl/f6Jz7bRKIBLWamEwu6k5MAW5iJgni1p
uLEkVoTEYMpi14mNHwO4glSY8YqBikEsnB6sBi5VHDW067RbnbO11/q6lgs+c08L
nUT+1FKTczXRsTj+MZiKEqA7Nb0NMovDkHEqtbIhfAgmv3KWFs8TieJWRSkqgxno
5oI4p8codUeTbtCW4T4VzBVkLGfiMytogJz5xAMD4572wdya0rnMnbn6YzKwqSi+
0JE7IR9Rbox2hoCOdCBdp6QShuinqAXZo2mWapzhJHEw3KuqnPlK26PpP0Ef0i7t
QQ+5dgRimkXREAHXDbUM64/xTAVFFGCytOhZaxpZkfKNxQtDrCYSsZ7DMOvs0gV7
/pbf0AKQrSeESC0vgwbih8oVDhTh1se7pNoLCyfQEqHUhTzXBTPFUlBe+qdNioqv
vYZLgjWh2xd9FX9N9zOOsJSVfBrYTgwOOCw1ty51p1VwXEdUFXFXphPhIZpy92a/
RzIdG6YtT4ck3IhkTu7R/2yEfmGTg0cBeJ3jYsK1Pgq+bq5jNQegy50IEU19cs0b
SO9KvIXBejwhwX3x69DhoF9nMXW6YjGbJr+gO2lratR/yk+dU+n7iXXCF7zmY6bD
gE3K0KbkaNwd1tq2nId7SbjnBDHntIkIadruzmO/2i2X6PcyMQQvNpwEuojh34NV
85IUpUaumrfYsToZNyVynsm3LjgB1h5AI3xZf/W3Hj3iCbiehAQhyXPyMeCl2/Ub
0R8Ky3iAIAus4vB9fN3vZx6YZJ3ToLuHicaIISVAhDVfBFwjBFYcDYivBWRBhJK6
3SUAOlKf+TSjjSRc8DyxfEjuxyQQb9/WpHcoBDv3tw6GoniGxd4j/ejKIR0oxY6d
TKlKx/g1fga1YE1G8yitoYKRPUAS+BcfEChFpCLgJjoCWfE3hr9DkMAlF2sRh6dB
WNFm//e2gnn/wXj4mT5d8IVtZQJly0Ig+pbwRapMTiCXFGaHL6WDjB2QafiX3Ht3
YbJ5hv4sd7WRudwfsjIHWf0sOrSGR8TGrWMD5EIJBc2tOsfGCTxfzYnZ6uiPPpZt
q0pJL2yQQcHT9b5Ntj3MkTDIuKPrtWiwfjuxn09yGbgqb85zCKe2L4cp4i1NDRQL
DkfahvfIu8sAOqCD+MHMhZjnCz5Ze3tYh+HKCCMzhodtpcbWpIMuhAsaOhLb8MkY
CFobs+I88M1g9U8vGw7jrvg0l69+F2l2N3z7d18vmtiRJ9yLz9lswPZYfWgbiipH
e7RKHgxku14XvFlcwCkMY2bRX6ymsXfe8qycMYUkvPoKy1mqmdZ6GUicq/3eiAWM
HEwt5+xrlWpmCyTFJck1v5T6Zyr1Jrh62DTPZQJwbgHroKZGLwg81QXgD+roORcs
WjILzlhx0zMuVIt0r44xEusuH7beB8FHbqgD+SwkO+DXcpZ1XTwlde8Eoz8r29jz
UZ6kjfyp2i7CUtBJhtXmMTXu+6OzwMamU977mo1agHS9VjOuBXtuEwoNVmNAlSdJ
p+brgPCqwBeQ3K9N4hLobWTww2MyWAXYn3sR9kjsA3/9jVKN79OSSBatHaCnQnR/
CHGJyQoYDPdxMpi6NTE/Tuca4aLn7mmFujpoBuPM1eA95BbXlKgtSe6GYeIo2pS4
BSMaCtU2mNjL87CcC/cznAQ+RIqgs/r858+3KssnU93Krq/V47AzfttxeLcu/sDx
h4wbXUxr0oDmSVWKDuz1yo7mTDj2jm0Ombei0BBlX+L5K9oL6sIl9ArkbSpx7zhz
mdzkBLkpDucmXG45BRhPuodil9EZfKxnBisnKlN1DsgpGseQXi/Kdn4/U2LRAWUV
6Dt788oKEdMeU4NNdwgizxn5OYyHjgB3TnE4lAxJdeyfYPyQ7P3UiTJhoopjJQ+q
ccEI6qjGFnVax0giaKawgghi+EqwpUKKlwFtfjt5d0APgRAFaR3oJ5hF7YFTusiO
k/BtXxSqu3/F9pnwz3L+h/LBPITU9lStDvumQgKyGSvVRq9Sdt1WFoBS8xG7eNNb
tc2FvkugU7qqhIuzywg8WeLaPQK9WdH2/Zn2IMA+taBRfWAdihGBYiLDS8AWxaxw
1lFuOEEUTeL0FeXjphLa8yCTrshv9+RJYjS34OtVUtw6aUTMZejvi2zkeGCLrzXZ
myhgYXZxoLKDg98we2GTNTZ19poXP/vmwumhEz+xk1v5YGzUOSLRQnJOv0unmeNH
QuobIU1WZ8IKyjvHjEibp3n1A4ajA5uYyQ2rV/hMnerstTWvOBmVfP8/lYxKiqBe
gkn6ocQW49Q387AcG3c05ScWFKLWen26OJ8cYv+hUXTXD2wl9mOnxgPvK37r+EaC
yz3UJxjjZT+2GIGLYDiZHAu3+T6z+gPbedUVwSbL3W4lxs8ApUAfnYe6tImWb4lM
O1p87D9IuaPhTSoq5Q7uGSU2kjuUaUhv1F8iy9y1vG82X0BTik/me91pBBHmB7T2
3xg438sW3+sbDRO+hAItQJKXivBo7aZcN8OLTj10YlrR7Zs3yObNiuo1wEBq+r0c
K8CB7pJnV4X9AOP034qfOyOz6t+/waZo5osOATG7irVI6QVhe8/E+OKzcwe+hbmx
/Y5Ha+fvNkpvc0GXRImxQjpQUhAL6JznmXPaQmGiDAPSjy0n83DeN72w3uUXISL7
BtT2YIWAmCweM4+6sE42MbocfN8JsftraFOQIuAV+JgEPUCNNXFBDI3UIQGZaKW+
U3OnZeaRaFWHWrEaQWPk2FE6Mvi8L/3aoEQ70zhiALxYZlXkokM5TNIxGzS17T+l
RW/YWbuhllmRQAdoPmUij1/DRnowMTcUVpX9bWon1OqcLLZpeb0KIqHUNtXLCZY3
6hNTOuOWAsSNhIT2vK9EDaG8cxQNMUyHViAPMrbl5+r+XkRoxGr9Ruj0E3r2pein
LSGLKMAUcyMQhiSZU2qzqOJEWAwNwOg9qn87tu4BTa+STgNgkETZcV89mwGB0x52
3eWdIvz6583dkZhTCFZDyTFezuikCWq0Byadr4Q45k7uu3OWY/eBItZ29pBb2ucm
hmxiSy1Xrxad1Wy5x53fLHia0FB0OvoQ86ktaNPhyccTE+MbSseLnxwZf0ev6tRl
qb/dD+XbLWIELF4EQ/NdRVrHnhKekqrjoXs/t0L+XOY4GvfWHBUQsrPnfdKu+gJK
EKTYxcNuAa39+4Bjpe8tYXTxqbV0NBhQE+zNrVIpppae89LHBmcZEo6avDOfXi3c
yU2EzXmyyQXO5izQ2l7xbrWFg51Mqd5wFwuz64HduSTpFDmSeDyGB3qr/kk5dK5y
hftt1ZVd6GBPKf4HX2G3fZ4FTRoCq49loOcRXNmkRwoEMji9k7vS6t7Wpqr545ye
8z0uJUGjV9hV9gcE/CW955Zoe3VBbZZD2TwqVWIFzR56FRH14CWvSF4bCFGFKq2b
Wa7aGaWP03eYG5gqvTVDIRXGR6cmVAJEX1hLg/yXRd3khO3ySdRXmD6uUp4BefRv
blb3TDttWI6LxuoAUppp+GNGEs8n8C2v0qg/bu3eteplBNM6AZ9IkDxh4BbLWvSE
DGGDJrkLK7s7k0lYnC+FA+GQUxTwbbd5pNA8dtOpyeqP1RqmZyF2uamRuhlJvrtD
dQo02iskLY0FgVVyAf94cX+CqjEYew5RYxAtELgAEu3WqxZS2TsD5ZSe1kYHhBTk
2+ONqSNXrnoF3cl73qVy9huF1WWy6E4Zdx1q+vs6OK3Ul7OweBGYzFjU+aitGW3t
2VREJXWfTyU6HtFZN7E/m3lx+sNJPjE10YpEo9MLxsSt0GCdEpNTQfwf9/YnbDJ4
TXD3AYzUqVpFZ039SwujCduTqMrBBg+TR7TQzvbBC+vEk1WQYfxeyGFhTisGEXFX
ltdgp/Gvb6Yl7nsGVYPf9wiLPVBJqKu4dxn2Ah3zIYCBALvdi+L3hZ25yLVjYALf
g+dV8mPWDxP0qY5sZxWd6RLd7R/39nkaxuRgmkN62/evmsqEPU13tAORVjEEjczs
g0nqL/WEmRqpKJEZ9TFwGBp+0JfJYA08RKINA8egPtNgGp5JCVu1Z7t6ZAqpgWZo
HYxfChONl7CcjLPC/M8wkYLgEN/3Z4H4lquZHv5a5omsrB5e2huLs5IpS4RjTgM3
os4HUV5Jdlzg7FW3Bb/MXfoccok0liQWCgATHrDtjv8bisvUayfxGnEsGyHo5dAk
OJ/8THst5MF9ZWUSw13sa37o2N1iKayCqrC2wM/btPXtbLT9y9trYRhwZvG9yyYT
Z/zJraQD8DSVyE8DiGktZ0wkgAHbmJauwGcVS7ElqxysbALVGkT3l/4x/6oJ67NX
gyj3juRR5ymxtvUA53scTBqvWFezHSyIcQWbNsGDN419oanYcsS7TOlNV2sF26Dd
gryaaSSJscTBij9KYTyAf9NqhSVVtZaFyX4FcIl9ujdJohaBC2lYZ7cMqph4b88s
kUvEj1dq7X2JQEmiO97aJcx+0ZOU64OR3kC9DM6Cd9N68d2JLTthu/1GY6Aw4p7R
g6NsrbUsDaS0IgLAtovl7eUWxDAdsBdjJvumQVmqdvV50/EYDk5z07BocibrPjoI
Uq3ZVdNu4NAkzVHNvi0p84SFyH1/RsLATTr56CUf4AR/mpqESDGFmByARQNc3iob
JZUr21r2cuvCzTzHWmQxBqLx6qkoHhTqXogZODP07zW4AAFTQkLtWBeEwHZAfjew
xoVKYR/RQq+BQ/EUAtaESAWhH4RH660/txnonyamyozWylbw/N6B1Fm0PB143oCw
1hh1v4YlqJZ1Pp1FA2RiNYTjtKiq9MoeYXBPOxQhsE6zC3UjhNYlnUlPPhtmN4Pt
iDW0EJG1rjCascJs3c9JIWcGXMEbFGbqF4unIuMxgNqPJ8oegW3cTmPNNwOOVCNm
KVJMiw6RltY9jXs+S+/LU9KgRjZOQsWHb09Vmp6dcu9SBwZZ5LbE6PM9zB3tVr71
WoQT4CtNATcX64Y1LUELkfZwBQf3g6OGJjhVM5Af7lTqn5+dM5z8VJdCpYEN1U81
kqrsobA1nOe0IgxTOPI1kuzivVG2MAnOfFS8S+n4aEenlB3/xymRX9s0mj/tFkUB
5WPf8hCDVjSRFNlnwtsbsHSzrNaTJ2gm3vo8w91395orIJV4f0nHSsxwZ0r5lAwC
QXE1og9VPwaBhdWyozjDtLivRmB6UzHgbCwfrkbk5u0gzP/667+KBTSEsbQrEFXY
KmUaLAas/csYTTbEAJgZT82BXbf3J08mk/Rg7fT0wIapfrgKXgwVauZpl7Wbk5cD
5d50lG+f+0RGYAgm6GrzzyBXoUDIAr+KEjupAHJw+6/sy4hwSg8sGp4fL3XjQilC
ZMJ9bdbC2Zis2gKeJ1KWRDTRGXapUbfS6omTOD9DSF8RWCg42T3acAJMgBJ3pUju
5hIXjkxvv+FaXuPpIm/1YbETxADj4cNO7ZMJ0yN+Z+GgXGPiZC/B8li4LivcpP6z
2n8TC1lto6aPlXfZCh9YnQ2rYy+5w4DG17sJGGqb7ciEm49T5w7gf8buHVGPSozx
sG5mZHXYbFAxpYHDoQoEi24CmzsFJjuALvwBw2flwCJnFN/GJt0D20rmdBTGP0dZ
SaBkfU1E6splRAO0/OCF9YqTSafA9kzqd9QPNRAw4E0gja489pLEM1wv2YyOKujC
Ihil2yYYAMlgWJTtA1IBfmNXcl+Zez6Iwc2XMEVFSuZBypwVQfXv6PG84AhygW5j
1usjHnI6tbl5m74VYcklMYLQtO5PmETXZeMAT+Sbem5OR+vjrC34BxYj2i4Bgbib
j74u0h1NP5HxyrZc2FYu0AMwWZgg0ZSTHoL7EsEs5rQu/JGh3yAgyQokyKaGFdXs
/K5RzYgr6T/WFhTl5cTKByDqsbByI0n5Ei4Qe13ZqA9YW3pYL8+7WMUe5vaZ20Iu
ixh7xrhQKZYNau5O/9bSq7FcSX6hpwth/4cPfB9Ycy9aNqQblRDNNhBFF26qCPRq
RD44cuEA8+XFHzACVglGrXYDI2AGHnH1Ai8G3gqJCRSTypAHGJ8q9Hze/VUbz0yD
Y6WhMqql6aCYwHL8fplxK2wPmJRfHeDNpIb/kAnZMQxVvHnJQoMS+V9luULAwn4w
fGHtkxzL6PzxBdPUjVPhezwvxVVZO+rZBM/izcd/W2VfRxtaiwctOp46CO+ogPgw
KrNL5JRyHJN8fq3YtxN2xEcud+lNo0RmKLtrEeK95P5M3ZcyGald1+ZHf0caoI7g
vPzEcDdnI6cqAo95cDn2wGkfZ+PO3hknazKhyoQiJheob3AwucDlUVshCw/hBRKk
ItfW0FjKvnfbUDU17a9Q2k+khqYEpmvlFQkgSV24PdybNBlnBmNZfLDYYq5ccV3r
3ld85NMwEVpB6vLeT4BLQ6JpZBF84GimyDEIQ0dTlAMmPtDY0ZlxyFEeH5iXzZ2h
JT+DaWB3NV19oC5FkN0nYz3e1Hd5bas6W28VyxzP9HMN8aDiueWNRD67Fc/pzuph
agS/P0nsq+07hLk7b0tYyerFdqclIY7Iqo6la2JLPpHhv3mMkQd1zMDKmULRk1Yk
8wZ52HkG9swh9FxtjZWRouVi4B9/3F+Nh1fsXGESH77Jy55/TdnsA1+fi9axomQS
aaE7htFVcKdKqB1IgIpZN0aa+xXfizWD8ueyEk2INKlR+69VSHGiIgBbNsYAutgh
ai1HR6p3PUHjjRE0akxW8qFS10yBS5qWeqbWczRVtD9E3WJMRMHVymvGqMntGJdp
EHMgZHhgfDAntxjJ4W+iymDT6HLCo/Ki0967J81tF6UxEIsaNl+fVzuBUtBdqqws
4p2U8VbF0NJRUTADU107N2OdG1IdZOZTGAoMcOpfLDvXpzdWQjs9XpGqyjxsXHYz
lc2J0JaCPeNeDpcAsi3LcwE4ogmvi7/EisQ5gmV36qzBEQ1v0MYFS6TTtfWRpSPT
Zbo4tVlHO4YR3/1r9CgBvHVOy5hi9D67yRO1Q8OV1lWyvKqxDS3pZ4BsHxG8OLGZ
+L3zJXKzsF1lCvkPQ3Ss0MXHaFihessHUE8y4lBDEJYCNor9RItLrJ/MmZngH6lS
RkH6aLRRfeRgw0g90D5cbq9ONDU3X1ZnBXGAi4utFxaBWgAUfQ8V72wUuFkwyJdD
L53qtBCbMyYitmQZJg0BikJEyBU5JuAKBwFNVYm5b1JYeh7gZyxevCxIQ1kiqFlz
vvB2st9rueY1VmwSpow6mA5VHAZV5ENzf0NXoZKQeioSe5QT71YR2DwD9ehL1Abj
nBqd1dw5zfShy3yi1VQ9hFq8aUmcn0gN/DQM8fAljfNxwadbW8GMMsRtlJxdwH7h
uZbUEhaCzuXEm95/vSfoR7ijIafjQf0fihEwmkgnWeCYWt+eM/euAljLKZxMl8S8
eH4Huq/Qh/SYSAmEyAtXI3acBWFvvWh3S30YOC7fNirRKuKxEX9FmuncnBE+s3uZ
C8O7XmhVgD9PCx11KBihnM5bUBhlschXhbIk/+g1kPxECa9Rs9NWTTYCbOO8jWrg
OsHIzxVMfP5gqkzokvvQnMhGCS1vQVC+8XgljRslTVLzPh3PMm6v2KB1D+hA/Ers
40hhuDJtS2Gzt2n2JJ81dIRx3pQNnd3xIsCeH/I5nZ3H92NxgBzhmRFnU5imkTqY
CJmNUjYiS91xLAiAWIkbTO03U0l4krq/2tML1YbDsc+ZGDckJiRaMyDSfJYmE1fY
UFcBddfhAAaMSu5KmETfv1BZo1sfb9nC5jNg+q138F2ZoHr4l5iKDW2Ay6koRB5p
bqeemRTVziCguDzTj9SwWTiWSX60rsWZAgVuAUgb/rqYkmPro802iDsuQLQfECko
BnqIgdDMCQsfAKYHhSnWt9kPx7qbLHrq/T+qLcseIYrbia5OfddYrp8ObPg1+674
i720uta3hpLqzdmEu0BtfYd2NpjKrgINpoHaJyshQP+nnmKk/6E4deGVjLecGDO+
X0BO9HIwRcVBShFb+x5/KeU2onuM5p/orQkHWS/tg/OhAc4/3llzk5mbWcDjOXM5
0/3PWPDXUAgQktZfa6AVSn5piJf756iWlmD8qgaBF9N1Ty7vI4UZWir67Q/WJTAk
s7/btAPFb//FPL7aAJ0MOP6wlB0SxJsHmmLuIbj3kheJfZZ6IQJG6UjzPm5XRa0H
asCru+kbp/l2m9ILC60lMQnnDYONFKaLGdHdSWvfhgE7OdgeLZ3fOau+BtxqaqQq
z2wLWH6ak0+hXIhx8/7fSOVuH1VrOPtxWR5X0eMn4oPe4FuZPY0/mOjaZ64MaQtk
1gulyRwDBcJMyjZ/uEew30lsyrGqtPHNTbtH7e8+p9Af722MCZoEYSQJylgytOMe
KXg5epqR9gaX3zCvV+6yRA9gI3e5y3b5lKtUz+UP3upbekp2NBMegOEXO286oMRj
LFYN+brcK1njYzZ386tMZbMoaXYI/f61C3WTzy1NbxOkuTaunhXVQnF6mTM5zJHx
ykUDDF4VWwkA13bY7+EK2R/iPsfPiG1LhpAoIJTFSYo6VS7V7xBjRwFITkh/tEZ2
utjYzFrRTUogl3hqtbqwVVPpxToEc5fXJL3BrWLVFM1jqMnVp4b+K+U3Lx+IwYke
D99pzcK/n0LFrAk5EOb0E1FNlywsfILwq19HwxhQiup3+QxwX3mLlPI05ZmhHFuN
h0krOz5//qSdhWtk9EpezrZaIIu88KQMqoaE2CK0gRzRA8EHhE2JYZfLEJH9f1O5
VVn3xV/wRmCKeN7fJpI1JNT60lm7hIDnJJg5SO8tKB1DGBZDa1S+pAmU9JQSG87H
n26K5jCBBUXnZ3vd2VNw7MXZOzY3tDlpSHDtp23u5WT6mmMKLbKM7YZTQ+Atrrba
QGWvdQJmEoZFrHbVIx3hVObF6/np/GUcb/krdrAM1DtIlrve0RPLEp9xFV9pqzm6
d82KJpH1cMp+rpN05GA2UxtjvKbtEgxYdSO8Y7OXZFZE9Pfo6x9rTYdjHHBGtUfV
DD2dcW9A9EKoGBmDeTlkw4HhpWhqAIA90xml+blnVbKuw/9IGlHxIAZnciI/UtFL
8kZ0E1/AJI4ezEB9t+82w9lTaZXUft7VD6kterJpp6uocGhi0n6zXjda7bIPz96y
kKPXdCM2NaKEFPYadpEZliT7gXsSSW09gz58Xr9x647nbFET8eQfaRjGOFeOy+yI
vbom3kM0lgnZ2fTerEcfkAFSdrsA7pxhKJC3DCdLhZrljQqyURoPGONccTCnm9Bs
x+ugxSyuJFwpvMZCEnLwNGygQyJ3uIegtbk0Ovo7dH1Xxus6R6jXqILp1+TK0r5K
Vuq3znlIpugmsMjpGY5/87cCz0x4OaLlZvqI03ZYfNy/mMhnrCF2NrRuM05Uzeju
qtd0GFrR81DgJ3/1ScvhfEUl55p7wsZbx0QQY/ama9XDkh9fYHP3LqNwQluyUB6g
vT08VgPqMRfnX4UnVqqkqvhsgAEyCX0OtlloE6k58dMZNZgQH1WC8IUMIa/AUu+n
ZWG6h8zfH5WPwm2QeXR4a8luMyayQN5YwQG6MDxbopk5SOE5ttB3WN0jmPQkv3aU
SOnOEDuIb0GIbk+WeJn49pphnPSbhUJ8nJe9uidrpkZiqcZ/gCGyy5WvE6fEiSLw
PGA/W+PpRN4/5MZ0S9VfRvCRqFZFL2e+R7MDodXYdXyx0KO0NLFkeug6UnR+59Xd
3oamHNSh3vViMk52r4e/kH/BpH+9vx+bGWWDuaskvGZ6Wsd626SLIQiqs3RvgCno
80SwUO3RQDiZiqdpj3GtVmued95cajjCf4+JJ3f/nLAZ7SSwE+ZwHnqY5RRZJQdT
pCkoBD4XDEQNJjgJmaKQIWGkqfWoJNHYiN/YlMjl+FMDX+fD3HbwOgwEfQlanYYC
NTFGH35Ze2dAlO7XAQMwJzaZoeIMGPUiTsmm1Qa+MuhrfCYYHg6ckRmpxZUPIim1
goSIR6DniqgiyQ1F5XlTY+pTe9wwWBcPZO3q7VFck24qhEYPhCb23OunlPekn7Y4
2DRbKLt0q5HtDURgyhL+cW6pJLwow5kHrAag+rRW5Wp7jN1QOMzsWj8y3ar2Hbhc
BXBcO8oHV8062MzhZKduEsqoFt1wB6SyC4vYjU7awI7UL6wSFuSHrHMH27Yfv7UZ
AHzfxJEzkfU2WnIGAGMEFIS3k2dxdVACfgJy/agT07i0nLRejuMEiHrw7FAUqxKn
cqLtC0pH8bKCW5NAOp3TKmtBBGuxXf4jzNiD5K349UVotXdn/05UpUAX/xoOi0A0
zg2d3Y5Bjq/LqXxkmX3exM7BKoGshW0QD1F9mYbN6kLB7GqR5YQdkoukyd6Vd9WI
OSc8pNm0ykfuDTBiMdyCIfEAoDdOwkXor8kosg5oDHs5ebIK6HFCAK/U7jSIAX7L
rzsfTW66j92wWJw3h8ezRhacp3h3y788no4ZP8lqitg1LZkJ0qRRIv86XJZrIGGB
FP4BBk1g+4h7ZV2gvI/CD78KTc73zQlgOxShsmTfKehohE2bKC+21qrnitiP5U1x
6DlgIyoj018OSy25RdB8J/TGAdNjC5uFQFYRKfaCSeqhJp91JWW3zbtSnrrAoSJK
wN1rdBo5J3IEDwPwaFhVdavBBQi4S8LCeAbXDtfO3ZRUpVOhebHnvkwGYmZ/oF2G
UbdzJ0rv0J4OewmCV4kdAuZcOw5qgCTOIWYWxEEVJtWqz+q8vNYk5M9QvEZrZMJO
iun4Syt6R96+lRdnZz3w4WON2Ahj3Bix7YILkzOUYDAzQLG4yDbmonIqsaum0w0L
6HG9fOx8Qh3e6nEULbo20P66MR9GqYFFsUCyyQsyninbgXOvdJJ2QvsDixjbUpge
T7/JK1K7eDPyqVL/HCyYfLn91ZtOgAk/ywopzPtFKcUMCg8Wjm+rri1k4Tp6r4W4
SG77/vBSuYKjZEGEZhb1yzLO0I6kwETbChSrpLtqADMelPGGQws57UuNed+SWGer
lLCSLhbkgCgeuMyTa1sRF9KKSJ3gz0pc8h/01efQPm0MIvZ8rYlhXqOAP1VXbxyW
z7hcUYS53m7QRzkrS8jbQkZxoYGNj3H5gAyp4eZ4pmFhBMTRcu0lx2VatI7h+8FA
L+GP6TIPNw9lfD16REV/Cddje6sDdMWn3zkECNp6FAuzkQ0V5G8l1WGt2llaFsqX
BmEpA+UYOx+17r38mXQ8/TPTrnSQ++gZHCjT40qSQh0PT6esKqn1LV8VVpab0SVR
EsfrQXZTL2fQZcw8EKHMdUiW9KIamfAe8YWFlGQyrmAkpqDYAMwysW5Bfb4ypjJy
VAMhxzZuFxaHl5t7l09ei8N3+CvoCSTPPhO/jbRrNCbrRPc35ZNtSaBYv3vF4McX
z9yzOT4VnZJhUO8Oqw8UxNAniKxPPdCY2q/LNnAq+uraXenkg0INb6vBkgoxA8tQ
m4OrdS97BNg5OQrpeXhLSpFEYq6otc69HrTgBiXKj1u1q2kLk7iFqNkN2f1s6t+9
8cewHf0reZyMXAJ+s+EUCzXFJ435F4MXqzzQ6npqGs8Wdcknh56kIxn4BOzrcWYx
VDpDJmme4ZPrbWVcMU/GuQ3/uhbxqGt16SqfRbB6Rf4rnYXP3SkgMYIDHqFd26Lo
epYv8YrBa2D0VK+fkHosf+W9u4DVN4D+NDl+IeatcezldFGJJVM9VCE93vs3UBkv
RzgtR+FajGoYrWhszib3ydpHelrzJ27Qjc2foABcTWxw06lnlSTnSQy+Sqjl+Rzb
nxGnDYcUMYhzWFFINXD3KLeUchI5r8qKy7GYlRTgGHC4QDVOLVDHEHAZnWAUN/19
ZAtmS6YGE19OQGqrrBhHCphw8OMmmC78O+fEEFxlYogC7RJJjyCE6Fz/BpmED7GB
QVV2HohqKb0vm2diy+YpRnpSrX5YBy59H/Y81+7GmeFVdmzNVHxUOfueEmQy6ZLx
4UFiKbSaJmkqdnBIgbAaZT7oTU36R9hfI6H2QFjluVPZTTQK0JO7ivMguZ8AacLZ
b1tH0aphvXdzd++r6z4EYHjIlMEyRdorHjy9wgKjhd22Yb//muo0XwWBWZnES8iD
Yk1ghKi34mCa3d0u6076QVGfh2SFrN+JldDieWNaF7PEBIi2Z6H/LCexaSJWuLNt
fWnnhrq3NLgnuDSj79+t0q9yByY4xHKeIGhOWebvKv5nXFqOgB2BCwV5vecao2Ld
mBpJRoaub7VP1b8dXWXb2ivnW1/BPazsVLvtQYPM1XDDimarjPhdPe3Us2BXhQHQ
xHjtZ9mIb12k7671bJoyg49tp8TMimaKPeSxPem4jMahuJ13VhjhxOpibdEFhRpx
gOlzZmKXZLpObnFUUKcVifyV/NiVlOwhLALaBcs2NbBsHDtp7IDzz7BtzYVuzHGJ
P62R9H6GeFefK6vclxEKPb6xhWSfjoB0MR7cWWAYu0wr8t3nrnOxL6wDWbJmuSlQ
yyR3wPuKJxZWS3/G18O4SHo3Y3BPTrpOTvYdMvEwaqhIARUGOQWgCBX5oQhDtlgq
sLw9DFHG4r65TUN+lRQlLdQAaDiFcCwesUbMYzSX+KacpXnCq5/Nwbm18JnsmRrg
hCkjZ9I73uecuAj/xUsRTefmwUmS0Ubl4w+tZAf91TDr2gSVliefr0o9XHBSyhS/
2BcJMlyf4jM6CY0X9jibqqRGhKJ36MYF916vAu5m42rG0BszQH6LKx4aezIVZ+5u
J9gir2soyEUB2PbC1+gtm1njA/fTc+EPMvAaSiDPuoAZ+HYxVDC/6gsAmjVvt9/v
4WeWMIQf+hq2xFpQD0W3Dl/vVZOONcV0EzSqMIsDR1wmXhclgRWebyjzid37m7Qz
rxSVJOzqNtNvw6sVJTBrivxRuIPu0IXr2V/Rmhu7qCxztnDtP0dbmxFouatwM6kR
QmeqIB+DEaF2D2rvJEAb1JkyJN/LPEKFmdG09d5B/KlUjl96UVweswfNayU7dPE7
FZcuz8VOloVJmxNBEEkJHPR9/LV/DyZpjC6kBA4fjccOIkX1SXgIiAS23OCjjGww
KbvKzTejm8bwsI02NRPiU0BOozlay7Y/rz+oKoKxP1G4GHn6H5yLxXfWb2oweOw7
OnfABcVsZVBycfj/PYb2ExQLqwJHF8pfcLc6Jnx9YmSE0d/XkiPaZLVyKaxGzQIJ
GPVRZD9U3aM0et4SJ0Waydqap23sysCUDBIbAoUR34koJA2tbRKB4SMGsrObGqcL
j4mZ33QVl56nKd+uOryEOp/qh3KMmYqZRXUKz7MTWCh9ihWloO9OpUKS2lKdesA3
2xAbdLGVG3pSM/QSKXvU0+Cy9YqlVw7xj0oZgTGkOWdktz/eDbdNR+ICqWUZ2Wul
9qjAcaau8p7jh6iMw2nqtUmf7uRuZ7mY+11GzNTOmQ4zlAtNl7TcHtsoYoBcMcxT
nK3TOOOlxNnGAO7qj+QXdROU5GEVTQcyqaPzKp84DxdYWSVhGPg9LNjqGOFS5ns9
bZpAhmQ8kOQG2Ce+SSBXahE5STA8A/EKoVx6IYjl5RfpPS/Qzjpoak8jeqLFashN
I/rZvn7fECr6+1TZwZt8FtN+/dfaqcwX0kH0Ad59OcZ4xmIbJGvJXbZDCty+ya7o
nRl2S0s/tGvRNsaYD3vFzCv8e5cJA3tdW2eH8M4yZgrNry9uP1U+6DUO5q2jF1VI
4iex4eDHHWJS/M7z7Nc/DvfJQ975rOrfJo9aDShSoMpxYV0BKHwTK0k6B+7DyDNi
mjsnqMgGtWZYmhYZhWvZdZNDj9xsVta2Dxt1wVCR3FMTUmZ1nUGI7Nume7ZZ0VGq
eKx2DozUc203x0ekszCj83a38fvV/VNtXLLaXdstST3MsbVrq235R3mc5DyHEXtq
3H+ckgPe4HFFBjhjLfyrCF01ljJ6SsTYlsOKSaZeHhCFo7j9bWFHvP2Ghx0z4c7q
LEH7g3ihfvXH28j1MODYaENIIow0rMfagfQ/w/6ZONYNBEyOYSbuGEqTD1inxFYK
10fJitfYIV79xi++1xgoF8JJUYNAiF+kfDkzNCIP3vINUD46NEB8Xiww1N5sMJlO
32tZbMnOWUzHyNnpvzso6ZQPNGdM3W6P3PU1atbHyy8mZgLY3FGyOBI8je5LPHBq
Rfm3jZscV1Mlb9Ow0xqgpPFYvr0jTutPuwA9b+lLehu4aXcvk9+aZNeKkStu+IQl
czNwIO8127EC1ENQkZUb1u6u4f5+fGF/NBniKX4xYNkvUBR4UlA6s8ZXXCHe3sKb
qukOPpqy8Lw3xvEcHTeBmMNNlDJPBNYzDVqEutBk8X7cmlXOdyEERC2fIpcrFCV1
pNc3pdRQPMSEKn8Z3oU3mmo6emvDsJ5qnViW3IcltTf3rT2l6+5gtggI78c/LGqQ
BxYvHC/piWc4HonBXjxjEQfxWZS/iAAo0wosZysnKHREVgtfSPPFkL9YxNgDj44Z
cFNixvqzqJOp9OUrYCcJI9TAD30kmMr59UivdC94LX7aJOq6VoZ3zy2z9GNOZk1N
xIafm8nCE0rcZaAk8F5KUvprIS6ftSwh35COo8hzjRpY5+Lioe3PeYkRNc9uLgRQ
fzkT8nxcKZxmCmjJ64txOwvICgQqeoWZ4QHOUGZ55qTNGHEmyathgtKiOgG1apyA
6CQFI+z/2zN5AnAeEByddfmu5/vZUauhIBwchWixM4OqwybI4M5FBS4BGCTQ+Lt/
bwVjuqna84VgKpkCiO8v8Ej9vaT6d/tlhpProw0hO3SXxIrHk7zkYUseKit8zFBu
7Ker1g9+LvFBXjRP14gb6gCpGu/Ekmw7pKHbkCJfTrf8DMAGAsvNupclPY+ZsSYk
cIji8qfFV//6q350BUXAKf5jAWnoKDh3E6BJXm9AjWACFoRnkqUTdH/BXXgPag/e
4h8aRj2ltVUqy0hjYeAivEYFOuwzd81mIe9mK2W/rFQ4sW1vGVHORu0zEfwYK0Le
R43Yy9Mjy5XxB4EZut3PmEAJdMHp8o+MqwHUish4QOcPakvGLPlIK/I7dLpAvBhB
C95ia3KnDoOWoYUDIY/oIBqJ6qL/cwJlON4L1cNLXFXSKQ2nJYkhFUXHpN7S7+FL
pvAdR1T9YJACnGgfLskP398x5GgFeaFwpj6EJ5OtjTtrk4I2iJOoYRydOjJMo1Bz
/0ypRZm3TWGXlrkF7cQWGRminxRbObzY8QuGIsAJzZ3b+5rA+81DjoYYaZqkSBtf
I89xAoxoYl4mh/EzZaPPri9PAH3y+vEjv/0sBHp3fSI8oBiQSypVD5ue4bg2Dneq
N5I74xI4mz4OWLdcPMDN5TTcQq6bxYetjGtXJfq8VYcOkvh/zim5KPFJq1RaYyLs
ZGNvsbFSBeWK5vUd3gBMECxhL9dJno4s44BCoBhVLsPByZQSF8OKumc/UTV7191Y
aEmmOmhf0tbZlOMBVoyx8hpRL9+E/dCZqeFtmAHLWnb7p3iJHRd+P8/bvKzIt32Z
LjDQqB91oYXmZVPh/1alzx6aIfnPTGQugIt223FBWYrNmbPEdtsZ0E82Gb/C+jDd
X8kw+IGIm/dj5DHurksxc0eBC3Erv3qKGbx+95pYfvE94z2Nq20zqYcBybULQ7Fs
1sAIl+DTCB/EENSAGETXuJSvleZWzeQZ5XCoF6MAFBaVxlhO3aJXB4Ngr39djVDh
aQQBRa6FGxRVTZ/4MbiAUgE66g+UDrvfykwLlq5yb7Y1trmVIZnYHucTOjZd60vM
YUpkN/Oa4GzgkeB/gAubme2H6XRDQvtqlgHKg/+YIIC1LEaD0IIVla35XCpxcuvz
68n9nN/Cll5FPeBKjwBamcz2RbO/XTCP3Dg04F5257NXJzpFSgYWPV8AKFv7XjNZ
ag0v7g4FMdw5FsLAg7f/MFoY8JNV5LLhNE4nQz5BOdIZSXhMrvBcgFNwNce7yRgW
DyrBgaIRrpdo+U1nk0VoTatLhzMCR/QLKGbobTdQ6Vi4tX108MYa9PZ4V1v76ey4
yrH3YpgYWaF/w3tti1l9E/KHkNLQs4jDFIp/WdmniRbJecMYZa8Huz08/ZA+6Uje
2KRMJrto/UiR3q9lqGz1czVDFeVkMoTJREdy9PZYCdTE+jLrc8dQA4Nch7II3TYq
hq5ACcnHBSg6t4JBTjGStpicUiUxa2twvOCSQKvTHktcVGs4Ju4hZyjtLngtSBOe
/ysFXqOmq+hy2yOlSE5/iBEy28SgHYjciRwQbDZ4+Xb0mtPNhlSXy6I/+AkbwWwa
ZQ2YcVeNl/iqXW4J7fjmji6kIzAgFc0bLVwbdtk2BjxZCoLCrIeX+QLpTyB/M2bd
pXL/YXGRW0rGTL7mB8o35fUF2Yg/8ygvm2Qr1O9d0Tj9pim+F/ng2Q4YfhtFE9nc
a/Nv3b0nwjQiz76VrRh3rKVRZE6brxJ4iPj+qzaOeDwcUonzHc8FFeJJ8Ed/kMNZ
/YjEGYme3OtvjQMsDuKpXHwbt47+paTnIIyBAffPBo4P/ZDoy7I7nfw7iD6R1rj9
bxHWtw2SgHYTYRsoqqWxthLmHUgYSjrqkdTQwU9xtNUw5KSOjnxEoEihtCVDye8S
O/VG/HdEvc9zdEySzwr+WwNBxC1WOw6boh2GjxVFoiT0LtBO8TojYeNUvCxTNPg2
1lAPlHDFWXmb5MT+cCjC6dxe/uCKZbdZ9zC1qdyMfLo11P0Pdev4DYZREE7eOXKE
TadxtXH6Lb1or89cgS353mUNF6SpyD29+s3fQFGYhMQ2Bn31CCNzxGV1TzBv1xFs
9ngNhMh8wAOiFw8XUFsYRiW6yUNMpmt5vN595O2feqmkVPnfZAb5H5mQorcTHHJF
yPR4UbFnVKATSnsfACuKY/jg6IQqA2liz9GWhePNazMr+hfawJilamIPA0c1P/V3
8J16Gh9P1JPs3IAd6fQV+oTgC0jgQGPPEsu1SMUMB9+YPLwKVLV1Vo4in3/pROtQ
ZUnnexUKZqsQOuofLuR+e8yh2WEuuCwNO1XU08T+kAvebMltm8QnL7ZZ81aI/wQg
ZT60JUD9wO9WBrXrZ8D8DOgmMT0MXsnWzpB3z3mnM8PKRGfBGoGS97+LoVBkcGbi
4qVZln6Z3l8BwgJXWjnumKtF8tyRtmDR4EQcvUsM47Xn4YkWbU391PGD+OJb8SHG
OoFzwUXyTHni3yOSn6eXk2ifqTOiKdTp/wqrAZ1oJV2nXfh1CadqUEXCjec5Fc7L
BhrEl8PjI4aj8fQwAnaCuunTYCLI48XzjBnsPvfPNkKMW4jeJVTTwjHAqTNkDHB8
IKxLBv1RrHPfrINwAsvQ192391kzoUYEdnRz9bhg7czsiyE+uEJwXGedmKNItehJ
cRsM8zSwBYTgWPaVwNWOhKH44EzIP1DfryZok8oQ2RjWm2fO1ZlXf130qHov7afr
oz0LAPRG+o/1u65sRZRpKjTF20S89ZRO7bV7+DSHesqEbHW6OMGmT+7qFSNqtiiJ
v2OYqUjkH8qUwXP33L/1OCATwm42RqUacfPoQ6AezHiR3JWRgVtcjpgtxa53eUYe
v6Mu1saGuW5186PXvwXJHquDYIrn3I5LqT56MFyouqZOnzp63OC/IZ2ssLD2c0Hm
iT3RndllT9p4hpEi7whJVIc1U87wMLcOXLu1AEEbdxrEfvJBZOxznOnqVBYYQmsK
ovZ1RtgwvIHJWvEFyviyCPy/iF3dGt+m9QiYUFr4cGnQa4/2KV3+2jy/CEiPFa9r
zGaPclxJeZ1/hNKEeI9WLXGKC9tjv8UnJMCWSFaDqtexzLvClP7U7S6MUZNra0zk
RJrpQUwdkmW9+wmYIf+zsTbJ5lvHnqd1utRdUWDkzJ71vv4HVPKjC0EeaWG13XQK
KR+pMiRa68selcNKCeCsDtJEJ5RHn40X1vbcBgdvVfnidfGdp8TpNL0MAl+eu77k
xjX0hL40Dpt58bgFU+tcKsyjlyo2um5qIwh2QkNL4lOmQa65WPZ8TCPbd6Nmr0+p
YOJKbt+VwQ2xmSM9LyFA6cgGSzL8q4iT21wHWdi/8OJCw+bAE8hCZYpsa9rm4nLR
8M7vLvWhcVUmUhewpP/Vkt5WEZyUFKrj/QByDwTJh+QSRmSMYt943G9oFOGBicAS
NB5EbuQ8MuF/f/qjVBDzCot5peYBF015jVaULD+54OqJrJDX0ux8DJscebNU+rmD
c5YDld6w70loDnFSbcGjfnlhgiOuC+SY1qTgtZwsVRaf6Hz5SBz9WkXA/2AQJ1Cx
jfr7I4mkJPshrmZSxU6CNQXmtZzQqzJOgPwEFXF8OaqQzhCOkugDVZvjHqySzxRY
xVcul8JN+A8IsfwzOCDLT1U1WO9GiVE5u+zJswLKtHAvN2EBl0GKx1nFQprhhqva
2rKRBR9mWS0K/SO+qr6YZEuCit1qN76gN/dwAD8bd6xSR3AnNjLkCeJL8oWLnzEh
GZSZiorvNca1sr52f4OksuqQ+bZYJlqOLUM8gmUFAddaV0QEtqg9jmr65BwdVrBt
Oal4OXQBiOESgjB/y6RhDMkOjWQ8THc0XBTNr+EmtZmgN8pnmcQ9iQcigqeHJub4
pqMfG6gyPgrneTubUweU5kGo9PGwXh583nzbjawRRyYl39JEWrfMzceaSzOUCN8S
bo7xLpdogJXjJkGzZCdb/dursDvNH08YfzWGUo4lRqTcmHcBCGvjEdfk4cJxOSTA
lo+9Zoc/gE+vxy18c52yJ2jWV1myAHy399tnUTBHLWwt+HI2HyFo65OwLsJRWJOS
BFKIMc+ecKpyOt35M6wC7W7484WMWDaxlZ6P+qJq7NR628PgfxriwuHfW6Z9DhgW
rKeZywLWfi4CkkPKg8CxehEkt7+m5gqFTMeG4z/UjgV9MFkFFCPAd1dP4lX2aryB
2SEmNFdH7FSORJ3mjm6H89kr1/xCI7tGoJZHcVHC0zPtPwrgN+AvH/KZF3ZDsnJX
Hp64vt8idX/u/AdmdfypPJuajYPMum/izx91VkMSqSPcaZDVHmqX1mmq0ZxuiosO
mNI85eKsRYalo0aabwmoLM3aishsar5LJxZVkgKrpmxOA7IEySues2RsvP11G0hp
mr4ppG152zgDeikcnPAAekRdFs++l22tM2p1AbBT/W70GsNnWHKVJfEibv683J6/
PSkOHuu9yXNczB+xhdaHKVr+Zkvg8NUtsOp3gwo8WyFJ1+vuCJ2zIvJf+GBT7N6Q
R7JdsrbPjFcC5OFWe1uaKKTmmwR2sNve1rWu+QPCdzHfAJ1BYA2jTz0pWkaSEBvt
uH/BTow+ST5f8D3UWgsnOuy8DjCOy3Pmxi+FpHrJdjpmQ8y8BqPrp1bc4Y1Pb8kD
TEyXdFl7YHLh5yM/OxvDR33oshMN2lXrDppzGWvIiOIZk7LR/GzycSx1jhDfZ+1I
vcOQMEg3ySvUp/KSfi0QEQzSZTb8eW6jPsdhNT0C7mM3VVsuAAoaxvnVZR2qtvhi
ujxr+wEQJwkWQLhwWD5JeXsI/3fIPUqg5DUu9Nx0h8xIVF/PzZLk1mQ4D0tQBowT
Axhr7HVDOokXEp95UXNziLrMtoKhjv24iJKBzVJapQwtcGavMnhp983S96axj3dp
tkD2k6s62r8/fgxYb/tzzK513gbbQlR/RVPixRmsrRgjup31jRjUNh9oKMwqTql+
R4IfMs/eIy0cPouCvqBod6Vtpk+gNsU5r9z+H3vQ4k7TaQdbl4v+GV/5yQ6LZ72g
EF+c2eirvB7l/pLcsPsublTGA141z1qdvPuvtuiF6ueqGBde0USoUuX1AUKZYI31
BvdKJxkZ8+YV8FCBycKVMXrN70DizGZ4SSasf2Phty/lbwrvuX3BczeSYVXhNx+w
Wks5xc9o7cgk8YAohUpaqHu7/0DmVSYbFNu3QWLhirGr+Vkmh3V1jqxcYVe2y2A4
Sj42KkA/mGud0VUsF1GyxmCTQFQjQYqCFriRJluW34uEcpAW5q732M+2i5QMJ2Yl
D7tPg33CINCWfhjzqaPFbwmCXo7UNxtQOSavxWz0uVxNTkoC8i+HXcMkISsio6rn
Rn/ykJ5xEgRcwGKT2HSZB7JMu4kuxGGfOdozxrHKQ3FjQLcKxcyudPI1lT2E46fG
ibzTCPeHZOUhwlGi+4e963upIhvR/d8e+44bhcwisLxbQQL8UpevadZ9ishP+J7C
HPY3mgqsB1+9MXhIVjTvZ4ddkcFk3vqiNwbML5dYWnQDsZlmrFt3LEQ2SJW8gvH8
QxeokSmKN/C+W2ZD0IZsxFcnQedTg9WFtA6t8w/UYG94rlp53+/Cp8kr+QUzJeS4
BNzrBOGb7iZ3qqJBQKSrqBnQfTZFSZrHgxG11RTRYzaxeIlFkRXTR3R4YRLAGoqK
CFNS6tOO1e93iU1pkN+4RPTQ3qM1wOm03Tercm0/3/XKLSW/Bz/A0KkZww7Tioo/
veizUDKRsfGCV/6SJQXoWeP5+sz3gLPN8Ibnzqg1giDen9OXJdiSfVmMb+EQ8fFw
yTBCBkK1iLEIfbZrLuOjyc/oXP3S8S6ojncXqnaTYQYFXzFPiZOsBlUYJt5FmL55
DSVmtqX78qRQtc5VJv0AVmVP8iocTLjGajBO1wL3bsrTVHUtg/VFE1recGuUJups
QV/Ezgg5WaAlQwe3GT7o3appQtbyNbSROCtoZ6i08blIO2//RpECj6p3moXGHEZg
wpOPA0HjJOr5OR2IQ9++0zinAYnl4T5AIDZK+lokuiBXY0pkjHe7u8kr8tq2Ity9
ObhixgVNbAwghx1BtdLvVLV0Gu6ZD2u08fZuy5AFGylbFwE4I7Au2HdpT9+QttxJ
cU3rQnCuMRQRjmpIi5TptWX+GyBeFK5CM7v2G/IxpQZd3XEee6NnzlLaQzVO1SY/
77LMQDkPQi0Y3xu8acJ8pkxLx2E4FEjkQi2WBVSwH0CfYPv4X78JWnN9BdmQhvNz
l2vB2LzQsi+ieGotyXbeQRgv1Y4v0nHGv9vttIW6hf0gN1TN6l+/ve1tuCKepprP
52Qv2kBaH1e4oJaW3x9Cu9Ap5v4xh0L+2qL4ZUzIkzBO2M6uiIcHI5i1cNAeFOEU
Q3OCsMprTIifGne+cp0ovvHYbVRgKhnL3ljDN0Kh1Rgd26Bhs5kS2NZIs2rnzf7C
6EBw5oowmjMY1pBEpgkGFWRKkY0XLpFah2XVXuP5E7msl51kw3dnflUPFIxOFT/j
4lRZ+MpE14yyu18UBrTYKvEknuKZcR9NEgcjueV0rzjhJrbH9LUOTcRgkarYv1G6
ar+LiJEBqoGzrA+8lQkSy4kE5QYIxDEWNZ8/6z2gUVskw9mrxdObI8GPoBnYtUnU
DXPy4CcNZQjn6XcHNZd/me6Tor29cn7IfUxhSqC+VD5wOb2wHcp2kAvAfHjwn/6a
SDXhUjGbKhmOKgBSqn/mQ3wcXtC1UbiCLlsjmO8HQTrF3i271U0C7kR/uHLJiK2o
+SDXKwWyRcDDmH1fUSDQoJS2Ygh0gYVMdl2VgY1fpWzWGwUVWlkcKqT6trcHtUSF
0E74IVGGe6eM+F+8kgRTja20hYIwe2ovB/bes+0Fj55IktRsdQBEWM/gSAoXGmXl
SZr0EDKDx9LmYohWnnnjoUwbFPwinT71uMpjOdXhohIjH+mSBrOxw02z0yw3EQ8p
LKK84kxFcKS0gvjARd2dbWc2E3Hu2Sw2i/bYidSYJPRUJD2fi830l3TA2akB+/Vm
ulB46cID2FEWJuUsaOjtLLgtYWuOTZAZ0kxTaLt25W5bmt1rI2eSRTIoINOR8Q9B
0Q+5OOQZsM5NfwsAdSfVXwQHMR7LYI72wYk7O3QvF+nHeyOLK4wpd6YTBqSPW5JT
5AQ+7gsQDRlVpxV4iHGfOMpHU9pO7dGITT6jiBdhL/dh4k3foAdDORAhfaL1unrB
wh+QiT2h5q9ObV1QUZjlTWa6MFVn2Rhu48szERL5YiheAA48Q12P8pipMNeYQYJ1
2SdvtJmwouAbowx/5K18zplQm7xB0flztomOgWF24Nw8livFw36n4CeSO4qo5JYG
RDs9ydycyCGKm+P81xE+zQGCLqK9gOwhGbnwYF1lk9wKzhlYRIHMBER3n8scy6Bj
go5V3o9BhIp1l4/E0BD0EBpO6Tex+mkZj+Qpp/LKeNNzuV4f8mccacFWy5udXEwN
FlajuU0ghLO2/dLFBYaBP6CJq4SXxyFD4X+Y6JRjGc8jRqUNNgrnOzm0B8iEqzo3
jeRjefHiwoozdIBMO5fUozKBcB4de3ov2On1T7jgX+lZKs7A45Kj+KzXe1zhb+IH
8g7QcTrR9F/S8EIyIQ+AoNRg4O50Y8nctWYbPVb57DTr0yXxqIcmUepHIYOZMSW7
+l/EdW6xLxmGBGK51+2b5T1mGql8HrdYpkQDaBzzd/G/ZVd2V10K7Thi3MsaH2LD
pc34pObPViB04rP3GBAldWNtRBg2fryRJMxNMMFO5KelYVMgcWpbhlogktf1iIvY
AA2YBkfBqcGqzQcpp0sDIBvQBkLVxizDjOG6iDAwV1JHr5yJHr/FpKYfMh8dOGhs
eo65w6lQzw/+LHZWB5E/o4zJJGbkdxOfszFZiD+iqJO6PDHiDjwxymlSvtyslOVJ
o62ae1L6LNZHojnA3Y83fK/DES/GZbvsixxA6+73/Q1cgzMegzU/CmwVWYIK1FOo
oR3jp+THrWC5NU6IBMUCVtwHOUdZgSCk2KHzJQZ9xvL3ApfEKaLownI5ujc2+cut
gUeU9JqlimdfiqqhR8FQgFVwsVIcynKQ8C/fNik9OYpi5z7FJcdqAAV7Sa0Jqy8N
X93TB+pePZ/DiwVy2aiZPbcj4t1OAl+m8I5G0SWJmaPgBFpofjvmR6D6rwI4ZuLl
kEDshkpgeosHpU3ziQHS5KOnlCMopBOjgiV570EX4ur+8xlRMZFLTI2oz8+8b6Gt
lXBVu3Edb7ZMgcuz2a0wnCTuxhQ1+n0DNv4ZcPwWvVzsdEMnhL81XkkIlCWDFtwy
xCJ4USoHEnxoCPwPePrdwv8I3Ldb+0WsClHrmhk2NdQMW/NKnXut27bQOGvK70nm
dlLKzRBkJiEM1wf1WreJSgJX7v84LFOni540gLzrpTUxcrhRbo5BSCSkJLina3EB
fdgka5sfCqmdBMJg6syB1PPevVP1/+U/CDcWTBvDLwqKPrF2kUXIZutt4c5F51qQ
WQpkL2EKKfsATaQKv0f9+PZ73UEg/xyNa0DDE96zsfXMhtSDa5s46j0+anF43AyU
X21yUOOiCWDzAjhO8EFoCLX40FIGkLlCNOcooVVbM+hQDNoWSMkxJAxMgEzcHpCT
ioPoS200eqX+YBg7QhWxgDHTw2qC7gDSmMci2YYXU3vA7X51BOGGvHGfwNI7AnXa
QghZjl5NmeFcQNTT6y/le4LoJrbNqf4KhWLNcE5NAocSrIai6NNvgEDtVNu3juci
KhpQNbLVOZjAVSY6qtrWZWJ0zyqIdNQ83hBPd4+517U93ThAmeuScB7xLsj9+XR8
DbJe2FXxKfV9AIwzjd7md9sAaGq9KTnVo5RGQDn68/vgShf67002tglCNoLLPBBM
Q/JeMj+VpqJAjSFOBZQK1s4U0KhamIstt8V/wIj5GT7+hK7zGkrjiLhye1912Ibv
3x8+B8TFaMnSSlOfHye556sevS5ey7zFCIqpEV7+Qu+xy/YYKeeXOmjNCchRAOug
vUHi2IksKzqtV2WWlAbyPXqVE6FnCvBfYbc/vEFPrJZEL4ggXfLja+A+5/3lnYML
133ZVe609mtZHYSoiflxofhZmFWF3W1Jib4MdIrUljzH8j2v8ZyLz+95QPxwV7fe
cABHpqvp36g5NuknkHy4q/gpgye7JsukwDcyd67ZU8SV0JbK+tzXXzKvfGCVp0Qy
LU/qydHVf9SVymmzVqfFGM2P8sYKkyfiPuoY09/Avz658T3WdLS/xPgQeEK4fU3j
Q8Smd2QrELf9AHN6g0fIVO1/hf7k2EBSHPAPmcTkVSGByqEPv8x/peQhgMc8f+5L
H84JwTDt1JAQvdnBCBJgqwGpXhCVO9MCltY1mvgid6TUtzfPs6XGlKw3hvfJdv64
0pBtyfHM4DatIerFXInsABNqK2HiC3a1YeMQ1tGpsqycpf77wKwVVa6w2W9UAgY/
xL1nz23PCYiWj91nuRahaZZJbubayrqkszbHpKZnJBwq9qij7KTAWqa1y79p0UsD
AThR1DaCuzdHZNn0JTD12LpcE1E2tRDzyJtt4pmw5AHnSvdha/u+dz2lbXLgBlB3
NUfWBlRGD4XMvJ0bmsWNakgGedz9YpNGbPFhevB5XI1xSxjLvPY76EV0HGL1yQvD
/c1ipsJRYmO5xbGJoYGpDvi/3K+9DU07QGrFS/0yLASS5uUoTGBRvudRmYbsRUUR
btOsSz0JCjpgDhM2kyHjnHiL/XvPItY5CsRfMsMgpSCjl3SkUURmQQXL+QR3f6B2
zWJl1yTWr1ot4enHn52M+6h8R6iCBduEf4QYGtdXWoP2uJtcoiIhus2uRCO2l8gN
7Gjx2D8yZr0QYfxRJK74YfGQhlMkRxxazmsDELP4y3cvhD+zVIfuyQkPpzEo6DI2
e5ayoc2uGszHLHOSym6sc8Dk0lWHb1LFiM1K6ty1Hy37RqJC0PXg/QSoghaZJOon
DV0LiqQ/UEOoV0fH+OhK+yAxQqCnoOIiiZp53tb2UXE60yhI1vyec/XQJ8PDL56c
iCnPBq2dIgTfp8B4RVrHLr1PVztULaYyG/Di/0b7uzHBvBPtnXSrDGW6Pa06oqfS
1V52SOH1Ivct6dOvdMtw+W3ZfIZTNQ7sqGCMYDzWBTW1q1V4rYq8fk/CtnPYsC8O
tMPqiA/qngbTHbt4FFSd88+mqv3XWdsXEVa+sMDHL7McnUxqsOfxI7uSFif3PXLo
qC7yCTZq/t0OyxFftVC+mXXN97ne7s4OyYlXdZZic8AE9BCiU6S9irohcbHWVLMc
ftVGCa1+tciCTEj9BQlIKul2uES82PwQznV0pegj1emPpTdAg1HHcZg2RH3PcGu+
ccfNTsKYYrUTdxeARU5pPfFcY2AFoeth0s29urRlkidteCTdcstyDXOlSfBlwWSP
YbizT3YvOfnKF8CkL/hgvzKm0Vl4L4chrCAGjWed0pEPNzXbRPxmp+mrN7s/y6d8
+nCkbkqzWhVeEWDX7hRIjh+thZO9X8uguTMVWF9YQXfTY9Vb8ZIpfmUYDHIb0mxG
b2LWUeoyp5p7TrOZNoYcnjvY62mKR3g3/Qe/89M5Pc8DkxGwSb8zatmgsH58KCG5
hnY6yo3nHK4lIyNpkTiX6fezeYV2Cqk5iztXALwXeb+LiiFd5FvMpDo+9si4Hmdo
wlNZrTCb1rtY8D23Jv1Ac//3y7dmo7sv4hW5MuY7I+kJg4BDlSlRD6jsewTJuNsv
Db7uiCza8RpCC2yOur+aFmZfOIG4wWk4EHolydCUUYO4ApyUPIVTJN4ekO6/MXL7
0AQsgOGEsudUy1TDy/2F2atbp2SdVX08QUEPPCsGfcV4qBoP5SrehlxudKurS1OI
ap1mjuraj2zJKO8XGM22+Qd+1lyaJG8lZ0kDbJPzBSotOaHjMtX5uJak/ICcZjdn
hS1WCUFWdRFNxyzALWGwnG/8R0P5v7TPaQTpAhLReMLnHF9jiTo25HJZNIW5t6+E
J2fOGoP8Y2xnbBVzK3HjaJ7IRma8y4e3lACXx78tPRvL0Tx5NyYqwb5Om23I93Di
YX75eX241GlQy6EEiNMS6eA8Xjy+jbEG/2ylbKQmHTNj1pakkpa+qRKfo+xfmzHJ
D2NhKHa96fLz9+iMeSoeD9GdMadrynJEOR9+GebGzKA6aksOemmpRmSV3gYCv/fo
YSfAzAmScy5fKhI8peNZnL9Z1+lZ9TaboaI2L7gHrGKpD2Jm+JI9bprUBQRR4Eq2
JTzuSGXmVzabDayU9FzJ1Rl3vMnGt5tHbb2Nx7j7XqVu7COnXJCpBsrF9l0C9q3J
y8qWfG13g1he0SI5LS9wXAwrYkG/jb5xQOX0rgRZKbCffGuXPHAwB3smAtdtrFg8
hsSXxN4tO26Zv/6axZxCY36uycl0TnpRQqvK9dPU9FNAMuQu/u36YMkK9tUZR0M1
+aWz9yn4BBJUxDZiVrekycnXO2tU1PRaGu8J1YM0aXhg+GSqeHIlizAEhNYR70fW
62VU3WrL9l8murf2Kf5Ep1VrEhKsMh3Sor5mQlP/jotsb0yshqzjiPZ+61YV7uGq
MZNSgjVIYg83OWD9NR52GfnTc23UCTR5XoAKNPdz8ah4qa90Lr4ruwulfI5CqqYB
CAux3wXo5IoRFJmIgw/P2rIYMjr3XTjg4OZMwssDIYbOyhlaN1WHFk0CzDp0IVer
YLxj51yZHtUvLxOnT1pbK/EG2DBmfO+KsQIJyhgAQQ19xNkUJbGK/vhPfiuipPWZ
ZDosVqr96zPRF1sHULLzoD5UO3J9K/XLoLaqCX9ZMvOqmb2yXsLrVafd83xFPJ3o
yNyeJzu6Kl26yRvBclOJ3BKxXEpBj7Y9N+OZXpfPRuANUKQAplxp25cAHv3HasEn
/7WYyDvfq4J3WUOLwlFBhL2WPqo4JK6al9MafFpF93B12fYDdrrViYxjkMd4rgN1
i6/K7G7iS/t+S7RKyt+7LexXP+ALBI6VxhIHWZwks0oVdcydf/6K6Iv5Ao6q10H2
th5CESPZf2+H9BZCjRcuxLpo1GaAcOF1Ilvl7Ze/idqOYJVeNkGDnUeeJUQnJCd3
q49Ulup03Ju0ar1vE6+CszKGJ1g1WxKO7muHR5MZld7EwqB2XegRSaJZBNKLjJy1
biwNmjw0Ci3oh8AZyvJNIzTPXzEaE7poAvTvWOgzRgM7XzYPKO5FDWdPUYWir/t4
/elFiyg9qQuVIa1pSVsHs8y5pnvZ9pH3RDrG2RtwUoH7uQlkKExldBpp65PyTejW
Pyi+bV2Ydj9HVQ5nxQdr+EI1+U7zvfFSheoONAYWne33AtD4h5S4tZ6ScxgH6eme
vefFiJSD1/5kLAVp5WLsLoJJRS4HKYE7pKR+7DxQFXcwCgtOg8MPNxatwuGQfzjP
yOXXCB7wscirkwgMTiNNsUGTf6lCnyd/+/ThWmEMLb421wjGKYlna+R2SOLBW1+V
YdI7jFCOtydh5I4XM9uKK6rM4wDukhgwBBLFToNyofArvGodI2+irjzs3oygaukb
jB9YmU4/80R/tXO83BiudWL3znyjMXFbP14SzJS6oygjnsjw6jbTVW7rjnHztt9Y
RbMBf7O+zWsbuWI5PBViqz2AGjQEVFVO1/uscnwFsu7uILa9YMx7kWLas4+I41i9
XhkBmuACTyDUmfx0ZZkpeSHwjF3St97EwD8N2rDNJcgC87hm463ttNOZMP4lhsEZ
IDkUD53PiMY7qTfZNLDeH4KsknwhcWmXAaJMo5jw2R9UPUiDwEEqFnsHOiirXGoN
WOP40XtoKLvwUqJtZke2/idZs6chGr9GaE/JXKnA00zOAl/25ZI9nfBPDhydzFmn
vuAwceHa+mMUhOOFueNBf3uPbjGcNKTnHeouqolAPgVnyIXf4yrDhgfmwxNDqHP4
LDMY1SI1OnQ6vk1NBJS/JjBBC4OHYEMEYvKs41RwcnTgwb4MIR+mHXb6Z6M3UhVA
9pjaqQpM+L9ig4fngPV8ni+fIudNhCxZL2YMtL+Ap2wZ4SFuTV3nMJ3U0IaPnTcq
5qFV5c+JtSbAZlRPekQw6JYYFEBkj4VqSLH5frCfLrBdUtWwmWSASoVvoKCVYFtB
8BpHzSJzz/jJSLtvTG5QafkiiEg0+6/QCN834VJNy/AOj3LoNAxEDLGqiQFZlpCL
WyzxedhJFGsvwAipSRjSIsgJkzyc8OKX3PznJXS+rEHltbHszhncdDWzcvP2xccZ
6ps8M6sNhprLmMoR8jfEuKjRo047QF5YS5QC4/PUfyl6Se1+twuy+binQ8XqzCMj
WQpaqQScMfP7rBpVvUtKmvvNcEKZUHFNZnf1Q2wbxL/TXfTnBQ3nMjdk7McF5TIn
fN2ll+VEwbsdScIn9Xy7FpsSZhLdYOIcDjxx3e++sRNPKIlV5BXmE+lO11BHoghu
wT6UXcZciw0+8+DkOqcu5wpOoVix2wq80AMivNur05bK4T5bsybkeXs5+v8BUv5m
yPUxnw5Gvvr1WGsz0Yy3iLxPFnWcIxkpj7gg6y04JdttJKYeI5JOry41jufYqNwn
8eCRzxgjrzTrpTuiJ//87av3S4aKWquG4Z6paU8+7arAg1ABYJt+UHZynhTPCWmV
QSPQQWpy0A/S0006lewH/P9Bnge85kRtC9AgzBBxNa1RPVLiOvOQbajI6JSdFsUv
jbG8Yieo5Ne1OoFN6bbOpxbBM0OpgoKuf8upYS3JdwlyaErztlx0x3HsAk4az18U
6D46xJix0nJGBlBjycPJ5EQIZ+uv5wS8zKjY/sSp6zbx6dpGavL6DbxvTd96XAZ1
xZVF+QQ1Se0ovoKseZplqb6UJPhv5iD3z1u9IrXpHxtK2+LFi2evJEa3vqqqV1Nw
CoIwwtEMrAUiOzJ358yLwX+jcHGzqu2c0k/emvSdfQinNjQ+nYQ6Qz1ybU5YjYqF
m2aD/vffko5DaJ202hPz9KLhKvP0ZLJOsnHM6sVUMOagP/U5fT0UlqzYqzrlQ0zR
ksPawib9KX42WZ2l8ntRbLDkC5ahBYr+nUX5EIlg+X8G1/odL38vXPUh/IZomn3X
V2t5llgzx1VeCRctgrJ+e/zuVnKJqizayUFk8BZ9tDz0gE9UI0OY5XP1VESFKilY
D4DMKi5SlMdUw0GzwB+9rF8UAFqNSWDPWPp04RAaTtM4nQ0YC3Nhr7p7fSegS67o
MlS3JbwpM9WSW7Af0SQ6t/aqYGqYc5VJzZpf988hmaOov0Qic1tIksKDXwz6Yvmj
IzTwn3AeYBemfp+X+kcew9b+0FbnOkreIK60yDKJwMYJ5F0DPzQCcqwsgONu9faF
KJnQ1lYvbYoj9Tnhj/Bk6+uANKLcP/t/L41Z9pXwLB9xKULb9LnZPAAIy/QjKsiF
u6VBTBQ7IosNUgnEzJAFq6eZTNiYQwurM/pzbBt9gC8WSk3VJ9IwTY/ZVpyrXHmD
dnktlUqtEkvDpjN5kocaQP4QMjMcK8yKZx6we7plHMH6l2tanffXM/2Ro5DGMrSt
0i0zV6DLbx5mu2nmbOOU2CRMJKyvwzpxZh0R9LXNCypKgEpSgBnES+tQCy5Aw4D4
RSRWpq0DljChR3lS0elvTqh/3wqIL6pN9e+nKvgd1pHHQZWljxpFP6TR5HdtgPBI
FnPTMd8I4nJP4UDRi2m9rVtDZVGYI93x36EZr1MUIpCbpcYWl2TI5mD5/uaVNOIx
1pjzrvYJp+IYm4D/g6icw8sM+66PngYFdW7ClgFY4baqESfYfRnI4Kq9KhfkZiUd
Bmx54PhmU3UAneAxD/r6BGXmM01zmZoxoE8F1eFwqHtWlylREk2P7lYDqpkjOwtK
BDMbFHqP4G0+k5E1l/6bzOxXWil6HqXcbghwaKG2vLzw4bUlttg8aObw0s7FnXpR
iKXpqR0LXQPGrGMdtFZYemBNwl9nffjS7CeUzHmzJeCCqDQb3Wmmktxu9oukIEIa
OmnY3HnxpQmqAesUTJNLBaHlpsthrVkw8Q4bdTtdftGDpLCHX7HdbbVJBcJi/W5u
pIQtXKy3DJpuQwhmdfJgJNFORyB5qjWjqpjakLk2Q+RsEXJ+IEbtACVdlTBX6DVG
mhoupBoovLFt5D1oQCC8sRLcjfhsQs+g7VkZ61WmJTSig1ATjtkGSrPbB8um6GQe
yZVakj9Fy/kP05YMK5nDRqs9hprvcPQHHrKGUSR34uA0KWDk0DriEA17undDFkmI
TxFm72GG56iHslcCcoIZu69wVPgZSS/aF7Cn6YNxi8nz+YSM3aTewRQz7rplCQFz
CCUm5p/K+LKlToqvnwsAzphO0nggR6vMjQ/3mp4hZfPVVxekaj2z+BtqkKiZLrJo
AB5sjByWHrmjbRXENgLuiaICEPDEDzIKNtrEeTeeAvpyd7AHoE293WW89zYR4jsk
UK+iqHGcmOMj01IVn6kVheyswgRCBV/3pTiPorv6oXNcwySX3c6Jdp8rBWeCEPWk
PRcZAjY8FFuzD3ZfEES5p2i1+/hwCTh3dK3+QpyJbVowCrjkohkdcld2g4qaLwo2
PEdjz6Hz3bzGR4Taz98kz/zsWePrFjSAD5qd7osnrm72rV8VWoxeIsj22vczeyHt
825I6uqxyLGcoA/tkXnG9Zh3UrKH/KUo6VVnJuZ5DEeDo3zj6WMjQSN1F5DLO2PF
MeYaMPWJqKbUiS9kPZ9xiKXImVEUJccHpBeOZTGAI/tqaK57+nr9smYG63O7tHew
hFvUkOvRO5xLEqIae3GY/bWuXwWuUP0yZdPPNz9csJY+RTjOhdDT+34+69jMFWew
YbB2QTLePo9z119bDPtFIm9C3Hm3tHDf/gsXit7GokYTHf46NPEx48b9l+AFwGQS
IDqpBAHrovUAVf5Mj/SviDZ4sZICQbqlF1NcvyxsswC+6Xqqna0g/ucU8F4sUmKg
d7WyPrCKja9zdWhUdqlNLVg29A+iGlmHzS6knn5hp/6uxnw/6XWz7kvJDmlUix+Z
fan+l7yXMgFzTLufF/x4i6eKb2n7XKpsj+6uxhvQOJ6FMbn2qilqy8f1FhOxoQaO
3T9aDKhr++s4DA9QJkep0tHGNmh/kaY2FRIALF4tSBuHFboZJV73nBEYneaIJ8we
tOuF24A77eXzo4xA1zSsJdLbpJPivzVQl29/Oq99ulC691JfgdNVxxK+LILM/tTo
Crm0NK/gcUPRQLvnzZBCPJxJxmFHquo5ZEcaPct+ZJQJzKh+p2YegzimwJfeumWb
um6oU8cczjY04NPzXG6PB1ybRYbLrkAUbJdkSqwGkliJq5be4EdTt5v+yAyLmsNh
fexBERkeLs/ZtKIf+LYj418AFHBGHW0u7qZXGStFHeF/PCJNVnWxc/ZbGFOtLkCI
0HdfwKYD2n0wACLYlS3jagpC4/vri7pNbOJ0V0rkkR30Xh7RbbFSmQ+IPTWipzXF
SmIoeiQi7nhzZyN78H0dkvi80+khOHN2w9liE3gtnbDchJ0yqhIu4wcvaCWaSN/V
dEs7zduqMbr0F5pS4sg5z/Hy4nLMXdklHmVRso+qA5O9HbzJvNcB/RcQcBoKlb0Y
Jhvw+YfMXxTUzwMqrg+cklT79Bo+pNE0hFRSirz/9uZ77K/w7oXl9n+7hV/Y2Luv
b+b5IOOW0hl6OeCr6nL79FvFfm0Knz+n2JFnUTzFn6hhixNp44VTv5oXlqMgilS1
eaamYn2GVW9Mqnbs+loDcqxyypk4jfmh3Ik739TCQkYHYjy8RC+tm3Pxis2ZhvBk
62LjfprdUpO+s+2naqCskREHzKCSkngitn50TUROF49yQ28hJjdyY+CL5HzsGP2e
TTxdt0KIC29hrhMtGfx9G4MMkoslyb46o/wJtzCrNhKPkss5yM7tWqNOLV+E5iAJ
b2APv8gmedtv/Bi6SsdvVx2YFg7Ctorq0ZLAd8O2IZYPDKZLbFEPHvjcKgGwrJzC
n73JhmBPFOF7fe40l4MC7RERhgVytVx3Nipuf0An+D8KxdOwR70vaF6UkQP9YtiR
9MEr+y/S8R3dZsipaHbntCrEVn7uv2TJQulQH92lqzvwbK0ZXIubOSGfpHWGMXLo
voSx+TnG6QEcs8zGNMGrIwqwvUp00pxue0c7rAbzezLZw0a2I0U0PcaUI3tPx+R2
bqr1c6YeWhS/lt0Ob1UiwP1LHpTzhndwaaK/G/ltVpTNK11FrMOoL60V5yVfoxZt
9qVNPO6GvidEi4YkFScb1kzQy8SKkIEZkdfmV9QCriBNvBfrgVULhlGmm1gLJTDv
ds6P8ocpAIe7DBDolID/2gKdlixsHLREYcf+ndFUPqSawjEKPsqMJzOXDaSWngJE
wHYNzPEtkqoVXjv5X2fPzML9i1A2kL1ku2IbA8j2+XtuOofh3eKwowdqkX6VJkTP
YpFZdJBqPLYnd7LCOWArR0XMyz+C0eANuFbewIuT3BuqIxcjfrmV15s66x7kD2Ei
43XKeEaSdMGWAVgQWbzSHO+DwFAubkptjbTWeqrah5CFoTSDkf/0o9Kfkl/OvEds
/6CNr3LnWFroN39I5TnZ6QTqsBsTnJR0t411y53BAGpfAmxL0fI+1QgdGQGm32h0
117T1vu5BlP/qKGCDX67vAEvH6s91Rbvv4OGkWraR2+JDoyIGOKFd8UVLihOv/sn
beVnXXtLDvaATD/h5we7s2UN/5KMhPtEHAlmiwuhJMRoTKsz20rP6gVx4voWhVCJ
dZzXv2hIi1OsEVlsnrOisKmqe+GMMCmHMgsyDx749g6EDkcsW23BC9q+cJ6AK5LV
w7/2wptmXXRxByUd4zwoScvJctwpMfFWlcf8U8ynnGkVzjNbrKaqXT4SeNTEi0aM
s8jr0pn/hs+l4sgDCsxZk8eYlQfgWSaOfqLV6SCMrvu5I7UZyXEXqXNdcSknvbym
BssR56GVlg3ynE/MPDxIsHbdNpauLIRLkiusW9y7xZneR7+gGsIsPCdIAQGPHgpY
IWiywBvhBpBMRVALZuoq44b2tM+7LwDuEG6eIwCt8KGU8sZ/1elTmW//SULZTD5a
LaYj8mlicNJdSw2GgyBRtkm3KuJojgaqqF5tuW6VJL95yVOKgfS4KWzdiCzJs+bP
mgU5glZhnL/Aqf3yJOwY6QI5yCBxcgjPxAfPdJiQK2Q+WxSFf5K4DpS7ws8ClKrs
tFPgIca6LPkSLYHFj83QpMhqQFVNSEc62n+/ctTXnMIch23EH9ITOSL43dRhHd8A
DcNK24tDv4uj1YwINNQjLWfCcNyTG+4p42uXmDtTIagD5xQW0oS9JfeG8y3s9v9w
U5+Gy0VAP1LNYFo1mSmoslVBD2H+hWqDHnO/70h/aCrA6MVC7ScJvZF2Y35ktYro
tWvNtx/zm3vDfm5ouCoBIryLfjWGN1RdXLQOC/GUZi5Eq9hLZijuVhsAksGvoXgl
EhMYsdkBNFwyhFhrlyDDiGw1llhi/7S95xmi2dB6zQMaFcNqJV+7BDR2btdAJSzf
OGYXkJJ3wq2gtbdtTqSKzxUZPKvE8bpVGp5fcqt9ldWUgPvG0scMPXai3g5zmt1Z
C1eZ5RTXbJhEtzpLypx8HW6BDxqhpl52JRTmJZifSZ0VHto200kI9miyFwyRwY8T
MwBurdWAjikeiO0l7fR1kBbRuZKvkLNkrTN2m5EMclhryCuU+ycHt3Li3D0q5UNL
LuHxVe6gf8gAi9Y3rmQWj0AroZIf5kzA5RwVVQz90R4fhvetiOwN3LhPcnLu6+nx
O0pbCPtx83vlbWU/7Q5bsPQwYkL/QSAQsEcNX80qc6dbsXf2GhFIy1V5axN5erO1
Ww5+RUqFE7mh68IQuq2xCmsdBA6WLYqxs76segXL5VZhi2pthNduvM4s45S9QKKR
r5EcBsvzhbIKwQii3OpjDZXj21bEoo+eaGzhBQ5TEjHfZTywLuDl1fwrq94M0pBw
wx1PxX7A8mtlPYp9+I1T3XW9//veFwyzyBSeoqW23nu9GYjcGTCbzsY+QQ1oJfjW
Pcaqk/dyN+X8NbR7cTbXLzIxnSkZigPEvdTIUugInYsKL6e9C4o6qo2m5ihS6pDb
TKKuP/fR0BTCJMy7kYcfC+liY89009gd0ZvIshA0NmIyH/Cx3YNazqhnYRfV628U
bOrR98pQl4bFXvi6NcypsoXrd+rPcCCqacIJMVAfBtiivxoBX/NW72uw2D0MOBYN
e2FpJEI5F4dWqFgNFfdvABjycOLj0olANarhVL+0U736lhX/o+QkF2vH+q8lPxkZ
BcpJRvJw9C4uQ6G/aB8Hcxa1AWnbH1K65aF/feV5J6Lh2zYtohbnqvUPGyTkMFIj
2oFivFt1+6ocEQA2zbLcuYiaIDrnVIf3glZ1Lg+l6wc7StztXBIhvrI5oQu/G63x
W1iKlF9shqCColm+HFmbRDiAG8j9ySgEOjS0nbi4FNv6FotlNY+4t+Hp+4IiZbGO
50JuDQy47qbuavJYWZa7599D9jz7qDY8OQj9AoMLY3OALHsUJVmqiTCpWsdtdnCN
a1ApzYj5FvlXSeBdvqGyUAUItHrRU0CxmksDqSTUYNaBO23QzzkN2awnm573SrA4
yjo/B+Q3AsAA1+hvKnqm7djjjRFauPbE4mlE0iT+bgLW8RQtjvBBFym/VGDLoRFH
/QjyinZT81o02DklgMWZnxNhvnEcqdr92sa4t/7adHp/nTR66we/anU/Sps1Cu/q
9szWH+V1mp2fAqa1TDx2NiTV7VM6R0eaCS60m+Sl28W07rv3NaNL31V7V2hYD5Hi
tK863NLyzWNCG+/7Rh9Eoz/wYvi8dQUGsi68MOHrnZdcZdQ1VohzSdsJrsxesQKh
p8hCuQp9DBUGNN+GJ3gjtgiVMN/JrHLZ4D/AlZgRt2GeXshzPk1HGM2snZHr13T5
TwrESG8t2gQ2xsAu0NRsQKF9g1CAV2kND4wqRRIJAsc2LZcKgoct+EfJyyu7GUvC
bdCHlT4aOfJ8BV39R6WGN62RkwWTti1FegM7G7ASdzkiWgGl8GR8yfsqRTRgjBfn
Irg480jZ19cnS8s4SKfVwLevbod8P8AV+d6Ra1YVlBLdQvw+YWvcJYTj+HYJKEdf
CaT01t9NYTIDckDedKOGOTTqpmKxuMjSyuDQEBc27bKq3zjGG3VNdwVTfVFpZ5/6
VssHPGR2qzmmlHiHDL5pb0BWyHm6a6HEkJ3HRyaHE7Rqdi6IORGopK6yCvjAytrd
uwyvzVgonvRBq2ms/gzNZtBWOREy3oTPZ2Ypy5bNHv8QoPslkByWQrV+Pk8ijsNK
jc/MockSdRHtAAytl+Q17UUYsQgJuVQUcP+spWm4/boKdQmJXjst2qEK+l4Cj5ay
FAI8GDCjBgzaBzl63dbjC8RZzH7joW4q+s7Ns0ljFheotRw6xsg4PjbdwYUzzsK+
U994Tcka0xkrscr4M23kJLE+wwpzIyRokzMw4n3WPuvrhxRU7CmaYPpTbLTtCDea
fdgNFg70sxhIQDhiA562VM2RTKIB6SXyvp710vXj6YopV0fM0DjUmROvoHJsulEZ
5fc/D6rncdcTBDbgngYRgwyjcyXOPZbTDp04yY5gQRsDTAXqUhi6AiFIUrH0wZ0I
7+tcu6MtZhEe5TKlz6lCAHhPV0aVHmTMGNwX2llSpFUK3Wlf03kwCAQ45S+0+tHc
fhH5YFV6jy+TWPRnt0d/yXEyKFmso94ZT7YzXgoHX0gMHzqz6nrK5LFpAdzafGmm
MlFjw/YkXRkCZ31/2+KOYSmklNjwxT3sogkZzSvf+sfoh+WBxxIDffEI/zwooewn
kYe4FAFAlvsivnBLQMJ3P3j2AHSoWMEBsrH7KbSrhKf8buX2HzX4ROLVtXjS5dHq
3jnRdfXgsXA9sBLwH7pjrSLDM7NZIpVDiNiDvpc7voyeC4gQAdoKWpQ1nKCgKztv
nOKok4YJ8EgcPKKZayfPfn6plO6TlomPLvvlDAR98sdJQgrmvQZG2IviwCjIKWUn
1zF8o1jr6QG6FExWcCaA6wwa0W8zRgvLZvxM1OQehnbBQooSeTxVuZf4hDbC67Ha
UsuaYlLlFT3UR3NDtxQOgPLNQCTSbjGFMRuKBLHiBAu9CE3qxDqE5pk87psWBfU5
JVBe51MtHbKVT2mOcYg72WUEIGNHWwTQIOxoDzx5pVL9Pri+KUA9yKP+Ffgf7vCI
/rEjpdi3bbMZLFXqB4MZU8/svI5Y5R6DN0yar10zP5HzX/YozHyzBBe8uXQVkgPG
MHwW5xmt+XVhS6tBXBKCYEnmYDpcrQQcLW7pWLGORJi+tGueb6ItvTbtEU6Rm1IG
jzAEccULjqEG3b+xX/sCnyVfOmw93p6sNg2HaSV3b3mTz6oJRFO7lgegPeAY/MTr
8F4OTRoU1nXzBJ2McSMfs+dMwJxXS9y+Xcr47BQ1qTDLwmOoYMqYJXoeHLizXaom
CJbpqOrhPBbrT1qG3uhTexdjbvjlW+LTW7IxUhL0qruXmBr54DFBVSRiuvXF0wBH
zhpqXnhQCdHV//anNd3i7JIAA2200tlYY+c3rPE0AMUJorb/f9EhjhqvDu/ywRL1
X/XaKCuA5Ut0fFnf7nOWT38QZ4pQMzU92P0EU2rQbuOrwdL9xd+zqcymiZ+T4UxJ
P0xXMXcYjYjfKFJTyMOY+0LscY7f+v8N54xxaahXrweZlXrOXlsbATjC/mGOMr7S
noHBBVELCAqiqOCG3+TauhlYFrx+rDgL//UIa8R856ZfKoomeHUeJMG3Y7wOb+hD
uUmN5d7XYl3ccflIUJtuLvCsvduK7TAjQ7vMunvFPpMDSoycvqXqU+WhKJuRHHZV
H9RO+fw4oX1AUCJLE5BZTAyojP9u438fwWbge8MhyuogUX8dSUbjNdLGTNSaYyZc
nfgMg/545oy27ckR0Jx18uF6DX4blGg9h7KEi3L0mLwuzdoxzHm3YUQp8+HYyTNg
T7M8anYVLpz1licUgVV3QdV3HklUPpnBeb1tTSGEi2oK6CRLGBgy539DaX6rStct
gLmCGJCEtOg2k3eOfm+zXzgj2aDifTkrzxoPozXzMMwjuFSeTRqmHio+UnxgmeSW
xa/GiI+VyS5JR17eIBt2v8XQxgltVvPLMNTIA2tPFj5/EaNo3ZoD1K1SzafCSu91
nDAFImdXQotHSwcgy2Dta4fRvqpgYnE9XwP3ZWZnKt9Zxmq8EB93Ug/R7NUvvAmm
neENA0BhT5qlp0iL6BhGVab1n0v4+FI4w540in884D17tttUfCu4iX1q3cVKd6KK
/LEI+v/FWeZXGx7qG+ufTTpxbUjgpMTLACiyPgp26f8jn8JaQK6ihj1lZlfNnhEe
N9TQ5du3tfQfXrmME5StBHucFf6CrR03naG7+LU9rH/hN1ajCltxgOfSLoeX8Z+I
9+k42ZbsspOFDxs+KE/wKfV1TjW678GX4dhu/g+CVWGL2zxegDl3QF1hQfBl37sE
tnw6NWsxUP5pmcps1HVPl1iFMzEEjaClg0oZk9XDYAfMKDuLHMl8jkuVUDQoTGaH
Huc/L9EAn9FA8fQbO8qYLXMJF1sHHOUxiHmodw8pKXoxMvNMDYXMHeyMGXh3X3xw
gsv2F9iIqbEmvfhM6BH4rnA5Ia4QlKPURdqpSOy3HfDRfg/vUL8VDF2Ick0hRi88
ZyOfBdjeEt0oS77DrDh578Ln6cxUmvT/6xtIRx0WoX/sstyG5ceVmPQQ7+75yflw
TORmkTIS/qfWOpEl63l1udGC7/NrmcRnmG3zFemWH15I7NGXZDk3khTBGm7a7PyQ
SRWkrG6+yObuaSx1EhUaBlLXEJl5IieQyqPmh9CDHcRzkiS8XZKkLnnZs/QY4M1R
15I4PJWi9BQy+AJS7mqhpXnQWyaAfLllcbG8QlQbCounkYmESmrnHpG/8j2yUTwU
HnAZt/awsfFeOf2Sfhkzj25ipXmsq7TuQOjEFGJPBEChNWhnSG91fXKwNPa21j9q
T3WzdnexgON1lCq3hfVpW2Uee2krrV8tqJXp93jzzR3WxSVgEuo+YPmoAzIrkw8n
QfAiugr/sB46yNsmZmiyure4AUBxf4QREQLTOPOQO4Di6VHi+j5zln+VFGvX77aG
TIt//6TEqsQkvwr59tZTK1wqMChhG9aM+ISuq7/waJ0uoPYztTxjEUV0nubg/Jvm
keLVtwDwGv7jOcItBhbN2ugnGj3NcetjuKtND1ApFDLNfTrhqHdgIpsfoOXYBtLh
ziv0PgLjCchpdyQIk0MTBf7xikqsYuwUHy+L5++1PYx3S+1mSchHwLDIqio7JmB/
K2GlXQDw3Jt/Zu1IZpvJv5YUS021ZO6YjRhLLQJ3EvJMhwe7y0Zdd9gtCAnv+6XA
jMi3NIfcER+lJLs8HW1OcWdDI2/sYp+ALuY3rcFDS/cACkP1OLjYwOAHykwGifF3
2aAlUVjJWnW09horo0KW3dNeg7tvVU13NoDXNdhWzJ4uUzsklmZOe3uvG01JtyQI
nB+YrpiI4nvheun4AdnJNL+G8+NlWsruUWH/9yZSOgHwGkJ6XTuIxygM60UP1rZP
OkfY5uMapyQ4ExsS0JbaPYjAJLD1q+WfKx9V1RtSoBC3gnym0YyRTLWfFZq9ttP4
RepOeZnBpygBJx5xcPlou18mLKpgXzyeRCKA9r3T0SPYW3d2lemKqAFKBmpwA/TF
5htsU5lPeAQTTrAe5OqjRcBMizVfLiYdQCwwvt3TFwu7BLFQnZ09mSy1iQA76y7F
AaQl5Eoo9iFnSdDXk4+srvTa1KvxCNSRy4ybLR3T4GF5OxgGdasYRz5mmTA8MENG
rFGPmbO02I6HEbOwxuNo9ZifGKwIo7mABbPMynO82m/7QEDpAFvtMvO0bqEaZ53h
+EpsWQs/EGbcNaNt3ELksLV465vy68EAin8bL0eKk/vle9+VkR7uG7ISV8iXHMCo
y6I4XBEDXxjHuFsy5TUGxUBwqCZNKZDJU0gh1jCLOW38f4UgHJVIvRlPLaLZZmo1
K+anzxHBnjrrt4/+KKPAVhGQrkLzmu4dhG49L9wU4hRTOEQC2quq8K+nLtyncZ7j
6M/gljsXUXjKyvQjv9LOqOYgKJLKnIh4vE1vB2jumRVBBqLJMrfp19F9vUG8QNww
n8Eb7Z5peRffhVwLq34CwrGMETUUoYnPPspvIFwLlV0+CIDK4hXdVpX0J614wFWA
5hi/SCzks6tc97+ayVRukVbVFrzQNEAkBRl1y+JkelBaD2trh+yVEww4spiAWWd8
ag1O0X82huUwGmsjhTnTjqFH+2ANlssGelNer38msZ1gb3Vn8nyNRKbAa9ldxzAy
a1f/1OvOOTfOzEMM8LZ0Ujp6KfySbI814e11i/EqCw/Ckipn2CoFIo1LRHAo/5XY
jT2pOdtzZRiijKX4qkxtOzZ3H6orXZ5jmX4Dc7pNx4t2K/5fpe7PfMK3cwtjzp4k
fv4930QO11u2oZ7hN/q/2z9+2Qw2dIuiMToM+ome6Rr+Xm+0xU0uoEQhPM465Z5Y
mx/cZWrOeEurhum/UEHzvMVXMA4lqPmZxepUadw0q9GuduQNZIAkEH6vpfSwVSKd
1lo3QmasNi7xBgggOKMd4Byih3ftlAWVxXlHceddfFrC+0tnDZBMwZG4z1p6mhZF
SqDAEU7TjW0+2r9+Eqvq/GwJLOHp48/zQ8pA5RQVo01+YI1o1aPuIiwOvWANNgkl
niQrLcPiZDYXkaG6QKiSp2t4k+I8ifXlpnWs9rDGH9yGItGzyyCnCKkACvoz3Iu7
yT2tzeP/CW7jg2djasSzZM6MuCJ1tJ1SURbSxpL56GKiVHLuV9OGNy+yzDJIN9O5
UGZQE06sdwSHL8i7nSjR4jnGVwLZ+3pTgHQcAGpnboYLqgh33k9GT2zrTIgsvo0G
VgINGOgeciLAUW86C2S11fFD+fR/KWHfcbj+IwEPOEZ6dH70TnHATIVxwvr6tVU9
63eDXITWwGAs6TZ7ks+hrQGSDLXdEAWc2iiXyHnvIuEezbtY2liU1u/NyhFohkvV
NuJX34frY00u+0aeY67aYp2szzdUU3ZnkeqgiC5nhcaPKuVLmLNL5/gYylJKOlFo
zmFMAzS9jwivUmnFOm+WbApcTggy3tK+PLqDeua6V583qmKxrR6qCjh+aMxmm5Tg
AdJM8aXmK5trK86yTDUJ0rvoq57sLvzUAdz6vCFubfIH/RUu91h4LQendoeYSS8/
SXjVF8v026YX73zPkybUx7F0Y+jEcFtPzZRXubK0OsxzpLx0kkF7RdumEXtwhi99
t+TZYHhF3IkaT4IaoA8V8bbUDwrRNFu6W6HOP/lYKDuLU0fIQo7NGdQy5MhunLZG
3VLwCDgkKg+fSnqEZlFC97kLjyWZICFYD9+ORxJx8HOuJxNTz51gwa/4H/Ld68iT
ALVuJefJjifxK3UGIz/UAUAwceEF/g+g786jtOQJF/yLIeUk4jQCwm7SyAzXlB7g
AjLlSO2yVdZRo1xixvd8WoDlEtTXdHkvZBzqlJMAThRthzQElCw57VrlZGike7Y8
4JpmnlRMhfx5qh+pCf47srAISCGEUUAW4OQWqRMAMQQDp9U8u71bB5RO5T6JWYBD
Av/o+Q5755uKKp4KrOAHqnl0tp4H99xCMlvg5l66kswBjKTWFgFXZfFi+eLmwnlS
Abe/4G6sn5qbM93PX4QLzAxyOqlJvMr3i0FVglmSjLrnGO3Ege6pmgypQy/XTcbB
/ZKvbefe9zrLg9d6EbJqmvVyJ9fOPD0e/U3e1AMIk5/EnkzoSvp6cJCijG41ewFD
Ug+2yRKtNjcpnlLSK7JQnx6kZx7wgFgZ+u+quA1iqzdsRCADKtnJ7nDIwOF6fkLf
jlr48K34rhIyjQGa4IpxPGHbhKyGIPLdnY/rgBbgz5T8xyQc6SQWzy9v+j6qwbrb
iadwUxogd6NMgxG9GplucMaE3HFXlmJoPuk2dFNY1Ea2Bg5+o+wThvoihUmeUrmm
8Luq/ZlN6HoLu5El2aUyfoLj/jkDUWTJUYxS94rMW+V1mVFejhuj5E3meBjOtoW0
tADRbGPxsrxzkrD0cxbHZGjBbZ4xCKVONMGW9xIarJeiwZIujDlUwokI4JCJMIh7
AS2GN0Sca4/sw59lNU/tOiL4aJGO1Ne5fkMAcFRcdjrt/q5PptCiuhn4s1nmmtgv
8ZaXl6oXdDhdC0J7MzRCf1n94fZ9EkXefYIlqO5fi9s6xPdulI5TgawbZCII0I9O
l/57eAUN6bGhtmhVhJ19/jCO9YbREmpxAZkDhWE8nEc0jTi6iQrHUIoHJG8h7Abf
6ySlmIfdZ5NeDvU3sQcOhbYaT9WQg3+nCMrZ/DPlZRwX++XP3104uhqixput+lpI
YzHtJd7nPvYGy9RI0jKKiupEprjcuLRBqyLVZ6/b7JPdJb2kWfMpF2AnguMrTI2F
rYTdwOPylAf+rDCGuu4o7gq5i54vqwL1WkDaemiJ3IAIA8KNgNk4JiB4SrzKo7ql
z8TTYtaYtciCcffyeTk4BRA3UZ2Fauq077uvTOmguVJ1d/yEaJSEbDnMpN9Z0WoT
JRS1T3JIwhU9GPjZHtJxfNtPXDBcTUe4E+bmIPG6GqxB8pzrpFEz4tg1fKREUnaG
psHLYouw7pnh3kZouQoeAYX2sacEmGFoHRk//TDF3t6ZY2W58CGXnre7XLYOyWFd
fs0UqNVVI1sb7g2Md4NogM4HV4eNZ/PrXmb8UhDqGZzi6tc399GG1eNgIpjY+VYi
9Pp3EUxsnqIyMTHPFPy/kyuyhQy+9WAOfDzFKB4Q6j9Eo63Klmj9D+ragos0C+9D
e77aIzvVNrweEzXCFY9l8vncoKkeAk07AGRrQNzUZMaxcjW3i4yS0m94MekesBew
b+xk1V8Lzu+bhIEr/JMnvIUrpIUaiiDppCQyDGvBXb7IAa1fwWeJ8JXF357jzEGw
OGXfeQnGiapLkqEgVCfAwiOj5dM52WoO76OEVauNIaiMFL6VCkEs1kG56+6UV/0/
EvyVFi29UDZ7LMyPZywdN7t/XQ21XDCOiNZ8kZ2r+n8USIAF9pgLmAbjn1aUs+Nh
BuPjVGBb7cksPgN9r3GYitnEFkDNQRaFY8kQBgoMKe5M8XQ1gBPcl72RmF6qZ3KX
GjGvBRsJMayOmzDXlbb3Q3AvC7zM+9OGNSbocGQwZwZuaS66p+DbbVn2SFwS5Qcx
YkJnCwie0RCbpHZsJuGKSn0+6l0tzMjjWHZsaOFJdlw3dB0ChQOrHs7Hnxj+w1wi
sJ1ohRQY0T48eqz7fnGyWcx6IWfGtHP8alsQ7/n47TsiN7m3EHm2B8mjFit4+Mmx
phiG5EkaCkPG19TZ80xsGCljV7EeOn4hLBnEba2tH25CCECqpqP4BNsKhRboztGs
imYe9oJFNUE9dxq6zjQxG71hkz+LWJjats4lvBCbrpQZ68i98rS4TfLwDdsdSmDK
p6KbflPqT5tQV16QWkkYxpv36t2cPOXPUMDIkpbqvIUyCgIKeTm7Jr1lu8nQyPGm
PFkKuBeJmNhUbuGx02b5ZodiPS4u2zxmKLYx5MHZbPOB50+wzjmZQlfGhiGO3aLc
Wy66L3DlNPwjW00W93qxcjGqUHgCL0pL6oXZ6lCPFheRbqQuyHecQfdPw1nerezv
riffOzfnKXJkQDPqMOLY9F3N8szypBFVtNy/Kfjn4P+oONuOv8EmsUPStbJurDDP
gRvPcAX61IdIqmPoLLEBdBZ4x4EHTTgiPY23SDkp+F4HL1gMi1Z6gZtX82fc3LIS
q8w7q/OldTPPPsX1OL54MVCPv1xwpMAYOGLy1DlELM0D9XhY7Ps+4AqjqiSSTRsG
kw78rr1BFLfBFTxrnNCesQ+CAFHTJm8aNYe2tKiK7+dQysvxMWM4CNW59A3X8M4x
ruXnCJnLnS5S0zadMHBXzVvgGSmVY5xRw0629j1qZBY9VR4nn3FVzyKD8C10HAN+
d8wBibdFtWlvcfdNNnHhbAaBk6LIkZy5uj35JQqcNibn83gd9qjhdXUZ4W+bPp/H
yOg9Fy/OYJnXo3QMQQc1YdZXw2lCuQri3tod/0dj+XQ59cWezCgy/XbIFkOy3x9p

`pragma protect end_protected
