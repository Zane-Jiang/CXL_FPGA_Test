// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tDgOvacY1/0sCxyFnRK69SF6Szy+GCP4zb5s3R0puS3HXd8LM1N5JL4Y64Go
ncqQn7T0HNMBFjcXMS6ncoHeNZJL3Szd1Uxwxw7gU3gSeoghYqzKK5DVLVZH
u9ci77RrjASmn0xDuj0c9IHf8o4KPgAoplvi+PNaRrbwOlk2wy45fVfD8RoE
pdfjkjQbUb4n5wBBLYr1YiJI8ouT5myjKBLVkLPT6pAkudeF23T+LN4WVR9W
p7h3ElXKAJNaRrhvIhcBaSIBbEuaPD6wR5mCBciCoq38O28YWhKPAWkdogg/
w+sQMKhaJKMUcLNTqqhNbW/9K0m3d2vMqWPtq20gPg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ojhGYDWyYN0vbYBA44mAyvQopj8eL2Du/GZ7kfdP/yx/5YF6lf0RALIRvFrw
m2UTuVtylvpw+g5p2izxRQ27f/zCSPcGXSb3SZv8YgKK1iR5IOYtxaZQA9b+
J3E2Kd0q4qxKHVbYd19PZPPn6qqd6lHfNqxa9DnxV+lWKpmHsurBNP3006UD
Tl5Ttxdja6+md8poBYJPpggljbG+LTaVmZ+6GhOYk5nJLwEXI2BqqCZ89s44
YYPqKoDbWORp48fvYHaGOAu4xAOYTovBjJJVwQ4JlWrS2rKczPY4kWTwOCHs
jn/5VEd5W0s0FzgJ/IPT709frxFAqBGdOMv3l+m6qg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nXZblprU/sJeD1lcXRUVAg0+kLTMzrEqoN9ZsOY2hJnFUOH67dtTqQ+ppB+9
C1oBzOdPeFdUuWeEUyAXu0c+HTRHihoTZ9AAbziYerR4eoSwwUXuUy0WB5x+
LGmv6a8313Td4WlalYOfWF6dItc1CQAbTDiElMC88sMRp39bDO169rbeIt85
i67GGGzALoYCchizwh5GNHqfKGEWf8+kZLrtoA3FhW+9mqFUCUk3Xwk2w4pt
q7sB0M68oNwe3zTaxHvLIbq/iTpLRd775Zla97LPtsBuy5OM53UNRwXKOTL5
haE7T3fwqJy7etow/FDI/V5X2z8AJkebKuuL9M1B4w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ab2POd8+Pv8I4tpIURn1o8A0eJSV9RH3XBKWx2kqrxPlzvHnj0AmIZqAX4N9
ovPMbwORCukKYfaXQUYFYxTbQeTxpLuNK4JzsmnFw7uLf70voz3yv9jr7ylO
skln+XPg2O0H+zwOFMm+/dZx3DMwY1J8CkDlqZHaoopqF2pBjAE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yGv870kLifSWv02HNVR7q8Cyt/uajH3UAkWVCUDjv5dQJJwbHb2fdjoq+JnC
rk/B+9HPqHtOQrUqfTpBZTmUvCNuKTeGAPdsJq61p5YF3+kuCPZhSENVFt/6
mpO7lRv68q5NNf98MRPrl2c7NDDQznIyF5zrphAYFr6UtKYOo/WcT2ivTODW
jXyft8eQge0/29up9zAQiSmzsawDeiv+nemKA9ImHljHQr1Lk3lUlLQfOi9s
dUUcnExFFx7SCHlLS048xLxSCf7jCCe3Qv9ZqWNZ/crUiG+39Gpi8op/spGV
+NlA8s4K9O8098gI1ymAkenPc1H/N4wtS6cqXQs56Bt8zlxU2rvlp8exhEUU
xl0pkjhSqS/cVTDT+tZj47yHn10bzJYbJfvIHbgcD+bSYxtPuq0sTqj9VSTT
deYyMjwv3T07/br77LPjsKk1XBkHiN5sMNwaCtNMCxj/YeEnZlsKiG0py9Ou
m8pJu4nORe4MbeuD5aaeP/X/t7X1dqqp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EH3zRKgHWeUXClha7J16cBcMfyjLP94pa18gfrZmvfXLqRkiQLiaDSdOxqHU
4lhxng76sg+LNzMitiFfGEl+uVKDSGhwLqqG3Yu19flu9YoQevjj7yoQ9+qN
wN52xFr++Kp0CE7Ce2Ppl9aut3odnaP1iz4y5wK/E2JvX3t8WlM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mDDmmvvTf/EXEJXz45TQEvmUx5NWFLkrqYnFrsTrNP9Vku1d8k/o+ZeRc/TU
CSdpf0GDWu4iGDKGNTDvuMGdXK5JoEgyatKOUqj1BHt/w86B2hp2o5Iy5Z0z
NQo4kFXU5QIlDzW3Qwv05y1Pcc+6LYamLv1bKfpGO8wl2zgdsv0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8272)
`pragma protect data_block
+F6VGC6Y8fO2Rjgx+o1dhdxfbO1HyZLO7jUsQZ9EE9jUTS+KYX4QTlv38Wxu
5vocW2rYVN3z27cue9vICAc95KGVSHxBy//7JU7pYiCXlPhZwjyTts1b9q04
glYTjACXNrewS2Z28ecKxpYHUiAzTSQ/3w5tiUIPHq3wOkys5Ho/Gym8A7kp
P3skQUyHXRgVZeVrRMAJFyeMijVK2kKwZVhPiMns9Vu2ovAQ+H1DexZ2dyDO
oKeXPLhhAmBPiBf6Nmg4Hc2lmdt+kR4Dj6gfrmYDaCYIbb/lghkvi0xvayNg
x2mOgT0RY3OTo7lUvUIgwkYa0zWjwFF69dFec6L0x79FRP2lCtR/FT3AGr3e
a0d0zY3JQOaJW0gbFO/7FAYQz/pl6Z2scRG5CU70HQJl0VDhHNcHi1qmjnSr
unh5aBmpjaq0oqVHmuwbnTgNri/Rvt/I/b2D8aDF6SoiszFw9vZbP2msaMtY
BU0pZlWzGx3IB9E6B+uW3bGbQJYNolTbDJ3WoTVIYDft2Va54sKEhl+x9XHq
4d1UsOs7PKRUIxdKhh5uJR5gqNQWguIy9YesuLJnzj5eg0R8h0/KRTffXMh0
cQvr/nGxyRwAU+BaCYr2je4yQPl/igJa1fJW5JQpFcxkeGR6tkV62m9z2uvB
u+yWjFhEHgXV3HG+VkHDp/oEDq6aNrjA5v7g8CTVJa5O7sJxnmBZchnhTC8j
akBBgV7wAYCNab80MvWQb0nnSam+9UE9BulZwLPWPvyXNcqh4ObMsE1ds5eB
G+EFh7UKjyT8Vs2Jq+yrKPMpIv9XONuY71JV2JqlNXFdvbMvgd0jhliuYGbI
BjpkfgcyH1fEy6662uAmS9NOgfUGhsODoKjHZYkw+jGj9lTGDBb0gPG61KSD
4E4W+ybtcTRd25vwaW+gKs1sYucdrH2AtOL1ZVQ5O7dNNj6wFlQukKbqZaXZ
3h1Oyan+JXsyVPYocci8r4jE3IgtLr5AR53n0pUuEein5YU8ZOnEqTAHsOyY
gDW7XuGP2eLWtH44C6SBur6fOa3DxHhvpZOIsjgEepPN5l3qVvF3Gj6jIzbN
fCpZ1U6sJB5t1k7dTB2O5z/TjK0WbvN3HCM58f6x2wevmgE7QujSkHKa81Qh
2NDjdgj726vlsX0YJXcp0m2tKK4i2PKd4Q9GS/HNeEXMLEYtLxBITeG2dOOZ
/1XOCQDqWoWYHOIKG2KFVXqUA6zzyvKhcDf+2iWYZ1tqeMrnF5Rkf3LG2EBp
aQZ5HlrG9Zu06SQAuPdnU2BfByOkI7Y+RKmofI74N+jajcisFB90JN6annlC
ISFr8bYk5iPBWRNgiMf/eN4b9aDe41BqcIOzx5gajJRf6RqeWmkWIf04WEne
fuJTUSTvlynaCGRh5kAxv0rYwdxdxWXbj0xut8uWKSJxoGvH8YuQ4rGfhjhJ
X4aZ6l1sLGHE/UqxPjF8Lb53DvSBc1pgl21aXOyjM5iXIFH9w1lluJpKKQcn
92de6MtHVre1YdATdBAdsP6O4DGNSIt07wqkA5i3jtJteEtP/IelN0MKibsd
qWHGzvADMd5pfMPY9qp6debj5AkuPkPWfyBWDIqGV9uack8Fl7AxfuTUAFdd
80h95yVw1Giyo3yVEYJ+A1XZ4iwfuAAnwAwjSK5TL4Xc/+m/L7e85yUWHw80
BDUfSN4soHROlYQlF46agG2jkIo7StzMFXwtNAnbb3YAE52wLtoFa9paxKIP
CsMzUZPsCKVYHKuo4L4BgRGMAmrwZYw2NjEC/3j9FWppMleczKrBNb2mFILk
Jl0n23aWM1CfjeFTBEAv15Y1TlNXhNUnynTHiU9MDedrGwmA8yg2sUYiICdZ
g2KakQ1K5+eQxVkRSN5FCC5Pty2lbOGnSioH+0Sw1szjJWiQaDUUYju+90tU
4s89sZ+HUg/nMcOhpFoFsX9wr7yBAsi6z5O1/hnGTGkXRNpMRoginzjfG6uU
rLkOFafzjggW8ppVdBghjqxW+oKLiTJ+x75YPWfBTOLvui+jUAiJ1RVF1udh
l+TVZ5ur8BvDzj+cS0ejw4MkH8hFL14Xfem753FFPqxaoLnb445jrnUfaMzN
K9t852+mfVoju7RXd0y0fMmPVF6KM66Zir8Yfxirr2XAUNqEB79hfq6he3E+
mDQrGgzcqhui9OAFHeuqMgyxGMTYrseYNTHdeclM3rNcXo/pX9jwnNbODcZw
1MDd+KRcpFnJpuLHYvbj/FYLIexLAjshQJWEHfNK2hyE32/GiTeHV4WBhVOD
IAbN69hOpWn1gg0+a1mvLLD+IyHcarQ+ggJtjNySpGV3QQPeTaxJss9NGinY
jpNN7qx8mAzJ8wa36BGs8Fe0KUQ8I1pJQAzuBEImBNuLUdVNnB4SPUJtJ/7i
CYqlnftXIBaBoUwkGyfKWv76vnyIxa5JihnqG4UHjKmtkK1yCAOwKz86XZDs
8QwF1X7EohpiScE3PJH2bD39xGD0m5mqhOvjxF1kcV1zWFGElb13Nckwxq4T
N3tQuLOh/PZA3ISKB0bm3zlxqWtG00Pgd+XshhSfoXtNF2Xh+IByz8lrgKbB
vxNBTGqIFfubp+TI64a4DmPeLySxa+FXzzoh359/DDuLNSlyOgUiRHCKFp5k
P/HypKrPzKg4klivwRty9XobPu4mfPPlc2bGuAS4ykdqvqLt1Iq2JM+Uwojf
DLuAJq8tJECx9LbNFNyEvCxCuB1KNAVLy/B4OoW5xXsTGQIeLMJVXJkvyoBp
yMUI5JyG0sWbS0pw2YWPFR4Q3inPgZ6GlvQJyEiElRYC/AfJXBIwJesA/hpl
VtvSsxtl63tWVJJXNsItOA1V+AqpSBeGAk8QJzQ1PdzsMh8PcXz0TSNS6ji7
o5W4bIij3VJi65waxofkkcAT3rlDPDmrJLfpwCBW0DLcQ5o1vMnwtzigFbdX
Xxlb/7qi4DpH72mKaFMjVGqWZhDcLQb/1kFSyPaDjtX6jz1nkS768OwDpPC0
E8xugmN5V8AFr8PxF7xTgOtLSY3DhYtmW+N/kjkjY0AD3El+Jy40qRxf52qE
oXRfxfK0xlqx8ANtGd9VdYZtDTbmhriub719zIUa5NjcTA8LjOhPT9ceo+2g
zUJA746oybrwrqGUV+gzeZzWI3A693Y01COgPY98rmWJ+mH+4hTzgV7l3eOa
nqT5uiQ9F2EB4rxn+w8SCewQrF2P318df/GKGI1M7Wc2GKBmDBb2BYrHqyXM
l2prsmjX0uQ9sJY7IONLbCpdLrhD1IBebnI0WJ2kYnnH0/smhsTf062YwcYo
6f8/JHal3lPAas/ogipkFS4Bo48dQrGyzZBMLowethXGl+iK2ECHpkxQst7Y
Fvpwpwz+Dx7qFmp1DRdc2k0skgy0Z9TiRjQ1Pougzgd2aWQOLsxebTcku2Ko
bSn+viQEaHcCjAC/vsgqTEXTJ/coAOXsbwVocdw6nW6iX2gk9whMNk8cJrD1
xjQk2ZFi+PYJjwLQkoRhFn8+D2olEl6YfcX6G2fIYymdXTwltDr0R5zhg19I
sKBl5Q2wi8TZQN6+syuVSkChjLL6KbYmGL+votZwxbbTPAI9vLz7lF7HORho
TIR5bumWb8CC1N4B/NT48cHAW1WGe+zgmXaf8NJdMgSyZaqyP2U5WZh+Yo9V
0/P8VGERs07PZAW7jBnu6nyHse//EBhiCBCm0t+9iaLKj81Dg4OHlH6mRkjc
oUIRH2BuRi9ulze8eOMl6ry9e5B5QgYs1w6JrEaC1tRC8ODu382frTgfDDQB
S16falOYrnn4+0n5t4K9Bw9r5lL4LXP3emIEPVA2NB0W773ROQQ59ZY2yyEv
j3XOuDuKUgPUZJqfNPqxF4TnWhpbqlGgQQI3hKKuzGIIdmJuOA376OBBwrBO
peTM2+1NQK7lKZFuAqynEBSmEq2otz6o6HyqmB+H10zie627rS9ZhYWTLRNR
OXd3lRyAcD+0D+0j0D+Hfix9IwnBbqBwXDfX+nJkUCByL8GEFZOK3hW4lAJl
vwhu6QsbtCQAeikcpzV2qP8rDl+0NwL0W4yBeefEwtOmj86ANZq3c+JhN+GY
2oOSTbZPiYXanDFVgC5u2HuxvYmNXR3BzHRGFKsTPOIARRUM7EzKLre1zelg
H8UYpdqcPa9bbyUpooUdwng8N5o4QZ0hFxbCSn2+Yw+Z8oTWVN27d0ImVO1M
TK76Mcfxex1QTGG6htkKj2LIy9MBHJKxnn8oBlDuEfQCDtYhMIIdI026ETtb
L3JmQfpUIwEX/RnzWc94yYiN4wtTLu87hA0oL5Yf8FKSuGtmqdNd3fsvdaj/
jjFAUNyeCBePNqOeFnSGHOVTByK1w4Btl3LukPcckp3oQhU1qK1+6B37GVEu
KwbA1SXigxeqcuepmSR7UQXTpEwKyB8TA52Qtjfc4wZKLsTGuVrs1cozvqW3
79kCBgQuLyKhdVq7OwbKdJgZYQ8+6EScYTAA9e79pn05Wc3YFF79wBLQR8gK
7lnawqTHNKt9jT7i5PGIbVzYiBnAv3L6U0mxKvZGcqYIQn99tI28j0Cuh8Tp
zDbWwDf8ZVHU7RVvrr/G5wo9G9XGZTwZqHsQKVl6omYVuZiywVhH+j9A30uy
mrAh0efnjeaAzvmhDoN8UT98ozQWAxhWobYvKwnDO6z6e0mvVDtzTwOyN72h
oBM/mxAOhnjHsKx+jsCd39SB6yQamFER9bXj+Xmk7Ll1LiviQPemXpD0Varu
6aPdLzefQOOzmnpcnEu4msvwlgfx1H24ocxnhx2SfUK0mZsbbfSPTYALr3kG
9i3p9CtfL37qlTHhxEIFu1cypsBBfWp6+Y+6RaJPw9cIVHDXVhMFGaUqGF+h
UEujs0WnMowF7xFy4rfguFHJ5Dh3YIlZK7KpWM7xzhpq/e49/Ztd8pGg+Trk
CM4XqNLUaYqUYNRKyywlGfIa1tjCDnuBZwRgBV/sxVdKGct7fta7+Z1m21AV
Y4jd+RvvTTrC0iIC9OgxHenyzkBK+fMr5E6HCfuIL0pN0Pg+6ceR9pTnwK9Y
9sZNvv5YX3WQCCLyCFq5yeT4JgKP4zF28DUqqRykNKVoJLs4E//51ZTh8rhW
hjYOEq/0CHuV2z5acaXzsFP+6CfVoIxDsj6L6BgWvyP24VV3xZdNGCOcyDKs
ks+c9jZC30VhUGfDulm66kBzlcGDJiuEp6hNw3oKABRx6BvcbCRLXH0AJaCX
AobwabtrPBvsHYukz7CChwt1uuXFVLB64C7I3TBCPDlzBmlpKDmUYqA8OIg+
Af0ac5JznU5h2zlVdHbdXoyevj1dECujhrGLE+MzDwpm3kOXmyCUlx1tnLZz
jG1QNIN7SR+R8v5OfcB0Soue8VpgfJWFxJsk+1Ulm0OnnuOD/FstOIXRIlQo
BH2yx+cNKzzw8MQXqb/ZqnT8LPrgBoPF6TnVc5VW4W6oJIG2/jsStrJiEAEf
9O9JuY8A+6b9ZivtuHrY4asoRchC0+zrrSxaEiGOt5kvt9/di3/EMXk5vKBr
0McQXW+pcmqSXcusW0olXOZCCoChss5AUrLP2xTX6TNr15lUgmffysdOFKsl
xEaX3k8vhg8feZjgKKqqZ+qQapvI6koY5a3hY55hVRab7mYXaPmciZxu4eOp
d1TGmef4xV1vSaWc7wCU8tbytMq3YkyHr0k1pCavIGAxbY1odllQqyS+74yR
S/HJsLAwHD9TzblO1ivg4VvTiLYKGq+206tUPhBRfZ6ObQ6szoa0JbexrjME
Luz3UXETi8WnNk/+2YvcnylVF6kH18tJepJSGcx0QeTzSk0ZY4hCpBTStTvM
zrLVgsk2rAf54VSOpLebsp+E1F/PtZn0qDX3kab0/d01IHnlnTe6Oybdy2S5
fg2fMzHq+zFAHJbxg+6/EbINgVolQ0yN0UiysHuvHCSaQgARhzhollyGKeSs
GB2WbejTV525y7i66JMrhJvvsffZsPPhpNKF6c9vdHEg119Zyr3dPkqAfHHE
pT/G2Wpm7/A7ijZqs1eo8dvoijOv5Jd/Egqwmt4EhUQ0g9/Pdxm7EGpXsdjc
Vf5i8br+j1asX0UlZbUxuxowcfW3OF/EI4IiNI8/NXlUVIkyCqRpW8xCRUhf
cudjDN9NNxzeIH4y69c8/Sldxmc1zEP4AOdiE1blxAR1SeJPYMWEgdQO1XKD
fLtfXCvZKiGoxcwqXIQClR3S+EhrxdfeVLO+1K+OkY4clqbsLbiWUMY1P+Qj
8fFw7w4MzsIZiPpVdamyuWd/wGwIzdCFC68fbIzzXXnYF0bFGdamn7nHg63i
3YMRCHv5cgZXw5deK1WooH2+jlzsGieHICEzGhX4EoIJIcTM5LJHqgqFPMkX
b/kh2LRziloKEQI3ps2eEJtFdQp7noQxXnvZxXXfnMmo6TVSIyOUW3P7mFuY
tFCq0fFfqzNvQM9KP7OTiFtBC2amN+SjZXa6C2SCWXzHoGeXF4bwze6cKK89
2xsBSUZbhF3280R0Le3A8RJL5p4PWOL3hijV+nj3TFGX5DHOlYC6rCXp5047
6vvOACxE4T6tGuyZM8mrk48dQlAazVy2daoybF7qTsENoOFwJNWxcTFFCjQM
WZcrbWoIQUjnvFWLcuAgwxb05nsuhp96qcN0m1X8ZJAagVHY3k/EADxEA4Ws
Z2yEOSoHgNb2KQ6EJprO98pqBvR9zHF/1QHk+3eePjnHZEYU35bClB54xVWZ
EjMhFvZ+CTGZHN/DvjPC0B1Xwr7aQE49PPawKwtq1if0/KLj9jKZJyh61ZZd
X0Sm7ZUIKyKwZ8cosKYtkMc/I7QkGB9PCWpZP29MToFXRCLLOqrtk0tgivsX
A6Ry2pNZEM3swdrvorNuN+Cd565eQ3EXc8fQchkTdqICa8gdtSMfpuz0J9Bh
L95l8uSp4p2pUlucb/NcCPcodbKdZL0+fP7HSRV9bf2D0UXrRMKDzzjwxcxU
hJh4LtTryUbx3SYPOFFwRmAUNoP1Kzlw3wUOkVo4/TsVfNC+vcW4vfcMr5so
OMRbFyw28WYaE+5XdikT1P8cYGm8WCs8V/R3cxhrFi4iyyvuxm9Z1vmUj+dO
LaU/LCcRFlvW57Ol+hP/vJZriphyA7vI6K29+ygqoMKYTHfMS6EnP8cPL0TX
ZWNFJ+UbLYtWsfDzHpFTU4kjhrrblGIHKAhK8r1dXkZiL8gwsBIgntEJT1BG
rwGyPskhx/R9Pa1O75tdGjMf0qW17IXsRUA7KUeyGWzIo6BHIB3lxW88k09O
DtXUYEDl9EzUJtA/TxBtctRaXOK2WLUsqBtg08gn+xo1NAQ+eAcvb+7lu8R6
9lZKAEr6Ba81KlNwHHE1AdLb1jXPmwEkyJ6ojE903MBZyABImfXhKzjhnJ4G
8+a7KSvpHHbYQz0u0NmJRKOq1QCYlDk+xDmxF7aQ0gZC/qCaf1JHahIQDXww
OlAFCyXO1cOGzgqSAR51//CpA+hiYZvaR1P8uBFurlJuXTPgsnVq7Y38S927
zYqZcjwg7pFGwPAoudfXwwD0yi5DmESjcWYQnTu1y2/7KbrTGS1JAYEzy4tZ
5qjGUbKQazzfLc7Ag6gliIuZ3OHmCPjVnKLjLxK1KVSjEwShRdh5eQWG91FF
7ZlPFYsCmx1Yzzgb89ricOJXmg8ABCJeqa2eCRx7J/3rAYzgfcGqqkfnBCf+
PHW+kNIjHgofarrTWOC7MY5Biki+jeLz0qOrEecwA5TgEyE4pFBHCoVgiOiB
fEfgsFSJ3dpkFBXCQEzkIYE1V7s0H5KF+7mIHmnOiX0KvdeSNGDFQ4mMwxBK
pS9HTcXus3XKyqwLa69RMti8jHhsf8bTec6Zp3npMjo0+nFayvWUfBrw7EF/
sH/d701kkkIp+rMDQ0VSlS09UCwpeOX/vt/nm5vwI56JKbBHn9JmZdUC6U9T
7SXJfCmD8qg2/46rX7gRuqg0IxbLp6M+ZaEgO85GBc/EN2IcEioMtX+KP2UI
5VrBWdi+3MPrL/SpmxVBuGKHe/P/1b6gQX5g1ltMG6ER71TrOFSQOhtsLb06
zur99ElVNEgUi/XtoY8X6k58f5xcEv7lcXx9cMkUov+Ebs4rrWU44eXse7qG
JDzoC4c73ZfNJ1zXBGvitMJXm4gGweC9yZ+JAQAA93WoH5e8Z2P+qFHLgTui
13W7PrqH9HhAv6S1VVawKcjViGBmXiuXUapxR8p57s6Bh8xuLj0gtX+PQ+tp
Lz93laD+H7+iXPL2bL2fYVhqWW5pCC9tBxpr0GywRd2kBZYsFd0sekdohke+
I1VfCeu7DDqEYSlgHuIX9KZZGEnySSl6K73/HrNRLMbiBKGdyHa4atDKY0YV
vXaGuwa58J1P6/qTwV0zMVm1gPjibeCi/qZD+H+ek1NSet2wWKr/d5q9W9fZ
QM7vsavH/dSE5jC7gVtaUvHU5hH7t/vYZ5wOFwcq5sD7/q3ROGfx1a5bNyAG
aPVM4x0hlGTFXtdFZmUwgbSRFtFH5ivPeo3o6rOXPDuN1rjmjjodv6ntHavd
JD92WPAsiQj/lkUf6fkwCTMs+oJECWzpd8x/4DXJZfNYC8+sG6yRZLdCXZYM
qF7uMPKnNRyP45TuFIpaaorji2r38mUOR82V4pRAV9HnsdwdhFz63Geb+sZq
J3MgzTzgOaISqub+5sdanDjBuHh4CF86dP9y6AZP5LAIKs+sjMxd0byKd80K
ZT2B/9bTDyhrfD+LUo4dQczd83fQDgb/Teq4vW6ck7iNF002CZB5rw+vqQ09
BwmZ99kTBhCK/DsD+nCB2U0v90wYqHu5dSv7iiapgU3GIhc0npBLDrqlw1P3
3nRQLpfbgs+HvIOXZMiXqq1Q3jme6AcdZAhyJF4qWwkY8dMUNNyYfihrzzn7
8+mGmS65yZnhUMd4p8ZTrpotPGDysH0Y54+zUiLK+5Ca+bSE4F4Z/DdAJhqm
wV1HIJaw2oL072dnZf+0uaHzma5pPB5AiCeYjMhCRaNKAC1EdKz1EoEd1HFu
GMk2HArV2YncXmGRoelaIjmq3qtJ9sPpKAmYMHDpG9kO7n6L1Fq7ZmJXAc0O
gcZlh3OfMMPvhd7mVl+WAPeCC/+lT3xEIwWhau3mcxpgBe0H/KL6LQGDciH2
100W3bq8uQx1anXc/+7wAWo2v3gos1AP7asxnzfwjlFJk/H97bQyBKu+ZR1e
J9cFn3B+wnrNzgVANhS+C+jjT8T2TSFwShTNxH3esMLezsvaNvaqPrJE7bti
1/uI2C7ghzfhBqsFbMPdEGfgkt3W7MlKPomA2yNQmWYXz/FNbDsW6sm/CLfO
uvmeXeN6Wd5q+XK5b43wQ0zYXtRRNyRjZ3OuH0wF0SzdMb+52VRFG0WuyAVV
KN7cjjPsLolwm+/tVHurbsSTGw7Bqs9uuQpjKl389+jDww+6pmOg5DgPAKx5
Xu4zdFb1psAfCylemSaHf3QDgD/siEE5KPUqIcByp+kTXAq3YgXvuTAP0H/E
xp+R/tV+GbIHCRwAHJQz8r/pJwiou05Gbfv2krhzk0HCY9U9eqJf+U8qSm6m
66aujabDIZEtRxXH0KqMRwgEUWdktQeAKd7XqKMkUyf97O0uyI4oSALc1IVY
walFhKQPaTg6J8rXkiLtXiV3khgD9NMukWjcNoIAPH/sHfom9QWwRF1bQbjn
Gi3omO6Yym+lNEA33dxkBkTTBlzrA56AqAMdUyfznEVryROiw4IVinB0tMj4
jO+U5wqrxEY6v+Mevmu3GfxFldvu3knVWvFWERcYzTxaWQPByjfSG9Z9NKo/
mVrn/CRVd0PE0YKYQxMtZ0sNlQ1/RzThphOcctSjX2SJ5/WaUWXavQw6ucrb
q7m7TVRNc814VNYKit89Bu9Igik1FWs+ae1Lo8u+Q9WS9YfU/ofpEEU7hb9D
1OvAo8VUkJA/YP+HG0D2oLGTOsqMISjxdgACiMypeS3PSydPMhORvh6y9y2R
5T8yvSB4D8S/WqtU9IUDeOQ/cwyz2jGveIIojpHK4stM/dg61JAk9X3luzSD
LrOM8oqB9fZCCxsgFxdhX4Ng4OPGUxL7Sqf2hHDpG+T6TFlQNIBkGlJMnL9F
v5UbUro8RnzAz/LIrnFl+TaYY0686ASyQNHvd5zNRT4gVM/9LRul13y+mLPA
+t19qTHvRVo2ksCROaPWfeel/Tpqu6NqM/dOH8a25qEDpjgvzJ2FabmwXpIY
LwHqqQTBjGp2idXwsm5dFk08IN3kdjfb1kInQCP2AxKBv6Ql1P7hdGMkUonM
/IhBCMEZZHCSSfO08MF11yzfsq3b4woUaa0HyQL2zq1B7CxkBj7WNEos6Hpi
4V6g7bPjkadl5O+YvdPtyiP97TZ1xnjpnt/H7IIgTsbhdCVIf+ir3YSJwRul
9qgF1TwE95vDRRO7muTG1FLcizHgLq39IBvzaDPrRCJF6kyQ1QTZiITLC4Cn
TgUep5n2a5BdkJfL31yV855/2swoctGMhI/aJEmCq97m4FP4RCHzLl7Vtq1D
OtEG4nmwCzNNAd24LsXCCAT6z3LQbCOLGJf4YqjBoFHV6y6lMBkeVVIM9aMJ
6I2v8ckzS7q6869g/L31lz0JH/8e5K1aGbsJABZ7zva5VjsYVApWQ7nse+uZ
5/InYR3SLzZavNtmG10nNc4o61Cv4D1uCKH+1DSFP8SSO4TlFkJFR2SfDFh2
1R6xKT04CnydAnrkOMeA/f71iDKAMQv86H0IF7RQ5e5j/ihpEztIz6jhYO5e
rDxbuQZQaGVzRXA9UXEkx1FIrHTo+USjJtSpizIIFnE5Ewmf8ulTCIziuI0p
jdooKIYQIVmqD2FL1muU/cZke4Iz8Sy245yI1bbIoHNpUeUiqQp68bDC0iV6
+jmqeEiM2/gV+60ENwnBVDBIvhbxrbUkFhXhCABOy+I4tOxIPUhu2kiO7n7v
yOG2y1rrjDnG+B6lKhQ4sPNuMr2HQtVJkfoaWT6sid2D1CPqje1enPjPpY3G
9hakUpSlG6G5tNiIgT1dOrdq3E5phiM8eoDbpQHaHTawSO9IPg==

`pragma protect end_protected
