// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tQK7zLDpAepfZmikqsNVk3t6CLUniuPkQ6B6fffGfy4obSNhf2w/qmnarP7H
fRmQauHiufeDPvMrWyw2hUsaExtVFYNOKm+ju/CCOEQe+gt2GL5WfqbTjFNV
fF+R9s8fzOTLxqxSiElrP37XKrLNqt36PuyBWIrNgdpVS/RkRy4c0zvdH+wZ
XCzeMjYBR3GDhw3oyAbn7osgOkt+80JZMbPGiyJLtNclO1IyoUZ1SYhBpsM6
ml+/zlI9RP2dHmvFbrrEBaQpzHfF5O/Pkn57HjkBxCbVW48Nfo5VHLhyNkta
oyJkCSDuZgQZAOp4UW/nlJa7JcHg3qHdpbmdF9X0+g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
myG8SEgo4y+oOws8z1Qcbm4g5sIwRt/5u+G8FWekoMKUexvTl4fa+ob+Fj6L
T0prW61Yo/qGJTKmbPmjRfOvUNMryTeInpBHdlPdJMcDx2POf2m34A+PVRYh
Wvn4U83iuKfrevZ48RwBDt5zlYqIL5W9ckMKEqJHYLQDjkMkpVU5hnTjblFn
YSHAVQA2R9KBCC6rQocvsDeVMSuIUljX5mlsVPrqwgIpNd8jlcnZBg6rvxj8
Ye9C7bijlsyHdGPJAK6OiS7lr3GaEgZ4rpV282kY3U1z4SgCc7cBpymLWPRz
wyFwENyxLQtQMdXzViC/tQVniJdL0x+HkCQjeV/0PA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BnI+gDCrH39vbJ5N35ygMyqf1hdgvCbb8JqSXsE9RZgeiS2M3jpd0U5BUc9W
GHHOAfgst6APigfGPgG7/dCRaKxRmkHRKgfHxc3mnhBWmfAHZyNdu7b4UqfN
J2XnNpdE6ws2wLi8g/1R3WHxdsrR/eq6brhh7D5bX/KarNLYJQHYQhpQdGMb
XDjmKi4O3uj1n7Xg4xS5ZVB07a3TQinEdJDrVLZCGV1F1mGAryPcBwzhNOq1
C/wYcDEVAMHhcnJQ34XR3ap5b3qMrozm60Gq9xWSJcZVylTL4xBR/wYY2PtB
ohB+8WsE71PyBiRnhgaIxdAoMnsqIxWVgm/xjcNicQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pk/QQfbu4vyGFAgLrYwogIUeln5yroy9SL28khXzGiMgttMS73IEG9/AWL62
XtpP7/to4UWVosrBYrFvqw4eC4uxKlQzokZ77RRxgvdGTzNGjEI6x1WP0DhB
iQbtVLZk1+YJmMYlXYiAdFDPxGOdLYx8B7dMUTjjqwRKnnOIbf8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cRX5qsqCLi8riQmA7iLm+OsjaHBuJJOQKhPCca8rTecbxP7cS+7sTtmAhw3v
3keEQRfDWnl3di08QFL6TqSFfE1FLQ5C8SSUsN3qDP6XKfpjllJSL5u7sqZB
V4DFuc97/T4OFGXSaaVLUe4wjeJEL48O2FBOZ4jat+MeYtDWLnsJse/Eulhj
Cok9YyWv6Rv0d6Qh1rXGrlgj5rQOvF9MfNLAiICTiNGOuVpweiUnH+VbgH79
eP1ZaaaQjA6xqbBMJ8TtjUwGIUspJNWW9jHTthC686aJJ68vJMCOCa/fclcK
oTFbT0ZVP2UySyCOZwSTOl8gYoKSInkLxpVXxh3rCX8QdGhhUTHwS8QRhlll
fk9tGTmX+NaT6iRDGrRpWZZQp2uEryzzfBD7JNDU7AQxEe2izynGznY17kOF
t5Wh1WEyUYKXG7I2vRvOKC0Mh8kBrv4AqCQwGLdZboqVabY5em1a9QR7Nl0n
eDUsLRbdZBmY7yq+XRy3fXzPd9S0YGKn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sqFzFwkJ4kTxUSFjBQfz/NlVtifYxPEylIiEWUu/WUaiuf5sFpVxcZcTI8vR
TOeGTkJWrl01CB9uYz1Q5zmtwt0B1ZrHY+OFmT7/wrr6OnBnU/xqW7ilRKfN
WVOJ47dzX6/iBWllJmo8I9ErE0Uxi9eV1krENClvxgIoDDCV3wY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Rs8C2T2+wLDel4nq/nK8CttzGzR7IprlHZVt9RjetgA98GGd0RrWzO1W8rLA
gL0RQE6dm/i0DUryN/xo2+gyxDWrn5y9vv9rjQo3UTE8z2bGyaLF6H8T/6GY
x7uqrywSN1e8JcVEyuoJW70Y64eqLhpg06e4mZx0DEX5lxaTxIk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1056)
`pragma protect data_block
Qm/YTK8GnFh7eTtIaVeB3GPjUi+TCWFNnNPMV2rpvLCHCBxUM9wCliTD7Bv9
a3b0iT5CZtPEW7I8dzcWvtM+avQOyrQH4gc/gd3hbdYZBxOlsQ4tf1R6/gq3
cPCXlOImlh8w3sveRyMaMOWSM6givG5zF3UY4Lv+Ypj3iNMxnmQ+DQ/qshz6
FCRWLYt1+b7gvLyB0AfgARqMiGN8ZAgLlxsyRqq87TiGGd4lDOYb08H0pkCE
qcgrqVcIPhNd6+9Ii74T5LeW3QMkuLuWgkHPlEPI7Xf6gYIANPJTcOLq39PA
zt9Rjbrazwa4Mbjwncg4tfUBsBW+eGR5dldQq8dG2gzJR5R5LHMp//j2gRNf
tHOI+1cAtk3cg4Nu1uIWVh+hZve68GSR8TOx9DejCMengINzwpR1ZzH/JDmB
Q7VXAhowjDNOuRrv9MnleCJ1bfsD5wL7v80yWb3XeXqMy9rWBzxSYoaiwKw6
wencVYouV9R6NaISgchy0jgjiThsOKiUJx2SXYUlF+peFooVI9E80ImOVrmz
eNTlpeiijabZJDkHMdeU/JXkSRzWN0H6sfTCTIoBg/e39ucq6yzGvOSna79Y
5t5+9TNkRInd6VsXDiG09pXKB3tFR/oBFnHA1jLbMnl8llakS3MSQr2Rgtwc
if056cm1k8jDMgZ6EaITxnNoaeXoFBGaZWiBwI1a0/JNl1+Z7rRFivAYacT+
VTMxTEzS3lOIpDPp6WnNL8E/hu6nQYlcmBclL5M4c2cMrlXsTnnbmWb2/YMx
Fvs3zpv25UcbzOTpFIXxrBe0QI3jNKv9RJxfiT9/VOsHXt7PhjRU2npz4DNV
BKw6Eo+47vMT9mTUOQdkHZMBnZWKApUPOTPxHrALNVhZnAiCm/GRqZdSZB9p
w8CZy1RDu6jCzZ6ETF7NpBvIZiSDMfLnz0s7hl5rwSDam+zhulcgNwETjvN3
2SjXulMYLWe2x8OA0ftcGGxfVuX2u6pBDNuUfEObe4E5X/AyO5Gu7Xr8ylow
uusOD45ToqqMAM5uFTQQtif7EcVnH8YUyraHDkBLDWqFVoenOtZsODQ2pWjd
Ugv7DpKK9Q+QxarBLgCbxDG73ghFDFHSzumWIK9/HBRra62h4+fyAzlAmefe
09WizQxzobFbA3wLvbYqwsDNBhs9wwlASskjcfoozdFEGlLJlysze9b7jeei
pRZkHW2IMNvwHBVrQjQZCnCXOttF3d+M833A3BO5kb7+LjcmRw8w6K9QzVaH
j3mZfqTqui85gvuWNWJRKDs6/i7n8zPdQr0uWnniUM+QwK8zTBhob89i1HGK
Arx7oPXT8jAXBGqNPnFthENwQcVnRsJ3LhrYDiHjNtuSwXQeZIKqwSAoNQ4x
Azdp4rxdq5w2+DGVwtyGpuAiS79i

`pragma protect end_protected
