// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mazOUbOCuE5+Nx92wHfi/kWggdCZBWyP5yZWd9FnPXPq1Geoy2mqTbGOoHA0
v01/aRvDsC7ysLIoCyh3np8M86R7K8/eFiw9Rv2fn9SekhhQu88aa6r0C6+M
GqabRyfZHlXU3a9RikMREDFB4UBKUYpYfJ6+49kOMgbh7NnA2x1lli2bSBlA
lMAQwW5BlTh+rA3VtlG7mFkx1WgeDRCzZeByFiDp+3d0JL9F+Tbn/FbEZ3m6
O13rU6tYlPof71wv6FjGcAyRdaoPq4epKPcm8Uzc+Z8SUdNiiYjBuz3TA8Wg
b8t6n+gdh/C1x3v9Tf7VfyuQJd+P+1nPRr/ZRJkNPg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H/S8dzqxc7Mw3MUxKWVDb3sce5dD4oRJVtwgqauY5NdA7thCglsoGCkdSTFt
8tchz4WF04xPqP2/ICa2Ck0ZU0ZeKX9XIq2MSwaAs+D50hEN+d0wO6heCReC
f+B4Fll893VdNFvvUd44ENCTp98tOcRprOeXqiT9LLmztDBZMNQAifwl77Hb
6CbXWs6+t2ZK4wDzJX8EOgdgY2QUuJfifB1SljIFpDEOcah8iSrHFttnWTS2
jni/+iTIELLKseZbV5a8woWZTMXs4l4i7EfdGVSURr/S6hv4AL1QfF4Vk0VL
ADqVCLwnZNx7OKkjS1FRwhaeh+IlMrjZ1GgYAvAAUg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
B92thgsPsgA67HnPvGJMHsTY4O4lvsxh+EFasPpGrWOr/5fgLC6vRIDgT+wh
95lrj9fJL1m4SvaihZjFDk6RBSTzvkmC//76Q7p7puSKWFQy10zpfeIFOsvR
4z5zzJ7Li1k8ZckwYAAHn6QqH27l5+gUuT2nmm7Z3eNqP2oeVIClcuTfxskV
0kGEnkypRYc1GvYQxJxcsMYC8ZbOazM5LERcv2EuBk4WNxOs9o6Duo7GuTea
ZzQnLBA9+ef3dM9tVjO0VjQaFuKF4kqXT3Km+xjLm2ezqSMq1WFcGy76wetW
o2chQlTt8TxqUJsaadZU59yuYBR+bPQ95tUgNyp8Qg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ui2vVHb565t/NjGyv3nLbMQ0Im/nRNvlmsIbcEKttndcGUSoKBLltB4MJM7s
fjFmEDI5stQDZqTC5miguDXnLdPSwBXybaJXNXgVi47RmDdZf4TXftK7bTg5
PUywoaqkSRjAaaFSWUrSKbxF5StqoCi/Vigi/E/dI3z/XDCxx+0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xKDAPNE+PPHEKT5EHBETxbYaMlMO84kF9pInHVdrVFQmqH63cIvN7nHodwiD
RrS6gOlFtnc+H7iJZkBe213GsKomiQQfy6Y1gGXkNQV/eD3Y+0rcPEkAAO4c
cjiIrntdB7SJV8kCPdhQmEVlx2iqO5RlE91Iv9ZfS6i+S6ybwrqKIs2IhRUK
LmUeRNulblnqCZtEWtzXBwmn2NNtS6Jjh0XurLrHQ5wsuuZp4jjzhJEYax9d
LlvZy+LPabFe2u9IIUbSbuy2OC8DNczBx4iw6k9NalnjJaSN9/Gv+e4inAYw
/MV7DVu0+DRLS2WmpSXg4Nj2Jda/mAdsVhG5MFo7IZ46zm6+pfpZ9jFynphG
5JBzYy8msygnGtkYyIlGld6GBP3LVohAoqI4TkSz8J99LIJVSvIfG4Pq7Bqz
GjRWhCYD5r9L0HIcGBGW1AS0tFOaSPnqS2ooQNlxBS6TpvtcTivlcJcdyY79
QOuTGsPC3VcAtWmKCOw8Tn/dk4wNApOj


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P/a8lUdoJASmssgkoVmk3Hp5lVsnlRAjRC9qV0bf6S8yA0LTH3WovOdvNKSE
l2wv7eJKEN15uCG95yex26d+2Dz27XDJptYtH8uPd1aUDYLnL8mJ/5rbtQQh
jyipGajr4KmT1/h3UDdYLFoZp9YCQdMmHah1W3WQbZEnMKJcPKY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hzX30aVMNEmUYB5LXeYuyfn8bBrdrQ+pETWlr5uULxXA/DvtVMpk70hfKvdj
ND5Z8xR/JJR8ubzswNM54l4PNXNuXKe99FgJczjMsGp5ZUW9T+8WsLvCAz4t
ylHnUJ00Eq1gNFsvKkcZXoEK9OewGlPAWzsZJlDJRmbzoFXRUyk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 48784)
`pragma protect data_block
/jDRSWyYpu10XaaqZuKyvw0hXNhzxxG3Pcuwtw6WnZ46/3lN4KOLd5ZbQQEe
7Leg/8FF+qR7Ut5aaP2gPOtQTN683BxBfReC19m+UUgaWDpHEVnvm2wx7WrS
fC0cxlrAwz4wLv6Kle+bONe6GVD87ynYpLlJrAOmfSlceOZ9s2IyMlSwDXmD
V5JCJX3zK5ZVaesX5nzhC/Cdl28rgq6RgAhxZ2kI8vk6RxFAR2CfkCIvAO7L
whQ4iIUfrD4FCtRuzHAiy+O4jCF+bkQXG3rpf0aTtT6ObvhZZCfrxfWYDZ6h
KdyhRJPZFsDaT1d+9tBth3+VimAYuBJnDsSZiTVpRNeBgQFIjQB98jMOO+sg
+OPtbb5DF8y+8Aao+np1u86+q2JPox0WW4weOoo+i3lXjaJFlLy/XakQpIUc
9j/uqEaLuMljE26g6ilqkzEE7ZGvtqRT4rYY2rl6DbMYDd5Orj+BpNZoEIQ+
cVwqqXjbmCoJCB10AJu2FatWgKjkJJNsgnXngARcXTD0JImJ0O7icYMxWrDZ
hpz46CQgq6ZVHWrz9iP/YH5UmS4bjgLpCgg/jP7lhMN13MSeM2Ler7DZZ9PL
DYp72sh0aOjZQKOAKx0x0SaUM6J01FCE1LsbLDmUKENEmw/k8RZsVaZj7XZD
jf7Lw9TKyvDsHm6LwZvs9xR44rtuv9voUYbN4XEdtSfOZriWqDtA+rzUhTnE
/0I30b8Kw12y0RnCO0EzMVdc4yEM49o340uGfJX5OjaeDPjTRyt7REMnxhbE
Iv0tJZ0HwL3kuoDQC6NMzXMwyhU3W2lQ47+WBtef8SDcF9ukuqIjjnr2QXM9
JECC2cKTrrz3/37H77MYiUzkw9rmrrEFwa26dzwMyzAbZ3EqQT2sVl5XKS7/
oz7vmZLQ6iq1tYIGh0od+7liLKoBQjvlB3/p+6RZJo6Ml65OfdSnNCvdWRoB
FhuRIyfMM0TX9iEN9/FYZmSeOMxMjcbwtWp5+hv2URYpkkNwDTYaJFnSoAmD
d46VrTqR/3Nc6r2ZbFR3a15tyri+Fk05b2UgKT5K3RU5q9nKLZ+tDf8ebJg1
2t1jGxGVdkRjxCO2UipJpH6jyUzYOhtDmh3OVf0Nl8QGeiuxxOX8RcS3nZlL
V64Wi88a1GWbAijfiKAQkgXWQ7FYWWH5aRUU9GJ/uT1q+nhSQytVF7Yr2y+Y
QpegbhVzYNGvxT7rJL05XYSmr1MXaBEwKSEHIXhninJSYFpwO/otYt3hST4C
H6QsSvznhOu7H0NXMfLM+zTJOWlo9IFrA+pWFzdseauUf9kEhZmQ8YyoryBe
4Tjqo1mXPySO8zpBdl2RQQFdDgyx3+VIHnHj5tBMDROK/smf27u3ccGHM+Z5
oxDqzsRwBYIsvnKw+WXl0kF7wQjkKPVmnkJ/c3sGK7kEGLSSaAyfNnR0Jo5i
GF+mz6X3Mkq6xuVn++7DlIfuRLOwyrqFk3gGfN4hv4q8M0ER2RVkBzfJJoxi
bl6VSnP1mecKPlTPQVpZ/naluMKldOcrYP6FehXIt5+b6oriRwmohcITCRh+
2LGIrhFRIOQdK+pXQqucifC3MZmW6mNDswiYMFvGawxUq4LxXRptJnteZYGz
CwUp2yyJ0hKmmdGKZ/oSFSBSR8iLOvDLCvmL9Cl6N48EhlXAes7Gzay6cCzx
FEmSZeMVmuoJKNCNjcRs3bQxQXJXDVNLH/ECxeSFM2I6PFD2qHb5S+49/akq
w3VXEx3RBbh8W4uFNvW3yopIkawQWjZivkZAVjq1C/BxLxg5Rkn3biMLKT14
lAOWfIHA+2YoX6cNjqXIGnYDaba6DY9aXhMJdJ4f7tmDY+lZQeVPGwbBAwbE
ss5TT+kPo8XLBcuKvQsgZqMafZnEty4zcqjfLLbj3uXTlBM/cmEL+Bea2k8M
5nPM01m+PV9Somia76POqnK6M6sdHcBKl1gle0bX/3dA94yV6OrIEedEAnFI
D5M4IrUgtR0GcY8hnpfNz6cVNh7FTln5/zmAO2fGIsT3970P+oYxfY76Q+Ib
pbrO/Og1Uwwx3nmc7hk+D0QMa4dHvdyW3phbH7WWztvYuOplbE0D1a/wnDgv
1i1tzwXi9YO0enVtFaPdDTYVutpILJT4EaRRg2hukx6VTMF9xh1YoZotAlao
G/Ef4hxoSwe0EUnU++MjcpjT/0zQAuzw8lSfbwg04eT5e6Afhm3+GJmVTyjs
a8BaQQ/gJDzqltvUF8h58F8+fRNV3/ZkIpQw4VEd6pDYPtebW+C++UlNlryp
kBJKAWZmtaoZum4J1hpx6D6+3Mud9OSQnfPRZHIHkcmOZ3hnyJIu5BJORFqY
isYF60nGWKXUrkN1ff/NhGxG5e5eUSVQxUaHEZcNV7yVer1nw0rIVSqk/Gk4
SAU+kAl+hqchfq2MtY2DHSyREm5YaaOwf0fNnzmqq30WL7iq+qECo1m+XqSZ
doNO0ruhn2TLNcyKMupsnI4dXHw+POHeueBTuzjDZNdA4Av3iyYkzVFqV4MX
ZmQA/mZVlKdsfftTq7hmbjPTbVCaZ/YI+1fes3ac3tLwpf5Gi4uLyqi2QXg0
OOBBgTUmejQ8o/1AikvEe07uhmyLUrY1k/U40c5SsBtjWfswMnX8v9Wo7CdU
uB2l2gHZXPdBDE41KJXBUczFeGQsA0fYovGzu1kePymrEqUNWM/O2j1uhaMp
nBP+buF0wl6+g8Dz73IlmipSLocpd7b9GNuOELHogRDcnfUTUIQ87oMev7G5
FsPgElv8iA7ZZBzgvA32xv+W/Ngzca+LiGREQcm0febp8Oj32FfU1yugVqrM
n8LQtpeA5pF+AMQ8Cm6uJF2YrEZVAx4n2LMmqd7wwnGLZA9ssPnysnumG6DX
xGyN9pNkukyTPvpVx3oSgiEp4AAQcyXgpNkHKjfkj8uFcn8eDiOQECTYB4hz
JX0MUQn21mhznh2JsSPEvRdtOkaYKbSVlvpii/+NzV09hr5AIRx3kf5QgLmq
QC33aq6H/CSJ72vvdJfswMN7jVpfhxUhVFUkPWSV/4rFDt6KwL4DSjs7v+tn
CNCtyNgqxgqDgIZhA79QLSlOtKRA7/LDL0pers8wONjowIU1e/wxNE+4G0aB
KjXZ5wXB2NqSCMPNvAUofTzwZnw0tsjVN/cnNoEPkODp70VFg23okbDHKVhY
a/LdOdqR+9g8ajzGW6K18vY9aa1XQZ9KHDx5UyVo7Vph25hZPvjPTcDn0rTC
LIInHMF8gR4dbZEdhlpb7TNmVQGDkE/HZkdlM83DVAHKcn01N4KftQlv50r0
Uy0s5bNcu838OIoxmHsFznxhpKN5IYTlRCYy3hGFTfrqQLvivrFRJcn/OQcK
SfdxS2SrELJ71wffU/SR6RdgrD1fMdS1nb0JDUzURsXH0ABC2OQJkvjcovsY
l47EMws/+pNSFqNq3IKhoxrmW7ALayEdPDW65IKa4tbIKfJTQwHH3SHeiRvz
xYPyDvpwx/7bi614FQScGC1NHbrGBxCfAwlTAuSt93SknrXK+7Kf2nhpsSbB
zf7SiGqVX+tH9cSt0AW5qZk2mwwJTWi1pNEgQDmVZRJIJ4ZvH3lcFFJvuyww
WAPByAD6bn8eQW1XFHZXP9Fx/3BlvLk+5dRCxj7XP+Psj5at4pHMnJmYpqq/
xrw6gNmR1kRZ572xmVjxAmllUzFy3V9j/HTdbVrDD7mvJMLvQfjIFZsYUIcY
uVVUKjxajimudW36AskBUu6VGrgV+qMoMKqELy03lsYo97SWn83LOfGewe2E
iGgm8ZT7yfpw+F0OGv00dmaS+AMRA0L1Q5oC8BAMK0+0uptllmj9BrEoCCS9
W5tosMqmhAs2TWrIh2wCvhfdrHHiYcbdRq6lHa33iuaJXvgQ0slGm1pKRBpF
F41lT3evAohSKQwGMI38gz61/asMlboHYq2ElfLEMdcb33re8trQn4UjzsyP
deJ+2jsruuOVu2tGSXUQEJtC7ByYZkx/cK6yQEdIgZRVNuTEHFZA00z3BweX
26nKiLB7keW6+ng3B8uFanM0g2T127np3UcEpRI2XW3mWxSPHh4Kgyn6NjoT
zDCpo+meClvwPA3TAQtBtUj5ect92pnKiWBrE1rlls3LYSzDAYyZfKrP3TOz
l6H2eBpSqZiWz1LW21RiMNjOqfG2Cb2p14NkDA1CF9Y5feKMdCpQYN4SvDG9
pJHu+DH7ITg8VmHA/+jJUkSNlGMSK04n/9ks5q2PL8abQTr8rlJrQEiSmYuF
z2AfpecqoKkuwxCHVqFlQjXi0mRSC0+4RIcvB5owbCvq7N4IsJuUUkxUSjMO
kKu596mXDOVuAFFVljyRXlXT/J2QJwdBB+yGs1sXUsvZ05v8oHhVSmIZ34Yz
62PW4Zvk5XdHOyKZCmGfI7WvEP25AnASfw8SOIZDGCPWI0C/oePxxSbbaWcO
e5pKAJsCtfeojk9pZy9qxNIXQftYaHFWmrnXJsX1KJtOVZ8SUFEFI0Wjf56z
aQTT0yMx9/kEapymgXBqSqPShic7egXm6RAQM7RKH6TJtMXmFlcQ4pu58dBP
wnDGHFiy4yfEE8QS99jEncOf58mtnYqkPNRyM/2ZDYCKU3d4JA7CiUMrvZKV
5aRiNT2VEcMD2TN07sbm5QTyx4OcaAw9wj4J1ytXjAY8GzG0HDLIZ2KLYjio
1EPPYvdd2RkU3dgYglow0YDDDUDWY0uT+x8T2G1ij/3fqqn/otdhO2pTSkQF
VTVdqDrB7od7hiqsfqxFdXerAYGAjfUc27wwyCamPxP012h4oORAGld8EbBS
MreQW0kzeri6E9jhc1j7zAZwcz23uhspmpz4vxvlHBiPnO7GtDKKQWCuTJtU
xyUYBC+yT1peN5MBXwrbJBsWxXjao+n5g0EYiKT490YLexACXTUBhqcip/js
2d44rCR7B6BI6fpfRz5Zz5zTCur4ZsDpzbPlGfcynT2bl9FjVn50jITmBLez
pzfX18JmaCVDaStCc8XCRtOvgB/Q48T/hHEihDEkLb+UkNi3tFQ9pC6G60Q0
V8/Gl/YZjjneOfDr0O3RzSH1gJEqcfBpycZ1pE2e1x01soM2BUaFW+KD/I5k
SeHoRB782GE1d5ULXtuPJ/lW8sMX+Fep2HyRMkILla2BvS4O85PNnYfns0zp
4KRft2zZV8s3HPbeXAee+C0Kk7Hn08WTt6ahQMJZkq8s6ci3iZ0S6OdgYs5K
25jQQnl7yEYcDl3Z+9rsXL5RtlyYwLDkbsv7BVTofhtMW4vCHazMm2Spdk+C
PxvV3Hf3krRaXiHzp5RL4k4I04v/BIyL4f/8mvx5+ljt/smd83l+KECu+xg5
SQ7KFNifwR/GTfx+6I8Y4h3gmr1NH0WMUgsOJGe6yoOjaOiSrmEgUufXoCnw
Ou6hGLWIoqZVLKgC9ETrW3gkyV4zn/UEKgTWMoFWbHSLl62JT+s5XordRmHx
w+uxxR6cx62BHFJ+dRDATClsTqh4IOnddV3IZ0AZV4gf5qDI2FQ2TCPJhbmk
Qq6m6Rxdwu4HdTpbJDCABCpsR9GB80z95Zm4j3BBZpzAM8RnyZTbwr4N4uew
RtxFYmayxJI1dZmRzJRNHjRuyNtLt7UXDI5Cj/CJp+RBkVVRMa1k8as9saDF
Iyiq3eeD28WpGiPk+/sr3bkqdPHJJt2yb+F4blYZaFnLb3VBSwRFXEADR9Ku
4x/g5rKTbbNWKrQgD3WfnjDmjTSCqWqtRp3jJ8hMgtEQ+d3ZhBSMLtOKspmB
nxlxNV83UsRedwjpG0QpivvgBJvJM7CfB/7xo8WLj6B95mXzFetVc4VEg5l7
+V3EKRLik06cUn10Fur31Etgy527RQlZPcaZKkBH9wgYXB9/O6Y8qr8eFqkz
KoMspvZH+h9u2ejz+lz/Y2em19wnDkYcJvy6ZoPfKpvKqDhtw5JbEPqBwUK5
sioxnPf3asjs5JwrtdIYa7vRcB1TkRrq+H8NBWOVaws8YNxIJmqn9Pty6v3D
NOAtYVIubTj/KiNMfQ+rYcDFT0r/sTCFsU1Ukv7mdPRLYPrYRTtqin1onG35
nFLPrgIrRpGgviw8WSvjlc1EdKKrGpkGjrB+UVIIEnR1W5EC2eWraIp2d5oE
nfKAdzrMLJlZBENGmlL4EsTe0Wb3K4dqxY8UrtVGj4OoVwYZ3ijn6CI7v510
Ln5OXv/vbCnnPr6pUpXIR5xpwXin9Ecno7pADi+BL3MNbgYYC+/1IMGrWf5p
xYdy3zGz60RPL2h2tP2ytvK1kf0gt93OD+10EaQmGbV3wmM2qtL3AAAITRtN
tYCD8ZUT5BAzpcUrgccJlBtpdbxOu1S5pryM2nUE5z7vBwM1YvDDDHxv6DVX
eyNqfKni6tnKrC7V9DpjvyjIZ9m9uABHReu8BCDsdPHldDWrG2nqkW1mDXwG
SYobnVmpmV6383aRB+o1W+Qw1TG6d3C6LTY6vjNjcp20svHzz4VvpnM3KUt5
0oSrm+zmVk0p80Zxv+e0fSQtz8mSNKZD/bDhbzjZHmuwoAQ3B2CQNluav0ER
+WYhoGeS98iZfiP2qF/kCguSVyKPXBKCc7JaK8AakrmfN0Cu1LwN7ECsCulC
cI9JGSTDCcH/uhWAeZ7aWIdxlmPkUwZIiBBNMnl9Iqcm+vg0AXnjhzLyZW/N
c/PAmJmyyKRRIyU+Hanm69yrkwXxA6EqsueWFEeFqkLtz+x7b9sfugnBUcnI
D+ZA92b4ZwI2ZSWdZuG/ny0E8wCdsfTM1AJDhfldzgov2f9QavR7tms4bz9q
P1PnBgxQ5exwAbkNHRocZlnO0weZyDBRv9Q/Znz/lt08q85NXDoUtYRrzFSd
7jN6w0Jc0gYf9ojNoZIEfoqXwd2xpLw7gyM8coHr2SukVFJ/+grPRaCncc3S
5IvB1y6eblvIiYvO6dYPsNGMImR77DjSboyf8BMBKQM1Te8Xr3KVlSZHTZSp
ykBovOp26SMlqvgWO/paN5ZnC+yyJaV3rkX1Z0wlPlnYrmVa9ms2eIHoUiIX
zr3hzYMGNSOLK2twBygxAEEzkUVUmhjPR8bwvk1Kr8zkBExpMtcd7YIjUGMe
SkaRdUamTwydwwauDLjYHG09WGIPISPJblsHPWrzTo2hkHZq30AiXWkBiDgh
B6220ysvH0wX5GlU93uTouy+Wjj/gsms64ItzjX6iatXlnMKE46kUGa3cZAJ
UJc+o7D4qZodAKwYM+hHaKPNJ0p3fQlSMk3zGNDZPjsYctBd18/9Tcx16UgZ
WHMhf67/yAEiaLJ7IfHmjpSHzPZ62XHQ75QovLGnR1eHFdntCbfXoAqRL4/o
CwapgeviKpCU3Jd4SdcHayZstnEXWr5x8tlFOHUihxu7H0FeMEF9/KStmfK+
RDmV7ZzW5os9pjEs1B+GKyx9a+s3A3q1JQPVC9bkXgL3Y6XIyajIH9rx+yVJ
UW9mnkXHku0n+c5MMEfFLvpwlUqR/M7l06pY3qrGE77o4WEr3UwLDoQh59vb
jTsO5BhfvobXhMDPWA+Yz8ccK+it88IkVW24rcdbQQ4xxpQcL5nb/I4dsGuO
vkmhpAbeVrUYLDUgmOD7H3ds38XjpcrcJxDlQCMNaMUIu/+g6fLObEHLRpoy
Gbq7VtUJug6fUjZ3A3Bo7ES2KkD0yd4oWF4QSNrRpCTxwilPjak0UsYrc7tJ
j8x0nZs6ByEs46EUIvczWZNaUpLfzgLILptJMso451bd1MMQfwbFRJLS+0Op
DgsdOlhm7SR4mn5glJQwwpUGzzlI3uaDwy8XuSIMVRCBPzf6LGn0h75mfRdO
waGkjeaAuyn/fmrpqEteAEmvalt51lZCXNGpTeXo8TRkxccmad9ojJtxriDV
DyMIA+gAT4g8Febi2AUqWGh7tbMktIKBu2b0Kvu01nQgzF2OlHen9Hx2wqKH
8fNLLgWjrZlIDxAXa0IGqDoEoc/ox0zEiEcn5vXbghR+dzJsMO9iJTIXyAkH
4lGz+xuH/By0vIKcJcfBwjiWO9N7FmLLDjTNMpRb6W833NCBfVPTdNEAA8lb
90a5W1Q6dTHPoin6Bccv5VkYw8Yt8uvDE5SrldWAqbYhY6egVG42or0Fk99H
J0y4N5xpsejCxa9iEE9Jl8SVQl0IPsYfVG0EVntvZVTIC71/UAw6UmAhzVnw
kuIMpEMx6LDPQe4tgbH6Q6zu01a3+WobglLT73EyEJRSMtZynJ0JaxghJQV+
se6JOUL7sKaIiVTaWvsttlNwXNNZ5cOz2uvJYNyi23SuGtM1K0m5jxh3+AHw
A4u+8ukLh9t6OzoGP7i4ucgQ1YIiDLtjqOLdu7g14VHOcM6AACz3rKabxQmu
fyHl54E8aFFkacQskVzBneVAPlMAFr27JNHoCbD06USzBg+QYfMfzVa/3nVC
y7dz36W3CU4BK3s+lZaGfBqhBO4YFDwC4n9ShxPPJL/A6GOBTkRsFv0BkXhm
5GVhLX/kiI1wYAx9LVWua/1w9qB3jQvcuQsvhcbzj6fCpUPEnwXU7X32asPX
7L1JVMzR6NG9RTED9URNcdnloYvghlBLRIDkck9CDjd7TC9ohQvhmimalhLY
+isAZYpht4rfmgNB5dN0rk3h7PI6n1GFlgZIfpjd7VG81NmD4Ll4nPRYxVDy
ORY7gBI1UTZnayv3UyG6KBo5NuO/L+FXumDxyQcnos9EE7WC4eTWCEoKf8I1
e35t8OREJXFouCQJ/xS0W7hB99rhaWPaxT+LCagB6rzIu4HxqFrpT4FNIcva
EgW6w/fkRiOYSobLDSjB7gmIGfLZW+YjuHJ6QlqpuyCuO00ePyo9B19rI6eG
6grN2u8mFUOeZHutgaycIvPwDju9hgOZRjfMWX+8X3WtJy7Fqu2qq1AmrQbG
/osg3AVD2YqFoEwqKTQCU/OyaXiaGE07M+qftnqJdrh2xMkH66xKRWIQY05n
7MyysSx8G86oLMT6eAftmPjVhFixGI+4Di/w7DGPfknCmvBCGqfzgqZYm+1X
5kNJX/zz97qCflzmx/J57z4UzqQbvs+EcKOiA9c9d25DLT2xILzoRfUyRcpl
QUTvlVFIrQ5w65MvzWvosMMzYlP0iT0yDOr1CC+autHycAZElmdWb+I5TDWe
T5rbJPTze51AjFq6MQxYl2l0T+1lDt5ZdM1tjNkplsc3u5iEL1e0n00KTIHN
g+iNg+bFIjAsKvz789Wfc9dcXLnfcc26lLJpfQJEsBHWn4KbZiUec1tNgUOZ
Bhw3g4buyuuZJQl+p+/ysv1AG19p4f5zH52s6u1yO1qx3lXKXiuVlhT4KvQ6
x7JShLC7e1RUvGu5rWgc0Egw3nq6suU6WJPv1XTDzH5Rhr+r9/haxd14qyi9
BDc4cmUFLw9ahZL+cbohV+fhRqoVjRMLYrbHYjxV/0SUJEvJwf1dTzpzHSot
5NK9r/X0xGBQ87J2r1TVvIfdTPvB/y3IVaSs2g5TdRHwRVRI0U45xsnTKbQ3
sKo049XX7iv/TqLKXPX5Z7NDhumQ/ZB9GSgzG1HcYYfR7cEp1WA0Pr2W/qOt
lBOVehPXpYWeDj54KPs5uKXZara9KtV3PqI9UYsPfj0qryXeOSpmVVoyoZF+
MPpT0kjkaDFWLGtythKL/8QKaOVUVhmB5B3pnOKfxpk9Iq4/2x3B2WvU+SPe
JHqf6fUGh7+aZp5DdYGrMY40hZzYLFoxqbeQQK7DEV/hdaLg6dpCyy7qTWVO
UqCuLk2DOfIpn3TvQisiYHR67QlZ4sTUMY7QNZTe0vGf5aSZxmY2D6YoR3R6
bXtBYsoJ7mGUyJYcdS9JueITKFNqZYqxxaLMmyQ/VduHYw8l3TuM/91atzn6
xC6o3eV8Zk6mahP7Oi/A+rnNg8POnQ+jj7ordeubSJznyMVxs2o9f5SHBPPp
PNoy371un6GJAnApCRdhLb9qM17Zcu8TicVmReVj+CdhvOlOHt/f9C9Z8Z3F
Uc7rHgy3sqbAmHyDUTbtypUQzeS+h5yi6SPqTYLgAS11hLGtwjjcKEMEYHl7
YCmEh5KpUI8TQBOMV+sseTctJiR/aWSdv+B2asDcSAIWqZ1pD9YrpEzTHBQJ
9J1aZvIxp3owlAmtSx9rPOhHxcmvtrLxYwsR2+Js2vat7wCiLMG/H6wY62M/
wn/IUFBmWgK6PcoBjwMFizE/5t2ZmEgSd1L0GGKGJNov+zdtWMlm3nh+27x5
midVj9tFf1SLtV1AzlCF7WUfYeZcm5p9mfNK0e1Dwe83T32LGs9TnDF3D0TC
5hZm+sBfLqqsV2LAus5m8br/vyzv8qF3UpYg4C0/RCtBHcei2P769cbc639T
2thFAHU4i6GveydFWyUP0CqgDSqUlOGQxu+HfyfPG+Kywk+PAixpj44PwuYy
kiQIF3Q0dgsg26bb/itXoHEbRQTccS0/xw2tKbJz12R0LG3VEXOc5b3O2FuA
81MBEtZyVh73LZP65qb12yvYtKuYQUrr5zisfcKipsUdOVwhNa3xvfLdnSxy
V02zZXffUU8SvDyoTgZL6VDnplDA+pe1w/nZwewA70rpWOZHXZU8gWnijzkF
wnU853heh7Sqa3AD1xT9JXpZSxAOU9LtxGUKGWq4QAlWUrpbIXw1Bmxd96Q7
Q49oH5yZn/9swRJLYwQQnzSvvqSxbF1ujNoEeekGSv60AeZtliNaEU59BD76
4M+5vvwKaromtB1dz3yNNz9m7EJtquphSkdcMfK/Y56vIcBXaaa+LsmLH2+k
oqBZJxklD5AbRGhAtRfIsPQoaB8IPamqULS9RXVcAIdaYx61GJeRH3efXuAR
qAFuhMMZl14ekTcm27EOJvuA8tHOEeXczJhTWfy8hZDtYr+kHYgCCdweJOlP
zmQi17rW9aUpIDtsYrwiqE0MA0/EdrDsWeRsp5Nwk7/T5sX3LNPMFOLfb5ML
mVVloMJa50V8iLqgafdob4rHPLoKZ4O5+kxBjlx1F0FppLJiYgj11GlkQhbd
kT8z42pFMg2DLdrFrJD1FOp75YHBG5p2o3/qHpw/601AX43APuVWXYJ7zoV8
1qVjJa/I6bf8Kmre0daIAU+tcSoh7kwTTAWlSilmxiosFu7UMY1UtdFcFcJW
BjPp/vbTTwcY8UBOSdbq19NLUei3XpfqNi1QYcZ9l/FTTufK0zcs1dTZJRLp
YiMUsVvDjMMdS1dDkfoxj/mArjDF1Om9yko7uH5YMFkNEpYgwhKIVtod5QZL
JZnIxCLERs6RcyRv3/ZmWp6m6CreYcLNXWB6ajPg5sPEjor0N3z8q/geXss5
ujsRtc2poIzy9w8/5a2RnZaZEmnhyviEMkOoLhVJP1pYiPBCJADt5fRnkYsa
T0JzGjAHI9gBwKIGBDVfz7sHeNEAT+ITJDUoXC9QiltCui5X/MLB6jPF2CVN
P6n/ODUtj/M65ehFNv+IHy543PC5ST7KRVOlqIF2k91V8GbsLPST0nWPKUTe
d71ftCST4/OXGMxwVLil9cfbUoLwKILQ5nu2NIpFMQ8IxzYmoyvPFrT6FRWD
nlZIAf9BmSZHsCbKGUeLjB7fOKk57f7dSEx0l3mpP6eMEgLnv6xgjdLmBQiM
ElDVi2t9nB1gMg13GZKrd8DXm8MuckxrvNSq8PC8O/NNA4mymlPWD22OWUrj
yT23kCPyEhqlbPHz3ByDpUJywAsZ0lX070yYbeJ6DqA98uCH86/C12jAg2S6
yXqJYa4CdWHabvDcr0D4AkQgn1jbUhkZsAhDRQ3t5UoLEpyTgI9wTGoa7c66
hXVK/HboSQEWMYu0HqcxJe1uIGCAtv3YwuSzngViTPWn9yLK7jlyxiGLySz4
ZASzVGYnWxO9Cj7049EWww3apdf2NI1J73QoJFBU8/E/nUmvjSNIrNANL/Fd
eP55N+Xn/lcxGfuw+vKPIPa6IAd3fBs2nqps/8to950ZeVV3lcFCk9AP/HmR
xMRzaF+R9m/F6kdR2gKV26MiOofc+Zd1RcUq9zKM6n4SYKvPYJm5GbvF2HPP
HxVLXFj9f2tQIrA4/6sy4xuktsY3xDr55XXl8UJjW8e0lIyuXjMtGK3dzcO8
0//9NAcu2eOXECwkHZNReucD33eFAX8zNuzz4hTYeYidMZ12ndqkqoMKtUeA
mrFdXWeoj9k2TaTCAAJ8fEVfeW7nXPfr9VpuJlBg5s3TMg7JHOGyrYPomE3f
uiQ3iTzBlcOM3s4a3OtSqgjmKvIhiBLQV3adOQAqwBp7aHMJycCy5+0so3GM
x+H44NHKYcB2hC+oPZDMoGBhT2Hq1pNKN1sqlpKuEBDyjdWPS45SxuByLXlK
JF6s0ZSRXeXFkZLo8szyr7SfgdfuOwdz/5putZBR+Wg8e9w4i/FDdMLAzMB4
hYWEdyXUnuLdjXQU3qf7y9M6ZcEdZbsZMabgOHSvzZ629+EjzsnJWDYTRs4c
jR/eOfhtoT40QF8qVI0a7ca22QjZYy32zC84/kL4CvI4BgUP359psMMjAUoD
l1p4OZox6DHmLCiE8dZOO7yIs57Tl9eMs96RbRFSA6mZYo8spvg1AK7g9qlU
jMfSzN7TPyQ1sVGhBWP775K82+7SsjJnd+ijIVd6yovjbCVF8PCF4ctzbHr8
2k+6OQeiBw2z3NsoyI1JRDdnC/KI07lDdU4QB/JTJ2g/34//85EQNgcYGKW8
ThdVbbuVXF30pFDom7e4uuV8vD965NE8lsBLj1+4kdaRc7iLoe2FAnaaOqVm
NQNFXYDnG+6S0ShfvkQoLp0/uroqIkDsVtKCF/FnhmRWbyFMg78jfK+mghPZ
xmVeMbsv4jmyrONKrbY1YfRqUXwZjf21wqbaFLIZpHCURk9+2yJZ3EyZPKaP
KjVVj6CTG7FFD+Af+xczIcBgt7KnHHJ90I+osP6zQ+TwYAQxn/pr0trm45pu
VO70b3qzVPGbBH5A8tgQSpmyJwiFzEucH4E/i3Q4HHcd5aTY7RGGdw/56INl
TwC2NuXaVAPrJURlWjoeTXMs6WwEBRN47PRYLXXamk6vaabs+YsdsmlEosd9
/oGweDGo5B3cLPf3SY+7HswPYEFHiHl3iruQPpxic6BDxFlDiQtMVT2ySJyD
tPTsgfrWhB8LzZrxzdZLxiSpzYq0NCy1DwJHQ8uWYZc5j+1V4dW85IprSgDZ
yjtXtSiX0huTvLDUyVCvQ+ES6+rARo0Sr2B5Px/gT8XNA2rpcRFzv3R0/dpS
jR6V8w5k3hZawiNUX1qFadD3Jgxqvk8l2p1WTbjUlOpqSMgR1jdgoDn/7Mtr
QzUK/ddVdZca2SX7KitGVPxFw0NeZaKKNpPHodtwADPEY/b2AXoWhktFRQW5
SrQq/QYFcTV+RvFj1ddErFoWSDt9qWismhUQzG35XmKhhvrXBgp6XJ5tgKQ/
uD40BVdIF7Awo0RTEcSZ/74Sl/cfFAnKN24Wx8OevqHchOwrLAUFETzugixD
pMUeKnEUvF4uAvYY3e7gah0CRNTn/MLOf8Hby0D+v0+mEzg7n9O1n99+YG2h
Msob/YKCCcOLbFzHGeQRcmO3wugjh0El9hkcMRqfhGsx1aZN2cGsWFuaDDqO
A+wWxJ1J9cvIaW9z/I70KeGYVJ2lK010rH6ZB0qBHI7twHM8naW6xdJF4X7r
Mt1OJnI3QQCPd/7gn8cXNc+pQOGLQQ+zRqBiwzGFJL09VBhqm1D0jsSB3Ver
9+doAhdsTW8lS0fxDsfE2aEuGUwKf1ClJKKLRWnkaJ2V3mjfNVMrWA4cEsHe
HN5rbduoesFO2Uqq81auKhw+dz5UZ40evnEZ1WJEYIS7eGz/cMG4GDJ1LW1T
LZLtYo4i6mwCbnpaHN8gBBa+KppgXVwyU6MgBMbEjKUxCTiX/pOKCHtjuCu2
Lwzpdh1DYRPjzxgu3VLNupphilES2vzfCxtSwteqdhImc4KP1AQg4mVO+y8n
kllBTZxT4MIOVNY3zzzC88Pqb7N+FliUAll+U0TJFyiXXTU2zEB/u2HDfdY8
ojocejIrQt4+ULY1nJEs3k6T+dR9QeswZJOswCi7de4gGK0WuUVbLb0qWUok
gV1HdgjnAtJU3pKJKo+1vEEvTv9mp43d9yLc88OSsQykzZhwo/xxIZ+lJltG
FspS7Cc5G+Ikza6ITJtAFsPd6Hc+LQyq9u93f9FCt1W6CxN5wTeml35LSzot
g9idHWJTJ6UD4AiLnuV7x4fv0y0bcjhZBooPf9yRFmmQ7M5w9Z2dkhYmk02T
4J4EzlMhVlSKDyhelcnUHY3y2sVwYEtmi4GWrGqS48rAK1NWmmXJ/NtO6LmE
kSu6uFaXewFZs/F5jHvrkWHSNQ7rBXxsJNoqolv4N3XymOmdJw1Wdl/kAuex
t5CTHglRcy0SOgiuqEy3WYDBvxF57uHvk7eqfUB4mlW+2eqs2DL5vgux/bzm
UK6EXRtJEzElc0ZwTAIA2mcDGukxxekEfxIViw4c8VKCPZ1AQ0LhZw5IdH+D
ysNmcVu2s5AABVMZs9TACA/NLZhT/Yql/HEbJt9JjiK+mTKxSgyElWTLkM+h
+9YTGiMJ7fCuWxE/8N8V2OZFAcsk52gi5DBJMfzZjw5800bx08zPyYH52Jgg
N4BC2rxH//VFYe0Pn8+qjwWYVt5RwjFsJvZiDJKeHad4XsycaEF9nLhDTyue
kdo8YfApj/0wMTUcgYZVR0XuA24RmeUntyiYAyHDIR3lDW8jTeBIE0qxAjqi
oA/WSM47ie59Bfzc37XEtyIxP6qXEnJ8SuhWMbQ6uzmGlJAbGqL0kRdF5pkh
Xa1vc8WDc+Ad6QNRIHcnRL60nEdiht5P+NmGVJRKELsosCUvWQLTX+4euS96
71cEOFwwDm8m5OYld6fUVBl6EjGaLLrraU6VbN8DixO8ygQUCVG4Q2OpCgtC
7ddEIWmWY7bu3BJj1+O7/sWxSmn5+FY/gMq/u0jKYKY3I8XXk1WoUH+U1xwq
iqcPFod2GIwp2aU5WhgdgiGdbtBEzU1FrfG5fQ4VH+Z5zqULZRgZh53Ex5Cl
D0awO2iKCHZvX+H7GOdmQh1GEcFnUsVwNwX+5twOmcftkBkNci58ldIkxHR0
XH8dboX5lW85v2HaIcNe+atAudMc9YE4/pMEssfrZRruQpb4jKM6W1m244Wg
BUWTgZgb6XSh0BDQrdQaSTTCaS90pxyVJrov3WIO8fo6dlQeohMX822KPWHp
kdjY00EchAKvVyZbJY6bH2tVCpHL0Iv217UCgZV0f8IgaiJd/2PJUYt2obZ5
tlcWUTEYt0tIo0ZKO/XrUZG9cEKnRcoc6eTy6YLiGHE4dlwwoEVVs9HX1T2S
HitI4cMXwNiN+sdUWMmLsrgxZ0G9gDk8Q8/bEHb3SM57OX9PNyJd1PXDLjnl
v6AH4GYP2eueS4dMOjT0aNqDUrbLTK0amksQ1ZBdniZJwDAYL6EDn+KAObVY
4ddQHd2eztdmJWwXGzvZp2wX+9CZknOrUfDuTyXnLB3B4saTLbZ0fcm17+4v
b96rXswfg1YpX9d+3KR3c0fI0k9/q1jj905yWgN0ycrku19shATmL3CULqx3
puEDxvZZFTc4+idrHVU8hnEAcJcFmQtJLN73ZctsNuh+sq+3vyfsNv9xQa/P
np7tuWY8RJuQWV4xnXRKKb8KpqYwEaupskEAVtOCfqIMGvQaUCodY0Vel2Pv
aezGIezpBax1p1ghmNTO7UNVueOm/9H2K1pvRJxe+MzXJiu6moWtwz4a8fy8
li1tGK+F2Ei0IM5ZoKnYGN/9rWHutdEdtevwzHFC317YE44KVufqNgpdQnK3
6nFp1jkbt2FHNnskqoWxh50WobMdFHAvqeSW5GJfffUavi43/0MV4PvTTOco
hG1IgmbL8GcGqCH361mD2wdBL8eTlfmOcup1XYHmuaEl5nRu5yQQ7H9XwHBI
NbnndRqQG6kAs+lxD/tJEBKlndiGyOwVq5kOu1j6f+MMClFsSqBywTt8WeV7
jq81yj1cA3OkLsxNmnaeXB1q9XyUgU5t3b3N08VBb9TAlbqcg939F7wJE/Q9
lpj/06L1UAE6/Wnpz3LUw+i9xsIbAZu71gpQUYcUy0BciWGtYdEydY/7lQ3y
YVWGwqmolSIaF8FLkjZxh/4i4cTrdExT0cioNgjMGW52rCUsE+Yy5MS+sUxi
k7ODwHnjb0UUPdD/MIdnzP8D8WU/hwaTfoThqtKdxBW4r4nSXBrzs2gPaT1h
5cGW37sZYJV7YiU5rISyQ6WkmbRGJppEk8NpEJ2qka9Wy6lEdn5yOo96C8oN
b7dZKfMKeyUuYShwL3z5BouGc/+dcR+XOod2AkqtklJYdc9MTLrlecPDieZU
twZ72c6Bgx7Xj4TZr7cAJYQzYM/lvXE3M6/1qBxHGbOBTkmI5pY7O5u4OJjU
ve1FJXJe1DISPZeoopxx6i5J5NnzGOcVrMUox0ES8GPL56CtNLUTRDPvs6kH
YARFuH+V7CwT77/p0pl8ekkBRl7O2joWf8tVmyy8h2QMCnQbC/tjYIUroTMq
sBz4Dz5QEVv95cL9Qp3Meo40+1mXUPmVPlc7MmzwWbGHoOGj3HLc6TxoFSpM
yZynN4jf1b1sW5GLg+Rj+mJ8wTE9ChCN4uuCLRNsZ2stk1tjON3vVPI9/Kgh
nqYFI14X2PIAyz+JrkgUixsW/hkU5BbRt4KqwAqfE2LP6dCWqzrs1ELaW875
hjYzpxs9Ocvuakuvw402pObkn5gQh+cjHJ1mz1/DjZvH50zkuTSkSSCupIyR
IdDenktsZzXlHEN8xiO+YrPGS6PovCd/5KsC+4erzQYOFVsKQsBLtiXwT/Yl
Ae68US+Clg1OWnwSvwHzQglvwyG067wOcU7+Jv2v1IReTmXF+Y7weC5I0Vr4
3Y3WVTGFuAeicHf1u0LviXbHky7pYfvzqGqlB3R+aOIUksKWWZ8Xi5TVx4Gf
dV4pVRSz5X3y2nhb0CB1NV7ClPGcRIy7MqB+5T7vgFBjVleUPckfpM9eOT4N
8/Iz/eEtqjZV+zE0TKpbonP9ocPZF+C4vzQg1HVTxFR/mIt5OcHK3Fzya4eA
EKncSRGBxp+1oVKECv98yAMRIPAWjZBhkQu8tRFEqES86wa0VG3GrPsGqQ2j
BQvzoS7p9aHSHF9l80yMB6V6smRW2+KIw1hLZs0UmQ/10gNl4AAcQUE0uAdt
g1CJfcO+HVvLUtF8Zp9s+SfSZlmnEG8H49b0LZdWV5v5BrEopJJgVUNxYflH
phtcUKAH7Ed329cjw8C36sWAcouV5CYaQyZzqrSpAmv6DC6KtvIj3jB3J4ox
MAGV/MqjnQeUwLDYqIbWg0guw6O4kTtmmO78zAoE1NWXU3OD17xgf3yNNhx6
gvFALMShb3KBlIDIeReqSXt9xIg5VGPffBrJFoE+7egf4U2lvr2USNV1zXBj
qC4F+Vvh8rwj11TseUlAdoV1HXbfhu80qurXNpjWvfr96zqaG5IK7pZSwLH5
5tz7yyEGk9c0BBN2MUq+Pva8xGCmIqAO7Z6MMObKrBT5enXQBzvMnQT9pwZS
hpFQrG3bVZGNyxXVeXdNiFDrr2xVTqOR7SIpfrNZ9SJjaTHYsLVJ47KoHLNY
rjZ8KiGdXlsIXE/Rgl5+9lh7WjE3XJmc7sehLXAiADguY6rJW7zNgo/d7ruJ
s9V2l84TI5pWDdRX4DRdm2Nbui1Hm1EpuZ8cyaBJhr50itDRvMhsOmgr+hNB
1U6cOcj1oY7ANxSjwzWF7583zponLdpnr2NxDFub50VP9jpIMdOhJeZoJ1bq
TWf5abe5/AXexQ8DOR4h8ymc/LDiHoL2x7uC4xA/8oOYs9aN9t1PNu+xyTu/
DoqfdogoKyG+ABMz3DN2pF9zJJpPezsRVc+F0xVYBpLL1YeXlhW9GxaBwZBB
ku8c4qjZwAWWIexzF/86rp3/8hdMHvnOPX2Ogiwh7xpS6Xv+YbsmcoeeceBT
UNMQ7h3EeZyBK+Pb1io//35o7M3+5jmxr+DTusl//cp+oleBzmeM7wEmjAlm
JHLrslRiRyseTTeUmXuV5pYQQ6DiXkK6mlz8LJqteD9MPeMDmVa/Qu1BcM+O
MP2k0AU1aNeZBel0IaIJBed7KbAMRhWMN82xgw32LrLmkqj76XtutAHiUoLy
VwEcbS0krwR/+2wG8wyEBI9cYaRSauAn0bO1JUZWsPi90tLsA8h75IKwC7JF
bgdLGUrsZAsCZM6kncz10Y7AVkFeqcwSe5ypZlbHAGjnJE9yRW1KPBemApvE
9HnwnpiCtL54SUCtfijCuaWW8tCmEKdoyDrhsxYBeEo2FUbS0Fnm3z3x8MH9
0JgsrWjaRZpKcow58Zr892DG1QoDm4Q4Yuo9oiuUO+6sfmam2XXbm7tUo81e
c0l7hh83j5Pu+7XQbE7oGMvZs1WeiiSjUsO/Y2kKeaEVAzpmQvgq0OTJjLKI
OL1PdLtevyenq7gfs/+G0fvDGWjfV6fqGojk+OZR/EeIU30Jw49aTKQ9l5yo
uMI6nEd+Y5BZqD8TKG2ECszJfZy09x4YwSX8IcpxMxJVN8wApESuAkhjtVIw
KIZV+cEirWh5pST8Jb4L29lqnt1tR1hVKfzYqdb8SU0dM7JrL+Ng+lBT8Bs6
5ovlO9CklmltPA/4zSqAWL1TSxo8UY7uJ539BvV69pcC8TKO24G+53iSdBHX
4KDcj/4Eogzl+iug7zHXk5rIWUbyRboQXGXwk4ZZUrVB9gCoEcLhbWCTB8WA
X/xLQH8qL0s1u2z7qPl0tK2G1G0OZreg9AsPH1EUrspLUbE3oExUf7hHhidm
dXx0NCNQWTrEQjHHXZNm3sVAuC4sBDI5zwBKIxzgMkYs7YOTSImkAT5sE0WY
kwEJF51DvqpR2lGP91evM9CnfkzoxDnJsLveY7yE6e5Mwzv6CZmD3WFl2OSU
WmAFJiZ3JcIJ2tcMCAW4RJ6QHoFpJygMWLjYGb+Z64ZsKcPx1758nLDahMUG
lnDPwPq2bhxKICSmIqfCXYs/55hY1rIV5mtWAgbELoqKFqHiaPF60CC7+Vu3
288mxhOepxHs0ojTmbKnPTdpfbYKaP2cEzHL4R1nlmtIG+gUfunmp9X4MCU5
FPtxa7pziYiX8xNSsVat0LpYLTO+DsPtg6KJEwCeEkFxF8TPpd2H+N+6yS9M
mTThu1JI+bXABr0Uk84mqRLM3NQCSIBUni8ONAotehsgh1BNCpogHhGo3Ozw
2H3WnNZBVKDsu4zqjj83uun2+YReCZ3zG5rltBSytCb9wnQpBNXgedWoKI3h
9Ju2OPh7MUvvav8xByaoW5otLLxcAuh34Bcwby9Sps/18//RHA7IKs6Oxk6X
F7FLrc1H4LwRlacyHEqlVGIVCZT1oY5VUKA2xq1a9W8YcYupJBBxHegkTWez
ORb11KpxWsXc1li7PgX59xEZDnWEwKfsvaor98plSe9Ey3MqVe8HPEJU7tyz
/JhYiAhSoSaEMrE63JttSTHMsdbvEDh1nVv0rprV0hGqjAPB6Jn4asLiQqyb
j0iKvWXEyNnlAvhRjhVJlX7Zg5dnPrsC+EgqufubQEzO40QzcUqY31P9EZsu
pGGg7ltLWKOzVtgig+HTIzyAWNETHBcrJ95WaAL3EWUNzIC5uGtt6h4JwYnc
a8ZJ3fTpLm+Woik1BZ03YD0oiW+8ssLEzghuLK4YHD8SlDovpa4aJ5rSCTZM
/cRN0roHTD7cVMOTuSY5WO4CQl48PJZ30nvxWGT0ewnbM+S2nl/WSuGJGDOo
Up4wfiXo83+O40sbLy5e47wQNwuYS91EvTjzUA/n7QgCKvtnc4A4hUMm1Xxs
EmL/RiuwLThnrZEHvzrifKn/xyN12YkGSDgFfPu49Q28QM7H8Du0PAJq95v+
t7v2jWUx2Fw+ujQvMorMyh0ltEdFtLBe/aYOhUj+tCA8abK5x8LF86davS3f
64XvnLpdrjypUL+k/f2ElM9szMOwoFJVDbf4awr1lNNJO8KUbS9HIaQ+87tj
5cMKkVCtIKTIKRh0ZnbGAkQIIOdjCD/Kd6SLLNeY5UAAhFJQkX5vO8QrQYfo
tzX0ZubErfZ4QZl/CXE26WPsd3/wtAEtHgw2O0rDD/KqaJl+t5P/KWQfd+m+
YeQJbhnjWxgTzfIW2EGNvSWgg6MnstKVyHt1xPk7VkXEN8WN/pM6FwdfHN73
fPZSixW/jcSykCcGN0gI4p0nPySYTtJETwLMWz8IPnu9t25SG2SYEWQE6TzJ
cLXc+Qcz8zMPqF4QDi/OQKD3Hw2F1W+JniqJsJFoDxj8m/NaoPiFW+6EQR5/
vNQcGJu2/JN/0Cj3ybAzF5upuEHIZaq1O9wKs/1C63TcW02D0cvzJQWWTkXS
u3/jpcMiyWHAfVX7qIBtXHBCXHo6FoOGrddRzcFQvL2+kJK8sEXvgxJAyCZM
mR7V0L2XUPpmwcpp+RJlrnvfWYucUNnwhK/u7rGU/S1C6XigMNvbFP1JJK7a
PslwBPhj08CllByNbImFab5KlkjAZlt7Ue1cWM3W7nV+KuLim2VhR/dXQ4G8
ZykA9WOesDCBUO7MGzUvx8sq+P2T7h5uYZVYkqrcQobGhh34YSMC/xYnlnqJ
Xv0sRclYN6ZbuOttxganGBupOuWAagtwllGz47SDAybMA7TSqe1Ldfi7btCo
TBfMTMkUnlinzhIU1yj1jXBPff5bsHL2gavMCfSn+0DffnkgEgVL7cP1P5hl
D2ICCcQQ1XQzqcGHAy0N+cZRMVrlaLeCxJ4TSwePMt9SSvLDDKViuAnRMODm
DQXsK3eJ/iX8jbJo2cLjRFEYj+3ZQ3Jm41z5fSFZ8DtD1mM23pIWqKegM11o
AY2//emMgOKq30r7+Z60nRDcQjnUMg+CoG0eJAM5hR5jA3GuMdEAL9t9tDR5
eTiUJSZKh+UQYMnngE/MOq4mhvyCCIfgVcAwugy1XhhACHRGyq453ekM0fED
pSpTyDCzVJsU2EUSVqIErrc7v+OVoth4oOdgMv2SNPAW9V+YZMrAcNEuHoX2
O5zO6p94KYuV9J7JOyj6jxgcHITlUvL1P1OkS22bW0XjD8kaG8Tz0Quv4wHc
oIoF1UNhLcksxVoU9g9qHc56PX3T2rxcM+nNo60BEsYLX99sCnFm6uvv39bK
1qeJOflGnf0qZwqmteGgqfCGnCp6uf71hnp/SXCGtAenZva2OAHOjz5OXrZY
VnZwTuySCr7Od+gAfK2HqT2uK8RizX9AD0RPm8V+roFcjLbJUxXCPaWwgo4H
Uv1KzJqtScIkWXlI0w6GiAozk3PQuyS6P4Xzymhi1VdFQP7Psu8Wbn6+nDRK
or2AHb89G9TQfjygbl+ue4k8Kn3KyaZzCPEf5bm9x3qcXmtKlaKet5ET+kY0
j77G5jklngesK4cY9Ob19dAKoQuVz5ow2nU89PfCVTghlJ3RyqYmPZ25IczP
bMjhALC8v/f5LRUOFePAoQlFf8uzYFd3YCRMMiJSvXz6RLHu5Dh6d5FTSWLX
gZtu43Ja36Sa8FjWmP8YyjWzMYvKN7Z8+gsBBy36BZcB6WviWdWu2AYHzY8s
d9P4ySV3QUE/lWQaBV4rzCSwEGVj+rKkOkRXg1lcCsBc0wwiTIolLOFA1QA6
hP1xZInP/j7tRuN7HhmwZxOKH/wccHmssC4K1lsZKpHYaPcir5gYTqAxmeJe
EScQkbyNnA4kqpCJ6f/xuzHviILB1WwabzW/iKcl8ZCK+iXASSpBru1sTxeA
jNgt5txA5PRgesteoa+Q2ifd5C7t5LwVDO56U8+IIwXUVNxUpOpbzOoFDskD
R4Qu8G2f7KUjKCwagLe8o4b5cln73zTgn5ikiWSZ2ki4+EgoybZWzRJMQnhc
TOrctVSZSBs/5vPLLugi2T6BUyId9KsQrHT1Vorrl2NmiI1T6vp327qFLgze
ujBMRA8b0Gbirk7bsjiXoZhy09lUpi8PhWf34UyO033LQQgBrSCAAMsic9Ks
isjRnL050ZYdxGzdWqqy3c8e6Y6LwJRzBRaV8d4nn8+MTQkJD31AAhgxiNL/
6WS4jD1m3M2UujORCjT16wqblMPGmRzLjCkxmyAxOkFapbDuf4ZAuxWvBrqT
86ACgyBfPZrndcnnHX1TBdyecKOqZhy6uYGDCFupwdborAFz2f4Zv6i6vQNV
GTVaLi3zIj2YRJeYdddYJmtuiXrVtT+OCmdBSHrGXzn0w+Q4zEObvuyoczBT
sjP9ALlHSj/1PRhPUEy+QG2majVJKOxDVChC+Pb6NjzXAGBdT+eVqJQRJjNv
zApAuuTtj7C71EYomAu89F0JFTQuV+M2o3/ksjIju/bNuJm2vx+ZTqMKSgAp
XvkVZSQTQKjEJzx5TIKdXqAV6DfLuBCOjuL4v2ojhz4gQV0KQ339oONd5Q/H
iW8x4qSvnZKaoQLCxvDicS3pSek0kCgK/DXCX4+BwMj1MCUJn0L3tuDjXLQE
ujJDk46eG/sN/G2K2740ttL2TV7XtzshKmhSXQJ8PdIXK6ObUukqEzIs9Jsv
569wuk5luW0Xa+pFxp0NNYsXHNKpVwVdbtxAsUev3QXE7PtdP2zXBRlRANn2
bCl1+Qj+3F599FgYMJa6NuFzbuKZQymOv719yEfipire4mYwoQV602gi3ZrV
ZdMFOo3VnytKxtZ4VbFky+DpgI8RO4Q96lx309PNu/TKX1lbmnc5amf3oq/6
UyYq65BhCou+7TD5RjO86qk9FsfCLbPcFuUOjYB+AeQfakUMchc+acp/hgeE
/SnKHFgtsQ0Nt5/Oc8lkybQv6mbr8BgaXBSKoMa9ysCbO3dZS1rqoRRA15Rn
Iwy/MruoLYM7JnkfpzLjfRoGqMDDo0gNzPiCNQ/WVpCPQip+vvyc3akSmLAG
qj/kWgttrIVr8X1pv197y1Lo3LzIw2FxFF6sNCO03f9Dpxws5PuiKGgU9tOO
LNMIZtP9dwYEqnSP1+2Ie87sHEAld8rZzOHNRrtxm5GvKaXwzKMB8jmXzXC/
ou3F4nezPUBjl1AgfMX7rFjISpPeGkBhfJwVHff1dpWCjQ0BZbpFirvEFYWy
73wzxGB9sU/wcHzHFCPRVVqolXzAnpPsi1K8YTsIKhNe6TWB9V78ci2nhFoX
tWK+w8kZ6FwU2fJVcGXLMKRn2HwZbXYTrr1JiEkv2GjJCgDxfwRCqI15ZaHK
OEIpcmD55qHjw/4eDU8bU394S4UenLPO4JYo4tkJjfB0YlLb1SM/e60yqp//
gsd31Gdrrl4LOdAmS2xQ86EEuAaFfY6JqYMHMgDnNAdu0mgf8ghWOhmDU109
9VnfIn+aoIh6Pr2guQvQTXNOPuhFCATEhIOeejdV6HeDvVSt7RSRkQ3NW9nX
AUjK5oZC1Sm70SUk3eknONXjlYQw2NNuM4q8dtky9E5x0uK0j8OWvv2J8dNE
nPaJSpNw1Uo+ps4jIx70MRqhWCi8Re1yDCKq65tcnSNdHcNrfTmAhWtKRQRS
PZOlOBvyc/Flkje9CzxSNs/vCzskzoLmIPJUNlm41jeiIBmb7eWsx/Dj0B1x
DFgezXEpFpDPNj3N+/GKcaffKOuzV52iWNs+zOyen4WGjENjsLkzLPGCKSoU
6GAXXKsBmuA3YWUaULgDvh8X0uWXf63kKYTrsqDnrZKvArzSWWDGuVdjbJc8
6DkJoO0dRBBLN3O4bAWrqw4vOjvB4oqoEkAh5LaPg+sdgLDRYXcf0CKpYIRm
rltMvIGBRbPdh8bTijbQF+tuxUdc2Gzpvlwm8ZVbLVNxMXX3rJL4rIVaZszp
KZipz4gTTeUiHaxYP2xpg7tsjrlRcYASi+rV2hhTV4yoArU23Xe3WB+sDqNH
0l2p9VdgJL9edZAjoi3zsFhTL1bIhsfN3gnIQTZSXesagmAw9y17lrP88BRF
21p08rz9Q561D1d36hc5D+GhPAp9CFdtG06wMXOns8GQUlZQaPaiy9JIyox/
cfb/KZh1gBJfoaxkGDxPRrAWRtGSqEKJk62ekLDZpRNaPW19mlsDewD5c3Lx
LQsTyen3rSeBFMprzS4xVM2nu+Oc4DpjQlRueV3aug5h9fw8bhbEca633hM8
EmJIzdKUHVrlbaPD74S1CH95UXHqabizTQgFPmEFZ4PZiPvjN+mpFxtg1Itf
Gmo5Pjegf42gnbqADdIE56vWW99bi4SeqGQeoQiQzIny7rsTV6deRTxtdq0a
gLBERfBhDmFBvdzfvCD3W3k8Cx43/GPrSlbe7jrQ/T+Z2ozWEyd1FN+JsNHc
pYOLKzzbDoDr6DVARDmgUn0Qw5gdoDkIWAWySGSTlu3Nsv9LC9KrDFJDEIYr
xGeWHRPrl4OUZALJcKJQGfonga5Zf/rg+ZVsgB8XPTLaSkVpzbP/VPm392l7
zsR5f9Y9NW7rUx2armEGZzvpkKfpi1in8aw3r8Iu+k8H8mX8UU3bxvTW6uqO
xmHkbfqJ/WeQndsmONeGGeNu2payHrQ5+uVs3SwrUvQ9QaRcBQUNosWLoQwk
m7NLDXmKspHP5AShaidyVO2//5v2m2Stdbt70U0m2y6wLfbLvpk6wSB8VF0C
wrg0Mg18JOR+iHlYB6L2VBtYFJ1GFBqtc1dyYz/KxaG7T4rxMy/sklzFf/Q3
9jbKGdeL6tI30ZREnsshUyQ0o9GBMXYLV8rhbb4/BihKoK+/grEQglzpUHxo
D/OuVosXv+aU7M7bUWB4k2e47cEb64hmt4Sv9rPMXPui6l6NwY5/x0vaeX2b
GNyXqoVFEEHDB4Z7mGGKgIcxaKkjuHsGH4rscfEdmvokGwuonsLGhkEzYFTu
07xpPy159AqxK8kPHRxWRhRXrzYezQHu90b4xFNoF60zK+h8TTEwcV6Cr71U
5kZPhT5iGrp4BDPWmIJVYds07aHfI3nhxrAMGYHZT1EyQYN9BPZr4dkTEpBp
68BH8Qtqy6BBVOZuPrx9imKpcsPkCdhavlCAgVZ9fN4YvvFi31y8+SHui2Et
clbpA29jiJOmJ+dG4Uz88maxqMfsKNtV4LZIlek5GmGFnall2hk5yqS3eNBO
t9GrZAbZXeuK9TauH2x4NUHHBeZfH1qHtDDbKsNdmhWUHTClQgjnQZxyVdqw
SgcwZFJp66QO8vkXryArdZkjvA2xtPRBuR1998frCxCOioA4p9YmEglTfLiB
DiVMXGziHd6aRnvbcEHKzihgo2m5MelAy0DaR+SLqbNZYoIX63dajTcyhgcN
ws485TDMaSZK//147y/eg4RBQ2tCWU4t3Vtw0pXQzgVNgb5eA83Xz03lLQPV
q6gxVfTiW0dBLeg5uXWFu8xfFkrtHjuhFvKWaIoBXMgpkhxoeFu6+zjgd8yF
17r0y+c2M8qewsz5l74XHngDcwcN3xkRsoK/0qZoHdubqaltLAcqL/s+2wFl
cfdnv/kxSXzE6tzVwZ2F/DVITa8iQFKUHUPk17u/0W1mNKJfWyQNUO5foNQ3
Ud2Y+HKkMng8YOCYVUC1TznxERrtsU+Ov9xCB+wEJKkxnw0Kzm3o2NHJSXIf
pAt9GoTEtSzH3GGobP0t2kQ2+00UefrLLVcXTDR1VZe1wmKRMUXwE3hiLowI
N4dKODDOsyF5NzXLKDWcEYm90K44FtJUst8SJ9BivRGpGpnWZZdQ/AbGHzSZ
8sI6X0LPhQLyvoVIy63z6kR1CH6Z2TPqemJIw0HoF3aP4EbYG1whN9WmfjHO
yJltTBhetNGC6+RaSx9d25oWQGE8eskGH5mlYGfkAlq454U70PnJ8KVC05QX
nstFbZZFSPYjRLZ132M3t9ALfPAfcz2N3TcsO9UAMdOhgP5EScRSROKe+vsd
Fc6YKPFBg/Yh8zepL90pOwjbDLo0U+UDtfiY73wmhBali56pDRIslhYcj6SI
U29eaQqWLIgR2eTLNoVvlf/ozWzojWWBzP6aH3jEJrJMRlbE+eyEPu3ybcEq
XEaH7GmE5U0nV9FjIjZ1msyy31gHRKFlZIyC4G1X5ox+BT5ImJD2GWXK8ms6
BnOQYKO13Jxga5SPXCgD39OH4tbVbcD4xN1r4PCHg28QtRsgfkryuSpSSmz0
0U/yKxl9kksXd20CG17W27SXbnWWvf9/9rZFrhdjbO9oOpa4lZieiEMoivZ9
ZQs9X+8DACMkvYXEJvujxP8uBreuVQb2Bvqpa9WPtVOvzQGiTVcehDDhJiJa
S3Jvu3V3cYphz6JjRqvg6we2Si6tLJAz+uaMRjwErD5aIApLUpq9QkNdWTMo
BCaSwbUS+lZCF2SjYB1pAHX98hGye6fCDD577Ys/2DBjZfwAQyVsYD4z3og+
nKq2y8KpEclr4sTRafqejPKcrHIB+PHgcxIJy9H/l38ydpXA60e/Mb0gOZJt
Omo1J7Hn475KW1HWtqI+4/PwkM3rcVRs38j89Uxjz0UkPgtkYqUr3DHY+/k1
5/a1OVWhYk1Zo9U/oPx3JKAH+IvExUuK0zeSyW/p6OFqM9jdSv5PrCFVCmFd
g/jhFK4m6rIUn/oKVZNTM8nYq3OOe9fvfAZKOQeVVe5ro6Yq3J67sUpjMylE
+KHLfiWJdgEL/UfmCDFOwWi5euQvPH2MHhyGQkvfUQHygkItgyBNfee0uKm9
rKdYKHV++JTZEGUcmpJqSb81YvS7vDGQAO7HGJKSGtuadi/sirzYIAR1/bam
jWqqCnfjkAX77UKNYfd+32SkS1k+VFzMIBO68ug00yR4+Vlx75ibWy8DPUOV
w/R8Zw5T/NKQ0c1EoUu6e/lWKx6VoRuVvEjBsQ1fLen0D9mNpPKvPUeftleQ
8vQG1o8sim3qdwh5E9olgtDTcbSNguEGTb3uC0HT65Ne6aFaRmrIdED9XBtl
nCTXVNl2DeH/L9YzMj8XrbMjkIoVpCMZKBKjmwNvSRFcCaryHej6v5/U1f2D
t6oulwJ5oza7trcXfV6Z9rqsK8ApmQ0/KC5pts0WN5QOUc8ZJY909GsCeNrF
udcnOkdjgtRrj4rui9Kh/mmHvgK/NozenK2rbrgzGZX0GQFiWaE5BlN4lV+g
oRewSYk29Vo2mgPTdsgJOGhak6gTQDLbobqjbv5CIJpSZTG+WkNtn9n+k8Vu
4dQC0SsC6sW5DHRcjXRUI7j+vD/sAg9WsrsjRLbz8i+1IRcacSlrGMNzn8VF
dOyAME8yYFrsTDPYPscFDx0SL8BWUmp+V0CQ+8k9wAAeCSt5Wu0jZR7hUJr3
fZtBSzTBc7earrIQHQQsa1MQzXMSdG5ZTv+pIDDhWFfL9LO952qr+VfSnmPb
rvlKIhXCNHhTUlQs62BSMbiIIAubsRBpHXOtMx0e8hzlngorzedHp9jzgsHW
4hJhHNzN31dwQm+ND3JEbE0ozm40OALYAblTmvWGngJiBSFD9J+2OeuweqTE
hjq21uV8xBhF8ymgxx7KGdczHPOSrB5HjJshYvgg2FDQ7zY65WjaPdygRmGT
5k/SRpSZEu3XKpv05YmaGfWRVvDTCK6iGHFjTWpS/8bL7K/QB9MHLxXHB8hh
sQu5UUGfpi0jvL8VD2/HI5gMl2CYr9B1onTg+6cm5ajUMwuaB19wmcjgN+Me
cG8gykbmgNodJMMMHMW1yHjsJOAXLg3GT4iG4KiIDpYR3iubH70Rqi/+G9on
LoCLs6l4T1oDstUaYMUkMJIvD1j2c9R0U6yPKsAovfbFgksF2gxSJ4NGp+ps
i5n13k0Nurr0N6nouP58mhVCWZryhUmr6m5GzMo9bpeL3XC2skXVPybLtiOK
UE+xDnaqrNgN/D6gmiLSUDRt+70vr8+gKUG8aKTNujiX/MApYvnS5zZ0tb88
XIj3h00kwqqAS40GJPIAQf3qyAHbaxQBiWyskJphe8dQ9/T3Sci8AR3rBOc1
7gkkUP73SxC+12b92dnFOLFHUY+pEYGIaRSS9w07nMt5xdjOK2kfVQgbOOCF
YH/5Yov4+gsvlqyYywDOY3jR52gGGEZFoUg747L+qkj8tVIqUPxxWvRSYr7L
RDSXqiLCSDfBiUc9sxCNWkrBeHRqs+VHhMnYUYeJ8mlP/mg+RdNLCBb9wbN1
IvHY5ztsHaDIXnS1bC980op5PwBBFeb+OPDeeoF6aDmZAAKNPqtzmrUYaRiR
WVhr3tqyUcXEyxxcmAsLCtNUH1ewWtntr6QhG/BcBmpsw2c06E++E0Mp2IoK
ZTCkSUQgFrCDGTcg+W9/CvaAcPYRvqMegxjcBK4kqDVBfoLS3jFmfRe8O1xo
V1iQq2So0B5u48S5BKNIh3L/Ypwty2iQvAs81ptZnn/DImlRydYIiqOH2xFU
kmSNhfKDPGXBTC3wTqe2I8No0HflAz77yktGIhaYDkel7IgROIEEcuIDBjQB
VbHdD7Q7/CrD+bz1+u8XIEmEAIpgFkBxaa/k1aVjuWLUeXraXktZOlhGedzN
o6cbnk4GqqmNO+4zhgSdvz9sI5GidmHBtPwJDrg8XzhfORoup/ybAeSnQr2Z
5hlY2s7UZe00Ndi4zHBMyuKhMdbPJ9Zr+rkaAhgr4yFiKqgEoHczR2tYABL+
pUIUO2b9ctLkuDOofunvYPyFPbINMPnE5ZBKk6xMG8EyTlpasnZWK1+d68ah
oJb4dnSreGaNYZH3J8KtLD4pgYN+vNWaAtn0w80UPyZCaz/ToDFaFkzuV362
yuQtPmfCdwlOHVxXg7O3BaADPAd4BYhfzZX5RBFYnxiTqFT9ccb+fUUGbCPz
w6vXnduKqomPvQ+6NSlBvLoYy3x9ytlzz9D5k/LRzHgcVkVb880gXdKz7bQp
PYWtHSVLsbp5EoGxFC4scqgb0tnUB2W8av7pU3DA9sZ6ungw3xGx+eyNe3yF
/uHCTL1WtcKOcjQLW2WkRP/lurlMEYCpQzz7h+oAI+ydNjDFQmBqhNNB6AZr
QxrGOTAT/2iEh8hWWmEjRBYpTGg2ZBbl2sBKHcbjh2/g7FYR0iXkxy+/suu9
i7cDpzwxnFiy6KH7ZtS7AL+KQzkyT/eG7RUkcxCQPGZgh2iqLfI/ctRNK5ji
J2Tn03mXgVaKZPztWhptRHkFUwLOKGS+wI+cYgyURDLToRyKUOrEIEzVTQCf
XbQH5x7x3o/LnAPqiY2/8gXRDAgPFDIR9BSsBY+b55IAD8yXAogWA6lAmEgy
Y7zIE+mii9ah+uefBJl2af/yjnKlJUbMoEwJb+uhEQzqyTvM/TdN+8dN++yR
BSpcz4XhXGMg7VG7Jmte2gcqHZlLSnGbVcS2mUUUIo7OE12N1Hlqa3MfnC46
86D6dM8EkOm3/aunSmkpORrdOkMhJheice5JRkuuDw6P9yvsXpFAZJ0zCKpY
4kW74q4hFwxKfvhRyrXNjTCetXPLwNfH3mqEWS7AJ0IEhiFx8sFisyVjDNTY
m14wQNHa83zP6P9xI+zb//HSVJcXejjoO/GYVwu77KG9ZIOMIUFOjNWPiY+P
YRS1R2AFgpsU0kDvGg47k31TuEm/TpPEaAkWEJdoXkr+U+7/xebkhGFlSLhc
YRqGID3rCgPAdjZ3fNHks5Rxvpwo7r5ni8PBXaacBWUgBS3pfj+PuVxPD6me
UHWQ6VyjABYuVQiN+FeM7VQCMqM1bE2yn+yZXE02YoYN/jJGLOfd2VyucH8z
8ezpMgw4pLqt+dNfiUdCcmp4JTGOJhhD3H9JrAcrTjJqi4fp4JdF87GaEV4D
wlr8o9T65NlvSIEzSzADzI5XUG9f8ejhUwAqI59N3Mw5kmGBR3WJ/vOrnLtz
w4YJozNhM8cImL6/ZFfXXXr6pP2GpzkZqz03DVLr+ftl0KZP6MVPV5WHlhPp
8DnMuRZoSLhGNaK9L+7iN440psekWLk0O38YgQbVeg1m87t2vx5FpB8TQvGr
kcaXuGZWlmlyRlgAW4eVk9Di3jYIDohbpRPnnQa+q3dkBTo0es/Pe18hnpMg
qguD/3k01w6cJOvkDp4brgqxrtuOHFkzWZ/eWyCpZZBgJTyp2JFttwZi0rV2
RWW+N8DmENtpE+5Azva3l14WbhVyMOOy6OCHPtOw+he/xRV3hJlSgMWFQ2qj
lmP9BA3zzAPeg8QORGBvCDb7YEGkpMxRNMgJDtbzQ6OYPib3eSDIB3BYW18f
ywWsuCRF5ppGhq1fwrGYCy0iM8QQAvausNx6eWrWB6uxGFmnWy33ShBpblYu
i4AXt29DPDLHndhU3w9FsnA7E6jBZ7zbK5aUdBOaFdKSwIgmdRPdz/1MsBIV
gN8WMdDZVfR8kyYjE2vHU5i7BFAIyI8BH6Qa9cfFj8R1V1cyJ+rsJPsWVX2z
tUJaOQHbXAZO4VYDT7IyWBvrsudsxX6MbaVMIYNXoA8cbgH158Z5HLjD9Ojs
V1aRqt9qZSX3s5dufWpPSzqZheLKLOGYswCob9BEWLjcLLI/DkozXqpaW+ZW
3dLg6drBarGE6TeanakA/ofnaQtB46egx0jD0+GndzoW/zZ+KMr8wGxqCLMa
cmIsQaf+4iDqyHHq3p/KwR/sb/6NhVW70y2cjwAG+cUyRxPjjeY1zaeq1htl
sDySoBxMxaZfR7qIqYlSvFXjINxSmX+KYglEu+N4dgBKHempm3G7QPGmKFR/
B0Mz1U7lXxa625QApcf5D95ilNrJ0NCdghcaIaCHf0Ipw7mJLPmS3jiY0bXa
ytorVP8oRBSwFdbhLXm107gY9+LIkLEpeKXJrMZ2uiVCOK+TTE2yX12HjMEx
uU5tKw5yKCMIMwSuWzVWrYvZ6y14pcYwVOEFdyLtIPcPja9wIF0jIfNOiAQN
XJb4M0NAFaTcPagC3sSh58WHwsnGYtG7W3gtgUObLavKd6iGHjT6cn4RuOjw
d/N0dagYfDJaRhftZ+sgWb0/IDHuHbSQInceVq2qVE+K4vCdncX7nTMTTpJL
amXn9cx3WoB0gLEXF47CPUWgwDCQlqwCw2vb8PaH73g7kxcmlDMqU7qgrYjr
8qw6Ox72dXl1ddWMhU2fHI8Yk3JfS0Mk2GcMCOiS8uFyRmrdOVQMZIrC1oBI
nAoy3genV9yQ9ew8UU7hy7+b/MFDh9Mx+XhUGgqIYLm7PH3I6BreseAHEig/
PRV9Cyu0ReZvMsXpdvyGeDImJobbATxpIkRA8Q83aLjS5Le65RMA9kXh2aqV
vKT2Y0fAVRtZBPDdkwVB2swciFEobMxtVM3cn9pW7qG+dMMlEA2H2VwVKbaW
84KxWMZXUEPPlrSha7jLQ15SEL6UCYm7rhV+kRoU6Xp+OSIOgrEut6cWYY3U
cuuhY/Zzw+CxkFFclYk9e9hbRMDrIR2fuqFTWrAkbJ/0vDLk0ZXKeSMmfAXO
e7FO4MTroUVaz5K/Mkw0l5y+FUqUX+QirSR4fwUIXh2ngcXziDHC7kvJ/Haz
DtpnamuwuX1Hr89i9NJUgtseihyK4W0MPLYl6Bx25/PBlydjHW3T8dbn1dOf
k9HReTmxxM7rhxy2GHK3Zi4CIQtmc6fi19ieNON3psWBGgD4LdD0NuHexWSs
JFx3CXS66EthI2gO++Jr5kRjLfuhsa2Lvxk+iG/DQE3CCJjcJdasa6LyBXSn
9nO3WJb9yLH+VwQrleseiyKZlG9cqcewQXeU24+vVeB6SuXXcqtazMUDB+cm
gAkQo5cncsB4SXgVzYgozHHds9k7Uh5y88u5aeO1wWlmLe5M2HmARZlxtDPF
cDt1tYAtccO0WBX71yIjufFRLISiw3mB/hxU5c212zA0gr6BicsAZZi/mlGM
hvr0P2BeFsoW19dgt7B5FI3G8LDAUB9RbHyOkI4Q6rVj8xZ04vh+aUd2xoV9
+HFbQHwBwKs9VYPM+ptTvpisoSu5iOwShCn5U8hA8VsBTRkS3zxMXpryhdAy
H0Mo3lYRQQz7y+0iirwZ3wwufK3VEu0QX9co4dEiVUnX+Omvwtdqp9jPqhqO
COnxspkbkHKsLWkRJWKeJJ1ZFoUn4/cHEZdSWiGI7WQnFAb64tkg5jVKfRqt
UUbjv3x2c22NL5+LgR91ve1rIHqPUvZmZKrRjlfiMSmrZ7f+YWH9yZjhPAiT
6SFJ0OHGVZBcnrDN1/zYRn8GZk2CSbF6JPiXfXKcsdh+otm7q7zX/e2LgMdR
H1hB8Yme8mbpOtFotxPrXh8gojQx2bID3pK78wxRHE+dxodJlWcmocP29RAU
FPBbQBY9feYnRdVb4VT5i4IAGN39ljlBFeCsL84AZF43Jmys0W4AtJ2ZbpsN
IXqkZSqh92TXLmBk92kY3zNVPT/zn4oV1PIKdxU4ciZqrfstpKdyK0yi7nvZ
Nf0e+7tdD8dajwV/7mk6C7jvqTnYxYTTEPwXLildJoXrlW7waBkhIquHmh9e
r/xFY6sp6QT19ZD8okm1niUc3NDqFtdzfXgCmJh+c5kgu5B7ql3n8zWIkUYh
ApOIEZPuTgCinorjWc16Iki5SjTRIaDs1vKoXFsUqrOaeqACxioushTpZGrS
pYIDWehuPO+LoiJ4ZNQrkrZ6DVc/kZ36Xkp+LWnGAZiN5zOD0rcbdVv69Q/N
HnY03b/0Ixn1MQG2jH8shKOIck4rYE2q3CKD+EQw8Y1DzI51LR9nSwSdqnC0
ZGEPhMH0lQmwgN8uXCDC1EsZy1Ej/fdbgce/KIHp59TanH9Qep4rncU4p5GX
urD/VasgmFiy5diILWD41z0kCUSwtMOPAkJZ5n77/PN1Hj7cu94HvgyqnqQf
wt1+3a+Dw783LiHgkjguY1vv7X7DY7F1aYkiObQgQGj9bf6NgQGsPG4DbSgL
W8np39Xg/DfwbImDeDncjD5LPkGbkHTSJiWzwH9kAQsEiypcLU1K/wMoPh1b
4hit6DU2f3p3jJEN01AZfjbPG0EjT5bPKFkWv4cV3G38gnVG6UGBwI6cuFov
Q/UFUZleXaGkZcGyY2bagYTK/l2IRO/M0w4l6BSNTnwqZj7qzKfEfX5VNcBL
EtvYq3NCRixxIRjrlR87HmDUEOy+J6LNdjddm0wNxupdqkPUEljltkrlwgqK
jHdbxPs7tspg7XrEnDbDomn90NThKZb8yyQvXILEg6Hb+pjgAsmiuiPzNSwk
Yhi5gzxopz+ovt7NkGrRjp0w4PKvOIt3coL3jIsMsKy/Ab2ks3HObhNOid1p
5AkXWEql+xkvNFhpCJMKAggJNiEfWbY+aN5risecIs6/HH+O0lN4xLU3G5e8
gjVZjQ2jMowpMtdXLEopvBzJJ4VaOS2Ue7xow3xb0kvkW6358+8DSNBsZzbP
iHkeX9w09XjldSAoiIOlI+k3JlwgSICIOJ7fVTVFrQOrxmz9qqMyQVMC6W0l
GNBUPckKh6cW9SMfFf2drAlgU93s12tlrpl3iyiV7ddNvOJgirhVZ15sHzRc
dj8Tzoe76JnatrL9rmSTuovja5XcWe5rOlgeN+7uPBqvI7UhxOnpxja2j9XA
LnY4NntgGyiv6s4v5ozkaKck223ZXb2iRrz0bUpgVPFHgIHYMIJG4J/OGY+a
6C9YNa9JIi8FKqyuhCF6CFxQwYIuAPoUFbCau7v+fpAajJvuSTImiMOxZWkn
8/ZGLuCM4ZwybOA4llDoEs0q/qyvWyDb39H56D3s7wTURPhK5rXZMxNCYL4P
Vs+354irXEAzyypqWqL/G+4Dh6lSYwU+XsPP4erSDMtUR4ucXoEt7zcvAk9B
AlSSrxjs05LNBn9SoT5a6Nh8b28xZZbSZtr91/w7MTdlPJJn9UtFV8L+bfV9
W7K8JJBWzAuPfOKnHlgnKbSieLIVbOg6u/IT+PwOUmJT3KUeYtEmXrOdNhjy
HREJFaekqczgqtguGfMR+S5tthjge019NEpUBcsar7h71MiaNzayL7sonYGe
XL4AKzZTVOv5m7hfSz9BaYzreT2w1VUKbvANDZLuwHwgAisTaHo/Ml3ePDVe
jPEB5PcAc7mfTFG1K1282K5ygg6i+sQZpbiG4bFM/Jdj5i1+u/hs8KE/LLrM
qNrFd74FLDhWjkez5TP7Giw0kwdO4j0vG4tZCHLiRolQ3ZJ8Akiqj0yDeU7w
+ydJ3Ws73PfhALKMybUUrycKE6eErKE8Fz/GOANr06Tj7FnO7aiWjFwjkCsm
oGWDAHcBn6/HriZF2HpWQDR/McjehOMoL468YwiJeYIHPzmkB/z7YRu6g9so
Q8sNE9SM/a5CL7Qsc0Ly4A2FJ3iD/5Y8ImzWKMehWrt89hApSysbO5K4oMhS
6S7NaNDHH4WXzcf+3gkI1rCLd6/o77RNjeDR50JdwgfQVNfcxcCeo/4mzC4X
HIcJ+qV+O6G/9ReUMA81PcO3fxQqA4s2pG3PInyUgRK2tPup3p4BuLgxkbwy
7Gq9GqS5EhUEWcgx2Uhp6Cuz1ymYaxrOdIhx8wo8BQgPDjFa9/1PlCN2hWVs
buC/O4yj+CNsiR0RC7JDbyGuedy7LGTpc6bnd7AOUkaPt23TJYBYVw692c7V
0TrxpUaSUrO0TNOf7K4ZrYbjwrUbF/xdwZUdmSsUpvk8huJOewRcdxwKDUav
sNuRgjqLHny+QNwoBxl2M2exSieEvfbewDZvV1AlO+Hy46q1oVvQYAxIwChj
Sw6d8wQAW1K73+YKpHADncViz4sKABi4F2mZWskm+JBNreaxxkuNjcaSHzl0
FfylHPTxmcvXC0b3oIwzi8pRAapN68xVaR9cXyW8zc1xh2lnepP4hGJY2Tvg
SaSu4LXYj27MB31eh3amIBS+Z5djJ/e/ZXvniHt6eCPVaKrYoIaZCI7JZ4Zm
JKh3OOmjQbcOaG4WHRKqyYaQnQU3k78MTmSnedThND4mvqOIBd9K1GRC5R7e
Ds796l0/QEblJhBZzgK+yaSlTglvmfPCO4TGOOWoa+roM544hCkZfaG+nTO/
UjZ//HECfP9V4PHR/yxrQ+1NBvBDGHmd4hg5SL/9BeBrLrL94Ka7VKLHcvgW
qaXfrPM4cmyRL7sYxW3WOrzGA5yLZ7g8p2ZfbeSRTZ3ifVvia43C2GRlqLKj
UROMdtWEvh3QBRIU477TdWmWSN3kq6XPUUqCjrZm0wyrKZ6OoTU4WvXK0DnK
GxmwE2ZlRKTam5hOSKZIVM5GzghV9jKdBYstA6X+g/xaa7KC882nXcSGsuoz
I79gjpu/SZqlGCKzu6RHgWc2EbvfsVFmOqsQVuWG3afxcmKQP5NihyNjCbVy
qGu5mNtwQmKXG0S0D7I49SJAL578gKeE7vzyg5oBrFXDM15aaa6dyXRZquGs
1qbi6nxYSuIpJVvI4dAzAy35QN0zLaD5CLFcjs4U5IXZSGE7VgtI9/ZD1xIV
S1VnXpHefPGxZgfo1R1xuKwKyS5nrADD38htV9UeyCKsfSZnHPU70FnHqJDy
Osw/9RHjdxqvC6o09v38+0EIkjsm917iX8FFxD/9+aXdfPyl52a83ZTtmUqT
xH5v/GF/bqprmd4lPInDuzXKoqTaant15pYx3XFq2Z3Ket0Efziu+zmcQ4yY
/1RPRSG1meHrqomnc/LljhHGjxIR3AuCwbetjr0ctvj6jFZPJcs/SRZ6JxBb
kUNMNzHdeI5InkgOszb2S2NDHT/478/mZHnYj/WdPv6oMZvEIX1FvqESx7+h
/1fSOAyNc+7gKzjLb+xjSnSlq5ligkbShu2ZBYfloUATMtumCuGhMeppHB10
xMG4/BLl4RpGlMjrhb49pBEurUb0fRWgJnLuYmTu2QRN1Eph/5gjorCrTu7/
PUJo96LCsJhk371WsdVuDB364lMu4/917S7cmkQ6lqjz5TCB96LdpdphaIMS
Uk5yTQ85AHPxMgHEb8gzK/ComKc8ptyg/Dmst0zTYXNFvtqUsGU3R3oP22ck
tyofOuJC0u/KU09hA8XOe+jan4Fx18Hd+aW7Z3U75bvx10YpNehdyiaoweGP
dUOrqm7CS/4yK1vYkjC599flL5DLE/DENwIlxgAK4vd29UcbxsQfeBtiTx3l
UeThhjcxnbAGs6CAdWojglHeDJLmgCcOGxTarJpuMyjANM9eeWjkN3xgopEh
mukL1cKS4yVYSGTHDwvWeEPTsApMPnX24g7VhswiFQcpcgicLueFUIc29OoM
NclLlLbD/u/CzEWGp9Ir6fmPXV1dSph9sIjPSJM63gzJhDKKdrlitkEHMeYF
DzkUIPjZRC/iuwebgSMkb5+SrGtKryOVBpQEHs4Fe3KshkUaces4UnTInKtx
MhcOC+cegXafd07CEVoR/WxD2ycUnrlL2UNP4OefFswY53L8ttl/JyHtu53G
rJUJO3LStcDHtVNj/Tmh/83KEpD6e7WR78umfwx3tnDMhlorKdXrTr2v+0Gw
MId/4wAPgF8NbJ31OZEzFO5XkvjavGQGx5Rell51uNJCGtAr0YYBbeIqckZ3
nlT5dQFdjLEDdz6RpV9eO3Ga/xawVJUqtaL0wppg1HNF/F8GhXFAPp6Hcroy
wXvfe370NiSJ5zQZxmSwKAzVf5DM8WQ2Gb4lOXvqsUUY6s7b6iX+JwGLekZ6
LoSQy8BhekJfZiyCVk8vLbf68xwQfSJeMDG5jpdMhSRb8sEOoKrbuA3Zn2aM
/Z17IjQFV4bOYUx/FeagIZvUXxWUCSBf+/wC7W0HxCyH3Ly0xma+sGT0fRHj
LKsMeKFqPnBzRJ6k4qaC6xeuq/aJTSLy62uxROuwI23HKM7C9DuL8MAnTDij
G6mD1+1NbZBXJ6eMDOrc+E7jufGNBcFf/Fix9jjh6vuH54BgMzzglbfx1/rk
jIrZojsmR5wGNw2Dsc92y6aoRpXnLQeo1Pp3w+iNHu8FrJJsZueJEO8qaAIM
zllTKaKJajq62OSxc8hZXnGbBFTqA4UOywrOP9JGDMTuVGiRYLIriAfgADjf
VrVTzD51cc0msnF1qqGcNsPWpj5cMDQrlDqh8iFHfsaNuSZsLFjsAjJ6sedP
OcTyvN9hH/yXrCUuQI89WfKREuYdg3hNdb0GaDIg72otMKtrVQBRvpekTiG7
hTEljdnxUE2kwiwteyeqK7ct64TjFvvQRzHYtgGeK9oBOdqSbsI4xJ0n3ZUh
6PUMC5iauevmq0o5m+jCuf5wYaDxkxzT19hS6FIwmVOL+cN7z0eKM9usojg4
V5DvNYI5z9RcwlkfrZeB0ar0iDr5LJGHdqHSs7jD87heiAdogC7rifXd38aT
V1Hap4uegnLDHFs7vqE8cd4OEufZdfnnGHbYRnaPav3HyGfZSmje6JhLmtRH
x6sjMCJefwbED96IJ1ALBTpi5Oz5F95zvMhKdxQsDL68kinJtSu/IYazvKaS
DggCwomBzOh5AsWOVL1oUl8jJHDcghH/e5K1ySNuwHQ1oTcZyDu7PsYj3A8t
KVoHb7njJDvJlfjvY9GqB5OK2ZWNS0xWtsMjPFtKRr96xBIhFOQorb6Co9QJ
4ZYM5cdBd9sC02GF31wmu0pCZNFfJV2zJlx/DrXgZTTQlMDb/yXNCMp41m+d
K9GT0QN002SiHfV/b7Dc2/GQjBRQ7XhZwhd2sY4imV5xWIqQMvlD4WEAGjhg
nxAsd8Vouahh500LE3HXcBKjlJPeAYl9G1NVn7nDNmcZL7r2HTOkmw7cZDhI
BTVZguZoQDgX9ToeT7ghFmEvPGBL72wzprYeNjHLX/SUkVwjTEu20CiepN3Z
iwBYecYXMGaINiyGLkl0/nf4kaHr/2Nf9OX2t5FbyRcBU+U0PjTyfch/lKR7
EiEx7Q/5T7GHfQvZvkvMA3IToFA6YxVLI5H32rWPri+HQnelrl0NOuOCDPpD
g+Kc/ZMTktZ6CmPd+okDr8Ucp8Wxm3bm6YDhllyHmZPoA9WX1/oyM42DGUjL
Lzjot0eTvg80pu3oatS+Pldo8XVDjSiH8enXaPnKAwKDFPO/+P9WpK7eILVU
+J03TXnyP/aI7Q5xpvLxKCnhVvay5EVbStdJvJgHUY2+QrxR2uh+eYtBb3kD
NKMVJ/ggrqthC/GIsPDUHOSmpayymi34S5atSDv3MiV8rs0hzV3xFM7ifmwj
3IrRMx0h7fTP3T2qhCeTbIBur5Fm1nZCx5pZ2sCMZqIv07UXuf6f9EFbslwy
oaiTAan8pjORbxI1ZVKLyUcPUWo71jV0xNXnRFrHqK5TTVcgnTL3j/PlKeI0
MHfrHtmQqSZXCVKEfRdPPS0HorcxTpmJMbhiizQv46DA7E5aZ9VFM8A9IgyB
DoXS/VsMd9WJPzkdepVWM1kT5GSnoyZQm16gChtkfr1URX5qiMtgEbV0cetQ
VTSW7VJS3Ci4aUahXVM5uG2jBr5KOCgzPE6R5+ng8w/viPX9fuYQLSJ62MxQ
Ms7ZyPpT5CN/wqkPQwCylixlVgQKUTLzMwjOI7EqSW7Fbsa8YqqCOyphuW/t
XeC4TZELdzL+2sc4aPNK+7Qg2KfRq1iIkS/JcO00yriQ30kmX8nixHabUMc7
oM3+U9pIACVYwSuXqvV+09+h1cRtFIciVsip2EZmRb0/BU2jQ3rW8raBDQRc
CG3+Pw2Dd6TfNhG/lwvyCC8D1fPFTyLtxoh3zwn68OWjG1hxjmZIkp80CZPj
VtS7O+I6KmhAlylFq+oJZVH8sXO/ut2rBj7ce7BpYJIjmx0h7RQB3zhobQIe
HDgaiynNFUunL2CrJfwq+7BBkLz3bzMZSuZDoFXV4MNy3VRPFkE5STUZZYb3
eRNIR9BIls8DJWj7XNbKNlKyfPS+2m8KrwTHuqBVWwEQW0IoFvjXWU5yIdqK
3uAWRz6PWc6NVk5PU5HOYXf/2r9kfNuc+gkbMl2mLuVonkG47tPpf+Mynqhv
bPlR/WlMGLCE5THfy9GBhCafSUCM6GU0SQUltGG7mMgC/7crBqRPmYAe2We+
1p3LCta1xmK2ElZeb26rRBlZ0E48jJpplUkuCReZFiGQJ9SGZa0ACr4l38QK
b3r7oQYO7z4/qjECLA7Qd0yn33cwTePUqcYhSuMzIGLSoVaeg9DhRIwfv6n+
Ry05YrgMsno9cyeY+DKEWUHf637fhfFFd/wjFQHtuXzLjILh8P14sP6fDxA1
apzCZQIArMrcEE+qnRW9q+s3YDkun9TsMygTOAjcoGml5a96y8nKLfazuCp2
7yc1fNiS5yTRiQvYPUpbtE84L/SrC50V1j3P+Wj3YQ1nUV2yISZsBBBGaKkw
0QTT1PILSITFUAHobi5DIgvdJM2StUyPPo/BZDTgoU4GfkxBC1PERPPpZSEa
eqnUvPO+SMGP+svox7dhhfWu6XEqc5T1NMHcdCpbuPch53amkGFUkGulvU6K
Pjamg2J1bjxD08Icbw25C3/dyltHxLj5SpyPDyY1MkQohIe8B+Fyuo7LndC0
Wht+dfN90ISTN1F49IOnXiaHNtv4z+MDy9BRDxyOQwlm94J8vPgWmG1d0qDq
PDyyI58J7Ar/a0LBHV8RLLNI/7+Gl7GwnwbmiPSEbBCOQThU5ff3ULAW6G5h
Evkgxby5NRImaS0Pt6qpq1ZoTWITTBrlGUXulLZy3EcmW56X6Nba4eWIbZVM
hIlMuwctaiuiBO4EUC5NkZskrRsM75+U9MNiGIh9Kumrzw2BeXwdqtT3Bgcu
xzPXU/SAJoGZeiR9iUslVj2ONcGUhfw92xeFirYrs37heFZeOKIhz5vu7yAf
bSHkdXeg9MeYxadQnyJb50XkV9a1QcVnoSgNxmVrbQLp/x6ocbk6lJgTonQ5
ZUwZ/gOQhywpLQG3gMQLsV67LFQo8rZAMulE93jvBKJ13JyY3CidHiTnkdCE
tyP0JBqT6IL2FHre8KgAzjjvMfMnQIvZvuDfFJw2CO7NnZAgiHyzQn/6maBw
TOeYillab9HryyCipGZzjfqFrYykoE5eAGVfaJCi3eBLh6A7h01Yglx3dcm5
DCFuMukq1MUGFR9PGBR0/kSC3s9bxG12xzDRQd8cVwsGbiCTbaAifN/8QDh5
icp/THIDOj2kn83y9gEi/jhLiOcC8rjKibf8Z84cE7jo6vSHmStdCAh5Qzeq
Y+RlpCnNJYoAZmk3VNIEV5kzZgvLaKqI7EMDHrjVXb6+CnG2OU3ESaQYRmD1
jB7KCvEIQg9vmSZGne9URcKdjXDwUjALYxSJmx3/gBDjlrLWn0s5JA1nUHJF
zd3u2zKytRZaNkYZ/A15bcnSd0VGC1mkvQgbh3mmneeKLTXS2zF7CU7Df0RP
YYwDhpfSSWH+LLlu0X/GsVbrscxJkHXE1a9C6HRciH1wP/D6VO7WC+s1TEZ0
K2KsCjWPvy5EbeBG2sXOB5yeaX2QiHsoB5CITx+SyrwWGPhCB+QzryNG5Muj
HSL8gWjHCjRDje5oOSMzXhM5Q2KmvjwregTdhTgRxOnWxEzlk/4Elq5y5vO0
jlUbUreDtWOvSlmrQIjECW7mgzJEICpfClniRlT/Ammpc6KWCkg2XgoFqhrX
DmbModiUUOchXmeLKHNVtekv8w95PAxVUnI89G73iCbutV8fibNRqnIvC/l2
sZMBZu0I0G9TJ78YCXToH9pD5COcFHqxs8fsMsZYNx1bOWx8nrHQp4gXrUYG
WK8/KdBtsprc3eMO/kH5t7c5AX3080gKQ6mtqb0V36H++bqotWij/XUirzJ2
WCg6KyYdG5JX430160usaFH5DaFMZqS1MricWpVkQpMGqNxfnYnxPc/qf70k
1IMRVu1FInowo0HUBL/moruLvAGoc1ABxdpvDAUjyfHyE1mO1GSS7I9wtWOV
clKsWZ0FKJ+MN6RZTsNCQ7V+jd8lNQK6rATEA3SQ8nydS2q63BHABWYT0F/w
dCdTNqLXqBEuc0fSEix3WFOdf65sEnghlan/Kccv2OJMQHJ5DaZiarAnQMcU
yY/bohVp6G+0NYOFu25QOOqaUY7xMWz+WDj+xtm46kKwwSD+C7/wAuAdF7Q4
Tw186ECulpMATdPWvnpeCs0Z/uDyDC7oHN7F02obQRL58TmHY0f6W4q9Gt0C
vNgXYKcRvzuNuo0r+cuaANi8pGqKtxXRIisPZ6t2KDuyAo+kND/oMZlTHKiP
wz8l7Vgcbqs1GxyOvQk6dsIWDeJx7wKA4RS98YOSz2T9BxZj0WjP+3yP7KZG
01qmoNLycsjwakntr3EltdfrqhH5Ha3p1sZN6l8S5MvQ07ohz8Vrk+BVPUhL
Jh5iiOtOmde5SUNE9MHAKYd3nVcA1DsekIgcCfnOr337JYAhFswsYFXHQRvx
umVcjAuopmtHYAZMUv2/KoXnysr6Se433jYb3jeaGkFLj9Wlkcf9PTV+ACIH
Ou9myOBYxL8Vl7HTHF2Kq7WHa9tv6Q0knU0OPPnAvFE8A9cdtmxwqDZ28yH9
+WBkc9lg5PohEJNbRz3Mkr7ViSWawiQUEuOrZDPzD2TLNmjN8j87anyT7Hmb
Hgvn45XTKV3TU2HJDQbqIibItvMJ7VL7jG68fS5HhFwLPcJNupg/l7DbIAf+
en2idO7ulb4zrNrv1Ri8Gh20B1frSbQDh5PmOSshcCqMiITpBYsPj61bxNQa
8YyCnAVWYqzs9fJZ2HqRpiJIqNfXJpm8qrrioMVe99odkY7xHo/Vabm+7Lon
DcSv/Rg+ZKzOkXmrfLjrGOqCz4Sf5oTm6GGl+jfl+12J6a7IN35eu77mayBd
ZQsNGyWa/G5IvybWj8MHiCWhyTCUWlJ/CpCrs0XrR69w6w83x/87qjHoHRNX
7Ez04KJh4z8GcsPPHYUHGZMLei6AfXhYGmdaeZnmI1gY2qgydynlyuE60a1/
9rt/mRyWMq1yRw8zOme7TJCRJz6TJLC0CRmjcsDzfzeDd0cYST47E+idp7X9
dDwj09myPVAtjJv9c4cPGbe6W0vFAgNyODeGsnrEHsgi3By3RD9a7RJsO19s
saXN876SGVk6VueQ/IsdNggqn1YtnhkV23P2m/JNNZH8qHwYExtwQLTijHSN
AeL2DNApsYexbOi9fsxm6L+hr+5IDDsEKjWa7NzdHspiiXiVrt1nXbTuk5JH
qzjph/1a2Q5LAcp33kelnTjKdiAHcG+Pxo+finN6APv+rdFNnLn6XWyoalWl
CPdmU+26mNzwGAGcAdJ5a7kgsg9cjfLWX5bdGVPmcJHpocR/2aDVOzray+eo
Hnujl19F/AFBn+Nj68mL+zwV8d14OZQYc9MFy1h7wXFELWlYODFNpR/zjhlb
whGrelEWLpAVTRmsyxZWjWyJ++bw6kcIB1TyTczIA1pA+3Rjrvk+jcXIKJkd
ELSa/xNTgoQRy92Ccs/7wztFc8P8AI5iK3JGXBPbXeqpqTxGTIl2AHzJOTKl
EvOTKFmU9/J4xnnesEoM4Yj49N1y2DO5cKoXKQXG281ATEg2ZYSflzYYT3Y8
Eux5LBBDGcx0TTL9BnRae6j1zZSHtwq5IqCxpCqjhLfiFEvZQiRnbycRmn+D
G7qO2RBP7gXdI2X+OR/Vt9c2FUK7GdvZpzWcGo5VZGeKpDctkzzoFePnjzFc
vdFkWkQCHwewrdawDS7gNtG/JbeIkhgZlVPD6NTVsDxzHbwSIGT2j4RIO+3K
DOUB5LIViFpBoCx5gyjTCgwLH5VIJBuBjGWUGYKWpPy79BKZoPJJSbvN9wwj
TKPZjguN+myyjGCLk+BBrSqFkaY7gyIw9BP/QTqP0y8qlE8d7SZUjzdwsdwn
ak0Fg52tQivzTdrO9nesCY6ZqNSLgL/ZTAnw5xKp/GQbU/0CifEdaKNv02z2
Tk681t84fe6Bwvq1yKZ7L19XV+3GHzq6aLo2i+zxzMAjRxRxvTk2C+YprpEV
zjvADAYkr/I1CaFUpwgwhH8I3PQkcHIb2USOhOuGGzp5BF8s+6t8fNYFUQ1f
yvtZ+OUTtWM9bHIGWHXjQG0unw4G0pylhDlMs6sNxYE2Qy3cC5BqLQ4CHiUV
+8LuLqz+jBnQ4Vj8GeYj7o+c4Jz1W2/uxtWpSwxEh0kvPdHWeqL2zQjT5NQv
Q2YN1csT3ml4Bec70TLANx7CEpeFLbURo3JnvxOw8fjUnB8y8cq2kheYkZC4
9AIzXjiSomQjAFRmSkw8HhG7p/l5AlFcoxoz/bfBGGxtQhlcgpLsImYnpx2z
n6kuFLhzZ4dRxirKcfHdWwMgs8zBZ/KjvbklLDDNyzEDtBU/oN0UpD/XjSwy
kZXjjDbG5C9Wmd/J1VbGyeAikjgrXcubcw/iznFWeA1TiRiAyGCBmL+oLXc1
IJVMKBj3QfEBkioKdDct8Xbwr5321l7U3+1FrnQDbBpAg5QHjT8Jh2gfN+Pw
dU3QEAqfSxa8Qt+8MDL7TdeFs4Kz6jOaX8oCDDEVe5dH3wS0UGIwQp1FNp+i
PFODP+nztkHp6NI4jmO7UwfW4ML9J5QVx9twZsLbeeaCkZAgcMLGWRzSZWGA
zpBI8eGtxFkz1s0s7LxxgfzM3TRMxbXJISWB+kbE91I6eMShGVoWwQGD5/Lx
XME0zYyjg6SMeo5vZwMGjMZ4y2PCKiY8dUK8AhgYkeRJ469X7df4G1GOJh9f
rQ+GqKLbIjUZAxTVWoSdiEo3iLH915oIb5Gnbn41/iZh7xFZMRZJKdSCc9z0
iWiuD4RsrR0j3+dsiDGKUifzRudD5auZBDPgSotAgdhQmRijlKorcsg8w7w9
AK+Enn9PDafm9qNe4cIzmB3ViUtaTp/vvhIQmRIh9IHlHo6kx2O9AxYPv/ac
Onc2I1JvQ9jyC3jVs9zqoR9c6/oQfET2FbW2c75EnffLLg9LBP0vKp9wDRZo
DOBDj7hyrskP7YK+R/q2mNKI5lUafbeyxvY2Zxtvlif0v6bJsp+JXKMlRo04
qwop2adPchzmqHDzrCrhTw9NZaQCJHFyb41iDYV2f5oj9uAHYrd9mOEAyQb2
FkPgURlFuA98VJxlxz7JJOfMO13zeUsXXJVqnALPDNHh2HFYAeOADlsP5pM5
x+pJKAHbuvcQdIJmYrpAli5aS2kZz5KIkaXYR7HSrkRYNrPYvuWsgJMXMAcV
AzWTtItSiJk/UgKvJ3D8TwX1x+uHfXtqlUp7WrwppXuFC/mxB9Wwj3QYL+66
xZr2dPaSSbX65Dglgv/fpuTcSNHHjSvpSDZ+ZOV5ML6227ltu5cu4dhJ5dGD
/1uIAfIhAzdyJsVtWxu0PCpM2GJIrs+rvcneQBwFsBEFD7H5qFlG5at9IuT+
u2wNgdSfJ0wYp0JYnnQ6/LeqfEgNv+3QzOQ9hVnMZywWo7flfjF1Fv5dl1r9
UCEmSeuBelJO81qTnS8/mOLwMCqhaQ1c9XobEftTmXkj11sLaPV9pkRM+DKp
WU+X4s+dY/32VCskLp9OSlm/au7GtDpKOrpkR1oRYi3J4oYJbocO7h3CcIFz
hGYJ5XTRQSoedtJHiTMHn6rU1AMAVDhTxVmpt+0p5tF5CIhFR5TVUuhSuTS4
LBI5u49YchVxAYcf3AVr/sl9/zyxGxBew0uYSZrek8uiDcwSg94ag9Gsrhpj
FM5DHywQeNICIWWVeRGH+7M+uvO796HVVcbEq6YbrVhG5/KmFPwmgqgcMcG3
3hHntnTVHO7IWvogY098X+6l0VDT1qukuLT3WsTedDeGbuZDw0xSQw/Vylsw
zw+jS/cgo0t5Yb+nyMPNC5DHM/I3bV3dKmbkWYlSFBTJhAE30iam3toMJ9Da
eqHjJKi84EZ0mFbvunG84jdvr9aBD7timYNJPTmE3CicgFfOc3uuXJ/lrrTs
tLtHhW9InQ9IZbpcsbT3/HnF2VkwDwesynDyVPz7A1gLDxOb6fcRk9pPUZfC
w1f/C71wZIUa/KaYiMvIMgCiofojDYC7zKFny20oYN/2LITjRw2uSjgBlM5d
XwWjyS/hGwQ0HFILoQuk+v480hJgFCY4katLtSdGXPzOyuCebrMiOLKImXq1
PFzi9NAiMiw5uk/3WiTd7Qy0g1EIjzLUYXXwmeIc045Gvar3vvlk4jPwQ1jV
/Vb4RydO4I4kNGv59sPXQ+zBnq00eQFeShFgFN4tjB1JfSKi/SmIjN3pxeag
39SXJGRDI4/Lk2DOZ7Rwcr/BRFLJXuOp9idLurayNuSCU+WjBHdGVe2GxO/r
4rySEUfO3eFYIxUeOBT1vXE4bxEOw8top8+6Eg6sCm57Ad25k+WcoZOvrZi2
jXCgT8z08LBt5u5tVZnOJsXsmVQnAMSJN7u8YWk9AM1EBut5WaRZ8JEyxnDU
g+Fo6sH9beJKwLfp4iqAvyQMnbZLRukSFSv3qwLGY4dcHRqKU4cgmQdhVdt2
K/iu2msd55XhYzZsuXhB3c3jdIsylvJ1/u1uqWxypS/IU+bTVj563NdPeHWE
zNCK0TTyEfsL/H9+HohvxAtcoXWaYzTz601i6RK8SJpFi01Ak+D1EH+GRHpr
2yeLm8HJxH9ZK1+n3spHknArdF9IWKjmJh1WitbEgt5eGyjlOiukHrnn9dCT
gWXs1nTkkzWe6buzRWZwDgTzasi5Mchs6aZbZ5iMLIN05v/wU52Ie5a451tD
LvslWlUGIF36/UrooJdIhDzLl7GpnPWlUquG3tQZDO7zKnSqpqPikY8TO0mU
GSJM3rcb2aWzP56guCHRrbO9lkkELOUHs3CKMmgymgDJIF4y0Pg7LGAFknnF
Nc0SWQfWCLmXqn0uJ54AAV0dDOA6RP9q0KBnksYkQDTKt3frN/2Hx3NBjb0G
F/nEICSHZQDNBPXDbe6OMvMS3JEoFT2qqSRc/+43YKu3nOIw4uMOUtpDz0Uu
qhH7c+F3J9ImCEUNfLWMKXdf1vzY9/hKft5nCW+m1S95X7WMz2YRBy2he/yH
fvgCN5xND+Y/MU2il1NJAof11xdN5d+n0JpS8CzDRIynLGJ0rsHhq1BU9251
wPFwzfpoU3kbXLTgWq1QvHO0qVbdu9ALxUgk1XnlNRdODIma88HWpUDA2iEI
Jlq30o5JeIXmMPD7kpfawEjnYLBgQ/UOOSBIzOEp4+8CSL6oliFYBfy/vpwR
YwYwcDstHNQJn8/MMPbIL6d9we/XZqcbMufX6RDZxYSINmDhftb/KuxGIbG3
JCkJk8eXgC5VVgCs0d54WWnlTag2aDbqapVINBonSiTQmuVaVowVjYA4j6rm
C3OMYdGFPFKxj5WFwMd4Njg0buMhQzSggV4MfY9dUt6GOC9dwZCyW/BH5KjS
Mn1BTCVVTdB1l2bKfnxInxoY+AK+cg4FP5eCMIYwNDvDe1ct1A7A4P2rQijm
gB40HxI4rjPzeWDgCLKAxelUbiqX5gNmwC9qharl83BAeovN/gVpfU6U6ZLR
dmvNc5H05hBwMQSEWO1Ss12I3P1ELjt35S63wGYPjkdWBkL8A5l1N/SE5Tjd
MZsNZ/s420OOaL5riULxHS4LPA/9D4i/Q2OZJu3pjDWDXdAiXB3K6GYFYEeG
0UsBp8OHoG2GJWKK4C4MCbYlk1hEd62h6snYl2ToNJj4fhRZotrG4zL1fLp4
FLF0xPZ/WYIJhooRJ0jLCWLEhsN/tJpWKSKYVPEqAPKf6E1fyIodaqfHP9zN
rkpqnM61j9ZIf2Jc7I8cLlKtjl/LMsweKe/id1lEUBH9Uf8CMFVc8UJIXqTj
2BfXuXNOvjySCc4M8qyzbw1zVgwtsLQ7bDZthFaHBa1e/a+nwQhpKpS/59Ut
Q/wYl6W0cgHWWxSCHa1+M2yofmTXpyFgK9l9En6ebzcwxStRBfwxhRL3noAu
XeMoM2gBzert6r2Qfhf+Cm1LkOB78dVuradmXh9wzu5QcCwu+t2NggdLBFiG
NrYT5nZfBr44t/CJrzX5fnUdwF5BSesIZmN1LFE1EtjA+ahJrPjhQGtvLcqm
eoofSKpYOUgPb4xICupwrlDN5oRnXVRbJ8QknljT0TIRto6siVJ8TBFFsgXk
TvOkU/N80KF4QQ2aqSCtOtq9z86e6ijWk/gQIfjx1iOgyeZ4xew58D79rIzX
i3Y4OaLXjkg8V4VSDFFIiqW1/n5s//blXLd8EtXDsjUKMMtrmgtg/ywDwUbK
AjKDUPsCIT+OWVo4MtjT0J6bBvveWCvldVJeNAEEAc/hX6/TdZgkVDCFAXyF
oak8FGvCpyBZ53rkIu/yrAP3x83PzRy7YMyzN4uaxyTpfs2zR74sTuY9N+55
fu8UJP2h6rkDJ2PRrNq58KymFNATteY3WbhsWP2PJ43YSOMpSEIk00x/nfO8
Fiizd598P0MNS+CPkIIheZhowlVZGLaSR97vbngx2ssA0w4kV+dWfQvraNhG
J53Kk1z2pRpuSK5sXr3mFTACmH12MYMhzAQBBixScbAiU7ElzdEMf41w476g
U0XAIM7egNXy0o01HQ11kyxqd2wWZAVF2nYV0soguRUQw9c2QL24wUN2Zbrm
2bU4lunA3I1dOiogW9cn0Yp2dyGT4MdXCmtJYoWQYqD162Bum7MZwouIVtW7
OLBTkUJ8txPDpPOoLBJWBbkZF06pGMRdRVqDC6f7ehzu2ECimkFlcjAVJYI9
gTSQYpghjk0Bv0d0OstjCxpAIfe7fb3VEE2EsiH5lcATL5All12+xWReWpwQ
HG9nhiDJSHZjqEe65CTbEu3Ok9zbnkB9IDJcEom0dwqhinjz5BMgFhwr1CVA
ZNqCn4BMQSVINmGkLf3jNWeWNlqoupIjafGKjgNFuOF46AnAr7Fy3a+XJsB0
HWncl3d75tDrxvJ2x73juEJtn1PxiSdOS2HOi3hluTmbXQkzjxKuhCRxilS0
s4doY7avQm62FbHg0dSl21dhZMuWtNcuRaaOf4pUEuiHGctPTyi1xAMLbZae
1DmGRXFEAu2t/KjpX5vg5LTlN7Lh/6n8aTFPrcKtN7tj0v9+6lSFMdivjIfr
KG8uBycTBYpSsN01AtcIbjvPMiqR0VbTyofA6Hijy/3QaNIVn9lfobx0Zsig
Ml7uwn9ryKsY6ZiUm65tHJVvj/JplrdTbThltBKotGEjn3LvD+7eLsL2VC1h
CW1lPt//y7rwFtLRnphilQ3FzCEdkJeznXyup8nDMSebrfPV6UC6cZubKX0Z
Qi+dRViGI1MfeBYU+KgN7NgFPM4LsvDZlroG5MuzJFYC7W/5bNgLUyTSiLmC
hNWxhkX4crzufcl4eGisUP27gAUZePHZKjxJ+est2g38pXgixvSlEJbhtThW
R4JKrVWGyotOw9E4eniHtQ8c702HKFCmbP7aHP/WToOQgTDba58c6XppUpfJ
g6Jd/Zb6QztlQcUgwDSJCZE9LRec8hfxuiCRZMLXuEaubCy3Oh+dss2+87k1
eWQY2Qgx2iueFlXwwHigWVv0OWUq3qzAsSCklmdIhtjX4Sz362UEQlk5eJlo
RlTUDALPpBKtmKZyIj44Pwn623OmgOF0m13WDxxIkEhLzFn387c/59PrmYlA
p9HPxagO7qdJWVjLaJPtBwQsIxwToox0naQTuBHv+U5XOOxkSfE9K7D6Cysj
m/pCdkT5Q2LADrO+bog898iToD+bC4vXPwFzztJyiqRUdyQVKyfpadqHdrtd
R+YwYOI3I9NML4Zy+e8WYeI2llnDlpliW/qBIC/VBoEvDZCl16oEPAOnG27q
m+YfgTSY2y3ei9W+5hEOEfFcddPVftbAycLgNoAripYgMPv6ukkg2qszBvNA
bbJblLJz5jNqwXBfhfnZAoLxFv00IUKRM5xAanCfYsV0QSR2VNz/0noK1Jkl
wOtkefMZm7braWlehJyDoAhpONen78CbrEQBCjwQDRG1Gg/AJKT6m3zJKw0G
2wHa4zYTmyjKbU6kHVNX3a8Cc/XYcHVjlz69VRZOs9CByLPCOt3MHtDVN+Gw
e2k86ellVlW9jljKCaxZ/Vhfwh13pOjxBFl0SlPbWS/iPsPuvPKItm6oJhly
sRMbjAiSScPkyEkIWXgv9CyYvwSIKMpmjtFGQaDdXjMg1xWxwkpgg7MfuxTW
EFcorJ/uITCEiOgPSdpUKMzvmWf1hikfGQGIKE5h7DDr0qODLdj624+/fzbg
LdJ3M07c7bIIHsjJs3v31rUO+nJ1W73TQZZeuGaCCraSIO7kCM6cjXCoM0rN
A0624C/furlTh71ninGINRXbYiSWVmgCQpg4TQTuwT7uwyKKR93uyMGyaIvW
JRo/P68hJhn7YR/a5HRPmKnMgro7LHeETn1NanBsg59gTS/Nr5IH+HnbRki6
rc+sh8cKxgeXwFSW32Idd6aZlErCOY1IjgNZymG8X/4l7gP6BOwEGFII65xA
XSzVMOWZQyg8SgyW8/xUAS1UNNYOmxjiRwcPbY9cAXy0Y9v9bzkO/ni0u5hU
YKhN4Je7tKLUt1oL27b9+/KpMpNcuus4dZWwAXb4WgSA9EeFc+73XadBaFu2
9bYCji9LXfNhqNEVCipGzgDEPMEcgPw/+jxfkkSDn71SQTTRalRa8Tnbf6Au
DtRHMcTcnPfbABZtIZ05m89fsDl77lxo5yW478Ptqq1cVKtazlUeAW7LLCuE
o4qRT+NC36snchg6iNYZErCqkKBUF1MW04M8eoAn8tDCQfFWHq4Cr9myrrtM
FmxNY42NHvTKu5Kr1Bpf8HqiwGb+Vc1MrIPBi0ZSsyS3qFiJX+JOoAFC4OUs
XhAImw9PH33mW84XQs8n6SRbtXc8yKW+0HUSCrMZe8rgTTSGvEqbIqHe2YO5
8a2cSUX6L8A3SYobX0TEWMkn7tlraWvFtbufYX5vwuHjDwuWe6uCzeFM46Hz
96LJJxBSUMlTggIBjjMR1TbEepCgYaaK/Mu1CARHkA8NQlUn8YwEpjwmhNWU
rC5ydf66f9MAeYmWhcTzQFwls3hICoF59DHtNvY1gp5TuVCn61H0LUf4thmU
BJeWkXj8OBUuadFKbCFnQlmzEqcHBQZBHT0rrKByDif9i05o9PZKPPWiJ9rK
7TilInN2CJJwNHcVoqMFNZJgnBpPTBFk9t6oLOmQTtuLqRFs13p8trzmD2QP
FKGeo6F/ZjkTTPXAbK6APSRgkC3mOPCdFQmqwDoyH3NStxkYV0WkQICC1GDm
9qtRiJYWwnglkdDPqETWPr6/rjovfb7cpmbRuwYF07y2tn1dAKtpkjv8PWYn
dKo5psk/Erv0GtuSM9VLFQ2IWCt8Xx/0IVSTuohB0Yealbr13xv6k5Drp1q1
Qt+qVbhSNeGO0OnD5ZOl9r4bfwL4ysqa/J/TFOBn3PWZA2qnahw5e0NTk7sO
BtkP+nWVIbBypGWK6OimUhG2M9nsHImUp1edwKd41ICWYikvmfkvR24/8fE2
sarhM33dZZqlIhy/E8NcxD46RB00DOmn3lCx77hj3CGH1G8ViZovcKlEffWN
405HYt5H1GE8CL8S0nqDP62QCywm/3F4A1lErdxBHPVqQEVBRklSAYY0tTNA
iN6R7qVcqkUjj6y0S/9Cbim3rlTn5RPqDj6omaH3lN0GnyGYWjs3zmyWgZKG
pZZavcu9eD1JNfJ3f/KD/opgl86LQMAIS8kds43j4fwF3UE3Hpzx5LMG6LQH
7Gn+KcolX/zczTprY4hW9bgNqX5Po6wuo7dxbBl9tliFcoy62/w1baWg0rqx
vJtkUNINc7jVPtBP2ugwf0i5Dbgjbh7HQzPmawAlac84KIb5xHA3kocpNouW
e10vbZ4OIqutgJVelYFpPSBIXOti/GYH0HGjKV+Zo2c2hPbe0gQ3Agi8hA7X
r6hgvdRnSe4ngDPWZ1T1luZ4GuHNFPvxzaRbkUtpdNVcAoghCnSyxyMhIOWb
OC3Y5mrdsqto4KN1SGj8mxPManAII5Z3UK68wsUWs9GPONeDFt9y64P9HSGT
iqURrGHYBnQHUPxT6Rj/dqTQBuvodcm7j71KzY818LRZ8kR3kPknajS0EcGz
qdBr6UgjM9Awm3NBeHnHC9uIlTe3lXfHOWYQK7jC3MUHsA/IvkDNMjaC/Nf7
u36RqH39a5Q7UKk1NPANkZ6DVXTxTCR52OXiLsH2OMSN/Cu9TMn/sULxZN2m
Hrh/7csd9NN6y1yDGWiWZvJUlqNJpjhklKCZopOfKGXvamV1j7nNyWzAmvb8
sNJJi1KDu8t8hU8j0IdLmXPwTqIurAGdW3MmMG5FoNJuoTYXoRskrQxiz+zy
TZm5YmHjxO0n1fVj2U4/BG+yUpqu5z19JYrAVa893dNDDrnbJJ5jr87EBMVr
Ixg7UTSeCCziT1gT+ivvUxMDJr7UBtSmcmJI5uQyWrhBC3tvngFQr2AQls29
tL6zKzCFTBpOZqTuK1ggqmBF34Y5iWUYTy0ktS1xXxf2YmYNPzlsJR53wv2m
IiV17h7uc0XBj+CLUaj6+F06jFxJmgNd9DVeHn9rwgqF8R9JRGvLcECi+/n1
tIbtQ24hbuTFDJOckiX1/bE0LSZXYZ5DMoJc8der99VkCuDmBUlUZ5yY+hWc
SyE1Y7uVaH2rGcRIX8MorCc3G/2WGX+d3/7pfrulaWRA+mRvEshVIRkJWGdj
8RiYG2/XHbV1UygiM7BiEetAk+gCpuf5K24Pjj7FVWFL6SDd/xlQb6GPwm5T
q8Iqa8mlJ8JNnqjYqpvgScjuXXHRSnaVXdf8W71WqizcZ7lyk4z+zJ0B4HDl
NSeCSUESvAZw5rVNsA2cvfNXYB181IehHUNY8zAOPlXdG2QphbNkA0Ox0fGQ
oGCCH1hdOzdZvATll5IHAURf6mSs6Z+ofB8Qgg2TBw60V0znQMigEUDDzAiA
lhD/qpNs40bzavcOZ2mCxruaqG4z7D9x6QeiJueWAlklxEq0NUlFhe9Lr4Ww
IO6MA9wXbyoQRMZZVv5KTufhg0bR9VxVAHWkBeOXuW/tvH3qoggomIL35PdV
RNeK1RTZnMhdB5Crt1BQ0Be2o20P1W7yIC4h1CjtNPXzr+hNqMT08dV/cxG4
C9P32ig+KoiwrVhJRD4KQhp6YWhscj6iSV41+1VtWQypA0wRqQyXF7i5BHCK
pwjVk/nUTL09M2b4/TD5Hv+rJTxx7lO+W1HAuQL0bAsVaWouZyRiBhC/UizH
l9oAuSx0qCkt+nvBBc0YG/4ZfaukAabtae9ExdoHh+MKZlyH/ucR4bXkGiBf
qSZ3iHj4tvelsRplLGpntaHOlQ+FNZICn5CYp29obaLR/7la5nipivEyTZPB
IJaPAr2cCTuniPDSBfWW3oOZ6xS3kChKa84guq6y8qXWGWahdKTtxlaT6GCm
sNp6mZ5+2CepUNnosE1pFa6xP1OUzgLsLJY5LYuZdJlkRafYL8ZcxsBoHMF+
Rzb0W6OjRHf/M49ZRQs8jg545/RvEAbhYyZsMaax6wW98Qs0oCI7qJ8pGuI7
J2yoQAPtCgZqRwd+nlfx4FsdmgkDLXSOxmAR+JFVi95Vp/jl5ROKL8qoh4nP
LIQnOCdN8TuCFtAPCsKJzYwMWE9NJPlGimLUbYgcfOZysu1Hv461bKH7f0bA
5YpCEd6fTtE6BCVBzEc82QhQXPDpXL4X9gKgtCXQWNnH6z7kvG12RpGEFidy
HJM3tq02Dx558Q6bq7CJJaeYGBx+z8FAM31dw9NCHb5gfUdqmCK/Rb2E+L7n
TVb8tk0HQcvD6qSWU/Up7o6pos1ma7PNhSH5boJOybwzA15M/IDsixdPJjiW
pwchhrXawrrERXw+Hs63yRwFJUQ4fdG1PpfLFhw8wgJGotzHxL/ezMTop+RY
hSsl4OVXcgkA6ZMIKxsqC9fejMcWhKvyJYXAmvS91eEy8bL522TaLXBgPZLK
4nkdltZxDbK/xczpK1b/ltxvpQnaGSyxGo9v339cInGs5etV1Zxs/7i3i+hO
Ubyw1lSsOaaztYESFEpxNSQqbotJ1O4TcQmpm2wIgIkjSeMjB60jkAHn1o8i
Wjy9f5jOcu5q4MMu+JGW16ly0fvafucqkdCr8JvW1rPQU3YFRi9G5jls0CPN
TmcMdaj8CYhXr/k0puxolOSpqej50AhxQ/Q8615LKt8b0h9AVpMyLKH1nPPh
j4yI2DoqD11q0vtGsSJaAYXo04MbB+PfgKEzfv4ffHWsDSVXgc9oW5JVBuVD
QvbKYiigZr5GQAhYlruwPQdyLKIDEpbYXJhgYdF6pG1IFqB2BZGVCbtb6rYl
B2FGSBE+JhOU2gQwokRjXlzAoMBh1aOT9F5z9koVnsLdH1jTrKpvD6K1Rge9
CfVI/ZRvHygtIrv9Cs3TAVATXsdnLRkOSkhk2OeJO3CA4qEG5Nbhz7wmn0zl
Im0O2/hX4zfhu1PWEHY/o9fSRiw1aVAGbMjW2wLCk2GgGBQ7CnOxEP1MtSHv
5zzm9zmkeOIUvy42xZhNxVMUjUUnwcyiWI9kiuH4m3ecj5vGS8hJjldEkHOP
GzQlTV5P3epxoaN1it1FyWYpSuoR4YNdGYreY303ThEcSyWJs4EaeLSxw8mt
+L/e3kQOndsrwWMJ7+IqcnLXrHFg81tOE3ATBvRAsuv2f9Q0XINbhvOUWil4
+o4seSXRwyM4MwBErqpHotZF86fIh5HgoU0iyu/yYJLfHpIy7Y7vvWRZYIt0
yBS6232V4MonIEuIJz9+2JMnGmno5s/laRsl/JSZWgjAFgkvldtFVl9Jyn56
gwBPsIOuhbmps5kQa4O8eXMdYFkYLkvKWHypsesRvWXFGTWWRyFBwFKf76kg
CAi7Wtn6oy//wIADcS1uJT8c9Fr/maOTQivlunawmA/kEESSgOHQiDGAF8Zh
40oxvWQDwzkoAVJZ9ndkCxbzscIrRe4TO/al189FwBAPGNszD35L4C0zlOLa
kOSZ5ng9aLEv8i4Ye7gnuAhRWIafmXOFRzIKefj7SxHVGuIAX49ME1a3/BNm
2PNebQiNKmGJfZiJKApNxCRIERKsTc7pkxCZ4Cp9LF3Sv6Mcz0CgDm0rFEdm
NSI3ARZp4L7Kn2WKbyJBMoGHJl/RPbSHGjWBdzpFWDF4SWc1ofrY0itunxdS
k0/dXWBWBjkiBaFNZ8ksURjWNCDifP8hT+nJr809ks/XoiIC+sLW8Bc1LnGG
q3YwoFEsjr2xdWn73cH/IJJBPUNBOJFp3oty+2AYcvKb60W9LRkUsKr7W1Rz
RL+0BAu013AcUSGTuRpfGmjEWdeC/h9W4sdWfd71vNFSIV2+8frx+/zgZttZ
jaGEVVLXI4BEIhbF6JnLEFFSGmVZrg6/k6o2HLD5IIP2wLW+IRt10DadSyHX
ZRUschNOaStIcEUN/gTS/AE+ss+6Bot9VkYk9pb7AbHM2bWvKGMj/iNXoYpv
LYsTVNJW0FHKbz76DTLf+kDFsHbbkPe19zcdTHw3f67Tajc9V8ZOQCV47VSM
tIIK/GkfdMAA+aSKRtauUV7I3CJexbp/93TUGqtljBEl7FcNJYqJSQTt79IP
eb88s0k094jOyfjooZXcYvSA8EyXZHOkoh1gvFhlUsozAirDi4Ocr9S3u8AO
ywImM6lmlIAYbfgKyZuT+cRHgODYhwLvnx18MHO64FtMPUwYnvJm7ZVCkIgr
qxCiVhhFpkhSL3A/x9T5uwNx8ZEK4YS0qKWMmvjKwOWcLo9/db8Wn5gmRdKH
VnScQ+D8UFawrM41CZzUufI/UhbAO7C0nXCXum6dx/2KoPGVuX5fNH1Y1lpB
WZL35Zod96P/72im/+I8dTPa9q+bZ0go1uryDJArvgvtZcQX+wJudQPJlcMm
6XYrO98GQ+6zVsEYUsN4WfOBX6xoHCjsWxcqcp3oeLgqecAIJ8+SieCw5t8y
yB2C57Yvkz0U/yrXXDVHxf/8Qq21rbyO/MbM1S73y+vjcXL2XhYTAXYQ0Pq+
y8ljInTg6P1FN3R/9UbjXIfkKmM3MTVyCgrELyqfbqi9K4MhbxQEzu8K4x5B
qrJP5ENFrsH2wHLZSqaqselrs/tLLtJ//XnnQMgNZ+aZioeMYvur1NCp+osG
dwprG7Iyv7A6ex3Pq38ImYis0yEOmRIp0s2Q7yuqaCfTNOclbx+kYRrLibY9
FRL3+KhKqH6C+Q+5hrIvL5CVpvsQEj1cz7uBDpjEI0w/328/Y9x0wSXRTs0B
5idtOd+0d/sPHYqsLHuwKSSdPPu2nEj2wda8+xmniMFJYJ5J+c39e1VVFa1q
WV8jllUPs3FLg4kpmxIGByTmfhqwYAMmYTJys2KCpdIkFZ2QL0btWkodq2RI
nsUlmgB1+ogzNhP804Ibu1y4dZsLv1uLMfgSrvkk3uDACwffGrgAWE4kr6B8
5WxGLsMpRc1AuD1nP0H6Z8FcR8iZjv6oCsYnAPL46iKWV+6BTOSgd5G2p9hD
D3APO1M/aNofP0SEMuEPsefDKy4SEQbFA/IwTi11bhSPDzVc1ABr50vgTJfP
m7PK3iNlFkXTyecJdT/L+bVmsiCAb71D3LaL3zlZYLu4xEe1skLbhJrLcHGp
W3mBhiMsEEDNiYnuqduj0q7MIrbCNPkVEOGjmaGDaqnNCk++lftlX7n4HLb4
MT/QcEtpgSDjskpTmay8nzXJl1/O0yipbtX14nevO+vzFsTZNtqBxfML0XTd
h6sh9TiG3quLykFUuDg82Kft/oj37RLf+bvW3Qj5oqvZ9QTCr/uLADOJHULc
DQf5T74k0d6nR/I0d8dR3fF2YbQRc1Ab+hKMWHz8TKQXvLGMm2aEVAmPV5wg
KvT+k5GCuAsBMNj3kqD/Olf1KXBv7Z0WP99aAgjkf0xhZ1zU0FvBT1o9puO1
I22HGR9SH06XUGQ0/tb6C5xfrdRElLAus4f3RyqxdMOKpIIvW3bYqYcvWibP
ij310cYMuVvIU4JpL6beMuL7Cq0wz24668IC9DOsYw3KTGamj5iO1MsSsNax
Y8aswoaNGDlHivd/RzRfOJuj26uGdR5EGzfYnXWpg8isjBGHBS6cQ9UE+eJW
ZJzZXWdlTjR5dPxpeWBNj0KrhkxkPUYL87YdYoEJOFoVvCUCGS1BIqxu6kpr
i7LsrWYtiCJyDj6zhJj+Bex+gE5Jd1pxi9X5MbJ9+gMzvYyPL5XJhgZP9Uct
NUkUuvXmNTkf1SwLLQneBcHqi4emsIrfMP27RugKorlqfhEYyRgZuNQvz3AJ
v2mRT+4r/DwRA+8gLQpdsaBcwVPXZmYs089XMZ2tVlhO/ExfBRTh0HYNFISD
MdYohxI5zMqjExWzLMAMbkWKUSHO+rREdAm/H1iV7O1uCcGeN+ZWC6+AKWc8
QW9JeT82TtQaxhLbn8qAubV7TqbyIdcFKnXPjjKUY3iKlX7jIFcUB1+BafJj
ADJ8s5FzzCpJt5C5pXe/0HF2C/k102RNNEaEtZnhALA+l5u6rbnRipi5LKsp
ipA15ddLJ63XancinZ1UwP++Qa6g/IIoOxrBWPevmEA87rSLnTEv3zxXtBei
DXv28On0ydQO9+uWB9dfM56DCcyCjBym0B1uJAG7AnC/+VYvC7e5DDyeWKgk
/pQcUShtDjHGQhfScZIGMfQl0q6gQMoxjbE1CC6hxDsv7Sm3Owy0lug016iL
LoHWo0pV9x5kxIwg9cPMvjRBStDQLIecJj/B4g/KD/zvqMlvvA2P3zH+2qbn
gTZEf31jjCsCMVCHIeey41U8RclYyznG71SAILgQF0eI9X/G93sp2IKlf0i3
gfDpkmn1GNkK0m7chmOcauv555iihqmCuHuyE/75CwBMf4wkzjO4+QYVaJHA
CWb7hokkYF+blI9cpuZOOoqSqrzkQDYljgrBI7rgQUeqa7eeTVYxjqorX8uG
u7qqnG0d3sDvsX2FN6+1n197DXL7lyeSs2ly7hvFA5dLtkSgPwaTmD1gdKke
CU2BxNqyVFg7SzH6kw4akmSSz5zCf6FflMh9SzHegr/LD+f8M21jQSIMVTu/
TRVJ9oZrAfAGFD+VvO8MoUnVifBvGS4LCidin6jBlH+UvQ6O12R8SQ9ZHW1g
BOO6y/DLSFNQc+fFjIv2wP6yf5XCLvSn8HFRF/o1S0dtOXZXPLs6Y5ungtPO
tERyQGXhMrvz5ewiz93CHfVGb0QCj76O5lbyVR2uO0Ylr/UGJlT6hgrl9IIR
6zTSFf+EkCfec+st45I1guYUIsdvNIQc7prWewRSXhypxByGTJ4maRyyEflK
/HdPAtYwvgoMCYwzMjXG4F+CDB35ame+14kXIpGgvfBeVgi25q/5yf+dIU3s
BTvuwXFt69WVDF9eWWDc3L0qAy70wI9XSNxVOJEhps7U1ixa4wo6LJjtY/Zr
7BJH41JBCChSC02vbi31gkCRDzPWN/gd01udqmZH3XyV/O8WgtraheAFenXh
hJBvNSczR8WDrcN50TQYWAsbQVDWRWzghkeSynk82h2ED+9rTRZFgje9Ff6q
tpPtECcKXJxH1YfPmeF8XZLSyaGHkGz4yFm98QZYhQbuJU+J3ImdmSebPe6A
mpUiRnGuMkqtrQC24hByJ9cb5KEU0wrl/v3H+40q3MDxZOaVhEWv/xuRdXAG
Y+cw1IGZ7sr2rLRZO9spbR35qxhRDlR1QRDcoakaJj1IihiijxpyBsKCjbhk
setHEWyvTEw7BECHJkKU81ib7TY5zAOssnJ/UUcUWT7UCku4ID4m6sx3cG5E
515J2lx+apMCXtljRwcvQBGbWIcpfpVeN28VnaK9Eie1s3gffeqQo+FCq4Dz
N++V82eyFTFetGZRPii6Gaj0HZDg9MKHWbfb68qQ7GwVO/kIcqg6ihm+mzoe
x8Hx5RlzzGG2ew6S3LVsaGOfX51qqlujr6BISzWNZkbXZEmXP7xvWLMBF4ja
RGSjLa1/+g1DnhaVwOJWFS8AEBlDDX/9OI8EfQo8IBSXf0LayqV+TG5gxrd7
22X768dIxiaFdYb6LcuDQ03GZ0Mntq298+6wfBM6czenb+nwYG0vFFA7usTd
khrrv+Ctny60Tkd4uh6g73X98Y5Gb+6yjN/wyzb9OGXFlUVEVhT+w9HgTOuG
kYeI70PXNe7uMg/2BJOq38aE4h5lsj0WAgr7ymmaGwrXmBftjeV+15amohEd
z7kE+UjqglIsXtZt1CfaSXzjtMy17P93trxG/lxS3Ecu46zL6Gen8oysgrRl
DmPpv4YCnRgNKDntZrUQysUxHkmzqG67qRlcaMmGNiRJaUXaOcgtfteTOPxU
U6hql8IrzOGz69IQI4pPZezllW1NSj4fQVjsvhpihKtJclnFXaCu9jXCcKvT
1ylFojbIeYnO3SaYUiLYIUo/S6FxPHKl1mfqtxWDaSOT6Mkpjz7FuYcB+tir
bYp5embipPUeUy/fwOGg0G2MQu7tdwh7mbaDdefmAT8nfMHfD4+iO28jh31C
c9GcvLnx7fsN0GIFYxHwxn0QpkHKkrKC8S7XzAwl4VTDbGXZUE5+xBsTSypP
Z4VIZD0oIgknWOPGAAeG4ieMYkb1BWVcPUpP3zHfG7RYablqnZrYPHfFmD4h
BLsno4W5sHIZimGYvYSmVYow75GroRzJaZriXjiVA5sRk/I6ABenM98YlC8x
pVI1m+noAmUgoPtGEEL0A+lXcCQrMFNGG4ogylAYrFn+fnLkIKKYDUz5eIT7
HHeT/UScZVr8cCg5omLoc12+yCgRcSgCKiUhH4rSlYlNSNebIVV0X3uBzLI7
ydey16kzBMdHuNza7STf3IRcfopF39Bn4pmkx6x88exFUqcFqCZOoQByErXu
7Yg8XFcOzSmTp05iF8lCJLTzpldYMnmiTBQ+La0LFFOf6gQhbl5pC7phTpTk
IxcDZbDAiihPLMBvYfHOMWRTFWBDXvgJQejccCtbrJRc0/ralP+hJy1cCQI7
W2UnFoVa6wqH2akEzJkT/ithbjO1Jaov+koopwG++0yB0qh/qDMtTLMaPVo2
5/MCbYUJYSWYw3P1LiOjxefxKy7zKIrlQ/NsbbhWQfz2EQwnAp6wLwjPdNrV
qdGtVZuXTe0ChjX4V4wOcdUZxnJYcL8mkqA2b/DSlMKnAHYrG/38NhgbrJRL
x/GirheWSzWSV4e13J54IBiJjd1oTEs2J+tfa522sP9pM6gRYmugJnueKjvf
nv4dH1VMaDjlPgfRDGuURWXyp3vVx19pLCvIYTIzWp8jh5duFTls304DjZT7
gFuE3Ce41VWBylAkZ3RltorCYujwiK5ZF/nlLm2MFBqkLqoQDyNl148CoV+H
2tj+Y0ZAsKh4GJyMHD4K9p4pRw9o109adhLXqc0roc9hecUXSy7bAlKCmhdT
dTeGExXgnYxNp7jj+4wua+gTAV2BDnmpiiFi/9/TXjgNQ9CoW2t1Ry6imEuW
E/NmO3K9h9GJ+FG3nbfbysLG3ngtOdpmLEzz+vH0nYydzPbHrLtVPoe4w329
7FnmEO9XZ+ZKOLjefde4cOS5bb6DgHZ24cm6FNWi/ZiHlt5F1usYyCNTvqJK
8GxiIFAl89jFCd1lSar8cibKns+23dbAiOOdc8VzPaiC1FZQ6iDcaYCtkpQn
k0zd7PQf/vwT1f5JvDVfhlygdzV/6wbB6OEw9OMg4DeIUF57q09N0Gc/NlI2
tG0TX/RZ/9yCbgkjugSiBWw9HfBdVv27ej6SVsNzvkru7wE6f1nKGtmVM/Cw
kYibJrUDrUJnfAdgfFxswUwazknOIO+4zbuzKZGMcfcIiehOsL2SJBwa2eOS
jad3nXR9jj3MLBQuWfQf2VoOrNV4RzNcRVaKOfmHM1g5mH5+QrMppmnfi+jT
z8fhAwc5lmPCdPryHLMp6B87NOQ7Dttiur06DIG1WEX2F/i7xjSeWUQgc+yA
496FO70FUHEqakXXenGet8xc3UK1hU9UB6aXrXsHTczmEKIWWbEod5jTm1SI
AwOUGZCtwbOZzujsOCbajnrqq5lwQDmdKrIfd6Sjkhb4JVGPaYFxosDIwZ9u
1zL0GDzRFjGAULheoEkT34q5o78gKb8gk6N9HhwQ3fS15i6Id/mtBBv3Cy0j
+xOe1v4yfq5BseVqqRyCF2B3bRskpzC5PW74oRFjOwmGLUpdCtuWMKpAJdeh
xciklKMa7HuFlei9CG2AKO0VqxVK9arpwbtWvhAVEiZfzf42phC8/ye6LY5a
ZwpMWdTHNqhFPGf8L4S0b9zSs+uLDqUgC7HbJxrg473kvsZIh7d43zzzAtLI
xNqHe+uwoOVPjKywnqSrJhiIyYtRYp8Gl3pKm3YzVv0nSULNDtISbxmh0EXu
2DtyryX+9IdiXNJpO2Ju11VbB9B/yum0ND1rGof1mgePQlX5cqeCmF7YtJ9J
jSNws99M6ybFwFbsVW0hP7UaPVovckD34lHx3nGMsgqZjXSpoAv5AErIvXBH
n2x7Uuoe5M0WGmcNBmnko5P2CvqiLnygVpxOY5HyuhZtDZ+t4eTupWAB0Vgg
gEnYD800Pov59tPuUJBuJBlYhDJlV/XqkM7Mw1i5yG7SSrKBbUiWHTO7bUVm
zwQzER2zHpFE95/KPWR1N0oEbW1rpht60REbJUnAJTa+iqTPgX+PV2LlNdl9
SsZp5PNRJMnXamYpBnz1AiTgMwUovqafBMYmfyJXdnyoGz6OEEL0F7QEpqru
NZqGtQcvMEfIq1+WI9UGU9IX6oFmBP7J4W/PC+GnVIXKxS5VwgfcCWp9GZ13
C/S+oZxsQXI44BUf3KnFdKOUvYD+6kw6zz8sDi/zUEJrJ0cCRjOIE9d0NDiC
hENBB+lsKe4ovpa55JzRKUL5EVYx+ynNhP+m11Au4SZYJ9t3dAqLmb83JfMz
2aBPVGlUzLqRkjTfiKn9Rt8M6IUqWT5b9MRR5pNGeZ4nTZC3bLxwZub7obOU
7IDQTmcv8hRUPanbCyfd37FRK3Y2O70MPJDmjyGJCeV27T3oGMdxBK9E6vz5
lt08RAhn8eUmEFF31+3/7bPYk67RvfvTvYGjO+04URmDV6hhHAdK79LqMi6c
P+VQldXLX/xhc2Yc2tvNbXwkwxVAQFNdE4zCnTiXc6lsaqaxzb4+m1wQKZWO
rRZVvVGKvas3gD5OVBYY0exqbx8gsG831/UAr1cuNOazHHviihPaGVYpuN2p
DsmF2ngPPfxz9Z0vJJ29K0h4B/rwBs4jnyxziyFnZXEI7FP4OlN/TwK/q7H1
0fxkyIYA1WBHPKPGom7xy4wFvGFDOzRpAQs8hAtKKrj4SL+Y+WZau8yCeMdW
dNuhUJtHU9AE397nOQoiIaG0xnb1fG3VxnKh48kWnKQ9rXPaoSzSUQGc+t/Q
ZfPEiM14v/vA7zUx8Xga5wKhTD43lUnZfKjEkXcx38SmzqEmszzpRhnevpK/
NfE50xYgHYY84p5bnAyiY9auc7xzKHJb79W0/N+FzVpOyxTqJS042wkoXIND
RtDjUu0cfO4kZtwWNprJn0ygJr6QXUNgkPwArgqmm9kmj5xx+OMITmdwx9BT
9Rxgs5+cgXnd4lTlfrb475L7l7vcmfX8QFyqV5hfUH9NFFYiBvmkm8Vhdw+q
SememwmcK7eKCHNt5Rt9R+NlkbnRAYF49sbpiFAkXOzPAHywgSf3AggOzhH7
YepjEOmLubitt7i2/uzMOecfReGlSkS0mM4feQdvgTRE1GcsttKzJmWLZnMB
nU70tAsVxaqyCyzp94sMWlzbH0IJsbb7c+bojRdeYxS8WZpAZlb1SxZZbgZi
JaRPPy+Gui6sXqYZzySonnjtz31vunDLftXpf1LFmhCCRa7nOmHJS/7Mvh0u
Vvth3ZleYhLNab+zXBd+ouonBThqicD4Rf3VK6qp32AXlWFnHVsQkl7BotW7
3G4SE1h0aeLWOvYH3Avne6RDzH1Hp69EQwSK4TioXCxY6VRyKAAC980ZRsiB
hBfEhYydovvt55SYX8dQu5vJJYe/5/c+IM5ZBXQqkehKL5bfs4jnXWctk5DQ
cJhpvcD/x646nfqNUWZyj87gNvix+XwAeeu/LsJVYOisn7Katn7pxuwwr9GB
OOrMjlYKLX6zXX5SA+aRLEamvy9zhyh1JvTO4IAZ1Ab8CheY88FIdokoO3B2
tyllmjol1RRo0UkgGJdtn7BfpUvSFT8qZi1DKurNXHTo3UCxOr9DJUP6X6Lf
RejJ2h4MqTlNlahVRoJp1N8+UNPq5MM71qxvvQEmFTRN8oEMGegZDfbCmycZ
i7UDR7rLEy4rSsKjk2Yl/BMeNboRBxOeK9kunhsdBMua8VqnsRDf9kURqS4i
S8HT9qz28LsQPzuq0bFihZzwUDWsZoAl9FpAb+E8HScxAoFHiB0ybnJbnr4H
Yd+tGgzmTsI+i1+JlaSsSVt6sn4qvDDeYjQiaQm3Nbd9Bj6NOwMwS32FjfAn
2G4BYmqsFPdoWE0KEO8D4uJ/FhOIy34wEoDdSdohrEFLo2xPQGLSCVwKgeck
AFTWQQ97guU/30xamPncnKZELDw9I3mH3KQrwKtHkRDZWFKCKNX2ED5AfoDl
RDzlhaVqog7adi2jJ7Jx96186ZnuQfnTrgn1O2HPhqkU0OahEMx2fIrjHiDS
XWJj7nredKoLTR/mAI4CGKZXe78lb5wyiJMOgwnvZhPR+gCb+wHCsqscaDpS
zkhhWFwA5Pdmlh5ZGBuWDz4QD80SiYQsQ75818ZD9iVpLw5hNep+T45Wa+PA
hHuaJH2JBM8rwKggTvlHkSrfnb7zG9a35Qwp66Li2EM4vQgbnxLi08m3xfi3
G2gT5o/1HW0doUFStA5B0XYs8yyg+8AINSlSFuPN/w3ixzRW8yjZoFhcFTFM
wOlJE8Jg3YFt9SS0LMClcvwnXpOrsj+Bl1y5RHwkBAmflKgCCGDmkjM0qgTs
4EaKjXeBSCuj+npd2TJyrM9VmggnXdqZbDIewsf3v1sxsZaiBsHuLbCBtLEB
lq2pybv8ouMLDMQ2PrKdq6L198L37/m055/NNclwHjjGwn2BAwkz8r1vFHe1
RRJsSQFqS1/+GPkr2nuJf9f6OormuMOlBWjQMut8gh+J8e3ekCQPikQyDW1n
qpby7QzYpwTwXhhDbM4pNespEf5+sTHIMuG+Rs+N7AKzX+DHB4/Ra0yS5Prd
yLGlHzFcDxNBjShjrjFb8e8kvUheviM9kPtXxliR/Gy70+AXqoM8PlkOzZs7
9mPZfNR4hy1v8SZWCMGcgyANjwlNC5Ct0pcEfzlz4bBkdr2UhCSp2FPNFvYu
pDYu/XY/bsf9WMoD+t7tk/oDQ3c0DXVv6EUSWPAj04IpF3CL7A2/Nm7FEnJR
8G5QFEUya+DQTQWAXoGR+5XGKmNiyXnyu+EpmBP01CFHpMOs7gu+RSs95CzD
7Ztt5wvVgkDuI4LdSJISzL71S9xBfewmstDhGtrFJeyFtWCEGSGH0a+xJd32
DzQ79NUrvdgu9y+VAo+NubSgbt1Fx2vnCcTyJpnE94Sz3O63eMPb1aeJbo9e
22Ipd5YcVxlENbzz+9R7viEaqTg1YQUeggGXB+0c/bacccaiRACS/U5hfcY0
6Ikr8L6hcksVr9PMM3CbHZ1mIjjNbTGNEb8do+1saDl1K3yuo719ErfYbf0J
2NjKVkYNn8FgalJoKPz1OBmd2eW4vdEcZ/6uTo/r9lY6PhE+yQIegIJBDCvJ
inUWUX1QrcLoHKkJNA+MXzVIF3n/Tl8jgvTMF57Otlv4CfaVkZITp2CrW618
hrbP7GUjPo4IrLSCABLcGslahd2KrkxjXIdETF3azlQpMyPmGZdi9Els1z5u
z1r5bYJcF2vJy8iweFEQJV10ZsBuPvsnr19fl+8Lk+HgnuxtHp2zpS0i7Yu+
9G7g/o3XW+930MDfjy0llxOoFM4qWhbOjf1wQ5eMXERyVizHSOQod00Qz9pw
WuMrcFhPPelJzszXXKtjibqAFQcFZod2Zl6xeKKjO3LMDx05nPRHTSezjTRT
YO6R4BHb8cjIbJLA2mPixMzr5KOsTOJG/tyD/mpIyCdKFRdeTt89EMRANb9t
0U6Urlr11cMJyLulJTUuRpo8g4Z+nXY1nRpND6u6j5ZVjzXV5oopuf0h+0UM
CcZ8KRZtbtrE1HFKmBUaLiyrkNp1eqdvSV1DBpUqjyLTWKSA5U9D6Cn7n4C2
M1kleVk0+n5+tAl0qjBQgDp2D7sDBKByfXvt+aecNsNAQp9BXDbOm2JEbf/x
PMz01C9yf9W+5CrzAOdr1YY57j7mASZJb0ji4WFfKtjRfDv/6v2XWxKnYG2b
2zdewyPqneyphD7TV/HfHoMvpd4jY+8s/FypsH74CINQADLwZPk4Nv0n/43c
c4ASolQr0nKugSEt2dpFBn4Z+7xTWRU76nZoCATIBwhbp5ajGyeF7N7uJbCI
9bCw3ZuX97Fftli4kI0M202+aCRY15vaClfAHNwPgYx+4XNuEiXTGs7Uj0HI
ZQY4bgBcgWr+/IeBU6Ij/pklhObopzPBINRmiCHIeUUVx8yFjRIROPqmfHZv
zr9XLeKRsDwqzMMcQy5tm0BLXusjuoe/E4l6WJfRMM07ceNks0i/pG/fBTXN
tIXu87nc8mqQpPl1BiplT0VBdFVbZFlNDJGaSKAjO8gyVrLYGpuzR59QtaPn
or3I8WwRekHUu3AWAffQ/eqcnKIKlq+9QZqVk0MS9XDOyhA4Nv+AsSh7Cysx
81nrNLkqhYrjfpyOuiSEdF/vlOqLYmRTQL2acT4oqUyfeOJqxI90Y/Mp1/9U
ZUYCI+7ecGvvAwcYaFQSbA+sbYYRRhliqFhZybDDLLUFAqac7hbtjmjAQU99
kFejeKEBY9goyxWQ3mkS0+/aP/grI/kv3gzTMHx7g/YZzo6bHok+05R+pkOe
pdTHkdGQdvqiClrNJZ0fBag/QyBMJTSzR8XZ9RBgw15jOUPjVpHFy4wj7+bz
v1tKHqDacvt75FO4oGjs03OohogGiCxq4veCsn5Dtg3YerGt9cHQQbqK9a/s
L6a9PstFpWQOYVWwgX95Gk3LAxoP4jR4d1PX0M6iz1ZuPHDwQF0kuEan2Div
5N1SSt/2xAGLkHucAkh1PRVqRzcxoNv6UzHpASaFJ2juzwEbjWV4l4zWvowD
cnI37dzhkmaYMbVI6OhPD9tGDdTOIaByN0FVX7PANTF403QW+hYEM/iDar6z
yVUOAjqHYCLqPcfQ6RbnqP8ymBQAZobf7Xktd+F4OYiZFz4yAYZJznEIyEn7
prfsh02Q9rqxPFyjQrCiW3eqBlavXtZH+Fte4KSuxpmoP+MQqxN7JrOfXx0r
v2n99mEvEaGvVLZ/HreqUmEbiaTsGrpBfxrvL3DJvZCPFvkiTaPyUErwZLwF
zXn87XBJmHNxQqXBn+vcR/NB7QEsN258rgyYY4tvYA6QRJ8s5zba6vKsji3d
720yWA==

`pragma protect end_protected
