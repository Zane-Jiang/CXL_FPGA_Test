// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EuM/7yq0WGJ/i1VnQKrKr5Ra6NlrDjndtiba314uh2DQ64qlAH7tZg6dGmgP
zWyF7kZ2++92At7MQLWsD7bv50WsS7X80lhR9xZGu8/81M1LWOIit0p/D4dT
Blwb6BOMKkAvWyCTBAqhx3xk9q2eHyCjptxkwVN0SZwAFiQYO3oSBENpl6hi
G/befP0zbPnXgWKBdVMYAVSX1sVfwui2VYRF+kdPV2JPnXDCxAwdGeCt7bJe
9ltstq+IyGZyRZqRBThB4fXC4XVjanEd+xWnATWipEPezMajE3dqRAQDwh7E
IzhPAYQ2Sj6O4LQGPDTGwTNiXaXLTjWNLdGu7IfSxA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WQ0SC2+2EFda/aJ/NweEIvzxZIRoWNFlPlpeAZv60ITL9GITGclPp1fGjeLM
5Ubkj1aJ8hrdLHxSqLiP6a7r7QWbBeegpVYk2sNSzyAhDfHsDX13Jp4RwEtH
qXvzKwsz4bQqxrR37ESndc/viogNM+51Mpbd8mGwhYkISWQXJOYEaFuH6QvF
y94Td2fChj3DABCXkNbHOmrgcWkKSHEzqoQoMwha7bP7+ySPMeOo9B9bu3yJ
lEZ6o6VvhE0WyghMYIVYiIo5zAVDOzvkQDe7WypqRlqDzg6IUcwuzsi8xWNo
NwTXT/wnNCU5pkRGUr9U/ViQd57C5WajeMkx8aBuBA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RBOcoMIKWPqEVx8pGWLbhjCaXguYiKfu3PaWvKHeQ5yZtr9KB3vM1lp5HQ8W
zw50Q6VBXTMVShHIMm9BSL0F+dvcCPly9Oo+CcgO863BaA36plq0Z6oOFNC/
hrBpLW4TFzQ2esJGtLBAGWgYUZTOPxwKTRq5iGRN2/Ps5m6UA9KLaA5Ajxo8
M2XRBgcdsBzX7NyybTvzEoaGyWGD5iFzlkiptUj40QMTO0SClQdAfcUgYB+Z
6nXJl5XUBhD8Ut1HNljMd+B7oDbBqOegZ/2TZsqpiKrTK3a+qdmwRt+jAw3C
9bC79yry580Lp4uaZW5TLbKZs7UP2UTygtHyPKMQKw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LaIgEgsHly/0avwuK4LWDoMLnzmqInGL9Cz4NRfrOYqj4SH6lG6I4PKxhIL7
wS5s0etRgIGm04HrQSuQ7AcN13oDlWQUUvEy3OnZxl8fJ+lxiPM3uKSQVjCT
3/g2vqElK3YsKTREpfXWC/Mxpo1l6yAKDW5gl7JG6y2kTJ3fI1w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Le541JZVvrvof+bW0lW3jqLrfInNaH9DzMTELC/6M9mObLHtLthwsExfKbDC
ifCxUNtUODqacQzg98uZo57h+ZvKD2ONNanVx6jJ95XOj5J1IBTAfOUyKoTq
wgUuAr7IVvn/jzIRQII8GYDiZC6pbHFUHFFEgUBEPDAqPX+bXQPBK/wbhVPm
7fIEr3sZF6xlKlWVg8xBNZWerYEYQ6moUxJ/QIigxS8C6ytqcy4XAIU9fhDd
ib8+MIJy4MlaPC2LYj66vVvkMbitS8P+3odHdBlAPmI0ndL35y7UDV0wKV8G
nPRcw5yU1iBuPYgPihoP9nsLBtbEYliNB3oVGCqmQuTqZB3i00DuCsJ4+6FL
6+9RHVcAWTnkGdPYdNGR2fpXtt/0J13zIru7ef17cwHvkExHw4aVW9mTXZ9o
AmG1HNdphF80c4WC6gBRU73eZroWnLO252upkm4QtTqu89eut7HTVhlr1W+e
3CWCIZbmK4tiL+EV4+wJS00IaL7CSP5C


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QN+8mMRfT6HNP0SDbdkNpGMR9ICoCQtkEiUVTfjkZKGnww8P/4MO1rdkMBE5
tm+uGtyjVFkQZ5d+FbSikgzgfrvatWC1/2uY5UhDxWTb60HscbHZTiHQq579
cZ3ppymTa6seViJz4srbM+U4px9bSAEaaq4sMt0EwXH/dXtxWjM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mqrrtIrxpMnaMH0M5u4Z3shxV27iUOSrGJSCR6bgimYIogQgYRbN7vl4Uu2r
jsLCCtJMeFKtGFwMqFL274GTdSCSdFPr3IsU9cHAaveUtxdwsk5zpx7jPLJk
GngPZBkdbxzBcvtxCUpWx/b0NgwcLqoEeDqmzR/sXWU27zRCu4k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 26544)
`pragma protect data_block
77v2IRsSn7unB8itM5Q0nsaq+NFzcjfxuVwbp71IfPN2hT3Cap0SKaehuRhX
mOB2sVKZYFMTYLseWz8By+qqc96mYzt2IYMIcOWsHwXtJc+ejK3VluYoImcd
XqqYyfFU9LC0f/0aID18rH8dvyqCfqh3FRRTnsGmBf3Fxky/5IO30swkW0+q
+Be25UVgSQy5EyOMWLwOnfu/hDH7cNZNkG0WM/Hk+SF2tiT+O3FmTET1IXpo
5ZDAl+6QFjJASHNW8Jz/P8N7ZxPrT4lFpDHQKPbo6RIuhvr87hVdPtERCpHn
jEfAJWLkC8aT6a1WueE3VtjNaTm0LRmYqQoYrawtQ2fqFA/q9HPiNhuagGgE
mUii9kLpptrZreV7EqMfZ8yNokB+oOasMyMN9qV0Gqrxy/V9GNICu/q0tnBs
BV9bwKfyBYrDmaZRznILAsjzedAc+36jMTLfJ1NtPgQ5ZkeHcIV40lHq2TDc
ttUewwWc8egRM+4Ohf3QN2d0mTEaj17SLOyiZZrwcQRxoKKQxTO7bGc9rjTn
qHjC6GlAeCofTEwOPBdyKv3FPMFO4rqdgFiTnJEkTe+JE22Oa7KQW53NKU2M
ZbjqQQsRGRU5xDAtG8DHLM7e1j1cmoVsP7N7Q8EDcFDXeE3ulgd/S0CmpKDT
F2ylJPm4+uM1/Xm3nvwoCHZsxzJ4+hjABGOcKm6QQc1zvYZkFOyEfTQTCOxx
sbyjWVe8HtEIAlXgA0y8BCMk+fJardLHWdGI2WQhzTLDemyXLFCG+vjIV+km
6vCsADmZv4M0fh7zdqDdjy6FfBSpH1Ps1KMVAdGUPHYcROkzPyX92UIl2AQe
PfgRgEt1ER+K05I9VQBBwyXvGIJgRJNECI8jYbVgYQPNeS1yIc7qFsl9qKAz
1wPrRLnMNHdB19O4IjCXkZ6XfckePloDKBhTVKrbzVWHNG4Eyb6sNsCY7FJc
pFq3wuguC4K87ATxoudZRe2SBiEAAKL+tfU5oqb8iib1qxrZkJGqNXRqraWV
LYJrhpcXpLCCLAnijPTuLDoS3NLdnys/hulqlc4LXwzlLDfvJ03eGxxgdbQt
EwocLaoqCZwGe8QUd/IYVsvqxOLEPKOcq/de0Sdxs1AtPGR/4L+450fbOnw3
6Ab5q8NhWFrhYQMuh3m+ogBs/6VgnBFEj5ye4dt1eP210x8UT3zCv175r8Rk
T4NNuQfiUoEUQ19c4THSrWFRxPiRiR0m7/UyxN7Y6RDAku3wIEFcSLJRhiR7
QzeO74xFc5Xq3PI5xU3UHrxDZ1lPRom5OHVmqpk+EyaHJlAWA51OnOZ74kVu
SKWjO9v8Hk6qQiFbtG27l1hRnVTIf+z4oVgUJenMKzInf//GhGVKnylJA2aD
fEF2jC2UdZuaMr/OLpASJaDRFxMULwByG+gACbvxsxOLZ6gDSFrVpQqxjsXh
GSO7uEbtyZnBNd2pYxqVPfktrMtvl64yr+y6uQ8bIP3hpAu2uNy9I8uciVJ0
71gJ7v6IJX6MkKxZzFnDpCTP70f+/4KYxW01Zn1oxLVvlTxkeHs3cbMSwNpt
7ctMVn1va+MRb7MzYbok3NwmggJ4itMUU67PiYZqxO6wdzRlQULfMbi4XXst
Q969eJ8N5LJ3D36K38bsTgmx2uoz4zzxjuaoxPDjDPRenXODzKRNcdi9I+N/
+Td7/lcl8kTKlxWRGe9hcYohhm+L1eLt5tYos0lPxMbKCg8Bp1kWyrkunbxh
kl61tX8PSgo/1d9GJ0NOaxgwuKI1t39USEsWgjwG7Yxfb2tM/W5wfmCjnufR
Icnqp4RAz7ysQsUn835k4NYp7bAxIFGmfE7YPpSCvF1c0l1bNsJIttX+jKTr
pwgtDZI52rVkhH8Aa633O2byRbB3H9+rTZ+fY20Lcg8++SUlax8Z717n1kkH
+u1uFi13vpZCm1fq+nQooGqZcE9e7IA+58yyLefVGdLKoloskcKmWTFfBqEX
Ilj1/adisTZcx+1OuQ2oicOlk15ec2gM1p+ZcMV3gB5GAKJ05IN4i2HjAXmI
6wBj1SoLBSDOYpwruDIaQvsqLxasdNFtVSXhBeUnaoMWsc/IHS1/8oTXh3tS
xx6gn4tD4kv7Aq1TXBCn27aRRGpUrW6wtver5cajB4Ut0jJtGKOJk89l3tdW
sxSBVf5jLb0IF0V+57VHatD56DwCO406D3Dw56eEJ74mUaio2qQei4wXdrcm
Jm0JtifhzqXi1Q1qD/oFne4N252a0G1HvAIgtTCYrbd3SVKypBpMwT4dGQBP
tNkQJeSVdT92l6FaejYeO7f8NQHW50Z6y0LJDrl3l4oa8sQlUud4Cow12d1H
kQxVGbxGh8qceQaJernJPVXZ0ReWXKjJqlngcC9i7U1DQiN+verYKCCOf06R
SX5NMywvkFVVJK2mw1Fxb5+dWv2R4OcdKSdUdc2mCzl657x6ihJup/OuMPeq
9VxcaJQxEJRCVHBjlL51/NDv//8IU67AhRjLnuVhqEQjHD1lsM82DsOxISDy
phb8xCIqUd0MoYJryDBAG9L3wkXYv148NkB4JXpZgsYDOte6eJAomElTg6hs
xlM8hXm9uRaxNKhq4v2wNoANPoZzzU2cdnkU49HB0jWK3fFLS+aPB9+7TIb+
IfaGdvgBvZ1vQ4R5xY5jWGmvzbM1ajoG4eeHMLYEdO/2ZFiJq28wnfWpbv+w
oQEXDG0xELvjl2Fx+dFrXGdOCt+i/Ap+cCRCLXGhslmokIuTmPsrbiC5aotP
PBJrEXmSADKf8OOYBZoQEnIFjA7qGmfW2XJg+T/pmyAEbhkCekPZJp39vnc2
YOohibIWB9QKRaePWkj5bycA9xL2M9BMK0KKCi660KkTtygvoJHODleVho6w
0FY5Uz6wiTsj9svTjb9DbpxCkS3xsBeTcEmLyx9/HxHmYefs4a652L7XnxsI
2KwuvyXeKLSqduPHky+bYjpRjBYVoPrbSGoLZheElD2JhaRUdm22GbIfVvrR
EJh/aiJEPKVGCiEhsNW1S4uf/xp+8zYxRy8eRbvYcUBdgK4lbuDlHAKA7B6O
qhXYeyESNHpCzgEnJa4FVdtqkuSAt+UlnG3jolgfnOHlxui0OgoXSUjrK1ji
0tY77dP/qM15gYZu8BEAYrOTmTXnjCeU9XCbAMjICp9SkUWIvZl4oNeOxT4P
sKizewlCZjm2IVuwJpUtnI+W57nA6iTiVxl7JjCsKXNSUlNz0dWV0pZdWO/q
qQLMmjwQ5x4TvMr9Tszjw8oF2ZbifiH2tGuUaIvNs5hy0MCGWHkaKRJKT8nR
yAdbaz7Mols/vdxBYzpZOsJM0w+d3xub+rbwuYV391hDDiD5+SCZbS4ZM1op
vUzann/H0wh/bsFDF/b1Rq+gQEgf8wttEePKIUNMNW5vwalf/kDjkYweqbSF
Ilrn0FsPP75wfNiD7si3EbYfTaEcqRHT/9CnnThSOjSOTbvt60vYLzcyyuUK
PnPfBhcQqrRhVDMK8hOqW6Y0T4sAY418ebYMU0o4WgSnURu216PSMLpuNJML
X2VU7hs42aFj58mmeudZZdFLtZ2S+bLw/eZozKhuLd73uT+FN0iZNR4bLdc/
aA39hic2VNe708oaZwaJQ8xAYNQ7tN77TJox452/Zo+dJCtvrXfl2svNdpvn
5Djv7SC9BEO8wnaJooMFRU/fsKMUlSgO9y2SORNxTopdSwzv7O8NqyJbF12J
bvv70N0oDlE1MAGTtBooceEVr4a14KenUcuVML1Fdb2qeYtjSR1pCpgyOH1U
tU1h6ZV40kXlhrkTze+RAFA0v2Nc8HWLgravF6kO0nD4A0UVdzUBIv8maMYV
etdopGm84j5lV+0T6PkdYYN7nWJfSFG/mj2wMB4JSxde8ugFBQV+ZIbTGeix
z9U07L2B/Wf0Mvm1PDcJra64HQsN3f6rlvZUkb2pPEshCBXVQboOdsHsvf85
6cUEKnH/9p8j8Y1pyxdk9JO5kGwOp9lwg7cbM4k/Lwlo52XVfE+htDMFJpTQ
GYP4VOJ0umdyCyaBED/G6jr3m7hxnxDgjQujmCaavF4eB2nwnQgAlpZ8bHyq
e7853tKvHdkjXIV6sYAFETAH+Q5xLYeZVPHuTZ0g167nFhEY1NqkbupAxlVo
zNyj7rtmwnw2kMYxkPj+dvgUZZKd+1IhWlgICmjQpDzdv4AwlrH0JcjHegOC
Z1ok4pww7C7kwaI2ziAnQ7UyUcyQaQK+KXgGNLumgFBWQmATg3ZyH0p+nvff
c7g/86AScyzA8rL/Bra2/dT7sfJml68y4tU7IMIRA65FSgJpNW8rGTNmhfK7
VyfZlwpV3u+q0YQeYCOuttGIV6RN+ovq3UR9Xv9H0ak2MIxivnaLVa4Y1pgG
KtLVeTs9lGSCoshcdFxa3jcjfUnpN13ntiBBHlOuFzpZsV4Y6dajOyeA6JK+
vsLBBsGM5N+mn/dhdxKGXQA6N0Fn6mkn8NWpbeOBb/ciaNnWv5wIa6wGhRwt
PTEyw9JIxGeKez2bosmHvkC5KmTc/XDHwFICP8hjelIhUg0+oXLEaVT8/MTK
DZsdadI1uel0hhBWBFh3KBREoCdI9hUzQ/XhYPMwMXRffharcbHqIv+B1C25
i/RRuHOE/1zIwRkwC1UIz4P4Ye9BDH539ACGsteRBNmUK8K1vqTfrQBYtd4N
Jivz0xahB6Hl97kgPXO37EwowOBsR1F1v9DJAYwlDELoAaCuJz+votMe24T7
H7fwriK40SuqBiPSehV+wSnW2KkQqDtjpitXxFAITRQ6yMeBBvGK+rs/eC7T
nxcjIsgd+o+QSEdkHmdJrYypy1LhW7mXmaglSCLZSqGxZEjeETLP0si4C+jA
eqd1wacq3D6fBZxh3csdoMCPzFAslJxVny8Z+veLVOxSHR+z3o4JIxnLdCqB
FHqEfrsPMfZD63ZvDr2AKQPu1H1J7glvltgDfJSM8KQd6iZGp5NFvJwwLAK8
hqkoEuiz8gLXdC/sdwd6ck84pQntWeAYkw9iC8WnWm0gBSO0eABiWspXrTDN
z70/1PEdux5WGz0MKOo/CQwLZ2X/O5F0tXHxos5N8Zk1bk6JCvd4e/A8HPY4
DTLRWxdsPSDKB3opi3D0AqRLcwIhC6mf6MHKlZ6Tj4+wtUFuzASRd3rm2nf9
BubMw3nE5HpYB5AEELk9HlApDiGPhTNubDKAeLjCXGIBsqXH1b/J1juzmfY6
cd7NEMYOOdxhfhp+4DIKLqnaXPehdbyUtRNtoJT5ahrpda4pKS8kjQjQ/vVh
UD2GjZIgk6eSuMTUUOlhaUVX1fiM6+M8dGFqjGoAXzkNy3wvY3q4JD3A62Am
GNCNzDu6rx/n6+fMuRqcRh1SJUsDQgxD4vAX9b7IAI7/NrmMhVMNBNBzAdQr
p0rcb7b1IO61jh7zGDj+eY+PQo9N0KjRSkE/awcM/LuRgD+ExPVEoWMtTF4B
2rtbiaF6bU6sCpGxjeHHs8I8+2R+mC7AuV1TspEWXPLtLH92hUocYw/FeAYR
WF4hJ7hdtPkKK5zQJCZg6deizLWZbS1VRPeu7hCglISfwLDgHj53nUD3dvh8
aNbozjLHq8J/l4nalVuKGFpGLjZPHyhKBf2PMmqHvkvAaMGv2nef/gEHbrIH
HyLnctU6HxzsprXpXRNQSh4OejUI/Fj9NJxHPqXR0rSl81e9gvnqwarGvc1H
y7AJ+FugdrsE/EI2mldM3ky/+I/dTmLm/4eGY3nvvxZRkfp1UkMMeVRS6PGL
WYTOZtQ3H0ij0FAtOMIsgT86FaofsOwsSXN77dou5FmBDkaaqWagHV+ZsEC7
nAJhPuVVMR8IgsDgV75T345FWLE9dT88DnKOX/RlyPfl4CAtgk7RQzqHL7Pp
SLPxW0zKi3xsp1/oFUXsgap6Trh5sB3GoYPVLl+7K8Q1GDZa6jfWcoVFMOe4
T1jBE/qxi8AJrktgAm9tWz8LBxfjWpchZYSIIK01mA3vYpokYeVGRlHAkbt7
qVCICXUGodS2UIYxeTLnWt8Cbe3NR/jM+l3XfssM7xZwuFWWwbPoQ22dj2J9
cwSU/H6DBe/Ri2AsHL6oYwT8I2ethKhjxZZ1RPCfLTdCbBS1d2ow37f/YhqP
fbdtEdhFF9L7//SMc8JIZ6MfiB22x3SMUAfUf0aIw0twehbgwT606Txd6Ju+
01hDvRd7o1yuN6Oz4bhCoHADzJUF3gt6UfNjTLvAOlf+jXjkJWEH3vpps0QL
OdOw4EHVB0+pmmPkG4+r00UojL8KsGRl7EJ+XB2uaP4YWO55teuBxyTmsyso
e7w4GVi7Yn9oYbtLvU5cwrH4euwdxrY9wXvDxgN/1eai2jA/eqQ2l1tTAs6y
NkqAfXgTfEszwgJVHH1npVFvj2pi8cGrKyOHXaeoOzSE9VIjiM1Hc6vqw2pU
BicCoxTwIaGZRhaoORTZQYMt/mdXfEXWMC/NEU4mktq/hpa5a7Si1TBVMkNG
RLidKvNClTlwi7PxVTbmNjYKilGIEfnmU5WlFFYotaYRb7NVMGS/r9qW+ckv
IryQJqbTIVoVfykTs6eoGegkvn+5E78ApJiRy8uk4jaSJypWgIsInZ/pfMwg
YWQNdXmhkdtpbzHlMaCWTXuI0Kr0506FuIpTFuQA+Sn/+JmDjMC69CgqGt6W
Yky/yR5VyEHYPSJFmAokaQmVMAv2QGbf0AFpeXQyhb2NkDnAp8ZguE9wiz5m
IfvrVpIvWaWAR0MNnPMn3AqHtZdwjwhbiZ5qIVJDcjHpsw9Hp18y15WF54KL
QOZVaJQPcCEyAVvh44wBe/hhabQUX0Ljio8aOhWIWiT/xLARLvdTQRn6B8ml
vg804ofEwYU7izK2VFEXIOu5KL7mW4v9NfY78TmdSzi3j5Ux/Ddg57AY+1WS
3BnnqQW4I1iZUQS0Q2cqZxUY4ybY6fGRmpUF1AdgGb8wLfBZjJdW/gQtdG6F
oNaCTKMzyRzZNkFjePHdy3YVDHDSjXBXI2A8CHxko8jfadnEoeastCGcI4qE
E5BV1riPWgIOEAfnksrEWY1neVnZvfWZrcDFsIQWwxtXPXYm/16aTRFzUhXW
6yKFt+FO4lhKx6ttVY1WuRIvEe3lFd0Q5Gy2LUny/DCSghuSsLV/t7F2BZd9
zxAQ3524hJo8tmPVfeNdVvjCyHLwceEtpD9PTEvDL+8JeL+HsQ/X1PUWkENL
WVUseq9ghKeUVdcEOyTJwnmQktnUj//XmU8WVj5bp2PoSLAccbG88eCPWWrB
4Da3j+HXXpIvaoFkRIRjJT8SRyYrePfwmU2cv0SNu8yoVYXf7WofKVptWuN8
q5VrXqrDGYzjVHGcTgyykMOLzpiN33QS4w91YVj+BJ6ZHaYls6840l3kqH2K
GiFlfdyEppRf6bB41fKNqew3paadgPn9WozzR7tpuYuAFYhJU4YydTDZVUXI
uEt/N2u9uQ1CZuSwAeKs69NpMyRRNVJKlvY3w0j6Xs6X92qT4l1nn9TMtnO0
nl8/grWzY6iqWg5UZZvujzGxGmIBvP/BGI5Gj4qLJvOox2rr0E5v9oVs1v4q
fsb14d2nlLLi6aEVukqOAz+IGaYgfuJ3/IpMQ23UfLCQmruk0Z6B8ksIB8+U
2rgeSNTurzrjaZwe2nojzpptGhOz5l/TY0JlM3eV8n4FvQz19H5yCxMqRpl0
5HXXaUDYa6yIT7KnWOQEM517TlRJ92X7e8vj9QYyKSrBMT5e9oRX5ffpUtJc
F8Is+IZUCwYZs3bPxpS0i/BaGVMQSus/nTBbfz8cypgUkPp1UvIcvePMNwJI
t4L3XYYVJX2Wa2x2QNlMhH5ij/Q1+CRPqTCFR/+iapYhjOucXzSyQihCxVET
T87uUpbEqt8TbtzN6lnGSTtN4+FLbpkmK665Ykg/VFyEGgEsLXpWMbQoggJq
QwytF2CEIOrNyztZ5JxaxXDVwD6gW0qpyYXze44aTry8Xw53Pc5j0bO94K1f
FZqZAdEaq3ssD1pkoZU9A/b+KNQlDGm7Z+PX8MAC+PvHUCihYpb9a5q3xPy/
TuDP2+2U175lulB3OTydnRN5+Tb++LJ2UExXoZNkI7rEaPD5WkOaPq8bmVpI
yQx1mHrVWGqmnZCLAFIL8OPS6p0aghQlHrPT8vLfLnOZOZD8vpgvziHfcEch
LWX6KvVFwRuQomEfCA65/MSbAOty5qoStDbvhvCUCBwicKv+RITBHmFQnHTw
Woax3Bg1CoYvhrcWFwOT2VF71byA+XIxfnaz5O0Bd/4LgC/HONfFBPOxWAEm
+p8azxqCQBEbOzqmzaSR5SNstB+qz0IhzmWHFxR/wN5WJ4o+ywrw8W3qQpjO
pg6tisZJcwOw2HVAHTQ6cNq2yxJwr5JiLIEvIc5SKp9V9/N6eCNaZVQuULAG
oaQdB2ALVeKpcRdphQRsR0Dm1XWUYnoAw5Io7GXX7SqFw6o2eUcgMCA1H/18
XKBFT8G1fhEfDVCvlL1iu+JFjntQPhZ3GKiIbeYN49sNO3TFIieZpT7Ds5Az
0zNpCtHCuqP4CyLLW7TZYNTpjygQEBkDYM5vWsqAbikDhtTB+q8SF6IArw27
S2AlbI8XP/E09WSZpSHgWez1ceZa1BiKONTItD8oQxr9LejFqI1FPDWvQ0Mv
UzzKK24jtQsMncVjshIZHUbT/Lph8X/tX0f7Tu5K9opD/BqmCPVK75gVmfOJ
gMnojvi7wEP10ZmjGzQyD2U0fTayhYS3wjcPD2H+IquqVb7Yj/eqU4cU5oSz
4yaX9gPa1jd36uBwGjnrdbJ5SUIodq39o4yr1VTSXXT2ypAfwJb8LUNvZk4/
uLK5vF8+vWu08wF4DbEe1BSErbzU4FxLvULVskLeaTaNaCx6vhuEWxDZVeKd
XVO4vkiJ2uIFCz2TQ0jEyFbKIf/O3Zot5qCFDakz87uE6zK4qqYbVHIBjHOk
MsnFselEA/gU4s2kRNkR+xcgHBvIDwcx/ISFRFYWFoAK5Cu45Ghi7Aus7xAu
//9o8X1koUx1hIOTeCb8chVaVnBiiKZR4lBQOVIphj69f02Wmw7N9EsE0kV1
3TPdwtLJtEImKL05PSn57gZLio84AMJ6JVQaELJ2AxSJlaWOV29491ztHPbk
mDYQ4xStGFhZUI67OXWkN8xV8ZS/vS2deoe5tacoym576ZnceWMebzc27ml/
VZdpH79gRMT2cIblX9EcL0/UZ8hetvJepzb6R6JCIZqMWJR3O+pi4tSlLUoW
cMhK+jDQY1+0iRwWSELO4BUd1X1NG4X+1ZjSSVTduDX8V5AxP2DZEmEpemHX
eRagyrBJeTaYPusA5pDiCL0gmyYOkKzTSh/6nu9jGBo8grtQRwpxETGX+6+j
7AhmXf4ySfX/kyf2n43xVAAb7WQyhjvLa6F5ES0IqPg27+MpRZ5n/f/cO2Sv
u0rGUfFWawCpoBqol4Pd83H8ioY+oyRrZWv614RbFHFYe31RPZtiMjvppluW
Mol8BrVzUCFcynk2sH0xSkfJ04laO/ymDk3RzeYlbtR5475wqZUbL3RymSOi
JtetSQznBs66DiRkIiYXq7aXdxt+rWFuvUiv/dxXeaxU8TwS0aSUbG72lyb6
F2jyhB8sMdhVLJnF2YO/rWEiMuPskzR8V4tB5A3X5P+jkDCkakN3BvHzYeu6
9eWbB28M6kazjJChrhjyxQzmq0Hs9CfHFfdUpICcD6Zq8AOc5BRLiBClkFoa
XO/S+Brrsrz9u9fNKds1JTw5FVXUCMOvRRzXZNpqeEIqDKCU+r03bMsepR1U
8PjVki91bSPxV9b70C9R7fkdstRocxhObMSprWhtRJRcn6aMLv4bO5JzpNU8
iyNKPDPFE+wMct4B0x/eWZdkdQs8RIiMk0qv8MfrsdQ3xA0PYt+kS8i2P9hN
tb6+zvL/JaBIxkWFjDj0I0gqaX1b2OuV4J8EohQdBwdKgdCr62aZgKs0RTcl
LqeVdelDiKElQhq6g6xx5zdzVqUkCyEWjXeEdmhQpoVbkXtDUIukH0Te0x5/
lqbneWB5cst91gNfuZAUKxiEG+sz21H30Jyt0WRLaxS+E4FMvXy1gCwxk3x7
VrP9jYeWOXhtYUrAz52ARvJDh7qQzxBhrx2wbmVRZNpRL2TYevLFq+B/1D+j
+97IOYqyZ+DVa0k64TVqIiU49UVjY2GncU/rcw/r9H0rXEwiiTyR2jGl6sJS
h12VZz3yEdzvJ0wzrQeehf8YyU639V1H+Z5MKnXgIztDe9IvVRNCj7Op9Y1h
AE56G9KUW4/GT1CfIzdwdNC+zWJcj8WKVumerdESRfU+76yBJFzU1QvN+OL/
JDRbe1ohRRLoshYMOdXWMojiLNgxODsy5ksR9VGq0jKbQwa3UApBhk32a9ml
VmmBnKN6WQSU/rqEN94b9lTS8tEX7o4KNi1a6kqOD9S7BaNYay76C5gLWnP9
AQjTE4/iesk5c0hSnc5waqhkedW12jECdTBi3mj/13vaieEvNZu45/6U/QHy
wsOKwmXZjfV1CiJ9g1bDUIiRfwFRvdRCgretekrpYTLWRZbx+90f8NGYKJF4
KACsLDDmLM7KRaSeR6v2MmyFwaAKwngX13w5YM90YRAu7gkgJxbo0g52o75/
wuARPeC6WQ3dpnqgFwl/8Fit0BRESHoQTj6TsepIOqU6MOrTma0Q2MJ8XcFg
taGlL0PtA9R83MZbUlfoF1/8hgw3Dqh35IMUZfLvWHx6y3pJ3j27f2oXW8WP
LzkMpBRWhfPiwbY/BXDQxuOAm9Qi2ukjWjeNNLca+SvZ9b01d6iaqFubo9ev
VnEntxMVJwOUooDc/ouYNmgQKSv5EkQTVQSwmYWvBT5sIgoAPh5iVMploEEN
rRrMs9+11yT45GYhShRJN1s/VzTNRQes5iesN0KXPufPYKF/WZUOoyl/QBMW
W0jYD4fF23LsUQI9mlShYhruuslm91bDhlHjK2dnTQf1HOGVLgL7vJiuy/T7
vmXsdoo+8jBjLp6BdPWeqmp0Qmbbj38NmKsHG+CKers2JHw1loeIKvyY6RRu
w4hv+tO1nXJjhjwA9K7FIrpfXCIJxbnUvnIKRTgeATxH4tMC3Dt42+PAAGhX
grSmPb216akxi1u+6GLspXuG7svTxsmWEozbPGuNvVeJyHniXe7utmtyRa63
1R7Wy+LzV2dS3ocKIJOxNUZ0evwq2lXrZZdGA2jp/41gHtonEOccPCAPas3G
6g1iiKxHLdEJ/PKuTcBPWxiUmzp3tKiHFtRmFS2cqkgvBPOYU5vIsobBAlQ5
nJ5Yfx9FY10bMPFTDQqooF/QNUpmNTtAtkla82qa5DkU6HdGewfmzYDDZPz0
mXZBydKfC4yQH3L65J1dSGNrymNmTtF49xrF+5jiCXKoUxZUDImdg20F09WL
gBrN6jnezoCjOKPABXCauE10d2QcFvXyeVAgzLDxYw/JGShtST4aG+84Mgo9
GSEzvZphYUqnOzPOn3ZUn5v69oRPQ5m1FbOSaCmHj4essCu5X0jqOccdgSMj
8yu6oZeqHBGRXX5AysE9ACgF5vIDmC73DAGDtJSmoV39Nj0H+HmJi3yVAyeH
sz2nAhC6k4kVSMXOqKbrd6HB9jc09DBGV6PWNKZ58WlXwncV1/L0Z8FizNGT
XTTuvuQ+11SQCz3TKVvBQBod5m2mvdHlYXmiFT8GyTwr/ff96N1CujyYj+lQ
v9bbZYLniYsQKjy6G1gG6ANXyVdWTpWfBJCefMb/ajvCzX4MLmkHUeBkC/q+
pH70/cjOmQThPlYv4C3+/GS7RD57/NQhh/Jw5IKLA6fhG1Rv60A9LfZg2mHY
0fOAS7KNzjSX5Mx0jsY93vKUYqfe3n49JoAj6wavetncuRRKZzThy8IXFPYS
JFFwfP9Xs2q6lFIOCgV3mDgsSYMcs52MC+7QR8tXSpGS6wMcbdnkWdoFp9DQ
BpE4Cr9G/AD8JNbD8e3JeyO1zele1+g83T7Dw5/dYnG6Xqwwc/ciMmNImDQC
SiIateauXP64UqE7me51K7u8QLIHPa0DSJCczqysgXXdN7asLd7DOv5JnCTc
4/4LMPZYm9Cr/MuWUx4Yr1BmN6bqN1hexSlom7ewWs50FNTFZhHXlUmqlPAW
YxdHAT1FpsPIslDjete+Wt5jZZSaczTk1D/FiHq2IFuUHEleuN2P9NIBeW/k
igq6OEMh45eeV8B+w3D+dnv9VMqnJsDL8RB/U4k4waXIetjtoqg/n1R4pDUh
w9sKwhxen3jCOPtho9AfFbL1nrIL8kJkC643qVPqzlUOBWapS3TmutnaUUce
mYz2xYQQLZBPyBmwTTiQohNV0QvPgg2FoPdG9z0r7fnR4423A3zyl2JfHof7
YnAsAdXBZm00ZmVvHw38N/6e3N9vJsCH6Wu+uWk72p3DDSb6JdtI02MO3v/t
//URWtaiQ6Rj/O/+5wTrjLQ61tnZg6VAfsQ/qmV7JjFLN7RAOmMy2gDu72t8
ZtJdujBxHLa/GsXliyh3lX8iPC0LkjluBowHYXciC2uY/KtDHp6MIIevpVNG
MOLhgZDUrxkD0yfo9y5BvNG9AlxS8Bq0fBjS2YUFR+XxoFeeztc6Ku1ex2z6
kWOSXNe+JkCUMs8NE/GiEOOGGaZkPBy+0jBwnB3r2B7lxz4gzZ4l0fDgZb/4
h//M8CE/+MD0JIw104OSOvykNdItkftCx9bE+hyc3tQYHhwimkTlhq43vA3p
6umQzp5Su/T9doOfnV7C9A+a0gAvQWqrHIJtCsDMKWW/YmKGWkSSCCRuy4uY
HvkPiGQSX4L6xbCsk2gm0l/4s8su/z8S1qajqvPglgXlLMa8qEx+TxM3Kvx7
jfZdEOasMFuVS8l35/aWf/1DTxXVnfLvCWtX/akw+sk0ooQyL22cbK1s1JAw
exBqibtLGG/nA7bsUWycAx5CJIdoYfoPYQBkb3BuVlGCpU5Ryhffk1/wi8PT
2e00Jn8vXbUDDHlxYetTfstAKM32fZ7Mv2bY32pNv8oSJ6U1Nlzhj7CQ2VHk
9dB1iv94ORxtF0J4PCV3CHvNBDNSAn1Q59qSRp21HRGBbvHGHwW90Px3Jm91
ggC6nxugYQqSlSRVUNbwikT0Q/QLJQ6F2nasx0Tg+wltsm+eDo0i5Gf8iw5a
ZUFkd+aS9WQOANXQMqJAR4JhbxGg5UNJMkc0NY9bmfJ1Xbpc0C0FfN/mfdSm
cojvpKeOcZTuPdRyCdaugKii0jEZnwakSoY6BErghUKoPQQ73K8qRzO6XrCp
qCbC5G50kUD62gIvQE9WraFLejrEkUU8SEgV1gEabFvllAh3EMlqLcmqYbK6
tIKedcextZ3ESd1tnURTRiSGoqC/Ap1jMFMwOGfoSUWhB34c5l6182giXkSZ
pWdETlTCW9oxkU0NV9KDhbQFMI/bNq9o5jvOiSfwEKpRrFlj+DKBckYnYc1a
UefWzjJwc9uOwz84zPDl5EBDmbfJHrHJN/60CqjChSP8mFWv9vnDFXbPHG1J
9cUNDHdjeLYr44+y3t99ggM4NeAY3y9peTYCrYGu5RTNrGcn+q/7NC5X6S09
f6Rj4Ajzt6tmjQdHgV+bsGl6vnYWDQk7EmA7EB2NNIqAD/O+yjtgz0aphpp+
9l25OkAWsv+nB69ATt9lzTre9BTVkkHYyuvWUHfOWnFG+A3Np2KEXFsHWfho
Xg545D+CZ2nnyEhnZmJQtrGtHbmmC3jy8c+Gd1pMKp69bIvvRh3t+T/nFEnv
8YUr7XbG118o2rjoE2zMYsZu7NCIryItSC18fU9+6mT7d508HrMsTIqRkPTz
MrlkFMMxCjsBMeKFeln2DlEpHJ+Mdrd3lF2VwEDuHxqNR4Nlgj62S9iYdU8P
bxwyAFSe1f6xEb+VTYNuByclXmXL33PbQ+uGWWj29yKwXtsTmFEUuvPBMpSU
97kPXIXRxhZFh2nM8jGqVPe1J6SLAv9aI/sqzfagWgBW7+Re8t/BwXj4THgv
O5cyW+NTm48kIVrtd2JfNC0uXzdxFA1GJFzRuSjc++YiwZCmX3Puaa6G9l6P
zpJ8bOmAl+HOEYmdmVPtXaFnHsQwDlMd34wecstzCEQjTx5Q8pYOqBI/6b2e
PhQnNFyxbs9VPoiTvCM3UYHiuFqDdkfwrULpEsyjMd2rNzilv4u5BPKosjKY
I8WLt9W8+QAUA1Lryhmj6P9iRBS2hLDhrhTdZ6uAYOqbjEbSMqn5AKob63r/
IQqyT1WQSajtdjEBksOz3kWoQ6I//IQxVvgf4r5dF5V1JQeybmotxuXX0tYg
Vq615egaLrq07Hh/cR9In+pzofTpDH01gkpkude1NfJjbre+6QCGQRJPXvC4
g6Ji/dLuiaxGWbO8cskegQeqohvgfQ83G3H7OHbINd9Cj8Y1at4fbBnxuiOr
jiEG3+KmShMTr8uit3tzCD5gAZc8B8SgC3nqjLkYghiyIuwNanN5gW9HspeQ
bhCrUmJZiYo3Se1t5DmBOwS5dTW3CjYRZe1+4OXs0XAF3q7SSKXS2zRFx0fx
wJrrpmioLaWxoOBbDizKC43u9SLkSpSM7m1bky8+zUBZcjkELTq4AKlv0buy
2qhT8bZVf0PgexsbBQaROl7i1403fgsixJ+GwxO9Ip7D3IMXWF7DaJO3YAHA
mcqW5rmw1M393dlB1hfFmdUE4IiF1LDKZlDaML6uW05eVm4oBbjeK5AX/ZWL
PpqF4Q0fE/Mf3I90yQZPykiX2EPqHO6Z2xG+QXWdvEMHOyQbxT2KjzXmp2EM
Pz8Ea/OdmtPwr3RU+OQ/d3UHbHvzsEO0aTZJbSAIvzPxaf2tPhvqxeAdQXq8
khB5LYrPdUo10FHjIoomPYUwW2/esWgeWTbTdz1cs/qM7rX0OXVslWIZgQGJ
A4qb3fjmQHpvv7/gj7vNF28HeEZOaB8nXeckxJVA2gq5VwkEMa8zJLUxQmzP
Jsi/KFkk1HTBWJ6tWbtLko6mlcMPi9rnOvR5/ZA1xw/MX91E/2LRoAXvq34D
zD+vzxJjYtkdRI0GlM3IdLTxQR354SXZQ6nKYex9NEJTW6e1h/NA/ww7vl3j
7yCJOBAqbqo0x5ZpXKBpG3vrJoUpUIxcOpLMcZU8s1h7aaCRBy+JtRsQcLy2
HlkJlWtgykrhdLJQKVstlX8GSGuMh8T+k6uiTurzGrcBSpPa5hUOzBpV502X
fe16gfRLJ6GKruie5eWPTn67DJjgAazpE37WB4OH2yN/7mbk2mBsaYX/fnes
e1FYsgCX7+5MMTalzf01QnUmweLWKnErBOakdec4FPZ296yQJxKTgIlKI9qu
n/nFheSNzskYVoH+EXA1NdJpNgnmn2NRQmoJ9naUybisTS33eY6eukghzgTO
Gjkk2fHeS574bQlCAoIZ4oq1x0/T/lhFntPwm0vr/Ter9r3pvnCSaa/T5/2T
IObcjMphL7h2l0Ky9I/eYqSaah/rtzrCcHsHpugbl3P2DndDAfeleOZ3wZn+
yz3xJcoGDRuk20MrP8uHGMIjQj7W9kRryVKNh/YXMx3tEdQofubyE0qLdbVi
F4mqnDuwWWjm5IaX012qScY4hD40HYIG4JjPZcelH0X9AqCHvrpXJfq1ckfQ
aN48kX+H9loc1hoBOW39K0AsafW8LQwsR2PwsK4f6/wfa50V+7DiZMkW3SJE
AADZq/99mNgHmej9gmderlgqjlS1bLrgTwrrux5JREyk4Df+bRI2fFBF74cZ
WUcgdl5FW0hVRyPGbso1ml9gBs4lEKyX7Ht5SO27yk9WYSZNlhg8wc81Gu6J
kll+KkTTJOHEY6yQQmg7DfISHCBbkbUc6wS8eE0YwK0yJuyr/uRUTwUnAX+h
Etzin7IuT7mEoM7XV2R9HNUXQDLu/YuLDr7auPyJtCJN7xe6ecWtYpOTby55
AjErw8OjpwTU9LgJfHdKWW/3+bgQplVfR51b2A69B0j2L1xHoVk2OHdjcN/C
07VtCeia+ATd8zlf9fXTqxQCkF1QU1lhoq30PWg2DlF6/WMEQHHIR5EsIgFs
RJvkOv/g6XHB1P0IJZ/qmBOBCzye+qMF5afjj+1TrfU/t4xD1iT/OKwzFNHg
/o9WGtMj3QQ4tJOPL8UjElGEXt7d+nOGM1gltCd2Tu9ive7OqvIqfz2ePs/S
YbeVS7kBlG8KNe2i6axT1ALL8pBQNC3CHU7BS6un7743ZpyGNCqwl13plZf7
/WNvYE7VuB3L1neqmd2MCvUmZhptwYtMYK9waYcm9HSXuX2btCqT5zeb2Xh9
1oC9snnVMScDU/A6AAkhX9KfubMB+eZ54IAaCkLHb5jA2Ei9MUDyW0vZJW6A
4b5cJcRWuouw1D2vOt/Rs/BR12vcOBySA1u0ShERSwEX5iKaKo+DwZ75QLp5
r4jnShd6pioqkpz0SOGDYlYWkQ1SS6rwLQeRK+hoE4ZsR4d8orpY/odUxYfb
epItDF4ElzcGO91oA/o5KsJ2kIHZ9DEh736Yu6JTpr8kr3P+PgMZKudY9AzK
aV0d5g3hryYVCsdgp8sC31TxUBNVclyYr+GyV5BJLTOJPzRa/y0rpQrhY8QF
p0gVy7Fuhe5eMfodD/rUzPlaHNFWlBqo4N9YIhoPIMHsaV2JgVBxFjguiLOt
MHXVL+G+OGGSXF1mkrsluJ89zFSHoeV4FgqEW7+V2BH6e7DSjORq9fXwaZIj
AfG7nTz2o5xQR7fLBjKBDOFNEJKvlO35UMZeqlxwW+QTjygE9IbzeVnseS0q
d1wztPufQ1nuDdm88x7CBhLrCE8R9SQOzPYWF/zP20DDbsCCWJU5/7xVJ18c
VeCWbk48rLOOcvwWtssbFPszeDFon0i+jncj+KbpV78z4dF67zd0k1MDli+o
ItTbJDiQB1nD1Sno0bYycE1izlePmOUaJaAVXqieA8E5AK1LSJwq4s1fyhZS
oEFm6LjX1oZeyI6GqmzKrtnK9m3EvrL2um3jXEcol+NlFsCanm0X53Yq/hy5
pLqhSAPW7ZjqqdSJ3h7UBBfi/oaOd90M7/YTC/uBFqfd+uk+G5hPfZkIFiAt
GMM9Fiw5GPyvdbtVO6CxHFAgtweiLm7/BIYVgDvkfeBWAzCc142HFHYByL+H
I4v1joKwOt0tQnMeXXo3XOiak63w8/TzA5BW3HOPlT6VjJ+8Wa7pAuZ7N7jD
R3etQsJIzATIOi1IZZ7vrTaCkztEh5SBdCJQTCim7tcSt9/Lp6mgvTOv6Xo+
VpklGgB9nLf/6J7IW+WiKm3kE8zuOfm5D+MveoCCgX0yZ9579B2daOXzu11a
lf+uRlNzgrJwFschtFGJE3K8kOLJJ2syJeRDsv4mqVZFogsNYVM6ylHS6sdj
2yRsinMJgbyJvm3eRAe0xVFARhaGBhi/efXJXg4W1/C8xahe4SLcaQwskXvX
xmxCMG+idZYTro7QwzqavXZgGdjuB4F8acB2iWKinTiY3V77SaGayHZLujY9
rUeoK7ZPK/uYBOvT2JnjYegdQeconT/98vqtxijaGFRNVw3kiOU39Hc9sgxS
u8XXQokKLByG6lh548rCtMhdixBN6hlyzfQHrq+mdYocsk6V9s3lgO5/Oi1v
jgmV0zJTaBaeUtVxia24m4fqJsnkrGkv65SfGc5KR+hqnI7Gvdr05gShekXY
6jFHHuaRpVEJIj09BemLxWn7HZrX8CCPA6AYmguIxJ9jZU74KEn78slIFkcL
TDWp9EOjkG+nNyf3w49DGwPv8uuxLXFV7/pOpwA7Aql2fXmFpotBONlTo88Q
fNXyvu4YYF0w5y78JOvbQvFef+esNLkp2UV6H/DtFwglU7EAvEr8SFZBaLu6
ihkwLc9tgpitZ98vs+L5knDcXQEHh9jnwUga/Mk64IDWYuC32CSAarRjz7Vh
HmJtU3uanfRpbTqWCNszecmKLyq1dh2/RXGdLXYLRCOANhJOVbpXU31UV5IT
DqJMuaPl8m3zZDcj9zk2TbDomAEn8n1XZtG3p9GMcmKwNVjWvozUFSV3Znuz
LWN9JqOT85Gg6eiMvFg4tz54Vl9vUfbocNTXjCzoOhdXdrEg4oV998GGZkHH
V/fXhlqXU0fDUmz3vxj74MgfnPYN7SiqkXnxgwCY+luOSBwuSd0cGCI5itQy
KP6HMPtn2E63NsKKCpMr5EMpGsCi92ihwtU0flMbmghx7iPEtgvI5mZM/VNN
dywtNnq7eSupeT785S3Vl5fnHKREVSkym1lnJ26jb3hnnrw8ye0TA+d77aMh
VYhnT2dQOFpiGQ17K08yv3ktiVD5t0hmkiLUtlBHWTXKXhS59LDSv1vUq588
Ng9URwf64v6OJTXHWr0OvmwPeyMc7r5aNT7x2AmD8HvIP7eGgmcWyEdcEHbG
c8bQwoEhZMuPk5ygijw0SIB99nSNL99MXdmSf+Oxh4AIPJZiwhhZLuBAnfyI
4UCA3JkFMkOzGa29JqwelEJ4vrQJ4h/KyjJBu81SkC0Fo7/41H9ZNYKxWFdm
TECuspXi2aZW3dMKtEVl7oOxRpacY+EDU8eiN1XV53kH0TvJW/gOSJc65d7h
gR/93A/JHxgxlAhEKRd3aiYOOzRc0x8ZTkakWl/6Hnl9eda+6PVc/27aD8g8
cYWRSWp4kbx/hPEllXs5C+5JNQCe4SH8FKO0jmyiHRDMqgz+79Ez9VgmismT
q9hFVJ8FQ/zpaK/AL3B3sIYMLBMSUguB9zIdtjwgWo3dO7Y7cURUs97GypxL
Jtd1rqRZoYwoFOl6w7B0WFjwnbhialSOOYaLL1mTqmPm3gBA7ZsW+0nlKSLp
HV4dI0C0ZFfl3xyA74ll+CdXZKZ/tZ+5MSc5tUKZD40x5yBimw+1D59KRiEv
nhPRTj/kL8WMPsl7bAHsk9eV0QsprmCi2iqaJR94v3nk/0mEcbxidaFLa3MW
siLvM3tMYKJsARJ4lKsX3Tge3gsM5WK0SV/lDdBSYdHDIH+qCB5AIN90Nn96
1lQApyI2Gti+V7wya2Pw3N+wosDnpR8K2XJoZz7LXquma2sWGGzOPxmQpihw
Lb66ynR2LmLMHZX76MOJn+i8IcfRu8SwYyzWVE4slH5an5iELBEXuZrI8hdf
ZmSBpSuYwuaSifXyFRUxb/S8xHXIk/7cW4/9vqAX+JN++dgD5mbEHnRAqndD
lDbYSan5CW6uYSKbYfIpfQXhWgH42mAgpb/kTf+rjLTS7NBi1WIxMpNmC2Q5
z/I1gk0jRyoRJ+NekTeuL08O3+MUAJjwQmcUu+NcCM8pVZqnjEV1x0Imwysz
IaszFzlINb6Lrh/jPVybKM9Ai4fWHzCPNpZMz0orKcfIDvLbtkBAyMeyW2Y6
ISzf4TAyp4SUOgy4d6Doj3+iiDziOTzfw41Bc1Bds9okzxSMPohweqK4k9Dd
wlcGBaeC0l9ZKxztibnS2QD/7V8DZebV1dnCBX/bamZ+eqQiBqb3P94WzcAN
3+cnWIT7Dopp7o+sNYJZbFGKIMJB2AaeVaG7HTzOicrKBLn6Jsn/Jd2jGjqI
YNO2pAUSFqf0/lderR3P3+JaPbPLCC0yYOpDVaHfw1b3VV3OpQWkOV+ChUoU
7dL0+o2DrYM6hpHE6vavqGmMsMgMAEdelZ6mAKiKmPIFxUsTSF9JooasFBoe
cKkEMZCQeoExQl72iCv9PUe+OMxNinXTCW7cZvdLlTKJIIGd2CZh33kjQymF
/klGGz1A2kWfAWsF3n4Z8NdAs1FKjrWTv+I8fxNAdXFtRlCt3mtYD4udl9Qk
WhiEGw/WY1du/j0hSuqI7WCporuQ84oT6LfT5g0yzqFx0k5woAEardLJDrUw
El9ERSnIGCMlzDNrJAnnzectxuJ7wS6gBPEGV+XPTXQ5iU7gk5htwCBScR0S
L4h8GTwac+2eq2XBAghLTHLDLxWSOEZ8ZhcoqcbBmLJ0ThQHPTijDjIpmzOM
c9EQA3xzn8RwXVIJkq3krppr5Hc3glA15F1B/LvbuWXlgTOdkwiVDiBmv4zp
m5Y1S7xwV1qy+6Yz4K2qtIhsYPSab12TebcA+2UxivfSvSOkFntBcqZGD3U6
YfV8Pv5jb7yX+p67Sx59KrRyXnqoxGTFeQgkWpAiZx6sEks3YryODWBrAHBa
hPB4XnlpJKLd17EJC/J4CxhYhNfs4GY6Mln7U5oHvxDbZxEvz68QG5h6W+lB
6MkqGgChVp7ETo8Qp5tbRWZOspnVfS46VkBv85UYZ7nNAe9eMygcif49/6dG
hR5DG1tVrBAdChPbQwgZXVyr0IwlCUZ1DxnV5RRCwy/xYRabPgZ4yJ0JFdCy
ZLapM3ci148QbCSmGner1/VKEk24jHvl4XnvVDZyXxLTGRcdy1k68ao3uqAh
LG7ffp2b09Y2gT866j+4ucaV7CzDEhMAHwFP/9Li68jjkdnQmBREhLeVdGNP
xyADcv7tq70elkfaMemHiba0l7u9c1a8mHczDBaWrSyJ1OJorko8dto1zCpf
Ta4IxJ0w2dJ0TxH9N5/+iyP650XbuHd4bCD3WInrxJW9rEuUV4k8gKwhq9cX
VaNaQP3aF9Oaovk2ZY2hJi66NOfsD9JX85g+6yYRtzR5ftUWcabRGSjGiEvr
ggajOm8fkHRW8X/qQGCTVQS/SMgBxItYBDvplaka7ov6LLpyz3sggzr8Q8GR
NBKPLVNX9ohZ03cunB53YIUGL+xvsQGgxiPNGleLLaPV6i9nyvxlEYuw8GBS
7UNwauHSSei1EksmBLJeT7+Zf/8ZDVQKWpGEaWjRcjAHZoVLKx6tvVN5j+eW
JEe3/bwJ3RJtYCzhpIBoGJ6xOGs/lBn4PESf8gvTwmM/EYo7KonA3DxdSRtO
lfKU8gmc4Wi2zjBSYAkk3WEVmMVopQKr05c3SoWnAv1D+avyj1/L8m89Kao4
yXB+Wc6phXcdnttyn9FNoPcAJDbvkt95H3ap0zIt5r4bOIvoLXSMXmT2wDAB
z4vGCw1PQLySooPO5f01s3H5eVr5ErcewFt4z7QSGAbqy4BCms1FFJaWIWOc
kVEFWmrLoFVO9Kzj6PheaPJuYnWL9V0XWq6/7FbbdzkFfE3oG+O1sfGQOW0o
IFd3GvfRTcOHhOj+Zr9N++YF9biWjXkKXqNkXifEkghJZC5O8fVqrpl23UtU
bq5wrdmJ6KKuwihY2EZ4KVwJKCkfKwJKaVNaZ/IhQF/7gakWs3IRgO6GQC52
Q7BiKZi7RYxW3QnA+tfSE5MafDShUgWPNceGrfezYLSZ+mWekYkyNQqV3s2c
yyiW9hRIXgQ/EeRSgdSkU80JB1ZruyM9QONtdWZ02O+wG5S2DKs9exHQ0Uer
f1Up1zO0mSF5yfSyG6v4mZFu67eTrTugz5FSkbqe8dZwbPat1cxshBShHFrv
nC6qOGb57IHBwhcFeXb/gsyvRuoj//SXo4lRSgDaBfalU7wsEFK7JmZi3IUD
vd6nkmlrkEVp0DjDNveFnIMdKrUqRaSVxmkcLKHnW5heAF6R5SA0sgaAwAe2
G3blm+y4iBTgAhOxrQ4LF837bkID+M3vi69yALfblp5YZJclR2Hw8cnRGCFG
U6w5s3WYxzTyxSJiBJFQTB+Dh9fRYT5P/0P3O+BLVcwGU11NJDRLjVSNVftC
cMTZc4Dm7yum+uzlpUuxs+6TwJV8ppvWeQX5O1QyWuchC2YyO4UjAMcXd6gz
HJd92ltVDq349zj4J2UHGeIkgzlsziuxaFOqi9kkTk7K0V55hz1M7V1UkLC9
iUuS45bbzGCqi/8SY6geBRDrHynzSuGbqbNIBnWvEsdUB1zwfjou8sHY1G2o
Pu5luAbAztzYpReOaC7D+xBoqr+DzjN95YlUWHx5K+PdYIp/XFKKgYEuoLts
cZZCRs51kyM5jB9fdyqPwh9JadowUPhpMs9x9YVcrC/a/oEgVvJ6WmRmKX02
VDO2lWqcHPizBqL3FHQJtSkfBjRg++tTwoWLzJ31YnV7DMbCwcsQnQLHyPHI
TLbzy8/rLJN4SaP2Dct4J/vvUFtkfP69RUY97ciDLjlkOUzVUgrAdjOfPfj7
kCATNCrlIFwePF3JV8gCpUwuMqjR6YrTwqbIalOf6kFTDGKklSfg7221GYPP
IhiqTU7Xrz+r/eQ3dfaSOxtM3KmZkEUWy5r3rV5MMOiaVY+8aNeZPSWNmOXt
5EvlfivN09Hnh7KglI1lWk1SP9buSZoRi2oro3iRMOtAhYsd2nE9Z/Cwsy+l
lUnaqU319El6gkRJe2eGWDIV/EISwLLELLfdJUmGHPLNPrY6C4QpZMcyoT3z
utvPEkeqLKZwGuCPolNIIKzmyZaiLfNkvwMOGUX4ZtpYnsvqd3te6WaEuZxN
QkiDl8nNAcl3q9mtef0npiDcBwj9uSQjo4OBdlBB4UXu2W0t4kklbTMvW4ar
6NtmhqpTEkZKSmWb667/lzY1oOBqHb47HqmS6gdptGrTG8buHk5COTrEJaYe
N15ODR4sZGw9hZVQr6vC77nwNZ4Ngta11RWbFqGLIoLk+JqigZKbJ0FZAftY
R9/zmw5dQcoUwy4hP7qEomXXwuoOZZROK3jgLK+gbzljvL1ANEnXgzma9n+a
ZKgGz9H1HSfTiwNyLjZzv5AXsVEg4ZRiJx2u5+kQjoSAqc3iaxtlPlcSXS3v
3NIeA8QSvZDG2ISOm+IXeynejOtPdLoJRnYl94utwNs0hKsWfVx9yv0KVeMX
RM03Bn+UZDPLM+MSkxyzia/cDfsiy4I5lr8xwv3xv80Q0uKWmyGNXmSjtv8n
g5nM7IG87hRw0/ldbtxF2um/83feQbXDmWVjeKSM2ju27gLYMwTLReoFzHLB
cYliyaQiy48ZLim+q9CirM5zdXPesYtCjRjZojIO3qoozfr8QfJD8K6xTGlw
QS2X07IFz36hXbgyvKwGdha0XmTj0tdELvBVEKP3jriWJKMA4ZVao477Z1oy
SZ3Nb+PSCCbNKTc/E2vL4//27xbIndM107+p1QD6nxmbynl6aKaGNp4k1qHE
WKiPy4lddCivDozCHr7puG8YBF/vuq00jNKV5PGW2aML+R08h4hdB/PvQoVu
MOOt1JHpvsoSkQDtOFW4av6CVbHoqZfAxNhwfrH3OiOhkwfqCPjTfTiL8YWb
rNOh8yBFsc30PYngkDcfTe/MI6WbVkDOAZSPtmrUy4aFHgTiVLy5kPBRNcf8
LxidfHh49a2Y3nMaZ7xf2YGOt6h/f/+F8cWzcwLiBoKZIyOZx9i0LjQe67Z0
OtQLcanxCFGViB2G2XBRyH4VrVyiMXluN2MaGWyeGUvBXkDnWaxw0sg4sRk6
1E3RA8q6xwoeApccJKp/lbiP0Kcjxb6Evw/zqHaOs1tmWjB99ZgM+S9Sa0/f
5mSt8y+Jy5g5B1qNP4VhY7DoPfavjhB68NHdW/Mjby2rqom2fL+svxyKsrYL
37qm3HnMRdBT2/WINGmEJM0khPy6F5275QCZtJhKxdwrI22x733eCYKLEOvU
zvAZTHDWKL3rp06TyordiOevFb96oMPTLebEQvfYXLAoKOUBvgus0xJd1qFI
oBxAiShc18h+lnx8SqXITaTaR2BV9IY54kdCbkVnJmP2CWRzaSaDJHbzQHdf
jbYpqBWadqiCsj17CJOgAp08zxCTzIhGHlc+IxEiFXNt9rmQksYj/B/seg55
AH+93TmZqKfYn/BzeZQQwEAneFHIyq5DLvDvT9ipo7liQ1PhlqNQSL3gqeT/
PEIS0Huz8TujazoEGsQjWWBUQZzgKviIF0A9LRR8I9QtS9id0643reSgYtuG
Hhr9tKWr+PlcdhYxBFay8xpJ7b/u3qGYtBTVqWG5FnVSV7lGuXlag9y56fYI
mQpAl/lU7bAqMoo5oG8gWKqnrpgs6SnpdR0+c4Ydqkq91OOS8iuQo9FX0PIx
maFCaUKOjgwtQfxCWECAST8GvtuL+1MGZjWuZUFYSSsY5YcMB6XGLlzcjmlu
zYrBbXggfDJlMrOHTgWa6ZIzfU5HggWEqn0Enzj9HtdVuRfElSNi++bRQmMo
tSnu6muJ4vj8abO9W5jL5J/aBf8zMNaXA+UXuR5viYWOK1BBtZ0khJA2aNXc
oAdi9VCbxolwh35HjV6VC0ErVm/7sj2wtDyJmjQqxN/C7yZsjYl0YPwZ2YV2
PvZLFNx0veK+gpqKJsAoY2ECzNpELrIsUqB+MV4Bc9H/uFcdaedsf6SuHvdn
ahbFbiCkP+nxSxMaMzLXDHS8F40wsZV5Zssc6xDj6ZKaXyCiXUYvGWOV8NER
ayg+N+l5+IeK2AXHvnZxsgUvRkUvrFNAIrpVnUM7Y0JzOPCd60lveTvrixWX
58w4RYJuTtyOSmZHLLPXGL/PSamnek87xIEylslQNjMDFj6UJEYQr2ZmVN4Y
0uCni+grVWhdQkCf/uQFV223gz1+HIcOvYyLRg9lHU7kr6NZgW5bf07qdghW
hxaWzR5FpskpYsOXN202oXTshLeaiGJRamZvOhmOKSdqm2x+1CjeLCcg7AXr
2znPODv2elXCJNq38xq62Ch7e1c8DYQ/pqZe+K4Rli+UoJLEBy3fm8RAor+1
RqgegHtmEwbtBCvRApHHe22vHNGbAiDrIlF4bA0tmxQ0uOvn5Xfdg40HtdGA
y5OUj98CJM1Q8vWjIktH4/IIOTHx2Us8vTZ/hNd+7QqtroeyLQq5pP7Bz+/f
TCAam0gSewX36JA7xYgFueCfcyLxYCUDHFsPeWLnwT0i1+TbOfCZA3hVx2Kz
knbEYWr6nE99aKXt898ezsNnvS3MU4LQzyIx/+0Za2VlMcsYDojRtkZf542I
Pv1hHtFAgOVBehj06J1jiBZAhhVcf9Kd6nTPZUjNuR7ZlUApq5m6Os7oXf2M
NRJjdQUNLBlDDGpQJwYHgXlHkOs7R3pwLmWDyoutTjHWH9JWFKy1ggvFj9+s
F6wBve5HcHQZ8wyRSzcQmZxtERB0VMkBuAgBSQBSJ2AZ8gk2WDebMKcdok9d
TkbsBoiOg9oRYrWhiH3Bv9+l9DjMw2qcckJYsQ2m7kKyC3xDWCSK2Ws/Wkq6
tzcIi/jFc+hbnfQmBM87+keOwDYC9En9RRpQGPaO3Kqgeizb77RV8uqtriKP
wIpxOyqEyKJJZkIHQz4UvAj4KhPBfUPRftNGw1ktFAhiTfkkXOdC4sd4+UT+
KCL6HoxZc+okVFWkI2IEs6/E42KYOS8j/wUEIhmDY8tC7/VaSqhH0MwC7HVH
tSpVP5YmMZj1IRiKV+iHilgIx7hIuNzg2g75DxmBJZEyT4QifRdn9PHi6iZG
TdYAYOPotsfbmez15CkcPVMNl2Db1IhLpcqrU85/gpvXnW9B8/ICwm1Y+O2o
6t2lDi+UWWr/aEYwSDqouVliiXE3PwlWTf9SrrFC4RCF4nZZmisYkcKLmObs
fvpOiricZWurhFLAHCO/pq5SXIs+2JKoXf+IT3JmfuV4rGJKCBZy0NNW7o3g
4u/6TH7GaYEfOxChxSmnP7L+jO6Sju9m9ilVlMYMMR562GzFvAjkgqa43QY3
q/RMzMTFRTWQfJHYB1bClviAC166ZNFl8chLSRHZxEFz57jJ3mB33DVEbqpi
QwPV0ktYiF9XXVoVI5snjsbqF/Zf8We8ulQlcvSROCNO48An4KWkzIIr3hRB
AcEERdhK5i4DQCjiKe4LGpnUCVrkalVOqLj1+Whwj2UqucjhgJa6SOu158Dk
W6GNjoBo4bfXzX9mqZXv89JqyBbZkVelgEGjCwFKfaiBTHl+h+D4v4qq7rqz
ESHXCTH6XfKwZEWnUUsNAK9W41mC4gNmFSjnpIQfLbcX5XoyL5Xb8FkMNtVl
oIBAWgR8sPbbdof7ReBiMRp0QmCZV/RwEcR/HQEKd7hUhrk/BXrvd4mvC4cf
dfoGRl7ZUDwKniYGrSDm4xfJFWM7s7bGpeVuu9xPSEAKFyVa9nH+mWfc3HDB
hfXkoLJ8SifsbXGID2N39WJaUEFd25SYcXEL13tuFiMOKo3tsmt7PupXC1Rg
FtoG4aYdaTnHII0o5b6QWJd+UCuwJYowLywFG6qzqAMkqG0KRrcbqUEzOwxt
4zpl+nYt37FgGPfL1ibSyc4hllV53iyqG7FDBzwLMQh8xcnFvi/5hw5cV5wt
cwu5cXmA8tMPCdXKypO9bE+6R9KZL7BE+k7BB1QsNa4ZXAWCp1jE37VQxxqc
pFPCZVry+meB8mY89LOAHOmzGPrpLMstOYwFKuoExlO+/jKkzTsZtMtpefL+
EVxihTk4ybhioB1Qa6FclxqAUkb1IyWNWb00C7g6COe+g/kZqNGoSAOMq+O9
b6G+zVa4L2KCgbFwS1JCPB4E3wqDkm4Gqyv3pB2Ge037S/eDQQQ6bM9hwG/A
OYNvRW3ccG6mxPDXwhqqiDaeYu8rtmhEbnQhozPW/H8DcrHVjY9nabitv/sO
9/g4sk/cOCJ9ZUN0AWUICe1QlfSUOhF3nt72m1MKNOOe4thEQzWkLjutHezs
x+3O+1/wrLkG4xJZWE7UO5PVBqCSgL5u9ik20N2A7TBDUJW4/X5kQXup+vSd
NDXygKJvJq5v1fAM6lO4Pj/p9tBgDO/7xJSV60ue5mFMB91s0SjLJDzCekYE
GpJT7mQ/c20ezrhF6EOMuxAnodIuUzuIxm50yYwhwqbsU8YcXkSzYY36NwbW
vNRjoVItyikZexpXIH94Eowb/XgOrR6jiMul8RQjgm+BIOfg4i4Kg1wQSX11
kmAzvK/iOSvRh7oinBBtOxrMOOjb/62qaH4l7Ek/3DHsB5/Q78nMSfON5RPH
exQXL1jTrgVB7+HjqsAdsCGqgBGIPKt57m019Jsyjhwn7wVWfT0DmPH3YvE7
cPUHswNGolzweYE6VsDcunJ95SCVE31jdZqnS3LTgKl+ia3dYBvLVYPe2uIL
M3JaW2wOCyR9p3lNs8mHnt5W6NTOgqu8WVurrDg8TTeXtoWsoS34eP7DZrtW
qHEdvr96vfURkwy3DyxJS4TcSJn6wvoKtZoIo5gfeyPNKwtdNta9S1EEPo0Z
YljdXnEd0Fp2IG6keNa0yXxmMrbctKlkGFQeN5oIrbyoYQy5l1HPBkvoOjLt
wJifW5Q/sn2PxShzn5b+fzajfzh/4gFdCiQxFFWE2f0P6JqdUaB9APfRzVng
ZtXynJRaIS9KSpdBNfWXqTNU4PQkM6W396tgqxAv3VTAY00OfqG6UBvjI9Ze
sytQE/QKze4YqqW3eE+aT+PWMqJg7eZO+VVAQhlcUomSZSmD8niMEAUogDk1
/y4EwTwvYpjKqnBYPKUyGVzv2iaKXJ8mIDALNrjcowecfY9jq2DLa6LsnmdT
+eu7dxnDX/Kl9R5jMJT3JwdDK5N1S8MMrUK4Ce4t3ejp++kzMlVOnVkQgOFj
h6NKwDmkVpt7ErpEZ5pJFVb9LJJIt+29HyfkPCoCqUIPub0e29XOoxIXZISC
RrHwqJfmIqajsFp8n5NRl/aYaYXsZ9mhCWULOS2OrswggKwKEZrewSBH5owi
JAP53hdrCJjbHbYjLFesvw29Jw9gOmbam4oIBFtAr/QWXfadRGDgNhWVmpL9
Fm91BxXoUN42HuQNvf5FbeMdq32U/Gklte3SGs91SrsiYz6ud+XFa8qQXso0
8W5ktno7FAMO0Ydcw4OyzYqI0h58Vazzmeqt3QtH6vAfAByBIebMTeiBY7gT
ib7w8E6kn5aXgRAdxL7FxKQTIngZYzERE/G6AdWnnfCJJg5I/VM/HttA7eLW
QiV1EHhKszZp3f9E5GmikycJUlOmYJMLYfCKdVsvv4WyR15TlnHsLwlDP/Dw
gdvZeHAOBs07fhEvngGIWGyILvLDXvykLNoSOGhzLvR0gj1Ne18i+j8bIjlc
n1gt57uEP++SO5URco3c7i4VcVGm3O0DWS5Um1XJUwSvGnT03sDOKQFjkKyi
juplrltfTkSqNGzh5EOO/V3l4/TBNIIoQoTlKF6fj9tZ2OhuzFh/ezqW8XVi
nXIP3MeRLMl2M5DdbPMzqaeKCCC81CTKirKAaiVtKZqeh2DFDNssNnO1MhbS
/IfCn+WsfeTOBzA+t2EKoKNH+3hYxT6vufhVhUCoAULqcKQTiqTEcA/tvsnq
iBj1tVZt/LOVigchL5XWzWcDTHlpak69Kl3Ihp3ihMhH9rBRenUDYubKYskk
XjDyJj+hI5OukmNG0rWjRy0+yuV9KB62wsJnd3ypr9BLT5kAw5kQpVXazNBB
g4MMpp0dkNMHt9AMjOpQcCWpBEBaPl7P5MUEiMVSHSMdDqQ49d9dQfPjNCbU
eZuuUlvr0d8q00nS04g9eF/4qoqxe33uIWqDy5W4jAGVjfzzr7CTvkFpUmbq
QNIaXKWLqkzJl6q08IuMn9EbkSEbPCM/wBwlpZMyzIQqQcHTvaJtUHHmEz7s
1IyaclMwi3k6nolyfsS1y7zKisEga/C6WnjFVCdOwaWsxTh5mcVTFSa43kh3
diLxSLDCVNfpIpRf71jlV4VWzmEbWXHuhf2+x1EsjphIm0Wt4wAQd4HpYS8a
Y2LDipadDFL8l/RmK8ZKom4y81WBY2ekIdvKlx55uG/rsUmHkvEgmSzLPoOw
mQ/Hb9zgeXDp5WlJeFo0eqeefzt7jkX3CDoU9wG+1cXh7+IkQemyezJlpAaB
AB08TetyaSkT4q18zEdhwVeuH3XHJIpIepPsmRd/mGxNsiXvfUE84AXwu9zH
I8to61w7C9DqDPZxHNRF65DkUypfvHAMpSa7VOpeQZsd24/+1s5oZRR9Moj/
kpMxKeGxX8eNsJYZHGxKOrNE7686mtijir1MBdxTCi38ZZPc1py95UHnpwOX
aSsUPAVSk/+4k0E53nBY5PxqU9NTRqRdB6D5Ko3fsnVsAxxYCZI38Og3Eec2
aN7pZhgvGcLMsAzaNduAYiAQ4ZtIRnEzO51F5G+/wDueL96IrOogT2zMF7kE
l1ZBH/ellSoXZpTVymKpcu9cWUED1D9SPwJ24nIZz2n387yqpUgIFXbSswF2
ucAzSfilxiZ0/Y6LiEMVviWgiMK6COMiurEC2fb0aVy+0XbYPnAL1eXR3DNM
V5TaE51UWxQZLspyQMY5ZwKrp36faVhHPKm8C9A7txYfiOC4hNbzuKUlTxnq
9g1qlWVZ4wPKw/yEuUugB/qQR05uFye+o1dI75a6TJCd/s/qRTY/nQ/dYAn8
pfMhMzmMBHvH7pdqEd/EZPBfxGzcUZjqtsm7uL3qAEQvTGyvYCtw7D2NQNlC
6por7CcvqbX2q6ZoBeWQmw2d1cDowNeD7gYTws4wT1vHs7XW+1kKcReR3x4K
KHVoqGcWjeUOdvKMjI2npg6Eu2YnP7KsmPaGh9pT7pUkkzndCQat4oXcf6Qo
QeLIRGwEqzG7Zg8uLn3yKhMg2ugb1yT3UamCWK09UsQ9XW2rsAg7ij8xQzGf
RYCdyzUJN+MzYOA2oRkTrWH0FLCyb9TxVjaBtvnKhSY5kCDyfOX5pfxhEBwM
QyzlsvT/aej1uCFaYZ6tXJRqhE7CHYyGyNHLO1Lg6oF7ABTQdZAX6SXa7teq
zQc7WUusN1Xc7+IoQw5CPSqiZ8Hn3T9WK3dfufyv4sEWpDQnUWs/xUaRSVnT
tKfJuTa4fLYpac5mFgNpqjNMpzW4V7fmyP5xFBfJztS7rfsM1l5ay6xl/1Ju
TNf2JWEIHwsVzIZXJEG1f0o0bJZkm+b4UyZslCcGH24W1hMS+Rv6irostAXm
oDuckrmWQ6gzoO5kRqiz2DhYrgDnPH+GMfNha5gQ8gPY81kQsrEyJLmiJMBq
lxoJbcimUASBWrMcgALmaon/6Lctcn6f2UYgbClXp7u8NMhukwo1JNSfHU/Q
bYWnkfLm8sshcOMe5QNLCWT+eiNy6MqXuIWb8RzQp7mkdW5GbGu3InYruzq+
+vXLA+Jcy4EvTwpc+93C/cP/T1aZHsvLbMmgaiybKRkbzRrxecRSUMlf/LPd
SCbn8NnJoOG3OHz6AQ+n2RgQrc6zJ63Lmq4ieGPHdM1SsItDZ/a0YDRS5TZd
fSzp8wM1xGnX4Szn8c456ClJOGxsV6kQU38HRzK+xeuI7KFkwQ1qGIDAebhA
sSF7M9xiEJT8K8LQF1jJ3DfdLmcpVED9ZbAx5yOYBeYfBRmjeenN7xzjBJfM
oO5xp0oGY3DfesXOAP5yMLvHxQdxvTiEKhE5qPb8R53f4sWn2WW9/b1fxEgP
I9pwFqd6nrpBi+hhJXEcDnRp+TqKn5W32p0BGibVnkru4feeFL/HzEJkPLSY
H6egWW0Nt+3OCWvKEjJpJFG2kUSIexwhM0jMMtNxgOMMS73T8jr/JS2cL/Qy
IOj7nf4u+zC2xDhjFMb3jd0D5QiQx47Ud9Hv9N8ROF2T9sqEsEXBFTAr0li3
4JZN9868JIXUnHQAVjS8HO+llgHmPc4uo5Pi0vWhOJqbC3e89ZBjQq0PvbjC
dr2NeNPrQw2Ha5Mv0rUVo3mnx/iXuqpl+nDZ1RmoWUXYMdW3gvHzdzB2vHba
xlyjpjcgKmqBNKONDfQGbxnIXuP79GVIOch6XV9TJRfWP1ezXs3LX+VnPmgS
FlGXEtCCSXyCZRRWtqRb7/SXNFqcMmZw6NyeWQvJ/MPRe6J54NS8OugQcxLm
//qxhjRIFZ5cEiu0lFp2NKCarKBS95Z20JohbaT07fIb1/e99A++gxA6tRF9
+Ma1MOtmfVG2obKQEIJvVE1eX2mNsTjHK+gbJbhY1yUxJemxNz15pedSLn1x
O2+46IB8M3B7ENUrBTvNJp/Q1JQnhR0inBw3t9bgY+nCIToKqc1yNlaGCQTI
gw4LDm8qyVPayf9cjcFaqzLwklSbxbS10D0GmGyKn9vAC6PbRIVoAobRmynl
ypAgqG5Nl0fmewfMtp54m32eEpWEh+bZKAtdSEopY3s26ksgTGTEeuVd0PGV
DFdaLnK4JBKn2suTf3vjS31nIJYjlukJpOFYao2FkKrnRbBekIY5hwjixrQ5
c/BJn3rbALAZCKAHlCPVknsGUVXxyiIMpv0fbbCzl5z6qws1KwnvmDVpF3JW
GlS2DHPUMtEFyPGtiWXET8VYOqU0R5rjxs+UlgB1loN/hm8MojXcVkAa22Ps
qRp6NLBaLsiBXaBduwo/Id+sW5ZzUiVsFigbva3+jCiyAcEFhH7mSduyHNYN
p+XG8YxZOZvK7hx/FofzPpQPL//Azewd5L/HXvW5DNQ/crQt7qbQFAy6xKBo
r21xg4z+nFVmWoSKI3gFeDegs54NgE9IsCJs8+p7MNiotJpPJI2/TcuoUmtl
cIkEN1yz6Zbh4ns1Lgt8+AfOaF5FgvRp3AFQUI6BC+5t0VLXndBChdi0jEhh
sLR2MxKK7Wbj1ELritYuFeZ1Pg4kWyJPyOdKf6bIOxAB3Z3SLEFo2jG0zCHA
GPyYsjxT4ENkQu98E8/wXoPuIlFeJ23WV1Hz9sVtLY9WDpm6mZLI+sYozF4/
TGjbxgqwD016pOUYMoDNqR2YpQaolxlbVHZ0qCMqpdvhEaHxIHhPzhrVBQ7G
IbJ+VPqvkKflIiAHjIeBnshXNBgPhjJewYEcufy79G1KgLD+7EzgK/ZfRdTW
nrXqPbeg4QQVa0oj//KLf/me9rewm8DFRo62g/ehU5UeAxQPhjAh9hFHdzam
oJUcuY0Lq8m0gsP29aE6d61w0MU9wb95Ir5YJywz1z/pPZLdPvXMdecbRpAB
2v6naq5qHE6O/KqUbOsSTwr4S7hXJVv8kQbfVoMCpsYLPAL+/n2rQGl6IXr+
H791um3wIWjaw3kO0EpogPeUad86z5Gj+2McEXx9AWhQrdo5LI0xcrPEjncv
dC6Rv6OAw4gTXoxl6J85D0ZPX32cZT4JTovbCBr/X4f15bUzdUWnufpoQDPr
WNFr8pF5fg7o2g0NjOPsa4u7orR1kmJultZkksmDe2GQKipqqcfUcXcY0CJK
qkdl5A7SJyqaknrl2rdifDPjgJOSjbzii25aCnnJbXqvJdHPPOrgvnazK9N9
1K3o4XXuSI/0OKLdMiyD4tj95jGbV2tpt1tqvfoUiiR/me/7NMmW+o78pWuK
2c0bxFW+ns0yJoltouYz26LIQpWue8KAbFOVSbwUHFMXXbo3L7zxfNEbsgX7
EtM7Vl0zAR+wca8CGYgImOO+lfQtEEvCRDcH47XxM8Lu03xcE17lFPNL0Ij5
ZdRpGOZbd6jL7HRB7BbazJihfwv5tHU1MbMazeijBcXVgVcKX+bCgLfG2XGH
IZ8Pmm2fFk/W65J/mEVd8vF0y1jKBKFlSeQX/PZbsHKw/MxuhA+ntiPqys1m
wHeNd4/BmWkZUaw1KGCMP+FOvgfRJe6mYYEjKXGVl4YwYG7aXkS+aYQZvnP9
i2js7iGUE7mkVOmwWP+PhXU4u9i2DhGUlM4KA3Ifh1Szx0hWV77amufAJafO
l3yf/vgjo29EmG26x5V71YW4NdmOG5NoJ+JD25vuPtrKc6NIODrklLnx+vRr
ZDqaefvQL1kSzkpwT0roePqR1FEL5xc9zx2rtmzUFdwMzTzYpihD0GTA0zhu
0E6/YdOqvEs3iFcX0V9GZ8We//3VRli+IcXFUQAjPI5hCipo+HkpJB98yhIR
gbRtL7AudszygMft6w9s7VjvgE7l5D4hL+zPBqUyNpGSkqDwsWZYv8K0YdqS
fq/KlRkYAXLkN+8EDcJTZq18WelRJMToLdDBF9PWEwQ4+/ZYHsrdLBjBySv5
AYIhv4IK7MvxyCjGeGnK8XR1SsEBNWIqjuAhfwBiGiOlwNJFdtRwLMXYDLgy
lPsxVoPxLt5t6QlujhU56x+BtxXDKeTMKQUR9VKgD4/ubACdGDqgjQEWLHKt
XBUgNE10POTAgkufkHL9qLaYVDB1YySSVW1sJB5b+eO+xYHLsVQP5tMch2jd
pMV2WjvGMUo6o5NX24Cr0zOpEHA8JJJURT/CNV7An8MUhxX/w6topfi6z+Mw
3rf2Tw9CBvfr7KQV4GyI4RIfyyWHEVMclEAcmImsw8tqwFx8+QqBnQxSQLv2
YWNb233z6z7p9lQd3nsW6n3K+nua8UR252efE287Qu58OZvbXwu1SLGbxjka
r1MJIWv3ZsB8wY5Tf0WqjSNTc2OZwQmB0IbrQFzdvFjfgVNBu/nlnBTT6EIk
IKETxuVH/KJCoelfY5tMJo5oFv0Knf1LVQ1P9hql9QGIgqzBnlzC4eFgmKMl
fdrxL4E870SjQb1PdpgjVqG8RHmIFUIdrUz7tkrlD6kA54Rm3mKAPBTmMntT
BzUVoazvXtRhX4L0T2/gGUD56Z0l/TFsbQ+4apHPhnaPG70Fku9iP1O89Lo9
YypqOzciEVidMCms8Nbg1uuSnNTroR2hBKZzvcHRFTO6+6gc0pNJ0tDIISCi
dynerTC4cqVW2qMRbG0s46pJW1/VF2bMFaKdtRE8eCd7lGJigt1qPjehhks7
2boUxPUuQdiu3DgbhhOe027sKYHnErIxSBwiKqtdnWHRzprVJsfMDXFgDPCv
G8V7VkdVrmfMgzIkD9wkWkWYkMXwZCw+tJ1WQX7xMAu/CCbOi+Frv/Qov+qe
kZN/zABQmzPYyM9c2hEK7dqe0egEjUNTxqPal4Ic6wZyy2XqFUrwjevwmFFj
B2ZLO2Fh5jJJWs3+tBvHT4bALzCoW8XJRyqxUGkvx609/7AMrws5ezS4vqR+
KxKBIOKb2yHAyrPsAMRyuGPm2E3zhsl57eWSCuBrg1B5qcxopn9uhRzxwqB9
bqUM4b2d2ZxdAWkE1rvxDj8GO5jMG87iaB7DC+65+fAUyj0u3NgiTiHJzN7Y
Wlbgue/rnd9g+qmhm6gN6bjyYIS92wZjF9HvO1oINadSAun9ocORJYHYKzYg
90J6halRXkj/pcnQ8MUCQqWrMq5+FGlSwUlJpMhV9e4RBCNJ6Q2AlhCL9rWZ
XTzvg3TPhvoIgoJu50yu0/3GRuzsPM6GwtzsvHMmu1psLjIic+Ts98+5WDPP
zdb0rKzgXgws1/jOriy+C6Wb3KOuvyyvGJNQxjethKcr6gP4U2O5BUvMXZ4e
t89IC+TKqRrcDb6YojcCVp2N0nt3LB6wewS71kHn8QJcIYb8LEy5VauyebJG
7yE9GCC+uCIVUWx+dIaD6ytZhkV2o/0FTNwBB1cMKhhzPMzB8EPRXdSDB7Xz
MV1UboVPUadJOhJX3qomFd2A2QWVBGv6eGBQ2jYeKHb7kHTdjUFlXwt5G7HO
Ih+uCDQS6Gid626hkH3g8oQwp9r+JTcmt/yRi1yAcstSCJZFaRUXM2g7Y4bY
R4+OEsjSpLW6WRn/gmiC+SBDca688OYWLWVNs8iYiwGWeEgoKQX/RhTLrEqh
v4lgIltAOQj8ca2RiOv9Dii2BkJtHlJPm2EBxUKzcudX7kqnqW04LfwumHHx
tp3lUPmTTmWsEMvU27Ew5QeC1y66TIVusNkpyx+NKHLPKNpFZkUaqDtk//63
39bUlm5PLLda/hOkV4ZTBilKDCJTsIwOiJC4DQhw0pFgCbNaMSkj0ebzpdiK
isB0FCcn/+nBMAQwIZwxArsiZKyEhhn9OG/ob9NsA3LhrgtoEMYsiWj0tj4N
jqy2VIe/BgfvvWEklQOMrLbe8ury1AGadaGZhApbJFAAd1kc6yc7JvpPm5qo
ivLYrv4sztS1o9zt/G/1yH9nYddPEd00/OPJPVM62craF6lWhlrh7DtZj8gI
Ep3/4aMGzzjkt8IwWXhXHXTdAhdSfhEOlyIasvGYNBzBXoc1RAiLSli5AH9F
xWM+5v4uCR36h1g5dZaCc1wjn+zdEYvwiT5ldmEIOLQ8eqWMDlK2Pxf2+mxL
ottyQDV/rpk03jFq40MjM1IRVyK81cyKhCbcOq78P1PbMHWOZbln6rUbhpCl
1T7mY/OZ0SfLale+dUeODToleo1JBmKgQv8Lbhh61mLNt/t2+hlLJqgeVRg3
2UD++eC5AoneIoB5qFPlOPnGRl0PdOzEVqoorXZyVhFRUC8YUWUAYq5guXra
HCvr9wrdA7sMCGNSs2pIw03o3j5NrWG3tKObR4WMHf8nWU9MjMEcdwpkH4XJ
CWWo+KJeZW86xDhA3K2HjqT+qJ4Y/eoojoaICie/ssmsAFww2ZeQTO6dOYd0
kJk27myqfY1bt+tP/AfY0PmyUzOo270U1EJvCJlazQSSOOQ0UgwzhvHlt4HF
F65CHs+qXY4eynStppppDBlKQDzVwekMvX+wDCoGexRDnXHfemzy3n2MlLeG
YXaj91QLRaCGVFn8CV50lPjV3NH+h+W8mjBJAUY3PIGuLzDdz11krqmGe6tC
7DhE9phOpSfU/NZWqeE/5dNDUQNMin/aTVeVOvNFT1iAmJZm+M6F91pi9+oM
hcXJPOxj5ZZQ6XwtGIbKJpffG5wMZe6S4KqiM0UeN/RJVIEybN3T

`pragma protect end_protected
