// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
H3UTB0sNZSu5dCkVrNPRauURorn4pTBhcUWb5pt+WGuFgl6tTyJcQXS9rgoLLxer
ifpicY7wyX83EByhpiZptDzrR9YQgOmFS4GW1ltCQ2BF1S4FcHHFIYPWP3HFzkcN
yqvX5ne+iY8gqlg6Q8vA5hytqaovpiDMw0FdpLTxlZpVbKVQ70nliw==
//pragma protect end_key_block
//pragma protect digest_block
d08oHSHjjjlkKGJXCyYDsiCDHNA=
//pragma protect end_digest_block
//pragma protect data_block
R0u9TUtOKgEshUjZ5SE/2pyHLyHz88PJnh3K6WVGowMJ+CpJJ8Usg9hJIsASfEU8
OQlGGWTodj2Ay2zJ1qUt7S6FknrTkl5lToyhzZ2HHp3Y188Ttr7rifCcL7weoLio
ruUJhw+41y2Nh8JHrVHGv7HmV1ELfEk72I+I3rAmO/mTEODPPToX6plXldQ+iooC
Xk+YmwaUcPN7OP8Z1MtUDVcgrASwBpBmq2nxjhuFKYmEum3VWHMWU8n+pZcymXze
w2n9GutxSFnVDNHpsuSLdkqvKjG638z5xiSDdXhwE/2J8yOLgWZgcH6O8qJ4ep77
F4DRXVnXDa36vEcMydVGpYNuMzvGDYSKK73f2Aa+Ixh1r896U5IZypfxxEhE1pZK
jXMl9adtlF/Lcxjd3OazOf7P5XkhpYxzYJLz5kfD4u3ud6yY8omgIHKO6rEe2RZb
51zrmWC6zrl192W3uwlHwwLYm4GYLGoSUyW6SzonnXcVX9u30PG3b1ZK4R3qd98D
S6DUqnK4FOPeG+vM4OkZk3+byi15Em5jovNEWs9VFp8I7za4rb5I4m9G0s3hxnVN
0LoaNcNj24l9rRpfWWhp60XWXkT6hnSY26m61KarHRMCXwtMuXvRpmUyPCQfd/uX
rgNqGRlKQfclfbu0UEUfHGKGUWYUlmV9me+1wjtIys3XDhUeCNjrYhV0tTmUOzs8
sOP1HEnCX4+CANOKvzf5OSFxfWSvKIdRVodmvyqAnnaY7CnVO0umdnmU0W/1/rOT
sOfMwabjsMasA4EDJCNaSSGlGKGI2wZLxZ9aM57JRpaA2crxxjvQYMZO2McNEFCf
jFrzOeEMgIrMH+XPbEH8CUtX+HDlDpJHZS+aO3KrbmvCftxuKeA3Bl29BPLunHYX
XofNG9b7m7rI0xBLArFLNDGn4Q3jjD3qjKQPhewb9I94IoAsHvkH2lRFqf/QRSd/
arqHTOklR4IHlo8mgXTEv0fgQBo3CokOFLqyhan3gFDCGp1jr03yDJFM6iuTYFjF
mGGouBKF0J12L8v1Fq3PTrifj0EKln9qaWghHABhSYUuslPYKUFsRSx11IHLZJ4Z
Xadjh9VhVn6Z2SQ3PQWsK2WIGKM3DzmEtrzzIVWa8a0LB5nIh79r8aZ8Za5enUOo
7h4bq0cBfr5vrkVqb/0aNUlSEeveSleSeTrxB65taz16z0Nctv+TwEnu1WSrG/Ay
/Jo9F1DUXl8MpVzN10lPty9d+qpDyVxsL80iPSI4R0ONIeT3k+wK0nenU07uSSKj
lmGWcqsWPFDPNjsdY+qNJbPB9l/qek0Esx8FafdhLleEYZAw9KPjQlxIM4ZDDhjZ
SIT6zJg1l3dE8DCnOVkL6RqEpdQHDHA88f2C0CW0rtOR97JtKhKa619DY4S7j5Zk
pamaX+d/0ZM3Hrvl6WQMyXtnhtjeRxYIzoXKZBcyjHKtc3UIC9XDbGzUId+zldvG
7IE2SP7Fut1QBLPHE23DqP6DNUyyfBqMs20uQ6NZqoeYp/LQ+r+aY3dcDRKRA5h8
sE5qSFUVDdoPq5odD3KYX6MZVUrtBsRV2QoMs0znW0aToaUsRX5zsxcY5zw63StL
KtvKZcvIVJECfY+0sX91FOZjz/6RFmH8EbBrmZX/y0uombQR8xPQ7Bzt6qHkRe8w
dkNDBaHUmTohoOOT2sbea1lxygd71Gk6Ttv1y+32CZAAq/KQQOZNthNs8svLUHUu
e85eQW7UJEYRKWO60S9D6HfmFd2AQcpUxktWvL2rmTMsedjl2c8l6Yj2GTUaYRX6
qf9g76IKY55y9PQ40ztBsFvINI3xG7vciG7n1ASZSZEKZU7DSCIyYr7kK/pXZgC1
JUtPYCfpaagufRzC2QPeV61UG7MWSyhQjzhFP81WLhdVQiZxYvkh9qxZrdO7ld1k
5xAFXU7WVQFFIvIeCn7HrKDzejax0biVImEOjoYrP5id31Bv2ew57B0DSZJLbBiF
cWHD+XjXrqEfYJ1MJzAOdLJR3/5NqOy9G3DnmtGMTMGQ62R9EBVWw0CthCg6dn2w
LPf4lRJSTQ/uLTBTINzSdu25TiymRjRjUmtpDLVgHXdP6CAAC5K1U2T/GwW/AY4D
krIABbBfoe+EhCVISHa4JFVvvBMyf3+78qGEEIqV1IUwghLJd/b4Z/d18ltUETHk
G0k1BlmATgbTx5YernbNOnTsW+XUU4rifNPAbeeVM0RkleUPhcJlF4qvvW3CRU9f
USe0Eyl0yeBKMwbKqQqEhySr2wb2hBtpSCwgdRhduVywTCCk2wp74SlFAeLnGd8x
hbIzpqZH+b8IwN2rp8gEHmPj+evGdYeyK1X8m/RYsgBsdoWAolL6JHqUlbtS+esH
/FSFpYnLUNH1HgWxAcvQjNngYqVEaVVc6TN7nCP1e2vqmKIPrcIT5JUopr6FoP1f
wJg2KVpz+f4sB2cCn91AOJeo4i0ZcKRwYyODB0jV21A99WXo17WdyyUrsgS4TjtV
m3FEDnE3mk6yFgv8t8AjN+OORPTknR5mWv5OMgMC7yr2mhO32NOxODZoQEdeC9md
gbyc1avQlu3VfTE1SUF9LYphJX3aEJ4iPNgaPkWAHFigg2jzlWS/K+VoUfW/lv6V
mJ6YfBC5Iu7gqKRdizxffTyjJbWrBq57cmhANyfPioyaDfEbXzCuihzef7U3ogL0
gtv8uBUoO6pJDsTWH/OVn+PDaTWQHse2ykXDKSwwW8B0GayZ9xnT+PswFzK9V6OC
vhRFMn2/Qkg6gMGA+rRBy3tDxenXydjT3mWxgvRxAnoJsOFZt/f2cgeZhqjMkwFl
GSDhHeFiJocHYtLCLMpsjEPhjaorpzZDbrw/njdSOi+8mBCFOqZTcEFGcvt3fZh5
tOe+wb7xwudodLvGZIYQpxwAFJ7+tUCbGuf1Rk5Q7R3vYQn37Ts5Fj3J7TdTzBQf
4P+HmXIYODC1KK+oZrvIXmuqnUnjXHKSaXJmt3iUMxx9Apkid0AOWke7jX2gV46B
JTlSBGvhVFfQdmVbgMhL5mxgFGOPq5u9pzf2Y8YQD0QKTuXRA/JOT5WyoZV+E8aF
76ZXpcHUiss/KFGhfZ5IL6JS7gSWEPuqGm0wpP+iMgezsUSIo3EaWKfT2UmXqpUc
61+yOm/ZUzrkZntsyxsM2pdzu4wx0FzQnYFDY+z9O8Uk05ze0yFYUtw8x7AW92BK
bLM+Zrro/EW9lyOGwYI/cO5rhmEVEMfza1GG6bW1K5ZHGu+rsIqlfjTRd4J7Hxe/
SYRmElXcCEtIzDzcmdZvsLXjypVOtSKRUE+sWMgWfZZTpEZYFWre4OROXYM6Qx/m
w2l9EulG4a3g+IhmJf+DjMOyDgqtGjgO4hTEBZuj09gQ8iU4C8dMjvgAXaNW5KcR
jPvYwvokvox2yhVyKRXRBCmkGGChMHS7YvQxCJtrAEeIZWmGDCSIrzi1Q01xa1AZ
H+aLVUKtEemxMa+957Ju+XINeBvqJe84GmkFnFVArxXmeEslqlYFbDzQHTrOuguq
b+tPtbkm1N7XgiCXhFwksjgDXZCKEUj7ia6tpNHoVVQg6E8lLteMVxzCidll+Ag4
Cuj6PvQNHXlQdDfCWGwSa8ZYTYatJ80JPsc8I2dEt/12JBoI3I1k9bJCPoJQf6SX
pS6zTkndIUfqLH1KCeICo9a1Hbpp1yKNrudWXq8clq93lnznArLMOTIpnVYqxq+S
6fo8beiXeJV473Uj/TxkmJPqxvsdtClBMnWG/2hd1/Kl8mRCmMxVpTGXJCExtnpA
kTtfQh79gItY64kPf1JBAYVMSZP15DCGiAeR56kvb6JvdQHCh+C4XAjrZKsiGZfD
9s/JCjVH9osu7s4Mnej1Q6XNaupDG/Zh5tbRpF+nmpef41z5M3aChPCS1cL3FaBi
/hynbbrdhfHJbrlNgjr2OF16j4zO4Iyna9/LO36eyb3nQuDbkdPqF0jITTXXZVZ3
9We9k+GR9ITGFdCCDLZ89YtHF2maeUU7XEhOhRuudb9zG0+TKzeihS4DfEZh/Yd+
kvD61k20yCS2EcOENOhKJ7gVxm8gD4lfvd/qebdaXrC2DPPMKKpnzxg4V1+wJVmb
35twQgdGsehm0W1ujezxjaDioIJsfVYJmS77H/BXFEdG/7/nuH3UElctM3ZuNOz8
M3zxIJfkfLIuECu2HLRDyA/9v7Kk8cNjmXVVj9GnjMnAoe1Ki/6yZ4taKDnFGf4F
IoczVwrH956pX3hL9WlnDZy+uXTkefN9jigjJ8b6/HkpE6n1tlRD52Lr4EhzMx6P
E3NV5x+29NPifQ732DVy5pUQIEI1uMexN4uQ72u3DQPBrDSCow9D/TrthNilNVqo
4SnqwfXB4fxcQfD8iGBcPHjBrKEoz1vaaXICNc3B0WxFWkVsXmA49n/xNlnQI9mP
i1tvOzDj+uXjYV10H3PfQ24lWbDYYAqg0tZbzKsqODgpTPWGR1YUgYZQ39qEQP6/
29+VGnP4W5DKlBQKsqJoguPOuO8sB6mVCiosUOChssA6VysxS7uIduVi2/sAIIzq
lNYKAV+OP8nTPzUuEei82VGJ9rPX6m2cc2aJJwEMetBIHE7kGT6C1pcKFueYNqSm
aQELF0DdaFb/LEseS4wYg3tT6BVyVySL/nLu/SKzQTyZdhg/KH0e7w6/JrANA8Tn
x1p8Ies/l9E1WsEZf8ENmWs0rNXlkRR7lkRRFHvT8vNOQBeN4gd3amTJrwetxxof
Puiy3hfC+faAVXPSia/QeCt7SqFm2CuT/FrYZDL5Gn0GKNsA3ZlgIAsqtNum/sTW
0WMSyzVr2HhgvVFFo9OA3t5oecgjJqC2diUTQhjjAcs5qC7ivmQhI/bDp/6q2amL
RIfQTfk8WwqAZ68X7Fgt727gTZdJ8J/t4Oev7YnK2FpMxOlUKmAX1XFANauXOqJe
mVsCX1rfEjXAy/tZGsQwwHbe/CWPDeSF83K6PHlV1OZ2D59fihmKsPISLw3T5yjr
RGMDeof5SdHQC06mXTIkEcloxmV4KBUik2pc9IWYCS120mUSui734jxscFAaLbHA
CBHHlkrAPMUPotUosEU6VrqQGz7zkLYFbqJW5Y0+V3ugfOKSsp6C6yXpHd60tRk5
EILgUYVJsW4l4vwqJ9heBeF/Tyq3mnx8mxuNvKgmucemQb9CwrxGFUIhxyOu8qsL
cPmQc0+aIigETDZ4Gg1H8s2ksktiXmOCyVIEn5Ttud2o4YV8OZIkFBtsk1gJkl6e
IM2rE3MxM9MAidOGGPk2O52d2sGJOo63fvnkV15s/vgXCMEoMYeG6Dv9jXhW7oxT
SRZud4reiOpCeCNkibnMi2IqgkK0Cv358GhknhMAjm1Yb96p1qQ9l/xmHYVSMEIX
CNw1hIi1hbhlH1IMB5710KL4hAFAOVHNWP9edGEUJYnvuk+SPY9AZ60b+s3Np5Gz
MY0pER0ApvStHW0sRiMH34AfKvlBVant8lYXfnDjdU7r6rIMWf2hlQWgemo+fLli
VAAH1KjfEGrXiZIBcIY1ZOkvD1bAlXaXwLWYykBO/AkBOFleQCm8+4lixZryNQoO
m+6xTqMpAwW/nrUJ79d34XuHQWBe4qxmyCo3tf6DW8NJxdCv6oWl5d/xhuJa4HMu
xNMWeipXp8nAzkGDPJWjcn/mgdRFsUuOanydbwDWXMnpnd+aO/TMEuEsJ1oXl8ht
aamvyan3SYceypGy4aavNsHAdNbrpo+s5lxdZXZ7uCXeps9OhT6908vuwLZSu3M+
jW3ybcuaZwflPcShb8PxTFJDvFiyLkY5i5/IlJ5uWd5IttIr0IbVM6Hu/jZ1uPPG
NhnSFrN1yPmCdHKuEFzFAWL4ZcnGvlKJsWjOngrBx3iobfHdHJI/SA6Xxcj+7dti
1a1k8ABd4uLNtdf4BE++o3S9/yvAd+i5FIyLnU2p3iikdOj0lxhshHJQ/3z/wd7T
3oxfbbMLbJsUsSIB60v1IrDABSMC75We3JFqlnuCCqg2+FNBcjKqG3QHOEskHtH9
Mf0OkmyqLCKoLyJVZSej5aoLRJOA1UxCl7szXh376Ds6joeyzIB6yKC7+6XhgHdh
0awSnyR0ot8SywzkF344+ep7y2cW39skukJehBOJbCwSTi5fd84/3wNgTFHHpI6O
TqvbssHvqgWKrdPoA4BFThBgFqIrxuqOmPjJKVkM8X/xlOoulH/GYC9WdEj0sQJ0
cvMaLMdmj6E1cS2O/9RnQZNUia5Td1KJUQEEkYKfhnHgJRUaWlHb8spZrEOoPweI
+L/e5iN1d/FEeqxT8r4ysLJ0dWgmZ3/w0txoPPAlwbwZCRHWwVo3PC71dJgvaaep
Koa6fC/lHGTld+9dbGoKI14q4tgDfNSRwtoOVugyWN9Oj519H4+zQq5ihxDE5JQH
bTSqXbLoHyB0JzjX6l7VLumWFJadabe8c6RNAI3aIsObq/O9TYhrqahsALbN9kHT
vQPX1moo4WuO4ss4EUQy7MWwRXrvoid06YrCQ0Ao8y6gWPqEmABe39jUpEZ9A3kk
TjprmqVWMyIEL+m9Aswqxka1zd+BBSR43Xy/ZSWLZ/s9YBZ8q1fM71ygGWHnJ7Rj
tJgJCFGkLgNMfHkKaYoz+m4j8SGYnLxteIzivgeSzBK27bOZDeKFiI/v+UOyZUtx
Ecgs4eaA7VwdGQqVjD9Uzts3jWHmXUEHXk1D9adw2RNDArdR0SjeoSuo9iKvG5JB
NtQBXbhEUq9EXhX5/baBBkfpbMA+fnZYoWw2rsHTyAlab+zycgvst3tDOSCIbdVl
/yh7YvNdoStxbeDZe95gTrDXq1XxF4utxa/bfj1ejb0T0L2Z43zd1p13EdsyIFCY
jJoUfxef3B8aS9EdOJ5lidE+FWjnvREkv4aUOOpixLQC/1aFhlDNhAmZ6GcQDhHR
/sH357G95mTr2S+Plu7Lcu2YGMfmy4Dql1F/Q1nY/B1jJoVrGxPUPwsdZl4gnNgA
i3c1jis9fy1h8PtzgLSW3qeZpHN86xt7Ivwjgq6kTUPo0PcgWTKpZJB+ySxWlY1d
DHDKV9SBoDr6+dKOCkS4ouGvFz8VMkALoVlqrbZlZ9tA/lBxt69jb92CMnTDnEJx
Ql4PBJdDa2u8JenVMsnc91kRr83UImteMwra1BWI51jUPoryPM7uPU+9fquYnujG
lpnQ4iZ+DazSEfvlVtEVOByNgekuKoWm2c9UVio0SgL3g8OVsRdIsrUzjQUzV3cc
2aq+AKaXBFMZvqjg2p0L6hukdbYRU6kW306y1WisFDYYYTHHb3ztwFFH3lxYTVMJ
roa7zbL5qegEueGHnq9Ae6v7Ov3PnyJtyhIWpM3gvEanTgiXH0L2XR1A5Gts2IsO
+uehzUbanBUQaY9c16tvBzW5qCIqi4glmXEnpPPECbJxSfw9aHHpPkn44EnsV3X5
9dhDouRlhTZ6MC8IIJhQCcqNkYat5Yc99Ln/9Unrj7f7t+PixajfHKrqgxLmw9V7
A26N/dudx7BK/h2LhQDQIKSoRL1Plyu+dEYREJWELE+Wi5zTYFSY6+sRsBL+oiik
yzobhqMJaZrTQFKE5TX8nH6A7QW/d3BJbCKvns0H5i4/qfF7d64iZpRpyOjvUMtv
vrfSJt2/XOz539CxKiD8wBKCLoz7oTv30p6HH2iC9uVVaFBwgheRwmLGDNXBkyWT
s5c12TGi11IUqJYMOsWPmvdGdHjDQklsT6vJ8OQo+ZeuG1cOOkPud2X330y++4GX
u5tOcIcyhm47GcIvuFFLicNGTEXPmXePfKGMjSdA1w4h4Z2pQGDx9nTT8B3zp/Cy
u2F5l9bVNLN7122ZDvu9JWZfGsruGwdQ0L4YIQ4x/F0+XrA+FzGSoFRSMoqfe1Ry
KWjfKQBznKk18d+XDOQLWFQ4n7+heiAQyEViFoXsTk8d9rRVpOkM6LNVFRGI1tK4
15EkENWdCUIGWkioRUT4tAWdLAzLWHG6QlFTpKb6OE/bz18ybUXuzM8GEBr5F4+A
0YXl/UZY59ry0pwynBs5GagWIzaW+JaQqp6FqVx6fk3yJO9ipEM4fWneKh+LZaYI
2jjALMQtUBHWlDUTqbNJrNGk4tqvJYhqGscf/ZbKrWXFVStnbReKl3rrQNWKj8/e
4i1dQ2XbTYdHb0LAE7T3u7X2ILRMhPLIHp5tdfEQjFkDa4C5lSWy53rKiZj8XUEP
CkmL7hshIcVAfSnEKZt25CzvOmFPKYCcusMUIm6yg953h+z8PvtgCiCXOqH5p+Pi
NCjHF4XdH5trqTFTyP8BE+C7NSCUOztwIvWB5dvgSnW6PZcLINwvYidiVr8cWh1N
dP/fcFZnTqFQKEMMYfZ7mp9Fgai+X0tmTjhCf0zg98WPEibxmqn9/Em+H4g1ckQT
QYkaoy9MtLoEXJN8KiFiUg/v8a36R7QsKRKmgTuJhUYDlWv/lag374hGe2P1XaIS
OLJDRJz8O6jK0jKoFdtsX0Z0WlAohOF6edm8hS8n7xk=
//pragma protect end_data_block
//pragma protect digest_block
DNOVIoza6tdAcwvTL815FR8IgBc=
//pragma protect end_digest_block
//pragma protect end_protected
