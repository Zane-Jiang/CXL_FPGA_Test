`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
QNWSDJlwwbgW5jnn3YgPVEpfQ3oX5LRYiUbRKab3vmr//qbHH2nsWrAFKmzGGp+f
wASdno4ZBU4d5KUaf+m/5A6xVXDMMRpVFJYDgevXZQ6U+eQrqT/xkGifpRDmh4P8
Y85li9cagyDUgPj1Idh8knFTIMN4TLmZx6xLrpoxDX8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4032), data_block
rzm7lZyMBm1MYatrhSRPQiCbwviaZJyAAGNlXgzC63+UFZKnO21Vka4NeCExxgJf
v1SpV5MRi22QmSVwUc9w4N24hrfFb+0HImgl1PPzOPH8blFLfE0IMSFC7cik/dyE
ZUd61zRP6Ulsx03nOUdzk+oA9t4owOfp8i99Ap0dbyha5PuwM8cuUNX1mZ9uf3Oh
QfvhnppnyvmXA9xMeDK81jFPj54bckspEmqhrbU+osCEAAWivBD2FjqVbKwlmiU9
ixORZ2aRGbh5gHbVcNqkZHrl70vIUA3dktWeKo0l+jKe6Ykx64K3NZaoZ7Zj7Xql
q7oUbr2OazyuDgqm+/nlOHcswG3k+h5H0lpgMJYuOMnydEPuK/UvcFNj53ID5Ke1
0/RZVfaOyn+LhnUI8KFuVvT3JgGgE1sKOZ8YVDBZPHdFjSsEkjBs4ClPiUCj6Ay8
NuYIqcvhJ6+dNp+9btg/qMtd2PusU1J8Nw6keREG5l2hc/WjL5fjAQPz6AfJyLik
PIx+VeFtCpNIQjWYClnbni0ZQiGrRreioLRMhJIx2llRgrl8yMlGg773z9efXVtB
fSmvx77JphM5SBsNgzoU2lIJWsYBjJkHAHzwnNE40cFFpQLSXcUtXWwnCAbcMQY9
bcTwBLOUZb1cURwdyJqqJB8QiC3Q1NMytP4GDx7iQErBrftR+gRuugR8CNjTtyYS
Sg8VpbuaeLuecp4ihPzm8fCveyjCtKyQpc3XKOgppWLt3yKfTelQYrP0vLs0vgVn
CpUuMMkZVvnn3B7AEgigeJ/k9JOuFNITGX+vdRMhiiIBbfyusF31NuceNf7aen5i
npRWh36Bn95sIFs8GExC351TKPsxGMgNChro02llvlejB9makn4xH6DxmrVfTASG
REEWOQG3br7cLTZkfIkHQnsBuGfSIznpyF63QCOnkEggGryThwl0bw5jwUauZ/9f
7YwASwCbatg72ioIZHxLFZg9DLy+Va0CYWzyo9D5q92hYqvP7Y/Z7AZj8SdlM8Rm
OJQ8MWsFbncWNaRSuaqb5z3z7pCp/RhgQlcASKkLzHyDobj3BrB7BZdK7YTIsgAO
khp0U6qR0EFztxzxblbW3v8RBDBU+z26m6lpPLbYZhz/IMyXDOlqSDmrJ+thnctD
1S8bmttHIGhMyoRzpxp8qiyK7xlm+xDV1wEexujNVhnao6nivJIfQa1DWib/6Oju
KT+Z3fkfRNTxLy9ib470bLtnAGEm/J3tGQ0NPMqYwPy4FCMUUbLfnLUn4iTuQHTU
6hpnQoWsEWtu3krzayz5xK7gR3+jpB6uyx7AyvGSApqCSARh9XWtJJFmXnBsVMx7
+gPxAo2OuPUd/DzLmkvptmnc/EMYunogsUia6X6zaeFBSpFYUM2RlOwfR4mL/7lh
puPWAh/uGJUiDC0K/Vu3KpXNtqnOIBuXmHul9nZsqqtab6lZKLog7rs/oZrOC1S2
elzrs8Iq004I8bVVY9yAueSpXQK0MNk40MePDXLZEV06Pgu+JYcMQQRnm7y7Ix1y
1DUk43E/Ebn2f57vE0n/BTtSxbSU7mame9m2kcor8bKUFrUtCT2A9eCIDK4LSJUb
EzJaqor6H3epzWVKEWvRaJ2Bo8jTUWjmc4FTSI99/EP5mQ1C5I+CBUMCaZSsyHno
B6IQ4tz6cK7Ng22ePBFIaQ7T3kqg/6aDt223fR0w3Cm0IP0WHBugT5d0DqT5U5s6
wy50+buFFcE4HV5UyLzpWKLlKsjezcZtqZoR8I54JFetOU2fuO6R/MyFGqbi84aQ
c2Sz1H3XhWap1xujyXCjCPeYVN9MT8VhFyhItvrlQFbeiMvQXsrEbIyF86MvZe9T
GKj/pSPqiKqjO9kc81/JXmoVAluDo9K2vRnQ1fdYtPEWahNtRLXuZhvNNaqyiPFH
Yt3FN+Oyytk4/IA4E9+Tw76pjy3cnN3bp406/AWhOHkqmyqtwXjgldIJ00SgZcs+
+VPPYt7ZUqSeaeBmLoNv0MEdvSRxossM8sAeKm2178xIyey1h0H7rLilwUHpPsrQ
a+c0pn58CHmSLLUK53qSwYh9m1St6bebNi8wMfwNty92zQ34lKGkI+mFzJI4LDhB
B/USAEHQfFZXaXN05uXBmySBmv7XZ4HCABEoU7+N0HT/4uxd5TSF59x57cxT8Ygx
o41IbYlIRHBAVaHkFzLbUXUmM6LmsptsKQcI6WwatYOxESvRfWPbJXnElz6f6wcQ
KJDXNFXvNXoicNVsDo+V/arLKGOZFkY/TQusUpwPzsGMtLv4luNvkS9NbOTH+0i6
l2eFFHRJrK8wSbEOlCLfRyDJB5fsORoO1id0N8ninTW/ZignRAScGSPIOXEEgTnj
VVyneEC/7DKYeF2Wwwst+nOZ519QkOtOc5oMGZldwNWve/W75erTlTrVGYTztfk/
+tIl2LFOqcvYio+IxJ16EXBwbTO845YO0PE++6PUSB/3oind6X1RsZ0IREOzJMrk
qcBLjmd/0Wk4nAu0WvL9RBvh4LiL4DngeERFWjRruDebw2YHXHdoWdWclq7YwHQL
B3ok4aCpzUF74PQ5CvgVv6EMLgA/LMUIdBbD/ldfRKhtnt1fu1cpk9hOel/TCuaa
v7PbN33mdoIMr/AaH9b5WmkPmHSQ2h65jmwbmjcoTANEp6WeeTPhwu+iQYEO/zJq
W3XLMtzb1/JyHvaP9bIBrUrGNwhjjJOiBGTY07slUuOuQfXaBXDC6oFhG5Ilow49
GkXMcyNpGOodVkAk1tKaeV+DF0hNJwEcx+GgBNgQaN1OVlsvL0kfiZfi1UHzIZUO
0QbcElyZ4+HieNO0fjdN34me/lM7RtIgQ/OzRde8xdoSiQviJqHxr3YH/S9PoNJO
SJxbS9H9uDKFEoJzRhPtGEVyyPHkFWdu75VeR0M1xBzf0KALn2pwnwYhjAIS/ToK
PTGMU4Dt6jaZzjG5Z3aDl/LnOTknXsm4PyXefOHsoAlomz5nIrF+nsHU5sIHOiX5
Z+jjtzADo0VmJ2BwF8q224aZe8WjiLxnPxqes+LCtah5buQxtKq5oKTKyT3Dp9Lz
LCjrUwS4qkMXVTxchWucYf0aVfP1XppKERLxCaVhHl8UlHsA4KxOttRMLWnS+Ul7
4vyCfNt5puXzfO/z9L969E6qQt8/ZkUBer60HQAr91qnQzMJIPg9M+2YhjTEF3hd
vCvljofSwIRhK9Lfr/xPAngh2/YkA31oiMqxV1O/l08aij723tFHqx9F3MLa7Clt
yEyDZNfmHa99ysQApK0SZWUwlGMwv1N+vyETIBNJjU18ns0Z10fVgEVyihiC0quR
F5VA5gyNW8/p0G4l8PiNL8WrcP1YIZkiqLfoL5Tf9K1d6fNT9NN+Nq8OWceqoM+6
Y5kWKpwNixj0lWscJZeIV8ifgQnE8me4HxieQe15ctkJtACkXsPLVLsHEAemAdji
D/LU2I0rNG8b1kae2dKiqekHApxsRpti4m9Zdo4O1OnceXPlFlOrzQdpTVEawuPu
6juf5fTttizL711XHXk7pi15YTlrP9RfUeZ/wjE5iSbCu1NaKu4OADI4x3aFnbw1
1CHhMf0CNx56e4iGiEIaUa4x8cXmYyy+u1psVD5SotUjEJiuoUqUn44tAxF0nCMw
Chd/c+C9N/5PAuN+ScKAGiYYMTnenMJgVRimxACDJi4A138C3/17sMJnXckqtIoW
jb5RjwuntWzcJjDGPDPRrTiHVBhHEUKppocGE+j+dhWxw/PpGgHochMIvhnMJqtN
kLRe3URJF1Do8GZjXyaS5wG4lJv8uAszqNpj687MZP6J1XgffjptPkyYUU4vuHW5
vMVQqi5suBYjAFMiRGq0E5c8TU/qDWvKoLmeFXkzTz5N20rGIOIasdsjEB7rceGo
DMMiGIPXETwgbzOqZhg0O4WOO3MbDWKn3MMvKGNgkdpAxqz2rqA/P97EVoM9RZEM
tWeDhfGxFZsr4jTs1hO1isf3z6/6aPHd789FKnqsBS57WoQq+T57p+CGSvkdREYS
xlMQB5OdzJfkTYgnVGiwZgotmhJxP+R2ZOfAPSZQLIp6nINwINBmArBI/UE0DZh8
UC4tsAIxM+u2w2qaOcsiDcDDMYwFuLIaCNe+ViT0cZjcNscbgaXjYFtvISeJ1kVh
byZpPJAiDJwGLeY9KOxT1PahAbnjJqRZcg1+TNIvO48Y7M2tPhBrBQ2S6JAudpN0
3FO1Gi3+rHqjPzS3Pg6zdaUlbO+OT2rYsjxD1h16pwAgSmXmRkPIy40lWsPB32OP
B9EYxHt1GeD0bMQ2zuER+SYDcisZ7j+g80OQUVm958E0bc+9kK6QgkTJ5Q9BMF17
vwAp9yb6GVWa8nQFfoP8kcgf/E/STCS6RCJ1fLlXMFgjjBFFAPYwkh/XuK+Eskhp
0kmpoAl+DjCIk1Xi3qjzslp03fbbP2BgMmq/bCuvEP+OvsDhIyI6LdGoXP18MZjo
7XRZXP1bm9EreuQaNBMWSZUN3c411Uko7VDU+L0AloWpTjQfl5Tr9w3k+JplzCII
VALhDGIoziXSovRnrFyLZsCPMLUWqtlYqRebn6UgR0r1DjnFP0ykqqJJP6mIK0h1
pi4Sz38HBy2KKdESw/a01gRedp7Eg/r8yYZXdw00+kpnr6JyorZA6Iyo0Bbo9tLO
n9ES9UTDLtOX0rgrszkmDndyHRjo7FrISoZt6oq/GXc1HH7hFdk2haaYC5YaUH8i
zkdYVy8ul18CzenweWdwyMU64yk+PzvZPUdG6j+ILg4UQCvuPwqVlSl2USReVPk0
5yHLEUXZw6d+hv++Y0Mfyvwc9cxhzXErx9RPj3m/GGsV+zZyAAJd8RGwpKqAe+wT
6fHwXRImbVdu6xB8h/6qsYbFfc0Yu6ry91TQA5EN2M96bA+XIAeFSYOF+fiFKD9w
/bMPTPJATKDvS4O2fjumCfpslAEy6qW6HknZSoT2/OmHrofqHJu42spKarpHQqtg
3Wbw3SmfdA7sTU7wnNXi9E6J/NK+OIgQTLvh/7yQhdKYZ/TiKGKK1LhuZDnfm8oA
wKFtHw6zoddKp/gbatPt4v+ozjk69EiqwCiWDYf+NaxbpEHs5YPLlTsSdBHJ2wf4
YHoIoKNsC99BzRn2KqeC+5dYPontXQywqr6uL2KxvJcTlQMcPG+Z3ijepYJOPsTi
cvykUfZjoAVJtQpLlcHhysnnJC9k0RMKNCDrRUwDlpDPf/5T5lHi6I42N68TxXxm
1F+vQmNtCglQpk3CA0CunA5mUdiMFjoj2k6y6NxGK9jAKMRAlcgL/imUzVuvK5Cf
nmmoVC0oxj4gPjRQOmA3y4pBc3Rtxs30FlqsBXnvBwZ0YozYCO6yI9d3A/dAGYGE
`pragma protect end_protected
