// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vAq7QV1bc0RxwnERPIddk5leFbfzdSdz4LN/a/hW2YksY+4l215uNcHPFvEk
zkHmvyr2w8X2zmbhTa2blOuxK5feKZ5tM1Pyj65y8xxHXbJFSxWq3leoVl4d
WnAf/DwDbsTXJPPTPW5x58+3R7DKoF14E8Mgn9wnRCb67LoMy5PqK/0FY3zb
mqcImNt+A5iwK09vZjlTC3tN1fZO6BWFiGRE/+76/tglD/wpwfdgcWXIoPUk
rP7WfqeRLZFdjYMEcbn+t2CCPeKtXhg/5nK271oy1B/NJi/qq90WlRWJBWP6
DhLkh43nGHR+HODPAfQo14W58Ewf6/rGzShbA1xvYg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XKNuEEPcNT5V+Xp+B/7IP/Sd1sgUIDOlZSffnD38n0OV5tgSrvYZcuJV3ysS
ajlAnwFB1KiGgU/I77E/lds4i3Yrz+ZseaeTuiA6EKFOphusuR+tQfkNnNPO
vlJMs9WOQlW3VEh56A3EW8nXeN92Mh6w6Rxp1OaxccCmZQQTpQ9aehTNhYmR
HDkGoDsck/paQZszglBnfFxWskYaL6F3R04nQa+UqaygPSUEOBtzyHjUxKDG
6aizzcjbhVeO2SfvDPdOQ4467R3aaPO/M3fNvSI4ZoMEABqEDOY/Rzu/79x4
iVX8b7wGGxvDTycpbwlhyT2RPBG1efVSfN2Zd/N/6Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VO488KPZSXPhRfZIgl/jf1R8y40KSW9nQMPc3Ux1rPO67A2elD0bA+AptiZr
0EhtTdLaP6rGlPdRV9B25Nh6hF1hYz2rNE7HN7CUxU/jiBT7SQBPd3uqCvLU
leohC8t9ygc6uF9wscBR0QNyHxXqt++uYLAxEXTjKTogQFzjqBPyWCtCXE6H
0Cfj4cNfNgy6MBQiqODra+UGTBC6kusJ+A9tG5PpoA4gxLjGhltgaZmEdXiS
qkGs8+ECeN9lGP2X9+U5CTmpj2RG44oDrHwJZsENMJrn4AEePCJDAa/Pr/vr
s2DmOs/DXqGK+IVh+eeRv9jNoUAd9+qgxeGVplQhvA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G9MsbB4lgl3WaOKwvXpE3k9cn8F6om61MvpYxrQOF+ZLomBhAQ7u6ALvZoug
79SPZ2spZ0WfOnS2Ti3mv/wSS+3JhKrYsJPgaQMT0XvRLczzjXQiSSNr1Xmd
oLF7wOLwn8JkxpEO4XdtF8kBFv3CSqh7p2Ve/Wh2iFqgIiMPgnA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
TSWrPC78w/mg6FHJvVNQObfpaOT1yAHl/7o5xXgiWZkQMpKpn5azvl4hSR8l
DKvBZsr6wMlrkO0rYOXQtmcs4KbG8ZudlQUHj454lldVI0p7kfPAc/qWeQPv
m1OFiI4YHmgTJrChurl+E5PiI6UjfnVp3Ky4wbBEL+na2cNqcKI64gitE7vK
N7cy/zFGQbWbparr6TISgj4sH4U00LIFP5A4L+zPg8t6pwWwJ3V19g5Sjukm
Kxw1RwCFGUX6h2PWEwgskYaOdOaBUT1EwXUL2gL+DrKyw82+rCry1d3uXpvd
F8OuuU1zxJUbwb3x8OB5Y9BhtlpPfollXGXLFqGaPviJRzU2ybrjZl2LWPzM
JwrZDC1MeDrW4oWoFUmbmEpxQTalQwV/7wobobPKmJpCx7IDqo492eRMh6YG
7wA8CKHhR/jklr3H7IN/QNSpQfnfYKCrkRVtKFP/eUcSuMIvNXvxJ3rUBI2F
j4aAFyOOa2DVl1+vd5qzuzSyY8xCzg53


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O1L1d/iKJJV+clDQxM54FcrbQxRM3pFfaw5GWtmei/eao8JXhuPfW6Q3TACw
gtDHVF2HecDzSxS8WyXtUu4kDLNDaJm+FyccnIRT2qdVt0Kdbu2MLneIM6CO
mP7ltsTNjtuLKlp+HnnElkvNQVXYkdCg1pt4l5uwQ9lFcQZGn9M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LJI6ZJ/B+ynxYuUW5ZHj0X7f39PqB90o8ur7pEOH5u5nUcUavAyrN1sjMbJJ
LYCObefHepVRMek5QOtc8P/6RLv3F8ge8p1sHXB5XuCd4VtLELse+KJlHiLF
3Gs2wAXUy1vJ2AwAOkvV8UmOnkzDzZu8C2/UOjD1XPEo9S1LWQ4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9280)
`pragma protect data_block
31Rfqs0PzLPEDWnWv46kTB3mwuuphI4t2F/b1r7S2tLaaRw9iDYemVs3vouv
8TT/Zq+hFLltQL/eCaC/2GlxCmnBTDFYsABbRbbqLc9LHlZX8uHs0KPffUVv
u5ZsGHOBZoE99XVzEIm2B7Y9coPpz3eMjd0B0Wa+eJ+tnzBjklwhDuJIgeUx
jMPGyKM7vM5kRfcuPWDvcCav6LZIRTWTAiL87RX9SkXC+a8q7pkikZAf5/dV
rsrhqozmbl7wdJED1+Riio4gOgsaXd3eXpqQUMLkEr9wjb6ecV8S/5UjxKfP
EoybQ0ZHP264Uq+YOXUSQlxO32fhhsDxZrDJzXNfoAW2M7W6jBsGI2FhpqMO
d66qHP8Z2jf7duzDme7JmvkaQcNKN2eMlAGcgs+YQ9wZBqfDsaJV8DOcaon0
AgCUDCK/ALHaUDw9niXIOWys9QDd+ng2ZQAeJ48h0+Dvl1vv4dhjUpYsQrIa
fCnpdc7xNOfuXMpBarMbqsAFComPk3NvPS6zd6E/0dQsJJPCjwTgNYVtlP6J
Z6iUQfxAsiZlWZTU9J12d//QEPAQZ6jUgoECn6YJX2GnjNpJx5QfnY9gDfHN
cZGHglPhFNZRE7WmzSumFeUI9QlSE5VxZFEpYbGVBop1EWNjbsMX4vbuoRNE
jk6+g8zAuRRwmxW/M4pd3OHvHDox9bZVYGq4FO4kWiHrR07CGXa30Tnkw9fU
ecYlP1QGDvZZIghy0hHSDOe/DB0NZ+idTlgKJcMOVEf4DRGtO/hOJopG7Z8g
+cscvDOHdGZthZ9OLbQfXLaBncT97qulfzljhtyOCoCvLJqb+t2k2nc0EiMg
5aWu2L9I5jLMWPDWBcRkYLSmx48L9MAEtGHdqfyc1tj0oaja0dBFn9nk1xdd
OKABMvl5aLtZJ6FzyBiXO7TY0pYRxQOyZyVEZ5kw9eSAhbp3zMTWt8X+UpkV
6B7goA01MdVGXCl1EO9Yfa0qKvCBu6EwNSz1JePc34zai+ShsSMg7ZvqMIQF
baZo/C22HpjgxCQ7JPdjJzyHAycJ8SJTUY+02YaqbLjArHfzX+xUe4lyKSqM
rclcXqehdTQPpiJnqDMpOag9muPpL7Dyt5LYCvLrYTob0RPR3b3jugKHALrz
zvOjYRpWSaV5SGyM3TsL3MjiTNwgVct5XHCgJ5NAPmhNW1A2pGGAGQqbBoZ9
Sn1R/HuJtfrsj6RxGnpVB0EN56xGCKmMWx5rpJwotz1EE8uNlDfjfuytH47A
KzSCCQNLy0cSu9XAynKqULWPpOVAt89wfm7E9NR/Tdqdwo2X3niPxLmmaS+S
H7LZ4euuX+S7IScxL5tKDwwD9U6lwiJG7mXhzV8U1S0xD9gTIwLKc8AiDAcu
VMz5ZjFKywT+N9xzEsmcaPMGLGDyCINuV+AZRXz5zBCG/7zWxrkZsTxrv3vt
aLBbwgzGlOgsoW8kKPeotIr8GwtC+wR+PpIFquDAunRaGA4Syj4KDkw7dL+6
EUZ2ujFx6ZfH4acRclCAU+QOg/vjtb/c7JdvO2A2oUY1znjkDUFtTDccGTh5
e6T/fPlOwsxgCSA9Ys9Y1B1lpC5UcBiZQWC68VU47zWxX5TJ5CpJCwVKwTiB
oCuB3y1xztjUDiYXcIREmRfpGLU/yokG3w7h6CH/CApMEabMf8UluzQ2caCX
2KY9fvoPNA8IktYzZNe8qvG11A8AaYVnqmHTEv5hMB9KGcR9Ky89JEQb4zXK
TbH6FDEz+A1i1Ti+57DSKfh2oQPWbt4R0I+mWWEia6mQ212tS3Uff0bHwHTQ
EI1TkcAf1NJfnqJCqCjX7I8v0Hhd+9Rfmn/tWlO2t/6vEzt1VnZpB8G/VAFP
RB1RezNL8W+Cb7GjtawAhA1F52zkSsO7ukXnwCMKs6fquvHEdFcszdIs7kT4
LTbJp7R/TO3/3ZDOh4yJxszEWM22dR9G8dM+rffzoOduCAEYlTxHec4u0RwV
e4C5vZKFbk11CXJB6NsXfrxENIZqFJKujJJAWdWpg8KZUB6smyjWzdlkNMNx
LcDdtjwTiMDdS6/O4POOLPee0zFoL259AnutM5OHt/IcdMFQdz7vwP8EuWpq
jUjT5E4G6dfg+hT1em294yX3R7nTUetwuScRdiGhSFaWtlKBCt7fIiocvUkj
Qr4bvBEW4RAYm0GItzs863PCfB4VqM9+5a9Ua+k8hfkFpoWpfMame9EWVOFJ
JXyJ97WNP9B/6Gwsksvd/RBgeb1wnrt2/qSAD4lU810/fSxdW1egooP45sCm
/Tn9TVB8qJdlswlJPlZ6Dd9ITNy/ASAmvhD0e+pJ+QFPkEdLcXxmaXI5AdLd
aF3mADTLamZUQu9guibRgFg+nKaLTkgDsLBn3mX6oKC3IHYDXnHX3aiXDqpo
IgRzhMzqV6ULcf8mUvJRgWgXhNYUmf/wltex4ds+Hb8VJcTSg2Q+I4A2UDDp
sYTgOxjHF7oYkYxuZ3wYDGIbqpbMfQVd7g4V2TYQBmelFLEbARv82mpS5ALp
Bj32GRG+SFeAZi8Ta2v/JUQmz10LPBJLC+hHgvhcL+4s8/hdhkNfwTtbbD4V
AxbvJ84v2z+H4tzaIwOAkXMe9SJnBjjpwGpIfYkvFtEZOOTyG5qfv+caLQBE
GE6mGd+AgsFVjtf+kX29PLIpXxlyz7/poudAGwY5GjBBpZnjPchJ7yb8+S0z
kBP6aNV8foMl1CmcqrcsVSSoVZJ1aCXya85K08V2LuFte9gOHi5fjZmd1qJJ
rY+lUqK95+S4SiIZDW+igId4T6LBagYG1ncs9NYTj44wVKjMW9TvKhlmlIn8
ICjcem7CjWbwkMdaxPkUvuEtZcJwjDCCBtdC0VZ4/nlYOJWulpFZYR4Le+D5
BeCZpgVqlFFCZYmy5TeeISn/7jfDnqxWJyeEwFLRIfmhAec2Z4qpiwMX9pVa
0QcKhZTGIXWPmJ2WztEKzbAxuJs2+7omraEI9o3sQJEvfI9dNsczqXZQXckh
xVpeqwGxy3KaD7KH6nVYkLsAPDHJ5sr6ue7alWHK/H2QuO3TRUW69wgeDoXT
WoQNqFU/GCwfIAcXMqYYr5rJXCwlrPUEJN92qbcLPXg+enqRDGO/AmqgAKLP
CHkHKQ6D06LrNEsNQ7hgj4aX0ebwIO6DXzs8o+TVfhrBgA6+ggUtSfdTkQXg
jj1//eiAQ+wDfSGb00EZZs+FiU2WtxhDWBTXImxy3fkdhzxSnl/YlpmL0VGg
CNKeSwyyCVnD4OKGCoNsaBSyt10cdt0xorYaCXZA7Y32n23OHvtVqscTAa9t
bDZ5kbCyY6CgcoelwNShQ0KDSIkKz+WlyLOE13uJsUbS9lmyvlKVbKLHpfsT
swSUAAF7omQMfkxtME7gG3MUe83cTYirEV+L8/u1X9TT0sdKb4N0j0vh76Cm
lGLCH96WANaKz1kpEjbAxRPrJbMPHMZYEVosCOuEZCbzbkIXX3XZWwVU1Vns
DYA0Gs4JsQVIRa514wOWWz+R8ZWTLFoQ29sCMxF6g93aLBilBbGSCafd2ORy
2q3L96oGTGb1qfFW3SaAbZaLThy6O8ScdQh8P6LZmxgQ/54NyUxpT28HNThA
rpu+QGeVLxkFiOs77rEjAXy+wq3p8sbECqkxk4hLOYGxEwqd84Havs3uh/In
B/GRgpPW1h+9ln4y4cCcbvoMu8ayTye8bu+BWAGCu31POC1TJTcCC9EK/DNv
1gY1j1kChNltHh7yyJtOp1SQgDBIV4mAxL7J1Mfvww0TnY/hjwbyWaG9pef+
t21bIectBB89Nz7Nlr0cfNBPNJVgjhtcShZDeMqad4SDm68ZnwB7ZkPYKQTx
LsyUwFT3+1GlvYYfzSpvfQx/GohUOvXwnhBckcEVL3CM2TjRN+15SEk/w2Qm
QxDibdsGVw03BWer6+1dKDKsTeGgvbuN87/PHpv63B5H9XUW17vpF6Q4UFq7
MABcNqMxAT6lexHAVZ8Uxj11NLegs7tFOCUzHui7q4TUvg1FLWUHylrnfu0Z
pY5PHve3Ye5+f3bBKf0uxJbS5U348LrPjxRaNWW44lSFdmIK9ZIh1qVke+4Y
JdAs4w3x0OsJjk05al7LGnkbKdJdn0JGEJJ0atdXwssDaBZsvwMjwVDtx0wS
MT5PFbiqNmqnLw5eNpAqSLgGpttl74m8k4NS2ixQOfUtgaPtZNarCMMdySV0
lqTuS3sKEvj1eJdxbUNvpCEkSOgx2ZM1IK9WLo9u9n95v5rwCVGrmAU/sP1G
rYXL5HcV92QkZtBWEai+bqP+sGau+XhjMeXLlIhq2GUHH4zwjUebUIDzSXBR
c9YEvyyoW/gPrEmhxBzwm/OCQZVSz2MhPMVAzsUVqsN3Eq62wXSFLIOzmBSY
vSS7R0fKdxtyQUq9Z7XMiHMa03Y2l2i4t7YNIfrH9J6wMVkVpIYiz0vcC/UR
c+RxVzKJfhNFLKrdZ7Bk1Ewqn+lakxYJiXh/vRYItzFfxT5T8Mycq775TbWy
xUu//nI3ao/RLJZCtax670Sj5sEoxNc4FgDCmg4HE9cnxCX9Ex8luT7XOVM2
sKOY6KNr1titdaHztW4qhSPbtpXyyduJYRbOAwlG7IRX05kvm4/wphtWO2/F
qgjdiTPSZyMIpA1k6lIucnyKlPukfhufW+8QOEkgqCjLgcbyRCGDy4P6l+Lx
oScQV7UtblEcZRI31Cqr8AMgWL+JAykKSh+4rCHEo1HjgE1Uk8TWNcFBjAyU
F6fnR3yJ05Fo7I8kzC2t4osNE6oAuG4VPhx+9n8n8VKF85Z1uT2TDNp/YfN3
X8lxqU4IM2J3Bi8YQSI2k9EhL7h7djSYznbj+8xN63bYThSA6SxPYoSZbtT9
CVaTTuBmjlXSBfa3uIoSqguupq5HxZRY2UzvDTtODP/U2nOwE4oYzd4L5R1/
mAefuASd6yD56MUvisdMjDiXqOtan4yCE4l7w3htcmvxCnFmw8tSwNTjb58I
lA6JMBGKmfe4cR8k0Hb1BQRa6SU9K5PwMkt+6OX47XdLdbch2ahHyuF+GsCH
jCCkSYq1EYCxISrK8fp+OwvoRRa4ikADHrFyGIG7u9X6EiipgBdXLgwb07LT
/dPot2+KEmTP74PRBOjva+472a+o+fdaS+6Sj//+dqokUMCD6t24n0GyqbGU
2oJzX+r5FSznIh037C67JTaCQyohu5IG0lxIvKCYxC2vUUXDROZ3o5P3ICAz
mmH5Mp48zS/I6XVn+svZTIwfpbS5InXdTMbLPggLaMSUS7+f2ulURpi7D2Zt
awuf4Pe0iDlU/dDZKZqirvrc+iWfBry1w3P0qeJluXySXMdvJl4Wi/C2M8GK
pXrUpluHEQTDOk/lzSR1jKXmquKh/JMBFIHjr2olgalD1M2HEZOWvsMPAH6/
vJMR4I38Bzrp+LalU7ByUZTsGZ9TLPcLLviyywQaSJLcpvnED36nSC8tsW12
MPZaYnTlEgGFOMxh+krtEaWURt4r2w4++GwWR/1kXUziOveej8DMglZs9C6o
kJHuNHbDWoOwOLJr6qKM8Qa7ZhkxQaUa07tuDODiTOLFVxphNJlrSgDuf5cm
43r49P75YRF7VYh1JUwLYNfn7QnOBU/FIWFHc609oSpOgJa5/1C5YHCMg2cM
4vP8vx0s0jdaIjDzYIknm5EaCDasFIuvq1J7ykjIrRkArN/UqAUYKNqBvucT
apx+H1Q56pZoWAmFPSYwL1OatDaNj7Eiqx+pDL+P54D1Gow1J9CyGDkmTRTd
vsWkEk7BzOqrsgingldTCyAlcrSmnu7BijF4jSi4OFHofAjeMBDiVaEq018a
GYr1PKzLgHYah1ovHNia8pxcAg7xBcoB16QTMxi6y02cEFed4HvmNeG6qtXl
IzN/4gIER21zNZFzjkA81BIfEaF0ae2oCmG4NF2iiuzgGc7aNXeC6TrbX2/q
++52XUee/Hyq/s+P6rFqRJYmWebAojIHE3kLnRlBJHoy1jzsop2mZPgIlpMZ
9xVE7odqtw/PRZERU/ocMQfgjIiv+sXi82sJ/hqJ6+AvRklZJvAQJr/wsz1+
oyVCMjT9rXBAlywS66A+Sa5sbKv7pCXllW3nC0BlXq3/+uwEW25AujfNfjv5
bHc9Qkf4kwxzjpS8kRfWlvVpre+OK0YuludZliFYwSvyk7alm9tWly7IGCJx
gzH8MuwQ3CEY4aNo5JB07NEXe8wmeHPcCsYxULQdB8jjyoou69IXIGiyK+8j
QUeZaxSEweDBuuRbOVmeGTzLvfjZnOg5LtUDgyX5wsCW04TjPiLM/TNi6gmW
q2S+9h2GabkoYFsF1/4w3MBtpc9pwPEu+bX9qpYHyy0zZs+ig213V7rQrTLO
smZYgDy+zlQFYB3TxHEA/jgamyiCQsvUCbvwhAJlEQPeIPD6Zd28bHfaNiEH
sw8/duVjr4yiAzdwRgBlF8LRjiodW+3VMqq83nKbCFJHuXjqhSJoYdmZwufG
ZP2HoD3lCrYrumFmJ7qRnlEVsySjRj3bHynOcgbSAO4WUf+ssJY0UXaF8KGt
u3Hw5wt+TmIRYlrxVyOodb8xlZrL4xx161Z9E8N7ABRYGgDEYW+/YCNGoKlR
ig4eR+aC9l1mOZ+AMog1r6HQgmjbsiFhZeBGIJ8YCdnpeV6ElW2JZDnK7vTb
j7773rc81NwND9ahuBuyt8ZOVR/VgIrU93I4ohVK47aLv7nLSQTW014OxTgE
3w51ryGdrMp5AYJwWwbTo+ICiF3JGKR4YxcROCcUcw+m9R6k4WHdoJHJ90Tm
dVph+wOoivGDP1MzTcmTDgRkUSNRLHYuA40iDvVBRpMWfl8pFfSQOlUKjS/d
+0+5bdAzbB5B3+H4NgawwTcWD5FPcDQpi8THDtjkJaWQQwUceLu7adzdVZvQ
8HyAhQFXmSp1Fyy1b92cqGl8vaud/v6TMRX1+pt3EyGA5d92vcAN2nt3Vx1S
WVnJmup7DQDUyarCfKnp6as5g/l5bn6h+4GxgIC7AnNMTPp10IlHYkUrfsFB
dP65hdWTD94h+3sXnZPH0TAmePNjkmJaeLISuJ9ER6UfXmYPmwkLk0Q9S4Nb
OeKrNrwd4eCBeqDYBNEy9hWXHp8pTrR2Yt5qFLJMWud17VB3OdCnQ09hpd9s
jJq6ZY5oE63g+WQkZNT3CKPn0vdSNapmaMfFg/0OqOg+uRoYkVxFfU2V5KH5
+9bHhnPlZqLWCApKmzqdQ+UueB52QAik0FUiLgo4i+gaX7beHdoueCs/vt3S
HHoHSYrE5MZ30o6zgR255ucWCKKoeyu32Snn6aY3gjIZqtZ48n32VELIOGPU
jN6kToC4mBiA09D87QjpIK4O7myO3uxQRnXvo71nPXAk88GICPzOw0hYP36S
2QjxF3iVoGD1w9Gu6EsMG5uVcJd/QOV5L73I8LOk5H2sZ8cXX9xRnDzJ01wy
QY8jynkFrSwf+TmhuCi1N0HYLhV4E/7xlHSlqp3D0rlKcljyyKdfWIwH4XV5
uQ9FakxKADZAba4n0m3cWRFZr+UNUaz2DspDtMDhaZ7+y6aVT+JjvwxGJPVD
9LjrMTTBWO51Y8Z/kcAzDIxBXtaE3iAh9ZZKxsI1DYLB/4AmBfgWFw59fgm7
m4wJYspjllgJCJVgFBx2UWkJdVwibnuPLYEK0atjNq+5YGxC1PcjuFV9kEbK
ILdHDhcm1++Tbb14kOUAAmyXsxd9qIA1EvuV8XhhvHBuJRxY4+3iQkQdabe3
1EO9l6SDq3K49I9jzH/e0KsrAKzS1nDF/ng4tYsVcuoYotxEKmrfuXlUBvIG
5l2qIVOUB57CxT79WY2p9oevHjcb7SH9oaejAukAQqwEP2AypApTJZx3ckeS
BE2cAag664GqzJdC5aM6fGqc/gGZcCM51rt0AsWIphwzudpZKvyrGtAF0UtE
PhZCXXHgvnltMdcdhtNW2KtpHDmEnegM6lmQs76bLmcgWJaBYuhlmiZIvlFl
NFm5L3qJxjuwVzvQKCTa25YV5N7C+d2waLj9xD3WXJurihaddVucm0DT5m64
3qk3r6lnuQj3n/ql8DJd+O/qZgIGop0mlY2DZJnCJsEsXawqSj4QO9hUQGzA
vM+cSFbmO0QuxpRCDQT1WRRvk4xti6CsFAtobpjPEfi/Vgybgi/2VQ6GZdp4
NbvrBqUnf5lt4LLXfYUvI4Ema9Y2+dXm5AnPzCE7MQYVYokQ2jD7uk6/jkEC
+bMSSPzEir3AASs9owb6E+ttZKV+7C6+CkXoapdCMRJVshRftmxoEE46WBYc
9RUWk6e3az3JwB0+S/Ga8h1uhQDKKd0m4vuqiCG0vaPFjVcbgsGEELmt1c92
BhBuPmgG55zVJfwFIlDBrrZKK8CPckVvY1q3YwN0PeQpbqMU5TQXdYphvkz4
GsP7MqkMfplZo2jp/84uhelq3bEeyOQXD6QZUf2zcUW6zWoVGLTFGzOwV51p
GUjfjl5+2hyaFepvfY9i3pDSftTgPhYVEfXJ2kuvq15bOGzb0JaRG8WTvzMi
UI9XbRN5Ofx4gmJpV0wyups7v9eSsMcQSIvGcNV22KwTUgP+ObKGVhvC5+BR
iT29SWsl+pmwK3tvYCkLTtDBJYef1Dy01WWQcclZuA9CRVgpz8yghjSJ9fBF
iq8u7EmKjDk+1wfi+OoXY1g37NxJR10I2XmWc2RcD3Uk+XGax2oZ14xk543z
r0LxMVhR3fK+qhqxELMDPV6TJJglwL1Dyx6O6+YHqt9r3gWlilJVXDzmLDyV
8SnUD+UG5wUqkmzagIqx3hFsMOfPnhN1u0fHL7LZZOBESO9DHojxNARUR4uU
49eAV4OkGqADAcEoe9DTL6Xljk5DrkMxfqEixDp/w9Nk4HvqBL+b036QUogD
B2mlrUVuMiZZH9Jb5uJ+8VcAvCvQdow7x+jiXjOdrFeEvs0CRuh3xwiFYiKc
pdESQPA7OJgJQIb7bpF1oRNziW4ghIZKkFOY0w0103dclqe05C+4wJHjuFvM
bAh9efwg0xzhMrZDvMRoXSWw6uMjEMnLpHCryFBold+YNNevAqEzXiMbALws
IC6GluC0LvSyWtHbm7UmJP2GIy5HoWgwygdJ0GjLBAhE+AAHtHrVoHZMDfAo
L8CRc2g84+5NhU2EaEbRX732enud8j9Injy/nYNYnisUIHhfBjmcJM3e3fSM
yw0KmFXRY/8kqbAPed4TIdsImMiUy+MnHlxm8G8KRVeJmSQ+QB3wnGB/BMGr
tk5hmYTL4c9TV/Q4IAModH7ObvU62LVJ0mDZIB9sorAkLhXacyXJjrmsKmRC
yDWzGmDSfQ0uQODsAKLgCQJgnaABxCSo/f3RrpVJnhavv0NyaqZOMof4d9Kh
sQ01eHO/yuVC/dm4qrlbZiRvNWz/ZMl+2QwD36zY22C0RlV8/+sDqRklZYJZ
NZpDBArPd//o8Ngs2dUt7YrcNPGSBlDzFs/46ksiYSk5QVaw3VvtSFnKuFI5
7nIoV37Gqi68hZKxQM1WzxP+wa/+wg+i3yZKHbQgssyxoImm4bsW1WSwLhr5
CKvCpPtj5Sp+uE2KVrGjn1qiPBFYQMJNSyCO49/V8vyAOqTKO/fucdyenozb
A5gyNAr/s9i/d3huBsPa7ZVbOF8zjCllY/xfYwm4vC/6QtUhAiImP7Ah1fjf
qTvEM88Pp/OYfFuUdwU5XMLS+hHy8LCV0doJpDZ+2raO4qQRabMiL+QGsQyh
86QyWjBEEs8vfQrc/VrUrPamwlUFzXyRCx60Qt0DUjeSVkhXeWdntjDhEJ96
cttXJu033aQy78tokraE8PNYIgAhwQooHyc8EVL1UcPcGyAjqQ86tyq4KT3f
ITzEcModZPh4ANWlZ5TznKbO04BDoiLhu1S9qyI0NbQvk+rZ7n5UgkH05b//
UEU85kv0JR3JAPPcJOrnq9sdxEReOEeX8MOzsIKCy8Bulx4uLbU4XRbA24RB
ayy/OXvqPsGNYGrknjYCVTwjJwgaKwSLbDv80c5P1c2aOEEMS1pFfERWeVLR
UnX45VoCSRcrB21WaIMIX5f2pJCfhYUH7cuQhZ8D0yb4UZvLcHlDGBjt8848
ouCipK9AFqEOp5dpgtcWoSJZDAPPNN3Oyk4se8Vg2Lhalr7Iw7ajUVmD6BZq
fskDFtMQHyKOoxNlwyyp2aXosGWgKjuV8NpDa5G1mXqcu1pFq0PM3fuqjdck
WXboFKZYgNo/Hm2JeoAs7zQgxC6BCngevSuuF0fAL2o/goAz1QlUNvh9tC0E
fssWpRMJSqoAo9EqhnpSlg+iKS9BRSYUUcpF80xIhec6ZxDll9Q2xFVcBvet
eOJaXXiPUa7KD1yDiRQQNUAq8cTUBynp33wD/mL6b1vLrAVATauFi6JxE3Lk
nhQrSiolBC+FSKqw8xbahwLJnMzpZ1qvNdHaZuopT+OBWNw6mpKH5HmbVIgw
mRcxkrdtGXgkGmKmH4ne3IP5NLwfRSWLI4/C84DeEpq29znhaqJH7ySLtizm
aIMeu8P0ECrbD3q6oTHBlgKtLPm5XEHkuYP/wfyNt2iN0K72H4w97+Q65gDQ
IS/qnPeIu0BaCdCfHvc/DtrTn9gsuM+hbvWBgLKRMC1GBrMHZQIMddnDNNgT
jIOJbl7lLXZPnR6mZLkCZwua/oMZ9F3SZ/OCOyO8B5FS//+cOL7Ue1o1wyBs
AnqJr6Aud3JfBA6R+GCE6BJ3it1OUc6jjJYtxhL3UX3WbgoUupJdVfVEl0Px
7ilb/xyQFumWiBzDnWrVj4DAowszvdeHSu8MLk6ZsLjrStSNbf/8LLeodISn
yWxipYFKegZngaMXLKYSDzucQm9VtIi+9EJyvrT5dQhByA85nyx1enYOXsAM
OaF44nM1sNd6Js2waBnCgSVqJsIEjMQcB9Rctl/kmWXA3hIve31O9iYnK2O4
Sd6aFLKuZNAadNZumoLH7mlbdh4d18W4oHoV4ZR0KC57YN3khw6k00/5Q049
bl9oJ7xLuO1iKJayymcTGa6YfpaAUWt1tWwSgrYRyop9dgwgNG2q14c6YN9c
OMc2BMJ3b4mLrXJiVYGonDQA2Bj4+t3/VwiWVxDUTTdLXT2sd0s10oO2yWoJ
nTeXt+UfvMSzQ8TaY4tugJHN+Xt5u4K0X7hZxM+ZmaOLlZTCzsm0f3+QY3kP
0DbwyENRdgIwL52vnBbdChAyraNUe7C6btLFpEwNaLCcQ6VroiofsKsRWGK8
VG7BuNH+r6MHH7T3bKut0CnKfhgeWbbLHjEWRIMdyFJgvExwR7vBoFkGxvjn
vW8z9O7p1Y/OK+wo6axZHJZBnMTOMYUNAexQSPipsqfSem/xdb6DH3nTERUm
gK7SNvqZ4Zu2bJOmyBelhd+7QhvD1hfXzCeYaXIOIQ6tQUpor/DAHRVCRM+U
OXS68HGL+BQoLJCqQyhKo3qOtfhbXLmSLL3assLNUj/cYmHqmzwZw0HvrSa3
mv5UyzkTSXmJtA2pFO3sLjHewo11ZbppRS9pL/yzS2M1xvHnoGNflceyYZr2
29UgPBBL90B9Aj9edagVbnegykVXc5V/BgHdDGq7RmGJM3Qp1I2HVTiA2QOR
gQ/bho/xIveTlwGKizwOWd1p/YfJuNpIUpfuXMBwmHmbrksG8qAc+xvj+p84
kZhmd6JhwE3kApWlhHLchWaynpVaYFhrR67cTesnGh98XhBJgtkZekPy5Xhp
l23ZcxjUSwvadm6l+GF5aaOmBHdxFrutV5scqjaW5W5Rl+a1QcGqsCr9565O
mTOzz4o1AoYmgg2gaSm6XDbyc6j3qYPZYdQEH9xi5pLy0uzXRHaeaJb5+HSt
3wsyzchP9/eDarqQqL5njL9Mk3tiyeR/Z7KCJBXXxzMrhGWKFQ7Pe2DqRAod
cmD4QGgKsGc9bPtfokEcHXQWRMC2ym7mt7RKd/pQApxcyNzLqXfhPcsWJ0T+
XkgX734aLJ74j+gKgqkcn2RHz2s0i4KWA2cHbJG5clOY7Vy7iALW3I6saX6K
vuZfF9DG0WCdC/Cm/HLEDsADRg8MSmrgUMSrvQlNKPE/QiurCnpajnsSjatE
EQNVfYaRxfEmWBaVq1DD/DuHeN8uuqV6cMf2XwpmmQUuyDNXn7vXZwrSwPbf
0OEp3SMsHCfT8xoGDT3vLLw+jDTk0F0f1w8V+NodFq2phTBBBhb8Ad4po1Tk
49TX5eKmOR5jzUlPEIf/CvtwW96lQYtWAEpPQNso2C0+lycRmsLSmU78Hz0E
WXJMvn03K9sIgPULstenwb49l/0Nmv8ZGTTLasKRdVnDtr2ulvZ5uDVEUtI4
v2XduAm++1yTLvFZmMJDWagvP6dyCkd+3SxKmIfO0tHjQRvlO51ltSGT09YL
ajPS2PRlCvNFVw==

`pragma protect end_protected
