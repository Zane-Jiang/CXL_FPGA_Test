// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Whs7tcKQTmfTeds1hlq7CX71Iud2HzcZEiraBdibO7I+QK0bv7h/TLp55Kc+c4FP
XWfyJIlR9Ztli5f+K8TsJKsLfXbnWUtvlU7h0KXX3i/ItPG/AZCYXSDHzMhcb+Rh
UbHxqgltaVLxzJ3bxnVtFxdjOVJQ41gjgVjEhho3VcXHCCkGOb30iw==
//pragma protect end_key_block
//pragma protect digest_block
x0FR8Ni5mXQZOcc53phE9KfQAVI=
//pragma protect end_digest_block
//pragma protect data_block
EtHs6EsHpVYkBC1qd23457cXRoASChLmnx8q5etGjqgownRJN6myfnwJ5HXWbjW1
LDSjIBWNmzyk3D03/O028cCz7JYMLOCy2ylA568BsoskzDcc1FIZpT4g2b8PSVre
WveJFFQyWnAtbdUXC2ZbjPv914TUymHh41sSMi6gPh7PmvpcErJhuKDybwGBB0zR
MxUn9O5PzB96ysqqnW9gk0tCebuo1QTK2c/i5hAJdrAuYUdJms8J30hT3C2UaM0e
xUHm7httP63/WbmPaY6sEkxguFCxQi/a3npm0Bed39Q4BOzgj+Ekp2uHlbBcyI5y
WDEHwo3dFpQU/EXTJPmYyWB1adOVWj+BDo1cABA5g8KVQXZwdcz18jmjkZkumGHi
ydFA828+Lpk4024mMu3WPTkjtQHiFmkjwF+yRqikx66x21bUTTJPT5qWu2h3dyJ/
QegbaJArKjK+O5c1jL6Jo+Jpn1HgrnhjcR0bjfwjfq67S7Q/5a2ZhzAv5HyUG384
KZ446eK4KpN2N1Fxav7C+YMK3xWj34pNSh8la+uKqZaeW7J35agXtfkVg6ro6PeQ
MlulCGHgwdrPzwvrP31e4KxNCx2LgXThiTqpnbSASQJR95LeGx7TaeWy8x8VQ9k/
HUR+xV7iRBn4m78h8olq2roJYLZXQnDoCX/5WQgVlZiWQ0/DMMDxa/+ukdn5e1Ak
xmfPdo61MINFktbUl5wNrqhNcy878WxUb5gxrb/iap9Fj4c5k+TNdLQnT6Xe3OpE
/u6NKOK+eXoYCglK6+3dfompfyUo8KxAT8ITM3MSxVhnvUYrTndvQa51W7G93x1Z
A9UoEaoIm1ViHEFe3styYBzT5M9CveEQB0R3fzHuKofnlibw8Gym7Whl2D/SPxLD
JNMWKp+eDznAFCnpAT7ZBFGilL6lQrlSQlw84/CLY36A096ufHswWMT5P7W14QkK
RwLRkXDQHxXYojOMW/w77Ldb756eGggw2chKArPpwlic0N9YDTqwyV7DWfguX5X0
4q6jeSQsyF60iM97m6x9rjaO2bj5AedlLzvxOEIZTUFwfiPUJt0fF/1oBuK/DeRJ
9Ooq5+RNA3gTjB/4Eppiz1N+aTwfXjoYfIh9WXgQkDJ+M/94fA1oWSRcjtco1fhX
vNE2JbJ480EOYnf1EOhhZNBlM0jcwFxWQOc47iNDCszjvKVmkPcbC89KPpjriFKR
uvlas3SP3/xDOWEfqn3pkbb9jlsEyFJHBNcM/150T8pWnUAwQBmKy0r09QYp0d/2
0HjJwUjc0XYmsp+g/n9Mb6wdcIpiLCRix4uc+UPyOCcEu9jk24jE5pLlesIRxXFB
+k73e5Sn0LS0atGSozDW4ipIrlwBeHpwgBnc1mJ3V/nm0XH3Jsa+p6vZWxjl7MQv
KFrjdiXFGNuVIvHBLWji5RCs5rFdeZ3RWmSmCGWKInZvht+MBJptzBkw0nGqnGeQ
Q33bGDU42DyiNI+2MfLes2scwpivdmxrNo0w6zmfmwpVLqse8DvR0VbfaB4CZCWC
LVCNx66EESgY8YoEbRReXflmg68EGiKh1YTrIclxIOIeMU3BuicNywmAwL8ZDNAl
pjkoI7yd/XrzwybRTvHqRY6MfxKOC13m8043s2FHhISmUWvGfsvWzk1WIgnm3R53
8XreLvKh/SXh3ZK41GN4QJZglXiUIgXX/pU4q5950w2TGLTEknB2aKgJhQ9nmQ+w
SqBJTMuQzO2cU9CuJylRHd8nNBcwTG+xZM/cO3xZUMu+VyjaZt2FszK9nWSe5BEP
6MysHroMakXWxZzBSi24y7yNMi1Ck09VgXDOZFcJEZxDZo55SUxuDFe+5OkMuT6K
djWHHdFzkzr6nipyDcn1D1OesKl72RyrCfX/MrKPoBt0k+PgRUmk3hRknEBkfVdq
GpcDlGKkExYuj80tfABnKNlZwUvkRaLwuhw6ui7x56CJDUVL6kkXfTLKwfw8MuxJ
cmTVLX0PqoCSP031bRBNQ/zUIoFtp8AXNcfFg4yZrGOMRq30k1zpwkFePVH6SNnm
u83oOZkMDwpf+U34gXhE+eW1CM799l9V/U4HIuahAvqxEtRyemIez0d5dQxRbJmn
QzdGvmtcAEmCTwcHfgZ5LvwvZhJdl7SzYVQVAY/ypuWGHUqP5I/8c9jKNWUpQvsA
TXCp7SJnP5Jh5vYKM6AWFGItWnvRBVpmRr85ghBLVqYWqMJhBR/d3z/Q1SAsdNMv
Y3Qq0k7qfmr8IGDA6KMdDL9/gYokmV5dUuhO+IaPs4abLtU5Zya2zPr1VFnN4Sey
8n6xbJqTC5/6fiqyC+ITlzEIBOh9t9iNdJYIl2d34OZWueYE3TAwyuZQDrVF+8RT
eUrx0BDgICuCigA2ZAngii/HtHQ3hSTgqQZ0M3W3Ec63q47B/HNr53IFaliTxlVL
rSZx508glje5ZUqAvDQWEiNBpViGYZf7JhyniN83lJGh1ynXzQ3jSclEOcQdTHth
kvQiPT2ImiQUXb5L8DCfLYVN47rWTcmjkwHYkHyrV0p5E/tU81HT8LR3ReOr/lLf
Pi0UfARA1cAeKWwszWAArXGVVGeVD8aiFGp39jbSLDGl36OQDxt/oVzpBmGAcXH1
bPlZqUBCnvJ3727ILDokyLkjweouuHpM/ExhWQjPXhz8uFaHF+X0oy8qDae6dWZq
6l2WaU8JY8CoYO02vHwlAbhsbpNeh8QHMtpqJuD6WDct03Z2BY2WCQfkssRnBXMH
hkFhSrQShsg9J+cH+ewUHvwgSBTM8P8oJPLfEhMKLnamDgYtkH/PSaAUtQjm9RBa
Tcal0l5zLYJkeydXTxCBuINsOd++HLkt/5jMQGkfB8rv0FIsYdIE+v8/DqG/MTLR
5nRrTIAbDvX/DiQDija1tYInA9DwtRoO3XaUw5csP+3com2x9qePPJuHRygIC1Ab
dZXUmat09dFfSDsDbRGpcj1xmM3eo2hfCFAaFFMJPdWr+hyKzQSSxnvttStNKPLj
dpGlQdQyEnhRRHVba/jIrl+jtzUOrCy1J7Ab0j2vwX/O5qV14AUxCqLB4LPwL4sp
dD8QZTgxWoKcsbFliDbKGPqnHxjHgnCtCL6NR/0Qy7lEhFONx5LtOoqhNNAlToQ+
Mqa7twzeGsf0ScShykWPpiP2sLelQnMp2o+6ftnute+Ls/0SXNvl5IwZ6/wrEu0t
RosheoqnxWQfL+fWI0aNPPZswJ7INTuMPvROwmVzp5o7GPMUYXEJT49XubOj79xS
0piLDI2RJwLIhvVr6pG53D0ohY4snTWOFMMxrNZ9+nm4cMxy1/PaxZOxm/CmF2SL
Fo6QL/orOt9FuU3SUCPi32JDIZ8bOkixhPwvoaLP7qMYb2azhso2CCTNH3t9wc/j
srRWu3LHbLraP6BWfaZN+eIHrU7fah5HEw4jyTuqeTtdH6mXWbTRlQJWloRR8wq0
e7eua38h76WlQqZt1hWopZo4F079BjR/Sg4348KHCSmev9REL4TiVWGHxl6n40OH
+pQ0NzlrFy+XofRLyDwKmXYMJTUFZUNfxS/5SY8g4/k60XU2n6qHJERFWxY94m0W
UBGgmsqWspnb94alFttasgZL/P/O8x2qDY7oz5gT6cSvr2Fj46oUbgO34lsGitpo
FIJz4eiLm1cCWw9fU6wairWoAa+oBx3t3owbW7ZCFqgOIzHHnOblRieHTleNwe9z
9Bmg/SnLNo12uUkEmJ62o5eAr0wcBcJQxNj5Z1++ZS5/XStcdOXgAx8gNxJOJ27b
L6DbLaEuyFbmGBq2FbiFh4Fp7yrrT0tzVvZ0wzxUTAZE7C+Qjdyg+qPsd449R52g
krl+6K0f/WH+4NdBjA9GAeE1YSIID5JiXXjAm+BDPZ96mx2fBjxK4EYTz/23Nd0J
QrrLBGLUj0BKhYaCDp0UE9bJG1GvYTKmaVPZ2fs9iHsJmnlsIElf97ryZhV3kOO7
4L2Hxm0xJbsKFcqtor+elSbC1bX1CasI//qH6xiI9kuG0IhJqxrXonxuQyK2wYSi
0stCWVM93mmCKkc5mkMmpxFQZng40GuElVlS8tkmanp+UQBWzHuGjcVPgup2bVkm
h+VlUAqM6EVhPq8B2dsjK3xq/QtMZA40CM5XG4+sjYr5TlZh7fegB2nPR5HYhvRM
d/7Z+ge35iUzcwqb8vELLdm8bzP0aHIU369f5mu6H6x8tzg9LZBu7ERloEnnqJtx
ysegP56gbmLxwPdM/QuqaJORmYDXKGDRZXR0NPscrEBpb3x2XuzVEYpLg3O96Qa4
QwyzBBOSwAhMG4+v9NkzAGDmtQSgt0ZnjpRrzcjr1i79ll2kZbAr+z4dGl2YFdYj
hPJKTNthhC2oZczfrg+faMjCZNxVosb93ZST0QiQaKlbpVALk/EdmT7TcStpvu9c
2Wm2L3T8lUIBd0gDeQPquFblF//QMFyng9FS5iX5aZ20CojfOmrg4vVWbrEElnw6
vRnofDzChfWbBiRiEw6YJkL4KiAp7+BCCh1Oi75cWnHP5AGxSsOF5vQF5P0zm04O
43v/anKOtcvFtgzB3wl6D/ASE/KmD9bwCHac5pBy3l5vspJA4oD/PkmIUSD/0CC+
6pn0zSBlKUz2LL5J/zNyfoRGck3PFm2aL6tGD6T7bkbLhwPE7oOK7i5yDQUMVznc
DRYn8YiPuS8ympgBTpgXgPpMsdrWBPebVSsPwHKUS0rNS+T35v4BT3RiGqYNh4XE
naMucHO/yUut9YpGAYYE3bpkDD6xnp6AlJnGfgOG1Ax0AZCj1rVrWJZnDI07aQPb
bZohEVJsD2UsdboZ0RLVHpshcdsNcsOFQqK2Ta3Y0zBsnh5Jfg8LoxttuFXfxbX2
dbLFFGlfroL7K/9Gi0YLI4xw80weWalhHHyNL31ziHujnwtOKbMslkwMDEsSYmJy
NKB1l2zLPaZgRo8OzBq152SOfuwjBHX3KetUZJp/exOodoTPvH4JPffmH1l5YUY6
HaOFyEfGjOhrgSBydDQLREpIQ+/GQrSy58kcflCS0zcsMH6aR2aqtdVhLOYw7Vee
mcjvID/qWxDLjVVoSX9c2fd11dlUzBTWeqvR2sKMWBsB+FlVH4KUsZnPctNO9Ufu
hEy0Os+/pMx29BJ/k2UGymuiS27cUwbCmhJCcJfg0db0GC6sr9jcynIXguI1qovk
6zEc+VIoUvEdkIiZtV2ATyI34lVPjatpLPKiFWm1LFTFQZJkG86OhEyz4akwVyM0
Djv6enafrH1APzuls2APdlkivOgXJxQ95t9xzp+isBEytqRlPCO9+wLUpjo3CkPD
0Z5PbPGNK/VMakdpLQCeeqBk6GdSwQDv0IgDYuly3D7kkXuigdFzH2qLmhWRG7eG
Bm5UwzAP72UvcDBXvA7DLYgSG2Edezrj5F+qPcqMhKVBRL8CLC7vbjo4hchBliaW
xqFw24cHJ30oxg8KawGTwNJo90jwDNk+1z56JRTg6foaq9oQqD5YA4WHrugt/HaJ
S7WPyRKBS9kGPdvYX4kLp7uDVEgCMtOmNDRr4Tv/G8CG52QHJCxj22f+dmFu5PMS
XqS/S2KEhmDGXPbXn4DFBDXx6MhJQD0ktC5ctCHsG4MrBC6GtkHXqXu7r47UM8AG
y/86D6+lXqoElHFRN/8OeeLwwMfRnuGYDebMH5iQOx6VAC+paC7rw/18tkK2h7U5
nVV6b/kUwHwSiA21VfePeWqxqx+ZwLC6o/3YaKH1FnsNNkp6RYmZoIMbxyJ9htl+
3vhPElYoqHigrH5PwcaRPKXeWMbEJ6vZccpkAtQiuKIfnMMT3d9HMo+1mvuBL/po
7UdC11mCyLz0cbxNfDAj0agia2BdH0Bwzt1uXa10eHn0y+DTTx1biYlbwoEFnO4d
2A7Nu8XQAYr8cBm2rXxNAY5VBl9AjhqFP05hqOBqOgqG73fi/q9Irveg4y92G19J
l96frVQA0GsN/4GDm20OWmipvB0MaoQH7YWD1QEVYCMxxW+dGEUZoNB3pqAFhyT2
hAMDWGktiOHZp4AS6ksyoidHA73l6f0xu91PHZHSCd2MwuEjWKuzgPWxd2cFnhJa
QEMRs/MPfCPBgiRlHAhGFh+n311dQoJ1Ih2n2W9kqp7Gep4llZBzS79+gLV95oDX
eyMQUJQZ08x8Nr6DpRVaz2RnTTgAexPGBfb4xD/EF9v3a9XTeaA6CjNnzHvh8Hry
2LqiGuFSOYjdlWPLzSCXEUjCbXR+cL0qr4dEkK2L/QtOoQmVxeXvZW/cxp6rZo9d
HJ1jPdkUsd/Fo7WP0UadBCh0k2CukNZB5a6GE0J7HjffIhtWLexraQCO7Qj6Dv98
GUDCW9SsFTsv4NwLSi5UllvlOwZCrvDcdNqmVCmcFdEv1HspPTQWrrkdVBI5ZlMX
7wsI+/437Hepn6+2dGhmFxIVI4qzc64yTPDOaDSxplwbHLjLObwBc4zIjSTG9ILq
9ZzsrtZ5aNHmQ4InxRFw7N+z3HT4k+mOXzhCdZt5OrTyvXorlDTVixLD0NyeHkpT
Qq2FkgfolyEElD/vv7FMRGrUtTRzwqAnonvDZPvwdZmeeJyfjCf1+1otzBGLPGaM
+622pGXw0Pi4A8VbFWqgQjHhJwHzhFdIvZJDFyfHGW9oBOvISSthoIsB89iadGWa
EwtlxWKGX5jLxVXP/eZGGqjNvfHboAxo5lkg5oWIUTYZzTeDqUM91s5NJfLJenLe
Rh3zqGutGcsGVfsHYr6+5HPRtHAHEZdsqc7gAsWgXrjksBP55/V/WjRYRdFIZTzh
0+RPmEt2oaiWVVuNaFALptzoYL5gWUJKgXDrGxf47Q8400Uw7fopjQOgC9Gw8T1L
fVXIMucFZmPrPjG8hWiZ7bUx5lPRNonkGZyrS00P4052Ov5IdSjjUX8u1HIxKt+T
zA0xpHZkaQbaOyDNuqf9dDaOgEOk9z7u0IVtNTDmsMJdkA9loxiWbBDRdld3ZxmH
Ayr+1oB+htZVvpePHaGZ2d3p7QgeoTMV7T9i2reX1N02pf5GgkVOdg++GNbq7Ta9
6kVT9fHUHTfIfxyfQway7l4VNpjasYhWts/QAGXglsgSoLjJo+Dmjhbn+fezdiN9
oYg9qRSmWdSdEWxumtlT2Jn5ZMbzHmgKbbYzo1QPrt9WsL2tDUZ64jcf57ZRZHDj
X5GM+N146KFg96gknhnPmOiqIKKqQ60zxsa/AmzYK7GUjIFX29moNImDxWYE1j4G
58x4jgRds//vLECCBh61PD/rcZmR5uZD4qPj15GJtxSfYH5TPCF4tpHKOmw/WwsB
NzUqWCHdZLODxHrqjDVOWx48D+g+IfNjLqVfu6J6uPfCj+7SbSK1e8x2Pn9V5g/m
V5fPZZ1PP8XKFBxruzXDbzfyo56jK2rXNOTjDZYtnZsYJxubDNGT60u4Br2PmSfv
SJDVCUMBGLXrHy0HFoZ/PpSIYvRD/SMC0ZOx+8t9TqxwfzPfDlPeZSLuuPgUJsbf
tPXkOAxQPAo9n4Juovr+duT9fx+HoQNqtMV3FBIzimWu4GrVpoTGBp5shr9x6945
rM0ryMitSoJUtUvMhTJvusTyYx1EuiSP73vl0bwpkPSIhHe1RzSvq4CA4g5axZOw
Ocfet1259E4W2pg17KY5nPyn83/11NAX3+gAWqTu3ck82kkcxuHy08oyJilx8s4/
z3snCD9PdoY0RCznuPZw4I0DXHViH4LCcNJQRtBD1iCe7/3cviGX6DQU2gyyLH+5
Wfpyu07xow+9q5/nkiRszwHDJ8DRE+PHZnJEtpNIreyZ6ZaYpV57M6HFFtDDh1L7
mRlFlOOTYj2j2a2YdIkOGl/K4F3CiNClsnZZ8fZHxn38bQ6hekywptNI2f0lvxpz
IsKHG2LXS/2v4CTnPi1BC9t6709eU8i8FZvKZSa5ryLL5lYJPJZ5sjjCbDjrMw+r
bfLdyHgs79/yVuLB1wf4VkEAr0SHjk/NaFWx+JdRYlvl9CN+u5LrWuqphZ3WJHrJ
SHuYLjIcSJdi1mIKoopjcUf9ORZLiMLeiSX5cgGp3bgpD2BuTFw6A9D5dlaxBU3U
qLYgHsU9hFAAA2PeMYJuwDMaSBI5+k2Z9tA76oDUVpZ87WS0XkO/GyUXAu+D6T57
rKOi73GEwT6qGNfCK9ql2yHPW7Y5aVOo34rYWI7h7UriAPUQQtOHOUaawQwF9+mb
mm0MTiBCsZ0O3x3T8o7JPBdHrKhvRyeKoZ3dVaNcge09kz1o/gxzFaBN8ju8p7yk
dymbyOncOq9uqzzb5XHpwrIpBUTsBOyNElcCVipoPm9Wg/7MXWYz0k/QQzOtOQ4n
w2ktEYSb+Anclk+pvXfrMIaMZAuvtvMHHImgLgbTXFxQd7Z3Yi9Bw/spPyFTCXHJ
2BTM/4wDjSrmLPzv+/ypOtbNZmCgF16bpci7kALOAEVy/bEVx+1xU844gsQ2V4Dz
QzRTEFxjF2+zJ1HmwdAhl3PWcdd4Fkvy04Hjc4DDred1rlTR7ic99b1ANqS+Hidb
U5T1Y6zcDu8ottySM6ydpxWKfZ4jlY7HxvC91zRgU6Rh4sz6LynocwBDUTmixSv1
UIb2mFsWVJh3jXi7oJoYUczbGzUD3/z/GYAfuSbdFNuw+jTKl5mmjAmCCH3Q8CdG
1EMauJ3y3m7nvgrrMrl28A7XscoSyY1kjCZbulMl4wpyw/6BkRJP7cccOR77GuJR
WzlvVFNHp4hGGzbXrp0YIsXk/eH/BK3fbLoSHXqiOhjwjaWJdm0EZ84+MaP6N41H
FyhR3bIaLrReAtM/xpNyMSSuA2T+Ls4ne26LO+ZhfiFxTpqHw85xcUVm4PMPeIvR
050NgPsNAOXCL6VzYoSzDjvxYP69rFXLtax6vk3YoaD5X0+GkzI02wz+oWRqIJym
hAg7ul9MQjGzEoknLX7ff/VEki6cKRAk3+4xmtqgm5VWFmHP/C3xLLmeAh/aO0au
7I0S7kgMFLG0CaYkFjVbfQrzu7X70Nbyt+3RU9QQPgQq/GSNrYvZ2ejxiX8owFmd
/4cIAHsavHldwBvEcAor83d4hNByUckuwUbWwOVefmzYe3YdxkF+cGRFAzTRZi0B
o5JnjzxlMlTuyp1oCGCBiAIBfgKTNY9RvzgKQ8SZbJSdIXKlEolbjvOwE4LViZQJ
d6iCTUuBSmlyQrIjHTOhQ0fIWPAsVb+TEccYvBQNKV1EgC9OkQWTpe6ZZMNFsoO6
Uhk1sfrtlMaCPu/LlZ/TOAVomnZkFVpL7hYHNpbtDrgXAEOF8GnOswxOYTb6nNpR
W5DjXCNklIrVe+uVM0Y/k9Q26wODKO0Vz5eR4pW48Mhnxr0SZ0w/cV0Qz78Jj9x1
8dIwNrEoCQvOPQMo1CPuhhFsypcC2cLA0e0qjSM2WkRLFJXt18ae+z9JcI3/Wfq7
87Q5UaNPsuIkjNoO3uITuZYkDfHZCY6V61CEcXfvjGAaRzyoxC7jVxtK4BTkawX9
we0N9YJyz2w4xk6n38T4sGcJqcBY1B7wtipqX7WIsWjCukM9LeE3E/K/gr+XI7pY
HYSP8d1ktGO+RH4Utt/7HSy/INFjupV7FY4vQ9+DP6cz1VBzHbQ3e+SpP6yHsfuh
Wnxjs/g6XSVrGIYkLFPOIAVwouFCQF3vVAM8C4nLT59ryTniuV2vh3NhDn8sJOhX
F/svXyWlU9gLjE4SX2Apw7vmD591P84jhmnEUBLU1UFVXFwM3NROvhaDgvWaInjH
7W5wfD/1mzBXK6gk/+cSjuwPcdWFK3vwBwbiri2XT0eLoBXZjj+9SDlzXkCbJVSS
sp/c13ZLiIgRzTli0FVnweNrE8xT1p0tslrLUwMOcYZ87NbzyvP9qiAB4hzxwD32
nFc4P4y2MjF4dP6ByyXmO04/nZRa2a20TmKNoBuFube0+wDB00kTnoaNPkL2UhcU
KjetgiaslxezLyFrxo3UivIDnmXAhzPRpGNEGV3qimuEgSMLjbJm6/RKz296HKne
os7S5VXcrMCA7vXkhSYbuUH21SMVFL7F2lZU99tbzlISNzpXgujU59ED7U2ne7Kt
W4WyffOPExlnf/KiAJRFUucVP7zh8MEO82AJtBywiMUhrRy/qPbfx1lvRyLuQ2y3
qLnPTJIuhobUk+fXPpSKmE/iojg9uYbRGDZu4/zxa/Qa356hI318LE/WvOVMlbSh
mgMQtnuILrRCgCJMf33FmjPc1M6DRaSE+Iq01vTUGprXUFl9DWk01PvMW90l9Rrw
5DiNAhZnQ+us8HTNMSJOerkT67gpvkCj706txwYCbza1CMEDAV7bqejBdWKPmmgf
/Uw32etsA/KkYsBo6zguIOSCx6CzRRBfooCBWUU1W5AfRoKS4uWFH+9UiS+6E3DB
m5iABMezbrl8yQ8lwtnFtEowWj/rO9veaSjTpg/9kTfIUmd25xn2BJgKkBDOmaCn
8Krc8ALcpqCW4ASHlt5FGHbKNCGkcVeSvoZz1u4P2QGnpoJxgeHCaP2+6WbYII1A
3BXRAmu9I2Irgww7gjHa9ofqxmphxY2SqeNkFnoVGDout7evlUdfWuwd218/G9q8
E2BXhFcTDCPNk04oPKnbY9xZVOmfU2Il9cyXw1g3up/+IvqP5kBqU1g/fSrIVbBk
FV4DK3y2TTn0sAlHtUEhBoYskGTEZlZCxMHLd7rKKpwsHfSQgjJG3UllIH/mocxC
jUSl5HZA5PCvusBbRiPUcO1EtFdF29yYmYZGrWDdr9ku8xMjV1lyxCmbpDSKMg8B
iAMgK3wgCb/UeQ3yGJYoTzduzSj34IJ7ekEC77K3kny6MQcU3/7abR1gCppxGpzT
c5jliVMTfy8JW4hoZ+HNOK0Dg9vahfEW7BdHQWwCtvAnPkaamPuPYiq/lkRUnsyg
vKOBVUU+0YNrq9qJr5zRNuQGlL53RncjbwRfz1WhuYaKIs08FmrBIBR/5zv7GHEJ
tiLDVEea8HZxEgSkKSzBiIi3cHCNzayQSeFC3uV9zopeiaiyxmY30wxiFUxN1oQP
BBYX5fWtrBiCi42TLXNwb/jCEfJ1goNp+pcW5o63nzC41f34U8VyqvImE74mzDST
kxGDlxvJNPSqeg0yCUKROkx6cBJi+M0MPX2msCMdZzTdgxMWQrAuzUBOv3b9IAgD
w8xqjOJ55wfrpEpbSW63j8zkCvqzQnHC93YMGuqznIKW6uIoNGd+BLuKZblQl8H3
vvooOcGqORl2R8v6OqmSkNHoxg5md0xESAW4XKOR+pqqeoTk3sdl3V8iYBFPhW5q
pNSm8Qj8b1an/Zxao8rgopG+qM/rjDtwTE7fZf6fnLfjYXEiB61kT0TReQ4kjMUb
Wp8Aw3FntMC6HBttLNJ4zdJdNfB8zuJciu8JcX+OHQ1uP5B07ZjLqVSzq5LbzIgj
LFwr77VlB1EX/vSb1HBfQ4cM4AJBaxIA7FV+MnoKG0RiCh1SnrXCTAfTYKfFoqE5
6f3vEg50ufzPzTWpIoic9KnhXv9E917ikt8YVWWtHJuF3jNG95t0tUWk3lgeLzga
TvloQrR8ljgvHV/2VqH7VHYcUYvx8z0XHm7qLCPrVU00GOB36m5dQc4lJsxtI9zh
f7Ur/PVkRsZ8a/dVTyYG2CTpphQKLmxMGzTPpBjrbggt75Y8Bh4FeZyVdEIb91uh
KiSbrJcv7KY7FM9JIDvi0KxzVe1OwnpmUyksPoo+mVmSjJv3OkSQpW7BbzskkfEI
hHs2jzdNP7kECUTS3fnoto45zun9kVQcce2sQE2btvlgzXjnZGPRjq//k3O5kODy
GQ6XtmTY3RLeb8x7a+5LOd6i0k6MElwpGS9uLIAOjSBFnOw6q1oFzZHXc+u/2iFo
IeOzv2KoKmGug9fCqgjbi12RtOWvF/zj7udVLQ0lT0Cn+GAYanshp8T6PQ6EuI4Y
w8uZvQPzAsyYdujvFdqrTwyYHgMO+XShpx3OrV+TvegoKYwnZDy/Ly6prN4a3duZ
wq9O8dDoxwWZqlbCLV3JTFfGUA5wB/dpudfwLwCFnXDZFU6WPbUO5UeFPpBRdsjM
kbGLFPDl3pcOXZsWnreLG8kZLhbEkmX/ng0O5MBTzMU807Sm8upe//TD1/L6Nc//
K1Q2fd7vCyFGFIC5IwxoOQXaRtTORrJOI7FQcfFno9xPkaUU+U17fbwh6zyQUz+E
4SoDYB7NTPz5pGC8wD9RN5a8yp9t0K3oWL1u125WUIsWSCf8e8jcz08dr/hKu9Tw
K7OPML4OLnA1KQqLJS5u6wKEKFmqsEmCmLJ1MCA3J0RA6IrpnY3L/UIfOhaEjNoQ
tLdsq6nO7VEElFCGGSE8UpCERjz4Z/z9Cn+TAM1HnarWo1CVo01R1YP2X7v0h5mP
f2I0yBCFQfgw7D0uyIqNZ+sE9i2YPvuE33UahM82MF1qBI/CF0DZvbb/GhRLf3qF
s1PClftiHdC8l28kVWie2wCwBs9ocsg1iM1m5+uNoo+oW5Ulysy/WQHkYX1XoTcr
YQyCgp4fMrOjTaxRoFEZLSs107zQlFdXp+4iJxV1POLj0f5fe1WU+gJaorVet7vE
BMAhbakFBvEM26oVG5S/s1ce1fFom+oPWNTQOwDflTQTti6qsk4EMuoCBuaSFkYR
T+UAViPRUauEn6ZLIoo3QIXqXQiecf7r4yqG68pBriSHvdUEhC/UZnuQzeOlbaDQ
+sNVTIic4TcaGmxkib9d42EeD414qS5pNtNx8gxgsPKGI0ZP9xGwBck1dTeItl2A
Bin7JNz2DtmBzjY/vM33BJR0/GYeD2BUr48DEUCcDHpS0JL6QCMw+KgG7PHOdlp4
vnNqDImuYhuZxGCnk052TbAy+g2TpMzyfAF00yYo8sFiQ6qNHkL8bCL/VX9IhStp
BzqFNNy0sRi0gqQVkZ2x8hON6AvYSstMOn6ECRLSD1wEhHtTnZ+9lWqinraiES4T
6kFi2CGKu6PKGq0UlVb8Qq3RsghH2LXw7ZIulg99nkCi3aki9e4x7mP8zDtB+C4H
PPy+4uAEmHN2n4SpPt0fNxGwig+X+Fevto1QnwX4hGikAi4lVmxaVJdHwQw5UB/y
Hr2/CBLAN0VN7de+oJxq8B4MPIfJaALY26/WFxBsS9yt7rhtRVBE5Q1G1SPwxLrn
EeUPMKg20A2JRle89PKiU1cbqVx82NAK1BtppIFXPmVlpRysNg8E/2V73JTjERhY
jnE+u+olhlcAvF1ulYaeqjprL0bdTFz6vh4IBcNz3zONRqNnLzgbrqJHGhSAZ9xM
E1eqNDR7LEImqs+asAmL0y/mK5zDxZinieAbCUVzN6f8TM5DydbmcK4y/neLU0xe
4xjxbR/EV2cgs1pJSbdnk+P7rf01dj8zWXGxVkccJXvWhNJ7ielabkTjBO6Lv9Hs
JMgg6ffT3rPFCCYsVtsgUUAAOZN+8u+PHzA0BlB4JPAwLS1WxgrxDEv9BKMNpAeE
0wkqpZp87oNhfw86vuoxGuuBsW9BT9qLL1DXICKn+NgiRZhoo6RL6aCV6OwMaxfs
yOaHAXFuTMRjgVuhu+XFkd9a+u0sFqB0nUz6b+Nm+QTtOG6Oj6iPcTcMlcf+t/iT
FvHWwHooAnsvzkbf+hhDeTW/bPeiMum4qYbcZNkVg22M2mxMr0Wu799+uj/CAm6a
eTvlWBhUj1PMbmGjoJ5TBbf7F1m/8l46McAEtyn+Zj/hg1IC7BwXH8Ct57oesyZq
nrrgebmEJxbF7EJEueXQRJae/5sW2cnKB32gjPJNP71seRKFlN/VjaHJ9P52Yvlv
49GDiU6yY5pLtr+gFqVXFIsCDS/H8l1fEwcHj5Da+F2NgllVzTqPiRjeKVLTKDEV
0kacsN+SjdBAqtrZYw3TvVHK+RHVGkgNenrT+SUzq4iikXTVVL9bLANWNbUwobjU
pCtWOKTiv8lGVJ0FMoh/GLjZowj08G7mMzGyYUtKnGiL/6N9z3tPlLQNBC2GHSvd
QleQ4li6TYUThMFV7J5/U7yULyESE1LoR8B+Zk9g8bO7aXJPjpNmG05xJnaysGJ3
SgfoIKlG2Jpd3yqNoegJEv1QAovfHLfA5NLJrJ9VD/k2fT/mIpUBqTJmYKH4UqJq
oTWpernfDoV7YKAnb+xbO67T7rPhn0eikj9NXob3yWPubIaG1qpVL/NU2oMJamWT
PQhZR5CPlv3eH1b6zd0dFJm5V06sx43b4jR3rUXT6u/ShCLW5/AGm7Bk/qWWCeh9
kZX7aMgeJnEZNaaSYJ2Ecc9qXjgi23E3pQ5k+sIzrEAm6VSYKWcJ7ebL4/1RjRFS
xc6II5M28iGVbb8zHUUACN2PJJ8wVN53NrV8Z/L31rAeuNJrPo2Z41U+91gI/9yY
muHHnaGCXkZHBK9SkW3MxpdfMyIkKi4y5oDohmCP/LOi5+iYdBXC7Jddg1c66pTE
FGf1Y2x0mDNWVIoKHTof/e36YDEhVj6adRxGBb7CjDj5XauxgBxC1wWSEFRrdAzr
PB2uD7h4F2xAH+xfUzmz6WmgOV6wwHmkney2ju/owk2ez+7GOMwrKo+2KB9v5imZ
WOLxDfCALF0lOKDuX/YBzibljErPlEE9JtByceWK6A+wshC1ZySterNgB+cJiIJ6
SQq4J5xtiOIxB0PUGZul1o7ik7Kjw5ChdgHOCKFP5SpxeRtCcZUerRpoEa2zYg7o
42WqGpnEOaFq5RUqnPy6ASVPt8V7uIIDrSmpvpFZe4yeFqlQwMkwwJKx9aeKbKyT
sFrtHkfR1/JW0v0bnam/JSh2qfzTvwGHowvvtDmBSkQACF8mgSVnCGNtopYpEjri
fXd70nERmRz2V4qSZTN82cwR2VAtYA26th/0Fgp8PXsObWa9HpiLijlZMOJetJnL
jSIaOviSY7Ea4h61rGUAFQYcsx0IF6iyI97OB9Qp8KJP1X8fadlJRGII4saMVzv5
5bM1bk3N9xqKnchlT3gRikpyGaHsukbm8Hc5i1XvrUGp+V12ldgy4Cul2+8Q7IUb
UepSe7fcJs10IpcpPmUPKPgCAtn0zv1X2uungzR37Yd+LMwcsAPqFCwid3GBYcjD
AvJ5Bss4WF2OVAHQEXvRdW91FPgjQZKEP0t8v1mXkwj7mfD0WJlbarVh2SJ9r37M
V/53T3w92HcJr4CPOuw8LNGxva2myfIzHcQyRlgzqAReDzd/h9oNdjyvW8O5w8l7
yVtQ52bXPYPtgNodXSQtRrQJlqFoE+8hSi6BRYtskzEgc1x48rJ7okDB9Rt6kPqC
5g6ErGj2Hqd5DZKa/xhFIGgkQxG01vf5uku+9Cfcfz3tSfHZmQUJeV43MU0MCjDB
fZnUa9GZ8YNPxGbRHr3TYPQeaN/cmH/yzQdYCOI3GylSqx15kkUI/VbIg9U1gmCL
NCwXEWFmVDUfQhXUgt9L9ZSwHsTAi/RRyHDzMfu0D8ph6Zc46ZgU8Jn0w681++zX
h09cRtEvXNmjs44VyYq2+U/q6eeVH16ArLOosUp7MHC7R/VTS/KvGFCXfoMHNouR
pSJ8lnJM4RkQuzACRFYEDHFKCMz+itgdTGVXCAQvYmPo/5LDqM1hLJYVaHyX67WQ
NWCh0f2b+VvF0Yu2wBVMxJdWDsEP1mq4mm7CaFrkH4rWTgH4qjB2L4HzKqHVMQKQ
4gMweW6PzlDZ3vvChmLrK6Hm5zsMvOufzjwHxN21gHdY0hd6KxOJn9bnEzFLwjUh
hzFZ6L9etVcBFz17kYVA6bPriOZIYoTSVcawsYcQ6w1HTZylt2eEnzXd9SpGKdC7
xhlQDJkoyNAc9saiOQ1Zk50nF4idC/Sfy/7i38BAmdu5x6L/LptS5aQIgDm0zCg5
jHtiPkfWhSoV4TQysJFCITvfxQnnSI09sM2hHLHP/OIi77UAL7LRZPmSFErv9DML
Zh+zZSZ2kghoSMti18Kqu8ku8K442MZ2NNDYDO/Rz4ENGdsclII0vElNqJukI2DV
TH89C4cVxNycQWJs2/ujE2m1xyVFhIJtlhDp+kghwBsWa9OatrKrYYiy+QJUdLeA
2zdVZDpTXJNEhMmaWcgkbOMTd/Z88jqTuN2yNwXvaYSzqfCSy/Bj/ypt9ojkrfVb
Bd6qh6MfBKi6kak85vIVCKjc5v2oMX7fgUJvURXA0ydpzQ7/bbXhzkT6hqvj02TT
aVx6qTIMLJx1lXWv6W/d9Aq7bOAyUPYT8H1/u0tQuCtL1N5TLRbatAT+W1PIMjFD
b3T/8OWx3K9jcUa010+grTcCcEkYWWMvSA5qkhuyRdIeuvYLigUn0lvZ+jmXHfq4
nLiA5rn8dFEiOLsSSVOsr7hENHN8s+1ux7Dij+nBajSyxZjxgqH23nkHmkgIu0HZ
6cN45ewHyTabz9b6zhVcQ6q+Dqf9h2mdAWt8kjxqX7FlKKsB5OJxnnhO9epLeKwb
OcfGx1QC+uJmNeFqk6YQZP9rluEw305ct7EJYVv8SscZcGCgXmC7cz/2lPr2kgSk
WOatzohfhrM8ElgqkSvEBryZtDFN5MB9g13m7TuBg3yZuJQXOMaDF4wE9EMuZXs2
rYr3Nxw1m0+IDLn5TrldBlsPZBUdGyPThju1YtBJnYrJH6lsXwE4EbIlwXTsMVJp
TsEQllyANbdgP+pz24/4NxbvIc9uGll3fnb6uT/TzeqEaapif/M2X0Eqcw3HKL2z
+d3/RtFmyGVNBbbghNftKgpbPBEbM3GfrQ9TFl8CcA6x2UF8KKWlL2so0QbtbJT6
xx3zfqKrYafcyiLi2HZ5gXLObtCu+S+Iwd0AruQ9s7xHOJJyji/nhfYmq1KJiXmR
UMBTeKYWk7zn0Q7XFXvJ+0KYxeV94Axj8gSsodOf8teOjYEa+z58PNs1RKyrYA4q
vKNvXLG4YIU/7jlbEyoULHNF5mW1bYzn30OHDEMD0Rm9lSyxa3f8yO7ojVc32PdF
ae/BZDgzmeBooHbKAblQkH6f+HQNtunxl1Z6L85/57NDvSioS1ZW1SerWJWUmt5l
4vF3k/57NPanTujqLgDJ6cB+WoiaCNHXN8dacmsnqLOpoQ5aZD1/dmBXVSJX8SKg
Rr2t93yRKB9//s2sfqjuoQ9UXqsAVcWV1gWzuMUPqSTaKwP+R2LHLLlq2A73HHMN
C992VUn+sveH2LM5qdZrV0E4tVrM5Vmdv0EBSPNxatrvnui+rO7WUZNnsZfWDyZt
DelWX6zpdhJxWX/G0BqG5IjBBgDyU24yW3YQHE5EuIA9hGLX6SSFu/5garQ+DLd+
sB6uLC+u1jWXuocUd5JPV9qAANuSAqhHQwX3/FntvX57iqqVCG1PeEP6NrfgEalY
E4uQ2pUBogmYEpftyuUUmT840AfkObygWxUtTHbGJBJRogejB/4UYR3q5vwp3l/j
vuJFPlgycWSpEJGTZ48UoYDWlH2O6XGUynfLnYIQM9dFLh1jaNBSEV2V0/pulG+M
qZmrcxo//d1BnyIMpluw0HYKOR1IzbI+viW3GvCvCkrxt9kdpiUOqTZVmQTP0xhA
I+tCCYb59jZSRNDYB8uHE+xhOiYYTp+51/J0UeCOxfOecYmbqhXNvVJ0o8cCqRQo
rSji7hM9IwFP1WvT+J3goQFPNVU6SbjVsAV0or6QVR0SKQRw8YzjajZ1zBYcTNBS
n4YCNazBFJ1Sx6ymdpzOvl0QG2PEtKYO5WnIjOMdkxAKO7pQhLdYLGZJtlKYV1JQ
q3iJxyPVdDdIZ3zAFa34yRMi1L0QJlJI5q/ibM/cX+cjkpjNcdVp4w1UQ8CPk5Br
qF+F706nQlClGaS37pYYu9HrdbbUMo43YtzENM5J80IBuitewTW/nxfxIW2r9hhO
XwrhTQQTxJwaBZnq/RxM/6gFircf1YgLQxz7vmEzpAN7L7OE3Bxp1CEPZQkPGicY
ID6/WTTlrRA27LcbuDzVwIrGSfvPALdboKjZEjM2xPwI8rilEwJfyYPAZaCujckK
wEgVk/xgUB5ZVeaPo82cW1A2uhicmXoiZn37Epn75OL2wp3ye4l0mWEXp0QKnBDY
Mv887OgiXerxouZt8jLQl/nPllPHUXNw1U0Ja1woTOXxygU64B21AAhtMM5BQeDL
9ibP7T+VNdbuT8qrcagNb4ca7/yZG+C+IXdLAW7NwuKqB3bGJ6mCsXKCrFPqvWzh
yuX1F8pK/5RlAFv/nIE08EalZowlRyCs5RTz0bpAnYtE/kkxGO0ErMGrcxMGCUeO
AQR7KGmLNVOo758HYf+5FqiW9gWt0cGJIA63TeKP3JeS9ZOUP+39LMwtgeS2lazV
r+1t4z4u9sUElo1/+dHbb8v0U63wmVwkLZI901efKVmFEzssDRbaoyTETQge9RpE
EaeWSnwJJmU7vmKHH3sTctIqugYpLO0O3rgW8bH/j23JXGy6oXJhheQB27G0p3gz
LrQsr861kuS2rLpa69ZzX2PIAzkoGir8BR0AvsrAIJ2a950JtprrSBg4z9bpf6MH
b35ZE1AMxLBMwZ0rKKOcb13fAtkEbZCUILmR+3OoHsmaQqWY17D4RteUXWXonc8G
mj6XpWJTwk+AgS5KHcOFSOvC3pcJ+6UghfUoqRSjDpmEjfqO9DrasFQr7iFrSmlm
yNzPm8oHTEir6FYav4k+VGtlJfbovs9CvpOG7ooXsONgbBV/ROZ5A9r4jhwOeggN
gzRr7Etl8ciGPYSvLgvwG3kuF/IdPdPzA04niRPtmg0rrLwv0u0eUppitRoly950
/arlRHsPXGEuw4D/GbiAGaG1H0rA72R6C/Ktrvx9apCHqhsyKs8fWqKXNL4WYUo9
3NnFnT2MtsNXER+a3a6qDQCBG6FHJZmyONaTwTgTbYhWl7ikSQPwYkGi7f5taENe
LkFee7dASWDXzvoUF1ce+nd1mQbn/5mGS3EJ8Pcy5LHDMKgp6ZfVazlY9TeSRltQ
imFZ0KbTFmSkxm2HhKLvcax8q6T6bdEeaeuKJRXphv2rVIuUWq2ZDekMRky3sWgc
vNdcOsLnC6fsdJSN5OhHFsn4LYePssbW2Tqj7SvJ53d6Zl6C0zJc0lm97A8Gu94/
dIIT5E8FzliIxuLgPQsBKR5aFBHQHKgxGlqo2Ptq+DGwcTUcMe6O93rkYjDYCck/
OkE2VZtj5x5Md9XcDVexjijlcpRAXsJospUkrhaMUMDn3m/f0lIvKH+rKfwDpOjR
sbGfM7l8T4nepIspmEamA4U463m/hA6HbftZgnn7zfdWdlEXwnARd6hMrM6okPeT
yxlQldaJcMPqhbygmsmnElxiUIKxN5surbxDITwAtHSiTTWAEAAtKhhBeYc0g8Q+
61ENBQjxD4TyedohRfa5gBM9UrDJPQ0KbOFKB5bH5WAgO51lo9blytHJkxcomRDr
lEclqMy69XksCmsSlZvQtIx2g5c44QH1yDMcipLxCeVwMEW2GqDGCM7aRq5bo7zg
KL0EFtLy6vsf8N3b+N0375YsjxgmasRuFq2zxERPWlDckBAGua31l0YQRaF3OkqU
9GBwVZdMXXL/MpsG2gq4E++VUoSdT2gX1IY4ygmVYx1GqPvc3mj5djT2K7K+VzK5
Lj4uJzdKX55O/7p+J9rgHVMOaVO3ctnl6spUL5nJdpX3hBLpLs6QxVGQq8Uo65uw
/mBnEqgEEMdM4qyjSlX8RjnQy2Od1unEs3wYKm/ROdUUKOj/E+pp4FFa4ep/HkIP
2071JnVpX7z+hrSpaE7Mkze1rCZGL3gVFW0xCghTg6WKbEVWtnsbd7eFQG/e/AEH
P+J1Islm4buGd5B/kWb6xvujQjDPl0HZI6rzJQNBdwNaB6yiLjODF9VXpP65LmUB
Y3bGwCc0YhdNXuwPE0BEBL1hvTSH0CgagQ4ldR9P7GFI5QWFjvprReVPezJWnCHE
TYCiKwsZHeCbNbA+Kaa5+0Ij4lYLv5GUyMnVytl3ysmEJeH4ZuYvMV6QQjmJuROm
mI3fJ5KR/92EaOy8/zjKDC02eHiE4aC8s6xiI6aDPC8Qo1YfuxJo26H/Q7PZG5V5
hoTe+PNsz87BcP/SoGPMI7mYh6iPYIfeEASKPz82ZYtvUdhU9oz2j0BH811Hgn4U
ibxmngzlAGntxs/kyT8DfWdZfX/hbIVAxDCKUbNPy6jSf1Vse6uIaDQLkdaHb9v8
lZh1o6IspoT8MTeqKJOPEBrZ9RHnDKrCV+gkpNhPvgNW69lCD1QiNxKgbaFA5ciH
JIiYltwP4EOPT2sV9pYWCzj2EfuU9bQSub9CGE838ToqZ2UvnGPAunH2zfabd9s/
mVd+je6HV7X3zuzbB4596uuCN5T2Y7zLcC17Wrzzv85Rhfg4XKWyAJNWkCGe2whE
2LuAc8mGkIDbOTmiqh7RBumGFMog9a01K1/SIO2u6RsnplnpCk1hWtHaZKaCcj7c
X1s6BPcwRHRgFcmhk36Gck4aE7hrvYF4lCqOepPZT+U2eB6do/AnASv7BrULRgZC
HoegVTBaDm19GSbTY0mgHqPenLfa/gaZoEXsQw3OVVJ7zsWHIPGQAhDyAAWgn0bt
YwX9voXqM+euGF0QqEmcKa1R3Q4X9IWG46nEoyJy0gn88LDIXpw7PRZi+JGw4dxx
kJpI/JRnTfvmzkkNzkcKOnXbotQiIzi1Q010S0K+Lyy0f48Z/WFm9YWQBehV+6KT
HZdBSlDgAdyaGds7ODdT9C/GPvlEu9Jotz2MY83GFROov/jbmFKKFiWOmnU/z6AQ
Id3Ynq2s6mqX//CbKKmcNxXOq64a//7ue675MIoBX+R0PBDsLgKG89hQ1UPr5kvW
4JwBmu6VtCD9+TUv/j9VF62oNxzBmv/hq3AYDaZRnw953mJ/5LYtzdYyiaYNGPF9
EaKBOkF8FBAH+ZOzZMEU9pe1OeKM+cNgUJMku5HMy9do9k3y8XrYFsPEO9tJ3RKr
1EPKWp8CMYq6QE+CBvtInpgmRUvKNO3KwP/0UPXyUl40RDCJJbcAWBfC9GpUg8zm
EvlDsEoiqkujaF5p7jMsPvDwWsji73CrAn1k2j/11tyQOZ61Qm12duJZsCrDQ0p4
weqrOZt+0NsBmbPRkBIaVrioaIc9/OgpnkSI1r7T4m0KyJc/PghFYjM8+YDsW8Sp
+J63RSEElL+42tUnF+EfICrc1kgv0OimAKeFWm2cghbstpG8vHbk7dovI2y2SMgo
udXwlPer2b/gP8iegg1eLrXAC7vazMwXnCqutTcBorYUIqcm3yZdIRdEfmPT58Qu
fr81SaAi/41Ov67d5rPkI8+2bf0uuFCQQA2LD+AB9k3I74j2YhNCQh8OUUs2htNj
0+f1JcPpDqOy4s2HZCkG2uR9+T2DMBz5f4nE+wkT453+Kv7LrIvLDpl/leKeDpl9
bmNtUa9KMBXHruTnLN+NK7yoHX/BrjMq9Ql9YefP+k+Z5D2BqLMZ/4Y6L0PlYC4W
fNl5SJ4uNVP7aqPGOrB4w7R1KUZFEv0cWegY0Vha4w4fJZHAJyCepwarpdccp8iD
2j83xRuF65GFfLez0Pz3sHbxw6+ryXNJbvb8zuhjWA35iPOyRdCBZ8s7A7V7H+bI
j9g96yhOPelvIElJAv09Ao6QFRSfJ0tSUESwwyUGNiZghpvg/5XPFkBzlVqBOOdR
IK1wmv/8HxHut4vg7Kcl40/m26ow/bw2RtvTXylqKn7DthVvV2BuXEN0bs/AH460
swAQJ3OlolkMiEQfOhqNgqImUNTQhXRHXAGIssH+tEDl9Gmd+q4zIHiMlcFQ1a2u
ecO2pNFi8lSNbBOalYsybK59BE+qVZp2YsrYxuDxIFXUfZ8fiM1E4+RXlBjTh/2C
YCNQWJZE5CPKvXVdApDAQ6npBVojgDCzaQ4e++WaK1f6X9HPNJCN45Npe/hFdeyW
ku1dR1OxG3g3kJ1iYI+Ziu2t73hE6oNrkrByU9ZfUoYBQS/6d9YfCtdcTlRM7BIE
SxVRwuby22W2bICQFzAcu+GhpW6iPAyLgX6lf3qU1uD5ACEHq/As6jZ598gJylW6
WQ5b4IHkl/ZzevsrYGjj4q1OmiFtXavxkjRFmBYlNQb/Rfs6iQuXFvzEKPUSdQas
yO08Id39sCP/kdZfqhpEY3wkpHkaQQKbz7KSM6Gxpa0C3QNTT6He7BS7PAnfV+Z7
iMVa5PWzE0DS+Ntob8ZvHwXnnt9IqkB8Y8k/Q3+gF5h2Fqv6Nu6cMBTViDOONj0C
mJjA47swXnPl4RIMQVUiaOhCU7rIqZg/6vizPRTK3xZQX/i1l8CCefDviEVYHcPU
Ov/a0y1yOMRJLErAw47/S91Vu+2gtIwx31pDPuvkidnADesqUxvrfVeflOnvo3Ae
QB1u3rc1FTHtBh2PAl1qcjEVNsnLqoETA9LMuSprMHE4bHAfB4+CzZDt7VpHoKaF
afqBjoov5+Z+o0ylpqo2Ua2Cml0u+YQN3dZanz1+F7sUKxg+NOPNnIuMy0A70//i
9k6l0hovhKAiwP6PyVAOYv5HAw0ca8NHbsqZnCTdOnZDL0qchA/xZnvcNv6yXHKc
2+pwNwSrA8fuGRCHnC3+4VhfAWzmL4UmD0uMjvxMtsn1ezBK8sGkKdm/quyfE+S2
3AJf2a6+ssyojH/uVRJg3wP0xPPPlSrxVlFHPz63hN+SgdLBfDl+VtG3Gls0+sk4
ib7I/vZdx+kPdzUTxknM+TzSy+bM4B9E7OTCz0+GL0JCQFiCRRgVJN7b+JNEo5mK
c7mnbTNbYN1geBtFJ70fBIBDxcbKKQBRn2f/2mYfNTLdOEgOFyR7Z9PER5rqdOIh
LCSNzkdEdVXToUEbMDWIkb5MGKdo2mMy0KnNNRCPmcgahjsFa0lHkMFyalMp4cE7
m0ZrrPliBxhl3asOwNsoQ8bN+93Bs7c3btRz0Be4yEUuxl6uRalpyzpb7qka85P5
OnXpbMImJ1D+38MpJgHE+G48yttmZA/D6R/iAGB82/CaLDzqprxdmsxUphtn8OeL
fHZM0y7cWLAzw2stoR30nZjX905m5hevNV54y5tCIMv6MCsSW+wQcvhzVF5HHXys
zT/0eoXHhmi7XOc0y5eBWH2zpWUn9zKB+izDTmGbtnAZCu+xm53JGaVYebNQz8bc
4gGLgG4xjPuwgG6k6m9Z0cgarlW8aWNtJXQ71J/9Lfz/7tzha0xYhcWxGmR67b1N
EGL1yqVc2EQ8XAvUCbXrNec3ttl6xj3FMtZXiWef/KG97MZowdjpSjewqaglzKEN
5erikuNxWGPFWTUukpK26nCud4g4SIfLpkdaxtqVjZlx9lrRNTBAHpUqjw4B7jCt
2l1/qLHfAAQQMmp4R5WpgvrDUi4WmbGf7Y6AwYSy2lhHVHC6pv1r4O/uBjDpo+wJ
+3aOjOSAXkgeqwbHmT0sz+8KV5y1HjK8SVzi2sKbU9xnq4dTxblpNWFxqbzCe2h1
owcWzLsrrDptqTr7Y7Ke4L8+9w6wFoK9odiQU+kGcXyKaUWwf9rgH56Z1L2IGNwz
GyDIxVkdXLbs4gMdYlrRW6nS+y5Uwgxml3km5UDdwCbCsl/StQAqX6q7CkEq3AHL
Wi52qS0vCrD+x7MEzJQ9AVCDKvGDfqNGvNIq5ggBtXWTQEW9I3hmyndILcxouKn/
L+C5KFLvt6n/9ESBVvgoDTgdjdgUvpXJ5cRNKMb1ojnN5lBiEuAWDT4pSAG/wF10
KDpEBcmCtC4oRiJ+5v//t/QJKx78p9ITmf1yV48JO95v2smJ2XOuzhQjbNd5FLNR
H8zPRnHEFjKEl43J4VhA2NjKWtvjmKbxHemJDFfdYSETL9Gqef6ERPxk0UqqnGIL
bW5de8IOWNWV4/eYB+6ko9U2DXia6n/OGFbyOS7Ah2jRokf6y1YS+YSG1dNJFtu0
2SUscfagehaSjj6nDG81t+r4q1qar7NxVoRxumjEDW+OQdrzPBTLuxSfJAiG3JGj
kkp/hK1pT7NpWRZV+LpX6QS6dEM7YhhJyKUnH8Wp4gpaAK9GfXdelnEyLaTs3+kP
UBXN2i+tHRUuaE2MEUbma+4x6flWcsSQJoaa6emUkDZddXAF6ebEHmM4ZQLF+QWB
L6ENrTUUSOoLc4iUalwk5aA/CL0uUPpOuNBJFbboDSshVQ6duXSEW9vACc1zSQwD
7Y/+skz6W/dnFVTGnNjMAXf9zm1KHPdJdG6h7c4q31lIqZZGZAPvkSU/t60VmeNt
aaF6YnL56+IlXfQFbKsSjOtm5nzrGkmqr3S4HQ1j2L+KQV70ybOTP1BtvIvNE11G
KU/1aj0cpkymC5+A6ghA7wWLkP2eDHEJhEQOat2MuL+M5guJbcegJaXN0mXV8W+q
mLwwamFgLOvoq7P8KnRxMIq9FI1oHz2TMtAzVGRBfD4TGmtSrlFQEaHSYipu4jz4
zoxwUvXk942yxabie1U15a/fCF8VKJ1ecyNMxQ7qmNeRTr8+OULmQfUp8uEQFSaG
vwa2p65PrU2ikt4ZxWLEYh1T27DzfX9wjIFETPIGSGdZilwwI9yP3dUTRim1VmVb
QBRdr499bHAvKY2ga+32+HlnOwxuF84ypYpWjF0phO1Hw7x8CqSO2S+b8IYgJAG1
ZPZqsB+6YUFN8ozoMmBHtr3CBDuTOykrcQUAtRpYGV+BfysawAuRA3ZJsYNR9P+z
yNhMD3INg5kTpYCYUDGZTutiMCOyvsmXz3XLkkrXnqMKoTenD9/GR9x5SYEheZ7F
8hQt6BNtEOagXCII0YE3kWdgaIiUSkIHzaUk3JDa7dP/jcIgWBCgD6knsblbIzAV
hoZ7TEqpRr45qJKH5a9lCt2mkaJ+LFg5evSyAuwpHfgFDId14YhQCSk7TLFYT7A6
PpYhSTw5uA8VWs10JbluaH3uwKxsg8zEX05Zgwpha2FSsCBWK2Zprbq0C9I76zLS
EpGWkl5vSizvh3DCc9YhG7KMiReNkC3bhoX2+1mT1AIVFljwEqM67N0qgITZ+FC1
Qx7b915sKNh8IzwRwtfDJ+gXwFypBdjbCRAgXnnn0mkjUzJ4LWngU52lTNdKXNhc
1Aq7kUanxgHz4v5KTRwjNGwLhTsY5dcwfe7Vx9Ir+AxKHMDHQUQ1nS4vwHiq0NOh
Dig/aGQbomooyaCucsEU2KwP9SzGpxYjUa+xxy484/tpY09MW2e6/K8Mwh8qJ8d+
1Ce1oCbBhrSgDk6pZKIhC25yNJMUnCpWuIDxlpBgJ9+o7TXlsF91+Cly7A6pa2HJ
FF3JTmQxYWtiMOBXWYRkE+5Gjq+27TJacvEMx6LJkN6qnR7+fnrFu9oYAJgbZYQE
y/fq1lPDdID4i4B64ZufSYNih8Q647IQnseFRNhUN+72aNxP58cTDYhZGVlIFOlM
ptMDVG0IklllxOVmCEPKq9asuR29F8MBoIYgqVIuKH37zNav9b9qB9dvCMyfUP2B
Wpm2w/O43PSk1VW78IlUEwpWXX8IhTizFZGdzFzJnM9bsfeGj8PrwKvmnoJe+Igo
MWbIIA1gONIx/TGakoJMLYEUuTeE4nV4pdpHdxNz3T0Vbv9RloXLvF+2wfuv100t
2HdqkOYMojGVfp5FFp9VmerekUXoN7d/bOHvFwlEOFBDNo3yGXq99h8UDoTL04dL
uW7E/2DW/ueCz4xrek2yfudBs4EQ9dVm1Fx1Sj/8/zn29AVuDxItzAcymKeCpPm4
26nnAJhnWG/sWrCMU3zvPGywuhp0b2Uh+Zro0PLTybj354WyLFXLuQ0qmA7JhCGi
w9Kv+1ggVgyNYy42mQL8qjQ8vPu/2grZ9gbYRauLJlwW8mzqeK+KDoKiPSg115mH
b3fJ+C5khixOzKjGntja91jZMontAiQe/aNFljxRmKvsUBfGEHPdTf0va7tgVgXZ
o9ctQheEciHABCZT9MNk2pZzjE5a3dbfm+swTrmosXyp1gZ5xMfBVhuu9IVCkKjy
D2GDc5nk4FYI8IZwNrbDRgprCsEihTs2jgJ1a92B9be2l3zSOwqufJeaDl6yVnKs
mgvYNZUW8mJP+gB7O9X23rD+pamqI0dtzGZedv4paTldAglqdNUKA4xPrJrYhdrp
RC1070zLwupvIZGrwpvp1ESBqyFsd+0Yy4PC0Ibd5QoG7gUQWjlM5or5Pl/dIHfk
K79YIWkvNvNhk1zsk6az1Bdlfap42gsHDbkPDaTOS/WJQQaKzQBibG2y2bm9wFl5
R9MYeiah2ces+YyK4t9B9NemfDpqmUhRyigF+6w9pyPKavUYzsotzmMmWsCpuBvO
9H1zmDCQcPwTEhs9Y1Vv4bTa5r2wLT8VDhJRZWOY5B8nnq/KtCRTFRg43OTZDhca
Fp+GEOFv5hWArA4gdVdMkl9Yhp29Os30HHZW8zgDOElnGtZZWjH9HgQROQ9lDVK0
5TCNkc7oX8DjcjzUllobtFGOJzwIa8wV47AcBue07mvuH79IcB6XdGEZ8Mu/VgI9
aCKEMyK+0dpHulKhoB4lkvx0kxnhgX3F7pjdqg73rumoTiOdodlWjFtTWqiuzIWc
AejX2pT5zXTp43W/E6oM+qSmlxVdrrlm0ze/F7LYoip5JBJWIGZKjKr/cNE7YBnq
8OY9QO4M2dG8n/r/ZKsuz56ovFS0LFq+QPxipdZDFrQsa0tczQCbG2cYumYnRolR
O7Zx1sjyMBUKfO1Hn7fTsvlvAVwU+GtMTZxYnSAioG2kO7wxj+GzIlwulQ6JwXJd
tSTXGUx91lyGPKhG6F1p268x4PMYSYAZ/yFHCPs9d+UmI8LS/lggeOyjBl++ITH0
hlEpPjPNxfOv/zly5XXWHcuD4hPEnKj2Gqhsg5WKPaIVpuRHWI9ZTj/ivROfguyC
yWGhaMFhNu8rFJprOXc8mzUwONeXte/JoUQcExwqP+SYwrzguOcAQ0PBuHrqB18l
YAFRC5Z7i892IIJSY+SCaxleiZGNg96Pb+vyn7PsilkHmJ0lJpOjaAMcxJQsnLFr
yzfbkfE8izzAbqqcKK5N7p5g3pzQhwdU+LtskQa3l5OmzKO5Lam5Y89OQv7b6Qi4
/0U99e9iwGePtLeHx6sLf8lCGoW9KKJfrrQ1fdnkbtJvHs1wIAGG7f4kYK3knQtn
ZTYf0bfMTRPQDVHwYoZrs/KlwLXlBidNYymZbLpVeY5rJwd0aew5sKHZYlwLl4vg
w6koilnmbRLUT6URmFOpgZ/jtu+Sv7ySkiy0EEKCYLw8gXUyKqtsaxHTctSxiJ3q
bnheLJO5MTpa66jBSZGlzT2jjb3Ae5icTmN3wKMdvAbir5Cza82E6nnRsLoIDTEr
HW2DbyzJwubmeXX7cOtoz2SZjknahtQCGacClXZf1J3B55doz2Hq1+E+DYxixQmC
JFHNFJcXQ9Jpr41U1u4xBkkFU/mOJRGtHfPV2SAFI1Hd7WNJoCUacgiNstf+BYrU
y+81YqFCqP+F3DU6jiC/BqAeauZCuufXsAB/dTbJKMiulnOFYOBvHb5yimqNsUbf
cZ4B62vZ4xF24GWx6KcGbkmUmILdVpuDiwDkihlXI7rF/kCKs5Ju9+8qr6bkqrGf
mNL7aGyM6HyqJCPWdPmHAyZe7vd9x9haAcvAE2KEDocD0m71wS+MBOqZTkOnjlAW
W1AcL+IkzW7gyhfvnNJ69/WNIrotq+vHP0jwaDkdKDTxfuLoBAOMD3U27SRxs/+I
HiF00zMCw9VnevNXRu5pL908hwE+1iWi1Wx5Hj/CC5v56tvcPydUISrV+EBRZG4F
oyr1bNnY0PY3jJU1O8bgm5awZOHETECwUeeDRyBQrT8chuDHS8pgr5ugtXtVwTc9
d5pxDCbeVyDYHYFV/wtjGcxyTQeACA/JHzG31CVWDfCo0DFOynf2aTUaSJtlHcbM
DUjq5huDly6aWOkvBwCOIXNAJlWisJSGS5g1A7fAjfClZdDrYxeCFN+3vZ3tLN16
Aqq+yHNpOHem/1mJ/+T/3EeKku7a5tB6N/8tYA4Fs3IuC6Xkf+YQiCbMbOnF4Jlv
de73xw0hAKdsuBFXAVXkQZ92wmwtgotZDzbFgr4WWGfabLVUZYxvNiMGpts/hxgD
/fHo1otCSfsRqR+JEsLCIPEpBhbhNjZVUuNxfCHJwK0noafNVFSEgrQcyxIOQEdQ
JrohxbZKXBLtOAuhybyGP/pZP2iVz4P158RP+VgNbgscP6As2bXMB3WEXOXBaN6V
zX9Gl3/Rkbv5gaLzBzEqYL7NXh5wk+D6pfWramPlzz+1rb34v0vkhM1ZRcDYC7K6
gdw9seTec3FTsWEkvlirCUYRHyLe7ZUqZXZLg0AANpG7O2Tg2GL4wYRsIudJhh9L
jWb05bq3kpNo8BaKxnwikMniwKhJn2i0ZKYFd+PIzpVoeJAnL9O8J3zNpZY9mW0q
HOUaCFiALKpwOkXIJqnbkEA6enCicXxJhyw2VFSXkrNVxAuPf6rQXTC0E05jcp7E
JdqecsE1RAdDjsIjHaCakyTo4VzscJskRny4ou1oXHlrBmyLJswWCk2P8nQH9Fkl
lbi7vjKvzfLB0iq0RSVL1i6tKVOaDJUhtI1WU8Ia0TQWXXLb9yW8H0057WdBR9jb
/cwDgIg3b6qz7U//NXHo1EmJzY1ARNBEsNBZuZ7aRhdFW2+eXhyTu7DBlRZMmKyN
v2V3kDALMT2jNjZPwovua18gT5qT9P5VOdBbsUsEJNV4VwgYWDj/Oab10BATVPKL
6pWMJebESpBCOQY0bbOrK/xX06g0vo084Jm1GGd77vO5qVb9DlNkAYwVohSjifQB
rkrdtzYgBhvgCV9aVhPPtRvsibrzOUzFTJO+aNFu9xkyVtDyGNCT5QaOEmqGQsdf
HkswyatExBfyiEnOQTBrkveGPPMBthmHc5dhG2vPDBjH9xr6U6a7fNtNuUKBglMr
dCXUhtueJ8qcG/gRpzm20JwPj5uzk0s+hIby46Hfu8mX4Jladiak5xsXwQGyPXQb
7dvHQB18oMA9N3om5OqGvXSd5kQuyILXphZzUx8f9JqVm5754HNFi5xzckaEj/zP
BC/bFOODzy1rf4LEmjlWmteU3YunEcNF9fsjABFSauvNl3F2S3O7zVFMmIiC7MQg
LJFVpSU1DKxPSjnt0S5ivIKVtBIkZZuC8vdL2u2UqO7opQOYqYbJhc7j18oDfj4H
Mnt9ZBZNF5Mbsi3L2qrtjAovQaMG2Cu30okpSlg13edRqUjuGK2Y9icM6VslIJ0y
X4kc+fPyt2A1WnmjrcX9NlyESDCRRixnEdBl4f2jzWneOs+v2B6gI0qI56FQcYzz
1dkdZoa5nq+4MRDO5+YtTipPocUeqgmZlNDp3+Ca4hOrn3BP27lRXYyBuG2M2BGX
7ysSXV0ra6NM3fzV7QOq6spCHlcDjvul3Vd+mwKeltC0LEeDZ08UdXyYy1/UB8Ak
CF5+u1CBZMztpz6OVOeBVMhmfqUxO5mtPNs9Y4wvJdZdheVe8abe3FowmJCo0vTe
CT/t6CutIimoW3GJ4AWbBNp3AHeNSLxTN1v7Mp9/Y6nrTmcRsiyfiy0WlThKSjG9
aPm/u6PMsXyoeRNq+wlpNKQpVamVuOIyh4gyy4+p1hcwob73jr4XSOGfMTsUVrFa
AwLNnyzFxOtPjS94vHNBCq4uMYsDqS5CtMVneBg7XvK5jI5Br4V+eZdE6wgjtUUg
6Tk+iK6W2wghmKS5BC1b2ZfHYVd/oZtAa1hfdIlgl1kwI2Lwfdaga6E0f9YllPeb
JVoz72gcC9lp1LPSMcOdIpDjTxyUp/Ltk/GTITVTZ69Cik4ir4v1d0Ss7DAUly8i
8M0OrLGTtU7U1Dl0mng+wgTYdhIgjpdEw5D7wKp8sSBJxkMwRz/GfjCAjgyx30/E
DqK6Ahjwv/tMgRXTkWCIzAhe7PBV6ccMt76vQ5sCQ87pQFXt8EyVDjSiO8ww6eZu
oMTdlSvFU8etMw6wP8LyjO0UAEFzW4MZEs0u6oEguuODy+zXXxK0cqojXV0xPQW/
lXJ7HZoa8ytGfLDbFL3FD8EkUajVOAOJv4wvYlJSd/3uKSRhw+bAGDNG7DhMou34
/qxJw2cMhtv2625KlkhCo1njOII5YobufWFQplRcsWsLUDF7YOffs9Rfx8LmIdn5
jRxwrS7iJWqdaObq+O1xkrjgTA2yJtEIHPF3JnwRnO0cLXP4x5rHEQULrvTAYPHO
vSbuQbKYmDuLALtJ5sHa5l6TOc0/DVaKpdd5BnoqiGNuL35B41YqRyCXdeIamXUq
MO/2AnLa7KAVO4AhoSUvF/Z75UWCqjsyhI7EEQYLzT4cVnUk7QX5mjwDtgqdnRtc
zgcKmN3D4M68WRKPcFhpUX766vjPTYIAfYpKlk9Kq6lshfgUEF6UuBl5IvhaAEBj
m3qNnj975aclka2JydGn8oiZLrQry7WBZA4REp4xGjbsS5Na9pePNkqIZpL7jria
NJ7ahqpoQvnfFvPt7XrZjJXDsAU17+zc2G23Nt+feHuVp2xuX/tS/0O7MoH6APZ7
t6jkgUTxzPSYabBqac34H03ZE3TxJUh+CUBcsgnfYT3qmKLTBSRTnF7cvYuel/qp
7xM45QHOPEPhbNodv58UKOOsfcgO7m9RZKtoiYV/bJGfQ3a+Nz/LpqPjNzuSM2dq
25R40XXviZJgnqhXyAFxzB0G6cxSKpyzXnW0sxCWbq90iF29CUYw3DDXRxcZWoSB
c8PELAIjnbbwZ+7ZNELPPLRxVosqSoVCI/TxziqWoFnuuGcAxGCrTakB20xReaLs
rAXrQlvHZtWY2x1VSELRzPDRURVSEh2ykm51QcSCSZokypoDgT0O6FuiFlBx9QVG
W1IXVbvdeCMQDKqrzphkcjtSdt2jROeIySk8ACe31XpkG/F/PsASo+spmYrpj/L6
XteOyfLDg1dBVnOQzbzOT7iyw/KappxPKO0gfg63mCUtasgr+KP91G+gAGa/7Y61
YJBLLW1fFi/CkWRjV0J47Nm+mp7DqGumK/jXocNMLr/muklhLqqTIMGcBd8E1SBT
F0YTapy61eQDOBgv/ioeen/MbyCqdOXzIYctEUzt8xM/Szxh0duq9yeB3n7dfcfG
991oVx3uxY/iMJagbY5CCmYRho9IYh8jcz7jrzsWyOxdrHvwD6g+Inn4ABQquHLB
Yij6kvHNSW5aa7tgyh9lc8FvWFKW2ySgjyhtJNSzfLp6UmIsxcl4dr8D53ReGVWM
Xc4sEuNcTeYB8sVkoMBTR9FE3JAyoGovka1wsFfPnnvSb6zQI++mlkCn1P0wf3Cj
z2IRGeUoyYem7egdy3t4gu/FeCu+uDPy9zMMx9YzxiPILCEkOG2X4RLmqwBX8+/6
hDsVc9q5jnf9V75t7YU+uiqelyO9qmm87NuaRTpUic2AkeFPcS0HBJ+oWTWktduK
CZp/PEl4O04VdXvSmHEfDxEc3EkPFzrdBUfzq4EO9essTejYR3Mrx49zKN9YBMaR
5IL7FOVQtveAZGze/kmtK9dZawC0wza+g0co39WB/qQgCAQGXDx2XVl/9wX9OOw8
ADMBQj819Vwq41ZtPCH050Q/OJ/KPHJQit056Q0iNXXad/ffJrHRD+90q0W6lD+g
vXKW3LpO7AunvSCipH/2VhqbmjaJauFuywAZiyo7lG3uIX27N9O6QUpRbK5ncPxq
dpOX+g3luw+dn918eqo6LKn1HuqdtJ0oJZoz7cf+fRVQSUuxDjjokQurdaHN0Sne
JH4pjFXhHUZ2YZl8rKXmfC0dUwc5YJvPwWxTOG4U3cz7mfSUgidC3kXXrV8JPq8G
Q3PR5ORdnSJSR0S/10QsQz2GcQiKc9gcceyLz5WHV+73XcoZOPSiqsVDvhtAl5tU
qspVf3l+Bne7p3n2R/CrXc7D0dl62RiCLmB8gQO1ttXLMhf+RYlKq+GDsD1JDx4D
BotgFwCTTCiuEn/aq4O8TmfhEdXUXeb7WLEtd1QHgEveaZDgvJHDDNcFZ34qvpzu
y7H1uPQ6Shhy1aICGGYi4KbqGkTaCm81j1nlH7ggj+DVL3fSE6+hAvfn6nzhUn+F
kFuqg3Lj2nC1eSiVOzAUiFTkswQubM/SHUWLTFUP4RHqMN0L6TQPR46VXpsYdTjh
xFNLMb3KnE7e4HP5Qn1AG/NBJdP7Qjb4mLESs5YAFDhqaRPN2Ihb//uWdUey+8tc
4aiBQ2R/6MdpiSML0zeRpmVqV6/dPjdl/m5g0k0h0EiDDLPiJKYJhImkbwikR/06
s8DhHhZwa83yIDWlWIddUeBRT4LBmeo0iaVCyuFjPSSoXPLvxPBLH+Mdbp/mwMSd
SMCD167K5W8gFD6jFzFIUshBbo4gc7XyC7gvIQpqxde4SWUp/2x4IfW5MtZam8uB
NJ7ODU6U+b4qRNljOy14Y6SoF2swaYBgKtQO0JGIneDtD2fIu+NhRDYhK9200EpC
on0w1a/VZ02IXUQ2bM0GRzMpTA2ruIKgdMq7SCgegoRj8gUPM/q96gke4Qbofwdb
+mrB2lgXWGLvQTZ7GPjKVHCbn8DGKBxQsCD8eifTOo9OYWhUiMoXqRfWjDuhmAKp
9X6cCmODmZJpFBtzwH53R3ZtKttyCNevSoHvi4cYJdnlAgAWPjZJSvaLFmgfQLro
hUy+4a2hsFASEgQ0Lq3rjlWGByuz9SjwQsFlud6D04rDBlDfQ0aChUXbcQedUkeg
zu/ZVyFo/hakIKXewr2pwkf0CKlwp2GiiWdN0hr5q9SqFafR7VdyvgZGgtoSL/iU
hd0i67ml2w/nO4VBwYb5EvXAeo0rF6JglnywxZF4DQF6WS0B+WPMrkBZPWKElmAU
RF0gvKd4ckQfu+OPNg1dodGHAfeewmSbhphmehEiMKGYXa5DFHvUcuSD2ExQD6AV
OoS/+Hp4VhySUechVKvttAYj5E3sLWa8Lp5j4BCRv0mnAs82R+5oKRaElSo29gPF
dfgExAz5rB4qpD3QdgdzbQlXMWZnJ5DgWvO6lIgFbPTh2NRSXcaDgp4vWL9lcBkR
14WCx0D7c/rvO3E6OuC/CYfbql02J8q32lVHehB+ISsMj+6m0S/tRt/q5s5HAS2v
lPdm6sbCAN4bbZmHh/MCCXYlEXphQnXAM9wiW0ORmiMtw9qtRkKBl0YpoHyTzRHw
fsUDBILq8BDzn3gNmvbKxrrvio+Lyw5HsPHgY58ngl4awY8ExtbZXksSzUrdVrm9
5KhlY3FMlZisHVyNTn6cbLKQQpdpKkUYewqyQLsrdCrzziSgu/t8jBn6RUqZ3xaG
zKGKxJFPvwz5XDWvnLm4Ecro614y4K+NYiPb8xyl0R+2mc13qtzi/7/ohaqdwihc
+5wgd6MKFNM3oFToqesbE/klIySW7SiWlkfhZ89uBZ8kMTB5Xjb0SrU3de6+k9qR
fJqz3xLqbBZzFcKh0QCdCUmeGFjCp2WP8ev6Bx4uukzoU36UH1w28q1uZlAGT6zq
we75wkEoXqUOMf5j4Tavx3ebsWIMrSlixTK4p8/Ac0vBpyvpMqNJOtBhE6esa9Dz
cZ3IGFY/+zPBTZpLTS4wvbqWjAjATgdh2aXge7qPPll7UUTaAsOdLf2cpK502Gsr
TEEtTMvFlViAP7jUhkXXhaOeUvu+4WnB8aryEPCa4B9H5diynkAM229g9RF58xHO
By552e/yvTt9cYTjE8RCVJ2t6105rQkSA+F8pv5zqMHZ0ax5ohyiSjANmSc2p+P0
fEjYreoNCWST76Un/AnEie6Gx0Ld7Hspi7jy13GtW5IiJfn9L04lT+aleS7Tot8z
l3BpxPl3NVnP1V1q/1jl6hn4h6XmKVI4C4NB98Kdzc3tJ8bA27uvz3UnAvriErMT
OK8E6wftOWeRggChnj0xUk2OQWgn457Y6qwLtINT9NJSZ34bV6bPARPlXOcQnsXz
gqHspSif/HWrv4ZVVQZlYA614/ixazs3BrjM/u/MCgdOQniVWVCiohS5xdeOJxm2
wp5RQufVOPalt2wY+xh+ETHwATwILgZkSpdvbC+H0pboOuh+9h+HG+BPFJ/sSbMM
8SdkMF7fkejeWxDTEx0KKgzDO3POffPUmZyZKI8p+VX0cRKZFfqnyMLTVMBKEK9A
Tl28NRq6O8IVJhncK/M+AGQbuo9r3DVA+/busMVYPqHXlXyWkqEPK9xNkCUKEhdy
WR8UCm1+uJBOpErLDit4WEG5I7IN/Gy36ACu/QJ28kpeD67wkYS9MyC1IuclKrAF
nOS3d93pOMsher7iMcpJ/yBIzptPCtGfNxsON1SLTuIKs6Ltkf3iB/4O7SJJgKj4
/Dpi3G144pbuR/OSpbAqxmBpmVcNPyAot9KeDrmeorz9d94X9wQUy8u92xwvYHrS
eDaG+/d1y+Qu5PtPoo9gfaii3idptgCc5plZlp/nX2Ia/N97sUrEd+hlrFpD33po
i2HBc+gea6nWn+r1AagQZPUxyJ7uve//sxlH/25jNPJTtWYcJNwF+E2fT8xr4UtE
lFHC3qdlycePY0R3/RhNVMmpBhuI+spZCb4KzWi6VSzRIfjOc0abuI16v+Am82GT
YTU6t6F/J+v1mw5U2dDAK/ed9Mm0v9aaAMEZz758R43FxtHiobNrDYG7VWfLIatv
CZhYrSYfkrMwfRU1y12Km3cC+GVzv/oEXm/VnmcqxSv1iDAsHeCs9pQ3+AKoqEcO
8rg7EzS3sgCt5OXeQFgPg71zCk4RCKxRi+Ffy34Hh8xikZPP0QOY8nJucaO1b4a5
gCqmzOiD4I9FiZABugvHk/s1vB29bN0LecFImgUX9mGjH+JJgtJw30WgtSDqUR9H
n9Zt6w6H37c0MkQLeW7JVaKhK4DPAm2IT6uRjO0m0leAZOd/pbcWa0QtUTdEpolM
posJuLcRJQoQ28TS0LN8Kj6E3sribexc75R+67ywzD4ztYso2L4K83M4R/i7pnM7
0cYT6JsAiIpESZBTun65s1ZwH72yhx4lwzthcKuQ11gPLboXEFCwnWwk1TqwIJE8
fwE1ohcndgYCx7D1btgfySatGBtIp3EsktxGH/cZJA6cxkJML1c1vMWYyZIsWSXe
HlPhxn5NLT0SrDi5AfjAxJQBzTDLMFq78zT62KEaYYLxE6gMHtlj7pTGtpJ4eUAZ
eEhoeADNeIdh2kfIqCHlY1xfggUAbbT6EMJNnt2IljBh+bxBBv8cDNMUBkOPijMA
A2/xO8DYlyMTYloIr55QGi3rzpXWtJkX9bJy19woauoxyI8zy4a1YIQ+rkfQsOFx
GraGPd6MFQt/vCNaXnLe8IT02RIBX08gI9EZBTTQFNMCMm0/gFeGR2VT2u7Ps4u4
BAJeT3HXmfvVjUzr1wHfWVq1WgVrP3EUxHCKlUK6pNOArFBzwi3MoB6tI6xZSOvb
Mw48syvgMGCljP6ANdEZOBj4QO9p/0dZkEpMvFk1hpGED64Urp2926mAOANQRqNW
Zz4hXNzeYEVDhgy8nNK5qM9l1QPHo021QWZWv3JuZW4Z/kYE+mca10beUUvWQSbc
yfsLchjIMIwrsOa9NHT2598Ouri+tk1cgb9Mf7w3M+wkotK+1ODdu+kBPTk/aDov
nUsCSn+qcIzzKEdLX2NAhD3QevsCP8hlO9XueGRUs/9ogh9CxGuH2tQYK5yCW9cO
Olw5W8x95yQewmruAtCKNPDsRuv2mEgiuNkvJBbMmDPXm1xAbYPx//1SP6/WSLFz
df+LioZh6DH4onUoRlEEUZ1EWSJjAjPP9yDrANsRqUQfkXCa3knKXS5Pe5T8/kmn

//pragma protect end_data_block
//pragma protect digest_block
XvGRgg0iYjNoguOr7fBNVdxCgOQ=
//pragma protect end_digest_block
//pragma protect end_protected
