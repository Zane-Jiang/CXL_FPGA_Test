`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
FDvp3Z8pzX088uBLdlGkBCWyjg1lgwi3r2pSGYk3D7oGbrZb2YkiXyqcA3cM/XqI
+XuLRyS3U1FPZDhl/fa6cB4wjou1dnaniseMzo+N7CbO2X1Ybgy6hM9X4cnTORCI
/psX32ExSBbvJc6hRTLtPKi4wM/HSUj4FXw+2ApVWXs=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 44944), data_block
TpSbcw/33xbRvxfafmaRdL+3EQ1XJVEGeQI6hZu1DycQkfG4a0RMO8aJefL00fUB
SaO2WmVDheB+6xTodj4eS2QJq8FXTkMaf0PIsxDBtxr+xsrbOEudDpSbfrI5HqFs
oYu89jtpA7mmrWvz/D3IezO9sGTz+sHhhOkJLdcT7YTDBaLUI0htDDSivolNbE1h
4k55cFUTGkg121VnkzvAg9RqrXqntgURUwYLERswan34/VqTjv0Xlbtr0bQm+kcr
zv8xiWKufUd6NdleGGvnB7NQ31JDLM66qPe4xg2IEyAzuv0469Z5ThGQ3zES/CyJ
ud3WmjbV4jFx5owVAr4733y4pizQaSnlaPIvelXlot42fnzSXCpL79uDqj7Bx8o6
J7B3SRb3CqbEjHRA82VhIrCtjidtQcR8d6iBNX7ZEq7AOa+BIPNDqYP8yOvp8jmk
lZUzrrsgMUSc3/dQyxn8Jf/jfTQTqA2Cs/LxO8tM0lGV3ApOsoH2/5AX0nPQAWdq
pv/dj9kAMhzvGbQ8ZSEYgiO8QAGs9Z0A7M9xXHvt47xP/eWlf8Oflcu/GrBovflE
7wy/zyIanmW88nrjeHHeYykDuI9wX1cPFQOkMFUh1kcwD8RQ1pOXXttuBwI/iIfY
7Y3qgtpvuSOPR888vygcCUlaCCITZ5jBRwKk96vcD+fEBnRnv1KZNiuQ2O7uY2+K
zyyxrWYmROJndZTQEPXNl+qG0FdEe1DmlUrQDaew9lsAZ3fvg79Z/5ArcYdqAxyb
1uAP4A9BkJlkK6jZJ+m/5w08b4x3uT0QL7GukvhQxuarmoo5Ql0lm79F7chqbl/P
HiOFrXbfGHaF402HxM4ee/74DveRsL0/scpy6/JwVcczMtWSKJS2dqaGAJMqs2hC
rZuWH198AI4R5bhm6f5j40CgLlk6ecPBBnlQqbq8gjCT2JEDaR5Yw+wrjW3Vo7Oc
D3P4FRCbeS4UT112UontRmJCYEHPA3ie0hJ2C13pbBJAh80EkqYLXyVhbSj9qguD
67sh3sLUzcbP/4YESZiQE7wPVGxtxmZ+UZA+7oQT5YAFwzetVYV/ZFQjCA1ZIAVm
+3U6Ouw8RVF6UlPBA430rwEU6lXpIZyBJL1ntl4K4BHzJbd8CpaL36wcOT6EeMQh
mWB6x/MlS+m8QiBUMq8wJvGLTQS6C5q+Y8dqkuc/xygNKdc/a7whMcNxItp8oimu
C2BAcIAA7+Ad28o0gFIKlQZ0CwnK3vy17d2KsenGEVytGcX8LoG3cbWJ6alZ6ynq
vN/ZkykJ2NyiTK3Ipu/ayigfHeIXlonDSHl3wcMOgRVvq25ZUajWS1QRDjt8HHQ+
Gxz2CLDsG9kRfpf69cMnhEMGhaMsnX8n3ZqKYEQ64j3RNOOMYMGZYDXWVS8magi3
jC6NkpuiCJx32Yf6pTUdC1/SdinxnmoJUCK8mJxf5y7eR0GnwEW5mkXlI0XFDN5x
R3aQ9iZX2C56tizurwinnajrzV6sJI8b3cCIFUMbo9GFdK9Ovd4aRY+2THSkjKZJ
YxP0/iT4j6fcr4FhszkRw4mbXyquNSqZbGrGoJ2eohAoDh7C45+1hRUKzcrZoDbk
VJCy/aBOzSrnixjevwNcW8yQFdqW3YHzquPx5+wJopNRVQtXeKSxF/dEzKmrtWzW
OlqAWIWwf/y+dM0E0shnjAj2xnDtJ0mZmSBym4fE9CNgcsmIlF0DI0bUJRdlfCtz
O/wKmMaj8AlavYvNy/eJl5Mx9QKEk0Np3wI7l/w3YmVD8cX+txNX8Y+uOr1wa6mk
ZZ2Be5ZG7ZelaqC+JqqA9GHkuDH6AJBgW5qBhEGY3cr07eB1GuchwIvIiF6IenOP
h726C+dh7M8cef1JJpEZk9WiBYSmy/sZ/4ufZkhc7h/nCQ1/kbe/VfP68w5Mf6G5
xrYOAy7vUkqTkMMzKqOlAV4KLdM3oPff9IinEkRdzuLPU6k9eGctOpqemJtJuhQx
4eT9VSvZ9DaJqBBbhOE7/XUvBl8vbgAZa0FSbo368cEtRfiDTC+S/rcd2cFkyz/n
LKx7tOJQJTLCc9PsuEBxvfTA8L8x0MJ0naQAfcMgtX6JXQTSyJMiowUXX16BE10M
nygpEAFZaVorOHh3kdGmZEBOB5lQ330pIhek4jSSK6polp9XVcWm7vuAZgsmPqUI
ti1ll60a00+Fbq6ZYDUeDXLbaizId9sR7BQOUpykbmyzcOBC0LF7KHVRNIeo99D8
2T6o8N1TonDkKZY8aadPJbrjwL0P7xdVqfna85a5yrh7W1mmCeKrEt/ATRYMNEoK
RKxTh082J7tKQXx1f0wDvPLtw2oZuA9jj99bbW436y8QpJCByWs8VPfRc7T7zpkT
s6ChS6OX8Zxr44U7PyLwnWfx+arxK35ky+bRc6JHRwe1vF9w1ryNW8sg/4BcUHYe
C/1mhcBD0sQESOmgzwmGQPI4W0dnKdugV0KyUa+zLTN1rWWREHxujqkdyLxZbWOL
XKvuT/iidzA0oVstanPSBzbJvpkXrnSUs7TOz5AJikxRsXziV3bs6xYjSt3AoFBX
+3fu9HgwZSzDKhvR2HCM4P2+uWjrdEy/T8lpQHFr2CF+Kv5xtwMMQD7Nu+XS7+4X
PgNcC/p2L0rVUdBT1Yl1laZnYm848ycytFdqkp3Lm2W77/9Wo5tdbQx2hXYu8hZe
7Iz5tlZaGL3xo0o2RN/gajVAp4QYhCBKgIrkmPZr9QyFTNHObCXNdvuSvDuOO/TX
KHdm9Dg7MieYbvWbn6W8aR6MRqfAxuhOddBq/Nr4b6p/VzeTGpHdAekW8SkQu+EM
cCWI2rPIzH5uXCpL9MvBLs5yKf0DyUfbo65IBsOJ/egZ+gwvSCIJ4jlZBa1tOW6r
V7WU56AQ4+rT5rElb7i53+2lIge2DZJDenQ4rFUKLnHNcxNXYM+Ty3JLqyukp/SH
SQvAsXahqvSjAHkDVH4S5xd9iWxkLYeVKK5CILaVBIuquJfXK1an+E8xiLSEysXM
gnA7wFqRy3CbPJQYqIjgWq/AcTuyIQGT+HloNwdjJ8CziDAeHUdxqbgp5iaqqiXw
xaICp7pdroC40YT+fqeWa0o+n6Q4WcE5DQZuozIifEQg/eGdgMMkW8ZKYjjwvUJn
txpcDFJ3c8FHEhXLNQZzmjglYOZm8k43L5jOJArG00Ziux0k8Lu/fyG2Jzew1W6O
WSeMD98Uh7hZk4cQI5FFgzyYg9xfTE/4l8zuPU62paVYRqBGyzqn7rNqyG9tvTvj
nLRcsm2eMhTAUB5OLQgdUbCjLOuDVPaE5+APuodNwqd16vqMywxxrs5Eul10vuzW
kDLe3vhwsmtdlS9hGu3YkP+CS49hz1051MsPTT4AKyuiFAf3+dlANakBkfPLSAU9
uDgV5Qv0WzLzSaAJsWyzhPvh3SPQp6sOldnTJUxDCirwANbDB8v2vx2Lm19EnZVr
TKLC1S61CSH4MRJPwTmsh3t/fkfsPvyJ9f4Om9FsbJI4GGbhYiWJTzl5u6m7foH6
sNgTwOX1JDy1bB2oUvW8WdV7PUdR3/9fA1oPoKmJv1QMWKThXTI+fiOnOd/491+0
9ey7LOluTt3CSiLj+K5BXWU1nqjsQL1w38Ex0THmDmtxNJ72Pa+xkuUOLaUJWrWu
IHagRlc6sUNfnMmK6TJGH59R957LeDc9Uf8dd1wi36TaHk+jkVPtIduGkqhUsjvq
aCcTONbf5d6Xc0+u2Dc3DRywSVWDQLnbWB6nFLKac8fPnNP+fgYzT89hbBlA9u+N
5xe+pZM0OTPbHef3e/450hkff1/Ztt2LiFObajhVz40tL/PXAZeqAu5aNVs1MtRz
poqx/oeTSyeOQvWMg3s8s+yJwe60K59TFrNHINElpNMMT76U3jAvkg9wOoK/R9BE
Mtp9DW2W5s3x2LI4RbkLibWJO4RFmO5eS2bcBXPtXnDmcZ42PRy2NrzKqXTZo24r
migK3EsEdwI7W3+RBLJQM88FjRrcW6RSiAbxmnibmqFLUydMT1nLtJQO7HVRmrtD
eKDNd2/L/ayplbSJvT0Qvxxq4GUtHrF5+p+rQBj5POD3HFMHYkofKxlbu9nTeVff
6FPWqgGlPWjCtPm9v+1iXWdZTgpaPRWlgWUf8Gu+OvFxY46RynV9K/y/TywtlyMU
sCsNC8DkTph4En61sbqoWiyMYOODsQ7j99Z3pDJtOTMVFtZb761i18jzdrvFSQIt
siQMUgh9c1Q8derqIdlrUWJSlC9NEWIEcX2dg1RlWiyhnDmg+2NonADldQltgQL7
RiOiMqVJnkaBGeovTN5Ks77ZO5vaYzyKc4QlHTrRg9NJtQivJDkPNg+WEto7Wtb+
h7hgdOv/F0MDMmDb817OIEZGFEbwNyng2Be5z4B4L0ftqt56SB3WYPF+95/1DZYM
zPHU0YKZxuXL5lsV9EfYNxrGEtwF2Shl8egIkeDNxEzbrOhAJRDM8aQJ82VXtF5X
Jua61mfACJGXl4Y4LYSyekNIeZjwZv/ek7PlltPcjnfsqMPHyUlekYUSSH5bE/n+
AsIeURvy3uoBMDcmM/dWb7p75Fiigay8POQ7+/GZ7vYL4ESoRdV+8EgRstN+K8PD
GwT4q2Aoe2F74fSJHO3Q4ot4CUv1+O05Bv+oxdIfS4F4NE5/Db2awd09XpBHEbgS
dN47wCpbNcHpB5NPymIO8t0q1hVgwoa1OfMPKe9cc5j4t1+q8aTkxSOMDbIO+ekf
4Y9jAV/QM1S5wcAfZtWm1Rx6fckL/R09ZXWVMVnv0hh/m8OVoc1O78438uyo3vNh
dHAb450CX1CA/RVIq8faS0k8xeVljUa/WpQxYUUz9bB8FhzgVJHApV4HErFmjlbc
6brl2ffSvc8noezWpymCyUVNRMK8MZ1BXFhQTd9/6qUPmop+CqM8oCUIJJOzjxTy
hEMMiiUoFrPq6BxtLCPaZeDHGC/e/SIX2BHA+NDRvwbd0hi47u0LFXQGsaPGB2Th
Nwv0MZdR4AqB7gRobtNM48fNPNyCdWqJsUBuwP3fvGlzzVO4u4c/5LQgddl5Yfvk
bY/qFK4q7/m5TDEncn+g7jQalfQtObH9cpw+or1ShTb4G8/e+ngDfdj4UUjp3DaN
xINhqefoZ8ghNmc3CVVZGkcc+4tw2qYOyYaZufavnGmfE5lDEvi+lAKPwpzPI4V8
aJO8o9gT2nHff7sJueP5PL5MZjrAY5CZHzUXYpp8kJmlU4apMVJ9V8FG94gBiVnY
yqVI0hTvqPwFdQk30Wf1wYaBQSvIOySQS15VMn/65F5V8/upPyst8FVNSFrVc20J
XrDLTAKxxuXMFRQbnXdZIUpMvdqLbieJkHhxlp9gRhmtCDHMuq3t6i7mtMj/HFpm
NW1+SC2VKlLfbz0cPNmV3LfW/tO9JMHQdVA17OGhSDLIgsB1zkq5KMsWil7S8F8e
NZh20rf3VDGz29kDw4uG+n8/+6v14lh3KTiSbfzd51U1jRrFr5RP53s0hhXPNM05
ZUkpkrmB9gqT0eqP17cylyraivQ6Af8E5fZvU4LUiL6VlaQs/rnzaHTf0J5xmWVS
mI4lIxC5MRXMli78/MBh9cI7e+7faXJ+bPAnp82DpQ86dU6/VTYXD5w9FAZ91Yyn
7BBqJ41fNHLfF9WGDdEY5RF+UEpIFxgH5tiKfWAlHBoLBcfb8dsEhvWZi1rha/Oo
tRDVhyFa9J9ZEioeIk1w7Ayxxva7zv9cz+nSkyiqmOzeNeEkrkgdQV7X3Ff3mhJQ
0NtJZAGxGtDgt6LQCftgnxtck+Bc5iPR8ydAJZWgKT/VXv5/o9K2+P8lrtD24gjR
qwlOit1xE9UTgmsK4qjr97efjXnqsBS59OrnIMthPKIfParON4zsmoutyoVkxp2V
1m09OSYaBcfS4j8rwaKHX846Aztowlcd2I5Nk2jVqEjZqwz/0C+tciFL+xazUF5J
AKOHP/DodLd9kUYhgjrccutssJzmqddKjsa2UNCy+O+ufLhpuqf/efW+HjI2tYWu
wN/tRpAG7tvfgy+FB3Qk0qtdEcj6gJuF9JekHrc240mJF1JiCp+CCTIHNFuB0i2g
q66kWz+pAjmXKHi30SCbyeaPlcDfR8IVQjP0OOSCa0L3AmqB1b8hpoDndOCeKWmS
ekORqpUcJBzc0lQn8ZHZvnD4K7X4ZweE0Et1rakqHzFvlxidb8zoaoPuxzFiHwg+
xVjooV4L6iWUSI7KC1/fBxcCtP7Zcgyp3zmVmfrSWrxBPsOYkaN1cqB8Puq6lbxU
f0pvW234to2hLWdQnuAortAGiqX+rw86vdXhFxpjjfXiz84XbLPTui0VGBnEKHn0
YHJTiaLOrdwwaUFdtopDVf7BMh0ty30HGKb/4QGfDJNxj1EYl5TO1z0mg/8Qmjg5
qomPcw0tb931DeDDlirDRUi06DnCTR/tIg1JtG1HsB4eWRcM/7Vt7mJLYFOcrdhX
RKFaLOsg0Km+Qdeo4QqNVGXErBXJGK+qH8EX+kFGzKF7i8J57yQGIbCiJ+QcYcPe
V+vVsqeHMBVas9IA749zhfSCmzw1FMsmcUjH8fJwAywzos9yHCBommpMgHuRqNZV
QGAW8523nI6ObB0WmjYl20Y96qEiTqkNuorYwJ1YHskZmdpO/8ZFRSRwbjgTaqNc
K28QqXwHbFMpApafRuQgeaLpzvXWQ7c2Bq8uU7QcZ8DYRZj23flJYPFFBmWgkKKh
LqXBao2pcTTOfI6w1OQ7aQP98R7K5UfxEjqF/vzrwcykcYh8Tc8mizXbQ1yIhdaV
qlaKv3zadMk8sn8STI+Z3ZmhsJ6zjgxYTIVvdYYR/YomTRyvWxuOSCAEPlbt3ELG
TnPhwl6vXtSG7rIKLa8NSqkTaw2nhE9pkYJKErESgNNwZA1ocFR7lrPhQ41vSAhP
2v2UqgIJS0SE5nF7F3kWHfdXANWOFF8tr2Sw5cAtqCh1etorb+KFV8exn/uce1Zo
5piN3dw4/sIGZoW+xIu+8LQCuDUkAp/t2S5vIqqOARiKepBC+H4X/vI9oswA3VrI
7x1ewkRSMl7T9TuJ7BVBzV9XkF5FW3CgIAB/ys5ShgxAkE2ma91V5aX9IIw8y1SO
Lfc97oRnA9b8Qyt3yfv12b4e5U5n8TJ8dBXltX10gPQzshNp5PiXG9iVkUROI6yg
EhnJLWK2UvGAz8rRwwqAiH3si0kG9OTuHKAqASPLHqQXjeNWuUJBu0VBXgppagLA
9e/H2AXhl4uqVP+OHuizwIH2atxQfSBEMOSCO2ZblZjJz2H7U2i+FHychLH9bann
372U1/UuobWJ4RKCwyzZ3iWlF5N1sPJN4V4eiN4soV0eeWIyt2sVD1AA38YJBBys
CW/PrqW21CcLLO52oY5BgtSg93GDDRVkKUZjE9RRlW5GIM1mVoXKMWMRQKzSS87Z
zKf9YFIAhEcPEO7o6N3QtJIY9pj5YTOsmIro+ZBx4Uv33311a+HSkxNgGVVs0zrD
sy/E5NeuzMQc1KyKTKNww5uTkuA1Un+kdfOU1As+ykhsfDkUgQ6KSDcpwV83wPag
pl2Aqs6EMSaqERLavixtOYLnlVJMCwa/CS+89bjYdDJtWjOHgLeCd4wN/S3cXPIM
kcrrz/OZ7P6kzxGJA2reDRCRyyl/SLr0gQpAA2GHeiyJBw3SUhSrYzVdvld+IK/K
o1FcGEJgMFeLM8bIGea7yiKmR0EDvY6Tkkc8Y6RGHnJSjfnQGfq75GbO4thg0EgV
5X63y64FtnIKXh8fvzi5ybMdUDXQb1E5hY5427cTqmNKuo4btmRgllQ3oW52jkXL
ShmN39eStjDvYDwkJUJIU03Di44Wq5hnyU3TDgJFGu8bpTxJJpwi4NMxwaFfRaEr
JhrTlf+pzXYn/EN+TiGqNWMepAJv5oPCWbC6x9c6kFeqSC3vuetL3XxpzYfh+BPA
Shq6MB0+u6JdSbAbfVytl6ycYqtjHlrB4te6IWTAsrh7zA4wVphsuyZRMquY0aQV
qsP5tp20FXg/xoxqiBQAXsn23OwEhr/iXV1BjqfVcxjz9kvjJmUZxqQTSgR/O/Ta
m80XkHod0p+LC2QQNxe/xSgGg8tr5kBmJffnAJ2P1239EeKKtOA8wSmL2Ux7PAC3
zzpNMBIOoPTCOxKTCUU1s99cjbGZmGpRcjcxjkK6NUMNjnfQp2BpExtSdkyjlnb2
z0dNnF3GcnCU/LvM91vhHqus+P10GE+Fih4PvfKxw710EL4VG5inu0asxZ9KbY8c
WodMlxkjJDNtsp0de2nZXr7nfiaqoEzXGudfUVxYqrUqaHJWNVbLV6N7ZUYI3GaW
uLnSki37qYWGRJ59Yvh+aIvkOlPKM3ZHtDJlB8Mj65pxHXcDr1w13m/Zd6H1xfxi
GnJAgI+ZbUcNFPPJbsxH623Jew/115F3H8aGIxJoc61RNQcvO5M4SmcVwy3ulAVj
/hWp+TCJ+m0ClXnBeBiPEnbbjWFKY/BuQ6EdxC6Kw5pKVLjrb3Y1pa9YM7abxjPF
g8mux8YoLVHd7PRx/lvlrzWB4EYaFX2Y64kbUE9J0OG/eZijGdCm7rX4h6/ZIKU9
OQGCct7pNNlJixVA1b3fJyg1VLBLsIfhEEHdz30oGawvEppnS0SHZlSKbRu847CM
eMd7DvihQsIF/Ps316NzOb4qjXB1l2X80TWpa2sr7mbUk+CMYyabWrpINp4E8LW6
Rke7w3WtBlQd9hUtsLIF0Jpza1hbK3Ugt+VhjaF1nNLLohLKOOsx/txy5cHaAJkq
nIU6CMHDt8jDuhsGgycn2CJy+CY7ShgP0DgHqGdmM/BHy3GQBVNHjm0w6NrOqdL/
J+oT4zkeGnfMUxP0tqDPNR/QKSixsexTJNmEE4W8GVJo6SpHPypMFe8qFhLPMxlC
10U+qKXRwFYduSFR+e9W0dYvGsags3aHc8+I/FBZr2s29V1RKRJyzr6WBIOERgT5
Hx/65Zx5ufc88J3VGz0Avva/R3urRZJaWwl1tf63l3ayjbAZDnJYhqJrcwHPLm2W
0zln5IRR7ys2U0kdFM0JiYwRy/t47qIroYGUD5OaC92+q2piFiTM5XI4BPyf9LFf
Fr7R7qNopj8DTUnhdNenlCjPX8QaZRzw82w9M7v7UTR/tw3IsWJ64mHr7V4K7ijV
yRofoC9B/TyzP4+i236x2IcI2WpKVw2XWnIIPxiXuL/gNpQMh/BAqP2qCxew70Fb
mWNuOmukLA2fHzexKgGj+3w5c72wZKIo7M/wTsVweCuA1praLEY3GIff3o00FkoN
rQt46y7tUIf6n/DxOR4tUhZepsPDQXEULyeEQ6wSmZ8SNWijKSfWxXi6uXlzNerg
hI7E7Z0oIadZkpeAz+DsTNKSJ2HfMGDwXo1LrI1t8iyTaZfH12J+si1kZjt9eN6I
HIEDZSdCpvsQkc88lkxPcxrxgfMTXPzsBen5tJamcokdWISXWKsGW4CnyfUnwVrx
HaNKt928tGwx63DVZQmstjxf2UwBE/KZ0dJrUscQHPd9vjNb9Id15oUf0t3T4TWX
A/bAZgEX00ti8jh0QYv0JX30skGXjHUEKGIE3JZPKZ2dCnqy70QY9g1p+Po/KwVK
TkS5WTQR1MWMS6oX/tJDj0XH0Ae7tevw6k3SxXuJ78OqfT467ils4GxmtCbGuRI8
pfiLuPtuZBtZ8R5+1ht4o3xmPCWfCRbMUVvKoOatGfNIe0jUYPi2w88t3kj+r5bu
Qv5sWrhF9sRmsnDkbmqCosu76iYmtuJ0zYYny46qVs9zc2OYicgjkydO0+quMYcB
bXZgBjhjuMjqqcUb8N1paVxd6CksYUEp8OnjmsA9xkXcz+RxV3JVW8+fFrhx1R8k
jGYYCR4HsPU5eHtkJKQI36u6v1Xk3jhrwudPVcsLWCVrgfUuolKJS45HoHL0t38h
yxbL6BDjYIjffGya3aWbvZu5nEmkdIl4ayezsZyuO3AsPwW5DcBUttDdvwCDYdNy
NWdCoAcGBmQ9jxnsfPbfyTbRMM6USwi8DG/YoAoWTpXyMzSNfPz13AbotSAplz9m
DhODk27u9rcMlGDy58xlnknoLLUGgIxlASOCfFB+wsd4xUJH9++En1M0PckuKKbw
gwWaZBD9R8emUznuvMMTKxTY8Q+drFnAC2SpJmWXro9mqJ+CZrds2O73Bur2tGva
FHgYN1kX8d+2xOFHBTN/v4xGC28FZtFzoBbYTgniR/qPa01sd80JyfyayQPJb2+I
szXVZCEqpQRiIsu3I7limLUQFDWgwCNldz2nWogoyb1W9iv6lsyf19g4iitGansw
RoZ862LdmCsggh/wFaMzKTru3DVEJDoArSkDEOEo8u5U7nFIIwqfB2gmxTq+qxvq
so6TacpOkYS5HEItv31mgoeehUA/6Z904rVmSpHxc6JfvYL4kpcwQuknbWaoEa+R
9uQWIC27Zk2YDgYlAasC5s+EWSsg7W5TZpGh5Pfa9KslR+inFqB/Oc9qsZdM6fk4
lk9l2b1maSO2FbXqKAmSZ7a579fEPoctVt8iM24xe5Scu+lKlPPoVC/F7j/mmgES
Cz/ubBNy3YBAbuapldrqy0j4TMV9sIEw/5zzL29vIoqeeYKFXVoET5TB05FhzHbH
b27Zj1ntsLgxeyYF/yaQ9in3cDxBZd79+leD+X4yF7GJbcRYYOZlY+ET/koGce+U
LDYHVoOe18LjfuolKvtpO8WLjUfrTEZV6pZcn5h3R0AzbgpiIO3b/b8da6KWg+Sc
gf0TQg4024Vs1/PyzjjIISw7Vmavr0R2piq06vOMC/NLF0UCVPnCItSKQRN7AfaB
RiEGqZ9BQOFJr5xG5esjVALS+WUGJaKIhX9wyG00AuyHkZvAiJSQOj8yOXncQ16F
T24tvVu+rOqnIYtSEF98Fj/0Xw1Aj+fwB8aTSpZrjGYcvurCpQZhHXc19OR+sh4X
83Z5yqBRj2jK24Jnu9TXBJhTD67/Du270pUUFXfz2JoYl5/gpOyM0QgMsJnutpnk
6rP3qnnuL5Ge5tbNAMeHAv7kdv0eP/pMoTcLxI4oSOHk6blnlC005PXX0cBqw3BP
D9uketxxkOPWSUiZdjVjAAUcKW42/EzwVVvfsUNs94r9Hio9yPX4JujSseU4kITP
u2P1gqkIWaweNSH6HIWzMBmNDQmpsEIyEqjUykyM+yBhKo8caQZ4QUOGLsCifmpI
dT3h1O0hXdIW9eWVcaxdqD0gRTgu4yYMqj6n3uWMOyltVXam3z3ScoNqxmkf94Km
i477/oFbEHmpckPZLDeQ3B765IZ3iJiqnVf+pu0GUJXoSOQgjksodMOZnMXLBSDk
wkucwSs5lkwXcNhGKo90NRpIkCeDuMBQJ1mpkNppT5Qa8JmLoDAavepVCaTIfbG+
Y5hC+jE/fVQWaCs2U56H9w3R24eP1oxz5OJjbGEHzzuVUQyBGy9TZjkRb7gcdP14
gSYY5/niDJKHgMY9J6bSOsDo+IT7mZig7QywfSua7POovqjA4sUgcoqsnvAl7lQv
GeEAKoZ0ifi9X2mI5UEZjvc1PSkYtEpsPkWLZhqLB0YjZPXz7SYbqfhpOtuKzMPf
7LvU+aaKtTCucgg3bJ/Owsbom9JqrxoTGbkpJfjtLljp1FOU1aF37BpxVq/zZNUw
7APKZFzP59+5wvGqgxQK0t1RVfQOv/TjwB6Up6Y9fOrqmR2CxxfXAg9wH0TlkgC2
iS5qSFHJtJbjmCDaivJOyb0rLGa2qou/E7HFSogaLua71wtiGlJxZJM280xaiH7Y
x393h/bDHW8GYFmFcgJ5pMnSZk3h+iqbEVUnuJcfC24vwM2smg86/wonxB/RFsHm
7cgLZhRP4EChSBwIFhS/S9P6/piCD0sh8p68J6UgY0XugSLyAPkTjGyA1ZQi+4J3
yFUQpMOHl4/sxn7gATb3JgzrQcGFwuUvA9LHx0H6CEGTY6/SOFPa8+9OQWVuNvkX
GarwsUrouBY1Og5WqiUt5CEnJCsTIKfK8D7Ij0vGWbspXTxPNOrTsrnTNCY5925u
flRk9z4yB9eiJ/2bUCfwiCqea7QiAguRxTXT3j1idum8U0YSqVBggZXgo8e3Y+Sa
KOg4yyaAW2azKk6mu60TrVnokJF7n7zdXDVvfHXmd+JWplBluPdMPXh89ZxqvR6+
nV7nrqRHNj5LA1URNtnP8NmextaYj/edFbNm3+2NstfG7jV2hb3IjWY5gGcZUq3b
3GfXgToTA+JnFatbjTaL1XQkFZByGSq5CUCpoICzTed/y0pKAvO+xQZq7Ydm8Ra9
evHi17/DF66Yuhue/9dBYWbHkuBYT+YLQdBLTUhr+SQfktN19QO4KhArvU+q6eXr
Me0wEla6pJswJ6zK/pmVkWsYuB/f7zWrO5tvbdFxqT/I/jnInidvfQucakdOso2A
42tCEe4ve1TClxuI2vFMRthzfy/fkPAm7krsoF0UtdJNisGk8Pfom37M09dz/Za6
FGX3bSOzD+OTfISWi5V9HtJVlN6VxCe7lltP3754twChQ+1N5EeBGVhWZCcyQN7Z
wJO8eJeMU1SI3AFYUwU4QHTXxhuzhOSYEtPlWEV6S9n+aT5zqDYrmQ/7TvWl8O3E
2ejQIjrg5Bm0lQCev3oeUBSXm9JSQTKE6nqt6F4+iU7h9GzKCKZySpkGTeJ0Mpja
prDMBsK5GKurREo8eBO3kJFtqosMf05dH9GUh+PruWtOVLaKirg8Od/LStw30KSI
VpWiWYvJpbto71URniNRqdKiHB55G5yYssWm3fZ+gG6qvPL8b/Eo+x+do1yzLulI
OE/oMbVV+7VmTVPoL0hFtZhCqC091AnTGkgjfwCnFeUgfaqS0Wr6ZciQxjPsAHuQ
kxLp1utlpkhNENY6wxC5fzDFyOchnfplx4TRmmpNV7PoCCFB83fi+0M83nJrSqeP
X/x0JRlR0sD+V/k+wL81heku6x8l82mJGXzzdcDt4KbuF/1iEIP4UAnTUKUOzCFV
1hprWTCzBq2WVLLgHISfeX89QrQ8OanymZb7Rvj2bFHIvd40N8/OJ74eJ7jYrah4
hZXWegVhCKNfuYjqO80wzFyrIillREqK3nXXx+tUYu6MHOaDbkT8kkCY2yCeKPFa
TC29y1GlDpF4H2VbyEIJ4es7jhlb4FrFx3muWEVpIXX3RHKDUYWR14P2WR6l22aj
gYmABDOiK+tnkehIscVqc7nicqgB8O1jsxWeAuWgWvXq7ZH4ofTPSNbpchV1lYXz
N1XcNa3+9brv8Js/QrpWEtgDqWGdRkDb8LIDWu4s2sz3xPxFOVCqd9Rdqccrk2+w
WvfSILWkqmm+UTQghi+bMDzK4jWzx+l8MhJv7Zvl2EZhLSM/EZNol2q5n29uXxb3
bmfjkjbtqaat9r/Fb6DA5hVD43n8HZj5+UJoE+/GDcC4ViWoaJZvFDgwEiryv1r5
FuYz/zKIQIJRAAP54LwxY9n6BM6rUfBx/2nJfKSlKR9h99ZMVTESueQyTqLIVhUh
MKseLSHwV+cNPqPNZUiFCeHq1f9C2W4fMWIqoLeYlTH6IG5NBkxAwtPFM7yyN7/C
Yj3iQ1VqwboR2DPuQLKmUBJRqJ01j60Tw++eA8G0IhbnUQU2iPDLEb3QRXwyOGNS
9axw2ar83rLSshT+3dS4yJy7vxgZvJwp51ckDO7mEwL4U4omtiNvJasCH4MXh3kA
W7OGBAEj5rmwaQnlUhnCr/5K/HAm8l+WefVXb9SXWYQvJIgUvwnLc4hI4hvjPHo4
hOEGttCgKkjsrf4JbH/2t+B1lavi5qGXviW9YLTsIg45BuaHObdQyD/dsBDpK3+b
+x4hiSzpKBf1TwJdSEV6Qf9Mqw0ZuMFiT3b0JrmnmxzdRkw57jTZhBZNY3+/8Uz3
05NTby+/IN3f2XG1th6ZhGW89dxF45HL9v3o1T9EFCP/zZaTlhNmJYqNMAFdDWYn
o3rWAU37S8bIDXlf6zdiAAtXJrbg6M9bfJsgH8ERaI6OvtlEWIVRkzdSI1WruIqN
JZKaLR5BzxALl/+MyzxG+YPrCgJY9EDRh5vSAwRCZCg1Yw/RNdQ/+FEbmhGDas8f
F6+J4FqftysrkgwD26eDwsIcS1NWdPbvlxzNdMdlJsqn3R9VnxDH1OTH2eewLZEq
wAgPOouBZfLoD2Eh9ZJHCqUqpXFWxt4rtOUfKZuj5Plw4sZwpqOlMGUi2LAJvGwS
5FvLJJicKDPYy5Ly7wo9GXqradV7/f8mPFgK/Vc4qgh0PFDsbRAOub8CQK6LVTuP
fsAp7KHBXfs5E/Q12IhIAPjkpbWO6obG8JKTgqD3Y5UDx9LvMcysW9FapuGCoU2n
MsHSeamKlUZiZ91WTk+BjO2KrQKRwoxEdWkMez1haiPWJCPqs7V4CV0bdAdp9wtR
M2Sm1QXGLOlLafAJ3czKCZM7WFZQt2RMB666DbWiCKgstioM/fWrQbda9iXVOhsp
pQQ4ID7JTFarPyCG1pocONOd+hJZkbQq5AAKF1+QHifTe7zbmgl3sLjmA7ywOhd7
nW4H8smewcAD1Fov5kDbwHv/qlvYUkiLTbcjbOngQEk0Vjur8cRRhrd+IAgggwV4
ee33f/bOGUZzUcIrJ8C6s8nks4S3aGs+eFQ8o/HBRFKE64JJ8tPLj56cUYhMoVBb
hHF9hOdfaRvmTLW8b8DHn7wU7sxnNUuQk+DwaLhCyndbb8b/FHcubDSVf+ITDOjC
Hz1rYIALDTC5eyczt5utm16dzJfRRWFI75fjZ0kcpuTU+lkQ30sTBG3YNFFaLOvL
3ght0pS+YLfi3pGxAeNiwnBHJGoE270CCcyxHn9n8vcqfJ+u48xLYBsPI2r3Ldix
oF1OmNcVVmCETFdxMuv/2ohUApXLRtJPgCgULGL4uXmmeJ28dwV/2dWJWFn0V8U5
FhR34C1VZltogITjbUsqCz8fRYc7FqmoTX88zZwiPi+yju4Zjq0xw2UklARc5Q9O
iMq+eyNJIYp8KxWWEqy6vokWpuw6jlVWt1HLsr0sphi7+P83blGB2YkAw9PpCo2D
Iv5ngNbdzp7ykYaRkaWy5hKms/788zBQmgzjgPmfg+jz6ukoX4LV0KcxrnskM+fG
01OJUyeRnkorujmtI0gEC1GFpvsqDxw1Rj5QrdNY4rMx2AzHCZTBfoSyYeSwsgD8
bUB5fj17H+S1VYU8B8d1qJBVBFNimZVByhkA5ULF6NZSwk7uwY20Nbak0ToeFLAF
XelPFMbs7XOqcmZm4jPOssDfqTfL4qkKbSlI/88uFKyVZGv+xy+2mQgxnDadalHl
6kNOu+HAHs72HOWS7YQmaEuDYbJd8ky9EFAcKycNiA1VSMd+kILcL8UCOLw3LH1L
LW9AVVYz2sIAFqovFdPep0JbcFbWdeSzjN/sjn7CxERT5f0f3yweiBbDudfqoxPw
oUMuMbIS+Fk03QczcFTU4SAonf2Qvtqn3JpYclhnQZV+BgTTWOqgI2TunfmeO8Hl
C1lCnljRzNqF4BERM/iKBPP9EztRlLbQU5iuwugP4E/k7QNI1wa+cm2c+CAJ6t2T
phM0TLavxgbIlBVbVh8czzf2DXKMrNVCd1KGHnNygARTFGBueQh+otzDBwmGTmmZ
l3f8hnkB8g+5kpFubCsI15wlZHjkHz22JDvJ3dKUZEfmx9EFJkj+6U2ZbyOBRsAD
D0puFL2f/p4CjiZfoB9uLdOqbb10dwwkn8njFiUJYgGueJVzuA25xEhMErJUOXcT
CkG6ju4PhEg4TI1TGgtjrJxkNvX5EBoKaZ3FbFjhJzy2jMaC/fSv2J4/tVVT/AtY
e3C+PhxJB3xntiK7Kn6U53bIbqOi/52p96Ze9c4dCcpiesYsJuuSeujlSgVwNGD9
tnf9TSKAZ8KCkO2Moz7ysdqNwoDpzTFTJc/xqfCkmJVGPPbnwFeD90gavoXABf50
V4ipIJKyLeM2FFylp3uW+lctZ6P8Db4qaXwXGry8BOMD5vn9OSKxu48TIcpU0zIR
J0mlB5ljplchC6P1+QC4Bff8fgIgu5VKbWs33ObKVnYYc6JA7N5Obk2wnioh/J+X
RIG54BCmYOrHP9iTHCUiAktHtWFi28tGyRZvqkAT7E2Dn0mUqamktUl1PSy/s5xY
a5eKEViW03cJfKS+ZjUCjI3rLg/7yQ5IajQQv/IEqGrgNL1Zb/QOyOiuqME+2/+Q
i+bj58Mt0YaXiRU9x+3/ZtYgCE6oBy5FhjaNU90jO+2Ny8A/JDC/cXYHv5XhPsKI
W+d0xZ2FifWFxxr61KThPxOI3O7RSGYG/wHPujatzvUm8xH55ZThuu9cvrKXRN+D
T6c6k4bQSUfJvqEpo3IJInfJh7HmP5dMoOijJQHndHCEpJoyPoVt+upKx1OBhkrb
gXnedOmE15NomAx/svHWOMrURTgT5UNzil++vCOBZrHFh7Y1QWUigVbXZYsbz10+
G7ZwZ4ta+E3gPIW1uOpu1eIt6r8ZrKH8ZE+PHmKKvrnyWg/aw0oeCZA6CnmjXN9U
cZLeHqCPJ/vDIjHA6w5xiPH4CfQdqmFYTw8bU/d73zcaF1Xc7n4jE9go3oC5xIY/
asty8GooX1jvBKn3n5jC95OWcOb4TyMVvI6HFvJ+ZAbvdfZOfrkEISr6I+0EjPda
bTuDdfGDjCeUds+hXx2dpMw7aL3vCvj5+0YPureiEB5vLG1TwkxNKmM1QkvjC9cg
Ztyp9G7njnbwNYUNEPtPqp3X5LQ8uhecTzLUeXfUJPaWvKOwLJ8naKlY4BIPgdvW
ayDjlac6vEsJ/OpabECCDzwYYHNzJeS2vnQM1ePRy01nxAm0pyAEKqugvuCxS9xN
pJnAN6wLsq1prDYUFAgfthm5j/cK1R7QPebRHCvdsKhAeBC+EQhMpvrhzKZTtR0c
Z2ognw6ODGKEYdJaZwyfuvDOihwYY72vRH9duAFsHUWtOWlGCY//syexlur8M0BD
MhEgmEaxDNHdBSP+wtYmSUyaoD4x5B73ZQgozqk5gEsl8Ydnm45hLikNKiGDynJ/
pQY1I1l6btCleuXOvDo5ybBTEmdBIV3czCbhiLMbdcRvs9KjYCqF2XgGNNJodngB
fDyKXoWMkcjxAssf6+Toc9OyHvmivVo5UFHkGdHNQzXLVny9dr+6rTWragpQF7Kh
s7I2StVvrp6lVH83NV0oxuHDGjCImR9gAtCMmvBLRZ9XrLK0cP0w4vlDiKat4Zxk
lceJwvHLp7QxLTawF89dup2pZyBm9hHX3/67slJh36Z2EL7JgAXLxgw3zNvb2cT8
EoIg/qRkJt0Sek/BRKrauXTHDgskrhHacryJkXA+QHGQMa3fi59WXee5lSV45047
pRHjnmbZNMiiHOtqIR0pRkaKzY0fqi0eqY8EtECBS15eWdlHz75JpMtof6QlN6e0
o6LsWqY9faSPQ2bUt80vhI4Ao0R+cKI5NLW/IOTXfprCl+DXjfBZYm9mZ5MgIeuh
FQOpUah+DbYM6Q3uwT6Nw1/Jv/xvH0binSgK4qWE7UhfjpOTTrHSFLxyMcPtTaxk
Q/nOtmCY+8YGl5mTIY5qdwwt+bsr4tSrwCTG1Oe+ksh5HgQ3+GlUqpf5KtX9H0qx
d0mKIQItb+/pMVxzILF/XcsgW78XCmx2XvJBt+mpvRh54JJgeI3n5Iq+bKe4BVZt
ZBf6XRFgRb/3pxybONci4HD4q8G3mL3yh7PPIQEna/MCR5CkLCOc7cbhLBpu3EqK
HWl3nPwOSjlW+yjTiAXmqJ3S5luuyZtf3QPqetmOxAjLa/j8R3bj1fIv7spFOaOU
clb+6gcez6E87cR1rW7kW2ZoY2Fj3aPYJtoAkyXVrBi+k+M4rdtSjbkK16UPxTiy
qElEEiOs3zq+bZaM0WnvVptr+KWFXie/Mi734dXbsC7lnobYnPqQl15WpzZXwWBg
9sQNiPVAaqKQ978E+U2+DThqsG/upZEqRbOuVJmYFAb7g7JM8hqulhU2kFpSqh0l
irXeJv+nrkpCW00Vpq9aMWDQi4BbeLqTXwQ1ksQ0DmqNQ3ti1J0KIl5kIvh3CBR3
YHhi7qXSjusnZ1oGgeB9UcZ0BNrbgQuq1E6SQTHp9wp3/FOoG1G4AdTnkzC881VZ
/3RbAcEMSF24rku1nh/nF4OtLNwle2eBFTJkdlv55Do38M3k2Syo5Fn5BO/TO6x4
EseB4xe34wMeXSYhtg/korle4lcvwUpIdUvrjZLTX8mGKJRLM/jADUF+TJlaw6np
PMGGmAThQs/MUOnSTJLMZNK8Fl+Aj1fh2aYAXLhowYGdqvGPYiY8se86sTafbpCY
ii66bdcd3588JwsREJTE+F1nR34UREcCuAwhBdGFsdnbZpCtOYVa0I71bPb5mE6i
brhx4L5ei/ppEsCV9C9BwUGxfLJ9vFTiUKnohzYJDmb8TRRcmk2WcN625qif6Oqr
9t1I48Vv42RPuyiwLwjhnJb8jcvmrJHLycH/ufCnY+/NyqNosRmiFMa14+L8dAgG
pPyMIoF9lX28pT9VVhwPHqljtO0eRScwCJjPiyJqbC+S1NwyOk8wdhnqICixJ6FQ
hQZ1k0halw8QGO6tCVVWsFatrvQyOonYuPJXgGmALfnFfDLz6GL3F1pdy8q5Edqc
qwfRRv4tRZyHToKn95ZJYBku0JC1AbaMuKhwZR8jQbM5SwZ0MIfi3+Nc/q8BcBlV
BSHwIxriG/eJNva9mfRVkPWEVRar+9Ww78NwzqLbbyDBNx6FPzHIOlxPlVbdRvV0
R7v2teWP3Kv6OGLU0cEwcU3g/flbku9iE1IYfgTrFRcEkptJpO2mXtC1A6H9GKpG
OuxxQviGGoALd0sz5RnRclMEaioaJUP0cDbwXKe5U/9qnBlW1vfqMjl6hi1MOx1a
HJeOtbrp2tTSWAL+u1+w0/24/kOHxdEidv2B/WsmWVbJBp1y7xz8KE7KmKkhJd/k
c0QEEeJtxbBFyw+HaRVKY9lkuEHWf6wT396VKwLXn+o3RV2n0NhxfkA5+a4E8Za0
KCCxNw7kyQv7n0ySScaO43rm1GW9OgSi3S6ojwGDgi9CKi6tBWITNG2A7L24zP0Z
+F2Gk+KbvCPUZr4EsL33U5f1wPksfD4E9y3jT4IEFnYYSeOtuLCIYOpUWbPpNEVT
LqMogytIb4v+h+lMJJeOZuUyUHJch1aSBopEuGJn6rU6d/mD/AzzjyGZ6InRzg8v
VsEFEecLGiql6QOyLOhO3lO0sfEQ/0Bpwn9ob4l2FDUanO1rFLw4NtG1qY9HZkfp
wX9No3avLeokVD2WlkmWA5+yXCSftKoe7KV18QJnqfMEKn+kvYe17galDaySr7GU
HhuvPqpBhmY6eGTn+B5bVjZmlj8C0LyydveYUBUNwNpmbh38b9uD0e2NX+iqVvUs
0kOxhfjsYozkcOnqncVdWJGWj05KD48IfQoHlB/I33AvyU2OvLFT3NzQ6sv06Yew
4eSVGGWWZKXOTvnodb9tdoD/b+NrPp3o1wRrCZImAA7/TbygHLTc2FH5kpKZ3VO3
vZXl92uLvZ3uKlt30qkoffcZRHDjW2LJDt2IYpa7OPwN0gvBk+vPJK2K2hSR6CdW
AhCB5qZIcJpmz1wl+F0/Wv0Y4vAJtj+K1LKH8rq5P7kx7Onx7TVdspSMsVh1goZm
odtaDHnq5H0zOhmo3kFjS49ooiDACT6Qfl7xAspjfYIg0WRDuguHFYryS3aeIU9d
FhnBfuMX3UIo3yMBJveAyrXQxN1yOBQtXN5BZ1S1An+eUIRm2YKwkjwZ9ESomgm1
Ka9QOF15Y8ymgUpA+iS0iIFEd2QE44hPAYA3lz4PXB+og67vDjPz0HWE8eARezv5
JtLfcqMo5nXf9dxA+5BDMoOcipGRsKl5zowzoDco+q8JYniEfffCHoN2npvoOMjp
RJjtRp6GGljU0S5wHmoZAM9ZWg0QMuFcItn6GKamMksrLlSXVDGWw7JIRTtvGPOt
i9Mk6z5nxNJy/344EGWf0Y6L1Mq9/QAsMq8BIL3Lm6ecImGlzv+Uq8hV6YqMIL5Z
ANZGblEfw9/T2rneFkPPbMRP02PSjE6MkDbk85qCbXb7/IFYf5CgUhMxm6CRvIA8
jN4pRH5QMx/jMJfBxzWgYmjS7dLq7p2XIuAB6fUfXzDNikafU7Mfdv5YuVP8g+Rb
GGC3pZqTzxAYg33Yy1GSM9ruobuhJlNsEjT3Su/TwuN0GDUPiNtkVNG5HidWqCTW
7/GiRjxFVdnCZOxpZxQl1fGn1FMeeKH1Jg6KTYewB7pTfAb2K4liw0AMPv9M6Xyt
DHuWL97a9V+5RwKSLEflbyL8H3r9ZSip+ZgkbzDc1XwuZZr/0JOqkL1Ns6wwXPuA
Qxm9E3FdHlOl2B8j4tfl+ggZ6URRcVqqBvQssUE7hMuvy0Jm+wzRFfeDQTKxCn7R
AwU6SgA1WNGu8MoKB1qsJQMxRznEeFIOCb8pJjalNuWJOHxl+RF9cUgmdIiqYLaz
ZWyglCoqmMFFHb7f0MzL5Wk4NrMklTKK9wQIXot/gahyECg0Mj6RZMdZeTlz44gl
Tv+jGp8V4njVsQ9ITI1nTzLZZ+PAlJCjdy5XDpuonoYGjlQ+YTpYn/+cvTBWvBMl
ITvzCq8iauVpFc2FsMFEmSOMxxQZUGCbn4J1TCRL5YbUqFYy3dhopxQ6vg8iot5X
gHLQ0z++5Cbyr0DoDVifQrf+zzs1BZmzamPPO9JQv3Wch/tM56B3XFOFWh895BzV
Cww43T/kt3LFrZSUox/Us8jh01yqmJeG8oOJSVxoWbuiInWLSUnUmdSjeRPgtnmf
FRcK+lesvaAsTTyX5Igls6u4Hkzad97f/0TUyUf8IDRgB9wegdZzPpDU2Z9iOn7l
505p/aq6GVLVNxIMq21KQ13XfJeebXV5CnqxUM7N3VFzlYwD3UJ8C2v1fQ5QTyRD
Pd5J/nqhbQgbdp6ZxJih2KC9s6vxY3E+jnX2l7+czFAi5Daan5uMVLSdJFbgEIbP
/AydmIst981eer7JEsp4W8T9mrHDuzRInTxs1iRJCvmSt7k/D/SNqFcmaaz5EP7z
pAwQQbZlgCflWlXZQ84Uv2YAEb4thMSq6eOd6zQTsZXUI/DW0nM/iciqGNdbAKjH
YJ4QXq4ecrWgyi5Fn9vz1rxXTMZvkrnnvYP2lqha05gkD8bzwSdt7k2Qd+d6Xqpj
/bWTpm3CMZ0JnZf9imPelsYV61EqdgaU6GHBQjKfb96j6K80JXO3CZxzZEhgA85D
zVEEeD07J15xWpeSWPtsiv4+8U75Umz0g1FzPp5BZmu0Q3sxIxD09VEpCSKjpE4G
aqkNJ0jPevCx6cEHw7WMa3XJ/EF19+LiL6gD4m66kJ47MyAZ1hP9dUmNBRNc5SR8
qYdcVbQZjNfkV8GTIEsfPN/Tw3K4dgHqBZy3bYm701boqnmZBnLHVlRnXPBGxH8y
j3gVJAq3ob0hT6ngoDhTGnjv7UXNiScl6+jbFH6fuCn98Mcq+5UEEaFN8n/BxJRR
NRL28PGgUYXgAzjy+3iTnvR1+YPQM/L3JsPfGeMSkREV4KsHA6Ch7GUIp6OinDbn
gbNtGkqQTPUtRyW7muuhDiohyvw5P+0Jqc0aXQkvRL+iOYfaAAlDZF/HcbeIFqnT
8Py1WQ6wjhDKM/PMaMIGb6EibgvyScKbmMbyIDtSF6Acnr/s7YnCfRQBQLylg09e
pI9TnU2Pr4YtXaYqi79Aq3c25wHsRudktdvBLZiEWlYnkruyE1Hjt5idNOKw6Kle
TCBL3HvHpoQurhjH9+w+VCbWrO6hpfFPyCKpg6KtJAenUmISkszyEVY1fdl9vAML
m2u70Up2gqpVDc5UE1cFdPkzlA/d6Zpat3btFHzPjP/nHSafZtQ4XGx9+X2wX7v6
WkJCya29P06MRFqsJ0M2SmmuQH4oUIuXO95IDQSLdlvz0J7oX5LDtIu3SHev2tAs
9+s8FJ4SEfqIsPfbioDCbS3ZHGqG9Koj0LthW8de6ooQIplzDoSoEhOA4HULvCE8
KN9HVFV+P3bF6duptW2G2z3ktrCsPn3KbZazoYujqY5P0f/mKwW5Kh/BEr6OwJR1
pNlAHRKOvrpDJvusRmdXNMVHQDcTGZkwNNnGrEDNxwigBCc7kvqhWPt38jkVY8Tr
Mb1C+6qnaQMpEA1JlqWEeZDUpHU6PCNG26vs3fjRjKRr34sc6YUeDEwrMTwn3IoH
7pVeMG1+FReePqtRV4sXoduFpK/QyBalut8VsoJdW9eDxJA5HwifpC+hXt7EIvTg
QqCEkXPqTIctCN/klUZsxwNoZjhoPIJDS9gxgcAXjieOhwKZ9lek8rl097mMr0gX
Nnx36k49z3veC8ZxXavwJK16f3BUgmN3VrzcGUI78J+g/p5nV39BoX8S7kmua+Fq
6pUC6yKfaN2MkvxYmLlOMZdAKC2eJnOOqtvoD1uQZNJP+goWjCqjplwPH82A65ra
nYNjtbyettEDetkE493fPRdYQ4GzKCpnZyIjRsRY13vgErVCP9bvlmgjopwiCJ6q
wIagvogvmZvWAUgRC3AoYwBcmUYLTi4ldCaqo7Z4qJH3gPcJmwem3XIrdn3G1+VN
Yi3QvlbvhrD5h60GS8L8kBU91aPxUjbIe+kjsInCuAl5I3hJyX2Cqr31PgQ+iNyQ
TvC9kyoAoNTD7qPJW6HiU5hPNJaeRB3T3PTbAAkwIau2YUovT3FvuctQSlfKZnz9
G0MjLzs+A0JcVqJxdpuk4zZiCllq9Pyoo2SZ1XCSd0emVDcoL0OouZ8hyAf0jlB3
RDwCBu+B4soIXdJUcrXNXjN8hCAhJydBziz/A264Dv0CTXTjHUHcpVzTLRkdZh47
943Znf3pjZx5LiPKX8xhpGZqfnBG/dKwzWYZ2myjsCBaXSUM+UsPAbZ35QVOICiX
JDiYydGkwCUPh0t1juvEOq82/NJQ7D4r8kNGpNmPqIcYprAxASx21IRBRwuoxk4H
Q4vlug7TaKAWYhRKUhhXOOQLalubHuNKV/aQg7WdPqBXXeX7oS3dwW3yQN+v/zfw
FVCKaH9QSmo8qFHk+jRtfjRej7OWMBlnEe2cXnBCg4nABPCnhde9x5aeDXu3WYtv
KLg2PNhDxn60q9QkBTWcGvP7SkZNfY2ALMH25TvYuPbdaY9HrlNSMq56fhsvIrWk
ogqm/48gMAdgzsFGtlxpqf4LIzeHSurCBDEkDAXsXI3wcG2WVRFZ6KqcEstETGXH
F7xA94qXOhbGD7W8dl9+NFWL4zLWWs2u2CBGIwCSS+EVLK5CNFraJIadKfRKQjiq
laUFnPo0pl2Eq5r/UNCaVAAi6vYfglzAKC8GsWKWACczXe1oIW4iM2VEIVZjgv7l
/Q9yqRssx9Wg8uRPdSCTfJLX+OICeJIPyVqBxsPlTjx8skta6GsZgjSOW6OkZ5z+
kuYlogjLx3sQNpFID0c9GUaj+mqME0d7J1Rg6PI1hdLnObYPnL4VXWRnEYnWXGR9
0ZQmnzhmgPbZJiFW9O2YB3A5nrVSRUxX09N6qAZCPMNUs7CjQ78lp1dYOq0aeZ5a
EsyjI1f9WBvc04JdQxH5PbBkVlAUXppBf2S4UPEbvI0vcq8/xqbMHgbxZNOuU5w8
KeX2T5eFxkXUhEH0gR65lPzXocdqqkNTUvwkNMj/D6WDMddoSGtzeaCHI0PCNtJl
4Nh8tewCjnlc2aROGK0GK8vydrPgjiaBaOL+Km/rRMd3eZNzkZHPFzqtufbzgXNH
g1E9dlqpuF9W3kXxWpXJUDpVY1ZJcUnxR6P7uYuz5srE/cdLarnHV0FXo2lJMn+7
5t49re92C+/emRfzL0N00KcM3g3EIn+5hqGyFCf3mxZkFdHWY67TlTRpGSSXLmfM
zxRM7AZ6gKZdvtgZgGYU5fvg6HuTz0ecOmu/AiT8AtJc81WQ48Qf4RCC3YEZvKTN
9vpv5C/Hl6/JYRoQAl/0OsNtOxPTt21AbQvACXjbf/z0YJt8Uj6SLRXpesEZPNST
RskgPdK7mDYcmVV6xAFnLlmB/BTHRQfNReYYfa+ydGAB4jEE/V2zTsFe0LlLuxcH
Vhh3/Xzh24gzJxe62T3pxi6WV+vgwoyiucRq7D3mRN+63dgDkCiGO9w4P5fYTv3I
NT4WD4UhiwElTBiNfv781ihaXd+ZW+ffta0B+N+bgrxW4LdrpV8DORXJ7CktXW3S
6jJi4c5JVIwrdHw8j8LNAXDGALKV93Jk+7y52XqHscUYsOvlwAQDMMjtZCIPZTZs
VV0VwGetvf6go23oKXwNElZ26/ZjRS6VbMBNTFKBo5gUR/lMjNZdZt3nz3+z+o1t
VFOCOSN3HHnPX1hHQMUr7F3gsXwplNddjxP7dX1HWEvE06HxooqbLWThn8/ssJYX
3Rj2CAnP0SBicPQWX2hVHjOjKZJz4aMiMKbtm4eFP4FjLFXilk7azvhcWW90rbV2
NSQohRCh4AbCrbeE7Ik5riPG7pNG/yohW8CGnhlB0k791EyYdujmG7pYU1pHwJo6
G8ghZ3DyO5VRCKRnCV8AcSrpYTzx+KoMIYsRzcY3GYvxmFXJ6UB8ZXUZeiIOAXY6
aJJhx3rR7EC8OPyaq2t3sIT/8LvIrlHlv1BM6o2NZBPMwK4VbfjtfhoulfjXE5bg
f5F1DYzvL1NjFcyySPQ1+I/qDzA836xtRps73LVFTwIcMlenH7tfmGX7cksRJHXS
WBl4wciMdChYrywK/sMjHum8V8BfM9iSLwCKPJDiJLRVhvT87LPpfrQyHLuUMORL
nGOPlzgV3v7AVAxVF6P1mP4tMAMANE3XDPM75H+S8cwVCIgdNlMnPd1ygwxds3Wr
8v3MQo/437mqi/WzSnF5sxmfIev6+rLnHP3n+7N0nyjr3OLTjvVq11F0he3qSmqM
8iIE7OeOX/9SxdDBHOlt24/FkvhKc2XFA2GgJWKkmcXuSqFvnEPm1GGUjk3g5zHJ
Rg5iKDr8m2HsHWa0npPhNk0oOsmtrKZtTyIXZORYJNFxdX+Zjkndx0aq3UOe84f7
9BOEHtc5YJ2KJzM8UlcKjfYt++jCtMrKeRWkbj/8Imdegbr8i/uGrTxtNz8i2OSo
sxjVtuNSx0Ou25tNBAPNsfL29fu5ux8SGw8f5b5F9wF0jo3lPmRn6/8CLp2dkTGd
jNIZcaZxlj+dXybLsMmiKldvUQff4nmVF3S+pNkQGAIJQuWr9j/PQiuKaXCpno0U
9vMF+0ee++nYFc/xFd8oayO6m7f41jCX8sGI5kwBArPM/FGM4JTsv8LDI7x8vK0V
UUS9O3ueXYcUk0C3R+phT4kWVv2ffIIy4rx0tBWvMihe8c9FTQ0ej3vXpfCU4rVm
UyS6xRYZpE1/2QxhUcy9gp17xPT8smub5HnGVvarHKdGXc5xZZqrZKLSeTWPuAo1
ShoFWQIZNFJiSu/yxJkO5A1iraIUJDUAONLjyyM9oYVRwpjBHciZskoFFiE9pqN3
pjZ9K3nmq7uQa0tp4Ow07lc18MWPWWZ27Z2fgXXPWub8bx8hOsBznksDIHWlJTmm
wsVN6To65v2A/LuoKWFHSMGFn4E4V9cqwERF9yoX47aKWyB4F7sY4yF15hZb+pd3
wyzqWfWkhPgB8WQVBd4ETrG0tiQ5IbpUQajkQ/+LnDnGExHtU1Hqw2+UjN8/nzzP
IcFeGgDDWJsUoYilBmCSwnDCJVzWPVfYK+99yZlDss1qp9D14Uaka8VTRIBlMPLd
kBFA29Hv0pV0yq2rUbY7zgns8UtJjQ92mrxx0PXt+aHt/MYDu23XglA2nuZ4hdTQ
9VpR3ySvfilwGV6JiwLPLo3xFJuEH4X4xvJ2HpeHjOnDSupKAjOrbfiTeuhEQ0po
fVcMoiDO8bzwC/ihA2Ufc50C4Jne14wGgTCnMX43iKOD0EE9Gtg0af3vxY4A0CFW
dnBnWkYIuKL+0EOBrFqqs3ERRYyIBiUcGARxvjwS7FPAZ+h+j5LFnlhvHJcf2hHP
WQqtlE0Lg5lAJae7viHgOXit3Kku8UuVABgP6ZeFrGnstFDu3thJiMF2kqHVuuIg
jSIuEowvglbChkZhDiQrhOBP4mXfWZxb1pwhFPXeDc5S6EbM8RJ6DXBobWf7zcCn
WsCNi/rX/AHZcrf048UTc6oeDvevUQAskcfZ1kpg4bcAgtnazGaLNICE701ByF8/
SOgwNGvMNMMbEWAlOq3Gum08ZbNlWAQX8ldblyQ2/spksSeKls/ybKvKmcHfXU/R
ojrznOA1/HXlO4v3kucL9mDwvKywvuQ/sawJBXue35NR7boFp5U1oEEn0f9k6l9V
CjslFFzZL/uJFq3rOd/FTNHbETPMTPe24sUfE8g/XxidSBtJtCmPsjPr9A9Xj3Ke
5hsq8o+XNyee0rTn2bIYe8GxITNsAIdENwTzC6MgtnuxT4lhBLv0SLyMhas+rWOX
32hDbsPswmi2jtrH2nYFV+gg4G1+SK0xSl7ic4Xi4oVu7MEIIFSySWdg9HIRLSto
0/0lZfHq++lc3l3lORGyzVmDOWj8zZsnOSW5BeDpYbtyeMmdoq4OfwqfFvSFis/3
4+iMWFbipd7xDODeesIgjNYP0Mq3HTH2j4sERjL/o022HBIbDns00NH7iT2uIIuw
Mwp4e7YsIp7wA/mFbDjUAqf58l9oEiEShY6G/cXUvl7fwAGlnvxEltU7vEhvlONp
0B16V4waolr4sxCWcux2PpHhsU6sjVUKEvaEuJ6EvFbZyGHXkDAon8XnjUyzy356
IswdoZIrFFehGa1fdn09zuPxJEO7HQ2qCXYGtju0QyqMq0c2MMwQiYrRMFqb0O3g
oEoPORfOl9gl4k4OQcdzdSdTgkgKlkk1pa2HxuYkwiU9THQFQ8/+b9DcQzLqqRD9
j5hvEfcdwKvo7WyPlJL8J0a/GDGVxoHj5pnYXiZdkH83NiRWcFWJ6JBxPWRToWXH
VYYhuRmvr2zqsZCGcWwgNo7XybF8wOS3Tzo8vvV7PgOXK0V/gN7TyZfNigmRnj1k
RKmrfJGsYfztKj0Pz5EaePTydScbdw8Dc2ek7KBG2uRRVWn6awyixu9jBi18YyHG
Eik5L0nli9CfZODvUVDgAKCzB/WG41ixG3y4HKbrITYoEw3nnGQuv2HDCY41Z3Y4
DOw17vv3Xnenz1rXEyYgmZoKKHYwekG5CBwPVy/D2i7SHBRyw7hU9Kuw2epE916/
ToKWthlwNdTd8/LGwzeJCLs82N1YBNEuOndkDX9Z+jpwE/s9DBuq9SGOgS93l9mg
wL7N/UVlHHykZOZoMoMm5i1lnz/IIZMhme56zpd8RyBE6Fu5ui5Lkws+l2NxzlNC
TaGdCWcfSduYBat+DGEaO22cYtnaFTMe49+qro14r448yftpLrt8haf/hcn+o7We
EAi38M5+NKyCAC00TFb/M7w49vhjSyo/aQgx8l5tcCvTDiN03iFMTdcMUcO30Iwg
jSyh3veaaFav9Mfqib0e2qkBn54dyZ6RfP4LBDEHBOwYX5W2NvQErA2X1Tm+FhBI
Ux6bMZY1x0a3O04ZH9dqQ8nhcHFr+hZQl3bt4Df47j/hZQh46Dnto8gl8tleG45k
VXVe3KlaEJs5QdSNz74IKYyQe0AyPsDXYALRZOzbgznvBOhF2qUWVgMUtepZSSOc
/b21T67BJrM+CklJ+Lu7vVfjSOmjYBmQPGbEeO782q57rgdMACcUoLWXy3vDZV9y
cKpxZeWPgngy36j9fuPej50HqIuvw4sCQvtDwFa4Obt2NNRJKyrGDHQ9lh691sPp
pdDFpmghcj00W3d48Gy0N5IF8i75HHNdt/PfhaIzBwqgDMVVIv/7DhJr7Tpw/MwC
zzClvccNQwR7rwFUWHgsHuZA8fs93ouPBJO6v6R8SjThspVJkLwKQjX2yoDIol4V
MITWEOEUd7X14i5DaiSiSTDIaRuhiNr4XOO8Lm0oE5BhzRof+sDTQPH+cWGrT0Iw
MMrHXGJERAAofoTDDpE8qVPTGtj0x1R+wkx0LlUsGCuf77Ief9L86ainZeFyTRgW
NySIANbGcRbIfY2hvOKj0KL5eroX++imOApPDgtjcfEdQnRibMHPjSVaKvIVwM4Q
Lv8DcQYXhHzp8tDoUVB5mMA2Jufn7xTW8nHcN9DBhdQglnEtzcVX92pwt+7hyxPf
isFHiFP7aAGU0qEFydW89Qhgty9Q6IrCwXTWLh1PFyvFnm0HhjeGT3qTFw+T85S8
rtCqGzwiUPe1WbSj+TAezTU490rLGD80nn+iEhn1lYFIrPd9FExBp/fzKE+XtQCw
P3/gaMnb6sWgrXvpJhs3PzwuvwyuG+t+ob/mqlSZQ8C7HoO5PvtuwM4JZpQ7x4r3
bE7qZOFK0M7kPtQjF8c/beOYkQh0abc1yKFu1mM9Klj9u0c8W73JQi55odDuu3/H
Njn1DiFWZcu3IDkb5y21EVM8HAkT3TJCcfSPFkPGkCfDQN2dow1HZ7BCUMzHDrd3
XV61v+/6sxLOWBoTrAeNpurB77ljq0jHgXae/zeOJQoMtIHtYFXZ88bRSxd6P/uJ
YHEDW3JapJ6bU9GAYfyKXWzppvmJXhF2kM3GsbgyLgGoN5NDDPuwXy3qiVQpu85a
6G24dGsDAp+oIauyE/ht2ZJ7Jix8SO/SbM+OUigP7EC9Qs96BE6+B6mExWg6EB2W
Kef10W57O7AySpXupeLBD5krTgIqjn6J0VaKtHFTKlpvhgq5LtLFKpXrvIzrVpXj
x+7CKUaSnT4rtfCwikZd0Uy1cu7m4GQy7G6/KktKByLdL11QAP0WLV7cjkPk1+1b
z2wXxDl1h6Tuo2FUyVmFBFCx+bs/YmXTahrGHtFlRAZiShkTke+Lh4Y3fJ3b1Dsr
GSBd5WTNYmeuLui1CiTno14kPo6+f9eioqYmM499/ySMurP6TF1N1Np0uR96Z3Qv
tlGD7wI1Jl+cFvyiA4GNM0Zv3Ojp1IWkgU4V/IoSFMqCzrhDwpgNcUV/3NM273h8
oG5FzRyn5MDsUpFYHzCAaogzzlQZYzMRLx5biMgZ5jHf6Sh/bHjlYM0ozqpR1Nyo
67e4SqZue/LsmcoynTUHSslvOFTYSpwIn4FH1gbFfaaaNmhozzBhvexaVM8L2ivr
jbhw0HDjiUCYmfDlkUqyS2oDP7DTGJRxTbuLLThdfMt5uZDtzV9TmOBlIbe4fEvP
WhQ/e96omMXc5pQyOdBzQd3L/89W4MCJ41uci3wfoIzrE7PkRRaLSrfHLk5DlXjC
FomobJVdGM5Vscmv8dEgfF/lU0VDOX6Oc3KTqODv6aY/F4TkKcvgHsZ4T1nRb1Eu
Y3YtvahmsU4g57VApG1TfsBrWPWqyq25DzrnUDDByJd2B7r/ljye7rEvtSmFbq70
S4E+8TRLuezvjrzgkmW6jnUuFPdGJFEdE3I0jxI++n8OvgdBswAGcpkacEVPYh8N
36LQou1f30oxOCFLLr8gDJBszzgDHis4zOeXAfIFkcSwshlOHDbAFwSv5TOIbJni
Em2tTOZdLJRj8UAs80YEPiQS5+RHr7gaWcZXkRU98YeeWweHofVf2Mcc4EXH92Gj
FwMmqAc0cCi4uA82FhrIX+/0RvLtb+IKqqBZLdwP+C5RnzqAa56CB0wqFZhMcPbu
MOsuY1jsOQ4MuBeJxNVGMtvtib5v5v+GlcI8ARDsnzwkPkjOeF066FSGSL/3Ut+F
QPqYVx1eqT898+I8a1V8tZc1uuP+ARFf19h09jRmntOKZwhPZ3TrkWkQUHFnGb6u
Z7gEQ488ItMGnboH11sxug7Kc08fI0KmeeAbp8ZoJYFI66zMw9/XwKvHW101Bnah
tiUmWL9wxlcr+DnFGHOvxiEhVs+DDW/kUYVF6mPi7MvVvVKuNtrzvCqoi5F0THXC
qIbFtfcNaBlxFjhg1PPZWre5JWbogUWWObnVXPp5Jb8JWdenx8iwdcaJhy1wiuBd
isSIflDNODk/Pzd5ez+4rax0mSDPACC+6w3t2fNIeBIIYELSBYftgKOOAL0kAZdE
nFWjN+WRhvuOuOSagTMjoq6PRAtYV6FIYQPXSFFZQxd3apYj8MN682fmk7pMWk4y
6GcwjHDvyZLmwROKsFVqRkDsfBikHxVp0MiWIsjk5APfAsLzWXJAYG0ru/cwNVLj
HAPtBq2t8GBAS86pDOQwrYtXR8UD78zoXTD26CfSiTzROHBz+QHoB+3gzrkrK8jt
V2F+joM5YbPfvjscwKBRk+sfBd+rOXFwz1kC6lwOubu85EzSXL7bkA68NzXp/kvZ
az6OmRItaSEvsZe5jiU90v3h+MYF3qaDwBsdY/dM17ajJgJ6Kn9IHZS/Zq8YWMXX
aRhs1Z1tPfAfYBsWQ9gc4NjO8QD434fcPBRSlHs5gqKIQeSDRST2xAwNQHxcTZLN
KCkmgjpt07/Ub6kCBMdv7HfjOn4J3Ghdc1xzxEGiEnCp/4TrZvuwIWLE95YVw7rr
vy8gffXv+7xHdVoBDYFG3nkP8BQT0E0QykvW6440jSDD/cEhVoy2EM+oKo6otL9K
lKZhyxANWbYOP95yjq2Wtl8coHJB66jaKzY1mGwFMhCQ5LhOdTF+xKd5qrDVjVGO
zkozggOxwPLZzjnsDmaIC+ElFAfo5/29loFGocbwVeZa+qXB2NSCfv02Q9Mk+Nwz
3KSAzwiBRxqBBNmanW1urdU9C6Vqq1SLl3bfMMRdwQa6P9S1CLu+SCOOXsm9zMg+
l63zOVKAcIekkz/CvfudAQ/xPHVzBwlEHMIIXnfTo3eaNs4LIqLK8OvqpQZIRaSu
qK6mmWuu+K+cCwMGvMP5sKEcMlrEMGPyLaRKP7LvMoDDCfiN2G4AJeYdRkJfkxa3
qU5JJgRE76mAT8G78N8hljlXfrA+5MTelOeS2x8XHdAYNy8HU8bkCRS9StF5KR7I
1VUjNG68d2rLSKBUv995WKkJNWkVaVLd60tCmvK26P2pKWGtunocwuCnsuGmAs0C
H48Cw1EOwkrZ7TzcY07X0OK34+/ParkkxSil+b6KkNBnjxIPpyA0zJZJhbrcnbjC
wDCJna0/hB4y1SrZxK6JS1SW0+yLMDFb2SO6g9fa5jAMWkdvcuKQDLAZ5U7pchHz
s5SS8M8w4UobWITiXUgQUtywc+HJiLNG75WF2sefHmxh5oR8lICkKgE1kU7vHBb/
n5+r68jLxwp57YopvzrdKQJOElY79CBSHy44pc5AmcSX7XLE7GKYWnDgKzv0FOEk
+BT0BlcSu58XZpyw3jw1XdXQmzfA3hX5CP7xmqj3aFsYz4jhCmFbcMTeM3YMGgXM
VT2zEu3yVmB4tbJA/KE8Sw47BybL13ypnpuQyn2+JdqsgknTUN98Udh2OFmnyeT6
2qCzgYYAsl+Dr/yHMcczpt+UxY7otjAjPEHUBcCiiAvj/JtfXFg3fh0xjfT+2j1I
2YoHIqZGMzCzj7TbPCpWRJkmmLHUrMRtwYty2BDhQkybTd2CYZ7mAnqvwLFpH5FV
/X2ymDLDGCZuxbJIYWqlmgAFb5HMX0eC20DZb0DrgOQHiSPf4z+pfdGlVjhvVuwE
RUAFQHq1upW2y7OKyhEWKLp8jEABLhHbELRM/SPzU9zL1SPASwzOvuoU6zIpLdjv
CUYkh0mgdFlYjpmkQsMHCOQTboLCLxUFIVwxEvUl73WsjE3qotAHBzf7ySPvNebN
otzK6zuBcYRyA+MHAhWSCIOM4OC/T8DMj8LDXMSzc7bPj9hGLgP1EiPFoKnNB6T+
ngZ6blF+otlF1fKUcfUgxAwhvnAA/uXwSBD4AeuBrwni+uxt6OAjMAEDkzzIp1wA
Gnf+xFnOQl5aQtXS1rrawRIhw6r5w9UsDdFQ0A6R7EzKIG/RwMaRnHpTaRcCUNh/
CHRks/or38hmF3tbW2okDZonue56pNTheC9hHqEFMVAkL806MPkyvkhr5Xn56qjx
eIl04H31rsEy7Lbgykb3BWV0W/dVqiyFb0TMnMTvxrT/tr74IR90U30EGagBiHpE
TPmQc6vbBOnrh0FPqexxdzFytm3+iJRsRnUJrbcsSC6WYeG17TGuFDdXfX4f3qyC
sGFRGCAlR1Y4sXQf85mjzr8yTovWUUb8NPtxIHjAvV7l3pUNbe4wHkeoABzhZhw4
YHp6Di4L87qkFRBiVbIbVi0iOQQT/ZxSKMYwPgk2+9UddtZQvW+lTbRyV2UG4A7C
4EKkvIddt+dwF5ZUBhLPlmiiclqxo7Ew2YRn1pHAkQyiidSQlfOAEEHMqbUp+TLj
cYNfYV9fImbF2yfgSHw42kgclCscCN32cWuRYA9J3Mc0ylPXXmL5zW7/mIzs6yl7
h1GsG2GUYhjDfQD0B2HiBt74XWj7xKDjmL6gV6nq6iV2NzrkXV3N+Dk9OoypeQ5R
yqEGU64qZxbS4Xz6/q403pyzZXkkBXom2QHhDWSCuWbBecyVUT8XZfj6QyhQ1/I7
WtGkNJNJRXKkTpk1kcIguRDo1SArdgXj8KcOBD6CNKYP0DDxxRoZisk6q1m1HIyA
23nJO+1KcLIdl/F76fqxxy3zX+hhhb9Fq1r73SvZZeWOZYl44RTjkKsfK0EFimjK
dlxDhKYimPiia9R3mQuRsBotNpTS3GrEluUkxoOp5H5ZbJeYYCeT6znsDryijAP3
C9irj7A66JN8UyGvKZ/bDXdEZ95GVZFXn9Y/a+cv20VnzS33AxZkPB6EzsEzBbyX
gJmO6589Ihu9LJOkicSru/h6D/BHPVYLz+SUZ3DOKzZIln2dhYwXwWdIjWuC0eVe
03sVCKSENa9J1TTBvpcnmDIltbIu2kRNsv799EQUYuaX/3icbnjCO1s86mtlAJcb
dVYuZA39T1y9FkYpdY6M/DgoYx5HVA6Baaa/Gx489ZMDnzZFzmlMCd1Zg3h2ZgDu
QaZuHqK3AkWbPqBNsnfatYI5k/1ocP7AWv2eEHpcszVfzV9QGe1Z+g9xQOIma01D
ltI5nWOM5EGahBk9cuvZFBb76nsU3HXGbftothZro+hCrCmTUKEkyQKgRuDtE16B
Vg1ahxzN/xlhjgrSYnBhIzvtZvWgO9m6ol+aLp84tGmmazkFtr1og5ZvVE0zyP/p
c8vyVq10d5xn/ylrc91BPzVI99/yMnVkPOfhKhPAoehGE3YwD79w0Qz7RSYLws8B
pg88yWyZi6u8kKUo7hWIj5gEoidTRE7H7m09ZAt3zRMsnry9V3L37Co1qgF62ClH
G0vwHGf3qzlYgha+3UVFt218U2CBLRo0t6wjtsH1HkIm3YRaXSflSkGTkAwrb0f+
4gvUsxn7kyzUrK7HbM1o00d98aYrpmamkbrFqSozwAAWuZEfKxpEbD64kjd6aiBt
PclC2TSr8+P0i/muRTy+pQI0jw8z3MPkaRGdLISfCfuP+HyC5JD6hNhYbvYRlPlv
NCuJNqc9w6t1xWAc/gI/wiEOsHCnZ1s1YXOwCikDrPRmdL52bmKbNNRay6Xxoyk2
pHWtqU0xkXt4CHcTiQTdHNU7GS031428jjx5hnmoRAaOpr1EVduUUVbKuGsjNOoJ
sHYcxI6XXwRvZMKEMfFtW//b9D333FjkEHsJOOYsITSpqd5q13BTRv32SOGtyvIK
iJi/vydGwuGqc5GLbXkOkMNrBrPZrL7yaOWP6a0GAr6s4NkVREt7cC1wLcgi3iHj
vs/QK8sUaElxcXRa1By/nPphX0Vt7fwoCRi+ux1rIQ3TTxBKtIIyX7DKn5+XvZHw
i9Q2Uw46LJf98OrO76l10PUSm+WihM8l/rFqXkBdeSlYz7WqeADFGw46v0N3yecA
0Z9qrpblflWiy8o7TN4V+bC5PfoUZ7fYmwCUs5A1D3pnE/6wPUG8i3VXFijzKxWN
d7BJNkijeJ4a9YnGtXvVVhqNTQ/fKOnKoYvh8GAfub2D3ZHp8qID5XX2JznACxsZ
E7UrdXXtP7rCXCX6VmnhB7C89WC7eBH4E4r3pP0IDOpe0sMddijNC5z0PEHnTzKc
Sr8R4nCZ8SgRj+R+hpxmRWL4NmwqZh7bokGMpqoNqkZDR7fh+7ZeZXHfz4t/KjJb
ykZwUK2fhfirqC/b+izuJhbNVh15AgFwOOJsikH5BGW/qnAdyA9XRlUey8I+gYIH
fCxpmP4tCID4a+y5WRbnJAI5h4/QCbU1XuXIsto5ykKSVT1nz5UOqE6l/7GDmJYs
Ai6ALeSHWa446VE0k7L7IAa4Im83YHoqxwOc2WdeR5pYC93phdu1CG7XigQBeZkW
jDkbPhhc3UvDWzSE/4xBQWe902FzbQfCEh3ydi7Ws0dgCEXMhS+tNGUeLk5PDEyG
2qmEGivFQ1cWK9/ASYDzBYs4ysrzxDHbkqBK2a3cYmx3URR2hRUXfeyN87JbryQ/
MlR8BLxZRGHAzRMRlhQatBNlQoWMiFaxuOXq78179ttwbJjLkUXCI4ayOZWGhH3R
R+lgj9d7Gi++3a6VTs/wRadS2hEj9z2zEPKSXI+xRKLLffyWGs31uNjhAaxmDqgv
3Wk55+Q1sF1rTj2b4wRfiwI49EDI5oWIdrZxvoq7uzlzskdNdybrWFBQOM9PVY4w
mBSqeQ23A++8BW7i6byrya37PeNM9nC1ejxq3rkLb1aZTPcNnBwq1KjsElX4OBTh
Elb4npq9MMAIOi20BQSjSKULFVS4XenkSi8A46rOK05WN8CYlcf6NvxojzXZR5nH
iAOMUFZGfhIg93Z3QvCalKz+JN5ynQXaLsYszwhlBAMsJMGapCZaYz3AK/ylu2aC
q84gsYei/KrwFVIgcNe9R861uovYyAY/G0S8hAWChmLOdbt6vpWn0NYtyuaz5yUt
Gi7FgpJqkfhrz0Zc5Gz4n8DTfxvycAhFQytCSIl+YOVi8MFsTaD1NGiHXU6GP8ix
9/vVzJGvPomDZ051UK9J+0PdaCrk1MKd1/rBPZX/CL82aKpB+yttq9j86iT667XG
dSyjsu+IbzQA1idC/mID3AKPK48F7X7ae2UQDANlrAWKGK4CfMhtf5p66m9TG9gr
J87wJszZDno6ZIqs9XMoB0hvcCpN54+8m4e94+4qUxzJ40Nm8lxcvK8KHVPm5qqG
lO8q5OSE5jDZhkoaCGVF0pT+E7RRScikcjqm4mgLnoL0HpVHA9W36yAXIuKeAhU8
ad3XHjqoxHHIjnBQxq70Nu0BVPYzEs/x6KJ0o0m9h9RoiCh01pQIBmW4CPen4B+l
Swbu5HGtRXk/7KxCdOSGuqKbFX0i3kWImMF8Vjw561vfYq8v4bRGmRvlGW0OWnE1
7z4gUQYM6bQL6xMM//P1RoxrvH20dJDZcpT2AnWz0k+dtJ3VkSxnBV+XaZObOi7h
5di4UTsNVXXpZpjIgehX7bX2oHF7l6owViEvm+If67buZS6CUEX7NC4Az7xXSbnw
1JiadEA6Z5KMgp+XaEQwb0h60FFJIN4RGx3xSyTHkaLdurx5iIo6cSbb3VF7Hm/k
+a0KKMiD29Q8yU6IZHK/f61+EzcT4FIfUUkTEEXFD+qRGovhniwG4cc6/sn0EQ2J
gALuBpzPwydIU+ns+uWl5dIpJ2Gzw7BAEb6MEDf4vGDXBqJ40eS85Fk9wM9paetc
PozLKDpZH1P37tndJ4wThmRSZpKu9XEbe7AZzTjqxAMzdMYWUpHL2yLqN3zSHX9A
HHrZV8ewT9LTp0YNU+7r7hE7necYjJCTJLX4bnQ1RrUlEMa9iIyTKWmkqFGrvI+q
/Dfa6VOmI54f8uSOjUolBlZm6o2B74jYjgOLcBE/GgPiat2y+u6DnXRtGTJIqFFW
rzr3od40r5xZDhsj76LkzAivEhDtt/cRH6U2fN1rhJEZY00Ju8X3fVdrOvbwbddU
halyVVOoo/UbKwo27pQNTjQ6UtjLDbDVGRqlaYT8ai84DZrrVZwOksu1CUOwlL2/
JHwe+uP7Duj7edmaTKgB5d16yfihNtisiss6nV8kqIh8h62B71RSxr9Vi0Lw/aKW
7WcEokvXdhg7TadPVyfL1t9EzXSy7Q1z7JtthY/aUCAOKGdrRpKxnSOuxvUOeVhS
Ekc4DTacuLsXlflpzYrBKmvGR93gvfeITWeTdpe+uQtRhPUMPIM3Q3sIy9x3mUUi
K63zi2Xt5FOO14zgy8gedn/IRNIamtj2mdCwWVBmLJFOX8jp/oItUoXQaHylSjll
xY5xzIacYi6ajJ3qNlGfqAEkhwGHxGI8m6Ai44Crd9CC2resK9LT+71Vo2A3dCxt
kGhdGDT1q4PhSZQJ350s1cOng8n8O7VtB4i2oIzRBC6ze553kueQiUPUZVxw7Yaq
aoBO3jdQaMV8Bc3KkcHQaygxm8CjVp/7Swn9CRm4UvlWzKI6Z0UXIicqVYcbgeuF
/BqpaAwoaV6uPphGtcshaiXrgbKxcGlGeLNFCeJUfVz+shpr1soepK0s4n7nmNuc
w81DmTKIUWFs5ZDT8WULkNb2aNVsF5u63KFVpXNXahV4GdSgbvt7tEhTErrCDLbh
4uN85pXuzEaOYXcNvOypoNqLbuA1F8DMv1zppytfzMWepFHVg3a5c1npY3X/5tZQ
zGLq8PopLoZ6J5Hj0FugXU7Zlh6yJjpR+MQ+H0b8mDCrQHZCCOuS+/UHPD0imndn
UxxWgMy/ReoiaxhygtPOyf3QN0Scj8F5XbTcNJSCWvG1Z0HEm/dwFT9Aqkg4JaxP
kz6lIbZYblkVlLU6vQbGJ0uzRUJ9ppJYSVN6tj7edxV1xpbwSHhM4xRdhYxfknEn
DluqdiRgfo6XhZm+MWAAVRl7zG46V9fLtGFYRKGLq9JCk4eyvJK5+kRCLnODFSak
Ds98RKrikMuy9Co0tErpaDTXK0zP88LdwQEWq59kK57cg/wmbeOLX1kPPpQMBprQ
cq0G56pg2AVIVZrV12LUd9U3s7IQU0igeY58iPxCht2PF55fqQN+gEOj1qa7agjM
8TLzVJQPZ+5AdinAF+/G6/kfQ0Kqn+uzcec77Uwym3RLdCQDiaJeqkWzB5WU8Ef+
1dUmYOeDYWfk7wPwpR6Bq1HJrSIcmGygDnSkaqqn7t98SC4uX5tv3kmR1vn3h2xF
drqUcYPToLHBSzvTiwLKMoQcaQyVeY1N/xE2ryWZhFIdThkZl9MYUQHVVL21EKeB
ayLpeuHeWt4ypVW2VlC5qRTJXez12Cx4HLrMPx/XVCkSv554mbFG4m/FFiKqbr1i
WHeLktPTNnaD5vxRCq34J+sRj7iU7MJuq9rYBlDejjuMZekAFwjMfmSBWtXZOR9C
w3AfBXUsrjTjy/x/rT/ZMNjEe4bibqqeXLednkGs5Nen9d6NdGfmjawTe/JkyaMA
jR+jnfmz1kDPtBjP6CEad5H+/a5uHxE+dFx5h8ZOUAujY/tWKodrPUgyuGH/Ompo
Mj0GJTPwAivSGIsagppaq687csVbZoSWlq9Yq/01NYvzu7bOqNJ6Rx+r5FX1veev
zz4RcOVmGHInm1YnlAmvEmoiDKNhlcN4jfbL/9ViiH1ENwJ8tGdX81i5rc7rYVsh
VXx4N0bNWLgKvcd+cdTcJuT8lvFwAdLCKUCB1NRmGJo7XmSto5ahNGSa2GtBXaMS
ywhBeXYjyNIBtk312zs+7F+4wdG1pHXX5RG+O48Ej1Nqejjtzw9SVYvRt5ZhpljK
MeRvabHziv0d1D/oJmg5vUho6O9gArp9GbfJ5QANtC/R8QfEcosXv3kU6WiCbHrH
E8TPSsZMjQUXGos4cHWGHN9f5HPQfD5MgpDaPBnzi2hmu1D6Px7hDBCSdlFVB4TQ
mA4+ixl1I7W6nSaNehyEAc7jKGH/W9N3BZ7GqSrDsehKg88sdHTpVD1EwqBAxZfp
Ee/pRvek2ShsNlpg/0maQU348ACV6OJWs4J9nI+BKIqcDXh12beLAcWpai/sRYPS
Wkg6EfjZe0gzPoeGzIfvkjrWt+lLucSp/aJK4C4mqhc7GSEBDCxYIHt6x6HC99OD
vZ57iCXklKExSJSnJ4zG6NSe42wLpseWyHMMZiAnAT/QgY+Pm3XzMFXj5mfuZB25
kkiggNks/mWkP+5WIIdhx8hZKjyXbjDaDN34AU1OD/rYnsp48/uwYy0ZlYSi6IOi
MuV1UHgqI/rDsnKzteCh6rk3P60nMWNibtpZ7t10QFS0aZIOnYpJDQXxM5A8FIJp
rfKu9zMnBYk1+75Rx6/pHzVLdwPEIxUdtppXC9TOLNLsGeJ00g/SGN1OmeGY9rFh
bXdIY2NgHrp5bS2TVjJsW7Clg9iZi0coUG+iqgATUZOuSFh/jBoKTjIeWraojlV4
JQRm4YQyyYNHA5XhglxT22BK9WCtxFqjqahIjNMEfd1HthLZ13NYJwP0lu4GcfX2
z9EeEhWxmXlq7vaKa53S9Yk3kDM6LatTvlfKzKMs3AVe5eMCk3D3qSQWiJiwKdqf
cKIVaR2TlWf3Qt51n20CT+GqXfiskLzFgm/Afb1SizBc6o+pQ0Xn9AgNXub1Gso3
ezntHTTgc9GjIZuJyoD2moKxB/7ct7Fek3b6v2fN5ljlhGjZYCJuimLKzYYLJIiX
cf1RjS4Fv+7uD4KH/mvR0KB2UlvMV3hq8gV0X2jFLRkk763k/pErIUVU1fMcC9NT
Qtag6qd4hvizVcY+yRs7NG/7fbX5rGWBoMkDxxJ4awO92QfhYY5yKjDeb+waFWt8
9s+1PxnPkRKx/zYX5UllnoY4WQYenf0HgS6MjMlJzAHrzjvBisGNf5MNMR4jZXtM
/k4QbTgWgoLOj2/wGKMVYzjuTkTWaIZmQu90U9GbYb7o6Frz5B/P4UpMkTwPdtQE
alHTIxK0enmrVDYEnLGaosPmKL0FwPdRWoVJyyU+H2KHn/zE/jl5afmXjJR8PyUC
JjaFRCOcTIJ2Fnx8vL5duje3yzv8PDInUlnPxaIJnj0SRUzr19XIbqGCB08nD+mj
lS+CT7h/1J1Hfavplo5QjV+8ZaYeWRkuEwrnJ0FxAPSOTaAjoGLkYupLru613+lo
PCTPvtkfueyHBqy/aIGpwN6jy+J6/sVdz7TkWGfc32VHrYV1a4kn5+APhUorj8LX
IrIt7yO4zrYUBzcHOZ7AEtKpuCgiNWUhoG9Pi5NDIPzFsmCtB7h8UEy5h/Y7FK9p
pCnQ6U/AJotC08XgHq4+4KPDejzLwCePSW/3NBmj8yjG1rrp8u+eo8RF7y6nw3Fw
i0f+TH60ivBv/bMCOD/i+Yquz1uP8I2b/JWXhQyEASwZbfkDkwwXDTs6tbOc0OOI
RzKhDVFU/r+jsYqa0C9AEiWZBeu54xP7PUQXBjW6dGEb6xYfdw359Uv3cPixjjNs
YH60GJcdeMBS4xD3ta9kNHllz45W8r2qkO51hP5E4FqDMwexqeq74oSxQmAF1LcL
DDAte+KTXN8Q56JZBq66mDJyCf7RIu1gx1uUfGcHx1Es4+6iqD/IZDil7nMd4L5C
rLeJ3LMfoEUpMvn5GS/u1JffiKgdzsrSNOr3sZbBXrWiUI+tKDCcLz0j0chIG07P
Q7nNbL+yyJ+t1yCGImM6z0d8c7vPs3Lcskn0z2vfOWpJ012Ji1nxZgxEBvSJLmlo
mhtHoAl98ZKqTT5aU9rV7fR/ntemRHvSMYXPuFj1Q6Tk/tPAY8akq8fknpX3V/8w
frn1BOYGDJDiJW6c/Lo9VjZiJ8+eEzMMtkAFWUgCcfLFyjGYTgSJ30lffHmURYhD
BPd6DpkKw0aZ/IyUTHIgWLiSO6fn79kHmj302sO13FzG/rttivkHMwJCl6z2ciuX
BxG5Yy/gD7QAYSPLT9rKKJw0QUujyDdmxFrZpAy0S8ydQJfNIXDYjD7kpvaB1cuR
yc6tl8pdeGzmini0lAHClkn1aVAKtzuWuEAoXxWhDHWncUCHo4vDqGeyjlEf7fFk
JQUMu/Z20SPGtHKIxh1A4ZtGwhaMoB4KZIQ6cER0hTNe8+zSa081YYICnXuZu5g5
pbCNLiMd9DXO0RDcWmhY5NMwPv4o4zV3rfl6sUITqaHGSMbEZJzfoduVvNWHSTR1
cNdkWUMY85ZGl3K5+pd2K7hWDeLqvtnqJwaHornOGxNH0k9eEzqycMwP0aswLDMv
a7PUtqNGdMlPp/GuZU9jgrUYUFIWmItkryVlM8/eEq8suY3V0VPff7bmEPtlBjho
+IjSPGrt74upKliOpyZTAj+Mrq8PzMO4/qlNOkmW/ru8tuauK/mrOzRxdombtHtE
3hKFzjRfs6iK/JZ3DdRHiugwHa73PyNJYQIyvRWhL7jY5opIH0Ux1tC1IMXYS8QY
1qR0JSCwwnwF8uF1ngPkyrEeE0yUFININrWmG9QmWctxx7EyzCTlsc0FaEw2dUEm
hHLz7hxTMC7gq6dPXGbHxwemhca+859TX7EJcc+Jbvlfwl34qhcv4A6G85QK2WCO
ttrXfQSd03q3y7j3glYtL5oBxL5XixGGlXBTml89sf4dPB6mO37TBsnrMOE2sqZT
8H/gQVnP7XqoEM6qyO2bjN3rGYpuD7ArJjWRtXaG4WOEk0P1UvM2Ss93JF7Cm/lM
UprlpMaz4l5NKvUBiWz4nW1EQUp+skyBazNPH4QIF1jLDFzzahNrdQpuf35yiCAz
TBI429EtdfSNixeYmjrM4+QZOB+D/VVIHxjHkWccGJYGFxTNu7AIKP34CSWO2P/D
sWKRc4+1U1MeLk0k+zbiWi9msBHmkXEyK+iO8eXuaU0QERXCxDsMqGA7QTs6ypQE
dttM8I6DBclfZVk8HZBA8EqZApoAwLDkasUeJS1dEwaMpWMbCMapMu9PRDDxUlki
LIEwAzAmbrKnG7k8crUToCoISQm7gmMb1mW35M8Ctm4mRqatH3REi+2rP0NkqgKb
hEaBnoWzB2vWI7NH1Vu2hKhgWJpXv/P8nzuMRIbIpGO3YRJIrtu7ueWtQ69i9Uxa
LaK1ZDHFCrhADNQAYJoUvXLKiWCX9yfscFsZeKZGO/55y3+FLoO7lQ6ORXnv+ZZT
wgZDvn/SpPvu7gyeyFP2/6mEktNu88aML6mzfxSmjbTub0UEhbMIv04b8m3RISqC
SfApd56nWIA0r9NTnMxyhJCLHmEqUF3KwCdBglv0zIq3wfQeD0QDPKAlUwiUxIs6
O893vvPnGTlXzbWTX5INN+qCvMcN2vsPAIEhvRudQCof2zXn3lp/t5U/KqfuzkIF
sW+1noVpEWuaMihyfsEKPM5BwYTrjkezwRuseU/F3XO62EkBdxqjZ7Xq04VmpCIy
+7r3O6OSArI3cnOw6uB3wqDoX9BHqizPRsUhv9xY0JZk3aOy0NozkmtdtcqyUV2E
kgVnwCgO3BT57P5z8pJmueQnk/vClPK4nItGTVC+d9V+2VaeBwga+Ncs2zKhHvRC
wQkVUbIhB4nKgq6S/VcS1EBJj+n+qMqxaKQx2MpauwznuWFxKffTysnb0gIbExdv
V0Gg2RQ+b4K7m5yq7JEO06fm63gP9thRTsJUUUtzDYo0732gr8JYabu2v1dUiJzr
kJKMX3sbL0nq+La5YVYJi5AcFI2WSUHfxxrMJGiMx9ja+d8CdcL8nYSMbYtBYtQ0
Zh3j8J991hpOXJGtU28eeCFJpWiV7xJqz/fX/s84JoSBhKC//cBT685eWmBftvB7
sRSezK/k7fiIRyb4UaFaNSSOQspSVoPbpLdf1AQ+aee2c3aSWXa7iJ0u9vVv60Nt
kN+UzGjjGbLm1qFFjKGX1MmSg2q5jKtW77kync3m8TcVHXszofwvUK7om3kiFMS1
oJinP+JaFXSawxvRDtbuZdQYb3m8freLS+7AMiQNbTAUmKe45Tlxl7b8Gpj2WZq0
SBFO+s8534OeXphNJ4OaXlqvJTKt1vPqRAyPCMrMJC4zK8EubtnG5xrh87hamwlS
hTOLu7nBgfBvgm7d9z8d6o95100ylz8Htu6oFWwcaMin8EXUedFs/U4q9aAh9qch
M2tdJpO4yJNcQjTDjAvDqSCB80lH3tIeT49ohT+vmiZAsWOtUtQsf+eWxdrj0m6u
mWLLCxL5sD9A+duzifFOo5PAUAEEyAAxxYzwuVWHF1Wt0Xi1bgCdrXTM1l46Uvoq
R7jl07vGevLrHQwnmqG/C20OC5iRgqJVbePgn1qh41/5CaOvTHabRM42wCKWbDg7
fy7BDhJhXYwaOEa652IDIn2h010wIQ/phm1QViNyg6Gebw5yZSLDOTCQEWF6oqQB
FA254zfuQ4Bl3j05wFpumPZZx3g3FRjww5wRA6YZUsw0mClCbWuTIrUwQhT9pGFO
agJWRbZnW+C/HTFntKUTKf8+WFjS6yw8+RSJgmcPH1uWhBFcd35ZoohBEwhOntIu
UPa0zT9nDbVgLuA6XhavkyhxE+Mxrfb3EUt3UTpL+fA8ThQEP1XRlt2elPS1Z+h4
pVmTZSgRZNlDdlYfVQT+rN3d4L5Jl5TUTP5TV47uQLPpF/RzMYpKhT8YwCMHLdfM
Oj7fNjGRnt9kgduJtUGTn9hGtNcl0zuRHnloKYjl0a7c+W6Gw99g7MJ3JdviSOv0
yunzthIdkQ4HAiKWImh3dGiFOBO994eoLPeXa6CYfAxPN/Tc8eI+WC9Jw74YErmj
ZcG2AF4SptdenP5Zy0ps5ai89AJ3O+Q8rjxDgESGiQSik6nmMy9/VbqfHe45Fr27
Ky/7qVGWbc08V/VUI2Lku4SwhTS/VyrOZQH+CAKaXImZLOEFPcB0vfpLHZRJy6HT
EnqcTFi748P/7vKNhAjrAN4Ph58utslY4Ps5iMpSs7iK3ZcIlKD/gUsSaYl8K2PD
EAtlxHCQ7iITA3Q+tPym1/0L9Xe/WfZE44K9Lop6nPvvjTidcfBn7nkHD6EYa5Zi
7o+fBOC/U17Q/U/5LBR0odYGpngZsh4rRdBl8XnGXmQM712NTmmTtnq7AMe5EPR6
OUP1wqeYrceAza5L0qOvCFD9HjUdKFqSPazbOIB0ZM9W1Ymyg2mxVybp5btKV5Lp
n7CgS+gUtmbE6b8inkvHD2UIF0r7H59RgzLXlhw/Z15sWLMwJz71R6tlYUzX01EN
klX7U6gA3ZZ9lmOtURasZOw8FT6p80IGSgHR1v3kFMfieNWJtegSwPsI1sHsHiQ7
gG052w4yYmoBJNTtQtt3JbaSYevwZ64GZg2VB4SbaaX2HR0C0u0jxENPmZNScH3T
/6UKrpxN5GQYkP70p6ku2i6soDwG3ABQ0RHk2mY0MJvn8gWwWUmIkUG64uBXdmnJ
YtBiAST2OJgG9ZPazMie6NGKen6IPVMb9LvLlR3c0+IIYpmx3LScIF7kfimXqx94
F3UQFaBuAZh6ieyrXa4oOjRzfI2xzDBOaMMCU9M4ChGGKfcL+4lNLdCpZZRM1Jog
3IhZCr/kBuzlscxlcq74doalAQCpR5YsVHY5i2NFvvCWPh08o5V5LowT8MlE4qAE
1IDIMJzjF5Jk+rS3Tm//wGO5Gh9YYUmE45Y7CKvCMKVQ90SthtQFQ81idnzHTXWk
wxsdnMb5QY5lijGdI/JvPj5PFzbNfM7zpn33sh/lLKKlEvtVKPu15HA1XOhrGx3n
IfLYZgdXtG1NNMyt2K/ML4cuZhneYYQKj4ViYjYzlB8MhAm47Oe/f8fTWiM/2WQa
6JnZuesvO0KTm6r29BZFymCF4WUmPjIdCef62OICMx+JJRKHUdTC+aAKnqJ834W+
TWi6XR02fmqjdAXkx08D2nPfD8jlHS1iktyjsameKXHXNbKdJ5B+Qx30yWmioYl8
f2s9q/rbrc57v9GFvbqhByJELMXoDI01ZHBFZN32MJ2UUzLY8bStv4fOpYPCHyHx
bw1XCJW2QAEVf5dV3EmxCtdDhkDI3u3EZnRDkJ0Ex6zsQlxCPKLNdPgwyh0hKFRd
b4Z2oGMVdbBZK5se5q7G4lV9uLYdsGMrdj5ZjZso3suB4gh7CM+UzB6QeICILUik
UOP96SKcQx2CrC0a2wF/9TFjLfnegI5zhZsXxCXPiyeov2U1IWSaLZLqQlce2IH/
65RD8AAL2PE1+Dldfm0D1s+2zwys7U5U/hvHci4wifdhDmsI8PcP0fsTOUrOG6Ou
V0O4gwItqr7YT/ZjLqxhJFm5GL8kUvg28+QZAURTFLgboNehv5tuZtOTvip8mETK
qedhCOhqEvkuxsf68cV0ysi3wPZxBokYG1Y0oRliN+gdD7qsOpS/HL7bvNJxuaXH
pQkNPlU2MrERPf2lWR62AaHjQGNwqRu3zHVn9dz+zYj0BcLQ2yvJ1iL7rlbCztZI
DSHgC0XULqF5UAv/5i/Lpn5lrJn/LbytEFj6k3jpqAg3sugnoFUoCa1kzifl/KX9
Jk01wOLWjJuojq5KaZwGNRtuGGrJTT9nsP63nReQ9EFPx2KgQ7FXvbMHp5etVFWj
U/BomgGBfwI5Vtt3Q6nm1+OXh+7FtV6e0JF6D1EG8/a/XCLyuRTNr5xavcwnlehc
8iANymdLpzuvzYY4d0GSvAUxE37Y+urs8dkUe5VGhvO6iU8QdMveNEvlBN02xSir
xLc+1feE1oChcPrGs+JR+r/nVDFFpna387X9WAPTWwHHM66WPSXnSph/8YtvFxO2
S7efyNRXIWjHrb/hUvX93w99luDPvMTctllmo+WkMIY2/X1w/C/vgS38KJjNyo36
mX+2HLvW8IDbNiKtjFFYRcNsts9oHGykZbbEb7fzZath3p85+mGNRUnYo3KfynJn
klTZA1owa1G0ZlMnZArDEaMPXyqaS0W59SvA8hTnLkl9tudjNJJYfkCpOLWXGPjt
NTEeYVSY3KsZ9yNIwi2AhSkFfi/dgPCf52p8CU2LDUF2+Wr+X1GFa2Kz72R9DrI5
APdYzP7a/L9I/BSmYi4WflwqIU/TxLaeZ768oPNTIqcsLIWNrt7fF8F8t5AWOmft
N9Lr0epXyZaO8p1XOzGOE/5MTXaU1qtgKRZlihpzaf8xh5VMV6pQ8D35QjYXi+v5
JVzjd8mkBMHhZjd0LQzIkWSDNh7Xgj8A0jLNC85W65aGzZT7C/q6FOV6rFDnvJ/S
Gz50VmDaiQ7LF7qOG9xMiHWUjDkKUsRTSk+nKjSPsmpE4rfZe4H+Mb5PVHOdmj0h
5sriucHu+V+3cnFnpjqLuKFzYJ5mP2zDQoJWefXotS0SG+pUPKhFP6Gy6Js13Xti
G5abbUlYbrKCGN/2rb3y+cOUDAdh0wmmvuRzBU0K1IrRW4tE0+0ZuMZiG922rjtb
MTqxLqz5RPuwlyJEuODtB/+vZPtiHVEO1imLVLPCpf3Cvwmkes/nEfgLxCSQkj5N
T4sUMNACAKNhfjefU6b42nflmXSXil/sfLAQqSoDY4YDUTIecdXcI1w3C4/G+YfJ
Pb/30ZQ7gp29xpiT61TDEbzOayOX8QUBI8iUclalWBwD5HtSeEIQRmsW2H5TPCYc
s34g6ssp0RMPluxUnqHjpUPiJOwvpW114oQKQn4wLutME5id/FImv2JUbVHFw/ay
Mtj3R4i6EfRRMSjbZh4qbxo3UyMF9B95gJCm4ZwKEEpCEYrj0kU1T72fXhFhXfR6
Kq5rhl/gUmZzSW6HN1lJ3CwAmv6r4laHa/X2buQ/xC91+/69kKUlVHePccUjUW9B
wBiRKGlh5vyZYSIEWwrH2WC94ObPw/ZvCH0qvZ9x+QpPa9IdZcf5soRacZxYzlvI
ney5tza1vE2FPEzwNLAA59wa1xDWQgCprgJGIs+F7RHculxyNjdMkUWweOx3y+OU
fo/5qujIDYhXOWK3bAnaqkl8csa3k5snG4iR+Ybuu3OsFk3BV6FIiZhn0jmoWEhO
T4b5xe6P0Vh5XBBRpmL/5YdwM580szzV1l9X10w4KehRaVvuGfGV17Gc6biTu6ho
Nz7Q36X1Y19J+wlu539zL9kjA0N+CexirGTUf2DoImCgbD7ihkvakePpm/U8yN4C
FpaGZaqM3n64UkpKVlgU11aMub5XtsKRWDMOwZl0mGb2JM751zIU3nq9nFkiq9RD
M/OmRMWcGYaJlyk8reFVBlEB9xbLrdxq/YT4tcpCcMSuZWTTCO70ysWN2DZeMO6B
jsYVFFWRIUU92pWvuTpmHAfepfExccgSuKedahfd+2CwiQEaTv+0wdUxK8Ijdzs+
fBh60NGzYJdqZyvtjePCrgB4GZp/LEpcg3My1GVvhNYbPaej7L0wQHCPGnG6F8IJ
pRH28CtiKpP12+Bwjx16u3xDAnkAhgEpQyKW9tVeOcDB0JV2H9/yJsyFb+6SYpKM
d8PnHNzZtok0Zwp6BB+L/L86mUd0wKdgfmyzaxj/sq6QJ1noe8lZv1uNLWThBJ+k
GF0IixMmEzglnLjf4GF+kofgQNm98EtKT/b1OTpwfIxqI4vAVnrBBJsVRZU+qdur
mqZk9hTfdz3Akp9Kro8r/d6RMjIXhy4dTeIxFJn4h2CyltXRGJPlvbR39Vilioi2
yVQw+D3fDT6VPruCG8cYb4rxnbpF38IT9Q6IfYlX0CwdfNNmqgm7+O+Se9bsmtYc
I7CXCxmadFnEle5rKMRNbR01Mpxj71QA1XIHx4TFK/ZZwkWMBQAhdk6emiVs+FCa
rmreg/x0zkdYopUtXhNy2kVJuXUOjnRfCiTTCSh3bZIFuhTIrcprfAA9Fj3r8jvg
t+BZDiB29SnUrDm/l0zNC7GL20O4nqifulHCKyJyobHSdgXHnwllGy5ifPzncsIl
2dVAie3P09JY4Ao5Rw5HlcBmLhXwursZFubcDJ1BRvQ+0iJKnxohoNpS+T+x+R84
Xugu9a7v+60XfGxtVVrFXdZSgxYUMWu8F17R/s/tj/T7SnDxlDoSNYBWAtCxR7A5
3gcGc2T8e+q8DK9lpqrJKhpVdkymAUdAdc7I/vMs63ola6lAHsvQlT7jTMlYV6Sy
Z+2FJ7iz+ZY+7rl4cidTmwZr7Hqq83S7Zs8E2YsS7dVzlpPPxF+ZrhGSrwtw3fgK
8sQtHlRmvuRxfx073wkFo60hSlulFTsNf59zQfVHMkmI/h8AqDIHi00nRRhqKFOo
KfJMyhC+hDO1Nwqp20vdSvzgux8cukELKYLu7SbyBM9naMbWx+81ztwPWvHS9dwW
8lUVJaynCys150uvzYi+uxl3nDued6x3SDni5ucu9HkX98SBWuFYeXfFkpfnzkUh
t5gfDa1guv8dKyNkmLGKgAwsUQBRJ71YX3iaDBv6SKUeDTdTD+MfaKM2plIXZ8ho
uvcsFYQ+HnntQhiBt7QjuiIEFuBQli1e8Kkiv3T4DLwRIPSAIoMECkpbS+HPFSq2
C5av7iRKGSvUldErsMjogd1MS2OaGG6XD7RWxcjLwi2yjaA387cj5gE+8SL2jSZt
PG1uMnv/fXKHvN7wqZEuXqXRg7Ch0W3jW8bZsAArqwofbS+FwuUXEmTnAuScK4m9
YZHZMw9k/1BaWl7YfGi2WqRiU2QcymTMGKqSGfx4aJagqa7PjHYvFdWUrGBBNwl7
nMbLU256M7x7FAPhoOHagWz2mSiWYPFXeKIKTCVEIqilyB3NyKfqMLHO29E8VYV+
8TFiCIRJP8fLQhncI674pc098EbXEDHoIpYaAbCU51B7DqtTPJaUsuEaMp4U1Yxw
7vHhgmv5lH75hW61BxNPACrTnbvlmo7IrrjTFI28lNgH/KoZ6cIhtMubN2M2YgJw
qyEzq3gM84FKZ0PlkQ2DAolhoS5QR47S87iemw9vGWMgSiTvld4nPGSdL9uVfNYl
+ewe0IwgZ4d2SvsXH7cYMZMHY0YelUqYJ9N89uTPKyhFqiUMtSFW2NU3gxudmsIP
Oy2xkEZ26v8vE0mBJ3ORaUqJhlK53I545KgegHarmgLuYG4AQdEo+lF2oLilmHL9
5VsETbvnEdT65Th1Qd5N3sGkQSpTX6Ugv+vajag1BxtxWJMVIP6zBPceWowtNrbp
PLlMMVeQ2Rc+6AVUEmvdvrqeDnnU9Ozn2aOP4UEVGSHxY/HE3MaYrDl/Fd8ZCMQS
ePw9IlFJFt5LSWaHSn/tSr1b3NwFbavW8JRf3YIYChRrKnej8MBPvcbS6meqPxOs
G1DYAxq9ibvuAOqdx/TPR5Cig3sJE8pn7OoezZvyLZC0rXzrP2e7jdQ6/Mt79s1n
xINnrlDrEZHZmTY7w9n6etJ1mCV+XoW4e0d+yNrnpk29r/5jJgwN2+VpgVe7o7Ye
aPGTI5YpaNZ8SQYZ91RC6HFoO2s3k3I27iMupIlcZm6fmYm6zdfuzjUjbEsMRtWz
DlUL5UGU1+H28/LQJk7Qsi3lXeKP/8N1l8ExlKLJHgyr8vfoCffK1QW867CR7lMf
7kJve2fzl98wyo7AvlY0/E35jLKk+y4TF5Z091qJ7PMNQGAQl9dJN34Qm5Fjk07H
/Z5KUtUQ7GMZ0pv6E0U183Bn3hhByWkPQjhLqH1iamErM0XjijGd0A/4ggkUwfsQ
JYBM4EDF71iUdKvrkmKY/F1M33ISAz15ShNnf0dT7vCymDCo1ofELWMNWarccQ50
OjLZQEr/1eLFOBO0dYtmhnohs6aoXfOrANPVfjv33UntTo34vcphmUarZRQRsqHz
u7IVyYjLkfdFRKt6nxdhCDLfuUHlsRohKStg9DGKMI7IsTnpWNJUPK3bm64B/hYa
v/IO9xQNG6IH/SWF21Oy58tSkAhqPmrlQSbkUWNWOJshjqUWBUAW220jpR670xtH
lfnBE9pKkeJqzOG5Okk/qN+EdWT9Hdk6oZRt4jCWEi8G9uaEbdMgSRdHrlCm49s4
+Vt9zyZhLT74Byweqxz9mOLi38kTBVUBW4FE/WBfg605QjBKYR0O6ma/89P3l/wq
sjEuPAXaMOg9gRhi/MjYbmBeVbb28txeAxWlrMVIruC10fpNrjea/38TS/TtmCp6
4COBCOf5ZhzQG0wkge/oQhpP/uTsNNhp62S5Hjri8BScmOGQzz668CbuszLWem3O
WuMQaxuoFIJlPRFuM1B7O5Lfw+Q7Wz/ScuXaxelb2S9xmV7ucJwF4IHp5Clms3Ol
oAc/9FLYkkrxhSfskOR4J6hzZsqWDmRKaN9U7HNhVZGVmjiZHJXb0DSTgs7WBEQu
xuAKMum3X0Pb2+HuOeJvTpqA42ClB+MkvkbyzdTQRCizp3ggKjJ4oLH66ppKtQ+3
PIHnNgMjf+q3BcKoqb9U/ZOkKgHaQ6GrxlR942OmIARHfJF7pzwVyCN8Glhp8uU/
SMxIEwhhChX0CdiORvdHZCFVGhLfLhCuIuLll8fSaToyh/49+pIZmkT4o1NJnLwG
2nGEW80Jho/A1zXajYYKG+HLE2CazYM7WNI00dkC8oVf109IEmV/Zflr7hfIMKcG
24wAdeIDvYAVTSIp/OJ6JrRVQyCNBRwTWD05P7vfT+7QBwCHnBZzuuwlXX30yb1b
cy0sXXF1tRnDwsmcVSiKCgS36D70UP/Ds9tBRMPbyhNbOAsPRGK/plMa/MWB4Rxv
8yzi4xMAXjYpdpBs9samWLVkGyyF89t1bAmrrP3jLwklgapC6ZKQ4fTr8jDFWcbc
5l+5x8vonUd0lb+Tk5MBp2evRTr3FuVbFyCqWI4wuUMfTje0/aMn7RqyRbRfrVof
XiPvcBo8nYzqFiqErWUXA+X6C3gC05TgXMplZL+nuiwARXe6McRX6+fTnCRxbUTN
tMj+OeGD970D9CLdZAwvz0nXEqehuN1aG/2cQmkLZLgtnL6LlvBn8osQU3I98yAF
RoABYog8c7cVSZJ6bWuv1pMBH8o5uxMo1rTrEoFIEnwTnlARxiLczzfFW4rRADX3
I1dwzBw+tG8d6HGOIwK6y/M9ctgWZQRPZx9vNC1sa0xxPZS0bZWJmOSpvAH5OL+8
sA6HSkNFUaqA7wAS++UYxaP2Mz3KZMeLDN+q2ljUaCDwOua5gnUcTkzEmgejwnbi
8naf16vd/dgIuH2tFFAr3dO279RaIz5vOXdUZ6Ns5/2GtXZP6k1k5B8jJmn3TCRZ
/5A7fSaIOT16LjOOefj3nAI3GiwuuUzeqk2xlUWSjJeFocQOCuPJ4oRMODShqQpx
reE+IL5xkEL/uSEOyOATL4wjlX6N9ri+/Upkmj5h8y9lw6L9Z6hNu3M0NKErx/MU
Awt2yzox5LqMWSx9xunS70eeOzFA/Y7GG6Gf58gdDI5vUTJJ0ewbSmUUqIj4eihQ
DeVC3BLU8adJNkyIwQjFov1xkqStu5kGbJPo5/NWTcTkm+zley9lFQOCN5G6moHh
vOReSH+IcpqmQ2n3qKAyI80zoJpi6shdrgxErhO/GB/ac8gVN4wdyXhmvjT88pZz
oEj5oIjDU+Ez6xak/7dGzyIx0+5VMqACmJvGqz15cLsaDB7f5VDWobw/b9w8Dznj
HHfLiVhrunSVkCB+zg0KejIP/v82iQP25IGgUwyyGlMSDWIzY+48m3TdiOAB0r9B
U2MX//HjglswJJcbiHFbDPo47ziZERh3UY1J8KjFDwkZ659cRog4omOx8OKNTJ5l
brS0APqSEfgqUBU4QqgoDu8kEe6xGQIxW/dHKp+DaKcNT721Ltg7nPL7HtduKJmG
zc4zqee+8tlrTH43vD7xuGSVlU1gjbGtGUvUx9Rbs0saOilo/MRXFdjguUB+lPN1
DdDlGOhWL2Agns+dpU/JDLJb6MODGjO5ruxWXg/kv7v6Avcak86+nfbmOn9lpAZt
CVIIhfOJi2+ioWCChQ1vTZen90XENGV44jxh07Wdn99u2a6Ccd589xY8sC4jeWzP
eVIUaZDI9j9/OtTXCgcq3cI43MXPi9+mnUpZj4mjibgfEYYmFBERhldsSw2pSd2a
VqF0QYnfd9sItt9W+sPGguBAl7wX/K69T9tVzmKc336OdyiK3XrsxfA1cQCjongo
7s7Dp5Uz3wfP/s76wAEFhzxiQggsIrIz14bigu+XvqEvoXaKwmqp3/IKQBplSY2t
ieCIcwkzb/KQ17CFCdzCEo9pemcj+d5lZmj/KzeSJlgThBrl5gjzM9licxJ1f8a2
Ph6sPldnSPpLe6hQwuI4WN8JUzjA27FfrOH2YoFIqV1itrZ2muUKrwYJNEjM1I5f
AsiERvf0mLZWa/uDy+FAkBXP36qO97Ot9O/szWHDsUbi32ZOW3R4d2Kkiy6zR2+3
jHZ5vrAJl+l1MfeIjHjfiRKALigKC56Qcar/j72vUmRe4GX2rJtOhd+/vlOzTEWN
g3wCBM0jWbz1y5HEBe2rE79Vf09KDoNopgPbzOy5QYwGQhX1O8xrtzfWPx/SmHD9
ASZLB6hyLtYTinlvDl+iPc0vavNnC25QpJ9lpZ+MbPvoM747d5y5inFv48qED+bR
vmYQp1dcIstLa11h+SlT2/h6I2zvO7IkZ31hVB7EnBniaysrM2jkZi99EMgystYq
7at/dj8490nx4yCwP6MhxSpnc7AXZnCRDvW9go/aWzDGiUzDLDOR4QrNIF+E8xQV
/Nna/BI63s5EIHB/mCJf+NE+U+gvQs5r+3P+V+C0YgY2caUrmsUXc71iXFdK/XMT
69k3iwejV0OmzTgls/Pokj/GJ14ywgvPZSSgG7Ue2VLWWRtZiQkt0BJ8KNgQbcCu
UyNEtrjusVX4j9yv/FZGltf0tAcYmMl8Ks2yCvzPp3ZUzRlAkKYWXfz9Q3XBf0Hq
EGZH6FAclBj6KQo/gwAY694226PXCZXvS4zM/x33AWpYUhox9x+p/XrdVYB35O+D
WB1i3lOoZqUYmMZiey0XOb7AXLvrAdu3Xb9Fdls2SkY5spAF1wnFLXf8eTgie6s5
kYg7zH4Kalhrn6jRcQx5SlpffX5J3maxs6Phjy42BTz1/d0mz1HBA2Pd+IswEgjk
uYiSPhLvc6IY395bOJLWfhp17zk7vehifo8GFfAcqYbRcY/TxfztNaHlJd5O0tQl
Ssdfqa4VhDYzEzYAxPwlg6KVv43kEyLPOpreBXSFcCQNqEPqHmiLoIIiDzjJT8Bq
nY95xCUc0cobuJJ3O+A413JYT3eQ+5x0OcouDUYGl3+UigBqzJ8bC8Fz8LCO1s6M
b7Z6yZMdwkccSDRIJONFjBkxSobFt4eYPDhCnsRQqVh5mNh/LsmIjisCjCCRHZNH
P9iO3Ih7lFA9s7JW2RB/rqsCKEzsxfOmV2ud1ykIL+cy6/cPcusqqhJd5xmppcKV
k5zQYJvfh03XGCQ4rDrswJ+XSnNF1caWDWoEGciTi1TQurkbr+YyMYCIHZTPI9NB
opB69yvgH8+6a7+zkLRWNRrbOzGuNcpyJp4/iwAkI2g5b3oYr91d3m4bU5Pe3DpG
EWsbiEcqULRM1D0pf37bLA5bIoyBeCwM+svm96hPnKOPXmAZSfuRKhgscKT5ev1H
BH0qVgLkSYisDA3wngXFrWXmA0gQ3ys6Fg9h9YI+Nh10RVmfKLVLSRc4bcJgxIwc
6jdBHYIiy7U6hu8oyYAnqvJX8Sf5bu5olBNN9VwDB00j4dnd/KTdeW43mLY/btrs
vt001P7sIrtJSee4YxMDJVmUnPorQ77fIqcqenadxq3U3DqPHS9iLVNwmps6d2Zm
8J2xhxRW22xhYbV8Z9jj8CYhQpRjR2f/wUdvmpf0Cu/DBeOmqpZlYJ0bxAOvaLbY
Cf+w3k01qYFlzJ68Qaz4ppSc2xvZKfV1cvuv2SgHBeAYz9vJuAIrd5vaOrza0ADU
51y8T2OwfN57NGx/C1JH03BOOKhZ4L6Do+lV6H8+HYNxDXSwF5oJC4Uq9o+DiSWl
A0AuZIg6MYvmAT5tIWoH6uwBggH6fRLbU8dyfP+xNwdVYz/GDgsNQuw4DOs+Gnrv
Ivgfw6T1lZa4/+UQ7aDAQ1SevK9atgoKwPVcqM4Pj58iUCmsQpd4G38YPtnhki7U
V+ZaExQThMwt7nyYuVh3aRf4jEyvlswJRzojaI4ES9ubzFGj5V73mlvgWkH5Pjch
sZginy65ljLHcPL3e0Tvwwlr5iQzLZrqC8T6T7xeNS9LY1UQLssWNFnRlaCLAJnc
659jUcAdJHuki2N2CEoj/xsoZSfWjhIOOApd0qmgwH/rPIdz0Ee4SSgBiJEQ0AHV
JdyoyPxvveryzqCJ1YVYQSbQar7MA5y4qAvPUYIgpm2NoHu2lRlkRIF1Z0kQ0FD6
OS4OyHimoH2p4pn+MaTt+DfLCq9mj1K6Pxk++1YVAnNskta1s5+d5HJiW+UlnoRJ
3X6U6Lww5UdHS77mDNiHAMjtIn569TaQkLl1uTOzwHvp1pz4K5ry5zyJTXAeFli6
+Kw2mvvGopSkhIR6+InYCoiSqJro7PSYkWJQHy/vCeFwQmrdi1DiZjmo+Eut4b+m
aqp1Je4V3bucbS5rZkexhSNMfkosDHQSd6vnEeqs/fqVXBHI/+4G4MUt1/9PMw27
5Ph0jAvStNLmfNDCq/0gxNBXKt8jxZJZ70k6RYjhB/W8tcA2HLkCP3KfD1ixg0oj
jqe672saV+4+fx0Ee3cbjSZknmJqN0Du3UfKa8vU0hqLztvWIGdSfEGFsBS2Lfpl
Yihx23NWMdItwrmhGlpOyX1g+qbLsAsqcD+dgyWtq3qqa6d9j2Z51tHqwnzCveS5
ZfRsHb79hVoOM+98QXzlb0ZRqPzqeK087xijQJdvxdDl5BEL2zK8mX1w4VFms0+G
oGE8ZzDwOQ5xSOXSOf7FQ0YpHqGjk8X7P7YQ11dJJTD4dekjIWNBN3YwR2HI3kWS
mBXn2DIR8mXl5aA1jC/UM6jNylNG88z9UR4WgE+fP3n0SuHhRuDgojX2TXjXS8Rn
lqVXGygNhR0wzo+TCeD8xsJinOTZIXXjUHbdY8UtZ6xcsFwlWRuni9+yFj2JvP+v
6OXuIEZj2QisaNz1LtObJrAFYtNHMdSqBO8tU8u6/zwQhgv8M0Bj6At37ITRxlP/
GBMMdVgrmw+x2/h/QvPgs3OU63/sx4qFGYSVxf+buwaq9/3sEG4rDYSA2P7eaDuy
X5n4i3yfyeYQ5u/dLHmOK+5QrcV2aFNA/8bdBD0K2A7X3cBWrU+Jug9LHMUBGtdi
Q3OsVN0DtUv3IJQfcXU0nFv2wME1gqD5MEwC1IXzG+hfdqlx6FGM/LjfEJsmhLYJ
ikhV9TiSJOgEzX/j8zaJbxuU9SuXxjANqVVQ4mNF4SQeXHA2pmcu6jXKN2+NIsGQ
tZsf55cbxTi48X8HK7HfgHEOUl6u2DCuu+m91V+5EGfCS++mN0EPEWvVwY+SI3eh
JlnSvD4apJ98p6t9kyB/8EQTRfkfdLMrJQz5esXs2IlBpersA4dUCFZqCKD47hR3
yFyAFESW6Hfzj3ULZ2Xs+YvyDSGGMJuAKm+2WekmN2/3ovMkOGwFzM7Mb9i5cPCb
1FRC/oTV9k0zep1hq5MROBlqrE6eyNtx5WKpR949g70CI6ffplNg4SgKvz4euPfu
RDZjYaSRNVi09mBXQ8+SFELUGpDW1EcytQn1Bse9R+XDXjeSd9Xde0nJ/E/5KTpl
LEWxi9U5H0U1q7qvS1V5FC63o6tFoUFIVFEN0taVmsCcBw5OBs6LQkmVhyqzmouK
jM8JhSN+YncKBfcGuDl9jeDKY2vOD7PAxgadHDV/8JfeCDI2OJFJ2SWea8mF8m1h
TsaeVXZSvV//IBWZw8edf25s9OsS4xTGmlGE/jLujVvzMt53L4fMD/SYgDyFuVPR
SrtytAr8bmCfiHtnsxgYx+Fj2sBBAFjEMEEu9DFJ7Kp5Wz1lewZpMVVjov2MmKWm
KmZYZBFWn3x52aziY08SgbbGKh/wl9KThJu/ppkhqgmcbqDpegpFyCFPXlLThY7K
naL4bcE0G9VtNbZYJzDhFCgSlap+e2dcGj08K00pNi0yUL70cBHbR6guaWEXcGnY
JqW4A5iuC1zVUnykH2tgQ1cSGZm7BQ3WLt2YALJZgdiQBeGtRYMi8511mJoQDfeX
lenJGyRKt6ZoQPKHHw1Pd6pOoGWWqADDJ1mMboIhBVCmP0KsvNCX30Qjqm4R85NI
b9s5mjND8+0eoGWOsutHTa1P2WC2+qJlYLumpi8Fd53CsFv9I2RyAiAjP2wHr+0X
YdJbb04iJp/hyDku721nTdW5ER/2J6cm3m8U/UZJS0qdDwpvE1bJfclJVRUN3a4k
4gTqzSa6H9yiqzfvKnfp4/rlclv+066iVTl8E3PpeL8LwZuwkbeZ9Lwwqc1i7eYS
XkRxNTVdCPIuBj5Xlzx4r5gg0Y3DDcufF7w3HSVIR4j3QVDJNElAmiUGtJ6qTSdl
RAEo3q1/Kqu/tSQgZXuo+I9loFadqlwCK0b2uIpSPADTlIcoj5cxemGHK7Q8JFg1
8+LnOsPfnptvyMW7NF6LsYCcBFVgCDDFaiNuqfmfN742sTaP784lEZXO9YN2+1p7
0U4jmwj3dL8HoTYDr/vPBgUi5ijb3tWEYoIhP8OJarsqEf2t2Kf/HKBSqSKFZ5S3
PTpfwwrdN4Ta85/yWQDoYdsOOyLlYSUljQHvGC1zK9La9JJQjuIPeNmUQ5IjJaoW
eiaRrPDCqtmVvTrJYJoScn/ANY8ncDIky8yt/5ek54AodTEQPMY06bCV0Stiy6/i
/PzwloxILLCoKzMJXlldk/AVMMGqQnKsIFGlWQML+eUqqKbQiin7CiHpSziWaaRk
WeRzPOguBKbFG2oUGv811nCJ5nAgXowrntVXIPvivoadDQX3CbVOJYRiwhw3rAyX
/M7CvZWX0vLAs5Iwu1kHeA4yTGyaDAh1KXh/yAl4dXks9EeQmMX/nwgLsqnhm4bX
FOXlJZpL/I4Ymaf/qqAd+rRCNqMwbFQP0AhkF86TiaZ00Q6lalquOIkAzValh3GB
7/6Uq6fP3dYyD40Ff1fIPojnRwJXFhHzRREyR2n9qf0EP7P2iQee/QUdYNUqvN3n
6/GxUJQ+MVRYZPf3fpQCt/Hi6bf0H+Hs36p5d1u1XfG2iCA63GLWI66/x8743Jbm
OF79/aW1FU3lYm35eXhdKX3LWONwT+FGzPgY2T0ittNjD85GUKEKpzGqyxi1TQXL
x8sKM7VFvV8bF1hCLNfpU3aSiwZJhhcKuo/0mh8jZ0h3RV1c7ZxNBvPxM4xQtdJJ
U4J9aLgOcOd3b6wDuSkbtFuZh9GgAN5AEO3Psx7rF1KJ35KiWD4CUNQLotiOkBu7
uHlwxYu5+G5L7Hnpt3fG47YqnwDfgQXy6JDAtlCywaML8BGo6RE5PmOjdIbAEyUu
9wv6CtGB+LOo3oRq2L1eudtCEXUlUMq9n7gd0fcwIerDCv22auCwd+C5ENKL5BYU
1xahktFPw1RPE5Xrp4VLYE2AGuaP8GeOvYWwW+lA43g5tbrlRuKCs0a+6HQNwOX6
jVobPHLY3JnbYFWVIeXKd9liEK8Vqvuq+eATbVSciAP7A0GYMsV9SqqKEiDj3dOV
tRb7+eIAOaOe7KEtU5YyzF20lrMmW0IzG8i+m98zV0W8U3vwq+Zeh2e+m/E0zBEz
8HNr6/D1m6AVUWFx7RrNLEyXgnZzC/HlEjVOQKmthfKmiOOO+VhBv8y56mDixs18
9X3VGEQmjRNrnBOOTQjHdCz0j3zCft3uT5KZEAvweOOo6aLcv/5xQ4QDdxB3FbVd
MbIxP9ctmJPRMV9OCGb2U9ZqKeaz3NsrTe1KT7abVfUI2pS0daAm1rf7cETpebTF
Db7lMpQMO8LkRJuKvciEWnAwBnQ5jjL+wuhLp1wIH8t4M4NK6+oOLHJeaeSKgkGi
rvbn8hFWeYgG7Y0QTBNRUWb2Z2w+tyWjV+zGKAByFUPgyKXls6aUhx3k4b+IlfUI
qySUMX98wZts+BH+1/6Ow1N5UL58OBfTc1tg2Wlg3T6estWxhHGxUvuSTOJUgjvg
y8DEE1xrCn10+W+ZhQyQYZctldILbVaR2P16YGNPlvRMk6UA5a9XdEhMpQXwGfT5
ZvLuP9d0lWnPbrxHpRLvPfgJQ17NLzOUSZwSGLMaikO55D0uTcUyw2yVXJBxSxlw
c0HsDWws1HssGKegYBDG6KY5XtICUWIt4EqJj4YdEblEsPZ+WSRbfy5kSKAPPRJZ
f4yN7VBO/JUGDjwUk5bkpqkdkUvpGePCf+yhvocRsirTQQp3ZpQxe/Sz/Z4qr3Or
8wE3dzWtdrjG95IC7oRSS20e//6tdsPL6HUfNbVqdxQA+UZ0cZXr5/7ng7Vq6qQr
ZniJ/UtATfOdrWUW31Bw4dIyPZykJC4u7GmEIrm/w2pGCgNnQFHBNajChudYcp8W
zwrLCz+ZHABAEvkVz90ARmVPSgPm7GY0yKNP4NdKp6IcdGut/U+bCCz8fgx6eYDb
J01CwPCHy2PEc+fpnxOc+25rBomDsixETgivR4NS+8XImx3UjB9XjmHCyiXjfjLE
0bLUfgt5Fq6xJsdZ6pCWOGEb9OBkVYAcMuHg+BQvBZUQnaMxrsZAMgly4lvq95dv
fkUSNPJQIi3M8jDD+5M01lPCK7kvv+7WJxEpCuhHj9qgaYt8EFXqY7Ur2LpBs/uM
ndN0sGH/l1rVZbrmuKxZIqfDHxtjnvT/8t9NdkhQzj0cEEbpfd3O0OEcTzi6jtcH
HajpQFRzcd5oDJUD/x0L7pCS4kOF50ubvDxbgr6L8qgJ/o1I9jztgb3Ov3IQUZwV
6xFz2MUFcJQ5J5iZsIqd/wvEDWd2zTJmEnaPyQl7QCFAi3gVvbrmvBphXfuO8f3O
1EYmBcFOGt7vtRf1o4b9KVe7NEjy1LcEvGpQRMgnHWrkeCqUIEgYQNQn+wlb8/RJ
e2a+ZNY9Z83MxUmQt6kJW35RPD5jB0jrGl8mSEdSRqGDAEASbCDr4NyWxHHqN2nd
KQy4Nnwl1gqMuh0hUdKW4z5YMwTQhZF/wFkN97qhQyLEt0tgCj16b/RLJVAwcOVk
DrqI9rmOg8PrikOpQNV/YsF40+Evz8I7Be4nxGicYF5aJFBZH2soQdT38FcSTHAd
q5DKCHprxkIg7BoHmLUKh0biyZfO125b4fSOGp5TDtTAKh/sv/beohvfeoApiL8G
rM/HaueQJD6gkpj1LiwT2Gq1ZYHjj47sJztqV++jOfNBSnlTL4fVCoEON8J39Qnr
scnvKLOqt+cr0M86xL4Q4MqHqerI5lLvsrtjuQH2zGKm5Hxg6QhgGOykHCGheQfj
6fdLhyQoIa5N4QIuTUnU3iG36bHxJKjX9R9OQliO71aWZHEihgrlaZ3OrVQPJNqI
+jfoIM9hjQ3JYLw2JzSHCnmdv9L6GjcgVYL+lTwY74qH+DAJ9Has/I4HvU/EWYOC
RPGB7JRpN7cFr5D7QMXIdfsL4SESN4OahZfi7kuCw1McQM7+pwrVvscuTp52Tz6u
UYqL1AOPJP627gI+oq+yh+jV9kUideVMOxOhZQyUkpfL/bKN0OYo+2i2dwlLvPy/
6yWfe47fQZ9Ixd9h/q4kL5afFve0xNHetb98B2vdqtknuXB45Xbwt41VpazBDZkF
yDLi/wWDfEuGymBOzgt7Up3CAGjfLLXIQXS0JuPtP6jFL5+IcvtpMhVGU9ZE5xRJ
P2mVyKY2BQmPZ0u7n5n8vM8hC5zcAgia8cb4bn4lzKEBUVfzi0uLMBEO1VVlHOqq
7pZ3V+DBR5kkRIXjB+FFGTFf8uazHirh5GIKZMDXmPg/Mu71Utay5qTzoSCTj6TE
3Pw7t28NeS5QxBVE2K1CxPw/MyjnNl3VuSEP4JbsxLVFmCl699hf28AfvX206GFE
BMvE0mwq6uxzKMTERfos06ce0gGgs3w39OILMK6nWCuDlCk41N58gIPdCoYuH1IU
JkANu6qGQdclKj+LuABQRu9biuzS9PJf+jWa5jjtTy1oBB0BCmH3O9w0jgMtdDrX
JHwG2Nbfn564gP8R5iXNbiTRconGzL17437hE5JZ+edJMlHH1hCJ3cteGRFuPYrN
RyUZEO9pvNmq2meukjnQP/J3lpjLDl2nptQ82pyOgQyb+oMZeY41uHhe1uGoZQgW
rL7f5otyC+M3PLRa1d1EOhoc0JzeAdMh2WD5n25Zm5XEoZAXnQA/K98CYtwkDUC6
zDQCwvJRJvetT+hTUHENnmY/Dc343Rl+fNYLnQRQ+erforbVs0/5CVHfxhCcNZMR
5Xm5b3mulq9abnj0F6mbHRHjNGByk6ErDeNWyhEXKkGPRSELSFhnFqjZ9N8kQlq0
7L1wjtcdy55rROFIG0gwwVf9Voto4IvSQAi0OnaTLeHiEf1gkmogxUGJdR7R+tyy
KbMO3kDj7bp8IQ1/ErCCe33ZmiziL+96YSHPKtrpCT4JTg9Dg9W45TPXY9NZ7Ri6
K9M/2GmZGVL+NXbKL+F7JWvPsNUU3bss4611cthyyaMzZKb3l8ykXfDYTxzqw/hE
8+uonpcfEuOt7eOyFa+ZXEPpIoqxrJy3doA/DdHL+tZgFTho5tSL2B5ooi3ghQ0y
Cd4RQhjSGq8YXrRedzv0/NScEOPB4IcjxOh/4vnzqf3JUi4Y5CQfoNg4GqDpZ6mG
bK1rzuXvMuuPXOM+Pkn1QSwhX6AvojZsEiNjQFksswGqzQ+RDRyhfmtR8y5aTbsL
EwhHArZhraqdx//6S7w2Zf8VP2DxmoSDrzinCWcbnl6o6Dt09nP/I4gfc5bXShod
bVBGnZmJQhfaofKsodiwLzYv4iuxFHa2+kcJ8sc8bfQzlOqGAMXYrv4kjCANPgB7
XahxzAgE1k8ejjFmi05oL73GR18l9gjbyOxJTCdG35VXafwM9znLR1uYDyOpL9eP
VZUViOgcsBOlqvlC9z6pdNSd25Wl82amaUvn5QicIMQpWVSoXV4H3EvYUswq6EQt
5EOt/RGAjJBDEFgX95Dox6HCTlo/edFSREyNyreXeWOFnqYHs5q2JmbNT7G9u4pV
ImGpD9O+P2R8gjhZHpPxwisr77unjum4rlblueKLFVH/oKvBz0f+aRwuj95ggMLx
XCltuXmHdj5qcRA0xgBhqD7JK/FlDOAo69tAA1sr6sCz0Vn3K0rHytPzuIHkcb39
wTYvbilAlkokbp2ci7zU+w==
`pragma protect end_protected
