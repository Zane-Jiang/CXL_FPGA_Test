// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0kMVKw3CRyVmEG5lEDqDMAzmTAP1Uu37slrUKIAxuYiBtHTsirXNghVZevG6
i7zGVX6p/PBgYgtJOFx1hyt16bNMndqLdNrwXbtI3jOks8lxSf7xvexJ2jtI
rfhTTBTDI1PRag1PWk8ml80d6J8HeNZfneIYQvEhkd3HC6+bFQteWeCdB8Fl
RmViAS++1SPZ66d82GQ5/DsISz4WIjwaMepf5fCREtighfL3wUiBUYSfVrI8
H9+nilNepKUFa+CigWiMNeDhwOOIywYTL5mYe9BBOGpV68Lm50Cwzo8vZCCQ
Gd0MhHuGC021s05Bp5AMmA5Wrg5RWOlqCCLZQbOs5w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e3umarmfFSF1oPCqRhTLiTcNmDNFzHd7UKfpK0qfArRIXj8t66SavesXsuzN
gvaBSfFkT+SkSQ6Q6g25Krd+3xkY4V0oc+uEsD+w4/X4pHt4Tfq1XH9Wtjd8
05y41hybebPI97DVscONSt4Dh2ZUP2DPP86D7JwEilsRhUX3EQmCU5ZNvVzI
WzdCCwFCsEAwVGHOZ1N15qNtZMEHHn6JXYPdEUgYOYm+rype84zd8npCE8t2
xarrEeDjCfSo5ZEZAEkEnUzVYTYDv3TxPerXyMAdLivYZPi/lhaWrMFNbSJV
rZbeGJ5OQFH6dMchuQpnwJ/LaTP0U7ieokhD0/qnfA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pKfqN3+QCcLOKdCwAfjY2IXXe0tnlQe1i0gWvrqKLmQY2F7G31xLs2h6tTuK
PWOWqAvTt5UJzSkkhUnUKwPzPFFQZCMF20NqE3/TF5Lp04q1+Bff5N0paxHF
NL9Q0XCgT2Zf31POMHGpiUGqEgl/wHUuPlkKcCt3GJVk6Vtb4UQIIwXPaGfE
UTYf83cAat9Ufy0jYA5EISy5J+Tt6/jFH0lvl37+AYJyCk+zzghk6wqOleAm
njp9hQf+lyHwgbIFP/87FgGrQSVW9+ucW+4rktlo8bDBMDBNWeWVztOyN8Kn
hYzdzKoUoMU27fcCxcA36gZwkVA3fFEPV4BE5Bq6Qg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ULegO/docu5EZ0gTdinmhlDWu/zQFwYza6RN/TFzwqfktflKa7XaEHathrcc
qLXxE1iFNvehhTuNvyr5Qx6NmyqZdkSu8EiRmFHFGEO1asbQN/oa7ZnLUep3
j+BYlyDg9yxObA9fbOgVUSGUhWmqph3JsbShNB88GhFf6RHOY8I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
U18iMnV9MyLrTNzZ3FqjSaO2smN5/E1NHk3sVjwhpZKXldTZmbPqcaV3PhPi
9JbYTHuWNCrw+UxGA8V488BwjSclrUGuS3UsNhORYWC8N4qCIywVYE4eq03Z
998GxaFAUpMJwQF5mBPJ6BtIWq/Bbd5CUbj4MZKWoQzaTvLJNsa1yR2bdTEI
tATiU/NjhB4LkLoPZ0B/VPTsgC5MRZVZbVKB7tIeeHud7hNeSjUsU38h8mLo
twvUMbiHXEyC0ywx4XC6Fj93f0JO1edndOy6P3SZPhip8ksHoafp/tWn+RGP
cRTq3ds92YJZLOXn6gflSpqSW4jlyyzJDabnqfP4J0aIsITDycWrvd99kYF5
heEhzIM2C8QmHuFD5IWhLPY+8WZM+b/tbySqrg1AQCs4Ycwmok0ewhWbhUVT
Yav71E+7rYr2kZcA+2Cf2uwzo5kuhdmf/fkotZ8HiRgI7asfkvT2hd1ZmsJK
thMxri3dA0TPh0vI7CL8dkrPnXFM+BpD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eyClzJ5nUTO+vUPTwAHmRwtGkiZjiXwsAgHHPMz0HoRlhj8DWDljmJ8znKNq
gPRKLt7V2vvfYVdtZihMdMOQ9ecgkScZsUM8Zrz0JVfORjI3Tusi/8NupeZY
qDwlReK8nzBgoPSWRA73e3XvrCQEdoRkO/MW5Mqecyv4arcGSQQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E7mT/h8WzPUpv9EtYLrqqQf2Oo3Q66jPnHbLQCHiywlYnDGCs2Jm2JqwiFiG
vNVHbE4IT9I0doPz61y8oJfJ6rJhVolLvtlKmbEIQsYHgloXw02rIz9aD006
Enmr770NQPx8a5brxTF6skc6J/rdTrCDAFWbhdIsCdenCW1BDyE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9808)
`pragma protect data_block
rMhwaujzA99tQzZSfaaVatVc8+FsB09tsoDRnjQ3eRGL5E7STjVsXBHcekr4
yliSU6MjlPuEhW5yVjgeT4yOc2MxoBh57s+/5r7pFyJWihy9HINClTXm2RPo
wDE+4tlRNtIxEKuoH+R33XImu4/Vpkx8ppeo9tHzhCRlF0PqlGZtTF8kpMfq
BjYaqItMdak3uT+YtTsOr79+VEuaDTl/sBNy+lxldtwmc08RILf8zDxTb40V
G5vVFpYsqJTolTM7dFEx9ln7cDgmZNAeaA8avrilZ3p9TRIHqTe7QkmwMGY7
155ntOhKHaPM9BUmleQjXk6acjgKNm+Cz5JlVcD7H8oeON3JuDwjWuPueGQa
4Yik4cKIu0dgfjaHSLOSWrbTSB384uC/XMq0a98w0CIUezyIocAUsNmoqviy
trHaQtulzFUGfmuIxg0LvjpD5ZoRIJwa5lNwHdKPBVC5vJgiqY10Vae5nmKb
ZJ0WvwgVwqx15MfvcPxzpd4IUlQ7kbm7VicxYeAHEAN3yNjeg1e54e5MY+NO
gjwNNz+i43x6nHP7/dfrP7UNbHKvjnxZJ9hETvUH1eCz32ouQLHr5QY+TgSM
WzO6xdwYFC+l0UDZJOEbsxmXVCrlWas4E86qHazUn1o8K94+NRYOwG9y5x5A
BbzG1AfkVxjNCsDAj0Ckj8orQlaW7CiYgmM1JHFSB9f9wSTYkTJvR799zxWE
JWh2FWiDQvq436fLe9R21rG/A55B01lAm4QgFoEho1uyUtU/7Qa2llO8BC6N
lMPXmqY3MjSCpBSicY/iZFBU/jSOGtM2LmzTs6KK2sppLLiSwpy0uIsQU3UB
jnvSvs25v056ZsI5DbkiMa3vQqMw56mz6wGhEq5qe2oWWUuNNu5f+7SUqGFx
WiGTJw8Kac2z/xPmmwZbZtjNGBMcPtOr1riFl4xdwT0e2NGKthxolmZL+7KO
EchJHujGMVxqHtbioiZdCeGyAqFDYixZ36VILDTyyR/CQvY3JkhXI7rRPYiD
fFruwVF2+dzTFlOuBTXiIsd/h0iURYeWu4F5S9vluMzhmFisewH1KnqtdtAu
3PkeZ/ZLq11vmGCTiiMDIaYeK9F8W202ftDcox1ibLZuqQJdD1hURNiw6clV
b1g1BkImhj+vlrO4htnSbT4/XTv9QSPBLOE8j9d+/N5lxwHRdYVelEenzyrN
sb/X6zU4DcQDDpmiJhl15t8ecS7y6ux/1pRTIT0d8bCVh3wlTK4QMPs3xdIE
qtQQVhIMe1erwaNkG6e30RJzOabbMxJV2ZasmMP9O2CzMSAQdsVxheDHdUti
+YxJ7gYmMotGKxcIRH+u6MRsxw0BmZUOIpA8ebSdQbKuTbsObpTgaQs4dpBL
QT71iDpqACY8NxzF4AcnYI+xGkNHsVc0Ms4tyUAGvFE+x6KHXErQ7RuQYgxl
GGb2lhnN6KwtoC+KvQPituEB1Z62keB925OIEMkZkw6GXYI3Fvf/UtIIAnMV
J0LUBhFraZoXfWsh9BjlHIclc8CDRG2isKPdR3wVN5so/spVdsO6JYuRA8kN
fAZfUZ7W+NG7xyRvEPYqq3sJ7lUwyRFVkB6j/TwCuWMMyyEFP8YwBeaVEjp8
WqtHiVlNULv6qnRPTJm3d2Kg8NS+HiwfA7rXZ3Fa0/ghMwxcrbvbwAuBMCg2
5gnkPGH7yu/6YhHMNQnmdKLXLfAGOMO1nF2k4DXoo/MnwVXKA3EmTMN3fS4/
mRmhXUGAJszqEFzeHsL0acvFSKm82jPZikh+8ueVg/hSyT8uso9bBMhK5yaK
8Y2m2wfodp9xXhhBL8z3GPBW/aONp1/n47tXQyfPzZnP9o37gBhc56kNPxaG
osJEXXOzlYwe/bWkukJTM9IK/t2476bGV6ys5u9dRA3Mb8BjY3oR/SuNe42E
8LGb2X8fyCQuqWfJKigyh36smNUE8Y80ghgpYWDquSm6XGxwBWi0eCrnR1zR
wHmjQP2EzDvUIgEuMRHpw/BqdIlCthxvYVGJxvWNZFVV1vq4mVSX0XltRmy3
xQStm9bP6iuOq216+xwX43YAm7o7FMqOVTBUS2wZ/ELxkoAQMT3cY/9JGI/e
Eji0DSqRZd8/pe5T2NwhVpFquRXldKwph5VcsgLoYPCP1P5p/sPMlnebNOwo
z5y5NSkZzM47iCByCtkpOuwYJ08wRKK1W2u/PlVpC85MKwo5oNRLH0f/lDO0
mVND5PMW4cjNYZuIfRMhalE7qE1A9zaDEVwheKT6jL+Zyr3NSAzhucUe/ATb
uDxHMtaTp5mwl5TaKY3x34sxFr6WNiTLpacfwJHO6CPmpA458/1ObqgPcvN4
cmM9YJSbjGrUWDY3B/V+rBU3Aq3wR0mUv7KtyT3e1TbxJ/EoQSdAKC7DUWfa
ESleP+hwxm0zppJQ/b7SGJ557CKSf6QrQ/ytaAKpf8la4LeEP3kTvnrQWlAV
C3gcOGpO/7SzMJ+AmnmDxZSzl2ixTWtcnlw5fffMpd64n+Io++MxnyO49crw
D7SU5M1hMMb4lYkPkfxrIlpKJvV2i3Eg2A96NsAAvb8tgXthtgEV9+YJxVX/
qaAvntz8RUyPoOeUvYqliJMuD3OYqq2BBrQkKLHsdzo3sF9wzHHarz/pjhLX
xoDRfSe+eQQhFathx1k74/jqvFtRbPHcCTjSLBahHEsrbCu+wJuJW0OYFC+x
PeEy2j2u4vmkVUQ9cTyutZyeF+wQj7eNx5hh8y7LfSNqvHSX3L+YbqTxyazN
Og5uuL64NwmR8IZ6yPEhxZ0AJeFJaMN4JMsc3bly5SVDvBySJOEKz043si+u
S437u5MHqoj+lxVlXi45032aDidRiMjUlsTqjR60UU5hnwzEfH4PiF39cMbE
iV61zglBKg+mzShyt3PNIO3YAjDWR+nXEuEOTFiKxh4jXanKlIiVCaztsdz5
72/sKET/r0EKmB/+LOjyK7tDf6UiE7DGvQnwqulcyl2lhMvETz/LjqB2Gva+
jYXnPDMlf6Qzx9xQglvKLsp9nhQppzCYy3jfdxD+saRvU0hz9h/oz7oWg9OT
uw3FVW7L8/vK8jBjCSq2K2bfys4XC0CBAUR3Wpfwq0tAfde9IH9M9czE/MqX
cN6SN5AWeZxSB85aeSzLjKfFtjklLZepNqZQKur5BqKfEgSC8EkZPus8PoMI
w2hTd5obvpH6DUjuliF15zPdbZdU8Um2BC3hrnA56AXmiGXQMEb/D8mQF/C4
8Kk9EwbvAScH1whZ4OOdNeKblJuxCdh49jvV6+1BKbEssCPTa2+KK3sThyxt
RsUvGMJUB4VPgF+oVX+L62xJvgSF/qREkUE0LO+I8Gr0zaMHB2sRzM1y7R2f
VUyOeOYevmefGfEpDdIHZejSlCcOwZC4Dbf5p4/VY0mfxQ3EgQkGHyt3rZPQ
XwZ3u8vfbiFyFUSmhFxaqtsvq8aWwsduXTIgNTdYE8NLFk7ijhbjM2L0mYO9
N6vS/ckHCd5nuDL+eGPMDCYscGOp7wXF3hjbd15qjP9Mnf+1Q9/PFGuGPpPf
3udN8bFJVDvSuZ4sCHnuvtI5gM4o0VN+5EVjRTxVw7+ajrAui40qN6CoOJju
HRddR7r2mSeYzwmPlqM+8NSTGNOQOVWrRbFLYYNQgpXP58YyBztW5dvw0Ktr
A3h6SVyWxEQXwZs4xltf8gYYM9iAR1zX7N1rHyP4yKIMtAx37X8JIDw6uLW1
PUJkcZTW8K7NYqG0x6BtYD5OQGcoqXqehdRMx2tEYUKKAqHn1uRlg98fHYD2
tGTBreiVNjr8DAWWd8EozPtUnSD/AMwqPIm7FF9DR459bNEHNlkcOVhaH2Bn
ZyAUCpUfjX/0pROWNURvZeb6zZwwoi7wOhU70UGZffYXwA1hnn7Pk1Jb2ShP
Uc/sWVl2tNIF+UnUmyZV5a1XMvrTrg+vWIWz54vAvKgzgOH+QK27Q7cNKQoa
t/kU9obkeIvJlCoDRnYVorr7AlHpDhVBaBy5VBKlwF8ml62IpNcAnTd508Om
VYDW0FjaA7exsB482cDggcWG0oEDA/oF68UcfYwnUn/iL1mHxOhqjx0yr6Ot
xfIALYC3s17xR1OlBPiwMQpG08JlqQWFRbk2BOvNUjCKzcwaArbf6xL+Pnc9
KhZwa9A34yx81tIR3FjgLk6N3is5m+qqzotc80bCHjD6fVR3I2vLE6E75kJk
IjRgTM92FFIALf80FFitukHkZqPyI6/v7thYnPDdHpiQUCjikaiVcT3+v6tW
ff4Qt3PG/78VuQz7k82cZsjkYSjYF5M5U0OSv6oAe9TJbHIpnYxePmSQYikz
UUXzumrMO2LcSl/wYCF04zAXcREcwERaYffyIy/Ib/gvPunFevk9EaG4tbpH
Ujs8/IoeN75u9lqnkeRS4P7LD8S9Vkvgf9ROktcMG34jJB3l9ojxNib7L/Bz
vsKfeFPwobOX6EMwOZKXfddlj3mkAbvNGR35Gz5PVviGcgOJM233Eq5MQkMC
g4U9ZX/b7raMnn5W/c1WVSZs39KQ/QtCPE/tRamXOtxmwFpIpkk2HRPs1egn
tf4FMng9TntuTJANWDJX3T1auQnDynF18L7L6XqXAJn+KszyFbmR2GjNcwWo
v2vdLJwAB7qQkREWIXXEtdTkqOBZ3Sm7e9YjN2z7xeksuXiA6Yj+ceHYvbLw
x653Ol4YI4CwRLuFOYk96D54h3l+6r3SobunMn08tNKel/9yrlE8hdobYFtH
kyE2PIyS1ZVakGtiMwGHiYCd6/ksZLLhNU1uNuM62re8U0RJB1BJIO127wNC
YrRAfPXRD6Yn6YfMRx7AAszfHKOfPJAXJbVByFKvhlSOHGJhC+9GnLAW6Wu1
kbqeKl/YEGRqM0WLeVO0QMWSDRn9qwXJ3maftBAvxWhUMfpIMY82oy+pqxyv
Hp9ox5l3pSDDGeJ8I92RVTllosWtSppAlix2Z2nEWb+fRTtY8wXrDpNrVMv4
vnfRJcnsuysGoW9mvmBzObROZD65PS6H2C9gEOVDmNgloDdEQUlude5ya1Kq
PGFV9JU1/CQ4K0mZMGuWv6cWi2xId7qZL0AnT939xUWZyufgb4lO/zOoD3Uf
3TVnKIHX/rVPQqcAqTjnpEt1eFnnJtFsaAOZY8kgZtOL9v0tQgONQFRq74op
kGQ9ABk8ZNP/RL5uZk6NIsR2t3IZOIKDTetNNGA47rRtxAu72v8BBNgIbqkC
bUTHSm+UJT8T6Au59Hge8vY60yYs+2rJvnvVQrhS7EL4bAIj00FrBwB9kAUV
dS225I3tkkrTRf+YRUhivEaDgKuGmzz/Z6NopWTyufccTYADcOS2E18SzV/B
mSb2lDx5rCDZKRm3kIPsR3xC1BhsJnMQDev03nvCEf/QpaV2TXOuShBt0VUY
z0VF7nFqt9+zMUGezxUmXkaJIqfDEJX4iqL6KKCtPT68Yr0eJz3VLfPdTR5h
kkdEsv68PT+yMLMVt/L8YkQNIa8rVxzU+fL9bCBRhACcXOhBdMJAGVA1NB3X
qlFllhJW2oAUPMkK0pWygKdKuFXpiL1MNDDaKArN2axOEgnfrw4PR0G6pwZ9
/Ia9FeKShuTKTa64+4HiY14MF2XFJXvJYc+2JOIgw3b6drSx0bCaYpuzx9Nb
zQW0LIgR3ImZKLbtuTlQ4yN9orSLZqWntxaVhE7BRJ1WmhryuFpDgn/Y0CYA
g+tZcU4uo2m7QrYYQLiYhSukiEMASegw1gLX+TV/6tyg6T7LGZiFpENH1MXI
MEuzbmD23s5kouhDq8EwdDOndEWjimc1LuDAApNrAqrU7tXOpJkQHY9Iqlas
VKDjQ+41IF/oDBN4hP6YGBchiJRpd+0TwGV5U58SdkGpNDs/xi+suxNpzZ0o
ul2yZQoHWNyS4yDtpSwC3fnjIO5mUN3npc3qLqN5vBiG2yxvNyxfKKrSqZJ+
M5w57o5TCCIg7ZEmrY6xYqZnAyblqEnPG8koF5bpgQdyfIBFj8GA1KjTxjPC
wedHP3v5TeNZrSFOb3nd01urxLo5AB9DHQ6+6uJBwYp4VpysNJN801qtThyw
2eZeA/k4IHnBQRjhvFV2tit+u/7dB22JcoXxjaT1KKwNdwBQkG2/DCcQH7wg
n2Ch/7Nvt2CUQ6bl5m0gAp7V6skxypGyCEpYflNudXS/fFHWi67Zv/pm93R5
EFjv2I/NzPyWxUiacxwzpCcsrAiH6oqttA90UKf4l4A768j5SD1jWwY07/AA
P7SX3SBJqNi70utjeYxyRwB1D/8yEMKoKUkHOdfcXpX5uNsW+bAoXm2nmHan
CaTW5+ChXqjSjs3tYjGlvbDBNRCeBSlGM/5zxdCJXBiA/RJIqMDWl0szFZi+
HqUTkvIVHsCjzNw/GX2heEvG19LfkzxMOOGXNFbG8a5BfxAuHCamjO5cnfw1
kt2M9LR5GxAMzoRWgRyUr4MFnf8INY5rNN1JHLbSm/CA4X8RpmA+l8CNFfun
GfGmag/6f7wPP9WJO0h+58Hma90zSVQDgF0J8mMPjYTgRoGBUDKpgghWDvxS
JqiW/obZrufyIotgBn+PwZ6Z6fO7iojFCdXL+qrwgPdDO1du5GRueMutTkaC
wx3klrdQo7bkHw33UCQ3FYoUTasPSW5rkkIXC3lFBkIo/XIxPCOe2tZk8YBm
PAr2eIflZL2VH2EsfTuem4FgIP9xokc3lZd8jTkP9iqWvoFjY8LUsqJaFbpb
gFynAC1yacGyOJbblraE8NsPTf+Xuy1BaIZ5DGSxhcImLNyX/tqaNPY1tUMj
LEhp0dWTSwDdSXAVxGFkj0E/MifUs9YSTHfZrueB6vyMOCfgvuYIc/JjwEG+
H/7wOsHS0ZpMryAWkd4TXD4Od8LJxnPHkhON4LkGQKlCsyhfIl2SsCZI+xRL
ZUjiMQe32nLqGJPfl1tJJj/FF9f0ykrSJQEEfYP3a0wRSkFLj2az++7V2BEn
s5ai4dIklsZWz4IxSbxRB1BgrRaAdXpRYB1+L5FjKd+yGoNamA5w8sIxxNmh
O/nrgLZYqbgJ6dNv+/wC7sNQ8c9Y7moXOiduphid6TiGxzLAKAiLx7h1Zn2D
TktSut9QbigUdF5e2YHA+5KEijk2lvDMChY10m+u9Ns3q9xZPzKCXgW2sIJi
o5sk4WpkjujVy+e8eTrU790Zo/L79uB2CKlf2PWj81zDHjF8x7td0aQ9dpXl
z7WD3DDmHsVcXPFR0kiFRKXiDKjLVrpYwv92e9Zi0eJi2akHivsKFgaeejEC
cxJv3Rzu7g1Ijddine5RGcZbemtujdH3wQ10rFYDsjAolMc16FUC31loWYtL
OcL6HuDu7/ti9qd5/gSQosTfq4wDychY8bKBzg7o7goT11NKZquHeWhaT+Zf
NDWSnZg23s5ALcOXRTbJ6bJjCQNBKWZal+fRIbBRL7hlPoCUciHfOqnvCwDT
r6RxDebMDKxqS2PtrdI4WrUPISIN1ZCgnviE9qkQiTbtgNoT926Vi1gVkC7+
wNjkUWOY0yz+fwAkcx2txzGHxUgsPKv9BzdsRYpYHEgaHXDcw1GxDvpEk/yN
6qW6BPuSnYq6/bSFMt9P7rmHLYvHqdXXfYvzenyAOfdlqyI6qUmhv6NN3Z0Q
Mi70KzYOX05+W2++QI2EvwbPRPaKLFA30Cj4alhnTbADF0ln96R62z1/z1/R
wSqO+X3QqWZfNiV9iS0qTQPDp01woSG1Y8NKn00WtwBnItmDMJrqNMV6JAzd
kYC6xI5AeVId5u1a9TY2u2jYctwH8VmVO0n2l4Wi6AuDKV3MxJHSFdG6DCED
xO6QhepvQXOlvAzUesyqNnhXes+wMDd8ihnsxPIQSf2TN4rqBG2no/2yFXja
EA4MomjrVFHPRudacztkQ+wICP5W2gJ5LuwDExZ037f9L93CjllxlZKxmYlg
WE2Ny+0IHh2UcYLNZmnRVt2BA1usfHBF4I7YodalfIWV7/dnEqwDadHHLHpM
J72qUyaho3uiYjg5S68kvz8r+WbECqVFreFHwvuO+RxqA8RBRriAgVzLNnw5
CSngvH/rjS9teqFqXjLFz1LNcT56qx2DKSrPyz4Tg3SSJI1nntzWTzPJbZuV
91vznEsI6LxyzQoDajB2BMEFqwt8nT/X5qP91B9/oO+q90vwDMgNMig0ve+x
G/Vsb5PNLzQAWG+oWeDYoMz/cJD89E0J9NO6qHqK1D2dXXVrB4jlwZ9oEXuy
OWd7j9vGfzIyGMnxqlBbozQ2uOO7V89jSUhgprT9RDUQJJNsbQraTdjhNUgD
SawsNP3d2/vL/zH3Wz2Leg674KcEuMNr1dhFpwhRN/3KBRXPMfs7zSM2wIgW
SyJFvtwV3c1SlkXlvLDHSC2rk/j82sBWU82JFfFdjHKEXTlbuKDPSEhvMQKP
/CdbhGtcA39oDlbTv3t1uKyDbzHWH7gYuqJhy5bKJkeWXIatThsd9J8LIhWd
n24FMGd65yyYlTVOzcS3CgcoK4yc2cSxt9+QN5ko+pzEV2OllateACrwwUKk
JyWvfJpdWXegDLmqn0EyTCInqcnjrKO+wlFoHck4g90AkvPgqEvcxP0AnfQz
Zg6O+fb0mkQGLOj+f0/yCILaoIVv0625Ml0l4ptN6BaPL38RRd5VrpJj03Rv
4QYzmcEFx1DkipKCkoTbbXBdvJ3s0YaAkTlH2UDpB8NDjwgHtRgo5yFBEdMr
ivk9ZwsVfUASQSLepe7RQxIUkk6dBcU8KyfOD1Mgohtf4jKs9Nv/818+JbY3
LA4Dg5UuIeOQMAORHj9zpBSgpC8fBWuMlTX1NpoVMDyYlVLQV0yWXzuY4wvq
V7dgdmF20sr2zgHSqnYvQBbnHf1gmgevLHwoI0hsDSTHVtQ356EyPrsD6GLZ
xXZpUUuWNtGLc0UmEokRL8GcM3Gx0jCMmRY4s+zQvf+8Xkb7rZiJcz5NsA6d
80WMKyol64PgO9s8eoHYZBm691utiQCQHg9SNPCz7uHvtPfBI3zqfDSHiu++
3QwQ9G/MdBGK6jdOq2siw47/jfrhtOppfZ7dZh4x1Su4JnXuqbUTV9P6PoOi
HYcNtjV09GgCJJUHERuXH72o22uMutduobxECgywZr1BcdeTYZ5yIq3UlQt6
6dexxhi4gpDJKvBXabFTMHOXVWtSP3HoQau4Wqxr4ZfyZKW8pbXuj2tVcJrQ
1PW9JgpJdwi3OFjWEfUfopByBTNSblU/GvwTpI/W2oGzii6VvvpYLSpVeqLF
1LbnurTC6vv0MzNg0mdOQWftx+fJq/4xFdO38j80pNfNJe3YFewoSSU1tqaG
6g51HxY6eZkPIUiPt8mQZ8sigsga4FX60MBSaodT4C3BaoG5BweLIyJm/Ye9
dpYIvtwW6UfM5EoBLziXuiSR9K1KdLEuayslzi6a8TLPtFvZJxAU3VvA62l3
3FSUZCjmI5PvortWBWIMDX0xw8eYiYrbHW3myflx3Hi/rzUKym1oaRM7pk4X
GgKgeFMNBi4ymcJ96+iHO7b/RaxsNyVN6W1aDPlkFLM93qiCI//qhJyRJ4g5
rMULzKRHvTEOyIo7Ga8ZUgCrqkUdn7UJm+LXKBwVUwgdDP/CdDanZ7QaqwU6
32CiLGM/GlzLUbmS8ZvtshqI7/RTHqKntmPwrG6raIPSLvhSgS9LvvAknTgu
hrlTIf+Ou/cNOiUSb+0vRPXPuUPq5pPue6OIBYHPSyg6Lm93K60lJQN/fp1q
YzjT7ieiGrk9onjcyFbYCTo9a1lTiL9t3EcQgYoIbeKgGcv2OtExC7K1Hvpb
/TvYRurz4iR2sy/GxX+JF1ahczwTQ+bxQJ0oY6BEEsDiSiQfW+P//icGoJUb
QcZrSMrk1IkAJfMtzIm+6UPq3YBTAawfLity5MfL2A8kn/fpf+h9/yOZ5e3r
lhkUvTLb4ay+OShZNrrTKF0LQFpIet7H1mDe3DzEqVJFOkIsgfNrKDPPN1Bu
eJM54UGhHmq/gRcSgHodUdgT24uSLTRl/Xk7srnI7+GfLonnTtoadw2Q2Oyh
D5O/iMug4ryzGVC9TnH2+ON1wVF75gLrMLekP05v4P3trX4qmadxPP6nwTrm
aG72Z8DtVPXuUTE6dpEDSY2Euq440pJc8Xy/uDq5bp+i5gKO7Peyjpz0ZCZb
1d6BQonEJUzu0gP43Fc96tMsESqzg5ro7+J3siwc0SyCfplpS+Ss/9KY8yoG
hAazIkeJry/Fhv0Mo1508yl8jDB93zjFL2fOsswzNtbBXZsMO3/vZxS+zx3T
qhKFF378kzCN2GMENOYp02tTlRd4gabc+2lXq9VII8aLdGrrHVcmRmHfJW26
wMYt8IEG8k70zzZcrKhnRrg4CyoqW7SEa3o69B3j2ButZWvUHy/I8Aq4qMEW
XedtRS1zGLNM7Z5nOyugM9c5VRzdoaA28l0tyqZej6acMkKtkXWzvRuugK8d
J0u3AZ8Vh9TaD6ymUCQGNudC5tE7sm0+bTpFgb/vfYi3y3nyBwU41swAIli+
PwXWJqop7Bklkp8GGfpvD6FdkG7YL0IJBJcYM+4iyqq3sU68ALF/3ScW6uCh
wezK84f66s/yQZ951TtNivCV5dvX/iBCZiZ7j+0DtK4eSM5uZoHoKA/McSxT
geh3uBrYZ9pCFD1NsDCx+VXw1korvHdm6EKyWnrA0w8GWxx59REEj97rqtOX
HlhjSdSRLvq58x8pti2JpPOw1RTjMemsL9NwQGQ+l5l8whAfSsxo9IMDLszB
rlRYJ1utwCux6kJwJ8t/lzjJ7kksihwFOHcpPlsO1CYTesHPOLarjlqjD4NV
Kt4uHTj6ATlUsQsiQhqUoxz4+zZv/qKYTznv9lFb2vAX5yVbjCJdMBi+QcjQ
cUVYwSwcZ0o1GOY2f9iGXwgRnIzlZLhC+Nqww5zXy0ltuedPvbru3R85cEV0
4nIeGFrYKXBVKa7sIgWPQikDBCO9ANfsTYKYz+OyaI5mI6mtXFfPwN70m3Rb
qVp0GIX3w4xybd4CodcjTT5CrpWDR49U7OFcT9nTLjdlfrAYDcAYulKnGKu3
U4hjLU2vG49EpHqxBcU6ACfKC5wSWYjJ83EuQZ5MMMcT4ZyHd6fcMT60KiCb
GSpEFEz+SKlxJBur9U/6mZL7s7gnpuNolqxgG52NQt2SFIGGMIaUpA4GQOyO
EC2SCu/AcSeyF2C3Io/rw2PgEOqAea/3ZKCFiXoNHQM3R7HxxF36HU1SHXDC
4woeCQfy8X7xHOWSuS05V/tJnjYkfHlCk/UtpyzSt4L8x4GMAkRf6L4Fhv5A
1yxoOh7vtVbA2jKZwxUM08Z8ye7/C7YO4MdeI2pa47dA0jBmCvr5tSDkldvh
nWtTl+ZqIxiFgZElOIJY/PiKhRfluPVBXQZtLKIm+3rNaGSGLBu2EK8gZi57
y2zZbwryhg9U7kkCMIEIZutTBJiOFP6Hm6hmrY2jPX6gEeqFruFdWT7E4gcr
g4msNhdFpDsP6RgQnZ7lm8QilcLziddjc+Xgp7Ha46skW31K3RU/PLQJLQFR
cxuOR6zUmveYPy1CjIlZpTIFTJbm8X7hNHTuG3OGFSZKaXn8gULT7VUOyZHB
HKYO0DBKXIFraSfYmsypArtx0XwBiosdPSx3p8tLj5AP+icsVphw3XspYSph
AfkehXjkbckc178XxFXg4Ox8q+UNfRBJrZ8AVSpgCt8a+6PnOSrpmwPEscnt
M3+CZGy/mDY7pQzBmDtpfvmE4pgxoJqryWSRw+jE2tbfw0ZN5iNB6WNxRNBt
RJySp/oKz2PDsKIE+ghKyt2HQ8WsX7SO/0VTc2yZfaDEQXcsyRA+K0I2jA3W
3A889BaOtTVCf9gMTeLc8z0SH+t2E4N+R0zyr1F9PphCHQQF3bQhCy9v/Afu
F4IJClkk/xFfoOuuPVZQDJ5Q+1/SP1StijzCMpJa40sjRJTW1Gn6kCo8/RUd
LQxuJB3gvlAQvQPmuCWaPRgpxNfKtKjQZWOBNBkV0Cc9AJ3ZQnhq4CXpdWrn
mkPKKR3F8tTnqSAFLrdSwEZ752HjbTM4zUVg5ySqWo2Bny5YLtKoPH/RKtNt
79wJnbyZVY6iG+pDICm+OODvo4Q4iYIUJX+sDbJIW+2BXhS/gLOXHRtIrkw5
NMuIxex/7kuJ3NCFEcyipAB6kEL+lZIC/dqmjiRabFmg8bqvxjOhg9GFnRG0
47/3r+iuV1/w1HGyul50FDSWapX1+2xdRXmQovazWlzvk29X49OYkTDzijse
XLMouVy68LNyTZMkPi0BzqfshBG/G/nn+UU0oMTgA6PuHfj3aJaFmg5nfF7o
w9QsldxngZNhSEioR6vZey7EKjVsMurTzBFUOIsK6y+SDx+22OiJgFmT1IO2
h2oS13Kvum9htmH/COT7Ead9DguIpyRYgbNdJjxyICkFHOn57HoR+6A1JxgL
DEPinKOxAKkz1owAj8v2MoZS5UYYJeJxaejiHZ7xU6v7fiZNm6EErHV2Mzr9
QQY2+3EOZG/HYPSUWWuclihb6shQxOyCtccx5y56dtXuxaE4wGiVIDKPVf6e
WRc1dTScfv8wX1AIq3u/JkP+ub50LPrnN1e3zLyIw8aJzC9So+qXGInFTakg
o0H+xh2kW1hQDs4wYcGF15HgrrHG+0gtHE3wtT1vzWO/NwNs1X4o3H/Rkcjy
QDdiwyCQ9BHPMt7Ve1J5FKN2WNaZLFi0wVWydpQYuUSlsC+YEWrfmdyOM9Up
g+zGClDnVM6V8OnzsDHHrwz7RkCbBd64O4epdl4Pq3bH1haOQ88lcHZQBHI0
xrXxgduUhLK3PBoauIlJ6eONX2zV681DK4EKGyQxch/XyAg01W6r62xXknTS
hlCxzMy02YwiKkxh+uvSLRatTsw3WgNrzbJyFtfmK/3WE6w3iNkd8qz4WQe7
mqVHdSqotDMlU8l3x8S8lVCV0IZMjbNvNK69mJ/vGBaUK9Hy9ethVs0Gb/as
vZNdgn451Sm8QjKcBD4xGKog5OPXbyPVYJ4bW/HYueOfjLtkX6qMQuX6LjaB
kOVbE7g7tAOQftYvx+pVMzB2dGV9/z8gua2EIOeLDrO0KTwmzswKUl3lsg==

`pragma protect end_protected
