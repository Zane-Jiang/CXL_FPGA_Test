// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
sFrM/8WdCPRrqlDtD6UioJFUA6/t/3VSOIxIlDHf0AKM7JO4OlxvzzoJCjCXIh8n
A9J1HRTtiYzEqRWLYyF7sOichEN7IZ60QZmBWcKmg91xy2BQqIc6z3t+esH8Sa1z
aRbc0AwX/GZs6RqMflwoErAsLVp8gEjl3gJ/LrZi4EE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 22736 )
`pragma protect data_block
6u/6qEqESbeMKcYmTIueQsEhNuPa7BNjKDXeN6Jg5Po3+yxfch6Z2TYztj58V2U5
NBFZK9u8Chz3bX513YNaZ4QoLcmSBBNP3Hy9PXXq2Oc4j1oVFctMhLjg0fA7UK7G
gLHxcMuGjiM64VKMH+RxF+0r+KNPCjEKTVT06VOCaTx/ECeUGfDDDpOKTk3rELWx
A18wWTHTQX4vJ8BNHZevcKEGtGvfsCq7wq3EDFmqJxpSktpUdwwen/mgT27eCyCa
xpG3Rd+lCTvn+vbwXG+i4ILJP/whQwIobZMmuBmYu8oIXE9fT0wv48x9+IgUxNw5
4LQQ5iQgU6nGangUJCGtpsCU8HhJA84Vc8CB9zi1rGIg4m43ADiwnuM7qwJadlFK
rhMsNaM4WjBBGmmsGBINjEVO+AnHPuvusoGGft+eSr4RDa9kfhvKLeLsoo0Le+a6
x8SsrkrxdH7LICl0XNhIKwVRtXkYbrWiRvv6udV/npG7hKKrAt7vY0VNr3Ezw0eK
Us/+cDKcActTpO3l1og1MVZ+Sj8sd1d/lkFBS3Hw2MO/qJazBVUJ/MNZCMI4TS8X
PiJeasPsNtrFP32Zl4TvtfpvHfEZ22mAFGbAqTC443TCJOL1SdBy1lrfDOZcYMml
51fsHZZP1iRDxBx5So4/cOkA1hsAyMAM8XvyK3JwkISfmr5xXFBp5jO16zj0Ygl2
rKeZgXWjk1muQsq/35AGLoMzO+CwDijnvVnWV7z7gSx8/12tLaSRv0udhDnOlHFA
O8cqtgoAp2pj/fVJHknlqGoh59bi9Vxgj/E+7QnkpjFSnJ3RR1TTcMiT0JdSb2Qj
q1G63XycEUhvLEr50f7Fw0es6YBDaB7UoHE/0n3BO/YicgCA3Wb+h4BEpuU7Eu3Z
MXZlknfSm2rjd4Dwu1CMiDa5URbxV0Jll57VffmAdR/N6pViWYK8aXD7LzkwQFMJ
1f2UyxCKuH00uH/HnEpYp+JSgUDXSHa89r0djh9ufgEb13PYGU3UTH8jB/DceUqv
aTqpnHTG/WTLLJTMKl8WnJ5ZcHaS1A4ktZZLSIOXkq8R83BtjGZstXT0MhH/ISJj
fGasPlbav//KEmaBqPFEnnhyF4xraazhMnpAUqAFAVWpOUpcQUZBN4HU5/XGfs4+
IaSQ4axTBk5A4U4ebz4hppfm2GAFicDWlYvRd5V63Vm76OnoDgmDiGQMqSCb+KZ4
Tbd4gItMBXrE7VuOcoXfMjtAADBbImlddxmjJA+t7TsCsUqNDCVeQ6g0L5bq0oBc
4sFAbxHtfzsMqAvuuS8na50jKK9LRcDuHEuucZgo/wPKpHfpuamiUc5cnH2TL/QV
kSxtWU++V389t3LlXoIvzyDE1GRI4BUBrbpQf/vDqUJomkfcgob9HF6v96nxSMhY
vQ/7DG3P16TQv3wZWqHi6dUwYysPLzJFANh1yTOMp1tH6h6iyzCFIgIkRJc+3sQA
uQuhsn8sK/dqbEpk4jRYMNFuJa2atArwRfTkE8yB1kekt4Lj3dIJ2I1wPw9dac8J
/2FwgxUGojZtvuDXl93A3rkSsydj7nE5LQvhfhOvFidkvsmtiJ7+cNxrUpUQ7Lna
WYYbASLYLgz3NgNu5ayLDWcMtpEz1rCtETCg5wQ6Dx3P++hCyCWlAGs2mGt/h7pY
8Rd6Qa1vWb9qkeF2zTOL43+vVeLzr6EYKUOJE5ksJ4zYXe9lTotbCBp8FjFuh9C0
cOP7X37DKSz1OQ0dbspkYGKq/YCFx5q7vMieVP+fvpllEm4Co5Wb2tFtAaX5jdO0
OjBAfjHPPNmokZvfdGpMGWg/4OaMi8TIynxn7k+wVc4a4UsKXi+8nIaWHPc/ReMF
aSAflmNCqTjvEPRAmdTlOhWWdObLrp0GYIOyCqp1H3JWux8fpt8MPN++h0OQjuh4
w35dH3CJfZdnu1u2wDmgNosFjGPM3fXy0QQ6TAa16Beqtjq6xyDBHAIuvse/9nDD
MZGxC9WwnqsIhq4ofzRWQ6xw7kYN6oDbCSdwDvVECku0hnJPB3SVcaOLX9vn7WjS
MXX7Gq5pDjv4FBD2PJQ6eK3FArEKxPSbCqCfhLKcFQ1BzIDsmfvJ099qrHVk9Fh1
CnOQ5C0GHzSgWzO6aH+/8f39M4CA2o/ge1VqqgfZ0ahOs7AGzFxjC9qqR202BidQ
6GgtZDz8IIbLJUFSxkbH7P2ON97/r3TS1E/oB/5BxcvUqGgpFoNqzIr10QileyTy
zrRIKyzaOGcCPwCQDqImhwbSR1ZtEqjFia75qQnxa5AdWqor0wCCvCemB+sR+NEU
b5c7h7frSgb3TtN0oeLBCtTSew7x/IXDRrEK3NeHp89lONReqIoHtWnimWYoBcio
yDkLr6XbeyoTfAmUpjeCDF2B4gljTuLPt17LbFgl3wxtAHCBuWFLe/U33GpH3D3j
s22T83T1JSzo7pWti6yYP0HtPlGe9R5PwG7zy5xfGS/6hOSwO9uk2JotaFB6hNUr
7EbXcH6Uan2SMVwYGt+reQOQ6QrubPOTurY4yyDEURLjwjaKzNMlh5HF5K7/PLS7
VhfzBLmblOevMyioJRlYdAPS6AqYHfyboIC+P25eXfM/9EZALtrOOhJPQ7/F5RRY
xrBiUajIVFaSUKkcFBEXgiwC8xfl2LgRjADSsix5Mwq83FwXdoBsYQxrgG3XKKZt
7sPhJKqx40ohSd1W2z+v7Se91QMO5l5HR8rKmqyL0frjshWhWyQfgc5ydoszcL+v
kOjbk6BZ+wEVjVWtT2JA+i0gLOwQ53/12dq+sAFPqUUCjMDRlHs9FPOv+owqGki1
KzAMeJWYilJ7MIEtxHRvPGjrdQedyjRrXuoQ16qKOIAujU0hJvtirZBeBadmFgAU
WtEH/nPtGWym15FVj7+0r5d+xu/Aq4xEHd2A+Mnae8qnNafhbhxxScRDRFSNqOZG
izB9/DkFtvryuMjOPZS74Jyb2Ir8qCiWmueFUQ1DIrFRtFqliDCNz1M8QDkG2k44
5AhVxpQ09VJLC//9vXkuMoiH7LXFU9MknIuxmUbc4AjJXkvUbBJvE+KSzIpbNNVr
1slMTHRfDqymXQ+/qzxolz5YVK5ixEhuH/iDOGOgWvz4UcQfi9ekucVg30O3YYFf
mrzfuMzzr2sRCKuG3Q115JacQT8hprx/lSghO02Wg/YTtGOi/bG3uiTTf+P9gOUt
hMI4X6D2NHeqrhQG4jELcRRtHU9UFpj/7DKB3kTeXXSe6bvJFPV7uDxXRrmjWP4G
g3Z2vbGYk40EIlRwxbBuNf0BXlKRbnaollqSssHs8zQVRsaoTPdPuTVRe49omrYy
gBD6Msz9+Qhu6lEuccNSKCAb/EMXSd31OHNhEZZxxmSRelshfafBbL8nP5F/5Sba
YpIUALQuu2fNB2zA0Bn4UnPU+d4PVigEnQ3IBZ4o7yMgmo0tFQECROWYMk2xt+xv
eu/yk5+NawGjOD/YdKEyNHE47ccSJ21qI6MnvZt4DowAKP5z4qIg8R5u+QUPaqoi
JMRpGQi9xSeEOAFODXc8eu4RlKOIog3d2IqC16SOMm9m0QsIBChDuZv+W/GJ9gpO
euvr1rckeT11ytyXLwnDwVYd0e2BVJL2gd1msGssNqYZSmkO1xs7Pg7sl+IwEP2I
rwdmYy9Tq3yOSvnex7X1Sulz1nZYszI2LF1Cs+Yp7UpuVWpmVNAA15hFnNAAN3mY
cZP9YaKXnl1rYbjjq5K1cXdI8O2lLpbOu3ethFFRG+JgUmUMCFH0ANWYGjOAwDcf
7r97eA9dR/TDjNWsFpDV5aGC5vZgJVjvemqDkAFFSr11NRe9/8cSz5rpnosHHIJ+
nYfGZt0+O/UakEIcy7sFpBOCvhRSvj4kctXqkYAdxGk0vo+4pavvfGRDwgb6Guuq
jpywbb6v+iSQUDJPiwzzbGRIXF1stjOkmUQEKxQ+YcqppMpt0nopCc1YeeKGFmA8
3SlJXLEa8AFhkYhtTir7M5LGxjaKsUfaJ2OTlmxnC8GNT53dxojhCje6UG4Xjhbu
rQ7k60mSCB1Kms8dRoNxZL6ZCmlchPPEf4vVMfl+MGY1jODX1xvOu0NYHyNIbaT1
BHk8y2u0GVwn9CuYnjSSMWfLpxaVKZ+95FgTS7gJlpZrlSPEdWiQoAIWn8gjBacE
paATkHXrhiDw3EP46RWvQBAmTU8OShKlIijcWweU0BtiIQCq4BjcRilVkhMJbeXY
ABZMWt1gF7FHofJisKCZwmSEqld2KnouPhoiDJKef9TBH3/JkQgEUmiISmHk/mvx
PjIlL9DkaBNzDQH+2wBzfQCewNtYPwE7hG6blJjI0Pu119XXO4BqnkGwB7ChvP2s
JJX/5bHyCIW/jZDJpxcT9YBk2CojqOrRQPiYuGemDdxRtU/L6gvU9Wyj/BLUYK4H
zv62Sw9vyVYqsH14SQYDjHlWQx3B1B7WvoB+86tTwVVZcyR7Xa8SL43H6qj0IqEp
LEUQzsTZ7XaHprXovjAYl0lNsuS6tnPRWFvNFDG6DEzBXrY6VbLfu8oNH7eHSdu7
JJjJ9rEkhg6QBOmGks9MEYYDL6V1cFwOsZEROKMNm1WyFhKMij+OwdF7iMBK06z6
zl7P/actTgUGd+Y6VsRnT1IgWJE5ZNeFW37zss9+LQ0mM6swihyVwLe2HqVyplu0
0QLG7Rr59pMKz9sPfSfqtQIpVD+ZKClOMa18W8ngqk968vXcCWX8br/hkS98JIug
l5IynAmswqYVUQdxpo3dZgSPR555ajzu8mTjs+ymhxjK1VeN+Dx9s2/I3iRA8MK6
ArolNkwf2v1zBcFQrqa3Oj5TioB6ZT4e9TvD/3S7F0vt97rZnRU0jvKjHtAZ44UJ
h77QknDcOcDGYF1wNOLk1SGA3OgG5tecFVGLH+0yepwmjTW985XF6urgo3BpaPQn
TvGzo+DC6rwppzD7pQVlpV1c/EB9bxxITmyRhO3llzUz6F+ZL2lMLlcMcuVFAGjX
mDMNKbpraJPb85cdZr35yG4JkPB80xNqCwgljUo4ZCF5N9BI5zkVCb7lZAeC3JDJ
Xy1X+SXgcX9FWIV78zT1O9MASS/NsjghBQlBNQYy00bk1jslO+6xhnQY/EcqPU1f
mEXvsd5FW1nBWpIw2NsVYFs+mrb/hlq1ZzmNyIWXgxQKodu4UA4o81ZgdrRJs2IL
VLQh17qULkkmFPg6LEN0+th/HRRDU7jsc/OqH+nztOs86Kr2j6eIWZAEmaIpX3Tc
Jplj2hWZ/j9jaVVpE4D+NboOSgUJ8HKd4s/Nsij+lARApUT8gxV5pX6rWR01WbJN
Y9qysVx4tWYFgy39Pdh+uJYeuycCQ8U52V/JcF6WXHF+vtYB3q0ovexb3aDFnicF
bDiIIT7jjco+DbJXfF1mXqFiMWIuSgIWL8Dl4PozaAaw0Q5owXCM42Hzq13YiwzJ
+ObbSvT28g/ZToPOjQg72gNAtNXgjNUXHpWVrLjhFYXf7OFycdBof881G7lwWeth
fZth1BP4IbBkxU6hRnsC//N+2Y25YMG6XV3aoSxXhyjrevEmi2TjmCLsgRhE5iSJ
UoaVIBLqZGdEDJegDTU/3hNy5seh37Duf02AhjBjBOhJxcJnX/62o4WAqdd8dwts
XdwwUV9OJbnYzevuMr6kBRq+CrZx5sRe1DlsxBGf6qv7hahvqL6JaoqEwbAv5b/f
3Yrt+gk1v9F1xyECvpIqlqDSJsmjozDeJj1GUGFEPpb4mNEXuElPLg8gF+IbOZzC
jx3fotxRY5MUbDa2F5JU+Ap92BsMNDoAAJ1ek3ZcwqYdbfMlsrWeImiQ8xue12TH
i+x4koSkFgBIbsw4EIiJUGvkkYEWaHmVjpEfm0UMv8Mcu5/Fiz3rHnyFIXKiJHRV
oVvSGz0d5Aj8zyTuMn+/kTYgvPt8l/ZtONHW6LydnerPmaD+g0lh2vX6biZO7KkZ
frGqyzhOQ8pLlseX6PnXokBJbTxRdgzHmuSYjFBzgEtxkySEZ1FAQDnD3fuiczCX
K1l7wBvR+PhCLlGCU8XjrUZPUK8YTE7Oioz6LxHbqcqmZz5s4bURvF0hUn9DYwXm
xNjfgxMN8b/f96HNkcagu7WatAlDBfQWLRY8jZRhecF5AzanQpK9qjvrayCT5scK
7r/NxDp/o/rbzs74QMge8ykPcUNu+ILzvQHTS8HuTQhfwYj5PLd9JNW5UPxqE279
vWH7pEgsP/8T5JKotGXNs8f+zfAyz1llc2O8tCmqjbwaI4Z4vGr0pfQyrO1/w9oM
fYg9LDCvDuXmK6XhgYQW7DiyZOESxki+Q7+KNjBz5EsVlS4QKkDEqF5xDLl1p1uP
iByfYOiX10s3sIhX9jCNqYldVszi09QKT26wMmzB0C47w9FV5BTRn6PJYGp2VEk3
R9vkxLIc+c1OHQa0y1ze4U70Wp0LG5ey74QadMZgnO+5eIFIqWGT0gHk4bdxNYFU
zeNeMS7dqPPczplpJB2n0OrEKqoPMY4M/QbtT/H6XNkL1RqwsEh4q4Hevbt+h7yo
KuT7gRMlqGhr/YHctw6P5Q57ZDQYRYS+2qa8uphhRajwZTGQrCCsniCs82txNcZs
hpEDHwn8AEGegrVuIMV3SulPHu32n7S0ylrut3GVDxNewxe0wDTm/y3MdylACQiK
eah1Q4z+RteJ1j3P3XpfZQQgJ1mddLinl9nF9g7DZEj+BaZeF4EEzQ3g9EDTHTfS
P+0MigE2bbkNMm1f6/WZTN/3wxXTNm9FYq+LbmxrqatqOPQZ+OqBmK57Ajjugq9y
A/+/3NsnQSawmuplQpB0eFlC5B+oPxbbgeD8Lnph+LulsCp4WdI3Jd0FCPrqfMMh
Ok/yZkZmo6TIZDhpNVeHxiaZY5E6NTGiH+AQuR4TaOfIZKsv8WqESpfEHcjAEzC+
GmvAIBKJkjIqtEyz359FWawfXMKk8oS/h/TmJUuH9FPTWb1aaxF6/vhZ0USO8A+A
RhKztfImFBp4lCCTY4mKptD5ven/gcZS/9UZvBqmA0hKfHCR9qVvRIM86mi1HL9p
o3T0DjcNNqsRj9p+dzRPpbCtP7SrujD9TGB2yjRx34GpRuVv4DTwCJ/Sp7E8QqFt
B53l0O6Xgi22zBo/S3Cnt7RcBYAY4RbqcjKO9qKCG6clmeDUqLdW1pOayxTYK22C
VJ24eBa5NVCQHtMj2y9WTh1Rc7JJrFI33JfNLrBUzZMzEEbs1UVbcoD86ywAdjYQ
T6UJXPtJiqjW+EfTYeiyqX1NzCybmDgsEjLI5Eclcf+Yaio1tF4tx2MvvkDwLkkY
qy+Zfq7HxukVcQf4QjSWi+7QRY/3F6snswyrTsim7C3b4vjTyFgneH/l2QOhHMo2
mQWlQUE+/yWyK/0BqOTOtEQRiEgLCoFX5Rv3Ie6931SGh1SCMa9x2jmiP3IgEbpt
l/7jZj1/0YOeehs9qPA7GzjCRgaoYkJQKE1d+lOddcD/DgGF3E90060j7O1x6P2C
eJBjhmlOiG1P4VwNJkf5O/0x9L0lRG4Lnib4ygdl3Uc9D9iihqmMV6/OoJp9WL0H
XoVthXpDvhK0u9n1lIzgojaZrrD/7XwlsPY2KalRKowvwnjqwCIZZ8bHpfqTeaZh
wKEAXbdTxoqnEjST+UjS6c2ycoZzw7StCOMokNF2R9WF6IA9dt7MR42KbP6I+Yr7
81GmcRUfm7rMxmKeYRi9EN69YCuVXV4nyxSmAMpqGuqlaMBGnsZt9Kyl1K3B50n3
RqpSsaV/3KTrJ7AxgtlOH3E8CRHy5ZNtiCrH7A6bBifOMA6o86Z/H6/zYoh5XPrg
kDK4pGR1EGfIO7Mp5uqQ881g/O/XElUywzwr7c1kPqoOl85VPGWm9AnQofIkehfx
rBk7Anb5ZXyDGH7efEXEKlqPxi2/u8kWnUrRDs2+n5aCBM+a5sft7GB6MkEuzKbV
IAF6WwdQTLjEqqiFX9mbYFNnQu4PFD8xz9AJAaprLtbgBJC47kU46AmjsBzrEPSB
AEBfQhZTY1lKq14BeXOwYMbnnKrcM6n012kjlySOrz7v2wCpnFkw9CEUYyb6CSy0
ELZaZfLbrpA1VAoWvArm0T6SSHwmR/EDX30zUahWyXGuhzevmNAb/3YyxHgUplJL
2VDDrJ0EtaDye0FeSkBn5bUm8/1fLEuWqpvkWtVjTtcsFYSIVOlbryFHhRl9kIic
TRA4r02/hYAQ+kEUiKJGDMhaUtXXg9sqB0JbJe36njbbRieA2or6oYoWcXEnGtcb
8qI9gwBCEZ8dPZgfbMLaM2B/5g0uauGlj9PnvAfaPudf49keRXzdjIuDmFtY0IAi
C8Dc3Go/g7BoF3ah8Ev7E6blALC5n62wm4ngJPniQozSyxQ+PX528FkZ4plXcMJR
FzffT6fya9qXUnffrpAkTHQyNaMCelXHLLR2wp/cfTiMcPYA49nC2FkyNNwFvvSl
Fw+dbToqmoo2TBNI1DebTTe0BE7UCfs/OT+nvD0jxWQ/+Ih9uZvhZjf3bgzAtUZc
jfLjA43TlVsqPHEMkQD2KQrgl3jtS0NgwyokvUfBiQjVQ2+fOBmGM67tyJYdVEmZ
txu6ubSfoJKxi10aDY1d9ESt0gCBEKljAHkjMTpzW+MYrmruJTvbnadsvksXyCPj
zRvsd+Iq7Epexr+EMw6S5tNNyKZyMqpGYFErFREZCg9rxakYCJdBj66+FgXyFW8N
5OL8Yk6MVpEIznxA2VMivlDyy7GSkIt8Mt4pdJFXBgmNgydJcjBWMfr01PnnvHTe
fe8Ao0JChNKoJWr3O2KMPizCNquo25y1cOTWiYLb2mGDOi9OdB5GeZ1WIR9LfIk6
Innve78nJys7yj1dP14XCdFEo1MJxJTv8MyBQgdAsAKJpilsyO1d8dKMuflELcxQ
4aVEvSnew+lnooHA1RPisRpoZCMaBLyjSNyxZWUWZitAJFJu1QVPYDOcKKNFbq4e
OC7LOlhthN57naPGqRXsqSE9xDPtJDe2iQXTSJX2bdMaAA6kpU9M9UNiM9GrPDLk
K/omsNCZhXUfYRsc8sw78YOHAGS1YSzkBdW7F/VUYy5qPiKg9fOoJ1oipGoI38Bv
upk1UF8WojUqRGjq3IPeuxC/sijQIaKA/cr1IqDBel1j2r8TY9mzPnXLrpPOGFsz
E9gPxS5ZT0g5WLUCQzunkMAIemBUyKRTG8Wl1wKhtT6BdluOeGRWAuKu75SHoY6Z
gP3uLMAwwfo4Is47Az1woZkd8FZefHqQwMEm/hQuLjiJffCWDcqeQt1ZF5p7b5vJ
vslccPkjE45LX01g3avAnJjf9g0U4N9xOdzw9dLxethpYhdgr/j5DqikqaVBySLp
69D/tqLUidor+RnDSE8a1A3o/cHyYe8SnFFjfRmaAhxDkz4aOdl326dSk/+dfn0O
3rROxuGe9BaQkXbLDwQu5IunsAcOXnHCmJpr07xZ37qND243/uE6qOJcUfQN6bTe
SWaWSnid+SvZbhDLuDlaM+ID/vqoHF9K+l+yemxZzL9q4i/xnFmTI76B86tdj3pr
im26k7hx2HuCPYTPR5+IXk+zWn+gDPuLcZbE3ZP4JnM4BpYBrEANL5t47XG0HKU4
PhAs9VVN3KwEo4Mo0pqyhK9kEzZ9jKm2/HNN7tybt11v80ERJn77dqivlzyXKmn0
Q7wiWR78LwRimGYxdnS/3L8aGpj2Tk4J/fLZqnPKWge9plk0oFo08rGLzNZ4/iUO
5b2GZo8lXJrbUK5Mi9Xc/reC4xjXrlNpGy2iLgcVfbnldcCqr0jJO8iwXsfWafWx
hRC5xquTjNFGkIEOy5mJ047cHWyXbiYlSpMGaWJQCsmW6Vg98fp5TTYvPEQ5soia
Zk1+mF7JectmXYKyyS5yTX4wmOMNAH8LW9NCawHFd5usAKM927TX/3RK5Fdn4K/J
emzxtetUuxuOerZT5/r5piVBGTpWDCNYXEzlsUjhjXvnltHbdd0aSh9jXgDRx2Qt
8J0f6LX82mhzxUYpD0Viwtv23qHRjN7k6V+vw0SsSPDYOhqEE15Le1/355Y9T7Mn
5lI6GZLqO6gXpNmyXM+YMhCZ6/i+EO2pEaFd+4lEDtmXzTp9rAGy0RBvrmdqsfVR
ZVXyIYDOfNS3IMzzP9q6kSS4xjehZdYBkiBFdmdIfMYBUvYXv7hIUghhV7qNO92j
iR+AZgUzZjxxTAUdUIxHYOTufdyAVQWcIcLRHtfXpKSkfpuh4e2hWYYnE63yLrQq
/Hpsz9QltiX+OvlazYMxuKxM/oAPnnvllovo13bXMlfLvoyLXde+CeFiP7iX4OK0
H+I62xt7C0GTckw16IgkSS74JZ01nug/+H1OwLs1zcCtktr72tpcosZTv5xJmW5G
KzbEzSUgs913gg8ccpg0+BkS6/TH/lJwP6WGwQ3Em9LywM+xy6vwx634P4KTNtUw
DCiTaGkna9DuieFjDUEO6/ToNAWu25vLy0UhQyu5Ul97M0EnKaX7fkqbjhOx81yS
Rkikwzp/i/gbNvUzUOspM2ocHibkV9BAOiXcjvwE7o2scpgbo/gBnUiTg3OZxsA6
TRCIK6vL2Z9UMny2BMXPlLDjQom8iWk3hJN157dwT5TurFWA7bDHseWIhKLa/16T
w/gfaDQfx2Twe+GJWFS87Zt2YTwL4C1WoVu9utl9DLeVGe90g/vSa7xOnmNpBXxv
04exS6VClyYDhZElgfwXL+j8PyrDbborkstF+3Fox6rrD4phyLhuuSpUfhDbDp1W
so4ruvVPD4CjiXakSK2COIuLPfUPRewyDiKPiTXF2oyKZ00Yh8DXP4te9+cpCqsB
//faUtzOccVz1xo6nI2zbNSApB9/iXNzYoiN4mnsN7q9wdJUiKqswmUnsmtku5l2
aLKM2vC95EZKpeGjgqaRNmRFyuOJABcJMVutUsw9MHUpxI4ZOVyARYtQl5cjW0N4
F6D8bDXfh3jxG2BmiOKci43tRIut6vNZL0zXGS3FLd8eqxsMXpj/MuN8Ubl3VCsW
kDJsUvjkaaylk+gB/sntIrxy9V2mmo3c66+9lHu5D1CTFsVbtC3mv08oNyU+8t0n
84COwi5z0BEMV2MV+TEvrUh5RLOtAXHXXHqNiUfPPeUGWlu5kf2ZgpXz54Kj4+Ce
dhd9WsVZwslE/IQPPUx+5bKEvTw8vekoAJLp5yNI08roBxM+XAkHr1FP/EafBaDo
muiIrVUH2oqxMQFwAaBReH/w8q4RHzMDjTK7Yilr9aj6s6lYYLQ7AzY0CC2esED4
qBFCVidh8jJScFcOnYriKK1slwnwIXb2de+48mPNxuqi0k2cZ7r+xfFOyKZT9kYm
dWVxta4dkynCZqLEN25gag1tnIvzDqKWGtHqNDYVXpw/w1Y8xUAFHWVwDFp73QNI
xH6xHYb688y4+ljj5QwZLLNFsx8j700lch+LWedf74hkzoL+cHVqscBwFV3gi/ia
mxG+5G+qL0i5l7UKx8VEGkqIUtZOyMW1mT5hSV2h29TPO26poYB5VHAmagsHJwck
CojPXFV3uL2jJetz9IIlR+gpOdjdGHZ+8bSQbx08Vq/yCV2Gbbfbb3Op8slRkEW3
Q/M1liO0DvUhNRAf+Mi6mNCcADkVzdNTQ0txjXSLAmQHjas6b/En+EHp03R6XNOa
K05u+zxbUqlL41lNNFTMY0KeVQv12rn9tpkz7lQp0ro3Lpkb6DpJ29NR3ZdAcFu6
T40U7XpjMhoHJowshjR2rwqoeidWqPXGhBYl/DtgdH77tUCnhdze6z4g7ZuV6K97
nCKqhXpAOXXK9couEo020g2df/gFwQrpvfVvpoUPgYkdo0+JQtGDQEOP7ZUH3m6w
fW+AkcjiGoOViUzN1GGAOves8jOovgB94YIEF1gP00OGznvKQcU3T5X/1U6iu07r
6/zEVFx2UE9U4GZ5Fl9lOpnqoyUsExFkawZcoh0y6StRRjV5JWoCNHpH7+JcC0wJ
ha5fwj5qT9E4f4FE5LSjsufzTPsMHrDX1vvR/d/LQoNDQ3zzNfh7QqM7jfC8TmUu
Vh/H3RlmP3/aZz5Aw3F6EPPByUsTjuHe/7pYKZkBT9DwS/aW52uDZSucpSvXcJWL
KYOXdUUYsVMfzbJXaokSyf/7bTSMZKMau3QXuV9xjwGZQJGThQNpvtIZTw510DvX
SiNEgV34eypeDV65r9QSS9Waf3n3S7jAsbV2jiEmEsFPWnMZHG+QjYzhe9e4jFhF
wkvOCtNsvXTlDJAnk427w85oITB9wGHU9yAvN8EDY+h0Iv1Shzwzzf+OJjwM2ltL
mYp+GyFhIiCS6yXrxQpXpKvOcTGBycmxZ6lQUhTe30FTVZDyvcybsb5RVnU4gczA
GR7VDPgLtGDO3BV+C8X2FIAhw0L2WHHI8UINqaYzKYoDmHYRnnbUS105wGhI9iPB
ENbrzCRQZmyoXEmWjgTJ58fug4bXTcCg+MkWJZsYjUE39CMKFeTDT8SNRjW4Sf9f
d78Q/9pPGYBmaflrK7WMu6Ef9mB4g60Gr6q1B09DUdLMhwjFODm5NxyR7LHqOF4I
uw1XO3XxYr3XugRSgIsU/OuDVjxa9//kayNaIJKrVC1MhBcgDEivzJ5YSQeYHFsZ
EYQ2U2gcTuEVSAyEk4JxIDtr+aK6m+tgrNUUfoUkN62sSOtIuP5T3OMQJF+oYH1L
BU3qEDRNuQN7FZDJq/f9KB7Df4ELth/qtTXGzk/tBcyUkFqhIg6wY9FwgtUmrAmQ
sJNSsR/TBBs6zkGGJ8aj0RK9Jp1fam+PTzk9HqQUrCaIPdHFjZ+zVsKRel+7mAg5
6XlGHP+kxcSqlfnc70XgAkiU+u9RmkMIfAKH5bJxtKMhBaDtQSaKfZS2Y+/UnKYg
1PgvguF3W4rNOVq79XnO4byyo+Q79EYoMzbe6MTmgmYnie3SnrLPTEeiFL2oycUS
9Wkd5fc3VrelWtb27PiI1PnsDnWVZwvfLV4hbKXafEyPnMAbCn4zNiruQcbHaifI
/Dg0dK5cJ/XUj6mgXze8jhJThCD+AI2ljfsRj0kYJ9KVjuqSFLD6c+oHEh7AQsrC
m66ZQ5/VwQhlqTXZn49dQHD9f2IzabM0+SddjYkqCf8I5koxU55hwK7IovVASjva
G8hRXJ6K3A1wJuzKEVZ8YVwhReKVbb0IUQnG4qOjw9e6T6at0wxImY6xdQc+ezn9
0SRb4f7faqgmAI4ebLGOo4tYdrQmGnK5IKbBNvCst847xEjZjRV3eYrCxoF8PCCF
1mLAfKSLv2AO1CyIs2DfpjWy3kq/QJ8BBRfHF3Ty2h3wcE0a7W1anu11WrKfO1I4
dni4/39Gqecl1ZGuP2aWVpZK9hVph9BeeedHFmLKxPdpuCKYAUcbG5T8UbbdkTtR
A/B2vzfByq25ruFHBTBZ8TuUMjAVsnZnXZfrf8vjwBKdpR0N7bj2Z6ytTEVx4PfA
m+1R9AXG0fGBa72INvuj2jJYvX7iPWBqkdkRKAjtBlTF5pdGIvEw7cGWx7KqYLHN
ZVgSisLM5ZWEEiL0J8W4PHL3e26xd3qu3i3Z4070BgJcbWdi3r3QXkNhagGIsRqL
BhqLVUmPWkgoBEivkFG3v+z4V+FkdzjsmA4nW6ro43RnZDfdljXetOWUFsw5rYn7
1CxyDMb0SGi9lhpV1jYNuis7YiJc43Ftz6jQ7u1z4UZ7HPbQFh7KKGsTox/lA/zj
w+YDboArWxTbdVcG4pNSYkvsfKwMD50M1arO+ftNVjUtG0zKdLDBl/n9AiBSW/ry
Dp4Z95J316etJPOKDPYSRipTKi5j+aP+QVu/UQzuYQHfnJeo3LBkKTZy2a/PozZ1
6ZXKSFZM1iD/x0rs4BbLR53MYKMyfty9A4VzgQNab+4h1bEwDhGDwYU6Q7EoCFHV
wk9dmWaX0y2I+a9B/DqHwMaxF/YEZmY/D6+oxNJaPFaN/8RQ8RSliG82RT3fkTjS
I25ackJyXEcrWF7i6prdyCAPeWZYkr/zT/YjJXLZm3l9NzSIqzEqH3THqG//sS/M
xu1DGg4CAgPOaATNRaLeWovO9XYdY99j3K005EishXNvEPvp/5Pw7Cd7b6IbKhgN
1kV6tAemlAbbUfwF2e3fTqmp1gl0EV8+dYEWh4bu6guK+a8RKYD0tIz2S1IVBGPh
mLjMj8+4/R9mOBifvJ7gFFnFn9Gs4AUfYsRzen6af30tXLTu8VnxteXerTf4dCTW
7Pdr0DmF6B5rd1ZbUpGLM91wY3oMz6gzRhUPLHtbZupCFDdCmGrdLGqH+derbGk6
dQ94hBrhsVONY1SCRnwUVKlBxCkX0DmALUZkhcygAE/W+sb70uJORCk3H0FKmUvN
UP784gRrJaG7cn0UBZsqf7f4IJJQcKODWHouftXj8SC8+RPLsdpjSwDRHHrJPDt7
fExwsfPT6/bl+G3efQde2YbIma7FW4iR/jerg442l/BB/NqR32BvfV7OWo4JJe2Y
aSlS9P4dfnOhdqUYkMwhh8Sdox5+g0ys7UuoJGio8OXOTPeP261xbJg8+kE+BCmx
lb1e1mOVHMKG3v+ZcCbqT4p9xFpbGXUXyRQuDZegP8uREFnXcHK7CM2HOK4iHUmm
xx89h2nirTeZ+V9hCYRCaAhn8oRtgsL2SoFjDWRmqx9N/MA0lxC0rmK3LIaD6RV/
oD25yI+uRhxaFafdZ/7fQEPd1vlSVHMpPNnX/Pxrm+wRbwJSrLiyDJ53ptSExYWh
Vy3KycMfhy0AiGH1Bax8CKGO21VwwpBN2gOQsC0HozcK/QvtnJbChwclVJF6A4UR
gqqWHvF5ntiysEQycZZ/SNdfzREt+u4/SCEign3ub/7AmH06Z21AOK7hSF5DJv3U
RL3ztsBKJzwg2tI5UfTxIUZEXAc/K/GrpMQk39BYRdwyGONzWTqxbcNNZqoneqzu
i2EipdbDZ2XT4IqjFC/7b6cYNtOvLGrFrqNhVSSjWRi0d9ehPvIWFJi+3dURoRQR
PC3O6VSVKYua/iCFhU4e8DdNTLT1GeYGWgVmpHRQGKalOkcJhfBty1Pzdjooc29e
g/HQuafTztG1HqS7UkcuMlGhwtL/UHnzodMUSVzopeUonTnvDCuMjQ03ljNtxNkS
rhTi7mzV9tg9VD8HLl9S5JUFHsQLkCySIWByf+pxN6kjhn70DPm78/LFing2IOXp
Xm8T5IkWrKrtO7ybTCz+qZjr79ucJRfvM+heX27QG5RYVa0E1Qvi0VWRyFBsLny+
Q1cRaf8JUZjjdw+/6uObW3CPCyf7dkueBvpi2GTq3sAD3y0Q/JSOt3Yq5CyOb5Ly
Zm+6iplL1y0OIDoC4NXS6CSP1+7j0zoVXfWHx3oiKdyGqvaG+KY7MoQPTyR03/jh
RCjd6qYbxSSYgDI88w0YnV0NjISEfM+0bIU94aaBJ2NGvHSBd+BDGQzeSXfxqv4X
V2EmOeNnzJFq4cCn8KUm/khBG6sDao/AHCxymViSxhhIWPLn+z01+c0em2qDI45q
T3Z77KvgPbXhuHYtbGqHotyqxEdtrTm9RXcmLcX/98ANgAqCPX4uZ6CC66ZyD17R
jfJGTImo0r1b62EqRPlMB0DcznXGLB8nMTuI8WGVCPBbn4h7PLsh2Gq6ogRlhRg0
BtCxG9DbDl7vOlriEbDRmo0QGFadAbdQENxYeedMcE2MKjJIarAmWQkYZo0RYsp+
A3bNgIvXQ4zOXhWKLaS+4hUGoyO08qXbxXEsKHDMxAGwJovK4MQnNmwpU0mbpmV7
DeG2Z8Kxs9bWlQKSMe0JwZRA+24fyVHW/ykatPhHwJcA21A05mWYq64XphGsYuCh
Vfy+5KiruGIqKWITwqjXncc2nF/VH3dlGWnCco16acMJUyZj3M1qdW+dj2Noecm3
5hqKp9TP4rTOeXM/Uwwj19x3i4GptBDgDF+bWFe40KfA0SFoRepUvcDiMcJjaEFL
m2a5oo2++WeKXFRLoMeWaUxpo1WNkXbBkiN6yWWESvajGxcQOVausM+5Mb3lZEy5
E0UU5FkEUQre+iu9tO6c2ODXFZWK8ylBQW/S6+xUlNGnS5bQYnmEXyOheK43Xp1W
WVPv+He8woYElInH39ybtnI9DrveIOCzjswifDKYeg66uWLxDHxvxuQCpTa5A3ur
tkrKiHWiAoWrJD2hC1MUC+jPXOIMNppE28ABQaPhVAT1/S/3PSQ90/iVtDS9WFgB
5PN2w3xRdh+z5/6AXtVMwVBbjbP3leWqwuT7TEVXz9bcp5sZ420vk8T2eTlfBKNn
pwGrZJU3Y5J6CLuZzzUqOg42Ks7lBNYxieCOcAyDGdyc5Fae2daVkBePMirYMQab
9nCPZ8bH9db68ZjdDZv1e8gbavyd/JmGmuqzubYUm8PIuH0Hq3auk6wxoA8LBJ1y
h5i7pvVhfG9Fk79FdWBXoZmUGR7nSa1fgG9lgEIWe8gbB8URN6fy4UfmDB/PUxL2
REAC2Rtc1v6Jxj6ISjJ7PkMlFwNFrZCsKe5/DYZ1WRhkr0RR1NdlJYYGv+bBKCDa
HFnYLRSc5Bk3C7mwEzsyFtMttseR6V1ujlMK62wj4gamkJ3sVw1qmGlx13JN4SE1
AsG1bEGtPdxQpsAWKWJPTu1jfRuthbmwWTBJw/ltsY3tq+AE5oQYrX/enb3qYLG/
BC7m9zWcgDpuiZ6MYjGExXyneiNmwPb+dvZZd2154zwCr5G2pkCO+BBTUDb3QYYp
gsQ5TjN2yrOyDfZxlrsoj4Y/LbkwKJJUEL+Ys2djatHyVHHiPExoquj0j8LRrH4J
azEGCgfbQGGQdZKw0KE3G5PRgt+ZPlsg/Z4UOdYog2DtCP+xaB9CrcZLh8vprzqe
EvPSU5JRolhfNc791BS/I2L+os2ngwzxwTiXkeDra4kaERiMMh7pQnwm6mHC/ypo
7BJa5z5f+h6L8VhmOqtFL+IkOqMLAtGQDT5sR56XKGpVdXS0s/DaefkN14hp5te7
SAMseiOM+yNTnCXw3pZS90c/PZiGT59yDuorbKCCaNlVJUQtXPgiGYaB+hdI1mDi
uy74PlQ0qCOXT29d7PU7P/LtbuJaDd4rPJZC5Vj2qL8qDQLS6xDzGlAnU6VrAvaf
RcWoYduWLPEoNMLVJQBLgPNzbTbiHQPI0K2CLjSSHMInkkuP77CZYIpA76KoRd3l
S6Iv40vBo5UYEU8o2uIZzWIKWfMi/PRJEVJUsoETbyKWUwHM2y0LSNZVmexXxGST
BGA648VRHEs42gw+U51HutRU03E48gP0mIlh7ugykcASAF3Kz0lMvMRad7TwdU6n
qBdcxOV1e3iU0mFEsLDczUTquZxdLXxeVhnP53cD+6z3lbDy6h0ptFwR/0pXSF2q
jkuAL5vKVlP6oVUD6QhqH9OKjwZRDrXZMy6Juu0+L2yYhfnkXYZXCbk0xWmbQdZe
crb+F1R8HXxI8qCYKtYs0uZZAFITKMiVydw6D/fPh7V4oY/tttY92rmSJvSgzrbE
378mYpPoZTOWSHi6oIOrRje5C5muBWDOk2/Z5N+YatMS8nG+AukTkq2aGzxXaWHa
N7IGJHfHTXpmC8xl3PloTDoM0xOCm1TiWIfArY0rYKQWlxKF8n9UDMuLYQeeSRGJ
f/+ouMHlWCLyvU3jHuUCfZwd3wgcb8mt99TN+BPErsUrlug1Chdm4ucz19VUh9hQ
6RSrngMisubusJbqdbE/dbj8zryJyEZfqhpy6eb3ZYdmwY41Q/mPqKgIRT3s7l9f
0GYgdGPPtj0Y/SpnZTyK+iDisX/S/5Kn/UErKPTZeTkIZnicAV2md8vfMLgEbGpI
irzsW5pmHa91svnoX5Oki/gwb68L5yKdeSppdVNIooCLM+QdGkoJawKZvHB+jaOe
4LC+ESHEfAaVY93SQYKq+WarLMBu0+5jYZfE3fG7FJEs/9EN9D4i4TYDzpbT1mPQ
FGEL+pQfK87MMHaBwC53lFdej1X/48FdugCD0EkRgBxBxxBs2ZBpCrRVZp69x+3Q
kjSaZPkoCkmwsz12k5Jw8S36h+oBg+FyPRELlH+zJHc0Mzf0fnQJznplf2Ipn6N+
mcozKOnsEJAAo0u1yeFkJkF1OzGZoN5SjL0VS4X2+605hdVJkWJHOnJ6PbBQaezW
PYxRvjZ1QSv0WLW+pcQKB/5D5Wvff9R5fX6n8moPduSwZsl7BpqS/MSxYA9J6c6d
C7augvTrqplGRwb8uV3MJZRDkCTEiGTobLNw+fn/kA4igT8nJug1x3CPdnVkBknu
cVKmSDcnV2dnF0AnAOyqi4BpjkeB9rd3UEUNDWgsNW1OCSqAIMTmvtEgGyhGatuM
XJFmqezxKt4IPWIpRzVOLsrBaKBqYUX0+uDgrfMlYPQGYnu10cv/pcPtPUCDj+U3
IZZlLdpV4xv5XYLoi2Grgq/PwiAfDAltJmp1AFcE5DGMQnF4b5tMolZ9wEoIA7lA
mme4SfJACaPYA78J5ijPfOPK4dk9sk7qLGmkXT2tXy9o/svr8sGgNHBi/52c+yxz
e8MpgV6++fEhS341yuTLEDBRpt38YCh85ke/JGo5hvqPbIrYnRbE8yLeaCYKcMKB
XOpLaMcGQPET+0QdfcZcedFINLK+ix9wCu0WKuamDMxvok3CqeC8DGBe/QxVpQh7
fgplntl/OEbjXBe+MSxZZr9fj59Jq8s7KIBZY0j9BslQ8rOw0+Dkbd4r+B9S6IRW
3BHiP6jP1yn9pYRWmN75AwVMoCop+kC7vbH/NV3MKgFViEE99z1qbT7ZBQkpJkqz
4QsYhSSN5PzBt8keBroBKyy/V1N2NGlYB9KZhg1uktYVJZMzEvPj34veguVyrs4q
lN1fW7Jrob6YwIRp0qAYCvQfa67hKq5J+6HTwpmzM+jynCCWntDFQR6lVIZ5Y/s9
nn5KniDS7LrZObJ8j0fdH8htFqfAOKnp8uwBpHlNk5sWJ+SEUNbVsZORUBv6mB35
rB1t9Xngfk7dCl6VM2JBEVj0VzJXMQPqmA/u44dl7LAmQVJXpRCn1nCzntNV673J
V+LnlJlq+gffftky3t5XVAIhrTw3tTnRPx0nXOnymTfW+1N/uOjx5x2h+7DFYLKK
0ETNymcNcdm32fduryBszlr5kD8U7PkzSTnyWwF/fnBkeO8FDKZEdKAFjL0e5380
4iPVheAMapLstcxYcpBjKFqQ/XP+hKf/+1QA/i4EXTHLUGyDQuuSqLKORj52tsxE
N5f0iO/PJrCJnzirtsjvhCA+swYT2XJVrvnbvrj8lwqPswjavQ1ew6TBgjXDF4sQ
s5knVVm3VzlsFafK5J0AW4Ss9+4zmsajsXQEASMVuU1Br91FQhRSx8Lujlts1EhA
tTaH9M1gbJ3XBiSKM0PUzI62y1r98b48q2nXNWg2prYLRpS0bi2xzD6gCDYONdgX
19KRUL96HTXQTHaia+xd3HvjVynVHnSLdM9NxRkmJe81ohWozmbNma9GDtINRubJ
6kdhcpsateerogXSN8ruuBI/zlXvnw8wSFfNwFKOpsBZr3154eRuk7hPLxTvyvPK
Q2O0yroc2xvWwQUzi4tWfinXWZ4Kd2f3HVL9+lA2ptBjIpV87LynrmmutH/oXews
4w5HrHf0iL9zhECVRGhmi9qV2W7WHrNIzmU0mEOGiIogvElZ8mQLB8bVWL5wYCqb
Ke0dO42eKRNW3zLR0NnJ676SydHtz2JavQ1klqsBcHiacUODeNFdokpOUXXgoZIl
9Ux6UdZkmD2hKJ/zdJg6HXIv29fyIpnpd4kJFXR5wRsIg+F3U/nB/2T+MO510dBw
WYy1V+sVmO+qLOb84G7OLjkOhRvY3Wll+L8nRMHQy96Ua5SK+2PZp9HGtssEIKPC
6PuBUd55/Jizuv3g+v1nd7g6mfNLIq36X4khq4hPBgtwUyTm/jvQzEEExofSbq1n
vqw6hPH6B2foah1XOUXHSYEAT/axDN8Q8QqiiQRCFDhu4Xc2ibWhmCZkgAZ0hByI
bvliVEHDIAh8Jbk8lqrU/WrXjhOovNk1+prEzUimwKSvCA0ArvtiyF1o9jzvmNi9
gFxw5FF4Die5++X1Zhnc4QU4A6MixNS9JMIauq01+JxTS8T6jZO7vclIdlCV4jzc
Cqk4cEi8PlfRr5nKNCwoVpr1BDwdaKnKD1wateqr/+kshqbXE3lWfCjd3LZFzKVk
A2PAI+OUCThz8G+kcg2WYBRfEsgJOrOiQ6S7lNinkj/k8S5ezy91lCxNkPFo24v1
hkkJJuKWZ0DPRUnpX6dIdeYXjUQS8vFICLHOcloQTDTIeTTXlKbI3de17sf4ae7n
gP/tDfiEZHqDwItNee/hknrv/l+ZsNuR7T5/g6/ji5zJsUMGZmXB1EOwyYREaTK8
A8M2Ww7MP/jSaF5Gz7eP/8ILBqmnM/CcUniutorsPCTFfyD5c0juDaOrGdwefZ1Q
+ESCasbZ6SaPkShcu6lJownZiSAc+JI122uGZIGulc5m2zvANkjqgVq44ZMka5yC
xSAuXKXNl/j8xgbgkeP9AsktpAPCe+ozFGq9Gcxz0N8vuRU16kRO5FC38De/DuIL
M31KX06/HBZKdyfbXegbFmMab7wkavoWJlxurEgdtsHbMtIcV5zHaqWJCvqwrjvg
+rk/EEg4A6rY1GWokaO6EOaEuaFnX2HvbFhHs1fTHbqPNCdQSlb2/U9QooQyt0/b
eTpPgmqNO9wZN/cYs7nzUPpfxguOGQniM2vSpo3Da2h8kCIrJbpF138jTUCO2YaE
RQT0FhEmyJfv8jsJL4ZW28oOz2tbiY7C+dk8XFBI8gaNOGj11u2k90Utbus36m6+
TbjCjrKnarUvPVvLfh356XtFnxH+Qhy/fa6NnowkpnYFPYMU+SuSqGKfshKveRKl
jkzWY8heQQyAyzsWLSdvpiE92E7KLEdytpAhiA4gwu17HP4bIiJag5Vj82SY0Tcv
HCkb1CupL8VBrLVqI3xMpH5VIU69iiXMlQ6xvaAe86nG6YlPL0h5Ebh4X1AyCFxd
aMuciyexcDD8HH+uquojblvZwm9liA4q+ChzELsxVPhkA6ZB/gH690e1+FZHEf7O
M0SGuRWmbCEFKYvXnH27iGbLwMVXyeOR025Q6IYvyqPtRbuKX9x0b8Ta/zFEU//V
u6tbWvn8uMg/Qa+kEnFHbBlWzs0s+O28/bmvZLX4+O27C47PYD2h8nf9hh+eGE4G
hEGEiEzhuMNxyG2xOfhyRJDj4aGUCDNsg6SJ6uVJVUx7QIDvKhrLe3WhTCuajFqG
6K+kAPo5+fdDpJVRiva/AeJwMaE6ZKPHqYHao8X3Bx9VAdVvUGCiUkSuYepQqjXd
VPUmyuhgG51zq6CYv0UNIamoMqnegrUulR6lSXmUEUDO0lJ/tcfeOqG7Q9x5deBG
13Lgh7zPTw5dYtOwsfUp2nR6WPCwD1fD/4cMbQQZ8JfbB6MrNZPx62gAVpMlDx6B
90QLQ1yWWdEOl9wauqbETZDuCltW051sFQL+QpCcAlAAdG7MfIuAncGVuD+c7R9o
W2q3NqGL2GuWXL4hQcV8hIil4YLpPzfRed0PDO/p7mpVrIL9hwyIsfcj2juAUxQL
rj+/FA668P3QOxTa60x/zykb1sIR1IOmgmdmIwfyNocR0zvha/jFSK63kKCqwNWG
lARSxP6dMdF9+F+UcvTrh6QYDxcrSmS7X/YKAmDkQZjNn56hnN+nODzBz5DXVycv
tn3ucrwanB8mpmw+KYzH+BSY2sQkNiSlxgwF65pVw3MuLq/pMXyYVbKF7tpyHi53
o03Neq9pnmIHrwILHXfi41Ln4Z7lOvsoBZ74BxarFJ1FQRXmTR3jkfN4XGo56DvJ
1qSfdT8gXIREv+tk2LMLHbGDLAf3RvVfHxy3tboo5qwC0SlQ569VOY/sA+aZVWUW
ycI0L3AoGC0ccS1BvEYgpvD12sBdW65ipZv3cDy14rYRbI++H4c+9DCeu73q/fbf
L0iOld/ziuCupIa5emB1e6qZ3g4Qgf1TNLlniIEhtdudpywQNC10TYJlJc0x6MWD
CtOp3KvzwbA+eFdw9+uhpuJiizaK/MnfYk3EtUh/LJppHrMugxrB7Roe+Z4rPKE4
jywIwbO4sbBPfOmOj1SEuAaPljDw/8BBJOy6/LqALPVTAL055+rIpHc5NJ7C4081
yGp5A7s4eG3E570nQroSO8TCVxJLZhsB0NpEFDuwDGBahpVbRMvoBxB2cbtM84HK
ZG44IYT4IW6ymSjpi1q+NH8/PV0YvWfDW0/9rQcyQWTNDvv4DpV04gub7Rqst3D1
6xSsYM9N1CITSM8tJdQvZvyjbgVFQ7bWpyvEYK+n4AgfetmEIsb7hG5rvNLWcPvb
scYmqn90oUZr3yXnUhlyo3rv5YGtK8JMdPaAnZjeE2agxiHwBokXj/aabXeCZ3hU
uGVjSUxDDAs74pyvEFOFKomiaI6T+vnXGvzmgpHKkE6z/yvQVleOH/Jdhupdw1Z7
Q94QnA7B6jtbuFsTthYMV6iCSB/82bHjELydPsFDzP3Tce4gucv+1mdR8NsMFB6N
Mi60K8tXZPHerzn5G7LZxMY7ZlkHSm6IoMVy8XVSVKG59B30lKRhLHzYAhAgpUsV
lNEjuFR5/IzdEki49jsxbZFcuK17dPkrPO8DTwfa0UpoEIuw87uKrm+cWNURtO6h
SphLRpq//GFtdW2f77NKjR2EDjzRcklpZ/drMui06mTkdVuFWWW/PF9KmtLbRxZF
WGJMfc4fzfXTYuf031SUmty+SWN0FHATajnmVAlBuq9DJpNzPPKGHiZQVIBV4djI
Qtt6dhDVWLKff8T8nB0deDoyAzra9PDPDosWQmV9IaiERzz06eEIADuWBChv6DlU
JF1TT032DPrhOKhsmg9rzsyIV8SYfmbRZ2roSJwiecIxvkdGxhG9PJAHugv4TLEA
TllS9DpU1l/YCSqjisTKz0n9MVnrgz/FPE21dz2oj7gJH8D5sf18GjhCkQqQXlOL
I/uaNWsJUBPJmoOKsjAgDNfwZqkZj4z/oI1NIFS1ZegUS9WQjw4XgQCFcUqsIuhW
eMquq8dKl1Nq9XTW74Eo0OUUj3LTFKfD4voe5dIRCxad2rEL0IhGg2foOhDhECKT
29fduUVAjEDGuQohCmHnc7Z0N2aRpvsd/5Q9A50pZfZZVP8RgnJ9RUd3pMNMVH0W
v+6g+a81z9AHcfe00xRmeMclpe6oIUycglIUBg+Qwwjy3RreKZhDrfzUvaZEcVEk
YUwxjmfZpllC18QJCjhmFFiSB5tJpHxsr+1IjbkfJxC09/6kp2Oyba6nY+/sVEJC
4ply/W2YxKKTetLpMzofPUqyVHNLNxM9awdT15pZ3O2ul+Qo3ZUIpZ3ihimQYWTN
RTtPqcNey+ukIofwoXhB5SYon+Zc9rYRUK+ajR812BYh8pnOP4YxUs1u+c8a5Yqm
B+5II+s97pzHOvr2+dYSy4QJ4kgIgNcN5cp96DmU6lWbEprjaGo1tJ5evx9PPNMM
4OGtEs+3Vb5W++Q3/ErJEgAcFPMhhIey6VL3a3q5owA9WyYAQBad5Wyd3evYhW5H
isp65oPTidgLPJxRLJjavN7mzF4Yw4uonbKLAPBBZfaX0Xa/mYYIubkwOAF9HH4O
nrYgC7f/DJ3Wna1qwCnh3tvSaws8gfSs5WN4PwNXCXjrki81X1UJ+XZQtBOV/ckU
xfOTcYr1kBZUY/u8XyyFO/EkR/1q90GU25i2Efz8eOJoAod0WzToJeEphTxaQPYB
LeFwaEwNvmwOWFzF3EJCGYkL9I4xSPqlRvhE6G8oelzU/8Yod6C0MK4vOvuXJVSf
8hod0dkS23/g8gq46bBNJT0GHofnn0aUwUdpbocipX9LpJOYfvKubItu7AINIgiw
Y/QEHH5rmanFpsChnYJnOmVvSldzSUeSlvXqOUeSBS5sjedzUXxE1qLVI2fK+7+G
Ghybit8596E9S9mNjnkwa6gE3xkevPPDpeIWMeSdVNrlgkjjOqgbf+QT4ZAGlGn+
HLM7nJk0gDO+3G2smxuM9t3LuEvOEq+QdmwHE+lnqcxfna6xSr7BZ4lfJi8FLUHk
E4CU780GAjcIXqgmEobGAQasfqDE7rppa8WwsrY4o4mXONK4W5yaZHcHt52zGtdv
XvvDNAf52CueD0eUGpPrvricTWgRV9tgIWQjdR9vLLuSsJVwOsrHyrqyf919uFkJ
97ronGly6C/WNSZLzY5x98XluhpmEevnxb9FJDuSltJdB9IDDf6VpLieutGLnMCG
7qCaP14YwPvtoGXutcNl326cqg3vYyyCk8XJc+dbr30oXJisxlGtsMewg/xbAkQi
dhJMJhoYLtNVCO41lyJ29MDLbx3/1zBdn8UzJFwpsgcneP9c9YczVt3Jpd+IN++t
+SSZBtZeqYd0IseoZja/M5tcKfpAfGjBayM0OBUP4uw95utrAsw4nBK2zzY+UylL
EfTypnPVt2sJ+s8TzAPxiAb2/RGQsxRNB63x90lOBVVRTZyZJLM6U/hmPBocspnw
MOuQR6HnqgZGh+KSz4TUMOcbHU8hN+ArcvZojaPvnqC07qrlxuHBzWjZzw0XBsdz
eq3opYBX9hroAtjLpfplj/FNaVRs5PUAAOjTYGwfW0fPaCozEtuiqxoBWcMNt5/A
DFIDH0pDVXOoT/IPafUnHMkAEJPHHCp06jwv8x4mSi5C4D1TUwR3shbjiooYnngl
Xr3raMkxMB+CpeACyry4WynyZ0Db37nywogj8G8+sUL2Q++Jjv1PnZ/eIOFAcBU5
Wed5AH8DVuBgEKPQZcHceJD2w+UIqHDiFAyOLggMJWh5yoYDp1nBFYhUcFPCpHvh
n5Cbp8qbQvFHn5ve2nFxj5i36zkvvUa03PkjMNIpRc+x1vXfqog5ZbWOSYRhQ7hB
I0QX6+4q9N8PK+6aPGWWPPgpBsnYyPvftrHbRdg6QSlVdjpZWKI3b1/7r8TVkD2i
dCzVZ0vhdoUeljYurXRCl//DSprrJ55BRcbqwshqZQhke5Kyb9acBtOzBB9j7/jR
B5MPjwAz76dKUDrAGR1kyjYpnBQyi2BJJ5B4PupFTXVrYvrBPe/hGXAq0ftjHVHc
Y19IZ0i+IPmSFxoOJFP8+77Pcsq5rxapW2at09W2MgcPZ52z2fBBunYFiqyHzCSN
el+6mwcHzp12LaafHko/oDjdRa3WucG4/FHfpq3dHhrJ5F93n8l5BkTwCJrJLlhZ
4dSvlPtoWp8jrEy/4EA4DFxm7+KpRH3WGBVMbORolFxJ7hzn0Twpu2H0iDGOA3pH
MdaZo1o5QWTz3VZsHl00Rp1plWhTyCWLRhojBG9/xP+0h75wotKXWDAHHGwAUIdN
a4ZxJCwW+dmnIl0VU4Lj2vBCsC/20HF0GIqPGgMk+S0W/82BKRAYqvZPkHTDHMYA
A6CT8TiITkv83Rb6ooRvPSvJs0YxiSGEdERNSU4BCnDRVle5DfngfzopHyz+8Mc0
R1KIsI4fIfQAms0pa9K3hdaiUdVt1Ly0HyZ+GXUMR2n9i3H+PCVcif+qf1hh6pjW
1rHCu3iCnEBfluPMj7U7V88LFOXcdNlzUhQZGbDwQnlglcsjB6GuTb95LiOHmSZv
r9y/UJhv3In5S4uYWKPsnM0lM6G/L8f3jMX5z/MVFjCmAKCtrAJULO8/ukRJyxKI
dIgk4owuRu8IId1NAyuRuudFEpuMdzGtcy/N5MAJbp5jIZUqL4HDIAJ81Y0IIjdY
celOpkdZ1oO8mRTpr9jmL6gi7pAShoo0haX2y2rcoAkInFphszIo29TTnvLjh8SG
PQWIVTI1i1V15GYfZ23vkbnkun1uwUR4TU/qzgyOYeTnVzhmfE9BnZtB/D713VFM
VsHhAlsUNS9PKGKYvHcit/FBdbm7ruurM4uI4hrmHfn7aNrv4OhCFjJK32JO4Kna
9rXGLTXuIxpf1BJw7QNC7xVwqP7sLPYDwStikL+s0vEm3tIpxLJ0Qc7LgeempA9r
pn51edTjw8Oy5/SOoS87AP+2pZECMyd2ropSf9B0BNa5/Ut0OP/OObZK0dNTG0oR
ldXDEXZr8WWk2Szp2lJGuhNrnXgcZvFUvQ0DeaMHqMOXHa8HGbFTHtwAKvB4NpH1
X1j+v97K8AmZDJX2dGKC2bAH+Us8DYTSdZAIB9BP00OIeNUkmgN5azM9g+P3K80l
aHB4nwICe87I7TbkiTwuOycu0rRa0Wcm8L8gBttl0SzqztU1e/tJZFVrBlwVgFu2
edYZbq9HQ7QxuRBLUcVgjxzboOpWf1Uuo3BcqBfn2vcdGRE8bpnsO3W+2CPg23gw
z37Aw7EV2bvfOQ23vrcoz1qWLYOETPbCZxgaxOGrXAWrWhqTFgdncM2TUtEsVL/F
yb7XfIZZIGh34QmdAsV+3wGDVNYoek+19c4cxbxUlL2MWeFzR1GXufO66ivO5d/p
TPPS2VNJb+O6uRy3gahMIXPGagpIo+FoNtB6t074AxZ4IELqapAe37DbfzViiJ3s
8Q5/opQt/Za8CNFLpXxGcDtF8NMceVuulgvFbpQP7sFYX+np5950/gVy71d1fPh8
7u+fJkRd/8Q8VdSeZ/cCIWEAnxChN6+aPkXOWpkvfimD50AHTDbx/mKRIKL6wJru
wv0rdPmT+6zIC1zYF3NsC0zwgG6qiBnrMPJHM8CYgFmsAgxubneqsMuzBHmtNVC4
GbC1UUmkbPQ379fo8iSI0GfIT1EJHXtWfeukXe0aYxQmx4S95/BgAd02PDBXOnWf
cJa66wQ/uA2sw73f/ESL/2PAVfI8jbr6xS0o/xHGw1TLjLU1KrQyCDyqam/iF20A
uhPcxea7ULKBqSfyW3o/aAofd3cG+lRVtuP/WsmnZXCgLAlzwf+nz5n0Xe08Sgen
75eQEd1xKIzjMjKYpXaYwoJZACZ29sGRHAzxvAsEVz3jBRHBmJ2sq21hePM0kEsC
kpnFWMoo8gZh097A0PT9W12aOu0xDvN0ALwxrk4jTJSzYpwBsiLEQsAR/WpYBl/y
JC5kj/gM+tLqpTAFv1Gk2NzZW1imTipiR6cYfNgbGpKzVtGvTCw1SgeaO/QcXRfR
4weCkDxsFJMhjuDwwZmMk9AJ/Rub/P1G8mE/6GveUAIF3ROnSOoRY+RYaCBFreGZ
9jAwd/1PSlJmkzRnDiXH0F6Nl0xxm519zwWf8r7um2IJ/M4F1INtepy31eZWWOmN
YKvnuGeSpX8jJqctk7coVW83lY/7AfSYfQFZ1H6BxCDdB4wGcswF9JNM9mK3ndYU
0zDnjjUI4xxEBRlln4gueFQIadk+oL2kh6VuSlORqPXy1IVoJjuIbbSvt47lqvcp
Jwu3YV1qB/HSNIfP1ky5PQswHqPc31z+S4tKL2u4+vK98WS8kTnV9EfhsZi3xLp6
25fivHhRi0UwwDYwwwtF/j8lmEJq7HjnT2dbxUl26EPLV6aXqFarOU3Ys0rlaqfO
2YxApVIT7DWu0B9ngA1FzyTK05LBjGrvPD7vM5iX5gm3X55mnXjNBiKqOhQj2Bjc
vzA5vrpWoS5Osljr8lKj08wz3iMKhktlWB3BpXb39iip6AytqXArD5IraKyAQBAV
hoIuFfWLvZUrFADEuwdMHplVci5f/PvAxG2T7m2Tzsi79Nj1uGLbRORN6ffGxxyH
Q3AXZEMbaF5ccQm4wJQfcBo/bI7FqcVCrA5m2vH9OTfrNQYmltA5DPzDBE07y2N4
xfUhXPmUGD+ZXBfh4vgUYx16q2rk9rq7kead9CvF9xhslD4Te1OK2jdg2iyGcVdE
wOTkQLBmlHMJBfg/RFyIAVXmknKCcYNs3NNbP0+r0G7nRDxbY7v+uF0bNXOYqUnU
V9pvMshK2AQEYLL+2DDNReP7suxCEGLFGA6Gxlm/+p673q4nMIK9UXRJxtTBQXHe
lc8GhZpfmwgywBykss8Wtj6l7wqMH31fwp6sy1T10F7VlK+kA7iMae4ipFKPbWvy
1924XSXaKdiNfHAVR4XgdJh9dtfTe4HP+Veh4gEXmrEnbhvQARJzXSZqpbl9yIiH
a8cgIBM0wjL7NzF112OPevx5tgdfMyuDZPp5EiTsNE2G4u9oZqtJ2eT/zjs+F1Jj
bvLRz1RCe/hM94W1bSDRdkA4PjLQEd55Pc7S+8PFvBXxZpBUpVXM/CVM7i7hCfd6
n9Ae+zSn0YUMR+u9iM/n0vNrOJwuqaEbBetwBfiPLINeUqlDSU8sRumbJ9XLlXBb
CdvwlKHVN7uaBPwWqEe00S4FovfB6yeN3AhRO4ykBzCyf2TvEW/v+zTbpae+iBdf
pfRQ4X268OEx0VX/PxjQtRAVETQJ9FVMjz1PSCaflVLTCA1O5OCmnyjRAPtnydQJ
eQAOLdaHx+mByLjxDGZV2m+ofI07Td00GS3OmA3k85v6SXIOu8jSACkRtJp+WZmY
QCKHrMqYuulYaTZGHyS4OGYN895aSq8RgF1mGjBpaCshe7bOKoXc2oL+qFn1fTg+
sX61GS+wAMUsNkQMD3O8g1wVF1oXeOlEhz/SpC+imJY6atpJv/0oXbX1aINiMIcf
vGO2EI3UaIMdG9rjUUJ5xBxiAqjiJ2sgCgMu+ASlhuXXIfTm32jewIDXwYYt2Vzh
IPuKw3mI1A131SBJwFXPnMdFLjU7PTa3x75bTdk0KF6gCHoho7ERHGvseDO+30Rs
uttduRjDh6vBpV/vgI998yyZouoO6qqlUmriEM1Fm97r7xmzDuxS6xMVY6AHJ4Ms
qyM0EP8GmZtdmmNnQ5yqw3CFHLZx1p8Fwaf2BsbMvmNs/h+5jQI2ZFo1Nn3ZAOMz
vGj+FQckRWGYuT+qJbv5F5LYMBcp0JnQGNJ8ohOhmVuSB5fWbBm2sb11DqJZQtrN
MRKsA0wOfd3zZZ3jY3oRORffuqIvxr/mQ/IepZz4n+2QSgkLdcuJiE7tD+bU6kcf
laCs/wxZXQp1yK4RW6+lk3TcjX0qiE8R0ML11yCXl7RE0a4OJQuzg48ByLSeOc1L
9Cn+M4Ajuj7GqYuCu+V0SXUg3oYzggvPEXP2MQaOnKgrvbSPBgiPziZr4TFL9L/Y
Jy1lUVBk2pc8P9ENGojnC6Q3dlHSdxXFgZZicPksOJE1wT/8qEflhmtL6jT79YWZ
h4lFxbZB933wZ/wr1DP7ZGy4FLmT1dA8Dfjnj88OvkubjYO+2LeW07kXwyrB+fjF
n4IerV7BkjDI4jsXZcD/1XIczyBGYZg3utfeB1vYVH03guzR6odDAeJ5J0ekp0WK
sQVfflBacxz9r2RwSWkVF6uWATkQ4WVqKBiXn/QqjXVLyj92KSnL5lShcJ2HurQe
Jl8nshWBIjNmZFBFTUY2l+FwIFXz3ijCWyRNT4EDKfYXxzF2DDZ7jeqzc03zOA3l
fJXEdp0LZytQdqky6TB/wfe63lMAekkkG96Jhgu54t8xW+MgZ1o0BDjc/fBLM2IX
xaUNwO2U2XGrTcIFbB94Pz/K3tX184IBjBAS6X0h3T7ojHPE28dIM65VZpo4UiWh
ZLtCkH3N4rBLD+Beaiaj148Crd6/+fPaoQG9eixKUfKHn/E7NJE2BUoF+tiM0GYV
IVmOe7wW7kG0i7gtu6Ma73gUKDZUapbp3AjrYAxe8gIFvhK7ukDF7EnEficMdwCe
D7Pm4b8341goTTFzbUhVXB9wXErkXhhHXPOaPmDIPMpFlbMc5U526GWucPKUbJRP
bVAuvb37lcvGNhNCXj7YFZy0jU5Fg+9TlP2fjzOMRB8as5A7WQN/8sf4I5TMqr9g
YAM4i6hpVBFj0y0qdjC4Z3D6QQVBsjnLP+jEcqGlHc6uE1FqucqzE/acJNQfLJCp
3UHhdRJJ0rExDgObGt/diq6aTNbAVUN2v+xhrSjvqEUrZGh2ybZUhNCFf/kpj4/S
q4QjU+1yyu3cOPSPmXeLL+smKnl22Bv+2yp8Xvu74GqmAJEz4j6z3nKNGXluEq1U
+DB60pIL7BycFCQQ72VUD23rs2iXYfWrzrhpodHAY+Rg9i6Eu/l0LHQL985ueJm5
/h3qvE5kuaJ1L7NQBL4yEhkIpStZuV5wx/HOvUh06kSVt29aIP8PuUnnD7FAbPPx
nJTAla53eqAfYxhZUD34gO5GyafU/axqpI+/xgUR3vpBuweYV9d2FL/kPETPn5UB
oakUQoRx4eglX9ebIi7RCRECSCAOt0vcCVBqye9KyBHjBJH6gSAcbo2+oXSX1gsT
APwYSXSD1MjrJ58NaKl6AoYU5hwgk9ZyvLVVFZDgkp+jBE0ZpalX3Edk5kK9H5lY
yGDGqaE1Gk76iie5bWBC/RMkyVU5fUTJ6+NpwKlxQQY=

`pragma protect end_protected
