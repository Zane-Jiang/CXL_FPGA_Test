// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
86vY+VvhwI21HCa3ans9Qcdr0s4djDEZ5VKbgF8Tm2yy1EMRFf+szjIeCwyAeq3Y
rBKewmCst5ypHoNkqKwge3zK4pVGmS920phbLNi9ERu8fRevWr+qr5/vo5zFGzn8
8m90lxJynEUE3VHmdu+GQm716y9yJ56yV30eWxuq8I8lmn57KZyd1Q==
//pragma protect end_key_block
//pragma protect digest_block
FI8FLPGGPJXIldjS7vypYgBE0aQ=
//pragma protect end_digest_block
//pragma protect data_block
bWQ/VLDUkXuNMYlcEJ2AW9nmYvN+tiln2VuNdstJjkhJfNTiZlJGslCJzBzAM+Qp
3auaLCQahBqAQ82OjFVDCAyjVxgwnzccmUxn2THD78iyZky+R11AlVUO/QNdUiYf
G3Ke0vaRi13lMhr57sYUy+rsrXEqnM4G+yisOxczsz7iG6g/8ZT5R1p5S+xYT3Ds
5ExtTSEAJTw++llgfC/tVHgvtKvouumtGH+H5N+bDNR4SxVo+wK27Gylhrp2vO1s
4Jk3PmOZO/Q4BXFAho7zjJihEAMhttd1p5ahoXAjDbhvh7rdhGk7wZXJf7qeAdx5
a/cz0rEA2lWx4akypOzCZCdIEq1L2K4LAyJ3TaWEFcAF+6Ngju4Fgep1iAexi12G
GwuFZig5MrdXTGqQ78GjVfD2DTHwJs+fiDfT8bKxaZpd6Ik8V9lttyKpi7gaGJxX
NXGNW5kY3Cr5fJlBuelKTGS33wnq83NopmUANuctO0HV7twqnKhZpY3msYtpRXXt
0IROsME0Cv0uNe+I7EHgTzhmaKx0Zp5/7Qh/lnl0AZfV5n5F5xbcwPShE62nOym+
va+OCMkM3i0SQNagWG+fQnPtGHVkqL8TtXIvKA75isKcPWeE1IRJbf/rHsMOMd1t
/FK7+gvI977dTuzprNP54TdJWOOyMpMbHa7U/AMa6xYLa6XOPWeoMnKLM+0QnuSK
TcUIE29BB1BblsfZUutQRY7Q+C/23rse+hqD74vjbL2SNDYeqLQhq0AlSJB7RLIE
+x4VgYizSdKo0ljkTKY/kjgypCwYgBXLjQoidpirMMmcidO3EwOUMqWgox5bAZre
StpDlUYtoSoZ/B8PdFoEvpfB5jChpxd9TII0R4kTpQEpso0VQfll4NNuLipqW+PD
zcaugiGZ3Xp90o2z74EEHlrUaJ8HzWKE4Fzv0oSgp3FQ3mmtcjPorov6syTQNJKx
6cus17sT7ee1XS3u3ggYzx7WMMNURekRyz8lGUrcWZ4BDWI2h8udyoBFu5n0pzIz
eo0op0bgimPIMxyMa5pSFxOqvDCmUAAe83XBuWzoea8ZbO+/OHDXSe7BQx3EneMx
62PpLDIg5FD9SP2aXZviie5mcFwZkT6IFWjUWU0krFsA/77qqCguBFc6/QTTLylM
egtGxZBQ1nQXXoETVper1KCMeQD0cszVMcXvaMC3tQ1uG8E0L6xDNmUXao/i0i5I
+EqwazoupZWPVkwrY1qntRTlXKuYTmXQMkXC15LHy4givqO6gDM9Xk6bt3oYa5pK
nzeiwhAs/M3Ncyg3kCDYAvKMIRQl1csRkfJPdrtRQnGAqp0vo4ZKapKMheJFbmnf
TfxcraR1fO+bMjsTZE4RrNR4PYuuibOL+emBLkeCiN6OsOhLytNrK1mdCT5IiRON
WxttQVxG+sVi/zRzbWnrqUQCOK4eDDji5P2EKQbLnvcgCJ39KgcoanG2Q32A8iR+
AWWbF32wknTnTD/EZ/GTvL/8Aq+9S4iSaVX6hfEAmEO9JFaMbai/DfJTaqKOyh9I
OrjmqUm1PSdriFkc8Dp0xz5TvdlYSFl/sFlMfFSRWNgMO+OhmFA+7c7UAwRQONwZ
HTk5HJzoXMwUz6U4ZA21zBZKA6GHNTCzwsAgr4E81R+vTlWruZWRmKkr+p7dXBNq
RrsBkp2CsFVaXh+nyv0Ji+rXlsM3Wxolzcx6NQKfLOb/DYqH+d1XEk8T2S01JW5b
GDGL3p1XUNj1uwoy9vwxbmWnsg5NFm/OroV3gIBjftKVT2/AmOO07Yd9WjqUpqoF
HUdOrpnLH1vV2VOoF7TW/dfqKimKEo0FLG0NhRr8ivI7mMfqK6qHqEyCu7a3r7wl
SBjCCi+HdCR8+tdVc5bQ7MrmgpEa+UYcxvEwcedyl6jjT4Vs/Asw693MF9KKVx0u
gvOIgvOzXyE97cQjXeKOvb5qy49xBZluryvkxWYaNHqW5kbjV8d9c4SP/vxnRWco
sfB/PtL6nN9bQry2O/RtsVwcPCYKuCR9isdHlZurO/rfgDJx+Nwms2wcawwp/FkW
piJ8MgQDXfyVl2IorIYTEY+BZ7pVUvllux137ZRplaQRUpSgsMh//IPoM6UdoqIC
kD2gbT+apz7vfujWpqN72IRXk0IQsVj5D4iP28b6jab9PAGxcO5iDejOThZMgtuv
8brVuBf7wvqPdG1HLth5M58n23RzWaSyX9b79216H2t0Wjc749FM8ulnFR4fJIPK
zCaZUrUYuR1XW8yM++KAMI7aQfP7y5GpuKxWqVRW2QvYtbhvHMdH5JTD1KRoTese
6IWS7n3yblyUrBmuNhHgQKbD9I0pgeWpBigldoqOeFXLGms8BOHsscR4zaIKcINp
DVTQbskGUHRhmIFP5Q/BZUvUBoJPQJLnQ9JpVvoUZKqBhDuoXjGENxaY9LrvnS/3
Gis/YwSXUc6ytr/r+eqhetoYqYo+KoafaIpNTWD+1XfoRCNKLMY3JHBkyU4GHPw0
PWVzbcjqI0ZFY91IpaAvZJp9W8qkiWBXeyUrq80o1uTgk0LZS7sbAzC0ywn+L8T1
G29Sm+xWwcB8Ku0699Nfeyx5FqNgNtTl+WvokokGOTHuOSWGYxiSIK/wJXbIsWBe
t2me7X0tVR2jQd1j3ldsFGwndaTuiBABPwLAJELueAZqAz/JpcBx7s+SrvtDPivQ
Vx9DK31uZlg7JKP93tEyuFRZ81BUcGdzD5Al9Txg0Q0eKaVMNLaRY/1lNw/lTjhf
Bxzdf6dw4uqG03+QJ/rkg/YfcJaH92m8zOTJI9KVNTRKK/a2skhjeUfkfokQBsS6
HV2LvuMcn0GJQchCdwZqPpLZVC0UuyHKWgQkDcKbK0SZ7s4muJ/wWSmr5kaGewIR
fPpJ0ndFrGcELJTOFKRArgzVAGa0oX2Y9VjO7sOc2hwqeriQgoY3qjd6II+pjPDT
HuMwvEcT0xQwk592jYPySg3OCVUbgujgDBeInbUysnardBAZ3Pqz4OeJ19j0yDvG
EoNrdQbAtW6zt7X+xQ0vX0j3h7zFaw7GYI1ouF+woA7pqsKGsRDn18/wTdLuCXqx
xPFGjYIxhqeQltANxnS1Ouvilbn03+C3eo33vahaG9JjwSVgZb+11vzn/9y9LCLP
CWrl58luzRqOmMulUeNlScVP0SERUDMRd/TQYfkHvHfBlwxVIGwOmHG8QuFakazk
kTfgfL0wcGLzA210zOlDTTP2yDAU70YVsHLEnF5UzlRgN+DgvdfV/xhHEaL+HyNK
jUQ15d9vT3qd0IT7ht/n0ctaGAJbuB7WGLCAHnEqoE31GxoapZozuU0Wg3rFe8et
eDjOQW2ATTfAiJS5nFuIY9FF/cNenEf/ndwb7bv2MqbfegOjNaodRooItx41CWqO
RRRn4mKU3t94WrONhaodEFnXF+sY8sN51TDueJan8xDAMkHnaJNzJPFGrEzOk7dd
dgPGUrX0ZV6YFvvOo3FWA9rer3N5f72gyt2++MJtl3HjytPOiyEEcyZ66xRyPs21
yUPVH/t7gchzt4A87riArM/Z6G986X2I128YtOAdRYisEJS/Xw+dtYjbGohnj2vQ
JIJcnrDCMW9PxERy9nyHYVdJSBY7Ey3JP/yzkeCL08/5lbIezG78Y2nCpvcJJnBZ
Ryaj5NBlj1PipsLhcHGMyf0J51MmqxBbu2zDeKqeoieO2Yl5cXFJ8BIZQwIdBYtk
LV5JC3PonvJbpG9cTnMwrt4PFU2Y1m45hLM6/abY2Wh7MzzbiE8V+5JvtNoGHdSj
wAX+efEK32Xd8Py1Kg9Yz7AWnLgl8FpP0RMrYmZviSZzm3kpzgOhX8MbhAftP1k2
wxsCiIetLmk1gKrzV7mnnG6tmkuBsEHsySgHVN6cymZW5tOE1TIx3EAMBfJXF/+4
61tZDQO+RS1PLlE2PT8NKvOqsvQUh2/bVmDc9J+ImIf7RcgA3N4NEp8E/WymR726
2ub93mvVO9dFekl6vekDx68WgJvWqJKy+O5zbGK4WGvil7z+QjhNsf5ZHqeD2ody
ZlWctbTAyR0mFveZoTnL7Lov6fesllYxh4qeGKYsWE6mENTKvaYSGtHdlHba7NJ3
2xfWGZY8/klB5N++PWZVkUTOaZTTRvJoE+CvZY/uDstwqlbJn6PQd1xUseBK4PRs
BWVlzhAfQhXoCEDA5LlnWgmIYzrSWnKOXrA7vjxbLqriVdmfPR3Frp+lv5ptdujr
xMatYvb6mQvXhhN1Y6M3FdfGSDbqo0cJ5HMSoU7QJqBLTdPqFp54TBlPoAu1dKgG
+GnOzOnE77Zf3ukvqsDXC36vT/S1jZE9OBeInSiC4IlfYQmjklDA15H2J2BNOVHG
sAokc4YuohwVOHcuVdv6i+DSQaOSWHwkNYtuDl/LOjNnOIJMJf8Dkyg57iSM4pqA
l3AF48YxvZBRs1Aot/iKdQgDNGCAq5pdjOwwB6pCK1T1XmAqO2WE8yZsIRueeEQD
vQLJIdC/gM6KmNqXmMnyrR2cGjThObx2bpqR4teCEWtjIzPtFYlHPwx8yi+ZF/nK
9FthmIEin6UXQjwyWGxJcEVskHuUXccgipMeX4fQXoCN0DH70ioZCmjisAEKZiZY
fcjTC3nqctBF0/Bn7ItbipqUlEQQu/K3pU6FugZhTb13TavDqMV7d5YhUwjBQ63C
I9SFn1m1PLhhn3MU89nVDz9JMEI8V6PMCZqXspYWBdlBQElrFF9EyvqR6pqLeyE1
TGUm6j2dL/VCsoPkvblhpqawcBWaTMvg4wmbK9cK9G1/dWKoR9W74TrQiTu7pZ8I
49ClfMouGrtsa4kwIFN7L2DsMTJY6BqX8JFm8bM0ZCtS25HH8YrJhxnFYv4vno65
GmvfdzF3pxQ/MHKJg3t7rHE/3XU0bFmS+a8DUH0bj2hxeggSGV8Ai1wr7jmtHR3z
3cndkypzHHJhT5SqxJuWwlYZ9qYqmu6MEE41jtOmUpLe4YqcFMqAxcSolwk32VfA
XGkYhe60aq5D1ov2dYcVDl5QKPHu3+lYbERCPrgmsIxZX0fciLRJ/M8D+Kp3RD7i
hZnhJJ2UjTbumXlO9Ff/QVGoOafAxsl+ot7jqCq3TzXjbGo/XykaF4Wpk/aQdWLU
xeIwzbQrDf7OexpWVaCRvEVqNKUeO81yI/uChqzsa5R+zBnKcuansGfBokmSgOMl
+jj65uzOQzmZ5wj8ccEqAmdxDAsr+TvsSGwTQ169k6TI+WAI0CogtsxI1g5mSenB
MfrqTs3ScqwcZp6cUGBokYzUA8MHpW1yqENbrJVFkPVVt53x/MvKbyXIQhmGsB7a
P0o6QX7oWfuYeF3f6qooY45vyb3Zcrox/n0ZHJkM7QHkELx7tI3fB8NBEq1i1L9T
SROS3fB+Nxlmzd/KlVHJrELRGcVxS2HTsCu7DJY+7cy2J6zdxz1QbGloK2nnLqxA
ro31YMSsJ9Gvdb+pBlSqJBKSvryXqmZjmaQAUywiVJzytV/GZJbuOJ1EHWhD7p2i
/MUEGL0DenUkMpYYmj9PJx2SpH/2dTqYRQjeVVwnosNUeGQbNZQJs3t+HFPv7G9D
ycbZbmFMN097JmwinXGkTCSXLEsjLyML82+wN5ZuZLlvomkR6Dv4ghr9moPaBhGm
W5RxMTaPvOvdvwPVqs0+vL94jzVY7BsFhHx9IUfQuETAcnYxH1dEkgN1t3TPBo7j
DwZFJf5ovqCN8j7rhzMtsopvKR1jX5gKfEKwtV/eDwTp2BlLEPC3aHaFKGszlMhc
+Kt/GbXyLSbk4h2YN+/BL+LsizwAM+fwUDuC6sLKMqn/8ojAPktmyuQCiZ6WAqfT
Y6cigyc6ogpex+TOHi7os6cd5LZd3j+lcBLinO7+CQTUuBAmQ0Gdgfdpwibpe/oK
1c3nNVclFxdgl1jhePoxFyK34/RdI7RkyHMwoJCociEyBTRLZnNq27K/V/w4/t24
HL00JugS4VbQxbfbr1i3YeaSfrCWM4e1whbLOb1xv95abYoIroyXtWfEz6YBV57q
k8q/YEJ9f5DdnxdMFm/eYHa3Jjd4wvB+cxxUrYm7Dzjb/pePb4KkWaY76hUrFoAu
gGO7SuQDc/AAt9CNzx/VzJSrbRpxN8hTnaYK3G5C3iwQE8oHyL6Y/34Fu329dK2P
L6807MZkIqH6fSw6BsqjdHOnJmflV4+fL1o1dzcSxX1lChYoWAehfbtLM/Vhuvg4
AJcXXLeYo9ydQkXMMHe1mGLsDvNxL48dP0SOOd9zv97u1UEqZkll3r2Jfb1E2h1D
usJcpX6AQK3n++ENW+HTzpwkEVVP/VtTcbKGAkek7E8QOLeB8C9mERl89UqVi4gh
Z/0xJ26v77xGJeTaUgFRqRZ/91QhFg23lgXQ7+734feD2ImrrUjBJ2zsinCSlcLb
pE7rYIKB5Ipwv0a+dZOeGQ7tf83rmGRC8IT4gGw/n2asASkuzzMsuH770FZOzMKe
XPTMTFnBOuPS5dhyivnOCMptHa9f1UhczAINHTvBND9szVXPTCxdnpyeKy3qOwUK
ZyTTDX/UHXOijc0jXZyo9vVS7XCL7Ee4uak6OI3Pwv26CX/OH7jkAGNb3xB7ilkU
AnI6M1ci/XMnwzmx/dVA1QgjipkiIYrKjDKzGs1fUXEO/aicxPr4X9TLAPtLu4pq
ZVhjivyjydhKCTrUDxR7xAzgzuPRyb1xw+2WfBjv39y3LI5iq44+slupcOcHhYbA
Qc80hNSWjmutZztkclUFxrQX1JyptbGgV1iy2GmOkhnFFhv8T7FFqNrE0d4cwnyd
VEk2HPTJ9jWfbebEenL6RrBpv9YFLDTRlpY7JoaX34cf93hZefKe+9Pt51SEp3UA
UaWwwnIyenuPswIM/GcRY1D38qrzLYDxICwpDQo7I/Xy6sNC5I0qlPnEggtHmXXd
tgcg/HLbBLWkwconIEi/+IvZvraFey2VW38rYJ+01nuVrGTwGQg3OMdkepZGBMgX
oMj+I4b1pMw/YrPZhHt1Wa28+O+e9/daaFfdl3hQXfaxKV7tB0B5tkLwO+ZoZbqQ
3c6uKbFGNOFJfQY5Ccon5TIX1l8QXUba5rUPIupk3BdGAF/U0+1sSQSFAO9nDUyr
aGylb22MQ6LiGZ4LzVczRsfH7aE/++pPo0H1+d+tVlRN420nadP2n8bYFzRxLvkC
ATOjNxqLy+/G5IcVx7gSEptveLu24EmDQKoHQV6Msl1L+jMZMyBrnFOOPTij+E9w
ukYtRPGtWqxFQFIRd/KBm3wFQ/018lSo8Kk/dNcXcuy+pUuvmHvwS7+9tKsTdFYb
/Py9g434YRQevPid9sxBVaNr6XOnmOeQntLMk271vXOBigWx1kDBrmC8S6EqXQi3
aGHcBqvRi00OnAOujGGYp9bHQXI8eVmRYqk7mOcWEzXv2OIBofM42YGd796VfXzT
Iv1Ay8pCv/BJKzHodFZUEEl2G8GfmMaqdPnPfKksiNVmzRns2rqYIrivq7p19xMy
DYCGLvOTIdtWxgAGH3y/LjA9aktQpvPumGHmaDSmrDKR6g7r5VWCSga9LwNv0hkS
8Vr+TNe1FPtyU5LRXRIGR/DFApoLTf8XyY8dnYX/L3xlQ2X6kJ6Wqwz6ycSTmUbF
7xVBGuSRFeL6HiTLvn/kCaRmS3sqGNN+4ad/HJ9gm/IKR5P+VIq/4NKhsXuRixxe
Gd7s0SyWOjWE9aYC0uTKGb9GeRm1PJ6anGIM/m9Uw0KZDfAgYAcAR4xqtjEqQ6wD
7VwGSD7SJHEV/7nKcx17jsywD1QZ5aZupZWX64wsCdJMVivsbCpj5/UfGzrx0i8I
vqQaa8Y9JDvE31b2bzKKuZ2djDH1vbpTAJRaUVxyCxNtIoYLC4iiDop+VFleEPdX
3svuK7DgU6iO8kjsf3nbj+8/S4FMqNyQMukU0Q7iK2y3VOeyqlpENpZLe76SqWgv
/TBRHxCSytacP5UwqHnYqvM9WUtiSx4LYg5n9LIdJxzOO+mObz01m6jKBmG/asb5
L9/dxt4XeXi7pkVkbUetrahvrlUlG/pZyO8sfktd2E73jsi8w/jIcVZwngnnJ1nE
ILjGlfwvGUxWoCsylkERzmwT+61Y4HRnVVgdpsZ7Ehd+5xf5f/RqzEN+yzVjLjNL
UL4P+njH+C5n7x3gNK3gcIBwmZHlU85e4HWsdcWQylqhy2ecNdnB/MJE6PR83ooT
dPKAMlLr5VkiVpTsoTVO78uxFleS0Bp5gkue6DL6uQSEQmnZ3R8YabDsUzQN070g
aakKXMvnEDvA0l9P+GoEbKkgbe2eea3lN+15EJxNYiNna1tRPiuLGnSuVKecNGEX
+aGvVtEM84oFHFoEdgDsQLHJTBfSa+4zNK++jYf8toOeZ52mHFUFHZu4CeFWI6pZ
L/7zq+0ZhPcFmQD5nIcYrWUgvmTxVDLzr+QNvS3rBcfgsfB9WbIHDUMOjFHJ7jv1
JfNhwwPgCOH3jFU7mZC2qpmDfhzL3pEAVUvYCM1v/H3HGsUYVHi0f307omJPAe85
9D+u3qFKBtFC012F7DDwg5c9a/PymY01qruKoUDTu5se3mWOevHPFsUTurJkhcu7
7mCHPI2/s2/y81gxETyJAMmASTR/r8Q9JoDG7lQiGfYVIJb2nBS1hhWEytq1qNxe
/7y1cmctRoMWvskPt54Z/lE8skG+z4KyWfzHMrdcnobVHvWO0EpaNWidLHMiX1gR
TWE8i51QcpDzMGm+ki0mGHFUwxXn7/ivE0KbZ2pYE7H6X0ceI4I+WaUFp513fsVM
uOz97e9NfFljHwT4y32jt9e1bbv1fPedLq7lAh36lRX9ULmgzrjOituQlPw9uX2u
K7BNg06TTzeo3OwfFFmqgQXT/oxTa7WC8YUJN7bhJG2LjMjjX8Xb4Pv9YjzN/oBf
X8q6xnYEjtcoJdcWFrYUW1SbVw98s0oR+Hq06r3ktuYEh8F4HxZ41X0B97N5Cma3
a/7rg+8wsbkn/cZeFl3XKKMydiiiCRypNA++WnPEAY8+c8964HN32aVTSythcim6
V0zEasjlMiaC0vaw4dlfwZQ4JaXBinc26p6A6lI4Yz/Zhi2dBozuhMqUQG4jbM+W
IZsyI9jeDOZJZHjHtYinmLp7C8iS4UxxrGSxOp268Yv4pRzKxQ3IFpUtRUgo1CJQ
LWCSpJ+1GAFaFiKoq7j/iI1L+v5AfpvQ8DxiKIerQDUISp1981hkr2Nv5XM46U33
ayjN6smdjn+sfewVwfewu6vlTpzE6lLNrueoQZabzmERiCpax2D5pYuGjD8W8F4U
E4S/bQowBbwHBknlxhBYmQf58atfE43hZJOqQjzS4nvMapOtpp/ZFyXqW0C4onF8
75Uw/6xBZ83DP5/FYvpiOPdapMGGzOUuzhBzJzgHFonWRB9FSyn/EwfXQQ5EjTH6
EFDBxNLG/VgdwNRlSAwOYCvJnmwHwdtabMaJ/SSBeWoAbG6CQ56nUrGRsTprkZp0
vvCScinEa1pqzaZl6EaDCZ8d4Qm3ezVSasjvrAVFzJIdLASogz7WyYRXjkUO3IQl
mLb/24J/n2FrczRQrhkY//afcmS+1eEXOVtWVlIZ7jB5I6ips/uzN0a6binJsCOB
zqh9Br1AYhRfPicqIQxEia4KNqLYHvQXY9J0FqXWn8MTT+PrTpboLTbkx+Aqsjfb
5hEYleDH9mcdVmcZmUGd1xxzmzwJEygoOCl1KhZIKkE6zj6TeCA/OEm/o1Lhd6dr
BtX6azN8PAvLpYhkxdPyhdEQWMTZPhnjYRkRX1gsx4kmSdSVnDQhT8frC4LX4vxy
TmDc6xgppamcw3AG8193NEZSQD+Ei3vWzGXHrlrVM+WcDO29KzQDjYn7yeWVFItM
fAyvgi5/aCH3vIBeNl2q2DryTvWREkhCwfrE+1atXOjyQkMl0aZCEHeJ80oLEOCJ
IPKEXUml13tnjs6LraKxeNgVq+B1SHAJEIs+mPrywucfFimNTWVm6H2/nLX1dR2+
8A6ogqZbmsmU9DBwSSmR/4rPAxpyGMbMTRKKFo8b/nAtIXfr1LKH1kMl3g1iNSf+
1ZtAtX1QmcCpo6H5I1u6ukjyqIup/+rIgCgupXW6VhLOJw3Gg38RPuWJtPWCDxsJ
NIIVZTeqX/dkqZ1/8HhIBMdWEfbM0czKxzsA5H+3eIyjiLP/WD0w0XbAg3N+SvjO
yoGjd/7dFfd/IP5pAkCLYiK/V2aEwzWOiQDu8stnkbCg8AoazEvw7VZ5w5XNq4DE
sB/2QKJJgpkAZ4NSHhsdQX76BubFIA23FdgF2cDPvvbECFvDAT/xxpAcItCJIpJS
relh4iLSaJtw1LcZtammxa8+dbfEL8j2la1J6P/kCkbEko2Bd8DS882xUTutUcFZ
bgqtOH8reHRndOrZJir+m1YoxCBKH6ZdUpxTFa8hHAqsQoOGI8ihehYvKZ6RWDFW
7usS9QdetE/o/0bGfUpbF9QNSfdtFQZt/1tAdVLD3INIM0aS5TLcLDCtZocw5dnb
Wy1g3BWrAGblJ8uhm7pDlTw6/sZ00tdW4rpsj9YGVY4urnd7OTcwLOfQDV/oVEXb
52nqN4CDSjQ52dCMQhQGpmaT/20o3eOr7bo2hHH3cGE8kf5C5gYenQsBxyu57Rtk
GOmDACLysifdyDg5gS+Xl+1wJlZ+INAckoS/CwlkA10n7djEgGzFmp+6NygbXCxq
GNhtsLzPd8ExCANI/QvDPsSHw2KqlN7S9Ey32v4Crb3WQwhNz3mRkNousKprTBIT
uqH+wxsH04n4jcuOEc31ys9j/sFoMiKeDZJy4SSVHFOHuu6dZwmpZ2wP5+HNbcxe
cz2QYMWSv5PA87irx70pUCHFDtAfe6uuclxP5TSZQEXAZzpWuomYlz0WwjPWpckI
eKVXvFtC3UjMdToITCB0Mzj326KI+MmfC4ZKZcVP+/jglC5ToSINnk/kQihv/ZN5
JAnZjlvIMdImsElsTv2l+ULErYAa6gImHBhgKnApAlKFU1UfiX4tdIDAdGYvwSAy
MyWv0tKsDuq+6jjFN3m6S7CprakWQezoz5HxvtmrECvZeDL0YhetYEFHiZtIBFGF
/riJGuim1do1S4ftTL4V9RMqfxpLCu4RKUaUVgL0bnFOOE0hPhawnLJqFyLktwWb
+7t9t3YTaQ9nqwlWiRyAY9u9wuJZTlQUX8bsOHGTIClcxujwwmprDS7VIsSbKBB9
BjthgFkdOajbJmM/2YsQGWQum/0xNQj+nku+YQ+oNA+Tg++pGTvl0t3rJznM+Z4D
y32n5rU8TG4J/f0Nvjv4dr7er0M7bdNMKUPifQfQ7w7PptDFJUg/yzrx4QCJkeYb
Yv6qV0tBZa6hEiKmcYlqcEPV/IKTU/rq+ZQrsdvHZEUDsGl7si1aMFeElS8yCm98
MbhonvQMAnP4uKbceIiLrETgGCB3QfPFhfDXIearYStKyf5uFzSdmewRHjmaQYnp
XSyD8B/ZejzawoJ7TtnD1JEOh2vyLoWO1D1zrEf6dHQxhGn+dZiwQWU66nyy4aFo
VvlPMYwyRc+ixVhq/yXKyb+DhyBWdK6t0J3QKqpn3Xd2lmbEy7VMRKIQjjiNj2bJ
FM13vZFb2yMyg+0LjtxQpbeOw01I10bYPKnY/KKE+vNWr1WKKR21gRKZYSUWWN8N
0VhQysguNVIidsk2aqGwiujIuKdfrxVwF2LriKnuvBxTk52YCMD5SNL2ToEjl6FP
71uXW8jPWXm8SUGqwQWb9i9D/27Jbd3FKuqNgOAZU3vveHS1JXbg8ZOgtzHNmOZM
MN/X7BakAYn3L1iFKwg2m7mW+CViXLgLQ7IDPT0CyIO23pHMY6N+jokOzx1mVy+X
CmwELvDAoChol1LJjjw9fkTgKTkWHXL7X/Zov7vnRXrmsQ8vbsQVgQGcKWK73KYA
RF2jOPOhz6CMHV4fxAz0xMJs6gyCeaOlmH38GmB4s/hTqPSQNADW6WHvaqhsmV8n
LgJx15NQZNbYF5gkxNq+IQV3kqxTG+O4e4IyMsM+6fE4/nFtUgFhxlRG1EGpmrBX
mNB/6AhtcRzLPx20VIKGHC58AgOGsllRrRSKvb8w8jJzmPx32O4auc0XUKJTlOTn
yxgwtDbgxE7rr2zeAQQQbXVGdDBti2vr2YKfQv4pxeJLU8wDU+63f4ig2IN0gBA3
/IdClGeLwkA2ec7pMCr6FGm+sndokNej+yLPFfYkz/FPY3d4YqwrNqCQ7NnWPpmS
Tpin4Mu/XgSmIufVxWF7pcN3nTAMhANhgl7cJwuxL4dstZu5ppJj8y9hkqC+U0ba
k2lgP95zuITjikdQckXJsS086WRT1yitqZ2V8/zwtG+tK4c2zd/y1xrj4UFm9Wtq
3Rf9z2v7qL6W2tf2s4iyShN/z/osGx6GK6CFh28dez+7Ji2BDfyqFGLmpvwoT91u
b+9qbfJzTpjkqqL/ejAj9Wmpx0FQ+OERzXSPITcjTbAAgnzgkqkqhfQXdW5aYiFh
ANEaPL9Sj9GkgLxbuHF6NkmgxrYwzf76/k8ymBZJbTdu1bEe743J0if1HCNscQ+t
M9ENPuIlH0Xg52RsN3KO4BJWGY6I2xT4+/dPR13LA9ilVxOHsJCDZJLLAQpZRE7C
8E33PpCLQus1qRYtqwiu1OSorA+Hxsjbt2wUjJhxGSWCnmr6FkKtXxF+IUTEvS41
IARVWpvEM8mJTHxaawipJp6DufqgQ/Cb7+Ka7FKqwca4XVVXS7sNsfhWkrur9GfD
/cC6dr8+JXEoKolWJR1VlsGz3rvecvyylHxQOqzXPq/YKt/gGuHA7GUyz9fcgtK4
rI9iQqPhk5axHEDt0lpDsGK672Ou5MRnyy/FTQSP4XbaSBbmZ58EZQrL8DK0rEK2
gIBwvTmVdKyGfc4n4adf07vqA6G4AroNCaiRS6A5fQFqYGunjFXwRO6voie7cuwa
GXRYCsAKmICrj3gUelatmPkAbJk5GjOkuA8IUOzPVcBl4LKKCsNhLWoNa0t5sRdW
Bhi4H26Zsaj4COfcWEwK1NE42+8dqLD/xda67ngZF+DzmtztVYMPFu2vJ5xCsuj3
FXtG5ZxDgzaU3J0+SrCflslm5l0e4vGjhIakttFbC1MO6Tf9akYlvQ5GYQo5G2IH
K3AoyxsX/eKCAOgZpz//q3NNRqF/WDH1Im9TZkJ6rhYYOpxYpx2XNUko+4Lv4G8S
fle1oLFqx2n1RCQ14jAyvOVJO7pQchQh0p65v5RMlK7qr32rwhqaKUP9Yjd/dtLb
X1xJonsRgv0r+LTGwxvsd7TorWDIA0y1Ht5VuL65sFYvrEIxnfZTeybADIkQHg1u
wzqbZUy5aG7f8mWe11qtYU3YKnf39yrO4OrtaUiA5voj0evvgmEUL/Ze3NpUUQGU
Lu0I+FG3/nHSXzKVmU3UVbsduQbZAf+2qKOus5Xz3HNea/LOobQKaY2sQuSibmFJ
ftbmU+5M9Brf2r+sQ6qwu4gSi7uCJ90mhx9YqZ6Z3nhGhGfrD57tD8P+ybzzt9/d
3xif2Ov/oRT6J1OlmNscQuxfNjSSDnzTR2VbPU7BXdgoYsw8JsX61e5Gf2OvZkI9
bhZ/6CzGskhCkkZXg2KH/zgv3imxa6TJELnrWbpdBdolQEolCnjYCc9M/9djNmdg
0vzYkKf5qMzAJFvjX2xg5NRo3zVxZZQQULixFt31YhpNYqqzA0Jcx1KX5tti9Piy
fR/PWc6kboYFGUmOMtUtY946apG2jGUBdHc+f0EH889yroAPjaHu3tWNAAWUDrWw
nW53fQ7C6ew2nQxXVOjEgVj28sgP2MKyfGspK3ebhdvJmpinIvqKYfxlz8sswUv0
UqOVfJ2X9/ddNNpW3JevCDdG4ktnfqpMm47WO+qYKW9nLwSFHF1ka6msEqUe8/T5
W0AE4kcqPraMIPidcVLZ+ff4LjNDNdPOpca8o7ZLjxVK4rqUeFt9DnAokKL9+ECA
fDA3Szc45RgGZp72kFeiCXitkf5NYabd2Q1wgkjYIcnaGZzkQBjJXlK1vxrQOb4s
OUNVyxuJqE1mz/+jE9YVgGzH9SSlaMWFoZItvrER1iEy/Mx3xeOkYzXA4pg1lYs8
KrZrf7beBtVs3+qMFmFqn9BMX3BYoutVYDVccrG63yeU2JRmmS1tuyAE+Oca2Bxr
tN02kdMtRMPhBZsubq/xwwBrrmovohVqGtmil7QRAFM+NzjRmF5PUBFTdDuF61Wp
pWCvcEsivwV8uCFn8W/DAO9uMK9kmU7vwls5f6XrN/ln0GgnCMb5KOHWm0tqjaY5
nI9z5mMN+RRG1np1zGRae+Shzl5LgONnA3D/1GvstYyrbjoT0Eb1AWY1YB+1nuwP
QtlCcEhdT/r613SjydDyDfC3FJg9U0gribnQ/hrcDQ2P1xZEyO19nGCbGe/fK4F9
6jbCh02Uy5MvJbS6B2m+dHY0sUKg05UxhTuaYbfVo/OnybAt4/s8kEeF0a/9Xpkr
8qMbytr+LJtKzEYf1vixxExl7vAV6Nuc0P9qq9GQsMDvEF22oj5UefNuoz+nakBS
ZMO5fjwsQv0rl4sBIQa2MYUnhuqB6uft9NTNxzBdqeKCz618QFGHtT97T2ATBcCp
6RlKPG5e9HTo19CZAzW5nBU9GHik8PXQ+xbydoNlnhSK/bOpebQDTYV8AMK9rRBr
+1HnwEP5wTs03IqhbhOUPTt5ca/ps1D6KrYvrHJDpbJ6d/DxtaLMGU1qhYQ5TGZP
gdp/+1YqFNE+nqAFExLIu1K3kgOBu8NzmD+MwriznZW1kISM9vXFNrXgjEvarKn8
FkcDFav4ar3b40kBQ8HzUslAcdQW9kazFDbaDel5HWoOIozrXD0sZrWqWdDUdqYw
wS7AIR7KdqUx0palX2JCghkWsNEzvjIJEhNWXFn26VDmF+W+RJ2Z/RUn+5MMqZIr
g7+fp36wg73PpQnAXs/73pWE+2vaOz5OseztX1ED3hleuoqQsyWr8wmSIM2BZIa1
ot/VYTjzn/EUuX/EhQkEb4KtmpHPStULjByBSNF2+YjmAbbUOVY93UbX5XEgp2NC
EfhwQjd7pz2o1o6Tt/JUYnXEfabmeVuIKbDYY/gv+S+q+1Sk+Xd+5eKifAEs4ORH
SAO9B6RIrf8HCZea1GmsKuzaIjywK+K86/qSNtehSFuFtEYlj8FAdXmZEQJbnrQZ
V4tjWpZCZNwIjDk86cIAvoCvdXD4b1FR9DfIKG7+aerD96ZQ6jmJqWU4RROtEFo0
nplDCQnuDDgbGJ4UWku4lq9SrUNrVvOjEfhNMozRrGUe0lB6pJyI27TMC68PuMm7
8fLqTXvo9d2BpbGh5S0ebkSRIgM9VAMzJSBz8VckLGiceQURHvfW/Skeg0mNNl54
4f/uYQ2yehBjdneLXGROT57b67hoZkRnFqp3ZWlBcUbBCkXnSZCJdr1HLVm+NbxP
gySkeJxwIYkWUvdcB11a8bVzk4RGdTyNPWrwRK75tobMU7ZslvPE2HmgbzGUh8Uy
CAwzKUKcOVb3tocjuOTglqQBRFbwGW+3v+XBqC/2V/7m0w6+HvpVmIXpzcPT6zN8
TlvdMeTo24QIu3hhALh0yMV27oOp/q7n8zBN+ypwq4wUgYBNXU9taEcta4hALvX7
BOYseLr5Eb/aUZKFrnU4/o7wBupknCrw6TYq8/6jkOphjHl2mT8Gk9i6UGlvPv2o
zorfn6ZD9ry337y7ftfiZctj1z86VoxsuwyNjozmjczRhX0k34utX38vt5XjKvYB
6Jynf5D7GlmT1Mcb10y+d+AU8/nwQOPuzdNHf08FnevQ44LyKSDmGzZiSYX2z7j0
/I9rfZrxto2yiVLVNG+FJL+q2ATdblBEiRg6u8pR7xSPUfQbFMZjdz7wqy+7JNNQ
3ZjwNo4JMDycRHRL4N0mLmUD+OjgqA2g0rQ4YsZR3FprTp/LdKG3HjLFkZeLeaTj
rLce/+1RJqX3VzxEo+BR2Py8cqg6IJAZnoG5pJfqBxGlBj/zVIXYkOeuEhrWILwH
dFKmrUc0HpwV2dmlMSHGnoeAqxgw+XNHgCk0TozXJV8ToBoIy6AE6Xp5sgGM/pek
b9LSxrchFKwecxBBGs3Z/nP+39wKr0MiDW3GsJwkNG4teuOvXp/nLtzb4nJc9z2k
04Oekl02Vg5aNa9PxNgV7vuEaWlYVF6dsoKxuJLag+SmGHNZzAhr7z+9mFSG8St3
R7RJIqVXmODRYnutX9UfxBHq1pV6ZdPPbV4NcjFkk1yHWdfsPmMxrTjytkRNYbdP
QQuXKzRtX9borMUVRT+C8SodWUKu1AC1PUNhTD9DV3LZrSYxUoo7USCw8ACp5Knw
BaP6hThRUpHoOaZy6rGWqX4PQHKi2wc2YR8uIXlwsA9irOLWdPcqbA1K5M72NTHh
5y+8tnSkH/ZXpPCuvp6aGWe1Cr/JTFf7QogvOdfUyzLjVBg1/7BJ/ppq4CHbruyA
axasyxtbtWZfp/X0k5Lp4PXMeNXb716LqI9jH0tsl3BbuBQ3IlFtRbDISOdWk7AX
aUbcmmWjW3xk7oM2zwepKMyas3KK95UOlvIQ1cAVv9D+Z3utGa2KouFvBxasKXsl
C6v8LDKzx3ZAkYjmYWR3QIPMjpKUtqPRDerQhdHBrSBRdJGjafNHON9o12EnS1UW
VA2R+2r3a/kx4jIwFGZMBBJxfR2dFHvyE5A2WfBiAjsdF4CG0ZSi+cooqKqO1yIL
Yt14EBFZsBiwXU4HWsHp53HRtPAI4Azz9icIlIoww7A2R6yRv2ab/KffgzmZeeXf
QrMqte3/fMKRSGrBzab8cLLW2/522F5WqH0QHeiowDSLPwY4aYJ1RU6zY4SQA4f6
l9VR9nEBgNttOQhEwAFr9C24S66V8Oj7g87NBbHiaAbkTUzmbkBXRHN/yiMB85Ss
WIv/WFDm0+b3iCzliy8ElmFJt8XqjY7gc7zeD6O8qwj41K2CT6xo0QEJobdZYLOg
w56rI9Ze2xyUaMNAxO/ZYJg1QLVUnxX/FNOULta942nrmpTSSZeGZQMsT7J5wYUv
DHFj4ig8TmADx6M7JN2LLrMvvBnFfKjIHuFtrD7TfbTGpazRWHOOFFKxxwzqOuCT
e23e6IBzDqhf8ii33DDT4GtWEEpEWD9Uo3zwuUk7uJGH0ux1+WykB51cWbA++av/
rTv/yrvkZOCs5n+h5/hL6UxCkX1EYAAJJvFYdchWFYbjPVBMPbGo5/Mapg2P/MXA
hZR7CHlVAdjOltR+55iIO1owCQBCRDAK7wbZVkIPykMDjZq1BON9KA2f5r9d4tds
Mk8PVA0qQQgwr9TGAtfvZsCthbRQZ3oB8vnjsJpVIdiyZUU9x72pOl2/8i0cN2T7
YqpH+goPzEVtx05ytmDJ1EqP7XUBc6URlE5iu3NE2P3NshQCXSn79bdTvnj9aIeI
J+ze4FO7A+Hd8YfFzrVhQGVnKsflKtjdT7SmCHyPzfkwpH5Foh/As6AcB4mm5QMW
vFn6dYeiM4gxLhUeK+jUcC4dAJgZYqDonYkCDpXoUHmfyER9evFNgThmkBS9lFij
7zHFl+2tsQarlwQejQk+yTGLNPZUvbADjGPCHE4sqgGAtOMwXb11absFvjJ89X2x
y3ukYLodFMauiXrnR4IOf3WW5P1VVKf8SJQQwcVq53DBEivRKRhTGEFvbjIIrP+Q
Pg60nRrgmC49qqebulKGZdZsIb7Xxq43xvOwDOkomqN7KIzgVEVIvdDfp6CczMQe
8XacZBWqSyYmo6/M87IEJWoB/0oMvHwutHGqK4MN2ZC6Pf59sOjTzTAR60uqzlGB
QMHvD//3QixuefkOne6wcALOs9TNJbzUpc9RTZHUPCdLvLwu3HflE2TaoF8erihh
vblpxzPCoFJGWEI957kLyJDbNmMi/qb/vebPF7a2k2IeigmMWykhn2T6BpuQAFVa
Mjtl++oBpoPs1LzCLFzOnDzVpPkx2/9WKa1rKzqoGTBQTXvZXqyO/Eci6NUeFeGz
HkQivoozd0ZcjnP6R/LmDAVOcCEwccodwzEJ25u7EX/deN0rdUIMIQJ2KnQbfM52
YdRT7z8NnMBxJFgO/Nnlq71V9U9eYIQEffTrWfy/PHtjDm9ndaoObaggAfnPXL32
VgJYmavhDWq72fcHLHFildpbWCvADsh0XnJsE0925Xe2HG6NcUarSLZiUdZqv+Mw
JIWDh6Ppt1xDupMwQDR62QxxWio1SEQ5RckNSJ4uNElcAasVlSMJaRlHqcIwS3ZK
0ECksBVNTR/aMlXwFSgDpCX7vvh2WbQ4BzRxzpkllfw7d+JmxIrAxxbKpOgvuO4k
Z3zJ2QedKLQPy0E0TojDeP4VYifScE388uW1SCGyXDfCoSiFqqXnrLTtzeNPs/2M
jfKDNRRY8nyy2Ylzi0iq9FX3KNgoI8rhY4IP6vx7/KF/6C3XKrpdgMHKqGBYs3/u
4niEfIxC7jjlH8NvVi4iGR1GG2drFGcQaF7SvoGBhS1lNTdjKf17s7yzXJKNKozZ
RaVTgaTUNC7cwlFRqqnvY4zgtbAA+DMpaMMU04vIj/S8UmMS4mf2CCCm6nCR8e08
WimcU/KPAcVqkho8NFlL97lHw8GwOrGr3B6ue2kOBY/fth9a3TQzTdll2zc7aZ/A
nIyjXoJhdsF99wYSaZ/V1RMmQaoSU8F/+/iIvldFIZapN4Gia9G3sZcMbQrfZ8I/
rPstx2SsGv64DVyoMevJGkV6M9K5u7Rl/qo875YsdpTHhrHyNoJljzQ+THEgCwjL
erQptRJgsKW46+kWC5j0/ppLMLX9AlDC5cjK1mX7tdlKQfpHlUvY3Q/YYCbRKzbo
hSNeR+P+kpPtDNYjz9iOb9L0zTkMzphvblDp0/1KZcSE8bFJrsqWj56EFklnf7vQ
I/b8tYYg09YHPNajwjfguDprjGfSifYVqZix0eilJugMLs9QriyMfKZ7uM64vv3v
rwN29qqUKl4UpYX6w3iYbYJ6gbVWy1yM8ALOVcDfPwotdUPv0DCdG09c0dqFCPDg
OD3tXxGKGko8GSVNHpxjWuFfBIyCYsdj0kJZGsB6ai+89us3Foz8LE1kVeq6mYQG
aGHs96LRCHBoHc8ouF2vwTciK3QP5nERPr7o3HXpdpHZVIdXzxQ8bgqcDsjWv1f7
wwK/3/3Ax2ErYbJ02g+WHBBuxI06y8FqpZ0jbaIEezc46cVfaCpvSZvwTdnBtGLS
noAyh8+ViriWa0be/YI+xwAJXBlEoNS+Mzke54ZS4f2jSbrk4m7nqTTWPm86aAZ0
26yBnbH+N8tinNlHX7Mp0uoA8V+1aD2aPEj+nV8el1oWzgZkjl+cUqoa3N2vmq7o
Ffvnv88G6ThqQBLDyOhiaY0RK1NO6gUbsa5YvqocZxAoGnjx3WN8l/YYdmdWFzJf
WmtvTBC3mFQo2MrUTHnqSliLotY13RWMjhdVpfs2rHXSn8lRz2B7yYOejcPVNq3Q
Im9YJ7VYnDLy6y5HX39QWRBQJtZ7opfQ2XeaabtfppvCAM1/7B36T7GBnhyNdUdy
SmgJwCicHbwNaEOTcambqN77F0OraPRM8oTy1Z9/W33NJ6hG62ZyEEY0tCD7jhH2
mPeBeQcUGcyEjxt9GPu5m287+Dy8FpxgWN91leGtis7uAjHL09Qc7m9rYbRqgpwp
MI6eXm9n0gjAAZAFmajxVusNN2VSdcMCEi6gmRip3WoAkUWiSA+20ZnGfSC5u8Np
H14IJxr3astQ0bO2wxChbLW04H+329XdQvn1OndGVH75ii6DHNe6RQJBE/FWBs2t
9VkL5QD9NrdLgU8s4CIZ4rOi2pmghjBipCm48sC9R/lmpZpHNv7iok0Yx8he3fJd
61T4+Fjgds7ixf3R1PbPalEfq3T8F3jCWhged/Mpkin+aeZvYiqR28uAp09OTQ1N
M4kaiWTF/wRz375U1vnXKDijqa+IWfbymAoud9LfDnocW/F4lWL1ffBdxjqltAWW
Hd+vP+2G2t7LxXMm/n7gtZRoUTqDOH06FhR8RBNVfpxFD7jyRCjMOIhIvo5xq44e
zIl4zGewohrIoq31NxncQImEORBALHUy96qkSbjlEH1ed8FTHs70CR4eqs5BhSTy
30VW1NgzXbQbi4oYQH16QSmEB5bjTWUSdMOeB70Ia/CmPkv3McR5gOSkX1Ad5uST
3MC1aDrfYzxmmamYuFbY15L327qOvt7HHGbyC5va2divFVtbYym8cJ0wCHEggh20
p+Dy6eI4/fe6Ev2t2DMx+aKURwKt+qh2e+hTx/ExEL1aukKbDvrw3ykvOebIPSLd
S72C4zRhJc6IfErc5IFajqoBEosa83BtHyAgbSfYq/wEPrY4LnD+Zf/ZPmzlypRk
AxO8imCh3YnFT6OeHzU3X8ifxePvNGIyRjpUnLLJp97dzRTwCQFIGZR8WalqvkMC
xuPHN24BArc5qFi4h7OQW3Jx4IHNIQxyelF81bS84IiWskHs0Y5gNoyAmuwdbb8/
Kvj56aLEOiy5d2JZvaR0315amIzlV88FhCLW8ugsQfiWnW+LB+FuM+TAl7oCZGGe
dxBI4ZVkv1kqaBa9SJRS6+sFrZBNfrLbwbteL3MAtyZQcfxMxE1N1nf2wP+V0dsv
HiLXh+P2AkYpmZ/o7pDqn0M0hNqrdGgoH2voKhI9g7JsaPc1yR9lkXCnRFQccRPa
ieLq6mpo2O9ISI9pUo6Dw6rYwznslQyeF1zGpQ2+l/tcRAd83Ocy2M8wW4iNlMsd
vmB3n9i7lrfjzmKu454t1bIgnJXmL7yXYeZnytdjgsDtP4/7xlsxWFSBdGLGM17w
/Bx6Ev9i8aGGIJ+3W2dwmg6zIw2d7G3WF9t/1920lGPpP1Ad/BemmNIO3pnHiSv7
P87YsHDOjxJQVmqVtgDt6EyIESveh3hzHoQoWoy/CcwNAsTnG9by/CV91JMtjfdr
/I3g9aafTB6RWqWXj4BYuHGmO0mxFPtt8ss1+5XcZNTBzuCt0YM6RQhc5fbv/TTH
M43CudIHpz9jwWyRLUQvjWGVgueaLV4joV2tf07oeQ5vXQQ2KpQxG2Ox7J4nDj1K
F2mkRxOdHPAZEI6NfwsvzcXUum2QwHmDY6chdBZU7cIKqgHvjB2SOY/KngWY7/LY
Fo4pPzR7GjlTjZlAfCCFCcxvtiNery22cVC8ecFpDbsRzKT5j26odxbd8cAdJ1wi
QrnfMXq3/QT56JySP7f+nX8CMt9Cwqd2AsW6Q2QC4d42TwSguvc/GgiLP3KrQ8rR
s/BbQsb4GovZOMLQgGNn8f+S8mMHxhL8GEF4fMRk8MYLtbybrp/EL4pIVT+EPLOg
PFmfnMYAhoNN9+bRpBMjjzWhks9S5uNtQbq7dD27M0zZyPtd6XGhik/e8yNbYGKC
NvCSueyZf1J/u8uXgBXtkS82EF1iDzD05HOIMTk3DU9R1Svhusc2H/K/zr77LP4F
sP7qsjv3ZVUWr5NVkjigfEDtXujm6Hs/XeURC8v0N8w7xnDziPBWgLAueNeWT/hM
/0SK0jdD9ahmqTJ92PTbr9HwOQ7LxamqgcI+Pzp/H+hjCy9a74wiJKFhDl6Gu1jv
z5q2qGNy5YRpQSkseluEhHSubMJh1zLe5uXev72PTM5pld+iMg/lteFtY74WhYJV
wihVcWJPJ6/xYfheZrRjveicgHGkMjqxuM6ZleITb5aogpgzWes4KwtfX81+Jug3
TmWJmwoJZi5LxVAa0SYGI5Ng/e6lL7cmbyjjetaJTf2SfTNW2rdNMHYo8dxV4GMS
d+ZWaS78wccp0q7GXfuKiMSwzEWoMySU2ZL01Pm1r2sf0VgKwvMBX2/ksq1Op6Ku
OrlYIdJGOEwMdJHHwHto9P1vBE1Oq8w50phR9G1FDYDZAXrWyG7eLXINxyA9SJlo
B6udNp7mr8ofRVtkoiPD+HJHzLTw8zATNSjLi3hTrVCIWfIXk5kEMKDrZDUGprRs
ZYBsUCtUAPepE/ZuwFCHk5gkKudEy7o3X4KHcQnT3MUC2QOMIvNPFfog8ohU3KaU
rXjr1XLHbIm85ipKxkXDTa7nm20bDqx7Bf9wvtmTRRJYrrUdSEk2MPj2q9QP4N2y
JyPxXcU4vH61pSeYtzNC42B2hazIxnxPhn9E4uj53QqBMBzpKfEercTl2ugpDulj
jj3XGV4eOtP5Up+jZTULtmzrRymeDJOr3Yk5RboZA0eisDaU1peHGuu1L7CmHX1D
3qeP7w2yQZ4l4I1ETdVQT+aDIpeHG4/cRnXCtWZC/vp3XtwsgMkLa/fRCiMYx/rq
1i52TTA1ic08sCdjR3tPFmJ996kNZykIn9dtGihGHyTZXruWshBQiFTOD3/OsV+M
BYwYZIR0+c2oFMx+2H2XVsMFj0GGsK5HlXbaRc73YghQqLHVcQU3kyAHVWarwMom
6aGHXO+3TNj4jDg5wYRD/Wga2nXpLyJlLUFqRjXL2P6GyorHBmC4Y/U667ucvVwF
YnrxEYaIYYDfz8tnKfki0bhk9u26+dFR65J56C0SduAgGvA2YCCm4zzlfCYFJjvU
1vHW5WbZfGli65TxYpUhT43unXlZJusytRy3eu7cn6PN7ER+sMOwD69vh3QRzZFF
WHum8E35YeoYctjH2P1jlYVduvoDZ/CSp0EJxkeeJqFQZt3y0ebngVO2RkSKwD9z
mA12vCx0hNLMA63F2fBFR7Yu3APmSug27MKo4/A1ILKLuOk0EmmY7deiuR3Pev48
48vXv39q6cj6llVIV/nEoOIH8JTjizEcfjZA3Ep12Rbj6qfH5R4KIFaXs62njWtQ
3C8q5259Yv//6E6Zzg6QtLbb1Aemn8OKTWRlbl4/hbEVOWIaPjnt6QMLU9u6Q4wK
A5h+Aqf9G8MlSKz2pfWECNMxIKSUJTUGNMjMwShVNBjEsvG6MmJV/WoTeHHT/Szb
B4aPF2+uI7VzAYCPwA7xVbiVY4yjgvNVbvIfdOtyxjHFKaWeAdnPY0oQMlahTSmg
NSaeoZZZyUMnMNt4BdX2wt4wrUP/dt72fxrgjlMC9/WtXsYJSulxkH7j1GAbgE7i
xN6+oh5QAPYeZcrTgWy6TKg4mr3fLjJ/bhgI2SKvmV28TIYlmEWMfkZWaFePiBz3
JztWgEP9PE5zQYR8GMq7+InoFIBOqEBLLBzFT86ANX7uTy3NdmeR2Tt7wBwGYa7J
Trj55zhNbUbtbQreIYi9zerxqJIRX2gyW2gAVG63wFiYDD0zu/VkasioJdhr+Wfv
37cyhIyej2DwLAbVOfmwk8MlCrfgSHHIxsrRqHqRPT34q5EqN3aeUmDqQ2gP53uc
S9ly+sD0vpwqMKB9nEsK6NKgA20tTSRfIXWvCp2t/it8LScrMTwsDWYeO8PBHHfb
SsE5ymgLtiAVgbUQH5iFXprVOo7GlU0+NuuO/O+md4BViR2En50iwVYFqmxMgcVW
Yge0c4QZcBw85XY/yVA8inqC0/P+3wUt+W1qZuJH5twuG82a2BHYMbOs4O5kRlHP
PRlXzCFapliMuZBRhPK08IYTlBc8qJ+xkA81WJIrmgB1XVUINzYMVoWBvjxYWydc
px2uqqeo1Ltg3ydGXzqcQvdEhoA04lkGqcCz2K83I1uRfRQmlzajPIPiS4BVStKo
qzfVsrvsRAqQo6j4NY/8dBNC0FPngiNTWqDL7Nj6tXfNoJPO5ydnW7mMu7l6N8qY
pFaL9SdL0a81Vo1sSkfjtgcaaESW/Qkeq2vNwSCZ1Ms7AThhgaIm0mTxtK/SW0ol
InjxnBk94p2SwiQ+2uAwosd+Z/qj4fE9rUZOLx4GrzB/saUv6gEKxYwclx+KAzEy
gemUczhJS6jrtZLaFFrRsp5efMtGQd59IFuAsVXv1TQt1jCSa3PDxYdHgPRgcWfX
n6d8j1fobWbbbRFY6kSMSDL5wbuoCCWflemnSQ0G8by+0HpcDej5np5/WoiAzPlw
cka+n/PHGKlDuZPCvP73sgqzWV95kGPutFW9b6u9aHTCDuIwo/i3rnFcEprYphKo
F4qNBeQSK2vZ61kgAl7sHbsOLGUeXnJS33esM05LhFmDTRpJNX+tYkqUQqK5ob9a
GmHMKGXkUoaEvCtg9om4ULxD+s38E+xVE5+W3w8Zf9nX0P+sVPFiwF/EV0v0XAz3
V70k602vqXS6kmqqJge42aQft/ZjnrPMvthXjqjT4Xn4HhF9nEQpYEfn2gEumfQR
ZgWoWxb204jg4h87dw4xM2OE0BtXOM8w7DaOfgKSnfV3nBeSLmwS3DIYDwBGyEWi
/MQXPj3hoshGl8jKALEH0o0Vp6k/QisVEFV0L8MOAnoZOoKBJ92K+uHHUPnenPke
c+FUDpOa7qwYZvYlgkzkijH8TKbEM653o+eKjdQEvu+SGRScuxRw5lT1sTBSL5rS
R7wqisjbm4x8dWb0OIOrzsEjfQdKWYuV56+p1Wm2wu4lWCVqPaE1SpsvqTxXzeas
nuqCp06wjtOWbM6OsgaptQpMhgyiI9FY9BMe6HYTx+wbJ8Z8MgeaGe0mvSnV2tv/
47A91tIjVBqFnoYXHn21IK/khY9FLULnEWAPn2cu3oja0e7CIvIJbbusAaLldPI7
kB1+v/Jk8YZtWXGd3AZt5+aJaISBLGE9IHAb4bwkbWYz6TPDx11+YoQOqMde4Iob
0/+o9V3IVIOVJX95om2dhYTzgv9WSM/KZm38pIX0q6qdPkh77mX/t9QOqiVY3FZ4
0TUAcDUYWEGFA14ZK4UP6eEQyhJqQkfhRDhnfhFNdiY/GAA0sDiFReasYMCiJzxX
uuyxtp9bGTogrkZStxOVzGMGzAxCspzv6oElAqnG02PIFskp4GRJi9Jn0TLCJGP9
mUnqozT+qjxuzP07wFZ/V6ayriRxNPAMbqut30OkTDBAKkPFbQhgaiGxgr0x/8XS
t19NWaagoHn78fv3N0Q2h4HFFFZtgehWWwIY9ZSsXPovuRnPho5SK6VvNn66E0EQ
Bh8X/9Ka6FRCVZEkb0r0GVV/cvFfd/tWWNPkDp2tyVwsFT0mXZdj0O4nPPEznPxK
3VK5c2a00DuwQIrgHugxvgUNp2lLlNIfR1Nta8EWx7jwI+A+gZ3S/FMneu1dGFcS
QR54eOOZU8pGks++3rA9P4yr5zAije4VIdLw8kTgQXfkoCV524EVQGTwY7t+lbhb
VX2c/87AWTeLkQ38viw4aUHAxbGgxensH1mIl9TFPhJmZc1Tja45AN+/9WvGC3fQ
+J1J/gT7jPI0YOe0bglmdkJeO7j0EufDOQMD1i1K2gqZXIf2Cyq8FxNGFEqbEYPd
8lVUgk3YxzVQ8zqsgkEBG9pIvnIGR9k/wvIQzk2p2SSNg2rzGWVTulO1VzSCieiN
7TGfGrVjC+jBpMMne4M/B0sdLPAMbl3FPQxECKZ6OtoOPg39fteZkjDCPrmm0Lun
ZeQW52ZkChjGvcN5nUWm7DSUTSNWdxkQ8vpkeAl9jvfdnAz5f2HDwxZmKqlBsyOZ
U7bmczKB1NKkKzCGlfWuq0ITeHQA49EPkO9Ol6o8If3c9Agb8FSgpKt0uHSuJFi5
FLvsIa8rBjMFzeE3/ttVnQN1TjFHOu6BkOed2FvenM7qtvHEoX4wKV5DD4JChmgR
JOpZC9knGoQ35cQ+mNCO3+Lfh6I4xthc5JxOM0D8JG92bfbC4FTGUJZUnyKqYDcC
LOO4G6bOclWxGho+ZmICM/gKUydxGKAk3G9DWWVtuRaxV6QGFNxCzSu0prO1PyiP
Dyv5Hfb1LdMcx9Ctr38iOZynjhyYbz4Z79zNdIjvk7zdHXr/s8uC8lGPkEybHpqb
EOmWu4a/WV7inRF8s8TlN7l3ZZefpXBluY48V4e/FgtAm151PBtA7J1VoFWaH4+S
w5NIbqyErw1yYuh2Z1rkUXPckzynYsZxMaCqwK67s82S3IGuOixNe3E8jZi7X6fL
EjO8KH2JVyh/3mnlNDSiCuM7Gi/mh73ETUMk2BBvVmI96ByDOB+wy265RoOPH8QQ
7R3k7fYYWVghTTS9sSVsj8CPiFN82CcA661ayDVMj3gNT+6FjdkTn5+qycoN24Eu
LMzIfY6O6H2kIUFadCATq1owl6io66KEt+b+sZUUSeiWdIOMuX4dYIVFAtWX9ZH/
LLMmKOJfR42ttTo02uLY6EHlC9JXRrpBLsZe/XZsz/wBYjd1t4BeQR9yGdHpfQ9a
znJ/DBNdGfCudV9F7N8zb6zT7YxqSoc2kKcU4MlpvXLUL0F8rjqNgKl2oSksq0iv
YZ9MZ1KKyCWhwpx9Syh3F0dtfpsyGmeOkWSMYB9WBz1vw6AdobkBoyAVg7PGbP1e
liVvxV01BxodYFXZMkhqe68hj+dC/UrPMwbKBAfXy+DcOTUCRPeuRJvyUx80VWjm
+juSZV4S4yDgRCi7NWnoIAHqsQ5Cuth7n87+MfvYFIPmRGl7HjEYWJwQhoMRvquO
ZOKCnGL1W45+xC9HGipRy3NOiXxiQJesvA0Y9fPkhWvJNWL0auomMMdY477XjMpg
CC6vnkKoOs9L7MMxktI9rLZ52O42e1ynH0HqtTIpAiT+Tdt9qZt2joXatuuRCQQe
PcRj8O4PAcpXOFya9D+diM10WSlx3zvz9rXSMgJs6nFlFLbV3KAgRpwjO4PaZ3ps
tFC5Mn0FhM5XCrhfWkXRIftEu2ntQkBORcosMCtnEUgrYHhjeCnRyITtqcC2BDwM
kmZDKL2XnqCWjDs1pe7YipoGnAwSBJLum9w+cJ3v8yvd4zUEkir9BTYpMogO6WQy
UnGi24shI9QVHAOGjWDRHk5L71x5bhivPLQaS+Uav4g3PmaT+VCk7XdDHcrdieCf
QZcNOFQ3AK+EQ6FKtUjvFfRGKOijW73F1BlI71V8jWZ3ot9vXNqs0gCZgcVNsdgc
L00jYW4vus+TlGrSKb1PDmht4hpWIRd92SsJ0q7g0Gwde6NMiUyCiVKUXFPV9It5
Gp7uXr6FiCuNJoGnwG22MjO7pXjVkFwBBSJC6E7rCYOdC7LtncZdPUWcIoeEVDg8
924SsdJAg150xRuglLcUpEXf3NZqKMCeZMnrBnHdx+1wbQ7S/UdjEOk+k5sHSqJU
QLEbxCUwiKooGVUH0XBPRPt33I6P6p0WJolwXWKnq5Hnm//2DtrCewJKhdnqSKf+
vqQ7deLwjwVGI6FBlPSHWYOUGjT+fvQRSot1QBxBTznn62T1MAyHPgIXpCJ+M1re
pZxfWluk3Hv5kBg0Jyt0JAiDXahWbPs68F9fokmb/ARktxHHQD4GOzoB2ZQm1ACw
w3YgpU/AFhaiMmgwuoMPp7IvU/h9C4s5R2xBmOCEMDNn3gD5sNs15XJuABoTbdp4
ukPgB6daJKA9j/TvdNC4rv+9EFvrOK3Omh+RWLMMBqJxdXyqkIbC3hae+o9O2Cbq
CUySh5tp375TwEMhcmtQ7qsqrEyhu+iQFvlRcqenEnVkIq10uAxm+4wZjl5PLA3j
d/SFZSd/l20TtqaY5AfS7TRg/J6Y+xN8dqzScjeEizqY5yjXiTkviZlLHIo4mPaP
PMZ6JJy8N/TBbxdvL0bk9vd9ZmI1I9zCoyl6lOG8+wRZJvMvDlUSB/tNwqezPLFs
zkqTmDkwFx5SbQAmCECMwdjYZFqzG8q3gEzuFqPK/D+fSmdbVgTyy6V4pngeZEIO
IiO7F4W4T7zpUxO4mUhVyHDSJ/jLe2/qBrTVQWndCWAouCSRUDmvHvTsPBt7ndl6
sSKAKkBfpvxsRDcMcvGxvLrGfKgp6XpCL5tfNk+/WtW5WHqp96cDqJUH0hezNxLh
NGmUHT6bBQobF/O//xC1jShxCTzHKKSz+vJZCgYOuNJxDxOZd8laOg0cys6edMui
9XS3SIKWvRqjN16U29STPu2EDObFJ71Su/wdqFescMvxphsbW26sRYwync/iN2G7
Tx0Sq3FCR5tQ75jy327f5Jhkgb5mpiqaUhZWGHwKBvr+JyeDltFN2qE9sk3vFmz3
X1qIbmWEyCVwYvHnbFnsD/lgb0cq3ld3vhvOWGCGTx5y8Ad1kL/LUho9hXCToKGE
q98f0Omg6oLzu4jO6zEqDW8wWHPGCcGavnUs5HgHyr4h7xDdclH9SzfjrO38MVV0
aXWgqe6oor01S8NR8XaJzwGwj08TT7ooKw77PhI1xY8DbonSUhubkuXD09tb4bz0
eq+B6naM9NDFxFtGYoMSL0WB4V3CVDbR8LsftUrXz74LnddyJnJ4AV3Nugdm3Hkw
R1KZrz+4hIzKh1doEjVOZwfkTllE5fwIY9zBKmefffiLg2AqfkHFDNi7xhVg3wjZ
8cChZ2AaWP0q4zfDsAJk2xs1dFa9ANw+4xs11gCWbas42R2gRHtrGc82lsX5w2OE
xs3/2JE59orCqKDr3qV3klVcQWc1QMv/v+4JJNRaAITSO0dmWA3rDlZNuSj0eH9i
Co430V+/WoBlpWUXO1ppHNtT1lXu6kf4XF/0s8xNpcLLOq8uH1nL0J7bf6tGl2PD
52KO9dZUMlkQa80rHZ0d3n/X4XKHmkNJ8AIpjhcU34zAIPrNSsdvZTzZZF/uYNJw
LoBkDkDvOr3oPLBiki3zTnWWmoe2zG8SxGo8qLUNoZhtsZ5jgCsaXq+La0PeqdbQ
mZXClCw1IWJTp9L2s8MxramYyK+2N0o757YcdZqsojVlcz9+KuEB+TQCSxCQFZ7G
ali1KbVL9HrvflcBASgpzJhXe4Q5V65TcumQ7PF/+CaxWfIQnMdmgpPeEl756AXC
nMinNQYpJHLNPkBBesAcKM4v3Fw3mW4tCWggSNrH03LfRrVwCAbEB5Vb4MKUPhME
VjE/XT9G/2LT0c1xaThfbdytU34e5a5lZkYWklfGm8Dvdc4cp2iTCfsFFbDeFW3t
THtiYktG73WrPakBn+rjDTip6ahjGCWFoIBiOwBFyd7cfAOhztqdAWaUZD+z8RLL
eocz5tzPkasiq4kUZHnlOBYUq0JNDD1tmjX7xlyiQBNnExO+MiyTX2Ai5pH8Xm+b
0GY8oEhgR0mRSOPiFrzplQMEhwizGlrjabY+0fB98ZHldu/K3OuFsdz/+3R/Sz8r
k5c5oawM6gfMZ23RBXtCbAlQ77oZSkCeeOaqFkx+vinrCTtIAb+L1+OuxA/WYT6n
ESbIBrPsgf/Bvnhim60G8XE4uyN/TigP3Cq0+jsXl7VNJINA4G1HR0W6iJCJOfNY
pvWlcSZRdWM3j7wZnIDkDoMMbIlD85lns+gSrZhOtUf4YrYx3LPFhyOxZaQKLg1A
PX7/0315kIPghEB+KRlWx0QsDZUUdjKOLjYsZQLQPzNPJ9Kob5fo4nf1lMugaiNC
tUdCkILWLaN1Ly5gvm5PGy1GoayQ6FVS5YLfW7j7eZ2+sLvkljd/kY0LDoMEFPYn
N3qRVxAsWLPHwCWojrbfyMRu08NJk6vINKPQ6NDDIWn1puIJvn8deMgZfisWY6xr
02B1E9eVhgWUvp4u8yOTDys0XlLh1HOuMURj4IVhTd/U6NdxESC3X/6KGURbrCRc
zQ25Ey0iuHm2E1bBgruAAzVB7liwkObXnvHPalvVRlid9gLtwvTbMdgLaC/q0jBM
qVVMmYED2YxmGOclKbi/kfyi24Yrc/e+uxBlM0VZ1OMrv+Nu8rhIxOIoDXe4CJ0j
Nds1y9f/fOf9p4dbIgvPWgoVL0eN4GpuajW0ohanTRAtgo214ZbqrA9gagsB5Ye4
JPNO1AKwLCvSqXB4wx9EV53VEGTfa2JGHdyq6TBI6cpSwkdGWla7CjpUafVS+I/s
nUHsBwsQExHD+9mFpxA6Uoi4Q+aJgmMxJsxJZDQiJ2d54ac9zYmBkhfr0jxdlqGb
r+piTlrCtEAYYLCFd2upQ7zgk6Z7IawklsFEP3UAOHFwmMLxphwkNByHgTVVCiIa
AnPWxEtEYjvs2Z1TY8W8zm05i1hwMOMGBQdRYF6XpJSgfKiKRxJznI6MNW+ii0DF
FwrOWZbyKoujlTYGBuOjpzxjSWz4ilVfck8lmbCW2Ln7iB/xQ9zxL1hMXC4+tIZg
Kf7eSqwuL1l89GpqRNUt9v2L3kdj4g4tAMlZB8iSAF7K3KJqFR7xT87kqlITcb3g
DXcm/rIaYWm1zd4V+Ycsc5U7htDHy78YZhnmOs3lLgeij17IaTJMMUiPhAKoVOjo
RrIF2E8hB7gosKyqLWkJZhNNQmYHyyZuTTbi9K5gKR3y8SrUjN6kp73Eb+WMVhfJ
GyATGa7erazAn155tTCwAnhtVpouunGkGYVUoYFWGkFOxRrSl4uV2cWvD6VrPItS
0oKo9GaWhCOi816d8hmBN06axW79nhhhvBEjVfLFXvbOXmJeMTwQ8qXH/Ct1116l
6bqwg8l5FvuyfSgdh0V4iLH4RVNq/4uUAFHCG3EyvgZSgc8dynm5o5EfY/MIBL7O
Vp1MrwXIEpeZTr6bY7hOVD+akv5RQXveXyXP+jQ6BUS8ysiQu0dcTVC7zRg35gOA
dX/ICBKHzLd1hrmK7Em8wuCMzR5iFN73GXUetvnfNUNav1RA2n251jqvBeI2FQmP
OkNz5GU9LzHKP4WxjJZ/1ckY2zXi712+IK8kRv00eyu6xlR58LCxs9Fd5nkE4LyH
WU7mqxqLvQ73UnfbtdzV8Dw7g0G48FjtnLfnR/bFxV4=
//pragma protect end_data_block
//pragma protect digest_block
9ORQHBFYllO6+ORTe7kJR8ecnzA=
//pragma protect end_digest_block
//pragma protect end_protected
