// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
WdAJQnhv9Z7gqRIVtH5j2m5hSnkFhgQ6wQq/OXor1+ULTiqw3mhppP+p84GPPFYe
2zgAvNuDiA3QP3Hcnq7YSZ78zpyzMae8trNp+dmZq57XPEbFMiiUrjMGhTgUF5ub
+pRb536Qb+UP3bjHE5TXEDpE2K3iRyV+1SrcdKjXHN2Nm1E3jSi8Jg==
//pragma protect end_key_block
//pragma protect digest_block
ADzzOczPZB7Vk5jv4WpfCB7cdgw=
//pragma protect end_digest_block
//pragma protect data_block
YGyupO3lYRDlCmp1M7YLl41DcNV2du+1hoToYIRWH84KrgryUBnNc5z4jDhllpRF
CHlS6LinuQvak6biENxdg10W9WbhNM01+Cs/g+5lfD+a56o5RnCko9O399MjpjaX
NDjVnXUMgsTXiJUxFR6Syt4cQdTZMKIcpWb/bdOGRRWybo+cflt260zZxrv3aZUG
1ctJ4/g0Ip3beBrm5xbXlWubC3DllUfzbWTdzy8XkF6hOPZfigxmBiOWeExtW6Kj
t45Znwm6eZhoXkXYVhFnZSoAa6jmxp12vZDWLNizs0kqOR5WupWF6Z/lz2+Eo4xt
o8HqmEL/4COzDsFyD5Wsz63JF0rRVMfXKGULYCsXsbT6o1WifURFZlnIf01s7qGd
YZcOV8saANFgsOBt2YOJqRvuEm5//YiQ5uxtbkXCwx86ozBXp/HoVK/lVgsB0Gva
I0P4H8bZgrGA+/h8tprdPWYd9Reo2QlYcxVFxytc+SEgdUj1gU1OIj9ZlX3sI3e6
W/pRsYGIfMDjX7WQWkPsjFEkVWr4DhiUOu263XFmysC29zz4XVsM24O5gfqgfQBZ
qAthwmb1We31aund9viBoz5vAgcV5Th4FYmJ7xQQ1mDWvyO1oPNhkMv55iif1HFf
vQry3vL0ULQ1GjW1XF/k9/6u5wU7ms6581L9CBaFrzt3sKnf5d3Mt58qeC9vDJLu
MJEWytXMuDiDXAu+D3D1+v88WUlXlcnobKWuiVG5reil/l0OOt/1dd/w7t6vKvAY
42wVcpEYnpf5m+Ts9Tf0/JLLj9ucDyb/Abzx5NpcRcV1V3CamzmK1bCKMM9qYrZd
ISdHBcbxgpT77pd5eRvIKRBoxXctld7uDONoqSzrb0pI45RIilduaAsNeTx6OiSy
c+ydWqLaJZsXRmwMHruxeJqJlq2YrNmmJSjimu86xrYeUrCQIEyjUgd1v4jKWEV1
O5IhnhZMwKkcHctCdSKeFa0BrxU7Ax8FZRNlmSX4ehEkR+mWOTkNm95U9yVUTO+6
A0ks5FxVnVCLKJpT701rZwrCnWOjQadkgnAh/qLuwnkIzEMgxSpfYkfh7qqnb6Z1
fgfLIj3EDe8eB4dcph0Ox6OYkgXG0TnJO66aAKSz12ijBJJ16mZ4UA3pLGA83XAb
tID+e2l1TR9RqYw9guFpSjJy5lHuZa8Fk5rTp3kusExPDSkedzgHbV+3EYNopXPu
I1VzP5sDIbzfyzTv4izWrpECbsxGG5FnAN5TuZKiP3OdbLrXc1dFHELAKB8TqPaj
EpVlVVP8lY5ZwjmRt0ZXk/5Qq6TOa+YH6VwFHREwc87p6YTKBgBp34q618sYImzA
v1wcpsdMcHg2dt2DnPwr6vr5K168oi1biSps3CPeLHcYWSYvmGpdnnhsN8OPr2Gk
WDL0SvHXXrv1LPCwFt+tjZhmaYMIBUszXAqvV8WJmikYOESDc+P7tLUf9i+EPeWs
XWDwy3xKwDrFNwytC17KyLL9EYJg0Tmd9w9M6TTaWw2P4ZdDsAkCXcItLwB+vSUX
rLKOomJorqteM8bQH0T4WlKHJpRHgwjtvbfXlTEw3sPOTlqbh3/dfrV9Ka0xShkr
dEZeHL3UuaLeEjZLHjkLjyuQqk6jZ8695Lxu2ZRKOhmMRrlLb7LRMB4/PiJ1xfd5
X/DhPZHJaNYwYBKm/AkMRYfnPlXJ1+XZHAYDp/eCLjngaK5HLSPTIXvmW/hwdnqb
umC05cdLil2H8FMKmPsYJXscBesZyPKELdvndchoapLVHsWYyspAWGdRp/P7g++1
82RXChBgiA/uLryW2tIZnM9tf4nJJb4vEdaH/U3MV5JqJM5IpjGj2FKvMLmOgfFf
9tQwjT+WHRW2ds80G3QwzKZJx4wu2SrhMR/BvYFpx7rLe2Ffj97swqPL6d0nuTjK
OzFZzympQNE0OzBhlKt/p8r7rGF6GCpcHDUDeLVnZI4jeQKuojCvMcepxWT7tVhk
DIQL4u+Ifkdygzx1E3fkTL7qqlOSiT47H0GJ3lRU5xpoWqB0iZTHg7gmvbyLjHOO
ha5c7Fh8RXddYrUx6geXhj4rf6r+6kwP9dMuEUXdewggIZq0orgwYzim6eFkGAmA
scX3AdQiLzjDnm5D3umzEySbIiQHB9CK6yhjTBkbSGNK2ftzDO2Hi0yaAKdOTB1j
JcRrBz1tIl8/bIqpGWqG6tXG7+k726x3bZeruTL11eJK2tfzciTeWL2MOOfXc4p/
/3U4gvCdmzkf73r4iWczv57kPUtTluA+3vVVRuYLo37dWHox7voQzBkUmJalmQ6M
00rDIZDPwfXTAZ+YhXnPTlMaY9n9o1Y3BGuxbNhwtoh1hPopGBZiLXj/QuyZlcLC
sGpMmrUFhgUBtAIhXEJcRk5zPOpdQbS1mRKHwWNYmrxYOlONNuGxp8O/y96GekGC
GEYzWjD7qXqQaNw75Us3t4VWGMpsuy8stEZaxV20KLTEGeZlNnOedvPKCrwBNlGC
pYeoyp3JERTHxxZ91zlHlqcjAvpa9vMVLxVz/0d4MTRxINtqFLPQG1AbCcuqjr/B
/4/zX+t5fWv4mcKiodfDg70y4b72nScdtu5OKRJBQFTmOisUkpsDXjfNU+9ex9Nz
bY2IOjYch/sIfNnqBQHm3mvyInlAnt5Clptlz/5CJAy+M/9dYZcaoDVtUShgsiol
ybplh+8AEOL6qeQ7q02dWVbiKP8rLf4KcTMFH308edYJvMore2QV1vOv3248fnwM
GP2/RexiFFfozDEpizp6oTRoVXElnnX+BkqykIpVZRgDkaDWFdVvltgsm3XKBHSV
pszLuvTwXkqXKet+pIFuisJ7uFTIamO+K/AqZvib0C3XpjenoE59Os4Wn9Bs0tqL
rD17bcU0G8hBDmUewcZ9ZJaLWLrU7Rq3lvLMHcJVnX60Pp8Y7hAHn3nhIdZcHjAH
YfwNmvDvFk4XHz6TE+2i749dUMYbhT5F3WWeAnnU3VKC2Ir1GSSj6/8DCgUsyS28
StIWVpUvA4wr2kZSPI9R/Kp+roOA0di8zoBqZduQGe9eEZaIgnQ+Vg2Xh1q58Mh8
xLMQqXjL+C8zkwScYrz/m6lt38LEyQnwzPcRlqb6wWhcmwmNTvpJYoTROaguHOsD
R8cLqyJpcjsFvna4zwGlYcNQe85lcXpp/ar9/+c785fPxXtn+8ckTIcW0DVWjPjM
cvV2sWYl1thruBTUHNju/O0IHNMLooOehqO9hz3YTQcNcIiZmL6/OjeKc4eLJNyH
9IWgJ4aEq5gkfHJLdk9pOtJGEqIfljKHwOTN5yG4JtkUxX1ce7nmJIQ2e97LKjal
LoDG4hwBR2+m8DswVtIZaSzq/rD7Ybnx08O5eV+MsvxfiwQM9o1ogssCo/RCd4NZ
2TKyUmKae+Gr+bj+LrXg7LcBp0Ilgxwa66LoCNlJ1KDkpD8Mif5Wkf3WQRm/cNRM
9oIKlDEw/dAlfQK+6C5CLyfZPtG+S442ggA0YBLexuz5WnH9P6WTILO1NycWy1qq
kNJQ2uZDaONOp8Z4WgagjnxSfhJWyx0zJw6wf8IndfYGKDjrWSdaqRDe4ALM2E7t
kDvZ+kv6SzK0E27KBtHdkK2F/Pv7JTMr7RhVk+EfEj570oVQg1sp0Bo9fOIh9Glm
tOGT4aW8SzobNQCH7VVQRgX/YngQnT57H6cujnQ2tqJRt13rWUalHijK2hNNGQXi
SmlSSlGIkZys34JlwDOqHfqTP6D3cj3ZONyUBQ+tllTAhNvvSkMLApiSm/KECnu0
9nnlgxZe2LD5WObCTOoVISWPDNDGSFwZBcchQibMatrSlZWmdfuvkfRSWXfsdMcO
oWKp5a4o5D3ExHJVRctOeUfJ/AF7zMu3TJ+ycoLA9aEBPc+Zg9Hsq19DL6JzYqnt
wj+EkkEaRYtvttE0ThG7pQT/Zqi1mzY5cWbmdnqwBH6IeHhaNDdUtnom/ounCXJu
2jaOv5p1cjxYYQBoccrM44tOJkGMM3c7075dx3o/z5QFTlnQYUjHBATxWoYFGUVj
gLRcH4Ei9LmB6KpgISA1pfx4i66rZGaXbDuMgpSmWMwpxmNTkR18ihDSm/ccSVFe
sT0tVG2RVwAwcfuJsdFbRVAUq3LCXFZiYnmnTksQ6f9k/GeXsxc91YYqerhuLTts
l5UJh1qZ3C/nAcbi55A0M4QyapGCUgcp3TKUoHl+XMXGt5Iw9WUk3d26LGjtjcLZ
OSJ3q77dR6a9ldgEI8PdVJUDqkZ3Lv1wRRCyRKBneDIGP/DDViwK3VQdX9Fvts0Z
7qorbwRocxuUHhAZ1wENmtoUknYZlw++8nt0Val/38vwNCiLV8WN+r/pdIWeiagE
iYlhz9Xq5XENdH2qGYYSXCDaT+RVyMD0oFhwBO5feuCOrHM9AQCIE3Z2zEX4jr9l
b1BeqtOK+K2jHEO+LzEOeglu1YVxKhlXAjQ6ET1Jxnc5dzyfsIPUHjf6eiDDt26L
8xvRQlcD/yVlbePeHSxgfxlVwCiQdu4rTf6zV76AN0Vpizuv4cO6h+dzPrnfPmQC
U7KLxNzaLR1LSHA1+mx4Uomy0pXnVPbbXluZOgkupElpDXLNi8rKR2wUicvWOzoh
1zV++wrRF0N351RUn4Kms2bVnfxO+hmEhH8c7vE5G2754izNCqPPkQHEyteutDwR
QFoDHK8iBlzk6PtcjghRuqPKAv10JvakOIjM3EnXBiWdDqRF/McrKY2sXJKRMq3T
ZBk/P0Iwia/T4J40GIjtkiUtepGNvxDu1L5uKDZglt1GIU2SnhFFik6acLTeTNar
DaC0h+rh91KcW6Drzhk4Pov9ugv8iVEPgjMi2Vt7MS96wc7gT0jzQySU/EHeahQD
VbZ2nC0hVagZiEyOyRURHYcG+dWnPXO7SYjcevUw54IgvEmWtFYViPgPz3fLxw32
EpE0cu25Q8caX2QvPjc94EpLZ/VwCVR+GUKQjX/PjnMryDcfTzYQnqTP8k/K69Kt
6l4YfFkRg3hVzKNbYm2l+DEo5MMUUbZGDoHHf7F8pFgv4HeObVBHXf3QW5grWRvC
mORXBZf3jTIROtlw4P8NgLhTtaAPk0VjnVNmG9uT1Qym4HOJ5Xqh3220JIivVQB2
O0Qq8evEuEzHy7v53uxuJJfpI9Pyi34VbQ0yy96kNk3rf4iWo/5dbyeK3CP/Qrfe
mqG8q8yyfVYgXJih6ApbiILyvNin80ZcXDGziq481N1T2g/7aeOoNW2iz7avFxQ1
iUua6lZsp+taC2n26PRVqXtTHQncM1OO63p0p8mSh+aAzxm27wxau4lbYJUoLRxa
ve29q6V4dQRz3e/7bkc4tWpWaztslSfypb9qwFiC3UboAYYa9dSP6xy463Lrkvpb
X5vz0QyjJFSsSsuO3hqJ23yDr+IdBE3NvWfOYb4URqHVf+2cf2w8IecdyAOxtHxE
jhuFhwLXUphC4WSxLcHY4gMRR9mPU/cEf8mCPLcYsknkEz/DXuDisBDBlZFnZURR
id6blejOnC9mUyBVyskTrZSypGtGt/0R7r0iSUm7dDtycuDGDF8wSYW/v18gclUO
9m9PSJtJ/yBchjzoMbFaCwHhItrggTFzFC66xuKZYd5AJZ6bQeXsFMvnP+ME8VNE
aw4c4O0FsjAgcUM1FT0ivZQhmzvuIPJb6gZmp8p1gwVEVChx6TMQ5LV+Lwavl0gR
wsfG2weIkE2Z7SC5Q2MZu92HWfHfoNDTWUpu7qfMZC1Bn6pIKzLEz8yGYce1sWL4
fwQSt9UWY643rMX5xlxkCSN5tesbhQY1IY6VDYLwHBzfkiQynUhWlzQ01UKP/qIH
KYSW+sfZ8zmeqW0nkHiCKMFi9rAcUn64zm7G+jdskUHXolzjn8CMmdnEDxOim+PV
mhGknlL2lODH78B1yYXeQmzHg4pR0RfiFNO4vC/vwA0GKlqkwSDveWrYV6AVMOEX
zz08rjuksf74XTvPUi1mvfN45MR5xeLkGp74HVHQZ+rJv5yoqnFweeghJxLiPiD4
/99KVX0g2OYSzhHxkusb6YIE/ayJwulRJtOLEUNL9g+IWO8NdIJZmd6amJpXzUqr
bvhovDNDKWIl9gzkAh0aTylxLrnkTAsGDMy++2H5+V0gVF2oyE+N3WWs5EQl4j8m
EG1R4IDendGcxN7ejX+YdiC3hn4T7CySaFFUdEg8P7808+0M8Grsub510xk245JE
7TPTZ2QGPu+Pk/ZqOW6Cx5XTzfd3yuz1cFgDDTPYut6s/vtGWkh/o0gExngqg4gA
mbMQkC6b/0RjfEPSps/4erLSHu3ZGtLJfjRvBLQhdMDTV1lnyeO+4ROMqxlV/ogf
awlnX10/0BOPQMN/ogw98aaIXoKnoI+x7YZ11EAD6Ckpa6oJVS8JYeTLaG2uYCnR
Y23+MFdqLjgyCsSN5wE5IPoCWG9iW53THG+NyXCYe45ep5YgV5NxRakjaqZJUtYD
MsFLeV7xoMIHFtCuN9gSsalAZXEr/iCivZp0BjM0Atv3wIIM5USubP+T6c153PiN
7GIiPmG3yfZVcTDsA9zeMC+lQfOrCyPHAJOoncFZJsUiu4V642ZBqUCfBmtf7S2M
IbPJDtoUzgwXA84/loPUuOy1gYjH8cR0ybcnqq77vfC4wpf6kSCqhXITJuSfWLWM
dmCGR1tE29iASOOSoyTtLM4cGediQ3nduneiUbDNoZlIR2cYXQ+dnophcjmGa0nU
k1LE2dE87POkthwcVe5FZJhXAKvQo1mxOKv4V2djT9TH3IZZ2eJSavepDahiy5GQ
xLe4uglKGO3Am8UXh6ULxUiZYCD+0kh7JbVy0pCghCj2HoPTGzW4xgcQiTvsDShb
FIWRid+j37RlDgwQYzRCdMrIvEmGPpHVuIZKSUerECIR6SNtj+hzgWEDbk5zTT64
087DsUtqApixciNLck4LeN29yXydyYAsbhxxH3MhnpZUzn+O32gKbDpczLk4yMEX
bCuocjd/xqIzonk+qzmWlYm8bhKjpXkXwErphB7eK6Y7F+7G2KaKfnhTZ883zz5Y
RmAQs0w9KirMrQMfupLWizFE6zSQogi6wx8Kdu42VDhuZBp6ur0oKEcwLN3ARVPz
kpal8rcbE0WOTU2X0JCz4noTm16wk77Eb1/u2BKa+qXx98658woWOrqw7Lcjpye6
6S28oGV1NLL4+2ztZFDZODxqB3/6ouzwvEXJmqub8KayVysNlnhG6tvvF4Qxahi3
MfRp5z8g+i8jbLZfVqWOe1BilkZWKueSNEXbXIRvBlPaYg4/mjXw6oONrFceFQC7
n5MGDH/6fFliMcW94MBdVKRtSWD+dOgtLoS3Z3d+cGd5D5JMC4YOjIYN6yZ2KrQs
PLSOmttxUornFnuULI379HC2DYxmHO5Jhn2aojasXbm7KMTA4gVEGmQde5OH1bKw
27S1SSXfxS6WQ+gN3y7czmmCc/yVEtsBejtRHpfBJHOePxHDfZCskCJnC4gqvdw7
qPipvO4ZXIH2ebs8m6P0gPeZImyZN6RUU4S7hb/100Sek+Fqgqp2ro/5A7pwdI7Z
IDTKyK2iM7bYwkKI4b5U3F0npCLC/0GYS4mk/tZn4VVYtAqUkFm1B2ds8wVi+nWB
23+esMuOUOp+596M2tmh/jFfzpmSOEmMY/1QPQI/1jgemvQ3gVVWo5NOrD6wqzhh
gdy1bkt7zEipvdYnfLzFLhc8LSO0TtyX0+GrS8+5qDzXrRmYHjbKZlh3IG+fvurS
iZBLWiaqA2g/vsav/51U1gobangz7Y79w74yfczA5j6JoKT4mnYtde20Fo3ls90S
Eg6UegUVhemC51Z5VVkV0UzmzKx/+8yldwv8EkzgRvg+hWlLIAJAqLdX7YgDBmyw
b8fHD9BON9WcD45fpdgYfH8nQ18bjuexzNjUw3feSB2TTsW+OKFL3FWc6nyysZbo
63uyv9X7mCdymxuqI3cBBMCEvJbh9h3N47pUKxpCTZ84XVxdigBGpr0d5d/sWN58
Ca9dmcAOLZehGUP3rdfpM99zI6XaDhjJeoNE0S0SoC1klVWVPhuWeKra/sQjdLCD
88hRsw1D22uZbCrKaxijdrT/QCN03ZuzypQ0gbf/oFSqLhBpDaS6OUfUkW6hYFpL
C3Ytb0+9TG1h7/vnhM1OR3HgsUIv7dXYKejGrhFOuN+G6zB7UWGoEbUJEBeb70Ha
Ll/Sdkd16YT0yjOzR4O8r2YmsVB7kpuDQowdOERetBMm7RTG6wiqQkb2uI/3dDL6
FUOZsje4VOsqCWuYVAfTVUj03+/+HhUlI67+PNPjqDHndqeaXtxbxdlcm6VEg62j
q+UAGHG4dmsOJFoNNGNsKd+yv3JWYMpasMmFuPjxeBlL8Ln8M+35H/dS6YlqKo2U
3PHeFwiRNMSN/Zy0zDfPKfP5NGEQ7r4LfMRRIGDSCznZ2E2ayrckihhPvkOcCxhF
bmIPK1nP8jARf5EWbLwS4WQ1E9M4Df4rwgxRLLI71KkL34kxJMl6ku/DyT2S+YXT
Qa7nYIrpga6WTrYY6D78dQEfcrPyvl/u0ogi5VqHLBHFduOA6VyFtG+qwp/KYC4z
QL/fp3pNUset32UTypC4xQwJ3b5E+j41pxQ7DKEpvWkO5HcRWrgzzVhuJAAYN4kD
zM7an54gPUzOl91d1C9WBNGOWIR7sG1lBTTWQ1A+aOeDY1odXLiGKhj4ZWnSzGEw
J/6ThEQWzLfAdCiol1nxzbi12z0P82EfS7OW9iSmgCmWVSEss04+OJnzvx+SZi2A
cFikGI2bPAnv5ocBWvyFVaT/DFeto5b1w84+JUVmTMRL7U29i9aE4CrOXE1MMRgu
BPS0h+x6HBgvXLBXYquY1YWe6ys+J1sHPUeVk8JC9F04Rgw/YKgzb6317uTEP4TH
AWjdVAXOKHpQ+HXaSLG+OBnnfh0GgpVehQdiBgdmtemzImm9KH5eaudBqJZp1/dk
PLwyqRmH4FrmJjXBjeFt0xEWS+surgKhWynIVF/cqZtBATjheMR+nN7bQ4s6OS5O
jDFUa2J7FRG/1u9Hfznk4jwrZw3IPdvD20xjSfO1j9eQYD8+sSxa7L6dcDpUido/
7Ph4wDibxSDAh9FwgmYQaueDZznPoUXYkXUNWabmtdiD5DiFY/KeEBJu26IC5+ya
bVokIAvqlrK+8Tf/8jnAVsxiSRtOiC3s45rApCv4pz+JWzYH1XZZnAi72I4DYSAa
RQLxMwYVBGcrH2AdI0vnNWJWCF/mU3PWjvqqICfWWnvM4ED25d20QBvAraMBqqpT
FslxsG47+67N2sQh3BRwrxxLzuA8maLnT/s4AytQaJUSXccfWfzSzrAdhLkhMwOM
ghrHW0pJsc8BFPxswJVNAWERJZ6yBPm870MA/kyOPFnCdqOdbrOWIPmSFlPJARkR
F4tCxIPS1TbDMhqycT0eVE5XEVlj2mRXlbJwwspurZxSaiaJEWAJ8t0tO3xwpzJy
yKwoVkWUVt7QpAiBg545k4Ze5+Qy4p8MZHBgH6tBfJl9YVEn3z8QySyfDDlzBU1g
4mw0AQ20XZojB2FqljhQcBvpcm4G2yAVjJKM7MmDNhJIVZxMhJMF3IPloDM/9W87
ll2Gr3dZA/kvLeLO6aAfa51XQuWScsT7hNB/pYr5SBRsW6hmqvM4a7cn8bxVpjRZ
6JQTpYHQ+5DVj/XzDHkIztPkHGcSEWSoJkOKrpVsdxC6obMQLV/3CdYxi2BlIX4D
zuUZOassVqsEISFMNlRFq/rQwDtXzW+7aKGShE/vYUKRc1uedApn5prQIHuHswdQ
oprjRvSqKLBoTaxmV4h7r5Uvc73g5EubwTEylxZgym1nJU95f96SzuAW/vyL8UHb
reA4ncWDsxlN/mV5Xc0Xle9UWD0QSJ0bA3HV8NuXm6JMSwcAxEr+ldQujNm9sMRd
mKwJU9vtSnjOn5mJGZW0Ey1WX/LAl8ybm9N4/W9V98lQZv+vlakgce4JkuFnhix5
7oWAt/JAH8WuV4cZrnzeEb1CKM41xFSiwqt+kTiQsxofFZOwHPmhl03Rtdf/5nWn
L+Z6V6QiUg9i7phsXz4xcOx6uTRbhzV0vwVSflsRe1KRf52M1oNvKOh2I68nIh5T
/JKGfq2iW6Tc/Wvrty0V9IoV6lfEHNlMqYly95ITNLY4VQFPC0O3Komyfhqu+ulf
YDoKwz2dYYc/KXjgeNVM/0Ank1meNNXij+fWSjYW5SP44wefYh2tGah+60xgksFV
XRLwmBR8W57AoOu8AbtniQrC5wVCtJZPFzXSGb2atTBoepb5/5PpBgYI51y3qZbQ
GclyLlX9kLxbQNj4Vg3+Uhq0M3H8lYj2Wny16KvtVZe1midJduLsCvGX4JG88wqG
H1HVAyadBXbp0y2thp4BvIwrGFoQPOw2ojkAQr5xAPuZe6KXhIVgTiTCRZjif9vC
H6/NqCQKrVSOmgun8steMHscaCFEa/VH2j80t56FZYInRliU0/jbcqV9P28I0RnE
2CfWJayJ8/5Htw6BD5N5GBzO1nzVGgK3eiA957RwFWlIKZEfi8vPN1PArmjqwJg1
HqGGJ4AKKCjzW9W/8ldwG8kKLqHgKdsET5BTl3XDkmChNGTiLTMxbCAeEbzIBpJh
yTo9JbF5xHVfGRk5c7DBEhMUgZlrzelflOSoemja8cJU4TQg6I04e8E91Mw0/87J
OMBu3g4sZl8N/K2ErkmoFdEfdjF7y3diL9lPVeJkm3KovN7olwaqhibXdSJ4wi+3
LAvXt9GWhHzBsxrWA4lJhhyekRmokuyb2qkOeb0hQVHt9WfOSgxrXBZmBdezaJ8r
qlpNIGdGrGyX8QDp2dhK5s7Y6U6l9PQF0Dg0ceLpJ7RwZqyJUkS7kUg1TfVXHIa6
gD0jow0oj5bZqadqa4k7EA18htUD3tS6Z6ITMJwDDXA8szbY4xpjpQIi2ZBcnt/7
WyUDQZu+hGswX1LcTd791rk/be6i4JZLvGaapImWLf1B+qJknUmDQ9KW68O2ks3i
bbKPmf7bVyuTRwhMb4H8rtNA/bj2dkr4kpJ24emJL4G8jsAv6yxbKcgS4Vo5TJ3m
oaE4nlRSvGlxMkokAbPvnS85JcxATCQ6uvF0UVH4WEvzSgrVLiRb/BZAE8l6me44
LZtOwC/SF5mCreh/fPpJBhWsx3xjfvew1dK2WvKMJZwS/leE1F/OhJaLtlwsqi8d
WEQCrRltfNjPYcw3PYHjsNu7+6oxL9at0VjYdine6hs4hNo6NQVUoCp4TZTS9o5r
vhOxNRGvhrPBQGsMn8gQvgZFZY/1A8ykCOBlE6sMo3t6ZLuRtsLfADhWAXKUBTsd
+0MglzmngqgXrluZDwE46I+ujihgMQfi4b+lXZzVxnNj1aNFNkIveubzHBy8iS5y
regY7ORSxoZrNwz3Y0uMdqtum6OdmaGtpjgfO/VjtZ/KfxZGCFIFU8eConzmsxDD
DHkWsLYMxJwlaF+6Ch43bBzyWhMn2tDcbvR75x61zHFXPEIlksCaSlQmX4IcOaCz
ZqAuie6NsUODpHlMF9WNtTWrHox9Tjy+QMa3Q8uhUGJDSvZ2BlV2G3g64usUx4P+
QN/wwOXzCdN9yd4qfI5w7jqghPO7szoMOwD+hs/J3DNqDlYlZ92NDpDMm9rdK1uX
2j/kIFaQF+GSs17BbvhJDgRbSi06uHLndlHnSEBfO/k2UZ+jV7WFjc+Zrxw5F4Sp
Om6h2GalCASZgV3hlRxJV/mdcWpt1H7vffAjQgB0r6elSIDcAJnSMzgsh3TZKy5i
4vGtHaWIrvK5GEqpIzHVQZXWMvRpjPwhqeYz27uQS1Gi3M/1RpWiGDwsypOxH7eW
e+AMya2O5z3g72XBSN74EYpt/N2V7oekd2PeKlB9iRrOUPsojDmMNMKfHQFa7wOL
W3f+5TlQvalY1pf/hTlfkinhsEDk0WMLUUH1rI5fuxD9BCM71blyZXNjQijmVFNx
Igs6OXlzhfY3Kel19HE3dKdKiBbnk36YWmzrbDJrwumNFfjNJRp9sbxQi7SG1umY
3wtJZ64RztTYOgyQaw3d0xioII9jnKcZsKP8zp1jerZrCJg9qp01tPENbW3Esuwl
CIC2/XyVwAmt4ypdXP+4UcWnrjXdfgODYBFZaSgSJ/FMeIkIM/AXE9H0bpBOl5/K
CRoPbF7+yM4cKIEpGSh9yALX2wqJokg18eUgQAWDqWU9WV0GellWxEhCqcFSsDlR
vZyVE16UHEo5NekpBGq5wa5POAGKucXntrtkiTiNMIZCKzeoBc6J75CBEYPsyypz
w76e60YL5RaGo2gvT+BflQ9SFzyIV4gYOGgON4hArJtmTExGCWB/1FujKAQ5zuWn
c9lSFIehNlmOceOlI4eFOD8Mk/VgVxERY4K/ZbvzpG6uCA9fW2hmfe+yyMbLBygX
qF1Vxx72OoE3IB8fxxU7ggnlGC1P5nmw3WJxy8ncVBGy5/EkWwHVloEzTSYBhzaf
9CmeWOktxVIl1xo97bpyT6dHMGgccpavubB9//DZhkHLZbA9XMBCw360lQ0aoSP4
/w7b/l1B+1eVwILG5F7jiTYNFEb66jPrb0kzUkY59mWGqIE/33OTIKZ4QUUozZZn
gNDzMccM5Ye64Iv2k60tyz0EQC7m1el6y0KniGdjD08ne9jdJ32ZGWZ9l1xTVJw7
nqnie0n86xFY7oC+XqJ8dePSX2rxCjyUzbjx8FSWdvO6x5NjdXpIp4uaahJyxXAH
0nbBiuEgf/mh+/Th2Ivlya27YTSG7TNsAElXFi17PF9xac21hxqk/UJc6kqsRsNT
NY1KW0G/ryVFKZupfF6UZJ1dhTR+c8Mj3lvGyWcgc+Cov03FXUVVB2cYdF49K7ts
p6j8JKU3emHrLXi11EQrx4Vbjf5fV5wKRABeWTbbyGdTdD0s+gDYnh3sb881d5s0
ighCEVxBckNqd22q2gTgWS+6LKfNY8wgckUCiqRC6+DAEK5ZzJlQzpod2KORFZ0L
POQUABg0ZTaLyLNATs6CWLDHO5YRxIDu0i0N7acgmHPzg6A+6zLx9K1Yf6KwYfvt
qwV1Iuqq0tW2q5u7xDuplGa3EMWXmn0gPPx5FSbUrDoTItBPvBsyznxpqflznZVM
codaaAC6cuByJ5+dWbpovVdRwm/lQLB7VG5Ls8Pq9pLUQREn1zGEY45Mahnfm2VS
U/no4rFliPDrGXzbz4lhm9PSRW/tFsfuH3wDPGsUcldvWZUpu725yyvFyobhmTah
ov0tCcJ3IH//d1C+5+rYYlspJULjbsBGWRnHEN98nQT1Kpxol94NccdwdOuDp0tM
95rUVVew+usJ3fan3K93xh7IRnHe4GvpmdCvebzV8400t1YgvgetHmvgmBLettyB
C1bxdrSOKjLt83juKomZEutV8FfpgfhYVahcdbTMv2dZPdLogkYVHP94SZYmQJKm
GE0/YWqFofR336WIQeb/U8UtcZ3WsiZKVstEO9LbTh02cLC5gEJkOMS0Fou1BYs7
O1Jl0x9cHZ+HHY7GwjSy2tJzzc5Phka/cfXiSZrg006wB51ynW5jrd4ZoqAQ4u9Q
ACmyBljadr5rc7kx/Y9K/ojYH8dJSnCjldyk46dnkr35uNvquWU/bnQUcAA2jXVU
oKzegTTAJZolhwD/te14sEnlcs2kJu7jWoxx75HLQKqjhZKnCj96gHCXQMuUuZeL
AxCegUOYjXOnE2NiVVv0k6faCjjcvF//JrJyGrOeMqiOttyU6fmWDbxMonBJq9iV
6+ollfVOi7tVCsAWQLatyX6SJELnVcMu2LKegyK7AmEryI/o02n8gabOtw2YbL08
BuqJqbQa7jwRYX16Ri0P9yCHapD2J2P4FRsvPnxIzP8iuL3I2xlnoh6uIPXxARjp
7X1LwoaKFOwVGmbylLgIZWAlI2qM5cf+MwMEizRbn0QBxZlpCh4LM26/kMp54l6p
lLh4u8WVTxHE/NqoVxxzhZxp8u/EQnDHB5Q1h+vbJwohiQNUIoZp0QkvihvgS8d0
wckWu/SBXqqG9lC+5WNxrRZiGFDLIxodvh3dwfproGQw06q9+d1HjsgmcPDBjQJU
GT+61yMtnPIm4QpQz7sQjVVYsMu1XQRYgtzBNbA8ekpVXWJVwDEnoBZuTnbVmCD0
IPXp0FgqdXCBzuJAu08e/HlTftr5Q2lzhnjhAuKFlZUOE4pakKjDcx1vO2OlEY9A
yVNaFZPq4yTPd0iO+l6JgjabXWj50xbKzqi+GQ8bYSYCM8wM+C+lk7Fl0pyJMcNY
5WClJrKV76LH589sfvS6/2cmDXjtGAqXkIUI84hqPxezYUoXlEEmPWjYaQUisWFZ
Lud5hEIPNOkJ8q6z+upslM50oFjBLPxUf981CbvAy++AFPIY0nvdOPWCwvcWOuRe
QTvO9UN9DLISZ1+UH6GqLI9JbjUcmQ0fgkAget4vJO6FEbBmtnWPTQ0zyVrXFLin
25UFghwbSXM1K2fFtHs2QAvmfdg3UHkSsoV+xe8+7qav5NGnItMELxwMC2ZVugdG
Goe15KTLRByQNNTqgXFYDo5YuZDCU+CQ6n2eEgllADMO+Dca4OCS4hWqOGACMiVz
jn8oQu3p6vTxrT5Vprl723UjU2eYIo8y9gz/QxOpvzgDRv8JVCHobzLHgLolLXIX
1UShl6+Ygbd+j8pbucuYVyq7Dgg6q3w6iPHPdckBCf3Oz/wIT7uQ+NH/doDmblfW
ki5wuemJhSZmCcX7flMkAYnhZ/NeuH2RE1+VNNlP05ZnqxobiBjCbqUbWsNeYsQg
0T2E1VInxIkXcQ8jhOYGNk04Z7Ml7k+A7Yqt7QEzh9v7gJ9TTL946lo5HC9naUMl
CAGeQ8znb3AwyhGQeE7DJ8cQcuyFKo5Amn81Pl+McWN5pS7Hki8eWLORc9UPzEEm
aII2CbrnfWkSx2Z5BRFeMyfUhjh10qGXiDO8sAub22W33xdAYXa97HJVJN3UwfNU
FKwTIWucmSslVtuiuHKe+HAD+OPhpmTxwVARd9VHdPi7bTf6dawGsyiwm7T3fw/Z
fxGulG9SY9pj+eT4C3LSbCptHZfUv5vfhs1AjR6KUT5LVWzjkk5ikeyjjwXAtakl
k2pB5u91otcR4k6cY911q700sDnKilJcmkXbKFkuTX50iZBtTgfQJj7I8MdoahYS
6kqDIJlVtu3H6hG7RpBVD7stToPbhkqXCvTU+WcErXmOdwVXDlhx29Khr+h9R8Wj
EmXO8GjMueGBnasc2Is9mbHkX9ljaLJDxZs0uEm6tDFHyJ9QcMp8pTieWYKoQ597
fbVgLkuTAWoYH/PpfFbqDV3nfjCnMApTNN2yAyaJ32uMPS10abuhU1ZoveKi/tp7
baDsVPZ4PYXgfXT4exl9UQjSKm2hTRMLpcqBKoF86Y9ax+SPfAuobfTpQse2Un/E
EPLP/CwNPVIsyJt/PlyJxfg7dqI5jmFqIsGGb3dLrlbIpLiGVqAZpKN7BxRwjTzL
uNOgnTFG0uN8CXYKcxxeTtSFjoNoRUiaqkfLPZ8n4H8vxiOwIeCrAIRSjfGWMkJ0
MFffOCg7r4iZW2brTGecJQpI+zkNv4vhN1oH07i9Nb3gzvmjS+DmWZnlifaogMHF
+uh+CKr1g4UIyCIF7MDYbuxYpfQ9wq4mLDXuI+TE2tHixvaSUrgQldFobYXxiuDd
hToHWpwvksEyCZ/gcX+ula9XYDBMMquQBSAP3OwQMHRolRrI8OeFtW53LGgdcdwu
KOf3H2t5QLY7kB0oorYYzhaIxGliiYAIFyI2vROyji54jtbIPFwOprYGdPNCuwEP
7H1HQngLgDE0U8Xuaf1yozR8pwBHrQOIgMxJwAn2BVZMkiYnXpjM8Ij7yeRTZg+q
Y/NUGtnGf6jag25tkhD+7Izb/Bt6RBRRUx/0THlno+usnx4fg8SLo2i5R9dWQiVH
FnZcEcoU3FvsmlYxdI9v8uEzJw1HRbCxpNllW7fUDcJp8dSuCfcepflA8818wXG0
dpmceKe5pldyPEGgkqVrJ7pwEuKqJ2yvSDTnxRruC0uwzXnNkxPm3WOBF/dtegDt
ubmmIgW8+F0AwmDNevIyOUZjbw5vFBC9IVZBCd7veNpVtOMIc3rZfIYiCBYrpln3
39jPUZe18mW5AyqRxleAkxQvt3wA0Ou3mNmcXhJ1xMvhplhwwp5Zm2vhnU5ZBt8V
n5pCHQFKbre9Lt9AmaTwmJgsHuLLYwJ5ua1WsmUNNLhE7mUYUS3e+e+sck5YFjb1
sxNlqGL8XVztwRJ4FxCaStnqMizN8dHcrXCwu/R/lePsjVjRxW2XN7AvzV+oPGmZ
WfXmEcPntk9IpxFDfCdvybAyrxVQQ+kBtKnXFsW+2TL8Bp0w3jMvnQvxQnh5BvSJ
bFMwAFupMqEoptxQoUvNh2B/SGVCEHB0Jk07wK0nZTVuiU+tA35M70PP1IZDoRvb
pUx1VUpDskMEYeNeuSJZgkdZR3bLSsNqrCDghXytrkkAznCF10WxzfdM0yfDbAjK
5xLWY5P9nj6AUgPFKAbmlK+Scfk2qJeouXpqh8iulqnIuqvgllMLtRO2sShvng2r
dkAOtx82Rl/RgOwrZ093ZGPsdVEJoLP1in8+9z1HD25K1hhSFBDTwn+55H7uhi/M
poSV+3bsPF6kQhNrrKM3XVzQy97FJSlIJmAQtBgXyk4XeSXr2Q9MgGOoRulqyTRR
McdAaktW/m37ZBzvwSDLpp4pNwMjoELEzNREeGrlLWtCJas98hx4MFUM+qrFR3zZ
TqyAGE2lVxeDIBNb2V6DD9GxafkZuDGkA2YWT8AWMG2KkkZMjb0L1DEUAHDpnK+w
J6UHi5NwNv7QqJ4ElfR6/MYEII1ozB8xGeSWltVkenVzoM2oSDxHVwesDfBFxXcF
YX6LfzXGDfpeZEq36CP12Us11Yh4FJMSCwv8emRdQs1KWeubBBtg8iayFlp2mfMp
HCksX53E9WoNHv6j8lcf4uTi4MckbMftQZZh5tJxHJouT4Okg4WbZf2NaE/HGhg9
fafGhYUnBrKONFc9vCgFEolKpvPshIMZw2CB9VxfuW7uGgqkXeaWQKxioj2phy5t
Ojp2pl7PPiDfJdSU9tesirZELZGIfL+q4D8eA8khJ4JltN761XimrGxAfrC2H/wk
BC8U8viovMIJ9drV8tZK+ua6/bm0ShSBonmAbrkrlz3MbLCMF94f2bD6FVLUYbXu
8aqENliM4Xx0Gq9NkGZgMSVY0l+mz01cV04B6gb1D85TIhK3AYgxstRutXROnri1
JDfmPgl06ANBMqMLt78GYmTNySJP2rZdu0WUOzGfSHD38GvYfmlexqDg72v3Crfq
nrgG988Jl+RjtOdetuUGV4mdewE2w6U6va8yl/FT81EgUZ7ePYUVFN8E3Bdorp5d
lov9F2sZOc4U3nfvmC3TqDw4sVdYXMnamsjsEfmxnUeQ9vEuGzV6zf3goc2M1ZFq
5+HrjBaa0aZpW8Vw8DzPQU3bOIqZCOgvLZiUcpsSF1/NpL1uyHm/x5nnyPoACC+J
rnUCRPis+0dZZoBMkp18GvbiGycDaFBdaG0rIU67WlmLZdQvCoPktI8ZfEgUQ22I
AKp3q0rnvi8wEVnBofvoXcMYiLR7eFEWQGlVYIAbIEsc6ns4gQt2bJDEmX32lSxJ
lDaoybCmeBVEDtbGXYUUFfJFNo4ikkv1aF2ZX01Q50oNUtOdBMAx2wVV3ibBJRdD
wR30oTT+RPm4iM1HkGGDLM1GD1M0duRbtC2C2J+LiUp/4UVoL5aHAG0n81m2zwsa
499ZldanQ8Yx6TbBgtK8BBOUsZM5+yyYwE8E2c3AAfUYDd/u1yEiEUmr0cDcANKJ
WwyTLxDS68k1mvYTExK6CubqvhRZ0mpZa6xR5yqiH++rWG3W3w4kXz1UQn8CaqiK
fw02DKzpldXD0TZ2M6fRk876r94bQwEXhATkflvzSzhDxnQAF7j0emsyVgEIo/uT
qI2ntX2rShuNScpg2S3+LbLMmVeLKFa/iYK8RwXI1gGuat6vy77zYuf/VvzpXLpa
e5vXvxZy+iP+OOGEa/kKfSSPr60X3uBYQE0/uIyDMbZ7Xei+hYggkloGE8Od7IXf
qd95YEkXUK88r7bMRLCZ6kCW0jPwqXcnKLje2pGHoeyTg5nCD552ZI6j+R3XcPdv
rBl50z9Ayh8HUSBQDwAVKERdEjsdTGeixwOGYSGSD40mhAaC7IClhkgVVK5hGVN0
N/eLtqe/IsJUdcxVKyVGG6RxA3BmxicwCWX09ADCZcCAhaQRD4DF2g47l6xlkyWk
VQJUxuIA3BAYgdJFOc7oxBDpCKYm3WkUl4yVY7xB72RgxObril0LKwTg3LxSkdXg
pT0qn6vq4Rwx0Ri+j2z219g/DWN/7tKP0ui0WqbsnsyIehHKLX1vAeTFUlH6Seb1
aRqT4SwajfHXC9T/Sf+0g92vxIvYTT8H/2TWFPhkgQQeRbisdsoVtDTqITPVeAdP
sf8NqdHWWI5X3xwIrpsVtOpEYJnd7GmF0KjS677WHFC3jx63UQnt9QNqciMb/n5S
z23K2JPSMr4H/sb1hV+oyb33cp2uHwUy6H9BJq7c5HLQ6/2pjjvRMT/SeSufxV6K
JctIN/VHPGwRXMCMJZfyRWaOspqvP2HtOR2YY7kVGUPdJnYjrX3PR1T8FW1o4yBf
TrqjiLmxpgQePXBuBdi4CbfPVopyUA+xrh9cVcXhBW30/hZ8MpzCg/XOHHDdiQyU
jzTgWd6CAf3GHwmGAEql+aQ7ZpxC5grLgr4i5wcpdpyJ4IZZk4jBklZ3wudOLbFZ
7QghUCHe2rnCmnpF2HmS87aYDufoqw6JjAJ1S3XtOq8bwLgPDJ7xTtgt6MKQm790
CFSAGDKn+YnA64K+4rg2kjo3uViI5DpumZ31e4s5FKru5RcRwTyusQOvNk1r/T9p
g0ciyd7goN3jBBLVI0L3J4s2atXBP9HLbZLULja7EEFf3weCs1T58qtkoHdR+fTq
yBHfnGymWWNIYXbb/NEbqhU0svA8pa0y72S2x1vowGOeKqj6WpTzwHI+vU0Myi8d
nLzhiykdEZ3q4UuQcbDMI65YG+IkSy7LdUitW+t3C2DnrqHjBQL4w8gBgJLTZcpG
MDLXjGSOnJNAzEGZS9rctQ3E2nDi3sH/iuj5GXf/1dcJTNg3EQKksAv7cdT3n8ry
qR2GZyzMhVOpVSpIyOFXwjbFy8rdaNFlKTI6zH5AlIpKtIcR4udIe6j7rtaPHis3
9QO5uBCq8d2wYOXVU9C/HKWlU+T0BdQSuOo02KC8bmcFdKGpzS9ekzq6PzaYtE4G
T4DJ6yYop9x4xgHX6mC9O7gJedEpcUCHo9I8qsaoJjK6vZlZgvIgOWbcT1/PpQUK
Lat6/4tZSgcAlex5ClQIgQlssPxEr/9iOSsDeId6q0AlnnOrUavunPKw1Od917EP
VsAGl8sefFyr0vfOl9sF6okchZQwxjYqdP2gZJwB8FHeqMDM7iR4tQEhu4nyVG/R
+aBknx1+mFvKhGZ6k9Z9HPZbSgjF/p7s3nlOVC6hGr8qwZg+lcZawONXKwc/YtOp
5Nt4zGP55I3ruwK4ohFj4cxBsLA0GQRno7tXsLxwInQcgnwT27gqboQCuCKmAaZk
ba9x2tNEF+WvTi5TQVZZmpg0V46PeIj0vN+w9drwNp+D1wCEo93LgB6QTRlc18+o
svKJyuB064NEmJaGx5CUHH8YHKtSz35bQu7D2Mwc74Vv60T0TzkjA3WlamG+o7NM
1ZvO7ADf0yc+s+LxJ6ZcKcQ32aKoXzPVQYUE0+CDXt4XXqRr8NyTFFPwZttOHVkX
WpTCVItz19fzZsaS1R3SRucRn2MIWEwJ/Qvwyz1QTiJM2E1pBr6FMRisdmK05vb3
zeHkJoJRJgAFpdOKpkyjjAXU2QFfUt/tNHlJYpHaL14u88scRxlVLInuy7UqnjX0
+GCPuLJyn56zJQOTo8yubBl1J/SaW9a9FpuoWc1F5wTLFrs/kHX4TPR8XosyJ1o5
xF9119hYga7y2oPRwNyTy8cn7RJAB2Np3v/yeQ+ooX2UEjZO9zQi1y0BLDU7/V9R
QEByg+tEyaHxvkYPS1Dokc5SYbywMPl5wVoXVrbl0745KjKXV+ArvfNdHkHVzkoI
dtOVi4t+TJF5s1HvjGRvezJXKtA9WxGFuurFqc2a8nF7kwD01nhn8EBSBYxO6u2K
/BWw2OoCb0iWYS6cp+5c2VCHempF536j09hhFCtxQWoD8FIqwpi31vd4cEJI7UK4
K+Uhw/6bNoozcjZYL4SASOv9yIMu/2quXL08v5vJ06O/Nk/mt+RuJEVWoIbPSy0I
dt9ku+XSSxFljMk/PHchcU9wVKmd4acUx75CVkT9xFKo5kuk/w6ylMSlBRxNnh9l
rOYF4gpbpUM+ujLm9c+rJEZVdSgorcBhwQu+PuVLZPqQX7kBpFdHDr1Eltwjr0e9
HDWu2OUNSBZnduXZIBivNwOzSwTDEP/DXkfWggRQLyEEmzNbISNO2hSlVJVpYkqv
IqTyLpujzX6rH4i7aJt5utuvhMthOUgnKFj0hHXLt+CHxkT52ECk02R9ghQcjBf1
ORj32cs+NLJ0juTWHnm8IYfYK1w52zChLzyp8JJTDYvowjWj6V5bz3+qNn+vaYKC
OSs18DTLBqTD7efnwgUc9/kv4g4fT6j4HM3HPhil4Ls66GS8VKFS9cgIlCiOHJQ/
Vd/1cZcX9ejVxcFPUBnzKYazSDZXQ074aZ1Q2Ds9mUWDwpkHVIlBWFUsqAl1GwBz
1JBwJU5hDMeeyWrP7TrfbvmbE/nOLGCASC2+ZQH8ZJb1naq4F/79tYG/8QsOlzpw
VJCM9zlUdPnQoixSI4jI9zTf02zAncTQmckxEg3ivnwTBPi0exiuvTwzj0a91gcr
ZZJLg2jKythvyUBGd0Q8wV2ZUOdk5ioHZymlJKq9LvcKhpGeogO3zCAmqChXrK2+
Sao2FK3mHQAQKescQbvtXiscEKFA/z4n+b3Xg8OXR0XwGmIqOq7rmSEsIGLclvdt
0kW0n6CAcPhF0+oXi0INtjnxSqNaYuLR9Fk0115A8hWuMVBd0NNnR6a61inA7SBM
UZyL9Fk0LpGakqXVQZKqrp2CAzAF9Udp01plCZgmJFvUd0UguPhHV/zNO7LxpqHm
SyBg9PSpbh6Ju5J45JV/GtqMx2sPf9X7pvl5gsQjvvKwLik0RF3M0kn0P1eiwEOB
cPZdehza6IDi/atctquiRZgyaWYpz93/Q1s1JQEYV/V4zXpcQSXx2dlc/62uQ6yL
s31+hD+OE9u2Ytqv44aR0q3Bx0gJPxqD4H3VM/VVN9UugG0g2qoF/hG6TutnnQwl
wF2KSV5J0DtWlOkfEbDCX8yebnA4YqkSCyyYHYCgFWGcGI2juTzyiHxOtG1hFm27
dUwaI6qLDp9Nt3Aw+od47slvK7kXPb2PoGIgG+KGoVW2uUfRKnQZtRBIjnrpCJC/
BDLRYxfVKyuNEmGJnIDuwq8YV9N3/Am4SCWf4/RFiLoZUawu+g9tC5A2JmvqqC+f
A6L5jbYJo2gX7oKR/JT99Ww7DdIiTY+lKxAmOz5p9M3Kuy3OcsNWrTBL3JjP1vvX
U6FhZAzkuDbLaW2DEJfVNDTk/vap/bRl+SYhIgPDusiAiI9eQJIoDqil+mVb+2XZ
mAFcktfUr/8I+n9h2ouLerNxlF30f/CaAJZvVWtpW5dws+TZoZqS8xMv2dks4+M5
FcOqJ5Ed532PRRVG5OG4hSE8zr3xx5Y95H01mSGHpzlWsh8+LsPlN+l5bi5kk8dn
uSO1GCQpiUpDNbRxyw8iESRUmH/v2Tp7/gtxNIJkxWcTibxch+fV/BnPdAyYh2L3
ofFyotNw7GLGVY7cYjc+0fOerSAjua54yVf0SsgKxvhb6TxC1dyukerx7Er2kyTd
A1Y4m36TbbW/6nsJrEaB7NMiX9Kv/jfMC6NxOO5NWt2FPlmPxEptO/tHPzjsr0Da
mjN/rpPpoUCD92AQcQYllwl39GiNGvPAhYev13Cf9wCYSKlm8Wm12bvthWjLaYg/
holnErCuAZY8nLJTyXmCTbRDMCX35WWKoZm+X+nbi8Z2qGnQ606ozrOhFdEX7hBg
BUSa7W9HMUNu7Ix/THuCbY/KV0z4fGuRPfuuNCmFchfRxadMHmQiNkHYGGxUjZSi
ZEeU0/iLZJnvRaZQndW/qZbPHJbPy/KZhTz4F6Yn3v3BVxq9voWmyuWm+OHJBBZ9
Gr+J2tz9KZ8AxNcn2+pcz/eR5vnr/+IsobS1W3nuw5Jk1Ibo6x8teDO+erG9DEW7
7EaoojVWzNQwhn2T+8DQqLoC6mvAKoKh1cWWiOeJHN4JMrQE8/Si/7K47EPSNhqw
IPTcwROVNkHPwg8MBxh4NsXOWHLDEoA8XftlhqQeESZ6JeOh/GU7CYuKT1F4pDLI
eHu8DmJwR3x9jdIDqggxLct+WRaHYFFPIWLES4s1SnZv+0NB5O7rAp15EGEgV+zE
jjawjfiObsAu+pi7fEyP2tbn560DQ8l0CMtCOWGAYqEr0eFEpuVZhBdDky72UpDH
kScHczeHeYXzdznyE4qhwdeRwbgLow6DopT37UuksIAnXIF1nWt9JBuzi/bvzcAg
AHD1fxwckeIL2Qb0iw8OoznrzJ7Gq90HxX0IMZH/nFzuq+CE83Px+EVeqA3SmWwj
dtD2jk1yrI3Cc45prcN0NeYdmBODFifB+cYFrerm0cDaoRhpKcMGTp48UlKN4KOl
9fyV/R7vKN8nuQHUDEEJdXThwaoaACZyrx3rrjxSh446i7l03fjjQCn6liZn+eVX
0B/mm7jmEAOWZ7NV5bNRfE4QJ2aXioG0n0KdEr4Ak4IhIizlizEOd3b14h43UyXe
5ForXarAjOqbHaGsAQ7IiHV47b/3lKz3tWQAqxhO0IK2T/Hv8fuV4l6gjY9k0/+e
H3A5jC0EQW3tdqR7AY0oZrW4MeCN1yzUhjVC8b3V4zzbx4UkjoHx3+cNYWL0gRWS
lHhRDk8hSTtWXrVO4RI/ejnH0Ipu7LrqkqFf56fekQE7yZtZShvhaiRE4tGLp8lj
uF5UIRi1g3iRrCliHsoiIh50P2jBn2ciJMBv+lzWzTlBSlhGVF7zu65UWbrzJ0Qz
CFSwWZbmHQc2hTR0+DiXu7bjS0K5JI0NlGU34oi0Oot3ZQb5Xt3yhPG0prjOyTvQ
RLYhHzu+z8ANHvhBCFHm2E0gQGzvtQIJp9+Jjp8YD5QN6QIbuRRnQgIQbEVMlJj5
ZFUrm4JHzmrJxMKI+abKXUkqsEOPM58Ky0J3g2Zu1OdaZHhu7ZlS4Yvx1hkijd8r
75fLnUVvSpkwa7XjBw1delR0vv1dxNKiboojrAqBR+K7gXNDvZZkRD+d50sIIDmG
ErbvCt+VSMJQQ3YiagoHm8zvntDr7xPO0en8vQv/0sEwvpjfXcKVx+DXy4oL9pxw
I3+XLd7iotM74EiZNu6xWPmK4DzQJdgy/+NYLrSqHM9BEhx/+avr7bfOm+L1Urgc
xS01Mx8+7znDgNBx2kwxjw8brFIB2ThyVxibvnJ/xP5+I9y8wd9IDk9p3KrKowHd
elxgXIJiwbWezbfKvTdOSDcaGzBqeFo/9H6tJxwjhWTWpPcSHb9k9Pz+i6Ll4uef
MnVvM5F1vb99HLBy3ifLwVQHKZIc77MqLudRDAH8M3/sngTtrjXbV9kCmFcbSrnc
ibh3q03kl6NTEzI7nypnF4G0gmDM3PuAH8aJdGgmVF4ssBycYXz2ZAIYPBX+DKj0
5W7D+Hzv4ysvnfv9+3vpN6l4nJmk69EWwm1PULXKJ3PGT31GUyhPrSFEVZp7fxI8
dI70r957wzu3PpuyOPslMnywkXcCLWjTVbpb/Hmr1MORDCmGJ9xpGqiwVDtgLu5Y
tbM+Vz1phgycU+vombqP3G6tInyT1lLGkH4SIshCApoM+bt7bJnAGZQMvoZZ+yC7
XsbWbntK6SVQC1y9ilsNoZrDWGbGCyRMzPyqIBJ91H0dcrv3+AISu9/jLS7yESdl
++0li9bk5d7kIcQp//dneut3P6lpCA5HbFQ4fFyLR+shuc6OIONTVhFV3CVLCYmL
XpNfoR5HlJTgV7PJnOy79Vk2BQmzcSCnIwj5InCig+PUVE/Fh9UqJJ3AkaMFjrlZ
bwZ37tLNgp8ciyDvh0sy6guA3yXabpTxiHyDaPiYhbhs8W2IIEEn7JH7VWRUtm9r
nvVPymzhEftF8E4AGT02p0m+Btk5Ibc0Y1rP9HP9aolB9X56NU3OkwAQKnpZECED
rUESnDG9vLkkJH7sNkmlrXTjSPrMoXIRvVrG/QTLRNh5vpNUSX7zCEvJBRSd7wXa
wCaN5W7+Vbcl3NqHNeGUltw+lsXFzOKzTUXfTocI4S/oBe4gEhoKjFIVav66ppIC
fxzP1jUq7Sjgs+Yo5cll5/3rLW8Xjg+C8t7npl1MVOxgOr9Y+h4Bw4XG9y0uGY/m
RJ6q1FoNQa3j0B0P+eK7hyWHQ1iQL+NQKDasX03+JGzGj8tQz4zDmghyOLYBGjpJ
Cf4GWkDTAyIQ62qQ80jgebmV/bDf9C65RMPJB+OygQATx58hu47MHmR4az/96uum
ACl2AbCN+YyalSdxAFxCEz+qSF9ZQxf1/eEQeF0wdogx1w4NcbaRuk08BAfjjQtb
KqPFnuWZ7vnS55eV0jbTfqUcS6c+WqbxQ1g6Llnp96AXOvNIk3adls3ApSpX1rYW
1LZvzS+9c3hB8KWePa1uk9sgqPLhCrztR2eT/s/MQBP+Q7BykNqL82+sEypc6uX5
YEtizZJaK/2DPxu2hF6ijkqkFBAmQ5BkjvfdilVmUtQ6lNJbuu/4IORjhGdg+20f
KF4gcZa3cZrpt0L8Al41dhAI4jQZJZTRqh6o/ocVWA+Gly/fjkAlOovvVT79RZ1p
mg+YhjWz70Lu2w6U+7GWJ5Dny1GaK3WDpEbl5J5s21VVc+gNXAjADhTLWPgpp105
XtCzsmYnWVML1QCc6AxPGqwevJrWxye9R8qdzpUazzpOktlheaZ5nEm6d13N3mKJ
jxYxRDgZ5yhM28HpdhoMnC0gBy6Q81fV1faKOW1Cf4FAbkJJQotBBqph0jmYZ3xX
hg7OR8LkisvR87jNqtuENYc3xnlbk47nQpdLPM9/HnJqx9fZTxoMXT7K4a+v/r6s
oQ6xKO+DNFu06xAMvvrm6lTPEfqx+HIFYjcXIHngSFzjicWmjvW2E1Z83ULfQ0rD
/+2bC4maWZV/ZaUd87bzBlGwG/pEFpjCDll1IHtDbhBM8y3n8DQP9rehBZN3tYBz
9653ywDpZY9qs13nbC0RcXnFhbu7c7Ar3z05m6SnhdD8AdFJlGmW6Mr+uhiQhb6Y
at2IYvXhVRgIxBTqhsCs4xK8lMvQzH7v0EjnNUYD5PvaHNgjLMGsq5WPozr4cRij
I2e5N4DE4jtDbAZqD4d7FnoEc4QxuZ4uEkCN1uGWUJ5c7BRkVIg91OYqqBkKfLZG
rcap27yZmQtgUCbql3NfOk56bFzvrRsLpbBo2i/QFV0BhoGWgr+Hr9eqzL5rs6JR
6dPh/Q1hODHKK8O+WSsEvFYXCv9ibWCOBArf8TjyykaQzhbXfk/zhRhmdsLEHTLc
Fc/aeLRjJProzHtM2Owfp9qqnPB/qO5UiRT2xUXVK2k3dmjwUTl6314Ymy/Jb8eS
xU4alc3qp2EclEy3lTvNo/7Jrb4cCHIshgtMsuTrG44IL0eQ9z9xJc6XqsQvBWo/
6tIEozS8MdgXFNH0joDwqQ14zwjhms7jvnayUQwgEdYor14CBU0sYCU2i989LdXf
yemjVoStZJUMGqzAeWJwNN5l+jMf/DM4rqmVTW2Oq/DaYlPwVawVL7NQnS76JFYs
lYBDu13gu//eO7sdoqdsqHis8t9+nvTIhWpjyal5gVNckh42j1JnCoF/cYK9Uv4g
FWs9l2EW2PDSBESLhvh/+EkjivdCr3nxzDH/90CStTFGckScu8QUDqipNDmoT2Ux
mH5I/eGv5zDPJkeGgSjoqQtVwojEE5Pv1Uyenppxp326RjFCoAy54KBIBTPPMm92
PMoOPDXHOSJhtzpPDizM7xK80m96a2zMwrIWHwd3YuZB+zHQfcayvqipixl0rq9y
rv7yZxDxl0XSG8TxsvflPGua1SF6UxhmyVsFYYnRFsnsdDpG/GsQ8jhD3ssywpzh
2xgWKxr44EI29n9gPfaOAqkijrp9oCJyChkZaoimjfEltIVkUTi6ZMz7uUzhUlHZ
SqXcsZFOfsJyrcgGBNMN0xydoHTVNN3UTIn0kglHTfOzvSSXusNPKiueCBkWobm5
tyFnHbr8nfmL98tQfh50VvKdwnFJfj6bGocSOgqnRaS824Bq4hLKbwJYXEalmv78
ruZPzGnibdCs+hEBvN3GD9ILTYf/pZWfXuz1sIwP3HHtTEWdgUkPnW9a1JWJv8JI
4yu4SXMsix5PGR5/vGuftikmA/oDWWMJs7DUw+gYAVWL7LEBF1eFV8Elug7eQAZl
oGgJrj0FSCaUJWVTPBYqSlaPzdyGrscX0DCc3bDVGGWZKlPm+gDvxbVWe0yFLLSm
7mgFaOycS1WKmwVL7IiAYtGUgDcCAop7VlSrcXM7lXwQ3ELuQ8V7h+9VqBjng1Qh
tQsVJOY1iwlWnhYFyTHy7/ya2Yr75pO/zi8BSWnLK022xF3XEkBIwmgfPnkkdAwi
68CklNoqAl/q57YLpAQmcva7EfC6OOyrpeAT+GMhZZRpVp9CMDNzUZlYLmqDOlMM
peIKR7KGWUWBuuO3j0SHr3J1YPYu4P9Lq402n9ouCQlISuRW5qNZ+CftKQmK5pQS
ccInVatzBtXJPS2QSqiPofTSwqn3rzXwBgXkSwTaTonQ+x4/0EWs5tTWUmz8vpij
N1UessY3lIlNzcXkpb2hLFhIsHIuMdzvKI0wkWeVfiBb7f5qitHAAo4kweCznluV
DA1VXPSFFt2yNgrGkCVFdemvTNo3A4fEOPw8Ti6R2uC6rlgHxdu4pTkRlDU5aneZ
v/tjvB07LWzZ6zJxQ0aKaRaNxfWyL1Jn0OE9VtzX+Z82goFwj2R77CmbzZRjOaAs
pFfORN38BFtw7Ovh7KDQ64vZXEhlc5Q3LM10Z7onH2siN8CDrzHvSRG41W55BhnN
gxcPGnZRpIsQLPq86v+nHde3vDLpUbQX7Yuds3y9Ml8Z7rDRSz8z3iQVMh9CaO8l
fdee9/XwGaHeu2UoSmiqc6+FfzqdmUwRSAWKeMIKJ7OwZCHzr3Y5bXMheunQ06l/
zEPHtVLfhpfxAaWJi27H03DYAjsYddixApdzcYm5YWx8s1BsMM67QDTB1cmK1DDv
1a2+Nr610VPIYJCzbJ6Fzp5n2+QWLXT0i18C5dTQTW/oTAlmRX0epXUnGNENZAw2
5kOe3XZGJWTTa9B1og/H9I/CY/SSsuJstwG1zKpTZuNE70dfBJMNruiVmLYgT6QT
4KnSrtEilc2eeVsvAjjF/tLFUeyR31Bh6njHeY/xcFJS1khS+yi7WBTXAkw4ytRv
Ai+DMJUa9tXa0bkoam+vmGXQcK8dcCex0D3dvRunyzt6I+7heL3DfxTjmbfuPpcX
9kcm53VTUVCQZgcEZVBNDPl28Z+0SI2c+r8YaegdJpeaTyOUjBhnrx0OWHrxxxIh
3Dk4RgiqeYxLqcPVnSuk1MZdB39J7U6AFJ5cBRyX8sRKRDAjXBeB3e2OgsjXQH/7
RmgZmWfLLXFyYKvUGYdWOLPblj/KKpRMwpHrJH5j3nBpmgFHBgHAieq5MAAAINX4
qQX1v3UNNq+kO5XYrQBj/31K3nEh4WzjUqpL+wjRS0gBh9V3qc1cXNbH9QK0AAtC
qDtKbnrvqamAXZ7GeJr9+RinWBcqLQR/++4ubA6+j+cVpRdCS9PBVnI626ACE6HZ
YsMWYTTuTGgS8GNITaknWFFU4+LuX7wnr2fo8oC1biuxlB0nJAuWnE9gcv+Gbl7m
3QnIVKh6yTDhJrZtpTz+qH1L1hTbzbW3SpS2+Y9P89TY8YVU45j7VnwzV/Cm6AH/
kZxWZ47PSzcyYpxo7zg+PoGkFV8ZMfS3JNpNlZDvCZYuQO6W7xl2zwuy8finHGDk
ROtucxQt7ltmhhfW1hUr0Yw1ue6J03Ed0GfP8sNxeRLMYcG4a5ubTehiSu+Ny0W7
19s58sAohn031FAZ2FbCiFWEtx2VlvE60NwkfdM2/W1NgsdPpsfHzNLvg5mODSBg
13zNeBETUpXmrVLGGXjlam5vacgnRynDJiH6BKtIvCRDhyn8RphwYCHPq47JteX+
HgnGPAk4plmBCZMGh51jKRGufc0DuBO5msGX8LNLQOP0Xps+DsNsp6Ck4TzsGa0k
AkO3OjUnzYUGs2X7W3+uqSvPlZikQYT3izFodlC/M9ZS+n27iy3noNrorU4u6343
gb0QckXy9hPozWGW671MiXMhjEb8CGjxYkEgzqyWovEcj+rg3OBPdNWTbFuRjBT4
fXA5hLNTu5dJKcXRsolrVmn3PgllVJ8hDudvNfh98+I5v8sXDem+n3ErzBeZgcQv
ZjZG/j59mIoR54AdXlY6BTShCZ8rdW4Zib2Pab509PrGxJomWfOOp3jPACPKdZc2
XwWpl/0YcsuJi5U11w1vYAUF8PsV32WJm/TxcAfMWs0jqOTcUMPzFWR9d4rBYxEB
u/Qn9ON9Iee5H3ouR7+hjr40cUu1av0N92Xjh1YOb+gaPE8vf1Ccm0OdmEDNh2vg
/oGHzRhpZxPf6BiFIZvspikeB2LtiW8uXp8vfSo8TowwrkmzWxMElTHhxrtWv6K0
O5x0nvhoDSJcqANuZpdX9l9g/S2LAWzdfSF9bauOK4JUPmgQF2JjjIopiwX5Rxl8
T68/FNlx6Sb8wHUoCjjK23bnAY9piQSAg9z4bwE9U0IyM0EOrJv2tyTuqpTJTQ8K
WlQh06+SQwBFNqaOeHq2AvWv7OEudjJTKV7/99FgODKvT3me/VPJcVU30TSk+sVe
rOUIhw3o0yy65fiywnph6UsgYpTfKuIM86E0ewSqWPimZtlWo5bi7OFezEyXFXb8
xE0AXeBocuGYmKU7PhXw64abnddYQTBbUuxQOrcGtJT0y2pWVPaBwRvBLYhWjoKG
5vSwz+pPhgUkKBrJ7XZtq/ILKfW+TMp6BWE0j+4AsjtnRvLN9S9q+cWjzKKRMkbD
zDpMWa8cOSIQKeauAbfLdSG7AqdOr6ye9xtpZmc6B9mpMBUPPT2bLwnEdOWA/EX2
VrK6YHFKmOVto4FdhHslA/sYsMSpmOqOxyK8I2mfxn8PmF3fe8xb5nFVHgtwVV+o
aEdS3XPHLGWoUvQrIit0Vqtr6wvNGB8WekKUnEMpjrdCxhpigaa+MmQIxB2suMlx
3IO/BGRBTk+3EaEg5sEOQ9a4+JZXyh0YiUE6K5+Ur0++8P7C5tISwQ5AOW6rVwJH
vAIJLAZkHCbNn3IWs/U+lKfSnA2k/ojCysV/M6OHCh5SyGeFnd/xhgOwPeF8HHBJ
r+yW1Ew1lcl0182YuhVITZOjedASeu0VEYM8na8Z6EzGGO3eScLfRfPdU7bqq5DU
IPpH/OhKgHrMyhBOc/PBE8hyxM6RRKkPEYudWD1ltRJgvz9FhBgXpTr717kLLTKl
IlWa7nLiVgE+8DMPWicXlz0jEJdP0K47Oe4zwAzv6RkPvICN7d5DMBnWUuzhO/Wh
mEhz6pArmr/md8H+hJu8Z3ZXnn2uzp2I4LgFsnmcvnUxzgP4l4wpTbALuQviHjjn
8BfZckkLyV5CqXB18mcJ6T3Kdc/aa3YWpmSv1ngV9LeQntmbX3JUGZ8vj0NeBSBT
FE93/yY1lbkKeP01uyIhNVuMpzXGflxpHrcjYGZurX4RDQ4R58hK9e+X5T3qB2/p
KqS4QwazMpCZyLTAwJ8cJdZDTjSIOBblmmb/6xw3xuYCpm/GRGMNkO+gVVVHlpOn
R+CMdQuWkGOx477ZDIqhs6Emvcm6d+qbRUfmqnN+ueCqa1O4CebFV/j4zSCkuOIP
peAHZD6IHJpyhBy4VVmzV5FvFY4lTIQ1v+HLrZpLABL2F7kh5gAzs5WGQl75w/Gm
jk6qSLowCQ/+Pb4bfXbzAcQ4MwNBLzk3Jnn1+CSd30VTvkcilVdmZqcA2vmyP1RM
hIb3Wh/nFQSJIma4t5LN2qU5RcRAlsQupp53vYUDTnCosttk4c5l+TqxiMxUbV1e
ToY79DgG6hRTJxjM5+98vavk30s0IlXvpk/oTDr10ibIyknBCK8FqOHNBVgpt1Sv
mWORJtifLjRFx0CKs0tSf1BMg2jLbi1xGSpAARnM6PAbEgCluP37LUQ60oMOoSlA
dHkDNpKPH7aBhVCIW2LxRbbTVrKRnug/4J5I/dNENIE/h5vejefz4B7Y2ZpJNWTF
VDOTGxVcMXkflI3MAFzhKZ4oDBzYYGpm71lCQD9QNHUc2cc+T+EtiFJy36d6pfNi
hZMMnQiaUclcNlOOxe0yYzn+sbTxh9Zx1bVEZ6zsamD5p7+06Y0zTojP/u2rnKjc
/UtSFYJgGyH7D3lGVyV4kMyyG3JMUFcznyTmCHLYY2MrfOQueULkyahYOFzIUCqz
C17wDe9eolFy9te6sW3cBarZVeE6AwTLl328MGoCZIdFQPEG2f7ROevrw7g0vRX+
KB1ckqbWuyJMiE39YdYPUkhyfbnBifykn6ZAqvQXSyrl7WNa15XoBxjc7hot4XJb
CdpJNapao9XCo6+2FMGH0AdiKqlqbWMyNUx25I8lXM6lDHweXnPL5WtSxNK6LhvN
uB/tIF1f8AFKRhRjf+g1WFiHEB+9ELcDP+zEKVLYuQ9t4w88fxeil2YKweIVT1lt
smuprvhJaW9H6sL1xygM2mb+2HnLy8+yhQxeB9+gbrZrHiviA5mcHQ5UV3nMuDJ1
3czy2dWsrvlWdT5w3wHRaC1WNO7X7B5dzd0QxyWzUidK6lu2kmyeg0hWE5SFnkzy
fPJZzDPxBsQJyjh58t5tjPIv1e9gkUWkL5E8xtA2QENBXmdzZnsBD9oViW43I6Xv
qYs8khvR6UALBju4pSQfubmhwgVstvev0Zx0+1MuVm4dDFkK8r6pWoEz6MgTzBtV
XPsRr/PGf4qzvw/lFKOga1mG6nHWbqOJDP7u0WNaWxT9sG6gsDpQKpQzpPI/o1Vo
1XBMbLYAE/psPnVEkiNN1r1ed2H9ciZPMsm9n34sYVXTRqNbKy8pqBdfQ/cg+nUC
PUHNAzx5vO7lZ2ZPjWCt6+wi4LkjmXScUHQBJ8xVsuLjI/Dq+bOIbLaIdBZVp4CN
qgCoQa2NEcRb+wSXtg42wQoROH+CLMtTzEzAwgBOQFdO3ZJuemXgESXJtmHKEbPf
XkYICS9LFV2JwYgJjtqbgbb94xDXRSlcKKnylt+RBqd2q01/LaJpx5xt2jzg7Tk5
nROKksLYgy6hYRoyh/7wzEHXOoadoam4PH8TVtFJsaW6vFJhAQ0vBJeAWOOGJnrl
GpDch9DOVx2CJy6nRO7M2I3laGVfnYa9IBLf5yGF8y0HK8m3NrrdklmKeIDDDBk7
vjKe212kcsCshBsgYVyXTUu4McBKVRbur71iyNlpe1/K/KK+orPA0b1e6rUcKQnd
AGmPrxrnaWmYWpxaQB1Tz9xtGZ7tnIg9Qi5K+IRRrcCnnBZKT+OekZHXUu8JyMSN
Hgc9ZoqtFBUoRSOXa53sWzBor09iLs8ko/Qtox86su98G6haq78jSzyr0bKjxKuX
YgLkPoxZVIVuMU5u+kprqkCZRADTUnjDAIa4EJBOzH6yblbNE8lpwmCdpKP/D6OW
D5FWFo30a/6HCG/7hThj5e38oz63rJJJgXmvP28/HmR0vTUOT5ii14umQ/nlobrh
ulyUo61LHGtPa5gFIJPXBxTbtyVYeK4C+/dpjdtBCYho9qOmUHhim0ZpXQAcWI1i
hQHdtJ4KUqjJTtTwxLwQ3q+2htO6dOxci5cw09CwpkzdVkUmFJ1CuoXmudsvTYCG
pxv6clrgBsfsXgAwet8HCEC1C//xyCI2DwzNAwVPvq9eQ36gImDtXvNu+IACDrBk
fsVjHhouy+jVkuW6LApLqgIiTNrDvDROaUVT5RHftDlcoxop0/fBVgm2K18tBMWD
ThO4xOQ7CZHxij9ySYe+M2hq2ZaMfgFwHdNPV7TLoaWVlvNmiuv1o0c24tCTeP01
guKIUoWWH9Q5Lqywp1iImYvayjzYoDby/hRWErPXoIENCH0hlkzifD5efFa++bRK
ZhVI3MMAHXr2prSC9vSsYXj7YUOMJF3ScQKdTsoD1IWeWs8otZ+i/mAUZlrAv6NM
U2NmChUDq8REylfo+iGhm1U2eDaLhAuVzj3MEY06DP906jcMzAodM5tMo6f8aZVh
PjosOOs7sF6daGcnB0f2zLPCyFBbDSfdFb9up76rpry3AjTDN0FZbT/v4N5DV0uZ
qm9RlSbfHySyNxNeGeL1+3TfcdeQSGWGKfoXIyYbtRGeQ7VM6BV9Rv7HxilNs8iH
lRp1Xjii/sye9dM+xYqaYrdjA4voOfEsmD2LFrFd79yFIxTiigIBRsbUJ5yXIStF
UfpYdtGMRRPrLnjRunEGW1HfTm+eI4xpa5q3pl7ClgbgyKTQDPwjVdgyyEc5tAzo
Yz6/nDu8Be0YL+WIO86lK128EE3PPkMBrzCqUD2FeBB4H59V+JWwlUdMGMmgktdk
E57dg7+6kJHn298AfXGpdNDoL9MN1Q7wqo2gBUV5T+iktB0hI6CLdy5tCrsG+/6W
MenWxRlK6PTif3rXtTSX/vU2dAm9SFEFU8fiYsj1cKv7BRN7fOPoSDwvU9PgE2Y0
dnwimQUHGuGbRl6WpF9so+rtMHa7z2w7UZtWJcCG3hEYhkxPnquS6hlzROe/dD30
TMYw+dxGhLAeHQbH+8pqMUl87rFkCWmdC8O9DnId+h7zMtDikWljF2y7xreb5Edf
zzFiWe5jxd1FnJ3rJR4/g3ysGWq71C8zZRTuZWSxQ3NFRZ7T3Uq5AJkkwGJUX6qv
fBw+vaPPD38AR950Wz01bcZskt9vm11Op/iEFT8ALKMpHsA4RAZNOlcbDewDc8fm
nyhG2UwPCIOB1svigObZUgAZuhdejp+4pfWST+H6mmDpOv2TDUgAoElpvP7cjAgJ
RajuW5rTp1rugOkCiB1xJOz5+TrkKnog1sAzDB6izTdxsFBMlQVvUqaNWI9kw/lv
QSQilvfnC971uQJ3pTYWqP9LC9DV7bypF4jfIj8TXaDba48LWM7DQyWY+q0VGy5B
3OA6Vn1bTaKCledVyOKIRzqi9impsnV4aPVXdetB9zHmx59hRPRav6wBiu9H1QFj
yQUEc7c7RAA++QPD/jqRTl+dtUL2R4Uf3vPPq2j41aXW+I+7Qrn4yRW1+P0jdMuh
J+5lYS2AuBa4bxoJH/oBMd+okSkB8cucKwlgpfHolmig5VMmRr9gYUDe/kuGVUV+
SdrfkK0xucWcdA6IO0VN1GrD/REvZ/We2wK2ookPhm07RKkXtJC5iwhoEmj7v2rX
j1gnMHzMsvvtp4+xMS1vyN9EXBFpDyTE+rspV6f+l8lBMWFUBr5ixxenTrDYFx1K
qGBVd/BXJ1hEqNBO+p6Y/QjyrTjMJJWSDZwVSLxhifjqn3mto0k+OULUCxVrTJkP
71ZLcWWWXbKb+h2764LRLSc6HpkttE/J/RlG2gOU8BDSXKqPplIQpJxCHqOpfEz5
GW+nSn7q+ZYtq+FrQNV20K3RDMDJuKHjRj6yKHBZIPOuM6VDCffrBRBouloFMv5q
oz73lb64odXE0ElgVPK86ARe79WzyUQlIarPqrgAXIJU2bXAZ8r9369uYm02pYTD
FBPtWhPPtMkpuJo1lu/wicjUa0qcsM3z56EDW/LfTVFyjorJNuKaBbM67Eb1LEBN
NBgT3a4uMY2llzzdeIRDXfc+VUQdodMc9O8hQWxT89KRvaW9N2iD5AAlB1V0kLHs
y4x/pUgTo2gg8EB4a5PkKvY0rA5J/QagXbuy9jShNiYsf2nsk2fb5Eg/+2I8lhlA
9H2x1IdBrnvjKEIuaRin6XuTUXWxnUMQTyS/RqBDogOZf/+u4mhuToz9U866VNbl
nB1t0rSFIpNnGwasxvFAcJTRoQg2dq4NuS9Mfdq6cqJnNqh55utcrZu3Gis4SDXW
/1dqMSFXQiETmgUCpUkOLHmdV1MFfntEqo9xqu2yngUiYke4+4KLrGCTQ/8ZOv16
Pe5iMwVU1hHjAIpFcNbGsdceSxm6oriYIwS1qKawYn3hB9ZDM8ir9/VCHUf+/o47
l1tQzl9wNNadw3XrUWkTbf1PEa/9wNU93fowWNSN5jKcL03tTHv/ojD43maG3rR9
1xoIzmzVtrNyr7jcZ0jx3l+q7d70LppXuVRwlcAsfDfFs0lPY/MvpdoohfICHw9u
PlXNKjGO8cBOxoYT3KxBiJPZdYD04pcGDZwmHstgZMOz9PFXOfhNBhyiiWeq5q0i
1bCuMdXlNuwb6yGbIptq7PhbbqY9geeBOsOr91PgoRV3gvQiLJgPYCwPkKgT/TvX
Vx/YQHXHvN5fm6xD4IWaYi9IbjYjYFY3u3rJf4eddfacvvL3IfmQ0MF46Lddt6F+
xSgvZ+qn5Oo7nfi1AxU4RuNyJBEWHx3SsMik+EHlNshZV+RxGWcSWAsFWBPn/CYD
IGOk7sD5GLQcVlCT7JKSmndbMouiG4Pbtl/11liVi4daEFlfRDPVE6KTcDuDWf8K
bQyJNeJYnfwYn+ZNjbYsZEH3jMOXFGrq7Zz46f8oDLmghhc078BTe14bBtIt2CAl
coGxW78dZgGfNEbuvLQrEvFIBeDjFhsNCSlz2g1GZr5jRpkJvqznflQ3atMAnKt0
TTp5OnuFshEEl5szT2tQJZksPBXGak07KqooTRIbfil1dVHBdlMfopfKIkmfRbTQ
vWysLJDN7+ZJ5cagzN5zU/Q/m/0Lg43rbO/hwjVYwjmM/vTeHAPzjXd+R+uembun
/JY31tOHddflD/0FfLItJnIvLzHuIP8xduTn4nM1HeqXMdD2gP2xYfsW3xQNq9xu
Cink8k+MgPpDjkUkMnGelC0IFAl8tmM+qLBlKQPS9djc5aUIj32k8+RlKmU4387k
VaOpbDRjP39Qbszja1XH3HhTVOTt3AVXa9TJElLKVOWEGjVJERQMubfsngNAoeZ3
168ipMdjNTea78AyFJ7ji91eOGZ7TOhJxhMrieUnoYMwidlsFiaS3MUUeWxvaRAj
T1m3YzVDMqggnwmqYorVESa98RRNWW5+uehtVohGkuCtrUt4tic6cFtnX8QbhEwS
9FpVHGM3IKptaoQiIT/BYW0j6rBbez/GF5XkaeGp/OC8VnpwLaDCWWqrM6CzTDUy
xQ4+dUKvJVqAKxrAgr2ceYlxU288I62F976GfDLRH9dVZMX/6oRyXyYEs/Adbj5m
qPYRVbcN1HUFe5caJoTUZ8CVADKsMJRtCqQTL4u/72DC6T9X4wq2f1jgIrIkapTL
gvB8tgcq67P8IP69lAZ+++QDxPDojwv+cgAonCHsXZq2oQTaFOgNmGDo2KEDMZnN
XoHWTjTP7zDaUpYVCRzaUztsnVWCYitn/YSkml+h0lxwCUNT1ha+3gmMXbVcEWMs
2iCEzWd+tu3OSkTi49NQx3CvioKNG8ovQvG3IH2BVFe6rZnJ7dR211/v3lb/8kXK
yCDmGW7kHHQgk8INygl8LBuHCnBD3vfQ3MktbDj60VUt4likaYJY9iZbBRIG7Jx3
a5D4oirF2KHjB2tJawgwn/9/MTkoOhdsZa0bPpL6gDZ3ldcMEkra7sKmvgGoYUd/
bjGoUe9EIJCWH7qkd6k3r5QhMi45y+20IOPPTt2YYYFPtaYBeD2xXYyy9D351yK6
p5lD/Dyi04ugDxOm9i6UD4H6VlWdRD0GENCq5ncSOcJvaxiVWM7EuxIhMf9DY4Vc
YA3MrkpL2giYQddMhpld2LFGiYkNvg7wj/OWhyB4VOqyxG6Q6e8EyXVNtpsBg2l7
hbpFx5w3oAy4uh4U5bU8eZxSLweFKdOit80+V7r0ve4dNoYCZ4A3qfVxqcqtD7Ty
nKxFj0KHLGDY6dLe0BS36njZzTSP6S2eZIFQnskx8tlnmovoDDtfCm9xKywyl95c
atqDfQ5uEcSefX+mVzOOVfRwjpo2/sW6uv6EjvRloOs1IpbZcPTZOXhOOD151Jwt
ayAlVn7N70ntNqJqJPtkjfHKVupJdlOxaRghTDZZn7TJthFzHJG9StSD97uyIvDa
+XoaFtsut+dw1cDGRcjmp+6ntSHA5YsyASKTg0M5yzoAl913R3Xr4N5+q7vZjqlF
z1sJY1ZOS2m1CKqTTLECLqGm2vb8GYQ4In4Jk2EAaOoGCew+aSR+b8Gq3+J0Jd0p
aJ1GXpVzSOuRFSXF8+TNZLLKXdqdGvz3gTs4CKfQgzvHbNktUL8Tr1mI/CuhSYEs
06UFjGsTxg4edAQ8dqLBE2RVQP6OT01AV/8canrOzLNuIfMAW+YqIyUxhNQg6O96
Uh2F9nBMZeBC7CCWjaKt8/cqMfZ8Zp3+7e5+OSSs23tqIVhEt3wGbqHzvViJym46
hebKC+Yw0wU5TeYzpiGuEKHiGHAFA8SmD0py342/gvOkCFeO8+VTXTGX8Z9TTZZr
rzp66CJJKjAZFpwvKNh1dI4gY6zlhu41PSl2tWtVL7ZaeskUs38VzvYpLLrs0Q12
Nx+2/cXSC+iI/jNOkFwMvl0MUhfMh9UD/YzLZ8bzMLSALtwycrLV/MnphDqzxNxW
p96xnB0DCSLlDP9C/K/LESXL2y4fXZGQbHd3CSEnpb55o4ZeZ45N10VV6LmllsmJ
z7swMYK9cbJuCD0zEqlHMykmsoX94Z5YaNuovz2Q7mlO2dqOtlY6cIqXDhXfncNR
db4ilrnwNW0gy4mvRw0YtYkrnKw8/SqQ6Zd6BNNImsulbZzgmjWTU0dW6OTiZinn
ZapLmBwXvIQdLu7IO2S+wSBRcl7RcnTZXjJ6Ai5KJQMtXqPtHDwfS6GwDSbGz6LW
N5MUt6jc0iK3xqjlHH/AcCKdelN8r4627Kc3kePvySIGfplmeP18HWutGP3ZjM69
q3UE+DlLnmgTKYnOTn+81JhAlfH72WQLjZIH25cAxSjxmOj+TeOPAO/cfIHquqKb
MSJcEOqVwpSvNzUh+9hOO+vRMkiRog/Dd6GWCgYYQ3bhZwBkLakUJPE1XC/fYP4m
RTEU0iYlEVe7I6rQ/ys/sSo03zpiBdeXOlWnqp22eAHTejq08FPbApAY/53KBkpb
K2jPb03kv+CEuzzKveRrZMQajzb0PFyyhL9CmRf6Y6AKEXPPL7UKrC+1rdzjAaK2
EQk7H2aG+SK2R5MiBtTyiU6YJIL9bbivsdpTZhEbF2ah7Jh/vuKJ7Ol33XJfkqKX
nmqTskR00M2snO9562FWbfbCInLTSB/swbXQdyEepHe/XUxG5OoWBxk4kAm4raRA
EvZ8sIEkS2Qvi58BFHxUbjZlu2GfHBtrr3oJpheT8PF29KWr/WqyvGp/OJx37dqm
Ed8HY+b8lka7dlezX1FQfo7qOUe6mjZ4HV4/LMWMLXfs+ggvMuoZqufp0cX45AeG
wZgQ6pF+nwUNDqdGcctTMEACqCu692vtYWg3VUtDkAcuo0pqecziVPA9WvD2p7LR
Rsb+3WcdzKYbaGNdiFicZz9L2ex42xM6BJPQrMmToS41wG8Td9Ux786btJ/tj+F3
j1en6WjU5ht2Jrmkn0F9agR5ct/3dbumTZaZ3p5MnCt4q3hlghk614ScujqpmyWI
p6XjGiCy3Ogt5GJbHEBQCU8Km9bxe8Yns4PFlO2dvvnw6MQK3kNl/CHna0ABlBdv
z+AtuhAcuf0R1kqNzrQOVOUfnl5AWbZ4SF/7ScpoVa1FJ2RIClAcgSEBhDGXiRJa
HEAjg5eGfrRPzY1DhbFoRMF9KhaJW1/mfQywv/heD35cHos8T9q/IYDr94qIAFmi
01fDzA40jYj2gLk0Io3zcNX3IAymYEPZ0xb5AG7yx2QzNLV6dnCBSI1QvcK0raKx
npqW5bEp2LZ8gOWw521ZyKsfZcyFeb1c6OpMHrTs0+7JqJG46T7oW72I3acozP2X
ianRUAw/MlfPxr2lNPMM73L4F+XmdD1lFIfAgh6oLATP2d6/PTK8gbRp1N3RappY
k0xQrGCwFqvtZ40xBNqw/hEssfmLzd9dOTzecr3xjjNhUwCyIuXsM5bIgAWM4N+k
sk4EVV63IR/JSf1VLQdM/OlLvpH+Y6mc10ZCAcu/n05x35ZUkzyyLrdFTbvBmL1Y
Hcnni+nW6g2rCBd1i0JJWPyUYFASpbcBPLRvdLXkMCjAykdgKzJwiu5pJu2v8vrw
7zaLDHgGPoS2PzIERw7rGoEzlz9WAC9gbYseWD3WgPvs0lorH2l5cJbM9SMDf1KM
ldXamEbVp/VpjckZIa/6oaFq/vfo+lzb8W5aeyNVmeGmHxxqjcCeSFVbuaA23KLz
eKRW3kfIAGDmD0aRbblkGgYJz2FEpvE2JAwmTX7g5sDLSnDzhaDlNSojwGiFBodD
RxmElz85enWGdjlMxBk8onVqA+bsOiiXArTHaAaI1hXjD+5XmRBF0nZhgl6CM08K
iC9foxtuOxMWrH2lZwNGQCOxHsrFpr8vF54c9ucNm+yqMGJW5/1Nnox4ACRFNDjm
y5+vU11aPH6QNcOa3Z6JpMIb0GB+aCynXb4DNlUFr3EOL04DZALmoLFLHpaD1zjQ
wNgJXNoitjFbA5r5iIHt4ZIzzFonRQ6T+QFBjaHU9UnLFg2iajLmbOsctnXEOUEK
p4Spdfbw+iVXA1oR5bQFGSeXyG1PJ39L3YEYtlh6/O8qnttvk+PyWybinTZRwcwG
w356FCvkWtyDeAnDOw4miIw4aYmVw8oxcjSMNiXqUcChOz+8L1m2bYSKy/24n6GA
YVFngGyS+WnSGHD5ayL5E0Nm0R39CvRMBpaY1QIMntzKM6roq+nY/J0U9g+nBsG9
SGw6G8c+ieZHid0WKATLbDCP++t9ChnTe+fhXZp5TaWOqm4yRSk3xWa04FSi42dt
8xmlzKWPC0zUOBcmLtefplrWgyv1F3EJzsPXAY4nZF8HL2zbh1DRBKDqL36F8cFH
QhGufwny+3VSh3Wirs6JzaHAqlxOiY78InJfkttuwI9oRpz12scfD7XB5ITj+glW
F9XATq5sDHgzyS3Qu758ErFW77NfuqJ0mLASpjNVViD4WZsBvF/FlWO1id/14h36
KqcL+5SxZoXnxaOeACKSgG6ZyEKJhVAYrZ0kmTNLMpyY/mjsKn4XQ5cW1nKnKqaC
ZcuD8VGGlRDaQdQ1P3kEsmcrorLZnOKpjZA/l5jPeHPSXKLwxKpgKqiFgRAE7tA+
8Oh/Z/CtwXNzAHwylQ+Kk83MrWdF5onwojBS9oGEf0AF9xi9M8YMpafKF+dXG50i
Hx0XoQQLX7KCklcfK9dEkAXXTSRyDf2/gLBPV2jBd3VvSg2fgY/a/ThdbXkt41xE
194ujDLQNdlhO2J8R5AL/hEqMY5RhpqWNf1dc5F5QkMuNFnqzPCAs2h7IUE1Pt+4
/49ZeG756h57Ky7e4rPx38j2yVZmSF+CQepw69dmNI4yt/jimVgQUGSNXQO+QLJP
6WI4aRCjMGQiGKxZ21tvO6SpoXi7ppErbcgHNGjL69JQO7KUd8elpGinpYQ/XzAF
AxJHrGHHrhdBF1tT9OkhsNbm5jqnYhgEw9LrrbWxQnVLwT68/cOIZZ2mJqVyPHhX
KqU9wuV5Y01Q+FH0x2WqHycUzTDJ8FWeyUwCWJq9Tx4WRg/xxTt6eU1xKBfsVGT2
ywo7bRhLPSmVfFxDFW+cOGWNZXk0aWhc9RXk/Bmay+F1lrCp8Z8wdUV9M81JA3Qz
EVJOyoT+jrFnvt27kbY1IwBzt9WSck/aav5zLXekobEPwRY6vMjZM6Y44ZmPuE/J
jvdqTC3ZC+s9/0ZvMFM/FUfamBngtV3WoH/HPIURDSR8pN0yWix8c9bu4f9DPzsH
Boc9zaBLQZ5rZFseGeWJUwesDd6Xxk19oKSyAX5J591w6VaCDw6rE7wngBUpeq2S
en64ksZehaq5qlc2dBSsOocenuiO7JTFxNBnP21jmevqOvqEXTPJ2ntpPRGk5xEg
g7O2pA4qEozGAEnILWNWRvMq9hBhfMj5aZTkGWm3Ya0Ub03ycqIqaYH9Ogg3PXwP
RKBVlM/UBrbjFh3APSHUpP85scKw+ddErOKQ/qA/11jZfqCz2RpwYALBsYY2ApFl
3hOC5l28jlBULEFa3k19MlaurboK2qtYdRYkDxwUgYxG3NbOlkC1nNIxBxWXYcUF
4GMEzkj0/wGZ8+60R5dDZRLi3SggmEQPxA5mNc2FHkdegcUNlrjc3DGGWtfejFf4
rjeITiQxbHvzQHxUscFjbsV5ss34KG6IbpcbAbSBuiEB/6bKhUlds4tD7jfZweNO
jx93RV4ehvtSpCI83hrXip1QordI4icw5vZUVEczGa4MDBMZdFHlUM4C1msxNc5T
7Mzf/zKIzdMICNgvoWMhWqCDr59fRUfhtnYdwa+pT+s+dnzqSRUEJrIxv/kSUqM+
K1HVLxa01h9ebzsrjvdu2DfgYXGNJ1uHc+PUq4CBy201+woQqfI4ZAQz/mG1H4ef
AP7+08+ZHvQpUZjBbnHFHtEnP+V2zTYfrFyMEYRtDsDZNBVqK+IEHg1h89Nb07gA
xWy9gYuRrBhb/BzZZevZUgvnq/NM7FV9BesQks6NWqu2UNk2G7WctTf4CmWCP4W4
CDssLYB8Zha4Wkr9RMjp+nc478ecCgQAjK7b85rnDujbp2ktyj5o5tEm2SJLFkt2
E6eOgxnErjG6c0iRMwmXEqk6vRTGXIvBDSLbx2r+NvQ0C6jDDy/pExVKOQcnG+bh
476OQOrc25CQht8KYC7Ihu7r/d/ilBdrK/YIyUnCpI2obqXOJBZYzk5sAv8Nz4AR
IfzU8k8pDbWJQXco8HkGWPYyhPQ72Q0++ia0X4EERAlb4455HF8DFnaOW+Q5O1Pp
W4nvuqY7WPA030Cq7nmJjNYsSNAOQW3B6chpvra9wqSOwyqXo+II55G83HG/vvn6
XlIAGBQT3Bf2UifvFgOxkBMLB0C6Pr3I122lXr/CCe00lgWXarVldfcVygyZx1gC
mc94kpRnIvc/flmB/cKZzv5cMveXIR0ZrjYDkGVLvCKIjfsvwGq+q/nxlKYsVIEw
9DLYBmhuIvwBu0hvA227RfOwbxL7VpVAPHHib9KVPZrpnEHIugcJD4FZRPp1ekE7
wNlEvwieTW3WOJA/pv1H5JLJWa0X/HaR3M2hnEmsB3ZwO06ewYoydyk7f7L02HT7
koQBBdkh02E4yghgPl7xB43P1OScrOBP7piUBHjtTcobUBFNkd5VV7QARLC+gGnM
BJ6ZVA5AcG3K0Nj06dyFSV+KKP9EwgPY/wlrLZkABYC62Vp7wgGGmDUuUSyfC0VW
xMMZzn5yZDMphNDP120Mslm2Mw2gF+ajjPrBgBucbNvIlr/4bAKms7dzOaDMgewH
Bgw8P1dFLsaJIsuXu9Zv0m2Fhn8okl2BefUbmS8l8bDe5YGih1La/QfEAxJFkpc1
ZJqP8LDJ+3m8nNCOfGssTBMhOxWuv6fpgujg/NoMAWi5R1i4xPxDX2Lg7b9FXu+b
Xe1eUSUtHnDVpZQip5afAQJnMZsJ6MzGBwdCkvxJyvSwErxo3z9qeL2W37Uuh+vm
Y6gs027Md0tAR1d7hsrWEsQ5Xe7Ofu5cLaiC2woJL7cx3H+U7Dhlfrq8HMuYyDJq
Hen+GyaFjIf4KXFet4GeElM8kv2QK7UDEKhKVCWgaHswjwC+6mf9bVwOgpuh39Ag
+y0o09cjO+V0SftApZhlJK8bYmU+2voLIXtWqFEXT3pohia6DxPVaWiZZ8zhn1Zg
ntjN4q/DIhlOX3A9ETVDt0uqk4GwXSIDw/8A9zBtDxXAix9Me8ON5IiCw4+brl5U
o60j6dU9qQ9kLmG66zjBBF5z6H6E2SxUS5aSXIRzRjaUn4+OxnqmfyR/HQjtYc0Z
dBIFaGvbpYD0/SqY8oGJ/Aqj5rsvevxeHGiP3okvYrWclrwyTqULpK6FvlNxIZBg
oMHiTraLwNDR1JeqU+5u2jOpW7uVzOxGHikuTtRS75IKNnRlBV4Pjj1BUIqlAsng
Iir1tr6TjwIq+dOHDHtNXopoWzT6CcFtu0nizbQTKSZvyRA18GVxnN1ZLU5sabjY
z7Y7zDN7RTEld4gydMcL0LVGqFgjEbRGjweAajiuIzCWIIXlPXyVG32SrGhLPoeo
k33tegGQU9oEfRMQ8mP2iVlunJ0epn1EzCJ8zyfn8g13lorLuIM0pW5XnB5D0HHg
5YLaw9jRBoNCY2xFHASsfT68Q2+VDVrHoE72/ou0nFyNFuzfDw2UntnOGmoadorS
i3jaW2HOgw8W2Xk9HfhzSqFh8UCB0jgaxwcqqSy5H0NYaPBytSqu63IMbAfqVknt
nTpzhz5di4nHFA8cuIKVlrCBOV3HTYVc/IZBlQoT81oa+aO8ZAhDjXee3JYZ/K2x
T8DRzv2E8YN4C4jb5nXQdrmkuoKsRPIV94sKFr9DY9dbI1uFXRAwJSq6IMGeyOrk
wyrORdXCyw8PBEJOCUL6+VZVi5FeUrj6vUK0GqwUYhHGGTjmp7Dtql2cC8BKnft3
3qwJlafrmZAOsQcIQ46IOGZGdtr4tm8kSMjT0JeUJc1DHNdNTYROI2kRlILbob6x
KEj/GLzvv4c591wQSDb3yF2D2w2Y4l8On1BhGlNSYG8VC7v0xdTK+YlZYYO0PLKP
YNRQgUBlUW7H7kiSvqX2QXXt39wrO/DtyQAj3gDAL7aCjXQsQRqhhfEe59LiN8S7
fypHpqyukbXox62xi06J/ZCCAriwzqSWlx9FbZmmraekCA4l+4iAF2RZWvyMOItC
fcA8/Vq6/BlBZ+ptRDz1lJdMsQqhOoAe27OWSVaxWqPfyi/Ic92jVp3scEpllMjw
CgVABw2rgDkBlJbHg39a9pmxAeiNTxQcni++FCahCj4inDTGNmwqU76mJcXOn1Yi
Itk9RzmXicmcQ6o9ZpIRjyfWkQLfV8m+pMBGDWa+ELOJPlijCVgJc7rVjmoHPEG2
0ymJIRF2qvJnzzqNkEtocPNwK45UIYfzQtT0vTBi1BehgZqKUAdJG1NpuWEI6/O8
Lauqf18trkEaskpyLsDarlxIT41B2vVGjsgR6+8tPL3xe6L9uT79OYUuwxro92X/
3P1Dbe1C0V6VpPF5T0tP7HSQkct311oujLQWqnmDengKXqTsL7serrmE9qgbrRZ6
dJXrpBgimePWlZHNw5v1gi/lhhNboCuhfHuID6VtYnXrLjKgJJSdR9/w7PTKUpxE
BiuPlne/sfa0ch21nFxSdUTTOcQjmk+ADsC7md7iWs1VF9J6xbzd8/a+Htz4ZtUr
aZ0rxm3F9DL29fVrw2rgOKU6NFto4jZv2EPnrW/B2PvyAuiGJ/SAX+e0uYz5TWyS
zOTKRC2kxjihzZ6zTRQuOt9O7CiZKMSLxfNe+s3v5EwV/XkWDCG/6kNP9sAJMYcx
OS/XC5RnePCa1LNXP29KZSZDD8/Nriqx1WNqV1ZNJ8XmgaXF6apun5W+b3fY97TA
OX9jkkhhLKq0/yzNI3zsEy4OFKDGDqT2LjJjWitT92gMhggaaNJrnui7FrNZc6dk
K79NBduKLE0DNfFpQ3jBeLKMxuhMEykeRuM8HrJNq4naMf1PLhKGuXejd9YedWtc
Mmuy9wOsOUXPd0JM/SJF9v/oRH4RzHfnzlFqoER4cfooDV7+xz7LSlh+2g+q36oI
3GdA1vuyQXY6Xtc9aVHRfnxr9oedlkQ3MGb6jUfVBBMEp19Z7rXX2MxK/qHyrbxr
N92lC3ZZZ86AOnlE1vgJ3zQYvIP8O8kKTphYdWHQ5nk+O+v5vN/14LWA00r7lNEc
jUtqI/pQM3+Fgz4N/JIdPXsvspEbg0DDOsluNvKfDykxhPrri/eEvFXjFeRH5ioK
eSnpNuQMSaxB524GIrRR0tZOXB3Y8qft8UIpXMkyaDuaQmreL83CviJuEDuf7RZW
o53WQ4XY0rTBgcbC8Socvsp4pTcJtb7q8KuxHSuiNLxcvvxmc3n1xOTbCpBOSaXe
Xi+ZKivLQCey/PpeItA8bFVLfy8qHXIlLmOrbmAjbs6b9qdAnZxd5fwT3ZTULS0V
2H1ar6pan+Shzg8tbgM7o7vUSwB/pHlSYD9sBrNbjoZmeHdh8uEbxsKuXAW5M6eH
WWiT0hXb54qPnu5Oz2DlD0YakoU0BgCmiErutvX2MsayT4w9V8co8Cq9Es7cxAWW
isISM6vPjDDSnRuz5Vm+GLeM9FlLceE2qFpuacClFp9ukReM49kmZXB14dU+E3Dh
msGwGmXM1l4x36Id7BvSnjLdLWG9RUAkHcTm+hNniTbz2L3GR+5KlMxpnFGS0AEa
qPUbPcgs0Lmx6XdyU+P14gBMMV9WzZuEYVXxujKRN9kcA9vBHkxG3PlLQaDb6duk
c/W4zYg34OEqAuU1dO0wPF3j9TcLrweLs74MpnNcPc5D8DzdqFWl2wVtzUfEaYiw
1sOWQA8lHZkodxlt29WfcdkMsFvNl/kY0KVETXetK8PttoYSOfRrGKiy9ig8K1Lf
C/MfJNouHQa/zTP+REFN5NMzmExBAvzOs8woivsM6GKuOJ3IdnXrRqnluaeXqhhI
2muGMpBOCrj9C6AuTC2jcTzfzyp7dhfUNrINGtzEg35mFvTDJ8D66KF5gk0sc8YF
ZorFzJipvqTCbpW57f2Kb+6uEMH7E6InNQA1Hh5JnsLSMKtemJDozVlyWQCa8VwA
bYFXfBOQGBWghbmUYP3YVxUXyMxodJqTdY/xCcUA3ZKMLDUYh78cU836GGd6JuDX
5aYyNoDACKJfAAWv9BXGuE3DwoiArUmE6FatmiYW3NbpK4qqUt4XAyzz1DIgcFlJ
t/JP+lGFmHKI/712OfoDHBEgHTRXXu+ZcfCKAxIvErdbTl2oG0xbwuo2aKFiqxRM
t5MMYnmAn3mJU9LAJKzIb1u3Sc5mSRj5gvx17I+aC9XgrGgH7/xkySLSucVHBGK1
v8EDqPTvkc5LXxPw9A8JUi8RSFE7XEZWYMfrHVt0dUgMK1Jm+iK661DnlEWKWT4f
WHUpRrRJl86IhSTSks3Q4LEujVJnnLc81lInxyxAG6AWpmeR+vbe20yhtVLVG+uN
7ep1UNh6Xs/5edOzgmu6c71j3DzG8TVf7eOVraRAozyUw0YXW/irP/B/i+o8fLD7
/pGVU52rWI18QnH8N8k4+gtC6fJh5VH2eoTSdyBP5RYUoWRPiTbfD3nyKC9zZRQ8
8kn6Ogkkgi9oN3ikbunYE6Qf2lWdFaf3tgB8xwUzyGope54IMqCNuX8HVHktsPmf
m2ct17OfBHhV3b7MmwEZZqeCq+vkDmzzWvjqpHs8lsUxLgwvAdO3RXAzlS1CU9wk
AWU3sSfR6FO3tuto0O7one/iCRS9utw7ZM5s2b7FWTgkFnvjE5NvY6IRQe9Gl2r+
E6NvMTEsfRwOAaAsBZD17l7ye7efFq5JfxPi8sxZIGwlQUWRYA56IHR2NZeS8Rb2
mQwOKwtk5bDdbVBmw2o6w4cJjH4/UX9d1NX+vxhN3WVcZP4GOC7P6jmjgRjwkFMJ
kesk51CwfG0h6Xc+X/p0KIoQAQz69sLaI+JfUpnX3Mrhl63z3jl9g7d9IyA6baXA
B5CfAuyB0ahberZCshwB4fEwis432g12bURLfDQDVYN6XEHqq80Hls6LQUHFOcsh
3H+yd3hTk1d4jOi+2MJzAZhZCQup601pMRrokxRv+6no4dnxVRajhLpkrtFIoId1
ek8sMi2Jv9gxHNjX5JmvqB+/fCwn9OGzm8tSjrpqGtAPI79cTavumUQbEBxqTgpE
QSMuIzXTJuhffti3tGZH7OwjqohpQrziMvhTsw+xqejHXUzsxB88J/wqwmtH1kNX
tUYQsLqrfssksIXlbI0gVgrm89hW0ggbXjHk5sp6xksucKXco/3g9EAUM9NnUviT
v7kK/UqP+SgqYdz4So69yVhSI5bF4r+ADSYD/o5ybg2blBV3IE98EkGBatycP7O5
NAml1voWKEB+ZqielJHaB8Ldh5XYQc9JL9YoM8hAwr8mxDkvTycx2I9bfQBoYKrA
k33rcRnqqNM8zMTtYIvOY6tMjDSlfXoVKRAOtOZXuQcN8pwRgNOkOuTDKTjmaGsr
vD+p853Dfc4dEwcbGUs8bgVDZB6yLL4Bk/TTLLhwKDcXtOAf7lAQsAH+CjRU6Y4/
Lxq0fW5kwMSNPB2eYeoB1g5x8f6NriG4K6srzzc/ggV9bE/zBAH4eL7Exw34xL2H
qmtoH1IB11uVDei0TjS8QJ8p/eEysht+hysmlb9oUYBybZmXlvTl53ge9CRjDjUY
ZGpkuZf3tRLZnFa5ws3lGs0Oa/+fFYCYjlvbN9cbOY+lEfw3v2SRi3G0+m0eIrRy
zepUwHTKTEoqAoFohrm1VVzIkEzwFHBYE9Yj7RcE/mEUrwbEJt6R1zPLLR2fP0JI
nrk779J9Kyo/XNOs6RTObaZ/eQnvLc7MYzMAjAtfiIHJVqxE8kNjal4+FzfNusj8
Zw2l9TjE92DNbkno7qN0GMr+iAqPtG0OTYSbWzcYFi718Cca+48uOJ5i9hnnzB4+
xsD91RZdYDddEfpz4Y/QZyCZfpHbgS5+l8Qvza1gAol/DxTUhvx1gY+pEIoe/8yO
T5v3SPQQBs+lN79yh8R2SmFmPvMmb0bd1yKmLn2KwVFyrGvJPbgAoZCcohv+/1R/
n1QeUmWaOayZtfjS2SDJzj1HCh2/BgkhqJEpw0olJkRSNrijOJ+WYcQs/eq3R+l3
jAQPKsDSdJolV8k9l386EnKPpKCE0lCckNiLjrd/5vVVMO8MlI+etoyFyw0+aCxP
mvUbtKN3UR9USUYr5Q7LW2QG48xO5MYJdbAcvPhA0hFrLLy9HoRWUmObIFeitd/W
y/UNjEkmUpXLiabzqs4ToyhkJGExlpy+1CFowvTao94lo+0XwXZreH9hqQnP301T
AYJNHQ1koEm3IddY4UT0NsBwng4wgj+AcLvRPirTor12XcHF5nc+cODQIomnQ7zF
zjQUE+Y+UrnHF+POOsmYS7+ErhSiqG9lcdw3eoUYbiul72Ln/Z0yu/FGbGlOgNZk
YUnf/m5D4vQCsD0zT6P3tGYjCnSlx73fnAsOwowo3ag4hUNnoSbbDBlYeCnlIZB/
DQZmw23MQ+PATdEdu2pM4/dK7p3oJHEhL+QneVwncWIfxpc66zZY6aN2N/LvRR1O
liexIc6bNP9xdjz+t61KrFkhyeC+hdaP2H9eddj4PUQo95pIPS2WWAdOW49nTJk1
pHdWAsASQJiiIrfWWZrlUJ17AjUszPS+xfFFmL8/ZaJ5YQwBnz5rm05+1Q5gDkK6
CNIhzBSYYCdWrmmvf39lvpjwZgXuig7lCSq69nERvyBTVSvOPTAvPke9gzTlaJgz
4RLkNQ2eZUn3zppIvtBNoFoNnNyAUJdwWIFh5IrUekHTJJaahkHH3+1bkAPo8bsS
5KfsR40wz4rQ1wx/Qa2PNiFlBax6ooLIDhPp5Yukt4TuNqS1SeH+kZzaeiuRBqMM
MFMivQgerwMq0hld6VINv2t9Zngo6nQY+/nTzLeZbxzJ3r9JwgvwlNle0pruLEtc
tr2wWNyAFEob7KvRKVHvszswAP8wLSt1hiN3dBEUFndbMC7WkslPT7T0i/eUT36Z
+q4LZSzo0b/HRwnXy0/NISv7IDcwL3u9rnnm+9jjr/Wi2YShm6TKKJMW5X09QgEw
rZQ3pCnpkzgBlWQsRYmwhrynAogossNKwyEm1hVDWgqgWU4WS/7KQq9nFm3HKnfz
EBICVGhd/Kaq+s2PcPHIqKu4oBMSCPlK9EvWNB/xgSJWmguW6kh3DS7cwI5XjLdI
4jWKEhl+TBDnl4v8zNldaa6i91s2MJAkGMOa4nZDredsNGue8NWpwxa7olSCIYwz
LCRf7+6u2M1KuE6qK/uByOUB98lauT1wUzieoLsFLWP+05SDh2Lvzw4vOvl33UiG
lDHLV9NgLwq69nfAB4+w1OJ+iamq3Yp7c+1RCNUMj+cSt5O8d8k/ztJmSyZeiE1C
1AdYKD0wxRxXb69Fi1pg2A3aGN3dfteNKh+TGWdQQJMHDLU8CloLlG7M3l2FBiSU
ysgP3kRwjxnBGFVYDfe3T/crd/0Fn9lnwXmlbqrqPsjbEeWEpY8TiN0bhCYnNIdg
UiwOLbjBwxpt3cz3eNI6WS/XvpN31VF2beK9zchdWjgYTBjfKU8dbTGcXu7fpXZ/
6t9+Ya/c9/fidGaf0CDpGRDhqvkwD/y3+y0IHT4XAho9nffYzsCD/zlerEceRXuu
2LA4fSVTpQbEVp4clJxzD2f6pwj6+prfsGDRuXRvm+e87/X2FCkTlOpj6uoOxYRr
Ohsr41hIsQoBzfFA/MO+9jqpNzQCcppaLnA9XgGy0GEK7PTYbvJiS1j9Tlr/CWh/
L1FMne+6xaNlNR/xwovJd816JL0gOCok7gvzV+xs3TfL/2V2dw63S720sr5y0z6z
d6xUKRmAXKu1gEeK/SYUzQiUKjV7e10RXjgIYBbplj2XJBZ+HCXOmCdn9hqgTQgs
4t9lEgTHe7g3gT8OWTNIXit4fX45OYtk14ir5xpCBEQ99UGYcjLrok0jz3e2CDB7
JsEK68x5iA8zGEg3XlwhL7eKcG4nTcRmjOOG95h0r3S0VOodj72p2YLBAwzq4NTI
ZnHr/eLnaj6+P21XSFDeCTVZo410lYEgZJ9gERFdIkPP1mcRisP+8gMKCr0o0S7S
PmzP0hlxZUNZeqm6Wm+MbiihjlXzCBn+XmIzT6szTYKdQdShXiYfr8UlT1kbLNNh
LEArwgHKrFaIt2Owl4cJ1ZkJU09O911HNFbqSsro8yeQ2xGamfMfjWKTVeByCDzy
sT6SkpDhKa9Wsh8nib9AUT0eCdOfGIHYr2909wUgaaUuI5ZYRZ5ieUARJGhM0+5y
Ka8gMUatDHl+MD5gVNHXK9q4rfpEm2F7ef4nJJTZj7AOnn2HbIZKdVjwse7IGeDZ
ffzO9yAluAcTmDwGGi+fkNZWITl2Kk1EGf7ynFBPswwbh4rI8dhs2WFuQ1J8nrmb
qJGr4RiFcmwcprPrEvmrcFjSTwpEsiX3WPqxb/g6WyqlJrHxahbZrny1m+pe0SW6
4XbN822022eojTslkT1h9FQM7vHlVT0/G8GIaklRzDdESmWTNctk1aALB1VlGyBo
I5ZqwU0TmJXL2lu78N+IFBsN0OXzKe2CuJMxvENb7H/ZtrGeCq64ATVMpnj0I12k
KZSWHOmiYodpRMMcV8k0M3SNfnXj5W1iBdNamZN4OpIsrggttOeZN5ygIWry1v3q
5PGgze5QT3YFN3wrDzwqVS3OHysIgHdWWXW/RmM+ofDr4+Qj6Dwcj9QhkCnN67kx
/Tk9FM4WHig4cJtSxUJOwdpnelEXT85LkrixKCfr3ZOisXQLduqWSfgVNJ/Cxzoi
ZnwA7sSzK51+pRpBCKGabpYqo8rurG9LvVD/0TuCEpQVVGI49FRc3xDZlw09IFs+
Vw2e4KQiM/E4nJApu2/YXkbp/vPiih8fiUSYVBYmWCOc5LslaP0IYCL0d/25vs3M
j6AOEJYz8t91JzUiaC/NL/HU0sWANNMkaFXvBhcX0NX14hHzr0kZnLGCfin8lskE
UGaJ54muD3AudzFEen+968LTsI8dU6juzdE/ZFib53tSYYqRGO/8kdnNBCNfR7jh
e5vQf2+jZe17AADbPcrdGIlx6cRSDnDY8jewmrqaruUrFIYMEZqY/MlNsqZ7wVeP
EULPH8GtjuYYytPi+BdWWfk5rFpUl+Gbj9HHA4yabCxtHeu4bMYEKgn3yqoAe4mg
fLUVkhsPQOt7e5LEUkFrv5m6yDeMBVPK0m5PK+6vbQkqiSotlr1x3y7NJQWmpkza
AQWgPRiWil9r06/hap5Ct73eDuek4FGnIWHrtSb5WxkMFQz+gvpWPzM/Sem3FUk/
Jo83hxSsoDJzAsLYpc5kO+s/T/JiRViLX47IeH28Cj6j1cTQ9VoqjF6oIYbDiKqP
KWotS98OFInDSVA6R3HR+VNFckW7Ul1b5roATGOs7K/SKNOuZjCly0PPsYQ1eVi+
7XMWN0Bz1geGekex1QUnW/Ja1WgJgOiUvNYY0cY1sHNDy9U0esRJxojgDBobY1zl
3+D2TR3F0OiyDDwMB0yVeGdyAOpOpYjIWE/Jaj39UXveU6DBiEwEy1rK34Nazkdb
2p9f7ymSWjjMAwxPgmrl2JMp3lv45hO9iivQ5g3nXSNoYcDUG5geU37B3tRD8sKE
YtiG8Xe8ql+H9d/bqFqoQKDUYsCL3ukMgMw8r+Kksg/lSq+jzYlL65Kw6hcdYAqr
xHKbtP2exeBqVE6IKsZu0nCIDBcV7Z7nEmkW4GfUulyvn1fNJmH8NT9Y1SHUF2Gw
HAr5Kmb5+jQdKBEvzRHNhE2d4AWsyChMON83WmCwzjX/NfMFouCDoUxKkBFTah8r
mnJilVCwlGoPePMBRfQLHyT/6nS52mbZZAvkFqzC/c42Z3nJdMQTUcA94FoiMwwI
8fGD4sUu2l1IumWnxgHj9Wp9i8x7exiLLtvG3U5qCh163zgMl5XmARGg3bp8h8Qf
/i7vW+qQfblpTKFDXU9e1Uy3kfIogWFfpGCWpELuoB3mZz4jjdPGECWLoVx31Ddi
ApbzRlvG3xfM6ySh9O2/eud52lc5LPx7aMkJ/f0zHYiU/2QMsVsjTopUYTiapIhi
mMQpFeGF4bbT3Qyk/5htqUtbN+1BYGMLz94LqlYACwWWd9U6eMpPf2EhXkeSUKMp
7PJn9c686q+tCwzdqXPOithu5K78nMlops1eYMuzORvtpPlvXuUD/hCN94I2q/Ep
ZCIpagdTBJy1oKpHr9+MH1VrYTGee5w5HDF5V0AK1aVHcFKt5SEGvebXDZF8IPPW
gpsjJMxZSX8mrGUUiNAgbwienOdRsBCgeGUdDwgIcN3Ec0Q9+gcYDG2+z3weCyg/
bNGkksZgnVJHDOsn/zYK/mkDSyhzCGTf0Nym29dof81gV5aRCIfeQVHp1xWCfvbh
7SMbGmBrI7P8/Up/KJkDzwmjKGilsUhazK1sPeVVb15fI4puolWaHTzUaLlWAM1y
E8MANWQ2yvpeZt+kS4kIcsuz+KDliWKTow1L3omXKgJ5WoQ06Pt1SRFRPBjljLL+
dNi/BLBi6AGTPFFN6uHqMfTGpWIo9FBFhUf0wL/GyZjsatsC3VTYUe3SZ2oexx8m
FvyrXjUMSQwIrOO13tzU2kNth5tq8t22cxljLZr6s3UnAMyP94kNYkMgw0A5shdE
0SGw3eUcciLFaRmMLeUxl/VPAlBPkBVsBgXIL1Dcq6iy9RRRsajwDX3BY486Z8d6
HXXbQrOJOTEOtrd1+xjYto2D8dieTcxnltnDyOPkzG+HEQHHhGLwa7vfyriooHkQ
tG5PHj7HZW/S1UfML9NiHShMdcpnXC/A4ketsVNU5Mhmu81vD5tndzWcUk+5icrY
QsOBekZQdyJHfZBqzZAgo7x93Ezvp6rAjlvTmO6RQNQ10kuAEzS9H9sI2Xqpvpo/
/lW1lRwLtuyTucWMU3yfOMZdNOLcIF8f1bCb+BBLIQnP33o+oBAX0XubQEKfnVxT
3hEdHtdLp1IguPHEexe9nU7A59DBs/Sqv/Sl9y4K5jlxVqTTEEGK1Ph32otk0S+w
q59KHcX5YR03nfKK8qxblXC1rZp0Ng0DATUXlgc3M72CHzXUqEdNPL7OyRMVuKfB
zqQ6GpfPDNAfzhCy44au2Q+Xg+LBY1FirAF81EpukpklR2wpprj325eUsszU66lH
SeicXCnw32S46kvf7ATN9StpmhNKZw/nnDD5ZrTFyUJJ0K0YTupI5vUwNLD26Wnq
D3nPneG7kzmq2F0bPylM/RemMt3EjiUe/POPquXAsC154zmqZf2aXEDD/+JmVwyI
V1SvUGnhM56oy6mKhiu8vANn5V+q5+/X4p0frShIHH1xdkzQeeLVOBZduK7FcIyN
hcXAkz+zbWz0/kOfYmg0+rAiqI4top1gq5Fdg38X2K3JsKZngHtSDAAR/ZwBvNsj
dJ3KKqpsH6VPOJEJN6Oyk87SdT8g/alXvu8AeaRM53CjnNRJKIhgcvafqesSOY2l
SxSeGQYPvFFg/OItplkCAvJPP4vpHTfq071jvzPd9CsbeRRin3s4w/nqU/CTD6ZC
8P5WZOn0nz53YP7vEx/SQ+7aXw6QLii2DKTLTWQVDBTkdYLwvV2CaESSz3nSZ2GG
ovOWIipWbPUe9S/CLHmIEu4BT6QhbGhAQG6od3Ms4MdNE6Xvt7e4FzSqx33FqWiJ
J+4TA/r4ZpMuUNhvYeGuu1HyDPAMz9SCLsnOFJ7rg2exrCYbJuQXTLA1Fc9ZtvjS
I3sAyyB78H/axnaCCvRC9EXTvx0NK9M+eTpJCeL1tavw7a05X5n6/0gF/Ln53G1H
vp8g/i2JmkA8CU5GUxs92MtEd4ufw1mGoANOCQT+zZEXFA0fY3z14Z2nd4B0hxj1
k5BsqBxICJAp/dJM0fmqytjyimKAAx1PvcNKMJtg6QNxyz/WKGVNeQCepSCJQ/WF
MfVJF9Y5C+gWwuwNQJGITZ/J62GEhT7uCDd+Q3jOF7JlPyvjAe6bGe2wfG7r2skY
3UlGPZLU8N28qrqVR1a1l6QmRE50Xes05RT2joTu28nICjBKDz1gfv5zYKub/LGq
c8fYVRsQDR8H3gnvPI8JHCm1DtlYes2SC/UQKyJyz3f3g9M0KiTOztSMe8vyxIJ+
bk/lCcywuyJsMrVayj3QAPEYSKsmIOgmHmOCHGe8VfDhr6ExzfUqZQG3yMwZJmMD
oDSKyCaenrNHHx23A5STT8bQiwV5MVQI6IWr+h/n4qRYCd8KnN8LWhrjR/0bCe/W
V2goNeWrVhBFnONhIrWfLMqvlX/LRuzlgQsVkMmFlXPlrp/oMA4kvifyKhTTmIon
/kJ22bAVj0V2sDIQb2iCJUmPPh1h4/lxbdLung+jZX05Mu97LMXRPaq1AiUgtmHe
gAjYPIGS5XjDgQ3L1/cz5oJh0d2yMs2XV90VAlNyTesOsBAZqt6d3SO6bjc3epht
ayWWmlT/3P/rEhXYcGPii32VqvlmhkMx/F7hrKJuNCXjCThv4zdpkJkD5QNzKYsf
e2FnJPryrqIGdC6POM84SWcJpsC990aUJ3gTNZp8CKzm0QADDyFQEcTgElDYRpsZ
0io3vbJ5n6k98y+mF4ghbzbA6TuPqDY36jUYYtAGxI2sVbkbIqA0muhFlw3iLqFr
GKPlRZYdslfpF8VyE9UfgobBq0CwxskdFnzvfV1oxzaEGAQu4UkUZ7dqGYwF4vIO
qet0SSHE2Kv1kVggAogj8Nq8Ho59WatnNBMQUEW3q6RNa9ykfT+GSTIeGJQaB6yy
fAcxwHEBvKqv72VjFDCV7UXnb0P4hLF0jGJpGqlNwu94PnghUy2YNwq5/vCJyJ+9
Iml2zQBCe4wgPQpa99n/L96Gml6Nu04mlASRS7tZ0hHcNvAPmC4xkAQR70gMzyHO
F0YUMdRDhB6jqpNgQElae9K32AM4wukSMSl9nX6wS8epps7IVwygSkDTZrGcZGRe
cnCMc6x0539hIxmAIylkWxIK8IG6UY/o3C7efA6UFBEG0x5vpOgSUtOFN7vkUFqp
UPXKZy6fw+ok6Jemkb5lB3IYUpsXeijyQzsubIB47hP8q9Hd2wjrb03GvEv1xmsT
/pJUwPGExYgLU/ousq56i2pY2p+tiS1g7j8c4Qn4sF2Y/ll7ISLJPFMUT6RUdZLp
8yyLn/zpqo+CQiPF4EWksjRiIMKEKkM5pT8z5Au1lWJw1PDrgz0bHM4BiO3qGzSZ
5iYG8poSms3QCB18ja6m/PKvCUgODwz0RnNKCFfy6iWY9msHy9wTtDCDksyjGqfC
k9rJIUtt7E9Ev4D5OSC2EQHtjbNum5H0NMb3mYHQECFjCJ3PSk4D12+gFZe9kLo5
V/aXf3q1FgLxUNtV8/wbu0StpBBCaM3RE4KQhQhe6n4/M5kyW47B4OvcGysukt9a
LeCaXT3A9GjGSNjSZ71yIlG0fbyGfXsXScFESXIsVb2a/oKANVwfjYJxCs4yb8b5
YsOP2kiNKD9dudBEsoxiP0AbNst16zNiERIw+x15BsI4X1FIENhXF+p0Rms6SmlD
GhewInoBoALjUodafrir+i+qBGkCNE+VnVO5IPkpCb2Xw/yeSKhuxjrFu7JyeNfT
tKo2mVND8PCNe74KVlvCA+U1GkEWqXkkHlFuT14Ch56WomZFXrk3RnmsxtyMscBO
gIoOmQJBbKgZOcNV1E4s4SugUV6tBCLnuSgJsVIukPM8HKN5Othu2bicQJzAZ+hW
VT/LTsPbFPQ54J/JpYDVV691Au/DMHMwgCOjr45z0gc9XTKxVTCLAwynCRj4XfpL
HZC8vBSuwX8JiZYY3l5bJIaLR1GKHlu3W9vBhYyw9X+E9ATFOZHeo2LOk83J9lke
YuoKGvaxDpH+JmdqObzF/mAIcnPsnkYO8y/KWaHcQCSNoYGiPagMcVqDuiU6nDAI
yrFKOgVZlV5h3VewGfIGkXuV+uea0xtBQwiFl8wSE+grmP2hl8qHjUDMgc+IEtzb
T2UnjC+KmK1fDWXf+v9Xd5N9LoWiLQWIrfw+SakhCU6UrFVcmCdzficJv2XIi0iN
iDPuESu2txqS1WFFmNn0a+7da+MQCWNEPOrOW85NkRzTD+7B7haNKSfsRCaGEZKH
ilr6GX/XLc/LI5S2NyoYPhKDh3FDWpq5pKF1h4ubj53+yPJEhGcvVAu7QzVVZ/VI
dE/1cC+8fIGA+CRWavSg9MDraehM3NIr7LfWgkRz1YoxzEWDBvRsz/fmLdU1HH7s
JqfKD+eSwIDT2bv6yG7zdWQkEUECfxXwc3NqkE/bNyKrMXokblUocrt7mWwJYKFw
VA1/OjUuSa2qqhuSGEKmTKNJq73Pt/04nT3tshX8kRQZa3e0b10s9kdCTG8QE1vR
j0MnT5M2k6tonde9nEzJ+P+V6welKUmpsBTeERWxn6MtmzkmqICwY5xEPhv5IU+a
0zsAFCpEdex0i7UwFqw3yuKlX6xGXciqeuapolr19nAKFzVtHok7YpMOsgM7rQuC
MZZy9vomlWkmkqceyf1BGm9PHoSgGRi090C5kM/UJrxhoKcBjO9fHVjlk7O4sUti
f/LSFe+DfTF8OF+FX1rTtYR667QmbsGtQeeH56OFimZnaymq6+0e7+JSJyTUUUNH
sKrLQ1BLYfj9l9cW1LUVKk1avIcP6s58x2sR7LmfboAGK05uVzTcju7odDob8T5T
fgrozRQts+JY8U1wlPy+m092bNNz0I5E6OiOuCEHkYkZOcElb9X3AK9/4x4bGWqS
w0JR2X3ihCLslNWJpb1xTI9U2pRQJFZF+byOF/cClc9WMJWq8saQ1P60BRNxEwEo
4Y4sQCxYfFlIFhTyWnviKEUmuqPm15Sc4rdXJmyUNW631PuCaSZmkxosoEGEQues
5bYjES5G9yUwEorspDy0n736QqXYbGWjqCmFgZIdoXcNzf0JwmU8+QZUST4ZSmOr
0WqqrdglOra0di9KIUDCE3KzdRZsoSAOJc+4SXIYRec98XXJvnmuEt7QE+/NvDXL
LZ3hgszTu7hu4Xgwn65ua8JyusppW2/osdjtQn7Fq4m+Sp675hwqsWX4sIohPkFW
AKz0EkU5Df45lFhYNOwN5/L6U91z5ka4XCm1+cxtEV4Z6u/duDm7oueCd0Ry/+hz
neuo0Vi36TPXqqcs5q6tGbwbm8mRYssT7U2FPQMfsmq55FK7yUpcNIRuN0kWfsPy
AlNvuM0RdRZzjBwO3Pt2K/jPUQ9YD6Iby3nhEnBOmFW64ROdjr/N3m/zfBprBmAS
zCfwS1aUD3/KngpI4vaaLVkkjCdTPJK0j07+XNYzyu2FfnewZ3EtZkAKKzi6RgSe
MdAfedWoUdTf5w4zQU3bwHN8egbCuCnxHhlXy3tQjVI6H1UwPFBhLpI0588Sms2Z
j1gH6oNs2vm2DrYZN4WMgLBP6XtXCB4688u48IJYxABbChEO4LwFN3SClIyvK7R5
QGqu8EP1G8u32QhCEQMOnts7BAWwdvYxLVKYWZwcfPyxr+B00W4NHHJV36YvqRiy
0+/lkaA1ecQ6Fv4+/oLs/MCEpRbwhLygJ07rVODHQmm9C9R4MfunCg8Ev+X+mXEm
q9dh/T9IsFdoMBS0sKG3CU+gpmULFc4U66ey6cEl3jalZ8Xil8jCOJZWHWGZkxos
CoG2BYEbv1FVO5CoIomyPd33+odVjL9YGLfg4Qfsxzersd8Js68zRynsr7OVokHf
PNZLu0tdC9vLeI5zsgBTiZGr1J5e/YJQYTw18ZQ4yi90c7QI2+FzWJuwM0EcD3T0
Frqv/KVh1GdvlwwKJs6C/DbQ2QCZuY/ayjsKhJl4SKpUg6ZJKdtpz3A8yqom6osx
5O6dBAMYpSw5EO1OcRD5xGmZgM1uRYYUD2cOWUvPJHvxoePDXMsXzfN7TYGKLwcP
iFGqzHLrSAa82QoTLtEqtJ3zLX8pHX8PfzvL+frEFTysRX11kEb2UGlQ0hbMoWkp
HL5QH99NEvPNH+UHNKEj0ib2WcHCPqUbn422PYGyfDCvc+bxQlDLjOuIQzyhD2a9
beAdNPEEtdjIdtuZqylYYmGbQo5YVESWcD6+th+0kghSnqVKsbaINbtNYvdwhB2G
JmPyLLPiF2jZ98KyY392fZSXVcPW84NjDX3sHsx5ni8isdk20LNUI/5br7ncv0WB
E0pqe1oUqtbRuU16/lmpXHfk+7mQ947L6xeulAK2hH4zykr7mHU1uGS/U2Vc01Q9
Vwtp7tlN02+RXqcvEKmDKDWRyCR7L/4HK9xntwIIhDnPkJYUXtgBCV++G0PmB7p+
e+QhN7/x3q/Z03Do6H0+FC0Un3wOAtQI8luACBWy5XOqbKqPHm2446e1WuBu9njc
Sos5lD7n5I2vkPEm0Sg7k9EI5Q7mU29CQCeC08lpYsBA7nlUef4Ca8qgTP+ig9OZ
rH71Y/VgBZuVRRVAqJBrhUvyLWI8W6zeMrYxr9AwKJiQId4nMT14OYj6cSX5if68
cg/4hyfzrHh5zuj6a2Jg5ren8QHrN082h88SbVfcTWsJn8edF1K+u0l4rQCVHcCA
w3W13sDmz+aPZogrvkxGQRApwQYnN6EunWDEgsuTUA4X+9p2lpioVJw4tma87z6b
XFB/auRczE9Y/ZIuDrr3Cz+qI5w7qM0KepXDTC0jBWzTgqXac04g3vX8gYqCpUIt
EBiGJ2sSP9xEIKnv2WoVNS9P2eHXKmIn0AdPBh+A2lhxpUr1ESf09aAqFkCEIIaj
Ys/lsK2tZNokyTU1c/vCTDxzzGCmfLZwmpI0RiSfiPIN94krHMJllgp9dOnyaBF6
8rcC2CxMO0j5M2dxwsFeVZ+O61751HjbMqWu7jPGgxxinDbhDW9H0K3UYNajE5WB
Vb08c01du/uvCkA0pW/awZn+r6Ur7SZ9bL03io05mRCM270V44mHeeKQmP4+96JR
H43N9UNHnwcJ2WDf/t4B58I2iLdDirY3HomwGv8nz100bwFww+QjFJxRfQMr646d
0v4zYl7qov5iFbHBW6SZyW+sljrHmAydRXTMwlvRlSPIxYgZjMxgM+ol9laPU+Qr
n5zGa4xHkIkfW+mhgSDaNIcauB3jp6uepwtGuJX5wWke4kjKp0/Wvxu5RZVtUVYp
/w0vLAjOSsJLTxZdsuMito1dmyXYB7+UO8ZzHpJuA4UTlQ1SkarAcmI+ejYNcUbB
exNOe1v9n3KB+qWX/pRLNoc0OuxbA7xd13wHQ3+rsvo/D8lQvUSlT94LymNiIw5a
62bOm8Zxi0i5GDWd/F/5/5FGyBRh4mr5trwCzv7Ilk2JVlMrJoJcZr5P/RgzMedj
OEMW8VJxI7NwKqxJGQYtEnD12TjAgKHsjR2+cq8VF5k/auVnTiUszqy35Iq5ekEI
7UV73N8JabfSyVgQNqdBlWHBJMk2/mLlB8jOYDqS/jsaL86q2JB5JqUNj8BlPpXh
Xo/vs1NZqhgIoGD30ahOrn0UDyi0InQxkiufeEx/TuzaDRK6akxBFY50LBZ4o9FA
aFP2eo3ptgccOf0gjffskz+vsR4ZnjCLp2rNNYVQ6H21iD/i38+sNP06GSHJtjSG
0j3M7SjaSdzLSApVi7ZCcjYO/IKl1ydCavUhsukM2FoKMQYEStu8Pke2ku2JCS1g
MWQVYSdTnqEPYLS2TrlXezFOS3XQTk4yxyxaVCLDNQxwBBx1RElzqC/nC7E4C+9o
9hF/a9hbcTjYZImNtY/0y++9Zy0L+RCYbckqKPFZgfIIkhMiP59I2ILBJ9Svf30W
0peYUsCGWIA073p4XeMQO+zRh+i6fUVvvu3rp5AqaKgMJHKVQYJp4X+tsMkNHGKH
MMZsmGmmS3qw1l12Om+vPog5PGTRfttVIc6zEkbS72/YQlumlOl5b3W8q+1ESZKi
a/uZCtn2hxa26Ib9r5DV47IfahC/TQBnCHHsCZEyynXHjZDbTRK8LGBCR/exPFi4
tbSZ649Yl41VunW/90nV9srNQXCA951GfigG1nqKCfblDlUrhZj1c6m2oqgygUVo
Ne2l00mxgfklNcneM4ZJYVT4jWvoQXem3f7G+J+w/fzRQcDnZfX2B727c2hjKkcs
tseaGfbNEKCFjCXoqpm4hPmc9UR8xzFA9sJX7sZRphjqcUpzQi7ZEj3n9DEzh+E4
bqPTUaAQE5kKnbRkHqivpA9NTMrRZ8H2jdCzUhE68k2Bz26U91DVNKo4FEOYfRCv
hJr2+KI+U60INueoRZLFuAvMHOGzhZY5jn9GdoXEiPHzFCCcfQzkgq9UXcA/LG8N
xbsjgquQYo4WCmNZIMZ+d2O9+wtKQfo3Q3cZBF0Fi6iS7Qq1D20raovlCUJtFNX9
sL1iGMfXSJeMfdC06aH8+ArU/0RQ1CgNuCMumVfBrO6UVSi1f9Sve3A0D1ehoKZo
7Sq5NavDATvJlvZ5S+IGOFgx9omoftWHRM36axM9thjdEW4vD+ESBNEKqMOrKqZx
+rSDQy/bMb/VMnIswC+b2827QqivxSDn7gX6L7OBuBJPI1sFi2CM2l8P3YQPmZPV
fuxuFINBgvH6bOv75U7V7QYa3DLq3SaFJB06T15KSUD8Uvwt0E+jyL7apWAxB4pP
GWUsL4V3bhiUzdiTY1DJQJVB7RpvFpEn+2+0846gEmE35btVSzpl1PfcYtyQ0XZT
iSRH7ND3bq8cF6JkScNe3Pb4NKa0A8XraZ6cIIRTRNpDMko63MblJ8wfRlBoCV3f
2QesY8fbujdYptxX02C3/HyLF9aVZ1aV5Q0/7irDqhw1K9lcOzszR7pQzNMk1hto
uSm7iFM0344w1hElw1JC0VwzptyRJsJ2+Spt5kinCHscnEHFc1Pz2NEyTkViaF/x
fKQMoACWYwFZWp/5Ww8KiK6JAAzc7vupZQo/ikJXIlOzUG6jE8z5jW704fCLHJjg
D5c9KhYgpGWyMoMPbLNms27XV9YtiPeT3jc1ePh4Uiz/RhWdqFDi0mdms+AVi5Xz
J4PDU+rfz6ashYOvRt+2cYxdexpmZN78p2jAh7vXtaDpMqo2Ojo15WcQbIP7mVw7
3emygxkzWzpiftTUIRdT5QSJLASxIRxT8oSFd6zcKXiAI466JsLXLOH5TQExhE6z
Bo0hhfyTyMLILO0pvxqOj6O2BR5u3CN5htJ0iYrb1w4T8g3ABGeX/dcv2QMi8CWO
84qWLapXH0QKPB7rtA9mvA==
//pragma protect end_data_block
//pragma protect digest_block
trGpVpp/dkD/rOGfgUSh1+Hpq34=
//pragma protect end_digest_block
//pragma protect end_protected
