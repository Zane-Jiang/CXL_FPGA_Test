// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Io6wDCJ62HRQMZ8DVyGTDVsljbeqldg1vSR3TRF2ZIFeESPbL9CHPjMWIeQ1
vU9LHNJPtFCyo/LnEdqbwDgxnhQGjTc7CDgYnLJaPgZCsRXfCK6IjRRBxwXn
+wtCeQqZzPhf7KC/WHI9d/YyzIfRmuX3CGnAliLWwMiSXWQdEzUUu5oKRwUo
lkSNmuEKGVuPXNxuMb+DVyNMCAHN+9nQmJ3hK88DNy0AwlNtiOBGc5LYvoPe
160dG3bVtnNYmJLnc/SmPhiKIEC4X3t6jq4bLUwxb7qyZozJ3K2v34B/uwUh
9jqsO36zHAHhC6YcFMqvZiyne9kKNy4jjLQeQwPqZw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LGqMfIYIZ4SeuL4vekdpxRYc2Kyp9CBFWpH/q7rzEN6hCXCP1ysPl/Gno5Nx
aGVHFzi1+vXBDEM9eIErV0ujTu3DmlHpupbtbl77ZOw5OBKD02RL2gN+/UWQ
vFjk8WY2R/gP4pBxJQlhoNRh/DKWig62THcqxeAQL4KntWLFZfIq8a7rnOwc
EU6OpqM2CseYrJbppHbglD8lJVwYmAadDD3ieFiJuEo6Im6lz1ItxhCzQSyx
soxtGy4dbjUEKB2ko9ksiDknvPy4LtyVW4a8pTWmt8QWsjsHVCmDQVgOyL0G
Z9ytuY1t5/nShgIXQ227Kv+k7Q6xqiCwYsihOm0T7g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KqQO518e6Iu6Fdqbl7YYdAntIdJs+cOlFI+lmjRvoALn0nhzd8Fziq1VzBiP
CT975M1HBqR2GzpcQjsZJMkSbMo24DNdC55xbfZyrcCPOhwlqWdWoY68A53A
LPI0tr7fHRJRi+5fQ1lYga+m0YLWGb4JSUQrntVjYMxW+KQf6WXy9uhNcfKZ
C57gZ5spmGpVjAWNRbBTW0U4BtzWNoq3qsUEYoG0SqNIDjiBpTnCBTySzxUE
kx5nE6rWO2rjfezRVLzyWMWEziJs71s5A0EO9CJ4Ri9tW5uqUR1MklB6eGFu
SXeG7rzDmrbSgjuLB2Ta+mNB0BSj4yst9dXyJ1YA2A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m2XBOU/1HOw2J4bIsUq8fencqExNSVO35f2nztnIjrRehoLvI+NAWIBtXIAy
ZXjVNb2e75gBMQS/WAebqOAZWzvPKzS4lGs+7DrxuJrx3eeaJ6ZzBLHUwvng
BDWcooGk0rO52XyuBc148wmqpq8LinqewOL5VUjDhqJ5DWGyqPM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mcnMkRjNG2M4kC2zQk4ej3zim+2jrMxxZHtVFuuHs9DK7gmzT944g84G2gXZ
92gD6WNeFDhK2qyA3KBxdsmpF5eb7V1NzvWuUUrWgXdC5nSiVqZDCnZtW4/b
TQwBw4kyjrZ21rUprZoY3DJS2Exv1IJdUiV1fiPIMbqQ5d3lhFSzjc1Wf0XP
27Mw/YRMyQzqCzRNyeIqaSRgPlykqs3zPwKT4mqBF0t40qH27HRYBD6yOiMn
fJjeI31BLFwFVLL2tRWz9FcsFZtl59KF50sDxPrlm+TWKPZMUFzslklHLaNf
U2QlS+nd2anyNJQWtnuzsVieJBm4DpM9DnPRmYHX47zOW6iOfcwB6qhoKylY
FaKkgaKRMgMbPd8vrR2hwRvUS1JPiYXxas3sTYTjjqDL2ygI7nEkhUSlYV5/
jRehIp/ZTVXXiPcD/k92rSJ2gA4ub1E+qxE1ZmIM6J/EjeT3aJc/GfUMTYG5
efbrj3eopKmC3vwSAO8J+PB42aUGTc9E


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sLPJncDZ1hoijUeLyTHpzrRbMjB1gV+Z2wSYeaFfEZ7+iKp2SToFAaTXSE2a
zeaXRWAgxseFUYis202kWQuev6qxhWWPewH6SzGoqbzP6xkIQ7x1pmchOX8I
WL1CVbd8SGlNuL5BwOqM4UvPGPy8RTrrJKbvJJI0+QqeHRarnAg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rvNfv3Whm1cdwK9kOaSh4FD9W6uR9dfSP7pH4Bp+FiTFLRPrCLgLxlvV+s0r
VqL0eue7tU/nTbtGMGAK3bUBmX8bTScmdia2eU6oheN8t7j04xSn6hqmqz2i
X1rPiS3XvWM1n+9KUVHtkYB+wVOxTSDy2bO07quyFZZ3uvsyPLU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31120)
`pragma protect data_block
7XcLCwEcido/LSL5VzNRKQyBZFwUBcANc0YOImeLir+712diPiGng5YqCwOJ
3ao7MzzVlRCggb+mpb6UnmIXCzOV+0epJ/OSTsuyigmwNxoi0ZdkH66Dahyk
b0+QOj3+/Xgu3rOIuFuGU219LE6a9CXbjz5Ab88FGr9nVABd3QnJVN89Nu+5
SL4DqXdx3Dfs3AWy9uwMg01jwanoY1GTdyBVbrfunlsmxZPLDIwv+mcNCsoj
yDU1+H5br1gTX5LsVLhjVJCL8scflIDVPdW2QTuAZCHG8dLEOkd86MTBRHNN
awOvzhQ2y+6PlsIceatH5CvGaZ0gjtUzWlAh1Lmq5Xdl8iqXSoslJr4uyynS
dgNs5+iSNzbZ/6IZIv3yyCTT5K+hRMnxxWDUN2EUQEOXMG2ls7gUqfhuCpcq
pIpzV/vHsDTPlCYCV2htH4poebEUNp1AoXBlijk22FLQc9nOlyzHJQhJ1NxM
eV/e7gRfGANCSYhZCgxCfMYGBH7z5Ad6oEqit1WYy08G5IwtBo4jFXfVUQ5S
eoZCHHQfqOMydFVVqwfiRPFjhDUehMeuf2Q4GdzEQaqnFswv11hsAko1HAXI
we+A+5UbFFFJrijjiDKN9jW+VuJz3insNOnNLf9e2XXZulhUksDSTHv2H5fZ
vzk15lJSZAS26gJ9aQxOy1YPkCfVUsHhk9tEFilK0p4wqBpRI9b/2F9QWraT
GHhYIkQY8/rUkQSHbbHhYTe5b79Ii/LsylGk9xQbJjC0dyxTUXH42UPny0Hz
vH1KI/4BvgsHIXtIIFBy6nycNSnCZL07KoGO/5waZtqY0fvzU3Y5SQ2RadCh
04n2I8XANwyJ6yhqQmNCok5AZAD2Ffl8sMvOgknfbfK1JMQS9z+geM5UGhQC
YjXZ4UlFx2wrbQ7eiJgnKpvONwjgqfcqt8UT4KtB2FYs/Wf82Knh1hgTCv5O
BpCu2EoSgMoajGiFXf9ppSxLmGkvbw5p7bfqq8vWWZJsTNsYSfbCJZOXB+dY
ykUu+Z95/fvu7ZsVHRgx/mQUhTTkEViuFsgGWkdAw/raita27eWmAfD6qngS
ZEpNvktxeZgsklqNBUmbkQjyHdSRl5XZZoDBgKm2rG0l5z7H5yFfribfK7Vx
rtk22DXvoO32S/1tNY0WWvaFKL1q9qYADFTke36sxxIC6nwBsk8bON7fH92x
qpPbZdh8CJnx0Fz1JHYOTd2uTyMRpnNTvw4GkNKJoVxHQQbRu+AFsbSbocug
wvcvcIKzFn83EVlAkY7RY4StGvjG2VydCiE6CGdQ3vXwqd92tKnv1I3ce125
elKsLqKTdAuX2D3+xyHfWe9C1UjMGgBa7iOTGqGg+pXsHtvo7r/vSAvhC/BZ
aCHETAABICkUWqQ4QOS57tnuX3FsHeto9V3KEaH7Iw5RAWU+ChqNr8muK0uw
7zwMNKgEhTepAVv3fo7j5aPiwhLJDwC37G1707XCgXKIZwbVvxUiP+BZ/P0c
QoZJ1OtSgcWkrNQ6YEAYxcnE/d1qazsoR8UEX1ntrlIebNXFWE/pNZRC2QLc
vArtg2kQULxBu+BoKvK9cfjyQ8cNmB+RkOiTM+v6lyJrWIrmdO0q1vJ2DEUv
HoBESJFjz5aYtkISBBe2+BrOHrwOOYY7iG4bA3/ODI4D3WR8A7umXMa1C71k
n4SmEqAg8HtEC7kYWHSVHvn3FQKU3LOPp3Oqe7E5dmlt80YkXWldPACGW8MN
C5LuIzOlbeeiBYcfSz3T3P+jaEoLmjQuv2N74XwOjW1Ue76TuvxFTAxdLGqc
BLR+28DUQ9jounYQR5JTG+MyBUUphdRrHU5w1EVkX9ELPRTkplhsymL9h5Ij
8ZIDumoTpcwz5/rRPoMdcXcSw4C9A2IA8J37O7pXuwHzS+E08RW1KHaN1Z1H
L6XuhkwPX0dP9XIBpNlJUhPOtnk97NG4Scxe2nqtwqVLRcaSPpZDDwrzKcu3
FJWsSe4xEP7zRTjUVY41HRZW5kt6Yu6FVpIIW3gaUJEl8A4MNPhr2im8EpgG
LvdaseiKj8hMi5fAbBV5+IehHE7EWtluuvRllpY2ATPePb+5ghRtfQlKGKQ+
es1IpSxaBNxLsh6jJ+fOfEtUBiuJWR7u8DX4aNSpKW7gKXl2stOWCNKGIylx
dY7b0v2V0YQDAI+pzyfFtyZFIlLdifK5n7b1GktGsMuVjY90Dw5fgvu0qtDp
gmGw7bu0OS6A4jFWwBG4inQzy9GLKe6P8z4A45zaGS9ErnD+FmowzQNHr4tr
amtcxYJuT6FnzaZDE4t12gvP2mnd8hfKqMO7sQJMfESEjuRhz0JmLwoeULCq
fDznosMF4MjQiFpxBskKiquUmHySR5L07Vyikjzu1oxSoIR4mCDea/4EzpjN
HCj58UGIWgVYNeukzVYu5xGMJVEksfDKkXWPPSEQXgmJJ4S0gt1WWjKXkbSz
03KYaizgxxlojp2/gr57Fi2jhp8xDsn8HTuPjc4t5NORn2fB7v4REmCEfy3s
M5DSp6gS92Hm1pDiP5vv3/ecsV5jrdVt9ob6ni2iKmPe0nPIGhT2HUodR+Jw
lzmWjZMqA1Rc+nHFWss4VRvCjxZC9OoQfLlmwfPhBu2ao9pfa1aFFkgIPCLk
I7Nj6YNJvgv56vhpPvTLVHGjSry8LLLTqiy2FiuDuoPSmngn4RctwfIlJyaa
KZuCDSbeP5dH+b/WPoI4Xjp0hetryTBidJjeKdWvLzu6g2uVzsU5utw9ijqf
o1It2b7RU+dYPRFTHNiF7I4vU1/5NWdvheNptWYu6aej8C0O7XW4Q5SCinDb
1c7hd8a0UiB/o1DfZQzJWLA5EAFO2MqgUAzIUrdbhOh9mSl983wx7IHpt19T
AafrbyysAjKnnSg3NS7YC7sj+laX7j7Og2jLwaGlCDrPzTTyHWKhuTNDNBEH
ziz01PSdT1d38rOfvAjC0snKmHtIDUNsY/FJ2tB1NBoXza1iEAJsaUaEv0rw
TME5i1z3JppK8Vq6QJWkHIn9TknYqCAOaPssHt+GsnSbPKJEZGgqDL8YfPwv
Q2qg0JlRI0KOvhIGHS1A40rydTgWuxjUylNoYkD8XtaT9aGUqqPDhX1WOVhy
tAl+CNGtCwfyNA8W1Lc/jbBt69FTxCe5kBS8rXzFj+F7/GikfqxDwTA2trU2
1pr3NSrvlgHtXMSMXUs6RU9gUf9gP3ycur7YeC+McaGzvEfDw27CLtdMU4ek
n/0Q6KVBUHe6uMiOKEgsaOMgYn7kB0GWdNm5LPHeYOZCeGEf2Zmwa24k0uZX
JZ9pWlH1iqx2I/Ka1RkUIVzGRy7kTR/3+qDpepji/+yyh+w/HSZDV+5ip9I7
snPQrVpJkeUlfJfqoEt4p/V3qAxtt2OhfQka3bflmT8zwaaMJt5hcP7UuaRj
4oIImbZuNP0aRyZaHlm10+mw7fesvxL3Ytq1YKSTWVCnWN7FPmOvvv0iQCw7
nMBqvIp6PTJCP0H1yXMiug4mPom1NqEvCh6J6An44Bmk0LQVtphxOOvm/3oi
3mFrKFNk6dIKXSTCZ9IrebCAVwps2H6XmlAYjLs+MVJ5OFVZqxsLREdRaawb
tZy1Fj+P8xSVsWkuyfajLJd6h4MIgu/lGjD4FzxQ0Sz1x2JgH7LQ1zEE4OU+
sdpgZ3TBHCdF5SHx1AbwDrHzQIGWduAHvsaBcEME+M52Lw5n3S0/m0Bg4lgw
UUpuNOIRcBvRRPeJ8d24uMAJI+G+OUiC6BRCX17R2PE0lsQk4VbPdKnt7TIT
206WFIdH+yG9sb9Q8/awj0nplFrAcCSe8f7Mih2HTRhZI3dHaKA03MS6OLS7
q5aiXdNh9yZ7nlJMXyn/ClgR619Ky1CY8hAuG/vO8ehkB5pE0agaYcu+9z0K
9z4LjY+a9n2+u0/ECjM+RMnlrMNO1weQXzPvlA63nNLLo4hGneoTEFqNS15E
cAzPyUpOn8JA4FDe8sJIG3lKUZZEpCQvDximSi9rBZv6Oz9GSXUgyVOGg1WK
s3h64VKK7kJvaLJDPByVY4M7j4L/8aADb6oxZPsWI+2hXx1TKSFz42J3kEP+
NUNX/HjSRNL6lF0wOdyXv6fxcZCoyaHXxOy2Niu/aM+8UtnCiGwJ8dErqgZ/
+zM4LgdIRWBh+3PumPmCgZESCxFH4lE45J58f5YKa4vwGyt3roojqnB9bQda
Wsa2KdDKqreqW5/ZBxVZudQlNg9ScAQpT71VmGBk/bF3omIRzlta9d6W+UCW
zaeusNgMVKCmbvRksLrqOqb/qyLlfGRuVrbWouDMxMN+Hb7e56rksshAVNqs
UT04XPmWKd0ehFCm6duRu/VEfGl1RF5CHida8IhKSNJa/cHB6/aQ2YSVsw8I
96mSDYhWQcK1l7gC5IM/fat93qZ6qoIpjnRcLWebff7xG87i4FzSTFRs5Zo6
5VXccOgpwla9jYRugTSFT0frDQHWh1eZ4+tQiRKpL/dAN9T++/Beg/1IUqdQ
T92BJdJq9KuEnrvV4vzjQaX/fQZ5NZQ8fB7cB4hABdP/ol/pzIun0Q8QEXej
qWZnmMshBoX8BCPlsi0MxTe/s5FM/72GqAqvfjeJJWw2JOt+sisTrBDRC9jx
6geu9NmCG92V0ih5mSP37ERZfbv7IykInbOyRsJI/zoFoy+F1Uj/Z/xBvrtH
9u/Id4yEJr7G6As4b0+ZN5WFzCNgzwFwhMCuuVVBXs5B7R9vTdX1vnzSqHc4
C2UPWqMwpY4WHoeAytDa9eGM4n+RqDnz6yMoN2P3org61/Jxq6PiRLiHnMSn
3lkxDTvdlQiHdG1Y1DCab/sv8d66pkKFCKLYrv4KR9MPP19VvnqB2L+Ea7iU
wnl70vKrL2JqxNGG61Cw2LUz/zblm0Z0VE4YJ64WP6gLPHyQuq0iIZB3WhOy
g+W6M/5pHrLHy1mzQU1baFHUi8UDaAOK6WeYSUqOvsVvh2T/ox6GkRGVWeNP
+iSjjNQu83rwLYZxTjAGOkRwdYwvHwOLnep2Jcb8gazNlCofPyWdSrm2Elr5
7OIz9VQlJ8PgaRxXhiG2hSkIcu6v/JQc5srYCh0d0TFhOXcS7gAxvrs5vuSd
B3mlF4xQ1jIi0iuNnoDx9enePrzUNGuPlyTokeOzO3trky65fLewJ45kkngG
7ul/oVicYUpbC+8QiafIXf1Rdc/ye9dV5oJYuV/WTjGOoBxtPCB91sRds2MB
YqPi7TPEdTD4LpYSafswNAPKRaShkxszgMysO29yOZkcdTylVG9o5GoKvjtZ
MpBlJrM1datVTaqXopzWvjf3W2WAZjkLcDjv4JbtxYWZJ3csy9WqFB4ggdWG
cWApHuH/fC9jb1i6qG6YsbxDnx1zeBUQJauzYreq4SZV9Dcrila4S47z+aB2
9EVUW9ncRvj1nCfUNWCfqLCjCJk/7zI8ctpB1C3M0rlwcg1NcontyAd3kXVF
QNFme+ETxj7AoaOcNluk671cezNs8obaONcqoGBWBUUCgSGBhEN0bU3DxU+0
3/FrWL5/V1L9i4dKsL/M5Nwy0JKWmLJUjv91DnK0XlQCKAV4fHLXulPraa3A
76ihhYTjSgMGBn2+Fb4Dp6say9XzA3fOj2lUignDpAgfjiItDqbElKu+Miol
+sma2BsbLIjWtZ6VklL8tILxaZbarniMAhqPSKFXyAowbuZ+rbYvFv7Brd/T
S69DeXm4b/MP05S6M0za6RdWoHlFMpd6fIaIHfXO8eosvYRr0lgoILx8mwOB
HXBoukBeluQLQCB3IwpEQx61m84SFTacmbRhGwHAivq1vGoLrtV0mVD/mQ15
8AvK0WdiMa2Z3JARvdz2OPtx8YlKYViPMK9px1yuv7t4KR2PzUVlI1qyhKv+
zYFf1nBhVLZzXKwIPZQdTOYDC8385NYpM36g/fssrBlZMlxoz+jZnPjfLZt6
8C87CF6teufX74HZixOYKrmFJ+dQHw2VIwsCpFlqWmZbaAWOFMp5HB1R4Cq5
/jjqE+IYpanZIjshEmEZfYcKSqfX9O7b/FAY8mtv0gr9pSXXCNbBQdJ1O1vp
QFXtXOhpgRFTWppnnLm9Ps6Zxob41wEiMQblqIR6kGwkdtIDsowghcgpMA3I
2yLiwNnGY0UMLpYpNa3gic7Zp5HaxlETaOPn3jHmKrfiGxbUPY5ZjmyF2dI/
Cg0ixZLjbyAjNxwxQgCt18n3q6nWaoxZOdQS2EHIKiv53XsyaIoHAsNE12om
ALIsU1H8wmwDlrJGSKLw0LzsA1zqMmUC4LYgwN6BCIrnEcLTerbSo+3HcoD9
TM4ZiDjDlHdhSpRVR7x/kS4wh24pfGBc2QmXflwx+6D3CPohbEQAX/lZqEBp
0mwejSpUQWkOFtNPechItKVlPdDp9q1PgQYF6IFRmQ5GlqIGEGkLN0Dea6Kc
e5rNIAielbQoRIg7qsl7ojh5p7it1JQBIKJRqY3DQXIrtw9CDsut8iMhggFP
LzlVMDjq7DOt86PC4CThywvKXrn8ugTJI4Wdje+c8ZGEqgkVimyNLW6WFmMc
v2R/DHNmWockygvkVHPZ62+NeF8oetLQ4oIsauUZxZsQeuGy/ENv+1LPY7La
m4bOtTdFR+ncGaH1BJDGM0aEsUO5M1gLx8FkVHCYfQj7pkaEtUqXOc8vgV7M
VHIBpjvSe1pb00WcyyOsin5WZZ2TSb0Hp8lhCijf+Wo7h9YYgkZ6T59zDqeW
jRY24n8XjSMOYJmp+uaof1AX+ZGgwDLUXQ20qlXAxZgHF7Ch6iQYyR2w5HvM
w+DYB5Qs5XA8iZ+yf814USoACh+kcBgsqnDtSyr3vawDgAfxbTXiJHB/SXDL
f1DtpTfYphMQ5/B7kFBFeJ/EtUaKpQIFBUZqESJixSrKF1L57KXs4cADAmsI
+uNnAYKXJsEfagG+RjiaqkfyrLDFILWk7LzkrbGt2N6IcGGBmBjFosTccqcH
AnlVNjQTAf9rDj8DJAKji/VSMV4QadUxOeA3+n2Vc33Y9r12FjRJss82AORo
Hix0FrRRlRyA2Wi8kqYsET77hNXbIyjhrI682/uWDCtMGyt0Tyh2bDEUaceB
uYaIXlzfk6JfM81Ngth3lX1C0XapwzvBBy6CGEh3CNupSkw6WnxwB5Io3uhD
UjE5rt6fkOE2WQfy4qmKKFMSI71kNfTeHaU7DTralWlrkyweT66mQQGV3lJE
fzQ10EWDmKeHfFuyABXEWnkadCzcdUfQN2fief+FHXW3VTLuahWupfr+Ua3Z
EVDnM4/qgWz9N4YqnlDrEWojzpg76DA9ea9oFhOb8zP9/c61QP/5QrPMSQ7X
D9kylnhsPXcDCa+ne/lBtJNlMaImuEN2uHN9ZcG7grtFPSsS84p8eTZ3Cwg6
zwjACcC3UKpatdVExBEj9ItuvChIFrXGrvcYNcJx3zuNFbGUZlmz6qMOnoLn
ziYseM8UGqKOh6PuWmX8fL7JLzG5l09N1thdhd28KdKlDWhKU5/zHSngwDf9
IEAiuCqh/vPlp0wO9Frk9Qf2FXhu7/g8+rynu/5BoPiplXqQ+ai3nBEEJkCu
h65BWWL9KZMwuPimBrNZvnPESrxR2N6Ar+Cwm8ir/UUfC/x7X5bXF17xjCPt
pqkrpzOPjK3HLV9abt6iwDiZuk9R2N49WYTwyaE5f1ASjXP037XJ2pqI/SpQ
Z7bGAzUQe0sXG9k99icCcxVl1F3KxNwQTTj23du3gIF5TLtKy4QjLxmBWtje
BK0xWmGjsh/+Z4oKdYbnUoXdATo7LMR3/Vb9emwAhxOo1q+Pl3mH4nGgSVnz
ZYvk1o3b4CFL3H1bO+2SVPLWC9qk805Tl4+KiGjp/xlDoLMIB5a9Nnxqqn4o
PEikT1BtwSKKv2tYsrG3Q+5N21+FqOaMGs/EKeOxeMtAvAjsxJdI5UHjILHS
VOxoPm7AiLmQgajyx5/WqMIpmflToyjcp6njnWK9zFoL6GwLma8YcUN1tCtg
jrq5Ak9KFErLdQ6gB7yTXirXVYVwNqu9HHtoVGjWN4zoCb6UzeDaHnoptX3w
znNEEKNtR/7EOT7+2bs636+pUtzxucw0ZKx2wuGXpNwxfkuZn6+5R92QlbRN
7BLwv7jzwoJpLj+z9thmdqRkjqXtBdxz9kNq3fXZcSZ/3rovnSe78Hv9RXlR
d8g5a7cwNYf6i5e+/YAeYi3vsI5yG5ExUEA40Fqpx69mmysekzyxSeL6BtSR
3uoYJbDkD9NzwEOmdW8XF9SH+10LSeN5DmU3LYZgCcqN6coANE+BVncDMU3v
61ff/utFTEWWcpPzBoo8UzSbENm0E4047B52Pv469MwWgNlS4rsoa3p7mGp9
oXDcBu5EIe0oOxoJ5rQ7bCZpfiw3ljy4xiGP1x/1kRSRazGQwdWdTMgDbpAS
MtLmuzonKYGnAtSGP5lpOK+Ecmh8Gogi7PX2+dn65QoE3gRA9YKre0Bz1UGr
j34A7MJXrTc1ehFam+ZgqmOfNS7Ezzk0ggDM33gsnZkQdf2hIt+fC/W5uC9J
gKh6CtV6IISFl9rAG8wMnZmackiV6oouzV4Ocxu1FhL97vNN+LgldUxn8xD/
cx+DE8Cuok3/ZLQysAfgENs2SvU3ttYcMsiVdSWIt1f+BmquobfesdLyMZiI
IWzR7Edok43W5rvKB3K4JeCyBwcD/hlQXUkD4N5+m8c+3OWHZ89QKfp2gpHr
0lkKOyk2FeIjEozuY3wIPhWJF1u1QwP7gSLl03R2YHyJRrsP9keyopO8FaZd
kLor0m8gTzwolDmBomtxY3OrV0kAQsN85fQEH4BLr5A8KzCDU6pl1FmzM4N0
Bn8bmGxvWE2O017b6xvdwcKUQqNg++xURTe3mVjfp9yPkUMQJolHkR96d6C2
BfMdgoDYdrRkxOKrqJBGHCBh1iUX6QfXqzsTLJ3jwD8/AZtpx/U0ljdmZtTh
HutuHjjtSOyhuh0pOQi2NP6yPgo6jcwlZ0aSOdEd0YeTKBTNdvb1pXbc8yK0
LPYY8SWpFatT0tZ/Eyt7rWjtVa2/Z/5R1CwFU7LMvwqx2Mnf/X02+avQfBRq
2/WRD0MjzXo+GJqKY7mlP8FpUEwg4xEa8qK7KcbrtZu1SfdjfmLMfmh7OFJN
flz8fLTYGywjua4I1e0g1aJKH56gVg1vjWMY/t9jl2GXi3ffcfwH/wqbrfo7
Ggp/oujrNso343qpUUAmhX1G+Tfus0jLT0ra7ruhL3YEeJD6gfUimV9s6qt1
RoxS1XMK1dW408hAkidvPj2Rvim8WlZSNxfsZD9SxGNvZB4zasKOwGpcZnRG
erlnZ7t1ALrXNBoJY/ccpyI9dqPT9n+4cP3ULavmjPqDASN9U8gU4Orb4bkW
Xdv5XcrJJppeph3y5J01FXrQNS+E2RktV61/JaKG2taDrxaUYbUAz5+kqkuo
FPrUm7zCeWQPVZVBIXWoTOmIjlt6fYq8jR8Xpj6fcaQrcua4oZe3RDz6mRYN
oA72FCfafxrfXWnetK6gL42wsbQXc7v4nN6jg/jr9fItbdbVbWo69Un+EmEl
DEu5cDzamZBpD+0DETFl1ZaBQuz4GbTM/JZEECJXbbY3wc2VaI9+LvmAQCPU
59yeSBTSFeuPW5jVLpCgD3DZMgq9aXSPXaYHVzKbXNEUq9Nuqvx83zE2JvyV
Nrkq0SA5KCdT9Q8pZtLUv8p0EC0WTBwgnec60UyWfIUtw+9F37Ty21dY3YCm
f2WRn1WYTkAo2z0kzvIt5g1GQOP6mowVEmqh/BOTdk7waB2lCpqZ+FmQb2V6
bJ/whmlC99iHASHtj9l0mxCXOO2aKUZnLpPb+JBIBeDiMJ/Z/WHjMkuWzZhY
jj9e9hOSuZOXlmjS91r4Z0MJFhbfcYF02Qd5wUPSavaQszsysqmhrkV+SqoL
6uOxrXpaXMO+hipn+wqaaCRrwkAwCkdiqbzZcr6TU0/YzTaAcQf555w2qQsw
R96culi0A456G/pjJ55WGpDiu9wgPiiiPEBmmMLlHnEQUJ5g9ivjsP3WZK6+
kOMsQJqgWdAAk/FKzBC9xVMz/msYMOSALm7XhcGHb0LZ1QTt3l4/CTL7Ctt3
tYEjC3avJw0D2fqGK5JaHaBl4p4H6yM68NoLjxg1JUiZW+YLKjLOXtwSeenr
6ZH5GMTAPRg/saXbwA3ZpIb/Wb4O5TjUpUs1ZyNBeo/200D7L5wA3TVyNEms
03HJSPrsqMo96jfDzPupG8xNgsfHFvZS5kFnpgvZJIXXVE0A3ECA3fzvmnr2
fJqXWWkRg/LxVmWgM2XyND96S2+B1D5YQ2jSVtAfh2VDs3zo/UAdl7Xppnar
RJzyrg12QKxYNU4jVP+FZ6YTyeNxI7VSdCROrTtnfmSGPv258kl22ZCT+LfT
90Xa/NnpcO3/fRpHyB0OB49R/xnWC6d5+LVvDyu0PoXbMhkvimeEb72S3l+i
IIy6H5DobELv9SrCZllWZvsUQGCOTxiAweigT6WmbQYFiF4tnkqVNagRGmxJ
TqVJ6ZtXUjuwK2J4nXSqAO5DouJcM0FXsk/RKqUQe5hIUs5Qxx3I70L3eSrm
p+a+UebkRY/tZA6AXQbyZZdStuk18/zt7pDbec5dLUJyytmemJ8EbMyhABci
fPg/adW9xdkB3WNtzCmbx7TXRAdwdCGcAnlK8I0teiHY5p66PqbHnkZiZwIT
Np0M3h7eWInTzbzkp7xV0ICVuDsoWjhNy3T0oB7yNWwGYfNEIbZFMayNo80I
UC01zBMcCdzrHjB8LJjj78+UJ4yy01lN5XxY+yVEm9A6oxAnAO77MlHpKrhc
yxQCdp7UhotOhfx0K4P6+ZZXanTAq5LOK4J39qNAgkNEu+DrY/Xk0jv4z4DG
e/723c5v9JVU0fZc9liyjAifYJJRqC+LFl/PSyyxJDSZYQsFm3ed6/TQ00Qq
g7WzU0RLbVeqECxZAzaI/r6XMSsJJz6PVXoOTtIxSdmNmJnfFLJKx7v4vF0D
lrIr61UfWf/59bPkMHMOobBNOoT8Zp/4l+V8D/Ana5SPvVWHrmqx66bSC7tY
GKbAs4JBlCjJb+N7IGRUep6ZSI4xxeKNuEGZppwEzNOEoWlZFuNw5ZPkcJXh
aRExC4FIiYVUiRFuGkfmxnXzbgYBEbipIHjQXiuV/dBWIyUXN3q06NhgkTWI
6aaiyQg9+P+ug+H2FrrwmuNbCxKyLLwJHV2UeU4TQcYSXIYEM+wsONHo7/CY
X9spXh9K2T6/eFEKQABQY/P7HScChCmai+2yNqI8KaQ9HJqTokn2HvnpaTMM
vd9xUz2tMeko94otzAdmCl/YMeX/vg72yO7dhAaIYAAWAz+WDhhsFgsAG8te
XUOYHwG4qwwA1aCnLXZjV0hwfAkcPE0iDaVfVCMr95dNhQ8WEUK1QB+k8fDZ
gNGza3Eq6dZRbyRcsopJ+mUkUmv3znxNl1itb74i1mRbchoZs/idEozZh/wI
J1c6Ku70iys6HIeVGS8xgXBoL3Jt8LNLFiQXdDdNE+OU99KvsU4bPuYgnCyj
zJRoq+iDxirOnXnrTWXqjD8YSwOjOdu7B+/y9FqgDono2VZ3dp/8CLSZR/BT
ARBGvWb9cGh3X0j955EDlOYfCp+6+uR/XEEmyoVV6uM9ybdQfQkIycXRFMcK
jTGnCQ2A7+a0FTEc/M1HDmK5y9r81vphPG4tGXwtPQNrxBdYP9PvTXJhjXTp
jiPh2HulJrSD1weTdAjjkhad4ojD6O74gfulS3pW+OmCMfMOkZbMjQlNFAy3
HzTUtMUyiqFFVl5I/pG4/xc9juDdZYcyciTWs+iRRNKm65k4gGAd0Jk9Fd1W
gpT2o42t+Gaj7JUfS8FqOdq5gpJlyLCoesNVlklW/TTfGSymqrDKi4gvIhNW
VRYmSUXobFL+tW2f4Lj/Q2/tgaur48gdH6/NyZRpO9/MeExmRPIXiEw8auv/
tcTA/nxf3NERtWr/aXnsZoXqKI3J5yb/Rn1Yw91KfBL0Xv3s0kq8I2TzCCP1
2t5f2oqBK8kiHCNVSLakv88/hWKb+IutQZB/iCx0p1ziF97lwhdazjBrxBnE
KjB90GIrZAGpDYuTMggCXdFgHDwRz6VS5un0dL+zpa5G3ZdpW3+OmrFhqGsN
3I8h9qWeBgoBDP1zpon2aQwz1ZNZgadJ7SX9BHhQoB4mGp0RTNrZ8oQFlsU+
07JCla1p/KAOdlOKPWCk4bg0VQXAuSfwqUSItRczZLjjmA8QdqpRZfPR9n0V
1y6FxFrfy8ka1qv/Tp9+XYoM7Vjm+Tr3rumwAjOoWTwLpaBzCWIcBVp37Thu
INhCqV0fVuShvh/xu9EV3CWEKkjwOqHPy+I+3OVo++OeLmUnwn5SvkwQxvaM
5jhAiJRNAq5bb9l3mz0Ld9P4NR42SFuZ39h3lFCjnORPRDizrOFK9QMuTa9v
OdiIdUxxVmfBjcmC1CfSp0OaZDVKvIz2GoG8z+1oaWAhohrVyCLZctwu6wAi
s6Ia+WdF/V8480zGfnVorW65sw7jy7YltPzC58sdi3DDw2fRC6Y94I4Nlo93
yksClHq/PAchVyQ4t6V3GoNM3CiaDmtqWdJytGUv62fysBXdCVUF4ooCGJRa
16Wr9jyEfDTTlJ4ltxIFaawakG1Ui86bMm2E77smX2/Vk1dqYMwr2BXGYw6b
yxLdxy7T5NNegORGcCc3blx1LOUfYr82zWH0MTXySRh5hXF6vreN3ZDzmtlr
6QLgH2rWgfFWettLNLrNa3+1q/UoCgoQIJDmOGcSEjpQW/xuY9/ngue5vVAM
2RvncTMmCqHmhZcULl28rnykuugsrbEW7+bq0Ev9sdH6eerUxNd/E08ocXfs
VMTitjjvYQmQ8pxn6Cb08gzdBMt2yAY3qopn60PKt9JQ1klhds12biohBZEq
rP5KfnP8O34OWTd98FRYFhHery3Gd8ytguF/MoOAcQy/skS+rNVJtYbRcK7n
lU2gPWyHMyqURL6xbLMofhOLOC52sJHRqBBtE1sj3J2yMWCj90EkdBQMeSu2
cWCB2OhKy4tgekWA7EJtzGj+cF35G/mFGZn9te4/p5+j4up8e+zvI+H4UFOu
LL1TkLDW7I/7ElpEiWhVEWTYRNg9OovAZFDxGk3G8ftjxhTl7LKQyhP1mBC8
nXIAwAm4589EVU3TqKnji20E7bq2MvV76kQaRsZz4AprN3ZiTRV25ASv8w/U
YwbQHEGZ3fvqrfu4mHcSpjnvxHoBe+l4XyVkUVijIkGe5p4SKehwjmh5Y7pV
EWKcZvzqPrcGN0DkeeICCl4773CAK1yxH4ppFt7VGtqdpGRl9Hht+8xuYuQM
0QheTSTDU/pTNMxwoEiySTuveTWMRNPaWfPXbqIAF3fPZxLLgkMTxT366rxP
qgktomrcHOuI5cQtAVF8ohri1/FfTNP41hI7ZMdSRDIPQgS0+7RWS+PakRoQ
FNEN2XVJNsG0AOHno2ixxFwZkVYYJffg3sxkW2ixRGlMUnDq2KoxQOSVj3ln
5ysUeGp5WcT6pG9z0FX4Pgl5uV6vGqWTsd0lc0ecOPrLCWa00L8pUu/O5FsR
eHky8miw8P4qapKlw4O66Vo3/A9b02tOwBLVYPRmJZ9LVbaKSGtt1lxdd3rZ
ZSP7gLRM1yqiZ0lxQY13HsfboufuAlFbE6Ixvp5WLiGqiTeJYrPK/YSotI1w
kFmYM9nK0i/iNcCjCOfajQg20QYPbAXU5ZnVt/N2TDECu2FCBmA7MbxL9QuU
x88Ldh16vp2cLAkSx3x9jiODn8e6d6C1xLZpFp9R9jLXQ72Ir8mvDsN/5Ijp
9TMfsW0yZ2hotM3yt1KldVy5Dj0SNI8bkWnc7BD7NXTm4OdiEaHQ9pjzs9ZH
S4rPtygUYwH3CuX2UfHfUlME0s9lqpF/K3QXDL386U+1a8i1HA/eoqDZM9rl
qSzKY9GqQaPCvXZvuBrYpg4omSlMcewzsEw9p2CA4nQ5BCUsffXw/Loc5orU
my1SfUGUt5D9fwSysxclJrDN8GgUoAGeYhT1wEWlYmTiQoBQyGsU6h3QeVS5
7GmC6Fk/Gb+JlVNjf8weAK6nQZI1A8dq+wpxJH/eoxlRciJwdBgd2gv3lwmr
IF8YSCrotIh3jsDqX1a06BPxkvIoRgcFBuDdrbRZmfPJmjGIM8bhG7BbxP5G
ajw15TkKPMFfh6sLlLNIx1MnbuasCosTabRp4/4hwWGlj8QrZlRdasnKbUZm
+t3dH9E+NWT8LnRSpLr5OSN63OsTyidSPfHUJt8qtqLlVprD7qMvE76SOCOa
zWxlN13xu8d8wwVClcxFWd3xKhiNwqlSJVFHgpT+Qxvwy22m7Vy57bL7uvr7
TFWdKCBryVkcIpgUthvCYPnH0XtJp9SLB2IdNsnc6s4GuAgf03DK8SZ50Tan
twq2Zgua+SWxHLF2oPDGYP29RzH8lOH0X1NcEGNxha9tMZTdFzL2/Zkpa4uu
3ozqTGyU3+59AsDgjP9QYesq0MEasovYKidA6aYlSUg6VosNv4+b36/EdhG4
H1lfAFSM2DRsxb0IrGNW1q8557H3PhmItxy/xxcXxKJgCyy0OX4+jk665k26
yoYTQNsURlr47VGzrbYK9PjGzhlh4uL2hvq9llXdZ71hGSGnPNNEmCBa1FDu
qg7uw2bA3fcI6spoKzPyWhjuRXQVkuRXyFr7IdVLUoNkVvd+FF7KU/e3cMPi
DozWpmdB7zImFt0Ung6HNLB7AX4x0m5uRhyKEu4wwd5yQjPuaoBBBVRj9y4U
oMWVVVPMMQEITHoLUukloCdIjhUlLeURfviNY7GqNU7X4GzkaYJfyz2wL85V
hslYHpDa0p9yCGQPlqSuMt66/iYocpNMpzdUnVaVKUaopuoYSps0t06u5Av8
KRI3k7qC4qOtFK+apQrY0p1o9vLGs693JrowyiTNlJdA0Rfjf+dLeAJ1f8NZ
YkSQ4kQsrvw9K8RV3AJhnsjUXWINlUaVpNnAAJ7p1/UqCRVhPv5zk9+f1cDy
ON66pvd5/22qTnvNbzG7UsthTIBf5vVPCAdmSYQx6FEAVQp4+RyMzr3YThBt
UtWM3geLBJzfBDoZ8Oafx56WqCbHxvUuCQ4i2JpOZU6Xj2yaxzGE8DI+4py3
iw1hc2WKIApuWpW2vjAHGUesAUi9kqEf1hgV6Pa01G6eDLz5KS7cbDZ89fCS
d13kbfctXKQsw51Dd6gjR2NSQ0xX9zkx596OrStYeTIXFQ/ufl9E9dU5HYin
fyNSNFWAHPsb5oJk4AXXOmK12b9XI572+rh/Qap4bl0I/pH48/fs8XCqk729
1jD30dxSURkYNArnxx1NHxXDRjgquLXzfmWOc+495s4WP722KLzaJrizc8Ji
5tRe2vODXZe1AfMIOgaGCmUZLBkbFmK2BVXL5u99rTopOr1MDzngi/VTKgky
zn0BH6/3YOJlrWFLtg7w3BGdBVuRZYudXs6p9tbIkrbeq0pOXMCNu0z1eh1h
4n5a0n4lkfnqA3bInMJY7n47OImd5XU9ARgG2z7MbYTwqLt31GBUn6XLLoFd
H3J/2cVRZEtmEzIM9QXrxQdqJBw8J2GA80pa649X3rrPABgxEITVQysO2EYf
J31WEnJPedBS77RX6dMoVgnVr4F21cAwEznzd6uRMrcVGU68uCsmGCcEWBkJ
h6doxctJY/NKZHyU4aWsPsagKxVluF7zeWio045gNNJTd3KczoqAW5Pt14Bw
okWQ1ftg+coo8ZaK1CbyrYe9G+WaFCNXDyM6AlJ2QBWYvlv7cvkCETbym1gb
dpdXhna2tzAxRiBTh8FImlWVyT/9De0quq6UEWoMj/Y2JWSwDo42fhPL4axi
hOZEJPWbJD63vxxw9B/lX6CoLtCRSYxc+fSrUOJeKYZx545h1ZIWmFDf5iEL
FJnrlmpV2hjeNJYQWqC6kWwC46vtX3ZcLRS46o637zAMQeKwyannnVTU3cvf
FEkMgX1tELY4CHKgyzCh3lnaoeSkOTAjQyQMR8mYd2wiXTUgo4GJKzyTIhut
SFG9T5f/fzX2HRhrbI8kd7SwB86Xw5zS/WS9T7t/S70LSS56do0bz8Be9Tb8
sNmtswj2aCbKZH7HQ3Do2YaEWis7OodCbysv1eQeaIluBDupR48DvB+Wndg2
zHo47qBrj2hpHgCRWxOmCNCkKe/z0kv0O+Uiua7CovPqsO2I6QDtn5Cy+8qi
JSRBlE+aqlvHi+FRbpDpxQaMlRTSuEKwLnHpJkuh1ROK2uYPHPN6GoogGo8k
tnekUKwtQHMn/HCMF6MnSeSc6x09QDRSniZSt2UDVsk+w2EZEYloMv73Jlwl
Id3r7B99sWHGQ/fYfspMtuOkT5GdL8HpzsMRWPVMblaDQwC/9fq3RuT7uBv9
oym4CZGGrU4QeeyI5MmSXsJZQfmfQZpH5KspMOLK9OWBLacLkDW7tgYHtWsk
/WOamQ9gfHY6afVhsSyl0OxewOiD+vf0cwsWnhbk8Ee/S+MRp/m/8cR3ERgS
hPtD8Kb1jzFsxoPSoPnVrzTjrV78OHEto8hVZaMxc/DvAx9NYaraa9SpewZ1
jmDa+lRH2iZZRLW8XIenczLOJAsNIBL8b1oygbdT7jI3PaBg5nQwSA+DDqC9
81m+pe2dVqCPcg+YU0dnBJFsAnz1picADsqtqMM2TmlIg4bNguzx+zxHezwV
fI+Ugf6/QlJ45RdrNPAxlWguEwZzYUt4ceZHrujG7XQMws4abBDqYFiBopjY
HVYhZeeXTc6YnwBZQrgW8/V/U/OHIoSuG0+5ccbmNUS8BWmVVjFGWeO/vQ4M
7atrwdHO32mi4iYOw44zUlDWd1uLAPvdt1sIbbXI1uWfL9NY5m2dqE2CJbDg
UOPgmDeo7Oe/PfQ+PpA594gVYosWBjyxGwamDqDmTopAUqjpFJcMmWeS/oMB
+mdqZP+5HnkfyfIGSHVlw4qvlrxd3DM/b5RX7BHIwjw5IjTAxk3hfkb+L7Bx
qnv6e7nB6Guq3Gc6m8yTiYAXh7T1KWDADHS9bXWIRpJoLu+lSrhS/ST9x/hd
R/13abItNDaiQmPEbVnH6f7I+0wkf8FA4VYBZm05jRvN/T+28Q8ysLCE/TDY
j6gXSBzr/ffmJfYjCVAmTC5QvF4GhQEkcc+SH99YCyhtitnYAyuDXPFOQGCf
++JmNkNWU6jIKYsRcdUgY+Oou8VAYNIRnAa5nH2qYN95Qu3F2ccKDZ5QMqFs
IHHqriw95Dysu9bzP4uYTc1ZJx2u3foiTcNgJUwFvJEoOBbqAe57XA8ud8hh
IH2rgqYOWMFGqSvmlGEvZoSc41ptA3pNuSfb1LltDYiY8iMtnsU/+SkO1kYx
ZjWr5mcHSUeATjD/5VUjpz95cTO6JnmRWe/ywLrySO+muJMjiYV86Hp66HMa
0rpeearDEDkECz3kDrmjfZz/H1aetRPryKqjniFIfXKFP7vrE5IqFB+ZaoS5
1eQ/FlP8mtoK3OT1LLhk8NoyG1MLspK6Hmccku+drNC35XLZwHc5BTGi7cB3
udFtIwLmS5J7T9dnLAi9y6S3ASt/R6ab8NFzR+Nz7G+xQ35BHIDQ9v8sUVTU
3BCrTTyddNeRJyJiYpOOtIkb6/ujRNL9kqygK41Fky+KMLUqLhKCQfnl6wmP
pFhucAdZpILx1ZaIxR2MWLskv/eQSoLT4krVUrU7ZfArNGVmh0lBw9m5iZec
r1AysQPjBb6a1SNQ+eofEpm1kNcWw3hQp42WWrGBrqPG6K5xQaX5uSFVsdjt
36Yd2KJj8sAOlVNo19Qp9e+4P4KoLY8aCpznUY8Lsz52FkWHTHVBPYIbFR2D
BUDRFehBSFRxyJdrTQpWt9mB/QrlSb5FKX9oawYnzaofIV8zeacgL/m34uVs
Ayxy9cDNTRA3jb63xYO2zLHiNM6u+j1U9gj3tHDLeYOckhgnwBblIOarkcuQ
etXVAtT6VOxrExTDRZtSdtzHOf5ioGuKLLZabUUulUoDfPDDSe5CMlti7nnK
9hAbHAHSMehx5j8wON3JVqemaBycV14QFkhr+bAEAm6/nQGo+n7R+EwooQsR
ZG/OvxoORtH/6EiPl2rthRZyOcRWifUnIuSqa80wRQqBTkR/m6RCzpaU8RCv
eFn4ytx+vW4Knf6TBnExC/8yOI1kPk9FPwkVdqBTsA/ArbRvAuIkOx8+6Wxe
SfoOFQTTOt8FKy2kLrNU06GuER5/3NCGUXFOVIVRTMQP/0x2eCPALq32+o3X
Fh4Rv7mysrAMM6vXiFieEaQAvIAtFAbpOxvOPalCjhDp4itsYORvm2+qli0M
qKWlmuAq7Rq5txewQdBL/Dv6iPm0zeojZVJ4vq4TIxAPxJnaMyXM/l+bzP7s
CK6+2eb3huRkeGloKCTnDx/GYfjoUK+TFGNXFAbf+6gSLaZ1+uGikuMjqItS
tNgVUhVSXn45VukfjXxj+a4uKOY0DX25npqo8UC7lawHMm6rHzZDYHkQqm78
J19Kbdx33C4Y1yGB0sbxYIaQQ/3Gh3uViuEjKMWhb7ZFryjvS+nD0IAYTFcN
5cOxgG7OS16Jsh1Iulxppq6PjwZrhzIbUJHebrDW8QLHi+eF4NCzJf2No/E2
3BNJhqfkQQJ+keeH/7JoMoq6Bvq1x4wQFAlb+Nmecz96wRWuhjUbIaddSNs2
nI5dSDhcZ8jpnZOicY+QN/rR2Rxa/NER+oqf63UzeK+Z2nLwKyW6lEgQUXWm
A/GHcNUuc1i54QYidWGGurAEvaCQ3PXpRXjDmncsDa2Cdp3RqMY9+vv9c9bs
cFUJ1QEzFwG2wim3ntuC3lLVn5TuwdNO8FoFteZYFkIRF+0+aStINxS3Tyxh
ppIBawa45McErr59/76a/YkPH8GYPGDptBHmBqX+y52UjvqjSnUtPPylEq4b
FqjVZYSSuXg29ktOqua3djgIWGaNqSXUleqXVJ2krOFSEvnQ24OLcYZROY5p
Qu+j+U07HF3szWtonzWP9VbPFy5HIBjMnEWzMYVnCr/y52OmvckaYDrt9V6N
fSgeppnuk1IA0o0dK0rv61zJVfAAyr0D8hVp3Dc1Mu3gAQyWOAJZu4fvmGVe
zNp0ygGisZS1uy34WvqlJWZlpqAeTCYxLw8R0aTFzyGas/f3FyBCb6+qgomT
5BmN86tRtV+dIix+Psp+9yjXAcg6oQ36t2aK0VMANfb4Z9NL6Jn7gjmgbeVI
9rMAD3wP5SO9+7t8+kwnoAN0J8XpT+NiNLrK2S0Akl3jKQKKAeYcHdCCdSMk
EtM3KhwSnacMc1ab5jPIDn0Cm9/wVeH7Xh53HNA/TVfjC1N5r2YaC8HrfQF+
Qvi7ydkUmbXnesFhTMmGClO4bbuolIF+Tvq668odYhyHh6ciOmbVGEPLeHyP
I0W6jYG2EzxhUI6gQ8/NnHRJa2WFfudWdD7OtjjgTd8Kt073f9lBSMDQTTRf
WQMVyQ8QSCYzL+u2tnA16umYPxryCeCKK854hzCZSj6G2U7Z1FUHxy1FLQWk
apxI00aD2xmWi8QsNPCH+4FyeM2Hih08K2aTeYMdlICSP4y/mxz4oJX9XuXX
gU8Vt8UwGkTxvOhIZ02AFHDz/OD6LPDfseA/yVpAuQPLkpc4wF8H3dbMk8N2
5OlLgcZ+VI7FK+aItJfcHVe6YfXUQ4PIOLJzJJvzMHHsac79p+IC98WXvgLg
eK/S3mh3JYlf5Y2brmd/PyN3EJCRz0n27PP4805/uw4B/1LjhASxC1bqw9YP
Px8igLYJnw4I6Gb//ilhOkd5WLYt4t/E6QOHExPEWSArbq/8YsMFQbzbSQLT
rF6n9iuZYIl3t/Rlk8TmO7b1s8pPBOKhYyoxP55N+WwM0ZL5RsJEZEYLTCNK
9aU/TDug6ZBibLD61C2HRdpNxnxbQGc8zN9rylYEATMM80Mmc9fN63fBDluK
5LOtGrlqmHTVBtHLTRYC+SMWIWwN5KZkJOhTQWUKoI+n9XKoaNSjnfcIddeJ
LC3fskg75NXF8Pm/vdOYlhFHOp0fYjC4BmaF+xDR6yM09q7O2+R2Dy3p+/oj
MzXJmdh8v4iZhhSXHxk/hqXQNf4YLCMlrxrefhgG8d3c5Fi+B7LvFEdB9V5p
UPyuczh6dqR0vInYh9A5f7tylX0hpUKt2eytYBjDsv4FIGA2uBNiIeh6oEA4
+SPfDNGFxhHu2aksgEwzanmR9gf4Y6+DNMvx7N6ciOejFHw5WTQefrkxYnSp
0W0l8V9u7NJ2ppkEA8JxykEE5/+NScXb2k4SRVSybNatTIIfSytj+VeF/fsK
NoTox9OlRMy5CM3iaXHW0FGdbqm5xpD53VZCNefo6vyGyVByYvKh4kHmOhtC
Q6InMXnrkGXC0SuvyCWZ636hC5evDUgmrh2pBGyE3rtlcJPHYCU6pa1G+aKg
V91rdz2cPIbZwJox5ofcCx1qNVDTKr8WOWAbLS8zrwvIDpXnTorAQ0Rv1qPP
StkIBO10TXeA2wDlElrMcNBKjHIbyF4JqItCWFcdIby19lrn51oJIf8P56Qp
pb/PEc44Ke6wPCMwBlFckN+ajFHsqgCbGBYLgT8WDCHeYAPGDyjBVtpgqB66
NEi1Ldb/1vp3PnqCq3dzRtjlH13toV6DYFnXbRlGi2XCegFoX9aNvWaOEK51
jZ82fRBUg2/FxTIVcVjguLSwgZaKVBcGmFy81ggIpfrYe04ZO1CFqvMWAWw8
0A5LUKBIuo9+i98Ua/C3X2DxT46xETJpODzKU+yamjj/j9/J9Tr+D0Qkwon8
tTDvK+pD5jGUusJ2fKJqToAS+UGRAUMcETRj3qVLAfIdqFTyEfiWzTv6y/pk
VC/hsWqIl4nu8RMwzEO278Db6NEMuvnofI2z6UDxjy0boGnKh4p5VdI/4cd7
D/GVB+Eo5eJeGffPzQoeQe/9eiwb6JW9ArF1kQpqfO4kV2TCaihzaSoCT9gP
asKNhUhBlfyjXGMfDluevAatRhHerj7//83xhWhQPFH3WZAZYgWlJVQENFiJ
TAjPihG+tlWMLq/VFVJONo8RlE4nQQgHLfL8HGy977YXTGdpUMqdNQHhs5VH
tMrIfsElD56qHYWFDuxhvTaHGcjOg1gpLMeqK5Rcc5NDiSV8dCYIZ5yumXmQ
wa1Bl2jhBzyxdNEo5H09QGfJD/8Vhk3TuvTBbCtcsst2R4eSA4z5ntXaOUUD
TCnFTlloltCrD81dQG6v8Q10+oxd4qhs+utO8csScy9E6MWIk4TdRxH8lDqB
8qje5EtWWuRgedcQhM/Z822NcIkoBVn6DXbqXFGYJm202xfRpNy95RIU1jek
CJbdVcas2x/h6J7KupTpQMjuZvWt0SpT6IRB3s00dDsx8da7OG25gxiDaSy0
G+K8fSIZarT36BJ4x+Bw2n4+ILDn9dRDmypuaf1uxvZub6Q0U6y5lAPqQIAy
5opaCBGcuM5h1ylvlNkUU1RB7LyyvxIM1fMiHsa9Mb48mqZgniXidZ5m3CZ8
4ti1az7cnASyXxP4HZDxPhRGSigWj3s8rNfbLPsTZoaMCX1DJQ7UHI4cNdqt
1NwCut23aWWGl9h1xVHdODIJ5HNbbCS8qgoY0TzaAsDW1c3juXVroDDx8yW2
BdZzosWnC5jeYESirJOkf/jtIQE7MjLmxRy0SGn/yq1JQrFHED0vvZ2VK743
ELhy9F4hFi4BffQz8hBJp6KbegmcRMPxAcWIKaf6gjkOSmFZ3Ox+nzeMldbS
qaDjCWTSpIWAwdWcsGnrw5UM1C6Zkseo4XG2jw7076bqrfLC8fRerUEZLXdD
or7FhVepcBiLwRgHEg3ad8RCYU7Q3dERm4DD0kBqrlfuOSyxcqeVyZMRVHJV
1puyCbMXSDJLw4+m7OeaOwWAzC1Vv4ejO0mOwQOnv1IR0UXWeeRGuuYBMv4L
BByBaUSlmt0D2Edk7KzYeNl/kwavlkngHXL9kDxlKvm+/R4wCOiZYZueQ/tv
fX8Q0B58kbQi2zLgzd8N5MlZDBZxPP8suA2kP1yX9qH3IBWUmv6XQesv083R
Dn730DkID0VTKXvl64Oo5ugWNIWIsuLYdvpRT4Y/j3t6tskRNoFS1lSyenDH
VvGkxRnnXcWanFwEN6Gv3jmBoW654/YmhtAKD7soFnj3atRWeXFcE41E5ERZ
lmHmfJsJypiuhCL4gdIW4v9qwGb8qlXr3XE/PeE3shcD6k9EgwoXOYg6avp3
tL3qt6J4Vs1UrvD0qT0PAt6lwMkAs1xCJf5Pqi7oHpDEWRbNSaJ5Kt/xTB27
LyoSgljxMl0A4sBZL0JETgvgtq4cgRjszv6HDGtSfsOvDStJYRh9GJMLu/cY
hLHhQJaYpHpie63Yo1nwBABgaxsKsg1HdZ8nigm64aw7K/iVP6opq89Egce8
GM6lLdyXjDqjJIMOYlabkNO2CVWaDRu0bdT5TEe+Ls96HT+Dv/q+Ul8BP/dl
DB6YQFG8aopSvY7ElUVup20S/kB4G3M7XHzsyZNy76Cgb6xqM8JfFu7bsbJq
QYwiYkEbgzctQVQXOYXkyx1kfCeuBzBFt6YzjV3s7p+i/gxjTxhgcXcucwkx
/bMiJ2vfxEzYE/7ybDDPIzOKz4xAlUeioB9dEcAP2MVBbwhoOF9BQ1ihIEaQ
jXlpSYyT9rpcHCvSgD7VuLon5WmAcb+C9rRF4q0hkShbykrqM9LwuLiT/0pk
/Hf+K8YceI2r0Lf4rCG2vXiLLQdxmSjZ3nyQxW+V4csEdxnMzq+wTVEtpcHG
9HoDDpiPN22vf264At5+jWTTjYMVRCIj0Tmno6aVUYlMBIhgohVosGbL6yLP
VQ5arw1dyngE7RLfZ6jkDKkHnhaBkTnAmmHk3cVPMT7lUnJl/vE/XzqI8qSy
rGpOJRCSaE+WnCX6IL6wdd4+7UtLUenslOnA0dP6ZB0lHkrBJaC3dgXLCbkk
FBHZNuKQVslOSv/LqHUZhn3ns/MSSsxoB9Mr2Ewvb8ncxg6h8eJvm+a9WUdQ
GobwZhVnWfs2stgCoWAhKLqPJaqKJjfbKCkDaq7FyAdSHhb27X4PMaiFnf45
MSh+iDsazISWaox9u/Dr99LWUtvMzmFUDMJ3Hlq0eq5LlnNUXmKBNJQJnOgu
zBSi8GJAE+MyJuY9a/6ZvIkUEgdK3vdbiZoFwiApSV4lbh6rbcXZM8rfe9xn
ECJkHJ+U2MeyHBsfnNRjOatCuoICSDcJ1/S6c+5PkpNxX8E8MwR3qlg8WCcX
uRp3d6g99euxQYiAyS++uv8FLTCpFpYhjAQlOAMfDT+X6vLQ/rpG/Mf02MnT
051ZtGdCNQ+wC1aVIa70TApJhAcmtL1mMBx31lGbPOwaYqDMoqKebMF4rVTs
bjmMHR1xXD6+0e8pdhi3/dJswWn8ezfNXP9cTJpFvh+Rmdoi9LfrqUoV5Bx2
PIdQPyXN6xbgbfoVbn7vgqwsh+KhPjpDhuRCmippD14L5oc5QNkVIIHOIO6M
5pFcx//jMTK/KlreFbtZqMzV/WciPV3JC3HcZa9slAV9rtq66lomWjaOwqcv
0fp72e6lJRr/MyKF5cP9T864CQvjymSs2BN9Zj3lW6x8OzTRSRmNwW4ZJT9X
xKSVu12x2Ku79tGnW7WzLZdoagy35lgzE8LPKWsmmBKyCCFZW5E2Nd6hayUM
Mouzol04dymWDawoFr7XGvHW1C4rYHkn1D3yDGMObCKHKgzw4K2SJ7RQMUpi
UPG2HbKaOtiRPrubMTFfTinkM4zW3ekuNDfmMQDm+co2BhuKQYJooHNv1ioA
PDp7HaDmZmvaX32T80PEFqxqHckhf4i/ORtKL4zD2RvQajLODVFzKacmiasK
KEsi8LmbIXOHSv+SAcFaMsLd9ymTkVH6518wj/IMdSLn0mXcOw4HiiQjglHx
KyR7kf9F9+Hnog1Y6vtRcbuLTfywKD8ctaiQbA4vo+ANqkXWVrQ8qEshkU2H
kru1TtUvwVvcqg2x6rxU5yhtV711HYqQuEuqJrr4xHn0Q3bBEcpuoogo8tr5
NqZ7nGiT66xS40U9WfC6a1f3cFms5X0HaMhuNeye15HwtqNzTd5cRIJ8ER8y
Hqygk+KjM73+YMxWpG7snZmjCyf8Ozl0yb+daQBEdjkfFlWRXc0n/r3r28FS
SnA7ACO8LZd3kHpdWxxSnv8LYX0RAfk47hdiZ56HDJ7DNp3jf3MDaAAb6m5q
11HitNYJ7thfsNaLFl1Q3rlIvApHXoFzwOcxpMMIv/hupM5kcD39Ni4ZMyUw
Hdz3hFByR1Onqig/QUZgGMGs0wHXnmz9y0fz6HWJHUmpqQTIHL2CINw10HPi
uKhgBS2UD6TMKbOmRRdTTQZRnxn79DPOh4OyZHr11rhre/N0ZD8P2cnUoaly
AbNUg2ncOF4XOnb9S1y4d7Bt+BmY+hqLM7DmL+4B+J6RmwhN0I6Cr9PQKw/L
H7FvJCXPWF5n0NDp4gahs6eh9p7uKT+iIbhySNdnsX5PWXnUtDPYZardAdls
Hikm+UfwCsogCEHSoLMba9rNIFMzfkMPc5KgPiOuBti/b/hpzAH75FvuIfp2
TKZdxV/vl9LyMdt9I2429mFePr8mcXoXRNcbpKIL4U2owaiBH94g/J0m1jIL
UBEF+olB9xOHpg3Gv3/ZG/CxyZKDvgI0lYEvl5zzZqZYlOp0Bgo+kf6T8hWY
/4DjqG9Etj1rE32odkkRfQSzvZOJirEeQuYmTN7oG+N8X61KP+i/oUtdzlV1
BmdITkIT4X3FhQ1/R56Ua4IH57ZrXqDhou8nP4flgLKWwnw6ZHjzSUzdvcSv
trzEOGe5JxaKNb0AGgwKk3afPLfTwr3Bc/GrYYPjuOkz7Z4iWSKhqZBNf4De
WzgGcRRuaAJs8xlt4Vf430/2P1QTyMsc1mcUVDFd9QZJGK6YfXPMavqDSUFi
pBiks0geRed2ch5NOiZNl8TSu3u1crDEj7nuytO/OIdet4VB7j6iL8ZR7YVy
yo1woxUSEHczu9FM4uPGGaCMORx9KXf9dLTSMV0Q56y2WHdUk6KfbVd8Ygrr
cGF3wGOFbJHAlqrH8o/ePXuQpoqKf+VCRlCZv4bpQlV5fsezFhynlr+vK4Ia
M1zhyc0bujQu77frBAGyYrCbzDbGjM/zGjF8Ao29MZmNdEiG2pNi0DGeGsQZ
WUcKt8a/es3AThmG5pE1osG2K1L9bWLV/GEOhG4i9ZcUegf6TUkZrNBlhSha
PWq8yHLCPGFSt+xxeBIXgSvFQcBKvtqvkh9j4L0Y9LYRlf0XekEFNWFA0Yoe
3MrT5xH3NyU9uTZW0EyoCZReFQ2w0m93YuUppF8Je/BI2s4Ju+rJLIiKmtVS
dx5EAwlpDAi7sK5NZJOrhz5O43HT4A5h8Ot+hytU7wHv/k5V6ILU2lYaF2JN
A6TKc8u4paV0WaClM2Nk/gkjx4uVQOE79qIxWVCpIl2frN+4GxJhUlKcTZQU
Ouwllq2xDeQmkQZPbXlnSKWqILER0PmO2eFd7GPicJDZMCtsSEWEYx4fVuDb
SFzYT6gscFdyvZsIfHGFR15gXADWTnjOJ8+pHBvKDFZyFFXC+CM9k58ZLuKF
cDWr/jacACKTFsyV26XNvwJc48+/TeHhjVVFxl4CPtfjaRUtM12s5mPZUm44
yiBPvAbvju8IOVmhvtzZhu2IHl+c5KvwvC8qh0ciZFKR7zsRfk0anjbnmOw2
bv8P9MXdgAUaj4KRpP2glaxnz2HyqxRn9Ay3CcaeZ7NnAm/xfpRBnJdBTMFC
xkkC7GflnvsFt1iwVDeG2o8TQs+ly+dVxP1ZM/4kFgZzYW+Ot8Xw1w0YgbcI
OGSgqLGdOqds9mocTvlBWAVWbcRntC/nBPIdbAP4RzQuQhoTBxNYImZZThOF
Bz6jS/+V5QvHSXrelHygdRsGjlpzaoWZ5ITcburDNdj6GMYnkDnw41zLREFz
s/ZXAbZ8AMzCX3kA/NDKO+q6MJ/fOD6rzrqmQHIm/BfnRzh6xqwJMHrcDV/T
cqBoF60G48+PkJr0RnotHFoFCxHkbPdWCDSc6Ql55sSHvDIBVbDgqVrs91y5
8pG+yM/LXeV6+nagHwD6ZCCDym3PwknoI8nIRZt3VpJ7JGS7QTPPSBuIfLzb
90WpxTJA3NCvSTaMyzb3Gyjro7ACflIvR26AyTm0adqbV0oJRK3D86A/U9c8
C2TIEmrvWJtsmauacJVNKfW8vEqBIByD8PbCpmB4uBkF7kQiBXKMmoF3/NNe
xd9LXe3K6TTYLEoJAARlyfl05TGLUcUikjaiV1h/5094GWarzig21VEuGqNO
nQj487I4th9jM1sHwvoLpMoX0nvm6c/aYUmyzGawInl8avauf+oYx8J58ZCJ
6za5fF6XqUymKV7b7PazvE3u1k9adHasRXkOhk0Er1WWQgNNYY5dbrALr72H
Jdl0jvdCYrmdPs3vxzxWCAibgpLy4UZo8J646AYZo/rh56pa3cQruquze2BM
BGgcv+f3dq39Zd6avmsGwfVJf7yzG+mxfZboQvUVhV8bKgsIdOUBzDxDI7Ni
rPJvVgMkuT8MmJMWOQ+C4mScw2GvyPuAMCuzDRXPLevYKTc0vfslD+R/pwjs
JSdgy0LBGxBRkYsns6SqQxUKe/h+OEKEM75aD77ItO89zBaLoQHeNWYix2Zc
oiPw0EKJTBg9gNvCBhW9oVlgZEahZX9TQGt+1/hDTGA+vIiwO5R5UwP9MrD+
U/H9HWwmZiPxH2BY6a+sFCflRgK8Oe8Y7grnjKyLG+ubAzXDVaenvw33ntmo
BUfKBCNW4q8cxM4JglGivS/x+2ytpfPz7H2b8WcqqPGhnf7IAljkJTlJ/QGY
3VwD+0TBuU86Zx9vZL39BivC6yFsS/T1O3uoY7ZxODK3dlLPpV/g0RXeKkTz
VKYR3MITVkafBV+SXQZOwFBc8Muy6HnvoRzJxsbOphykQUBXl0s4If5uRKFq
PYaYlKw7ImGq8+oW/jkTQmUaZmdmyfJs12A1XqcTzN0XfZNr7yD/ZnOPpH4T
piH+lYtAU4db1TxeR/mgS9wflMJlD3/NWqVSKb2sYRz6EPIlmN7i6Nrno1tK
ecqeCErOd3LOSjEp42Pe6ybDjkIw6ETh8hGqHpN3zfiY2zprNg8PZ8lpXCon
xdnXWtC97SxIZoVAsfU9CMktyHI6ZdCSzaEAhIqQL3v7P47hIQuOeTDRqeB0
kr3iyQXvVOQ43b6XQ1JlenM7Uj7uHvInfF7I1/Ebfa4MoCs3Y3gkKFl+f4zg
yGLzCIjWsqraxAJUJHDwj748DQxLOmjVvNabYv4gibk6u5Rf+gO6wFeCNdIf
4Qxvy/sx+wScDpnZmbMk3OHBPJwXslZkjKv7y0w3RmuRV6RnATtOwB8j1Eb7
ZlG3ceFno0XKivautK5/ji6eC+uVWB3CmfdYZAZUjyGCiCD3/3fWltKMk9YJ
l/lKuP1tyojKDmaqtut2XRppptMEq/H8rVEBUtduTcxkUNbOQcUsBWuP8CQI
fyuLFmcPK2DizjuSHN9VhO0WhxxxN/iTgsxwp+mXSCofiRLNlEVO4zgijWW/
5MU5fDOnzuB9ihN2Qv6Ek1Q8866g7hhTpkVCHCkChg1EKUpESeUAEraQN9lJ
7vTydcX9dSw7RDn6GYSBmPwAcjKMYr5+LyEM3aGZoXnspRLVy3G8BweXXjp2
qdIH/YwIaJCg8Qsf71TIKQF0oebaDcu3ba6RTlxwUnJqu2JjQoBqerHWSUtu
fZlo7Xf9TrwX7ikX5QM92Y5nOgaVLzLAzB9W2jpnXLVNG1PWWnn+Frhki0Bi
4/pa+s4kvxmeUSkswr37YgnNEMmCbdXncPURLTgwL6PDt7WIKBl/aog1REI3
rOzCzEC7fj9Urh77Q9NI1xz+0p8fB+GddlD7FyzNlEX2HyNOV6vvwBToxkI7
WV+Y4fUqEVdSXSEaymJuRWoMJ/8FYN4bzvefN+jGN4QCxkqUaURZ76UfKK89
a8ZE6UVkcfCrRRUiXFe3SEH7RMHyECVSP0+gxFKnPFrVSAMbAXlN8bYjuoEC
2lcC1VPoZgTlCiCL5dmbCx+6jEgEmNmRmXUyAc5V54wxhcXw20cqIgHEqxDC
OP7OroX1eY6Gz1nLVpj6W13etZ5RPrhsAbJFg15J+Nqsa/McLgHVa0aY206F
yrwFhIviSYgzeuPgYt/DWbXchMbo6ckqRQHEFpPoJrGxeSzqzZ3dOazcSbhR
yogwEAV/a5yyz4NFYIhBaU2DWC9dqX1JywJ0JFvnqgu9PF0VfBPKwc9UKOBi
OGEUMCwt5Z/TqCbQpTSXIDdYxMLjIozB+XjAdQyhzhy438U97+VG8QSyrjtU
3oEVzLgsLaIhp9W2u408np2BBYun8zrbKsyZcoPyBCSoBgvlRBpYGycucom/
uve1/wXMyM1h0rbE4OLfGYEDhrPEEchfyLXZTzX5q8Od7iiq+EPCBu58B0+k
FfMfeiqOl8otmTz5TEQoril9meoRyWGm+n+MHamxdEzI6tOZouXNFjWXkYMb
YfvkUcZ6TwFTi27GqHskYWlZwvdXAQmcCGIT3iaDlk9SPFb1Mm1SnbicuFU7
iAGwTqv/0TYgvcfmFvdhlT7dfiXZuAP0F1eAu2A4/r+anGpA96tUf0zQJBwT
CdVuYxRSq3xbnG8B2xLpzt8MeZgsyZoFBjhY54pVrO3amdLBY2S5CzUhlNQe
D/eJiaEmKF1g4mmqZ5ta2DJkJqmOnHWpv2vRGmmUFBP1Kdg0wpp0gMuJUnWD
utWUiMH1YRmtERuA1PfKCAULFv6CUgDtoliE3afzG0k2Q1hIXSqGFeoAJgFp
e5Kqb2t03Y5gFSINwwkUUWY1KwFX/XcvCcu5ZLBTeFXfcvMf95rF3vYmovtw
q6Tcf81jd9m0FId3TYQLQYQhSvmIwVtvrHCXcZHPQPqDy0tSPXC8yDtdhcoE
0LftMJrYw9iKKr19hIoyVomZNAswYmr8nZLEGLxX6/TZ7J96XytX+M1I/dvP
xE1KUIgaajP4l4BgVccZUAvWX8TAPACb0vGkfMmGFq70C2vz2qbByJOPTQM0
YyMZam90WeW0WzSEjvKw59eYeF8U+XT2Esdddq5SYBkljFKFte/w3FP2X4sG
0b3Vp659+E++HTTobhcfEOk/zHBF42KutEVwI+o0V7tGVVdY0Gggk1FtE37v
aNm0CoIKWxBfsQlRARrWgWQvzQwaX/x8gWl0RjvZo+TPzRIfb6Tn/fN5/4gx
578Z11aIj0AwGEngTsa1x5w3A5wxpGEldTYwjoui5JpB2WgblaT/oQmGha56
gCYME6/1ZTVfQPhTI7I4V/LblNNYq7M1XYWh/ZiU+2Cw5AuCIK/8U/to3iLy
0KSUDja8y2Fr0pwCBDYxI+5iG2VFFN7CNMzE6qy9hcsOpbvdsgqHlnVY1ZPV
nLPPb2OqvXdNeaqf8j8X2zP3rt8x0KEklV4iZzkBEnTHeXZs7JPMzxV5lvC5
rAexH//+tu7s4jskE5uN5ayHdw1UJpy3xJ1dxJTOxiXDi6sVaoQwNcqLS014
YDIZHe1kU7C0MD/SnqyphgO34Kle2azmolwnJkBTNuHDwSaDNIo/Pjq9PSph
J4/6O3ywkFMTcRVolhzAoTtKpMOTiXSGqT2UL2xtVvR9l/2qswednulmlSCu
MmVvJSMWeTfAKYfrrWrDxQqD3H1yD3ou75b4YYL7+SAkIiKF26zNKErRlNUv
wlJ4OD8QnyHUcKs8VNNn8ZLUMym/ezHjJngU5Uh19XC24+pZlf2kzAQDD9oF
srP09Hfwg6iM5SzYqDYRwZu42cqDaMKtv3kTvIxNdXn7qwcw1sOnUtqFxeBy
zO7gj+JrI6h/z7f+r9qw/FuFu6w0XIzAY/1nGtjIUyjQemjcVnGdIjgSAodN
YnuIt5eUy+brY4yyeQLJ4yNovqQWpNYtRp9PcUKNPRStkwM3GDHB5ni+/skp
Rrb1QS0n6JFXDpBuTrcF4cpZS8WVwUQ7FXOdF1/2vnEOAf7LwwiJDNqBJP0F
XNvW74uXIMQBGOToyr5PkQmY4LO1Q3Uj8Z4ksAhXf8XnkT9oG4zGaS3U7UWX
m3+mjKnJpo75sz5Swwut4NqVBvH5TICD0BrCRPuMJz5PyZaBoAz4yoJHP1Gt
ENzgONnWTb08JavM9QIcjX749Tl30y7bcxa2RjvkgY3EE+mcxLYviqWwKXug
gPSoykDnhdqU4QMYOggziQVb0C4IhWJ1KC3e17N7lQwEjFmvLkh2quDZg0cI
hIsi1HszeIULYHyVgg33En27pryoZl5TiG5BG9X2SpyPgaf1o5T+pJGu2iV6
WrpRA9nSH2Ut5fy+sUEGsOHsHDc+N3cIQjpnQI0d5nGdE9wXODmtYXXChqUg
wUFf0mfqRPHuS5KhVg6rl9HQIO2yOT2LONYV65/GWZACO7pgj8oPHn/hAR07
dPIrIhTbkE+tjjgfhr3JpShKixkXdBxBmTP0/wFonlPeelVT+41x7YCwKN38
sEzQMLxSpyGU4ncDzOXK56Tp8q6ryL3Jebnggt+nnT1/FBAOCAji0Rz5Rkwz
oMq3ma4KxNRG4V4CqLwpd4fGG7vB06yf0oHH9NBsXQXaLwimnOIeq5aO5tef
GiaTObbI+0wMiJeBgepUfn/zA2mqZjU3zhCni2Xh6MnUqlV7cSHnVYQ4S0hi
i7K6ziTJDHl03qNdEAro/M35FWOqu9t4VYrgSBkzvQvPY41DUKHE2q8FwgP7
o7qSqylMZjLwvmDgk4nv14TEli5TQ1NeQI++j7mHNADf/O47RCy7Qt9tHE8f
ISuadJGsX5tAeAvTAL8QvAV/3Ytwm/+wAnYRbbobxI3rqriqpL9BD/sEFKke
oT5Ku3XfJhUZFPDlO+U1fSVT+UbRbJp2MSD6nKVwVjhuTPyol9gvwE17usGU
v/if05f3JFVKOxnB/hzbgah/zb1kn04eDycW5Aqwed1HS+HB8ipb3r9g9+TK
agJfOxPV251udrC50JG1B9g7cSTVZdhte2QheuWdXMNMvE+Csz3ywVI+W/hQ
xqS9mvYp7neOhVU73d3+5Hl2KOB9iZHdrA9XJ5IC/LkzOj0Enn1zn7s2a8t1
+2Vcif3mWLkbdR3aQt/RZDxGz+n/imrooaN/gOWLyHdvYUah375TSaj+SsmW
ZerSPkedIHSV/w1WNZrynvAGZqOJJ6mJkFG+oqW6z4OCEKz+A0Q7nDeh4Xbm
O79g3ysii5j84uDSoPKh0puS8Mo8b1lYG3O6du0JkYp22m3ugNX3WSqvX5l8
BFnJGWm62PV6K/yNuowPRBcNQyWfKohSCbuw9uVZ089sBN6v1HFdUf9ntacq
71NlofzC4A5dh65sIrcV9l5A2ooGyviippe3MJEwwvUrjD/OBXbS5YqOVWd8
MmAA8G70U0NSOwxwIpNsMLzRcKOZgJUg16oCP6Ac53vzSQT2yxgzG/rAlAaC
HSYfDOkpt9i1LZ+Z+LJQGKABESqzW3plO1cNgI0JpUKdRCx2XR+P/o43ptR0
14o60O7u/mOJUVvuSlm1x6+1oePSGz5kx5Mbc/3Yc8AmVb73ZKWyMileLlr7
hV8uoK1MYwqpKX6V9zigWTZBPlp2Nw+R3g49gtUSvMpPWojebGrRcxWxkWAh
O05XjEtn45kf4sihDSpW0yMkyKofAxOA/7zJwcTR1oe9tI9+OxVPE09DmDhv
5h7GsGnZjWzV2PyhybYsB5kDP0JHt+0fjryu8a16fRJVTxUdNRFUC5BiuIu+
qEEBnqbjjLomZRgmzH2Ot3vgL9283eOzvFibjnqS+iSfWjUK/jbXb/oHgIdh
KUdIWF4mEFccacJbVBDAsfLezP3eIwsrWU8PDpnoisQRh50EEiiKf3WpsPtq
trSB9Sn/09GvsbNeuK4m6wAStrig7m+MZbTy4JktWBLmf6WssDT+WHqcdnTC
vvLzVktv4M0zf3kRO+EIOYotXppWnkfifsqklmM3fBWLEGcwS01lF56RsA6e
mz0JShtHufAyOUPd+j2y2jBw9UwcdvG9sZbvD9oFkJeyEu33wN4iRitx+UBl
HaAS7HjJYE+IhVRnh3H7ulifsL4b5ThQ1JDGNTsqiYAylv+ffP2jZkeOTPe7
jTLEyQIuJNo94GLj7lRR/MHt7RvvSUh4jmTLm9auSfPUsBczmfgk4/u4f+o2
a2Lmy3upiLOrS6TWuMm2HHNZRkze1APf7QFGdRUzeiq96H/bRb7NNNAu+aES
Ye09EesJrWlIH0MpZxFMtQ8fxE8f+H92QnyVc/iavC/G0q7mEv0l0lMeqlNx
q5MVgP4nrNoTIm31Ks/7CP1j0la6A54IQSHPZ68HZzGv7GYe0x29obQTNCXo
Num4dTrUiaG7mNjA+apG1Vzl22fRCXqZrMwb5EF2F6KN6JRXe9AcLgu3I3Jk
lYxn+snUzGoiH9eUCspfoFy6x0NvZdlkluHbKgZsfuEdAStj71a5pjBIX7B/
eGihJ9SLHqtv3x7WQKqUHgb9kKpbLXee6KOs66AZW9MN9pdY5RPJzz1AVACG
Z4EXbLjQM1jq+1tq/tPqESq+VvrOI6LY1N28wIk+2jJlPDHt0jAz1SaExfbJ
2uXwSszc0bu3iQwCbyhhcjqLh2B+MfOmGpDUAViwTNbN6R3xQWoiR9S7NYg2
etAnwFx/Pon1cAkip/STh/GZsFEQonHkZoITZ/e5Gvkxp9zcgnXXNUpurrAc
FmBYUIrqVmeg1CKKgg+/GhG7QROToDI5hlXjU7rDXG6Wiy7zqs5UA2jeAw4u
ZE4QfazER7cKSuI5fSIwgsZnG0zokWEQi8xPSPE++0/cjILbnx+94BGB8JCA
nbFk6JYQpNiZa95q2nKwQr1P5nYtxAS+uSngWqV6MBjEgrK1V1ZirriUZIFM
vFzYVnpbN93rNsFJh5IJLYRkssi6aYAD0ehlBHo7DynoGJWsIxjPjjQTOB1j
plwYoGU6Mivj5KTF1Xk7UeIFyQblLopInAWRrLRQzycBD5GYprGEuTltRsl9
DVbtBfSwi+5wfZRM6RqDP9Lsok1dhd5GeoZ+pZaE2K3bPdHDIqvlEeZR9yJp
a+oKoMBk8n0FGyEgc0qknq+DvG4XIjabsqylBVezR9HzDTODVFfDFvounoXY
lgLUDPumU+eywqQ7WdftXgrai4pjX/5dhzexJJJ+cuehxUIgleouNRp1krC0
ySzsAdpKVsodawJPdYP76guxmlOvXJWONWhx6KSb7yEgLljGJgKY231HJhwh
pJO1ugaAh4EzD+TuKAjvmWa8O0fJlwHVrFx1aycRcV5qRMM2kNx8ZmeF6Abw
MZotsq29xQ3NI8vDOkyPVvS+WXUorSq7Pc1yHhY9ecBbWuG0LHeJU2kFWa3M
v+CVfesD2zaJXr7GxCkXdEXNhSfjmsnSy9SvOcv5/+Oaa4Jwm95167Xg0kdi
kUNzybUHheYFcNiN6qHG8a67iRDjT1agHvBf5JlCqcz1fCg6Wv0ogiRdKqju
3bEtJfhWTOkeSDD3IGSXOe89l8WDcTNTq+4RUFKuWsSY9nLFE1gF+mukkSIt
+q/1uJIkxJCYTQ4NQ0GjajLB5bQQAFVK3RI+NFj3mWfaUgOmg/5AXQKBVeGL
9tn/e+pvmqJZbkOoSI0B4TG20kvxLebXYNMkyUBg/q6XMt2IUfJRqh29E2Ds
8OlOefSIpkx47QMX8kQkt/iDS3Eg7NK2KIBi+61EK3iov0O2MSFtSIxAbTk4
L+tV1heL78roq8I9ZcNPQ1w7F1Ed6O6HUWHVhYBoOn2fVtRE6/C+gcDbUROa
qJRlADqkj++yWrnysyRMkr9alRQGhXal3Uy2G3Xl8l3oo1xw8teu7oP3itdd
N6DzddLp//KN3kPX3rSBaJFvTpr7pYKo5Ar2ZOFVZ8T6fWRlYpsa5RvxXfLs
59tVvwqH4NBzmjPzcjIdf+77oULif1OEyqJ21ylvmItE32QGes035+pbktNp
KwBIspnFCZbLgnoJRqA1JPTk+a3/BVfXr5MxmXitrGjBeufh2VuRMwCF3/8O
VCjLIkWklSp4+eouSGwtMT//xLShZosXU0ODF8F0YpQa8AatLtk8Q8NymtiW
kNS6uXEGzrRvfHIKjYKSX6sSY7UxJhfp1luViRfdiknlqhuHb+VrbWb3o7vf
r1j1fJ5Y33VRBEpWrVVKbrZJEBrLxBRxXPEykHh9dq8pPKX8P51SZ1PIkdOc
gzys9N7igjX2LA2OPudZvUedyxDkRYZr2ghyKfCiai9qLbo+gTyWhAiJ3fMj
TEmM5qayKvA4AwpivjQq7DRPlO6tkRBb1sxBquNXmjUdrNKLD1qJSuwpB0W1
ksloN6LgpCLIpL1huE/T7HYbfZYPIGoDY2xfaY4LQjJiUuF2ymY3g1ZcRABO
i9byt65eq2C1meeJ3zWLabJ8kXsdd+NM4Ij7AXhUjHC6tqoDP0B8aVgbr2+3
kqukYTw5oXJG2J0I62kxsWC3JNqC1/i34Dm28ZObhiI9hz6thbrxeCE/Ej/A
S5ljt+NwkVLMMEDZcCZ1AovDq2qCa1Zatks7BrPrbSykmwvuGKgVjWH7as/R
4bJsKGxlRdGULGXkqPgaFPrsUew+HY+tvkgQHZaScs/8LydaTM6zPIreryxs
cEQr+k4fkG7ZkHDZ4wD9nfagYF3hKPJ1rTDbK/Vp5jsYORexaEO4m8Z4+b91
axxb8mYrkfYt80LNzgDwzojgp5rOaAGBoWOnuxoyyw6K1KtHs+g0hp+9b7fQ
LNGWABVKU+VdqsJhHIoMY6ESxlgC+OR53jR/BJ1dSAetkZ0F4gXe/JCF+GT8
pl3wnDEFs/YA9SiY3TbvkB8OT+UHTfs0ReYjUZkHzPjH2Be+Nhx1x4rPSjGz
MsuoA/AJXnuBjwFmoaizpB/mW4pWpqFkcVlERc5+3pqNcJHOmhAL8x+18wJ0
bbdmmXYjguaHYOHUVs8OXM1q7AKz7T16mVrbpYzpX4gr8D1jqTOqpvn+aNEQ
i7I8s5NvL4Q/vM6kM+R9U4K3QrrkG9FPVIn3TAtj7VB34k8UbPA9Dr0IBEsw
vyYb8YniGDn0Hu9gwwTD7cp/4JuKhybw4Oxyt1Ka557swuUtR5X7rmRQODRT
gyIGTgpkobLLXb2ZBD6oQousRfdv7d+18plr602lZBdKWlkwGyRlPIVp8EUT
1J4CK2oXUSUUQZN1Drh6L8xlV7b4HndC+ZFWxdYLlbRoV3GNveUlmTREoIvD
73qO4z+cglYsRL6Mpc3QlyOXOTxPxCEOpyPL8WrJp//NJFy8Ha7nu2zPlFPt
VCg8JsBzBJbqo0lAPYqSuhnqyahJx4AooJZS36dT7VVDP+wYnj2VI4h23qgz
O2ijKEpmpKNnFblPi0iZU8xWMkpCTofFWXAtvpT8nGJW8kezz5AHKsbqfbtw
6sWfoXk6lMYbZugTm1jDsqr5Tk4ynGlmKnDEkVjV0WTRRC4VCgJlHfI9jxcm
R8VtaCDLLIq3bFYNfMlRadg49rtT8r3g9G6ejgn91csAQ+akpN6/KopmVIwl
04gdIlG3yVnRtnf8lWVD+LbJcvAkniqDOVd6qA/jqT2nr/NqMuQBO493+pMu
FREAsuBoqfnfSs/ecJ50bRGpOuBbIsjQF2pwPXfxZc1Hl3sh7bcfZuLsaTuk
jDq5+JiiI7RL8mnR6EQyr3wXBr/fs5tEOpN1p8yWbweYQhw4r75RHbuwcuIR
Y5CV/34cvrWF0/G1ReKrYaJtKSbqzCqMljjAMId6V2SCeG1FP9Jd040lLSdC
+2IFIv+allxGUwve0PyGH8HGrCxwVc4WGu7uSK5rBgQ+FccnxpkKlrr4CzWL
Dwmli90vWcgem23fmQgYOG/2R2d3xOF0BKgwh2My5dL8q0eHkfL2qBGnV4u6
Z4zqcIQVurhaFSkq2zJix+CGAwPgeCKX+J5nRr/6d5a5ofcfhlCYs2vS+N5z
q6kPKhqCIJFEuBY3VR80kQDGjY2dsB6uhztvwsY5lvHdP+MQPHJAsNj3/gpm
jSFpjA35XZiin87DJVPANp0LaVsdgSGL46oPkq9id5rZHqfLUxzR1al++f1y
PLXbHOy/83JiXLm+JQbPSY4r2uBjSuK12IyeZXuOjHrGKhOrOmWtxwiT6BKo
y8fQQBtQZM8tM1jMlz6B4rlSwCr9TQJgxGO60H9ISz9e36JdC9NFaiLWw7+w
svxiZXXUBtJw0QEPJaPAymkJAZLzBn9rOnwNUgW9maFsS3I9vzGTxxL6qfx6
DqFN9Ywo+Ev5IAj+uDt+jQiAzfBCbVKKjIrXfeEHCwvb0IUKAUZfbs3TSoPW
g5VH6p3XzBNpWn9Ag/54QtaYgctybmaJX+v5j5KaDjIeGwrH+cBuxZNZgPQC
+gXz0n1b8RKLtFcWoCtCoW0bxXQYsXy8ph9PXDhdpizHGCo0RSFpVKiVHNHT
zAd5oM1Itfq1nBImUYBN5oQMnS/5SRYVnUT2c4r/sxe4c4lpw5NWfqge5O63
qkMYpuuATpx+CB1Ywgvf+ttkDmZhQyf3eGnFIADKpo9juUXECiYifQfAwx8v
HK+KKj+K+Mmr0G1/PzY+tJqne4E/jYadp8aHxzTj5ojz0dyCaVL57pAH9ns4
4fwIrcv9cP2P2ml7ImVrfiKtQ04HkAG8cmr3/Rs0Jp9DSnSe/2dI2/SmnoFu
9joiCkje0KJOCivQqZXEgch13hGj54Pl7KkJRj4yAywzlvP0KdNDmVFAEgAL
8zSVc/Bt+r6YhogCD4kLJpYAgdoO/BMf8fm611Y1eC3pLIrnRrrn7Nm3wh3r
MYMPj3vsJdL3mCe64P0m9W0btNd4Qv8c14JLh+YDzaWnHi1KnxzAXdnYfKpl
5Mw/qEHog/cfnDQPwdxgcrJTW38Z5/DPscqldKzb5mU8HKyYrRQgxqYD6QQk
9hs73LU3ZGiP4Uwwnb8eCFxRuEDi/V+Cbbr6dUXA7wyVCPS1Pe5hB6kLr0Wa
HGfYDT3gI2XPYqDmN5nV2iEw5BKF4Et/54DmUxkKlVc3Gyh9Mg4Vw8FGQbhj
pnWfmmra1Wa0l5kazPIocv7Or0E7A52tbGUGKx8snHJe9VP3Fp/aycFEnEIr
IByqAffMEZ13QaYgdGEBlKbDaFM4Nhpmi90gtkMnSuJ/TwZ/kSP0bQ94P+Sk
NSi1O7RA2FS6myNWPhqJGdzMNAk8iHEoKJSp2bcQxOlcbz/4bLayDQYRSTvP
1aT5LYE63yrdcZ0MxgYKAgtJRSNkhbm9Aw1Mm1EyuUc9DWZ2sia3URs8BmrL
4KQQ23kpyJYAvWxABLfNLfRHbzFW68rW6+Och/AHEqTGfGcZdUvlq/E1mPAF
XWg9L0n+qaaHwQCu9PIvZ0x8d/xeein9X/s5a0VKn5vm+8SQwzONne97QDgd
thoBcKBLO+JkKd2TWlJSX/J1LyLPFqjkIoCs2mx+8egTac/G4sOSN+AZay9n
nwE7HUpuCa1OKBTEb9IYYHW/9uR0YJ84VVTKvTVrvMMPMYh7WkzyrZPVOdm4
kNFD45diKl7jBB09/AEMk5KepSQJa3JGGhz7/LxiQj4n2hNzWoOtsoMQWIoB
0j6GisSizj3ysu0UGjm7AIh9b/bPhJdhggTtddqOHPYuybPWFyZxrftGv5ym
cClXxUvdVoju/keOzqe6yR1DPrfOFg/94aqBE+d8ExwFVpCycXTgBEj063Mx
jBsI16JMWXVO+4JrBQuSMm3zIiN5GJV9gFuyaeN5wYm3w4Q82iGfmHCiq1yd
02f+IHtrUtTjkdx8JOkC8nkW8UNIY5WIi9CmHtOvM4RU+mpUz4LYqkvwgB2l
2RXw4Yjvx6gIMofC3jWA/0CDFbBp3CoqJbTiKo0ddxSuYxhiZ8XhEzJQAa7A
OovZfu7VnLYw/AK9UgWscrldczxtUQl26agPz6TandJCvATbJOqa0eHaTB9e
lj5kcm+1J7bYukbXvMXOipfTBZdIOPW8QFB8+WqN5ZgeY7ZZ+/Z1vv7XEoYV
WXRPynLS+SOjvPAoOr+6AvoMO2tONw8Bq/ybuqYNjx3kKIH7iW5E/EEXr7Y/
QiklB1qLWUP1ScRnbRwuWrHjp2sH2GbJiQ27avOLNBmP6zAkOrVLP5UChn9S
JZWni++DXxt3REnDxlJmJJKexsb1BUxOxHiZw4250S0phg+ldKTgZtjNXaeE
2xMh7RK6BACTyBVzkYklSCSZsVRoZa8fTG07wuiTTzfbt4dlwF5jK9CUhG3p
/4M3ioopRwjpuylTUlDw5EVVlxjVOFBLdBrpUg4f7wEyt9S/Yot8CWOfLlW5
it05lJyZ7aUJX+vXRF31MFUVRAI0lRccvLOTIMOgFeFdr+lH97aaw1J9VKLb
pegt5SAYOWXQfbSvE6llb96PPndE2hy8BYhc/GQ0BRGTHD+8K+xP5y5o2U8h
rAyCkHoEysdQVoiJ51D7c0wL/cqCSuDrKzYZmUg3621sOwvQXqRARG3s7XXD
JUoA46wifoG6rYSkie3mvnvHyfe+98h1ry/Cet1zTa3kr0a6j4ds7GNJQgt6
KJ8l7Pq89wgdVAQzenvDAic/SI1dJE60/dJuvF2zTbDXrzULN2+vqu0OlNqz
pOn2itdZtS1U9Pv4c1XOobxCRacg83UI4NpvZV0IXLvAmqsLc6zF6hqYCaF/
qsyj+yVrhB5QnK4Sw1Prx015UkrBHKQcyjwYWAzdSl9Tff6r0IN+yKS8OSsp
2vRxlUHjqTiza4qnezyItguhyFWheOq4eNH5mqfWPQ7m6oNKfNpNLLw4xwwr
jUF/tXkgqE4rk0Tb3Okz8rpX415CweinTSRLFfT0IoUn0dXiDWG/2kUzIPSP
JkUcyyIwn4fiqUet+x8s0McAAJC0FGkhQxKF3eKY88k80Ka+9tZiSpeShF3p
0CxtN7KeX4DU6k/VtmgwZS7ptBjcbG5l2mi+lmWnJXvPIelS1zPAmmRmR59x
K782u3yLMXI9Fhi5A/yASI2Upp7WFXpgAur6n1vFK9VDgNkE1xlg0z44KH8e
oVupeSSq1wXD7aTzcxhDcyo1chDUmFksm/G3aocKgpqdGXF0TP3pvJwOc/ru
239SQk7YtS8s/I6sWbUQrH4D8BoOumLCAZ+CpXzqHzwPFszsTCNBgjGc4wD1
E2GmbGUAlop+ZQQYl1U0yX/H34gjPBlNVg4WXIJC/kqxVR2ORwbx/6R2t8lJ
TsD/hi1FkAMAB2NB5Lq9qkRpgnw4Ah/dPsSD1VVuPnn6zxHCj2lXiNfWd1iB
CroTUaetlOTKaUyJFLreZKoElTVNkqV4NTUJZk8p85hk3llfpRDBC93DkKwo
ZgM//x0PwUnMujbv1qw2zwgEtKBDrwWnKjvTKfG+OLUGrdHziDvU46VltpPc
mSflixhpxHaF6G0nxMEin57nY3RT3Ak68F/mR1WYyCtttWkVW3FtZmCTfuxE
dFTaYHY3U+ire1r0Kr8UL2SndlCylgTGZnxPnllmqOFRCdOUbsc6M2X9K9vi
g8oxac1ErpfBkWLetYb1ZIBE6O/U1SjsWG9g4jW//g3NUUOR1mevNusYmpCV
QkCa3AQX71i1lCPFg9w8KcQJqnCDb25Xj5XFG3hGrY1VVD/HudIRd+xP+uSt
mMZfTgwU/HoXPG37o3egOz5Y2ZRhmkh/GvD97VmnoWNrcGwbtA5FDClHL06G
sfqepEDOcJyCKh4R//3pRDwWUeeECn9NRPi/NgoG7THXw1qgKBZjJuTXeiJh
hKXaG5ahpAGECl72b7wJvEw66Xl2Vf4YWFG2O8MTBvlehBF8ap2c5woA76W3
ceQegcLiyyu+LZ4wHlfvGfLQkOV3vYHR5LrjwCbid0XrGpSIK0gl5e62Dnp+
XFw1cJxoi8y8e18HOSWm5P7BHN8Sbn1YJwkAMINxZYFdNuNvNgsdOc4AeP8h
VapyeaXP5pK322vZ1MSIxQXWyXsylgHcLlnFVF19rJsAK4qrB4ycRkhIPXQL
JtK12Nmiov+1a7O4vxgZVBrQXuIYVcCenwsJmI6oTcCXRYH1J3MKpmZxe1E0
lrUkhEbLymCkYBPP8m/8ZyRwDH55am0l04dRj85eoDO3fFC3HLsBFZaMQ8VP
8WcKbykvYGuxdzoDhLobBdqhZdhzkYeSSpaHgLcn3IC73ziyGMYmMIQYZ66o
xE1gzJ/OCiWBpptSbEgbo30Fn0ZvWx2+kFcyOhCIiwZlokS9w3zb0V0IqQt3
k8ZnbdfUpo7xQxX2HqbrCxW+ql4lBKveB6snuzSs90zpR2LD2CEh3YdP4Zhc
QI43L/1qh13LsMOLGMShInO4gzRH4EuKZ/aqcaeVMgAQ75UZRuOVG0p+KjIO
q1OGWBa120qK0580pnmb+K724qO8N/3AwW+ptIgVEzO09y6K8BNhvXtn9Jtp
u89Rm13KVwNj9FO2eS06+HFkWTNDM8sDJ6R6Tsvv1R+xY+wuah17M7ihvpWa
icKIltnGWClBTpPKIEIIucJG/+QVHZys0e1V6mu5KF6pd7TGsQdsfLisAgE5
7YljiNwfBOjxt7xRG/VDXH7O+3Yya2jcB8uVBQVkZf0vmlNFhGjuU3qio8B6
8K1c5/BK80OJWFT/usMikSMJTRIdjDEXf2oLDc9/SUORHcApzU5ZYhnCfEU6
pZ0NlswJ67iNkVKeMCidb414WEqtanoLBqgbAj2KZGEYBHT9UDhBSp6kSR/8
Zw5azxBIfjMiPYvMxFsxJMHAsX5KUBt89F4PbRAylh+qqKDd98kwhWg0mfSU
mbtwxyVfyCSpZQznF3h87K0/o4RUW8MdTFyCu/A7/wa0IYX1Img2fHHN66Vd
KDDg4nULyr/zL/hAAlW0IR+VVg3p56CZ0Ul/ce11Y5bACUUHIpsnrOqASEmJ
I+y90hkZ9DIrj5JMzUrI84haaHP3D7hJojhm+JRJW7oPf8+oRpDOyBc/faXo
6httY8YUvaazcItsniJeR3CfcDcTPFwljTx1F/RhLSNWz6FX0ITnnbAG8mv2
OLzgvbwOZUxKR7xe6hiOp/OvH3yU0yXd1hxO6Ft9/FRsI5pD0exWjVs3yIrc
qHiuNCFzHnIsz07lFRKkLvzatW8NsiE93cm7zqw1euzS6xRFdNdbgX0SZHBm
qeezu7ug+7t+4v5NN3Exn/rduzkP46MuFIGrfadr2QyQfpCDXac1GFmRLqwY
XhVyqu6tfeCEik1SmzuEQyiBS22SHA15NwRRgVcZA0hcivfH06zsqr0cbssN
YymrQfd2mpfTRnFKEvZPVS+AojEhnz8XpII2E3XFDy2Zi3tV+9gDEuKDzxID
aDZ9JGuOuRGNm4KYTsqKyn/LgOaMlrd3UKe99aF/s+qy7WzYNSoT6a0G3h8Y
7zV9NzHFdsTucLRimUXzNQhL+Ih+eoQy/Kl7422/+86PaW2qvxsQWO/kX3Hc
zEE2FAOXQfUoexwHYHw3DA9QPpQaJqPfLN4xT2O6Arkhuq+acmh1NTqhKqsF
gKfmczwlW+G/ILSVI83VrGKOAjziGR2nwQ==

`pragma protect end_protected
