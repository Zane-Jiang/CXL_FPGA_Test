// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ciy20M0RiS+kPlntHqAyOKoHmK3b7ZGFsFeTHHIktvJgBFZwyE2T8JX1Tk2v
HbdQqTBjPiVgGNV3mPxpcTzOZJ+IYZlJyPJks4kIqK3dLEevuDZM7r0d342q
UAcWpXPWWKO9tyrHEXlDltJS38AQ0/1Gf86D/STmsiBuw9cYu9JiA6Z+CDSx
LFhRn3BRwEAs5nnyxOLp5RzDz2kBHjoDnE5wRjLPOrYyfS/fExVBfNsAlXf+
0VgbTMfyKNTC6s2NqxYP0LpqRUsQ9RmC+E71FduBl4BmpU0Okr41jyxraU5F
+ejvxFDzCD4G/zwNV41wwCsbY+c9icWqoWP01l6DlA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MIBWSjgYl8piY0YCneNP/xZXkFv3tUETPmStjI2fQ4/aPLZ6cXrosODVffM4
wp695uySsUkgO8vFdGQDTuobNZsMw23prrLcbE8itE3tlmFzMYc77taxpMtU
7E77eiKPJYSScqzdWf1xx1SnRiVbB7n9in/N3OUWMFRKRjrzxeNIUOmrryK/
Ogk+VvhFBjrVVzuWWlLMLto1mp+QOiUKCrnoxuwYTdAJ3kKT8dLj+HSLwNh0
hcC9Xb7mT3xiYMf919hjAeAtVc1f4aXg9TvRwVeWiZ99RuNCsVtODbuEQxTK
UGLkDP+nMSAsIqoW5Qo0tqoapbairyB0Lh+4VyCl1g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dF1TaTW2G/6JKLAHSJMK9zocEcVei7tDlhZYeJyipgWVbrfhDO2WaDYABWL7
nK3hn4HUpccqvLywP1DyHwtWjmHSXuXNoP9gMJwJ0qXQliyF8QZCiUITgumc
5klEU4qMclErdxR9ffYDVIxwa7b5G9A3xaSRQaBGEloVDK0z9EeQCXcbQeAl
ufXglEHEPwfz7qCXURCcKW4yqcGyv8Cq+ZHtZgIPjx1ctQi7qwv+z5voDc4x
6UfTLPitg+KGAFMuJPJ4a8WtrgOuFRLNiMCchSrAOQoJ7q1VskJVH63C9znH
AtuPotzjDBbkf8+6+ogbVE672XEFejeJ76zBGeit2Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
V2g83zSgBWnCv6qBd2R992QHuxBdNb65mrIRlOZjjK+7VMH+EOsZkHxHuMNU
7RPcbIjsZ1/J+GWXV4m7jFS7zc3dctQKRQYW7BVz92ssRp9WJZyoZiPo8ZZc
xcHBXJaTwrOor9ROmFnlNowiiOIa9SF0xv820SXyH6XKRo/mHrk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hkDeMOKFBj8xYmqZzT+5PeZvspgBMQHSmyeE2i92Gj7RhoU9nQ6qUz5KBMRj
vkciaUfyixj/LvvB2QllNCOZCb/ZcVUNZ+FaBRJKdSGCxqC8TG7vKtd96eQJ
h0jV+U3ZCEbErRyWa+bAGuSscNkqRe8N6Zajc85cHN3iB/u0992hZqWnCGJO
ATCAUaZxUrgrnvAgTXiNJPDbndHzizJIDq/AEoIeS7mjMhfWVHvMiao+4d8p
Jngxd3MJUzVxLM+ADRSd7AU3e0kQ1MvgxlWEQ8bVAQgD9U9ZtrqxcVgQNwxY
5ouYd7tI/3bNkAjEuP7JYBRxplh2ErMDIyCUyWtmEwzV/4Y13EoqAsI0Sfh1
mmf9Xyca61f+kmXet9GH7fgXbgrwh8qPOvRiwXCduxpW3741eq+eNdH3Nq1g
cyyyA3w2FlWIJMcAmiceR3bjfBcJD4BXQWlPY76BsY2M1OFYgsWXx5f4tIKx
ixdrPC95uPjnUDrXJxBA5p8OMeNSzfbF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sNL9A1NBycebjuIffJTeLTjpCfOlaQlBxzkBAXbkDpI2cDTFHwD9yYRJR8c6
kRorwP8Jmy7897sTku2ovmvp5uXBgyrereuB10QmntgLfSpZPnF68W4N20rs
UUMMrkUN1f8FafCimkrLv+LuTUxm+GxqZdEoJQLtocIE6vh4VzY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EMGlnwsDfdqMiV19E2mhFoMJOv56gCx0mY4J9K+TAlK/SfYc+2wLxW1RPEuG
7SAaSydTA9OPYVLYLU/p+1ZzfxBoKyl5bH9Lgp/v3Cd72FTCxps0KZ8nt4kR
KM3LggOobg0Ev8g9z4RAFaErR5pJFMKa4kpyQaCwjaZMzdoJkRM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 143120)
`pragma protect data_block
QQoSIiUsHigDJF8YAMItHQBybwWs/oIOwWxHnwKuLajj/2EwVi8UCmh2uq0P
u0tuP9LxgQTEXl7n2t3avAdS0nLG/gYvQiejCqW1JJsl9SEkHbogitSgBCKH
Q9Hh/czvrDA+uWoNudUmJNGTz2+Fh9nuCfuxeREhWElqX/qgmyicPzLTrLoE
07bA+sHxVeicS9BifCA7V6+1wfp9CX++YyyDQkpSK+phUPKj0k8Ptt2X2t7R
pPN8nTimXFTm/akLffzT+8912PHXU4PVDLkmGSiy5ldYBDicoPIocgegxLmT
j+efZhEzmqncYe++koKIn+3jA2gXmsdwjgB9oCmqu8XmNKPwKB45lzALmG/f
ECsSeBy34w9LCcGDrvxO3C+isZB2awG4kb5EXnj8of/cDRHl7yhQKMMhRq8/
VD2KA1xJtMLAKy+iyY2YTE1xFQ9sdnida1bxbTjGHlKfrWCh7SkFnlnFPf8i
bNQ5Q6/Pn0bX15CTK+yogwPD+RB9g2kFkRdP4YDb+mR1BoaZ9gCrDGZvO6Ii
XzU1ZgqoisLPr5Yddidno50ggRFHG87r0fKGTQvswy7A4eisN6g+X46mLO1l
qhoJoDxU0sGqGOe8wOoJYIVr5hSih7ZJg18bCxJTFVjzomnUQiKdXVJJBE2D
AMn0Y/w35Ea2odMQo0V4GceNYaYNi2zWTUmHb0Q6cLQTImPo6qIPkdyPJ0B4
vbS/YY3pbrE5YnOUtcxMj7hKeffe83ETwQxeoaPdEyBA1xjoOIeNZlrxfg+K
QzR8xqPfS4YlNEEmBefFKm9MD/LDsPzjYC+4R5FiJqdYEmRmaovwZQq3lI7j
sQT13X29oRqi75R7ApsVzAkNqZn+qvV49ereFBj3dKAuoJ4xYRUnngCXQ40H
ag4OrBLLPXBdA3V2ffY1bqFu4HdmY4YK+P/F1Wzvl+vKDeVC48HcPtsiGSvs
hT70xL6jOB58wt1GxzHTIbapJUoIvleq5VqzkaZs1Vkx3a3U2geek+9G7xEU
fCKdD2l3qVtgPsOHaZk/vWnqlT8/TeyjjbuMS0t5V5HgErUqqhMjCEYVsbXt
vghamC28ATNrI+0dHcshab6iXZpFbcJTiQswpIA0eJIuvVaVA7im8D4PgjMX
eMuHAL9736w4JS6ytLHCxLQ6VHRFpB61koriJjDnfPYQs34etYaT/7GMZDTT
7JVsZYunNGevDVs1Py6aJtGA5SAoH/JHDTORk3Au9lOSCYvWgTF291uaEB0t
FbOWbBKia6fhndEan42rQGdeTGvd5NY1xSUPVIZJZNYNlN6taOKLPJZC5Ut6
dAWIsCYm1R8PkLqkz1ndpMTpO7KAIb007AK6cP/m2gMp8C8/azxS9yeviKh7
ZPRgm1IJSzuaSYs3k13cWTF4ain73W1kPAPdWaQHG4pndtPqj5fvAVQLnqGs
cWOvtLH9lUXkE6bTKiB4bk/eqofApMkmqkw3mgHACOmCJsxAOgnvUwSkgmd+
cxocOyCkxlnkzFoQk9EyueO8X7ClVqYMFX09ktzItf1m2uQfAVaLpQ/SUXOc
Y7FEySo03IqQPoiuNOxR2KVApj5M8422aHyOSUdcJzlm20g7x8FfCaNqh0k0
5YKQKrdQYJniBN7tHg1UolC4eWW/sFhtLqjuYCgGo8+iu7zpCrggSj9UyY9b
cd4ZEmXNo3s6CQhK8j4T9PYApn0S+/+MTi9tM04D0EJw1Q/yCZXoRgauvskv
LiICeO+a2+DEAmNylw7LK16wVqCU0uXCbiPMTBq7zdgsoQxOsaDMd48NI+OV
la6yk2r1FJ1gqawbvvCVsg6UKDKNvrLY6FPzZ7PqZQXxaNq2lv1zpdr+XkQ8
geflW/LYB+MSNti13SHYi+FhiibHtwUx94908tEVTxI2GrxU8P4jNoozsJVg
kUkD9QR+GmwBOX08mbzPbu4rvNcOzADQgnSWLLsClrLIV6SVu0wZCTLuqIRc
P65D/B1TQMSTvGDq7x1O6fH7hc8a4qEr+Ajth34CTLk6r8RDObUE+eoiB2gk
GTTUN7/fjS0a/DoDcg2G3PVavk/1hT9Mm4FP5kq05fYDa/RI22YSV+J2zWMT
aUMNPREPPoSbLcgiUgwuOabgh6dcA+5tLwE+W0Av4ayBTa7P5zn72TTSZUlW
/0LXHBpK2aYa0jKwg9UcCibCd6nUjVJq0zDwtnjwPh1VpnWEEbaKoa++wIpl
O666fVWQLpocJGwEjIZ47sW68TEaRfaCu8Ogpqkv/F1VnL8Z4gjtdXOcwyUA
1xTZKwJS4xrppTmuJHJj8wSV+E/MmjAITmix98PO1VTHWsnrfw90s2h5+A6n
RzTxYh+RbBONUw6cIVD39o8JuQMBb3oBKwF4HcY/gfs+d1FH2Me5SvVim6JC
NzJJRw8rgBkaHS319Ywz0fS8xEF5UpXnuF3VW9xu9+18IA+bEOmrmI3+PTOp
mK11AUXmQm7Dk3h/B/QlY0wxGBlcb+Hi0NP1vEOzjZpCdsmxUliKEsbjtnOx
a0db412Bh9taeVuRz8wAN6+qUFX+B+d4J5EiLq9KRebiTtLrcDxgFoXlbiGu
iOoWTUNAYKnA5WcjmqrzVZwykQ29Z4QihKlqvjxgLlUg3a+khbVl6T/KXnYY
WUZprpGp9AEtG5n97WvcxyRPL9iFW26UDT1Y6pN/3T2H3O/+KOyWH5DN/7+x
CYGjv74waJHUaH1PTlJ2CYbB2gpGazngBl+qC11oxRlmaikmJ0RCY9/sdicO
TeGcUKSw8xRe1ojMw7Dr6Qva2syu6UnAsNPNf+6LRTK5G4v8QSuX42SHRtyT
bjhUD8r1z9q6bYAW76d3t322W4oSwU+BTcDscBh9yW7QWumYpJ6Wkw4wjDk1
cDZvX5l435/W3Z23X3KTeH16MRQQSWMQd/XvzqDfYRbx42PrMI/xG7l5flna
fOQtDkvnOBAgSE4ba0Vy/2ontZXRHP+zLDckarNFqewBWOUHNVnjO0bDC3jR
t0xZfh6ohaGAwljCm8dn+sjf4QuxSXeQ10FrpepKjW9uGuVUHluWCFpyxsSz
GBQocAxvaPWGTUVV5POQ7giuLwO6VaXnLtoeQcDWoWG20mVrV0ZXc/EQ6d3g
QwPvMz4bQH9FRd9bI4cuaYZ8X5tGspCpQipgvq50xwk77Cl5vn9aec1gHm96
PzC7j1n9AOmDa1CyAyRZDv0M7nKbIQ2/H30lEjwkBqvOV/NTDoyIvYItitdm
lCP/xUJp2HHIfeK3Tf6iXByVt4NBC0SCgvzZYO/w15AKvT1OCnIzouDjctuE
3QfLkDa9Ybntb7UFnJnwp4ZsaNzJhg299W3OncwTjcvLBal6RLViXWnBXUau
wxzwyaqdpoEUlJXmJqUKS876NLAjU070GMcvUtWGKahyqGhBoeZey6BZz3wX
H0EmLilP5Ibc6bDhbQ2iFCGk103AfkOEy5gXjL+R+SjXNW9kWzAsRNJK2hRt
Hi18+jUHSzCs2uBM/XzfLPMfvrrffaZJTSA3mi/A5JafkoKZJLzokDtHfCyH
cBVbFtsrjZLigMr8s56tk5x+qXCNOx3a5f881MNF4xDFsLhM2qqRRLyQ7fr9
nUsxep9ZYV4+5lY1lHV0nUJjPpLv/E6hMEu67bf06QWIwz1oZDNkzUuIBAuS
V/SJQ+weWL5i7MQIhYudTQg+xZQxWtY6JPZAnVU8VI5Nc9NxHQ9u38RoO7fI
5phukbjQ4sgSsYiVRzHqk9DussJjnlC4FWqqywjhUduMzMND2uM+dj4KgaKn
w6+cC8UkWyYT7VvYLI139yyvnlwifnHWSWevb37Qu4wtbay60SzlEHD3e/ys
29aL6BjEzlvOXrgrr7KZROJL9fvyyOB/Xg8JYYAm08QwhzrBpsgC/jcoAcZF
fyBFKjrZ82ycgOS79JiUxBeoXg5rLitEtSDuvLllFAUZRsyfsm7Qbztrn5gF
KfTdvsxZp5dnRet11jCTa/hl587St/OEY811vjqpXi9dczjbqc0PYdltsiAt
z1QMzZR0SbF66iLrEMDK40He35PV8xTK8z1jnLuNf807pSYxIUjt2tNLADUt
CMo0cPpjc0NBPUu4k1Q4/MqsDrhH7mZynAmsrGEFmgWx0LcVILdWU1cl2p4F
nYlPF26WZEeSzBUtqJL8mMpxLp4cIRkRcW0jmxdBqFqpNj1v5BVUrBzzkbrX
Hc5eRwvcdEPiJhsHtZyxm9BMIpgtX9mKYMkk4I8kpHDIv2TgQ4ioH6zSJd+D
27MQb1NLjcpudDFo6Q0CXMOJNPqsukrZK6TLE04Djq5MEi5DYD0TGJj6f1g4
sXKcIdVF2SwThv2DsnZGXq4uusnLYpTyUC/Cq9/vRHWUePW7I/lzOF/WR/w6
w481ihZoadHgNqLLhQ0uXtlvywE6meHfvzb8TLjFsJRLzSw3tIGVmgCVV5WC
5cH6MnB+Bq3fPp1VhesCYunIwH5rEI+smwDGjuDjyx68QGNKcPgg4SB0j74A
RXX3zWzAmfaq37feQuxrWpdMxbKiCZHMLgeoNoZmVc2NmZWhuBayod1wCMxM
5ibDuqjzxP7PQRQPuYtRTv3r+Pfa9BUoDx5xC8EO/rvnkaq+JRzrL9dhPe5/
LaK6oXKLZ0ctZIXcbQllKc5YuclOKUxFlkeWSDp0XfhEBqpM7Nm0NbtKVRmD
fdVMmaZcXjxbJ7am2tI6PfqToIMUPuD2JPgXPDab17mjejjSDFdInTBPK5jW
DGZ2bdmGl38bbztf8mrCF/Pw1DW+O0aEDVsrEivk0JXDamKKMJ+aRlOa1CFx
2o2Dhh1A4+2eoLNtfeEXHCit7cQ63dEU5Pul6WltmGf4mfPp32+R7RP/4RnQ
jIvyaaA6L0aRFFuTGkZ6PaBXcfHJDYr+F51r+OK+0hMBgRueNh0bCRYuLN46
BeVVoKIouP0/v8h5/WB5hgzAbnt0lVDdy5A2AyjGsD/jX8O2htLC4JWlrrKN
CKnOXyCVNQI2QVv4AXeC5FeNmicxTkrmLx3TfUawg5iGHhAmWKtYOLfnRqDJ
gfeLAauFWK5BY1f4fojfeRoo34Z8Z7NYOqVBrHQjDT/lPorNjxzrhCxPGH5/
dXhDB9SUHZ2Gn5TuV9pTlGkWBOuClzJoeG3UzjnvufS5uBCiwI/I3Iqj3++6
iMpw4d/CfWGfwX4Ale1zd38/kEalp8fM2erwJdCOcN3imE1lPqd0wjaavUj9
NhKgtSUCM+34/7cjFJsO6h0hbFgo4Ksrj6T2UhryUuepqEb+ovlJKL2sQViz
YHFxU9YZOf0KJGCiLOhREK5dsM9nDbxAI2tYuy/uqiqcijqLwbkt84LrFbi+
FWIXT8BDkRR2R6BVGmIR5WfhWgEVBWAAPP0Mlagul5JPxnGPmky2eLlx9P7H
7poeS///Hhz2k3Xvt9YyPnGe0ApUZohBn9igXeTX04F/L0qqmmy0MHtPLmp+
IL9tNYMat+04PsYIVxqwqcY3IKR5V5Mg2yk2BbMd+7Y37NuWnZoRBvGMiOzH
p4nSohu2zeCqxJSslA+QMzKi8B1cqUNusxZM7T7f5jAoe0TD/M5oxcO7sY/6
tbREE0+OgpNRV8YMpW1RGypED94paVjEZNSRxLwMvp0Pjf8KiG7ImLCcwDlj
ACtZgYHOKRoSGZ/JH3rq9nnDtN0zHqoAqmfF1GMPE5yxmaZIMVFQKAU7s/GS
avZGxFEzZTUv9D1JiruDW8jl2PfkhIq+1S7O9ytQCmhEwgS7jj8BOFQCZHPQ
W8CbPdMo1cohRGjsl6IXso+EQ3pzBOAV/7Wq7fuLdExhDgOrQq3VncRQPteN
Fm87qhY99WTPXCjhwEBKvOnldUyKDOd3i7v0Pb/YuhdDG/yvqv+o9TTacPvA
UzXxnixIRtxu6j8KWEPRm9BuKbBrWMAAfG9QnNYLoQ1L2PKmIoAgA05QiNub
cZGtn4L3FLSUj9bF4SOiCKtfNUurY+C6op4Po2V2bfc1TXL/j/zZUueWcdk5
tIPDwL4Fz0hTAXj9SwZf8LM4TS8gGOoIzhglmGwj3jleUmVrUg22HdWMjVqd
uG3QIbQtkfG0eIfQ/AARgZ4b22vMx3qsmj9XbAE7AqxbZK/oGuiFki8hICdj
KJCrf0WiQXmDG3pFBEIFryd+qA2e8UsHIyap14B1F7V4cchQzPJ6yz7VszdY
4TeXRPOdL1stApTCBpg6cjulzekQ5vaUUomsxVCLp7dUfIJ0ghqh9d4c4mG+
FRTACp8AS9tFLlw9AyRA3NUdVKcDnxRbw7+usi4/sTh4gxEtkA03okhX0/jC
67xBCVchuFnjrnC4glsVWJk7O/4ogfYDLVVthTqFnTTxzO4CDFCNnQytcTnm
tXDjsQCREhS6jo0N6NqqeH6/GmkP8wyvqd8HRHrlPh4w8wZkGKrAgwGnqK+x
HRyAIowReHlYa20960oE6zjYsmizNKpicTWG0tvZOh9d47GFYTM8klhPko9E
xTpT2cylymoodNDaDXUq+eBT2sr8R6bTV2uy/rtf+AXfNLWncZyezwqoWwxq
D36m/d/vTRYTJOM3Rqu+ED6LDuBgSB5djAGvmGSkr4mjsB6IZu2senJsB0OZ
6YgTFFRyeJ0BzgSEOwMCQ80G88iGPfCSn81RVf7f3mITOttk20KtarzDfEja
p14HspC+ELzYUmFPsJrrBo61dQNANctjeEYcIPd9CpHxw60okIT0jtBkoYSg
WUY/G6vD9FDRL6WyGDoYHMUV6pJ7XbRJmYmA7Hj80unvcn18NgvtbExQJvWq
NSNIUhQgYUo1+2ihhecGMmiCNFcvltExG3shyicRchka3XRP5V1pvCgrfHkN
y4xSIMV6CDPK3f8apjKnpdiMWUgHTfK3BAs8sjdNSyEW83kqn3No7XZ6xshk
4FO0NUaJUl0s6IN1qyHrBliwxp6YVuYjDV5J7WsxqlD8AvC3MF+wL5CKi2gF
iTwpawpyWVn1Tb+gLtASmar/uV2JmRdnrg1pR9YNDubbEEEuQxweXmZClytm
ot0YGKgySOF9JfKjTYojnM5b0hC6RqnGCvGlmlriFxP0N05yall5El/cNdFk
xeL5mT+c6qO7ySaJtPDQlwu5XIULeADe7PGcYhkP4Sxh/gEzkESLWraYoWCy
Jd5NC58LB2wNtZcT+5ggqS4GbpOaj02RgnV3F36C3kcb7/tOkESBDSs7faNH
uFevgiBYYrGhvrF5zRalZbKOBM4kyU7wmuoG7qLFLuwpccucy71U4UqYdYzm
dAPy7mCJmUksHc5NKnxrXfs5vHOrWmOKJsG5k1PBsgRkKGDGqHHoRA2VMWs0
Dz50HP+pZKApdBxP1ywV1BMYmp4yhTQ8LuREUR/vwHf19dOf+pzDfq0P3Mfr
x9xvzriGu/B3Nre4np2Io3lhXFP/mRvwNY9zr/ymFTTOLKGt1CQR6dpqs1ks
+BNhRVnsA+PojuW6VmQEd+UWDO3xUck2azLJSbEHRgk0OQihy2o86zyrdtZa
zXSVsFpu4onv/DffqtAGbDQnyLd7oUWIiuadCVCDXXjihRCUEdNsZG3WMgOk
RPw76tnRQNhU3Km+uWqgjJVx3dRqurbnSd3Dge0U7z6GDffKm15lTZiLsN7l
vqP1xSGtvI6QcE4wmB96ByEMJvLcQB9pPV3x65YZyAsrYMzpeQXrIdNBhrSI
Iez6qdUIGJEZ/JNuveMMc262zs55Jkkzg5W4xJrmRBxv50b/ibY6qe+6TtRK
N+6L/zCcQmNk5j9u1hZ31EOmdqYMwxIq8P1Jic9h+Gef96y/IaF9cwlx5UrU
Zq6gXJm2KLcGvlKQqqIlwM1tm5WALc9R4D2FH2aqORHPBm9JAzoBYCCGd1UX
BZkHjAooB/OooboVqrfIRH4gSOjMzGM0Jp7DSvAI7br+5qi2KT+CscEwKX//
/OLjlQaj5mHS2CHLmurZcZ6mTagTae1Tek875K21/6UA9Lu2zIIXsonWsmR2
TXHj1Ov6+rOhZAdtWUO2h/M6tDFCddMBsnd/QdKWw/HsnEi+BmHUQiinL0Uz
U6BTDWuK+dblUMG6d3SNPWRHMpVZwUctnDuT5LveKU4rzvGKRUoVKijQQR8A
95vHMYpZiO+jI2iERDjaLvJHGqnrfJ+d7+zDQd29UnYnM4vO239KLjtVZVXR
EMMtCvFDrjO7LqG53A/aa0TqGTcEEoHUW7VXPb5m6MidRVBur7/RZnJWs1zG
4ejK3Cl1fqbhZtHYf5H2yigtBd0gc3nbphR5Dnfp3VLhBY6Nx9OBg7zY/4ar
TM3NEoruRSm9aQ3mzF4b1+HGuw/7iFbITyyB8IZ9E9Mx+92soV0fMt+Vnr1i
AS0x6fNoZYdtyhYGi3TyIVpl0bJ9S0Rw5nutxtLa0du3NU3o8QbNJCPwXv20
NQoKAFKY7M8d3PsXvN7A9Rrt8cWfwV5I2l0j+vSIW8lb4JN0Je8EUkR0DuMh
Eo6YTNUf1I1VwhgK94mkoA3hV6nuRFLdq2ypd7FKMVD3YGpSSKJzyPlmdFTm
XDEeyrl20cDy1koT3zEd6Yi1Cf4Tag9D1sFH/tZavAWjeKzH4mqa80MA+ARb
WM9My90a+Wlp5rzn36BlHiHO3nuR6+ijq6x8IqRySLNGIJXAbHhBVFnZ10hr
UPCrF4pPc7iFe/YRY2aTQgTztsey5QVt6CgL4ukj3xzRzXOaJ/JurDgqaeLx
ArKRtyNEUz3wKw+LrSyLylukOB9fbwUaOIOTtw1Ri+sb28H+FLqNkhwaJ3lz
l6P7SplO0UdEBW51ZMxmaDZUy8bpRHNqmp5E9qMsGpUE3CuWfnQ0WfsAKsK5
bJKk1z6RfRPgxCNudx739CCAzVTyp5UddGwNVB72o6ydX51Jz93nIuADBdcm
Gflaqaef0Dw13RB1Lkc+5d/E761kv/iledcSpgoXkuLoEzyt/EBvkCADiR3B
vJN70w4HHbavX00nBHWfI62o+lEANbzLV9O4ZGMtRz8urrf6XhELjo1MedP+
bmDralc8xS6YtBg0roxWWvuLCFOIVH2wxWzu7tjUo0hKTFzzuJoRsw2CbsNq
e3dFq+q6mE2EAtWMzYNVZodm6nourJImWREc1kASt22e35CffCOG0hVuVYOp
/gTrunRKYHYPI+MzVEjczTQqQSJmKLWB7+umZggGV2MaD8Vfwe1W1xWRmQLz
iMEz5mQdGcAI4MvS81nFhMM+UScwB6MZ9ii/ewRjJTm37VItnojN2mpbFrBa
8BKJBfKvsa0gPul3q5MnjBmHU1RivmgkNpb0OzSjix00V7oOEtZFRQ/3Un8m
ONPz6bPtZTwihwUweYXOHtfneGoJAIIgYdGui09kc5cKurUTVt2qrzH0UDn2
kLDJZPMzaCNIyYtQfSb+yup2tPoXaWdL7oPTuDnwlF8XN0b2biUYS6R/60xA
eUzJJfXknDIFwdk420OhSVEMj4d0R1c+Yr7VThCZNO7sAU5P2hZ15q0oydSL
gVo5rPudgsi9CgXPM/eRpp7wehTnAlMCG0iHkCamjD7fpP2jNAeDGQUGL4Rj
nAI7tZL8jkB0X7oLlAcHg1eF89WAeFLW6DvXKeKDeJDbZnf+bx3wpUHdeN7h
9Juhl1f0irFLKB1h5OYd3bz3mE93oyCROYkqOS5fsPNhu26j80f/EYC2Ryu+
Vqd7emlzX1Dm+TTdfqxXBWtXgy6wC1xVGEG7rnoGds9X0sdPkwwCsfvV8KN/
dHtsOvY3XZMB4fCuUzwyrLIKEVPIpjnPH5i3TyGtrk96QwxhXJu+6hvTqA73
FAbT/vDAjE7LNn7+eaPh6rmYTIeloTuoNnTD1zExawsMcDO1TNzZtObQmIYV
bCY0IN9ciujq7lCA5BEiurJ24iIiE+aYRYwR9SOErFebEcrI9Q3obBE45Hnz
ABWIfcrmNf4ngZCZwsgvKZDFBOpZP++9S6aJuUhDY+m3PtfD0sqXp5rnWA2/
OutB2Vz5CR+nYDY/dTJIn7r3WQUNO4qhVgbigEgXSbiBdDgZShsfOU493xkm
yJyybWuUzb9J2dcaOTuznCn4dXEV9Ppajcv7clBWOj0gA2gRDbwH0GDtnKay
KYTpPCaSBi01tAWJz8PHY4xHRIb10jD3VqcaHO9ckhvrWjHnpeudTdsvZ3aO
x5hdg37x04Kzozpp8nWdhF0vlun9/XmBRfLgxH6B48ALxadqO4ElDHMfir0n
KoZxU8iKMS1LmhPmgbEU+84wIzrKI6VLqBIBnjesezcxQSqboMG2nDQCmCdG
BSvSPC+g00c75by6THXXFRfOKucaBWzfneaQx1XiNhtmfM0Xu23MpViJnNDy
MoF8sJFrtT4WhNymvJmUhcWB6CnKuX6TO07rQ99IwNfq8CukLJwvIkMPp4b6
OSYGXglXaKy3FnFpWeo9F12H3zovomfDF3ktUGfA+YvA91ltpkk2FebrrJ9v
H1e1LRMjaqL4XS3dOexDc4mmkVW97vQEhOVCiftQN11QozOjgbw6f5AzgcHA
OAm8JoFDGTeU4iWQSUdXnC5ECgyhK37+BKKvXloAnawYVDPvgqiqrDPAPhbj
L/5swL+PjPM0B+O6ON2rL9kLuE2dCPPGmZg64p5x0WufKTDouGw1FDvDScEf
ywk89fOLNQXNewxnu/fBglcHx4dAbRiCM+BKMDaBiB4nx2NbzEq2EXpYgHOd
kHG9nIEUvz5+1KKTSmg52/BHjNVX9Bh3ht3zDEV5LNCV1vFQuWT3NgIeFxMZ
IJdLg/mE6YF3R5RFgUIzmw9umPYmW8X+tUvgxht37EAW+esXLzNZhGHnjZc6
EOgmUnrGCbf3D6uZZPoIV4dg1NQMaR//PtUSODCmdivnLI9SzlIYIhSEQj6O
3qEbzWZyGvDcuKYuXOzYfvFWSUTVLTVH2uxK0DzTXhNkeRobUqzk2Xg7/8g7
NrdFDssC66vc5mOAvBdBPnD2BQSnIEpjsd9wgJ4azkp3fG/3SiBGV6eai7+K
lefjAD5tbXM9mL7lasE+XPFD44TayPXW5WappoZ4f+rKubSfS00a6PeL9gLY
3/NQlS1UgyBmi8wLU+4eVxisHIJ7IJebMxgIeYJkoa2mGmmgtk8ud5w3hLvV
nbhIwtA8fmUSHi7CnRt5Rk7VVXBRccHgOaTzrwk2le2gyNCqWlkne59vLfPb
wEgAF6lpurX9G8sq006YjwEtGJJkoTE3GgenM9kHgD/8alvohc7Io6+Odb9r
suVR27E3Zu/P3XWVP93TGG54QBpcPbgDaHEh3hVkeeaMv9fjhB8QGLeTZApl
CV3ynSzthlIxLzbxIDLN++MPwm7BXN9nq44W4jmjwwvJ5+vTE7e3TXUcu05i
6VuhDWAlEy/0V4vX6ECrB2nBTjYdbx+8zGRz725cLeUHlzB3N64qcYNy8Iqv
r1H9HzxNgrC6mkKh/tWAzVOOgiRslyPeeK1RJu3sAOYTB8Vjmc94JKXmxc+J
KdbCEVFBRAivCp1kP0JOHinP+NT9a6zJN2WgIWp5iaAWt53aSmaJ8qfYbdN5
oRfWxYI7iUTmr+yyFae7gRTOzXVw76iq/p/vJ7SQWq5lXnR4h8I5+cZTIRoT
ju8BrYW6K9oi09o6Isbn8yTD/0qegWu6GM72NQqOmjJ9p6V5uUAT/lVAcGYW
RamPvb33OBPW7ioxBSh08YDi7ZgFl6IrBC4GQdUnu3QhcuBNO8c6Mxr6KiIJ
Kqf/6rV5/U4Cfq3aMHPAziSnXJ1H16s5ZyEz6OGOzSxwvmY07rAqjYZQISm/
plt/qhR7y2j+czO72KUio4iooyQY9D1o7DcU59wFq8FHWHyxZxlQ/qplHvNP
0vS54sLva8R5RdbWqXIeQqpJ632nkH2qnR0cenNYwUINCpfbfiwPBzv91CEt
oJAhUhrw1K0AzQ5HH9sJfDHCsONxiXA5g2dqfNyIWCeQ3dsdNOxyGMh+R+6/
5Bnpn2chyv2HV178XizoKKnJYhPKvt4JanHrxQEEhpcHl27QmMn0jsjDTuXA
U6vsf82iIuOWSnfvRAWHiM0i1fRo/RBWFITjtiFDMkP2QzjbhMJpr7mh5OR4
ALS2laIN2FqjvDNPkSOdG4do14bgdJVcE4xr73nz0ogcvwgK5BulvtN3odMk
d4aS1kg24eE0dLtOBddP3pu/i0EWyfbki8fl7KDP4cQN70zH1po7EF9Berbz
DE5CDCEY1unpmfvICaI8lJJ1bItDX9pe3SAbTjtE1m68yLdGvjBEddFku2kV
Fm/DAJxem3f17NFc8A+Xn6Sem1O0x7Eb/fm4weLwEzXBFh5SUD4bWGkPYPpU
Zbb32F1P7xNqcRFXa1VFinRCJDbTJMDcuo3+6Ti//nvUYBeNoOT03q7e8gt0
8wB76yJh51vPERTh5EG/zvL8IclYQz8xrA85QRR8tEkfAdEKOwAs/rhJ9sdm
Knqzd3B8Cz3SBG7x7IwABXtWqacmlQrko7qjR4dcBJALqeI849iw/6jfVNhB
5brWFeVNAIGtwwMW2qhzdJbIwqeEOKjfX+cm39Dsn8PQE9cQSaZGmk8il9DE
tZch7mxThq4CrYcBdZqfQERze4CGwoTuRzTRpvY76t8n/DtyfFJi4TS2WD6b
uxnc7Nch+JHz5K5adKV4Cij7ci59imcClMUQcchv9raiXoQcpTEruRGilZd4
g7lAAuks+6ezQYzL3Bz18oj3MZ0Pfeo+oNyep6uzNH7H5K9YYK7gwCwvfDrE
Cvtr6BAoi54dDKocP0/W6XeKbAjOiGEKXGrLylJxEfWFlbeF4FUUMlgQfc8P
0dw5awwVSDSAsbqbCNDCbiOOXAZNaFlsWYI4q3lyOAHtKg7ddz8V4iRvRcep
0xLXD71ZnQOBEfA7sQNn5wK92/n3dY+XbS5h+w5+7VIxBcDoOhH+aJfZwtQk
vKF92yRwMEjjNYpRBakq4CBIy8nluKvSi6uUcvZRFeLxl4tkwfLX6cGGSvE4
Raz7PHOyLZ4JgyNu0bkpQcptB92nlcM1smGe30dYf4r9FlqrTeZLpw5LpPld
JFXN4syg95XusW6OOzq14muh/0QdHea3WdptNIdntIin1J+PUs8M4MoHdkXU
wjuAgUEIQ+JrhUKZgK8BU0G4oi57mVcPmDCwRfoDF9UwVt+2eu5Q/gPqdd2Q
In/I3nwfUCMDc9g2pnhnnLvRhm6EDyh5SMnsvVk3OSXK4u+FS+4HGUDzROIy
/ag+5r58cnwK6bSmmCOFKxEfuQ9/o4nYAeKN8F1X8vUO07Qstnsb3/jHvcNr
dC4iZJsszCzfgEtT09HpZ3QgDo6tNClCzX+AKNW87K52QReGm7/AJDk9nT4P
g6pZ2wrw3yiZnTa8Nd8zAqyD93b0IE12UJT0hi/kza0G+KFskK/0lpJ2dQQ+
PGgO77I3J3ekmjg2DFG/mRh8B6wM1WLkNK+0vG6pWCDuOvi0J7fbBSN5UxQf
IjDq1btZ04DCB7C3+/JBi4tlMrrdhGXq2SnxBt7/feQgBIFjgm5ne6oPyZux
KMs5q0SWLBk3i33Ye5FGvFkkbbyC+zZCcR1BIOZ4M9piHNojgsmsx6oJxOkq
wx7P7O1u+aqJElzJCOSOjw+s0M4WFWFR3qjD4Xh+WJ34DAHxn13+GLQqZ8P6
B15o+I7RnhxRpQQCjtKkrtlxK/oRc1vIIj8dO4ZUGmSbR3/Sf8BrUOMIj/Ou
mA/Th0nGQChTiKsnFAA53rYlOG8PxvaDoh88fLopaYnAslUntYy+Ac7TdWOM
1AwvsNZwShkowPdL11oC+lE3ZP4+T6EF22wJ0JO3pfPs2grPevqRjBr7d4yr
8XR5ibr1wrNKBqwzz9vp00SmTP5KxQejrq+wDS4YmM/CAcT/dY/JhrfMfQ25
ux2dgks0euNHRt5BG5cYW25maaoaRd1oV+P0Q6Mu8JTnLSNzTZuhNewneZlj
OC2tsNSTUpfez1lGgQBfIeGIFXOqZ/ZLV9Qc+On/vfxREyQFFcPQFFOt7peO
ckQuZV2H0CPqK9pZK9if8i1apf5ZjJ6p2HSpmwP2MlAJyfiW831zY6CxgUZO
eNgn/bzcg+sRISdh5NxXlKUppdPowwuRtbZPSc+FlHi+eNPyZUR0vSAjcbNy
swkqLhwyTnGFaM3mZ9BaviqGTWfGCKFCuP2k1c2XjmSZUygmqvXHb7U5qI6M
ZiDdjb+4yPFeconIj0Uxuv3E0qlZjZkhQWj2iY41gq3ThgLLpXFI2c1/Jy7l
cUx1wN9FTX08XHN9yau8lTfZwmhJCadP++sQPemVsIkS4YgiikA5JUjXLQ7z
nQmtji8PAxOCEhzEWBQzexZCwJuzs9XM+81YdxtR5wtj0L52b0aqZ1ButP/g
mySwgOUIndCFcpBVEK0vSLSfqf+7YQ39p6vNbZH9+kCxTl4u0xJZfddpwFjF
s2JGA2EXHD0pYzPJwyY4EMVHeYPshH/6xJZgyweGxMYOrNOeQdPU3HTQJ2N/
yqi5tgvIW2gBJtvtkbT4VE+V17Rl0CZCrbWJ72m+Gn8j4nK5tj/BRn5Y+DmH
RUk4v/Nev1ZF7ioQzFsgy4aP2eMhjHAzvVo5sowwVX5qasCRyMky5RtSVEOy
GgCIehSRoG/B0NwoxogP1m9mCCs2Q0p7wAZk1EP4VxQbcnjsMvENJNhZ8cT3
3M3CUOmGCiV4agxa33PMPJlPoc5UCOZ0k0tACc2BbdycgSdf8pv7ZGQohBwQ
yn/x6Rk9ESvQWnPHJmV4UDC3+d5F+JJfpIfyvWVDTCqPOhbjWKyEWXndjCV7
QM1oRxJMUw1QB9SSkelloy3ewmy4mI94BZ4UYCb92wTQ0Lpj9oyJ2ruJmnl0
DrpwHlxJUAsoM0Ybzn2cnEO60Y5VGqNa2j/Q2OW2dbGVVKmb1YQf6pd4NU4W
oDkQdHFovpLPKjvG0q+lt6XoJeZ9/ijN9PXgRhRFSKNBMVpJrsJ5pHi2yVji
iro2oEeqVfrHrxjt/zWHvvZ2F38QaowXdtSE5Y7q2Azud24WHmJ8Dk6eU9CN
pZ2LqLJL+DkfGrxne5SdOVGrebjL2UGgu79vlHiZOjovm5pkN9M1F5LSPw1h
0fQ+vO2qt4PkQOPWpbTLQQpk7d2oL4IYgq+ekb0+CFqWwRkUbUEB7V3yk7b5
usoOOtnxUEhhrG0zH2oqzgcJmnZPiVt0MIkbWohkaSN5RmkKZBdr/Ut6+yvY
nnpJ4DFKjXC31oTggl/4KngN/GsC6CcdMPRDS6GrhQm3IxarKHavsMgkdrh5
QeJgBaGOSE4euDgO3WiglI6CaVnQSeJ0ZgyajZii3I9JJ4cLkID8NRwXta+a
YjFG4dW4tez0ZO/9Fj4SPMxK7ARuR9yTaQc6Np3qQu/nL2PuxmckygJFStJO
ByuNWSppp74chzEHbNV098lms+/sEW2oMUSzK8b486JFlL+/qH4QmxIlss4e
ptJUBXJePX/1J6Zg7QUeTO5CdPalwr6UA2bnQhyc25OH+Cz5iig3O24mNyqB
n7nSPq3uZojp3vmo+Kruu63PWPPZMhFyLKFBQnchQRb+k5o71KB2ZDghtIdA
kyC+wHTdJzuW5jJ6mgNh+HHqsaDXTVW5i0bDPSQFdQbIP6GS2Yx6K+btcNiR
pMlHb8GcaphsZv4gnM4N4pXXf7Wyp0J03ljVnm0hBMX33nw999JfUOIS/rtn
GQbk+jga5PI/mKqtfDIkj6h6om+Y6+vycwntj0yeh2Un7rn0g1Ytbb2bX10L
W0M9IBtyDm3xuxGqUJ1+VIt4K4SkWvZvm6N+U/h6AZil64JulCDkAbdo31Nu
GLdIAGcOQFTgwsy9yNGGW1oajO2tCGQwyVGqbqTx4Ltvz6e7Q2sWIEzOep/O
fpEV5Xh3HuE0rYcnAvqAyC3+52GPLfAqtpb0LpioSsh+6eiUprDSnW976QDL
aihQVWP5iHZ4D4VqYW8S8qKYw/FZn3VzqCxZulP4Q4LTDw9LsQN/aAQoQZOn
DmzPglwwoHedVYKrYLDZY05PxTVtVwUY9fMhx1JqVhsiC1TAIlsrKVaBle01
KKl8lehfEpzbg5TBiNRIztQxssPKklJocj5fMhxe9yZZeiyQEDip6y2aCx7H
8IC00Q/WEWcIwNlqCB8gRRV+S7bkG+jqa26MfFUe1IPPAr9CyGDXHM8SYRmM
u4Nb4OwpvwGqjC2/evrgRnUokniazT/gNYDeBZNLTDD+3n7ObWMF1QX2fiK8
t4BXIThgfVoeDwdNMx/AHZ8FZ75ywhYrO06wK6n78buVQtaZa4h6NZhoz8YH
MKOm016uMrhirVu+vtCN02T4Ti3J/wnYg0fiB851FSVkGjGvyc42/ccZ2pct
FtGmD3sKzqtv4ZxzXDIogCY5wRe1T+SonrIHNgnBCroZ1ZevSyyf33964q5A
Pn833hwGxR7pDxu0u7e6Q8xVCF5SNn1tst0yWv1sf94YargikDwAOXwg3+R0
Mp8fYMCraRw8hjogy15aMNtnrdxTYpmC7OODJdg8b3fQDiOu3zX7VE/iYCOw
66rXs7w8N2vrK9AfvfdDlR7hWH4OTH2DtEXdmYqMM7Ao9/Smy+e6cDArneoC
7n93cwjnkib/lBLW9GNBM1JfO/xQaUyI32QqQ1tIWyv+9rjRzAXxCqM+0D3O
M9PuJQwYVuaYa4AAwsXLBSrDWj8k5rT73Nzq67G8u+CoBoKD/Xs3B4izwAfS
O6eauT3DZOriTS4rG4i9wuGswiLP9Rwk0FGi9FJRYhizxfXmfYyJ+diJ8lVh
ciy6FlbgFhGXmHZibIhjxggiQco04cGSZa90ApVP75zcca2SGfqM/bcDCSRR
CFGUQSjnu8qAXxP5+aaXPyETc44utncu0AnE7AIuYQsSESVYlTZ86j8B3Ufn
xhsUUBwpxeNVKPh/Sf8+vICHvWfmLy/Qq1wOvr6uSicj06C5NKha/XTTAbbp
zJUGp3BZkNaO7iPVsvCO+gAeITuNferpyZJ0psAQy6wxLIQHUEfHNNVm2RMZ
ADLrh563y0HJ0GxZbJDnL9ev7dgmo15iVi7i9thxm82ZnQl8vlIt9JK+kfYq
QYM3hP4JhT9xJaEF42Rr2liLKv012exOCa6Ng2/ZvacRRkh3yuIqpStsRV7g
QjSZ7h4RkSRq7SdfswMNVve+xxh+zU1c1Plk3Z2WTVpDlbhHEUVUYXQ2CKS7
tfrTDhCwB0ORizO9CCwij8izev/gl+Dq5mabx2pa3i4X15EKVZVEVnSvBmgh
9bvUJHXpI9Deur4IkFmo1NqaBwLGKndTd+Dvns7QHO1HeSXyZ8RQgsSaz4vl
Rj6ghR8Ze0mFQXPB+vbnzrxPlCYzpV/QqZx9g+rdbbovIsvJB7v1+PsSOysa
IuUzJUwiO/RC5I6bqwwrgZhOdm6hY68vxcN2RXPPN8+D4c0TYkLddGfKrThH
FqB4k1fgeJB1JlwSKKtXSQDdyWPuZq5gviCgwXj++Vv2c3jrxhRAOOsmsb4A
MS/uNbb04OEzfwlULXnYIl/YlXloPNlv9+DErh2Jj9UBBtX69NNUzWK9mFN8
6SNw7TVDbIc/xa8r6MC7jEK56oPfREr5SuhAgbC+bgBvbo84JfvuxyU3fYDE
Kcyg2hF/3bMNxmR/z2OAcyiG38yUL0Zd5E99/EayfnhxQIyXVuhLdMC3R1xm
HMFdUkd7ZvHCr5FtxL+86DZhnHYCBM+Z3GICS82/m2BJgFzyFd84uKNufBad
T598NAp8jfjSPBMGJ5+A8Txu4x0cVgKFtMp3gUCx6RXLwPn43bSU9NuTZlfT
M383tS4CCEKddU4jmjn8I3xaGxm1zdywrmqOLXViQ9oRKUci3a6mO5y2H/BL
ixqMGJLP050A2pt4wiRjh2lm4TLSdWZjGRZMYFVfzEO+6WcgfNU/a0qS6VAv
hMWuhhRqqsI2oydR9pl2/3fs+138/gapDzVZddD3Cn5umAuCwiBkC8ljRcIl
LjXGGhJ1rQ/DaFKiGIvuJiEcnnTzFa2Ecu/N+Abw4h76XimMVuWcfkqCgu8y
vKIVgkQ1f5kSG7qtND2BgJg3HI/hE5QINxCrOiS8LZU6E9IbsrQrEFN9g3wR
yWJP/hjsNzYzj5KCwWIBWA57X8XHPKPtCZ8IiICIxCeGmgb7RRLvwBUIBami
xFNFijc8kReqKoVL2fHwUcYauo9f7uws6EW+c63l+QBSPrWuwnENBowsUZn5
442hPxrKe3T7qhX4Vcvuq9bYzaPqC04c8ZkSh7dHkYVqpR/3QwPagvGnDwCJ
n9Gw/7jT0rrrXgtGax7EcZrXqi3VXi3o9B0mgta8kAsqS0vem4KQXGsyGJ4y
PMgspPE9fwZBdlN4LiD6oUh908oy1ONsv897lS/lSnzKfuW+KyQMBNMkBJsk
7YIZ/6icK2curka/9K0QZ6DJrpgj2MZMWxOKMj5XQ+AP6umbl2a77rIo/zAF
nPfz9Sbhfb7e/3yj/P9xfQTgPS/KQ4Tljbco8botLqW/aIgJ3MrHko4XVXxD
sxzuRF4esQ0Qer0s35nZJ/iRV6AIQs+MWNyxZOgwUHss/OJudBckqp/40ROZ
zfVVLj6zt1CFSAdWjrhGZTXwGYpDwKcHfTH+B27dHQ+sk8mVRGfIBUsuzUZI
WcnVEkA3iEV001TkPYMcSSTTO3QlOzc5sVJUK+8KctWka3Zv6Dk3cY+sAb4Y
LpSovtsmAqeLu+ZvEZWVpRooqRw97CbKYTeSoflp0DGfhv3da2rajZ59nTmG
DnsMa2QUlzBeGqRP1hT0HNYLj4JuSNW08DRI6uqM5yZFUIZa4+MyhJN3nJ9j
l2qofiODB7V1C0USuYRpdnbIcMPrYHjUie9G2IRcrKwljo+m+qFuHDpKppQg
wUVxg0O8KahZ6T19LJH1g8Rma1PhzBB2uUT348S7F+kZmzbyfCVyvd0eSsVV
K9YLVvvCkWiRsXoEBBe675+cVfbhxQDN/QB4YAnesUa6+/qUbz7WI2Xs8qJJ
0OdQEypt1juo/nun6ioCtYbbHVu4sxi1j2IsBaB3NQR0x52RIbE+ieXP/TQJ
kZ/XbafLx8Mc18/1KQQC0qK2+sMIFnCI2NxF1Gy5iWWrlSM3PfxkE3hbdwr/
emLfM0OY9NrMhAcQeuIjDoniRGSo0gbnFf8uFD3//WTFZq+1JQuXoKki5Weu
QnGB0rhKe7EY4Kv9hXicmvqArlHzfTpYSZq5x40/wFfi2KS7V2JwO3QvQjTK
slUc2V7SxgrBRlnZSQOYhso9fhoQ7xojE/6cPyv5AZO2V76nnT3vw4soe6d/
DGbwLw71NYgp0oeX8r8icQ8qI1Y+QdRwq7/vnQkj1dmBeSHIyR8INhHen4ql
EuX67iEb5R7WJO9xTzDNTBGDvvYF1RFmdOMBn85acLVia/elXddPfrDlJ1zS
jh7jcO4Opxv19/dN/5Ie2dd5C4ucMkHgAKM2XcMG+kqwkT9GNUU17D9vXTDv
TxqCskpdhb3QFsycvKjfR7d5VmY0hHDkr+vtbHQVMIYMrSzHuX9cbE0Y9sJf
qMybmS3pe3ZFP/Ywc0fuZYHyOuzEXXm+jri5lt/kxM9OIZpGdFdOS7mOSr2z
pyEAnmqFd20uniH4bq/kBd9PAWc7YDuGVomq+6gbBRPkSogPYagWvvUtcGKr
L7gRwhsq2y/1CMFryoRDnmbb5jEDHJ7ypDwf9t8rRkTeRCezlPt+UIE6WDD4
3YE+4S0LmVSA/VoAjJKbybRbwOmC3VEG4kB9ZGEGULizNNAxqyCt10cdJdKj
23RHh0/HrknlBM2EQCuQxXk75LHyk3Hz2fcZG7jSxLnou2P63R2tY1VRA3wZ
gIHbuwONXyBvQVY4SvYNdrdpJQYvxAq0agXTS+2R6UyytOJK8AlmBsMV8267
/F392ygbBXNrDhu4FeAgZFffallwlGH5qdK3pCeorm/OCjVgEYiUqIFq4HSQ
H9B/1fPKq5jy6INt0EPyl3mrQXlaV7PFychJzzshgC+skk0QydU150D7S7cw
Y0HMrgzkGP78UzSOGkBhLKwhtIwTVZ4mtiprn5KHo4xKR72aJ5U95Avm3UVb
WsfUlaMJR2ztXyOXHeg9s1A/+FGnsw4mkoXD89zrexDNV0HosJFutYdqjX+s
0+e/LJIOiKiJk67a9fCJIQMTA7fcFz8y+jkVh9sHKK0iMSuukeUhDscJ2Zxz
Hp3lmgWWSK2mFtuxtKuD66XXZ8//7yfpQgVGkqmKFydjE9uu3P6qYKj7Sqyk
EvV7gmC8VS5yhGk2nhi/kwUu7Rv7pU8BroqnXCBTVgXFS+POmO+qr46RAZES
CdtZ0TOsflpnYtEsLruObKfHts04R7m5x7vVQPqcXFis0TXJ3DTxurSjYYL4
/SJyn/ZkVYBK0YUgtrHJjT34equMDqycfldSwUD7iRxHAC3VS1kx/Td815za
+9lDAb0Y0Szm5UQASKmZsMBlVDvy1/4gxrv+wQ4WyCSLvuupcIGHRefVI2cp
+6+GkKpqXL/DimCW1AQ6lvWDwv68grJjX2PZDWcKSh09rL5BuF4xHHq+aKTA
3LcjAEuxZ/5qsT6xvRSpWxy5lvlA+oRyQMavnYeP/fTGD30aSCIOPCvW+PxE
HobumuJ8NYNDMc4MIb4krvLvORAAOQgIdt87t2WY+kyzX8OCVWOqVXJ+qMBX
ubmV85Y4cmjRm3Vq1WFh9QuXol3XKobDzKyAFv7nhfSLwp5CQShjkIFFZLg8
tHUirUa+8dhz5ebYHP3K3GjzOy3Jy0I8jxRcdEOFr6ec6aCHN2s0Sd9xYTUA
cz18wsaTuOG40dQyfghJf8KttcN9B1BxwfQ8BLhbqFQp68llcycoLfjhvKmF
VCjyi00zFLNM5HOMk3X0x6KfDahYgDcWNXP4T/+SMw8CU1ipusqecAsNJhvp
2yoaarJH8CL2TfKlpWe87tRvXB+234/RGhbqTuX6Y6W03NwIl1gFDi+4RlDT
cSFNVFawIE9GorA4XPBpbS+bQchuc2+2vMdXoM+UixaUHGn6bCHMz++MEox/
ir6SoUBu/0OOyiUjk1YnZ7Hlfa0kTaA2qqiQLk50lLSfExctX7AS42/Ta5Bx
F61ylpuMGDtc1Wi05oTljeog4fINDHtUCMsIjCwHGNvcbr10kPRUTeSOmgW7
7WR3/fvMPAbHeIuSXwph+psz/F74eedmJxL90S4/v71FlTwxvGDzLQpQvd2B
Bu1hx8wsnlDIEiOgfqLd6T57pkSqfFxmukUK31bwR0Zs4Ndx6PSBusZk4GnF
MjOp+XU+gZVff4L+7y8l8GtDBpwJtIC/oNfkVmM/iE8qNVWzy0GrAvvY/98Q
RwCOR2PO1NqU66ngZzw4PokCZ++ZSYh4F4qwnNC7Ss/GOfKs+MkW++CDAqp8
ocbtsypuTIotWn0+G0RQxwpZ53I7x186rRtMB8NRCrqtTucv27cTFYTOEp1Q
N49jTZyfDTsU818Af50T64pnrg4S8uwGl9GTvREBrji1A6ECPbc+VO3OcqGo
2U/A81AOgN/LLynOWJpVZGc6/zvtm0TvKFkYpczqhEJ7Ef73m7I4V7ti9cmS
xSkrTT0G2U8rEdl3zCeolzc5cK7oLA/Qt4T/+6yhQmnrCZCoobTcizSA0eRl
8MmWGwKXNDrNvdSDZzHZc57ERhXlCk3mF9ZwvPGbiara3diMKftsDSDPaJE2
dFTzqLVwg3X2NR4V2Fwg1uwms6lwXoPbpVN07eqUH2DZqNh9A0qnDb5PP3E6
afqCUKyFJacf2Bh6t92tmiytF/D2o3PCsr37NKdFR8fFWyCQPEUGd4ej4QuM
m37Brk24AZpGlBT3coTVa3MQeNiNLn/x//kVSbnqkeVyi+NNu3BRipkb34Tm
aPqh4XLjvoGhowW5q7/avIVB+0Um5EkMO35JWZR+EVCoxqk5PDrhsEaqIWrA
Z8Qrla5ivWJWWB7tj/6nH1rdj14dw2OzT6q290kLrFQVXxdmkL7rtJJ5kqKH
8ZhfQi0kfcYfxANCoigQaU2Ub8u0oJXtOl8e8OP2RCyrlw+HrNR5Hs+ws28L
KwqbEql2s2Nc/+EwguiELyLvgGJ6vHExXlOyg7Bn5+y0wjB3724g/sjFhGNd
JO8gnKnQnChfh9LW9xUtLtneX3wMUR0Rn4L8Kh5DHDWqM9Wvn/14MkSrpq6J
BcfHm5Vbo+oPNAqQ0Vj3N1yRQfWFoUkVYRFlPC+Kq0FBJS98r+12CkNDEavg
sx8v/CCN7Y7ZNEtVnPMc3E7WSF9XS+mSKM/NkmnxB0e/qcrcEpjza+pRH8p3
youK9XrFXp2k3xXbzD775CogGGf2uCVjYXQLsrEwgsAxv+Etcyz26Sbx5DlO
f/rXdlvPuijosoDdL79mWVQaHZq/cZtJWncfTSCrIPZrCGxARtpqmayFRzzl
jvHWov6/1dKysQynXcvf7FWaaB0+XfRs4agbHtfvGaXDPkmvqFAFIQFMzMQg
G+pTHVUJy+vLJm5lpg8DPYLWidY2kqGSOZQtBdjfMcrEpFC3dcuW16cshpOs
MG48cp0OT6yz/Yvpc1532Is2tw1DVE2LaRWUOFlSxjzytfoYjz25VQOn0DMK
JAnezr9YlpfZ58YuzWV8lvLFzJQsmiVroJOdixSK4q9pnZ9gtVHlNtFps7cw
ghFyg3e/6CvjQZMZm0yCAPw/1YFwI3TD3UgY6fVzX4uPTRr56XonnZfKJdJ4
bs3Rb2sbKFyWyasPXmLS6jQA5WI/QiY7IUhLyx/G16P4Z7604ENy+AhmR6Oc
I6XPhQv6ER8xvlJOJkV7YkieGPGH5AELXKBV7pl6pYMVrGwrSst6KXKVkVir
PJkrm+15+ucPMvP58Wj2M363gDbHnZLCaacAMRA03wWntPUKnhSKYJ7jeSDR
b7PnjmfyCzGW4O1q4aAu82IYPlYfQ1odxv1Y6q52K1NEzhR+f0S9i9f1vbeJ
aBiKmTILpJ539/vaHwL64OdZ2Hap/itt/ZDKt3nOKnI+ywE3VzTTxYU7QDB9
/tzPP2iUX2CDRjd8+G87m+XNqDtAoIHejeoWWo+76Pp9YxJo4mHHD+QaoTt3
KL/W0T9FXvdGprsJ6rtNtyhfMQ46UugE4l2ZrF9wjQnDsdpfivquqvfmr+av
v02r2QU8niMpGc8DdOziWbVwNNDgx3DUDG5Rw6DEXhoSBxgfgy1iVGR9S7NN
N/c31Ut+tFOvJzKBYXWeAM+qJG3ZfVlwo0e/VBoIPUheivzygxC5lWkdJZxP
LXCTeIEIbrqJm4F0njhwzl51gwvJ1grxtrMo7nSQUqGnlNNlc4fOlkzs+Jff
V0GZ+tBAp+b9bcYXHezmQrzI4+l/BooAi1ShLATcKSjxetES89o8SR+XQJ2j
f5vwpwSDSpykQ3+rDsU08mUv3A72QyJN7ast8MTeBquiG5nC9psA2v4rNVuv
rC9GnhkeG1qNmNCZm+HAnX1HSa3iS/eFFevNTSdr7gKzFMHmMpgZWPYmRstn
nwY6OO3qRwLLBglTxTamE3mGMETPTjWrWefLv2J50MRQ5Uf250qiRPFAbxfj
baIYgY27QF19Pz1Ip9/FKnYPZWtB3iWJybboHnxyJXrLYTbc4B+NGSgtJpPI
eKj7hnu+23VxRQ+8MF2I3eIMzKcRtvG9O7pnkkULNUvuxpzPTnwhqbQ3eSxp
qcuRe2LgTHjJ4sZr/a9OfWamX72aeM4D6WiPtMaH4tTltuVaSIr+Fy+pkkq7
CH2GremE3Eun1ya/HM2DjEb1mRhsNYnhVaVTm6xPvClkWJcBeQVPmuxFlvnU
thjTKdVLgUM2bfka4BGJyUttypQ2IeNHv2mdH968FNnTEjuAD/mHKcRFFol3
98UD4c1k2GjDxusMR5xxhh9Ka9ht6/6WQGXWd5CPNJEClDo1xRj/2e0omXMW
hECGBp4Kst1owP81n/FIPyFRwohv+0BCfdDTok2Cd4wAoJYyma5MnuPQZlJO
xrFsC7kQReLbn3fDmruw+lpBfsUV9I9iui5mlHNhLItX/bAxB7pUkLKQ8o5F
jCBNZa+ErWFPI2YZ2UohcFsjBGTC+nhDCkn4hv5nxQNziQTrfbZD0YjR1B7P
BxULXXWg0pqWUlBAp89m3ixGJJhRg+cyOQdMviQFhj00MKC0WMJxrNVzD4Qm
BswxBVV0T4u0DhKgkr9SlF3Q1QtREyhwrl+/pIU7eFf3URIJyTNfmf4m1QWI
YUQ/wR8zKaNBGIVh0b9LpinXJaJvJ+NpW+y0ZJ8yTBxg+/+8OGxcQH7IwIap
lg1HK0bDygYlJjgYraX5Z3ONjRqvvFhjuEVnYSMByFdvrcl0D10Gv5lxWa40
F5fy1/v7pfTTHSE1IsgIBnm+dhta5HMv6oBku3/F5i6rzbFPv3SaOJNyRkvR
7LQmNZVUcChpNXP6DfSx6ky21r61cOzHtxcTj+gOEz1Ap2W8QHi3THqsCr2w
YyHM2/kj9HcWh6Pu8UtO+/Ps4q8mpxpiua8FFzJuoxXbu21Ovgi0d5mGowO8
lbmdRPJp34dj9Xm7xHddUY9xid0jSoIq3H1DR23YL3m8p71t0XYnzvOQi70m
yzfFHRdtVikccx92Hg8Us5xOytrRe64dHYpAD+Lvcvw1uI7MjihOrhs44Dsn
NXxUgk68yptd5KATXBY9fKiNp5hnFLdnOzzxuYvWW9+KkHxRS2TXWqlYfab3
CeyIuZdA30MnaicaS/wFxTNQqggFvzbqZtcKYtIjOVONfu2TMeBnniFoPhvj
CdrcWEskCBoClwUoIggjOE59ADnHIdVnW6AvIee4bM/BHUbL5Ie6X2wg124h
N+1ial8A1z+TjF+qHKdT6Z6q4yu8cDx//hpQ+upfNicYISoqNQHLX+USe1VR
z8ANLE/LyUuSrwkZvvhCD2+b9wciNAJujy4tYtHtGWVN52rPcvh0lPxh1W0w
wZYvdAJKrXQ+ZWwYyMj+lH8JZN5NAealCjswbSWWV6CmqJedB1tNJSwspH/m
0FgH9yFezMiPipbEU0EcDlEa14rIkI3TMaCoCV+kE+TjuyvFhgLZ/EaDP80F
zytjI+GSOWn0f+x2pkxhgWZ/08mGMDnfViVvBv+3MnD5hciVheOUb3EYV0bi
URi7W6o8c9VIiFWM22fv5rIEJSuZw8f++RPTup+PQBTvTPpcSM42e6/VqqsS
t44QKpavaCqvizYzc8yFmUxOb83hLJDKvsM9X5J0tm+xEb+6liconGLlfNz5
flpTzIdMs1qScacsV6VGBtP3w8++pAV8OlRuMU+c79xan6JOmKDgiOnkMWf/
ZfDg7+FcHt3yW7w/7tplsbIJFO9YrHFttAv26gj3gWUtK4zlCAthrA/LAgL9
2rBmhTdIaG/iESSKfM83e5BcJMh+zheZ3e4VqOzv5MYZavW/FTXbin02bwWy
KRgYIrh7UyCiGs7TM9bovkVObsM0Q3rMEsuniUDwaHNZxQeyZZGz9SjCt1w5
o7eA+0XnIE3JSPlajgSULd5WkR5MlDWDARx1YHeuRPzHHAvT+kC3M1kEbg5A
wEEpDna3PGPW4n7mYQK5deAo/eu+XgO0yQf4iqvp+B9YHOk28kl4J7phh9/b
7xDucBENmi9/SQn4RjEJvSRiYf+pvZpOe7kIdNAMGsPxV+BqP0qfhhJH1Tu6
1i9vZjAeaRDHw1G3sTUF3kRX9EmrEdh1QuR1utMo+ZhmBkMYMTDhT9tarpLX
bxExs6gLmWFNe/6F9k4PATC7DNy+T81vQfEvbhHTWN7DUMNbHoMqGvpyy/js
jqC1VZbCGqvDXhTuioWQ7Cq9BaTYVP6Fxpa1xWcRE3XNjvhxUXvmGyeZ8JkT
NyFQRtgXOdjgkr/SY+QuNfZapOdtm/wDDym/3I8QTaS7c91b4UlxaKZ7YuX0
brbJ+RyMZPhv/ibsznNgXRmBzE0cF0mLkgbNUaPDtzTrgSw0TCuRvNOO9/XU
2NZl932VuNf8o2yVXPpDVvS5185InWWIdSBBfKY/zgHLx+n6IsKwuUqrmkta
6KwnamiXyvXsi5yC9oyrxy53FHsXMV1ex5WONKwBPFlQUKHpf9xXo0xBcuz9
vhIi5UVhobIp7vZXgsRt25GbRAObO9cP495PYP/lQYUP6b5qawprZrREO7aw
+IVM3ymJjfVfE1zkBtCgjyVcATWsM2OvBZLSzvWHHRIdUj3x43rFLg44Qe+j
23g+R/j2g38jrVwjJYhdnnfMKWcFw+qW3lMcE1TsC/7vZlCTiuv83BSW67Ov
Z1s9aSvVkwhPerkeVbQgUm3cAq2JcB0dD8AsGrtacY+XOwWkQNf5xpvqsAlq
0nFecLILeHmISbwrn1iQn+Wyna1qiSnLhyv4u27RcPYZjq1qO7xoMkVvwi1Z
uWx4FIKRGQyq0XE2XpK1HtSuJAxQ1en1SrOsSA3s3L1Ib1VCgtZ2Tg/ZFXLS
JoFhUraOtzt/ldnYPf8Eb5l8unZJy0wxF9czJN7VyDUWnHhOQkjakQzjt4eb
51/rEv8mMULG/VWGmMR+BwlW0qSpYP7fJnpeg2Ivl0IKmn1jsjGtWdXbn0Wb
d8IB3aqdAuhIozAIzFBClOsmbAynfiUxcAQsL2bwPsLi2bwAGo6zHLi5n1JF
9j2qxy5lreUVg+uTGCTGhyILDR/y+ih2UzEiEeZD4GLVBrxCyscZ8Wk4wO0s
ugKwmmvtu4H2HWZTFz96YwfE+tBDssQ8hK2qdF4PvAgGTsFXQiKT14k1VMTG
vRH9QjDesXJNaMb8JXkoMCelV9GexofJNJWPQYe8sRStSsbWkgtdoh9D0fSL
mSUPETljLgh2t1JQathSB26oMh9CMynhIF56S6OfhNfOl4fGOSpZSo3ycU7+
d+1gr3ppuU5veDIvgWB8Tg9zLlxE6mw7oLQFTw+Nb6T+PIdwWn5SZKAptOCF
UxnsFgN0YLXQV3BpfJ+l0DBK642kL5TthVac+43+DNrfS4OYge77VCYSu+hh
/vkJMG6viU2R5BDPX1AWc2VyUFVsSB1fLn7ZURPpRbNRqMbBhFGR1yXIggoP
+e4ewOILmhcQFPmqErzETM6SoQYKjsMfvfmBrU8iu1PU9TXMEjllrTIjG/Fo
+D5uFxpk1SKFSiU27gZkFEs62rw+HFpSf1o+A4vxf6HmfVJ82ROO+P7LS8cY
hgrYoVAA8E/0k/60ujaBCIp6gaKY4pQOXhcFHAC5UH0ZBg6FdyslgXB+LfJh
jdW17YDKrB/T6iUpT3cNRbxh/VWgj0MKJwhpBGTJKpBu+Ni16saTeWDAbAva
0X+dSYc8YEFm8hVMfUnKAokW3Ph2K4hnMGwyxmtTpUXQxTfLEZXhPpVOLDjd
gSdymQQoD+88Yn9+F16c4e5uP+NqMr40eTqu9BLXQdz36/2KI/lBX0x7PQhG
YLhElJhxb3FAnFszQwQ77W4sqMLQaddIDnsnphWnmwMXRRplW+HYekvCtzdu
4BklHkCiZA0yb7I/UEKq6qJT5tEcDEvUPmwvWiq5ButNB0QXD6vCClVvmjb2
uqVy7mw59HqhfosfzIn5Z7ztgYk/CP1PboA7bxQR7+T6jcL7agZpkwvWXKG7
I/YQxous3wavR0wOlSV558lZtAfovyW02D52JwaWQnBJ8Ppxjra2VyaeHnnp
6ZWfWVTfj/fw2CfQCCr7PcROdUUDDU02vu63BE1sPUFSx2bZuSZERomA2xfB
eNUxL8WjDlx8vlJugUWu3ZbvFsMnLxzyBOhBtOHaXJXdN2jbseKC3GfS+5sD
MWp8T9L8ENXoCSfn4G2QbQNTn9r1osJR28gtdkxdLPWEaOk+az2EXMLdnsSs
zsl4ljb7BK6S3X0Hi+Hp2d8JgK36Wb+uYdwzZwOV/VWMHhdMYHJ65dD874Ox
Qoy8YZxHK3sfzWezyhknEs7yfPo16nD05jQnTCCVMG93FcxjddFjE/HxDMKK
YgxIFBbk8jZW9DwtodpGCyCsyKtVMRdCDS3+vbiDV0iCGyySZHC9+wH7OWZV
nK7C+ZQELluduB2jJ3rVeZYfOmj/LNBNJWhrqtSyNlnKk4o9NuQxS4eKCkYT
iNYQmeA7z2Haqz63dWPa3LWoSD4J0rXSE5/rQz8Ws+Q2G1C6vTjQffGZO6/S
VJZT7pSEufDahKLlmJ5k1WOWyfx4G8b1DPccgzA6GUQpSlpFk2d0fPbDkA1d
oC23UUdnm01vois0p8q9oBZXnDXKsOSOyd7Zww3jMO2/OvfjPKw4//KyA/hY
9VAJ6tuZytHH+mNCtiQekiFIZHJUpTW68LkD5wvhRKh75Kcz61RdFE/n9Ir4
FPjN+c2bZ6UKjG7TPzQcYjj/TzyQWatsYVqADg8zNtTguZefXgqQPAnc1/RS
twWQsB+FWxVejpP4qpTR9eeZWLtY0LUFAnkne49SH7JSmFLzfDnz886juMeQ
6EBa45S/HSIUNPoFNq62BcmIvF9Qhjyc5yXXxla42n/UZVFsF+ERxpWG3FhH
X/rQKEM4wb0lH8juk8izV7y9t76BgjsvhObgMLVnA6ER+21yQ+2nxvWWZZa1
ADoJKYfoVQBx3mTP23QvxwCNc6X+dR3KV2+IgLtnsIxg220pVVEkpKoTQhnA
SZ0/iDblyabBLUnss9toAMOYP5uEQgAYgEwdbYF/yCQjbHjezljxoGRfdPvk
Q3rw9zQtCzAkxtxK6mrGH3U4qLzo/t3nCZZQKl2htOO5PnIgeZ8Pl1s3QDBS
2RoJpsBx4Ji5rwb604CkB6bdiBr3wkQglE+GqkCTRnYPYvRfQph3lMiBualh
R6FrqHm4bxshJde/4lOds0Du5GIXsuVLnK1YbfTl4ogY6FhEcL/5pjwgJs7P
2RcLSC/saULc6VclyQrUcOmCUra2a1TuQPL+m8kx/1yD8LWReQhPE9ZM2hFX
noRoV74zWqpnWBN757Vr32ZubooNBlngnqtqk1cHOe93h79KZmOUJmpThjQY
q4EQVW39/QObqo6Ooz5NyNACyOkwfkvCzvGuxXzp8uC3gzlyoIRwz0EtOvX2
F/XNZBTxANK0EOVizTYprd9LxO2trlqh5Cau5bjLMnOHsquYa91Qya6NuYFk
XEK/M8xjM4anWH7/DxlvgMoCJxbaxq1SbhP66wxT14cDzfKUpzfwhlccUS+h
JXoAmOVdOKUU13oVlMmoP0a0ZzHWRntGzj8vRP1JeEs/EyAh4x/uD7oxCHJu
qXU5GgGYlP9yGb+cKWYG+e12BNh8VwyihRBUzL7x5SACuHlPb1KngCA2EENm
gpWUjzEiGaQHneMHDRKNgZ1oBauYka8uVsnpsyv5BkpscdEm30abQoXlqIh9
zv9/9KqkozM0DtfMxExwcMNZmUc7DXJzYg0syGc77QpOOqb6O9A7RF7tF4tc
+X0osU0Vy96HNVm4l5vMn0PlvL1DZbnyZF7qObTPF4U+IBMb1V2xBB5LKZ1r
QNzYxWMGy5V21ed+By0vG85aNnGUe58i5XnHZeAc5V+uGC8VRmjZry6i6Yn8
6vB18yvz5ijSkEN2UEd1gAMbCAhIwr/YUJBsEk6WBLxpLKpLLO1C2fyvkALY
V/hpqBVbdndSP+ixMyghMDZZ2l7efQYOSDxJjv60u024VjFaTBTRGBHKYVYR
tZBWLAOh0nhXFItMeamegLgkJu32EVUnhXigKL1uH8VX6gddRtU3C+ufwyVe
cLsKaAwEMB2A3nGso2gtqxAyhIKSsG8xITlt3t0uPCqob1m62gerrI9jKdCo
RSfc5LHYkt2efWgU+2ga9PMkAv8hajTSVvZAgHSjH/2jApegraVCACuimU0F
hENusiTfRtQvHrs1ahqjyfh7yYqDSRbsSG75JCdulSM05Cj3Ge36W1gQU+Pr
KpDKAIb2YKAFmyfXhz2KmocdnlJ4bz7pgx7IOsQiI21UoZbVwoO6jiiesbHn
LfV4rlX8/9oBPZ3I9USpgN/ZZ2wE0yPw3p0prZH3RJhbhGOWaYBtvHpIdVjj
CATzAHbhEWJNpC38ytXx47meXu6g5guJXyRev9/CMoqhkLqBH5zB0cdIlZTM
YUJjHLgfWOm8ENfbuv9pm9BDRFgkrFEo1Z425wF4h+EJiyQZtpAW9Kv2jlrx
kvyYmpxwyuF2wGdpc+mws2dtoHq4gMHoQfpP/qVBRY3sW4aoUUHM5EIt/wSK
Af2OmW91aax2PT1yzm4TYHnX6guKEsgFxyFfK4xpwFCwucKX2j+j2I+lPqwE
z/3Lapg/avNx+INXIVi4tbHGZEm3KO4+fBqf8Zsr3fgumbtnBsskYZlLeFz3
1jEMA0GlYQKEJNbBi+uKgnxMUOi1IUhdMpKaSagVBPu5i+z5scfCxL1Sc6Gp
t8xu0G1GkPGoalq8tIOFp7mMtT/YUHWqlHNe5J84Ve/o0sx9uDjLY9cjjpWG
sZyBeOxsIs2Enz1MVRQyw5BFXYNT+b+dPpqzX50pZpjvtLXmhIbo9/wtJhUd
1AwsMw4CUntG4BtMaXc3sucpMpVqZs/tIheyfaCsc6w1dc4Usjqju8uyidO6
IRh8fJdGw+qMfi9dquS0Thfh8en0I2D5vH+38f74MuFmIrVXACV5H5UD7p4L
8XmmIzHq1uBNp0KlW5RjrIFR7TVo3KvYpBEEiMb8g+ojEm+dA7pA9mDFwP0f
VmjK6LL0AQALQbOEHS8mdAXVGrKCslaDHz77YiVSRoAY3C2AzbWdYRCprIiG
LkgVnOZbNyivPLf/wABvQDgolPllQ3ij+zM27cSvaP/0ErkIc2rkdL3vOYyA
0ZbUXIzXa3FzDs0pq4QmmIvW01Fpld+C2bXhmnF8WHZgHCMV78PQd39/fZn+
d6gXMFkdU9yUZnrjKd0Au9hYHTqnqy2GSHHD3j9rVsnVfVKzdp3GZFF0iOfy
LR077xpTbC8BH4DXzZav/HWntyU4ZAqttJm5GnJ3aWWKvpDejCwjucPCpdCZ
rQKTEo53FWhjGfCQDe2rMo8wQAG9cawkSyzSyvmQ9egPY8XzbpZQ538suTDF
UoevTg9DsmcSbvF10kTkKVfywQB3sc7Kqhl7iRaZz+rmx4p5p4nEhF4W7DNE
dm1eXGLaQKKVAVIl0W8Gw/R6/Uws+W5uV2hrNkxFB1LLo5sGjiJy9Ji6aRwj
sgpHlgj1TWasYKbGwqTvaqpbYnspUMGxnH3pRZ66hc4YF/jxfOapAda9Btpm
c2X3VD9LdcGesDr9m7LsJpJ10x/GZbcVd/ucbxW+b7BsGuGGiwoczYMoz/sh
hljQYiqBCgrg32BaIa3xpxOuTsap/x9D5s7sv0Ysfx7Y6y1WTxJI3r2sGPRW
ALxy1Gv4sncLweb5wuwI/YrHcewab+T/8VzpGJo3rwrDWkbJVbUUWXkSiGNV
fQIEnTCAvy3PvdT9/Swzh8OWDH79b1ExmnLTqz0BxYLoXcJuCWxtee0272G9
oNI8tAqZ7lCqz86WLCpEzcuFJN70zVJ/8FWCFIc4SIcgak1ke3K8+xvmhBXj
IrasgwD70SWUVKgfBmZbR713QkRuonqMZ8V9knS719isaaEvlgji02xswfxC
t3kvhYt2PDQML+4+3NYNRzWW6YS4Ei28yTuFJ8GR5P37UhzdiumZ7NtJoVnv
IVZaoNCzD4v0enim7VksNKDNGjPckwUdOTUr5EOjTgV2LTGwnEwRU/nXETAY
JAoW7inM72Ux7gf6hncTIvzIEeBzv5kinW4+JhKQN//1sErPuLStIVdcw+Lh
bbbMnXG5MJbe7tEXvYAs9gzrltJ18H04mQunmb7+RhwizGN/Esj+gnTwqBJq
1wPVeyMzdNxCCIAKLsS0BKK2cGUghjEbCGWLXSWG5d0oVf2BUMITx8xBWuze
84X4j6FJF5AE89IVhH+dyTvba1JSQsiJMnKOgcOozGfdd2PUBqiipZupfAmD
nauUjsSwadDjdv1EoWKUJhX8dycDAR7uMDflrZlDdvihugKE1rknGBSANgfL
U8XPSFW6gk6M8oBPCeXcSNFK7oDuexawqfVMmrtDgPFnMlOsihtnTr51KPAw
tFNIe1pBJeVXtwMlUSYg33ZaFkwfZuHl3lUjE9s6UcGXZMUMLmXJsh/Ku51q
y8JaRyAQandXsK1svb604TIUbG9qGPwqfFiV4AA+Jt0tHO+X/XqTBrLaQxy0
McSm0SNFz/TxSedW/u09XXdwHvq9S9VgzozgRoyUrf4BcsLqDFYT/5iY/qnS
wLA5xpX5MfgxFLhUYLKbNKNvSxZA8/csJS0DnH/iLEYC1D3tyIYhXk/dGKco
4WqY6LrpozFlmUO8NBjwosNIBUJPWhJlG60lMHJ0zTlNVD2TzRnZ0prufrWd
ks0NSeFRQ7F844IhvRve/EMdg25DeEWj4Row1P5bsiwF8VK6tFAYeftqbtKS
j6fsZBNbSrAJuEpQYcsTZHxQiXL0SwQkcqli8cEFVeq/3lAs1CtWIHjW6N5O
0kIZven4M+ONqXEp2avZjVMySUXx8rz3gubCsyUX2O7qFcGSd6an/IrUbHEn
gI9SlOkp1RcekuB4t6EACg12wCQkgivajznIpqO6rw53pi/Ay7HcLgT03+dj
E6DgjguxThCnwIWO2BMOXxL6Ielr4FeWdFHBijML7ruX0llDqk2pBiRAMr51
RabvvXBWcUNiuw/x+ylkwQ6tnc846qts+fvN+A08vOxSNX4IcSGLQWA4saOj
byPBbVTJQOPuoIF8v7v4yMvWxONKKmPGlEX9u7a1URTi9gao2qAWPL5Or6kM
Gv0A4KfT1CoZddgqdS/xSopI6YNhRqjya7f+io7cdKV66QVzhndHQQfZjfgF
BjS9OQakan6XAkUyGUYEAGc7N7TNomH0i6s8v4+pCbTdq0sQ98GrkYEGfaDf
9OBP81/QJ6zCK8hgs0deUF8tBc5T10legG6gDbj0xI19/3KzqWztdsiru5+R
6yuZJIHyVNnkQrTyZFy/ztaLurT6y9HRmFHJEdUZPDK91zq1xOgpJnhQMC9J
S1+y9L/iGB10iLTtGnrHBoT/bUIaxe1rqmmxwWNz11c/Nsocl+svOILcS1l5
QFJUELrmPd+zXJYzporarpxUHYBerFD5ye27BdCdP+VHEbeTfvKdvGZv/DW2
6XJYqk8Om5JFJYoGbxuoTHa/1ORRnHJCaO8MXW4Y9IvMbi00V7WYJEfnKJxo
nRvdD8IdBYZwvs/Iitvp2n4FrQSFIhWA+NX96V2Hb3oav/dHLgxeVABa0ety
N8i7p/z16dhqfibz8G8mSBczlaNQ0QAG4cYYVmQmUjVCQmnLyOJds+UmRx2c
GrE3ffcNNupUgdp10y8F7Ka6TuKtKBjxyh1hUb9g8sEHNcFGYaeQoq0HN9gJ
3qd3CL03fdNI+jqHtTLm3K5I5xPaXH4KHFacSOJ2nAug6akY6lSVqfc9GcNY
3+PY09sS5McIPi+uDunRClyOxTlLYAs2twLbqfrz5zRuORbFWmOnEsDxVSVo
/8CMYVZkeco3MTJGRTGHxMCQ9ycxK28XKt7Tsi5Ot07+NmHR8tY+m9rFVijo
2NHhKXLxrLBiY9QjVmbB/S6p8yyft7K31fVfdMc4OoRTYDajj3CbSswi3lLa
UZdYtUpMklr3MXC+F0l33XQFC5zFaaVOaOc3Rr9oVXUpt2xAoe3hzfk9QSmh
rWGccHXAtSKnM5g+/UGDyVpIRGj77D/M7/tpxOFI2XRLt5pPZPCl3yczaCw+
Qvawr9o4tV3TAPRhTNey3weA0bG+l6flqlAaQr2Ps6+mIQNTzhNBPScOvIlp
fqMSeip4M+1POrFLV2loq4rKz9Fw6TjSItUJKQRF38m1mqXcPWSpRMFn6aY5
Q7/Z/5WqFtO1582IeiFcSU4RxUjD/x3ouoF8P6wOtqqBUQ8JEt2byLtf8JX0
Lr89kMpABHDFvfA1ipf8g+7/y/BXHk8IG6YZFuvrmw3bib5vlhRfg46DPlKH
v3EthlC5iviIsJrfzGBzI3hTzA6GTOqv455VKQerrIfff+Z/Gxqryl4jdC45
AvjLNosG89ROVfncRz6ERE9Kdldkyp+TGSyAHqDmRWCcfNwnaz6s5XtNITRL
Gbj5hbP/yBcaPpimOiWJzI4KFTSWY5HMcQBy7jFnj03xX6EI1ai644A+hqWp
3n/O22Sq1mq8Pb7zPCXEwTlxZxoviWdndRolx5msohDRw8ZneuE/PAyWg/OC
43924DcGErC8q5KG3/kH0bHJ4J/q15x2Ase3cBSIn8C4MNVcervHgmxYFum6
9IabFSRZPpRA3aamd/1p0PfAgYe/p492tJswDla3NvmENgJvztw1VUwyOkey
g2LdlAUtgCOteIdTVCsu4nl+KCbQinlUp7HwwpQoR5ZbUcBUjK0SamcuLTBP
NsS98ud5Q/MAQX5Y5aG5lAL4imVrjGxIzeAgDzLEyujdnlxcw+ugATjW7lZ+
ZTmxFIS2+tJzaI+1Cm1YdCv0htJqezF9Dl68HiO24cLp+zyo9AfV+V7AVbT8
hwRXm6hz2B+Y1sYBBysol7Y8TaKQQFeh7dQnDJzQecq5OoiT00bIaIpyeV3M
gJCeZLMy1c+InvmX4QCJJKnJRlssEL8uACg9BbcTK5/HCY1crNEWACc3JYhy
BL7hrjt3q/jF0yBdDREXLIHtnTQ5+0QAmhIYz3hP2aTrVfsfykjgYkS6kL+q
oKbDX3f8p+5giJmEisgZfcTm7wBhAhkuUnAYNNS4DOKAs/0GCOPz8EDmEQ5w
sm8AEhiiDx8e1GXWiZAzP1I3vC3vjFv0yucgHvDgEffVEPTRCRw9rKKO9t+U
D4K3/Xena7kMZ4O69SrXPsorWabgBl3elUXx2ncjaafwR9h81ZPNbioiGiI2
gqVe+MHi1/yHT6XW/lcEOao6MKo0wwgo0eQ/VT4Uso8zfIW83fhGoTUvQJ9m
FF389erraSRsIQguTecLbou/95uH1sm9hYV9qUXiG4r7rthk+1SzEbrKqlik
e+mNQ74opFDnQEk+Iny9LXgTpVHljeH6vQC5qjVQPXmDheg9iOfhx0e6qKQa
njd4Uw36fXaIDCR+goiZnb4KNTpT24shmKfwXmMlvIg7nB4iejJ+CC6m56Xg
MVw8bcNg8bEKkabRfaYP2JqqSQhZOmIxTEnS6m2eCwm/Y37QuTxwzI0fvX5a
lkdRqwV9me9OpThRX8BEX1Eh+776GD6CeuarGpf9x+y6cJ5R7Y9CfvQlrXGZ
9TUPdoa2iDGDlviVeWp32eZx4N9qno0rqK43QuEDi3GTN76XbwXK83/kZ95E
SVfYd9m7TEBikA8XQ2P4wLnRkWgcOsdWcptJaQVgONjBQCb1ARFdr/fj/33j
j3KxoOOdtyCTyrSCRA5m1y6UDncbM01dXDbqOjwDYlMZUf3sJYVPkNF9biQN
LSkPY1SSZXUwOllRNKP8iPaBNOd6YxAGaBSINXKC7MTFCIDiGS4nt8wbYmkR
IqSxfcJ2F36SkC9WFtsx96tkEZKN6ezhdDIevuK/a0LyLl3dkzXh/kyGKl2+
zjjqrFOF03mRLF8YqxUE8HIGocTCuyAyHggrtuqCJvQgmfaufJ484cMf4SjU
V+tgVW1cfKth0H5LQp0Puf7sa+Mjt6zti05E6JgKNYZ20sabvHST6izzr1FR
bn99eR4nNE53W32ov2RXhoShkKrGqdA8Kp5+A/rg2NxharYfWZ5vh/iZdftR
pW1Q/xQxLcK42yn3g0JKjcOGSeHb+pBIV6XhmHZrulBoPxbyspWRvzY6+APW
zQqez1ijwZ51+4lOQ+Uuh6swgagLxiqngTQEW3uNYkiX48Eqo74YeU7Sqj8c
agr5q9q4WkALBj6Si8ahi0dNJfHwXvipYxMiZVKm1AFySuRJgeNNB80oTfFq
YM3FY9Y/FskqsrW4hwtZ1uMNTNrJgQC6TjLkjCMiymcICpMDR49D0FHqQfyb
BZasGpgAzs4ZnhwXH3RQXxSDuevvze8hyCDOgAF1/SJb8V9oO/3YYw+BBRfs
1tJuAoPLSXorelTVJwqtMFxRVy3WrV7ddN5UE+JqU/g8clxjqtHEsbi0UbfE
qbVr2Nh5nKBxVIIeltDNv0xnUpMY1nEpDUdwGhZPkHleOaGxxRxgM0mwebrP
aQKotwOctItON5DkFjrxd/Wv+UCArAM7xPqHdXSiVRiMq+OVewF/wYwYz1s1
8rCGOVZIGKTWy0qwglhQkEo5Maiqoad9XK9rnK/zEp4+39GDfA4sB9/V+kip
ovK/wmhv9aShSrBOC5CGdI0kgbc+zt4CHcBqMT0BVzfnJ5PbGDh48MOVYWeB
8fsreVQ2OnMvoe3/jJwdySUMnvIHF7FkqdDqmOCbaZotRhMKNtMjCm31UJrs
Ja4NqI9vN0mTdV36x7T3+z/mbmhkrlu3Wfz0IH/cUHPDVPAEoTTmmNbaixfY
3zreIwLifBAaR0DxXKhGbtPGcup01JgSTOopQuydgfj2gNtC0rk7ZMTN4mt+
nIC7+iRf8XMnHQFPtfgTJ/KnrpPrFflnkNPtwUG9i4lk5y4VwbukdMBbOkTp
rmF0OnSQRu959LJWCLbyUBElPt39l4ih20xAYGVHQ4FNs+FkTKhGRufthHgs
B348doxzVOX0A6R1heQc5but6D/zi6tWUg4FLqPZeNmiqtJhy63oIBLgCuQQ
bybPpFGio/cQs04kzV+NhUxrDR4VqpzGvHaf8x0VL0H9oOQFlc4LLiacb4qZ
hojTD5XrWU8Qen4RyFiKZx5f/+r2ls6MAbewx98+FXwR2AzpfvHEGiSzEPW7
q2lu4/GLx7HH+7Rcxp0JJvYOkJp7E8lZaYo5HzSUkR/6cMTZqie5ijZ2vO5X
yUT/yYGdBsAIDblXktybxQDm2vk+6lhEXRJO75jbZ3fjXhyEFzdTBPHtliq3
eHzVgP6tRCCvS3oTXDrJMvYAiiVbXxUKSjP6AozKFLAeEnwoXvAFrYIA22n3
ddHKwVzOXoIFR1JO0NaVLe6xxZl9IjH+59d3hm53GSZJ/B4dwB1ZhW3bhNI+
aZEMPStil+xu86xmbZbw/Hk3I4Q/Yn3wwAvHNGOZhMLLhUt/5mx6oIMSm/J3
pPPdI0Z9/F4it9GyKV4TYatV2PzQ5rqbf8Z2d/tzCJeF+WO92Ln7Tt0C8fQm
3mh8Y1axYqXaXljJZvGQY7EMfpXFJh8nUpmvD6htmty8gv0KI8PaDcskdX5t
YcwGb3ce/QfrjFN3CoYBTGjcwoKifEsmKrUaYXIC8tBueOnfksAxRTrPaqwd
Fqw1ZYhHkSLVxXCyR9DkB7VvxVq1blow880vngGw4W9Ggyfu/Dr1e4VVCG92
LQTyolxKH4RaysvvO94Wi/Lb9Wc3d5WVUs4/8LjRQdFYb6R5BJrMaMiwXbxU
nEn0mwc7Toboi76LsEMVxIDQNJ5wLHA0MoV2L/9AeGIcWHfKeMVaL7DVWzzP
YOpI7kOo2roX6GbaZVkn0vTgWWU2t/pJRc6YdtQS+KzMFJ7PwHUiBjO5hHNU
SMhAm6hdsmzTUXR0abL1yIYlvqRZGuX0ujDJuXrDTR58ZJwy4gZivjfx4kP5
3gLlieDV8h8egXzJP7U+LXr8W3C4oYP5KTGapufMVHgmP7SjIhoLErtgYDuV
+maSBlxIHSFcD+Wq+zL/6MzEzYovm8K5hbDelLZhWo4GwEn/cjFAFppBcb1D
P/JmOjJNO8nuN5WXP8hbSpVJtaAZVt/TceL4ytqiLg8i4s1C3IWSoxYoGpb1
F68LIY1fzLb/BvPGmyJGqAYFS7yXhox3xu3Wb5bB41blcS8vWXYyDcJ1npH/
l84kHW4ASHo7fEBHri/XMis8bRidB0CRHq+uyKyP1cD/s4ZzthNxKdH70XU+
gjZ2KI+Y3BcAHmlVd5zfkmAHRSxaS/oL2wA9sRteJQiIwy3dSHjGfvtcUdyT
9s/gPjRfvgTMRIXBGSn5WF4O5ohfkNGE+k9VxISfSPF+uxX98CN808ybgH/e
3OBKGDz9uqSBTK4Lu3tolSFX0V/piznHw6DUpGw/4JljV5V2ZdlrDfVGNryU
BFbnGdLa9OxIClJZMO42NBRr6q94t+q5+obzfrcT5t2sshUlGT5CyU/jqf3I
i+7IzfzvaGeGk6eX8soqawD+dlm4RZTdEwoLzBbJQRKsakCri+vV4d4S3Xq2
MYRGa3h2gxinIdkJj1zDjPQ+v+naBu2rjyaok/LG3CAaUBw73sA43nxO0FY0
SHY1hfpOc3RQSifoEAp8i2eyRS+QVBiA/CngCuz/YwRdDvPdo4L2Tnwz7MyE
cIQcLl+YjA6AzEEF6/iWdvx312kak+m7uL5s3xbGugUq/NkdKBCOyyVl3duE
Ta369oduDTey8ngUV+WGj1FdAQaRZJRi2EGe/dfCT+lUunJEzzbYcdT5ep4Z
1x40Mwrb2zTMZbxfyKOBqAZxxNcZ5sM4cgiJqyJqFcPHZ1tbFjo40NRAVGJE
btLzhjcHSqPwTGe5gpzEvmbhtPpEHUyNN3tk7+1pk7zndlTsFh8EUWA9U+vT
IepeiNzb2+D3R2WX7qSF7361ZJdxG2jneYKheyzw1LqTJ3zkS1KL/LiM3rzS
U2SAkT6URnQZ/HJk8PevnQ9GlU1nkNweNd6p92qK31AVfIdqJJXIDTeJbe/W
dWrUdYMObEQidWgxGkqB9IVk3ElXX5PT1lAPwcGDpY77Z50B0kgqArh8/4sa
8H69cNNPSUFX3n+LgCBnPL4fxUcbix0G4a+mUrZxogpCMt9l/5CUrz/gnUr+
dSgKsFVlqdYViVyFYfWoO+PQSlCKlmusAFRjpg0DXDLtuTVe6s9t4U9bu0Zi
T3/Dux8y8Wpd5m1TW0dPOKim/BVLV2G9rLVUz+NX3hBDxlh+rgzyUfnHWKOt
cP7hDYPlMSvSTiIIs67ZZAlNnWED8FlLnm0ew8k5nMtoAHKkQI5M2k6MfFX7
c8xq7NgGd9Tz5ewEYp/cq68dkguW7O6PhW0jx0CrPf9ktU3a4y/SG9bcGF05
CSat36OJmBDkh31FkqR9948YLpwY23Q0M6nDturBrU2R38e6BIdyWyWoVJ4j
KDuWtyD379AXWPiZITTPtiKJ0Ij6NijHBQKJ9WEz2mcL4khbFQYygmiKrisK
zbot//GxrVyXGnenqTYluM17xqnhcMhk1jy/yAbPpFijqogjW+h7Wqiy52VG
DsXu9cPbea0TG8JK0fXcJCvcCFPyWCpe0w9SrAad8GJwPzBRiXyS7Swacibw
Rs3WTAwatjBwjW6uSLY3qMSDfeujljikyHmj10LycREli+MEhac4QRAupMWv
zN9RmieeSyMecScIIhfdBLCLEQKM14IlvV+rfGLL8UfTegzfxv1EaVJodIbR
ObnnHOZLwohg7MtfIlAnxoyNMcSJqNqfDQ8wnbdBhJigncjI01vkxxMicTY5
NNyoUQY9BwVX4iezfhFx7h1QKUSrF+JhA4GcDMLBB0ZMmeJY9KxA81tiofrH
9GMJyDFLpT2WHaQs6fW9haIakGBZeX+8b5a0JC9LI65BZ6z6tBgfKVcDoGmB
gIfURqHEm6xdjH5M4bdPcmLsPGPDuSAFloe9qAYPIJSEU7VHumXVkWiH0z+4
bkpFxGXk7VDtatlsRWXCFYFiOYS3HvJCZNq4AVZlT6ZVBIz6SxlJTcBr0qqe
IRQxYre6m1w0QKaqy6Js7JmQSYjQ4VvQjpRCcN8G+R4dYqbeH7v08LkcNRhD
j35fBwzDOJLLZ4kZeUAVLaKYyWO2Wbyt8KwOFxJp/CpZFZbHYIJq/a3VZTyg
WSjRju48N8wbzbdnCaHxbFZ7pL5RO53JfeFDeccRPrggXjiVJ9uYmRIIpBtc
Ww/1ND/1pjVvHFAtZOP7P6OjDzDNsst3avqwvXfg5e4UFWQ+zq55FHVrElAY
rn1eOy2avxeY0a6i8KDBFfMyEEdm8VAbh1uK8kdWLer+ABvorKfCpEBqH/hc
qEzwis8Nh5MNkjeCjgoYGYITH3acXLJbZXm+AogMSZ7nokGroVsxqUC0u7fb
KDCMdl3QWigDnMuzWgvGP9rdZ48KFh4TE1uuNPZafAnETIcwOUZ2K9XNNjar
USjnpzWfNQq6OD0d/YiLS4kQctW0yp/hV7xwDOP0/+qK0Moligh3F+2Kmh7n
8AkdEPx5KMgChMZkIeVxnnAQUMtx5a8XkdhBMYIIWx8tl+0BOSqPqiHYBGeI
LRG2KIMKjaRY0S4tTbM5vJ4VceNhdghaH5zbPC2/7LGXLlOLxwNoz1lBcTS8
4Rv0BtQoxXP5Aur0HKqlfl60d7+3LdCBEvJANSrfW20+3/wvxC1Kf+ZxxZF+
lDBRTw5pXtIun6/8lZPk3SzctzF5xYApqow2EoP5T2OQE/0jf5i7RK2wd1T7
Lyvm2PyvC9CpCp1XEyAVujWvgdzFsqxBxqhPnlFamG8VE4Gy6wSBzvKEXyEu
71WCg647wu++iZLpGQfbjaI8rN9JoesA2wiuRCM9a7sDtGVtHVkBYSq6yNL7
NRNji3mWW697uwAVTDTP6Cmj1wsM5YxkrbEfakAqk+rYZWTahM43o4M6LkeC
+c2DYHhMt3rym68rMPBUeMGi7NLFkhXzZuLAZFiEJq/nC/cIw/TJWi7N6Lwb
jXXXRDL6spvO7nSXG0Dzio2TI5AcM2t8HqO5w+p2/kfZsbAQoJ8dLKhYbcEZ
Dt0q/R5hHX6HWmn0XUDji/WMLQ+s33TB1k0pbozK+BHGidC8gJyRXRkWJMrk
tUX7wzTq9Fb2hohMPLtvn0sspaaEf6FWO5lzv+FWy0RdhOSmqso0HUJZ+Pla
cuIC7vzrX8q23c4pRJLYzWJPEDHlQw3NPVYuAjwbHIvF49YteLzjWsiT8+kD
1dQqN9Qyg8l+bhxvUn/WyuHxdu02BD/qvRMn2TrxQTSELb1ZiMOUFpI4TA+G
Y9JNoNLm8XSIG4VWNl5enx1Jr8gX+isKiAUhRTgmkDPdGo9dOGDJEbGA//J+
LcweGkt3EBt2vYyCf40eqHA3D3orR0UIClWc3iNleZudqEA+BYqiqoq5I4xU
oexeTrHOLsmAaXawFX1A3s8gvJmrFFRnkQybaYc7P7ePC/pImVe2blx+Cro9
af0AFO/lNBln1nmc8X8xXNIKdyJoy3ZLrXfqLjDdP61uTMSiobEgjQg3PHv+
tXT3eYrydkvjizY3ZDbJHZk6GK92t9uYa7tjxEc5MDHPUTr/bY+UIDtwu5mJ
eXIbOY62VW7AlJWioTku1a/G48JLYXmC0ngCJOebrc/OqPY9LWAcr9apC0vG
7zoy3ks/e4I7dVNH3EyG5BmNj7EcBjdVF148Vzr/LaVh99JAJQxMWbGApeU+
W4+Fl1V9oqjiouywvg8ZTovyuhoycEJK4J7AB8x7Vlht0D6MaanPitrQQulG
3L6n0LF1HcfFi2TljQYisDC9aoJ0JN7U6/4rJvfcMxPSox4bko1qSHTdVJz2
ptSjYJM/HMUcfH8tT0YGTPS9q2mshO9iIO4KFW/SQyFVNL5We+gwBpdhKpJp
Sleg6hbguZV33hd/mDV915mc6gQSDtO3FJvS/z1tagNsyeJtJsUpP75dnmQR
WDqrvOHGzfEvNUNptuDvsrL5cIQz2pN3U3BROIjl6LpZWx+Dbo8qRLephJrm
wadF9AZs0vIEY7olTRrfvGHRW9VsrktLeXu07gGTqum5yKw2oWpwNNy6K433
H6JgX21fGHwINPw4N9UjGATwcFpeWMnKTD+Y5GWpKzi63X+TmEQyg2ShQpQY
C5QEOdjZRjOJSl5JLbf7/osbGyWgZMRVzC3G/n3Nyzd/7MYF16cc6qR57rrU
lGWzuFXlhSvKe08WLF/pv0ZWSD7X+IZanH+IgZWnGEb0XIJrn+mw6iwTxWUd
JW4FkWIu9bxgCCtXsTyi9LTpyuGgSo1bFtbX7oVkSqTLLY6D0btAgXnD1Hol
0lyTXnzQpmL4i0d2L6xwKHhgpaIfqRtqoKj214OT+fnLBeX+k9SJn4lMTfYL
UkP/LUxcwL4gStQ10yAnQmcBMxfU13FF428cNeeQ268oFB2PH/HEOVhGxiSr
C502gmuGVtYtozNw1tUg85/xU7SxqZrBn06N33yQZDDQl4pjzJAJeoAQHkFW
TklK7MWSlfnYFauw3iD87Foi1Sw0YkDMf2LauV85bc5xlta6oxNXUZACsWbQ
5NVGZcjCk4wl8i7xgqWgkMckt1hRGm2n6NLgn8uwlNCCFhi97xC9Uk5zegHv
yRzF0J8nT0rS4EW3nuKZZHekSgSfj4gogNKU0GrE2OfTskX6eS1av0/qRK8X
hQeju4E8PxrA7fCW2VlM21Q6t1sQtc01sRTGenYt+UDAwu+8GrjXtGC6RB0Z
eg+kFELGAaE4+wCks8OOZ+wCZ2qn8Zx/xjz53ej8cMrd9/PTElBXRMwnblr8
WHcvnKfFjuzima9pw9NXOgKDC2F8ISbK1qaKFCL8dvhpTxS7uOIr2+/KSVuJ
9sdZbyfQ0YfXmBeq0kuv2BANmZOnc89OVrYivVnCTuzXCZYIrVjNz8nMj6yP
+k5+jIRUw0Hi/3xRi9RP5YYJCefkn1peLmBnmBe9ySQIAqOtBSV6e7MIJHUD
H7O+4D+t2DRmaTWA86qwWm8U0klPgK9xn9Z/kMpaxAra4krQvC9Um1F8SLe+
j1V+X9p3NmBp4bHH9Ojm6RdVkichHcx3SAxV/n8Q/KLqQF43BV1vuG/yO8IJ
jXtuMr3MC+1OpJawPu2+qdJymyh+a9VywTbZ17X2dcRpnL7s/l+uhuiFW5cT
+ZxqL97Q2eGZ9nTQNMCGaDolwPByXxCKbN3pMLMRj7x2o9smShm9CCsHaALl
RkzrbjbHzm9MKNJ3BM11ydfJ9UgBfskO43+5S3ctVzGUAXsFfFUHxvGA7jxD
GjEXVyRn3Cxhn4VBhuEj1zUg06edHZs5ylUTynpt+VzAnyMc0tDkcT3Oe6JF
yfzQzcC/g7QJi9hfdTrpYkULqeQojA4WUD5cJL2Ox3X1Q0lDx1D5w9BOeTS8
u7nLWGOSYegln0pX9xI9g6Kg1WvuWDBPneFHEP0Ya11eyRlqEz4aB0ra4eE8
rRNYyPwgeWA3JlDNVIEM8RZRcX4Cch8Pg4e1Zzy+PlpijwjloCNSwpylyryZ
i5WIU+CQ03LskQZCrE7ypqjFkUidesg3CpD3J4gEVidGYc3PY83m1+w1duP/
ePLyjw5FME8oeRyCwG91uUOLuktNf6iOaAeyNYICXaAdYO61hyUNTB6jQ1/X
MKxTiCb4izoX468pO7FDwe6M2hB8ovNNhqqTt0SKiuIwj+731RBLepYq8mci
CH8oyfxDRwS9kyN4svgqJavOia6yxO2KzNtp6wOo0fEJZ/tgcPDcbxuJteNw
4m66FW1zJEpPKdlDkfIGxM6s4ouOdFRkHUbx5s/v3u9653CoRLr0cychy5JG
luFPbnJYXtRc7vWBVU/xHQw2OLKKO6OsOQCFSj2gNzKvqKsaEwn2b9nEu8m8
GR4Yi4tiqAuGG9D4TkRtBUJmSWZoesJ1usn3iwuVPE9HesU6h2KhOHl0fBb6
weewlIU0ABe/rKIpocGqsugmESOlA7yw1xxWpySC8lQzlJMcKXYB8qihOOzd
/MPF6OVwYnPebH2QuNxF/5YkC2+VhgaX4pv+oIBnx3r4CMYXTdmMRiNcRbgh
16oJz3y2O+zlDVcBpuEfSXCNxJh1QfBZJeX1ut+1QFWHLDHk0An0NFosZjFZ
unXYbVvw6LhAVarhcqNyS83KckVbNOD+kV3Fw4S3MNnat7/AncGmLBwqIn99
camv5btGrd+ssNKsKJNtnwPYvCgpf3zDzvi1X/J7UGfWt8zl4aj9kNf50maY
jPIJbIkeLGvKccpeHNze9FmJ/JPaFUbneXQ2+dY7ZNzpU2G3KJ8a5tr6m0fH
VIv9PRgxd7ZJHm4eDc4TIKdxTjzNf172+OHdRQYDK6LCHql1TRShE1AJRiWw
3kScNSYlG4xBESYtlqKsf3bMxbeVHqU///WXj2JXqIKoTZmKZtgjvXrp5FT9
E/hoiX7KaBUZYdv4ur9DAKdGxED51K9nm3ODhXoPLtbWv57faULaCO7hg3mM
ck8dJgxCgQscFv/CP7sIWMYAITuii9d0BLgfkPqt0pLBBzj3clOO+koDSZp5
jXyi90JwJ2uyUmyqVg2mYjoxqxZihchI5EWc3KRc84SRrXHfAZrOia4/tPkw
gngyihpKVNUb9LPgAqT+x2tKthyNdjhHUFciYrftC0dSJxGi39aW8A0JWUwK
/FhdwVcZ58gJcAId/l6QpGhcIUiB4P1OE45xRGht6kLNohHa4HnngEeQ1XKJ
FLETD4F4qJMU6ThjS1E8BpYSbraHtlV3WsePK+1NOLzOeyaBdaDvDyiqpau3
mW4N1ld3niPCc7S7gyroSp+9RK9tgbpJNSmWVJ5i7KTXsiKPm3GAgbFZvO43
nGJvl84GxTJOSJ9CPAuWkfzvwloyhLuPtM+8WVS4nKFjolaV+o1casYASp4Y
8Gd8oAsNg8wDcqT4eqTTzi3ECVwURg/QxCT8WI19QewZ6Z+wx6vlQ/9k/Fzc
pimVB1CDD2vZpAft8A5uiK9EhVjicEYd2XJL43NSKm80fGhLnS3px8lYI2Al
kqEieJSh08ngWLOE8F9G2S5Ntz7IQe/7PbX8o6vVOAwtGU3DZyljAE9MVcvP
QOwGNAm3oTtBMEvFYwPiuOphLCkiQ44qTRjULk/Z8X2JgXG3Wus8wh0MQGsk
K8mi5uf57RrYp8mgAh3Oya0y+X0tpbbkoxqet74cVAxs1D802mumiLixFUQK
l5hoVxGVF57bDjXzM3mAcio5NNNdR+iitrS4yHfO+wsIvMIbc7wqQ+88vRTa
WY2M3XN7wmWVulKxRbJaXl48Za1Ofd1YjYGfg/Ypf2hhbRsHT25G0CzeWiu3
LSox8STUDNeEmlh+Yesv3GCLvnjSskNhMKlPk0LxlYdbSRwXjsjGV9zWdomc
0QgoMI1RcGeJYWljxhmWO2+08Z5rTOUrbZWoOQZkUwpkON2Lk7WlqeGyHlBm
b7vMHuTcGjCErXOIuJWhDW6uNFci52/LKyf77qGSI113CGtTH2Na5K/ZoQVg
YL3UUA4JgyJkfgFjHyOYtf552ijITtx0dhWvFut1cn2Tt4ZD8Xxsr3szSslB
UcmmxrP7Ndt2+w6D0ZaLwX5yf7FbHL7Kk/Ja9S7JlRY4x5tlL9q3pHlQHFOt
/5WFbr/ZeTiwLBAii1Ovspjj+T23bAjOLwbJtD8BIOfYAKXdtsSyLSFDkjBP
eJMUKSlPLDfgC7MPwfwk6mIG/YUTFUedUyTztYOvTbBZPpd+3m8xdpwxUxJT
BoRIvQWRlkBbYTD+yuaC7ewMxPjOP4eUUDnsnDq+EtyGLX1HgHAzxi1dPdPZ
hL7KpBST9zLVRmeXQzZx9PJ2xZXUU5xk+5BGdhJ6LxlQDvqUkR9xSk5iQW4S
YWGdcwVYJtWP6aBHbCnemrF0RKExDU2hz0uN4uhEGZH2bLL0DL9Dq181dLVV
U9ysUk7oQV2FX0/y41ypPCn8l2V1OKRkMBBUNDBloIDYHzMiv1uLRu62TlDP
7qhtdU1TE6r7GjbphDPxwoh256XTp50/ZBZTMbvF7FK6acj0AKpeZYTWhNb1
C+tjhz1hlRWCbxl0z3TQFthmFD3dOXCu1bPVkQ1vaVMszK6CUHfyvPf0Sl8G
/NXlrRi+q/dn0nWxJg6DdAq/r0fh1mlTvJaWM51bGx7HDozOyOA+cMqRiYoW
qwM+quhCYlYtJ2F6/WGCmgXx/w4CDTeS9zFXvDN+JBHhGcAWQ4I7oJaaUMEC
hnCLQ/epKGe+PsRXrGN+RzpJR+g2V8elYtxzzO94Nl8viCzJIZRaaNpc6HzI
4+YPhrhmhhpMHowCYurK8VAXTixtymYSuDnATB2ye7Agnsqqu9HPh9cjEwDy
a1jC6b8usABVl4+LuBxG51WAl1KX5fI28osS7nm1xoKDM7StvK/oVPS+DblX
3D0ymp0W0sLMNVHM19Z7Tw8FS/xAAFIWIx+3+2GpWDIRwK2B8jKIu/VkgmCR
jViz+4VbxMjur9HAO7A/UlsCYG5gCQxgg5v2gm8zUP9kVhI8AhYSpZBlGeGk
q+t13EU/8UXOej/XP4a/LlT+qpdICTKeGjztd4Hi2OrdF5NxxJNj0bYtLavz
sSIKODnWuLFDeNPoYJkB2riC/zcKqYH01WcUW0rpuKzBTK31tgMBV1572UMP
VCeu07YP0grZy09ZtIIB5dwTzVvtqN40c/JCMRr1EjJoUZgD2gmSoQYWP7OF
YQaRne4Wl9FaeVrgJ71viMjF7WMjLVmgPlLFycL3Y5DygR4/NGS3PSdbYbrC
koDT7g0RwmHUOiPsRLZE9LTalKfYdAmpa5sSzED+sTSUx6XCyqWJryTGvdbk
Hnw1k4sSzv4CmYXXIcoIioJ70KBf/Qr0j8S0OMg/iHlxE60ZbnuGCek7dCol
gRuMtDAE22MDs7Hm3CGzZoVY0178qLkU34b8NXfFDvHei9mqELFYXV0xvczr
KI1LXz487qPHaMu5W4bsZHzx5VgQL8DITBu8Dej3pDA4eGOKd75hUyMGjXYs
3ehMuW6xvTdmrqoBgBKkYYlyjFAcDYuYksoj7r+63tWZQHI/3toCq1nofFUv
wGz1fqbJw93L78h30OvDhFA6Ladhd3rAOqM7v3ihrOjWNS60X8MbjrszCqga
dqx4psIkhjHK5MMRdSGUDOpaEDEbb41AxKTqyZE+PAnuyUtZucl+wCq8K86A
CyJ7ycBtS1HLu53Db+vdHDeHzGUIqfgC0kofjkFiupWK5649tWy03vwe502+
ewTK763NgRG3iCpWoiO4REltX74wcik9H+rmbz516OAJdVX5Rqfah+/1R84U
ZxQ/UKVoUtYxSf5Yt318ngDRm0pf3c5dK1WlAeEPUrpm/lPssBosH7XMq9UA
D91f38t4K+0B1yTIKCjIhAnkexbfMB229s9oAb3jI1NSQ4BC7eFfGW7qrUVi
p3w/L0qsJXsIwjsB/1TmN5Nz0onq1mVDkeDe+R4urPh7W+x6MDC6xdw/zTuE
2VtaTpLfdxBAwPyO3kY8mvD/csjhMV/vy3hDNYy6Z0gsTOG36PAk/0wifarL
wrzpylJPpfFFuERvblywkq0dk2QnfjBkp0wNILI8SvEBvrmw2yKfSEauTx4R
eh6HwX+dtNyXNlPv0SKcnLaIhqpupXrHOHwDuMScbmJh4LAYN+Tuwl2x/3Y4
vvgprZ/9nm7OBM6gxdEooAfWHqpPiB7L+HRyeoyEM7gcnnzrYFoZCKcSzhQS
w//umXLUG54PSml4wEBXneBW0EoaVvH5B8fa4YRHsuX0UYdxIi8KxqpK1CB8
mPjhzidCrw3LbtQX6u64oh4oY66xththoePe+Tq6Ng30ffvcJemYVJS7o+ol
j+SAtmbwX1UjMd4Fe7dJIqHj3KUf0uVmjXjssQx72hIQyh+DaNMQssdrMVfv
bdCFOeBCuw6FIvFS6KMWIOCY0ufry78OoxWq+FolbfIDzgdWNu+xf6Ww1x/+
JWI2+3k6jKsQbVrhA6f7UL68ce6M+Qht2NfOC8+ssKYNFll6WD940icExAma
oQ9UT+0refmlE3EXKS3Pe+medKGeVLgzQbr2meB/xLUSvuMN3XxyrtIuE7Ph
ZilWd5GiEjI+hhxWXtjd3Fe2LECbIuU/vhJE4Hdc1GhfmPQ7bawvSVE6/z0l
GIXjUzOOkC/5qzltkx+uLEKcQxDnEAQhGAlQHZicks5/cYrGsmjXMUkfDQL8
gr+FbMi7oUMs8Ss9vfOV4cSInJizvSY85XOGKLndVgYJs7day1F+nn/ice46
9H8bXqbmyZqm/MB0AyMkEXozHOvFNqLUyhNlp3jTPyWK8ZPWb0SkTDXjv4lp
8reQRj5WVNRUA3yEE0iq2vOCW54zlYjfWd85ni02NPHwc2K4lH1aMV+hxDbU
EMTaHUjadowxecRbUlA4aj5tkNuD/VHn/5sEA9lJgKCdNn769zUd3w2ojiLq
ncssioA7ejjj0817yEJ94zpR3sQXp8i2/PSziDSMFJwjIPdYqpT5TLd44Kxa
oZl7Jg17b5ON6vvF9s/GxSBBny/95udi3ozbQIszHtXUepvmK1xuc07V0vtz
ZleLP8hdgcZng+DtSznUCaO47Lk6hKeoehQTrKQqbOczWyyPVdXL4CBlRJrB
kFK/dYigyA7KPt5tBZBMQnUhUVAlTZZImyNKSoZ5aQ6MMKIVMeAUxUyf4xIu
VvTAwhXmrteyMwsz8NF0bznH90lDkjYvzDGGTkssjj9sb+xhcdXUfYQswkh1
5q0W+Rew1kAgAGstTP5hFKILD4UDEPJMLBHvAFBPbwxLxAdeKFVX/AJ6MJc2
jjhnssLhOzd3ghJnVtgBkhXUJWAfNjOwajWNUeR0NIMphR4Z/3rH+ZlphNb5
88OTJB9OmfzO8AJXviuoKOMIFpbyTwgDTv1JMWuefC91AzWzGyF7UCf7QzKF
ep3fbLLwC2w4wIsSeRw+fCY7Nnya4tTv9pH0q1RqAXEnlEfWsCfpbp0cogvF
Ti56CBl+PS5tdIWbbtI7/0Mpb+8jiIl5kE1sOrbQfs4JWg8QzklhjYcRyTi/
3viZJNY3+6spiQDHXEIgj6H9BJGOG2r9QOklqA6gsj5bvC0jzYqK47U5dxLb
6TQBa9/mWejCYDV0N8Mua6odShHM3XofRfHAeqaFjWBMMYaT2K8ae5U+pycW
JKP7KmVoaIrm1BOHdBCuRUEvSfO8LE+HSdb9niBj4xub6xpVuokNnfbw26a0
2q4yPKEMp9y/0gs4BxYzdEgNjBXsRgFh5MjXJUhtLJoOdbUb6sxj3RO3kbEa
2pAyXFfmt1Orop7lBMITl6PnXIrLpvuxHjzzHyyR00QXbD1JER+GUngK81FM
IGVPvFZ8M9q0XIM3IZYd3sJS6Sr2COBn/RKRu3hVcz+m2h/ECOleoN1xH/QX
J54Y1OQl/mrxqw5T1K+VtzF7tKJ+Jg16vmWkR9GMuwnyEtKKTVg4QG7rEnt5
bbMWJxkrO46vmNJIms4aCkwrK/lZp2xfwn61io/LG+8rzn/mhX/4DMRkEtBu
HAOVrNo950IoZ3TS+DXHBjG7WlFuzaV73nu0GNj/g4GE2cRG+FNlbJde7sTy
Bf4JxqME6gUjC/E5cM2SygFtWvkT1NEHpZS3gNHeg6na+9PqeOWv+5senm+f
XXvLHBXdINbfkuu8OFU4lkjEGYabjfePkCPElJo+ln9M9/HpGeLDdC61IeRV
Pys1Ril+lYJ1evRZsuhB0J4RP6br/le3G7dVTTao6pAqYtzt6OEBVSUxkncA
p/FOwOj0aq6rE2c5slXapJdJZR1+YQJmGnFbKYsJNcY9B6fh8a0Rd1ITk8ux
r98Kqluegx8ke5ZqjOShu10XQb6fpGVo9ygox4VO9uVZpgJ/HK+A7aMaupdQ
f0r/cVeZ25AJbkGjZ1GB581WKU9s7ce6s8Fbva1Un/RYffHf8QYahYGtikUP
pfUELL+/bnZJ4oAV3YJ4xnYeL3Md+m4cVLo06R5zDTVFrWMMytNTUfYXf6JO
k3VL/tUQ6tZt4tdKCp6d+EFNqWtwCOBoaeNbmNDu0uKq6ncDDfrJpJnoAtom
g7j5trhPZfbrRPTYQup6sAHucQyJr6vYceVABCbptuqNr2UvA8ggz9FUWbcG
Ggy/pzb2gH0sh9uURyzWqeTx+K6frxkUTgXYWjFnw9XT8Z5UN8Za5vD13U8B
ze+dP8sTWRVTDxoXEPQHT/H0JAoCqeMaEjXZIqGd4u6iqHIxQpXyRsfaqPlY
IO99qDIf5Aa5TXeVWoWfePgq4PDQHC6npCQathu6Azn51egznAycn+anYOEF
uPkF1z0+xzlkUFiYr5FiWu9lpAldX+5aRP/nxzy9izbCQQd98eiPjm0136As
YBRFzUN8gp55IlDeWIfpmtcpcFruifbC+4eeGoQQ90GhCSmtHYL4vYedy7M8
UA5b1qS/mn+eQN6hwADdh2/AtEx0uzWwP+whLW4GGA0F//F6ltFU3obIJBSB
Tnz/xUpWzkoiBj+74QqKdwhIqbDTT4I52m2CyNVWKbfPi1skZWelH1pfvUmK
Kc1PZAp0GkS8EotpkEvOO6uYKWMVek6BnNHcUhM1Mv0hA91FX7tZ1nL0frry
3idJPVS6iFBC8QgdGPKZ2NbEH/LpWPlo5Bdh1V3zDNO8gr/31h3jMZs82JLG
4dtcD8DG/jiEdeA8DdHbIaTVz0oNMHcZ8H/Si1rIxXnhfcQAKbO5EMkRM3hD
qIMu3CI12NDl1Nj0nIJBl42TTzyFUt0tsbr/SBcBPysiZ9T8JjhdiGmcDRnP
SE9sQv3v1pMSFzJc7PBb0pQul1LEkWDH9idLdXvS+p9X0vuqZYKXSqYchG2N
jv+nDaPCao/jwzhUEHHDauNGKOJg0TPY1LLrpElwYiXuKriCDvmTdzkl/lW6
IZfuV8dxgqQg2AfWK8NRLdXLwNCykg1bFLjXUgAXcQyGHf89Ev3XubgPuQh3
Tkm7YmcU4//fCy5Zx3LtjyeIZAgU0cupGeHMz1Pt5jbR+E2d4F9zj4TIna8d
BXh5cAXTI3aB3z8AvlICZsbzdMJooxiDImvfsaEyJnZi73fyGHnBcq215vsJ
jxRyXml4U7uYunugH5gB8kIK744nvkpOmePPtTxU7msPxT/MCq0FZ7EwqRi3
bEYITmH+Ei+VOxQwo2izQEuKiY0a9mPBPPYdt0C2aHIcTTYZ1FbLqLLlM7yF
tl9dSDKSBYrttObxs9nBWqA+2ZXW4BIuKPh57+IlTU6RiJrcPhzZXfEPxuXS
grxvPzGInCiD3P+Ve2tehM8eY8wrpl/KmojIay5HZwvcvAr+3HmCG1F6lP/3
3C1i0dbohLZc6bYbiFLnlrdI8x+QTdcSEd8+hSm6XM+V1iPC7wzhVWQtOHsE
y5eQuZs2LBaDkLJyGbKYo5L1ROU46irUVMDJ7zDIHsGenyODCgaRXBZagcsI
ynKBw/+cmQvtLNk9D0qZ9hoSlxwS/369SeN7hAP/YjQjEIFOMJUKQ9Iws3d1
7L0/b+Sjmu2qig9gseRMTos4JBZd0set88DA+bTuE0SZW0v/Ya6e7y6O4j3A
IQXlXONO2Ku3XxhUsOZ++vS3zlOyPNhM68P6jLmCrw3Q0JNPHTpcFYEe9cOf
ljStNZeNPWBruaKbzm8QEfLF5SD2GhK/UrViZia4rVJRFCpPwASEeyNn5MAE
7Bkdgp2O/Ok31a/Ppi1ofto5+58Ih2FMRn6A54oTkHatBzHwO37J669oSIk3
unC9EdNc83gCsdmuwoC3QIqd2gAYfoWgizhuHZeN4/1UVC+onwJ6LQ88D4RZ
LG4kDtevC6WPSgx+eCqgTvp882oc45UtNMKUm3vbXrkMLW9YZWEAZ6eqNktz
XdSYJXHOQL3zsygsE0p3JhTl8/LB13vfoAi4cYt3GsmHIkXn8Cv/UJcbwMaJ
QIjIqr8M5TW9SeHAaPOaDgmgy3r72iYWA87Q/DotfFR38gjQb3iWr68aP1Wz
UGqTZ27WPfEtkgzRExBiaRkbqeOd11PqK9qa/h3U7LZIxTpcpQjyefMSHNcN
63/eN54+NjeQuVrh3HJRZyea3CRAZSmxvTsjSug/bI+shxl+LXxDybsD6lo6
MqqVL4sNqJcR1CKeM68a3pYPCa7iXpGk3gHG/B6RJ/iRqt8rUMjAVwfVZuNg
CIRk0hKmeCkpPH9pE5LMFAyiZ23NVxf7M/2mLRCrpZ+XqN5c1eGYxp9z67Ah
dUl0FSQq/phcto3XM0yqAnJA28OIygmqvPIABIp+udzll+bu3Wge3TfoQwHw
GUipVXEhL4U5rT6Ysp8hjHuvApb0Fmwqhstn7zsH4RmReeIzyuP5XWOLsz1M
g64xy+3ydD6DzePEhaotB9qFKHmb22ZjQxiFqYS1GOsuIIOC41xJqdRsY2VE
zFnFD4ioJD524+xwIKueiB6tIAyBsvtGJ+bXrkmGPwnHVc6c9xwpEju6zPmB
1aa5y9X/zMSPDzDv4XZQaVXihiCVdfJ4alcwqshKjOFqo0QixayQLfI5DqCx
WBFNDw887XA9EFF18dSjAvnIKc3J035BAMeMGEYbUxG2lJswxatzENVsUzsL
98KWSiSYIt+OGYyPrDzpyhP+kwtkgsvC0UgiQdYtbr0Ey5TbAMKMyGOLMZ8u
/CpUnwskschZacyECtG9XSRKhXf6DOdKbKwrr7Cvbehzv14tCp8j36k2+qTt
rX/1sfPUEFO/DIQhhZzwMfD3IINc9F9WBiiKOk0DRddqCs2YXKIMUqW7uBWc
cgotwWgJw+MUY+HD9tBLyb5jf5dbH2Ll7IQUei3/waNcrMDOfOGlJcvDbQE7
vYWrZkEq9OqmU7rmRrD/XEznnuuVC0oDloFel6CsL0Cep8QMS3Y7zBK1gDam
ZiGR2M2vLfy/AI3VRRfHAE58v1Hmh6p/pvpwpJe4JgpUTxkoUVF4dbfNLYE0
AoNI2H8m53faRqvrWusPoG154C83w1+Z0jMdsd+kU3IDi/voX4pbtRGVa/wT
8+PKFxzPQLCO7PoXcu2W6AwMmoMnPBANTsprByfsZvAWO7DBkIqauQaPT5aV
Nr/6HKkvqPPNquP18IQRlbopoX5Aec7clHytBUKPLlDQ2slYjR5GA7CWu6Qh
4BWRLRASDLc0grw3NxeqQ9+3F807kzDZW8OlL+SuokxByevAycp+X4IC3DBc
riEOpWQrpVJfv7f2u9GsjvsXFF7jNz1q76gRKbtGeqkkd4cqPy2f1DeG6gs4
IwOEWvapy26s2vVBUVmB1STWQY9m6hVS3Z2ZY9qTUi1X3ymtmVYHfHncaw1l
dHIxAzh44vfpB8Mvowir+H+H78VYn9BmnjIXVPDMbhJMyOB7ZuyxZBnyoCgD
/cr5ziIbeIi2uUr9mNIZc7cjU45arBEDBnfn6bXNecvVkVetkJY14daqq2A0
EQ5bFL1w/4ZqJ6wbWA9A2NtvfynDOei/7tMrCw9RDhD5TmaZNNGZXTwcwwsS
DGRCLj4NaUSpdmZJDU1/BaUP/FcHYbAelOWwn3dGngA7QALzjTJwAjbHcezH
YH+646Vorx4raSNKtwPt+hSa56Lh5yNO49tgoEwoUzbUBkEM1voY7ofu69XN
YRhjEEv7PXf1bEVIo/hCHxWqVJ2lr7W7J6vWQaRhFeaGzw+H7D5uT5DJF5Hq
NrQZWhDO6zYLiMzLQlgbl8m4Y/E6bTUO3qix0AcBANlPJAt+DYxigoRlFcy3
U5sRMnqDAkp8g6eAz1s6gYcX0ZKtUBnu73isNmKQmnjR7Ld6cMFUkFOVS4l/
DRJSQwMVG+erRp/J5DVhSRCH/AZK3vjMQb2m2HVsyoxv8JnXn2G6ehdpSQ9I
M3X4CdFRwch9gzQux4OCc6BbTg601g5gQ8X4QnKu39nuQa+MXmtBMJofNQXY
6zDDpOKr41FsJHBS/Kbl5k6XVDzzAF7MEh7b34GtvW1VY5FG6t8IcFDDDpME
RTCoKeDzC1hZJczEPvCrurD7WoFOC1SYFJR3SQu2DOiPCOL14+dkPLklrpK/
27/oWSjOFhQZl5cIMZiA/XDiW5RfbvNKH3vEP266zONX9dzc9P22u3iXdtg3
AtTKbbEWf8HrEtOOjHFAOioxTkIGTGSeJzJcDJm2kYhs/uuQti7XmZCzYwxF
1vKZ/IjsH4lovZH4EjuH1bOdExIl6OsLXgf+Uzjb3EyPGkonQ9wZs6+1/USl
ecyOPBA7+JkoNpFBM4I4xgwomfFPLm1yXyTrq5QdOX2fe7vcQIp5CHgORAqK
yBeZprM8EoxBU8DNtz9eS5unGx8aJcVzSQTC+yEmfmdwmSxEBJELtr5K2BH4
WYk/rkBJgf4KMIKqdMd4cm3SkgSCzpg3aUb2acts08HcnkOFpGn4gajk2uJX
f/8VoN01nXdgMkVg7H9APMA62MpZsVgnQsrRM7sLow3Y/flyJ8MQtuBqOqda
JVLaGK4i8a4PsVPmDMp+ji8AmDNCJR2UmCjixsnRjMfoq9JxYRh/ihj3TVCN
NkOC6vYMSSBfk/3hmDXuJjQfE71Pksn47mBifFncmQrDEgwf/jY+xZodclZK
lE8BopSa7Jzmm8uqvzA18L1bO9hfGqQaj9ORjQMuoiAyoRhZ99gUcAPm955p
1dCQylW2hHPjw/3PBaaS2k3w1Bcj7dAsc629oyszh/BUuIrWwCTzYBMVmjt3
4uCiEZoOqDogZy/gv0CdAGVED7IiItUOP/rStE0lvB7a+FBU6PksA3tSXEvH
bY0BCd51KPFd2CSKbSCIwYg0FhoT+f8lFNftWdXB2UgPf+a+JNqr2Km9Q8In
2UCwuQqH6HgrGk8tfXaRLHDsb/YPbBo5mDaJmSRK7VeDI0i2N0WZ4g+RdnEc
GPKomtuCNH92Jza3EuG/H+QVIit9hUI5JqfLdVOXzkgbL7FvpEqlheV5dNur
N4yiyoCi1zjZkRg+k+dKWvE9EiBQUNoYk2ascZMawPWfm6NANwC3hx4hNR54
LhcF/e5TXFY+l20foslYaf927JZp178kaGBJ44+56AvzaE84cAFjdXak2ovX
g8t9DoRtIV/bcpooc/6EoCDPekgEIbEJ1Ui2JD88kZKj26HLJ6D1QO1lVpDC
Kg1dOCdO4QDgJfygDBAxl7jkAAw/Uh/MR1qcus0P8QnZPQ3WliWri/S9AZiw
bHfOY3iFK6ub6ZBBzEmuSNANoCrIx9uIdElyelihtZ8D0TNH5foERzkXYujf
FVqILPcuQg3TAHGt/6uo2f74HAEaXK/Wuj+ANnrU2t6Sc2dnLbDlDDYMcAwc
d5/WayqhDU+iwzBpFONHNx3CdPHKh/veaa6VYuiFOi0NzII/ijLySYwjEjn+
TlX3KgsNM6TCQMtcGNHvpjGoGd3S625+e5uzwlfo9+jPCJjm54AoaQ3GoLEj
+wrf2PI6hOaoI3rzy//Bp5m1fNM9k0uDXhtdADUWo2HHXIVXC8K5h2Ij2lRT
QvJvpGiRkOWnURAkeU/vUisUgWDXOfBO5Po2h82Q3SNn7ajXGBIPNI3eJKih
vZguZsK4FyI8pi4S6IT05HKqbLa6/5a3Xuv7qPZ1xbGc2erlSyv+NIHV1DhQ
WcevCUsz0E6f5Rosx5nAQEOIzz15hCdCEJVb1aTmlEUFrzGgXWeyuiPkgdaY
sewAt00Db6h3JlJIjTda8p+RNEWRKr9jN5Pq+QQRc9fkfbYqJGX2VOveWKqz
aTCe0byQJPGwpBv0cRp42yWNGw+cWnmzTsvpMtKI/aRHy00g10b+anr1SalU
sEgy3fLjFNClsJUmY/PBGKzw0aeI7Ex5AIOircAkm6qHqTbyW6gxP1nf6plz
GJ//fqVcunqD7JuiWSsdt49vQ2qnzAFEOevZasdwyDwMi7PF9XehwIhU6zuj
TpR6lTOO/PxvZb1pYhJ5yXWvBQjwmUoe+28EIbVc0cAU0Xmm62MsYc55Qaai
thZ7DgEeEsJutldBOBkAyFw60Q12WN8bL+DB3MXLR9/e+qhQBSba2UP/ghIS
IUk/eWyOf87xuJfAEatm1sN7vCL3jq+I2mwrc8iebWkxiWGejltsrAf5vFn5
HJI/WgMdtjf5wddJVKIqw1btn2XH6Q6de0pkh4sVjmeCB1bXilcvNO1HS01E
Wh1CYSrpDrvQ52Drx1w+fyQ3LF+snmvzMWPUklKkORRvAg0JE4RPLeH/aa48
By32PD+pddwp0+SpZ1RFgETCZ8v4LzDVIHCgeqt68DBCw4FAwjHqi1fFtBWl
yb0QPYtfPXiawNeg13Iw2LA0OTImD+qx8jXhXKNPG0Qzona54yB5Y/+FRNGw
QVaLKH+18MDzn+rq5ldyyh5G5/17+mg/dEjPT8UAS9Tban4hRx+WWdLf/2LR
BX2di01Le4amHPs+ZZ31WrpzCiluMyxQ2Ta5S8LrOz+E3VdNohrzL8Ls79ve
qMXpg9jXRa/siyZkx7cxCIV2LzrvYtp4xIq217ifr3+PvO3H9X5b8XxnSxeq
g3DetuiSo2jQXDm93EAJ0LUBEI3RzTc989qKlJfYEG+UcJcXjxr+Bg0BII35
cEvg0PGzV9OcXfxC65esLJ4jNJPTas+kbLuU8kP6mkAQY4Q7aAzt/j1orwiQ
l/wUEnsF4eVeJuk3dMNmLzAizWxws3vdpIGVu0WaPWZEDV3HItjmss6XCHWA
gWQD/JIRfQreFJPAb3jgXplYHMxiIVTiKRasVG4+zvMd1zZ4TP45ra0udmJY
T0sbhiBY49uzFDq9tNkQl/n8qYF7XzPnwUy4GrvMorBRUc8yAjC/FedmSOlo
r2s0DR44xt1cx2bYm9JIt2XcgPRfTg560JyDQ/CWrP1yqGY1/oNQcZKyumUL
SluB2GYBK+mPRZmFa6IK/e1ITsCJl6GXnS7S2DDiqx33emTYNsQ3sF14IeIi
WVlyyN4AMXR3D408OpCqK65XM148U3zPjYyvv/Q/LVPhQucwi/UQFJ3WjESc
gUSHqhPR3eyOR9q7iHTqHBtTgpCCZMEXDXl0rhu7Ex7ONBfmwsZO1F0x1Bk/
HpBNIdaEEiJsmUKeFC4ZeFtCy7WJhS+zDy6AT/R2YXrWZHbYPtW5C3W2TqZ/
9ndoAkQss0Fv+U64njc6qcDrks0lW/YTVHsEnGq9aF7ckCbarB8EKF/k5ZkX
BEsqEMQK1i40nJ9zdA10i/kFqErCvXhhMF8hT50etiTZ4jeyNLc5xZFqwvuD
Sg09S1uP66Nl1a5JeWe7uo+wC6qODQIoJ8oumNxylH8EiOGHKJy645QPq/y/
1+eRW2RqWbGsqgHmchE/nje/T/GVtIm+N1iinAHd+9Pze2lyS/ITyzFaFIqA
AD13sMPpqAj4poqjEcom7yOItizIIiPS9wmr0Az+G+5S/NRxPJahSfK59GsU
ZohXiOfGiWykkKidDiSQWOP1WIzdZ9b7Hb9mYz+J3uJ6InT+T9umkE9o/8KE
POxlhgWeytLyW2ED0zZ5SmutjxxatEwboeTe/LU+/0pnf3a9y61wOaLmdI7G
y8VYZE8uJjArlwOswg+sf7+eosCNBAMIc0hPb7TpdNgMC720JCWqGotYdl5g
drRSRsfjNJ6L8HbvEIlamVWSFuwj+9H09uQ1PTfC2nZMIoQaP9nnkwZcrtKs
qOTU9leZTOiGo5jyy56q29uPM7/Nm/trxr5FMtqv5gZ7bRMegJIx+vqVaiw8
J41OJCXpifBemBEgh55muLG/EhNVji9F47Sjom6ECukACfERfLMyGeoKRhIv
546k8mqEuKKwDQvwETFnySt3SSWFSa4e2LTIICRSkZFR/ujJNqSr2rf+YDVJ
RbgvkeCVECWBPgrk1f2lfhrx7lQI5UgyybWlJtaDsC32o64oFsCOxEGQbqcI
898dQL0N86zqao516cwxLJxGCJZxwo60iJG//TQSnZZgYNkVFp05kGPZYYIW
vTz5rUTJW398hnUpIEzF7/9wAUWDrj1DyNqboOq1c+ynmf4Hk6gqyxoRVbpa
NqLgjzYDxZptvNzbjvCU71arCFaNRLVEFtfooqqXca69NZfpGOiWR7BKJmwd
uSkGVRQqX1EGHMxr+GyxVvoAY3iiEoZd/PBmcSVLA+XDekQE9S2ObE8GPfB4
r1nx01/iwWRWizCwjbVLqEaFJuANaZMvjgQs7r8JQbesYfdDVImgqhOsxK2p
aAnnhsGteRnyYdjhGd6fUtn6orWVj7Ki6BvC0STC120ATFu8DgwGadLUrdLa
BLT3HlYb3yrmR62meU7vrfby2b6pAYkgp93YVj78RFV195IVVEiBW+TikrB9
lsF2PR1dzTnwfpQa1UHg/Sg8OOz4JiO97tVCNoRhILGcPaSB1IzK6/D6oQQs
uxWEnaHWgbzTBieA3yS2drpqMM16RkwAQSFH6cSz7wcUc1DeyVo3j0Exf0AW
AXoxWlQc3YNhvFndOhyP3Q+jRSboCi68Q5cKVWt/LZlqeyU2ISfKWqmUHJUt
7G9uIU8PWHmJfzPQK1/s0pjPTtHR9D+o0zyx9WTwaoE734a5xGWFf2T17wwh
nut0c3on7DMflBGwiuRy2GvZ/EWTl2TJzyxrHjnX/Bqv3PAAoW6NzWLlJsse
RsO0i7FTCeAFChKto4mosYdsY2e9dobkFiRJU8tmGqEXtGBNeW0z9bKPA7YY
oYxVCnCwacrlRIvDqCnb3KzreX9lPcWlMnqqL1s7BYW/pp+K0oUv7qD1N9dO
uIjEGsLgtv0cfq48+J0ffGGuSTT6H35c8j+72zNVB5sF5+MtiV/Ifh+S3fcv
gNIZf8rk7R/1X+ptR4xy6Qc7kw6Dm+GpiX/Xk2aEqGZa1OXxYXof0syHVxHj
icvdjzddZdoFGb8aOcjb6vjK5CNVcve+59aUNkjcmd6v0kFp9LvyejpLvQss
6QIkvrWtVR0z/8xZynzmER1teYHz318pmITRYkAdbD8AikRfUWKo9qzelvkY
dDw4dVKrFoRRiOoPSER+U9dBLqKqsmWzqr/eROv6Y+2ByZNTVKyqMn2613EZ
/1qMRrOGuOXvOj/B3JhB/78E3n4dxYM3Ig7aECIa0mHPOL76W1NoZx1v9Jet
yATu6uedmVRIkKmDpgnuUqxZD1yUzaiOZvys0QEwRkmNlD0FZTWJBc81sW2a
qpPxqMo4Qd/t5Do8ui9fotb4jWkqEC9EFC5j6fHzYAm1T83akkbgCKvgPahC
G5Gysa31RW9vTPz4qg+SfmGmbFueMGmEzpxS5PNf08dGpP9QOHwBrpvo2MnW
J4jBOqIGHbBc2FSeBpBotqs/hkscD1lDDrBqy4I06eXsDsrtG5xSZCY2SG7O
RH4mDhiWBXdXG0/gZZiU7U86Cx2vxYJVcIWXICudEcKeZCR+l5Qyuj3y7fhF
20ia53albXDA7xAcIfPPxkr4ToI5H+xIrDDv8S/a2Aj0hqPz+r4v3Ah/pCZo
NAF/6aUhFmXAuRCsly51DbBYaNwpRd4lAMQor8AK6v6r80qeE52CoDhnrYCb
NWuQxXnjvhSudzNghnmTB/p95oNwjVVz+FVR/tsEPhQpVmRTOTTdmBhNLOT+
mkq8IxlK+SxHRyYBkTpLTShOWUJs1oDCG28pLHJBMfTNYngFDEpqrqLkFb2z
IWxNe/Y834NKE1BGW4OL03aIUrEhLy5D1qL64untc0v+HaCxXAbMP0T80FcC
aGuMvt4xlw4c5vqtM1q4V0BUJIgpzs42RbrIvmV+N6+MbY48V6scDJXJfFg6
+cBA7THbYnL4LJGe31QjFE33b8tQdtSv/Ih4ybxmKhXsHCo9LwiqKazWlbv6
OguObJ0p3QdV3rDedeKC90efPDzG60vi8nBi6SOWEKb0CVqW4FFr4dtjfUNY
rqlOzqcER9NGVhmMzQxSPJ8vrbzj3nbiornRifBF9jumIXvlv4X8+mRA9I6v
SHZ3SZ5gsk8yzuV4Nj3Hbffvi2SDS/8B9iPW2SGfUp8ydJw8VsEO8pQUiO5e
LrKJYT73LUUlRLCSB16lcG0DBu3qVNiIFSPx5FP/XVD+oLcvSAlng67VAsml
5ZeetRG0lPvaro9FwNRC6LwyPO/pryIBcNYrVpxr1bq9tiHo4Pj/7Oxo9jTf
ZN8oaOMJk1VU5KH4Nop3rlOYROeyPDfoNrMaEyFq+e8XZHuVn4Ehf/riWFlQ
J6IbfIp/YjPh+WbPbq4rG0OrhXQJKqfMoTKj2LLo9ewYclTup+Bg39RG/er0
8Amx27EywZGdNp5YoKwGl15G46nM+510girGXwIiwLAevkyBz9zuMFeJBzAx
nYdTCb6GbCOlAn3aSjudU+YcxbG9Ry+EbnIvSN89yNjtWsXA+no3iSuvoTLi
GWk62vQRISTbxmzKfX99kLA5Hi/U97KyvuPj7lN+rYQNwpF7APttsuie6F6G
d8A0nszE2T0u6in7H0V2zLiiD/PiMzamgdNPoSV8yNxlsNPtXNP4YG9FSK7Q
2jwHTYINkGrlXuIaXnJ+QaI3xT4qd+8qMRxOIshIbwfG2SFcJwtaeYLSYh5D
AkLIR30gH94SU5gQ1UX92kad+ZWGUQ46ac3bsLWg9DXkOAcGs+feOVzEu451
yUzyanU7ENCPJ8E75//bQ93chqOUowTdC2FiymNHmUVVBvjdW3eOLsHTopTu
F5FbaNupZ561zwwv1vEG5absyiv3Pm5srGen/1VHFOMcdF5C5wDDNKPoTtC2
Sh1DZEwBZ9ownSv47ip35KdAOqqA02+NMMM5du17SVIAJYJmZcZhs6Z7Pzw8
oyob0xlW6ZKe4U9XFHvGkYJY+3mWEwSsWDmo3bkI59ygrdaA0BX5uKBom6VW
8EBGt1i/f1h0pgtTEynPvx/7Zr2d9GJS1fKUpaMs5RB0sEetG/P5MTPkeK1P
sAHKmKBIWdNllUTBuMlSi3Is5t7mVbg6I2qsDGSm/gJ85fLw/TXjqwuEP5wf
jHESbRRdJNA8bKPMsIs9KVjTd8fPRhrURDBW4gRYEDM0NnceykNSoO+cImtS
5BxIkamP3EPbrxiwNdW4UaUq8kgVKcI3z9rBvX6ojxiyeDkHSi/DY3Y0PhZo
afCqShTzpU82PIPpvlGYcJanjzenlwmqrgAsAYTAtw8KUTnZIUKVYIyk+z48
40uPXWZPfdrMhzuMfR02kDUDzdIJVIULGwJZdqeCfx6a0kenMeKqpE/314Eu
CCYiRj48so0ufRKp0XzhgRcCzbw69fjxq2hON2pVzAto1nXghSMHDduSUIa0
bEVv4SdG0EZsmf/fgeP++l49iiw39mNwLxsfSkgCscSr6Wr6/w5tjDId+Yij
XYrI0079WR/ZLVvwHku3YiBhlQt7qKDubJiRhVNX7MFvgkmJCVQcRqDKrbQ0
P6eEXYnv/dcwfhueilRnnv93zka2kTbqfxccbUk7mz7lP8qbUuCSenITbF7O
W85c2HRzVn65kDLvaSW6E0vBSbwW4Z0MTbAVA4xJAlR7Z9SLH6/M7oRbAhJ/
53KGCdBE3AwvTDLOz8/oO6gsBLTLXwoG4pu2KbCjP36PtpFxTgkuxYHevLTy
TNWK3G9kKwwk5e9RLfb8f9aCRbe0c6JvO5c5ANAk63dwxH5x7CD+aSP1TbqG
mbw3YtEK2LcTOyHNaWGf9K2SVqTKMsXaJUpRc9vh947meu5rUw7w7oC+jTJY
JgMHNyw1iCTUEg4ve6VXPqIZSjM+0D8TAabXIlQ3iynLfLETTxvbRbcRj3U8
vDRpjs84RAxt8zvxqmoBAosFJjAaeCaeGF980/yPVhoDUB79TfV85IK4/DuQ
/c+T4iajwp+p7zZT8NxTdM/WbG84vhIl3cQv0DovUSTDHMMF+T4RopyquM5j
gCXaUtC6xHitbFQd9gC9TWENgVmFf1da8YFRHqDvDPDLN2ZEwSdE2Q18hqQs
y/o37zFHrm6YjODdIbCSlm+cKsrVyrlunSUvKCkpvWGw4EYngI6bgZYqyU+c
YprqrUfcE7zy5rlF1AJGcpKbjgBof5OeHGahB6BNiRr/3c0uu9I8S0/iXXQT
w0Kn/4dk016kp7JTyORTd0quQ/wtQlSNC+ld/ueslHvl4/br2JpscGqJaD2w
gmQR4IxTeS/1lx+zZ1N6U1XzyTU4C24jZoW0T3l88sTzdd1mKa5eqBUOX826
lDUqS3v5VceENGw+ojNE1/sUfSt8pPl2thAL/SZ1PTCXy1Pv77cTOSEOOJHX
hxRQFMTaRB19cHsjD/buR57NYIDYnkE6e+DXCehfXgjOkTUgCxjAqf+a7J99
pKJGOdzP4N7D/rWJ2m9moZsmKMRtAb0YdNEi51nZ8in4wgIo7JWzpT10Hf7k
P433lCMuqW/pzrU1UJG1moFxmOl6UbU4oeOI6zHX194y1FgNxgRQ+9ewYkio
YGUfgWTawbEcATINskoAmivY7+WxUSEnToJR0R0KyNZ4xLxT7Oegzca0tNcK
Y6i0mbNsFM3GJbwCj998JP0QRYB+Hi2+bgH3zjPmQPv+XEjc/UF5W9rc7Z1r
P9g2dqVKts53iVa6EtYYsWelEKIlL3CDq2iyP4/AXdbv572wfDGB2TErI6wk
d9KMLupHWDcfIxH9JC6DGYoRZKL6Sr5iU65Sb9O2A28LMfyhl7nUiy+HnFul
zuqspABOA8DR6qo0C1xGEYh8HlXnVuhaKwvF2goX3IL4zXU7bN5++b8bcMrp
HaZOxzSMmWyrqfKBiPerX7kYEaYmwJyBfLx08O4l99s+yyLqfe+WW8v6argZ
CBGTvzBWyBRNP5u8d3JD2A4R4LwXxwePz4MoRshAt+JD2qa2TiWI5EM90K2M
kul3AC0gn1A9WNn7O3SFLpmGOrUdm+M2yabv6qjH6bmek199+BFjDqhV5j4n
mNQtHP+gj7fxLdnFMmwYEIu+hlN4zBSJO+kFl+ON2ug/3FS+3ADaWXKj9NoQ
XDoG3ymPsg26PGa1fCbMroG0p4FkPS8EKawlc6ajKk+T7M1EuCp54Dg2W1V/
q1+7REwuHnR8/7KTfu2s29g4cGT7001Z4UW7dvX9HK6HhX1c1g3++jsmXKYZ
a28d0bjirnbEROX710q30iYu59Kaj6U3M/nwN5s9UZbbqi4IskKaaI7vNLyp
37JLWqD4jn8s2HHTp+4i9GwaePhgLON4shgAQPHx4cyFqrMA4/I0kHguS3lJ
Lf/ITSJFBlFMT84rxhGDF00RH8PYWjA6hqz0Tc7r31C1brYD/EyuOBUo3WJp
fZB7EBLszQ4ZphgHNa6bn6NTPCZdwM2S0fb6rzEqoGU89H42bGN0GG73bbZD
C9TSpkSpvHfaXwTOdM2K5y2TaZQLwcjpFE6fCaT3LbQ4/mS1rzM/FY5dtTnM
VFb9FN4xauCUBVxVN4i89wWXp3sxqY1ytqe2pMSD5NH1fH55qZ95qZUADSYW
IhhDWlN4dZ9fqum1RsnIRP8SU3HgDFw16i7Ak8E7pGOje5+XJou0KT6DJAjy
LJ8+k+u9uERgfr2JazSAXZgk0Ja5sYqbkxmcUSmlDxPbOnwmkYlj4j5lpJ+R
Jbhf4OgCSwSYNd2r1Fcbbw/RbfiI2Takx3d7hSWtqWbm3MOgYszgyT3CHdva
zzjbAXyOau5wy29Fh53mi9e4tpmbb82Y/jeaQGStwJjtmARrQW24/DMpE4wS
C6rh1ArbAuRSSC3twf/hLkZcNj3a32II5+H8kN3khY8nIxf8l8i8lnoipucz
tAjDqnXFyZWKcJ6KXHX+wkjJ2I1mrmzIiQS4oRoTLkCdz4eyrrrsTVpzaOkG
r3aLcUkfl/UBWxCG/71Z6/ThtqO677jjJsWv/k/SnJvrlHe1HQiwRtRFienr
Go8WRDUzppRBLujyIOXNT3ICULMxKs7zNP9GJAcqltpqQmPpzVjzTTH6PHm5
araxxC7XgvOS7JDNbQXkBnBDVqSOSnTiKGltswtAeRGTk9SMzAgVWIAM03sx
TwAtOH46fq8blSOrXgZu5zXFWc9MG9slQx+HJWP4kk+bLxRysx8/MZTuzb11
66kHRE2QN0+PR7CAwwGGJA7Ehn3lxz0c88DUoSGcWdvc54Za5s2DhOc2v93C
AG6OwT82lqk8x9VQrC7V6BYIqH2LPoqa32VYlkTOheIUEE2yamkp3tIH3zqO
x+NFZO35OOtYwlqhyt6P7xt0ekJkCKl2EfoxhPgS9ckg3H9AZKFfbicIEjoQ
YeaC+82k6okzCL1nLRYJib3aamHPibPch0M87p3MuJtnN45OFvkWsSg8CE3y
JJmcyqUyU1HEGUsD6Rp1kJz0ji3iwfL7JjKDXgMEzT/+ZtZ3PZXMQSBYdn80
54LtEyR3Ef4ogLkTMhYZYbWMEzdBFOCiO7/HODD3eLdm94pJHTVEjAlNgG+i
ZjkI9MF9VOOuMSP+mozHhY9UBEEVK/JcjgkKUmxLmSs3XlWo8hojdGf91wbv
ahFtHrHqr3ZT80If++ZQmIlhV36RnFoy4WmZF3E/IxwVI8N/L4IlnLPwyKQd
5D0+OTG7d4YRTfa4v3YxC53OqqCX1mQ9fdLy8aVHgMyBbzajU6e404MTCrg6
gV58PABfcgPeN9/6nKcMqp1xfTZNlvXcOVZzWwcUsVy94Tvrcd386ItlrfcB
2u1YmP36kkU2AsuNv0bVsaUYvI8x+tV6r+rSMzsEMePXwI4anhlWRVZTGyoa
drwVu556+Ao4+7LmVkKgPEwllv71kK0H1I5BqwQOTtTI7+YXWuCyA06eFT/v
zGukkCwsL5S/R30hn4t8Z1ni3glufLPhcHAj8J1LFgKUBqkN8eR9m6O4upPq
/XFlNhGu3EObMscGpscj4LscJaR2zbWt7l5Gd8QOoD7LGKOFxjMCKdd44TJa
Z8vVbV+mFkpfH40GDY4O8EYtSWpgdJudfEBxIZegpPXqA9/2JZH8ixewjFRs
7ceXnmljvMHvIfoIla5iIfVwDVPE6/OMv/veTht4r6bSrFjiXtQzP//HtcF7
qJ8Xx3RpOn9SnuAOmLXhVuLj9uV2j5VMMqsmaITlOTOVU2rEoMQjRKcsaf2j
SjStE3WcmNe8iKYPlqQ4IpY7od7SDXASJ9GOvUnKr2lcNEiiiU9+EeY4PWgb
BdBNPAojSeKqBeaOZl/zA3nYQYCSLrr1vOFxMr99mrfPtf6DNh9AHHQiLFRZ
XHhQ1tMswH4dWiSC2cK6qYo/u/6N0SqI7k+iRXWghQcEAFQaYJ48Pt8QZOrZ
dtSd1cUBm+muW37hDwKVnxsGtWeYStoXFLAeNCe8ODszDEzvE+Dl6JBVewah
8D8yJpuLf4pMJanGNyGkDMhbw1wf/kdTrF6suq4sDW4efzIuzQ1bmOTcea2j
AJYiqop1CnCytFhLZF3JD6+SQN+o4mxN3AAcN/biO9xHCfZD5Hj3dWLYWdqf
TOwUYLTKP7l8t0iIu34qFS47ltOdLG20+PrXUs5bPRsFFc6d/kHG4SU3PJtZ
pfqw0TEU+uZ9hg6rWWxMDFv/v9alH3/7iRUMq1YuKcsWdfKS9+6mbSPvbh5i
3KQk73mDxfP9E/hNy1XewCfue9pvl9s1WM49/e87no7FXfj36CTQsluKqznW
CJSSr1AAvJin6ElfRFPJt4LRCzt/eV3xQHOqdEKStaSCeTjwsiiTxxrCOkcM
ZqMPe8I6y+aGVYwfcxZ3qJ0an/7sYTYBLVpp+DRWnf9MIjGTXLrgDDgOPGZK
77BoszVcR8qmLjgRXx1VdRd+vriW1pXfKDgGG0+7+ASsPQAeYteLp4xj6W/5
0db6OeuTR5Q3B4M5EuEJWDFNdBBUhEj6tLGTUH7zYQUBFlyq54ikSaMzxNgC
P4W8uDgBQwaGG4GKvU74R3CAnsTqsdKy5e24RWRM+DMUE/EX9onAzIOIlZ2j
xfwh3gbR+69HxvQ8UGNCoZ/P9e5mxzjYfMMiIpVGrCdjvWMiV82T6I9hhgou
YO8ln/GvxmKzefrDqdjq6xxw0R8LtpN9Jb2g10Us3JKsXfBoC4SdQ9xCVEcc
o1LlgYXLrNcp5NHNpmrbwFFGpbYIet3VHmanoknPHJ2eRyyzEFgb1wVkj8QM
DovTa7urW5ewQs5PvxJmnoo66EuQSZdB4ZyDwmasKDjGM4Cms0lARltPpoxC
2M3RG+szqyN9A5JJbK4bIZy0Tl61e5NKwjPeC6+antgQk4UIB8UPrTMCJBTG
dHblrocKU3N23nHNeXLgQi0podtlpaKNyLuq77PWE5YxMpwmr8j4gHL+Club
2WZBGbTiVc3KDkvQJaSBIhKkIjHLQB1sFaQBNStAmGV/UdXtjfSo3fYIKqGN
tCJczdeF+igQ5SiplltIh00cUmgavDURzT7YGEExtol9qbt3JPBV+sE5qQz0
iGL8RhUWR/s1qhNCV2XEEvnJvkRyNcuu4HFIXtI8nNH3Ujm2gwTMnbFj1aZQ
tkBbW18kDV7Mnp2endVQQ67WqkNvJnEvbQLArmW8LvhgRDeyqdQC6rwNqJeA
1scqMXX8tmKL0baiXAUungSsd0wZHrwoIt3GqU7hw8HFlsLHnMHQii0t63WG
N2QD+1CRyK8bAKqCOm+dvGJc4lvOL1wwC1A0GH/aJej/fh5aayG9KyCGR0rG
NCr3fTn3+Wi8TWAHkyM94IO1fuA20zQ86CeNhdxETsjluY5Gn6U5vppSF4Be
5LIUm8br04qAdTc/NyZ1fwhDZvNPHOpL7iGBrBQsAzx7cqjggebyGqje3x6g
GPm85LFFrhLe5ZWMQnaSNoDb/tnpnidffPU1S2GuPIS6zbsL1W3RU1e7Oc8b
D6jOtSuiB0WJkgs8MUavjs5VZCrl+kyOWtCGe62SSccvfuPbW4HvN9MNzeQU
irP4Copy8RRnm4O8nxf8qNjeBhhfpWLO08ZI5I5N8G7oZoPQMmeSkzlY2egi
kDURLTdt61Q1emJGEN4Um8uCyvGWX/Pmd6koBicKIYDSzIbzYRFOoFDIRcIn
VrCtc3lHxXsNlWiUabfKjnevGN9KHOxEA7S3C2PJh+echN/jQJheW2YLW7sD
b7Gssn4XUrZJR/BjcieZ6HABFserpvFUWHXAOL0ILePvi9seN2qBaSMlUW28
BxVHz65+8HYugt4S3cGh1ztSDIGXnRaBSZ8UEMNMc3OhKkj4Cp5GsS0l/QqO
MQ5pYPgLx1MJMf7w8RU7Ojl+xi9R2NBN64GWesXnlOO/guUpc0nB9fWQIdYR
pV+/bIm7sA6S/7uxTmSG3CMuF7pSCoOB1WUUZfCrxYZeGLg0IUtJ0cfp/S7Z
nKByzYOuQYZpkNQbD8DmhtFslb8m6xAhofjD3urNzIGjMqo0IKare2uze+t1
O/qAG14qjAYPDg8KiV6nD3iNwt7npO0k1Y//9donq+85c377Vbs9kyl2tAEn
P9kotc0UppxWF2ITUnfOhi25mZy83bSOCa3ksQq03syWYS7U8ZZMSjSdOdA9
nmDSzqNz9Sb4fqcY5M27Gu+ciEKskYz3wGcg7eMaM9CIeOuk7uIJYd4SN56d
eWWZgmeicIo/SCKJ7P0CXMYBNsPzC6YJIwnpKKw441bwBJwruASH7cR63oHf
8DBKD8T4/vEidZNrb9mKkfezNejQ38OgYD20El1tgCHQZY9w/h5+0fvhzQVU
A/ATkaDbQFt4XJyWPJdVY9Gazd/cE8KPIq34s1dKqBYQCfLvlO2e3QbO6uUy
/NOVYqDd19Qo0KwpcGeRW/1wF3DRgNAbL3VN95gqJdj5ucNVTV/XHPE9IgTu
G6BTtOoJI8PPezSQR76/2N9LiJi53SAsmHojGfc6Ps2JtaVlaW2gz6UZSV1X
UIIcTG06DWK74yg9fXkk9VYY2cT0KcEA8SLC0BBeb+ihmDJ5uJj/qN83W04v
6tgIJeLimGHVuuOBJ0Ds6iq6xHTKZFk+fqkIqGEIv+UV06mdZuSW6OcwGM87
sVKGWNg2tW3fuwzZn+JDqbEbQ4lBOuAQ7wtdYNEdLaOzhWL5yrEEtUK2TONb
3tZWJCLaeUFaCrjUFtOyBoNX9Fl+FCiPsfoDddlKOLI77fUl2ErqoSyTxEsV
fvjJ11Arhl8v8paXTb2uECqnA4+T90tQnH6Gtr4+odYuupuZ0WweCDI4WCUG
R6P/CrrDoHc/UaeZchcS4mzowtLEYbTnDLv7dOiAp6vIEskWI+m9dshws9Ak
GqK8hwg/EhjM7NzYnQ7QIFh/P/UtRPYNvOXQ163LFNQXVvn/2nlYl631lZ8U
qImjwJG1PFsiSmRhixfGm24xMgMqxqRYL901oxpADw1OZ+qiSrlfzpL5nR6Q
UJktu+ea75BOCTSHyihbK+dmSUVjxjENDXcUdw6eTMYEb6OHd7NMIrvI6p20
IGqqCR6/7sQDmeoHNM7h+gmWXtD2oRvf++JZsAUmOqm6XhMa9qQRBDfWCwvd
IGn+zKiRjzmdMrYPLREhApmEt0UtxFkZKDUZQYNIUqz+g4H/wYMfjUtVPmlD
4RTKA7pZOqwDPuq2xpktIj+35sa9OPVPY9LqpdqUnh4NLY1zV/omASRdUpVc
TXnGXn7TFpbCoC2tTKFTdotogAvAiOnydOjV6B/5p8NqaccwN6oQiNMvAWNI
3fjCtlepiJ0g4tu+A4TEOfEAIoftgvffvCyfbQA6D852TJquzwgay7xd8/r/
K+2l/h6tQJGDpNAqLNYabftU6UWnuA1yRyViF+2lkLFhX0xe0nku8iOQWhmn
AYdiX+UOZons46u5hRAO4jOaF7QsBYIm0zYj6gFk9CkkTRsZIaIwrP2DJWxT
FnT5eE+p5yHdJFYi1VnxKx41gVHZTbMnTQViyn8cFeCTFOsLRipakVoWyzus
L+cMC00W8j6Xny3fXfFFoCionp4gEMZHdGXnEPPAUMAI+dGmzUjjPeVMQXLK
J6FBTA10Pc0UtDMfIZeEW+DM3/SCLtkt/ikOHijJyPBLH1TSEc89utGOaWTT
PmbvsyLi9LnnZQWLh/09se2aUxa83Fy3wbH5pIsQCfKrOO33nccs/G1qw64d
1aXkr3MikVrbMr3RcVOyVlCdU9/73XsffeFQWZrSW6UXCKbF7iAw+Pd0tc74
z6SpVb806RzCvi3uMZEgUrkZZJ0kPThFxjRrOQtgMByrZI/A3saL1nP46yS6
SQHFjMlLz0hjQ4k2aUxD4MYQyDjR/q39Zq7QTiMbgyVMRY8hwkLanXJuvf66
Zq1+6htRTUZfsTFgLrWv9pLYal2UPDKywPPvHIqJuULC4W/q5ONenzhc83OB
G8dXejx5NoGC1G9ZGGHDuhw48NYeDTiRALlZKkk9gAjZnTv5OSeM+Li9sAom
aOVAlMmwgTyU97+2Brn75+hFDWSY2HeC0Tir+V3jN8BXyrAMNPPwHmtOPwtu
mWQcGLdUbd3mtC+A3v9wCSOjuCW46JnJPpsY9IfGQSGSQkDids85U+LQS3Ui
RLxno8HVBrYkd9fZVxbjulpApTEOc5KwpkQ6KNVkqWqbDB0I0zJvEoRdUzUc
i4OJC6TeiZkPvbIXZ+1wsDLFvdv1G2425DJ+/L/UtxozeVW3kvNJ5eMdBi8s
r6snCpkez2RcMajJ/3mPKjf/TmrPwM5jbuqUyb/KJmoDZetqU4j9H0o0mlRd
V+m81QbejHPOw4oYSol2siDpCv1zapP8/EhP3sdgAqHubej7kbCtpM5wxn7d
O+Ygg9UTF56VehPyNbpGk8QgK/HRGDrp2DV6prpBwXfbofw40UckJz93jRw/
Vjfg7fu2lj/w6PZLicCnuOhYuZnzhTbRufcDNVOV2ypjm7klChMRbXoSCcJ5
/vhmfrswe3wGf7/hYFXT1TzqLpe36Y6brdkWuCPHH84IEIxB1rkqpTxYvgsR
8xKHssf3LEFmQ4i2Hxa5U4vkGytKUXT8cfXofE7O4+MWNiGyX2JS+TwK5FNa
+FCm1LVRLRIXuA6DkZ9nZ9ibi1+6piz6D2iS7VAk7Vu6Y7BdUJDtdV6Ioez3
5i7IG33tPNirNef1vUWodKYhtsC7oIShJq4UhfHkjGE/VCBlPUkgHkJ9u4Q4
jrRq7AjVEH0P81ggsJpYs6N4KXrTm3d6nWatZzOqbyh5pr7Xd0dfhu+vR8GS
sIrJ88g6OO0JXnBwVsgVAIdroP0l2KgdBDlN1Z09Izc/CWYXb0bfdTNzwKIp
RG6M+KkIKCSApmgbwBwiafM4Z1znCNzvbnabNG9v3IOVHbwUyYe2C1r8F3Xx
2/W5XKYUa17bnhjHzkxtt7h7wf9Am92idyNh2/Dp7tLS9yE25KsWCPMdS3Pb
MDz2iYsgyXCPXT0KgPMGMR3Tg7pp7DRaDddMVjE10H2qx79D7Vaw4Gb5RhP2
NfYwsJrx1+zamSurSpgeFs+Fw2i2Wchx5Yz8KC0bdNBN9IC/T1TgyN89NHuI
DO++JOGnbtTaQWZdGUvo6LNGEM1/4fSIUAQf1WCh9EKTt8GrhO3lGrrr4/EX
qJ+KV3HWHNZcZEnVozBiQumcC3abk1HoBv3bBw02M+IBAH9oDBVWRF+28Bk4
0FJYxl1sayHGkjGQyBEnRNF8RwAUl4iMmi4HKx+E5P2EyAZKFMCgZA7cPAfQ
bv9wCrGR5EK4dGQg5ArlLu/GuyemQSMNGyDyU8MuTL+duWTlVDPo4Q5JscSy
xCJe9YRXzSOqYwrTkEA198m/c7foQiSNe5UYHkTC9us31rzEFQpx/dxFKpeG
bUIxONgX9/DUpRRjPgaDZAwnGj6g8RnbVLAaO2e2P8+a3KTnejFU5ewIOXZW
QKBdIcQ8bjEWGI2ZyihbPm5EoAmw24NkBFdt4vYlVgci66qCCQVZkrrnnyRU
xmDZnZ6ItwcGsqC/fwQqrqTU92Q621Kt8NGMVCe0pZBEFP2Bv7IrKZ2hDQy/
jSqxxkqokmRRO+pEUyV1ZcZ7nf/y5yIFXs6cr3q71fVKI2Qr2wDV//p9rPY6
zD1b+McioqWJ+73W0TC9iRKxXVlCJQX58IKGJc/Aq2pgiogO4/JVWTZreaFs
Wb0n8+HC/qxkEl5PToSXJXVMg5yHcz0MGA13zqo/HqMm/CfCAlSCvRo81p/X
gOYPdeHm5wrrObZCx2af4Q8EEkj9kBMlpORe9aleFc6AhPbkmuUKVIoGSccp
KSBdIsZXGaaOTVvOIb8G1jEV9PzI1/3ugWZCSmfe3dTiQomZPhmD4CD3On3d
WPHzbf+RLyYs6C3xsUHCyVFxqhnj7HNmKadMRzDmIZtdq72+tip+zHwyE8M6
UF62OFO4MQpmBDxHOpVVw3gJX/XFm/wwW+SVEO7O7iQzkP5Ddbm3LNIsNahd
Oy7An8YOYtAMdv2SIYpORIdajyPdiXWWBDoLcwvsDUaOmdiLVPjkT9TMLoIT
cHZCfpbPLTERszLebU4z6//M9WC679OFeI8gdV+jlwom/g5nY6yG4HNChTUm
fe6V4NTsIGZTKNbgurpxLNdxA4PDO63Z6s2Tjl1M1e9nKL/krQe0s9X5eNn5
w2QeTj/Uw9Ai4OjcWSffb8Z9sbOa97Sa1fasVYdgMg77rdDmZ1wA2RI9cPNI
shUSCK5gJi9Uff+qH0hORQifi9CWAzTgfpPRKUrbJz26nQU+nIlizSkTKjh8
vpwoVYsYyQzoqPy3U1oSM7NIK6e+WfP36jQc1eVtdZW7B9b9kJ/YJv7+olAq
0mQkMVHIlEJwvjxghlVjlTljqms7FEfsEDtUX/JZndr8KtUQDQNC7fbBZyp1
ln0h+s1q9UGnirOGH6/s0xRjj3TLo/StYPd5LMiYHG8psJ8fUskBnxmeDjz7
4e/y+q2/+zsMuzjsUxN3l6J3F/6BZcYDPPrvavlxprPhv7yW5II4esGkOdEr
wZ32uyczRSe0Mqt8F6Jf1egohZzTt68ktkQaYZN1NnHntQItEQgzpFb03oG8
Yat0mfyixnfN9H24a63Wtan7zqy9b5vsONphVzAouhahDmfKyig839lNP9q0
vrCxgW/x35r2UT6I5ZwG0cG4EwOFW2IpZb9le3z2rdbBSTG1dmBcmejHcyI6
Lp2Bi0w0U45fVEFBqVlZ/StG3a+gRqyjV1EQr1yKC3gfW2thpxO70T56OMhV
WDsNSuvnrdXiPCCAzRl1yWaIzv42gZ1UnUkCK4uGLzyAlA67crYqKZu9611t
BVjYa+HGPkZQY+U2xtwqQ7CSHchjidkC50L6lmABacngPRcPlvOAKqrbr2lC
S29NpPbu4keJPyg/VfHwjSfVoxCqnnvIcT2TCy3UYQhJbuEV/l6QxS5HUX0L
Pi56n+21Fe5745aT2Aj84caaCVOFimPSsMClL8oML8PnymCpe6Z/MhF5NhmM
EiTpG0AuA0PCzGtL37qI+whxugeBEEiJbYJcgzI+OyOx4/Z1/WUy8u2GgMvP
v+/8N0wxGrBPxvYzVzOabgKjXxLH8k33oLCcM+qrHG5tgdB2QdOtVDISGNc5
Ht2TqwUj23a0nyZE+a1hajKcqVSJ/KaeddnwvSvGW+R/d1tUtgNXCcO7S7+B
Chkwf5wBQ8MCgnt8pX501zdw2vrvjPSErq9p3/T0OyHVVprXY6EcHj4AuA5n
fB2rJ2zNrn0/kYhK5U8BBoa0dl7NauiYsfJB0lgspXzWikvwsDb3ew0yR+c4
kHtFca8RrDfcuLPSbuFKLgfgNZBfLxl3zRvE1TZRd6zRtNoFVKP02UxKUF6d
I7nKWbqV1x0JAxWOyIlggWAxULt4bqj6UGqagYuEo7qRgr31B7HjVvjU1CSE
93hQRgGWIfkKgRMGTo7mNCkwYwG2sXMVF49ELBHcy0oGWORoLwRrG0xdASt/
zMDnscNKlqH5aJEbC/haUEWvbfuMv2nLj8XSsOSNdrvRC7CrtNJLsEAMTp/p
eDji6LZzLlRtZhnyfe+ijgm1gC5CMPb3LNC2ji0M62hnIFaYNk6pNEWk2tSJ
zFxhG4h8Mkmz4hMVZtOS1Ahe554xogYvJGMtqujvGv2ZMBwK6LhWlbqKemQM
j1NXVILHHXRNBknaYCc/V1gs9kX4rYDf48eYeCUxiYxLrpvszobrH7wYf0DM
nDvnuqoh1E97GZHuuHk2Zg2eZjLZ6bOwXVSD6Fgqtuy/fFiX5VADrFjQwNlA
FAfI/mL3urKb4c+sh78qOEXR3vktEzvEdSuEDTtcNeuZ8EZD6fER0t87T2eu
TFZJvm2pHpkDShcDWyYZKSQp7BtaN5Yqg4A061k2DVvgqcOsH1YOyCPW16yd
ey3hslQiR/N8oJbJYV+rY3XwIFWdI8w3auAEkjH9K3dg9Fo6gDd7eT0Ta2MW
wP43OmTSGEc2lzV1hLttVuW34eozlEi++3uRo9MBzF1EOll58U5oFpRSZFnU
R/Bt7VMPn6MXEL06WWpsvaPoj5rB9nq86BglajF1JrjLJnzGJW63N6TyNfE7
V3Dp0i+IGzdJGmI7tvKpIKY+5yI94PyM/X/flB8KOyFPsl6fmxJVyymJ00/y
UBghmpzk+PeTQmSF6tKFk86sjMYj+pRwH/CviYpWu5jX86kZy17q5hE9/uWK
UfDBnNoC3xAbAPntTUB8WaGMAazVBN0pVLSK3M53B+Ws93qZwFmlVxHo53rh
cGnS1AHsTQG4b3i54utw+Mhoa+G2IlofGwIX+PN1cbJOlQYVZy8DCB0Yc4Il
BKIOAjoxvIcpyLBbn3ppI3VR2LP062ULvTBgR7elWHlwa9GglkwiTg1KxOQt
o2+GeOsyJ1zQ6pp3lG0Nyym7V6cT2EwjUXadk6mXnBVukmnAUTd+br5kQ5DG
n16O7Qu+2ZQWYOoA1nxYyjFkN0P4vUg3NUdakUYaN97yAGkzc9TLB3Ts5L78
4EfOlT8pY+MXvBDcpEwWDn/9mMBKAKAjnToGgqCn2yvskeDyI3GuFgn+A+r+
NCn2q9b2WKjrot5FnIgThX0ewxB4/odWempf2ZY2eYYzgPk+v7vx7FjrLj76
8OOcOSU4QZFLb8wLupucBH1lWKV8k1qwC9qAWjJusbzvaWKpMdXMt+p9G+sk
U1Q2KjSckFqeyzlrZ+vv7+aw7AQrBgFBJd/q+c3Uxzc8V7CEMK1DeEujItmj
ruSxTVuGRSiqRVAFiUnueZP17j34niz4B7ngiQJXc8W3C5QeEt8IJ+dxuAwr
Y8BPpQwT+nzWRVDRRCbaKynXvfiWyCTzE51RNop87AzwRs5XDPM953mGT3YD
XBynzgH9+e7NTY8VtqG+og7VTBnykEDdOPzblQixESbjYDKNrVGrupR0LkUL
CVCX8JovZ2HtWrzQKAtt9Oa+Wonc+H10QPBudptqp+jpk2yKsaQi7rUjDQC0
8JXTXn5y68dqtZAMTTfTJOjKgM0Vlk+T0ldzColR332ylCXST9NCla85iKd6
sp/45qeKY1zUZsEqRNRlY8J9QS7jcZYWCSAlbCJWv2WY+FWGECZunc8Bf1zo
3ZXGkSVqnvSOe+ivznx97XY8YFD/YSZxYE4ItnT0npmD3NnJTq+aSIervanX
Wty0ln1DoGrKWSkCxkrZx5d5JUdL83wyqLwAZtP1aICtOXt9fzuz4w9Psxcb
CK6/DFSjki7AwM3IjOcQ0PfnvyY1gKnpggdbzh9VUks8bavJYHo32RZD1l1G
aOMZ2wF35dSd59AmiaFbGEptSBafQ9zoQdVqCcBq8ZhV4DjW5f6/gHSvNT/F
wH3NcD3zsxw+Ur4/RVscKGdtKxlmuh4a65Pd0SPCydGqjtwk2OjsaXFT1XMt
/p5J66ztYBDttAmd0wJIN+awd7kOLtM92cFrZntvol1Z9F8oRRItvNZkmA5E
60hLoxys+up8Gj94QZW9Zd1dXHgwCwkd45SUwJZseh1RlNwUL0mFlVDaUGlo
PruAMxgrP2KICKBzIjlxc+vWtZLcr3T/Y+EfwozRZMfoos0DGN1U/0x36rZl
w1edbbY+Q3Fey6b8ogWBaLVDrs58awPQqCc8KWy0DsNGK4Hcg4Q9IZAc+gRL
lXdcdVgksDB9fFmYOufH2xaDWkarhelDxZhFhPno4hbLKs0rD6NmlSi+AH99
tV3+ICZ8Tm4YqfzmrxZNFE2moacc7PdlDF7RLqawutOGSu4yEIh8H8avp9mI
I52GT+d+GhuWMwpRgUQB4IrU5BJ0COEiEb/O3VqZEhSkbUTzPPc5/Ywj962K
H+aCuu/hh6tuW4RNC5h/puxLNPMHZLHORCeZ8whSKKblfFi590KWtUKB+VtM
e7AJrqu7SaEl0fqdwimLuC8qmNXIeFU4ogwIoJ51FKym1ToUnXUGQw6WA6Ib
iYByEe8xgmgOb4Qxjt//3NcsLjFkNIOAtVQuLGyfU1hQI4KAF4xoAyuKpO3d
jSjJ+od/LxPMjj8m//PjDpYEbfVVx/MvwX/oJBfxx5eIQKLy+Mm7I4tIB24S
L3yEpXEJYhQKjKLI3pG1V42Cl8yhEPq/LLozxqR2hGGNrWXDEuFRBP6Xojrs
6f0GB+YnMLSzaqU9wLv+rSzMRLIKo1+DU+af+CnjMztvQlYTLgFb6sQiYEks
DkMX2EzOoh7PwNBxmCaZvPua1GENy0kW4CJRkaSPVSNXqQZNSYHVcaX8sRZw
0/qe2h8wNPcJP+wvLCYZ+HX3Bs74hpvdxhIzSkuXU7+nyDzqJTrDU68d5xzP
aN50HhEVOohCC4puydqaACVZhLjPvUCc0UexpXe9U3bb9zdMNQy4Y3AtjBrf
6zMi+YRsxbaQnxbaxJw23rR1IrYjI/crDKSR/zgcyXO6XTfXqRvujkWP4XkJ
yD49HvR9UvdI6aF9LoT7R1pUTFHLNZIR/xpVnQYz6r9ysHuVOpVBJIqozJqj
8Zck9pD6T9vQWUHKiYFxUveu1QQQGXem46cvd6sQiBSpTJyr2jIUXiLLP2Vy
/7rI5XSTOTVZ4cm7W7kO9EN93XsJShO85EGK1vlKhMq9j5bqZfJIzpAtu28p
yQ902kjJL6d6Ol4b8HzudrO1/3UW6extPidfkZKU5rmPghB+xp3w8wm1IEiF
RVRherQZRkQhssCljlj4w8sj8CKF0ayCOd2N2m+khJXriZsvqHsrTPlhEW1g
FGBikBUUs0+kcMrIk06MFZSJHUbtOjCmBXsEaCK7Q3SPexaLoy4QlNZQ6H8k
Vrf8nutMrwvY/A/bn3UrazLiPu35JPy+vE3K8Qx7+Rcgw6vh0T+nBW0Fr8l6
O37YPjEZO5q1XaouvAIBoylWrxrcTljUPrbptackoMcqtBh9PNMXcA8N/LyW
QEvexR76pbBYsk+uAPzMLdbSIJ2TZddz+Gt3JiXqinPlpu5PU0DiRWS0Hvq6
gpjJhpnUswkRhLcDeUJ941hxTrIDR2BT+0DF54ySRBGUl3csoAE47YMD/O0p
KkWm/6Acxm6s15Sv/aE3q2gpFOFKVCf0bg34ZVSeBR/3xCPk5gs48WjROLSx
dawN+KZYPUm1VRWCHoiIIY9t6VEHipPCSD8UFzEvUPnnqx+z05/ObC2W/5Hn
9os5BuOHc3QAGEVjiHClAzTO9n99weoxpR8tBKn4FY0UoUfuIOtxaz8L9PYl
5Wdnfp1n6Ig0T3NDx/P8XOvZUszw90+Bz4Ne4DI5RKUOSPNPeK23fa0HsaHL
YNo0QCFZOWcYCdz6zNcYUe6PmRacbYYiFJIMn5MMWlnOrn/zZwRGUN524cyZ
JHHp6CtHXLEdtif+Yvam94EutsVxUF/nSzOftyd1gQOXCBXBsW+P9kbzBMe+
on8moeCqiO8JoEEY5UwR/nIjhiCIrMcvNOfDsmf90/2320eZtQ0s7I0nj49p
iqENPvghgBaMrQjums3l3kMzh3vrkEuOcxtketVKGuYGEi7OAIg7+Vd4nk7v
WT1Fx9vA3gR8VuxbEKD10954VH5STh29EiSlLuWuLj1LyGTzeSvUqQkLLNf4
JeWZGEBWCQBvyPXAcH77xkrWOzFI5sOMibvCoY3Amh+ssJpm7RfkG3S3L2/y
4zghPivCKzrx3DVUu4Ty8HQc2rEr54oxx0m+ddErErotswRobVFV0g/jXeyL
XyXVcVBtCQM0cvB62VCGoemMm7wQ9KAKGGzX+9UagP1Jv2q8yKTq5vWvxpte
PXUhRhyent+srfPxZR/WgiexLg0K8qXBKxsYb30XVu8wUMqsj35VkgbUn2E9
jxpl8vpNS0KfnglyMvJF5JdzJZtXibB8IFxlc847tm9wQu3raf54XOz0Q4nc
/Bjwx+guhI0ZXQy8fB3QnrNZMYobruWJGHrOZYEN3gmVtDXApul929MgHQYA
jpA/qjPaeigDkx4Z/PVMNzU9wIwHaxMaBiVTWSxqz3NbzaWtaXsQusyFCqql
xbMR40ZdmO243t5sEVFN5KFSa87U9nU2tDseYaT/RYo16XILLwuFUtQR88vG
PRAMn9+aoU2jPfFyfZYvG4KKdLq2rPVfxlbllgMTIsZQvbeBSyjwin4ij0mH
5LU+o9R4XFc8h6NJYqS/+e9XAQ6y/UonNdJvbN8jMSWUhUfZSkjvVQSJ1bap
c3XSAHA3mbcDVeCWVr4TjlfegopwSxcspIKIykIbrtvhAHn+ncdIUOnROOA8
KRmIlnJuIa/XPrP18Xec1F3WaTBdWMoqAJJbRC4wkRG2y4QzSVfY4pF+mBXZ
//+RnuawH5x54Fx9fn6geU1Qkab+miMasMC7r0U9WRHOqos+HpMkzjrRAsYy
HZSBPK6MWkYxMje85PVdtMUUaY78D9jKM1V5kf/Fu0gmCFsrMec1Ofj+NJGE
6BDLX2BjYpoh78FB1X5+dwVNkWrcF1ZhkM0qc3N96djcYRXJrY7rcy8uheN0
g6tqt0Q59x1aEncLG/vAfB6V+eg/x7t2fpPGYTGdTW7UMC06tBEnJQtfanX3
/zAhERNdhpXLawDYb21MFg0yzwEnzuTUFFMPqAbXP7iVxgLy8XXKLH1UZFKV
S/zwlfYHRkECvuZ1qV7EcUj2J47GP17BKMYtiV4j+AqA06vkbt5MsxKiLhEx
PblSxmmeqrTyKhrYdP2QkqNNDXJ52TSiY+TservEECBgnu+CEwC41XOLH2qp
pPvktU1bkHkxLZu98q1h72B4q1+HBy3X9SWS9/n0lsYM7p5XrCm7AZHZCN/m
eFRseRTR1M85eylTk/FCAIS5+ZZIpg1zKKbZXNm8r9lBs3JP47Nl6mSRGmoI
pLXqJkmZU7Iza/pkMufT9Z+qpYn7kUMfPiVnW7x+HHV7XHAq150LkS+iDlWh
3Jg3+/Fh1MBF1fgfQZfRvy1ikJExufAfkw49posSiSaL3FgmpGIopSKzRgxr
R1mUvbzQXg4sGtE7kLUtVCL2adsh1DR+CBA3mgdAEMT3N69ETDSIimLHfqjM
4ABFQinkOAx83NTeWwPbHaPPZDpdeSlFZHMjIjZJUZ22T7zrjFxTJT1ypYHa
WY1/9faptZqTmGwSNCsJrMF0MZDNCWsbLipZUAWyodX6vzP8gvflGed+RlPX
l3va5EnOBO++3iDiL1grZ4krPL7qCNFaYa59AudLSrEuwyg1t2EdHlaOS5NH
jxiUIqB+jtscWhpxAJLfDA309ZF0kjtdzWnG3EUNl1f5RfN2ECDAcDlLv3RS
xTs22Qg7joVGWRS0v4nFKg/FoZ6IYAGfHq6SIRID2nw0EvEnlk7E335y5tZ3
nD/dyOJ2ihpZ80gy0W4sfluBpwdWf9zHIjAEa+i41Hd0+/ox5MA6qReapPrU
5vQb+5K/LNkrgXauMDy3D0ISptqclfeiAOdXrUbB3CgostgVhihwyC7pGaqo
q3sLxu/MClrlsVLZIclwC7cAJZvU3HC1BTAbyxDEMBN19/vqceeg7n2Iq6qq
jLw+odLtxCkT7CQOKPrvGYd8tnLaqgXTGcNgGoGRqmgZW3Z+fTYCOA9DTRRs
HqsOqFx7La1z8CJtJZjstm+YiWSsUBdglCSiJT4kgfB43d/54bF+SfvlBJkd
9ZAGv7+8o5IWgsO6MbjYaCiCuN9aKvxSpc/8ClYusZwjUoWuopktuUZYzhV4
YQMhOWU/obML/EweSWpjSaFlyybtrX0b5Hc2yDaMI4iyiJJ98Q/mdmNW3DBG
IAFq8j9Ox5gZtwTQN0XM79rmiReXOeiDEwParOVKkffQRk3j1QpGWNI9pFMN
RpmFfJ1riJLKmYcwvjn5ptDQu/C8j29uV7nsS/cPvHFSNKSxlt+UJq9RLLWQ
A1X4YDuGhAdhvD3bF4fYqcCjeEjVBvRwOM0PIm9osaY01hW060P31qOwWG+2
Q8+iGEHhIcBFNOqF9dmRnMzRnqqK5rpjj/rY9Wv3LRI9Lekg5+JOks9bSTZD
qDT4gYi8KuaL7nViWvt4niQXuyjwaFqZBqBn6OkwJb7FUo2x6fxOJmnj6bGH
ewRGCbTCHFQOL90gECjNpgDwy6nopHWT84A+9+ys6kjEgthQ9BR0baBGAAhx
na85rrZ4MUfgTZ1Kr3DE9P5iMwb9N7zGWJ21ay91ph8LNfAWQgb9j2rSbwEA
w2KXf2XN2U/LOQVOnm1QZKQfs4ijh+Arw/7zyJ2xNrsJQc9Frx5kDTxJW8HS
+mP9y84eK+6+DCnDOEreEyA1+Zi8kZGetRobKJmg9zT4sEgh37dXaSRSX+VZ
vubA05R5ZqlL6ykyCYOkFQBSdQ73G0FAu6f5FlqwnqO8XV/Pc2XzXoRVmpLP
AxSWA7lo5Uze82ro3/lNGS0bDTGUhRCH1t4DmiMdAmjgiyF2y8Q2vQe/pMp/
cwHACmprbpIQ4xVffFXeBPDabDQ7jXctRHwbp625i04aZ/yioj6fiy+zE3UP
COw9Jl79RTRmJX5Y+Tm8kPlv7C6jOiP/2dTEaBzcRPP4OnA4PsXVJt3BpXVr
ILEaNC/qUjlE4CrhptLtDerqEDdW/WvoWz7nPVaNfDW310S9PBIqWceB+PbT
FejSte1ueKV2uLm6FA5O9u2RQEnY7bg+Ph+rhdI9uCPbFyXmkLs1l1p/B91A
XIrc1WjXEOOhLgGG/5cXvAquotfij9ntLhjNlbmhuZ623RE9qHOV3BBUJuca
t6AMGUkIsjAMVk8xIpjhwd9yRkkjmIvMaD246PwMBYVW/A9P4k2uiQsiJzZb
qMc2dAzTDiPQwnJJGeaPPmB7PLem97/jx2d8BkEwdJnh/yBlQpqv3Paln/pI
YHRjvKFe7jln7Sp6n4iuV4ibeE06N/54WBSttGQbMfAsVq5gVpch64w9AUMY
TN/tYnttZAf9C2txEWQj/QFRVG+wFlcz3agjB+yQNzLtlScvSaiFFyKmuQA2
7R1MJ/CzlvGEC3FxrorekZlI/Gy6C9e6rkGOAS06IARhsJL/kMGS4Yc+CAUx
z4tAwxtexzpyc5rCdUDAY5Rf/PflNorksRavSRyGwkjHsaB+Edw05YQlA0z3
NI2fX6ODs4FC8+sTmQNiYcKFwDphlodPBlJg+fGNmwtfZEokwU6y1eKO64fw
AhJl1OLBrOx2v/24YM3Gcg947vFRZRlJrDvEMnhYKFJs1+iac4Vw60E1SaW6
AB8d+SkVPi1fCrJq4wb5qs3a9JWharslXuP/+uGCrwKMNQ6WQJXbsAmZKw6S
t26gtRahcSHcNluGS/TIQmIf5g1vUnrVIRmwJu2Kq46ctygddb/gqvJI4gz6
OchvqFcNxPWvfBtyo5KbRybwLoNXyQDOc2B2vASyVbqNMnMR6LVPA4nDXcx8
y0XTVzyyS6t7JKYHsnK3ab6lmt5txNDthdcxisNf5HdwS1YX4Qv8w6gT4Pj2
9I1W6sdCNRrBFivDB/rTKRYOBsfDM1XUztbCrPNpDXZJU9kTt5WZtQ5x+umU
+JxWmRx6deO7XZ+pAIGrG3VoxqEdCBDhrx2gaW9z+0eeXW9J+RaPcYnzQA4z
IEofKV50anY2k7V/L2HRr64zvaLeDovt2MAwdaMH9rghqRVJWSqgvvF7D1DR
cLeK4oWZ/xBAnHHAP/nSpk01NRI2E1cyVqgHbJCUTksl2fUOnq+lguDmBdu/
g9SrDc5oJHnet+QUHbjJ+ZAHBbewae4Rn3LYHUTTNvQEKRNP1Cz0T4d3o0go
ciuJv2OPXDmdNJuAYNq2SKo0fVeYnmWaiAYdf1XgPna4nlZHcPzoBVjufF7N
MnZ1yG6z4Isyt29EiR55CQ8Hql1KL3ce4vVmsmRWlW8Znhhq0psfAvL+NbM0
ksymxF+IyQhjQ7o9q3fgtrriiyNT2Lx+1b60WZk9eqjnHCGKWaUCymCRRCJl
p0gSRosYNLrFoVU6y0HySa9G76Wrp4bsA9zZ+gBlHL2wUuVfr/8L6nBv6Hqq
tWSMgpHMIStk7h/Mox7fTtNucAG1yJS1VOu1lCaQ5SIdyJbbHDlTqoZ2NVM2
/hFxjRvYTJLeZ7t7Mqq14MLDKRnYGZGRhTja2+6JuWr7FXsMK6pS1+zA9ruc
svwdMcSGvBfLdWVJhyRRbW+dXOQNuzjGeTQnKp9GH6fTQj+f3CZ5qmo+0z2G
V5BFXSB3MVJIDj8ALjf4EDXNgMa9dfByai8mZLuGmV7+jqG4/isAI6CS6uWr
5B1KdzIIzi+qEVl0ZcTI19uxsNfNLk14xYmObrmBvr/yH6p7y12qXycgL7N5
F3VNEAzvCjbbC/+I2dkA+7Q12vdemyZ6GtblQHdj606/G+z454y1WbtzAqY4
O3xdUNwQ8Cs2Wh0HrVn/Pi2rMU4vYZL6UZmXcRNa+tWKO8I5iZAiUp2qU5ya
h98f+s8/OklBF1mnU3I8wTXEnAo/Z6a9a6JGvR1ZaCn6Jvrl9EH3rgaEhuIk
h/GVlDZchcKrxJy2tCarXYEF5h68tGoihWCrwqMofC+3CVrG7rfbUAwwURaw
IHiYK1cBZVal5nAgfBz0IRD4ofaJZb1djN42P9gBURS99ALg4B/zRwYOmSHQ
qnSboZOvlFnFJaQmfBdrWZSjY6/p1SDzqg+QpouXLetmaKqiJxnYpXxWBasc
z8gIgMQ9JuKqf6ySamMqkd5iy+sUKhngQ886Yqbj5S/Zi+yHLoaq6ET5yLff
AY/qut/8k1XzMo4aRh220Y3JBUs5qUbef5UBc2iRQTWavtQboXfBUloMJ0Ol
srG7uLsG+LNU27CYIc6GYwf78fgfCuaCnq42W2WCWaOdXClHrr3SKIY59yE9
3qe7nrLujB3mP7imtPJlWoUNlQ8dThOeKRuJb8w/GwzsRFTN2c7kaHbzw3/5
zVAH+fsUyD1wyLczPY2UAzPMFscX1J//00KSqF2PtmILpxtyG00BkedIqkV4
QFt4B6Ok//pWCvyhVipT/yerCIX/wh3ReDUaQ3Kxuw1rn7s/1hFI3D1tyYuM
7eESd6kIqgk8qrmtzWfrkOYroKkXVkNEqZTbtIsCTS7XtB43clRphOK7aktp
hjpEFzJe+sdAF8hV8m2yvy6gxikxFA8wSzUEg4mCQxIXkjubtYuoV7H9wODm
CaQLpWkjNhkC0+bZ5FbJHnegv6PHPV+Nl+8DzUSr6uApKJNnAAPPL1UUnz1J
mJ66kMgLy2JZaF24IUl+WuQFZcXhxO7tysb1SpRBoYpwqqpBFqC1lNajKo5z
UWCE+eUuEf2udSLLf0vgfdcOjt221iCYTdqcYTDw7BLyiUqnWAvPv12f4hhp
CvjSr7a6TCbgNL8XMUvxVJHm1d4dP4vPj6v7SlpAr8SIYGt2mJhTxGRDiZPB
x7rYtnQPVdj1x6iPlubKLyqqTzUdL5dyCwX4cO3gEvfF6WkR/FEYQp/NQ3TG
PNLaEBwUmwdj9P0sY0jB6cQcbCQnzmDHMv9RVQYP8QTF+VcJuPG5bMzzs0N1
45PYy5I0UkNvq/7UUlVsZKaJMrAhwbb43W7JDwVjf7Hglv0gMuTK9o8mDxcX
YQEt7ZVqwjtmGzahBTqKUq4yAOfqNCirY4cG+oSy3HoqIhh3ScDe2ILvXIad
lY5QTmZx4h0IvcfSmp/prItxZ+TdY8WoPrPRDVVDznmikNN2Z+sgmGkHkHrC
vtOMUtSjINza3U8WHOVAKTPnSVbrUWoOZOIjrFme0WIr/vsT2W308LipXM9b
l8C/kLbFLTcCWu4hU+Eci/UPlIYIhaLwUxvYGujXxi5VafntTUdCjqIP+JJZ
uoUExNNQLfQqXfurYQQslYyGb7yNL4lkrEOSjScbSRFhIfHvTcJ/OERkzBtt
h5K5QNLYoNBPVQOq+du0sldj7UPlKn8FMsGGI9Py7zuY8FmI2DPs2vrDFfhd
5H98FxoGt5HENhrEDhNRxVAxSZQHL5zFDZnK3Cm8NQGvNxg4giEW/oXePWh1
Vm8Bz3CU/ufk9yxEUNqbwoAolqwvcTmKi7DAMCR2wZsbstsZC9VQEhMeSoht
ALrPROaKux5wRE6DhKbjNb1yZYi32d7PQC5i0smCwCLJD8UtINirIkzJJPuj
/tcHqqcGZIIBowxgVqgKvaGOQt47qqJ5OK+OG/3kskLTno/ULcvYdVExYOWG
SLyWmmArAjlQhWHLXcYyFLgDaLW1VXwRxXw/HMHN/+YKzrvmi+gPYApkUN5V
n6is6xDgdD6WBOi0WBIVthoZL/x/Kijo9gSmNiYA4SBhT1I/k3H6S9MYs/0X
FLDufiwKfVm8T3N0zf8dh5cr7OiY7W+1zJgiDb1tQgA+pVCjC2dCyGI47OEV
5hN8C2G7gkX6uZmXfFsr1VsF6k8O416spTYtZQZBgJjL5ZzUcHV4kNghY6x1
gpIqjlVrpzhcbBmKI3ltl4MozhquYUqv6ljdkL2iOQAOEcL4Yc3iqfbzT1+W
urtNBPocxycLXK3IwuHbT8B+VWH4gK/Nj1FQ+vDRaN3LfG0Rz9TBh12flMC/
+bALdesldleZiCP9n8Ri69jNJZeQa3XNgPJQxb/QJfdK2hhJ3HGR5uyyahUw
Hc+tnL/Z66v7i+Hc7jHZF/Xpfnl1wsq9FRejwFTxldz9zZenYclUYf5gyq3J
CNq/1KAviX4dIiZWemelFwBkpaPuhDxwb/7I4VMyClAbf01sl1V3qq8YeoyW
U3ykC6DeY33y/AmfNCYt1VB+cgvzjglzo27qv+lCygE8+9ht/UuIWpshylmf
Hyjob5kBeSDxryLCqHOcNV2lLdo8FxmcXHkzOasu2ALQzylHX4e0WPX6hfna
hUaMjudU7UzXBPaUmtWiSSzfVEEW1yIDmdi5nFB7x7zy0nqZwSbUSXTmpuZk
dkPAFEcwQShEjqOCqfsx7jUr9KNXX5vMNMytDwnUesG6rllS12JhGFP0ZWrk
gh19ywWDE0nFf2Y7SF2qGWp/DlDCTbPYP7p0BnGyOxoTVAazGiBxFE0JtYjJ
y7F4pDhNn8rB/w2D/tqcpxdNe4gQ1GhkNk3qgqgS7q1svk/E/I6k+l7ekW/r
Nwz47/+hiAADMmU5KXGIFHLs2TJKYSDijmIeRV4DjC2Kp2xiU0PJak2jbET/
S5XNWyCd7M/eQQ5Kv1d8l6LNI/u7BuIkwkq0wu1ThI2CTqgUCRkNJjU6eCfv
02U/SIR/fa2xGpWVd33VT4Sz1deIa+gToCVPVWIPjXRkUztCYYs8PmyJtWPc
SG8GYB9jujqk4SX0wFVVjEC3BkYGta5G5RLwuAHl9DXlaehB5QrxCO5geLTs
6sKNe9jOqYVSDmiX7COHfx2ReVAGS6zDEzR3eH9yRMeORqCBWYrc92mzRUm4
LK+2zwVG+Lt+pS0Yx6f1RttsORxW722oXh7Sa5GVvS/EOz99ltdL1ljyF8Ym
OWfe9Vrp9e1YCKpZMrBuIGAi4RNc+N5kqXiTOF+5jjdNos8eE/OEuosuu+Zj
TZyrle+KSS7Rnlm1jh8MlWd0Rdv2FC/3g5UNu0Ko8sEFApYYY4GSJVS42X1n
wBAg8poZBUXjZnfE8kqbTJeAMAoe6rLHLDvdT6SLzDCCxYcSZ8Q/JwYes1m2
LtwpY1aYgTNO4BWnvYSVgyxGy5MPbk9yuu8ao1TmRIYRJ/SP7Ihd6zgHFgnp
GzSIQ2xggQwZco663N2Ht6goJ3pPlhWGzcP8He+jXqvxf2kAFivobYZEllg8
fDUTJVExjq5ZwqX0Hb9zV3RDy4UzbOEEH9+M3BgXDDnNjr2G3brrZLLmAjkR
xXaUTzPPqtYT85jv/avNRYrI1N2aSPaRTnHUfHVPnqmcokDePSNPcw++6cdR
+TXlRWqYtyNrIPgE5KKlo2gB7n1QyL5c+2EfVs1gYoxygL9QFJXrXVpjpD42
JcjXfpyQoxBS61hdlgQK87kQ7feJs/Ml9iOPIj0H2HHqmshnAd3A6HaRGVbY
WNKveyY6TUntfyMSeNG4rXZQaUIQlMS6kVVOGfUejr7tdLB5gidSjShfH28D
EaXsqHRkQTZciOfgECppe9baCM1sXNKJMZ0FJlrJjk8zfdimocIvvOP6kemZ
D/Tl3j8yNg0mGZV1Wfc8Z1pH8qb6TnZyscPiuXZOqmzQYPkXvETtVL8qQcnO
CFDTxQR6kdZiTUrubGnc0wG4C6LYCammsX+Z0VtVtVTPxXgy8doQeWqLPere
thOjZkabgxlDhpgtxr/5DDvf38DEdtcsAOBxDWLto0YIy6pvCX+HyMqye8ak
mzkBkZNL51piqY/wl53TzBs94q2Pz6PeYDhQPPxngvblzX29ZgAYdTyuSW/k
0Xh8Y0LJWMJagMdJCSk7ZEcyWlbRu14vmWRVsKU2qftJoR59I3z2s/NoMrTa
LUjZ8fcim5L5D4OcBu80eb8eJoTTP0ZmgGkLEYAqE8r5F/sZ6WqnSKaK00Mg
JuIN151h6SpRV4WN/Q1It5C/pudkDftw4Gw5KMAPoxzrvRtYLmgrwnCB3qkD
i3ztgWEh8aJQYoChamKerL43mDPdlC7pj+/5+L6M6IpMOPJUbczCKBCpK51R
AMEU43rQISFT+KUWpO56cjBqBkDG/iQbTIBoHxVTMmLMDNP/2txsiNIKpkys
mmv8lJqEe+zJjV66QlxZuwaTsrSEsD9oud5H67rCoiYXeMAwxU3Wk5Q848lT
sktWWnOXn5qPrffrjd6LDozM3eDmKarepUomQTGsLxgOtvN3ALLFY39C9cep
65iTNuimMWMA/VDe+UrWUs5wO6kU/1QqiC5mPgnUla5dyNnO9RvZfsDSjqGk
u2lPW1n3ZMzFSJ1InOQbfGUWtSMf9Y++9tisWCzzmR5RFHbDBYX59dK0o4Um
zzKXoyoIV31idI2jOjsgOzKqWjVXmAw7TzcC6yZGpvJYx3b5XtgyqzhV2m0u
roXppHoenvGHWGUALDVp5K4/jQTZmCpecQ3wR3LTXZaeSx4pXn6yiPGY0wQU
s/eGe1jV1gDCwrfcPXwaXAb14QbYR3xktMEFFw14umIw6N92LHF0fjWjKStY
k6HKdMIL/JdLAklzU3JhWqqfcpSBNG+veSAHVtP5jdWq3EWi3DL5EEa8i86/
i3kV0Z5yTRyEr3sCsl9FSP0M40qBgd/ccZw7/D1pwC2zBGsrgArw6NlMTBKS
HquguarXlaFah/CVqqXXKXTl0VuwtgQbyspYMYIvnQJzXcLJFtjtsG9Agkt3
YvG56CM/xkz+pSPGONUQnNL99cA8OudgnrOQD42d41hIEEssNI3TKiWYFg5R
UMClcePh6ahuIUfAUXxu3TF/f7+hRJX7L2zayyr+BD16NXccCdB31ka9Ylu4
OVV6PVmXACIZ5CwkJaIg4DZxFImKACpfA6C01YiEzjLXXHISfhiQMdEu2Bu+
dwjcSPgDqi9sgMKmdyrrbp0gM6sEHFRn7na75eoHa9r5D9Dg9KQYJOJPh3Ky
dA2b2haUDyJYyC2u1Kt9fuap936bjU9vyXqJ11XogSdX8jQGJrezmBgI1tWm
mW/HiXym1PABUDcPVAL02025D2B2i8GWiYd1OItmA1w8ahY2sRnwIJYAnp1p
tkZLmf8rnJ2WfI+PYj6mpAG7BZnjeUA7HD8sbaIkiqC5zr8B4iqhH7Hz5fnT
nxq91J3/lSe53D7Skz40qpTu+SDUbe+L1PBvN2owbtQbHW1SGsacqZAbJTP5
9CD4wsSoN1qkFU6bWSdy+8R9GBV8iz8/edRmz0LD+25UJZ7lRD9MM5cRfNFA
EO8Dn5LD56d7Uq+Kb1QpYtkwgIOEt02/RcUR/qyQwlNT1srIRrjqYqYhRZip
t3XbQNYzkiIsS+jPx3DvoKgY/aE+J8yfrR3YYy//R2QH9yYHjL1OAEkasDO5
8dYzPEjRIay0n9emuPVvZT4o7yLBSoKFeiOhYx5M5ZR3v6mfjWTLjxH6QQQ3
E+m5sHAD5e/gTc40O6RWLsbEFtThNMU1My1ksZ9wfxdD54jLj4rNScqVVnZ9
KafRbD5zmisPaIYyAEbc+x6dJTpTwUzzsl4Wagu7Z5D2m4H1OVF1QMInD1JF
ZoyeWP+p+mmBeaRTgXOKOVBflBuErY6ijmfLJPxegPzRSSR/htLRrigt5D8M
9YAqmENEts0yEALfUB0Aes8g1Iw49BN+svlTUo363OgP8VlaQEMXrLxQPbA4
cswEBZCAVxSSBJNEG9zvm2Ruc43u0BuTQvjHD6MsUFq7YQKyCjl3jvqpDooJ
vxpv+5ru9pRWd56NX/tP+yGaOigdnFnWrbvempi/Kpc/hB8cqVsVVxp6wt5H
+pGRnCly3h2InjPqrgQyGEqHXBGaCaYVnz8HmiKTeeGiTmycwTxILeIR9rDj
/P9LZ8gQiJwO/1Rf1TcoSkWZYv5XmPtBHbb19O+ZyFyXVqf7pedO99R4e6rg
vihYMWN9tJuZPoc9H/y6QpB9HcwEstB5J0wMUKmWqNXig1c4vDc8hIYM/F1x
OdPWzCmo/xVpGzbV5+H8I8dKhs1PTSnWEiuV7R3NI5atueTFe3fzT+wubYjG
6ObW55Hy95uY6Zfs6RHx09NTz8K2sMtloMiPwCBN2it0/D9QldOOT36dXchP
oRay7NF4qaEh5wCJ3hBZtukL7qwpGqSfRzY+AsgThGTLZoyaKYpiz/5nZcbb
Y8Lb3JI/MA8tKxRztUCtYpbXOGhExQrMTv5bP/SZSGD8f0K53RSMbAgMjn0H
2guViXwL1FLw7WFFoLCv7vUXHRj90MwmRXipJe8au8ystvb8hz4suD1scWMc
HqluBHLb9FJCAp0nTRmv4j03QrM65LhZCHAzK3uA0a+D9SOYVli1GIHxVqfu
alyrYhNH3jkE67YKnX2hOZ7Nc0QejOGXB1di2EafO9RmxMjflzFhxK5tAOv0
2lISlq9AymTf4itymPSC6OHGelYe9NAJKnfxCdDS0rfFuhxf/ZPk13k0ie4s
ygcMQzLJTWCSyVjcmNj2qtKACAkVo3HJlDpy34/A7N2LDxLx6LYT8KSr2IXt
Lpimp52QKknvOowda9TpmL20s5yg3tlQ719aUdN+ZNCFyeYXnCM5JnvdrDUs
4ektz6C6uark/2ikiAHqb7MUxB3ZU/PTD6YPA42sspXVCh9axAOc/SZuGUfM
cDbAQ5cr3oQiWgQ+lLCS3KnEPw1bBwaOUM/1mlyZykYC4IIlqurMVuAYm1q3
5IqP5LkbBMCI8P4eSo9z831YULoX+5sX0CM4iazMRTjEIwuXRZwiePiTRFu7
/iSqcpHyK/XM7713fXsTGB4CrNHp8PwXDK8IoLfrQ8JdI4Rafc92r8enit+/
TbSGE0XPVvjFN355lGOEEm2nuv47BkTa0L9vckr+RKenTLzoCxl0Q606FitK
YbZV2ZZCGOKItcR1tyvcMPD6Ybf8oVFX3F+1ySYzE6Tosft+EeJFzi59v+9L
TL1aDpMS1XMYCEwZ0IEZawzumhufG9XhbdBkZ30Jp9uTNR8qN1TlYBdnaBcH
QsdcipIKPVQ2naFZQ5mmBBZ1BQX3MQbhx+ayTE5BFcC+C0ctwjirpZubs2Lx
eNIuap3sa663fZmGb4Zstab9O2WdAGN3K9FeMa/intJtYYbFCaxbNRTqsanB
CegoAPKAWHyuGcpswRbArK34GIVOXt7c6A/LULCM4s4boAcen4IkHgEOaG9a
fl/saX08Jzar92NW4IzwKurbMj9j1cf7K5DQ0k8+6RST07ULfHmZQa8zpVrb
J83FnA75wvd3iyUZHyofQ5vLKEgND/JVl6xdP/JdLrIbHbsJDZRuYM/MLVib
RM9dnpFSaA13v1rKJksFONGnU6X2Qdclt3eo0pMe5B0v5E12jUkxUJA/n9c7
xO7j2e893Vyoyx0jRGoGC9akc3XLBhi5E5ODrlbfCXL4x8rnspJYHrtOPbPs
s8QWKU5sRSyMsD1vAwoNqBhoeuHtgIILDKmhyYnUaQZ0NfWQsUkgIgx3t7QH
q8SHUFoCHModLPqeN+A8yM5CMtaOWw0mZ/gX8dYCGsCvmv5mkEzCr3402rrS
l/FvZATP7+IApxawMdwH9OxoeO4ara9ZRNNfUoTTN9hXGtsCgsmhPdUYY2AX
3aXmwfUd7DQIv9AdH7mrv3WshVanqdhg7gHUPPNA9rkizFWtrBhXI+pN7MYQ
q72dEvh8kH0WlPXzBqQ9weHYKM7Q4pdD9L8HDtmA/FxJ7+CDdCTBVxIR0pqz
2W8xvEQ2XXMh8Jj2tZIzQYpSf95G/w3WXM624/RVv9vXp+Oq6xuAV7e6Whff
VFGaGQn1aqAF0neBCamxSZ6dJ0LJi/6XrLCbvD7Vhx/X5Tulal9Yc3CSicvz
CLm9qFw0AG7bkoFVWBPTL6UevBm/u155EqYLTj9XilJFl9dZnDKn8FAxlrHJ
T/Fvk1W8MtQYtW5+1DiZp8alLNSvEVCRPaW5D1nEaxzPy59fAu6xYKLYX0tc
ZRvIC47wV6giyp6UsmT/Wo96vLiyC3dIqZBtHzD4vNDPE1h51UUBhNuiI2qn
C0YpPmV6zr4jb1YbkvDzRqvr8RIJ6xvrz1uMYT+Xo1ssR3BKf8QeuTtSSGTt
7TajJfrJ5sDDWqlVGWEI9JxpKtqaHqcOYkshexvboD4YaOKx/vddJIC0YAvU
VoG/GLlWV+JVfd+mA2SU4edO073M3wYx6t4N0jLuOoYo2Cwo/VBJMw8AL1VR
Bnp52ZnYKVAQc6EQesxI8+5yY+9N68Wnrg672ofPNFgNxDq4FI0+0FDblDIq
3AZ7HJfBvnovZD+IyOTi0tl5vbZuKB6HQ7M9Oi1yawvRsZn5CAV5D/sjQ83d
i7ADJTmNCmOooy7LnGfLjkccjh+3FeqkTtw3x1yIrvm5nIL4nvujpqWxlUmy
aJ9yQV+HvRb5XCrORnGyrP/YeUuxJJ/uKGHiw7uWF00UcURbdf+p3pLCDVb5
D4yXZ1+Z1EYjbJgiNo8GUAnHv9P7OdgXJrliz/q+MGxCzGCgj1pZIyFSlP/m
JBPhsXPE4E4MlUEBXH8A9eL5iMwH6e3jZdxsPV5DH9SL0NLDfAjeRxJAiE/s
K47sE9Fz1WTIYKbI/+vLPX/WFEoRSZ244/+Zk1BglIh+EYlJhQE9kskSa2HT
bQgpmVWi3qxY35kLR2xYan+8Gk3unXAG6Va+WAOcP1OkmRN5A8TWdEyNKsLf
xYsyDQOUSOWBOG4Kw3f6bH1YKugMeTYrN+rOS8EnzLBo5fy3BQV7r9RayR3z
VbbwTUmw0R+46lSFzu5vqK/zYZcsKHFUC/3AIW6CNMW1LB+V7W1dnGrKLAew
TG3cCTOGIH0DcDYc9Ny3i5kddRGbubB0VzzYYKUms02nzsYAGaPURTKSMfCh
/EMuQYNXE4BJx4y/8grBZK1OqK9Uw71cp1mXs8vxaUe5Uzlom1HkCA4G6S/w
3bTW9Osg092tVjNew4duOGQBixfiIcODudFDKeMges/nTpis8CEKBp+mdNT7
KxSv20pug5gDw83tdGmUZh2zXaWCz7MKZId9SspTIOcvoaweSjSo0+YohOZJ
v+qKsojg0KfhCW7M3H9Wtr+GZDT8AcCdaP5eBVXQhaxVw7Ch0C+2kObu6ibe
q5pJSdztgZ/7e3obwdbcI+n3A1uHQEnaWqnj1N056bT4anwL6CzC4T936/Dq
z0GJp9FJ48tlvmSujfhtwBwum8i2zEcXxUkJQhbi0lb7McnCNQE2Q6f44/pW
I8vXhnpol7QU9GAJh/lJfYynjt38NtsB5gOHZuhGcHkGuCtv07y3KynlboWB
QOVCR4ZqG4Wc2JNzk6HETqT+0NGdfllK+Uq/eVesnxQ3jCO6XoWCNoRPAdcf
NdApcPFHC56cnGD/ceIK7xId/5MHlTFTSGy3KDehQmX2JIn3H7rOjqayUbKT
ZbU+0JRqEwrop8YngQ0GGmqdf0EAg/puLmaK2Z1QMQN/IKAMSlrmEMqW7gzG
PJ02f2RtxR6xPqkmj0TpNCrtvTkpDf2UW7vvasRWHiqAJGLrbSK5cjDqR55k
y5Q+PBpcmL3cgMUIKAeaj41bh9XaS9I1i7hqXOIHhYYjNXOXilhBpSHv8TQy
zfxAbHLt7bvjGCkiBySxzYEFsSEi6f6CzA/2l897Lhd+NKezThK69cRMx39h
GVWHKqqyslq8L3qGbOzcixplLCpFIjhP9Ajj+RkIGFC4RNfXWa6wjUpFLPSv
qRnB8VtTu8xPiax/h1+V1kCIchVFtgyms9/dPIpUpjDT3l+Mp4p8/6dGQeKt
HnURMK7LhCE1xIKitglada6tiUkzKV7w4HrHOkX0dBsd6WvWEEg+a+/IXlAo
zSsK6HpznWTAKg6mHR7IKKkoN4UXUV9vNbWl4cd3Dq5M5DNk1Jcts+zJqvbV
u3hIo64A7g4/8liGsHOTCsm0pgWX70UfuOkVpSLsjLSBwCkpUR+YgoZ7Y13V
ASQEFZu9a/RA/2K4VE/RpGvzsoEmydBc9DM8nmybS9MGXdFEtpLucnuDqS7S
6r0l/uGEyPQuCUAiUmk/bQCumrdGAyu2FWEDUNtMGBssUM5jiKHTTAw6Dgb8
osx4B1Lxnz42rt/Pj48iTzzWNe9EGNjNrbEajFAYohgJv1R4lkktsUWIHy0J
a33pKt1vO2eQiKmaXS9OfUj9n9WyBkpl+umR8dhDX1Ek9HVIInUCxrmEjdzz
NuFNg8HgZ1KIaB7QVEG8/EvLgNMSFrkSow1y838+bXyUDCYi+5s3JfwS4Snr
dquLA6Q/8jL5s3QtdnjddAfLkIFMbFJNF/7xqAYjLS+QMI/ME5MkeVB+n5u7
2q6hG7F08Q4+M+BUAB9M2mzxnCGb5JGBSRQwV/Q+zIt4k7hytgi0jZjfbUJe
nz+f8m9EUhCr0cdFYEIwtFnfWKRcIWvIPYwC6+PPk9IfHZFUBTh5/vhkn8SW
6x2KLTNQphFirHZAVrZ1FkZ35L2AbPHx/rNfjWK1jFR8MiRvzq1bNNkedk/z
bL2Boi/AMNM557+onaUvrSn5/6RTbKW1AiIlkVtnaNSL3wIDz5p+HpOa/0wJ
zR8Dh8Oz6LOxZffAIXJt9AyNOgtPLdPCAerwnpOo9nZI7JY9UqGL1VFp6Shg
jD1Nz9McPBskfbA0fafo+6pda+M1rjW4F0GnpMyqERNwOiY9WKpKzbaOQlwM
MpVbz5Wdx6knIHKEiyonqCbaUAXJlD7925Zp+s9bzPaQxUX7OKirOg6JHt2O
NaIkWacV6s/jfoperF0sFYjI9fwXXMw4PzrVjaEQ8Rx/IdpX1M0jrp1zrLYV
pGJBy6yV+KMKY0Ru1fdjO06SwwB+0w+Mx0PLzAMy3WvC69ppabR4JgGRVZR0
qw66CVaM6KyAZyy8dof05aL3RiSVm+nRTute+MwSn2gJ2+5DlTSAbMa5Ci2m
qQKYO318V4gcSX8KccXxs1YDAyAc/41rOHlhM+wyEE1/uC0oMAwRitPH4mDa
plsW1N7GbXSoanilhJuFjpTZuFdNXrQ+S0eKmOdJHP3pGZDC0yPdHMIu3Rs7
VauSV4OrIOXU8uk8t8NjxTcD+cbR/LDOL45d2232ezX42NwZz0frZDCFZRdd
iSZk7LfhwLzW5PxH2+zARyl7aWyccLC88HfkVH1a2YWBCVywkrbFon10nNh9
dDAe6FoiTROj5yUunAlS1XlMc/oB7iqTitgviEwv+SFgQRXmEYrX6U3ILfzf
ra5dhe1gbUtJ38K+RzA74Y+ZHXDfpV7ctBCBwr6QkuEVLwWGs3+ltAcMuMSB
zzyMqaoWnW21Xt+hZGT96Pwfpv4GqALZjKphXJDGtaSk0dSzQShzEQ1eBOxM
Ji6p0L7gSlBXJh8AC/YUrgN+IOlVoM+fKx9wKJFvkfCsT4if1uNTHZjhKbNY
VZ52IFw2P5XPSWU6x8zJqgTRm6OR59QercrdyiAIWfUciGlrTbDtQzR3yVtI
NMBuCRjr/WTiTqt1+8QQKiaXFU9uzYIChhXAndxcdaVnyctO0TnniHX8pxmz
iXAFbsWup5j+j0AQtfy67IC7Cvv4KGaqGnj8FDKtEzBFJRV7fPTT1fs33C85
kXuVzf1x8NpA63dKO8nRmePx90BRiZNw/NNrKkiz7DrtWAqK2XasETpQA2SQ
6TKIvMri90ZR9cxukjLoBpwI9BpYy7SVwOuOREK76tTpxXP/tB7qx44MZlGd
dZWO60jRlULsMsQid2CSfy8CL2+FgqVgjoUc68SGs4SnDEYtfbH/P7gkWifF
CA60JHisaGkXcE5mxDbkbQ7RXhlDAtRGGUckBwvRvZg+rMcGdCXuEC7Gvfrg
lU3hsyAtIk99cjP2IqyoJGl70NiL8bFQCr19BnwT2pvZ+psTBMsUMIJKsK+j
cVEYBQL2FQ6WvpVICt+MFhS2MqyDaMJhH/uzetzg2GutF0BqqhTVORFCd9m4
zKH7OF2aIjL+0coB8+ug8rC5YSXynerp1YIY3DtluQRa9wNW9cQ/aFcJREeF
GAti5c3BMdnvQ8kaX1eFt0Hib5WVD+IsRB96RWlzyU9ZHPRgyUXBcBlVJ/YR
bJgQ/ejlF44HHaWz9/8ABdPfO/7PUJZNly1orAVob7wBMOLTw+mh1oIiKDlH
1XaAvHXPICjuuisFyhaTwX9XMI74XPQGyg483VlnkH1VqWtE2HJMaZtUGKE8
DAvU8V7wUlvVlmu0vVjuwypS9Mr4M54P99k45wHvEUWda1PNAizKEVLFFNYT
Lp5InDtfvCZ76CCiBh2EbkG6j1HlwPfy/H8T6hz3tg0RubBReYKBM6Xa8YlB
r+MMT/szeVjw6aue7CxRgRLseybZjt2BJ6Q1Vb5b+uXiR5b9PVqMd8RtIBtv
GD8TCkPSs/4344sm/ejOCH0ZEVaaC6U0FA3VtvSiZAu15wnZhirOEYYjTffg
d0opkOW4BvH0x9iO2o9+/DBhMQmX01cQwuvtlZNfiOXTvtMhAMS6PgSNJYiW
6wmc4nKK3PHrAP7AL3O9JT0tvCMDhzUFHCjWIMFmR+Tn6uIy2EPtbH+3PKow
xUTlVr8yjIIVr1JtUVhVBa7x+MRts8yiVHevadHKzcBUx8qiHqQGaZgkiI89
OP6HY7mHMfCPxUZzn3ClnEBCo+uB081vxvTvJo3qm/Hz7Ia6u9thlnUuOsRm
iea9IOQzsyzOo0iUUy9kolG7m2XBWP73UvIBFoJD8Ama+WiyUNmqk2y5mpyO
ZnY9Lrpw8bqPexWmz5dNkMH7RWORyjIsQ5wKqY0V3eW2L0ndQZCGqePttn2a
k5ro7V6hEfGqA6Qd7+txDHQ5XUln0iUCphc47Pur0cxqkLXJI5+IKWcMx1a/
bT22XJri6pAFI/bbZ3ReIG6/w8KQzyU75LTAorsYdZ1YP7+ZietNDE6ZvzLJ
n4Dee42Lmg1SD/yS2vm1dvjjAwo8QMVykpPSgnxgpgM5I9ONJAIjnyg8j87Y
EXI72aJ6qgCPyKNFfk7loRQ+gXAx5gEdosbDx1a28jM/uFlbPYYjIwASmm0Y
jZytUrAumqW6b0+/c3yl1fhW/TKAOuN8qKt9MjAHVg9EQponCrBX2tgH6t6t
w8j/QveBa/6X2U8P1Zl/jHKPsbes4ZFvkMiLBP9s3XdzVYTGMceW7ZG/9Gy1
rEX7cyTlh73Q00FD6IFAegArL18j/W5aDMw1FH+EJ584D0/ICB6Qky9+uSeI
TsI50zvjry+yvRtndChmjSFQWjVdg61ATup0THSzWZlOHk0rDM6GGhHPbxHY
s0Us3oHHeaNIBIPNLiqDX3bhVdvOQJ9Aq5wExo07SQWJtlr2zfDSHPWHpw6f
va13ECpAPk/E/A4YAcl0aLx+tUJ+pni0M8Oj3X+t/v6uIAQHulSJTzSw0kgq
FVaSM99scAAPtUuWRcZowKARKFHzAvfSpVU9zRKMRRidm5jlEoVnFV9RHt9g
kqZqTOJQ94mpl4JmosG0F5H7zOwVus2+qbCv1CerHS7zWADYaW+QabpEejXh
OJSSVAQV7s6GsuiZpw4wp6QoFFzhoZbtGE9H0LcmFCogrnSVloi/1pIidE1R
ZF3bf8gkOQnNlmcje6KZH99Ih+j3v9B8+ZbwZl0E5ifRKeowQ+9DEfuJWWqf
ID2vZcqd9w89ACq+ikwHOQb/SbsglBqmPdAnTlurNLlF+LH3ixcXcSavqL78
dUrN8E/h/nQsTpyDoyARJ2j8+VV9vzdhsnuX2cokYZxXPp2VWkjpRWGvPpxr
WZakc7Y14NSN0SkfAVj1AIHj2QXiWtpLUMMyaMiMWfJiRBv34cdxzdeam811
m9SLEQys7vCjO47jwkoHIkal0Rf69h3bOoWUMfhUEKv1hBDwSf/DgYS1Q4BY
6N1EyUPp1ihfgoYYMrBHuRemD9liYUmxZwq1dreG6dlLEZhMQu/oaBrnagQC
li2XlHT2YZk60+Hea8IlClBF0B9kZURawFD8+BAG24ZiErryC0Owav2HhZzJ
E8gioPxAcYvNQwkXLNvjDlBpvqOkbgn03UgSDW6lwxz3/6yxXALqXYJOODJi
Qm768tYy7XTKQl+bX5DVgktj8lTE64tMcB+oYO1kZwmBo8/SHhgbAvmCYh2J
BJr0hDT3xRPDJXlwWVQoHVE08K1GIVluo9fjupShsMEHK2GuFcqlyP6uJ9zS
btnBnve3vgeeZLx7FCWJVREkkMDbswt8bogh82SCRvGC7n47quBZTS9Pkt99
QBpt1B1nm3FLJiYTa0jVXWW+GJX72Vn5IkG2ynFnRix3FCpiYlbRzPfg51lW
u7M2XCCt6s1pvrgVMFN2yWJ2hET3EXHfYvvWggI6PN1BmOtnW6DhrxF84uFc
TOVuEOGgXwM78V5bVa7K7CHpGh//0RtNhArOSSWQTIJRa7t3KvMXHr0nE394
U6tDwtPVWoM28ZkmqTp0qwmbu2a9vz5TJDU44eqJWLtE91TrFaUvr9yEYpNo
QnZPLpqVk/AdTFfT/l1fNCq2Hg3R9cNQdb2LqqkawxBpTnArYhwhkhJMAlS5
t45fDsvsZA7Rqe7Q5+hYRjL6bDvs+EX3Pz08GSemYzNU1mYTYTprggEVMlzT
bL4GTT4f1z+aADvLSnvgc124ICjQVdac5t1HwaIoWW01uUQmNj6/TrJftyUC
0ALaxdSjGUX+rxf7Cc19lFo2rgHrr7GhzMIM5Bjyx6gu5IPmVHU1N53RuYzY
nVhEgB8qnN7oBnuBH2MPbOE5rmO/+b6QRnt4pImb+ZpVxsrkrB2EsEumVc3t
YkSNc/T0tLWUy2dySmujOFT/5CvkB3KidDdiKMpLgkrZ6LZwVZh27b84nmUj
xJDxcJSbvfTIS5xHoSQUAZpPKPHR0TAROy+3pY7rKAiq6Led8klA5RYgFFXi
YPUyZgc55RdA0V4Hs3D4zzbGEZIGfUVZebc5ScOZ4CFrBaoCFGcow0KMugKD
3BZoM0ixFT6LjtRD7vLOjaO1CSveEgZnJ8OK1BgwlUc7Fg51kubIN3osdiwU
r9DXeU5vc3G/2lV6s90v2lJ3jrcCzDzxlIt2ZRNRA1ti1WGY7LFPQFGxfcfb
6JfOUApf0ReLbxZpWULc23gSWHBAqNc9W5qs5s+AhoK96NVfBQmDKQ4fcNy1
3GjXkbtEvsAG9FVWNYND0vrxq92AXCSCXMsgFKoSXDC80q4q/RHRQvO7ZyVK
Us1G4/mQov28KBjzMlzPab6xi63uF7ZwjufxZbHcAonvCs0fy8I3fhF909tN
Tb0vZwS7/X2zA9mrK5oBMmf39Rg1wmY4b2PqU2g3+xntl1PJCWu9pgLAAMAE
qVq85FSp96U60O4/msIeMAzgEhxrrTwq8zI0XxjGDBHdb38Mb1ABirZNrBxp
dnqv/H/HktxdAmILQDk1RE39qG52Jo0IUpxfTvkPZTggkVImqI2qA+hToxHu
rafTfhqGDj/jb6HyK/yCK0EJksUYvJVwOO6bl6nIPMwUwuBRf1VAuSJD/d3z
mAtZmdmskjJeGn5kTALjnYYRQ37Dek5g5YuKiW+w3jjHw7aNKt/JoUVsfWUG
zHNGX/1RCtjjOf5dzB3R7Dg2SB9Uw0faf4Gv6vC1BGmlYV3c7/DSEmRXS8s1
vgDHhIQ3XwTFCXiySBXhiR/pLF/KVpM80M2srec3Zi9Sq3fg83uPxie++uQc
xASBxp4RukujRPd2e1Q+9xWLmNqWdfp+IUuMEwflmz6LVkbPx/ol6abazDif
DZSqEHU0qTbVxDuHygvH1vRXRnyvAuve2oBVgiXhvuanHKo/mBFf12zOcA5R
bfHnYxmn9XP4mumMMyoBqD1NRJcZhC6yVan4I6MYE4079sPKx861pDEhRppb
AHw7CP22fQ9e5mZpwTouGGNB2pu8uo5RIC6uVlBtyoasNhEga1XC8YdW5Y/T
qoNV3WsM10rpyGxpgxkrv36kgA1D6snEoCpmlE8/6+8Tb/AcbY3nb8ogPkXA
sGjEJXExgiJc6UtREP6Sb6hTcPOfmKJ+rSX9s2dcDSLc6nZRs3qpPBvTF1gD
LDe532xpAr79zDI/ACxNshhIbzcWgmBc/VNht9JaP6zudnUtWx5EZ5sQp8cN
arI05UBw9seuiTOT0h9Y4A1Qc/F13xNs9UiRYOrK8lmFww3xY9PdzdM7q/Jn
/+ABCQ+S6W9wih93QOWxGNnCrk0x9aAc3u3uap29ZRyahd2Ej03GZP4B9JSo
D1prLbQjO3M84OQzyWKH0g5PLiwxy2U7W41OkznpM/VrqFSymkdszhFbda/A
ivsUB0yvRD/beu16SEyn3hS/QhuBHiTOQisxfYV+ktuw9/R1/QYoBTPAxyIY
+oVNCthHAlrDq9hZHFpjtvQQdgiRBMKs4i5yopc7znVhJqqX9nqerIrsMc8U
lsLn+06IcMDtb7jVyD046yyMKcazq3VEMhXdLiCP5S9UkorVsmo1SdzTSbfG
A8Ro5VpYnHndQt2NXdnUg4LmFEtBrX83seF5raIj9IyGEMmTzo2CCjuhK0uA
Gbd7ZbP+zdVU/qjhw19uax3bMsC4EMV31OTqJMJUfSa3B/4ydGFFcRua0STQ
7ZZT65GK9EXtzVqW3ErAGgul+o0moEB6N0fdqvjkO6BdGLSVKQgA+AYVspk3
VDp1uuCnKgUOpXvku4oDI4HIDaki0eIRGYs/G9u2sbJsSMURkmKHwShwadyb
7shrHT+9HtmV48BUbJ3AmC8t5DcDLEQJJ0pV4ve+dZmOOzOo6Q2kLIGiCx12
Y7JvCdgrJBW0STfKoAQ6/ywymg/XtMcCaKj8neck5RLg7MdurlY5zLYu52ig
lrNCgY9beQT0My5yXY70Mtr63ItxpM0a0NKI2YgeT5jAB2JuoLkNASR/cMrK
xBDrBjvxDbNI5hZYR4Q0Bcys2H4WzkHz67PrETXTw9RTFx1Vx+3tHVFqqJmO
ZFtFiz3SdHJ0V5zQyIWxkdzErwKgUmOaMuglv+fCt4mGGEgRHORiuBDPH9HJ
JzdAoEK5T+gnDJfbXpNtQ200NEXQO64FLuxL0jWcKSuHROB/NM1Yve/2o1po
H32/H4S48jSGkiI5MXosp62jQBf33XIp6FYiZEeA/OMBHZ2HbKLJ9bldChx2
8NLaDGefryO72V6oU/hPpQwKI50iICBSBIYS7CSX37V1S4BmuOlu1WI+Hngg
hyjgE7vogJHTw2Xc0EOiAPWNpdxkhzO59Oq7a/KWhNWXKuiWgVwVxzgRRbq0
B4+e7Qr/kiumng3UPX9RzzrWAONSAsEuzVWHbGRLt1FwfQlzRv/IIOI+iAEp
FDdSJVlhBH8UE64ovYx0rUzrPMEmdN2wNlFfmZ390WJJHnLBh7aKP5kGLlvl
AxBm3sdYc2LSW3fBgkk6BJyESQDunOnc6Vfa3WKRXUAXOb5RnZfEg8eifcBy
5W0C39NpKsbz1fzP0nqzYO6Q1/4tX9DmmFCGzUi0VKeOu5d6vUR55S+mnny8
D9RzSU+NgVIe5pbnw1bZ+C+K1uYJaRgJhYjtC6URnPgWBbox3LaE4SdYCtvk
J+8Y/vassknhlBl01pmJ9Vv6b1b74XpvT3Gzn4PyOB+X3ldSHDiPM/VMjp8Z
kof255+P83sEOMwAWvUK2bWciTO8z3TNn6VyoslpRmjmjFfXWiXw3KWdFZRS
AKDbo1RqywVzSeWSebmlIsk1GX8aNA87LsSgJvIybKLR/KHJVVtQHIUBwvus
77rxj8NBG6pem1FxnpZ0dGCpTdoggyFSBLs2WPLd4G4WvL/2QkYjeigCKagl
HDG/p4xIqHIXx0hnVyI05l0Jkua7XsdnNOmTjWdxQlmATX9GAdgqbbcgrL8p
YwkmjyobzIAOGWvA/LVZnOugQeQxJc0+iJjsjtce4EBqdzFEqi5Q410CimGB
rTTB+7cvh5lbhvN9iggGkuvW9P3qorzFWUiv0XdN15tThvnGQ0HAIyfBktiu
uVzuMo9OZdqg3Qw7+rZqAe+0nPMz3ugvlCZ4zFWxHc77cZWrmExv/M/o0vGo
OGW4nWzVfOlW/CViI/VrbUjLgvpXFLGIqHv3yHzv9oDFaPPzEgK1D31A9ewH
OUBkOxKlZQSAvWr/EZKIfeCnGm222bmYCaNl/8FDWNoQAiJl5O6tSr8NCElm
52S0XB12NQg41KWcrje/MmsG8HwKt7fT6rQr57IrizVo9Oaqc021cehg5bB+
fib89mizV+VzDEcPzyPIza70yAwmiY8GppGpe0VbUrAGln8D0b39dd8Afqld
LIVBAaWyLIiKMHuzPwkOzx+o8klk3zXGhpn/bXGtf8SujmpH4atly+Nlk2EM
rGFaZrGpJm/rdrtFFT1ZRW3tmUb7Luyc/0WFzJdR26XoRqO68zBgswVJG691
5mjGc6r3Uu/Yvsd/SnAEdAnpDRaqqZQug82/z2Cdjn4vAJgnyxxuKc2dW4yi
h1z514lQ1/VNPvTsUNw5NFlIRzHtoCkkQLeFEItyINSciBwpQe5/FtLaa3HB
fpY3sM0GaTjpJw/TxH14/AhTd0ejp6XZeBLNu85MZcBlyw4f7IedjirgltA+
VVh/DZvXOW2sc50yMxXdNTgbB/loOT8hSyjIg3Bj/haQY8SI0d6U+fRTaE6W
hDqZ245zw5TsiNCMDjNcY8vqVm0CYr0gLiRzGGdg91PWuUMCJNmqUaww7Zko
qKx4b5k0rHFQBkNnMQ22W/oIQTeoDtrzP5HuRL3sUDVwFxMe8fLwQVQ7pb7X
Bbg1nUwRECy7i8pXst9EfT92M7ScEF9oykIoOIKkcswZtQNxMMWvya2r2y5s
8lUr3GuZ45XaTh0Vn07tiPWj8CwsnLIEfafDya2G1zUH81WAyyYRB0PjjfpZ
gvQ4xb7lLcGtpW59EOiX7peyEQy1KQzPyx6YFo1OEF4IK/oop+S/7m/MhevN
TgMgIB6yh32ZByluZwpiWBC8LNHb5InD8QIVS6HRbkOUuzPq+am4sdK2Gsh2
mY0TwOXA4xRboVsDPO00KvGC9d0Wm25d8a9IRZUCfk9KaIIHt4t5xW2hz7Js
NqLt6/Wlnh+3GwwcMOUYpftPX12wenNfiiYKAb8HIWPHWONsQoko42ybAx0u
ajSOdH7+aAzEPvpo8DzgQa0NYYhEbIWOuKcmW1CpflsDdnfJoF20uKq8+I8h
WtvnSJ+6RnUXfL6A7L+5NVATh0o5trnY/IlY1dSM5Hi4bpPBwlbUe0H1yvy5
ufzJjTIdeMupWexGJtz3F4UFrD3xw0ki0iudXECwxfnPBMeIH41TQUmUrmAd
QY2LJYQVr4XqM51wxzck2HB1qsAoEl5orV7xr9tHeWc0qQg3KTzQ0a7XH/kg
1BYhPV/qwnSs/Rh5mInNaWo3P7+8JZIt/ufQJaAEs8h7XOYkWrEMPj3A9CGN
6P8DDyMZry/Gd2h+Qq/C/L2NbYCcFWJav9Wa/jcIrPzeaQxHdp2a6zyrqppJ
hzmtQdEBnF3Jmf0bInvxakG89/a1EYW2K6ohcPJz7id+7pPgUBBs9YLXMuEI
d4wKHXM+1S28kbGiQPsa4EObSEpvR0urwMQd6Wbg6aXBG4mutSd6jFYs7kNK
nOlurN1GFjHRs+KtUuGiFXcMs6M11gefENbnZnyi/K1Bl/Fh3ZZQ5mqCBPTX
FT4U1qDU/xvP1FbkTIJrm87nkFMp6OUBzFfF/sG9virtualax5sKdfxRyhjb
xt9Yl854KqvM7bqCp46o+UrBV4G7yP2eidLJ13PooQ5E5X1tB+s4egW6h2tT
WH+seenX/KWES3Ngs9O8kq7WrEvKJygVNtqKJ7TM+qh1N5MCmfVsPldh9Zjx
MZgcoi7THXeoFSIzA1ZvzdM5zLxEbW73UhsWayn5hC5LoWLmc/aQptNK4fvZ
3ed1HioeulxKJ2bBHKHxGV69fMT7BrelkhXDpIAPpYs5hJjppL0SZ3yvBAkU
rk1id/oNkJvouez3lrqBFY82yqcgmzhQStIu/myFpnAk2ywRGEuI5IpUR+M+
D1KyVnzxStBMMvbtt8qVqQhmmwBma34D8L6m+RvAFN18XD5NEc4/eCuoP9rO
K/uBRdiCXq2GFYBoj6grfie3i1JxmSbCAT3mMCjJByxccpiEOuGIKFJJK647
X+urY3knq8fHUTa7dGDIHFLxyFzYg9j2RuXQ6UBXXNq676qkFY6j0BrHQSUz
6/tY1xwm2tJDjCRXZGffWPIOJQURuW7Wm/uP5LwbFvleJssE/xgGPvwyTYYG
J7AdI49SEXXTyEh1lvPmnbYgue5HCfMi/zHkDZGK3za/1Rx9q0Lj/SIY++Dz
L77fDdQlQYWnk2N/yKTEOa/2kZKq3FhCH28ub1oKfcrqHqo457IRy9JdW1uZ
fAcBWu7dWQXHNNbwEaf/b/2FucdZMBU2PZLwW8Bhg9RT9pshIBj3RvEJYGoL
ZvTFodCTmAte4irkNGZxW9X3WILCZ1D9HwZJ0Fv6Jp2qez1N3nyLSSBYSK1x
heo9HX40XwOeECbJQ2+GMMR8mfTrLWsqRcolAt+zAPWR84Vvd12mY5tEajau
XR1xGc/unzS58gdTdZzYEhRpBGXUQdnf/bKcNIFdA+uf8exqjvIGstDsDiJp
gMSq171LJ0FPHrtzdMgg/NIyaQqCPyWT76vUpyMATzYaSIzjET0DwtS8l1IK
eswwZyccOvWCyD7vO/uCQ+6FQD/4436gCXi7sAJB1vRoxS8OgojlLCQenuzp
5gZ86zcYeYamvvn+7PW+p7GB8rXyRudSHSS1V3QuHFQej3A0m+PSRh2N7tM5
g0WqYdBfS3nk86duAIT0Ry3mGhkarL/yqMAeQ9RkA+KMkpRRmH93Np6BYSY4
46xs2XrPYM6npThLvlFRRMEDAYGobf8I8RQh7AeFHT7ibVLa2ccVb+WNIWSl
sSfG6gkv03/Hm1THpbsFLYKR4iJPUzEuH2Dq01jWBZsKVz9oO5CpMwGcavhW
wqMXNh773MdqwMtRgSc/QuL91T/Geai9FgSR83Wpf1748cXZO1mw9qr5QXmR
22Zw3FcEDwtae+W1OTNRPNT8s1Wwvp+eG4RB001UwDSXUFkpFTmDspgaHERD
SjzCD9JvCfhmT5VQZQihLSRfrXALuW6TeGRyYJM98Rde0UsdZZmWP9JDFfQl
uNSxo4uSsPPoDEfUCiTY3UOxlNOWqA/036OJ4mYgJnWu6937OfMQknmAQOuT
X945CD1e1VdQgRXikOyXrV3tFkPXl023itIk3mHbGbXDs2qBybByhHI5DQxY
efMc4O+3lL74N3d//aKbpQU70ObXVO2SQLYFDSgpqaqi9uMmX8WwpCBgjLax
i266axRbYlPz14et6FQcD0rXSx48xlGuU+OjYmFdITBh34VFRcK6kIxYuo7o
pCoRUlaSyUQNAOiqPzwMejjY43uQRxvU2ZJs29urk05ws9Tl21P1wO0NyWHG
iQbs9gWjpEoc4joDpbkh9A0KFs7zJylf1hmXD4nMEI1oKCohIotTWWmvsWRH
WF3Ar5nYR0MdsW61wE5lVkwRqyI7WEWr3YU9WBJkDbTTE+ildgz9COy4pr05
UH/5VJimhZs8T2ZqYJn0q4UVvb4omQoXLQSLejQZezP4ebngOEIm/hVoBgFQ
jNma+4Ut8A7C+niXxV/rRcUOBqFf3q7BvZQO28VrOl+Ubct8hHFtSB6YwOJ4
X10axg1oDAP27T/T7ShhjNl5pLdf1dA2zQAeskrZvkKOdxZK1v9esyXebUIh
zhOx9rQ5HO+FpzH4dR/azTeONg/GfvWeUnBhZL6WVYSfL/xwm/Ct7f6226Ik
UZ9dtCfNN+b0PSUYCGRtY3F3TRE0ZiEiIYC+tuPP2lSK/5/TcICvaIVQARLu
ekryRQyBQaOPyU344yMcVCzHuN3z0XS1RYSiBgbAq+Bz9dAs85nNOWPmcv+T
v9lh0gHUqv32v3vx5O5eAR8Df/M3Qsg2OquE2kgcwQZfRa/IUjcQ8nbnGmRh
e+Qm4R5cNztaip/6TkcldsWqIbsGfRVhr/LKVKGUvDJzSM8zNApTqsGjLZWa
IRWmENiPk+hMZwow9YFoqhshGY3eV/UZqyByQGARcUGs5tkGHY29/lgywlvx
hqzxqrc0gjV4C3sUErc6xi2LKVqNbsUUpYLgIvpTBwDUsNkYzYEnXyjpMUMw
AzyNIBsZIqmDuf5hMc9EJQ4IQguNiJnpRulWPXRxuhqky/bTCRXpGr/VMATC
KYnPEZTez7pCWLZgjy/hRy2NLrYqAe2jbS9P+hSWa7r0mDuFcecpnP4PJ/9S
JiMQpY55dyF9/KWQKWwkD+TQocznjz7kN7nuQLPmvGUf9InFlmO8LzxqHGg8
UoPgj8LyWFr08T94ym3C9gZ0bQKp2I/IlwTRpHGlykgLNUnU6g+oHMPb68lF
EIHwY6jYQsAzsQk3d6SuxkjDt42WZTy2xdlyJ0MNhe4VnDfgXT7zIVGW7o3j
CEzaH5tsA116NSSkm3N8IPs8m0N3qbRd62QfGdp/GUXHJA/P0aT+pVcialCt
LMftoxT16gIAzLI+0gIr4RDiPwmIkwxz5VHCZ0eac6FjXxr7P/GvueBzNKv7
ba5cLPvlD0ECuuafOc0Du+PlBYPdogWpt/A/Uxkxeytf+Yh7qDmLxYULhdhD
0QMFchndWzyi9mUvNHxfkebUDDeBbMJbrHPChGK0DkqnRrCAzQx+I+JCBX4c
Wro8yJvn7kN+cx1gZxR2eTM7g9fJ/SK0/9siub0lg1/LbaAUFcmQMvPqrsas
Ffee+/tz2X483+LDCgiyNpSVDV+c4iXm23rECP92gRmQzWKxzmnaxDWCLfZT
jjY4EPqxN/UL+JjbVBCeb0DsojlFNFsK8BjFcIClntGypnXc/XljUUAd6i+E
JnHNryIN6VbRmdR+PY0sl631H+DsZ5q+AtHFZkUUKp/UdX0G80/DU1JhKT8L
yBuUkPmztUDg5Iq3DgcXA84i/10JXsS6EBYgmEZ52oevg7AJJEHIyPuS3yfL
UCuf2tSmmG6MAoMogU+2jZeFf2dAnTwXP13UcGVSwv5whKjSBW6gwuKvfxw2
Ue2RynL9nas4BA3Foh/816YlLsdjEvFNfL2vc7LkdIVYfpoo/X69p1Ji9Y4l
R8qxhtkDUIFFk0wzFwqzYIx2ubsvhx3fVotF98kDQLGJhNwUqvyUdG8xWSGZ
0QBu68iaQXBKelhNKu6fv2sC4RN5W7hNRpYrH5FA1xb23vSK2uJnyV67tDEw
EXFr28ePKdjWy17zUoIAPYhfI1HVYelsYbJq3LBAZ6mmgsD0P+1qoj6ixqHJ
O0UXxo5WHgMrZXsre/8tH6vuy10oP3yoV8F66Yeg8ROVa3WqZx1YNCG0wbnr
kzmKl04G1GDAvoGoZwmWXV4S4o1wXyeyYh01odZHrhP/K/wv/0gyKnx/OFLp
xOrWvmNxZgxvZ+tLo7hGSY1pzm6rJUfS+OPyWxI/Y65NZWQB7apHfpInQBVG
7cqkQPulMNPEqA2+KS+Dat2te45oKaoNYAtDUA3ADwxSSO7P/Qc/ElIIUlmq
clWqDCJLTsoVHAx/2/mSVXvEZ9uFYuPVvIWSBxATgYymq4aEgAaW3Y5ZdW5t
85p8On6L2RlXqyLPlDGqxPV+NwjDJiROo93GrD7jyyrGBMVV7DmyN0YyCkWc
8uqe/qCDWAH8/cxR13H5hb/uVRnE8T6lYuchog6ZWQ4cETWU/Hqpi5rJPTXf
VsmcT48PnrsNdpfeA/JNWc2ImOcqNcVSkJFPGpa3p4cRPU/QstYm/njSsxGC
5cT5MVw6APXGN0JWbpHKclVY/onzGW6XlVCAwTY5NpTXfrkidM+6SDnSydlv
60oT+/8xhUPBNIQKomWHlAixKxQqrQovlquGaRPY/NgBK/7UPYxJ506ekfhu
0HSdI3ynmdR3c7J9HNzl+2xVf6xwzTx69GJRa2UmG1awy1XfDTSoKTjNnzte
XDlCR/z8+8mCvkzA6WdYl03Hjiqao4L633fpdnPRpkiDaLkj5Z4Xh2Gw9+Iq
34TKSkCaeEe/T98c6UNZ8kUlyc5yVu4nL5hRql+F0B8p+HIa3qE1kFWdp1y8
6TOoc88bGCb8hkXu5Etn0+63RMfyJL1c214VjglCnyZ0SfrdhNXdBaAWQkrx
Pp78salrcc2X6wQc6ZQEwbUZ6gTMwuPXQSRREbZNXpEuYH+CQ3umo30E6yS7
BPmGnnYEGik7/Mm2TiwYsN/u5R4AlKYrAkMrCdqsqCksTY9FI0BNId2Pcb1+
+MLyTC6flne20Ni4y6Sj4hQhzTSqO60BiIWk3bAXwhd4XECJpWHXADKLINW0
b+JpJuXtjy2wnZga71Q9l6BSf2H5CsodLxnwOW4XaroeP/19cqBKCwrTBL0d
pdBukoLTAZIypZmvEwZgO2E4wV01kwQcNtrdrocpJCO7KbCLrasv1YwRfhFs
IM884+n4jqY1C5Ctsqh3Fkd8j64uSmXW60LYVrRuQHmfdipqMEt+wpNZN2q7
etX+AE6fUoqHp9ja8FmcB/O0fzf817YPnK0RM85778muj1RtOmKBj/ylpv/g
Fam6XjYL4lkV/Xz3T/4eXnWGsPtEl47UR9aqlZLTL6BnuSZnCi+MojbeHxCm
xO1gSKJ+sZCXxWTPGah/X6+1tJy+h8ozUZ8/ptWRlepXhKf5JFCFmAxJSabB
VNsAHRNzXyW2M4J315dxkVEGJ6OAG2ubtmdhd5rthKYT+EKuU8jApNUSOTUR
Cq9xCkaP98Vlu15RVc4xAvPtNhHcR0zdmsYrJPRuW+ZM840pOZiAhKkBJtZz
6siZUaEGQUrtu2l4Cd8s6BRZ5jKzauDWQHhRI0bLL8Srd0czzKZopTSvFe0d
n5/nYtcawB4WfUuHXIKCqYnqBv9Fy6v+g3j7IrI5r5PQ5paV8Os9bFkTwcxB
BWz2w4DsgudalnfqtbU219yQfc7Q2Gni2xkuRA6pF8ANIpyacyef4xd8BNBZ
2FpbB/4UGk+Blq7ris5itQuMpUzg8m/em4gPC7lcW2kgDwQ8tcZElmZGGkP5
KQlLBGbiEdKtgZBWK7yh7jHnM+ijCG2CrO0af5cD00dOiYDuSm74RTGu84Fy
/0bRC1+IupAGP+IPqIuTmzv3rmYPRUHqO59QnKhwXqhKJXxrC0b/hJL5n5FS
c5F5Qnv4GnMatK/c9CPJd8LiNzj6KNLb4t/gbAfPkEJ7KWeVfojMO9XdxlRi
p1CBs6g/IpdhJQweaoyBDt+veG4Wx+6VZ9chztvLPL24TMJusahsoSL2i2/+
JOXt1V4+95/cfruU5J3qxbgz7I2GSd7S0hUn8SzoJRxPDkcFS+5Tuhho9UIT
Yc6yKKWz2pL7NwnafawrozKDP9D0tPnI9jv7ZGCc3/4KGEbwaU1z0T02ppbw
d5AaqHrBb/Rks8nuLq0SpqdM97FGSBmWH0rL7kbzgc+AzHlQxDFNZbKqTmqM
Xe6NswRAtOl5Fm/7U3LInm7aVY1ubJLcQxoby+Eixgjo7XwBptTQpA4qI/BM
J1lWhdXMQPsEsZYLfrHl/U+3vklM9C4eZ0ZC+Qk3W19QVZch8IpVjH0EhhWZ
4yjJvn+lArLbZ/qSI3UDZ6vMiO6kb7GurrWcNg3mP9oZBo2jU2gzFJVkK2al
u/VY6FZ0j8Hq0C6ULRm19e4M8+j9J+8qYsGxp+h5YdBwJn0RnD+f4rmOO230
fzGMPp87HuKg3sDMFewshZdRv2Q/DsJl1GCBoaRleTfyTJADf13bUIADaVdS
3Q7caDkAwzj7GLLGdFW5WDgbF+6cZB3iazAkefhA2lbLjtrXzHQ7Bm6a5acm
UTwWkKPoE82Yeo92ONTY8Z6MkqMXsWcHR8cggcAsrvLwo5EZ/sxGh+R53U6j
9dqIq7A3stWrk0PFgwfc0gqFL3oFaCrmwAq8Agw94X64QKQrjclblWnDqNXs
gYLYlvW0moppWEn59JNajXZt9K0/5ajKCbwQ7cfe/3Q3CdlGPVTDeAOg+rsD
mRdZ60AYKaPkH/dRr/U5nJtaS2U6CStoevYMC1gspOgoDCoXJ5t1Gt+yVFeY
Wo7By0vfcYsv0Bm7scJK/uiNHa+EuUJoMWHfZeax8PQQPZ5lLaNGHxv519fU
wVmgE/mcSJGuLIYIYwrHMZUKE02oJJUU3IJBWDwhafQUynQZfVvOeSKbjb9i
8vmPxIypH5Oc8TKmNO8zEU9yP4C0N/UWA61KZbGr5FKjCKWyn+Z4vW7N5Dxd
URbtD/j8GkuDOPd7sHwsCXH8VPejf57GpjMT7iblLkJPQgQ8G0kwszCqZvfX
//AA+/AaZeu/IasrLUHP9bY0aahgJr2OOfwFKZ/gZ+8KkcpxBzX7HYKB9OHU
1T+UxzJ3lhTCItUneOY0hP33znBsemJmZWEEahm6hPdErAZ64FhMEIvcUuxq
YW8ZYe9u3B0eGRLCUCFBaEmJgtoLYClPinsjHWNUridCSQytAbrVLmIeWmac
aM6rtdNRBjauGJ0Uz7AQ3HnCxAdeCYMZtggJ15YcgnRXzBFeOo+1iBP8D9as
eYNSV4T/woNZv7pg2meRVm+9Odo00398559Vt334ELsT9G8TrjISxJHOGMMh
YzgiPcuQEmzU0JUdL/wYzpbr4fddL23TwhiMqstBL4J1ZWRvWh+CXOEbZ01Z
TgVAxKKn+oJs2PmjCny+AfJbRp0q6vnSsz+iTiOO1immMgTQmYA9zDUlrvjH
uD1E2VArWEFj/vpYAqrwQOIO6aouDRb3UfmeYk0BliTGpRwS139Df9vMgJdI
Xk9OX5xIOF661A0bQ9BAwwqzeEWfGl0uUYQexPwRtHdpB73MU7IYLEA3/Av6
aGMPOUrs1mCxByPpxIh2cG9SYEwVYrmAanGLlukiji+ntskc9gyX5eK4f/ox
5WjWSXL6g7zWbZBQT+7ncS2q9AW/blzfDad04gEM3y8HOAr28VDOvjcXvJdK
gRo4neo5h+FN3hKvey/e9GxdeiVU+PCamei60IL8FqgIcobxL8IieiSF+5xc
K4ubhZkzAYOWs6PBwm0v7ZDEICCAgwNYlEugt+PihmV/4PoFUgS9ibKlGsHF
EkX7TVSkEircDTSFiMvB3CODbUt3bcLk+ScKAhv/SS9rQjWwwv+bmnphypJv
REhbn/PemJOALnXjCsqJqPPHfBYNv5A7o6dESNH2aRQftlmrDc8muyFnojXF
+WDJ6cqyWSVk44BjAwB91MiDVi2SKC4VJAKdPVYRdqo90CiG8AZpbav/v21s
YVEFkqbxBFOMcrmUQxG7yRaDJad8h6foxbNdB2ogVh3OY50oVZCA0RkcBCvn
qxUUH6WRwem+36jlc5IVaHqUI7xgClvB81jIsC59murZwHgBHW6tr8GNkrpZ
BpSS7f74FFSclMFu43jRd3EfhE/Df490xz78ZvHWFO8n8YcxnYOtIrt5jFl2
JkyB3jBLaeeV4IgvMLIc9R1XpQho0h/Z3lW2jqmTooRtu0nx11vzSqGo+T2j
uOd65ocHUy5X3a7ZEU+7GnbUtKwvYyHYghhqeHXLKNXawrwotWSkTb4NnLfu
fov+PRetLmrlKfTAojnaZKwdsACtC7sOlnZxx20mbvcW23EUyV2jU81LXGwb
Om+AxIRKPE0LCcuV93d1Pqf6Hk7CNK8a3aNXO8nIP5a0+41Dpi+GcP/RAJa7
3opdj6QqKl8Ee7cRS2R50OJ0GWOF/IOzziIUuJW4awj5wx06GzkE0ur+bnGo
IW6Cc2EJyNj/MesHPqJG6ZW7DbjRkIg8X3SlAzsWRSIooHfG4k8tdrGXuRBp
fpne2LVhRsTdChOMbxD0lXjLAS+Cctx66u7rjAzbxDU1ahJnp/buzDwANPXM
Q449+pJ3h96yvkQ1jyo0szPmaS+pkS2xYqsHj4uLPUsYoI/hxJcgbanf+724
JiWLDDyEgcAdgaxdYrgZlCrDM+QH6qM5MfZw8NbaPvOuVu5qFO/4FfnG2y9q
e/r3W1kE7muSrneTIIRuof+F6g1uywLVLQ2zCUZfv7SrTsSawFCuppMXoTyB
PLva/C7izPIFV6LgoKIey8QIZTNlQJmZFdMOV0GOwDRLs1MlxSOx6ItQ/XKX
5PMyEURAYOQxzR3zBrOoQkt/Gm5677lsqDvU42t5O7yJ9XF91LInZw4nNZWX
kU2UqWU2Bc6CSgSxeG+poB8z5sx3mdlkXC++LJT8KqKttZSj5sb5op60GkNz
NfoHgwb2/MwQ0VGS/qSGll36IYUfMwCnxhOivHyTSnpSQnwKnFPiAWi9neY8
+/InyFEWt1qMVBqLMjBh05/WbZuMT6NoD6W08Ub61wosnfpqNkyx9FJGDKbe
gm4vgsNqWVUpbPTn+sNoDe0IEpOzYe5QeeJCiQSkXc7aNTtNGA4VJfprf6uU
DP/B5XIfqY0Z8i3kxqgssBN1UHZQ+FMqIxo91Bixggp50I88Gvk0gbVeOuEm
BEIPr+3BUo0BjM7ax+gldcudnyUydV2bI8h7S8t+cOp1pmtGG6lsxFcDdwEl
7K8Z9MvSjnJGXrD5VgmdXhPYZ+0FsDUCtmbZnH8+hng7j62nq8xr4IjPUBw4
AVwow6En4C67aQ/EN5rggkJgfx9LE40kZL7kBW1H3TDlwTJLuOlhcWlgJJaj
ErSh2leNx8b/GqbwDpuPg4lwgZUohU7vQBUadb5ULkSEysylvyaG4T7iDjYg
X/FNyWuegjd3AX76XGKO/br5GGSiIyasFyTjSQ3WgDenFE/umWOnT3h956dO
EE9Q6DdZI3enkwSfOo7INrFSlZqRWQf65WDCBgbBAs8v1aflLosjTlDK4Rdm
G7C0mhACa+yHHCTdMDbeO9RjjmScu7h7PJcEjJvrSpaJ90FYTUdGiFe+MNeC
LgObQ0oxUBw16lxm9xMbfCKxvUJwqasUvsJyXJD9G5KVOuvsCtpsMmLQxRAY
qtCSmvVnapxImXW7YvpV4UgpQy1gxhOFDE6PFhzBTjdtfxkJWr7p99XusseI
JmIicf5tJURc5NiPBNEQizJY0UH45EiBsSQeYYZWl/yhPob3Ilez/nzkDjxM
goqt6RTGPFl8rULpwiupSB5/9Okz5BoazXQb8fy32M/Mxy2UZxE+oEi0Kkph
poTsYNLdlm1rZymdUAWLr4hoC7pK3ZgogFQWjQedCGfwXdVpTH0NPJ/30Rih
FWgqNvYmNFj+vCx+/3LtNQMnwvRtkrBbkySstiLkUPzqzSqKDuQOrwu2NyEm
nIZr5ducnDU0Y5/o3GTrtpcrRRRSZszwrFzspr3aUeb/W95T5YXF5x0hpK8T
gXCRWlcTFTc3ll+mKRBPjsgLzHqLCc+48m4lc0EVwiKaytzHB+Ei9YIN4L4n
IRRyQiGRH7JJoXHZUh1VBWHjeatjeWR+DEMh1v/8k9gbnnMaf+ueO/gmpgUY
EiIuHZeB2hWy/wDT/1+R1S6wyuDAemgi2ZqK09HQBlz9e80fvxOR2dOrwJXG
UzcDVgTmyT72hmHzUQI0LBfTVO/KyX7Qmc1WNx4fKivjKUapAxljSk48ojZl
RIciYTEfClSl1f1v0lj2WMBoVGGNmR2rGCONp68xgnSEfm0wPf9ronS19yB4
DDXALB0Mx05OA1v1/Q1u4+IZli1mg0lkaFepYeW/pOdE8Mfk4P3Al3nMxWA2
J3vl7qr4E6r8PxwTIQs3/k9kHGhwG9jp6pLS1topeWneoN9Sw+em4B6SrdPC
TQA/GOuigztge2FHS/KuDQPVTe7UAq1YvlrbALkYyE6yda+78WwGg2g1sbHw
dtScVDkd/tATlUIscSj7ExJlxCWVY9qObqFF0D1rWq3oF6ZtU7qrVXyfEE/+
LAYhiBuzy/eV+xHjVfnkZTnNEUaBJHoQtNyg1qzTwfJKkHhdmRce16HJHmIs
wy3sCN8TwYVU/NJbYpAailUndm1IP2EznDpwEnlvYQUQX/K2qDRUgLsQ3MRq
CTOzRQVHouQEkzZWRcw6dTDzGNxn7q88f0p8wQYC/sSK6brB67obcaUdyq6j
HT3ZhBjc7zAo4CMUeygMwZIJhHTdkFjOhTdqX+Oppojns9egG1Hu6axrYOuY
KjHNQ507Fcpbpm3n+7VKpzMu85XMsjiFovMXygbIT+wQxDruIqBzBaBRLM1l
QN8lZwUsscvPxR06r9+q6kpoChW47wWmAARbxJMEvpXrfUpOwswjTPlN8SA7
x+82o/BOqZ8+Kr5Y984I7+VRw3sZt3BBTmdrw2fr+bloFoz2tdxCjnZFhDlQ
XxuCa9o+Alp5uIOgSbRaekoQBM1LZ+hp9kG3tOYdbShB6DYyRrT/V9qf5DR8
WQfuocgzJi7jCEe4O8GxlYFV/5dgJFCXuga93+S6NdZ4sMvwINgFSkfO4phh
k/JZQvbhwmAopwydjApaxBOMqbMAEMyGC4c+FKuIcTYILqnDaJghmLqYChsB
5P21g0LTUrmyI+3pPazyKUpCZh9wKdctnneZzZbpnwwfogRoz2vucbGDB/nb
jh9Icz/WP8olXxwPKj/nk5d1BvpdNgCw9xXR602lViYPFdg4wvuca8H76Jc8
nCTD7ZOqg6VdTEQMPy2sd4c6hByIGfAbzFPuAZJMQRDWIBeUupOygUhTgTly
/vVrb+BZ2UUhlMCzIRhF9YLfQTSsxtjza6LauI7HJL9vsVz0Nfq0vp0dMXy4
ANhuqcpjH1RxXpZi1tyPb9ROOdYBe6fzgiBGGS+BO0oKJQozgrdgnci/ZBmL
U57umHlsgeIusiVVD37oWTlNsW2KsYk2Z2IAg4GBQA+zf5I+vTosB3kwuBUO
Thn9xDXD8bUOA2q4LkhF3mRTIHKft/9LQrEV4GCc7ndialXZeksBkEEchxoK
wy7xSy5p9IrZMl4rZ0mci/T2Jzo0kGY1DcfpCml9L/02M45sHqVmOFjq0SHP
tje7mAVoYsY/xuF98GI5zYOia5dr0fuCAXLpiiE22/2JrM/5lxnihnCDzxle
FYLBScAm1qbULJjlw/DQhkA5hHiR+AiVrqNe9hhma3k+GqIJCmdF4r97kVKl
bbo/Vuoe6XtJaaBiYE2A0T4gVy2NVLjjBe9UuEvhj2wCkznD2o3Do+k3Ineh
fVxmbDSFdSWZmYQZEu2Cjpc360BtYkSLU3XKS7C9oyAuv/1iYjr5gGNDPAkK
lvvHpR+wPxu12p1VuZqYXnYA5y1Ul9hE7NhYjSMmaA50tjuDLiw7F+QbAfnK
pk2V90WghUktF73AgPIs+XYZmJtfvobqRzd+kgu6IU2sUTkV0XjnhXCGiKhL
3lsZYNJsLzm6/UY2A/1qb048TPnN5IA9MCjSRREwE5+d4RiMyfgXleBU15yI
L1BuoMyYTbgQuivHYc0jctn9xv2OI96sh7AS5WZnlZqya34Kj8kEPB2lzRuQ
6uGptN9uayZ/3bo3EzddOugXXEftKWBb9mnF/WCJhrdNc/AelxDNcKaAzMOL
J5teWr+4xFxBIsrXDSvEij/x2CplV2H7BampzT0r4RILGbSZ3A/x0XxEq+Go
cXs2t8e8LKwBUo/bJBvIR3sOGglPZ9b5k1i7q1GpslQGfACkdijA+DAtAIpG
L44ASNwfE1yj8KQU806X7HJ5y/ZOcPZPEF2lpUzr3iZUckyNsp1ND3QG2AFY
YUdonpRkcHnZ11k/Wqrsbv1+wCrFPm7Il0izXrLNLeKwT3yTlFe2W+8f7EM1
DSut8keJgnJLXSJxnnqRMz3G8aYrzGkAAFEUZB+JES1j7C6kDuQwWZX4qR8x
z7WnlkaD2sx/6P2sx962XFvmwr4n9RqvW1wRV7sOaRyZLKsBwsDuatyyBkgx
9TsJXCvIPAbxXH+/YMcQ3DxFke0lQzzFjxkxLxruQOger7n35mes/FSkHQ8k
ZxMf6r4oZxv9zWB66tO1rjEy1JUaYxo11II4cJ3wyaolMK7O7SirjqQ0P/+j
yo99Nw5zInXV897nGU+la3qnPI6dtmwwRA+EVLLlqXME7UkR5wouB2cdDIM0
HhNuKi8VHMncR4qI4eiZ8w5/b3hnjql583UIdyOAAs2wCbyPZBaHdN46brIq
PJATBeGpGD0ce1Il1jE8yDmjNYO0V+TnOYgs+trs9qU9m3VDqI+/inMilnDn
wusbjEm0uATJEolNFH0pes+Sz+K2FUHoDeU8US+5v2m7qlM3YLHqZywCq4kl
c6vu/Z+LSun+xAJ7jqDoQ1jZiJeWbWsuJCnZ77By3jBCNSpPvTOCH/DUY7pA
4prpIn0Lt9lpOVrnpt8sImWnTxlaxNKTZwwoqnUZ3tjQPmuNpVKEaUKcYWPp
vCAjsMrYy+a0TwyX8QYplVOX0HLDvVi/HLnEy0ZcomCHD0f6Nlfbb9Mip6ub
fBHWDayQYLwze7oQXXmMIudwbP978EsjKEtykxiL6H2k+Ue+hrBRFGiz+FeN
/FZYuUkxB4z22tPdzSmgdW124hbo7qbZ5soE2cAnbv30U4JvCLl1lZjvgulb
kZxs0yUlab32GDXm6QhF6OtPGUCLvLj0ZIxrrTi62S4+Q+lZ3DcFzQSG43l7
VHIp92W0p3Sm8HMtogq7+U+vQVmK4a9nU21XMVfTay59QL4z8BOY4lUFPtzM
9lTzHbUhO5uBxFBPPxTof5+kRgdTXWU8Sb5hWzYuc/uytYuyFSE+6uZwT8Z9
4RXs6nJJe5N15l49qHtYMRLDH72xKWDW3R7fRYAR3iu7nQAu4lRw6RIYFFty
Og0aVAy9d7vV0xnXVSpzKdAju2JxZPXkWiwJZES27nUczMDnPy2eLIqr4Bfp
wz5D7C+iVKDKcDzmfUlCztrS20aJBtvdIJOdmtK+/RS+Aw8PeKZor4iB6wMg
nPB1ZLZXLDQairWWhY3fI0yiZ2qnIUjvG6N+T/dzqqwb/51VfYU6SI7WmPTY
JKdbcJDdAiEHtUaZO68lB/8ix/vjqzcAeq5yHq8TTmBtfj02Rl2bN0/p6R4Z
MfHyxTUD4hggv+4mGJgGAkeH1j3NbuwqCq7+cKUtBTk4E7enRfN8Nu+h6qSX
QXxJM/8NXAGOatp+uTgHU7yJfNP7ofPJK85HnQpKQYLkoXF6lHfrp4yH1FaX
Z/7FD2nNekDEDqbLXAa34bMgkfhFpRb0lZBPNn3R5YMGGHNXbW9E+L608GRB
GTwS2FkgUgZgsq4PmFB5xnCM7bBUqQDZVn0aaj0FfD1mlgPtk4phKyX+fTsJ
kOKZU7djT+ieM8XjjXPCYG01p4gwgaDLg6D+hfGXtxbp0TuRwx6BaFXOJTLp
pTSyBRXCMvzhuq7RIm8/G53X9Hs2431IVLZLN4xMIsHaPGonNQU5JnB5BgKj
bcJJ48n2dSobCssIk28jVwVuKv6oYRocU7VGRuBBljgaEu43E9O+MqAoiRfh
dtdywmC6C0iTp2URhtPq4hm4SWXaVNvBRIE9CiT8W5t/ClkqzzfGy1FGY06I
J4Om8Ra/1MMT0YNzPuU0NP0wClUI/UDvmWR7UmuAh1pXSglXFHz+kuGv3aVq
DjaCzm3ord27V/tf6e/5/y6fNpU9u2qs43x3/B1R8RQzd9N5e5/wdGdypkbT
k1n5y5wm0i10u7uRFpLrX9dxzvwvvXiBiPYT4sTySz76pRPoTHMPBwXp/P9m
YEbiPtKT7oHhHRgMuZfrChac58ym7HHGEU6t6bc081L2BBNipJEvBaflHUWs
3qF6WHrJSoOOQzjMFxnt4SeKnrI3tkZ7yIruukM/OeK3nVcqUwrtYqVCxDJo
E3xENyH2ZJYCnxWoIMgyGFUnNQ8ERYYh7J2BOnStvLqXSsxn7aJCsDEqV7WA
NHMJntnHn/OlbiH5gSRhPEL5WN85Smri1WVPGtGvKD59voCkHVdwX5cezKA7
s0umqhEf3b/SPNcQYHudv3ixgHAEmqL1vDaCigq6+60he2qSzRznbLHRyNeZ
5e0ak1Fn547CR51FtRykkWTZeGT7ctq7w42tAaWhdkPG0lxqXPsk88FjxHD7
hq35LCNrZDI+fM9RuF+r6Zj+dKBDc5nb/EDJBcHZS8plsJ4g1N7NjD/B8y3B
rZBstBkoxML798DNjJly17ofazKTAMMZk2ujFrELdVPITjwcq3h3iKB6ZZYf
dW1AP26Zu+2p+8qRLKdjss/kjqmBNP6luGgvrhXujp+NWXDpugfOu8f1H/NY
1z23VoJnPB/QzDTMMhMRYTaFaysXes/uZqSEXp+Nqx5oKjw3q0P99UQgUSZq
nUlM6L8YVI1yA7zcYcqpHIHJAVf1jBzKcVbQL/CnpyauJeVhg59soebFC3rp
nF0uho/EJqBn41Ayj6iCVcE965ljlaKjyd0ofuf8mwU5w8czQ/A3S1ihgT4J
hONCyTG52N/LfB0MXxBOFCcuqcZCW+6MNnnpWuRvRMISZn3ZGbVo7GW3PeyZ
UR7PWuXbeNeIys2n4cLYuaHJuoMiLj3JECbnp4/sOppbGmaFfjzgvkBIREsI
YUVaDRpY7cMayVoAQvyK86gZAUumQ6i6PBU8f7HOFMi0E/7Jg409Rwup6Kmp
XUrIK+duNyYbdBZiCT2s1BxpB+nDCqJecyTRgO2UI0HwfeBWWkph14kNcQ/j
qaDkhZi5Vrh+ZraPXgfFTj4YP3IrHfePTg2RVVceouTanIitx+RDHHJ8RKYN
APHiLvDmuP951mQOrZul5555LGeS6xYMhbqPlQUTLqQ2Alkscl0zTSFDjat8
PdGL8XsxEWzoLPhTxcdCCE8dnS+tm8ellkkb25tuK+gf6s5wtPH+BOeehl5q
Qt4o6W6VbyHNSVLRyYQurS2tp1PM+VeS+jkOfv3NUQkDSF3rt9yLcTxGLj37
ko5C7mz6ONJV0tE6RhJrzp83NWESP1KO5SCS0NCiHKMQQs2TZSlp/CVLrVbo
QZP59hlUFBwlOUccCkFn69g3DzVnpMwvbv+jNwsbVDjGnP3p++0shCXaR5bF
XspUU+7NCt6O9em5OkTAq/B5ywQw2vpbcIn8jEFEibQEdOp9Sys2QbKhnW8o
OsquQoxDQuynJC1NsNceQiZBJWUCUvS/raCBsa5iG0Xmt8c2xJOBpZH8jEEB
uRepw4PlUxV1bMup1N2bMCJ0CZ3ysrRmRMrSwMg7x1NQdUS9zXQNJ4T5YrkU
I5CVwCVUFm8pWPhn1GERysRtwyY3zKspWnFDehufl7OQJtH8XUtW/AEWsJRb
TIxalbcMjRPwAhsi74+/Vk3vbOcSycNiv6MpzMyACEQu/UgEw4fOXnDEo+KI
VU3AcxfFfx/sgeWKr0RrGahhHqCbQwb+1Y/jTVvD9nKk8eEwJzJFLDmMVSyJ
ZeJG75s4ZmFPaafswQ4twfNlhYjAihknQlZXwETguM/TYx3iCUaWZ5o2OU2j
uNtToZz+qqT9gTH3RoSVYaFrjoE3KSfILBeBv63DjYzrH5m9SzJPy7QYtnjb
Db+3JcyBSoXduGCJ6R0GU3sZAN7QQORNF6H9RfmR8pwdzowJJcVSzDWr2y4E
VMItT2NSY4G/kuyEDDUTu+Px5+i4JSiRV8dyR/uuNDQ+4KipnEK8IilUuA3B
lvd1d51pGPpy1tXI5Ra/JeVaM4BOQhEkGK+yhiiq/LN980kFrDMTPdJ+ty2N
aQex1yTICSCaNP6QvIwkNe3Gc1yjvQs177zfQ6EhhljnfxpMt1+pPM1wR0S8
BWMHMoKmojPb4UlHg3SFfSFxq/pUawLU0l9dtHrcXvvDY01unPMgE8xm+J5M
puF4dpDsFeuU07Sw3fvqAnV+A1tIRNj3Svpqt9gDcVy6PcZHrVijGzAyAbn0
7OUnQARn0D5auFI5CwbIirSh/x+56Nhyz0Y7PRTYS1wcDQUau8evwgfi5avL
ZjL9T4DQXlhKHNlSRQOwCNG/TLq3GZA6NU6NqJqPCza2eB1tVD7/0qwN8lxj
yW1h09LCNnJ2o2EA4NIvr59b24g7cvLzZPNGIz8uqmXlf4lo2TIVV3FpyqA8
O+7y38R12Ot0PIPxWnlTUltkqBoFx34UQQgdTQD4DPBMfyX1E2HoxlR79UEl
3jpGJRWtZdxloGkrBl+idPou9wKzpRHuaOFsWziuRDKlif0/2P7cQlwrwVI2
jUyiprIn+i+xhYcMzHe/hT7o4imJxXQFUczazxC0plEm2+IJIfAl8+Q6aotb
Bxermc4nskvQdj6LT45DwWmVK+J8nXWy9Yhnyy+EzVnPYLy+XWciXglpF9ev
SI80OH1dy112ctFkd5CaJ1v/1P+MloxUH6uKcyQchDA80/59YdifSATZUixJ
Z0uQIZ97QMKgquzwnzwxeEAUSzbs9I4mVixdHyEQ4xfDEt+Hjl5+5TCBLLa0
m9GLbqwXvwksfTIZn4WQMcOTmGPY6DYLj2xpyBKMPyDxF99MC5WXH14wwCyY
Vwg50C3yWqhyMv0iL4fN8Pn9IBNJsX8KLRdN3qojCbR4y2OaxDi+qXvdxiVO
WMje3WIu2LMC7/pugg6rHI1GGmYxgMc1b0zCabNO6fSLCrHMP/XrnwtyTfg/
Q6DuYBt+Rjf5MRimBxoGoylm+YREHcF15xZNkYqTl4TBve1HFJi1hhOXsyxP
1VdZlK6QCBMkx//sta7ORn74zyP+SU2rnospR4YQQW5NUMgOlylHEe+2QytY
r1HC7BKmBorj6hdT+y+clgSWvdNDw0J+28yeAzmwRC47KOZRdrybGbAUy0Zy
gWyVjaHT3BMdcy0H8wdiCFWIkeFlbKU/Cl0LfjKa5wSo3maN6XXid3FWRLWQ
Vgb2xC2RoXibOiM11vOMK7znvVzqaMt+xQirEsRnDA8n/xxKHLXJtVG+/FJ4
jxhsgLF60CooFzArXtHgYWx8ZRt0rHUexZHyHbTl+coY54C5za2/zJLffUEd
BuZBupv6Avv0Mzzgba7RyFy4fe5XLBAM1J59ow3CRI4yVSw9WQaYTEzd7pNs
ZIDmvg3LAzZV8oVtJZFF3YZOxM9QVcCfP0OIxRnh9JvZl9guKpSfYI4ozCQ+
fEM6mK2Wt/QWsD1wxjN7AwGMVkUn4mBepzfN4mdg1sFv24DQxziLRKrM2Itj
u1UD+c4kge1GTVpSS4YJhM091YxOtvhJi+y6XjBfcB/9iYgrsa8+ZC5bKfys
RHHofdss3p+3Liekm2zQs163nlsvrR3CpDpmR9gN3vDzjCg65Gr/NZWuO8pd
k8HRKWwL/bGPSFfJeew5lg34QTN81TtbNNtw4uBVnS5mrYYpd60nvwL7tMzV
xSW7eRUevQx/hHxIL2wl5qpHsHYNB3MFNqAHAkbwhl/PxD1afuh3QUeMRg5V
tXqP9kQ9DLUSmjypjiwptttrWadYR5gkJEr8WQhQf+p8UXEBtT4qBLGO7lIc
kp4yhVyr1qS/Biq1tUG371Xl6UFg/QNhQdqmiVLQyuIg4tN+9U9YcBXDAY6J
iZgvFWfpmh2X3wWZIgJe7j6akSwz83cjMf/3Ke54qso5NBYsKIhWGvJgQiRx
0TAct8w3T4SrXbpYJsv5F17EGszp4ixG52IhLCghupaTE5idkBsWTY3aGYoO
WBiCz6bI5w4dS/KjyUn7Tz/k8xpQMqNJ6BKS1e7UQWdm2Eg684VJpto+FHdJ
8UaawnIiurQRp/+SbrQaHbxUd6ifQGXPUgeVpz0cEqSnqii0VhMK7/zSRJDU
lqwO3wh5ifNG0NM8M5IigqT+DII1CMjuVb8QbZPeyvWSJ4Tduvpc6LVnNjRi
bMpsFIkRXQH9MJnP2w7KeSWy2cMynSwnuFBgVkzcCeF545hHA0bYNDqyhYXS
gU4ZOg/NCAbamQmF5SaH2r2g34Lz4DltZ/q7Jrh+nmUts7vj3EzJm/g7DJmZ
fZlUxyM+e5lLPb6j7VgfA++9NlJ4t8U4wLqTXHo6uVlMAsY2GO3hwBk95QyZ
J3/9P7ZD3o5HbFL2TLQdxELZn/Ui94FU7nFW9sjIyOtLIrD30h0STM7aSANK
3+nnrf+N7YrE7ouWIz+VLAnCF9yblA3D90R0Ai0ZNQeJLMkW2g1GxzQiQ0HN
qZd0iHAaTbxcckaetx+0V043j/r3QmEb/Ph3fnmKBvdhbBdLdhj7wszrTNJT
9qlRUw+oy+dNldNXwon1sDB4scyXr+eKfhBN4WFYw8KJTPJi4bDbcgOw4sof
Eth7omGXz3exd9kMeUM3+q+3l4Hf7ihyskecP3C7uTGfHN8xj8FXAsc1Mcpf
4AfEdacgaihxlJs1sDn4S1pyIlo1hlIkIVWbzNix0eQuUw7l33fhGOAQVyC9
lgQfFXz5br5D/q/RcR1F5tfd3L8o4CEzEyKXjhQIO3H0erTush3Tf44wU9xH
SeFMICyC5yxsMsbpaF55yhNkb9fGxJLr2MwvKPXMaK8s+B6fBLzKPD2DMFZ/
rqxx09ZiYXanokUyzHaF8Woq7/32ubhDFtP3StmKsBvjUPQBheDhNuEKe8kO
bfHw7JQ1qlzlnHn+XrQ1cHNtFDqjXzSf7HUVJKQY5KrSctIhsq1yf6qgJN2b
icwTtfaCeX4L6DSut7EeSm2WrsTAg6T7wWGy4+0KA+NZyU/JwQ8ApV9N349T
hcyRoElzeMb9VbruvQZ1qMy/9WJveV2z8wyvxq0+J2ergFTBws9eB+eSLBTa
4uDIP9oWxPEoVtGm+qwLso0V6tp4OF1TUoBwF5EvY39XjKfmscupJwFuJmX6
gArNhBVeJLqQ1yhIUhthfnsCXdBOgw2SBNI6Gtt5wjIr9rgo+b2M/LnlqlA2
X1/ZtF+ODV+0yjVs06cRc9JuFtMGY6hfHXXcuOvkGJIKykgJWzbDaXaeoUZK
v93Rnss2NJs74d1NKv2PXhc9xootx+TYqwHhUdoc37gTtDTkDILOYhS+P22n
TgirL35dx2IlgBNDhS+WuiEAcTuqCh44r32DWzLOvZ+w+2Wv4g3k1dJU5sws
yIcl1a/2qJaGr1yNxxiwiAHpazmtwKP9FjlPuls2uRwtKzyC5kufHx6QnGFr
cRSQEaGKGA85beJ4LWKAparnDt9H3rb8WdPc8vZwxLlC7O1oPVa43/RgCmsr
gOXL4z5ylO6VdhXa2WmcPr38o6l165TfC04+M9pU/LREC5W0JnCHPehSRKY5
7haKGw3ApcIbGHpDDer0AooxeII0L4eGnDmoJTlmxJ6QTfyaRJeMZvd3oTdZ
CVinaCtPWJ/Kx6wJ4puVxn+CvJ+3hPjeSkrTRMBo4MAzFh/qmuSWpQiNDZaK
20OweVcbaYzTWmH5DCEVzS26dA6X5MoEABQVxCu/4RX/VOb68C1AsN5vU3e9
YyeQlrvACWn95fCaaxFdU01CS3UMLvKXwuEClhN84JUc0vWBE8OWVhVzRezu
hK37FLXNYaEXLyjtYGA5Z6uR6KAM/nJsYbhnU6gA5Rm94PEbEFkYhsTOy7nz
VRozAX0C68PTkPtKAei3Et4EPTBtaoA6NxFPP3idEHPzAif+SVFnpiXhIu3X
FrFnKHm0VM3wOgG8Ku/2gJtrg2jQnBVb0sWEn+uGn4rT0Zx67JaD7BJmDRuU
YnRKMp1C8KX3k0OKpfqpe3VimNKFCfPJdT4tGapAn9SzsCv9uxAtwxa+Z8tX
/5ftT9EUNYSpxrxgxKo53I3KHHeW7a45nq0JbIeS6u9bDLc4XA5Zz7h7ucbX
RlyyA7+cgUs13N1Zus3h/2uImsoZBvWVARDjMog99VLBwDtCYRpm1EYdE77n
QItx6EExtiU9+nD5TKxorElorNRkFkFnWxvQ8gcyFuWotSo/4lphxuaMNu0/
J4S/IJe8yGvxydKbZ7t6ztTmfxG2VbS76ZXsEQcJXqHj/Ia7mkcK/nVvxK46
p0+m4xAsff28AeFSQbS5Pk4abJcJM7r9eEBKGTBX961bOpjrSvNerTwh+959
5yv84ffEiveMNLejLLoyg6WbJCmGUd7gs15CRRQuJAYKdjn6Zxu068TqiniL
aidHBvMjBoavdUsIqJz1hmk2DK00OEifRmE2RtU22m/Jphj1otTYkFt/rkKf
8c8SGrxDHTe9pRTpabxbOiEdDWv4gQ+nyL8UKULzUPDf5qlQGF9+4hVgL47b
l6sYAn37GFWllv8qrWESuxbxPZUlHAjy7tAMd1swKc9q+2i/YTxmbd/3h8uY
1XsYnTjiYw03MffZ37ynOIfvPV2BlgeSXiW60rdWITfxbPOYaZCyMXJiWqbR
lerHlnhkGfRiDvn+ektHFCh0omBnIv/OffjbTZT5bWrTWFw5BsVo+pe63uSx
JFU8SEbjWaPSeFQHlHEDpq2iCPDZqF/bUWNfwlwgES04Ub+4rnWdbsMQvDoA
radWzGrgWegQGtaejvjl0WeN89N/+tG2AuSyc/MLGXbYRI0dtcM8To7S782B
ZRC1JCHtzdepmgQnd0cgVDpkmyfs8MXnLtHI5uCv/0keCYISAP3sGq61nOwm
1V2/npQYXhyqfQIUpq7Ys4aTL9PeCY0kQ8g9qKZvMBW1Hqf1BvZkF78jD4fb
gKA23Y9EjYEf2XKAj68jSQJS9Sf2/OHhm7nzKgM7hw2WdimiIlmZKyKh8dmJ
JJg07dUjRQQy2wwWxxUVb+muMhiYn8gY2djzvjXL2ICZ36FNUN38ZtcpQbZn
kJm70uec12GUoU7At9oEBojnliTOUcbhCo9p9yEGjj1aiO9ATUV0anNIr1zJ
+egcpgKPCa7ROWe5l6/Lgd9KzGwon140WlodGlmY6EL4x32/jUxWPVw+Ux/S
g3YUSit8EG7m9WxSX7A7fKL78j0V/FFu9hKgkV7YEGnSV/pErXy3f1V4hhRp
FzJnA9Mry8GnFgCAT969Q8GkgSWpavbcB47SYe0uTWtd+AZh6lSSc+BkNt4M
bUPIdc6tJazHQxEY5yVfHO3+QMtiMI062JkucqIMUGTEKvn9CiEfmt5Lw8t5
duf2uAs0Sizl9a0MjXqAJE4DvLVBF7F4hFaz2ROo832qKheyeYuyj4Vb1vrK
0HlfXjO/3aNpTkQdBVQe4NGeGUO6BqLmd6tr8oCZa4SedP4ovzMaVg7RdnBf
i8yihEn3bjomSZgO6VlOr83nCU/zmQJNCY5JsrMvrTsQQ6F+P5k/CorLFknb
UzfW3D/4DZGCMnZ3vMf7BePcBu027cMimlPpPg5UxyoxdXZodoM6r7qWLKTg
3vkULJ6S5/CusT/ggLgyAbq274ynulmPXaWsJoCIpmdA6d8+mLm58XCRBXRa
UUZCM41wuuHDFDaGivxto+qr/IwrmLO6XYvG75paNduc472zC1guGo1xl+sm
/t1OhaJfLr/shrcxg41lq9fXXu9zK2iLXTKtTYADcl/AskoabhSclMhnYCS5
F39TIEwd7Qmwq0Y3Br9EA4ytzNaFEvIsvswtySDmnYN6GFUvvNMyVLIL+q4x
3+4dOqYMtKYBunQqX1nEYbEFGbXhup3G7oI1HNJoUI0xVLG5MBw3NO1WOHp7
jHe7fDMJ8A6onSQEmpUj/23CZAW7oYLVCVis56jj+j4lXZ5u8ToejtIg19oW
4crxDBfMowY1zKdvqfMAkkEsDUtob6jj68o+MowwIQUU0RKAn5uHq5p8JNOz
kZCp6UJo/KrH5RMosckxO7PskTcs2HAnONhFhC7ZIG2dJ5JPxyn4c6ddW8/g
n0L83TP3V2etdbF1vSLcv17SfveEjrS90zBCRBosYw8R/RL7D9FBZHb2lOcM
SF/sy7367xpc7Gxg9m5LwmO3AVHfvIzNC6hVLw1RCD78L2dm/cNahB8dxPvD
Ve2RlOtZ9Pp0NKpdwv3eRHDUB7+2iP7qE3uNdzhx25iDJ2tHA7ZBNWWwbIVX
RCHZ+I0+wlL2gNBgHwywz/wkPBiJSpY2hDYC3lnrH0hPdnpQNKCHVOQEUlcy
TTQy+eFML9EOTbXfy458eAkpA2HQ0jKsoqdxcuXcoDyAL7vembrKM2haxNMQ
/jIJZ4w6xx2DlrJkhWZ352N9NSZ83LImsPvmGGFhHmkJ+ZroJxz9IR2IxKSB
XSDaHHmbHZvOEe5iMmf4mAJXrhOBMC+LPLjqGiWIlxDX4uoleRMru5Th6D6b
+3lEFMcfIaiULiyuh4d+k1ERbRkE9Q4QSdYk9WcqOcgZEBd4r7VNtzFPbZs+
JEXcHe2WrS4JQQg2OZ6r8c3lPucPVXgppm47ruZ6HP9GJnucOBCmfCfOnkJR
YfwmUhybkHwNvqijcbcn5RPWc/ofUGEuA267RakdTNrFoZZ4ku2DeTWzqVvq
Hf6Pt0ge/3vKFuvlkGvX95+xPN5aY19CbSGzDn2xiro0sKWVDCSFELgXw5Fi
L8noq+CxBCrMtf6xRveivzwJHfsHRBN42gu+i5qrNI/15Lis1HIICoShcX3e
4TYZcvmOJSzLMeth6muiE9XLWuc1uO5XuSAsQbRHgg/kWwyRi91P/W1X0uFd
6Lr83iruvWyvzzOGANoQJEe31JxopKj9i78D23SJy5KKi4mbAHFM2GkM9M9d
rfyZO889z0VkvPEbFHeAh+eEeGqZdh87ZdTevZMafrO5SJFMP4eb9xiqeOi+
dhRJu0nwvPLVNBVeD/T7hqNDB0M6WbiLpsrEn8kfJPRV6S0uKEgT4W3wkomu
zwaLNEGcrCt7qQEuNKDEwXDMFpoCh0j7itwpKNgUNCQieOd3M7DlXPfetBFm
i5VL5F87v+guwyuz83Ynjasyuf2vC5mt8E2hOyYCA64Ct0aBhYpz6niYNsNk
AYHPB6yZKSdHvauUuBBpigoO1ekCK53u7z6Xb0MhOSBUM6QtSSKtJjtt/eeU
Og4+mLf+/J2Zm5RRjCiVR2GXQkHRWVAfiOBqlgbMOmVpX3xhxpaMJmHpd+E7
7LdamtrZdZanBryLCTyRw9fkaxGHeDtlnkTUJRam/BOO/sHTeAGOZCiIyJPg
kv6aNyEx1blHgSz92IRf8bRrcopKiW8iSnErUJRLbUxKhWaAeUoEjdTNnMiU
ixfgUhgmHDfvVlmBqY+UKVYZ5nbRVVoa21aRJuc79Z8p4n5UfMMieY3RmFzh
XXAdqGvZu2BNBMh6nfOyO0xrPRX7eF7rps6bP1ZPP7wW/2pb/eEQtUUe1YYw
LnP7l2LCTbKqzXcYRh9yV2ce5wseO5OyKHqRlQxYo6ryube6RXnCb/YRpxpt
hJ0Rq1pYdHvMzc1ObkYPj0I9Mb95S45zmglOBfUJjyfLxmni7OmHtChYh/Gn
HhyVUye8dPWzZ8p59llq1RM3QTbfihpZDnfLIluSXWtF6R1T3FSWKQBX3FBy
u4YBg6J5E6s5XBMcUObyuTbb3DvYyT8szPu0rmaYQndiiRHGVFOk8eSx0mUQ
uanwDQbZh817m1TReWolyhGumbhvFom6N5imCopkWYmRBvoDrWskloLhRnZY
YYz+isFbIdhwTDFBFH1KBNMzSs7+tYSumgSKCiU2PFGlQQ0ljPBntFM3wsOy
IRvkLPQOng7UW6eEcysc3gQf/HPQ41VMWC9h2qThDEAaupCTiP2fRz3tGOz7
aLwMH6ur7TbUCmSUZv7y93+HRvuQF1mbUtudGXBeY0/uv10tHO81gTNPci1f
fGT6cUomyF2v2EM+UwchYFiy8aGmvJFc2cBYgFEpDA9nKylv6jCEA82ITPFW
IT8uOFFLtniO8IkeDeig7ZrzMpRR42TQ/HSU6JOpK5DAEmbzBZeLcLDJ3F+i
2Ku6yy1bkYLMFjXHSnbJX6pD1gKZLj0ZG8D0B9wTDQR5Osy8aN0NpXxYC+2Q
8vw6L8cN88UCmoXXU4W5WdjWCjDWd44+Sg8cFoNPw7tlfarZuokGVfP3FgCr
5Ir5jEz94Cuq46FH/+SvcXCe4j0NOaDSqXKvtb/t4C7l6Loggp8qvEYiq4n+
Gtye7N2laiik3SwnZ71JztkskOGzYCZz8yTnLi4+XwfDsw+kCEaiaaCIjDHt
SRUlIA402FolR9IJ4Z8l04tEoj9ra1w2VImJaiYnE7kAahSY/pAOXyMZzn7p
kZDC443vOBxX/KckRfFf3pTEgp32vDpfK+o+AqaeccyJaPKFT8pFh1LurT1g
N45nJbziefGD97Tpb8CsCG/bZ0b2FapuAoba/33e+Rgk4L+Dyxf7pWNLZ4PC
3EpD9QMssFR1rUUZSBAWbILsk1baa6A+o1uwMlpWUK+0u3MOF2rC3/vUEX0V
i4ld+kqgjhe85hpBoW0EHydo32uwL7xexhHa2lCnkJKsNO3/aWc6vcGFhhKl
lHzNgWYrEwNqFOV0gy0Sr7LOtHzuWRPMc2JJeprS8aZpAQlrrc8CY9CP1W40
yWLXsxHazjK2OiP4wUa0eSz3GjU90sz3tYad4AKBYbQk6yFPP+M3fx+ylju5
g9uNZBgCtgzKWejHRMxC4JZF8cj30Xlz3SoE2hy5Kvvmx6OATrvkpzrQL39s
AJJMg7d3EqiGdlYDg1eTbEeTlvk3rWTI8a22P/vyN5WqBhwXAuPfZe1FWALE
IRRddPJop/6zXP3mXWOsaqoLQV0FVCHCLcq9nb8ZPEBJPnm+RZVqijB4zeHL
FcT8DXBFZ2tPRw+pu7jHmNQePYAl9qS8agSgw6I+heb6V63oCEcYY81v3eNY
2XM/+KhCysQyu93fRu6BjNUTU2+4Gj/hZ2JvmsHC9DBo+88dwK5qGlQpCqm6
zqZAzpaPOcTCsGNM0t41yWay8suxj1cW6WFMsa0YiHE4vP1hZUb35lTSVxzP
ZC6tt3M/LvWiQ5HOLg4BBgIhEvm8ZkDueTYBFNLbFIod/i5pE/MsxYc7Rs3y
1VfGcMahRpwATIaDl8p2JJyhxJfHwfcE1C47ioEJ7eBQsBNTGTRsEt+H0PTt
fnfegYmp4rvYqYDPeHtr6GSn7u3Z7RqyZrz4WJ0xB9HsioIf+3SmRavqFlaJ
4Mtjz/KYfEvCTHAE1Dup3jjitklwWomwyeofs91J1wOEnVxEjMYcom1DudZG
QXbsKcya/qXIHKEi6PxsqLue4keMY2AzMpdQUbS2DHGrjcXSUbG0WYB/pdv8
2CbMIDn126cugqCdDzN+3ZburLK5wxtZUrQ6o6fhMEWa7IAptX2tt9QNsfK5
C33w5bkhpOr64C31eqQE01JLk9sn6UbMnFQ5PLjAJSqH9jelZQUzdq8wY3tQ
6cqvADab90HcVuHlS0b0GHVuVgAJ1APRK2nff047H0r343mH1C/jjA1M0fFP
jxuO9ZC+hDLC6dHD/BZX46n66v19gJCfGso2ZAKKbxLH/onDxrCLXwjByfkF
EXTFFp8JhDZQdLAAYP3k2lTzhs/vWzAp6cQGry9kzWdbWFctrhFKQzSqRpEu
Ms9HM1lIUdAdI5f+bDxsBfu0QQRYDj8YthoU/KsgXuqvM425x6lQ8Y6f5ea/
qhe8W5xIVDCos53b+iZMWorm8RDgV2ROnokrOqRIwWM//zRf7myqFckCUUpB
evMdOQMdNh4TzZo/7RFnoxE+qiGVxpZ6BnQATkQICuCN0vwI9aIVJg9DrQ6+
wX5tgrWeigRLaCTDAwTihaQ5RO705xR18d+U57COoJHKVREPdLbcfxD/MpRO
7AeqRJfjZjf6UAr/toJc24Avmlxm10Yqjr1KXLgPoS7qHpA/xRCWnxNXWnRZ
QNuge2j029KwXr72WnjXMBut9kqmydl6kfwvvH01f4u0eILIdBG9KMAfJpJz
pbzLZJFjq4gnQvF3K+1nnhk/P1byIQ7GLz2utC5ADzG4p9K3NREhLPy3Ut7K
8jELHQ8B25HkhAiPMWGaNOHGp+xJlRIKtQdxxfTr0rclVa6cuE4mkJ9eUc2l
r6vn92ZYloDcsR2/6VnHy6+UcvS+l47itxrlUEsSs8zpRNQyGQvuXGizJVbU
6CO9tbyJQoQuWfj46Ks4+cnKnt1TxZUDGss95EbwUwBpeu2UUOKCqfZwGFrC
QH53CQ1nxmcc/zXgkdRSU17wskEW6mUp27AorfiqhYf9TPdLN7n4ns2zZrqy
+HI3vMD0q6Lf8bSWq1kIuOeFdrOeuni/xJiT0Iabuw9sOBx4JeA8+GFSjclG
xDkkuQCtIR/NFMenponwlFhXus6inRpzETBcaOQ6X0pGqdMT7qrgiGk+Raod
BK+VjPuM8AKu21nUYOwhENzJsVD0R7dZLNcl4HT6Oh0MaE3xUDjPJUEBD7CT
gzYuEB9PfCrcFo+MPJxgdzhDRRRgc+wEMlZVZ4SEOcXL0Aqm1ltqAuInA6e9
KCElX1w2tsRpwB9XIt7hbG70yu8p3GH0CdU1aw67uGsXw9v8GLIbVlhXyWJM
5u2fwQGYwNfEZB8G5BBZtR7P+fFStAay8kQNcnPYegQqA8X53EkyKmK99Ez8
GZh6xhDTQwhQDVhkTxbzDAUnlwgPh13F9szCWR57Fwo1XnxBobmps9ZSMV3l
d4VQ1ZFjlsw0XtDFXDXoQzxLGHWYwb8idl43cHGL1xNwTv4VmM1mUJ8PlH2Q
0bqcrNBrmtLe/VAk1+/lLQ83OvGYkrKsb6YNzWSpfa7+jRg6P+0OT8YnsmRp
srbWGrG39UHickhLEkW/IGvkmWxC8ss3IChzNyRDHmZubvHxcDuiUoiernuY
K7UwDuIBY8YhuRxc7eYBxnXi1I1gNdNYnrO+n6JlBTfCA/8ZJuESE/jeSo57
JtZAL1Joq7ryeF85hBCoKzqfQMxPbdMDiqyDMe/iQKzdt/SAHuU6q/5YkqSW
n/LBd/0rhI8H3H04fSeBzInNy/vFJi9640eQ/HKL+OGAA2yGnSpP45nI2zFd
CoeuVNpMxgiscK8nloeVrKs2k/rNiMZ3+xmxcNbZziVJZgeUaz6297Q2ArAG
W5Ewh1SMWkkC+2ejB91mI1eqaR+UiejjCulmJX2GTfNIuIEnkEy7yRK0ZKH/
eFV9qSMyZjgCGdqX+ESsgRG+NnC22gATi+9Ruag10AqnO3LKXfk0yjhbKPsx
n3UFE2BQM8vQs0hyAmKFNYSVMBj5u2Dx7dm42sq3y6v0B60sSA7U3SAQa5Ns
ZSczRHIG/6+Dg+R7dDE/lhBOO4cenlySS/60pTC5IAE1K4X+FemalSo2fxuO
cK4z39HSa8UGdjxP9l5dHC47cF2KSrTkpT/KsRQRJENGO+8bGh3bSdK2GVx6
vybxNkUtQzOYOlBBAdep8vIBzbY/J+Nv20aysU1Hn14P/ZHQwzoYDki0rR42
TlHZDBW1bD4yOpP8wuSbALtYQYYNYHUPp+s2QUXEfa2oFC1+zO4QyeZD9ico
UUAQ3GfAsPrDrPAB6TeJZkWiJ63QnZlbqNuTZgPdUxPydPjcYUAOjnUsLHL3
aez6ZNKTuuyuhWfIxFji1VT57vSd6IqZTaQf/IQesosD3VkypAcz6zwoF5pC
CdNofSWEUvzwYVGjP7mr13PF4fuyUKSN1TFCMRQ1Wa+JXJAIwhcGCNfR+ROq
i0ErfjsOG8CJ+rtEAvjmm8kSknrTMtSW3XrZY/uonZOkg0dUG4Axo9KgU9bg
oJus6uyoLQMTP0+7B3JktFzAQ7Wu5ut1tpLMX5nhBXlW6BCxgOjLvv+m8y1N
v5jGexDMmyy8jnXojoZSAOCnccdDjwtAav4uMiD6b1KNAu2Xhvdyo9rbweng
AJjaSV8u3bOOtxBbYCKla8/RY/afYUyf+Dof6SvY2ev92tMD0rQWW0VoOMQ6
7kqULPGsHIdCBVBjqKBaiISLmJWBW9gbt7j+lfv5GbM1EvhCuw+2CBywc9x7
jk30a9azCUj9NnJtNiGVomF14BpIdvFJ+Lk3A50nebX2f8g+KlAljMiqmdx0
xfEFuKnIo3wzC64UG/djS/MvZNBFhQZYJ+T8+fx2HxJc69JWU2WTiiYcdRBN
WPsVHsEtf5tO76SpHZ4Sy45u1dhKTo+wAuosVMEEuWpnnJzGIUCWdLGFf0H3
s3WxmpQpVPVeCRi4tnBEpiLa0J2Yiv9YpMwBocj5y+Hx3JMD3nqQO2/pWldC
8/axLcRodH2ySN3diAbJLkov3mXI24azbfVgxgtkF8yS3ZnjHUjuQ3K0u1it
D8WW8iKAtjkH5FdFtbuLGMQZextp+2RiGkAkFLsplXxVY3tFx12zGOEBDBzt
r9jrTj0l/sGQ/aVSPIG2ACR9bFhlYhOg1lBTkkPcgsaz68GRcWxYQpKrwxNY
ZwBBhjYpAAxbVMfc3E0haWoUdIKF5kWdG5ZyNGIn6RtbWzHd5O1fL3A74bNb
s0fcCFfVr+uhk0IBLU5Ixr49FbGeN3YiAeqsZiHH5XhIA5JRoPJbqLtzGBSo
BTRkXfOuEZvkdZTZg1a/5kO5i2yjHjqdSAiZMtTqYS7fzDl63soI8aahcMAp
Ysrz24z//872au7wjFoqTiJyxkRO6QnNoJHzfBGcYeQDA0qNMyQU2oJl5J6t
23zgwtcv3xLChCl1F2AMMQ+ijdb/kf1qTt5WOLQxnY4+HgbHAPkdVKIucuNh
IhsxqOTzFL7NvM8Xedgj1sGv+QGY7D0KOK1zXk57f6TU9Fe+ZFuwDuHH1x5a
ZP0J2v+uYWy1xL93KI8Ovfw9wTyjYXVaFZDKJ628+lnOSZWFVwpRJR7vXlaP
fMPw6+LeWSuopB12wG0128jM/TaXVsNvzRkDkUAYuge8h3NfrX9JFAYo3Dga
rKqOY9o0BFhABuhnC1ET4W7eb4JvuR6lsAPGqo8jTlrnXju9Z729bjvj+8UM
OjhZa+LflWCoq+2SQkEpVyQdUQdAbdDmEkvsFkkDAa7G1hvw51LFmJlV5+e4
MVyvZ44CNFaKnNTgbsgk91xAMDede7RYX2fpYjjNPobO3f3ErMMyCg14gkLf
tlRa5qcVvSD6ksEDVR+jDLPFXLeIoBgNJEm7dDCLXnqJ6O/IuLsOpZj1kI4t
OJhucexhrrxWYRnEnqodwqHkZ2U7IFjDMTDd43nMGKxae6pBInl6u36qRs2T
bFImm4XwTOM2yPBW+x2JTrL44dqK8XbEk1mQdOdvtN+rUETRBKnE6tgsrphV
8xLRgF1TX+LITgADPmOoSRuDYkYcc1tKvLV2q/RxH5ZnU+Ys+45VqTsE97fN
CVskbDQfW6u19ecVW7O4M+/YZ7ehT5fwSDxN1N7Ve5X4XMlt9muiKTlxwnUa
MJDKcP8AH3/7sfEAnjBPv/kOamv5NXH0rW7NeV2SfQhn1ytzZoeoOTKGzL5U
6tGZ+7mszXX1PpbOi8Lw1x+2Mcs6W61RnC1HxLmOL9aVh9glG1YpjgEii/Z3
kSmGJbVA+guO50TT7WM3VgZcz6E8fwtG7Y0d4jOPHrItHYhJn2B+kJ2m0FD5
ArvNkHGfDJK1FMf3TNDMefnE99Bw/7jSUSxAx2o3/4hic2fTxCd6RHnR6Ag0
ZHVn202YELtNnUl8xblTe9oONlQOuf4IG2soiuFEocB/6WkSx+Edwb6eXeIn
18Ydayl4g5H2jA1sC5G2ByoAg5OIbzV/xM4WJd82tJibBCnaujb642lzrikU
lTfzXhOkXcLq99dUDelLLwlpMsP4cXrFHYhU/v9qzqY0HV/A+fig0gjVhaY5
6O5Ab3+Epk8ZAipyCDf/XxFX41bz06GoZuBIR6/qasZmaH/JeTv+xVWUmZnM
UzJ3qd4pWyG8LKNoJHh/eP1M1IgnS2i8uk50TC0O/mbP8QibZeFH/6C8MoUr
DJWUgdf1PY9MtorNl7M6VQcsciFs42xoQ2YtnUudGRGawjeIDNxzSvCW1Q7Y
TSxbPjBHjQx98xSaJvXJCAR0mOrwL8DSEb9wdhDyojbyUniR1HV80lkKw+bn
u70oQtbRtxglS7/JIaSZj7ttyQTdNm8tAdyMSqtktUhk/yWq7O9p3l5gVswG
TfX1Qb65ZiPAYpU3W+msUaaWBD67jllKMQBLrIijz+NxT1sxyb+Vpug60XnV
p+EpMWuYLEBjeMSVKqwoRFIZAmbM+ypN48ebs+3imj4oasqDDn4m3Ao1nlI/
fuwUQsD/9QgDIKDG315g6rlY/aqeHuGNj/1tAuLXnj7TU4FVJcdEeC57tfDS
tmA+PgoN+eGcplqj4fNB2jBZytOqvI5OevgA1SvFPcLrxAdI2hoQsYrz4Q2T
uMsmRyeNy2iMUm+9gTggLe+hp2wL/jLV7s9FoqbG9DRqrCtWRyYN50EJ44qr
/JZv6mcIXIwuKiia+7KZe47o/Pgqb5fHAZLbY9xNCio1HG7ftGoTNUSZuLw4
YmJJ/7bbIywNETWVyunJdr7uITPgJplBTLS8knVgTVXZ/40IVUnwvPFhCSaB
pMJpUbMg/dIGDoA2g5KP//ddKuKyXLnR8RJDZhz0z9m2g9AqC6mMtUfrj0pX
ENeVVv+joCijAlXixWrgvRZrub/NNJQPlVNVFwGVZwt/+e9mNTtTNf7A+9b6
FmMG5V8DyfxAWfQacIwxqt09hbeTu2L4crsHtoHadZmDZ+HiIj3lbid6cWVe
gjT/kz9yTz6Gr5Nasxf4czToTc89GrdxwdU+plYEnK0i7SxxzgKVoRggHeto
0clVjWa6H4nbPyiHO78NJJED8elNsRp3LBf8c3XNV5CM/+L9NW/hwhgIV5pb
4U4qTLx56C3M+fDcSRtZ016cgf7LeK/ucb+c1UZeGhccH0KiA0oDlGiV1XG9
fCKLbK7l6nRn7ZX40q7iDlXjZfF/sjU7ZMesvG1Yk8mr7fZzz2UUUXv+w2sV
6ObhWyXyq3F78+AAAYIf+urkButZhG01H9GWAREwW9JUBiDReapay6IANH4p
53+VzLP+sxkQRGvrKg2yc4vjWofdnHlq6kicAJpqJtG5zODKtuxE7dkvwVqV
WRiaNwWBJd2XVqDjgH3iOfuTmz6P7emR8aSDmrjdThZUzxIen355wgeEpXig
tfo+CYs5yJCgbl1zSzCwvaoImgmjioxTt+cMUIt4ekt212DQxWAibJLdVN2+
FYcAJ4duONrUt4cI7Z8pRp6CVcxoIswwd1PI6FvTxEYkiRAFUOOkn+3Mvi44
6BdShdIKDfs9zDcXzrTblY6Y6PdNgxAOzEMcRF+XiPNflrk+VrelEXa1czFW
Pi9jgEWUXrVr23O8yj+KmuKoHF5swGkj5B3ju6/sEyoi7rvu9qmO863fXTPJ
2io5Ts4fw/CwQ9+zOgHgCUCUzZbUzjrpIJPnuHf9w2x3BqK6VLRzcEQfHxMd
N9zaRKwpUXxDPtvmguXT9gNFguHRciZOVKYNorWTvLeVuWKmvcyU7YQYu9DL
3ghqGYJ0eRtgPL2L8hYf6BaLPLI8QF18XiaInGxckl+CrBrcyPEKXN6HaM+s
E3mYRLJMV6k/Y1iKHCnUF1PA4bIgMndFSUDt36i3XyjJv138cMJ8Aczwbzj1
MBRwEQayHtx76W0RWeui8Td5MwNFCTmOlDrpYnMDa/32WHEUBlpszghjoNHz
C2lKMsPxPdkX7MQ7dlON1uEu7bfIFb95BllgzDxG6KBl3MklRyreSlXGTctg
yfzm0tDJTmiX5iUKCjngsvXxRCAh3EHKa7O3thHk8FRxAxjOx3+iOCT59/rQ
BqzWLNLyx/Ygp/bKK3a/wq6wa2flGGrMOWuURa03qtlrH9roez3+SX40tcK8
jGlBck50xJftjNh62pWRy6nBLn0IdV1R/W5SL+aODKecp+X0KIu2LV1HKTnx
r6HhCwTfv2ZUt4FS8zMo/XEwG7YFyB97N1gXb6071gvZUc2E7gmprBzOjz6O
Pn1PEfFFWAlsNzk9c3sWoRKGM/Ay4dikrXCCpqWuVixrrXRuDwwVcyO5QF7n
box4uSdyD+TJ+YJCHVxySWqQqDncftggqktPpMdMUQJdMC+W0Tm7eIS5QrIZ
b1KIWbGAOLTG/NmIFBYoAd5vqS7vazs2Sn0IZzhzqO+TLlbIJmU1bHdn1Zv0
/mo4kJRSIZmFhkykdD8T6shqj8xzLyVSR7VGhGfiDEBcM8vgpbI/kWQgKGEB
jRyBZ/S/aG0Ikk0ER1znc/1dBK4V7CeydLggHfoqhCO+084+8KlzI/ak5/EW
djvB+D9T1y/KD1MCqFhM7FQJoaZYKGcZgVSh/B9UO10jLerxeFK87si+1zqm
Psc5h0nXEU0H8Qijz/6W6jQeDeIoh5sDUrx1f0/pr5CJgxFCO73tRxi5mwLr
41spbVwwhMDe5SkmdOKcfCDDcJU70KrAKqiGWHf47w4e9AjCl+l2WBXY1L5l
D7bhxhpVJFSZZzanqlgNoqGpf765D+9UHIqVvqLVWcNxY6TDi1NZeYcyC+HX
4CVblv/D39diLN99NSSTj4Phx4OcEz6j5D9RD+YImE8naPL+fv3/LyRxs3+D
1ssNNN557BVLqUpvcWH7Yr0yF2XeCer6PkXQNnlAyoboIFaWkhhEZoI6gMFH
+Y6pe5KZfhtQx4l3jocxFtJxqY++iNwHKhAh/dc1sJPbwgZko+im8E5zcs2e
/zaYXxb1Ixe0Ix7SxNXn6wv4unh6ZP0OljJVt7ZZkZ6yI3zYTfjT9nLSF4Xq
d2obAR07wIIy1GrCHwT3iT+BXtlZ/IKEgqcBVmhD80ud7IVwLulnYFPHqUAS
gmCrQZ5XhzjcnispallnmVcd9Kq4TQSsicLDY3KrCf6KbREM8h85y6aFa9Zw
Hvm/murIC+URlSBCpqI08imCHSGWfmVXeUOzp6aqKUo3kNZWRB3bbiqvUYdu
az4zh9Q5CP/T3HIksvz37EPVhSVkcaIn4o4yFz49dnvEWqTHTtmzBV3WsGyt
GWU1DL7KbsBoVlzKFHzgPiI2YWsmXcVfEqxycUvrbTRKvq2mjIMGaQFxiPxy
0mj69lksf0kYIonAqFDEyUR7Yfuy6yIQEyqtYTytR5WAxyXwr2m4I/8S9gFl
MieGmALtWDnqYOVlSqWTIoZ2drqznE23J1sC5Rnyz7BT3H77t0vp39P1HhE9
DG8wi3pJV1uEB6h2Mv6YH/Qp2O0v2qVlMpjY7PPV6c4eBPHM4niRHDxjeauH
Qw14jtG11g+parQsqFOj2FjQLC0hjnyqhsbq+expa3sP/+O4TCZVihMz1VLS
xaIGccwLAtT4NJcfkSEGps8eXWFd8JBMx9wFyB4eBwH0i2Mz+dNqfscrA7dy
H57nW/I+DBnyEAzntJ9YjoRnoAR+jUrBH8oLfzcvKCTxrwB86b73NRDyT83r
QSdNemjs6TYrec5CzrBjIXPoF1OZQbyQ5beYjGHK1sM0eNQdumJds1wdi9qw
zLfeyoZjQBrBqGihQ90XLf/JTGRfA114WwBuBOdI3hsjSTe/aqTq7wdC2ZwS
YGDoNz9ZW7sogDUZmbtgdCPaaGKpvYLq+W8qP8h0kov7AiNPlICzLtqvsxwy
3qrhdIMiIxw7E2PGGxk+mqrYOibHjsG//B3Kuqv7mjH4mqMXw61+nNICPVNH
XF1TeKZABlRFzn2sc/mMI4XccotyI5Gx0EBvXkEJONYguU0D7/M8vH3Cozgh
ttPwoiAE5x3IA4Tlh/LnpYX5nNaT9EvYMR4EBI1bJ7vhL2NGGt7dCRzpoH9D
Y42q/HnpEu5IMN6eeRgA8x92GCMj1vQ97sZzmxk0ynJ+Wk7XW00Tek7vJHtW
X8v7L2eSn90Ws4t4J5/JIRWlMuXOyRWf56Xtw47SUJbPtfElk6yeEo3AzVn/
xtZnpLDXku4YxWS1eY4QiTaiP1n9Gx3lpxsEfzQP8S9Ct+kNpDtp9IjjHG5N
bdGdcHCFy7q/48lL525GCFb3BwZztpaCcNtfl77t9Yfgtxgt0cRk+VHriMtb
m3Oi8tnW4rIzsd1lMiIat13k8JHsgXiXCoHFak8rqAkJEpU4eSY3Azg0sZAQ
FEQaJm8efViUHsWhmBAyRrUF+iOzqQ/1RpjdgD9Joe5CD8l+HKulxXf5s4nK
fQFpX0yAloikbft5zhP3Js1m+w/PPOsnPAPwgdo7sz1FmuFsrhK186HNm8KM
6bzv1dXxSA5RLfH1syBvLDzYX9nPMC85adOX2tM0yl1q7hv+xiuojb1sNQO1
I9HcSXptEC1YBYUIpRRK31tOsjm0Ju4JDZ7Yv4aRYF+On9WXiAsZRl/BMdb4
AWj/EeagcvnF1ruEMrSlfTI7WYprHYLWF5wLtZlEkLTjs7qPQSeAJoqDeiKO
oFyejeT6FDrs4OjmbgA1XtzBbB9vFKcJBEmhzMdBneF0nxcE40z7qu1zbpjS
zY6/AFM4dB4OW8KbgPXy0Fz28Wku67rriq262x8tYPCIQAESpcGppVKLZbY4
yF6Kgwg/4WFKQJDLXPcGHIPXGJCGjhvtrCA+SMZhlJcgG02NYkSilwNi0FJX
i2MxMIUYrqsY+rox1Q1mcGNuwbYQB9Ur9HS+wRRKqzB+BlMy3ow1WvkTv9Q9
pYNwvpvSTMZIfWMrbdT19ubyV5sNqZ1rAWi/iEPm01T01AFReUec4Utx0AYy
6rYJuuh5JHtMiwJZPtV34Oc7vNvqOIPX9ZCinhvlmFZ/ZLT7bM0kVQkT6DU8
zWRhDvx1IfE2yqONtSzYL7IvnpUtBZi5ue25tIHIZx2Askc/aLdIWxa1tvha
npTzmmxA3DymjC7Rbj4t4mgMvKN4bWZXNvzg7fckqIaMXgGVJJKGVCwmBMYw
Aqnx6mmOEfD/uhxOooPCmKHynr9att5OZm8/Uv7o2Ecdk7GkLVixHpOu0hOi
JKW/bEy+rM3RXhu4eZycZSar2bSdP96WTkHJUApKT9VPhEhTLvXVDwPQPUKj
iCREHduNNr7jneRs/s9dTMfFTR7nAOabQxcPnYspDRLMMo0rsi86vxzivpm8
Rz7E8ImZQ4qXm01FKo3Thg/trkdZzuv3Jsfs075hAsXdi6prxO3NwSosz0zY
NmVy20tVijrugbjysg/P91QmGLlRQ9sYypXkVoQj5IXREH4ToVbfhBq9HmEM
go1Bsiy28ngOTLSZIWKU7nef0WDtWRs5uZM5vzjuq0XXQzmAB8+Cu4dotXj+
3VvE6cxLzIoLhlVThXMSk3Uqb0Ox7vS5+I0w2YhUsEXzj9y+qqrspn3DBtFf
b3NFoQ2VC/3uXAxXcEW7ZzlINPdiBvIn+8FC1FgcYEL1qm6LHh840DBwQMbC
9lPNXVKeydiPLrn3MWLhUZ+AtljPZA540Bcm4FZCYt79H+UcvpstYCcrKazs
CBNH2WCCbUKEr2zVRcHwfcDJyEldFssKzM8UkenkdGFyBuDkHDP2KC5TvtAx
ckmlkvsXcTQTVH6L565+s+W5B8XEGS8mQJ4sF5SdJSj4cpjW3fxSgBuTBT9y
QgvyVXr1oBk2PI60UTx/FOiIvMss4D7v7gmlRXWSjUt32ZxEH2SplVf51qlj
vzYBrXLLajENydPmODe6F9XkV5xCUyJQ37XoN4KAFQZT1rbYJanr9YU4lG5h
yv+kJMlyDlD1fmXZVqqpgr+urzIWCU3TiuzOimkNRJoKde9bu/fngmb+ngDx
QsOL8uZB6ErPevV8UG2kscvFxaWQdMW9V3s30AkmLY5nT5fbQZRmiRQRIpQs
uO1tpYgDBRCt+AMHZ8xn+aLt6CvWrWC6Pnyfn2R/sDlUChsdtbwtLUL5UtUH
dEu9qYvHJiuOWU2Dg7UeOgwS0yY/Ck7sqnF28XrUGt2i/FjvY3XtTaoPr441
zE91nwaXtIxz3UxlNm5Ig0VqgfPoLlLwccRCtKB5F1Q+GAosmHRQrGwkPjj9
lXiSgKetAuHYmsLYjoqnSL3u3XUJ+bCDiF2kNC96531X2CmCdt9MxKbWL/cz
HCeBpHECypI1EjWZEUXyEi27WjCJaSrMYqjt47ltNJ7xcwFNUZe3ypndrl7E
llYSXRkxWSlLMq/Quxrhtk+QwdwZXOSh1/IpeF975UhfScFpLk6LysBksXGQ
Lk4mG33o0IaKqzgR+B75Xf7zE/jP7IPee+TplRvlu/wqtmOe2ve1sGn5L1lv
hJMwYooLQrsGWyZyFVeAU6fU3t5CTRGk9eYb+9b3d3V/Fz5sBpWu/HGtxj7T
+IUPuxt6woR70lqkV8KtJtVgYy2bNSR2U2S+FDUTpjpx0k7W5xHHBLQi5zUn
kVQDK9MYrNLBJ3YrE3JThtSxgnmR0dstMd82yvxX+U63Hi66tKbpgSuR36fh
HIonEgxkR6/INnGHA8u8/C3KcsA10YJBZjMWfj/R755AcavOapdbXC14nfFL
pGj7caV+sSqufJkAXQLoMuZMKvsF6zilVEIgxCIbcQJdDMi1PEmouMXuXj8w
+Vxl+eyB7vGN1oyxlfYqhdZhPEOxdOa+9EOpV0vLpFEyRd8JyWgJDezTuLmH
StPQLDP1sLwsSQY7mLFAxs1/4qxP4vMj2d442HgWlj2G5l737VAg55CZb1UJ
Uk8wU/fS2rqBU7C2jRef3vsWga7hElniWwxn5KZZ9idJxboFTyaT85hlbv2p
JHXAb7WzLYgCHUWRT2hi3rdlACk1nSamUnTEar5Heb83yfMF3E/XjF44rAKv
TnKtkzM05Pbdd30junDuYkvcb/XOHjEAngjJD+KQ2AOOYKi9ROahrFY+zS4V
oCutKbLINETaWosrmGqB+2jUVnBml0P7QTB1U1iiMMRV6j/YgNr0J8A7Erj5
NStxQLEw5JtlfTSeCTRvDev29yJOw7dW/K3bjZTSHv6YM5r3v+k9s0mGUmQ7
wfyXyIcwvyQDu+1EezOQcQwoBN0DScDME0bAtWSxoQmdoWI0dg84QRs1oPpd
F/3Go/n+p90LQ7uielg1CrB94gs9dtH8PrCTJ+nxq+3C3nBr7GoJln0t1UJI
vSpkZxHJKCrfc1L7BmZFtiukbnP8KL6RLCmp8nowWLCLbA23Ztlrhi4J6zWI
ppKfXQzqyH4sLtKOWIXP3j7lcSR8SNcTyN1vvD8io+r26dNrJYIYZAh0Frt5
rH+u9FxwHVVpgbSwTD3bvIMxB4ZOnjtZl2lgNmZD4PSAyl2q7aFWjNveLY+Z
mItndTMHhnCjlNFglTQ8aA7EWQ40qSH3fPrzINNamX38WHxMvzyZgSXIrw+7
agTiC2Yzc0yiZwOtzezsZ0rxEnQkwHokKUG35D+UeWP6OJIr8bZ5wlS0tkrG
42hXxyNsKb/tUTPSoXm8G0qZsZ5UM29YGAgId7WCporP5O5y/AMuorBIC+Pc
eBDI1xRueP6dv0rKN4ziDBs4bsureammecTCu86cz5+Ky+dj30ll3TP63GTl
xiiu3lHwy9bDzqL4Di6BTHtB+guiH/aX4ztmbtWiKxXFPVANr5khvsbHOSv0
JQOlkZtUxV7bjitrgGOZ0CRaMv9la5w/BPCj0k85oHN8H2bYr90awkqOoFFJ
U5wxC39Q4OVCPuimql6bbIOpjwd+bsyDaK1ctPaTLeXRIC5ArjOoMnBVIAiM
DLRNRvjFEUWEDacAP5eJu2tBbRp/oOWNt58mQOFSrFFM3jbMc0/nG0y13abK
+h+EKHLivigV954AKhYw4v7BLfzDyuP+LxDQVQaTMOERzvKrM1bEkwtbsnUg
xoiS3OVznLhN4GD0iBjFNMTX7q7zstgtZjCx/8F8XIjI/LAoRJjbDDzxVfKX
s8MKyGTs5KM7pB8hRkdFZdVigNp8POXjjWcKoWHKKbpn3ur5xRpvdDKyxx2M
wm/Ni04vcRp3lhmm2DYfypvCJVYM1eP8hLOtNn4tqYYdWwANq1w4rJmPRYbO
PqqaYPoMJHbjC7ehLr78CZeahCQzspUi5iKu7u8yygpi2012O6pnYS5hapNf
WdqModL0WL8rMuHgN74VW2aHBMxO/vd44t06ZodL6pY4SdtlMDU/XUOMoLB5
052PmiRWspdIFiJGsOb2V3KxDx0KhIOIlQuxW2h9tn4Lt7a7kwHC2xZtTn5P
mv31NfRatMy5L5IczmrWeX7brsOE+znagCYnx0gG15paZnjpKWPDhTihkS3a
mi1RptBinusDhN6NxVKWqdKTtUje190JyCqmbg70eqQFQOW0E4LyoKvBitlR
H2wMI75ACa/FdO0wrRunro3O0ZNfH23wJ1AYdnt3GzRME88h4uoB4IbbVH5a
Zov6wN7gIKp24WGKpy3lPsHfHvp39Htd0BxmTqOvSKZBFXzAZn2pkBiRAX/t
5dRE0iv9zCzHt/s/JcshQaxH1AbSLoK+DKCnMAvGkzk1VzJTbQ/GiI9xhIEn
eXBTaFOglobwxqBlsf5D4gnx63oqymxEokLCitQP7H07/1qXoxQwHv9/5KJ2
G1BWtP0dkYrONS5rFZ3dkzMRiC4eED0mwckFntBlkO+KmGTdJPogLN4g9QAp
dYpVIE8v5Pl6ABAVHawFlBNcP4guwrP8Nxu1mFINyUBih8UFJnZ9gvWqVdz6
cQbkbZ3Vi2zfyX6ZGSjptTe/Wi9W4Al7CqlcwZvaPkJBM+nFjFHSZeFS0vvH
zWaHpfNE93ccdg7eHjX4pUkkc+u2VhZ1/nZcIAHbxoRgXu+aHlBJaAR5MRq6
9AmpD405bfECNpxz7oYePhObf/nneWpsEqW00aVn9nZqB3Kig7UNRKmHL+Pq
h4jvszjLWIGuPajGZNkXXNHxR67BycT3bAUoGQ+9ZxmD077qia+2WB5ZXccc
V0WxLeZ7UIyS/7Pk/OhAHoUI6p5AaOSqZEDe1i+8L4kwWdKyK1as3YEEBA5k
0lcs8ThIg3AMTo830RAbP+bG8anq34Z4+D33Tpaw02v4H72k5Uei+QrOaSXW
tFkQc+6KuEyFCeUVgppaOrd00PvaKDYIOtO7tzX33Zw4U/GIG61pNtXLLKNR
hX7IaM+ihB9mpBJmfIUcjId8yMk8rEGB6fRTxCpcjX8Q+nQHlnZtO8j6E9QU
CopnF38WvzDJoHNDa8WYtPulDLIRuWvtgT8T+RJcPaTDwGMi9DhcL/oai/HQ
2Wlcs1Ck4FYdM72ztZOryQrcLcUwiRtj8Q9GWISq6VB9qkWUri7/wWSUY8O9
Q527pgmTNbP8gyg4CXpImGpciCLvTPLsZAuJDmJaE1QTzIqQcJSjRGtzd0ww
JpOIQTB48QX3x1LNYOGF4n2X2AFDiLD5GKc9CwEfcKYsL9qEPsrNDvEeMtIO
mDmH6Bh9lmz7qduMgTHb3RjGmx9hZT3LeAnAnjMoH1pBO7LYrfucS7PjS2C0
y9wpRtaSw/1pyXa20fRZzeIu2Cs/SgPyzyDrEDsL3mnbcOwoTvAPUqj1dIoT
9c8k3mksRKdEW/sIv/ihIVZGWPknzXchyfShhI8Z5Vhbh/1vmd+YBhGwXWUK
RL1uG6EYYbvL1Y9lNsyNPvSw1vaqCbZCvhQuGMqYqc8MhApQ/WOQmK9Lgcc1
ihjruhieGC8XLTifVDPuR4Fd9thWPO3lk+gP5dLxK9siHDL4mBl1DTgnZwpe
q3dnqvPN1snuESIxqG0hEXnPJZh6T8SU5C9ahpF0qhbc6KpHqQ4c3gqPQlAU
DSDjRYegFydQbXRniZ80eItPzSo+LeJOgmGhKnHcL/flhyfNKUXMOALSsr/p
rlTEEEKFT7glFUy+lVqO4hqDDloSh1UHykMrIfSHyrN+5OmDawMw3PkZjrda
x2059JJSkL4kTq6bHYIsTrggc5eK3fSr/GC+m4LI8iEUI0kSTlv7Vcc1MlfF
sp/1bJ4EpCDiyr+On8x4isXvU2Hy7+0AdR72dF+db/k1nKr/LbWLSZdEP59R
PgQCgoGVuPpdW+lCYAr9E7v6+I+Q5F8XLlDJYM2bcCNmTZrP8fym76IbYPMG
9iZyaaIQPOK/2ujT6HDi1hlmx+d54mFimh1Gz0Tw9LAlM6hsv14yR2qKzkPq
63wwlGVnjZa4QUyWC1TsTt/uhzffil+gsdFxSGfBdfNCcoK4ruacjVMfwG/G
1taZMPkkf2/IhvaQGqFqE6c1nPY0MHHzuCeeDiA8innsF1pYRXIJLPgWy9A0
6Dw0W+eFbP8oUP5N0GX/191lH9LRfNGCLtMRZfEbxipOT9Ps0IRWN1ICg7OR
pe0nnXQUsop0CfbGrxuWjbrTQmTsxz3DoLVdw2lTmpARVmcJmcpGr80Bx/mp
5B1Ymkz/Y0+Ab0ns2lMYyQw1SmjnCPGs8KmYz2sMWYsSvmP3UabJnL3AT4ra
4KuLFFGGmv0o8FpKE0n32MLBVgWeJuNMHVPS+o39I7b7j8dqI2pS4+ZVfM+X
VGrgd46Ie5h5Iac8Ed2wwubYYdOfox1+f7xO3mKgzFK8eFP6TEwWmvv84EUk
FwagpVFyV3GNauGTRxGGjImdt7i7O7FmO3BbvS9X9b+VPdh1/IfVFVBS2ISL
u3hES1cYJcyJIL72JTUe44OMjMuFyVkj+F0N9RZM05iRCIgSHTwvtj7WMtzU
ec6daxNlCu4TalqxLlH1TRQIVsmuU1tOIgSbhF96RlyzxxLUel5hc7gnRuBg
RMZxAeE916c497ZJC/V3C36YPLhuXNaZGyQz6AuYCE1lJOpaK8Eaa06P/6Q3
o1nvbWMgAEQpMhvb3gSCxGoyLACvhrxlRWy6IlF+jKwS9dUnDLpZIvb8EU0c
BBBToh0s3s0ZAxjvB98O77kZsgb8wFlo/8rj0lx9BTDv1ml9L4PajOVf+QvP
vlk9DFOCK9rR9l8A0l7Cx9NYB5QBWfom2+PUMGfRQ8asRnpdjtgCqnbwIvGb
FpiVJV46Bg8tAqdBOZBdILEmryf2Nyrl4+ML0gRaQpCxlj9vVFjIy7gQklfh
+wQ5rgobg6PTQxXKYAbremtjELOpZ/lqLoSG297y2F1GcYp8jLMs7h1bGouW
7jDSxCOsyYBYEkv167j+B57IFjccOBwN8j23Lok660tRIIyLoNHYMlWdqOL4
6p7RwhDmjfrm8jxgxYpDeUVzvkjYisUs1TwY0lCr8GsvuX3hqRritxVNJ/cE
2WtgOaJ+YIhzFQNMusteAjaIwMmCFKkE+EykrVHU5tzSYMs2LGIjkWRBMTBf
SaYHNJelQP1s63JqvHUzG0kHW8tCfEy+xvp+9eCRLbjSXNWTPLvdR6s2teVa
CW9T4kXruj7GkWqby2HtdXR6GNBvkOuDK1N5uCRSjv5EBeMnFzjmONU6a9kl
2BNJ6CeTL7Kkw9uwdh7ebha7lmODBWYtGXjz5sK8zhtHyXkhYQqEDuui1S22
cDQ9LheccUQhY4+uB0ojeKjmvpoefqvHOzeiqvINtxrbOmP1KnPk7M7iQR9l
wbVf7Pd/hwEtTKFINN+b4eu5JgbA3SV03JTZ79uotGhdaYAPTzypCTzcyCg6
jnhoJo+cdUaAAq5OdT43I/AJGgbiPfaBENiEt3We7EEBQTO7SjSPqgRZRJW2
tNp00ueAQ14xiKQYxT6G5M3k6sVVl/Jhjssl0WyFGBexz8csb5gUoaieMLAr
CKyU+XFW93q32BxPs7Cysk5vAHTsCThYqojjIL1vgA9NHvgGOdo0T/c/u6s0
Nt6oCSQ2FtZXaLk/cgG/w5betn6CqZJHJg1sPHQp+ql5rpnvhbVsfYLBsJ2n
hTWkfr45tQAYdJ1KxJ3Ct/4UnniGERTHeFBlwSQ0AfPHDlsjk1D7p9zNc5qa
gtnZOLkE5RYvvJ9++xCK+/wXiaj6xEHkKmMCExXLuKQPbgYsgpA/d5Ojy3V4
mWiDcdKxh61HDYeB6PPPd+3j09hk8BepxW5e9XtPEixQq7eDnWIg3CFm36cx
YzxU1M8cZnIFqKVM5WTZNtCQBWSDKyB75YLB1HSTnQHb18QIqMGav3r46Uvy
d4hJbige4YoksDARXFkKIkbfMwL49FLySvRFM/HoOz4+FmFZAZSDjj0M76c7
ZapkKPrh5XKkwcVML6isaPc1kb/dhlzJ8ihXMGtaKq8xeFKP2TXGWlXk23Ez
rRfKC5hj8yR2DMljsQoOeSc9B4CHZjKZUcJPdWzfSRJprNVpThu996Hd01Yd
Rr4EX4nhdrwFvSs6FWD3BdoPn7MeTc1zY9XjOYqn4hYP8PmqlhxMwRWDAvYu
kkU1hbvO9rVN6qjH4KR85IjqJfTngavHDtZTG81CBOo8sE5PfNwsEFKrnL2h
yeLG336ZuyXuWBY7ORyqxBQrWnlJD7kc9Z8iZ8+I/8d16ABXi2gE3LYcQNtg
Djy5baVc0IfXiyFK+uxri3hoLhooeKoJec85H/zQcz794JUwbaUBFSQj4OIG
HJJQ6rBJ1Z2PU3qkUCaGLF7D7hjzfP+FV0dsLN8xYdL3lDc9t2RkkfMCQmn9
uAdZ24gqSY8/e/uzfXDmF19W9WYrMoGaLJ6M47NM64Ik5ttDLlp2IXLwGkkt
k4Rya1kb9+c9la8jvRPEcl5hCCy743dyuLebZYJQZRZwMU+l3L741mn3uKgg
5DUf4hDjjInj3Q0ff+tTHMyVr+2XKnRrqiPIKi0659R7Hj3Lpc7QczWdEQPZ
f55vDoYI+sIjgMrILoo929i4eq1gFwS25nK3igTG70alVPbTymZPayOvO5NI
QTLhsYGpsSUE11QdRXkdWirA66Y8WXcs6FMMOJIXnEcvbOX6NSAOtcwZ7KiN
HDCjBT8ujX7rm5N6okMfhztZ1XJWSGg4N23xnL0O2I3LZ8CLitRLwt2CvZLw
9AHz7/3s/74f9FtaXcxoLYOjzp2Op59szbWWf10UW7VqdyAF1K7bMTZO4h13
Wwzxj24rMtBrRndQx5jy+db+DrbfRy/wSUxv7xAlnXv0xm5wyxPBUYI9tGV6
UUWZ6zXrC/36kS8yXgriIT2HUZ4Q9s7+HvebaBeBRok7A9e/Ups40i+ZOoU9
CN6Hf2KVvxcrbgdAFHhtxQ+h0QUi4caooUBwYO0Yaiefqyd6EUqEIHbjQSE1
tVBv98lUKtKKaeEPFRQK84arbskIPRCUc+1ZIbZOMcLCo3+pFxNVOKf/O+PP
SL2v8Dv6PHQG1Y+2YRdC+F3wnsUPKU2aw29kaumj+KrExX9av15MvgVLBg8R
1IdrSE0S93uuk7s8OsvF1nhB6ok2uzPcKX39VB8D1osOReOG8DIPzTX5aWxG
t62IKwXFdKyYKyjg4k0cd4gTkxoKTjtkUed1hIMcV0/MWoSqXMjjCsoxxwro
gR0K3si77qzrkQroQU+qHz2svSfzp9lRlQlmRnPD+rS3Ghip5lUBD9wpHi2P
iMdHzfUHgSOwJLNLrv6SdCiBcOs4kABuA4XlCwC0Or1dhMCHs7Zo1uiZTfNS
zu+tmW7f0RR9VOVeSmVcG7Pn1MSY/0xkNQ1wfL4syW0h9hWqTnq6U2SYcZO5
7BnTPl/+UEDJaKASSzZLbTDq9xw+22u7jeobQ4NEGhKEXlXlsAF5z7wULtEU
eMKT3vyoItIOS71/20XQbRKsWDbnZKuQJZiagSO1T8a4LHGKF34iVP7RM11J
5FonuI8tvkz4OtSv8odI2Z/zuvINPY1xDIh4SKCLMfZrHerf9d3ka1ca6+4T
MA175lEbffPinLAs0dd9gNOCurWTcWcId5p3uTPPBri18RxGYQloH8szP4Xm
0VSVMN6KdIx/Ui28yQU//moiRYZWerKIVhOpiXGQYYlYKtXoUCSk57dK5Uck
cHGjGA4QuHiHKIYuTQdd5XBh4OL+PvhvMFXnczrgSfED/vm2VtprO7W5RT5n
j3ycWVPnionYtbzOe1Op8dUK3rRfaKLsAIqN46CLiYRz3eGcKeN9lD1u6BTq
ppp0JvtOmyYMhgTkM9GFKUz14FaUpIdCKIvPq/kCaDt9OYm1cBBnCiCddHE8
wMf6Fg0b2Zi1rMFQ8cSjh0qLwsq1mF6NTNP8Dh0tSx0RvCW9Mo/y41wO/QLq
ZT976RjeHCPg4LuuL+LEL3kfakSAlEdY3+wMTrvRZqLMheZmOqMWmbh23M/J
VKZvWhWmlyRtFuLltIaFgvZHfMTVGRFBpnphhiLqObDPGG1Ya94AAuKMyC1/
IkQq9ivBerCtDfBVib6BvtCdI8V8K42ZNv/H5Z3zG5MofXjIYG1WwB9+9fVq
crc8JWWgZtSrTz/1FgjbeqyGcEX8fmXVX6Op8EeNXixxrC6msiU1YJmR1a7c
1SGR4ESKjvokdPGXXwnVZj44FPa/2/Cx9pI06WX9wI1yABT861+HrtnxZ3AC
po76TRm5BO4tnQxN/mf8rUyhZ0LLFvCV0H4qUHGg4dBcfLvVAnvWvxfYEc/V
gDGWYZ1HJIu3K/PIvLOfhTYOF/tIOwBJKvhsgfQp2dvDXl+2CHCAgR/m40VC
kWhLPyQODgOO/Ny1a7p0lPJ5L4x4SCLPaFcRrRgb4AsSIZYHWpMWBiaCu8wb
dEvxilq2zW6DAJ1W+1/NgQ9z+gf8H71eD1PcNCIEM4u+TJ/fpA6yLUnPMVau
yRj/ApXzN83UeynQQIZPx545qSrVSNNQNP/VF9aQleUal6qedcTBvLPYOTYa
VWE7exxjjoi1iswWy2o5zcIykBS9QpBbdUZBeIn1EuqSVS56HxKpLYakYBZd
3Tc1fHb+7FCKQLMjPmFkfk8lSBYeuOLisBT4pYnalLVx/I6FZQPCqOTCmuj1
0hv6udIHk23kqGgtGvZ8xj8JGUAowJLgtl0ok63SQycNKithXX0oR2+oYYA0
jU+yj3edqPFrAkVhP2a6lWW8/n3z8MtgAAdLDLcUZrnQD1ypPn0wKksPvZ9g
UkPLbpQcb4EC2T2bj6mHDUxUJOzhaObBsGfExr6JUk0eH4whxDB3GCFEg1lB
WWJ2Wth4SZ12ZBDn3uTQO1+edKzVElfzkCi30HkWJaY6M2RV6ayi6gmlp2xb
A5+GaCzYQbWc6USK+ij1CRDamiWMmMTp5tQUxtNyXENBFo8lJ0w0wgHS2yqv
fmfxlngmuaZfqc+3slD0YR+sarJHtDuvGpiypSWSbAtLM73jqHLnNYNTJbH/
4cEOXTa+jmVEfLiZEg2gcdWNKTvajwPmohRhdlT3iGNb8CRssD/ORq+I5OOz
akbRLk1QfUbvklQHUvi8fLj5PO0BP5Oqvqnn8p/tNV3gI6BRLPlIuhSMVvoP
CdBa9u+T3sL2lf5LKBdAszmILdcbNlgKZ3XCsbvdBzyiEMrLBUkF4h/PHQ1f
kecDeM5wagQYay8qyg4pGP4HjfA/wrGVlRbGf/b1USghAeAD4XlhxwPmQuo4
3V7pT/bGeF0c5nZYrJ3CH3rCceIYfLotRtxLl1pfT+p6/Yl3TryfdY0uNwFs
IVOGB0GT31iJUjv2e1tcG3+rkD3vMCqQ2Uacpdor0sqFKv3xJdGOCr8ZjEOK
aBZy4MbS5ieHYqLRnBml0DKOWoVnktW2l06AqpdoHiG5eQu+4gceWTV5Lnah
1OC3++gu2Yknd7GYqZ7rpvGPD1Lsi4vJFAJBEyls9uRqXej167NIn7OOIsL1
E7mvg6xWS+OdEw/90BCav5bQSZ+DB2nsyfdkFx87h2Z2jJYpLC4MrpOrvFpH
dMEMbUemCtA/QMtOlxFr36W763ZQC4VDHyzCC0WPvlLy4MUrZde1f0ylQKax
7MExs7hI+Av4doJq/6oX253w6xu8nTdsh8rs6aDrKC3NCKOp+4hRL9jvjj0K
Q/i0vsL36u3ORW47/SuVqvXgFnA7mb7PGSCQ1L3bf7RWBGWmw7xb3Lxsn0dD
V6CNpdbRanSjNTQyL/f4AS7duJckoxjHnYULyHgFUZi0X7O4UR581fB/OY40
WTeGRgN+GmPnVyWwYjq5gnPLBSldhqUikcHv3fKYu38JJQOwskYZonHnlVQV
pouz1xAFbWEEF73EKxkT7eaXoCRBGs2J/N7xW98ZXBw3ytLHePxbA+ioI1bv
3sS6XoRGgflaJ/2Km45Mb/fuI0Ms80oUmnWz8L4gObWaEZsCaiioVUniMSNu
W6gcI3x28Hk7auq8gh5T31sG3Ey2ZTk8FE0hVI221Ta+hHABmEccyfNNhc/v
velbyVwc2UBOui4pT0H3iEn1F4hwEpyIhkXKP0fs3nozEzaREBcyhLqFKu8c
n1SMSudCCSk2V1Te0yLGW26VoVlpXUcTv8U6Zyt83YCtg8BfajV/fDoxpFFF
4EB9dVbuPO2oq6zmnOW2t2GVRPkISYgE2ogYcSS31bzEZSUGlyRoyZBlINn5
i5L8o3PQ7zHEpfYMFdZfnR1NVrSSqb/TfhuK5Vae/aw+DgltHmhIME55aR2V
PV9J+jShtZMi3mckSwQsCUejFqORnr0BnQgGWUHNYv8y2q/fpYHDQAjHx4U4
o1Qyj5lJ3f+PNugUMFM47Mf9vzMu6HSJAGB5TeYQXP9hMJ4HCnAKcYwbVcBu
v1Ius7VzZh60vzMTUbidTWCLo9KQqPjqFo67rW2YaEq8a01dmQLZR/PCaTGA
tjtdyCu4KK6d6MLJ0+8gc8WCxKuwARJj9w854lfHIU2p8XksfbbqA4T5c/wO
hnRRK9fsR1SjJuvMv52R1xY95UXvSz94SZMdQlmdMlddjBfAR9spBX/+jkYv
2wjdEN3q4P/7/u3gMJDvLxkePHsB3r6dnNufff2BcWq8SQU9/LJ71XQMlcg4
Zbvzu2ALkvO6H1dZcyIHXDIpuBDBaAhbgc+zVhy43R7y1Aj9J6xLJQjFOaf4
224O0xADiPts1TgZaYxtxx43yTEp59T6ILEYvczzYC6Ns2RekvULl5KIz+J8
rTit5JCXP1N7MQRyqTDg+bmr1MBojMxMyH5oU+GQRO6bRmXR9GqlQ1zLOQhR
ZLZJHoi26EfKDW25vrDIqAnbqzQbppANIGD+zgfFlXocQUrTZID6goejK4Ay
Yv/SevevC6423ITrqLDkFI9tzdQCztW6IRTvlsRsgxzTYEZkGn8wJBqcdNMX
LO3YGamHFdFz2nbt1mSMEScdilnECV93QzjvZykj3BYiXxnRDIcQfiZoIbZR
1MQQX/1z2FfEfB8HwHJHvhgo08/mXA/Z/lf0ad3py/wD74vxyRr8CjIil98e
Lgo0YQOvT39na/LbfOpKeycNoJ81a7j8O/ZwKWJiP2uL3J7yDkiuVP+Znx3M
Fi1oIuTTVqbeXGXnUnthuDcuVkxpvtzIvPYbmhUCwNZUwnB+VsVs6glZBQjL
udOo86yviwa7PH91XhebHCDHRQKhpO/bo07lY3ZVEJ6zS22HVV6ggCnbJBj8
RRSeLW5Aekd+nz7Xg9ve6nreQ9dNFYrjlEOv3RXg2vNNunlrAf9rJ/dacBrO
Aos9Htbmj+NGq+BbW0d3y363Z538bk7VYCGnkxGhk1Zfx4HCXaJpVBQCKu1t
5H5Gvs+KQRiOE4/f87x8QV/xZ/7wnp8c3egSFsqa0W55omSc/hvpDCweRH9+
FMGKAsI1KN9vLuZ5BTianhufNjxp7x4Q1ttBXCE89m0TIbgjSPTX/twIe7Bf
ZmYbjKhPRiNWHinKLLk67fyxFea9CAbNoSRWL5iZVXhFZHJ826Yp7HzGkANm
v5sVqlz1s0vSwkM2/WnnPzd0lLmQc8nRUxTLoAZSgWysuDSTxgGBnvyVMFs6
+sk4UslXUjCGZf6i4G8E4MGhyuHUb01R+J1mEOS5eyVTbaldLMUcai9Wv3nY
rh5Zk1iw9/Is8QbtFBHHWHxNPb9MZHly1RywvsKVC7XR8407qYIJnsKk+/m7
n6RjFwnMa+N7/lg8EoXMBBCx+D+7DRsTOuLR6lw0KzjM6RpbMyIdatnJgkyi
cxn/OSYkcWR0qmVzCf+y9Dbt9al2h4n8W5G33+6fe3KQCBWzss8zfphsEYcA
V0LpCEcWz9bVQU9fU7UIMpw47pEDJ/uJMEiL43eL35x8z2DiyuhKNoBt35pS
N9q3cFGJVAOCDmMUBeNNHzXToFk8h3PLKmRZlvHotzYLTKP9F9RYqFGFrNVg
WmzWrk7LDHwQH0F/WTOsdHbKhWrnRB1/6ON3gcb+9FHPgl3KnrkHk31p+AS1
kunLijN3EGD8DpKARdw89CRhGpPRrXUI6Xr8uvaSP0nUrg+U32P19Z/NcWAt
ADFUrOCEQ7MVrZT9eYhI6zoa7GGsqF6j0lBfdPA4Me61yQ5X4M8leTH0KCpY
cNeiJxC2AMDRqbP9W8vfD4pWa7rT427MB1yXyUWhtzsX9R1DCOKo+WKEMVDs
hQ0HWO8KTSx7TW/WR1bMhyT0xOWMUWtBntS7vu1nMEr3doO42XV865gAg3Hp
52AUQ5BhgNS8OqShdeD+WkVYWAWyTBIv/NGFBm8flMYic6Se165nZJrArysm
HDJEonltEqyyEjl5JxUQI6EaEemF71AsaoAYMZ924IBAU9wXNm0ZEH+RZ143
D7gtLprkyejcIHMdRv2utiM4l4NEzZuWW5lRfltsBP2I+aaTHrL1QXd5lNKr
oiBlnc0bTJYciQCpf0z/eVwoLfKyJYFCpiGBc59T15Wi+r6ShlfeF/+MpxNi
bV2Fdthyr9womy9R5ajgX0mb2jHFxYOjL7pTdue201EW/kPj3x+KPlUh/AVY
xeArlWjZQSDJcyykxR090UEaVpGROvcZzXs5flGEz5hftI/ElHlNOr7v4cJq
JyEEAIjKx9dq4ZAzWtJO9J3aQhBckRsovm7p4AFDW7lp7vnLUK2H/SHgBkY5
WIj167q2eIUQM0q5qLr6t9N5KJ9ak0C8Ip2Pcy6EvBbhnh2tQNgyiynyM5Xa
Io4vSyNcm3Z5+7BqH2MgTEDY3IWRTYjsOE4+yYy/9wETaXkF8mRoBO2iY2gL
5Xve4yFhC0SCfJiCaktOd3Ze5OJmC7520p5ZdMSKDuu7DASCYGGRrOFC42ap
sWTiREGW9dhv3OdHhzXSxOR5OVrNgq5hfYYY1QrLxi42JHbBR4crNaNxOKxP
HLSq943/ZUtzUShqeCewSQz4dI9C99Ltrgk3v31vDjxwtoeOcQPUpexzQt2P
o3pGuumvVMSYfk+afKvIW1FWcxttBgb7jk+UGvJVZobjgDN7pQEEyY7MgLhR
wh6qb3lEKnMVc/gx5tMPgSLLlN7n9LTKJ8N5eHmEp5h4yMDVFAG/HEnG2akA
SZO0+i53itcAfvU14R3rqxoiGP4Zku6Fb67e6yUEtFyeA4J3E60/+PnrBmnZ
xpfH2mP2prEHiRitzmB9/QKAzg30KrQzmgGYrz5iOecPDXq/7MeXe+P0fMLr
d4uBXX7eqxeW7u/UCr3rkEIJcst06j09U9ZS8twtGHlRDizMACdwDkSipCIs
Ui/NSmA8CMmJBmXPiEU2FdZ7LbwD9uVdOnoTpB1aUYg8oXzR0c43CWPpXeDs
UZPyF7XaV8rumKj/iXJ8ODikGOkH0pX04ODE/xQSqxWOutYdL9VbjCyKZX6F
lHezZPXdQeK/zGtzu7tQO/mZvuB/AayvE6o8NnrVEmU4h5LBc6ayclw72k11
2vQCkCBYp61Y1K8gmmpxCjoGDWHM+XB52p3Zh8MlPZ9wAYTuTLvx/Z9bed7i
kMTG0pJIovMT/Ett279XdsSzMzlkgRx68M2sJbKBM2eoEMvxwwPcMoYQD6XD
P+fuEqJFWGRljaqPEgamJu1XweWpP2tNYdSNn3QzDR4cCJkke7T4rhqKDXye
GlprzI99t0ZLhpP4zl43dAUwU63DlQ50H7Xdzr2ZgqkH98Ohr+k65Uf174qt
gnfvKo10UcSUZOHKj4pn0z6ZD24a5wf+sbKsEo/7n8iOAqZtVIErzgrwN0Ah
52hbz4pXl074uuY61WPGZ3/VKlBgQRYEqlZqnlukFXygbV8MiZxKV6ph9HM7
IaNHM/J9U7E425dYqmC3HBsQVB4g1NquEKN8gDEn013CXb3lxrxA6/8K9iK2
KiwGMWdVaw8K4/3CBW1cKb2m8tD07+Ws0wJZF19r01SnIc93N/o9i4cGaG8t
SdqOtTXQrMx1XKAbnuD+ADqNf1Zq2FJO5DspTiNo7oiOPhs4zoyAuM5/G+BH
V7x4hxlQ9Xed2TxL30oJlV+fedOzMOF1bRSUIW+piZjUYviTcF5rLugm2PmB
8ErjCxps9HcIAiWBCwlqLLFvNXp8HtAY+4fi2w77J8Ee53rVoFgmvz9dMq0R
ipuw2dRl/47jr9kwxoay0cSdVTjKvWqFFxogEWK/bMfdo/T68T4o7tCfBMOL
tWQ/WyJrpojuq4JmtPPrCAcNzfOBwsHrMy+YRdfDwqzSYj3EqAMDgxnYBZ9H
lVhojM7jm0vo4ZmduBIVLudtL7MWWcrSptIeZGWZxAhKOGpQ/WQB3gUJTMcm
UKvbF9TqEnRd6CKagbNmkAfFpgn6PTxuWwS33HjM0k7JHzMquxU2mUuHrsT2
XJ/mh5IJHR643Fr5dlsMKImk2+hlsjR20wIZpxBpLopH4wlAkK+fJk/esrMW
7suFvsBi9xp9FqGNMz7HEjOrlmK0PgqfkN+gge3qDVSjE1Dhlzcpsz9BC4pY
vz2jzbDNVRUJzoQtjs9t2KmUgClGqfHvekx/X2CH/LR7o9Qg8d8Ntb8S3dU/
sk64cSoiJiDuk76FTjHTc/bvTXwQIDywMCXSxLqXhq039+FO+nuQ5THTLoAI
S+n0GwFYyObVA64R1QuOIJXVnJ949DV3YMN4YNMdbH/zXwf0i8XCO8K71Msy
Cc6XWE4BalGqZVQ1N1nNEyJzovyXZV0fhFnuNf6nMrLe/SUtUJovG29rXT0R
P+4O0vvHPvtOgBy+78u7Co7f9YVXHZZ6Rgf4KWziMoNebsxo2+UprYWj5VlM
uTA7/MNM0rqb3Ey2nv0tTJTQPKI2mCwpG62RtxXoSD+J3gVpOqigRrhyYxYQ
mRSkmupZVMZ9VXAIZXn+jQDxFoN1Adftv+eJ4olY7oHtleRe1bLkADVZm6HS
WnTHPz9DT6MTBhXjNVwzlpgvKegzL7lOIwTBRNNVvcnyUAZs8OkLVVsMwBJM
ZERpTdbKkiNrKTPzTomjYLsEiYtWp9Urm1cGkBFXiN+AZVRvu7UiHdTmCRyn
X93IzR3qw/avIga/9N1pDwv3GxjXnjRAMy2bQbesv4h6GS+i7Zdastd2Rkf7
clRVx/a5ASpHkmoZlJBcQZ6CUu4Z1r/+NjqXVpPeFmaaDCDe3e6lCCh1Poir
gorCXcCqCBdv5oo4MBHEdy3zCRMs6EAnsvu34RdnwxhaYZMHbZFpQBTQM2Xw
zGxfzsZPqN2aWypZY+GGG4Guk1CnAq4Jx35wKeY+ME/9bX92U3rfgY3+OZoU
l+NOtxWg3gNzQUpovsJQMr/9Z9VDr/FuH5q9m13xrvbKNOaPSNc7M2YJ3x2k
n5kywtJqaE6ohoY/2KNVu1l6OTkV0wuOhD8pLwNdkFtsJ+wjZRAfayhKI/1D
vwcmhGGj+x14ilTWH5kfsBgaYBw3X5RlIy1TMDK6ELse2NJsQdCf4WR8iUIr
/tvtdHCkCGtO9fAWEbNlYCuYnaVb7xm7FTPmSFWI3R+DVLgkCbqdXztIokQd
52EOdcFv/VVRpXwhhiIgoNrOfjzmgtu8gn5+ec/1k1gSk9RPdCXecYyu/8K+
zbS5SsOqv9oPbGZHLK4LDRKRj5qsEHkK/8yxlUcFnSH3m47IsLApPNIar6eC
aDwOvE1/KZFe8kfQQpKJQiul0eyu9tMpS0+EKBaLMuicC/y5YGJTImLyvv7/
zK+fainsAkOYiSeabmUOw2FgfQAvaKIgTQD7F3LRpGPCmFEK9HzBXCkza2n1
+a3M4NCK0LlaUbiwkX5twyqlgpfK18gX8pIguoKR+x1vF+kQ5yr+WBpUZn5y
qwIt+0FgS7cw7zJRb+0rMeK7ZgKnCwhLlHHKmLLQOIMsuhQOYgHvD0sJRGgA
hA5h9BVcInHnHV7nZUqGdpzFJ5t990U72trGTY5DZl022b/1bRDoKUin7LdI
Pi6dNdaCsvknLZjXfo5of0yzOzEjaFnOQNyHpkcWPQyO9x+xwKRheArBR/Fa
H+Txms1eUXtjYL6t5EWPwWDDKBQU5VbYuBmN+HZk3wfXiTxvMz2TV+P9O88e
jJopyWCd8Ybf7u+TFVbQg3FWOOwKv7etE9XGbYXqTcEBvPDtLCgCQYmYavaC
Z2PvqBX0i7a7MY5AlrATvlg7QOv1P1yRlP8cIa4824X/aPv7vGDH5qhYUgAC
BXVoNFeg+1KGh76KJ8IGynEPvpzCJVIy5qcAgII5j08c20elnLs4gufFUaIT
krNm+6GxRMdFzFWspZ9YVqFBnMYk+UbXyo7tmE00EnqiOzbHb1gDVrVsM+Vz
m5UcUZOT1BKIIkwZb5HpwudVaqRbjOeuRSGAFqmYvpEZHc3nJCDzkhjob1hq
BWpJPBivZ8RxNpHJ/McB2sIc+9lz5ynW2bZwInBinHT62jbo5QME6xN/s9Dl
phzxtuPb0zCHYAzo/Zz+b/LvFKaPyNjZn2ffhhMozlad91VFUUmbkKvIN2PE
q3tcxeg2lw0dRvJWROLf6kdXE6lhSFc0Ga43rc2KC2FHWCnJBsPJP65gupog
GFuVxWnnoOn4hsBRB1tburqDcgspUOzI08z0DKqMq4+LZ6rO7HwuiK29MtlB
eTB60e1lN/H+XDuc69WZW1RtFkrmrjI7B8vu2xYpG/NFGOyxpXkrHkUBzAfY
Bc3llc7b5TyUeUQ+rwPAv5Sh1548shJww89T8xEcVwmX1DeEx4fxzepVYsXv
ocB4Ti5Hqnb0G2LdzEkb6qb4iDYve5J3bIqE2jaOA3PXpdhCULlTqxrp8iMF
CctJMlEH5OJ0uAIgFIQ14BeZi2ysc6ROxhCQka7keg8jHnl3dYEur9+3M5Jz
PRrJqkaSurelCyyZmRiWbM7OHjkROpa3AcqN1GSLnSP1NK0ObXIoG27ewgb9
s9PTkr065aYySeOw8NTf+bpwJ3XC+ULj8it5SzVwEEbZVYq+s2AFZBzNWwj8
iJsRtMzC9vc9If3/WA2iEFiIbGEMWgzckxbHAakK9A18YVJX+Ekbexo4f/CH
GajcpddyxMbWtW9ux8ljxXJuBC6pnLo6+lhOvGUqVcizfD/optV+2o+uhMyh
oNa3eP/JSe8GEUh0J4GHYl6x+88kyQ7LY40+bKEShPoA8sm4SZQ1CWsOCO4A
g3lttGI9hQONLbalTJxA9iL9L5FbFF4OTPLCC916JwoHEk5iVnfdGTwik2dV
OPyLKvnyw3Dr3T2eYSsxxaM6FHvqQR/Q/fBZlCvFymRQPUczGBgdEtO+OeUO
g6Cq7jz2ebE//K0LB35T+YV9JnKkajAzMt8d6muVzp9Wml85dhk6COXrxTIO
0DXoTC325Eeh1C/KDT4pOBVg62wAfu0/nP7rDpFDBFLQequL0om0O7bEWB4C
EMrBQa+wXHEJOoc9/3TiEZs21PaSwxMoX/CzuzsBqqt0hq0sUkOYWBR37wgL
uj1lskVPy0gDqz6MlB8TxcG2/sqXkBy0PDWRs6gmT0Jm+jFdMdKL9eV8+IhE
RMmFqgL8h1NZEbjLlBxFksS1XpNEczlfgSU1HvmSzKLjrmqnNylqh86TCII/
DjBiK61bD615iROhztuCS5XpCM1llSMV9Cn5cFx+hBkFqFxSekCyrR9E2TTo
dmQBi3VBMvRNLYco9i8wiEson1btDpZ5tmADMruStIt59MMF2mh1xiHMAnq6
0KC/H9pROvmUPPdQJUlXUdGtgWxk9JHDLsLYnChDKa4YfCivI8UrCa4DuMwr
eYc8cSJID0mpGMko0dGncBhIUTxVhgwb5NFoj0/QqA2Sf2TsV3OS/gO/2exr
NV4A3FE0VQcYRLl8Gmc/NE+iO+A2N1k30fU9BmA+JsuGyUvs6mSKobB0uCXe
J3KKFJIA6+PPaFjsD9wUXQ1uRigd4Ju+jZPCMggyd3qHRgjjPJyVMUbf67Xx
9/ifWU//j5b2oOCjgVPepBBjponkxcCa3f3VPrdJ90ZNM0xN2BKnxKPziPYT
TTRBnvbcmSGMlLXpUivkUfHB2KBobyHAcfGmyj7oDdxCqHyT+PSQQhTZAREZ
WFyApYGQvary1w44FGWQFKUVIih1dWLDv/Och7KhCXhK0/Bl1s/U31u73Vus
JFUvyVJ8jkqs+uBx+ky71yZJ1L8/CCYTTpDnx69NpVueQqF3J3ly3yzkYnmN
lmmFHSdOzsS8vbITl8IU8S/UDy8hywgck3wAuBNCKd0IKLRXRf9IZ+IEx0px
Bdc5deGno2sXyQhqzhxB7XBlpaHGD++kAtjQQYbCZCMjx8jW6xDiUzsanPqP
O4UqVvGphqXEOV0FDfeyRpcmhX4cyJRpnrjCrKlc1wgxhOMj2FXmZBPfjsKz
d4aLmRd9OFQrAgo3S5PnbB+iZ3p+sFyNi60uoEncZm7FopfkSADxaneMzebM
Kab7Zdt+SBLTa5j1dSNdc8JYeUyoYxOiowZ2PFahPWZHyTKx4RHYu504iLfK
U/vFZJ1fK56UuO4nyxYRxreE2psfGqeGuXerAsgIYF4xm1yPtp3yT1hdU0Pd
iPqdVvLOLAb8LpgvYFTv2gdyA3ossO2krhMU1+if3mL9lSpQQpHTpEslFhRT
F8lKWqy/fUYYYHySBeU0P6xRT9mC4I0c/S2pd1lxtSQEJWEV9EMpXQERfa2a
bPazPF/dO47AkpizCduJWwmgY/EehP9vSKQ0ixPm8V/YXqx2/4Xyd/A7yKR3
FJUbB56YWFxBGyNl6qmy8Ff1Wx/mBoy+e6iNb8wSR/Q4dZBplFpIJRN62oDa
IUIPbIvI8ejgp5TT/+20OPNrJxp/o/OiM5ifpJxnUlrsfmsvx9jepYCTT6IL
nYihzGfxUmVqXTTmxvfNQJ1EbAkK4HoYmtQIJsPSYsJOw+Wh1ucpgyVuB0Kk
eEKrpaM7dd3iHhdCNHc9xKERvTbX/clFePGq1sVi+dBzfJ/KS15B5UqqDFaA
d4d0VtI9MWYzUUFtWgmzkpERE4uhgdHxbyDSjl8XX2d+CFay0OMiRASZ7i9/
tWwZnjxU/2fASaOt9ObM9hfFKwtZYpRhizLecxebW3BHITIkGWxmly2fu59V
qRckbeiFb3oxs6nIw82mjxs5YcJ4V46gddCv481kT/n7UWZ0cb/QX8ePmBao
OK+hgBngvym/RLjLT4wojtvxGBejmsc4D5GtMfVR2m2Ck66LTe00b7VAs4yc
qznI4H737PdYpW43NE+KfzUjtckdHiF8M9PzBd0OiFC7C+bC74c7KycHjvk9
7cJbdPvENYOT7VtMXPKZGzr44VU/c2aUh1ijIvpASsI0LTQequi8H1NyPfmb
rV7+ezinQSLxkhAsPyozLZEtzx3HqSd8ReEeS3wFPrS39r59RW5EJ3EYN4yi
p7JZGRwsCG/4vGVkcviGSZFBzj4fGRhE8LcmoVenEVivHVqS1QtSbXE+nwnc
71TIJXv8o5tWa2mEvOwXnHv24QxXnR78SzY2ocdS0Js7LvhjSPDro+idKpE8
Cdj9xeNHeCLjtKaoWB01DYWjAzuZsfpmwrVczpQZB1F0GMURgAyTmNfx9CPN
64bKF87aKZpdzxEbjtmRjeGsfkal1wbWBuPBiSNNjA1MAmgW6cHbM2q766oI
1WJ6chEjgN2saLe/Xkr8fbN0bMgBoK6efzyvgCJlsn0QQdXUIAk7FlhXVvCe
YQ/ojPDcchb0f/HAk6LOB5r7NNxqc4JTEK4pIa2B+/hSTQ2ChAodrwJyvzEC
TZKI06csD+1PhXj79JtpsyPozsXYOzCqGOdD+xceqozaYVbabA0GHwS2o5tb
yqAzQUCXxG/HrhSapw2kJMuKViMjXmAc1z8LkdwAtq3Zy2JSE1/IPsjbvGQI
RnZqmgk3zAqF21qnfndx1H5PVuLkCpR/onveZE/zuRJPgHPUukltVtqrO93l
6ib3MfBboAAOZukR6gD0hrIqH7vPjTB3ZetvwVyS5428/0Ec73ccO78nfSNJ
nKtwM2s9iPwxxvaiH06eL4UHqKXEhWmqE5j+7pTsR86Mr2gdehnNqX5N/VVH
26X65Qvl+CSgAVcsPMm0m+zHLdWLvEi6PrajaU1Zfq5qePSsIrpxaZZ9c2DU
nyAmeyxwtevJUu+g/4CwPDGZhJ8BPfMOJ0tq6gXbOyG5HgyBUdyyGbwoBzgN
z+vBJ2tBJO1b5NUmZgISlU9VB5mFiG0a+xuaa5UaIbV5JbT8EAWloCYrFUZX
LT6g6i2m+Un2TjX9edOFubw/49MG2ogetaG/EcNkwVSwZaMnwpRefXjyy/4D
PxPJtlnhxemUA1WB2xlDAdCwDTwJKNt2wwrGg7cvwotcCnmaBk/J2sr9pl8Z
M28qwB4wldkBL9ItfYdSSEzAntdd7rBXKA6Wl1YcoFIDduH9JC6skn+ISxol
AFh3ptDwfxlYCa1VzEjr1bJo/gcrJq1KSpaTO0DQ9vcu41dQ1x7Zwc9UYbyB
iHWui/2SrfRF3/uIa4e4pD4uBHlBBXceWWyHGx5lEFae5IkPdZw2JH6xQ7Zj
SAN7c3Y39Se33u8eeN3IjdsHSoYVNju7OnfS72dmYQlWf7v4FN9V9Ck6FSzy
TccsNAJwWDO09DEPA0gp0i31z65yTtNGkdnTF3/ytJMUewN+XQzrLYdXKNic
3bijGKUMwsZoemgwSbfe1BD3AmxEuvvzEmhPaqphBbbHD8j9EUBymJfOW2Ba
XbHJdmbVwWxZRioPlN2q7ubc4l5eiFuTRe5wwpK6Z6YjkC6Wgx28Bp47Ka7o
fiTnaizaOPop07BNZuMP186tilV1xEMclFu/7WcYiXXgEd9BeIO3VnkWpT4X
Wah/TnjHCrxPiQnfNK8tXuihi8TOaXqXu161+Tsyr8EDZQiOBJLUDhGCjE57
rrJNSiypNnV5RrkI5oXaXKzqnJaWaQFfdWNG6n+H6pRw+PxiVRVCAeDY9udm
QZIpQmp/ivWQHBhr9rqjpNYs8flMUTwNQeYnbh1hYfLDfXgwhr4J/xxJikb0
n04se8ywGaMQlmXUjRgPPJtheuUKgjLI7igFWOpRsGGXRhXZAkRbOxjXoWj8
xAzIsanosj1QNChUb8Xz2fR6IA4vLMtINJwIjxMHqYCu37pTzK4+v6KpKQU+
K1iAHJmWCNMb2pb9J41QlUJu9tqz88WRuHkymqFNm1G/zSAgVIeEoVWSnZOT
7Ey7UXl3aP5ZsREcQOXK/pvMk8rqEp2ntq4iPQBXfaJOzgLg0gG9TuiU/dyT
dDxlw+RE4uhHVOrdHmWnM9EAOGZ4FmY5+fHJfARYD3r41XKybL6UeGE+XaIu
ocIHhxa7KkbJbiYoG35lZ2y3Y9zSWFF38IFLB4jMe+w5oJHXQR9U8GP0cgQr
00IT9Ff1o1vkSce0i2fxNgMoKaz7giI0lZBY1VZIHzLJWzZymycJN8jxpA68
HkwsAlpFnhvXMbQc7JjkiF1HOjI0JYJqWRW5SJ6Cnlt0XgLc929bAMHAnMU5
mExsTkjoQ6+r2Fh5f8BKDH/HyM9WEmjsEOwVZWbBhNpEBJ/11iNGhJLCkBB/
crLfeHBc1Au+QOCgqwsxaqdY71wetgVh5dAobpkqFDgCyx65NuPDUVm13hAw
uDgzh1H6BUiS1Oob1OIHOBLVcbkjhRWNAZq14neLVM/+0NXnuXhhLjJPGhU4
XG4mMSFrMXKT9Qebx2gQBtyi9aE90VcF5LvjY/QlQe6JH+f6GMIXZyNWRZ9q
F9Re365f0WEfqiYTQ+tz+cm11EIOFnjvB8JDFGbe5mmndw3k0n0NoJa5GTAh
bdS3tgDuQSLUD5n6qtbHI7aoXfueIyv8FyXmihzYsakhT2vlftV9LXRKZdjH
Ltmpp4UPJBGXgeJIYzVs4p8nEn0PAdcnz0/BJhq2vcQpQbZXRd/HTORrXT5K
CQBcyIREZsp2y5vMZmcpGUQseMCNEZ3oxRlrEy9dj1M3i6Tt9lMRGXmmKyBY
xtc2M3eofCd8VVNklFgmo+i8rekuK1PZuKHQHeIRQV8GLkOY/EtRoS/i+JxM
LiVirk+6a0jDpKCxBd5vgrjxi2GKwx/C60eRxMqAynnn64s+QVykdumAHXWb
8bLsVkwGpqFesL6sQ9EvDaI/uj2S3SWEF2JMNYRMO2wk5aXMpktyAXl7KSmS
AqvMCLoXB6SL9e/dPbJlsktLeKjjfFyCeB461K0RWNkV/I/rqJp2sBiHXAfM
IBM1qgiV3sl4Sf9jTXTOV8Pq/SEAnbeI3Z6Gp9HYD4xytsBjiR4p3roTIYBf
MvLVfUIPgMJZCo4lWI63J63yROT1VGh3lZ9TSOXPJ0yWlU3txdOOCJF/iEtJ
sJ/78ixwmuPlLm4H0eGofmeGaZAF2PCTQUdqFUPX2Jg2gupISZwN5kkGEwRY
hem7Se8zlaHZmlQ/txmk43MPdHFx7MEsgsvUNkzHcbwmgTRJumnPgDclyfch
PZrtGavQTKOLhg+SNIEZ3I0xw5oKcnM1Z7VlNowR1OBJI3h0P+iuPRWV7enV
sps/81pUcNWRIY7SyS8l47aRsovFAiMFbNuo0fs/rf4mn8H7OGuy7AI5C1c1
YcDng2cnHXoqXb4XoGvhBe3a/3MxA6J4oGuXZsAWo/0KMD5v8fqXt6Zb/2LH
wdbv02SkJdC6feje5RFePoDsjZoOi1176JmSg3SwqDqevFwzaKS8QOs0lJsA
zWDKdwMBXjGv+yt2IDjHbPBXC38MKBgZOOkA2pbG2l7OwsZHo80GkW0HlW2r
/3KDviWNsn4OQzO1CH8ayNgP0rXmo/N4pVIXRbvJT42YizwNqYcZET6PR+6v
BruJVB49TahypHhYImyUAM0ymFoPTnBzRFhFF5S/7bbFcHarR1oEm0cq4IiR
kMrkuCHNHvx3uyjOLP0M4dLKyV4b2lEEh6DlQA3pBKa4fkpni1dIxK3+cho6
jE+/MqOVLL3ibOr60uXWjCvu0e6t8S/IsJ0xbr+21uWZjuqdWj7xVq/crK+G
YMtx4Hra7v4V6k7YRrpuWOl2gT+aqJ/yXQeTeSYfvL7RIzudS4T8q5MT7Tih
QbnQWyQKHcMKHEvxqc1LdqqM46k0wr7fQcJ7D4mQD0hVRwjFeuqDwjYSYwWj
wUT8CUsTDcC10tlMtIJnvw3buYJ4tmiAQbiSqiJG8KgfQp9HuKKOo3+GHCeO
snUP0KBQjfgFwZ5EnLSTimOUxzWPQLjuramNixzdMJHF6gQzQzgMYVQPq3ec
mIK8xVdBVsiUUPk7RSirMLYxxf/cis7qeKIpmVqENav7HceYidBFz536midd
k/MMz3LKARCy//yWO2eVs4/HqMOotCiuQeotfg69QgZNNM/gMBRGscOD88AZ
8/KEpngfs5jDZyCJYtOQkgdypRpSq6XV17mAZGRJqNo0sfe9hNnY9+wSw2os
ZGZu6nkfyLkWOKBzxfuKlI9KWjhEQmtdWZXPXkIvVDcmcxvI82G5ogqqXPHH
0lOEJK9hruDhQTH1PhdZZ6IcFTdKDFftq5kGhsPjvj5FkoZYMbvdH2Wz0P+I
VrV59xf9sPeA/32x4wbQHTi6kMWqZtT/Jf1LB5AZXlCzjbBMvru9X06QJEgX
14T4JEV81g6jW88ZLg9AdlubW2fdEnT/aKEEY0gH03qo28T9By0CJ41ALuUl
qZkKex34UI0kFMENQGlSvZXYM6wAW3fkPK9D9P2Khk4zq66LMplNh13hlTQd
8fDDLn1iHH/KKMMeDyieeqkb0qA1T/wAYMYeB/f+CusN0drpa8K4U4fhz2z9
61ieY2MbDQnpa1m/4KTlQJkOsd+SbuvpUuNULQEzf7uljKrYy+bYYoxNYSsz
q6dm1KmK/2M7CSvWwmon2ZwaDGADalzsaPULe8kQi64Zg1EAX3sPVTKgUiOH
InrS0FquXhnD9vB0+W4IvTYK9+GJw/1fHO3uxZUB2HauE5P4XqdUdWZciy7X
ItXSuLhX7onIt7MS5JcN9bdY6RZQR0ZCckEJqxmERCq0Pnf+aYZsih0EpAsD
hRQb7149zIxsjJkonB6xKiN16Tmb6tRMkdp5qae79CTQkb2Q9EkE/mkWkrVz
atd1xw1BIb+vH8kbyDScA1L+QoBmnARMsjinlDF7+99KDoObt+mrW2Q1ZZZK
Yqj7D4H3mObhUzMBmWTWfWrfArpji+xOyZNxYWPXZ0DGkyqgwUF54g3MuBAi
EjojTiUgxBbpTQ53MX3Oy/PDsJA21sYoDV+PiPhsnD6M1ovm6xZmOK1Pm9GV
ik0aAtyAweu+wOBCeg8Pu4bBNBk37tTjr9Wg0dtsIqm2aEOFzv8dCC4eRV5j
q7mT6N4zCh6MxlUTB/wTCp79mq6cwVeESI2wLanoY3DPJPd0g8ZRPbkk0go/
UXLGI1Jl1i4KEl2Dwdad1ERAFj+OuWj5idxP7o5EbKKGBx7kn4L+xOUSrY8L
WkzW6UwGD6UkYoZcPJidYdKdXEwY4N50PU53x/pqB1nPktNFZ4RQL31Fnuwv
wPH8obyocsdGaEDCCYwyO0VtH1rc5Up/W/PLA7ClWLzEsnJtRFZ/TC16MO1B
DB08B3KjGjlQhaIkdyICWiV8PNbGyDD8Z/BcwWqeSkSUJsDDCGNLcfcyx6PG
TyArOsNjkOhU+wu7bYoKRY3/7vVTnWzZtPhPHGHVtU8JzLtWXbCibLBy9+nr
mFLn4F2r4xlaYuNR5Ikezm3Qg/1r/UEkGv30HlEVU2Q2pKZKbW0PWAMVkvDq
OdXTTcYa64ACKwpsFZnoLph/HD/rxN4dZN7Zle2LNVyHt6YtTg732TzqrwPK
aflAF7qZ/lDqvf5DbV21Yvu8OsGr+03koTtEGKGNHHKwSWDwaut9L58cb5wG
YEgSQVAfbvVF/mwzQPNvLzj58GYHvJLrbfHyZLpiSlESkTLOkTVJqXbfqx80
FdlqUDSV9qQ+Dko1gH7XloIgeyC/IOhxhjvLRYTty4ryAj8/gkGnEDWV+Aub
XrXvTKr4HXOwdmntwsLaZ48pyPU7UA0a1g7kT5X16COKk57Yohup8Ww64hPb
5UpSPp7i+fsT5J3JDrW5KPzWy0IidnYasN9tZSXtCSMlB2l/4yimlXoLiITC
Rm/0f3zdmTObQ+/or9i/eInEDuKsOh2NXnlaZ0m1tXtUbEW5XKoQw4oKVr7A
R9tlgN4DEdhFAokd6JBOXry4UHSBQri1sl3vMvc72LUExcdXDMqis/erdCDU
hnMGj+Y9PSrS7xWHW2/L54HDB92oYTDdG9JKAANjkzIQwi+AqpZozFoOJWaL
rTbzt25a/01qjIdY2B2I5gtdSmjAza5OyoJYLrwPQQXPDLu8MyPxbxNliayI
FqN9p3q8wdpiYfla5M0huSecqV3sotAsENf7WTAys8q4TC8wwNfVrtOB4EkJ
DRswjtIneV6+XvstTuM67IrWzsYKBzr2gxo4JDBMJzq2NRvJuJQRNkcfOXQC
UibSYFxYd/wDTJ+16QXpTEhC1UibPjjQ7faRjyt803Xss2/dic2SHeb2x1uU
uuJDTevaGfn9c0WBiydA9VX3561/h+UyYyyaYVvLlMh8TV6QTzaATZ9YZlmp
A/kOCcbNhLvpJcq9igKN483UhiocWMmX7lFGJkUpE2kw9n8gMzJakkP+BLG4
Oo4JrD7GHuns+ehtEF2cuUi4Cebl3EZbn5tjKsNI0avQi4t94dKyZh7kWEAk
g/SXXos1Y34QNWSShaCE2Hn7A+SFdhnQv4aLBfWssC/je1BnKiAsYugd4IXN
vyz5Lc83Hct8lw6MJrmsoz17z45MgAUPbU4OBSJcxfcns6GR0j+6OnXVuVoB
1hPxg895N3N0PMltpj5rXDPSAr+dqzosZXbgLS3z794Xj3zxmxR1jU0sl0k8
GiV8zCvWtMo9WMFwn5Io0UGer0F8FEENl9gBfjTFj36h2gnDWuivkxQaJAwL
1ehC8CjrjI2x2L4477Rc1UlRFDhhhbwKlSUcCO5/oOkoeXxYILlQ3McBF8cl
dPiIDEK51e4DcYupW51JYv67BiSAhOum9hUOLpZD5LWH1MW+cRftG40Uj0XD
jY+DPYj0Udl3Z9w4/uk7kljxG6rcflZVzc+FeNfUu+5SA2PRsnZniF2dwXCY
Ej6WF9fCtEa/iJLKLJf5lA2tZ0ZB/ORcBarF5hxet6rSUjDRf/Xf+BgPUBtN
HBmrgm6T+YPf1DJyF1gNL5HtM9c38xq/ZeNJoQU/d+xTwJ8m5wBRpaC+cbDr
M+wiiVyKJSlHHEpnDxhjCCEqJjfSsmYa1BsQOz7esj/Z407/jsWGLglPeGGX
dUhEilisY4YNxYHaS7xokI3IjJw+G3+cMWbLkjcPMKtPsT8lRkT4xNUCIWxe
5L9u6bVtS7gKFmuC2dkjsDpie4M82ZWG3BfKxYva1ivSYUHVbtdjb4++kxnT
znW1btTuDXQY57b+NhzkO/6BeLIiIQmuTre1m+g/HVDzU4AHg3OB336Z4t78
97tppzv260QTvUqE4ZqgEA33a9ueqoSxzXWHFhAkFuG+FvoXuRSmFdrLj+8z
xPlNUQM/5xFIILHJf/taWOltSJIsKMGKVRAzW8N5BtqspRT2fsQu1gTYXVt3
3+bez0PQpxlN42ggeCOyvAuKJC20/0JDFR989+p/kYQjqoqJOk1/irgJ4V1t
4jbCNkxK/efNm6Gce0Ywpua+3Uc9Bj0iNEu8ZL/nf3eR8WhonAiiplF+sfdv
2SyvV9Mu/IfJN+wceoSlUFNaBWqueHjkQOukq4QVXzQTdY8RHiPHV3p9uHi5
HA/LUb+Mlv7r9muqREtRs58J92WvsSvpi7eFueMu4k5Or3aw374LHWI1cO8l
77wdwem1UFpkktyBYPGfyq1KETJbjW6616hMEqYplxtBkTt2Ln/KcaJIyEys
jB4aNdeMxLtA3vZEum6XTqiTh3DBziDM8U53jN0wfgDrKyFNr63JaA7H5H24
CerL7FcWpVujU+P9BVnNxC16pGYmGuanB7j4iSmHIyQrV062AeNO5hkEdJ6G
dRZl8bFhB8Wp/8a2ZiI8F7ggX+Uvy4qslR7aaWWa0ROboXvVUlMSz489wotU
NS+E9D//zfI3z9V1l0QUBVtosWvmXQ+h+VZQYtiRDIFLLG+4qYrz0uI6H2lo
v7zvZ+HMvQROhzZovNlxwQSereSUJw5LAtB74uYIsLtFjlmgwX0EQZMgZ/Mg
qa8ejs8XsrbPjkYiejEWwYHJjFR2kbovB6WQkeD/kpkR9JY/880gcpg5qOcO
bLOpulGnw9HmHjJcUzc/AzCUu9xnyCRQ+hbLOLOmt5+czoy//40C0fopfp20
PDudIqaYf1lk68w+ocuC8sS8Y6Kx+rHThc61Bydut9VFOAaWjiiCtVoqkBpa
c87vd2CLKp7QSec0V4X3yP0u0Q2Me0Me5rF0Cd2AkPA9lx7cJoTh2YBumyYd
3Y84u1XpeQWxXHmJyTdZ0++Q+v8RCMKqcG6AAtEp1Adp6cGUfUmtV3bImj+z
j9qa3b324qMINR6CFzHBul/v9A9mPXTsMxeQ4/UcOcq/FqgJl98VBTj7AEv0
8ujjPd0GIUOz2WRbbtANSR76BiNa9mPIP2z588qRMAF0cPmon92+LBy47krZ
vrWepffTvkuuE4/pytdSaLWSiwcAaQcv+wcNqsCbPxApQrEUdMc3YgMOUstf
h7twh+EFMDqrs3id+z5k7O4Dh2lIxNqd/J6Nd6s+VQf7Babv4pXZHVsnjt+G
igku8z8V0RYypnAd3dKXjTI7qSWIxj9IgXlhYn/aoTm6nJKgPnwbpHzs5KZJ
XMUphxkytfyPNHB373DJgsX8EyNpJrjKwsoSbob9XaQ23pN00O5cmy/lx0q1
88qWzELga3D5+7z77cY8kNvvpel5fgYdT+0gbdH5K0CqXiKwUtF1gaRda0At
IsS9grvZD7G1pM4OayNmrwj2y0npfbO+dXVg221n9tOUY4ux78Adb4H6d7Ti
EEanbzU1Nc+vwdb3XOmcKJU/pK7Mc4BAG6/arOnrZmwW/SMkIRFMtnsw6rdR
vEZdGG+L1Oa3j1j1OLXRUq6a3FhbTf+fPwi+YeSyF7ZX9rPn6orBSJe8gzRl
AROCA9odlKwnW4JsYPlxHBUb4+rgwV/EAd+e4wV+HXHnDUs5G/8MRS1/b4IR
LKD8yIS44noh+C1aKiJpxSwaLeQGBop+CIJI50HmtALx8T+vxOj8g7Obot+C
07AYqYBageQdVdTYzKo7XJQfFcxsJWTDnKkXFQgdOVadqPsuAN9TYTlXoSQy
3jPOV8Ocq91nW8eeIJHqCXppHekVOsna51R+hW9+ngRv01hpnaEXXrcV4CaF
oRkeLnVB6fhFbltWKiVBBJXBuRp6DcDAdCbPIPO1wM5a1HGSkjNSg8m7Z5h+
dZ0Yxu+4znxmUdBT7Rgk8QLidRhwiQQUTNUnCUPAWaHQogvQi5wgBKYNYmK/
kwMnwIdMhOsYwUdQb7Yk17sqRmwCyKztWC05pBAziAh6TNj7/3U3Dx4X+WcV
enzG3WU2idVViBRcOYg+TvF5iQ4iOK0zyODvM5xpYS6avJkp5LWWV1YUu/p/
V/S5G/D4YvYhH6JX17ltn4UENX/ZLWp4lux+azkYr2JrkKlK/k8DpjRbGr3W
0Q9JegoJGfF5zCbimpoIWv2pR3MqOb2ZOfGV7w/9l4r9kdwZH05cuk/vxwWV
8TJUe92+3Nr6RpFwLmpko14No5jTKsvJqCJmqbAhGZLM7c0mlSqiUa2EjbtO
J8CWz7GP7mOUD2mVzj+lWp4WUZs+wVSleUC44pDveHZAJvOsoWmGxmLvBKGr
tdqhqhd4AN0LUcztRD9YtvL9vCXSjGx1uXDd8wDwkKCv+e8CkfjvrKg06isV
U17HhoOEY/1NWQ2xzXyoYn1mAJVO9AeBKGPbW5jIMogmWsd8isgHqDZ0oTXU
fEbJxtCjeIytX0lTiTqqmZBwzcsHJJDpuc0LhVquPJXGMyFhr7PPm2e8eAPp
GZkcatjZxCNN85LcAa+I93BB9+FtP8Ev08MN5bq5vsBKcu+GubhEEDLoSSq4
d/NpnxIlUSllKeqaiVIP6YlqAZpAjautmRmxhQYOrW3HPBPc+G1RtdgSREs5
d3/+M86Lv9gMvLPDARELjtrdZf8kMN2JoLdkH4a4u++VLS1oQ5U1nv/wz/CD
GgsLsG4HiilX4iZvtEkAj6d9zmtCXIUV2zoanfod6n+73VFtVli5K5Up87Rc
jFAIbys2Dk80tQ+JL7ccbmfMvjEXO2gnSRs2/P8YpwBjhMp+RoX3QDnA32ed
65bbBAc5mrzNyVdsSi2hw1wplt7swnvZmPz2lCNjcux8M2xL0vWyBQInSBJa
zqxAput1bTD9jKPgd5k5Qb/D1CwnIKPObzqZXrGQiqrI+GzVbNZ+ww+zmcYt
KWAfASzUnZKNa3B2vImLGA5TsKjg3HSi2o2wRA9q8K4ozIgn1BoGMGXtkS+R
0wib4FwyK8Mi1kuFKV/eArZhYLLl4Ax+tNUV4C59g6mCVYkr1MVAzcKDH5Lh
osibqr1zTcTnXitYf4mjMhuMo8M7jSXV89x4DA6rpoxvpgXjm3cbJNJCm1lv
wCIvz1cZhACjVcXu8Hh4exP4P/EHn3Z3D+HRdgesgqGuKeGSk+nFU/lAvLWf
8wovcKgaUOPUOZKRDJhsVIkK1Vgb8DwK5dddtl9woyXu0ESs9JC5eBVhS+D2
YcOgjTyVc1NOnJ+94c7IT6qSK+MdneGsWzJ/i/w/sNq85QwN9uMiFL9LrEGS
kFiO+KjnBe/zBTJQn1u9n/Ww+kUye6cj3qwiB/EvMRm2AhKiw8mCVWsOWSBf
do+KwdVn9zD0qmXBQJ7Bavcsg8EXPEoBtebRJ5XmmXglROmfGN4e+YmKzsuc
+2ilxXZRL2XNh/RYqbAkjQA8KbTRHp5unfKPFLP6Auqm8HEWSLMKISjoAyB5
c9wG40tqCcteeF5M4OjQJ9ztP1MWe8p9q/M21juepf1wX4N2ay1Sf+tINptN
09u6b7Z+fj/O4R8rp0m2v3CcIinqjgkV1Y3IiQRlIpX2FZSnRNBbGiK+rwyz
rL0qDmz6QsAQGAtvEu5zjTMTIBYKvWQ0YLaS3NPzKD6U7x+g1eHvbQyH9j9x
u5rYXo/pLp+n+RmtjURCuMSK+qJO46ospVMY5R7TPYwFXEmncFH8urWOQLpY
6w382xVoKdR64y3bFl+1NBRBlugO26CqmWJoqR9kAsuHOe9K9b1PdPt1masc
jajfVyNxPLnGWipwJt6Y0sCWqIWW37KX2oloxm5vQhn1BOFmTZsXQ2KVjXad
9moKB35cySzE04u1uQsbvXnlkG8UKqttfJVphZrgzmaRVd6EhxJL8gl6eYpw
CCA8iuoFIjgqIIvCKv+38vVTZhr+0fA/cXe8JdR7E/zTjdQ7qWPuIAcGSH4G
W1BdKIWR4bMRA0cdNzbV+fdfe3NYGC2glxhk1R3QVSVbbqKd8orNcBcc6ZCm
edmeOrBg7nxeDyQM+LtD0N4O8xuJ2d7WQeXkNw+o1O7PRxaBUhphzao8Pv4i
MUFIViC/RTEm3+FUvTvxkhtXC1Fiau9GFf8utMrEggoHySbPNBETT4Pnu803
C3n4ux72hW7m37YxLLOhot6fhNR7Crdz1FJUjLZf6VJ887DBBqhUgZVvzcoq
IUoK0SkH07w8PXxbU0280FeU2z7iZf1fiAGj3wWfU6QneAZZm5wX7DNnjn5f
rptDzO/Nqg7qqAcWWBkdXgfQeYFJfNRAOKNLzLm+bBAhNr1mYqwJJ88cYhrP
fwgiDfWFleWxIak/1/EKpVY4E/4nsmT4lJuLNUuSXYzRTme/wKRnkhyclLG4
hgbGZn213FIEF2Qfksvnwpe9/LaLaEFGse/A1EkOkcK+t49ouxEVnvGRM5KO
uUg7X17vouEomZ3Cwf4BshU0o9Xuqk2yAFphkUaHCVIOpFXVRkPvDo+y5eG0
MJpBXMTH0zmqndSu5NNwagJLlFhwkdYl6Pyq7IrJPz9WbSXAU11VxvIrZe9v
r7PSFEAccFLtHiCgTvyFOX6gFoVHLVmzLnyp/qnMYtrmybdezNT7VUglcze1
hdsnirjZpIIO0D4k+e4b2Z6hYID6vDS2s+LngW5g+fdPC51tBhK8uEPwJ7rq
Ga7u/QFISlYN1Pm3+L05NLDcen9SCbfiooTSAsYguODMXqXCpNRPajdAUi47
G2jIwAx8H+Z1BAHiW4YMDLw1OWBe3u4W1WnMVHImVHCGOlkdJTOPOtasnhZf
sHJN+DgqkYr2Eu874hbTjcsU32UHGDXcr0/9gBivZXxapJ2D7MA6UFlvZrs9
ZBBk472vZoPLfK5rxB58PFAwGrNpvkb5ZlwETxrKTXa10/bPKjeH6NSDtj8N
HVFGDIH2hPNo8u2yvua+0fKrCJ6xJ7VK9+9uBkkTso8iHqM4eFy0f2bpUTQH
O84BcKOSUgNcKz4u++gka7gTLR+57um5tQ7euELzHI/ahm7fxQdTWkfLzHyo
xl3TVK4cy1o3YRW30fZaT+kfnX9RSekQ6NXoEs5K/N9yNEXAm4T0vTdGFjID
SMUOjJODQOyGPjHhoJiNcg5KHp5TRuvqsjR3u6+KGlFXNLpCmXDqP/RwKan6
81GFZwI6spJzhiyBEWQ9hOa6xTvITShDUtNaMrm9c7io6YSlRLyD34XFDFgK
36V3wH2IvSNgOP2TAnj1lespcSmEzo2iUgNJV1YaSr0KHLJLeCRs9fBw9+Os
NLwRR3V+HatHyJ7UJNVokqM3/TzpUfEevN2kiJTSnxSIi4dkaemVJTWifZ9y
+p5GGAAFGDlzVfc+b/0nhMhe/qPICynro16jY5lm6Wfc93RJDWx+XxOGqtmV
jT0wIO/kUlFSXYcqBwm0NrIn7c4Eomr9noyZYRO2nWFpeUi/hKOnu//gz4So
jA3qUHa/7NvNIqWIrrHbJbARfAik0jISvGvwZZ+hkmnsLh25h/AYMtyOegFc
fukwGLQ1GkBkqNBhl3bkQ1LvlRpjlE//EvCcFzpaenAr2MW+XflwNVu6q4ge
p3TFFPe29f8qZTY6vHyJopg+WyAladLpgXgrjjh1/MUpKokM0QUi5brKkgwq
fsJqvlcwvcB3pv5Znjeuh/3gRIw2AM3gf4jzVtiTJmAFishCwsqgd9jw9lvZ
7SGZ2df1I1aSEk0+c7mSIAzTmept8Ckz/NuaylWRssDB7PLOGKbOoJ3z1qH0
kdyD6ad2BwzP/PZ0tGuId9E6oWvVj+c9Ehs0vVSmzf6Cbk7YWrPXfqH8dc7X
msKuRldytDizhZ4PSLpYhgZUBHluKPvMrB95ItDogGrPeXYH22IiMDj5B7ap
fJXeHqsunN3Kdv3OBLTcfWCCTnDt9QCmj72KAYOr1M4zC7Mpvip/C6f3AhKI
aKwdLWWCQ5f3tS4hSr77CEspNneiC2oCz3dA5TwsFwYZv1926OvnM2eLiGtR
EfQdUd2Saae/0/cu6LO7vkEUQTPZZlc32YB1ySqMi+5cNVi6ON3ILcTjBjJk
bjlmlAsIKdcj8E5VOwB/x7CTULXHC3Tty/eebUaa3EScAswRBGXb6DbjEvJi
0YrDVRfZbPbyYD6lfvST924e3l2Uzd0BTD0p9v+EnqaOGqr92Haej04sZS2k
nCy8964njcqG3T6EM60tDabtmgH04BVYzsBzSe8bjlM/v1aiLj88K9TkV8Fx
K6kF6fhkA0GStQgG2LKOAU4KoRy4IZ3bDZSjUADKI+ubI6WJNKriLCMDsqTe
qH/krom+0JBe8xl5n1JUsUOks4zB++Aa1yguWsigsaDCjykIHGut6moL+BQO
3xPq82pDI9RLPp5w/VUuzwRh06xPOO89d9xRcztND4i20RSTW2Z3wrr4CpC3
cRiUH7Jqt4Zqz0kQq2l/aBRtObHIB2C8I7D1CxSt31RUDvGTzF63xnL2XAhP
8RJyVutRVeHjPFBcC0hRbRlUF9GyB1Qu/RI1GVZ2keJwyBebNRZV7dA8UdG2
2ioYAk957b2v9VT8SwDu9znLAqOL8rHo7QKdTnYPh/W+uFPaDYbdsRTnicHY
lRdYne375A71tiAcXx/bZjVI+umte+0mlaEhXVAK4fpJJVpH48kQRhV62y8V
SOvURB1nmLczdQNpS6rjL9FIGdDxUyYpGSchvrQmalLc5YBScttVMBSrhArK
eU8HSCG8aR9g+gC8baTOEnVykN66YUFcUeiHL7eS5VOlkz1StkBluFAq/sLd
J29FYcKOGAsxzF02AnT0NcZBC4YMun3Ic2MpIsT3PxE37S7P2lfbreMOsUnI
K3vUWTEi5n4tzWQPxGF7HewCvtkcws6H3ruQfhBWqOpoLLRZ8fBXNJvFsEXL
M1eUiBq8SaOB+leAy+enZrMTW0Oj7uCuJtrcfV4W+gXH5cUn+1aF490QYrrQ
gmBCoI6am5LLP50QIaqyRfZbT5BIoWiLaB7E8uDfvt2LKyNagZ72Cto2FZMa
aY49qnEyRn4ozn7v+kjhMQqMQ+rdzBzskC0ZZVKDbIQqYayQa3k2hIttlpev
ByWWRLgXWQ2DtbRksKGM/qweAqs0RLv0vHJjQ4KsL58mu/HYDkxGpDoGRV0o
IvALv7dqO1R3ewtNFIPIYesXyvICcfAwjMPLvTuETPylk05DCpNCmUnkoxvf
q0lnyQdIk7WR5cMgvwuTc4fq8LxSr/ZDm3TM0TDmtVu9ifsK58Cl4OM3dHqX
2L1B0Q8S0alUpHD3Zf3moqTAUT8HdpCWxF31yIBWiWL1FBues5vSCEKQgonx
YfoWc8recttsvo0y+ob4I04UVmZS7cm4NVTUFtMcw4cLU4SYpuN/qw09U4Qg
6bVUxK8dpWTMTA6mRSt6sZeRkRIpPpDv+6l1giGlPbByMEbgZ4V3kLk4qq/G
0s61MTJRFyrkuB5Y4DHCoDEAbRndUJAQ39YsMgireZaeJKGYtt93S2UFMAzu
UaYmRhXW2sXIwD2TwO+Q00Uz9513/eIp0NkGHz0ynEJapt2M1U0z7BBM/+kS
CAAFp4AwKcW4VaurWktbHf/H3rTivryBB6KLHSNomJDx6RLcgj5h8pVGBGq2
xETi3makhJ15w5RujzhAo+vIaOFlMj8wr4z5D/76YhnqAlx3HVL/TvuChOvK
XTTQY8//i21LPvIadlP6BBI1y8vvHoNfgv72aliqCoOtMRE92WZiHzpIZFj5
VfxgYEre7XGeqs3EY0J4KOdX3kFxpz5ykdJIZPUet+RE6XMZyEOb2alOiVz4
nfzA9C2CJosRbU+ubFwONe9brbHlpsTfMikiWEo6x6NS4GHkW3gShJLe45Eq
qBjuhp9W85lza0ZzT0pGCxKmafofRRGL7DiRZd9ry7CrxHi8ARDVuTTozss3
rZgXveZwnu/ergEqsJZ5RbpvvqNcXlP/OH8AVLQeR8AuDgW7jpkh7i81zo0g
KMnUoOeEVXlkeSgfi+ldpPg9O77aNeyzNlODj0AXMTQrejuS50BZ4VSrFrJA
0pTwnSWa4PlJRbXZKvc5W7MQUjklmJdbz9rbFEPAHCaxIDEqROqaCLWpHVLT
4knMvmrn9xWEU3Xxmtz3yZQ0so8XIrtwfyCp3txXJjqWspSLOq2j40fHWNHo
ZZL/EIu4jy8QZWU0xKe0EP5qPAuIpJctimRepIeSl44ZhkOtcEZudmU/oS76
KhWKK3WYQUvBEgavaTLEKLsy1PEcfP16oJKPrQgPe3ezxMTgzuP3SvgIzz+P
rqAibiNVwtkKiiOIMjx4hTh19nSun4D3LO2hwrnAJkhztaX5Mkotklt7RkHD
7AsIm/a+dNwWBa+fSTHp/AlUEyKJyr94tSrgaPjPG6CHdXejzXdnvScquc1h
3dMjI3kTHoSV6wotrXUbbrwMan98LeY8jZ/a13EHAkEODIJZlDgTucbWsx/p
QTuJzIIe1yuYUK/m0ir3Wf8wqZLjmqNODAa+JPmWpqZhF+qKMQx9CfGn9NbY
Um9VUy0uuCmKYMgkrnrne+XrZ98/axXIvz6WP9hPzyBa8LsJYDcZHmw350Av
yfs0JfXj4Ajg/DnSAn1LuiUmeU1eYHkPXf/OzYLYAzevoef+QgsiDvHZ2RhF
ggO38kR+bcv+a/hmrx1wyuObmlrdAxGXeBrK8IO4Y1VFRG/xiKG2V80pyQJ0
Mv6Y39cHKp+vLEW7OorbdchzYXP7JKOmvqkRk3Tst6w/QhUpKtrGDNZNeGoJ
kbkK7NjRMGqkF7NE0zJpdwH1qB/FshDzrk6zLLhapAIQsTZD/zUEwbAdtK8A
vMAhVMQdmkdq/R1am2I9yBRMOLwuXCuyylDEdNwOcdv/YN/GX1Ejvh162sV1
BCzUPRRl2qZp7crq5kF3EbX6tup/QeKr9ahTMJsPm5k8L5yho6VQRUF2Nyq+
Q7ErPnqK0LzFnB7dukHd8Kb3GgNQlZAYQ856oZpxuTIPm8kz+IuSLQ8rUUoj
9+0EyLdFvKkUqLol61PqUp3UEB2PQdXC+/jL1W+Uz7nnTSq/fqm1eawV5tT+
gsZ+xNj+IbGIWZPWfTyXtYbfryZpmsRiY5LUnGfmJNr7ieZSCRigDRQ5ldC5
xV/cpjoje/vPBj9jv3bzC6zcvipY4I4SijUqKySZbVdw/1grQRVI1BWxAZiK
Ms1o0FPJFE+noYhSG3lvemTSSNFaqOIWQfp62HcHRGGwXAz5gEECyW/A9IUV
sbJcSMhgnN55rhH4bEKsoMAEggA72SxlE71WeqiRqbCaszVMJkHeLxO0vhCR
JxkU57E5mtDb0vmwVfrrFj04mRqbm3POu/7PMg5134OiGqvPePtm1Iswc58Z
DjDqB6wgS65TLeQtxLJzpRnrB80mgwwHHVCxb1K2XCyxJtutMOfOxK9MTzaX
K4c+//4UbI1rntjst0S0pAkjo8P26bErxUP3gDjTMwEuWE7kpL1oIpTv2ZFL
NRXGpN8i1XtAL77M+9wy4qIj9fioJx5qo1DGbyGAQNzU+mYuvNhbjHy69Ykp
li81jmKSjvIkoJ8iUaD4feKYyfwZd1u/3r7tG6EerqoH1Gnv+eJ7xca5vkBO
+nGFccgcqosEcgSPvu4fO4mSbX5X1rT/IZRguqnnS/HACBDt3EqADHGe+Wnc
6gMd+6T5oc9MXLVHzjfHGzlEtVpPC6esCGvhUBvuqQBz5dV9wwIqPqNMe0zP
8hjyCOQaHYwhauNJNrP2kkbaZYW5at8SkIpSzxJZALIhq/sMTn5xb2JAJPcT
JPmYrCoNiMydY1V8X8j/cM2OcA3Ez4tYmoFFiu2DZb2d8CiJZjPfQ1QaMpW2
UhQoJdJS+MaWkV05pVscBu3dLk/3/EPk8opptbXXj9TvqL3OogPRvxmVWVSq
XWKtey9CuPaOSROP9s0vmsLPJfFnvhY6aTz3vjaAcCjr6S49DJN+CkK19+Xi
+x429tLju/W0S32L8+NK95cWxGLzR5YEURkXlZ0+MrwPXqTXoP97jgArnFJD
k2w+eH4V9YbEii9izGo1we/uM60li5Emi4NL9VUNljPhOT99wmp5fkGVXhgY
hEX2rB/4ObeYRA/DIDPmahR1aNFCvWt2KZMdGfmeN2mJntz8g4PDb9B2eQlX
NGanTnC6lwKpbQFinsDarkz8ERub3zXMaz51Gi9+lc4OnE1/LB5Hq2pOMdnj
Z59c8ZNHgH4ymXXhLf+xzOdYrPnz1PuEa9d3EaWhjmmDiVYKxqj0kirShhZv
tK26wsTn1eXpEOvnmH42yIknC3u2Je69e+ND0XdeRyOazK2d2VC9HiMhrgc7
FQKCp9vruzcVCGcSaJQAjmBtWWdr04k4/RyJB96rdzVW3cEYL1ih/TN3XGp+
+yQ1APqF1SDnhdOtCdkJD0qVW6gBAM0GhF5CXkgBhjSM1AyA0mQphYhw85wI
aJJtfqmI9Dg6sDchOfJ0EJG8bEM2YU7b0dJl/6FDQ3nof7+scSH65LZpp80Z
OW5Jperaof1KDHzC3R7hbFMXzuve8HlQQibma/SbuT+Gikrt8+mtdTX2gM7P
6hJAia1e5bhKTov70iP/17fEqwCIYq+7P0Mf9e+pWNzOgjQhq34gXuLUwQZq
KqJVQB3Bg4Da3tPY/yKMf+cks21uXX7TCQ94DReHd2r6wYTy+pxsSd/21JiM
++vefV5+0bKJO1UMCBy5+4BcpUr/idwTe5haLaLPETssE/RNmKM337Xg411Z
mtZzxDyWD6ddaWDF/2zBGof7BM/vgum5Ka9C/CU24gD23nujExgzLHbp9+/I
qu8lhQtOn6ZLCfqrkGULNgVt9bPb75yRRLRrpplwRHS/eIG0BAXCEgFQzNzx
xyk83Bil9kJdL0cCa6iB314qvAjrYvd4afDvNtmET5mzwwkPLkYATA7GCNeA
WhvnzJeZ5IDkX0gk5tke7w/vea7x6znQNyBiIEPFIjCr8Un0ZUSO/SBpRel9
dZq2LKeaWa5bufBzleisY5Gr2tV1m7/sjuUwHdVhfEpTMwm73MJVhxqyznqx
3P9P2uZp3n2q7USYkylVJCzOgfM2PeRSzQoUMQnIG2Y+bpsLSMMB32DwTOKb
lE0+klkm49j0BPdMTGAix8E4Rjj/nEjoADfWd7M9Hk5pg7+EDcN4pWS2EuEK
Hhc13tbVgaoKj8RpRPeI2SCNMiXJQT3nyD9LqgAJJ5YA0+E+pJu6XSKnijQt
cCt8EHAPWASJj22BxoK0GGSTcmEDODFQ38J1O9cTNZ8X8qH3G9NCU/djR9LA
Jb0n9aSQAdwdZnEKFZIiowYoUTmVJRfNM7TDwbC/Vxce3NX+nLp4tGUUzVDk
75FwYx90suXYpReJwlTNDuGragrW3U9grGyoOsnG7kybo3MHpts7+Of5Rkbe
jVPONvMJIzg331jv0IMzh74PMgK/O+eqI1XhNntTKIHS4fpebC/Cxku2UQ20
1lwidyCCGk2V4KS6uQ8eRWAbM6rmOIqlo2WZMQEfSDUb7nvUIRMa1j+p8rWx
D16XQbqfR6Ok5Oftftc9kSW80o676BNLqpM4e+za+ZtjqQpTv6KQRrzZT1OE
f384zz+rsh0Qf6aZPkpxF3Zfrms+2IU+UKdbVlJsjz7qjplBoX2IaxEPCBHW
dbhT5tAfo2g1pybz2xC/IgTbVWFDtmdXs+7cdy/ZfORfvGt7zcyRzuTTEvFF
veDCkIWU942DBM6lkkAP8YKTv89w1/rMTZAkSTUfetml0XOC1YByIJDL+lDP
1rEBi6dxCkmskH8Pxah5BQTCy4qqkO4p33DFOFt2BoROQnq8eYD7mGrZ4R7p
+YfXOwyYAUOiAHoDbx3C5X6oIhW2gw24SDouZphx0dt5CxqjgP2TKLzFwt4w
Vsu3GzNHNQjr+JKUA7DkcC3DsM86NNRCKy0Ks0Iyop2NL6LsoB7tihJxKhdO
CwUve1kFTTfwfPru+Zkho8cuzRmSK8avznVlmpMoBpwsMdYCn7JxRUHbkdGL
HqWnonJZD9nuB8i0zHWZHEtv9Hi2oHnBE/fdxsARUsff8rzmFQQz1usZmDpr
oyS2S2YPxKjSx2y2yug+3PxCnLX5z4oCcBgZxbHGi89SFU0ms1kzVth2vtQF
cbMBQRP58JJfr3aYBDaFycAiFlmnzEftqVteTYZkxzCp9LZQ9aYybDIXbmWU
EuNEAi06K+C2a0l1UvfbI7uAa9aJDK3yV5pxj1gepkCYbN0ZCRG4XyDJQmeO
CE64Q/ElKiWB7tWM873OoZgUmTh95QISPX3L4jOvhCBUu16OzyH7WBro9/Gr
xH0Fr6xaAN1+CbWQmsLqGEfWdgXc7OpF/7ZesoWwANw6elO65uGTTjmNHvzR
0A6SjH5UT6l90z3nMcwEApFMVlB3o1y82/8AlXwHeyk5UhEFTCEM66UnXCZl
hB3KK/qsdjLbono8r9a9IBCsKvOAspMT1DX32q3VI/h61Ia2Ujs1/XZKUyKB
I6KRU3iBWIY+tIXYYrlD0Aa9XJ3mcXEpI+gH0W2MUTahhK0Cbq2WCGtlwemf
CBozrEpbZ+DVvoAPKoNQ6TeJaPf5srpgu9TNH9M+NsjSxTXi2bGj5NL4ULKx
o80f9IyjeAbzZAQy33i0/L4nKur3xkg7NuLgbrNzMKWo9tzRB4h7TekcyXkU
Ru0agZqrCsgHffVMNIaDk9Lz9s7fFt9e8ticc32eyNwFRxMcobrm+q/hm1Jd
oCWWArRENYr9H5Qi02lIyanR7mk+oTBjTViBIFvXhW8WuI5TqyuKbfdEnVY4
o9IvRXCOaKTBpMD4MSEqyTStprbCLo7BHzIhURlXA1OkVY97OxU0RPJFglAJ
ZBVmmAkW8kivKopVE8P205jWbBjKU/mxSdwy+7DC5Ocw2aoN4O/RT1HST56c
NIlKhF6+DP1p9n0IPSyxMPcq6VmAcF6E4Wayq7031ThaGC8x+9h0GcrBsRDt
mrK0nyOkwc7bSJWZ3zkn2d8TqzzTZmaeULL/FGixNpggFbxSXU5rUbMbPhNa
ITBQnxHnPav/YR3dbNNlQk1FoH5hnnz0bSeUaVZGek7DIKJ6fJeuYcREqhg9
lIQLOELN4ZX1Y6YjcZ9RnzwBYuTcaqxsp5LatmtO4bh0OfTBAbk2HQ8Na28X
IqTBshv5kUJCiZKMbfGja0nj1al5PTybNzqtgkAqTt5sEAXi35wtq69/5GFo
+XxYkuD8opkY+QrS4WFOiL1xvcMiWIE09MOMkRrHzjKGDH+O/2JMveC3umQ2
mhTV/x1CfcCVcfnXdIIW/3ndQBG8CcNJXC01ArGQOQfLX6FBmH4tgFLWhmNE
O6Qg4CX2yT46NXv5v1gOJPc71Q9GyB/pLStVtLHOflOsQZkoht2rNWgm+KsG
sxqkiSOVg8+9VISqqHJfJ4ss7v9+nAVe0BssjPNqPVvSbjYaqZ/GLMi+bTdU
sD/kF5V5f0ze9krlDArBOu+OpoOPc3wDvm3N9wF6p6J2RaFZ7j7FMa72B6Al
acS6AMysUGpBeKjsQxR04/OtkLfpINN2Vs7fR9gGxvyjBnKFuNRk5++1yJ/r
9rXTHsq+Qfz4AUINkAFqNaJL98WWSb9QGI7K9OGDvv6n4qVMCdZAEwC2FtS+
uHuEhkxxB3OMGHGnoajNftGs+QuN8Z/30x7+/QJHISWl70tbMUH1ergs/UpC
iNzNJG1q6frzWHb73BvxP5IB/4P5htRgeD/3taLYTKyhYhZUh17uvql8ZtGe
jxvyb4xIAENfEMGbEus40vhM13VV29vFEqQLu5Uu8qFfk9U0+qPny6NFzgek
hxN6z1sUGxUmdefv9yG0iDsbCVLmKin0ZMXVhjpsuvq+1NDnncWXMF4YdHxa
omZALUoWYChktDg9QUV2wq3Vt7c6mcX8K63yZp/vxsovLJFQt7Qztv/3gIty
0dHzDtEdG2i2ZxfX4LWEJm8rTwJzIgjn7cdY40xZEIPGBVxzfDuQlq1Fon4c
BlHuYBEHSq5LRJlEjfhixoeLYVc6ktwuj6aFcqi5IbSBIIn3+WncLa/8oi6m
fiBPqYHPwM5XHdTsWwAoC5+VQhKHrUDx/nbTt1Q3A7ZjG7fHs29wXOInxjEM
3i3LI5o0kE1FQnPJOTyKQjrL/4APEHXTpFZDprmau8nYn165Snl/ErX5yD06
Y5GecQ+qcrlH9dVmy9K4dZeDFM6wRRP9PSGkC9cgDYpJY6+31sol8zsgnaeX
DsXKs652ljkJSif+M1+C5nPOiPlWNIQ9v52RvycEPZe93SfRBNsFQO+Hs8/1
mWN5lV8tbhBK1Wao5cPBTaceXJLUPTCNzUG+tcvPc1pp9YbiunmWHw1XyCg8
IT/KeZ5lGMFHq9O3OVtH7CCSPMJJX3NhAabK+awQHPQIdSi20sidmRV4kREC
LbJ2BrLuNblz1EdJo2lZCF9zgPit+dpgLV8YmIgAPA4sH08KUaO+26lhCcNZ
rOOnPHLCaltUa/5FqfjLk+pSJ+1cc5VLP+znTMKPf6Sxnn2PLUkE3gjHU0TO
soa64jzPiHS9pzul5+v2cGd7KHMTXzlroLUw1V54E3cNxyYLN13TMnMtDeYx
EeGQW2qRzVXjibZtBvOvtcAOd6MBtkuSCWgmNV+dFjI0QnPSZ94W4lKMI6x6
i+/ST+D9gqWwV4l59lcP1LBJKWqc/7943Nm7dHNYNHzqUI5VcEE2UYg2BW8l
AlciTTBeBx0N5OG15hd9Ijw2oP+oyr9vaSLxK367IEOs1maoMFCTyeReod1i
/woeZspgw4zbPWVVrHwCkmGoQiJuKj693BUUUeBVewkd1T6M/IWNnbqUlbvW
rWyBO+smTL1tmSd2cuh8szkPVzLs9df6picTzm6DbkRQuYC2kqO7o486IzK1
AhPr2S+OKpN5S5BWsx/5hV/vqLT6fp54DKHK6eX7iEQRbJiN338tqhmlYHne
ajQ7dKlllYOG3FhHWnI8O0h0CfeQKSCpfUQfq46DGqIvBrhxuOaLIvY5qZw4
81L6Xy1d3lh0ZXFQT9wlmuO7XQM0tDOymzrNfitX/BXSr6Kol0UUW1z4mH3D
MlXTquOVmYmmm7NJPQRZ/aCfogk2S6T/9C4hslfxuzDRmBzoTRKctGJpKpBV
+Ncw8dJP1rQR4Hxd4N4EpnF5OBGSgnFZb70sc33iHtnQjdtxsNqseKHnBp2M
YmhjkXKQPUClg2MA6PLRTavtNCNAUx915Cz96aISsasCPxEOb9YKj2SJeMaj
6RT/jtmsyEvRqO+6ye/CNaTrtuoaMRc4uiRqqyUR967xK6cp2i4bKfBDN/5T
IGegqzIiZuB4yrx1b8z5T07CYCzfbFJIic+o+C1xRpERXmaMDgcjXSLroxhX
R3A5C99FUEXTwo/NaCS144TnhmZxlvaxYNdsqvD3/fuLSH2AWNiBY9VAte6G
k+4o0LPJjOaTGG+1PWzzJPDVhWtKDjbSspNi90nEz29MJ7xxrGBeETGJ+tHQ
DmM52xNn1PnEpOjzt8u0GuEB8Z2Z0ypyRCLQSb71O/rnf0m3xSXG5nYPuU5p
UnECFWb8B5NKPUcDlM8g7BYfWnh1SFcVTLc2aNnlv9x965+kJ/9yVqeihGYW
WoNAhw5NbIW4tEstzgqswLNJOTT5MC6QkZGXZ7vfgVpIdVDAnfMaV7bdojK6
CbEA/KQw4+5OFwyagl3wrdlB9kJu+V3es5mFReIFSnrtV1A6vpvkLc7rXyc6
PiDGuMYQuRyzk87EQS1rR3L2W0hmm6GzLzYtet+M8IgQNPFT2nvgHFtDP+Lv
q7biEy+S7JvBRZ+DcvHwrg12V2xI61sx4NRryvSC7qfoGCBgorap8KM5KavC
vL/lMuQ4aFEjHnqEKPJOuMFhMKsmiQMyU6pLmpR84PuQFzyinNVlzFrVN689
Y4FHmxAj02buuG7LGWL5kKavxwR+hrPbAD6/N99cfjDp7gWR6a4KAyVJWRUs
VCDZwJ9IuPIKaaJctReUJ/8pcM7tr0zOMeiF5R1jwQAyvVPYY/A0ecT25KmR
jxugLxJkBk0wlecEAjg0KD68a7pv3DdvA5zoR9IhYIeC9lorWczCN/QSml8j
+aJG3nCHOgbK8Hs2PkAwiYQq2WTyRhd28P/f+loNKd/+dlCxgwPUCfooMI8j
ZkaOSCp+Qpw4njRwJbC1TEAn9zW3YKytZqGftq4RZWzADiqrr17ufO7a0hHZ
vY7hQEnqKDdoBG4k6tpTcEPA5YfT3kr0FyLqlVPgSCvE25sVWy0A5CsFdA9A
9WhBEWYmjx0e0HfaaB/K9AVpkN4ZUNue5Ozba0r5h5l6uRFri1gmXFnc1t3+
KSuRm7CEnKKKw+qyO+tXZC0IAOzXbS5Nn+UjB7ZmMU82P3o18TIRx/HhhhgM
VSy4IUrkuWs7VMZNLUk2YlCbLPD4lCVHt+QKGAYLiNo6KNAW/uFT12D11V8i
Xkyq/FTaURph0AxE3opMxyionDpr0dwd7BxHzm7+L1HFiBV0rh0J5Ki+HyMO
BeV8zl+qKUdLFR50rBPM9u55TKwx9UEdceBUipu+THCtVwC3/92SA4dInzoU
XS49nXO+Dqn8j1+M7UBkhygPxqMFsaGU4dcxlnDYfJEDeXl9SYLh161969os
cSxwp9/nA5OhyGE0R+iJhjtgRz5XBXOKkerDwFiwvMBp5TDf1UemwEakKGRM
yX/4/VUJq4lnsHtazNzUYpfQdkp++NB+9reHUC8khF+2p9stDjuQ4AkdQi0x
FPbtwseMCA9vzOU3kYTu8hjrteSVc5k/prpRaMrh3luFHt/Q+YBVOeRq8Aw7
7UAO8Prak509lJtry/1Pu17DaxJFFqW93Mom+SfCOiX27xW5vQnpe5+rKDyx
lyhD3VjsQJUZ392ONa+xwwyGFNSg44lRHW8KV0oupQhg6Eq2X0oEYAggVFOe
ImgN4LUV3L9dpczvi0qwaV2pVzuus14vG1TzYn5GimrK/lelIajhA8o3Ne4p
D0HlVebrXcuP7E0ADyhw93bEnmnZIEnISBeDQLzrDKVNDdMQJDdN1L/p9TEE
BUnVErerMUVbWENbc3YQ/kLarcApcrgCeMlhCCUHVAt/KewMCz6kSrPb2Zf8
Jd+MJTrSLgJuJmu+Tm+YAJlnR776t/pBmaDZI2cjljYK7rDyE9QNqZ8Ji4av
EJiJbFVxFg+n4vhm7yDRuSUClv2kbunFsoAHYZUcAUubj8GuPzd5iUjjKfXv
ed2CTVNQJFwTnPUEpQpljXp3DvaQN3hAPNUbFDqVfY5PJ8aWnMC1i77lEzJq
/76aetQqXL3GowB0wvcqjhkhJxWygtJR2u9LSMsvRUY1Aga4Xu2tyZV8gbUv
6G0Gg7Y2hh9o0TwZS5Yl74mDRmu8XUH5iMsNC8uSkLhv1lLS+hpJxwU7+1ET
EzRbwMioj6tCfEPeXH1rUbdZ0C+023t7AYOtu3+G/fx1CEoKO6vGAq/AwtLB
yRySJqDrRjNIxZ+Gh9Xd685H7azT8gSaSJeiADQSsXITIDiFFwV2MEfmZaf7
0fakEQKPZiGQbhVx330dNRTLIkHvC+1QzRcxloIVzlcVZ4i/yNZ6wg/ctKFB
PIplXxG3NacTwHT1HFi4k/opxMy5KhKcxDHIkvikLeXFze8wb0qAhP+fE/Hv
Q34xDM8sqlZy/ZoW4usu4gOIA27jOGSEOgUoVUQ7wjvg3lGXFqneSqE7X0rI
sw9NXw2ED9y+EGouX6aMs8zipNdHNfAauAJOqR+qEveCJEy4IObgBeDtYSjR
OLzH+FGpF08BCNTld+V0JXZekLORIpO/uYK1E20BgXlwi8NkCanmpMsfcdje
9yjk86NGced+s3xiqOEloYteZ5iPyW/rzKCexc5hbdsb4pIaIAOxXiA6uHj1
OhZtUD6v+tPaU3dab0zz9NbamsZzCPj6VQFJN5i3qERqkL+TxkNXIr3RfNnO
eIQSK7m7Nb2dbtI6JRdthDiInZBLauI99gSZ5PNSKjbXFvoly3jk6gaxN+qI
KIFPBnOaJac+NxSsuneNjAO8jbDxIsObKJyY4qKA9ljw+uCEhipDoy9txVbm
qwW+PCkNbEQTbbhhCv8Hy95+hn4vpZE0WGUKA+UGVJVultZZf51VcqVdVOpc
kqpAfJPLYUnWOHazeFkV4TS7JPWmVKdZo4J4kIeXklcbfxHOXUR0oIsBf/3H
FGP/+d6XXdLlnHlaXABqA0VD3LAmh5+SEcXQlvJ6MbrryZi8TbeHcH998Js6
NSG/FqIWicZT9VOFyyD6VWO+A25NdjcTC0yF9CL83CXSWnF5ZPIe1x3sxshh
Grn40e6GPwLTnlaiEmClK2E9udP24DrAY0qc2+e5mnVwzxACa2m1au21Tn1y
plz3UfBEZ+hC4cTH6umQCb0vVxMkYfplSpYlv6169SAgQzKnrqqJeHcieSOJ
/MRwDOf7tC3rHFQqxwjG5tSrYOjD4e/cEIHW1FjKpkybg9tB90ujPynimWyr
p31PHmL5CHTp+SD2HlMkYxbY1vaDzoPIXadJ02xq0h0zUFWx7UyMkz2U2tpx
XeeI2K6XJsaLqZontt5XQMstThOwC0uwpWbRCR1YMbB7XWnPYFjbJr7lzVVb
EHHnisUus/F0YDeuJJRSFmQfFgriwuQ6lfj5JcInL6e5pROSZGm0cDgVwxcC
NSB5qkgmGDiMyK+MaleyWqat5JFNqDrKTJe+meU7ZJ0a0kvxninZTysFJWct
uSWPKLbUCd2fWDxjPtEm207tah8PzpNDz0U0XecJROC9LGVdNwwo/l9OTL2L
MWzRNW/xaFwZk5z4AjeF5ywhbrUwbVd3grx0XUYZicpEY+POA3nOswR9iGhl
TOZu6F9EJwCQ4w1WJahimUlsBKduCWbe01RY5SQYwRNQ7XIENqamZtx2JjEE
FDf7jQy7zBaHhOF8P2Bk+90qbpjNJnDmNE1tOPmQLSQML1cddWVCjKDhzCAO
NaDEPLlYLvyel32Ye9U+FdbNYg+L5hit8Zbu/H2MgW+93cox4ANSFDPfNJgF
2uiiEbEJrD3frWpN/KUWDAzcf1D02JfCnpVGWPRqR4cpD6fjR/RhGYU5hdlt
4qQ9G6LaCL0LGAe+VcTS+A/ZfWtZzeVr4RFBZo05s27I606G4jxl9h77ZxEp
aneb5ClHTXj+rLBNeg7tdL8HAJEPhnZQsayEyPCsHM4gFB+X3YEHOJ2BBF/v
0VCQ7T6DScBh2/3vRXCGIkbd/c/xgBuEsyJv9LSVaD7GWSAoTFLXNXKzrs91
Y8gs5HvBPkc5SCuv51Y5NIM0KTTnWJZShYJQyIfRaiktFDoHszLITziQurU/
3gHAz3mjY4rkTewl09C10jVmY51D3s6utL8NOYegtSE4S+o6eHcuLBqHvBKN
/soR0z7GUcjZ9gCwaZ3hBzzzXQcGIrRyTH3Dnrl+vEsm6C79yaB3z78Rmen1
GdX9XizliP4cu8PgazgpGom4MW3saT0whXn8HCoQrw7/4PpazGUIOu1jJJJC
a2r6wyU3tVZ5kppXO63nJY2x/lYZVqG9OETl02UkZCh4c2cXQhcZKSbmu7pm
igbbusUhUk11EL16AbdD64eX7qJsU2V1YjJFm6wnh/Ze3uGenSbmes2Mzbnb
jX3QzgE19gUnDyfx6khJCdJJ9RfcOKm24zUBLdy7txxisqD2Af5ZQTxxLwi1
a6pKUTzRfXaSOJ5lMDja3lAlwfWm8fSr6JLshk425YDaEX/6EQVPB9R5r9g5
5eljGrZojX3PcxMbKOflIU0+5OgONUwsdggK/lHoZ/hejS1/HqFOMScftsBb
rmv+ikmkOCayxlk9J/youUZtMqwCFbIJKSKHCLswMXl7KYHyK2pnXeFNn4S3
5wGMzvoCJodx73UKqF3gtq51o6A7aoZnQzizHVwo2jWdaF9uftr/BGaBHaS5
C/9bc5Hm2fuC7SqGsXfwPtiI9YN5m3zYA4A39ua/F2mqtuaOmS5gmZxXmYLR
Zy1LT/4nMZBumOotKJ2AxWfRBO1gxJAgmQ+9ZVdtCb44VpN4Zxrp4r2QWJOt
V/QCjHiDStOHU21BGlLO7O8Bp60VIgYyg4ehs8ShFGzdUFXTtu04mcRNEn2A
V0YPPn2d7gamo5h1yoHqOGQe4NHNO+hZUYQ2NGP0HKTW/1x9ue8td+oc6+co
Qjtg0OWXRdS17zDBpu3sL+35CIiOE/u9oyarHGbqTcptqFkk/QYgxIwAzTs/
6UyHHbOXnQ5HvuuS10WjPdy3mfAKE2lLFC5eEBK1Ql3VVEeIPHuGQKQtS+EH
/yfaudMT9JUYVIAhUVdZHkrodzoh1mVku+nEJR7EU/ETVpKsR0NyhQCtYZ03
M+yzY3QwRsD7JnSnodRxpVG/drM09ZhHINetQKFRNlHVFuRir5PxL0XQXIAy
nq+GpnQyE71ND5/ymjtF7P0pSd6Q8W1fUjNPhQklXFj/LVtIoAIfNKaPaT2q
8X88LWNKZ5sWnSDbE55uMa1y9M8OSDuf2ei2lIKxNAloF09ds3V/V2wUD06B
iURHZHQcTEBjGY+AQ2AaRkF0ru7D0St1hg0FYUwCXSoWHCTUVlRo5TgUNqEH
4igcag+f2MYcsDZ0UJ0kQh2hGglnpyw3xCLoQKiTct6eX1JcnI6ho6ThnuJz
5ZgFyLvqhtnnnNMJ94Rsz5O4rCzcxd7NBXdhvOOj9ppNcZmSOoKnCSp4pDND
4qZASorXO1baNOZIb48AMa5/1u8Ixjr91Fr9g8gCwUZuwShVsig017otwsu2
fuYErNupsCkfO9Rxv9vWr4F8u/lIGvECFvRFSC+MTk0vGJMGn2SVRg3V/oz+
Z3SSx+X9/lHnO0uOxvfLN5QhbbMPuTmuEVIw1wtXGtX8oBR+MhSRp2hr/nKp
Uea1pLJBTfT2JX0MqxvXYYrnsmzp3mUCA7hCJFwRItI5flsJG+CIxy+GCJ0d
JhgnTEJMKH+qZhpS6NeLAWllNl6CCNSWjvHpSTRy4P/u1FMZjuffl3EjuYAx
FNl3Ds4rOjlofr4cjy+a14RTm+MtpkSn4gBATw3sWSw12IurJnPzeUVa6R14
h0W+79mqv9hlgikLUGdRBRs7A5sea7g47qswz1q5E5obBQ+HMAbbZpwKZoqM
13vtVRSCAZy7J0Xnc8vqvv0DthDY1VoSL219T9zHxEJDo3ypmUFXqG/wHqbN
xCybpRop9ABdG0bIjQ0R+NrZ7gQqEoFZ88P4JbRxLlF0AziTsnsCMz2DM9Lt
qNStEg5ltfDKeufDFT3PnRXXKSaTFtvZ5uBL690c+anJHErfy/OsEZWkL+NV
PzHfZP87e2a7awbpvh8b7aG7vqHblYE3wMJueEFm+nZDds0TypOac/zfBowz
kpfqmbawAlzPqXC2LlRPt9kb6fo08Mzb8RipwwLV4vh7RUfKnZsWK3YNvgI6
RdwMCXL22X93y0L8S9NuOwIEhb7ULmroPGGb7W1q4dGykq44UIr/IRVyNEyJ
q6Ew38UaNg4NAX6f9hCVhK46BQefgEDd79n9fm+AXXrp12Hi5sr5SWoXpqiV
MNYYOxC3W8chhY2htuEspq90ArwdbT6BnPvq/kjDN977sy3dlkJqOsseq5cg
8n/GMbbpjhsqRRqUuJSP/BdKX+kcxtskSPPFYQztVZJmd5RRgET+EjVcoTJR
uPzhx7HUvmo66Okc27RO7eDh89Rf4d4xIftKJHSlkwqGiL8l7zw6uMle/EQg
SX3hG0fC5pMfMNLals9YfLtqlHLvuGaZZ9mm5Ksd1aMT8ivm4eOaBaDLRXv3
CARVW44fx2/ytKCxIJwLiB15IaSjGd0w7AO8hGJ9uFnIP+J9CWlz3T77SGls
c/Stf1+rPgrBuBNpprr7bOPNRzWyUP48jbdTjXe3gQ95PrKh6dQKOjW+W39F
UJG5GBTEOn2Onw4WppnNIo2w9G3ASV944W/bJVbdLgzmmLzdv68QBiTjwvaW
1z1qBcJ+dZxeX1E4UEpXsRTlZ2WEq4tThoiDtlIja1a2tcBQC3vmUMrM3uXV
QoR+uOHiOy9ATQwlr4T6WhtYH9nbY5X8cTHStNYDkPp3B+a85zYtziWmkl/s
ntFKSebayk8VtGB+Na2pJtUanPzr9+fA2N3mmcQg9xZTbmDT8kxUz91wFzQh
ts3MvMEXyWUkYCh60j4SUjU7tQR4HwYN4gsOGcInVnHRWihTr8o2RTTgJBzn
1NVA1OdRPzDPI07lgG82w/50cM7r3QSwtNKBikvMhaw9T8DuAG/iwYnNpcwW
iOpiI/ep6XCOYvbu5q3XUqRtEvt8XwnBpS/9rL/udM7Y1FR9HicVGzrk4bzo
+MuXiOv6QVevwlcpP6duo7TYJ+CeG6omNL388RUJJLabkiXaO8UH2ggmWJrP
0q6TxS35Zl0IOtLdvLd5dL8vgPV5YX0HQLhdf9UGstH0pFHsLffNbPn6g+vf
GWv9c1mhx5pVCMG0EVAJx9LuTt+wYGgMEZyZKAKSx1Ba7YIjs8FzdCsB6R/C
xPOQWciGS/8k0pghfzG1d0TORWeyj/bQ57r2LIlDEjhwX3Zbhber0IjbHn89
Ll1n5CbyfPi/qFyjgngGhC+DGqnh83BPbv+kNafIa5oG0Pq1tiz6urv0yuW9
SFMgy/M02QeENg42E7U1e5KSZY5EqeO5d2YoTgnLJ2hWSOsZzniLqLL42eGj
SYYH4W6ILOUoyi+W2B7qzbQEfEZdUREBiAsOVspXbvAolshqQuOBnNBc2VML
evOizYCL4gNBz4uNE8OybZinQCet6uawTfxN5KV1ZSL7tYstwIsmhTgQqxkL
k6Kqxer6Qxs8/2LRVrd27VtjGNszTr0u2zMR4WnrXLTAyhkPXTchGb4XoWl3
BaqysOji6Uquy8BZM/ViF106NR8L5uazgqHj2MMYOJ0XChKXeaj+61jQZCPe
sjv2BSSGmMFHkEOUmjbIJH0GDUCOuWXEr6JBK20bPClOqR3gvrymNVA0yrac
vO5gvS71662/yyAdr3PiPjuU/NRdan0rS/E9bahtiBBHOOZQdfgWsr6Qz4l5
MSji4bB6O1cT6216qRfNfaulP1IPYIOAxJsbm2077GYaR9hWTU5uUoTQwuNZ
WmNcstuPJXNGfzGOAJkVJt6t6rjan+gdG/XKWjSPYgMq2g8uBe+klHOJpAmy
VcS48iciAldO+MODz/PiB9hyzIlO9G0gi4zxoNTvHuUgmsfw99828VAZKlRI
VAp8aHQeG5dnufK1dqD6VTKiZvSvONvC2jEZP48XAzBur6LXnGSiiWOsc8fK
TI/5KrcHycUAZjwAzLr476avqcdMqR70ToXMORdLzmmE18mgVJ9Ob7ZMex0s
l38BPR5c7ROqxZWzuYDTqHIzGcka3Xxqaev996rJGXLh1eiBhHESH2l3oobG
MHHuWTb9MSJ5OUrq3oN48uweDb+B4EeqreWJ1slAIeTvFqFqbxnaWfBI/1kj
qc+7z8jTfJ3GMjOmrzO7fJBi7n0XlRv6wyZ+iZ/7ZVC8TGruplZkEvNnWWYz
eQ5b/69VwvDkB7I749SXo68XPw9IPO0oMWeYEVeVOD6VZOaXyLI5owEeejcF
deNiPcD5dT6ei1kP+mULPA6EdZRuPdk0heT0V4ydcoc+ZmYW9npNN5wEGLsj
4HrkI8C68Gm8R8veAuyrTxts/j/PXNPBS4pTdkyFYzwnBeTQuPTRTXoREvL5
K5ktCME/OOhmAok7GMCt1xXbK1e7ihkkGc2SFi1TizXKl0X65+sCSyp3XR8e
y0cBx//79X3Re/6nXtrDKhhfyT4hjjhrGniMnNiCHOM1EndaeGCI45t8apNW
ygSAScIbUcy4IWVVXIs1p7W9AJFmr73wCVu5uMl0KybLBXJI4azXMx118guV
OnNQaJzn33grGk+1TlksrgLYy/8WynonA/FKB7X444VAHVEsOfBvxSqsksOz
c4RezDloQuSokVHfo9+/CW250DP/sfNOMGf4wdPaAdsTg7DmR6lfefy+v/v9
d7ZH2RFSZcULeZD5JqNZDUfabznWPaKypWClBWC3g9aOSvcCvoQoKsU+TrjL
Cx7JmbL05o+HIyQoYNpsHIto6+UhRAs0N2nHAOc+pb91m5kkGA3k6YYlyGzY
WxKeMd6NxkNpnn+xfsui5VfRNZbey5P/uO7JiKzeyTOFTCnmGGPqVjc5sJWO
3onJXSCdKue3iPnoFYHNbdduy2K/EYG+LqResMZF7TLq91pzuwriV7pU1g7c
l4uTrS9J06rZz6FVx0tDIJSjcQCBghGSskoHPmphCrPsnRhzSplH2c5SzNwZ
INRtbcDqpGtpNzPXNkjH3SkRhfQyteUeIG8MmH6VVaV6vFLH2z0dNSTWKHdz
vlSy7Hqn926/B0f7xMva6wBJTSrEgJlW1ZxhikbFlha15OIo4+ztyNEFNWxP
Nz0soraLTtYnNA+P8avFiSNtIsStmYBkPMtZL1Gt9XNmHs7+YtTO00G51vxw
XuHasusFlBe00AmOvqVPahLdJWZj+tfj7QtJ2lqy5MLxDk7DxM/H4jj+PgJX
i7kNQdftiszjpBQhvlYWAAbqcJuKaKLh0/3ycFhnL5rHOFvDlMIHuVFqCQ2O
pL4Hh3e7vs0ZJ2NW0H5pPQZazM6zG2uQoW+QL4/UE1X4JyaluY9lEaxrFDlM
UVTuSKJt+KL6kOADvw8bJrE5lG0bTK8X3QVxBGI9qI1JEDXEuPJ2mKMl1Xtn
gKlrSVNmVGSTC9n7o5qd+DWSAlzYrWPPfzZ4JQORGv40pq2cHslPBC3ftAOH
ODHf8l6d9Lj8Bh5DznVY8UTZ6WR6JU2j/3y9iu/qiGOnroQSvcqeHoEEcXaB
hbulmOQ8TsMuTI2SYxPFBCahRiQ88YkpNoL+7/2bShkPQlmMbB8gwnD2m3VI
HHrZaey0ONm3A0KVZm4GXyJ6fm6KkNMs5RXkohCvycers7YpliF7HSVTheXh
Uh08MycbhywqZAv/Bx0KHoWCeqjGhmklGK/Lel1J9jckOIuEpjjxGypzCeEL
eI8+7hlAfI/P/EuqVQoUYHL0/mGYf+RPNxPrM0sdAKx9He61gfZ7qntr2XOk
hiwkSRx8zDIjgrh+f2X/NGfJicqnWgyIVSCc66aG1r78aeqEkwqukWXu7W8E
pq8At0mVCQLEqHlhkxEGWPpomGd8c/Z4n6Zi4ER/ElwLyGsmlan/6Lzym/SK
Kvk9UspXb9rdwoOzFRJjlM5JxOe9hOjhKMGfqFcFgLICE6MPAigLx0QCueDl
vaaoe+Lq7yis0BaUf7/5wYAC98fIrHIfu+0gjuMtO2vSvGH3MZeP0vVuAhX1
2i6gy5LCsap1Isjd+lo/8e9VYG76Y6pZUCTtwoey1OZpcnhHIxY00Y33xF71
IFuGgaBpk4bHLBJzthkUTVSDxIp8nDQiUA6O5npkISALJa1LqHVi32iDuDc/
y/NLM8oBPhwEdNkI2PUgeKRpl51ZRmwgizJSsZWyIJjD9M/NsxPJ4QfLvuXO
PsYO77e94lMmn36HXblr097vlV6016APvAbp7zTyyc9O9ngNOg+BOTob6FcZ
PJXTz+zZHf7SWIVlzl3vcvVlVeJ9NZw3tVKzFDuiHxvRYSfHPr+CTh9/OfjK
FSypxXglH7ljCCTKpaV7gzDsALD3hvrEEOhjsNA16KpGoE6hJefclSYMu+tk
YCsc2maJKDiDS3GpaPJNp7kijipkr5tsmsGCwEOyllKNzC90pcARNs+sgkVb
noXTTmei/OOYli5Jcd/FMJ3MH4pKGUEdwogGmLCmB3ppptvXJvh3/es/HLNM
q5jXAWQoDt+ZqVf/yGVZpz5HJOwFzqx34fFZWWM1l4mBz4ygi/9Ovh/Gxo0N
JSnrk+66S138WUesuXmMG7Ht2IF5yO4g4p5u2QEcvL0miIZG2DqSDzAbqbyi
FpizwsygmfAj475xbM7EC9Zy3xdkKJ3Mzc5BAgUFuEec1yZ1TTLgBVYL6rkh
6AZCgv6b2EpBqiL6i9sAeQhsG64l9Gw/Yy0PbIZ9qcNXChSHhaYlf2XLk+MU
5CRtuRgZABv6tG8X8yo43v8zn1qdZDEnrxFRnLw2eN00NvuTLE9lVWiB05/+
tWzlrF2RLiNvtA7EeL7om7NQoeic5WjK5O2Sp9TliHayy8PGC6Dyaf+Vjsyz
PYUYSOch3syQ1pyLGSrUiVCsu2L/nte2EvGOcJw9mJwcViC8KPov1CkTjj6T
rCosMeQhNoC9d7m5cnSUIpuZC6xr29hJ8zY1bTkAd4QjMf7Gz2KEF4cZetkI
j6/vxoPVj/mOP9Z4ydKwq/3hMRMgPgU8NvYNe+qXbMbUkxZU2Fl62UeOPNlz
DF2rLouj2bstiUS9n2OJwBNg9MtVPTpH5zqnCfFlb3KU1ZXOZkHvh00s0vKB
jPTjo/WCT/byT2qjYzDIHzLl4mx15lgQoSOgcRJo+4A8QaoCxI8kZyk3yAF+
R4WCxroOTjLKgc8VyEpjsX/+OvQvOFTwkbewNjRQXMCsGEyCVq1egmZebje4
Ewpgfi4BNuICHAMmUYGnVI8EJTGODmYWpExaaVa7ssYRJa+W0Vp9fUp4HGlw
SEM+J6GjUNj2thUC09Ls/IvVv8pyF7rarZ7P6DFRpxlPJSKH5abO9adDK1ZA
eRi5daR91rUqT3XDfcsh6kV1Y1tu+jNsb5w340+gRYh1K0nqRrLZtiWZ0QwU
dC2VJK93K4BnD3F9Lt4uf3j7gv69IlSx9IPf/KhXLMg9IWkxEqEvw11NW4Bn
bJ9sXKRJXe04Hc+9bQneuYYfhyPBKOy3YF16Tj/ql9gmeVm3pJnZew1+0ouP
3rlE3L47J+Awfc6w4py9OqOYYivhNcqa81GIIBc744HQCtBPwUiIuGPy1yZ2
GrUgvZEGYczXzeZJHwa9taCcD0c1ga5Ty3wEhQIQa4tzOBBewXrNQsXGTuqA
nnvPJWu18OSMdFCW74occOjKsuR38Unv+GD+baJbyt6HmJzGR7YdntPPaEY0
YlAWi/GaRSH1auZuSaucPK6aFyzoB/tgfALQfVwqv6oZLr8/GFPmKWc7YTXI
uh5gbPNjYvm7JzBJwOlSeJh/dAKpT9pFRMTAD6jb6AyCdJTRKd4AuNuYh5Ti
BpguTItthNS0GfVa73Oemj1g1lyxc/JwuLTA2vqEqOMJp1oYdFjNPL6CwmPi
CxmsZGwf5iEaJPAyHlCrR/hW4O/ngtBmYOftkuhr6aOkgufNVxZNqIyYbs1r
ugBfw7GFRadEK4J73LLNvJg6TqJKF77mNr3o7amoDtchgO3NmWIu9+lJLfmO
5MpAq/vx8S9UfYl48Ej5R0c67PUDfdHaCzgvpDvwFTxbn2CU/Lg9InoWqIWE
soUSKaQ/i5le0tR2r0bfRkzEwxHRXN7RQKxwzrKzaLW1+Q6363L6w3vaBmKa
Y/6in7mZiCnd0b5aOF+JRY5+7zVNDLP7G81HUl5U+IL9q2QVXKmq1wxwDHf1
zl91M1hwg1dwbj+TIpmHQy6rcow=

`pragma protect end_protected
