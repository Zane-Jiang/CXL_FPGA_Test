// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
aXKoGRohhXFZFcWRccEUn9nQmsgY/gWYLaCUCj66q+Lt9mHggwCdn+nELyW5BKEBYUkQTL8yfrA6
Lec21WcXZz8YYQ3VOGpAjikguZoS2ujW9LUVA+bo+b0iue/K6XoBvOVvBBiexfL3JRIY8FsN0Y2x
DCFcfDPIFGKZEkKZ68yb9mdfBB5D1QELi/hpOgY1Y3/dnHR3OCo7iZZguqX3voKQU+kVdOJNvgnS
ZvKAj3Bpsr2cES5uBp2tDVQQVtpbU5tSkaF5/3bvFQs+hOpy5hFbTuwjIwRkyWuQEFFIA8A6sHsf
GRKiQQqD+nQWRvxJv84HD7nnUpjt9hoL5dO5Zg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
HMhvXVFEjEEfO3SRbebFW6+JDGPtsYzliV59msAIRl0qp0lP3OCB9QGgOdMDDAcfsMlcn8Cj8a82
8SzogCUmKSqqiNtjK8SpaKCvQMTBdo7Npnm9eUvhrVrRCeMMD0GkIlD7aN4jRGU+P/wOfAMnS1uA
tGIsdlI1nHQkrV7QTJC9MSGxg5p63ODhOSrC5ksjV0wC7OtbGlP8sHK28bPPb9Ds0kpUJc00GU9d
uceWy8NgbCa+vMW/9WPA6nu66LawMPLkFaN7BU3hhhTW34hII2aULXa36/uEeu2MPSw2lO7gDej2
wfivaI4AItjZpYbhC7/n9DopLmGLDIC1z/3ySUkzFfuF21JFx6tMdBHiNw4tDIF2Z0SLwR0f45f/
TnSYtLheQnQ9AoPU03yjCva78aMwJTSTF2ZmBuifmNfBsVksASthKInz6sjkeRtdr+LxOt3aYWvx
QYVQEAzKGVuCl2uOsNeVVjH/xnq3wIwB3l7dtZkrlfZbtPGgNtGC3s6MR5FWkF3Q4go/yFoL2MEM
m/IE+vpsemS6yHYY5vyAnD9QmlXduTw4MC58BOqvMaz18FV84J1bJBNBi3dx2JxCnpIGOAGGv3Wi
H8hhzkQRsGEM2R4Yo0C61RquWJv35oub4GyKoxdN0EhBPJacr6gmioM4gCo3csHvkfA089RIdK3k
tDgsZI6g3NWM25/bblWX2kefq5k3lzMmVzimWS0PgcghNTCdlxxEJNEo0apfoWAIxhGz+a5Uo2e7
G5Nk1VYZNiQa3s2F2XDOTl8rr3n7VqIhqaV56BYzTodBE0zpuU4qHMR+UHRfx1LcPndUVz1+jVzY
L/1hMLK27aqRMET+9E7GOoFwVL8WhWYigEBepy9z97ply+k+UPtm3LLGElM38k7BDOF240PBy0C7
ipUUS5Ak5ybP+pIvBZUOEBIavY64i4IHVlAiZRAJfYQXIquHNxKtxbAPijxwlCK8Z0kbrlsIKZBO
dzwW2w3caxjiblIHJopyHHMYyxWIhzBVKgltD/GHj01CjSpcT70z175AbmOKNI8UplqrfrDzRc06
sUb+NIiW3toKkOgMvi/csyVa1ChVHx0grA0NpUWIjjL/xvcJuXdkFDIyTf9ad3mPcI93GPVUxeSt
RFoMRCTDJQ+LNk3bUHaAtg9LB+xhPui3U7YDoTG4O3fenGKp9/1kTfDrneSVFYIXXC42eNRq3gGg
wBOhGcJvXHe0LMU3uehCI7tSjcszHn7f7GnoANd4Aj4XNC/XHUaibeGXSBOGE5S17gWp/g2Z3Z6+
cMOt8UyeamMu5kNkycgoeFDFF7HS0fbgeGD20khkhcY5fXCUwKLF1BDZb7PWHO4WGlyg4eU34dBR
Fzcy36Lh2siJeMwmSil6JkewmD9W8jTXjCvL1NOv8lUv2mS+yCETseAigiWm7aBNt2fmJ4FNzpE9
gJJocf+h6fx2pmxNv+zJMrmBQiJkEMlskC/8mTdg3WTmV454RDp1issKYVQG8o9QbTtEiV05P3vv
298dq3iIXDCGSALclADWRBS8YneJN1l+ZNkMNO7EzRH5jSLh4KMHMLS/pekPK0DK2S2Iyis1mB7U
+FbsXjbolhfhKs8b+k+1JSvOkRQE8StSeyPZTcYIYvn2CHajZULGafsO8VGMqVJ5z20EnIz6JRLa
3FY9Vik9BsA6S/yjiYL0xEU/wr0q4vPYf/yhkQ1F6Lb3fMaoqgOqnwYLNeG0Udiqp4nxc1mnEhh/
9sBaeU2HkFybETZT6a/spE/pWZqw+TWjMHlC7CrZT3TazdxIwtnQfXwUIKkhnqfliJG6FUCbqzGi
hTPJdl3phwsb46tRi11ecZ6NN0i5qFRf5jFBD0DhuBNxVI+Htz1dnQPtGoETjp/ikhKjgXtcYAk6
cOs5+zYxFRHkmY8WiqqlMbovXROGNAHpcjY0cdjvTeqgfCvy0D7Mhf8imGhMeY4zmbAh99JAq0Gg
p2vrgCVWY0kv5rpwlUD1Eohs2V6X6LTmjZmPpks42k/ZYrPpxcfMByzq4/ElpXTZIY5DCpj0bLPn
6V6EPKenq+iEl49DQIFTRaIPaY3iy0KF1Y+v963aqRhJ9pk8MHKxeVusCHXvAr/t3gYbKUSCRKu8
cBDIe5ALxhU6Dvuhm6CmfijF248kjfvsAfgLi8WrEvhh6R5PAaMF+UiOpPnaHDi5GwOjLDzpFXcy
4FRnrZ+oHaD0bsWFB2S9LrdwOxhqvPDvEZxrHCG6f4k/KDxAHmKn2d0rJNhj6/98tVSuTcYuRw9f
Fo14W+GmmHxI21mM/j1oqOA9mzMIWHhg2J3LNovV5GNxmY7HGqBJdUAzhtuBPFnXc7vF1+vNMzLA
xSlroKHqs2np9B8OlNX9a3Qtb7prvi/A+2/AifIYJ7qiFh96t8B6O9cU78Rz+5RM0bJarc0D0mPC
VDKRRWAS0XbSO71tW/36P00z92Ye72doTL1wPrQ13HjNiK5iLN0qmQ4D8WA8HWS8MIPKIJ9y+Ujz
EtYg78oDICvlgZWDlD3FMengN2ti84YEnNGkPj5d/KBBw7PkvailV39ClQBgD+b14o6auxNFNxnz
2mDDjvtPDWuSAR/mbe2ICRfMnT8vPDEEyK3n1RfQMIejixm2uqNnyJ3h7yiyMYhJCOsHno3122up
qpXj4NHRGaIdID3LiySo8voCOUVPUU+aJAMp3gUne/fhWNcDFd/ezfLcLdalJkcIFUDDZRcx8JU0
Hh1moAbdwP20+WtaGcnMbXKX6uyfXO+EqNswD69eOHKXIrDIw2dLBcLMBzep2P80iY7BYyjToLhX
l1yfdWv0wQsVNZSB+ZFUd+4gtJE01uuUjxK5iGB9gyzZ4pth6O00sv+ngmM+dqDK85XsfKW6Bw0y
ObAzOZHcrAx0o9/iiDTLiWzo+iSk385OU4R/axY6ERw89JqfDKHZacRcTEl4j0dxFJtON2pZXZec
PtVISXI7xdy9W3CFmqoG1LwH63kfE9nt9cG0dQ8zPULuUGAmICEX6fswe3/Nly+NuMYOTXJ/ZcnB
L0Fu6XKBuXe5kbo8chpur5lzpS3WzeGLxHY6scy+s/5wcN7DHL5b/zPvMDba4Tfw1G7pJcnL+fkH
Yn4e1YET4bPJtcS7GW/UVp0wWNYCCjLrcM2JQ1E60f2YzQMqcqImsaB9MvI5FjomGtecFyJwmY8A
8tXVZjkx+ZxULY0C6/g2exIbDrb6ln869vmr2wJDXdlMCCn3FEdSGCvPbMnkggwGoOYSRBu3MrAb
IIXogpVbx0TNY18iTWJeV2T92wAxvME46otHT890ASfI0cxhfShR4DN9AlrpNRdAqS0VkNdcgGkt
b90+Ou360e7RwYAA7d+H47oAl96/mPWB+0zJgFfiTn0NcfJFAfW+neGIg6knNQhE6Z3PNJ1AB8Ty
NNdObre5t6OO3cFbFcmrsHc4iz55hBek2NctPDiNn3fLkGhVjZb1qbbv8wyAFwUaiNXsj8xrk/o8
mLYp3tkiOsoQQfXoFlV1XYogUxxJVcSOcyZvJETShLBW8L0g8ClvLJxXhu8nxHSBX+0mYwRY6Buz
+W/RscG4yDgfll4IZjC7/V05s0bfFlznu/m1bTtfJvHgwoDTh/MHSlnw3lAxIZ68YsPaShtE4YMp
N/tcuAw74nhQNQoNjwGdyRRSi1gq1LkokvTZooa0oZep2+BVyyKG8NKlA/83+7nm2eZUifMtFbSp
Q/QmAg11B0RJqC4yMdxS7lmbLggDNFEXytG0qaKyqgFi0gTcVmOU1uRQBBaUKUY4nBbEUMvz6JId
fwolN9viRvUUdK7WrLpi4vL6kJB/yQBO079l5FMvDIe+xDvVYUrmr0YKx9GwGZGnq9JFVwkwJNKp
tUsJIpXf98u9mmOjG4StaGDRcDL3ht9wTEamRsK/wZQ58Z/losyLLgOWTcA2c5sxM3GaHCjseRHO
QvNtDvbncYoseC7s+F6zixTGjbvrxhociZjDJbzMgiq4maMiDCPfsB7dEEFEyzpqcwbyCLGlfGaz
ciOgjRn/tf540T00G4o8sd2IzUREc4K89NFJ+3xQcc1x1gnRVZyfXZpkP1Nl0UkjNWRQWnXqWmGM
Y8DudAUkK6me1yalpQCe9fIT5k5WZKUKhO1nj8xq1UvZDtZctPM3IGzSj2gWq27W7mc5EFCgYp9h
1eOtYMEn/2H3VAYfSYepbDZUGeTDkbr8oRBTwojDylgxCizd8F0DOzdjRVyFKerbViSHNGz5I+zy
0gmMPMhRn0bCXbP5M0e8PZmo7eVXBsiIjFbt3ovSY4XF6pfv3AHzpe3aTrK9R/zU/PoY5N2IM/IA
B/CiuvXyW+jNx3v0R69t3YDt7YxTMn+mjFkK/TU3fWECUptBdltpN/EYIzmzlheRYvdQl7vytdTa
Huq0olzCa1/pMsH2zEbl8X3p97Am5Om6HxBNzHx3AqpiLe3W8QXDhHoAEm35zRgohrS8pytPsInG
X7XYyAitv18LvWuuUIBr9YFKR+onueUEYR7KxruQoEnQ66Ppl4HS6ABjbMMHg/eerq1XHHDih1TC
ufePQJAD+kwer7G1WX69Vv7KadsQZcelkx/5UwsJpbSo257GEgpxmdpKcZo/cV/jCYjdbCWcm+0b
uyRFAcNONSnQ+VUXq4/7mYzipZC70ky7ilZnmGaADEFu6rX5EhkgM+zipNkij+SHdnZbL9/Qx6XE
C7EPg+U+N4MHXgc9Lwb92sEqOHfe+UXKfStxzkK/dZkZLDv3xpa6PRm5K+oVALX7BMkdsZTkXIj5
9O9cfhTdbqfmnlsNLgFisJ38jSkPtfM5dPssaBTaOL//gUpxN2ocjG54PlyRouZn7eh1SFxSV2i3
CE+0RKGsTz4CoPzdfoPKGt+6yPnq91FnhjavBEDp6/MbtisrtNTnrg98p6uZt+KCa3TibYdCTNBs
vENPRMvj1zWffxzyxIbhPWDcq5FyhT8Bl87XYuAYAedtkaCxWIdZXwFK9JVog8d5KGlMnKILCu++
6I/k+voix0Sh8qA2vemtUSyi7YAcffyim0xi6osxZnI10FVqz1JbVbDIrfYz8AA3oPXHR1V8GGRv
UArh0GVuDd/B2sK/pFZ57mb0LYUi39MpAzO4Pkc71sl7WppdJRqYMD65kCxXQdE25R7smkZK+3PT
VKQ//yUwCyh/FKxUDnx/u+B21DxqDMKKhvfSVw9S/bCWiqKqReICY1PMe43bbB46+ofqI8yFbO3F
ncLcRk0/feNor32/lnAbWHXUZMm0LkLry3CICJ6D3pXpeT8bXCUsqVHrvAtMSZg4ThlmVIid+tLQ
Tmey6zvkBwaCm7V75fWuO8q3xIq6+qMq5OwlyfUiGYEenK1yWwgQNzlYcGVIKpTQyYv9YXxBtzSQ
ImZOLneYKGUJGLQzwcWbpDpOhb3Bvs81Cm3e8S3+yIx9iCyKcIQSugoelf83HUbJq/NrhjXjTCR6
Qf1gZerwwrRjFspdcu6v6oFyNwoyrU+iQtPkLDbIFhIYtY0HpyO9NXTEIUSBIEaXNeU6tqw4rX5h
RT4slsGawfkKuVt9Yz+RaiKOztAsinRL1pzdIkT1AHeYYzkrFTiTINT6hh2emW5E80dD4FCRi/Oe
ZbbQTKPCCzZ4AQ+rhKgKZ2vFRh7FoJ1XQg42FRTUBn9sr20lxda9Z2Ac3b/Ev7Xh5UL0LbHGOTGq
zIz8l91+ChLM/zT4kRup1tBMY2nU7xNf0cRp2nFHnaCG+Snog7F+nwyK/b1hTXkvCBz3t01gqEsz
JWjciK5eB+vdGGfVYQ+YdU/n9uDHPJ+aSTtqX+6lClf9aDRXHl/M7rnePIYnlW7ebtMuEhby4VeC
Yn+1R4tPOVNZviwbLJN+cw0dUubct2wfqD4q0b57yStBSeJqxk933VWFZO8ZU7+APhr6x7GEP3BI
EXMAlC7FsC7KnV2u9Qy3GcBixBuGXJSSraAnnKxsW+wXkGdGF67YgJIjwbMaQwv7FdWCh9d634wu
UXZ/gyZM12ZM5IwHgzeSsRW1DBUJcxXpJGqsvwX/K0+O4uXITjDmmTPsYzuJNZk3XvoSpjhjCVdg
Ol2VeA7VuI/YR/ME7isBPRuqFijwYD3FOPfheWb54xq+cPeMKky0tg8CUEhio6TTMANkRzl74+7S
EJg0ahta3UlyudWqX/1yr4QiIkBHOFd9iN6BVYHgO/AH7hRERRegyz4x6ktmVZushtNwKTYWhBYR
68YfIxmAo378l1LW/qticKN9Qb8VuKX9viRzcTwqm8lwLFaO6xeisT7Y5FcM1ynVY4fRvqh2U4Ke
0a8xuGUrt5Ar6dG6WCJPzRmq2p8tUz322Ig561dHGV9Bpy0hcvDQphkQMKkeSypiwGxZLHWFOpYR
pzWoKt9r9D8JNWHRNagmLGHxXtcWnP3Y/8oJEDnjgBzn75QEivFePxFwYnsXZfA649GWFIPHBNRm
68jbsPEO16lf1/zHVggb3YKAKFtHGGVPJQqGqHRYfH4G729A/s12gD8fV+QwhLpNimlCYcFXt04D
x26W3QZdtbMZAPy4EaOsvwdgTaVyfxNG9x7CGBLcsljJIrpjy8ErKpjyH9twmG7iPn5eARjobYNv
zWknIHa5TfqhGroXEsAIhOc9UY6rfJC4KRrbcLhflXiXYqz66TbdWtKKPUsRyauIXVN5mlZJzXdH
a0xcFjGql7GQeGOnNyEWq5enCeKBzg6IUiEBbMHnD438ETMhSEEjF3sW7zW68MF1he7yaTXrAFAv
a8KzJiOQHeLYrBf3u0EU1Ilobisw8wrfQOtmc4BmrWNk2of5y69FaSIPpUljJQDivsx4ofYbGZvW
JXhyJquM+/6ot0UI9060AbI+ePEwMc0NBoUZpC0ZXGj7XdVsG6HIWIR4clWfFShserj4KyCczJFA
KlzkcLpcDlWP8mMrFerQ4nlRkh5CCXl6sjMkRuWL1nxT82m9jCJ5E3i2hKYnN2nvnaeO3ZOxPBnu
/3OZCi0HMl+j27z0RVJj5LCntVCHah4Eo4zxB9kivK7ORva1h1cgcfD85joF4wah9BMAaDXF+BgY
0qF59NFSieFWuLZVkb5I2xdv+oi9jKJedrfgLusMKfxwXnvBDUmiw86y5Pa4CHYypAQDwFq8JBVf
UisD5BeQ0PrbcrsCDNxcGa8RFu6x0+CCHlib3k+h9RJkFFaVwuliYLYjmC7LmYuRlQFacVGHWJwN
hjBCpq5hfIBADIw0XoE+RnoFL6nxrqIgpnO5c0OGd/pUyo/CoSueIEjmlqkrdgosiaMBAAXRAPDY
rvOUQqBiTCFp1juUxApKQTKzHZHuw+9poJnWIJdCBSZ0GZxKzK9NRRer+CvcJeeRt9tgvw8eDJJZ
lkeNtVobf6Cw0xeu6fuorA7k6OJHmAf/ArefgByMUynAnvx/N0urhjDhh96SSd0EF3cU+wluwBZz
KQAAsAUs98wixuL4uqJYfrRY0Gh0n4Eq44fkZDBvZcbZbxSroBGgSQBfolMy+T5gapq9kg/3Jqem
/YOPhOzAfr+otkwNiOvZ6yBvjAWZ1Bby24xPzYzTAmpW/bsxsbz0QO2BjhYSzd4jBUEn6JJjQR3w
ujHut4rPRUQuaU+iKHnzpVtJJC4bIc0OpdSzMLrV/RR3ZsDeJhRVv+SD6pCBkQTgSTWs9eRLVCX3
2bLZy6NDWtWTedLWkVO9DL3amqn2wmV2reYnu14nlskxbjc/zV0dYXbL0ad6y5XIetPchaQKLkFT
I5DuzggWnMdOr3w4S4unQt3I2gKkaaulMyRTLqBvNRkX5+ZOGTLRWz9+8leoY6p2mTlBgwj8g3uh
/d87B9o5eCSFwrtcvtENwJ+bBaxPqRnKPkqWW/l4hQZEL1wZSeBxnwE1ir5kDdWAiSjjOBaTCGLw
CUheZ1KQgEV5B54j8xXALdsYLbWaAlJtDrOEBVC4dGOkJWGl0d1v1mZkF9Ed6wdK1yb94aSZAmqR
5qltARUMtBQCx5Jadnwv5WG9Icknp7JqBLpXq8pBq7eD0sE5634P394qEKOljbucXxY08qDUDuze
HOHXoZ8G+u0nwS1Axm2+zNCMuHesqyDhw7Ov1C+6BJsQ2hsJOwrIgwsiqQQRQAMueQebL6WMdrBa
MFO8i0YNLhOaBBjEgIlLZ9ptkD0d8c9GV7TzaZTWa7lik0oQr6wDLeU9XoQ22HszVCTsWLJVvI/u
FkxYNMF0doevGF5E7wOfcYYZZrZvI6ijCWz+WtcuLOY3YH1w9y4JvYJMmpEm7szEAMWUE/9jGS5D
bvcUtDYwb0xJp38zAKzxtJ/EiBmosmEysRALoICC0Fap9JiYpbxoXcd0qVRS16xaXTHcZZ5muT1m
YZfF1fN06q7m8xrphRIPqfN4lAkzoCe7u5SLBrvl60DnI1Y33/WUYDN4/yy5g8IpMTFeAG6E8Y3f
GMS0ZM+jnSxqyTC15C8VuqpioQzQVi3wMxTSdKSuXdUaVBZZApy8hq+1m4rNKJXVO2XrQfGM5qL6
3XIbx7Kyi73EjgEk3ppr71Pv+cQ65M9eNm4Dc2v9UT9yVML2v6b5eEi4dSEVhz6YasF2rR9tstGz
2977rnm5IIh3boPqosfHzvTvx0Z/OR99xDXLYQHOXC5kVJMe/cp/ZqihFAQDgA6ulBfp89yV+v0l
Td+kGUrnQ7EAwRmvfeKuhf6b1ieJEAParUyQpVRiy/+mCV+uPxw/FbiHRq8NVgqUf9Wwej7A7NHf
kyMXXLORmki11omgAny+bwJGVYvrdz+0tngY3PWfIm3vVp7MohxjW5duVAClIyssmzeQfigILMbI
HvLHkHSIiYpzK8WzNy8JMDqkZBG5crBGR+Ra8vhX9BCtTGR16/Z3OUAR3R4DNy59CbRcovvBf3mn
fl/fMPpvZeiy3RoWbWXkrSrSW3kTCI3wQqSAETOd9TEMYXfV3RKRVAIT6q4QpT54m5EtvV9S3GZr
qPWGnGr86fUrLvxv7EyhNccXvAMxxzSQuMVAyOOmZDSFIHdCyyDBwChf2lGy6GO3J5Ky+4jgOXne
vnQ5y9poF68rMaLKOUARheLdY0n/TsaKcENnsPpN5xf52nIVOR+nh9CLzCN/o90JAbPEgt7lrZIO
MnBI2oyqX+IlQoTCh4k1XZJ4dIg5iCZiGLBi/9TWDTTy86xg5drNto8A1xHEBOKtqu+hq5S1OhD4
RWuaaewCBEChm9g1sZvDPixJywk6RDVzpdzbOEpiGSRwmZw9C+0KllOE3kJKnnG2ZKnv9WDZaqdd
h1fZ3WIAdeJ3O3X1Y873v+E+PmkbcR33dYH6Ry3ud6B84HyoUCMdQpQGJn4wL2epVIPD6xpCyg+o
AAcCPoVCeDVWVDPWMTJt6CFqk5ZCOZmj9EM2ygSaviwkIPbLJkbRJ/DYtkqxu8bvL12Xp1YJTQx3
AOu9meUDvdxoqghewbemnVG34Kld1yEruML4ugwxoVwIreKTruMXvPYyaSBEnZRuEGNAqEU6HLr1
o4u+iN8xIjuBOZcZ2gtFOl1SjgP8KftDe8ojmTVVobC+X3d5BuYS+OftfbSCxtrR2PWDs01DNMG2
HVTZ0k8465pUJ8MzZh+rKrxZB136u4XP6AiAOux0E4niI/htqt7mqtLHQ5KvhQakoBohUAEC8B55
sBkuyMM8WwbkLGZ4yzXhIsF25wNuklBT61R30TYmUGzyljVoCExVWHyavVXnz0CBdyVRvuSLsbKF
tFz+7QFJJprYkgt4L5KdCXdQjlQBIDqfbpL0auUnDtxRs1QiDFST2/9g6A4/XcMHLqZjrWQ+5QEQ
lfs+pH0Ioh0uV5XhyrDFLotIqygFJ1NbUG/f28IcyauwZ7KtLIOWADGd9+eU4bjvHVd00Gx3YlcX
sf27IyfJ/nOjpz39BXtpZgNe0Il5HD/vnax4G8HVPiehNEzqoO58eXvkoUapDDGWMTl3jFxh3Ykg
GB652Vo+v7rt8tlZQIY2cwXjcfywyURAOeYLldNIUPz5gxt8ry1m5JHP9C4/9DtGzdDL4+cpGkFa
vBGNgshPg6Qyh4pGd9Jo64MvBRPOorNujrX/8q6o0tGrkFyM0NjD5qD0a9PUigHTcdyEdFOshTO5
c0Qs0Tv6S9hwwJEyKGevrPc0CoKp2aQvTqwBNQMrK9OXcs4ttf+vOFz9cXQ891gvcZJ+y/sdFtfF
Ckl4H8nyDeIZZdIHWY80td0P5nwJOrcS1isPmnOkiAZaZld8mcIlk5PSwwa5DvouWxOE2BmykV25
Fqf2pKvBuE08Nx88Lho8rIsVPP5hQmjENOvRN+MpR6Xj/HkAD0q864IZoooJU4Nf/e9EWlfbZCi+
A/GP5squ3j4nlYZxfY8qwlW/L1qooruW9YusWPYEzbPuZBmwwev/Pw/PTwM5Bdupo8Vr6frIGV1y
79sDm2Py0tY4KQvzR8qDNcjjFwSu8hs4W2kpwTJhPuyZkyE2Rfer2WxMByy+a32Cyv6PQWbfCPCx
jmap1flwDJzs5Ef1bZznL8t82kuNBrdfpvf2ecnEOjrpfjbUIQmdboct8C6/j+OM3g9ajexF7PXt
Mbr6drze6xDQ3cteD6mf77plTuCWHJmC33TtsrKFLqkRWsaL68jgL35YyNytDXfMTWUkbYXqu0Fy
5pEdEhrGmvDimyHD9xjxLHzG7xH/3fovDZALVohpWkJAUCKoZTDdhbSWcwefxsqsvrrmPpe1qAVZ
2KKakN3d4UNpzbpNGD7e7sckn8VS0mD8/JxVG+dXXuOo1yEyO7fUErPmIWGKDXFh7F/Q97Fgi1Kt
yRypmBpdLyuNwiD30iQS+bOruzvUVYDsXF+31nj3tOY4IO1s3diEjq7WPl/kbeHg9r6KNLkwonu+
QFvpvsdRWr5k0xK52SZ9v//Q9xRKNc9RbMoNW6EIj9hn5fmCEk9OH3Janww/nMq6CuceWBBJyGYW
VE5024iFa9SitUpXqgPdWpy0kvM/5p5X1DYztnaT7x82PafIofqYU3QezbRFhPTAI/xGYDThz6a5
oHIsl2g8DoG7y+R1+tNN5hIuPNSH/lRL/40yfrO6kM87ODgglKowzew9yopbxV6DCEOTQIwLW29W
5WTSJ+jPIAdQxOm200StwEMtK9Es9rRGTYeQCf58EM0YFJiOv/7j+liF+y6AIJTKkfc99334+fvq
96zc8Nw913iNEJKSFJkGuM05GZXcq2vq9FcOVCZOpaXPPavhqR3Se5jIgwa7h34/NkH0uSvrQEQu
WfdN1c5M7DgRzSLcRwwE6T05qN9W4QGy+ZpoovyQGrxBZo4XiQS96QICPp1UuS5zxzQ205ysmFsi
TcDO
`pragma protect end_protected
