`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
cHDca51msxZj1Clq8H1tvASwn21VMVw2EZ713QtjibBVtcDHNjNhWsu3JpaUF7yS
9jRwJP7FeUapMkt+x7iauG3q27wT92wkUMwKnxxCsgZi0cSCmjYWnJ+G/sQr2hSI
I6UNj+tn6haY3TNFsISbHB+yy4aWpkqJvKVuASazQpo=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
TIE5iBFnnN5cBQszYzhyZRoLU0AGYhWhoD5XTMlQhSivs78klF0pvXGmbIuIyI+l
iU47m8U0B5ENgDT9Q6MVW4kUMaX5uxocTakV4aZBQSKDFwqtnJb6OB2/GclJjeNv
L6vbDsdBuJulu6Eh1Bqe1L7uDl77pTNR+fixafBzG27oQiDQ2Vvhd35tQO6UI3Rj
tGHwKf7BmLEmYPG38KOif9OzV+NECHsM6eE0Jgd0nN8Kr2lCPX0OGHzKFLhzBeOa
F3bCc4Y9kxxi/522rWZm9qhie55vIFvvRZpbFzxBIy5SWUd1GoNJtlzTOKafF1Ri
i/ucU/RVUkInO4FlFFwrGwEy055hPZwvvC3X+EfsBKjKrIuTd+/UgQtVTnskXsHZ
WKx6Z2c4+di/cGKFQQKXGv1BP61h1935G/xrXWMWpo4avbUBGcK9s+kfuP1Iw+1w
OFOG5eECAcrIYWWBltWKi1EckHymzPz88GcNOl8LlnnYOkBSzcywizIny8ssNaG7
MST7lWRqk99S4PGIM+IyN6Ke6m1e1+p6NKRP9Z8bFxwgIBJHdvKcgQdmYwtpl5UR
JFQlEqP6CLwl6xc1jtE8SdYoi9afq58joiU+wYievqFKH17pdDHPBGHOR1BeZOpO
hTjrZODM0eHpjLHBqgP3wrCaneW0hOM0BxXB5adSFJZhv02SEAvYf58xNziywiSK
qdxbbHsq9lv1CV0BpEIjGAlp/SH/EMms+8+dggyd0R34/XjwT7oDSuqmx0NbO07S
FU7ooJlKOOP9IAY2xveYDEVPPY0tckzNY5CtAtCRKeGTw48etk413QNyriWeH0bj
CeZv1O9MndNEIuEK/pHaH5yS0Twh5IWABfN3GXFxs699twN1F16o+R3Tlv3YuKw8
O+BEotweU9YhVFqXa/lDXrShFn+7UvGSqaGnzczHsyCJJfrLQPqM98UlfaiYdlGF
ipIQtkWUNlq4X/XBDIC0FbHMBioFy56iP/0tMVUEC6o9HWK7Oji4he2FuEUU4YAL
EUR9QdOD2xOdxgplvaZRGYx0IkPMDtY58rWmzrFSWYvpSmPs/qPtARId1KblXDBy
E3vFS3nq1h1BKLJHNx3h0AEFQFwMjjE/HvgwfvjHEO3R2+i8mV/+RHDLNch3GCgg
04VEb/yrXDlBWg4HwTm2vWDHdfMOnO1zIgLJ8KZk1UJYM26YhUwsplCbmLZE5Rfn
zZVtHpohsCl9j0ajcWsA8s9ASnIpqmRkU7Zy1pgQIq1T4/18jWv1lrpcumHYGPrH
2ODnDOQaqKcebA2HSTYC95K98hft0PwqODG+cfez+VjJib9mo4SQQckWe7utEM8s
04sjsfOyyG4He2Uu+AKyr2IUjcNQKl1u+TU/W7XURyNLiK8tU5PEx+gIPFA/dgiE
i/iJ6CRJvgR6jYyO5GP61EWE8zJ6VqZeOAvtE9tYFwTaf3xy0vfkyaDI7JtadBZ1
pJGasdtkZuQmQnVmhq4+v4cC9hUYm0bwLW1S9qGSDp40b8zZQK5s76HpAr4DTlkp
ceGK7BqdEMY5+6+RRjkQkJ0PQ1/nnVzWcqjpIJtNeS6TaOHHusIZrvOo3+i4yFDP
cb+fSH5QhlT4cqo3qOwtncZWxOmrbOLURwEwT8KK/ThlrtXI5LL20qDbhvE9cOGz
LUeEWUBHpXn0IKuRX36dINPuV+YuFLCd2oQEw8iGU6DqcbV81LOFhr53PWFIYrdZ
SkxfcMX3JMtMe2IX/3m8Xw358NF/xNt/MErxiKQx8tEhSzT68lpPQovpYxCgBAUR
8Zq9KNEnkv212B8eqls1M4m+JQMyj2IXl8QDrJD+C4NrUhmuA7d6v9b2brH/a8M5
1QZ/UOIVpxN2AxS+Ts8Ii08kkLcA1+GutIPXyRHxdApEbyVQYeUWcDQ2L8lV1YT4
wZtx14J2msHYPFKkx2LqsP2l6nv1rXbqq6oOKOC/iglYGXHxv64MhTeJpIC/eWXv
xr+yy79wQ2RwvjrBcAR98BdEovxdCnaSiRZuUBC9OUrisNZ2+IB3LgzP5304C5kJ
tIQVSH5wG1dcpmFVwTsasZZK6U7Hs3O1BZi3jMFjqsspIryU8GmJSTKQoOEBkqoz
wUgnzF0ovfN+eU+7e8QuS9kAQXwfiPGWu2+vk2HWnS22zx/0y6iZZTsJ0B8EwReS
5Qyfil1dAPllzzZkt7rkAjZZCnB8ZRcOw/ZN+wgj0iOwdVuF28sDsehHLLzfCSXN
34C0w7YXWJjlMQw9qcty/rC4i8j+JdZF1rugnYRsS2yM8UAuyhDTSC09J//7sSb1
EEA0mYaTUvXKE16/HVNnIhQsWwkGBBRBiT3v61/PIvp+RN3/GTe+W8A40a5S3mMj
MviOZT3kicNwv8XlPRGG3Yp00YPaMcJS33KhEjuaDZvGdhKuYpinFeIQjUocrG99
/F/6juaYSv9j8agQpll2PPHYFcUEWyT1tE8mKQCM0lZiJ5vPQwVfNabr78zHwDNa
J5wZYcT+YKDFN7uyW+u4gl770bvkx7AhSYnff16aq8gqJw2p1gigADsLSXbR9Hwr
vtIZurhFy6ezfrUGjEEi9XOrZ3wf+U3vUGq6z1L3Rq1ndKE0lEtH7lPpdWqm47TH
i/ADyFDlZM+VIUXETbBYHsBCW9ae1aJ9f6GDDlxMes6WyvPbBMy9w74bI5SRCVVL
pnIgC+V6m0SycXpg6UEfE/NlWClLrIj5MF9/2RrRj4WL0+BI94A0did1XTfa7mUv
um7UnHnXKFF/rdhhzIVmhdnXjKh/tnDJumduppQB2k51WedG2jf/SePskomzGnPN
HWD3TeW7wWMIhWoLU6PYuzrLthYOgxZDrMJ0JLQTFdsaZf3wQY1sbA913h5r2zzp
q8EVVfdG9cgzDFTj+AFVakgv9t19+9dE/a4LAEcDCUkrfhiBp60egivqmp/3Fc/n
+ku58cE1SMzEnfa4dB2x5SeOkzFAst7XaAvEJubDC4w/TnEdBvKcUOD/h8stDhh/
RhoCsRehVRH8iavZslSg0OV6L8eFIW+mZTb8ifFq5tWE/nynYCR+CQyweLRVuEwU
iRnqCTmjTJb03Ck3bMuuK9pupieGV6scmv+1vSk9VqK1/f+ys7kFEu6VlnOUfClA
KDtN2N9fApqSDEl+mlBvocXhDHF2Q/xVtqpCJ1PoshqdQm8BT25eRMbvcDD35jcZ
BGqYwdG6Ic9DSZN2CxlpJWUImwqAVfrcsfrRZ3FCKE0rJ0PORpOuuv13Y9J9kzet
eB2yjkqKH0JGENZqzh31O3tKjTGjBDSAjvoFv3yZ9SCoSx1WhHFChP1UtZZa37jk
fe7Sdza4i+x9V1c1zneTmS4df4oLh6Ywkdvn33Ul3TSV20w1qXffOhjHT/rbnFuV
uOt/+9gsEQwG3hff8beFxJ1Nw2YK+Kc1pgFAXksfnw9xra1trOoa0hVvn4ja1rxr
Ktw5avovh+BxZecWeElKWyT54C+AqW2hDJ+E3zGzLJzL/hYAlwOOQWMMLFzqoy3w
0sOKgxRBxwV4yDZLE1XUkOpLECwXmg2gRav12Ut/DNPPrz3J8AwvTJtt0D860pv2
30Hp6YQsEtsBWOiww1JjJVDPhoxCCXPoDiv+7zIrhOQSNYXAuY7Mg1LyalITsx8P
x2M5DXO3KJg866HVbwqRhtaHH7qP8sOFQPGCowdAg+RluUOvamIOhVMiiWM+hWIc
zhb0Q63Lx5ypo77Fn+RhMCJXtz7TaYF7aRB0Ihdelk+CVSA3m5vzlRKzFlQP3AxB
1X51776E01kEXKsLpO5uoc7aKASxoWhBHlwwnVyEKatS16zDRC9IfTc7SBPHhBVC
Neg2Bl+0suRoIUSjSKZLS1JREx+e1jVtILhnFCu3QFhW3x1xW8v1ATEuZ68HzKwc
EJhad0iyDRRju2wjlHQJkof9UBMcWGJx9FE8NI+Jnmeu4VhHoFkAlmafUxbDrE7K
tl/HI7LgnEXSfAV3OL4l9wL00VySK1nm7cFRQO0t2/wxQfJmP37TgKdVB9TPXhHJ
p4n1WaupxJyNSy+xmrHvfa78liPfWZTsxMbeMeMIZbdP/UCUSefaIqEXOd/oppIH
cf9iqp8Om85qvIvUBEcgi93+i/jec3S9Fcqw5uj4eGoVIexcG9qoJKXsfiUuz6y9
GzKRJ22le1Uy0I8p1SDmFduetvGEU1yrqXOfRpV3UHNYNd0hsy6ac5CKjb+XJ/YC
5i6ihBX+MqAjUMSpi2QM1yjwTF0hFMSpfhTCWCC4sCI+tqZ3oh6o8tHPPlE1J2oo
e1rViW3zfKVFc1V/WkZq640LQYuWUJf7bixt7n885Jf9jw3esF1k3yguuT4FuDrK
rq3BPwznN9CSnax+a5lijDZRYgZpBkJQEz1Cm7eh6DdDg6SyJVTaCLlFjveEL4sK
uU15SG4Q3VLQwpzOg+o98icmRCH7zn5MGeIhlagVt9QlFHYwtsXLMLG2edLoHj5f
QtEPVFeZH3xwI9zl6ySFohzJ6fgiiDCLJLqjp/4/MUYkwzX0QH8UTDL93m7q7eAn
4rB+MP8Qb0C3RGf1CuPSBHz1SQ8iLtvnbI1f7b6+LZ5osO9IF5eQeKWEtqnVdGXZ
4FEKwZMKRREi7CgwR9QFPGupXuvMsSxu23yKXGJnTm/i9TjOviSRZXYOqdYdQ2Ei
yqFubD1VhqWF7HdSGiyjjT0HLWTY1DmSopjqvhZjYCfDjP/b2brosUMfDHnTz3nI
FOn3Jy1U5zoDfwDRTEQnjvnIuMg5cPuBHVeNq6rX+StvAKC1Jw+82bzt+YipGOC9
LF+twP3X+ZPJHneLoX980tFv+kZQzrweqmiMyN36Amt9K3+JhVLZanBKSJT5biHo
GmMRFxCeJw6+yOdRSNeJZ6JIa//r76K6fUAsTcaJ93cIylG9puC46S9swYEFRAsP
CXL75SCVkMgFLVFu9Mi0YA+5w9ArpyxzJAwQ6NZVDLUL+Jc4WimpReV+B1TnWDhM
NnYMeQKiJoP+s2TW+knjJP5JhofDL7X5eYL3j9VXWQthDHTUPyNvmJ1/qVo+idJx
cDv28pcPbtkziF5I/WXsF8FCqLA4kn9lk8YKSRS5sA2fu0zUw9nP6g9jS/53wwFw
6Ov5O+ZFXnxgz0Zvd9oRMq1rcRaCU4mQulVDw7DW07YtO5nIOYfl/Gwl7+z+oMqc
Aye59fM2l42A2rH8pPC0qkhp93ER3EvrcYNjkhsnChoZq7RFtAMwHcTqL7mmIeYk
RLa5X4rl7mUQ+n8BB5aQRev22Tm0pYIKhTzduL7u9es97s+fMM5sf8udfl+pc8tC
dyOZoKo9nUJ2M1yu9NuY8bRepZOzOGbOkFfaFkY3H+kfisXLJnOrj/qCkJoZ/Qbp
sxXC7pwCVsm250RzqngYcj7UC0w2aNCkVkfJK5uoj8ouD4K4UQ/VfDne9E7q5J/9
RX6CdkPZhNVv9RvWqIlQc/Zs+8ZtTJqo2nt73vG28efRkq67HhpF7oxaXR/cim3F
xvBQ7OeMR2yWzYAY4UuEZN/84ZUVVDysHR273kKFxdfCGeUQQEu4n6fp6W/azM+D
SlfTDRRuDNlrnKojbadxrqUOUHpImGQq2h0gpMiLq99IoFCH58iwO60j++mB0Ouo
g2rzvl+TZ7wYKu41e9ol+w9r7CuZawFrG7JdVAuWUTjl/YAP5LybtbjCmziaI/cf
wpsL1CZtABHoacuw429+qlYwUcs4r+BFzAjeARafn7wQ47LaFmpnEaP2hrR76VQE
/oQtGr8QRAl4t5KUhgS8XLeaYXP15uvl7aw9cs/ZnLWdjunvru68wAlpgv5QE9Xd
PBvVZ4s2csbLNimhv0AxAxoekc9JH8d9hxYxDBavqvUiDepvYKTgEPJCnslkAOBD
2c4iuZCql5hyHhqoePcBuMof+hng3Ntpseckpgn08/+ysbnRHDPcv4pJDgmn7clr
v4x4eDKDj3Ndi3yWBbICUO1hwWOveTlFkKx9PEcrmRSj71X4cSxGhjBev3nqpiws
KhUs21Ud1Vew3b8ZlcHkImGHLjJf/XOSJT24uo+2a9xPjh8EIbizH+2y/pS7xNsp
jYC4Ool52j2WfMgjg/NpQqLn4y/7cexr0M1UpuEPXevzPJ6zAoOnB8mnOwQockPY
oGsowlvk9dU2D7UdUxXmQFAZFps97npDjKlj2ApARP/6LDriez+AgUA29MrZ52u6
ZybddsukMp+LgRnfy/s7n39tuRJRKCOHvB/3IFS3ryzwgxJ/SZQduLFlA1U4kDvF
KjpzecoFsrVO1arONgrVq5hEgRaCZetelSe6hEVE0691LMvZn2qQb0XJitWAKB35
phNM6USoNS9ps1nViZ1O+0ypPQN05gSeGp8UL7eiqOYqhn0MUpVGLOw/N8w5Eeqi
3PoENVLbemZcFC63DqzYxCuK3tXWNulZeYk61HFr5ZZ0AUsIT3bYDbJ5hZ4xJuPH
qTISwDSVQVzYTOujFeHjXLXYW8MFCid3t3wEUykl0FSmykdNh8bzBwnmZwpt7+5c
P8xw5a8zqgh92IUCKpob0EB5RsqaNC87MQU0VhZ5o7KXnTW31R+Gt9jIoUFsvb4I
JjN+LFSGe8t8jalof7GhADSD6kdC6FOUumMyeViqp95DkkR2UE8tPzdDVqzpWff8
vVygFPj0GuTu9eoGMG8XMwWfROvyzT/+c/jJ7Dyd61vanwNrJKkijko2Aa8AZ4xU
JeivfqCLuKKPR35BTy0ixifshdAmW3pzfKHI+qdzGMt+Gvv7U+agdqt6JLB71KJN
0HsplGy7UYekXXJVGR2NgaPYbNYB1ShhN2vdDUsokm0aVS/tjKp4oCc7aZYKbqwm
P9wC+s7iBQw7mEMKhgMd1bMl6nuvOWfXNRqkWMCcBLvkfrTYqe5P/yoGyaazbHI1
mRfiuR3/RPmW2m/JM4V0u6uYXYAc5OB6iUPifE4wRdysO6i/WsZVemm9PFOuWh9Z
jhEb7WRB78+xEDe+9lcULVnzhTISdt3/c/VCJjivkw7f06z2Cn2Nv6lchYh0GQKo
WoWHuilJfxeSlJvmRtDC44BoBlqBmNKuGhRmWH4REprrV6JCsxoe3qqexpA2/JsQ
a1pU/YfhObXWlBWkv186ZaANMw2vj0+BaAqueq00AOXsLW71aP7cwub54TYzvnUB
Z8jlqNi7V75qb3sDpZR9jHs4GFS2fAzxCPipOMnAY15/2AZlL0IuQn0yMeDj9brt
ceEuaZuj4UL6cxJie1ky7njzTfUOH0pHRis2dA1ae5f+lE/4STnINnw71QEXY5De
8S2287hsCSu6LTf56RkHtP1Pbfrr5GK6S3+/+l7jf4jTpOF3XC7KBCKtKRUdCXTv
pwz3q0tLToQQiqkVLtS+h0NIY4lmAnlHfVzbqVFqJ00cFVBPHGosOMmT29bTZkyX
0s8G8MItzoSh59/d65FVUfkRXwL4sHlAD9bi/Frnyg+4zSwWfRvNUqGGbANd1wwn
ZvfzGRhjHxD0R8iXVHroEjj8XfdybEUeXWKg2QPR3pJuf6tRi3155fPSGRWfB4+6
qECuWLAo5yZuskEWNeA1Qg5wT834Glz25dkH3b/tBd9CPPLLRccsq5C2V9o70vgI
M3QxaXc4Ojm/w9xElvnudwR/K9bH7CUvSf/386Wz2V4LLf3TOHj55frsZ/EIJMJj
RpeGZG38gvgvo4wa2GG+RnQUQnAU09yn1v1CpYFbj8jKsukCx0BJuOVoCtOAQQ7F
N9W1kNvj1s4GHxr2kUyBa8g4uyEtRdScOQD6L43g9dYa9F0VKBAzwrL7oZuNWUuK
QgxmANsozx2CLZ1xDpNVudDiLyLeRSD3CYqZ1RviuuOezMKumsv3Iqd0usfl8Hff
iNg/lq/40mNXm2CZ0WSFEPEj7CAnwunGo6VIdutlR4/UV/wqKdwnaAuZ6zM3aCtn
sYTIMe3mOAnT+2aSmdBUDyquNjz0r2J8jnMducwQsKJbOU7XpUz/ssw4/a/zbP39
5FKaDK+kjtNx2NjaSvtTfQbGBsBq9CidLKVDu9cUbWxslSxeC7jfjxiUFUV3llBC
NemsruMyGNY8q1KTMWnPX0NlVyfocYGofyGJRYXB4HHZR6+ZFgkIvQbBjBP47Fn6
9LsCNt9Phv6uxeQWcHExT8BhSw25UAIQqaj0J9GLiYHA8QTiczAhVjdGV5ntOxqT
7LviGrmw5oYsEv1ug3ClflZ6gj4O6EVvYPfrXZfA6Xffdbbn39SkxXKaSKqHvSt0
3ETY6pMJPE+2vLZqbxZ5KvJQEM1XH3e/kd7eWdwRrSKPS9cDqK/70XkasPoyNDlU
mSO/558+uPxDTFCfvQM+xlQRPKBNxA/JU2yMy8rQVfsQsZDLIyutdOWXU84AKdgj
HWoGD/uzqZEXU1+uTV1DJTVpJL14a/PnNkoQ9MWdlWjoy+o/k3sXsJvlKTAL37WG
wDjXFpOdWVe3jPyhE25O2owkjek9N20ft1qmGuXS16OejrBilr9MjLdqsG7VcXuP
Y6O1c5tWapWrFF/PKHI4ncQWo0dqPVFCM0rgJjg4FJMO1ZzmTXmyIyeQOasU+n7I
uQYPf5dZF30Dhtco0HdvdcTkOqePnHto4HLxiMHcdzV1fOmYRVUOuFBxPLdabKlI
nZsHbiYofzDqbTaQPn3NFmaHrpHwNzD7S8id7XbXpC7v3tmNnDAVHEQ30lD1AXyr
52Fl62SFbe5Js8LX3nlJcuI9mFaoRh2qLRQLPJafujZ6GmOFho1TUT+qYaOp/vaS
CSyCeQIE3Y8UinJYKtEbKcNwV+yhak174kDSEpaH41QVn0i2zEj1FarIkfe/L7gH
OMBdU1bmfTj3ZnywQN30uEuiQ8vuki5icyu7vKhryqT9AVd9ML4YGHUT2B1/OHGE
6SjKQFR/zG/AHd5rWS0CkyArcJLD6tPHTx04seFfbVnptZKhgg6V6baysIeeacNB
JI0+5iQxtr0UqNHNp3LqkpUeGZOkgIfM7s8Rq/9BKctyNEaj6cp0yb9xFSG49H4H
d4ltpwB3aVj+IxkXsE6LTWKRsj1FXRlDnEyuzL6mYpNnf2mskI2XpkI4csFFWFky
YYSEYV3QPdwe9dJ7K0DVcRW2lzjD7DNT++ZW4w/RJQhqVWQggGAWTFRHn1/vqdD6
/uea01WtyoPZcCe3AIKoW0mf/a0DsOReQ5acC9X7QzhkVVFHhG0mtYEue37+HI/D
SHVKLhZUfkHdXGeMJGr1idel0ZNFoujQh2+Tcwl+9iJY5SEbATCVxIpIYXEcx8kK
k6EavHdhRCQ8a2ssu49w2OymV6P3Ceb0JNK1COsjmvbFyqQapbvEkrm+2TdGm7aK
H2dPJdEhDldy1zBvGF4EA4htW0YMotTbxiPPMFafITG8zycU2+sWl0XqSF5xyx3Z
5h7EBAWBqI8syiB/xlRQJH5nKYpxlon7V4M6qmlctWAAa+PcnvATaoNfH9Y/1ZIh
YMsppUb2YBBaWsM4sUEKleTz3F+zDQYMn1p0JTF7zNSXkd/rnExFhme9S9FME95Z
geqIG/Rm4YEZRkQ6pYqoSksVd0dSKalyKW3J4BzS+aC4Q9hNsbSavbPAJowxN969
i7YV6qp8CmdB70PMrlNUvij74uWj3A6kg2KpmBOrLG6/Gsy78ejQgbJLOwrW7TFO
cb0pEr9kx5mVxnMHKS1zmQMU4wwesQut0FqAiOHqCInLwzeSezs0cdDNiAe44H8Y
mEhbx5EEWkFj15w0D0tjcADcKm6/qohoMhiDikAMgw3oolGB6+mNiTTCRCE9prvd
5p0k+PBwi0AE+LXi8C9Rei6R54p46Tu4JTOQBrHJds1Jn/JoAEGf7o5O1i//Kgjd
/hQBTEtykBtXoR2tb0YU1nYvanqmYNx7kuBRP4b0yTA4KYHse0F6AMyxKIH3mCdv
Awx+955n0Llz/yQL17dGaX7ZG41F3dp3cSsBafuskjp6DRMiLBXTpPi0hmIHOLxH
HqJMT1sekb4vX4qYqOCEN2rvdU7vO+7L2IGNe0TLPn/8qd5Tf3ft7sUe6cPxqeWM
6U7XFFjqY6p7CtIBkHRIGLUxpwOQwfBGPIiXSKVV0SOKYRoS27rxzTF1lOXib3Te
BSuS9yAEjGrFViEpvzflT4F0lDMjzwI78xFUO0Ye7NBf2GnnmtPMrcWq7DfB2Bmf
nF7avvQ6k2ZZeTUhwznf/XpLZs86atDSUTJuvlfq7pxKcNAw+VBX0ASMZbgmpgN4
7TvGvHHRJAkuLhjwTnD2ggKFteRjRFxMe2EDUK4u/7w6Wf6IimA1aucwq9U+IHNo
sp58Esn3aFFMfj+XJ7cHRa1AYvclaI+JYcbgngRk8NTA7M3J2UBVQC7f/TGC8bra
KskESxue93FJlyhOj+rA8VYIMaDWBn5sDyb/14i0I5r81LUBiOY074U+ccnNXN+o
Z9xVXUH+rJOjIai/hN0iU8b0DzAXgKpXhKSeKq/osYtHa3on8XtN77C9+zGsEi2J
jfayESr33iPAwzJZqTNlHugDtojCKu6ogBcutLYt2hUZqPOkhgrA5nOLwWKlG0dv
ONRCsU+8+zAlhCZd61zp9Mvlz014Q+Wq/ToRl9hKdFHsmiimRkW+D7Z+Lz0TB2+n
ybAq/wYnFf8sHHcgNsbh1pac9z2RAk26xsxJtrq55GF3CNS6FinywWbcWjkdCWpX
ts8P3iogl2iHxP4j1G8+vLgWSA7WpwwQ2GiqjzTVvehqYU72l0UL3Q19eUmQ7Tii
Kiol4ig72oNNb3fmaZXJ9GnLVcMtAsAmtv+lNqFOKY1V/SRQvZ+ojomdlFrU/VNT
d/+Q7ZoT7XoID+Ep9pvU9AygXFFo8Sk0oKkwhEHiOiBezVTHQ1RveykOSFpE2xYw
zi7ozdBQfzQVnicLo70+TiwoBcb1gzmQY2mDGy+XExvAOQiXcppwzT0MseurxaFu
rlhvPJZA3q4MDyXMChmARtXrBH/1ha4SwtQItg5rBN7kD55d1oh/Kh2DN7zemly8
2xVzxep2y+jl04M2YI1Y48pmsejmfFzvwxRz+Z4tbsdZaQBMRCfnA8LiYjupsURl
y0kt6N+Ieuc/hvgW6nZrJktfo/JVWt67wOZg13C8Kb2oKKZLJa/Ir6p4FQO4KNlL
g0qAiftw8iebqkGTJBTY6IfOatZNRQ5rbGqY1nvvkR58VOAFks+lS18vUMmy8MJG
wR4uXHYQ3vK2OzNOzCKcliLXqageeIoWf0Hy4Oux7WV7puXyUUBxMM6+GD7jGfTL
g25G6Ejl6ii6LFFrrj2Tqsqi7ch2X539tDstafrlbwQE01iCyqYVeIv+0Y3igC2x
ZsV/G/xiMYRSNKxxdIsAI8axXUL+lLdykW63uXaFBYzvxhpYCSwmnQ9Mvsn/6d9D
mYZgAIofQ711n8tdwJ5btyGXxE0ReRta5liwUS83CuM=
`pragma protect end_protected
