// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
nquCKoW+vmJ/ODiZMvaxW9Y2Kc6mFG11g4ddMHmi0IJu3s1u74mY86AdBaBBR3TV
91Bk3R9bbuBOUw7HsJx++BCvt/wSRfNAqrufVDlwESBe58WKWG582r6Ha8st9ADc
TlNFcBkNXr0e4/MTyp4F6OCD1hE9NmWUxVSXtfHxDok=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1824 )
`pragma protect data_block
v7a+I+RAi1aM+kaZbFPGwt9/g0C2I7RQMDBfDCT61uO+LQ+Ko7tFK3s1hiHet/ek
pXhXW11b0nBgZ+ijnmdsGyVAWlwyn8P1gxO4I3i9XNgPgej70JOA+SgZSUhUlc7f
j6msmFLycuuxsLk4XxfnMUbh0Ho4dy7KO2LLmjIDl/KLOlhIg3yJLeY7lx1RMxt1
4/qotkzrRnaXpLSfhmg9DNOiA6pRuxwNOB6WAhgHZSNgIs/h8FfJuiJyKLIRC82u
98ovUYoanoGwhUvDk7vx/hD0A2FpovsgW7RU4+DlQUQSdvFJI7qXAzLCmdutozzs
havENnbZCyQ5LFKih3RiZuBCN+A6q440we0JxuL3tqL2Xz3XySG7m11WA6g412Wn
BVfaU/pbctQRC6NMvhlbRwLqjTq+w9Jek1KKE2QrmeiP7DELhqtK4yvMMBDnCWyU
vZgibZ3jeXs18QOP2+776SP1tvqwLfGPEY/JF2BBzYnEMax+SujKphypqPSYw/PV
T+96OMx+hv81IVOy0eyBrsrbJtb5ZJ9KjwSOZPIn0RMjXDPfecXwKs8+jhcsTNDV
/axEiS4u0tNEy6L3hL6fIQxh/9SyAklAVIACqxWoHaSY5soDxVhEk9nkVW7Ewoju
rMNF5y6ReX/0jwHzKN7iSJioZXeRxGPi2bxRh3psFcEJ7KxpZb9heD8HV8AYVvDa
/pforHz5DcM1dFRMG5HraNfKrDoIJBTHiJtvoi0DUAQFeLkxosqrO2SQgxCK5IgA
3ihKhst0wnzr8p+4VmwKh+TNgdxk2fmWk0l0kNdxWwHusxNHvKvM/tcxM92SaV95
vGYVuVu65bOQ3t+Otynu9ejSsTthHZ8TVi7I8ItInP1Auwtfn1+SxEQkisjU1DWh
7fEMvGnNcu9xLlh14+nhQ54yk0uZBV05v2NBT5wuo5T3+rdB6G0ANjUMKlmbIBC7
9WM0YeldHL+0F0k2O2+5eoIHHxqHbBYnvaBxue2fu/NBAmQ4/rYR7NkkgcBEL1te
8ll9QoGmkkPyGkjGCRJhUYkOu5dxwVRyAlxrF/GhcxWaKhPMn16bAXe2F0IbYg11
lMTQxFzs953MLbz04TEefPQ25vwGf4D3MOCA7OgmJLM+0KgTBPhloIUN/VY9rG7y
ocN435Z7GXLmns5I2A6gRRh4taOBx++UYeMH+y4ayjqMC71UDxlF0JAxpAZui0ky
wsKDj53OHrcwcc9fkaOBjwgQrOoCGTKHJtn69LWCVUzr3Zn9BZVZK9z4I+Sh0iID
qyF+Lu2RQ3RQDGoctY8QqvZyi+9uTeduo7nQoLz+9+qzzsUola0iQHjMYb2F9xf2
onCp8sZNpBKm/uuxPeMaY5jej+71wxYpw2vIfQq48UigMhN+rpcYqpPlb795jiyQ
Es9bvG7J+xCcNfe0R16XSmsHLgsQmjPgtyQEyNZMAVvinGFqPdWO07fwteFUif+K
ho7xUCS9LrguXRGQIknl/eM7LiWeq1QOz4WhL8xUAVNf7LoNb89CEB8yQZmfwbTN
eFMYa5OA2aeNM0lA8cppib9GLq25OBmC8psaD2tp+hyQzWIuOqwGQtNpPIJFsBvG
fPXI4dk7mrx+/SPbA1FNiJGWsR7DTRKlvWu1THeV7Z17PIHwiaef7s8uEI1y1/oh
Jnxsw1KDFH6HZsGMGBTXfy9gWdk8CyAmXjqYYLTm0d/0eY07VasnmCk2TWOEP0vv
nL/AWWXMLfkoxxe4TLRWaZFq40KS/Q/neFwRWoQHaJic0SoiWvWUeGutj3CgBqW4
gdb+qvokEQFjPMBbgEZ5PYlLvATQDw7Vm13aYbYDA+XpPEVM8jBDRkl5wBYh4dZG
cMew5L0L0Q6l+nr32etAxqKzHwETcVABLQx3pBpYakJXkeYbM+VIcYRNgVh2ox1w
IwzmWweBHj90+s0MRoCbS4dZKQCegC3Z2gIQiWec4XmXZ66dn+yVjOq1W+dfLZ0L
78LA3sQQFyeYRoSw4xYVRiRy5IHGz0w3neTEFhjOPMFh4jZg+VLDdFGE435jnjWF
7xCl2IxdHVZzhqz95GVsc0Hi/pn0/opXhH8UD4TOE341iuRGp9AVPdeMWT8O9v54
5d7/NCrM1ef6iSulLUZqPosRh01DRo1PAK3w2HHpOvjPTWrNDgzUieULX8t23VGQ
R2CaPYu771AIHr4oBMcvutIfb774h/q0nRmMUktxEeoU1utltXQNQbu/9vIa5Rj6
3iO7l6n1sN0iTq9Avghdx8JHRuWbVdya3Ccoh4Tl+lU6V0uwKRLVthuEwxMkngAn
67sIRc+dkcCCiWR9Vkhxph5nvtx/RQKaSIFQXlViFP1CUXXr6IErY4TBY3/EC+xo
pCnPBOv1zPCAdpxRo4fUhxVo8FbTPuhWD0ANUSmXCl3WY1eks5jI2q1JZRn3U9V0

`pragma protect end_protected
