// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fZ9fXo2b7uVLx5mtCSpTe2sjBV0PJyVo6IpM9HcslT92AkUFLoaswFMinpIS
6Y8X+1nyZWEubygTUfTfuRQ0tyAlT6FtX7qZHA8ZNYdQGPcToOjHaNpgq0sy
P9QfdeAq+Hd4rFg2fpSGUvNxPXBRLGaG5lCKnnsb9omXQRQ+dORBg73dvu7h
O/7ekaBH32TUx2jddaiu2LEBqDtemKYgsBhCNb0+QxXO/wHilphR1C+SHr6V
HAUhEY1wmOzkxjT/1d8I5H846MF+FcILgyzRGhXRoXBbRMrM22wnw5MwNMea
8IVRyilRntSNw5W8KGzKXyT/9jScb1sIM7FudYKgfg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oGSMDDmaeZ+M6z5q2UMIs9OprrBTrnMW79+9V/0Vjjt6X+BkoCHPLUPyMIKe
Hm5RoFqaRWRZP5pfT9OrW5B9dWCCwKYSJl9mfoBdIdsXqtmntJQu8idzg/is
ePbrCgaI4CxHhkbLhEy4DSYEOc6cSat3h9CIPhLcRYuxWEzWV2pFfyOtzkP7
lGZe89Q2ZEcBGFfVjqfI+iNEMEJKqOP7jqVlEoTvK/wG2RBRG3r18iiFfNEE
6lEsAwrWeeqFfskKkMFiHXAtDmtURMzGMht7XJduNG0ZYuD1T41mRZxiM5N8
wX+6bfBTpdxeQ5sKlzuhhLzNRIAjBFADx+9y13KmgQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
arLYDRZoZWNmt1AN0ZLqmKoCnDZjxtkkoYF5QHlxdVtlSsNJfh4fTbzzB3/1
o4cnWQvn153aEIgyCbTpCV2IvnAhVKy3Lzof9FYX5TlALYsVocA9kuXNfjHM
xYoeonvpMk1zXCnyYInjaTkp4ByigKymuK5IBM34de1hOyHBB0L1PcRTo0ji
8Y6nrbNDQNIUXgLvguxfQjVFMP4bFRNuHnfYRwN5pHh0raedjqaA9T4AGQ+J
Khz5fl7dmyGP3roI7ZbqhhYy9xLamCjR2uO0lsF5VrP1sYEsOdKxp/PjOvSf
bq8sxnSMfiA9bM489D1YmYIDNV0B0WtzvZzFoWJb6w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Nz+QhAKvL1itzFtDCxM4vpiYeOJseUsYpvxtN4I98eLYOMSTP27cZhC+iF2b
lBxVSK9OjqAD1NbPOJNTdTXs/8phNAjNr0c4izCB7ueuEju+lSPY4XKZ2WpE
Ht/kCzAJ7Tw12x6NBwWanHmHOUTeQRO4gyYGI4bym8QwJ5LbTIk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
R5v0kZLCcXyc5St5jAyg0Xg2YjOfkBcReGR/2gXKC7IcVaZh7JITZufgJwSV
Dwz2M12p967uXyFx/iSCwTUe+53KrWMg3XzpFfzrJyaJpRHgvbwZRK1CKwiC
V8e9GNyZPAg1D0FHLWxIu5wdRRQKbvTUOjj0Zp4K3LYvd6ww2cwFDyPMI4W8
lxJjsu7LJWhcCH1b2C0SLkDsv2F+gqc0hmwtwp+uCQGkrqLg+ovgL7VHMWpO
1Pq0nNpO6YtHXkOGhx8xKb1OxE2wxVDbbZAWsI+F6WdcbGISs0eSMvPIs6Vk
5rjz2Fi7msZgZzoQy5eYPeBYRNmAXkHsizooQAIiT+po5v541PsrdTKKBbWT
D0CIiPDQiFrvAPoZ0SfCHbf2LmmohHtBtR8bdutnglX7qLstsRakZ4tGU/Lv
nuMAH0/WAzXKOnPtrAPuuiYukHr6eQcRBmZhPw0MKUMTeTozvJK0leIMLy5j
Tn0thxrj91U9MdxyPiUHJWJ5L7BNCzXp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W4gVX96zL6dnDxxpUx71S9tiRNwoKVM75EHaqQOQr4n9nMvKqbG62dA86gua
dZCBOmnNRz6nK528dc+sT3vDzXYPDvqjGENjZH/nuhoS7I+kwSPszQu+wy9U
wbrhwp5168fg3/GMR9F90bB6Du7QP1uh/V3H2v6mbPMdd067qQs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hn5TwfrQfLuj2ISsf5nuutAVrL3JIFtNuKkLnkAHmwFu5KdFBlVt/Nu4aPAf
TmCQ7yU67NFvkWqPDam/RvJesC15unjHEyHlwSgyxi4JJNM4yyXS2ExHz9Uw
EKHQhe+VXOv8YPDJXxtwp94mzOkZL8wW7T5iN8glYbemEtP2DAc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
BhAkxHYJ/QkSap+nsG7s1H1sVYdiqsdWK85HGkSVOmyqOaxGxOAxCoiDlM/k
mFMO121kIq2MfNn+lgl05Qw2mQxxqlNwx3ywMVoUNDaBopXejuFXRWigKYxa
g93HdnkIoKeC5Nj1OXlT4V96r+sh7lgRvyFRtvigNH6mOoL3rkTx1jYrxH39
kNDlyLMKaJsM19BgR/WqOJZeoMITu5A7GESVdF0x5jG+k56H2RhgVS7zwEr8
hjasJnVRYKeJXI6tMqsHCiWmKasKQQdol6LBHm1jWMuP19rBkqvONxaCUpD+
fUE5LaFOBn4deQ/WXkp7xGf57WV3HwMxI4MQ94+xf5DbCXTY5RHsl5pggTDI
WCuvri1aJe7fxB9Qj0GLgK+GvxXPYoHNI0iHl6HDHapTgQlv6L2aPhWtqzQZ
D/fEYUbKs204v9xvFuwmRURZXoexm3kOFa3R06hyV5/krC0JmHosoVsdQZW4
PLaZMf1W5d3v+MgYP/MBFtlObRuc26GpvNxdDZQfc5Nnhvborat7I9TWEpTk
zLr/mcFuenyvr9/RQnUBrFIaydq5jx2RAkFgIahL+c+TTTEEtMxfP3zUDebr
bOzQqA7RD3mipfT18jScMHpTpvUn8dr0mTx3Kba4uTaExVQGpfY7r3AyOt0i
dneq9+pRg71fiVXF7ueoaRLWG7+76fCbUtNiDMECiE1cWsP+eSaUgoieEI6b
D/LFhOfKVC1j8xjJUSfy+RD0L7HgZVPUcJC9fJETiTE+2wu03OLKvBydA0Wt
O79e2pmtnrJk7IGp47aL2O9Wvf7hBm2lqQ7b9zF6blhyLdPWaSyaFuzg/BFW
/jti3oBEmo6Exojo7oaX8QX+UkFwc89SnxA1iqOUTaXQ1C/kX/OVEQtkE2c1
4H30Xc2hqw/JlaQ8aOtOrE/421bcedyfT9fUk4xRFlvJ5gITFE6ocImot+U5
6xrKpVT0T0atC1/HMeIyPYZDW80X88mpqUNH7IjY3SqCVUdpg2f9luLMG8JF
z4ZmXCaxQ8y8q4S1URJx4EVBK+uaMFlOSog1+vGWX5oXuSf/eQMH0RpgmgwH
ZAfGq241wcDmj8Zbf+q0MYuKGM/qx2NGPp31t8eGm9eXOLhOmLPjJ2aDXwof
v3ZLLZaXALgOiluZxBfd1HYACE34zclM+9TxICaJdIl0K1JQShdsVbHIclTw
wz3Lx7UvJzsprrfjSw1fV6yCyeMlMQNd7DLwXluby/K+SAHg0HdySWbTeUes
4ncs3n+60pt9ESjSi7/dMxwoHh8TKWWc5JYx3uJTMQQ5KGD5vmXwMxRJ015g
R6TDk64wz3hjLxe3se7Ue1CyEcgFmhdkcLK7Ami5kfgAxYyIznehY4fo1JHA
zTySgtU+aHgapmysgEwhhWtrYGLdgsD7Zl6DQ/HLUSdEPzdl0AeK/Qh8ZfzI
RZ8MfMO1k5iy/QdraqPRlMhCrN1mFARFksQbuDQi9JsifGjbr1g/D+Am48GO
zeFeuW7KbHCXnWpitibD6GsgTIhSlX13JPV6BNkiPgd2BNN6iw8I+oekw8sz
tq5kurVw/dVJdkYL9CrJGRcUnpvKf3U+R9mdh2Mjh8KJ6idMl5F17xRE3bX+
/U7IuM2AOrDxXAHze/qrHOsIg0307oG2i4L0lPswn2cX7aSq/MsDsKEcTRRM
tONi4ivY/E6KwoAah3fIJkc+dRd2Ku2WKstM7LXZrHP5hRvfAUD7d0E1j6e7
nw+SjxwyBDuo3kYZ5SbhDpzwL1hUUe5zESFm8rf5eeZ5Ick96BvozE8bmXLy
oLEKAKurUJg1HpBHtSMSHNyygwoBP15ceH8=

`pragma protect end_protected
