��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���3�t���x}���u\Si\���b�mY$�o)��o^�/�Y}�;�a^���Ih�ʚOqkG��<=������/�.�]@#�֮K|Y�G8��Ee�
+	{��î~8 ��#X