// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jHBH2H1wi90eOzBbHaHRIqlL9bN9dQwXKMHaKvECL4xb/SDkz4XqCUb8Ufpl
2Fa0Oekp0icV55TTYwJc1zpDd2bI0wgmu/W05zF5Arf3RV17pgPapu8Mv1Uq
XxlrlcJRXCsN3LA7Rozo/cBC9jrKV4Mzun0AQwLJh+bIoIifwaPIoFqQSS1J
24DwElW6y2eor/iOvNArkArEFGPqN0aHxwzgBV/XMREpJbStjuVT5Zpkk+YE
4G+VcRgjRykP/vb0RIAYYA6zsDiXSTYZnPUHrouFtFW5KXzOQjaEKuFl0tDo
smiCVmOjbUz2QQEWXkA7jmSESqFfko0vi1tniIVIpQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qxDtenL0WMQpmN4T8bMg25kCfJ9CTrC/sD8IiYqqjyJ4gCrYp8WhwFAVmqca
pSBSS24dvUvaIG8wHW45bzWX8LI3nhK+gtFTmq6GcxF2ZjwQBo3tbRK6bUs5
BHLdYh6eKNaAOpI/0DEMuJc/QkETj/+SjZIl0dcKmO5uYPkvHsHHhP85sion
bL10nBR+lhhjOcNmS5cOGxsAUjO2N3KuelBwFzsFgqYM/D/T3DW/GwrBI6kf
ZQMIbdzLn+OaCYorfusHgUBjTUToHlh+e+jwWs8ysLG7yXd2en1+Fgpkvp/J
MmVGykp/rkUWERB0eusJQxDpMKCmlMeLQXX9Q/nOUw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qRpNDW+HWMzFtHnpE7ITYAZ9nB8mHAYUX15T435mAH03XuqKaH93UFVoPYdN
2c0WIOGswMlmKkTS0iacg6V5C66Uti1NJCs80YttB5R7MdqCJ/q3Z5Uxp+dv
iOgDeTdPS1x5NE87gU7b96OLOvItDMdtZuhkbfhA56tfp8r58Ts4mWoGulVx
frEZ15vY5ZqLqYGO5G4GPf5862+lNLBJquQ6V63yhkKv5wI1ptCtstm/HIV3
QP5bZciAjS3PdyyUlT/okv5Qvgs7+x/XqY/zL8YfMV4f16xrlzdwdHrvdqkQ
xW1j4pIwMyXET3ZdtzYA4ASv4xWu3+wCZ2v7zB2SaA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gWZRb0kz2KELgbLSRDlXF596CN2zBDRJYjb/qUUbs0AcRI/ROAb8bB9vesqq
u7i26Ch/V08JxFzTNUG1N0W+CQygylh5y0y5DEM2tRq66qNt9E6PnsGPLqJS
vEnXZuiSbMKT3e/B7Zqolvv45XDAonGXvuhBF+FLmIG8i5DocOI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xZq9J2l9zJKEx4a814ynV3yODZWFJ3NuJ+BhwE0Qx0TCJNNxpO1DZGkJtuSE
+56vc4oLESHnKXEapFUY2POzqKoYBEtoqY+X/xHadRasLaLePVBzyY+IR2+I
PaMC//qjhSq+ya9/vxxLYAI8VkME529D7Xda5b3C5iQyvd7VAh99dlFFPlxL
59DaaMsLLuZpubZO5Epc1gdXUMFNwFjhEOn2uranyai2jr7QGoQvs6mjFVIs
SzMRlMzt/b5u8STcH+gXP+Z3IQ6bio3Yko4bnhft9U/HElO1+8Chqle5cbab
gT1aQSuNU3rS4+SUDjn/e0Q85fFZmYxU2gToOGY/m7y7unq8AgahcsDwTdL4
U4W/+BsgBc+S2A3lMJjoh0ssnpYM4H5JH6qql/4O0odREE9kSurQ/rYTq6Tq
kpEU/yqs3C270qMUdRaSu5OXi2duFxNP3LAKiPT2SKZAvsugm/MOHaQQtkAZ
r0TGvlHwnWQsPTGHtsOj+mH2Lh03RA02


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SKemt5kgL8ZGRBhUbFKKSLlJk4YFuv304UUP9pMro3peESHEfifagsJZvWXS
X1inixDBIOV8B1gShx2cVy/NZTC5pOCeLRzw2zm+CmRz9260/kjFrBcSdE/b
97Vx5nrnM5TQBRvhhEkJmrJZxBgtRL0+nOTzdEwk3tkFYPG62JU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g9J5MYOqzz1EvUgRtCIa0lHox3f/nd2BhYOXUZmcDsDGuCgNZV1SgcUvsUKa
pQGGybpYMruOCxSUOELsk6YOvt87XTIC592GAUJ8ich89JEeBoOGgG6kvUbV
kUvla7FU6YLgGqNI3/5cuCjXG4t/KhkyYKuv+Bt3FgOCK4HhXWY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16880)
`pragma protect data_block
c4ZpnSv2m/pnd+6be/EAz+B3dpfjS/h7Z4cWI7QlhqfC0A50FHvEdCuMMRip
4ANtAjChTqjWRPebn1sAEOyvmkccQyWlFr7h9scM1yrxZJFgxe5g+1SUiIiZ
FHh4N3PpQa49pEKZ7SyeJSw6wwH8/E12e1QM2wF0M+0Ayr+0A/WuwKwbVtwS
UKsg0mQ6bM38EdFoSFNv2PUgBIN4tizRofyx+lJSaFH0iB2zw22jZ11jiHyI
45u1jOv4So3Urqs3DXV3HnC1ftMQTd8/f0lHx784lQN9gXvd1xy8IZJgR1QT
StTDunvd3OymOFWL8JJ6i5PvBwq7iYnZJrU+ipB9W3x6KCLNnNnuDnzTY5kt
X4g85l1Z2OUIkAFsiiDi2O8pAynsnZrAgN2vqYJiswr83iWW3J42cIFQKXNH
GA0si5odMyJMzhJXQd56Oq3Ll2iWaCOvMiNcxr4FHCxhOzb9sj2CDDvYOOm4
zvF7596rOaIElcDcwdkzRg93nGrxSp2rT8do5tnTtXzruVcLyig9q2AnTRCo
35YE9eEf/JAytIGmyqvQibZHYQroehGPMgmOKKhEbQHgYolAWD/kXlLoT/s8
s8u2+oHeFjbZzfnIRyFWN2Hfsk5teqrJUGU6iNzE2WiXrEivjXEMGKZigCQc
NGrKsy0MH4zhDMfMWfbiqJZ1C6VZF0vAZ2ulQtc8ZWsR5U0Cqc0Gj3CHFFT2
3RGqJLImUzDm4bQIwcK0U7GRATR7Ef1SZFSWIj9IxW/UxMf6fopazJTw4Yb6
koz2C2qKXpNMhUU/9z1ZkS5BRpLDVkFLMqBUc/tppu25Y8M4tauaOXagzzl+
rzhAFiRRhXFeeavf5wf5VEep41yjfvbUO4cvj+SZ97c/u/X55uir9p5RJQtf
tS2PBw1CWt3fDVpbunt+IXmiGexGNuIf7Goh8z3hqFo2BYRXXSNnGQ090MhH
70qhGyaKqBrmHSvVEV6N9GzAV7Rfh/R7XDp6D9OpEZAuGYclzw2neOIdBYFR
8A+lEWITFHbFg86nkLWyn04wCT96YAl8GZ1VQW+g8lkcd+5+byxGFX7ylRK7
962x8qBTt/vbqSMP4+Cfs06QSoyQyvEdVEdAGBf1DtyRCmV8y/bk74nmh2t4
G4aHbbbgUjBxLs54sABNWD0n3wNQDdK7hx4O21FFAQCrl+GDZ5bWN3+2sjUq
nRZakLWwBY3Ljh+RGejydfkyozQhdoc11BQ8fHv2TTn0MXeGp/Iyjg5pgY8V
ZYrmyDGhAy+XiFuzY6SmeJTQCh360jxp2juSorp5S98880rmdi8HOapJdL0r
LXPCosdHLniDUH3Ly5RelfZuN6Lw9XUEPMPYvXjiYL6ubm/8kqLi4mlCcf8Q
5o/p+yoQhTBtgA75LZ3SfDS8sm6xz7nZSkJBI9hGVIpdghOtQ0wY8GXTwnjI
YfGOrJfBW/930DYnk3i+WP2seWdm7CTWhuj6qsNFtWEcrrgMiloSfxVnqk+I
l9691Rmotq7o1rJgEuJ1rRAWfY15BucX1JYYmalTHgmn3SzsFOEzd76AH+YL
Jj98bF9M+Awxqgvxdpv5k88YQJKntnNiVLR9Jws+53KjRf4HCRZncPALicok
D34geUX0mjhgpfoUOxAfg/3m2RquLWNAWHqa24PGDPIvJR9drWnAYb77dX+s
Wez7JeZxZYna3URO4ZTCmsNkJONCCmlzwllCqnWavhJYTR+q9SWJcYBSmEL/
6hSoT77NmD1NGuOzVMoDxIQ3RtO+NF2HOBbwTn0TwILabvLWcj6N8jHFZG+T
a9qSKWS0nP7kFXSTZ3a+JpfHr9rkwb8EYCuhIdIePwzXN228KG1VJ7TUkQn8
zOIT26PP/k4YTPSE7qPq/sh8SdkohtOVLnO1JKmhAFfv/5cvL5g/opCFb71y
PobOMmj9IgNKJxGFFYVbTIyg+M2PCwXgC/sLABBKj+nQO4wQUhsPX2O8SWKD
o6WaLy8XMxmvPnadCZFGylyxb+p6m1FzezEqm/N7AuurE5+Em1CeEQFHzkXX
9QyvJnChAknN8DYdI/MovyoxQaxaY9tNeAW9LRCwVIlv045UOBERB+5iVeSL
nonKGvzU9p/RnsI2r97Wo8ZwjvteWMQtIw8E41v6kgvwzvvu7vKsTx/tMQeJ
kpKylVCXVuUQ3PY1YoZ3+YNo3t+U3/CiZMC8zZxG+xw4Y5RPSf7P0AeEHuny
IjqNR9DzlN5YZn3anh4ctMtRYHJVQAZ4pta7TmFM3W/WTbRCr9WmkRfNOToh
DLBfzmEAYVdxLcm0YTHLsOIbFUfiUXxuRZekuEd5fozpqVtYPQv27tQ1qjy0
P9hlSe+qVFS8SKYU/YAzKOnaQgd8TuF0cIrkNcHoCgoVtktsqz4xDUkQOHUC
90Sd3eMCWRpX22J/Ko8sc9hZ4Kn5YeoITmGst1Y5+cAZ5PSvzrz1v11hNKcw
TzH2ycsg/uOardGwVqYELf1U7WYTkoOM8UTz0HmGw9kkSwdtyIDxgF7afxu6
PRUYt+jIbiVYbytngRpzMeHB67I35T5ireYAQW5VAso1lyRhmM4uJ89pWtR3
n+CojHLNtTHs24VjSTUTt6WPPF9apkwSWsJFQ/A4EKMj5I2WWHplOYP+reA+
64On1SHw1/aspiV1NbF6fU7OBrhrlul4Am+LtOP5+AvjZsDrmdhDW6pZqbg9
74nwhUzX71ZUspaCNqY7BP9qGOWIhbwd8tDARpcLHPdHCJnieVAfAogr0u88
NMGt0HD0t4PP7/NkDr6SaBZOT3Ijyqc0ENAb1Tcq4msTQlPegw5bDx5/DXN5
lfSmps7L7XXMsDycK+a3U4pxL85ejDjWJtUASisxXkIC5PFFNgu0j3PZ6KOh
GGb6dsiQfuXpqbKGt1U28zb5aXbIVqJEeniWBTNCtGlPl6qIyrXTgq7pZcPn
bASh3biG2qnDfQ3ckS1RRh/XImnigEy2+JL21ELellYBfhLyPFl7Fl80ojtp
Q9hNZ1eSN+0c1HqQvD7WlwrBPIc+wdEFrm/KmQMNoMIILNq+jT4fOqpeHN7w
jQXYcveetAJiEfCf/1xgS4ko04V7T4gH+GwwOVntvVDNVA9rXRdkub6aB0N9
Twh25L0AujDU/K98z5LOyCiw/5n6WzQQ/tt+5bIbNhn8p7kOhL4tLvI428KI
8HN34l03V+dV/+drRn2AhXTWjiNOUvNnsgVK5JLu16TE2sHBxCUsj6Q2mqHF
qwpzXddgtN60+66nABSvTH/C81JH9AxkjH6dglqHok6q57UFxDePGRjIqtsO
XJvGCPKTAqDQ1LgdJN8rl5jcw+nffWVAUHkUBGlx09oxRaHYkUGdvZaFVLP7
UzQjIK4q2IsGroing6qQ7q67eHld1juxWUPERM9JzrDtW5XTT3+75C2yCZnR
JXmruwJgScLgRGxsb5C1Rmh47GOg5CT/66u4BpiyDPvlrMNHsOvRmSx6qYTo
W+ASJV8kW1nRQk9NLKWXJBQlun5pbhofHAbNZv0UEbqbPVtd8QZPKbBzZoXS
en06KzHkYas4ARJbLdNDkzATc6H9Qe4PaXBLQv396/m394hamhm1g9ZX6c5I
CLJORQLeF5OVw/18DVFcwI3Py6gIxdOPzY/OeJouiLcGuct3KZgvYVPMUdPg
wVWwwDXc0V/y2rVmMZ9K4uFszPCXAm1+/6AtencGvldbteQ4z9b6QmPZ1E13
XRIR3i9DLcTygNycpnc+S8BYbVVNrMj3IlxXCDELyxvadXjrpZ8MjUBsmIl6
QPqaUxQVMf6WsbuvJTjIsznfmgvmoqUjkfzUDpiBiYN+uT4MrSedBMXAbumG
KJuEzSF5UwJupJYZ+vIjRvLGHZTgIr9Sq0yj6dnX4ePlVODtdr4Ju6xE4ftA
SrHEtAMM6JywWINtrLp8mJeo4zhvxOrJ+tbqvXUO2Sv2xn8XhVqhO7nCqarC
PvHPeghN8McEYAxvieLkkBI0lffZZ1nB08Fsj6ZD80AWD5y83J14C6TpAy7t
GL+IJ0CKzsi664mK6n/7KQb7j9gHmQ7hwBUcse8hbVq9DKsHh8xsMQ7Z96gy
tXrlOA8eRSyACoz0tdnCAfdU5PUUpt/CftRr5bV1NiOdu+Sq2F4eC4RTqJkv
22NglzIPxs2wb1dv3umhVlmLyY0otpQ2lQMMjv6XDnIYe6q2Jx+1nTkSEwMG
/5ywu9mpy+kDKLaPCgvuWDi3dMeysJXpGPh/kUXTWh6KvSs+5dx/Mk4D4T1h
ViOgMTeI+VWB2RPRFcJT2raGcACCGoLUoVQXStKWWT7/1lZ4EIL5t3YnCCWx
OUQmHegFAQ9ZJpR9Igr4/S/tobM6YWFt3AGRBo5imDnE8xbPlZenSLaWtH7x
NSA5j2b4T089bQScAUJvCN1PQP8dYLKM3t4UkJIY7ySXCdcDkcPnUO3Kd/1F
P8hwnArYE1w0UkGRwdotcSi7TT0+QUViT01amHY9hcMrBpZEri5HC7woag/M
iNkx5FB6eKWVLOSgMyB4AD4htFd/PmcP8SMkoqMEQgo8G/JLkIZ21xwAbcFj
pmX+Z5s7n/18PQf1FwLNPnf8XRP8lTHY6Za9kRtcIDM5a2+uPpg7F6I9WwBi
+sAjqrPoiuHlt9YwFaVtI0MR9shryszSBL8tmj2zIqgReEKqDnC5xGXFT+rI
2E0TNVUfNRLxjUSPKdRqJAbptX6DSu+PN4A8lId4NOeC0GCYVlccTl4E6yTS
zqhL7+6cKDjiYegNSKLvVAnV2qKL50Vto7w5AgZ1FSyKzLtdM7UOIVL5iG/V
ALtU10/jcOzFqYOLw3mnbrQt+E1AXq0Gl8pOBraBXWPOrVkcKoa+EgukctnV
l9fHm7arpbssKWApsR9alANaZXPI1DKNUYBD50oM47StnahfDyzXpmoXdccb
/JpZf5pv+XBOr+Z7O4Wfl7Xn4IktxzmnAwvIVBUlUBLCJ4kx2dlrsjzStouC
laGV07fVU2m1m1hBEabmW4QkJUd98VtwGbUBB2PSZlGShy6IR3GlvAEjESHa
jp1Ad2Yjhzr0zExT4x4oqHs37n1VWw0h8ftsK96m1rMaXEniovqfsJkuEKCm
8g+Hdnhvu1F12jxZsV73QcPRuK10QXf4EsEYYB+nxs7At0Rtzl+e9AcZHQYp
P9tK5kGtZIcRFoocw1+ssTsCWyJfW2KnKcWIMq+Ef9lnODIDjqm9UmsHTt8S
IP+9qnl3wcjC02mEcN60Or3BiW1TepgycBwA2XU/1lk5BjnQBssigLxu7cJ6
jMQ6EPSNG95rJLZtV+2s83UtNupRyJ/HlnMNOCv2fpjfonrS2a7m8rA9iSEw
er8rH0Yy8X28zr2//bIDMqqMAkxXibCGf8j6IGwNABWdTD2OT0l4z0QoC2X4
4/N11kzlfFXmg5LbHbmDgztTmm05vvz3tHhp3W4Q6scuR4d/BJEWKF8vAf5Z
3fGCmYaEvhyjAZfo4vwtDu4CzR0L4OVFDmadc90S/tzzuzXVIHTKH9GbrXe+
WVQjYusOY6S8ix2CCmqWYhKaSE2hbOBpqEZrbnHBD8RQ1alP4EwiHadEaQ5Z
RC2IqBmo5Pw7q2yC55S4nT7fiboH3RLiFa5/Ea3sy/VdTEw9KU5t3Qq84TZl
DPaH6uK/NTbxYv/gRQOwQ5VZHzAn5eHsUT69dU/Ms/H3vuORYY1qGultqWf1
/dSabgpjamjEddLnzxsN/iuSiiVnWapkSCDgtHgqKXIcSuWlzKqDj0l1AM5K
vdD+dd7y5TFXKM6iwoYLgprX9DlYgW177Yb6E461pfaXF4rdYf5VYpEMOADX
eYCxw3jiyJtaf34UHGsUDbUwZWaBPr+pQwRak+3hYySpxl3dKn4Zm6Z8zgr/
0GbHglvWynUPqbfYugNVF9qark69gWoWYYGO6O/RZ4EWROe187WR7ueJLevg
sAwZ/RciGRRt+5NCsSc8qgyokEwh6a27dIbSuL+O3BTn49frC9MeeF1MIdZf
WQGay9O1z6Gb8RnINezF+MQihY/2+oea1mbTwkCGOLTMo96iW24lYdt3zE/w
zECbS4CFnLzyQli/U5cywstTknJVgS/us+LKyv5R8P1xCdpo4+c1yUBB/1Cv
4d/ebeJ2Sj8KkqymTASkzbwq1qETiU8yYi2VehgsBhBzC68ThvJcPTz6Hf9O
aOz+VqclFLbHQvczqFIM4/5Q+tXduMnyZ9vCaSGELNSW2ui9+wZgvjRQ+8Fh
GrQndQS6Ij5ntNyIMU3QzzNUm38SnWOGoz7h+nk1hjQ1T+2KrFlRw04mbwpq
5ZiOCeLI9/Dr3MvGM02OJKZUjicyI1WyeBdrFBNVr6ela94UmpD1wMflhmh8
SNeVFCxAhTmFX9+llLX8/CMo11N2l9LDJvvqbxb261DvMd/Olx7d2cPPMZ8c
r4FBVipYLaaXAGT5V+swoanZs/U1qpEuSra9iQkNywSk9et2ccy1ZZcpixsA
2jzuhWL9UcRuHo3Mx4isSTdBuSV9Cfa48HnyjlYRLQqBOw+539lLFyKjb0qX
GdfUvJZgQiKixoDWZuSQiRgTg0gm3qD1zMqc22cJZubFfJA8teOHUJ7nWk8E
0lsEUnUURBQgB8B6fN4RO9BIjffOBhKGp725oHjDWUG+TpsRQAqjoqI4pdWP
FeL3BF2WpaPhVhizkfxlxs1DQJcwoiKYF43YxW6LBuG8jKQDKgszAJjm0Imq
uDRzvxzEBq9mJnaBhz4FDyXczQozx7Oa9B5BCZ20/BZWCNCFPj9YWOrD/i5t
EehSqp+ks3yPXgFq+rkIFrBFDW2S/RgDk+c2U+G6yfAtHb1qc9oi7rw22buh
qD1ETLmR5+s6oy3KNU3sFwFTxQoUzJABkLabkohOz+86udnfZRAz+dkKRKpx
PbAKLlf9VBnfILe0s4atrqF2nuWtJVYrCIwdsa1JS+aoCUhZUyycvE4zgi2E
MCeGil9thB6cwvXpdOLrWSkWGPe+4u5o0dAz+NAX9q5n/qPPJYq0VvYbPo3U
BXWSnFNLOuN4Jr/qxJ7lZJYVz8CXAlvP10OPVMon6tAM3E47u4o8laOw8m5r
DzsQNz7zv1ZE3vMp11XbUE84JQ2CW8yYfAWFT4mk6mW+LsLVTQ+KyOfWq5QI
dlO2QH9o+uZU8rDgaaVpIDKgBQeMiZejpf9BbeOK+GODuza20i9rao24f3j1
2CP9iXHS6TyY6ALfOFLMjaZVMgMJa1+nEUQOL7suvVWjAYslZBaEle/8JByL
izBmyKaFh8QuyIBEnYMfNA0TEv31gjCF++0hm2jpjICiSrlTcj/2yjmnwbd6
Y9V6kk0ipmlPPnQUI8ehBgF+h5q5S4QJBMygbg9HV3SSs4rC2SY0W8bhMcCb
+yBg4u6Np3xDFfqRsUABmg7JESfX+oYlzTGEFp3cMXFNcRABVZmNOnlwSF9w
xUk+AN0X7wA5Mrpvz10AF8lQPDwHgixhjMB4S/MRvCk60r4KlZX4Ls/rwMJ8
LGrXjoJi4jcaa57gpBLrYaOCQiGOTE18fyfdAsodg1DYX2eczlrfl5Ls7+5M
kulXLfPZiIEyLPH36/1jW+pFq5IjpT20a3EwF0lzRC+gyqOIplZRytzJIiIq
uCufh9U9xfCbwQK7VdJx2nQSnq3YXkB0I4FCIK0M6RkGYlEDe2ucimJSHJrU
r1ZEATxTvP/bN9PhhDk9wyFj3cp+oURbIYz3iergCdoMR1rb9QTGHDY+TrGH
0XcEZKPRgfFmaJ10gzNjrmSWLQXf1MlQkyoYBO0pvRA98xcqIH4eS4YK1/xJ
S9Meg/nelIUSqiQwcDpQwKmp5LVO+91IWjwU5U14FtHsPOlRiC2/5+JzBAv7
EgQ8CDirbW8+blH4VEOwkVPoyRyH0EFnQiUDTXmi59KDHLjJajNmbdOzbEup
Lopxg0tQELYYHGc4GskqDIWHydx7/XadaFlaBEyrb70EmCsm4ZFooDk+XSDi
AlANYZ/0D5DqBrtLmIohsB89VTA2T6S1LbNY/mhwBfgy8uDSIbCfcg0WwThD
1FmeESQ3OpH8lZNlYicKilpAhXU4FYUgTEZeGqoAok7hh9vS8Z8IUf/zTc0+
ulf2I4zJN0LQEqsM5nxglcUU6yIHV4145B5jS/pRyVOOOBGjRBe2eDc+vIX6
Bg/ezkRnFdnsbVmckiOT/KrpRt0LItsqwbi3hppxYZplfCGuq2bESMqeqeIu
wb1H360r6zcU4N2yG6wCO/1CKMLDdzVB2+XU54X+E1gNqtTkJA2GPhm5ZcJe
rc6sCNLUu4j02JuMh/qmEC5drFGUU+yKjR1XvqI2crbfU5AoP45ZPbZxbSmY
iMf1lu0jBrcxBaxN730RILKZT2A+3fZXT51ZUfLyWA9xdQlr7OhhMm79ycOk
4L1CRvfmkZg5G3/7CsCP95BWZ0U7M0UeVc4u0ZNxhTZwRhgiP7xGQ5L6OP+L
sFdakc81+Vd72wVA4kGR2hH2HxCEjOj8hysVV+E6L+wGnG8XTpAMTyrgom7/
KogphJkM0V1EEJzxA0pdw0MSpbhBalE17xbJKAqNFHbni4iYJIUgncOXCTV5
ddVXfTK0Kp4zxe/TSNn2RU0WgqGFfpIRV96+04ABME6RFSKUCnhmmMYaAr1W
C5l4+tJ4jq9uw/6jcEjzwG2nhEQxw8+8qw6eEK7i2rYSaJ/+TLQTP1l8WaAv
XkR9eh92Atcms04MXb3KQ64XlkJziWloxcrxT2kFMKi+kcEM0FJ7U43F9d2d
okgVFKOSzFCOR6aoNYuDhc5m7qe/8Gj332RA79bZztnw7dw3GAy4idG4FO8D
VrW708ybGW5d1Meiale2QQ3FqEDCTv2CqxJ2ueRmX7+7SDIKMAlccpxBON8w
D7siDZ2mDToglV+WPrI+zjxf82R/2Y3WXa7meL9jLZgET0iNQ52kWyAAsLfz
zbD6rOHhrq++2BBOvZA2184vh90oXrTxgZWQiseEbB29wQ/AGiTe7Bs9l8R3
TW+6bQwGt/BMJDR1WsDZ6SlY2beaA/9DVdV+ljMYhs0ZYc1I0ZnjAMyprog7
8uqd2oq831LLG5wjhZEcA33jV0hcvhEcF/f+nhHbLDnzPVLyLrX/VjHV35W1
w8YByGx37Ljdgf+JP1juZI3abe11znakR2GgjML6BI+Uq3zBxUpxTagNWMcR
GV8JbsLorbcRSno4avNNtQkwnbczvYbT/O6k9LUJPHVu/qNupJ6APAKnq2bg
49DSbCShQhwP/Vf3gjifeDssWXj6Vi86Gm0hD+Q/lQRgQuhrLPgtQAaEZazP
NSxnUfcXiDzPqxhHbqyEKbqquWBX/JLKhFmU+MF+EWcp2kX0RQieLEGHgejD
OEfQ34aTwG/OeVJGU0MRbfB53xfaSkPVgeFJYlmxUDe/qA8ZXDZWVSg4OYaP
a4UAGhPfOARr/pZIaJYopHLgGlqLacTNWjLiI1m4v3oqvqydA8kWlLlnM4ga
0PzvxpOe3Fd7Q51ZyVWXRjm7Ny5jHJxJmwjuLh+C/tHzbSuCP9AsiZ4ZeWnA
Lzbv3w3FTaKpkaJDDIYxy6oD3BYJJNEqX4PTPFZt0rUOOQj8RIqz8H4zn6HV
Xv7oj1ieweVN1jRpjj9h4OK4P6on00BMVmW7hL9289yk9aJ4vY2vHvysh6G/
hACha4Si1VV6pePh5ag2+RUKTtXJgjrpUzN4FTy1sIjdR5g5sO42KVWR1CEj
eCNXOF+QwMuPHU2VXu7IfQ65qqdM75gpIzfkpwBW/xBUFsiAzlvCqOfBmQK3
lMqp4XLKLYwyJhpPpeZS6GbSTTq0Vty8u8CUdqtFVIpCx4NnKc4GEvYBVCmX
i6aehiDqmPbt4KSrCpanmehlt7R1N2IIViyugdnKPjOLAxf6/e0ewI5zr8vT
6f2pdsaAgPJ4hd5rS62HT/8l14aKw56RKjlJSK2kjkXVnK1C2r1fYPnPr2h/
CV9Lsz63N2U7F3SriePmSlDgj61WQUXBxg9ga4AB3ZXOZonTIWUu3ZMcCdXd
7BO/0ztIQkrfKLPGSH6r6RnrI/M3pG/8nXS2iOsuRGEBqzCyIllQ4BcY8h/7
5XfbzbIC3S6xOlq0OSmWnYzXkS9ruy2N04iPlsjdFww9oGCik/etVO+c1SV6
fYnjIwXV3oH3XMrjKS9v0MLmibblRRiNyx25gXHD6zVbfx4/LbutUxvQ0Zgi
DzLpEBWQKEMg7apdIniyylbi1y0Cj4dmAcGvQZFKpu64ni8Fgyw5h/SnBo26
aRYiyO014F3jJQhFdnlkMcU6mmRHxnXcBnEcF/R+x62LUWyEP6f3VBTqZtYN
hJ2Qo3AV33kNTKX7dHrNhmevm/GqLGBGHKC6UAxSU6zScaKMK+uZHvml0hSX
IB/0TmDnyJ4uAkxBx3ifNFQfNForn8FYwXyzbJWx2uOAEqXhQSIqZLLdN6hI
l7gyGz2e/Hp1GvxSj4TGw+NDnMXGzIlK1OEeV5EvuPTjnxu9Lz2QRFC74jUi
zIwICBucUnqS6ULTZKxN8qW0E7AgryJoOlEMsfALUF/tJn1XcDWSe6f0B8Fg
C5jqTa2v7Kg4VQmgsiKiAK43AtIwGTvLaxDwcsg3aRZnqxGPYhYU7A1zAg++
ugDxRM1aaiU3jsOPmtxwfTyb1rlPy8J8S0qFiMWQj/AFI9JvraKt/RtTg8cj
prUOErzP5ooOuecaSR1zpJMR2HmiWdh6E1Crle/VE3oIG8NxAKG8AvzQPy70
t/mzqxUBEdfqbRJwrcRuwAKqQYfrZ1E9UwygGEX58Zn+6p4F5uCdydPYRap/
exWUTTZFZkTPly4n/mwcdM/aakTk7td0Aa6bYOX1HxJMDVeAeRN/bEMMJUUn
uBGYHucFjuzeHaS0TZAiif41AwONa1k7WUEn5Nn39r0V8pmS0QKbuDlfpkdR
27VXHCZO6FXS6X2TYUTbyZAhOP46SHMVPp2YWDkvjjkWUJd/Uz6IKK+I8zz8
JvMudUnsCDdi2HVYuRSEgt74E+7z91jeteCeX7d+jEk/v36pmJBGMr5liJP0
nU/6TqA4Kj+LSGm1O+PmdfbK6e6JyabRse29lfhk0Hr1Y5Q5khmW7WRUwsw3
w+t+HcVNPEkPVB9HLDeJQgNIXckj/Q21qIjrk4azPFkd2xRhqcyJ5rDErLVS
eeVaGoqOQTJYMS+0CH3fn2qBN8izbz7hmRDFt/M4bl4e2CBFZmGV4jzPxoAX
tOIN4gtkkH+DOlf7HN7dTCcWyIPoGmWo/2QFY/0ieK02N7PolclYR+bO/IgC
qRwGY1xiC3mVN+dmwMKINS/INORBzBL7mtgG2D4dkVDuddJdjD02tiRitiP/
bzGMycVu/AXrxljxVaOjxXuQR8z+SCsEzhcIGPdLXXTVwAf78xpQZDnfDbLB
6u0IHUu1ijSgxJ97jgVe/XtAA3vQatqCazX2JrS9JQgs/epXkFyXPZ+hDjGJ
Ed2slZDnrMn6KfJmt1FsynyBKS1Sf03JfnWySIICtEQ2QZADTwKxDmvr76TH
FgaBKyRkqw9F0c35QyXrSnYXGPVXDzYFCufQswg+IsjkKPf8PjS7PR41u52Y
Lk84c2J179d7lXg5ijTd9g3YX6kPhE1lizPcKLplXyYXYyd0K30h1lGt8luD
iLIoD+l6jvhc2fpWCCFOStJOFotMwecJNSqzYy7OzvNhzZ84aTTme5+j/mP4
YdU5Ik/tFa+U4DRrxMu2alvKoTMlqplshHpzsjHEuKTNf5qLTEIyLY6n6uSL
umFSPqg3FHaJsZTsYtaexs/yzqGgVRgzpzAJ3LnC4BwIOn7rcv4WU9uBOmR1
QYyJI+89dUw0OQR813xzTfj7dl7xor2WGQzFilmSZbLkmtboVTJ37EqUinZK
B5OcAOyprD8hpsDBkCuWFll9K8tYwgihyEDaSBpEjmLKNunHIg7gQcBB7Nkv
tQylHbKIlBr/YV2e5MVAPHiaLLLhf5bzpzLeno37ks2YwDLqIO5tY+SsZT6x
WjseX+Tosx9+o5fajC3T/SNyx0fS8GrllEErIB3ISwWt177LYRuzavVCEAkj
9tdAPmoiLP++URsdNMrqYzKX4e6wcI+90r5bmbQ5Vfd4xL568kVJGFxP/OUv
HouFKNk1i9hEXW+W9c9KR5sQpyt2RxD6pTr2INsUx3NFMMEL/DSkquecJiId
/RjQx6bilijB5XGM3VHJ46W9dAkEpZf/Io/aI94Jm9tq/++93ty7Uz62Zjd5
fsofXVTQqcJ8nGuf292WPSnX2Gm1bWNb1YuKGfvj5qvJz3C76MQL9sitI6EL
cyHo4WMxnDjwBKc1fUKeZfM59pL542Iz4vGHmiwjoJq6QDl7/djBBu2Yxj4c
vsme6lA1hReOkbmUvqFh+riENX/soKG4Ye7EGqnpoDmJ7olHKjB/wSN6LZ/R
qVahpCrhq7Jfsb0F2O8xgmMs+q7F7PtS2FoAUJSxkX0oNGKv6foGjsjjZpyg
8GH/LeqYrMOJWpsa54vHTjEQDexvLuqNdFHqUuRV6eH31dtJZr8GW58axdUQ
sx2nc7mHmbF7CkhQJCZ7UGuWtwtFiRXx7vwTgCdNU5zraQZrceDWaoqw8eeG
dbL9msR4abB2kM58P105YhJ7XFqpmT6kxhG4rej3fNKOT1XOOgwhro7rJrQ0
BtkYKPI6BQDSQLtSvb3KWH88vke7hW5820TWrW5KeTEEZyfhlLgktiIY27yZ
QAt9aQ5abQBJSZcyk0tyOTG9FswItfTaWatfS+sgTTyinnK7GmaGAKqS+1Wx
kiy6/Dy4DbXizHs5AKbnxD0IW2tpLMzyFcUl7xPln4nJa9uXfyeICF7KMmXD
VkthOo1V2O6tj3xyY57vwf9nnv1trXOm4yP6E6JWXCiR4ux9etKkBQq3JkXJ
HOesi2Rbw4yqxlWgyTLO1bJPKXFtmX+llqYBXcwM0+aC5qDn3+1+B4yyCLr0
O+e3wq5pOtzO4Ce2OmE2wa/Fdw9Pz2F5aph1Z9Qwf/CG+9i4R9wA0jI/2zTV
lev0ZsYRNUD0qYUfr5084mi86w6KCgj4IK8Mu9HV5uLEiLezVLzNKqJq+HpL
DMjTSnN2PL302DXKwqrAyZ/3qbFHLNhMEhNwbvxJ6Sw1S/2Q/S+mWIriXx0D
o1T30TSta7xs+U5R4pMF57Dcd/TDWu92AMv0kaM1rP9smlj67NsP5vduDWDk
2w5PeqIimflLkAKH9D4HAXPvY2fgpJvR1fDOV8UO+9Bjr+JXJnnomm/bsyBC
e3vsNQlSjIba8SCHBa7t/fncVXJ0Gx/iHnpa6koCLR3usA6Q+xpyCwaSckD8
GUMHofxiU8zhJeEJ2MUBmiN0bJ9ZVTi0oK0+l7JfRz1HKKvVPBwU/wY8/MqT
vhoV4fDc3L/6nxqZR9LCZiDVuC63q804Nvx02Vr6VXygXM1YWdVCOQR2BORV
hoSleYUMU0JLECiijPLJzUyqEQPlA0E6JU90EmeD0Nj0W2Q+9P4er8inpWmI
sDA7sm3pW3vyWAdMXb0gXSrgaezeqWazLi1+woMn2GHuatp3F1V0e7pQH2IQ
11zLohvr8h/m3Elcs3ngsP26hZn8M9Tm9uY7tXi3azI9eI71ut8auPNqOGlZ
lubkwCZOdgAFRV92OeEzybB/lW4yLKzJsbAqwcaVt8d5uoslp4dwE+qerM8W
Ioi1q7LZ+H9wsGesdHQWKcatjexTNd5mmZt0gmvJw/rCLE7OJkRKJkdmWYFs
XiuisjaaWBz+qhBYx8F0WWEm8vHHzz3yMpkPdceLdg98B0YdL213LUdnu/dc
4yyLVOGWFEa5CawM6NcWdE/5txFC+irCT6H2KJQiqN46At+pl7yEddOC+MjU
30l7ObUK4fOeSxvGs27T3DRBiQ/C+KkPsAAMVgKhtmAErsL/gMi6z9Iz704R
mNHZ4Ew8xkxSTnMwjXU9IezgcX8v026Gyaa9MFNGeijFPWXMDRmnkvISb7U6
mWnl4mLaRMyVhgpEQ7IGHgKJ2OpN6s5bkL/mHiHwDlVn3zIzRsGrNMd98lzK
9dX5fEENOyV8PA4nF9/s9gksnkZ7aaQeud48AggHeicaBncoilAoHnYOWh8M
9xJIba1I71mniXOlJQLWBpPmRmzkrpK2ZpIYifNdsHPN8hkNhtpuFM1GwpDj
zY+VdUyln3mxDMdIRs9riFFiuK2f3WSakhhGP+9xSSmAl0ed13AKfzPd3Y/8
6yMmzTWaC4kpEqbfa3OEBlH/gXh6WkkMKcrwaVCQEg01ynIeNkV50RDwmFHE
heKRjPDBUcsdcLg3uApqzQeghI/cryYdIELYVAtqTheVekL2E6SzZYdNhslc
35hiI3HOHcn7a1I6KTbnJ2DF1LIVvskt1z1aDvsj+21honujPmu0pO/iGh0b
/9pnxJ+qzvpSTrPk1uEcdydRCIKGye2Qo9DyY9s/X5kmOjWCIyvjaClq8eqK
NlVT4yxuVCP2RRx3J6II+iy7ptpQwMsfajEpyF4Z+4gYNRhF0xh37p5QWNI6
uQ9CPl1C17Q5tHFdvYA+Mw5v88eRl/kv89ND9SNKgbAZiSqF4R6MtnAi2bQ4
hB5JLQDVoOMCaKJhcHpsahVro+jw1puRBd5JNxGHeRRefkYUbUaWZIRgO5c/
U+/p9FCV//vKCg+uOx3sGNPdaamLySNkjoLY0db3ejTxPjSvjSx4QfLq/UYs
eDBtgALoCHu+hiO4jptmYA/XIe117aRoGJ33fceHKF7q5qNC9jxnGXms88pJ
4X53k8lw0//9JBVafUt3FVRdEgdF4xvotJA8mvhJn1dAi2KEplnpS+v1H9YF
0RUXPj1ihU1CCzLt8DJKZmKFv1l95TEKzluDA0LqyzEAK7u3nibiqN5WPvh1
qK63nQlEneWX1LeWhuxJVDWCpn5gIbtTJpDFo8lm7XDv128+Wr8P10y6hhB+
VKkUNyIpVt40MC7USwOQCokF4VyJ2t+zItNwIaxaVjIO8VtwWQ3OMurCZZ6w
lf3x4uG9kudhfc5p2W8YV0c28SrFmdLFpmU0mxqp1v9pIXP536eMaQLFfAw2
JRLn+o7fZw5f97ebxPBOwcxK81s4ch24YtV9kykNipvJ9Y2q8UszQORpWWfs
rf7GDf9Bpm20ifhl+AJ1AXBj0smWYRZJQUrGqwjr9QVpJn7jjkj7afORv+fo
e9HVZ7BZ9nPzp/XsEJApf1gqAH42aZYe3D80VpyC6ZNKLsWVng6yTqmF3w2z
UMD+9CvbctIU0TAXTtC1TCabwUgSnFDAb/BjYumTlBBI8HjcXgpKBA85TALi
ALmC9WPcANzjazdboKqpXT4hHZLW4Ir0mxyUm4rIR2EB/QWl3HReyCAEZdaa
an7B5L5AALvfRgTnKgEGFArr0LF3WqMM15ZDlpQr1Z5Wupbmf/1ZgQOHpna2
oj2m0DsH1YND1QbXWKU+OCx7djYD32Je09fs+UgWOALT0JAvILtRSgsiezN5
RqpCThvdl+2PGKzRrysc+H6+BXow2VIPa34BIuYsUO/y0CQ7FwLTYS2DDlIb
0cL7X3qwT+7pdAVAXWvGt8IjtyqOxZtNiONWSJ5Cp4UmSqKO8eUBO0chXuO4
s4aggbBSHn8WpqKAhSw9cq3v2Kstl0Eg56zGq/M46zuYqlp/pF9vnsATKwP2
Am5xFYmPoVl+AgwV1zNcsuRxMv8FdNe99zLN12GtNr0dMdWamiUujPPIWqTA
zxrcFpkDzI9XxwdCgihB6uq4bMo/1JbN5YFFcT2cC3t1uKTSXq2dh6sriLSM
n57+aTxKVRkOwzTngyjhfxdL9DWkW4fF/tiSaKHJ4j71sjxlLsOwF0GUh5wf
lMaDr/m10MrysQrQA5ycRGWvQIDAZqB3tfyUjkydwKjufL+fsMTuFHwpvNH5
6UwfBwJVyOGh7j4NAizPCnjBFun1Nti2ZT5UGcKtWBplRHMFAbe5Naos/Y1Y
xyhvD2wePgaTnNO6BDDELAK2VlOUkgO2ZRHSVf5QFrcwuIvDCwTEqsRIKAx+
DBuoMxK/IEV3Oq+4VmwTzDOzYZEK3DauLs9DRoF5MyysHZ7FshkRcdApn5ST
HhizJzEZwi8kA8LoDnrYAx1EH8uS1bQI4RATIrFGZSeu+pIzg4CVsi3/DdTN
+YRp396ceZYRfyLntf5qDQTxbacUmBDTB1TJ2ESju9lxjVA8qT96J732pVpJ
PZ70Y3BVcOxJPjCxXCPy9XPSJ+vTrdO0fVaFbU83zfXkyKYX1xOE1g/Kqsad
b7umot/u3OYAeK4HdPRNXJwMfvMybU9SKTeWMJKQfehQbdqRuO3quqv/G8kT
I5YzCpxrhu1nwR6uGWTXFAQMZ3qjfvfWL1MyO6i1mzvA81FAouTWKX0tFzPp
uLX0BrRZIMf3U2d+0t/735Q2bblpRK+h9dkyJHr70oVeLAytJa9BYgmt7Xga
mL8TbkDYZPnvW+LGBRSJ4GWbVonWM62bnOJm2to2v7bKai9j4yLf0SEbJfda
yT/98xSxD0LmPWLHrafLlSdH0dJkkx4l3lEr2nVvuV6jhNbjk8zXEUuw3pD+
E5uxjgC6v9mQs+VXSOhSF7bqnMdE9V3j/LyTPpw3BCPDx4hoSaMrNFKEVFZu
fDyTYdnqVAVFHLc9FtwLTyoKEE21bWu1FyYSsjAIuPNrB5Ww/C7May+pNSQU
wIRJ87L9GIZPBXp2eXrIUAEf0LcQ8fG0F52o5kL2Y3+fisfgS3bt6CZCW6Y9
CyrmpBTpmMZ25ui5yH941liSuetyvS4Wck/5LvJJLOmDU/b9WyDzCwJ2Qnpb
P7Jt/3UHraCsuXJ0DdQw1mIE593jPYc8fni1GuLQ8YK+qa7EuiKn67WyCxiU
sTrsdHkJbuz6V5j3pkJxV6euogU0ePY32sG/M4ZrdvMm9Y9KDbHHMLZJYD+l
nRQqmkQzRFmtKFlNDvN7fLFV0UubO6L3e3+feUqhkG49q6bB8RhVqgK/Anls
NgHS/cy7i/NslzVvRQ1H61qQOJDePcjPjOVynTxaN8/YnvxuOUYUFo1ApxNB
2ZB5sJmuWGmJQ3bofH8X4bXoq64UZB0Hk7DQF1wTGWPCgpZfOUvQsn+q3B7e
MDZOPjvCz2zX7H+qX1BYAPlO5UkS/V8HFg/TJ3HgZeY8Aum/ZIh0NXQVswVp
ElE2WeSstMmJDz4WE4gPp8Vh4U/VKjMMz6c3JksnEJA6a/3Fo4xCzqCXPdIe
iH5fUUDE45tosjfaS0V4GSkh+iBMzLkDJzFRJUZZTvauREwZEXorZQqBG+b1
2uUsXQ4qprBBbkRWtqYzyespzKqxtA60+7cQFkY7T0a1okAtSLrdnHAhXgg+
TpWkL908djrDHv8qt5RqOBCf1RY+gYUcxJbK8oWEQDhKXhoEa+iajlOQO+ja
9CfPcPMCwgxr67lr28yHxIC44tVkF76e6ESBWry6QaNxJ50yOFzjkVtMn6WR
qSbODo5CQXFLr8AUth5sytrapMW5Ug9HSDfkt3OOywrOVndAUGPzsjSADmvM
bDB7JIBw/CB9lvsrqRqOyJRuXYfNWvGlNSZj3rPlaZ9KNyukWLlIX/P3pNAm
DbmFuR1s7h0AZ7mGWchSi/KV2oZG9Tp1lEOe47ltulg/8kICM0Z0z2k95FA9
gNCh+Ao/wfL9tQrjx/vCIxS1Cg0MD87W8tq+8vcfAsPZ6yuz0LyX3GcXtvPp
suoaW9h/X8Kafm1pth7LwwzP0vljDbWVPYd4UnsfoD+HZF1y9r6ajeuvSk5Q
LRGGrL2JKqWR6h+JkBTw0aIFZ4dfRi7B8Ri9SWw8YrtWO9cYD+ejYXF6vG4Q
XlUadNaE9nlWhLI644wK92IZkiKrx9zZ5W5FOOoVf4KWm75BxjHXyhGlMKwJ
O8oiGAmAVktCFVf7EkJYTnkB/aWbt980tSZXHefbFZbHF1BrXH379UneZe6u
srI6iyaQLmAQ2gIMqoC8ZslnFkb/umAOwg+/wXINuw6NVmML237Zh17DpZ6/
iIYDCx/Lka4dxJyMFCZZThzqEV1ihrjrrkXX0Dqym8scLKHFaQo0KdnB99lR
DExb/ov4vL+Fyc9wDc3t9lOt3q74e+3CbCZ02aKBZj9e3GutWZG9gLwXymxw
Ojys3e6BtCeq3aY2TD+N9RoqWSLZ7/OJ9tnMLz5bkXLeG8707I3b2zw0c1cL
JwnH8KZjglvekyl4JwnR+0jejkOdl8X2uOLdFZYGl4kc/WlUu9gGXu/SgwoJ
7ixZuFMFo1md9XdbWLF25gttAOxQbA6qPgpVfqZ8+gGdKPl1X8Cez21wXW3s
3iF1Zuu1ZHOg1EXPiUhKVFTPBuJ02Yvjdelo7+uJzPnmWW5oiKfLuXfSdGJg
r0HDuXMAYuBQG3Kx5YLxbloWS+Zkq9Liq7vYJfdyzWUc+y/ZwEq6SChY0bS8
fcpAhiYqKlRzZdwzb/pUHZjTrFWm74evzDkppwROrGYJcoAZsXFGg6/uxOR5
jorDb+rAa03UOEoPq277/oYSrB7Zqv4UoL3SlgTXH9K2vadnC2q3Y+Olv3m7
yptn+Gk0LqKFWoWn+gZKeR4ncQ7bWy0a4/0wuJ8t3+bt4RnxpCicVAPYYlE5
XzZ6AfiUMxErfUBBYRY1jO48GN4gVE7efk0U+enOKUYSieKH9VaMNw2MxWOI
2h0rCRGoIq7INnSaKDluHxHTdjxOE2TjVf9/lkwgKEs5xRNoNss5UXjM4H+n
NZBUgUBdbzfpPmhqUlPvw8FwSbH+oAN2a/xnYoKkq6IUjQ8SA8o3We5cbdzu
92W0WbXptdk/2nwmj+5Uwr0RnSXeZjqWMChOHhusGOQmVS9Iux112rxUPN2f
umoZZj2rgsyBOK9Oq2kO9j3CLNLie+/rvQ+HBA1ynAezNripjM9QfedLN5un
QgOU9KOpNCYLvyheloqKdDOhHti6vzv2L5YhvCviV/VqrlmwAkw4H2sQojUj
K5syKL2p+UuZQwLyzk906iTnd2/HsBOPvWIXLYwuBHshpwy2geL3j/cAZ8xc
YMf7Xd3K3wMFZaMsclvl2niApTyjy1utNf3XKV1TsEBfI097Bb5Vycs/PkAV
HP6pKQ4r7cuTol/IWD787pyVDozKlyZHgFecde1oi3DRW+q1LpvBXI11ebjM
f26xorIBfXwF3Z5eg8U1Q4Fk3P/QmfFMkfosV/gLrPyEWavrGpAUZgisvSHu
EU9soMucNe78cwA0zY8BN9BjxTmskicSEmxvL/riIeW/EanA5sF5WH6jZBRY
2rZMIRPyupIYo9Nr976MmJghywZbB3Ei6Lwpg/PQVhNq4HGsxPCCd4QsmkiT
pfQGfIj3Oqhi36NCHgbwMKKlgWIL7jhlEGrIefUTZMja8uY9+z95UF5urtkb
L2n4vt8JtoxDfIaLNTpe/wL+DqDok1JaWCAV3w03DwTTYD0VPDEmDA/qDgkQ
7IKR2fwb5gPyb9U41kh0FxXwHv29fe6+ufx5LhWw5m1hEGem1TDKCzRiaXfD
846aRLt0eUAGeiD0wjOajz7ZW+ccu3lpG6Xocy2EOS0nBUQXxzlcdmaLhjmT
dkqE6HkdDYGff86s5F043p9E3qn7hCn6ocaWWlNCYKkvS5htZJhEjQwHv7M6
o41x/lL5sizouLSPiTkctzdO+2oZ2EDh/KX+EEQtuJ7UqKd2vUzXeKtP5A3D
gaWGES9zNnTrnTu7AeDKE6qViOxFtq7flY9eZ0gN1dzQH9oGBpZH/QmbZVqb
Hi23DnNU4m4b5hDwRhr9Xceqay3UZCC/MGjE+WZRhEFvKCvUUOxQsTRzmlCn
AI4vCju+IOsG4/OTA4cHXZC7mjmM85TKiBr4AKYxv4jyAOtN7xUPWHmfO9yJ
D4ZenUhMHQUg3o0p0Khm0+1ZH6yznOuoAIKu7Lb+f2i7rE3fN7b6K/xazmLz
SeU61AvtALvb76dHkBzt2SYYoYMS93MpBgb8bSFohlSVABi59w9lAL1FMaoi
4SH5M229aZRKDxunori6PENvu37PY83P1kFcjiRlUMUPviGvRIJtfXGI/PGB
5jZD6S1JKx0VY4lsk9WWX9Iv5xpZXFNEU7vS47ezbiHagoS8H5ZYV0uboxRz
o7NsBJgcskocPSMQ+4u5iwW2VfCVp9TC00hs7wDjyP4Hy7RiqnuMfqKdYGTq
MLB0bHgCTMkeDMtanzjAjuziD3KlVqdzhaBvV3uIzD38da0hr42TyJPDT6Kx
65zogFbA06qKQZrS/KjIl7WlsgF8bXF8aEyWgiKWtuUwM+84vR3Z1sRLtwAW
nrKde+j75i8im98vR86xpA138YaI5fWP02361/LFfX/+AsgNScJBwRqWWyt2
0qD9DcDY878S7u/2mFThXRty4NU2iiHTFVY1hvePQSXETvkZ1yjhJ9IJJ60S
ubZOaqi8uUd8fhzZ17MyEa2NIEgHAkzumQKsCZ5h1e6b5Tnl+xOC+iCpRNQO
M8Hq9qtvJa5lfQCELn+cDMtfjrzURZK45yRQVQiSGA82VUTxwYbqwVUgwkoZ
MaL3TSLlTiuoGfEL/Up8+XAI5t2coBuihRUXRVE6LqySI5mP29M9O6ytQHIJ
g8dNqnO55dFcB+jbJ4a6Ws8TpcC/W1xhYn/Dm9Fh0+PdsFfKWRbj7uC0xycb
Ts/lvhGQWYBR3NtZxBiNRnKljHVeTf4ZhCCwpwUS08EYWgP4r57bWuyO/xMy
xmzkqrwLJNuSr/1qHhNpxPZhT3g8t1ZOB0hasXryJj6DZuigqpo0F821GZMW
PJh7Gx5Lw0y+rI2jHCjhggcUKpuyf/XMxhhqokdrdp6DGH2Sp6IOyvbQXE6m
9EP24KHIIsRMpzwQArq4aM5Uc4nxQBNI8YefhrwoB/MNobt9VzeKfLbQq85I
cZMH35QANQHc1X8Pa5AstwCqcEWe6AyEINwHTfN+damx4zichwtFcE0+1RWl
NvF86ANniv+iOdba9/Mdfq0vSOffx6GU+v6FqCZjVvM7UoBBrg2zIY6eFudT
1ATHqsBcqQmT/+H/D8HoylB1pADXcg6RGmKZR4fs7X4WrNkakp+KQ2bODRQA
MfZz81/IMnVBd8rAtxJd+Anso4d5M6CSCWnp9iZ3sjHV6o52Kqz3egL++oLC
v93EmAWjNmUhx9b6raZkhVShTolZgRATJYRRbfKj0Q2QsxsZBz12fu4CTamt
7MNJ5TvMe7s2CcX3ON1espQJdDNjDjyxbTR2O4pyRjBKu2JWdhvLLUlxynGr
XeW4kTPnDX+suP4i0rAuz6Ha5+6hjinONcK2+W51U6sdfRvDJ/lmBtOdAoud
0pjAT604XkJFHuwUDBWNWhbt4LKzq8xirUNv6dtFMSGLcXnA2l0dhEuisHlS
HWMY71hpz8DI7W7OQVgSZweqQFsRmyPGMZw9GPINOJ7zn6RXkuLQG9am4w2U
iFriyvQppNbjD9LLxlglRPZgwCefyjmEfIs8eLmymqyh8iV9mTUlAtkwoFKg
2/5TaX7FpPIMEd+BR/KA9QmrMFIWZHPWYqvIJ/3pqU9GqLH9UUGk/9ugIZkO
L0ExbNQFN/0I3zlK24/FET23daQnWu/+MX6QADdUnRzSDejbBAwguXmub6BI
MgiJ1HR+T10l3xIx8U0KZ4DroyTXDX7dZiar5epFEFSbKMq9F5g+Kh2mshgo
X961CXqP1Q2vkO701qIy5s23HyQk9LXnfyQ4GYwEB8grtItknkwqVyQf201o
Ba32qkCBegXAZcDIQG4un5ZmFunDBQhkjJfZxaP12W3pSuCh5bJ5E+Ca0E/v
0IpEKh3bopWn0olT9QoMHNVo4TDbevWaCaDL/VYzYewEA2g/EeabYXrCLvO7
aZ/AjEFQtLrh4iCc63RgKliwcgn1PvHd+LKNh1dJeVYOAQ4DI+Op0Y8rKYHO
WIBNA3T4LWgxcGqx5ZfLIg0uJvBGR1E6Rxm3UPCLwZGf16STnZaKUBnagE8G
mFGDmwrspD++CffI6AgWwD6QkepA/fiByFV1GtdxvemE3KNrH7vETtXPtfr3
OBOCgco+9wC6KhBQ+Zi/ulGkC2owNpadwP8Tr0cumPQFdBPX+AB+MI4T9CfI
xqRah0DgO91gyz2jX7Tu0kJCc686t9EzbvHVUHzyQv2ciTXUefjYwCMIcD9a
JFNIhaup39VAat4Bc8rioh0uYw/kFdwspjt52YZTDi67jHrUnVue4AZ3UE9s
NIWLdofzKq/YRebNpERRTfnTj410YJAsugMb3ZXWwOZKjSchFjvyxk0xAoSa
6v364WaLiAUT7afn0BWNhs+hgsmxn+IMQbIn0NoW4XSXPc+8hvl999qHbMuj
Jg1Jlh/pADHjozXNgGDSw59cB0kSTT38+cRXzEqz3zc95zuanh5I6XtTESin
a0fK/Nj/pW1XI64baPK+3rMIajJTJGHKM8n0EUkGGG8hWKPKkivufo2KL069
4ZyE97x9ZsV+VX0HGmvyoTQMMZkiEMZye+bZpU3w43eGe23+NM1T0L0aqnGJ
7yjbnWU=

`pragma protect end_protected
