// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
guuEM5Cr9ULym1+/gIJ5RcmzC0AzGZKIK92oXvb8BJFM/DCR/KTHcZXNVIxp
FoVcob84ydbwDt+gTe4njQ4ig7pEXn1lSBT/8LAo2UNw6/oKOwv16M2IRQzD
uYqBjyiXjh/rEwCmBWDVdwgMo4diP2aKVYhaP6OWlLvt/8MH7kvnBn9L4CDs
0qKMewfAj52KP9W868dTAkh7fLblRUNBqu1qsvBbaam/FpEwAdkBNrznoIhx
9Vc6o0Gp3XsXCuf0NCyvHtNuYIiJ1tb8KYXMIony8i3cOzr6io2f0CNb6rKv
Q7Krtqa/FFzacXEi/f7tzG+y0OMg+Bg4obCYpmKqxw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
isk8YfIEMhva+md7/8oAeA5hFc6IsElEZnyflDyKsAfzjTZYZ3C/R8yFkGMQ
mZCOByEJpdVhd8jgZ49Y/D1BdoC6dLtRBoXN/10flkL2oPtCPNaLyAsl2dxn
hvyV1eLFDt3qbwYgdtbDEvKit0u1ZWFN+Sm3Rgsf695XjDAKKi3TYY4adwRO
d8Ts+W8/B0gbEnsfdFwSpZG+gLV1d+qJLjZtJJROWn6xC3NDl3/B/YXjFKmU
c2g8QWuUc0ZJkGCFCFLivv91aLg9tMLvFZVvrzifTmH2l/SfeolqUweUl1oF
kOGdZ4wFzj85+fhOJYB4Qu7OFosAKjxQP5aFK1hZ+Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hZgN4sp7FWhaphJlowmG/HTG/txnzDlG/ggR7NfX+lJFAFXFZH6LWTThlJCb
/hO1m3QoTU/6A+Vks24QEliSiyx5ePcjaAbTNCtygb0tZpObxF7ADZwkzWyN
VMCQvOlyEiGvK7AtE2+4IWwTPojFDs832HCYFVcanDHLVzT6E2rMEFvDenw5
KXyx0qbWQ2fCZCcKB5IoUL8uuj/8nlYS5D/zZA3o9R2/OB+e3XSURu/6ITvX
X5hsprn/EFlgXnwi/6t4oCUVoRp1PQmfkl2r4rsmK2FImCU8Uy1ZUMu0Bl46
3Er27e7i7IByPVYCAMgwz5ImHoUARl7LK50aXjofVQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ExstZRcWvyMS5fpWdB1Yy1emLJ5ySQsdYFG/JRpe6kZDn4fR+riSVqFEeJ1X
gxLzfKfJx8Gko75dkU4SZkl6R7t+OJdBpsfwsGSJsiMA+LQRQmusQzgpB0bg
yYwfvo8kfo9+SbwKlA/JOo5H4CWrKE9vzdI+t8UvEfY29I0pMQ8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wW34INpEp6muckIsI22Bf67XAE8mwI+S9emILAss6CqXlW1nST7TOUi9008A
Fa4XsPT4WqAW8uXkHjtCfWKOZSDuTs+rJDB6iwSXJECWiNvY7anHkRQv6Xos
DVsGseQT+940Zrwvsz8naGWw4eJyNnWP1qTQID4l2O9pciX6rIYoaVTEqGkP
4q40PkUQ1aXjB/k+giNrKLiSCG5lPs+s8N5hgXrKZ5TRZgoYOcpxF30wN69V
DVeAzp3oTB1M5okQfZLmLruE6+KT6Z3CC0utRyMwcRYPyeB9ascs2YIqnuNA
CrDU614xlI8hIjA6onaEV53vSyccbDkxIWP4zLsqer9Hitz6skCbXa2lMoyq
MOYegyUGyxRG2E0cQkg57D7j1FgQ7QEp7YP/kAf+RQJ7Iq2cVgaNEXnDM0TS
KZ5QNaSod111x14k/8Q0dpz9j7d/CUbxPVLXNJWJZ4cK8wyiZDzNgjiZe2Kj
TGlQQ4k00LVxi/a62ccVenLdYm0wzbua


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fkD2l0pS4obVp0A2X2g2GYQ8Ou0k48RYg0bd7PaX3Ru4mTvnENr2SceQG+k6
2riR5hDXkzxHoKuXhA/AfKyAoeCRt0+AJ+Auu6JbGVmFN3m/ufJ+550rcoSR
FAEvewUsMc23mPd24kbUc2lODj8h6W/Xs937SG7G5BH5OU7cSoA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hWoWhOQM8mdCd3qscV5eGPG+hwDSKBMRDgRRNKe/MwrsLBAOHYdfemSQ4nuk
9ha7V9S1sPULvrikk7GZT7BCZsu0hrMMrHp2n0ez6LYhKnaG1hMsEXSHhO+u
7bL7gt++8C5kzS2qaSPbwaM4uIoRMxcDy+vKvAeYB+Jf2CHQcV4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8192)
`pragma protect data_block
t9g1F2RELw6vjaC4QrcrsnLc8NWkZG5YYC/zCJS/TjbWpuGJ7JxEITk92UgE
TjqtgkURG7AR9h7GwFelkBmDZAaY5bmCenEdUJPIVCEnKMok2QsvULi9QU5G
J1ii4VIadnKp/4gmr9wY+jCthdULxg665aVRwv0qstg2rW4UF6sx/ds96usg
Y8Qq3U5mTkLifxFGOT3EsSlzVmD86NbRInx+Tef8ZeOxb9inI+vCrW3lDV9e
F1ueqqJloroZ356ezPqxrNFc5/DAulIyXJ1rUEktMJUMhI14LDPuqLTa7taq
A5ktQqZOxm4IRcjWGU42sTk4K8d7x4Tt1ksSIKmMOjEOQl+KW0QSvaqJpGi3
cFD/lTDzYHex/vC59CZ/08zeyeLGWspxX/bY+rJHSERa0UZvdGl2T3UfhOFD
X3vg6p3ol6xnC1KiJTFWzcbmEr/vcYhVgjDEtSw+gommMHdX2t+9w7rEC671
eUxexXZHJ4MO2eBE+hxZ5swpmDQoRVayr/6N/gG16tu6IRpkPewkVTFXpcHN
PF2VrWxRIrB+YQb9IHZ37JEcgplW5nmHkSdYByV+0geQc4oxzhr1IbwCcjF7
l4f858PG2hpDphvBTg3lHm6dYnGwYN3r3fFcUo+saQNSTF1sAsnpFMmuA2lL
pEIH6dQUimtMmC9yvE/1jQMap/2aTdTcMmS2P2DS5N/mIdWV0CIJkhdwjXwG
g3KAIQBBIryS+ngAy1glREucRG2lBusypnvEOVuAn7klJWQND14xnZLZ1VHu
otmpskI1tyWLQt/K9xsH/7X3kcs29lt66PV6rCZJh0mo9RmcdGP0/algzEqh
kOnogKHjWCVzsEAb70+FkGiWQG5UhlzOv0A9g6iOsIYqSnR8qc4Y5JuDfNsr
hn2SonAHFipCG1BS7+9dJNwiXrFJxBhZN3YYgwNF5Q/ryjybsTFp86tob1GT
XP7UvU6v51S3uVU1FfuLJtm3s/B6BRuWCVP1xk4PsP16BM6lepM9Asj0ld09
LVpOjBElq+LFaEbxNBjmu6e8lQxPIO0V8cCodKw37fVl93YbM9dlL3HDMW3A
g5cEmyYPDmv7TIW0rNqsIW0kn19tb66vLhIqUrP2KeHEjNixG0oUlOC4iKzB
7E+M6nlzxjSMTWTA9/qmtxGD+zNEEo+w7Ow0JQf2NhHJlPc+YEzvYbiQA40k
UH4tYsuoC6XyoZSRR6aJ0wc+CwnANJxyniyvHIKer34xd9uVXXaPI+Qr3dbg
gmlh5wX4cNVFErYjsomt1oblPE04w5RjUfcsDRdM5WIvTq39Wog1xcg0guWN
LUB9zDYo+SjE2O5EX/ZHx/EEnzyKjwqSzQ1a2MO0Ozdvk5Z7d64VUb0qKitw
EP8fpYWxoPq7l6XHEEJGUBPgm5ugxC8dH0kKdvBRNp6VbjrUHNYUcTqdY/36
t8iNhWCAcUcB4P8qAsEMmqYaCoMJAEZgb1OpInPeOO2JDzfF1udxkUWxc/pj
bx4ZwJwmiaKte8Z812dCF02AucFQw5mSmeRl9YuKnzUhWmY1UWja1KtHGQ7Q
3HMrqaT+SDjc0MzagE0dge6G0LuTgO2jj+gvmDTGYJxh7H05TLATGi0z84ID
BpvGejvbzgF0rK87yhLmE2h11KTMi9gx7AkfF3BTOLSTrEAgRxtCNt43KgX0
bNPUZ+MayPy/uJEc4tzyXAIQTP8tVAdf0bkQ+CvZ+ioNixMo6RSHddWwxxAL
3PYjA2qAdqh9j8L2BVjNRv1HkYWX2K7L2VhgPBFKN08gyLrI7re5WqOKrt1E
7o9dEwlYvQJyUNalnEHHtkA4ZcTxfhtpjX4sc6ruJLRro6DCroY/099v2yjj
pEq+1k3NIkAZ3jsZ8FxOJefQXOMC2Y/yY4VC0bCHbmaEfWcD1qI5LrkwpG3o
EQzm9uG4/DlP/OwTYlTumM74WKhrqyqMnACqX86Lt9LvGGYU5aY059kLbFre
XFgKsk1tz+KHihF9IILmdormnHDKT4g+aqu6rYOf3zFc15AVfABIdZm+KoAC
2l6y2rtghYO8yoWTU1hYCXUgJeNzT+iGVmN+wCbWlOjBl6UyA4eVYw8BiDlu
O5s/ELoiHTa60UnfFZRwcTq4dDJZjcyZ+M0+SELTLgGPgqz6nD4XRC/zLXf9
HPKDym6OAWRT27iTj8XGKFTLlJ1tVnSpZJC5i4LQB7ileIgfDj4XarrGQs0+
sl+qwZSjS3iE7C5IhgnIWftBFXBf497MyXzw6VB8Wty0mK4h3PyKb/iHWcZQ
KaJE1AvL+QxLusOOK73+x9e8Tc/PuZcCGWv7FnHVsg9S4H39TiwTOw1nO4GX
H4dWJqjtX6PaGTkkJQZLBOPC/h7v1o5DMGyzfYLrrRl7UWJnZt9YCB2Ahf7n
8KqRCdnFGUqOA8Zwvz3WcdwkDV8d3yqc3Ot3N+6vQEsh+rSk0yf9GWbY6vjG
k+IQ+lbNR4JwamQd+JDrtmuDBlaORf1s4XkzwobEzpcymFpQNBm1nXpQAFpE
ABHqSLlzXpLCeVaSlThYY4sjhAnJoDvLPsx6yCM0GkligcOqmH3kdlAx4Xts
KhXRhJM3u81MrHygPhVSBglOyEnrj88jW5A9eoydHMd+ygHYr/vaMj+QnHjy
QwZClxJTuYJxZEoC1ZmetBQRPspWS4VVxApf+ljPixD+ATfMR/ncfpJOKz8G
zm3yF4PXtdN0gwTWLNSpxP/cfPwJ7cC207YgZdloQU647tGarifTKZlFVajo
G7GCsZpvjxQ4NOSeQ1hh4s3qTo+KnZ4yDmngur0Wmn+e2YC6+zMmK+6GjeyM
NYrHnN1ppzqs32mGgBepbdTUjniw/Ahp3AGkjNm3BmrAD2oi7HBq0K293C8B
f9ppgS8GdDVjp3IUqzBXoFMzNjXv1VFvviCBlSNoa6QmdbdZ+u7e6kEavKL2
TQJN6S6Z0Q4+TaRLq2pE5PDAxbCpQqKlbXMhyFo0nN9l4Lqr66n1SVLIAMAO
Fdmpbmsc4XvoEgA0fnliyXetYgEBV+Ow/avJvEUL5wHLHsUiKS1W1+AbpcjE
xJHtRYwp4RjaEacT4b/94pRuhXCKHT9daXky8UnkDlzZJ46CBtrFGKzJlzpG
KWlZuf4c1S4JZs1f0WzHwsWMSW17C4/T6D7p0V6M8mGzFaqPbHQRWDIzmJTp
YskhMtVBBHWIWOhCalwmWnO7oWSrCENk9SQmaOPklAGu1+vLkxqv8nRT/uv8
1nuU80YOjz4HBhEsZYUJjXyeokGpv0M0dL9O/lcZ8mjggeDn+ZCqvtFeQNtt
VoA1rPcBULHph7isUq9MuyaORa/6pW/aAOwXER8MfpiJt4WBB8yxYExRhjvt
V00POgCzuur+7cGf9b4D210i/6qZWGpYeV22/boTIgTZLpH7BU0ZYcgSApXc
m3PXbx6440wzvny6S9BhH4O+cAbzLR/Lus4Aw600YcYeprXxKOQekrXf/hM0
hG/aDQMbAnmG3yBDmOnxLoohyitKoeRGR5avfhwNWcNWcXuHayOgfWPU14Pn
nJSVmt0CFHZKMDy79CQph+hBdxxkA0w6S9roij5vhBILPKdi6bHggzg+xGqb
l0JUYuOuDpTbMYjhWlgqbjLKYPf1EJgrOztjhoLbZXYDG8UOgYgZPwVTSbnl
3F48akoAlFma5O7ulnHnYQ35W6m6TeL7050AGKzS4/7155HLGiMuY4dUtYT1
h3Oj/6/nZumqx7qj6pQcyyaKHT6J4s/kX4FrbUjZyAyWHow0PT3535Rr0d6H
Fr/vAxemcVHL9/04z6QWnNkqVh1UKI4osR/YKJDvs9mEE+I0u7jxQrnbBSxF
/PfBfUg4SsicEMt0Xt1psrgazpREDwIS0Nx4P/9ImaOCfnIsArv4zlDlyPGc
kVoGz5RasdGPhyG+TlJSYhkubKH8sTQ/u3aPx9VUJ+K0cuQ4GT6H5GAIj7Hn
lyb8WSovoJ1vhIE++rjyB5c6RqNYrLZsH3nz8cwE2YEZOpNUElVohncZ0CBW
k1sIVowpEXUvKzRKFkPuZWNTNa7CGHPRweAiFfdQoRYvI/a3au8x31t8BDRz
8ikRg19xiTMI72+95ntKOKcCvCgAqx+e3qkYHpjPe+dHtktM5c6IXyuj2bqk
T3yNR17GIkqT5II7PtPU2sXWCDFnE28lduHQ+JPLtTVujrA55Z/L1Olt/AVP
vumKXlklHoEkJSRNtlmg7vneFs7mu3JNQkeVhpFp1qRcoHJcGZfE6nCH7BLK
pkJdsLECvZGrEAKJkQYU4SJlRvlYfMiL/otBxMjOX3uSb3stxOZIqnJqit9K
I8Vlavuvh2Kb6ObYfj1QDUo2jsRD3w8hfhz+eP9lyJx8t2rX4QEKy7Oj+U5N
U8jYgb9eKk8z2HdbIjB0sPjNt71K3foLdYrZ2aW8bYIZ+dQhPSdRvvsXfrbl
ZKlernA1TyzAbz63A8Db4iweZPNbwRaCjJGv6+TGWVHCuUcVCXo4S6WVb8JD
h5bowHYr/2RhQQIq4VsCZufW0CbU0sx1dFi0RHLEGG92nqnfGXw/sMkFvndn
n9CmOeEF/9ncPyh1rQWiVp1dSLWKviwiqafq+VmtLTJFoWVSmsR2kBipQn/J
sCIJK9QkTPfoKREBPT4k+UNAt15rRyHzcb89IK9HFNNJY+JiYeSbcUKAO5em
FGAdZbbfZ9IxXLzHc/qAO625MMwNOAy0YipUd4aFvir08roU2Prc8tfoAXEd
qeGzYXtieU7EvZKKt/ys1FViGiOtNXcudmU0hvzT2bx8GQatw/dBoGNsYomr
vl9t5G7XoH1deDZnnZdFEuetpy2iyvZOQ7g1oMiMbVx2/C7qyxyhOpoIy4to
WEfJvkolnl3hsOMoPP5g6O3WaezWUThMe0TbECkKn07wj2E4qm4+1jdiauqP
kJfl6bOI6NVIHRuKzI9YAjkm7nhL9UKdVR806fDhGBLGw05yryCTILAiJinJ
oz5Est1s6j4UIFPXh5l50GKm2nAULKpGHvM8Y6yUd58PQqubSUpItcHsaKTI
L4np03E5B1YUiEZyKvM5O2FAgGJb2vrQDYW+pUsYTNYhwI/1T/8T/db/FGkA
xbIM+fkclu+Ntgul/QfvvpEv2l80/ohBf3EUcd2gjpbX7xveFe1+3NGx/G0F
joIjnSrc/6blGIMFH901TDLy91Wvqdew70PzZi+2bVpVzvUMvs3pFgue9fr2
WEzI/bT3VCWWJXwtHaR8dEfzzsgJrxBmk7Ukbh/vYNMVCCNy6uEu1hHXuuWD
e+3KN/fffTbELLDsvJAa1UjbcXNsnEEMWhm0qvRcHOO1Mxl+tVM+tdDWFtXs
k8XXypXDSCTw+VdQK13vf3Yj+SP+Ix6JvJDjRz2EBlOeA8Ku0DrW0ai+qYjJ
jUCnRitGywdN4xu63kys+UjgACWgFAdMrwm4FBHQZjXzuxS5psZzy04b8O5f
Y3ywqPdCpw0/AWh1Bt3NzfhBJwI9G2hGJb++/kYeD8/tBVfW75nIleRB1v/9
fAjks3+Dt4HKCry7sieVcW1y+OtcmMbVyu8UINkYkjlkXtLmuz1Cx8hi4Jz1
b+sVmV5YHgmzVo3egbUf8Wl3lJJXZ2qq5H7tRFY6f3+vIOWo+X9P5CFOGPAD
CYRjb9EB40+atfg7d/1aua8C97cxz+2oOhMXZhkAo2Ujh3Q+DRDsKDa6ciLQ
uKK9R/u9Lxv2q9kHYkTw+xAe1TmWU9Jsb66W+YK7zHhxi1ze8fIKqhSulvZ0
z8GOwFvRw2CkM9dyG3EAytR98IcwRckjnuNoZ9q8vm/QdUdYHJYDwVA74qjs
/+6bxYkXcFfFgQoSwxwHAyQV7lNdU4c26CWwrmgnkDe+ZQQ3teWueOzM+v9C
Tm9iD/quoHORPj94n5MLEpPSJXXxtXKOOfUyuYze3Om4nbwx9N1wD6K40fjJ
JGRCBKZh3mlkwzFLtLMWUfNNGBYo02BgbnkkR4wXZu4wvzWMDmh5HZi3EoAu
H45JLSPfoTdB8dNFe48+XNP8lw3ReBhkijXjdaeftghAmrakJe/bTAKZ8d7y
T8EJ7kQxMG78tbP6vpzRhvDmrbzZ/m1LB4wGzi5EaDYsv+C8yX2s1PwGZ6yD
SRz47PBVNGaF9uFOesVKDezkK5WHYTX3+tE00eQYCQE2WvH+nus/FxNJ8vun
rPGur5jnv74goYZZz4wMi6iBHo1DwDCiyR57ZpvYYwhbykouQB0zn2tf3JP7
fBJw66eeWlsnyeIye4CjDHGeFJl4pTjafuk9I0CnpaYqsj3/N5ItEXVPllKO
bBPgd210cZ1Y0UNyRLUa6+oE9Vbv1pOfCeHoQFwmF6P1nRq0J7s8jCYBxgeD
cjwW8JH0HdnGkN2+gpYnrGXrOMaBwrr4Pk8tvoka5+ZRotngAvt39y5IN9Az
4FaTSuz1DN8OnK5EKQrhFHxwiXq57L5asWA6GwRYexVwlJAq2TnQAM0aIZXM
wesPT/MYsSoKjGRuRRP50zh/L5u4PVeZKrIeZJKWP8hu/v9MlyS3tkVipue/
LxsJ+Yz6KET+7Vx6KMwtbM5Gi6v23TIvt4HZXCMFzfjFMEy/u/XED6k/T00J
FD+zwLJcJfbqTEcUym9Si/C7uodtuE660xs4gbORI7LjWJfMix4cpfKQ4kSo
poZXhL6xANTQRsFHE5sIiKTatcspeaS8E11aVLsLHLJW72luNOOibydqfION
6jmV0T92aN6mcLzfiBdwxuWo6yYhjCC1QHd99hSYPPv1DYY6fTOYp1TDWgsR
YDOVmVzUKiOWg+tNVj2Vy/Hj2M7gvbSy89OvFY+QAOCKProZFdTO1Pmc+LQ1
wgxEQo6jaILxScQI/IRA3LYIBnjXNspYAu45v2uFTERyJlPY2oWg9dK0A+NQ
JYPeuIDDY73oZCMxvJpHPLLE9LZaxPUNgFR9tljn1B+SJNGQyMFuhRu6RK4Z
zThiH+nF0SlEbFKDoKvTwwIvfN+uQdvY9CCEzcX+X+k/vFFKGchGOFN4rs0G
VleCieCkACPdsmjIhyx9aAEE/1BqIsnS1c0y1ydqQofmxjuhobYT2/p1jbCM
swNvS4RDGPdQ4id7BjslALh+1zuDWe5Qr65v5uIOAotvuxolQeCNFwdnor90
WYO8I/YKpQGj9MT0Y/1j7VKuzK69f1QFV7l9Z12LaKyizyaygq3Y0zvp8enS
AIl8TmygXqngbMaP74PLKUSeEt0QYUGHAuS5RtxPfW1kd0lXzTRF8XJ0u7xe
iXZxCTZ0hHvR2iAKqTC/goIcmm0a2vJlc29qrvVltjHi1BRxR+XApAIdgNR/
WB4HbEQcREDnki52zavn0IjVATyZq0WIV2/1wta8DPe+UIb7iKPL85+VHd20
AcMcnH2VbTzRuNQlRLHRNYK46oN68tWgX4h1FtzhB6PmAqyYi7ziHJUQHli3
3j+bpVnKJLgKi79eGQsGmcPfrmcQiOOH34aLYjrFsVt2NCqFkGEtn/7Q816x
uGTgo8NV8PqZAfmsXomFm3QyQUP0buRVDvihnIvOFKdMlK8sR/uwVJeoYKhx
h1ujD6iVnK12IodzmgZpm51q3hghlqjK3GqrMqxp/Hoea/FiCuctWSuA5JAS
S+G5fEz+pQERAgIIpH3PcPJFz5ulU/Yz/nAumkWw+JKCI91wnmYbenIYm+Px
E3OFeRUopSLxqGtxD7V4uhYnADqRZlf/tNvuLfr+ciUEgNbJmtERbwSdXgZ/
EEYsDo52KR8dfjTanbBoFeSlTuj/jzB7nyvq+tigMS2sottHjNfmy0w8BxLX
v0PexrJmoe0hA73iQRNScA5drQQgBuqBSyCKTaE79yS8ApfXZ02EzJ8yv0t8
Pxf/4JSD1vxNd/HWIUCfB57+URv5/SMCaIb8y1bswDXSvezn0Rauz9d/0j/T
WVugVYiJTLVAQhLvXRbZt/KjJloUa/GEE5/+Nr8+hhg7JUulnz3vFVv2kjSQ
+v8Gcfd4W+hxx/2ho3gfpapxrOArnoTSARbuzn4DZCB3yB0l4zszc1ZDm2cU
axC84w2XiWEu5MaNvFDNfEVS1f0CuVyVxQwb2Aoib2qh70gPr1seM1eAANI2
bwpVOQp5uEdMiNwk1zg/ac6en5f4ws+FQLYBd4FYacnQhv3xc7hKibModdx/
SahNIYv+MyTjxHARvG1llNNQdM1rRfnPEYvyA8rcst/9XlPO5anXZAcdYrsd
BarI4kPwqPIMrIkwP5Skr8l4aZGT9fCcr45v/nj25VvK0tl+QkufAdMvgiqm
Cg6dCdux84e0ai/xK02j1srzM6l4bUIE04/7Z/R1VQU7dbumwpbnfXiKVnz+
mb9hIVj4jR2hyZ0PbjdrYxJHTVhUtA0EOQYh4+pWwUhtcZNvpMXhroIF6GYG
CzYtlGLKj6Bxa/8BGWtcjvEJhwPIpqewjhqjvxq9eXMxwM794/a9Vywh4XcT
zm/398P3UetBnvXUlfEHhpqilkd9l1vyCdS1BpO0YeFp9E1Z0G/UGG1+lDUA
fbK4OmrgTdvK8DHzea0xSMga9mMlXUm6V7ZIMsKW5HA/Zv3CT0Uj20Q1bBD8
KPW7Ex8LoH9SbofGapP+/IrkcAFqqp4QwOE3nHRLtlW+FDjrVf/qDm2HlbK5
IWJPX0Y8ieifAZD39mmDinZXPCvVQhCrwdoJjMrSA8Wv2aNFbhchWa6sQOH2
/Y99ZHnpxjyH39zHsYYqKl5zuz28u0BTbMz/N55TJ7eNH8cyF23yFpWrxXXp
EflmkQwFiQ0HlrWf7nvnUUgBszCi/3d2d5qeWWXifMrGZW2UV7xtNK0PlMIR
RAl5IkKfIBK8ce57tjMcEvbUtwbfIV1cck/9Ge2KyDfT8efTh/Izwn8YqDdE
adqz4Uq+DY9vzwtP2atESJdm3VMLarRRRFAac5OH2FdrHBIASP5hkrO54I+m
9UGwPg37BeRNxLIVeVGnjAOMWf4fAQ2j6D2hw/7wxF2aQIYSIN4dL+jKyYHQ
NJQ5QvB5535CIX2R16KlsfNTZNl7p0qWXUnjOTLuE9uLeMgWpJEI9AueJlQe
yUfvLcyH22y5grysqo9oeXP1m1+PCpp0Z8BDpceBwmag8L6Hy3QsaAfWw5Hi
xjkmUrIz39SbcPa2Ym3BM5kA0RmAE3Xzcnoei/kpwg2n70J9OX6E+UdFXgCl
ARYJNq7vtFePF7cn39kxOIxPUYEa2Lu7g4lZqPKxGX+c9+b/9GzTLZmcVWvc
Kn5rNKPqMeAzldKbkWth2aPoEJZDPdys4wJOLLRULwERAyd4bkD0UN5TLius
ZRYzCWhBON2np3Jq2BAiRbarZQg1JPthMA/aq9z+jlJ1+aXtqmkPUyXXwJO8
+ihNz2SkboRM2w4DtGPGBItYOMxfFhX/11JJalVnOVjfblbjg1BQyNsNJ7ts
bX3HaJxnb1VyXSIGGgJZ7grL2mEtuCgNGnZIzBh8K03BkU9U7zINXiFAkdlq
+9PFu9lBk5jTec+AKk+PpqMO/bGDkgIpEb09PKWi9tTIS1E3J5+SgKTY9vDc
RY4hh0Sq2mhT5L89NlzbAWYnawM9OOU/qAIoydO7nk6Gdc9BKn6lOStNxNLN
DvsbvMSVvcn4omNK35W1s+7i84ahikjY+iSYm+6uzSMSMI6aOqAi5ITtcWQJ
VJHOY/PtZ3cRzLPPNv9NRCueP/SPZMqU9hhYedjmuplRBzVg1XcMqjafX5yi
ddt3hjQzVIeOTcgYC3MeAOrdbKxSqnM+5t/u2LAyYhN9lfCippl8TpF4rH6+
IUjv+uivFyRMGe8594YBflAn3xtroKyHrBp8O29F3aoKbaE1oE/ZKXGI4H3y
NGAlgiOkDqmLwzc2C1AXfRP39jVchqQTXGHNnfN0Ped7l3jyXx39wPKw5tfb
mn5rmbYOV/dVbxOswnJdcrrYvgbHcAWDQ5cmyh07ZKshlOktk6xkO8166zx2
J2Ac+wAMlAkRy0EppCac/3FshBA/9wLwr46F2QgR9Ccilh/w2G1YJIgp6WO7
n7h4csLhulXiTYZtM4ZStfBiPwO9iED8KyVEabDFBjxh+8oiuVrLFGLxZO4m
J6W9qDc4lfzDjYXcV0nQ1yaaewMcVxbxECFn7vHpnT7JyiCnAiry2MPCR3u/
dQP+B6Set8L8H1w+ou/7IAtA3zC3mok7zyeQSS9bAyUIZM3F5S4q5R5jomqw
5zYaLcWuoVMT1S1erw2RV0JFvuP9RwBOOCB0ivKxZ/MFWcfdRG/buxt8671H
APt0ADktBg8EqJ76aCgONjUO0KQYL7vBtJe1DSt9cjbXTUCe/0ASn3Jga44p
AWRy760sT80R1mTcE8jvyry7jLtDyJsoxTB1iEKNrpxTPuPy4PIzDwiZCJ/1
Dl1d3Y6zqFwfdLppjVKh08F2xtQIRhMV4ewObzOLqzcr+SqvPAV+OJxIyi3x
EBFhJly9fbtuNCkabuxFiLhnBYJSc1XZoEAVsNJoo/BvBv2dAVRB7p+B3D7w
s5ELBvJ8jqSw2F1mJI4iW4A7nezZViEKdx2jEyFBJoF8NJbWXL/Olu9b61CJ
B94h/PTv6KjRsMUVOgRJF4LvgBYLzZ1yu5c8anx47CSgZihaMD2Xxu2XvJU3
Y00Dgjpmtm/8d9EvR9HSnDgxA0OoUBSVipZUr00i0howuo+fxzDSYlkkk3RN
lxCsZTgflj398u0kUkINGPQjEyAj8V4Tg8ebvqqXGvsK7U21u4SWzGrLFNyu
Ydi97wRCPC7j7R0nxNjChQBLGq55gBDt/6IF4hcCp4SfcESTjiHLyCy8MN2v
fJPsUR9kxsS6iptUqLZ1rIwQSULTTRDWX2/eb1VCySLTFB034tJ9FQ8HoEwQ
qys4qneVITKx6rHegCu0kkgrA/HJt0Ulo2wuU0B5A40V4iEsEcMPxYa+gZfC
bdg=

`pragma protect end_protected
