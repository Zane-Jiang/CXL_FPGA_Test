// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rBh/OSuoNj8Boxr0AxGTV9dRjfPwwGInXx7nkQprPPnMHqMWmqYfKyau7xYF
RWVobXuhNQONIQNORoeFzJUaoGTjylVDayuv+el9vVsmzepBaqTaA9fQPH9D
UnIAP2tMMbKk7Usgx2IowHTog0oFwpKhgnJvQVmjyOtGcebfJUIIRslGBGg4
Bja4Ikkc110A0bPc9KTFQ7LY/K6WmS5ue6uqgzDWM9m14DoGqIU4oNlFDsKw
ljCX7NHN79197nym0SIKGAYjgJV2PLkNxDDkD/i6ecf/Bwt8eb8Z2JpX1h/Y
+jghU+Jkj1nfSkbppjGdXs7O/Xr0drXd84LP902SBA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UZNBgszFZtCNnC/IkJJtAu25Z3XcqUXGB/ccO/P6AIWkTpyvHI4+VmU9ndXg
ERcIoXoOuKnt5nrRxIRqMgGUNDB21wEl2T7V6EyE0SpGTqWcroCcC/WiimtO
3TaZY6Qeoz+9PBTLm9QMpCIwWBFG2R79/j+4n+JEpK3ZSP8dIasl3QzblATt
nowqWf5GZynKZZ4M9XJv78YUtQw1YLEHzcmQgtNUaTCKSQAxWQGVCyZ5CNA1
xDA7CeHUFEGo3YtALatwWnHTplr9rV/EcWrSi2xBDQ+kUylo5pFlM+hYTHB/
r+Bwz9MO7X2dAJ0QL4xfrVw9HLx9VwGEj8VL9RW0Rg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kSczvRZVxA+ps9gty/hmnjPsIAWDW57S1zXGb1hEP0rvvtP6Yi6BVA4LAH8S
oLQEgSsVd99dcErRoP5zLTiUFDqDS4+m7lSQeWc2DTPakF0nu92wTLkrhJVS
F5TNzyXlUMrXJLGdpPtOB1S5DT0DEK1O+zk68u7uCa8km0H92pghD0CjV0rZ
CrLLou2+yRvSBpUuoGuLTyQcy/e2YpcxGg0ymMow21P5UTxmqqar6lgacoxx
zUYjV3IZ12AdLspsMx7PMdULYA/JQcOy73eO2wZJEhBUaF0vRDPrMA5Dkg/E
z8CvbeXbfUfiYTJMdkV70wPPPxxOFUL2znDOoIJL6Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oa7EhOnSm+HwpZCrqN22a6jx1ulx24qfaaRlntsvHtHl/snexcpUZ3o9TaX4
gLwV27SB99eR9t9TqDIdpjBM3FJBESF1F/sqgMWruf5blJiVDDQPiVWQQZBq
bz9g6Ns7Sty48HO1caKqUSMzjEUst3G/ichogbwovc9C995HPQ4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
u2uKEoJMLbtZlp8r5+DNWJrKwn82T8pKk/vKU3gpqyC9E7h96CjUQob0DucD
6qek8nz+TDLKhLvQv8guR2ttAUM6olsBcosvEOaW/gh+YIJg150TwnswPM6k
BKpnSqB0+2DzwESW1iRlziE4anhv+54CDJ1WfhNsMbwM/1do8P9nLrntaixY
4VsiCL3DcHF+pLD88aXl3+mLWkRWb7o3IYnuzVqp5svEbrIqRSzBfxCxuBd9
lZpROBjwt47RS4eikyWr0UcCI/JCLjkZrcb7JS9ZaWil/FDssTzZgC3sCFML
OZxDu3R0ciX+wPacSaeUHAWJMglhXyRVdiIc4zMoREB9XuJcJl+2L2nGEgXY
ZQaVAZ7zkjDpf4Fd/SFWFbDX+SSpxTpfP0q6RWgIAjhS98hQu5twGbIk/MAe
l4q08iprCoO0BmfpAuPvZHhON077pU4M7VeQO8mVUq9lPb32WQMstMp8IXVb
C+wp3Eer1vBlD/LdbnaHTwzdFpbs0Yqk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KdirSwE5C3m1DnItsVW407UiFVE/CB+tpNhyNGpi+fzez2dPJFOJmlhNobyu
lQHSEn+QEIaUUTCCL7HNAJVz+VyfoFwQDBNhO39wWudW5t1XgZdZKFF+EdVS
dwMRRwHw1ghhRKIP0soF+AosDgTd/60cx4Xjyp7bQKhQ3of5OP8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dhPTjJ3Jcsagp/43Y1AlBd5M4n+lG0OSxq2bXOfxv2r5zTQQCIfHl0+tXZkC
OFYc6sE5bNzF0TkOnNy0xclNdRB4+QAKX1yMbxcp0oVQSdtDtlCBb4Z20olc
qX5tjGWUwVhZQpC+U7lJZJlUz/rx9F7iV9K/xTLud6rblI9tXAU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3568)
`pragma protect data_block
nsl2q8Erqx7RUDBDZLaeqpyLvkaf/7fwWt6eXgOz+rdL5OrsKD1wXpgNkIB+
RQ/3NqQUcKrnJfzy+DNuVSrwz7FYrBx3rz/CWi4SlXs9LGyazTVnkmOnY+Jk
niY0/mE9VdFoZXelf18azFPM0W07UEY455ru3ik15NApt9D7RXFmejnD8uEW
mwv3xlK2LgZULz2FajeBrQAX5U4JZifb2RkG68Rq+mB5tvoxh7CUJF0e0/jX
wY6uot8FIrzIely4UIQ5kqmrO9iNWYT2xusxsFiZX+zNcSe5Tddk5cocsoVM
a7i/wMEsMrbSpRXcK9XM1yDdoHyr1FTXwUiGJzj+2OBuiH48qgP1Yu5KlQR1
Kx8ROmN6tMr90OSTwOAEK2ovXiA3awPzBwG8umU8lZvyrpbmF3qbDlCz3OVn
Dw3Nxuj81seNuZWY7+G/YEgK4Gq0VzrcyNtuA7SUjrlnGJZXgtqW+zlIkL8b
I4jWhYMlg1gx23LrGM4t4Zzypa+1kL0S0gP2l1tMgpY7ERT+1k5mrgiO9qub
heyYMIhTD5v1w4BESGu0hkHSQZ/a9sBZhkTd0wAGmG+IOqMI8WYSQK1jZ7XH
wqTs5rN3jY/dnK6sBMB3g0h9KMWTA2jTVDObKGhRVeSaT/GC7j8Zc99HBos8
hOu9bwUNL7ZIC0qOuvWHJ+f15Fx17m2Y74BbpJpgHF79VeoVygo0230DVELH
gWzb4wPdlAbXAMwWMTNczbyqstzvmv8X+22lgU3n3SiBIRQkmLaBcgVibhDJ
h4ajRcaw6xPqf5KVufFXEqzWhGgdN2X4nfNfL2ameUbs7mWVJoPG5EWBZg5Q
fQvkOSa2DEVrqx0NdK7lOHyH+1UQu2Zu7oNUKn3oPij73ij4VkPB3whrdefc
qQQlpVQh/UnrvKvnvxozbXQ3O5Pv37uGmLV/RH0xk7kHDmhoiAZyCih/UDGz
YTCsNxa9Cay8h0o58WF4wPi/8oZChzQZpZ9nHEcrjpkoUhSymgsT7OsttvtX
FhQHYsgegxnIlf6tFhC0BDNCSGiY4fNr97C/oehZQqAsKGGKgDrAXOtOARNU
n5sT+CJiHdUaeY1mEiy0tYKuRHTPsf5ZxE7pwolBzZNlygO/9G/jbVY9qQHh
pBaUWpEkwDFrKQ/VtBHRzDH5jKs5YIw5oXucwzPmdPKBX6NUKGvfL+UmMcnU
izcKg0g6khYidzlXVzqLQol/DBm/XKNi2ObxTfu9J5O2kOZTyPIvmW9W6dFp
Tm66MPHJzQSmvLmlEqfOoRiBNuSH/9lkyxo8tXKsvUlJHqcba7XZl1hbnyw9
0oRyK5qKjBiVNbU0tBPnudVf+L8INxuM2+7jJvq9s2SYs3xWvkSj4O62ZFPX
mifWDtywDl4NR9q4Krtu3J4vKpg1fRWchhj+E5+gKBXFX4VJltTJ+/IF1nhg
6BPnJdAs5KEWkBEgWx7YFP501lzyHm8S7kfG/NMdPLeJLJa5Z0WZBmVOTX3f
Bq/2CODYFQPz7FeEnzW0I1xTM5XIt+ega+1vQ0FTD1M+giOXwOaDiBiMS5zZ
FbFPtdW5D8rrMeM5NAaq0ze26V3x4ocZDINFkRhbwzbDF+rdmZ0mQekPKWjP
RD3AzQ4wfACk05ZHEWXaCEX+bv7qjdmVNw6zfVFjYyOx7vEhS6+RqPLauP3o
iBVQvwZ5/HW5ZWaFi7rkNgoaATaSZr+AWcgsMs1Zz7WMGj2WEf0Qm2/3msMD
JJTOBO5Ttemy0n9Q6NHcDZTViVFKGw7DXnAFXAKKmH//KbQd7LZili3UcNxX
WQkEJdVg/CQ/PqBO8Udo2wTLwVQAhs5oTMTJf+lS/sU4vkmuZWcTv1prD36B
Lr7f9sIDpX29LojFwgy6GNat1k3oBQML5CWR5NWGGlYt6L7NaVRwiZXVsF7F
idumAhKDAeXkGK4Bi998GP/5sntcq1fHlF9aGzG6vj69PFj6+tnDBWqpYHyc
khDSgfMOgtXtm3zWc0KT/5CEsAK1WorXhSRxacYazQcBpqmQ8e1lykthvVoe
8UzROTCb5URD9g4lxHhWyKzERPXOvQ7djTDpIUILdjuSJlIpOeUj3zwnzU8n
VTdYdaU+Xpd6k7SxxhD9lea8H7YttKYvq9IHnRKJOYeOcWvYlfjEUhLskLxi
BYduVSorNLNv3uD+b+tfw0tan7jVwyO2o8iPrO3b9aM2LD1EIPi+DtKK4IJI
qjZK5POp3tO5D2Z6lj7nWAtKK2Ee0s8Za/RIA61KlF5Yl0MNEA7AvPBv/NJC
acWTF6KPzOl4jLgrA5cVfGxMWg37730IKdaOVbJy/DsEL+aa5vXcjCgaKhpY
hsA5waL8Rk+8ZL+rz/F8RcX8svbSYqymFN86b3Rzi/imr2XkJDwnfo8LGJIi
/gTbyinYImQ+8n5XzT6xZgWUujDNAUEmaJ2Kzxse69ee1wsIHTsuPoWQoReY
VcRvnNp63vW5Nj2gQs8eR1zETEHwmdtyLoNDyzRKnogOTajVu/W55otpLUxF
Idwt9+SV6kxrqMmMozaZ7e8dsNH0A/JK01Q5CfnlwbjdVXZlyMg4E8gR05Uk
0Ml70gV7GDxXQ3o7Fs9NlkisMKilGfizjEHfBs2RK1bYBkgMyr/G7mPyMAJy
cAMqZ+xHhDptO95B8X711cukvfI88fLR+JBwAXlvZO3RFAzAKBNG7FblDmRl
lu+iNzq/9SNEzdNjfAMVVE5QJ5j82I44AX90Wm8bLEH+JhTPWVQmKgUnssqz
fDDHCMyrSHgFbg2U+Ycm/WTFqxeQnIaM7Q5DBO6RYSazcjt3wYilH6NeG1Sn
kdL0OXTXBcjVKAkiOeSRlgJ9wCN5+P4GDsMaCwE5DcpPy2wDgWUVaH+jFh3Q
O68GorcIilyfd9qZbUr8tOigHPBfa10YngAiUHs9JdOG1OUGxQnzgtfttvep
0+XqcHhYH3nmXcm73JgSQsX/e3B8FOJNTFtYZqrN3vXr9fZHhJaexkjb8J+J
0zwT6TNeJg8aw/a/mBcKlJarMETGkXcVJq+yDc8cqK8qzcxxBJBWqdpTonbn
8jxaj40WIhg0nZ6t6MhhERoMEhPeFj4koIruySrFMpxmIyvJirmz+bprKRhY
BuyxfrplTHVbiQGIFr0JwxZmqGfVOmatFnJdSTsHG3cXQDJTp0FSYAkYxZUI
ewTKu0AB3lFbyqa+VaT6Vd6ggqschO25AeEx6xxesTl2iq8k03R9CpFLzQTg
neZUUEqKX9yFLcREL/2MM2g0JOo37Rb8YAlneiaKQ9XuaVNLxwuhru8RRpxO
NzrP967RcKkWftAtGlNn89hKYFFs/C4IUUI5FW5bKHtuzgUiSLkhy3DB2D4q
4Lurhck2yoT/PqWI83yCrwpbYNJ06JYm1ALxDEovcK6y6CcZl0BqO8mBZ7pX
RdQ1/Vt6TyRoINNSL4YdifGSxXvQF23OAXVFfVUc0hNVyyKz6COC7ejy/zju
XpaFwJFiF5z3beT/rVAMpXVBBI/IY+lkpT3IPAUp/i3uQnqDBaJQGhXobSki
Mj9UYpCzeo84+5bGg2fxjtPQfmGUaYXY3kOKI8PQgzhrVhS8foqgp4TCWRoy
agJ+c9kdaj9ETUxY8toE6dFtArxrV/Qzk56qkIhfwAjd0Hb3mx5nov2ow7wY
zs2k0FxRcsZTLO2/uKpIsvUK5muQrsx2A5aztYorDf548KVyGFtjl+ef4Kju
MNZVlNZdtkiL+PVv+TdTmRQeCZSOLYEK8lOuaJAtoPo5X7HVIV8LvvQKHM2Z
FjYpbedYBW9LJoQfkR6Qe3gIFX72opQvfmjbFDrTlOzqmLJQ1ZjFK8ujHNAM
3MvIjsyyyjGh4U3rW2hmXuHh7+MiMDEKgr6Bu4qMzmK/8eLrXhU2O/c+QdKW
d2LrE7BtPFfOpUehCGtSsFS+vLGYgoa+4nrip/BTTnlGw2lzTXAqbP6nD/P7
wtEhRRdDvhe8yIwqbJKBg1iBsEKiYx/lxkdNmMULWnNhh05R1h21YnfcCnKg
HDZT7zhtFZgZw11pyXAdXyV3/PfRc98XifojVoPRhHkeBFPuxlkZab5sYaWQ
+4PIhIlXTsIvLSoGhPijnVanaU3EieL8rTOrR8GHcagmISVfdA3IENxU4KY3
Yev/CU4BrBpfuSYqbndZA0UC6HbJnyknLG8x5rHU6Pov5+YBDSQ1iQwuDpFI
ZOrKS+etEWykv8r137I7odt+azvEvZ766XrOEvJUu0Yk5eubE3GFTnbRbW5Y
1OsISj35kggA9Z2/UjQB52hdOFZCEXywSTeBvycdfS7+PgebJjhpBlTCYI8x
ozF9Ds36OX0ARkLav9TO14JsHlty+9Kro+REAcZHV9DF7OOeXumqXO96Pxk6
rPeylTKDXdlgYEYFmaZhKpvtIRcxL0sZPVEayjRoaS1llqkBb7LQ3OOo1qg8
8tOvM8hXS7BAArjHRGUMVT1H5x3tOR0UblueLui5FPctc7dL7OPGYg4TNPi9
6YeUGS9LFhWlo2z+Ao6P4HPBJAFPM8tMBpMG5IhkW7GbsUV7PaLFVFOVhkNr
XCuJw0HOf29vlw2oqI+Ut+PGL/2B5vMeOxCLxO3K3w22KuhJp1amM3yTpCzM
J7WFKkVKEsP+Ou/dJmqLvh/05JYarD2LJSCpzWRV5RWLlvcByPkeMMfaNedG
T3xja2QVgofvHZkuNwU1fNaE++3zHXHPGraZsWQ6Nkd5t1JXb/34YGhanxa+
zTcGybzZHpxm6bPtLA==

`pragma protect end_protected
