// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rW9y5/TGo1B3sAnyoIneOevWYvDeH/rb7nSlg4CIPTQplWHmmmABxXtOPRH3
7vSwgQfLqzb2NE4m0IkisuMiZu4kfzeRB9df0LzzrnWHp8eRWDvfQZ6WfQmF
JYjRNl/eytGKIUQ6UEMvvul7PdFJ8dDHo0tjkIvvlcK8AwhqQfcKdA4Hoen2
T02hLrdW6gwND2Q1U3CHew6m7A3WzTDmW0c0Bld4olQF3m+UyVSkD4na8UAr
PC2HtdJJEYLxAhhjcR199lQgMnlpVW3tcA/gLZzx0QTrGKOtQh7p90gZK+qF
g+aN/82x9BVAkVHaBVePFZ0WnXcCWLNpj1vAlyPxXg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Dex1bUbsXBytWjMeda07/fjVDOI79NrJ2gEuQ82GVSYgZPJt+zdTHvq+NjkJ
VFLHa0dp3X2ovbWblPD3Kox++7NNlPaGbBnwULbVmpm6FNcmYaCkIKJtSzIV
ldyHhlYe+Ob1jivSXJLyZBcY2Vglr0WM92YvpcC8QQI32iUiGd09W5o/8jr0
hSVKOEtVZylK5C9LELOljUEgFlUgeqTnvKUf6vsKS3AngLh4Cll6RJslE0Fb
HaH9Nqtslqkxdl6OzL90i8j+fBxrPvSzKzF7mLgwZMbTZy9GEiteUdEF/b3D
clKuXTpCucgY3qnsyb7GtEoerGk8/d5MLtYKgAV/7Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pnec9ZDUy0ILAhdl8CbCOyhSHN/CtV4gZTQcI63mrSqrbJ0RmrxIvw2rx9W/
hbgCkwzSLgnKUgp0+EPuq4K/wzLnElPL2ropuWg+PxuRMo6FoY5CU+s8fX4l
PZBRDvm5CyQQafTK5rvOYEgmP6bELEeIkT2LOAk6VIJETEEN0ZqWZZ2cL1j9
r4UIC3ufEJkkOchTRyz5/WEhjgs/tJyJ6lDuFKobioRoTc8F1dEexdfA64KP
NoFVjvdJ/lXKGNyMjf00pL3MJ0U0eNiJf+9FXAhVevfvtfYw1h2hKS1Y1Rt5
48NOKnoVbg+VVvtLTC/DkEcsyvQOaOVxJNgoaJl4Bg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B8uMRZCPTeimATOg4u2QxXFlsV5IaYfcZe3uWTvOPeFP7lKo+NEm9WwlvdJ5
w7tBqbboqB8iQ+d2gJ0irCcQ8psKKbDLQZj2fhtFZPhE4r8xPCx06o0n/c3y
t7fvJ4ol03YtoebIwoPhL/YzHJRcX7ZytI/IYZOJaSdHLcpTSqQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
P5iN+9LZPqQYzLPVowP9Mebe8+EMN/fvfh93Ani0goUKFERFGA1aW607hM8e
m+WeUMa3wFcIVXOv5DDe8x3yj8XCH/Sycw+0TEamTaPhOqiBA0uC7JcB8dtS
Urf1wgw3O8FGqm6eI3fmPzIfdYfZ7oGGkL0iTXPTPs5Wkc6XLqIeBYx2x0bD
1fVRQ6kPIyXZAeFMNjRcsaBc6kyc/S5U3HpXbtGUaJlav/76YbXKY4ZgjU6u
t+3rNuWp3oj8th8a8cn+OkG4lcVQTJR+GEUKhcNhCBuzhgu8tBYTSxbamdFE
o3VLytQ0cGZGRqYxI277F/+ukMfDEBplbA+EbA/FcQEXJmUnNXt0OY7sEE+r
HMq2QKnfyGECiguXrq8qS++kQuxjUO0GlVDh+MssqGgqWKDbWdLyehKXwoJv
Iap48crlQlEmqi7ri2z/McabEOltr3cx7gh3as/s8lnE2pUlwdFK/rTldjmf
W7pYixsHf8ar2JVrTZ0X5Cj8XVWFwakn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TaX2sclhjlAbXr6ub6bLGkrAh4IXE8EZNU03ejtADSDy1cX/Bizj99DbKwwv
39dY+nZxNdND4MQ+KSOMW/WgYVnU8RrMP3zQL7S2kjALvPh+ZUvIHbaJvcI0
cXNhChHICE2yVea+6+aC2BfUoUviFLuOjhKVEQienpczGzaXefI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LprpV0UKf2pXDdq9fS44W3g/ERQmIG43s2JDnwPJtsS+InH26v92FeRWDaJw
NUbEg1uqZSR29XhrSzRfpwf8/Atwu0d8/c7J5pwlpuNTbrtsGDSllfhlSpTU
2lhhYr6UcJ+Pdq+opoqJv5msLA1g6fGHDD2xX9CLhUpTPd28X68=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6752)
`pragma protect data_block
1tgBrwo030+NETT0En3+GggKgRwrnC7y+zsdAJGVhhNG7eI3F6gx5ZcRXLlq
1bwqM+Hn5QT6DvON4B67+jm4cBs+OWEqIeGP85yadRxz1Zl4leQpMtpydHSv
b5pI1OVFroJZDc9dYsajm2lw8eAKGmrnT3UHPoWIojsiT+rwXHoMwJD+w//U
/7/FU/o1aTOCyVKTEA2UHt7oT4VLWPD/D7HXANakVXXUt51wyFJCuhK5auLk
E8P/3v9SFV1tI79V0JTyPb8ydCu8dWV0SFBO4dz1kbofk/f4uW2z1iuu5laA
7l8K6i+ZuNviHhAJAv5CgRajHCrxVJa6QRXJfOq7xIbIKQ0qX/Pv4csR4DXO
3w7xNlE9MBYKWgV8mE1gG5X43ZFuUeLgLUjFUzA23ILghCM2JvC16woQL9Zl
2OWRSGKKry+XxDf/pKAvXh2TYGHW6KwgAEMqt6A49kRrW4AVHgmuo8W0axKx
/j+BrGcYj0Bd4C15WWwCzhRRQYisS1XITrjCwnGcdfX2vpMtPxL4WENUEtLm
KA3Q6FAuwkuz0ba8TVrUmpXLuhl5sGReswZN/YLtwcvpZ+j5ChEdTpgXC2rC
ps+Wud8zj1xRXJKjYL5uZDBv90hlvzXbxyKlwbZhwTZR6hdP9Q2Xzx2YR2jD
eml7KKPKfBZ+Fso0QIMZsj/wjcbUzVtcKck59jjHuzl/TVgwjS4faRppd4j6
zla/4xYahrcuRx/eA7/mrxUBJqryFh/hVUmzCUJ8J1lJrSFbuuzfbX6ynWWg
F8N/tJjMOH7W2juo7fnSq/9DGNXR6PQPtcM9PtEgFPp91wvjwq/49PalGR5B
NBpIhdgZ4HooDV5I9YwdTJu+VrOcz/jaBbl6vOZqbr/h1PZjCU5Sx4+Lr53M
EF+FVhO/QFVtmj8dM7XcJhwuDPXzRU7JOK3MpSy+O1a5mmcfxe6VqhLvqaHE
1q1iDNGPgfCVsPvv4ag8F0zT8FolmXp3VOjGWxdzQfps8dQl993HNyOGen3j
QmPYKc1opEQW/STVCdYfxCfZnNLac20DU4HUR49ERlsaJzggWAAByW3Ot0I4
GfSoYMJP4hwwu+meaD9ZagwA24ISIVnO0S9edmoCsBLqVLY3Pskm/KTxdjhc
HZ7L++2Vu1rSNyA4AnIeW3PTTh4gt/+9aUwS+lVugH4QnAUSYmc1KHguM4BB
lP2e91yOyHRJVd+CJXHf5TMk10k1UdqawMVpErTfE2UANAngGwpIIeHAei79
XOqZGxHedab53WOXf9fhYNef0qeqysIJ+UdyoRAZUOU/0InGewrXwWCu+YM7
IFebmdmQyBFvTC34y5xZNJeEZDm+8XOXe6E5HuaWmxfqRT6tqoLMdCaaY5w/
2Vh57KQs5+1YmXyTqzcGBew69QoP3ty9NrpPqVX5B0wOAKdAVRTzX0XOzYCt
XsiCdNNvL6kl17wwFjJGQzyBXFurab7D4cOltC+0pN/+gpAhn0573q3UKN36
eewcupEx+lVzEgzgQUE65CoTGMnhfOGmnK/uVgfEiAwt2WG4KRMo8NoFtGhy
ARcfzzVRLXyv91+UEuWiTVnbaMNYKY7GsPj8PZ3HwqBlIsCuRJAytkQRIraj
ISML7XdFfLBHhK7nD4ENse/icK7xDeIKlPIg6F6eei/demJ2+YvJY6H0rwiv
LNZJdXNLC/qC9DaTjAeXYPlsp5labH2y0K+nrmUfpR32b+i7tQWLW7Gn1bQe
jqGRFDmNVwOIqbQe0qMkjIvNK7a/4HHbwRk1nArha8SrMpBR7fNwObpUtjDX
ILfsY9+sgOchi097oCaVFbeta+9GN9/eWwaYxmtMOhGaMuuGDZLA4kAYLbbT
92cAeWjp7nnbwHRqQtQ5UqN5nl/IFDdWOGMDRSB2KqlmdciKgWnGHaENGR/D
2NjqLUYAOyqP+nO5nnUmrd2Mrz2xjrnJnQzyLAsUVKhTx6byoZ++90GPuTSs
+Q0H5Pf9irfEgRyMtsUee6jBd5tx4F1LfmAswjENM+wCC3pI8EUU8awfRy2S
std5SzYRFSZvEqCkKGow8zsnX9KdkASnADpuuhvrFhJAFIvcCeL73pwFUlym
DN3MPmLHWFNh9rTk+0BezLsVdncMWekkdD/5BNa+dX4CXxEPHKRN29hBS6jF
vJ+IC21HBC8psApIeElPWvv5C+cNpnQBd9JIlhW4zSxEfP3oaMeSsguUYhAq
h3X9OAMSkvVOfYA5880QaSlEhq0+2yQpoTDzZyZOJfXXBrXTBnUaycvVwqRd
71K8Mu6HLIfpXBKdWMq0WYrzAVuHvfdPkHLLgmCYtmBk5AaYSyNKQWHz7fw1
S6dxvz3CqvaT/V1Ba1nqA51DVhoWqJLcqtFbwIRgjq98cxo0ouSpJeA6OYNc
TTxgG+Jm/0eK2IdMaTh6zbHzeIm5Oz2GqPISJ+aJ+HjKPWrIGzZqnK6mVlEI
dDwucb5Iym2GTnDVGeEMmjy4eIep1WuI/1yA7QsmPkpYxxAjIpiTe/0WJMN5
IuOWKE+twIFJi96paU7/npPSNGREiqRmaeqiw/gUAQ5NBmX2uicmFbZyDwiF
kicwOrhkGDvW7iTUtIPQvOgb7WoNMKB4fC1OHTQ7mmHkUY6O94NxIVGUvaft
5hUBSJQ7tLHVF31smD3VxATujC1P3W0oOjUgifTI6C9RonilQMd624WOAvFZ
kGu6kO46sEAPbqq21ZMwSyr0vZYYkuJLeoEa/bFSP/ixjyYX44nNsJQOYh6B
tf4ThJlHqxfPtUUI1/L0qqsGAJukuLCWctgF2jfHC28sVP99FUITT9Akgd73
F3sM7UtwL28MLe5SrtqYccPYkjINKlkkAAGA2dHGP3m1SwGkBG0WMFtkahyD
pRiQxEXYAxNZv+m6V+0oBMY+e8uGrPTBZklEQ95yjYZCMLYGS4/A2JvkfVDc
JK4oeURTawyiR2Wy3vZWfXtYF1DgZLIuzc3C7UG/IxIIGNct6hHnVI7lWJVz
oZ/meSwId9ODhDQICRg7+vwQB6FxSzZb8t5BGmzs37V3t7LWX2fmY6dPjZuM
j65awUHIN/plQkht3NqfTQxyd83T0/Kogs6MUtpa8Tjk6f21ATPmqzq4cEOY
CpZWZy5+GKdHGT/BFwjApNgRT1WVLjK+a6vSY/Knxk2xD6BO7YpGSRDoVvXX
fWs39f1Zw+1LZ7nZzXeR2qoYziNJd4ifSqETJqUZlfwEVd+9j/7l8dJ2vswT
HSsbpH+LLitlG5nIBP8Dfi0j0caRBDZHBMM0oLHVx58lS3Dh1wOs0+ws1PsV
Etcqin6oJmruqKinSMpmSid3ODhREP7gr9gkuBv9eerttgP6QbVEkW+sHScw
hyQV3SiKHpcG7GHXwo3g9f6qzin+arAk8aWSrZV9EpcDrNgWD7Ibt5qshqqP
1CjOYMEbVkQiwvpoWCeRD93rZb1kaGxOgG19xVcUOYSZ6gCzx2fbq21kb7l9
6pY0ELrizhP4PbcjI9HpGjwXq22FRkohqPpOTWTJ0uEdtajKjd+C2f/wazZS
Yn9dfMm9ZAhxvn36D9r4wylA94RitTEA10HCk5TmnR/T/20olA3oDTXOIA4/
S/FvPZbVyaM+HvyVuL2xLt4asPbEXszjK306/rPKYO0meoKevHA/AglMxZXD
os6rEcibepKB6/dfzx3ex2p4cTsl2yH2WyF7+In8nsZpWnNej5y6NpXSAgVF
ps2ICuwAlocwwx6fGlJmo5nVO+evbtAfjzeZZWj822rfw7dozSSSKFzFN+0o
COhlVWBQJbR6n/apl+KjhbqQBCEh7M6IiODtdUDI4hmsScG8zpoQcS0wed3p
j1+MfwYJwxpX6kfkq9xfGdgFOhb99BWOCy4O4e2cjwPKGXp/BGy3JDVcdvcH
Afnm8mVpS154EHgNTMpG23jC34g4Tj7IOy7LtYr3dFn5lcgTus/Hl1yjRF2L
+tfiFELkUrdZAclwgUashA40qwOTc3qZl/HmeagzGOXr27TlXD9gU+9JEMCx
weLPP+zAhNpptzmXGoiZpZmTHHG0NxEHLyjeGI0ujd1dfEFCmqLL2XNTpvhE
xpDWCdUsNTw+QDOVprMnrohx4NGbeM0q4pbINFOnwmR7dOZe3jj+0mZQiCbH
m5LE3VnCPGiySZLPQwxApTusjqzB6QR5jSlaKDGdswyOdJnOUQOkpHXA7gzF
tR/EE+FpoMjAeHOa5Td88XuZR874/NcKKFaavd+4xk6snCDcLutLEmkZwbr0
tHwNTZglscUkN5iN2ueyZztf7XLUHEyxAri48HCthLYouZmxKMpct/ewUSU6
FfKz44U5Zl6v5Lzxd3+wwFBP5DA6gOtkUkJYqEDN95csCt/DGZIpJ28zsljG
/q4CZh/phjQt9wNxyFcLyQC+mQHs7qluGFEz5IHI/ALPfYglRx1z+WWiNmw7
1syp/hauEPE90O4KR5YR8s0ABqrISMIT7nyZ9E+yEUMnhrryyIfI/sBm/IoB
gULSkatDYsHvtV7tvYFWVN4PW2SfwQT6yxwD307pFbvs4sLGygwDPKYAqHXe
1YvpkObvFuEuZzfHt9QGa629HDlfY6ciKWQXZMRyFbbjDGiURPYiE7kxct9Z
/KxkaLnryQgRQkBM5vCrqYOh6KPuXyUIBeeyU8fOjdx+T/VOYGWZ+a9xo68S
y2d9nrPsRjTPQfwQCKS4XMAcCEB3Nq8d4hiqSmAVNlpjhgkdVQADS0Wq8Nsz
rK5Bf9+WdjQIaNBT5JYVk80Cd4FbC/1stgMchOS7N82IFGbakVgPv6y2r3pb
l3Ka/JRECAcNBV6OwN7GJr+DiOfLWlyMcI19SOW/Y7reaDS9TSiTsLkmjAtc
cx7iUJC2vvIA9L+3dqrvDwhfvggytAAgqOKcmm4xE0GGN2/pjGL4aX9K4JAj
RisrTvceXZg4nFlYCmdGNU6YncH0trXrwmRlpYb5tOeW7qWWI0VDZQf9q2AW
nJdO0uJH60/tWLX7pOiXCbfp1IaOMkjjVzceaMtePa8UjfoorImnAhWNA/UM
XjJAL6kbNXiRXrxuHOGhNebx7VcYFFeNk3M7W15W2ZBpXPQ6aVltW5IGE8rj
DKasiyaLT3Am0+9w0ALzEDJohujl1b6bVeUl4T33t2DLf+FsItVCjuEhA1Zy
x41o9fb0P4bBuBlQ/cgvSKHrWMeIWuhVNQ15ykaNV6gdSQewDBJ045fK0rDw
mLJfmAx64fuFDIrO7jE0k3g1btul/SqbuumcXFltR9vtOlmmgFth0C3M3R2S
ieAGFBm8d6fRwhvihkXQc6SLbmoKHRymBaEUaJEnbUap0qWhja6SHhR211Ks
7XvMgLxAUlbS06PAsfxn9TQhFgVtpJaj5mHcQeoQvrm2wWXwhe3O53LMMZvq
iLDgJlcoqUvyA11xlblk51o0UwZyirsgsy/i0KnV4lkbpnQ12HSm4RCRzeKG
3Rou+EST64bJoRlQfuiazbswXHPJChZWycqNMXDvmOCwLzsEZ7WwNS/eq5Qa
LFsbsfAjT6v+AF2q1FXIQIN+QTIlNF1bxZCJauGsoB5YU0YEvaKF7cO8lCV5
CxDHByEG11rh8Yul3TdJGsOxuVvNz+iEIbRm6POdYYL1JHX1+zGD4LwL+qeh
6tMtH0t8yHfC76Fr73XFoKeLnt2sl+hXwdGhv2Q7yd49YkuzW/anVC5jr2IG
SESpxL4bxHmnXeplt3HPn0jZjM+uECRkX1DNR5W2CVSZScGW56OFMViT7xW4
BG3J+RScDBueifQ0WL0F15nUuHsyRAuy+0CgS/JHglpWNwTyBy/cmrtE/Vs7
3WEkumWMOIfLz1Kz2zpetUk+N0EwxvEkW9Q9O0vu2luam2ZH40gltQTSNJRu
nx7/XuPHbzNrmro0yno+Bklq09ufhS8xiOUjRA/40b7tmxCHmpfqJnFNmBeV
xzVrM0W+j15XDMU8bibfdZ49z1Nd8KOW+bSK/Lphkks8QmJyEwatXlQlH9RS
FOxDvcg5dCOQXI2505y7iHu6jd7VpJivE0ZcWKgpFh2Acn6FHAthYx9XfiDd
DyHY91ZB3YYe844Vp4yg9Y6MZsgywadznqh8Kj2mJhKorYVENqDxkcPSduLE
78QQ6vp7QKqSQ2LGZfOA1kOtZHAU9/k0ZAIBW5weZcHDnY7nnAWxjQwmJX9a
ajM23KFCVlSdBxOgvEr4tNubktBAkXH+2xqE2hASuBq0S6/bL+QWJTJ5ye1H
mLfh/4wcKkxh3TWL0CUhztYyZGkpYHfn5X2u5RB+re3qF3oaHk9091nC+QXF
DtdVymk+rkGoW60lhSnucXnV5iIufT0vP9Rg6rNW0wuhJ107FCmHk5GfiULC
q+k9rDCtHiJK/7GDJszgLS7ZE0TMJKWfrb/UKN1cYvrKINq/MBjsad8yIDdo
bGk87KiT5JbZ2iWHwfUBO03wwu8z4k99Ec6V1+GGFn4WxqGJ7yJ4C2PnVv0v
brvXpdK+PftBRGqKvDBL8fU9+kxqSiMwJ4ecBls9sOH8ihQh+xjMPCzBISPo
BY82Y8NW9VilkpPhR6HvUQAxd3Py4JOlAstpgkURYJ/URSBPjVSOh4qigC24
3r9V8BMOsfmVu1Epc7hHcoCXWPo4AkMwbgcmLV5C7gq7K0Vma9nShSx9i7Ix
S8wPufdrgsvuU+rSxdzKjulsOgmPQ60vJ13RLPaLT3O6UiB3Dvq2+8AcxIzM
P0A275YW8RZkcGMy3Km4rif51thQCEBYSrcMlcXveRlxEUoyLfZJqAej2c2Y
r2K4e3xylyv6xgL3It8IzwAGbnWrH7P5G3y/9b9xRMgSu0Fbrcuy7lypJYdK
0DwUbZf482gMHts3V0IJXbBFqfR63r+UH1LDEXvy3h7iGFlbHHrclmv7aQ9J
TrRzGb5vQ/CumZcfuhmOeZNa0qkybo/7AFuScw3YogVUx6OV2eBqpfKRGJ62
bB097YoEAOmjL7lC9adzcY7gjq0RSsFldEKPaQPbrrTvpSyVA0UiJwGMo11Y
lrY2dzQGsmCJ5jR8bhQ3ezcJYMwBhqJqytck7f6MICksyneIpnLez0zJDuaa
dz6dg/1yaBECXjtIk3oiN/2uO0JNMx8OeuUcjrGXfpX6/Iqfog3di+FQLran
3vcgxBczGZF4QGz9et4QhpktLmeROKgOqInFc1eAK1Ab5coYCPVjZDLJnmkn
Zv0vQWGOkKX1FJVIhHNIr28XzIPbDUBzKmtq16qPbJo2mbYg3DZni82ptMAI
4kDSp+Y5V2BHx7/c32YVDafWapUpvcobuR/gFnDWvZiNB10oHvA5bE+Bdea6
D7scflG0UbKqmowA8/Vn9M6hxaQZe3tWdkqRsoAiuOtunrvUSwPYos/02y48
KEqV57qoz80Wo5dM/emILPXp1Q9quvsFMbzJO8IRbYs1g8Bj+TT25oJmYbwM
ytfjLcQ5zncWs53Wf4YB6qVcWvtb3iUQOdAq4LmqVqQYRiKdvQdE6agO/IVZ
yJ2FBIg9u5egcOaZlb+TWYUkIiMFOQNEBV7UtG0AguXiKEy9bU/Vi2Bkm3Vh
bRbMLLx8BxrcGnk19Kljh4piEGedkCuK3NxUahGwT3Crq94DFdAwLyk3msbc
CGr2XHvi4hrfqglYAm55cMSh4PvNLoEV8oTn0mZZG2Wjig1q3oPBtZuiMja/
oEsJs2Ps9l4SkE+/HDqijlw5JImePYVKOeeNGk3N7m9S943DyVAfGQ1svGic
26Ykwvo03ba251cEIdKyf1GWEgSeSaoqIKqvUk5g94Jmm6WP6wUmc/mlGLxS
yMppuyu3UuXkXl+Xt3aUYYpYnJJdR0onRAzGlSJR2OHEey5jsjDW8YSAKsrQ
geCO/VA2ajCK9m9nLoWahpFvfaTwlvhL9CF0u+J6Dg4tfv60pjMoYEgN/zjW
r6VpclcJGnY2gRjD5Mv/BGegKigB9AgT/VxIjhQg/PEGMwNupy43lqHxnJza
DB/PGYa7yYx/UsoK+BNgKZQ7BUT/OMHZrHFzp3gcM37eLYboxyM92nrNmN4f
NOF3xYZYOQxazz1J25YCSk8Ls06dSd9YIb92gqHgifbeVabuGIfXdj0gaM19
wNs5mSwrY39potguaJkn6IRZG3JQNMZxS4LxF9zXzFHfQx9ik0sUmIQkgMQq
NeYRVoLDn4e+vEHNgJ34vvvlyG5r+EvtYsxYGTPB2EKY5KQ/mb3L7lFx3jr+
I2U5jMD088pUchtCms0Y2suVJkn7mzcfd7iD9RGzPeinApiIqgdehR9zwQD7
c0kOzJTT9d6ZzhE+zvXNnVeLpnL2XYlPNyoAST9kHjbGPr2k2xdzmgMkMolp
0plFhtjG44mgrAdRPI7KTVNCBGvyLpZo3j7nhWOfPJSsopGGL+BHFkxlIYjX
UJL6HhUQe1cN/EH2QqQDUl252gj82PG2fV8Kdonrwa1xEH0xHqNLN9hkEEto
+KUJTxYX3Jpu7TpKLGGdswizqKtnBQTLRdwE8118RZ7U2FEdlLv0BQNMqBti
Vu0E4uCSeeplEpwrNflW3hyg7ymmfU72LPz1ClXDqXGzSt43zom3hdbftD/F
u1O4xzNsfBkxS1V5k2dQKJlFIJCSHjr1bFkPpkPL45tw63orIW6vK6MPCEsX
bR4jnig59RrQ4F35Qo5APySxV0bwBlPfKxauWvKiW/WSobEbwQ7HTyhbfp55
d6QoEIj+uCrfpug7FpP4vEkyCihvhdstjFg0N7lHN35aMfX8Lpk/8SEGXo6a
/8RWK0S9ylrYmU7PELW0PwZFE14i+tBMR4SttxCMuuKkKOYkJw9a0VyTW8eT
Si/WX1rE0DT918dJ84yV9388ST2JJ2T/Wl0F5Ts8mH+4yrLoAz17anhgb7nG
Mc7a9c9FF/GmtAQvx8aHHAE1k9u63aEG0nva8whJJmDqvrQmAi4UauV3QjAE
LCJCyoxUf2hJSKMBIXfkemCuXK6g0bzuZSx1H2PI2MPgHZ2/fa3DMafg6GKI
ufE=

`pragma protect end_protected
