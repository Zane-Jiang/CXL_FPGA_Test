// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kixM4mLgFaTPyYQicxjZJKaLkn4IQWJG5PlI2xjnvnrWmcNK64JU0ElOhWuk
c1HfAlAbQbrp3pUB1hQ21h98C9CNdT75IsXGyQ2I5NVbtbX/8d2y0jfJJNdn
1i4uCuDDQJ3jPAEsHuoFQR+D3Ry851+KoaAV+Xd8V3ulcAii3s19NTsY/JaF
iLTOEasQUROOjIiSgA8zce1GCyckNVIn1heRQunHJTBKas28objyaRctxtB0
a/px8b01MyAb5kk6q+Kv1qvIFDY31UDqeAvQ5zBTAvgp27qHEBxny53J9wee
vmMHxV+9V1GFtt2pvb/f9xgKw/7IUlo10u19Nna2cg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aJyN5YdsKBA+eX8C7FObU5MtMhSICffe/02c4OpXOg8p0suiy7R/uw8+/uMI
YRJfvUedVv9SBav+hBJHwesagMn8tXZsFZ4Ugcqj+cSnRdCYHCar+4x3OUl+
+zyRBA9boVM74l17JKAeBusTHoKS3AgzEl/6pUAa0frp/6+pMLy1M8i6zdSq
1GIg0AcJBAHjWvH5644iDRrUBjpO6BAw3h5kzO+vhVYe4WQHvwSC9s/QEu7J
M/H7okmsFxBzyQMTGWpEFmHb5UilIYogCBOCvxdO7jmNdDog47hZHVG2l/Ay
GkeQfOVHIDIa/D/qAUsccqGg435T7djjNZetEbq2jg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YPi5CisH9TmlkP+LtwusUb5DU8jjiX+K6dPNkNc5B/apZYRY4M87TObGoqMx
sk3dGsdr7ztutnRiSTbAXLUG6ZIGCayFSk9z17noFZygPHhMe3A1DyEi1dTv
zl6nAPlt6Z2bNM088KbORiT6e6t3vObCIgLwOh822zI0SsxPDj64RJNsK/hi
CVJHZJSDWyI1sq0zhUirMHAW65jAJlwM88JVk3Mh/lpZv6TpPTEFsEoBLlWS
L8bJo2kYGZM1xtLVi25ovIxFiuylfZOPtRKEPHh2joTOyt5Wf5sfxmfcjjG6
t5aeR9+4z6NW+6nr3XeiiYPBsuLik4nv0m0A+sNDdg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SFV0K6XqD0zHtIkGNraLlg813vRUl8zm1+qZgajS2Jm9vFmR2PCyW6PdU0I1
AhuoJEjkgs6+K6Ys0LG8x1f7e0BmVdWOO+adwWJj3Jn9Cgo2TIG2hytUl2CG
qJjvxOqrSZp4hpBimBDKnWo+59xl6GxmsRjapgM3S0X0F1hytc4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
u/jeLRMds2QeIE0Mk/WU+ZeYogUf6MJq8DXQffkTUhakbnA5THdE5vwQDmEV
m7QkhcLoQD9MJAEtc4BgpCNwKaADWzgJdA6xncmadmbSaN5Z/7LjvHVf0Z9E
kliGXU5R8qxRaIat+dHcB6RDN5Eic3XH3GXpPZWczvSIQ2kuSF8WunCCnbTx
rOSO+GDm4uhx+MxXynEp3vxq04NKf3uVmSGdzDCYjI4d+A7rrZ9Vgq98kMZ0
z+FnmQmo5oQfAno1C0RvlAc0RVdkfGeOKDWyu4BML8n1eXQaANBFxvmCgeT2
r91n2vyQSHUrUd7LmJ4XIS71HUJ1xZGhe/hqp3fzEi6Uh4HjQ/m1MwxKbifR
MI/xxPG7MfihxpqlKWiAssULBz4DYLuXdilQHzd35nCjecztWJ2M6igueSRB
0ovn0Tlosgr3aDBflDTAgcvLhyTpzkzDf4iNOPvaWL8ZXD/z6r/duEs13jYC
iWGExV20dKzF7gj61FA6JLiHHwtDdYcO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WcE+u/W+NzGmStibDX5/xFdFthx9IjidvEjBBTKcsA/NscUJmQ0QXgrNNWBT
Gq5gPlbRzslAy6pJJm7fst8iKIucMVu5TjhuB9Z8Y/sQLo2OqyH3LrG8NJSe
eg4qRmnQmFdKDgbDc38NmhbVno7jsG0ozfagiLK7TqLHu0Ozgfg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jS8DLszB5iCFjRm6VmkSEv/kPy6kzIWS/yQzLS2NprT2Po/gahgXEo9pCc+x
/2vN8FU4a/nWToc/vBxEobT19y+/tCXGfvGoA69tqJhE9HocMaACDjVCNh9Q
DEUlPgtw1/YNgoaZ3/Vr2NLic9n7NuY84TIJfBq4gkUe94IWp6g=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1344)
`pragma protect data_block
pPJJKLt0Qc4T6+yNM/yVELyZzKqJXCOtSA7l30ndR5E4RrMmS89V8XY849rH
ospu3qC5oJ8P1GOFAYcQsVAALF3Bg0HZrELpAV6ZT0KABBQMuB9tChi92d29
Mp0RLVnKxeW2QxJTl+ElNxAmuNOEDu0KmkSwzrv0cooJD2rtgiAWjOSKLIRK
bL5j7k7wBIPdIdfu9JUU+5RT8ySVXMk/UEhm7KsmpGpSCihJ2OvHxf139i/E
xiXxgZ2ScO0XsmWNZ+KDJaqjmvrrXFRXtVhVkDTyX4kF0cmyFnQwKxjkz/an
qM7RnkYCIllfq3G4sZkimIAPRHDt2vc1jr6IluQZcHDn8n4vKApj2fv2wHOb
Ysc60PmZhJesleTQCF5McmVHkYAW2gjkpXwu3DoG8bSWyNN2HqyuEcndoX0k
MZLYB3MC1RdcPqEI8Sex+E/iZQYH3wtdoEIuqgEulJ3QcT4oLQdvp573YiyS
FX0RXNcclVjIba4jmR7aMFJj5fWd9Ik4xDV3w/iBjsAi1DpDbQaY4psUX0Ja
Q3AOrlUahy+dVbik2rcOJ35h62kqj1xZHAULitheHXjOWOT0eUEy2qXx7sWU
c84aAV/Uk/VYckeVuiCMVH+3+wgdWqgCF1rWbJHyyILTp8iBEU4WJWniMVLk
WeP077oRgAwU9b1Kr6v2/BZUdAinOZb07/v2sEYrr3FGqM8ahHunNmOKv5bp
xeXbD5sJ/lWYkEQYidA9FoQNSnAfl4BCWXYj7G1w1N7boY07sdmgXh5nTH23
7vBVHLRdDq4svnHjStlGb3Tc+S2H/DvqZy9VCFhSrIwHpnyyxTJxqNGocMh9
OhHcbjV5XUaL5wbw/lmjiyJVKlBbsGDVdGcPZ2eDW1+2l1u/sMIP1ZbW9x99
VGKeXfSIVNOUxwSM+Y2Mz3h/p/0PHm1LgKglCru0NQccXl1gha5k8ASvtYeV
9RSmdbPg7MV0mkAkt6QsPOfKvm+AaZht34ni2zhsz8cBLAOCFSC6qJ+e+H/T
HAlZrzzzzEY4xvz5NXvGwT+L5WcsPB2jU318BJNipRy0dAofzt6aNxEjPQjF
8MLiWYZ1r6/0Py0QymraHqv/ga7xTwn+eDwxiRd0AvYoXAVR362kMkKScOp5
gngFG7aNlKpEdZIgxrpONPmi+xTpnbwkudeXpb3AZadW2Shi2fKC3bJKffB0
SBb12xN3J2RUlgwn0K+Nm9kv0j4KD5tLtLfwVnoWPE3cetmtXPNtb3pug4NP
GM2AEachs249D6IJiDihVm2jU3Mpiwa/61qkU6ytwG0r2J23J4FLykBBIago
5f6APyhbgcQyFfykdQEGsRwcfwRIpCNPVEGaO8OcVm5yHHELgpQT5ueU47nJ
gOsf0A2T90HGKeikm9jGjb2Zxml5H3s3ILUgkJJHinqirBHz3ZeLdOZ1SjPM
+Ehxs6aB8gbq0j8SpVWX6r2gXQM0c8XfcQKdTCjEEr/rtvmPTsW8FfC+qkhm
goRaj6TDNW4NP57Xc76H5CEBkIbNMFOGIeBlcqMk/iajpSYOq2AVT+DxukgC
t74Um0KnSzS/R40t6ctZpe4ElepwbO5CkNq+LphCul8bkbZxIAaPopdoxl5Z
EC5ZxmL/ajmQDI7dQ0z6O55KnIWWNBE5xKhG/j0NQEG9Kzyaorqz4UqVGeA1
rhbE/lLap1YVHUnL2jTofw41ljNU77Cs5yPK70A3NK3X/yq7SlkMRxXK8Jo4
BuuMobO4PtRe2PErtZD606pGrf9Wkv3Yz5TQ1kQzwGIqEnkyFcuP

`pragma protect end_protected
