// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
f/2s+fN9Ly0cNfhEoNJT37SZoRrLiPuFWGZjZpkrAWQao47LZoM2z+ez+rgf
TgYWC9xPqD5HeiPnk+J73eMAlig63TB56wRQE0AD7cJlabeZPc57w3fP1ca6
Y+vKtueIdf8hRxwOoBP9HOKOKoeqV/53LdzhM8bYxKY0bzuyxh9pNAPPoCxC
1FgPufXtb3ba9cQAg7SQGMbSivposfD5yDk9k+6MSMgTvIq4MPTCfz2FACcq
XieNByAdz1l4dnpOL/M7XnHqhoWMqLo9K2zvR0s9MOeC0jF3bfijkU80wBdW
yUrMprMX3efY+Sji9YSTciuFs3n0ibPIDgVtg66+HQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N3onFo4hdI/+6M76TGs068Ap80Qg/U7wO9DCs/XBiWUoF9bnWpvJkFXsyimO
vOggrZcCKYMPag9Pz+VDB6dbf8p+4zxf9yAAKJRhgSc7sOK9/K4TsrS8ia5J
eQiTwDTq7SCcU/ZTrCX22IjyWRya5JNhspWFpedOeWsmYfw2O1Q68f/N0Qfc
f/ROOvnnbj/x2lEOazqeX1zQaIkmM4V/yj95TnovWo5qzPHI82aW/o971Fl5
PcrSjCjrVhPis+Mva25JcvCAtuIMfRBuwN6ZNXo3leoWFS7MmpuVCd9cDiOc
wilsLUoKadH1uE+D+ksTGIbegTAogyX6JRMqkurbMQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H7VVtBcPSG0GCEgfretAuQoUWGbR0B9WkUtgbNCaZGobuRnnHYVIdOABq+3v
vBmb62GpX8qqi5kLdSbIqFuDD2F+fkHY+hAH2vfEZlqu2ILfbKVye3uZ8x6P
u/Alr0qxWN2qO8aGRaGCYrlkfxjmNNKLscThEKNIviyLClzJuWzWg7Lazs0J
MDMTCSl6KhfbZEssqFfNk8tRq2PGNbGWvjBwIaLMa6Nivvyq2SJl6D6Hgdsa
4tWHwceSetmPK7F1cQIrzbYIoYQkLqQqy9wQV8MiWbIQ11t6iB3mPg2RtbuH
1qlBRusMaeI5DOx41xNFyX2+fULINnzYWxMyowLseQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BEQKUYEO1DncJb+jwk3WN2S0JcNV1QoRTxhsaFR+zmHQx7V4f79hdX98/w6H
N+5bBYm5ndDLWfdvAgdIjM30vxO5h3j29kEzQouiD1M1rrTVJKopsTRbAM5n
nYyA0MH3nHQ3yrSDHMbLocVDADSkTYk7CUC5Uf4y3HL866ISrAk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
vzsv6RR146MAi/NktcRU8V/6KRuY9bBrR9zMETc9IYn2ppjn94PY1jCUgOpr
E47M65CyoHgQo73NZSowqmcFk+nzAiWSDUH6qxKP/Uc/RiM98DYIZVC3Sez1
RsiW0rY7CANpTKu1KTQAEBT7AYTrjXl6yqJaLQdUlaBrwRq8+jEmRhIRNJeG
7iziMyIykhvmCIb5y/H9KEfziWRQgr0mf6qoK9egKnOi9rpieeS8f5KKxwEu
0cmHQS0y6I06SKBdXKkErx7m10pl80PWXasFNc2aJqlJfgZbctFVE6Lueqqh
E7eYXe8dyUtZTu7F+o+3fH77Ypwa0+Ik3iUsigrOPUTgiwlZSFk2gZfC8y9L
ny39idK6WjWYjyfhx9yw321FDfbVcjBYutgNcl/a/bewTECX1dfcaGYyWtPk
MiHfulhpj/nxES0/PZIQsYFsdCfd00rZQws0W9ePEAVMkwAZ28/QV47lZ8dx
DuTdzxHRuXa8iPuyWJJf8gHldmPio8Pl


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ag3/acIM/i/EaiAmzUpPGIWZFJwicp73GxvearTTKZi8uD5qhjZaL+8VexO1
R5mIm0w0Dy8E2anZ3cvqhhuI5LoXrAF3WhC5KnKVCYn3jLOpH9OTd2pgiWMR
PcKm+pGkTPpFSjphS6/Wp32soEWg/T+l3bgwieXOeSYudehMh8w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ewbpqoLpfRJIX+uvmT+ukb0VPuyLG+zaNi3pC7TZY531ATPQwvCs2c/UKgNp
DRbfVsOeltRFAcHXcrfbRUAQ6ENl2JKd/1TxR7x50z+ttjSzBrh16PdrXlgw
05L4WpgbvYbIVXO6D0xRRMUJUQBfVRGZ7uo9GVLbMWGibz7yxSw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 281168)
`pragma protect data_block
mk+1PCB0wri+oE/1fzkW9XSXmp15TE3v9x3gXMkVveTGf0K/yVo2ZXReQ0ZC
nOaEU7cJlsMhf8vyCO1FEHkj1kyn03kpdt1xykXguUtXVu4QxH9od003xO0l
FKcjcTI+AFJ3eBAjEyrR1lrXUFl7V2uKQDZIohQx4DuYIzYyaeGNy3FKQtjw
6+F8vcPYunxQFwT5wdY45Ca8K88T0/cltaQYll4UQ6BrPDLjqZPW/ix9qGi8
7AJ/c72Y2nzde3zFVc6bJ7ReVy4rlHtWZy+GL9sYNsDShuqDNUfCqynO0O+N
Pexwx+qBZGWRjDJv+k1ziCidsWXP95Es1G8puxjj8417ZU5mD+XEJONFNrTg
1KFy6zeqAKW5I8bPMs7jxbm9u60L86DbNHFfhFEbSl0a8ldwNxayKxSodrxl
V2G46mAlNJ2s7EGBAdUcuuN2aphAuyVIpc+ZC2p7lm3ol4QlnQyxSdaJz3aN
fH3EWOusR+tsTHqqsY1iOiqbxz7YCsTq7gtbsw8CLUWnGjuMGiO8EONzdOXG
52uOl0OXhBQKGxD6A/rxhuV5zdkwYg75bVDOd3noxAPeWULvaejFvmTgykOI
jJe4GkWD81mk0BNJ9g26Cwe/if6cFLxFZ0tmdtezexeLTEY5Zjb57BwznM89
H/m87CR+Xedfj+l3sUJSKNLT09xK8DoihMST6UjPg1gJvwF95mI41I0sJoe9
rSQ0DLF5CttKqJk+E1O45QK4ANZBxuEr4l+KgBE5BsMStIFOCeJyHaPGXPRR
n0qjA1nfd+zUwdTg5Xc+O0HX5X0CDhsr7XGd/iAhqX7LRFVYOAcQNs+gG0mZ
bgiJ0ozhtvNVjOTRVCVhGCzMIWFTk0Va5l0+mdWT+lJzp/dJyT9zAkpSTBYX
XeSMVEltM3i0VCHrti0C5e6rOoyVlH4w7KOMuHmvtXbyPnKdgLc8Dh1I8Kuu
NvwZLSdmftQyGipX61T3WTrTGAe0kRbNGDbxHEib0D61DWsKHgr0ZMKSjMJv
vQr5wrm7BqVS5S1eR75miU6K/C/nX28wypyi0r1ZO9UY/CfAfFDsn6DoszGi
JzW/yl00aJK5yO6tow2cGqTMyUseOIaem+67X2wqIeIzpDipCyCYGf1dPnxX
1aNhzn14WkiPXC40zDDGdYZZifQrcbxBEGBG9iwhtmX0pDfRfDryKxCtCeP6
kG7vdve1MC4zRZtPaH1QCptMhuIyWvOjnSlldW3ls6am9gFIX34qwAyuWO02
MmAWTeqHbMdL4X5mtBUjgglU9pLaEi7IMGVsGGh0WTl8xzzFjZSAxyyWm2qQ
6grWnPCbPm0mrhd0EONJJXuZtiSV3mW3IBb56WVhlmFXkDj+sREIcN/db45u
ZA+QxDkVZ+TXrxbDoMn4nkh1qqWBe6YEmj/BuvYsG8rCBhV0qCb7nS9khgNS
tmJkHBd64/Fldle2l2r3yu5UwAfLtk+m9cV6EFpxW46dkqlCPyfho/ltdKJ5
lZuZeB7ETAq8dyJ2qtpT0A/B/kyB7cjG2GVpkk1Ig8JQMrX3rs4JhT9IKwcd
hp78iLtPW8AklZu8vzzW4X1IGQsm+izSWWR1CyRq/Nf7hYycdX+LMWsKwVK9
kPGdNvnDgR/XqUldlXeK4/f9FRtgB8yEFfzxbhHcQTmLKI+JlgN78c2APhVX
htTn5EGk4fd0KEKoaAOTKN86BDKSVADuRKr+30njnxA2TkQ78VSSAp2VHy7U
qNAi7CMs2VO9T5JAp+MoR3IiXwjdgw9XeuzhirJSobcbB7C4vuj+T+02F9uh
XKq40mJVQ/G1ieP0ToWau7K3R82q0z7vaXMITWSoBuG9onsR8rxXunWJz89N
jx3O377j33xelYcZz3djS8YnU6pX9BGaNE6PwhUs2b03zWurC2ajseWrdHFx
cu9x+mJPoPAaVr9eym7tsOKfwQViQjeVclV4EVgD5QuX/XWH+JYU1FjKY6yM
pQaq152C8IkIUjUdIXYSscpdVjwDkA3MHqHk5N/HENII6ev/CbMx1MX9tikg
xcPRj6Fqd3QZ8elx1ia/VhdC1zdRhbyOd55xNxkZltKZ3TMecgR5XNriWuLr
5vw968uR16ot3B5lLIxm0riOGd9d4WksOxJQoELqELDI7SIo3yCniLewBGi1
JnXVVAulzQA8QxegQx3a5GSp6PTBcZCCrPrnuz940gRWpq1Gh2oT0KXX6tJ4
juX2yTM/uZ+p1kT93bpssY9WkgOA+yPgO/zOocvLV/u9xY3gP7K9VglJdQxa
QQBV38xBeJ7vWwGmVYmnLmGhIfNi0Au50pZpzd2VpXh9vGXyn/LcPnEGmBgX
8s83G2fKIOETRqmPA2DYL5zmG5HUVaZ6hhFZZ5FBtOxFJkOEs79KnCxeabpq
IGctOl5XlpJd1No/8oISzBCOdO9dxT54dDJXVM3Rs/AFCzZQqizKtu9E/fuL
yx7h4+xbeab5mW04t+6SxnlmVEZuGs412JMv0/5sPcFXTO0En6D8SrKoZtrY
Me8Zu25+GHb3wC0nLokTMSCG7o7TRJ4joC/3dJFL95udkbTap/zx3lP8rTqX
DKr6MAvwfcgtaBrwtig+9W0fOrausjkgHrFei1dSi5FAIDDMzRX7ELvSwEtH
N0kt5KIRlaxM97fHmIl5SPbLBl3izhMxCvrsQJt6M3igEjEhfqFw/K6Svqt8
XBFCs5rKegXIyhqo16BJ70NHamqJjTWqulBU6jQc4qQ+5wMzGtaCJr/V2rSP
/cX40GPunu43PEibB24f4RgxV57j/QDHfNToWohP5Kagtj7+qaT+C2UjrRSH
ZWh+JgvyHGQwjle1luiRISoVVFT0/2GV73z7Svsvl96Tul2EsJVw0ubezEsv
TeWGnyxZMZgyEQhSPI6E5+63xD1BrGHz9h0RbpeIuqw3PPptfZ7Xe+/YfU8D
rBP3ZFXt/xF4coZ1SiQY14NIiA9dVW+8cWiZocHztcXnvkiV4UWQBXXiGi22
Le+iKOob8DVpkXcMNuYFpBqPfLbwHT39VZhGVUXGS8odAT2zxvovBmTU7Dgf
DT07rD2CxWlWGi88PEM5XVRM3TnZXxeD0eFsXSQFdjKHHZNX8RVW8G5X3QQ5
zmUvPtqfSdZobmuC/CwH3+67jbQU6zm+ABMcYV0y3zssN6Mj0CTYA8VE4hgm
VcAYXR831qEpwpw54jc16W6SHS/vP7H0x1ZQR9eT20Uh6wdppiu9j7btM4JX
8PpT/ctbH6eHevDxanQQgXkuAp3XHC8xKM7i4ivL60NtWjWIxy5TVSOcfgcA
qjZto30PrBMeyXxFhltU0CE3F4OwIwE9CTHS6adsuD/J+fR0/S5hnh/2ICNV
mfbAdHugonpvu9kT4AkOmCJh+RfFbjh/mP+DXrZuy6b8yZ7zTOX1OxmKFKG5
HnYNyCAHp07sY+tqRcANCqigbeiyNe+mqsz+JVpwL6T7UvNsImsVjuyRvmIr
aJ7To23NP6LL7RVfDaGyLZsCF6CVxQ+CuuoPUSqFMUOqdTQisW6kpAeM3tjk
bNMTnwn0yeyPCm4pO9yenSZNlF9Q9hOxaPFamC7xfSiTZ4G0vA7Bpb9C/Pvg
jI5wuwID37HxQH7y9s5XeAcwzIpzx+rcCWrCtYZUAeptGuZOXC7NcTf/j1GB
rIei0b4BolCe3oH08CXp9q/5DuAh44QLKQUz2iul5XLffwLtbzZXKbo6bMQH
urEZ3m3OHvXP1WuxPXmV48+mIE6oeIXwLWlvFQG+xD6ar+7GOGGhI2yw2BcQ
DZOCFlCNc7S6Je6fqAdDODNxWh52vc6FSIfpGmVfZb3zOHxPn3DYr49yoTdT
S2sdLIbbmGYXUuu53zVUMI9K8yzWWjN4x6cmHeWF4ik+cGmgP8KLkl7oblW8
gvKo2OtNVLDkbVPZ/SAkQgQ1gbk7qfyvpWzQDo4xAgLKnMSPo+q2MLPyR7q9
B/22odCGJeLjp1BghGKf5lgQ9PQH7mXLysC+jepEc3e6ak12K9q8vdN7hWYj
KYwMXhThoRtfMfx5Caopbzbrnv1MczSLvUK1QpMThcW34RGK/exXnfc0fanh
QcahrvlobXUbCxH6B4rrO36e8zp/oqf9IW6Nnck3mIgbxJoRBFFFBiZ/8Vhj
K0AlWB7n+26Zy3HiP2cJX5iBu5UgFLj1LUMTqJZWpkaGx7XN4jHnDDlLCBit
TvQZpaF1QE4q/LpSsK/ptJqx7gNLdZjKAoPJNVwuak/Oop//OMSyt7SmuQ7q
L1VrriQYd4E7F7WrI4Sa1LRSjw10bMgzd1yS7hl944FSxIi519b+Z4KyWOvH
Q1NhDFeI/WAwb1d6NHxOVlZ54Ft0Exk7W0fEk08N1sdoCOivUgtIa3VUnSCW
l6J4czc0rKVEU/wt0Aa3SJrvrgQBMmgbfl7HmLUoFvlTSS1sf/QaQ6MZ0zsd
6M9WXaLe6UiIjti3WeC/OP8jo+S7CXHh96ly1Py+PNeJ9k47QCa1kbIdCcBJ
VBflfwlydFwrQ4OKLiZVKcCUTc2UDCQpKx35oHWfi3GCiCRnpFi1kmEwoZ1D
x6HT805/F2H5RoVhkKm50mhFHKbU/gw/pWDQqHDClFQ/vuZzkLKPnOSK8KHo
FuWuZ46aXWn4VbqicWuTa8VGMqZ3vJVxiYkMzWpdJer+JY9HzkHthZriRE3P
90eXPl7+F32g1LIiJKG2sElck3h04LTDjn2vPqenHuW/dCmD9UrWb+62S+oX
GoILYBvgCuqPlbRKQPFi8l/zyaCMiqpuQ92kImuvzv/rWGy5c5ELmhY7zccm
9aqOXcr1axUSTzQNE552Q/o3IP/Rw22QUd1XsM0n/d5aKfff+jRbdKsaIo4+
0DK7R6Yzft+FqkYnG2vOFcwFUt+lUlQxUAd/oBAKG0epB8MgjFkLtU+e5z4y
9sn7tfsFEokNMno6RooZ2x99ighIH1TH7urWUy+evnw6wUigQ2t4n3riKmIK
aFOJ1QNhzUpfiAdS28t1yg5vLJBx3xHaaf+tjWWp5HkK4Tn+Ra5hekzV4EDG
WwiKn9xCIvXhFPSmBBK0V2nwiL1cfrl+XWvQ135Ak9EqqlH6dqFMJsgwuoGT
F/3Z1JBV/y0S5cFD2gvO0anxSDxSw1+G5AvnaVcYHvUCef8glf6LeRt66pNM
JjGNZN10yp7rah4XHk1ui1g66eh06ePK8LkOAiUQY5OllyYesyfjU9dFaKG4
J5sbwtmfJLx7Xwn4n1rP2OAf1nLEJxzvwBvIJugzSNey549uHpVt6KI5cRDj
PKZnujWG1gI59z3j9UB/WduRfMPQMS2l2bbCKrvMXRqrAs+RHJcv506pBB0l
uKVFMGyC1uVWhb823rBWZYctvH8htOEIATMNFkE2ST/EoLwmFpzUHoByBYkW
EsU6Ki7lYvw72akgakligGnSNnRyyojVOjZAgrdSuMbZpSOO41a7Dh4Z1ttD
q13LaI+kAqSDDlhJYxUDkSu72Ug2aCNCwDrsc+zVOhAQUEZo5pD2xiRrZshB
SvQkM/UzEoySkYFHRfsDjZHaXzgt8ZMx6xftG2Is9KyIQMDLZ/J1NLCUwAcK
Lqu3Rw+TX9Ia1re5aCJOg3U110bA6utB/fVcRFaQgf7dPc5fE625JoLK+QeK
ENEZKUCF658SlQwIMvf3ONyOCByaVy6o/dDfWEK0hLpIbHm+wAlPIasFWKPq
sHdS+R63yGeAPhnzDzde8PER6Xu3/uiHyool+qVyAoVZ4ILpAVLMcoTMYbIZ
Ut8XFn9dQvauRb65Br9FoGZk51aYuPE8+eN7W/JXsimFDuqRTTbKXBzmxRUK
3NykBLLqgFAe0jLkzW4aEPCSyb/Nwr5LWmn6SUOwCO6rQc6W85mEXE9McPPv
e1Es8UbfMMR41tTMguIAVVGq7kgt+zKv1oRvkKicQKSy8zIYR0uFbnV5gjlX
Pxkue0HL/e/RC3q1/V1wBdSnaWIuh/OwEAAWVot5CqqsjSAE8iKB3iWaXfwr
/DHl4iA3R13QFjAoMDuo0faAc8cB3vzgSLR2vQ+RKrhC8d0z+8EaclHtKZXj
L0e6ntsV2hAB8FHQd9jVNyJIFEXqozYzhOYQu0qs2sxUJOFxNk3SpPn+ctPd
a6B2qb8qUqJf5XYW0Mxc1v4ANH0x8PKfjR+bT13qBWwCb5tM1NTORPAUnc7p
Y8asZvB+cKX+MRd9xRdQi/GljkcMlekrYv3jpbEBxEGOdHXB39bkg9JjJy1g
0ZXK2rl2Hjw9b1x7XlrzvAODNQ3xL0xGt8sR4js2/+ofjrtplpuq06tGD3x4
Cr+46AsCw/6D1Y9DS2cQPrqbUwXC3T+nc3rKY+B7WNZEo8XH5fV6bWdZLcVK
+DFy3w5xD7/EFYcXaT3jxv9xfJY2an+0JNeoxJ/lE2Z8P1o8lHGrjuJ0OH4l
7duExOMHqzxC9zSWePxXhXxzoRakAbhr/yWN9q4MYD/YEBdj8+s9lsQcyXsG
rSW0lS1Q4NmoMgEm7C5kIPW5B9dRGpEJUb2raQSKNMXAVYu+vS45oMSanQkY
F6c2Fr/iPsJydhRVjld42+4NrXmwdIyXu1WPCjUWxvKs/7IeGStbJHzWsTxK
fo3A/HGnDYOSrFdSZpx5exISpTxjq5vq9VLFDltoMYNVwgZWxITIcM5H/Xwk
ceu+FFJna4PIkzwW32pfjn7STVHMJ+mti0cjy8jBxwhNmzB1f+z6r5wFPDVL
8MCWHmQWbU56pz4eFf/RKn/k0NDK5UJw4Dtyklr04cHv3dBaZxnFEOo3ldrD
8cXjay4b8nGHzNsBE6gT/4eXG5iNslwPxydziGhgfu7BiV9ahdIrZBIe6jgl
oxKHcWlPax5OCpTTJv4wfcQPNRGpnYIe59xWruRFVtXkzGRUC9dUTwiaJmS4
BJyBCraSFFUNe2ESjpwnlkhaaC6PjvtPEDyYVJMfqNCo09SKlxLpCa1vkL5K
RSqFuyNweP/oadQnSQ+DlFy45QSAJNof+snBO/FGROkRhwq+t+tSV01wT+M5
gbi54ppsn5lgfYLfFJwheM5+DO8VBG7c9ovE8TicnbPUgGnCSnMNB4OnIfnu
0VnYgtpsrvOhmCj5pVe244KTT91CC4VbiMM6jr45RFK3SzJ7WCQwCz7ISKyv
Ikzc+6V3QwOUVdFdgN1z4YVpV2IzYPdTKA/wD9qiK7S8878hcMeCqaBEVL/k
DOIT6DEHNpK/njJgPZX43c+oFrppnUXfPbD0Or6gBzZG/BQV0ZjBBlP5pA9I
U95WJHMrn8RP82/HF68/dmCQva4dkiaihxJ+LbGjj/dQTFWuF72ezKpaIifi
qh08xrPqz3QcsU34YlzSgRFuDpXM6vk57WnfHVE11Pgthji865UNWB09cgFg
xVhQ1//DctgvDOwWag0CNl5xIkAFFxLGyz9O0x4N08jhqqe8jpT5aQgNk+U6
j8utz7X651DZZq7yctiwlDylvnqJRQVQk4l5MF4y67jc2voC0AAwdSrzBKu4
p8Mq78OeSnbnffZYZ95h72IqHR1fntog3M6biAVFNQ6fr0OWAfObqFxUpLyF
QxzmkQwqgZZ5ddkzw9z1jt3Y13Qc0oDwjnlf5mKc5Q55+Imw1eOiXV05RxHH
P9gBdaqdssnmsE3/Nhbm/AZR4XvNfSTuY6ssrHlTf/CDqqGTGckvSC8J1ooF
udSFt9pAyc68784BSPiHETwZrdq8iZ3Itg1lFrqnPPYHu2xpAT4X8dvs2/ZG
/hoxsY9c/JnHPjluGaUhHcekE96WY4eWMRX5tEf9v9U5Elu9U8ZIzFZKEavX
ylXjYoEjW9lwwZnS2q2iln9XJrlIXgqJQLFNsZKnzHMyikk4m0Dsf5honj1N
H284v3hNpDatZvjIbyVdVqJAS3KdA8T36wyxXebpFFSf6ekW2ge1QgJhNyhU
68zuttGAamhPcWOHWB+q7jVOoqXWKsHFBhbt46kpSLPvOj5spEhZFq3GXoQ1
aqIQv92sdhTha2/1BlPXdQcVzGvqML8hlsYXzaGijYWPVDjYRi5cc+/Hm2S9
N+jRCbjwF5lwSgW/XNNPVrKNCstRcmjwlHqo82tNiaiJF3qnS4e9k5OHnOTG
v4li99xVwiBRc72nyKZ8aNvC9uNiy/r7VYEi2U82zWumVeOLOEbAIhVM6jXP
MHIszl3QS+mk5QNu4MnTJK2i1vK+guD3J0ziouf4wIw1kMFWcDWa4m1DIJs1
VBhHkuZ9s1D/B8LAZX17lca14mA4VlNvW7NELWiQsFAhR7iSuTx4zm+K9JzX
LUofAny5FfWTwP9oUth1M8oIA/6+S5WgSREDOx/bHq5S7S1QmGB40zH+6LuU
nkoBXAfElKXTEePu9G8zUCunon+83uXemrrUJFLOX9MAA/X9Dk6mm8fwtpSt
+uD0JF1VXmJzW8d7b2nNV1xlFEkNH1K2YlcsQ/qh2soQDepf7yZf9X0jfYi0
DVYAhXV0ZKS2506idpUQNrjh5W8QbqcU9Co5ntCoHs210ISgrpiTi1yXV8ez
5fq/nP7WCdwWIErZy55x88aj+Ytv0YvGnioZ57iDZ63UtecBAQFlvufW01Xi
jrP+JmJTGIfHQFNnnUYa/aCQS95LYQPEgLIo6O7tSaqN0khyhvepZYrEihwn
SGBmMEmWeXsz8WJzK+LwXPOR+y5Pfc4kYoZxBI6rlJxtyHuX+rh0VLDMwlPB
IiZKz45G76N+rpzpiVsfocyufXN86fSUdakm5fkDpejPxd1U+48e4O8vVWUk
nwAVGwYPZXzXBDog5RHB3q1KOE2wpmXi/IPEbA7KvLw22Njn/yedLvs87WbG
2kM1nH2DmYlOHsDIRtjnCXysh41sEVLf+36pLuH5OiUCkoChn/+klTHDPTa1
ggNHcCisYNs/OSlFV9llEzVOSGQ5bGkBK3bEpiEzDEK/5HQK4QTrW4qPAUJq
QUA3TvgDKrg8i+bDrH6IzykKbugU9nbIKEaEYlOrThuq/5di46Ch6rsZpzkK
FJgiWx13LiwlOXecwFCy5kNH9XnkJ1IxfZ8qxMvC6rfWrZyLS/AvcmvM+4F0
y0Eq7jBT9XNIemd3u9o9JICu6DHtulR/JSH9GJ+Ae8BM8AV2qKbuBRVTHwjp
M9de1QSd2KIxcXt76U1M+dqJNWbvwYyrK6Kr6dU/cjRsFvN/U/bI+WEtYNdH
aItENdJc6bXVKtJUyzbGLtv+2L2EkjuiOcAAjSLJ6+9pzVpMCtwK3dm8J5Gd
c/SlbKoEsEGmQW++8O5su5Wgf0CabowNFovehaALvbiEeNQbF97oe6u+DWQP
WJJx9ICnhq3qVxYXWLYrHFKfaRKY0gJgswNBBcC9g3okwKW5dnMV7KxRLCsP
jWu3T4nFHxVWmOz/owAAZMl6xeLCiNSnIAIf2sGkcHji/gwtrCUx3TMsxJbS
GJ9x/9HQ8SUqh7cC8WLfu4iwFVRUrHVTPDBOrMK3emLJmsUrWWKI9A04PM57
BL+CD/aKGSg6FPvSvx6QB3xat/XubqfmsO/cBYLiRBDKW9Lql7dlUM6W+OK2
fFCxsalW91QZ03t4l1nS+0oS/gkZg8MIUnuKaicWnJ9sWJgICmXvZPk7LFf9
q83pXlSJe0sYF9759rdntWre9fF6ctGBYm0IwaLx+8NK/lbiocGnHdzKy8Nn
vgRzi2Z3gDGFfYXvjT3G7hZICYUUZqL9xY6F7RxNGwsUwr4s3qv1CygdhzpR
0GYM8z+AvxiMxFpkpqLLKfIdFzXOM+JB9xZio7TxScaPXnmWLXujw7Osnewd
2+iRaAZBrZudKhGqxoPxd0JC5XRMS8P2lvGLCInvTQbBPy62EeXTiSjD9J87
SPBocrzlkQq56lKsnjBUQl0+emHcBHklOWyStRnCpHwjKSmu3tKwsf5ZVXQ/
pCs8JBreJnmaWRsyaemzjEyK3gi90nARM+ci9RTIiBJ4ty+20Ti2haQ2rhoY
DnNcR+0QMDB4l3JxG05ym61O7o0zUPuUiIZskV2z9zfx90JvoglCReolg+3W
HJRwe7I0MIpfjJEVcysvvhYFAWvZgMmAN2VaFa1Iu09oxoAnekBMr6R4sH4R
QVnY+Hs94wGZLF8UQE54PEalmdzxmGPVxgFfGsu63U3+YGYVqVOfTSlVK64W
Ol7QYnzEtLkEsmuKJFTaaXD5jZHMCr3Nio/xStxefzAVMxGIGW+3lqJBfOtb
fqh2BDXpvKLT1trNuOYTHYgu1KtDHtvxT9OeHXhvlePyRPPQXd+jwAcpD2pd
QYsulimhOu4wuqtiDKo962/uL2f+EqCSC1+CG/w8w9VtsS0q5oGTZ5aJpuOl
FQAvC9WMriMf3stdm9JtBr7dS60DJzN3m5VvGPMixhBbdvGG7CrY/5ikLtrQ
e9H216QhqUcoKN25WgchFZeYCjt5MeLfBB8fYOJsm0r6UjrcE45ZJG+bTeXm
UINNbpdWDWrEWjPMEp75rql5jwMzIxLjECad1Vi2MfxlGQ9177EdjSLozv6D
oUZrSE6a74NlTqzbQ6OSH2zUJMzdlFo0gjS9jQCHkosjeKZ5u8vJyTLKM6sj
nyOiGukHdhkf5+qCivTwgPS3oC28Vt2gPVDAxtjGilcnlA2fbjYjf7VRoq4L
Q1DpP8RL4q/o119nNkDyL36YaFlX4zHBFwY3d6YMkvN10jkLo7HScRSVQw5e
9PvQIkHsI9w8NkNhAjExsocMoyUzaCuh7sYBGHCmlHbIr5aobchmteQ0B5U9
RzEnbioMW1aeyn7YdCNDKWa8BeP4b9lOJGUJX6SdbxrEMzWpSyKpX5kcpdRu
NclGRQG2TFgKKj7Ywd6Xq5qcyiVeBRj+MgxPmUyMG8J4CVScMNZhuBmESzyR
iIfMhIfX2AoylEOp1LtetDsfqeDj+1dq+s7r5fGOXLWzN7LaslZWNxcbgzq0
B9BS1Nj2g1qggsWtB+BVmRpXoyR8YUCC99UcA5XxXTRLLPtGaGRT1eaGvV/I
k/uxtKBoQYN2cHpzyB6fl8habHGEqFbWKTesIT5bI9elNT8P4nY0gi1lXwK6
VICutK0E1IhSqdZBbxygztSCCVBcYLi4hqyB1e5RuhPXy17gNflF5yIjkeR3
2imvswYh34ieFGODlxP2NxAJFatV0HYAkB810mFrOBOm6SLuJ8b+iWLGIK0b
/8ECEtjHy9G8aACQzbj8EMz2FukD3voeM9CS/0PsrRRG0g3yLKlnNzR01d6x
5HLFZcUfpOEH3ew78N+u1SVozBQNC77AO1OQN0MM+quydsNsw4EbQetn1TLo
CYo+TYr/Z8Kl4Jw5DycpCCd/AugTZGU3MhkQLx3bZyTREThG2d/y6sKkDTnP
K9yqwruLNeKdNjqVxlP2ZfF707qSk0eAJCT4vVr6xkNZQ7pnCjLCY1kKfqwB
c2aTPOUiTtcbWzZCVoA8azpDAWmmdz1xkLN1WAbCCtBHQdBr8LX5TqEvME3F
Qa5EZxjImwz/X6P+H8y9/cjx8oC6CdtwL7V+/lPF7yVs2yb3hWPoqysmFhHd
JWD+Y00zLxoRaJSNjYisiG2VLMFY6kH/+gn1L8qSd3GH6HyUQV+Ek6MK22DE
PxW1XAMJZCt3nMy5Xf11HPRlBge29UW5ePPcGDIK0UE8u34MtY/piflOLLB5
np0KUgPoznsNupctN61XIi/q+bfUaUuksYI0Cedn3GRmKiw00XRMJdoVbng/
yYSF2Wgvsm/Qj5mX9Y7wkm9OsiaLaRBmjAikM1NMHknkMJboi3BJ1Yz2KpzZ
hvSx8bTXXbq8+Mb2NCia/1Q7LgCQXB+0v/vmQaYoPR6s5E1FLUvQ/7hINMkc
b50Wbt4WvYe56kqvoLvVgzKuA+O0ZraHJWDtHD99rBFoin8KZSoHDYifawDT
afP8Qwwzj7Z5c4RFAdkDhHIFLxckKGSiXXq+ODX9DRmGPEhl70IHcLziopV3
UcEADjdVx7OVsRNqezXSq3G5uo9xbfQGlBb+qmV2CKbxvsUr8tSFPzoUDOrf
d8ChFj4fxN9FuKmQ8IIGCbrKZB1W0Nb4lTYJZ3HVr12uCY/+YFJ1Q0PNletx
U1ynbSEHayj4sadKvtiY7FUKlfVUSmU1tOxUGjxP79KjDyvjr3HaB28vyi0Q
x7rrtVoeHJ5SbCrbvxqnIIcW747/BKxjn7wzRb0MTP4MD/tLNCFChs3g9v5N
yHS/acXubtQH+rQKBItJ52E+ln7ALNbSnkfO1axEJxdmxndPJ48ZjjGg7qYt
JgDIrhq9bDpsz1leBjXUYBkvNQKsVtCOMAJ9kD3RceUOOJHR5zW3mPYNSQ6x
TjMU/an49DFTODyp+Fv9FBH4TxPrB/qGuwp6kBvKIZK4+9uUUXWXlOmvQaUE
UE8flXS5vRTHYqRxJphCnviWVK8D5uGLE4uN2z6AYRGrd2T08eD9/tPKXfXu
QfWd1NQhLIvToxqvgKHspJpSa7hDYEslZFWt69jkOhg2Cufip3GDh3OcSkxh
VKYQk+vmBNa8EbX5zbDDJ6+3HoYISMg4bCw88nFcsSob8L2zjWk77spxL9TI
7ygaqMTUDiAZNYUcX3M6PWxnx7bcG7f2qZTD+g5fNK43KtIf/ioF9WTS/QuF
M+iNrTOVXLVqK0u2nDRDg11eW8wu2AtmXx99sYKwmPKb+z4Y3jp//F5RUXc8
1XHxLqvuUnQzFCv11I4TXrurHhoCc/Y+dq8oIeiopmnrgBHIOh3t+eOW1h86
qHdADqa7WT0DrPbhXtCVVWtnx4cRaERoV6tZckvWwA8760kq973bKr7Fr1zj
ict92nbMQYLO5eQbVGYEIPg/n8xUBsKjoPemBRuAGYguAlg2SABY/uDJag4J
9AjBijQ6SaE2MnS8J7LYGKW486kuFsGoWxjLZek1+cPV9MCE7VOWKU4ZX2EJ
fwOCY4cfoKKtI63DeLinRTclRMk3TnA0q3ut3VXYFoBnZUUz+HLFNMaHZbEu
Uu+NZBzQ1n0yBo632Q3lq/hulSB72S/u+m91TAsu6al1kAoRZARvmcDB/BlE
J4DeV/D+Jek5HepidLOZ9dAJteb3+lIrYlz2lX8CpMDKGf0IKOS1hxaLm3Ft
WMY2jVMm6YOOv6TiFPeJEIsBWdi98/X1+N5tfoJmHVRORjYy8Cey1XhJoLqh
t+rv/1iQfHCk723X3jyxmS2bXcGflHfUL+AuPnFpERM0nZNHDPWwcIuxqmpk
g2b+vNEWwMio4+0OujUefBJe1X1rFPph8pHpRdWwQC9PeUGl523KtJ7WiLA8
TLzGEa+7BEBzRQchJieV0H8gOLcgVMWx+Xe5gGdeS3W6Bm/g+FGcqdJrFOeX
TIzAbbvm63RSYNqieDqe4UQuX1mTVhD+Msnv9Hm820XJ9ZxW20cHleqq5J/L
cHnp+Djw8lEvug56Wb5oW3889weCH4QUZx+HXV6E6N+n5m5l9AcG0rZnq8DL
3/bi6bga5bKDTEWnJETWjUQwjc/LWGR/Wpw8n4xqRNgBPEktU/3EsCLJIx9V
6uS2DGg9vEHnHE+X2XUYEkZzVfdGB35maF4110alF2wmJ130W7TIBkJfQOod
Op43naXbSyn1z6mS7VbRjO6bDZz7R+O/A+WEEkaBdp8dFl9s3FXm1UJ4VS3T
ZXkn9j0Err2cAymv1D/0XvagJPjnDYeqWgTtDPbyzCzOwTmFwMMkz71mTZut
+3Jj8FXsrXPIaUi4jOCGtZ5fEAi2nutBbFdr3dBMoQHNPu5DZSmdxmzC1bSO
CH1/Eai/sDQ9mcIToCaHvH/O7/aPyHxEcUR73rY2D950rMHd7oWfzlvVu6Qj
e53Z63lNxZ8ogEY76EuhcI1jlzyaSsVyAZpTzK6aoZAWV7k9QBMFuXRaJp2e
lCsm7j9YGxlCHUrahPRftRCDOHuCvrECp5oN0TNRQ3mffBLm4yOTft3Ld5o6
rrjjzdwduaOF6+RFQYc+hebkeSSEh0D5tfbmvNbZjcnx6Nnu7g6bTbunPNyx
pAt5NSCl4AKoai8KhvKDeYRbl0rBL81VpMnZbPiXxuXA95oJgTzclAPU7Fu7
pXzp72Mdo6vSBjufqaCeYC9ayFE5M+kAVM5gRfMAit5h7Dds+DbHPstbN/Uj
kK1cRZKw3UblY23dk3iWGGvRHKWZlB0oqVsoIiOzJLd6vVkAvUjbrcvkXmi5
kh074eA61qumTy4O77i8lqDMpjOBGdKPlnKuHlhx1CEWqcfxg5OEW4J0Z8vd
z2pAXSxker99V0RxZMXPtINbK84DuYUzC6aWDubJ8eG2S/ReIN7zDJO+fQD6
cVXelKmbZ7q2oNY2CTSskxYq8AMeW+vJ9qPx6A0HavzZhXn63cGf0U/GD3X2
aHn59T/w/uZ6dpSmHbCLR62GLy6UFr0cDXZP2GzNGzBAmejd0QAztfyOA3wB
s0pB4f9qM43ZzkPThBTusHZknhtBAr+v2Jh712Jb9JnvihcQXbJ6H/rzlXWf
mLhJYNkH71/0CvH+1oVN0hpDgcvmtxXDTNSePh88A4mEZxFKNGE4otxIntNz
5ClELAUy3WZbTdkDM8SYtRtrfAg7hs4UCCWzpwRC3k8Lan+iC5j+OhjeEKcq
0kUuNj3umzySSN//YtDOl7VwVC/wfAivUqBbyQN1/LxVFuxD7lBwqRUkcS3A
CZMPoz9y6Gn7ePzJt4CfT8/yNk0tbQyQXECSG+m550wH5nOWXkeiRWeOtV7M
ekL6HUFZ3lFw86iTfx3MAATm1IpS1kRvTSDbyyAhoTivZPoHxVyYuvVj+26d
z4xEdavdFgXizL+4sCqn0wbyDpuzZ7nin5slqIXVUsh1mtjECYbWsPFxVZIz
Z/ki9x6X4p3FYpX1bG3lvAhifKTaKlfBz8jTC4akPRk3OocQDOlJdB5AQscx
3kmg+7xByvyOpaLNJDIKOHCO0mStMrvYy/AqcgtH7DJG10LXFNEoICXmAn5b
GQDZEDS1Y+gH6NI9d7JymNdgdItXW1daNsuzFZXpKuJN6IV+djtbe7kNqEmd
FeAeAPDK8AZTF56No2c61QKTBM9fJyCBugpG/QbEnurkVMvn3ZmuJOaZGaSV
xvVz8PGem7Kdsy/nhOqNp/GOOM9Bo1ghJxNU+L+aPnjCXqhOQ/+sEG+paKNC
EtgxCaqrcvEobpRfpAeEhZSFpfN438qsUzNjYNxL1ywuUfLjNLZS8LyoA01z
85Hac7mfI7pgqxqNj6eaKdQDHTeDtlegfX5xjnIaNgfTd59ZVcfOAs/Fkg0Z
RgouZaYmM7j3hvMlrZ7S05yx29C4COBa4oTngvEc/JBqxOtfPgYWYFRoQgKI
tlg+Q4PUmzpSkuZqJLGeTPtCBGD5+9/1Eqw+3VOBbLMajtqrWhV4ZAntSgYm
jbRohS/FvcxFn/0LKPr0acuVi2fBpb0B6P/yjZkpAN20HymiouIiaPQNVwuO
9oK4AU5nKMyiDRctRXePIWwnOJPxISx8u7pcfuT0ytc7sB9OX384v4T8qyvB
PZoTEWgMkQqhkTnZ1TV0S4pJDV0m6nm7XSSb0KWqGK42VX16vS7eAcaC5+zE
PjnT+wD7VUwSM+PloGztvHuyt9jnnIzNof5D5Nmsk6W0xK96Lqd8Zg3GA1Cy
RVIrT8+Fx02x+uJ1RvPa8sH5ZrVOsBR6q24NaN9bTwsz+I2DMaHtpIF8Q46z
j8I14/8/qI2pFdb3vIn5fNhsV8pX30iagpWIKEzz5Pl4fDOINctpKE1YZ5+e
pLIn1UEej52+h3bl5DIqx4r+gdG2JUSORzLUFd8llXueoEnVqVqDMK5ycwhr
WZNZLWGZkB/xTX8mgW9ZhIMdHPWhJ6ml31bvuDxRznldFLMs/2JensGVikua
wpLTrNvA36TlaqQDeJY5fGdUGCYmpBlKOmu2OkP1OQwCAo2P+nHZdY3pizxx
XZq2qjVEOaJUvebhf14V8tipLNODPmDLtL6Onzp+vHyO+IEGNfdaXghnECRH
pKYR1aFyqOO1YIsrz/CIr+g18kwLi5rZrLCZordsH8iYJiZz8VZE4BlEcDHp
IJv/Nwha3LMJ3YBFKCP9iQEOELhYWxPFMytr37WbK8D9rGsEGQcNg5KvTExg
tHxHAWVPunG40IWajG2LkeS0KadAVTfiFVxVpRGCG3tl848gk+rxNnhuPFVL
C1kfVJO4nCHaQhG4kbwFEZlKQu8YCahIATzMnaxLQwnarZ4pMRJZxdiISZK+
mJlBO6JFbtco0Vp992kV75KTHi2ENL35gq9ktb+kSpw9dcoVucBneUaNA/Sf
N+hPwdjJ3dYzYVSBW6NLcXu1clRwhPKvRr5ivZgQOL0XZjzhjfl2X8x1gmnE
/jP2XSimnFZB6ALwVJB0Yx8zE3d6ZyKlG5ZlRvQb6N99D2W7fa2Lk1HbQEHt
yV2O683tNt0DOJ2/uiW0SofgVFi5n289VUq/ZT31/8BlOO0U2jeZgpaQgVvc
JnARSMECvRpV4yq14D8LclkVvAxaihqp/ixAv/xnLhQppbK8IfZsENvhC6/S
3+f+964/+c51XcWdG/cqKBL5A9Ca2SQ64i9nNL5Wv5e2G27nXwD9aFS4+dfT
a7YWmVY9jIHPOnrQcJgyYY6tJE2w+XlcvOBFG5zOSaKRGEjN2m8mzs2JT7Cc
UAT8VzqvSOskF/vqbRgHqn0ruFj2UJJTWt1lHDDxsvScnJJhHZFUUjh3NYSy
knA5KY0EdCmdInoE1cYlgj0P0nsWD+Vo/Np+ylOR5Oj6xeqRdLiMVEcFayi4
7Or4ltP7LODlZCeyt0q1c5qd7kzLRy7vyKdNrzLF0aMtTOLHaXdIgpsPcLVS
5vwI4N+xNnMlE79AhCvQOe06lBkAMwib7sEttc/JYb038d5YbJjaQgvBOeVV
M6IM4rrd8yjlIoG+ohYMb22HtyYcQT78KoG3ItZMvxDVGXSg7sddfm/PFfMN
Ecahhz9nj0DtU+8Pmsptpw08E2MXxuYFc0wfBZcWjUnCuEjzlusSxTDTz+ns
5/swjrkZMKHnKT1Kf4DknQ8rlznhoFLWWmTPG5U1PbEuQnxdpjGYAYJ31YN+
kPkhiC0JBpMslDcHIbXkINuhaJWbbHQgeP5yS7MnFtbh46MpENPV8XDT89Hx
kZhDLm2CVFvv6pS4oqTfgXwY1+X88y5iXMnOGSmZtgVBoS+Qx+XwI/6ti3uS
glW61jIt+8RBlgHZkn9qB2NBAAucDiOOaUwULd/lAK67EEyOU8naHf2gpwRL
8xvNqfBFJ0iAvSCqGOLWedoho9Njr36uM+VJ3x57yOq0mr4uBxDdbnCZMnHc
UZSqeKvg3C8BF8ybnc/0BcjDjLP1EXRDApVjdQncHCgScv6WycBK15Rih/k0
MDp0Qbl0Fz2+JLExLTV6Qa8Fs8+v5yiYb/AWNWAKNCv5VRl102ojT/6RLkIc
R66o6enkxu0TGQTy/NwUsImewsukeoSySIkFI1MLfiZaqkI8A8llOSfMrKir
TysgsnVP8ol8uFOXRPJxftYAnTkhtyTsPR7pmHhGP6ykuvMeYTigtT8sS20/
8IBERXm7ZTqDCmnWumbudIG5SxXCYtyRkjl9+DgHPMrnxyZ7b6msKOFpOVXp
cCt0EUvQDnY1jPGZV5xBKlWBWnJhdtF2ydlMegdPbaKOEoi5a1Sx8d5NBHsY
gVkbb13EZIIg061JHTSQkGmy42mFxfqnyso3sG1oGqMo/5BMFJQM+lH2K++E
oR0JhTQBeRpNK1GV6qqPOyh3iDUpeghBKjLAbqCF7ntnuwLKs43I9BD7mTNO
WFP76z7YxlNjKZ6JVJ+WXPEollVFw7TzyAZhZ/ejmHPtYYlqBOp7vO0DPcLD
wcO5YUnNtJJ6y0JpBRN3tHTlm1IVdQC+3DHNPrp9XhdvKplci1l+JKBUDxXp
26yu3Olcu3wi0tej6EU/vgFWvmOTebNJz2QXarMTujvpigP3WxWeSiw6xbkV
HXuHXodamcRj6l7dyC3nZJOly7o0qRU+xOaHtMNj6u9J2LeZB6ZoiLS90Y7H
h5t4dy76+y3gFRKKlNGWmvQVNVniUF7n4lv5ChU8Ubs8JO9IRakps7w6TnuC
XU2wdXQ47NTTaGNq654TEUStpRXMAni2aiigyYCujDUr6JHZp+YdSHRzfkmf
CY5jUsXGIfIFYv8VkMFHePldai4bhFortdvjJjlhbTWKhVWW2Hj+zRx5RN0v
bEv1APvXvyMTe5A/IGjbILwLY1P49HSpDqWLmorljxm7AppUfuNdJFmszUw/
5b2FB8Oeojwn186x967PR5qxIGWFs/ovJ2+lb+pX2dm4YQbU+kkp77oJT4Ny
OyOIFcQjcTpyufn/lIVqaex+fIyUDgXoZ8xmSHvFNOu4mLVFrTRYLlwkpRgT
ul8w4on+CCtLCYh83RiSFE2uZ+DqyypFCB6ltn/CvVl7UVs/6w9tGme2itqx
0t1dD8noRDmDFa9We8vI3WVpwJs4xUNJBhI8dry6ADG9Fm8rfVKeD4imjTTF
1V/XhAOlehZOFAz7mfAHcTmV++AE8qbVklMFsRI5zdkfjZsE75mPJADpZXFd
AgeEKf9EvWCFIMhXZPi4tsiHccWao+AaMupgncLFOnMism9bVRd3t3Mj3KoF
o36nhaULFy2R7bYJAX34ohXv9fKOGnITuQkAIK+tvSKGlrli/d7UvArzJD4p
dbdoPusZmM73jBf1vh817iLsyJCHFb4N03UrFfTc+XUvd/O5LGm/Ty9aCFlr
21LFLuuCRxS2kkBsUfsthLOkSq7OQVfSJpkNSWlWwLu8gEO+4z88UmXE6AU7
OUDh47r7yHdI/pNk2BWWsrxV7sNgbjG2vRxiYY69jZ8/I1FgVDp3bT7gaW/J
4PR+rwij/XuISNhznsikzYxjuwduiyrboXfu3i5i7eb++6UByDd0KECY1hbZ
xKur0H3g7A6StuBY7cl4zy2eSfRIMQmUaGaUuUmHpDM1GzFZWqp3VtDM0zGR
IfGwKnSjM8PxkctbUXPeiypYBCELSAnXtyuqrn5Ci9x7O3K1oHTtP6TWTM9m
tR2OWrmvDiuRECpfJAfgj14quKEZnhU4bNpjBD+NSUvjugbKpWdXTOv+JV5E
WMJFDPX/5sDZa5VCaDCsgTzhCtYlp6E1N6B4mpGNAkMGyfY63MUzDZwlZHG6
xdSGnZqUgkFMXGZ+fzxoR7XjQhDuC420et52I9PG5QCnvzQElZ7eJF55xbOX
Y4TiIJEHgDNvqNJ4b6N+9NqwLv9UVq+PNQtnOOoIeVsSKiaGcCXNX8paGSaS
Zp7Xyq1tYMdok5XMajsE4RWFzBLQbUeTykRsdVL5g5ATht9Z6ivsbFfYq0eF
ditR9aJfwnlAMy2bHFAvh71gqr43tXJuKMSXZwxnRFaMLSHx99+hKVkFaYZp
k0Nol6X8kyaBpRYhoq87TJ3UiS5Q7kEJ0ftUOUGvftlxVswYErFhpRQKk0e0
OW0AniJ3/n5ENkf8SKguTdX+z3J1fttO/JSxYB3qvZIYU97T7AHr9HgkgFen
J311gGYUpaDmkGE79wBsrspShRFHa0vE+6e0tpZCS/zjDSE3jirNRQzix1Mi
uQsIsxsqNzxLWEFNb/GBCz0CJW2BFyOx/Ii5ZdjC183/uOMn0eOBEQ2DkYa7
5n03M/X3EJMm+8bd4seVmVj9V7cIGcvWGrTNvaNfPIwvanHXl5oqJ9v5bCt8
BYg3GRmXU+2KyRd8+zNjqHL1BD5b8h9cGSvfiGgPSxh99eTVK+S46sf5gzyM
aYwlzLaLMz/vxq5BbgC+1aQBPE1SUiGyLKFhdvpQ51WyyL+UHjHXmzClLFZ5
c8dA5znujDVlQYm9Wvqelda7oRdJBmIkb80ysI6WaEjRyFEZFrFxvodoS38O
5SUmokdAiWsntMM2+RGuhi566+KcBZv7Yzw68Ua7X6jGKfz8BJnH+LWTQH7V
f6Gr2DcreBVr3mLl7k85YAgpxEV2qu8Te91HbPvQFci+3naX4HqFgIho2ceu
5yTBfklf8UpDKo30ps56dAezhVvWJPaxhWxyItc5uDu0Ki9Nan98eOaBxanw
PpgmtjiCERmP9Hewd75XaL5iNqhNWbK73CO8jgbVrp8TmPm/1pNlGcAdPumH
wzXpMcbFSSbX7AQQfxE1dplk2OmTUD33wjRnuCLBHgHeLgMse1ZZm1S4Ynfy
qLJI7GH9J1/VW2ZBrsyYwGLj0sw5eBdxmyLiGlyRoLVd+JrqYud3eVXLXNZn
Y+E9LQInxl8IUskp1fmgz1u9UTrtZLDfKr2LMn+Fc2EZO/hA6PlR56HHZspL
Fse3WswhMgbxryn/qsDUKFR9rOTXTEwCr3RfkOivNsS4MOZmfuvQtwmr/EEm
me4nHbnxSxCq5UNT+W3Ht5hcbh/3AFVuod6FOtfdNDCx/bb6xx2vf10mhJst
CuFE40e/KsOygb02F3fspAP5j8QOCCzVrY3mD3B33mbzKC8pLURzu4yEDWgh
zmn8XwjM2nSLugqrVcXhRlOlddBLipcorAqdxO88oPsEg9mBU9kPjJEHOF+v
4LzasTsRYlBddcthJhkHidUkbCYWD2Ld+Dfpbvp15IbfEy46K7TPjmOecVnz
Nu8rCtqEDf8GB1GVhwd2cOBKDw69rxwzOCnJtRgSryRjhmu9EI8poCeXDNwt
qkSw9po+3cZr5B+jkPRei1LJ28cEYIKNeA9AOhAWa8rqciZwv+SRRBeHbYG8
1I4Aa0LWcBeoqONhJXtzlRmRrQDA96w+r8SgeXjB86s6HhVS/QT3oJ1dsXap
Yj6nbvOE/JxfbUyjheUPbwfCzUimBrFUrkCzBBzoQiU7dQ9bKuqqw9BVnyv+
h1IFwlhAHEP7D5Mrh9m2leJwbDfzevRh833G+SKFdiff8LbCpylaYT6Ia7bP
kvW8Ol7aJoUmJxf0zcyT2Yck8LJgxd11gjAkMYNxFq13I/sCavqHE+EHqmxP
eFtpGmRpZjB8b2CDE+mbVpNx5eLLyZuDKUMUd5lD37uvYeL9O7bKZ+EWBd1G
sGA8VVZXMII0z9FMfqkFiChNOLtSOoiab9QM4esd9mq+6JVfbGyUb+F27TVa
vBrAowqYjgmsyI4G5heGCse9TFQYj37474D3e0a7L6eLrYRzW8yfmaajg1ML
6WSbJLAHkLgUx3rr+7x9Nl08ltn7rmabRi+4oP79w9vU6EW866424As2z1w9
pMWkoAg/o4pS0esqDYROUHFurkzZHoCDNdx0t2Qcl+082I011K5RytCbZGFW
fNnJZHInZC/WazXpnUtNQ5a4UGjupCCZYKYeVH4mDTPOwbpqIvWx4bPv762C
SPO1u4/oSadiYO45L0Uyky50NBFTkxONjxzq9uj72FWVExYOOPkWrfEKkbkH
SOm2DxeOd6y4XFKwiQezbWUj/Ay6EzhrFZGkrl8bHKmfwV/oacmBpBZ/p5ll
tLsyZUBsvuAHzIGRUaZu3iM/gW2N8nxfROz2Yj6Ui+6DnpN5xmUPEiC4FSyf
LeGIKZbwCnusDk8bZxTbQtVCAJRS3L60r6BC2FKviQb5SB/Ig8WA26OCpOQ4
Elk6V9HD1J0Nau+IaTqEEsObaIPs+HIPy+qo8/1JifjXlSVcloCVckCNtfaI
zENLIeI2/QK0miZeo3Cb/0XB5uuT+l4iuoGAGewAdBeewMR4UjiBlTZHFBrq
jlZxk+x5MnlRYVRYWAYtZ6TGKaYV9KE+L4BZlUD3f8O9rvP2/cMfnPH0S7BR
bM0eL/ZUkfWViTn46bQCt17g5+P02q93cUnCNiMN17YlGx4YVyBliASi0QxD
W+l7TVOyJ2wosParMnd/QB10yxRpVpc0SLapg8GnsTOtB8Quhkj+Koz6h/Ee
c2AqtHi2xXRoCX1+MbnDErQ5CaBykCfKFAjfebV99V1Ij0osK16lXo2zDDo4
53mdJNiI5U5OjIZ9B+2FqDT3usFlM0UiHvE8+igupvjTl8FeeeJON/nREj9c
Lj5Ojft22YZbnxrDjKjqKIsnl/OQRWFwUvvz2mlKmftGhW/05XyOl78fGmcp
DHNaoNoBIiLXjfcudNJp/aNuNeQhqMgikPrlTFTHEY8EXg/MH8yAxRZWox8W
4rwgWMR+7D5gmKNV1TUTNH9Wa4QocDB8dFmqDegpepTSEGsR5VZ82e6WOsI1
appJO2NPmEkp/F58LSkHkUIGVoMg30ZvlvItD2j1+CthW3VpXdv8BMZWxc+k
zht+Bf1E6iOUT+RwYY+evbNcanDqTCoxOTCXVK2aILycpBQezH0xeb4FCuMD
eCD2EeIU2a4uLwlL6gY/Gm55QdbNSkZOI60a52OVNaJ05ugJONbl1bApyyuj
zX/TxiCf/bYlI5+DbsO3ajacJazVLlLmJF3FtUtZoRlnSh9Nux/SFrX1S4bL
7CYib4ZSSoZ5rYVNxadSsPx7MimQMyYohxs99+dJAgkg/7itXR5OGhSdxafq
yPoZlgs8oNVnJ0FUPsZKQ7Q0zAqnvLHybVlwIIVz0o5iz+0z05drvTowbXiz
pCAfy2BEhWlaFDhXYXzhtaGBmTFhHuJdD5zIMzPlO9Yzj1vNKoRE7qXZfXhf
Cq2wcVyFOdXvPaVCtzFWz3qqAd05Kyemnc1lL0Vc6v6QEXya+Edu3T4M2kxv
hawS96ev/NSXlVT76OXEAlE7zRHWqBNz4ziyGYyLxb6Egon7CXSEZsLQog9m
s/LgDVR3jJ2C6kjbNLGusNVeXfClNEIG8BcrCqSngcdJIbd4TOexFMPlHHuq
mQBhAWdKFbvYAtOorfigpqdNKBzGkdlQxhH7PEkjx8A547tjRP459Hv8Og89
JicLY8azajfZa6omy99ICdt+6c+eJRUsQfT5PacV4FNXEnuVW0C0qDcu3aBT
1crFKvz2mOHIZ5MmVbAwNQc2E1RC98tTgPv6ew/sFjw4ipa2DAFIvdsdg9+I
KWpeI10/Gpy+llcOMVQN/0FTD+WMc55/CRBedVl8lD6mlARg5EdvOaWmYpy2
ZUY8X7gKV3+SiBpqDoxbYui5SJdaytic3jVPGhCImuTWDGz4yJyWos2/IPMM
cZW1nSjbZKIO+aDnClzKHmqmW5XOuNyoRWX5MGE+hhGGic/GjklclurBdejk
0dO/SJi0mrn/K+0n4UiylNW1Ac908fy5DLMiUh7hUhR1J+ZKootNMO/2K5Hu
h5GUIzim7CtffMdJGpwGDVpX5mDDweitIHQhHFEMvper47qUnPAg4n08wEPP
jTUt+bgDhui9PODnyWMBM0JtQ1Lc2PGlbpQmMq32b0nJpmfFlSryNVzzrabm
RF2OS6bjQfcp5Q6LYyt50mRx7pzMfN+yyYGq7Ga2stH8qu1Di5Kg3cZJSqzB
35Buyvl9LkEPSvwGrbTpGUdQKkeQ6Slq0rmKB9i294zMYFgk2qNKkjN5gNDT
TaxoRC1TJe/kChHmsshN0Z4/vehndNBidvbAZnAJ463ES7eoWFT7N9wVEYOu
ZRWvxO3U1UrcDJ1LwqmXWUhbhMoiI6T7adUiSv2UcI+u2zkHDz3yN+3jzoBO
8WgKMRuC2+bqXqjrpHm1E0Vc7wSpG5mTutPKl4mVHoSEAa7zvIu+6I9LZJT3
pvxLkVav6lFG4/04CMKr0XrPJSeLX9sdrf05v9i97pRofxQA/BGNOGpfgq7/
2DN7qLc5bD4J44gIeaIu0SRr9yKlMttyK3uVgz5L/wCQOJrr9zjR+3LAieS3
xuHrvGjozjSyOhjgpkhJeybtAD4naaXUJkKqv2t100wtd5j7M9yzWeMoo2pn
S6PYJaswuuTewVHN3wMCKyRxdiv3xfMpxtpBkWR3SXovhYaQP00ZcjM9uFqc
x1ZgirgTnFDRjHe22s7czjgk3y2CbF024xKmUD0wRvGnAj9mUNVBtfCQpQ9B
OlukWkVPrWY1Hbz5FB0L2PVzKqE11dRZsBZRgEZX8EbKOw75m72FlzRdvCvd
gQq4RgPQ3k7ygK84dfEvwaT9fE1O58eVhWlDK+FPz9NO/flpQmC4X7KALVJZ
FJWcZE+10rk1gBA2LPsgjWhgvv9a1xQ1fzU4vKLRVNPxU37tdTAxbWWehA/I
1qd8spwe6bP1IoGLBSVOk9RH8wAMUTY8KxB5SNadkiqe6NT7OLQ1xqweTT1G
vPIVJxfS6gg/nGTnO0Gp1FRbI4LzKgsREFb3K8A4a48Z6jSntq+cGX6T55Si
7RGrRuyBUmMcE8InyxUCmlC7JxPMLWBNxd8wKrt1Qrkb5jCAeCZT4QPqB76g
VIvstfFzOakKllXnRtc9yQQ9DYuXFMJIg7F1WA/vtrD0aUnORms9587hgtoz
76T+v6CKtmhWm/l3zC8OZfU4ErrITOm/tIDp+qxi9Fg8nnt8XYELT7tG/6bj
m6idRWGoAthS54+f716QmQhjYKq8z0XnoFQDvXsNFlzVT3DhtIWa/67+vjs8
90/xSeqTVozSR80jXhZ8X/Fp8RuK8uHW3WcZUH1HuL2FGqKrW7r+reAXRhvA
LzeuN91XJEWKODQ2igAin+R4MEHj7/kTrU5ZyHq2T8nHrd1gD//vrUnnybla
PCBdDPaPpSxUemWbYLnV+qfYIouVCl4/j0uve4nraBLZEyUio7M23a+Sebao
Bs55LmaB5+AWK/tRhodntw01fUwOkTnljvv7FwIRJSp6JvTF2BQ9ocIAeYzC
fgl5LErYHz6MztOrVFyEqRhzVufm6q1VUQNfL9ho+y3ipQLx7AYwmXDpbJe3
RTj73lzLyk636zxRwpfXnTGhDN8wLjNVGJX+QFHu3n7WaNV+TtEHtjQkTScN
QzeZd5dZ+xkEzbNqradSqCR/otAgi38k4M6lrrqa46poM3GxHsFrsL2tD37E
ljmZQLvquUlOW2IXxgdy5+g68da+yAJEioTEP4B+J7Zyv1zMGIV9/qdhhGs/
+ALi6wzfooJZN6ILKmTKrLGHvIcAH2AxJdOQSe/tEJczufc1afyMjg6MNXC9
NPluIvGumq0mkITQr9KUW8BBmtNadekWVGuyLcJsJs2L7w3B0tJMUmoVEPuz
sMRBTcnVjgPLBgRI6qTegkRTzINxP8bOmxRuE1j2DGQawq12xA8hzJLg1cdo
yyp4My6KlsshgNO5JlhEU61qMABsrxH22zY20c+7a7RV4urefrH23eb5jxEn
zpE8LH1M15ZXNqsqF33h4D857JgTJRwVZ+yctSZgMCgZEZZSeN1KkhyWn372
VNmvrMETUV+m++jzzIDmhqrUXyIsFKJOjt76rFPxe6xSGK34HEm4NXFJNaqX
1Jv4E/NW7/+bjMQQDYzE8GJppkHZJntmcUxgW5RbmgEjf2aqHMGZhohQdbnp
BlauF+Ln/vLzjOOj4urnhTcALC7W42J52AtrP5XbQeZjRFpsnSKfxQPsgS8V
Tp1/zidwLf6zpv3JyihEkqE0VGJ1B3TH2yZBKsTlM2m2ogN1ybTH38jl+pRt
zQYpeHvP4VflMYb8T2mujdNQsmrFXS6vUejb3zTto63b4Dh1j7T9F2KGXaDw
HFVzL/PxwAHuhmr+ce05SFZzHfvud1lSqgmcGBQITPGVfzV9abfqRWMwE0vX
TyB42rFTu/pQnq8tZ4Q7VoJdPAdI/p5gn8/Uj7TCrha+LxBOn9k8coFkrNcC
bCi5OqhYXydU5TbaJ2DDk8mazPokozukXyF9bKvnlpXbwmWzWKKbDvnJBk9s
uFSLhmDAdg4LoYD7Vv+B0gJlbb2Uvf1oS8hCUeJ8JoGD7k7+wwm//dVWyP7x
XtKg8OziG7tSIGwffjZ/UeDoZslS58oVcsIwMN/f604RRNa7CWFLRkHSczVZ
Hdw2CLsWzfBZj0rXaMTKHjnsuzTuBUss2Zx/0qgvtJOhAFBOto1/PZBpiSOI
nK70Wyq5hylE0f2sUEHLUpJFXa+vGgkVkx+O6Ox7HnPXd6OjAnR5gUp6iOyz
XfzoT+iRh99unEc0NarGtJf9ZXzKhrG243STDVs6VQxHLMTEMUngCX2n/9+Q
/7/U8vxFshsLvi8c/UJEZEczHwdP24CPNin/kjNSSYeL5ymfqX4RwtLSq/X1
pfbVdf9CJ2S4PJ+PNDcMCzZzgr0SlC0FVZES1sUR3dkH4Ccua2G3I0KIl9e4
MvDn0jeZGDIFnAtzE7aNIlEXQc5PnkFmJ9E+IvItl4gJTggbioMgVnU2UwZs
l8+UkTdv4WmrANBUAz3IQbFdQOALpv9zXkMs8rWPZlG/Hsi2/hnD5jMDhvAD
a5lZRfcUEDu1HwuTDNwLUbeNMj8CGLyYdDTxD5CrDOhYgmV82ZyxLcCCUH1b
a7cMConJOECvgIP6soUylsjYg5YctP+bRTOHj7PywqQDFJ8QXSwe2X7GHhZf
58AxvDTYSIC/rkV0AP+iGi/AB2azvmikFz3nEasaZsUX5y3X0XBhnUIKKmLS
yRupUUaLyGq5ptAH6aq4PNQLaTBp7dWCP7wRauBeKc67PezBMNBU8U/HWG6Z
7NeIKVbQ5vFBqAoLOsb2WrfJSbyfuZg+JC/2WXkWh9apJt2dS2VqU7W7Feym
GURVR/ZUGS+tdTygDBqv+TDP/HrGYpRvcmJ2d6iUeOJZJQK/WScdQkd3Koc1
yCa51UUAormySxtKeAAR33Qdbjp4Kh1zCe7mftRm7W/nHUvazyyXD6nuCdAB
aAavv3d39ZVrF5JzwJoYPI5utjTkCVtyhL5PD/CDL3nr2FecroNdaBRH6Ha+
DbdaWil7GWmJHjVO9HA65uCNt8eJt+9tGd/IJ8JMA4gNeBKtreTjTHyXCNHz
VOE9KHnRTvKQ8LTeTsDPe3DTqzfpvNGfKXS39je/7fivPjIu85s0AQOH/HZP
rNcV44c1dudb43DQeoIb1nZ/C8+wvlcLyCRqviCS+97k/IsToh1MTx+6z+jT
jfuqdy5xsTUy0HwHtQ/A79xsU9LxzI1XiGm3nMSH6Ee7oE+A+vWsmzKz+l7V
WFDAs1ZqJ4xLrzvndjxGD/HpMjyiP3SmwBu/01nvVj91UsWSboiucfCJ+IZF
USDu8djaNJWUQ2+4ieMVpC6fEUMuwwsndjNu52Y0nckHl0fAv8WW5zxYNuM6
IOBW6apP1FyqsPZ2q0cubZ8gnw50RjI7zAq0CxrRQkNzbMxeU8jQ/Vp6m6m8
IohZJlgC6axuJCGX98a5Av1XB319CpmP0u3Jqm7drdeU3pejh3m3IgRk57Vc
1jjlUk+0nshskDy7ZnwNoPidpi0eba26dSCYilhBIG0F2aBo1BDWQaxlKuAI
Qk5Haos2dNf/U9h7meL6l4gWAHg+E8JXR04r9YYFS39gsMIq7OaITU2rMij4
HvrvDvlfjP62ilxM9y6h0tRcvz0ZCTXtvJVcix7ZGYdA/+jNaqYyrKRPvT/+
5YL98WOLMIB4WyRvgUTtDE5V+Nw1KLmrHqHacLnJ6It0VDZXEJ3vHrZPsEPy
tyZ6l7GA5cPLvABJYgQ1CCyZvjId6oPRIa+odgCmEy/5AANPeu1rr2iBYXEG
JAOL2yy2htxkUUrNJkmWQpDFcYn7RGYs2jeMaGzP0xTWCBU3izC4QUZiLZUv
ESDbM0kEC0pLewJEr+0JC7MjfHIGc9HuAXaz4A1c9RH7M5JF7rbAgY+7zXQf
Ft0BRamBU/LONdqOcxgyrlhg2dit/ZrWgum1jngVR1o28dtyYbuBksnJhH6K
Vkf9K+9NAJ2Pd7cqX6iZAiDEUW6OslyqS1AOHmZ8RESqrb066SlAfZxe10y9
8+7L0Dccovamsp9Wxa9WKopdfwfYsS96TTnGdIu0X8NDS7D4fOXcFUzFi1vn
iKzMam9SNtspXJYPq2/Jm2lMPRAv+QSe5e9Miw7QZv0+XBkD8vIaRi+J885F
/i9DYJO7drIYy60Jf3rykNWihcVYmdM1Y/cGgE4taUHSBCrWVMnURPNIpNYr
QT2advmiGsqRyaZweCDFIOThoXHst5mI+v5+JVlfn7AkFSOY8Ma3jC3OFwgp
X2ttbSCstoaIYoCcKG1VV9aUXZKKy/YK8s8RcPHXpCCb3SqkGDs1mshjTQa3
ZYFdmLJVDLLTedvtBwjzCWVMd2Ql8kaVfy0fR4sLlmnMUVRINiNeAm6laeOa
PaZ+y6KRcUp0KvEc04I+64E/D89NfrAPLu8AQHoZmXulFQ2fWsKvplJ3PbtV
FZ+axcNgmlNniFpIpUeNsKb5Jj/dJats/TGJSsGlIvYhS0ES6wFP+qXt3mTz
LCwgyZoGrXI8eWGTn9pQ6wmqQ11RNR0ui96xmCme30djb2SSnlzhNrgwKkNV
q7XCNk3xFgX4rCVimYRxPgT8c/o3UKDIKCM8MVp5OV57V359zxFom7HVZQgn
fGPDobrEsqZJqYympniFhHmnwiXEUwe/v8fXF2h7Rg19x/OsE/XA3hMs68hC
mfXiVy3A/+r6F0K1q0K8EK8qU+jQIDDKOXLDFog5MN8x2RG+X84bgUorlm+I
ChEWsSdF5nUARvoRynVng/UE5AA3dXpfD983MjwOLpuv7Hah4x0clrStPeAX
8EnAbGeQqT2gfwfbvC88vBx4Bt2yK31MJI/WQ2t6gR4miHG35m13B8/aHzHP
N6SDu5PxcFnEnUPWZ6D5Xr1ukjxhsATMlsVdQjPqIc0MAT1gJdLmxJ0LqakZ
8/1fZCvnxYps4MqCOfENKlewCaqSDwi/6SlnB5X1lnGz141S8E5XtZ7ECV53
19XMrUx6kr52cltgvc4bIc4X2t1LyGvtdK0M5AKEQthHQ7XMLSkfCjXjPmC9
vzUT8KRT9q7xA6dVtEQyydjxsTo0n0QBQnBLsv69/un6qC/jyGgi2fIrulFE
f1Z7CBGCQjx/g5Ml/X2rxht/70XQleN8TEXCmBPW0zIZJBZNeZzxvxrQMFpP
kbDYT9A+oFE6TI+lyld/YV3xa1VeB1vkYGMVjZUYW+ltMB3q8aEge91xC+FQ
YSWj6FiNp/IT7nh82PxNau4Ar0sCYXOZ6Z89f3aJBmx+ErTRGtAPdX7JWT2Q
1EFvimrSyqxiAIpXKzvf/52FnbwWi4dwGUgpzVxwRwkLbWb7eigUhirP0pRf
tZGavLik/tPuDVMZvIHdRZg0yoo7vsO2cr0sZMxhzylxUlYK9/WR3NSsTZXD
jZQbUTXevoLtMnbTBDcubp46C87oAkDTWiGAn3n5i8SW2ETz3iqpJbijuX0Z
CgURoXZt0baZ29oeWPcSu/5tyKjeWmVynKHM1KAtItWAYKoYiQJk3/sHAAfg
HZGIZOpe9xOrt4h3nTbNBNhKl3G6qbu1f5rCqbnuuAfOsw1hZNNRs9azU2xi
W635RxU1+gjJvx8yctp582KXwjabZoI1aKcWAP6IfXH3x7U6OZKxhHqf13Qe
7z7sWL6R6wkiwj03Gq1R0UXgrt0daLpLys6dPPnqM+qfGg95zT0RNWhi6lpv
pmu4UiIt04p1C+4K4pLCrcCwx7tKmWoHaUHaKgpZNbtY0JjiHOCMjxsF8UAg
vv/7Um6yXcp0i7s+D1Xv8gmGTG26TZ8OeD1xfM7r6Nt3yOkh5yoZHn9xr9Qd
DPKueWPzIo7huGeuAc2la31D0EppANccghlxHCddB2r5Io8obRJXujUQlqpP
fXC2YRM5Sx5pg1s5kc4Qzs6GZiKsPKvNPWJLEZT35CL7L+V7kwpTP3UbizoI
zQLPwy0Sqg8y7DagvmQvSRMp7ZeqP5XcbtFgteYPH920BXdvMULNjLrAFsm/
ToRWuTiPrcOdEIHBUluC0ytL18JIL50hkEX4085rh1LyzwUTgU3mi+S5Sfoy
GW8c3XWpdmFjDXGV03Wy/ldWhzbRrrrbfwzQDgbhA4a3jdclhngR/NmXS6UC
SXmpGUT8hVbeobgXI0xluC/3PzFIj30rp3EQDba1zZzg01MBVR45/cql0Eg+
BJaBvYeQLDBwZSEPbpDgTy7yl5/6ypasNdL7yyGR5VueKtvEFBEv1o7NOxjp
/8FbJYe4IyzPKo/cXVvj4vEsEBMMlPLkUJQ8qbCKcd9nV1LIaHGmU71fIg9o
h8+gauV7H1Ly6OxuGnLZSOzDgoBXTJqC+lw/NGqA9Kt9WWYviN18aCuZdZWn
Yj53lTY78Y7OqbfK767e1DHPSCUSq5AyHD0zB4kPOiyATATT7Bi43+3gwp8r
YgH9gz/PEQUQIJupTAhtWcKXSy4ZyhkYRRY4P6c6MacEGw25xPSo8vC1MR6p
JoVZib80gaWQYdkrTP6lH3OFo18YLMPdmqRSCxhJGNAlWloLX8XISMSF38ri
DiNnTIuwvzeIM2ZyYmDhjSbS1UXHU5/VV9/Pbhw9iA2GNJCefv+QMdplsr7w
qg9/UNHWVc2Ta9ORww6gXHovmuW4m14ZTg63HFtULl6SHpxJW/o2rzAl9zdm
z549OvCsftLgVlBmjbUVso+RkuMsA3YojnaUvhk12MdTU8/MZiMI5NGvm5+1
FxdMqd7BL5Zo4q52XIygrKcQ6dRa86rJXrYLdWv1Gamvn/rIz1SdtknneAwW
AIwQojd2pDXeEhahPkrhZmbEKWW4mEWF6O9S4Peycw9ppBpbV/D1ID5SuFXh
Xny1tmLYKxwJCSR7FvHSjF2thj7TFSqX5YrRegNiMiyz1lzVBpCak0uAZUvt
Kulok4VyH1lviLJPpOfjZXoDBIsIHKs1/a9K9zEhe5DJqU2cPyHMTmtpJkmD
MTU9UDT+P7GX2V0oAdAs5BQ0Dq8IR4/RwUeR64WOrtrD27SnRvmayn3ytDIg
UDKD93RvcIzRN7NYv777XKnNkXeh2rmlL7f+VqaSamJTtSZ2lgQy60uhQihZ
SLWfDSymcLNg3+VvklVrzemqzX9VCUHv5uCuALQcxXIvdIcaMARZKyZkVs4q
iYJlwJwXEfJkldbM8pnLq/ZTARxR6x9+JgsOgVVSuAgGj5fC6hBTe6vSI4uV
PfitqVbAGAzROqunjKTxK9dr6OqFZokRtqGBqKH3oitKa0l8yF5Bx+nGKm6U
2UI2pCaQ7crOmCfhC3BnRRcAlzgsfMRCEHWUBjfVBVHq8hO1MgK2Srb2MSJv
NtHPanRwMQmJ+ZhUu6R3PDKkat9OWl9Ov3UeXVudW1CGfJHNcHHs++fNRrby
pDlNS8an9dhkal6w+uGxfIx7eDIUtWTs+9RQc8hHQYSg+4uoSHXwvVSNSEqF
DxRVKIbMBk8SCqk8pOEcIU7HfvQOFnJPnaKU+DofkE5EsP1pwLPvkpRNBCHf
TI0gdtuagLjjdM/yfU2rSQAsAXnTnzTdn7hpyMBrrvVZMzG0pxOJ5J/1oMnC
1aPG+/lyrwtYWRIW8XfMk4Q9a5O4C93MkAVMQeqKMyU+w2zhXsb+z/d0n6HI
IKdjA4gbWI4eGdX0jNzh1QDaNWNfJEQHr6w2dwlJFprvREUMtXKwatkkcPQL
/OUGyR5AxCOpKg4z7acq+6iXUUKgvX9qmT3wtNlq1oZsGD+xVKxH82HXh6Rp
2j9a1ElMF745OCW1VvZVRCDk/rkOZFCGRkFhlwa2y9tnWNwyRRuAt5XdBwTc
Kdgwxp0Xk8H39njvXufjz+zXOmQiK8JGHCY+8t4EKKlrgiBnooUCGTpBJIUG
2UIhLuym9MrbWyiBQaH5YMBqc8hOLEDj8LpRaExuVXmSO88GlrFAO6swKCKN
2SbCkBJuRHz0E0IPJsvRzJ9cU4FaaD4eCv0MLmSnsi5sQEYYBKMp/GQEN19h
P+RfvkDWFYMeI0MLAQblm3mbgEqRQfkWZugqSEWtu3zQzPb2S1FY/EHWqr7C
hXxNYV68N/GetcbTXMpTsw0sM3qCnD04lBxXP6yIABy2NoldO7C/saewPIZ/
JH+vIRNSB0PN+czlf8vLMP7tJjBEZuKrl0djeUs+YowL0Zo/mP/aeq75xYS7
k1CQWT6+FsvW/P3sKz+ZlrTH2g8/xm1vPeyyBNQxd0wyp4QF11VhCL/jT1S2
7MTTppwTs8CI90zDY7lne0HROVtfoQmMEQdDdsu2zArQxgrry3rwS7grU3UE
la63hmnXE3lfbDDQ/Q3O1gxrq5v2lczKCuEBKDv6K9S10IWz/7zFoxAj9csp
nlpFMa/DvkOO3zkDWLZ+BS3Ct9QE2Tc4zI3WsM8NefB5+XjTkXYEWOiZLDPV
U58mO/daPeow2zILvL0iEJQenbyV1LrV428MG4c8bvum5YMof49e2fiXtEUP
A+rrTnd1SJjhJjqUgQLxMgvnWXDrF6khZwtsoE6Arr9zUgFGnBvbg6FOGlUz
xcutZOS6eKy2nDiEalnEkte+pKCMLF/jrK9U0Cjzjwa4ydAvIFy4M3rffTDb
KNf1V+0HesJDutvI/HRN3LodYDsEZHMjVU3Q3Z3p7CfngiISy+HmfIa2wmG7
1rsydRuY4Sc6f26/RXlxq2/pptPi+uTjGLphAJJC6AksZ+i8IfF81CgFpJ4j
GM/HBjk3TGu6+nNJ0JzA3CmZL+LSuYXZeyP9tsPVeTjupM221UesKM+k6XLJ
imYIVV/dZFjh+8EBIC6dsvhE1CgSQ34hX0fkgyLeqdJD2+t12WYnI+fN0yBD
bwcbSYzMzMP5gZmX9FIn/5lHOinAJ2M1Rtb2mQy0ChvQubqoZVtTfAyDcMmA
pDWNtQmW854SzdrXH8H7XikmNrsTBtqUKyMbkK5VJECkHhg39EQ8d9m55hht
rl3+Asfzm1Pg8Qjr0HmOPTPdtTzK5OJxEfo1eGUDFpPV15K7KoLGD0IeEakT
wfmoO8WfhxZo1mERdBLm7W3mGNOVnYc23MoMpU2ivFGgV7akBRHeJcENfZX6
W019jNQ8DdBDDtevd3xaDuSKQa8abigakE7DRtWbpuSmOIFqNrzdhzRdHgo1
DEjAUdcqhjU61+u/QnLJyAtVIeyTVojkM0vE4Vj2+jdIoKUzI7nC5jfdo0zC
TN2zpFvMrEW7pkUj+qgk0GX5F+7/5lxGcCo2fag76fdDYzVBv1d/ksOjA5nT
Mjvo81J/+cJR2YJOUhTJ1fUSQcMcMMUvUHdjuJW/jE59bDVblOd7apPuXCuj
7pRRRSS9iab4NuQaFAKLKQXDi5ql8MoYHL7ZIRelEZYjQuqyKkCXqFdIXUbj
jbYZhYYjMl6P6IjUSqH4nEeikuR/Nup3fKkarH2cxGjQuO3YkhZUxV6nI/YK
ObnkDyuW9GZrR5JN4sR4L1rUD9oqFH5aCddiVdlVMbGzpv/IThSx63Yta1tw
w9WivqFFMuhJMMYHwwLfj3owBLgtbqvQ9dy6+fN0Af5br+GuFXhXEH80uHJY
LTnCNAwrQ67dDgEbA2XZkaK4kAs0lHwsOeitzUaBRcsHe+mJjA93JoM2Jdq5
q1wCkaHrcR7xytnjiH9SFCUIhMTIe7IeRPFvfIDYO3LTEB8Tie5zYj1Dqa1v
lu6uH+qMhkhjLmRNhwbBN/nJL5pqHIUe7nSPO4uQSWl1uKECAYwx1n4fxVhh
d4BH67ebowj7rmgrLVzqBz395neiosq3kW1vIXO8CIstfMC91IFhCj7J5VzX
BBZG5ETA8yVCKG9V0RcABbSVhyX5kHNPqvaev41bJKX9OyXE4XL84zpNc/1T
MFG84Y9JXBQgHerIfd0rdMftS33W5XnPXYs8qOl7yuKwHHvADIRzvJUdWMXs
Mu5tWtHSl3Uo1QOcoo+Am5GS8Pdsrc+pfg2fKRrs8wxDcTU1rk7MWN7u5PcV
UdurdPp3fxT4g/oR8SxxeFJuz4nLYOo8jhH4jkpR/bM77Y3gYKGUu3Z8RiKl
vftw0IX+CDoK1vVNMe3cf7wiVNwHZaMoDwvtR7hFncJMkNBSk86/4KYG50m6
hhCJN3jN+dT9QoubtfbdfgU/9DLpmoqhX2yem5+WsrUB0DNdmu+KXxHG7UjF
FXIXqfMDX4gsxzzEbo1WKMKMjsKK6INUFV1OVbdvGdpnaTlXsbeBsLgN3A0b
k0foHtrjameH81+MsGA/EIg6bIeJ1rwAzMelp7PGqn5aEbxOjF5J82M31+uF
HSSNDXpmYq+Wk+BOjWJ3Do49rGMJpOr78XSR9AJzFG8UwVE5kODAgapY5Vxi
z0AM/8kQ1FlSOd5I0O2lCGnykJpk0MtdQYTfNiPZ2pWG/Cb3YmwSv/q0tPuq
pIs3rD5toUhHcmotAVuAUHrekDSCwXPa1gqQArfrTPamusmC0LQLAAIa3UPt
wuxN1GhT7jKmqn9thtyYjCdHGVP3A55Re8EFORbujWvT5oe/6spxxHp871z4
5WbrOpjHd1Nyh/LB/AMcWDurblVHCuU7I0+knkaATdrGegwlGJHFeNsVSy6L
tgIvBevERHRYssDJeb7N7lVEWMDGZlV+F5RgLGQM8Z4coH36AT4BOW8S79wX
+FsMPpSXMONUJJk6IsjvLW3urB0HIzC7VJusnQ3v1Wz2zht/Vj9pTUHpC35r
6ur9xY7dqLHjg4j6km9rY7Gn6ue6FsHBD1n7kcXSdSxdginRT2vtWuY+/F/g
byoy5zzVwLfxgdWfWxjfUBLyzdZTLuhwn4Lx3rE/1qn9WR76jcYk2CrP8eue
ObefU3SY5lnGE5M0tNegtQoMc9zuZmHSntSni/7Rj9RAJGQisZxRXo16bPH+
zvubf5DwR6izQPW2V0hR2ycahW/lGUbM71ABg0JuE3eMkYQSFmYp6eBqUuYR
w3pvO0VTPFUNmFUgFt4dT48HlRvvknZ4+x0dYhuVmntyaYHiJRi8BpRrgyJb
HekPflmE31U3X4eELIYWqyfxZ5vwQbjvJByUl6dY0qF4XHE7wWQlEowHTqDW
16FV0abzPYSsZMehRsGPWo4XdoZ0asTBW4lYGp5AQ8PcDvfqqWs3i9azLeI0
llTHgZbEY613PFCIP+3Afm69WGtFP+D4vLAl9HhCBq/mRKYO57gAL0U4/eLQ
10m9tEI/owke6OFtXN/leN4L0+ZmTaU5j5qucZbJ3GR5hjfjhkKqKEE0Kymo
/UDQazvL9TVmiGr/3MfAAyjYen5g6JVvN9STwumXBqmtQ961DIy/ue/JYVG5
ckXc0AEw1ckwVkmAfYEa70tcaQM3upcgIuxjN3tNWmZYLkX9m3ZPTuhtXvWj
45IzPFR2NoyvSJQdMLQeF5iDRDMhdsRaln0ktM4LB/IUEHhXV6k4mPC9cm6R
BHRoxo6NQzc2/GrBR7WoT+i1dx3pymaUrNLUHRHhk4VgBg9DZbu9RilQxrwu
O3H6v0EKHHQBcpZgnvbALYmekVjKqVLB72vvFi/mz5BZKgAay7/AsTYz2YRE
ST3u/zSj590npT8c5x2hReY0MdGi1kicdqDN3LMjBhbClEUP8r11jM3EfE7X
b59KMEtVhjFeSfM/sVPvgUvceNRElaLeezTytpJ5uf5VUPooNNtL1B7WB473
7YSU06d9efmEfcPINr3YzMa6sPegiqwFzNtGOMimROJ0JiKGlAL3pigCpKBI
SHTZRoPat7i3hnIEW5TXLDKPaxKLPtXn/uCBB7ZiUf/diMtrsJH7VBNqc6MS
q2z9/Wo3pSPaJyo6YtbDr+pZV+MvXSSYK55z7QSfQ2nif7RxKbj49PnjAh81
g8adSCVqBkpTfGQjO8iTIvlVbX+M3ls+QBoOAiXwiwpm5WoDaCFnHgZyIPSR
m0YsGrUJgIqVJ/5SoMM8ww0Ta3wRx2oIUGEy+MaWW1gTLtGLa073rc7bg7o+
t25byjPK8Waqly7cUzkWG/ODDGP+EPPbSCeWkpAQ3qlTiJebCk+jpn3CkP+8
GxPu09qd8A35fDZ5B7ruqy3Sx4KpOOqDI726qvCjdU1wmEmmKDmRuNHr/a6g
qJS08bWlmX2k+XLOFlyKOSj0Fm6/k09tgrAtEwRBhLTWdwYP8RM/V07rILzp
Gm0vR3vekWLoPkT7tJqYhNAPzpyVy0CNrhaJs0Dluz2J3P9mEvu68zuZ8z4p
EI0132hX5ythgUW0BzYbONe4WZwYPe4YYg3fJpx32l6Lt44DDlfE02vWDIGn
jnf3O268UV0/e8ilMoaelad5tEZ93m1pHoQAS7F5bW1Zmk0ZyBWY52aZmXfz
ZHWnY3tfNKS3bOkVCppzMAvpeqIdvpVL5xSU9JWMxmIeCd+fTxJDw+IltbM4
8Rd2MAokG6XSCvFQ/poSxejPWg7FbrMvPfr6HxttyN0HXNDAhE5YqrLqqekY
2CpNEWBWn6RY83OD8nAN7lVW11IWNNllzSG2yK2ZZ7qs2aexhLUkjYFvFadp
FJE395sGtWK1e6XOprhCXUyH82Giz2yHvoHqoQsoN+Z6YpqvAhl6I4JHptze
0bNmh+os9DXNqI1assgNULDGnLJ1H9i4X+AhfKkBlPCyAvT1ykZu/EOBi1RR
AE9ln3M4y+/VLajqk/MzBl71l4kdcK1QBUp9DNiR9OajZi9eKL/BODil3qQW
tcoHksLUUxNcpXSjkQsn8SXuxe3HwT4RqIHj/L9SS+ux08CUk2Odvei0TgVV
8e4UiPP+DIlC+j8EmdYNUCRRi+XjJM9h0V9w+QtRJgKfjRCwzWOllUcAenWY
401S4OxgmKbvjNa36fHrStm8Vx9jqLZPz6P+rJxpGw0wWq+RpBV2xiQKZJ/A
d18c4ObTrFI2ZLtKL8TYofIGh0cWO0lumyAHgcxDh8mv3Ez2PgpwufrHiczq
edtvhhFlpAWVPugU52lJqBxELfhJT/rmA1vCnIxEetk3XD4JmjO3ua7khkio
nc/UlThMB8FiAiCmeRgA/L+MEXqU1EcG3Pw0pqeWk1LDEl+87lVecbL0e2F8
esqxWZCsv+71OETQftaFmO+LqCQ0xzUewBQZYo689CwHLAW//IV3bltTdcTb
KUwiCEESX8tIkeZPwBk5mm3fybNB8ZsjbK7dZSxYtxJbdyWE4CyY09y6gWQW
Oy+BfH8M2AOan+RDCAlVB9EVkBY/rXLU6O1kIcinlE97Ph0hAmr/hUHa33n+
ctekghEMk+n6xGn/pVMPoxLOGBsf5mlkMQ5WF+hBopDV4/PRmeorWkw0Qwqu
OOOwiwZFUoSbI8F22+z1FE6l3o017edjBFbBmbuBpKiwhurQl4n0zuSpjsT1
VwCpZqk3nM3Hd8KTHLKXWMIxDcZEB2kKw9rk2bqrjA/q73CGbGXloYi4QGuL
LYE593MNe0VFcgGM4HWByNgs5TNuGs+xJfbO2a7bu8y95FfTKTcH7aD8kQ3F
4KMJpjDtkQAyy3JRsgm+D838gLWPLDklKDXevYYAYoIMkIjF1wJLzWvfJM+Z
r7nlDEdpXs60MaXEDFZdKbmLf0A8Ff2FrBB34YJQxtiIC3ylQ4auUa9plQQv
3xfTo1FWKzQZBoFoT+8Uyn9cfMaGZPeDIR5HqCxmJKz7L9tMEQv8btb6HZTS
J1N8afT3JNYHtw97MYwb/UF7eFQm9/zv6DRW99nnUSnbJuzZ23PpIPbwT3QV
RMFy1LIdXECHEcDkPaPjW/ZGYsRkfBaNUDEp520N6hc6QGMLeoTDBWI530mX
jx9EqJL+h4RG1Q6j1t0vbqsZxtvSh8k2f5GK1nexiiywSjEMp70w+oTioA/d
x1tC4saWtWyI6HC6J0xXcv0Ywhk2SDMeQBiGEzepl+9V6ZyOwd2lvuuxvGY6
TLbgZpC0a6UwfSc1P82aHkeZR/5OhCWP5ex2XKyFcuoYEcOvunyp3Cb1ROw2
rVKmVve50/g2HQLl8OXsIcxfqKM8uz18iuFY0CmS+x7Zg84onP7Jq9CLsYz4
Rd1EZkGX/tQcS7AZGTXa9/QaRXef12788JwrUDw9Fn3NgHMs8RKPMB++bzmM
9LGxVnZ2izH7H9AQbboiiqqmWb8Gnw4k8i9Rrf+oxKa80y4t0pjzK7PsX6WK
JEj7LWbSlA/knRtv0kI4V1knMh9H/ikAhQq6WFVq9FC9hWKR20W5rWw2AHXp
LhqDJjsLlQRZjddvfIyoF9XZ2rCZYyz/xrhGwOgkC8MlegKlxvqH/0Re6iKF
5OTsDqU/YecArEMjPwR54DPPUfNrNmBCt1wCXa21+HADNHF49v43EK7ovv9/
prwaMrME8MxzGkbb4nbxsNQi9jEyAGcMNqzzO5R98mY5OnsULS6x0He525iH
7XwFpDzzcB4K3lYabi7VkH7OInlcGwDXQLWnOUe7pQmOmc4DBNJi30sUuHGw
fVBeN7cwwDVRXrHj5F1Pz4NVejPlndTgrX79wJRFX1hFdc0/K3YKd/kAI+F9
LDC0v5WQKMCIQKVXXAHK3djiv2oW5aAnpI6FUWmAzJ9xhQ/Vhwt8X8fKIThu
o2KRieXD3rW2xcWwLh5xkic/hsgdy4s+a/oONfDl+zZ9cmGqEv0yWTCVfZZX
2dc/ZVHYZPqn99SwffHiXy5+asNVa+az3jJSt4ewJ7hSLid183MMSLhCws13
gz/LUFjMZdqVp78twTgm1RS24RN4IhlAYpCl5OzlHdCcovSwusYoFMqaqCGo
UJ9L4lbEFM+FNVGnzHxJoMvqMPEzL/2gnDvsFbFC9aPRw1+yIGlW9jMEFO6O
S7BI9ZAuYSIAhD8BezdWMpDm1e51/Z8jEXALNfdc9d8s/V7utyHvxXzPRKMt
jWlMuwk8e/5yn46GL+TzJohoqaNYvEeNZ93uxMCC4jR7BA5ew9j6v4FVRpLn
LSVpgonAyreaD5qEsrKdBj/a8mO9q2GjZ9a8cO3WhcSypcMMC7vHx9PpsKbw
UiYn/71mtouGpuuP/r74T2JwVQXvjEE9ftAMvO7pjhN2n7bvgb4hydXEmA2j
nQ/UTSjGeqETdM49nf+KojYE8uGDOdf0Rr6fihki/gPz2Ur0Zf9uLhhJFyGY
OcBYW+5K3nRV3x+6MmdtjGSVpYPYLFLOuwqSy5lQW7taqzWTx8vadEOGWo+F
yzVvGVtUPwKss1xchsDqdvii2LvbLAvw6iHeDpKp2PyyKqZUEYnbRdmJgKuf
Wu716cHv3ZHxUNHCBFR42hxnNCOENtbuORRysPpSAaCoccK8MAimFku6hJ3N
MOxjoVcFszfw51tTMYulnRte9SbaLRdkcXjqE4yJ02D6ivRhkmiaBOcVm80P
Bqgrj6O2ST/Bwsb7ElFrme1Nf4/XKPEZ6PYp1ZOKLGwzSrLxAFuU5dCqwcrl
i3L2qxD5I2nuZby0jrcOCh6CmzhcnJbJ9tNJrIBz5dPC3ZbB/Q5W9lJFlj3s
vCkr3G6hf4vL7vIhsn9bqdalS65dj5+Z4F98C/Ee8d8tNUP+WN0kjAY9vAxh
zF0VGoCFBkiiC2DlEaWb//nNU7bMVF9GMsMCVfuLYf95UIofQf6Ubq4/olxB
b5ostFvrJfhT4fE6+oY/BexrJV8EjWkbVK3CNSdQeEfjjs8TTSf9I1LzplbR
19up6LyO/CPcyhUt4eUybr9tqCV2OAAxHvmD2szNGc88k7ldQi4lWlv44gGG
g928FHP93XJQ0vjB8CKyEF+Eh/5oIbvoCBwPuYHSAXThSYFkWumiZGDwqVJT
MACDxSPqQFFFE07h8ASxQD2wcRST7r6wBXUEL3WDYBNfefkGLP4HA4FbnZt/
jMqmdpw5kHi46RGF6yyklhM0yeCyVXl1zFIL/J3/MpFPC4kjukIeKQztP/ZN
ownstEcErIQQ3WJC65RQLrafAKLPgyvp48hasol/Cxxs9whJBQKpNgEq3ZV6
scopB+4UosJXLqS9DH1iaxnc6TVYmkcX9hG8NwnpeX+r7rzbyDm1CNpmqFXZ
AxRUxTENTncIlsA6YbEClXXcs3U5Cz6qlclxWrvvJ8i8Vs8KsEy23ngV1VKI
BNW7C3DYVteyR5RvibLbdMjsdl2yKPDvgDBnMLpFY1r31TY73ZNZshRCAi2o
25VDuwlNvR2eENgRSXPEv2biZ547Fy36NSNSr7YlNGkLuDdTQDADCu3vLdCQ
qpKiRwID3JChc3Ypntbih8koJoXz2Rv2LBLkqRjtHYaM9Cc87ci8Sqk3lEUt
G6L00EfXSIJdVYnH9PRl6zVj6S4CX6C8gykt/KztuacJ7i5FJ7h8G1T1mi6T
0F1VTUdXYmm58QVOFM+Pdp2JuMCMRgxpJA3GXq/U3dTSZU+/I618J4Y6RUr+
mB7Z0UCbdmlFlFk/C30KaCB6esoB2lfyLCD8TmxByB8PKqor5A7sC2ztfPXP
qktc+BqJmLwJM2vogbKffVI+W1yC9K3MfoLvHPkKWn6WLxRnjg5cC6+9xS4J
VBvnheRYoQsC6D9zX/XFz54Qni3Cjik8tgYKeYP3fwGwXaAHBagoYUQ1M143
3RBaf6AlJvOkS9FJLZXwAxLUS1e1z1tkd7z5dV0V/XjpsjEI+H5p2evEqdLz
Yvg55WNxW3KD+sqkbk/oq0UzkfL9TtoXg0N216rNh7rVNPJ+zaQ3xJTNhh27
DRP8EBQKfZl8W7j1uWJIzU9gzzsoVzm+fx93SWibAClvhf0N73KDSC9YYRwk
z5fqIyTnDpvMVAspXChVYXkEBJHOxAEK/0eipkyxwv1OFLknichQhwzrJbLh
MOqLZ89dmSUddoStErQ2nwUwTKiFxq24w53ABQSAEXUDvNes+27LvQB53L4o
nX8rfBInxwH9wwMPDWIw7uJt0M0f6E6Wd8Mi9iGWrRKAeOmaAF/YPzjuPryp
HSzAylKi8L8jTtTGdNplYP11K0ZuQwLvcW9tfxYamLXtmrX77JXXbV9Gro5C
2JCig8Ct40GxZSl/JerVl2suSwl0Fq5HeKOUkh9orKtu1VnGDDhfkc1Xf6ee
r9msI9BLHrXcdbhz0wHpmj1fD0qH9waMYGzx9AaFlNCnVKY47qZnQacdPMa7
AMxjnmpcpV6iYb/8DtTlahSQzrgHoP9TP90gWA5dalBYzj9NI8SDXrldgvKq
lZ0uWImsKCo+2cRsAqqrzx5SXeM89YPvhz1l0itarKIG7NQe5t2QudPv41Yq
cpTpJnYmCFIgk3dlDMFphX41QAStL0TdmJEIJhTGAgtz+sFz1XqkBh4JqqIz
wSv/ScArh3Cqhya6afrpFSCIhuWlnLCUDPkU7rABG3BYKHKDrfoPmFQhEURn
LIjlG7mJrhC8wpyOsnXy4UO0LyWFcEcS5nw+CyHZN0ll8OnqEDp8ZkEffRdo
4jwlUvkhBLn/XaohfvXB9CiAqpjH8MhbF1yQGu56IT0j3HvpJiFwDgtTRqfn
7efcKYWsp+XZkY5r2qmn/M0YpY5BgpPJgtF7bJI3nf6dGYDO7u/C2rJfz72t
43z5Fr1RsiY6FIm9IZ0GRE++s5PEDCTO66ryO/VHRykxEw9QwXYAVLjz1Peq
vC7FlP7Se2eo399gyXwG4iwprkCNU/uL+IYPvSl7WIKib6VdmQ51hohQNk/n
VxpIq73h+7BSmGXCZp4j0qJ1uVFIduev6Vv/46mbz7cARwi0rb3Keg+WNfxd
F53hvpacd4kIRwdBguLDyUeZGrKN08bwbHAN27mFP0ObNr9HLj40pRWkOpGH
TIJMWJqhgjAJ0yG7ksAJA8yxfoe/6b0TzgalKXGMPJxV+BVCNzvtgz111UkC
33+uZoalCRZctez32nsbe+FeEQjjc27MZ+YiOwR7mMWVOO0oau1Tf92u5jGW
g0H38cNsFVtpX3/CKW0fqnGUiKBvUmS13SHJk3Tm7pBNMxWUHbN9aGNvoMsd
jgsR9jz5+i0pviXsR89rRy6DeaqX8Rov4aU+5o2xMhJ3zwjK3rroomKB4WhM
nTv8Ie7DO7MTBN/ccpqrtr2hbZmNo8n/imOfBzZpc7JKaZP0MItgzgBzlEXO
1UReTg2fzIo0tZettKz8UMUa3PEZ8uLw7aHkrBnnUez77zGp07V2lI69ScVf
vusRJDLCsccgj/lY5ptXEzLolW1Vvah9Q298ZaRtmSfpl2eX2v7uKHrmj2u5
+irTNPy8AXbn8Kt06/Oee/lro58C9IB14bYn1Em7Ozil0vgAbMYT7/8Cz6kc
sVg9Ql8dmKvRAewpWaGh2S4lw9BdZy/7/BoCp2lKWG1GtFoHVlXQ0UPRkjxO
alE6Ks6Sr7mx57Aumi2NHFk8Q661UksXhrdVopjJ8ANn1iREVm96d3HeCrqH
fUKcKCtM/zNu8w0uCybcWn3Ulxz0jdp0qoKCIgIkeTvupccTEFgmnhAAyPJk
O1qVcKxs+lgFXca0GW9NQNEXNXk/LaE8uSQ3YjstwyV2z7FknZCJFEZkQJCP
e6ZgjApyR6PSFP2p+XEvLTmiFoPYtPQZmBXPAx9n9xZwf44utI0EQV+jXEvw
kOqFYGG38PiR4hGi3dUyC7vvpmohkdUQUjgy0Y0/ABRq/S9PNgMZRmCsTf0q
iknseecPbSV3YHNfBjXtzqgutmTh4BCJuETcZoMOUjd3hDJw5DUDuc43Hj8+
DwAAMrADctW6mhVuVHXBthHhJgHMfGoysVzJFBR4NUAuTNT1WXVaTu3Nj1wf
OQVCKAjbTHeuSoD88FEG98yQ+d2VwX0MDVL+mc1HCGQH0oiZiqaIffgVMth9
yRZUyWt4sozfhX1PSpVLz3Wv7EwW6h8NUzaYvN59oEX0+UWCmYZ0Huw0MIyP
OMPX/spPdsGc7SYx1vsNy31yIdHn8EzhN3q0GyikL2aaUo6LIyBt3kqc6U8/
Hseq/esXrBOo+yUkW8jUUofZlgJuBwMTvilvsDoZ62UcqrBBarNx1Gg2s6pA
zwBWaxov0pR8gCcC0ZcY3n7RZRKCwdFAJcUbEXPiPs9s4KrhT8K9Wdtwe929
FbIdi1dr/0k4iSaY5NwaIalGwQafhZC+PwzO1QvU3UAcIzUIeBFUP7H4jVSz
seNfpkne3wHoFMdVJqDn8wuYDRYXlAP4ZAAGzDvj3yf09MuFDDWnYq1g97MJ
7kJc2KgQct03zc1crr5wxUl9tK9sUaB4dbM6T4l3R9U2bWNxki1nTi0EeadS
LVC4mWY1WhyvbecTqcTUh4Wembe0BFq6KetqQjXrbUdduejMsARp5YMA4kGH
wc0YaXxEt/JNEyoDGYJF0awVEQ//QjL/Q/giHHx0e0pIo0xtpqGlDoJuOiB1
ghok03/DK49llodNoUMAbuzFgvBwQrmXRMzucwhVafCeFf9HwQSAYzHt8xcq
REzALN1slYvr4SY7Y7zUrw+fQfVjFsFrwYMb/cVdaXkwZmhFoTQEQz/0GfQQ
LAJkL+fMN0geucbEerGC2Wnuay/RQtpSpi4XnHsCdGE6mpWAoJEg3U4ey52I
cyjF+LvKh+ofX8/8xWLUKjnmK/GzPk/cp1dTbXsc8mKo18N7i+llhwKVMpio
tfQljcevOxIamh1T9PMwtdHPuanfHu4gM28fg2jf/dzkhhyBPXvnTMe2GShN
1MbAGiLsN12ce6fHPSf7ivE5pWixmUlIVAD9G2CzswChSOeCJSYCTVCPlRac
MZSaOAGYEibtjlcR7XguBqBobaKR2pHPYD8bzTk0++/h2SLGKPaQI6OXhrEd
ZCwLPaKAO4NYduYYSdnNg3UKk8MouQVTAFXgdhtrToiLD/hO39Pub1y+piph
ALgQD6ei5l88d/yfU6TQdVHVJjym6CvxlrdpLewiTWCX9SVoSI/yYu2HCZ8H
CKDWPEInthLIj0cAG96sRYGbWKGUWySS8kEv08G4OoDGQYMElaHlpck+0My+
a1Jg5SK0MWkA1UrZualSxGaQo+qkLBwSVk4+ADZc85EdlQHoTkBSMeSszdlA
zVneo2DRIDZe8ahfLpoNZtmUUMeBnqKsUA6C9OMVK68+fY3MOcFvlGkNeWnN
/0QlBFBVqaWoxQ0ay1hgVpvoXVx+aAQi4zEmtJoWrwO8/rqqzWN4mrBsNrew
0hV8RFR/AiVTApTPyctxagXaMaIF2Fe3OZHG7ZoPVxICdrzpvdb2IIX8PCxS
x8K/x9g06oLr8NaHoF7ogZOz7mYpurxDv3cxpxmHdiH6oWPV/Q+8xeP+Fq9c
GTQ6Cb/cRKK+C2TlChS6kMX4hFQVtXq4nXsyyqBQ79AQHjk9N/kjn2ze2eZY
/USnQGpGZTdOqrQwMmJCTYI0x4vDQfMdeH84nx5P6xEvj5TKCwlHWI4ERzYh
1C/VMK06+1U2vaWkiKZI3SdbhF/XUIoqAPPADx1r0woaQQoXLp5F2BwsdQAV
L2ben3I6xms9Um91tTPn1Yo3Qkp6PkKWe5AAWlvRmn0Ru6Mm6qrFeN/BgvQf
NLAuOzlZtLQZhkQex4X0fu1xsEiD+RLClmORqxAySWhKpLPWLgjae4Xu3Eep
JR206T87rDKg536ZK35RBV9JsgpRpx1/mjYiEM2LQsGe1TQf6DZYru+6Xb3k
ZKdXLf+sFLqToXP+0dvvqg/GjQSk1Ngmp0HZGGL3j+2SaVXxqGy7eOPJnsnk
sBXoxH1vh5+DB+h3Qoa5H4XHbw+6rdM3UpBjoy2O1daojEH3LW5mhJvf3iKP
Uce5+5MleT1GQayiozgzJEP9adx23uHudnl4Dt4PJq+eREDtNilBrlc6AX3l
hcKnZ0poKNYkRyciLbtWGiXrKFkDDScrOMuHSd1snGCJXKwBksh4dTcL5QRA
Cc1Bz0m4IqCi1/cepMjQZyDqDS+AsjFyTT++x0hr4Pl/DF9VkErSlqorM6C0
/+ENgFl5PJfsbdy9qJC78E8j/v04f1i9lZNChnN4IvDIajhZ4oFlSdHByMz3
JRrOTr3Cz3rjaXOat+us1kEuaCeC6gGAIEfdrQFxMb/Psjnt5qmvty2rxm20
5pc0OKmbhbl/qnyz5t+q3cxLHP4N1GyfMDO6JzVWsamOw7MplBbg8lq2RXOd
CKclyQEOhNhew1KHcvrrpjN1QsNh1XXLGSjJAxxeZd50w+LDgjYH2yI0vfkV
loiQ+SssfOj+PEGalL7VGDuZzLG/7JaKAvgcyADfX93bmW+WrNz03ReCiNEg
KfUoHyVjENQM+ijZ3CTv0VUOztVBTD/cwWY0WoErAFpCI3h2kLIyEUBxwnrV
w0MUm8RZnVpjrhyMuLdjG7IiraaS0NAR92l1Uz35rzOl1ysSLpXcv+63rskl
LxotswmIcQv1fHxdOzBjyNSnYdSHhWuVzQmbl5dmgqfXdpHXnncaEbFteZq2
f92qbLOQ6O37VyeSx4VUjrBCXSR8gIlux8yTZwB53ayNtRuIIm/6FPyvsqHL
p5mWCMmBf2XWutO0DD2URrzhYsj2q6lM1z5gbs5S5471vu25dwtEIzC5Uf7p
kUDKsKVGaqkUL+p6bO+5uxiT5Rqc5HxKQyRBHINSKcg35DNepkNkq1iPS0aw
FM//ys18mAKVIlmuz+SWOo+tJUTH1LLsterfxDxgHoRkwWr97iFgWLax1sIM
GHLweeus+kcnEdvjrc0VWVClvq7XQCkmAkAcrSkc47puvHgyY1Sd4bY3Kc/h
0nk2hSopAzeoXTctsyefFsbuXw8Fh1D/wXFpOXBYPyJIFEUan3hUZk01Vemx
TQdr00/7QJ/GAzISvO6w/OTO9iJeRvRIOXcyXsHjZhjmwZwVH233m4jwZs1c
SrnFuFgBnwmbhtWJYotD1kTBFBXvZ7GFRvnI4qTnyyuyFFnTaEHD2KQu7e9c
NJ68LWmYQI/uWAcTadr7G2Udb/6vKqPN4aAp3yQFu8SBwNSSIEtSx5/2FPtj
87lnKqWdzFDy+IhxRGpYEzNhOjRhTaHZfLVnCyVnfQ9vRQwHhOZENcTkohYc
0JMVgt6X41Hzl6ttL7LYFsNr1QugRIvTPNdNs3EPPafKNnvOadDf8ds8mBF/
55RaikptMZS4i1UfNXH5yeIoIsFflN6rbV5vr+HiZBOr2PCR1rDrsa68lI+f
H9K8+AMeLYZJykckztMFaDafMaq2aGKoNZju+uvZc+Qi+qEAgMknOO5FfS5y
buQ7e85wDFbXf9MDyEOIoAZr+ehoXJI0yZ9M+2z+dAa1nX30DCrq1YzPanK0
dsuwjtwxQen9xTml+2Ue8V/9+nKpe6zrMvLWjCbnAZtNyjp1NsdmBKzesVVh
xV5GlD4JKq7QLJjQXVxG7sBaDOugN5OgG7O2l2bOb/md7i1KF0GNtNgmZgI1
stL6ulXuHRVLX+KKSqEZ2ywrmyw1LvjPinr0ro1rng/vJeu7kvyKlGx8dMME
CG2QDg9yxs2SuNwBMxnt0B79p5jnWLGEO1VJDQRcVumktD7R/Te3fG6T7JlE
VF4Ftt1OAVhZS9Al94LvELjr7i/W9Mk1NbogDpcEM1pyvmHKyYChIbkROkT9
kXf06iSMi0pMhiRqbignOwwoTiC82fzDEGp5Lx12rAn9czjfRy2WFz+7kgw6
WeGk1oNm2telZiI42eR+xklOwPDuULwQmshA0Iw2rafasxbxUDh5Lo3ep6dP
qTlhTTbiB/lQNC82kF/XOPpe3m9ZhyULNOxGWHs8MmrbZXAv19OxdxpfCS3o
yoi/bPSQN40HnC4MKgRCI5CXQ9zurCMCsLBCgvTzGQuaeSigcm+0Zn9GH1o2
UQIRWqc1fQ9zRVpciNlm74qAl37jrkq+XPsXlh4+/aEf38BgxUB78CrN00hJ
6+mMOmoK4HNCcAY7uGRieOF5hopOPzDC+dmsdgMzDCyYPBDDaeYYetBeUiNX
ZLmtq/yEg5J48+L7zxS/6X1YJ1/2c8hZJq43x8P/A/24thSWRMNlY1dWjXGv
wszB2LyOZnkJ4pqvf9xMgraeBgRIdcDhi6rPQE9V+JIfNUgbd6YMvAp/wmQ+
G2DEWqcv3cHIuLIVbT/lxtZTYJqy1owlJDcxZeBPCBEf8XjnmmpRnXb7exOp
ApYaLplutnRCxrIajXVyDC2PcYQE/QP8QmQiT4rFG2Jdj03E/lYFgdiM0ISN
W/k168ASPFoHM6wuHUcZJ+X3xyBxQUL9ovFMk+lqshxaMKy7QB8P6HYpyUpi
fPwqXnq8L2xUBMxdUDuVSrsZWUdOseVn1td80G8Lu1JQjK2OidXcdzIFpJtv
gdp3wnjByMbIMXSLQgOcT4sbKNCsyQtnYezS0Zl/HV4BvOXaAp8vj1i5FXOl
3X6VjixAhS9x92UP0cjjdUO3nmUg3mf9iK1Fhd0d0hXsnR05jWcEbvb3920u
NFLBV+zBr19rg/+GSuK7frrS+8VWEWmbk+Ms4JXGBBESC7pmGxOKE01lNte1
8ron9w9i6B9qx1oBCFP/hiD/gTMjZN0H8KOC2m82Ofjp44E4+yrsq9RVnbJr
SFU/VvbkKemU+FYnyb5nrxBoZmIxjTYShx2nIsXSfekzm8xbSh7Or7l59gfH
zLJzMcisXqyXdMYNZiQ1vfyfPh45rhtO91ZFStngLfd1zDLSY4LKnY5g7wKA
SKXSxLVijqe+J2x9LUra1QdQ9JNnGnFEa8cB7ttpVtmm3XPm6g/d/YXjB/w8
3nUO877JEOKPvp0b6qLT2qA0AZ6mDDTwKdYkYK9X7A6sSphnHQXqHuXZBmHo
1DOjp1lRHf4LSGFA2zflx7Ugh39xwZJKyWTqlHWRIClSE/qTMuGcuYqGdhm/
Vw2iAk3+ZKR1VhEl6uTtYr6UvQMWAfZsus11ueeat8bGGL3MNmX69OE1Za7X
0kxUf1KB2c6ZGNDLFs/wGAkK/PT2owUdn7PdBxHzC8xc79iQEcd6TUybKQL3
38esWj+9n2EWfmwOaaWM2uDT5Oy1jaGIvCAJgE7s3uVfZz6wmy6zIHHcTF4g
QrKMM663KmCwgliIcz8mM7a49R01Dx8plL2czVqs6a+lDZ57DVBW/lE4/TV7
Tsk6CM2VzoL8LkX2+A2/hg7uGrFQkzlhF2GZWEOTH4QGvdch1V/5Mf6cL9iz
HlanwB8h87Nf9IVJSPLJ7RmEok5MkTgquGCLeWWuhGvv9NzguRbrQwjVGsqH
ORzag7+NKRnP8JT3e3kCPbRWdQ+vCHA1XKpJwemp1dtvxuaywY2RSvmgHkUN
UyksCGL6Q8B8Klq5kX9BCuo9Yud3rWrpOxgNpIFmoAvtKQ/V8QOjSTaZ7nDq
PXGbmgBY/lvm3VCD7TwMlEWWOqfzT/oOqszPdv74zC14NrhNvHhW4NN7HvWu
DPEpRSJBZBr+hlmxQUPbi7G0CKxR3HFA5R7gmUe2RkTpDQ+Hb9I9lH6aSI2o
g1Hw4v4J3GCeF+YVX/o2cgLPhuS10lP/R7gQoNOKmchzbPPbel4Wq7vw3wk7
Xs3YA8nkA/Wdq13qv2gXEqtV9NQUrInuippWz7Kw3vIP3T68qlttUPogZVHj
5cGoUKm5ui7JX9XcdAhVZSvmaD2NhFC3HHHbhGmpSwGu3XrZI3b4diS1miqV
kFZZx21MfCy56b8cXB6kz8XMAqP2Z/X7rtwC9QMaYg3TeAocisO3t0X8o/pY
WFB1OugXuESkUlMOBnVGaC18Og4K2VfvxrOooSyiGLCGYi8c0ZFrsmHhQZ0S
9WZN1dGOktzvKHKARWqfirwyq3/7tpKACd/MRXKdaGWllqm0bo2z5PA163qN
KddOHqpNsuCU/0VydBojyn+aCZ8HiazbbJunFFsCDUKA1M7YIYl6zLo8v0aF
2Ma6LZLQCdpDppjoaTra5bCCsOG+3fq7/7PlxVcMWle3wfXRa4LkQjnNiUgX
xOo18nPLe/s5Jozt8H2VTBr1UDX6oam4q58w3CyQjgmRzAyVu16weIPZH0RE
FariDsGTcb8YGJlpHKtXEKmG1oGIldyz28AruZki5L9XByuGvmXnpYQTI8I6
Cg8lj3Ll2GqxnG35lRYpm0cEPheRGkV2e1YtW0rfJ5C7pRq55kHN6W4P8Mf7
aUHH8AThAr2pbmceaD9SEzaF0r8e/PwqoDR1qiLJqHGQKUKQDgZUtMFuhNJa
9vrfPnLyB8KmGzE6qel5PncRnXxQ8zGRoCjuOhaiaETmzzmZk3FMikWf/d5M
cUbSLXnKz+TGYenVrtE/xXH83FXi3HjtuGEAg/b/PmneckPkxZ1RWPsk/VLZ
ig8PvT1O+6+rpBUqZgLsvgQJpNjg3j2exDM7MljuoIK+ObZcIAnP2AFYNTCs
3llREJ1ea8QFY8n655T1CptVY5wupX4J91u9aSS51BlF5VI2O3eDRbHhigOX
FhMQM4ISeAPUlFnglpcBkao4u7fu/1+Phr1o6jmymcFs6folcgV7Ttogl3gV
lM567ITPOeMOv/4Pb+KjA+mS1JF4W/lEn/TDm+hiWGRnab8wMl+L4UGPWqR+
+s1wG/obTINPm5k/lF4ZqK+ipUEZ7KM3ufK1V0/rDoF/BpfutdnQgVE6zrGC
FBALvAGJJdIlMjmbCblfMRUV1ffYaKyoCFiL6LN7gx7q/Us72w5ZN2Lk+a3n
Z/2xos9HLm5xBT1WPOirDHAn93GMqzOaoIr2Yt6tqKUYZN1tl38iUHQKdpmz
CiYs8QOcwJlA4E1yg53tOr5b31hsW/ad7Z+IsGT77QhdMdiCqLU3xy0o+Bo/
Zfh5kG7skyMrvcMx10IgqdAQpSkZ8QX0jrJqyNXgnn3cc6ABuwJkjZWJjWen
8Qc1oc9qAJXbTd1flAF7iga0WdVh6Qn4ZNSDzUVwWtmhicB5LZA1gqbUnDpJ
8X2O6yEa15vM0HvjbohYcG6t1krqpizGOuTh9UCOFvN39exr2PNZ9EjD2FPp
qvtHscw8f6VghusZpVDHRKv5IjA4HYT3ebCVAfXdLmawN4a24dh+BE8x29WQ
K3QopSyR0BHePFfezU6hllSyHPP5cO78eVeuuYzRFdqOaFOCOH5hIvirycC5
ggNYTMtYfQm5c5NUbXzYNdHuf3/82SFq7Jh1lq0vR3biSnT/GIgtU0JqWVB0
MkblE64O2m3Iqw3UL89r+h9xZ1mchKp8b/TsOicABSiFZrkjJyRdJjjSQS3n
s9UYUqbXWzmjeEIsr6fuWWCPqFZIQLAxBWYbgbQDgBh6iRhMOTaPDPi2L8FQ
5YLoEXVXBmoOiO5m6smnEJr1UScgHVPJr0xz+o3/C8J4ocFcN5fpXaCPvPkf
2JtW5w5WUR/NouSeGiaBcHwNNPcnlalvRV6zD8IU3w6hw7Z0K+ClZSgrHvpq
FnPuDr3cn1L325eFJzcuVDZdpGC9jBWgXizpY7EI9ujd0wvkiVtS1m8bLjap
zOioLbcwWLZzKxmk9BG5jV96MsFgVTyg9srFSOI4ReMmNHZsTKrMf1Qns6MP
6hGykqaBub4bpsGnYX4iCh2YSB/aUmiyc7LmB1MecxQCD9wOXio/bbSU7ti+
X/0k4pzq2Hea7i9xrif7IN/o3sXF92ediper+6v+K87+CANj7LGUwVNXmiRS
AJU9KyzGkm+UPv1GNm0E5KlxMY2QV0yxZ7O/BMyCfOMLwyF759U9Votbw5BZ
ASrcyyAUSD1yqOc1sqOsCqw8gPr0setaWRyRdXo7KiDlgzsY/rtM6LZ5OGnF
isKP8WeUxv1vD4EmsW+DjgP/nYd8TTHHrTVp7BtbGj7gBiaiMCbnV+ZTDtsV
9MoSltUeLIGSq8920MvBmE/YDN/nH1uSQiTG45w25s3t6CIecW4+OzEbkQ41
RIYsecKgVyXIygvjQzyqlInQzD6wyrc5+oV3VQjQEnhCQJC+HonFc9nS0TOR
pgfEW2FJPyobOrBTSJVbdCpgik/6m/EJDE4N8nrazwrT3vBatviJhL0pWxO4
akyi4szzDy9MzZG7diGdNO3gTE+7+RlROfCOrAFdilog7h1XXc2ynljvvVOQ
VQArbetGYxp6eRU1doay4s/vGlqSb9h8D3tzywF/4PssxqXLjWcPzIYDhXVx
urd0xP/cwRlFMQRi7oEkzsg5hV8qT/KBqhfYAnc4mCHnb7tN/0JXveBev/cY
ygG2CEIlH9imsUh3bcgek4ip99seDdzwycDDyNtrpvDGh7wSbH8qakW/EoBl
4Wkvp9b5XSoWMvuEbg48sdLZokK73Aq+Bqou5GqMNsZgwEhzlTrRR9UUTl8Q
wLV3AJusgHhsKLOZrUrFNfTtMrxIFmJEUOCRLIhjbe2JVU7Tl0cJYMtNsLKO
0D+tFo3yyJsRTL3ijgrOQu3SGPpIdQnCK0dNU8pfBxe2TiXChdy+QfuKWfuw
dQouyQAkwLXlt0gyLK/hAvQJxKKuWKAKGTaGOA/CLqiN4D3Ce92fCzUwtZch
Ol3BH2/JF1ZFh/e1/upYxJfu62WjkoNLqyYhjLsVtMCVBGjdfTizCDBQSyym
2wZMxMKNvnXNenfP4UXuNv7nDSOEW8rgF84g/m1lNRbNlv7DwCfruQ1E5mEr
yyibulvf1jpvIyRmEfvTEU3mL93HO0iKkfiZRmCfGV1xyiKxUkFNjuVpjzbe
C+pXVtMMqD7Rk13BXkR+nHfF6u/82zwxoXZsxqFsxXX06fJVR/NZlczxm7Lq
4/0mWfUIm2bn0YfQ+PLNFjAz4vw9I/rEgLluiThh2qjJT6GfYXC/a8P4ntTo
Fmbk+iHT7AyFwVnY+9DEwkQllH4Oz0fbOvFhL0ulgl/izFkbhROgzZOVveIP
ktnZ/vZ9yiUivJ1RrBmhXrwo7D6v/r8qmkwXHE1bhPvsjy8oXku9RHTordkf
EGs7UW4IaN15Oq/AlendJSNEkMOfnm21r56UTTNM6h48yZ4dlF2UrjREhANl
VEG9sWUsMRIDV076kqSMRPaSLl6yM7XlUgm7tFlU3pPF/a6ShVQ7vS4GV9l2
xya9S3Kf5Tb3LUQ8ncJuO8WD12DGMjzWAM2b7JYYLKi2Lol2Rl1i0mH/T1WN
zC4BLt6xAc27vTUfw/9D05RcsAJK3JHw3TqsgBHov+x2vYl37NuKuhYGblOZ
iSsT3+laMgW3UJrwaa/Dbd8yfhFokfClKOAOl4O9F7IpjJPGdYFWtT3Ol2aN
P2PSP9l/mlMTehCUTIMigtOxU+Lsv5Bls55rAEn/p5Ywmpns4xGiQ1uTTISo
G1amnVET5oi0O62CMEGF+Q4RFwCzB3Yg4j5f1/cD86OP4Gj5ikBgTDyqZoQq
e1Jzx+9IKgup0tu+sroU0xJdNpsk2C3EjTqBa3YZFxMOWJF3p7rvlpEHjvep
AcioZs5cE1Cok4VSbCNr8LUvP7krnkjVRlsj/bXwLAaDJeaOTjZ7zIE2ZQo8
3CT3yBB4aywSzqzbbKRlx8MH08faeZtv/R0cUGL2uT+7xO/DOJQBNnnIDoDc
XYov4FSLg9aQFQ0RRNI6gWdksfP6PBvgm9odUSC4bnE1cAfvkyyFEIeVVJ0W
EDJZLyhOfwlzX/LzBIC6I+AXJI2IEAyW3FRTK0Mno4EHfRb+6UeD746xKeQk
4NsA1bqP1yNazKo0HUYHFEphEQy97z6Tu/jpCSkKIKGoAoDyeLJR3F6LwGC9
vdKGa7ahM1IYBYlbBOwSGG0xdyNHGIQ8lHrE88Wk6HP1iS3rItwN2uqlWM95
WVkEck8SgcQPqVEKRtrabbRLLg++nWzJeSDo7cPiJ44heJ0zJG3kXU0D/R2d
uTESIUJ26AVSMO7EDTEJ5LWcDlUQeQ/SxGYE5Fm805vBSjMGObYLrnFeBqA9
+nDjQRcIlIfH7hJsYAYIo4Umy5xojX17PEzswfRWIW9kR4OALH4kP5WGCIT5
1qf8wVa2Mojd7cWmsrauIOFVdU0ufDvduQZ46X1gDvibgEgx/29zjuIat6t8
J4v4v8+TleMvuOCqnmd0n/OKtR/gY3lKWvT7+vLbpUWlhAwCQvrYPv74bZNo
MLAwkhMkpMxR+oMueO/qbDHiKDzZPnj5uTi1vvhHlr1SmnTgNegltkuZfL1d
fKVwX5HLphk/5Of6rfUqHfPDGwpu+YEcdemjtkCnvx7XfGE5anknYFwj6ynf
t4JATDM2EpY3aAZF8T5afbCwm8vO9eGgCzv0auQ37SrfPcsarqggs23o2tHd
MotQLVMRdsvVJsfI1mssM9Ke3ZX3mmANRBJNI5b4YUcSlmCgJ8Jrlxir+iuN
1iITOjG3QaPyCwurJmj6+kyZnM52tKPJS9QjeSWELeLHOuFPfP+/lIxMvLMZ
58fGWHRtb1kyuJLZZyY5B+/iogRS67ZPhmzzOla+jxVZTcxmCIEdcD+E7oOQ
IBusnN1ECdSdD0IDQgO9jUxoELYUkTeTAeTz5Vvtb3se1bBLV65t4rcBbLPa
H/qx2t3XGdgXBcchs5EehyES+fk9K2kpkFHQpiqXPWy10ugTAvriXUaEn8jh
52whlsWmmfNTF3C0SIIOQqsMFu8om1XIUtmgibYaYAmjURB6Hnj7INz7pjFg
ZO8X6Wq1g9U+6aba8fDE+NbuxMMMEjS44p4u/u2qzaNWpn4PVKh6b92SesHV
fV0djZEYeeSJcbLP8rASId+aFh+gBMY7Ol2ywF0jd1f6naeOoF20BgZlC7p6
g2XUUZMxmHPat/kGuDQpgRTmQ6BvZoPTMtkaK8tCCnqveLlDMth/QdF7Sj35
g2Pmlc7L1JcXlRGoPi6gUO8TyJ6aZYGSEPzlOzVZcqU8zGHmpAn4x/3E+8YZ
sErWu9h42O2GQFlGT/vpM6TRlTaDvdsjzXB/ug3hyBSxP3TXi6/+ENbew6TN
trTaz2shKpCr27CG6M2f55vcVH76zMjFDy0E+ewFyNyENVVIy8pfw5PYy79B
eGE9CYGbr7d9QA3qjjxcIhs+ESkudZEftj3u840TXb1LW24aLXWNCOBsgR8W
wxVivNq40UZNyzoTR9GzmgYZmkGRaKgcjDtrvP7EQkHWDCHqVL2RgFHbZF5E
AlF1TJKBFITlO4OZn+EovEhyH0RlQXLtAaR5DYw37exybS6drL/HqYZBI7TM
UbaBTuQgVQu7t8ScCMlfrCw4OvPiQ1dTpNv25yCjzOmWnJCBzjemc5diD4W0
6UGtUpCRW14oDfwu847HPpCmwjlsoYqhiSfoB0wmlaVt/VA6CZdP59XjjQmV
fuEtU1Cyf8bJKJNyXejy10lNUvB+ScQtaF9sYcEj62ucGhZd9i8mBwEqgtFF
9mihkEPh7XN4FfUvVBtQYMu7W6hR9OMItOxKVwXxzwc6XfUBcCeWouewhXuj
yl/pQSlUt5UqfEptCLfMCXT6Lo55hN+NyjtYGK3ebMXYtxvlrZnawt1tyxlI
plXKDjw5B1ZhaTdAWhTcg/T9WIrLO/7P27ByqkuC1D7/MQ029co/W9x9wYgM
fL7KClM/f7GFYcM0qLfOXeAtWmohj0ObPcAZ6Wfyn9bHRoLOx0X79PQQwkd/
xnIR+v/AMELT1Sv3M8P1acZcZaVJkt0uVHGzXZGxv9kw6OejTq4RW/nI1mo3
Dkm5mBxtvxQkOe11wle9aWlimmDlAZ6QMeThJRfjbsEq6yHwrHY73yzaMwnS
PW1HCrEX4CSR0LLt28lhHyYd+hdeyIYiCocl4GNcbBRMRa9gk6dYKL7h2Lt4
ZjjdReTL8xiO5aLMigB7T+3e8V238+AYk2cSqlqcjeIqSK/YnCTg3TD0VJzT
+GuqUgqec48omg2pAHz+ty/m81Z2twzG7hNlOz0UUD3hwKI0maQOpWy7nebk
HqbUO/YoI8Of7a1vy2XH1SYq83bQDked6SeYv7UxpPDS+BZiS0k14tSGHCtl
SdvhcfMe8ptw2qHelC3tLpFioaVntOedKYIZ2eKojrrDLjBvWXUhxK12sfVV
o2n43WLv2Mj5GAvoXdjkoJYw4PJsXrzMDGv6TzUhSONxSlaIf3yU2S8T+4n1
4ujqgCh31XoEIs5L4OO7mMrjWkkv3RAETYN7KyViCvRAENzVFCnoI/1GGvhV
pJ48dVaDg4/9f0X8gHhL9yjv6l84hIq5yZrPIJiXM2D6XhcUqRW6DNqC4OxN
VLksY71hppqeNjvAVpUBF+TTpoxBOKrkVeh8YughJ0e+jHrMoYnF+6W74jrZ
YnjzqscoL1zvox4flxyCnuehARTFa9BIW5T2PZb0vgIXq7YBv/OZZ3lItjdC
T9RCmm3pOOEYNwvLLY5k0ywTm9vN2ePoejtGgdihhxdNj6cABvRgF8tBBY4W
8DM+oOTStff0aAIDjlF7Ud7Rngg120CplStJuBl8WKAEcG1DzxHiiBpEnn2G
oZzfWbOVKqo4D68igUVSx+V+3HgbBNB7FKvE+1mcWSg7uRNgPioxGtaSBSs/
0AFSKa+PjKYc6su6VpL4xqfJ3n+slQBsVWEpeyscTB/9s0AR+onwDewpxpx9
A6sPK1XLcrg8EsSznre40/g3f5nVmPenc6DtK8jaX5xfX6ckAX8TjxiXL7Lb
KOC+PMpm5PZn22gemcpM8RieXG8C4CUVCwP7KkFzHJ4fRDKeoHMmzN4+3esX
RZ4yy72c5lk+KX/wQyV9DV2CGoyJPigBgE3J/Lb43bzNXtLVt6E7RD2PEcuA
QwniXNSJAZRbN/pjBZnlsW97jO2VATP7ZyL97lKg+s8J3rceQZV6I+jvWSrE
3T3CI/BXhIcHjPfhUNBdTqFA1yKl4Zqtphj/dni17GH9HT8iFmXmyOj0rDU8
f2ZBIzi+X6RvzPejcVoxWhB/rcvT9IbG2gQau2VxpbCNPOSQ2ygWIYcnoCRZ
u1HPxam7vJsjrKiZ8m+7u59clkFqMQeYltP0x/G7OiJ2anZenAk/rL4l7fZr
Gn7rTXldMndnZIxBbeu2Ol+p5pDc8aeGQ07H+G4eUzVNIMlr4Tjoj3AyM9iZ
5F0UjWWNN9TRDwsQ7GKjWgYr8Feimbm3HB4ZkItIeW563HkO5TNl2yByFVoN
tZ5sVGLFLHyc8z3S6d5Stf6jBgoywHnQF7TmV9b8zHcBzx476oMuLcBFM38Y
5jFnT+7Na/e7Ryf6VMI43MvgVLserNaDHJl3UZ0cKaEbrOwnhZetEI1d2ZIV
1e9TZw9zV9M6O8MhP98xQUPGRrTOf9CiqF/pDDyQDoAu6VrIw8s6iDZuyLBE
bYhd8S2epB+qIqOJrldSj8yRnrVBwuzUpFpzFJJ49D5xj3IMU0ugrvwBSfrt
blZYZJdihFWv+9tXmAZoZo0JY4FgC3lKtxu+Lfo5OUFf8QwGcbdTF6rqZN0t
vrphXSj0ZK89afSF8nTc82Nv0ifLLRyg3/ZbBU38o/cmCnD3nxFjM6rHSQas
0OCSuqnGRHoewVicnDCsRM9SOvRbaaFxtfbWLCSGNKiPGIBChWlE4s0a18EQ
Ulo02YOCQmHz7O/N5b0hW5VQ+hBxopaD+syBDhOMPQLlv8IyA81WNXgMuoJX
hbKUkdxDKDHpik0MEeDy2L8gQYTqSOLil2UIG6RjtNISXo4hnfiXOjGitXGC
sAHAeRO2hoT1RlxHz9CunY8YKSlf4PUgHOn4JvvXAChLCp1UJh/TazLE0AAB
u/+oQxmnWYakBZ9PuGKWUEivSJFoYeFMsbGzxAZ1DR96dV1/okpoCspASTbW
Nv8Qu2KKdGtewjG8Qs3yMKSlCbPaXS2xI7lo9tqqgKFcbaui2WgWxPxuPrMV
O1s79Ge0vMVT54KqTzf1yrYxuHFT0J27tEAj+uN2r09n64IUyBZeYnKvZEHt
6ivha6Ji9MZAlfEBoFawAlZd/hXi33A9wZVs45TNB4eGaLbshGb3t5GI4Dxy
uMaVfqDOxTOfv4PyY29lg8E6KwCB4e7Zx4oePGLo1uZjopg45yj9rI4oZx69
NvSnAUND/9jGhv76XU3Ky7CiXll0B0AOfosdMKfyW1NJegYiDdojWZj5elFI
LhMuS5HRy7UdoAciELa2r9aDoboU5DZ706wEJO0hBK4Fv730kthhKHHmrGVB
MDDGMak7ZkXImc6B5m/+CrjnD4Eg042fB2Lu4g72F2ECutMMB4fZhXqbtLYb
wkHgZU5h15f6Nqzm+Iko4KbWlw5M9BlZqy7lq1TwsE9EWegWY4KN1jDkrRKx
KiyGpzfrBEMCMrfSffzwWeBprrA59laN/yc6VVBfR1Qx/XvhNLBujTXRv2Qm
7EZrz6V8f1vpvuij+nyqv/+S42wW8Tc2Bn89TCck1UzMx1p69SiMRGCFlRAZ
KDdI4Ci5d+leTyyEZpy1YNU1GnOXBkezbvPgn4qU2I7MOrHleYf66e+5okVU
zoE0wjBMA9GUFdiJsltI72eJo4lNtOwqChHeoqcMw2mDuJrDUC8uLc9U64uC
nLxiLu2n0Mr+ZcYgTtY1Yt3fdHtk7L+/QrKBG4u837hrH0MDYl5tkaD0lD2O
aXDAYZclJ9/OIuSdO9Vs4Jj9FQAkOlnj5oPjDE/gRtymQI7gxEJCZjfBam3W
jF481lC9WWEJZFxp58jN56CupkzwFDy/hyUWvY3Oaf+sJcqOueKCU1fjmgcw
6VM2choLvw8OPi8EhMIEFsGO3WT9d9gAw3UtL++ffL+TMyMKmHRDpxHllK7M
vOr+bm0PSHwqpWaz13KU5Qj36kk6/uggeXoTr1BeWKCpEc/Uwga6eRM/UK8m
qkbQ9p2bp3dDKoKUWG9wokOkv6EZaNQM1j9MGzrXSMNit1YZlxn1DA+sRCHM
7R6bPZGUXi22YpBk4Rhcq0k+xHVXqaiNlXwKExpfJyViT2VXcA8AzxJjjz2D
cdPIanrDdGQnsFNW3KCa9akV6hLctBJ6OKdJxoS6pXsb685nhsJeKYKyfepi
I6GYRp0sE3OZKxokSe7oHKF6JvN9BeAcJ8BktfLGdZF/PdkE8c1P7KA0M2kb
NzIKr/BGnd7JtwPE/xYfAGUUX5lGhCFGmCE/dxwpuR/T0ylkSj6tFH4FUDH9
XA3RCsReahtxDugY6mLcqytc2+DK271td2sKm3ODyX+znNLhZ8GnLsBWq8q5
4O/E0dGL6t1sOyugnEgG1vd54hRPeavO7KUzG6Hmp2cQkUwhtE7huvhjf/VL
5nvWGllCFUske3mA3TEKZjhsZ6ZLP9Ex/SnzsoEHJXEwnqDjWhcMx0At5E3i
cbG6CsJPf+Rek1YWNOUXPe/16QUJHkHoSTvifVkq52+BOyS5rVXZLBTB7QC8
aksjHU6dyMaOvziq3FCc68x9GuE2dvtl7VkZySWIZjjlkqsNIveQQKcQ8X+r
ajfiBe6szBO7zfeyESOD89PL9Ae+y4Ntyq1n/Ba3/FKxf1Ue9/+gQacgCapi
2XafHGDXzCKCzeWSukv2lDPbWwwZepOKVtx0UZNpp1nbC/g2yDLz2HzFD2hc
/X7TBHQfILpu9uqL1HN9Q+qL41D5EoHcv1IYccJR0KvFbLEQdCAOxsZ3Ao5x
FhU5PG8y+DzjzmH9YAbnFwZoG08K/G8WOljvqJq3+sjags4LVdcNam3YxHHc
DEMFujmYQ5bNaH4UAxIqmafTrOm6Nwy8XuS2CxCE60GuPO5NK0pFM7C1mZwy
cc5x2rXoJ3EXbsolyb4kFWXWtDZD8BQmYGh1WVZ4MqQ6rsPoEPj68Ev4bJlb
7dXYCDL+/o4i5o4hu8pde7JyA2xHIwOVHYuUH+maakqDjKNFQ12/GIufwQdC
kkxaXxCpjmyukvS9GV6GWPtQS9x7bzW4MuYxf778scR5Plhp1lCzpqcGpbGu
U9SeGTi9c1CKyWilQAAJN9MplzftuGpmKSXhFokepxGzU7hMly8alZRTdZfU
TIQT+xMnMefYM9W1xNzHpMTQC083/0LZriWi8ncPR9FU2MUFd9A8kd+2NW1r
hMX7XVMOm1KkJw6iJYs+jXE4iiBlhdxQ3SLyk+iiqCKY+Hnk82UGf7mmyEeX
JrU/8a5VOcd92Oxy4VD6zKuxJYHGO/0jzmk0jwF8tUokknmqF9OC2TYByGLJ
M5r5q8dqdba8D/q6pChB/IqxUSX3TfcEU+fjBGOVgPhfqosugSb+OF9BBMxm
ucst2UUACuMDuGNG3qYOh3/VB7l/OttT2SQqfo4htorpXnC0Vi296HYrXM6c
JESIIp/gFujIYWm1mHtFgIOnbibxMUVDIrB4ukMu1v6Z/SINw8lx9vnP14W6
QaS6ch31T2xLn/DZKNPvTDbNCFT9FmWrSV5cRyPky/m0kqpGFAtZZCH43T8U
Oa+L6RC1K0I8AQduAd6GG90p8Q6FLtNWx6hV1WFh0kGIeESilHbq+Ty6STea
RghFedC0SQDU1691eJOZC1/kDO6ourkt5sjF5fThYJCCGi4ELM6YNeKKArW6
CxgsE7wWA7a67ONfsx0o0eAp9csCMMZKXe3mcioH+sVEO5DLraXvjHVqMhkz
KdaQK/tWFgemBsH/QjDDKcS5W4LP1P+Dp+yqZA8q1ua9zyXcgh421/MQUzxZ
yESbgGOfeeS5fwOo42zA58ruStfnDDP+znachkR4v9G1OREi3iDy/CmpJUea
Rf3nylceETTYKY4vhOc9Sh9VeP+ISCXZZoXcuc7bjQ2F8hwqZZr14NEzE0sP
qZl0Qd5cLDcZp5c8EIZ5YXZSi5rFp+vdAsL1RgjlNVBvL0qvN2qgKRqk890P
zrpn1Co8raPgquZVWzX0DDsrCUy2soh8MkyNFjWJbkTBwpQP0N8qHGhOicnO
kw1LyHwTiNY2Vmisd9p4o80ro24W6G1kKLtUZ3AhD7UwQX8EaS7AkBIGEX5F
fsvKVxXVDH2bao9YBwfVi7Swd5jRzAe7iCHKVqHBexpFCOUFhkBAtlKfNSO4
ZTxXgovCkYaY9r7BJ7op34zu1ncWAKPdAHlm0oGONrpuv0maIhDp6cD3DdvU
mAZEnfMAHsiNDxZRPbx6iQBnDIYR1xJeApBcGaEkZi5hYVe9CMjUH6dwSB8J
TqSyc2tgQ0ns+7X56rdRvqL0PWO/hvZcIBz6oi6UxRRxxgGP9x557wtfVciz
roCqnimxLKJ5OjKalGBSYEZXkvUE/ki5BfZ76bk4asgW6liZAsGkDDOkbdRt
JWB1VMWqOsk/v1VHExsSJ6ytX1rdEqx2Y6h1eURu5peCnfTAQZMD06U+yHYt
ZnwHd0xzRrYLCnxNsb8/P7fXAqAbX2OGNOMTOfhtMfS/1Qo27lZtiBf5dX78
Xsq1k0kmt4xfjSbbNKWqFf9MEJwSgfBl7XczPB84ZY48PChcvFpfSzqCNMvm
nnyOJBzLzhA/D7LuecGskiNvpiW8i4O4lQpJoPw6oFosXqHprsR1NAXqH2tU
33uQN5GbDwzO7Fw4RXDQW/2aZfNnogKpAlFmTcncQbhgvyarnNkgZ1YQriqu
XiQiYow8UBHPAfroKyzOZrjwj7l24UOZbq5OUnL7WVpa+N60G91i0OX9BgK8
0NM7JdssD3wEvoZhANGeL1TpKw0SY51mLBtE251q6LZVB178B5sG5Ae3oB4c
JrlMcqiLKLDTpdNsxRnvQk8zjnRTyW6UCWShOm/rI8PDl3K0WsbBi0CmS2k4
4nkwUKVWfzYzJURtQ7rTnIy7I6lABnZ4Dh1gIH65DpxVaMyDJWgZ1feVYPMg
2aK4CUt2xRZX02xF33v2Ons/sWyM8XKKq4k8wBYKvBgMNsX3i7mH05FppwTO
G7a30Xg/piVBqMndrSSWNKRuNNpr1v4mzmnBeJXyH4vTQB86x83UYeBIM4JP
dt8/6x1bjM/GLyPaGzlWCieVFFVl0Hu0SYPVgEBSDkyBQj7vSyJ9HWx+Ihew
+RSe6vKC4jAm3kLNVwQwLzdw9roX6XFEVewwT14dQT3Li7ieQXeduuyXJJrH
MjG6u4OJ67SuGTDZefyfJHIg7+6+TJv/gEyMMPRMjapvmg49K+JgVadjiWuM
qC2Bjy8NdUKWYKY86JIWY1GVTonI+AXSj+zQtxdVRZTk5Cj9pMeRN4UucfNH
uQX/UKJVfe53EiBXvDDfqCo2cZMQxBIeMiHqpYPQeHcosEOumY16lf9ExEMN
en788dub5S1wRIgWr/YVU9mlzKr6LLrI+F3rJZZbo2QtcDkKgXI6/AWjcejS
0imIXaqRUNgWBHZCCwOl1mdDvfLJwQzA3OtdjYwa+8XWmsxZ1zWVAYsQU4ni
OVzrFPdMGtOU4UGhTRx9a+5JlWHTikxcOSS34h4EnT7xcbs3FmeKONwZbaRK
vUu9qn+INaMea7BH5T7xp8FmJ8c3OtEBjSg3g+/Ogafxj8i3vHToZ0JyS07A
W+mEqGjyP5mOvhqTLiRcLstdJZyGAr7u998KKvdvUtTmJ+GmLPkTFHSS59xJ
S3eovT2qs1+0g8RUqs9Z4LNZ/+pen7LptlUnmvFRqPFwjXerGvHdMrTYM4fq
1bIs9J6pc36ojFGE5Ayh5D1Xoh+W3nLvqJgneaxu2ww3oP8hfRN8r165Aem1
zPpUh+7WME/MNjeuwiev6UH8Th3DznMZHZV0XhftsI3qEN+KQtRPdOhaH9YH
n5/lAR+lekG827U3YxMbBEZKCs2OtM4oYt1NRxtB2WqGD1f09+mAsPK2eGAy
JXxIE1p2vsMUq70+KjORRcOnOz0aWTts8nsI58MKMiTnWMcmERO7l3OAkk0A
vPZBRF8Bi+pr1SjF6btRv/EhP7YjlYYhGPOQXxcZ4OUSNnnwHdIF74iv3Iwh
c9fJbLUcucwsAMvJ7ea0yB0qHG8hvP3aBvih6/KJDsiPuCjViM+mOurwdKNk
WOVKo0UVACokVgCj4q6KSHh6gEaOqf3rRIBBFsUbYMW20CFWzN6FcVqDSPjp
RTzLIS4LRByXEDqo0bZQQxb57xqAwW9wMPBKgh5m4zkgH3hChhEhtv72ICYg
uyxamDwPs5xfc5kPWn/1dqyAzo34FaYt/uwrHLUKx4LPNJqLF6I5TvEYK0gZ
+F6ENbEOvx+x9TZ9knrTRmgdTj+SkdxFh73512RAZDFiwwo2okpT6+uM5Ksr
bpY6GbSpD6hRVHtd1uxk8Lecl5YzOAfYPZ5YVsD53yF0elzoc5WSLK0pCr9V
h4CLLPEhF22/mdQJbNGfwKkGHD2opwETArY7X6sAwSNV+G2+mPvMwZb10OtA
Ldcwfb+afBs9v9pPXrhMa3xAlV14J/pW2AzPWzNF76MhKVsnrLtBvkXR3eCM
qRXAzGecOV2JbafVZyroWsaDBzRM/7TbNkGcEcSblJvBRxWMeHKTRtiYYpGJ
JqkNV095LuMx4rZ6612sRSVCj5DI+onYHHoLap1NctxMW5JVct1GDi5a6J1m
Wn3wJRyL0N/qMtCgwRq/45dozxMZYU1XYDnRv5mhgJORu5V7rNBqGWoA8quP
YrWUiLc5vw+juV2NnheKfIRsqsUEOXQxVnzNHM07NrXTn8e2wI11eCIHmUIW
2+TMdyJS6CNEWKswBfEQZOCfs9J7pKRJkI7/v7YnDXwXu6LohsoS4asYgorl
aPTU0jmwKEvt7jd3fvJjL2MEMJj+PE16m8vaZDuN4iQYPMOsDzZOqrpccw1S
ng2NQFa/XPSwspoOXnKLgLltYzXA3vW8wXS021+BFiCIZsHnihuEYhFneTmr
WVjwL8CxO1yBMtJgHG6hFiizUqyPVod94UvuO5wQHt7oK6xl4yrdpn1CZDCt
ccqWOsjrJcAv+Ht5AIxZN7r6BrLk3iglifx+Z1anTUVZz2zpnKn7eN8DGQaU
vcbnUiDPTmwVmn/Vm0r8qJbCVECIsHBrqpduIYJUdkEDdUxNUJ/2Zmx5qARk
p5cjIqx4g837K36gHhoHhS54aeXXP97PJhLylS6nKhB8c28VN4pWteayElxa
jU/+GKJ15fcMLi7G7vq3mTi9r2KpGsTVyuWSV1CRmGGHigo82DGG1S8YNfv1
24m0h5dlU/gUdUQsj/52e8UfHj4+YVrWzCW2s36w1DWzNTDExHJPiU7HRUhG
Qa30QQrirkrkjm2/mJ32wE0N2WivDr0f5wtV/5SXiep5zMOLerZRNF6YiKqT
DU63FH2QH8vPE60t3VHJb7+u1Ze4dnVe0QoTdryjvKbSd2REfG9WYv0yYoLq
2pVhcyhRtUMUNnwVLX6SJveEK2kUjBUyOMVDG52WyjMcZOj01+Bg9vfmbbzu
0ASTr2292XJgzztiSqNL3kppRMFPdmbn89jY93z4LUX7K9r/ImkMCTjp0Etg
X+S+QSfhyBqTmXe/YGDNDFtEVbiqPDZet2hfJ9lXgQm/M1tLh0Op6gDoeJJa
xwC67wBGRFXML5Pv8SXJCVc9XaXo+l/l//l/UoHI4L0aVUQNsRR+wNV+qNwp
Sk6r/mM9gyvEayZr0CJL3894i3xzN6YZPp6iC0f/+LMeFt97IoBDsZ0a9c4V
AyCgQEBuEM7kgp3Bp3v8S1/YmbLh3ZiaLwSXunPalKDoaUANyWQettrtL+nJ
z2F0+Ube7oKu/G+IF4Ji47vBPGiaI+JXuFXEManf3sJYr1ChGap8sW7rNQuq
O1Mm8TcgPRfofZr9qssM1+UyT8gV+FWwsbk5KlXMsOQlw7JEZOl6UYxOy6qE
3IQ8YfkUOUXI+P+yyE71hDCZG4u5RuUA0ayc6zBueZno6leKQauYE/jXXKyH
X5i/zhxjuuLujkHXU1tihRK5InClIrV/JJyiHURWWn7X2y+yWun2Kwo14O5A
PDs8hRD5dTJVz3FI4Lax7kGFAicRZ3bj0PNyhp/zpiyC2ruHKdF/4+Nsu97X
kz67Vn2nGvAkPWIy5dHrVgreFwM4DwYtw1VD6KXmx9pdX1I0RHhJwUCVbAsF
lCu9yT87813uMszS3h7xDoMXyNnwLzbCkJoPSlH93sJCIbhkYSfGb0AALItC
S4SMTM9cDVITpqNrgJFwUtpUU0lN8a25hYzB9amdtUo6PEbDYpSjomDRro+e
wFQUv2RGBArohU/QYiHY8XG9cn8sQl84dVYNkwhzEz/vsfc5V0bcXkrFbno0
dln3raihd2nOpwvkhXxlJKZlyRLqJ53xu9H5QRmga3PQxRtTpRXYkNZgV2VL
5wjdoiFdQo7nyq37z+gB0sfggwA/QEhM6GKMFt8MfNaGyqCR3E83b7Ul84Fg
+vd7wY4WN95farhQeZ8w8P9VykhQE/dAtcou3QOoMRMmTvzybblPZ3uBxf3o
mNf/RK6h9exViL7xKYmyT83n+Up/STwPOJTm7RLMO8cJkGQAjtweplbWguzH
ikGoTn72SYbmqf2apIeG/ERLuo1XSnALdaUajJC3zMUgvQQPOtfVtR6xpn+B
fWIXQfZ7fSRpm4c/b28PUvsDl5dz+oTrl5PODlea26jbN2MMUqeb0VxcffIs
tTCD6R0gRhUpjFKBczMDEl3TUweFDFzEbazIAVE3CyFzTUS9ffUzv4pE2/Ex
Y/7gqV/L4E2z6dt2EMVGNHoLfDZf88kJKV0vW5netWCxxYhZmvDx+C280ssf
yUubR2iDFhqAPn0n4CZpVv60aqXo445S1hDdKyO9KSBKbThUn5vCFLkdCT7i
SZqXmxTsIQFCnI3ii3Ic7A+4Em4Uvjs3jlNKiN3nLwHjxCYEAByYA+/n/dOj
1N++j0IvrGmRK6qbeyPVmTJJOTkqTfPLOSDIJCXNFiHJsHR1u8sUbCRvA3DP
1PSX6WaF7jbv4S1emxjD9o/KHn9STieLy3XVsCVW6Rtden62Gu3QjbzB6on7
lYVqC1+qbKi6C0y+Fvb3KZFCkP9+ag1CDS0zUmSczTJNVwgrqKtiFdAcTmNh
kiSd9DkjFfiayRoNb1kEilpuC8I6kP1SDnQGbgvE2vO8NUZEJXYhpxX8VGZJ
5bpdBi+x76YeTaqsT52+SeB7h9PwzO9ABS1hxmBnKg8aW/OoeWC0VdfuPj21
phmDXYfUpnZ1Eny9p7I5pwL1XB+alEyKL2vwaI7f7eChPqBbzmWTjakERfgc
P80HP5IRSAmZ+uQ6amdme2VZayfhGPeOpi5ZcF6R6f0738XQXE/BkZ3eZsJ/
uB0UlPNt+NJpxIt0b5MeXBLJS8vcMX36MPSsTm6hamo+8E+e4uelVCd+xjsC
WZPDtLi3ixfnbd9fXLIGNNSAOoivwr1dWUMpYT30hvAR5+nBfHFgRigoMEe2
zTx6XCHOsQplqnw7IfUYSGGUI7HugplVPoLDKo7DaJ9qkqrn7Pk+rTyNvYAD
+haSlDQAU9j2/pdztXNrvpHeoNNi4NU9RLkD1kegpeYMSORjv7KMGthyYnMa
c7tw35y8BFoDxY54r/eqKH3D4xO19QYK5HTXL/RepvOGACv8ZZdS2Zmt1/nW
9B0gkvyoZIbnXOwNy2eupJyxf9ylRz3hQVzMYE3YVaNbHxtYBcW/VE5pXtk3
yk43dB4ktvqTJaxawMzuixB63+1g8X+AyOTWp+ehyPAYpQnAs1F1XqYHjN/S
047PWHXUX3g88gjJHymES7WL1krZJFZAUKEKvtA4xpUz2N+D0Oio8GwDCRfB
LLQNoFSCvA6Ampx8JRwMOPDbNgjQDw2wORAVOGxAn1ctnTbh4he+BQU3n1je
YiKtS0bEUfI9WBc7oGObwbCVo+m0irH+lPFW+74w4eJn4sXcQxBXdkZNgEA1
0XDNVf3fsaOAd6aQDbi8i2FGG88qyajdOb90D9T6yU9hL4HadC3cJu9lpRfR
9izNqEyb/JoFZcJSH0bt/Zn987d9tT7PMGxRDM+JXwtMuVBg64558j5if6wj
L/YcJXtVQfuuVpQkZRiFnNogHp1q3/akCOsQpnjRlvXJhx7jMKS1bpasNyJ9
/Zf5zXYsUzFA0Kk7HTz0QfUjLyhoGYnJKsjrIpjOL0riilTmjVURaV/F60Ty
5/2tgnPNjN5XBpqUspOXOC1ZRSFVbb5ugpoA7/T6mRs8RB0oYkEzRPXD2RjX
hQ3Fu6sMpEI6wnYFYnP8fiRy3B7MIOc6t/PXR4d6yaFsCiR+SVxUE4zjApgp
FhrON5SzcMeD5XaEPpB1vrRlstO36u7xv5otcUjFDTGcrZcvsPlpW2PI5Xn6
wYj+d0cw8VPx2xjTZjueriS6QK503Ro1qm9YmZGMRHFZdh0XKCVHVg3S1mYx
KrjjdTsZhGnzpfv/KLxoPrYp4MMPJaEhi1hKPBECOyqBxKwU7q53lEjkVosR
LMJrn/UFG1y6GOmS6G2Ns5rQQVafmIdVy38FGwf4cwEsEBRXnYyjoda7VSLq
hvreOO9zXe8AlzD7uHMnVkgS1PCaI9tK6zhVG7M/5q7eEhSt4CxjH88N4U9/
XtdkmnQOaayxg5DUNGVBz643NXFSDSMX9SzJMtJoitAvahIaOsNiKHd1xMhL
pFFB6jYLVXy8UQC7Qm2uj/PsSjT8+vJII+nxLidLuMBeJJiLIYwXWk2iyy58
OG49Sh/7q6C6aq82wmi5p2TS5Ubt36LISbpGS5k34ebhfxhQQQ/S21/W7iWv
buCHKZeniIHrUqZvUs2sXKm0mxbBq84zt/WJkin0b4mBR6USTCWNauJ0M8PO
4ZNtOZgUuKT3Sp5s10QXprnI5K0v1594mq3nCR6aV68RASokHOs1LUeuF9Uv
b1zfvzZM6TwD/QFgAaSRDSZuULF5xjTAD3hakUCoJ6CATWeaekCZzaq7mNL0
ZrgELXL4Ijiu7NIJPAtyoUIIgiUQD4ce3xRr+Te4YB/iYSwr/dAIIsiHqZpZ
puJu4P8E0k2hJkFefqHCWaY6onEP5c6EiWghmgRpSNTUdPGdXz5Xln67L0P/
MEtQCmJ+skq6cQip7lX31FShzCrV4X46XTL1xD0EVl877tgDIy6WRapSLmio
+PYzJLdWZs6dTjWceLUOrEzd7NlF4ipl7a74KN2OYwaaAfuSwxZlBXkm8MRE
t6XcveenYX11KFDXWQJUoDBVb3SinZxwInTI1Y7LaXLSnLhpFghjkCMtdjCm
/aos5QVtqaPfjriQMvBklpamb3ISpY7T2zmrEkk0CoelFoBoH1h/Qfuxs0Op
jYAaBL8XG+b3cJmX2hUkf/PdXcR5XIoPK6z0r6N/zjE4UN8VlhDS3mV9vrf6
v1UEqarjsdyC6QQp6KlzIB9je2fjVn4/AmEiAr+rzcGKZc9ZNdMIa5gOc0nD
VwRE6XV48Yukck++m8OXaiGE9VdWVVdcJ2jjW9IdcRD6/zVXLzx1ta6PNXBe
KrdqqzRX+4Vee9DEwKd5PL5zifZLEBhG0MBn127WGKIalFD6EISVOql8qcov
IPPH9bxBRo+5CUz8osi63nNCcues2wkXNVAutO12scAa/1RtiJFoxmH0XohH
EBdBbV01yxeuAcCZ8gSvFWdyvdJXC2dzGPfbHsoz1YLp5CRHsjpZ18OvT2s6
8n33g6rP6Li7LPkOJmzipSQwnThMOLbEzurx3kdZMer5Y2+XUakefuROXypa
dG79pgUuvGt9TQDDH3gIj5zppj1SVQg7L6GxDnWmXYeykkLjEHk8dP+bluei
MMnMIdY32ylD4IM15F51IqdzIl0kjIUOMr1acBuKoKkhljfgJ/i5gr1wy6DB
VgE5zMj5i/tgKY0n3Svx6bN7dKWI9nJgEwEAukjkG96blLLtYD9OUtaic7F0
zi4Nas1h8MJCJQCKhOGOQ1RUmyxSmz4nk3Zu5/SkUlUXmeqLSCA8JAFq9gto
E7IJ7Id0TWb69MCp8fiCUlK/ZhOjLLLYTmskfKkiIs0xoR7v6oZKFuHKn5v1
gKsDiOe0F8LtogtL6fBcn0gLIBNmKfS7IuZs9PnYYtmZvhWbsSVoUyQbOI+l
cGtvdkp0UAcYYCgTYCR032P8FWYdwqqKXmTU62mBYUHDNMBLz5/FfO2WVIpV
M859WPLDW/+9ENYMUS8FQT2Fr4TJ1lUKvWMsBIcuVzhlc62XwVql5+yed+Ca
1nC+2HUM+eeblpwO9y3OsyITHusuj7c6hQl2qnDp5Mmt3VOnRN3TiQBq/j7D
+gKGr+wpF1WosdRBY8KzvaYJ7miM/CMHIA3aEZb2kjPkHdsYUSAeA0Pkb9mw
okoo9ac2vKBpEPw7RzohFrg16kfAEt1/E3kQiq9RAE4+6vDQ1pC2oDeNgyfA
33z6CRzCoy+1gHmoQ5jy/AOO2nlNeGAjnqFlMsUfOJNNUunPFgNOpRPwpGgt
3LyZ3Z3t1Huaw8MRKXZvu2PLgvn2+jpH4IfQ4MqRyDIrgtyPdPD12peWnAZT
Uy6Gd4KWoQ/K3eBx8HnwX3yem+3tC3IaAsS3K0faZEBFQEwh59n92mqw3aTc
ZMC5LUhl6qTlc5xhnL8e6CuFCnNBChG8FCgekbJ8CN3b45/4fLw1HET31aYW
7CEC8WA9HPtN3PJ7oTwSuuJFScTOazvjC+EtDFpJzqrUg2e9Yjj6zCpqF6I3
bpmh7H90+4E635tfr7tMpM/MGdKH40sLtVHjFpi/aOHbQT/2wUadvPTMaH8b
XsNsz/1QG0kaC8kSzqEEjyPpTa7UZQBNl3cv/FZiQh+/wY2KDFQd0lajMrxd
s7sPKnt2N06LS27EUCM8W7pAQZLP08bmdEyVWJGBejP4913W0u3ScT2oi6LL
ciJe8oo4ATP/SHCEmoJLubxPwXRSKyRSUT9RaeY+n474eWEVte6CmG9LhjM7
nZsIkGk3vr4+fldQsnW7UdEKXhOwdBwJlwLE6cZ8dKrjprLRYVwgwl+xSRsu
BiST91keHk3S2wDjUzeJnJ6Xv05P7FTndeIsR2apq20BEdpTgCtfLr0CxmgF
8caoUuv5crtvxBYNFmhXJQiIUY4gUT4sPTBtL/BfRFkncjWslUqPmXJ5xPgn
f8SMErMTGIt0Bz0xgQUi+8lwl04aIp1OwSkqFFtG3oP8n9dcJsMno7/rhcja
RMRTIUrH+a3fj7T6F0K3Nhch7vs3zZ5not3vakft5jC/EUk7eZYPHJ4o9+y4
S0EHDpBY5F18HLFlauLGv7fxkAgVXwvpczBzpVyO7gP7r86vcXetW/cVlkHi
f5pwOHM2E0Cu4OPW3TfSjah/RcgIY6MZePd8KkfOq2rgAsq0aPTH8lbIWmTp
rOEJsVZznGQBQYDzJY3CSfxvkv1uDEHhrWAE+zwRiVTxMPbrZbr8HT2jZwgE
Ct7qzIBPKgfTHE+b1JTnrVPuayx+TjjN25HLQ33SFiGUPEXLyeW0tKZ+EBR4
H32v/xlUfw9fDzStsFltLzkRA0/hqBfUVKaUgagG2xJcgd7c8n7ivS7bP4JX
JBKXIf3M27SHVgYB8XgVbNpYiihZF/XMhApDw3Lo9bn5GJIrzInN7Ib705xG
4+3WJZgOoSWkDF8NaIVgnfsp7puX4LX31OG93YPMgh2ZKy1AXhcMi1PdSyr9
fcjY/1gttIHiVF8akPssyX5KLBoN7FWWEzfvQPYwVYkYr8A8XaZkbhrge7dS
Qn+WhlpIgcAdN27dBl1IE6Ujxua4iksWUs3G0k0LceQnCEoprVQnGHqgAjRd
90pgZ5jrcipm17sVdUYvRVKka5j5qxAFhW8K9gSG1PxQcwSgiSfIlV022Fqp
/CZq8ODTczds2cQtyy0Ym9er+ljAW0/739H6/mwFtPKnQCrbAB1RSkmApd0t
GKoqAaX/wofAnabEbsrrto48X8mh1gRWuCJHZ9aU9SrBBfwnugZZECFMOi0g
R18Eec4euXjpI9aVa/5PtYmFS95I5vl9SMQ3WU3n2tcYOLhOybVzjmhXRcTx
ZFwP8aSu3gBM88cbjLzoiDo13SAg+TG2f1KYsYgmzneYSJTHzdt6FpiKL02E
Y/EAib4HZxGv9tzJy8/UeLbr2hydeLd5ly29uElaCT21T4zCCgWYriT1Yhdy
dflglPoLaYt3VbOpBQ7jeSoUElUYOzvqRvLxisJTFs1r+AW6WroPHZXnZy0h
VuTCEaL5jfeTmh79okhdROmDA8T/p8GhOe7LEhnu7gg5sK3/N0I9v1Em7nrR
hJkwSvfXL2puHamwNpi9bCVO0pVtxHozMZHwc1DT7gp8He7wUT0MILv0Yk47
ptmVYTwBNHpMs4exD+g9I1pSQcJDctlOYExPsD/bMadA83tYX6h1Nwx9fk5F
bsIoiMjK7c4cBE+ckKAIc7Hrsa3XNFL5SPXtap7V+UbK1UGLPLH0GDoYMK5t
Hb/Lza5e3rbtFMAef+ajrReRPhiW9UsDXcUVWjG+qb8YvPn11zL6Q2ahMMLW
j0+yDrkJfSbyRWjwFSVKrIUI/8ln+IyEhZllZ8VXW+MaX/MRsm/cC98yPtkM
Qgnb5GLQI9/Mpx16O8G9qn7OxLpWmgYRWlUjbSCZyfrs4YzWWd80PI4KuPz1
kG6V5V9BSmzZhLSkvycm0ZzLwsXNaTP660AOUxh6OUw3lPMdKh9Zh/xz/fq9
deRBxTJmQXLC22mdLZvBDBs1FuoQF0nZepld+xzfyFIj+T/LJSKGr3ccuB0q
5jVjoOmxmkOE4gyB9xWgDkzIxYIz7WNtY/BObhgqvembmdFdLYHOEDYqU4RI
cDK85n5c/S4PJIJimBlF57vqWfZffPK37Z/pKACVfsZylz1cAsJGDRASVT8h
Nb4bcLHTOmINTDC3WvTocORuHrAdo/CcDtp1m1tVR6wQWwa1NvLgT+W+sDpy
Smj+V25FRuZBs6WvBrVHyzQzS7O4r7+r0ihNBQTNOHDBp0a+J9HcxeFDBjJy
dOFhTAtqzhbu9lqpXc81AD6LB+CEtOdzC7lfz5U7kOS6cG8CQ/+mbJXEO5z0
ci57Ix+zgFo6d4vx/bMzP3J/EugHAfxs6D7Feekv4NVimk09CsKdjZm88k7h
2uiAzMICxW5QQ5FfrtqtKzJfnYpAl4tBw9IPOC3G6WI2bvm9uzH/Wjhdn/CW
f338MmrEn5qUgBmO7aCGgxvkdTP+lPCKpzv0zEEL5IkkEAML7YqJN5stXfwg
uUKfBRSkzoFKuIUv6FFJ62/ecA6ciladTfwrbKoXL+u/hFLUPkcG53n2DG6O
USpvfcBnQX8LtqOfcZItSCc+d0+/OsodWlISrzHXSUT4HrMUYNrvdrHOIGbn
RnksV3i19KzGZrjdTLW4GQk/MFcLKr3bEa9xeDTh1dP0ghf9R0UTbKn71Kge
lPeObeIW3qKkWPleERCmO2yY5VlRJlG8B2rhq12/D4sunjJp+2oMymuEe/FS
2ok2QpWp8+PrwzjeYrtFlXIwTQlPBiMVBSTnKm7uZSG+DMgXsWEhBooIZAfE
bJrjfI9daCk9Hhy9ksVXmgn0Fp0HfVBk+pJKIhZ2HKdyoujTO41Q1IFn8ggk
ESsSSJh9rEAwP9cgUw7btBHrp4WZAZ6yS6g4w4TK16U2JhQj7CZq18KUjhB9
dMbY+icwqXGlNbOoOOJ1Guyleube3hE5pnNxfOJ5OeuAP21TBvPsv2XZO2Tt
eYxUmHJV3hxUZSfYc2IZu+oGY1ZWce0DwTWmrKZcOLPL9B3+UUbCZ/BXIEyQ
ZTWPvNExc9dU9br0qleqVrzZj90NhO/KPmAddoXEAab0MtHUPrvPc+DL3oFl
aImvS0Yv6J20TgcCSWQKqXl60OD3PJo1Xv9G/t+QheLUzP0LQXbCbGqsYz8n
LoJeHlZM3DO0aiTt1CzrregiMq1F5Rfbu0H+DdRy+MZAuRmdXaV9bu1Q+hlU
0agUrDoidfvbCp7jJQh17p3nwwTsaHaGx2bFLw3EBFRD977uUf5Do6RkZkOw
blwqGd9V/f7MTGWz5TlFi8DA0gYYDMOr40JlP7jUEvHxJlDFvzVl9nLsJh1p
h5XVqX/MmuUMJ5L3Ljcy6z2/T99iu98TDvX0aMkLD9BlkZ3O655OJycAEbk8
vdXSnnBkOLT+pqxNLHQ7FFmdGyL4CAezEAgEvNLXcLzKM26Oz3IdEm+BFPHX
koHcl6HSNBm9eBYcBMdMVGm/CA9VmU0+v7bnS7qjne/lmKHBKjNzyAN01fgG
NCGdozqV+AVa677+V8nPzMSUZeUlTEwphdEZFG1jjbC2zi/lWZD5CNrHXF3x
fdem3pdljLaEEVFwN4owj5ksMhcX+3BK6qJn+3YRrmZGGW0RMV2CBTyNHbQK
i8pTf3D0EVsy7aaz12SOqw4QHSKzebkZsMhe0Jbj4a2Ktxqor1eipmjP8bI/
QS6YLu1STGC4dm7mCjXmDGC0WCbfGzWt/r5txkW1Z/Sy/BZycnuHDWtYpxvQ
sAVPPjDIFCiswO5LfGIGJuiQQHIFUcwzYHFTZaDel7NjnprqiAQahmOLV3Dm
R5wa0wXQAXCjp7Nd8zBmF40BJlbYnGR29CSbqUpqaicbLM07pbf1b5h1eHrO
TkydY8aVgc3oIIcx+N6bXjvC9rus/at2T/nhWd2ntBI25UQZKUJ+owUW+dVQ
TU9wevoBuOKuzU56STgzoeJYlvEv+PeatW89UX8tRkV03Wa3Djcd444zTl7I
liH+3eLZsvc4s9/8bLSjHHNqnvs3se2PL9/KNoZrlUrXRwIlUizfndfVp6uK
o5PsEM6h+zfJuRCU+ePwiQy9Yalq/cPX0EJj6a9sVn2XoflIqRS96575y9X/
cFbMgWImFP4H73jMky0xeqi8ZO2AQM3b/+A5J035DetX1GNr0M7XhBa87Snl
jJYLbAZa6nUJUxW/3E4J3KCVgoBNx4A0pHyDxq1rt/bQwVI1DBETnN50oRms
X9yYFeaU/ff6wBnlC11RyGRPotNMXn4W4KJXQ7/D3w5F+cuLS3Sz0hjnO+Sa
s11vPW8VmRg9tNDna9GD8MbbGA825x2xgcPY/wvZh35II55HK9EBPpu/hmnh
pNfstxYzheUvK8BhpNgZ5jTEfLp9xXxtd3NnRo+So4vHMCoQP1EElIcHkBv2
yNLDmSk/rBsNmgSdi1S2QOZHxruOVe71tjhmMUZZ+o7jaDCMHvrXoj69eeEl
awPLCtpMFqg08I8ZvXQnfQbLYJEObogHTipSMFqUV9GYe8Mk1AOIfFRy6dcJ
RNrJ/FgAmNQP9od4uc8GO4/pKNMCLEA0B6KmfAfNBzVqA6F546qwnKO9EDOi
n0LXIHf72a2BMi6M5OJ719medH6/AxgQVMUpWkA5ZqV/4MIZaKCv6Kbm3V6+
g9eSPCGIgigHtbdOLpFWHpe3XUS1CFkZUrdu8ymZOn0lkVYzkqBz9a26vSvt
Hau4t/n+SdKStbW7FQGtlJBqXVCFcDyFA3FrBKjbzyJgRULqV+RGjp8yzVh/
gyy6uPq/46VtiidH8Vv+S7dwQTt8Zjnj3OamQu4Clov4grEA/KGqi4Rozntl
IyTp+Sdxxuf5atwZioIeKEkpFX5pLV+LV2ZkDBIsoFjD77s7O17pNg/lHRMH
gUGJ4qki1pnkqT/LVbItS0JxrSw3oDooKyPYCdHDlBUK1+hJNkvrcHC90nG7
nUoTXZT57TukYg45Sqk6wL45c9s70XbArjmQSOA8XEbcLfM9aEnrMSH/IUaE
GhFBCeIuKnCQAvM+MF+P/La0Bew7pvCvn8BWETXNYdjoerKAVM8D1dj8uLj+
y4rNydJ1HIewDJhoC2xKxD8mrjGqHFw+oEmmrfplJdlfChBBZtNc2lMWimYk
8vlLoqFAGpNGWNBVVKnzoLe6nM222is3X3dV7koS7zeEvMAOo21/LnLd7SeM
xCOnxHAD83wdGFmXz9dx6qy/AXzSMr1IfhkpR12JjeMbKZWP/ZAsY3Y0iLyi
eNpZ1p8lvIQAmoNjsIDDEI3h6vgGekH7Gd9oALcwE3zjgHATM/4j9Vr07ZoD
Dl+tEvGSSHfDqD0T1DPxSucKCsXN9pScqoswkm1d466zBqmBpR+oWib+Upfi
iYGN2u5pdY8jTECE4WUDM0NS3UlNNqT/anpHn/nWpib64Z4VIk6eGZKRgmtn
OKxkFXdIwnl2ziHlaP+5HC8vwldA5AvfkEAc2S3DB0YWUhH9m4v7YHzBxHKC
IKhxKN5veTEuaUUfhB59RG/xhN2P78OPCC/1BhUhhjFpNQ+nkK0cxzU74YE+
UR8pN0i4sJlo6Oo5AztpVTCAooZ2dLAygnNVOyHnL0A/VkbnHGTMo89mRku3
HGvjklzaiM34ds/NutpPIM4A9m+YOYIbqsA2yLIUuR+ABSf0cQnr6Js5aa3V
JDyV1SXHUyBZUC0oY6yVJOTN1A6qB3gZwrgIF0Q9YBS9TpM3uQREFNHvefHc
86lk2vswV/izqoFCF84DB/jR/RFuu9cmy0sUtW92zDRd1vseKl8SPyk96DFs
JDKoSRh0639HMQ39XJeMbzj7hw0PnB5go42OUoua2NLdygUbevxA+TYonJRF
RNJ4RBHgrkHAZIgP5wEisRtSitPE3vmTDSUr+B1zb4BC1n101pueHJn9/Dyf
Mr6KZIBAcGYx9EC8PmiL7wcHuL4LLcERQ6jSxlEGgZokC0cIfjheJoC45FgH
fkYI8dqa/TLroaybxr+jFgEcHiZDhQlXE1AeX/dRZF4qRmv6zpo84JOE2V8m
Q3ARgh4d5OzTsIpWcDvacg5o83JbLcPrw25RvTH9pjfDuChmc8Zr01trhjk5
L5g3VoAfee84iYVCS9csgOcSEh7O4C7mpq0hq3T6KsEMayGkhAvwc/gQf+ww
Eb5dNFJmd7Aijkay7i5GnSpXJu72e+ehM1hoYDmMvSvcR7qE2l2PbAl1i4ZI
ajoNhj1GyeB3F/jJHw7euIBrmBqP+2+Oaar/Lvotyn9MYTnI1MKkFAQJzT78
0RYXDikZXG2x9yGYMJf1V3k48ETSJ43Cup/2xnlATE8bEaqtjPdjK/f9cgMI
3y6ZZmS4Dk0RCV+oXWqWFkn7MKfTngYq1mN8UggELMpX5G33Cd3t9efqcAta
lE/x46SofNYkUl8hfAYVRkFu7zjpRkpACQW5vTmVnrlDAxBjCgp+6tzYqYrq
VkARNOrS0GyijSVDwUxWAHzTQtfRX2jVAP5FX5wei56k7SjZkN2eGt3qqNO2
4B+RXPW5qjIFh9iBgB6l48A3Dz1bU9zI0IvAmUL/uYNTQI0X0YQBjUwrhRec
RwMBZ3yK0rH/UVK3ysMo2Lk0SICRqFKZw13H9tf5Kpt920el0N5CPMr0UWWO
SQOCgcpgC4qjHfIoBqdqdmNC3D7iL32opv6njBr9Oadr6MUtEI9IVGMLvBx2
HxhZAyckdfzg97YTszs/SK/xVDGEBklvaGmSjiyW32bSHnU+IzdtF75xU57V
pSdX9FgLHO/ua3q4ErGFidHc8eG/TLpUz5bOzF7FzwldFTQRjlz7bwOPIo3L
AuUAFrS5xR/LdwFkFa+AcYcevqY4ToZL9I6dbDGMWRsHh2zOEkQ6O3gRZEeX
VQSK1+tTG1JimRUPoVjqpJVJ3J0Bu0DmfN30RXnlNb6+QoOOMd3QqTipN6YF
A1UgBdnMbTetptdtQg3A3wsCcVwQ7Vk0eHQW+lNt+BK8PKYMmmYhwlZto40H
HMKEp0lKEx1qg78hHsOsYFCtEdjoeIFJYBHWZy6KPi5v+Xh6KsL6jS6YPQk+
5l3ogpbxnMFyPe6bZWGsoKPcwNUoPl/+EJ3IQ8ebhTXtqQQEP4tztCaNAZGG
JcGf0cxWwRpBcy6Dpjc5+e7yUHhzo4uTKwRd1l22IRiXjMWnwjzC91U+XkdJ
yEuKi7tzI9PbXh6EkAgKNtNFTsKnQPEwccWZCLQf88ePDcv6dJLDuubj3w8o
rsjWH0yW1lUMPHX2UID+F+eF/68KoL3SakGBpx7Y3J38tLxoLDb+tgaqH73D
o1FzCNknfe22ETIz/5VPhH2N/k4hHaYT0PtlBYkysAFt6yE3oABggV8gTtQh
7kGsX2wrYzdxVK1yTSbUvbw0H8GgZbVBLU0tfeXkxDg+i6JIgoCuCbiwjcxh
ErvdSQg5F6usHNkQ3PJ9CoBYM5nC0kw0Hms1kBQBaqq1OeH8BZrJtFzBiHze
0OvH8d9fDavSDzERCsAgfT7HxtGnM0/fcm7oQBRCLF78VhKRqNH0EcspWqXC
0Zxh1As7xROyYHpuu8S6VIA28Pu1nRQhv/NjF8JTZ2r2EkVTfexk8LLTalGL
fbkYD1KDwwKvPB+cUd6gpEBxNU9n2UvER/K5ucxLGj0QgOYFmU7G6tOzCaHH
LO1AovrGOfESFrgsHqruuyxFVkdB19nn8HMjaHE5U/SHbGxI0nbe9tFAdTY7
ArG9A7DEDxEJ8jJUQOH+eB2hTYPP5AwWQGISkY1XkpTwkLfldVnm40a8DTOA
0K0/XsZw1CuinzCGoF1HzkUy/fJQMVi7kjb2zKK7+6tBGWY4ScGd3mfETBtr
loULKzmDzPyqBAmsJ+S4r25FDHqvSfXxLbplfQvfxqSQuzs6ZhuL7P2taO2k
hf8oGfIRKme+KqlFTn7n02de6qEUYWUZbsOd0W9S745jpPjpnehb534EEAFo
R6sqiRmnJck9tKHjBl+SmUOeCp3nsTJxVPDoiIusn20S3bbh3q1PhttN2Frr
/cqRYgct2CNE93s6KRW3r2LMKlmM7OEE5t4xlZ14NqraxC+ymeOq0WfMpt7k
FIGvr/Pf4udFI8zuJVZXa1d1Jxlk+M0RuzGTCZZ76Lhp9rS0IH62n7BNZQMf
cICSf42T5YbyxnXcMHaXoOFzdVJmblei55JOsrtYAifIRNb5QMPUu533PoqA
mtkLMnvGGJ2FDtTARcU85sLNACBit5dHAEszYyvkF8bUolBR3gIyacMVX/u5
uYMwxv92e7DNkZ8sZBC2YLG3+mKgk07rYeXXT9uvH6pp5mHWU8zHA9d+iC95
lgraq0FfMzBsZbRyUFTMhBNU882SwxDqhRVaS2QTFjxgJKTpgzOYiOfTLhQU
C4nA6cPGTW5y6+dWIOq9CKrfK3T7dh/zSN3E7GCbQzlxQ5kwViVdQU16I86S
PAxk/miMCnBGXEEvQNju9gOqyvYXRURsz7nv8OAtPs7k/3GYrqUbAan/0Rqc
JcDc1/2cxqnc16GUJTn+8tvL1OUKa7oNKz2Jm5jhwPUZQ4AQJE+RnmFwXfMB
0RUv3fCaprik41X2rrhjhzDyUrEfcujc/nLnvTxBTcLv88XlPFcKH7vzQqt0
gLbvIS6SVg4XCUXd7r6OcEWmcTE4GnK6/nYul2HY0k8rMqOBlCOWZhw1ZPgk
10dNXd4kK9IFjZB2/mvnE9ciTtYEG7oISrm2jphh/O3eF08MU5IYSa0cn7ED
50g0uFP3uomyrSh4VSXZWKgvCvpaZ52HsB6WFpGK257S/Y36iiGYw8OyyUXz
V1HqhBjQgf9XWOYWSAVQ7Yq/wkXLOZbW65VRhle04zVVynDP2xkuW9McL2L+
Zw85ygmacn1WFnw8lxX40hEpOT0uBIiufDwPtx3FKdX3h2hVsuYMppv4OWex
yKHsegBSB9pzLdyx0lW85do3nrbL1wISg+05vCUll63LZoLWblfuUr+M1x+R
DDLZDc86jSQ9qgQLdyQMCvrVsj5stLzVBmf7X1uWep2MmwQWIbxWJFHv3Oj5
n9WchZsEhgd40yen2EpY96JlLYiHIH3Co72Lew8E7yfRhgABiP6Fx+AO5MO4
GaLz0O4ljR1QyLph8097P+ANYsWt2HYAYUzG8YBwTShcxnRT3Ior1I1jxl5h
biY/UiaOf21vXb0ohGbJRx0Ed+q+umWMIzZr6bjgyx/1q/0bTET8PZOmcBKZ
pUK0r2TPDN5OW2+UUTxIqZ9Wtnft5op3YiRaGdAnEDB04ejQXAgsLNRaHZ1O
mdpTdgxbHIWPYhsuDjh8kP9z0jxSwE2vsLttjzqJ0wj40L1nm/niSiZxeb74
BZ60+7My66JI3u00Vvy0B4ZlXHBgslfDluFL2GtRFwzWGwZhag6gD0g15O+T
OowARTrZdhM4LlIeKClYlCk9Y3WAMA6nfUMIT7UqmCE4zatcqKq3QQ88PLOT
12oCddCiOJLP37H/wKY+m1aBwcpN7gniG8EuoSCTiRNZc2N1vNzyYNdnbriP
7NGyBpHg5uP4Acg1jJn5MXDcggZkEcmXEiz53LmOtxNMtMX8o+phfOWHJcrL
KNBLtZWPXo0VZYwEojWzE0wJ/96ypQpDqKdG8FlYS6gaDw8cfmyUVFWb6Zr2
h3uQdcoufOkdtEiLkl3fyPhmW77O7fZpW38rY7vhJDey+iR5TAWA3tMFtuKS
61bXDkO46D/8CbUHDtjv7whQNcKNjY5jBYCOjZTO5VqzNQho7TqGRL8PG7Aj
BaJ9p1tozMjUJ/CIpmKoZJq7V7Sg9h9jk+0bsxxPPPXCILsjVSIa96N4Nil4
eHhlKTb1H+wsqu5Arx2qMjT7AFk+xHZXIINv4Q5goxZmj+nbSlKLTpf4JHZc
JXDdCRa8z7l0myzxx02phU5oKS6vQih8byRPhzeDp1JM5tTndBvMsHY/5T/J
QljeccXQDs4OUltytOhoXam7p565AbOvzd3LV3s9QqiVuKC9LNACZRPTVlyk
cM51FOq4NmtO7KJddfuImMcT8funt/QTwxuFLFu+7qXhvwCdVqCM0F7MS088
iI+LqmZCi0KjKQvAn0432vNQOTPpOSRldr/MJDtiw3InEBHU0A714BlGij4S
BARgTBcjYLfQ2Sz5Xjlqp6rhwlh6eUK9g3DiX8yqKsJVjs4hBpeXUVXRClc5
1fl1Gh6Zlq0mLV7IaMsGcATCKrTStKANt6tB0aptJfB5353PAvWvaQlxJYFN
MmH3huoi95F0o+YThFcsrhZrfjCjw4sZe31wsQVEKKdU5dZje/0EC481VRyb
LlqeZTYe+HU25GmwWJcfeqE3tmqQCCDOaJwPcYFAvX9K36DhJrcsBHd2t+So
LwpjkM7nsJm21spy99mu18Vo3h016l/p3xlsrl9NH2EBZP0mBekDwMVBRVjR
2P2Xr9JVkXbJQqnqyoDq1YmobvTWRVFgSkPvhokO6jf71jFi1t6ZSyjWibyu
9vasNkIXrxZ3XE/4CVhW/YqJ635iVH92dwosVAVKovsRMdIe0O7wlXRcm2Ju
KYnO02sKBBkxlOFTA6JmPaXmgqmkW7Bm8kyYksIiz24woOFneao+mMAHUaHj
yHqJIjnT5S5uxUDGLBFg8H93bPfowcRMk4a9x4NbAl+8OJFKqZkUwP1lZnvX
ZBeOa9MMq6EBhO0mqbL3uj/rs+vkpUaWXrO9aI1H2ZueRrrt1CKh0rbRtEV9
7w+nLUZkIHu9Kpof+mncJ3tJoE0DE9E8sNTSB4RN1lQgWBGNwrthaRmo/mR7
4zDqaCkmx02l/fr4+gGUT83wllpo6xEggKIJvRvyLJcNVxrauo0fSqh/5SaI
Veeizu1QSgdCf36vy5dAET+CHg2fvFxtsj3X49S+a0ox88KM28Gt0t56pglh
u05sjo8yoZFcloALoYXsX1riOngbvfdJ2khovz7kg4NpNFYzGZb0GI4mzbeI
LYKKU3+KuJDiDNr7YLfzZAU6SIzyv4PQw2UYsUEufJA/DJT9qfT2QZquWDL6
TqmhqCk4fh1rNQvYioree+cxNMiBDE4MkwrwiteldEXDT2q9VW5cqTH/Rtgb
rLdJ5JHwrEYGUWdOw2io/iuIoXRSrlhieZQGF2pOselk1P4MoYTa6iVvdihE
roCdbPgrLaCzQpCqOHr8UZeJpCNNlbMGSfrCdpvR0MuAzXrc9g5RZ2bc0fig
Ow+1zFlwmtiA/+R+xmKbIqLSxk2czWVrSp1ClXf95OKVZum6YgWdGf3+Ugl3
s4dDN79Hy3+nIyVlE1isKEfhlHcUmmasWbFu+M9hSxhDIaO2mMCY6V6p7tda
kyqF6sivRwMQZ5emdCy6zNmo857HZGNCMfgAHiq+em4yOCrGfMQDBybxPkgb
4Yn1o+uMDrYWGn8hOBxs53wcpfulv++79bp+Hl4P/1ISnjt/u9fse9wJPKVH
CE7R5KDVmGuAi1U/QM+LItu2n3munGmorxUzkLZe7q2DvkMMB+brPrc3SPQF
8FZy0TH7t3XkYPSYoP6pGdZvvIQgW1hbgvM0ZiskbD+E7kEWXpL+A9GMbnGO
aVYmvV/zht2sGAohZbmQsZE6Mfh6PDh5AGraDmEUw0YGxFPXSCn0H4QG7Q2I
GY5y9aQyiJ951auujPOZvKYtMeOG/BRmYbQqFvQMseOOiy62CsE9REtI2btl
GDEHlgBzQhx8HPvqPeZwGaI43KJye7SaLW0RYoVbo6tmvo6jyrUJrMFTcbmh
bDctxDmj5R/Rg0/m3ZoG7C5mUOKBJ6aXwkiHqw4aIJau6JbwrsXG91n73PsW
0LL1AA1Lyukxbq/OzWkXRmBAfsx8VZSDfmnRFKsWvHv6e+Vu4MmCUkjlbEOn
aRURokXjTXsybPNkKXL/8/3psPaiH9N+XxTJvbs0oWVD3Rn4GjTBh4mdfPb6
orjrcKzymRoLLDVmSH6SyaVFFJU8pEZ+5MJMdcPgU6KbO2X9wtfKDhaeMND4
W/X4ChyRucSyuQjQ092zldm+EAVBx92LmC08Ae8wNhAMhMlz4kfL4EMif3Bv
jqNwCi0Yao4dhOIOy7H/6ca79mhTvAOtsDA0PYE5Xc+aeoTkiIsbhB3PS9NF
e4LA/h7WjctIdOZEwHzAGVKAnX/ldUNUuWhN0qhOy1Sf9/51c305jg2jcjV2
mMu1z+wubDlSJWHu5xA1feLTVyANpLVAXiGnWlDxSVAhYyv8SxPQT2rum7a2
5PAsZrX1UAXZ0v9UBprLIhrgga7sMwiw3WZpTkyLTaTZXFFjznkEXGGpvC1j
qLyB8sZ6IuvXr5xObrzrvxyhk4nfbrPXNbnHCK764Ho4un+hIQK3nbQnjoO1
YjBeyVq/zTbLUTOUTtohClVSzxGpMjp6yLCp990pUH/rQNYoMCMkoeNFZ1nC
qD88hqZ8NWxi5z/rVtbS0NM2+NYyQvEqiGhg1vSw4Thy4pFABHxG6AC3NOfE
NUrM75GU0wkzqVb+Ekx2wlE1zzRv/heVYLylb7RG0WIg9+caQyOiOfcWQ63Y
E8xPYQ0mZakF9BjkhqHPELmb4Vhhz8fA6PA2FIaoz69hiodSNokAjXXtxx1o
1B39EP3SczTO4JHUdgror+JYjo6BmKtzj5URgivNUCr1RAXhCxkWhZ6I/aaF
vNrCARmnnQE28AGoPvjR4Yd0AEUVCNIA4c9jmTymma5GZCf5w4WsHn7SJH30
mqOZbvbZsDuX6JbwNrkeCfpvFWBwMF0EeRdCpceKSgR2JzSj2ypqPstX1zzo
NO/WAFSjTvlA9hEdkpHmgiPAmViqvdCR91geQvnvqlIistxtWAccVrt+V78B
P4WhCbVZw7+rylW1a0UedBPqwOytacymP7T0MIZc/1zXnX4dqsn8yoP1jkO6
8H4p1/KQeoX4VS5G+UnBvpJXscSbQN5XS7jNrZrWJCZT5m3A8PesD7iYxos1
/aGjeZPS+W4aDVTQDZ/dx3rtEZT8huiXFSSfZTNlABFmHOs+RLoBTo8p0BKw
g0zPSBoM2CzCkGBzHFc/iF81Ib30yYRHLjsFkNK+X9apzcWHFoyk4Lw688AZ
NeIoEojpgNDPiqT6d1ayV5bDRCZNmmQlOpAGdenMtRQkSL4myx+GDzAhODIO
9HilITKXW5sAfm/b8GaiPlIj0VqQtbgemBuewHYE8pdA5Ghbddrb3i8jSu2S
CuC7aVAi7oow4bL3nfzuLRct21M6T68EOv5m231aq/kmK7INylsC5yBr/PYn
iHDxsudkxywGEoPv4bK82niTLAzSjvEfLJ1F+BsG5IMKJPjEMIkmYKyV9Owx
owuVE4MNcjrlzXUaPRRaonCSd4qeyZtZzrGp01k9txX/keLKGs5k2zYKyXgD
GmBhU4BVsm+INRizAv0f3qIva91eU8/W0oEJFx8c/+hUBHnRaUUAr2eI7Fjk
I+iZOfbYgRDGXmiuCvfTWTL8rf+GjU1C7trY7tLGoeGFeqwiIaalH3DnLBBq
K+7nnmM4LUShWSV/uje89ZAFO71dUA+kdYO+e1NvTHtfWB5ErmlzSCU6Aibg
6CHBzK17JtPlZ6XPhNdvfBTFXuFeLMf6V7iEz/ZHJ3EgXXUL23mmRKUSYbrZ
mwf/mujvy2D+0eHwhyZYnDHPrn7pb66V33EL8GUxgjL4CODwjPPIGG/1ImwH
YZBgcHYd1LcovAbcCa9SWhW60Z3MI4rlJmd2F7tyykr0c1Sv6rTV5TxmSAyB
ZVxDGZe5LN+FJKNtU1CQhuO3ZnJPY5mbII1Te47xEzkJxw1kEew7SuqVeL+P
ElF1HFpVTt3SzeglTQaohtvCvAW11PxMXrTVwATTkpzbx8ej8HqlbNwwhgLn
CbjSks93yxwRQqdGkoq6+WkPNrM8kzyfEAhfogYaErPryLrdfX9yKghVCyQc
viv10w8/Pfe6WjocDPNrqntDppp1QEbySZgB/6DpM9l16vWCUleMgboCydKz
N8yx4ANHo136y+KQxMmYIdNwgFVWMh9ZXqUm3slcMBNq6Dm7xRCHByutTzwI
sf9nOn9y2JsyinLdMiINoouD/MM9A8gaVQsEMDaIHLY1io+wFR7ENQwzv9R/
oY28FvehQ2CWOoSIP9a9CtlhpunVwKPki25MaRuHkHkzmLdVqqTIPU2sMkKA
6fKxCKdYbNEz0N5PuGLFtqgjWYpVZFbO3Y1esYaDgAnl2gqitJbVnD1zLoAk
1iQxD7LX7m3AgUWgB+3rZ5i/CB1bNi94yOHPrH5MM1Skd1ZgzN6vNN3bKefx
IeWnpxFqMU2ZsjgTWZxu4VarPnmk9qXqNFJzRQYkjrydWScXtVoV90Si2VGu
cYWhHhQxQlKCIf77ozk4FY40jrhVdi7/IBs1VUGkk3pHFjQiAyRNwXFDcb5Q
ka1QNINiB7lohYCJCxuxHPJB6g55ZBcC9vq7hILscxoQwK1ZxgtbL4D9t+kA
O9edymrFgBhs8dfO6Cv17/4+e7V3WJvEq/z5K53K+Vx7nLI12hCJOm0OGLn1
+ddvOgBpELoYExuJpy2mbRllbJrDTj8WmmX3+a4AgFWl1nko0fBkYFLO+j3l
R/L3Y6qOwWfOqhStuTC3f5ZY2gjSQ7UEZWhfcKw07lBWCwCenSKz282etIBV
MzIKKnZI9SfdALQzgodd1IThzsBTkWGnUAYGeO0XrR3QQFUKnPXDcgm08RQg
vG1rSwNhXvKqzVeTgbOSfdweQigihle/XHYC3J0xPE2u0ZhdQt/v77ToUGwe
X0yNTDWBUV+x0XC3WRFIRSNJtpiZS8DihgLOb6FxHj5EKLtliEplum6yduIn
LhvWaCleNCEf+4OJKBz1dc29lB6cloNhcxjYjR/32DKV0q/5HKUbDRw1ou77
3vK0ofEWASwUqdds2M41ftsBQcYCatTSNAfpCYjTFR0jZaD9vYOfFum4HkxR
T58uCUptbcTxl4Wx0vCe6zjH3KC/WZbs4fKvRTFI3+nQTz+Sjh0VA5jA8eHW
1Tfp8oNdgVNJr9I28YoW7v94NkTlds2mWwd8fJ57im7a0+ax2J5IZq1n0GY1
SYRmLgtLpoi+hIRs+0mrjzxHiiyegoDvnB9pdjhU457wJWv5/RzSvZDkNLdP
CLEvgHhViTCAmrQUoQbXi7nYikxB5TdvjGUss7HLCdHsJ2VkUzMKzj7T/0ey
4qpL5Puvj0soW8T9WMpRJpigqTirgm1PEvdhQc0Mn+dUElk/b5CniF8sI2lK
Sxhy2dyqTtrAeBxOELD8SUTyeJImhfpMP2yy7cV8/tfGJaBL900XToc/96w7
bo2jjsBmwP8R7i7HPJduhWNP9HvDXVx295Cw7jFSFGUeckPZpF3+aRFhV44t
qF9YG26pFyKdVgpey8ShlyDL0oBhIZbofe9yH8TIoUUBijoAyApYI2DEcNg+
FjGeJsIJuejzIicHrCmA6YJ4C6zYsJDOlOoiA34mYZi6I7j+uT8Z6qHAtaP3
fdJacxgBGevB7iLSDU2l3O4/iT9jdTunE7hn8zuIeefUBeRSrgUYk4ZZ1WNy
zrGOVfC9LtnX0niJZK7JjzSxhgF6b+92KBf9l43uXltD78tqjq0F4Cx9/A7L
z9sbMyQw838D0km1jqkasLq4G+is28CE2DiKcPa/07HCJFg5B9TSDkesFwXn
qbJ4gQsPBLGCQ+mhXVDQPnKl7+4XqtfZoC90S5dllFYyJzMfDEzauwKYAbiu
jTL4Kf+5DptcpasMyLQ7U9uNeS04926iZ5+Pk5/SpHGkOnGq1Sz5wfpzm5FL
71TzDlINlKsDpW7xK3GkoSUgYPy4JtMm676nNbH7ITUjXj9GdxWjWbEVj2Rz
csJlOipMUkYYeg4ko6SZNViKjTRWKvNyIBPDbY27sastw0vKKqWXq7dVmLj0
DqKrTorGYYaJB88l5D3kfON5VVdeUKtct4qZuSrYhqUPCNzxdQyIn4FN8iLN
yMB++7m42sZOLQy1/krxePa2CzEXCAeGV0eduihLfe9mCbRNPBYQ2mVzBWe2
GPtp2nk14kYQOsqWw5okrw+heP9Kyj4XozyRUJcM8/BNpWfarFDTP+D8eJPz
xlIGflE+jccRAhp5ljGWLDWnup5Ql9jKx+3aHSNSgR3ZVSu4QWLPJfSsFLI0
rN66qIQamkvoezvX1/R5xWs0tPIor3RNbSr2wbfY4GBhCflT51FD08LJj4TH
imnt2kIrOy/TxQuAI8NO2vyXMuIVHu5LN7Dv1ZhTMa6ls78x1q2Aws9bS2vL
5zPjxTUtp01qQwQamDqCX80GTr1Ug5NQkdTCIRA784pCiT7v3U/Gc6DyMyW8
28WeQtdXZ9D/iLZJfJosLxWtO4tmHB1hOtlvLsza/XX6DHJFgAMRjqugLykB
61c/TYXQ0OTuSj/2mlHdxnH6fqLgcqfldJLQQcUxyyqVgOAUUdHgic/7tru5
woExiE/yYQ+k5vrTp17FP5Qf58DjkgFhCjWkcQblgZUGB+RzhXoz9X/PQ0H5
Ue3ai5m0pa4pV6lFXcOI9UIjDBpXgTsDVyySnL+zqj0ir5O7dKb+MHGwsXI7
EygDCT6iiYUDIil3LLaemBOGlnRnSNxWtK2ByaYtsxLC8EWn1MAujMyRE/bm
Ycyg+Qs7xvhEwuqJcXhAJfWUeaXy+aDfa5G1R5ECHARhZlgBrV+9aPtaYJvD
u4wspIiiqyaEfA/XSrgoPqtJ3iHJRSJNnQvjvH0uxK7FiuRTS4eYSA+NUTbY
BZgkPjdFk655b87I/L3h1zdp8B0tFjO7jbkydCdd1G/Sg/BSJRBYL1+PcTFV
EFf/b8s2fWAAxD81zI9H6IvSRBUUHMDM0ut+SUse+n/yncEafKGEBcHDxRQy
AOhX9bGisL6kimD37CoJd+vvom5ivrTtLwPSZ+MNzcg7TFlHEVwVdOWd5b7X
z0KPiAU+zIlV6aC4bzrdRL1s0A6mcYXRNlVsPnxKfToKXKt9qSmw8w5jCPkH
hSSDrWLO4CDSz5r0Y93L4s9Nc2wmJogePBqPmUELKQeDwEGh3BpeVgfzN0pO
OCYd+stEpY55+tK4r2fOzckF9dahe9Ca+ObTkn/jugztirzLSmWaO7dpAsbD
SWflfBJLDPRumIJrCSt9INAxntL4sTo8qWg+lfPX2htaPqN8CePJEMpnSqm0
+Ql15aEeRTz02kRL3U6tKDvnnI+0aTC/6y9qNwqT9/Tb8+SX/k7Qe1gDwCjb
CngpTU1NIzOPBs2hamFL6d4b9CfvnBq9tz7222g0hpHEsyO3bQCm73qW1VSW
M192aLniQMuQbqZRlWFBHMoqn3HahAg5PAC+9DYaKye5z2LLjlZ3gf7juzED
GJiW5fcYiVv3TEAsrQCTUNfER40VnJHpfIFlINLCdKZHylnvXYoK8+VTHJBg
fsT9MlxpsD/7Z/19WEkI1i96KHRhB69vnFoWuSyfNXBfDQOqz0JCTr5m49Xv
kiTgpIOkBjA2wtEGXLUl/b0DMFoXi/S29cSJH+y4WKvtUSpOkZXV5xvxMqGd
szWgmnk7L3XFJFUBze+C/stvtvZLHB6sfXkpSgDbOuWIzE6DMQGekXsoI62X
NraQ5QY0eGLmgBDC7nIqNETMjGdYdE9cqBVrioSj3T1pjEL3srm9AEj9NbR7
sdAOBDjb+Z8XBQbzUKvGTEk/WhqrQl5Tejk7tHK5bocr3b5ERgSLZhdTqMnU
Fqtn/f+TqHyAUEoK7bMJZB7aNU31NEXRKLypoPEUhh5Pti9Rl4mPlGPfX9FF
HqFLtciRY7dJfKffHAwlVJm6beyELXCdsu/TMbkMgJixlmTNSnxxUxn0NPzx
fr8PmKm5s8QLYYoEuCI9odZ9sthREqwrwEdhThoBdpfJZ4sU1iP6ardRmTAi
lddOkjQBKJmv4+CkeGv4hjv0td8Q/nXdW8XewYQooq0zbolr6aBMQVWOYkRZ
9Eb+9xgh5lSlDHIJXS4W1UMC6XW+YUQF+LaEjmkTP3Q1+5HftBZs6qrfh/Ab
A45jclnDw0YAhM+FKEkAiz0/KfiE+Uf53uE7K907UClxBxvDzxhoOIv3UWXb
PwCGOsgrwn1nLcNEAG7TiLISf+zsKLvPoDeL+7zSbik28P7iWp6H2wSiCCLW
/kNR7Wv9bpeXv5c04cv2SEa2kloyO24kzidAnX8TliVQcyXmC1QdUWBpmN+M
Td6vIKEYLqEJGouNwzqMey0/AKIzZpguV8Q6Uxg8OeSkdFhIsOVBY8hKNOq3
aQVofjMZZ2nqjE6+8yJXQfaZk16kuepN8NRU8V4ngmLogjJELT+H4mhF22Pf
0GBec/aOHya6jkalPNux31vIjmm01NwAePWxIaBFaHAHX2ijm+Hr4THawa+W
hNV9++Yic7FZJEZnc/jk0hbtxMIfhZWfy/Yu78a2EFldOBkhpOo/wEoZ+RBm
AvOqT37nmKn8VnxZys43XU0DbStuJlhv233ZZVu9mox+4WIaMY/GI7ypRh+9
7ivqkcCNu2YUI9U4oiiR6+W4/WwpqVPUEahFY14FgWSp3pVrw2pSaQkhWlMT
UKv6YYUOtTZWf5o9Z7Rvb4wPGTMyLDD4KeBafe7dH43IgM7SBinUKgQssQhk
x1Akv3TTbayueoEsAxfP89B6KGpLkG4rMuaoRO8vS5cQvMS5niVY3FYOLQs6
foH9CmB+F9dQXGRHA+znfmmRved14/cpFXICG1b7u2rTjxnk1WJ7zhGE3M1v
ZJwU+HtnwRIWh6J+jLys3VbBK4QdNu7e8Xmbu1YSwPgmp0mBfvQa+3O0UB9K
UWbCxkFIOGcanbWunoGcMVjApjASHWU89GaHZbnf40jKfK2xw/9VsxJ1pQIe
ixwW9CmnxaGDclPy9ggNCf1ZvySR+UZiS+mmpi2YU3kQxRr3a+V4eivcvIvi
7lDJ9OE2+4PBzNVCBK52Ks2hOSrxK2rO+actWGKfmvZkIw20M3ZzDvBlQ3am
kn8seJlm1AbYXowomIqPjM+WQroAXFw8HlkK8RJYPHNpb//lw1MXrWiDoz8b
Dtz4n3fL3o12AmLQ9iBbv44PbZ17XZFJ4QG5R8BeNJ9BueHG3c9v/r0Z4vgT
XWdfOaWDs2+Jei3pqIWyDjCULlD7eOhLmoQKZVucbKCL+MJTXP/aH4zHQpUe
D1z3I+aTK+guavy38tnWSqwSskG0kaqpuxiJeYnJXIZl+sskKE3wkN1j8WVW
MEnVZJBPPkA10QOMKzyoTnrxrbK7gYPEF6JHkKePaXtFtgbyx5LxuCTTskZ2
3f/DJCUmgE4rqHCNstHulcg6XJ7aUm/4qgtxHZCSariEJDKE/TWpqXk+Dt2g
Tn45IXr9rQ9mwGQZIo8FvArorxRfTX9XmaOLx9XSzGwDXZnMCmFYyBYfiz4v
SqF+1bwOeAQ5HVwhwrwJ+T7IfszfXXvYrtdBgCXTUUuxuQG8N31NlHDcrFT+
Yng48H9oK/V8MjqeYcdrQIsQeGvjTKa6dwMtQL0vOSwZyNXSX4bdh1a3yjNX
WzSZ8Ty9KPSV6usbA8e/JEQ3/O1BxUL4prH27hHg19T/Q/3LgrH2MBA4WSMs
oCkLxQiZENgsTuUPPklaFeS9Kv2dpuYt//mK/XA3WMTN0C8vQvg+XrLe26sA
FDCXFk4jTIj0Kmfmpc5evNTcw3i+aauQO5d6OrBAU+ivH3AS8i5C2IFrPDtN
wWGndsBFJaIRpkv+Gi4wxE39jBnOXFtVzTJVmgqLOfybtAHiHw1ZqIAtnWWv
k/YxPeDAnu2H6//RkRNMZftYuvp794P0I2h5jiHGOVBYPbV0VlihYN2DdhzC
jJMl4wbGBWI1yk2ZszmFOHtL7KACQ0hQcVH1tx7KeAUese1DIkBIPcfzdybx
fHrM1ztfAhPg2M9IEFvlJ47uErtSSH3Qxe1RF7ZQuK4g9cSZqVA3abVT1n87
iSs1jHGXu8Z92OyIPSCiZKp9B/5u8L9eJODZTme+oizsWEdbebL79evBAvAB
nHSjJMCii40SMXi5kbOkthEPaBPiTwZ3mtoz5y2a907vBeRupfDjJpjC1ifY
TKSi7uF5b5gZIYRR+KhpqR4cmeAdKUhy1p+7Af+6bjdwjxjX9pt8LMOF2SVa
F2WW4PZI/7DUf3/cQ6tvyXbelbs4eA7qW8GaxKmHFIvfH9fnSGsPOXZtGBno
gftXvSAzXCZopgYVIJWI/QLElqdrZf0vx2mrIP3mJoIZX9PgOmHPi1OAo6sJ
BMPjerBawgurj3FVBd7vPUJPHaS7pbI5hmQ5HtkSLTNdn3thORDnfaRCs+5Y
UAR7lA39JxX1J3jopzqdSuusH7nz35lBd+Na9ydK/3j84n6w66bq/c4dW+av
qhzdhxL97imj97/aRoi/rWAqbG3kw9jr2hDf7Jgqgg2IoKOajA55PUvQg5bA
iWyNdZLVDUzG3lMNmjZuRX8CJFk+OzFBk0+P3neF2/waYA59GZ2ZqU4KqSGD
UHolyyx0skAMTwPOgH9vIAZk/QR8CXqNv579Yq0VARvpMvenEs0xnu2cjCS0
td+vEIGMB2Hnk0/XMg+/dxRRyqPY9lu5ftuc94ZW3d+gjIy9qS05s85iNcb1
/3yIhvVB2lQIlmgfFLSYNDK0eDaWAtlxtN1R9KPx9QkX4Zrqp28t1A8wlnQh
FHA2ebkKPMXBU5+ZE7nn/TdJPAhnSuwI93/7goAsUj9+BpEUkJUw4/SlXKeZ
wZpFdnuAtlqrVwmvJ5Xnq9Km2NO2fR9uw/SpALWvX+4eDQne/iO0KEZm/0F6
aMTHc44wSUq6tkMBBrdTSIhOQB89ezhcwAQJ8Rj1uY11j/V4Ux+wZIrMJ5xQ
spgeuS/QbDbdxL6tj+n2D6K/H3PS370wuLSuk/mytNgH/iUSMaOZDRnNQl7y
Dhr6ArBoMhZcF30GJT5xOQoZYb517j2BvpNBygHQM+fEBpLcyXT9b+llFoFY
sNNolVwGVoBVnX1lpJ5jEvL+ilvXNDuTExRF9owf9OOg7M6VMddx8sX5rXvR
XGaEm35onNXCJZaiAHcl0rOphe0ZvnkNaiSwKFqKWzlGRJhmLPFe/iUvu6ya
VrQb4DfDQIQq8Rt8qPDM/oM90+oZ393072XXDU/cscMFJVYeTUt/cpipGZNV
kQVFncb0DBbkUoLZvTmwNrZGWj1goNSnywF5KgKxhr2yB4Y/DXjAPj0dissS
XVjmSM12vSbXAts3xixUXhM7XrVG3t9u9PaupEWM3EG8ts+IeexcJAgkahpA
4+HuBaCcw0n2owCvOvW8uZ+3T8P6Pr9Q72eFms78eMrnC+DQTHKiI6TSAqMT
CwR9bM4+0rrQYlMY2lcYLsLrqLGJ6rA8P5RPOCt34i6bHsrqHpKg4+1rF0Lb
eKVRoVbjVq3h3KQVAtPGoOFnJxjUzyXuoBDN4aCici6XeZD4eQfhO9SeSsrg
wp8GoAwea7tq3WbXpRhjcqojhkSdICvCXteS03O2+cTcnf2Kq2jIBHF/hu2r
Cqsc1ryqXMYxR6TCFdADTS4UfOrRVV75gYLZZCTD6jxfvVNH+vi3ZXLKhDq7
4mVn7THxOAyzwn8dMw7/S2U8pGFi+PsJKGV8Sq4+HxLHUnnSAViy3/4w4hvJ
QtttQ7sdq33A1f0JIgbC90AE76eVpRNsbiRv3S9J3u+/OAAmlgtWnUPDBnTN
W2GizJuVx4h+8uAQzObjRLWL4F8VaEgxq+aT5Vp32enReuOcuqRd6bWIHGbl
tiF3e9Jg5KKevqQmi2Es+Wq4g5tOdAC0gkHuuvaEBlZ86GTryazaxjKEfDop
qcx89jucnE3MG47WF658EoOvR/vFRb92fem5ZmfbtSTkL19AtNZKDUTH9UVw
F4jsWwZAewIsNImnS1Mja2InXkjHAbuBbuIZO2LPBl6M8tLnTK3v+6333E60
spxUTHg3ADuQtgPd7bmp/q6BLfI/BXN8ZAorXvr4kIctVA+BdcWeKdxLNshY
BDXOtq/F1bv5tM69HG8BzeK8ZwfwPN0jNz7Py0m/TNlKcK1uUrcurcPfLMvA
64dwU9KLYDb/EbzF+4l5kzLkbLarhmip4PSwn7TEuGJQuYZZCfnjvinvtZTr
5lojtYKWRYP8gqex6lMqRexxIMQRGVZDqRfxyoeidXOzhNAI3x/pptjddLgd
8ZjI9IAsMrC7b+hWh15vjntmIyXTN339bYcbGdlilF5EaY8CeW71thuWwl7I
kZduGymiHq+WVxVh8fuRebxv+Jf5dvcQLcANXMqZrzhZk7DjDFLF3xLTNFSR
SkIbLeI2L69I5dgtPh+CPYzjf2j+C4i25aG5F+bDmBARVcd3L5no96G8WGHM
/71fosyLKni2dMqIpe+fxl6RSM0vVFdaon3Je4o4K0Xg/xAfCTTQEULYowwk
WSLAwFU5vJT9tY46PyqAN3zued3kJvcsThs1jLW/xYFS02yEJLNjiFD+uji6
nq6OspdihQ/iGrHqGg/6Uuf2GTl6yIqpvGJ9keZRVTr7tQx8rSzscYHuQUu5
r5huguOjgcHA3EwctJPx7L2q8a4br+kzsrMMZBE0X/D3JS7klbZmrF3TUHlh
CWUBJKbne4xDcvLS/WMJetjufeTAQELY444SYZrMUVDjYFZq7so2KG6Ydc7n
DDucNPhtg0nDyZg9Omf5tQ1v+8gpMUcaD+FkaNK0LQPT7+k/aduVZcVtIFlQ
h6ilsifOgZ1RdJDInvNEteGbwI9e48BIjYi1ofd5RaJaRdXQRonLDMjF8Y6i
cnNJPki3FIm+fsQOZanjT2yxkxhE+cX/+Xd8J7+2bVYOLK+JMnGrwYaCGzVm
FkGmIg0rUhKalflq3eTpungLm4gC1PdY/qW2136wd/OcI8739F/qo+K8Yr3a
fQttX/Tke+IVka7vljaod0w1+2AX0qGQQfvBKlMNec+CFMjj27OY9qqng5J8
ZUIq18ch0w8BEApL+irnVkjgHNf5D7kKVl3gUQ+3yC/h6iVYnCCT/axv4/FV
of3qOUJAYvN7qTzmGnOG+8JAMyLbZC0RyIqR1/j+LrnN/6ndHn9dJefZTJL9
R3zpSuHrjVeTPxjYL+ap9XACwpzHai2xlv0+pE0qHu0JatXzxrkZuNVRjMfn
eLsvgrb/R1u5LCfRNGAIPpp/+BpxiCRnQuGP/dRf8GnRQYHnJMYHRboib9Kd
JZhWo+/qPAazWe/2KE4b2DW9OYYA4FGxFtmmU+i8qYkfHCj+I9eT/w99xoSn
iAHv8vNIKZL7sdX+a2Ln9smVVp39tCIEtqESmxpCH2xAhC96HDKe/v94syOe
0LCB9lFjA1LMnwp8YojBGqG5QJwfi8AUtcrAAjlo2KhUXJBwuvZrJCGxfSD0
XQWWdSAIAzqFAkAubFGSX9b6pR3+3h+S0YiqF6vM2BC7m1awaMglhN/cuW1p
G2Gkgom3XkNI7Fu6pz/UYepq+19vp4NZwAJw7qLqNB9YYNkav3S2mn+t3B25
YOl8CzpiOkf9//oPM+csom+KaB9YwwXqIThAzdGv2UtBYPa3g4cCQTdafZC5
bt/NUtJYDtJnqQ5L6mTiFLMOVbL92W19QwkPJyRSu7RHt4bIVEb0xfQGe0pe
u59JwSP4xLokEu38kFnsMmYQSEs+On1Rt7cyMlVvWE0gfou8EGNLBAjZ+Den
qr4LMzdPKwjYIOfxUBkm54MOnsNpfsI3GtHRCZr+zQycmaQ8gx3JzwBjYSvK
XZySN0j4jWcn9QH1sz1yahlhvQVzFV7atMrm2gWoup+ZyEhRTsAYYa28gPsk
xH5Rk/J+WZJPH7hODG4sYJOyyfGj3KJJkGv8KzGJoJnrDl5X+t47DKga9L7L
ahncIu8rXaMJCDSo+EDvnXpWOIc2XwhWfl0FSLvIPc/ClnX2XI6fvRSHzBwl
fglvax1WOswr1vd0rtT+Qu4LMa0DBAe8bo++lMW3PcR4qwzmSFp4sT6V1qat
YhLAfbtE3hH4wEj5kIW+sA6pYsYfJF84I8L+l/L4j7PqSwfkHzuj36fnapuf
SUEyQuipJBhPjqvdgoB09I403gTMUYjs9Jdi58O9y6wIPpcYGBWmKFtZy/Yo
AiEePHI/Rsk4ug3dzV9QZNWYvye0UDrXr+Qm4yLANBWP7DteIQTPtsvnHwEc
xtmbTuM3IWMZXMsaspHmsogyQg3N2mdVk82eL4Ag1q6052iftaccbsOOF5BT
yOb6qYUDeFB6wQ9Kg/2xb4JdkIzd8KzAL1f62E0j6+Rtp7rIF7Y7yCso7dmp
rxX87o2Q+9g9dObBfaslZ0CviAk+e8tf26FqE7nHqxCJcy94JHNZxd7OOHKP
azVRKTwLYdpPfqgdEmHReHoHHx/Nacs+ZUyyHJ6beKYrYRONWOPv6+e09PZ5
TdAV6WxVQ3Kb99pqhv4fIp2sCEP6jJTyh027mFMyZvzqmayi5bnV0/9tjSvS
A22RH63FgkWtS+L1r9D7aav+8eE8K7b8UPAPo6Jyk9flciAxzgYn79xMSe7a
TgylmjJNCHedXwZbHOaQG6+SyoAgFOifZ4mggCGis6GyXu5mIO5uVz3cKn4D
7yEA35jQMzOlPCXgj3NjAXYB6COsKzrHoJJ+k0aMLO9k9XQmo9C+RGvcTlvr
o59exWhYDH0Df3DdBJ/R1bOige5IsrL8+pAU5tVbp/AL1yzOrTgGjz/qFoKJ
WvBNWJ1DIPxZU2m1/EtcEuSWbyc9+vj1nzeXWNC+mT0hCPEamU/6VxciKf6A
d4ZPJAo8laAKtAVp3w3AsBk7hZ3J2bSSnKFeNoekmkfzRKYquRCRMDLMJmY7
LgD9NZ4FREgBzSqVEASm/wL3HEUd8vXjJhtdQoo+V6hpgSqYt5hML4PREZnl
OUhoJQaIZhgwgoRryeuXwOceX3ZPByxg84e+y3YL/sB1aq8qKo/YaJcZjDyg
iCeUH9fmkK/8Y6jlJzrGF7D5L9nX4blaLxKuflbxBQ4TcdYVvU1eCoY94Zet
N2K53ikHEZ4zKnii0N4efF9wHCrySim7sNA2ENEWg7SG49BFs6OBnADOUHrF
lIyEeQ5XQ+nq+RAvehWdLIEeJ5knMyeBxZoVKAqeAzLsItPENNGAMyprP7/J
6Do5JrHfjmJCYxjZman2udZnsHn6+c0piPB6z4plFx8hZjqFKmZzQlEX0AJu
Dp1kHhjNV0LbTqZClxCFe5TUv39EMBGLfft4DFrQdewiV4eYcpMnDxx25+L3
9WQ1SHcCnkeTZ/hFSwnqnDA9jRAVmVYI7xVww1EBuX3kKjKEVqbqxkb2MzkK
ufWxmaqzNvSMN7asouPY5f+uTSBvMieaQGqAjmAYMKXZhA06KZspDnPXk09J
LPRyUbuQlHzh7pazmnjCTOZVVW6P/5HkRcnEn/Z7alm7CyDWh5bvEXM4AkYp
/yat7V7U1dg0Jb+TWSOg+FYGFDF6ibPs0jHUV8eMvf3R8W/n8OyjrkcVSk88
QvgAnrbW88u4G79NQ7ACoZG4fWBYl9n2XKDn1cQD808kANlKrhIqIcsUd2BR
ddD3Wjm7bwypiYqn3pTq0xvRuDivfZgpxAlkXYfsVcW8w37phqjd+Qg0LSZw
AEggs2d/py2w+XrZq70KeVCMptTFjt4hgtvJhKxdxa8AxWgMP+La3nPhAekf
Dfdzk9aSCQcOW3chVtBewoVJFVObNHNxSjk8ZOqvRl3kbZlGY/HbmdQg2l9j
GBmS5EIsGio49TyMgOdNH+JOssCdShWyJRPq5hkgXZVcjbPcDm1rfIuSFVnP
sXCV47NILYCPsRqdyDKUhgNRuNDy8hXcu1xZEH+AIOTrqz/DEN7Iufd5ozZX
/jtkg9ExLZUXjxfOgTPNUlUtALnWN4Ev8tdJI0wUU5zojNjKAx6sRQI9rtFk
nqyN4G3negrJUMsDQKik2hcv1FCR2NqWj7f/nJU+pFjjK6Z+xNDZ9oxfiBAc
rJGs+WHbLpsro6NthQgNYLPvdkoK+g4C6LUKsp5AJT1uyXVI4X6cKEwOtEGY
Ug5TKqTzhzgTlaINCGf/B6r6RswihAs7bnTbOyzNjQsK7Qik/2ziLtlRHikc
HtiWMBWmWnowo7Ul3H83qUeGpfdYLyf99ZAv+WKszNELwsQQRk4dwXAdYQgK
tXfjdXktDO+rwHTsYtVN6C7eN3dKbrcxLfpPUcqUKzbdRUW038Q/hndPfSnd
V4CyUBa+/XZyF/Gcx8cTyzEKfNbO8XgUrh1Bmx8rUhU3lA8P8ryKcSN+Vl2v
mGtkMqi9pnF+8hA6anzE1Ny6oUYU+1hRXiq+iga4ALewpi2edb+v2KyPJaIM
R97dM/8deylb0bH+jOvZo+wDxdeEuVFi/BuPby4h63jfTXB/clxCCdFxSMNH
bjjESO+G2W+IVWTFTGCJoEk6BdIvzFOlzWxrlBwxT1o3pqEGfHA/3C2otuKK
IBYeV7NA1M8YaIi7ceO45kmTR99sZaeYuY7m3WGr4gn7vYOlXDeIY04xSZJE
coVmXF2NAHV4EVaojT/6HqEGdHDPCuCRODfybYDmObO34Ry3Tk2Eh8fV/ufV
Hmzd83MV5dpxDUmuAlpYPpZw9qQ7J581ZeqxfPxsRKOKwhJTrtxwT0EPeddm
AP8eqVtTchto4KvWSuv98xs5gz7WJfaYAQxyXDeZKJHo135hGqDCZtnUciw4
RkTQx8l0ttmjU9wtMXW4xYiUbsfhGMaHVU5nC44ZtgHFvy2HEMOjFrhwWP6k
OOZO0whPITt2fs5FIPM/ZgQSuqpzqqxce/NxyU1ncJX3wZr6zAZvir7B+OMw
JCrqIigKMSdGnLBcit0D9DYKmrKUXq+DYxvcgKt5Bf3ikAze9BTY1R+PJ75h
dg64vVfj4Y+B/70v44j2B22A1VjmzCHw41U++Cd2XjC4+37opqxZ7sU3a99s
AFCkhcS5sylo8DQJS+in6WWO1vq22km8guWh4Ga0E+NpCOsEHfoZHbzURl6X
HsW1pz0nD6sXen2WXaGHoD7NRQKOZYrCZM1HSRDDLR+aHLdZAbXa480CQcwe
CLl5eyaRRhp1lr1HGv5GazYhQQVSUATVM2RwfWRYFBm1p28ktTXP1/sqSBWK
VviubFhlc7ZFTfznZTTQLfJjH1KUoXsNVGkDwVsyXh6tGhCjZriuPXVaphyq
GRYYnKmqxG8XUT4b4p679T2i3MyGHA2h7Mxx7Y/Lwl5WgEB7OwTwOw//3BZU
KD1LQvfWy2oUyUWtANdqZ/TrwJAHwUJTwMQDYo17aU0NYaZgL8KFOYrnf2tG
wvJtZoELOn74RP10X0biizxk9DfpMi6Uwr4Xxl7E/URBp814f9bYW7p1jIs1
DfZegdrb1xWAmpXX1LhW2tw54GhzRpL5KxbXXMrc/FXIi/mAXKUnHHWfQAK7
atOHaswN5gMutYhoTzfE99Wqox6Za4FNvfTd39KH6Ih4gi2xzLB2aAPBOYCU
ZiCT5odlWzGJtcQsjgJOtPCecVrhuZaGlUJugGXh7B90MO9Ts35DhNS8oSTg
RXmJlyk06vha1JCF9ot89gbGNBK7/6BZgK9rKN+iRE1aSZXE1iUJ4gOTnmGC
55RAtyT5wJ9do91vwNpsFTqMpE4XvTp+vXz5vP0THOW8ypGHBElgDDyic13m
0JsFIS58+ERecPtGv3Vu7R0rJAjLY44J2sQN2djkHrjKVYmSQm7eaI8JqFye
sgh5akQpUyAuFS223kNM7MQ2+xJNBQ9skXY/dyL72FN9aiWCPHpLT0nUMyX0
DKXQ5Uzbk8CvN5BdJhxQRYnQvGBDee0VF65RLzDH2KWbO3KwM1vq8hoUOUJQ
3AczvUdKwdYlz8Kc33Gs6Fxs+Xm+KCl+NOolMCrzDaPUnDOxBao/SEa+HYEE
s4dwUbASZR1SF+H2R7T+t25+TtUT4ED8b4HEIuKlX230bBpus0mLPNTaf7ff
sVgwtvbc91rm+sO1N9GtKoRRjLZ0A6zUvCIh/Fi13IZK89fcAv2W7BGTwDa4
nCUlBz9Smv+5CH/OYF+sC/wBu2si9m5Le4A3ocLy+w9TZjfncnVWXgl5lL3K
Yw6GkzjqgDgqIjmJyFehFvdLzjDA9B1vcU8JFnl0OYktFsR/R3DVqUlwag+P
324LyFV8y4qU4E5Dk9ePVGleHiXyVeBJS3hdtEW+BEy5sv+4b9JQmC2hwUcB
Z8uXaSInU0snBmLuBxiKd+mH4uFqWrR8HAz5YefnVpwVosVSZr8EinlxON/k
FtM0m4omlkOxUYXJCPQkqeDpaGzTRcR2ngAc/pxxF5Zz1vWWRSk5aa+3RHEp
5ut6NUUOr0Z9zxObiq+BU7JaUwy+Gw+LmD8fMpieL2D7MO/Mz7MSQiJ2RrMN
eUkSLJ0rlUdBAMfoUPk44x0SCXGwsYYbdtOV7xCTC5uRVi5n91roLu35PMu+
/JZF4QyPT7gidazU1TW1yq18AfxZ/enShges11IbOJpXFtEDrZAnK52Du6rS
9F9Ny0Yiqk7ZMGB1fEXdc27DRAdhWTPGKmMnh9EadhAI2x3z/dPF1zc+yaEY
53rx1IZ6oEDoYyFo42Kw6PbWcp/WDAoAJC5gOldEXebzG1GAOYEgeZoc6pGB
u0ispOPG5QEdXvTIT45eLnxLtvR2IRgd3JkKTNPI9spn3kFHdvMLUyvLtW/U
r5XDKefI53N8dRaChBD6UkVP2Oq6LrmQSrSXifZGX6O9rqIHapSj6jnDee/q
SJS5gtsRMyqoeBCdVq4XFWcHg0S6U78DS+vd1QI/rUhVcKlWNgM6XJSZjFiK
ZZ+hJVITV8Nc3BrqcfvGddxdCK78PT6RfmmUCNAzsKLYsOmzc8xawn1B3xvq
TvkW/uwxYLjEPPVoElEpH5fqJE7swot3VvZoz4G/KADa/ogDrlwVM7F6DFey
LvqrOKca/fG3PTL3OHCBKZlmjXEDTkAXUiOkT3HIaxTzqvUCULtj9YuHb/wJ
nRHyuikpZdqBOwhJNQqM6+nPxxpp9D/pe17ANNjJoj7zgbZpjYj9PCZ3oEmy
mv/SQmB2OakRC8vLV1rYwPM0Vevu0kFkZCERQiBFeJkFDOEcM8OrwP37vLhh
IiODRhz39luqZB7rPUZ4gwzyI/2pDnoq7Y6kPXxgRggU35ADuBWaTQ1HJvYL
TumSahrP7Hcbxf7ueDkgWfgsPlqG6SlhZwO2FatwMLR1EUzzsHOhawqtNIQN
BkLNAbN2i1NhQxXYiH/QnNcc3Lt9rurfrxqBJbSvUfotleMtQl9DoS38elLq
3f5QRzP+ZsjT5V8V719ezP8b7X6WS/e8FyRMC/2VANeR7ugezx4IZpRzUlse
Wf9B9OkUJZMYWm/3QMXy2nDDmb9GdlqPzKbCAkT8mId9wU24Ya1OjSK93HdZ
g4ycDeJCQyeS4TnGyyTKWUXa9kepQ83RwKF05Uq4ysoSMJvESPoxopohYySZ
yGdp/6XPKqWOvmdYqESqssCf9x8FIKAGyshsnufnOeFoJPIWwCkNJomCquCo
hM/rFr5M7nB+FGI6nzkEmjOfeVWUIZkomkvkLClkLosQdHaymr1ufkDo+c2P
dSNPe0ujnuOnkdXFxk5B+ob/511/eeJu+sPQAAZjTOHQbo0/C3UkzvWR9NKO
9NoIaVTsRywvfHz1KJ3sWquZa9kE/IYpCue46+z8AKNqA4ybr7taftMFETMB
MrbzV/Bm1xJp5dK0gi5KxbGVOqQWh9W9kTQDcazH3YX70hSMvXjLdLCg96pY
yzSRfVPEe9+wUrmvrZtciYeKDmY9JzuwLoZy+qS0P9CD6b87IcMk6M7dmTKh
84KuMRT9b//FUvLyvhWQtugdOtT24g91dPjlzXrRD8ftdYzHCkR2gcDTHyn7
s89475+n8lCsclctXPvlQnm+2+frYRHuK+Q6NzQBtNweecBMerT+VgqBEdDc
dL00HgckbCqtebhVuLC6QqtFp9Sn+eavLHAczQJwaf57eATjIGfn6Da1uQXM
1ne3P7qzTZXg9e6222Jyf/lBKHA3jNQ8sacm3a7Uawm6ST0ZT5M2/iXnz4xh
Wy4BDDg0nDLgD7tisnTLkLfy8S4yl7ijwZHdgggVTdnsVVgCoJAPqJ1KFiEK
ns/Fzqg13hTr6JRLLncOFkSsGlrtbdv/MN19Vc1hGJxf6Z2fR0r7bvldgL0V
rek9ypiE257mMSWP017InlCXjhy4mbYNUTgJobyRU7uMhuqEKGqWg3KMFSeS
ksl7C6hHUEvEHLxC9iIBwBIMGc2CAP1C6TCaLbzrRYR3Ua3mp5W3MbsfWQcX
LROrEpfFnSbWV2wP+1ORDlxE0sGbVpnSx+PEfMtVMDS8y1tAwHCLqge0SacO
oMzD//M50FFBOEOuGKd2e4/GXi4QXhlIqhSEXsjuQiPs3psM7hgDtBC98Ink
eMfEAYO7iDeXA+9vQpJ+yRazTUhlikwNseLP668mhVa9qCuk59pS2qNh+Xy0
6nJixC/lXKHo4JexeVt0ibtV6buGjM+XCONBWi+/a/+3y7lrnXCcnB3M2C7m
OzHmYP+CuMVpZ6GWK2PnrIAPxzKgBHEI4q/Vn64K6xWsIeh1DfYdwNEHm+3/
AAmAsrqLOQI/dEeXb/xSLWEUnV/wzaEWzZREw/iOU0tXJ/bCEPD1Ou8ujGVI
qhZ8Fwc/QYznEG6D9sSrHb6YemUO1KRpOAF8kGYIABDNCxX+zh4DAsDBjk/Q
WgPtP8YMUR46a4XyjhErDlM2kHV37uqznHoMUEjLw4N7ALiP2V4jRf9y5hcB
LEq5JcB8Bu316qhMV95E532xN+iXHKwqyxUxSnwd7XyprVzgkCpzGUbbnp7h
TalMEmFT+CSEA0oMFZBkvXD7CRa2he18wxiMtZXhavbn8Ygo7ij/jVmMBUwT
V2zV7tkJD63jMAlNckDj1vlXuapbpwmXiqHKeiO073Wg7FdLtqWX30gm1tSC
0iAVnrO3sElt/r6eSisMU85EkSCvDbpvThEtowc0k5LO2MvsNEGzjL/Lm8Qp
7RYertB9ESxNAXvnjpwlkF3SnUCMAHWrPMXcXb1e+KSLn27BzThyZ9CzCOFv
I7z8+NM73VX09gCKyXu+f/kt0t0flK0GvejiafOzINuRyW3N1RRVDmnGtcrY
JXjRyX0etVY6zTZdUd2wzd7OUB/GL/9GjABdOoD1EaDsW8X83M0OGQzmWjb8
rYPWtdTPxC4DT/Bj6Cn6nuUYpaYcnvf70iOYIlfa9Ny6J8W5jLdVtutd0Dx8
+lSvNA+4H2IsGOTW7eUu0LBJAFf6DpsAjk5/Tjx0d6foqxY/FyAZFQTXFeem
QY3XjwIHLGBwCB+6yc5oWEtSCCm2L67uySgfdyLP7Usn3x2vNxg4QHJiMfVy
jTQIH/QQJdyz6ziajCSmvrM+0vc40i3Clwce0Ks4f/a6PZpbbAXQoeJIS2PW
//Lw3AcxMW6Xm0/BMWyocI7RdXKuiPvfpyzMQZlxHNQ17YxH9zP4X2/1+0zO
8KP6LAf76FVSZ9G4HKJ0LTZDjgECj23zFK4z0cDTrKIrTG7HRsg9NZdJFH5g
sSZ0WLyTxSP8WQmIBNU/AalCSnJ75QlfI3DsoNC3Y6jPnpZThLUerX/P3B9X
VRncpqLiNxEUmd7bcECOnqUhgjuniyh9AzNJO/51wFJiz/6EHDzO90mx0o3T
1QkkpsWb87uWZu0FRgqqq6GnmGWDN59SmWCeygdP0oda83IF2ief5WkzF48x
3ccvhfAPc1WN6P4Nc9j2HlRQUR/gH8jjIOmeYRNbw/bUc3+355Sgc6Md20v6
b1zyxlyaPdFuA//qMuQjWMCT2ydFcYj/brak5+iN4OkiigBnEGs1WkieTtNe
PT7RiE/96Nm+NySfkNZW/9LwVZJGajD/ZdV7gddhytCSIh9jPjwC00vWzXeS
jtKwptS8A4Z4yRIl+gOxCDk607l77vOPmxXS06K/ISEHIRZ2lgYnYdDmL1lN
k7GRv7o6RZMBG+KkB09/ndmZt4nZ2jAUpOJZlx/gbRm3hhVLRixbmQfxntB7
+VlR9uQqreiJzxDlbdGpEOnX87YlIAiet7PU48zqDILhEKgtKe0odiRo/Pte
FJQ/RCI4MVC0q58VSgfPEnFpy9msIDFeTtRsKAOoR82CtFoni6msly6yhkXi
lnWFk+4T5dx7+Xn3jJMZKbnG4MWkBJl2zJIO5OZe6N31FpLcY12nTjAKQye+
rEXYT30i8kL3JW5aY6OKgRwqzPwKT2zP+ZkF0ruj65z/rY1/ci0W64qPFFNo
55qIj0XuRcryVutZukQ+vVF0ek7J4xtGWpgotHyn2LturVqcHRoSzuIBSz2f
WycpEbnP3RlwXqbZgyZuEYLq3NqddHTx6Ebu9lUlOL4dfsFscA93U9FgpcyD
8VqHvT9ookmKXfNNSBNiAD0gbsRrMhX1M1RTm7TkEupjo0WZ94pwugHK5BS8
GOSaFWYY9jySCt7BPlPBKDVIr0vTBCgLAReRoK8Pr1KBXT04yNCP6vQ/SlMA
rLfkE4CTwj2/3K+KcrCBXsA/yKGWTLvRegUCZsgH2kL5GABddhPyNOynbOEw
K/ByrkbHWET6pO96yHzp04cte07r4LKZ9GISzeZ3JBhMJNmI/69WtyDtsUNy
/O/6kqQxO8BmhCHUkr4SYf6YYYQZabBtDwG17Uuv05Sxd5p1y2ZuzfIaLpyE
niu5WlKkmYyLYpDPyvxeFeLRpL8PbfPpDWduvqXhxOXV9gUsz+VFVmNTGvg6
JNZWx9wTUx/ECMOJ+hEpz7bq5lDOMOdLjvl/woD3PqZM/jsUhldgE6MYgltT
S7CBCrN4f+HHB1h4wcRKlPR8Jih9t81xmmEMY9tAPCXf9AlD55mBEg85x9GM
/t//BDMis19pODUzaPJ2LqYy4AgUkj/WMqUXYwhTTQXvClEhVhtSfb+cz8Ag
Uk35YIXpZsOGXzOGy4uTDq4xEpLK+wbZ09Tx295o3j3lszk6ZE2lPZi3ngz+
zeL2g9uHag13z+Azrpqn9Y0VrSlMrs0oclQRgojlb93UG4xq72qAJkbIxgQ5
QRflES514JGibymqruiVdAcY6+S2HvqFU1ZO8YkC9Pt/sEI9mIFJTfwwRgyw
LZ7Fr03dmZmZi/1YCxz3FHuH6sWzFklgQ6Rra2g8ZfA79sgCPRUAVCfZ9ruj
0P12asTBKknwqSUZUiHHyEJuatD4AvIfFWIbZ28Op0ssWMs7/gNhE30HYNsI
635jnz/X73FM3wnBYfDvypHq7zFHbBG+YNB/CbS1Q/Y5Uq77r26hJ58FOdC0
srdLPLCWJUZMIHJTDlY1dU8pBH7pVKRABi9s6hjDSi1Jnp0/qt40xMEnAEu7
4cZJ1CQtwl65FjPgQHx4RPwVBaDOtvk1wVNF3ocXBZ0JZT8tkUrE/54leQq7
b6DwYR80EvSv9oWXG+HB/NIwjIiMVp8WTxQ166R8cf37P5GWnNptU9rJ19Le
ZuIMnrlmCISFuFg/5aB9RFgfF1b1Yn5qBtVeEmBTf5l6NSew7RLRj++23v4r
wwJS4Jnqv54Ljob5B+ObIQI5hxMp9pYDkB89uU5gw742kexNGU/zcfCxVQcu
gplI8S1nXUzeO3p1KlQ8DDeXCvanbHfr/dnWkdUI5YfJwxEKjl1+nnIXKDe1
g4aT7ZCvukzZFRALwUQgoiLECLvSr+j7deEjAX/27IWmWIJETv1LtE+BzCP7
KLNZd2gAsJLaDAdu2JOMIHb5LaJn3ks5vEA4BSfkEEuglYPr3Ln+N01syGE8
B+kOn1Q7BZ3BuRVeyK7b4PnPL+4IiCjndHP5f/CEwwMdelihGoyeEl5DfjNB
2wPaRYTNLuKuqrKOMFnl+LOQwTmSKeuSOBiiz5QGR7Fwq8FoHaN//pubXHkN
V85OIpd+zjqAQfs74tM8L66CH3bJPe2LqHfZvEq5j+AJQOO03yatKC7NqsoV
X8QJyB7rni7PFBywvqYj5uEdD7BKNj6l5NmYUmgH5jBDvfBA9vOumjLvGpsO
Ouk0Re6OOtSIHKK/EyUSkArqfFt9Rcvdfm0E5bDV5RvvUn274KVx2fMcmfa4
4XhQzwrvTWpYu0UhY7sa8hCw+7raNHfbt+X/HHrNj2zN57lHQQ/L+NFKsfRC
viy8a+JL74XlTe3cAQMce0ZxQq+YypSdbbHynI6b1JdvioF38IQMou+QYSrh
yKyP++1jFEnpojxsm0lyndXNM/48UiC+mQuZsafRvfx4LLRoPfwvqpfNkofK
QXS/IlsPj8EhFxxTofqobWKT5vPeX5sCwapWYhUf66/nrORDs9UX8P89kpV1
xvyCwHy0PVyV0Uj9preGDa3GW9AkzKmjzKPK1C0zwaH/Zdwbu1c32U0RnaeY
cbOxtnqGKomSH4azlH8nyE8zviOX8bfnBV3z1fThgl9WAitNhHtyS2gp06JB
Esbk9GkEuJo6CyXoUZUTMi1sM7xMLaE35wC1jzJLqt3hH253TxATd7NUPaUF
56f0sseRD79RmMN/06u4mIgmhuCOGKIUJNjqIUy7QIMSWzZgT7mwWoXyUgml
vlxq2I+ZEvBQH7OfKZDxjusjj31rwaQCvuPnnblyzT6MuyCccF31HD/GO5Uj
YrjxLJjfo17S0FyBubXEWCaI751YBWEPaBusyVgJczXq4o7Gslpy24Zg/ezw
cPDrCCcY3QQcqVZfBvQ62/TGJcawG8L67yq2NYnTu2GW8O6jcrov7uw3Okit
cI+HvlsodrVuhaxAUk7ixxmqh4gRHnW0OOdGhWnF06mFyfx0XTLfeq2puxl0
GUqWDuah7P3ZbPU+c1zfda3E7KQsWXZ5nmyA3pZridCAnF8PCsDJD0Dc1pDU
HfwI92bqo9eq2X0ItLjN2XGKNZy7rg0x2cKuQR3Rw1LfyFNPF671JMqf82Sn
eShrXB5xKnGZtFmA2RUpxmF5bnP4Y2mClnc6qVgVMcinfVgW0U0NikhgmJa9
VXI8dWH04Vppi/LewYovDTmQFLy7yt8iRlWWHTBrwt1f0gSpsWxgFH4IIk2F
xzCbFI9oV4RVJr3h3htXaVUo2euNUCfeDapHKufK9MDreLufFtsARJBA4Jwi
Qv91EzB8k4mSZ9Eq+vyIvoduFkVuOI5gzLRkmwS4SzpNPA/p+ZCwcT+9MNHM
01lq9GxK6eCB5UAKT1UvQ+gOjTHRP/HafxWDIoor86dNvTuBDYBXkvWlv9Ak
wnuDKHeZffCZuPSkHerl12eI/UP/llwGaZK73zldhdYAV6qemJoww9c0pIhw
Hh9MDBB6ov7cpwA5l0MFOGal7Zdi82wR27iHBVq/jLQrVGmgbocpVLf9ozZc
NJP4K6HSzBI/LPIi2oBquQXqVWrSOP9Wy2lEbiYvHQIzWk4soD8vJHPmyjZk
R+ZpXd/2JOBVCxlHqpxRbsawbHnAsbgo0J1BcFb7WEP7UpcdtO9UCWvl6eo0
zWO1zd8mh4b/8G/4uTD4bf8op2dNtAtIyL7FK0FCrJXU62lDk3ffawC/qk9b
4bkdQgpsk23LAsxKYcQlMUwwklBXZa9sbVbFAxM7jcuBSYYvAyvPdRmbtsMh
Rr5rY8KFzFTdIz0VG0BpMaE9bbs3/K1JEVWHn3RDQ9BdSkLb1XBrYRhVnKo+
yyIysCZHq9FuLUwcaxR+AUCrQsmTX0CC6gAaPljf8J8dSjxJjMREhXtDEtgZ
fKELznd9bfzGAvAlF/iI8z0FKunT75VnU8qt0r/UqYngKxMWyJcwNbM0EyNg
mPbbfIJWAgO5fStNmFzn2jBH/D4UnooD1Pbljzy5T3wjtNL55zp2Gd3Usug7
MCXaPkQq3YSQsYlCm+D25BY6qUHsoSN8qkkwewe05i1VscFs+2M7k5E1XH5e
9zfotBnlyzqC1okBh2r7HWeJLBu+rWMoRBuBfgV78slOB3adMUdTsRyKjGWK
MHZw9YQZHusQoe46zgCa/HvhuIaIMWoxJAf3bxoa5pTLlp2OCh4DpCPB2MRz
thjpeeQBiz1xfbhUwn+hOENe59SQ9jfzhaRsC4js8F5PVX3f+EqrF4ShOfLe
3MCS++9NJdlccyMQKjPYmBPiYwbPc0J9FNxUmyBBkW6ITiBopgnnLY7L4QGi
WzbZREkFiG267KRUWpLrNbqzBtNxtxZ+cqkOQZhbtNPLNrEd8VJPvcXgh3HM
MdZWGu7D7V6FfQC21rPl2MGJtlaJKkN2ezKn9ME7Mgy+k7B+Q3IfybHWJxwI
5ZT9dfV6F2sSP+WDU4SecO3hxqjjWNWEb6VZ4B7d44WGJqgDPTpJRgGfe2pU
dxWMKc+0w0iy2oNU2Sl2cKOoCmjUHAGXZDTzr0X/z4ZeYUKsXg7FzHXilbj6
J4t30Yg9dvI1DF1CLjjQCYJhK4OGf+a2C674Z67snZA7WQGwO2lDkUNllny7
Km4Bf/vfEdMDd+IZzmYhJtIUNDIWCBMSWIZ7zlcekNPpUudO8KUP74e/aGnE
acIkGDME5EW4gk7rgnXk4UdeWEnIfwY5aIkmuBBnthlUvIi6YoTceFlEyVuV
Z8rHe0Q/9+6DlqzLsGkny3rvc9p3h6noxuBPq8o1qEWlvHetvQ9M4AXcoSz1
McfSCIEbUpfiTM1GVzoymasnajRvlYnKp4QYqo1gIQkYjOGnMUwsbx+O59zk
yNywNtKCbeBE0ix3c96sbkZn8QsyJjhWQFIkzfg5zBFXDkapGJkIOJYREAuM
a5BtKwgJeRW7JfwdyXH+b4Vt6k00XxQm9+IDXEMozwjdG45LAgsh4hUI7aVu
sEE5DAblvDr97YX/WyUfUzhqFPMeMrKU7l/29rKhXEH7CPl1rhT/OW7+wfAO
AAcORSG+igxxk29KECEpUZQ3SxUI9reEjSxlXqoePmcNfI3RH+rVfkLXJ19a
l/166znCARPVekAEPeze0loTqt3RcTHu/Okm7EDHzwGTbZbTHKMrFRO1mNJi
XAPnHegsN9kmyzFeICwbI6/nn61Ml+mQTiw9H1dC26QmYibiH87Kgf1UtsRX
rTp8LZcYt1cwtR2zlN8cL3CisB4xhxK+jYjwPCnke3ZDk52E0+gzYFTiNyT9
PtvdafUvFF0CeCq0eGYI2ZRDPYFobwI58i7Yar+ncyIGmdCCHlAVndD7cPwS
EkTXaoHtbnCNTDTJCC+sRQKaksuVuLLb3Im+Au7uin7Ea8lmrnZ34mvHtpqY
4Hg7iXDQTfqJEbdztBRSQ5U0mI+/XgTBtLi+bZ1XhgpBF1yh7vIaPi2Epq3s
gA8iazuUeDAkHALOBeDqoXuD98Qo2tOSkXyx6Hfc3a11TfixQsoZiJoSb7Ne
0RlXmsSMwssw4AQJv7H6d0wU/l5VMpRXZWUeU5PeAbqQ7a5vdqLrz1Y7EASD
i+Mkt9rRaBLcvEz9dpxZp/WVAXNO1+sdI3lOCv48giudczNTvSi0/MPeEtW0
Dy7rq8R20dADl2al8BV1OZWeFmgmCMTUVmDMD9VCPDSwqhI1K/zvPNH4dGbp
LjMJkBqTeqAuj98UmCmjTUS5HoJt/IX3csA4bqW1x9XczVMwYx9cs4uAgrLn
51TiZ4JMw9QCVtuUFDEpq4cs9VsuEQAPE+EGL7w2M4mUFxZxN2VxGD3S/seA
7Z6Q3+tfZn66F+nktawAvjgQeUpqER9x1Dleq6IuUTMpdk0qX0kuNgAFN6z7
wpi49JeRqATB8R8SAZFeygYhfUsexmjseUX5g8VyXySZILkBctDXUQdVabPo
5bcnfCxlwMrdadtZueYF66OqeN2A+MJVORfWPWD/7mO772AMxCovayA0FEZA
qh0WMzqpeUYS12OC4bVanr88vSGIL1eiicrjns8G1ImqdOKx1C8DzQVkp1Ce
uVh0PMp+hmAv8P7xPttAss8DrRi30cOugLA8hIQ78WU+ss1qZ2h90csbmHfQ
figeyRclztcEfOWLALTZWQ8hqpxpXly7Iod3CtwpgQ76eOaQZRQDv31cUGYk
cWLDSeZrJ9d/Fejb9TZ8MSFbehnpqZIskgdgAhm1ervmR6EKw1+D8b9cuhJU
xD5Xr5l8pifcMkSxtYj4VH6pTZjJnUm8R07+DF/vUV+PjZ0d99rtEzS6Jwmv
zoDN6BnjKBfPni75feUJrBWMvyDpCdscryvWrUkQYRiRXndl2/CKBRLuzm4D
ManvRHnD/u6TIOV0pB1GGHPXoz6Sq/SgqAQel3gcLdQEB2e1VuxR3Q9DjWfS
tBH6x9M/HLw52CaZj8FXY+/dotjqSNSZvGNqIOQQn/aM9uy1UqYIyE9NwoPH
go8WEoEJJosWvmV0Ov1VFrIyHhapQuJSXNUZXJXgpYl9fEoN08W51FhI5leL
DM+J18GMpJpPgmJX4k3bdzt9BfXdc1ozJAepK8RzYhMCNofuX+2yMKDMsO9G
HEYCo4wD08rMTvdMYIPl9u6fo8/68BeKRbOn3P3mLs0bEE1p0rZihnXvYaai
y/dQzGrEk8L3dAYyUYP4qFK6XEaRGxG66s9WVYjJPubHacOeeiB41H48gl1e
1ojxwW4joADEjIq7pCF7e5uGYVBufCojjaQljaklEt5ChtOosSwNktt6kUkT
SzIjsV/oTHzteumeUD+KOy7M766VBZL3R1JWcgOiOtjvOhzJSRGdwIWIDcn4
CTh2AuFxuzzpSy2OkFTuGhww8wl2jRnP2ZZwZVC3n2CaDIkqiyzGHF+tUkRy
YG2OoCYt1lhsY2xHt1f1RN0ixm5ZEfKdcx4B8IGb5kmV88pwuoBvIHQhHNWt
WT4lKcgMk+YWjInvn/JXQykoApqUToXOpmAOzsPNQ2SgO6q8+zox5uU71wHj
kpBGsPYafIppgYDPkZe4dOzl3nFcdXY+DrJuGdhWycDR5stx8BLbHvxEWRTQ
adAktKnTB/Db26E2u7IxoHWpx7Q1fwet2WWBKx8M3osBv/70KoXxNrsTi+Ee
0/wbkqySs7uH3V3jqMM0v9gy1XHw0LMN4r5g0hD0t7PjFmbmN9odIPtR6oIm
+EmhdOexywX8Iv/IP592mDULh6L8EpIik/zFgJlQpeEan2BJr71TPeeb8a9U
f2AOHqJi5n50IOzTkgRPYlDZDcWSQVZLVJCqisNuUHmvUlS7Pa/xxXroaIaf
xka3LdtXeyeYipGpQZsmS1Gc7WItpKIUIOpKa6xJWi8lE3rV0qpekqMeCX41
EK00wjVIPGaFEzoHvewrl3xGCviRTkn+ugEU3HCgpYFiLEyHrDpP1icQ33fI
2NAJKr92eyEo5HtAEpVrvDP2kBFDCysHEKp93Wev0149Gd3aI3kIkwFmcYiE
1/nNhSeOo3k04Ij3IbxV/JsgbkTWxWamaoH+gerQWjNs4Mz3IIz+Bv2rJOSN
JJSr0fENjX72sz5JeHemcL6Mmw6Ucrcw/PCWGFro2ja8RbnS9emWuYTkfLMr
6ryesZAOY8BviyQugXNCtysssuNQfJCFXumnBChnZCsOf4BEfH36txSum2pJ
OStiJDE2cy9cMtaiN6ndLOuEbFUADG/W1E/P1evAO3TUMaJI85/RVSujmRJ4
MGKmtt5xSf6yoyCg9Ufzx0DlSxcSpwW3MQlmOj94Jvf+bOmtKuryYKIiVDXA
a9mlzPwux7UcwOVWQuOvBAgHcXtdi0nezWTBp5pcC69cOY8MnadJj78BhEO4
EFO3Qa1PF1iAr0eOyTfqtNJsddSjTIRjp6zff6JodbGs3PapSuqVq6VrzuNY
Pr5AZKuoNNzv0pS3I6SFHmDEx/aY+tmWLntDHKtg2CHcqxAXz8w30ZDlDu1X
xj3O0EOUG8dV5qYutSwJyX5oGE5yOvjQ4nrDXkict91CDK7pAuUSAgRXZN2j
vN/KsuhlP5MP2j8wc31MxIMnYnXMwYSR6m3QweKLnpSb6j9IdrvSRhyK9Zsg
K9I6gTOhFEMswmVXkLQnnH/OIBMN32SLB15hoBzGQ5pfJMdTCCuXq9l1+yLA
MXI6SvFD4uTFV/tQGdwaLvz/aI/ua+LxsaG+4z7O3Vsgk2/7Hqcb5YXU7CLH
qBMuSQw+2pvhmk8Z6yZX7PN3LGkNZMw0YxcZIxMAleNU2tpub/3rcGxAPWk9
9p88QOrfJdoFolwwzlhxC6JaOtGhshLAkXZIjnCHpj79JHlndIYpZct5FCKa
finhzqdMFOhrqUnvNDXmz50BdvXPJKwBeDtfVVYYsF150N2ZnohmIYK4LBFC
vo+xKlCUBj0PawlWEvnBk86lkQuLOoWwMtIooHAng7M8bFHYbmHfHuOpkbrp
9IqVuqpV5JSm462z/F7JKPHhhmcQFdAmytsK7a0xJzHMC+BfMDcCbiS1zlLP
brMeWuy3TUzXBmBX8/pRDtNWMZdx36Z43Jn8hCIm2uInDNPQMv5dpy4FuFmI
6BoKCtqJmx3gQnjFu7wi4ZNeOn0UmYGP3cFvGMHl047vW9/wlg018GN+ZH/p
UxgM631TUTOiwfpiTIPyFRsr71GgitIxyQ6+in0Iu8QaOliyzfhN8eEiauXa
TrqUBcrMfNGOZYaK3VbmKkswW8z3Us0ZJ4RnlAjwc6FYZz+mldYrbTmFZzSk
5o4cTruhb59MkxXKKPg8JMHmrsZF2so1NohqZt6d2wEwBQGLulFNtAHg2Vi9
JiscXdETOPEhSHAqPlQmCGaU3ymMcERZql4fKc+rtG8MIyIb/vejF2QinU58
VzUQ9czFL5BearfnRkVEupKFxOdv58C06IAlXl8PfHghvrB3GDyS8z6S2BVs
8oNyhIq3ubO2lVfABX2CGRNXdLAQfJ8afoUJFs9mMHodY+kUN9zQ6W45ydMQ
FqBO/OVUw8aBwWNt275Ry6mkGewZKRpfBsUh6FuhI1zHF5Ut4eaCSg2UICkI
mT2hU9V8LZEJVTojnW+DOK0utG5yF5A4BON+MyOvam0k3UImAaoh6DaHZSRL
wjZXnYxmL+Bunq1I97nwVR/9U+JjWUvFS9gNPxQbMZJaOYoVlFDrETnUx2Ai
xlEY+zQ1wKRc2iInxpSLgImTbnG8HtbG5HW+munJImVCyuVujA2N9iXcEaDt
Ulx51hMehSV8daaT/dxUi6JGeyEkDyvzdiIWQ6OmyX7F75Xz263tW81r4bLY
Vtndmw0PmRdomU7nJs2UT8ZsehZNBTaIBzAUJZsd4gIk5QQxvZ/WoeozD4SF
8NTyMVSbE5Q1go/qHk8Bmk7cLg8xoCUuAP0oXptAwN3C781qFKEhXt/I3g9E
e1TgCp5ARiG5gaTvxRpNF16lPv/T0UPqjgShkZElIJVfNGWyqI02DNKSzrEv
jeidAgpys9QyaP/Jc6VK+kGq0bUJNdAevaj3iijaSZnL53qIytQrmRPE++9Y
hKALFIfhktt5XSK7GXwsdrDMHxa8UMvtvOQejddzv09vx4PKlddHMVc+t0CI
SH1STv8bBKplh5N+4ueNnH4BCm4nLgRC1XfxEbCPVPx3fG3kcewtnjXM+Ev2
lmIbOePwsZ4g3MdVuIgfgHi+7NwE9+nfujkcguQdDKOJDht6u6IR9zmM8Yqt
vGCXcoRw6jmP+kWWeSE88gESME9ainhvTB3K95Y/wZEEOD/X+htgBnv26OXP
FhJotHyx0OEvelOMbZhly85/khvbmSUfDEu8/Zh1ow2Yd3U/TgfYMN0huOQp
bVW3sAOCTbePymzZw9YIDMpNasXPHdgPyntaC92i9ET52UI3sdFuoA9mVmA9
7sMkANSxWuKArjZ/WvjXlHBFFzhYRs8irUkVZVpt2CNoWHiQOcjp0VePESd4
w26+EBTY0Q4MOY1vjCYHT6DvC4k4aK0zcno60zcsO3gUKeR3CObksn6Epctj
zQTnwbXrfuLkO9LCujXhs1BukXs7X8BjQLhBe4AAexlS151bmRNoxKEvCsq/
vhN9NKqQNuYFNTYVBgTB8y2/dEIFws5yrxBEe2dO0J8m5crB1VrGQ89KePEB
IboSsKV3mGOEfV0iiVp+7AeuzjDhwb5e3u49CYkXZJQmzPiltKE1A/8vLJ2t
zCJai6lTRhIXMgOFknzI1EsLEtnRl8jDLqGzHH1iZ6yzr/qCngindJkkPG19
wcjA4GaQ9puyKntG6D49wCIA7lxs0Gy+ly9kUWA+uB+0v5l5cTatp2GQ6b6j
du+GK6639I6ETNKT/FQxyj2PERZC/YOS98H/yGabUe28JLMQFnkVkAHxnNsb
zypaesm58pv89Kam4tvjIim1HqCscj0cJLMGIeWsRs1goJZ8t6ppMfDcYprQ
GpjO3gk9dfLnl0cgUr9w2pFV9Lnmab+0Q46SmB3xKHASQSmF05t4OjCHKFU5
uNd5gYO6g+U/rRgOR9J8SgBCA2g4GBSDgfClRaN9eWV/4ae4Vd6vK6x07r2l
mj/PTZimkA+Cwuz8qB8uw1vb7c1EwCjMMRXr1b7YO33HZ1cRovDUkAhlxRr6
lmJunwUejVR9m4jZpZh1JFXY0Wb+FdpB8oERGzZRiGe8EOOacqFQ0umAT/SH
/C5vsaIQxbXuCpRnqqj0GdazelwVRNdGmoofz9sW4zgcuci0ly5lBtAjdVU9
LDJq3dKSMwPwz+t0Hb35Kx8SVvfe6oJykwGHNsB+gDSxy15opD4ZY5hc7KyA
cnWC71lipUral6++1re90ulRKccumL+o8HB+It+MdHUUMFvtu4lwK54eGN2i
WDCTa1xkocAd/2LlB0EPhz7d3E89NJPxNBhVHJJSAoeDlZd3KcpA8Dm7uHMA
jdLE7Bxqtxawy38W0xy83UvYh1I0lesH+fETdZQJ7HFG0XvgyX3KQpyyS2DF
JpaW05XsEByQq9APG8YJGsz3DnAjbPQxPLPhOH5WEgD8d7BPowRSJ6VeaR96
WwU+Y1jmdKtm39QBwXcA7NG8C+1NV3NEe1Xm0BZkrSEQBHUhVOtVHb0nqt6u
mlF/ckGEVZptIQYoEF9RwJg6eU+et4Zj9uh6XPQVAwAR5bmNpQzlGzfL7kcC
f4kkhUqd7UKI3WjayYb2LsK5b72ivI+X4/GkgRxRWNA+kvSKLJ9QMI/Wtsm7
MFAoYG49/N5Gr+FUlnpx8Pr+6GSGnSWztxZLIyqN4m7CVf0EkGIvKReXvH7B
b5D0jlrepvehdUADqeH0AmJfiScbx/lRgQwfEGpdwlPsj9FlPcIBMqZHShs4
gQPkC3Mxz30HkJxIFwBpcjG5UlFpKYBsByqVfnADb5LhBDoKCwjhoiA68WY9
EobkCIHhbb1MF9WtZi0Bm3JER8udVWpp5nJRBTrEg0YCgl11Ri63epzIh947
/ND8riJ5EM69Br9jq3r5PvGe8/5lYh4DRErcHUuegoBkXZWiq1TTBYN37Vqn
BdspdxFYsNq+r97etdCTJaMBCGHyPSQEPxJdBZkb/st6/O2t6hnZ2aIwab+M
HXm1nYOqRXboKHkXU8WfT61bRW2a5o3A+4mzpenY/K9YKe/o+ButFaqeXybg
VfANqM2yX/AxZh2LkhCUCMqFFeWlVZtch5F8qeawZf3Tf5pM5OMtOoU0B15W
CthV6UJDoaMNsNolMIxVdQvAslWpPXFFC72PnipPuZVm9U3Xpcekh1OxjFQt
bEcPvorz1ErLaipGBrpmv0MmlQtZy2qqhYsyUetrCNlsMdgLNf6NczY4zXmI
9UGPXv/Icegk3u89DUgdnYgS1iXWi/huXkG571vsR43TMH1IKHZyK+Pl5Q7E
SvZUn9Th+NG3VDTVrQThLkj4Z0OpNBZCBu2D4jPFevwVQwxJJV8HB7VyUf+W
VvuJ6gvEsOhbXTmYQ/zdnzmjorE4l6cMZcrcrRA4uFRGYQ4QmkzrV90/Dv2L
G4zZ0ibNxapLGZWF0js+xvrl0ywlqwDulje3gLk5aOqOT3jj7dj8j2IEvKlW
/5QJQ+oDKjTOGeSYmXummdSa6XVCnrkqflt3+XSvqvMCXC0x+AyOK2f9Gakg
sP6g77k1/UoQF+jJ2uncJKwmc2dgsSxBDxBzoqXhVtM5zC6uGU1m4M4EqDuN
eEpf1RdgIm4BMYUxQH46+CKyhIIKlPuL9V6VVLp+1SXhGdpUMh3q77TSyD1H
kK6S/whGfKrmvRBni+7mnk1qb6uLkOkOp6+DmZYIvtcTN+rALGS2o2YOZS9l
L7lTY+S7p6nQ2BoBsh3ZQkr1Y70JcMkFOEyrxs7644IWpaTWoGy3AjQxuRaO
u6IlJpZ8dt6Br0BDIj1GcS9GGqtm3q1H/0fmVWdROZKn9F2i0BYg5J7HV3g3
YKzX5W4Kf9lMBC4dFefnT8VHYcya4EgtyG/2YDFBMbLsut5BIYx65VPhbgcf
ceqY9KxqWUgypcGIN0axNnFgUetFKjd1Urb+NJXC6xtTGsWXrifynBwqR/MA
6AZhxfzLjWyKjneogVLVzkZuUb6WPuIp6bobQ3XU8eOuXTNcaOyMG+imPu5e
cSkMEI54eCNNSHU8bPcQmdTK8dkCdPf5+FPc1rWh2+Dh2pVukS8Nj+vv/aTj
vMNdFRpM5oXlHmdl1zdbILxM0pbZ95SlutfhrbctO4K1woT/CBpEslFBlJRU
jPQD0W9ExZRFuhrBHNh4MsdJ7qUr98x/oQmiMAF/8eAa6I/9phkjRhGi8vU8
90lPy1tgOU7YIAiexW7AS5O+Y1rWm15pz+svf+ZBBcG5DsHfpo93QUHaBhU2
cso8WNW55KquONx9/XeOQjBIhqyS1L80E0WyGcD01bM4nSyZTDpHLwX0eYUS
FGnpJrH+AcAMe6BpnssND6TxqQkzW+vScCZ0YdhNYv8fGzLTpkmRoeTCVttg
IGNlk8wcGFXc8Ahw2ZJChsPhuNSYhamFAwWhah7jck3tHI/zig17wP7ukKzG
DiluU7edDy+lhzp/5CLgOIy0tm178gQUkFZnkjcgRQQJQEO83f48Gsv83uDO
hoCVoM4vgoZu5oTntbFrXUAuhsR3q2sRtY4yE3NgeTWghe5ItwHkb27xpE8P
vmsYs9sJL+NDSwNEarGJTNPgI05kgOyxtlxeVz6REYYfUr1n+p52HSVvguJs
R1N+la4BfSueexgy1nwkTpGOoTaMyhnKnEGGgFn7p3KPDzgN9rJDT2tpq48E
vGG/N9WMvkBbkR2THAwEDYoAyTDAEqeWD6+xJ6a0DIwUDYeOfunZkFlgHcXL
ULlGjHv3+wqgAU07ESUQvygl9WU4ywEjRyoNc82ejOq7myZAeTQ8AK61wu1R
QBO15expY9jdF88DQ2ufqZMqB0H679B6UQEFm91rPgCmKoVFVtLDGjJS7Y16
ScwTG4WDQ05R7hQ/oXqLtMABuoRC7GBIRUdp0lC1nTZKie25FevBdlopelks
KV8mbxYApIAdQ+PmvzAswVDHBfJIIJNiXxgRkZpU89irGvwIBw8b2Aef5CxV
n/1r0fMTknBUCh3vzDOIX4gKXJKT5t+/1ayC5qjeF20HPq4HE8UrsN7u0KGM
Lu1SiOZY4dS1HqU/HeP8r9JF1dW67mTavaHc30t+BzJkXIU32IkEaN+suAC0
bD3IfjpYQfWflQ7HN7xXL9yBPqdH8Gpv2O85uq5s+7FWh4TmdzzHdRe80FIW
JQDykJMlOImdR+Z6i2rqR7Om+yVpv3WNk2ytG9LQIpqtuOlNq/W0ZGLS6JZ8
qsQwj/i4vmrggug4YrwJ+RCMCzTYyjKLCIkHcI4Nf/r282WgikJYHJ5GUiSy
AoTYecILbooZailguWxfydnSgVYQNw9LBj103hQ0QIRL7CT7K+UfPk5aPbwL
R/9q+7Fv918RT+drjcw1OWiu8jdlfbWJp53Aj52HEkhbp3cQu6EyvBvZ3CWH
imSirEClAB6LnELPeVxQwlphbgo4A0ZpYxYTdbPDocyibd5d4kuNNQYxuVi/
xkKRLBZOhxkORbjuJhtlvMkMtoLjwsv3fJ5TMhGodgjrZ18Au2v8R7MH9sWj
0ckBXdtyd6N/Eghby+9ZBk/EEaS9iirHeeuqExhV72pgPwvZ2r2lfDvSqGBL
2TW3Yclkkk1/X0kH0Bz0s8w7EX7olDv15qxaxqDzZrhzygC+rqW3PM++dDbB
HbEn+OS2QZPzw4fAvzc0yL/dhvx2Gs4FDaJf/VjVvqcSQP6j9iwZb5fXjwbk
BEEAoBWZHp0y+PoGmTW2pR4KhYRxba9XDqGkJ9V1gJLvjHpN4Kuzm9drQUsj
OJUg2Jv1kzEftcwrUdT4xD5d8oR/HBfX3wYWAjqaDLnLq8let+gYXmQwwcF4
Nb8DEt7/LD2152FDbLlqh67Ce0pQhJf5CZmxalypXDf0nNi5iw2RAX+FsHeh
pDSeaCKyu8F/en90IEbZzj7N0nRwhVVCrvxb6PsXFgSVLUglsgHJrTFn3xRk
HbfZ0IZbRbJrRbZQgvB+mIrx0zcpQYkOsMsbfOJ/Fz3w4S/Y8qaBb6jjSryx
dt83wm6l9kQ4wBH80SL+7ePFHrB+YAmMtmcZqV8UZGmfqCOr7U2qB/XiPxj2
G48sPCIXILr/12gr3PIui2D3fh2tSLLxrFmXeVd1/+A/cQt1eK2WDxyse3ao
xXIebZCeiLzD5ELsaArRYPOZvSCrZp+Fks98k0aaWvKGuW5qJ4pT4jByRZeN
Vdmtc57g+yw6FwaqIyI+TMAvBiNYryYYDrY2iXgEKNeu/GttdBuQuFxtAWXQ
faezuqUGgbQSDYPOvWcl74pKcbABNQs+HLyJMGmas4FoyxVBvmsTs8h0I0fJ
Br9bUdHt97XWBNB13T9I4IxfKfVJzGQVV5L5ySLF85athcdJVLOHKI9JssYK
PczKiqrSXhrIjAfp+sdQkCLNFI5ixTH7iTsul8ggKC92eGp6TUQ8zBvWCPCx
2PWyZmu+VEkwol7iHaUKthebjZT5juoAkz95IQiPM+lka31izkLfI2K+MeVB
ZGyM8QCDNBAQK9IOBnsPgxxA8yIfoFaNzkhbft6UUM4YsrBZkFe9o7Pybenc
sTXC8nss0SwEhTy//8exsQ9rWPq1ravfWC+nt5+BOmoLhQCiBsa+o1bExRUq
CRJJr0HDB9sQZIbFhIg1g9pJMjhEZ1P9yez/Nh+tyBe6wHAU6+MrzDVvGDvU
N4Goz39gkP2yHQcAesvHBxCeBJiT4qdhuqRPV/IeKCirdzjvFYA3cdTntF2s
n8QlOpN2gs8FzA3F/4YuchGbcWb2Lm8QqpCdfY+jFxjyOr+98m3f+cPt3cIC
L5kGeViA4zGoSieqDwPr3SoSlE8vY3npXsTkFwQgSyuoaNjalyLMsOz7SiUJ
dF1djbgNPPvlbu3xwA8yYy9I0BcbVYNoTv10DpNRyi0ESKOsdgdir8Zdnd7h
0Zvh+gt4PFJFRW2gkcUV8woOyHLmSTYNHc5gHC0mAzEDqPkbKQ0AS/6SznQT
xgWH4MsQhCQsrznuvBnRbaGkYmsYq75NAl59BE31aW+JFikOztp53Awqw2Vw
l/eUZREH0uC/EtEbvsekJCi7kpjV3Tf//AvdIa+jg+lpZ3iq7riyb7jK+T2H
0K5r+eVRzWWw/BIE6v1BmGeCFitiBE/bkYhP2Eo6rJsLD0svlBQ0nOxn59nJ
6grg+f9QqfVBHI2sewpHzRZgUUAaPzpg6hS/EjA37PuDlCfjJdqIgmmFBLmG
RETcpkzpeJRuTRAXb9t7Fcu/YjLyLAsO80uHDrL7BFg+tpnafhA3uknTID8U
DPghgz81CB3t+WQ6xeozAVwg8WV593u+KXfMOnySsML5wbZevBbtcxFPLf6l
omhFC2HQFGzT06X/sUL9DNfZkx0QOUEaK7obmTM9LqTGrOA0vSLjPRvzVApi
D8AuXyaVRjUi65XBw76/5rFdwuRVxx/2pXi1sI3QgtjufVzq4DZs16xOfyxr
sk+2f28a0sepMEQ8cYhEV4pkiAD8WPxYct4koYQ9mTA18Vs3exjZzIolwqWR
8m9N7XJnDV9R0MhVsy7QS17PEXxlmlQQ8kIFHkmM0wWU6YwRtr0YYFfxw13F
Mr+M5oKkFzCcGPOQrU2d3Kb6UXVoqlXGC6YJWHe15YWhN4JoSzGFakNcbzz1
X5bX0QyPNWRuSLht80qdKz5LCup5EHOgXDDCyaD1jnDwCKO8fFZk+zIeGeLV
2zqpVvOLL2xxAi1TtW5u4mtd74lbAhx9JaFAS3znw/LST1YMzp/YyK1m6RIp
56Q31mZiF8k8Iu6zcTfmOJVkSeg6ZEHgA4vlUk3qodvwZ8USMZMJGYS37V/I
1OVO69s65b4Dxr7rOIJW5QdgXE0bbG2Elkz2ikxwC7ZoSAPHYHQ/7F3BAJjx
rlIFB84KwA96Wzr81H0YGpcwCoJSkyKw9uuKQz0AP2Zi7hVIEltsvrhABTIW
PQjwvgGCHHtF2TCLVj6vYmA9UT5QY/N9Un7+wFrItgq32ZzU7Fm5HLkJtM6T
HM29EF5s+cx/1/X73WCBBuAFGSktO/gn2adppNaTBHx5wAs/hQ3xJiPBmRHN
0BTAs3+FaReEZso27nQf4K7tvhYBYr1hmxbgMkR+fnM5bYX9tpFLTyG+BrZl
bsGmovIFEZby05EPr9VLsDS0/CRQaC/B3zcdcOIWdF1QXa+9AnLnNXfNKVDd
qu5Dhk5TL5Ai9wdLIYKWCH6oDgveGtIyY+9y1YBFHj+W6lKv4+XH3AmmOC9Z
OeQpcxu9UW3+L+5t3VtlQq0Z36xNeeFJ45LcaoHHAaIP35DHfU3/wP8pRIgk
Zxecx5cr+FCgOJ0iP1mqI/dMAQVoiF7idqQGjDfDANhj26/MZIdl7Nx8H8tE
DexFh0N4nSXh/2XtbFevp9IBzkYfLQFaISZV45yysQx0QZIWdj1L4Nn6HYoa
ADTgrRhA2N4BbzBNZrRdSMMp9XVAk9VKn4LwM7Txi3ENT5LTo4VFPY3KfEzP
Zflb5IhO1xVoYKI7zaTEAjxhh+gaQoaeT77no3JnHQynmpv/Ie+HNOp0Aw/r
CkmgIBq14g2H5bXBRjtNsI3HCjXhC8n9p2wNCGs4v1HhmU91BKgSiFEkG0o0
+WM2M43GQzS3KnLeE0QpDIIU8PoRfTGuF/yruWCAlfcbPAbq4Sqrxgdeiztg
gI+yFWhFgM92YIvJKtCk49BotYumGZcsp0Dg1ricJ7M9QnLTI8GxjPQGDFWQ
CR42Rjc/4ktospEumlnOhSho20URZKioFa8BxDDlZJKdLMMGNDPLTnNu1k2H
ufPBE7QH9pPNe6CfuYveJ+i21cH3y4+yht3KhGVLK33vChhB7jcc/QGBEQSX
+BIv/PfLQm6ndFm8flVQgK8A6tb+bFFBNS9ACo9jPT9XQNShL+5ByLzHubpF
SJ0sHpu+Qn9MDH3XTv5tN4RV+++zO3VouUBDcGeMt8UwFmXXHRyqMBApArD1
IpGZrppfBr+nS+QNLPSUw0oqg8vKw8US/XtRm8P4U9hN1Wh0EzfvkxBYTd6H
PTzRW9+r904Vt7Yxi+i69qw0PUqn/Hg1x/fWUXOod4vBqXZGYPptNmaES55O
MBqcl4OXt1gvAtRLwokTEqzdvqIKoAjdYJrz0QMn11XjXMj15RD7pQNcy0r/
RynwgUpJiwtj8WXrhe1evXWtoU57wq4AOn6klUgtP2vpeXK7mMRbii8gsI1/
TIj/stqBN1ba3/AFKf11KTNja8wMuU+DARwl1BieIoEokOvrAcCqwZAW3/bK
3O1Im0EXRPYkY86yxe1fc43vOmJNiXr61jeaK5YazFN2ewVt/BzPUIdy/P4t
h0624/JLo2QLmnW9dv5U/ca+OF6vL/7zX4GRnzyLBIjZ18LwI1QcpmFEix6v
jZHibYZBpiImdAmFe1fpBvcuecswX/IhCeaTFcDWxs8iO+nFYT2tIl3TKQXC
6GNUowpzU6L4UbIc2ELyN7CC9NB8ZpDUT7dWu4mcPTH/d2BrmX1Tb+f4jPdX
nERZdS67jlvZf8RiNxwXblNSC9YpjJfG5JdN9TThlFtyI2zQap/KQTMkNrWF
MX2VYVWI7r8XJexlhE+MEJbJxly6D497U8GmNFRLJ+v8VFZnlcxDyS2Z346a
NqkMHUy3PF/4XXG3awMHfR5uOPL/Dmu8NhRafN/El+SR7J4D6bycnl0uyDex
0gyfAA0QO+qd2EkBE9pig1UBd/c6GsNNrS22LaUuZLEtUA6x+8bwLj+VHJvT
tv74VuQTWTe0JOCW14YXeLLwgrFx7oIhnLHzcqbV+bnrnmYO3Pqf7Zv2W/S0
6F8qIpzeWeXcX+6vxkPYJSyVV57RR6wqVGL6X8G2pB2lkGqj+PZULaNsNMr6
r43HkNKKQVvP0XO5kTTz2mPxl3Qc3updSS2U8GMqv7ImwrognrseioPASA8W
PhBl9wLqABxYD9UtwYOR/S9x5nNeSWm14MZa1Yp+VZvGCmR27o1oTTeB49gn
Q1vN375lEHScGBNZ3bfK9K4RMWIHruvy9/GuTWO9hrvQ3GBPauSc++C7XHkm
ull6urH/Qwu7qkHWOeClbteTNIoNdDMFBJKzgk0cKSCZGifg5GR6JCZmSPvH
Kxa5DXht4jNkGwCLxLhHxEA7IB42aP3e7IIUWDFzIivzNF9ajtcnLGciHv1U
Pf2CoflDyrK73YnleTvFl1iVmZwoP/90HcXZjs96q8vaaOYkk80GHvuANYBN
NrDPHT+ku6L+WXima13V9+yJxxnmSDDN/CfBBaaHZdFrU91ca/P4PetJgXf7
2FWU91jz+N9rnxYJVjup8KRUCgqyuElG1ToDXUUKnVJ20eXpMd1M1ct3pmEJ
ndnE6rnR/4Ew+LTQNk0SR2EB34MFjD0/ARGhF2edeKqZgYib/8AiarJbzapl
pCTOEOjq39j4jSeiZwfn2wQVtatp3S5LYgQszvQn7OFNFqM0POj1zCp73umw
4Uks1X2b0pn1xzOmnpNNl/XAB1xtcKO5VvnKW4e6EExr1hF2oG7XHxKQLbCH
L3jAm37OJIcNTJDPbO9QdbQaB9YqYsjnzdmItzwEcfmv6QETAJkb0L/6mptO
CXV1JDQkTtUUFgLBz9zAe/hxhXNEdV3wshvkO0W8G57I2YCuNu7hzJ64hklJ
PtLpbK1TiO7uslACvVTfjI4g0vOs++Yvlh3KL7Q82zOJ80z5qAVb31M/8ovi
9fzX8dHyIT1c06uqR3UlTPWvO16JL1UseLYCce1l9DiAJ4JmxsH6mOPVBpPP
XQaoXLx5y6ZV66bW/7+NXIiiXpABc6BB943u7r4hLBAqscQL9ldszWegboDQ
TlQ1qUxtXaV7vEMGR2cKjcEKTN6WRPfvoyzVIePNM4RDoUnVJNi5RU4l3bar
ssROlLD6EaK+KGcOH5nwJpkd6ktYs3H0goINl2opNwNKMVRAq78QypbXRwJn
Swrk2AcS/bcNwiN6PL96ng8mu2rWFQRrulvYoZ+U+1ozM53tknqioIg8JN8c
mCaSYHS4IagNdwSuvJ0G8Jujiw0Ni6YbjPqIU/OsLSE/Lz7nrKtuSDsr+4K2
DIUksUOSKXFe9jM2vWoUY6JhEgaxfMn258z+PDrfWo2HEYUwbq/PjGNl2kgx
Mwq21wMJdOnGnzW97ABGPcVwphUBzc/PU1TA1bbSpcGCkI72XVVth+bqoPqX
t5Nfs/A2flpJFCdXwrVl46ojwzlBMpv8EnoXeMkevxCyjdRk1zHO+kBq0750
ICiUqp4H7jlG/2hwPqh8+YIttwRhPY9NCFtpeTh+dgUoRc3sjnZr4vHReqGc
U7ymdsu/iv4Mu1nm7FW5cVvvEumg9d4Y3xqfZAFFkOLNalSCp5uNga+AIojI
+tATzFHeM4klT17X+7wZceDysSZ/lwYfNGpM2PolJJwYINRaHhjpbq1uPjTX
vXJ2Eu1qr41BuTHRmwI7krNa2LidoHm1wgJCVvfuos/6uhnoARp0K4o8x5pW
NClpxGP1VXlGbe1NF7MXFjwuTEclX+r3azQkVxDesdcDLH/aprkUV/sFBkTd
HH0WyCjyiDme3CYek2XBuHk0H8WtDegRNgwlQVzepFhd4O8Q/1ZRZ/jvqVlA
GlOYIZsg8vaIAidfz851rDTWnYMfV4mid6Xaa0lI5UfP3gBENUk5aeu0IxHB
MjX8sdV4dkpRa8MxyK8R6NpgnhynDQHi4kglCoyPwbsLiWNFzMc6zkdxx+Qw
LSeJb3cNiXGGolBB3g9LXySNdO4hBg6cEdL8ktWSKUbS8DeKtZOspJhpfnSO
vpQLXP2SdVubi7mwkQdKtMLhcnSMqnvRVbbC0AjVPM1x2cyZWOyE4AqgwzWQ
YqfHYjak4yOKZ8KnnXtUoMtoGRKyWvC55VELtz6ClY9Jd0NQJTbGkvY9Tn6s
8MNDZ/SnLlG7yBnPZ/WqcRnziWsDXTanlDCmBSFRp878tfwRd23uhC3VxiVh
tcLmG9vqASpXG01JxbffJvGx9kKCkEycVottYriIDoHgS73h7XVd1S0ufQFF
uJIBvfkmupKtThW/Kkbu9Sv1EKhCpiZv8cG+tb1VKK99caJTfOwkcKtdXxBY
3IDa/6AM4bujYyFC764i9pOoRTFy90hQLeAZV2iD3POFctN6VCTUWifOvdYt
ScCiijfK3zn+F8ZiPg/5Ua7RIrpGEIvomV4C0GiPoZX9OH2M/0HEAnJavMV2
hOOE+rVhO7awFe6skkpof2dcLptxF4IeOnB1kzvN+kuDMFou3dgrMoo0ci84
EbumI2lUbf2zHN9R5bzV8cKOfuhvmANBFrTDErGnutXHe0GNwJ1TkKMaLAOg
wOMdLNTxNmV7L0NiS4m/q/V3ORV/jD3KneCDDLFGeuW74pmwda8zXi3A44Wg
+18B/GTkI87iXpXBGg4botkV5qc0DcSk2nMNZGaFlCD6pPymQKDjyvttXgGj
9Yiof8FepSNaN+ODKP+3DvbKasX6UjNaI80NURXaJ2mDnYr9GOeQeaXF4ivI
QTobK/xImdicMyjWav6zj2QfReL90wQFbnK68Gw/H46UcRSChv0qv57BMEPZ
3ayFH7PhpBDJumLg0Zxy9JgaZXXqOXz5rrfjOvaY3c9TPrFrROd4pXCrBQF2
90/w/F+q7uu5Jd1FKDltSHtO7zGcuLeM4PCgQoWDiZLyzJSky4iTF0sOMSFL
AWosYsLVsqcKdI0cpGehOBzs49KalqGAluAgTUrQiUVe2yiq0sSwJDt++OL7
9fMF5sE6zlhbaA0JnOhGaYrMrjObB+yIBM8RICFHZwqzxNi2jVrwVI1SLvm4
FOOju1Obw+ii2CL80asJQHCmG5NZaiOK8xpvgx7uesAOBj1vB+okEBy2f9A8
BSA2hgKXz7M4NYU6LgEx7HUbNUWXTG741lncrpEXzf0Z6CrFFgOqOMB6HTjo
qNTzgdO3HTeU8puuE/KjmIML30XwGRFmItHA5Fp8mVhoAN8mGrSyCu0zv2OF
h3IKHPsAU1t/0nUlXThQDIUS+e/n0gNPDHoWv95cPbCAX8XU5MGP+PVUx13y
b8IyT4w8LoFZCFEokYTxgfC1Upc4B58M3IvbLHxUM5+hYFNewGFTU4G1zscn
qZYE6dyEGJv4zZZTeW2wr5TafCyQyJBOelLi6WHwY2kjcSzHSiZAG7HjrlXE
h6a1TlriCXobr7bIFR8YOR2NcrXN/SzsKFf+YBgA0hqwISPi+qgRV9wZxO+D
vELiupOb8iFqxi9HCoNAGjCJk179guhMGm1i85rv9N6FKRVqBDft45Z/+wxP
i6k2Qrmps/VokToeDNPD/WqfsUSz9mv2owwdnwAMn9CDLyAvJFTfZgWcO8d6
/7/ntfNB5xC7u0qST78dMJXQwmWpLvTz8XInyWwbqd2n4f4gwoLCTHksG5SC
P4KdrQBfDdu17Vtr2sfKI6BESB2ls63qjBa38EvfQ0XkrOWBmAk6vy1RHZmK
W18VO9oBmXruEO4SdGCCc+gyPsifDtk9lXMfVLbGBgqDxFGs3i39X8oeAYtg
HjncEBYP4oo0LunxOanLq+KxaIzT/k+iI05yJgqhAHY3Z/Pwp9ic+v94B9wP
rxP8ufks9VSzNgOTkcd9lysSJzebgWYIxAyCEA5GXbDR83ECVJm06r5jzW9o
kO1iS68c4GJrAS6e9RImsRF3rdx/8RZ/yG+qRYXe1q48ZMxbTlpPSA3nS6ub
usCAmTynJfKsC0U56W6Zgk5ZH8neY405V+ow5DVFZjiyzTWWEYTrOSoYxD1z
MbBGNfIyMxGzkqdc/UPS4v60jzg+BnA7IIu1xDz45TVpCitDPa6CpOgvodBH
dci0TDoqAG7/k5tTnEbc6oq8C/GwAHdlfbJp80pwpDk7aMXTubO4hGH7NUQq
azY3j7yblyMeLw6R2TwFdTS5QYW+G+9WihpiJ3cL/1nNU0Q9mG3VGHAZ13dz
nxJuuin1FLDYNfQJ6Y6duxW80eolptYA5Q9mtQ+zEFdPMxJv2AnHi1R907RB
x1sn81QBeCRhkaF/z9k+gDLgdQHt/bUfw3obTFne9UBjNLowbgqdokYgi0RN
svp2GKgHul75CIHZzvWXsm2JULxs+AjXYf4CXkWlFunsXjVxN6IZ/FFrC80R
vCnr6YYOcl1grsS49a0fbvHKlflXtVfxmUDawVa521WEI+kWKtn6lRb2YHoG
c5J/LWzKQpPMyQDyB25LO5vvzI7/RSLX4CVBUGllXPyqmScJkvBJb2sfxg+U
hQh2GyvQVnLY85soGC9rAsukEtZz6cvK9qalcHqxp9stvrqmZboDkJHMlESu
CcZM56P1lVVChpDUdkSvBnSJ/DiOssxysCqHpFKWT6xm5ySKGlzPwQzfLjcQ
5iJEHfHpyN91PpppDxPS3KulEx0XQf/OMJxAUy/Q2BRAd0qr9my2Fn6mEbm5
oCdSNNfAYaqhkoBETrpeffPjes6K5Qrq/tvAmvfrJk4qTqgZUNeroChCOjQM
4qNHdnet82vmZ9himn7CEGveXytEFEuazYB3O7iqQdBDDhbg6Xpdc7sANstf
ckC7wcTWR/wSOJBJT5+uCvHgfVbB07SBRvHpPqrtFAI/7ArnfiI76EN16YH2
OxV5fOPGNmL+YmG8P1XkHX/KCJ5m4RK2Oky8+bIHemUqtFK9JF/SLoATK7Xl
nXS6tCJolymTdOu8jC1DrF77zJMCkPugEC97W5O7VHFgGt8y/mw++3hSp/tQ
5VwFAXyKYXDNf0GNLxV5geAqH1KpXrpPn5NsVbDK0Nup7EJPONsJ3sucy8BT
5hQIeVXAasI/K/5DV5d09iBUy3ddVdiZ5/2vtXCt0mkqkWiXU3dHG+TH2SiP
qC/aClk1rDF4NnPecjCF5wqZZqn3nhZZ5Q8AQYAJcn7bCrqUsoobS1ptSzX2
QMnN6etVehBKJUhAhNomFHnhWibaOEFWtiYF1Pl5lzTT26s++m8kQK5hJf7R
PurTBDK22vWpfs55yRJA1iCFBvw6X19NtnHmPmFdEy9DKiJy+V5aZpbhzJkh
kGonhkciAcpXLQamt8Kgydj0a6w7gfZE6kJjouqKjTDy43d+FYt/8Eq8WRdd
M7She5M3tOR1t9CjlJykbB6uVDWeW9ux4zoHtEXIh5WAFHkgNk4WnUdgbRWm
aUrIAEUpHFUF3ULaEZYKpGUeXkID1mOs34b2MYqfkdx3Zk40+aM6/rEck+k0
X21WXvgPp3ssEVIwfIGp4uLe+fOgW2p4+kFXYz5jLrhD7+msMLHIMPLKCQZ3
qQVgSEnjottNWWFpoIVp5qhtE7kf5KBCkJ+RQ0j+hW3b2nb/z4KJhEkKpriP
NY4XE5q88R960GsZReVP7j9dIps/Of0xD/y7JLsUEPy6R8kGlRgjalp/CK5S
X1tT07EleGvw6x4Npdqcn1rDBCdqjFcqNpuT98tKl78tUH7p5ABrJDzlZlmq
SRPo+IBDY4LsdjTYCU4T7SfjCIxBliOGp7OnV1qKQCydW9bkoDrnZxz4ShZ8
miqJPpoHevEzpU26F8vaRE8v6b/Q8Hc7wheEOa9MNkWHTE4he9qWYXPDpL8E
4pQ+4v4cK6z3F7oPZuWInIn83OJwDlSmbFNYPRtPBIy6ypT9Z2SfcorEfA5U
40ObDI0ANqrES6hwbMO9oJdmLudvXoguU13Ozo41Q6RdQUasiQSjyPf35LqF
vgWomQ79+PtPWiHZUaI6pUpYa8VWWGPK4Fjc1LAhbsoFRUgiuU/SvtnqsO77
bxWpi/2bFBxa/JUKYhpv70S4kap56op1kkwS3Ov9s4fFYxhtHFWLkNZhoFR6
hPmgA8LyMSqKiFun/RdWS0/BPReIzu+AciYz5tI2sZSLybjO496Lhm271U1D
wRGfukm2qARw+Zz9eAJVv3b6sCQ8aWOzOA3L4pAuqpXOp8MBZzwRND/pv3h7
L+4Pf5hwe7rvKOuAFDu7yw1N2M5PP03P5SahZc6TPTPrswAARxovosGbRloV
PtujQAhUxlyIAMGcsAX58EgC2zbcfFEOnG0rdGWBNxOyind7lOGKh1XBfoY8
CT8zG6yHEhO4A3rjMUFGtSC9ikrcVxqx6vLeMG9KJi5kYBmBKAemjjbf2EOQ
j3OzVZaNAjjFYQoyfJnI7dQSdWDzmj8G3Vzj4I4tjojuS4zex4Ty0nYqGnCZ
msV3AG47fTo7jHklO+G2zQCZcBkdVd7NX6HoSMN1NnsWopw8xp8iPFsxDGvk
OUIyzTK4I2L2nnhus0NN1MZPpGF5m2yPsToKSNNFsaXB1AlB89rP5MkIfHEx
tpLNQheiY7tpvYiiF6/sSF0qZWeUeQIg21lCiB4bpY1FTxTUtKbWkj7mxgQN
5hue4VEqbJAUgUDaWZugArh5CuwWi/Y2/FoVd0T6tDLFmBrNP/fDTVp8o+ER
TE/F0LsNrmXDRt8bPVu3qHijliW19dd0yN9Udl6nTvupRUl7w1W0aPuNpNT1
agtL347/MMISOe0OUX3DEtM+CqM3J5XGn3PTA124NsgImMcHFC4xCusCQAwB
fN6PnLwk8KU/Op16iuTp2NTDl7GrTYtGNpkYxtlBQIGcFkh5Qy4ej8edhl/W
tgCXf7dK1vqAbNLkTr2cShtviQ86WwF2TcDotLhJbtitj5Il4XCqVkUpFpTX
5RcKdOgj0bqbg9fHoxcB2nVmwYHyHPK9r5yzw41YYx2UkM67HoBHXM8rG66Y
+IqiErfo4jSaBcyvsyHO7f5oqiIANe2nCRz196xfeJSxfK0YKe0rYp7bwJtQ
SXs6WYkOMTrGsrvwTUGrHUllAlMRo3ciXoJ6S1/xjqRZd0x+0RqXvsewMicv
4ETzg5T+gZRyFEeWYbM3MVxWGfXZYPZVSWOD7tHo5XjvmxXF0R3ciXkZ+/e1
DpqgcBT9dytMAjXasK4XhlOAN7UiaLV1jnlPwSwiJfyOKrHpp2BrZYp8doL4
/eKWt2ldrrPW+LhMRjNM6kSDleW0uKH+8zh56217Kxhgt+NGbD7jr3NuwAji
sDu8XPL4Q5UFStutjUCbDeibCmEnPnpySI++fYid9utiGO72mER111eviAml
f/BW2gX3PbuwWCcZyt7opaM0aiUcP9O+26cB0vhnnLFx/Mz3rAXyHtyiTKII
Iyd52vmFkUv2cfgfjB+BZ2szQ8Xt45VuDQiTcwc+/2ADBgMo2xZJzlHqqQAq
f6Z34yrnExHA68cBjcXtaHipe2oN6AeF0mql+iPDvvUfmEDYpXsBx4dOoUT5
GH3znatWSeg72DZJRdfRtrWYOOjee6mlutMqWxBBqoLWNarwKXLUKYchG4b3
Mcf5UD7oSIbcWgZ+McwKfk3y8pl2ylSc/Ru0JxTqVEn/E5ZNnqqwO8aNv1Qm
b7NQU+MFteyTyYPkJ/W417kJioBaD703dyr9tMZBbDSCY6/JFu2tMU3p/M9v
o6YIIuvKSmwHXPPdC91LMHBHPY1yJiIUDzSHWk8gsXm5vHAM5QlF/pSk6DAo
LRJy0IX35LGbXWlgPr1yAK17ve/jMf/rCG1zap4wXBqvm09qHo5n7rgevEwf
DlcUhVPXRf4qRKroBF2x5+3F3KX4N+u452DRRSJcPHb8lSlZ51BlZicBwKKH
j5r37SGiBdE+ZQHCtc7scoe4IXkOpeJl2EEvqM4Yv5J0JOs1n//ghXjooMEw
Kwyv9RweeBppcdFKAala7RuEJbpn299ii7IiwAunSgLn3jK6qfyHDm68sEd/
QC1H2FLtNdxD0C5D85Fm0vnO5oQMxm6e2iLqBjymliLdnTAtwgcySMiV/zNn
q1ciaZ2b12wFGgaDTIwpQ5M4d6k6QKw3bLfZI2HPqffqlspIEGf4kXWdWQI3
YTBDHb7gVzpDfya3FzuVNhlvBdnnaLZblsAwZMY8QTNh9jY9qCOmWglcK/h+
nH/ZZjLij1TzlKD+Q/QyJ/By3aFxr2h2y8D6uq8TFedZAnLHSNaffRVVxTgQ
IFwwwDGM4vjjgghjkk7oTFQsR6vXB9BWnYr+9VYsqb/9Mvi362MWEE4nvdaD
VdGE4eLsCTxhFHXc6XfeBdQnx+7wJoaYmVF9ImjuTz6BKMGr0IQaN1CsKmlT
f1gFLqtLW0XaaoVXF/ktSktsE+yKNLJb+CoohsAAOkINVS/l0nzcOL29wl5B
eULXSgdz4eyVUk7cGH1F0MVa2BAmyrSAvXbqS0NK8GSUvUo7V/lBKDxM16lE
8LxokVxZbFJA89r505Bb2pupEat215Z0ftY2f3IrmfiO6XMBfCTdj2V0JZoA
acmxebvMyRV9q+QwLCpxZKIlt8/dMPyl6cUbSf0Oh+a8o6ydnYmqNd6WhGzn
vVat4XVxpFWQM91icY5DiKr1npzXZtNmtMoMnxHZhHm8S2y9DKJn+ugiZ6Zc
GGZV0uobacDbYs7KVyIuZw9s1vDgxLwfps2FRTWwtTG9sV3G9tOWHNuSpm5r
4fYsjC0XZHpRX3XVR3V9yPNL8HzC/wVAIVDpWRpLPHD+WkKGTMfdwANsMibB
rAskF/qek9x6a1SbHsHxFWsqzKdEmSIEWkWK83X1KtwDsIzI6RUriBCtGlJ+
JrWPmiEyS1yuIgg4qRxESYA2C6kl7hDmH1ZM2QPK+lHg4LIIbyG6Xuwe3enf
/phw0Dhkaq9WH+2umvfzYirL7CmjGLqPk5auP/lKjREXDeMcmwDmG1hk1Lma
cbcCv5FGdrobboChYVISGJ42bfqHOnp6KXSh2gSx4fylMQJ8YOlHnj5GgvkF
UVetmU9My6JuyTGANw5K8KArkLhVSfhfWFE1S0VIiSaYfHcgAbhhjehys9AG
OFXDKE+MZqNia7Cz79uFYO8GvrDz2U64DHqUHfhpwR4G1f2tvdmFIBZJi1Q4
z1HU6d9MVwDZhaLsB/G/qk0D637ErNr9+YEAzWvRjmodIlmUgWnt4/nhssO4
Xy17wgpMzfTN7ihaYb0y/JG2Ij6FPaleRn6HyNhWiPv3IEXWKnRfhRJW0h3l
mj0aROmxfgzT+fmR48Ek+jXUUtjVdDt/bz+Qt7Pd8kQNiAEfaTKHZkvXd0Yg
Ki8bzm8jK2juj5ppSwLw4qB4Mgj2F+nTqifG3LHcwOjpROWGKkQx4Pdmyq4P
JeFLIkFHt8EIn9f+UoMA6AgWRU8IIa+asYyF4Cz0nkKFe7YA1n1M+PbgBRVR
cfH7km8iZlRvywmN5xgKWLmdvDRj86sckEsjO5pJdrs0ud1kLDxU/PA+qrlr
a35Ymu7j0jfnB4wvP7yGHu0cR3sjKicKIZhu9SJXfSa9UWmHAn0mi0zezW4I
oCYjzQN4qR+BruRq5F0VaauissrF9tGd+pIY6WB4Uu6Zwiakb2g3igDibrGJ
vdlw1RZU/NE1MoDT/SG392KhYd6NhbZSN0EpjD3WXcnpKYBQsKgDWEtO1vs8
lUjSWYuZAhKa8to/AzjE+I8seWapG8S/koFtrOt6MWZnQQsFjDsWihfwjvtz
1UJNyp4IatfqfJD0j+GQ8VtgbT3znUSc1gKETKPRV9xtBgOjByBsccUEat4W
/0y/UKZ9p9YB0Dqhw6msfSiHxB0s1URQaWsheTsUT0T2VJce9nPU2Y0orIJ5
hVAqGEaIb2XlhSXsSo6ulBTQG5JgO2Yfc0Mu+si2RaMNcOLUFh6kdbgMyiV4
olA3QG41ZSot4EjqoOvZvyxYtasBJ0a3it3z+e5y2HdSq+QdQVLGl4eWwE4t
4Q+QtGn6EsE9/PWsgAcvAE8O2QVmzv8l3AOwjIXp7QKb9lu8hySlFI6hcEpY
AZKgTzAY2KHUEpIM6KlNQbtzztSxoNoC6CzHr30nvHY25jJKUxLlq3gY6Cw1
xcK/ENlAHypAjUMEbTYtDqf9I+lPbSeE27uR2XVl63krwqyKOhsOFFrKpz+I
EbFYy1caUhNhX8GQuIw/ESlApa4tdF12yeizkeel3q8rsBAeW92mOINUj55p
yxVkXY9zgLeF96Xadsc1XojBjXf3vLRKPPn6nx26DpJFVEwAca/2P8doRR+K
YLFTFedNoVcKusGY5Pn3cp9XgkUDTSG7grOryVSoi8SIEgjk9zeoVylUjSNc
ji2Y9dZMu4uKUZy2hUmmSSONVXSAmr3qg52TJ+8kI06YRe0rXJgW9W6jwDkG
GvvEOtftYNsa/9QBkqXS7neaEDMwFy9Vs+gzFUpk0CHCwiCkdhYveXEveA9f
I0sO7+0bYSCb7Kcf6ZRt+JcJ2jCf777NdD7b8xmqrYH7wY31aUvwIjCjeZrA
W2uB4Fp6LUcgqyWju8CQR5jnyYwjlmisayNtha8LI0u4BELAdE+obSZpyd9j
ycmUwXOuOeZy2SqM/2Bm/rEFEjxdKCWcYEhLb6mDQMrjPkmFokPOfnvr1YfV
p0xGhoqMi7fTI9QK93SMYBxRdfo2sDwUSkcGwUGTcLuNAIZtZTXShliIQEJS
JlxdwVfU27NOCb5bjMEsje+mVHva4hSDo602Yv/eKGT7QaQBqUYT57HepIQz
C8bVKvxcu10YoFaoP9TnnND9AgCgScGyEFIRKxE0dsQJNeTT2PnfJR7F7s9V
z+vOnlCkORlZ+z50/yFwDjNteaqmggTgtHa4twVZ7DoP8joY7srFDb3ggts7
t8pnoCK0hMe6P57ZW4he1QskboTzKA0gOez/5ypY17OZkQY8PNjVdebE7WRO
0XIWQuZ7mh15YpYkJPepsbhoq3Hf62UWRaYiOfUplJdrLWwSj9o8kTVXt2V9
H5Z8spO+Asez8wldu3pVUH8M10YP0nclUlmL7codCMk21vRtS8vMBDRTqX3/
sLC9ETUCGixBMc8ZvM5LGqulBXAUuqMP0eSWvzcdQS35C78xj4oXnLTYyaOG
ESYzhbjPheLqTW+vB5xoLyhR1X+kbkzx2ct69010NW6anoTI8duLvJLKgjQu
ChWjJ/gtu84JHR8DmL116ZerCAtJefa5rJUH4FxMYrT5cFcYXwjCIS47Dur6
yi3y4gck5zG0Zpzr10hgz5ldQ4XFfeyHBMlEnMJmcrko842O1FvukrGu5L5V
+6+xYXZmgxiZgBkVJbzMDa1Sl63w3EPZ8h5qUvwdo9k0ZvJpIkWOeZs/Xitg
jMuS2sTzjPAehXjwRsiGsy+oC/sqTHVqQJpBC7sE94VkCfq5tTF9PCIBA6/w
WKwfyGg/l3n4C88rVCilO8rXmv9wHrUo9niii3SZ9wOMRc6/Y3kXSXba1es0
Od+fmWTl909SH8YQKl3cu+3tTarxaMbUVQ9H0DN0VHtipEyN56j9e9V6FfE8
xX3t0vFU2EhPJiz05IuLKucnYUBieoxy8uptltgJnDu6K8APIV5O/8N/HpcP
WQDqUpsyqZ+8nPZvEBaPbmCHUHL4zy/Q6AAti6uUEO7x4GgtfZJ7joAlsJxM
wt/ztu32wLq79szo0dOW+wr1pSKPsFs7TF5c5BUVqrqlq961m5sFudPJJGda
UBtrCNMR0dzrZQNFmUldKzzdUmQT3fCQ1BusycX2Oftl6x75/ZwGwqov9aOe
d4Cu8F6072MfTBJWR3f8b4EUpYe1bl5/b3rTmf+2yP/sDxCRdkyukD483KF4
5vA1swd2Xjy/JBl8JhO9HY2yBHKPYP9byrthETlUhfckiATL859wMStp+NyA
UAjVhir6NiLaLR1Kb1cgXzIad1xE8fwth8iDfwmeXtqZWBUly5eyaFlr7PGP
c9ftWK+xoOcIwEPy9Z/jzpnDPt21NWlu+22258wxf77JpvWekyFXebUZipTZ
/pU3nBYiEzQRLAxmFQuj4C92s+QNc/IY381I/h6IKWFFmj5orbdobOKi0Lar
00zFuXk5NcDDdxV4CMDoP4YMm+plRI/5Ge3cJPwzNWSIuZw/QeX4BerQxgwy
qmYd3UafK+7DRyjZ4ZBZgZ3Sb5sol5rBZFDchMHUkX/gienw58KTqaDpWYA9
V4dMA1Tx8cns1NgEcP5e23gjebQ1UndmT7tq5ah4ihQ2coH3wdMJf4XNA1kX
a7FP3cBYsx91m832G4XBrgNDzXV4dN5pY9ov7UYbwlSHXfoxCXF8jCr6PVBf
pc8yRQlu9N4LG0vL7d/8WSusAM4/5VfbS/qERCKd8s+jEWQ7i/gqqBhTfYQB
H7Xk4YHy1t8dMgWTCKJ8gprkH77zMo49zkopkXxneDyj2yBcfZqVNqna/EJy
2vyGE9yLbK0M7BE+xOwgBgaecO/Aatw+ykU3POR5iTvKvz9JGX2qFC06nIor
Ty1OTtOzDWGAvLu8qfWPVO0wsdB6gbcVa0twigHAYR9ffW1MYxPfdkWNt1r2
nnlzwo8IOrMOMAdS2gLSoY7sD/d5+6Zm3BS5G3uN24YnpvUKJh18ou+9hwF4
cDMGXjT2i11r8qu0bZ+Cm7VuZ5yqkKilzVu97vY1HJswsqNmqqklm346jQ6P
/k5Smp9UUkJPNmPbaYHemhRE4ka8ZwcZaYYSIAqzcD0Cd8FARaU155cJyCEx
YHUg9c8rL1dbOIQYIXEGx9YVanN8VydGvAcqAnYaRlo1SDMTpEhTt69pUhKM
OgRJ7QNVYlheblK4M0+p9MVOOijfVjRSqghl4W9ZAKHFZvN3NxlWzMLg+EaJ
Tue0GpAJr1i0qVdK6MI3mYZ+Yh+mYkOqATlOTjhUDDeB8DLGHXUBhegfCd49
0kyYu78xQqmn1XgJvw+iGvwXih76x0fOore1p9ghffWCoOpj3QjM2WDB14qb
jWY3bGAY7r/s5w/+OLF0wZ4EjBlZOM9piv/dP+llWANgI7oupKRRTe+ny5hg
D4D6/FikC2CggNoEa4U+KlanDQatunlPzJgaM5OejRHyyMrGIfvqJfWE1AQE
xxe39nAWkx7J2OClWZNjo2zEIW9x0JBNWAabE9m77RUA5qUL3bvmXaDYgTZb
6d2+S6QD7lH/j6Oc0VkmX8B8XBxNqeuTIs8S5lRy/X1XKLvzVL5OmomLKqfU
XzhY7JNgUH90+bXVmtt+j8AhV55TW/dwaxEAoCVcws1eWsbSzcSeZiqpXWoD
uGYTS6TxosOgEzRmnOHCBSgCkcwPbuMFP9gb5RhyzRT8KkVFkWSClQbrrUTi
d85/plWo5Tk4PyADdtBaKYuKwhgGH6VFbL0/zd1DFhxS4LZVd95A3qeRT8f6
NCrZ1vG7RQ+jQ9JARWrkUx2+EvLTXfmH9PQ7FBrhAGu7qar7ZiwhREgv9vcl
E2IjVs/c/fr2b+oNop3eNglcUiU7OURbRDUGs3EgjnZoGHF8EHnNVSajXgff
+mKHHLPtmtwXGWY0js8SaSCbiMZnEHQlJsjWnr7Djev+dAn7Q/2u/m9jLuxQ
6M7ooR1xlioWTa5NIZYknyjs0bh73FyK64VBEMArBBiMBsxpHEZZ2WrgLnk0
z6DNherNZW72qoPy7+ja55IqECyowzNkkzgHJ0gx8fzK+5BvPHI5muF9sTd4
HGasT3EaE2moAplDUQvAGNojcLM7lUk7A9JsTeo8hSGHgHQAgsYrXsf2xXPG
ljEpD24pxTanW505bmYRB77QANuwR31kK4YK/qztLFMhsxWLxV4/+3Z3qNkS
dJEH+qdYy+QtbgK59YXzmjkCfuLGcE0TYPxUw706/bQK2PHYfneyyGiiWXi6
kgJbS7V7Q7v7GtIFfeOq5FUAaejepYQp4of1L513v2sGNhvDivM0dfqDE3x0
RdV2IxkrsDV0osWF2Fu8p6tMdscDaeNUHwNBxHcMr9s4ZQrZjhSmrwW1CVaa
iLivLI3ywVT45Pb8AKtP/p67vG0wd5MzhbM1l01fCNvwWiHMAWZCigJCoXCo
r4uZO1loTqTejkG5U6v+ZU3VkH9A7oTGOykS62We/7OwigfioLgQb0ZUYk82
ZlZdKIgShJ+3YDoPDG9H3skOfDqAlpCXHX/CwZPu0dLZHZ0ZKDnC8kDRv34U
Cknog+51YlM9kM442wh1pyu6VRnXf8tFEW6z6vKdUX4zrbPvP+/P/5YMeeS+
0dg77fmpnfpTF0xaInzc5mKWKidVwKk4eSiKQYkOwE+1/pa30vyMhbdBIfL/
hoq9kH5WsbvT3RwDF/MzdhMtyJ7y0rA7eki2NPUfBIWN4f0T+LR8NockJqB9
448AculHGHU1JzT0qm3ZlVMnG4FBLzIxIgCLfwiLPL0AkRuj54J7VI3sCIvs
mnyA3gtT/0Zeftc36mEd/O2nmoX+flAR1uoEYmnP0Oaq7y9acLNV1ZtaBuYC
q3WgGhfGSmcSXraBfSqEGSglmTrVHF5id1sQ62BLAk8JYj8zA4f0M9WI1z33
AIl9aZKBwyY1QuKLqOyOpm7vZQmHh1iMVYMIiR2xwEbr2RLXFDJrqWmyq2PL
0Nyo14o4kQomnjaGkiTQ3DMBJYm1dlBxETh3KE8FKyIbJR7yq7APUgAfxwP/
DV9rnb1/x9WSKFBEc0eoGe4hebE4bsIP5aq4jflaTzQ6g+j08rOvyYdwxS4r
J3Md/njQKdO2pJspm3GtekWIi57whNGz3fIEhw0qWQSJBJZq7fKmoMEwog39
wNspFbH/GXRKvixcfGVlOtkp0QZj2U47SiWw0NSsbvENSdlm1qIqiI+2aoBw
MgLILKL7bxgJ1doiukXBA90XPDm6sqtpp/J0b5velzeM8ipSC8WWVXcVZ/08
bMrjBFWU5j4W2gTQ0/OlTmhrNAh51f2hJSNWVcmnqxZsCRIek6lIFHSlEm/n
oMcrmhLPeXqDhWw6j7FkEsW9sB/iKxxhAQF4mxWhoSCpp0+JVbnShVXKkBr4
IZ1d12o0JkFesKOWX5oTQIxoFqdjjVoZmxay7fPDhnl+DbpiuudDAN+MO/H0
+IecbqT0xGNgjUNjD+3BYcXhED2YSGjgIK5z5fKtCsT43+1JYBXDdGPQr14l
Yv2KRMy0Eqkx5I7fEtC+s8PLhYcOZJp+cwwbfL+rbs494iID/tDWoaiftWol
QTHSkRLhMtyWFLqSgGbTQ0yb0HVVdgqxpENW158vDjXYqFAMJbBxm4hZqVpQ
fh4lUwbl6qJD7EnKE2+l5TIExtnpVqZVTcdRKdUL5CtrdbvBhXwVKFTUk6Km
5OzB2vFeXEDURRCi8MqtnSDqRmm9yp1WPv7jR9qougY5eRvXefnVEH/YRZ93
cqj/TI/8omktuI5p/4hzuNmQGuU4ZQQBgJl2swX1LCTNXWkkXz4UvyZVUb2I
DUD61uJV/TPzKpZB8xq4Logw92jV2+UfAP7aZwa+lGtroywAPSHY22+SIQh3
uxgECezWJEl3fGLqw4pFYChqAeuTOAG+Y7iJyV5Lh3m9PaCFc2grOieF5tfw
qYk75KGh529MC2Iaefzpq5YShgIqCwWZa5TEqYqeTBWbEArSVHqvuOeOa9G2
+HDM0tPAX4oF6jDl3kE5V4Ius5LeSwS1nPSpZe4TD3iDY+jemgVNSSGknb1y
UWLiuBwKO8hOghGFghqOlt6OtvYb8zfr33RVJ2/ex6eSa+hOiHDgvRr02LfE
4+U4OEiKXBWX6DHBjNPvIB1TYvQ5yOKGXBfrzOVu7RcYkIDe0t90UZ+cwe0R
nAZ8Zp1+CFSd7e50qvGiJ7sZIF6Nl/8GsldGyi8BSNq2wecr3OFjCHc+H0ZE
MBQyjN3mRsz9doFZjKkHHui7tku1olIENBe2djFCB3zVIoAS8qSI/G/lOUbC
nHSjo2b1uvcf/Czt1wVjWEEgFpD6nWsb18aAuhgzC24i3nk22wIx+68OGoow
/ZofcUe2dMwNSY5u4Wrh3cicZ9CYvh0GE3dPGRz72RE3+YKyGnIYUutxVANm
vYwxjAfWwa1h0DHbHCrXMxw+VtKgGezSiXGxnS2TADar0O+2HbE/qEGabGB5
b2v8+AU/FyGt5Ug1ihR9MVAZdSxJlIkPSzVaBXatrC56z5slRH5zFDjAZ+Fa
2vMqTYsXkgRjYm/CM20tZGJ/n5Cx8P3+IcFE9sLRcbplTIGiHUj1sUwaCpRM
DvbWasIqWz39y197WkpzWBPqiWv1pc7pTrc+lkVfCQOs7Be1zjqF7/iD2sn0
Q+m662dPYLClzdIFxsBZvi05/Ry//TimszbmCMWuaSkqbNme08aijWzw2xu9
2GjM8NYc5pVBCsDxdhIxY81DnhhdAtzMBvJhKBactelyizMhI5+UnGvNcXl5
K0Z6YsuJuZrJezCDj5EPkEPTV4wXu0FRqdHcHvZdn/WAUqy8ui3Pol0jbxFo
SfzbiE3Yt6JBPECC06OJK29DfwCC/joTpDxO1jh6QuWkBEtmdAgs7UhCpSvJ
nTF9m2aQBSDTLbzSidu9Ml60ttVywNnPbWybwdUePuRwPf03ZDq6Wn/eiTEJ
2I5bQQ2DmTdLVOkkp1F9TgIErEomoVTKnb8JN31peS7F3OQbhMuYsohWgjoT
o78x9g0MVGKRKW5VSV/KsP1OmBbUrFr6Bq+3xMdmMOGar/xd/ilIRuo5a+9K
kn5lY7YxylcsEGycfjG4gDOwmiY4rJcqxi34CjPCCOwhRWndscysCGPFZJer
XeOEvMUPSTraikDRlNDrRO5jBqezOayOkZy9XwUM0DwcY1xE4vfsdkN4Fj8z
fYB/QNDaWV0y6kQK52PX6ofeV8oJgFuJBFEj8aSpTF1n8XEZRNbFxt/Yh3Yb
+sEiTZPN6XPoALUl6aBGfdhVbsXHgGKca/joMMxryyqrG319ukaFLWzJlCVg
e8xQp64GUzqixnt4gkMn18tuUZUBos7sOMz/rGYjCtUu3C7c9RsTBFDVrFfd
w3tmKULQXBR+IFbQ9D7JxdWnqYaWNkvS1276pMqjDm/hPjDhYus4dhH36k5f
w05ym5d9QQ5cClqpQRXLaRVk7wpEzphukmEgDQI016Zl/fCyY/ypAfUEKfI+
GIkecaNdAQYPrZYayAUCE3+53Ec6lOrszXFUIMc6epNUDqDzzoPGMGb+jMT/
jk65d2r8KJ4sijePEubNXA7Osq5pFXvZc45jebBKr7RjWJ9yNl6ZKH4SxMVe
Qs+0LBq60d/t791ufJMQwWL08+7kCLMtDp3y0IN4ZYa7YI6+74La2P+qMSwP
PAS8v8BSHlGlts3WdqddICtJMmpvfz9Quqo/jCaNKos2n6zb/ziCM3Kgf4ic
IzOP/gVlKpEWXFjjwpdCjPBV4N22qdqV0e01rtZUByXlO5Wc/RiREgRaryhg
r4C2n25Bu7q+mqtsrbYttCmmhJVIuqBd9jklJ6PCBFAyTxTcpm3qbEaMetJC
cI4pfQxAQyoUwPAuRdT10tiVNWGSM2SQFz1MHieLSyQ68G8wifgda6vF4bbt
iKizEi4LWJCoC4X1eEUAk0LeSzffFSFG65h3Qq8cbkK4bNvdn7LgrIOoavOk
oZxH3e1ZhaEAwKIaTbUeLZIhR/KElNDIGF5lJEQtqZxW+QbqA2B1D0eOGaTG
e0DkS61W4+0zoW7H31wYMIgPqkV1Aa6bcn+dCkjHqKA5nPAgIgfkLT9+pMFU
lf7vOVVnqlpT2/EYAipPBVKl4w0ssckFH7+087vu+nnpqDxnM/2dIUJM46Sm
NS129Ux92baCdM40oQ3t8YK4fjdOVkUQSdZD1yTrBfHVvfFokt60Eo3H5tBR
Gl8lRqFf1rcg76ILRe9FUJi2GtNLHJYCkbkw546fHkYC+8MDTeV+1yhF9Adi
/96BRwZf8kcha9+yF0mUhs1MF3KYixsYlCZbKOiusmt/wfXxY1FlS2LK842v
BPY+Z5MjKUhZlaiSDqJlqLsnXNZvKGL42HJ/DCEHqIrBniiCBPKzShPxRnFK
2xva4GOQgMdceYxvwFlB9c5Oc7J03j+kgk7N01GfMfm91pkatB39fXZe9OJo
J2Ur28GHU3aJUGkScz8037ejHORfn4PEtgayKjaI6ykfJ4L+CykS9JgyhaKq
bXQjqDAKo+DmrSuXwAI87J3IusZmuNg0qN50MzV9CWcNE6H0gySaESStQO7q
Imy47F6vmYLka3pj4lS+T72CtIrnxBgF4aiKAgvvk3aL2TJFdkikgpeY5EwW
7SbprDfsRnyW+KK6bqBmpHfcxVT7+cFOVmX63XOUH/7E0ekEUQ8mu4DAwBSz
Kpja5NEEiAc+uXjUBQtrFDmjsEykPbEmyIHuSVEnT8e+sFxVLY1yyTm+dNOI
NCdEuegWnHYfr1AIjAQN/eLcS4SOnN/FErS3dpA7G0d5AdPIzT1l0BAxr1zY
jLDlIXl3M5XIiKJRHhVEl/O3k4IUZvhm/RSnUbgcMyy4reNk3yg+Q+QzyO3e
sbgv/ANP14WqsmpuOpScSosWVofIKJwOYaCA3sKBv9gGHuIcJ9HmorLCaEfm
Z9hYU+XZs+sm25YY5IwCLlBs0eMqB75r8vC8m44+grbFp4pOR61MS+k0Lw5Y
0/ccq7+J1aOMqcN33iDf3H1QRB1FiXwE38yIK91icY9Yom1hZOQ0QuI57CU8
GL1Lwgk4LX3GI68BqOLhn+jP3ecxzJyDGtlhQIIWpxKdlhox0vuZ8sdJPYR4
hRHM04OOBN7nBZPT0eZCDfNsAEMi8dJJWhEsGppBtPLreimUAhRKXrDP31a5
hyUjOQl5j4EHZ2uNOjhv+axXnxIm8psHgwz3+VAI3UZDh4pKcjR8jZJSPRIB
fyLho6aSOPr4O5beZoiJyFsCGxH8r2cFIbjt8aINfaFRJ3XKJhRy8rP5L6TS
maLLFPIze2faSfjPA8wlX4IakK3OSpUL7zqQaUlPNP1rP7SVeFmtEw/Ww0gJ
3JGErYQCKbI7BNRN+CHCNPf3cVbUUSzilO6HQ20MH3EnI8ck5PWmM/O5xF+4
E9CvMuVxv+XRKpmh2ZlVgUqDInOluHYTr87g/no0VHmzcG/vduOefFipPo7C
HJx2s8FL9O0B5ky34jXmZDz8hYGOLgx/NvOhJP6K6lCCuscb3ZBb+g3ihLd1
6SBbX4toK1LbmIBufmMCh73dyLrTgidY3LdcXk51Eqd5zjgBH/ZJC6DNOD9a
7YOzH5XVQLlg3BLLbYEQ4r0LXR5Z8ifviH3kliWWMRXvTdRa7/W2+dh2OtdM
fXrjG6+CTQLvSfilrnOl0eRJR2OJW30cvr0IvKT8A7ZihfV52DCCjBSoiGmz
2Q8SA89NdU3Bm+2Ys+f+Q1UrJ8bmNcehUheEcIumOJI2FSP78467IsHrK6Vq
TT5SqwonbcnvqiuWZTi58PWTk9Dua1SlUKVDKHvPHV31no3u0ZQorZdSFfRQ
2maZ8bCZQ1rkwgQ/8RNKW3jRNIWmHzMGgLLrL9mtDo7HFjJV6/VZHUwMyYCj
tTZJqieKxtBcWnNgR1evYKyMFpULg0NAeMyqy1bVtPOCj7WDz164WF2nC99g
yetWbhZBkcaKAe6LTZwIQRjmvKxlnsrJ+ZZIuZqW/9GhjhH3h3YUI1Gzm+Du
k7SvfNyqYOSa7FXmVPt9T1TMF4UVbJw5xtP4719ipjLeM72hyGmE7n+Pa+7N
Rlaw5nxpf7HMeaBamfhv4HEKhemiOohhLnQIqWaf7g/2kgvt9rumh6T+6krA
6X7a7Cya1fz6yxelbMQcA0Z81TGQX5e+z+iHlQithJcoSi+JTmDK8gm70nFf
HmVPK5S6ENsGEr5Y+gwsK7/zC/viCPSWL2tF9BCPZwKA6nvQMTk4JduaVGuI
LPW19+QuEEOZbqPFv9c+jG8pWcq+ZR8kjr8WmNjqOd4TEzWwn4OaB9k90NwJ
h5r2f6ja2c/S4xzT1/T3SS3VkuRgntfrNflWErsZW8cIPKC0gtvQ54R1JxB+
rUJEiaIoTB6pDdcxLn/eTiYhtf7c1MWGJmnQygMrlgYZADOGr7dA9irWwkYv
8YgHWFMqjXy/wXUYho37+a3eg5Dsdqr9iIhtTcIjJyls5Mk4/7+xouqxBYwt
8PZh+lOMbzppuW07GJmHMuBT0uUFu9yBMfByFe+zrjMPdfdG0IzBHaedMRbV
1IoGBqR3Jpv0RtJMo8Wsu54cO5oRWKvkLuu2KHhhGAZ1alR0chaf9clRczbb
mQAvBE6WepYTebtdBr7l75x89G19yVK4msLYqvYjsMzzEmIfv7kx1mnvnwkg
uyrQQJxc9TnUkotk+6fQW3mohld/xCJ5kXRYBnAnk8W3CT64f0OxkHhkFG/J
tZZpuRz2wIDx7N89A9g9QUS+7D2Ph2FGcqIrhpEhCYLZsP/NETvy2Gr0zZjI
DzSIeYZdN7lW9KCk6QOFTwLY4I1Dc3SSSPH2I59pYUZc4ftIG9QyYT4Nrm1m
3uk7zc84Tj08lm0aRH2y/gyMVvjrl1n+My4EEUO3n456HBnw1aYFSsB1lm5e
Ovk7cD3POiGt5kpUHfI1D81m6tbjlCglxUI0zP9vFplTjHt5ONcuXSi5i2aH
r7l6mfhaW1d/P5TGUfXSZPKjovPw9iGrP+kvyWeEIZ5yK1/T5p+TGm+GroGk
wfaMFNYsLf568qTC6LIyJl6nr3O38aSoT2QDkObg1aU/r+BGVhBBTiw1bKM0
hQ+fjrPWAwJxcoAy7e4836d0HxVikrTCNFHdenTy6Uli3ifrXY6Yjar4pA6e
VkoaLXM8E/plZl0EC1Du/d0H8wGT20TyixcPN+E7ax8i4Djs0uCSSWyQB/YN
Q0pOnnVgIh4RzqeK38dt19bkDmcHHP/+bgQOeIwP9rX6zaoZ49gIsHYAshSb
fzCdA5WGReEmbQtMhfC+zl1TBhdd5UuAZpquZMEJTDhE90o5EUK3DHqPlE8q
RjrjDlRv8N4jK2RWQSM+CZ9/dWbbFwZjQWMWyHSZ3yF9D2PD2yuJefaF6gQJ
xZncpRXA9JsVEjnqN5QKJLuyqu3DByUZuQdHBiNq42b47nvcaA2Mu8dK2GQN
2KsdP3bk+ZxFB/KmbbmnTf0D4w0Z2DG8RiHlcdnUNbgx+5Ag9yXXyT/YjWR2
uL5s4H7qH7z/PsDUH8eHYQxaRGdgwKMLkOEFwh39BI0nTU9Ym/tLtHcE29p5
Ce4CTlHRYzDbmtbMaWRfAbqgYcyrPajVHVsrNzpMv06nwDIE+yXseCCEi6Ro
d7E/UTBIdL+ltpf8D4kvXALz96rk8XZk8JCGt4bjlJNZDVJHgqaE3Tz8Sdt9
GT5ccSAwXSZEtuWCHDucxIVlFxlKZBxBqi3gX4m+GW6L6X3r6KG4zU6FHPdr
M1Q/JHQrNl4c0h5tEA6YPTqHlrMwp4qclsCpV46kB4EkkI6TGjKAHYozaoa2
3zfwWoroeZmVwnxqXPJW7F5pX+OFrAiOeIF/F/yP8ztbOpsAiV4RkyJziLsO
4AcKXfd9nlU6YqPMH2trx45A6s5kXjE13klwJiq2h6iwAk+7QOxWhbbIEFdx
+P4jib9zXJlPAEof2tUBF5BteoRb1eha8sZ3sopSg+2Xa9QxNPItuReuqO1m
1EQv4g0SNWntT59pSwe7gpW8EZfRfVkfNiM1ScM10Ie8sIyzpveXgQt11RSe
tJEhtwTilc0l695ZeAi1FYMtc+IZ4VOjLnrzHBW2LsGR5bpPDOXIKbVElME/
mq6QGaD9gcdigLB4qJ9mlMkiyEBlPhwmxjgPnPsdFS7G70GLMEvqNJAcVda/
QrL5QYDkXu9OZMDniEyFP6qKsM16jOJtYvQigaTTssdZC2z64m9t5e7GIhdD
PkztN0Sod/U4ijXMNlnodgPG7t1MH8LN0NC2XK7ch/G1hYBcrk3vRDVUEH8q
zfz5XwmMVNfZAb8cgwwLzBhu8nNQno5QU9tCSMtkcCXD/+v7LACCsze6TByS
4tKmkwpEuAhjCZKArUfPQmgLCoU+FbweaXpNfMJuncEFCsJM09Q16jsds73c
rLmABNimI8+hZk1pXpU9UW6h/+USLIF4YR2tq8O2M1eEP62tBHkZXV3PNrsI
syUJBhF+WeCfRTUQqFAK9AoCuC7Em5DI5wq4JWuwZLfEAz2nO150TbEh6qfn
vSeSQsB9BDfaJ4iqQrs3Yfl4hiasYHAz330/4GOfIGJwtUnGh455cuL3VVVi
+IO1ui6ctQMcSLja70AxVgwYjfq/T7Jv/d3fsIwGGXlaCQekBbF3NQNoQ+xu
LnNc0OD9CHkl3m5hWTjs9/Lz8WnXFVaWGSh3FKjS8zfuv4R0W7lPSwxgKzN5
DfGHClbr3QJzaJlZBsBZI5xXj+80Zf2R6v8L2BIYhCWLZ6EEyesgDmoqnhrp
Wgqlk3gwMIuQXiDVGqf51IjoA+e6+Y6zIJyciM0X5hZeHgi8v/kY8qTrxp9T
5YSlfxeiKVukTlSS2WgVbUqkrmID/T68arCZroXwC2tagJ/B6F4Dpa3LX3MH
dk+hJsZLit823CsWnpYvY5b7hy6UzduGS5mCnZVNfTOEgoyM9lPSzkHtbCr4
a7VtNzk9lJMiwjYYrtrI9bTf0L7hGDu3vfQC2tUHsX/qvKYxb/MlTATkASYn
LmgQDv6cMMQWxbo7OXaTO/Waf5cx4tVQYvIFsBW7X2sCWpHvFG8j522m3AEe
7yV588Pwb4jVBUsHgYnAa2/rkBfzmfREYaxwQVOfvQPXLbEbNOSBNJGbeY9p
EMi9ysO5c2ICYOgH9oyEv5KtdqnFF/whL9+ncoEqhM0+VE6sxrN67SuICupA
CQKzTDdp+WQAsFOupb/tShNqL82hTjQBzF4wupfn7PlLUpsNSa5GEke1cQCV
CP8cA5seIVsLRmtTGJumvc8GapZ9QBpTqJd3RryE2+XzFrYrrtZBjcCkIhw4
jgz2ecSkiZRmS6sjEPLiwdwesb8o8yUqHXHbj0TgCCzVhc/5sIbfrVh3oCma
PR15mZhLTw17aqh3kjxQXO8sDG9RSl38fa+NfLUw9t9Js6jEaUk40Z00Z3VB
ran3grrMf+Dn+jmAXskSWVKFzByqUnh3ekmddNatrlUeoIIIYXz2KbtT5BPK
MBHWp/rrCdHOVyRhrxnChNX3A198BXZYewRB5WU70qz6rlwOTeb0d0B1gfur
/ScIfWsqzw8pYlYl7fG9lrdYQa4bnq1O/1ZnSG+mAe6OtjMTEvHQNM8HT0YQ
Am2vSVVGiH7sqfY/RZjPT253ShHiomhBl+iEfNQTnyNCFYgkfVSvFoyHg44s
6BW5i/eIy2HbRSIkhOXxD9qFeO/daeHhuU0K16RQatZ2JD3qkpNoSekmPo9j
smC0sCXNmtiU3QiVlmnYJ95brKqaYs8Mb2rTigTw+mU8NSDJZzVV1buy17jT
pDFXkTgz0vKKWCmNTlXcntLtExEjYJawEeld9BSxOxj3lGtimWaVmPCRodOn
7hlm2AZiW9buPf6ADxjGKrw6wDu66DglIi0BvHFZWPXdAPvWOmpbG4uJAujD
Ws/uq9NQ/7yn+0SwGFEaERgKC7j4nsVAfJS2bM73hZnr5kngO2CJUQ8V0JUF
MOOLRbuvqYKlrI4Nj1cA47CAPZm9jwUWIFRD89zkf+MlGGxdPulLQSxtiXv1
oF1dCUdYzE2lvjiJH5JTXZfWRTQblVlZ2IhFdPe0DAXCPlp2wG0N3oEanVHB
WX6nkn37TIBnRIM7R0VmRXTs0iMgd0rY0ZLw4i6Cc5kUSJ43XE5PeEQvePoR
fuhlR/xwhVPteg5zCzPcqqaT97xqa0xPxi9mZMSPrHoex+YUky1K/UuIwiAw
ohZQZDaFjStQi691nEzuZPOJVWVNxyCEwGciewhExz6TvN1nIPV1EpteJkZx
RVyr78u3VFBG5AlgYPyKdU/bPIQWNO5C1Qi4bJYL29MKwu35pfcSDvX+7r0c
wUvioOnspZKv1dLd7WhMhDkvFNfbvFxOqnGt0d5x61pW0l7dKlzU0+6Rjyu0
8SqhvROnslYApR3iJxBAQ5HeCx28/a9AgzWDYY3wjWEht6PgmczrktqDQH4B
B9kdq0dDkxTVULCceZPc/1LK1qFhGkBuE6nVkNHFBnAkuiJaeHpV1RxfzCO+
kVOmlphR4HSOb0rbNfC1UMAM9Hif9sxm+GjGUNn+6NoGXicS2P2P9c5pTvRb
Fdu2dLfIm96hePUStKrE3cLnzE/bS3OB2l+2DUOzxvaDEb/orbV4z2VYJZLc
gEr2Usq+NjIExHTkJht/NC9YQgL1jTxZV8J/66U+vRpt+EEtN1kOyywGa3fc
7ZMXxWdlxI3zsxZ8Zh3AVoN7uMygWNQRTbdk5liUaNRuBlQkivYXZhqARdet
e63/fc3B2VdDoO6XvzQah7LEj7YXtcmeXtlzaLi+zUa69sUUHfB2BsQuAdlF
w0twnrHfYCfbt+qBYxAIoEr7YxQsOYebK9jFb0S7qNPCLpz9tkSupvSfvkcb
pgzQUJ4zYdMVVtUH8FfRrvqO4rW5Rlntm56pEkZrOB+DmTk1oGLD2iy4yvM1
fTM/TMrGKST+LBp3+OvqsJepnIPs/6OiW8e3lkYc5lLO43fObHyadef32Ztf
qMibNDGMWhlU3SSg1ysaZ1HrqSCPJjSJsfFm1MTJQO424TqH7IimMhCdIpiX
N33Wg6ybzBjZhftSrTwkQvGeDJOxl3nMawD/XXwdYrH/q5XRrllT5eUfb2M1
mTqHFaM40zec/rztzdH40oKUgAmCXG9IFK+d5A/WjuD4T9Gh4FTtTPrcLEzc
/fa3KjRVTUrW5BWrcFZhPPTGiqXzL3mh8+Z83+RbEo8jTX6u8Ful6px91uk+
zU7r0wTKf5OUvmqV8EdT7niOEPxG8+/mM53obVwKE8jbX7wpZOx2YsLFvBgz
CEyyANKKXunGx6mqz364czLLeMQNxboM2/T9q1xT1J4Pizs5TqgA7jy8RvuT
USYEt0AEhpgO17fTJT+K62DTvErMN1nSJhaqOqD8Z6GOWKtC245H3bFv7nFQ
zCwG3rZ+FO0SCAFFSfg9SzlsNJmQRxNN9KqZSODZMUcD6GeErad4mD5u/e9B
3B+Ypx1wguyhusEhPvFOow0wXRxA+4j2BEV9oiK2cW4EobAEKnVSB/tLwv2c
H141P/gt8rPvXlPJJ1VgcVGoeJRlHO+vaQR1XcCF8HLkvlgzSkv9LlBN57/E
5FyPg0UBrYvDm84QzoSIfT/To89hK5tC3YkR5cpuQHFr3mS6bfEbQbBCRklu
5tErWZWPHYPUToesxPlNhF++zj5T4wIZn6V8iQGYabuDhpZCpqM4F0NFXr+S
DE8PtlGtlGSHfCXal34P5FSuGBY3sJCYNIuJsr+weub2lphYg40eSSAXHgs4
U9ao/6g0BNoEsfaABiKB0qIz5+0GNn5RkZbDxp4KNnz2S5oGxz5loB6cCe0F
53rhm03X1lRoPQF2ioGT5q5FYiHHPFtbQLkf6VJtcogD3t7rKkX26pfOILY6
8etUW7/OUPQSopYzTGTsLKd9KQnpBAfyLubdEAwfw5cWmPiixVjF4Seqbrwi
vO42/f1jJsbR0bHy6oZ+j4wcPX5XEyNGlNvrSWWrybfML5PZ/8ZWIyjdgHnk
zn6W+zdR7q6gBVqR69iyNfZmZvbXe1P6ie58u4rqKimB4RcVymvCiOMbN2gR
L74occPQxsdSCnk2MaC0Kf0uBeazH1paC6xUFhSmouIgrAw7TZG9nPruX2B6
TvmJIRziwpJwk+qjslOZgqMGPE/RjKsG9kF7V/7ltnexakCvDlPemriJV2Z4
N3zpnnUQudqALsdmXSgyWk/i2fyL8OLdk0qTNXuzYOU9ICZRoXaDZwlWvz+O
WY8ZYDhp+cOsrtD7y6nXM+ASUUuzTEVNHS7kzVHoTejb8zmkyT1jkMaA/lUu
sgToZhxzLFX6p+9SCZm4DTiE8pYbxGVD7RfvWybCROtmO2XrRoIlxKAcDR7/
4VKZyz+6Ry3t8h7hqDG38GVDi4xXDYb7L0CFI5cIiW7+obOJlqrK+7OXVDDy
AQRnHvYDUy4HWZ0T7/IR0WhFNXB95RYWql8aKN2aarnDBcfZt6aDWUOjm8Ns
w5BPk1+ITJX7qAXdYYy38FjK+qKCYfIOER04wR/9o3ntEMoFwmt9wkMLhCMN
kq3xLgLcczH4ACcCKXLmHgbubfTL/liCIsrU4UARrXIj4vkoxN5Nh7sDGyZf
xOBlDss2IkxxNN7fraK3yKkHPOtV/w9O4yLZx5HLshoJzFHZLRWcj31hvR4q
n9gcSNaqGvccYob5VqA6YPrimtjq8dFouOzXGInV2ecnIKv2TOuruH0LnkAd
wogLzBh6xrfIs26foWtgiqwplR2VjrP8ux8D+XCKmofXKQkqKz3xiLAPIqUN
YUmNiBQ+T0UjMIz1oKu1Gz85JLjg8hSzzOdxUwBXgrFg+j+DDeMVf4f1mKpo
8Gcgs86LAjRsXktC08bJIKEASAI+PuOFerQUGsyHVsyFmpSXkwhbmcDSWo9x
TDFEEeS8ktFHdqz5zErvR4UbPD+vJfrB2h4AnQUEA53nkMFuyZ7/ASFi+OXu
5nKNOCgp0mBJvmSnuVu9qOtauXwJGmjL3MioAkMoozPCAGElDJM6B4wP+QPT
5Ic3R/UvMgAPUckoN4vq6o9jHG0z8sdCpw20fHn1QV/vJMjY+Vfb9XyHhnb0
5dxwyhk5a82Yggfgcs6pd0NqRmNjJwbMld8wXL0o1kf9SUD5jub7oGaeR/Hp
jHUY0SYzgHtL0hxzs9BRy2/+MLtuR9JMSZe01M1gu/pYF4rfBzvpGq2lpvNE
b0saL9cmIPjMW8UmG5e5N9oxZ9SOziL0hs9Hx/S5CQK8R3VJUqcSrItat8zi
mtL1n8Ml7q7Pzc7wF5oJAZgnvu0ZhWOVSccuJf538W6qDrB4AQ5MKSA9Zeh3
effAmQ38uVXZCEV96NgvSi2r5V01bNd9qcpHBU31ncXYydXlyDwpmrDXysRP
J4a3k3NN7mr8pMYKULptizM/PZ9Am0uwb6JDDdzFe2i9BJiNQPj4CrOrFQql
leFZ2JBqhh3YMwhwNRkyHUREDrV9Bg7dCD2KpJHm5CG3AmxZMPVrkX9905jH
9QokY4twcQaJHbhAGfEF/NxAJm4bntCZo9rogsMLA9rBZ6laO+BcilcT8tbW
3Ag9pvn7dReKNffZbhf8kQZRIEFZMo9OeB5JNXUTh4qVL+I9Axl4uRkpG2lo
EWENJKQgHjR09I8dhrp16M7qRrGRj00MdaSbOpESFC0PnZNzN6MRCX48NZH7
N0kDeScJrUQv3T4y8qLC/bJx76Dnok5XxjaeTyjxHvcbY55zjPaRVmxU+B4O
18a40F1zh55hSEiqX9FBNo82DHmvSmO7c3NA0JVawDO2xaE41+u8E/4wMOSO
tck4kh/4gyjYmlXifAAcnWLQZOgQb9JwbOgKaviRacsfbM7Aof7BYkRGnslV
PPxMcaMoGt61jVO++pidj+jago8+Mgab39CBCrBDApw3Md04DejNw1fcQcwy
MjaydpfwQ2GVDFk0jYDJ6F7+74N0CIT7OYYiw+B67RSEcrZXYTP49W6RXUew
uYL5lSXkWf76fC6UNITKI2mH+yIw3WUJksMvYuFNKvpZjTqWurr2KN2hcIe1
bDfk1sGdn1unalU/H+kIzeJiWYTuGwISTkIjbiwDpSrWOZMv4Zcw/kAtt25B
zXPb2tRZS2DT9i+NlV06LVNE7ASEIld0i22p6KbFpSipBhr/L83CVbTh2OCk
377NPg7TuvXgZY/bC543SQbJf4Dw2www3IeIOg/SuHrkS3zlBkaGy8CxJ3Y/
LM2r3L9yC90ivGtkcI3NW42Z928AR2HYmmkOZpgSObVuxYMmqNEGPK1R9A6+
BIdWaTUfDmdpdhah+ooMw+nWoT11MzzvBj39qxnFmx1Iq7lClXemihzNTu6u
85O7aRABfIiSw5NndQh+fj2Dg9eRH7RB9ZzcPlNMQthm4hJfFx+E1Eisfjx1
guxC5pchYb7za8qoBcOJCj/s7h8N2fbYQhtCzbeaKgbMKnnzbbVBV+PpfHoa
MpJJFt7ela2iikg0FeXqEzQizrLzwcOq74Xr8BwRnE/XEP1eU+mnq9ECiQbY
b6uNO93OEeEDCGW3ZLxGfIbjmvhhFvgEfiu1r3AGnkDIN9vtb3zQBwYoXHNx
6UMY28HYeYEf2h6NShZLhWfUNFbVhFSWRaO5WTtkIc8+qnUsCxGH8AX/2Kzi
ta7aHsSMaZsWHnRLcgAKhc3UlKyo0cAlXXOcvqh83fYXXWLe2W5tXwFJSSbR
f/W9PjPlyJKPLITHPCxCLvqv+EmXQgFtqxFlRKxctfYENNohQng7ZeJO8svA
7YfOSNZQZIa+v0r/Jk9+bmT34uIx4kfsRBh47iXEVA7A48h5ADrdEogQAltD
c9+z8lhtZDy2OwSftUuB5ssjwm8KLZJJEeRBGAxYYMbIh81FElRnVAzZhlcw
HmcIDtkAXTaSSel6ecr5LsWBsWbGfI1DMQ2XO2kfXP6H8pctV43tq8yf1Gd3
Jox0H57168T4jMXZ1W+nLw5aZJCBjd+QDyo9UNid2DMXsC2hmz+QmzkIuU3+
ni/cNJgTW1k6bSeFLu+w0CSYqldmzFZma8oVSOPnZnRTRI1C0J7domj4Zwz2
q47aRWyLY8S2nhMld1OU0KK90ct7bMif6YJ2izFHpMh1Lgk7k8FhlV3YRwXD
bApV0M8Q3o7BJfaNOYhtWtRMQhte+u1A5ilXufJR3s0/NEA2oUacOujxD30F
6XholQK0ZcwFlROiJ3V6avkvYgwHgqqPQ+rK3ouEGv6J+LlAx4grvETPzsbP
4c7kPNlcDG4nUdAaj7nnpi4ACleIrqtIud+LoFow8y7reTAnScYOVOXbCtbG
/pMUBhY8qbRi92ptTzy6kGR+8ma1B/tRb6R63P7Hil+bC5qVTzlaZ2x/PFis
PbK1sYu1UPt68iCxVk80mYWQbObpeTsh/90gnOE0tUNIQOzqHa3UEtwVR5Er
NGgfRtdHRVHIt8JKVkncJ7tLrMDWRUYdlKSTl/WVIOGWvXUG2doDyzZ3ifDR
ZxZyNC10bVKks7OODJ5jWHyBVh/kq9hcnW4ZE+OUFrxUPRnBg+YRIqA3AMhW
gxkI/n+EeG9YK5gYPVSF56OK1+Yj1oP/bBEBuAL7OmGrFlFq8Or6zxoUznDH
oGk4m8l4mUjgUP/JnQ9c4Pxs8DbK8BO+KYnIV8dunGDaK5TJvAy2xPOHoIQZ
NzsEwxuRu7nA+5R/+0tjDDptpzit7gJbp4kp4ChqWnhwdDwrk5vXjVxI8JA8
4fDkuJvn4VhALFbfm80VJQZXwRXdfp/TPr/9EhfeptepJDyLSGojjGeA0QIg
Y6grWLghRuDtLCOZsMXZRxcLtYSdmnxx0uz/SlZDCxWU4r6JTQcR0AF2bdid
Mkm2PZviFXadK5CJy3GGdYaWfn301yTmR4JcT9PnDktHWxA9PJ9zqw0c6HuX
PqyS/0Ros4K+TYYdK1LZoiIZ4Dpj93HkAUr4kMQq1CxdtC/LD7zOsBZJkCMY
7ZVjslq+Zcd04EI0s7Epjx98LiTG1YBj9g95YhrCzK5c9HHtohzNbAxLCMYr
V/jZnbGlu5oYITsGbd7w2jSSqwouXDhOX4F6az7Umpbzto5oCv5ru+xehawZ
dCL8vm09HSSs6DVlA1EL97VZPH2yg7uWu24/awNpAfFQqBNIh1bDmMkprwI4
I6EE+pjifT1VNNf2U5Xr2z18pzD4Z6zp5Pxfll4/6qT/EraKuiRi/Y2GhFQP
ozpRIY3ZyUK0UgHO3iPVdxkiEjt4P4oYstBMR3QS/oLVS2dxH4tp1+8jSGf1
J0y2Vf14vkiy6ES9NPHEu9nvOUJrCxiIGb7vlD+lyrnlFI9lPszqq8IxJ29U
hD3vu2cOaD6M3Z3Lp5uRQ1TuVSjGWkPLCDGrDZxAGGJZK0L15FolR1XOwcKl
mB+imb5y+RAy2uiCf/p0Y6nEYCJYbxmh867N6ddpO/besWctctQThA4pbO/U
GbWhOhQzBwBB/ouepzYmA5M3E/HfcjlJOst/M8HGYANICzOgiicyzFWmbnHh
ZylDpTIWwPye4KCubJlhq87D7MO+RRSOge41vbpErxCOTAN6ntuasH5dCtIX
R9LUggoqRxuxiZ2SE0q9DKOsHWPCY+6u2UQuSMb8UDC2TbLxk4P+iU/hsIKr
RVat10btQqmhxiqnbs0pp/qPtUoG8zUo82iPpTltT3cYHkmXtmsyeD4HzkuQ
oaKDCzwNEDRdi3/bw5XTwXjmX5V+LG6W1+H/3JzEF14LoQhJOA+kPXl49/yG
reKD1nNaZ7DHmel9cvYZK0B3CcyzPrMCtD7RUFL12TQpAE7fLXPdnEWFEQAz
xWLjeejjdItw9MXkG6puSIzfk0BPpitPOCddLXer/tyE1Aq8Nco1yDkJHkvO
0H22M/TOdmUhfG1gWT1/0jgN5BJw0TeMvsogSeAJs+SjqlApSihgYjVQW+bN
tzcjeBteVfUR4wfww3HxbtuZJ3cv0heX3mcgv2eH6usO5mKqwtNRWqH0tsyE
K23UjsK4GKWE2Nr8xVoRRYbgMixXzCuloItLu6dtNlu36OnmT+5IRobVyrIh
wx2MerdnV8Kt8LdZS34cQ0ptAXA0NOdYwLBFZMf3eA9jpBjq9pNRUjrgD4Ro
9VGDnHI8RB0wZkHdUEn7kzmLpjNugB6hvorE+RJG+yfI4Gi+mrBI3KrNCF8i
fyRAfSqj268yRYGiQVPd9jco0aumzlmv1lgEWYCRVFK2UF6Iu/SLNOwHew9b
R2LV1kU2sznykw1GVJufgyNcgMPkgBTCjRSu5j6UTiwmQtJ5gu+xNWmbmKXb
Y1uQglL4ffNpX1RC3lSK+Un3WhPKQ2NUGLDeehoqYXFUmsFiInYQEwTyPMs8
ubfB9U+YtasOdlDr6d6rXvEV4db7cKYQMKZepWxbF/vTka165ejMVnVnuShw
oF3KAfdLumFLq4Psztg7TbrLrpfIjzSpehgg7kgnTsVxYWNc5KP3eYLCwWre
9FySeIScE8ftZoCKyDx86SgiU/IBn4zisYwjOzs3eKOkvHkKAK9IdKZHHgVq
099CNYoXj2kkK3dxuST+DQMhFBsfj1zoBe0sEBBkQcTx64tvPBtvAkhGfsw3
jFvwqNtzbvG91MQvgCIL5aJuskDm0MMWet/XjfS3A//n1Tk3djeSvVJjGl/c
QN++GwSnyvc6Xipzc2ub3ko5DHsYpyehg06VYiLEmjmPNhxxJ8qReSQpdke+
AHZ1NY4T06q+p7lrngGe14WqwZzE0SLYKYSnTp3mLGhDL+Lc6cjJ7oa3xDQf
dsgorMPrST0QlFUBtfnBiKT5AWB/SNfHghHdV3uctmT+ctOHY+uTWkojgmlA
AtFU2BNXEutYSxDuMt4umbVmZ44LADmhl8HIuu9ar3N48oouRng/0tEvuTUG
X3xueCqCvG2qM3imwM4G/kFPCSpebfDiStd6K07rGVGIDgCv5eiadU3DkoIu
sEcNANFo2exMphbFmq+3IQBIpxsCVVt8MU3wwHQpq0lHGJgCVhgJHTZsH8mb
2hA5z1QkjOJ/nBvZ1vgcJ0Fb0ZmNmrE1eIOS+Y5xDVb1sUFow+WdyE3thZ0M
pXi3RUotxUF9/9w8SBTU4WW4A2bg56XowuTJVSetu6wFsLe7KuEgUFG2cTIU
Y+YUVjHrtNfEeDfwWRwvMSFMBd9dmpYP4r1UW8G1oEw91kWQTJTVdpyq8hQW
ZS/XH4JhqgY6xrOVIOwt5m0Ruj1cPjUIWn14MPpNa3/kWd8iRTyKAvzPQarr
RFp2CxgxFT9HikdnUEGTjtWTmcy4xihqTFfNXABxPPEbrIl8PuP7mJwe1yCd
J4rRaJhPAFMm7CDj2t4221hOZ1eBWCfgzkfJ5DM5Ax2Cp9D6WxB7QKia8yZJ
RLvoxqe3iBcOWgXl6XicOtVFBDYOjAsS0SKAg457J1y+7l3MP8Ax2NzGnMxL
Ijoom5007wnSu7aH6HDZxLTmycNKf3j2LTPEV0aZo+mlf66asf+aJ3frEgPF
z87ePutu2xj2YA3gtzxt+4SpBYTEjdTe6fOtPbYkhDJOddT4eDVJEiJ+ECOV
AjMrjRh0Lx7EAgYU/4kZn2HRDdCws2L2nKC+ybBLcrUnnvbAGM5upAr8SbDm
h8xTKLeIHL2BYBghAJnNOZTR4Pu9VbAATZ+fr+gLW807W/xn8PNYaD04zbvl
s9mRqkzO35ea+RF6s9xZm29T/nSsp8YvpVmoQ4N5HC8i9z44jsDt5Ukzhxd2
rA16hmHn79+8+0SPv7U4KnFbJKnvIo/o/RWFZ5dOO0uBswZSSiovOn2zDH46
+2/MvbL9dwgdsDxkAbC5n+pPJHx92SGiRjtHTRbJ+bX/EPNtgbj/OKbaPQYo
kJSd/h13qU+CRmI+b7KA9x7oM0J6PWpvdQTJl5z5qKrcE66HwXKBtweLKqNz
A5hBEMM9D1dAJdvtMrcPu2RZ4RyktPNcofmEZqMWqmt+xZTqOCh0qxwJ3vhp
5R1gUjv8MIpSCevvkHcKSkWlvyAZNSIxMkC9HfAUfA8IiBtM1vrxL9DXOhbn
Gk3aEsyUCD3Hx1lYuBtbOztWFYm4Lqw/QukrbcjWXEsRJGL23ZGHaKvSnVr9
itsv1YewmStS5RqB/6b3Cagsar69TCQxaD36IT9nAIhtAJWIgOKBeC/YjXL1
PyEddmcNANelKN7YHZV1wLv/ub76qqaXzMGA+tWy9UbABFbDG+RfWSttLRc4
s88O6nJdtzqtvwYgFk+WWzDWygNsTvm927DZT3GXszshIvqgYRDdUC0a9eYK
WxE4+4xW4SVvotbiu+Qwl2U1WoSBkO57Y3PAGy8QexiYBzKPInFbHxsb/MUF
fyRbJbPil/NkkegYfoiswEj/fNDVaWE/1U5B2RP20/h+GkVK+M0sFkpconbx
+Q5ZSFUKxPhGT91I5mT2HprQaFvyTFs68Keq2kGeBbvNrx9zMXFn6OvoBtM+
Pm8wjEQDOZPH4pBIBPjL6TL8XNt86ka4gMotWk6xzGigTCaHYS+10FhZGKuP
7USJaDleB9KqWmhAl/IBS66elfUEXO3BMxzRA5hM5jRewXMDmmYXrXi9Qpqq
PfkcbhMrza89nbj2DfQJpUu1QLlBV9wPxNdsx0G8CAybfNWS2zMZoBTw9bJA
e2W3peg5XGRN+qTVySv7EQREfLrDwXbSKC0vCPWp/8PCIvyxT5P2+bNNYB1C
mu6JZxGkiNYgLO+w+fSQ6Bdp0fZvv5g5yngjomKEFOB76nJIdmFZ/1LFaeo8
+S6zAazBpyLyGoKf6UUv7bBUT9Bw7rxa4nNPI0vSVZkdk7Yq7GiXF5cleJdo
1JZ4evhh4Y+h10VVzu+gPDteWa1zFv84IMWV9uDPyF+XLdUPsY1PHFdXdTqZ
0B9THVEZG+ge4ZQxS6dZ9ECl8VZmhQ5YcD4ftbFTI0K7wfO4e7He0nvomASG
UlVQcUTdN/FMVyqTPsmScik//6F9sgvh/LbPGf+udPjGRW5BTBztG+rwahT+
PRGEu9qaw823ETK+uAGEBVI7KhKTI1e/ca+R+hAZxBCQ+6jzq3DEGCNepl45
tNpJBEollQJpW2rkf+kceeXCF3H2IfVDEYcfRk2wV/19FMu4jhTQSAzZ1kEb
aYaYpxUqYsFWYsWaJxaFlcs0NG55mpFdb1gWCdeb+ueluCoIudCazLntIASj
IioIR1r8lwqs8SFy0OsEvpvi+u0uyfrhSyJLWnYH3+1EsYRqI07r6BnSrPS0
lO7G12Z1bu4cTQMjScF3d/rG0XRSXYavpPO1pxVgbFqHc3fLU9W32Vz8Gl4h
n4ByFGiCHlM+y0Mpcjk+t6W4+t08OPJRLxVjtGtePsUVj/XndsxQ5K6jbErW
ilbwMBzjgqQccD8qca11Q/ntwV5IYJtHHjXwpM62S6/UFTB/F+k9mZjcn64z
tYQ9IdYWg7iJLBzFUt0xwtEq2VTImfDzl6YJieI3kXHDNN5Nnaahj3pnO6XK
qKMP5vBWCwzD6OS8N9T8i6JPtq2By/7K3uqrHLM6vw2G3uIiHAc/zC0x/xAb
smesPiII86sCXFmNNMS/Vu7Muh88//SD0gmkkaAD1zgX/vr9BBaqYllrQ7tN
4icKDpgnTE0w3Y3hXoAxxalY227bU/heaZK6vuDH5z/iZuZPK8y6NaCtjZrR
FIyNxkqc1xNGyhjOw/tZB+XJK3179oTam8QpZ2YL4n0D57RUUDEICrX8WoFw
CEPGk2mOX64egTcxjLOa8nzC9h81KOCpvQBsI6EFYiBk8/rQt9k+0vkCo9a+
ijul/AIK6wKeN2YHO2ygRgtgVfJrUYsw7/iMMjhNpCBtBpEM4ebSDoP7v3X/
DP8Koyu2MDZeh6fiyVTqv/ERIrZjkAcNIPJp2cAO2WBeZTrTWi0k1J8yr572
n/uzEqNU49QZsixT944zr2SHOV5y+3knbZ/Kc8Aksz+V0ALgVOH6HF++lQYt
WGe29KdqGfk/zkwPSyNLVA4NfCgdWsBxenv8to+GpDqU3vwbgKVGnpRnjRID
Dke0WflCyRwlA1BTRe4duN1Xr/sTur8JHIVJIZevNOW07wYNuwl04ZhO+n6W
cQLRiRjaNs0y6k+azYFe0uHsd5LSjhfGiWyyap86givLoARMRzS1ukdTVjKy
2UMeHz2mCkVTIFxuH8QZNpqhpgbejNd2MNKY+552KsiQ+Ztbzr57LUJbGuof
LRbcQJ2pysioz2eeVnrAezG9AZmI4jztJ595b9VToA4aykrAO5DaC2GI1Dwo
SK22nImVMqZkXoOd6Qu1zUWvWi+7IMLxbxlFAbpA7XotQAs1Ub/Ut/JrAFej
ynOYlwW381SNdkCY/tAhEluizgWy9pVCGuTK8yXFzXQlZH2lCO0TOM8MJ7+a
7h7yc774JKbECUc6p934CKpXFS1zFsNL0kwPEXzOA8lJFU30lB2b4x+HPYGD
DAiJH3kJ+VLWg9XhTde8Uj+VL7sEZJZykUr1xMM8/QBHTnweTYfB7a1cjIKJ
2Y8wWFed+v/coPIFDbNA5czbaWJL7GqxNVxjHVYX1QfddC2AYDpChvjG0x9K
94mlHtwLpw+tzDDNiRGk+CjXJ2OjHQiCkcwJji7aoD7M+YyKBO6IDkl1duGU
29irXvHaIu3CAmjSgnVZo3MdHvmuKEkks/zi00Hdg0WjKJ/HL9wQ3EZpS9tc
WFuNfl6VGfyFuStp4D0nysmUn0t9YUVcyrxJ3fRTtSpw30127xuwPXPelYLG
YqJKd1iz496CQiSO541NBHdbyNXQD4Ml2/F/EKWnpCDGomi+DgK4+ONOy8PU
p1yLM3op5euEasVRiJaZYYpT6qsqCxAOJsOhCEL+UyKpjvlX2h0zbuC4WY4L
Rtf0NrrtPldeZaBDKDP/Toe/4cmop+noUF8wZlvedTfT4C1jfL8olr7QkVuE
deRLyop5PMim9f0DXfqRubVqxNvfOf6ocUml296uQvNN3RUoiE3boIFufkjs
REZiSKR5lnVhrMcxk/K2/S/sVMVaS24aUpWRU3y8K6Ld86s3esQw+67qyiXP
u8Jw5jGhpsYWsQ1LgHv7bgkrC11Pp871iF7tNDq9+H4pqqTDItrdzCriE0eB
lQR1kU8aewV7Bt4/3kqyTO7x6i2fXOxQdyCoCPhyLjhtWcOK9RrNghYjH7Ht
CqOTh5+YDHMbUKRxLlMlwoqlnuRhrsBYTlD/xwISXQm45RQCQuDCH+4PhsCK
ZSekFS+muvj9bSpwbwDuuy5R/My68nPVj2tN0Weag3/soIKFlneTLs2MQfs/
hg8sB4mmBY0LIvu3GWFEi65DKYTNa2BD0gs/W5OE42EtHuBYUxNS7mwG/aMZ
8R4IajAmHnXrwG6Dv0DFIbyxwlgKiE9ViiZskOSRGJJZo99TVUqBLJXAZf+1
Ri44ppRzxfyN5hcK6hrQahLd91z5+UsuFzUWQ3WIYiqxZB96pVTzj6D2zdso
umZ+iqBuIzJ+rprOSSvLI2tVtW77F0gr4JcngOccliBp0/iqdtGCWy1hxRdH
OCDC/Yvlk/XZ/d47k3n/UpJVoShubfhS0P6MaL8Wc+BcHLPEYHWGTTdqvdic
m8M51sjfjXqDPSZbJTN9vjhIjZWV/vwWaP2HI1dzDfU1TFCh4gxO/a6GTkAZ
EW6THD6t5f+HY8oAgIVOtlLMp5olDcUg2ZEBdJFmsmR4hkn44Xdg252qQQpy
sRndnefw0I5PMLoIaHGV3+cSXN1vylDHj+eNF5GnMqdMksBFHprK0yM6B/Ul
sN1bYUPlODx9vT/oD7J8IBTG9Xf4QUZ7kJxjM56OdjqcWbi7XUkJ8Nu0F0C6
d4Nxie+h9tBvnb5fprYYemsV9uOUsQQE09CaHOJ32wP+QoZjQ9RI087w9MAP
UDod1Ol0pYsF6puz7aqb8ZKeUJY+9+eNwhjUXO0lUHVfTqdAqM9y6CRs+0dm
SITgWg7XTLs+NA9iKOOBMPZ5qB3y7nT9DU7XuDY5O0UsppfZKciUCUpngzT4
fDSkHpwJcDY4t5o6oTG1YsPTGk235j2byucDT897Ne3quukaTDBWjOBGnI22
zXajBXk5B6taWxP8/natAArk9fCl/HbxxSDEEKEQ+aRmy6mU2oR9I3M3miH9
jwQP5M/BpX79S56lamM70K9BnFkk/c6/GcqTHrdv2AsiQkj4s+zfBJXqmdta
ywN+0QLm/f4XSk7JiMWFeovwVeONQiRRGSjsRsnFnYQUYtXH0cJwA9UEVLhw
8RdPss6kt1zbPCk8u52FWr9gS/nP+ud6GoCsX24qNzDREsIb5lEm3X26n/Xa
lYMzC9OKzGd5FRF5Sf+l93ezioE3WO3LyBOBHG8IRTv/rmGufQoWr6/OJ95u
UCZirzGZe+xej5xDvwmlaTbsZQdnyu+hsd3hjf3PiO43lYRak4O1K83tIgse
gs4tWbZBZ3/eTWNa+NKcIsrXqpcJHAJUvTRYOmR2kJPtNhKkdMOMzXMFqgTa
ApGMWHusAs+DjyGXaWmPNlYxmsKAAj8gAtMPVz5pxOopfvoZKEyRT82vdW66
JZa9HgMp11n3v2KD8el++OZlTy6THI3MqM0G7oMDSBR0SCdcdVTq9NYPlky6
XjIqcQ1OGEpQzazDBoAFWiC3V/UAqQMCCwyUdCS49JlBbhhtcCM8Yi2bRVgW
Otba5UbGbEdk4mZWsB++u55T+1RYr17nS/qV77MCarHhLOspLNgrV/j7EgL/
gYgDOep1E9LX/HHb32ABz4lymAOpqV6VX68m0intAsCM6GioSQ2bF4blPvoM
RUXvrR1FRrXvO5ngnCbqoWxzlGAaA/kou1P/3yl2Wgm6Dr/MDOWS6ZlhhIT7
sERm8gyrjyYYbopcLQsniSN0hk1Nn91ya2kt58S/fLOLtXNU6VHygsXMNZSh
yrOro2fPaWHqzjdaijM4mrtB/8zfFr7HvSm6TjpcaAQSdEBO/cFRrSrqx62m
l2PHxZyteDue2ubWCYDntFGN/WV9RGHON8Fi7navjhp+8O4T5mtfIHXDNJRj
86JT2ybNSri5sfXgVungXIy7dgenhj5xkwD7WduOysDkq7cUZlGOrMiucL5A
Vlw+T2LrV3Jkll8JKBi8qtuD68396Q9ZKGsYo+2AzhfgpaD/xiHerTunrKbj
Yz3Arhu3x2UoAa9hK+sWgsf1jQPn5h03/ZmSXyaL2LSbz+/f9pBVhHgMAFCj
sCOf0o1YEUfmXE3qAhWy4rfemfw9sCdLxV6NgFvB7Qs0FApF0+gDfl+FE7N6
sVQxMryyTFZCsweRKlfEmgUdA+psfV2tB3+xF7duwERGDeGTOgIdbcuzSSVn
GVb9+AoEqKbWLf44ZL6OAYFRvwVBXHNS3Y3BFZ+za/UUvU6tDsq1CCwAGz+m
8x9ZsijF0yc6BEfyfSqdsxrjR8YdI2UssEatoJgbPsJPvnyrzBB1mxhXiuKK
ChxTfPpyc10yy2qF0UIsEXoO07OnbAnrWxJ/Ua/yUt47qMo3Wz4LGWTuvGx8
njXugmOwqqx9yGGx3hMpSDdFsV7JygLBQctKJzHKtt+DRn41rGCJaHNzZ5tJ
BYO8t4hQ7K2Ag0sFApeFi7OqOz599PyAkl0buYVC4I9uFiFQyUqpCwdkSHlg
99XSZdKZhLiu2idv8iTUyHDBhuTIWMwFm1SWqUIAJgF/TZmzqGndEf4TbyWq
1SJ8wHrSs7398cabPwHkD4hb9k8DGDHd3HMdaqoHLWrab6HJzo/kukU2rIFT
ZhyOvrux4u2NJ+4kSF5nZ3dL3TwAd1kbt0ncMNcWAyJ+vk0Ba++MT3qhEwM6
m+c+fPocwETsbAztOMbZio48QfNLTGRAKq8UDYLidmj9NvD2AIKXbBRk3jk8
QsNq75lWPT4hd+lcQ6wEgZcHyqfyTOtA3MzOu267p/d1LGZCGrNbx+rKr5nz
yJ+ZGrmrrOzpLDfeGK8568QomXyO75VJi/JEZtM6dVXQbIeflJ6RDsdFsfuF
JEBKrz2YT2KTVSTXa9qYNPSLdy2HHGXIpSZt7JMq5KcqyRYsdPMVAhfG3OHh
npnLXL+WLC9N9aA0SCjNLZpAtO7TI87FlEbplohONWGyz3bE9mRieQGIMdcL
rs/7TUop/w+X+JchLfTaRAy/YGEKZ6V2qIz7+FT4fKu7YLv5VjHbdd1ajo91
5xmTiD5jJW0si0b3SubRVlnQqdhlOwPj67CHzHN/6sGWLtaxFvqmY/zFin82
Vt0AZ2X3V7Td7A17WQ5kDM/F1MW2H53sl26x/CQgOt6Oph3w8h6vA9/0FfNx
oCNOwPCeEsp0zU34hdbR4/McJz7CNjDIsopTFU3hyT+isizS7UvvV9ksnMjG
Tl4/qX9oHu5xN96mVmy30s5UtKhUwStOYbTHWxFuUpTHuFIA0HxN6qUoGNbk
w0X3Sg8mFCDJ1+9OB83IAZDnI42OuhEH4WFQWaNrhfCxsJxEWQ2CwFGyehzR
IvtS4uFA3yrg94DM5cH6T9Pd8eeo7DAV4If5fJjhjdvnzU5rMowk0DGuMj6j
604pgIpyDckDiLASjmREIFlAm3a007fcsSh7UHo1riq1yqfoU0RpnDP/Ifv1
CGHABieaTEVcDNADmWnXPuSVSXC2/zn9IG1R4ReeyhEPvvP9joBcTSKDZQGg
JVNKNQDODNFBk1P+hd4vCmLeVNVS53/Zu3YkFXh+7WuqjKAl8AHwC4CaWRM+
L7arvUUTy9OXWLT8T6FVyMm39ECpbT92gFBQto0WkvY8rMVfOvFZR8nDr9Zp
xtH7d7mR8qPwcZW2ZBn0GEHP89EJaX9pGyA3Z3h2maG1BUmTpVHmJwOa7J7o
IQEBTDtT/LHMDfXUXnO8N2YMn+dfx9GVQCuIH8fFHyZYHTrfXARpDhY5OzqN
Cezpy2ZP42uaZ6G3cgxXtoPXQcW1gbmJmLFjRIbMynoUkort5otVcBo3CVmN
PGBYSRRN6/4wa6hLsy2myKQfSSeQYT8l70DcdY32wUpVPyavlKEEpmhejS8G
Tl2G8cPyxQNb+iRBjCY9iyWw7Iqo8G6HFI/DfUCrO4Xq+4UkhctOBSmMM5f3
ec133Ynd7SF0KJd7eMTY4qottW48PuLt7OYI/ZK+14+sT66xIz9upLwU6bDu
+7kqKpkkDlRGlezy4IvU/vlvrosJtNu9wE2CrwSb0Jz29pfW0f6tpIfH3X7m
GjY0gh3GZ/Y62/9CJqQ26xP6IDiOjlWIpE5tRd2BguZb3U7U9tJMBrsTLeMx
7gTREzVWRlW/xCLETsrKSSe9/QnY/f6lRGNDlEwtqMRFSdnnT2o9lTDMU6dz
4WelQv5wFO2vEW0A8YfyF7+bjeoYJfjrEHGC3o6i8oiIO8CaaxMfMbExZi6B
yUY2dHgenhe0IS9cKIf9G0LKHeGtnnTyAbmoe9W395H9Nf6xwH5aDPmLY5+N
I2YPZIbUzTh0cM/5ydXVkgA5NwP+2/FUZSP8YsL1tx+TTPUrVumVDJPu+mi6
sJny4trveiXCl2viflSS+8rwP0SNXCQPNkPZpWLKq9rncuXKOWPIAxg9lxFX
Fty/EHJUI9K4P0fPbLXlaaWzKxbZQYWOCW5hzkwzwbJs0sL/PyiCeRuO7AER
Bt+iJrqNMIe1U1orc1yA37iGA7+074lTJmmBRGolDdRHMPc12+lHDQ52ntKT
gkD/fEtL8tno274rL7A9R01hKz9mfl5C7QsVAFWUNjPToEEgJ3tvtcRBnSeW
v+DD1M9a/L0xJ9E77YlmLsgs7D02eJKrmbCifaS6IUNU3U6whP+ahGY/B6Sb
CIBNFcEYCpzDswZ01zhM+UaqnGnygNs6qnhn5SGpdI071jYTtIo3gw4CDRTB
V/MFRDqTM4QB1dWfT1ppNJEUfPdHq/Co3p7pss9JrkeoEEZK4CM4pSnFxSuI
f3U+mRuwunSsQua01Y6FOfR/heuzCjYlEx8PwfbeTM7eR/VvwV52beHo0Ssp
HtH192KomEFFo+JOU8eLBRLYlxAUYMKlu2LyvGEi4Hh7TnmDpnKm8rIm/JXj
Ch+nkKV6sLKYw4RnHfaCz5gDJvy8/ITtI36cJyjP9yFtaPjL5gjM866e2wIZ
x48237AzCACMtliJXcOIoKEe0Pu7nZZfS+vExi7BRxGcDIC41W0/NMtkFeIx
OVkzoIk6So9rt1pP/bSIahqOwsRkhwSv858YDYvxmDFZVMc6uPlwkHJ8BPEl
wC0OpxfinIsO+WF+BOYUash9SRR2nZBI6uu/BhJGlmK6CB2xFSQ7cVI1/OM1
L1363XTwcGSiC+hM4hWA5zEY14UxnYrb9Lj3KsGSw+DbhDRya3gFUWMJoIub
e4/cOpXwZTBTTPC2pwRLRNgNpSljh6jFjlKY9PLZ+Bd7fopXtFH2OvCSt+Ja
rLSADjUO1QpLJW/ctyFewkX1+NBnUdBCqWQiJSn3AzoagOMA26lw87mklqzH
Jn5lW7PWvac0MXV3tRR3TFmdMwePe89Ahy5AFJBSle4hL3JOD9gwtoxK3dWl
cx99vJ0QDwYMN8+1KqKdwItUxTYuRoy/lBvGJ/VPkHr8NmkS5yKOQ9C4Q8ff
9wRUawttoHlSaQWy2QIkjhI1SUS5nP413qm32TD38GwXkaw1evlH/WVyGipq
DWDozB4ItGt8CmMTV7q22B2x2+jzBWB4SZ8f16x/GCESPJuddOXBlQ2wxtYg
H3e1CQdkdEM9YbvE+NCfjuv0vEzk0hIGqX4EIQ9oHS7R5Y7aOfCh0B4ZYA7U
GHJTzccUHene5dt/uWYZdO//WgdQwheoO9I0nHAHDtIqnMJOYqlXAGT9BJfL
fDRfbD1gnP8RgAw+SBX4+TCXWYhTTY95gtemo79/lj/2TI7b6bUe3WhcVtDO
pmrWCRh35JSqyHsoPDzkIB9G2cErm/MqllphxQ2NCt1Y9U8/fn8GO9XDrMTc
2c89cyjiQnbpneU4rsVzJyy1jKfHOHL017geuFYBRFuJjkKwT23pnctC8ykc
iaH3ErJqEtgUznLbRphtff/gZp6Tr+wXbI2F5ynrW4Vd9h0q8nB9Mc27DjvU
BTRziIO4ZA0Ov6p+9dcY3SN/6M77LVFbF55VleKkivl7cXu6r7KmWspW2Jp7
G1yRCK5vYsK2vDRE+9gVxECO5LfWmAHT/ESQ24GcM9yFbO9Q79pdpsOJPRHN
L2wk72ZsALgXf37m/dvrV3k7IrG/hFaqhkYaD9dtO9/efbslej4L6dCm8U64
oa/40B46iCf+aTcfAmK+BkEFTbaRMuZwmFFVSmJH/H+LdupgsoN8pvv4T+d8
ErStVXLcP/553NqY6AHwVS2zi1SXlpAthrpJH8/CZfMC1aaldIECFIw/881g
yJVPTfgcGe0BZWOctw2EEX/524ejcNdrBXF9LbbVQkAgjjBsAhXN8q9+2SBv
n9aXN0otovjMWEjv7uVgU17Cj75whTyZ3+YA0wioQ76vFEihn5c7/JJmg+qG
TqPch/fuAbov9il+EJPiz5PpZSfP3rNH/lueOSzHXByLQJ2ekYIxkBgbnV+a
lvvpdOyE7WBFBhovL+Vr56R02fF47Lh9uUx+taG4WdHCcuRhTKTk1XQLepL1
OvJD4YjgduvNXDZ2mk3QOH+zKi2IMWsSdaQaqQ26Y+6f7YitcXeDXiuMzPCW
nQMruGmdEpQM49X0DA+dcsf1rGzlH/8xGLvU3gCJPtgEu+nVzD7lRQ8MlVdl
UVklCoGfrbHI8Gkl3wNEved7V7G4elbHv3RCizK0nwFbnKR0Y+5Zh88MKeJP
W7Lg10GCn9bfRP5JFiV+oXbUPrpok+P/4nh8ahoJMf/cTYQwYkZIZnWjTEW9
kSukJsN4JKVMHkGW5JXhUwnwzgOGuNiJUWClNYYromWgbezQ/RV9V+ZtPDZA
m9HSxc7DXki+/ewhGXv2yc6u3yobSQctzt2StW0NK8lpAcE8hKJjrXS5tPOp
IedZg95kTkpBFiitew4kBP7x1bECFm8TMQBjP8XsrDiW3U6G6dDILTIYzgZL
powGeFKIrDLYg2hmYU9nscKQ9nVKFeXrRaJbyQ16KZwy+M0oM8l6wXhhjhdX
ylO3Nc72yMEkT1M4nC7MHFK6LH/kXmI/f8GOfP9+y4CfNqkewSDyrsV13vlV
JmZwE0sIxNXvu04Qf2LSKcF3prWzV6xq0DEZMx/kgMMIIwM+wO+JPFe4odAd
NPm4WNcBxV+Xcudo/N1EKdloUaTimKchX6k4PM3CaIEsQ0/bAyGUOnKoiu6q
WuUyqegNrZrNP4KjzM40mNObWZjS00GFLEYxOiR9qp6o60hbU5Xm1nrZPDwc
0/52M4fHFTuLs3T+JzOWlfK7unqnWpfWGSajHopA1B7tMy9IvlKcZbSBxVpE
BwrNfPb34k1JO5ymELIqA7qVDZ9C46Q2bIFSXXYsY+aFuuKq6FSoy7BucPY+
+DNzE7EoVjVgytWA0n2oparXfAaXoAC6FgQqlMoqZotXS18WVddOh3ABSNJ+
Tzmkv1ywzWJcdDGYtl4tlz2t4XK1YFTErPM5nQODH4MUnFvgFp9eyoMuY2jE
gHmZP0fO8uWQXIv25u/0YzNBB5sLk24+vHfeNXGYELMA/HICGwbdeyaUESjf
a9e0tQsG00QsoQYF7xR8Mq49WVGzHkkgyy2p154frJCNek51crQBQQt3ar3D
xV6NxsAm94QHR4foiP926AkMQH13R4jf1xSDQEOOQyZbQmSnpZbwlgetocZE
tj0wdaZpjr0oX0h2K3RFfQm5qv0kI7HQSJcSRjhSzBZ7cgUeJOUgbUs0GPv0
hkwRaPOfCZLfW5LapQ8qFsbA8r2WjKNUu2gaNglXLkML0cX/SAhNgQJVoQmB
nrD9vPjn5RdLYaGQthojLVpo1aFAVHjGD7SN0C0SNauDxl5MYolupD5lUvM+
ux5QbnngdsZ4i9pQR6pyeHplfdBIWOY5yLSWoXGpLzurR2k/g7lrfxkxg5ti
9/ojUh348tUDZUsk3/NJwYrvxZCwP5Wf55DOJNjPI8Ypb+1YUA/mM+ZG/jA/
vuTSYt7Valwhizybq3j+rpqEP/lqhI317yC7TIox0SQRMsNUkdTpAS9tmi2X
0BX1Jk74d/YjgLPcKYDHFeA/8Y+k4XVm4PZHNhCeVwQk1OJX7mA0uqXCSpJ5
oD/UzFo+WFIgKOnKN0X1yzK14gxa+Ug5fEdtWjWMctJ/2QAcxhWMbtgsMvMw
SiVyIHLuUiW+pkCS2NwVq5FbLenfxBTEy68avhvP+cj/Rb6t8EoCt79bwG1s
u8/OZ/r49Ve+oP9DiZlVmgG21z8aaE0ELh7DwwOsEvzGpYGSuHiqrV/0cD9y
dGmsA1oPBJy8Je+46HD9mzjoTbdoibHA7TDPkGXowi2aW4p9woiEFJWaGcSf
4HoXQkllRyQH1HloyhuuCo4ugAwxrG94sMXbzOk2ZhNdwIjT7uplVFF8MBXF
005DKJygvzR67lOsjSWzhVTUuZFlJn+9FPRo3T3Yf/x1YGHDbyIZzcsOCnDJ
y/sFArtwhklGc+o2iYx/V6moNEg+GvPEqxz1X57+WhDZM7jAf/enpHDuzYk4
edh9KJCUxi2gBpIU08D4+WFuZIfo5eayZW1d7yd97uZoX8KrYEdg0buC0QML
8RlUNHkPyw3EY4s3jZYsQoVHePxZQR6uxdTtIKr9+JK5RF0FgrppSvbZzYiF
0x/rjwgHmfOivho44vwFJXaYr+S4lXVLoFa0LCa2+lraOmrV+9rzMDxncObX
c7b136n6sMs0/9aggw5PSPEld/M2HMoxAiemzgWFwmz5v+fVoUGOF+icsf+0
au1dGgFwgOKIFqF23kHKH+sIdsuVxReB+V6UWqwSZWgspFV9Rfnl8PT3AJ7Q
vV9pVY/t/vKasgoQfID7QU8Atic3v6SHkZ9Rs5prRMaUOqo62FXHvcvgMYyL
29ALPY/dWI8J99grinZz9j7+PEAhkHga9MF3ao4AgInhVQIG7WtEnOwJqCCS
Hs2bybxNjX5F1q1Ad/BOs/5ZHKV1wmBZUvPkXNDUZGwckxTRVOfeIUN98J5D
WI99hRPNmqPtHZ6NbWTCMFHXcoNS74PCPwqSCk3tOMuJweVrHXLjqdUw8/mc
pvIdT0V67PniGCQMb5LNBtUDFGkjPxmg+tKtV4w17Eyt5QZ0Rr2NlDebT/HO
5k0X3fRNTqi5KOT5IVm1ADO/nEMw5hFhUq6nVQXVJ9knCmE47ReoZPUB4Khl
WS4oIQqTcEZo40BDDtAiDcSfEcVHUnyRUNxF+5K7n5j1TA1qjNdEKpuJGZTj
mhm9urVVhI6rBwszrUOYXfMguju6GdmyyJVgwVt5eACydJaj57IjjOLogl4p
FJvbsD4baSuq5nTSj+Fho/nRqOtRwGu7RrjFJvPQeBdSB0/BSAQcZ0iXepF6
XXAeHyl3pqNKvUX0LQ04TcBujz/TB2Dz1euLEzIi8/dr4xFQrnYhKSxGvMhc
tCPxj0fDvB/FD3qvTZqrclkiNDHaWRtOgqAJDBAj31MLuDWOQ9mLTf6R4iJw
lAsS1LRV/innOmiWVIwp37EX6lw0PzDEHf90AMVOMVYqtDq4uVaVcHOwv5ju
AQ2Vo+GjlWIB+gPHCjVYVBS85VjotfzxDwKqqJEgupw4fE8HqEoLZ1/K73Ng
BCx8NTT5RLdaDU1X6UIf+8c5TVkhV1XeRiL6k/0irRlstNT3+vKPQeagwrwW
nTxdUUw129+8wAC2ek+FuBTv9Ayv5TMpdVYWa8dathAFFJM1jNRzv3cQ+tqj
6HKSyLbtn9c7kI+euh7mGDDlOfPAtbs/hZBp163lsFTDZ4kA4FYzlQcUwJyx
bEl1Q1ZUG6lyGj9n9V8pm1/5Dvq/ydWQivKHrAF8XBhncHTOvauAP3Prl1V3
kkiduihzQKKpc+pbFi17fYez9iC2JAU8DXxiYgsfUhfxGMuiRzw2Bjrgb0KC
xqyaSlHPSP4J01Ocu8TNaFRK6mnuz6kiJSAOqsc2KRqtyaJKPVcQYjDD9taf
7v20pDvwQ+8lMaUc+txmkWdnXlMgV34Tin5XQ5UCU/DJhr3eT33WTUrQxsh/
BIRW55JxFJCpCRPdJ2zwXPrbiyAm6omowzAiCVwETO28ObRlgag7CQBPJcgV
xaHrZ8HELMOdytjx6Q6b0tzawAjIZqQL1S/ItNULOOJTuWX/Pm9H+EY2BIZA
rg4KOaRfMtyDRywZ8b1gecgMiR9nzS+SyXQstdUstwOr8rdISQCSTIMd5T1f
NByy6rtJIByAgY6EcZBJ7WufVIgXUJZlfImbSdQy1OctY5v3ZyMZ6/14DGPE
j7fPL5M1N0eT2jM3AF2LodSe6PxVT9geg048MPbkL//lOuCK1fZL99fDmw4O
2JWvgJCzefrlZH0ew4FaKjGjkrnLOn2BLk3jmL8+bSDH+LbayuAzgr4su3HA
7TjTqmf9PilxUBPTRjTpRo/lA8Hzs94X+vcH41FxMkadS3VgTA9JkQ3IG3v3
hRm3t/aO58NeErrIrq8emyMp+e+7xCRE5imegwvBJ0P9DF+GAkIGSQxNrdm6
gVNHljGbhaDuEkfqzg05vzDB1liHaw1q3H0R/bCvexvBXG+uDY5gpY+t7fsG
tFDmWo5qG/La+wMkb367IzAW6kggBVtXNIuv/+pBy3AWPxlcN+KyYjqKNNEK
uEvXVuaMZO2fDuC3PiV+snif19YC4GUgbV19BFRWiAYkKsWUma8M9Q0zbAd3
4/M9BXDCd4h3KZvIR4T+1PqSnXgs6FG7qql0r/+p65mIMP6jsXUgSlZcXMBV
Nk3O9UwKRuKxUqhFaAQTnWxj9DpndCQu5LCPVjeKEUobg7zoEEfVG6LnQ1lT
g2mdSGYkfts368dF3zfetIqELkrjroNfk2xY3T6FI4Msa+vZ9+bvbQKViT6G
kdAorMF1roPsBQQ2MW3LyJ+HLF2EC8g7bGOUOKwuUYVe8jiesPxx7YUp/w68
vvGhPjTPn+5g/HqLdrKfC31oSYUd64FLfGfY9J9RJWoEmrEu7SNvB+doU+Pb
8wsbBqrAeU5XIj3C1OO5XumddcNJd8Xj5gREDY9Zn1kFEsx0372NSKWczYml
V5/cqBXR2YFFVCy03D0GNvl5yMtIIMFw8EQXbjKigKeb1Qrz+j8CxdSNGusC
/rajiP4tNp0H3+yQahSU9nB1iHPZgN/K8FJt57fwV9n2/ysXcmPRfsnaYSd+
S1eu4MfgWXR0HhG+FW+s0lSWxmXRIJ7VbtYp5+pxC3nDMsVBETKhokj3kS7e
L7QUCZbA/pZYFc8a+HI8UQW5ot9/l43zwlnmtHJG0EraArLtB//+W5RuSV5V
4i+dc/7DM2g9fVN5JdvWGnQxMO6F+7j7GdZxqVrNjKlwdmIJFj0MaZ0FrFlY
hYWWeFwcizmlt8Cs5Or3VCwK7jplg1LvcWcAus6hF96pWQM80AYlT9MaHmhf
7YzmcgM3cWfIRiHzqM2rL0DPYNb7sUan3adj+49SSmBHTNeJ+w7hCnUZAmKD
bD/DRRfzmtHT/IKcbUd3uw3XjB4aP9vDZiRBOptVsxs1V0yqnWMA94MoVS0X
O9Yu91O/RWoN2Cy6Cuc2cfmmr4pLWGUNlsUVRSEIVS2f2yiEzhEYFXvcHJWg
VZreYNin3ywZ6ukziXzX736HSUegygmffEgeTOX22S0VeauSsyDVyKCLLTK4
22FM962x7mnEOvTK9jaj36ONAofIqO9tnKOsKz70/nazRCtUNoBhFKq+pBLZ
439Geg+sI0xsIq1qKHrbt4ohpBsM9hEO9DThnrodrEDcmrUMbSZ0E1P8ZKBY
Ql5471z6zowV/U/fNAsR3ZCkIbbcfPGQDAydB25HjCMzM8n6WwBPBLu9JhDN
VTLzpGcn64yjqs29NjXcdVv6g5rjKTjAefGpu+p5pHYRj+D75C78DnHcuDtp
GxZxMzktSEgCq05R72neeNFaISlXt3pWjkFBn4b6W6yeJESSCUkEtkscFMUB
qNI8tUNvr/nNZcaikOC5iTS04a20bC9Wni+gyWQActqyTZIynq3pvJLjtnGb
YQ8n+qhDLaT/qXoiEZ/sM1dDbNyzPPMSYloVwMIOaCVJ3+TQRcHbqPzGuMAN
q19ZkoXd0ZbZ/2IZdOw3Rnr4ZSEb6rWx/aZjmhYpLTqcFEoYZnn9eSkz8FGl
1lZqJWDntwtA8Lbm6uxCxt7k57uwVimKmdsG3A2R4T9o/YZqp5nv/SMs4fqs
OYkmxBX0FBqgqLNr3uKuhvFiES/BudhZ7YY2CXv6MythT3jEwnV7z4Ftin93
COk/nacOoBOItV19tA0jx9ne03lf2WsR/DooAg86LNdeiXa3V0toBfAnB+/z
F7O8MiaS43Jl+Pd6vz4oQOF5j2yD60gR9iaXu+GyImG1Nm7+yXpaBerfnRfO
gB7nKHCHq4KS0VisygTtJ4w8e9EAS5H7Elozja/64KFNtyhkESymJ8NpBzKN
6C3r2tCWJK08/REXMLEKaNvxB039DINAKCOB+AM+thIoKAtS5wzt/XsbDUw6
sjsetLH6K+rRnu+A4p5+ymJs6eGV9CYBfIfkCIK4JgF4TIBeKQUQsba+unkh
efvXuM+9MMXBjoIwIbPoN5gaXCfYP5FuO4yvbBbu9TshBPl3LNj1PW9NEJ8D
mhpElmLXmusYSaJjCMPW6LCUv5yfZtO4hwvdkYjbgiGmRXNcGx3a5P8/LGl5
07BP7QUtJtQSK2EwqK9Qe4MDVOkSp/6sbina8X1nV5iAKtNm0dNMqrZvTFvK
cMZMX5Pojq4rK1yq/yo3OYDXDWZ4ukGKJsg0045UyRTdk9mzeKPivIPbp+M5
umtV8PgIOoLxaW40pa/95kZpM+Zhmt3yGqIeHyjbRJXyRRY70Z0ObRSLK3w5
Pgb3OqeFs2xlw/c1iUZurtG10ZeS4yDp9SjvTERbqEi0t4lkQGpU5w0t3HVZ
b8Kp36nUicDM9iE38k15guOLBRphLgyZzB5A8bNlhZbBumV4P2kt93hkqRoT
7l47L0GKvi3uhuz7quhpahu34NPOf0BrmznAkGmjTADqMcrLRBKAxaFv/Xxc
kVKdrlZifJKR/n5tJo/nIs4Dm/iCCl+rNscjEp6rtjjdpp6ia/gOE2gNhbWt
7msfoUz+WQGunUxqDoy5y8khYDaXml/bif9HZk8eSYnXsck9taC4+qgD3Iuy
+LkuRT/z50PjI6C1K7FK3xfJoqEODloJeSyMZmem2YKJ0qXhCAK7JykU8UV4
rtR3g51wVfyYsqrnynmmTsqctydwNzEzB8lpuZNxbr1sDwj0l6TyPA1c66vs
yLIhMOUpkvYZBG2/8FVRMCCnIG/Wx3rdEEH5Co6wTQh53jwVTtHfqopT5NXA
O57TfnOwwqS9qatQofRIyO5tL3yESz+lvZ5i3WQcRHFqpvXSdCflUejS1RVu
0INBwgiEp/0H1wSnuDc6B5iG4tx3wn42hgXp7fzgkqcXdvMAEZdcR2VoQ2fp
DSjmVm+WLTPvbsziq0IbtfMNcobLJTBg2CnqGd2UxOSVT868OeguUhQ9//2Q
Po3WoheFZ46Yf7DimFL+qkpGiqyEvGd+yPjPpmlL3XxBwkrucIhQQd1ppIFK
MxQB9Uj8fqtHmFA5B5XOI/XLCrpPGTcO+UFEX5Ns7BU/KxRW7BSaEofipeyG
feboeK327rr2qQeFv0PElEgPPzNr0TEY3PD8BbqkdLjvBQeQa+ClatBxOaXV
UwVMCc/SAWxiW+BHNgkKfS5MCymX/f9H7zP4npAy9DLo07fxtIddqEZIadbW
sn41rxKMzDLa15WayNdmW6y5ZI94jYoZVt/m+bhuBRyJGw0ezLNTOHEBV+AK
8WjHNUAP4W/gKFwcpTjcFCrKvbE1ZFY4nNxVZBdE9S8ULv18coO//KCPp8EV
okVZaoLvev46OUgoo1T394818Kw/uG97n8Gm9g8KFDaNBm9kjeiGdnsAd7cP
leY+nZiS287BzhQSNHqaS4Ndja0fMvRqfJ31pZMblJSKgrxhOIesht8Yhygi
efAV5Zwm58Q4rQQiPR/F5U9DZ0upVnHrmvtsfpRVJ1wv0q6PhW2RjtboJQ4Y
UB35evhLvFhPRi9DGrw3xYj0GyzT71C8huCVCfBURIYNYfyAsTrLOnNVUu+T
Y+98y6RwU0omcPx242vbOuWy1D9F4yPACTV0T3eolmKv5KRmhGDTG//IOlup
fyNCJ6Vep2U5jXSvCoUZP6alt2VWqY0fy9BjT3rAeUV/0bEuEERHoVyfthYW
KDhAysGdICm1rLV8piX5i+zT9AJ+NMcRJFNhiKn+QpAwdVE0ziZOzYnZANHx
t0LMrEq9bvyeHNdU2V67scBab9hSUi/wPH446n6Eex03zr7A2RwSmbS4T90A
jlfP8Jg5TTrlSh93B6nkvOrYunF0bPYUn/1MBq4NVOkgahGdXPNuOlAnzhTD
/a+UVfF0q92fZWjF73yoduzQkJPD2udggt9VGal58DEH5BkJP5tkztJR1dEt
zosLLiLc/2YiiUuYGKwkiZmbng3iQpJJgWbuU4z2Kh/GF1K3tQ0r9R1L0ER9
KbBWbID9/lVKjAPnKh3I3/ZglUQ5FJ88W6VIwQaEstfwrWCVZe/yhjWkPyeR
3K5VznzhTZk64/8XJech+WoLLf3zjzbAtVmUHG1fuu7+FeZIW575slcQZOPy
NlfXWZH9857wFeIOFhmtwTo/Nc8rWVOH5dJqmTy/f2yhBfLgq1rLtmruFLFS
LZXi16fmaeb8WxdV6S3phDa8s0eMv7biWd7wT29+xjFFTZKiuBel0ggVJAIH
QPIcaTajL2dIdYxwnMb/seMIJfyM0aUq31y5jJm4sehiao8XJoK1JVnKMWfz
ypER/fREYCrtCrSvSegHmMsWZ0Mt1/GBPNu05wJhuEmxcmYs4q5qgG9yKqhk
Ypi7hKk25iVz+pKqyYZg1osYIuVf8kG6OayWUAu3xaMS4z1tNUOZDCuslTKK
AjKOje0x2EFUmAc1oOUaBTfjoA/g1o7WUsjLe5hNPUacPZe0JqswUJ640SOz
LqWGY1SZ6j4+V0vrWnfdl0w5k7Z71et4TB9U2H7P5K1dQHZKDvzENX9YHLLe
bsXKZ33k6ATXuAOg1J4fDxxaOLEYmlIAkMbj6XsYcoToBdZyKzOrCDhlmLfp
PGqtB8hpI2iHUZyG5j/txgC7j6aA+ZYJ11X5LSaScABhEBY1Zc6Tbvzk17Cv
Hky7y3WwISVgIS8uWACToAL8jk5Qcu0pTyF6A2t712Ass/oGEaZDZllWisvc
IxsmZ9Lfg1eERm+rYbqOrStX7qoD9XP6xxWx6mA6XJ0+Not2LVHSgGA3Qvys
hwNV35lnyLIkfAhClzjO5Wzt3XH5prtlMY3uQ+5ZKDCEpQI6tEMUv9KzoYxc
AtzaCPlYIWGRst0nxuCQZ1uBU6D6t+DmWcK7Y+l7lkWmzBt9nN+LA7CHBwCI
pnMaLsNw3Br/XLt33PoEV0lMTB+46FMgz1Eznq0SFKWw3171bW+5FQ0UwnSo
qlIszH+I2KC+XfPmBwAaMzpTF/6xO6CUrVN59gPxhodnvcp5r6ndC/cwnPvA
617RqlSj3Aj1P4bmsK/Y6nyHO9vDDlm4FxCC3KFCUkrNw+l7q15wm57G5Sqz
Dqcjyny3AevM1pNuICoeuNx1dm9F9gVrpQOE5metCRWjV7The7cQAPZbi5Rn
tnWx/tCb9BbLHFN1Vo7WDq2okh+VWAlD8kMRWsjuJF8JBSv4enLQR4kC7BWP
JjtPFEhbYKzRUJibxSjDcfkdnoKRleDkPKqsKAdWgMjIAfjM51La/kDQ1TIZ
0kbk1vT3euRdIztKJF1p3CNF5lj6i0UzQjuZDECEtlUVGPK3xnTQSyz+lNHC
w+bM3eDWGTMUGIThKzS4T56TfB2/u3FWlkMENz4QUeTJPkxTwBaq1YmI0rgp
cMYF0uH5lVcWbJRPIDoPc9WM88m5xd6qS3C+izFr1AQGeYQK84S4APRzHvs3
F3kx5Z8ZSEFGscopBa/p7u6vp7WyB6Y9LOiQ617GYN5VPN+Cvpwu6dG7cP07
z3rnoPgQXwyu1YV/a4zkSKdWMjoJI6Q5LiIG3h3TU30jxyRlE7ek3cmwnh8r
c+3aHcc9BGIKBT5FTwH9yerNHfpOAs6J+0Qze630qGhAoehkpwDzES93ok6x
5oYcxn6hM3zUtkiBnGcCfH3Hvd/sevlzyRPwqwwGfBZ4QgC/WkA70d+bJXi2
YTzSIsldTdMTfAN42vSXdcTS/+dZjwldqoo9Qup8/xhmDx/n6poA642/ESGm
GiZvBNVyjpQDPGOuHwWZEUJoxLMQhQELrV4VYVTYU6nuBo+chN/RoQRhXEu5
JmoJxPTsYQEMOWMGAw4bdMnxuM0KgDqoPQNgjqXfIWRpZ8jfIWo4+mKXEoDw
2vIxiALiPOXpB2z8S/lrTpREFLLRCP3LuIME1q1KCAUdM51duF323iu6O8br
GCrAQMnNZ8LSUj4IwbCuQD/NSH4UbdwY9RX3z4RfoyY6pBitViH+0ORcMX4a
as+qRa4UXE/sCZoA5Li9lmtYDeBaYZn6bOTeHAoXEeEg31RKjECT8zpFRGjQ
dO1GhgNC0bI6yCVJqsKYmV4ki5pswtHNf6zA77cQ/8gtVC1HXuBCzShB6PgZ
cWr4A8lhf3kbsEQiPSUQeESd9TasvuPce/fvJjoIvtYF0KMgUkuYYIzN9MZQ
H7MMakK5wmE5qDfvPQUseRCuVbhQ0cUOwH1nodAtpbo2b9RK1rG+NnIZtZvp
rqnEHuM+Ae/IIbA78LmqLYpVcdnLDGxYO3rTz62Lvm8hg5TmtyQRPZo29fRJ
NDvv4lu82y87Imq5iNqiD/VgJYP2h8lTg5WXsB6hrLRlfJn3iTKgGwbHuRz3
xuvVEHuXd/uVaSjL18rPM8ytUo5x+rMFynpcxrYj7XdTLSkC00br70yKBFM2
ljdUz3esAjL1QvdhDxHC448/vsvKPN7B/yyMKRFq8uV7QNRM3RBY+WXNwAqY
XWdzd/7n2o3PjkwTr/zzofCmnVeUyJ7O4g6I2INxypRSBrAHf3bhn73zCmrE
hioTqn4rQEH5qDZK6tVXEB8jAZ8DmCSSQSxeYk3X0HVe6XI0h81butcKXIvs
SmWtUgSejojV7upXkTmS5M6tzFe7fhquKOCwP0W5VmUzjySoeMN1xZYjS2Vp
9s1Zf9NhES1CouMUa9qnurXY1uwqiEsfJ6ecSGlEKPjzBmTer5y2H4eddlNO
ffMFHtPSOPLmcuXEICGIp5nmO33vnPEzFx9EevMv7A2FykeymWkQcz0Um+eZ
hj0MEllZAWZr6OYEf1+XRUMutRaxKxIn3UKIebT0LmheiJhkxx5yj3/aZA+y
/yR9tEU780SUf2SyXgbdtslYmFINlEgbAcBe6KjPUIoNrCk1SNgdXfCvg1jo
H139CQyNU8UNv2/piXN5AGIQ686/gkjIn/ZYB5tGp/311AOKwxUPy+RXXP49
/EwSOXmNR/AE8NHOq1ogjzbgNknvB/n/wy5mZuBJOGOOCu14biZDMKoN+jmY
ST3qMIKY7WG4yo6j689onHRfL4MhdHcOLVAO50R1XHM0/x5fhwQioQwiqjTN
J08THInvT/nFXpaJQaNjqmJnNO1ZrnFZVa3qqBJWVPhvn5i9T7/gp7pbmzQY
/iJWVuzxzYklUVLKZCidItzsI72c+rQhbr9Q7W41FnB2gjMFEUOU/QjSWJHJ
DdaoXs2UzIbRdieS84qELbdyYquPZxpXKIwDwZAeaVSIFCKXSAxFGoqbGMr7
XEcFngekKhsgsyh9IhCFfd5TlsiKmeYg1GUhonRKOQJweROlXI/2PTqFbChS
SvaTWQmnS0pRzK6VmgWTAfk8PBO5YK0iWJoz3sLNFKCihTGnHpEqDhVrxHsN
rJ2VUEr5Le0gYN3n5kgHQIRm+uhyLmAuSUNv9LZmaKTR4eujji5VAkT1gWxl
1Wlma3lFpfNQo3F81halOPzIWXj82VEeiRcNbwwe4jiLe6xBAduhtdnOM9vT
nJKsu2xcVK5+wuYupVU/QbBEurJiWjMG12Vrfqz3ZyO9KsVRjIj8J+s/12+g
7fYoxrwpQpOj3/zup/g+3EpCvvbsMpywue6AFfbqgJB5/FMxkGfqttYQR1xm
BBLyO7aMhzOytYmeeGg6v5pac+cNSTjcwsMmpZatfGl3W6AnWp2dlciz3SDw
MHAkKPqmNtTETsSnJxhaiJDj7pkkevVnwJVIa6U/ufL9/VrLB9nwwjesL3Rg
s1sZ4qlf2fDNguXt/Sboi/BUcFHLKN05heFxayoV9DAQAwTK/K/K3UMH4p3m
cce7A85R1VOsMq9v/Gkx0RKxvHBgkxzXNgkxV7fBgt2GI9kbeYwLxcYn2aOb
kCTpwnuLxC/tf8KOWLIcoM3GJ4xmUIZmQIwRfgnmWRE9zmyjkK6/5J5wg9rC
e7k23XHBZRSV07HcNk/ep1lOxTYScnYV2Y0GC+HYw78/2dj/Tj/XQ0AVm7mt
DKvI70z1BoE1asU2KiPOtq4Afl4rpbfkyoBVXs3lIq/3JNd4ULH0gmA94q7T
OhPVXwLk1SOcmGJKrs1LsFIWj4dNLHpGlT4I6J1AYB9rbR0Oh8b5h9C6bzKc
QHpb89BXzG/s4PXvGeXsi9f/r4wFuUZ1MjS6LONWQoDs8BMHPfFUD+xiZoAz
zU03hQ508s5TqOPiIDEZyGqPADeYoQP/qUkw8A8TQhsNmi3EuI2TsJbRS51R
tpSGa5UnBSjS7y8EzLC4r5n2F47ezE2txvj97QSNP4rMq6bdz0XixxaRROne
hngg9l27fMHarafIf7pbwikgCcVSVG1qhqai8JgEcK7nUZGXkAmoHVR2TJlJ
Rn+JUSOWcg64GmP9mg7ZSVaOVC4SOetlS/UbawCn2xfmDU7K99DmsvdULF4M
pFoMwipRqreIBkvcmW7ETNTf3/8PIqj1XOfx8lntqYTsatMv+opIRdPptS2d
FkK68sTHRz2gk2sTT1e6R1zGq5oCI9zOL4G8ymVkdJ+cmq+RhwGUlNCo+o0v
XGMb7hUHrRNHpga+kPzq1T30bSrfwcG6o9R9ctyWRcL8pnGjZgyoTbGfGPry
bepYuZYUcdWGceXIZK33ik4M0s2sKpLzhyARD5LVZc3vg+OXSCEpwT8K8alY
UTDdSdlMki+qWy0BVcnItfPDoLZvqXgkOjx9s4j4t490lk+/AV6oy1sbILVY
f7dSD56hLiUoUgDSmttcvs1iGu4VRpPrumfvxFyks5zpk0Q8hcj4NOpncIfZ
l89tjnAM4FiCyOtgsFBpD4VmF6rKCwpuT5aFrAcuZ9XAEcBpkCoOm8YQZgY5
D/DShyMtNIxaFJv5+5Qo8XIKr/NVV2jzoHfgT+0SjdU/kqZMxTqr/Noysdtu
2nSj6teN04UcfIjE6AdJ8siE8lnAgYhOmNEdICxVTomnoYfzrhrja7xq4I9Q
0t1Ou4Gg2lvUaej9OG8E66mKTCuVmW87y8XmmpwTw0W7hLfijv83DmYwwSqt
o1w4UNoqmrTcgBMsLTurNQIjibUor+Qzrr+PKc5BThu/7BpIU9VXk16j9zFP
GWcYvj5yhg27ZsVs03hRO3/QnMdCH2CfQaEVaNcZyS2tOz09fO9w4bKgEych
0Kd5ZGN2g8qka14euYe5Goj4oTv+EYGSUyNrsjMPFgti0TCuscYxp9MrhUx/
U9liUw2a+/n0PkfmVcvuoqOIE5cTZKBpavHc7PefXwsPKUg06+PNfuKrAIVu
RbGqH1bxwFQ08wN0QcPX/rBuDMesKubHDuOyHnMn8qArm1tGjGdt9QvTvPAn
gEIhslag49qOuuol0hWlEwg47qHkUrcWspBPturyMWxlBQw+pvjt+q41Op+S
j4lsymAINljwmzghuiPBfKfnTK5Ihe7lvfM09wZN9Reeirw2HIN+g/nAN+Cd
7AzQGvwgeLiseESIGq6JyXPsw0izVB5mTVRy67IF9yR5siXjgdM2/piYpqrW
FrSH0e6+og1yy3gcAuxtWj+xDXsxmRQFopGQT12m1psulZu0xtw6Q+7v5USh
FeMmov9djOxiERKyiE1MprK3xL0pXbsZH/xNRlPA7qGzGpVZfSctoFHDSUl3
/li5PtLU+yEz+HClSOKagGTYBtRSxT/ZVV9en+OAKzXgaG14FdZl8oQvW7Ca
13gmCIv1Axl2AVRwkK0rtsGNK8IULIv7glTj3lhP2FKZnyJuzq/rhZCHXTml
fWmb4gJhG8asAWSgtlMk8jzi68uopzBkBPmC63dnq3NNku7DrBf4Bxg7nVqz
XHBeunqrbZlYSEJw/sDyXDcWFtSV+7c1iaJ36mjr0CPQ3f69XBAgTlyslEJs
b/57rNuOf4k8SUMWADLLdlu3NSyGmkgJ4zAZkmhPvp6b1WFV8zzV+rMbqEsy
Um5zsFqpXJ3amHlkwL51tI8Lirq1ahv9UMbqmVlPJxhjjnIs0FJu4DfL++R0
NnLqIwRiXP/XJ0IOW03PegAwRg4l6AlGY9HpnlmxXFZKBFi3GRRUnjYY73R4
G/n2ARxpK6q0/XxYWB4ZORMwSpeDfM/x5BJsp+3pmQe7bSdeEvatQ1QWL2Ci
ChvHjFIUEHwYy/f8p/8pLeNMtY7SS2BBc5KfiS6SpHmg6rkkSBKRZq7myYFM
PyG1MTJy+kDR2cI/3zOKkN3K2HCzU0Vp5WA7aIMn+nMzuPJqmr5KRpVowbxn
YPUFrmwRGEaZuVwBnKpOAxIPh7USythz/4QYlT2bD4Q+56j39akXJWXwEKhK
b9Bi+C2QLVSWNtarcMkxRqEIE6I8LkF4ef4gh4gaoyRmrjg3F5H6LpF43jm9
5AKpdn35Ugm4BxTnZaf59RbgUoq1MpvyLDyj7hsE0B4zHaI/iDRGaq3ycTCe
eoKFseAIr0a69x/GppAqpVizSoIOi2574djGg/8dPc9wc+60d3pvWk+HtdqR
JmeVDAMAx7pcgac3/X5onjD84x2F7AZPtH6T/judcrFSg1N5Iuj7ZJrtmBOK
BLn5YiHleVvZz1GP0qbIBRMQkNQZsEghKKQwQG9wBcUfFNSnULXTv6xLOD6z
WFXOuKrzydnmTqK4mSwclBdtelaxC3UE3JshFdJxmg92mNIP1PwJPZRsv6iP
nznO5rnCizqX1ybSHynvE7rXUyCkvYw/+HzdZ6ECGfDgCtQFDRU7TOPlxSsH
7ku179PczMAs88wkdLEOEoTWFJnmpsyqqgQYmc78qsufiheNtH69GqIh98xg
knkizr24kIwsaL3fmm4ZYI5XdbKsg53Sbyb2jQrhXcyX3XOBFc9uvy9z+jhM
3tS7dMznhrssbTmBWWjHwrO8lTu29iV4BCDoQsF+UhbbeizERyDchrz54fxw
L3aDoDNcHk1aTmVCVyGDJ1iO29GBoxjfQapIEdUfKu15MZXAQ4ha9Mu1mDpO
qIv9v2ZncurkKORzZu8SSyb+VbTBJcm0YwEHyLb3cgxNN5IftLSPu2G5vy7S
zjg4Oo6ogRmCaHF+m0CPgq5BtZ9Oqmo8LjGQ24gTNShMc0/nvItS4ZwYJOKo
DZ25SAn1HTToLi5ccvqLqkO+h+6gZCiFYsFu/aIof6VwJhGq+0ymP4HfTyv8
FunZ6N7KUhELQvqbqEaDRTvTzQmOKhcB1yloAVN3gE7yX/Iju4VO0Ua6Iwab
Yu9pAivKGWVHTUYbHBjwgv7h7hkaOB6KPSQm4ErY6dO2UdGQ+uI4KAe8nFw/
im5tm4VqUgCTK4xxuawtqWShrp/sMMzc6sM9Utjx0pVRN6A52aQN3/kw+1AX
/trnrcCygPaI6r1Z8dDIMlsd0z8xclTYAFo/DL0ZCHglRxBkoYXH5NW/KIXp
ROfvh4J99772H/HcGOHEiuCRYIkFfoNQx5IwzIjLPpvIr0t+eolx8AGrYdFQ
vIOFC0zcL4RmQG6zPv9u4emplHrbJShYsN4yRFbgpsZtCrGJ1GKjgYkJ3IfK
urcP+X1RBzinqpbWX9wXUtyx19wMaXGOyKn2JSWhf0GnfmuQHA/ww45Nq0a/
VKb5gS2JYvwNfQGwexly/q/3nMGflL3mBn7UaKSgE+umIuRaLiOvy3JVMDU7
vG3nYVybZ25i2vzo1qveEPbnPtN+EBZNIbyFTd/SmEmSjr0A3CV5zyyQfyMh
fCFPbfsyJoU41iVOZY418uaYIELcm2OYKPumPeMt0CaMvc6jA86gENJtdB3l
7o9N5mstOpLLf/E+MIVv4wdG3VnsHVCvp75iK0maP8nb5L4E9IHJ0dnMdxi/
g8Fxq5TSL/8kXsxtfwz6lE9VVbiifrjhGMRv2bF2jKcwqeXa+u6xY38nZrzg
4v9vjh/J2kb2zI0cQagjHF+4PzoG9g2rx/DkZbRSit4EeY1aY7DBBbbf+m/M
EU2WT9a4MOrCevey9ZCHR6M0QIH8/YS2sTdNmGKIN6EmFAg5mAj4sIWUL94b
VAeSIDeoS0ZkqKlzktgI2JyZiOHcEdWqEgpXIp8KrE93rztkeLWwp1aTZeFU
RwODcoQ/EuAwlxWE4CHZvLwkQJD2gvvhx8c1LX/joZjnRCIC2Ul4UkLBxEDt
liG2SYweVo7Iax3AvSn/t1/s+aAA+A3hMRtmWJ3/OHvnFcqBhj4oDaUXcxb4
2z/uTyrumuDTdjQ04ClEaB/ChQ5f7tswqlPcG/fpAulgbkwAs7bGfKdM+36S
KTUapl2TP72ybaELU1rH/DXdsfgn0GQvonYJU1vtKMgSKcqVSGNoMfk+PhEL
pSG4ZqzsiMsZzBY/QRMnppoI9IYS0oX/6907h0HdUHFeimpwfjwcY91ks1k4
nDSxlYxAtjQ+4N0TtlInrDPI/kFYj84C771+4zCBGWMY6t3nlgGdtKFRi+Xd
MfYlMCKbRpbXJQAAIB9NB8Yc1JY4T6AStH1vAxDayTXGiWyMU5ULNuodyGKB
1WQ1lKz8rNKkL/yp1iHKYFtQQhwtbbWb4g55ByZnfuB863QQAuZTx0zUwkK8
C+l3q3yX9V3+DnFiUVTb+x6+lN/1tn44DKP1DMOtTtEoKTd+ouLLw+jIsyD8
7DV0o8ksiwajdUCi2vMPgKWv6XcUBuQJzAH0YVf+WhP535UxLeJzavx91Z6H
Opi7l6dXUc9agISNGhmu1P3ZXdUeZgvFAoNCUi1C9CgOEsQEA8m9sVkF6hEF
StKNVoOLgPbWDJegNlCSFsnk0zoRuurd5/VwWx3VTWBGKSQEXbN9oSYckVzb
8Ow3JSZJD9vHDPBYjuxJTXvtsML8DZxQIAYMkI325QOqMk8RMQO7o8E2mj3A
1cRQBa4/HyawZADSBYYfBB15cb7UEt8l+fC5chsWgwBZPLfcncj7OqdKZcTI
Fg/i6BWV3PqXMAxq3KzaJWgS6JFl9tWI2r9/G9n/zY3IY5dA2y33uH8hms+l
yaUH8W5lU322uwBo96hBvhGn9orRbcfCBCuBhaq5U2ZTJTTOQUgwrA0Cu/zI
XW/6bAH/hwmmz/eT8AKlX0C0/Gkulpk2cwgikOZksAFSFmsyz3LI9szALz3t
FLKUoPKg0WCPdUubYuzwf7XdZGS5TB5HMFtW7fuferVGeFuhRtW6raAMWgew
4DNhdpB/yrGNeCWQ29RTvlOzDLMvFi7H8Dm0XmZ1bAK9byb4jA6cmLVfG7W+
hoT63ZgXjT6LYxrcp1ykAgsRXDLtesotV/Tg7eoHczu3jTXGhHANibXP9qZ1
ZX3Hx3ItV8Uzhh6JUywjWaadZtfSOkXlW5hGK3wBvNnxrNTScyiL7CnnVZg+
2nFYOlXvinfKgVvgYAIup2sxAu+Eg5XYLAiGYuOJ4byDndCENp+f1ZfHMRdW
cp+ZmfDo8JtTAnR7Wwrnn8bDiVYFQ0tqeBtP0skcAOl/ik86sXe9dpaSYphc
CMifQ2riQZYsgrlRwlZx6CK5MK1OuZNpHIB5A/GfP6cJwRuD64lVggt+ebdl
SLBBcd1mscX+wjiYSUZCeQV7jh8+wT+57tdia7E4EH7Rkrf2a+GJEpRafRvp
RQc0d+gSi7XrB57k2DjAyc+e9rwbo6QmdgrEJuHoWJLA179wyAQYD/26FsOF
lkLCkELgnUeKX9rcdA89huOsAHmnM9ygPOxUaXz0zXbC8BR+MtITQOmbBYla
BdzWDifTwXp3kyM5FN/N6pzwB7Y9RmLS8SJAEC2cZ15LCyMPAackp4cBCnj5
HGeYAxKzJ+Iy3gpc4Qq3DVY7yK3PoVzMu1NLllsNk2ec8g+nzObnfk7CMBM/
hRIwvIyMiNnHlmTRSO83VM+DES3+1g/TATg7woQz6hQGQCzuKSX7Ynun+OR0
2wdgPiERtyt7Y6CXnAJJiLwEHYDBcrcV7vJByaDM1+SR7T8FclFnfLDxWkQq
fzjcck2/1LqIr1hd27T9P9LDZU/Cp1MsHDLE9P5VffVYwNRfqUAgw/BGnAdV
N0s4BMEweNpsY2M6NM0HqIXLBE7rEkfEjZPCVetFEIJO5f5Chq2O+AQBvFE3
FMGaEAwVm9NGexa2iP6N1liku7MPkaqBLcfeOIWxZzOOGz4JT0ofXhXO08TO
7cwJr3OF96CrIZwaMgQt/Rep4bGg12TSYEcJzkYIoYpNdr10jHRy1s3Kv7Zn
ehq9WFolHczesCDzR4tt21G8X2b92OW8kX7/MfnVdMQHvaW6GabKoA1FdFvy
Bjbt2xTTFW0HqJEDPQZQ+Hl8L0qfrkoG5+I3cihSOc/T502USGznKAWgMph9
m4a88zXwHPlaE7VBzZ6TNcF6F3vVSfE4KDSG2Y05WqydkzJ8WOQL9jY0lV06
jPThNW/mdi+NwwkEHVFft6LESQV6a/mNSWopgmG10yjwH5d52oQah3D6FeS/
rxJwYBYHKLSLY0Ejy0a9DW5vVYPMkDO3uNOHgKCq7QI/ttrCUZJqVXseVws/
a1kZAPFhD4krhDJdF9YjdvmvJ2aWTKvMgpSa6VSV0nvh1hH6BiLvvVz317zT
nAgaEDPSvhUMqJLL8aA9GrmGNjaVZZI9l/6qBKQU5id0bA3/4woZ/gZXTWiA
cL0U4mesHw9RmSWS2UrPt+q1QJJnPxZ5m/3axz0wPwKnofY8qmE8eiet5LH9
IXgEN8nDcJ9arhUbNnazBtXfPY+jqQ1fCsDooOK9n9UKz61iMALfEt+RxCSc
yf1+1fCqDzYHWx+XcpjF2KTX6q37YCbhI1wW4X50wjocnxMs6AZDOeDNvUhi
6MI17Bbdou1OT8tyH1jkHvAWce1hucCf/BRDhqm4iuHTq4+ZawV/MVeDdHCw
TVvUgPQlEh5cYYnv7bo1iPx3mHZZWGbCI8BhzcfE2vOBfjsHmQlr7nOuRIbi
vyktXu+D5+B/JRXduPq0RrCOe8fNa7Q4WkFChXsXdfyHvbzHiLarWIB7EIsf
9OMq76ajz4qZFNVwAY5ldIOi4cUKm5wW4857jpQxnr9Je7nROoWYw/FbquzQ
/u5kkr2N+e36O47zGJw6lGVEef1DhSM2ikEhlJpX0nI3hO1+OghQ5jbUsssb
7JSZVVLja5ISJ5Fls5ZsUqOIdOI9kUWzDGlzs/spQMy3efzC95+JgX4I4LH+
tgRpdJd89J5p05Ic2YkFHWMLEm2swh5vM4WitAh4BOzHb6rw7yDWz2iMTiDQ
1P8iUn7hxu5y8ab4vbE8RLTxqxNGUMRUETo/czenf1Z3m0h2+gLO1OlkiyJK
NJqHuFCXRt3GGz8agoTXhswfPJP3cYsVyJ9prLjthLq42952OwsNDIrp9hY2
cM4xBlF++NLt6cOuhlJipdL+QctiEsbamJINyCHMf70YmYx8uHzkadQfOv1Y
TSjwnYsSAsbkRn0K+zGNOU8xWknr0FFsoDCB5CAlMtmPv448KFDS/BvVXeLL
y6zYYpjOgr3ftZo/VezQqKZiDpV4gl73o33lR+I8K8O/oSS/mYWy+DxAGnGJ
BWrzknIsdTsaBpdKX2zN/F1j/5Dw7IGK4AnbF7/iR4mjJQmMe2oNaHTw934X
x3aktp4ODwxlJ2nl++YZt6Qg6pZyqp2QswS6za2p6owZASSU7mmFM8AQuLnv
77rYwHOxmSUFtgllXBk9A2luw/PCeca5qmzzkovTmSd4+fsvtXdEZ32FgtVy
u9HXhkOeOezKMdP7tu3ybXjrQFmyDfpdX0361jKvBENiYlBBjXwQREBIGmP+
zotl+fkWE6cbL4CfUnAKQweuI5voB+hntM+2MQV8+HxjiDF+U6wocYih55Gj
AxJ5rTMw9RJ6JaDfqwm7aZ3vxX0MWvytbStZeAiMknhMJFfJDuPJeId+cmKK
v2wHjj39SQA68puM5xVuXOI8amYMYT/ajFlvSI4/DeYOwK6ekruiYxTzZuOO
Vdtxh8YxTQH0gGcsjS9dSN/6Iun0oKyY15Y4gitlc/pmZ8IaUlbXJmECzA2w
7QWXs1MFg6KS6YtLs6NtC6p6kcBjZlGr43G+kIFeznAidUJTQTZfYWOGFvVq
Tw1k2fFUcoNJpyv2tbJyu9443f7dO3aFzb9b4KEHltqgIS7mCTC05zXFCssN
jQ6Q1oTv4XkJ1Y0XTM8Fno8DkZH7NhzhPue54XeVhPa7YXNrdHAZZ13WkOk/
McAffFH+avv2Puv5Gn0Xwzql0makGhkpnllIGg8L1Og2IDv3WMtiFBtoof6i
x0aDRcpJRt7UwcgNo5xvcEBZRRthBhjFjgWOKQJsm0z/MxUqQzLDCylXwe+A
d1brah/yPaLwMLYkxLFtJzMSw1YC85LbYGe+khQlIJbSfko3Xm/ZsMzZvije
noTlx7CBjTnSXWEI2S+Kcr5KqWsm6kGDguXs/VvaNodnyDodXXGsMB1mXelA
FKY3mtV4dPUfFaUnrsxhpS3dlYEyePSk6fjJgsH7jXSkRCU0Jsee3YYIpABa
9lKaDZ6IGeW9A71fo1ekWbdTvBkNh40fD0+4V3lnetnpFW9Y7Le66O8fI7n7
xl8Zcn4LQnRzNYp65V4+gM6zRRbGabw9WM5a9OvtYOJpL0jyYQoKy1uXWCFq
acHnmI//9IRQkKRAP47GKwXTy411dhmmUPnyZLWzfLpbQ1yG7kpPUurD6rL2
xijtIkSRM8/Pn8ui7sEZuTIimgspRzAvxUSZhrQuxLD4D9Vg4UFu267AyKCJ
wToGOITxlM7x350wXOZA3ZOaqN+1eY4cs3yBCIiEna/JKR0WjrejkqX9b+8H
6hQXWb4Xbu8dXUsCVQsSBA5suMmhyPSN3kIv6GjUh/zVh6PRufYChgKQ3oHO
D8kugQnCQVRZSqBk36gd97ARTeHg6r1L0L6/Gyuxl+1hmzTil6FPEFDEhhT4
iGM0CVPtyvitjnA4rPpW5V0qbRzwwPg1S+bquxEP9Eys9d/CyBg35/PAo8vL
Yi611LBOoBpJRnwJv/07NeoOUKtilT+TceRIEWLwfe2aBb0xjfr74AEw9eHS
TShbrL+W9le78VTYXdk/TgycwFMxY0KFtGGrhUcweAzfIKfBuBAV61q1u6GS
mU5gWx4YRep5w+wo9n+1Y52YulfDnppZJ5HByJLCspJl9dYWLisVQoeGnBUE
MUkUqk2mq4g2NrjYitwah5uV56Mn9zTRjVVquzmnA2+0zyqXYjDO137yMKs2
j9NeZJLCweqo2OUsoxEYLoIB5+oT+bTIYJGs146ix9F62u20Har2z+49Hv+J
pCu8oQre9ta3vhz8bTw2eJW1Ze8vbNNzHIl1sYFbcRmNKzJYu3gIvnjxDiur
dD4kP8T8wd0SPiHKy96wfC39l6PLWvQN4JZz7jGVG4Sx5wzvPK4tENwK4gSq
NhbZusLWX/kjdtYBj/ORewJab8pfk9AcmRhlUzt7BJ5mXiGDVOV9XSmutsmP
ftka4G4dXHO+2f4MN0FOkdteRoF2kcnJja6IJhlP/nWbIygJ8cKAwPjKngPa
o492DzSJY57+4xt/Tca/5MwqqV7RLW/I+DiqIkHgI6qL9pBXCJLJE8CQuxDE
7Y2J0vS1C4npr8KZsL0QhUapgoRdtSIsJpf5A+Xbw1iqoW3VFRHNVAmZf/nU
O4YVH1HobUWWyL54f1qiQnBvDDQXbMv32bLLxG7UpfJhmiAzjR08H7HSUpar
w+FyTCfFHyUtVWsJr5AJMd2SGeO+TrIFmeCO0xKlmKyrdlNG36MGCuWI2p4j
JIhexvn4274JxFp7XJrqVqT4ncrzt81UpVOzGG/qLZfrnJx+NQ11rrYjLN/j
K3I9u/73AAtRluG9IEykooC37t8/wuCoq6jWLC5VfKbNP2Bu8vdUuhiuqoSQ
WD503x1f+0crusjUBIyjvaw9ofj8R9sxeskW2L3UWopvPTXCQ56JeL2DVm9/
fx3s4R7UM0fv/oSghj/G0xdPpzjgJK0JpNjG1/Jv5YGhpFlOejqybp1wVGGO
gjPKD4EV5uAj/UEr4hT3xLdlU96eEnqlN3/cbhOAiRHcdQxwRtcvieFZhh9r
LiErORL9MZV6HO+IY89Rcg4Fa4q2wIZfgmW1i6Q6XHaK/v8ukMKAg0xLPDY2
4fi/xamAxzHXQ2FtY4hyG5T3ZgV+O1sdNkm152lJR3ZnvyXhGswTeeChK00w
HKZsiFbgqHzVwQiWA91KM4Q+Q20v7oj3ymEJYnN6F+B0QefBTZPsHJXRl8eA
1q4pH8aKRid0VQ2d1uzR1bU16603uZ8sPFwvTTca5MbnnU/Qdbh3STDpTrGP
xmQvEWfhOW3n/1AGqAhIVFltinIPY+RFwg9q8hAvGMIMMrqWlr1neA3om0fb
rbEQMgwDpx4Es01LClE1f/wtQKwKv4DxG+85/iqAFgiolKbUCV/LPXxW2/qC
aK8aE0d5XI5JroIy8biSm0bs2+SoxSFABOTRgxHpgtqaM09s5tlYtbKTK1Xa
o49BU+nD0Q0HQo3ChxLy9KCUqlDjoi/sCMnC592G4/NcVFYjVsDIr1t/XKwp
duDXfARpVxhKhtU00NhnAhljEjuDJ2uF3T9uLcy+5KhxuO2axacdTgp9NW8H
gV+c7csgSb/WbSUb1MC9T6ce0MXc4Z7OTjT6UzNbTzkVf9EYmuzRHmyBiV4Y
HYSgCwzwN7wCResdW+lKTh5aK3+YbGHnL1OeDAtR6mf0nNsuYOZKDiIS/kyr
AJHuQTVYQt3rGwliupz6VHyS8NMWGUVWeVzMf5VCLM+LDdALIAIxnyD2JtMa
dTrcv1hQoDgJV9VV3XTU0xCyxYHzV4L5PRgqkBT1RnTKl5lYYmKZULmAcAxx
x0AizLIvmB24S7GL9osjqPKHSqj6bP3GIWtk3SwbS3f3uvyDSf0zQ8vtFIcW
gcSrAKkD9rcTAoWRL5mKNEyY80e3+l6okh8l0KVzO9mbRr75RoIvt3uouqgJ
tgXQpaFxoF9qsyQuxy2XT+drYUvVuoLSRP6LMf3FfAVdFiuhhDoU6zn2LKN5
hjyjIaIHnMuQu1LqOOrjKWhdVEAyIQONWDa1j62ENLWe1BJH20aDbMqk9+kL
5i87G9cndOO5Vt6kmm7CeeKdPoppzIJ6AI/ZrNz/xFN2TVPv4seay2v4g9Y1
P8sstZgKRoEz5ayEuy6EAzRwXDiRpRk/bjW5GlGtHrOImhNbtmmP3G1jDF2q
9lJ+4ylaboebw7HtxI7TNM3DGsVpaaE+ka9LQtOp5zWO5QWU0KFh8O4QM9VI
KHdTmVoAmmPNTdUuvFBSIq2vLYxfgzuH9x/VoGU3XOkN+2gifb4T+5/mjoxm
nctSn0uGESKi9m89lSZLWBWqAWMxaGn8uFYmH85ww15liZ68QMmOgNASxlZr
zGuRNaIjR4GDGIkmJxj4a87y1om2FBnkX98qFW1x820Sj3QneO5sJdf0h6XV
AogWr8uoTbMZKBY1KMHeHrC9vtyVMy4uKAkbAt/RQUugnNvTfyIyiWE4k5bf
k9/W5vew8CVnquOXE9vyzI5xGFEnT9ljOqJBC5R8ryT6XsYQwBMZ9AojAn/J
DM50pCSOJVtjLcFpZLCiVAEyvNPJ/svn/V5EvUbrZhGSmnRAlAmH6vmlxY/r
nZ9nf/O6MkvzfXHGEUaYkP6A9oOowwS25XpcvNba4vLECUpzNEcmNMkP606Z
VKTIwSXE8DTvQxpMQrzM+rrR7p86Jb6T9V0TGETur1NF2rmgILNAcwPx4jxS
wNbz6QCuIGcR1ceOrrmRQbMekieF+cmnBMMVvc1mEHIT5ZI1MvKKTel+6yyA
X8F3TK8cYzHfLAqyUfc/pWbMflQN6Tu4HqJhcpgMEhlUPmF6pkQTKcZHpJ1g
Za/BdWsG42E3UciEt3m6c3I49yWaElr6gefTpxDvgEPhylDZKmAHBt/cSsl4
7CVyOtx7YJDoDSqjzGvCK4Q2x9AysRBBm+HO4K4n6yTCKLQXmrA2SSztcLpD
3oCfv9ByG1RTl8DAT6ue9D7Hpu6G66H8Xy9nbuZ/lPPaDBKZL4LES8xK1mFL
KAF49fxqluffIMMLIF0vwNMsaeQX0JhOwnbx9V21c+psexWylKDtWdBtn3EA
GxAWq0NGgTnyGHzJMQeZKZ7sghzCX5NAzb44ATsbieaHdcPABC0FXlX6ep20
Ytr3KTCDJjdUrkR4zBETaa2kMfSjZ9LUsMg2tjLXZsgeHYA8wsj2/3XmucTE
klUCxdcuUNj+Q0x4NTXYMKeMLtERSMqIXG8bxNgF35AZXOr9NV+6hdBWjB2E
gnur2xBGzH1t0mPGmNFbdWummwcso+fIJzXJcD1FEmnQvP5MEwjQP8N0h0zg
RJ9gK5UgTpJQybXXw5U53sFXvDeHPE6jDnoxFMox1U3TWpkeyggpUadl6tx6
Tx1iUd3Os+ezci0xTwY0wMthUc0rNwxH2QPGI9RgVrVcnRBzEGtRQmxGBUQu
tToOR72DOkVSE2Q4UyZj5LYQU5NXmc6uHK/A63MZw/MRJcbVOYMPAtAjhUK6
vUbGwuO97IyrsQlAiMaai+YoqjgbLV3Fzy8CoVRIqTWjDFvx+cS4GWlu/yDy
ZPUPZ8CNNVSH7EFjf6bH7TDcD0cLwJzhzJ7Bhn06uCD1JLAOzuVD4ifh9xOZ
OddbR30WVWSigaO1TQghQD2HLIneZvC7+kGAy8pcw9LxlgLQMK5wOvttndEg
oglvIeBzSrI+tDNYHJRD5WXlhHXN41ZebsqMjyLkCt4qESdfb4/61ItHasD0
HIhNv9XrCnYltmAQqvCMJNjYGD0eh9oHYjI0ef9LLMBLnllXlxmsQag8SHP1
jUjLRafRdmjEmPmIoOqWTbrxSj6QA9ZJ600aBmUbzF6PMpGfxLBB8WYuMj3I
PGQ7H+BVpKx5Hsl58oOVA41RwfM8WaSRQho7+aKbxEsc4Lo2F9VdawjQq3Z3
gIYDfmXjUOpIJYTIC1D0U8Y6Ths8hCDfi+uj4cB2w0A6Ns+vy+p8RpcJNYg7
MP9uEGV5AOmYhDScOsQxfLT0pCPdCKqhE6OZA69GkjgX5ESid34k9saPiMpD
F5PJoUGY8K6zSFQwhkN4vLxXQT538TAvkZHVbb/Uhao6qHWz9tX7vcfHhXop
IjEFeNs5OtedlLudvrFdj8kiYeBCyX9DI39yu7Nzmem4xQZmUXLeusE6s6X2
k/sFQA2ZCGm/ZSJyDJ2NOkTMLJXQaK1a4HUXHuXWf1XYLDUnb5Htfl5tTcY1
EQyQG1DHpHIutTRaZjLKTCfJ9d9I+JuRJ1L93rtEw4bOdxtFjrSTAxQCwDxc
KOICjak80Yc3agPF+FvbZuoEyytwOXHAVVQw59tByiRzXdazZsdWf5ZSw2Qv
jmi7BY3ACQgP72giUFqO4AUp/E63E/dgkuVmUaHWqGBFo9V90qaMDohW1AdR
0aO4ebElecKZR6w+5LiK+vEhukywafqqjnmOXCUxHdKW+lFaUzfsTZvIWDRj
y1nbRiEOz11Wph1PrMzLt6Gg/BmrlkUSs+JBHtanLPIH4e5P9qRNjoVneZCE
G4sC4vGDf8X4va/m9vrGyVcrx6CsyXTom2qqenamXN1bGX27WLFvjTUG2JbC
SM/v08ofLoCrwF1Mhcli79uUnhgiBb+Z0IOu2UBNPJ+ix/7mJbv7YnyB7VnH
VunCJ5aLkKEPjVC6iseV7AytKbck+cKDwTCM8Fl/TTxDyvVw327LcE7fH25p
EyIJzkWsejXScQbs+IMhU6p8FpPgOQCTq30G/pqCnQIcEsVv0raSwx/ZsIWs
sIzPvtRzIDhig7REpRqcF+qIWR2T5w0C43/WqAHXhaBFxkSLl0EPzyN1joK0
jO+sjIN+7iVlvmkgds926RXcDKde0O6CO6pjv57PvRMZMALWkNw+fvyfGjjD
68lhbEzUWir/y9WVyx9ZNz2Y59h6MPnv1ikkpcM/BwBC9lUFdGzAkR+D/OIm
oe9YsB1aGhysRnTEsthtjafTf6KEFgBf5J0XvSGw5E0YBwkZBA0v0lMV7kYN
JyhuTMinzjE9I2sTY7IYnTXmbYqQJFKZfdg/I63AkD7bI+/WFR2WaJtmwFKz
T1iMJYjwODKJ6TFv8ZWEQIUKuSEhTscme4yRmNd8r65p1huxfhIAPLYgQjxH
Wy3NfLjGB3qC6SwIv0UZYFcda4wykE/j84jt2qIL5X2l2B/tQlt1zHATDwSg
I1PP+CXnd+p/0Iqzq0BMqMzaby/L4YBKFyPdjlr6VYNM7Bxu/8teLyqBA++k
83DY8iPQgLqbPr/6gVgt/gYLZ2f7eMJDYGNdoy0tYgvRVfw0ryQllWshPZ/b
sx7IV6BoABl4nrrHrUHlj2mi3BMU96YSXp7Z4I5YsE6RmCgvufRX/+YVSFS6
CFUbkwKNRxt0uLnHKD0SwyXOrnhEVIuHzne4y0SnjK4Ydm09CRzgHONOHjHg
rEJVEi8Gl5HYC98FRVMhv3spvWv4kHXiDRmhRJrt9u0FgOam5tEKQs3agvVC
4kGSxP+hCyLMWFNSpKbp3UAmd3nIBiuFBnn4nzWRsg+VxgDyx8GVeZ41zBed
5F7wE1aMKpYvTYZy0rMfAbchthLXnn/g1aGLasIKLZEoFgnsMyKo3CFPe9+5
nu1jOEMSG/EbGaOal5T9ufF2460M6t/6ow9z73eyVCJf64VqzMCIYYPNcUWK
2ttqkA0yzd5+dATJ48FlCaVY1r38zkRcgbBz7AAtj8clTyMUc3d1iYQ7fACg
Erhd5Y7iTrV1uraTRVNNKImJfOrvFfAu80XJN/JWTg5ExVMWrgSIl7L/CAz8
BAc9WABAlz/mZq0SCbPXwPCFw2gc9Ee9HE/1kD7DTpAYE5Ac0Yx3krVlu2wB
syxeioaTGXJ/B0kVzIR0Pd2o+OL+Dozw/i4pmrC7y9Z7Dvdn34uh4knfDFX1
jdN5KCDSIOqQv34/hPsDy5+CKUK9Z4ZhE4jq7wmkJrYT4iin4psY/7E0GbRZ
SLlRZZ+M04z9ujl5JQc91aF6cTtbNy3JhJzbVeNBX1HzRLgVl3ZLeP8yuN3t
JIgyOKMnQdnU0/wWPxeN0ULC+A3dx+JOHJXzHdUH15aG/6qRNdoyZcLukRjS
BcuWdkdVvYplNjoEFLDslDwJhK2TtntYg/8aKBBsV9cj+FmDQoXaCqBEUvfu
TboxoFp+BNxvOmX6c0Z9ciI8+4JaUatON+p7pDA+8JbQn4TwlotFxFAjKKJV
6w89KpkJCnsLvrR/SBfAhDg12icsH4h25bP47WEcdrNzJ/+GuTmBoOPWZR3R
q906cq70Wb+E6fVUflv4FYR/IkSNTinWnxIuuUvtYxe2dfm8JfGh/01pEPw7
cOXkpKtieLkIw7s5VOyHu5ByqfqlIhTlIK8Y7VfHcmBlK7YozSxLGpOJVSeQ
hsBmMtHh8uHrpa5cJrqRJTxjCthY5PzE4Cdyg+ElTo/JY69XOcJHd5srd0Q4
KsCM1zFnW0f9vhip8G7P8d+sjywRU4fQKsc6b/jq2+mgG7/Fpg9PK/kFUge7
Gfglah2LkftA56gdW5NfOSaVEuIz9zqR5lG7G3LImzErcPUOYvWrgjA3yH8Y
gjqbdex9Y9d3n2CXsFW3XiDvzOmFtrqn9+BMf2n+oq5bXrxypYkvHpBKZGLC
+lVYiNEjgFPfKzVi3jXkXLBIuv3aaPloeE6aEmIu/S95jA0KzZvfVSn+kYPX
VUY3OpbbWriO6f7jPJIoV4FQZlOrt2UXLQRSGt8FR3T034yF53PlCSOTWBOQ
dnAjhhBnOxTPHvTJPrhdyVa6PdZ/EFPTayTu82l4LZfMuI3WhhDwOlMsRNOn
L/x/oRL1MRZFklMO/TfNzMzHiJvI4emjKVyzwrUh51oWD+CSQpNT9GeZ0RPl
DWU6hrBfVTl99k7mjDieTcsQcBA8BRFmQ6SHUUwv22lVj6d86HCWP8pB+8tP
NwSQZygmsC6BIWiGtQTOdyUKeeHMMQap5nDSwpvOL8CFPblPwKnbjbjuXDpB
XAp5FOWokdemxqOIjUptcSz+bW6tE8ngx8bFm8PUOI+2GrIpSnRfL4kYe+fo
lC3ktnxSBwtcQVGJf9MD5QtyYHF/G16ObJI2Dl1Mx7tcF1V/awS27NjNLuAY
3U279OC4900n1lYObgflhOOUL7YB72v0RZGEB5cQKmz8l7nd0/cbNgqE5B/d
8WQ66QrBs0asKXBae/XSsFPFXVlN9fCu/vP/UFaeDZv3G3A41T7mYxn9076V
U2astZ1Auk7puarcX1uLMUgSYVl0z/7Vtf0aL9iC5FCaVQ0AYnw8hNJuAy6Y
ww4vcPnIB6D0wUNFeqgzOrAUOXvLtjry3gNlEyZWwU+nZlVgLAgzowCCxu9l
rbicO3ultvPxIVu9TXQ40sHF/myowm1tK466JWgZV+QxWb0SQT1mv3p3Ovcq
CVqNhg4MSyGUh5q5xr1LvcNQ5mvpYVODCzRzsrV6IyLLyJdt1fDH+d+v9p+w
LbO4bDcbrp1BYEn83CSjn/8eZ+t06lmdcBJDyxVWPiS4QDZ50SHHuYDnKYad
9yBAc0qt5Evkra1OQJUYGoQ6ypUoMCcBMhTiMNqT9CA3EbnbrCH8oiqmOhdM
l0Sza+ukSG5FhD+2OihsBUiWCuvY+nyHpXQWuSaTW86cksK3qERdtrea+NdN
1xGLmTLCDlj48qzNK4o+dKxAUqqI6tIVHj+5Qv27VVF8rz3EDG+7tkApyhuC
y1ai9bpKJztZFcO054XCnUgSHBigbKXlSYSL0Io2C6U4LtAc7Eq93k8b2VTJ
HZ3awCKBQ+lLywGHwd99jMs/IQ2Q44rtGochBVLPJ669X+YG/2ETfp7VVoLg
EM7uQJP+XgKUd9xLfJndal3wpAXttkIWMW13CNo+By8b6egd8EofuVaBXVJv
QBTRchN4GCXHmKPPr63TbwQzaslSHXZ6IY4ohaWH6rInAor7D3fvxHNLgTkA
8Wh4Oh9WdLxl0einPGAMVA5ZVWEiHBZC/7LvUXBpH7mrzTt9mqEx8CpL/Cm6
BX7RTIHqtbOa1NUGIIZz7TlcTnvo9g9K2NgkO3wfMO3x15bAOFF6USGEqHBT
iEdZXjTAFZVTbWpikVQr68j78L3ySZbWofgzrYdpYPwLLvZEIeAqd2U3VAQm
zTzIID3hmDr+C6009S6xBx6/SLkZXzEEsGi/so/2j3N3KYyoRlzP0T26e/rD
N2tZLBoRwdrG/D7Q9/jWP1G5YQ/JyY8vi0+iqyaeGS/NDfzeOmRoeWk4bwyw
akDbDsshaVv1/BizhHm1o1I7nlXdssoiBBkiqav3DN9CvtKC9p2voQtZx1tR
1Nu4vhT+vTbC+O3SHajI1pfMeycFh25m9FrbLlzo72wIB+POl5gsTBo2ZtP/
GJanOAtS+uZ4CJzY2io1eVmZY3e3AtLxKvsEUDrn20DATp3Ary18008JdgUA
oqD4o6R0flo2HQHuf+uT86BM0ZeYlBnWL3Cxkot/0FRaePWahMAR4H2N+UcA
HgLf5RTrxLSOVWwVLXdh2+R6NQObBeBI4JVmmYNyM2wEiH4dAzJxrDaLChLr
ixEb5XVjd2NM2FnOOAXUUVoocoU90lgDhUEq6VgY0YASPBBgH3vM/jKon8Bi
olhPZgOIAg/poD6WTWbvbG8e+poeZTzV88+sqgHcMQcOmVuuqaSOmuvTT7AB
ywpEhKCDsomFGYNUeCfJJj30B9UwP4N5LOlFHrHrJsBIC/dfKqdPqVwYHVTj
iE3DDzprCPFIxhj65a0dPdCcvzxPD7NBw0qIEm1dEyXl967o+u5YaOjeZyqd
nB9yET4kVDtMEI+jjWyEjlEi+IDFjMn8gqfe9klOWETNW0aRKge/1AoAKeva
kLafzBJCRBk1bnBJK0JZ2UUYBlFYQF9ulxncaVmxzyhVmSWRrT+LSzz3MPmm
0CxbAyqZg031tRFXzETMTwNwlfQ+LIBI9L5lKPZ0tTflOUmA4TZKfEP+aCJ7
RSDSD+AE44HrEG5ozstYX/Bhg4i8OlV3kBAV+8nu22bIIW13amat1YIIzZgs
RhVkYaKhcg6SN9emO3mKrqhAhOqjrIXiJ1F6GMUBTer+8SBE3oWLhpl43xW6
ABiqqdybdMujQuOHxlBoiMP2VGOY8RqBBpwhsaE6fPToIzWsqRuXwWXtYOuz
KpWFj77Ps22wyxy3u7VxQuca7lWvT+reidQkc0yVvlUaqgxMsd/bHIMBVQd3
CJZbDld4rE/kevCmllXBlhlbqqB0vdeyZSSoWv2c/XLpTuuIHWN+akU6Q4lD
zi5UcQ+kYaRAbfb4EVsKI26S01MYMugg/p1cxluOVBYM45LwfgAsGQBSOLET
K3i73Fik6gA11mnB2Kc7Vt+QgziOLjSl0OQ87YiprfHQHudiVB17PaiXjANq
KAuvdNNmchfvNoh/RZe8RPq1vQ2ls22DXA/KLVvUSrpS50ag9jOM7NuRTfdG
QIm+yvj87MMnuLFlol6yFWIpr4xImDf6iq2J+XJFt8tO25D8JYPQ9LPJMaVP
CVItv0RmfPLs+QwZVd7dZcY4JYdDQvSkXG4Gc3B5jWAM96yVAobU8/rSiItQ
HGaKM7uU4Gi0Ny9E4xWL3h92uB8CqPdwn01WzNvwaHJlaHKczdh2w4D0MXoM
GKw65kzECCDKoJSB7ywI3Q4/8Xb/wsvAFNCn0bWKRP3BbH/+WdXtlqkbzODx
DvJz1VLyCFF/WiF+1e26/seXXTX+1XlNgSLdWCrUvOd1cJKGQQiqbyVrnGsR
FzW15pENlNjCollcaR4ISRU4aku5we2IoDBFNi3KQQX/TWza8x/lfO+ZiZKb
4qW2282gjQaUkkMHFmtp6vubNjDrOo/un6RNGyBw3yuckHUJqD3O51VgCm35
MA3IkAlI7w/ishKR1Jy0omaqfSddGPkkwciaXHfvWVIl8KpiT7bJBzYHvsLX
Oxsgej1o3xfSMS7ObadksCKgqK37/8TzjRA76/zO3VLDlhfHs7UMRWPVLtGH
j3RXSmfGwcYIMFu8ROPt98QfVcJ/tclwWZaafcPNouu7wXxOerqbI2TxV37U
JXodPBijzlnWJPLf7Nye6ZT18Fc0+MyvDUm1hSxWlgrGTpx+4CqJ4JOaOSS8
OSZB7DKC0ikpQFdzpaOkFT5+sZ2yWzqqjMWRBXBSzVhQRIw5OvaVBdqwVTC+
vAREVUOTiug1otRU5HLwSh1RbEAbX1yUENbsQDlhUj5x2Se8PUugOuPWWfuU
QdhoHgjicjrG2Qenog5DVRMIL3x2vjaXwqmmwfSxPY+LWpuqR5birab5kYD2
MABq8IhFr6Xe+Ze9f1H4T0M7IqOE3AeGZ0W9wDdIO0DQx8UfTBfDh8g5EXrW
ZI+PbONoZPJ1DgDfkRQm2obgjFrvwGK07A+QRnTb0ZKsgoktjMWHMxak9sX6
UaQ3NPcKz4olk6420HSfbgk7wQTTzQDW0uMt+xqlwhiMW9Cekmf5PmH4vqHi
M+LHEHWkIBKz8Ts/Lz2av3E7Chwny/cHk5WGUwHenOcrY+DBg90f03oeAw8F
EKyv2gV6NxTcE4YyguAXnKON1JTSft8XItZDZRIKQ8L7uN+guKYO4onRCocn
VZtbG2lUSQMMnmhx7uI5DtT81lLuTT7Nr4yG/77p6hW6ocWI8rHwUIwUR7w9
aQUiSDMRLPM9gzOMWd0U5uNKa1k3Rh9kKDp3F8v++ZHXQqEJHGxO4Ndo3epw
jNdp7UXqNNvPKkEALLgfuKvAkyQ+Ln4lIhUZ2TQwqijXf1rL/zpWGi5bOzyV
emOLOqqQl+a21uc9wXsh2OMbqQi/O7AKBiy8lbdx/1gzrHwK7fah7XOYFCkA
n4N5h2p1zxQVkHZlcgeGM4GZOeKGDBLNl7VGmmzowKPrcsMHUIJvG01fz6Gb
2POFgN91EHIkKoP0ioFvrQ+aAryVZa644g3RHhpncmirr+W4sbUBt5rWLU4R
mg6/WKieZCUMK1n0gKoh/yhMZv+GmJvmbk9x4IydHL5Jy36JSBI6JDsZr+Ov
t60cEkpxq3OJZoeIB7viqRWENnGbg7J9VEksw9Q7hYugNQf5+l8i4E2UqCwi
1yJEk8joRp9FsM/nae6bP5fGqqGoPgxHuau9AMkinRwQcHpBlSYL7Up8+CSj
6I7LfIkgKWMTuaF8Apa9A8LTmYdyusHBzbQMhgRfLlggAEPy8cCwnnzjEsXC
nR+3UFkdGwjsc44vCpoYsPTn6J5J/L+U/PSLMuKJYAEQKy/QPEgysh372oyU
54c5UP8jXUxMDe5jqdJrwO0hCwAY2B0xvfakD6oEbyTc9VhysETavogNR97d
hF6BA4kc5KNwq1dVS+XfaHOWzSn1EBQRUrDDlUU58ARljzCs3hzL35hWSC2F
bwRIKhQROe1HzQUsOnrR7sSV3iqwu1vTUUSfxSFL6zWDTI3gkfcTMxrWZgJl
iByjcP/Blz0fLHN5PjYp7gsGJTy0Xayk21McO3RguMXxPHJYV0sOhvbuwzrk
YtU+cvXS8+k7TahwIUiXtErhUsnvsipZEEk4vpvltia3YpB6+rAPB97vvRUq
LoLcspejfDLcU0O0el7dpYr1XnHH4OBzMpnWRY4WT6fuMjKUrGspsKp2km0c
JOI3fmuVAvziE0cvdYfmxkvrbp74tegCfm6cSfoTVfa2Pnp2HpmAMJ4nDAz7
EZfuh1OZuFPs7QcPWC/WaLwr+Sv0zKQ55qeWh5nkmWKrcN2LF5gERb7Y4zXl
UTkNtQB1WdjDkI+YK4qSf/Whok2Ym67IVj1LZt5lPZaBetFeZwcgnxYNYM+y
BTCKD8PApG3HHE1orDlfHlWqN2OlxElaUWqwROJYKZZWAMoJj8UBf6l6a300
19pAYs1bFvbDvxzCJpnCYwYRicDkOA/m5MwKxnQUz62Hj/aFPIXX3Xrue03L
OMQ2cxeSFHH1R2J50Wbo6JKh/eyAKnmlnw2E6pd38utjwQoy6Zd30n5JFEIN
Tvo2+Qgh/6DDo53qbBByLNLvoYgNmg6b6kkgAraPadEnJp4Lth+Xbdlot0+d
/+EQqhlD0jZ/iv5GLUmNZUQdTbZe+An3dxv3/U99YfEmIU/GvnllE76Eku7V
mZHrDlfBZLaPkwd5jwUP1ZCGl7OGV2V8zkrrcKaI3aose3/YGePCm5a5tZjT
F9sTlAbG8+0HQbp2NZW5jQ6+hSo1H9iW7KdQ5HRiluica7ztzFwebTXjpf4g
PTg6pefDo8mNLAVa1/rgckf/RyqQaCOEhtgT+5n1ceG6YghvBwVZewRtHmdI
KMX9hCStDqmB4/OvfI94TBfMa+37bP+KLEPVVmYTCltfVVctv2Dh+/l2cd0Y
Hw5v2qhce3h/hfQyukvmLT170Qz9736zBQgP2YCYRGvb9FQ+gPFDlowY7Zi1
3S3N2HaVnZTW7lgmlxs7IO3DMJhJeeddDV5/5qO6eRk171EWly5PK0n5Itcn
nN0a1PP0uo04P5NrSknAsNULVyhvtjAAz5/O6CsO2DB33+DUo19klmfNhmRC
d4vP0k1bPQBEn1BlrFpk/jZZtF6vQW2Mn6qrbMJ6J44Bd0kW564+xwTsx3rg
Bu4DZ+WHMamRcWT54rLVj0VduMBYcq9fSkmEeZjUCbV5c/s0Guca5G8EUla9
IzF1vO8v9RbI1hhMhXtOB4tTczpouczOz98XFUevrHOJLu7TmjI6OnLNnoeH
WRbTnKNWnHl32pBeFd8N3qY+HL9DsC4KZDUiYQmj/DJiuZJWeEzA3qiQcLMH
f6TOQldgC2qT5kyB39xGnLyyN1YRWwJ1sbuy+GvhEDjVSFMZWnfvb2F8LC0t
qP2WbAvIkMllj4FhaBvCVY0M8AP3wexafdit11hzycfHgEE60FNgJm3Kaz2G
1Tpew6R9DhrBNdHIj5i9Hl/ulO9oiX6o99AMnkdvT+fQnNuclRW0CjK/F8sa
2xZvqoaW54GDv/68RtzF1LYZsyjRp89enSDigzCnAgG4/eLFP+6HF+JEasES
iXGlBFK0iakmScya2nd3XM5If945WCK72y3BvENvhvEYONdb/Smldke7iA1s
01tt+NRWbuDVuqtqg1V/NyH+AgHrQksR/BcvR8eBwBcLfMxbBN/nGrW8UIop
cLbJzrpZOzrwsKlksRACeadvqTsbXnjdIyui4vAKde5xth34Wtix2ie0D+ZK
6j4oGzSi+I0fLRV/ATS8swRFjNnZgfoPYuuIGxbdcDPTF0zZhzc0gsrFw5Wz
JcJRLUMagPm8c70UyR/ZUIV7+lvrzS1O8tB7iMq9Gz8etgYrbn6N70A+EY1e
kJlDVeEBHE2sNF6mzP7jRh1KD5h9FdIywuQ7seWMnztBgQNytEYT8XPF9F00
yJkkNsGHu0wmXatQEZrTk24aNokz+ZkMiML6gIUlDEf4e+TgFyfYFO283fHg
h6T6kMQHVkiFzx+58nstfLeVF8aX1DlO7YJtEy1NyTuMUz9tRYoXPqXTrftq
8vXbIIDf6VpUCcTTErzLhIHYvJ6GlYIdqWdiKvLaZ71XVVnv8ez4p9LS62vp
BLhMHI9Yyg750Cq0kv9sMIqf+Vcu5bWN2fQvIqLCXHq2wg+umol9dC4Oiavu
VJt9+GSz933DcLW59gEWGMUww4GAJMb2N940woooL2cNM+IHgtf61ksJmn60
B3cfV8nRlvk7RQydRdZmoa2U9C+4uokU1DBjL/HL1PqHHUUcig/bjDZVbNCM
dSXCiCYBsej1smac/sVpi1/ItUgS66X72L07m4WAsp7xMcfNBr/nlNDykCB8
mrzovhXUfE1xLZBvqm4GhSZ3yyTicGC0NQ1vPhir2DL+VgTIqUuBjHhgxtQ3
cKLTMjRl4PBdzndVStQ62dnn9vlO3bUflMIRH9FvgfftuZCfCHsV/LVjFIxg
JTr8u+PnVjQi8xVkmlA6VHG2dwIt5i/Zp8YF1x6c97gMTNJu3n3S49LxP6n5
6BIag8rbJmeb7NEezGIddxEvpaNknFvIkLkqD1rxMDg805Wh6tgcKC1gMCUn
szEEjz6W/8KE83bI+Zp/m7+a5mdvwhKv6yZrTtJyXOXcbFiSYZgBp6apdoGn
9I7t2QFW97pqanURW3nSao5Wc8fqT1cN/6Qb2DakEwwbsEINEwESRe+GjzGZ
bu4jR412CWlmqMdR6whSZHdultWs1mpx3lBcWJXub0/xKIOL2+PvH48/PDtz
ZoYgv76uKBUAPNEwID2h4gGbRbXMjiHSu9jNU8doOJvOZUCKatEg3qpIArBS
3KNsJ2XV/FqwCN0TCl8QeSCemz+rNWQtS8ajns8SVI8wNXrDiT8b5PD+C6hJ
538Z7+bScjsaw77/KKbdooUAXN9im4n+U1GzbWoL+o1QPWNzACtcL1Q6U3Gi
DWy4SBfXz7m6XbBEg675jfrFtZQZ+6LJiza/dDR0OPvrljdfnweBrOE94p71
m6qok9PpPnfXnh4mMDzlreHvfzA8v7OdxYrQV1ekYFXcwsrI/VOIMFel0tuO
PP3bqnUXwO7IVOFSbhJ2RGf2gnjiA9ukuo5246iYxjPTOI1PQJhfXvz9Oe5M
MgjFlT53wMyHMYFNPhM85J9/BQm4NwwCgTOVvnrmmQyP+X5T/aUUhO3pVK9m
QAtVOzr4e1Bl8Z1G5rCyxJc2mg9+LwbT6s+2/DnkZvigXIb9ernxgYMPr1Vm
alp8aPJ9zEurDb1igU4Lb7GfGg9rggWYXUfuqT/3FnpE1Gjiz7MO+ztFmSyR
PqU+weKJ028QGEU8Zq7/swoKQoSx43bsZhqUVWFjpr4dcayD90uH8O2xO/cB
OJfpfkGSbZaR6gnSax41/PkVxZ/7aYq9NMmXZGFjR1f6wNj0ZSV61Qk8NSy7
EBvkNa9cZQDpcHqngpVryJmJVIg8f0z93MrGpuSftFg0F1e99YOkif3Tlm6G
JNs/xXpgGQxdL0tR7FQwlbQyotw3WKclq9ZpF86PoLH8hSIqckJkD9Bhrt41
8zX3fWkRgWQWeChII4smOh6GBCzUDKDSPP0BVasIhGFLjq20GHOsBZ5GS43+
sUgetxjCRGs8Du1XyxfpIATk+bv3a7is2IXjHo/MkWknY+OTI552dnQzJh/G
nn0uoHNQH+yIpmRVGgjpX4Y9ISh88VNw+0KMZlhgHUd5qZA4e7PaFh3LGsAd
ioySaIPKFXOjA/8v3PFBRB7j6P0qnG+KmgO6j3b14xg/eun3YKg/yoP9C+1e
26lv2U4VA9yH/rlbWF4a19oYFD4B3VgeUkdF9sZB8wCUc+Y6XqOm4AB70u7+
Csw1WoT839BA+NSHGAxwzI6hQuxp0nHI/V8MoTBmQuaM/LGkxhWpM3A6hXxr
NMKHb0j1Oj6hWimApJi9ry36Jx0iyvSacrGt3NvkTdwjQomIgN7wcipkGqvr
9owC7HlftP7aU5ammy0rfmekeUAy9THv3dYij5hIgX8lVlY7RTXzS7mKOebi
HeeovneRsfx/con74Glzm+zILzrU0xufiZ3oSgzzBCdqJvR8t9wB6CWOtg8m
0jLb3JHDKS77OLPSvGonWavZSxiTnuYM6bxVdQz/BUgeSSPGqJo1AKRULGJE
8fVa+Pnpi28WErh5/qJbtHCSpbLupJRFVI6pXJIc5pRMcYrD85xnfoOryS56
JlrK5gIjPKbf6S9Sk5M4iPp7KeEO3HMrFf+IcdtxxAPP22Hng+YAkhZoEPu0
lS01yjIiUK/UomUILEzKiHMFCNx3PIFttAQEmgRCr0iJ4jQva+JjN+gsHbAu
co55H0WQ8Ldl5YOj3HRs6Oi/JH4nxdcloxwW7c9XoVc1R9ibqf8qyr0HiN0p
Y7S9GywO93/1bF41OD/nFkTkjvX9bwGuy++Qc+QZMb75GRE/kiIJobqgKqAR
VgSBM0+NkOr0QNsFfGUbSOZwMUwxsEh5Rml4dLggnCqeKNz7SgMvsmNNi6je
iZyghgvkV4wvEGbQxibTdGJQ1f60W9e3ITRouCyyOKN1Yx/C1Z14RZIvZkCs
iJw3iE8uSRQ8Woz2hvO+7853N2JlAuvkSgsgED2FzebAFgwtGAsbYN0ES39d
g3Z3695LXMzhEuFri+U/JDw9Syg91nSAj0A4igbEffpPvZNRVMCah2xUgSTU
0GkSF6WA8uwziFLhPhNtozePfQATBUaZ++J1zkaPv3skOz3JYqmqqXy0s1CF
jcLNUa3CIiJwuN6vw2DbDTCsnjr34qzmssxI7FeWEdQn4HJ9iuGkJLNqUzqW
kjaLjIxXQJZz7/YFxI0zS5qiqtymon6EwrNXjrwH3lmNSftHk3mf0yZYCOTG
Ar+yvvHOl4U1fLh87ZO9iANoOm3NruDuw1vZhdfCgDoo9SEkM7I9ti+mTp7t
wgfwFXICUekI7ANjfHAnFJB0Vi7ehhyZmQJKJn6lYyr4DsaqfUulkTZ7DI3T
Du3wFUoIqHFK3h8CXIYDFT5u8wLICq7l5in/FC7iQs9cvurrXqgYSB7zmyNt
/bcp7OZei7g3LFAhq7++XZyVMo8ZXsh2LWWr7UWqjBxISZLBd9xP7ZOak+eT
zdZ4qfsr057DEfXetd4I2GZIY4jMa7WCZriErZ4iQ1wrU/NAfjAZGKa+JAmw
WH8ti06w1CsniFCGFfNHL3M3SRfM7NbSNSOK5Hhr07R433cbuNyUA0mHYze/
qGViWayOGH99PcFiV6it58BgKy0oHVXeRcMt8USXUEwRs2aclYQufMJH4eIJ
y0A9duKRKoQEUs0EEfGDtx4De32DKVGqni8XC3iLiHl6iLnsw2U1NSBeUjHI
c9HWY1W/o8rID8yg08S41wzzjnS0frH7Wx2ciB63zxXdEfr3TDvmPOKUZr6h
nWu+LvFiIwogDx/gS0VXLkl4iqQAzudZykGkyh6Wn1eGSNNK6DZa1W6Iznmq
236eYVyXT8bIEMGNHZpMW2Vm6TPm07zUJ//T0CZah6levvbFKv1yE4+nx6BB
qZdySR3b7zPWs4Pqo1i2mPpLIjsPlFQdU/BY+PDzDS3puIDApZkz2CHgfOk8
0BnXM4LpUkqpxk2AbHM0PZ7egFgIZ65coEZ6c/nAyCqHO5GGUflFe6rD3MqS
0ANH+cL6jtKxRQGQy6VZLm7PIMIIfjvZ5nC3slZiqoHtDGHbFVqa6FnSQKN8
+AHEDMcRfoWl96D/39gKJTzlNK2cibNBD+68pB6qoV72whijRzL1J+Ds8QDd
TO+2xJOW8R/igmlQXSEZ82WjHNGNz4P6nUUEZpoiG0w5YFb7sQT8ovkBKbR5
bFtE8t/p80irgCogwypbCZLINqbKGGfYtzQ3owYZ8+o+6v+MCJ0oD3rqSg0w
xyM8NZqRvuQ2i4SolQpKUWFCnhTJdLmdWj5t8uZnjNiGszHkksAt4GOmeuV1
3VR9StY2wBf/fUPUte9bFa2QsUfYR/lpYVUBcIXeRiqTwhENtn/dwTWB72Jr
MAsKfS+fQEYN/h/dC1yovEDMbwF5nbE26T6zWNNAmh5SpvE9EoONaCLU7m+e
LLMaFNGRVg73DivAyJSVoEtN8feq9Zyfsx57xtbHtv5jWLdoY6VCALmbxSpe
7FSyBNpm/l6OSdsizVAhQtnXy9toct7z1yw/W6u+yAaXFvKyliqOXpSatLWy
mb84u9QkM0yp9+4ZHeMaQnc2edNaFtIGnoEloztex2C70U+hQq7ANh9XUFgu
af319jE+mm/UzA/3jLtmszNY6Stlno02nEtoOLyFKqKb++8BRO6JaibMp85C
al8K/YHWW7wETtqIo6VaI5kdH6TcCwM6Cq+/q2O7Die5N90tqVklnLoi4W+z
L3dX+ALi4Y5pWizjNvC3LojEUuYzKLTXronlxMMhbtY+Gz9F6IagSaAlWsuL
d9x2iczX+KiebR1YSBwYmblDK2fma9mjTAqphJ1yaElPwsagffeCAMm9wvdt
ZPQHZihAMTx+yI5q4+A2PnJHvSHdSHL/5Jm6Eel7aiqxrNt0vo5Go/ZU9hlQ
7iXyNf6Qcwfxn5/5zDqw/dZS5ZN+T2T++35jND9amGsPGxPw/yUVpRCZTNfF
PBJmCoATx8KyHq7PoRzMVI0GnP0xiqb+YqXWd075vF6//zu1uyd0vMSHfCWI
yEInrdkqQT3FibelaIU1tCv8YXX20qZvSJnATJLEr1CuxPy8E+rA6rqRewcG
eqqmJ6qp5x22+X/nxT850Ul/LhSjFpzHgQhcKs1UIMevFTK87ANXR4mq9l89
VeMOBdoVseIcSkxVNDuWGmQDpDK7rjgKeqAIHRvwqR9P0k5l8mzoLIAOQ4xc
lNKVp48tN4tXRC+q3eKEgssMmJJ7kW8wFewizFQ/EkQaFpuZKffuAKuE/oOH
UJB4fpR8nPLfwLpknsOH/jf2YnplNXNiFBTWmP/cXDKPLUXARGvv3vIKrNOg
1P35MaoUIo/nQJUaKCMgEsswVRWDMEb5I7DMfB3aD5cmCWPBtSGcnaVj8+wu
aHmBd6GhSMTyO2UsWIzYrdZlYgZcd8Pg+JHMbirYqgpPZR7ZiW3epl71/aNu
e/eRPynuLkYvzhRmL6ttZs2AyB6Y33JKnyJ6BbHb8V3Dkl8o51BgMHPKabs7
qW8/oCqAzN0m/Uoc30dP9mpDfys6kh+Dt4gTeD6vvCR7lhsN8sMzYEs0v9Rz
bTO8Dg5aL6AJw55Rk2id9OiW4GR6gkLHIoHcl3PHixBuBFFgAMFvzsdY+Eqb
/3RxrejkpOEtaw7U4VVmj1vU469tUO/kRc17ZGm70Ri1RhcmI62bi7/wueg9
ixbbvWvm6G4N0Kl8oGQabwcIMknHy46IGDKVtJPk779i2wyMqrI9x8kOc5db
zQYUb+Bf+ev9xcfgrWCNKgbh6CXY7RMZIceI0kN9mK8zkQYPKbxQ/GqVgEc8
5wSbBaCrGO87o9Mg7XmS4xdNTPHMKufCnERb5eqLvUev+9fMt4ustFluZ1G0
XrAV2Sz5TD6/flUUEiiCJ9xj1+iHUb0KkzfBg9UjIgeGjKHqln/vfpQcPUmu
3dNn+ndkyLc/Wrrw3fJabI2q/wW6zZr+x7K8mylD8l/7vOUa+NO3527noVRv
mZKPNrhJed0D/6DfiYv7KBXCyG45bIpiVnzyNzmb3guIxf+PXBAjPXSpL4xn
ClE9EDrczLU4ZTBO5vpDydnihSw4FMDsa1uFBY/wwuGWlJbjh02XP2m+YhTY
S2Wnxh7vbAm6cWhXRBWoPcDhWtr3L549qRioT2ZgshC1XQe+BTir0n1rLUAi
sos9oWAZ8KO2xQ2t9n9d6vxWzmqOBe4/9JBgS4+lkH3DTCPfg2omr72D2XPJ
uSLpGlz+nxrZAIJ6H+4tN7rN2rG8hMU7UKMSo66eOsK518uEXbv3ORF0ULw2
IqpJVG9BvAZsZvMqWYi7kUbv4yV0S6QUSfFnCcQwuma4hJqIPscnG9eCqZ0Y
OXyine3Ot+c5MATsjjnW9Dr5XE/H7rEHws7KmealRZVpGY7kbc2wYnWT0x8h
tjcTDeFFmXUqVGrDKE2F2xXTvzSYHMxu7fmwLsj2xDE/vEOkBaiNuxRtNJRz
vdcLeLfOwlbGTu6muv1POaM4z80YO5eP66QDIK27bUA21F03eXRngIgTIx0P
ZIjx6+C9v82EE4BdIU+avIB84k3HnnfNzlEDnza329oaiag8+IaiTU6M50wJ
fCOl/ZXmUaTIVmHpCz9vA+I9DPPcvB3IfEV7HwmGZ1VRcW5NQh35tylV7aeS
feJX+gKNtbSdJoaNa0BQ3wYSTRL79wjFOp/1hSUcNPp8bLctMXtv0HckqxGL
m3tT5dkZ9WpXIEBVm2dW43cjdALf74PJhvEpWMqv8pTlcLeS82Da+wijMyL6
TSavpq2rNBm5kh6/YIbO9bVrNnnuHltcrkm+XYd3ili3fdjGg7yAuxVcgoph
fGCoQCUY6IeWKqRm7pXzft562gPRaXTw4exLlep+BeqTrpUakiSR4ln2dAqB
EO9fvNyMmOJ3DA5ek9GFwTy+tandCHvk7uo/h8AzPGy7FSfqgU9bUwbOe++k
ei6WKPLtU6aRux7alcooLZ3/kjYA+lggTojnya0wCOjyF2DnNMroRuv/aFbO
IIPhHTt3511puN4ZxUHsTaXjOW4XMnKM5P9VkNWjcqvdKQpONFA2SuQXqSHL
peoJ+Ni8X+5BmKv4hi7/N2w/2gXhKlUH3xPc+hAgLsodIKwGuORPrMt6O1Nw
9v7MMTyfdYoliHtKnOP7IJgGZtRq7G3zP4okVDwaXca/9aFP0tbnFeQGKej8
AGHA31FUvkmDGRvxOhamn98N9Dw5lVGhbo+tfNbzF6kOIwXVsYTV0/deDXVb
WeyWFa0Pt7g1Ib167e2KuLm6upi2DSsKHMJ2IGUF/5g0s7kP0Ecmr81FISpO
qN3AZTVdKwmvx7X14RmhpnY6s0WzFoGyQOT5DKMLaMt+YDQ789NB8r5sfLAY
+PCo/9qIxy63s7FgNrj3xO2fZL5pCzsMAH9+L2zQo/bwI+bq86g76mcNzkKQ
utdPM5dfaBIt9kSsnh4dV1cjg99m/jtcMoW0UPeMcN23dM7NYcVVftXZ+yeG
7wdrVghFVFQ+GEUAlEgSvzCqVx/9VfOzAv4cKNzW2L2gsUfa0Bh8cHRJBYPe
V4n41RGA8N00roAdLtHWqWiGq6pPITtM3po4vxEcuayJd3AiRpDkryPWWf+d
LNiJbXVh38IYtsD997cmLcCKhxFByN5QYLYUTDZWokspzIqfmX20N/4kBFvl
Hjcx+KY4TFLttYHplfR6KSnN503NxH0QNwwvdN98PI78yqT4SnaJA8jtlKTo
59g+PL5DB8ak2Dv8cmZE8D/szUo+bn3ppWLL3RlzSZn0sN8LEaaqPmZw5Lah
ZMZaAsN7TegoQgAowzyVX8oufqs8NETaDMWBONSjUnOe4We/wpMW/43ZXUSh
t2AdMVyho9Tv9aNujzmZRdQwEh3+YY3NYg5ss9LunRNIqM2vXUJJwhKkqXtm
SDFn7hf1f95O3xV539nCSlD7wfGM3zpv5FVvUVUEBrqsPLMVvq1aJ/evnXHL
ZAKtV6RJoKDmsdVMmvIIxrWKPgtpCBB4LTAsHmEh4KbMx33qwuW2Rn72lB4F
EXJ2APU5OevAG0g4eVOmk5kthlICc99SmNAhs6v1gGxYYAT7IGeurknQFPB5
tXnXy8DvK/Ue5xvTtPqxSq4ySKgKkMBks0/FizylvuI0JTHWCwdCgALQSHTj
nIN/Db/iG+DPFFahepFOuVfs5MqpKsMi6D6ZOVuaBKoZLbu29OJY94zxypt/
/qyOGKK/fw7HcNSsVLpQHA1U6x890GKnS4K4jgnGjn7s67wUbiK0vXzmhD7F
cinSSreUNqSYRRaIsMONF062jCSw6CHRaS7wNWAFFlVGNKwEpnb6io7TSHT+
KSId2BdW7kjM/K4OIiBwD5zSbgQ++9nNNpZATl5BEca1dIYHDwq70VY7BIDX
Q4N9ELPAZCUQgwSmfYt48oxT0185KBTyV5l0fRT7PPvXal92EOjHcxYIOrRP
onDQB9U3RdMewVaBtsfI7Zd0plQgZLR/kIvqUrUkG+Uwl8Z+QkbQwF7qVORL
zmwktCrIlokVlG3KNoYdyipsaobPU0IOlbkNB5E9zfEzHRRdb87u5JTjaxSJ
VHn9Kmhn+AloohsvYFO5quaw1OgVcEAwGEC7alp4ToP1XvEbOvnwvDGYA9aC
9FmfYTjVx0MRrM/H+dQWTnlE3foBVB3PHthMD8ZMw/p44jztuzCMLl3BvKzV
uLvcPLOf7NwH75fjZ2cMUSPUxrfI9EsUJ6y8tA3WNNbl6UQgKfLINptygb/n
BoxsXZbWz1Bg5QvXlbw2c9hVDfNHqlHGxdh4IdvJOwyp9XMnuX+OYg5S1NvI
pPhWxpEoWXcbBhLQsKHZ/HfcXVzWKORHOzsMJ49/coGc14SMvPC5xMndzEss
L0FvZOJJY4hRTcEIYOaYslLJ72auvnye3sSjvVe8JH6YudXt53Eja22DzXX5
AclX73gLBjAX/EVuzerWWwdeyePCtr47omPqZJoEzP+T4W9wLTAudrdpR0+x
nRaSPeCdSTK+VtYq5zfWUrclZ2JFf72BrBsrXmtMp0FpA15WntxEV1sos9hc
jMo0CLSypry0OK1G+aNP2ZJnU/8bvoGwNe15XRiayEOtHl7ux88rNaznivsY
/EIW5Aqhfum/W/O0Uihg+DmUSC2HWkQpYAR58Fb03eVcy3giEMnm2cU+JOJT
PJ7O/lgF+WGFUdOX8jjIb/SFhdKBDlyQTCNaH9VA80Gu4OIQ9hkC9cbknOfz
gZCFB2IxDfZFj+fVYvKz1IGV0OeX+DGgsW08baoV/jM4/ovKvSln7GFxFB83
dn39wqOlNVkbOK1xkmHfGMfbFGYfCC8v3LWV8OwhrJgg4l0u7wHPLS6iy+9y
tM3JsDd8RieI8TXSu0tRdvKblaQDZcMQDIW4bPHSI8mrvsY6zsGo+hhu6D6P
C+eys3rh0Why/ryitc4liwg3AKd76m9EpTbvcQ+UqB6qg/3W43R4eiDFGfSz
0GPNvHGUp1p5eE27PNjZ2vvVffLNZFjvvFDeru0hNhOzUikRgDizGUS2vtB9
OA5pgAtdnCsLQk6C3cDFc21ZAtDGXW7rltjTNguNjLKAJrz1j/O8rv/x1hTY
r2SYCZRhqIEk++6xHTQjlx0Uli4mlyg02KumQ/7L9wAtP+d5lv1D5A1bkQaO
p7d6kHujJX9dIJBhwTqdhbsklKY8wd27RLRBfto/bVQ9HG0Z6Rq4tICDJzjt
IKqIGWNVg+G0nkDbT7r0dhm9FXNed0ObUIONS7uAabjPAbvGaVtD9xhuRo/M
PtMzDXHnfuyM7PB33VceDPCEalSbxlWFaYfhludokFmPwNh8BMi7cIq3WZ2m
ymUEEYBeuHvMIiTDGwCGU1FvJaloDwpsAJOFPd1P6boVQJni9A4rYAO4Mgm1
jWj0N9ZvKkP4HaYQEQEyJKGKzfzU+c9CfKSk7y1y8VoOJJ/WG2DWr0P8+taG
RJ2Y6ygZ+SHIKFhZAWYBuhtTcd28nHQ65BwFMs19U0IlI83khCBmb85jHkd6
Q+eJQR5p0WCVs3g/jxQ5DVHlOt2mpmpnl70CJ1nRPWF0LOT/063XrisLYd30
09YjNQRQW+ZvyVpryvqH/0JaVzJDNIONuyyFQ4KWmqgZnGmrG3+ogtfvjjXJ
1QW1TZkJP9kSP7rZnwCwwDvgCwrLoy4kL3V5LfaXc5GUpXQ+/CcweXjnbTqL
CFAgGpr3vknOvA0gsIrhKhKYwC3uCHRgEkZVC6tsXAuJ5K1xc572mIgUB7OL
B/LNWVYe6s0SbO/aXm/eRUqYONj7W3NqfKypHiCnqmFle3ZOBuguE1KsTGSM
GVfg+5jvlXtI6wQy0O8faCSkepTzfkUJbm+ymd1uqiblBGs+UbWK7KZsoxOy
c12CAAZtoiI++T/fb/c2MM9HZvgjVZlOGFQohWkOVtsCL1xVDS9R3wtzuY74
R9PT2EyYhGfAQm1vPKS/d4QZA9nJhS5gZpzACEUiNJ9M8JE/d8S/j+lzLbwx
udfZEC8e3UwkyeO3Ua/u9a8GismX73pvGZ6nzJCrvpYzpnwysHzba1Py/I+3
74AQxMi9sZrxIWCcWJ9FGQ5MmbylImD6CAdSi/8TH4Zb2L36E13z4h9V5S44
lQYi/SyboD3/gch+JEypaAgT3ugX2dakZw++iNKgEuccq/DyS1qTChimxmpi
pfUEEfWiz6Hgk5s5zBRu7upwlco9RYaAO6hY4KVDRsDKayJhJnyQSBKjdSZP
jOIHTlmVwt+a64QInnFRhdySSneX9yRMmN1xfQSbRFLDf+XbRt4V/FngqF2V
aX+/hrNWfAgIoCTOY99Lga64B6I/qC/oXHDfl+UaQgxRgt2zTgH28741hbvG
oHyM1Rxd/ErnkRN8wlFdDBE0+OxrUwnqJZYQdIiqKULaIJHGK3DuTeVkcaRj
kvPbeiGfzTI51m3lDqC8rqxwNhESeasi1Rhl8PCbnQbK29NqeSRthTUT9UiR
MFBjHm3F2Fh+76eK+Ty1DL3ZZ4U9V46pYbXmaS2fTsHJ3T2LE2hL6wmBTJti
LDLx9HgasLEfTXHOOeP8xKlNOpEzqykyQ0Yamyw+dGPZGarHJz7FWSTHzroz
dkWpcqk4RtbZEUbwLyKa8aZKt3f4OIGXL3QggtPfzx1UUYBp5KTFRJ7q5fUY
ki/6+nTrQXEgGOxs7E16yHYbVIhBc5h3yM20H0E/e4HAlt/WKt60nFTPXvri
GZcyb4EKd+JX+rymIrACa6Wd5LdyNAM3YjOTgNsWa+OUayS2egZRvWkV2pl1
0HAUER9DDgdg/uDDNvs/IB03CDTtIPrhTjQvvOAHa4sTxdw0CZVBaJydgrd+
yYhKnEApGasT8rvb61suTgxuVvk0tEnVx1TiUah/9k9AtpNKRLlhOBXzK1kC
ljNvbU8Qt2os1vitEjvUMG24e9z7xElBv/yoObWYxfQ57AluimnPeNDOQ022
XE3Ut3pGhfPkLq2QfJ5z6MOgGfbndmPsx4mZRpIL31LEihE35xNUL8pMR8GC
B6tSPd7V6p8UsVnQXON0NuImUgXCmPDtuD4+1LPfUS8lZjucas+hObwAxFiT
OkuGlhaLNdm8N+p+C83nO4NxUHNzAaJnw77JyDHCF0bnFucKtfiCdzbWgTPq
bnkawM0lOxXvmrFJ4fCVNZAgb7e+/RcnkSL9jREe3kEsAaGHJWvW+R1Au+Jj
hmXvlkQxQivZIeAjsFUKtDPjEAm4Jgh9190DgoIT/PWMqCZWtaBGzm/LAvy4
er5VUb2r7OWwImfffAXc6V78MwKEr1zCpNiCI+wIInHHOFTpUgVj9VUZDace
zaJinQgdV8KmdqbmPCpm4pZmuzHTar5a+t8iPc6ryZ2Ky5fKEkX+oI3b7WDf
fk+0IbreZ56wOuw2DhUoZxjBCGZO0AgQ4cy7THJ6WRLzFR3PsfDlsoP5idnT
0I8oYZkXljx9t3GO6Ejmm4lJuteLJxsB7CqZufCgavypHCcEw9rXdnmDYXHs
zP+Cd8gQrIO5ukL0mda2jyU1jMilnp3w9YdUTO06C4df3hkRhk4jHB2rLwa5
KdzWQ/MjBV46nySvUih6HC02ysJG0m3+iRTk6vNWNTe2UoLF10Z03kX9cEgs
5ZfqqMp2d4PYE2QHVtyMlW8Zb8MfZiWKQOajA6I3s30XaJD6vqGikMlYJX3D
gM/kSBohiKox53eALnbIHSCR0fYvYe2buoUghxppXJ+EWlV3BS3lqNoQeoEV
qBR2iUxyOugyKQz8Uq5gWw1L0LSv1bz/FSFjsP9rR6aUH0P9mHtDqXH6vFzR
WNThi/03PV8uxj9EyfcvLrxzk3lUW21XgUWmPiiq3ZeE9Ka+ZgYbrf+Zawqh
QdeP2nKeWA1kJojGiw0khk5vaTGedNyBFWnh8Dkw3Hx1XzLe1vE5CqYv2H5j
UvHl8DhKv2AB+68kCl1rl+Rv8A+gFzD723/8WPz4wKWis5qrtykI6cIlAniQ
zoL9XLH4Pj65tF8XAB70hmM78Nb5oXzfVjrzwKgRV9OHAEUJHSfuV5OG5Dgl
v5X+C2e+TBjtpJrmVb7hKCEnCD6Q6NPMQgYaFK//9dA2IOjzT5ai+s/TlT/D
vk4K7M8UZn9YyFn6nfx+RctM/R8x/BhoOSwzEbTcoKFQbF+p67Pywft8qu/Z
8qkk0CgTzQwlKXEi4SdOzR6yMnIRqSUEmtQ4NmIypFRPVRyNLrAkPCO3nq61
uO8dCmwdQd+5vnNDHpOm6Z3j7JMGf1atAuAYPJJ5+xC3e+40nK3SmLxY5ldm
K9dGOwva1l48fOsVsUY2QtKO9uQi7f6FyOhahN0Y4NMXs2Z54R3SVU7jomtV
PLvyhW0JbIQ1StKG8CxAe2QcQzBEwUvBVKN29Z/t2UGFj452C43NOQ/7eNlS
KTCe40bUBLzABnKQOufVfKd0ZEGWGWy/k2oRwyzvYbnq3dnXI4MmeAAnqtMW
uvVvHBN13Ca89Q+pLQ+y4zULPAnCMDiMg0fwxdQKjgzU3fXldsXTRYFoCzoY
Z8byNLiToET4pms9/G8RNxEaRSIX1SRYB2kod/7LN5rGpVU9RwWLWtE5OXhq
KJDIQWQmW2fR2OfcYdosgm8x70rltj1OXI5usVsQ94eT7+wtTvka3xYzMUuG
NOj/fJdpswNvdImlhDA2B6utKbHTMFU8WzjMhZlGDApREPcuxVLEfUG9kH7S
KH6+K/FGJi0PweM+UnxShLpXAO0fUesoXtwJbckEAKMPoO5u+kA7Ur8ny3E8
h7mI+zC2+VN7EsiHZeAfEhUfOCmkrsBrgE+MD1u1tuEskZJglFx8Ap38p1V4
1Wb2XqGhN0LaaSp2eYrYtv9vR8zQmFISRalWxLrcVGafwzzkG+SBtkjwTWKR
xE/WEWUntzCjAj88msumED+skzIu2wtUtJevL6F7JUKT/qbZud8xQ/+SSa3c
o082pdQyjAKJvnu5oKVSkrruLA9nV639onGNhmSRXdZE7Y2sGqivKfdi4SzR
LFKhfUulCrLkG7JQDo43FJ0MCNo1cmJWjnkS9KYk6Pfc3/fvgAwWsYG6Oovo
iARHt57ahLMP3y8PLgrWsH2dIlajIaoQhzFP2XW1fAuFpoIt21tK/8kenadi
AMgP5c2GRD4Y79ZUZY1cwS6ll+EH9UR8idB/Oezvv4I8kta6fKREz6XPrKxJ
7LKRGV3fY+mM3Ft9f0U8m1dAqMI8AS1q3x1TwBQc5IJtdkdbjWyZcFcH11Xy
WBavWCK4oqo/Gps6Ei6n7kNok2OuRxKgR8ypMPpabdfvnr2R+VS7I92XPYLW
rN6XMEw/GdfMsGTy0sZWrkuChLTC5wS51YEn6vV9jq3mG1nbGQviUHUVu/wp
2jA2F3ZrbR2076dl1uexiCRDRaZBMBgDXe8vYfpRmh6VrSVbRCHZgZsnzh2c
MKQIecgd0zePRmhcYE18ZX4WxXe5i6YB91GoitYuGlga42lG8J0ng5Fu7BAz
+p3sEUrP0rQ6vdx/6gHJDWdQs3jsWIQ3jhhprANUiGXFLi43VoWpHNdPQK0z
vvLwBUf46sz988iO/SSWgjmy/aG+z9ZOZ6HBx0ZAfk8nW0Xfd3T0Ybvqbkoh
W712/NGyOVK/8HnptKc71B3ae8JqvIzSWuVUb0S/TQeVPoUnH5xoxkDUjW6J
jNfyX96PXY00ZAlvUs0+Ci/NMjn65xQEhQhmXb8es5HxMZykoiHAIRnh0eX+
UY/Vdp0F5RBlgDJ9HM/ulJqSJIhrxgOEMdxNxRAB5uYNO9MIrWTW7CyAb9uA
3d9ubephTdWoJ0HmuCXwFGQTvrYy7gxXqSNO4hAfH18kbwpaXc08AsurrWyG
ntbhIScOamYiV/ZGO4VjwasEkGxPWOOniZz5YfxHGBYdMGEnB9071HsZYXmZ
J53cHv4G+puXy4C1TER67k8+A9ND2sj9wU8SonD2PgCvG4rtKnuv+VrjYqfe
W4MOfrQZsRgyNfptviUitfX2pkU7nSrSjuQ1KY54Z0pqbYQhLsTi4kI5+md2
2f0w7mluvlk8zPK7I3iqJMhV1csfs6tB/s5W/+hkB0oRrSe578wq8v4/DTzG
IhMipLY5/OaZHGN/Y6aHuKBGs4HXa8cdjjuVCwtzLH3ETw0jRiPZ3DiJqIT/
5dXQ8IScw4lsC4mD/DeOA6MPgsP3f73DT7+UYRFU3g8/dKGeYg/n7yoBLxvM
HLud+dKOJVPlY+n7TVyv7+f45NRIn3abKF8xbNknfzZlWsFSg/r8lW4vQpO1
94IYhy3RM1xqGu2tAWYELDiu0Wwefe4Ka0JPfeGUdBfJWAyLSCa24O7+/phe
UA0OiA35xcoJGkRVkOLr/VJblwJwsEsslol9kAdheS0/VZQ/4MqCgywbexMR
CPg1KP3vEts/343G6yDwer5Q6bdmNo/HGvy/RczoDpY0/zP35LjnU9MFnx1q
ofLYAfgo8pZExSBFK0xJ+7Sa9gqI63QwgJE9QyT8KeTjNCE2ZZMMRVRGNJSG
3FZyh6DYdaV1qtNnrdktfedEWkFPwE0AVNZRdEwB750dCRTPMsBY4ZAMA4N8
lR7eU8rmnbdB73wE7QDOFO0ur5kJxTfh0XFHZ+J1wkLyg4HpkTgLhmS4KxhV
zso2oCoo3xMxXahtDRKw6pUbDG+cZXBtbuBxGUbUs5c0B2QR0NoI9kIIWda2
jCEmX7FNxm7KivpP5Ps0UcxZvaY7UjateQd2t1TaaFKAJtql+LYDqxQTIRAx
Mgl1sy+PjJDjpDRJRXXeZGZNpoqnjpPY1Cq10Vfgm6tBEXkRhk0sWyHbH6or
0Lsczp/zIlhcFPexK58uNiStT0gaFv3uuQGxUdhF0jaJ+80OQMulgS1kcPAZ
m2v/0BaexG5KgTQR4tqTWkYiB3G7cteNiNyugBsdsZbjzFR7Z1iN6ELeVeJ8
g039v5ZjojEyJ6R6R0oqCx7hkjBzDQUZPmcMQOoFLnqgT3UzJPo8QoY1unZQ
QtNtBMgWVMowcxBmRQyzhp0ZhvmgZ4fJS/Yja0Qw/FUdxeWMKbhCAayQBlCN
8WeDIhQgQHqOedaoTsvApP7hU+gbxx2X5XZ1lGhLwJvcLURGSmLCDHnYh29c
dlNbxXo5MeNqgxy1OJKRBxok6lDjntLShug/Td3FHR/8NfRMXP2DuQjuvWXV
kmExQTVCrg9IjjTKm+z8chPjBE2+8AzvD5oH62dmgw5qjZVufKLi8rPhpYQC
EVjQ6F13L8bl6r4l+dryvDyWnM3kVJsNIAq9nlipDVYJF+Ht1Yf5/bc68DX+
bs0VQtecbPk5xl/iKu4OLJes7t1c9NKVOOa1JGsTKoEV7n0DM4bhpor/L//z
/Nu+B3kBotzjoP2oYKhFd4rv8stBVjcScFwoeIFlVqml5CTlW9EPyhcZj46f
9Sk0H+iYR5b/bmkRf8uDvJ+J7ceLVpikPrfC/Bs3vQeqTKLgFAHLQv1TEeDJ
KuI6DHw39fOIOIiCLGiLTP0O5ZtQdiVwvEjD24n+j2RCN6b36DEz69hfTkNN
Sa1b1uTeolxkS68SXe7fT6bUvP//G281GFjcXypVQQim0VJXUyEtgd2Ot38z
5jTc2p/YuvwZGVerqVPo269HcNvbiLKVkV4JfD+YiPz84HrJFtgehkWb9eOf
f4EAE2v/gSZVBjsL9K4VGewHFqc+BMocI/4Wlq5NF4qd9k7HKhWUGVDUgMxl
pLaUsOyxjxmnkBrW+Wd5MaO1u2Ltdkk9rR4e0oFeOO/qL89/4UbUI/refVJZ
c8FQF4zIZla2OxNAWh0qmPyUzN14OlhbrkzdL58X8PYE1LheCFbbuzD7oS9k
pl4BWSq5MWTRX3d2iZBmSoY04+Auf5ILLKU1pWXlnA3L92vZUpYM8XHtSimT
ibzvu4/1+PfvoJbI3cKsDB7isiaTgsOyqJUNnwNLlCqWOClAYqpvdtrJXLMS
MmU9YONIL0qd3AjfEBNa4xSDj9wAWuDNmJD71TGjewMqmw7JJak4y0Q5GY1R
vhCJqtjWHbn+09+jKpBRhKts/A8b80rJr3FkQ6YkCCm1NZngRXzqEyYiXVIG
sqC/VVq6cEvRq7u7x/nnDclOjOJ4eVZ38cjyGlAKJwiGTWw54VZeNY2H7h1p
682E6wF0zGaz6WdgHAC/bXyiV0AK9EtatmNxEjWRGaaAX4YAfJ0yGgJP8Aaj
CAK7ttE1XUF7+W2tTyxr8gAd1TuG2BT6EXngTF0E0Ijahr3VaIpthMY4bqpY
ognGG4GmxHzH//99eV3+T11aEhRu9eEBR76UdtWkNWhTF6ISP4J5Eh6l2qL0
LlfO9vhEG52h0QPkdP3MjLcFx0eBQAiEhxUAb+EBr0dUZomcwfino6gCZJwt
uCc7yqMkJY4wXVCjyphP0cnEThuCMc6hPckxy7h/zTWYUb5LANUuVUDpqfq+
CiB9gB8B2mFzWJez1a2klX5LcWNHMuerpytgpe29yDqMU5fh/hkQDQyOnITN
F9hCrOcmsI+nLN4tC47wrXu0VsglDvg4f8ZuoFHusnngcwV8YipA0NyMwjnm
W7j98stqLsj96XVUFmHu6PJxC439RtwDtQh57WkxOI+pr/ydHNlPUyUL+3OU
Mw5rtWRu96ztuBJhWrFwVLGsxbuTk4R5TeTmPrpPPdnXjdQHbOGTbSSgVGJ8
iFNQYklQnJFH/sabx6wcXO9YqI5bvDqZgu7st31GUM/8cLj6gMWbAlqxHDTF
LW6wq7d1HuRL2tsUMKnpNqqHq388YnoDuAoMe3ND5DK/sdlyDvS5aF8I8P2b
FnGCtMojc9UzkbGS6BTzHClvpT6b9U5N05Dd4ki6wvSEt6OR5ITdL/5pW+Ik
D1WeBmpxgrVP7Fv1GHVKAhZcQumGIYChetaZ+0KUmRpoiK9+lopuY3tzWs7z
RJ0q4yjchbpRQV3m+MlCeAD1TYyxh1dfbX3J/9KiaqqZNaqnQuVjV4BRVbA8
rJy4L7k5kNDBmJ88n0Y2xdTmkXg1J0K6QIIFf9D5L3aniNiKaduPemOPyNZL
1j0rzQ5QHUyfOeCDmxHh2rBmPvIEWdG9D4Q0VKSKFbN4C7WvSv0w9eIPV/ih
fLfcUVOxVyHk6K5R4RVfINnMx63FuBR5caSd2FFK01IP8SdL5XzIObwA2xKj
+TFOQPXXSYEJI3Bhd3NPGcE1+bSBzNATKwPM2PpQdAJZI2YbuMSlykYLS/1Q
5W4T0eMgHnqH/aBZHy5/9HOQ5c+lCJn+yok9s/d90/KIVjgL4rYHxBMZzT8W
JQooIx3MTr8wN8a5t2oJUHyHv9v/OHJqoPFaKJ7gy9UOihoHj1hDKPW7084G
t1P/omkDVKl5QOiknrz4twASRULWRWXvdLYMKNxXRIiPjzZhAJkshVpdyW4x
GnUgbnIpCcIvVUl10VLmou2YdYMi6s+l4MdhIdGm1KBgFIjHixhSN8KRpmc+
prxvXu3ZnoSEDneqdSZNUGLX1un9vrDOYBag5As9dP1q3cmzW3BANgAOlfJQ
MFU2OfVcmVYHV8jAbdA1HJRngKDc3MrIndzvqmLCnuibVyBVYk4sl8jMW/hO
nTYPJ1ptbN0h//kV+up/vz64gp3meynvkDzd60qjwTyTKQhXCiTQXDyYR6Wm
5qt/tjf1rtpFmjb/voVW1bvp0eAqsjUZ9PxXMscfhMdQMp7NA5XWq1KipRXL
2BygnGVOqsHUSavZuvT6WhzvGhhYMHNeanIufHgwsq6sulv4e6DDIhLQvsAC
ChXeBSOnJZVaYzOM1fs9RtqBprFhjFUQ6BbSr/QK6XzHtNxU+lPODVnMDGuF
2CE2E/kvF8oZqcSCwpZEai1CgExCX+9eAkhJv26Eo1D7N1CxWeUAb2PtfRYk
2FPEA8LsswZXKOKHqblS7z7JTmH1Z4kPMJ54qj6ixqVFR51KbOylXBB5yeZX
rb7YcWmYYVTVOLEbQkIdJhv6dzu8dOyHGvp9FkN4CSFPij9bRAsz04dltDqD
Dy0usq4JRUxGLgmSbrWMUzZiHDZnqse9MKbSRRHajaW3mVuvcN/ai6aHgc+E
L5679NgffXjsP5OGfb74nn8USw2nT8+hFP/WvNbpaKjCwDRB7yqV4mF7FO3I
E5KRLo2w8Xvn3QniMFOUkzaUn1fdJ3k0vJab5GSMzQHxU4od+yWXxpV+lD8b
8oCQu4IgzvJc0enA7j9Gm4/ulWtPUPV7ShtHbmY2z+UnDmCz5MK1MYbucixy
oiIvvQDiyasfpuZX7RuDg3R25rXcn3IPwqapVOO5oPTXUPdq0wen4cuOdmqT
3HpxsjeuLy1CHHh4L1XHpMktvmnSMThoUJI0w+f7WyIbksm2Q7ZQWOOYv8ZH
1zwaLsqy92lpBkiF58T14y0hYaMEhpMm03X1OzLQgAloBusB5Wn8qPMubgKP
9OcIfWAxSqotGT99EGSiAknXjnQ58gmmIph2ewDIBTMRSJIIJBfOC9j9+Y95
75Le6T7SUHu5BGIhuVQlLPwRL8VF9Qok4v15UAW04AftNsyIJgsYS+lBzPbw
hsakWq3RzcOiocpFmk6DZrtdUHwlNuHnyZ82Y7kA+U5jecqLWgVFdtIAchQe
5xuEl4jfhCv7zJWN9QovloEM+8H5lwo4ykv0eK0RIAjTiU//ae3uXqRQlFrZ
/2moz6qTGZHyPsMx2xyUZawwKxdA/pBqP5xVvMIdgrwQSUgkUXOYtL+GPIAh
6dEui7O/1YNgeFiZT6EAFv9saxTGAL5unnB0u3te0KUSYr3dNVVAicseajBB
vVvyorwsqoEOq2De6r053Csvn25WN0fNH7chIDBjRz6p1g8KBGUOFWMG7eV0
RL2Rtnf7AFRL+98eTsr6LXJn0fwT12d0WIQOxb36a7nfmkwT9lf1EpfXOvUq
LVuch5CNE+zMBu5v+BVE/UyOeSUxlpOQyWXm4dKLCirVlayFTLCdHR7pPqgA
n5OFDluPkfsza9aypGjmsqY7hlF6D+Hs9OButCk33fW3NOWct+3Jp34wxVUI
EZNblhyMgSsLVyVDaGvMu6vNpHh+v98bUj92UybCWr0a/CV+WXiB2HT+MQaA
hlnvm2skZFDjccGKs4l+3deEyzMF5GUiZWFTqZwG1YgjGPOSixTwUXx8zge3
1A1jgK5525QV3j7J8xX9PX1UVnapUJFd0j4cOoMw9WivXUUObx8nApDKfDMV
a/HHfSGKoN7Zz0R6EftTytbkLl8+Udn73RR45OfGteqhYi+mXKYKVVIgqc41
hs84jYPxJs6YZd/5kQPpzc86aoL8mUGXEolY8sLm0Nn/s4BrkLkB9zJG/8/L
zI08KqNF9qL3QUMrp6YzZmdbFDIsEkYeF+cLyxTNbi0aCNvchjwDVF2OeaYL
bDr8WsJgU2yQgasXBqcWTPN+6XK64XMKceSF6hL0c4oV/H3mNEcEq58FVk9J
fL4/VHUfTsNRHU9t3oltoIuwUV90eypcyBk29svW/DfMAFp1OBeAqKihqI+E
/tX4ddqjGwP1t7ID0jaQZ1i77yo4yYScbu67TS7AjJ1v36W312jxzPXhYsKy
m7RzYa/6MASIIG+1kWSd6VUUu3szR853rbWg0rDpAW4vA2GD6rOq39RdK7zX
Qp4EtrfcojPcEBzfmzN90sKRb+xSuh6AHsOk+8P1bHzwkgu+2NeLcKeWYW6t
so7AQtnWUATc3xwwdupkYS2LIWORf/8ruoze9mYcO5p2Q7p+nNFCynAeaFhx
czxjeLTxLKbW0qIapnfonQg2w8ekBhHJw7s5g1C8wWjATXZBHZFatL6lsqpB
dxHLbP1lv5LE7RWfjeRX5Azl59SEJW8GP2+UAJ5bZUb0I1j9kA6gjbj56m3b
wZ0wX8Kc9rhXJEgsSfYTrqEgu7MvQViu+H6CtxiIwRsowfuI1mtSNR2fJ8kG
cIYmlS0k7ZD75wpIXW226EOWJmW8rX+r18hG0S6flGuJnbe5BwWzWeZ69pOD
6kW2SbcltUz5A1kskIb+Exz7uj67Hc0JOhifnDXSr19TlglhEBbgfYKKFpF/
J3/dcpt371KoQjMF6eu7NQ16y3TXf1PK5snrvMP22S2eSqwpdMck1o/YqRYN
lNPfBdqsvaVgSSjh5MwuaD3M7pp8plasO3Av6pThUCX2Mz60vJz1o1+xOM9f
vfk7SKQTemPPvWLSv7A/gXmRN4tKO/quAF9cW7sg5zxj884/LM114BfH0O+N
JcEc7qvoDuqpPoahjnnpYr/FCTuhllcFKrTKoCfmidlPAgRNe7nuJdVk5r6V
hEWNhrjnI5rDWfwmke2sWydnU7kaox+zWKqn7RDP/YSVBNV3SiaTmkivAlm6
pRpFFSe3qdNYfHiCSXMeKPW1biRm0G6GxJ0QoQE6hTljMi86ORLQYirsGew2
/ilXkWn0P1ut0HH46jucCGuQKRdfMURqn6WDnjAUUf5FcnLjRB6Ufj+PDdhM
YWvrZ0YwFZz/c89+uL2EMbOyB1QE8/yaLfPKvVIbqAptarD47DVhzAHJI09a
NacyKUm8xTRWespX85EXbw13Obx4eoSGogprWt6CQhRG6UyAJVYWYdWR/MtR
OHsFg/Z4A8Qz2eOOD/p2Kq2ffi6988oDFTvMO8MhKBT2NYUazv4TAcbUaC+T
2Hb4tNsCdLk1A3RswmK3UERHNRP8UAxma2zBtsUE9+I9VKeAevTwbr0Ez0+I
iQjMXZpRXaNOR9PDSD+TZ0CmB0rd2SQJFuiHry8eHJHuHe6w/yF92610SeDR
hpO1wPPHyl0GWKQVSgKYkPEZeYyBeUPaUQ+PJmQsLHxQutUnoVwfmED65cFn
vybQxNBAIrTsRISwluqKmOT/g9Gp1Vp8eHzXIFF4uLrqUeIuZWOM/Cwn+Xm6
pmJYyo8lg6gC6pukw9WeCTXoXLSOHJ3eWB+Z9m/mJg/lVWPmfIDRZ/dFLRaj
hRaPw+bAac89y9hMvjIZdV0wx5dSi2iAlJVoXFowQo4U8aCF3no0OoydRIZe
OPNZ/uVEVLup4ogstj53+RgETNCGJnB4JGLQ64TqV7Imvb2Trl/MfZRXRpuy
CaCaeFJTgHxAoCbmoLWGn+Esmo4BqrmyHbJakeazYWqhauBLf/VG2bx4UyxA
Fh85aYD0j03v1dhF9ea3msDFaN0pLd+X8Qn9l28QjEu0t0oSj75tGGT30vfX
zCGT0ufnuEsUSEQiyjrY2JKelXJ0QV0TVtfT/qmZQ8Dv8tQckJjjgrAgo7yH
iU9CfAkTUbraILrSxNORkdzBkBYsp6AX//txW/HHJmAcsGr2gZF3LQuHXzIz
jnmrUDCMSoL9iEdYQFRU7qslVEcPMJFTmuehYuJY90RC9VTN/bX9ZoIIIOE6
VUh+NsFZkeCARQbxNFTA5sqUpNm0rBvgLsQBPtY5PjDJ25/6K0j+Gd+m+w/y
OyaLprBrMAM1ZOO4D2HG1BOPGZJ5HUbAx5e3u3haztiRWiTlw6yUM9/oSg7k
BYbnU0v+i+sG1R2eDhCQlWkJOLYUMuhZjgyQ1KjlAGcb+G6lpYMDyiG0GaAB
s1Je3h8A7a8Io5m0ts9tuqyml8VchW/OdSh5PhUW8mUbiuW5HJ2ApZYnxB3X
fX4NDandvxQldJbe812YoM1l69YEyFgG9nix7xMGtzqqmoxjYcW0vOJI6S+I
Ofi5EqT+RUxhW9E8tiPlfyuP78F2A/bkPPDihY2yR41MQt/2H+9gtgcq8K0w
/FVebdSh6P1a5uQFBQdGyMZV0UZVLkwqh312kdkgNupT5XE6xFlmGXfWGvDw
3oB1Pn1gcCVFh7jpRyLZn4yRfiXD9EA6UFC4KAj6c/dsbPt0GFkT9ED0GME7
l2U05+sjXO9AvPKU2UkUOh9brfqfhXQJVt4lE/icFyGpVNea45h/VE5c1Izd
JAwi+QwDk/2HvD19q57RpVF80C+WtcLCrNde2kbF78JELygwhGCTvNSBZRHx
qAVA+ugZxqJcM/NREKEjOPaYDJcIaw8M7IxP0pQMaZqupunkGCCUysIyH3gl
DVWVPpRNrmivIow5ZbCWS5wde7bfHS13xC/1zXgwJAOaNtAcl5Xn50rUPeie
n4b703BIQ5hTRhRuqldJhsugOlCXM5VKfTz2EGv/my4JmEffSi9KItJO9OYj
sQJ8O8b+T4POzUsgtI4lW0y6zgRXXvhnJfcPguY/i6qdMnouPGPN5De7RFm/
PsfB0AiD05Sd8vxrukzNuL5Y44fc/AKR4L5PNAGe7KZdcXuNO35SZKq34AkM
VFa0RihBMUyCdzWmqOHwr4VcnjZMTylWoKMn2xlWaMltaissimJCXrYbE5XZ
DTVL0jkXP6EmW8Lzp37mPCKZsssq6CAunlNXq/r50FlJOpzkc62TyljXpXPZ
rXIFmeLC+uZFkSxXvaqyWNLjdajXH699jPHPwIbRMtzeqlJ4kskl15F/l4cD
9oBmrqjYqLntmC8EbDx4S8xhPo6scO4LpmehY5d5K/OWGybcUz4OLK/aqO59
rry6tEFeIA5Tp/0ZbAGi5H/MV+Z36r7QHdSYsj1+WGjEQPn1r7Cj5EhFFPfo
38hbgLH2i1KZCdNKSTuFwXcNdrvBYd8DXME4bcc1TXdB/hlX77VAyj53c3uB
Rr1BU4BGtIV1D8D8/D1/vTfyjPf/2tLlo1wIKxk1SnOhtPVVNbpf/byNqooQ
ImPZWC2me5d5t+3xtKiEunHqsf7FhVISKSKh7PzH7vL+6MTu+O4UZtZotmv0
RkqS+hSPvKkImwL32g7UBhioqldXLhMu8Rrw4WGz4PU44TjDJzhk4YKpPie3
L03ZJDfrumYH9mTSjsXk08StbupsgBGNvORaz73HYmx9HoDaj415kfdT8zVI
KV3THifZ2X+kGwKspsdc+C6HLfaFU+SV2PWJ+jaQe4Xo+SMmJkLpU8wbEJqz
KnW3jVasvDODHrJct6/A17UUbQy4KqEBqrpAhYK2zTa42lIaN9WR2zSdCcII
YXO3f2r7FfWxNdHP4agsSe8OJaqACMnAxRM8wzmwaM9DuO+LD+0xAMFFb23R
1hy26BgizTc6tX2gRJ6R+suHLwiW11/g4hLeaU563jaHKSKGC0zf9KB9ptsS
tvYfvE85Qj7NtJg9erDQTtQAQuz+pSDqRqzRNYT5ARqtZZ/jzzAH5XPy9u/j
yS7cwOVQxD+t4uUHKnGupbnWuzynANRMtBWzWwtXHVrh4bjrilPhh8W+zvI7
1Mg57ZHMAWerFfFeU19JTvHR9W90xJtrOgg18rE8sRHpExyMTV96V0HGqnvT
Lno/4gLQ9FUUnYlzdKxHHDLHTM5J/Pcgy+rHqnSW6uMZZz7Ez8XWO5KhFjp0
KvUOHljnQWu/A05fNAMiVs3yorShm47pFTwRMeCnIxxHdY2Xww0MjRkNNCox
gryLNzYC2BFmB3fisgeoixRw9HtLiBf89LokfQsimsphtE/nxy+OU109Fn0V
QCOHxx1bOzOurLyej0DnPay9RfJ5vEQ6BMkxrcU1U6wKmAtv2MqfxVpMT/4j
xD1aK4a5OXxaIrYe2e/RcA1ltINJwr7vDD0Ri2WD3srLUU73e0/IkEuZA/sv
a60U2UwmYV3HB3XnhIt8B59VFCUoWtXpDEvCquHGlH/oFI5uD/5H5T8bGHi3
7MBZVlIyJoqBRsjITO3YeQ64AybP+5sjweSmDgN9xHngG3as3N5JKMztQ7fP
yLJZiia62LX5YuRkcMEd4ivAPXT9qfpZUUwIx8JNImQxiyyiUpwlAVUzpKg7
Wtbi5GOukCogXWmAXJXAVIugSeoE2a7K4zU7QrPlbP7/trGCtaWx4EVB6t1e
H4+VI+iiFv9ksRpJv1qquWBx2vx/ByGw4LiqsrUJqPxb/wkwNNC5Yr1SYtcV
PwM+FPI8HIm1Tr1+BaV45vEg+qbRi5dV/kXqbcQnrUCdMo/PSUVWEBR4ea5T
scXGkWY20mGrcv12ZA8TIQwbS9MCFBh+BUeywLdd+lGjUL32Yy2QVrLJ1Kar
35CNN7FWpLQTf7fGlkoHNpHC5YwIWuYztr+qnbQ5E5BJy5Dr3F5HWa7mimBk
ndrUbyQftLypB4/0T/B7OHZheHdoxRY/ziAyTY4ShKscqehRr0PFcnqlr5Sa
Ia3e6PrHthIlOUC9CQTopxnLhTVj2Jw5W4mDiP7JnUtx1ZcyQZXEsVbShVDF
kf+t8fzmC9v01DcH1NHfyMvNBsAr8fUfn7zEz+DvjaS36vH2U36j/nET4TC8
7Rhl7yLWvNqNHYrFH+78Kle7Hi3nGRxA6tFJqVLcPunpfeNy4ezE9+2nIfz2
hdBvBNi6dMalwjilZHS7aGIIVm/rJjRtvszk25ajrn9R7JG5DrfvfxYNbLB2
KWsD55ovpOiCRITZwBHwN99EntVNouyvBzC7hjPirNEnBQU9ej/KJDBF3Qaf
VSN4kc4GWuAnZI1oSt+rZnkkDVxCEFS+Dt8y9cUFvD3U3vWM+t3gnX05trYb
c+2EPXq8LeDC9JQfxw3XP7eC9LQwygDN19J3Lf5qLUaH5amuTzc9O6TqGTNW
ngewVvRQK9+7kXJvkNC8DIeWHxEbe1/jyHMExkY0ACcbf1wblKr+uru1AdB1
ZMKHmCGU3J/Ra4oQGy9y0ifHnItEAW+NjG7hq4QiqwzJ1s2190LVrWkvurbi
w/epZS7FnZt7bsPd9L6k7M9Z5ZANIT3DbkVM3W1D+xfxeoY3N1Q2O3Cau9P0
M0UMljWuvK/I0ZISy+NmXg5MQ296lt1xSR/UDApDU/jktR5yCR5sPUP9QRWC
nL3tFebAXDqNSJF7nHfUBJWv4plD3XYBnDEkX4erHuFYnyEXZ9Fjy043O93x
1cR6/xZWeug669OxNvfVfGHOarlXeyh81ryqkSY6CI/YeJdfqFW3VW/3VWhN
UFjVE3BY20EM6M2EWz1iMw7I25fP1NHmHvs0pdyASR5A2mmGUmC8T9F7xFfr
sH54mW5o58RGxXnTZPqfjtj5BhCe8vaPjwclCD6mjuLimi/jtILm7Q+H+ZkB
8rsSohy6QLQIjpX70wCb6Yq3u6sJnfZ6y+hen1bhHq81LA0v2ciWex3YxmFp
pMTSZIw4+hvLmmxJuG+XeBJS+9tbNIFv9b6B+au+1mQvgYVwdfbdzqapDW4h
70V8A2Iz2XY04Wvv5qVrKTS5yhv9R7LTZLWB6EfS5TbO5oUmck0fPPlC+GRs
u70GDBWdYpQpCi35WP1VBA3hyG1SymRw9MsYWMzBx0kD+16pzzG5KRidpbCl
TLTOx81edJlkeoyOjOI22HNhbZuioQ7jXV9+oVChtCQeF7oUuDnJPtXbiR7D
S8Wy78z/tsyfMXqkiF9m4ciOI2PgKg8DDrlvhvItYrr7VK0PjvK5ptGhFB1A
MdKGGMy2/mtL+6bt0l+n7cXpPs3YGLOYkj/u+OaXShEXw5ZD/CR3Tb3Iv79u
AopQ2amXfhq4vYqIvabV967zEEKkS8Sc8lbpXwnykKj2kPgFj7wh/EUrhFkH
cCr5RaEXBH3Tw+j7yRg5jd/3WjpsBrxgftKZeuVRXi+ikoYnoO3p6H7ggtrx
NBW045+vr0rhbBqaRrzy4GEAUwbJF0Wi+4Ao8e53eslU1izfRYZeuq7aso//
2QuC6zqOe3HwHZ/GB8r6yhShFDII7aI0hP5JyuZPYZ5G0PymNm6Byt1XYzHI
xqk2Rc/Y8fgs+Jkh0WzJi9eA9sd88T9b42BI/UOHMQuDcamvY+8qLjrr+4nK
hPRb1xoRXn/nlilxMNZR4+/9o7hdLnBf1Wrji/k5+E6eZ4seiWhgrYddgIxh
bb/ylZOmts+XPZqbGTbPPHx4X9hOjYcnxRK8L00DlcBR4kJx03Kvzypw1TWm
173DujW1mXl3RuHc21jG64CiOprK9VRHIAcbfBRsUPRGFA6/ZJMhrQjsnqKD
UPfZmA78byHAhICiqxJee6EFhFTwt0naLuulwvK6C8ETrY52xzu309p0nwkl
u+F6DwVDfAwznkuqTI7ub8j3VrXxbYB74ESUq0B2KtSC3fQz/uTYQkOvHZhg
43ZySkHc0i4iTFtDHZrrv5rSRQ+wZRPw4SY3oDzfhMybDYB8QqqRCvLuq1Ba
ILR2BFK9OuSP1oKEH9yaghf1pnINj5nR38tVxh9VlXxbDCklQsu/mX9JnwJM
PDKmECkihjvGtsHBL9sb6nHsCp2/B5VRPw0Iuqo3l0UqqBasA9L6U58+pKYp
XC4XANkHB42MOWirJeSzgEOe8gB/OP9p6KnzwPUoWdLjtyXbpjN+1fFAEJQH
xXD/C0iHP146nTY9LrJ5jUKR5V0plPMo8jfyf7EcsPH7e5oWeB53in1vwXHc
B3bXnj3FIOCApt7IVAfRQ5BJklpfUqcc2mORe97PnoCDCKDz2JUIhcqHoJP4
KT1uqFLvlQgk9OJvvtA3Kbds2cFohecimyrL90xn+1pP/uALa0F6hiJOdQSV
xZRzw46hshMC7iPhclkVqIAvjBp/BK3GJvm63DdM2VKVZFcyaq65gRTBCSnb
NCEgGd20pt4mraFSEfzT7Mrlz9dhojchnZ5s1+eABfKuy30sKxsEhmVhIpyg
79CpDI6NG2oEMAKh5iOPfi49Z9km/AOs64lQRR6vDd1GJbSHi2nvUClbshb/
EeYqnKt4RxXXx3tKu+bjJIyEcnhaHDkeWe1PDyayTqxORynYsMeVN9nCSHut
yCDxLvhG7skrLrY81tHckqjWzWemangxNEiO9TfOXDRA005/xINDPaOlS51G
ff+73yLDkfJUQNju5EwfX7R2A6WcWISZ4cn4WVwsKvf7tDq9ubEJibLi4Vt4
KWMr6ELst2mhBob/uwyt3U6EKYQ4ocL+2fdQaDJooPbeqlDxodSG5AmMQCea
N5vL2KPuMI95rYGPFN8CorVgJ1DztrYsKNbutvTqsg1NidH6+3vNl9JeaXKN
h7jULIRQJtJZXHKOTrX+pl+puPc9+OcHn8BwXsj/OpNB+11SU1oiQt4rbjsD
9fMlIXwLaa0s2K61+Vfr8QnmTfCEtdu51DoFYTIVFRKLwN0SgzioaNkBAF0F
rZl5nb1phlNTvqqIApHUymKZ/KuKJMgWuw5TfwkGi/okl0sKnH0VgXVW6PkF
8mFKfbAmD4hZ28lNpm1hRMcMdIU9+NK6GjXPStO9OGGkTiyNj+dacWJejYAO
0xokcrOMin1W7eZLIPYKkH8qdgwRAlLpPDyNVkhbYOSh5+r4zPazcUoY98vP
c4L56d/TPtZN8BI83SxJjkrTNX+eT8WHX1BLSZFfYQe88oHZLqUOdmGnswdS
IamgVm+yYjFjH4l3cvX7/fW3Vz8DXU+PWWNPJxERN95qs724KuRQAGDaVFR1
0ENS0Q9pykDcmbRccxB8U8KvIH4nZoWbWz0MN7T0jQPl7rI2ZCzZlmkOe+sz
INcpZNjS1o8D4nZpAR2zL27+JZvkZCzaE0JL5FueqTu4WOYRFBZTgOwtURO2
jAUWKQ4QtmpW/4I9n730RPurJu2AqHzqalofBHYpbe1OG/0r21aYTtD/XObk
3Verrs7UdDfvnRZuUOZUXjlokNzsgpOZq3iyV45IQGAURLDHZpZ8A9fMz6W+
m7HShXOU+vXrFVfg5tD8JIkcDWGfo2xnKRNPIyC8u9IP8KaAvqzjnwN5+vAG
R7dfUKxMiOGSzquhiuVo9TnNORng8Cn+O4mpC7jaa/iegNlVS0YKGUbJaaod
hY1pzUye71/+HVpHKKW8ijfe6694jikeZbit+R4IhUx8lNF1NAe9pnU14Vo1
9PuHqDjmD+bjoc+TOcNQa/tWcr4U5JaR0oVGgkRnDUS3whNo0SFcqdtczbDs
uUglsOLXJD2Ey4A8AHayyKYwCasNhmfP7JoONQM/sTUijUKYw5QR4Gwcvnfo
h63hi2Ol+80z0nYtOMKl2RKsgyVZC12a+QRWnVRgoAhk1xAtJ8S0wbBRb1gS
1XQj5XEcEuQVP6OrkSYRhp90McgWyLHvGNBut8/jEQ3L9CjNh3LolsUzMYW8
MqIvCT6khcMwMMgvKkISfVex4AOqTmCiphJEGWPyCWMLORNPjqwX7uMhxPEp
WFTAbHNTQ6zL2tUCzvHz8p4ZJktUT/3jKcvPvdMR2d40YGTh4//2mP6D52G0
WQas320yRY2jpRYlpvVIpZtjDlds86K/sm02J6lPrWVzFAlxKpsvVe/Ocl+x
G50N/E8i+QhBgRnotxCkpAEI5K8dwBKBnYRcLqjBmaZR/w/SUtm/CLlMGQ/l
7CXkesrvT5nyRHhDbeRn0cNZ/dx8VEny3J/3o7iu9P2SNc8TJI/dCgH1YVMX
qglcECZIVLxHddzmC3yk16WKXN4ok98GzY1n7jb8JLJIxgcE6KRnqKwJMroM
YxIFZhVKdWEEV81NCGuhrfdceOJd68N6HC2zGWgxWXVBxgFC44D5ZYl1aqml
6q9YbIKySUy86cxtCtd3rLGOqKn0S16hEkjJrLg0nesLZZmxaWsO2ejj+xjN
r8mA/KmkhqMP27f4kdS9JHoZoEXfYwHhkL3v6ysJsu3mk/lBplNgytasKL75
Zb6URwL/2/3amc+qts24lOv171w34+Y0nKXA2ryGR4txQ8TNMhG0bpKceeP8
JqzCfVpu9aDBPe1jZqu3WFPbiTJKHiI46Lew0sCYfRFuAQ4ejJ8TuMsiTDw2
5GZDJv4VvUCW74yYQY6om4cp/l+LE4NhsMZtq0vKVqOsqe/IT05c2BJAsk5x
Q+JsGbUNggTORrJgn4MHNZlA/3TnXhLvfzUhiZFx8qPTPeR9Crw43RB/QSIV
g5wkCYGT0oFkvg2l/YqXQ3Vps7XTkmuxWhDKrpKlN/dMM7ruR1NxRVePUrNa
IEZy1DWIai3SwlyNpWg9QDA6zGCdOkUjR49991ZGF31jdg72UXjPZteWXYAX
VPEkiv7YtMvEQd5fNHsZdPN8lXvy8wd4iuCt1i1izLP0SeQ0TDPjMofmOog7
qOthL7DWtV5j+wgs/BUPIoXPnWglGGh1QuNxv/LgcHfcLAFrim1hBJk/0aMQ
rzpmjcFZUEvS7vTzDzFGv/1lhM3yyxIl9gH/0nmNWEkoCO3Qk/olTnP1nRao
k3zVPrFTWFjrcE7WB2dfL2LUgkKwdRFD9Umw/MpqYP31eq6vdPZGhfmkei15
m9b4ssLDMizXu+S/5pD6e79Skab2r6I2LunpIsxa2pHc5w20tICwfdESOWrE
qMyxij3yu5TNSoE/BaMyqirPmiL2F9tLDBrzZkrfkQg7XkMezRwM4kP0EAou
J1RDH9vDLUke6RgyOnvPX75ceTqr3liNv0gUfTXwvLPa0q0IT2f/eX5wppOn
WQzUzMFtIxzjFwqM4SgznR1cGGHc7FsaciV/J7LzdFV33qLJ+1GlpGLewOlr
CbIUfRhXu41irR93cJ/5bep8AbvM9ZHIDINMl875+MfVPHl79eMyuOyS1VD7
+hvflVQ+mvk0L6XMrlB2J1pJbD8HiMGlXrjNehpT6aROIGZw+IbsRfCpTF8D
0W2g0a9zXMOIRYCn+yegBk6i/MiHCYmkCj7HklqFTXYY/a5ghARVIghxW1Uh
Uxto4gfaBdhIK+pLHK455ZOTGjOF5EDmnHTJINMC/CN8DkeBKra1yxpvNDWh
v4Z2IdgTkf/3tdCDo3PnnyqdFOnEX8ZRt4Sdyl3Zi2E6tLZ56qgrzu288Gcb
sSoPjgcMq/X/Z552N//5qyQuuBkmcDOI+xQBtoQYkEyETiWDUy3S/6kPkNJc
dg7Ux9bMQpC0HsApQKGbVWFDJItW0LKwzJS2nGQ0ePnic+zElkRsTHbDtaa9
OSIt92MpiERjasrX88sJocTiJfri3muEf9FDnzU9RPfMYjcLx3O6DV9A814e
pAMavXEoXPqwTLNqvHDcF8EnhTuZKQHr5fN3VnSb1eWdYmJ73j8IP2OSRfmv
ivKC/feR/xJzFqF37Yl9KuWHU5kGsXUKnKlBs+i4kb8b1ggmYR7lWxcJSbrt
NSxxfi80p7hUiKWAdqReuuD0YQwnwGHiPDEI9h/EQkiZt8b6mbmooldWYs2H
7sQ7xpBmOjU0g3l3s8J39CPbIYlp44j6pPK/5pQ12vtTv0vWWH5ygOtTnAaw
/DanCEd5M6cjaRBvl6fc6rQ4oHQGw0hYZKGpI5Tz2Kw2/ya2wBF3830tmoFV
J2BRnmiTxHUhpOrYv25LpyeNcA9Fub6V4jUdmuLDlrKTUCl+tVHWy0yhixS6
Lh35eyFksNi3hajiV91BOVzL6XwzGXpaAOTOtba4AZp9D26eaDRaCATrRAOj
8lr/00kvonSiEsEhK7hoyf+xeaNCVJegUIDpTIVTZyXAay7Nu5HdZmRC7tIC
zss7rV9D5YA+8PaCL40PKRkthycLW/KGFV/L2SSGbLMfWM0ddD1KS5Vrqeoq
99DGA/Xv0zvNQnhWd/LI2Rq81a3l4sjVS9xlNgaNnou0oYZ/8PHFy2DdpSL6
tLzPeebFafJOPImSwuYJuEzM4jdTw7+RzTn6ZDJ4eCU8jkKj9GwIA56ga1Bj
V2lX6lj/i4w+ZoYMGZYQDW0cObUqr9QwmXYPOnc0Vash+1GMRd1vGc2ZF6QL
+a4wywrcyTdYdzxBbQglcWHwYrP158MyjPMfQGjH9dhN56sjVug0yNeAhMmd
vsCY4j0ROgA1tEBJB/V0pIgRp5M1BSX4u4Kr+hGpmLK+ZkEs9+XS/lwlwsSt
IIItT/fdFpwW0Bh4yzO9o1R5DRVOhH/mpzinJhpPw0VPtUAx5+r5VF1bFnTr
HUjLOMi1wC7ygnT8a6cPhxATc9Ra1jC28ftG0b6xHhLJrgYgbzb2Wh5RoqIa
GszuRER12ODdVrbtLSk0C2n1SjZHvCcXajXeia9b0xzTfw9JZOiR8aTaqzOm
wi9jANvG7IDVDo1WhqyAbVyB/h7fkVrbb0Ne9rbES289pJHkaQYiWdoGPZbS
2OwiqbvW3Rqx6RElBFGwjjOw5pNpWutpCy05Rbnvzttbdoh1bOrXf1oKycKh
4dBnoODC1sZrU3rCEJl+A+mfANWFrMZz8RPc20YVeKBHI+0kb+aaf8un5N7P
IHxZxPRmkhDvba0cVP0kf114h03iWsBEZ56+f1e6bUvarzXXYvfjKSCXbfcf
3NK6vPxKi0qBhPWbTRAQ7ZZhAkMJtJ6p8RBqe6rMO3hRBUwmn0zuQF1w7RKb
IU1LoRw4EgUpZi4keGRWUuUB42ekxUXWWcmN8xKB0eats2v1K/hL2Fh0Y8D/
mcUEdva7Ete2q46/Q2CwIWff2Y3OoM9mCqvXceSr5/0v72xP7CSQa0vQF7By
u//ysDlTMyPnsFJPN10c3kZrwshxWg02+mZbh2zIGD6/VH6Z44mnsb2SbOwC
igO3Jqp3Yu2wJLg8150DJ6613TZxLRwk+WidfznrOjAax+MtAMHN53sGuTx5
mMBaP1mJGGWVawt0ZOfsk3xNMCpJwAKLwOic01wtz1AxML/Ne/qRJLOMYnin
gZpdNyRPWAykfVZXPhcBQxUdQfiZ74Gi28uazpmOvJfYaECJqwpEsNQ/RABY
VidF6UfailYv6hVQc5ux+6JGX9+UELpdwm3EW4u3h2PMvnvz0652k5nhB3zr
QOy8Ear+l8DaY4wDsUL5rwb4YiOWpYLuhIYi/PXVGqTPovXsCpOtw0wySbUv
1xI/yZua1EAqUCrVC3PVWxCQLojhoRWJ30T4wLpQj/aBMjjRtLVCDq5mm1Ia
c2AzSGDVExrrHELEdogB42KjWppSRZ6g9jZwSAWn85XQIVjmYMp02sES5hMO
oVGikTRgU8EtovtR+8/vRjc0AEHau8WDr7PZ5nWMY+jt5Jmy+/0uvjqMibNn
OTh5Hoes8ZauSuZTE1Hv7HYgJXSIIoIwBPOY/GX6fawoJV2WJwSifJ3egEse
H8yk0gdawFfGlq2W4mjlXAEFY55rG6G7uHIhSV46+Wb9gDhGLSSzX1t5ZhP4
1WSrQJsfcoUW/f4Tmnfu+D4Bqq9iEqd8mFSlJCZOOsIcgIqWLPOVarAXKuX/
sJ5716BGmJLWv6gcvbrNKAMHG1IiqgWla53EKx/8bd6Mt6OdsUR+7kYz3Lju
SYIiGWi+KEHlRXc64RsU1DhH/q8McMOR1D/TM1hea0bLOcWWxIbfCdjFugqd
ncpgRJTYAt6bgVNlzcejbjJISnrw7J6uyCpap/jXETCsLc5Q+7oA6G06Fk+y
7YkpEfqeJgMowUs2La3ljdOLDEnc012CnFCCdCOnHRGANBI/l7H0x2/5Tfpx
l1q2Dg+/FVwbIfJatTpanXq9RkB6jmo5zqJf3pYRI05tIoA2x0hUmIpvOt2R
PlkOH7GkgAk7lj4YWMaDZsaku14Xhupnanv6TeQvjiLyZJVWnqx2HDxoZGCs
Uyq3jtGCMxtFam848gHra3wbob4udNhVCvIVGGkiUZPfXtmV2XdxQyFrDxOn
vIjXY3FctUBJfWhpOqxic+y1zWbXtvUyOu9W9k7nmj98BIWNmmfnV5XhijlQ
ber44fkkyJQGqNEKO3xAnE5mSAGdz/3G8JWO0R/zEDTCr4RVee9H/CLEtaXx
ZzF/Oh3fS7U6Hq2KXVmm1MhQ9IYMsBbD7har+kddQvjM10XDlG2RJ66X5weh
Z2E0fap1NT3uu046PBqTwVs56bE1oNXMrjOkNATOGvQnFtsDQvdEqfz/ZYGB
AdB2qmcTPDcNDOKslUDB+ItK77JNDsmn90+L0YxpCtN3I6J8CoB0KadcneWn
pXTa30bRgAxnpxLWNhG2vovWxfYKNtdwhSN2DVb7cM97W/fI148EfL7+6NWB
XhsVZYYcaD+agg0cf0BcBNxSoFSYdKRfOSKtZOFKCKIAEePW/DZtf4KZZDTN
G2h4LMaqdpj04qLZ/u6mPpPKsLbqm6O9l7RzHYQUOXuZErK1RlDBROTDp0Gf
GfKTO3DIdaCrkOXWeHPOdVcWp+F0WrPXuipi0J2lgGAg7R417wNXHLuvEQWa
BTShvubhxi1SbBpcJi9Hdlw23eJIiGSGUG+g4a427iGdESFeixKx2cNLUuHA
POzTF7T9Am0AfnqfuC4BuWjOaXXqfqVemYRHK9pFl/2e+0ge2ccSpWznbAZU
G520jNT24lhJe/8I4oMcB2pgyZMGuJqiyeduWsCym5bq6jzpeofn3O9E6BTy
NnioHHYdb/HCeIIyNGtfckOyOf58WmJAqmpNJ4ieenVH2i658MrMMsjmbwtq
wuTABibBZJ+ijQK9G7ACuAc5UO67LN1rEtgGUv4f+dg6QQIeE5lU9heiG/Po
j95EK3I+yGCP6wlcZRAzmBEUHwTGfLRh85lpxVj+WPqoNiCEU0suSan3Bruv
40YGeO+Y3+9OnIi7wxvxGQHqhaqJps0jTpBsrGSZYjgWJJbVby9IlOKnr6qL
cQoyLL2hIcJNkofdv+fAp9tTBHEDQOxKofaDyp0fV+ONVrqNvF075Nntr3p8
QHN7ASAxtHbLR3wYuoFHCWB7dl/4kIiF233vyDUJJPHVkq4yPY37isPDGYpr
5VZzkFUAPRl7KhdH5P2dRzK43Xgome6E7bpc9Cp18DRV41tOn1seEFmQ7IOs
yWLo6ZDc1kaiy6ggeV3RnxRWdqTGO8nhB3Cht0WqLMBlmNVvlw49GIOMkmMN
ojDbjDCbb/JUIRlHZay0ZjC5ZbTFynFTEOmwdgotP3G+ae5t9qF9gDYMi0aU
wmK+gn+WoN0Eu+VZ0PEpTApOFdGziQMFvXl29SywirMHBr6tcP/ucntTG6h7
HdbsFkDijxewtKr0xwBvcZHZHPblehMRfbZfBN0RMs6GsOormrJ87AshCee/
fyi6KtzNLSMHUg/nXzVDALcDcE2XImVCHZDF5WCGSFNQR72FymwT5usV7maD
7rrL43hY+HamVbfMWtYpRW+N+V2QICLcZ18obCmFY1jkuj5eWnGka0asuoHu
xjOUkfRCMA/m/tK+0GLQd7/l8/4oetWWBkP1T55Dk6EO/9Ds4n5UC7CW5QA3
1D7lK8jP5d6VuabebHgUXLpaLpegw1ZEcPrN8a7gur0qEcC2u2PZNtPi/GXG
/TifrkCxa0ULFyTmLqyDJ5OuzoriUdc09fy+OtwsTuuA5DwZEX8kxZkVVj5V
o15M9kPIArHlvMbH3+vceJrqwQ7NtlKCIcIbLRMqFFG8qWdsYpC2ylWMO0ob
cCAHtg8TFAVw3x+cz55mdv91cVC7/UPujvUqWrLU1jSx6Kw3Ja0ys6rWlSmE
QZt+6ngztF67ZbfBATZPyqKhYOyLc2KzT1wM7iedVYb6o7rq/lpWDqf2GdCS
vOVAQ7nu5HmXtLnC9S9YvaUhRh8q9gRlhzKkPjhqm3GwIwRS/qT+sHJmXAyO
1Kv/BWQD8IwN19hPETGaKrZ6eNMxLAARBDbzDv+xiHk5HxScn91Dh5a0ropg
6hP6EFAllM45s9vHUL/2nM1GXdahiitAe1TPvM55iMVC4CQ5djZdNbPtOGEK
q6fnuAyx8nPK5qdTmICjpw43mjwK7rDp7H152l2YXrskbSI55b2yaGB30Ck+
gB9UmHPQ+gfqNDXGCZX2+V7MCLECatQluricjlaZBzucnnOheCQe8KTZJ7yW
9rMiOBZ00rQG+ibLuYX6PjLyorc4aK6K0nU6TbtxayOr6kVqJzVjDXC5XD6r
DVetR+pDvrmQsXziiZt78EPhsO8JZDorq1xmaSCz/PtIFh4zWMffm7bR7R5E
F3oKHha8qscMpr89RO6vbEbsHnoS/TAeTHKtxFPjCbcN0N6ahdHXLn65WQ6m
FXGTjF8ItbgNGB/v+sRQ+21bAYp2WN0xF+6ZTnsqFYYxVnV9tkJ4u/tXOnFp
2SiIuwz6ybiy2QdoBCx1W3cdY4dLUnkOxr43BUT7C+niRQJYavVHHp/8O5E1
3mlPs5TAXmAV+odoi8v/j7+7lBz67UJY3Z1CO3EaL0JBfn74lZnrCEjRo+MS
r6oibs/6I/hc8q2LWOnRla/4S17Q6Ni5jeGOonZkTZujNsFcfYcdhINHgvFq
Hp+7QGDqvc0VHoBP/Pk049HZAgH+3yzCjjhMrzxyLvv3nVN8HY7scfOG5C4d
L0EKyOcPCI+cbJUm6z9cwplL0cNgMHM4zGmqrHQ7KQO1HxwUOpc187fyQGjB
vE5BqICoIYubB4a39oxuBVLXTFUuadBSFMMhi6YgtIg184Z0Uwk2vf/uWwfD
mNupCOco1Qzi6jvrXQzFJO0JxSe2iS6pRQyJYqi5nLCi6DVXdJWEttfd8+DS
ggunLDQyO1ViApvILb8KWu2i00XICdWwSth1IWZKShuJEugnPE9pynthQmS1
LQ8sAbFtBkZ7ziVAA/5FkZ7MCDyZCMLSlUd8dymLk1i8sUiZNK+/pH7nBHEN
uPlGHoj3dG/yNd8MkY1Egelw7dRt3JdmrMj3Q5vf6eXozlfSnjibbYGjLoSQ
5Fm0RY8yycpzG3JtNwxagbvmelRsUXdQw4cRAPrw7KuYIfYCeILSzrPEFq8F
WgwgpXKzyYxvJGRN/uffvxzkJG436JRMfHBrUhr6AIXDuaVY2MyEiO8dY16o
13FJiYmPztRTODUpYmRVKgFVbFXCnQ6lH9MRLB6zgQoWMjZ1g+nThDIJ8yVd
PTf1UI4asQSeqsPEv0hrMRtvKymjYrYPnsJidEzfCQbeedO+l59rkfUFGEMf
6u/dAntogmrdovtq1fp8xlsot0SJS9Q7Khl9AEGBjA59cobxXDYoMKV5AZLu
DQ49Nbb8u+KXlgBlz5ggs45FirRycnyE+PKHsF7aQaoQtCa6iF6WNXvDhcoM
CIXoUpGCDf7lsxAQDj9kSwwJiVo7ho8/fc61VrYPIkhOWW4+WVDqOWJOEBB8
YYle6ey2/ietnPH+RGJK/DOaabSjfCdMlsrPcyMDVKGLoh897aEKLuZ+T+d3
pODlZ0lblQfa9ZPmjZOzKS5OAdMUHxph12a2KuuyzZ8sLPVp82jXqd2OQSNK
HxZFsYdq2WbSE9W3lTe1+V1IWccbbzPsI7iPH7hOndjfTEAoWiU+ERScm0dG
WYDMzwz2yCpLOs2Ej4Nzdw9XTmtv2Q7AGn57y4EgfKaRLnccDdGLjZQexEDf
PyQwn/02CfTPvsViXdmi8wFcsBZHhuh83R+4g8ehib9qAWDNeLySiGaSFWBz
x/RNwPYUmWo79af4P8pP/KyR9yPiQ5wWSNXdZJ+8kjlMR0kDrWEJgQpf7SC2
TSCZ4NiwFmcSC4qedD24q/ifyCEe2bh3Qmb1qYtuj/pcaPXWSB/wkqTcIrs6
9QzyBkFLQSexFXqPPlvHFRV/FSC7L6V+OvdaLkpiRrXxEATwOimGNYFqbZwh
jsEbu3ZQXcEmGqkiLOASrfT3YymWjzHokH8qms1S2YUMb3yDO+w7bYsPnv5q
Cibiq7cZn9jQTeGDxm0laHzAlXbe+vMIECHamMXNFqW6RrWKaJP7/5f/7edd
IVEDBo/p3zlJnmzdVXNCJBAIvGwBiMVmF6WbqHLeBH0J8RQcw9qBC80zyZFj
GcosPExurBEowGKfONDMnCuZ0kH2/g22f3FTuWrvRsITI4Y2A9fuhPGWvyTq
tU7bmeyxIUSfnwqNhQ7a8ShjKGhyt04aBOZiFgcR1xYgrVNhDW6fuDkNADSX
54UjxOZ65WfKL4ybf7ydYjy49ig2SbdHTC8nqRbvEMwH96MBiJxp2n/nAmza
djCvkqcM0KDzBZkqWGaQ2srws0t6Owip7yaqb6NPtdzTI4m+7KVkrufUqDCc
EDisAUQVEWtUKc9ByABpT71r2hskci6fYE7TXf/3NtwQC31+PeDLnFIkL6mH
jHXLYPkLZ2GIYn44G3kYxk7UXhl/SXaTugvISIz4cZhYrBdVTctv7785B6HQ
KbmBB+o5F+2avGw87pu2lwVmwuG8Lyc22m9DwB4Xcu5+4SWz7hPCTfafnCbX
Q9U8LLyCWuXFzqUWF8TUr935JpAp5IKNPOdZ6o0S/+c2rQtzKdeOz77kfvPe
pZub3QWXuCGyPDansQWUbAT/6AxKHmFA+75nVv9Cw7uEoGn85rlmjr0+MoEW
RU8VuxFlMb0pNidNcmVPJ51CDipEsDfL+2NS7lOLtxZ02QpfkmTVQlx+PyoB
pw8Q3TVlH5uS2nAQ2e7JwBRIEZkXk5k7mUbyveH24Nj0OPFs6BaAOq3PvqJh
DOvuK2jv3c5pKQLAfGSO7oTfCaGru+hX7ug2BLi4tmA8l0t8eucI25VdVAJl
AvgEjfxvfLL7TET3/7DFfgGR0Ne0nzJ75beJlCx4SYzB9UjnqRGKSVbGvL0K
RBBx/FoZsEZfjo33OWCfVo/tntXMgHq1mJ88278OQDD7GCPIKhSIwkfq44P8
iI6Rd68512aUgqTYm1Z5PSPdecI85P/cv39YqXA+MG/7MTbLIpGJjrvuk+e7
MuouLUc6VBr4RTzowgl2iU3XxCJkBex2DCsehk1fhMzY1TPZFZyooN31/MXl
uk2tyOIx9DSSnZ7x2EOYWIWgswSERrvN7FI8yLgFuy+EQmn/6ZjiNdxWflTr
5F0/yo6KtkfzAQHfMUsGwzztrvtFVKkmWNMNe7Rxg9C4LuFrrnKlkuJHSbuB
/5f0lknUpysXfb97AAosaSTX2nWBgWgZ4mAN60VT9HvEQ4Vlatyh3aTaR0Sr
1hmKG2iyzrvFmg5V0oUOdsvnBnqHZvp3HJQf5KDYunQNZh6AJAo5IBjit1bi
5P6RtaWJjcaVur1Gbo6np58Ch4lNa1uhrl6/GVnxQsgLEGflJDRRWX0hIPGJ
/fSIHNkiOJ1mKr+iELItaKKU7MdVFf+iwzFYHhR+ajSlDcW75dpvNEQ4R4Lc
4u5aOLgwxIHCLqGdGTYMfWy4ZnEUobSSCK6DuNCTAyDYFxfYhLTufwx+cleB
374V1iPeF7qlJvnHzf5jS3c5YTiSxzA6dalK5uZl7QX9/xxMaL1HkdwhZx1m
uIi1AIMqn5yoa4olaqjQMCeAdxUuBOFZr6k39t1X7/NKusCxSx9RLuAmOLb/
jUAhhFafO/1+s+o8NZefmc+x7itOm/EK9nsJY4XkIybTEsYZm0Jk87jE4LlG
oQAqA+I0TSKnFbZMJFZqRGlke8a3dWsjCip+KjnbDgSrLvr/J3ehypWTkg6t
cprLj73SugCcPiAbHyVhihctbBa8+W4qYEyk6CeQkqoe6394EeZmm4XwqIwh
tinqlCah3IBJ8zg78kbtScehHBxksoPgLuXyuyh3vnlMK9ecOEryTnZSibnP
dWuXqnlPUeoNrFmXivgAmb9DuttQ/UUi65KFgHWSXiiApV95gdzcv6Dm+Aqv
xMhhaA75e4lshdPgmPTpEL0TffVYMSz3X5wEC2UQUKQI1VCXjB+L8SAQIk/h
uhiXATaCzLJdq3MEUnaYrAE5x0ZJUkIKVjOleZ9OfYoaRjPris6nPqVuXM+s
TozntmD9T5wTkuyPvq1tUreKDZqZt83vVwY49QEyl0goG2DXWVp5KLc1YhvS
aJpdZWQ8b/kRGML4yWTyE47HaimHr/uKb9NI4qprPI9CtDnhxud5RgZoB/Pf
Jiw1gWI1MWLmFbw78w0Ml13NZIsVPjqGejh4cZ+Bsk6mStKZzYoQ8U+Khu/4
RCyFAYQJeEgBJiD9wGr5bY6pE2+VfkfA2gE3oqsW8DT+ZT8Zc5P0RzLx3ZbB
QoQXxsC8ZZ3qiN9d8SIt5FrGz9exQ6TZbRyVmt7/I/iiBLxshrla3lt1D6sh
ZhxNCX7Kk0sxXMgmvh/i4tCIExW9lOBDIoFzKwsDER7wI4GUqaswBQj4iQIE
S4SPoX2imAGxcZM8xEj0w20IF0x/Gs0vTcrJPRgcry4mhe9QyXpz8rBQTSpM
QGEW9xba48PX/f72y9g16rf+7k/UEH8eg04aarjv8rIsqLuxpl9WyKM96T11
/H+hI5ybX26gsbgQc1cMxbCPA8zegL7UU7oLR7xToMoBzvEshPuE4nI4me82
7tWfRe5xlzOYxrYTU/LaQDXgq4C8CkYlfSwCpeQTuGwJiZtO/YFZo1jwe1GO
7WWaKZPPd3vxJaBXCYhHsJNSmjSGEthdV/MR28jaAopjuPz/JPNh84Qh1h/V
U+QqSb+3/w49USJwTKg+AD6s6TrbHG/w2wg0zZmoUpF6IECYYad6wiBNyHEd
oORmGJ1PsEfDrawj2sYI5u1jxCU7/CnP5kP/EGvGaaYNwwUi5JhUXHD35Cfv
8XDdDj2GmB34lCxYNmmAZjkQ/Zd1A8k3lj+7ausjQki+jHPXBF8lk02A40eb
KpLrJMdFW9bfDIrSsbjIqJAXk2tuQitWRJ37zkoDwDfApt9XH0Aa7rIcw7wQ
dx+bT+eORzAtyQjriPK54OM/EPGheP6pyOFJtcj/Lxa+FvWn1RnBJKZQAd2m
0ZIiOO4OVk+uwx8oTsWuBHO44sRjgy+7aplXI1DXdXcvkj9R8aY8FK8wqpCx
eTe7NB58vARwitTW61YzngXS6DAeiTc6b8YZYLtOVPpR6Av4CNZwnEc3zW5g
i2ZGdB+CDrsk1e/pcYX9iTAHcDgzKqpxffKIkvP4DnS2M3wpXJu/jdytfpw3
Ey6LIYhYh2W9GmmiTRoehDGlqJ68TxOJS594sQXl34f8IKq3UoLj7syxC+E6
4M3twHonH1Yl73oqRP2Guqrhg6965jdggnCt7GZFeXczJ1jFRyUNxkawzf3L
dglCbw+Hwq83IYKfTRNqAzVxBBMo3VQMLubMv2tmAN6ii8+aFUvKU6gvpwyV
ww23/FptD9J2OJxKBkbbvtOj4LOe0gqHWQ+4Aw5kV8b9j3sNTHrVESFcPzSc
mW4k/LoYM5Izaaecw2vTmRQ7hCkOm9K6u8zwvxL0Y9P330034qd+zpdRu29f
uAE9rqYcVo4iBGJJ0XkD9o6KDcq70yqQBLR72KGUt150pMR9CWLoWMnUAOTo
I4KIqJhURnW1vc3EI/sRRw1DTEO8GZ2l952VR5Mxe3I3jazbyY1IFD/uZjYG
B2TkWkIgu1TLfchuGL44JQJahpcUiFEbdRDWN4kUwgA6UNhCr2MBFmubAoq6
3Vr70NTa8nowdIgM+IUhnYImSPozDt/9NOj3//bDYUYAfLxa3B+e3c9YA4sv
DjzkIIMGic5qW+DcoSDTWFbVin0+lS1GoMBYmFB0afbHoylUZBu5OHejFNJ2
ikAGWCumDXt3pAVdkO2CAq+ELdBXUM3ju0ADHSs1HPcYR4M/jRfnxRlnJ54S
WF+qMF/O001ZDQB6pSA7bQAwCqb+NqiTTmJrVacz1I5fmo5IfcXAzq1QRhZU
bzYzjMRPMeprZX15i/FXLcxKs7vM1vmbqS/PoWZ4ZRJFifTRwEKijEQ4/vh7
gIK4Fs7H7diVPbR8Y8Gm/GRoQ8r2M1x1mmD33OnQR5hxekxypHScAm1wQM6w
EHkkEbgAJuG4YfF8bHSZsjkEde0llevlWO7lwpr9UQ67DsvljuCWigy/T9g2
1ktfXkumIZtJgDaN7O4Pa0zwQv5LvTHAz/aOOTpt8JmwTkJngqFJ9b88rZSy
YRJYSNRE1RPZHVzBJtzxvkUQL59280P4AyJoX4IZO2ArfAPPDi0lj9miGEmL
PkETKJOEVA5B2b7m7uGrOnOoiqQDKVhKV4cDzB5WouRkoGLLYT3iC48OrbKY
G62mOIwkBILwGXwfgCmcIaUE+M1jeEajbbi6FWFxSEP06sgvayMR++AbG/GV
k08+4PIm6qIEF9IRjVyGSy3jYdMwP/OSx3HMp/qMk+0SxunOQzVkBDN5qqRq
EhJOIq5dfytzLu1jLHG942bPjt7pUD2HyHFkQrGZsQmSC24X6KNKLHYXX5Kl
poYEBWaZ2sPYIDjc5CNgsdvuvK+Icj0riED5AdZViwMucIYtTA4aVDKJnZfk
WVUq1gK7n31A4uLy9Ffkf4WBIkXpzBbtG73tLTaHzONqXbPaGZ+OvzNrzOeH
5HNEtyUONI2dxauu4ttgCdY6Zkr0vdEi1DSeXt0DTrB61hhS83kgS/T4UAE5
GyRjuVlbHJnHOjHeMAwPkPagUnxsVLkp8zQYWk2aNd6gz/od5kXjhn3zaXMJ
7g3iOTKFX/MVanL5fq46DKTj43DnEnTwD/7ySGdxrpLBycew8iTdj+1kMvhS
E/bnw+BmbIwl2wMyquT6lkC55XOSUmo80+n6/1iIjf2haarloMbet93/1m8K
4sy6vs1F3RiX0r7W1ZMJL6u8b4Bbssp39lkLO7b7qhj8IPBWo74Cn3cdwRP8
dFbeIc9XCmRVLnlJucvXbbJBOTVKD4flH76PgTG3y0YwkJBoYwHa7JqlHm5U
W7ypi0FFRnvJPNSey8UDzW92/evad0zbXIVBvK3n7xmH76iddcgpwNdc99SD
kbxIE8/SdB9iR94AjLo5Z+gKdkZQ87NpfA82+s7yaWsFq2zn4n2ZnRSnNq1p
ZMu8CnJQ80adXH2XOH8nLSBjWtvKDhTY6+j8blvvxg03nskJ0h2HIJEXYaL1
n4uhXPYtA35DsSEuBq94eCP5QhsYi5XoEiLbfMrXWxC2SyQ0fOkzjM7wHl0g
KoYPVCd/VOwFYFMS1dlGI9jEIYOUrK+YaZeAOlTXH5fgcLcuEKru1hF2xkii
5s/PWvkMVPIiwvZfAOnmbwcHxrz6CzkIn7Ph8sE6T3re3qHl+8oLDcPJK9zC
oJcj141WahdPc6rmXOF5UJ5eiwZhuKWdr9o4Z1jUn7AzInlEm9ZsnDR42815
lUlLaPo3+Gr7HVcRtONjZh1ie3tZuwRHsAgj1migkqSTYGFRc3jFcXxjyQj9
zjpwwkPyo3dC1/9vr85LOBEEvfgPCd9DWWVR7pzKB1/nnKW6RJsp1sNCR+o2
ZfHmrsySyf+0rwxeTfHEyStXRskLbRkEEPrVXYONz0Xqsne0iUZvTp4O/A6t
Ce2Fcy+1rqYdR2Ud3Tw5LMXtSgwK1uC68Ftz5W2yyY0C/W1eatMTvA/3tTV0
V8pGeLShIp8fHQHluxOClYCH+Ltw1w2h4xyQCkV2XO0Yth7zzvc+G7tugny8
cjTZfPniuNY9wMmSKRbfh3D8M0OU9GnPB/OwVR9NStyqhn4RB/ZjXmW9Si0Z
EW88+xyUIAlFxNr136G3b5V8hPvZPPqQrVvgAWq/rWqg2cmtYdqqdtUUcXO7
N1j33JFGSGZzJs76hRlr0Z/XkZGlgOhvI26aVboX7Y1nbdC7TwtwLBg5CsTa
5vkry6IERGg/lwKtP9BjaOZKW3FdZeumIRH1i8fndtv/1e7dGOW9FbgjfRsl
CWepvnhmlq6tLEbXixkn2Oc4dpO7X5PUVtQ41lL5CJm2I3CPphNTdk6sNxSs
uRsLORlKW2WBsscdoSOvfrp3eVlotVUzIzO/fJxmEn/qSP9UUVLSktg/zsN4
pLJ3gtmvY/t5eCZA2DnI++atRT0CQwTTwwIyuY5I3AXV1ds8Hl8VYkGeFBNQ
9MRwf8PhpYH7Eif+J12aBMd6Aj08Y6+FVopQlyQCEvDzH/J1wZ7SKUipujYX
OsgTNW9kyfSDqes/iqSW7C8FpqpRWSmIWHWA+9jodtiORXVb385mhIGEWkB+
Eu4gJeMlevNtfRtyxDUkiL2pvjxPZ0LmqgnmfLxVkahDZfQXu/bKuxZqdJIr
pMk/HjE38JtJeVlwzKleKEZG5MYO7wIIvzzEVmgnzTTv8qKSRkTR/brkjhRf
xqElDYo9DVe8313WNdMlMY2LiKa55ccmftwK+suHIO+tFNE7Oj3cr0HJ6/7h
ULuvIpm7+4YKBTYg49JNxV88DRbhnMmynMFV4sHdDKBzr11JkWcTbaG/a10N
nsKVmCcpVdzemKTY88J9RAQhi6VCEMX6jpIHRJqErm6dIUF8sdm09Am7vR30
rw+eK7HnCt8Ju9dpYDbwFgh/Oi4cUHwnGGYlgBrLileEVrRAjpnryFq6Zx+u
dAJYy3x9cBJfRapfs/uYuZVqd5QedUtGF/x7cXg4xMJZEyO/gbzkSlk8wGZF
mF6UpNkwyGec5IYAjDdU3MeZYyyM3L8kJfqGaSGaHyvQjsBJ3grgMvp5HgXL
oWPnNOCeGhaMZQWqAwkpu/mPAcecCgz3eCNVlPHAuIJON6yOMn7ywo5H60pT
oZqOgowmEVBzktk2koO/2dm9f8SBsEqnTspSaItPjMmWBo2Fkk7xyjyfteOg
j36qTrTAtER+7KbE99m1hNzeXL3ahegp0U2EO5MEASbY66Kb+Xz8FN48wySj
l/PKVwUfeh7koX3GLgtLr9gKi6OqTtgUZSCJdS+fJ3eqkV/4RrCWWH8GnO39
+ho2zLYjzkJINUJBCYKvmzV9Ghccf2FAFkNz4q2TN0q11h7QLS74hFA/CU8p
S1Q+DRuiBHJ0j/xTFOOBYMbwdbM1AgNMMMsPLxmDJQ5meTlCN3E/P2hTBmaZ
ZQ/DVCPM5asBF8Q0MkpTNIyz4cpoJ4+KTdVdCwn+S7gVUdg9b5OAZddIQAp2
WgHCUuonEGMTP/TeGuUFCBVTRNXfqvhU+4Gby8AveYWRvgBLjto7jMdy060F
E6CVcB2RyjRpnb/+CzWaeVLySK3Lz6vFUCZDEa3/+B/jCS5OtAQBZE88XAPB
QydQusyYpInHHb1orE4Wi0aKwvFqyZCIY+VF2iHZVfwK6sIWjs1tQZt9tFql
pgkoOCwsArqahdqY7N/NqfWoy9FJFdUpEFu7mlGCe3DcCJXIjG9HI+nPG1E/
4yhcF8qAk8gXw4FKT8ucnhlSBW71L9F5sxHvIC78lO/exw2NwEtoMgTzmNWB
TDWCVn9BAISkszU2w/dh4KcNe/cmKFnu3y1ldgnYM90i+mQdMlr+Hf7wssFX
/poF2oJSiNmPh08SfBAsnGO7oGjCHeLaC9fgolutQ3LUV4XcpobflfQobXfa
9cGkE6Urn61ZqgvHgHCQpUVOKCiUllNt1hGXRZK3RafMfHFeb9AK26VSyPdF
izfkO3X1WFlu7DV6TQnpWxS2XHLqV4lBI/9lqLmRlgSiiIutLjgg55WyXiiO
vNLy3Y28zI1usTcYqpGxboVgTe1BR2tJQIc62JyKyfmK891jR9tjGq6Q7HYf
Wyq87Bt/ICk6CiFaKqn9Or99Lh+vk7Of8Y2entxU76GJTiS6EQaUxi9a57yL
tW8haeQGZhVHgwaxjNbEb3l/YN1020oNXDu0io0y8qqX8UAEl/XiMBAKhZW0
wC5EH1rQEl7YzDyf/FOSTyPbcO1rmNBKVNXRS4Yt4kyPkJDkGi9n+l26j2Jo
nQvRg+IpnhfoPP7FzP+P3hkG/p5+zN80dfCaJLvN9OaXaXCraOzAAX9vQST5
w0/DoFbJLTtcxvFmCyC36xL08E6gTEKx5uJF+9nPgWYcj+XAJuoN2aVQm1t/
6+yFRt6IWVMLkEFsmkQuzJwywMGurlaAXgIfie0KPVVQDDr1WeIvEbi2aHp6
uzZv4Ac3/c3CEW10e7DB4Wrmv+r2tR1SotGiJUyjRejVWG9kngdSsMEE4sQw
T2hvWyHZ25l5LihCBfGblQ7hIGR8KEFhEnS2xCMMavfJMza90VD0Ng/wc9N7
K3+G3Z19FFSCxhmmXQjh10Z3wCxxOi8iMEEYCr+xz3Qi1e65zN3oO1zl1Qra
Gf8INCM8+sI9x2I8emXGEseed9M6iyIC3Ih0q17FRaEjoj2fS1H5ExkW+xj3
j9C63LKkYSJS8cHsh9HaFqp+4x2dFWUXSrbm/ZO39HEOIU+m3MFYSMheKgcE
VPhLghhbLU2ejTby68em8rgOcMXh7BKYMPbUk1sI+oRNAMYM2lL0SQL2/ZOa
kRzPqfgB7X17NabQPoRCxqiSzrXBX0UIabemC7DiTvqgVQK0eqMoIMWSd0Ty
96MqYar/1Vcktlrrdie5ShdJ6mjQlQYtqIgsFA72R3puvJ0zrBFB2z19R/cR
4fF2u14LRYd97ZXibolhuDpTG5MNlBWGnqUT1q6e5T0j7ciOFKKYXHInZLqs
i4yRRxmhEY9Av5fc4Q7OhUREQo/nMMkaj1GAjJZDjqqqe9Wa8p/cfbwiB0yT
qaUCIdOnaa73Z0P7dV4AUgnbEFk2cHS6BdZm2RfT+qXDN4TwqYX6lyJnS4Nw
+3R65xQnHUvJbdj3sqj/M+iGlmRGc+MsKNnnL/MnRb8IzcaLxbQxIiZQadOF
6gndMLOn8UsaZTNa9RhNzBXTADluaWpGVLClaIPL6/1HDX+otmXe8vtNwpdN
apP9t2nvH5BEGPBzfuSHserlB3NVgeeZYJQTR7M5VJ5IS0dKVo94Deo0ZM3H
cJZXks/RBkQXI5hrgIrt89IxJkPwH4l/pzAYXXRxcdxDM+Um/gAxzijhR6TK
WnJMCziLiyHJ3UmM1dKfFOygzGSjGkQWmUasYsXiWV2AZ4jM21mCaUUR1c/V
5yMYWiuvQnASCXrAroACITXWcdpjzvw+t5DYU0Ad1/1xyvlK37M9dQq6mqMs
GMnWCmnZtLnc6wFqCQxI8AYQNl7/6qPcsKxwL/RJIpJvcgz21t3PkjQf7ppr
nru6Cj/bHU3BKP5SAvEZtQn/7qxvsoDmfwuutOTTDNynQNJ7WVzyg+WLcrfj
SiVFGdRFb3DLC6QiFUul5v1vybSNQrsV8M0A2TSmpNcv6MRJpDC0mEum5J2h
5IPg+5AhyfqCxYUqVpBnv6sb3auxrpEs+P4BO5GHUlGtAkAXEUODdzZJLy9/
e0Bie7Ov7cERQWTxQsDT8Yy3Ttqeg5kYA+QPzR2VKAQ1FcSuGEM68YT75bFf
YmdxM8ZamXcPRNLn1GEejnnS9NwdYMTU7K/UfSik/xwBJkNdsuFz9TnxI/aX
4tIyQpgU04Rluzg7+l0EDC41FNjVErpUQUQvnGstjdvTSfucaJh65/w305H2
dXTfCNTGzNt8ffGUER/vxikwrvsWzaA8qxB8E0PLRWHY8Q3ij/gGz4anoFFN
lY0WLM1tMmFF89B//NoKwJIJFmbQiSMcslERbyUQWTAsoXBo4l+pXlyH+F0W
HEo/sH/oPjO9gxknRh7iDBgrMGhKLewqIVhM7GU1MWDks5B3gZoXOfrMKsU/
fftPYQSNWXxXQJlWsicL+dARj7DOohJx7GQ/oZ+OYkvAtvvgxOWG9dERs5mL
HVprwaU4+OA1+8RFxTEj9nMeihRS+QpJ09i564fkIRjwHIruJ+yziv8rayKo
I6LXfoyrGZOw3Kf7paF4aGiKsAHGinGjxeO0b7VQS9CMKA8Mvs0jmWs1Kox9
0fGOdmuPjp8duvz8X7qQHWkZmQgn9GBYV622e9G9z2ich/opqUZqOMY9Z428
v+Ps88+N2KBlE3ekJ9JcAqhF1Muo1D2jmxGe+q8FHIH+WfZC0qO7aekJXttZ
jNiOoIqSzZQfIJmDWzz2o8VTOWx0HK/t3BIjDTbflWDlucMslzft3jAJS86F
G47fDI+XM4v4fjJ6KSxB7HkMFPXT098LRFJTGSuEYFqy119x7ZiTgKUJoluX
BXXh7hvpZ2D39noAZukJWBiisVREkYCfT0yjXi7stBtSw6bb+lc/JleQvgLW
rjCbnmO/7BLjfXLY99/97WbPWOaGsixAwwtCHgB8bxdQdYU7sJnKGCaXxvzk
B8zDkxnxH6t5YVdgLrmkxRr1t3MC8MHL+5V4gy0dX5aqihT9g30IRgREPDAY
M699Q7ly15k0CEdRpw3Aw8FsN+LrUbatV9uHhxw7wLHR6LN2ihmmjULDOik0
Wal2qiq9N8g119KXOycB7CfI7hHJmmVjhM0rW8ttuYhmCvp+BZlvb6EWCWy6
rPp7hX20PnpBGWKtKLRKf1b5yeWjSRtjHPz5JL82/egf7w57M8jZ+NDFV2uH
BPJPoKBcKpO1wMtvtbLOVTOQhQh86XgaJbRTk6CkKQfpqGzlpkY+bdoyyCxP
Zjh2+boDEP1a4YxKAy4L3ztdDlGRzFZsqhBPfSXvrfgHYpUKBbyRZ17yD3ER
jTyxlyVkP3KewSNuYaSOIxS+aV/3PV2eX37ZWliXmVQlNwoWriCF8JxwCyOZ
a3sETGF79rA7Ltx8oe0XIEp7SvI9DBddKYGBuKHJCcPuYSbef9UbRTbnqcoV
Sr7EF+HSIHZhj3QCVKb1gNFEgWKKWhKzaXGGog2ytEX2tqRERAGVM7mpJB0J
vNTrDKZ8OEEk717m8043twvjJj31Wh1Ywn0wVlo70fKhULJfU0wXxUN0oVzY
t93Trl0Zr37mIw0xMJhYTg8FGgsY6SXLzHj1MYLeZa1RxqHSP1MPm4am1KRm
JkrlUAbIGgxO7XXb+a9LeYJEFErNWpAxlvG/6Uw0rh+s5QzdEdLt4tKTF9SY
Bhp0rA9O3ByA/iQaF7uvATwHpMoRsHKMcsveP7LL0cse1TAVUB3GLUdEh9ZZ
w4Jwc5T4Y4avgllmxQ7+h/TF4LpfJUVo3zUAagxnLYFSR4iJDFFO8FIvqfU6
XnKlVE1W1vLs/MJvGd8/lmuBHoGQl68OS678FNwehXLVNynXbVjuAN7IDdGF
QDDhvFrBQTAKtX+ayVxMpDDraLVJjQy2/G2H0eL/QJGBx2AYY1bmcSp1rEhv
WfA5YK1nQRrTJ9v4+/HemLNGFr1LBZ06gzNTnY/RQmboUsdiB2ACmctiUc28
+KxTktKPna7nLkb/0lfInCgSKUhAOXgxz5YcTkNkBV0eZayzCzQdIqh7phSJ
4wVyw6cFo8aX5nkEk1GG8nUGUwdN8mtpxso7CSgCPHAYZgrrZ0nJVDmZJqMW
f8QvJlvKAGphrMfJA2YfwMQjdne4Yb87lKhpZLlwB8C0jaaNsA9i0F0nhyfD
dgwSVzxnNN9TJEetMdBEdiRAEhcoO1xqqtWeciumPr2yuebvbY8S2rt0khNC
wb3oEaeFL2zhWv84B4iJ8DY/6CZAdkmvtmH7iyopyvpB+gcIRimT+oYv4DTf
yzuRinzsZqZl+JRlSH+kwngPgyYjnejqTW2J1bgLxeHJUWl3MOx/l7J78vC2
y46gw8sNGaFAra3HAly5nhHUQAODTa2URQxqPqo9noDyk6Tanvtm97Mu0p/m
PYLxELGJmTePZJC/2I3myNUnJDaB9HijmQQ7wJIXDFyjyBZRvA7nlAiFFdWQ
X9JeAdNpvm585edm6lEWWewp3ah/qBhPT1pxumXibyB5N6WQnlS+7t1M6gp8
8s8iVS6DKxjIlbF628GxK6sQIvnFOLtf84PmaZLTaHxHaOKnNadzKnFAiAi7
iNqrV0pBIjxdLrnacp+3Xq/UrRUpZKiqQmCIi1JyhGGSIc927qImZJ/PmYnB
mME3W2Alt71/CLryXSDvlF80omKuqRl6Lcq7UnPLTj+VOiTu3Gn+gauIUbaf
NzRBRpq6QZZBCEdJOLSVXYLzNZOURYOLfryE1hFkyArJloNGTbbe+33Xaabj
yagTrvSyFuujMmjFzutVJGQntXtJ/YjHrbw+VtyblWRl5iDmvY5mjDmewA9S
EZ4W6P97sZpRRoa/1FLPwEb5b2g0JcR7q0AGT+4I1UeTa3wT3IBz4qVQLi/Z
GFTbrobg55YZc+IEyO7smWV9a5OJNzhw/gQKdHRSYkZ8nVxz0AudFa7ohbJi
Gd+YEvRg5Ph3xZECw6npzzZTuoa2GMQDogJKnN373sRn1dw3Bmkw0sgBfeEA
l4vaJc4f/L+oK2G2WDPP5GX2OXt0WG7zoLzI8Bwag4nS7WFO+AFygma78xyT
SbKB6cQQcbPMNAysXI6/w6SWkuaNSTPkbuzWouZ6CUZptMRK+etA0k2PegBf
10ub0qWp63VTI+3tr3ILJVnfRdK2CFGmMbgc015qVEakK96M0u0hVHUgN/nQ
vQ00nlINqupss2gnHgRIlPsAYtJs6UCXu4+yY6mXCS0D0d6KQvdTQ/72r9dX
JnlNOAI3JGvJiHWc9QMsZKadf/YxaGpsNu8pQ4Isu1JKHnqrSS7Eb6nJLYxn
PvGsa3BXveyCRDfz6urB5Yy9lmObzQRQB6VSA/wJOUOwL136DxyrK/ppB/a6
s2LwT8qcRawedAzqhXX+IuBuhk/c7IYIkdW37lnuRGbhO4zmEhRIVvJK0Lkx
P7HxQr+YOSBOT5A7QLZZCvthzgqccXMorAVeJiyUacy+VXhEisUjQnieIHD2
NT/XVt8d83dWaOMNJ+dYltHXyix6geIx+Tv6GWHheEcGP/Jtxd8BvSgpUWAJ
T3f8rvCfIDE3k8+YXmOUkHVybljCf5blbu3Jw2OtRZOU2B+kcQIo3A9vyThe
rBxxJv5/shMjp+9LgWNOSW17M3JzbpsajksNhswXp2P+efpfUm4maiDhd+Vw
ojznQAtduT+CPINFJD4b1bJGWudrJi80LyUqW8ibR3+qOWZZKFg/sPQg6coG
3J1V4z1B6ORgaBzMIDRAqnZdWTW5T5ZhrYTdfGafMZcX4hJGP7n5Tht2W/B6
PeXcs1rc/RaQfbPphkWNOuegiyeNRV2tW4Ii5ittee8xHKhloBghPSlTKPHJ
qjt4r/SQvuIm0EWSRC5m3Ckx/Vexxq8UCHjIUhpZE04y6RWGbGl5XoDEGnJC
G75GmkUvEb+Gyj4PRvkc0LDgtRl33/7vSip2GerI3ddXyXc32qhax9hWeBsh
DJabI0sK/HIY7pjWvXuEO4fC6gK5rZfQNEgSZOOQrJO34cy67x6gidqlvrEH
kDHrHBU9S2pCPmq2lPBPkpHxAYoYGsLUGmwJTvXWf2J74h6/rEhOXVKlrewA
ZGQ+r2fRjaEIvwV+uY8xHoTjQHKNPFB/azxRNcM4CLOTkg9PkWDowidpPvMg
adqkPHBMCKeAohplJUsUmFd9dJVLUQXTnwx92/9AmWfFWVuAiGhVSAsQPAlz
Qy6XTUwbl9Nd/hj3inhyMrVs+q0Ig0alYBSx6RgldSsteuq5FKf9/IwExmqK
CFCpIM2hYbuZ0qz4Z5pNSWdNK6EvCWW/nB8nnB8yn+B8rUK4bnLJZ0lD3PXs
UfQJYWh8cTYhZ5ZoqXANEPH+jgriQ7bEc989RDRDrwv9nBr9tWGcUFg/TXZP
2EBDhCks8meIDrnhZDRWNwTe/lPieOSQDfQdSZB7W1JjLM9ajAhRZSk2qsC0
bBMOwhAs8DFCikCITDEPE/5Bo30b/sdIF/WMnebr2CZY+ghNbQv/U+HWV0sD
4NT0VB03OGCDeZZyfOCa7flGxAepPmLuYWiD3PTy3Se1+mfuBaSF+iNyEXx7
xcZH7eEQH5Orjnsu8fhfqIEDhffSKhoPR3rIf1uhV3KjSDJsrWnjxP0HnkNn
ch0xTygXnGx5mPzEtkpE8iIfzLCCKclM1V7I2FHm9II4c91S9WswX2GU7rYT
B2iJlftXH4ZGLA+4ATl3yQttvfx2MoVXbfIfbqMNdRsDUyotrL38FeoxpAbR
eBp0++SeiuDeqI4Vx7glR6o/15xHUdWnLTfsepipt2qafdVeLMmcKPKDwVVT
6PuaF1/JWwElqHEuIVvapR48MdqFy/0/9aLvyU6loGchsYuuWG72dcdOVaAR
2oP3jEG5P3h7hvivYIWD0iHlYxv6JqBaCPrH4c2Gh43S5IrDduBev5hxZnhm
uUBQ6yC5VyNV5kKcEfGCWJL56POd2748HHBGPRD/WvPRdEB5M0xAX1w7vOEr
/KL6cPtb9ncbi5oBi11LK22jO2di42BHCf4XMsTBk1MX7+XeuUkFGt5h5+L9
OcSrybo5MLzPM2S3FV3gy+nVhKotPzQteXjZPiAUJKqIHK68EX0ZTIdkZyKq
uE/yQ3FlqxS0X5P0aNPUn0bQCDsjkWurIe2F7bx6YvdnGvm7ic3lPxshyp74
pLd9Iln1r7A6F5/fDBGBo/jGSX0iqk+r1mOZdFupyXmpZMMl//pCtKbhvluv
Kt8roRpEKRe88knuQevcpZsQleSo/vXvIyswnNECiLGX7vlbqYHguLbBrMS3
8LM12uyEIIqvJp0j3PyTpsKjAqEev/0EoQXRlEIwfeh+IV0WASa8qLIvibDC
Ep8iAYpDZ5sbcI80cc1hLaXZZC9w5FE3hup6GXxDjc5g9+wrdsZpoggIbcaw
/5IT/Z/t9N1bnX2gjgANOF1kZ3tNXUhxLqs2vCeOdwXd2ZFdBXrSVx6K4/pa
mFmYhDnG3wAPTOdl3+y33hs+9WpTYXQhG1BS8ulXFPcSO3IH93nBVCETqHj5
+DXdBuF87hXgnI+PNZPEZ+mLIP3xdiRs9IBKV2ka+fLxA9xuF2RSpGpXjEr9
ogTVf2TUFCL9CmbM5av2/i1M9wB53axpJcmr83P9HSXEApPARKvxouENl9ol
2XBTlh085EbAqRHsGkYN3/fkzb94kELbe9Vp155t6C1JuRUliuWN+yjG7zYQ
cC7G0EI1KrVQCXrDUegK1sH+Thz6/aRVH5rnkbJl9HlEm5jMoGznNL2vNSVC
GFdgflLB5gRH4OR58EAsvXv/rrLf0KqTig7hN0oL92JOtkqWEgBw/zp/hQOf
pZBZ9UaEVPti3gUK9/XBzIoztjRbCbwyswFoCMkH5th7CarNszTpCtjrCihy
AG3TYzxhP8Paj24FKCCyf7pkMnh3dgVq+Z+YacmMKdzKyP498UUL5xRUc0uU
PLZBVJP0wQ9XDa+Lx4q9c/pxPLqlK4Cvm30PNnJ/bvl0fSkfUOSGApduaa6h
xN/c14dGGgYYZdNHHYqPjvdZ5qRshjPPcDPSLZD1Ov9r8t7SxEXIVxxbXqZF
aoYk68xEYKhVHVKSg6RSqNviMgQHROseidjWXkN1uNP0439GVF0s06auzZq3
4Y/n4iuegB/1dWYGpumROZ94dZtb9RM+a99R2UX7Ja3vo/E0g9m4ClAM3kwG
5n2SUyNYDh05PQzLu+GDopl1nQsG8MgWO7Qa/8Grp0sZbjUw05fBxl86E2ag
ChvIwDWazxvzEVsnRdxtjJyUa6gclSNXz6XmdEBqJrspGLZfbehYOKSzJGGz
FLUxF8k4dxEEbee6e5DiJTBtrTu4PHr3p0FL4CYtOphfglNp6KeYFGwzuRyJ
bHmY3y8gtQpptINMic81odYynCq80I4uEhdxOfVuXzEPpQsttyuw27HvIQy4
GWVy/hjcR5tpnPRMHLI5b2u2jhBg4H/Mzt+QC2ifMxQdxCAwg8NPPk6uj7qX
jbKhmDi0L9G1YbCeP+7+8zK9EMC86o3de3sWqsvCSuWQ+1geZiYgJVHtWLWh
FVNQEdax3d+Au53SRvnJExan8OHmeK7Q7Rg/84ccSJV6+ACmOj7D+SvHECG2
2XOdWJllq+2huisZaOsFlnEtKg28SP+dayxQXlvn7rIQNhlVC1vy079YQY6Q
KdEybyHCtO27shPzT7Zv1XeQHyUiYqN7JpofIrgND0TJWSJufnCCA23lNvg1
1qQUqYkrqoTq3K8unTUF+QR0uuqgW1etGSU/IuLNwOlsXTmTbOPjYAgK1A3D
ad3IJpnwPrV1Pk77aBQ2IRgUgSN+wKjRg6vZvfaUGWR9ebSDGs+KUNIsqAjp
gp3BPU/5niAEj+7z1C79cfDJAG82G/YuKA3QvRexm64xMNzQZtPqOL4U8o03
KTFOaxWJC9Mu29QdNmLaOW+qbTKEXEzTGa+FOlnjhqrQhso0sZsnRg4KNKPv
FRQzy7W5NFN7aMveWIJ9F3n+JNECerziTkUjFpB9K+1CgSlzW0pU5397Oal1
uKs937Bi7PsH3cUInz3VIAaUE4A4lwYraP/9R76Zt6Ia5dx6JQRwLqPxPKxM
mM/aFvr2C5hZNiVaTlXHsxuNRV+VL+B1S13kHlsZ+uonAISHHhv8MR/UTl3r
Zbu9UTtb6aVroIEXqsAPu5GZMm3gc30HMp7DqkyGFgho2AkorVEImuaQtMZD
p45yXPCqo6kJhkM4EjZsH26/BgTd93GZyactJRoNQ6JY1X7t33esoyvQosTy
ghjtwwZM1gJzRkIyuExhL5fgEMCsuwgZF+S1tDOZzz49e134y5GRIH0ljMgY
myBAypXaTudfnHFejXV/EFhdoLR2qxTRxZygjpZO8BR+MFTPsYw4dOeUrelK
+/5V3clBGrRjFX8icAaAcec8Sh/ZyZ9Kf72j1ANzYqqhpSbzOUu13bVB1gMH
k7lZ3Vgo7daTpVtXVHuA4XyjNTV0y1GFTZ8ecEMsuzIfzgJEeJTr2XUnE9ML
nXLvODcA5C1aZxwFf5chP+HUJB6aAtSeL1jh0AuYiBszwIh5pRGz5icV5/am
tCCF8WXf6vTQzFvsVVoRfJ0FPxYEYZP/PPjggEI8k0T3LmLeR4NmywHJcL9F
VZAtCSeLpWJL6Nfg87Y7D4tdH7ddxXp6swWpyVGWH4fBQeZAOW3IaOX9n2ZO
/7Kmk35bgozKSIVbYsc/msgwnjRvhRvfEbu6Xswz1x88MrN3DaBYrO3kS6DB
j+quqhVhywYIZIRpgnaJCQ7MyHEOKLXnu+EFK2TSzayrIGhBjTp+qLUgXadY
fcqJcAMV0HvFim9Mlgw0I5/KHM54KbWqcy3TSA1ccrYkEQySkGaiwU/lOJAd
V+NYeoAURUg6lV0lfCpIgIGOxnEjUKG69piR4DyWSI/+SMk8tTp5a4E1Ijsi
nSKBrZ9HvnxY0xx5ABno7herNRvYVgbpgmSQg7WSAvujKdMuWRIcc+/5V/TN
wkxHMdnuN7bHjzoYrsiZSEMmfOzabFfoOOTjIcdkikmvPCHmD1xG9uaCC9HD
OU1+IVcmnIvi321apgOwbyOB77hncK8ffs9iAY2NEsZrLYIKqz30mNQxh3hL
aPc4+DVYElir87MYNJldCYa7sganJMW+pL4wgvNidnCdzUvVFhFTvaMPY2LI
FJ1tyscl1HJBsSFYjZ0+aJV+87HgxB+rLeAH+7gqlgVMYJpIEumXcO5CmQtc
tpvFqr6s7GcJmQMeIbzmncmuRh2ijwnFA7HTf0I3IDxQWqN4A7h0nYjYIH4g
3NEXh8Y2w5WN9haXcKXdKc55XeloJHchv3GdlRZ4Xg7AZjEKksNVjS2NSyyS
A0R21Tgcd0QcBsXMtvpNWRTDxVAASaXXJDsm9dZGcywUfxvQYGFd4dSZsz2O
1om79USFE3FUIwyhqgEJsZ7eSAnrvuqcXBGNMuyuHg2tMf0bV1WKmTpM0TGo
Rfs2yOyqiqnQN+uv18fA2NQbcFYwKG0SISpG4D2K0LlpvhnD2hQS3pX5A610
bbUTHuvkxWcfOLvUzUnfWwnmJ3Yccdg1g9Plxbxc/tNo3ulq3Um6UvtfjLxW
Ec9LtihZRiyE/RDdVMW7DBo2OMOhv5k16382ZCrBKts4QG8M24i9IqqMxkGv
9f9f31YLNaNV4rDFe2yWKedAxGg/Cbuaaj42o8OFXsaDFWM+WPXKMn7f9vkV
704hItN+LtBKKHVItFravIFLHTYDPnR8WUNPPkgcnKfHmje/hnr6RNrDDm7P
OIdpWn2V/fw951fCstdV4jNC12JdB2k6NqP+JV2hCi+DXAWpSOF2OuHo1VF6
rCSJ54Zg8I4id4k7Sn8M6V9MEOe1kn19ZvPyCzL338KYBjtFGu2fG4V934Qm
mfatBl9z3XoN9jsmRCMy/+Mr8UMkO5c1sigkKeXUhgxse67AKSc2jipXN2FW
F5VHpkY1vQMa5hJoN2fSKT8wmxxKA5q6ALWuiH1RaEqvXmiZnpdD/Jq7zrGL
oEUUym7c5HwEMGGgHlNbss8ApLoTELsGPEkGwcLF6IrAnBL4HLaFCDP+0M0O
tz3mmuDELOU00wo4Sww3NPelwQeNzzskV5fyuhK8XpNmAW+dgvDGQzOrRDoF
+zbGop9OmBoivmexLx5nsCztoOm9PcOm74X+oJSSFwPjweZ8IiFlvIjMBh2J
ouhZP1VE+8qeYfy3Jh8v0RHCGx0OBhetVcqojKW66N9camSp6ajubc8wtEjq
QXunn9f/MKPRG3lQ5oxjCSF+K2OtfiqRq8WCB6c2uLvrTGDm/p05okQdd3ye
7JS76f8SVBSGuMLJN10zVWjTU60iaJPbYupn2XYLIU42n5xqybObdYI9i9rW
tVWZRb+pkWbuYNUdi0qg64mNItplkIJ+nXlijNV8CQsfgsLuK6YVPBeHiaSG
KyY2QA0jRVt0f+/kDX+rc9WhF3p1ZHntOnLfLiO1jPHWSbZMQqr87dXi2sg3
/GvL+ADrWEQ+KI7r+SrkLaNFAddclHeVRZKjLhGraUmw1fVXWTHQz30tCeYU
VkT9oH+R2c1ywXu96NEdWJUlQ8ffgkdU+sBUKKdiKULZM9e8IuWC5il3fwWV
60cfEx24QhY+qgBBapit6b0qaqIhMaAlAlsy3pluU9t6rtdl0YfZxpk77muD
LC9yJQTxagLiHTpm4fIf3LLBMOVEjvSf1YPFtzf9hssbnyMZQLRjFPvw1rI5
jcUrwyvaJodDhjKwAuLBAvubwd9OcnwUyYewR8+mCEAgEo56qTgCaAZVHtO3
NUocDeQ+12ST6CfqXnX9byFJByVeHOtncBADSFXDVch1U3mmmagZkzV2+R/h
V6jsajsOba07QYcipYEpfKABByMeQPh/PdBumIcDVJ6znA7EIpwgjpH6zezY
WiQB5q2amtJrfeVZQgWTl+/FahTgmysrM/r8uVFpGUeBfbxvuw40vOdfRD31
gx0qgLt4/U5IQjKpPqlN2I+RI70KQSnVtBPXPIztDIZnQl9YmY+wmXf6d6xR
i+bGUhHEBcPXlRbmWSaStwGDLmfKHFIxQKLoNulcCkfs6KTuj2GaqL/3D/0u
0QGBNWLU2fWv5lknLwcYuzCVWoGCA8lM+b3+XLhDEC8/KpFHr55b/SQyOtH6
QJEzzykLZEwp2irYIvvR2IV0jBe+BzmvVke26V8lt9kk0nwUGwxmT7agsXfj
CSYqB7E30ojl07X6ABS8YeRFghxsJJZqi4NCxE3Pbytk6JfTonkG4YZFw4GM
69Kl7PL3ZamIAj8fG872NGHNIruODKtYRTbL82BPGXySfBMisNoejAbhi73b
j43MqH5AvX4ZYUnItLEyuuuwoPMF7qL82Rjh9qXri2/pOSY1MTzwz1SAVAQW
IVTYBMmdNZiG02SetURrEIV4VcqK7DORj0s5WbWZIIY82YTAEwh3TFVk6lHZ
Ir5Xk4G8ombLDBopLpSHv5ZAD85daRdfmSh5WFIfSiem488cpAurTomBI9Ju
yCI9ZlXPpgwToGRIpDIUh/Uoz1i/VgkuWrfKscKTG2hTUFUTsl9PX0J9il3V
dRByv9Mkv+T8QEvJ3HPy7k8d2btCoFfLR7cIyZzBLs0wMFsUcBxN4ztLJzi9
R0gUkkGP58oSt0gBfqrwHVFHeHFiN3o8g81c+y/fGZ21zSf2MRidf4pPO44w
64f71w4UEKLVaZ8eZ1SRJCn7N53kUTWoOJFv1zeiLhP3VEb85j64b9LYZqAH
+wwcGgNK5oNO5janrQYAhUWzPs6Bx8215wgT+qokfLHOW227iPbFXbPPvrr/
Nr9idcbnllaXOaz8QGGLCav18cUpM4yQ3Ss/h2mXZkPifwl5HDFFQTq5lGwh
1ErtXLxqjayOyy5tgpvXKjlcHy3egmLMgXPUV5lQrHoAhlf9QQ2ox03F5lAM
P/FD65jke8qSGs09xvBPpNCBYBcbVvN7oVBz7sUxRPh9Ibf/Ia5yxN/umCub
7RfXv+LEXTmgFnvZorWbuTsoHrZYGS579CDHfCyyV4vbSnnxSWNjo2+xipbW
XCIXf6Ubdhj7CZSUqIfv1hdsC4xFt3K3bOeiT+yUoDA5xj1M6dGE2vqBU7ng
WnZX8HWe1Ts86EhwiQGqKfVT3xOwMYT4yKCGyI+AwZBEleeDIp5IkJqtMVpv
15xQ/KnatmLLc7TdcePF40xhFcHAYYx96Th8EloHK6pyMPu/5rlDhelk0YR3
bm+wXO+NLa0ZOu0pjLUN+/Sms0oq6MQYikIS80Jto+ydAk3MUSSyks1PLD50
UTfE2owqXORopWczJ7mR5ZN2VjzA32WMIVdWKalUZ7Mq6gYX8vl0roCO+y++
36hUjSIO2wrPs5aCVn1YB5Takd12UcFlXQdLRoR0MgyC+HOgA/kybnTq19Nt
AhNP/Zb1T8GOW/k3LC0uk/9oz3/3lVZ3ZlkUqLk9UhpUOqaTiHUvMe3Cvd7x
Oo6mjBY0X3I5IwXcIoz7jBoOj1so4y2EWOVk5Skz7n68JwtZ1/n8jwdXxz4+
8kcdNYiW9LsKkdMeduVULOxhHmDFsjGcSXpwRRfcL5b9dPouDki8D26TCTTO
0K7fSg75nj4m0okI55ZfVoMrwXbNk677xrbmPRHOJznJdwXyuHLUIbXjHH2B
WiaArehh+vzmQSRHXWx9TL71eBPSRsujZSCxGLGS7SgwalURrxJ/DEU04LzP
kwpDNzRx407Ob+JoApcStgY0ymuYrvXvYahZU6fDisRM/rUbGpoa9KoqLtyI
iYFO7rJiZBQn5mdKufZlilCSXu1PkqcxCUK9fFG/X1ymHUiF9l4AWqP7mhCo
8lNqK/x27ybswApOuiHqNG7iIENKLInVEYkjxoawifWUEQQU3ugO/FRk5qT5
TwOFwFbbXlPbJ5PCztLLEmmASq45pCHqZf6Jx+NWmVmGuZBMvB3Z6vni1EPh
AsHNrEIfphLr7kiK4UDtc1s7uqGfql+piPcYX1inBKK/8yRquwivtNhdmh/5
9Torlg/WUFHFUyT559Z/HJkRbyVofxsI/wRvplbCS/sEe5todG4rNlcwjDuX
U6U+dAN/SViStomObOcvCpMv+OpXdfyqGXKsSNxMGQwhLEj9oJriPNhaxpAx
a4Uv0tY0lGR13nYsONfR04rN16NU3q7Y/6Zvfe8NtoarHWrqu3wJENd2EyIg
q56XlP2V6/lwnt6TRCh2P/7XK96KDf5QZpqztv4k2VLnBj6WXMfjJMZKT960
9kDMy/xm7ZdrJhGdLZE0kKwSFxdvGFvFerT4ZDkn93vCOL3qLUDtcAsdmCuF
ZN3j35oF+d34o+llWkVRMUux4koqHHt6ydB82I/9i/1xNNaG0wEm3zguRlCT
8NgnWQnDOIp0Nkkf4hf0HfDIP69wtmCdxZs1BgJb0mSwNfielaeLoLkB2PdX
FLe/9/DgggcOtrlRTB0hYKTPEl58CJmZeCVzsdC/y4cuNafTAFOyp3Y8hlwT
w7ytNAoZ0RtpN3neNKWODPXxtsZvsUmNZBOloV0ftueJt8ijFAXZAWMMJRsC
JZoKYnvGArbCAYaDhNF4t1+H0jnz8vgni1zr4+AZG6vpbK7AKv+YxXu7CvE3
i0OGhVWEdn5AsVAsKiHfk6q6rw+TphZ0GatGurxi7Wx5yAvl+7g0Ys8HyDwW
OCuo8bk4cR0nE9+l9baK+DINJIaUDWfIVkqEHfMBJ5umPR2pFRDAprcLEo6F
bdP8Qpyq7U07TmEcLgDaSQNj9s61Q7He6ZyAS2sAKtTN5CG/2HhVBCV4uM/l
5h625vGVkepLo7jz7f0ulnUYOUylj9hECFrku37WzLTlDJZa0C6j8abo/Tk2
YQSJgOezWJdyd/om/5pINkRJRbhknKVJgck6jSq3TinVe+84cchleYmmcYsS
qnbW9tEYzkDjXcnMSsB5VDply63KmeR0Ycbt688wgR/7cPSrH42MoPoGmbQn
CkH5zjBb8HM+ZJleqIexgLyRXF+WebdjkO/LZR4o1mPAPm64Svy8CrY8r+5w
Bh+MkMnCRkzdKw0CSuL+E0Sji6ZBQThHlqD8D+hg59lRGHADKFB2GbOfO/rv
CYGJDpRUs1PamcL76PqV/RhBxxVWx2uRvtxcOz8T7aZesp7aK4qIv3BBjKaF
b/JSEwB76Ql9IPaRhqK20oLXnp4rRs+HyQwmWhFJyCDPikQvIe5a5H8VfaZs
KUiO/JWa486ZHy7oXCx01emtS0V9Vmvy/mMPL1U474piSBjOJcoPxFWXL9P1
4VjDJeZD2xX/Z1akz3I0MoUHbtH2h4YJ+Qv1RBfmz1dRcHsMlnTAcH3YVAR/
26tht1yytvQC79qz7VutXKg1vphPV68Ha5jIT5JYxyHLb5NVZ1+/03lLpSE7
q31HMPAaduEsCkho7DfSqZUvvcy0hl9Fv32BWv/szGqDnfytzTkwP7zuLq1D
+ncfGDz3D1/zobVC7KHzgrS4oZcW516R6S6vzLUYUpX0KQO88lruuFgLlTUz
h3Dgjm/l/Nf1dwG1xSRzZfMS2tcqtqZWnVV5gCuEi2fWQ2Zo+H/EMGD8V+PX
EHkOkpiAiJpHkdqszAj2v0v86P3e4E9J2tTeN3+b11pfxAc2oRjTLBFWIRn4
o3+CEyhRspPrTNj+r3SJHpzgGz67962QpAKBrPO77ZLi8XhxAWOZbNmbonjl
/jf/gKUyoNUwSgYt6paFume62PFrP5e5DrutBkMKxT+qCORjZ3+tfGEF60o7
oisZ0cJ5BkdASV6hO2+JTZqk9qmnEh41u7Bd8GrfcHTTT7dNJhO9/ONUmY4x
h1z7my4ZFid/p3LbBlzPtA2wNjWVtXDaLqw6NGInZ8Unf3ifpKNcBvusx4DD
mgqHaITxt+Ma63S0ZQnuA9Vu0+tLhxWYesi7hBgMaui96Tye5+PUl2tGEUV6
FNXPuufApQkjNj5vnH/YCriUSiC4QP/3GKzvn49Ey74VLvcg+OImK+e9wSjd
xgjCCyJpXq5PGhdRADxtVktYsBgSsb9FuvPwbjoFhtvEgbT4w24jcHXtbSsg
45Zpy5rs7rqh0AwYVQWcxfwDrtmUIEutf5eaT/4XGKwWjyCNo76O8YgMLBH/
0RGqeGOcb04kYmvC2fsFkzAbHPkU2rSr+fU7zJ/05Er7R8zLgsf/vzYo16v8
+bQ7tWTGD3xB6B/kB02fH07Bb7azkjcScpxLsraDdAv5XkA1XAgEnROGuRP/
5TohFWakwqJfcqjwMgXcGQCHBDVIHE9UcfR/tCPpw7PDYGy6zcfXYYzaYVnh
eEc1ZlU+baMSnZ/z+CcVuy2ZzkJwxup/xxRjvhfY2nwzCSI/ygHmXEvBJyrk
MoOLQsW0E0Vy8+9OuY5c43NNkqfqrE1nbN8aopxZltCRfCe5aGJPWx9bygqi
B7kEyiu/c7w8c9vpH2pqC1q0G0jDhj/4XqSd4u9NAAxWWi3y38JxlG10I1gp
n7cL9Ngoni7Br4ar9QjqhB/k9nf1d88hsUZ11VC9zermcZNdn+0d7iiOwARX
40L1YYAZEB99DvFr8nfSIrHmvddPd7P+mQhGqfdFl9Z+90T6O+NVRZaWcUlI
gv1dgM9JAoI1V3XnaYK2EEJV0TTCBnfYXfaHd6g3RkRLyraYBthkVXqmno7A
KR9XYqzFH2or13wjshZGUf4SH7Dv97tGgIOnKgj80lye7zqveKj8tyPQs1GH
AnDewI8Vmyv0Rnzlr4yEN3ywHzXx/Okw2Vt06Yw3jge7/aZwmZu3sF06jPLC
spS/Wk/cZ+s7tfQJcq3+8s/dReja+347D6JrpDu4+KNHR5tKi0nxUsrXWFEi
ku8+UbyRDtQHXUyWYqxMtgJYJkB3SxS7Hg+pPgTD7L+co48ENIB1Em26iuo0
pCoezgpzbb6Blff9ZwHrMEYOjXvdRS1PmEw711YXzPYP+YCCkQ50yvRaDais
tAp74XmJrmCeqwAsSjjzJDpktcs28aRTVsDFREQ9742Ww3jeWvVQ1w6XQWWf
YzDKYB0NDtPZMlAOJHCZ38RL2adeiHyYLn1mNiQruBMY+IbZrplldAgRc9rQ
e3UyR1wR6Z+YaOjDT1j3NGtqq/wE8tjS6RAb8BSIrzE+oEkm/WgsFIyfZ1dE
bt/eyV82yI4yzs/jYQCld+/wpRH/BQke3HJ54wgwfHei1x0mlQUiUIP6lc3z
eJkc7WhJwyU/9UIazDnqJ/gRysMu8Fawe9g/tg2Blb++gP2WFMhhGN5sCT4O
gbiCIBwb42TfXBokuhpbwa3bSXQJfKMeOVMsjIC6bktI7ub6iulROIV9ZqHK
pprtChFgCjfzC0VrnnUkSVc31giwid/DHYMEVUUO6BDRnLB7P9/0xj6Jmim4
vn8p5h7flHfEd0Ha+/0da0Zl+qn82Fxtc1kXgk8hux8UgUhAGWDOBInrdoT+
2FH88Vb6lz2MoVmY96QAoalZwCpm8UoLw6mVtoHC4V0oPG/O7GWI3CfIjjss
6vqgK8xKysEVFwy0yI7Oo7R1DJirekyuqJVInUJ9+tZkp53nWXlUdHrHdg1j
jFMWYv10cwS2gYATEk26TmgzuqmO0+zi+LSOMYJBVJkLtmLYR5BacUe68CkK
xJgAB5rf9pTAM5w5B2z9JnH4ScYYsG68KlTfH8dWqwNSwn542JngcwDQJekh
ND1sm2mgBnfQ3Gi6AcbbKrwizf0ewC3MCqBoRTXpw5wTNEdpZoZyQsxH/DT3
3Mi6GxdkVsU3NiFlALO86a4paMveXAHOXWfsfihqiYppp/GVC/8EXRN2tNut
XEz3ZkD744xiaRC51Zy7duMZiOdMahYr1nLxsCzs5rXt0+aQTyFx77HvniXH
FMEvamKqeFeYs6S78tnhZtYoYMmi/Wqatv3LMR2czcNnghoQrGmwJuN2xnlA
g1N3bRwfqcAAt2bOZ5WqwZpMv6OE13guKZfjPKy8uWqkuQ9NJ0UFVV8cEeKn
TsfnyRJ4hcrGZSEIAfpVv4TNnI5cGGTgYdgiahE9SWkb6DPXZ5iLtusb0JXO
AHsCqBzyuKE12N8WCK9WvvRrs01fEJ8R8k0EX4cXTtV7WhFiblrqV3brH9hT
OhIcTeg9jrkgalP6+6/bnIk5/lEMxjXjmEhXRa+IeNJwNo/phfFmYhvUAqwR
dbTElIBhquhl8MBeDx5VEpCw3x8M3SYhmSCcanmidz7OGoxjpwMGAj2ADUKW
6gESvOGm07UzqyB5JsOCoEAqQYh2C0rRcaseRDWbKxEn/S1zBhA6WjbzuqiC
OWpFfcsw1ns3EnFeKhnUiOjqIOCV2fo/iHt2HBmM4mXbLJzlk+PIg3UnZ92U
y2JEGai0xi06oQkjHx5oLMLxb293LeQeD3An4893TT9ycTEs3fR/dR4ieK4p
iXR4aEyJff6ZDIwc2UnfQzo19nAwc+cbiuIo45rkLByMgihOHHTV/gdKjgnZ
cJwFBf6+2GFqmMX1jSOzbotFa4gh3LhMyWeQr5LuBivM2SblGp7NP6JoTa5G
5q6hEe3bbSn/36CGP5mO+hYgvSzkK4d1VPGVcnhbd7wSG09Ay8Wk2aUZKuaF
S33EBnrjV+MU5oW4sz3pNBK1yb0ifkj3qBSzGRR+brS4H41ZnDJuhocpTRoL
NWofJ4ps/qe9bA05G41n5bmnIWrGVG9w1Tyz0M2iDfdiywFyoUHvIIM20YQl
qMWlWEFcO6CMYHMm3myBGFVmaeJawGLswNhazoeUyWMpinjyW1HQ/orGgnfi
P5y6qnFq6OVSPkMtWhuDGEDdW4Hq4bHnKTNRsNGimCcJNjvzqxcQHVK60Lkp
0LhJd+0YcuAIzXBmucOKj4Paj/UylB1Xoq+ABjgW+kKxB/m+6pooU1Em5X/3
qK5I9dwIPvICC96eb973hOhtkb0mpXBcMVUcKHrOAF+Dsch7mWmh/A3964Hu
UpdGIxJ8cWLPaKgJBi6Bdh+U0xQjEVCqox08jYWsWqehV2qBlAoCvGWQBWJb
EhhBKxIexez6Mg0KCj7R2BOdpRfYZhvDLh/v6b4m69eFvso+UM8PAAqmrgRn
k/Nl8nqgZX6Kv4+jr9g9uuexAr6pvWPSyxm3k/C+LBrNfbLAbwPpzYnjMSNv
2JQuja9OVDo+jB5GRs+DOmB6caEC5KPOumeDyVB4uMAZAEd7ffRKf6lXC4U5
3v8GUfoertTFDdQ+R2g/igI71pKBHq8r8NI6aGUeMczaDGDu3MgMD1GCE6Gx
HZkVG/ULw8s7JQAAP0ByvDh8m3WYmE5V17WedbW0ZJ9GbGbTURBIYC4D2C6o
L5AXpOAi3bhRanwwIgCxUh+poCY/lHXFs/wtFPjcBFw/kxbPT0yOtj8z4Zqj
J2IqTzjYEJZ0fSM8HUT+EW7cB77D+Zn5nfy4VgiyhdqTf0/pDtDN/+wFwkZq
SMQd2RL2XiEneA+ceXE7eBZgJdDyWoJ4qYosCJkGCu0gsHHi2ZkwAuhiH6g7
239ALWmvAZ2lVLya+XzfwbFs0e3iXKueB2KdHUbMAel/24aq8nTaSzunySW1
ft7UOoGqbOiwiqFBG81+b8Xb1k+GQbQ5rfHldaLgNX350DVevkJC2XMqqQBL
dyFzowEvEtao5OZxkf5QoahTliyY3w5ZHGHCfYMrbb/qwq7arwwXK253YMAt
IhoWxG0V5OG9Jx/3f1f4Kslyk+/PwqTTot8QSbZhQLMLVBbHOjP6JtYd2kXY
BHJ/JrxALzckTaMdSREhZIt+Witg0aeDeN5pvOD30gOL0rS8qsfKGTZxtUb7
7d5LbEF1WUy5nATLLQM0E0hdrlRYzcHInMCgzXUAUF3RdHgkW2XC3jxgxUju
577HlTXq2ghICXTLAH5yoqc+6GklBrL8/yZtPJlSVRi0UH7NXHjTf8gE39Ja
yBtQqcITFSFzrbCsaIgo7JlMcQ/ojBXHsds9QKESt9SNqNZd+86BBRF8VFso
VJagSBw1gbxMC7AhJsZ98Y8UbDJH8kZO5WFuAG/hlyZ0nYe5ZFUrR2B1Lyvx
6ez478dbVvsQazWEY+rhG4PSkh/LOu+eXb56zJLFlgYmh6fqm1fe+x1kPPwN
qvRz1yKe72rlohZnT8oe8QdXkj94+a2kWgXrEUHMQ2sGCndrlLDLMeprXozw
z5Wy/n/pOwlOngnEBKb/+4vtdioYcloURoSiZjJdM1oihHYgxkp6cqnDEM1O
zsxhhdi6+il+jiNK/9RCMy9if1L+ldNtlqOJrJLqf8fYJAk1aSh3CqAAD9FH
g8fVTClgUwT8NYsDMfHRSQnfIeDemZrZ4/te80au42rblAWHRRYR0QayN1dS
TsOnZB0O8mdCyh9V64DmR+lTE9KLJLeXO4cokRbWvXPknjhIIoTOVqg9r4KQ
EBitSAmL2T38vkiBDsZ/bGHr6u2ph5VGRbv/2MeW9eMq23CSsxSBkYuI/tMV
lXipEvhaiFAYy4uKXxyElBajzoGYEhy6HeVYEm5gbmzkwP7BhgBar2ByZu8G
rsWiCrnkLE0uZ34UvB9XbwTIvV0wkCKdDPCLKkoZJNhIP3x9EsOuL4Ant61o
usS6KqbktmGuF2VMj2gju7JHeM7TjwvU9CgOLaJMLej88VUZNf3UBPQ2GRIS
hMI3fgkTqa2BpJ1EqIGJI4N9zOXKhYiiNEFSlx0GyGUTTVztIVl3ltQLsafu
rf0E02STRhcfmAnB0/w5+mhrpO9GRtU/cydXZ08X5c9IBJDBM2HU5Q6G+wwO
CDOU2nNDW9MppnFpi0//le3Q8zVyRJzEQ+nv1MbFumhTjVa/5m+1nXD+uUbe
GvLOrt/6dBD4RqSIoYx/TkvEMtpANvr6u/kUx54LoRMAnaSM22iXgRYVco3R
x6Ee72/7oTdjZnGZG9l5fzl6VAf2MNytQsdDcviTnIKVogxQxlFchoijwkwn
c3gK/jD1t/WXwgKrQUxXSyjYt4YNQ0MSQPyedmSzPpPZp+g/4gm3eLoHv/lZ
2PTWO3TsFb0ErhctcrIahan14x0deKakQaNc9Aq5iBcz4MjfMKQvo4mhhMsa
rMqQQ1zetEPDjCFVEtTR1PLjg5TmOcF0AcpHieiJ3LfYU05n0JrA014arEca
4O2NN6aDRbvYx/HDI9wtoK2KIBnGGy7oWpqVsgpFWEpFfXZpTfKBL0bqcM0/
44LxC6mvC+7KxKo6P3vP7utbl+GuL28P4eiTFdrFlDsZZHMt3q89l/Na+M3G
gy/SsSMAtv5/rjGO0iy7k6osI3qax3vG3V7lwsfZ1/G3x+lr0aAo9kLm01F3
8dGGKS9mlabtmOd+VVPyfbWqgQkDaP62hZh+boAUwhgvnmNgmFArBPH7yU6S
GOfr/foUl6ZpQgj3tUNwXLwBVSnBLyMEdPBTdMNNP2TbMofcmW9xrEpe+2sg
REIXRC1Bb2H3eqSgJQV0FueKOk8dKzol/3tzFAIjQXq4R009LeQa1uQ4pUUP
J7zizZlC+R9xLtU2n3N7K4O7jxfs1fniKoU3YZ+5t+3YOfxAuuAbSdYXkpZW
ZESiORpDIqAbaCLngD7CNHv88psxe/sTDziNM0PAfJgjWCj7qt+nB0r8xY2y
7nZeGnbCu15t9ypGQRg/RCdwdV2VKU9hgTjG7KNwrKbuFZ350UOaMFoaRdRY
LkASLOlMMjuUn16+8++6il+qJcXdyxTxw0J5xtg4ijT8terlK79M3EIqI41u
Y7PFO8ccS/UBK3wUN6J+uTpD5YVaNUW/3vCcfKZ3OE/MxmymgMV+htayOFUU
dFe9ymctRmkJdgYDAOWVRmz+5aDQ8uswW+OWxUstOZhwO3U8UowSgingdm0V
7RvaYB4jbeAgnGQBk9qYzcou/SFpiFduZkMdknTgVR+NMAB4wOI8l8CtNPS6
vLUehD1B1yMOHf782Bc3+Q7cHK+YvkvyvMnOX70pZgdWUYv0TnAmyOIpyAx+
RofW1lxuHeuiiL0VYs4KF8ZwJrMh/Fc8yWEzwzbL1OX0MJC4Fn6KgWBMARuZ
+ZZkv29cmTBkNIcwQ6M1OiQC34I2v0NJXM4rDbTFzy+DJPk01LJ4Avnl6FMA
jRqHbBfab1mQX6Sm6O/q/C/RZBkHW1LOZ4OgByOmNk5kqXGscpy5j58KO81m
+T10+YTZtXn715Nsa5fmNE/FHxrTT+Zy4hv9kXytt2ueEfAHtY/sGY+r3d7R
uA73zswxRk9x++g2sjGOzOppEmKZbTnbefBXRmt+6O4sx4Q+7g392u/2yg3d
DtrqaAH1OxavVUkpvDX+zmKYcFq0Di+MZqFS575sgoxO2tUXTi+5N4HCURMk
e5YghrIBdKG0DYHY0IU5Xy0vmF09tU+5BVw8f5FP06g6ojQia+lRJsRDBDMw
rgQxkXix83X2GEr2cRztJXbCASHcuAwnPo2EJ5m94ohWSSof0/7BBizVaZbu
xAjIuY+0m+ruhQW7zEN+cJbZHIP8LVbl1OKVN29kNQaDfMCvN5WN2bPts527
/j8skgtu/t0mhD6f2U2yjKsew5QIsoR4dGyu6rmlVA8Ffx+8CxKjBHvjV5ow
HVkYVZei+MYEPkRHrObC8UhVMTQ52UYsma1aOqgJRsrCDY8SX5/JQl3Kh8GB
duW32tL2M4ysH9f7jvjBygtWI+cU+H8VCx2aAFSdG/PsLl4HwEf7jdBIzUrd
224V74lkS4mW5cdSIJqeSp5bdXjdSJJBcQiRsVowSsMsxvxUQap/kAHcEn+i
9lUAkUVhvrJ7heYR02leHVWhFAY/1cwDvSouJ6ymTkhiwzL4R3waEZEKJyGT
Z4IigL8XMf1nMKd/2zcpmWHIGC3UhcAWE41E2OBesnDfeDEH6UTsKwCrNkhp
tZwkzaqh46MCsnqrNIFo9OEWXuw/hcKKH245OdJJ/Su3FBAjCuJtsHQIW+me
I7V8z8e8tRlY8tAtuxB2VWYcBr4+cSdrZgeBt+qsgoehceXLYXFiuX2Uwwr+
ZXGXGiltQv3lA26dsYO/GqQzladggW0w7Fq77V/JZ8sIsetJSyrC94dofeFc
vQBike8VtNDFX8ThbQL0PgLSPyFF85WWTV3VWw0GMPzKygp1KWjTQFK3l4FA
R9e8MEBupmChe2sUabYxtBN45EgsZvo2eKsjik8EWzO1yn109qeJN17H10RN
bJ2qnlVeQx+vZricD0OoQt6GNNNQh0lLcNTgXlPEE/QRsvJUyaio0VTzFSzg
z/qhjmabnXuvMqx2+J/JmTM+Emwntfce+YtyFTfesrReM+c5QbKruUXHxdZy
JRyOswRez5TA2Th6AB8Ciit4L62q0itIsGpnTbq2FHsTLFrunw+nd2iWjrK9
JESGTebj/na1YAVbOnI04zd01mm1bP1w9y8jPvY/ur5y/g9AAqfzk+aeeJYl
ESsQkTPjJOSy1fbz9O2XGI7XGTAaBAFuGvJBvmyaDuBIK12HbfG9iLXTC0E5
EwyG+47kU9559+QXkvvvehX2dHEwbPS7cVkgQ7yqwFwGA2Mz9RP+DrT2S0aL
h4P4VNNdT+OBdt1YrkBkjWL8k412e4oIrrNI2sdECkLT7UThn1R1zrA3iwxH
tcYhSH/OwCd15mJA3ETZEoQqfEw4k2Jw0epe3/R64lsP5R5Dwwcq3QdhjbEs
xEH21956sNvkkF4RSTq6FbxtdNFsEXZQIEbD+cno/g4NP8jdfr8ikDSreHyq
yQMu+ByNF3A9THIggna6UcLQpypQz1xqCspnKRrXh6PKnMg0fD9uba9hf26F
M77Tiy61cgNZIbcSDVKc0lGg34tvJWUgrz2lNZGePsFhI6W+65Gd8IlktToZ
5bgcuhM+vE7+aSFCdP8tlX/Lg9cGsOFk4RzmkyShp6TB2nn6HlYmAgL0CM+k
pw5F8PK3pBl+Q7iFH52cIb4o4b/ZI/fFHYBj/VkymoX2mKISzMc2uki18+KT
KcjKWHCOUKQA9mbMcYc9dD7yAKnOHzDMZdc53Qf5apu7IPtWKXGr0b6EsVgf
mOH3ijJWovRFSDbM/th4ha1c5mmbG+Tf2IprotEbgeucoToLqN4ky7rsRDen
J8JdOL+odbjTgirxqKErp/hKtQ2B89GOi8im8DVkUrkxUIQmT/2hY9k51lwC
vsqIDGsbYz3M/eg9P4HmutMzfBdzD0YYgPBViE1TCi+r6IDNAHj7PkKXARKj
UthXsjdwOYMBEt8fPhg8uMb5Wf50t6GhD3klG+a1KyNvD72+pkhESxcyruBI
I0ASvoqSVpXaLTQh9F4VzWXwCPeVmfzl0n8xbuMefmNua56X4cd1BTM4mX+v
kcWYShXWJ7GYHQLy6FULCVybMySdVRtzGfNX3uZQBRhrpfZt7hvos0e3vaH9
Gl3tf7xeAIBWaaaVhasgHmvwCrRL/qkYrSlYpqnTdKRoZGvxQl4H4S6aHnGZ
wY1/noxmClgBZ35wQaY6knglbq/Y4nDDOQf1rZZAg57CX+fIPJplf0LG+4CK
7pUSskyUPye4agZZN5lEjmYPiSeOWr1kSlO25MhM3Wmrka3wb4PBlW8MMnXB
J/UtKOhgN25VrRVo0Y+Ha5UZ2fkRDNwab65Ju4U+dUyjh6CI/i1NSt2gm+wC
RvoLCB/17C+30OEoZlydwwBHju0hxnUvQWhvdB/LIf4KsBC5XtWnInlguByZ
cI2R1c0qQRKDZ8ZHhTokzq/B/SsanxDPBdoWoaXtgVuxHVR7125WUW4S1D0y
1bkh2T1GiRq4TsOHvVOqHko71UQP4Idq7jzOBfhVjq5YqRg0XOVsN78D+b30
PibOVxTLuzs0QnByrkBjRdIaMNaKal4u9EPSMvLABtcAmtQQpomsLscY/gOV
/d50DiS3dWItEmHeJCYsnBW+mlK/Pxz/XmBtBRPIfgfLTMpIhnc0bb3pboT0
rlwCO8Tfq/Ep9HigdLRW9kX2GIyk22hzv0Nr+OCHjp3x3qYgwGuHP6GjEcb6
EPbXlA+trwcXGuT+81p/hmphv5a7W8TCRnk2OOsQ7IQDQJXrgHmmHkW/EntK
3Oz5qJlALTQBcIAj34b46I/yia7iT2TS8b/ruAVfH6V+tF1FBdp0joDNkaHa
aWNV1gEwcTub7dSAsn47v1oWMGwDwNUnVgK3WeA3N8rsGhXG6C3IGix7jfcS
MVsZ7xa/tyA3mpluUe+eS90WetLmk31bqOALA3oi3njbm06UiUsjTPyFg6WO
LZOO9YJr4Gte7epOV45+vQQgsGkwYGzJ9ZWZyYQ2WxE3B+3PC9Qr+lJkohPk
Sh1fIIvthUzSwNnWZVI0R1IQAY6l9LhfCX2HocfMjb2vVt7/r7fSt66kYIW+
jWhU8o+CnZhS7tpux2+yhBaz0jCdx4HuQxz+J9M991qOzeRlxSLBBVTY41YQ
O7vL8dWuKNHO5KJFbITCIf4JPNwVjY7i0pa1JvZFyFfjlQFNB8/bSTYZIVD1
2Rz5fBAx+wKBrdvd066OGO4zF7FTe2eZTrXtVe0kWnwUi3EFE7ZKdRTapX0c
/N1bjuWoav9jXDlN3YM2gPhO8MbrS3sWlJfXsmzVwYgOs61Xc1zOz7qw8N/i
fBSZH3sGcVK+niVB5bR0QGjJNwruQg388PtNrQjNPYDFQFi2N7/WQb9YlgHt
Xcx7rZ+7T3ucCVSNkLJSOlpnCRhjBbkLALeOcf9GrIRO3HJ9kVo18i4453qm
7oT98TOGcSjrP4z8IGzKfltwu9+ihrd8Ob8EvxqB/9Ahs0xJuGOuXF7G8h2A
YYpED1Y0EF68dKrMNjuOpSDobR9tvvdZhMoTFZEDXMtZaX3drHqY9JHSiO25
QwhFoZUtPhE6IpWK629a5B/fVs4s93ZwDs3A0AqZEE5rKCgLw+o5r5PSyvZD
wiNTXavTFT2cjUdVIq2qBnYGu9/9WWUsD7YLj7FjV1bNtCZ9VsjaOJ7MQxAz
L0E1UQeNH26LmLPVf3z2A6pyHKqFdyHBTq750KIYVvKFz0TIZU4Pvv5LCo4C
BnaO0/we+BLFLdc2Psm9UXHJR869r3TGySt6tMofcsYU6giY5cGl5F0oNVmy
ay52svagdOMjgCd47TFq4xGnRzkk99AokFKy0nSPTYyERpEAxD5bhXtf3YRk
6GnLLdYNwSA8MY9i/AyPqLHJt7fQKlmaP0JqNEyWRxwjsW2Nsvhng7wpMdQY
4xgoeFxi9Sub5ZqFa7MKXU4Q26Q/42s1+qTcL3IIoiF0IePbp8cvnOp0DMsP
kBFsJjs8DV6s6VgO52I9fUxiNBNkP1Xt+aiKm8kCi2nvrh5c6yHc6oEpp+1U
3C4P0fRn+7lM+eKa4MWzfzNHWteTK0fzTTbsrS22rI4NZOQspYHACNKcfQo+
Bl5tqW3LBgc08C0G4zp9fDBBr8A2yf2OHSDdaOOc/sE0XKBSbj5h2IYdWd0w
LH2bV6ejODHWYYyuI5I/qduyzlAD+Y+DXG9a5cQ2/Z3QbN1lA+UKJWDkoURX
dD55VeJUACxgZsdle30aPrAOny9m+9KFLKbtWcaFJooD1QGcuPixuA14QzYd
OVnmp8VN0RFnxpMKkIV4KuS7CBAi3GWqX7HBlLdyT0rxC9GKP4/M+ei9vgOS
dNLnRvqtScLUV5DmfUBGUfgmDavxqyCW1IHbVzveiZs4MN2QLHpNyWCr7pe5
n7NodKnujHzhSojZ55hx6lCnk+U5yYOWnj+w5Y+i5Qs3AnqSdQ6ArIDloa92
gAi0EjyeLD7bIQ26Ux3H65h8d/u1F0FyoF4iNj6S3JZqnSE8nGe2Eb5u3+e+
toOlMouS3XupILBO6lwEXGPdPMUaENwHID96RbkKsPtfmLYoLV3reO8shnyw
rDqYQvBXcjuGNlYOTS4z8MnEtz+eoxxbl7xJpjgYXlpBz8wqtwzgqIXnFZRA
Qmsq7dJuCsx8aRnkuq1+SUqbXcHjGQkCBFVS4EHhiy1W1LVzTgqrkjVBZpKr
0Ph/9k7CuEcr8+iccr2ql1yfV9iKuNL6Lmbg2kNW1NsHBFgmJcADiBXJWYzE
PtqjUe0pGaPJmizM/lFveZnem+LqPsp1NyWHMdhkrLRAb8/ba42gLxHcGZ0e
hswW705FjifilHlYGjDt8X9LYBD/dtVHGfyteZJZxlddyMoKaOhAvBbbJeOB
UmolKwUEbFQ9fTGyy9tIOinhtLisZ3UzjyZMvU/Xhp8Y5SHbhd+1N83UKEAI
xjHDqeXL6X3hkwd/3ILa1NT7YAWWYETsLU7qyAlK3OPe4sEbwfzn0V4w00gS
kDdQPMiO0D1g6RuckrbkxOVprbTLUtcjMw1OQRfiZQiC5ycj8sObiMnEbdag
OlUBaDEOBj5Hb9/8gEu3dSyuCnyMFKOoln2hghM4B3NavlIscMneqGulX/cR
OKFhvfH6eNhl6CBjwit1PMTp9XyC4QtIN1NEqDWEUTHNeiY/94XhGy6yQz4N
KBaMkZaMlC01+NJMjpXAXxF3Ib3nWiDLSDXUU5JZUBuUROo+uFVXZ9H6hnPk
UqupsJ4u1QqCJ+0T3gIG/67qRgM3u0cQHPGKhdjkRrbWlSMXCydZWtll6888
ZNQqgYvDMsxDIbo8xEN9zOXNhyZtfPBfqs3Jf+tYO7C3RtR0xa0Een2Shsds
voYWMC2i0p8ZAssAnAOML5Nx4j/tWdcru0Mg8w5YJxrv6AOGZEhVrkP0aJmi
0Ny2rfJJm4gbGEkaQSEtlq+lyib3ZCW9HsiqqUEfMuwhbPBab+1jcoL8jnid
0HYweSVwrLVPAmslzq8LSUEwqUb4gwfjLEdqBcmzFpnmmSEHSLKAVBwbweAV
cLKAIOP3urLwAew07ViK4ARUYg2ozHGdUjSk9vlduMYv0xIjx6GQMACELp6i
VTOZjJXHKOhr/fdipx+lzN+onIhOJPXHLyaeGbD0eCAATjt4EuOEKmDdvVZL
oSKRerRhPWTcYS7PvUcdQNgQ02x7CckciJ6tngOTLDaKerjoKbCMvWlfvnQg
6bemG5rex0WCwgSabRT3LQb2FJc/kYI+0MYS7UYR9M5zxToI0YiOlBKssjME
deb5NZJ5eHFTc7G/BLMzVKAXl7zhZseeji5oNKPX5i+0HUQ+tjkrimV/ZQN0
IXQTlCG5DXQw7FImPEQ8RO/hHpOjc1UweKLp5uDZTzQQY0kqoWFLRZoV2oYC
vr+UVPkcU+znmIYOtGQiVD+vIs8YMD8aQIjBRP75CpK9O0cZQUK1m4qQ9e/f
khpfKQzMSfRlRyjNLCxp79GZ2zMIcKbWoigOFqnzD1OeRnhwcu6kdsTggLJZ
uC57gIAgTRfyROnvhXnuCOeBj/mu7tBDX0jWgpw5+H2EJMxW9ffesogye27Z
cVVReSUvUbzrj9Obtwo47cYZeNhT8e/vu4y2aoRF4dpj7HIIdwq8BhvBRwf7
J4/Tifv5ejowlX57YIZZGS1oR1ZnB6h+B92Rkrea1oFacu7ZPVCmRagAUCk0
3WhCV9+Cm7XPfXqBIHlFysDfRR93G7w9GGDNdmzzmQb2zBOBFonPJsdBdPOC
91JMPz6MMiP9XH+KS5mqutKr+E2aGwvuhrx2twa7W2PYp8cVasERF+FpWPZo
wmgT7Ln2Ouj0PoYbgOwWmTKb8ZAKCeAnj7RjnO34VlJPELa6hbM8DSqzHgDt
yJTjCI50KlMW3WDx4zRnPqG47jLP4ZTsV1JUIFqu2538DTrnjo7KDHhcNYPZ
uAIk1K1JpUpeAFKTjCXue1duYdpVRujqEgs++jEciByE9tt+jtfZO9NeW6p5
1zT6F+J7IWLnkcuxAaI+gbmgk+HWQKqEFtWN1Bd7vr/eO4JfjD4cZgipk/UV
kJBGIx201FGysW7uAuLCfzhWwM+NCe7GepEekfl3eK3KGnJNx6lRNpYSObQM
8HzkK1Gdn8OlZXqIk7Zdpgo3JlOuifcH5zkrsKgMgYl+PrrtpU4Qdlm4VbWl
LtpdyP1ZsAzbcehuOM+0yEmRy9sdv0hGFEqS5ZnfHjKTYM50lFTTSLRRTc25
9+G+sQ7gQsgNxjO4O8GndO23O8fMWU0Mzl7px3gY5rW8XMZwxfZaT+8RENbl
9KQtZEpB5DCk8pe11T78GxoSpcqmCPJq13qPqqB+hoecU3iLnOs2vRQ/hXL0
JUcF3TwziwXK4LVtGCw35egJVMdIMX7BekHZdZDVgl6dh/GBfKjg4N7ax+O3
6iFhlKV4Hvk85gXc5oGWEl3X+zQZ/xYE/eMM23It3v/BX7Wio+3W6t2L1WYp
Cpchm9oPDU3MhSMUn9xQb6IVv+QJRQG/+AZDfWo/KdZfvo/CA3FjR1YXGYbq
hYZUMmfZe+WoxmHL5Bq2gBxSEedqkeoA8D/Pr3OiAcG11gmyiiAaiv36deYU
fb3qbrqmntWeYPW5KBPkTLbeKBY/QciPxgnl09KSJ+jtatBJwQiM1/MS5mJ2
yiUxLfU4+3jkivc6BRfgGNLHzz7Dd2ueR6jAgZ5aicKP/dZd4BmAx9l2KKLm
5n8uDiHY7iOBIyT4ghhyayLvCDRvEUv8iYtLw4EfywUnPN4/tDzqv1nqVU8i
8QasB41SNgbBjQAiq0T7FCDMTRoCdiTEs7YypKwfzSFNYKgkplBzBa36vB80
qXWbdk1FGoMI7GIHsljbEBdgsyaezV4lKzouuhTjnUrLbUYgmnxjrTpX/F2p
sTBEX0m2yPWKiUmKvAAJrzlcXZE8D2usCxXUJRsn2yncBCQ/TF6wk3rC6qYc
Cu9KXBhhKCMmYFs6RFS1yk+TiYcdTfSCDF1Qbnwqg4ZfHsbPCj1rzgrbGs14
PVfMcb6TYSHgohEXFcbW7jR6eyWzL6H1GqEy/LIEE+ymwsTDZqkzz8/dek3B
0PEZEqaFpJPeTQph2z5F0NayENAAgAmSW0mUpX6K/kEuVtkjolQrls4b6UBJ
mcaeQNHYUt/luwv/2dK4Lkq9mc/8FpyG04U6tPjNdCXZTC4W4MDBK3Ytrz9i
2E1+JpZ9MzdWFnVR/DN4PH9FzBNoJ27umcyv66xV8gg/v5Q47aYBaod2+430
g4VeRb3uo88u32feC6w//kOj9+2p1PUEjm3RUfwGrMXsHDAbT1Jp2LkJ+2uV
EOWouhY9s/fecoyLJ3lG0nHwJgYaDBO+anOZCL+lRNHVYgLx6a7cLlLDoKg4
aOR8pAx9eXpG0/4Aw/Mv0TZ8gvhbIEKYeGBE/4ZARG6A3TNXCFvZBbvHvupy
8BOyif75Ur9fR7gvhASHhten9kbejHZuwLzR/g3E4jS/OdeO4y0Gp1Eppan/
JrQsziJEvpSKmvangHBEa8tVsL2DflLf/UNAQh2jj2gOPBQhOwj8stPwhPw+
tWJsF574ES7vxZlZ4OHFoqmM+/C3GDZcK0uz+jBSvldUTPUvRI00ggT6TVTG
On4E/FDvviQtUDej5PR2o7VX2FYAS7oAorcgAA8opstkUjnFiN1OKgBEruJ2
lkSXzy3fhh9BmYyUY72KeVjuaVIN5EKyHj8ncp7ZeZugPFvjDLHaiO7aF5xd
G+O8T2YVJtHHfPXtDmxuaA/02+N3IL6Vj5X27RjVQvMb4C50ik7lU7JZcUgP
1dnjacEtG5UvjiZqm8LAFTxlrAtmOqkkT1tniCUjtCIZZxxL1XcbpFBHMaLn
6EuvEqe3rHwpfdHWyKNZjMvqN9KY7VR4qaKhgjSvk2li57dQzj9atoCRnWBe
ksAQbEMEAABsUHR+6inQenRoDCfxuoCHlNSgasd1gaDEX6I/LkiRC3+E513j
nD9TixPEb5kmrDpTKaj+ym0qo2pXDzZX4pW8rGkDprVbGq9Akq4QqZ1rjPHT
R2u7Vq1gCA5+7AfXr/KZIa2mBJei8DClaAZA31Z2rhjHUbM6kUsfCxYNLSEQ
o2S8Rn8gJV84HRqvuh7i0otls4LalKxWrYJs/jLI9QNXEszGfyfzRzQpngtK
Z4OgneiPsopHgTJthrSQG2ugxrMlOQ2ezL3YrPaHByS/9lU7bQsorzDo9ZD7
FkG2eMMfJo70e/6KAiqHSm/x7sclR6UQypWZTHe2QpRxkY5IQMoppjETen2i
bQdV2O/fcbS3+9BAW58bvZr2PtU1WrUbRebjVaymeWW7DPde2g5RGrvI29Fi
1RzsrCJDyhV5WJc2QkCyAZMtmRu52mXz4J5bPwy0Xm3ZWX72vwyFzapYT5XR
4hIMEnOFzvVHfKPeg+ZMUSfjfqgaXhGXnGNa2gImOJvCYHY4D9waMRj4J/c7
c8Xzj8DOY4zclGYXlltZIf7TeYybvCOFX2JjJ2sZP1Zd21TGGc8HwT2EaIvq
wu690gpy2ihgoxt5lRW1CYOFHApci/7tNRNK4IjCiRXSWFncHuHV2B4bobue
Hg3vi2OtWihraXgCbh/4tniXdp1i4fNINtVoeaYK8YN3ttHOJx+nwjJmEiSW
1W8i8XNlNQSafvcI6cPEihdEB47lFZmpAo3qOH6PSIBz8JbYEFz1wV5qtwPr
aOQj6j6Eu4c3RsrG52tuEUznk8VBWnIUnIh19S23xLXdcEVVkLpoywdNugUJ
GgmqgpqwKpM5fTEEmlqkVoy8AFd0hA2r8TFXZHhW8RE1AAOzIhWwTvm5rEO+
LPKYd2UV02jrNMjqeLz2oGPmwo64IvzqnYoNYC1mUydYdvoZhVsum7xRu+YN
jug4i23v47FkVOmSW9Zimo/ClSUUjQXZzxeydrzBf29lYEgZGerOZXQyjGOT
9/Ior+Vy5y4vtjHLf31rCW4lVWK3cjEukL344Ty3y1lnwqQYgGFkDPeq25BX
xqK2G6ZWH4SYkebjM7qPOIHoxZorauV1GZeHnLYAWcebCXgEpm3j3+8Ztk5U
YKHmCS+0CTgniymMeqmxlX3LFJSz68AFiHb3ZUckGvqoGbzfzPqqCxgaveBw
ehrsHjpOQwiBFC1ogv1+yCGewxnJovd4khJHgJxU5bhg9LBQfc3eubZCVsgP
09TCFT7SOEjDOlxU3QhnW/1/XFondzusGgdqU24k2NW7L32Bz3uRp6ELvbem
UCP76hxAUdyZret/WP1fe5Bej+ZbdLx8IShKK0exLoWZcB5ghfOVHrDjqAA3
CVT2ZaHxFyR12QAIPYAN2uxd+InDiKxcOwKbbzIaLgZXOdlNJHN4WSoj9ZAI
q+B39dZuuZZVPMO/1cVss7olaj5qMrdrKIYgn9VSQC0cxY91HrJBbEEmnS0k
6vkfJsiSAY4FJbDqePiXZOZOZRlteqCuMS5JGdSesVGNUbpNU3epPS9wDoLD
nKJ2TR1zH2UOtVvscdfenteUMqyBEvYDEES3jAf/xZkFefwPwyfko2DTfJ+f
LrlENML1yrRQUK6IGkH+gseeazKBXAYsy4KsdQ/CKI7Z8iBQrTNZtN6q8pab
WvmCTGFNqvlEvQ6Q79I/s/QRBsENY4BLwKsyAYUk+HpO7h1YrTL4vHHz/T/u
600B2xz88Zkw8F04RdivRCKNEqH11QGdmlIaJckiAPKr+D4/UOALPgTxjpu+
Nw3hxHfSh5O8CxPVw5eldyJTh0Sqyv8iu5lhhZX9tdDS5hZZ7n3JbVozYv3u
jWcZdph3zj2yetFIN8y7PQIJlJIBedXacZRW3/4Hx4LfwQfFvS3j5N5txymh
3TcjOvz36VGWtyx6OosmCcMlqBki8uiXKAbdF53rOEgWyYB2mD0O6X5ZgQZv
/4pS9n94bnESrTULCApWkYainppc8ym81e00jg7hLz38bfH33rbMLm03ISB7
QBgQLC5xXnj+zz2tkNYGpQ7C/p1458Vrl8AZ1Pt471CJckRMQOFszQs4aczU
vPmddYDIAsnTRf0NqfbQHKdancAzIn0viycEWD3XDN2pak/k4RcWzOJkOCii
ijt3I8aLdpTn3FDG7j/6ICmyoFJ/ZFTVAzWGhVrejSXrlZMieIDIJY5k15rC
vT+6Lojqn1UqWGiXjErtkU2XA8sl9JO63UN0xVSIYrJXt07Oy630G21Kl6WN
eCOYRTVOh23Lz0TxR6P4ryxU99JJH4po2FY/k7U0PTtm+5Kr/qk0/VC2XBdM
uzDzRg38QCIws2kRp2P0Bn78LvuxIoqRjGvFhJ/YRGSB8toJkmXXqjUa4V2Z
IJ1UkRsnbON77MdzLUDHsmS8viOdhrKi2hrnW1Tx2jiqW+BXmFZ4CaX33ahj
DcZGpmNe4qh/5te9pF9nH9bfciuGPW2LMiOqa0DDNkuG+NLtJDdZNmNjxqau
oS5AfWVwEUOcJ9FT4lszjQV7qv2nsoCQENpdhoLP8L6vKPZojY/2rMH4+bGi
5sI4hFu/Ol5RKMsVaNkPttow4wKobbV5RiPkZeT76DVAtTk9kQuVVWdEn2V1
nRZcRhqPDW5pB8FTVUS1gpMQF/xz/yHzRXTDJM0XX1UC291zlQhKWub+AfOS
LE0jE4HHUTLLQg4lMBQgUFkwro/LbWYSHFzT3jXI8DCLPdq1sOr9RLemN+2d
uvtejnf9hEWMhnCl0LQdKiwIHzi2VXl0DFzMX25D9qjkpsSEAhKfGPUGFp/w
g1bnxghA9xBYX4tI9vuHrcX8RBqofh/PS0Ddqjlaw5w6KYiZ+GuAwId9ZdDF
MQ0CW7QKVlVy6sLLdf5sd+/YmebzFevUP4LzC/GfbE6uM9M/y5Nddq2SswpH
ntreCBveARtMuhFZQBX+0MWsTacEy0IrgRMhR2FlrIdgdXd94QImeeJEeTcM
f46/rdsYXgmfwYO0N3D6XDWbhd+mfhcadjqplhzVfUJxCIKt8+kAN8cPhfNT
owsnm/j0ZVw6MCnP0LOf+XzTB9Ubbf2kgIs8Ikdhbh0fCMqCXby93KdRsETk
aLnBGLg2KIkzyHaJHLry0G/sYK5rSz9SGCa1IZrX5gtwKCpkduoF0+NMr+u0
iYLrzZUe0bsr1tpwF2HJbQDinucWZ1rHUf3/vuo4+86tzm+DOVrCjKNV/crc
jqXQYrPPtVw9qPrxmUloyI28HuxWp3I8/do0QV9mZ7zYYWuMeTnXQC7hVwRk
8a6HhYfmRbcWF+txgX5KFe1IBk7/VlFLXjmtvG3I4wcdpCuKfgoDCPAPSvbJ
h3bayC8fi/drm8rWCJc+it8jT41AZy8UgsHBke1DGj1xWjTBXD1WR+agdAv6
8Pyt9Lq4fAqB7cpZalZSONKNuhFXKbwdJ4Vj8RcDIs26XmQK70lboXPKZdx3
MryrFLd0aDaKch1JKACajW6IkuQRuewUP8YQK5HXi+HwQ4ORovFXeQEvOs1H
u43tv8/F08WY2YohHWAnnGc2ztQzMXxwiN3ztZ4Vot6LjAFJVU/0S6nNf5I8
Th7S3eEUWo6GRa+z07OBunp0cimbXVgDaMugftCUuR60LR8YjsByTzkhz3Z/
9LnFPYE+SGquHSoErZcXDkG/S/yPqWANJopFv2kYEyGx2jhK8Ee4l7nJbih5
saNceX6j+SRUsk0PqkKCmDMJ/Qeyg8FoeuF16HH1NinBOzNkkCWN+d65bktw
XyfR9/viV/Zs7gL8XMvayV7032M907aWUyH3kAhX1sgURsSTJq5XPrmx9G2x
w7pq5Fq5EOVnV5CAVVOMrzeh7VHZSduYNo9BNOMHG4DY8cf6Nzfr4vtfgvAK
KYI8KEyL0S5u4Sx/ipKCJqI2Q6owT6l80oTIl6s4v9gDpy55MRwhNiECMUqk
dpuvhdXoJO6Q4v66VG3ISfXSXK8GBMAMzCT9s19cDCZf8IMmRzA1k1kNM+Lt
Kiac5QJgyCOLttjOoG18w/+URRf4cZOcYWSL40ujzVExPXomq5Wtn9EtlToN
os4kuGj5/NHWLg9aAyBWDeGnWqML7m05psH604/O/kIF0sWJFyeztMcMrk6z
lv79yMf2RO1ju25ALE42BF58YQBzYHHdO8mD+8drDmh4Bgn+DeIUMbwnK9m8
IlyZ9hlQy03fxHqcj/JrBPFhoD8YGw+H+XRxvQcKsRFznDbgwwu+qeAJ5Euw
AKCpEEmqPQt8Rl5D5bEflhhH/S35rujZBjs4034GVY/6mEwxbBXxnzjdCyxN
y524fh2xkLI3fIzQSkyNhHUIXJYvkGQnyUmeB9vJ1DTYn1jajTneMAP1y3vx
uD0+3L4VQsygsKNDFWYc/BEeRaDhiuBK3WkiJeqzZqMPcAmG8RIwi3m7JYsO
xeI12KHZFyeebhPMVLukZD9lSkVJ/sbFykkZ7c44REf7HFiDSfS6lFrN7DOA
+Cv8O6NX8V3NFPdJRA+3Owc8hPTWbYG25ud2aS72xEwptYDaDm2UBN2gu/8P
IezQE3mBKmOpG3wMBteyxklIEDgeH2Pu2448f2Xk5f+gbaH9NxbGSisUFyNm
QMyY9X3Z1O4O+Z5tMZBo5EDmNBbLf2gsQXLDeIiM6HRtyJBq5Uv72YrnOcBj
JI9QEvxOcyOU9LEnz+yH541rCR8lB3ZzNBzOgmaBPZfsmS1Rp+nhXFCuN/15
RnE6QWM7AJ+wB+h7D2vlqo/u8C76QzbghpBPG23lndp0wlNE31T4BK4zP0MT
DHPZ9HRMWJM8ICTh7WmJTge/bsVpAfWnk00XiMnv+GcZvz3XiPwwtHWrhqw2
K7j9yb2H0UmL8h9Hu5ARnx3qwOp9BlnqMWUIW2GTlrfJWtZ6F3KeOiGBXxfC
hyCxtQWao7fklCvV7uFbZyO947vx3rwk0J52QtmuvCWMQnacoBPIuQwwePZ9
ghOddVdX3MX/2xsBzIMz6Wl83JICDdf6m9o9c6fVUfiLDpodYvbmO0C2HUz+
CEoIUEto+PlkQ3YBR/bNS8K9nOMMIH6YgpV+CshK/fRCSMsH7V9cunm3DEqW
iw0U5AotcuzOOeXqGx9IHGtd5zt7thi2a36agLIKH3rHwoCZd7N7YitAlYNR
imCbO/O7Bd4tfSUIhc9uQFSkWQuEi4BxR64BZYflEfElt32TYlbYJOlzWdr6
42S7DBdcqPJ5nXYEGz+SfsdsNwxynLgR30R5AG3v4DSU19tkyi4kF9Eck/MB
06UhmwG83hpGdphGev4qyybA5Vu/uwfJvia7P1GTsN2bVJr3E+Z+4R+ZPLD9
jNiFPKtKJ1H6o+bRgdEnioa+BjHhiKKTkxgtOyYzcJDEf1TYHfj2MSBpqOfG
kEdg81/1vtsYI8p/8wkN2kZkmw0ilxmCEmXUhOLY+SuuRsd8rTGwNcl2kE41
aGGv7rnUBDfuAiWcpXhjId6V+McT4p2IQHDqsVUIdsPIh3D9Ayo0JVbuGyck
tpDKTIunLsUO3k40JfSKmUfI+OC7Q0xezHstLOGoe0D17Rnyt85nfk7mo5F0
19TMabrQHAtoa6kdy99b4Cs9f8otUQw4+kSRhF3O/yjq7J2o/jUBK1RbfNWS
R9yglxBIu62ePzPANG/rpPcAVCGSkq3iVXdrlTclTTMSAUKgdAX0YZ1VOhCh
PRKWnZUsnocSfguI5R6A9/UEFH/qhL3/x8ApxT95kPUyM4tIYs5iCf2rdMwK
XrKdwvUlCFSl/PmyfVgmfjc+IzEvOSrF7Ozc84eLlX3bsqSF+8ANcY2v+NE/
6AEBqWaw8ZU2PqWxMBsXXsbjUO6qJKbtb+0QXoorM/OidegvsiL7VTFn/P+H
9wU4K5Tp4seQ4fThmz5eHpWD4YOFeZwjDUE3OntVC1Xc0adG0acUz/V6kP5r
ngPs+hgGiyv2yNpj8Ut2SS3N5Skj/vM5ymVZL1lQ3RUp0QLJSyZ1sRZuwpAt
PP+JMxPS3QefVMWWpyQQtRhhDc+2NakDZ3P8byqYe6hifOHW4ni1BOZk67ss
DF9AlivUZCMUUD0f4xSq8ILR80YGIXnPRdp6q5bS+V+WnS4naw5G+cwS+a5s
dj4rTZI+waucen5ikuvdBqb0NX2YPFvVi2Mid6pjjiUrXdsST3/RX4kqrbcz
ZKGOIowZIm0wjnWEtrBRB5xo5R0unmGjX4VDGsv3fLTT0HMaWKJ9Cd9jsWi8
ZxY7IJtneYtEV/LGItDX1KfjWKRhlP60GfajLIJ5ZeOUu2kvdsZtV92v0ZuB
ciMwFVsxfI8MYU4Mu9nEiss0pJwVQfhrRzHI6N+KAeP33Z38DkcOfXFkSUR6
5YfQp57i4c/ylwiXCiYbLEkZFB73N/TQAeZeAXKZmNUxVoD0XBBKNsORRgm7
dpp+zyPLhjoMMvzIT5awnSYkAIBVlLBd+SuGiT8tLuAmK8b+FVJD48gmtFn8
1eXMBkrMpbL3UC/FQyFAkfl8jegYby1qB4/DtLy5vkd9U7kZ5+tsb+61EB0I
tfdsgaE9NfROu0KiI8GeODCao4jAaNJhT1bmcft0kWFykBFfXLrYb0VTTTBk
YCk4vsa/UQrGQ4c3qz7scQVwwndUnvTacMJir2DWKqENPKJ2nyM8QsUnSZ9r
Jg2sqHuxRuz2D8iOLo3pxvkuifljw6PG8UCCf8uwnehDM0c7sSmq8FN9gKU1
tcMD2RCgHEJ3CEflZAmrtKG2pcib5AdAAWWVYeikHTXScxnMpw6UgQGyeHEt
h/kWHrzkVxMlXQmvp6NnnQcUJHf1qiXQHDOVwv2yeAe4wz48NYApcj4VyQI6
XJwX4A46OCu7XjTHuZR8Kl7vICrpieRH3uw4wY2DwCfaWEkdmQFyAyqlJzZY
l4igTfH/vuUvBsMyrvFfSkdDUh5hg+jcIcDuazRCLM+9u5P0bOnxH0shjkoZ
IiGBUbfUbAq1qI5clw/J1l/OBCwcgM8ohdgghYqlW5g0JsapO/kylL880x0q
APgi3JeApKqInQzW4wEc3u3BNVVwNoDRSid/U7KTqdr+2/YYe3ca1HtfGwrz
cNgC5mjDhf5kNzYMNXYJpG4P2wJYmWVH7x20JXKID+zs3Q4Bn85P65Vi/fqa
uzdS+dHcQAMFldZJLWXMk7sz73aT1C/914OpVdtypu/+bno+vLHGlW8lNfLO
GPp4YYgWte6tz6Tsi1CNCh/4GN0nzmq5fxs6Tc/8VV50pa/Rs46qjuQBGI2i
5AwfyTzO+5RcyEZHqrXN1AMrjxrObV1D1Tqxry2ZH1fZf5MJI0nNjGBEUU11
y6d1zWiii7PNgvN+XDiSLxa4hDfDI0D6XOpJXNlE/WcTtxiHBZtWjCggpbbF
lGN6IDQQrO+ze9oNue8LA566lmcpWw5yTAgtKL16PcI7JjqPBajIw5WYdkgl
x85/xYMnLhTCPHZ4Prm2okIAdEUwOSt94F003hFDgahqvy1Gtu3l3NsDb5Ep
DSpa9xjJrVxqlTYGA7OJwRf+MDHVDS520tREfEBYwJJi6gCuyLjh63Wl1b56
DkTtDTgvTWEuQ30pzcrgAID3bwJ3DhmRb+fw34vAnaGIUqj+c4PEaEwI0bLI
z3hqsIx1Mr2GOQglarwhZrp7G6vGi+9oU1ISTEpRK/uQhD6sPyfdH1QcgdpM
5t4BdElhlWiau8Msi9IkCj5vVN9bX5hu3HJyg94B95W6RuITDc6TImy9qrwE
dHGt9VmAK7HvhGeY+N4TsmnJMSn4pH1aYmnlgjLvNDPN2Xud1oUkmDWSsWuR
fMewyT2J+rTnM7MlzZNcQFhty2t3+ki+EpRtievLKg2p83wTlEqSQYR4PH4t
FVke2dkJR35fi9XUJ3VIyN/alJ1vFSIDxFxzdWc+hoy7mhV+chkmI5PxKGiq
TfvYyOlCSNFAu1mFuMl0EPSPJ6SO6UpWTOUnFzILuQUAuJbVcqsnuYwygd2U
EPX+R4ufrvA5uMjwU2jTDReLFHKg2DDdkwqHpEJmoXUU6xaKnNPKc3TVoW4v
3sLVCFIPfm1clC0RRQehJL3J9mN0UGTsZS7gEnvQDKyRBHs5GCQhPTBGxw+I
MPL0fpO4OZGOb4JDpLm/mcE/+KosqLVvCajtHV/5CjnYxRA0Q2cgwdD2PZmD
MUP6PjgRuW3BJyXRmFYNpoWuzQgg3fU14vtmaSdEDsr32YaYkCb0K0O2YsFz
ObVm+CukJm72EN4V18qeY9xkxDQXTqxIMkyzU1tO5La5lOSa4K0UrJD7Nbm5
eHmz7VFt15tCQsE20vkmkxvCxt+Xwj5Q6J9T+fuTricOxaaP2OXYpBoJZPrp
N6T2iMhTGhuzKvDOXwdqlAjjR09cVEm40SmsXE4+3uTQMc1SC6Z1gcZ7tOVc
WlMWRYWcR2wuNZnBhVVZgayqODUrdlT1KZv9I93cdmrNoIdrSC1W9eQ0ex8T
QoojTIGM/uJOAt+JUdWBE37eBaKCZ4JhvHvPpyg1JmtfGFRgePS97QSPWvAp
9jj07bv+FW0SNu+ARZ5NEQxay7BF+oQbUiMny7PcjWuehA1rE4+kQQz56JJO
G1eFpLaurzMgmcxccA7o1Um29VACrDsFbQVyqck0cJrKgbp9t7bOlNlsrmDQ
fdSAblR7M2EC8wB4/OhEBrQfzbCBchfEbZsC5DwPTioZyq3h7aQKq89n4yZE
RK7iYwIsaBipVDe4+QgPHm2wqyV/xO1MfEst+CeJXZi8biv3VkppHu5bJHLv
BZRZJgEV0/BpqHlqSuuE2xBDm9GN3LgErABZ4WbSF5lcoRYGry90F4TBDS+D
LGSv5GLZFVAZmRq2paNJ9j9OHnUDBINMAiQguV9Co4H7YjZyYFqrxFi12Hzm
BUqlfUdlQ/fqZkiupqQnhYwQXVLk2rzjvIZ+17Nb5nMdsA+kJW2dRwGYYYMz
Q3PbDPZ36XWcq2hyJuCm62pts1nq//14srQXCKe0e9B5Cd2F0eId1Ql8UtTe
2AnWJJxAHIGICB854n0kUZbE/pznGOOfYYDt2U8RsAVzgB4+qIrqcXH7j2L/
M06KYfyiUJuPyqqviPnynwfOfsACGsdtLXYjiJeV7YFAZE4L3VCVwefQVfNp
4c+Js5Sutjcnu2V0eNEe40Pwy134KjMWxN0cxplwOdJ3O0fnr9Pw5oDEPRKe
WKIPGhn4YDSI3cFzBVUZGz15ZGeTOQjhDnVHn/1daO5iBt+sUvhFncQ1Oa+O
iiLB7z9tOAxxK59KVuyQwUvQXgMmB9AZY1nejFN2t+VeTyQL6xseNXTPRdgD
34nOn7jUCoK0HukgfcoMZFFBRNZuRhtk3nIf2S8xfF/eJfD5T4LWCTeGyRSM
sH/O1LcY/lGi8cuv8nMpyza3dkTIeNNz04JPwlowwmwT+ZnmDHdkCIuLQKoC
44wc/wvAxuc+boi4ZQN8MbYpyUoOdoWFC6EnM66lbIqSB284Am+mUFtRY1Ou
lqFx3KTM0gXC76Nz2xVdLvPGKLgvCWZKMqVCznIQvmCJSYmGwiMqM5iNHVTL
lBmN4PgLdAQN1s+y5dKapGx+fNqhxLAwvPNhUAnvbaZkHHAFUrcJW9ebDs8N
qZnGzJ6sBJaztQOSn5nYvW+oRe4WY7euh67umeg8uQ7fQQ30qoRmvgRWMZZ7
A0Z9rZmBlAsZ4bnQF+4FGedTnkladSSa+x1I3IswQIxa128ToRwfN8aH5Rj0
AIgikTounwNVGm0mMRBEXs/bHFbchIuBrbOFaWaDfCNBJ7oxW/nZLHz+c96V
rSMeQ+PzcNAS22Nb7Em9IcZ0doluvrr0TAnQwRULz66ZX46ey41c9ZxAaUmy
btJSk6Y/sh9zJaUkOFuv9a0N3iLG8Wrqw3H3RGEAUFTZ5QY4/+lAaFyPAOOT
eWAqD/qrl53tdaIUCra9XK2/LcAEcWkoOLvOesS8LiODQ0cbnxbKiTSHEfUD
UGxTnjCVZMrjprQRmAGXrEVHfk9kkwgLl2r8C0RFWA6Jr37tBrnB7QUuqCP4
9awldOeluNERwGjOZHJh4R7WoZdpzkW/Ylu4F1QewskJteBmdYrYENdyyh3u
0irowkntq5jlXy6fqipBxlX9pSMkvCkSQxXNvF1lmzhe45rLo8FSbweFhHZF
NeENNtT4muiHY97mJet3fnydeJQNDRNZNaywDif2rul6VtGObHim/QEpxHby
OLBpMfknmPbBZIrqOu1f6Ey0yqmz4wkgsAybFEKdoQLczYGyPHYWtHolpQAM
mk5y+TrmYA8Jnndoq2gLxTdlNgqI9WmcDqNEorDikvoRSFcBKAqXfllHlRBx
sD/QkeiusoBXmzjZ0Ixw6sfANoVZH3Oaeohbt/dwTA3ihod2C0QQpNHWSVj+
wXaY52mxkQQkeKp9LoYNzgPnMEqr8/jIRFlKNMhAltSS4mLmAlWs6qJfgeXy
akAC9BsibQd8v5c485THgz52e/i22IhicpyePlOUXTPbgoOJBdMwBlvpKaB+
9dDN99ZiPYCM6jN0VpIthiNhiAh6p1AqGKwcRgx7/+JlJxN9wmjTnIiY//ec
n5VxOwycw320PE7eTgzwpGG+zfNGrDR4LMSM9d1w7njy7dqbBz4p8Y/GTx0a
BLMXVejeqe0bOjmTKjqhOImyhbtfIkt4vW0UDRiCQxALhl6i6CwBkZGZMpJ1
YBz3y6CTs4vEkSGWoVX3X/hgHnGSCPcetVr/5L1gatKwxyeS1kDOYC6eR4gY
syVvm0a1XWe4R+UY9GEWpW3oRI87c67gK16via4y0p10GZQtd3B9TqXwwiJZ
CLLlDubvunx+BAnMc2OvWG07WW7eIa+jwbqSkJMfEgpAjjCosFfsS986zNas
9LxQV3Ah/bSpOgCTAYocumMVqF01XqzUwGKOcf7OK1AiuggxFoz5OyAkJhDx
whMUcKZx0jJlgFGXYZjzma5CH72tF4ftzxh4ZKIrxO4LRCM/4lcndFkdqv6e
XzDm9A9S/xR8atDcFTJ5Fmq2+wDVo5tBVT/2UJ54evqmmO4tdsGva9tnvQDC
V2tXm5I3c0ds7nerrPW+9K4jwZtYiIlMUqjHtY6GbEel6c5/4m0/PnRMwiVX
L5D0+OfmX+18dUK6+xPLlj4qkuJU1VZX3VUAr/X4qDbJWx/5vpWpUb7HufbM
gSYHvwqsYJ44luvO8pywLP8bZ/gpVwMAxuClihRuWOaCbC6m0kKq2zT5LGWg
ELJRNFM9otbtr8BOCqu1QeVZ6+ObBAgnhzP4EmN61/3SIg59NQzGF4FKxs9+
70IQZuEPuEzZ3OTcrBCa3SIbitsiS0mdIWZxlONKNdN2jcRY06a846vkqA55
mcIcVipKrO/1Apvb7mROf30QWXy7BfVc8DwTeBYAc8yg5pEozdUg64vie3ii
ok7UDJZlRKTU2dhqpSQVkA2yJT76ylm4F0qYBDDhsvNV70SC8zO1dR5KT/dz
s2IoRF/ub0a0/kC/1DO0LThjxAEHlRD7YyNuNpg/FP7EPVGOb7WJp6818baC
iKqwM4JT6MOONEDh2c4g6x6y2Q/mJIDif2xW3Cj5JPg/RcXS9DS+s2EC85Kn
rGyyrWmP1AkDqxv6+M5UhdJIS4YXwr2rEo0fXgwMm0uYVS8GuwoL4B3d8Vcn
5IHsvS3ll+kuDR4YfLw0tBXxP2f60C8Vq+Vkujzs6Fai8RI9oE9bI/wk+odE
JZB9tsJKwHJn2h3dkcr6+fjWUa+Xt4O2EpTuN+eB21itcscXBonaYZ1okvZu
Hsx8c0n6Q8SftXRgRjA+NyaHdysTwuufNkeBLwpQ6fIq9DV17bceSQTsIcN2
qrzsgWWIIB+/K5yDbQ63jCGdUP9N+DONAKPiHWFFM2mRlFTgPeCf2sIFaEMt
4JKAi5PKBd6kMBU56YGRtk0z3eQ3K4J3+gjO3p22QsjlEb4/4f5Yv5sD7Jg2
fXtTRBqPEdci2bxbaTHqz6mT6PZQnzOhfQM9Zbps1DMwmXU/vurmMLKfPzCv
N4YaM/T7EKCpgX/QIyv4eDqUAK2S6i52pBEfH4uRnwT+cXCvUKnA76POfd8/
xs/Tu+BJDKtFJrAfzmzZ7wpo6WG8yE8zqpT8Ku3LyPgdabSVicurET8EqWmr
3XTGinrJo8LLoqcbtWSnOBYoxJ1l/cl8pGcuxDjoA0+l9xTFrs3Xt9rI5aBd
0H7tTvnHJdQIe1i96hpHv8neO2DAKelm9DPuVk0/geC5LTo7gXASB1y8XASe
ImP4HPdi8XQ8VGk1p/MptVHLDX9sPtg7qhvjMIM9XPfXW9Hvbcab/2c9CmQc
ynoOvL4Qo2Qros4n/aJ1smmx5hoyA1EsKHu8qMdamm1A21VGlzb4wZ/FEGfn
Md4Ddfdahk+x7RGXdxfEoEtUZC9QtRqu46PQ3kWE31QWdaf+BLW73z1RjSsV
5O5NS9JEZazFbqdYyAFdZUEE9MBOP20qHwJK8TP6MBOXm7/j+vJO45HjHcwZ
efriqVAIK5dnpZlThnR0Z8krzPMrhhzWujx3GE7pYG5xOD6IMZfbZOqjE9NS
+387xu7gYYNUO/BrTP6cIL5BiHSv6kIPDgJYAguW4e0FbHeU5iKsfEulij8/
XN78K7NKDCYoIULuE1nAXgezDtCm1iUSL/qGzQymwdWIIXW+45yonAULyD92
APnq1ERsaihd2a3nxfPqwuY4/98ZY/EXrAHLa+6OpzlBXmxO78mwrSlf8V4a
36yjMcCb3yjJxKW4yahgHyo948CKuHJkW/VYe6KQJDXeOflzxuLgtwbT162o
ClKspcpe+xW7uvVxNkPOsP/eDEBZ8zU2H8Uj81pKYacgLdiAYqnUFaeDFtur
b/dt2cmy444aXd7mfFpF9yz7Cq0PvidbOnaLISqK5yJADLcK6Fvy6n+4347p
CVmNrHi29b8jymNF5XqhE0cz4p+r73KEsgYyP2zG2RzlF3oU3fKX7qER8HkD
zOWzr5vU8OvTc7eOk1AzR5J/UpVFXyFQ5NhbdNAA0au9aZl/6qshy9RlHHre
7znUcpd+wMlWoxm4aWxWT6lrgxuL0hZlGgKNRFxaRirirwjSK9LEpIw5PqPc
NcfOo+zYS0+8D7HHGKcWyN+eS7giW1XP4qYxzRaN/aO2fNs5tsMjPKHaiPua
TRiqB86YT0newD1lbfrOwZ8Afwzz9BR7FE5VWg1C53I/k3g/M5WeO1FynoDx
6+UYSH7vyfd7mP3SU6l9PdSYNA3SFNTLyOxGwS47/LdVnkEMst8nueHTCt9Y
qi4+2zY86HRHiwHJIHTFG8Ap+vlIqpdW6mOiYg0Xp8cqLTiKVBSmBfou84b9
RdjDqEaUN0ejTvLsv5xZZpcWlNZtrvwtKlRY1wRVbgoX55HcRLi+vIHujYLV
ubNN21XEAflxtn+fkpmicKPkBOSpuC4XjKkaNP2iHokRro3kTvOBHLNGa50g
80LRac/tbWW1Epwz422v83DMiCjJ1rGK7vkz6rAzaMTPTTmEAQtPgRATCi9d
exH0bIM5GMDz4+p6S6wIdPdReEbKRCI9POEye7ylWgBDQEH2hpRimvNZAi/I
1lxcOa1qdV8mCpcUj+li8fLppM3hllQaDFvXaUaaJMqp9SkoCgt0rHY6piBl
AZa6mCLPDi7gQ6QX3JlJgiCcAvdZkz0PGflj7ZCJbhElXplMXfJdC0eLQyUY
VNQAjE6vsDX5C4FIXnNrR/6TfkrMq6KbqVSAjsKI5UpPX9RPTfD3z0HtwOcU
ZUJD/Ukf2+gVYN11QG2EoREmuYPZb8tHrWOSFOJnitGl6Sn6qgzYjTMqrLZi
R5lgSTcqCU4Vqg/pwwcRh9Euad4iV7mKiAh943BvDLjODhoKhhCOs/oe0NdQ
KB+Vs1IuJ77EONJaxml5Cp5VRkWVQoEUiyrNxrrA5QlGtleB4+IO4k86xx+q
NgyvMQbM2X9ET2/ewrGig1hiy2PAHEBtorkNSKc95y1JeclTWw78yjvCXT5w
4LW2Q7GG8wt8QwflvraYQlpCQo2hnMTb/7saUELSWg99pS5MR7Y66V8lGWJ7
qXgGmoSK8xj2CglcFtWzZ4b8StFCoObi8eSr9njtxonsIkvfSeC3TdCq2H7B
kGF32APWtc/zN96vxHDZ0BAWkNSRNEtj3mRu0MqKmqhcRd84GS/jlDN5jUek
/okQexeDuV547mZzoBYSSuKQ3yCPiZ8Ovp1r0qIh8mcKTCKorvZLVKZyDGSG
NgC2m8t35cxpt0kK3PK0fSTn/n0yqA6IiwhPmyJ3A0sVJnUmUL/3KtZZkhWl
IqTsI0GyOee8VBEGAZidWD8DyMTzNIyW8zJ1CocR4DaPLW7Sq665fT7brWI8
esoPBK3EVpCle4zcIKUXjccJKOk/RVjhYUc60RRlWb44q2LXtqTRc5T3Z8Ds
txYsh+uVSjPC7pEyJeKO8D3bQ7b0McA50TzzWWENdZ0LivQN4Hx/xHwpFRKZ
cBcMxn6MzysVaqPqx1Cib0OWZq5QlIBwrA8hKnUG2pChkXD/T3c5GS6x6bcW
+8ysABdUShew7Gf/+HEyilZO93nG5+0HX1sg/Bbm7Pxv7qUuXCqcvTc8Wgn4
EjLQcTIdc7Rbf5/KTnR3yP1/V7IeqpU0xNFlF9nLUAcPer6tzp9OPdoP66ly
TYgBPSoB6nEsJBk843j4WDmU7kPuN1sOT+/hhJXRBd9cIAcDRhytW6FeLfxC
AwE2TLYdLQwcstNYjvNxuc6yRNfrolZEfvAhwLVPoQUMcFpzgDU/JZWVXOqe
EwSbGPp3/vJv/7ZKi1nINHx9CXDwBfmvnuEk6m1TUjEYn3+caHHJDZh48xYw
P5+MwdX2zADt0WH3lf3DWTUwTHp2xgmXZ05PNpUseC40GIAkZgrzZjLTB9j1
vI9WNwX0RIyRum7dO8Q5kNZIvu6r2ORzpgWVgVOYAmFq+S0MEY9NWTNUlyEK
I/7b7pNZGOIYB7OxcvkjoKvducrqz7CWAX0AS3sm0LzHmUKMg+7hOhD7rsXo
spZ4c9Sz+dr9iZqqy+y90s9OFsZzX5q/5XMQWdyZG4rlWLQvm7WoCzXVEkn7
Zcg6a5DiOdsdCBTdWp4vT4aMRBr18GN+2Qp4PztHWMXfKKi14tNPAZtSpISX
AgkQ69TmL98JuEsCGe9HrZvpyAF3+afEFZ2Vmidg6pAw0bvsJQSMbjnE3npU
s81aQRHJ1Tha0TxZYkmgd9QX5Jw9MyTdEfUXtJ7BZgWswawSKCWG2Gf7mF/q
W3XECLNlGhAk/HNOBYRt2dHsAwHW+NNM6Yn2Ws5o3zHeWZSzczP5952+1KXA
KQyNUK935ZV3jt4aULTBhaP0o18jzAFXH0wE+uHf4RUXDpboNNg7evgvo3YD
shHqdWTEGXN8lt+cEn/Q6OOt3mLS08BRwlioZoO1ASmeKB4rhqIKqyKt8z6r
+vsHEzWx3Cwf0Cq/Z/asqYVDaLTngjWZi/ZhYap9e+0gv/naanL/dTJk7dvm
YYzwLyplrE52yEutn5ONwBDtBxxPkeQBoeR2DAKdYzQwW9hEJHfFc7oHUz5J
eFminGeZJG64zUlq0Ol53rfcVoNmdbBysZJ6HCDXAiS1VrGEuDY6VItWV6/u
ymAOOUcNP9EN9zlBtWxJtM7J8TCmk6yuQZfkVcMDtWv/fBqZtP8wW3/1AozL
wvTi9v0JdsFUlBN9qOjz4ncSZ/nEoQjr71VaDs/XTLYZJ08H+Bb1UcpAtM6P
cmaa9l3DaT7jU4aeSoLjAFEnhrBfh+msruy3SEyQ+EmCxWpRWNetySobmqxJ
OmuiRyj6xEQBdGj0Rg6t8dFBtSJAvww7O4r7ascmodF+PKZfFamhtvCaQ3S6
6uu/NSetUPnb5IgDwm5Yz7j1hhalLENUZ0DpKMB0iLI40i2Fn0d1+MfqtceJ
f/Dgt5Ftib0/jRXeVoC5SPRcmouokmZV1uC7pHVXU44ra2noZIdi4qf5GhLO
2eaZ28ZHErIVkBH1vXO1aRmdnPmoeat1oKqFVrXHDulDwegaXTiRX2cOPZCj
HngUvLw7xywdz/iGS6cKc2T8OA49Vkblu4ng5HC0U4ohXy3gGjKIUcf4B9SR
c+obDjve/HDO24fWPXIljifsy6+1cqNVguSIT0qMwJ0UimWqDOERC2+ko4xv
g94Ckd9cIWiVyG9w6ybW23WxWrIR9qiVmUS9IMFYp1Ul8nSquXJzZGaSeRuf
qMh9AUIAHbHugwbXTNmoTaSAQC2FdARhqCa8XuRcKKLDBo0WMNwxJS/lINZC
Vgks583VkGZ4vxe6AK9DsMJI6wJoV88phPvw45SuTc/BXdqIIPrXYbwfXyxO
bxTSrYy3l5enq7W3g70+EN94lOno0W/9zFegS90Uxoq6fL6vozGVkiWkB7C3
90dABLfSb/p/BE3oREOt/WZu3RVgh7mS8K4XFw7RwwiFqO7xGcKWKhFgyb1P
1lOmCTE82Ql9HoO0G7w1Wlbpr1Vecyz8qXJlVDBqF6yG0wkgJZWYbLiRtG2x
gVab3z2ZlzccJCH50u9LRpwqLr9Z9+Jxj4EdVipEFj0yXSCxzRujxUDw5vZt
3rk3DyKMUfsx0txWmHaElXWhbvmBGnjoblTXJ1A5942qOC2O2Nb8/hI1Nhfp
+wsoDN4TWT8EA1GRsfyJEN/7H8aAc7Zeez/mumzFIfjpUYDYgv2JhpxagX+b
kjkBZfgeZFpK/gb4DohCAVV4cS4wFR0lP+JfL/hsRtLnNlzipP1nqc+i+eAM
LTDSyAtjlmrPasUdzsIOTBVWWCLu80cgmeSRukTw6xyWa7W6YH/5w2EyKvT3
9ec9gRTMPgm6bqWU6E4d1Jw7kQs0DrwWRla8YerXQjEiykVx4/i0q401q5jy
mOHeCWNxAPTk4cKKHTN3ZqNymPI911Z3lNmqnDYwUyoDLMof8gVLC9uXrawL
u9l/onWd9myP9QuZUfQY3RPhlOOZNt744NDgSxJhTvWgtocOw0xbHmAAt8Jv
eQFoCmv3ckeA21BNL0r9L8IdmEc/uZSQZj9z5IfEGrAGJM8YUzud3gv5IA38
tljBGUG+DcNLisRU1EBT+rE2a8nx4tqC/i2XEd41ZZVwjkTRnffLv/V3YADm
k+DuZzzoDtpTm0UpTXaan6OcqIpnSzeTXW+H+WYwoQotNwHczLacJegNNlNG
ZNciMnqYSXbRdRg6Y16Y6FgCMvHlljrHmASsk/7Q/7+kMQ1IvtYa7DrD280y
W/Mlg85pK6eb8Qm6RSUKlpKup48UhXfyv6o/5PkzPnBwG+XD/VChAOu/1fko
B8hDFzlHCXXLTgWljEqreAB2dg5kO7vKG+AMjdBIVapm4q8zB45nA6So0pIN
odfGpWGm8j8JeIzYmDcL2N/5scrx8TGFnMnWpigV3ua+GhCC7iPYgWvbTIk+
W/taKBElorCgF0Ra78I1YYC++QMiaubFecZiMrlxPCiqcPyqIpjSJBWNpiuH
NvTiM4ompv3hPh/9s39r/I9L2eR2DSf+D2eqZSIZvmawsDJKKSwxPIhw2s9f
CmTZAYx6+fZe0jWpSrKPiOTq5isPpIuGv3Xcg8Cro06FAXo97OpD9NRpFcdI
9UYLZp0r+9bweB0NXDLuNuHkQMbNT4Ai8vR+YWFwmoFBmgB4B1M9NLLkn/Eh
Z3igjSvVNT7QPlegS/NUd7AW8VvjPWQqcaDDZ+maAeLMBnDjniF6sDEPYRCh
+HxJbY91nt9jS/zWJM1bU2hk+CcRnYFNZ+emLGXX6o7nuo9qc7Rpo1JbFIXK
yurXT0Lnu9kLlZ6weyymsGLB/5Dv2X5fC5ao5dB/+mYsyapHnvmY3X/291HI
ptmFIeZjMHocVoK2mD1NKNnxQyEd+iiL67ggURoy0XIpoNn0e3QDXy7an5U2
KreOeK7fzzFX1/BDyTy1syb5IfG7iB+C8gLFjCIuqlyVFhmRPljyly/cn0xR
CgcmoTm1/9bSY5s5FTEHNHGgZC0thJ1SdH/jlPkWhzB6DUWQK3DlYjVxXPtY
9vfxl/YU+sV2iqAa+2N+17RVwn/ByYVDRch4wlTZNF2mUIORip1A5h+Pbe44
mVGm4idepFWjtQnnYD7+k29/PmLtSUdpHI66ZmV8XdM2p2jJB2tcPd03+/a7
JUXsiHozsYumECW242kjPfy6QyW4yyFyTZ8ZhGKV+MFqlvfZ5rlGNxwSA30o
sB3Gost7K2ECmBovbJviQvHmOBhmS3KR4OzpX0krb840kfc+SrGj3HNskk6W
8rFHKJV4nMi21nerCwLVtDZoPY679IIq3qk3ahRTGI/CuH8MVCcixi/uIr8p
f9wsnTNcZ7G9j+WARRNOBpaspNudYoaXBtLR+PBuX2sma4z318CBaX32N+0s
7xPxiyXEtX+3wPzQOCjJebvEvqDPNMBPeyw8O7UyC437Si+dvKWMqZR+nf2I
4ErbacHKK3T7HaP0b8M4E5x4cDJ9lqG/XHhX39REPkIka35sSNpv2jEQwBP7
pf9b5iOSzzEfQRzlkxQIE0VRb5/lFHGQPzE4SIQYgBibCRW6QIQqLZfCck7O
Qn6SafIyZ1q2WOpQrIhY/5IUqwDIHMEYXXD11bzRi0TDWVJpBmyTuwwW4DxQ
7caicHcZXWyF3anIB6kmhPUYoMNSNPaQ6dejCOMHn9l4gb3OxbasZ0dniXLZ
lSDPZ4u6kD4vPlxB2MFpGg1S+bU3mntBx3DT/IPOldmh9ENCZEBvL0nKeGkl
K8JlbRdUKdN8kA/y7Ej8FVOstpK83DYC6xOla1dr5olQHROnwQ9RXanNbrDE
AvKNPC4Zmym9pR13mxRJ/pNmjiuAk7oSvUi3bMtrmJEjrfzgdXtQsEn6Yh9n
o+sVRJFUTwzTiFGrFzQBB3PhLdDJLNG+3BbxKHQVspZ9LGVelyGH44xcIVjH
+d3a48ixSRX0xZ5qGM1if5X3UnCRJpUcIK1NcK3Nz2x/x31hF993fKUcaBKC
Q2MAZtjA2gLG2K+f7yB+wgfXj+seaHqeV115L2Dp8SyaR3mWnZnX28Wb1qLI
K2//fkts1BZNToGIaciLBqUMPXn0Zoq4GNiNz+vB2rU4BZKTf0Ztn3kujNnW
MyLSkL6CPld9jfHXpelfblbuaWUZuYY9442LAsviucMfYx54fw1WQAjNdiJm
52UvvnyNXtYjyYb1OD5JhG5n3kEmOPbDVvByd9bqMwfgWJy75I4X7eb21ijY
7OfEh7SGALA6rge/YdvKGOPEB0LyD9mncETiwZUL0C4+8mlhyxo7qWQzTgHx
bCDhoAxNWU5OKoqCtqJ8y8Da5bL1hTPe/xTUbiOVa6UC1JG5uk+6jOIORJl8
N2l9AuyUxgvokRkR9DScN637Bm1SlqxdquY9ZuFv8hWZRn03+I9e9IRm+ulB
jO5OBZYeejFUsIHYz/eK0WEkpSnREpaktEkcFb4tioc1AkKxdrKDEV+VcJO2
AKrUwtoe3DV3biJjssohGOS2HMZVvx/OYRstgKPp9f3oQNpQYpSM5Lp0cBaY
+QdTw5baQkym2ZMRxqLgddFk4Vft0PtQgT/HQNvDnMBB1LCLnngazJqRCpIN
5bnS0gPSiyV3qHukMBT43MPoMazkBnZafeGNx9JqBP8p1z3jWvJqKPlMZZfe
UwSzQKUcRx3TXzewFf59kqYl57pYcb4NGbDr0NxrDzRtvjfXDkj3kqEgbgBi
PpBK9cU6x3mJ7MJCuWb7eH4DqGxzrFpSSHNEMGi6tCC+pxYfTS1fhDRr7Y1p
6KYA4Xu8sIiNmXbEPUrVBuhIlbk3R9thVeehqtXtD8SBTlyI9Uv8ncJTSnxn
f2BdHDAIXxtNAzp13nUK6QdGSp36JNJlvUqElVbaePdkYNfhAULMx2SClUto
bUtpdpY1uSndgWhsVxZHTyda5JIalXbIUEYEma+ZBT/a4sq+YAzlEf2Ai7BR
c7JNrgQQMoN4dq0rOSJZmsP9ZDdPcM1U0bJe9UpUgzyga2lAD5Z6AGvTF/Hv
pGTLluag5kqO6zKlkER6HWgX6+NKsd2nyECnar5bCmZhipBGTd0lRyYhi3AF
4R7FUM6zl11F93tzkQfENBQ/lVdooINsuGxeCjBlQQejBLHoLvC7FPXzaGl/
CWZbzczT5J0C6VPLb7Tb/oDv9N4+w+POdVEqTHgn2n0NG1p/HEYok2zdq+SB
dGutKyQ2xUVGhYfocIbqst9mhdbdR0eKktMH5lNp3uKNh0rvqhtMM9Zd/6xi
jRSP6/KlkRMWUMQfqbwzHg/jMfU28eudHtbxS/hbo4HJaP8Bu/rGxgALc0Xn
OFusV1xVXOBeG2bkjNnrJ7V3cxMLtPRrn/DLXKuGmjL98hrjG+KZHrptD4Oq
le2t/63aOKcwXH7gtk4Q4gv95FtHvr6zkrlb4vNx93LQSUyAOUpwpCDw3rIW
5qwDD4hbkSrQgpHCAwem6XB6I56rihxauvlWPir0iXQFbpD5DAWv/un/Cvj0
7sgJwBLPQYeqShO1m8+8B5loC10/uLwOPJCTRoiaoA6+DVh8hIWA0LGT+kv7
dnRYSQDd4TsEk3BmjgdMk/AB6ukTE/lHBAf4dQzYuZ2WtJkJg2M4P5BxuG4P
XcxriAEaH660BSpmL6DF5rTzwVgwl0Afh43xn+TSI2VGq071SOpQIAncaoFP
IXV8sOSERoGt739f4XoHNgxSaLvUsFCwZVW24FpK7daISkrCPNoPrWGPDMcb
Wof2Ii5r19XSkPQaLK39UR3+yXK75DfKMd866+Skkr/fGRVnyXlTk67MuiB5
KWdHBuyiaIectHZ6dU0nfBQZGsoG5cWI9GKt+MhF72VoWy0SwwQnJET5k/5/
7feVL7oDztzpCWjvkoc0KVwTlIPi8PfzJvhuxPel/SSzUPNhnpzfRwfT6gbU
JrsfMi3L93q0feoB+vIUT/DjJHEeVJXcKwpk8r5Hf5QxVZ68PZXBb2EK6WJB
afX74/pWzc9dsdkf/lrWjUAMef8Ekc3roO5mBhgpA4uvhk8iDPzFsYKS3qSg
QHqQPn9XQv1la3/m7FnEW246ebXSy7In+FpdGifHT5vR7N7JlhKUaAThdWBB
0kyVbpk1FKWF0451YFiZjf/ro1SJX/51HGwZ5C9qztsyhvk9gFFo7qCGRBIb
kA7Plbq/Avke2qxe2bdTpE7gLhsl8u4TMltfAPPOxN/VKfYK2t+KJvFtVV4F
xOAla+wlTmAYQgmmh4YqXunzL/2uOkdKRBjVGTwruAQRunTmBvJydM47l8YU
AqPMC/41jZdOKexq2p/RSVhDyyGV5hbFS9nq8x9/G4Knzu8vf1uNIF1JH3rX
tJXEfauXTQ9hL4nCcHj5QI+Jm3EL5La0LlMUfCm1ZbrLVwnZjeKy01s+1xeP
KiZzaTcxALLQ+GgFAfTS9970Ur4joAhzJFx60Wqine4BpBonl1o6erqbeiP9
zdH8rZoB2gDcKzYuPNDf93tEyo8xLc1acJcXmScJvi+W3KyiD60/LY4ItC1q
IWVdcOusubH6k83Nu+4ckxbokz4UOIQKTo40hefbDFl3jzD6PBI8QaOa0fPB
DFpDVG/fLm1zfMvEPLFYT3OgtifNbSOb5fu6FzKATO6sGndyViCKOg1syYPF
fW7oiH+TbcZ5iSq6H+CJqVyrZlTT9SUXwOMTRzIL9cxoqYQy0OHJJ+24Cjoe
5/hCfIbf2jVks2lEJeuwDWCqeUiRn1zfD6fQJ092oIprpwIM2Y4Tu7ddHPC+
EU1MrdszAMOI21VaAe0YBd1OAPJcqaKnLy/VU7WLv/D9jaH9tVTVKBqsAhnL
AsXgq2cXL0oKHUV7++WJaJIkikaHcuKvEBm4vTwxfa1WOOKm6WghN3xolR5q
ReQ8L3yGKX678XK12AtOdLC1XW+amU6xlyptrSLOY/o/CG74wR5gypMLYafl
d63eHsl+taAuD0A4LpSaXrvGqu0LtUhg1Y2ItNXjnUchUdopTRW7GvCBdCU3
Ty52YtN0relQ2lkJ/ddTzNGlvNZ7YztvjATEXCzuC684rstp5x0+qHR2puJM
fvtLaobDWgVaeAN37ejU6YDqEB1dxwazWVD4YqS6KNtpvs2VWL90Tj23cKOQ
swVTknOzt+8bp2XUmdJ+n0ML5H7N5Qjd1jJbWHkHq+v4JafdO9hKzPW4NeS6
aQMBCf/KcojqY2zHsgHk1krBCNrbx9yb6rdEM7u7Y5MCpygFS0sgBXJG2rCx
uYW2fR/x2rI8rwTPSIG7o9VdHGWG8CAzPoI5m+Y3WJor9pKMtgyWJSEYsNtC
lgQV4tHN1P1Hn6hNxWPHIiUWRNvn62AlmrW35aK+oPXVtfr2mMwQb7s1jJa9
ix/8P6EFBA9qULCTFuDrEfMlOWyrn+5hGTQ9A6XlfMaIEIEDQlkfCSjcHwdq
8VXWfPYBxDK8H06uMWfCxzgdXR6hxl0EW1fAwrT5ytPJPmfXt+iroJUM/vYr
Sb4LJ78uBVRXoCimlCzzR/7DTtR6z03N5AZ2DKC9oCtBa1rzoMauYJHNzPTC
p/0bYcATmk885PmIIRMZqVZtYXevAyLRwt+ZkZupOL/1Kvxm3kVqiMLOCyHx
dENMOo4E/Fo00S+poTknOB5SRzWABtPv0n+l/62NERguRpA53FyJnyX5qZu3
THLTUmSK0VcaU7uxVU+L2gCbX5da9aVwsNh9cdKzJK8NX8Or3BhrpCrWoCHk
0YFgmfOMCrsRszYl/fw3yCqtJIbYuzwE8Rz4SNtdp/H1KmK/TyLk/KDJpwGz
PqDXmOI/qtIq1hkZfCKfyj9qYJ7oD5Vkk00FuDyVlhUPNrF49PEo9GLedjSU
zmTg8rwI8n5hWaOg7KLxRzH82NKKE9V0lLq1wlq8Hf2d1b2pf3Z/7lbdyVu5
9xU2lbnrHYl87dosuIYanKrY1+j/l57BJrnovY4PH4Mo13RtPTKMCi5umiEA
cALaKZGCpLM39OdiyAubXeJrLF0cCj0a9WVE7A4LUmZSpMDj16fWXNCOcPJG
0Tns93ClfjimX3XFCDurGgEDuo4tVaEdkbDyxhmqAhc3GuJnVIOUBKGugt2r
isCBJe9IcF8BY0roxBvpJbZDtPQaDyDzw2oSs13tczoak4sD9Nm2JOwHWTxr
JsA08y+0Bb6E9wKDf83o7st14BkpUc5JYY6BMWf8YJDQUXuBLCT1BjPIcExw
Zqb5/tnQzBkSAruQyZES/ovw0IrfQqfFtkkOfUxUDRTT9XY6dyJ51+z76H9W
87FD4y/nUdJbqFOOVKTCR0vw9Bbw2ZJmrVhN7b/bcjgPJ0/Yy9NIUH5LiX0E
lEacQoYUCucXIdM2VUr7tYfiiTKW8iD9CSaPWCOjRllpOH587HFmtbWQexqu
Fu120HPAlx6EgI6wIj1fWOf/5XXlM/QCVbZlw0WSpuU7n/s3cZmPrl8un0Me
8gyPDiGXBy4yej6Ois52OwIZCpLcKNBUb57bPwHWGJSv5rPGLJKHFMFJpoTS
gEGoc0X7LPl94/Y2pJQ+oObk7Z5e20aZtcgkfQaWgVrnH6kIFTa1tOI/NGyG
jgSzLJ19fTnQKZBIS5SNYKKTtz1DUm+1BCZF+2OMK/sx7oGpH0sfJys7traC
ffoe2zL9/LG9NAI8/2MXWefnnT8cwo7QS+ypqOOtxhaXfiZPDEkaZl5DyZHD
F5HCcN+YJA99lNPVSvQZNzqGxXbC5QVW9/FU2aAqCOHHsoZPB9i7c84g8bfF
fNuPx/ambA6Bqh4wXGHGv4/9RVfEFzFCDmhRHsQxaw0Sg003wuio15BigKPd
2VV1wW4KNccqraMaCKcJrI80rXHvnUvSYNI6FAstEwisEvU/HkM/55vl07aU
vajTFzLio6NIkvhZKNh9DOCpk1kskHJmLU0zLptey0N2ZpMVVAuaHvH19pi5
wCNgP6si7KtW329I/JHqlECIG8kYf5v+5/8G2KsD2+K6Y4fFA/0SW7gDjRsZ
WUShIcEwTVobp+YodSwnRGZZP1hCU/AYYF8py/STljT83y3v+CRq1V7lwYup
T0axEd7qDPz12OgMOnfGsC6UU2bFhzaUmyj67WeX8Ri4bIq/I9ggXxqxv4go
DAc2gLTlVmbRInn2f0LPxEUtF0jPFXIwPfGN42kAs4Ho82Y5k111AYGpKzlj
XutLTBtWsNlsAEXiQULJiffofwn2uTVbWofYfQVs/dvCZIIqxZQ3xHc/9DB+
DjoMouw3inXPpLSWsoA6jP/5ebAxwv9nTaS8lay1vFWPU8fko+2G5VWaPL26
1qriYy3xsgjCF6F7w8GsE0yPw0bHzTSAoTiuj2eK7x8UFlXWRpPC7K3v3BUi
IUvRQXcRZr/6WU8SYJqamJEJeLBmjLNUoWw7ptGAQngTSXL2UvrHew0frIQD
75vu5dcT+ZUpXPBQVycDE7qkfOmUOl774LEnMk4EaKQP4xujWh6EpNE4Eajm
5grbZ9WeSh1S2o71GosWgTkrbSgyL8CFj45c+F2Vne1jvax0Uoxkg/BKGcNd
gWEtKSe47WtqZfIkR2pxlrst6eGn7pOjHVc7Jn9aJ0TwO/BiBlSlF+TUL+oi
iLmkSmECmB8TNgU6CefHt2vKJhm7ghTIF627q/7XxoHXHqc03Os6Jq47px8w
cK0/cIH+SnNY1HV6hI0ru/dO/lMPos0xjvzeKB74kwFtJSncJlOeu6zoR8Rl
5v1GdOb6jZP9qPWHqmTTPnXDj+BC63Oj6XpPuz71lDVXzHR88o7zXG1n5+fH
tLChChB+IML40bTASi+M/gLAPUzb4/27+oaPC4G/Wt+4I3YnA0MhycSoyvcr
OpFhDiM92eckO8ZtZVoqxLjGRLkRn0ocoLyx8n9VFk1vMfO1fltvRILrYCwN
UWpYyS1aYsreViWJ+vL5fe+Mel8YZ9CkY4/QTpUrK6EIMNkqXIx0AZQVGGdP
1EOQwAKEnytjp1vOCTD8SgQPnZbbaq2kvypbpJ0bIJJzSv6YkNFRyWF5SuBs
Gze5JYyl9+4YeVhT3/WF/xLRaR0DSBApycUBVxdD3gaW94pO444W/CkSoadG
iMCFEJkpmZ0a5N9GaGNAqAmcfkw+NFxIohbqM9lCW2w/zwhiIdsl5Uh/sF6m
CL7X26+3xH7CsCmLwuw50yWIQZDnc66HrNgjlL6y8gxuPWWbIxSrnFD34TuR
JUZnGwwEsZDmMUf8IBB58KKtdW0GSGgHu3hKSw/7uhVtTCGeH8+WmNz03O10
jVxpm8NI5GupY7QvXRctEbqQP6sjb7CaM13JzBwX0diE8M3FXrLCWx1hCHEc
AA7dzPDDNEf0MOVFdqwcwEqEfq4y97Ud7J1UcJzppqwahJ3xmzM1F5GheZmp
1560fxX1NSCB2WoRsYEG0sp+d65Lm4giLbWdgsIb+/VNrJWW12ElxWFGBc3s
s4gSUy7VOcvc5z2f7C5baGAjYDRyIIS1+H9eEgT9XUwLohFyXyb6wW4dw0yU
lBxhABCHzJ83vg/R6C2zmuZTw+e5sUbm+1uGBDiitXS1lJYCCjKknoi6tXvb
h1b23oFF4cZc/cPj1kmMgc5rz7VC90CtXj0d+92WD55MeiDNwCUZtzRMw4ws
rdTWPBa2qa+desE/TT1mnVqX6m90ITDDh/VunDJtjbqeTwc/xKRLEJq2GiGu
jsHe8WeTEflHFA1qLKnCewhJuJqNOwXznD2Xsfze+H7xbThpXBB0fjjbYsIL
u3Muk2n6b+IJav10BijXNeIngCkaxxRBvy0jGKJih+hLAg3992R6H3HqBTQf
JpD4tMyAWNMd48wQCzSYwAcxbeMyJl6gWqHIf2Mh5ZJ2JiRURIxHmIBX5UbS
sTQzZ7WDVKgSmQolCa0b5/+b0Bx2mA1MxZyIDMIrv0HZouddT73b5W1p6rlT
hXHsOU7OCnI9ZI+GhO/3QSQFeG+7hPgQjRT70IknbYRwmJRENGX7AiOrW0XI
sWLxiwuYMzARhCACciYGi9nXU5z6m2prGNfX7zMTeFx6T01CmNKXseRCpCRl
AN1SfASY6p7iIUx5RnBql2YFeAJznx0FbdjTlr1GetWanQY2/HWBPdZpGU5u
Uqa8H8Jn2DqvK2UYjwM7orhed7QBqBQH5uESpMtvBqT7Qy7uFJeEJ/dfS4eA
pMLOWfetjTIgaLEWzK1wrny47Fxh8mO2A1+o3clruVSLiud3uv9Rv9YyeJ4b
XO2YAT5ECiAcfXT7dGO0NoIluk2Al/v2HsCvS4l49d+zVRsCqakNoxRi8m/X
Vc7lDv5WBhMPamjGQjJDzJY4f+D5MvpUCbOeOsSc3NwPifon8suRSeum/DBj
luBIVZbhX57ENsiEITbNDWXnJUfeQOC/meDBSC7Pcrmi4NhHZLZY0FqzU8F/
O0ak5Xg2LhBbe4RB6s2mz6jGMdL8m/qI9JrUNniFldk37vA99E7qq/IroSL8
iZeN4Ko/Ft6ot+kGDxb2HZLr+arBsUW4gvUO59RnLQhFlsABUVE6qNqZj6ST
nSUVglep2S98+WhLjww2Le52KRM4n24BtIOKcu5/2G73bPKB41RQ2U8fiZhU
k5Be6HO9owfQRnZ1ItTkIC2YwVptfwJ5ich4CarCWkfdVCIya0i3vr4rMugR
VQ7lOkJ+6T5SdLK3w6P6/2auauIJ+Td9hPWKD6VqQFqRqOHDo2MrLH4dulv3
l5fkitJCu895e8M9VSYZEV1YPMe8YgT4ABr1plSCdBWGh786Op6LwgYJwrs9
6U34FOmThSPJ2B5AiOP9KrUCVqN2oVNa8MfV2URAXL40BMQjiPc3WY7muXKI
dwd2o/HQg0zsUttBEB28nFkutLLS8DOdQbQtTtcqumbgk0BAU2cQLVH5BGUd
mhP0ICliD+6cRpnwZUi44TrEvHJymIV2wUag6r7WweNaME9xno2Ex41eIc9Y
HdBttFphWiox7LrWtuuDlE3dOJA+MBOJS4V7UKVudK9wK7Ga/DNmgdb7/N09
6IVufuSsM7zSzyEjvPNqxG1KH4kv3jIQoHh8hl82kuhJRM4Jp4fstbavVcjh
CCDphGIU2VKnMTVGj/ELcInwm+uFqIewVvxmyvw6EPsCH4nnPb0HwDT8NllE
9gTdcHlfC1zSQ8TzDJrSYxx6Ac0FpP2EjL1DXoP88et3nJ27qZ5GL/W9FftE
VY2K5aDuiqGU+JHNYNYVmtuCtmAnaHEM7frW/Pp8pOpd7M5mycILHBkHIGX5
+0/dNZasEPCiQAzStpFwRa1d2DF/Ml1LCyD3NwV14Y9/N6UtLcktWPqwcUS+
7MoIoPOXe7FIyEu+lzcKPI1xK+OOWPP5IvlQ31NGeWrWdmM8RkMeKfMJ+fp4
okPI7Z2AJxKyU38wxsPqPVdnntZN2PlOJHKRZ7NwpuZ3TnXTPvnAtaKqtV6T
iX2viUxx/5JrddzNEINAMqIvv0G9iy3ce7zBTM4w0Kl5Cj4OU9gISyDXW1Ln
WcIwSMEZIRIfcDIGF3saQu/WHS7zy+HvH7NsIS2wtwijr7tSkD3VfvSBbXhQ
XpFM3EjKJmZAFKnN1mkC9WWb+fMBbOQdh1BtdU99SpSXUrOewpplo83d3d4g
ZBUxHq7N2hGAPamp44Tgi2oB2zIXbT6oRI1zzLs+yKy5oc+/8iEX7M8KxRAZ
Bb8mo5dpJgDO+5/HX2C+I++eeDf1Vzkxyd7zKAOdfrkVM3FAnSWxDgpo22hF
S3DL964OvbqeAeiSNEWdtVN3CAPcRs2r7+18/8DH+rSCi/EuVAoZ14dQiIO5
7l/pnZZkFHj+uumIyWqUwJ8cOEUx6hyrVAcSFdD2T0PAXGUQHEO8rnezP1In
UxXX5xlUfR9+xve14hS7cgtEBP8wIRPq5FmuG0bc3G79/NoRgs3PabD4oEOM
YYgBRofItr4hVOIQj2PIj1HEVQzxE2q0DNDoXMHMYpXRV38kP3BvAIdJ+I0y
dR7goDXQCx/O3aOAftBCxFbNBCwmJu05Rhy+9hTaQz13jqNDKb/NeS8GkmP/
cXz1yxaJDBtzWA5ZPX0s7hQbsHFJGgDt4MnDKYT1fBQ+pi4hpP5jDVyvRifL
Ys6kA5c2gmEJjm9oGxu0Zk6cy9J2sq1WlGto2JPBfUbATVhIOKcAZ1djaQmW
/+lDtv0jLLdz8HIG7PzgjzWfwdFWu6HMaJ1Dfh0KC0Xf0l+ToZOOAg0XJPKR
yIzYkGWNc4ToO/hm5evk5UcU7eyukjyEnk4ulpJ7bVkerVuKrVOLepNA+dlG
q+neSfi9qM4IZY86q+F0lJAMhJv5YMSaALv4QKPG56+FL8aG9Sxdk/IyN3bg
vdYKymhFlRXvVO4pLQxmTdiGHCbvA7JFJAMOxhyOmrExUW9VoOu/HXEWnGdF
Xn1uO83Dh3Os9xp8CZ69BUSqyy84k+ar8+ISojf6s5aJWx23hyzL0VZRUIzX
6dRbFGFkoKtCY9I7nUUHaajdkNlaKfRf8I5ty0GJwDsISBQED9am4OA9sqdP
nevP08lsgEez5so8WYDnF3ogxSJ1OUsH1NniAWrZKTaCtzSNW40rAS3QNG/V
Yz9ULTmgENbeCJHEMH1R2d1+LSfoTTF5ljFoqYTQVhFmdW8XcXh0ANg5+6hP
UprN2LvPe20z1gni7r/wBgGMhglIaiCW2oLAr9KGPX2lRnkR62YRRXFFhpnf
BNa7vFzM5YOm5KmAKBWBj+4RDR86kxxQ1+9bJU2EwXCfMRAJGmKEk3+aUF9K
FocAT6kc//WepAZAN65CcXRiNq/UbU16qW5XivVwe8caIi0/44JhNGMFL71+
2nIDtgw2cd9be9bu9pQMyPB9Tl4Zv+T+g9Wgz0cSZN3F+WsBtLJc11QyAsgv
py6sgKfuUzQ0ISEe6Jl5n5TUG9D8/s9b5xdIdp39ttfgg2LScIumKANL06xJ
ULSnVuNBLBWBnwY/uXAzJ8CDmoW316jrsnBocTcI+uhv3IhoMJJMyJeiagVJ
04DdjZzE/6zZF+aNBmWXpM89NJHTYw7HKt5DDD54phRBZxSThBgQrGhbmOpR
3xUFz0jidt0GJjMaQJB+O1nRlvv6aEews6mWfKuFAmFHOa/6tA/9ZcHExTA8
bseOJcBWdhg/OtRMc5W5xGlAzJWznaRdLABoeEEAShJzFgwHiU0vYg73zqQr
HQ6pyQObzdDxDLWHdURz8umdsTp992oIxkWwYkeOykhah22C4VI+nvwXtNse
uY+rvImGa5jXhDGmfwwXVEekqbLys1fwXlbqkruM4xdRq5HPgAIPhWIjiyz5
CsCF5koF53u+7RzCucmtphY53tU21khDs37/BeEd0pzQAIoKLxc+LL6ASgcR
9zl+04FHXf5H9rKGwDFuFOLKxr6f4VUjOg6YmWLsg2JD+sO0TzE2ftlFKAu9
MS8R3WlyrL8Z2PtneykfiuP0wkByQS4WruZEkQfd6eV4pyaT5s0jM2gePKud
PHDenJ3hgj0tsEv5Mc62OZw/YVvf/SgQctl18bMWLA5fshyK/X5r84t44ohN
wegLkdAPMhWFX8bSUmumrXlMi1SMZmPp5FI87q6p17CDYI6q+E9Y1gvB3x2g
bDKgUuXWE+NPU3UW+4UepAA7Zo8p3DwJnpy1BhWIM5FhKIur90tJBws+nMDk
UcTpPopNnzFjb9tM5jleEWTwYcijVFXwRz6mkFTo0FAkMS+GEudYcGcbNTvq
YEvxmNfM0FSAn0TjDJTI3VYvhR2WzfbKn5rXfwMd1zxZwyIMaGjS9lWs2ntq
8pO4x9S5/B68AQduhvqpTSBOTlAaeI6TgF0kxmPxosoE+W1Wtm2P9aP+DLWF
lf6j9UZuv0e2UHb8L1P/dPCU7/5aUlN3CxlpIcnrRJM5ZrwLV4WzrBukwlxm
GnVaaYKCcdkzKD5+MxXudp5iRJcYBdH1Vq6yaoNqcq9axq1CwsTfWXqEYVRO
RGrB1a96TAywCrBTjRSejE3h8RZBNZYq1JPIwnRFpGtQPMBqPUt7l6lZmups
3FrZA5C5uRaMfnwp18Fw6EEffaJngu6jmuVy0lvFgoqlc9sfU7fEd4DirQSb
fuM1Dxmn1TJWL6sX8KNwVWuxe+0FxTNYELy2z/PwrmzyEatOm+qCZzePLP5s
4I2ARbrsx/09foA6UkstzIe0FylWdbiO6WOvHYvuy84t9hGHyWzBmSXMlThN
8ZN5CB+urZVh5HMFAYuWJEjmpLLsYXq7ZN4ueB7faeSIOKI2xQL9fH5LFJ7r
p6Z6vxAhlD29Nkq3+5Ta+v5ZheCEU5X9yVNenQKv3uxFqXOlVvH81Xb6Toc9
Me63bW7kvhq6iRg+FndkqG71MDq0Y/NlVwsVlk23gPJTil+jlycxeJEpaj8N
RGcMkLPJQcUuqslAALTFdjDuPA9q1/WQr/LpER7gmw+gcKub01brAisl+/5B
Bio7xYWCPOgSykhdqXHxXlBABrGfm+avhm7vsQCZvJ22FzYlNj2a8RBJPfiE
rWK9jbnA1D3F+Jp0nj1v0Cil0kgXXhElH62Mix9rMCBBtn/aG07m7qYXo8MH
XrutC8GQwvZ7HP50X+NxONpYq20tKvJr46oCOnIFnKRnkiDwezQEMadrT1zm
nImEBxhzyy9665fN4It3p10wyTyxeh21dOmZa55o3kirEDMQmzp5y796xlNk
aMOyEQd6BWIz0KUYQGCI/iHWhyyYZRLDKYsThkVsvrwxd2NMwvaxHL7Yktpq
qVT1h7V3Inff1m85AUMOI7s5/aaGR0KObDRRgDgHXoCsdIShveMZBgn/QZQd
vlvAtDae2W5M+f6wdO3Qu69VpWe5Zc04YckqzjxJzkzP+SvRzP6o6v4iCfJJ
qvHXeZiXCpMF2d+KwCop7e677QuQjYIOEdhzRU3tid0Vyktc0y7p4FMX4zwv
W4qovY6mS8VVEo2HNQCRYXqO4gvnnzrvGGb2oviLcPgmKR6QMPkaRYa2F6hf
DSePhXuNlu6laLtnTN0Dh7lvTgnUXtO/b9vLv0eFJhu3fL5kSTtYJ3EnIbBm
9fs1GL/6vYKl0TRAVXX/O6/GYSIUJ0jwhbLTQXiawYOhUM9EGo7i1JFtB4/U
za4beAkicK+LRx/WwY/aMLRc9XrebI1kAidckfZsLc1EK6a49mmb0Ymoba9A
PtuswG3pBz7X1Z3FDt3pwVJzFhe6BadyVmYx5jMn3RMGUpHAqOcXi7q38vWa
hAix4NrjsYSM/f0pOj+AESoFReJ5nNZC0n0dooKx76Ra3N/GQOUwWCW2dq5/
HgP/xbrcPLrHe9yBSOYHaJ3EFKyVq7ZlkabvHZg3wnwICHVMKvblfklEVd4Q
eX5T9q25T7+t6CZDFeO71krh/qjB1+X4vyp+BnD7FEkDsMgyaGHzQ8+JbqHH
KQJQIudtbddE2nn5txd6UFCaoC6bG/bLgfDs2diY6OGZN7MeKxWXhik+KH0p
O6rX14HrKLXbk4klw/6XNaHHc0GErWxDXDPik5fDc/A9MSIpdLHaCh5R6N1f
SN4TVtZcxDnY6WvCRLQV/qBUWSatcGfpCjp2ycdgc5c6Hzd6gxVFhDgRgg1h
n4hikJ9gSU8hlx62cFucwJd0G/koFhNH9B+xH3Tvvwb19X4NVu3F+q9hB7u0
chDv/iTqn+N7lgIUwwfwrCtK4IZ6IayyyzWvSoSJ6Z7Q6ncABTNkosuDRvlH
7Amb1SY0aGXwRlw8ggZtbhzbh2BrWb9IArZMa4jUYXk8a664w0UGI+n69bam
Adubxpl3W07euhivFCbFio6PhK3u0Wq2ko+CjS/VqQlEe2nDOQ1k86VNz15i
9/CGyncu9fB9967X3UBTnwyLGKZrsFjgDVaDY3dWiv6++GE5ZQEuI+ft0xUK
cbilkgZux8AHvyue6kyKOtJtdfOPqczg8T9usyEtE2QLklPgENbRV+3OHwLG
vaLD2yVZaepYDtM33/+ee9gsnS7nYsQa1+aFwXzwkKCAbdJYcT1w3yEojDro
KxduSJB+EK+q3e7dLp/XXV++kAYYwtNeZYdjumRZI+4GaqaSC6ImapdybhYW
R14n+YOBrNeyMsddcsc77SjjNl5KHVSx99VkD4Nuri/Gizx9vNHFgiEgtRmQ
B0nAkdtI+ADTsxInTTUH5TuvhjXOz/UfZq4H7zv14z9HN2rOSviphCrCWK4J
5lYImEoYLnU4uWMuUdROx0vfpjA2wW03WTAGeAlCObrESOKRWZvJHhnT7P+7
E/XWw//lR0/O4yNEMeQgS6Gg0S0wPJsUtpR9ba1yD6zPgNvETtFmvbw8amHJ
TaUrR+p+Q5+ttdSsaeGnPdRPV8iBZqVHtaCPYa1tHLGfmUkDsJAQulymnxqk
KFAWLhjAyMXHKKekQ8c2UFUoCqYqpB3pnKU7KN/DZA2rAJ38EpW+GqFAkS3S
9cj+xnapDlnr1e1qjnXYkStXFjhfZFRuwbmBbfSx4jGo8Qi/d3bl32f2nyvP
vlSNByKQs7Wt1VwsI4suQcIasQLdpF9e5Ur+lMuK1yG/ty4t9n1LYX/qE073
LSq2DJ+bpXuL/Q5+9dgDwhZKA9ni4JrTT1OEDSU4OdhCioFTkStTnTJJvAZy
AKqaOS+nZiO4bX1Za6xVY8CiLfMq3LvoGl0cKy/pjdsgVepmurSLK8oZaeH5
64AMTeAhow+cNeMzSMKRzNzYq1a/zqzD9swH5LRUc3oDH3eC5oUWKkdjFueO
GFeZtY3Al95fiHoUjUrmj2UxNP4OatleaxHJvEYaDU0xC/CrrvOIVnfSl+TF
YKG/hujpZCYEeA8r5Erwx41HNrkmw8ZTUtkq28vHZZonyaEpjvsBygg8kADV
41To1fOilhZm6zUdMs4zvJ/mLtqm8PMxuKxa+y7P6BkgioV8kACbSdl4m8kA
C4ZTI6fXsRuVasaOdCaN809GSFnJA2Q/d0VZwKTm3pxzFT5VLi2LDG96Uly4
vxBv2TxL4YrBlT9QOYSHk0X0cLCgoYw7CKOpNV3ATcu69E+On3JKObPZ7INn
o4bqXjuu+gkw/lVuOBqlFvyun+v4BxfWypSGo3l7lzIujbPu2y7k8rt1PxVj
Xg7XYtUSJccx+5dH4UkJOquDK9wjKmsGpbs1QLNIPGVlpWu2wIu1jXg/2Ujg
DnY8RB7oZFWbGD3G6GJOr4tp3ahjsNgNtNKLN7XDyMisEFLArBCYJE1DrzvF
815SiaoZaIA7+FtJbi86LgTVm0WfvbU/0V1syYswm9xG3m8oPY2/LH64PK2M
Co4g8V+yKhBWNI8ydV9wZJF/iK4j+MISVV323S8TJh6+1YefFWL2mj5p7ZvC
jb4H4G/l3sYw/oNpDQajiD65zgFTpXrys7RufLsLa6C3nUEZUlH4AE10ilvu
SWUit8foD5rObrkWkxzM2WKYTsdQvibOOIYF5nrogKnS6AcCV+imM+zqj/jL
8j6R7Kivo0+ZnSgoajBlh3MEwW0RC+Df+vvre/XlDjur8Y076T/OVqRkVYtm
2NEO1k+OeCxe5QuMHJhC5qmdY5I/8PsxmVobZKu9BcxRMmQf2JEeIcD9Vtz5
Fbw9omfTDu9yDRKZNB8CTN+0d9GJy7n3jmlbeWNo9+UKXaX0yjMtfofYUljA
LcQqAzq6pxRjXWdYu+GmilzPooGd1aOhM5b/a9XFNa8b06t2IjDFxXww3RZR
j2rU3QymlscFXyAxP6peVEeI8BU41HiP7AXlk6uvp5JXdX67Yo1fpd7giObu
LpZraQxQqT8p+DogF5BAca1xCRKUG9XG+HA+fEVCxbGWdYKV2uHIMtbN4f3X
TL6qxxgYVzyeIZynAO3XKCj2dSt6G8WnqjMByCW3H4kue+7MgxtJQe2NzY9x
vkaftkON5UG5oyqg7pYuqwt/2UTSB58PpRYkPSrOqf5M0/1bHG/NGogVFiG7
ZqlciU1YI/rObmDYmuuv1iqkSIoAMc0GXwL2VSsdoeYQ3p7SpsIzHQBxrIOA
3OhyTIbwHCAZD1X1qFwspbkDteboISIlI8XI7iqbTlaNqscSL8z+WUUwrfH0
M+VcejIwgFZdyDKyAODJXthQbO1yd54IGMSp0ZrAxHoFtHPXNGqibFl6rF7u
z/rGpD75TJ5r+cib3o6vuS5PdMoWRn54d+NvqYR7Din6Tz1ZKYezS6tL/idQ
e7bYIwGJYadlEyvwEtrdrxRcI8RJJpBdg/dRdPSpiH6iXLmuuBYbbE2RX5Ee
7kOcy6Eo7SSCx43nUZJYr4WgM1h47dGJ18ZUUeFUQIQMK6hjHqnl/g6bo+Kf
JZBEIQJTNQyPqcq7PEQAjnY5xxPsr+qs7rgh91j2zA75B88g4Y/JVRLRPzXr
wIgPbgtp58puIF7OE5FVGalLsqQ27Ff57vzqTc4dWoictJhOwvT63MlnV515
zRd2y3apE0UUGStTREINNYSB0unv/lcz1J8+YvaIhn5Ztn8GyZCfL5KB7Lc+
/+w5n/S53WMhoPqTaIOkK7+GkBTgN0T+yqJ0HqjQR5YnTK+6LMF7nmamSeFL
q71rWMcEat+Fdxs2fj4b/dl/fXIqp/DmoDVle918aKocP96J6XAzZdMywaPQ
tusi82cNXxik2KexLnTojUICL/zI+Irj1iiPfcTO4Mgia2t3VXpGXRPDPvO9
u0Hc7EZF6uNn/c65FNj8pw4fbPj8XpFFeOXAiVuM3RfV8BCjhYDE/IUt6MDo
APYTPuvIAmIof0j1xiXR/cxC4GZ09pxKAvRP4STWBqHOrSTFV7kws3jeg4M8
NBzAXaG5VFtqz4eDpYt6yHZaCde0iXUvzL8EHGZoQBF3T5/BBqHYariBIAaK
PlN1KI5kVPoq6INkzA+tkYxytaBgc4aopLL6i2xzR+JeDXegCNDR9FVH+wzG
2SafDFc/JEZtZ3Zprp1YVP3PDlrj2Npj63bpAHyoTwRk8sPvneEtYePa7IKs
TDHTgI+uE2/zL4KrP+S7mGlf+d3/4NwB1LUnw9HX6r3/W5y3MMYUqNWPZLAM
ZRrK2X10VG1Hkq2Dnbs41DJvtwaIotbNyZpZV8c9RTk6oSKC6IMlhsysTqo1
rE9Kg/u6xnHOdaywwWSaNUjVhsgBLuPAebeXJG4sn/YmKTfvd4YfyXjSzK+y
x/aGVeh/BSjPniUtiw51RIccj4Y1bTunidLMhaXtUG4SbtEWgxroc/4Rhy7+
asoFSrVsqMUbg9TrZxf4cl4aL1ay6vjuq3ANxwUndxpOUAX7V+H+dp/4Fzve
3QBYpRVQ4C25KXc5kx6SpEAXDkV5bXFf50dtYO7VbV5E8Xr32T5LLisuMjVJ
5NdG33Ig9wPRImRdwp5pqDF4PH76XJ0+dspUQendxdpsNjfIXwSP99QPRmTk
Q7X08Di2yLlyHUQUoJI5znRQ3tAjEC9FXts8h0UJ7xxQld4PfUKoB4md2Jv/
+rtHJDCCuaAweEDg9Fq5KZh+Rv/klzTOopeiw73jT7SBvkq0rsFvcS/AfiS9
rf/dbcMmwc3HVXYZ1+mJQTU8uyREmFvjcxHr5ZiilUuC2K0J7qf80o8TJkJn
VDfW0t9iS5pzfXgmDdd7sZBiEMRaQWZiIOKdFaH1S++EojDzFTtlssI7D6zh
lCWuNoknsdACQwkl1OQMx6ytALEd85r5GaZ1kUgx0Ex3dF/bm70vnXX0VJB7
1CgHlTDJOonMu2yeKOM4KnVtnRNRqMxd90QMjoarCfos824jQDAkPtgLH2YT
Gq5QX86qKBCBrEbFjyw4WyvltjFlGzUwb8Q+FhZWvtMOgffxr/CkO+1T2n6v
v61u1PqUH3p0xOnfujxmareKppEYU0ngE/WHIypFisu0vGcJ1SEmWKpfdcbk
m3xCj+kF28u9osJfRqhJNN9NyqzeusEK+p7s1eASRKZF0gkzaxqDYx8QoqBM
57cJffbChJh623yV1U5AFQscvYG3FrJOwFyB8wqmNX5Xu0X5OQEcgilRzw5J
n3NQuut8izAyrNkfSYeBTsZpetiSFGm0QjN4uRYTlLqmC9oyuUpaB7BNiIBY
gnmgHKdthGSCy/9sTzu7PKyohxnbTymZN2DkUfAdAIJaLiP9xdgLI5XnTtqA
PweAubfiZQeZp8ID9BwByKaUXEnIYvL5yYXiLty/Y4S/qlWny4h/q7p3wHAY
UK92HFJ3xZSixPaKOVBVZdOofn63OoAPNTBbnk4NhIONAb4mMh4zYSOHWrNJ
Yy0mjc16dlJLHRWufsSTi6G2tD3ObsEdKhXxt+xV8csXpAwSHFIdZKTQSxay
7T3YZCI8Klf9W50v9BQyShoy/+gfmDS6m1JgV7w4ZXF64Vpz3kCEodEOhYQK
s7cN3nRG1kqKbApuMFQPAhnPxMsEiBl1AobOEulLuwZ82pXqMZOuF//Vfvmk
pM0y9i/4XsKj1dTQjQN3oo6Bfq+jJ/bhKuTh60m2mtL0LNZTQ0FgxytehGSQ
5Ynzdi+I8XnRzdmgmMcyl3aCAsDfc6wa7G1odZWed15bGSe2rJyXUyLFFgOd
bMBH5uNDTqvRg0NlFLK1YdXIyEx/tqi/tDxzksJ0RlAv0gaXfuZHN/w+H/Bx
vCvkKDcJ8YZOmAi2fWEK4CjepxGPCSWztXNY4fVeA2CFMx0YqQVHeFuLmAce
FIC9J4gWOvRJyjKcEC3qKS06JaSx6mW5oa9xYhJA6kfdOdt65itSXqCz4+nW
9SO//z7vAtDzATvN80UvTWEv9Tn1tDgjVMA7xprsessj2jkOkm8fz7HPxF3b
ZtuBfySqgiYoNd4Fj1CkQUJj70GkgsrguQ955ZgNe2Ji/+77Wi9pmdjY811C
pT2OdpCXbaKMbe5ZGFmGCR1096/+oYlKkoO0BL33kVNKAwKisCwGitLbVF+y
BnWA8GUMYPmSxaoBlA1/uNd+DsWdtM8M5CJySLmZEFu76uxDHYxPvjqE2Jj/
h/0cp/unFmWmjaMDeq5QjdIfYIsvFtPBaBVaCH10wMR7ONRoyi2x3ZLAzboK
G6kXEvCJgcWC1UQevb0WIT7dM0WwYiftPXHiqzJWvSFGdQl0mqcfPOg0cGKU
YgrDtnK/7wx2Y0QPDpSHR9+AHIP7Lnaty/T9ecSv9V9RbhPJJRSC/OwXdHWO
Y4gR185P5yYEhOok6mjvQJ3+TfqImjdCpl1eNyulrprOZs+6rDIiR67/nw6c
UBPco7kZ9Ix4PiW2xY703OyieMoxMr266n9hGbVg65GNkxC3p+6YqT7fkSk2
Rkpe7XokXwwrgKWqiXCB9IWa9Ta3kFziNpq98t+SI2E+C8+draj29fKpu47p
A/Dv66zEFBEZcVtagSrCfvPjdLhbAs/tQu0Z5OcxpSL9KDo3HZIhZq5Jr9Df
qKOuSHLfB1z7kGojcZMlIx1q3u70HhwDOXNgbzSol0fwRw51eQwF5jb/NSZz
OTeZZrV9ESvgi+hW4HjE85bjCIYACEJifQX/r19OZ4/jXLfePpbEduwsapuu
+7NjYS3cE43JFbH5JTYoqpnj6B822DGjV9LTuAlBTtSAQ0TPDokOdZuO2zpk
uAHheiCTvnrrX9bqqneAqgtQA94HzPyjCEFSlKu4UPgxTuQWhNUjIRAVzF2J
uYtyZpux7GbJvbe1r8BKAlNJZuguBfRf6QDTdwHEP9+6g3bcHaqsHwSSqd7H
r2+ZlrezznZdD1mRzIU5H9XOpA9fZ6tbNdwi0KWC3diL4AZ4jTZJXGrR369i
7ZEqPSk8tTe3ZMWpo38RRRQTSd7xQEiDs2KstRB0PWJbevQUb2kxCOH2+Rlp
+lWNh7mmffB0o9NFVHxRY4ggfES47CmIMtCtsxCJwfwNdi+7BUCXetTs4o7M
z2dk11T6g1A6Ryt50y94UJ6mHkHSC2gYnyP4Tr1hP9JVVT5VMh2Ed+QRW+Re
3cwibE/0f7GLSnrdAe5prdrIcDYypYOn0uKXVQM6gg7ywq5Z89huOcPpWpFC
nkEikRhMnoUiMuDea/HikxVocz32SggEriC8UdTj6eWbaxkPK8ND2IAeYAaK
TfViNxfSaMCpXquOMaJ6ioPVcYDJVY52feqScfuKVtcEXzl0H5p0Uu5u5uqG
Zpx+kb9+zqlQGE6tHJ+DMoyYrp/l8fANdEb8IC7EQxqDZdxjC9+3jVoGgH5Y
wUYkEofvPzyM8skDM4Iual178RPu3AdvIfsnDNRf5t3jdVOi++d6wFmkMMWk
sdq5dHht93VW2Gmvq+9htbVlNQZBg8mTGh2pD0CMetrSXpWVQ7C55/ooJycJ
FI9fLG84kHeXIA2yfBwts3pWxZivT+EsKVH5bxZMvQOHEkZkFtpkLHNJw2zt
+X30gBuve7o07lExdkRRY0RwInK1X4RSpP1IyHNg9pNCU/cB67+Xhv0NgsCE
FbSDXe2iEKO5LuucpaYPOzKvrNNiYnJzqvN99gTnuURx8Oi2NUQg5NOBHyfy
YesdoovB9nl/c3soDusA+jieB3k2rX4QHjkskn9DtpQB79MTXM8twVu5iSc/
wk+nE30idIACc/b1mhFYyv6JG9Wjoll1e60VIi5Om3Bh4GqOqcUJ1Uef63k+
ehxJ1gWwMK6jeID/SBj6PJ0Z6DfEFAS1hXh6E2Qf+fnPe/DlENCRJE9jUG31
MZv5/rYFiiYWIW/w4qnQ8vOhI9jNfZC8YBCiBnmmHv+xuwm942QbT+dRsgPc
+aZDZs9Dizu/WUPzvotADjfkCYsW2plyt53Rkab1OyyMbVlW91UiKdz8h5ik
VDYd2eG7PuQ1eGeZdZER3Ual/dRBjeuLLTVzJHGNlKH/XJ3nnqkNaRHjZ9pt
+k3UfbjhwMpC991zpjJRc4m+Hnrto5/EkfEV14wPSzXR3Gdw/bIAjxGrNmRm
K0huSxTeN5Z+TLHbM8MyWjuiK2MNjKSVTC22m7gCF4lXCXICAkI9IHsHMSBC
SJjFtCMoQYO7ORZ+Wi6zQVGVeiXQV5+mEE11ZCY3U/naQeWxqJphkXyOiARa
gZBUzoTcDS1gi/925cjn1RI+CxLEdfy5BbSCuL3EGeiVfTr+RDTPUYBOdvIz
//gxzAlkOQiMNmmrUJWztIJU6v7YEijUh4c7ncu29RH8Eu6jf0DLiUqwFhAT
nPjxDeMhruZr2QuqO5GLD6Rsjw9CfRKFz/4W4sbN3u50cA1DbMaVWpsnYHGM
7L9Xf+jqKuy8RIOXWhmzaJgT4tXrFFbQ+2O1qE5JeUDcKQakNQi0jledu7PP
OqzA35W/HT9PtjyZOeFuFBPoR57RZnxc38o8f62nbQ1b4MGmsG5gM06Q9zg3
MW3e8/sPly4TsFnegCNy2ekK80nXdFYBqmLgmpsrghBMcOCEqTX8FXH9HvOg
TZfG5NHLp/4ssMTV/jS2LnC6A+Y6O3bwOcwkQ63QCZRXkHTPxLtFYJa8NpxN
la9wFZxGudOAKIj3N1b397kVnfAlOxlCmsMDgMqmp/QaRKWDSA3syFQHffHT
sYnzHYoAQ9lvcb/Kb6qQWlkPUaPr7Qo1t9WOVGiI5KqnybTEanptarixL6qa
yWsay94EERQJ8VcLhIigYGEPOI4HjQ/AlCzcE5vYr99fadfKliu8/en1+ATc
er4/05jzB9w2UlUiWacV9e+i2kTsX7O3Ka5P1G8WhArVR/msCeml9wLfCs+B
4usjrfqQixmiJLBiZNwyv710O8TDy3FH0RAzfKMtl8mXkBzgMkAsuT8Xkl86
xAlyxHws7qOMQuTI5fs0W5vXMW0Dwu7mmqbEdp0aUYmgJfwPt69VrgwFDde+
DfonhKXA/MYka/maGH2u1k/ouiiZ+B1HzL32vJf4AAUSlXNoklHTRLcZtoMY
IWGpPjZ5GfpQLuaDSqx8IHbOAf8M1s6iq1A512zdOO+yYjZD91ww8L8UXQ46
e9Yj9pxyqF3qfETJgu3hpnH/y8iZHDAyTXskrSFt5ElpOu3BpuMBm8TUvW0X
Zg2HifahG4XmH5cPzhFFo1Hcb7LHkWuxXo3kTk6NECBDVcqWCDpEtn7XjgaG
rJuNM3PYrgZuSYm6qU8TVR1i4p0l2vGlt9Qw+25lKKCL33lzJgc5IrQWDASE
+O8krYm1PY2v/PVXW8tQWXktznJI8aRFKZ/9E/WfdlKZSR8y5hvMmlExvMPc
BevM9NhQdnQJgp+MbMIbg/eLdA39fvGlSVo0UcGvxfHi2gdKnjY81jXwpyYO
1SaDo/+VLOxAHd2HrILL4x7uETtivkSbAYydT46qkv5IWGr9dNvfBwO2oSL0
dCHWVJvc/J8XLNi6vNwE+0fqLul0V9BCd7WoPRX6Z7ksbbSS3BGguxfJIOc9
LRvnMaZDeLMmPcaDG+Jj4lTvdTgKTaoz+ufH9F6EBJNk8aNEzK7vOePFL3EB
v/ClqIbrHyvvJmt/RAhy4yHNUfWRnb2rJ/CitoESKb/EeTkR3pP6zoRFXeo8
5OMSAWiObByIlqON9nMy+nMsOHqeshuKKHA4ADb38dv//7p7/2Oaj+ZhCGBj
J2VgXgVdgIWRVovkQOviRHYxa5gu/gLKRV3GpI7OTANgoTe+7jel6VtCi51t
vQkXNKMZjBju7uMFzuorHvHRxyZ4g+q1IbbkMicfLngzH4fNA6cfmiE3/i1m
bG3kf5gRk9HMxAQyAS+0ow57ZG8GwjLr0o1oQ4xt9CiWHabzG3V6ftkmTSdY
y+LGjt3KK6wp6DYjJ8A7aPeu9umQNUb63O4f3xrwrMcdKElzIoSMang++4Nz
Cj8/9BQm5lK8r1Bvxt/LvG+L/wmb181H+NljwkNOyo/e5VRYBrdESS6Oiuus
ee6NM/XFqzNsoUnga9Vxye9SwyMiwUMmKCcUrToxRohPbg1prpye/eCxJqLF
sqjRNZOQKE+QzFUzliEkQXa1+FG+TOqkxivKCSP3948H+fRVVLd4qkQP4R+N
kvKf33mg4yd5qKmErbuuOX8GS0zFXmXR5UrBUhOZ4lcs1eVUhpukJ8YcBkXu
HmDPI1TNZ2AvQ8TiYnbDNcMF6Pq0AMhn9DJBQ21hQBdiyD3hVrRHYC49zaCC
tVUUAj026JFwLYJMqQpqXzE3p73qZJwYzTiKkziQCeHMeseNqoUxjZroWNGu
ZUXH0Mlzp49EZQ98q1FTwaYV3MIkF0n712Zf3ilNTK6wJRseU1JBis0j4KvX
P+iNNeoT6EYR9QOn8bQSsIEsm+vO2pCl6TbagYDt8KWUoNrBmIaCIIVT4HOi
ZUcD46DU/HOYzkGo4kqkpPgOHg87GDyqh9TOkzyfwtnzJcjuL7ic1Hou9RKw
qyAXXYso7uPyVi/IL0xHXKyHDyQ7bzqdtXLI4ClbhWjARn/VCbQd2kDFYPMJ
WX6qvDMtQFDJ++Ludjjws1zK5Mh8/gurfQcF2UlXy7PV0tkFoAE3tp6PACoE
k+h6DIa6QchZOWM1hlf3+H7CBB4m16hxOi0Z8je0Uhiz1ugUQMo2d6DFSwFr
YjatkfCAHoYw89bFnxGj6aNZYWwWzzwkhQNl5k2pwI4GV8YVeizrPOYsxecO
Q4kuDj6TIrgzsF7A1+61WjWUOEqrooSNFYZ127SPcjbh2uQt345Pu6JI74/I
UQVFAYIQ9iYC1XYUWuJSlB+199898w9R6YeSuIYXypX/2oeYcqt129bcANhH
wFZ/h7qzP4PsnUX9nKTBWhQbC9efJmnZ2MayG0XcoUTItcvHjGkYyyq1bWq8
5taDjsTLL69XQvTy2dd+fyAYRCzBf0EgB7qluztHFzeYHwIs7S0DGGHPa4ZJ
l1bnjzRsEOa0N8l5BGYqnnSlfahbzTLVtotIjdUZ+tvtQv/DRo+0D7JwfkMQ
PSPWr2UN6obHZVQ9cWtu12GtYKhe03hSuCW0sK7gqS8qOgjbF6xRkKSiiV9k
tVXZZsY1e+142qOTcge/Wri661S2SL2wuRR2qFzEnjQQ8Xcffupn5ZlxAcgA
EKt3sYgrt+S4sYoj5xXLYLwoEor0s7D5B2/ytQYvQDfLWRMLFBMOqYbgm617
3M7jSOc0AH4lCSfpgkQ3F5Wc/fyY6sCgzgX1gcD4miCiCBKesCMrhV2GKCFd
lqpUG1iBrj49c8d5LEdL8wRFNw14QcYXf8RUTn3mA5VE2Es4dv8ou8L6lMkq
KkK6/xboqhQDAsfSDgSTTKcDkFB2r1HJSpWtuK0RZlBlnb/wAT7OSyLYzytR
I61qLZw5jWnXMbSxWZ5TD5xkUxKfYe8AYIOfSe5P06MydwiIl82Ze6ogNQ/X
6OpPID88vlP/3KSbfAnxoBKb6AgI3eHzlI+SBxqX+eGiAW+0sp2tZVH5oOZD
mPHqFwsF9TNSzp3CFnuobJv8TTe3Z6zckW6juoFee1EAmTtHinHOblRPXY6Y
xlJAQQw/3Ws5AXFJh2bDmrdJ92Of2vIGpcvvoH5MZLAsYTRZfkaEYsYDAzaK
aBnVejhmxjfsa3gkQSuD1p+9INIlFP4QF+k6E1OYLyUvNOnACJa0M8n4K9em
LwhD1zndl/GlKnd3p+knuGlMRfg2nIT9UpgPhIi6UsMms2Ze5cY3BHDwSVGL
MasqcJXEkm92xNJ0ha0OtVZQviKpkj90RAnXVv7Y+wlddcYaOy0OloRHnz88
xNDTUxgiX0uqRdT3g0PUsxnaGdGZfmQ+QJGWJK1oNqZA4aF5GN1ZFT/7CFng
lmFH0fyTFQqPGkKDWGN5Z+W1fDPtqLQs4d5IDZazCv+UsI4l+2eC43j2B3+Q
OarPViNAGHj2asC7bHvI3yUIpPbgvPBMcByvSDyNOOwHGasLNx4XVpELivN7
NxqQ4r1GBKgKsnz1W9R6l1YVHcYNd+pTBkkbiRJ+HgAnzJoFRGdDbCr7RyxT
Zx/lomR1fvGl4WENE6oJkSnt5OaVxHFGrqk1O2o9xb8s9qVXjW2UxMrWpZTO
xHUNYMOw/GDo5byWutSM+fDpd4FOduKhw2YS3LTUIpxc6XPKHKOr6DceRzVt
/ujokZQ0GcsqhL2V00vgljZ059JcQC/8qDENXRejgqnaQtBChxVaWsMgCmpL
F/f/TXLoYPxok9QNe21r9jxmJQw46JUJbBXJi79zzmxaEulzUC03vW4xHvpc
FYtqZT8J47fjKK1CtUtQyNSfG6Wyc1r9YxwQa+Mt3aUXEIuU+8EFQgxra86A
nb0gAd6RW3BX9OxgAmbVrlYwe9QFvPoRHMrSzxoFY1Tu1WSLrnHodLdLxpHe
x7+4eQBUakiWCMvwxGAHFqczZZihTxmBLc0v+juV6Jbbzw3X/+qlA5hdxGzZ
YTf4yK8mfu0QtbbiXQzoZt2ErcZDbXjBkyUGfWPTHeFGc2ee6rDV0al5DtEu
rZoYXCPzwQstKICMOv1/H3h/R4R5mlDo8mnSYG9vuAHKp1fylwRzDyybYrXd
/K3xGD0XzXm/PBCO35vxceXsKddtDd2ZLzv8HuhuP9ZVFw8FRAJgKNsbQoQJ
ntD1fPCgVR4oFyjjG+OycOj9ddZkHMg/Koad64rqS8nlPWA9lRkaJm4Xp4My
FulnZIo0XqDRNzs+W19JmNK/GGdeEn4v3ejAj5oiqPxR/PRJBkbsQ3G0sxQz
qyeNxYj24xQK3On0l7s2yNZUjm+dpHwfukPs38yfbCGvyJOvK65HHh16E46l
bwPrbcSdKzcpGyE+mPqt9QMyHXxXrQi02NrcfLpkpcWbui+ys7vj73kvTlre
JC8XJkN8QxBHn9V8FNBtq9Mj1bnvsuxgyHwYy7dUyl2t0dvFmkP6/a1VaZxC
zWhDJjxaIOtzrn/c21xj2YnoMLIHIVD81hken5044nPNOUXkdytR84YUnRRK
XPpqG1fU9ccsF4Czd9Ia2sOdia3PbrN6CPjDaL+0Xbs4FwdmhVDoUhbQeMJO
ApV0e9qvXD5dtZ2z9aq5oEaNf76TQ/1grMdGRqKIy7XB7eYwyfmb5mDoTBK6
sIQTCtmY3xFYjqlS1STxDJwN0uqCsIqldHnU40OK95riwBWp78n1movvj+oJ
BLK4CKiMdW4WnxJmwezGcD6IOuvce/Vnl3HE8jcYJWJF3m830ojXmZkcFDrt
ayYSwGO3SRmBrvUVBMVHk2E18PO8wFW+/effGgseiwFboLaKPb702o2wbCp5
g7eBSJkZVwCZPLeejg/xyui+ZI+ZeXYU/DNxt/NlbSpo3mAhA8VlOmOz/B50
KvOACkF0kGa3QEt+aWU1PMh+gDd+gi5TK5cZEI+978QJGfeAHDxoa8V30Or/
uH9hnnmFrfpd7n/H8BACyQ87s5lKwLWWYVNDq5goNqN/ySvTplfqX+Tu1jOk
th6+MLnVkJaQlXsW1s5S/FfWX12cv1JP5hVd1BNdphhIto9yWHET5/GjQiVt
B8b6fWPbo5z6LDmwcq/Y11lUrIsY0IikNVzxDpanzEUjCazU6kjnGbyQoTqD
37B7znD7xCKg24vspOhD3Ab5jYRWKFiFgzK3MtLke21bUeW4DODt4j+YQYyW
/9eKCqMtdWITH4qHZJWjuS9idSFPspvVsyqwT6oEBK4hjtXLFvPrB4fkw38e
4CHU/W449mWx1OZg8k1J0TsEcCMENPhhDftvgL0DVkIIrYrEDm+zQV5FriG0
QRVD0/g89Lemc8+1rTT6+AN1GxYDA4qmu1V1Zgphrl1n0zzFp8A9hWcCnfQb
Q3F0wH14guhPU0AfhybI5c/USfELNyyQYtvE7vmOOM73+oElHOjvaPS8ieBN
RbZ73iwhlCVhFEyat4G4O4s8Xp4dW/U/tx6midb5/DOwRYg45aKV1pngFzA+
sRyrcEM89TxvnAtDSHIzfWGkJP1Sh+mwykerZFVniTvFVxGoBQXdHLNbS0Ct
dgWJIlX36qJuc0nXqWYH3FFBGbJWhR0/lTobwssKpUjzpf07wyg7U2FSak/9
2LfxutWn7O7ilU4g872njXZ8DZRRhCCoahdhP9til1x59OZxrw2lNyu8Qi4i
L02EdNizyD+zcqCxNMAls1h1q4KWYFVdb6MD4IMQZmf+XdKfpXbusJ9nW+rn
mHlHTQedbt+AfQXsW3/95Gwjo9MOo6hdX4X5RmSe2DwjYZgR5RJ5VkrJnuos
UWvOHO33P9Fu6AQr0vuOkFdXJcs/INVr9KFMEM7+WXaX3VBz8D3vTjerZzfr
l5MbnJTRdlnCgG10UXgmwPbgBR1pubsmb1Z1S6ouO3xwa6Gyur9lsZZquWEy
gphwrD5C5Lm28v1YGOQjZlqendDPfapLp5DjxURUF0GQwCcUMWf4RnpTJoKM
KYFFvCQj/wiNcyHo2GfU/0XqRzU5aM5GgldwCzK/22pyb52hCahIy188HXW9
gG5kdsqwnvt2PJ/K210D9yWWnSv35G0Q+a8zq3j+iXZ9YZ/ZZJpYUMfkPwU2
iDx4GhwW3J50q4jhMn/ypS6bkICRf9r3U1CLaxjmK2iezONFDacXMA1ZGbEG
Qrm6DQi9loJwIknOr+lCnPRGmfoqduOmFWRT1JdC75Wclre+wYNrMpuMaBhI
XzaJ6ixxrnOGeTyQfQHoRmJSzoTT2n7wUraHmxA2zq3yiX/ThsX9sMrYG45M
BVgJDO0xTy0p6tPosnkjNSv6GxTuMsZjigsAMdnM60Ji6120ACDJ3MM106Ub
v2ymqYut8BvfUO/ClOLE+AQrSPwYdPG9T4Z2M20Yks9BmEJOK6Ur29TCD+P9
2moAtpLJmm/Uf98dtW73jUxb27etSmVuCeoegioXh5KNat+g/IE/jorZ28Ox
z+vo1nwy/rlsoqrQE2ZKtyv3OyZhkEnxCvhaq/UbGc2atfJe/TV1JRAn9Kf0
Z+cyubO0O0YchdG2ICKIOxC6FCxHKuS48BKC9LMutZrVBCgnMWLkhOvbGLBR
xokuqMWLs6jzbmZXInbTR2QPKq+1KcpClKb63pPRq54W9InkO+I4vCGGlpHI
23bqpqDVCeGWb7s9Yl4HpcrHjrOLfnVLkS8JaE1RqEaAsRYsChyFkG35mDjt
iEwYVzL4sBVKoz7g5LGd4SV0x5ZQr2xb8ZohGTUlkesTWfNAt+nCv/SMhAhy
YeDMT1RrnSlB6g7YoEQNrGU7AABEjCDF2TpbhcoSwkUZCbuiqbaejGodBmXk
PUp15o9hn75hj4T9g5yY2RleOe5wxdx04pylts+OMrWK5QIo1ouwMuKRCaUf
j00w5/vxgFS4INnj4G0r1eNEyD6xHG5E21sAK9LaZsMjGTxDGoRVmyc9YHs3
Z9rCk+KJi0j1lByYDi8Xr/yQHR1xod6tvvlxs9w//n0M7QpMj5Fht+4xXnHR
jbDIaMo+4slNLnS31J/lRxbBJSz+XpCG9Z7m/n4U8YEeR8WdelyfYsAKb5uA
o/87qSg7PbFdeq241utyGUxOAuJZNfDk7Cnc/OEt7dH7ZF65uotydrsPfAw4
jx5acKlmYk1ZvJJ9JzW/6y9U9w2rhBaoybmB/ALg8LCG0qcnIO0qSH5NeFaw
heBU9E7LmWCqSY2i6O8a2FXZvojH+tr4H4Pwy692KaU2pPnxSrkJyofqhCHV
95c4kbMfnVsb7CWQnD63LhjUKboteBJjI9IznEJZ1OAHEW+CWNp67lPWQlFn
RtBi7hBkC32BaH5Rzjt5TgfKVN4JBMEp60qRBbzADYpFQ/Z5oj1kaKsO5B7W
4niEfaNgQdAclU9CpESR9Sj1qKJtG0bAADMZwp6es3kBBRGUlZpM36INa8wi
OyhLXBBl5JjveS5MOcw1ieub6iVoSUgSX4RxBXHUg8VtfpOF8ZxB0EaXyazt
rmBKXo7xWcWW/oqavXe5Ur6Octa2nrFFlttf6/9PjkYkW7a+BsoaOI+Gdmj0
fP+dWKPHwwTwXDOB95tJloICrREut2LvoXWZD5erx6ExEdGhdwzdXBCp76fH
4McsD6Cqf6Kzg07g5YmzZAxU062xOlF/ToQ1na+A0IPl6fzqJYDzGQra/IeO
EZ2h8qJqcigAPTKKmyvVZqvJKiRoLQf54OgVVz41UvkX2KAgX9ppNJ/9xMm2
d6nb+6QQLqcwvkHXE3GOxKPkhZbNylGMU2zH2iv09aY817+z8EptaZR0hqKK
MowWRsghhzYMeS4XbX1U/Uag7cmsYws7xDrxuizG1+lJIA+dLk1vnJqOy/Pc
1FKX9N0pE9fWGLQxdg+5oOxYdDA16fW5tlkSmnGuX8QNEFpE2tf9GjvJJgDY
tiIHl7AqQj/QnctweNt4q5uwaBKBxOzsYWvfMDWVlWi0CzFkMWdc4nk9J+T0
8vfUVdL15Duj7YXESAWaeF0rnnH1POAY81t7XeHjeie4v8sMGOhWYx+/0WE7
C6fOOobAcbEyYTex7EpREAcVK+/n6G68UnQvxSpQ5UWJMmUy1GGzeqNdq3ts
HGOWg8/sm8M3/cJqYyZ+VoLKNEwHN6nqB00u0rhE0WCrEKAai+9GS8Vce9mm
+ZW8p1FhaZVlB0t3XifGi/15/UdhYv4R0Quv+BT2/h9bJ42V8J1FzR4HWqvo
/uH1CnOOiJDOkadsViw9UyqZnoTHzba6LAfeLdBmvIQ/2oESqjtbYk5IE8IA
i7WP0PhG/Ucc5UjIbY/xT8eU98X0CKLrVfSwZYUl/1LuLJkjQ8dMjt6g546c
SJVLeiiTeeDe2PNxPdS9i18LMFEvZr6vIiGMW1k44d/scUwraPEufKevdrJ1
eC0FcAQUVQcF126W4bArr6Q06eR0+FTimf4OXim7JJVkutYecrEOS9r3A8Pm
43W0LWC4ElcHOTwC7ljw658zpt7UmzdcP95RsSqhOv9e9Cws5HxXIaY0EifH
W4EdZ3sXCMSWnO+uvPdPEtyvzDbTDIcn3zVb1tzvCx2WnBHADM/06t7c1U8P
BKUlJiGuLdTZhRe+L2TZLPDAnJRfxZXsKYK9rv3n4rFy8YbgnEMgfUBpkDul
RUYM9UW+f6hJKvCSA4t06UaTmACPTIs3GXJaFX1K1I9BIR2/cZA0cUjDcGBN
98YjoyqLnhIsQlHgxeJ12wpL5ITYfMcGiF2jDRVjMf7w2sUBDeJ0ybzNFI3O
qfh2T4wJiQVXZ+DH8fIIpigDHnvpOmYXM1IG2QKKyCubHWnDVRIIlQ5XJnJs
kBqAIw5lCPoWQsFbWimt+kVcWNnNb68vvYMV3TP+vsAexU2ECYCL3N+hAqE1
1EbqO25a4tydms9YOK95uVAPi0M/fa7KqNUutLXR0Jus9wPvGaDH9oZW9fi4
R1zWtlLEjT5smgahgSD01ICEtxb8pswqxBlJH0XCWvoSjJEchel8PIzlzQX5
RyoYQFaWq5/kxzYN32EgO7FEy7bnLZZe6xtOIFw7Gz0vVHt5g6i2YIqb7Vhf
thICs26+5urlBci7tUPZj18RrvBQcHIC6r/kt++R0LPLxRhn85mH+X2gBYhQ
OsTS+sDnYy5RkA7G663BV0VqbjCz94gnKzUOn6VWJHQsl70y0IhBgg80U5ve
7dI91K603Dw3CWRDKEoRqCRvP6OF4CKKjAgwuBS22g/d4xm2ePtfLSrAbrSc
SnKD4z8ZisaWe7x3D03PbUljibZqYgArvSI3DO0l4iGT3QCMtcpHAevl73G8
PiGjAsv+lz0H/F4+Iyoic8L54/7PxHWUPAH3qZo9IJw2xImFhv6f0hWahh8u
6TRovGQYb6kT7E7ndxKf4BobEpnufORlL+JQRR8jWTZpqzN4lF5Hwo8Oejlt
lHMK1wya8J9OJfZo6PVIL2hPdT1Ml1c9t6Istqyfu/2i8Chhf+OXlY1dS1sX
FQNu1DfzC5qGltXHnhUJQka+gwxFVY2DTPzpQRQUum0swNhumQWOpDIOZWvs
frGTnIK4zJZFHWm8q+jSo7B4AKZcM14frfyk0BQD19LPShZi2Oqh6qi/1Ggw
Waw+MybgX35Ap0r19bRxL3ie1nAMAZ16AHaoebY0MrLwVFMfl2RksXqV22b5
C3htu1urSJeUrcaQYJmu8RfQ7e2cF7Clkx52sb1/R7urI1k1SSFwiSw4/fs4
18LaySGAsMU7vWG01tp6KqK9MhMojIen2AKan1Gi7So+japQcJJv8MrNJp+0
jBSkVt4If6neOqNiNjelLkyNC+BkujTerihMMU8LhOleeJic4eMQ8E4aXNAZ
x7p6kyMZlxbtcKj61okwCP0DKOvbMhfdzuAH/QHlXMdmbimE6Ye8YQrWEszx
rQke3MysjEFDboe+UNbDWxFIMws11QHYirMjwCDhQhLRQGY+I5xGchpyMRF4
0mZCLHR4KqVcyAixl7KZqAE4Gm5EaCaGg32Sg+rDvMZPNoo/bHzZnazoSCpK
HGV67qQfkIlf8eRUX3QQZQE4tDEi2r8rb9wFWVnMNbrxkEGNjcND1gqZTBUA
Uldsb1OPR/QZj8f2zANoMprZuexOl2oXPFlIik33mdZyURxOFmCBNHWk+Mf8
4VnjLYZkb3kjXKzWwNLwcB8JRPPLLu64jJFR1FQdb2ZgAV3YVgRBY2GZoEsM
ODE/4LGkXkAkYFS/D1X8w3DNsGnW5WA45Jt52l3Q5tTADmW9cFEESs0gS+dO
jCNEDPByHsMdJiAfmxOHuNR08TDWApbrG4nX6ACtUn2JEz78RoDHyCgmRSDP
h7LfCwuJk+Dxaa3kLXNOqtvSQ9IilqbURyzC8Bh/MwLGqN/b+Jz8+C6cib4p
9WFb8aX8q9AVV3TCIcFJwNS7PK9r6UuBNeveblP3hkHfJ+Dukssg/yOOj98b
kAeWAx7pY/agBBRtsjx41ItmN8Yy0OhO0GqDSmzX25NlYNd1g3WKU3v/HzgC
MArRYxEqLBLuZPw8nGbso13HpSgMP/Oc7tatVYBbtit2TB0pBEmmTYSjK9h0
fPvvPjpEX/Lmh3zUkgWfhd9U510hPeaQaqqp4UG9lICQTQCzMxvn22sWNe2H
zVmqAruMKZ+9W4Omo078SBDbRvtrOpnE1LPhw+zu/pH6fTamQb6zY5Ha78Bz
h58sCWI0vPph96AeYBC0kh5+oFy0/A8xu7dkMdpE9SkzSmqF8Nc1eBj88hFk
Ms9q3+RM0Catx9fWirWACJC05DEBvsZ0TLb7pfue9Eqwga8ySNuAVM6fq27v
9EfeO1S3NyK+I9eYyNTaJFix/lo6Ih9qTXF9JXP4GS44TJEftdpU3dt4AgZS
gZH9pXBhcKC2qs11S4NF3rqQ1sj0cdP/c7RXd/pm631TCBO+AQIICXz4eDBS
oMlQqe4nF9ByWr6UTDdlMW5Aw3ja2r2XgOq4cs3l//4L7Im1wryxeVz1/UHO
zcDSu2VZ61ZWW86zaYjn9ivWbP0vMKY9mXTry/xMEr8A8NyJJwXmoRykPdb+
dx8k7+l1ThnMWohvrGOHD090wII6luF0O66dyHWOBC9fi3+NqOxynfw5XgpU
GTQt+rJd1uQZEl9kp9LRNnG6e25r+tU6BbbqHB4zPApjVqm5c4k6feYhH++o
qyrDxlQEZKAlNxqPah+Ijljc8UkJijFNOT/0yWN32oFlavGzefQ93aiGMw3V
S0icWy0RWZSZzTbWwNStvlxCJljOKuvIvjhkMioFpfjUTgSGbZ+MaScy52Fy
svXRsMzb5ZXHF+ntCjYbbUSWuzSyJ0xCLFS2hKErcMyVfsktwbRMZ40yGgiG
QT8faOoDpDgqPIfyu3YHJN3oZIsh+R9y5a8GyzB7+Vz70vMW2Ln8UtFWTLEG
QRaim6WHMZFvlliPcCPm7LojQCyG2IEhhKGCL8tdYJgVxzhqWQ3NMx5MaPPI
fciQmxM29l9L8gM/1l8u7gqBbppkj9whQZ9u8c6Giv/GpeFWiqjhydHNiGov
Fn8jc7TDjW7tBGn7QgNJkSZ3H4fkKNs94R7TYgujgRcTIhZ8taFRzQhbNzAa
yc1NaLWJkmFQ3+IonHPbEG3wlTXkKjY9e/hcywkM4oJAhnQUrj1A1wTwA/m5
zRr4eBqUYFX/ItPb0Bmbwop526uYGeEnmlf8lKcCCVkxu1fnOHY05mXtAf1i
CGgnMgrNljNtVcudW87UKHZ5/m7DtCqRGRUaOMROsdnFL8SQSIKvJFw7BkCq
N9au3KHUhX6vQgmpkWpILgbRJO843PIETQqUVeGc9erWtyk6fYzgbj6oYmjJ
kY7FvOTgRJhowq3Ev4yth/nFrVyXeUXfdrNrRaTmvO/kNhXkT/9jbDm8BR04
FsawX8VKI0pfGxP1GMc+x4MRbu5tyo9tj47K6ymHv5Grxh+5ZVaT1zLodLty
aogyIhzM+IakaGnFNukXanvo5Amf5WVDdlP6jUX3Aqa/TkVYQlTLhBlj5XGI
k2j2msg977d1ElIsAUfo++TquWIkf7ez4QdjOcoQCgGs/XxvIaSrYXFDaNmo
O9ZZ+pdmOXyPjUonbPIuKLddPVJnfdEo1XE0DxCSPC4eWaZVi1OuZjbM42S6
GwYols6J68nVJ9csGD7kdxU0ZSoCMTQsmE57kJpziaPmIlvE1wSUvtXZ8XF0
u227CAgS6oO/5VrVzRA7KNOjw5vkCTxvYQBqIgVy/VPirl4Q88ai+ES8HrEG
OKlDSUjo36Pb+l0NVtPRBZMbfUighTplDdMSpf3hqM4RwEYFMvlLTEocIBJo
863fPIfG8aTgllaIHyZDJ4DteluG5aceDJ5HjV6H9HFE+JYvGwDSZAtfOINQ
59bfNL2PrHpLs0mGoYjYnhOtwkPhxhWomV5mkmhfg9dZf3wJTf7G417Qbk8b
ZedlW3BqSHWQdiKd9v/6iUerOmbuxDF8YqQVU084KcYMTEu5l6mSgwJAoY6t
+h2/kLcpt62Z8iQ8f8OctnxxxGBZP309HEv4PZu92xzYfnhGNXehZlzA/B2F
LE4khI6XUGS1hAZReBjAcS90dP+u+4XyP2BotLDXEiruoy3Dopcbj/GY+/tu
0Gvv8GjPSrqwDC5dHdJH2Vlb/cEElfLqipIeIUG/f8NcIAzOcXATqxjQZ7dM
yIHBNwY2KtMy8NSOOBozij74xPWK06fE90beGqggtQHRLCk3irxIVgfJFARY
akApgdCEA3gXxO81pJXHT3ZrwiQG4FeKOzUQDvmdvds85hAsrsO5w+Yi2ygl
zYjCZhE55dZtbn8j3TZux5Y4exMVigEpiB2UtkMqZgsze4USy3zKAq/tnlya
YF4L5AvjmMf3B+4YTxd3WR23h1pZtwn0XwVQK0xZwH4aoEEvXgeyJdGJiVTG
Rg2OuPItJ/C9Bw8IjK9V2dyqxzFCYL9DdCfEt7xr1Z5c/EKviYSpeplgLvfk
ojOZk6qw9iyXLMcOeLka7Vv9Ouvh3CYeedRnTElOd6ohLX3LVSIx0nmRfZEx
OQC8xkuUYllscQ7A9q4yZ/3CZ97iLEKfROqbEL/nzk8F27CXhLqpM8C424df
0lyT3Lre9L/+EysZ0upGYTJvkF9ojivX+BnmsDlQnmqk2y4Ws28akYgaz+uR
5P9ivIQX2DR6qlh011hNbcF/iPj+MRNIz9LAtOYfNbs2JgEDRCBBod7n3H8N
l3KxFB9EcpDX3xoxm7i5BlmV1GPCt6x2XaO6zjnPki0xpwPajV5s3GJpDsze
iYdebtV4wowX63Sw+2F35kc/zUH5G+ivj2cL6Gr6bvKaL7dDk2TMCirgg6BF
57lQRTJxU7SLGC5mYni+LY8YJgZRRA1lLcCdV8EAdPj/z6qLRasY/3QCMY6n
993yd1IyMlz6DniP9ziiRjDcoIrcHccTsK08g+Vp3iMkoZ0uWWh0jKKEpMVO
gKsaDOxCO9Axxs9V5lBTuL/p1fO1nxrHCZuGIJE/ddLWAAWTETrJpTmts1q2
Og9q+2dc12qVtlq6vzhWBI5ae1u62E1Xsxivi3vTEwXfKrLj+fuNq/It29V+
ZE2YMJcwq+gUaelb1NMK1OowF20+pP5dcv8Tuupx6jm0dcCV6IBHI30qJYX9
UnZ/YJWPpGhfmpOLOpoc94L8HwlQ0YZD+5769isTOgoEmo9TSWcrpjn0YXed
tXZ/s//uMn2d1FKGLb2eiB5WdFPfswzL7q8T4U08uwxoTw6s7MR+Ik0cJr52
abjdEeBSB3k40ISBhxZcCel61BO+ioVqpNDpgqMQGft9ZIjjgsHJLlhSDtff
mSpXyqc1e70ioz3H6m9ajnI4G9q7Ttyb2W2Kb58yOUuSpkXr9qRExJhAN1NT
7TlrbxVZZOte0ghTH9MrzR4nH809gcCpcZIRdct/BUmjNigkYhXvtIwsholQ
w14bdQTViwW8dYHqQa23S7p0W8iOD/I5Zf7mjQGssBRC/P1+7LahS6EBTAqN
L5dNVj9ZzlFd5PeQs/+hQURY3CWC5DyHhSehbkPXF8RLnXTytuGODTWbUV+Q
l2aiNfPbbBnZUXmty3ElPEvCcNtSFAOxbcEHmffh4q9AS6aZVIxOW32GAn3/
sW7k7MHHs4pOFCUnlcu6T5IXgAUwGTbVvXW7ZCOX5hkdItoBg4k4xLU0vooQ
frmHq6Cd2gJHu4dc+7OupEJqjsueWbnsOoRtAcp6g8waTuQdbZVCSxRHQXv3
0i2ORHJS0Em36t4HdR5vdgYa1Ndjbm6PpE/QIJjx/qcIBdpWx8ID7qdPKCep
pR1ue1Cr8vuo7fDimng1L9AAhDyQOA5lJl4X9v6MJOOhbvhnHhxQF4cbU21t
CtM/24bJHzHXAwJkBFQjoZj1DZX+IgjQqtOUOIH6GFraDUECaOx7GXXvfHs2
L/Z9f/bMMA0+uAEdDaiZT3a0Xv3JM6b3iKRJBKYtSrWybYyKANfQPj1XeNLD
haXU1X73JynHez0KkNiAgZl/hF6ZK+AXJAZ2snLMbG9V44/aK6MJv9pN3/u3
+GUnTSFROMpJaWiKsCT6Hix1BkyAH2n04nnkMIU5xNYnUoEqhsxBEx3ZYXQf
cufSO6bdmxqX8giT852lnMjdNz7iuNE9Ka57dMqmsj4n6ZVP4ZUBXzU7BBqS
pxvsiTX2QxjvuGzmPJBgKyC+rrQpBC1V56jaLNkC1ar/RlgMbxgoeojLzdYs
jipBCqmlqnP+REAeBqIqSoYDC4944cHU0IT9OjD5DqyFz4qfbAqj4WDVqcqG
T0ftb4RX77tUgH0bobWkkiaSnZUnT9MazeX2oFueuFl6wTBTde+OOaZc2R6+
jYleVgx1MmDNxI3Q5R0xYul6ERlLdHHscWv8iv8BmqEQVF9zahjxRX4Z5oQM
pIxVQN4sWWh0YreCiSlM9P1R/9rwo4HXG3eVu4VZD5N0G0jdSvX2Nne8WaJU
7wcTQgXo+sJ2byfFT5CXa2uKkwB2GKIpMzJmQXuOnB0eYiD5jUsAweOKLRxs
ou2qd4OHswb/9S9Xh9BCP9NnUkg9soSnBCytzyvrRacv4jsxbGp0SKIQwm9x
F7/yzLAy0LLY9miE7Q2caOfjIZi5zSI3vxaxJdk+GLK8YPMS/E/5VIHZgfEa
oLF/Uz68PydmDcPoGW87aPnTssiPDJwMvJYryvDtl3qsnbUPO0Y8NwN/+sF5
sRln10ACgqpeFxvwKgAhcXxz+OpkI/os36UGYqTXSWVMjGwHhSMeuSnZJ3zO
Kg4NFiqrostzBGQ+7Qjm5Tu8FdivFjJcU6mE3cTa2Y0UJhouDunbv6idpmmw
Nx2HpTWEy9OWnGYlphtq1Zw3tH4fbUcGs2GuTFWcfYsmfMD3uIqWJlZVrmRV
+8lCwe5MMaQxqbMJtpArxijTTYDA2KGLXaorOsEI8Q2trwL8fdndZ/3fuw0i
KCoy0/ooz5fKSpvHQ4o5YBLwmljOdXQUwnQNLkHbXmv3y7XmnMTeAJjRZprr
px+sawFDew58+8rYVPIm847eCnCWBY5NPqh0JQJ+uSNKSJ5DHMZeD8v73Da3
/Q50Q3SbrCVTnvrUNVX24Hfh6y+NldvdBINIGp/mfDnKfVXr8yTk3rI+Ulpv
yY3UMKZ1N3AbhsVb3ofl+eoRDd1YzVg+ua7CzQAeeSulr0NBwA6OwUeMdIuG
slRn5jPXNYheBoxDMtOU6zBAKnn5ZmAW4D9GCEmOkDJFalN6sdrIcNVpEgN9
dGYSiVGYsflyyw71cWMbwoakxoEtle41Z7/QtyY7el7PBHR5yuxSrc4Pc7+G
Hyfgr0nNGK82uMrb/qmtXN0WihTwQv5UFBrP2Jpc7r86d9T8Cr4CewD1kp/Y
uQg8NM5Q80Xl2vmFytSVlzhA9PIx1LYlyX6oDoIj6WtTQtewhGTIyJlD3NN2
UCKiStonYV5UqXNiGdKiMMWszDD28YKfSL1An0LCAREvA/JFX54gNqR+StvR
+U6V88aDDFT1TzSRsTcb7ARUPVCU8OoRM3wEc8frG5SrDqPsedzIqe7aJO3Y
fv7FWJ7Cj+G60M6MxmeqX5M0HvCW8B4aY5kdGuv/jILAYwyBSlqYL4hin7MS
/9WQ8ITphSmGieiVZ42f3ZjEOG0JkApJtJhuk+yCaZpTwziV0o7fspsoWC8I
iJIePT9CaRgLr7rtvUek0pcjqCI66kXhsKHdQPl45kzqSlujMrtANuA4zC7F
RvzivSa1rD69EZ0VC7bJHPNsBS3ylVnxMZT2lXS1+ZqE5k34GyFuSDeQAdZI
4O7QDMQH5X3VlDVTMEBLMqFCqzl4rBy+fx375Dmc3ODAA3nxnBSq7DiIupN5
Qt2QbJ3CaYddWSQk90gB39MSRLBErzHUZbTa6iiA0f9nWMgXzx68bthZaTwh
up0JPiQSFZ+r8jmNa+11/lWfQnBu+xNf/wloRTN81BiufhSCqUxgU4kv1Qun
WcgQHjYEcSChIzCH+FeAS1e4T1BR13uWg8sHavxUyunln3j6NLcUPCiNQTh+
DfGwlA0TzyyVYdssiEkYJiRKPmsBD1JvwB6UrTI5n1Up0c8BhQOSxEOXeGQj
6X+ZR82dHJ1nn7QANQtPPDUi9lbrJ6bnfK31WSiRIk4xwb/2+PuI16+VEtRI
1gw/WV6faOb/VXXClLS03tWjejJsol6hhrZyA6npcQD9XxDNz0nP3AONlkmj
HTVF4YJT6KsB3AInkYHuyjNnsAL/dcuEv9a/HFbflDqRLoiv8Sw5ktguR4DS
QTmEkg72gZ3aNzJG+83pcmGGBaLn8/837xR6dP4njpRGjcb+LGCFynWV5tHv
AuM2gP6LCq+TMTZI1KVHIsvcqabQ4is9cBxnCduo55QlTQkQqN33mzNYV/sW
25T+aWZ4sJBTXGytJ6V4XMv3aOAsT7SdNCgZOCeaFMJJQwD5u+d+Z2abqRiI
DZs+OgJHT0Odg4ih3k939U9tBCxpr25zNLgdGr/8gdW3r3qdyE+SdcC6+aqH
9UoneDAVlUDiZJAldCqFc9tIKBgeRPz+B4fy+0kOOw+vubRn8E0uS7D6t+/+
xZugAUQ8elOj/vLGJ+BQ6HXViZTmy/XG4STgtDesoSkbYl1Ea5/6J9rkfqei
9x00fA104NLfhE1ElA/4gws7bBosTzJpY3c/rMXtMh3sSG5e9uIaUZLl2/vs
WZ5UM2NWz95gcccLSEth4gWIcBKiQIES/W9xWXLJB4//DbuDvEYxtOXPr4u/
xt+McM+VkPsjth7uzAb1w58IeoNo3Z6Xoo7YQVNEB26SaT68DnPwx7xXJQ7j
i2t/FSNRZwSR25OwCowJ7XwVMdFMWqmqTODiPjjcms+2iSaoyJfvocva7T7R
UJ42IOnOjPpyygzkHvCJz7kUWB/Ir8QzSYgDc8rpKDKrTPM3rr5JsqwCNNOh
r6V7H9A+6VvrKncoPtBXXBve2ZhCFhqYDCiW9tqcARF8QH0eUF9BgtmZdIw/
EOzenolulVOkMbZQZt82M9KcD4XvOoMtAszle+LRcTioIM4R9H3eD1Ja3a8Z
LK2zqjDPN4oIrAA4QrFKnKApB9Raboyo8Ah4vHJcfOEjRY+LCljAxJNdZHQc
b8OBuOLkl51sCvMCBz4gRR/K9z3HPPxqPuW/SwS1XqUGP42Tt20Sq5i5yMrf
KP+PeUgmB6qEXjf2JFV9C3e6LL7GmYMEfYVUElSutwXWRd+cYn5r1spfwOGE
Qp+OvZWCy6CYp1hrb5CD5gyi7tfy/nPfL2Kf2T9Duuj9NE3KbZ1vQ6Ur+RXR
iKxBuHzIMl8y82YPNW0DblXbu+hNC0ojiJ2goJ0VMlB069QoXmLuJtWt0ky3
Jy54VeoLKZjfeetwDJSkiYlRkCDiRTp/EbHKihWiTfSjLZmDfELmbPUoJ963
TeVbc1L3RihAEIhsRokdjRsT4zVLHWnVULxCypcCoxM28TfnkBz9/CwIT8DL
OcwMFY0Mi4YjE6G2XYfGRcgGN/tfO0rcuTAUqqYXGyAnlqdOjujcQvEUE1Hj
OiU5fUT6DlZfRBZ9JB3Kmzm+tmM91kOu5hm2kbB9133xOQpB9RUAucHVOwiS
22YJFHGrUdxws/znqf0nSOoov26pFmCjeMwm6DrKgwdJeUiNmGUvGmdGDscq
Pclpu7V637k8dasD4yj2vFR+LqeHENLzrcu/eojpzELWwrYtGoXxC6JP75zW
+ekcnGMyT3E2HOk8UU/BzVV6bcZNw6MXbA3OCU5rBg7b7b9T4d9d+/rgGlN4
RJPGco5vq9UlKeUJNdA1ffZLKG+H+sXEC6BctvOf7EHijxonHR/trcWuSbaD
Vinv1AbnWax7oReVQgHm1dSbHMTJeXxfv1ESxwKpG+1Q7TSy289TO3bJWNQy
pVc7MpNO+l35v+pxEW94SzmnD1zKVxwTGQbJ3oFRUtzI9LdsYMGgF2MUFDGH
FCLdjaOf/E0SFzR0udS41SYqNauQmkOjQ+A9Q1OnI8S66gpH29aTT7JpSm4t
ebQ5XGiCNRal3KkmfW9ZKOeAJxLCsNYqj5nHk1PF9XkZ+OCc8bX11LzmQC5b
0AbKwqYfm3IS83jgybzXpWSbpug8nNe6+c9J/XkFDiwNggnW2UX5US2+Budc
kQOUr4DKATwaJEAz+FkO9wvgW/j1f2pzwMGR/vH9C84QzH8TvnxDLdDV+oOo
1NT007wCbNqwyCgrA7n4Vp0y/6TiLSorgYMraVSUy0c15yi5w1YTtIqo8zIG
4mKP3q2fuR88958Z9E91dYD1M71IRlPWxmtBLtCbVCTjW98+dmauBEa2f+ZR
4IGw/rFdJEXnoICM4Sa2mo9mQWlqgfPvlnijBxRA/0OrFjPlBWaXmJBlouGQ
Lr6vFbsXYEOhyPFgYRWp/K/pXYy7my5ICVPnuJL3jhe9coWrjCpEvoOngsSF
s0/9V2chabQjJmgEc3SU8KK50+wPIXLbBYTarE4McCCS9+91lgEtNn1TQwR0
aQwkL9sJz8XCxiFsZhI+fgKV39jDFe1zz8x3Fdh4Yz28hPx0EB6Oq1jx2g5Z
FqibzgAVjxDV1bUeu4fKapO9nNOqqYZKis4LJEICTQY+wxks/v9qrqptPbyp
JTgOimFamdOMrc9tnECQ3QDsQvhl95ONaTLukkwmJHTHhgtEZ62EScOiIrY8
IeHAC430BRKlumM+MmQpbbbSOe+/yYkbz073k6BdjIXQrixaMgKiQZj0EsTu
ioHm+ZvxPGMPBeqQNTTREUAQC2viYzc3pcse9ljZgJlAVOMx7Vk5daEoNdcO
k4fECd8W3vLyLMhtQK0oFTU+2zT4UXGtW5ehvA+kQ8XVCkFw0iz8lz07MeAQ
4NPm+eeqF8yUbfbU3ZQqOFnMfQACH8GXgaXJZmrOFhynYHB+zLhyq9KcdNBa
JoRtHuRMJy07Rc68aEcQsfNh7K24djOPeC2eQAoRnM1d1TmNWvpyHcm/Voyy
lciVNRD3mMWmARnQoRm8JBH7EQjGJk10FEL8JwFbBs9IRxtfxD8HLtXYbEkp
fkymy2c/aBlTJCa+GNMbvlWg/JYhxDQj+x+iJTPgktDhL42jLVI//r/bxoNt
LLdvg/GsTAOv40+nfR/7UfZ5ify4Gww/oNDAVdXB485EEEVrgjPIM+eTeKCY
nJJ6E+J66w5wbrnou2olavcGU4Iuck+NZVrLsTZPXUJHHCAnX6E6QYGMNjAd
Grvz69PqoOA9YUhC4O49acftbm3bGxwAA2omaycVg/iaYjUk4ia8PH61E3WC
u1ddp5amG4A634IHGEZfVI8SBlkEl2qc5WwJbsFhUARomPqdyIE9Ks9ukcif
xvZ+P4euuP4xlTgHEPkrDkvh5N8T97MTmc7MPz8YYfojwPIELaj12RvmqE+p
77Fc1fV91Pw6bT13+rNfT54Ep67fnd5DcrkDltK49L+Y9F3/quzxGfcYnsmi
yn1zGFpVvvkRxjkbwJSkd3KXzFOFlRmvbCPBj63T6hhd92LiLzDcn3Jak6Kr
yMFLLsizsV0AXmXrY8Jj0C4NTqLzP69Qw0tuypx6AVDoTkuF8oCiLY9OmNRd
OamwBoMOIVEh/AobhMGXpfLCwHLHrK8Ho2aAS2m6OJZEN5Xi5XZr/PFewVEb
FbqhxOPfu/MhIRiDgUt5nqaL/Rq8/N4NL32zPXVeWeuVdeKVOioGqYgfA3C/
xkDHZLCVh9WZLw80DIB+vma3U0c7giiBBVN/+rS5SGAonYn3hkaJQHlrkG3l
a4CXODeFl9Qr41Vr7FvvizNDmy7QBW5/7daPLy5ZWErygUM0WGIFOmjUB1Fd
Yaco/NYWDyTfU4FaBwhBV0jp6x7LzSPOGuB6THrq2rQSVZd3sGsgOmoZrqWx
9oQBSRuYF5V0ShO/MLeKaaeJV/HGLuFxjh4+5e+RrVUm4LOxDCCkCsQzbYfG
qGMyJJH02948kgEJNmKbXgHosn1mVhkODKKfU2tgkNXFjIvsoRHCJ+Z9Qrm1
UhMux8W5NMler97Q24vxdz67jyix0dYomDaaLtg9AtfUGG6lWz4Em0jnP/UV
iXutEhzjTV/SC10xaDJ6qeFCneRpzj4U1s9HyXXS4DLWZcuCiaRt8GB2aeLG
jYUTpOpKCbpIos0h3iRdbGOPptlHbTG9GOHrwUmOWibxewKTeXXa4HZlQgfL
wE/ii4RDMHjOBHqy3QahClGY8u3Fg8Dtv3UI2EE/VSfMC1afFQoyH/7WrXE+
GsKruES+GtFk7Yrf/CHz9Nypi5ynzFb7+1ohKQVuf1k4/shPIvbgDzCqqNKZ
H1ZrLC5eSvzSoGXqeBnTLWgQ4+Bjf017nMBG5aftlYV3ttpukceAE8DrQ2Jm
IXVXVOcU1gsKTvEONeJGCBRx4jOCdmX/Il7uercJkgGUiAK1hBrNonwdvo+U
jpaTRwPUEV6lHwlGbmedFMdYXe0MKs0kujUuP+BDn9y7a8lC1NCqDV71Zlhf
wT287fbEKFidRn5RR+DnpS3LmnX1GptWSz11su1JKBbkmRz8yR5yC4UAHsLX
20k5QZntM03xhck4gnRV71ZDZAc6jdCFZ44pY/KeFPH+DiZPuLfooHxfOMvm
H3nXdSuOsj6kER9e0MvCtppQyNnpHzvte16JBiieDPlKEr79VZFuTUhJhmht
xkMWn0k0QP1Yee00X5dhYjZorKOqyYu7acy+Ag8zHsGb27E+PATejU982nLA
S7TtwffQ4JOY1wt46wJEIFK2K8lilYFeBQdHp8Naw4UVbfFqqftpRepag6rM
Sf+mrvjxkSuo82vJ0788ajKYpoDASYP960npq+RBFtSVxGTSZMhan/dWzqSY
4dHFV2bpeGCfMPoTcwETt1OaSb84BQQBIFAiVLO38EsLCTrsHAQJtlm4FlqV
9OjIDeScKMTe0iaekxwmf2aPwCBx1NvfElSZ5NDbmj+ktwRk8UD12whnZRnL
FXlbVIe3G834Vkd6hE+b/TMhl1wA3t6HpNra+c4XZprtrPfF1O7E77G6aD1Z
Yg2fUAEAeOjo2kAAGHfNwVmrBz7h06waxUJr14kw6dWaY2EL2CbwLsGCmqGA
A7k5AzJsWZk+N6oItgLED2TR86eePPrn9WB0suR9//CT4LTOq+aPJy927rC8
vY4yxDFvKcKuAwcJya6sd4S1PywVe3FU4zq5silytm5NPH+2H8titaSqJ/WO
7zbY6TFCRmuxY9jpHZN5Ch2GjQ2kyAmkJdCPQmPrwj9nUEYqJuZN+mZ6gC3M
aMM0IBctHLtPdQfj4rDoapvrqmhKtkfaf7Zu54iCXGzyBDx0Ln6GsyccW8hv
iJdxlh1R4aqur+qwGrY2gsQ0+ZWhWT8IEmwfU6sHjhdjqLF/iP4wZethKLhl
Nu2m8Rm3HC+2SHaDso77tAux735MYPW6JwcbbWLDoSoqASmNV+0F+DQB1QRI
SaD7H0gDXcjtZqgA67Ks6DHatJVM7wXKXc98jIbtSQDctcaDIWPJbdFkO2qE
jK4VDn41mr/neoiyBPQndtWPux3Z2SbkxJ1gorInSy3DA7BmV34I+KDeI76K
mS6gNVQDzrZ4MqbNj/01OeUXk+popwq2eQmiVn57tQkIsaIiqMTSapPE1EGm
HMmphk0NJLrJ/nSVBEiMoErftSDlSBlOwqXEA6xfIt9XO5S8GTF0Tgcggcg2
5Ejdkhi1EOsGE79RXIXmdxcWvKBb0XeB0uEjtFxQER8ksp7tHqnHQT/5CQAJ
dHqLkuh6HZS+TeYWuIT/8PtIfUEyEIGq6EwwyrfE8Wks/WOem7xp1OrSbqK5
FwPBo1pIY+4ZzT8Ijje55MH+H6IIxgXXFbb51mlJ2zUudXHxm4fqKlNTb4uB
OkHIWeKz3aw9fEmTCWUm59R4PtXbP5pngVW47l6q0uY0LjOCStqfBmN0LXwZ
Bz7EY17Mwi832usaMxOQu+r2Z4gDWlEPggiU/T53948XSCg4RPcfQnyEiHpk
lT7x6Z2HyNIiIgxpMJ450CZ8EtkiE/ISp8//rJ+KNckdZSHXtC/NLxhAJaTx
b5GmpJ+6C+NRPwgEi6o+J+vAOc7cuWt6Vf03ICjRoez8+W+z8jIN0D4KUEYL
V85Cr3DfKYdQDlRJM1QXH097gXeXnBaNXPmjHeHhyspoJXkik4fnIbFMwKqU
RceXvPLN/zlQqJGk8vTn5l/32rM2a4jILsmfUhfni7VlommrFurimJsD3sF4
3Tcbb0nZEUjclPCTSggcWi3++dmopGZsW9X3GB/5XFoNM44PwxySoPrHr4gE
CY1kR81tCXiR2d1lsAW+fbFZ+M7pKBrb+oa1PL1yDHraGrCc3s6tpOpdKJKz
BGEWGl9x734XFefRMi4b5Wt/QjnuEWEMR53Qtnz6KA2tg3lAN8Kaqs3IQcAG
KH6wpdgWZOPnR6vDFTXJLqo0HnP/8XH9PB5u4eVnEwKMG0syrGCI39GXhT2R
zlAZUcQm3u2oNCj2D5QjZ7CslidwsoU2w8dwe0fzB1hbk8yQ0c4eoTsIP59i
3nnNuYHlt6/qRvpOdqOuRv6Bwpk0wP6vmIKL9ojC0iTpmJyj7w+rcVzs3zLM
z8EkQRu/qAzKHPT76DglEcmqB+RGJGQ5oWAyb93028VFzBMhteeASoBpzMz3
t146OUhaMBI2OxPwmb7XCFJCJe7zLFIaNrtc2q3PTa3QHclB+kphvvqHRNE6
dP2ZmsMRAx+aZXHYq+WM6tIAZZh0/lFauxBs1Q5VEpy7sqew1MOeWoA1GuUF
hQ3kb71S9K9cDNqI+ViCEYLLGH1aVwL9n6OzYLNi/4oIp61QTgmgOm7THIyb
4Dr0LQst8d4k9kGqCCkuIXlzfj8We4/8dQx8iEPvE02n3c1M+3wG/hemYluB
8vCUEA2avb6LKu/jGFnto8BgyNGatQ9SaQXgTEmXyjI4jLX7Y0GRb4GxyVZy
runaQ+fKKibgYyWBXl+D9pc4Z3ijT6Q7jkx2k7vTlDDkWdGEb5H6eG4riesk
53uA7l5UbVCoEUkvU+An3X7+gE1kQ9tX7jcOjTMsNi7mDSijGlRa0wL2P36Z
kdvBI3MIkAkKM7F1CqVwZMHHFyDdFgRMTlcrQcw8DFAIBvkLYBFnfFmmj6J/
kT7k4qj1XuQpWR7zi1+jWJK1Of02JqXsZZK/H0LhaubYyIXr9ir6QNUo6Jr3
J+cjMjT4EZyDSTJGYgYzPDkIyNqaHQymDQKd03ZriCyhCQCEh7KPQOIMzs4l
vLBuntKNsIzKqrhFmdzFgAEhGi06PyAbBbiC9KjtK11ZaYtnOSjMRgl5ShsG
nNJE3Vr8fLQJF8gT2ahj0zYGY9LhE5zwxcTo/vk/DmpxHKB5+7FAmBxytiQy
cR4ZRFmqBZDFkkQn+8ZE7MmxSh9vQzr17OdWd7Dg+1/ZKPRF1pxciWNGlsyb
mEs3eqDzBbsoBGWg7UYd95EuFgspR8M9ggqO1hlFV5AgWKqzFtr6t0KNqrEG
xB9Ybp7gR6emnnKvcxXEi60u9AgKIOsHX3RZnJFTslx1mw5xiBFgCa7K2jmP
RD+OQvStk4venrL+ynjfTAxOtHqBujFLQ552eNWlYCMoJmO2EIiAPbG0OL0Y
I/MOrOc/LXd3abdMVmLAvpBkO7vjOnTqI1PirSPNrPI6i38miTmm12Mtrjek
np8BHk3IkTnHchlhvZMP8ZmzvENUMA4YHqvFHpQdJGUUXbuRpyeGgRKzRdpb
MNq0uiprSocveUwlmh7f29nLhDeGN2e5PvjYc1zFUrL3wtWxZfZ76nCBJa0m
QS/vsixMDYrixbziXH48G+tjPQoZF24Y3t9G1i6JrkkIEiUwvSqaiqMl4xdn
d3ivq+ASTVyOOl0XYytQ3x/VaRNgh2jLtcSYXlOMO15B/HdV5Gv+qT709591
Xu3n++0nju6eKOTnHoXg92uyTD4OcWKiECzny/A6K8tioNVcmb66KjdO6sn7
ZhU7JGFrIvrQt1vx5+7M3rlBHQucqx5VOtjN4spOqsqY70Am+LPcYB3AvhlO
+ac4srykF9VncLaTKm5ft/S/+A/tHQmaLe8ngjNrshRmX/Esvx/7uqUM0MDS
7/x1gyaj4M3gL4ceTYP4p5mEW0NaJFzEPMHV8IAIIXFP8oyzQXXvC0yyun64
PX0KL9fPsQS4oGqhPjuOM/IBwCJJVbb2ty5v0+v3C1o+QlLRXsbXpN5qxFk+
9WK0PbKrIrDIjHkOb74uscblwYcL2Kx0J3Fq5ELrQr1tG5F76rE0enPUKNkK
7lXAr9JPicPMXOAjaAHgQNMo/WKh4hAjTny6Emifh4WB3smWBq14UXMjJbJY
/PP8fERjeGyWXrVs7/llVH+MefacfGzX1pmFdtcQxRRS4j/Qq9hpcKcluY3d
rIf5OZCsIvMWHwbjZbwIRYlXr0ItSWxW1bNcTa9HXanBxQjh1hR4p+RS19Ux
7or5i+h6EZ1ml0+8hrSbMSolKt94/EeajnDYRHWrxU8lrE5CPCBQxU7miDoI
YXhLUz/cM7rzIvjyR5Dhaswu4xXaZwWdAYBc1Kp0r/r0+l9CQw31N4VFSCBg
xKEaAIBvFnUEEY6i1kLtBTbMyp+fGUmaAMVHu+OQK2reppvCaV72MDhkwR0C
2yy/jLvHXlnAlZP85/Xkyl3NyhQ8d/tpnZYVvSpeWAKseAACbPA7FMjeHWZe
KtlaHwQ46nAeM77DrpKWFE/sargauHk24x0jomEoy850Ob0h+lQxs1sfLryZ
dvPK6rlWtDISAEINkP/fj418AwQ4g9waPcvT7tgilf2GCegV6qJ1bbB6R1L/
H946+I8vXSecrslC7V5vRuLQzHBv+XKkiwGAlLIWOhBog1BCuDdHOnlFGP6v
MTRA3uReGkiLmLnXz8+q5zbW+yUWDB74VIFUvrYg1kiIrBS4pZvH+yf1EY+p
nrPyNLtwRm6JR1iyvJKeJ3IfCBYn+eLtqj2c74W4B8WduFk8/Vs+6j26FNWi
XaZYubJoKMy8YC92VIhXwqKkd8QdU32NM9oxxs/le8XsCutWC6GMmAV0Ud6d
hNtlPvCxJGAQm/TVkfwBElm+ze5bCKPHAqLtB4xqQICpGfE6oHAlj2qbH5kP
+HQ+8aPU45Z6dGv2l+nsNY7sJp7idQEZhe99LiohQU0ogAzdoi+8hlW5FRMQ
/npCqbwtpjB6qEj7Km7uY+VHEHOjVBpuUQTpqgKpgcTiiXx+T61rm2upxTWW
QskggFNsh/GfSdMcSNL0Jmvw5icgDG2jzx+DIJTXWeJM6+zxCPjhBIm4q+we
3jOLsv0OEl6unE2Wvb94M3ZX28MoueufBRxKAsACYVlL2Q9KltlxegVWFQp3
jt2swbKej8Rod0GgeehJX/b0cOScOy7Q4MQujnpbnTNsdGb4Q6DxhkhTJJ09
qZ/KwsY+EKCdXPXEf6hqBSfzf+zfZKDmX4a2ki5yld756mQ31JsHBctuDvg7
W+scFYg+Mgu/KhzjUQ/a/cmI0/Tzt4ZNaJDkA8HyxcNUrLZnutxUwC3FoV1m
kip8fKB7Vc4D42tn2Wh7i+bFupkpph4xnBmapaQh8NQdYUj9fC0xq8sWYzR9
OrmhiNfGhXbxpAJSzjPUVi313kzgtEgAGxGoJFm6KQzq2C0MbuwSVcLFRHgo
wjmV0NNKCS2KEDnA6uJ7UVAXRn6APMNE6OmvlyOnjQPG4wfQ166UjrBONMsw
UmgyhrnLDb9aQ3zxv7+fHMS1WKxO88Za3pyA56ghdHaXGzz/tB+5+0AJLbwy
C+d9FRhJZUWUD63co/NSiehHF4TpXm2Lyfju81FN2RzNBDF0JA63QptP0RUY
HJXIvn4ckCelLSZ3SJxI7vsfoZcyBijfzru4sU+HJVv3RDkY29AS8KE3wSTg
1emNky9w9iCtAzzhihOBubvhw7os15aImSJo14o6B3S/ceGIgyPdDQjHQa0X
2wO0Yv4ATDiB2END4IwIP8uW2e20dPAyq14c4+ck/aD9A6hW8oiH+XNbSQGZ
kaVbI6KwEd4tyxu07gBFXSP+jUiiHwxUDXxWSZiCt/U1tFqORWI2ItmhdOoX
HyP+uwAyPRsWac02FH7ECqI9gvxGDHkTfdLF6U6cqTl1FcwZ1gUsLZ4pqYUW
iDebxgZGgUZFSmy9MlPjhWzTlj3pn7y2313CMT68PZWGQtXcUxq7xDPekKDJ
jNgWQQhFlVOq4PJuGs2G+1FRteXZoKoutCb3bWhtPPeo9keKAzMmvCDR0nZb
2LG58dqE56uF5WzMf5rYhyF3I6iOrggYv1VADJxJE1S7RDSnhF47kRxYVhu/
+knPZS1mYZ8GVRwXCRNZFwdfJyQODZBs68HM7ON/y1k+rlovMqf0M2uVJ47U
RXsSjxw3ULHJclA5iXpkdjafP/MephJF0lTKICV3sxaq2oTtUIgLIuHAm0G1
QYAIMZv+MXoRucfDzIuW7uear2fFuAo1W/NF5NNS60pYnSI7ZiqBqVBKs4Wn
MExfnSkVpSkWCl5vSXH+vq35+3Vpz4KmEjb+/gdprWpaM32lix0t2IanfvYa
65kvMvVjofbTFusTV0D2O3ZJfbj3+2X8eOHv7JpHvf5a3U3YFd+sN/ofHKtx
RrMHip7I1SXxBHy1z9dcnsWRBV3lhYXG5Co2xE4Dkb+4hAWvrmAUAHvoQ9VD
GNRqq8mEx/kpz4DnYRry4EhKB8GAjMXshHBV+RojatzK5kmpQ53c133JwuUx
qeHm0GqFc4SE84+ipbci/BovPvjkosPQFto6+LStcJZeiwSa8egD4p/+Mw3u
gAnQRU2akIzXmgbdVYWLyz6JkU2BMjw24R9i7XNRARu/iCF/ZpjXi3+uuhPP
lDN2uWrUxu1+qmQ3HybKGlLHvakp6z4KzM6Cw9gPu8Tn0hc62+C4sIXqLpG8
18Y4lNNPzTDsgdlrxxgMxZtGPcTu8rtRWArNqHzuv+RCkgJJNSq7VI8o5VXv
vZFC54F9VtQgc4GreoV2cZGgIOu7750dH0uNSn1JAf2rD4FAji+DeiepasQN
oKslS6mBNuiOyZVc+3wUB1wd9VL1z4tJdYCRNd4TG6V7G21oWWQ40nV6bMP/
5waO2TKLRZpcIUNU06BHbKXNxzzHUI6DWCyoGfTMPsh46uS8yHuv39+jRVl5
+AFNFS+bEARqI/VYGQTMBUUDBRntoU/ltefsvQA9kVlhGklW2qTi3VM2p6DM
/NoR6286QVOLIlwNMdY2VYXFbiCbigb+GbjPN6BJLBQ2PO4QCCHcKR0ywbd2
X3hVDRocge+zccC4SnEu6Tg8r9yNdCKDUyQ9LwAFH1XN46F3aRp8wDw8pOOJ
vFHKrZAbr8/9HwFoS1hjhuP4KNwfTRIAVDtQl7AcoZVHS+VEhG9PQYs/8Hm6
76yvST7KOfvLcTVSCwI5R2yzoquQlhJrknwHsQ8C4eMZvmWN1QFzy6UWluLD
AZxYq0CKpOPZ3miEYj7QsceGJfh362UzKareQbld9cmOEuQHrhxNmTSIv89q
1RKBanJyFTRZWhZPEq+7+LrZyEym/Vf+rwjevhzRG2aKDn1aCHr1XTe0owKo
VELFa/ozREEnJhzK6PPA6q/i5Qam+CfjuLJ4jrzQ4I1wy7HCApmNBmd3LppR
PjoscGVu6UUqbikejhRASxvDXqKl7CbDMWHhITkb/6tFLD/tvwaQxEzT97F1
9Ttr5nK5BVOkn0A6YfaC2B1gvq8SJymlnhzJDx9BDh6Ag0++grHwNlsgIOVk
OxIJGGsBmwI5BJfF8wEyVxwU7WLzdDvJzRAtxVBWsHnktvSNeZUeskTZOf5m
zsZDSB5SeM7cILozKK9UfhWOBwbITRFoa5VaMRwfqkggxSuWk1LNgQPnwYTf
7a+FxkZd0MHKZhvB3E0WgYU9/wuqlUhM9HTyoM29MJchoZtafnl/NGReHgVQ
41LCkSi0ePpsz9/8pZTakeeSnw3kISyY64zPU4/g8Nha9nhA0FKzlBCo6VRD
XD7QaUAScaSG16Bt4aFTMnSSDi0qdL2PYrzT5o8TJyFbC5NCv9p1BqnnLJCD
oufDG36xg9k18EBMybqQiXhi0TT2B9EYobz5LxIUIAgFu0OmlfJLM33QFCfh
B7U2WFGn4S3S9okiV4h/dshPI5gaswpSSQFhNNJsn9f1SvQonj2TkUFwvS38
I/2G0jn2LTMYMmvPtcvMjwFkUqlfoN5LgVTlEjqWBcGXb3HSDrra22PBxCqR
sboXNt/Kfx2qAEpl4lKwMctss4b44oogDxHhGJrvNlIdEBgGNg9w2Cqt4Au0
XpQ0oW7KoHsAZw4UH5Gt2sORRt5EXvdH3L6tjAp6PEgMSlvFAi/QIsQs0/xV
PKrw4xKuinvThwz74MWtQC3KmuzwRtu00JsVrzRug6JCATYnXPQxGluwWXE+
+7tvB7JF9qOoox887sExq50Hjibrp/DTOvUly33RjuYrUtLx4sLQUIYaOkKY
VY/QZJ4VHjrA96AzQlAFXMafaV1+qXqUr7ekK9eboGkFIure74pNReeyi/dU
Oi5QgWaKPhHE/cfi7fgozf1HmDoZmI/ZX73tj9ISWkB7/M78HodfPxc9zsuo
bmNk1MXxM1PDTeoqUeZRHqJQAoj8YYRa5JboqgpwUyG0KxlFOSD2AOsnAOWD
4ot0sSE6b8KP6ngj8eHI5OD9uvbHojSlo53VDYGKQyU09vLE4SdUnhe03cz9
Fvhhxyyjrd9lRtv8XY3Htvi4NS2eSAPXPN/Nzk+o5C4u51W5EX+J5hT3fvYy
0rvDbK7D8X31fiEa7f0euNMHqzK8xCSQ3Q52y7jvhfxZ97iV982/i2D+KkIp
Pwlhu+Hq1qHxog6zNQ+cExsrN9lHVCywOGLCBVtMHXQDpCgZJHr1W7ywkW1M
R8wdslve0Agqp7I+B/UX9x30xGV+hs6B4pocAdPdDxZJII4NiyHRrXg8O5Tv
f8Sbxdgh46hmAtRLvBdxK+ZaDuug2y2c9T0UvoyRbohBPKi/MqRe6Ba0NcPX
vfm5j4sdM8iwWuTToUBE8Q+K2TCgzhxiNRIhQVbgKLuD6ce9pIf3gC9dkraP
S6uQvvvpytGtG/YqWoQJ2G2oX+ob9W2CurR6iHM9vvaD7aIflS4g5l3qunWt
U+OVmZ/JBgcKgOyJg27ocDDKf+fqchEGhUzoOZOBOZA0RWp/SfBFKxE43Iiy
qHS7r5aSfCyei8kjzFTa4ZBG0Cpc540liX/qwAKDwWUTKiCW+Rj4fgXTIjrM
JEoZ6vXq+gtxYE1psHGG2TY/sZjrGGZ5FGStNPULTE0w1lH6w9Eogiudsr/I
h/AO/+Q0K6eCA0VPBpW2ybT3P5/QBrd3xjH15rNxUfkkBGJgiUMxHKZ98t70
czNhUK8hqVFvmN2Ksurt/XRPk3Wrehu4CiO0J9JU3SH/tdn3kJuJxq8feUQW
Rob1zrcoqg5+x06fnuSnkeRT/2qbbRmUCPgvcs2LfGzddgnlwG+ahQJgaZBw
MvZWzh0kB/xZ95UuNt117hxH79cGgIH8AixYOZ6pYLQuUiQLpcGlxRpl3qeo
UWYh8bnR7zQi14ocKXj7yLvkijqoXHTGSEZy0/9PoJ/+bRRVm+EtXqSrruI4
tA9E+EzG5RDT2DieAnxMFqtYTErw3gpciyf0BfTsBcIT7C01kBIoURQa1VLR
DExRbiq0/ukkUfOr/NbMRw8w8wWDYMYEniE3jbkJ3R5Mc0WTwzX98I0mfO7f
Aa8z7si7GGpdbP+bcDPwOiJYULcFZPghLfF38hWjKypYEdV0yTu9i/1t1ZKI
AL0MocLFfIrT3rXkPn2CW+AVUVWC1hKRI+haugRwY9KvmTGcg6GrR6pNwIZC
z4mEymbNCJ7IRZQ7/pOFaNNAZ1VeMuJyftZPA0+ezpe5k+R386oEFuaK9GUu
L/ByZkL+Zm8sD1tIjFyFklhF44E5oiZDqFnu5CAtgQGl12hLsqcXs6kjssOA
SdYV72Oy/DrGx/C5xf6Cp2AJYVRmuECJJemLhs9wsTt32aTqTomeN4e/T2Fj
SbVdVMPh+T+ZNXd5jx4G1dUUMOTbt9DJMLUiUFtm7IUI3qzn3meJasF0Sl/A
Cf5w9UJoIUkWgz8GzX5ZcAVoUt800n6fo5nMPRoDyIlB9t10b0x00WN7VmJm
Ei9rh6jnUMxYssxEW4zauj+Qo154EUGV0AJo+U0R0KUjk7id8xk5rfxYo7k/
OWWossppJmOGs/wDhCzhZmx9qzPXKBu8h/SZZv2CJBNdnbaKNZu1pdTjetTL
ORNezVF5rYy7vSLS3JnxLM27AIGdgOSmdbtXmp7Xls6fvHzSCVUN8O7YyJgh
MHWDt0pW4qkdOUaqGVAaTdwM2CoPuuMpBl58on/XzYWocQhetFH/d//xBUGV
Pro22hcMIdJe0Uhti7JscNxOheWlppfbx+ykwoMFZeMFEJK4Iez2g0+rhehE
wkplaclsQlamzHCmheqpZE7qK2cJm57IPYISAiXh55z/rhvhSvoYofkWc+bx
jyZFMh+DhJQ//I4QX4qrUcydWnKoZAiKInmduXCmN3d/77Z/Vye4XAnc3ojM
Mc7GrUIlLlaqU5ycVepI2uOriKVPfSOhsTITl/q0ml/guDIiC5OcMFxH4Vvy
tMlbKE4ORn3kwEUfsZwbgf7u8o/k6Edf48fegSYZRqf5kacAg5HwgRrhJPc4
k29qOGmN2f6QJUJKln5xnSCWXxhOyqoa9UX/xF/gOtckC7DFjERbAbrvXsMy
IwP/CPTip4K8k2eJBzP9QHddFKIjWn7NisroPvQKWn97WHTmxmiuW/0SBvSZ
8t2rfiN9j3GXubv0xLBUOHB7TsTSkt8I5nCgoTbCk/h53NWBrsiGlI7Cupu5
C2jy4PVdy2s4UmfPL5VjJXNVJlC2dNAsK/itI2EaKh+EOiSs/UE2DKmOtO6T
EEruCIpr6gb47kpGb3t8ITf4ZDFDdQgSi3X86BysfO1WLXI5KwcVJyP2dMtw
d/akj7uOQaMW+lPcqtQjo0s/t8KBLe20kWA72S6hsujuuDmrOhJM6TkIxsBW
vJ3S4+aR9Qcg/w1Iey7vZgrGlJGYb7aT1ZnFQxp79GWjgKf+D7IS9G5cx3ks
emJhkkIsv9W7n0Ao+fN/qnArqcdE9jgQwIfCo/YLGvg/p5meNyO/Q9GyHeoS
ykY5ulZMZHvfAUKDhZt9anWTTJ0oFmerJianC/mgfXMKoTLM/N2zQxqvzaJg
uGilmSzUOoX1zWSr44uKfY1Qn0czdVpCqpQ1wmg1cENFkSi59GnG/Uq9LPCg
4ATq6Otdqt0jbdvOTKMnMwy0ppjQf7KEwj4oOqinCQB4EFzosIu4CeBhhRQU
RpDb1lSARSwKriZl0pmidIKLdBKJl5ehmzPVTwrgQWH/MX32399ScsJj/zZQ
frzOU83GCR6xD+bwfeXtmU3UJ6X3cPMNzMdBXxlb1Hq2jiTRgBa6fp0ttcrJ
xHDc1QafhWB70tvSwj4d55Z10NTa3iKnbkNYAwy/zeJJ4zHE4yQyrGMBkfnm
d6hiagJAaB4LuCVQZ2YxLABnr7xaqIrE86A7GkhVAF0tdOM0HJUN5FsgOLEg
vLH+OF0HazKmfC+rONdfw4m6qn33YrnxUeS5TViUK32cUQcaYTzLMhszMjF9
f9Xl2rBFYasuYEPVsHaQ9X4o+EmDy7X7ZgBj8imHBLDWBQf8Epvp2oGfgdCE
0xecOys8QuBHrhTX71W2n2YZTCi9eIyvYwKiSM5IlHQkccrzjaMyC7tA+yEH
/vv5rTiHNG2+H1HDr/SnguXrSID6c5frDMNN2aBJXN3MjhSPYHP3kqLR48OF
d9JAySsliqfkmRheTTNZ7ND2HTbk9rpdEmQln6Y5O0jQdnjcaDj1BBIkNqaj
7mDxYz2xkkMI8vcV9x835LYaraX17G7oVQXUcFk/4fquC/R2Yc7yzKHUsKJ0
Zd7l/Pd5150XBRtVFS4+lEmRDv1DGp6wWUDvD+TcGkMZW6VfYvrRBLzhg8kd
Idcx2fKj4XR/SZrxigSlSwGQRm2bnK/m2Vub+tjKGKAM+VuJPjD1em09Ifnp
sx4PAb601VQgh5yBZZ04M/eOXxP0wTKLvynTAz0B6e8k3lobSrzrweZ7bChU
F5nTa2/WlVubKA9aIe85fmXaZM3JxMRN+EiWtmr2wwX+yz8nRs3blvF9x0eB
RbmMX9pPj7VQ9BkeEOH7n0eao1tCw3EApATugZA07qVPZl4qs3s/GPV5RuR3
2PPPF3fISjR3C96uMY4Ytka7Doyi6Dldbg+sXyFDEvqWsCt9nRAlbCUuNv2L
S7KGIMOe3fSaIqGP+pDvLVT/yDbL9MWeaCuyuMs57BrFt7q9TG1Duc3amHSP
4NMEMWmtZ6nxNTrp2WCYSiKhibwMFTdAwWrp/DgKP4FYBTf9xxBXdmi420Jz
Yw/+eLaHjEXIKyYF1rMZmdtGjtihVj5tL3IT2wNzpecjOReSzSA8Eq2N9wVn
fC7bDNaouaTOhJDJ4162aydH0aIWeEIHRCAK1VHOrMCGdBaZQWyvzmzV/ibR
wH8aiG2uv/QzDLFfSh/r09v3We9GLN+vEYkAh35iQS4q1wm8yjtzX6ds/ZHn
4gvl4bnIA/B87Ye70WK7IZ7eBDu7yYAP30MwMmIH39FpAOIitB+s0EQ4fTZL
rAejm87u1SmxGXhc1VHvlfyo4eWFHSSXxyXFOQf/YGvQwE/NFZLulSnmDlLH
PJcrh2Iw4eOkDZwY4aDcirc5N1w/6cdlhJbLKZ9FhVQJmbtcplvTAy1qZF9J
qncAptZvdk/4n6F1WJbJRlYUDrGb9D+QiQ6kgScKXLxPxGtFxWtfwSgFrz6C
69yq5SCoKCo1xDCikPwafpRgzNeUT5YnnFPoG7IpsLxpppnFVyFMHhQHnWUT
Bnyp7dOj/6XNfZanZFKxcMMVNkSU+SWf8buAMfMXZp6XTi36W4zjNTWJdPua
gJLdNA3ILDxsRQ5l3uuUvZtmlKtJymvWpjn+i1WzJkjEgMEwFZYrogU+GOBi
qBhnfM+otTXgYromClHjXno/0W1eOvyIRTA6UKrzEBM8kisH5hsYY6n2IuY+
SExW5AJ7HtbWJYAMlmYMagWdAWMmosNFCeWOrWSkVzO5dGidL4brtQkXpe5t
JVly4SLl8iF4/Bk9+0YZNM8CPQ8NiTEgcRZUA73ZoHpc1Lk1IAlooI7EAlqh
sPBxtgEYpTtvYpC2TqKEYM8qKwfc6WMtUJfTHctsnZPVFH0KZPgFPf97hmcq
yxD4TzSw2VLza2E33hOgioGZprpUSemvAMQDHTD/CsvxGKRat0z7rmqYaHrG
V4wsdS2vXIPcZQYwkgWge1Jr7w6vdi4+JrID0Cko4Bb1yVbPlz3fAGIe0U1v
PKxIv3TzoJV6rNjinMjd5Hsbve2SHRznxdA98OK0q474rt83C2MrN0ma8q80
ktYHMY6QEJbariL8+VUvUSSNPST921LWhrkS8nBoyt+ddW0pqK+D47BdCvgk
qRGHZSpD5MkXWhwRRYZjI1crmmyF9Asz/jmJYfxpfuZPsmVMvWoeQPzXAASP
dTcXPVkuMooUilP8YxB9u5zHrCXYbVLDKjTDxlxq4eynyq6/mt/amejVk8ua
qmP9GeHmsN+GhHygTCCp1LlnCtLhSHGkQWAVxgkQc7unWhAb3wXg7qrW623H
vqg7Smdxzy1Cn9s8s6Z9q0fce/GMily526Sq0xMYacguVnO5eDrwLHFonQ7Z
Wg0+gzZPMIJAyNEWVZJMYJe/9TLCEEP/5MLdLrNt9hJbs5PLh8Hgv8c6EfYk
J23MpOP83P1b6hWo1zYHs4zM8qh2hzkV+9P2ALm0L9raiabXeQA+N48gY/1s
IZFXw15/Z0Fa4HOM15+JQ9no3BbxRAaaJJR8DxoKivu7oRWRqU1wf2H/ADTA
540CTktVdtb6jmktFhWdtj2cdD8zPwDvAw2G8ZxyU4X9FbGBC6wdsN5Uk9Y8
WLJH2N5rnrLP9uMuDfdoulDTm3Cde799JClabTb1syz8nT1VZSwCOwyI7HzQ
3N3gjiPtKrIGsE7tnclf+w71Y2vsO/VzqzvjyIdpLYSQeiahY9di2BPfCsxa
OQHiG2kMPpNiC4W9I96P4y5B79GnPUyZhXvwS7OS0FPo0mBxMyL8bk8NoeXp
qD8CxJrbCjMueADUPXKpIoUUf7hZMBHmbKeoMMS4J5k0uCU4lerXL+6bnH+i
sP9YvTA2oVK56al3uPgAIfrJtKkSAbR8n62mMYpTLwLWIbtjgxDUU9NTdpFQ
p7UIWKy26jEG4DQ0FZtzUoHrWcMfDUdpTK0Q8vY9BIiZjG0nD3tS4gbmCgsK
9m15Qs96EoFIijkEI5RbowFrfH1YGIifbSZuGOwO+/cVdGpdDNMRvz4zZuSO
4VDykBCftc53ejwv5UUZin5HNcrUoGjGK4qVbvwaczg7J+Xl9Fzn1gz01gSw
13zlrucs64wB3qqYpn9IQWxPJ35wYkGbAwp3wScX25vs1QOGpDR/UEZxTc5x
lvLJrcgVwcta49bpz5QmgyGasEuA+ybNdFtZOpcU++Ljgq1sHnBUEF5+j+X+
h1PjhQRTdBGYUuJ9OmC2tSKNNoX22eRZ/pe6PkLhbpUPQ7/deFjWnP9bFCTj
Xn8RH8kuKzOELv0E/SgNeYB9VnZ0B7zAQrXiWaDpjx1IkmQjC/uJ6koNV0R9
8ZVLGI6LjQQ1ASZwKJ0tSBE3Fa21p9ldrGCUnLX3rb+tc+z+kPKsT3b0BrYN
Ne4Yz5zusGP9XHUNmkE/LDfwU0NRNYEb13MBxitrm8XEAYQegvj/YgvRvDPm
3ZFBdR9qLTXIy9eqU8J1FUyHNU92DaWexVwnvIkkNcrTtckyWwI2IGPnKQ4S
26LXUfO4JbVHj2iJE9/xkK3LD2LJExYN/g2UbeB6LQmzXXnsMhGZrM4emqxE
NEv/Hri3bDnC05upgD3XLDbDoV6LxowqGLjuE+53YeKMIajfRLUJ1jpZJ0Ng
deF3p+5qZlYpWMgwTujUWVxlDAJjQu0Ikdp6niBu1MPvEgs82lGVL5tkP7XP
T90Ld9StIsM51SIsTYOADBJTKXlMaSXkbmculuAcACcFyJ5XIg9UJCdSBln/
uO/jKvzEAtv3O5FOJrOMxFVwmYVG2G4wYgNlmL8NgqoOVgyBz5d7G3xKGizu
/dGcAUv/Rvb2Ck6BDi1E6ddX+tHguZpsHFPmpgdLR2q+hm1mjz/BHSQhjgq9
2X+bbV1mzcJxGsqTdR//8noz9PkPbYtMiDQBgLbhqSV/JWou9IJmWJMwY7RD
ISQkOsPfqT9FTVzUosMWH1AhGGCngG27nljMR0/PPF5zDKPYdVkyvC7x5hPi
w9uJmgpu5WEACxsSTWvomZmsh10JIU7IxvylB5Vwp9m5c37xN3JjAIF/g+fD
fEnB9JLda+mPxPmXZTo4pucAYCuYC17jc6AcM0ZCP04vCacjXs4k9cAiLUbg
Aip4lar6lq25Y5rufSIQWaWsATT1Fc+E4omXytl5hj/tMy4Z7GLFIMeL0ZAf
MtYGddefxfnvUhIXWcpNGTVqWYWqDBknolsTYn5Myt8cVCCpcllLxALs1nc0
Gmf5OF7cKIRiYLNLdlfkzhnZsVAzaMN+4Mc+HpeginXRdQVbgEPAq1tjhzuR
JhkLTYdBuBfCiveNVnOWg279GOSWJ6aDZFYhKyE5Vfh2WfetHUzj6hbges6f
ImTIjfz/1U9WoI3JYWGHR4o3SQpPyux0meJPRfwSRUn8zMy9zIt+hCNqXiMc
L15kaQcZUGkvUUc7alCd6/CEuGgRn6mg7IjKSLHhZOt+ftgTnXoWXUraUCq4
JZMh66sr0wpe0qRS+bcLqNTnRlWQu+irMEuWhcKNbsQjXoEBnHDrg7jSSvHy
opReun5zdPvYdT1yZGKje753EYbFcztfQQ+m2wnHMM66njRU0bgKPOFRq80b
KzYdoV1/FC13fFpqD83EFNwqyglHMOPgRpln1kn9EipvDx0G7sRl3q/g3EoB
SQ2FxFrqEp9Ofk1Je0U6rcZlmq0Td98eVWBYwkeo/9ZFgHdFGJ4y0WlPnSWk
CWIHttd/YpcslVVlgAchbd0/ldPg19lKnfD+MqrZj7nniGLGLj7MqIFtoB5V
uEG5Iqkw6zi+3zPkMbJYBxeXTNmYQhJpKAe0LS0tDgNTdfOkGGHYdG+oucuo
gbi6J5nnkPvafbckAXwV9C+d/2Krx8Vr47wObGJ2iOzL81rVHnpqw1ba2dgS
jkrV+KCfljpunfOZcMBu92eURhiL1nT7vq2ybE4xdlKNzqnVPQf3jOQWUG1u
qo+CAOk/XIWOWsvkyE6Lcas6QO4STRrWp6d6fxXeVwl8KLaOUeZUVJ2RD7K6
3fJlCYDvvT+tYmDoxT1OQAD1FaT3LyGPnEQVWHL6yiKAo9g1YfsIi3lvfT0O
Z6SERB1rs4jXjsIDpMWto8MK3im/gtm6UUC0lE+TLqOxNV8Adv3kZZV35SZs
mormosnu/B4KUBc6xCVkzqMXE487j3vn/wonoyndus8HPcEPtL3eifzOASV0
NjJ2T1CNF/56pTQ4AkDqHGFWRZ7dRlWDxG9DWb38OC8z8cAr3jySrjM/5ArO
HADzX77TPq2uxzKsgcvTkFxRM9h10dPg8HbG5UQhgJUDajNpdIuKLIHl7i2C
/XNmal4SHiSO2BFqGLM9jV2Tf8qJusAAoc4Ux13dfAeAqhDymy8zkhspEOzx
8LDBoPd+wDFnMEp9PQNk1FqpNakGk6+GRK8ODeTDntdL08XTwjNkNCfUdbYC
6/XnUmyZPczne77Ie1y49y8Ii6nhRiCwh2CecJTut3b9P3NAnl61PjsAHtV2
SwSS8B2dKpkE6FBhfndfeWqDRgccAvie5JCPKx24TvWyprutar+P8dZ1CinZ
vqCfB1bILqRIydj+iKO2jtJjDkPrH9jE3jntwI69AJXlnSXH6soAu0Jx+wB0
masc+HqgpBR4HWpE1KZPa85Zm5cDFbEhqD64luAurIeh/4CzOS4gP+oUAhAN
vekWnQVTJyrHL6j9RVBOFVNOe51nrI0sWtVC8U44yzGAXgPxNTlBdp/KZnOc
TBJTKtxVgSDg2gWofnEgga5Mo51BXz3HKMy/q5LR8Ib7xj5ZuqkW+NFw0Myc
vvQEFDRxz1YmnF5kr35sb1rDAV4ggiEUOoAACGyMVpsXur5p0K6Q5a/tnzg1
l/qEz16jFYPBhzuFZPxuR9meV7CTsu2v3B+6ykVwcuPgiodMto0I14AOLmbG
4LlFAMig/XVyOjYffSSUdLry+z/cCHf4wK4OUNu8y28jf14/YRDsN3Sa7X2d
ZnKsRrrRgdoTVd5Zz2l6rbrsPJd0Pt1KAIrL9nmGYZ3wti9NWHITG+OjlRpG
PFHpwhnf4rLbgNHNGknB91m9VO5qTYClSJzZaYWsjpxrL5iu+qrruAluyUGM
mrSsEakJiMbsr+upEG0Ou+jdASK0q18c7AsVQQ8SrYACiIA0rok0tJbGIdzD
cX8b0EP0ljHlhw+DwX4fRW3SI4+UAqxJ/dJ9wZ99CAf5WlhAn2FRE0t6W9pY
4zunyxEWLtsJf5NNqA5EEkqECux/XzSMSMmKMib496MnROGMvJF6BTb5F6bt
iaabrR265gxOaH/fdQ6L2iAjuOxALqn1Q+Z+oJEf7bJ1je/4TN0nxqr7cYNz
d5p8qDxpgRmCXH0I3sb2mF4Ma32xtDAhQU89q7yB0EelgfGCWZc+kfFMrwvb
5/4J/CAjpe9nmMsEIZnO+IO/pHzt9nC/LbkP29OyTVTP3qgvjBGf8CSiry7Q
re5Y7uiM/sXwWRYggdd48xGwnCN07cJYzE+5k4dz5HDABXJx1x1nZPVivlDH
jKmlS9/7zdmfy17AilETm6WZmZLfHydj5QJXFVU+noQLYF7aTy7/pbYab39h
wtQ6yqaxqai2uhrvaleRd649rzOti+P6e6wF39pE7t6Vq1dEJMaMUBLphkR0
ijXoKU0ihUv3G3FFrxRamYCrGync7/r/ZMQ6EBu/Gp9CWDSZg139MLyp6/+Q
n+DHqWCdd17PHiuXC5AQEvkeLfUpQtxy6FumLPOGDEhc26zwPfXsFDoielh8
rKb2XhvWlCpbYcagn8Se5QsmKMpH3106TpFu5K+lK49nDis713nTacJxIgyt
4tUKes4YlnIJFTuiVdrUCrgkKUj3dVqr94SdRI7nQr0rsO/5sKcqxNMZwEfI
PxBGfwsvLltu558lq65j3nMDHLX+16YbkXOqo++3WQ5IW2ZZ3CbcHha4oeKu
8jrYN/oznr72p5o9eFcVcS0RrfISsnlKxyIDkygg88qpIGHbN+HcRvhX1zPw
xc3nwZ5pgxhL/NO8+bFqL4cvHODE76ot0dtOXf+L/asyFLC1lEDJgf3spuzO
ND5oG66cYo2dNN50P5SUdcL4Cy0vOKPGbS/f3oqF0qaX/OyVSGv8xsuEvJR+
VXrvBNmbWTnUGhP5FI/KzW1W5JwIwPP2frNEb69Ws4ns3QHH8gulXhbwxxf4
tDFMWKbIFMC9+fVLi7C6n5jry2zE8K4f8tRoNtnWZ0Jj6kb1B1xTa9USKrhW
/qL9D9k0Sdi8k+kfDRRmPV7FndNi2W5BhxdexG5jRYJI4pnP4qMjoY1xnOeA
qR5yWqQzcIulRclnjHIYZfHYtRh/8jas+gEOQupuiwum1Ykow5Ql21pQgHQ/
fw+ZvlxRdcUHcLeRBYNS3AiCNnaxPHfoM71PKJh8Z1N1kOA1EVmo3xkSh1X2
YZA86OWNvAZUYjEFgbDTpj0pqVVFYhv7GXXkxMeLeAARiwNM/He+2X/uWV6W
yEQNB9A/hy5svRNj0Xm0mbAje77+hCbRBFAXj5K5//QeP+KP2w/l1LgsjtA8
8uq52o29Tj51Meyp9EdDOM0KnqmkrLpimTYTVQ7HegNdv0Lb46Tw9jXknxjk
wotXuaW0wmb6vN7L2/VAeIYatnF7i/B6uvlk3Cr2uYANLdrrQlWqTVp27NqZ
AB+VnmnbbBQ7KRjFuOfrBNSdp7XDMeMVe4hODVKm+bOWGjOEibnO5QkVUG2Z
fK7QUQ/ekMpShV9KrTc+/10CAeJLobZk44Dp0LA8wH0waCgkwwMrPi8vQ8Wy
RCcPg7HZ4aReCQjNv9VmTBc+CY1zklB4x8TLpwGtq0P1LX3nSr/Hd/UQtBYh
hoXf1Rp48hMzdv4O6ZQO3QDVVmzqYnMtNxAmA3EN8NVc1mhoaY+7SBaId5dq
CT4J6mv7YNooiOioAaJKEwTTT6ddlmq9YIx/HMwWvgyMXtJSsRr0D3svOEvp
zgC4pVnY/sp2Vc8mOyQzbvQndvML7JpLs9vRjtSkNsiVMrfMrcZqZhXPEutV
veYc6k8CLSA/NMV/IK6MPT8WAt8GpfuXRdkNT6IjLwkXi8AmGc1i9DSua1U9
soK9Nzw3FfTdlMSPJsbewOb+vcMFCwiQvimZSivYK7gdiAtAl245uI/EoJqH
CtsNHwa/wF8yxhm6I8ih4BXa/452eQc9KIa4l6JsTuG16Yy7wIR3tzA2C4sb
jgDiJe0lPD4BGnQM4OhVT+3HDtaB3cOBEsZbt7la0NPFJ8PhT6es9NfdkVl8
Qh913rQIooBm0xwtEbUVvgGut1iVdI0SHc3bb7WC86bjs+sORylKnJURKvef
+LjVqnrR+OpaB+3nFxJFNEs3eTwk1BdUdRtqta6T3EexSXmbu07tZwdhUjiK
YZMmOGdGRa//Z7OtqVpPnakSi5hr/b0xdssHWvtbZ5df4k8fk1VwU58LIIR4
fwV/BYl6ERH2HIJLp8BZXB794u9a+8tNV9RDoGMaVeEo9BPuSGkvL/cipShd
NdQAOPa1ImwgN8sbNPSgtPNAlP8c7oz30CbTip6QfdcwTFdYT4fR1Pr9i8A3
/cfCTes6RmgqeFVmol5wTzF7S/F+Qkx2/U1t7SGegMro/BnVC79WYwwFiRIG
O+e/Dw2GJndY35aDIqr756iGPVCcPbZeosuqE6OrxKkyTTD3ErzwtzFWUZDU
uBZ6WCIX6Hyu+iL+QoyRInsTIK8F+mJE5budRFA7Cp6HuGF/CnVwk71X8R6D
pcyEOegS3rQbjUgskyDvOQz0Xk+j9vmn7CDJzUhlVdr2Ff1kpFuE2oYriiGa
8r/tgj4ZNsjV1bPyEXic54sIb2ksbw8jxY7EEOgZF7w0sBspK9I/rJh/pbJ8
qVycP7aTbnzN3RFFaAwi+IKyWrZh9L4noXeCjuZblPclBfSgCbYEkFm5+T8J
N/xwB9zb1b0RpH1xilyugNWZ201v7AvYcf3tM017OGGv2z/WoegcXmrB9m4x
5FRSw/qSokrKI2A1F4yoH9KmxAL5VFI3P97N4WxUotHQTemC5Y0A0QB1PXFO
GVhW2Jbci4hM6DV6M4fiAYa7HoBQF8U5rwzyBzM30Au//rArSZH4iEER4KLj
n994eTmUsfAlOwSj7HEKJ9AsNvIzwegZ3aKsFxjG0FwlOPlGViHKB/LaXFNR
2HrOPV6zUz1twPIYTTSCuAJ7CgX3jDIAsr8fdRLse4HZI7sQE3fC6k20sZgM
RDPjS4QY6QQM+7taY6qEE3bLKMav6lS8gDcdvQTbuWdV+tcJJMkN26VYhR72
7zLMTleHO49Ri0PWDw7n4bOIoVh8FP01c75QzSEQmRd4oQTXSNqm5sYmwgS+
50mRBOgUpDzBez9pbFVlrnE2KEB35WZMorgZC9ZopVA+RcZCiwNgUbt3AnFg
GaB/Y69hgmPTHpE1NoECWNs0AzAaam13wKmq1CNbmm/HpbhZn2PDIVfnxE3K
NJccWd05+ouQEi0hOspLkHjRmjSSImdq9pSwaGbw6YznSSCdW7QWvKSRSIQG
dgW6xvACxzttZtdYW5bURxIyUcYqPXU58FtYOgYw+KmK0cNzg8e3NEe6GXsl
LOfdRNEfddy8qcTXqLj6TqSqy+aucd/p3IkzHZ/l5j9/JujQX/wmB78D+wRi
UO4E9Ez8q4nUEC4jWrdl5YkSNcNLr2Z59GuDDOCx4fPaXUZmoHAIm1JRLKPh
Pysyerb96+kIwJvyK9+P/qhD4i3K1z9LMe7/O+GWKHgN5+UxhRY93DHIAQ9g
LRCtAZG/UBIvZkhycWg1MzZOFHodYjH02kbpke/GyS75MQ0Ni23uWf/QfOWH
cX/FfzP225iCEwW6I7rVjVMM3oyu9ibD7S3QUs9mcPswFcRnFkY0ULe+CHCA
JHQOYgKymdls/NPl1njS2h2uPWiGvulp7Y2pmGpcp5r/goxts0BQzq+N7G7q
PiC5TuyfXLJkaUepQ3WS1KY5cjF5jCKfnq0l+VkIRAW/VOLgbjrEeHMg8NiA
qy6DhrKMO8WdRC3cRr9RF3DBXlcjx+mS+jHbqg//EcDJJIRWjhLc+eSfGhRK
t+5eLtyfCssLpqXQgiOmMWCJveGtwVRtPhctcqJFIwE1HfGtlggUwHcsik4H
hF0SIrr3tx88fAFOM2Iv12KS8WWQDOj/K5epjrIUPaw26sZNgHISQuahUBSI
RTDYU2YFeIWpM5qSLJXN3ia3TPCf3v62vpXGpoCzd6i9iNQBmDo1dphEy2Ya
KEg1E5AxQr2pOzoX6tRZ6x5pqQJ9INhAN2dRvtFWpCX1Mz+XxzIpG+urCcnZ
eL2TLe4hQwauPru1RAbVzKFwzHebQuWyLGJYQJJS8EHo8H57mub8KOzPrrNz
jTDFC9yV+nOi3g+uPukxFQk8VcCDRWPavu6Hmjj5tM4vKW6+I6uAfe7rHfMN
2gWFYgQs3kP/Q3rEr5uFA4uIIDqaFoxNU9ReIWzejm3S9zx3j1ZfqiLDoC19
baYlXXRuXzDBfPDbd/DLwAFe6G6KP/eCJEkxr9xYTSHLoWfBCdQpXpxwcBJL
OF2vOyW/Nyis0aUuZR36LOJ+hKj71g0JZdiZQcS0XXBzedD0qmU16gZIQCbF
RuLxTYK+X7t3mrqqiAppQcISngzCiVWYOeoCJfvdl1lG1SCsCjR9PaLCemC2
M7YBAJwsIX+iO8e/ELggICbQMn5K42BDLAiwTWAOsNr9eAqVlocGdaeAx2VF
5YMWcuZdh3Bca8moC7GKr4T2kWSZHtVFqTP08GiGx2ixpn/m/GHHWwIcylZu
9h/+wb2j6sPcRrMnVhtQi1iilCL/czxg6JzCQ5E54sBgdaiLzsQfd1ZgvFdi
7aFgTxjYfR+uW82uW1fLNBWD+YP/cXpDB9FwQ5M2NxHcgZTImenatgDdjSb/
e/wU8le1sKQXOfKhriMXQjJI0iSiGZPfAuVkAKBWPSK7Nzn89geI4/CDeFcm
dyz9ia5RcZbvfgAlJsIy/x3Vexddvi2hX3yQ9HUHCEwXV6PY5YuRgAixJsLY
ruh2ImHm9cA83MSGcX78RGeiDZc+aMQ+pcAZ1Do5AsP0FVBZLDhJdgUs5IxL
h/iigW5vw02yIfHILL1uw+kiw3VORAkWpaKYZuAxx45TMKn+Ef45zm/dTVzr
1tv384faPNsDCbkoY7JZz2mJIuiBvKMK6aowisM2qOlBlSup154ZNUIUYRsJ
PEqjA5q8JwYsLjXtv6dQqODaQxcZlY+6NeCp9NLPj2e3nEa3c7DDw1ET0sCJ
1bEGtStXnIJ5LW0aNZO7qd6aWL6L07t6QGyPUye4wjTshvhEJjk4kQzdShIh
RiI6hNki2DDZu/fgq2S7a1o8SBUQsOy+R732bTa0HqrbJN/0gjMcnIkgo2tB
eqagXyyZZdyiaFAiQ91A5ybmhPNgmVvvfhqij8v61IAKnKxpGaG4EUUOBHAJ
xbWksc17ASIeS1yXuPF+JghP3IQlJ48aARrSFyYX3sLskKP9B6a+nV4gx70x
0vrc5xIFtlMKt65F6gm1eQhjIFslGMOdoMn2/00xrR1OtdONaEabOon+yCIn
yP+ESEcZqZ5JI1YyGrxpe9FkRKmzLL6LM2hpob0l2CkOXoaMdzss1g607f1S
PkGFJwq0H+nq+KIJYhR3La4qHl6RLvvfhvR5EGYS8y7KC7QqkgOpW0+mNpt2
8hrKQwJffnifoL5xadOD3GuYaI2F6YpoUszL/sVWxbmE1xyLqGdCWKias+oL
yQT9WnQdeZS67Md9QaAIDRnQnmBQkOoE9jcTjlEE+2k/HkzIKypX+m/1Vq9+
r3dUl+jfYfLMJtty+/0ojc5c4qbToXJw7gY1VQnkDP5TA7zMyIn+7jji5mn4
IwuGD/4Dsf0MPp3AbzpSrdjeKfwAv55W06e6mXu74wK0+lJxKSRvrnE4iVi0
BkvhBQsnqeWn9enJOQw2pRmSQQdBXIuhWjBU9TCC1U1l1zMEBWZgVS4ehnx5
7ozKCbwh/VPXH03yWs4J8mEnuQ8Qv9jEvC1fC/Ypj5qMT5oKyhcxnTmDgfUL
EIxSG5TRc82zIhr8ZijwygVoWpvqB5YvcPBznq0HJl0q23GBpmonHST3iw0F
Eh6KzVMvpwHrS/FK5s2uCJPn8TLQfa03NoY6kWhPqVM/5tyfJdXH6rc5LUa6
Cc/MhenuXOEqnJZbAJ56e2A0DDs3TmbRZBTvSNZpj2C87dt74UJZb/9+EvdP
s25e3IEml9uKHR3+5Z2C/aM/VxD/cfVdpk4SpsOqPmRjlMt1DPOBIhKbz7kj
xcf0+IP+G4H8go+85vcb+E6t0zVzlRf9cNiul5k1OC3bF/jzeAwUOfJtw5Ug
rv1a3a6e1UKvnGF5y2TA9RrW8YUq/GyIW4v+n2iyDHONGkcuhPhFwdlIIzf6
x8Ybf0j0t2fx2j2exXABNtKUZaSTdFY19rsnmNnP6WspIytqpGDz6rEjV1O4
n1Q3yg/caz03eiNxG/Wi8X5MlbsNPG8l/lbjE5ngaIQE2nmz3SMDIM2XeiFB
AwrBWhU1J7gcujI+GEVL/uMa+x3u0G3eT8Rd3YxB+jjUgqFuJPmiUEmFVEKz
bfy80c6QfyA93ur7ud2qlfcLkHcmulqb6tAp79cEKZltVXYGpihr2tBVee51
1c+uF9YdM0ShYOfU3BQfdtodbkVDw8Ei3mIhI3KXa8+Wu86ZR9Jomd9ZFd2H
c9r6GUL9FWs6i6ccBG1XUBtgIomSOdT/OnNr2AlzSP3e1B06uYJTb74xeJRQ
TRhqXS92N0d7jCGfjgnDHZQFKT1ElMgNr1Ws9rRv4dNthPXu8/kU/0+lx/al
30uDqDX3r2Hewl05sPTFFmz3DM9hf6KcX+1erxz2z4kcssR/40deFLPhBXQv
4yrWXePu6K7M6Jvaw0IVB8+JubReTwFYs8qIN3OToN87S8h/uOr3aoTGS0LD
jDf2RfFhLntWHBMaOirNmMkBtHy3pFUchU63CtIAvlg6JhRuyLTFwL2LK9To
+OofvKLrJJRMbVwsbPDO5QZKpZAOkQAqTIovCkj7vGbC6/a+UykaV6g9J/sc
ZypooBUXX+I94H9MW9kOS7kGmxiE1E7CkkfZIWa6AcgxmOcb6tDYc4WcFTOS
Lty7zRGeL1oAgP9ZoeADiLFukI218iYdvkV1+nOUQNmXIdkFQF8+Z7xJaGkc
MjAZmVSSBnKdVXMBn0ks7zTbxiCgU9tseshCa+X9QDRNETqcz42p5WhPERPH
XxhQgxz4XW5su2vYMhKDFs9D/KYW6jIKB7hM0QNwmmmi/PlWsW5nYM9oQKVP
hFdugDm+30nASkN40MOlRQ0Q9ml5Sdw0M/pa08Z0P03iXfpB7+jHVlm6/lgA
MiPw9jBLZuIxIDm6IZCKVA61HAlVLsIEokIUTb7sMtDO3biHlgHunDWY7gPE
OwPp9NvoPTRmIxccjYGiHKv/d0qrRJD54lCyGo/iauNfUcciO4dZMQVI2HlE
4RSDws7U0NMcFp1y/wR7SRvK4Mz3kvkMClDnZoPoa8Csb7XXXBQzqVMQiaVq
BCTuQWeQro7pV0xV5UCR/ImtZKYILtVd3rRBWYvYucWS/Xz7G2MMiAhIzgrh
WUCXVtpojWOP7npz2D2inWuFaa5Mi5h1DnPm49aok1aBKkuvdHJRF7MiwKlf
8NpBrlMfAkezc7kAg740z+i8PzhskiHTLSEbuLDvP2+A6m/qz0M7GMYGXce4
41z5RRU2m2YhmOYCWo+YU4c6RUQUTR4Z7q5PtEoLNWDswNG45QBGxnXpJFRa
kggUkK2BdsouL1yYhdUluzmr4wJ77IiZap1fRxedLcbmDvO6GRV6YBUryVPb
bjZWurgFLy7w/Wtx61ymt4uZcvkMBd6gd8mtjvFiB55oHbNX5s1P/+eXxPoz
xBnMlKby6pT7m0boKlumjhzETSbxWSREqsxpUPgFJt1lX9MC6aW7xa0wmR+j
Po7f4kFrmT4VpeWA74LuJk+3rSvdxuARnob8qlQJx7CdGcA5Rc7B6P9rCyF9
uQx3InVbhYyAdC0IlVwyfOGtrxxOABaPdvEOO5K3fWipwFM1Inz6QGQF38UP
7wyQb2GO75OTz3CUlhnT0OsoI40qGpJTkW7ccGpTU0iF0zEIXBNp5cyz8r+X
cu6zG+xX3w68p+G7m18dNveLWKtMZ9aepSsm0/fZ6hdFEMpELNyEsnqGaC/4
QbZvYduxza7xOkqrDH2sgizinUF53mexRpZzrTESY9RAx60nln0gBLskQ2Gt
t4s0wXM1qwz31M0KrP/WDdeW9q0SUxTqCJIukdKipFOD0Kic8aHf0au1CDgX
qYo53pEM0NGULNgZbLP9okCeQC0IKj1lWPOyM4tIgtI0y+Bo/ynhatwKRnUn
rL/FtpyLBMtiMVpiXLwVmWNlb36oy9rxx9Ft3STZnO172pU5aXE2lC8FM42L
1CvXotvpoWePUhbII1/BbZfVLuWAeNUANNUow6e27LJoujg1+gzwFtRJfhLh
68g3MbD29rLBZLM4j0XKqzmoU4H+qBFpAI4T+mlj+ZEdp1bn0zOsW7gDc5g+
FaxHZK4HPZF20BIr6E/YOP5Cmv5ksOPLXHiyi1eBBoF3UiUVqj1p788g99aU
5VrN9e4qx9knqtrC0bNek4y1ykDV/EpbxNZs6VjFvIOebbmzyPXt5Cl5b8Y+
EmarmEfp/oaQGyOlYb2XqyEFjCYbpdmRniXsY5+wcfAR60Pdyxaqnj4JHrx5
NpoI8ERAGgUFPyo/V+3Q0XNXK7yceWFyA01xdW91qe054dC/Je7hwghQGMwF
wfmFIVAfyJd8Ev3cmos4wdErXJNlDI++5HYFVl+Mnz5+LwPVBYsM3jee54Cm
qvsV9IRKdX2vkFrjPBYsZP3rXOGT8mmxJ1lNMK1xZfYt3bSCe7CM16rtJqGQ
QOBALdLU/dlmx+P4lRP4WR24IbJBIptETNMBqcS1DQcXc5KBPojs/FvDhVi7
AFXIdiYqpkdve061hfwcmXvx8fja/vqGSr2YwP64YZS4F+QX1dOZ1L03oKU0
dPHsoeuLWVnHN71zGki2ERm12nx/02UeIx9EOPMIztWLPtlUIeDnvDadLwu+
05YrlxjNck1qX5Hh5azrtGEGIn93JPQ2oT47aNaMBbvb/vyxcxEWha6HgB0N
G9Gw18HydtIde/9bXqRGdhz5D536fSRC5b3EE2FsAUOK5OdZ7qTP/1cVx3le
d9Rjko0B6Xhyau+rAklf12fnu0xczgtFziHLlXjDVzS8Ue8bXgtH9tCkzdCz
lCUiiGBvHCXxBz3RjrIXQVPZX4jZZteZ4mM9jVBySxrrYXhGZrNAQyvKZfxN
Bq5HdN1wAdExzOC6tc7VsPZX/m5nVyeiB0LbEdMYsLpZdAUp3sKQqDwdEbrH
0PHqMr9z99Dvbf8evKdRo1U27lIkQiqgcMBGmvUAiliJskXcJP/oBQKafLgZ
fimJiWuvyttgWmdExA+vrZswIgdpTXOcU6dRXzeNpLqAVYy97m4A80I1wVAI
Ny5KJqw7yJQtXKvWOSUaZd7Wk9jc1Gp4eUB5qUUBHZJzNpX65ThjqrTwaI+R
t2h4aN3GgP4YoZ5JdJ84vYGN/1jllhxv9HOgy2IcLf9e8PMsCLqHro1eKyk5
kexCXBejuSJq43/nI4IGg+7dRAdg3MtaZ7RQkPaHNjyAh0gcwv7k/noncKsK
hYpz7BRdS43fYYd4CreSWjJ88/xJ04fb2d7x78rASha8Z/HbnDYnpGesyBIJ
yc1j08dUD9Wfr/to99jfsz/YTJqE/5IVCne+92gnRliVEY8ZJRYWk1+J1Qad
tVgubN1bTtYKh+heHMXKp669DEiI0KyjE7Axqm/joIEFgy1iqgIVSBzSYm1X
qarLZi1a2fqCeIGbZeZnQ0qZ6lysoVQq+daSeaUOAZUSq6LiPdnAfxZZCUGL
qyct46ltnp1d3iVzyN9I4MuU1bPiq2ksU9qojGCK8CCEFtmT1zRZonOz5YBq
D7ojv1BAlOae8AOcEVUexEP9SAPv0O0BOp8A87Xql/tyMJ6W6SjlLwo0dDgo
WCqd3DGrd2Mjg7+Cv1yMA7yZqdmO133Eg+Udz1N7zGkwRqeJOHp7jBoC5fzV
7pDz2LhExn348LWjI8XKSR8RW2BhA3J4jymvmWEFyis15t5q+2kHKd8SxQXu
djl8KHMATImlQWQBeBQlh2CZeNaXpaYx58Uj4Tphxfp7ei2niSu3apjAcZFD
7rHrMObQonWDwN3N1YFSFNt3rn8TwaHanyRgFlDgmv+gfqdMPSzhb1rtPPBd
GxhxKz1zWX0H9j5wYTKhGECjsdi+VzJgl5R1zMI2Ca+Iw/eT6RYssm9WM1C5
mnhR5+ssxnFMXGyins5ympDoDTBbZuVcU3PfP/DUlPMXNwMPDxZob2Kz8G9u
F819+7IUBV6IjB27tQBNQTWN5RGbj+15lPGgYtCZ1D8cqP5fDIWQrgLkSsQP
72CRrFwr/6c122kpo5Bc4BZTqpsH9yZXIujGYtC2+h5n7JbYTtr6lRNxeuEN
xoHwdYlgEnirqnLY9y2TLhyQ4TTbmR3Tga9hr7rVtuUBnZqbZAEIE0xf42kE
dIQIKq4TOPxOY5OpXNHNNX4szs/EHcQztMJqUNqQD4DL0z4nZcg6mKnNQAH6
VAz4y3PGCrv1ZggAZD2o6+c8TEeHojUDQbX2cO3Ra0dsit7Ens0crtlPAyg4
SSgs6P195WnEqL8ej72a+3wTOtXGAhAs57B9mE2RT/yJhLd5WGf30/2LV+56
HP2ox1UfJlu3cPT/BmE5FT43UbFQpogRdf8PUhtI7Fl/F8FNf6sfQM8jaD2a
UbuFNIe0m3VdOUZTL7M9PsmeEqANsxifhpC2yDBl3gWVOoPfmX40KCHwa+Ip
bEhC6VRmlkgoZHqo5I5VS4D5woHO2n4rAECjfqig51eHmUzQ+MEUMcVpgVx7
9IWt9sjebPGPMp7I5ks4fq3nZFwRJk/G8JKqrc1E+S4GPL/AWrSwp9pBQL3P
vE7NEadvL6aeWpg3waIHPF5PVf8TWwfzVA3QNe23UhsYiNOcvFybmDU1RYOt
URBg5XLmV0UlKTzdK3G+8+d6ecyaycHZDqhCwqsBB3aF1p4fDBoZ8CG+Ttee
g/66x/3oduYvdmSI68WF2cAxSNodVT4sfzgGlcCjZwhEYuMIKafopesOaJhd
dNDmLVS1kFcaqT2PVLGMlTKpJU68QS379H1Ncmk8FLDi1kxvlsuIOfT9/h2A
OwKIJcE0sMd1kuaGUeIxoG4okHV5GHWti3xFfOodac/6pMO+tppgFYumsvO3
O23lqTkZYq51f3Rj2mjQm/tez9y4iu5bPbBjEq1RX2/FbpPKuVbwvQCSkqZD
gRORtJcv/iovomUitX73OEBqWSLwRDBYrhTBEHcoXvyVxFuJMnvXnNuGqC95
gWdtPjbFAUHlTjIN3GoV7ear+rTzEvlUnrughvVYhz3BtBIw+yMWptRURhSi
dLgJQ90dlFDHJ57xDY7IHlSHxuYL5UShINFZUTKuRPXlhHPW32pxIUTlGr3r
7gDraPJA3F7MCniuHUHLNuLzA4+hw1X8N8N4hQgG1rLtGBo8hl9S0qTaPeFr
CocCafqKTqSwf8o4EKBYnPKcO6DnsAh9wxmlwjawsD70LW1mujuS5LaP8C8d
/BAK65ZERzx/bPt3fkUtAoBDPcjLT6pYjRG8WIn/nKzVAKcsESbe7/OKOaCx
dfgDIubDhuub+jgvptdEcjfIQ5DIfXrHFWKgbaiVfMpl6d5VzCOT7NJk9l0B
lrCzRU78SZVfu+XMFhcLOcTrN1XO7Avb7dJ4TZ3cPwNBB1+0i/YaAoVyfNE5
2BP9dAMg5jpKdCnX36/e0SJ5u1s0PiG2oKwjMnNpqS77nf/O1oQuPCUQ7XHd
xPfPZtkIdGNlXTRGnDOgTW5LPt3XgyX6QrI6cu3dJYgGZXHNU5CXEg/x8r1K
Nw5Vrk94iR5ITTHsNJ2kXKLlVbRpEYrmmrU+7BjvAzvneiCzG2s9yFABETQu
0gbFJohhw6zLjP6J5CP4t+Ydzza5g5aLnjzPRWzlbNNFxVni7DCJpwVEhVvi
B7IBbU2wr5Hk9hi5iUxRBYTBt2qy/EJY87P4Llz1w0bGzCQylkjVcRHTAygh
EhQb8fUDec3aBdOYhYlFmzCJ2PyGZOfTf3k2BJ3WSqh859zBPiPKyXTJabNz
p1wQ69gTst0djO6TRSL1iP/vOeLZqCH2/OQdlzgYV79x6PQlmi29FzSZUBtV
bgvv9BXooYs3Hbg01wdf1P1u6CyqHJgX8ixjQrX0yAFxz3AlBPhNpbUWpXbx
IdNUW/sSM7+C4gX6FMR4BCPIo3io2z6isFH+ofpYkk1bLUbobl9NrJIPIqYb
re0ynYzQ2MuFUfRyzumdEICDTLug76SQbaaOWABBBl0G79EQhjHkx3jorXTa
FxXQ1OV6xIVqRJm4ZRP4YQvFFVzizc7YYh8xw0Sp07pvujVMvEpl7W9RJwt/
kctkLU1eygyabWq87TMV9nFoTQxJ/Ot7cYNFvde8GsICi2d073OWiPuZw9pU
0DU6QAs6S+yrvGJtB3/gQsicn/4m9LS/dUCo9hyANcdcL9LkApDhpgan5Bhi
9/Czpk6hteYrziaW5djkl5ZCCsnNRJMv+wD875V5iE7Wm5YyvZ/2EJcXJwvO
64KlFupJNBKVBroLLnE2XpYJHdmrQJZw6aRONaE/8HoUY0OFMYV21vNW1YvP
5o14ic6DXsWNPI27+JNJSbr2TJ7CBm1ieiSmLnOe35X0vmvBt7WJqvoPOkVB
PT1Mmk31Mwc4KbgFpqkyTLsnFs7Na+NwdrIu1Aa2HS9KUbjM5HyoIQQGZQkB
65YRFN9m9RKAbtIjRKWo4gHts3jXNy3+LpOQ/D1bLpMtAjgiKPIyM8Yt3hll
LTvWUpLdhbkfDu8mA7Spo7W20TdGdMxSZOBkldiYqz3BDf7am4YQ39domoPV
9wyI+bMlDd6015YWjAC2jBzR3mq6jzgW7Bg6r1SmCOSmbLuaTkPHXxm+YgTI
VyIUzZDrjfYxdQdipklYEGK761tdR56oThnRYwV3RASFJGutwghcCnrHjNYU
lsLLfb8KW+KJjDSuyNDb9mNmN6JjIRUL9Sn51JblCXDe8XhIRrJXhOYvilMM
zcBRLVTAsxt0n/8hEUdum1iTEbb6sGW6uCWORJdROw+rpJ05TSz2z5LJ4TXF
b5SgR4tmZId0oqLrnecKNpuiJVSuwY/0iVwYGQJTxpcAmEyilHczr2yjJbcS
PKQ01By/7xh4tPp+q8mw5m+6MvhfsuMLgt5XCOzzeUBFQfB522un36Qjd/SJ
ddXe6bW78TmxXHVvCmLjiHCWtVrZXZoKxxxbZoOytrp7i2YJBa9WhMBCVW2N
DvmGuwwRgIro8ewy9SloWzydkvlcJlKD36kzwXo44pbAFazd7vx/mC0ZYzZ6
SQZafLdZfuYO0ouRKFjLeedIq9fS5Q2zhqiTwSIvvnDoIMuCi+6zwp427lFw
S2J4Tlz778bOiMWYUZhWlXt7GnIo58fd3Z1qYDjVbQ0FEWeMcH3Brk+3G2J3
Z4Y9BR//Y924TYCMYhB3bvhxWpt678GkUkttlb+Gt3Z2uVxy0SDQ4VqLeTQx
CQy3MjSMPpg6ZSKKp2pGWZJ/i0HFxemOgTW+zAfzBboTYYGXVpsfbm/MsD+j
S3yCtppSrhB3QfrZ82d0Yx5rbdQJYsKmNS/7/bNe3WJHrNSvUxyVRpOmxpEi
3INr8OV0ny9NC08QMKgmIiLdgp0QPVkiTyyWJoLTbz4p0AqXflo8l6i9H3cx
NVpSc5KCMkr7AacEPJFohGfg92GHXP0KLzKklgqc4XITBluxhFvLNq4dYeQM
A8puZFdiW1A5lz80r9FbNvO6o9IcNrhKuuf3E3vLO5O5A6JvF2AuoSzz26c3
iJFMeaby2kLUCHxi5CaVGWLA3f2lre5Uz+sI3Isvfiu4Renc64JekyNrAjLh
8I5oMQHcXfESxXx+5HDFwLTvKyop9jbETkX40DdB4qsY2nn9AT7ftPANAu9y
dkzlBSkzUaPOFQd941AfxfvNiXvshstaxh7KYPPE19EwxDznZ+AxJGb/PAOh
+n8RNBNm9p0LAQ+GKbwArrzaJ6tco6eNFV2bMNVLM1vvME375T9pWVR61D3A
hh4fuCU2nCqb6118YrgevLHT/VU4NcrY3zoniFGXBZmzox/wJj3XTAHUN6DX
bJut7eUsUWni0uZpgjBbRCTVOpDX7bZDFAQx9lbKksUn2s8PrNQ02jTN8uof
lbY+nrnyCRoSIi2zkcSPX6ZuI4BfngNTqzS3PVJ/DOH5RePQyXcwEfhSlvu9
UrXxSxzMeTIpPFYViLnZX8CZpF1VBjg5Hyvn9/LISYngm0hQUHOWpEFLcm0c
JOIiVufnuaf1LGPOW6uO+kHRW3opZNKiP/B2hSgnl5YDwCgBhb61RCnQbV+1
dNR5XE4e3nRgAF5cFO80eBMAxHiBCpsSbo3yzkyoERoSR+e4W1G0SX+eclrN
gEune0/OdnsgpbPSQv62ivY0miKW0wOnPQJ3hMdbsplhiGGJaV85mYCPha/e
p3VNiRAhuBu5Z09MnI7LinfT00Rrem4ZnDZmNyN+GJ/jUkohnordHIusYsgo
FeylVQAxfwH7gRvqWvCU6zihR8sW1hCLN+VtHSyjsh3BJuSxg4jU1DLtLhgP
wwDgvmINKwqaiUnAyQVCXOjMKjNM4dJevvLsRQhzYOy1glNk48f5PNSK9+65
g64MzFrmc6nOYLh7WhNNVnSLHv9P1sltPY2oo7CGOR6wtsqVsG+/bbEGJMlj
JbeTED+UyJUocOUcnPY7odRN70oJnpY2yP6Sc0RlEhGGqLKdMs75ekz4Pnnc
u6BoCZmJx/xAYhl22YOIfb+rY7DSnghqcrOrMTXYQpf/xKHYTWKFriftkbXM
4g68aTqmQj9MdutBs6UMYXKIv/dy5vUqXaNQyt/paZ5d27/YrKvcPYY3BZ2v
xxD2moa4ohihC6kdjxpEKeYRglsuNqJ/Ft+JW6hwLr0E5uW69leFSXvKL8lk
1qDuND1xTCZBU/pGG83ENqnh8Jd9WWrQbE1jP950qFErDh6n0joUVMQg3RuI
ZMBLgldaIRu4MoN7OSeMtt9H2BBsUKiPrcVxGvAgtx0LkQZUlQB3Oc/N9fbD
ywC/C5QdU8JF017ISyU9p85m4c2PJhbWXCHon5VsbvQIDOZKNRhed9o3ILfz
USmLSyUGDOMxrJih2wwH4sigYFXVCyhcFhSCuykuE1iHoMlSGTEC5x9hUktQ
BZ9rT7okFLsBBRpWVR+/AoiZ+Bjakyx5q8l0w9slRlPRyWY0c5LZEjW1vi2u
ppTQuDc8xsHODtYWu+FzihC9oIquVWEh2uUX1yccZq5fJmGwsNU/hi8b6moe
H6PJHuJJGrRfWahcttNkkFP5MLqvsn6c1vkc5PwlvDtA9NqIcarXYCxeTxMG
XMnUNRFC2mpGmno1dxjNIKzz7krRDSl+MLqo5X3PNBFWafkh63hRN7OZKTKp
nW1dM/D+16Vq0gKESAURU4XfsNvsObr9zJF78LP+z9q/cbwvi5qf6j/w7LKD
JFPrBc/hmvtiHBUSJyFWEl40Nl7gKFu8WRMV5Ug9GKDoIMD16PCm3OJmL2kl
P1040fB7NBed+W6lAYtz/NThBmZy6Esi6mxm4qbD029Fy8n8naN93ZX9U8jW
YInPFg4spKIrcRCTc69ow+qpcOTTNXLmEUtoC2EISRavjyjJ+0LJmBfM6ipu
ou2dYE1qY+eZ0GdYY4Yo7fsggIxfvZlMBhR9M37TJqRyDpz9qPJN0O1t3fY5
pd1fZSYrFXt4MG7anzEbJye5I8wFw4MDQ6JEWxFLouwDR85qi9za21BHhMtu
qewdhoEYsDRMO6UjW1Vpk9ae0x2/HiXYtNS4b2y8VTGPk6qX0j2v3+HLDYxw
SqCqDOHQ65bfNed+5FeWvgXxoNSIyu/4DQ8TYUVusss2qPzZUVyPSeMxvmTY
/l5Y2jkrqZpmAlvkZnruThXaR+dJuzc8FN8voSy9Bi+Wr//faGFDhM+OD8cM
bJraKnxGNcC6M526ohmvBuQnZ/bzXTboc1PHAuR9cxpy6s1ajJ1+pkuWKJC+
zGnJ4iqpugXMzj3erX6y5gG28aF0jVHhmh8DqKPHLErjbW6eGi1p+MjxftX9
n8QSva83Y/BhYU14Zm9csDe80zQkrcFq05e5feMSdSlCuGT/275cw/BUVoSh
L/cGigjDSpQfx371pXTkh65DHv8CWkjkv9qLpZ/Awi5ivy3dDyItU/l1NrB5
q7f2N7wmWRXfRFburHfU638C9EyDu3sWvSYHAZ1+US9mxqOvBvHI65iMYYLl
OLPvWR0zrm47W1gARP78AcFk/TFa7db1QyhZ20LQFkaYFa/OHTDh1V2iu4Rk
U6hvF5QCV4FhAtZ1d+/uPd9AFw7vWNhsWOgAW4OPEo+mmJcKZbmr6eMYPkF/
m6Rh2obXri8wVGn/l1pSyYD/tA6ETZARtFkltBkYA8/IMiNM8j5w8Dl00MnY
Qx2Ab7k5PGzYf+fAL6y88NtDzbgEtZlBfJsO8kxt2k341R+p12MaHRYv3y+h
LkxHpQK2aCl7/CSQ3TLJrBRQAud2T9v6ocf/hahaoawV6f9nBDibWV53ltmi
oKMdZoeDJuP68t1AqFS5j/YUX8f8zh0+1kjrQw3CQ1NIbOeskoGYfzK5A6fa
YVATVmaF4Mz2rM430+c3QKT9mJB//3c6x7m/tjPWyWsLKDJgkCuV97BNSggN
5g277fsr7lOBxwy13LOiONFDyKXpbI+X3mO1I+NWOGDHtJQ7reHTWi66NebX
YKdHrXUefUZKV4Rnu4ILSudDG7+MixMjZq/f4/gz+TX6OW5N6uD4angb0YWS
Aly5Lgl+NCRhA8tIASZOtmewON7u6CxsqsKIkpSEJdmGcGVaivlweBnd2PLt
Wi9sffsuxCBn/p+yUu97snSKgDT0rWH0Si/6N0/ezO1WTugZspd0CZbjGQVw
nspZQCNqQKqyY9p7LWXe01/zPf+u3OAHQgm7ihOBjrFZtumBlLTgskTIohIv
9/JzUklqD8QzoqtOZUWLwzF8+AoJePAEiGTJSDDbuZlSSHy0QyByL4zpWDBx
nGQzs1s2VBUA+Z7r/Qb0IftoAvxEzHAqQ1vIqQLuXdC/sO2Sse9ITih3mO7S
pzW7pFWV1bZ8YGdqfFRhJMSwnPAcOM3Q3nZop4p6W50qLe7nkeM7nzTsk4Xa
ASzHfSGfoa1qt7v4YP3nDRX+waxxv0GV5MLJolXFCw5CcC2eKtHQMa0mYcIo
Bnvo1mu8pAUVEtIQbG/egy8oBCrmRX7xdBARWeMzs2MEt5jCcKYoQCwKbqNo
VTD0urTSRsb95wwMtIwjMNdiU++/tkUjyur22ojRucZfe5Bc36xdVJjuvnHv
XzMQK7mD+eSVcqDaewCH+lFVNV6ppWkxyVaklodoi1DXNX59USJl4+KzDj4b
LPKC0laffDQCoPnz5XNlO9pIWvcp27xrDE+nOLOtTmaHbvjnUsrWNA4f8jZJ
MfT6fh8KXgdMpcd+tWR0FlmkMMvoJxVv5lrpLnuAMooshaQcZdmIreqT9lXz
5Qo8J4gyLqJ4H9HbQDk/BAf+WdWZTQxLj4V3ws6/mIkfYBjL8DIOysgIaNMr
Kz73bsvvRonBKItqMmyPw8DYk1ILcML8wR6hNjw3lOWbs99IN2y3ORPP0cGX
KGSQsSwh6BWK4YE+mNH8RKc22bsSzpn0vkPApyz9mCmDAsvCmb1wLPE4fp6y
PIELPdJ3WIT3dj1GQ3kZcGKUIuolPl7qdad1ny3CmgzyTxPRldF3Pi9flsUK
pRwYC5Ce4Msgu5qW2PGMuBGp2F6d+SqJnQQNLxYnHZeIgt6sR/MilNdVAbgR
u5xEedHYFp3fCM18UC+tjYE6hiMF6fDOWRbZnBVP7cmTCu/i91BrG3DDDyWO
lpBfhgdG7XNJ1+1ReZ7Iy/QRbu0bHsCzu7Jz4bTIP77vdudenun+rpQFZ29g
OIbkNkN1aDaYelfIlgrTDC4fdZfCYtGwazpj8FwxvB1abIZkFy0gAqsamS8N
/P6uUawbrW241U0O9LXdWpAQHtQgx2TnSVByiZjfk8KPFGaHgBfCvf0J7sK8
FcYsEtoIRqXPrs2cwfXXPRJDsJo82fkpj/fKLLvzKYg/fqYkk4LCLfIokLW1
jTAQreGSKxFh5D1G4V1MXn7nQsUamVn7jQfon0OGGyiGgNs6gaS0o3dsFf2W
GqHS3PM5D+qDQjA7y/GE0L0COHYvishUTzLHRlsC6DDEhF2F8p19VvyWMVpj
vMnJr5TW6/9y4R1EVbDuhRz1lOwSjoD+G7UOVjy0z9Hnc4eI3RGiyDRwb0j0
5yRnijmjSvZ4TKqtTJTa8Z5O/qk9/NIoLP/PZCpBbWlVyk+ODtH3y5y8ooSI
vpMKpKeiac4tR8DNyvi4RTgI57UPy1+3klSUalo0HP6Vyvp2Kpk27teWpTmW
GmfZQ8MClkJsiW0qxuVSw3Wrwjqy9UIJzSd3Na76naDyXe/cFPAUnb5GlI6z
wrsAYIXgmMauWrr4m7Tle0K4Mk9a7iG97RY048eYjTuVjKaNe6YvYCbbuyxO
xocg9E46oZCAW+L7MEv94H4m0iYxdUerq1lDjBWbsBBhXDsTww3+cMABeP4F
dzRNyIpoHXYuRtd1r1DwLXRlpmhtrDi/K+wzsewEg9ArNHV8k4T6axIlcML1
llie90+N7hDQHNcxIUfKGZJ9v3fphyEY0E18J0UVIZSs7lWEdGQhMpriqhGG
eLOgLu4jeHG65FWMepavPcKEVgpRsmehE1TvYyEp3WMKDM3M8QYu/ReT2AGj
6Cbix9Q/fdAJBKI0FwwCxtSLpTETTWVv1kMeYr9gJLPN7rLCMngl8FmvPzuQ
HzS94q0YjRlbh4XpeUNkZwVUtJ4+nZxOeuH6nWUlazkkK7KdNhpzykPaq0Us
1e5mRkDtGWDb9DqF+R9PcLiCInj7Ngi2pl3W3vQx2iLPINUoBozzbS5S0H2k
ohEPZTLWwsdqdVzOykLFxBPWPeAu6BcFCZHot7K5AJNWR7nZm/WLjFSUm1/B
ChnPLwAhmU86Ip28CyseLEDLSCrA3yMzaHS+JsMBWn8M8QzefFvhuyGLzCq0
vAnEWbGJsnLk+hwIDFrGqva0KUTU0ivGk1ZWbUHhdqCUMNp+09upfhHND4n4
294YDQW9iNsCtLr14vy59LklAaUk1Lbzq9QvXqe+Nb620xVpLb46f6D6KqPi
k9XpNAMinm86WhyT+yk3HstGzgB5VVcjFDpWCj/RI9SM7hxQqwCZAsNfUSWj
ZlK4T5epXVQe0GOBhDbWFUIySTpPpAuT1Ho3CvQmAweytouxwBF0svBAIy0N
D4SacFizufExLl2c4s/R4ozi+CjJQA8cBliUYnQpkg76WPZiqQ1Bju1rcj9U
7//QGbbjVAVld2053PnkdlshodR00Ufk5srDwGVPU2bqOFsReYiUf1f7IXxw
BsdMyIw8ucUO1nRPiku6KLTzPsKUusFLrUULxtivt/6dgFXwJWeutJOj6i/s
D4E/yLjOlnNR1j5KbgV2TDYJHd3/BWyFkXJ8BXM+iVgbzGr8YR8+qHJvPXYC
xOyD4LAzUxzqNoTaj7l9AroPtvqwwwj/EUBf0ikt4ejHMSyXQkWLlRkt3+3X
R2yNVbV/MFjkd6reEV9bZALj2FsKbOnV0o2FOtuC6PTN1MC1tSyEkA3ohLNE
e0byRC9BNdViXy3lbr86wAYV3FJIpukD2OKMUnFR/C5dvobZaj/duEKLH0W0
kcCbWVaS9VK9s3hTVvzHuIL0Fr07KgigpMArTaSMKH4ofL7bZ0n+6n/tduCc
zVW77L/vFpUpmX7bqDz8MDQSlrJwIcWf+lDB40aLsGmMt2pOHJd9ZGnBBPks
xNLNX1I1yWn+wmxeLGmBjFwQJdNjmSCl+zerQC7Lf7GyWdDiCguHO1DLw0JH
/MKM3sFqoLf0JlBrZ63HfZCsp4svDki3Zi1WMkUNK6/k0SyFkT5UH8Eaky63
tvxSkAA1ovI9ELaf6R2TrP94t6NPMy9V0+w1w36ia//1Kon3VZFeoKQwzY0V
XROK0fKhrrZvhX2tMOPlzGGO2D/b0e8UnVIURC/eo7KlEQvTZwuokXZW1iFO
CzHEQFmN5bP2UFPpazGj1VC+/fD31mynfRUnTkVWgRxtll7nWQF9MbM9QsYg
vssJ1UpqB8qJW+KiyrTq06gCrhV3qsvs10Cf76DawpCY82vnEmynspExCDPi
kZelfK1m69FDaVD5cQI56yK95a1t//++p8cL+19ur93NTkyaWt5jaRmgqMKd
hGpNdZc9AKjKZjUg4YWVHmDuHWyC3WHI2xej4EnJdW6nCecWqEhf1LSRyfhq
JJUZVjPVKMOUnzFsWFU2gQnenrjgng1V+t3OdprspMJtpOHQTLjYPY7SIAej
WrXyGUsYZ49xrGru/7JhLLR+sk7U9NZ6hqt2j9SaYfbF7wy5TEJx55d9STk3
TssEgPx9LodfmXCcG8WRtzB8DPrChQWp6xWz2v2NOUYzUAD9WF6Dls9kNSE2
qDNZI748aci6CbG56eDRQRN+cSNkb229IRqyNRIAloG65SlaWt7ZaX4v8r3O
kbclWM3DqsSkY/XW4/qCNre64w8n0dj4a4xJ4I5nRuPn8Lo0o07+P83ZgeJ4
tdzDffZyrCnETSddgn8GeblanpjgRYU5DfPTWTKa9SkaCd8rvoV6DC5CB4uW
MBBt/AfGGhY5BmX/I4ToJNnmw+8ramT9Gk17tC8to3+44aDvRm8QpTDzuo/l
U5Mx8toJuPFLY92t1r+rys6WAO8mflHNCJVhCuAr4bf7GlbDtnXSYJ9smWtH
4BRFYoXzUPWOpBzsExjE9U3f45U+OEOn+2TXB3CP/4k4SgOOAOAIvRvsHvX8
6jorvIcywJPjaJOKRWGfEtBR/oIM/Sd2DpkL8c2Vrl2Q2Q7CVv70q0E+b7WY
C+dabpHBMcu+Vdo37i9yID2P4LEIKGZzOHqH7JJT7A5C86G7B1MdZmSx0M/b
YNzbu0xvkoBa7zPZiW6CLFkgXeHkWXKKmd+L4n9XXZfAWCvtC2Qh2hOhD8qI
kRfxKk2NyLZnm4jJOtqb3CAO3h86O1VMUIh9f0sjdvRbsuX2qhJwr0bVwoLq
ha5SjArp4dM84U8gsMtE+wTE2TPm2xyJ+lIrCluAXrBvML3NoPx6BAx0fDes
iVP9trqZ9CdahC68J4jf4AAiuk/8ggJg58kf0b9yAkWBVZG2iuNh5ZSOiJkb
i6/wD4UBAhdZ7x8gTqciwikm0sd50xcd6Yuovzdolri5up25yoULRH0PLQGo
h41MAWPPMQTlPaSvoZWbdQhqtQ1yK3brUnArSHS6EhvhUbZptcybhhJEs7VM
DPhBqW0yMDzVpmyj+50uQjSZGd9iqDq/wmEVpxwV1Bka6qdCdKGGTOrDIGSd
DdlPR3uVZWUcXxLqQnHi6kalmzF+1FHiSO3oCJDF++sZGuN8QzXyDi7ggpDS
1Ve1kiXFNg4wlbhYHh3WCkS/fPAt8XFW6pjC1F1ulmsV1PifAurtVjN8+Bbi
70/LROPw1gWNU13z1Rb4JrfBZNZ4+SgguqHH2z3IIu17CNb6uOY42R/l8FcO
x6Ad4UY1WQlVcpTyaTNKT4LhzgbaB0UY/y8+V4IYVyn+xj5n7rJFRBfEcaaW
0ECFKjasw3nAtQYpMqTZctHn8B/HBUT26wugRUSawV9CgaKwTekd56y7YHYI
wViSYAQytnSLY9RuNin4F2igcOmvXoC+Ea5YVmLOJ9IsX61keR1ajEDAIVpm
z5zDmm0+NMroVkDBGj63ApyOsPE9A+mEPoRbXVN2Rrs0qvL6nk6P8nG/XpAf
Vbu5ZdLEvIMKdUHsv2LBKp7pYgE7XPdeQ6mnAAGW98Db0aW8RBDhSceLEUJY
kETszW79EhxHUfiS9L0AzUV/E0oXVQyoogplTfo0vdouDqBY/aDGZ75OITnn
GzO/XRjtUwus5fn5UcYbcOTcN3nbY3riAOjireVD6avetbhE35JaW7Ln5/yx
uKFiHTEqMBfq6nwdjvx2FZLN33fwuzqIAxMWGWeK7Vpr8oRjmrEpSSuP/Djd
rSm0F6Hy/qbMxT2/HXx9YX4m0oMgrHPmA8Gu2F/q8oQAD3jqeuWjfEs1Q85L
dnsXF32IDzvrT0T3SWZiR2qpLmZF7wLsoXxfoM32WgwMJaZ+w6Dqjr6a+YIf
N1HzyCsgS/GJXr4JTlkBQVY6wVuAuQvvAscPNAajx6Bc0IE8QzsKQKtxeFxe
v6rLvjviVT852AQmUQELVfqc1p2hWrCY153VSPooqEahYOhpefMsiINpZr4H
xizSui3yKs4xf2SdStZacPaPKWUHIn4e6mjkkGiBCDX6szUesSIXRdZZJuVI
uvsnli1wS4tXan1wXScgm2sYjW1muFZm+W3i3G6zWhi2UZQab6Wd78a1vyJQ
0i+5ZNqqbs4jQFS+LkKoEfNQk+A/KMvRT96UEAuziD18OxdX8V2Z4jvBm7+u
qhRL7AfN6n0VpWSnmzMYwE01WR85ZBf6YfBCVSitCLbXLoRj36gheIy3Olbx
Gppyhhux+QyHt3vqO9KE8YyM9Q+lmFVbIOlXkFhd3Ja3dKPa95Pt/ro7q/15
ePKf1bfMiDALH6FpyZ7j/1JPmggmTYdRMDu9ORWnuNkhDYTT5gayFglQ4kMq
phBkLdBxpe4P9rYXuYMRATsObd+JiAK2NrkegjW0rYprOUGM6llLTbSShFNA
nWPwgBrk/kkjYhzpRyqGgvsS7BvouYiQM3cu+B/8oWZZkvzcj4PBAwvI3mOB
VOjbB4IdHywtr8gSv+IOxrPldHvcwj8PFvhCIPyuXAAM+xb+v6ZoO56hC4Sr
1xecsaMyblAVxc9ubFK118fYmuRIf0dHBsMUJO6sSQ3eoYJVowc7+PtGRcbR
qWxGGJNQPA9q48nQDTBBa/VsJ4dkXgwD7gP+8bqFG+djQtpI27e+Do7Blwhc
sCJsVP3sdjkgm5J6sIQ5f4mMSzX0MbFnvP31C420dzGpJAqaukHBVN35ehid
towo8jSmWs5a7ekMlr3T0X7pM7rh5FGbNMk2pVREkCYJtgvDfDSia8iROJzN
8TWsX/sNqMqqbMhTLVDR6Pl5TZjx8HwHNR5yH1JhwAIwo7hiw8TEx3utDQxd
+TjyM7lXwPSilUppFEI0e3j8EJgC8uId/1RrKNW7Mvp0LsIJt5n1hu5334qx
RAPuzE3o4r7Yh9IN6SIRvGunpTnvKNc50V68WlvB0PaP+A4c2CsnoMFuNK6+
WxNkI/hCBtOEjrNmACAeiEqhjWdXgxibWwn5lJkcgC81/fLNKdHRq4Z3AzBg
zJZo660Rm97iH5EfF9k/MY10cYjC28Xkeed5gK6BCJ3tbIT7pbYsBKBnPOlE
eL75J3lh12YGwIiKMGvpdZ6i01GBfNZCaHfPpd8oowNwCUXZJ+P8alZQ764s
DPiAF4yzicTGWMvc2cLzwgVZlDchY5kedTpm6ayfLX5kWw6+iz+x7ghlIF2G
73sGPHjAyfe7mPM8u+EFkXiOheFFJ4cBmNlD44k9D/FqOI9nKTYAURkGSS+W
i4tGk0cH0yklJu9owFrHeGHhwjuUfK+ZpfQMU+b6VjcN2AtUAO8c9j9ge0NG
gRqaeKHhcWucg46+k9la4J3wU/YWjduXRvttUYJNUhNikuVGomz9Mwto3ZuC
pofek1w+5gwnHVzc7E456htAVDjx9nL+C9nLTvug3+gK5eiI2pXGXpm9SDDC
+6gX735LN3f6PaddlJz9OfJPqpPB5eRz/ehV1eeebp/lCdXz35L0eSC/PiMN
xpwN89FcliosVQCoU0wmwYujQjEQj6wtUNujpokPeI5o6WBTa7+SyN46hzFE
iucCbzhyVi37r/YthUa6kJpYRu0Jn/mNqvVPplqk3Gg5QAdM2kSeXUZV8+H1
dLYbIAucqt/6vNjZ4gMRbLmdS0NqFAhMLQ7GBTdawUSFIiMWUkyiGRsd9D/+
o5SDzyzHoCk2inmUQgSJQm0UHZBOeWzb9sWHNsQCBS7Y7j+hRQgMxDYBfLXR
khdCcl13tEPCHM88DAI6mbUQJYAO014gYsPGxtM3KTG6ctv65AToDRkb3Q/Z
Vg7Jck10uHgQY+NxKHhn9mob1cYd4afp6ruvEtmB/Qr+pMZOkXhK96MgVROz
MX8vfNymMjn7yJTfkSKYlz+tCf8MplfJ2aQR6HMm+hxneHLGvKO6ZgC3ivai
vBJj08ozBOw3XEfg6Ro9OCnKKOx6gVlvUIODOFXodl/62twanEoioSp/+U7t
/7PzBbQa+DnkH+Ju1valkR9Ril28cqT4N52Qr9AZeVjlg/WxuwhidysY+jLN
XFa+AwEK+RzJBo4wrSbP32j5z+IQsRQKuyHoupGe1j/PsqjMpnrUSdYDr2if
UpA/1v1xFWkSP2HO+x3D0XvDI9EJJUgXMzTCOBBgdKnneFWxBdGnOXiW/fcV
fbxyGrZRizFjxFYBwQaQjuJmIOryjgbtWT0tmsJDsyhMSThBqcQZE4y/APio
EK8X9V5hZGLSV9ewDA1/xV5g5fzutL+xubF2YbFPR/aEb8Q1CMhjOpyb5D6R
S7fAaThqTds+3IXABGLnRnDr/QM/5kBqBB75Q7d4noD6pfL3iXx5loxR/j9c
8H1pvciuOD5NcT0UPdBpF8FPTa4vO2vtRzggeNCQ8/zlXEzEdYrDNEYSKFE3
1XUKJEh5K3V2jt2c9BVDo97gSXuKXamd3yO9eBrB1sOVNni/i46NltY1f3L9
6PtIHVFjJkc8WYQx+0yDfyck/fxnmwM70UQ6oxbBTC8/WPPRD2x8MXeoTBJI
D5LYqlbPcCc0if4uiXMjAdhUWNwlqL0GKh7gvw6VY20EJOTPqBd97elc/gx6
YSQD1ZfBhAkVafxupWjMoH0wMuZosOgFqxyEHGQEG6YvX5k2D15jtPuyIhDL
Tj1Lw2d7RYEU03K+Gvab0HYbDnAR8n4Ec5i1yg+be2ieeB1anB1o7K+1X10l
Ye2mVsm548laHiyb1g2fG1ab/TDT+A4zcO73hCsNMyBU+qUOhBh3YAnNyT1n
Aug79D0TuMBPOAXcHsL89AIs43k0DWwKWyjov7lTCF68fdBnwwJJ7UgeC6he
8ypgWaCVsFC81XZC5vyyTkf2D1DVy3nDQ/AskSiu4tH1QwbFG7LS81l47f+b
80250XgmkhT+l1Zf24pIM35FhLWbTvMj1DWeIuy24lNYh+Mp/WYCH85mUhhJ
G3m3Uz8mVmX7Nq+TiiJs8pSSOlwHQG6bVSGsOwI0lkmKimeGLxPsdRRvqVZF
Kw8/uvsW3JSKdPujJkDSYdVJvf6/9XRVKRFYBFFvE9pgSabGw1mzq6bGclZ+
Tw6BkejWyoiJPYomoeGvsRxk2Y6O7gI+l4BZ7CzW00gK5baw9Ztf0LG8S+w2
Fupepyl4d6o3wvVGP+zVYYGbvvVen6CMpTtPaUQRMxCh1QgHbbcoaNgajSVp
nfWO9OiKDMWOcZdZ/Hyy3g/ihWOtZaCXLlvlJNzhrByj/GcmUFx8gsLsSoTO
cHYTzjFa8sOdKAS12wSqTp8Her/JLdbx6a0NokcMv2x1xU4hgXhPqArYjw3w
5I/RHWNlaK/qNassgZs+l1B0FNfjt4YJ65EqtpFi78lp0pv8hr69pPy60ssq
n2MISsM7rhq3w8UJnicTjziAbLSGXYdiAdEqggTOA22TVGc6FE+hBHgOcfHB
RVqkLNbNz/b+kjNiRli1or61wPv9OmgffUo6pau7v+IMTSRHtC0G0IBaeE+3
FKmqty47bTOfgx7po9/7Z4cQmf/y7ZPV89gvovyAhf0dUZcPnew3xl16EYFC
gAV+TGVzrz4Ha8NRvFOoR+6D/xktbLBLOv5YixZaFmGgol7Z2DJxEnQ7k32x
5YMrvCdi8Nz1Bbh0o41qhAuliHw2CEgT9dz7YVfNC6+e+qmsMbhSOhB/4nvF
uRkvxhBnXcYC6zJZHbgblR864QaiMEJFzkAvty3Jx+u7vVWxDLHFfn0/ce/9
iDcpNkgCwj4tXnNLSPRSSLsv7Tge1imr9zAqAJfKP9ojTAb/IOrxO8vXgDtK
EUxTthz6wtwTn85RW0BwHwPh8duL3/6A81eqJxzJn2KyHDtGyE++a3aFezOO
HEopvRArh65ZGzXarGGJRlYpv9UYiFX80JdujKhXMZi9VdKHQuXAZZrzTQPM
wVrUC2i+dyMDFhMQwpqEjS6PSEHQga3YMxD/d7b1Uh+2lvMoaUTI1ABez1GD
8LMhMoSS0ZsdmbPpZxYKVZEkgT4vzGtVv33U6AC/qGkmm0YgRkRdV2ZUI7TS
i82IhU0gARqX94deEde84J904i7yRoa4K2l9jNZxLsYI0Wuq1UWyoJvr6hZo
HXfNpH3VWgIT8MTAK1v4H0T8cOhl5PC+JxqAjMTIbUygQy45VHmYghIXBYlp
U+tMnruR3VhRlFTY+6Hge3Rf673eSOZ0MytSeYy3tal9Jhes4nGBQFwatJf4
Xi84a00aCbfqD89JoUGrOSNo3DJdTR2Vib1rt/iAQ1tpBoaLB4TFr7PyQ6fF
o2FoiK3lZ/Yb4ZK7re3Lb7K2Rhw+UepXnWVs28jba5L+Mu3A1UGyqOQoLKbb
4RHwViWLtfI2Jqyi5Wssroq+PR1s+RYSFYM7oC1WuKNbqp4disoLCJo0P1Dk
cGuPFzRvHdMK17Afy80huNzgR0glTClOAIaX4GZeOgUyde4oQwT5vqSQ79bq
T+a1/rFXb9u8FQLJxhz3gRR4BMvDx/TAfKcTYWHuSCUVBMUD20snI4wAc67b
Nh6JfjAIWV0celGjW6t7O75uqZzClYqDRaJKRPMYzUaO4AAKL6/ah9WHDf6I
Lxad8K1wQvTGXux2ej895/B/00XZuTcyGed+2LM4BUDzg7cFmZLGuePtQe42
gxpf+r/6vGX6hm/ea3FWVKpDcGJpNzi6saTK+UnYFOC3xDJYcE19SsHIRFRZ
mCnimvHuZVHK4dGLhomC5ZRmfYmxEEVzhUpQ323tAuLFd/6fjkEIdW+wx4ZO
f9+2VNIZhfYAc1Zyw3vbstnrcpDBfD2zyVFIZo0H6EouDDMRweFXBj5uN3PN
Ak/MFo2I4e3GTERt0bchmDKLM0iV1XJb3wYm8MhEzDxY7SYuDqCI+d8FajAF
8a3qsUEv13co/CGehExi9gpAFPgtdXkpSbxA5vB1aFpvhOeBqUoJ61h6LGrA
nwyHagCKWjoZ9LOZYoso83/X+D+XuaUsy6pg0qr+5Cyl/63w1WoAV34+Jook
D+zjVinX7hOo7AXEi4VWbBA1XqwSfYqzwoZqiMtGcRujPsJHuAItS0GrRYn3
vCLfDRzvR41bMn1ouJYilhUkQqiGgiZ0bQpW0wHPoTjwhtY6rrVanMbLlLBx
p4vjdvsFaEFsQBXuLoFpPVWxSlVwVWe2thXhyU3nztPZxX/fKEvtajA4hZg3
EzsrqfUDTeMXavRyiF6Vpoqrt4RtyGaoweh9Zp+bmHK0up3XnjYYK3jzngnu
F3wPBEip0CbGVljzhBbOzoIp3Z5sPi3pnA8vIKlHH3A0UTJ83Y2xUVPaU7La
fj625vvtxrlAZY29DZRfZp4hm7BPP8UyKa1ZSrF7tDdDWLiDhQ6R+/l9qP2U
Vyj+6K6zQrh3Pd5qxaKJ3ngxXpczS/OfoLMLv/sVhuafRjFW/yXkMb/LcyLX
/S5sY1YEO87xc/+1UxAFOZ3Eck0ZTaiu9eOe2JlEl1BdAglWX4d2iOWitWqU
TP/ci8Yr9/oxHT8Zj5jSApMEYGiLpgfLKu78ADpyVjO3rZsr70LoIJJytoI+
w2NSyk8lH/JM2wBgJ0fqAt9eNButJpM0NfXrk+8u6pRYcGRXUfhaKgcBnwZT
JUBKphbcgxF+nimbjz5xnVT6DFJsS+Ww+sk7WvDs+sy6+M03EI/r4PiYuA+I
b5fVKqmSmZzLg1sIDmMORXqNKrF3M08woYa0KBetBlx6jcQ7QajAJa6L3CKF
M/hFC/EH2zFyno5NwWWzYhq+fvxaCQVLZciaa0WLJlsxOFDmoxl/JUg87P51
ilawG9jBXzEX3mjvEcEKoaNFmclTyouyNKNyKJyEM0rGCxOBzDEK2beor0H1
bbFmAbeEmpFLH8jT5CeOdjmK4k7EQOVYP7xN4rhV+eb6jrTZ9HG+n+o8kDzk
JzJcogwvM2sbsHFIArJUax6j9eO6+nIFY9S6FzYasn6M1oYe0ZqlTlpSMoEC
4MGj7zgOQyhBw9lv4hrQzyhIfAUUY10A1MoyPNHDoxRvM2WbFpNXA9r2d6Wt
O2JVgZFiJMZeQcq7sxM8tFe06Y5+8AiGOBqMHThmEVTuXTKoOYjzgPqFdRym
/cwXhKX33ZeBIbuwcenya/H/bwG6QlvioMbop05lg0XzcHfSG7eIe0FVN5fo
7nRKu5Uunwqoj5dOPc1eoWD4IUVDumcMyt98CfF4hmuUmK7SCAmWAZ1tquhk
bKGaihfCtD8eFK4SDpzjpyUzw0tZYN7BVONPxEvI6KIq5jKy43wq+XQq6fBS
OMC4i10X6pT9NCfYWp8nQZQFNwGxzLyZc97BK8PQOHkNqZq0hDmSaS1AVukb
GYPX9GAEcI1nYpTh24LAnuu9893QoB2sk/LbnW2ryhO2Td6odzgCD53H8jez
8miGjyowjDAG1KjLovts5J9Q2dJf0ETA8riroUuG1qw/ZFDh8iRwUqXkIzcS
BPw49rj9lHVSnvK6jHcUprgqia+ETQjOP7Oetmun7DrgElMU6l+OLuvCmdZz
f36r+12KPaHw4oh96zBZhHwy/CctmzMT2itnE7YR4gvqIOQM5DMTtrUBnZLf
jp1TvcJmSOyrUA4JwiChiAJpVV4vlU8t4H/RzCW0YDreKEym/8obMN4Aynlv
FlrnWOUZVk3DhesgQhAiDWbgYOvnv0JECS3zLvvtQs5mya/Jjw1oMOCluY4H
DlhuVaABvt8=

`pragma protect end_protected
