// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
t/bz14T3kXOa3fHAnTukyde32x8IA5q/3QgMU2eFPC/JIqpMzPsC1acpuoXO
Ua0BnSd7c5E9CYHFeV6WqGVi5xXL89l2egLuOd/wJHfZoOVuKeneXRzf2tlm
r4LyPR8/ZTph7FgeKvhwI5Ay5vCJBUOxmuXjCbX3js5lVvczSxB+JFaPhcI0
FDhxPdeNODBBaTXtQAeDdtyVIvRlp2Fx1acnBV/DI8UXYja48JrxYQRIgbMu
/Dr0u3paGdBqzw588u+hyiO3VBWmpLHqvJq6qN1bkbZ1dHX++XYqUZRsR3Y0
Q6lCJ6oh5wBA6/oJ5a0wWkw09MzL03FzIx+4ytC5DA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gw2KDoF5fSDrBQUI4MZgcxvgMtQRNZ+ZO0S4pRxoEf4Fk2gKQ3069Km5zZQb
zgjDad1G1z98mIbtMf3FGhPAqiuFwR3H+CzVNYgB6O0bPjAfRaIwMque4Lc4
1O9P65b7Z+2m3I1qck4pON/afFZwftvBiUS1KTTfi4PHW4RY7TEH6EUYuyjZ
OaQJPaSCKccxD/b0Wn3hP8a5xNi0tgVjN6aR/O951FpVOKz3zCdC4u4qG0mg
sGHPcL4x4wkkeF33TKDy8EePmp+NpUTI3TRkpA+J/qI8/y2+ovpUNDFVGLP8
oqO3oCM5z+yQPg/Jld+QDl/4qNUQKkEr2vPeH79iGQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b19bpbOWMX4ZAZvyLvwsC3Q4wpARIC66TU2AyO+BOyXuE5Iwk4NGDrU6hAcM
jxMAuKPVqJku/T7n/lsKiRxcN6oNlPljTrhFk0714aB2d1v1DWc7IxnuNSD9
CEZrkLF5w1ddU9lQ78wxgfs2UB8MqVRkDUFNqdOE+jcP1BRWhJZIUAdpwsc9
IHXK3x4nLruJdELdJpi4aEmW+otBhS9tr0jM6hzFy3kttaSU0llUCVZxfAUg
vRk+EC9dV5fQ3ELT/T72XjfQPr4fzBYZKk5TsOEzg7dSfP4l2YoQjOuZexQO
n6YzpKavcHG9hDqKkvQDTbfKC4O1yqqaGWeGLz9ZAA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Aeb13AvJm6sBWePFxmYW2Ls5ISiibe1RzsqjE+iT0NAib1msuLfk1vn6Aq8f
WOfLwHa+zRfeuPV2lHW96yYUAVImjG2gRf3rT8OiHWFvyOiSdu6a1Erb91Ov
D84aiiCBDtI4yc8vh6xh13C+vVyV0V4Xcj40kmY3pG+7xihYKKI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SLwzzv8Bo6zQH0bEmPhsRYOEr9d0pFj1FDfQ0Eqqu+B5wPf7XnR2wPjjtMTB
7oVuyAzeBZ8oIKb8V00ik4ZsB6vrwOPp0J+E/xS6J158XEx8aXYcMziWtn2e
qRkrZl2cwlpQnmKwT52jKs4W47jbdyu0cVV1z0sFC26WDf14buq1zDgRhL/S
xy31/dRKHnbHPWkoF7nXHVy8YIJADC08HMsgpoq1WPOVio88VPxda65Nfpku
Ac5bd3DcGxLGVAQqK5NH6bu5bawnEyCTeM6MBxPl8vOsV+tBbTzf2k2aide+
n3giC7Y+DZdaywtgfRpCE37fYxSu6FxmwybHzfmOEmweIlG29Gn4WCP9B+Uo
OuJ2Zj3NnTgP5bygwA0WUxs1xzxsyXASiy//kHIZXzz+NIVnLk06YgEezzU8
JcEzKFUvp4OtlZxhTErm3/YBNX8OzHW/8c6uXnA+mUeg4bsqat2cYyMx35Kr
lDqiEo98kV98PGMpbouTMdfwI86BfmxV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fyLl5Ocg/hPTvdIv0jh5/xH29p6HC8hiu8vhGiIYG6GqcNOYbyxVawnyqUI/
FoIdoh9++Qb0YzMUQveDOXBZgL97nzuIfolclGuoZ5DNmE+lsOWAS9x+u++9
0An9oSTmgcWyATzBokB4G5jOA3/6ssccurWauiURbCWN7pMKMU8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fcTEO/+KboB2HuNi/Q+x43sys/cYzsqI8GOrMv/sfFcqrLZB+CX5S5hRtWK9
NetTodIn0zRJCxksMmtpdGXVdFF9dxf733hn9WBdwzlgwJdPdLAaWjM0tqvC
VN8+8RaBqdg8KnXFmRXPBbeY/dz5EqeZcp4ogVVzRZJtuXtv85M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1152)
`pragma protect data_block
uUhmNrtVLBGlcGnofvmx6L3j3xhMlWQUKQiyfnKFPS+H1CNJNzZUw5GyUhqa
BUVkY9hJK9pdQjOnelVePhfbYhiQmdu2NkivuuNx3i8nU8JfdHaqUvrewK1F
BkdhWCdjDM5oVKJ5PwMUjAE/qqr4Il6OEe7gEh3X0KUwvklmw847kCZ4Sqpn
Pb/yumKkjkuhkgu6mKi1xqOevUbNr63Ocy3zuHmVGq4P0bkoZvLfK3pj6owO
s3erRzWyUAFM4WbQI8nH3TAJkKKEPjFPrgzLt1DZt0eXmp2qRq3eblLX4Y8Z
N4X9pVXmgZkx2EI32fM8OVhziVW/ZTtmcafxEnKBiWglU3v1BEg27lqXKCNb
W1oSylZgZzwamtskEjebvd9pW3dDENQb54aAJNGG+0U3lMztcD/8taQQc67s
U4nYnjvg/YCMqY1u7qf4Cn/wYhhFPSV/8IsiOuz2o9oV+RoQGz86XcUkangd
fIhalecN2/gAcQ8YX33yYzEONlCLjgxMTw8ad57jtxIbHLXN/CccP/NcSIRS
1ptZg1J7lGPDCvm3OiGa3f6ERNm3b6aOc2ouerSXgQ4o6zPn5lb/ymPoRnpR
yH8vAh/W4PbxkVanM18admXIX1euwVDxulHqtWAg2pQ4Fn2ICc7UmsBV1fNJ
I3yEAXXQfCKKj8JEHe+PncOLFV71rsUH/waoJZcjr2cN3CjjxcUiUaTfcJCs
UcPN1aXSjMdaREW8HOXZEu55pX1WjgfwkUzZFYclBeD0AJkcElWhFdUPtHlX
A0kPIdYh9BJ1D8g7ADymJKXwzdvAC65q9EO+0Ic8duML9gIiwyuDH7O0sdPo
xLX0CqiHRnH1D8793JCaptjgplCXWEjtiy3CgrNw+GfzZMlCw0g2a/7VQ3R8
0Y5oNNdm0i+PDYRk6iPGaxddQOov19BTuT9z69Y0RX38JOC7kTfx5YrIctJa
63w2Y5tgZi1Pmsw+pVSgU3xAzMb3kTwSsIuOxeKn0BtUmhe+ChtINHhHYPl/
9MKqBInIEZ4KziyWFm9PQt0vqiGIimS1pLKV5gWENXeu2SNENed46QHKVAfp
swt1Q96Y/vbkRa++IlTYmY3kS1tHPFvyUZ5h6pS8IZtJA4gR2WbU9FgDKZVo
+DjRmLLETi50pGSI/lRE0Ynj8gEGsLNgiTIb97LPpfJp4c181bg7GRpTlrAC
w2Ph5W2B3JSpTmSBq576WkGbl1huRuY0hoZ+xygaqKZUvgu24fQI3Rp1mwMm
tXqMczUnkg2ciLPfiv44As6rBLOYTdczKkrphwopxi81tG3MVMRk623T9tFA
KdA6csN757+PGDEFTV8bkSO26K2lIMHPYASBwJwmNyJy+FIWs6u1fl05VLEN
EXEMKVbk57wR2b7hd9m1owdQa+Y75i4SCVEAXwy+1ds+ZVnKUF6G13ujfCxT
WE2fWfvuOagC1GthUkKIY27FknwV/slJS8da8IY4KdF6UQjJPsdLt7HrdLcT
LCdgcBX+nvq2Gwu1mvqM57PqCU33daZQEt3B

`pragma protect end_protected
