`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
ehYVNi4k5JOMDHvkHOV85T5J7AI6+maDv6jqOh6MKPMrEynEh0CB6wIz18Xr+tcz
TDwqm2Z1x+0Tj+5OnUN5APkpFujdfYjgzrDkv0Hl5Lo6hy597SQX5paSgAgu+7Bl
oLWz7tueSud2adLEgQs+pEZf4/OKyfq/7296QZQrRU4=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 5552), data_block
UVtsk7UYFye5xuuLzWmDLO2GGmGrgvCuqSEqdDxVMvjVcGHEnCouOe2jQ9aHHjEM
AD9EiSj3pX0wcf9O2/+GYz+Zjr2vUw9j+JMc91NXJ0MGAyWrRP3IkwvJbomVaH/y
UPPfSUlTfSoxMnwKp1FFWOTvY9FZy8NkdByHC0Eb7OkyvvFOfGo8qD0OAjh+P5Xs
gU31Tx371fwUqL7hSvtVPd9I7Ox2wmSGLpstCKp6+z64fk1UZWFL0kAs0ktUf1KE
sE8EkkQ3ZoZlVcOG9ziU8cLAQRiYLqk5LAQwfV6HWHSPqM9/ZGhVgC6EDcCC1Ybq
b/RNpvNdJd+PdZzd6QxAOtYV+LGUjchO87c/K3575BVOCZKi6yy8ltSGzc1bhjWL
/yMPfvIt+T5kyMeI24njAZ7FHIrhCA8WOFoMIa6DrIiAFrzA3mvY6rD1EAsE310v
cjA0/18YUt2MZGXYLZpTW8orHIq/oEAkTRTt7tmUrqijCn8yyyNnxfkIY/QKFV9c
+jXWlb3PgX96RkEEFeFXYfL2p1fACEz/Vwmw/I5ZWqW4P91I3X6Pirl9Qb/n+S7j
mJUhR/EHnufLLNIuGoQx/zAZKEBq67KDtI0Moax8gc75Z9HDNhRK9sLnCYOgNsRo
veg4mXZFVU4Rvs0hLlX0n4weMnaGbLELKFx0pi1z5Ytdvw/brf4plH7dVT2pWKBj
jrlAse2bwS7plASwMIgmRhKB1DiwpF7AAZlB1lTzRS11P6O9RMCGVEQnyDxcvw8g
Dq70h0mEZaH5GpQSiSXEQniTerZyDycVqkksLBzzik2J05HBx0lzXFn/2BOqI1lK
7DqRMxHeuxEkLWlokQ5pYGL96sWqs6MrQ/bf/5/a7n8mUMTSYgvs3bBOxHkekyJ8
SH4/bhyufahaYW5g8arNH60RX0D3pKhpZz/+X50nkA6X25ElIKtT6tflaEwzMjks
/0Om5j/72mJQ1RFiEV+W4rBXL/f84YNGpg61BrAEbWvBR9dlY+WAtwXtCyMuodwf
p8TX6cx0PvtwPNAkOEheHTdyT2b6FHNRcaJ/3tpo3cEhNSZjL5OGzQ1iOpUOTl6Y
XNTgx2Mh2eQCLOeSA3Ar0A21SwTGg4WV9z7XySrw0fpOT4dFCJFFS1YpGYtMqGep
xqSryOqYe23fLWGOuEjKPnX1VHPwIclRqwAmSi+cBaG33L88CkyQLyCtCmMYa/JS
XTGtBZdO7+4L2gkr/lk/QuBgiBXRO07cjjELY691bGcZhFushxPdSTfxyOZaX9Jo
ZqgbTO2DmihzneZR+a5FmW1TRRn4bqjWPBUqqDm9HMqkBcSwArHjSvvIjmE/hBE4
07eMTKsEDFDiVPoweQNweHXfffXZ7JVs1uNA0C0l/cGLaNFxMD2YkQB5FGnBprZU
14Y6YDFkf0uX/bCqBtYPZa60aScNVwQXyii8/890yLu+Z1WF7DPHrEqAHQccKmVJ
BJoeQeEDLxS/luqssviC+FPxsk35vZ6ga65++pmmWVUg0F5PPtLp5sZirM2CNSH2
OxOBvt7eUVhbmKqZwTwhwBkJQu+9n9tcZ1GvLAHnDUQJntqFKm6K9dBMnCnjfCc4
f7N7x4KmHhh3E/UhWX+xDmL1a+wGkhZyGG4C653EsDUBCaF+GX81WR1fUVpImqxP
/r+Rsq1Ul+QYDqkZ9rEF3Gml7QbQDhxYyGXzvtbSvDg2+uVl/OFnvpUoA+NtJUhp
WvRERVi/tEqDMNgzWCjOjtO1WSnvJWiEjt8qHKqJ4hqtz1VfUfMWMynPIrpulR0G
vMJ8teO2518eZw3s0APw/f7vHSqWeSO7na2773ROhd2xRgGybYE/C73bVLbGtdvE
ZG/5dxUVZ2DC/grcaJVfiKUi2djMAEeqczcZgJ5Utmb2ZrEv2IM/yAtlJFB5RNJ2
n5eJ2yQGK5g62BK8wFp1yg30UIWbgLwM3sVKswJbcBuoNIuE99Y6QCHjnsT97fuC
gSa85M2DrJO4wThddv9DICIt3T85gUvKbUi08FwljYbNLARqH7tYkpf7+hqEmhQ4
PXH4WDIjyAuLxbc6Uj+ldXGr0KxhfnS8Qp7BLXCnVOcdFlmDG4kBPtwLg3XnmY/N
GdlTC9eDU1S3BSE+PuCG6/YkJHcmZRY6+m0DUfJgjiFVp36Fn3Bosd8srrdmAgVD
KeMDi44OePEbzAgLAYuG+SzURWtq+ggeMicxcxVOSUxrjvtz8O1ONsQxF7SnZpM5
E2kay9hm6YZ1o0yORRPsTIU5UALnobb7IWJirkyexeoP2l+Kw91jWLJb3fqB/P7i
EHdB+gPRtw4jKC4geHuCZFhKWchODeS61UUlTlMuF9gjckcd+CwlidWPYB5Z1bWF
Zo8ckmYXKHEYyz9KnDplzqjH1eDTwsLzweUTLIjrEBN8xz3ccZ2PSPdb2Ynm2wNQ
wTQO8moNjwgIBw/fgL4p441oZdS10zHYjV2di7vnXywagIlYeG+PIorgf6FqDAVk
i9MGEouhlCk8w8l6WO7xgkVqseSnctB6pRJ0dL3kuIT9cNxWF4IlczZ88RY8yxUL
V9LSN/USlzbvRhE4s/Ocycm4aWeEPYzLb9a101089hHTQZujV62JVe+JxQ9Gp9bs
TYVPGdk7TfVpapNdsnlZsecbbBoT597RczSQri9bTuJacEYnIViFUwn9j1ez6qm0
MlIgfYnxbTbA4sFcQmJjruXetEkk6zGoNlp8oNdsV98XdQpKneJ1sK9/BlNEkPIw
hd6Owj5As8ISYpeaLCQWViy1M6jpNoDdflHPhhiniTlUp9tSHgzkSXmHCMq67qYt
9+BDC44QvRSW+0ahoMrevc/XisVT5Qla8FpFS4x0MEB9YrbW5Cvq6THkRIFXB09t
JmHBgoyubtDWKCpPlvOlnQUt//pGgLkP9nYeqxIl7pOqIxeU9f+0L2PxvIXgI/KJ
LW4n4WhTNdTCSXg6vdHFq5cMA9yAhalwcDxmA9acn3/o0oLVVb8yGUdUyecAuOjs
MncZKAhf9f4W0Mv9AS1mq21DHZ0PoHKUAYVr5CSnqXesL8HV6cmkeyXTOusWPxJ2
vJiqZGxx6Jv4ttAKORP5KdhRBQQIDO+cCYgWgGp8iyK5/63ZXGh3Sh4DhWjdR/Kv
p3l05/wHr+m2R93d4slLKrk30K7yzNl/Zf+rh/DdtfHB4CPowk9YjiUeCOwK8mtD
XVURsn3TeVB+SJRQ2lzjKbCNGcSymPht6+CLxvwvsUeUhGVklrXtbcOAMNOQ+4xZ
E1OauE3ADZgEBNuQQ6epB1pEsQiu5S2tpydj96ZBUACgkn7g1AbskkDL+Tdr+d2b
bG1Bq+bkadprbUerloUf0Ebpzion7mlQW8iNzfHWDf/v5RTURF2mdvZ6Yfnf23IB
x+Nq98n7EcVrHfsYsVXAB2pVd+iliuVCozpz/Nb7EW+KCmf1ZBamhfrWSfTmQImP
CvdBaNAIuYzjcrNzhf35f/Knuci3bkXXiqEKDKknxdMJT0MZzUViTEeW85YzTBjK
mZqlTMWRzpy4GWn0egngAAgi6poelVrFSXU3vIHzB8mgVUGK72KarMCKsKgLkW73
9yb+poNgcjvw9E0hopGh/wfjEZrSLelmY/op8+xpcvA2GVeJqKszrCe8RhvRg0/f
mmR6mvmiBSAB5iZerG08WgRtdvjFQsm2yxa1xaLCqNPuN8EEz94IvkDPoG8/ZUBs
swDQHo5cCjjgC7mRVGVi+uVnKNm3/675UgYoNANN/WG9Ed0qru5OGY64JjOikVRp
GIuyKYgjwoc+Fqt5MyKRE92CCPqlyTjequ7244YnNYwDwuFjoH2UIs8iR6KC53BY
vVdaMfrgzzjc0psKV+qU9zsK/w4eE1ylYAPps5FwOUtOTiZJuM5EoFYEyuwL4LsG
vI6evu0qvpkUidReKn+x6J5z9SterTtzIp0JzwFccG+qBoZh4CQYnnAJ/5S+BO/I
QScWIacsgSIC5iiwRvN8X5nbfuKY+xLaYgfLD9g3ANsKlAZxS+vqbe1CdBfLWVzS
AvlBjWtcgljgaEA4Y1U3Xr9Yk+N5YVyaNFbw6h2vN95S0PxZQVZB0g/QiCpnxgtO
PPwmlTwK0vuTiNftpTpwaqP47SevCjWQA7kQBgl3CtKstEE+hXSMe5AyP+cQbDcz
vFDxTGLdVhU/fUM6tp7l732zBNxUqWnHNJJjXJ0Jc13VtZtwpLewDfOm1TJF7Zal
pLP+eu7ZJEutEAR97e545+kP+0CLnMy/ADMNJdxNZPKWfo0aWaJZXBnQyyqrEOyy
qp+HcUe1hgmh2VLWMQben9nIEt5GtWxvZavIwxP6tBRS+HsuQPHfq6pQuq6/LK69
d3ghHR7G0LAnvUPObiE6+8Qg3sD/a2MB8doFo+TBmVJ7dbsEAG7ejozoEE0s9Uao
W82iXLDyN6/QH4CdBRr8UtAUU7vYMID5w8BE8sCRDzYVTxcFZq8OHA6PY88a3cOD
2lSa2jiOpCK0UJ9bnkyxHWNsSTmlveVlyJIU1pti0tw1WZMVKmlMAXFmWU4SaGwy
TyHdSQxYbzeInV9Wsw6ZwRrm8QGGyHc6D5zJEiiu0WbBkd/fHDG20w12nwH1/8tU
w3H49j4Hnxt7mxg8B22HzwRqARNQqKrus3qPQjiAQxGNr0teP3A3Ux9d4NxlpdDA
XdtZww8Zwh0Zf5n2oUkpl9S4CNI6/zXR3NCPEeV8nUY/3RM2MvVmLKD3WNfzkAGa
UcbLS/oVjND2MZdyzJ9rIo7xS/GHzJYGYqpARjqZPT2xhWRaTz1v6upzlcEg8OwL
tNQQq5dRDFC/tPwMXGvEOVJ4WW7QNzjB9/8SoS47eJQndg5ka3YWkfoOuMjku8+A
BdUOnkwvYk/sZCusVfOTsAHQyqsLgZUCcI9lkVdtHOyUrK3druFJ5p44IZU+O+yR
W9tmlT4sj7Um5iJrtVaSSFkGXagqJXAItYLiU2OThd98lzlpwXOSrYtTsZujktOl
hDVZxYauPaPx5kaVX9myzlmIugn56hhY3ZCsc2lvEwx7ao2rGL46+o4LUbr6xmam
0HtaWR+zGgsJqfloz7YkYicXjLg5xRXUsPJsnsrDsJ9+0jcOLSVZZNLgXXOSP86E
+N4D3eyVm81L/euhY1BpeH0mdJUy4Veb5pOcq5V3oMNvTzKV0ygL38W73ybVFh4x
+DbxzZfitch88sZglkKn8EN8KBzmASSaYU29WdDIKQd5mP7/ZqcuDLI45nTWL/bh
liztI0TBoaBHO+ZUOzbC+wSv/I9gneay9AMVVzlVshfesiX1Cmo5O8Nja6D1F7nc
rTj3ZkJtD2QwxOda7Ka9UZjg+jkOKjPO/rAABc5XaI+zHCveKdjwzhN1w7RgZaP5
BorpEAXqTFnI79bN7rS63otVfdrZNwbNQVqgU+CGcPF/01v+mNtbI1TxyYNZUndq
iszTZ/nCbCDQpu4U1KCWRjyUF0xJXZ6G0FE8mTWjTTWXvK6RxZw98ocaCTJZFAdU
bTDYSkxV7hwwWO7cD0bC7wptoYXS0pB4kOL0Rzv+TwigLQBNbyGqDU3Rd9yaNp1s
Z2KBBDmVYkR+utQafhjQFVITvQK+R7z9rp0wkFZBsztVfcLloLAYOuT1dwaqhOp1
xdohY0331rDX8iTOuGfx3CZZIRtgNg31BWfGGajpmKD/RJrnbNnOi9ANwyillbzc
qJVHUCk87Rmi5y5hQ99qtO29KHfuQR2JlMB3mCnarHh2gZLj+2+1SXE7vxBjw8IO
XyfLm4boSFRdwthHBFYiB+Ut7ofynm1IMJZBlzvnzSV7qTvgQYvSNYhmsbOISpRt
McWfXOI1E3Rp3HDp1biibjeUj3NgKCRzAwK00C8M9ULXFrA3XJq7ymFJNq+gNWWu
d4xoVuu+Z4VvLoLXf7wDpxz6jRRL6EBtNzurTMfqCQi5wAfFc9JhoSsR8KwFf71v
no3t/i3Zut483lfHOoXpLnZ69lfvQhGgalMiGfazp4iIu3//IUeAwR9dpu1asCLF
kFr/Owhs4xS8fY8Ed4bClMHKxfaMYMQua1r1u5kKCIecMJ9IVyfuqqECb6KKjhqJ
sGGy4DcX/neIH6vBTIgDEs4F3s8hDYHXcD3iBQtF9pL3WIMcG+mx7blHW/klTSL/
ZHzbCkPv9aCqoC6WAEusp/IjoV+EuUZfeasZMrgz7qIjShN8cHJiyJOw/bwAPa9X
QQXN5WAu6VtYcudwBg0xlhwDtW1bJcUyryjsue4kJHlIwCkjW1Sy9KxKAHsq24ps
AXVUc6kb3kaaMRpi7qE91uowxVBTm2uju8lFtNB/dGD8OnXE0PjWE40iqD7qSK25
uFrh7ltUpyqmiiB+F23OtMC4Vq4oRjKOGh1PpQom2fts4UTGBHWQmnAdmWg+Qo13
iCk9jm8HwS1VLDTeXRYFm0dVRYVLQcIBTxINmRemJwISAzW9qgouBmdArQYQ03WO
6joad5Pkua0YjXh8d2qUXLWf7Ju/4U9rmaarRgMPUSuPKUB+NlPwtz7578+1qYhM
M+ms/pQjQaiuMt7syKHZ/NaOIHJcTIUNqU+vwllRYMizGjmBjIukNsbtAo4eByMW
gH5j/XZS3JhYqDZR4gcm7rD+VCtvmRAObaBreVFzMcDkp0TBXAjdM+cLMoo33JzV
OWxwWQHKkLHAgLlvg5Iyta17PQdPhattUnqr7mj4U8SBanO3mFDOjoKmTmdXnXEE
BKA5rqrvk1/rX+ZzaI3fwJmSmllbdg8UWrpV/u8Vlbp2YksVsWgZm8VAtKCAkqq8
qtYTLe9uCj4TGaAfuBrkrWDAfx/iAEFkeTxDh6zpOXpz30Gk5UJ37yEMLyxw4LSl
0KLUx7yk2wQyY/qtwtiBU+kjmbhIkBTXppDdoRqfem/YsAykA1r035hHlxmvSuWu
w+43N3vluak0FQycyAQjvKhxA11zcDz6iUkDvPL/mdCWXe7yQKFbQoUueQcMjrBA
uOomNxAFfVDzw6Latok4otsFGtAbQ9zbSDEBDwQ2FjVuSg/GGkiElaaddIg3YFQN
A5wylOZ+cRVu0FRq2PL2RRHbH/AOX41OH0bZwamDiBtJ4HiuPwFkUk6OIWxlC3lM
lZNTt0GDw2HJqABwb/b6L6UddrI7sjqyE3lksjxh/sq4DDgcnrdvLYmWckE1lyW3
KeOcSjRetwo9n4THFcN3PFgthBBYo1Ok/j8N9y/EUSRrKlFrqHikaPQ+3RFT3/vW
Rz2zke3BWhh0p0+e+7OR59A53oLDbSAjCcXw1mjxw3Kv8qJzJhuye4Z8lyhaNL68
pSRL15+RHlD7S3n2hAPf2SWRzI8u0Q4M5Ag/R0yQ0aZsb18F/D583AOUylfhGGzy
LOoNHxQfBTgOMizhe4RAfE/4vqHl3Jweq1Vze3tpp4Y=
`pragma protect end_protected
