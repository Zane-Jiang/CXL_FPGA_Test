// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
ooi71whkRelO19JWKhzAWeAOPCrlJVLcTpgQ6nOwJhtJE0THsK7OVUBAopJMmRRT
AKpdkpJ8FWOKQFZVW0WxPnhrMv1BACcW4J5XgbpXQuFm9MEiBipAWckNKetv1/gb
IylPgnySwrv87Qa0JPicbcytLNij3zomMxCsZV0FofE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 29856 )
`pragma protect data_block
7x0wxJpSjGJ9rfQcEAQRsajMA9p0yG0DCCjlHecU96+ac73ayr2CN2rp76MeundQ
dy0NwQjnfnU3DZiz+uCuPGex1Dm+n1PUeRvJzxlr8R76r4REfWnVwTUNcxYD3lGU
NnD02TNUTmy7yXvdmrFMrwLosUdGW82jUNQGyxZPyo2qB6tdcr28rfM+8WHDTBjH
aVlRoytrSXOqqZX2IqkwaYmyfC72zoeSxMkxF+ENbNV44bzG+ayrbqPPmWhkuNQT
XZJaZeYZfP1WPa1dGpamMgXsPuUgYgKkRQVt4vsj1pYxF2E4fCDc7/faHM+P6XxM
SQai0x3f/BVac/bOwDE//72pwmz9V/VX5APr3CJnilVJgBKJW7vK4z6NNkcLrzls
vKSIIgEcXlTZTer8db49yp8HwNEIAWOhQ4sCVXLz4lZdgF3Cq4ZEQPjkORPSZv3g
FY4efro1ONEUlR3rQHf8thChe9kEDuHKklMI4L18UUGk4Q3SUFt9CD0GDuZUqo7Q
dqc0E87CkvLEDLyuRtvagnrdI0nC3rCVxJairTsWoE7Ss87oeFgGK8ST7W1Za48V
TtVNgP5vS5+LgiOC1do98f7dueAZjaoVEgbSIYKjL2kt0/Qb926qHbNG3jKU8Z2y
+twROjky7RYbGAsY45QBvtHoHcWH7Ki7r+kuvSgn3oidlfry9vAsnSNor7jXtrTd
4CzPI+HO5azyKa1LESaJbXyhygEzP80E+zaDv2vG2L+1jaip45qBV7xQvjkPaoWR
EEdt9Mjcsw3O7qNzGba04jmUC8+KHzWl0zbqDs5t5fpMldsDWgXY/2IFfeGHrieg
sRyUhHHmYnzas2yr6AtYlPXIjovZsBjWYy72nCQlIn/w72Wnqa3dMTBYlTBSjwC3
uWQ8xZzTN5ATpaXWN7xuKT0yPNH1Vk7+szahlO4LtuMDs2JU6/giCPF5T4Dt/uzx
eaNrwve1oWD8cRDZo+xCXlQXbI7BJh9ra2cceWV/Q8c686Xg1xHHW/UTDOiDkYL9
HlARVmaKMocxslms7yqwLIQZ9VnFFGYr+JfePu5+QHGtVbqc+1cm7P6uimYF/1bK
55+19w71cXatxEnAyLmiafU1NpN/FP9V1tS1750Wv4HJqN6JOXAD80V78fOZoSdI
DCZZI3Waa5SucgNtwu5LkQF29PUypKF5/UOowLVwaM0UldGL0RBRElPc2vThB9PY
vodM4gi5c2VmoRoS4FZdN7s1Q12r/KtXJZa3CxnhMaoKDSlM37Eb5+wHyFzW9mXW
/Vad27n6GOS5y4fZhntnxeCebZAqtvqgLJR/gZ2fq24zHcTuffVbwuOLIZNnSexQ
gMlJzYhepSSSs4YoXGUxd93UMcEuP7aoOL4rGNHljjsH8fjtL87GllK2v0c7xTAI
LjzbNzcIVhKrHIr+SiQ/wqgCQUbPTbGsU2bdum37ZH7uqriVVk2qxPTBFHMmXLkL
dV3v12y/hbCQR1Bmyw1Hc6PQr5MVlqPcU709Y96vQ0LjJDa37iO2+A0w3c211OA+
O017v7+1J8G59Hqa39Pd7fRQQjcSrAnCD1AIFJVT59G9IyHnleBbzrCT8TdCgb+n
ciqrvcdSIvjDrCNKhuyeXRUB2tBx5FXpWrfRZv1wV1rYnUve+deki0DiryF+5YT/
MEULEBRpujH53IFX2+Cz8W8vJGx2Z3mC3l3ItT2vh/XM9eXDnWSvXMIGWH44gAKS
t8B0P/D/GDjRP13TDLC32uXkbP4oDH9A0OIn6j8v/YQwyiLC4QbPWH2J+WJwDj7s
11zuTV/9RF+X8fU1GVOpj/dLXuejF7Nwfb5IuDE2FfeieQOKJsJv9LL9b+19E0HS
fG9xeb69XGDKNJEKf7oUsZvNYLXL2N1zgo5UcGF4++VYNZyyg0UYmeyp94Coycu9
MMYMN9ZlMWWDz3/HpB+71i7sqZZNro5S+S8PpNR+LsZGvaIft/1L9P9E8LmifdlJ
9DArvGSX2qyOB5yefCb6PbruZkKPphrfdUl7aSsVmpt/73IBe0MhxwIF99DhtX0k
85hBKvZepqyF2tsNrvtxzKF1Wof3RSKCKOgCDYlCMpn0vXPJUWO7x5xMa+RrRyYb
agJ5opwxarU6ZH5A+bfGMwvKmr0TnblTblp7VIYpUIhvIC462PjikFMkUk8AgAUP
rStNAKmQpXSsb1oAFBrmqUTOfPt1cjEQ8xm0W1bGBebFxA7D1KrmnRLT0XNz7hek
wPwwIcl2g/lbc0MqEtpeHM1tTn0lulu/btuCu28t06GOOh3GxdrzK49WTWEvui73
27qhdLvUsPfrNwZ6lmp81pjf493U+SDXpVIk4SqWK6KOxAom5uTP+ZzhC09J30GL
YAHYaHlh75qkV8HYS91AJX9SAHnF6FM7YkS6XTKlFv/4AlDnuwSOsHnpAmKjWZ0U
UOB7F4KuABcJ2Zf7P1Qi1GbhUsW72BZ+Z+KGCXjqW6wzq95XeM5B1Yg8oPQq9SWY
loira0Cy+XyU4pshLazyAbpfYoo//GRis8FWHTS90A/YDfePp76d8BNhJHBM9K2h
YvAG5PHaHkmZLuLdZ20K2/SW4lAedc1w7hlKuNuF7kazQGTiiO7/FG9A4y3aI+NJ
wwXm0M5Mlr1k85PdI4RGxt8PVX7Xx9jc/ayKxAwtyZLX6oeKvQmlCkaeoSb2cFh0
wCEPX35uxB6zVJ7rII1kY4AhzDQystB+gTeN2R84m2ZVImuBA1OqvALsPCTLQOsy
GK4E6a7ClJLkeOeRP41arGMLOd0PiZwKB+dE6NVHRolgPNTTyv2Mof5nj5jpbufw
/y7G5mbCadYdBP1nG6V1bhqZVDtIiJTL2FxiKtBQIKhEplY1Qn6pzKk38SkJctux
V56OLO1j2Rmhd8LiPs8kAPK5OIVaQJPoyo6GofNQAA0U1bf6D74zX9eaKgxdIITk
jYvyYH1HyDsCndd5KOsVmfh5mIMePIrEZCqGtUUaU44gUzhyDn1Ol6MNv17wHA63
xLw7I6u2S86Q+dXRV8shmwC7Zl/Gd7MellLfcTj7R1PB3nHK5X0yCKtxEaTszjxL
g7KuX2lHc1R/uEyKGta2DNucPZD5u/mYrIKj37UV2Nyb4UhdPEwUm162TJrgq71b
QW4v4QDKG1Vfv+6dZJmrr8CFRu4h55yemS9wZd7DFQ418ZUeb+xQZ60PjZog1Q0V
l/btG373UKZdg5B10kn26yjRe7jiSC+qFs0MUGAp8OQ/opBtdNXeBI4C6vmCAhv+
Ps+RdeCyN6lPJo8gFCBofsAjBCF2VhkVTnz+WZxiR03PNxj2e6V2C5dy9ETg+lrs
UCigtQBvzifc/4mWksSM7wdqef12EMCi/iNONlxmpB+9MqsF16Ln/Cw3hvRmcxVE
Jy41PTTMxg2Iw3pl5ULp2IlHpj8YjzqjT3Pqqb6RLYtVZTTxZpGLb63ehYp9FNGu
1dc8eE7dUdrYEkW7131Nx1l0wkgSkPUxVJ5VYrYs1FMpGU5hsiSnTU7VQNcILsYT
X4wP2EgzvkGJQHzeGkHTZfbhaNipTP4AqR8R1I1RY7pL0HLDSiIQ8sRMmUoyfJs3
DdTldxbVjHQaeAV0/HXw0UOHthFcBeMKeE7xiUDtrnN5E1jtrz4cipeHnkPz2f+Q
JSPvSQAD/Nzq9f+HXjMeq5khO/D+nQDqjGIKztyGhYyZO0GpvHIQcsrRTJr/Wq/V
rT9yKLB1EdJk6RYr07agzr26PRTBRUrRGr+cfF/CjUjCXOlUtA3/st3ffU/0Aoxm
TaCRQVIq59tivhYAuSheHsLTZ64PahZI1TV4FXUucWZM9YLyKGnrWFJYNOx9erXr
7BpQfG6wNY7viYlZC8QiJ2d8iCG+jQI8WftbbijWyMHiHQD61XbCPPSJedh8/ZNa
v3nRZkqWaVFYNSYHc8Vb+vvrvtbv0lxmebphiB3CCc3IDQVz2EM9XLltY0tk4HfH
bvTasgQH7qpsTr1mqp72qYy+PMG+93DT03ks66hAh2fat/VzIEAHdlzyswvRewA1
re76zikoA8RBQ48cJZJPsEjPfMIDMpiJGwmTF2a8CHld47OJw3EmVFKHybDs4QEK
ut+gyYvZZ9Vcqr66J97HgBYlPjK9sjaLMIv02aTV7Uo7LaTox2CSfT2DJPdm90VJ
wIsT73qJ/AhTiXFAb2TupIK+/Io4wsPG6P3n/D2ARh3PoSfJmCfCIFoj+53S1Fie
jV7BeFnZ2HHQX/UFZXRBo+EzwwDM6KdRjiEWyJzoETbKIJud+tjY2ZTuKUS3kPHy
xqYeRFGuTIdI/+N39yCHgmn5arQizT0NK5aS0Uo+Dm4hh74fn2yUyTaLgqRrltFT
yP+bzDYdLURoN4plTIibYtqX5/jfrV4t1KAZ41cDyb2MxaNnWxk94xxBE1dPMZlU
O7xmZooN6t/3WpyRjPbOyUgvh0rqpCQ/NLWIm6GsUOztTwsnn8Tl3Nh5QAzNKF3Q
gwfO2eg6GBjEVcj9+pWNjZtvm2DXeXx1oZ6kPnsfVMxTnfsHos8Sy6Ei4f0WXo5l
FIoFix+KdziiIkNCmatvd8ZZjOB5+ctc5Q3w/JBdhZNCG+mBn/OeQbcCE+iPkHaB
6icFY88AtuOhW9a14CpHk5I3QRZ6SgchUH8lQaIl/4g5v+Axpg2pqN24qfdNcyO/
3Q5QPSEuo7ltYpYe/00Pu34QwJYy46a0hd4LoAHmHNmnwq2U1dhnMNCMyy90VPHy
oBbsTL8pLYa18DbN4u0TYcADrrOoneYy8r7x9wsVl6VSmhMcwqlpmIo0dSqJbigo
e2+qWaC//mPJrGkqpYAz+/Hyj0f3hYDt0+EdsM5IQmcJsmvhyBl6AcS2IiRt/UNs
Nny4dW3C1Tbln3BZ6FDeeiYY8yYtF7QX+Jr390wpDXzepINp6bcwCbjO2b12YwY1
GK1oQp0L8pUQzY9+SjrnvRgAHmdtHSMdKCFbxYVmOgj0c8EDNlUfyUdhqeK5f3wj
/1bI19KwAI+BLIJROLYO/f9nZSHRluyM6HO8C/XMaNB2slvrmMo9n95iDkb7XoEf
MVUFgvav48CD66E87AVbM/Ag3O3yARLO8Jw+W0LIYRswZSd5t7qfpebJz1gLyZS2
fHLBM5/7jWWLD8JW6rFFjBV3iKHylcLwRdhDLhnsyGH+iEkeqP19CYHaC9o/RIwx
h8t4le/Tf8tkv1w2grOdPRdXKWUP5nAsLAV22vhm4wYmrfHp52I7yoyfiD/7NuER
PpeQdshxGx7YBdqLXnx/Hn+fHCTL8AqmwBrwzetlLD63Ew39Ni60wk+v+oQ2Csgd
wxPEWbd0kI60sszb3uDMI4aPTQ4x50XdOn4adgyoTHjPesJgJCui0AglrudhOQ5x
kSab41iRphzKviHfgsLITZwowLJMiLnSrwdd2Pu86y5MTmtyNNv/+UHdK1t3o6/5
wNu/M+IkwWtYRqKYlfVGo58sI+RcI0og5YPuLICq0jPeKo1/vTC5N+zHTrCgRu7M
ebvoz6FvfUtBCrQu+fz7HVo019StvAJeQgQK+j5gmpIYJh6MzkKJEwJ9HVk7TUIv
fl+BaVUM5SQKW4wtrU/hn/VGL6qhfsOhcwfaTZFHMYHEQ9/JPwszHlgaQQ18e4O9
BYb8DhMGPbr8vsvyIM/vTq1AIryfwcMZFyZSfc+/UD2Sn7tum/ZScC6GBg1VNcs2
cE/XWkkWePBAdsMHJgV6Kx65J+5MsE2W1s9GPVsXoBvIRUQeYZzxx6P/CHen9CVc
SWZUjD4QbptUCGQPout5lECXYZSIaN/BB9LG4NF1QpCSFA60oRF9c6IsoHCw4/ej
LwVCeEWFOOeHMkoVTHBpaOmKWXpMS9wmDxigVDYP3Tsa/ZMkDlwAkQ8PeUrSDcBl
2ebq49VsmYrvxAJgndajPAsqKw2+2BmomHUyGkYvE3y5sqUEjCMfgqiYAamE3uZm
6u30j62sL6bcEVrr74RphBIp489CSnkeIYdTKP41BKKPwqeX15JCnv1/qcCOO2cp
SNoz10XwrkbnM1csWp7/OBMDy4gYhxYhsnEYkirofJjcof38bimeYVucQwPc+HcQ
3p0oYa6Z/kZODu7L3IuwhtF6Olocqa1sF/oUcd2rRLjgzyaH1Mo6m83npapMMOjK
sLekADkziQLbcCu1iUUmWQQiqBM4LgaCH7AQ3O1rkgtbUXQ8l526S2U0JejecoJ1
IjFMhm6TG0Af9jAbfgQMc7r1QFVQBAxMM4OjdMs3rdkql44waHcqV99MTcYbUXWt
k+X0uQxdn2MkkK48o8Z6yQztmiNYa96jJhOJpldG6zOY7DuNaqS4srbsBeGtHri+
PZABB6/LrOCbgLCSXnNFgFnCaPS8r4QBHB+upsiEEA+0GNKFLHFERVWGJ6AT1LRk
jqu81h9CPrB+d3whEhPoIIsWoory5oodweQUqsrhNuHht8z3WtRcszzqxlYJe43E
Km3YHJ/hk5+ZnrFWijiQAA63DrU2Pfip5FYFadee7a4hsLAjvN/DleZTVGK+yHTa
RXro4PmuaPShEMiQOlvh1NEnrwrz2FuMSmtsquGuoCyTpqCyWGEpF6lcwCgCO8yc
26LzlPGM33Yq6esdi22uJGgrJ00pD8KEPEzk4Ru8MxZC2zbJpffvPc8AIjHbzsbi
JhA4YaE78HTLpBM6puxEdvZ/MoMIzi3nJou0/yROWaJBfNhUB3u3y828QC4OadsG
pI9Fa4g3fwrWOrWF874WFW/odLL60n8SPliHvyCRasyWkaqg5JjZ8TByVwO1kWRy
knIiqKSIIcE99jDP0ewWJJI/PIsli2ycXAXNVRmL6yn85KXuemRNEnuog41k8rUS
W5c6cG6xeSs1feqnUcMtTh8QYUu3/AZ5jeJ3rob2Njr1TzLhufnERbzqJSl+pFCc
O9H2/xdWFTXH+vcpKzZ5jHii/U9Q0K0HAiSmYQJLABLr115t8rf6PttXXTyKOx+1
20JYpubg1G8dhWfphyHH9sVMqHETo38CK3bEgW/maoIH+KkdV67zBRiT4XqO4ah0
KqzWk2bkq7DQ1YDRTOXkgHGq57+RcLqg4SloBk1tB5R35fRZTRVOWulokdvqIx1S
pKqpfhW+Kgf2Lp3uzS8jEX8ny8mUZKAXblx/W85K1e5OEH+HgnASvj0oUFR6hQ35
MmmUvrG1Z+G2FONR+J5dpRO6eEOBfEM1/lM/s/5m6KPso2LG3LzxLpKk95cL2/HE
ZjL48c5BHtrdjE5kJ99ZmRBNk5VpDPe8OnjKk9C89DqirNxXszjbFIzvgJl2sXUo
aG4vvR68BoPybkQX6y9WbbFfJwWMNTR+ADgb5N1a4+P4jRD+mh5wB4wATMx7rSkK
HypjyzRUBOxFIld8z2j0ZLBRR9FP8Sb3BKkBcAh37FxfoOKOkTi15MAN7xEbjNGQ
AK1TiUEFr7f9Pts1vyQchMEOz8Ocn9BL72nfJ71Lh6S4oEnEa/8DFDJ1Vczzte3l
1GJCbn2TPLb9NrHwbFZ3Gr7/Z5AEtE0+6BHYkBfFVAIs7gQulw7A5ctJq9bkA0Hl
e7GXcdjQQCJrsIuOLspmbug/TtscdU7/UMQmGDzEul846Wmjq7vmr6SPGRvlLTtA
M6ewr1qy6QKO6yZOg3IALcB1xdmry380EpT0Z2i8/BpsK5ToaOv+pCNH98vjnUR3
7QhZ5D1FvMue9A4cdB6/hzyDEKF60ROT82ycWDHqPWcpkhbZkrqyg4BQHCogOeKu
8A2qmFgTWUkltEIn9R99u60lva2v9giXDFWp0GFMtUwEq9cSRLV2IJ0O3p1Rq4Wl
FRTjHcBuC3RIeB2zgVgeejq92R6yGZ0gBzqVjwDky8CcHlSZai7cp/2h+nv/9L23
5ysO239NzdvzEf1GJK5a1f1l/0hhKFTxac8mc9d129E5tgar7p2/rEOaKM4OkezG
f7o2L0UT2tjdsSOeItna+ajzx8H/flrU9PzL1MZtP938dIhsVEgljKP990y7/HtB
I/ZslwtrtTtYx5Gj40a5M3M4J/UPm8x7gCkk4wmxPIIT6QsH0ksz2pmiGJyUKpHP
MYFcnzZt6Hva1MRR4A85nHTcL26/vD8vlj/2klUVVB2T/8l51mG23FI29sT9Nhap
HcQ2xTV4VrcNqBMqIXXJTz2Dcy7/y16rU01wzsaqgRj4hHHkspCcx3ryJLmRee7F
bpGonFnWMIcsFRlDaaQe7bkOGvsc+Cylrts8wvREmxPFMKnpmCeojf76Qh/ABSp6
bCN4uYszDSnw6b09x53CPeG+YALbGJ+cOz6KRfOk3MQfBRhnVj5+rih4fGcCVllE
h/hBMKDyi7xx3irruPPKoWDADPI246klS82jKAccZAt7jr3ZFuqN36fE2h9PVLMT
YUFhqq3AkdxO9pYSFOy81pEnmmuvyTz7cWeCaTxRA3trWnvMz5oZN/ayVQySq9xe
N2o5/VCqJZBTD2T5Mhid6bO9xyRM/LSSXspVXngVwn4kQhhDonEuRRF4/QoPSlcv
Nr42yfAW28vsqY8K534EfcQMfRjZgqHAapz87hWnLwB1NIsrJnC1LvK8CdJros2C
vSJx425nloGJBoI3Dkabxj6fJ6aeil++UjCYXtmDRNhDyDy2X8FWUuIQhWfZ/cvE
1/PbEN+bH4hRNqq8f/tdZJQFGtxzl04K/NRsGT5HbAC+ON6is2WewjWgFRLuREzj
e8tNABVH5H/YLEGSDVdNTkUlIuwS4FerpKe3oLwNzSh9edYrHw1S+jGTrWSnBVLO
zFHcneuErhqItHrt+6yeVaiaV6XfBk5ATMJwGL2RI9MjnhZm3rKNxtHVbu9+/29f
vQdnmayCkHYlOz0fnFUe3/oW/gJLcxvlUkAyuFwto43xjxtcN2x6LSmfMcIBeNVq
4f2HpAMz2QuVFamks0pP92/VP3B4Gj4tiYSzB0WbyzZejaIE4uhA7gzvmDtMTTr0
te2nWmtZauoK5+7tYkcc84VcoF2cxhGKqXoGv46MVJ+Ynl1z+K/8G7uJSY+2Qx3T
dFFu2mqTH+xCqpTEpyRLl7jkhi/3Qf+xnqCCnLXzjefSZOmDfLkeJTGzMagecTgf
wXCwWMAWEAM2j3smdZoel4ROh1EUXCOUDmNKZtEr94ehKVabGNO0na0i7N6+uhCw
uAJtdx/zlIAnbjXe9Q01Tq2OoVl+DGOqbgnfhQBAAUnUHzqKvejLYliPOAQ7Y1eC
f/mxN1jo6MQKKHMcIPLxs0LjYY7ubTW4jrtkHjJubzbZ8fxIFf8wpp/0/gew9DQd
gcyJ0xCR6HN+QFtiQ+OS9s/deTz0V103+5j6oT1Nu88YFoK2Nt2rfd2z2v+eFngH
io2sFH1jnFKpMhvPnd5LEdrqPfXq0y4xkDNyRaumw3I5hXP0BfmeAMtcd/Qr6oAn
HPlbJCCwGVVP+Rb2xpAiHKsIwfHL875EHyKzq6xHn3obUBneIklIgBXvWQdi81+K
T07tpoDFlyq1J1Oum5SYNSa8okWkY41Xsvr4MSx32g9p6z4DnYFK+DLm0xgrgp53
q9bhMVqHD7sNhAyBNr5q+wQqwJkIGCFNu9cYxfQCu9dBDdaDRBvaElmEKnHgdzMu
DTy9Gm/CePOlRh53exv/Pf+l2VbMBVtteNVZfpgDKQExp2LrKVx6lJYOdSy8Hoc5
DoANcDvm1u45IXZXJsDEK++j3X4gTv+FHYATuD5BvDONzQLxsxrkPLIi919Txeht
43H+7w/I8wCPERYzcTEz+boAu/rs209KnWtyCY8v8+tkIJHHAXY7XZ/OZK+k00rg
4ScgWi8PPdr5P5WQGCAacujKwd+LRNs+ywkIDh8+TQyDIs1VPlQJHKk0fnWEx2PX
5C0qlzRsNR/TleyUebw62Q7iTSA+Gp6DBCZnJwc96a7R0rKAbcB0uKDYX1ETtOct
woe4DaLIHUlHmEjQ4Mn+Y6kXYB6cn9AOCeozj/d57KYqij8Ua+anb5y+99Aa/aYn
PEEoeejtneyM4yH6Ba2svWbdQQPjW+9KD92R2gvz/i+a38Ek6gTQjxNhButldSXP
p9O9bsOUdqBI60LLh1vZtZq0t+G6W8vdrxbR1RTrExmxaAtJMXNIKHizRRpnH2vb
/RNO0bnwJFXaq3Anr+TLtrs2PbnKyf4q9a5dcYmX+9ABdJIX2YrxCLGGvluvt9wL
Pya4t/Ce3C5gn8yYzqW72ipnd/eCjtyNICB+yH3JEyfp8kHgfmFq5L4JubuXu+bk
lIX1SJST3BEa2stqx4Z6WGUPQO4uiY/feMFXjAgO18CcOO0zXUa/IYv0ukV+hBxM
G7wNsr9NOFwu/bYo88w/fRzeY35KG+6fN+4wq/ugDuyxsMbHvskpxveNImxvZBdV
lSut7ZWHf0jufKpI33PxznUNDdYbZuuJA+aEde9jtXKECdHTCIjK54JuLk66rqUM
IjcXfHcpFxrWXiL462z7ir4UE9Hui0hV9Mt4VlZIdNZFcS9XwROHaXks5jTuj1hF
OAdx0Z/UnzWCFK2CFzW1O9iy7jwJsQy5wF3KB5uLqb5H1qtnpXect2V8YaRIkWuG
lSEwzXKwfix0MDbU5SHfy8bQHlzRErOk1X3HwxABlzMWBB2ZVa4mCIfvlL9Jdaui
Ou6+1UVX8doIpcHYL+efkvhVXVxDDhYryMjKK0Xvn9u4UGbJUfId4ZZlGOt95HyR
YwbUhQ+60R8FM2NOHB71WUtXFe167Vl9cGEARxXZP2KlmmV+6QJ9JOg2PlFYYZ8N
ej8kSu+cGAhAV4oayoiUEV6qekXOFoXDIuJvZ7nE8addf4T3cfbWEoBgsRlU2Ndl
jjPkBFMCCroWiwYkDW5Muq65kzmTGjAjo5AQBxBMCrZgPzR9Y0jmHhk8lZjsjFNs
uH83ugGss180ItEenN2ow5792ZYNPf5p0O4pIozYdlJA6Af8UmiKVhKztsJf+tuG
I/nOMkcRnhI6U6X4jxKyQhgxtWJBo3eSsiG3/eA3dDQ/CgCbAyV0S4F9Ndpj7R0c
UEhkvu3n10kP7fmzTJT1GNNAqBykXLsU8eUdPFLUmKv+UV3/r3aeEIayml0lshOp
bp+F7l+ZNwh4LbQHveuMHma25nq1d8KFUWqvBPjN27ZsG1Bvel0MREwCR83+Htv4
gjwtkhRzb5qmSG/lrOZf0gWzQD0+4mw3gDrIV4ceIUHV4b8uw52JaiD1vfAPjtwY
mYJaLlSESwg85HGZN/dpQyQBAwXBw5elv1gqRoO3v0oCaqsG0VhWOqSNSLgCi4Fw
KK7chulJPPSHeywclLyQjZtwC5taL1YwRvcaUhzrOvzzo1Q+nWGH7TYPdIqFgrw/
o5iMOK+Vt3WnvbVZ2WqdMrWwfap9zzJQ/ZYuRqUWexyK71HS0nca3bPbDmt0av1D
n2c8J09vYWyBbslgBkpZ8DD5dNJbSREZFb+Mlpn58UcbxBUHNhO74V1rTuHr3gG2
09Em0ICDQU5Ww9qYiWqVRikaSVlRJKRI2r5ssrvVsVNufhjb/5fKBdPDMB8iToRp
koQhEMCnBMeguQVHFzPoZRScJeEloCqgaA4iUzs997imDUsTu8+GE2j6hm4lbhFI
CLi2AJ391Z3FsmXzctV+jEJrZcVDmNDKEGXKo/WpyTLBfcl/KSkKgRUT7LEqrSjV
vQT123nrTifDwU81F6Si1SlFXjvUSdqeEspDKd+sOdR7AapTCdBQQ/4Xh7ZXdFil
AwXsNZ5eAySHQkLbpfPCvwS8RWE10vr2Ta0g/PyU/Xcpv9Fe5VsPgsEFL43CT/af
BLqY6Cg3muAhKOXiXW3XmyBL4WZn0pe0+ZUP5BoEcPOL8o6uAjbnARXIl/n2lxHz
33+v63+YgDMy8inT+DFMODvCpSsqLR2SjkDMYsqwyuWark9XJgf85ZhIIRb711I9
YKwlIuoafRUOa+ios9+Q3OyoQtqW/8lpzySKVhp85Ek4juPWZki6/yt1Ln/2b7s/
CpZUON5MJZU/zW+0jcYBIZerwS5PzsHbIhRpRB1q9xOtyX+fyTNDYFOnKmLs8Rko
LZwx4IMTLXFtly5ngYXEwLOKCzxixMrGxPLb9YRa0v6mXTGBOFgW7UBw0cfnOWWb
I4kcECOshQTL4fSuDfJGtdq4XH6Ys9OXqCHC5CdqrZcadyhNWN/lf7xRrRHNlD22
xRrOqrekFlHI/Scqtash5Bcvks5NGgAPq3j71vlG27c5IPO8y4Gz4yIOVP7y3+bY
XGKcS97oM/dtW9wbt1GL7OzmdgVUr6UAjN2ORv+VZ8pUW/3cVRvn9VHGbybATTch
9GUayi7yqobmjQjPWNtA5hJuD7oxjatFN1LURFJScZ8i8Ac3wVrcDYs745D4PPRc
WSJW8osTaQVAiUbU88x7qT+aQwjrBJGbXPO3gwYWXYSUQ+/XOUP4ew4E0Nh1e8zp
oMt9wU2rRVKtmoXrBUWkYmFggXm3WGIoGkXQtvx70ujM1cs47exgODhcgLRd9n7s
9n0qBMpC9L9B1hfxqv3jQNg1KmNvugH2JSmnppBhkqzzmQIXT134wG9FC1tZBHEP
Xpcsfq5NvW6IyDkMo8CVmEMVvr8cpj9/Ot0TjGDpFQ/xIJRnxMMP5+8nIDSgzSCl
lHjizqeAA3WtyIGQhcwoLRyVnL4kUAYBgGW3Q5eemyikLESCDIgQ/UY5LitzyLbT
SsGpBNiaq1jJI7d6kTWIi06GEufVix9FsDxISFjhpnjgSRc9jU3AmH2HEoZJcQw1
e7XP1RjPrb8ePfOqgMC37qCV6jp2kuEGMR498inLo2ZIpCPpm6pwJRjRvbT1ColM
vssz4UUGTJiT0WeI434EgInMtdogmFod0CNuc5UVkYQxNi96vfQc02+DB03KXuJD
BgGR3OLmeMOBOAdwDdoFDgG4BxYLCldXVCxBuKAa+j8BVPMEjzZgCIlc/4/OZmjO
YFk04zjUT+jev2YuSJ8QdfFyCyBjniS+d13tChwEgzxtg5vRy2RHyJv2iuD4dJtH
T9EniLT7qiO7MsN15I4/u9wC77aiK47PLHH2TehoEWhd4xZ5js4X3FgJa4ydWcvt
/vhPnYfzu/Eihkqq0Ah6rZ08J3O7+IAzdbXKWEDPo1JSn0ZBVklLxOZ2fDX+20sf
5ziYEYKsnMYYQyALho9kVHTid77QRW/Rklq4YXtb7lmyKl6vnyrOLr2xjBhZYu+p
kCyFpxhKZWcoI10RmzzUze7/E0SzJ2G9DxfTr5K11f0/9+G1RfbMLGdrT3V4v6S/
7HZ6vBVGQt1j46LLvykzlDz39a0vrVmbRrdI/ju4NHkOBmfY7iwePsL7v6Ero3yU
/zEQtGQ2/2CPSfzZQRwrPmj8iiu13xYTr0WNmUMJV9tYGf6cplXYMLt27VZQmQv8
nXEh4mlRggrPUhcnm0SoP2I8EX0BdXNq1LtCtc8p5+q8/0T3GQ9TXyLXowfuJV5e
aQa7t+QcM1HMWkekOJ7Qpb1OWlUwy5Qaqx2lA1u8D8sCvBCbbdSJzhq0WAgszKdx
/1mkUC182nsDb43Pxqotz3JGP2/z8pPyhAWDQi7jdyH7hZJvYigPO35mcmytqwDR
lzh9NVr/g/A7jVipOw3pIDwg8lJG/T0nZsydRmzaDI71yPah8PckFJG8PiKrf8s8
/d/M3eOTfoc0f9eOqYFzxz/wavd/5OWrU0AUhCbDvmu/6ZeHp4AFecY4O772PU6O
WtaH1hg2DjDbU67QrgAS1qOcaptcoVdlggxo5aGnreGzmDmKXCbKquhePwLoa8w+
PSp16+n7oXH3G1qlwonRiO/LcIEmM7fXnlNGcVrTzsII+RAFR0/FVTrTlnwIMlix
YjM+2koC9k36i10PwdUlxPXRxhv9Nq4ueqYQ4UndrqZc5/io78y6wqppiuxBGd1h
IzegPnH8j9vgJrgo2KApm9YP2ZjcHuyJYyQlXvPbCvw0q32kM35AQgVRmHEvoIjo
sC6m2ITh269RyMvh4r8AxHPrc5STeEGhUyZxGXYpKNW8J1Juo6mnl0Xj5eQqB3cA
9+Q2rh2PAL5Z/VqQQG0BgB1bRIQQ214K0V2rzvmSrmJl+NAmZnFlBgyLoKRQXiRK
9daQhWsCcKykzJJxbB9iz4arSQdKIB6ftHOihUGUvfFV4Q4kjC2lEQb+gs25X5iT
9t+AqkaH/e2GfMOivqYIM5sUKibNBXp6z9cH+MFbH+/wyET+A0PkMkTf8Y0YFxAe
LDb64WoyUi6dotK7vVLO3OUDh+rrvdZW2PsuI7Ufmpsa5+uEt5H/L97ahpgAouC4
0Ngk/pT1p3DM1RbdtPAX4OCQZwNXs8/SZXXhk1zaxpQqu7gVYEnTGioY4rDgmFPM
HnN8vZSD361F6g7DyPEfvhU/jeC3yeEP44dQCQWnqQCHbWNECmbsoJ0KCCsEx0Is
goL6JUR3bPedPoFqoBZyLqKjacGf6L2H30EIEb5g6iXP5McMwYbLgFtTSdxPHWk3
NOSRofzhVSovmy3VkXwiMq/JVts03RrThL34tk7pA61oE/ak1K/JAVI9+oBTmVgz
ur6AxTL+Rd8e+cDOjkntxT9NhGLbaiGujjO1q95St4cf4Irzn4Ifb228Vx/XTsRS
2ga1VXZiNFuQjE0MBP5G2b3PlVPBL8DHIZZo27lUNsICTTn77TtW4tLcL+NUlWZf
eYNRFGIv4M7YQ2KIml6A/5Ez8NrjjT8Ca4U4csZD7L22i0Z22u6IpxdZ66I8sMG6
j7RGIDHF7CwzcYrqCovKQtfthHIpBPbekWLGEL/oxfL3/ZJT+VUlkRQPf6/xKLxH
RGf7wU3GgkJeo9idtaxytrg0fHbv0xzIDS7cJoSLH2Ut3LNUFlU59Og+3r2zfA7F
RBlh7gZa7TbwUnfqZnao6LYQFq3v9sBmnrSN8DIjtV0AgXVgF8/UrvxfQ+q3wnHq
nQHFI7ftgrTP/xfC+ZVNzpq0sg/ZwP5A6xx9xpEcGwaCpXXqspYcIqdEapMmDmh9
hRdn/jTFadIveMlllAUNXPBCjTfPfcoFQ1jwZyg1O0jQoVR3qlnezCRhxtfE+Tag
XPB8QPoE0NVrM/7B1GDrBZK37510xoL4k26SUqzuDNMlE6LK0b/9r/2sKVXjDb9i
p+6QWaFu3tLSC9xgOrhP8FndbmzAU58826bQt1NPN7xWgBiGIUwL6j2RfcPd6zWP
G9RjDr/4zNE7xpWQMNF58G++u8JgFK/KX0HrbIh9sEwu1LIVTxb5AYAwrCXhSUiT
yytqZ5K0mj/5OnBsJhfjHcSCwrqXycwNedkhswpeMVN8VRBmsjk/Y/iNuj55/m08
TkJK4y/sJYYj3PxfXa1OvzVQ/54Sgc/L2z8dqJD/pGbTBuGodO7L+APYh7eRluYE
pXMDPmUjS5fVzpEBLdd/RCvPmLQW8XDk5VWPQqFutw8OobMrSFHmmfsNK/BYF7xy
c+6ioIWFUSypiAI1nyuM/WRUShSeLs84bYcBSfW19+s6a8tqBVboV0b9EeXLUDVH
w+cJf/Cn7UFu1KZ2X84FFDiyHbazOepqlhfSLMUP+Um4C+tzPM+u9Eurg+wxFF2I
lDro1fU4JOzf+pdMf43Cgnli1esgsFs66yX4lABlXTAKf8Ojp/DMuLRqCkDFRJXu
4Yv9dPv6zF+E/FVO9zpgW7rDWIXynnIPw0UM03+VbcvoSCbvD6msuOZUMaHH/nt+
7y60ibs9Xjrpu0p1QIWZJkVXw2u8unIqWuMMI5Mp3KC+YaCROcgm1PccJwTXPfVH
B1klYIYcFTJcyRNhGdroyZ0su+GeVbYiBSkyWVPlNgUxkN7lCcPMWraJd9LXb66B
fM/6qF/3lw5JiRqWpyoEkRF3BdGuI/DLIzDdd3oiTxdzs1b80L/Cmqhk61C37sAt
KIrDPUut8oTNaMuCvtqoSnOCA0PatuHZBR6A7Ja1gxe9TeUesSku4Z9bGdc26pLJ
b8WMggDhwYWmGw3x9deRB5UK0GH3oWnLytd6U5cXyAFRF7loztDUqhrFCcr2DEFF
aZFNGOFedNsLHTKGhbluRPbpn02Ryeqzz+Yn51iCa3W9g98KxSN+G2RFQNrS59mE
53OHGd1Jq6uhD1uURjBUMDQf3ZI7NJp0xK6rdpvO7ja9Ht8RLGxSImseRH2r8i+Y
2PbV78ajXcGfmpa3SdoAJxbDqXg4o9nTpdWh5wH6yEPusVjRWyTCBJq/7xvSNwEd
34nuJgsd5k2v7+9ydeNZVXZ5RI9o149JKdZehqH/y6Yn8raOV6ln0Mk1iHWH32ZE
JLLEPk6L4hkjLStdEQqj+YJ5+s9Tozni7aEyFIj+Kn2ImdQx0+p3FmeNxEb7R8Dn
c0ryFvA2NcyzjIeZaUZC2PyeGV9lmxg4yr1GSeELmgWK9N0Z20CDfX/whm51ON2M
azbXhlpfUqBoauETTL+dRqRAzN1UtRdWUBWvuZeVg5Z8Cecupdb+rNsnK4Z4XY+1
AbqlXnUnKbO19mjzDnm1XzvHxAFiBLkZ2sNhnGqIAHqiT5LFNICTN4N4mupLX6cK
Th1BkDNmD+bHfNsi10TVL5xllerSjhW5r0nPeDlGGlGiAZuhzjODew72n3qWIAB4
s7gJTTaOSJM+g6ys3eXr+s7QJoQDwzwZepMA2f9F+aN3kHmo1I6Ke72s9oloCNQ5
erOi6mVNsTCTFs3hYu0dUCrKQzGbsd72HzV0g59va0zDwmoNmf0DmiInsnADlRak
QMtJF0O5YHN0xacWjtP85zBSBVxhyhB5J3+FFSowp9wiBOe+RLjwuy4jDi5r/1qs
89Kw/O4gZCJraSwpXKa0z5iyjzW82u2rbNuD3vNUhAMZo1/DWOhE6F/0B72qL6lE
ze1GT1/scm6i+z13zPDByekQJIKkvos9yjsy+oauTr4nbmtR4rhYnAjZPNcNuR+0
7HDJa10iO6PMgF1ORRQXv5wiRHmKdBGOQ6XpI7SDqoaZhCv2cxVxKHscUjndF/dZ
7RzzBOg8PBocT978QC21ZWcSev/In+M5nqyLRt1SmggMdCPA3DCP6IgJIegFpugX
vVR8uAhfSQDlJtefA0W1CX2BAbS175hQfCCRZ0b7MFBLDMOxT71ndIftsb8Phd4T
3G6RBIehQCctebce/WOukpPiX8gNcFsA+aA+oyXrlgr+W9R5yt5AegJk9boNTmLJ
GCy0tcTuXmmyvOG4u/A3vSC1qzGDb1AOpwDdbin5nAmWUJmnTqUJf/obQ97iMPB7
djgHoJ3s3LpwcHdUCNSGjESyotjiXWCjwaPkSGrPPrK8ncDfaB+8DJU4OYpoXGYn
NSiZc1QvTAT1JY1nMTu9z9gDWAIZUv6TSnCp58PM5+L3GtlDDf+BlUgQo7b+oU7v
N/++mY7GM2q2JzivlxI8iOOBDsi2y2yTbow2xUXgZEkp/c2kdTHnn2LMoB3X8Uk4
adfmJp19ciYFhZlsS9IjRPZnUp1cjHCCAGG6VmxN7Zsu6vNgFp8yq0QvmdJTSvLX
znDKTMmHoWNJXtLRN4pAhm+QnWzTh9kpVt8OH3kfQFLW93ZAoQk1iUhmeuwHc+m+
CjGMgZhw5thPR8ZhriKPdkxPJMCDZFFpmo3a2Iycat8Y0kY5qvrfvrb0wUw750iL
rIG5u9BDTWhKqxF1kmXj9/ogjgBqUbou5VJP1X22UxZAePMIjAEu0SjuaBYwGMDb
GHy/ipLx11KbV0raAx/WoxCMMSCgMKZBVwFFmwKHm+t253NIZlTN7hyacFu8R33c
Dm1DnNipRekiOV9cV+wvwwpNk2jAbP6nCE8+J9ul+D0TnhIW6IUZKQLtCn5/vDS4
Q80L7cfnOKj8SIuuAjrsPTzmCMxsDTih09lrPp/vxk4hlM5KLWo6uTV4+Myr8TGD
9+PxbQw7pzkXOtSqvkFSX1tq0lmkpcO1/4fl5cBm8XFy7yCTsyuI77VQ1TAo5lpB
ZPoA9DbenCJXEdYtJQo/Wtsgal84DjFsx6UuvkneYC7Zv2dFU9tQrkriT+6qoIp1
xQr14fxoqZZRoL147vhP/fsr47I/XIjrMoLo6bNMV9EdtNlNpPVZy6EkXyux3dFO
UQhdTlg6pszMY0WsqK4IvJClz1AlddIbo5Ms8Kn/onTr1xE1uLNS9GDiBi2N8jhj
iWIhbk0MPiqBNN75rnY6v5CJ6djRQx7fstWPFplUdHNflGYkgI7vWS+GMXJC35m2
fQj3U+gsOluqYRUGaz8JTvL2cZIdMxnu/mCLxlFM1uWn80TwSw23Ie/eUdK33Zxm
1DRilGReehCL5p89/93tDLL2QIO6QrT3eNTNrr8iLFM1/qwGY4x+dumXfHQSEba+
vJv3SfILreY/el8n0RwIK+sPhY1qTTIkHdupXXC8cjTnP6bppeUlk2P3HxBWWwMe
+AOaKyBnAqWMtozwmekWZGBpZsBI5/Uc14qj3hlcijWKsn7rPf+t5HDFph6rPA/p
CXbpwuQAF2c2Z1+7YobRGjhGR52OLElGuIcJlFU+uJaBAT+dCsw4vx2gxZG60N5a
HLpa1f5EPOG9+/TOM1yapqDauCInfADhnlnyWcVIyEJNy8RRAxtLGXyDpe+XHx4R
kLJiulq/tK6W0jKv0jqb8V6eQSXdOmaS4gWpgi+/GYVpNQrJ+PqQEKECtmMvH/A0
WY2oLD++UL2qLkdHXEayyaj3ucaDE4qMdXmdreC2XJ6PArvJqtRSDtYkhFQyM7OC
QApWn8BCl8znGs8eO1FL6sf4pDBkI02UNqG+jgNNRtsLhbs8yfMGo1MdWMMoRWcv
F7Eel9w1cUofFlWsiuQK5XRF1rE/PXqJejkOhLG4Ce8sNTH1VQctbjlJj7ZxI+8G
IzN/Z7fJW/wrkA/sWYAXWYhG/3nYNcqgmxoLeCcwWGHB8vGEfZnG+p2nTKq5ypJc
U9/1uhKNxcA3WAYjaUnhIbQGM3BBDX6wP+7mvkwfutj+TvKvzalKK7nw7WGANRYI
4HillydE7CRVLxf2NlXIYFXgYFjgdRNN4YtDpKda9qfnBPnV5YzzDoV5BGVNbktF
R3vg+BQa0SWW/gWDvGocD27cIBfh7xpWwaOKZKsAzjw42BcGx97hZsKYh+TZuv0F
+RPLngAKA+RKYOQOubMvjVVfvnIWEnVFIJ7nJlXmDRWpG4GnxMOu/4+DRDvk0Lzx
nm5wT/I1Hc5edYmFwpqM/614gMDcyZFquaYh5ALJulpyPESy2gdUBJgpnGIDzH0C
/6448RtV2EC+fwa6hfv06N9FTqaPdYxhk03Sk6LOGJUSJFoZpQBKJzkv5eO5QFiz
Jg4hyPRN/VvBhhebCKxU6HjBDO2zv7UgAH9+Z1vXFWFlZ4hzioEVKbEADNIDHixB
sS1QcFnjkaP21W2NkahBJFO661fX02vB+slwFcCD/MtOGj7T/Xuqz2KtWei+98UD
rewJmNFmev3xcoJH3zhwN+FC4VWLQUWARuJeUaFlmlY9BdBWX3y44EF5mcI/BPW8
i7+Z5mVxv4Kdki0f+YvJPp7Zv1L//qLYW3r+UUKQyNi69PgADwkrZ2Dx479PXaFh
wEuLmmyMvnkxJQ4RtCGwjiELI7PZDVRLvJuMwcsPDD4Fk2ocMgqyqvthlUNkxrPP
OnwIxUHL5AqSGXepux1D2teHDf5P2nRo+GQ3HN/d/Qz60UUoTkmw8wYjLema0aU+
THNpzmyonTfh5B9e/PV1U6+N88ORAqsDXBYTWei2z5iAuUTs0iey6RjYnAx9QkGW
6Ly0xTt0xWepD4sH1Rkuf8Bq669sqo3DgTyQuHp8MvxnW6qx2mlDmcUJkAplMjLv
15D8T3ehZvkXW/jGjraFhMB34g3ys6Ed7uaHUS06E3qyQ4pAe3lPRa4hFpEmcM4T
pxQM8ppDrbcIn7Ir9/0DCtlNY3cKChGEeMmHYhB1PoR8UZxxnZvTTKI5kB4eoyFs
l8MAwtrIVe5RC6henRCkemnhZQFa1QJDfz8WKAJTQ/mQBgb5hm/0Ygg5yWuowgmp
nMqqTrJdADrfXpPNQmBHFEsye9BARiB92bF3uVsUAv4WOP7Z7cAx4/4MnVEGUsle
adIYoi48L6HdRz3QqrwxgzflsTOGujxYGsKXo/EvU2zKcyMNURiMZZ2MUUbexjhV
BSypV/FO+gQdaZxT4bRFVt4otDtmiwr7smlqfzX3XgeUsLPzy6VAqu4JukhtdLBG
JPg7CsDBSZD0GN0hgo/BmAIw+XFtMLUpX2wHbX3xgOxGAcAfXvPMPav/d/jhhHHg
YU8eG7OZRiObZHQpuZ82lgAoluY/bf5wmJl7m+mOkAVZssJ6HhBJ57U1Pt4gu846
5etWXMTAAsrx4dERobKd5peJUjOZlo2Yo45iLDcNbPWzP40rKNibqqm3K/Qj+7wj
+hkCCCkj+hDm8tmdXALtLZLIjUb6m3OHbuUBmxNVOLYugoZmlQkMY+aqdhKFH1rl
F4jDggJjYDlF8FGfac88lSw3OUR74QBL/jS/CPKSS+xbv+aSASGc2LXyLBVI4W+c
aIW69DIYqv7WbGoHghqf5L6CPPETUeSvZ75NXgRveAkVBDtoqCM0JUk1xYahxIhT
mccWqYNXhdIDSF1gu2rcEu0HAlj7I9XDyEHP4oeGK1Na8fVY/ucK7vplcrl9TtXT
eDQVMC5Bybc6nlIyzZvH638Eo7tQ7uwryN3M0JThmeNkrukjewdK0KxeA2741l9i
slirLcOINPqsaiDM2vtMmJJoFdAU/PcXEPy7WMXH6jf1YxLBew1ll+Z38CCtPAv2
l5eXbcKYyYo3WlDP/rkccV2K2UgT0/YkgelBi4Q98GrJl/TIq/S4xOXlFSXqu6YH
Ta4dKYrio0VC5ke9yr0FmJPw6m8T1wvKTmiokWihdXLbDimLsTmDtAT9rV5/deuT
fdhQxZ84Pi5STaUD3ke8D7uRFYqpru9UfwR+pqjn7jVO1rg/VED4QPQdgDKilgkf
kBoWQ+BTvokeRuFh9u2YACBzPQEwvBJ8oGkjY2h4qmFVdkcIWc/eoBgMmkhee46V
ln3zdXxI3ZimmOUEzmUX3hulDq6IWehB26fa3HqM3Co1URaqE9J65Ffs4T8lAmx/
N1UbKHoC+X0xI+YKswDqPqDdAn0AnW3Y7skvk1+jiFR9xIvUSduUMsy0kkcxrNOU
2OtzQFp8s3/O5rJsj70fxY+WmiSgpq1ddbthgbjIRcnfpeOGkkYiU5eCPfgPFp2W
Hj/+CMhL0Uz6sTUxfKQ5aeJPTzqNpjMXUHC712gu9DMOUiXwy7tTEwgRcVPTEKMl
x0lcdPXL6cGmyYtyMbT6LOYVk/dNjd1Y6RiyF/kHsbybHXEHGum6CqCTaKk0Nd+d
C95xNejPZCW7YzKCm9stERnK/jzuVxpNjDkmFF0SG14tl06iYSnoNRgjzZKJNQgk
nC4zPUnAyHVl0oMyVcWZXyyAt03/oPxbTqTy4qNovIt416snBIwUuqm+UMj5QHvs
SthgjJr73VL0PpBWcsVxG8Z1Kzh0vq33a0CLVNw4wO/bWSXGna7tNxr5tVGiuNG5
vhqoAGEyjiGDowBNss5Jr1BGPYOeAR+5IlHLde7onNq+IhOgxXpr9pax1w4nz+Wo
k1d8oGSwB2wLKjTT6TSQ+FnG3Xtxeum/0ZslZPLZdH66OEGRXD9KdNFPE+Y7u0pv
lxCnbCynhKW4eB1YbZiMfqkXhUpKYZBBWfFyaRGl+ONGTmCAiBOYK9EGfwRnQdM6
Du1rtBVsQ58Bw7XJOpVml86yfOLBooFhx8PreNPBdHD+Czxf4+JSrtX3ajU9++PX
vMtSRi8NW6ci3oM6VxNDjnAX/0ujDXwlwgsXku4puYDabAx5XphFpV0MECRIzZHQ
aBtI+eTqBhgyuYNe1lcScBE0ABY0rZRhpIVXERhxyCsDza8XzwzAcjFPA4D5BSiy
OWfwbI5MR7Z2teQG60fGEOAV5cFoGhsQmo5F43OMXJ/YjnXta2RzqqwbZCQML7Au
dry4ANys0Mre/aEyqPLpht7na5Wq7UVMvrhSDmHp4bNNwaMqELRzlTRJjAg33Azm
73sQe5ir5G1xcen44OIVS/NbhLB8VHBclUHIDJHW6yG59qTaWAyRJtM+tiJ3Zgfr
e9tnRgR/vhiC4XRQ/omLL79iWuPXoMPTXuyF3RUiNT1aMx+jv/YuLh1biwZ89KBX
uy22e4vKpw9ISh097P9Het2VYPDoZ5im5m/zv9fyJj+2ZeCZizdWa2XDDQQK6jno
6MFK/usz/y2smloA4YxreDAYCwy3SbaUjpGvsz7rC2+p6lrvm2s+L1SPn4q/bfez
RT2C8n6c2u2iyIZNBGrk3iD2TjooTh5jXXEcXuKaD3bEpnmlt9mY+AzncMSoLTcs
nq3O6rxveBjYDM2vrbpZeeTc2P0q7hNcEKGlEgoILIhYei5jwm3QN5ijQkYL5CAm
UuhtuOym/4vrrUqUaKwFDRQIkcP/Q9p0UAMqOmAhZyCluRbOszbcfPbv8TsGmEps
iyXjwl/gDNacrSGJ++RwSbxjjWxskzCPLWWKrlWtGw8KF7kyAWy9hEq+yhNMcisU
k2zd3EtCzT5+VRm0GS/XC0VCdRZnAYEw1M3oMHcB/qoqi698iSiEAHVQpC/x7ZOG
NBc1/cTuyEgVRY6WeZphXl1M4q5DD/Z4H4NH0zohrt8uo9Lz6sKJ7t+Hr9iVR6SL
sn+pIXmqlu6TLLSW1z+E9+lomgQxDka+NYYo2WB0nz9IVg5YwFlH4NwGZT27u06X
rD/Fj1d1jbQE3K061pePHj1QGi5u2dB5qabu+1r8OaWyNzorLIsU0Uoy2E5YC7C9
F8kEZUQJZjPsuN9KeLKH0SvCfR3mXVbafHWC3e6fC2Z/Hm/I3YcsEYjh3sjYrX+u
7PYJOLJRAk9lPMaWgRWUDm6o7iL/0NCeSEW0aiU1NkL8SK03iUySobj/4DSk0qq6
UFMpNcNN9CdaAWZyJj5IKzK0Jgz5IOBc3zy/NuNkWjqYt2HMre9MyNnwpT6+EUdv
pItR4HGsHJO6Dn30hvZhXVcfgIXP3uoVoMnBdbog1RDw8i8DoTRY/xqQ5qP8Gxt0
yoNSPIhhVpcUkRCSiVu6kCCUG9V8oOP1Irlm+dA8bgYMxA1IrMEy7WCJZoM4FLMg
h3cp/27BgcZ717ihvP+dEpFcHJV3SwCMSXbN4hdjhqpLNgIj81juTG4ss3A47ezE
gjotf2sWS4bzMsgdd7F3pd9xXztiIEFsAETscBCtsDD7G9BeNOaGwRoJP+L/636L
4B5eNJ2kqnkEfIynoDMZDttGsxUmSZuwm8zSI7tNrzLKn/xyEf1TqG1sKy15MPUi
2z2FZmj+MCdrPhX4Hz0R5JBJbDjJXQhMoULqd4cZYqSv603viWDRNHjgfSElEZdR
nSAqGq1J+13kqoQsuwzuRkI9MG47G24MuHhbxStDG7grOq51Vcj5ikc7N0sM2Zhg
EothJawaX8Zj8v6VoKBuH5hYjKQ3JMDexSnNn67+T1THx4Eu2pv+GTNx2hdCFpmE
B7BKT6QhGYsRXeqVhO7qrRbYHVL8slZk1HSD7nExPeBiwGtEsbsSVz3/yNGSPvw/
K/ZS0CKjUPUb6ZfySRb/Cb7lHojWaO2OZpdoyAeTZ24CrmvsNOzQfBE8/7XKQU2Q
2aVIEwiOyQCX6H5IgoNX9ybw6UyRz2W38N6lYLqoSWpvnUP9sr70lRg9lzlLU6Oe
Ytr/ZLFY/l1Ljr6QIq3hK4Qc58GjYDDVn7USzzX4R8CKkWFknjrwrfaIQ2HOtAsi
qrMjDXU6njkC9uruPbLwNYxiOAQrjlO6Vp2+6IQvDIfEH6WCI0sjgCQv0SXMxvj4
ewBlgqyUO6rSDcIGfqg+ubCG4fc4rlPTbyYfvN17cW9MGIehnZCtCV6122tX/+Rp
KARbvQ/KPiLiTnx3KLJI9vk8rq4UqHhGrhy2URFGMiMpYY6E+jwyT4y4MyHGVzTQ
2vtN7cfNI4heppHnPiXYjdOnyYMssqR3oD/7miyeBi5TLaUVicouh7XWUzLNETkT
ssrb3ul3ABwHuMZtd3LA4LLKe5JCnvCDiIz0uGZxtsPWzNe+TzZvlMJlZL28L8N0
hytTXNpx3tCq2JYuJ51DfkGVQBArorUYdyiEOb2u81zCyhwqvET0HkQmIiVxc3Ng
m8DFaE0XUKP5xabVKoCHzFVl00xLo6nZ1h8luWPjOw52dT7UjHQ3871Y1JA+0iVo
c2liHCSrLFbPPh2PSHZFp6A894AhCRkPyNgt/Joj+YCxLuBkGerBhtJy5j1F004v
9O6dKZ4yAxDKOt/M1gejpkAf0Kol/pjcnx4L/JypUB2QH9Ego+J4LBqB6jDddTLG
bHe86ZI1/fvxUj36oyssnEtcR+O6UCspKpO3aP5PqQD6Rq0jULGMWQf1yIBHantn
DDVbX+oBaxPP/7Fe6MSEEw107BJiQaHSKEvHrXWG4jbD4rUAb2kkc9xZLcU8Y8tO
Imjp7AOgRne3lCqb4apJ0lezwBDloQdYHcVBsmWV01lxOehpnSxpht4KeYZL6aVT
mRE9tHBVdF7MpNt+xZ4Z86ruj81o78H+YRrk0aUCrToUCm2ha+VIDeEthrsWoIBp
dq41S545tXAxplTvOB/++4766BLkVq57LdtMP1nds9MhGHQo+TQhzTck71jxPDMh
nDRAkV2h/FSCIMZWxKBFykOa71T9oGqNE/lND1O6UkQjSqGcBHwWKenAPGIjS9RM
C60hTC//FNUxOqcuJVrJO8Cn/uZrCi9IvqPmuasii4an0a2/Yp5+TqCk0UpSR1DT
IzO4/s40tEB6/SyFPcjj/ThM1owxk72nPAZcCZpl2hJcDPoPV8mF66FuZp1pz2CF
QIUCBk7RPIJzL7tAdD2jpwl5u85M2TmG39Dl9ZwZyH+Tp3DwOCRuwp8mtgOQK49x
8wYXs0V3WuWeblQjhI3aYeJI+glMQ1oSYxUSF2FVVukXp5lJFyh3/u6v9KuQSsIu
CtwBC/l5QV9o9Di0KJS2btu5KzKpW7s/CaYTeKFu2SIQETTVLcn1f1d/EWmuW+fB
1z8FJLQbNNVoAbfCCpjVN8NfwG+XNBnCwbaxE44B30KirgwNhCnxY1/Ep8n1ZH8n
5d7H3Xm5TpT0S9xd4tgIKLBcnAN6GGpQnn6FpZFKP0AVSWsDwmCQff7X26D+kfP7
eHqBCxQilbC+87aRn+VcFK4/w3FqXFeoCAQiyukBjOiJhbw6Ucg78bhMcLND0FcE
4iRwt2ZCqMnMC0hk1WbbQodDGfC3CLTjyueccEeq/L7n+C/eOUXxcICjEUFCDsh6
5CKonpnnLowVLtSe2AlgVf5d4lwIlO76wVZFy/W5xmmQZCX8eYItKhfI3jiP1RAV
Ml6WlWElJJM2WuYkfhVFqHHy/HAT9VF/+gDZx22CGjh/H2ApQzbH4z1E0QUHsupL
e+PtYwzvLCGXD+PhEK5t/g4DjXjMTt+rP1Lfzkf8ZA5zK3ORkzc4MEnqM4SJNvGv
x62ogzmt5VKQKhXK2WH5hmCnztR0qqq1uoA6jUiyQj+Gmt7+GQLr1FV4cB9pmiND
hC9XxfV0+mwMwjoLWHmJTGKoTzqiVtD8osCG9iyszUmO4enBHDtnARmvd51SjorX
QcVffq8L6ZE9RnLJOQjQfn8sf248OROdIIy4viNxwdWtOd5aoT4Gp8qd48u8wACK
aP3NlZPy76qvuDJytK3nTsUDMavMTMrQiAU1MtA26wGH5ENHM9wzSBSOcZhPNSaJ
ybJAkVFWMKACnJCIvxCnEjGEgut3lIf1bR2hG3kmimIPlJ6A/t1OC+/mjYK46NXm
QGA45uCOjGPTyeZ6RDWTmpFqJYOHnsTh3luk6+gO29YWIaPyG2heeUH7/TrG2jS5
fpP9b0MQ6l5ZbwdssoxPi5Wne81Vsuni1jd8PF4xMJu9QsGFPijZLNWAeM611/rz
xVkr3/JN83KcjzBsae+5dbNz5jBOfMgDtrrLlDOap9g0rI0i7D6B+eDXh6lSeJ+w
5om19mJGvSW1D8HD2kZZ0rLWSBXdcOGuYzeFs2q5sg9eR6Ejy3B66IxitNx3lbcg
ijOUeJCOwCPCH2zwoVTgI228B8CErLPgak2s/I9K4MGaAWMSA/zovET6LzGfNpGn
fgo9cPgu/VHI5fZ5VyC6Fu5+MnlBdljqirhsRTNMwjClfwlMJnO5gU8riqhop3kH
56sFZZeQ7vjJRJzALvl4vc6/zTTomtZiZB3fFdiGuNKFgBJAZZ4/v+1Gi2gzEtUV
OGm+azkj7rUn9Fr4N1418oUX5wMESZufJDP3H4UpXi3/iXJ03pP4JZOo4vVOLiEB
b0g5nE4dS6pCu2ZUnjIkPv/YG/Ke7++dsJRdXkk6UEDWoxWp60GSt4fhth+hAtcL
Gfn1GXY2ONqz+DOe9gOGgChxhjvMOV1nKbbyvzhWq/viq7fto/P/HDBTSQPj1Mss
kTTcQqiZnvyNBwQeU1CSk/dX3Wd4lS2sRUAo5sivNNb7uYiPy2DqY6206usooR5I
ZGUhYfTiNrPsbHejWQQMv/m7/YDsqBxUmBS+7TL/kFqolXDmYcn4tOF8EUVNzCwu
nbZbSvDJbbH/Wlrmdwdybpbifnxi+5d3mBIJ6Hkibu9lNu9aTfmF1ndKo3RyYBBt
fTLRxkHU5tGfjBb1THgDxqGJtjKpkgSidzaqmwvstJbvQ7qt6Rpdmv5rwuMnNxT0
jbAT5jEKcOJBSuOSl43qdkP7ruzdmg5sxEbJE3JOSA7xh41cK9vIII3LdPEEbkVn
cNHrx0kA2674yAcba1QRJCEpdtnlpJFjkmotKQUDBVFEaEdmn6Y710+dJEpXdKbY
XbM8L8JV/2CknBrU48dEqmFJ27te9aseR+70ZVJhKefsw/1sW8QA51WRU+EEWhho
fL9zmYzstY8GoUptethKq1j2OXMQtQ7Qe3/o/jmumEko7WwwloxDI9z6hYLkbIQD
Y/bbvLev1MQHZkhWNdnwWcPOrPtfNq7nNsrLJ6QmYJhHtomDTWHvLaNU8rxMR/Xo
3QDRAG52Wbv/7n8ngZ3JQg2Vto5nYtXAGLqjgBd3J2+INKDcnLvO/9yRD5vgAQ3Z
WbGZbkJSLhz+30fYberPWD5KY6/MMbv5PKpKDXSz7PB4kkkAURjIpkFkh7fgMfJL
tOEw4E0MzJ/mP6h8r2eGRlQz44vmr9D/xI01eoWl0RXmf5oyDRTo5zW3r484a/TG
jyCJUz2Xf1UPcHBIbXa4xDLGXF1An0MVsqnyg7qkZzw0ZsdBZPQrPbwioiW5Gr/G
zTqZbuVClMfu6s9DqVbwRd9WjQoZrasfxuD6ffwgsr/OwqUdYiK11kdw8XPizVDU
HxHFzDB9oUOaKyueiFqRu/LG7nj6DdwlSmbGaq8kOQyN211qAlGMU5FidBVA3DB4
lHleMSwHRRbwkhQMcK4TZ+IDR5o3LNPc7k9tC04xVHj2BgYND9H8uBTC41TMh6qN
sOJfSCu5PyB8tgdsrVm1gHkNB14uLLPE7V9lP9/YEQgMRkaRixmyFs8kgN4VGaj7
OxyxkYa3N/o2ZLVHKbJkLq5BmmMXB1fsVH053pBY4zpKvYZfpV+K2iKscd+nrT59
3eSwva09HxU1Yuv1o93FG1kNwT+roVLIjEckhtwKWPHTvnNDUUbT6SIeCTowaEDZ
bhJfIYi53Q7UYvTeSvQ66YjT38dHhTgonf+garGE3fjp/EkjNsQEDb3VTP4DUUX2
nwjU5H0+aQdESWzHBCcTfrcYTb6Ogqe66R6amMJ3MieeRqN/bF7UiX5dO5c60QVI
+qizC/kRgoZj67iA+e57Raqs6174gukR/ZwEDYjcUruPRGZQGpyPfNEonuWDkWh7
0zfd8PZ1iZqQeTHcGef94mXKmZf2leITYzhhqb+aurVY+9ApElOaJ73vDIwGb7cI
ee0PJriaF1B/m/EVKJsrFyck9fAeXPrwrbJktR17Xiz7CyU0f1TgmFcbX59/i2An
msBSYOWMZ+BHcr/+39WJo/OYVq+YvARirOYq4mI4klwdR5HJzcI2WdlJwzHWmQqt
3PjCMOJlCwzRkJV/uipF8vm3Vy80V50hEO4aJrLr9N4azg1+gdbVbeekTwmUtzAR
CoEYDkf13RbhdxNzGMp8a9gqshBSVtFfg5DvK5DDNXWtlvJMUKE7cnIrbhwmAglw
r1evAZ7TPVsJ1oxw6BNr+J73LpIMIm2JV6yR/mIJHHzQaJdXUVCveHxlPLoPq6Ku
kJMMi8EVbiCNpWdvueQBss4bTUoJKlFqoPbpSRp8UOEDpY/54kgFQwZaGWMX0w9V
CmV3sGsIOGlcvOGeM35Zn5Q6wv6cdwS/UWmOWglN+TVA7l+S7CHH1gqSmsica70/
lHTQvxXmFyD5ye4N4+i7+keqlthc+otoSchWQH8koWlkmf5UkziXlae/S1bWxw/r
1b94ZHyN+3xKcLGwLWKHOj40vN0CEHZOFSh9gjHfkQM76a5mbrAGzAQS8QCF/Tm4
QlvTyoJFFX5hFSvkli+NHW1bEXUlMXF7GIbES+e1gTGNcwue1pzWBqHb0B2ox8YG
m6UcJCyxEAnvzKDEm1jC+mrTK/8k2H8n7QhSKnUQt/NVtKiD+WNa1R0Sj5F4Tge0
uwHphiWn4UsTAl0mk/+tHUqU7sXExNaHv+ODICaPB2kF1ed1N6P6+eX6pI01AsuY
IofAefePYD10rhLaKeZahmytFm9zCeePeShUJTNMnHS8jPQ+CPxC8SuwqVUaJJBh
gpcnKL0q2LgM918r375v+Ud/f3T/ZdJte9q/6+HRh1LhqftPQx4UwtEhAsfEPXgo
wBtUA/2c8jkqIB9y1mavjPQsfpGr6afYlE5YNLNhzVBA2e/drCnJPavOBnlNWYxn
nFChZgf0W/D0OD6x8tjeGuVMXDmzQhQ5eMf+WsDwbCr6Ikv08dD0jzg9ziWPsVZR
fE41waaqDqVH/J1QxN7s+hOKSBcQ5RXoaBOFDTSOD+GYATeV0x4FWmuu8x9ZA+1V
aXnt7R+Dbx5Z0maguQbk3ycOHcbyaITdSy57UWHgt5dMEreEMXhyvsp7zZYUmuzJ
zL95NfigqOsYATOVx23LYACn+QSfhNExw1GAZ4VtCo6osS1qKUVExhv1lqDQpNSS
rJLx+eNkvEC6RBiyJCrDgAciMfk3GkcEu9P3MkEAVgYx8sKkMvcMzYX+Sx6xyaSB
27UnQQyxiXNI1C4NIabLa22BpSyq6VqsGeXitC5HS2v9AsETBnbOdp+nQhwPWVkO
Ex2pHTMcgfeGwwUBur09L5S/sKifhOkrd5f0Fr31meU0L4XHN8FxbH2286HZIzX0
V6UEfCWyNqrPIKrpEaPxehx7Td5bNZyjWUkd7JR4s3XamoubCOI1eOm+A/8pLwM0
3Wu47x+mbS7dq59otY9tdONduCFDDy/uwpuymNao7QxMQh14QFxYtfDciNCDX3IR
Uz65nj7HR1fwbsjBO/a7EA8ewFotRmSaerkJRIVWbPDO2rGUhXHTk64do0oxb9o0
IErM+Z2oDffhNhtPZI+LLriLcxD/0jqhIkS4zu9gFjtuZHRIMeeu/caAd3zYMOAl
yGNuBqeuzBAcbNvCFQkdxqFiFf07ajvm8m79SbgeSy4Pk11Pw9GET5QwjW9LAjN/
szDCs9XPCUngeQ/bKulOpdyrRt6Dnj95lP5biObQus21j5T2SL5aIG2Ax5+B3hJh
tkshEzTa+kNJPMb30QKPSSZ/ZmF1oQu1vLsZhgTUafHrGqyUxIv9e/u41/SK6YL9
YUxk0gH3a9OnV5K7jD2+ff/t077vifVD0FygDPNPU+6tPrjwNewkk7XICYFbc3AL
Q4zkHG2oNgTKB+Kf4JRXpF1rIyW3FNGvWHzVYJSmfziOZGbFEkxUK9sTXmuX+mSY
O8iSvFhMbcQASmn9wuyjzalDB2o2NCKqKUXGbt0EUq8myC9oG9kJImJKM7t1jWZe
AMX9WgdbhUdd6YlbaiCshdSJW4tl2TKxh1KSlQt/d9+NwksgifJnoxFLJdwxzz7w
d59gz3c/Fmq/cVifzgb05Vo3p8r+H5TonxauRib/Q3XXaD7ZjcsqCsNrm3Ykfbxg
s95wOgVxbxJmQ1GUMJaoQZIdvE9hTiiNgrd0wS20KiC3SvvIJGl14v3W/k/C2Dpt
BMdZKjU83yms5f09zrY3T6bGtGZZnKv9KiWNG9kasi0ZO22fOix3wzcMe6/umWPM
wJkvWdz6/qjTKNiJ5oxV+jKg9xIAhieuHqUENuvO5MY43gUGuqZGhDskUUi96T16
AqDYpagBgPsm1zhQKlegcl7K4grn1sbK6BZpWejS48ulkamURnDlb4a0uZU9+aQB
WdCYLLAliB12zJYSvJOX8ytcCWSW3Bw/4spZQHlrL3Kkpza5sKJB9Q+R/GYdwB3g
YygAfXI22Br1ZgISCRhfG9M4xMZij2LMvBcf8CuLIxq3wjKJJvlJNLV2qzO4LQsc
elJki7Rv+8WIPJ9ZQV2Om0nVuQQL+CVibAhw5GxmzdvF12rgp3ZgeEaUXVZOQWrX
rOXSTS+//q0DPUnXJmx9A346IKLiImKiUcVLRhdsTlfAZUFzIGKR+KKCLErScEe9
KKG6pbaxMq/y063lOkKQIJ5ENbNj98l2BcTS/CJTcCIDeHN2R+qISySXbrcPNYjG
R4mN+yX1fFEOFuzWgd79n+QXbEGCh9Iyr3WqnNXLIHrEU7y628jNBz30rFaFwYZA
CofW7Ug2DkvfMW7/XSD8SlS/5pLL2v0PaFVrskyT+btwld4O4jetjIPOUn+3IiXb
Zgi43RUtzuq0tOMbQ52sh0WRb0WiYeVBGVwLQeW1Tsau7GokPVs2MQiJbhuFx7vC
NVZ4w1JD4IEtvCwPsmAeV2IZjlYdgPocYtAVl6q5d1JCUZ8jjyNSufHZpj+ViKXt
rYCAlTBPiwFeg7nItymuPoGHGjp7NTvtr02WN01cnR/ZtzuqZldBwtTs98h9HGhE
7xJdkmS4BESbcw/evaU60tTv1EznsQaMPWHK35QZORqJ5kSIytUc1KcrVYc8V+QW
BEyA2Ja7mgOUxOHSLf+3FnU002Y1+CkredWuILsAjzFAsKdzKaGW95EW9RlAJ5iT
9YZtzNErBgFKWhK9U9Sf5VBV7sd/qPHLdXIeKNkp6cz5n1cwDRActObZgMRletoa
uJNelGWG08brxH3DNpoGuRojULH/34fylD+RSTg51GMtsldC6OTZC+H7nuSTeulO
T0wJp5C0PH0mcJtClA6CftekzfjcW4d6VidLMSWkfmSK3sPjXkj5134YmE83dkvk
kQRh4MixKY0mwbmwu5e30A6N0Lt34p3uA7I2MNv2/rIWG+fk8nshm8fAhU98p9uc
lpPDGWBYrm/vx3AutEbN5zhe00hwX4H4ob1mqJbkOVF9t8kfrTa46AgmUyzVWiyz
N/apKnW9tcqlfGAYMmz9ROv3qx3NHoJPIqBNtrdkwLJzWV9A7bK4LBpJwj+G7dF+
bESXwQsocJ855mduDbsCUNNI13pmjYuKVB9eEwbyijVWe4+i21T2NK9PlY7hVoSt
uY2wsNu+nL8BRsJm4drHj69oLcj4HVbZ4tvZdkd3BUodpzu8J8tyAH+oqIp26kko
LuY8wS5azwMOpM5NVwxlNkSRjO3XdqOJ3KySfOKvxUcXHtPZCqSwTdUE30N/SEyT
iIcJysyhcDC94h2ytcI9jTo5gxq47iazXP9j+0wmfjezuZjA9EZ9z5/pmYsEI0Hv
07vT5vwSrfQwrmQ2n6lRDOTJFQHrelOwUUXVmpJJDuQtWDxP3RNjxzaPuQQInL49
RPbmDBx0sWT9ZI2S69bulrx+AvodrPljAjBaaGBA3LojCR5OqxWDI7SwVGB3Sigf
s8cDeEfEF44QDunPADnbv407XpQemOptkyWJ944onxxR4f7gKQi+x2CjOB8xEihg
Qo1Y7Xd9xp80kSCvCrvRG6K9gf7DpPlaG/NWBmsIYXmt9Glfo71yIuFNUW4245y8
m979MVKL20ui7TYIEHsMMt8ioybya2X3g1YHEU6FmnIxnmHbOxrmzvWKtFyWN1+T
8lb+TGKgJhri/zpEHyF2jCkq06xIG6w7lMN5jlCQSJZHpNMNgdcHf0tu2EHXTg23
zvNRBmSwSHdnDesAZ5fKQMiaPQxlNwTlr0bVZbkobyr/aE3OjqTzWeOYOd8xc7vl
0xC8tfeSTiQQImwTHIhYT25lVYDK7tDFao2f0OSz2qDeIh4Wq0y6H5cbCjqh1fyh
+3IxJlWRQ67RCRahu7fVcIIYZbe2CTmI4my2QjSaHZIWAuJWEzvmBvpSV5Bfscyg
41wSRxTKhzO6SnP0DdpzSqJFh5MpxN8dKPbUxHuTmCdvbLoniEo6HwJFscrJwn0G
01n+sScPhVIT83cOcFrYaaDFyM4QeuADJ8BpYuEn4UCswYSoDJnTDdr8vPiw7Yzk
InRKjsG1yJeBGG3D857dx9YHz2iz6z1rOHdj077ekMrAbUHUyQE7AIXB9oUvP1Jl
ikZrSlIZJTg082pkHIutBZOxpx4RieoL6JzV1yomzw/nvA4fTTHSxOluLNBHgUE0
Uy7ZZqACTOSi3u57euK68L5iZiPRxTxZHjELrKouImmtLHv+hOxBtGYriHEqLIds
03YAasnMWTO6/RnugIFglyuqyGik7ddC4bvv3KgWZuUeWYF4FtFiovQ4E4QFUvan
j+/mrwmCLvi5T7i6CXT3HmYVt2PN8+8XyWIiObWMsSJnY0y2gwQ9cB80uAYdpaEX
FnwTuHenOQPsX3XXEZSUzXH64+3P+iBXyTOoDkUIlymPDieIErUtlPx7xkXknFXF
djXI/0cBT7/2eUWZ2/cwkbGIZAnexPUqZnIY+qY1qqq09kM7B1uURRrmnuSWfuRN
c0jMk0dixXM3p77k0vwZHe5XLt3r4+Elx1DffodgMbfHZwit7wC4tzjzDJFVqfNV
CsEvSDahjIle6LIBLyLFvmDl5ZLlVtHJYq+KNLiuHYNfo8egoWBRhifXZUZnQRDu
h1W8LrqjTnRbKnf4wu6ldq9p2GkJ3G2cANRqGsQRd4HN6vuiuRDTG581Pk6iq3Jl
O+LDtRh2lR4bEtTv3WMYBzIWjo7ayZlkkAoCiYZgSwmffGUd1VC+fIlcPw2Lkksh
8SpY4IwsAuIviKjcRRWEWbmd3mDoNegE+FOmVd85ePXbXkHDqsut+ow+G6JTT59j
4wv3s50xcAAsgIiEXVyOXeupwr9yZ0JqNBqOtdILcDwcmWUiDzYuoP4ktQUkGf2q
g6ifsOCOzcSYXw1inNnpn7sNBmPYdyP6YxysoNC8/73p8MIpwpkNwgZUDgEUu4e4
Id4wzWBzZG4V19R8OcMFpM9qcBBXF9Pi6PE8UZR3BIVVFUsDnuCumUfpY9CSpCSN
9lyyrd9LzN6GBQS0mQ7zQFrQ4WpwjbspW2UwFvsPT25iQjZ6QIKiEHq9qqPmECki
L4ijnrLJBvEdKfrey6TX2MoVIgxaDUvmQ+aiCvZeLt8Cw+l/uPAoWV6Mh8qrSZly
Gk5huvZopsz9VkRIh92MnYSVZd09csRYHjDu+tkento8WhXgi1rcQM8KA4fkR8Cb
KURGG0Xqx/htCOyK0piy11r/b0AJ2M7BjreDCtBSKCLQEYffZGxSWfomwPbwXV7L
Omn0jDP8y3DxbPy/F1fc/8e2+DXaSZabaGN2azC/tfk5xCaLdys4xIO75OuGZvmT
dRJqQKksevPOIUIbwisHgsfefbAXCPEfr/ueGJNfQG0sCguokGncrWPqO/N0el/z
+bDLWe0t2+3LvkiFqLYsCtFDtMv/EoytqWjQ8GsEZlUNIuQJQw160+YDnYRKs7ht
AHecqRc50eS0z/RQpVzECLu2NmIQ19nTIlv3pXd+9yufhysbmszazRo5bCoXvGW5
1iHD6N/awVSV8bbNIDYF8VTncwF5eXzcf5dYZvY9qCHEMNzojmzJBb6NXyEz180b
tReWBtB+0YuYIINYapyJCf2rmM1Av5KmXpD+Jeqg3SkqyBNpd60BNI0H8/CNy5YW
DL6yHIGWiSrz6kfAOU7wT8tpa8uo4gVLjBIAbe49CY2RsxiL6DJVssWIizP8kJDi
WToWuxuJY6LwL+7ywjk+F3u9Day5Y+qSIH0PbyiqNVx7pZsY1dn4dcSLiWstJ2fv
JkRcYgegLFzahfb1lo5UaZZo9ITQtzKIjYwLkdtN9In44al/5DLx5HVCr2Fla9/R
8MtfiPTfD97r6BGeyA8qU14YYmy+3ykDx1gLdANtVpvsxya0KwSX868AqWGgW31n
bcglzDXmBZNkDG/0Q7nhjjUpbRbs9tvoDtWBBzL7+OeVXKr5sCFpaZ5yDdePMqGL
6v8SMPe53CK7eIVeCdPqrKDWm+Yz5u0f3cj7USuYo81HwYyHWbT6v7Jh7VPGgJzM
UTT5J/rXhPyxkSxWD/Vr/1Qi0Shvz/VOwh6CFAKk5LU9B9sL9nnF30amthnCdtp7
bdcGPzb4ZDp3E7BjZjgBRF0VAiQbq1t5IC2L2qEUYcQ6fPkLGuaI70tYohhf0DfR
nAz9JrDPHplCdPKdUNX5XpSO3BKOMuULW05LidHzeVD9cd457Idt2w84HZAvyIP0
+q/vJbJxZUDgyhKCdajddF1Zij6/rM4Mog6ZQkFt+Xie6C3hbnlD308yw6NLxg4E
ETWwvPyiReo7RoQ1TI1I8IkGJyu3nteA6RypL1oZGr9j5RmmhSSSRQyghDiUtsls
mo3TH6D7p/z1H3IPNtkoB2dcjVLDcPXDkh+W7PzcnzVYNKbVdllrzvR4a9qepHT8
SDIuwMZx5vy5nY8Wt1sMJpmvbAzHzTctqRMp5gNi0RIT8hsMRPB9lA5XuxA+ZcbO
cWD5d108fWh9pcG2BBskFGC+kzLYIokfXGVh6Q4syLBJzaXXcR+GHHNSrkROFs8O
F5TGWbZqRfG4QuuiCJyAiR9E9x8jXBBzoa4HWMW5M7fgM0+IB7ALjh24FdfLsgIN
F2D7QrXMuX/FrmqoPJGdpFE0axY9SfjbGngxVe4ya4Ff9ITp1yRjPSGea/Hhn3w+
RvnM9SeNVE99DUVFJTnyUOS3WLpy2TZ/z4GTbT7xpXfOiIv4XG8SWkKIRoL5ARuh
TE7J9UwnMp5dL+GsUk+ghGQ6/tMLz/5l6W+WVnV/2kmNqG7aV98D7X1Lo8dIpBQF
MdpGKERAf/aOdcN6wQmDOrKMo4soM6RQQJ64QLruPs7t3h7v43PmkFeX6SEQ6XEp
Y/2CfMuKbM4VTetC1QjQjKipNl7vk67QOfVV0EDZ6MGCpcsw6MOi1CGAkJiq3tPa
d13Mpk/KofQt3ReDsEl4R6ehQgktQCdVWqaJebD8hSyGN6MkFwUvUxUh6+YfMkma
iWtHtv3DSPp6VNF4vu2DpWGuld6ks9iA69bGZdicCyUL2sbfI/8jY5ZRbQWkofBG
9zprVBJh3AWI6/rgdaTTc5oPIImec+XjVBa9gecI6LmRcYMz33zkXIlc15NAluLj
Gty0JGdfSxeZLaOTRypoZG1jgx8eFeRfskanCGAECp1UcrrCLav1Yookc+KG0p8+
WxccTpTUGRVCg/gSQLgAZsyI10jwfMc0Q7kcu2HtLHpkniQOVpjZEh0E95UubMjX
RMIF45opdan6+l0dFhg6XoaUrD0qhFA2I3/1QnzJtwrE9u5kLXL2999i2ZNZ/YfT
uVL6A16i3oWv0KINXw/YOiUGegglWtOgfVQkBUBrVNXhj4WXVPMBv0eII1LKluYj
i+uFY3XQqzfcSNXgMi4GatSeiGF9S5Zpp9E+4Sa52evdArQ+hHpMGF6I9+/K5rhp
tvxLyCz1HSZ4eD9u3jpg9MPoMX5jIPuAn9u2lvhXgHe76coJvMtmEAkz947ZDQkW
GzNyYE9Gn8ieJnu+C5d6a8ykJ9/WrWUmA0xG8NwWjYGkkgOhYJQdPe09471eJdUH
lEH7rLZfoQE3Z0M0gBv0bjCUNR90J+zmIrwslvGuvEfV3ChtGiPoFdRYYNQmdXgv
v68GXadat+BURy6+XCpwMcuBxBgft7E1b5YgUn1zlClE6J3SuSY+LqkraRZ2WvdH
I5PnpEc3evWwc6Y4gEP0lfmOoFQdl3Rn2kfbk8vVGYqDrppzeXZRwaqJBCnVn4HA
ThGcilbDlOwh2+uticD8oy/yd1Ge8Q5Oc9C6cd9eCw/rGxRi+e5dDn8itUm+rXh6
4cmDGIbA3NDRDg/ak/o+s/2UZiQkRShEbcYpI/vgl1X2eoibZsWFCNKnuckTbG80
1N8BhHRsc1R3CGF43vn2hdw6sSOGK1rWer0F+edg+uA5mP14uRQ0XcDBVJOqo6KW
MR8SI+5KcDu7iO5GN+r29MCYlADDM0cxEPtvlUGMuK8bkwyyDnGbz2SEpDbvH0t7
5BYY/XsI5RNYBlOhX5psU9AnPjrx9ArdVu5roqPDRK/gFFxY3cU0967fgXr6sy9W
wMrW8uwLZVa3fNJNUBedtwGSLFg2Pee+cqliqDEijS7ccxuOq6+ot6zgwpMZKvRc
yrdbljBcqmt2wmDMWGOaKInUJtYoIOnt7UwnBquDjkMcczno1ZB/wdpNHEU5S5Q2
iK8WFwP/58OU78xfnbPj6N30NMOdW1If3EIk6FgkVwyBJCLyYi7t0KTefH1m9GV2
+kH6NGM5yCmwWes29feWnAEIzEc9OVRVS2ofpBvUOWwF1JhoVFganE/9R/VoJ7EV
aPSQZuNCiP/VZ9turjI2uwf8XfQfDgvqfZbdD1wC1kIuy5Rij/4b+2rbgqzJ9HGn
ooIAwbomAevD2XpbG7wReIyXsp5XjOrnhAgllCQPam+sHgkTA2RNj7R/+KgCs9dO
dTznGKnTR1xzfq9FT5CyswbsKv7qU+4eMtGF3fE332z1aCnqgzum51GTrWtck01c
nst81piF03sED80He0X4eiOGlLubvSMij4OBd4RU8sNFgdMchXaAczN6m0EfDw28
zju5WiKUWjn1G0izCT186FWrlEnEtfx5XtwkY3tJw7UWmdXViIL7b+vGkSYaKHhq
Sb11dnnk9HNxu5o7vs1SlNEzl2QguRbM58nsNWtYOtRZ8coHLTrq+9GlZFt0bvao
kW4ouqLcJ4taQ8AdWFoqRUkKtTIwoxUIcGUP7KVFaXHBRCLyUkw8sy8d4CfD94xB
Uip/eAkh2ym2xMuAVP0bEK/UxSk/O1Si6NlvZ/ruhooresekJq82UJOfy4ilyb2C
46SPZBbOXneXXGJhLDse0txRTepisABxp02q/eZiCX1IMV8xxYnNvB8Oy4UvmVbb
jSr/onaN8pFsW3lX00IVNCaN08cDzZbiujuPwurlYBf2Wbfa6zADlq25BYXG9IES
mynG4QCeQ5TALfyoS9BzwxjMTpgeSjQLHTpQsoabw9+RhM9/XwNmj9ravn9UwbwH
6nepZK+aLYF6vagJeTN1MRkOLy1diMRfEpCXf77EQn9Zpbz6KKh+eRbAXGh4yJMc
cv/rBbHzUEHPrUat3+XNxTXa2Eplc5lHPfmVYmfQa2T8DiqWJ3u/AZFhYQsHRLKn
4r0lIkpcMS5mktKXd6YvQDZ1TE6c2WFY4wMCgbnj7TkWCU0n8TbWatEYVvzplUwU
OsuuHsWBAIjWwSKDHP2t+9VmJOSArKbRrPdWcJJFC7XO16icxsK8jIgFGNwz+378
ThH18xRYdhEQ4LzGac0KKOQwPXXZb4uKr1TJR/TzztAyBJdZavs/DyBCM+bdrlcE
7DMc7ABoIwiR9zgHQ+sEMJ8OKyksm/yjCMGup6yzHkqOlGfXBngyz9Std5S8zbuE
QulBQxFL5IRUePpikSx+QUbcU5CS/GYebdePtKbU97ceiMXTfrtl4BCbAAVZf+lD
wS274vs7D6mSpIdmVdx2j1wbf0GPt8HLIE1asxXU6IfDyfkYSGVVGcNsYMbSFpEr
iV44isqa5xXXz13zZJwXASEvXxse3Ksm9hq0VDYlnuYNiNzTtzbfz7lLJqcRsEvJ
fyY7tg/3PdA5b3u3wc2FyW9beHZRzCfc9fbkA58SU7pP0owi2b6isWUOauXEyq+O
5COqBJGQL4UOQWEVjKCZwH0N0mLGh0PjjkpOqKk5bubpl98NN6qKsHa7Ps0yO7hC
4uSDGtqJ/TIUcHH2p3PiMaK78M24z8OnG/SP3DiGBS7a5Jexa+LVm/iErkK4N68v
ZUD2N3/O30zXv2yAASWNUglQ3PO2SChg7DAfEqSW1OEnfJqZ9rVWl2o1yD20Yfzs
b3dmS+ObQttE6HiAIq1Y0WKEQSb8VyaOLCc+Z8wrlkM4HcNNDllxmko3BKPACi27
Im+p5CsAN8Dy5uofWIhxNsDzHC/VvghoEe7G31bedhQw8nZey3l8cctSMzUWpOuv
27Q+ipi0GAXlFojLjr6wcV9AVQINooNCYm0tF4ZkPMFpuEH7qFNKtFwSYofslSHC
fT7hobqoyv185PunC4rOVbwtELWK+CrMcnuTe1OYw9oJ5JW7i6+7kQ6DaiHziX4X
9+XQZDphQoDGh56mqGyiSj509Udr2tMvx5MSpqg6N+CWa5BOHJLIUcdSia2G+c+q
fhI26giw2Sps6PD99hGprysHfpqqhxRj9X8Vl6fpU0XaxcbOUUhxVwzHKiR/u34G
2zNlVqvw60irMxXdrgEbdCMLFGGSzWdeiYJlc5KskPJJ4XBKSF5A+S+AfYSZdf3W
h1gdpfTa6K568qYy5jplO9FXrzyvtv82bQhm+75VfOIwlbu+xlk8pr0VIDeW/rC6
GPBQYOTaHhuedC0XGSzCgZkUNNiCN/OTv4USxDqjulIQ4TwynMkMbV1u/fa6Ved8
BcN7Cu713HZlBGhgN5ZVZAxfm7ESqotgB7HpZs27ZRXQZz4xWyY/v6daSOeg3g6b
uzyFUYh4WQuwbGJpImErEXuYxYzejUIQpbEaNNZ1HmiF6yASjcNFrn1hZs+sDPST
YZgx6udNMQceVlLfa8RHNGzZN7SPAWXN4L6bKZxDrjsgp7DA2nRcr5v5vTbzTodd
Q6iV3k2EwggGtkp67Ym3W93o6fVhWBo/2OIGgCPqisg2EkK7/SnkCEu1QrcDS+3v
NRNlsaaX1SlRjkD5a9NFTDI98qCSx6TAxJQ6td3kaBuqFc2btuMjlsz6TXn4oVlu
xRuQjLFIvvHlfMxwBqJqDkDPExAeH7k85kAGf6t2vygX818gCMwyeBtb/lnlYSmK
sN6Jp0M0VDEV+stDjb/FD6uTPnvHpUvJAePEFHDX8yrStDgaypTEwXfGjOFeNX69
P+npRAwgDOEtUgJeWeC6s7EGoDMZjLECqK5JTXs83WPoBPR8jJDAzrU9qr+nbTZE
rj/JFuuABBm2MCLAEJOIHJm0XuwL0qY2ymC+R91t4sozLo5cHjNFQd5qBAWHBgVT
cnDtdG6Rak6szoFeMG/P6J+5b86tYns7cVTolDLfai31wM9UST8BpwoO/Ty7CJ5V
fzBM7vKDAA7G9VvpfjfJMHU+oqmxsnn+Q5pl0NndvhvKLALk5TmGB2e9yCU8OFa1
37KDnn/1G8IuNGsB5eJtD1cMi3UNZL21bMOdGHtLT8hWs1UPwd+kx/cklLtFUe9n
MnFwbuaJs94YnIvMWNxcTWQ33FZzmilrIqJZGtjaTtQbgpyripEq/TKE4vh1v3X9
CpFCD9qECG+k9HZn0ttkQpel1tLg2xfP5RBXClfe+QfVDYtSoSDhVBdqm0NgWo6w
ta7edvI2c1pdLQYNJgxxD107JLo3uK8C5CXZNcPsDzgdJ/YOSBw9rpaiQOIEBdHs

`pragma protect end_protected
