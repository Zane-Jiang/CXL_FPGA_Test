// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OBsoIMuZGE0h8dFkod9cjFwxCw+TlHxEoP1xJZWhX39o8d54j8OmMhWpN0c/
mHSgiJJPucDmCMbMD/vG99iA9hanJvGi+CCHaFgjegTreA/lx1FAUQ53Qbxo
nTImPpMYwiPfMMUxD0LuLYMAbpXScCfqsC4NVN/aHxhsJ8Pc0Xg9jlab61qU
voJQu1BhQdGM2gVeJ/iGyzswfmjxcqQoRIZsCic2nNexHi2Z5VyMTZ5SQQeL
DlMooWvAlprYYxJYABkYd5DZWrenyX9YoDWVqMxt14BJWGSoUYxI5roA9wjq
TxkIhxvM5yRmpY1OGd6ZbSPEV/aH24ffEWW/PWHS4Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jIKk4xKbXN0/gfCXkIGRdCfQ3JByeYUFm3CJn6EV8iUg/gUksnb0Sj8smd4r
0Qyi94YfdlaCPPdr/x0RxJ2zaaMZw+Lb3oklGfQ7DNFyO8cCCx3OvDK8Jsbc
pQz8E5oUBI58Z30g69bIySQkmaUglFZvkOjckiX0LyKwwftGDkvJWMQ5W4GS
Xc37Q5HgB9acnjhzpCkH8/45IxmpaY00H58w0WQfnIkh9lAk22lsGG1n19Xa
qeRiWTAYPXeEk5w8nDoNFn8MO2+F8PVXpZOD/Ki8RcK8Eydh072TRwgA/jAW
R8y4w0MwnTqzmTafB76owXNPOW71/uSpRtmvgR8IdA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GJYYK4+hAuSg1IBFZkb5+ltIrnFE6pjWTl1hHyLwal3GpJ7ZN82yJPgp04nc
M5m27pZ5txzql/XX2nvN2FjPBoNicAFwtRXgL3Fh3NU1peJNTKkVkpZ8oY5O
4UVWMTH3mmQ5Rw03FRPF0jjxXbw7OTpD4w1InEcuYaOxGADx6MQ4GX+2MWOz
Rop2gri9anhnjt9QHNBgmVBmJOxrVlYFULTD9AJEiMC2Gp0Neb4wbZxh9eFx
y54/1i9fe4BwxcUA/CM3yIlwNcgIN/3PJAPtSFF5fuzIZa7n/juGjss3w/6b
XIdLwxI5HpDW/XriQ41TKjGZEJy17ZAkW95D62869A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q9pzjrWnVNuPuMOPRkqt73XGILTXIh8CJDZi94F+3bB9HADgHbQlz0J7doag
0wGNKDzuVqGN7oBT+KYa9njkt404ZqiC9WXOPdoBljtLmIBEZKjdGT3fFG3s
IIE0LZsnYSk2xt/p9iius9bccGkm/9YnipXxtJzjN6RPafUEqHk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aXQqsvcAiKBJlBxgGvGtJirmBr+S1D5Ml3y4y+3pBYJSrDYcTuRNidKHGlMm
Q1QOSdlkCKyy2EbeVMhCLnYqlgaR9Kshebt+Dl/tbSfxM/FZh/JrFNcU+a3m
n66j+bQC8HBRB0kqQ0y8gb50AeOi1gxjz4gJBYrER22HZKNurpnS1N/4NUbT
HCp7HaV7DODu5G07QyZ+xaVKYlo3gj32pcPunRW0M6C0VysCgmdtNae629hD
RqdeW8veS+z38TXSnfWiz8lDH9Q9XU3WN3vRU/LBsF2Hle4x0R2z6BwlkFfL
kCYM3aXr5QzuY0wPH6Rg0K7Fez09G3qJ6Y1vewcsDyGcc7w7saYz3fgGxSAc
3sp6v0uces9OHwoC77drrc8FbubTuNX/jGUCMOJim11Ym/xWNSfMPuwDk4c0
Vn5fYpkcgM75t9tIMCT7cjh4Z0aOi5nxvt0fzW2cC6XGBxJEx2Hz3PAG6ZOs
dtw8UjZXc9AN5yKo0ivS5YYnlpC8lLBu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mjsZ0G1UVtkiinvkxN4TELky3l6en+htJopK1rfnt6i9+CNzlStxsUA7fnhr
csvTzgsWQIjM7g8GlYy6yob0et/C/9Gy+W2vgLKSUR7g0cN28ugubWoKhQqS
EM+InwWiawAVWrIUMV2QhjyigPdTokJ2TPDkdXwYORiVoC3+7Lk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q17ZMZoVJ8xXVHrjtbOnV9Xkuv+QMPU3Yl8y0jBTNX4jV+TEx2uw7fCj9zAD
vKcGzdauT7ZpW1hjuxc7WcEZYiqUtqJAElFQufG/4kF4yua2V/rAQgfSu+Kg
Q3ZTky47gfw47Fe/u26gLHtCFYS1u5iioEiDadQvNdh7mSq+K5Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
Net0+Mmj7Srg5t4HPn5N3qorB9KyuDPgT21EhXq7u+KWHTJz8YMD9TY/SUQj
XQzScwN1Sg0guwhxIobF0KNDuWnT2aGAqbJDaCTZIsWLtmPkrIa6SsnfKH2F
29hAIrbRReOtUh1Y+o13kU4j1CySRsAw1QhOgKWGqthdWakNmAp1HygofGGR
E6tFLcw976SXdEuPd6Y6OvMLdOvKUW2LNrQq99Cskqdu6xQ/QEEGzLtHPQz8
ItuFohnOLI3pvO+y7LokTZmqi4GG5Q5LRbJkrdV1aV9iQhNIq3wnOfIa1p3q
TSDA5a5xJftYPBJv77OoE8yjC8AeUHCzkVf1eyoKuAF7c0qRNcnRix758Zow
bvVPgQNTDK6t12GuRVKx76kxfsTo+aoIOrAQxd2PtMNUkoTao7aJ0yKB9lOW
RFtFEG5qLxwVxN1wXy2yfGB//5mXLCLr4bL90f+JBskABj5LO6u5PgN44Dq3
zD2Vvma06nxU2I4bHmC+8esi+PsW0SC2h/9PDpNMjXrmF+KWJOVB2mkZS/7s
JZ6ZOZTfgpddhJPEic6N9DMFRow0ZMpvoi60XlAPWVqVUFh+1q5DKQIhiaBF
k93v7VrFmYKu73xtUdvUl4RbrRUCXf/lNo21ja6tXNtxKIq435f2p/V/mEy8
hD+jgd/pjgY6dysF6Do7NkYBLVpYp76CGNU4Y1Ucp9/CV3hPOca8o7baPn6S
/uLKfS7OdWsWyzpFaqxN8jZCewOwQbh4mlIsAWX8Kt2rSUqwclpsnGinPMkP
oyg/HXndPJAFJV77tQX6DBF2j7Jw4TXWXy6/pHP0plRQhQSj/iIhsDIafg78
HnN4g/m89PGjChutLx/rTmpmmfcMmtgqmKfRtWFu8vEoZVteMBhCeuFiOu8/
PMBoxrMRkpqsGU0zTdC9CsukAGB0xNhpE0trnXXkuPYlG4Dqwn/Y979G+a8V
CPEpKPZqx3Iunv0m7Xlp8QWXGMdC8dBQ6S6OD8id6K2pUUvZW1GxS/qD5wOi
2D9aq2FIBDiJiASPCAwMXiFYcVzANynGFqNSKgli45yXEkZC/qhvFMnfubtr
1WZ9Xz5eyyZkJNK0WNSZ/OZ90iTv0yAyiPvEwwvjh9/SB9sDExPws5R5O6Tq
MnfQeQSXgMpjwpbc8gYIwGM/2b2Vs5g2WtT8CPgvu79QtIMXQTIG6d4mfqaY
lLRS/d/WhFmIZWaIaC8U7Lib4J+yFhub5E2FVA0bThVjuYcFoed591fhTIZa
h88QftG3y6fCeiME25edn9j42Yc/LFAmhlo1x3KdTaHwyGKVWy2DmJveZwWR
I/y3sVpWKrFTmpTPZ1qpdv9RzYO/knYTsV9VWYBQCSlvh1g8YynzWeL1GlJ4
u1EUZow=

`pragma protect end_protected
