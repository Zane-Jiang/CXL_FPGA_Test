// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Cwc7HKBEJaLY3ZUFj+2PQkymP2nHr8MUFt7txvV/aEP2aEpBxZP8gQTp7Lkv
/QqsiNbJAPAiGR/hStBkkD2N4MSesHPK/YvlRnKbW0rhfR9bay3pbDNUoWny
3ytlrvpOHXGjx+PMaqVZ7w7RDZ/LiU0zfkazonURFpbOEL4lHFRlyg6s2Ism
rYJxtnDBN+r3rNlH4fbHWAQ/fDQFShQCVps1y0bZ9xgAXzqLh2BaNNuqD4QR
/dD6BsMZROdGaek1T4eNb7v2WwKg73cRGVpK8R85cBrEbqLBM0ZZzUKbm03N
MR5SpnsU1ah7qHalXUf9axcGnmNsXD4PX12quK3LKA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qSxecFvhnT9OM6Mtpe4G1RVJMlLQsKPPKH9tTw4kHXQPe81R4DWUA/xODXVP
OjSf6iNXimkH+kXbO43ZYXjGSXsL31n7UXn/656si70Nf89+nifAkvrXE5SH
OAKY2Ib6quVZiAxNOg/4eOy/u1pWiSDhMSTpWM/KltBvGCec8hKHsjgW+MIB
Wmll+6ENVZH3NqjKwrl0F2L0aEYqU6Hw5G0uVAdyicMK9liN1XS+PxDMCC5/
T3a4Rl6RAJ/HuWe3SffXlL4Zg3eJRlo3rjUuOnkHYh55TqqObfZ9bKiVD12R
czm7EkGQs+o0YAkPm+cM2Tv2qOIjgs0OeWO0X2ouKw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Tp+FEpvqF0TeqbtaOrQ29ojF3kGBnkzlO5oh+pAIG5dFm4g/StsfXMa8bPXd
wstWbgn+e/oGL+GZNs1f+SYCIcLnUJkxAw+dZFX7qyNLrsd03rg6KV5Fcv67
Wy0xTSqQzGl/RLN0kd+ZZY3pVMa0aUGQ/TAVcKYPEH7o7wmc5Z/zZxkTr8mD
/uj/TgoQ7T/55uKc1k0DYzUUJq3UNMxf0xuE9LyTjdyG1GG8cOE3bGK0DPNb
3Y+3G/3eIDNbyFSEN66zgxCN+GN1TCBL1LYCCqKRd8qhslATxxf9OvyK/1No
OyeDwLW8X64tcu5vpJBz7P4p8WOoNXNPvARynkjQLw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BdxLveM+mcXzzGMbm067kt2yRGij9C8fbYglUflJ03oAdt2y7rushA0YfCjG
K7C1M02nlh24qjlSaFVn5UHi2bbKdA3Zc9vOb9kk1zv3zbCdPxVdyHWLsizY
pHflHR1TGsQxog+HFa8DzN6e+KDIlZU9ub1bOlme8pl9/IAswFc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eXOLjNVZqjNRAHt7EKJ3ZArQA4EaGaKxnhzkfaDq7Ft/aMrMBFNbwjrp0IsX
ZIlvH6PL0NX2QBiQPTJTkN69WsiZNhARiH014R66N3P2Rl8rSxOBP6bG7i4n
yFxJ4kuFgjbo9R2JEtx+j+UNO4Mol+NTWHAJOKAZ29wiviKCxAlwsbwuwrrh
baMWew2JnX4Dk2+StmUA44RQnuir0MSR42fBuvoJ4kEUHG+uZmh1rH2Btcta
5aXmgOKUrmhCzRFnTuDw2IxKD0XrQO3HMQhFxm2NZgi1Q4v+JUmOjS1jtRWg
ZKBsKlS0uNxKte5d//kMz+R99G36P2/O1dvJ9v1NMORqNeqOZaiNUfbMY8KA
QApwZruqCYM/HaBC5zbNWcMemynVJSq8i3Lk2DCZHQ8w5E9eeX2afQ2vx5JT
NHUJ67Qfsp12Hnd2gHlMTZfed3LZAcCL/XMwYzebT2i+D24cdpn1WMUujRhi
AEd/F8C29FGGZNY6F2Ch9TWyVl2zlTPc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RjtrrIpieG3ZPQWZ7XULPH79tMW2rlJo25XCUuEaCAuiIvt/B4EUGydy/ziR
BBOiNGDEOgvR5nn4qcC69G0NnT45ugDlF537Y8qv6f4Vl7Yinq7epL3PCW+6
LxnwKGcIiE5T6omOoj5Ek4FHBGZId8QnoPB3FCkv+e7lqF/js3M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MshooXTI2QGhp1EsZ292MtWdFvTlbwm9qjZFlU3enSGMgYFlwMr3DoSSx0fT
OBGXPBpm3qiTo3qnldxhM0ogRIg7JLUZLNauY0I1FwaykMEfaqvsiXEwWk80
gV1/neFK6lMz/4ZfAJQFh4ljHyrhg8RFjLgTG2EiY8i9C6qOUso=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3232)
`pragma protect data_block
Fibgw3s8HizSV8At1PVILPqwbUsDHsoQWsazw2mitkwvUtARzw20uAoClrqn
sEdjMsTtsMcTTFGS9E8tM5QeTH1TvzyM9cHhcCn3DEPEUkVyZUN5tau+/Coj
ptNwG/fzSlaKuIlIH1bshibahA+jP0+2I+X4TliG3godDktLUYxyffO/UL2d
kE5wlG1cR4psQz7bSJ77J4KsQ3GkW2TY7lis7VRytopjmy+ZuSsZ9KTzFS1Z
hmKi6n7OQN968d5oz9SZwL/onEc8KiRIVRkS5JEMFELpYKzEfR1s3Pbg7/ve
a9d5Gu8aCVtZkK9AFNU2BytySSlQRtqGEaLf9iGw7A3ARrolQKTjfvfSklUD
cEcyl643wXyqEL2CxRMM7WU7cOc1pK7AzOSToz0bnbNnwwZQjscARbpXiCYr
YYnSXm4LVtS8jtEhVJ7QeFtft38l1uhFtQ9acnIRJ5IV2VEd3/Lyn024RGEP
l1yI+IkyGgMv2qTixUDttwxNV2rFCe0TkM6GplbwDiRqvBmwod7q6jDpDlyG
tfYKRTiP29H1LCFpZjNd77EruXOVix4Aln/PkCbZSBQGA50RxxMhXASCiGOJ
DgKcB4AZDCKNwkdDzMCGtDUmpi0pJ/ENcigQIFRGqQ+UsnTM/rpITTpRsNGI
q2N45JU8Z2oDWR1l50K5aKKDpG5NAJHNwgfv4qT/+ze4s1R4aQJdWpkVS0ry
bJe+imejyYp1Kix6KgtJYvyFmtX5omtKbR/RI/HKHtD++BkH/3gRTm1q1y+f
kQ28Ao/z4P0LuMcHosvNg5Bn5WtjB9w94POxKVqpXxzGCvMmpnFyjdgJPrCZ
NlGRpHzWfNFx3XidnTS7dVJifmh169xe4wL5DuGOwoE8Ukv3WD5eJPdcf9ki
NeY8HHir2dlnEsJQip0F4kgAK5cHLFgKDHGXqHKRyWtFukFgJngcKOsT89LL
HmBuDh52VYnPd+VuTFA/G7THDBPcxDiT+V3dkYdldC0AdNzU1DP+6FGtQnK/
SRxTJUaq90T1leR0kG3vHmxpWWK5QdH6kTGfa7gP5thAtyDyrQlMJKgQuDt1
9/bQ21gR0DDTZMLu5P6XtZ64FaHEl1+3PButG9Y+wfC3abukmyyU7qhHarka
iFhxHSunFQLDy1x/NebTbKnr/DiLREPuL7tHXCEiNVkUy/7bDK5DgEd0g16+
RDzjYpg+mkOItkLaoG8ikADOKZcIIPaBva1V+wY2U/qnhFkG7exU7FCz7B7i
qtb1I5oJ+HGryQDKxOxB67gWCbOqy31H00rsqxnim0HgjD2mS3CStriDp2ui
USBMRChCYpUp3BFy3VamJ+Q/Y7KsDdWsGnJ+Ysv/55s95TLPhTmTONAoa+jS
JjFZ51b1Cn78Aq/wcUEoTlfiwvo5kSh5KlEh4fq62jjWYhO0Jyv37Xg3rue7
D5uDo1OAskupN6vTNXbaeZ8/t1Cldv8fGLpBkuROr6WyhMPmaQ9wXx9c/DPu
kq5OQb4dv0Djl7hNf/SkO5/IWDUOTWEiVC6qLhA7Mx87+hDF749Aj6UJeCbf
XyI16cSR8WtoTdjdKlmcErFTb2Bilmlx1nhglgqHJrb1Pe6OtHMwFgRsVf7K
ryR/iRILSnWB8IgCZxUS16DyNlVihWfWey4RcFJKMw32IoORe4eJXjASUe+l
3WjJw8ZeEPi6sSTiNgAue9Ijlao2/FU+6Jdh2EhA+cOZw7pCdW4lLHqYm9zd
hZ8RPDgyq5cBnQXh69IvDfET5Yc8Ele9dUY130TV8f1wyPMsp1eMwQuFs0lt
tFP0pUOLQpGYyImq2GCpJpnXFWmGZ6pXMVikdwcCZsFjLKlrIjuZ9e8tL7kf
zCWvO+5aIxIWzkT8ww1JAdFQO//cJ5BPUNonPtH5T53bK2dLGoD84r1QhJSb
G2fymW784sO+8nmAWmVacLhdJqUnrxb8ych9eh5iw6NSun13sWKlPej5yP0g
4AAPKmwHr9UA2uZ2xqCvnoHowwn6PvnJYfQfBuRKT20T5I3FQhK5oQNZeXFp
fWFi8S1e3DBt9HzNAkveLc2OTUOVO//OmsBfm76j+Wu3mY1uwUB+/HT/blaB
oY3NIMcpCoycxALe3cDa7ZxYsAgLti5ShBFdgCvCH/RvY0xFpREABigowm51
ZxfsZLDKGxNpteQOHYen07Y0TTKxnJ8cf4NUZH9JW0L+eOVUZr8LklSptDGQ
SzTMyNZDYC1oMJ6/aTi1K1gyYuMgxODmSsVon86sWvX2y8UoYUMl01GjTwdb
yretI6WLh6e854+T9bBAhCRMkByuMGIYVIDc0Wf2w6kCBdbtk2NrO5X28F9i
g9zFD0vNHqJ2NUzHU0mvslIAQFhnjuBGBISV8T2JD67FnkSOI034+FHumCen
3qjSr6vwx+fvNEszCdSw2SxzSp8j1KlALBymxAbjthh2tI6Eh2UUUrCrjGa5
SZ/MwNYzR+hFfAHMFpCEquKyh2ZP0RtdyznrWoIBnN25zUCiS7kuiUcVFYXM
wdPhqo0/IBn2ZoWNTX4V6Jp82huuQc1bmWfpefveJ+xAGWey8UwwaHFCoq08
DMd9ETe584ctxmeOhfsiuP2zjgfV6Zb2RrqVBXIypdqUHxUQbE+JIIcKAmen
CfyJi/KAU1XUgEC0EOu2QN7WHPCzhjxdsZMjYSw64eqQyBFSDFe2ZSbVG+3U
JeB/BbHIDUQ6fZmTMYtUUH07vMSC3xqVcvyygYga0QoOqprRLYPKOXvhUMEp
ovq0/NLU9iNvDKoNU3AZigd9fSsxu8UeJmza+uRiqdDi37oldKE4iRJyEwP+
TJu4PojT3ebjsqeBAGfJNrL2AvI8MwBF+wmh6z4yu3viiSZvF3VQXa/LpbVF
zNsa/bzl4ZclOwZo4SgM8kZIUhQTYsOUYDjSgmwQJ/h9oRgUALEfLtrtD4mZ
tuns7P6VWmrNMGvE66WA/mPVxe9CYRPMbzS6ZwUO0jkoepf2vZN/JW8U/PzK
SbW4MtiQYy2FbwcSyLMtbv/qQv3c36jOlydZfmoDTYBUYJHhe3bk/Ro3JAxI
OwzeIOwupi26Y3RmSsly4YtXTr+gvGS9rUPCdvQa84eXc9/BvfG242qTARLr
3UIyE9n+Jwgo45BZL/2I/3Lh161D3tJ+F68ilFlZ8OBJmwfpVTAFnKxxZslG
3+MVQkuULIJ4aQaPpyyo201y7Z3NMt/1A4nYqyg8S+HMREdTVNHrr3q7xpuV
vEiONQeqXqtcVqgHkCRjT1mMUCNaECQtufmR7aV4mOwoZEH9Xp7BESTYaSzz
sG1kt9OWV/ssMIMzWIBXPBQPIGsVh3GGFTxIGKAme0fS7oBMYyA74q4X3QgP
kZvXobnrPO2ttYivEDHOt8k4PVyhK4yTwcxH0C9hl8U8Z9zf/cTNH3CeSu0D
+8BzKwKt+nZ378gCfXUnl695K63B3jUwB3/ATetNsu/1MVySqS0NhN3xpvov
Rv2YtD8AgBJMP+zTe1m4gAm2TTn73IW+R5ukrSFpY1Uiv7Tq2vwzvcZmyZWN
EVybOyxO8iv4r4P+1saZ8Gaw/HvEymF+6yTM8m9HxJH0FCyH1WBGMMVznqvR
QahV8PRD0BJQSKRhXab2uM/YeJMVSxCy9//3eoTmB6irlT3QCykU1S0xD78r
Uzaa+JHfX+V32QddaU+BZer0HFY4uoafzKpMexUoUCSUjuZXqLVQZktZE5ym
CouDgSJ/P6We0qYyeGrztDS5EIZpn9V5Ow4f+tvBguBhhBqr1XTA788G+I+X
ITKgFnQ1kuIjToctVjvCWOEWHu8K0sy3B5bssdkRvpYbhYJBCEG7IGDSGvuP
DMYaI141ABjLL0Mqd18ihPHf8zvpRRVIeBAHWBNOjKfTMoYmENCu4ilRCLvz
apclfMLN3cY83RNSvEjT8Hqh7uxdzsO5rZh0cDJG7twoy+YXuMkQmaoufy0I
yqTB7Kow5qqWoPghq3Jr86Ixn33ASeFmfVogxaW3MR3L0dyoEfWWIEP2sCbW
T33xrZdibTea+qohV6QquRQGOlyYgWWbdi+ZWh5QxSAqwgymJYKHe37rkeee
86ubwbdCxwEuvyBdHoSGmdxJqsRHOtAIQ47kY3uS3OckFdwrVBKjycXIXS3B
UvSpdkIeUrlPmWsDbXs7lbWy3jchsscfFi0+Fr+S/chYXZ2mJ+oCvEIXHD77
Z1zP8L08AfqfmiAMwbqaV2GwZY/dhRMwli3vMg2ZOizbuicH8397YaIc3IH+
mtkPXBrGc7rb5Bmj0AHhEGgNO/DbkHN5R0jR3JTcq0N+AQvUPw==

`pragma protect end_protected
