// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FYBlTGWuoHyl1gv6ZzDD2t9f40IIXLtV33HjIzPkWbeROowiPFfIdsdAHapl
y8YIOYG9pdCHuvj2xjhxDLUU5M7coFSZkpjmuZVlLogUe9rp5373lYwFMqCG
YX6LyZ1DBjFdllM8YKf7jlQId4GSJjXQhemwNaFRnhZcLyf0jo+4FT0pQ1o9
7wdieQTTIndkKeHQ52G+co1gW7QdKSJcA+rkHXGSf/pJkTvqkAdgkPrNSrVa
/ytE5+oVLDchQHQdLHr8qScji1yNiB2zn1arXy76FYCE6nYvtIPZAP478/gL
KWupXqRm7JFevv3xaJo4ygVZZ5Hankkh8cvE4Zkoag==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P4OEZ8PihPeszHjGjWHWJXJZ+mAZl3SIByOuTIEQpjhglxzYRLRriJoe/96O
4rQUSJrmMaUOXqpY8b602O5ehztoAe1MPOFAROKlcoR3IldyhF3kcnOji+Fa
8LLl2r6+/Gl1Y0XnEeOnSx9HaT7txH8NQlCYy05pspj1MIL8vcuXxntAPFMU
5IlQgsAkW7kXz+0v2CbFf6uwdAXs0q4VMOqJ6frFD+R14LlEJjIU4fy2GBX8
LwuLT9Rbv1L/n5j68qYXSn8x0LEeFqmJGgqdqRNSiTixzl8PpHuQnkb5MC5S
CqFmhztuQT2v0RNlXD2QfpTn/+gMoCjOd5HlRU1e3Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i7ST7sVgAUeFVHFDTo9Svwz5GJ6Q46HdsF8LlZbpOJGwGRjTCwZQyADl3Kkj
XPRiy1prAutGZyyKwpnpLReZcdoudFfED74Q169ctgEx0PKh1JlcN04ow94T
9Kf4JR+hr4dCuMIujpI3DdMqMdcQJFWVv+0wc+Pef3jE5OM/eeCQ9MaLECHF
KgZpoz48GaMg5sJ/CpfHdvpKE4SQWBOnJegRobt3DHo8VbKHmZmfyDXQ5Xmn
p/vaeLtrQ8FrD64zgYSNnw9zVcsKQ4Y3bxKaac6Og83rXFFqllvcpWDxGCxz
G7G/Ob7k1NjLeVdmLZ8ikgfvPxC5j3CR58g3o/WVFw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SC2ryLRRqRGU7S4lY6JgZwKqa9a1TOYG+zvyaS7f3bj1z0yTdJKoo091dT+a
ozcwlFo0a1IofmvOAojRV6PC5jT4uIwggSl4RZoAeAO1Qe73tRBOWoilsZwX
aYv0poR5a05mkgVUFHytdTprOlGQsEAekc9Bhx+OEzwmfEr/q8E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ewmBZhAq3IYuseyNAbAzu1fc1uzUWWZ0UHPqM+Suuh4JHEIsC2okBU8dCaPy
3X4L/Nk8iCKo6HX3FwPL8QBXIJF5EfZVIuBs88cf6fgB9Ji73PChMumIDHPl
AccF1NEzok2VeBCx6J4rWAvGt6kkM9jBlAjH9aHBoIZk6lf5qMXY3NhWCqDq
7ylGO8i6o1lAIdUZw6fBvRXuUja5K5ePhl1/JYyeUtmztJxOgLtF6pAOl3E3
WGhPJvtXVkgdzIB2IZWO9johp6IxFgDMVSp341S2q8kyM18hLrzYbk43oELL
08vdGyTHvnVXC1fZHs+hzuoqFRKdMxWJJINy+WtW5kBErEx+Tgs02wOr4QMk
qGcXg5gh5b+d1MVIdQ5NrUpZ9r5C59s1/I6uO3YD5ahsG+va+0Lku9LDYl5p
0Ww5sHDArDrV3ZUK3XtuULNCanRLnO2Z4pMmB2ggj1gWafaIUmzXzpzwH2Cd
KbX7j8Na11l2bapbufkB1aoRaDRhf2ko


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dS1e1IR9Bh8WkRjyoW5TTs00NobY3qLsSkDdzQQno1vjhQyEnHaFGx7bRz+b
iOaqgdmk/MlDeHG4v+x2VZMfy6eem0p2d06clYCD7IdHylwQDCRZjbdue77n
pYDzZ49kN9KEwU4csAraDPxCJv4qn+xO5c08l4VdQ+DfxYsGvko=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RK/R7lGPCGDOc+Ns7MNlkM9elhHbSADoEWe6h4rxSlbee5BQOsA9L+rnROmL
iSqRFFFIKBX8FNCuzxAEOo5dOfM0ybiRsmV7jHYnFb5bzBI/ytl3/xabVzln
Q5Fs3MOKIuVk2g9b6wfazmhT37laoBdxhDPLrpfb4ieazrqHC90=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12272)
`pragma protect data_block
6jHFLbgyIvSVMIgfD+4mqCSWHCaTvoW9ETTZ8reBTMX4nS81UgTDmRjfY7Yn
mIfpJYjEhTwoBlW4FeiCv/8Ew8jY9WlAf5pOQ0G0S8vA2DVjxlVKW42e9yBe
moC0oOWM4Gpquw3EQkz3B9f/RAI4rl8S6g86vyGG3jbQ1k3sMny+pfJ5Ao1+
gUT6AodvExtyoOnB7YZ3lfv8jPuu+V+1KLPN6Jws7AzoW87++veeoCrBb7lB
BFwqQRyPlF0+UGSmjUXlTXhBAhthLADdU7+ya14PMNyDVDUtl2IgcrVmlMLb
xviOkI4+bFHi/dZS9MSlMd4GF1HzniMGkNokTFCMd7YFwmX3rYTre/rINn9f
Uw6Twl4MteNjxEwTzgKqvF/hLEbt8jHoz934jC6gCh7mfbEmm1vg3rVzgvjV
hxP5+gJ/cthnURJlT8Xe7iANr+hBNgC0j2LaK1eEy6xto0n7NT4u2u4wSY/J
d29/fQjcSGUqpqhk/EtsJjTlhfREJbX4TzrSvG2vh4pe6uN0SwAmTL+qy5y6
a4gzLil5f6LpOQVA4eU/7TALlFs6hVxytGQ35deN2AusX4lmRKe+YIviMQ6i
NQdgL+OMPWtiv8CFpgG3XTVY7ozWqMSwSZ62/uppZPkSIy2OvkcP1JxzVgsa
6TkRlWFMkkWBMCT58hgI+CWor8n3ILMuxDOJK/HK2bzRqGjAuEGLovsukhji
syCHRmRgS1pZs9div6RHUebC/gE9WIeWUeE5ATiNwc0KNaeHNHwhO6oeb4mJ
GRTdJ2UmnVTKgP+lW+ZQ7+4WjVJ3dRj99opXfR+1q1+G7fJzvwHGlAl5XyI0
Gw8PrqzwZUjiIrFsFWF44gHUeTOsjhoevUfn/h9JVcm45SYpyTbjzJ+kTO5B
vGGS0tOPf1uL54N6ORX5yLhMOKvy0809k2vgS71mFUngIAXwobrJ3sbdlIj2
uaYU4lHL6oGhGoRvZKEPbkmKgODG1NRRU0SeK6LvkdL93xPoQ3lwLkLDRV2p
FOMiKSK5iTL8OpxCQOnw8+74luU6hZc6SwLEgYjar0C6jK01xaPTdJOqMjb9
Zaq5iOeUSXLNhXNfdW0FWyZxv5tEKfskMHqFoOeu1b2KDBbT5v8FBBWM/qnl
uM/+K5OKd134sFP677ts6Hx8oHey/RsTwpHetI08tCubQoRcwcLFfQZa5wvb
BgjkDBsyokW1kcCntvFagJStus00Zb7IOHQWGROq4Yh2/fNgzvwYFZRrp111
8SeM6wE6zEBTzS6F2SXYsqHgZUp1wfSLjEH1Dg2cXYrTnwrDBZ40CMDwGg4r
PS/OtOmETTHAm4J9LM8ox0hYDdtnPVowO10yzlRPuckl48waRhtVcdRD7e05
Lp2pSF+7Id1UB/6bklUJVzE07m4ulCLyWaEIkbGmZjSOJ1B2MJH27QJJ5TxX
ZXZ9n0gxxSdlTKZgdGhg4h1ff2ejhEFXDiBCEyOFEXDVJ69w28oZuHWu4NMm
DUr1df+j1zMIUL9aZi9+4YXrAAcs4l5j9kuopYNMBouCqGriaGCqgwFzEglp
glNlu3U+f5GalJJRZVwhKPNPm1ZIg97fcXM3Uq90k9Vyu5EsOBhPvrGE6Knk
G4VTAiwCbeP1BMJS6OpK7V3/Q+QWnh/a1/V/X/9HxgFg32azeVpnoNcq8R55
7PEFzbi2GEoy7H8x/OA0Ouuq9gkCxiHf7NYhHsZ+p6g1kbMWzAaXCO4TJQi1
eTuB6KA0lVB8FUEHGTbtjce94zT/Gf+iG8HH7P/2vgB5PfJYhgCI6oebhOXS
+kFxuR7HmWgdj4/thIu4NLdxxTKSN3zkhVyJiPXdFqJ8BzpQee7PFPkZdV0h
39l9Qg4LikReBqjpKzp/m7QQjCopOA82Nr4Tiwo4zLRL976/M0YLYNuQdfxT
stIYGS5XkmsBn6jvofiDPZ1+GapTYlkC2omIb1k2SWwz4lG05c06EfJ9H+5i
B7JiqY8qXsYUuHPumgFasDt/VQMjNJBGSZt985xwxEnv463FUPZFSOaCdAho
dlkJmEwx3AfoFUexSRyYenSFIZYufm9xKpD6iU+Sb2n4PHG0hVB1886Lrf71
wkAm+jLMXqCr2MBakF8DCA0UuhR3yUI1o/h6OXDFZinrIHPuo3c6dU3piLH5
cQgFJpQkUTJZspfSw7pk3m+GB+m04/5MAwTYorBc6M0usIZaVkGEAkZo8XTu
1vFIqBCuIRd+EgNSScOBV+OnrJejBjwTODWshWyXp67NywIz+1i+d25snhzp
s6/Yjf9gB1n2XOcuCzUwhi0WLSlDemw3MiNJ5t2w4/vCg9y8UBG0R8N439K5
3esJGjCzAi1wp7CbnKIF5znPb9ZeSpcPxRWvVzhbjz3wp+EDUpjDfv5ipX5H
Z8I4QLDXS2ycV+jLTDsmUG8RGVTu/r7xa8bFPxubd3U0IxVogwZmJx3DiAz2
vPUs+wkv2A+H8F7W9eq9gLpnxp7DQwLJk/u8H7OnduM0ohYZqQMEBDvTAl6G
d8NoyZMBW/RWSxmqecr4iyXuTtmg13twAKiE5WwnLyuOFM3GlwxpAOolk7tO
9GxHtieDWhSOLrJW33/k/cg9JLe55fwWjhNTmD8TihWribrx6iziWB2DAtFd
YNn1hL5kL0lRbrBgIbTScg2IVq/XLixNSUhXWJDllnwwQAcgKfw8EEtHYnyG
2ymu8PgFBBC4qjmhXk7Kfwj9W8jwJL0DfG2QY0cS2fqCVdxvCtb+LdlLC75Q
aOFT93kQHTpVZ5TwIVLrJkoMDvbAflACNMfHKVOT5xQNzReP913BelbO+wEW
tH5nxl667sNr6gZhi9Dfd9WcV8w249IbtTGsjL7AwPhVaoQuMY8gbqITRbV1
bQZ/ZP9E2PL6ZsmgF/7iSdkmdoK++dJgYXuexbswFZruXV6gjR+/3wI1+vdF
tnuJRzJtHoqhNXrdHimoSg4MdcPCVVuMagQttMAQbvfP5UH+/0mw+t6TW/Wb
HjrzqVtlROe4VNKMb1Zl2WTLfK07z4kHMDhNzLvx5PGig/rZ7rNFgRqEiM1E
pgk36q68xqmiWwe6SJ9xSm+bWQ475DDkEkCLZFzCQ4Q9mBK/2/NNrnmBFLdy
oa9JlDckZDhs4cjcuAaos+CgGTn+7aFsfyUM54CsVd4LnJ7yQ0I87Vnc/r/y
CmGSkmn8wqYj7vduBu7T78GS3bF9nOIVuTGasiPstKLK2RaaDC0qaW7LjMJY
k/6tvu9+NmOmy+ZNQEAOTHyuh2aYSsbnL/EGcBFdsXBHa1ks8ntEKGmmAUlY
VoU7vY6p+K6kpWVM8AzOM0fdEgvSSM33KzedcbND5zC2ub3juwnY+QJ2lxX2
RpV2eI0N94YgleMZYelufNL/tvKJ2kt4X6SsjMqfK0GFOBw6fPPPmp5moAKB
tTSg3BDbTAZ8e8cyr8l8zeP6TThp1YW2smkD1WjcIfys3/t1GFWoS9xAwquA
HxEyDpkEmoDShNkuU0w3HZ06eCzab3Aik0TMFfqFuHvLIMD1yhY3aT4NBOqx
eoAi4DwItoSlXE8PR03oJogd68zhKPWCdKc95ze6vJ3vVvyhorZKO4J3cfUM
ihFFGN5j6ZdkVci6xFtJpqe6SaGuxH8RhoOrbB17JXPQQGViFNvOZ1LEHSjA
JAUyhhmBilnQIuf+ZiLbtFhNW7+I3kpfkkZal4LPwu19684wreC8WHe09TzR
DZ8oOXLTEBetCvQM7ApNCFEOcxJcHVXdb22xdF/6NQMuxESgdprubCHbfHzS
o0eC0l6l3YzCW/bP2kdknf//jluQoTWDm9fdo/VIlrbC3/5RO29iOBVtgVVF
JDd6JJoZsygaA6+pN0IMzYmF7mV0+PTSM7gn7g/yhL4x8cV31/EuEMdQn907
HfeZ1dfnaSg8m9nefHzwaNIquoG5OdEGTKRSiYZ8dPfNx8QgYQPtvNvNI7Lv
owH4UqzvlymmcDCMeh69gBXZmaiDXqTkK5djYAZeOJirGI65+pNO8VD4SuJu
s0hriWmga0dDwo8BmF5UEs04qHWquEDj1P/aY5Yn7zPcg5ieTanLnA8eONV4
TwTKeCQlB/2Ua1ERHVvyXhjQmhrJbDUVERR23rRncFvhNj0GqfVuQL+CCrz4
AebAXtE6DeBqVJXMwJMKFco7hvkaQA79XiOSgiioLTTrlulVHx2FVeO0SzWg
tKKaX/4f2Bx+44GyV3HwoizpJtREx+n+3QTiAVFL6+4r3Qg5kNH3iqGuIUe8
KrRO8RkXpjoclZcjNAD8bPeY6tUTkSdtAnFC98Q+6bZrl6tDlkpGS17M3t7f
1jx63ymlFoaDKKNPpr1YoeZOkcC7pvlvSgLL63lqV25tdw/+36ZLPdvEktJ3
H8jGuuGJrHlzw7mSKupr2wpd0u4nXim9fW2ua0cUwvCO9LsJaEkZj0dIUJnY
2Pd9yGO+QP2jOfJLP6wRqjP78aMF3KtkfKFdujchcI2894lIXdN7gWJPa7pz
mPepDxie2doEyP86/83WtcwVVkmz6rWA7P2L7RiliYvIU4TNKu2/VWg/L9Rb
5K1MzwgKt3XKxFys4/lB0R6kVgokqZyJmnx27bQivadXEQUBiNSWSIKBlxsD
9zT8EFssJeukPu4A/JZsGcs1c3MHqIDHRR19fc9Be8jswr/4+spfF4qY0Djl
TcEz56UyZg0aJfNhYcpICF1zryc3kxY7upp5mnEZsVDppdhg7/qvdyByWfx+
QPUtJJ3HOJHhjjmfTQtyOJFf/CoFBILtkNZo5MPemJ+TjcGLcerJQu9A/K8h
h5rrfrElTMEI2NH5iC2Nl1IjA42kPRaw0w9Be1QDxTefaGtOLimfrSNRfnN+
VNuGmD8pd+HuRWQ5ZkMIqQbk7vz+vtMwtQrRvvlm6HNQLpONhVHlGScuBaw0
BDlJCXvxYVm7LolcFlgZVVMNSJ1ScU0yqDhZlH8NCSXKPwmrgls4QCF38K0r
rzoNG/nGnuKesXf7IgkCEzGHDLaGRR/A9TpOQ3VedgaUjTBkKkAiGdqWHWUc
8ryAGnY8c7iaVWbcVdSy20wdCh16t+USohe2khgmueObBuT0RW99jfBthq0h
JzDiR2rm9nFZt+teCp/+FDwaLnOcx4x+qrFLR1rezemnAll573lA3WwzFhsu
PZBuOxOGb8C8PujLsMY9xO7J8psyIdexBvSTEgKMWkQUh8+fZg1K+oNKZoOj
bZs7JxO5JBLMTGgEEnEfkgPvdL3C8fgbpLoJnMDvsSiYSLzi34eXLbLMZ9gr
O46YUsQMcvchOCBqz+WDBCCSgKFYhTQlLrAJFHoS5wqnKUmpCx4f1uDcAKUv
1gGMageT0Qh7eZ1JerzeNKiE3858701ING/2T0yF2kLru6Tx999m4CzXQR5I
4/0ujwNH9vE3DhabzqIsgHl1cmfElXTPyhALgfzXokmzqb6T6CNt4AY3qXGx
L7Ra+dV6n4nG7fBisUc9UP2aguoEPvU8BHcec1wD578IUayJOgWIwE9RxMoy
CdhShicFZGiAUqA2sPBDgzLyCPtx5oyGWREIDvmUtTknNe50p19Rifr75keO
x1uJJ4uxiQDbCFsnt3UYlcYagg0WwAa97OdDMHqyTnJPGUoFdl9XQ5sUBLqQ
3YdbeaTq9ARUdMy9NNPyN8rvp0kHIg1z9WlmBukNQ5xcPQmizr2ypx/JuFMM
/SN1qlkuSePLp0KVOoqqyc9Nie4jm7vPm1YFM5EhmexB2YaigB7RuZeoJR3+
Ow5rnMEw1DA12r2bImj7deFASoqINlIiYNOeRbFUqC/U6eOX4xFgCbUD0GV3
xrHJFQFJ0L221p+yz2Xjtr5P0ESuuIPGI1VDWRkdNI4mLMy4Ky0l1v242ClT
vkwGDMDEY7PNgWloliIVx6AglDKF8XceokVG+r6pzVBBSl0VcuJ5VbT69q4S
84JlZtG+XIWaVsyhV6u6uGVImT9RpLilwNVB9iohyWqUhX1woS7f/b4v/FhP
Ojz7sl3q1aQOFK5gqbuRTHVvCYRyrkyAvwzNMfOjq2Xtx4XjevImjoG0klXo
nPm4P5l/hs8EHMPlgeVm6WS+UX1u3zYMThKFRm0pkl2wlq9MnndMdcistfDY
stdfGKEomsdGuvkmqtNLmjFUHTG28DpgsrFfKo+d4tXLYEOk8upxXDCaEJG9
EJt8x9PNVkSGpqYLoKxG94G45YSInJPN0sLAX6gAydEpeN4wcZhzOHp622Do
WZbwMAYBoYEe+0idQZMaiGNMmkL0c2LOiWYh3t2ut9+C29+ZxQmDUYwWXoIG
Q2ZZcjY26qmGP+hitQcfnJlbh2zt2fc65HnbWkxLTu7x5k9zEuqmrQp9kF23
Sx+U/MLx7hjyS85dZf+5kt8XWhjYkpEs0I9UVhVi6+y7docLOcsK+5U7N3fJ
pdNx9WifDlISwSEpRf2z+4gXP+Ve40d/R+uNUpFFgUVy6AVQLlIU8KAXTYDY
XoClaRzFb2UyI7qLWfjNwCpJoDvqk0rBIgTGKHrQHCtbvMCo0bByIGE5nmdH
lBMbq7hc8BuxyifuhDGeKTarRRYt6sAnNqd75R0bWFe9shLvaNGI2pPTOaYu
xT8c5i2AopydqiGYF2NX2R8Iv3TfyeHmia8GCiWeC1RBWZMsisrf/+AReUh1
Xdod4M1MuITXWLemL/+ewW/f/s/BSfvgRKAzF1Bat40Pzfw1O5EOvrAN7ObN
iU77YT2mA6MEY8gZLANi0A9p/8YW0PDIb77FE8CZsBHK83hN8ZY2CvL+1S8u
mxONSUHL6Ol3C3nbDtis6gNc6HJm6oDnJxYoQlsWYAmkh2tMx7csJDZdz19c
uLzul9FvT97oxZCg55TS5FfRSC9se7c4/8v1EyktGgNFZuWQGuAliepbwUy+
BAontNiRMc5ezhrpN/GuvkJ07yHmblQ3f/3wBRtUiHpWF3WPfRnCPNltUmFk
gD9a9JdSrJ7lmRms4mXLy9TBGRT2vTA6We0HLVlAesjAEl4zdRy5rHPe5hEE
a2vp1ifZxszf/nop6NGIWq8R510Gxd1/fIs39oMH+MiB+6aEWL80XM7LKVDI
nqYxGoTMTCT+CACxRBTKTfOryGJllA23s4lkOensmZGuji5b184KmX/z6ziB
EgAs7uc33mrNiUlNb0D47DTrlbI057dEEz02qKUkWZNjPYEwNAPI10cdOx6H
FZ1/lDTL+Hb5BwaChAxcOw9IiLg90QKe6pCCQQxRNOd2Qt1kNY4Fd37d4ToJ
PoG12CFUtcb8X6yEP9ciurBXIKwHQ8FHJnzgSQI3VVv6jv9iT8v34O7l2xqt
9/a7LCqRWCUT71R8TXOnU4D1yyZaHCwduNFgbJxCxxiP3WVh5hwKq2Hn1z2i
wCAiQiHCsjebsHsuLzGPgd7lPk+bxDTjB6moptaapzuUYGLXcgmITjFaqyfv
iK9b+wZMs6BPvkbtabt0R3VG25xwqSXSkR0ZpU1cSU8qkavTZPbfC/OvAYQA
HLyROTImlITchKIPeynm3YbZmDOXJZ5l+HQnVPTiGVcxP5GW4jELOig8JcS3
qdPQ2l3r0q17HN84h/a85CbHhnuhQsfc9JjifMrAgegQDg4CQKsZtEDkPpf6
9B9CaR8xbOlr1ol3QyjigxESb1tcWMGa/pX4XO+10pOmzrcP36F095mRyOXw
WLIX8SN82zNenzsxsZNnW5CdVLrA04RZdSbFZxegxjQaViTKg9tbTI6Pw7vC
Z1cwJtp6mfbzaQE6BukhUWjfSoynN4iw+RQqtFREQUEiaO8h4HCZrI4rDphZ
Ow9AsmtWcAA7MlJBotUFZwDHQoCzoTV3oCHGEywAc26rabhPvxLT7ZJ7Lofq
jFqwypP6pyjbGwtNwWgwt0i9mYIpdWMONfweZ4C5YwoaBeCrBPU4FAGySxMM
qwJuTQYTlzlvQupHmV1DBrzrmMPEsgXPcQOH6hCmqTwet/35JVb/oJIZe2G9
Z7gXHwdfvNhT13jD5aeKa42NbUGe01DN10EEuEvq/XkhNeZz8en8QMD+TbXy
Nd+ANDrDk7h81XxVAjGW/4ojbBrgvRNYiZLLC7wnZFMhHD2Bt7dkQUboRQ7w
N5rydGE3m+5ieADeyim0yRKUF7r4ajh6xCJ1pDeawDhU7GiqARK8e+b3BF7N
CtxamtuJuN+0x7fSQRJlzTHFeRQjr+SU57Yo1m1okdmGLZcC1onSe/0DJyo4
1AupCKaxaRZHBjKLyxRzLfNo92riJMHPXbUNnRkc6MxKPv95jjfoK1dHxtuh
zv4hnq93n+oNyIUZo1PapaGW0HvtRQo8EANoQyTjNOs7rTbe3tdapsaZFU25
dk0dm5K3OCAlb3p5ZI/NCAsn2cgbrPyolY8Wwxio43ZsMs4ZE9dm90LF/LP7
D3V4NGjeXpac+2RC9WvR5PCxzbABGs2ytcgkSPy7jJ2kQvwBqlSlKh4wKgl1
rGKPcvWQvGaaq58vIEDhnG48etoPtSPi08g8NbzrBdX9d6TkHtTnC52XgVqm
8cz6vnXD+xJuV6uf0sY5Ooc20bQ1I2JihKSJVg6rEX8YqGpFF3u3EPUEX9UY
5QFmS6PdCKjNwECL1X5mxdV6wo7JpOQL4CcrBjqtJRwYpWZmZYTpWTy6E5o9
agFHXMLT/rp1c+SdpQy+JjfjGfLNgyfm+HiDpLtisfZlHFpAqoTjfIWUhKUS
RAGkrh/wE0Ya+uBtekq7Hst6fn47mRosXNgHcNaLConG9owDaSqQGIGMz/zd
xDTOaHBPHZGBHhR6Ut64NXi62DVXFiZxPCUt5KqVolZ248LY3IHBlAMU7DHJ
/Wj03p9p23otniu+U0e/hhlx80KECjApEZyy/5GLEG0fLLNEJjuCQA/jqxKC
csurmrSpAI5eIK7JuL2PzMAu0641Jv8QCY7SdJfRmn7KxZcxbSd5iS7MIQ4F
fr/n/BnCAflArKuPUodeT/R78+erQrQfXDBJA2cMKWPc3TYLUNdUAAhreeXC
fdq7Nx0KYYoRvlH0TiKN4Dy91rQ0WKVDRNcAZGkui+1jGaYaS9tuLxFo4dcM
Iei8Gg0W1yTzcqIWGMfLin1m0Vu+iViDE0Gkg2nRt1VM44MYN5hGxcBFDymZ
HZbmJRPLguhqYQoHVGAAvYe4eMGs68XG82GAKOPHuqjBors2cKnYdo+LGTCK
PY4qdedbgzQb6VNZtv9WTkkEi7RSq+eIBDu495mccE5bkrbEo15QXMTJG3Ok
D59YT/kFbcLerLzLyn9R/w4BpZHCBPZjjoTU+gZFETPBnq3INbsYP/RPVqnE
qWuyKGqahhBqK8ez7Kmufs1Tnfw4cs+2bxFeO3P/O88BfJubulbKiHKBa2F+
A2krA9ExtuODTfGevlqIoJEIP5ZiPKhTy5/VrderQf0gA6HClmMCyjYFErWa
O4LftvDHDvDT3r3qMIwy/se/xanfcq10EG7sQspIOR2e3rm3+2VS1peQ21I9
irwq2i5a23NYeTBKk1D9ICGqRraNDQOcqwPjwEOtCZaBcrkyFx9Esm5km3Yc
SQHf74CE73l2JDjGtLnhzY8PRyG9da/MKNqqtBRj7O1fep9Q0DbL6CXXCn4v
NJKyMrEe12d9BvngDtDji9d/56kFkec/ZZW/EKu82KyLzZfRr3QMyn/cmAqg
pec8oPWTLoegq5nNJoK4cEhujdtSN/M6Qtv8Ul5XeHvts/Nrv1euEf36R8db
8RGwWWoSJW1JyYoQK4ndzzK58VYBuzv0et/MLYw/kvBTZRRWS+K++msVmT7O
MFWj68ClPcN7vJ2rHjQOuYBfV32rVBbPYDDx3P11MGgaZnP5CLdGMqrw5GQI
FvtyoXM5K6CP/5qdy3dXFWlWXXZQYTDoan2TSYeCTgkKR0tJARMZJm5qIUdB
Y6Q8gxYuJ6gKGV/9sqWmvCMbjTu9Kel5EPbMpUeCz/fQ2LEf9H2s73c6vma2
UYPAv5pWirp+G+W3wb6VyrXWBWdiHVSSKdC3naMWR1V1zVC9yNUUYY49UkEw
rRecq7ve/VpaFI4R1m9oMmXZ1Nw6nqUFVvPciIdtkA8VJJnLCn1sy71VrCMP
0TpTnXPiT8hPC+XJI15PGDzhyCDvqxUjhk2lGDiZCrMMMHJke/Zpj9fNmKKf
N2CjC2m4yG0QpkUe8RM/mkEw3Zuz3FU4CksVXNbk72XMtS0K+4870bIYLW6O
jRN0oapbxfkym+pa8BW0pZ3tAu7xRWpBryOxR2Jh9EUisRCDrvTgaeCw8Coi
OePeyebV50bSJ4BquhmmkeABBouH54Nvpwyxwt7Im/uMcmYobYkMNSDi8c3b
Gvr++axxrCtLr33aH654Jm3AsG2ukbjzaYsUuI3mmzSVfZhb8Z3QBkCJL+iK
cdZbwYHp0pgkuG5O0w5yLLAuebo7MATiFLITgm0uw6rE8QdMOepr5QL17RTb
G5SnUkBTFkc88Eqm/kQd0uMHTgcy4zNR3/U1Y2Kokg+cHY+jvmoAaW/7n9GB
XyESh7KF9VELS5+P+NxeOdyml2/PX+THoccMuV2loMs7nfCCvMMXLb3s2AcN
tuDnKXOhCIyOmxsccgcVmJSxIbo4gJJg8Ldk/se7gGEwrWcKz13+By5QNpSG
yeL/gjB6ChgDYG4m7uLhGkMQSyDVrveB9Q84J5sW1b9rtFnFYjR++av+czJI
8xWE0BfbtWfUwiflMxYIFBAw3v1oZm5r5d29wGjyyE8cdMTLCI896iUl0oBQ
s7B0D2X5rulA2n/iUQb61KgbiDUUeVcv5ASG2TZww4e28jTO4/KLHGUGvjF9
98Vu6yKSQyQqVxGZWcXXVXmJDUQh0JT4n6EsHy7TF1n2Hnbw4V/vUmQjHGv9
gH1HWPmnEOT1yv43tt2q5Z8K78wpqMR2kFN59G6zFErgzFIRKO6XcXUbjVNX
m1Hyx3nf39BHPI7mD+3Ej6NmqbPvK9zA0EKHdV8bFRvPA/dGlOzKIh3Q+W/q
fDvknoM/KKX4RvxO2P+i0bdGD9XMyy9JeR8Q3uZ/oMYIEuxKEd/a2yuDT4pg
bel7mqT1z7G+AU/QwBWz1q8V3wsObBnJr+19nEq/g7znDUKwcc4tE2JPfbQT
2LqsFUmcqIJx9GLKaRfWUH9Wh1U3VDTSIsH7u4kU39+jmtDdpTH5LzWHy6x8
15WIeBB2S0be/5mT0OcReePt2z0xX4/gJ2uCgxUzF9JJgpBCmlVtlqiHyEdk
nJKxlxi+uECf6oX+8oS+YWs2m/QCoMUKidYDrZWQnt8I+ef/FHBoX30ZMJAW
yLbumRQeI50speIv01Pg5u9IiDBu+DiKGdNv2LhNms1HJbQuDijAuBYYEN88
2Q0+mbTW5NgaQ/NBxc2Ze1xh9XlqELsqSo00d3vksetpoIOMwHQFFRoyO3+U
ul9/jrfSwDu1Ey0V5Irlnk3uwMZKfPe111d7hVLouD8lhVD8Fn5w/adEQGzI
8aAtjWbZloeo0mwZh/U902/MXhwnMoZqgm1WVDy6K5xlDsa5e/DH3PJ5AK8+
xpuy7E2FsuBa0q+EKkf+R8Qn2tzKKLaQjWhJuBO1N2A1lbl6n7r5yA19g9Qo
myUWfvncLi8ZZ6CS9BE55KYw+xJRN+thyUYDrC6cG7DTshPtrUlaOceLHAS9
+8bbIb/iKs/NrXUn/aAes4Uxgbo63xL8BTxFSsNic5GckCyTmPHa6FKLBDD8
qlOjVTNIUN0hdJUvzdu7skGb7kIOuFLpcWnOqUAySS1f95fEoDMyX6+kaixS
+HUT8Cf8tpfxIkS8s1rC/YL/a1fH4clQ0vEWcMLV+8tzwB3ox975eMfrfKvp
FD/ylENfMumPJbmY7jIYFr/dFBNSzy1LeBujreHFaqy/U1JgXIf6BDGVyUbH
Da7mbzolSHnoE+XZRYEwcQTHfZxW7Topq3/sdLsrxEB0Llr4nXd+XdMRvMrL
FhcJt3oPfYBX/DLLAmuxnkwdG3PrfH/ZMQI5J1D3ag60ndj0lwUxpndS6Ss0
z4gQBd/6mn11wegUqP+6NklmQ0T5WvgtmwApVzlP2u13EVZZqoF9L1FGbcpG
qV6tz61SqU83bWmgE94mZ0s5SbVDkXD30pfymI2UQS5/cWF0fx245FTIDAjS
400DSe5DC4KwEenRhHc50DhNhfwkFZ10PUyoZZKEmECVcysQZHGNyNyo0/lX
N+wvZ1mAm6I4L+qW1mhijIWV9cHlFjUsYNhRhX0+iHbXwnfcmOIXN93mvCbw
lBOtOSF8ADZAa2EB+va3hsJsFUJCy/pK6Dj1QOQugkRA2dRpsOrIaxjBDtrA
Q3dBH8D40C+OwhW3+aleIOhOg6jzHCw4kYox/ZBcNdkMpVP2Jx2DY+0Ty1CZ
U3hlhTcnGL/GQlOlYzX3NgHcWHB2vJUT6oHij0WIhsKihl1HVQ4kBj5FFgcb
afY7av3rV7B1rmPr/Qk24QDoypcmbokhTGljPH5q3efpi722NkXaOaNTMHHB
pfJK5h6DToUo0HTtqZVpqq1coWHnWsqJG21Q+QFbgkxy7rb8EchH2j9YU5TQ
XjTJ+qXDM8C/a2uRLQjKTzG8KgabPj1ajQGZ5B2AoB0rsUc05EwhXaExIRJ4
V2tgXqgbO5WrTo+fSeYgRKq2lO4zD0MXtxDm40H0yiJp9Rdbv+2m/iVzdlOo
n9YrVUdtPxnq8k7sh0KHPKS/m5uYmCH/8GTsprTBMq+WQqn7ytq7sIfNXLSi
Cikl59xtP6U10ZPf+qgNr42BbXt4fx9+Mr6k2/d+CXkiw/udbsGad6m3H5XQ
w8ycVgL4qvnfuIUHKLpcjUE6lt5fkPVVYdl4fCGsDTCjpr3VVMDBqPO+zIdQ
RLToPYYCd4Bjd0E+1BqI4joRpJnY5n14aZ6VIlmN0awva2j5RmEPf7bx8SlX
ZV54ucIFJ7NAiVgui/WM6GDYyD7WKxMV4xXl/lGi1W3mUwZo79zZ679nIiUj
uvvwWYxBY1WDozxigbcminaC8hU1CX6w2TLsJIeXPduOcFKXsFgej4U7ZHN8
1gvW2y0FhZJkDDQGfcnYesozAVcKaBmJVbanIvwQ1q2dGGSeG0iV6+dk3myi
bhzhxPPgWeVJxvA4wIkVMgV32QDC+8Cxa1j2q7LwMh41OyEGsKmGXKGGvHpI
rY/48Tp1OdrhD+/K8Umm5F3LScmgpSnmly3tDboQXNo91ACjGeOeDH1wTvDU
IM4O8+prboYhvHIuLxD0M6MPrzEHtBh5K+Pp3wcWqOnDE3HrsABnK9N5Va7r
NGUP0CcFPSTUT1ICUHhbBRz/y98CURbgEhVCZX1r0uswNGB2LanW9zAbogUs
DWmxigk6J434PDhY2ZZX3cfwPHs/w0hcql/gwqvZk2/2NmFvWGqvwPGCeecz
sfciAVOWO78U+CaNY1JDDk73gfH/ojBVvBbH3pHIEcHRT/n026DwKUEMgkc9
Vt4ZHJGGg8KvN1dqZcOXMcuNxEs/SDR6OPRjSDfFhEn+f23FJtE6UnVsqgN/
ZQOSLKT179OhwEBbQBXRH0Id0rLN98BczlSWQ3twx2jhqTcQrlZ+CqgeCLe6
I6glNmXK1d1iIwdPTGldFr83LvoDhnVhYM8/maEVjFY+ZaHgdO/rnsA6RIMw
XBu3V4MIeRzLopF9918biNzfABe0VUspIhb0fnwM1IvkJK1UzgvsOw2AKZ7N
6CUYPGZgbITkUIXeUNfr9bZxp5oeCA87BYgCpAx+FvwxtZBoudHsE6MBsbUq
X0D8cIDHt1nIE9WnXGqj/DbSagDfCmQmljmySrkLHweslXQyLWwmVZzjHjyC
xvZepBvgi8IqEYvLbU8CCGaVXsTGEOgLoHq/GccSTDfCLU0ELXq5djvIr5bb
ipxEtfWMIQrfCOcWP9zrIvYyWbrhxJwMqXrMjMvC2tYjeA729iwVaExtSKhB
2UNp0QCw8eBU1SgaE3yK14qoPU3WyKZU7yzxhRV4QwhNLYxN5YWaqWGlD1Ex
0fSNKGtl/SuWn3jmwEGrScXceEh1slNoWBG7MWC5uzU+59KxK2709dAlbKPw
ibaDuwFoUh/HbC/CZc32AvPzTfs0O/rM/CMYWcD6CemfhSItOo/LAlF28EMJ
lQZk3uRT3cEN5oXPymoQWRVALWLj8QvowBDQAg3K6Njp/KQSuIDc/es9J9mh
/lNitrW/VhMQzHN8VO5NSf22jjYxwhCKSZi/leOAgY84kbHHcuahRFHhBAaZ
hLlyixpkzgZszW4fgov1n/QUOyVsFEQsnxXOR9rWWh6h4YIEN5GNNozAKK/2
woAMx3PIJHBW59/ees8C7j8CHJwRTru9jEtzqHA0fBazSRnvL6oAhc9hOv+N
my/d/F/AVGGjiD1oMGGAahkGa8wo86VK7ivqZzAAWBNuz6Fs5bon9BOZ3NiX
0Vm0E53uE99wZ1F0ymGWcNB0HrtufEep8qoRwplu7zywU4+1SdeGR6JYCFOg
1/wipQgkFaZSszfYpLYiS02lgPDm7l0OyK+kAF6OtS8SwxEXLdOEwFVkZHed
EchUyyTBFzAPKa693knwE53U+owHTTDpNp6tUzWkkgSGZSoo510rx4Wxi0N4
dSjeNMWPek+H1kMDh7r63LKXAB4sCdRm3BiJvbhyL77vlBOlNo3Ib70cerWj
LezwPjoS+foib2ySslgj0nvD1hizEy+06U+6M5lprDFlBEmeMIfSFEetiSaX
JF1+nfumGC0yZtSQyGi9THAbKO8J//VmpZcdUDrQEERhJz5vjuAz8/Z3jYJJ
zUOIsSVUb8AzyVvMfmB6Ey4piQgw2NPID5735MGud8f/ZVh9SRGCIhUsWIhl
HFkAw5TFJZVipzviy0I+k2aZu7nnhQPHK0vL5mV7xd9WREmRarHzQTsHnXK2
VWksko0BtbyhdUbqOrFXY0CXLrxUmad7YragihgTs3fajktaNyMZCDD80MZa
f7qdTT3Z2LYlStDAlfNVz4afd5P7GUBhOKKBl8dREsbl4Hh1XOdMTPNE9rDo
cGNy14Ces5dCyDBc7TTEO8kFiY1Z73vJjTqonAT2erD5C+mzHH7kq5j9jT9S
r6Q6JaiA6YMhKQ2Hsz0LhWyDUfSlzWYHFl1DSXBPsJ1KggG1liGDah6qUYSY
35C//RCMTOiIduPhMkexRM8cQUYoVSSgMcmUp8OKSnGNUVHHjfSUqc3F8n69
UmQEtl1kNS2p+mhiVaeQEOke/2yUXnb5U2+xxJ3hL3lKmyGMG/FSm3rxmvRf
lw4HE7haZ1K1P+/PN2BIWn+Ot3WqCjLBsLZC6e9adSvYGykXVd0KUkpnr7Tt
K32s9ol4Kgis4cn+04tPu0aLfsj9u/VDwCuvpJHOhWsZmmk2Kik7m8KmO4NN
cu3Ba19vSm3ONl96cN8MH206x7mebDldyqbhw6Rp9Bk+JcNo/PyZnE9qnIQp
M/JSjQaibKvQxDJfsMpPMUgTVe0+5ydVzJQgEN1abHat6a6yyIPvFIKP00cD
KD7/GMFpFQ7LKS1meg52i4YVj5ZiR7l/BPz9CpMNAaRg5xLnrS7js8sIhlpV
yNn0aG5posrocvhdB7nM1hpeW00zPzyRe0IGmhMX1QkZjAm3woO079kswj9U
qSVXnKNZR/93wX36SUev2CPILfDmJO3qDvMIJSJxHsjYwzTfGddApTDseuSm
l8giFuCPBmrzLLN4reCNrC4m75WqngghlSe1oVl0D6upTRx9jhukIyJcVOA/
JDv15CagK8y0XGEdff6cMdmaX4rS10LrdmyPBd+W47zaBPztkzVhzsSwMyfT
3r8ujCfzW7z3naRwg+tTVfEUsAu37W6AI9rG/3h9v5sNtbXndy0SYG4PbZ3T
lRxDX6dmfMWXx2QpxmFE1702LUxQtG+GO2uOutI7etdiR6Ctt3fVWgX3bY74
CnbXvzmH0gGsXoNk3NHTE3UZkKCLUh2WZHup3dmimwchKENq6G7J1AF7am8J
Ac1K7QFo5juAlZSzsT7znrOMAmyAdZu3L5rpOPUxwQ+mHJknVKlDPY4IiY+h
y9Uca0UyK2wc8BEni2whIzmJEKC4bgkp2F6QN/ufTLrBoFVruyyvFQdlRNbi
bfE/g9tqiELsElQ1lqSZSG8+oRxqBRZgcjgTbo1VO3EEptmPqp+VZBXUxCum
sHKQqEPJv3+8E6BqpeZ+H39Ft8rBYY++Kf4XKPvvLdIC9q2n/+cO6e6jRL+3
i7AvivngNzZQcHmFEuEWx6cmJt7NBFZNQRUqPZyzFeJoybPWHrs146scV2NH
zqyFuMqxUwxBl7f4LH+N7HCnyf66KgXd5IiFMlRpfl3SEJAfyiiCnmxITq0v
dp0s3tcQ7P/KJBMC29iQTFERY7c+swT1q8S6oEm0mNU=

`pragma protect end_protected
