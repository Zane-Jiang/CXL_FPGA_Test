// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
r3hpJDlAlWPuiHXuc76TidJovk30y8+z++b2VBBb4onNg9fvTDEeUh6uZYjo
bNtq/51HKzfRlMozXhRatXOGIFCck7a8jdjRvvtTDMpKwAGWSM+/z0ER0NuT
KFnedUijaXMTaXzpJEGdzyabmXuw0uhfe/lIJj+MtRo8rP/OrCAL25OYnf4t
02KvCCsSFfn+zOVG70RQn8MYYJRiDI/741m8g+G+mT60T+819kFYHfxKE/ql
s0bLVh0wqg5uErgn/2xjQ6oLIsqv3GzIPsp6Zsk2ZnPG8ghdRgrrZTtNJktC
qxPhwhkyfRaEfLMZGNIukZlSQ9Iw+WYTXCEj2sz0Cg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
akXnlBV2hvOXW1R3PIcWVWkdvZpSpYOn8OPnzFhRX7sxHRTwAOrlFd1MvNT5
4VLyWZOAxPoCgIm+hyp2mfKE9gSdVMSvoGnBSjOXnfoWBmi00CAVPbOJYl04
JRjs1WDeSwApFxN0/KbkrzcNKDbiXZaf+32ZnTIdJuhRm863HEHaZOxeVPJQ
rnk6OpC7f87VgOG2E0/G+mv73SszXzuqHfdj8XNYDTAy/xIYAe43McRt0C5m
1iMFs0CVyXAq0LR5kRGVYTh1JLcjqSMTcclpfSr6ePUCboVHNIpnpQJcXvwZ
sdh7M5XfsLnHnQRBBzpTaPJ2WFvnCpcO+jH8CFXlkg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HIN3+IieJ5imTQ5UuDh2jp0cA7/HYR6/lmWcC3r4KGDNlWiDGa6eDm/GrB8e
42DbiCt6raqhvBe+/k8uuUVlGtF+W0EFXLZCg7WrEXGIWu7PVyMw9AtCtEnc
TCJPnn8G10+RAYJylnyQZzOqcmb+bMT6lKNtdVC4VnS9oOZsj8euOwBPUCrM
V+/4NxYFQDNraX5yXHhFpYhvKEmheGcIMIqB+sswZxayATAp8Ai6/etEgycT
uiFeQXDHhraVUaQ9fRBr2bZath2yQ+9VrnXiI4wdYpeJEVZzqPNZhNCZHZoq
LE3tnUP8dWqbDfOE58+kL3YYO+aoFprr6fuOGO8mTQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MDBi2n8xh+bo4HE6yVXXc1Rr6r6rHxRlobPzxl9RhrUUoclwYbqiLvjM7PU+
du68J+ifigCP5rrcw6xwWEjQYYIzYOFeyOZJKn+Qc2riYtBHJDp/TC6U5YQO
RK4WcqSaYZTK1U3OXBeMLXonycUiY489yUrg2UtLbpdgHyPxbD0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JeoNRj+uw0x+13YgVD3bpFN/IqBmA1U3Q327xOBEBjK7FXRTwxWLv2YG+wML
U6xm1DmMQl2QgRBCYW1hPvlFK4ewcOOpBf1zotH1YViM2IFfmOzbkYcBkzTl
zL/CJB5f/AnBgDMhMaEOmX0p42ltOQuyB4xBCMJB6AarC6LrO0o/Y/AGR0SH
ORVSnLgtBjMXapiwmvCFgJWxHV70Jqu2ol+ALkQELsoFaTVMae+8Cz49MpMK
ycqB+lS06xqUDc/hL7RKwzsIsuwizhh2cFQxCsYOjudxFWvLou2nwy3p9wpP
InklDH9dJDfNTSNQqNeiI8+40KwgiinUJMhCYYiOC5VTNabVqChLI2UlqOhP
tz5saITbdgJOrGrstwBBiuIMpFA80ulywIw+mo3H0XYxBPOQeHYz6gxYNgxp
LbinO3xZilX2koC/s8oYGoEtSQ8F4ljZFFwTxC/GL2CQXMHSl8/9ByQRlJrY
JNzhJc/Z7+87cYbe8JNZH0gzrq7mnjPT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qC2qTbvlIPsM1KOCiN9qHhFfqpHpZOjdByblXrEAvj/svqrK1lysesglq39f
yruFeb2BirL5L5djtKmQMku9Znb+gKzp9uuFjS9QCVvP4Y1PnrsW3rl+HvVF
b1qkaMIVhtfsTX9WR/O4ei0/f9AbEZXuwkYkpYW881uGdfSuCY0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WCgI6u60IoG3CEnWp+cYTIjREs4tZDWFKM7a4uxAxWy4OeFjGs0MsCwfMHp7
0NCMYovAMQhcuGooucptQNq098XfO8TvvLn1W5ux2zgxK/X3Xd3i7FxXvR9E
G/iqKUw22j5Sr7ppIttKptCftNyORdIsEMYLY8gVM3gpH++9abk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
U4ngr2qBNXH48MJO8f9aslMvMU+7yPUfrB0ioTPCvRQGhAvIrxGIT2gvKQqA
UOwue+5Cv+V8UEUWuAPxigzsXuFnvhhfLBfHljkT6TPMJ3GJK1CeV7zE888D
TSTLo3Ib6R5D2IF6RFw8EMpgcY5Ygh+NtAeKIPJo1yFJR7+83qB7YENeD/rx
J5490yC2aEkF6t3LRzaWt2eIfCcQ5JmtfNSaVaPk+T+Qh16sOCS36MoY8d3Y
AC+DflsCYJEsw999tfc+e6vhPBQw6nvv7ORSmysZgKHYhj+fN7roEgjaXSNY
46cWdHxndi+4G3syOYxG9XWUHeiv1ONOfwQcNfl2tL6MB3/es6CNOXHiFpxh
aNlI4lHstvYUaObkp0OhJbnMVlDCgEdN+S3HR3Pk0++k7KMPnowDUOpyJQOH
lOOUgqZQNTYpoiQglrCohbvDbPQ8xiR3tNzOKTXhOQ9W+aXi91l2cQfQWGSD
njeOGlP/U/X3h9oWi+C623bPbfXd9n7YsU62oe6iMJ6UEcKeIxndRrYkqF7B
SrtL8teAYFBmmvADa/HAveZYsoyk7Zm305LXn02QXCBnzkZh5nq4ZP7T5fCp
VT01dRJ5I3n1yE2Sb79MY/NJRqfw48cMwUvR87pfD/ctWb/29yNdNCN2eyAJ
GqyltCPR6trv/6CnclZKDlnj5VmlMcfB4Gjvu3lRtLAc4Dvp6axT1xg3387o
/wq8FEQ8+NrHHjI7agURST5MvGJXREjNOuUAmUtOSjWU+9onzA2TD+Bgn98B
BrnVkXZHTsfIwzsdS/oayqDkcxNM+Ogg8a1pSCc/BDk0ZOZZURqnwbMnxYFl
FY8Wa3h88R8G5/olC6fIvYJctFa2Qi1ywXwixl+pAhP1wzPdU0ymmMXHCCkm
HntoWoNeAj2q7lOtSes/7MDi0kiNBZ3xbMzij+dg9v09iFtnqaoVYaii6nGu
SKTp03nMInjZ6rnJkD9l1YhjUws1ULlrYqn4CxNhV2bAUHm9k0XdS47uShWY
QzQdviun2sdINEq63YltUZCqZOADNTn8qbmADTI8INGzcyuvZgZRrK9Kvk7f
78udU9VhETke1VrFRUsWlHaFbWfnoHNGeoHdrmz9W5GtYLLC7AGGCCTTmXlB
cttR9pzRNWq3jWi5/pGrmlTRp5lot+m/+fdzUcQrxmDOS+DqKaf76S+vMGBG
OJGoA1b/VtUzM6nSnsVDgP6HozBKD0zhnm3cGXK+nDfGdPnp2kG7sqGG+Nfm
fK55DZ1rFU6AEvy7uhToRmzwVQReVGmZy8zosjkVYmYO6k0LyL/653W1KqNO
jGIW92M2eHJbkjL8/+nrwp3iUJDeqcgCcB7xv+tHjUTqqt+O/KLlBWvBhsCe
Eb0YAl8=

`pragma protect end_protected
