// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
AOnNOSOLg/k7KWG7RxQVc7bs2tmVJ2Rg7boSEkzhFjtwVfr/7rKAkfwMv31ub/Z6
ca5DM4p6hS9mqN0fY5xwAfnwV2G25DZ9ANNxwH7P2Ahlp2NdFogjVTXGF0sVoHUU
PIR4gXGjN4kqJrPTMhpUhOsHptc637VeAhvEU6VNqdw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 24128 )
`pragma protect data_block
reQfKt113UIBZ49vaghdBo1fbpFYMkudzrtxeTXUWa73i1Np5jb8LJCba2ziQS+t
QCj2E75ebSNPUBtk7jtPeomwYOxrEouUVQCZh2bhuEnOTtpXU5CLALLV45183V6l
CGQV0QjWZs99aERW7JD6k1uIRtXpjru24PNgA8T//yUdDt4ZnJZPGlpCX+bKhEM8
wCYnm3AwQGHlLRFGVcP0c3JfWpcCKdjSjRyBx/kJsMzd4kn059zNPU02LGop2skj
bOIezZKN6pbaWSwp5NcmagDy16e8jDIhcCHrqB8g0vUnZfktilxdSZok+n/itD6d
j11ugLe/lGK5bXWkHTIrwuo/91/VFdCWac++xTglWxOFSJkkk/vfhnnbA0VCbh3/
vgX0MFnx9gdvcpG8ql6MWlGYhB/I7HkBrBLVpY5lS3z/53aJNzmzu1gamFiTEvqD
3/BQ4I5zBMsxA1mqYuQfVDuqJzvAOE9vi9xg29zDGGoTi4ktvnrrgWoODlEpUczc
DF1daQEbbHIqnZZ3KAn+tlpgtbTGJ7lYF9x69XCKGCS67a6hW0DUytiDySxBt3MH
I65OfcUVMXMVjYwTqhRrtEMv7Ig8Wp6w+K0i5ycA4cXjKe2vPuCI9PQ5wYozI4pw
tsV+e4rhLlNTlDx7Hwy4c73IxxZQTqF27XcK3J0ROkRKik5Vjd99U9jaQgbdbs//
rff7EI3h8L4yagVz98gKnND69I/xAkYaefoTq3v7h5V/RCaosC3BcxO1z4hO1wON
y/3hGH/e23LYQv1m6PP4LE5Mxps9AgdFbQ3Fk4e0DRrHcqR33V4ZGnz75siuLkWA
TnCrNvrB/v5sl7ooRRcgqzlLls8YCnzl5myGXOX+FN6Djnc4EdZTcrD1/JA8aO39
QIggGgjdVgpUh+zO7PySRDNrWhsiuv+BGu6KOfOlHeZjHKV6jUtQjiW7Qkd4J21O
CNKWYT5pIsUbbS7f4mlh6QJVqBuLE1YONSXmZMNeFwEehZPdaDY90V2ESBFf+5g1
Qv/MDnvMLgNGWEb8+GVcfwW1pLW4ONzgW/i2ESRJlwbIrFK87qJG7bi+d3Y8qqQW
voT5DqASgmiz5+cl6TRs5xje4K/nveKxtF09n4QDg3YC7SB9UuVLkfvcQXrbsLBC
UT+UuHgxjGoG1cfXBRTgMOAZSBUTAgwrqXFxtvOEN+oLncPmomJCeeETg1gXYWAl
VsDVo6l0efUT6khj1kFwWNfKETwsqCseB5Khk2dW8sr249PgqpX49gjK4geR2ybd
Eoo5RRnNmK0EupoB2Umdf+F7LUe8HjzFOxZMJVlW+n78ReYNzIFQsMV16UdwRxau
5MggCrwSK8Z1Ve2S7mPjdV3RDyWCoqwnwHIDciQn0RZ5onkDsYuJgtW4IHS4ST5n
5ISoufKSQVa8ZjIz6jMWiuCviGQe5jb0wtxsFDbSoZMi+Nf5IXug/mJLWctYqMRk
iBaZm7RKY9KIJLVZKov9X+Go6SYk2M5ss0MJhacqnA5i/lOcwvvbP7ue7SpMJGRF
1Bs3aoP/Gfq7ddsXGbS63PQJOr9cPj1OiivEv/oxxVoTItRFX+9atnvmlm42aab1
GBjQ74tSPipwMf2eMKQPo5C1bP5lGMkqRmWw2J7tfmU5VmG4wXVCkdNxHEZGmLPw
IvH4KqwS6duNSB0v369DcEzxMNCJnr9xOFeg+b19Jv5Zfh9ZLggwk4/g1e0fFA0W
keE42mhs7qrtpnrs28VJ9dpmjUr8Gwvic6oDk7Sy2iMhPCIpL7teKLJuKv/dGIe2
bT3ukaGFB4BqNNtJCmXey7QfwlGzU8Ahovazi7dD9kxXRQn5iHzUJBko8wd8bZ/g
8HMTrFRPsMzBkBiCnnbSK+OFt7gaxceK93lANf4yawyVhhB9l/ie/Pr5zST2L0IX
xGfnl9ZsiqWwEwXeok4bDc3pskhQukFmAKOnornVv3KK8tgGcMJY0ZAELGSxj4dj
Egsa2fg7m2lsem4NRXaQgFdRjw5WcsJD/2WQaVuOJUSgmBP4EId0bZoCDEgg1rMP
cHaDK96qwFeb4uWLSbs68PVUaUHkfk7wV8Ku8RvjOaW3LIEaDhgvuj3DgjGkMzjB
/F0Z8Q6Py4GIrduUvWzT4jl/ywLRWZ4dHmSyC5j0Iur3RcPZ460xats27DHoEHdt
tp6zDvjrInZ+EZ8DbjX5CkxkD/NNe5sfn3mWkviOH3loHsFp3n/nef2h2WMz4/0w
pLYO9HkKQ04dnwOa7yecTH7bcf7m8Jhk08+MJ4+sVkvMY/TMFQN/+76vhyBC8lrV
z1CiVknRiO3MjfxR8/RZQmcEQRhetrquTa/TjusD9w6NIycXGEa9/I03ge0J+uvg
4nc9SGAhK48ByluLhNlnEIGLo3nqds50eKn5NdlAWvDJTEI+oqSZSgFC6JFokyCV
jO+v9YfMJlHMX2LbfC8bl2kFZ3BYGMETI8D7WNc5TzdPsFPLqsnIRI238BKGA7fh
Iyp8NqnLPsd5nKxCP5sNtUdyDvoIDatU5Phux5JV8CQU5vgkOE1dJ2Poio/2cEX1
witrbu8djgAf1QOs4UAKRrQG2zoezl4rUmaIrtJWhdsJm8Z4XoUhAQCOfRqc0vcK
yYWWo/4wp+cN68nhrjid9gUJzSCtn5KO2hh6LoVx/olf9vqfiilhrqxExlF2mhS8
9Jer0ID9hJzfnYq5lrC4B5n39bFF8n8O/FaXrMrfG5yE87vJOXMpxWe6Quvt/cHz
MbsuH9wOahd6uIdVbac4xJh51C23mCHZRfdmsfxa3otb1gbRDPntuZW+n5jnpxK7
0ELm4EnIkbREdgYdf5zkGjlBzw07L0PRhVznOJIsBWXrL237zkyNOOCy6aD1se1X
+fHgtJ2dJc/ZhIGtcbma/FsR9O9+e4vbzXLHU8ic/XrPrmEjjXaCjicxub7dSTD2
C+weUHNwFMzi0oJzsCDN4nWIsGenyUn0L1fWPJv3DJ720dv7waUT+t1yRS/x++hM
9z3EiAknk2UkQ/ZtkJQ6kuh6bRW9FqJgScYqwjo5hi55eFkTZ77AxCy0tbc9bzgb
6uRUaO8BqZJqWyX7ZMJw42erDGAuk3a7LpkUKF1lUnMlK9tJFqCvPH79W2uCDJbe
jjrgStuZwTZF6s0vVnFmeu7Q9hnHmfpiRvCSypHIbG0hGjDFr8q/aWDfPM1jL71P
y5Z3h2Lbqr8DkjrRGcnZvotZDQQmT5Lh7jGaY06EXNTrNiIbhOnDbgcBRew1PzTO
v9B74hHWal0y6Rcb/BvMfpBwx+nd2M3XbEaY0ae29+YLLK+AyxINJ0ANXRAukm3Y
r8VtDjuPElonRyT4nDC1e8i5ikWthPV/XbEKpqZaQIjgsxCwfxzbcFKY8kMHGLxD
pTDJruHFl1Fx7FRAJJIaEsog3qaFDC4ND7n7LWuS7p5/NYpYVjsiHPlZaKrAcUTF
UxH2oGFWtH1dLpzDQNZWwXNyF/q+juT9qcfwYTiWLjJiToZoXUDYIVWDqgCxyXvv
Wv/k6AFVXDYWgeVgpWv3S/MPIjKl/TfKNboOBZ8Zm7mznoQkRwh53bNwWXdRITVV
uCZclD0hzmUQhx/xAzWdhrfcwOt37nyW5QExU6sXdmEvjQg+JoxAMoItOABIwI5z
7/EkXn9QhMH7dMwzlTXLIK9U9Vsj8TJ+o4Dcgf5L3HDBnX3ZkMUVc8+l9yRlPpy6
HMmVguWqTGgkW93x+W7hvQdpX8UqwUbtOph6z3ruh5OlfFxCaFi80RUMLmh4ly8H
2lsfys9akdViHIUf63IEaoWctKr3rlNz9UiqR9YZIFxX30sZDAzAtPFLiTnJTUdy
arsaSpnjN4kosGwokLKp3wCW6zy7wplJASSKBCnJO5nPMgY404lfbKeLIKcwPZyW
5PvvfNiOuiCCabZDM2ph+TIuaIOEhk2Tstkf0EBMWJFh+ZlavRZKZC67600i3Rfe
WhJ8z7XbeUBWcemhxLqLnJGxAVaKPFi/Q/M8SC5ZhQoGd5CFG2tG8E7KiN5ply2o
Fm1SHpoR6RbZobS6TOtj9vVRAV2oMns7aCjTZYpMsvJFBXE5np7pLuy/qLBw/mWA
1CyeOq+FO9PMrGD0WgB55hWo+XSyb4H16LNK0NxlL4gW4TiUSvd9oTFTQJdceV3+
wY8V4BAF451OEcUsP/IMqjdvcIBr8XAD8IkdjNRunVO6vaPEV9ofd4lkgzsVM4nM
Oa4hUFOOPUPXGM8wYWqBFd9A5mZIwDYFQaCDyvP/UWVdaNNEb2vo3Ow6ustNqld6
LLXT1RI+sRjT2jm4vMaznK4r/xcfrspl087uujlorAh2q+oyRu0LU4mZ+V4GIw7n
tmXxHuJrvnF1Mngog6lnxODA3K+zfkaHQJS4qaOdtY0v8qODaNpYbaQKL75x7Tmj
H7aXT/v5VPioBAUNMAXjsiE3PVfWmz8Fx9HeItj0sxmWS0p28+O9hOhYSaJFEzk4
V6ZUk3I4Tc+tzQUr74POBHB6+dSmLEDoD/0PmgnDvYmbZjHymeXnz0CwR0wgTTP0
7pJ60ea9Kt3h2tYS0k6MKfa2oqwBh66cE6mOfqp5sAYk0q/nEk9xjZxXskwwoB5W
hKAfk3kjacqR0UYZ8f6Nwp0uC5jmBrzHO5C50DkrkVcMqUdCqaScELNF/FHIx2Fa
gXG0hvWCZoCYsoJJgMPYN+o1+Z0dTcP/MMRqtTaWPlePKui0IBWpGUWIQG7zTjI4
UM982RRE4ILFkZGrQQNBKDKolO3oqTdxGxBhUNHztoa/oq0BisNd7p2IIIAD9M7O
KWjMWFQaRxE/AD20M5Pc74P+cmQun7BqXpmus9RuIG+48foVlIaRQvHzD3lr9OyA
nZ6jb2qE0cFRZX4H/K4t9num9NaH7w9azkYMHg36eRkMrXhNpZVRIigrvkUPjP5+
+HisHIPlYgxcXYqE+w6H1epCaF/tht8I9TelG5nD0ApENE3KGrQ4uP1W8j43VEGz
SIkl3wB73h8uvqxyuaaBL0mFzzLGJqE/P3IIj2d0sRQB0AmO2YvO7uayEGBRmFaT
q168/rpeTIWVDt8Ovq+KrGwilP38ENz7bB5SAgmXlSRnGOIBuWqYA37fiJ/Mx4PW
a/EDAFxMGVN+QEAlDrkOipM3rR1V6bXJX4QURPTaHALkzSA4rDyB37gFcdF9uFsf
VQBc4WqcoUpHgdjB9RwFkaSNTKcdiITjYt1dWpeHjuwlfB4e9I27w4XORmQ9uglw
Th2ExhOkO8s51CTR7DvwHmc2TM1VTknYV+qNr6zAsZg83FoC3/F4zpTGwcrv6EwA
ZZL7c9AaPaMXDwAhxTHt6zeNrjCKdzhP9TG5jGevP7JkuHHzY8//E2mnxYTazV2g
CuV+DtiEbKFnZu8JHEy0pqn2P5aoC8tCdhz1JjqvZLTxKt5ASLVRyRvvyvBuEwfO
l3moXMxx81Vn6qyp+6C86vmA7vKpwLUBVFmT6sI17hda8Piu88etrcqfqSsO+Z3Y
EopCOnpZHzeXB8xU9VbisuYYBv43UgRWFkhPykZDHyTPoJKD7cbtDLEeccfIEmUp
UC8e0/L5XQni6ft1+YxrV9azagAAZQNvxQw2Z4yVcVCjJqdRU22/U1xDeFAtil8s
Vcw0yFyqEMsr+HVRKGzdclehrWLfwmoFbT8gnuGv1Q5BGtA6veAGefi4aeftWtfL
IkpspvmS982pLaaTYfmMEt+aXUruwAer1LNuDaAOiVuVR/0HVCLd9jByc1p+6B4G
eSM5S3ZsK4S0u9tro7jYIAypqGJcbZwBpqH5j07l4VMsv+DB2sWy2TsoYdF6SqHi
aXbXq6opUZRKktgjuKY1ZH6q1YwAvh81B+EUjDqwhLR1fNjbrcw+VoNsRfZOBk3k
IYNSGv3imAAJHohL21/x5feIJ2ZQxEmsJ1jWNncE5//6RY8iC7bXDvK1GAJCLE0I
uFglGvBaHXas2hlGZIWlE6wLzd/X6pxIDOwmmfrEwikwe7CMImJKEB1fB7+2SsY/
rM4b2L1ocIprE0mkYSOzntKHo06k2q0d2NFgMaU4M3XUwUDJTGGw0d6ErdEwYqBn
29SC+TpC8V8/voiIXROGbCII47+b+oY69cfni3tT1kqDNG4AHxKbSuoJzHKqHRwk
I0SE/CkDV+xIyBY8OcBthuNTyYNII8+dooUnexebJKiPzrBKIMZqWFZHQ+byYe80
17ScI995zdJQHBnBIhWMJ7yoOCpYEYi/ofcmuRA7xNYkZyveDQmCgcM6wMLetX9h
1WuS90nJeKyDiC+KqySdmWNtBdeuWvITv4IM36EBwido+egY+2ClNI8lSCFRnkoG
GImdBLDEroL+QNqua1JzYq+F33Rw9R5O2TD3aVR2DrLidGoxXUxAk8d1t5oEhlVP
V9s9Ia8/8d0iJth32XJUV5xyZvHz01BvYlNQVE0nLQqKdESSzu50gSFYMLlUN6R6
MWpD7Sh5auBHqVkSzurCuljs9yVQI0c98NL9YAaBL+dnRvAf2Mo5exZTZ3iovOqv
Ef0hL+Y4o+3ieSf9SUwtJnd0ZL/+x4fDPY62Vzxtn7yDZthx3zULKeRD1sONdDT/
rT+ueprjkmgcoi/PMuwjVTo/ATIRVydsVLNlsdCbQtWS0rAp1jqoljHqVZ+/e0RI
NdLiY6MVx+NwfORTcjRKtXFtEKW2bakbFxIIDZgNM6mEK67pjnTPMdIpsSSgVlPt
ExFeS6zJwH+gBR45zQyrWW3PCyynZY/ZucoN4322gJxbWscvC2BtNetci9+UrWy/
EUekcILW4mzP2xJd6M0tfHDcj/GWJBn+bx+66QgBkchAHJG+WzTT3HyVeFf77BfC
wgeaFaZRxQ1JJcTMXN9nOqO8Ppaqyn67acENFOev5/7iSt+ebCcnvXkv6+GWfO+l
9w5xjpNXUbaIrhPDH6/gFUc2B8Suxojs2ZWI12A24CwbaRB0YazXNc4ABrKr5FX5
XTTTHpfjOSTX30GBmpfgHunr8DVL6GxG37uGohvNNN3lBWMeGeq5uCLAujTrVB8w
T08u0aXWVV6RriU5QCg27wDo1Rjs/CW8y0MNw6qAnXRrqZ7SVQ6KkVDnNM4MAwKN
xP564986BiIx1d1afxaGmqM4aFn5jCa2CKOdW4f6J9LLMXwfJdL6bvLnkGZwPaH/
ctvSyI3m3f5xWegKtREkYILFrC7ED3ouNaIt4j2i7Xls2Tr03zGmMfEvebzpm4fD
cCmYxPZMxgtWDsDMwtqD2LvC2uNycj4xe8BJuyvTACbfAAFcoIOG64haTyX95Rgh
JrBhrq4RwEjnmrPF1oy2+5Pv8z8+N+RldPHs+egcHhQPDEo8r4ZMvQdU+Ds8iu7m
4XgUT58Z9bQYvSXfo+IriSTRy7M1LejnXOK2zc2FqeyTDQNKkd+Y0S9AmHiDcIf3
SlpVcQnKlOPZjaprhZPwGEfUqG7XyByJPnb4ZRp26IHnRKXQMka9DRU80k6Ckhx2
Nj1lD+WskVjC2eeLeouQKfGfJ6zrssHJTbYA8/O2uAhTLLngoX3X0ZEnyflVK2dr
+ozMhFAUYZdg1Eu4V/La7/ZT1OTfj80gJ0oLxOAD/r2LvvU3WmgELJpntq2UUVcU
5cUJdtDs7OnERh5dla0qJKrkeMMwCYXkMvl2S64AcKHOetP4IRMOPU35+ncewKr3
DFG/23UrtWSOd/QjFv6D9FeJv/E08SXxLBB59jR9YazyrJx4fbsMj3hJ0JbulsqV
qCck53KY03CuJbMqRsECyY5WoiyWSgWvjIkAL0rX9nTH1iPgEzE8DJMpgLOBz2So
kQwLwanrDlP+Ip3X+763luD2xHPP0+xMGB148Ao6e9A08T0Wk8qVWzM1fwbDcn5E
fW0q2WiSLXy0qVZfTmQYuX1Kx8lQHJw8GeWOkl5+Q9DLwyf3UnBLZdDs8uZl8oMd
QYuhHEMMtOh8cnro7NtVX14+7EAJiSjeaG5Jio/NHS152EbBGLsYcSKYc1khFtvZ
r6swwXV2OHHotdR4kGkTwOtE06kWmooySTHSBu+DOKn+BLZV/7bgl8Nt/vuKfMsm
oT8633d0YDr5ebgEATHyzEQXz4tL9LZZqP7V1dakZxZIiqeEOd5futp9603h0gYe
JZPVCiyWzQ/jQ0VQAt50JsJD41KdoBg4eI1HarjtHDBVjPUsnQl+xGNb/Bj4icHP
pWOkxqIREJ80R3+o0Zlb9z1L08O8du8DlBj8z+pCsMCNoTq4Qo0v1nYuPShg6x0u
ThKnWOTl2ArIhmOmgSB7TyfIeBgivkssMzIQJPd0MIApRMkjijZphhDki+9Zcgvh
zc68MRFApMK2Kt/AkMu1LHZGDmdgsM1lPPNPe9J3Md2ILV6OqptkPTZ9U8OE9PJt
6OcRwmbPOAXtGPb2EeHrU3diQoX3KLa4M1g9fZGtSlHMrH5qm8R5zzeEUtOXdeXx
KxQ0K9YSlF1ceubp8oGJU7ADsJ0yZI1CLebZC5oV75Pd6k4vi1XpvQDa06scffYw
y3YkDJzey6zom6FAXM5XiuQw2Z/LSOLYUEXm6HYyCjMbm7ElLOElN7/VRhV7/4aN
XDkv6atoQHeV1SXv9r5O3STmlyCdMoAnTzKLWf9joiCV4pzAWWl+N1lckDH6r/Ef
wC66U6+1oqOWi/FHkhImetHj76g1nfyGkS28R+o0il6mzbY7iybb43QZsywPMfDY
sjY8XFpcla/uOlwyLc/d3jZA0W/aKH9Ym4YFcSVvJW7HteH3WDwe/uGX30TDTJq3
s2bECObWb7Mi/pQiljWayN5TBj6NpnztEx3v2CkCR8cnkD8ufdufKXnxMyr4cy2q
Kc/z+EvBxBxK4v6ZpZKRteBvPNvFbff+71aM6aym6yHSjawRoPSchFE4MdOIM6lM
78/NfavPAdoYDNsvaDvOflK6sD20bHDiHCnGFRBl+tQhmCdQ0m+O5T6FaD3dlIly
Ylh0pDzL073HucNJKKgxz0iflMwygITUtamBsCBWp1mcngbXnNmOPjv3dTvYXdmq
gcorQeucMRECID2qfG7VMKsEtsgepV3+6aF3CGK0UqZfSDQFQvVRtUs8lcmaGvC7
OqzD62JtHy5nKNgSrzDgAn1BC6cLthiIz9FsNVEgsgLtr0g2xjdeous5pFbsHqYO
x/4CbOpx1v9w4LYcx/3XM3l2bPKUOQb1/SjgJ0TLX/xp0c7hfSWOEXup1dFolfsZ
Uz0Fm6ADFvgWSV7gmFBrPeMcQl5bHOINxVDXibnKyf6Fciwv2L+3xb5YFOg785f1
Vol+eJ/gRFNSNkCbgCPoC36XZK17Dzuo2Dz4vpM+/Q9Rsq7SajPeJgAkk7q4rS3a
gFhvM/cIpRkyaukXuzRZxD2YGHPP94zrdSkqFn1+UN/IRobnC9lmHbrPs6Il36Kc
LCqmtRiDiT6kk36Za4dkWsFWfq8VES/EcgH9D2QzFyV/GuIz3nVIw5zCRe1U4eLW
US8s4XOXo8plnPcY4wPOAmIl5I4v2jHzdC/f6C5DgN85MBxjz62tYh5lgGKWoZRh
UKIpEDIitS0R9R7Q6CgLpTI73bVdO5P/4SmvZiNrpPkSCxVRoFasshHlc4d+gUpz
QkY704733N3bLa6FmfuD5XCQsDuQbpsdPJM9jY/iYwO+IzIywVVc3834wk8lI2ht
0HqOaITaSxkLDoUu3bi2s558VRobw4aRzAW3me31VTFjNV2JqNwvrFiJjLBSLwrf
PXRoYIhLNs7pqX8aCpI+tNabj0wXGCSxuiG6TGk5rpD7YBPRQFTkR4xRLqcAblK0
9fYzqEmYT1WQL+CTiDmacy/J3WHcsarujbdD8eC0gHEM1uG2uh/TI9JajRXMyC6V
AKZu9uWAo4zQHQDIOSf2SnvJDWy+rlGo8Arhy7hZ8S+Wz48SE6o3yYhZO/ueaP4M
OUaj1IdEmvqkULfKV7Tj0xBuDyfm/l+WgxYam4ElHdJMN0OkdrWSgwu4tg8jwwBg
pnR0eett/orYi9AgE6O9Kokv4xe7i2OeNW8fgIrTH83ikrW2gRGy817x80KJPw20
Bne2JIMublSbjrGooKx6eNM+CVD9CSOvbsyD/9R6mGrzaB4PlmJfarmwQKAgnBoS
uwr62jcVkKBx7I2Bead27Z+EgEINPguWaNgzbXkdHNcEFxrNQ8ZAZ1ErElWG852s
nK5VufjEjZ0D9pIzQZj57F1mQvQM4rVmfvazfsBU/NWlTZD4Wyd0vjJmgaljvlHW
Z7geu+VjELgB13D4sWf0nHLcBS3ws9y1v8D9YIgTLCQX+FwKFBi25JgVO0akmJ5M
y0esPG0exFCmOP5w+b0bYGJ4cTS9g65XIKqNQBKzA6spqd6C46d1NCxjzywxvStA
/ZIj9WS35J1Y1nPBft7kMy8Wke/ns4y+EF+6TJHNpTwxJlGYoIvmbYgImEZA0XF5
uxCZmO7G7V9bzUwre1O1f07VH34BYiwTlUOHX5agJA847kVcvH7X1NDhxZ5+mrL3
jzy14SrY3AwIL72UGat3fynsJdInK2fC0/EWt/JwbjwyWS3XKOvh/KhpwBed3kRq
Dz0tDq5Wc6w1whcrN4cZR+JoEvBq0Fi58kKNnRrHplhHlKvgC0vVDxQeoIGheD5Z
NPcvXqEjc/6f1cJeUZjQ9imZgbKq+FG9kLUltb2v462lAKzfL4vj1wsE9OsDTeYc
StiLv4A41pSAdxnnWGjKqCyulrSXAVKPaOq2SDv6k68Obsi1wFanapmwR0EKTqfY
5skWFZKFJtHyQ7aMKOpn+gi//FCdwZSEhdvRBwmESWVx/Kbua94dHdHxAOBfFydb
M0fBhtuhbnNCfdp3bTFyLjW9u81+S5OOwtK3s/TkmkMGxnUbo081GprJgUXQNGtd
Payt/+RalSFOyZFggCnzkAyY+eNiKzk+C4UfrZreiaTN83i5sY1jYK3JtJKsH34T
ey33WacKNza4V3E+ptgms8NxyxbHY7M6bxRSWGCH1E2a2k9AR9zmwCfTyr5zr1dI
KtQyDSO/cFvyc2B6ccRoEuGCLHHD+Xs2DnS1XhgaYn8YWv364lGoOtDqCPEZ2nS6
7HneAYb+LC/88ZrMdtvaG7NyoXzflJoptJJ6jn80Oa3lZwck1ITiSDYMLxjPiBS5
dvMVbeoMKajeSngDs8JLjKBY/SbtybOTUgbSlvSoVSFaq7p+GsRlgp0APObyyteM
BkNv47xtrNtq7HSlN7UUaSvEDclTmm5Jv+wHWiaRZm5YMbZYMOqyfBgjkk6OU1n5
l8/aZdYrep7Sp2NSM+WUzBqIO3pazCA+KWgHFXewCS9WqfHar9gyWgnRZJqd2uQ8
XDQslaEa6BCCJ9iEnt+q2CZovu15zBUI0X4tu/qO7hb67o6snulU3CdSPBXwz4x9
uq2KVZY+EznoAEFp596xDpdGoq0PMSf2YUgOyWpyBnp4edS5o5fG3PO2dE9ARF/k
JB3joyMMv86uVNdTMzlNoN3NMRPVC95jM2gVrIccXbSPkG6jpH+Y3Q3xzegHEA3z
OFSzdHWcwFbMn+uxWpa1sFMRljAFH0nwmT9seTNTAlP5dDCvtIZBZFezJsugPUCP
hs7cYIEuF889Hgb+jTgn52/17PNDS+2Twl0tZZznKu0FKpTp6B318KAhV7BQ+byQ
U5O70/vCT0UA8QMT8RwhrIeXy1xmNqeATAflcI7FQJRMC2EN84CETQlWKolfxIpA
5VFeiWs7L4WEywbRmKElNwEJc53soCnfHUHolwoQkS/T6UdblepM2hgf4izuGQtc
Fvhm+mESBcIzxfa35jqfoDar/j+46tPwgwS4cQH5bwE6nkIizo0a++HgSLkDoKFh
G83MZDNzrt2s+EHs2A3Rqv4IfzbmsQWmSTGyoehRQKJfJgRprVk9PSbnKBsUTwJm
2vmTp5t1Dew8B1xHJQejK2XBgJx6e0WsrbfliV9HJd7rmgJxAYSvcdGdKXMqfAtr
YM8cXpQNAiN3wL1cehms2wTHTdTkCZhZ7k5azMXBvMdNnm523P0djxZqxV929wt/
DjIboJZ8dQ2K+yvYEC2ZEVQa0jaFN3QMdsr6R7+4ub89n3BLfHPSEqJyDcKELZ/R
O4NuHu8eOyullOf/zj5XYBWiZ0OUfs3/3XxH1DJ3pi/C5XKpuJkPgUrlc5l2LFcl
T4qEiThMr6ClQ+schoFyyQb1nFBGex8msL/xx+Pbechz3xQGXheTVd4aBMK74PVt
oewA7FcLwsrnqHmNo0r76mAnSf+K34cCqzqegCkkEMytnQkU/pJxrmbTLXCVIVXr
wcN+hcb1RKTLGuG/FF5zB9/msaLIxgfnuls4eYYIwoV6r/qjKS5vU2d7emfcc4Iq
WJawgjtDj3pWorHjAxvoBW2t50toK87A/yrXVlSFjxCzS8GvAjr60MZRWQx54KZO
Nyi2z8rPIZBkRY/WNhCII2c6diA5TnaLa+TDdqAziOZffTodMXBEylg089HdmzFk
IWqld/hOWBpndrTUI8X+buBbq/mFE9MnNGbChFvezF050vgyzPHNk51b18Ba2f2Q
ZiS8MBDWfMYhB9V8She1Qm+Bb0/424ssqMRYX+5/JP4FsIGkm1Wpnjw1CogE4rln
EoNn+Nb2Fhff9SbNXdjbrR38iemGZ7lb4/jX2bajAxMVA6G9gFtK/aq57gF3Ww7B
0fTYP71Jt9iOMAqO4jcK4oEO/uhkC2rJc4d4RFPFpSu9HVZBY2p99il1j7LRKW0Y
meszOybLaT1Oe59+k5vH8m2QH3gUgnrNFR3dG5BRqpIRMLJ9mKClIRqlWwZsMceX
pLoQ3hticYMBePZTpgG+BWYGVudmvRdihuGetnnSS6EBQA0j+m/SLx6Q1+FDGN3q
Mi/HT6Ain3By5JBRs89xCbitSvlmM43ik5Svp7PE8BiLUS73FcFFfAgcZBtfaqi0
/nWSGv+0Ufhu9+Tg0Bcm9bszALk2H1O7nTTWgiY81d3QUOWaO+jFVhqn4jJsE4FQ
ecTEA96Fad1nXkzTX3czYCHEPcW3V3ZAG1r5eeMdYR5C6OSqze/f3P41c+VF6jEK
GcQHww8Mv5h8XXg2ywvn82h5tWNWpZw2GS0BNxlO+lEt6ng1uv60VCATR5BW2AuV
G5AYOpk+T3ni5i8cUD9QTRnyqPkwWqqhJHMgnWAZAnLpktPkCDNWHhluetFBfolm
jlhpoYCxQK3qOB1B7RpI/AqYqxgOO3++biEkTKXrqzNRXY2ZNm5TP9P/Q1WVfOcz
4Lkh9/b+Si5Z7pQWcWfk0NUR3/rll/4ZaaWLtSY7359r3TUKxIeETt5W8GpcEW2A
a7lAW1riXOmjtmshKulwhh1n+cJYtYOXG7wdAZwCZOgs968AoYPy5Q1K2sM9g01p
Ya34Hi/CtmJfv+E00fmkzqcrMzE1EQfgWiPd4rDIJb+78NmL4kdf0uZCz57UFEo7
X5Sm6Sv8WAlPEFy5xzIJxyZUIGDa/VsAkEMCfz8s/biV3IFaxo+Du7AVZGl9ZNw9
INQHytwSuLwGZapNhOy88o32CEnvc0zrupVZidyzjTIDMLvrWoo8CoBCKhIeyIN2
G1EjqgbNFDzm/ko4AvZKWT3GFTVQ/jIEbS/AL1KBtLzG43QEYEjIIiBBO8Xddio7
+MO5lqQpGDnYLUhrpBZDKXEMp22jR9AINxX7HkWcbF7W8kOOgycaub5QdXkBsFkM
KhNaVjktiXuQen76CZOZ5PMAsV6AuFSUqxX1F+0G/YHYmLlbVFKgEG1Rx+o/86Vr
P6WAfob1y6lT/a5NAWhGKFZM6aHwoMhfULqy9M5FE2TbbLqLb3GgGD70nwKR57tE
6RxZhdNid1BcIQLtq2Ih9rt42Op7XrPn5n8pSsGaf3x29uE9yTNWSSBlX84bQKHh
1BOGmAGx97JQRwPHttkefS0ICrwebarXPWsFJHj2QS494z21wQtoQ6Iabv/5237v
vbylNxU5WqlMkO9NJeHLNmY1n/W4T/e7qEjFmDovOrR3kTnQ9AWLkSrhrkF22gdc
d5dk3YxXau2qUEUto4Ifxep/+Ke0ly35mtyboq75clRFTuUhZhyzKDZCYY8qu0+R
96XPNs6+OkA5zGaYb+gUBTy1vCqE15bCndCT0eZoKOEyFlZjbghBBavi7CQ2ap5p
r3TGYrPhnQa9j6m1TfEfPfKDxnG9StJZmGrLHBVOU49grg5e3deNwjC+morZ0Tlm
nM+uJ/cpfSQqrn8YiEeUQj9F/KOekWBEtzWfKCvGz8lsC8Jnp+S/pWVmE7/fIdrH
ounoYmuvmusY4BfxVDRvbmg7raVBYM4ciUc9Ckcvgsu+CNjcyKdotn9BXYSOhnxW
dJkfUiW02V+RzgEbYztYdbU+GEu+zrHgrj+HIc312ApjH/xE51E9Pyt3B0xpqj84
ijeP3NEoJK/mCs5rRFg9OhWkEnozz6nuaU86iVfGmKZp1HgoAtKrSriMRcCzJ5YU
Mv2fdLIgqNWr9UmUnnahufKwUdi5KJDTNJgZ6zBXKKIHWAqpf7XXSaQLzY4NknBP
CNebVNN+gbw+aF21x+/LybMmH7quERZz+V8cbLkyxm6jWHvx7jwOmP51/YUULTkk
N8lYNwyEk6+Gu9tDj2tQUKy2Vt3zu2hUd45O1FO/oHhvKJHPP5n3+/p2L8H3TM0P
U6qwRPOOPkdvnNpy8/w7pxE11Rlfqf0gzqlEMrbYRiNZg4GF7Ev0tDQjoj0C+IWK
VeuH455itQvSbStMT0WsuxCsizZmDPM8E0/jBRT0bGrhUVVXYvqaezQ5D3J+Mhrs
i0uLEkvk+JUOGEXOkfmSjn3h59NRjS6dMRggNASNRuGj54ky9OckKX959vGAAeUX
6fUK/Z7HUyBEXBeIqEee5bcte7dNh8sfyFhEjQek9GRlvl4HkUyBmEI66WRDI/Xi
w3r0DurkQYts3PdizwP/qS4/dLEr6zXYSiTJHZkN2G5SHY80gZ3kDWtC70bpRvAJ
5rL1BzSOlUu76rQLHIL/Gq3qTWgh6rPtdX4/mLlUGd+j80nUcJk3y1mlr/RiQwKM
7ghVWpf0jd+Jg7zFQ239xhFccQX/R5oe+RL4L3C+S89JmTI72W4fg8HI29oDIbbl
QeuPPtGR7oeAM1oPBATyIDcUEumdnPdcLhMc98q6g7mNOev2t8yVeUc2+akLAIAg
ciXkugknuZLAkXdWv8xRxz2OI20mjAlMWg5w0CGqFsMDRxRR5RmU+g/r6KpoUCWn
VKrCPHbE2vx/S+QQwk/u4S6tmwBRDzGFgXvBRTx+n3kPVEI7BjlmG4OckCInJjnI
iwFY0DE6hxyrQ/GPDU7KUBwI2z8KhLsVCGXcfTrs8CWanuxvTys8XWhlW5j8Tbtf
WH2G548mkOfyCdp2Xhc1ghlAkv8V9QJgeddz9u7qoe1izo/Lssf9ACSKYsquemnd
tbNrwXd6FiR0Wqzyii/m9sdVPqabF14QZhj8t358eJfLs5kwavhpLhcX5T4afOlh
iY2Y6RhHwSR/Jgd67DgGPzMWAekWNbAiyd2XTTNG+hbEEGLh/Bb5oyXxKCBn6dN/
cUw1YcjyCnQYhbj1Wmp8p2BWpsJFLnS6kCPaHdBQ3Mdm1vRxd9Rjb93CmoiXqhEa
tIPoPPelrCdJJ6zUhlkKy3IkKSckbUj0mE1832m5i8iSukqCp5QfNv4xnvyx67kX
3Yr/Seiu3cY8o1tdIFckR+5H5nJGK7NYUIf1sucfm0irU7IfV0+lI78EJeCgXsxy
SrvypdhCRGLT/utlGwaIFG76gkl0Y63ALGOQUGNfBOALfep0WXUQKnvsd+KDAHil
TVRfzjiRVOBP/FENDoYlvrc8VpEPSuHsTt49A7w9H+C2fxlifXhmV4rdSLvktIuv
PbNkCajS7IE+sWb4N2gJmII+7r6FP9UJMgOtga/ndkAL0qOEKU4f5n5VEq+jtaLD
4tl7eEMaJ3bAgRwt9y6+IBO+/8888KHsHsaHSZ40jAPq2xo6dohboSyGWuG8gOXU
3du0yQ05soTkr3XMiT2R5yjm35h2jajbWfPpEwUclsJpY4Y0VJ/A7YJlpbKq/f/F
cbY0nq0Gej+7Fdcb3hoquiERu3G611cOG8b8cQhz85tJyKVpbvJyqp/zvqt6l3z5
xfE6qyCTVUSgz13oNcov/4bz5jdAYj79fdPVSmkwWTlphEkURG/LQu3hwNrngkP4
lurze7/LbzOxlgmHWlpt1X1PYOKLkj0ZQrlUQqpAzFy7/wZYXwKSu/6U0O9RuyIu
UVSVtX7T3ITzBYqEj7p7/3sMXiC6wJ7anYFhfsr8Sovpag1RDk6P8otTYMojDDY6
u9nPVLHAJ3RLNowM3GoesIrdE77+SCt4xqeJb8kStZ0lZM3Tc3vOKrkdwghoUtAP
8AhkIklv2uWs5A0elCI6St/vT6EBe5eAw+7p19YXKDFf8OeR3w/7aqSOyT1StKJE
S9r8eJMGAhUqFzdIfIUcabzzeK1bVqVcGX3gzeKHQmU4Hwnzs4ufmlItHiznWfWv
MDq28oJdqi33e4OSnHqxLfeSP1T7Ett86XYwqZibUQUj31W41FHTSweUDJEJaMH1
K+kfnootjb+/gHkF0kVVPnkU75evpDMTf8285fV1eG4eJTybDLrAlUGfvE5sGzos
R3jioSTTGcXY5m7fXfIfss4YWu/apwlYeDdQ05rBpO3Vq/nDB02KTj/5a6bQcrN6
r4ITtDYGzNIQ8O3NF7JAEXq3TY+H0LAg6l7HyCBujPAmG1pSovN4BhKddQLWOabz
HhIGVTxvMgf1EmAomGqUciSmL08FDt7HuJKjFifVbfenqHzFjp57ZIKcyxkmQPyu
gCPze0OnLG86qxFiXx3sgy1ZJ7gz3m9ilUPQHYzX1hHq8M+bR4Ai5n/ZyEBSwLig
iztU8MWrVpU1Bh7VW9pv3N7vlvwYK0IxPQBYI75RFi+4S9/OEQHpwuK73ysRMXta
0U89BK0LfD9I+YNFgBjBqUGNA3ArglC4A3glKYt9FJnufA6dsSJB3KDPJi7PdUg/
2ELhNObgrwFgZAIY7tMU0904nXjynufUX8zBGMQjBHKGvPssxdaxRdO5YIfeOOlz
5tHqqa2DTYnTdtrsJ41EMJQ6Ry/DdwbJbjB2Abkf4eoayYZsubvXAvLWkYTgEZc7
3nQSmBmcB6E6HPhNUyO2g0JPxH87SgLO7FOR56r1x3l2u9SyX7BOCMWA4qVdpfUn
yTTUtkamVZndaoKcKE8s90OETJysWV1CB/5K0ZstgveTMKJTjEvi6dvw9ZXbH10h
CbnLlG+KlDMSMO0n45ROYyMyhPSVgs1oT+Rp5nviE4J9y9m2I8x1idMSVQOG3eJA
HnaGTgVa1oErPok7ia2f4RfzfRMy2ZyfLvU9ASVdumTzROung/Y4Gv3GYGmJPeTM
QkFOfy/TDYTvZjW1YLTnXZ3reDfMDLcslmpqlQ9dlj9dGgDiNQK3Y7URORniZL+9
b55YrgQ3BmS5wMJC7LzuBjjyAgtyo1Q5WgxDITQx6BsB9hmcPEZCZzXKSeoZT4Hk
cwTCDMvznsGWrA8jaVzQSV8vZ0IkNTH/WAwaVMBlry/ma1cfK/XHqEFqqR1xId4f
ja/1WLX8fUfWBbkgfBhP6ydn2m95K3HLh5bzlLUI4DDI7XU8VeQ/R5W/BamzXSAm
ndWVIILARGGVBkWiS4ZeAjcwgvxsihf7k0ONQ4QvjXLyU0VIyjNxrqxng8Zd3AbS
Uk4YlJz05qFL/Nagw5rspBw5n7dN2YH9N709lkN/Dl1WZSdyfwT4rB0wl42w2BfX
G/vSqaqRAMlmBxgPexyHvVSPqx0fA8qVRfT8IiXuW5EUnBxqflwIHMeLWQliJv//
pae2BM4CSCVtkBKoFALWxlHM9sxWATWUxc1Qm1udN35NZ3ybNzUJc+/5+zY5hm2N
PdwFbalwAj5oz1aXD/S2ZFlqJAiFwKJ9aOkvVtXbeQQBnTcNpTtcbBLRLAi+DBwC
67Wv/6lUQsudLNGV5zqYITRoQxd2fR0jgh5kLbM7uRCDJ7bJBfs9oupgD08xGePV
ogMugGLxglb3ogHDmX9/kRPfnfoDprDrGYMSzGaGYVlHHDoQerzSK8FCvclh+vq9
EPqL/kBX5tm8afseHmg3sXUTYe8WxbgedO9jyNilR4yc14jFsv8urXu2UtSaUe82
gxriEmVGNIbfcHM9Cg2xLIVz520R5HAm2nBB3pnUjT8ztIpf8J1bXMHTov4fNAe0
6Hi1fc/58BFZdDc+QG3jm3t8DuMMeZ/3YhJQsYUJV7+Ah4aDoupdTqmilAtbuPIw
Nu0Jc+KnfMqz5eADh0AOooSFfPw7xlh1cY+Zqfmgjq4PhMVWlIN+a7AeWZ1ddaXR
SQhZLtKCCUSB/4Ulubghj+mAFpfIMGn9L3EVqZ91VxY0ObMsvKzXSHpL3jo+q5MD
XvVMPP5ymwpykfDFvV4qnR4RU0HpAQGHyYmo4wspPDybqKLLJK6lYN/JJG4hH4Es
ibhAI+XXJ06DFKOTNIeK7LVoQMbu3MmCzjsPbFmgrEoCES3TexHJOvtkok7M7Oc0
ngX+AV8v1qtqIYfH/55xxWYckXo2aZS3bplSqWzk1qyqJxl4iwASBEXcrRqi+jzL
TFcMSTf8OHxe8Xf1cb6N8JsXfwdZbZaN/cKeAV00bVWdPEfxZtsjNaek8g4dEtR9
Nyc8lFfBhkC2W5qki9/GFD39osJCu72Qn2cS74nQG/32pHxenMn6afiZsoJ/F+hP
kO0Fbnp48LGETvVr1Bpc1SD77TbfzGG2BEzF6q5o/f9LdXTgh64mhmXmRlB85LXC
E+e0Yo84UbUefZ4iqdqqsaOkzyN8OORiATHkbSxiv3e5IsnNiJskkDgqf0Wh40sf
Rjzq2LWlr1CtkpJgslRPAH0tuLQIwBC83b5LfK4BOegvAdmlnsM4VEivmswJ72Su
2+Tsl12Vo+VIiqUmwE5ro4R/wMsThsrI3KXsCgrsp5G1EhDSTEb2e5hfvkqUZ6DT
yyzNr27YR8sVfSBm5wahCMPQjgZ1LtVu/GcLIdmnQmxw+NIX5vnCk0pgcABNRILS
Km9YNZWCdbTX8R4RJqig9pAU9k7EdUQ6Q641gWYQZS1RQGVzvxQvO4dfrZeBB1Je
FlprXD+ldpqn64OEqzbLK8wOf/pfd0Wh4+ytS0yaUA9bHHLphUB7RMIkAtQZkOkO
nsDAnWY8CoQ+aKhUpdL4O0F/vawaxfBXBT8UYj6PbcN7enk9GmmhF/uFnrhibI0d
gNMLA4MVb4MtM02DzS7vim1eMETOc/LFxFGOAVejUCUNoU7pZ4MRbMu5DI3AQixb
ADAvq3VYYAMHeIYfgRUIxe+0sVCccww9e4pZtP7cpce2x9giV86gz1N4ozVmXAns
tOP/Bqtl45eYW8m8ZRIj5CNsdMqZdLQS9RtnuFyPZ2h6zbfGVrUB1rVh+P02cYVm
9fuRtPGc9s2Hu7ATxTryC7t1LNDpLaXFjBRIx5fujDWAkK/vLry5vbcz6sKP95gq
Dl3LWfJv7KhW76Z2xGUXLZdnp+pZWLeNbSh0DzE11lOkC96pe1yL+r3SZv1VuQTQ
FFS/GlpL6h7ma7mAXMxESyScQ98L/npjJyMD+YxxjLbqjsqSSqpAaL+bKRJKLbve
2ernnRljVDfuAUwgThPAuSVGm0yvmtgruPXSI4n3c7DaZSDlMgUtYyAnS4gkldZB
37gdKHWhUJ3sy5DMHCaBnDMHEDsXD+caFkoaxVPsCfj2qlN/xHsoVRSJR3xh12R4
koe2sx9vL1wX0fQiB6CsFEfC0WId1PQZIvnjThCsNEZFE0V7xr7JCZEesotbqHfa
DMJqCZDR7lUk6Sn6xItchI9Sim37Ol1Q1fKZGv21IXm0TFTKrtOOeWDPYOQP8MXT
o3ubwJQf5mL/SJ1/tQLC062AWeIPu9BK2nprBZ7Doi4o0raVJ1opXB4HGypm2THx
LkDWxxRqLcQ8Oo4eXEPQX63bmVR6qbpwRBDUpO0F16XbrW9DnoKDkNjLHMHaRzep
GZvq0PIgTW9Dhkrp3v0WDipw66pFnPT4ERfGa9tOHcvwjdKKIDzPrszJqGlPdt5j
8LSdSd3/H5ocufDoEVNg/i/e0JWOOVBLmLh32urTxKd/h2onxag+JB1oVoBzi6eu
OWmC+enMfbYjArftfZtbXkWpx1JtdoNyYRjw4Z2MfNDvRYDa8TtbZlb6cvr0qUm6
TXQSOKLhO6mrSq/82gCyu7/P5izRNdQrjUCBqTcHYyI0DDrtCGjvdycJX67Y6iJd
6qIB4bb0OBTGZkjWMOSoje1vmfej6qBK7xAQsPY/PAjNm1YmfJX3656WR6IXPhLj
lIupSZxgFor7r2lcCPX6bzlUUvLKlO4dIitnH9cuz6/c6exrbtQlQTPE79CsOndb
iNEKaFSGfv8jFg2QF4A3ICbSnN5UKuWszFQhs6LfOP2VdfxKZMI4V5rR4B+A/EDd
9Ef13HVvqHGcSe6Vx75VujWrjkhcEDB6kNZgXd8rq7VOZ1gjBO6AZjL/epxsl1cm
abvFvJFrkyaqxNA6c9yXinB7dB/0OsAMWTSbGEU80MjqabWKg9QTepSiq07+ZQYA
jSNOh19/6KZtt1fUy+/k5eyz3phR+eyRYTKDip6gxcDOPddLJYCwo9RgKmrSUaxL
V95oCBqoCs7q/x3qP5C/13b/x1NqqvE9OkTJN3lwyXwvwLP1wYdzBM+orXImU/tg
wW9iABt4Ev74LLlpG7MbVfjgd0ZOf19gvwbJ4xABzpgUbfLRqmUvlN2rg5H6xXY4
SVFtWwtFbWKv2LpH2KtI9+4MO65D2qxUcvZ4JGA+cCRuavGn46J0nh0A7s6ezI8l
K6FgjKmogAcA5Np7fFwQjgogW5FWm7yWbA0iSl/4KXtmOGopHBb/WegDr/SXysIL
KeeVYH/LmbShM3+Wlwug/FU+mDuQdAuKqrj0f6ID2EiQ2aDpvebcsjKjZgy9IkLG
k8JkorEZ1Wi6kLhO0H1zptbr0w+kE41rS2ZgsJiwXXofRAMOvNy4YLdYvA7JJveG
706V6vsSSQuYSk2Uz5iqX9GFkIFwT1uhEVGFpbxzxgxRjGceYX+/W0wbskprIQ9k
X2VhsWBvoy7DvljFMMkf2AZedzBaUOz2nxynH+hc0foy2/3P08Vz+MLB/fcjyJgm
QpH0HCGz06vbI2MKmcj7VCYlXpzupT30l9VgyjAOW3sRBoKYqoprraVuGElrj/s/
t1DTJpnZaQZ4nHGK8jftwCRC0ncJOdzh/SnrZZ1LTr2yKmW+YqbAGSP1TN3VTFii
zEz6DbGaDEfPDWFuQfhQKkFmRzug5weUqMrPhK3WOcBcnvc8LOcZLI8L+JxMLGw5
R6ODsZQ8Dlrb+TBMUXzIRVF5MWCvGQz+e+lm/zr1IrQ4YSAl2k+FpcwiB/Yvlumd
Wkt+caaejisqfC2kGyRQDwnivzBPWewq9dmMqB3W5qbalV+GVGIjWvWECJOphnDJ
IMWnlBvudEGpP8Y67F2QWMYr3EoyM/jSUx+46vjcJ1/V7Cdlk+MeptSu8TnyOBuR
WFTdFCgsONZfv532jlkgm9rcEMI9Dk2YJoiPcRp9slyk2Aq2cbSjCatyQ0oGO8og
bODD1UBNh1nR4+InOr0FtuS+KVujUb214llkltcWux1jSrqyL+SfTD4ZWG9YWcXF
kUvUeRfpQlflmZ+oCBdhB6dWR9ZSTUCXnzewO2VEDu8M79zM4NjrS3+XvT6kpIwd
5mf3p8cYpj8RaVxM5RgSW+ZPxEfZ1GhUzTjyRQu/hpcVMzwJzfXzZMETv1caWGaB
/MuFTYa+m6Uuy+KtJjahl0alaF/CQtFYe9zmWxOlbxsC9ESo+0yb7lvHjREzLb+9
7azrfowlhT8YblnlYchOLUCeCL0wr+5GWiZttmvcPyHRjLJ2BJfq9Hb8Ibk6mzTM
Eyl0hLkm24extdM1svyv/Uj0+8zhvD5Lv43dc909Qxk85TknyODEOC+Kr/+9g6Xg
mu98vTtVE9OwoYgm0cFHOpDgaUdmi81QsEwsKCMTeJnNZbVS0vvqLJRWeSxaLo69
mUIxz+b54aE4VHgbeKKf43u6wCta/0hX9RfjGSfgLUpiHpk+j+cB9nxlB1RPtzzf
Rh5AcwcbyvQEekcTi/30GRCVefOuJ9x7d06wAMIA1dbIdOKrcqDTf/arB8YDDobh
hgR2B4ebwFKLh9yFdma9PSuzFJp/NAtahpBqnvrJlgvXORCqyFl+TtCf5apcZo/e
vmG2ZlG0XI6XFc7T+yoCTjA509feP+anad9WGCmwaPqo8MqWVTbOVjzdca8eq0B9
zN+MHLFOTgUtwW19jMP0zTEh0Z+q+ieP82x6VGhJQsaiUQoUVYlYMjTg9MFibzbz
jlLF+t6sH19R2J+zE3FGCPT4uk29ycUmNi8QyZfGCTowMCteGFSls0q1xEzyueDc
gq7CnUBlW1vLcn9x3M6hU5a4ziOLb4hycNHvm4Pvmiw5j0ZRlP48MqQBHqXdNIys
/td9SVPNDPZYu2fbImJ1E1waAFTemcfcXoMafrzqQzEN2K1zFTBMQNBcQepGuFbJ
nt3Bq4THI2+QAyelLPT8jRyliymZAMHAGf6PHRbt1mP0Jqqf5MeUzMAeSbZ+ORb2
VZi7nG3gCPdkR5CPCshv48wahe0xxPfrRovJRnBq1VCaGatsK5Cz3FlHB2Qe9H6i
H3nIe7Gd7NueGK8iA2MUih6BLxEfl9SynVQ0qEw3368L2gICmRXpwrAWXuWcfdze
jKlTqm97j0G1GiNS3WRVg9rS98GLg+2u+qzyymj7jA3HiIxY38U4nGTKFE+k7rOt
ltd6Z6EUYxZGZWzDSUwEsrqUQs3yXxB/vhAYs21yqVXb/zDI1QVqm/sLbur2xUxu
KhXCss7RKR3wX7gQETvyzet+p7h1Xd1ZhpcIQemvnSL13PxCiBlqL5bEn0VipNM4
9ffVoRUluzTW5lXh6akRpapKWyHeEsiTaGDlQJ2gNwzoP2GYvMljyFz+LjtmNZ73
1+NwUu4zCHwGW3IeLL+NnujBIqBF791ZPjCxREy/YtYmrJFaGh+IDTAOq/BFcQ9v
I+Y+0HklgKyU26wbaa3bLPo/curxGc6bSjWv5awjQxfYJyDG/iwdfHgpwSA1GVK3
56Ai+PlPn3Uj8cFKD1sJg03XE9vK2eR4IvspcKhl9JJMhIeEoQY20+eHsIdCFHuY
2EsRmOpYc65wkXlzBvTxolpYcuXHwNqm9sZlhafiIGyOYjCEmKpgYpQ+5+QePF9w
4vMtk/b2xkVlD8CDkvE0ST3i7ZD7w/LRRCBPJ/wzFoZJK48ZmFhtuv+X/LUkndP3
62Z0ha8/e7bFTLqunrAtOEYd7bbt0/Zc4USXEyy8APddPZaNSCYEPstmagsveZ1E
14jIqP43/dOf9ZgWNcoCbQx6BzQ78se0YZ+VMKe0kamtHGMTQ/IOjUiFLt/42B5L
UXc8RBEgI2X3S5asaquZZFyHuG7OQlgL35HTMHYwPpCKbAicRd9jTCyY1JccxzLH
H0JP2MTLbLPpVlsPP3kh5QrmMlx1eMkqqmVqb9w45AQZ4SdxscNTGFKLzWTSB/vD
ULLaSThkOvoGKXQw2byc34n273hCjnpX6stfC2IGVYLzSbj15dKlZ09pSuht25MA
e+jmTP3AClHNKiMzT44LZcbaz5jhIP40AGHKhqrgF2teqe2TsJpOj13ZOeDAFHso
qUoUN9E+di/bj8hfRvGuKY1E13vZ26Gv/9mb9uzxoY2Yl2R03Lj3e1myjKwnWH8R
BygjHaTti/lNtUEbUrl1zKjbCEL4jhITwARN9h0fEwrcMjx+ByzR/aGA9EdfjgU5
FBDf+4Vd9fyLKElNriMGhQYUwNKDQq42DmZ60/LMSi04Lmh7fzYyhfDBbs+DoLDo
JHsq1/pjCaDtWpTYz8imQJWU/2EGI4T959gdr37MyJI82oiGLzKnGuSAKoJWJEQ6
aHaF1xmtw6VXv4C4DAAUpOW4ealBLdL1PQUr8/7ZO1vRYVTl4YlwMMwYjEDH/Se2
/R6+dhBSbfJZ6k/imjjlA+76UaLUvFFzvWbB60V2RGvEu+LcgNh0ajcHNuen74Rf
kHTFzNQ4rgfHzoqnxIElMXn1JLNt1Q7Umh970KvXvDuu3s3rCfKxUsd98RFVWNqu
1zA04TwJ940tdahwXJ2eA73jd4hVxM5lrJzTlfX9XLtKB4dp3/75JZwRNkghBlCV
0G3YyahZXDhTwLp2Rv5wFcjNErBIdOFZ1HD5zKqyhs/oNgljurX+fH6+SSOwtI77
dgN+iO+dwiHkaYMJs4keNcXZeRT667uty3ThJyI6vrvkyXBmXgIJCzvPrsZhUhFE
fRQjGhTilFHM9ndNFWKVKIi1EcYhLXI6VLTyzqkmMvGCTKGvWwfPvbdYP4rSIFXL
lxgMMILSUya7gyk/KGBrVRGZ8iIBS4CTDWCvuvL/pwpGGXrIxrXdwpuu0pO0kyoW
/TWVKtPgpUkfm+Ydnz73ii4bgwWpHDGpssMGgHVl4Ogir73lEKSn8WtAEHaTRYBR
sB0NDXrfWUIO0M8l2XNX+MnRXEoH/87fjibGAZCkY9/pE5cEFX3ISCokISYGAhra
Ze6sBhWGXVjTl6V0IeDc7VosKmlnFhLF18PHIngjsn+u0pqCULLjZdZzKOk5NjEl
9NpnnU1ppZMK6a8zrPKhYMtBqDcYEpFOjRlPAQqpDw+bRprXChjBhKGnUxRpICei
wbBlnpjBYlCEZ9zeOc4Ojn5Rp7mg7+ttlJ3twp5+9z3oFbGl8UB+yJfYoZBqY/Zk
62h0M5QiiaY7P7baIMWOlDogR0F3ldRCSywTO+4Kp5zBvfa76L2mv0HOYJ1KDXvu
d1pyIGYwMIWyQ3lqgOC1d5iJWKvq/KeC7DuzXOt8Rbpw6x0BWVTaOtF7Svk04c9i
z92VdZAGk47hjYcTrZlGm+PgU0RfdFJONBkc1qcqzNTJ2y4zBdhBnoyo0I/1b5Sa
qcVA0ouh+FS3pK/tzW3y/KKSny5PIcKxLV67p4KaoyMTsvJOqKVsbMzN4J8p3lzX
UYkN4qkq15EH4GagPFKlkwwzJHXIzSvCPqKYDUvNVDllZhRTXHgspzCf4P1OHpXk
/6fFkhFuEsrU2MAL6Zli/77+c6/RuD3AcyO2XTOPs4UcL+CTgBv3L82n+b92A80N
P9Cttq+Cm3ayZPh5qyA/6Afz9l7PNpUMpTKmjVUn2DvKwCrgPg/zAUqWgE8cYymE
iNZNMihJWsVPyLo+qNX0h40EYH2B+zXH8RnKigkYUPPaigQvFQp6/i/n9tGdRRPs
4p2peT0qfJKzfdZz9TOZSekh2b+iOXfVqa3nZMZ/6q5icOSQ5P4QhXfXjAmEp4XY
OWGF1uAD66QTmMHJ6pHhWgANwLr2U7WUrKLI99JzuUmQ3W8+Qh76WYMmfJWAHGxj
FPJ8m9EZAkK8P4vy6MGDNwItBPQYuy7JtPsrvcydOwWPHIJFcSTT7/taWK4iathD
C3ryNIYpFornrIKDgepvsRO/RfKbtRefQheHX8zpRdydPWs9SPZMfXCezSoGLocV
decm7oLHxfvx4n93EPowC4SmoQNvWdVFi959XoUTL1fd7KGieP55iVikVkulA8M4
wD6FTTOhE1UQL8ZZcTQigs6w7Xp0zrSbpeJ3B8F1ZXK83v7K6PZg0nfVyubPjKQz
bfgzX5oJj1uQuW3pj0BJivA46b1ACgn1gRlKQcRPBNErYPMFx3Yh5VkfcShf72i9
U6aG7iICgbWeWesEx+27xZmG9POAdHYfzS/kWnzb9by9LOKhodp16VOCMC+HxfTN
ZIpEw8cR5fzRm1mK3lnZrFeQ9BqSJVHAEnlFLAQCulPmhMbiUh27yIkORDcGUdSa
wkpLtifVEEYZf1Xe/z/xbdOCbpnFj/A2VAhWpKPMzvJHuPW48cf3Aw9D2s9m5t0B
HD3esW+RDpT5I1TgBEgwzeOslOxodeFvMonlmGmu0NmXAVsnm/AHqKzKNQj7vReF
JcEeGTzvtkZk35ALbDVe0PQs/O0krQDFEJNrcSdvimYduZzhRm56rCgO4B2aDCaB
4dvup9/PMSa3q9zyjraOC4QECMUMsEY3djRkX0qSvUO7UziR25wOiVRpiaI1/SO4
Mtd31W19UKBpF+YrH3MtyjQq/iGp+yVilWc4/7w0CgWz2bHFvAD3m0Q1QraSxtot
AqelmyLPHjSLzinsrlknhwXyk+1C3Dj8XeE9226UxGtupaqN5KCrNb92vPrN6XI2
KdvzEOh7xvcLFzrkRPW96kXQJ4i+qfe94q/VkW83m8l/V0fFKC5oGmNsTZmEhYgm
1DyRZs6bOxzrR8NNb2TIzd1X0uzFo7ojqLlhJ9YjiZ7xhQ/9YFfImbRWIEnHKstE
WAOK/P+mncedNfuKHD3f8nb79K+80sP+uAhOLSSvtwW09Z6yGvGney6958OIu6A0
7Oa6q3FV/uSIK3qZYP0L2rn2fwLQwIIORJv0zoaCuba2KoC/nC3LnR5ClWJ1rt5l
umIKIFc9pNeFdszm9nQzGUpRY1NKrUy7r7ItLguvu1zQ6Bm5LZxx4Gf8+RwqJUVe
fI2XpCrx9nfekn0bPW+tju1TYD4c0Bhxh02BHpEXK8vGlOn5wXAD36uJDNhL/ZbP
7ArSDkgiRp4uBUTPEhhRIUe8wAmdcUDmTwGv41A8OmI2wkFgarjKIe05UB4bNeGj
WaVByCDnlUJM4VAy7EpGLxVX888lGkqmcoPOPKjXsM26d9Uf4kRIhgh3j0Hn1Z6K
zhHaK5mKNOPtPzjYRpuckno5A4sQjkdKDyZLFA6mGapz4hoS+UHDJmbxPEvbVQ20
gE/beSI7ZtsYt2cDnxLN0SXjTU55uv8W6CuX4Owter/tlXcxVrPtvv6no+ubukap
rJ/2IaXW6vhwt0fGw4+v9xUOqyyYqpaRIJO+1pUcddKgi8HyEoCOPq0HIFzBLK8N
MkLKGAq6moAeI7bUGHEWk/WPZewI2LwwJpB/0zwPfJtHyatAnbYmhrOO47qm7b9Z
/oO1/ithLY0V9MjGIulIGphTT3pDwHmKfu1xBt3PK6kDBSKNZFKCxd37NHl0jRK6
05bfizuu+i3fRaKmtc3m/I09AibR4tkJ6veYxNTjBYNj1c1gtSB7fV2TwrrzI0Xe
uW0vW67g0CpIPJQGaw+M58sd5yJrW4+GMxbj3ahXPC679YArkU54wzJ4uU/CiToA
y58cDFxyd479YYx9Jen6eR3Lb0imeEpjx4j2UCWQpy9/xDiM/j+u5G5kGu2ewHr6
lXB+zh+dhGfWC49xGJ6TXwkDA8LuNNGp57zUo2ns1jA+FIFV0uIf5G33h0d98XWC
mlGfVrLPe0bbVYl6aP1epUe8jHlxkhN+tBUsUkr0/WuGa8r8P4d3G5TRxfiYzUa4
+JeuTO9pDjVDKz5WdAsYx2tSkLKApBOBJjCymy1R2SyxbTsPsInnXhH5jA/lB7cc
yMk/XocSy+lXAHi0U06RxsDx6vTy65RRlDszVBY6v0570J5ZLJo0kl50OiSSADrv
Ux2a7H/4sEyXXYdpgGLdxh2CMvMbjRoMG2nZDRli/dxQRb2GjSeI4mXTWITwOY9V
FbnxKULtqBpj6OhhyAC4KCICQDBGwzc4uoXGZV5MACp1hHh2JPtOK6ETgXCv5+oz
112100TRQJJxIdrXT6wf+M5Rn1atqy4/IZEDXQn4McSUSmWBIbLvdihl6+JUfmFS
AqBKUoyg1c8+UoljvDmiQ7IwFhSoNCiRvhnQlX3UUsgytuNN7sLOd9+kF6v7RXLq
hMbZtqD9vwTDQ+2U7c52OoSW+Q9/JtSabolJyzWzo+3negFmNKmmUWQqVDM0ER0h
E9PrU2ptsRyAU22L3RjwTOafu4j44ZfaEEftdv5y0p57YoKEiHN/TGVmozrHSTZy
zBzudjgfjovDc4MhW3Fr6hiKitQKgk8y0Zpj9jAwlo6Y/+v6kY+ebAEGnvVyOTrx
/rOpF81Q6wrH16s56r9AOZuk4h4i5Rahc7w67WNh1WSCpVB74q16BC1zXfnQjdpR
5kW1E0w4lOoe7jX09SBRUXE1z5sgKbMUJ47t1d55C1VSNoZx11f2SF2TLB/3FIjw
pyfed8m2p5nEQqV5RKAA70f8+yVg17JrWY8/cslZ7Psm0HUMGp/c7M1usauVEEnG
pqmg5QvW0YfNJqumdWlNtKXvEILMUColxT73rzsZog0CFnHqn+KVRaQml7tAZHJX
z8J3MOTj4lQDgWYUNjUB0vCG0WM9aOTc6AkMzuOvUcS65huLi8fufyxe/MhHn/Mg
yBurmZwzlYsFWOV2kiWawxwF2aKAQdD1vYhNCRXNgq0s1k2qPeYN+vr+uuEAJ3lt
YecN2B+k59oocFtk0s+OxVjhNY0bCvvwtcOmCQX+oTD/5XlYUXOfpjd5pUMnWGkx
HCPxqsKlPpZ1iHWiMEjJb51dNzLPct29S4nsa+DxGpHgEGr2gFBRj2jgeqf3NBAk
1AJMLegDsx5hmFCSYcl+nyxATDbC56mSCVmK4V3Nl5xR3WbKoMhxKfr9tFnQ2Y0+
9rhUDh6OA0Z5DYuKxeWmdUYi3WogEYkUuqyTD2bT9sKnOHBOvDtv0eAJEZHOVhW0
qd+u0FQVo5t4dVz+y4VLAVQaElf7jJGY7YD2KVHFXN0H3w2NZQ/qs9NISEcxeDOK
PBVlnxmfegS3OoZD1UTSZONOI1bMn9Hy18KjJYuDIHHlRO1N66/qdImEUjdldVG0
YZ1QpoUrbFCVHqlod0IsCNy4g6wDxP5B8Un1xBohpl647dhlbe6lJWBStc0T1YM1
i4WVDFmQfbeMh+BdWmnpEk3R9eMLjrD4nd4REVI4GTZYvm/mCoJPvmdoMVA68rac
2WNrhU2HsTZ7xDb5TycQkiWSwtyU36PojOuZqk/obh/yNmxOGUtOYLOqF0+m4NMX
hiQq8PgAnFoQCw8NX5rZhtShN3BYEO6H5Mt71PjHTyHtxvGKdnqDSTX3jplc/Q0U
RnI81ifTJgOu7ux17psAO9U9DUqy21TjOjB04yJecp/pFs+KMnvWufe/+Y0Wz5WU
stx7Mg9JVn987TKOTXOTkKzJLm5FyLUj7wWFu0TYvmU5YZ7ta8UyZeY0eN0RobZc
EFHwv8cDwxrVmCI5BLZc+Kym+/TwOuFobkV5Ybq3ajDQaD+lWlmP2jxWD4m6OQW7
CHmi9d4ro3TQYbTFbui1uqlPHoX926LkTD+kelfbej5iRTXcs78w88EnNShCCIu/
5V6vnjie1eKrih2VIQxzvcqQXVWS14mMlm0o9jSFodkia38+fZTx4ElGm1ncfONS
y2GSEFWR3bzZ0IYufKpCWOTEfgnlaixqOnWSF6YHCPA3TKaenwQx5LbXz0umdcPR
MEl9lYF/oK/lwisgIHVSdQgoGc/iGY05ICKpajj5qz0EADxjedlXS+ngPrTOYqWF
+N1Hpgb2dchui5J2i7y9CxxbwspRKrdxQYXgzqb5vJLpO1eUoaYoQ4vp4uC8t3FF
WwdFWrO6Q/5wO3lmxRMKyrqn9+new3VrPrJndaKSDPQScbqWo777/juim08OZOgg
2+APBhi3BTe++kZlPRuM6/lpqwJKJ/XmDPUW2FUbqQcqx3xacA22S/zH2g8lJtTL
Er1Wpbrgt/xMWcmOaqdMKNFVOpfSId7SyXEhc1/855KAQMLVvGCljeri0qvltI3k
AYEZHd6LBcqsTlDbW2bxwJ0eeQLwLGggn1r25c4iy1Z7h39FqadwKyiRPRJdKpJK
1qhlTV4ChTraId7YnKcpieVvLDNWIxKt5TiLGxAdcWlMXSWkcmgWH/Z2P1BOejob
NgTxjqQHYfUkJDVrkllxpSyKoheDz4ylI4O3Va2efLFLKxiwalVjd1fzjonVjJIZ
KFpP07mcTftTPD2JmTfWlk0ULmCcquUgmrzMO1Uddu3rnd7A5XS4CLrfl6A89NAY
C5XUm8IV2zp/7OkofI+KJEwRLRluhB86HXEevGpL6PdLnoqEZAzxS9/YVhpb2eui
I/qzFafDjLSsZmayHeNZ+Eg3HftTfP7AXLrIcD5rqxLqcnbLmPj2WLsl/j3+BQt9
p1aSDGEdc1GF4NvukC/S1RaYwMphDCtPBmTi0meT53dAE36bTxvJJLfhlGBC9LEg
ctOYwIsFnbyAEWbCo8wq+uHQDB/VdmqvKqdZ39nGOJ07VgYv0wMP0TXX4ZWSCGLe
bSzETlpTqYhmkadQOXlxdqPUcDGbos/R2TznG4GXHvH7rSw9N3gC25iKWQ5w3yrJ
a4If7QOCTptwS8Selfskj6eYv0XRruL/yM7PFkrZ8ZSSs8uYBH4l+6hAgn2y3OZV
EmOsdW18fbq2IaiZR+gP3etfE0Kn9U6yXWsgAJV8q5JNtVWCmg2Fd0T/7PC+lz/n
edcprO1l3GKHopsU6WAir8YV+wTcGh5XZx3txtd4bHY4lmSSAtgh1dPMBFAkmhHv
HDz5jwxXT2UiQlyl9muCumkzYwVhq35QAa53dNJJovk90xvktBz6kZMIZsSonag7
zxD9w21X2Qv4KvczMkyiq9msKBRqsm6+FCPCTIlHaaOHnsugIBqqefRcU3455jWs
FRkWNoKdjrntO5Xy1UYv0d31lOSe3lrLrJkNctRu7FIdPMjXuQxgeJd3FMwkD2lA
FxhCg4wOjYFQWqbZaVMVNzSiEjew/lGlDBPHf7G5WXdLOMLZ2sFNcvmlWYhB9Uls
s10JkVy4N3Bb0Ln4jtNH1V/K6TDRjbe9DZn8Lx/ak8BtO+d8hy3Fo+DQRtEuSscz
5414OHhqxZutM9sK35or1PPGYp/F+153op7Pd5jVE5KOo/UL86GZJ/ggqHNM5ce6
bt9Gv2vA6lGRtXHkwcSk/xH0lGJIXx5vtZFIcOJAWCPszTeEa14phFQuxYmhJzg0
eIN8NRABYBc+IfaTnXumbLl5EtqarWcUWhU68Kuh25n7ZJqn+haDzUX4CDqRJ0SL
7L3qYHi5BTK1MsEnV5VIqmwsfWaw0BvpSirbBIKwDW9nPnncOaZBZwE1rYxvZ4kc
79u7fD9qFyy/XBz3bh8z2JG0P9VCH/o2hmBeNpgwtnLpXWdPS0GOmzHJpHLCLr9d
XctZMOYNh+dgVow+i1ddZsbzL+naJUwQFMcdkk0wO+36z3PYheylNR/N7ft5JX33
UeUrq6IMTnjp36bP1wy38nDmxz4xrWUzpDpSWPJUBX6WERYtB5xw7TzPMUUHs/HE
mOKfoyJtSVIV5iajUYojUdmacL8vaSmuDR9RQuc7Cc26i8k+Jz1s1HD4Hjy9z/XG
ZRMBYGMhGxVukXfqSG8LQXHlgIj8YhBrLAxD77IWRX7ECwL2spc3kUW3fdtm389w
ScoH33fA5AETFxIkgI0920BTabFHuXgAzWc+Q0m1yNAU2ccw/ZDhmPy9sgKnXtH7
MKkWo1yBxgKwmqfoJr1MXKdDCOZTIeRd3aBT+WdSFxUHzi4qkNTG6kXqDZHwUUSY
oNAuUWYGayFS8Re9Daqvy3NxGi4ANaSI26C9eSBxi06byLCHZB+U8zEK5Ly1x/UK
oimgQnvPAzKYx60K+bbtrBrDv/E1CVJIj7AFT3r7QBcq/WhENwl96KgJQuEuarpF
0vQPeDQNpYWWdsyS3xMknr3HUMSatu4MAk3RQSwIlTi4CB+qK3YzYiEt2r+G7r5x
LBHgN5++1MlVTMjBp5nOhy8xh4Nx675MLHaXjTVcDrnFpBbAMze+pObfdjH3mgVf
9eRK7/sCLixb+neIkTDT/JK27vIH5GQUW5sBBvtTDs/t4tZ0+RRj6oSQEPs78pr8
AzC09HJeWE66RMK4d53QLsKbogmFGWyyLCIzJryOvTD3UVFQGfMGpI99Nif3bXTN
l/gOIPLJdbd/bRQk1TQJtOgTo1naStjr/qEt3c4Sx+/oDdIyyHnVwh5BicuxYnvN
CpznDNH3Cz4AGRFXE0brhtNzk5+52QOHy/KrPE2ntIcFtpVe2rg71Bdakjac3tO0
mMMfb5j4hscV3k6RgYVU33+/66lpxwuOF2HApES2wkeblqsxAVsHDxzg3GWl05Nx
kTrSWgc1xS9WJYVXKDoZ4rfQe8m0kDiksIWG5lp8oxg=

`pragma protect end_protected
