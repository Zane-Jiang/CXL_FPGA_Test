// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
zf7amvhwXlSyp6Q6dl4wYxxQGyrdYf/5JhfmRzOLUTPbh9cBG7FWDJFjQjmTIp0b
WRvnIRTxud9H9ciVmuSy0dGlukQqipr8vyhpBGhUugZf4Rst05+lNRNPbJ9ElzvD
Rxq1mbPwKVyfZwXSqdCshA6YnyI+Pl/53TuOSfASdARhLjTmI9RxfQ==
//pragma protect end_key_block
//pragma protect digest_block
CBtQfYgydOLHG+uIudoJuZ+36jw=
//pragma protect end_digest_block
//pragma protect data_block
GecNNTII/1/R41b5BqTNK3lfAmmNBQKbeMpyYr/QeF4I4LTjCjL3CgD8lXiVxh1Y
do75swyJIlSwJ71jThUZWihtOZDeP73zt09Y9BZQfMxWOXFZ7NsyIg0mXUzH5G/g
u1JSM5AxhtAa9QGv2UbtdKnv5a9rZBOdZ+krYHt6EjB+TZ1lRrabgmpSJdiytHYp
NlVW/SNg60pz0W20p65Yn5DC1+bTXCyjw3IK13jmvXeptxVSfC8kZ7YkcVFFA78p
o3MW3qNbT1wMz147t8f5vjKpVrq05VGtRqbmb+iWxxTPw7yDdnZ8PNEdlrF3x3pz
ykT7aX+xutEtjiOOUaXD/sjW5Ffk0zU2EjhD/0t+0XU2okrwz664nYc6Fst2ZU6W
YM70R13tKwRB0VhtaVQZTVrt3xydWTs3tGDpf7TGGh8QJ80TeLnEf78o3cG5eim/
qfX4vG7A2NnaD2YhGH2+/mfkxvxIxh35YI9CU10D+B+C5xN+YtugbvKBEmEPH0iT
RqowFNR2r8WTXmlPtB/gato7wTHWp+vEtl0QXBXW4InBjn8j1E+sxu/2irRSWYKH
I688W/mwtDvYt3VTYF8oa06REMn+AwuZgqGcA/qsYvZAcDYBQRHWd7oBLvZqET7q
VKW1Y7btAxO5vXAD+85cKWk2BoJhzPD8XJUc7mgrDXESegkofACKvJn4vCzZAvWU
FryQ0wMcwQPjjbPVdqUvyVz0yMfKkoffPwsdoGP9zO8TzzpyMNcVCghCcHTcW31q
krpnrJ9BQl25sXPz+wmQ5AALU1jx5JZT+x7RLAs8+TpqSOcgoCDrZtZsOzaM92KG
ZuD+xUzOugxNYq2JyIm14yykEUBDrqu6bs2Rq5rE+phBXTSySF90g6pN2KowzQXG
4w7W1vGV0ht4QlV5lWULqEbU3rQ5NUpx7/o4pqOhCyyj6a35JqcAboGfgMwoJjvi
WOCaM5avBZETVRod6MZO6KHRBUO7e0cHyT0q2d7RMQWK23Afnz2RiClUK6qHFztt
/z6Lyo/3bon1BpuImEvFpXqQGg7MLrKTmSvKJTHm4OVtxxApxu/1mvWJ0Uvd6mj0
4RfBXm8lQ33dtbfVulig4RtKUoYNR8aB4VUfVosEIB2vWHydyJsD4foAm0syfRHz
PDlV8lsg7CzzI4ozPRbciMpvllnFyD/29UYEDXcPXIe78LbcYUxmibZ9WwmJydjc
qMokVcrfgUcGFcynrYbl473EqmUxbG54OSt2b1SCvTkn3K1KWTg/+HHNreST5Hca
tzCUMIkCLcg8P2X04QbXPMWnph1lTZn2PIlZ8M7JSttqqjvtFPS51fEz+nkEIkcB
XQoZL7ce11sarIZg/EYOnK+HaBBq/WIE+Ix2zT+IIDVJNakdg5g43kzBtLjx2KXK
rfBVN91M5rKVE6XcqTGsj2SI1AHc7CJ+MH0KKjoUTQvXWhL8pmV9YjX1EECcS0m+
iBKiU3vIKl8IVnTcVzl6eiwP5E+y5TZhuoSxgnLa2WrDaVCQ/2YYrr8pW0UjQkiA
5asq4w6do1Qg3VDd2RxIqjmfPeDLhlDZuIdOJURKnBaeKpsgigf5WMpwUN94BtSh
sDdzXwsLBgqmzg670BQud46PsoZ9bzY7yW9Esx55TujSYzjI4/yeM2CNWmF8cok2
vZvm4vejca2++Z66/Iu6uwYegtjYnSjqhRhQinJrt2ElCoKJVULDjx2EtPhH0m9j
WhQ2lUSRcxfTE605hldczbkjSiuw+b3KvIQjkYJJjFj3iV8GtN6Y/NEArbeXclps
pWnNI28l3HNWU9MWW8ymB5Ao8hRZntJeruaeX1yA8x2JW4BDTxbguFOu8YQIKrYu
sD4w1H6dwGPtO64m1KxB5vJ5Mc5QAsoLpfffl40VCdpFzv/8NprqjNbe4Gu5uAfY
VQB70p8L46veFvNZLLj9AltlpTcMqlAId7MtnQET35ryui71o1OfC9crYWQDKC+U
PF/ddtkVOixSKaFbPzGttndF6GnA4wZ0xoqVA/evJd8jUvnuFchammGGCRqrwhu5
EyS28xXJzHWYYSsdIEN5cR7DZuBD5aOgIBAZRiqUVnbYbAia7sCtGI0wIuAtpltg
bzh7T41H9goAGuoY3f739aJXXIBoDXPLVWphh3pEb8kzdS3XsYbBJc2rk7kBmmXr
4+cMFJHbaDuD/fmtuFyF3ViaYE3g5w/9dCnZpeqrsnX3PNomSOrHhLPGhxEZkCFs
zRLfS+rWbZOSaA0sBW2vYrVTkQrTpPAVdzMKlUF+XElbnC6YqF9hGP/UymK5ySIF
+m3jzXH1K3vy/JbxFi4IlAjzioSusgRpztyFKrU/DnK87Vewb1bNZGwFXgFYEbF8
a1ccWH9buO2JFAyfuNUTbdG/jfvnHaoKsfgSZTWgY3oq66oEW8xWiukL9ylewtc+
ZGyf0si3HkGoUASaA8D86+/ztCA/otvy48BykMDtcijCFYq+t2KZE9YLTdneRXZQ
8Ks/erTn+ayehwRv16eFvFA/BZA13C+M6vUCkeDP+Admt4p7j6sRCZU6xM9ZQplj
VgHnqD3YAOU8QU1e0wzPNFBHrDduXCpLpGZiC0A+nwhmgCad6GlO+Ba/2LQw98B6
LO/Qq3Gq3NnHaXEKkstK2+DJmxRMgaafwmx4uIYenVIC7k4+LdNoekjrUVJSN/DC
oRXMQL8JKFXwtqnGBTED4znamj5PuoVVbUzwUGyOQ2Q2SdXvnFILZizcNYW+lLN0
v+j1j1trmiKnwIAaPaSnv0JIQXJ9V0nCTLWtjMrmwusIT3EFclJr9u0hr9eqlb3j
7UqLZPZp0FpOZ6EUwCUogOsOUcNyJoAXSHKAT/XaBpaRoE0ujm6bEvdvgDhpk6Ic
TKGF6SLMwP6tU7NsomQ/sC+dBgsxsH+5fOnchStl/kjIKdPdzSV+9KR/v7OHygHO
uBaTY7XbHjiGKsUIX04dr5TBGzwYBv8bwamPXOTsbjYLECrG5/srRQ/GbfIZXMX1
tkG+mc0PTtls1NZBlWx2n/ninY+AEy9gwOzBfCG5BUC3JHkB5qPlRxwErffJABkW
+DIeFn5grxSMOuQ1uG2COv0xujuy14XP0HlYWxk0P5GnrGLKcIo7EYI7aqyVnR5O
LacUA20swXpKo73E5uHEGPHf9A8wv0ASxguwMs8ymOzJvMHN7J/zSS36yAsmjFam
00LDHX15/DxmQ6sC1RsuaJRXh3/BfrslKlHrJIHna5P92cMmdkGGoC/JYSYlPvyk
L2NnGSHb6l65OLhvneTOl/DFUQRFXJILE1pNSw33HFx8HUWzrBAXFriTxcYNBfhY
PfiYSrfHVPrMBsHOe8Sm387PITuxwbfDlYISGVQDFqKHZN3rrURV8oUfnC3w2zvy
R4rwN4KosrRp1M6UaD8zuouBpnh2pnNmNZ1XpA4ySknYKdeqyfOkzLO7fLE9z5ff
SawSO0zAYH9pQka9sZkrMvra8VeHPhDPwaQjBvsM4Yo3OpFkcvphrYY6CmgFDUvc
s6bvUs11qaj4PutMz63RrcI9wcrIaH+a1jDxSNXHe+4Kxkq3cJWQ4YPBCTIQVgNS
4ypISG0ReCAOzuX9i/EUFktNOTtRljg891DUQrLZ/kQtQtgIjSEHx8ZOWB3qU3jh
8a0ua5JCIoo5VEpDBWpHRFcaFqSyr5Avn8blN76TeicwF4smsCDsKxzNepDmk/GP
cMtnuXTiGAHYL8sQSFVNKA9VSKq0jEzv2LN0d7HRScYgCQD0InPLMCevJf6DWzQn
HQK2+0xIqe/N12YJcx8jLW4Mx2k30rDCfDN+mfX0yNtw/DNCkxfGe2wSBxIzkAJ8
eddcRgNH0t+nWBWnFJE3G95RJ25cf7Cvd9be61LbodMuCqZR9zDZCfdzuRqnIQ1b
ynsFIT/PIIlrS6khzsRSlpiE+y/dWyt15v7nwVXds860ednP9Xp+TgVbi6js69Dd
LwJXuwDhsMrflmTk5qL1jCWqTsU9qEyxCyiidRvUajxIQIAb2b/J4U4JQRAPv0Xz
+yhuPHbxw2/lAtM7swbnkSTcjMmRhBNQLdXfWGcrA3fdIWphVXNgCuRG/Xw2Vi3m
lEoY5iymZI3p/wMJn/+J/ylG0upAMMnNqRVGLmYwp0AHBsmQt5h6N1JDQZ/6LFKS
hfNp8ROitaPTaHBspjSA7VUNH7uM12d4VDN7jX/8lskbYevXmccusIaz72WYqOtM
h6xo/IZbojDKVg7PQIzjOJ0LDmhEa3Yw+jUDTIpALCJmDXRwrOCrG52QwyDIuAOb
DPXhWFDiJ6UDrhPtHmtPa5QtwBjfW1ikNGb5XRA29Octm+oixcEi1zXyxFXukDha
hRTaS8/QAXRwTCa3P0FrtIDcc+5TAf86q6Kk6QTt7+DcEPAmuNoJHPXeQpqYigBq
4ouIkSI8EjPMRSbEvmSQycFcEuIuTOWa2R/b4uV08dV1L61gFwCRdksYQu78IQB6
wsE3fJ2FR0j5x83jj50mTeysModx/itEFiuX5srIijGExjyLxpPBSgyltZkB7MR4
TScaEAotfGY+8/cN5UN+augk6hZVC8jb9VH9CSONfKJFhzts3rnORBpAUx4Dw2wJ
/J19Ekz7tvWYRXRFqfOi+8Z2bkjf/bskskwZO7yz+E1GT7X7rrqD0vCPHWyfBimC
cxITnr9MlYdXumByn4F973F3p7nTlUWo6YAWpEwhZ21vigpZeJBkLckohEhFCj0g
MSb/EZsCcFiRin6jJTPn8eVHb0VWbKe3L+BI4QMNW7tLsQSc+GXKIt9AhgAP+e3J
JVfTCUy7xnfJiV+KoDfFJrT90a5sYrJYR1ceHmCAO4Tb2TtZr6ZOOdzv/Kp195ZD
gXlOLxohWa06M8+dpzFB8SUXFi6IwhSu1DYKdMKct9cxGgOCKvnPHT5klhdD6Sfi
+RcsoL/QB5bOCE5O1N9JCqWy2uqEIs5cVjG7ZdsEF8Gr4w+eNb5zhkjVm7LCX+oC
ckWUplsKnDO1SiKuYnByx2ikqkU71Zx/wQqrsF5RLwXKTk/X8tvFLMBlzEBoKSKX
TH1UmYhobjCaVwPjaf3F2mx8rgAwFAbcq5lUaqUI8g3g0MzBFm3MWhXFJHJ2RobO
fgcQhpufY+tYpMJfHc7mIDis1SFmh3qGIvYZzdYmGAPwzLvn9VasVUAZWysWbE5t
rLudhkXeIKiDPuLWXXN82ZnaXodQQsgDHhuUwIENbRudAhMwCC+As5+8YYmts7JA
1D9o4njOLxGMuDIR4iaZ83cbAMpbtmk2NUwu7pfib9nEhtYJMFAUH3+/2zBNx1qW
ViCTgGtIA2lpXHC/4qK3bKBnKfcBFQxkge80S4nmXnifgmfN1+ppybsF2pNYsgev
9CZrFFOCQz1TRHmSuhqkSXFG+5LhdGTiJG0FpllB4KQNf0QxU/wRx/piKfdAQMku
FNs3Vv4tXbSQJtlqdprR9LUFE7VQNspMhJw/wQJqKYmnTBnTiDXenB8O3yWuPmDx
xsbKNjD0eMwmwy0lxAMCKQo6Qxmsr6/tjNWO97L4nA1mh/4nRYrcNlobuCuYYDOB
FPGWUkCJ6nqbGyKOuajnIoFIXBxuCzh2xSyPxtFFSdcMGfohuTPnVab3kQ0DhuO0
2Q3CihVBYQio47fJYaOxdfLzQCpAU0ah+coflceD38apgV37aslm7TBUU9p4rZTx
9+FzSyFzQO+uuntkG/DjQeAHBUl/y0I3Fxh0xk0D9BKq0QreYcf75/j370YOj+uW
Wh1Awk0DwgldKuLCk2FdOvSyDqsubmbx/PKrIRbuNn+HQPfW0VSmLEvtzzJtlaW4
YPbwdVSf4PJMCzA4EuZQornhjl6grYs6svLjIqaD/HSLriI/rrwCnLcaAtvy9MeO
hOQ0N03vdpJLZX0s1HM3zxEEBMv+nmkgxCpS0mD6/tTjl3ecOlp0KkFSx8Dk7+Co
8C2mBjnLGX4Rvb3ZH1GpkqlpsAUI3BR4SeH5DeXHcFLtxrbp7CM5uDkEAtb2Xbxm
sY6Ujyq3bfaSC02qhzjEVD6SzYiBJNsydnOVCLeWe51iJLYgTAQjBZe9OTqSDAak
7Lhn+8qBWT/a+3UTWMIBPBnVGsxPbVUqmUr8JFB4FBetXRBtc8oQEup6DhgP0bGt
ecZXe042ewz21sXGYDEkpzPibQwyf1EsbRIEgS0y9XgMPKMW9V10kgZFov2nbd42
nu4zu96IjUjbGE1eUIaZxGRk1dp0pCZh5y7wqFx9YEpAPYhnyOAE6UG7hQRw9027
rMizjIvmeW42o/+ydEMQblm6KoGTo6BbPbVONqhh/W9nwSvZOAhdha+zJUCmOvml
17y3yX1++mqcYQBD5UHEymjmuWvLzKfCGHVDBUYKFywM7ePsWKYZ6pTREyeNpIEP
qhX4nNwFoYSH/6oeAbSSJTijeu73LpDnAxbgQEiDvuzZRfqi9n0l+Z71a37hTyl/
M0e2UdbYROUK2YH4aVvBRgmI+2ok4GHouCsk6d2GsOiUzjOWmW/dUz5cMsoULAdS
HVKo33zyTVSpuyekjqVExUexhKTWXnG+Vb2UgLXasoJHYiqJ1DpNX6dNhf8jwvnh
gT8f4GixKsRJNst/xdRNP1DYUt2AxtyCf2spgy9yMbGO2CVS6p/aswo8+J1XAYQV
ny9SPyTExULM/g9/0Zv8CMqDaKJqJLzPIH4oTNnlpG3Q8b36LkJ7/uaK860qYaGN
uqnc1EuU0j+xSHJpSlkD72yfHP+RYl4W70a6PnAakgxhlVTJr1pRrjMZY3Choa+o
qHeajauKpOgRKy1MR3jlaSp7ttxUAtUKssNZP3x3U+G2+OF79Re7PIBb860kPq/T
jB7pe//bg6RcdlPtBrETSDciHVGqe6ClqB9GMJkotS/AobZ3Ad5h2aCOmsDRXxkX
iKPQyLy5GnrGoE7N4yEjff4RrYMWS4f9dOrM5j4BFqoXP5o0oawe99ToUYS9TF08
OFbIe2XpFV7Ycfm8BmYMp83fYmcMkoz1lhMLQgb474dahbYh7o1gupHnehM+7zuj
zdVJ+BjfJyGipMnkFAT9H5mg12tLx4v10H5dslmZn9DPQ3NlOo8Ge2GGdvTN3iYc
oHGm7OnxJ/m7cqnDDSNP8+UVlkehZIj0+zuFtNj/+KgEq4EtgtL3qz1LNH7feoEk
jE29F5GfqTV6g5ctGobJX+9BQAhewc6hVsZxJpWbikyjkiMZc6Ua+nphDkXs1cCy
hn0WPXJxPBWTZrEaZ6gHWCqIEGfNMNGTJ/JjVef8EjUCYVOYBM/IwcMsRjj8DHYJ
N+FVf3o7/uXF5ke/E2spXW++fyLm7ugh02Kj1hpnNcmQd9PttrJuIPRKTiCQZ0dH
Js14Rf5hiuwcY4SQc8rKzBMa5Y1X84sonj1TKdw+bdyx5aCI3UMoKcxMblvlTICT
IDRRNuntLGjzLnvHz/A1ykXR7IhoW8PVALJ2SX1G9A9Da3Gju6kwc7oWQCrA8WyF
yusCu1NttiZWdYswQp48UPryhWcuXHYq/E1dTT/la7nCNvRiFwVafNYRCY08LGW+
/wSPE0gfO4mocUCljR3NUhOp9I+y/1qvbyDa9WQDQ7CIFop5DfTI4Ttf8DKwFo4m
BdWTBFOHXzqh1X/tNzawxp9bHhOWwMgZuOTwswBpJ5me00WzLYaXP2rs2BLnZJ+8
R8iSKT1H59UsEby16bVdmUo6a7l84yvOZp5znXMfh1GgxaoiRMgejaWB1NFqIi5+
hCd2y9M50uMb+BpFMv9weTbogQk+tYfhecgcjEdiPI5TcBGsmHkep7roHGU/9/wt
id/bXuiKWdiRWm7UawRUMovXmZBn58U+LV8NntWRpM+CEBXL7aZV7TkWFqjPsvy9
mvQ1JftUKJs775qmo7O/rNkqxFVacsJCGcIlLr1SMRnwx2SRTrAh0UprPg/kUurY
jUzPuovw6FL11m1mQlFSaoiJj9MH5WuvSN2BDB9E9cXxjhfH0GTLvrXJnIkYlyJ1
MTDpVEtdlp5Drfu0P8n+mJkMXuzu2hRvu4m8ksy2rKxJYQChF6lPa2onFop0wt8F
3f5bcDRMWLFGKXc2IdC7GNGmOdc7xDDNNjj4y1wANhxAi34Heep44JklucgnUJDD
Nzi/nK1tkzXy7jduNx+lsz1wAhT1/e2FX+BW+3pJVSa2IPambBqDMyE6wiRdDuf4
eFKnJyFVJUu8yHOS98kxJp7CpT+IaunLKkoMPA147bK95jMrdiLqo7MEZdPGXWI1
il7Sf6USWkjgn4qGwDA46qa2hgM1Jd5XtqHbCZdxnpvJSj7tCUFUfHO6orM79URW
3PEzgzUMTVKWqKpZhDVOYEwBxZgqTVukCP9vTZOUM3tEaPL9oW6egmDDQ2pDCQrE
xD2904Mn6ujhD+nZa39qdm6IzUIAuup/Is6I37Gq/uvg7XkAXFmbBsJeaEg2agPh
i+MdYZAF+AfFo+mrMKwyDimqUPQGw9zyAOgcsH4voa8wVqR34B0kdwevKYPsU/lt
gyYMblqEEuVFdrWtMYaQk957EO081B8YYkQVlNpUWYc5t6oiouaYRnniiTJE/OOE
PFav9qtfqqpKHDA5OgT1s7uBoXj5IU6o4/8Q/MUxtkPlqFDtgTpj34tM+Z11n7eJ
NEgwzHoqGjfJYvOv9rrQlsQRG5MAnPLfmLmr9EsT70M0nuZ0J+YqikohrcCL6iII
psErB0oI0eRf65YW79nv+svJNWkVUk+zxMCPaW8zzlZZK14EcZ5zGMGBYUlHABFP
gs6aQlB0AOYfpozq3uGqSH/Km9I+dJ5RJY5M14Lt3PaQXeEWuiQKVq7P2CQ4nyiE
Qkktqj4bZzPv2TXNMcWowQEHjptjaPisjkTh/o8m0Y4tG7Z/+EXppqa0nrFWI37f
cLUatov1mzQbgbWh/rkAo4PNR5PWf8hj0EPTjT1V7ChmpAbQfR7/bcg0+leiUHtf
+b0VfWKautJUZ0yRysiYrbfVI4oeyj1YY6Yu0tpE7ZL7P8J9IOd3fSUWFVIHMiDy
K2CBEYBgOc664HMjzz7BC/fLQC8qApg6w3z2w7qS4NYj8gpV8wJTSwIy4nFjwP3w
n/2etwbyz488KExil2UedqJxYKAqueLHrSugMOGVjZ2k4HYjvhyv/73mOZznqDXR
Mol34Fq45IJjCXdfVyrEUYSVPLJrjGOCh5SOtEeJS1AHNMbO43gr3oJjafNlmqXH
slXKVVfNcDwO59BEfy6l40UksM114FHHDkT/50uctjlbr5dKuP3r+FKOgQZm4AaZ
YQR0yOQ0J0rzye2Z915O91KDjhUpuzJENb63hkSVyws8CYTHYnxGPrxY7FnU9pur
5JMxdEHEdRizL44LiolagNH+ExvQ0Rtj0DtM6LUhn0S7vmGoCtWblM+WDcujesOU
igswl0I1uIn1nxJyZpBQVVUwart6MuGDDr9TvQYi1q6rud9uNDG3KVEs1Zr2qlxZ
4qWzK6v0Ra2DceOdmfh2qip/f80u/RpnuvttovCmDgcHtQRa79wbKaZj/XyCubK4
ujw/jxkQxod3M+EGlOvMJAOr4pSu4r8/3OvQIYCu5RBrf5tsyiNHAsQ31G6sXK/m
M3Ui6q5Nul1vJUm1vEXH+qMj0GEYIPPHgWDOHXar45vgaSCeFyG+UdlclCU/mnr5
9hG+9i3wGCaisBf6s4OV4MtbKdFPqrkVmRFi6hw+UNr/aulkFRlbYAdhr0BRf3+1
NnzegEgikKzFHjUmW24bF7dccfehMF8+TK3c3q9ZmlUyaHPDzTX3GV/hQ/fE0/4k
JMUZJKsk3SmUOk3yh6ai7fb1aUJ0pyuoDYHISYW0LOo4Ee3pJE16pBAvdHkNqKng
i1Fck46YmUMZ8BAQqM/paUaCct9BkZ0LXAW/ArSgte4yrh9dRaKCXQLr6jtbldjv
0odusbmgJumNGB64/h1LWCHjw8RSQTkkxmX4bSiDlPZhGfYJu2kEAwmAjCJrJ9j2
5LyPDJrXPvp6oPdSLeTGVShAIJ1/jnq8ev0bSnhJcEA+Za6TNi/B5IiTplrnuAJx
FK3MSbE9Wqu4RqoLZ5Tg5m4b79qXmC9Tr4KhDxFvF7+IC6z7p5wz2FPv+4ixrR5X
gR+4EFu7GK47MfVJRKYWUU6clER2nEnzNEoflUuyBJ6Vrr21dtTpxxCfTDjmN8Ut
aSsxEOO1Ru/gybGkX/HvkPbAPPznBM5w3CLACEnP0yALb+/M+v/hYa0RcBIOcgWP
n+O0d9hh82sJxRAgiPqZHY9jN798E1EUWuKwwUGINp4KC6wW6ddTmi9c83spKOoK
VvTqMDuEEuF9DaRmn1/L1LpMtVchYjcYrYYuQ6AlhkF+3IPn5QhxYukUcoNcbNew
v3NbjVS6Xk03lz9xIwXwMmr2h4hF+/CgDFxYDvQGgeERZ+vDkIhy9H0gRY/5iTIw
2zfjIhUznw4gRXXINvjp2q7WFZb+YKaXYLIO8W0WpIXs3lKLhhdOs3I9oAA5ai4o
TgczX7/iyXXg5iZcCp1Ehu1jBVtNcUT3KFc9ufDxNzzvJBCFIAOzlE8Vf/aCTDct
vVuOokEBC4wpUEfeFb8kGUjAtGY7pBgA7Cwtdc3hsymTroaeYw1RINT71Nk5BweX
Fcxs7YI6f8BaCqDUnDZyjaSR9XdKX9sP/E41aScKQykAil9sLYJrTmORjGrdl6r7
DpRDjuH4C7jFP0QSlRn5eKuft5m4EaNBsJnnpgPcWbPN6Ku1YNjad5Yv1/zDmdBo
zj8MA5B8eijYHDc+kDCrdFoqDvbFygLP+/Vb0TThveXanrWzC9o0Nb6U7aXMBrDJ
t+qx0/ROy1V58/wySgrMeg37BM+mXHlOK4889kkV1aL9p8axqr8ySYT4HdwWXo1B
INHENZ9Vj8UdL3gIxyZaA9TM6Ftybv2O9g1XRMPH3vfmLUHo88oIAZ5e0DSmdz7Q
uznolNVSEfvMH3Wn/4Ms1GWiAvNbeLPdHeotBpNfLZiv3/q1fmRRH5uME6drgdK8
Rt68I6vz2WOGgMDlVpr/29/MEP1xMIxPcypbAlcVaIcXj7b/a0//4+5VR2rxAC4T
5LC1fPvMoc2soElfB/q/e3a/FNswXRlgz4x73NoeaT+IklkDJeROaHujncgHCrtL
LxmGyL7rOsRLRiKLSO9+Pc/2jtvHkxfVs09RFHwsXFLhzptDXj+ICcCtc/MTFGbP
FEUQyoqrgQsfDUQl9kT+C0kTMb+ZqeVJZlMbCSBEFAaD1/oSy7aRoYFGqqoeGO7r
6jja7LehZnYcPrtTa6G154JrNVv+Y+8Np2sEM0wcSYIQzd8zJERRW2p44RNaK5YV
IkPK5/uQFYpqayBHlXT2BSPVTcrR9cfehxxCbHI9xtR8cJQJqx16i+UwRv0kfXyE
7c3WqBDXN7WJcvtWV1YMR2et4Wh3FxtAtJr9poU8U/bIDxTryJJotZJ/HcZ5I0bf
nAGSaKpHnRvFlW5Aueo1+MoVELB0mqAyy5WD8YATEJpFPLjXoMcRWP0fsSGRgRYw
Ajeb9plo8LgG6AgZxCv+jk1nvvfGTha6LqpBQMmU8oUwDj3QUFF/lw+gec+QC59w
wTjrBEVfEIuYF9WIuIt+VaM4FhdMu9nxb2zk57HVAeyRsmNEjXw2zXA+uVWGFUl+
VS17mZf8NYGQ8ZN6apaLB5FOCn2lNpX9m0EcBWimzVV/CU84r+OrnAOBHO2rNCjN
5bHDhv2QdcLdJDxc1U8UxM+CKRJ85NpeIXsBA7lu3KK8xrdHmNSvnl+UlFBpaYoM
YaH6pwj9y+e/qxcOMfYm3cObIOPBpfkm/uQANzQZf1dlMhsU4R9Rz2ZQKsOy77Bi
nwv+xemYtn4Z7FqPOEu289Be+kQTtmgjt68rfNtXmvbQmxjdS0g4091L3aiixvro
BKOn+orXp6nNO3ADI+OfU7DFCbEEaec6OiGdssvHvbRVZoCs0OK23E/uXFYAYtQC
H73r9oSd5Q3wOTk/yfsJFXcfrTLbdr1NipknZwvemo4XVbnJzdSKmxIuLq5jItkd
N6TuJGCjbLDJWAwX2WnunSdAf9dur8E7YKoG3PAr3gylK0TOaTwZtSY6i6iMrj1b
iViiLVvlKRWxnoRfb4vygBsOwWs2EJpWhdyrk9eEdg5PjlSTakR1IzzC4Euc1zXx
1vEsUcxb2VCyp4CBRtVWtUBDnyWdRgsrAoOGniQoyf5mPc7yZtjMtSsNOCGoZjQN
7abxTdKXBq1ieyiId3kf8PoLVFkstvAuPOtlKNYaJ74DnrQkEiVSXXNsysYukTly
6ENHp4zQfUtRRwKSSy6Pgj0M7SZNfBs+XIVZu1yaDktCDagUgTXiBbuuMc/Oqvrs
oJCnvC4d4Yaf4+bmlO2bZIk7I3o0y1/PlSEr00MXXAzE2ZfmvEDXvesS5fUfC9ES
YhajJnLsNNJvqkPJh0FnhBJCZK75i9bbWWKkHEddUnWTBM9FxJyoP1+ycTpDjwih
TDexRhoUGq7fDO7LZUlCVU4RiGPgURccUIWlbKX2kqMtHje7kY79/wyXnzsZGuU4
U6U3t2tri87/1uQfI2ibKX2umtYTp10y7ZfEzG/KgSRVcMHhAYOydvtA3kBZmsqr
In7GgeLFOYOJNqyif8tBDP4pTGMZIAVwXaVb1tW4/Qs1MtgJjk6nVJZxm+BXB+PM
ab8WTdid9QUqJvHtBl5ZmcNWDRNBYY13tbbCIkMLX6Y05niPmvX/9VhInIt5UQn/
K7SqQpIvwlPMXy9ynJ3fVvsBEV+NJmy8kM2QEfxv65HJIx7SIYgHA0SZkIhsK5tg
YZxqkc9agTF+rRQDCO9i1g8v75C1azgbLL9HCfkE+Zk+2PSXJAuoDDTeqGbYmv+M
M831in9QWAUgc5zwYFs96v8RYsJfnkfwfpwEz5vbsFQ5OtEjrpi9EBYSZ1Hv7d9k
mTc0a7IfYdAJ5giCc56dy8kGoyVMhQYZ8YbPBTiDNkOPmpjcL0mmqmUHkA7zxe69
fM9moLvhBXglgecGv2tcwtc8cSNH58QJUNOZLQATOSbee4H2XIAP9i6rZUdz+v6u
f1vJuFTNnVYWrSWdcgTAqXAH7AN39o220kbF0CWCraJ4ytcUyFKf5k1mQ1k6BvUw
7wR4iwNc9Uk1MRvKRR0S6nlNJQObu972MREDmVXTIUp8we/8Hyy/qZTkd8FgqtDB
sF38QsoEaLw7nQVzGB5M3N7ILM1fpkFHzTx7+Gw1tVWIKRYElPYHttEVw85WrtcN
4Rq2ls363KZxI5l7y63tU4zFra+URRGKQ8wGFJ0SRuHFt3TNMq042gK1yhX/q31N
uyA9Gtp+VWIY2WaTcWPoOyaQ1ry++q6AbhR+FzXZvMkQWQlrUCUhPSx77NO+ZKUo
ET+1GNhM4c+DFEdApmQyJPpxgqiTH+W1qyKW98tvHJrrSvXCrpBfx12Zw702TBr/
xGxUDyVy8nImFzhv1oJ+DelX9b6yvSnnxxYyprpiAPe9Rac/DTwheXMz4OG8Fi52
r8DtcjW+yezJB2ol2aVrM4nkb8cjneMjxXWNnKJal90dXpZN3jUNR6aGvwKhfU7m
WK7mivL668sCRxDF9JTa/4sgI+w5k+28J38NITq1GMG9095q8Ghy2sWcURvwHPjE
r3JsrEzCbO8JSPVAGGFw84VzTzCuIC+AinXOrowEqM3i87YcgLkjn4EaXkhJXpcj
6T842mp1+I7QIAvBBO8xxlyQDT+8QpPLIVtSu1n30Rq+BzVnVRbHS6/Fc36AQ9gV
Cc3sAffD/Ltg8A42xEflobbD/dGeNrP5BQP541Umhf2JHlKtYigAKiZOJfQNobkT
oNVJVSr8nDOTDrHja5k4+muznUzvbSNRfb3kYdAHaP/XQgHi2QMcJM23h8petVwt
B9/XwzFoCtr8CzlsDu5adSpklc3GUGStAkT2ca/aJNcct7/e7Gc2BPQGu3JYQ722
K0RuxS+9LmhuPj6IWPJ5MUtevDKlZKimO3EjT+h3LDZQXutj+NZE/VU56ZB4hh8f
w7M/xNst/W7q3MzuRucuZ1SaRJvRFMxW7XCJN4xRUWTWjqgBhNyho72v+cLdRyDZ
BMbA/4ztgbb4O4Cqzy9bZs65fckhIgflFeR8py1YLer7U4sSUYrUUoz/F+U2JmED
7lFYWqYavwocm/ILN8ITu1QKLm86yOKaESJd+yIxunXqdw65Fd+YXgPLnB80qOqe
DOUNsqHqL7avf9Pyi8xPFpmaWaBh2J16Wo87gP4qFoX3VAYukoftWNn++huFbyre
FQNmRv41GQFyfrXNqHOcTUwfY/2O2uu6JUHJvyIaw+TcEHJ4Sg7jzAeZOQ1Ss5wx
Hh5k3BgXoawsGmbcjPyd7e6qDEtXxsvbepQ9tXb5BNmBJzfnmZttoVN0V87e/z8u
jNXjMBZEeNcLa/4ZBk+fnDhPBox1XQh3QQg+2u8MHG6QEFbbFh+7/rtKiSuthXlQ
2iPJowFFCq5Rv+ePCwpRH56qRQ7FEh9qTTyVh9yNHmskkpa7A0wQGAF6W7D1p7VF
8hfGd/dWCfV5YQ+1kyO4aV8mq8vS7xbMTgKdMM4XX0pO3hvHLU37xf2tUmNgrjpa
k6gp2ilbF/l28eR/jsBu26Tn0UzJ5U4eqlM0HPfguZ4UNvH5jNvCRHCj0E0Tcb4l
Uzp+g7p7s01N6yV4AqcFhtvTcHYqqzXEJZLpqH5jYXQYJXVkVMwqwSkU1dxdtch9
c7+QOg8ZYpMmCr3cBTdfiPgbTbaetJiu32Sur5f02yGtOjrlIh26HMqq63nuWbFV
vosAYyjNIZiTqXQkAGQRIc5t7VGLJ0w3HYgvc40zsLeuXLekNUP9kw9XHSAycYyO
3lCZ4p2Ch3UHNYrb8clgtidAoos4LQSUS5hD08KCJXHffneEfqWde/9MJnlMmZ+u
yQfLRl+XEhT8hZ+5vuAeHhD5BuWh9g07brcrfwnod1GtO9kQiSU/9dl8Z50WTlmo
8CbCN6h7xiSsz/vZNzvZ1uTyb1UwTA+S9R6UdqQpqDJNhCUrmhNRLq7RqTJuL28L
r2nrpqYOGSfNLf4cXr9JYYRZWWplvmUMj05hxFr9vrrHsm9nH1CUMW2SV2XpTozJ
zuVW0PNDAZVFjVgQqyYNWnw+bNzMZKYAF2Tz0x8vtdpJFqiwavQWQQeKgJP+ISHs
W/AU/9XI9xgv44tAnJG9AlJsicA8cexd993MEcBBQXNXCjk4L/xSQb59W/ES86lk
wOOEW/1TCXD5ln+ukMtx8Cv6/Ex0km+y976s3alU0PEzMVAtIP1p5k4frPo3j7JY
j/P5D/AeaUu6PzxRt9sK2IDLKAXTWLB55NpJh1mcBNm25dSbLDQTfjo1ZjVegwoK
E7tUl1HTJ1lgAHtvQAeDtCCeehA0UbJQ34lbFiwS948P5TczBxArjdUCdrpTqdSO
4ygxBdT0+k1Reks212J0K+ro5H1wTSGZ5bavrG0XvHyEbArsliOmS7VFwV+/AXOR
ELsou0+MQF+D8q76rgOgoGcIZJu19358TLBc5whmd7jFkYF7evD5AzD/2TMNKkKn
VEap0WGhqz++roL8af/QvrN0SSgY4PeyY2B1DIvaC6kWLA0LU4vIcBtxC5BfkztE
Xl7c7nBOh7csOx/lsdS80n70nIPrOHBsqXTwG+0sX+6f6QVqG4bY2Q+JEryGYOzU
/uVzF4/NylAymkVwgoM9FHjm1uVfzAcBuAQ3ey5u9foXBMx+XFMRkl6fdf//BlBy
nq32XzqumMwtnuU1P6pXFqqGw4+L83HwvEfFIuVX1wfvVDbI7zpag5jRo6xnseUM
51vL57S76WiYl6yuPZJm2dTIrY9XH5pxTozycpAa6GynNjNOcSn2Xq/D4K6/u++g
B29ON4pW0U8ExRvT224Qm/3C8FUhTfz7JBPb7uH0DQy1qwfF7/bfxb9DNzUWZ54F
rklgqhnkOnBxkQj4kvfyfl6xuV5EaODt47GmTIENU46/yVXuNlO9R2IUwdqu3Wbg
GwAHcHMwgRJLo/puEamRchAXJYp28EJVctYs8dfV4YjxxJ+2DX6UESY63/n97vMU
aL3cXHUBvqFdaQpwDOlN9v6nR5Qd7kLw4Sz41fsKJPVbmHdIdWaZXbr86SB82jqU
EpMh9Zsk9Xac+PdCckMLaw8exR2fAP3grFHkeopoNPs5hct44ip0YRd5Eq6nDLWs
dzwPwiIiCMlyw/WOhO+35KUtZaM2DPB+PPkyFogXTBxBYKKNj9bOwA2c/3t9BAJP
4UHZGeVa3C/StaujMKDZYvmX5lOCtV/8vmIfCiHsfATdFY4cjTxTBW3p+JqZ/RWu
r5ZztBvx8U8lZYZF+Irqhk4y14fkhsSdXPNoVAb3fFNFU+wRtOO+Myq08XnDSzse
c9kQwWvC6BXWzI1bERZ9DdDG85UX7cIgp4GidWXvtbV1vA/6t0dWKePAaUC6hU5/
oMzdxihH8cfnK6rSuLN9Iu7F0z7cqLE4PB2c1F/BQjCk1z4mJT1vx45Hx+hXUBnr
SPunS0TutRNcBu7F5PFiXbHUWiOi9ZEcpuM5hQ8Nh2WzbV7zsUlBPIFtbUs/BRx2
c1pkz27mPwmoCIEj0AxDIJFWl/e2M+Oo/Sif7b+KIwM8gNW3/D8IUM7aqdHT7F2V
L1SdsvZMqZZFxg/cGz2woMqvetOMIqlm6gsNiZJHTl3exUZSUh56YZ27Npa03xpl
0Yz64PlipY7xNpQNzy3jTGJ1OAYzK+CKQeT2WmQJZfVwT/heOQo7rLr7E/BIyKwW
5xvFRpz7r5X1RAkFUxEPdNisBCpC4LVeidrtYNnIaGHcFXUi7rjo7IHR3M72VbKW
+f8kpFRknB9hcf4f3vLp5zTCd6S1tDaw/lJc4j038OSkbmUS5lvaD62Kz/3j9BKu
hTYCiG6h8Y2E+e4KqCR6BPm3KqZ/niy2uhcQgrXUV1hTFCLBr3m5RE0GZKSczYNC
74Fr5NexCywIBXhNuE8pXtT9dywahhfEcyv4Nv+2+87pOuJNN1c7754Ip2hdmLpe
1fwjs5xvFgprC1p28vGGsNRoBM2w+CNOwzHDTFw9c0WDc6CZyZZMsx2IoZiJeC3H
SlQbPfdhsB1vmFoCzqmbN/EfjrLywxBm08GUnKswY25OHokmvw3ec/bBUuVM9I0c
9rKROljPIjEEgh3/6o4Q6KbENF8bM6fp92WYi8Kh16hmUMMRVGC/w+6ltzidH3a1
i/hudBYXTK4p5hOcF97lwAMosFuTqfP6onQQGfb06LJy2LIUss+euZ+yCEpz8S81
DfOfALZHHVD8WVU2G64GpT0do66MokKhOqnoD+4/TmLXK7B46aSAqEkMGPTezepH
nCDqZAuLoUkS2thyyePb/pXIak6ouBhs9rPHLGlkVbKFcBHEOZDxsMBQL39W5WR9
uDi300yWMJZ65p5zjhPYOrC6XW6/wUU6NIY7pjZEtrd5+phXG8+GONVc9zuYRWT7
1uODaRfj8KEZxGqmHy3nJ96gSGSd2QqnnvUFbLL9bQgPq3j7YvusBr2otm8xKeH0
k/BdrSlV3ymRDNqnvjIHX5lo5iDNAgbrrJGydUhAXeL+KjEGVbjutsZ5N55A74Ey
qGInCuk8dNAtveLf+UQg9j7A0uO8iqONhS/BaOgxCtGOQhtfOW8/1cTW/2j1dVnm
l0EpOGL5BGHxyHygiPEh2wVRJVAH3PTG+LaqRTNlQLwSNs2Y2sa7E0wTq6YK8dc8
xVG2xjZc+dxlcNdfP8vmUcNiYlZ7BNO3rcaYaDpagG1eURpWnvKzVeqSJ6JTb0zM
xokd/HGOqgad/zff4W1+mbAj6P9bHnEOV/xsX2tgtvgfnwBDduvMIDFzlW4pdC71
+BHRXRhLJ+ujPbeb0j/XJLftXf864tmkT/W73gH3j3aiPkqwHCP7YIYdT4K3SbcZ
mjEelIQzRB7Co5CehE/mbVcQ0uB7s5I1Z+nx4pR3Fs/cfL7vmS747HKa3sRI5M2Y
f2+B4UROKAQ/oOKQaY9FMacr9PBkpefYKg2lg9ur6LO/BGkZk8J5yxyTNHSjCaGK
QVXxqjTVcRF9wjX1e/g6Kx6PFKNjEMahMIgLPcQyjETAUlzXUhIJaCkmhlFHrDpV
+XFCiHAJ/dzW3qpWGgt42Rxe9XZV8WfrTCc4sbpQej9kfoBFOgaKTGq1mlQQoXsQ
KCD80XDHerwXGsermyOWFMLssNsiWmndNfFM1b98bLqh2lxmtm4JhqfpM+Vs2Ioj
lYuLi/il9IUlf0W/ckr2QpAdFB9o1j+ipBXYwNRmyrlLoBwRTgf/16b3j/zIelcV
SAXTTt/8aZ7ceCKp8HHP9z3wGkFA9tXFJ2ZwctLOuGSK9BIl3+FBRePx8CNR1zFA
4b+3dKIlvug17xI6V7c/tpsnACswFFgeej+vaK30A0Tiw3mesmbvGTMzfL15+i2m
8mEpCinihV8E7+Dl+RoEwaxiqdTbb6WxnwngQZMCMpDnniqbM2v8Yf7HKzpXWmA7
H9nPacmmRcqY1Ol7aJ+suzZHt97nfWYNqzhnpeg7loNlX17NL6GkpDAafISjp6MU
zfVs4gIDmE+NqqyKXRVCTcwuHDiNwG6q1QiqZxY3R6hDldoWfEYUk8QMClJpb40V
x9WWL2idVsi2eDLLuCffxBGKaN6YDCZ0HfuJMNPxPjeHvr27FB7sRNO/GesbhNkR
MSaDrXFLnvnNoXgMAJ+Mb7MZCx5GClMqCAgNqy0Io8Q7kouH9DrsPZ/7O3+4C26M
k2AuGT9uDsQUnTWghE9gQ8v1YC7BQLAaFKOA+fR0upippFO+Q4uKH/SqHH/51Woe
g88Gp/8ccdCfAWjvpsYeTyFxc8hoRA7r2n9fb2Fod7AsGtCE4z1xfks3/8aIVKVo
T8M7KaVmVfagfzG5H2SfyJvxkiV/TiP/y1xQcrKJ7MevY9V7BRkiBXU79A+lZZyx
5mpp6mvY8MMHopeOd+QpnmMDA25gX8WBw6wyvNfALkcz8LhR98CNLwNoBiv4hz5j
bfVToU/sInTKuNHAlHayUV/LWfVWossAssk9XMUGXmcau9eQB/qoVTZFDP50+b8J
SSZfnPz7fZ5udIY11gKA2J/xYc0yG6xJGU4DD33+AHtb5E8GnfZ8ZkljGjD5PHlA
EERYBc0tFZG8yt7e+Vl5/n0IgN0hKDCOVh0aPlHDio5th1B6fVw/1qU/BNB0WRBT
rnqnyADRcawb0LUVDHUFW67wrNUF7HYuomkaIbZNq1WUno5F1aYV8Wjx/IdaIE/1
ZeuecT2z6Z5Cq+iX+BQsW/+8A03WIrIdt9n2gWpw6VgoH2wn/fPoA98Z2GghZDRO
oBtme743jeYyXAD836Eqzuk1EIGnTJX5FArrhCfA6QzcvtcFzqMOB2qqpvVrLiim
XUt/EDD8t2y5z9VfE4/dkFhpCL9zFso5vVIa2z9f+SeSvmbD/UGdvRGh8A5iXdkP
vMnrbVO/8ayNL2uk0A50zwUp+u9HvrObGlgWs/JYIU/MsqZjOVDR0Pz2GOG7j915
Td8sLut59efcgmRu0cDK63gCFJSU+RdN0x8XkI69zVmpjtk1MSMSzXBq8bEdL4BN
Z6u+78QmHZfCUevNLImW1yzAlRzhyCkZbqq8ErggsDnR03fL46Yy4PLlordLvjnD
GMdZyyI3fJ3/ddjwUlsNk7fY4PnHhmbgkgMSJrSsjXy3mT2qtTWY2pIYZ9lPy4v/
9MwxaSDorjt/znw3ySZOQhKFXp7+ZhbLEezrlT+inSYNN7lUoLbyzMYKiv4a3qAZ
Gx7ZhAfrbblXuuJxxO8oq0Vbs/ejRZkM5anaMv35EvwWfvGmPz1uUqNx9+vnjIo8
yCZx+4BP/RM6Ihi9aFRyFsqeg6HMfnR7Yc4zBNCq1mnOjjwmlhB88DCS7Qj6cs65
o1axD7p2kivN8FC4Y8P1V5QiNVbcOydTKzhWK1qw8UbaMnxuEF1u3nl1w9ylb1+G
57hSy2GGh1CvpYTJTTC20yPC501LpGAKPya+tzBCN+wv1FoLTXuxhXB+faELOplC
zBSGLJkOrsJTLbJVx1Q/mQRCyV5MShtOVdLNZn5Mm9HRPWOXUqdN91ecxYiS6ljX
gOvnv1bK89/u2eCChjifI0V5B4antgimU+aoJamGP00iqBVg+nvojvpGJu2UsHIS
rU0VQ5NKy87GwJ/jnmVGEjVMTh7VyjV4V/TBLT1vdAHYlBo6LOwy7eGSaiSlA/hO
h4IkdaSwHMQDMaekaBP9jeujWjxBSEAeGHgyWs9cmZg/+FXnwkPKImTVfXhIt0I0
0rHWludrUVgtA/RN6WqyadDRdEykz5v4klqCmyQBFLWIki31HkMRy2tIQ1e1JLg7
AFmm3yy5KzXdi2lHdM2NCEUv+goDwWqKnZvsMD2lJHPhNmCoxGblLegIkF7v0koJ
7/0+yPqDNslp2MB6RQlv6Qh/ts4x3EzIWJKQr7n4hy165irZD079qQNM3zimBT8c
GmtxMOh2zQJE2LJDcLx2EjryhMj3pyDV/d0TOwUJV8ze+kkZZh/NT3TA1zIvXfhV
t2cJtBB8orNzK+4wJPERhYTV/qUPMrL5Wwl0TFexEi3eQvh3feNRer3P656qHixD
4BtvqkioHL/OuNvbFFbT1gM3x1L2wFhB3wzBs13Br0dLWAKNrKw4JW5R+YEltBpO
PDOxOWKWwrnYETtGnL9y07Th+HKEikBLDBmUJ/SWcNhxwNAgJnB/TfgZXXOcAhsS
pVSmXeps/nKG9v4QxyqHJULMhaTqB9TXftuQB91PNyjkqlGIUaDlarSqLHOqJ18+
bJn/U6ETGrscTYCqAhDtkPaRrEemmHcQTz0NqJHvMGKm9tlkLNwbxhdmTRJcX2AY
qGbSxoQnLDpiQQGa43HtUpgasbPFXQffSs2AJZQOxdlRBhGnPVAQMEcaFqnIdXC3
P0gGu9F0eXGdL1uKQh28bI/YbtN1XnB20R4sD/usgK3Vry8mcLyNyoS7ai9wmN+W
ahG91w3uP/PQkvm0Id5Jn4AcAw3TbC87GmpIPWROYDxvfxB6+qiqdbWisfjNyrOQ
7saOGhyuDeMarEuzu3PcpRwlC7qkMX4j4v2PGdW61iBDvNib8H7hIOlV9fCvRMWj
LnPVTHWxR6tJpIDESaKsrPAcOV0NYvXH0ok7wgOaJh8FUIHtxO7WIQaf2LKgJHBk
VjEghGd2w/S7gWGXT/sXiihS7N/zcwDVx4TEdoDU59qNYdQPZOxkuQYPwSY0LSnq
tsrclwfeohICa1jPXW0nvNmUyeP50RVtCO4AR9Ky/dDnYTaBPvXmzMaNSO3+tKRH
KuYw5Qyq5X552Is/DwbuNg33oLkOvrDMFqGwzTnlx43Gx39CPkdpoIy8z+ll03+z
VirEbp6Q7SlHaTF2PJMntnOTTb9ud0ARfY4GOI9Kansr524Cs3B7AmBqoePPVxng
gWna9Ruh5EG3m/I+8u4dmi6VXapJzxqa8eOnDMmAkXLBEmqOSNwXaOEEhjJjjflC
ujHeJwwD5RIE3442AEirlkszCqXxknlxQh5J9Q31zdNSPw4ecairXGCjHAKU5D4T
hL45Ka0+BNSTX4uJ28+7GcKg6Y6PCLxYFn7Hr3DESFU08JECRL6q1tu3OC1qmT0d
m2c4s3q49A9UQlqd85VNdAFOTxbLPecBYq1oBm+rDG58tf0dib6+pdXA9uuv51ik
PlIemSKLnBEJtnWE1Bex+ZGd5/rRuArl6uSQDZRzRylT3AhDylszhDbcyACpCdHk
uOP3198QtZS8XnVdUD53mG2V3Et6vbFtDidqwgcr/Y60fek4kRZDMW+Fim26KSwG
H8hrXOvF/a5i8B0KoAMx2FmNI6FK9Vd6Erm8LvQsBhZzc6EaHdkgnzEuhKuloQXQ
RAYS8/2XE7garBYffzc2NmxR5L+KohUbYdyT//ztnvCUaFX4aYNjWd/pdUbalgUD
9YkUsj4jycWDhaI1F6Zaw4Nw2YHcBQvo/x8va/g01sVgaXOF5iYIbn8MIHMe+N0W
jnSpbIpqWwRbMYB3eBGcrbyOdRDsa0wfd4J28EVqpGISS1B8Wu5poVjMDrlsgJdC
UjGV4U84r6zUROHbVU+UT7nTDGeUFslOegXvcawha+ikFZqZCqlOLxkGapQr5ieK
CLcqViYRefjVkatGDKoovj93yF78Z/IV9l/5QPfASLFz2MdkopHisKvQs4q+2n4h
3pKSEjjnlDqL2k8RF8d2HqYDqy940G3DJ95Krc+uJ3Yiuj3uZrrX68Hzuxpml/bc
3uhpev3LI8g/9RhMsG7RUwlOmH4lylGIrVQQDy0Fl+cLcWQ1kEZyi+e7leSVoMVf
NBzGwcZEb2UYIWQoHUBlVEi7lex2JSzcYJrEg4AP3SJIHr8Cm97iCWjHUdk+9Ihg
bgM0VC9Je3zHNzC8D1Q6hh9asVPBKzU7VFMXsq3RTtuJRq3teENvREoXmnZsCVfU
VeVB/Hi2lMeZt0++NhCeAU5/DYG1bRGYDzOaMJ4+CgKOAQYekEw7447hijiBze7O
2U/Ergnu6p9q5nybqoYEpUWhK9DmWYMg1miD73xK0A49/GqRN7VX3vOE87yfspWv
wJbZ2XNqytNqblTjiz2vYBJn09erfsYhUvIaoiKCBYhRX6ZKmwavhTOO2UveiyY/
OPVmDNZoU66xHzBm9f+jSqXpFliwquBPD48sX2T+bP+dlDEUUo9ABBUCKpyW46zy
HHt+vuE+Z0QvLbmqVJD0Uu+pw8ZVpP8RGBU2+PUNneXtyrNx4mFu891ExRBFCz+6
aQfGhImOkYA+vD7iplS9IOmE6/e/OmFZY/yBTdcVj5VACm5h81PY0HpKJxzM5ztv
ZOA9enQq+tETodTgRqjeI6BG7lCfCZJctmw20Z0pciKwZHtJgfuJchugq0/bcNR6
jq8fy20cG0Q1daQ1Fstbmcqtal71slcbfNszBtIvFxyvWatuLVdlA/dDwIMhCgs+
5nY8SQdUgS6feNQMAdbslLnOceodlytuNK3RT+YjfAk2JgAZXosqGDH9n6WX+TIw
6f5ogtA7dC82gUh32lW+znanZWK5ZNHqeQE+a/+OF250CljCqhCj6tdKrRi/0X4K
+PddF8FJ+a59KMFN+COsh7AyGmac0ntpPFzlEHDDCohdns4kKfZmCyfqQPDPKXmn
o2GRnkoLpsSZbgLqL6c5WIXS9r5lVnj6yB7kTe3Fzs2Ktus01QVqUGYPKBmr8To/
+MXp4qnanBEPx3JKIMWkVM0F8ukyO6Auf+gp7HlhNNqiNrRrTjLMK+KB6MzOH/a7
UJ3/H1C+2jI4siHntpPjpDPXFhLnFHEh2dM7apV+hU/bIiGP7idwcfM6Xv+yDDkv
tzA4V6XE4T4gslzZaKWeZjUP0Jf2qaedCXnjz5WoQ26lHrtNmT2k9oAFnScoeSyO
lTJhcRh8jze3A8ZlRnXYfbqrsklu0Qj5BUbN9TX+DceMy7MrMXIFq9PGQwDYPris
I4e8ZMzxxK8656zSo2enVdvDAAjJIciHRbIPiIhY53x0d8GEoqleZrg7K8FTF1qN
Ac2G/4vcseLKA/GDIP9ri3jivo9sOnmSbaV+D41Wq35BkZvtkQy+ZOxvW/iPrs4B
fIO5xfk1pumhSFfsQ/iT9CthdhWoWC3b73zYDBRCoZYvceoWBu0ZifxsDAF69p/1
a8KR0+pXAsiiZP8hf6Cm4VEKD6mmsSrkUUq7LJ4cpUFTqZPexssN3Ch1km1b0+ZV
Wk8vrrBn6vLq2Jy3zhhvWS00r3h5vrp/qqK0ZgOJSOU53s4uArHO3SH3hn2l3vux
IT8CVFbrom++7VUNiN3/ceg4VSFd0faOQKwz79evlFpk6Nnffq5VHWN7zarbF9bd
MLlp3OzR93u8d4zbCCfgEk2AysWExqQkzp9LyMdI3kFj3VdLi9xbgZm3Cn8C7DZf
UlypEuTXoS+CpbjL2SFmVejFfyfFJgANpuM10GjbEbAzbYuiojOk1zLwvhxzkTjX
yq0sPuZHr7rISc1yabHjLiLmNtH6Ji0S0l53IUWVUpVMkuB3OzRyF7VcEelTv74h
GdnEUwFXvQ0bNoNXSylPeJ9wEA1RjzWqTRJ/fJ1L8dsvmWsTfMAOY2fPmwATZi3o
wPhyC2EOLZsp0RSPSU/SqolMYaf8PfkZrdciHB1u0i+HwoGXQCDKEFX4qUFWQ5M3
eFh+Gz4O0Y1BZBhlbkNdj+u6sr3NEitgclEea+ludrRTVEXYAx+s7sF5Uq84k0wt
IqW4kN9038uSOQO6j8sLRSlwBPzR9HjxLqfk5kRPtz6Fb4YPJyJf7OcpcqR56aPb
mLGseMGzTNYHkHOGTkzpGRlV9nJ0BakTeto8l17wIQrhZCOtU03UTaYqxSnCL+gy
df4UlUORqk6W1kMjSXPjXV+kJHI87jC+CPQI5OYY/GOIphb0HnNglT+yv89N1XIF
m+p6JEFM+R88oG1uEqICmlEYdI4jeTH44LQHQETWupRZF6fAmj/gM62+6irFrFtC
8IwluKmHKlwTAMATHv1Yp9PPcMSCfkzByZGwRowlYn+wMm2xYGbn+oXJp2tyGpD7
EZpTmb9P2Lf1+75LkKTiXfjsfXmwAuEBD258FmH1d7/PXLvbZtHNT037o1UCbi4d
ld1s+5Ym+rLKcwmKg/eTrk2r07J7P/UGFOF1wx5/kbfL8M47DTYurM5sUMpV/AeQ
0aS7gU4o7mpE54Cd/0IenkD+hOHikhFvg166gICPmQ8x6/jj68aRLg0MelKeIxbQ
P5Qr8rsWqUHKGdlltkxpHi4WLXXC8vMDVHRocvyzXHfAloDKLCSUgNijLDSQgUqx
vm7YEAPdF4x9g0zdyuYtUlEKwcXlBQuh1PzDx4+zhorTzab5Xk8KvvsC6VVcJKyJ
mebTHwDu9eWnbJ32ErievtNNLdQOoovzkI7nR/ES0meywKarNRWTy/VWSeC98jPM
p2ZG+anJBDRZMeZuXaHqa2C2m0m+hd7kGlpXxIzFHxiGm+hoOIhSkFsDXTVX/vZR
WREJms7jfv28gbQ4qKyzbjyTjE4Hvxuz6N28gn76+4C9PXBTO3+n+T4UYaoe1hMl
nnsjIZrwd52n/y2lYka/fG2MECj9R4kewFd99qAA7Jg89E+9xFREPzlFovXfAI8T
MTsLbz5QmiB8APYcXRnNqNal+xP6PtR8VytaPo5W5flWlMIQyacmcYOvTi6CJJqq
hwrukBGCJNwWaSZ3aBdb0fixQeCC0Lu/nMzXRQdEBrXM7aqYBrbinOODbCDyjZ4L
3rgZXglJjyrj7e63GDgASV80lkgBwf1njAmDcRM958m15UzA5NOdqk2SVcINezCh
HPDf+RSBlZwoxsus8PEfwiQL6XFThySiTbEYUlH6qYyLte8QXvLw985f04wOcF86
YqOx8ZI8zV7T/ndOgkZ+u/QHSQALDF9VpLDo+GCo4iDwj4rFcfi+oA0xSQ3yLRr6
gDzQ7SHM8XkTNAXgWpoo14hDlmyIZMxXo1QUZL6SOXAVcEuYfK4ChpmkH87RxpJL
FtVXZajiAbJkMNkGFp2Xcm5556uTKtfhw0/cKvakPpFh9JK5QgpUXXp9DxWcAnQb
KKwc7fah2+8nOUhkD8WcINk9j+ZwlMnDcxR2Bzqhn4HXcjhSAynDsx90P+9Lo3QJ
7qpQD2y+sbn8pNM7eg4/zXvr3+uQSviplOzjd+6Am2/ZZIhHyIdnAOHDrC6C3B79
S5h5l73BxSfEj53u7LxOC5HKgkE+ATQJzZj1ys1uiQbdM00YlNjwARgIyMN+Eonl
rF+HZdqBFo7YWjouYbrsxMzp5IGLt3JNJXED0AauirVibVi16QbFjwmvOrqa1Uwl
3VbRidAN2EMP+P1lm3AYTOnW709eJ0fKjP49P7h52JI8xolT11um7DuLttYdgKcK
yrhmQtxEpRV+9+rJ+DLFsPQ1a9qFq5MS8h2Z0sS/TgbBW5Fi4MXiQ0x9I6mdk31V
Aah8GnU5a+P4T0POkI9qLNL/Dsp1scLAkiQLfvZFGYdqsIRsi0eJ2DXCKQk8uLXu
L/UJikovF5FZuI+MASVv5Er/qss80aUPNMD3k8M22+hckL5p3IxK8g8yNcROe42O
ZEfm+ZrOUQbn5pRP3rl5inNFq7DG2P57O7aDuiK1jYJdUm7/XNS806yRILuCIzKy
q+FQXRHtXaM4TeMqub000tiAjrELqAsb54H2ORpi3ksus1msG/gz6V4DyJ4EVM9Z
vlnQ53sOHbH/tJb3fG1kM+bq6X7y56vmshIEHIUIVpur9QiFOfAXdHKzj7ZRmuC2
+mZVDBeXk3t7lxhs2JQben4JsumPV+Xocq4hZ8V8XE+z+na+oC3A3bT3g7/uJqZ9
IlMAOBlX8/MesBKe0V3zyx2pJCa9Z3eJHbb8P+licBVCtnNRL4zmMkx5UXCXVmQg
ojIPb+gSCSZdMXRQIkyEt2+eozehs1EcoXRMpLncwlDggO7Y56YERpxBiC7dz+KL
M3pvGf9z0F0BGEwW3TpctO3DGDVKNJZ4y0nSfFYS7iHMh3jZrEb/2eswegh9eQ84
jVy1JJmv9jJ9spqtzwGJJHtm+XtWadTaFtrxmMC+GgmXs90LnyRZwW2dCKX0Y7pp
KjlaRcYKQ3+Ipjy5cPt5kcFwlNg7h6tHy8ihBsErSQMgP2/SnWCJlRAUxwaVukP9
f7/N9tW/BB2FJf2siYLzQrqn6AzaoqcCCZz7iXs2ylESx+79bz5f3pdB5+lHFXqF
MlRK5EIceEg0V3vwzjwF11pp3Fzl053Zzus2O56EFbMaNWNMRjt2vmLKnjWkSDyt
yx83zlKDPmRPk7VBW32BVcJ3VA9Uv0AXOCN9gV6rX//kLeLfisNYU/GhbW0tsyZU
N0NIkDx7ghyR4GxnqIFNj4G/aSbilHKO5oo3yeyneiAP3XkfObu5BZeeXQxUqzlt
6B2nCA3XQrW7K99Tjpzdbt12JxolEkQyXkvbNTkxkZMcNjzUyQkD+EbAza41LGOw
WeQWxXHG1cD1rP09qrntms7RnFJhTGJGOEeXwTjiKDgniRONWlxAln8BnSepSH7z
SYC8O+H9ytecMFXyWf6ZI1TnFWBaPizHhMiigh2IYxYXRzdctJfTPkdGoL8VYmY/
RmWbbs7GnS/Jm7dPcQXwbrWSNEwFIvE1TI0sIB+ZXrtdkJ6VanSRwn6w4JcbtQQM
fTxd+wHnbDVV74YpoYGZY9ix/kwMOIA+1gGvk1+PEg6seO6tz/uMbVkq3ei74YWU
FYhggxwezCeUw2I16gUhqm9OmJkmcwCvyWTRpO7JByifDyPi65eAz87oLBm3QN8u
lC2xn+uwP/hFRzrbKflSTMj/shvlOfsjLh0bJVKAgmXupW4pfOAJB1Wq1ixc0s3j
TLKjIZcjW98LRO52ly+zoi6gwb8/MWdIHVg3lj6JleeJ7Xp8CPy6Ra3Cr4JxrgSr
fTHPGhBocB11EuvzwI+0BZg/DdvPEanWHI0mv+TTLwluWisqWCdWqnLGdBXktqAf
y1z6rxu7BUJB00Jh424HAkVMnYGiYUntISviXdDJ8HdEwihGlvK6w7wOcgf2QifE
SyMFFZWokpk/KMKfzMXmScZSqZ+UYfHtGkTgIsXiyHIMzhXUDVD+s+5cw6pcb1cW
9zpsiQ984fk0bWcy9t25RczngxgVrZD+NNlJOFXucErNjWyBYYG3kLeNhvw1uJKd
Q+4JcTCdfkM+OsuAKQ9EAps/byYCAs8YbqFlVkxeKQWc/iZLWrsYd/g6QsF7Ed+i
hVvUcQmhxL7eUJqK0lcXX7GC3fV8dTIV+OPVeGMKfCihbslJgOH9Hih/h4+v/DWf
k+I/9mpcFH4XbhjViyrVAedCsYzITBHHyk0dNxoNLsyYOzCxdKHnBhxyQMAQaqlw
icbPY+otBZd/hf2zms8TBcVk1BWR3+pPXRI6BRGCSn+gSrb3rHXvSJQNnCHc67vn
LzpAFltShY5JDhvfs/EuDlXv3pWy5i8YfIjoRvUw81Y+OeLxDhF6eeutMGYv2FQb
ytxjI73SG0SbwUCGV+BzR4up6lt+5vj3Sxlzbyr1DmTiqUSXHGggGKEomAe3bykU
JY6oRz8Ebvh26mO4THB2ImoebobWmH8dzKJJ8e+N3vW049GxFVsXYgQCNHnqQgAw
bEYPwHyPmygateA55EoNrsm0Pc5I0GhKQTJB5x3fxSQcE/De40BWV1jT4ltdQs2G
Jfusdk2AojyHt/H8zD4gyyDp0QqZ9/6cUvaAZYQfVwk1/JRLL/6Jy/tpTmsPgO8i
uqdrW3JGiYP+d1ggEhRqx1iEOYVJy1sF0lvDzOcIUeOG6HtZbPsZq01gMsDduJw6
WaFrDAdR+zmdqSX5j0CsrfSD+sYWEg9Cqu3gUfQat1FQlTcbIP9/6yE7+CgDz/Jb
5/WMnUuz8JJkUhcUYi4BJpwh+vNAmVJ/tavRF1WxCk/eQK0ojcrzW8LJRCHUvdB4
9zGJ/pnvbMxufpywn1G2VVt+WZaivRZ+2Iqa6lAdzXcCoQIY+DOm7/JyK3TX/wna
1/ZbN0XytUCgfrTGIjlkvva4GvRC4ld0gk2EKF6BKtzDZuFU1yHxZS1p1pVa1mIa
heFvUXgSK32LZ45/GFu9w94N9ShWLnsfqCEwNA312K1PIuMVeUlHZj8UxJNlrfuB
Alx4ubzVId9/CvKKqUt3Pfl2CbcSP0MMy3Vmzm4qygJcBhdRSnMSq5aUeid9V8zC
2G1PwPU23ZgE1zCMAHFxW20VN+DMRi/gFwGJWaWW2eXXe3FsRIQVkdwEaT4OTB1S
mmz0Xn2mN4S+HF18N2/yHg/FBGfs5L/YIDp/Rsi620OcPQrqh1pYF044t4KjFrXJ
ZFIHDBYpApr2NK6j9Pgxqwh2IMQ7mXwwJ7RCebVSmfzlFL4WpF6Tc4fdP+skbB/H
YpOAyO5tiFYPUpGM9CDvonyW/6yWNAKSJv7mMWajwKFLwiYAh6dUwYGdtSemsSn2
Xn2NZch7JwTHjVCDRh7w3AA9xH7l30fldgt8+QzYfQCxG0Wrj1Yc2w+rylH4bQbm
MOtQQOHHU28Xqq7Xl4OUL7L+SVQsZBtP9p0dKcVoEA5BesfhoMaYcxoE3kCnwWLy
4x/NUM5gxnzBq0U1AfrfMC01iCCRF+Dhv/OOueZBz/X6dJ9U8Nc+UIyHFBKMDKMW
f6qljQZL/nYmtFNdh9XC/30YlqYaYIMeWfWpla6yK1HizRQxbt2njOwQE9Re4XKu
nPL19G2vkfAYNKcNFCEmDN3VPIKNO8JxwkuPajS6o4G5DGX83btvQWZEA4tzVXqd
SfVxHgmuxySvNS6GmyQhJ2LI7bbcdtvpGbOd7d+XWGIGfX3XODlEOhJ5vPBbRgoN
kFpR2vVbFKWENSa0m2/wPfWl7Q0peWppYark0i+xuRPHOK61Znl3TyTzCJDcs/FV
lZI8Ndzw9hogkh4+MfDqflOeaZ05IaSiM3WRyLTMyj8Vku3p+xnLH+j2GtJwzpjj
Wirs4CvksgRdYeHzJKxF8wIkguoX1poqN5n2SRoh3vbHG/cZIUBNFsfWg8V4Gmcd
r3Zg4QHP6MwTJGRWGsbMeoiuuxzSKKZe2DLxxYfozjLmVi54ryS9x/3ohtgI4uMO
yB+8UpgWpUNkiqHjfORS2oTxcHQ4x5WZH2XaxaVb/+INbEYzhtXy3UorCOIWrdMS
T7FCRj6SseXBoBgosW2qeO+MpYnaW72VuFEAjN4sTGRZBeR9Ffh/EBUBh2vOsygX
f7Fv5exGDflenaexg/D8MI1YAmpaPV21pMeVsPYImxTQiP6nvQHl2mJpnuEKAhpg
G3f2BZgFFMNieuPIryAFL6DxR0M1ZDX0yOFeXZPkP0mLPtFJivgD2826r+DyXGWi
j3Jdxy/enRSpGmFmKhiz9RCaVYxk9uK7b6lT8XENLsUnj3RmahKw28WzJAHWR5SA
hvs5j4nbwP941LpI2Ih7xCzQ1Sd3UzHIxuhPQl0sgN6FzhCXjn2vgKPaNyRPLWSm
0F+ErctH+htVOdgSat3D51ybkypbCK3S7Hbs0CpS6lT/0Pn12KmECdCR89BOwwgz
QDyudyrcW3uvTd5d+3mVvnT5LhvceKC2qI6Aci7C1YIP/k9Nv+RxOz9EWJa9a6mT
GjwX34xMAAP93n0p6T7FZdE/03frmBQ9VmWuxrFXX8Qp9k0BHYpuYpSELttBk3Qg
IqeKP8Uwk/hjGDQexEE/TubHiExhSTMNgX13udexeFFsnyaIxpBikO0dgroZfGrW
lZpwWDsDxyipp9BpedRULXjVtbMNhxjJz/+8Z3qbH/V8I6Eel1QqwE0Av/JX2A85
IT7/NmI5a1UKkHgC6ZoVe9V0WJi/u0cNwF98CrClz82NKb0POnnKlVo+zcby4Dh2
9aD4PxMm7V5uB0c7ElOTrcnHaqj2a33xMdZqOs8rl9V6zU270te0y8x82Gt68Z3g
cjotGcv1Cy8YvEj37RtCmjmB5nZnYOCyhipqtfgB4zEz3MmSpljqbTAfEI7u2B3I
iNxb0PlCvqEHHhIiE5qR7CiLKa5CBVQ6qboGX4ihicna/FSBFv0ZYAydw035OmQc
iHY6KlWy1qrvejYQCzldWv3k7WS6XsmDniUzQxnholt35mmkafhlSkHFT/oz/GAi
kRZ0LgEIulbMkf0KCE1rsuFW04AGiVgCpUgjhJw8jCYTJObSMnSG8EMGlpmtDiLy
H9SuWxlzVS5AizOhxR5wPQ7we7FhkJGr85W6o18mY22N/xPd/NqSFJha4cYLa/7F
JQR8MUSVc9xu3SaW9+JkgTuSjLRQkmAXlgfjE25Hbn0TjcWtIngCRUFApAJzwXhj
qFL1oj5vbn40J7cRquI5UsBe6gdyv3DA8g11ZRTgA0xhfLtNHswyysvj3C6/BaLp
i1XTEqw2Lewp/b3suUGX7ig/p5qyncH929gZ7ZJnEHZxoCa9maGRGwnIXTiS/Irm
lli2vc5fGXyyBJX2l0+n2NmMr5wEs75XvdNm/CFHOccD/oaq4z2PwcfJA/3FPa1f
/kL2/ic5UvcmhBiM4/zptf9axgVyk588+HYl6dqOxtliHsY1MlaXJscMj9lHBV9F
D4BzVhTvSDe02LKg1QRxPOg4IVBGu2ZFnztH2YWsj6MKVno+gVpn7BhDyJk75+vx
xjZqV/rVJAryYPrgyQTHjz96fLlEg3dkQOOY8YPHZA3c+3Bxf2f4BCPj2I5AMbkE
kWoTSA2mG/zzUrLXsVMGKudyDuJeUkf95DCQL2v7hP165vT0xdP7iXxcYDKRj5k9
pB6IHGoccuMB6A0PKSdiZ/Ii9vPsVv42CzDeHk1vpRtsJaNejjOdlIwpECUe9LcB
A/E26NPx/UtpTwN0cDsl+BDyYQdFolUXRei0F2x1JEF4K7a5jlDjfvWrTpgGuiOZ
UtZRQhKEJEz9MG0Pp679ThGK31JrBSHhdiQtDUWmVNjFkTWw4TXaqZ3jHGXqkx7i
ZdffKGF7zDwDXymtuPjJ5NXi2ecJNA7xexHOYou3i+zxvq+IVdRZ9kDypoVjV1Qq
iuqBZHMA6XzJ3VVEuLnBoyCLc39NGWm5mDzeORiMEU36mEJtt4qIpkbaLk+IU31L
ByxMXL3TkPGu5ewo2GMDfao4dfQkwbghEXrx0WQecQTeIm2Ng6tdvK+8cY6YlVP7
ODTKS0jLVMSkra9XQXxIElGRoADVlbvI0p5l34o2NZfEmKzNelgeX+3w7RPwn1Ka
g7ISeSJCNeSHfOVDFkNhX0bqD0mxNUyIFtF5WEoioSpsGYWB8K1RBtvSqtT2BA47
NMNR0B3L8AKmZEDx0xrQEIjBkVmU5ydIouOiBBDb1tU9aVrNcNOOa3OsaqwFv5P5
0aoq/FjSChdO9W9Jw3jVAOT6N7DPspRFy7W4YM3qJsXZwcSXOv7gColr18balY98
Zqb1jPmctZSj4jdFGdFQbu3Vez3b2cl4weDEYzjV/XfdHqiFUH8Z1xJMPYLqLRxo
6hs8b0dBxZ9MQM2dHU7zwVxsOfMy7RjiS0vKm+xI0ob2FJ4IkNYVgEmWr8mRrfgt
0JFFB2a4qfGBaok2iSMQ+Da0R+1YAlMyXvlkXt0F7uSfDTR7ZioihJcC8qUZvQc2
9cWb36i00gdzW7/zmXiiESgZTuoWjHTVcWfN+fdU21v86cKfFD2YruN7QUwUtZzp
ragyVzWcux6NTCePDpBidgKreZCr0c6g05/XYvy7aWEHW98a1BoB1T1BbgUI4HG/
RQnzne+XKz1tIQrSzeSd/5/9+PfX1Hi/rQKJaoSxd5CHxDaBbhVy9HmMbXqnh+uP
7MiWawijjbvsVqyjDoTMllU2LS2/6W3P7+qkvDig5wsnB+xXTuDLawuzxHFQtwqH
bFAkxtmqRflEQJ+mmhni800k0k/oVnQbiezk0vP0yZ5FsgbBhcq0rpawFqmvDGdm
hBlunExeXBBO984SdSgHjH8ishtbMjimikHizW27E8ddy4Aq8QXMpIVdf4ps57bN
WJPpB56GwHD7ki4veSJvODEWheHnKQPkCi1C42G6ZeRjxtImwjplLOEGuGhE5XK2
y9uZ26j5CnhOc13xQYGWySKK5hHY+7yheHlFUfcpqQDA7KIf98PwkmjnZ/dyGRDg
I7ZUgfm0zWAjTQ7fWAZyFTyflmCeeR2d019TtTodzsgnGIuyNnXWy0zWCEdaCKEA
4F6YVApC5RLUWQwzjahTnNg+jXY2Ko0kD6TjdJii7bON9G9DXN7YppYqC2lxAQ/W
c6hz9mhuVYb3dX+wQZEP0HbRjaKYAqiMenAk8SNfyXKeUn26KCDt+CtC7fvuQwwa
hLTquvwe76kbkrOgFMojy01cVT7Oe9/HVY6GYhBiUlqnmsTGapASnMP9xY5WyWd2
XovcpSN4ea1b1hKbZf8rJFCs9HuD0YuX5K8uGCAlrXhsrrETPxYSrZzc4WsDwst3
SfmHC3gTH38wCRztzrHZC6ZsK4iA4siD++Dy7VK6Ud/rGi+FclI41P7G4qkQTSrC
G3a7mW9gF7lTHJ+naNuATZwnkNWgCxvtvpNplQ5cd19GMg2eXUeFeLgcEARpTEvO
9TQgqpSAU7h/ilcZS5LPTo1lhlUn09rdwkmoqa84pTGpzeytscu3EYUDhJYM1oU9
yUt7NQsI1lWporYqg1PJogqsp87QXA3iVKY0+tptSLVSewlaRyGj5MULIe+Z494m
cV31Am9J3kge2vicsqIkWHgC2J1X+2BwmRLij2j9Q71MBj1iEz78ZCuzI+BADBOP
VnOMi0ixM6ENw8lkuqIFs5wsBzc8VhWQf/e6EiexLuLjk8wPNSzy9p2sLWm2TfZK
rMgsZRYw04OcaY4oyq5szjxQFBehmtSKGuJsP+/O5lrP0/m9hNHuJOjY2yziC90B
UrxePUINoOVfpsNcPkPwDv3TbpnGYE4ryC/p6wgtgKCQMt25TAg21K9sIwmtqR3x
3XPJcOymUEvayh0KjdmzpVMMt8CD0V11VG0IkK6pCpJnjJzh9VB3T6ZeRi4/+VfD
/mCRz6cVetsyFAWELLr8YRvHTyxTnHfIUVc592I7d+tyUf77Pco/qMWcITnPCJ7B
1GPTC4utVkMb2FvB6/nt28AbdWrWSVhzdx4eHTlUXne/K/Y9Gh6Lsocudx8UXKw9
xCxfa0y8hvlyP17oHB5Xhdle1mK8/LvAB3crJ5TfrR6Jwnhp2Ou+Nd+EEdjlKAVH
iClWkYJx6hxLzEQTLKYJAG8mktW93G84tJPNz+EjcRdUS/26k5vyJ4ldEpSuTP8Z
qBgWUgh2QLf6hNAz5EX1fkTp9l7upQ0b/RhZKqWp/x7wIXzGJMpjTOlmBwrOkmXc
vu/PN/w/ihbIjfcgzW+xXUkBQLW632pr5MPhEv7JNtcuZdMR3u0GlL40UGC79N3H
sHIg7z/1WaUShyDh9KgiIeL0XqKyoE7z6o0CSu/A3QLtX2tSBEiw0HwThTVIM2BS
GMCAbTW/JQYpt9mg0bLZ7uPUEA2s4oY3siqofHEr2QrcprU0/iq3OSFV4r3Q89ok
R3vyhtK5AJfpda3hE7HOFM39iwZCMmB4yRdSGrQc+zihspZSZwaoD9eeJhTwS8Z8
bnoJKYmKKwyr39GpO0hmlALKuPpa8qPUNswae3RaUC3YRsjhR9A69GYtu0IDRlax
9aedoHVjZQ6K7/JQtak42lTAHZq0DQElRBP8Aqm842f12x+kLNc0yKxynWyW6nYN
fVlVexa0O2oFIt9W0rRzpcGOHy4izh0GuaY/9tsKANOkbWD8o+FuF62ZmhrCwrsC
fsA3w48XaYX7Xv6qcyUqwYVIOVYTW0K+6FKdVi3RQu15Z7DQ9ObVzmFfrWx0ZZcs
xHAIsdh7oJzWUmn2eqNSLiFiB7ZGnnGOhMNy0ditFAPVfVlhzgzilRVgU6YmFrOb
XkcA+b4v5L1hSS9qeNPSPmGYHV6cyFgxRnJLUajiMOpNfmelzzNVUDSAAn9+bdQ9
9BsfixM28XfsTfftuUTTHEiHvgXJ6p/xrqFD4xaSHLRY7/CypK6FpJuIiEq9J2tX
8pX9dg93UrkAf6utX2eA8qZ7id16Ld1dgs3ntqG2z+d+8g+oS04HesS4VuNjVv+c
ewOTsZM2kZ5RtaHsGoetgu2n7ZNV6Xct3KiRR5M1jUnpxL65IhYFlghcf8gPLPBf
RCz+90QWSJ2Br1b5Y46VkSM/My8gtexJYAv8nDESrBF56VcfUESS/RlI9a6ZC2Bz
xM1VpJK2YLMd5szmVejkZaFnIDPz1IXb+F9k/ry7JyU5NI0Ia5kzYiYzRbK8Ea6J
4D2+5hg1F8qAUghEi7D1ia4JvKXVcpYGMyUvuUkaJAkmGHn6hhtTx/vRcP593Pwi
ij+9HLNFFDLq3cxNBWJArsI8up1X+WgvJhzmcrgsFavczT3jZHnKmOMAuuE2qmxb
KH+aFnD2cYo97K1bWC96ruWbECTx13TtoIjI2uQAaJYkqq1R8rRUe0AANI+YtlLb
e7PQolphRhVlvzla8l5tquHWMjzTFykwBXNj+OeakX412uNjsb+75Fp7YGqyDBaB
OoyB5fWy3mkIqZUExz3BcKBjw/HrwNVP+2Wcp6s8NKvne9gzm5xqSrYW2un4RPu6
kRLaVoRPAqvrmD3kW7Zf1rLLx2ugalC7w1b4rTHtitl9gEbGcHraJlxLyFVMfSUv
+JzjOGfeFzPEbwSobovSJloo7jjv59vouDJFRQmRltIq6a/R2q5IPOtz9hKdyNEt
gmjXSqKmIxKeNeYibuG7idnZ7lFczEkVOriSv0xIbBNrPcogc7/c9g1LOKv9FZRi
kRlDETqRYVGdoPnDj7lrhCGzQ1QQd8URjpzTG2PQUIYT5dJhzRJjmfio9v7fBQuM
KxXJch52UFaXY1kYd8MkLWSov8+fNmfFeIArbQoaXhuzueFo1fcS+1GKehmq1Rwo
Y1EzOAW3r1yAoCV0MEGjZl13GzTwFblxSrgbmnCSiJP7i2x6p1cGPEd20x1Adz3q
xetr5v1cwAmm3jMWlwSLtcmQIWpAIKv+i56JjS5VtVSW+rI4EYgr0HuZc0Lgs/sM
/nhLCwH0ZtJNUiybb2UKIQhtigPhl2pPrkHh3NWxGHKLx3D8PmcJOR4DYDRaiFIC
cedi09/OYj90p8uLpu7F5xFZ5GM7bwsE9WA9vg017RSEdAxnCfYXajU5s6XFg14j
H1uHeSFlFnqIL6sKhn40y0jcYNE5lIRMkJhVN9lu2+r27NeSZKCTAD4g86OOHTj7
oUNbaoyFxsaElIStLkBZo4dzQw8aEsGJz6AamDNZWYbj8Ev9Wfbn8KR5ZuM+2QBf
At5afQ9FK+JqdZWUXW2NbUwJBFBO/lp7xX61vHaAs5Rzgn1oOsaUJqV3/ZdA1uv/
FOZVPoEnbsyvw3w48jAkU/RCI5iRo579ipYC6EgLBDkvWROd6N8GhKqnLixrhegB
ylY42fjkhEWuGkUvWmpNwdHBEtI1ZehCvW/dqFTsXjm5w8HPUsZntNGnrSVEKEN7
U82z5uIW/fH8CoFAzzpL5xW9PF0P0UDc3pOzIjAWXx1/AevmZ/LRa9z1exxfjllZ
1bQiRBACCWUYv38f7G8xWL85EJh1XuqwFWNJJpfh7gwCG1hQb6xkzCAZ+ycNnZCJ
4NJnpiF7G4emRL2qxgCYxYIfBX/a0P4Z4vWAtSzJIUiNgX+nZtlT07q9MR3boPcz
1vrbzTBYKS26n2ByBOkMh9x9pUiwU0LjoAVEoGeMi/iwq4Ok28bMVDWwA4xgUq3d
KBf+K3TQlqMuriET7+vBKxG0pFltIUq9n3Zk70ne53oechVFBEbhaTJPP5adNsdt
PallPRAujqRjSvnLCd5ECoFtw2Bb6XzMN7YSjScFyBy6LyAVe33AL8RgzZjgoX6H
TV42+eRyfbRsc5RXDbOsUbaf4wHmYS+O/0s1f3zp8zyCV9ObSdz9nVb6wdG0y0qH
Sh/h3Lrjnl1zDGZzCucR56FIhpCf1tLa7uKcQeZ485gNA8WTE7pXpVWhhgdNDn8u
pfZqWAnnjhBqVsHTsQc2oAw6UHwrr+Qkn2R74Z9PA/BloW38W7OQ3RqkYu19e6cw
KiQcCigymZT/7OGP/8oQ5c1Ef5/sbVDthUeE4jTzFCsDLDSlKLVnVBsohW5YWa2z
eNvNVxH19JyG9Iy1BhxWSWdz8NTKacWf9FAirpBaWotP5wHZtW9I+k4to/b8WAy2
K4UAUXlSr6KFdSczB4tVZlZqZ9U6bXt1VxnmWGzw2Hr4WsvbBfgeUYg/WGWTbtQ7
9stL92YfyB4raEDvUTqxi+GrDJaidT5iDISysLher2akx9wl+mnBIlABnML2tI87
1LzQK42NPIWHgDgPPlxQ/oVCTwDbSzifEnaicAtBwSxPcEpB7UWHlObTnqi1ItwO
D4PmFb9T1YZtHCWAAWWfRYnDrTUl1ObrUbSe1yVxPGMlbcdBKh46G46A38ZjeY9A
p66Aodn6DQnYrE5ILVnFp3BYRY59pfnMsuVK7QqF4bTDurPv48mM9ctcLlgp+8jk
EIq6q6pFIMXJxvPwuqqfH+EN+wZ8F6x2yFBrwUhVKILsCuRkkz2Ioq3zYkZeF0IJ
CzScxgAWNzcSU8pYH5xh3e8cME/mrfJwT2o+DsZpeGhJNP6/KZI5A/KA4qanTt8D
KG+3hEPqu4ALVoh4uFBN/QoQROqUbRpDtzX5o3MuiPEFpVJXgwhhbdiuPeTxPNhh
U0tk5qNnZJe0O1PAreJDjPdYEfVGx3DsQjglGWTEpdzaGd41sLkvRl26sHGTylzy
dL7T0dOlk6v+ZjJ+AgREEw0DFE/WP21ofqtHo++kq5PBwnOTD9EVsDNyUOWHtN4P
w3gbM3oxjQXGR79qX5noN6LD6n3vX3m407uZBRhNW4ywYmQIE3U/Xx42VrjoB2ti
VVUFeQ4ERH7AB9HwCpDKuen1R6Eonl2j4khcDejKUvkP8oD9fbfT/sG3gaAfHq7i
nYXoXEvtSLY9aJT+zENaQ6RrGmJcxc0yOcsueqfURNITKWhH5crbn9xRq3B4UnAX
pqmrXx2Cv9AIzfwGMZ5fTy/Jm35y48ucSothUkgpUV0QK/UDPzpT1hzR57omTNCe
KmQPIT9qgRzGI7KG7aRrSE7y8lEBd4TZqERXLdMNJr9ut9voynTeRJ8NymnZ4LbK
aMxexn6r3h3bN0/FC5Z5/3RrLU1uCDccSdiHWmHXGWX+Qc9e6KVBYRa5BzASVCD0
axDrRDgYqk6hiei1SDn1VfWGi74zix3ZFaoCI3qYYX7aea+FxHuL2/P+GhIz6vpp
v5cFXfcx0Gk6/2aNgUZayCWHxLiRtp5GjhRAML11mlpeKkOSDXGYOj1R6L7QIWVp
fCSqnn4Xq9QMnULKAPHmKE8l/pO1ig54Pgzzkq6UW9v/qdrPW7uDJrkYIpdI0d4d
osL/tay1ma3J+Ewxp45UEimKM/qY78rp5ek33NK3FrXtQQvAjJReffcuWv69dFPK
XMI6NUMeSl/W7KGExf5y6pWZa2nkzU+TbxAKb7C3pitUH4GuQasFxXeCcq9N9KIb
PxKUM/zPECjSd+FJrIMKTcCXU/9Ix2kzXYLjRotmbJ9osyutRZe0tfciM24JV3s/
aEXgg87A5cW5ZzaEb6rdXicViOE5rCjEq+ASEQG2KqbRVLY93oDO0Xv2fex77DHH
O++hRE1SBavHb39pDo6EnP2WjgfkQfQ+Ev3TcBFf71WcjlKPRRjVJEDz/Ani/RIB
0UnuPXLzzNFXfCfQcGR8eD1M8EdqDkGZ1jC4ZAJ+vnGEVlRuH4PXe9ixFwMyxxrJ
snn53fRdAS3YoIkIwG++Cp6C4nRTpJDCYEmJE4AaXd28bEz8qiR6IO68UTJcHe31
4I9/lT0ZNj1XdIQlWtIt01mFQStE/58jUUEzs1cDDpGaFmLYj96aXfGHiyxpTNKR
mzKnzDiFlXSV8zGyRWMRw1N+JrXibo6MHdUF3sY+tU5Ufg0GZ1psaJb2FoiiyGUn
SyHTZV2ztULa1F0N7Hw3Xv1MCsckvi2GSMYmc5bSERKOHJC+Gt/MjEp4Nzn8ccHw
TbaAFFCsULKzOGJayIVVWrmF02LRNoRvfxF8OCDWjcnDkyjHRKxuyP9BM8cjYq0C
580hqz69T6sx8peiq00aEn9WC6QH894gQEE3lzx8BplyGQiAZ21rf0eVZFtAA9rF
vHxg026w2zCwg56BtWgQFYKJQ30Il2z0dd8mXAFBXNsoVR2pIJge3RrK+/tKr9TJ
LGV8clPkHRH8l8ExCW58qAU8TbKzkwPYJpwdxf/2A4y6AhLvDdYMYrgPuWOynrri
2ZR5ff+9CAuaBW+dMgLixT1I3+f0upusCzboG94I+w7moT85KfNGMGjHtd9rzyYd
91fAKQYW3wCMuEmQA0dI6ThyMQJUpS0mFdi2GT2gnbJ0MKQl1frD2Nih5P102mbl
iqUVPX8Fr21I3ExqS4iQvtsiEJ5SrYirq4c8AkTLLTuQEMbVJ9SOfjmxYntRfzE0
+aOSlCRu8iB4W6bjM/GpswIYcfcRD+JrY0GNbNXxESWNtaHsYFxWk4sBstyjwrY3
R2/5FC/YkUZccnM1gQSolojG2cBpkSr+O7m1l+zaLnz95FCKqJIjFO3ct5+zIOLZ
LBy2ubzF4oCH43hAr3Za32ssl6Uyo8hQFdSMVfhzYRKG6BnyjAAELZqpyKeDa1fZ
jmjtxjcNenvjgT2efBkSxAriTHbYRhMK+2pujTYLlfBG0bN8Df7YTkiA4DefUXmR
mzZJC7zuM1wZiTTzZKSppNRSF7Hj0adq1SNfA+xiStThr0DJobhDXDH5CIcTVntP
Yfc730ydAxH+QjoW/ZossDlogTgZJFuiLZwfNKGWgqQdtWZrVB63VFzMgUNEB+vZ
YgPdGx2Ph1t5j35vF+wqX3telLMF+hJenY6J2dSXkI6a7qpCZ0ncxFE7VVc7ps9F
JHK81NK0Oll68bR4ieGXdCk+z8tfu3rZOFvknrPA0xIYCOrk/c2LxSg2lzX54omw
5coq37J68EiEWgBLxijLSoJ33W8fNyWn1WNlBZjeumxMGGus1mEL1oSEyVUWODWb
pdddFMrw1NmyrT2c+aETOMKv6u4ACwM+k/rTAXsJ6M1ilZD3CYBzykkUx5dz9dvc
5GC7kHj7XwatWukdWhSMn85miJAqKcC0Uvn8hV2mg0zzs2PxxuRlD7cO7SrAtQTT
IKxCnWKSV9PlyvX4+tztJRvEMjUfeSEeQTYZPSPQn3IxTBLLBExqjIGoMQnkWTC/
0CQWC0cedWDhNYtol/fXWSuEJp1Z8kVzfL7jfzAUole/pUO8M3pcxSCgneHXFrx4
ENVxttJi7QoFA56FqE+jjM1yifoWGeCYLZiwuNNlVH3V0ylQ65Gx5J7loBW6PU/B
9g4YgycD3+py0jq6eWBBKBsK2I7K8BVHPyGSLv7mtvM2bM9AZY2fhiAUsr6QEp2s
mdoWb+5QhLwsDcSMSNFjZ/Q8gqxSlywT4GiFHr3kr/RGMGsGMA5vojwHbE+TkvfP
Gt3Zz9net+0XPpG4JujeBwuL/X9adrPk/guEsT6pDjKceKip6MOqFcJAb6JhMeep
1OwDlno8XgMOltHDa07zeSBFNm1MD4WBVJ1DvtKqDMu0hFZcSsjV3rOtiTzmPXA9
0DIZDNuC9Z9gEn3S7jWC4QGhTOX5H44vhNV8kAJoPX9C7WwHDKHivfZXRVpUytUz
wV9vGmy4H/MRefPZ3ciR3ziAG134pyYlYD1ZmLL4PJ3oDqe4dQEccvSYj7lhK0k+
vQVkDqnIQTnynJR+LYqcY6cp9mmw88mwQqjqgsFKe2nY4ZIVevG8+gHJVS1zIQuG
5Hxmu3/CWjT2myiqZzIDE6T/tzrtoobkzVSpkR+aCOXa8cBjDW6BfvCAPdLgGhzk
hcwiK4fv/j8IdhGniqwg9hBxlwH42eDRX1ZmK6sfRUxDd8jRohHzUC5MTJqoxA4B
ncaIKrW8RzUbnZZ+Kyq+RbsGkGwGnDrqWK5RqxUf+cPltv9y92FVNuLNpb2/l9ij
2DK7DZlKHJEekPN7tDiiXQVQk14pQymPKOPFhHC06N35KhTMoSpfjn4e4O+IjnqU
OFcaSAmt/vgl1czzmVAcNvV9ta2OCyiGAicYW61EH7dVrV5jgknOWzyvvSDsqoJt
jjCsXoOfgGKapRSApfYkeXuZiuXy2dDmbOZQQ3etlofZznq+s1CUN2F9OOQDc9s4
J0Wr/brashpJbvWcdYW0q5yD0OqvwwhdSNvWSq6imyd3Goqq0cQlehirlZYpYVTZ
IBzojyIysiufYpYD62U7/mhd96RrZ4K+pfE4CDUY3qcp0S0O0RmBmAaN5SQpfykW
GqD9vS7fjvVvXl6sGsuZLH7z00GywysNR0SGc3eu5i8PsZW0MKCqJzG5RcoSpVAT
0QJCiWNZujU5ideOLnhW8ODJTCYnxhl9hrvE1tfboLcVLhAhGg0K2im56bnEPTRx
ioJONCtNHdQ44/S5T72JVyOs+RkRbshvqoMBIGNNrpWMdCodVfgPrpikegm1Vt6P
IjxVckDncGH7JpAwm3jB7Bl7Wbqb1pGXTVsAp4aNNz5FcKCTrGglso7wJ3p2YgQU
mjIFfzAKWK+NLfcuMc+O3vdtTYGzXrl5LmWCmxT7ctDOGppTB8277O8JwDFkgtms
vhEDF8YB2DpUbHwWwua3+j24bdn5IulWNOq6hBpRZ/tJ0c7IdMWuTBoazMpTepO3
M6pZCT1inRE3uok5o8M16La0MSdmW0VxTOjDtUfOrzamzbC3e79BEghR4KSVzpJD
91bwjFJVj/9oeg3o/y6g/3VEbS8uafb3S4U8NzrTqvBwv/v7zElvfaxYW4TmkP1b
F0xP6u3q72N3yLru/RaKiPcSDeqNb0H7L9BXXXECwN4Z1ujUZrdAjnD/STbzks+w
+DT//A1d6VArI3ffamMRmtj6TPoNQ/iwC9k4R3qZGcyAOmdvxHvxUx+XR3yZFop5
AJ+o4a1q2XhkbMKmvVZx0pisAC15iDvYq+BswTt5sudgQe/qRUdTxWgiDOriuPZz
gkqMCBmwxuPnPpj27zlpEIdoLJMnDTXpI6b7Xv6ULR8zEkni+CEtffEM7JGUB1v+
cQZrY+A+PQQHgARvZ9/JnHjbjYKoMrFUrm9aqD17YDP7KyaDofQ/JNVfBT1uTj9n
K3z7xN/Eo/Bk08kwe1cMjkMvjQXcnOxO5+UB8tFPNtO1LX9jVA+/ZM07cEl8BV5X
UMsQtDeTybCyf+knYSAS5YMVaCpMD/oPKv3ItPqWW3h9JWGAQW3cqCsvI/aUDzPh
SnhcbvkBo9WeCZaEkZbJOKEIaDO7sH1ws5XgA3uAU+AsRs8hUKNMrkW922w4mfnG
5zlHJXDG7PqWvpqrIrQP7wXC+rQrPYk2be89pU8uoB2hoNw/AW3893DAoixVC7yl
afDJX56y6eVZM8rkuH88TEYalOxO1P6Ij1xZWXwcQ4rlVGWlflW2zfmzd/8/p939
XBTL5rmkvN5eYAjCJ+9+dEUqJLkEQQocYmL9U9AH7uq5otya075OAuhIgsDIgLHs
RJfCZbJ8rlfMWrxQic7qFxXIV8aPzjEqENaARx6CpjkEfaWAbrQzybY64bFgNaw8
I9M0FtzatbpifY/A68rjqbUyivGvccLn/BasynO6Pc3E95xWFCDfUdbhnj4ZH7h/
dYtw9BlJOJmLYaxHIPB4H5NNgefrXSMkgYSTtUwRAIGMPAVWQdPvA/JwqfoUqYY/
5yg37Ju9AjpjX/1eyPUPhX425Ij2VpZkTBGC54kZ8O9sgIHDZGtzsjv7hg8CgqlF
oWTrINYa8eFyiNVlGoQcpvJY7Yd9ed19hEClKBy/9IcBjaZZVRDLm+Gt2hJtiNtJ
+p/1y1UFXcWSgsfOYSipoT+XE5IbJBfc17ToGlGKoVkUTJPkmhB9JBvLH1uii4bz
ZhsI8IsHFJWmya+6RUFwc9FM2oov2koSSaNUQjzzcnkoGbZRPfVk4XvbBpGpmVgN
xjneGcVHZPe8OqydndgTsz9eFuFLMd35zdh9iaVrpXXSg6IsNoeKRQ0rTSNr2Ds0
IYrGbivo2oaLZksnrkEcUEBKa8HekhGkiqk9ruurM1i2l9urro+M7rwahfa9TXJY
GUsJUl/n2X0h5K72YJwo1a1zId1e4UVf8c9GoSYQYym4qpRIkqoFgWRyb2hvHLUA
8eP8Vqxw7Urzk0L1FbOVWC4UT1fMya9zUWlETKHO5owp8FcglRsePWGzbSnSIWYe
cLH/pA45pcy6kqUbjC4ODJH3IQaGbCVUP3co+XoJbnUtHlVWxlJ8YQrZ8RE5L/tj
iQUAl93kbdUB7RKSDBkeicwVmQHaIKIXaZMFJIj/0ML+gIJ6VjnrpNjyRPoW/oKo
9Ro1Z+mqthG/+YtMQSihd8kNQfwLD9Us+FeUGVYy1wkMXpGiNmWb2Z/GCvMA1Hj2
D5e8k8ZYXHRqOx9DB/E93tSSedhhGp/L8Ies9PtPInKiUvPuQSt672kAauFw4uk0
ChvmT6I0cPSRYqn2sgbzn6Ehu6ibTlh3D/xvAJBsTqQ1vY4PR37COZJKdZU9JL6+
5C32mlhU9Igxjy29heSud3bMxz0jNCxH+WbPhKP5DY+yHawjaaB8Ztj2l7SKlpGi
r2AcNKco6HdWDF6dMZ49GKecNqQ4o55rTJnJMRSVpqQRnXRWR/VfknEao3PyjvgD
K5drb8PuHbQxGhkVKXAA4juIH9/SMTiFIXxr2U0tPO+OvSt1BP7DyV61xecIbRkz
DBjZwftzqPLtkYahpzn2+1e6yLHKab/8crDZ2MhHHu3MBl4m79k4/OUP9t2h1CIc
OYcwmeEMdslz79ovjxCfzptW9pRfbDemSuhcG3xosYEQXoB+o8ZAHqyz6plUrzXA
k1wWXG4iJJeLyrW0QLxOAUp664D+4px86xw+/XI7g1hJ5RSgct+YehywC0zJHfgc
k/sjOZRuI4d9hPq9Q5+9FhzpzfjCPnhYzHgrHBG0Pkd4xDOVmSKcWzhBgEPE/0wO
tqIocH0szUEOiOCXdiegRb2ZLjJxlbFPxXvm1smbQ/CYdCxnymZhQt2SutMiBJFV
XLcYMhpM1DUhhMVB3reNk8zVx2zIFRszFXiTRphIrl+WsQ8BkRgIsWqtzPaqmID5
GMwmBcs62De6peAEjV9ZXRJbjkM4WKk++zyJ588d/KT1Y2B0LhD/wfm7ibpffoGz
HbDkbOcIIQ7E9A+ucERFdVtaT5W0cERpPVa1ifHFUnT5eO5H+YbeDcgSHjIZLmiQ
yi02FvKmAhMsmUfBDl+mbOnBiUtF7e7lZqLq1ADg2/foNB23lAsdOw6RMuyXYy8D
lppTB0nXfLCJ/crye/rZBP8kw9evGuXAh09/qMuIOeHEAcEZXGmRb9c/OZ89B7mr
E0rPhsB0PEkrnI3S1XNxCM4Jpsf1NlyR6gnxzPq9czCCNPJn5SsHTNHMKJ551QRk
5I5euDgLa1VsvLILfcRWFkmpTsPGb3600wWrnGI+keLCska849W7peZQoS9H5NOi
j4tzOuueW/3LqsQUCIemqGfMI4G6HQtu9RH4q3gd7FCVQHuquYjNUzxufiCV1U0m
Ci4hm7Kg9n/REw4K/PCpsjo68RSukkAeLRbrYCcUzUdY0tFhtwg2Yb7kQ/FGlXJc
SWUTTh02eA0EVPUJxhDPZzvMK4KBFihCwqe2Nr2f0oaZ0W/mHnymNBEwsV0zJYxZ
jG/y8RKuhBdO43gvNvqSkhELF+i9gDmubKElPknOozcXd5/ylw9hZdjl9MPAoSVV
0NgM2ONF33NJtnCNAgoHMcpCWzuL0D9/GASScBNVkRZSLWO/gm3CUKpMcw8Xn6wx
TtH8FMGMZ8yc9yf5VlRjK2uezJOehfPNmN3W1T9u8aEznSoiNO7DBdwy/iJLx/lo
LKD4eYa5OTug6Y7yF4TTtKp6GMZVmLUqQ2nrAdG64wKhiHtoV0GcawozCxjCYmsQ
/RWBX8cEvBiu/SaS7cmJcQnNBs7EgLkjGOGM3P/9ImBaDrTGkvVKbRes4hUUvBbp
XJ2oiOy7B+098cDPgLcc0DKzKp2RtMBT8oAN+uB7NylD3I5NVdMbea6YvTrPAJuO
1cLqKxnuS6nrYLWv2sHVYhxEkrx3w2fhIBx3RYyTYZuQ+fIigcbrpt76s+Lz1HJl
nwxyhjT6Nh9Wc+llejCL6edmhskPhVozliP1JgnGGLGDHVvpZ65cogGlIyxE17Vn
F5zO/YLIZljqEIHlbKxKe8nt0sRvTvPbxsXCNCkUw0zFZv28OEt8l8YFtD0yepHc
DOdN/wPr/B4L3kYfST3koK4eGQoluoJ/Sizi4l/KCcNUaMdBi0P/psACIz4YDixz
SqUwHqtfHgWvUNnSPYpczqudnbDL5UQZcMqleCsGfGSUwoQtV6v/Oyc0+OainoYN
qd6stnruZsZlDqLIRdjrc0JSYfAtPitaLozyyVh08Agaea7kiA44cfSkMmqZOlBJ
wSFIRDa/0dIodN21gqNS+hBIDUCLl7xY4yOBXHLhJnAkoCGILtwJfTaGKvDiXhiZ
BgMiMURtl8whK4hXc4XgJLq7ibnqy9o3UF16Z7JDRaZEwyugXFxAaYZYFxtnh5gp
f7intM9EIU1C3lGPQjFeDZpL0IA8W8R4N3sifhqqntX4yye1DkaJkePCS8HFowBB
KurZUVDcKet8U1zB6jd/tL98M5VVyamWepGOpW+wAxD5O/kn7oFJxalOIg6s9ZHx
qzLeC6qeyR+h2Y9GOziv9WVboOFHyn3kVIPNnrC/illAWCOu3AUTD4/ZqDOMkc4Y
si6SHQs52kB9RFCadFbo9etjlXb8YI0YtZnB1HsKLZkh6HGR+m+Mzs4fA6Fkzcsg
X6Tfr9fGfx1sMsNv9upsCa9XDKm7iDOMQiaGCgP6Yx87XkOYTKPwF3jXOioXWmTf
Mv5JFpwXasmvfe54lEhZRs01aZHlnEAhRO+Mba8SlHK1+7MIFgWWKz6LhhsF3aLE
mkwhvmKMKqWOolkrPMzMIQUgz/zbUx1C+0hnryjmUKu9LMhc8dY4aiwlY45qD3Fw
W1frug1GwicK3/ERcbi3iCG0eoE2arZiZ3BkJMnOnjqMmZflrZIgaMNMy4/iLWhv
Ju6AALTrNQUlMA/DX4FCy3yDMjhw+sSeXQ9nzPXFd6chLL0IO8FLf3TDvCmI+4uR
i0xzB8sUjMdQO4nGXxJIpEHqqCHb4HPHtdWJcWz1p3YAXGbJsxtmIiKRIWA9GpIL
vtbVuw7bQX7nRltNXBadO4qdm7toxp7xp+cR7IpNvAS1461BRwKc45zXqUE8Mm5s
YU8gv8EgDjQiJKiguk5Ofh83ecxtMbkgraFWMrWgJ2TjD2YqBtDbz/oiZG5F1NrN
Av22jAbU9DdQv+viqeO+f7zOnHYh1yOQHjtNh+bSRe0nRPuuW346Xstb1akCz5MF
SJ7D3AbTVprgXbwRicCIYWAVRKt5/2xtnNGJImCFMqTYe8UAQx2NUC1Co67ls5Tc
wV9brEuNiEvdF9ABCqXo7lV3JLJPe46saoYCd/q7U2QAV44cfl5PIa7101iSYAEh
5zdq69RrQ5aw+3VPN6Q0kAGZ6oKnLmYFmiv/XLqEQQIns4B1YV3aAK5AKOW1wCeo
WxpE4beED8SKgQ0ulZSkEj760mDv/WpheqPhOKc4c8oUJxhP2YZrxHgukTOTkIQX
VB7bvxAideKFAYys/sGJFXqh3YT6Y1ItIEsWVY8L36bx8JaPBb3ZoU2S87suqE4E
SGSh+E7cTtbhc2xjnqXjcgU4IAOGdu+j75SftUnotck8VohTI3k7gLwNJrKuM4Xh
o7TzsXdsCwe1NJhcw+xWnN96GGHAePsvdf5I2V3NVqatMtpRdZdCLpZPVwTHnBCj
kDAk3VodX50dGn23k4Sr909xsewKStycYH3cXRgBrR+WyhEZTxsTttaru1RAq1S+
vWxQiqA6z2B2LRT9DpPUb37oO4PLxdGOWwOReTYW35B5H/QUwohEy0SwMD0C2EOO
zmEymRTSgsm0MKgYVLCUe3NLXomgvN9xhl5ZW54rrsY/s0mf8aHtXh6rPspQOhU7
/KR4RAR+i4Ul9GjeHyKLeb4bDsDWSvFAbhJlua8ZeUJj9Cvpvi8sgdFVTmFMZAA2
ttiCMQL+D1xnkiGRjY505U1z5APyYCNHEfLwHnlqE2/lddGnxdEu1xbe1fG+eJK4
eWtjxQQQe289eHEEti3LEZWfWtw4W57ysAunEBTLi8yHg8chxxh//KbJA3GLkrbH
99B0GksEZGIr8NH66demIOlK2aOuiutw6gUHlhy+VJFMU/mlTJ7Emih4pfkgIMoC
2n+DvYI9Cq3c6mU1l/pbkQlp1UlgwDFOD+U14rR7NxPXaYa87BSyQlmdYhQ7LIAA
16IB66Rpdutb0YMAPJgY72T6GxJ32i6ks9Wdqp2TS3mfIzWpqc009Aq52hPA3gop
KeT44rTY41F2A0qvfggPS9FLUpFM1aZJu0mvAwEdFWKg/lkKhq6Knw2nNmMrSC4n
XxRjl5+jhv244y+gZeNBjcJPD0kudNmEDpGMpjCCXB+5XWLr0k0iWhe2znBR2Q5b
EZt3X540NBFYZMlOiIrYdg5J71tnInCZX046tqkeD1VXZ3uEiSV/Fhv8YF0gEfSf
A4DFxl9wwLfc7V9xL0WodLaU5VfFBuIUA03+cZA9aZKO1s5ZKBnYvorD3PadJG8V
rY+XJw2OjXpJXBdK6f6Wb55c0Q7hyuorxF555t1W6KuEqqF3DUAO4JPLtkWLlDh6
G+Ll9js8+lJPuvwKi7EPQGWwx7J32Cm9D1FdoEqQ89DIPbvehhWDm/PcNZcySWgE
svdbtOI5kaQ2Bwr/U6NCK7qS13F6C5p0xl7Q2N4Mtkc7UeCdgL1CJO9LezLrDnW8
jCjFracwjuAe3E/5Op7d18UfMETmLvoCDfyd1hRi3PJGYbIHsL3t5NHwXziBgANg
jaxqYG8tLFe+XYL1UKNYtn1wpsYFx8jIGDtFgOPrDz6ys2mgDFtzBvMUXtgDQvb5
dBtxCBFtJJp/3UjzyBO44EJogtzSF3bIQJs/4V0FH+b+ww+US6ZrwIZrq7p7/L3i
iRxa4YtK7hiDrZjNWnsonTg4WA4RhWmdGqeewGO/Nd00A289NRWDVLbPlPjjH5gT
AUWKAFEUGFDT7W8FEkat8FQ5AaKxD0qoHxwS4M2vWR4icuQ8GhfBSVMJgzgHJFkQ
WtsqRiUTxq++k+FmnrJuN/p4qSZkdbVtCi9zz4kHnGjtW3gXcg6NczAAKwwU916s
JvHqH+4x0p1zwnsQyFuUst0PiRxjiMKWRqcadjhyBeKymAvAHmyGAn0Pxkgik2+p
Z+Ct7PSz3tHAf8pEG8Ub9002ikB/yMvvNLDH4gaCuhGEJWxpoUfE3xklJuAwAWI5
EXWw0+Ns+SKQxdv9YBGhmXZhS6aPF3YO5nq5TaYTmnCY0fR0XFWqOdRejn2vEXo9
BgEPQqNQroV9lACwcCLuXG8xLJdOIUjDc2gvQJq7r7ibNLU9EYkkzCemI5CFoHbD
5B5cM0oCN1vjfqjhJ4wd91JWHZfUau9qnt/OP2oIVomkekvmRLRttCYWsw+FoxD6
235FY++9ui1naePtO+u0jnXRHLTTftwaeofPjJWSKv/U4elY6EMA5oBH2lDzTevQ
f4cOar8TciQ5u7fYKiv1GFrkohqFuZvRG6SeE4Vo5Bmreh+DBS4SR3aSFF4arEqk
/e+XqPB/vteiUA7FFOc/nLnLNpOXCZHrk9oSQnIgZGCfn1bH6LLx8ZOTLnu5aYSs
lOrHazFJ+iSMmIpfFHZmuzaQxozaIweQzfxYGepoA9ka/ifzRStP8QoGeWQebTm3
n+acVEmivjTq1Dg6e9SxsGZ1sfJ1xaTuwyb39cp1r/Dk0vNIIsAOnwIShfEa3kOX
b2N/emXjZ100JuqMPs2Tciqn0zn4FxgCq6RLgfF/BnU2e1OWQ912Dd16+Dltetdn
IoN907p4OHHVE1tFye9NNMrPZ9FnNiLnE/R62uFFl/860NDB69npzRjslUbbbeqS
H1KU2nNy5Qw0NS4EfNR2/0pHKvdqUSmCd7FsB5h8M72G0PV/nv6mzeZSZYQbkto8
uFslSfP2EYzLaBYuj9YZRrWZQLzyj/IkGCM8uNrv0bUENKCzk8j9yZygpKCYeYJR
tJ7xlcRu4YgU4vF/JziMDpTQAxo1KmE4awIeQSvoY3Uyjka+To+fB2+QruUCXkpI
5G3l83mAyPI4G5WkL/clElQGHlPZN/cVZjLrJXc0T5iYXk3547vh+mSmdbFLg+7J
sEUnkx04viBycJb+EFhJvK+10VXKHA9uHtu7WgJKDgg9JT/C9Ro9rkmYIvWz1qq5
TmR23FG32WpwQjze+siBMyuOyuSeEecqAeOHsV52oEVaDb0K0p0JPBC83k+y5+23
Kspnzzn/7rx6kfPRLq4HEQe/RYS3+rqUwl0qyvaJ9shNRqNs3F3p2F4PGbDukyu6
YZqfBzldghM75y4R6zY43fUvpKGzHZXsmAMQUOjCiUb6KuuNCi/XgeQuHQI6oI3t
Ey9bZXi+wTldjCp5C8/4dmVtr4jpD4BdQ2IUVzj5yhCXN1Ozf9slJWSjkcM2nRnQ
zUUH86vbyMYdTvj1XJkQQkOywHghmx+hprdU7Dyx5HwNfGSJyzrqpcLBUQg2Zizb
5REcT4cZaX+r5M6r5apKlCIucRn7QALoRI8P7yRRJI0tOJ48izQVnVWU6UoN4Nub
eWsbnQNTu1QNkawynoIE2vohjacGR3RIUB7Wd40G790gPlC/3doCgcroAs+GQMRz
e5KBX8HIaPaq3Ne9x118pdU0jqYIp3DBmGPTrk2TziQ5kGkKe3eBnnBSF6qWaxz+
CZhaIeVTZERuvtrVVGGSm4CgFJVYPzEcm1VSshMo9xxzTR5+NycRYoac1zyga5NK
8Hu3Ye+2FPaUtB6FgCAgvZsvKH26VEM55rll4PX3knI9O5eFy3TH3t9JBQBOmsiT
9lo2cz7biu27vOOnscRGPMdgxk8f45V6rhXTtz7mkjS6KWYS39YASaGoIHvCLCdc
Upl1329Rp4AHNA+iCr/mmAiPcHBT5MDwla2Wxg5kYXbx4lZUkzintlKTSzDMeDKI
0r1qwJSo0izcoSihbmbBEMTZCHnzgY0ldL3jWiatqk1HLiQbm4haFSLzTVt/iH0o
3tqKSwkoJNssWZQM4tfE0kUZ559/DIxXF1fNhBrAsYQBWEBwTTt2UCr7+k/13sU8
axx3OpiNaE8H21sg4F3sNsfCmJwFuewM57SmeRd1pbBZSvex2tjcC+1q7WuWELIL
txTEglqBbhYetDsjhcYM4mnzCZMa2XJVCzTztnOQSh7p9FQy5/V4HPf1/sPtKAzH
m2DfZh033QGukA7Wzi8ngGrlUVyHmXXQ9xrsJRl2tZ6G6B2mvE5Jl99UN3Nsb4cl
dFkwwBru87VAgZqukQ/bQVdYNfPkvaRvLMb2ORFfXtxNUJHgklcEzWjo/nu3YNw/
BRDk1RMCpv3XBtbX1V61XkVvjsfEt3D5PxfDTG1W9IoTV+ZwwAeVcdq9YAvIIZI/
dVXB5+rlHyel4jw9HgbOS7Tv86McwunmkQ+8GUPigGgY7B2Y3k2tZIRojhGJuXiv
iAaL73G58vn83D36knf4qoePhSwtN3RwnhAP2VpkWGNKHIys3tlWeKyodk3wKdw0
RsRzl6dFpM+7Zu14l0+v/2nWfWXnLPtifjhJnm53jAF2P+Lq1dJCDDF0zB17lvsF
pBXgYDMo8hML1zzle92x63qbrqr4BHe5HPtgTG2PChPF2qF6LBVGiZmrJigy37Is
MoAnk1iERyLfar1Cn+eWgNo/vUDx24vA+HkfeuxJgRBHP4sj7fCmf153RwFSGiva
96l6Zn6X7AVNeJSQqNr8PgRpi+IFiVDANOvRJStgVJ/sfy4SOW+XHYEJqnbKYwc+
G+WVEkJtZWeOnkeYccmXXrNtwDymricAIWIpGVB7Ogz4W0BUmDNgM+43kpIXhDHS
KKARalovpn975vUaQrzC7wdFk7lPv86AQurbAMr3w7zOafErXflWqE8Rk6WKp3SO
1IK1qsxYx+Z5iXztCP5NSdzOgr84sR47floIzTdQ5RUo6solDhWsxa7nb9URi59g
08QDaSybwmLQ0cLtmFuvYDQKyuNKb9IKI/CqQY5Hi0u3Hfqp09X2s7aCnJ1jbyku
qjfBgCKPw8L1Svb0P9N0QHqAVGSYiloRtVKADkuPjRX3SdHtpNb6yr6KX6m7BJfr
ywStNxMODyAws8nshjafnzAPOGp00AbQ0+rTFoJfmX5PR65fVRRdiK9rFtl0CLS/
eexAuK2vLgsAH8S5plza9c/2c0T1cBx9FeZgxqFtS41EdPnOFWEYPg0cISrmratF
lvcPHO9vjCKv0/JtIrcUHglJpLOWkDyUSlY85jE7mYXmaOKrDCXo+AJMNY5RB2yu
reLof5eJr1YfTts/GcrqzsV9arcxnuZRlaAtWu7NHLpSioAzdSRHh9lJPtuJMfF7
muPpf+m98K24qSbkpS5y5D3RrWNejOFen+k1+ocawU39PQtD3WFj6N6wnlKhIx5I
rqShIo0CDY+gy4OhcYGYZWpEaUqRLbA6HMkuFyN1FStY8dbQcja31UynM5nrNQiC
4arzd1XAvavZzovj4x1a/GYwU5/rYQ3l0/298uF2dJAS1/09TIJXnc64d6J8o3UF
wb/LwEFoQ0XL12FFQ0K71c2RbUXxGSPEm9+1ByS+og6Oo/xB70GBHHVGTHIWyezN
DYGLQTcV46ugEAe9AY4EDrNP/PQd0WSUG3I9IIg6Bf94EDPbwgxEWhmGtK9ZWyi9
DEgmI8opWmDXApq7JnzRFGPhhEN0b7tR49riSHqKt2COOSY0GL0KJJ6Pyk7iCtuO
2huRf3WTfeSzgJlYYmBV/581azL3n9XR5c5iehINQGOQ3F+AWu4RR+I3EzK1vgB3
9w7ji0PnelXWtbKM7pZ9P8pR0O8aeZZ3qrbCekHi3/3t56ZzQUl0lsktV+bUpJp1
BshxIF9qDZ7xbYhOUaaHHO3FftcXZiK+fzmYJTQNlSqOA/c+4fjCEwyIKKQwgN1f
w+vOuqUXn3CIkZLczzEp+X4SVmJmXmP/4aYxrVYStnG38HMaIeLHJvfVyzYxqxV9
G+ribDRN95/WkFl4KHcnW3HhAQ8X0ZYIxLKOf3lQZabN0rrS6IWB/RXAzb/MXer8
/BJYAHggGTPIlH6LkZu2NMM3zGmoEzhH8hEDyc/pHW4GGoX1+BUsuic9RlVca9HP
LOfA2IlGHUS7vKI0fvgZj5MWIEJlgEl8gqpQix0kgLp+WqKJHWaOF6ItFtiizhlJ
5hkDgzVpGfThME0P13HxGHzIyd/RYUnoTmIRQhW9hW1eADtB6kVNUEfJEN3o47hK
mwyiYubyKxROdXLhSMJQoLr5RorC+EQA8TNbMqc7KUEJ33ZanyRfpusLj3HRoSQB
Z/K9SdosXvgH3byMBwDH1/iRbmB2xe6mPb/fY9KUrczWaoY/m3htcD2dXNh3s5wX
xLNsXCcY1TlrpIVrccGLWvMq5H2bhjOHtSvoPTfgLRVolvxbvdYn+uKof1FCm/PC
EWcYxddQ2YkD+ohbV7C5Baz/FADXmtbuaJfSnERS7juVslEnnOWAIEAQ0HX/FT0g
cs9otfM1/wPb4cJvdz0MsA0p3SNsX9xtYhXeW3z5ePs9Emn0vQVDeJeAMqX8TOQe
4GMl0NtD8YC9tHlXqCPlQ6ip5oWQeYjK1y+0BOoTDap76gdqkCtzIG3zc+z+enVo
mRTmy0m6i05Ez2oYebYpVzz70ChKsMJQkoGBR+FTImSomZ5RbHwkFFbmx6qe+XGW
QQCmfYyCdU3gqoNG9D8Uro/U6LQilIrlzXJGXu3dZi5VBwMiEYtyzUIq6Cl5fVf+
7vFN8S3LejXdMu8q9d/AVVLBBoyH/Pf6gumjYYh+fIg/HjReUglOfqxUnc33SZ6E
+as5kumvXrzQcsxLqtwtIL07SSEXFwSvWOR0iUY+7moBBBXQRygMF4DB+FmlQz0O
j/BveMKgCAU3tdQhf6B6BR1vLqNuZgCOtrLV7Oru2AVd79VUN+bVqJYAF/ugzX6Y
uQmdW9ylxpk5CLpYnNfwETojh3/5tPso+hwF9rrYh7kx/Ga9CmL9t8A4ZDRnDt5g
ochmAsFBH0I1MvkB6sD+sYFz9chSIowRDQap/AL5+++JBYvfvUlO01Jq7nYs/MnP
kAvGGWKGaTo1xMt4KXLObnAbO+kakjahHzbiuxVFuvkhGFYqvmDJ86+F4SAEkcTR
z250urKmG0m7yjDMNzI/K3m3pvb1ZScOaQv4OHIBA2D4CPUv5kubsvq1AfIDZqLg
8jStWYpKojcVOGkU9TNFmPhqWax7lgVrMBfc1tRTxLQEFwH7HN7zka7vjtet360i
bv39Vik4EjNxtiPDvtEr6o21aF5rburDyOYwhydSaia4ZNJ/OTQ6Fl7U811SgsMf
K9umg44x2NvzUVr1Kb7Js89gTBR0maG5DmmI3wfIt34axENBsjkwZx5u4GtCMqnN
nqH5yjVDUm+GMPzJoHWpJOj4ZRzqYZVaUuhl/B8vvelWz9SX3keCVLuV8rqz0wcC
KChpCzkx34dSn2bInf3FkRq7iaaOmRGgNvcXa2VAoFg3A+D+4W/4s7aD0FFsL9kL
bLuyI24ksLRiIs9XGibtCBKD3NRUhgn0g1fcGN/jpb0Mw2DHG1awnxb4YP+7mKSg
jshS1VDfns/ZF4Mp1bmIqaUnP23MOUij0hznmUKYGlzfTs92R+NvDyf60PLmOyOO
IL2IT1MaIOw0HivXMFtaWyJ8U5I31ijam0XKS0zkTDCkUoyf7rH7zSFB3nrUZORf
IOP/J+tI9zsezegs1do8A6zTolNiaWuKyY+Dx7kVJQOjo4PskTBTX6eqtzzQVAfY
rowgLt9/N5xS8k0CvmmjV7ADB19i1Z1SoVtCJJodDotCdcid5/RQEoj3orrrk8h6
KcP2o/R0IJrAm1uEOZNo42Sj9PkUJaORjm1iNTPbujU3C4JX6+4FdWmWap4RSMWo
NdD0TJiA2+juK3vLfVSEr1Y7bONn0eT8Fw8v5l4l4y4DOiq+AKJiAqavLTWgMndu
1HH0XRMq0esEAd3JyubbXvJwNb8Q12Fjg+FP7qe5Fu0tSKEOjA5g7ejLHRJvakNu
J8D2GUq+o5PK+XYrLGGxu3nimr2ASHKBsi7q19OeBzWrtTkSTAFaqtvxblk8VWuE
o1I9bsVbRK2z7KHHNrALXsA5BkN4rgVZ2cuDjgo25tu+h1Kpd2MwOS7BAAUH/4Y+
TsaYhbcCQzsi5M/2wrAxj+MAs+T3+wWNGhp0x94Lf4lAhvUYc85nY+u5MVEDV7nT
wfIQG++4uAAaIes//G5uWR6k7Y59rufI/FODBAItBS7u4n6b5uQNkn4hbLQsN+5+
uN1MZUJV26epECSbEL/XaJil021+d0lAKUZ31bq2r9wBDGviMNoobuUTG0Fl8mDG
6xITXzPmE8tNi5iAry78EYoHpz11FHtxWlh2N37IQCxAlGNUi2B4StUQSXl/T0i9
uTmdp1CjUp9OhrFYJ1gVN4R4sAzgvq+uPAfQQapVzyQ3jTeaPUKjk6zidBuRmBX3
yadOQyf+7x/FVyViS1BimdQAtKwIVSKw3IsjAmh67tzZXeTwnjko7yhs70b6iDsp
Vtv8rt1ilnptJyQ19/J3Z17oFuC2mhz9j2krlZFfeXJAgoeEeNwa9bzvxd1+htxy
HMJn+rOFBVoApNnx49MEtTJ/kKWpUEsRS+7n9lDz848NXzDHAdk5BLKVhEU5MEud
lZm6sWhsTpbPROPphjKjdAVfJquZA1fdy8jbmVqI5lg5zoNkrRcjcoP9TgBPyqpU
Pu0eKeX2bLQO4Vdl7uUPRoovk73TKbXHHaRfDpwnrpzQzj/CRjAdDe34629BU/pV
QvmSxmnLlx6ErUtemATx4hAikIkUCV6n97+cQugoedKGDXGV/mQTHXwEUFMUadCt
bq36vQf059D6uRkLaFd1xdRMgtZ6WCSnlSQj4rIq1tMm7BotqcHMtmwZKQZyGPBE
/+cOvtxqkEzkYMv10EjPiOGIVPt/Q3GQRYignvM7RIWvyQUx2fEpUINSs141HZlj
XzvevzDMe4U6kc+T+p5NIulA4hjQugzkWHuTTQL/zi/1l95ud4f1pB/KHdgW7Gkr
g1TP30241gcuD1+Tbglctiaojamo3oZfEJ18G/Us9/WG2l9PeSxvqKQJHSA51+bf
GebunNAUhvVZTEq0cR8MDpgqCFZx9kye+fi39FxmI1zJyrewowcrJ/Lqec+Nxw17
YjYMs0XEQen/GSQf7e/j4tKoNokpKteYTUcx3z8u/MAf3OQifw9q2hjwXDU/H2KZ
DdLDzRbIued5Ek/8Dler77akegrUGqWiJpGsDhhWO8maqaicEkJVny90T5OSi+KU
cnsC7Wk7Y5LuedU+2Jhc1vtyj35to5/BNhd310bYS5HeCXvpeeb6VUflF+RNL7v6
KsKACL5v+ZklU7O4WVEYZWG3vInYVWd3Y1pe4OHsTmSgNRCEmNYd9O4lJ5ePXaYi
A5HHIrDzSpv3pL2QcZPv/5o18Q5wl0i0FugABGmM09ghOxSzgmPqD+/wbd2v5BIq
2dHdF76SVRAAl7STA0uYR8oG7bFYTIUeU8fsqnKci0ZWCdjntCyDzbWU6DokEkZW
1I/17Q89Mg+FVCgTKSO6MtHOMN1PSQW5CKVAZGlDMbL+FUgQGi0qAs33xcFk6GEc
xRUGBdaPoX8GO0ZbsesnYC45bjtysd/SWc1wKoS8AU5sBRf825+bDhOQXKZpteG8
dGB6FqSwmCGcmM8zsKAwAO61VT6I7ET2sINOcRbCYcWct+38CwlRTYCeQSiOGZJu
3Mm+xvyi04AOyVwmIWhzRGrPIjrXyoctSZDvBXWYva6fROb9tx5QL1HDX7XnJErE
8yzJlC3r3EJ08k8TRHjUGgXPG3aDH8LR+wXUmi5wtpGNuHfdoHKgujnemQI0WpN4
4eI4nCjcezPLLhhceN8/lWgqUBMLQI+fyTfsoWtvYrtUZu2DelW5D09pCD2CQupq
o+Kk5lyDrvF53ngxxqEXXgCZ9gug66mJU4XX2Ul5lDtUH3hGN4bFOWn+wpee/GoY
a/AULDykzRB0KZv9kNoug8zWD9FxBoiAcMZM+abCCuG2ldCoEzvuJZlUtGOfhkN5
f6LXxv+PaXk7FA0msUphXlJ/nEp7dzfu9mwprKClhUF91bd9ge8cghr5+HUOXxeS
SZLjOibL1km5KUIybAaf6JTCPzDsV8bXpb1Qh1O2OpogxOXvWojXY9VyXkMewfSi
0x5bMrKY0nMPqB4IlttHS0RtHSNGw1YGuLJwnd0aKisi44DBCjSGRzznqZfWhuzh
658reQT0aA9Lg1uCbAQViQ3yibiWrcrl5Ue8xN/AQhafg5ZXAGgvDqdRuB7N0yR3
P47GsZKqMhlLGgApoInmMZz1UuwASAI8+OQRSmmYuWQVuak2bpQ8fzvFOF7gsQ1R
2Bri5aLg45dYbG61dPqQMhkJvD5pWmlfn3Vp5Ogm8xs1buc+7DvJaMTHQL2vGH7h
GdBb6vSqCMFvmc6Lasd9vT87LsNGuLS+03gQwVSy52p43QuOe/uX+SLD3ddniAWL
kofmPDCxumQORsWm6m9w0gHiPvTzhU1OoDiwQjFD5ps9cpzq/6Ocg0QNH5UqKZn0
rzNXuIZ5ITYDf0B5kcUyR8V185yQtBg6w0qMxYnBqXeT5gUdQ5ne+nmCvSBt7Vur
9bVPsWXMBhgZ8NdT5xdyuimkadu7k9UXwmqoAGY5BqMUlKZ9nMKeDdqoYeITBnVD
/Dr8lx3hRZQe9fTV8xJ1GVeczb0FPWRjUPwmsS3r88LTWAxjmHWrbxk5frpZMpFX
z98Tf+1lOePbfB7vxLvTiQNqQm8eWvBfmMnyw9DqMmr5bfSZZoB3F3XW0BAE0wwC
IwmjFClUEKNR3eEUGj3EqA69mR4IPX96zO6u4ehbpn5xcq95vUEUQ844tVXD+D/b
M2oy5Kpt9CRKopL/OQlfJ1zH+oj3b2dBqppwv8PxPq+fqmg+tcosk+SnCS1DcB3U
yRfw5SXZDcARASYIv2bntmyW/mOm43JLai6hbjwAVyl6rFd35TcBbyY+JvQ0uxn8
AOGulIs+z2PIN0nnu6ny8PoU6LMLd9IhUps7+vuSij//UzXsQjKxKf6ASR+ks0iU
/c7jzPwBHwrk2gQOaCEnD3C2aL30uKmRNQwFY5IUMZ8/dSG0MiRZN0kwOM/t8a5J
N7p/7V7KrvvkTVmcDYIDjfrTYpAGhv+PMY5wRRRgQetBxES9e360sRUBIQXUETPp
XolTV1dx8xMRH4McyzVLMzVRFjUnXLzKBYE1GRXwubRiwSld50os2mDvEZpzYdyP
MALCxFHu0BXboZnDL3LNEc0u3RMHW0mgQue4veqnm8dn1aBu5sXfErtV8+8Fin+a
5TTsYaFQ5zPac78nWoM4Md3H24KCfsf5Ohfp8GIQj5VQ+FsCVAec024ano/WhMKT
9GvLo4UgKsn9sLeeM5JwkE5X/I8dWy0o6efHuWPEWnN2qxQtYxObE1/N2ZpfIoNM
n+QopNMET5xUmEn0gyTh9gnbnRiQ0syAui/uARfi/WxUgfleX8mO8zAC0wUkbE+l
e1uNfZi4KMtvl1S8NLpDaV+h6RmE4oQThqbPzNwil6Gn3+A0Dk9S+RH/NxHpAaSZ
AFXfbkYwSqdAfsy4wFNh+5ogQiu+OdN8gumqYFEwxnCZF8tj+fMTs4mQLPL9VUZ4
OfbMQnLBnw2TBxg2v1sd9/lvf3mVfwiqPWy2wQrTOjaI8Cpcv8/R5Z+ru+2jCZpS
CATrzBO0TKnaCvDzsTmpPkUvrCiaacDYvoJYjg84K5BP+TEFGwMP4O8tUpKPtFjf
ugu5jqOzlAoexIG95zVCRJiCLLH4gEv1Mt711JUC0HCDlfBQh7nBf0WBMEH1jag+
yFifJdnJaaPXL/ybv/0kh8HhJY4CPC/OMTcJhCYJbuREXkbBOD8F5VdSDX5NeAEW
Yuf4mBVMJNGGt8naz02BPfT8xUr8q1PJtIKy8cnNeffP4f4Dx4iJFSr+DUhvQmWl
BnHraG5+z36W5ZpIpO/20xbFsbO9cBPxpDqcaIhJDoVnZlJz2VUAcFPY9iDz3Nk3
MFJI9UIV09SXxZcN434eNrZB1A4lkFxrU3hkMmFADO+wJJsqZAdQsy/L5qlMWlI/
443YtZIGHF2kbRo+VlCl1VZzrkhnl3bO8tDH394hvSQDbAUHQT/AM/RjlNw7brJJ
9IpfCEVJQ8whyCMM3MIHETQbqZKuvmo2iowNvjf6H3cHXG0CnZIR3alBAD+NTAVM
+dwATuWzquRJ5iZTWpCxiK1RYPmv9nKXdRWZjHVIjxUSX057j4odkN7tN1VLKgHO
4q/hKPcwp4QtzaE0mB2j3SRtSsD5ts3J3vdWNnBSKMwsCKSyrgj9tV8YLKbLAmss
jhmdsmKGm+bQOsKO6UAbTs8LH/yUS86pRg3v6nKzx+/XMiJO+GqrxFrqA3Uy8Ifo
srh6oxezcgcfRaDyNRMAETvz38GRyjw+mImI4pvWcgAjrtRQENQsI0se5o0Nsrf7
irw9K4X5J21xFWjXDV6CNkLQb6F8jHiZK6oZgr085CBGg7i0XhCSuaIoUWLkEOFl
8zAWJb7joRQ3Xs8YP4KTj9XbbAmHFzFN+eT/9Lixn/u4fltqhPGJHrVE4ZLjDhjB
MfkTN+05CGgsQoN1GaLEl4k1GvyODEb9I31CjDfNtSnQ5adZ5+3nA6TbAm1T7okn
8bd6XmS7Sj3cYLsL06moHOsyIrbC+rFJNrIW2ea3GrN/d69k01t9g2Cx519hTech
7pzpDrNNNW+BabWwC0ov/xHYEL+25jMQjCUBts5dydqWDjTUuw7l622tpalYGqkK
uKw93CE6cKJJ/7RosEx/rmhKZJK79+ohNHxL0YFPL9gS2eaEYmAdwYU/vGhyzUaS
XcghSEOqpYRVtM0wREPkL89YDjIGwWwNBKCQ/FHzrR5fW4bOQG+ZeHyeYVnU7SUb
TtmQEe7i9oL05RIRTEiMqy22+uF5HGU0uTwWZpQywBnW84fYie6XGt71QW2hybsc
jRSBVj2w62V0FQfuPqsecY3zOzGpixq1Z4cFSbJMg4ZLdO3T1YLEtpXKUyQaL98l
A6fAtAi76r64puBok6/BEXRtk3IIVor0ieYuw5XCocu4Po9tSRjo4ahYuUiuqJ0S
/Q77CxKsPR+xhT8V81HknJ73SeBDlsX6R5DONB6h/+2Y9ywMvA3JsL5ejhYzZzzn
b51+o/oNtiGMn6W87GqoeK5yOcHHLE2yvGtQDySI+g9DUq072f0zhEDqwAzrJnuc
Kbyzo1M2dpuM5TUGgwvIpUGGYfYO8voCb8P/LFgPXXwBDwABlKDfGo8lRyOWIhXz
aJWyee8Jy3u4K5LE4HYRmsnYGNEhZ1xkClMrgDlbJVXedpTJQr+k6pBjZ1duMxW/
7Sb6TrY4EuB6MV7S6Fpl05mJf2ggoNVJC2P9OAfrSdTKuO25ePMbjz2oZSSZlMsf
QH3tcw7V346HXJgD5UyOM7xh8dUq2AA6I7Y17p+cYOeplF1ZaZZcjwF5YgIBuiAS
5R9qObpoO6mG2IebdKKy5rAve7RiBGZRVf6y5CK7yTnyWt3V6L1+6ofIvXVyhF1B
AL0+07qbbeCrmqKBwqdLVcPWNwwK1WbVe63p6NNLYAxlTqRZgOiEQUxEPZj7Rczg
nUOwQ4hwFROI0B1ROvtWwrRtY73S845eYjq/brbCF6Z4vX5/l/pmmu+K7ic+5vix
jheD5v66B4BDA6RRz2Z+Mc//0SrgGEggxgOpAw+vrbUBTAaoCfm+xO+To5Nltyii
NTkQ5yxaKAx4wMn/witgb0au3RCf0oCt7y4zOMcyOFgHgOD2hGDUPj1Tk2RlLima
tta1r6EVnP+MSr/GGeWOWB4MSK09BsqHeIw54Ad9j9EagB1VFjHc7FrlA7DG+FG8
/KXBOGFgNXnIlrJtqFd8lXhpSQg6Lh2mCc4zJPMnYMKslp4cUlw/3dJjmRPKejDR
DPo+KzwBzc5Bms4A6Bg7inc8zmLWjCc/knOWT34BUcVTL7IggtBeHR7m4NiV9Fbc
yaz5Guai4Vz+N/QU70P7ijH+OYA5N6It3nuWQFbgd2c11YMfoKkUyLgSEss7wqKy
na3ykXYBGEiu+qb823oNCz8wE27bhwilheCLhfM5QHxA3boJ6gvSqY257nOIA79q
PN/IDU5Aq+wm8bciComzEnkGYe/q3NbVlpLwTXTpZ6xVpwKDRHih1HzViIFqqYtw
KQw5ioH4mzZGqITrFGcfqEWHWNB0DKSK04XaYa8rFw9imLL5DnndRvcIL1UJZuRv
m+3PGCoMTT6IntWldW+QZPo0U93o5Kdjo5PYF7hXwJeQk3HJ8xs43KFbfnzQgjAw
+O+nty9lyabwOaH4cpvWy72zNGMYQdmYIIaXj8+YZ0UnyuJ4kQhfXes5/lVvtiBs
iqDfcCqwQqLzwIgQ2u/YivA3sDZA1rGPcVx9vcVz4r6HNP3B/MseOJk9Vet6+xGG
Vv4wUOG3LyJ+SjdNdWV3tNPxNWLl++l/ySdmtJxgzQQbFKCzjI0upD77aQn1OT6M
I/jG5IEgxzB/zlM7HZpGQ2Jf++jUmbgaMU6Sruq1S6b3JahwbGELwb655Fwgts/P
VwspmEeiTCt/lNhoq4+qApAB0c/bkjRhYoNo6hZkLDH4LcPS/V4qoXSZ/hQWEdz+
0EVyofFm/h7MWyHn7MhU/cYnG29pBBUZLIS4tD1usMCl2Kbg5FtWEv2MO4UT9uiI
Z814eGygzxAz/aWhXzEwrmOJ2+bTaAlMXYYazeGkQttaQ5n/frV5z/qe2vrZsRSx
+sgzau90CO1cJn28LiTTrhdK7bvnP9MeVI7UfI07CTY7M9s9UCheoYUcaKVEddaa
ag7ELsBrbRzdqJXTpdrBVfnqphat7G2NN+xVkW0ahc7mEDSsE8IWD9RLVIqyBYe1
Oh/JW5J3DpWwksagNBcGCHjZRlgmQp/A4W+wccZWNheBXSFP0j2mqw8TjhaBAes7
fHijJtNvoYoc6k/RRLLf3RXe4ZF6mOJQDWTI2v4TFoYgTzuh0EY6NXwl3A5nVTts
oANhEnFgYd6nKZky33GVZJZs6Zr7yD5tHMMNdqm1mYobhd91/V4QralKepkZW8Xd
JJ5wZDAV1EimDObPmM7LiC4GY2X4DhNpMMUK9AB6bNSnHS9DINMCUT8uHyxfrDw4
+5vTZ5fFBnHosaLsbNNO6uNhMjs/a4BOsf9GHgmqFvWxhVq2r0TjPh3paRB3FVTn
sc61J4Abj+zRSZefTTiXVEri6Fb6ykc0h03noigo9R6828pgUMh1YWW2wyj2unil
Pn7Is1m8TJu6cWRPcDoAQHcj6sgMvSYUmB/sKjhU3eeZM+37zez8YLBvrFSLzfzM
unjcUTxQQjH2EN24J5krSmQOHRl1YJj8lDJHrME1M5xLIThpqoZTACuoXviw9XaA
8K93jibpTuX/5rV2uczwMeufkGZvWOdJ5Rwa2aRB8b3mWHNmLEQY/sF7PkEL0h/V
DZAEMeI/SuUxnzUwCPDvZ6pHl6ovKKEup3aQblPWA/V+oBTztv+8ith092EJhoTh
gunKBBFcyz2yBKrolCTFUtjBxWLVaGVO/Y2JeslMLRWy1VpzII49wOkLfOoQ/cjo
zdZlsr5MLdnqIqWFHffMh1eRPsiq8XbC9QaKnKNz5CZsSTtYtggMMgQ1+7b7YJZ8
9Ry5QUEkdMPZoyk3n2W4NPiTR3knYuJOwfy4kOC1BxDXaGnwFNrttTPnuo3tito8
eQZj89XB6vcG+q6NSYlCSDqhQHCg27OMz/Jdv7R+gtLFmsS3S8dh4FH7Ts2FK6+n
36L30J7aAHa0t/w+5IdKykW1XmiMl/mcm47w6v7gVAKTYM0MS8Gm+abdcqDG7SSe
HaoMo1qf1LWsz9tbe7AqZs/aRxcuZHCPF9iJLUncDASiZ47XzAomNzoXe7Z1H5KQ
4gBv2BpanWq2imMHUK5XU+XYYNiuAqh8J8+kZArASwL/hZV54iafJRv6gSDWMiaW
XNT7A+FLgL421PYtADZQE+8r+gA/GEenBx7962UinoGS2QoF9RUvAwonu2SGS75M
6gUtqE/GIrgQzCCyW3DCaDH0AM5hCD1Xy3Rue3BFQPlSMeYoJJRYWQ0EuAuxvuV9
dgZRoKiOFroQp7FdfZWIbWW2fBVfuR4v+2p561c54X/efWyWRCiD2QZN0oFP/GsT
bSxVDun/RRuGcV3/JbLeZ8ygqxsfdqj0x+PEAcbIjjg2LMd3USbzZ57IC/OGPNr0
Qv7oLaO+st3vpVrWC2oEUw3xft/TzfQ1/Pasobq75rKJdvI9nnl4KfepyfxZ3VYn
LVjLimTYzMiyKONYQFSsYpIoKfZluMbsMyX8E/LovpYHmC7/QY3nRYa0AzdjQmaz
h7LQ+vcxWA4Hc0kym1mVVTb6w0pHnlKvuYCTzOUsvcg/LudmbVOBrBoEFb57RMAJ
33d3pkmTAF330K6iaFLzhR6XIePEMwNQar5rAE6AU/L+Wb3+oEscszj70yXrMtnI
WJSdM00OcGo+I10w7cQtuo4vS1UE30AdVMeY/JFDvZI77E9t+/U3KA/oPISBUKOC
VOiKnqfYMDt7mgTork07LkAfMp0o25gPW9EzwGzqZ/OECPrLUYj2slu/oHHoLPTP
cz7X+syw4ZvbNUgmKMqK50n7bzN7SO8TL6X++4NqG2i2nLc4hGy2K+D37G0vmxbT
iEogQrFUCynq3WbThWYGO26o+Xc8aNqwXKrE04EkZRyNYAD7XMBiLI98nPbEUbhT
ozx4lRFFTCASaz3cvSTSgljm+PZMsL9V7fGQPLOn+ZEXEYxiHCSarYmABLt1cO5E
kv78lZxKOBwPsXBAAyyGXdSXwzMuxZMV/SPfM07xVzkkkUuxttiZ7wsUIs+tdmG6
6a8HZwLX5zWxoqNaS2fEdPh6JU3tV/EhJw7h8jZhZ1B9f6N09qWfgEn5ThsE8VoF
v9ZkH9ZXoJxtzkqBWaqnsk930olaXm6v3WXBpKNJ1hC3+cXqFhiX+9X9r7p4GBQz
RCNrhzMH0UsiJgg0xWlwLJxi6Sai41z/eSphay5fae+g2jyapzA07SUV2HIjaVEW
I9jVKjbcC2mNuLgAKktFs96GwERekxolnGMvsxUoIzy4mI0zmDzBeV8ReRlESaNQ
+UlHgwqTo6GF7T8M3JHDTuvdI2Nb2E5cKWaB0zdgrUu2tHLP2dHR898XgMq4AiUt
S5pOoDw8XvYKoKNFt6yH39GBnc2eWntLNcJ7uJ5sQWG88WZWXaxkdLkllsY6MOLq
Mbyf37DZc+eBmepBeIiQmKLFY5qujfHEYKOZ8QGDjVUYrMG4qcsrvQzi70f7mhHW
bhiq+n27LXovUqW9pcRrwb6cCdGCPodA4a72fyrFuoI0GD3fX29jMpEd5xjMQrRH
gRYOlL73MySyxqwx4AAB5vDGm9YQkKc+AOrgrKAM/OZ/k6yTgvtoJ04nKPj7cVD6
ZgL/k+M5chY3i9gAwicC8chSWBal90D01aY/q4jwBvnbqB4qwEdoZ41cgf70m/71
+wThmUBroFTUtzuzSFFtxYkpbU+UiqUmKqtDPVhpHY7nL9/P2U++r6a3ebKPZq9c
+b4//0aoiBivgoYhpWol3qBw5U6+amF8AcEmJzJzX1AVlJd2MbHZQ3UXk0TLY1iW
eN2ybYRUu3kBNju967ImXfX0ykRwRcIO6Rj8DCoAzqxPl00lD/hVkhT9Cu1mJeRV
KC6BbFoqZmr+3qmEAysCtNj4+PIh9z2xeLCqsJUkSnVYf665r14sTioJOiFLyK0f
jtGUpGPXMCZu38VzuMNVwn55yIC36plpPrU/+lyw06/7qMH5PHsbxSIY5xdpIU90
DP/rQrfAl+HV5XiwZEmJAifgaca139aJs/8LMQPV3YSPBiZyu+4igYulJ3ZO+oHE
LIvzSfzaEs1nTqMfRb1PfiBpwRX7no/9G28FGs8XjCHUynAJtzTLTwuvgHcTGBTr
wrXjmnYXcqs038h0TuQXvi4rhyTHKMQg0fkQCQjMNSnGDxLrPyyp0wcdwqXqgLDI
AABntnYAouH1W6mADMOzlZVq8j6drgR8ccQgJyXr8fXIAIaSq4oJRMuWYFOYqARg
sxeNI9LiNxHxmnKQcEUEpv0PYdSrZFbIzUuy8Sb6iqHGYaqJqFti3PLybUFmHZ3U
5IqvgFTd8outXV5xMoKUs+UCDQyHTJGjFNzZdE6wHa/xE4j7dJ4ybl4lFZSE7wyZ
9nC9ikDWpwlZBsDWnqqn81QamwwXBntuH+jRSUJ+I5+980yS0CQYZpGX8fLZeFPG
eqT5kQJrAvbgrRxLuVdVAZqpxiO+/TdIwuKvwQ0gJYRXs6DxbvtO+CtE78Rxdi6H
6aatKe+G95V9XU2Y+E1/fDc7XfsNCKjJN426tW1GUpoJW+6+wqYanH+0IJxPc1xW
IC6G+3C+mn70Yxril+bWEIp9jKvrZFXWIZHOKNq/lXs/qhwGbrUZUWGRhRPnXIYN
9qCsQC3eqRJC3wfgzeZQk6l+GatB8DymjY0MXf8Le+zL41cahMuT2yaBPc7qrLET
FSJ0vjcjUwA1qrRt6EY9KplbTf1o4AJ5ZLrdJze/GrxqVv2C2hHfctW30ZK4OuG5
GrEgQnU2zAeYsbjRQBa6DD//ntUDTSJcAnoxI6P4UCBFNfa2qb6S19vnGOd5WTcn
/PfjffuL8nxmO9Jn14pEYZ1XpH0LRGU0FIto15DM5evV+2265o68f9odIk4QuP0v
Wd4v+8dYn3aWWn00JY3cijuMP76MAAQYnjTH1hClYn/qYxqd4jLm9C3cB4YsDYZx
AWdouJqY8oMA1L/iaeGsWw1ejqhgE0qnIJoj0REjM37ilMKQEUFfncqd4b7N0Gdh
KVFID8f/WnFzEe9TqiyrKZQAI7CRzC7W8eVTOiHxF8nDFQU2ybYQBDkU728kXqr0
W/02K7filR107PUIpU+sonRuJnxnwMAGKoiGUW22gb/Cnkvv5TAQded2s+n/IgmK
RS2XnpLz73jDigSvPoUyi7bQsb2y16rv+Ws9cCakJq8tTvKgTQ9xby7zTBWij2Ny
lhoaxEUfUiRjP3GKZeH3YRwc6yq7i5Ec07zVI10Ux+q2mEknIJ+CasgfCr5UMyRd
B37m5O3bVEzTzjRLRLyH/TKm+LB4fDTbvEWOkQvArd3cyG5N20p41Y1Cpk/zxBM+
0FatjmoX7tapnon6oG3LFOjKylux4brqtA8c4LyZcSQ/xatOA1H5TrJFK9nbSJ3S
TtGQFK67CWJYKJ4enr3K9HVZMXEYWjSGBcW4sZ7zo93gVvh2qUMuPuwgtyUa0t36
iDq6xWv016nIVFpo8SMlP0/0uUGzWJEgGbkwyoSQAJ1+qtTahA1z/NF6mHXgpdj8
fT14kRq2prtMf4cn5sIAiiXVPr3NywjivFpmnIOmGYqi7vgUbOGVC4saun+6a35r
ZcSDRXHK6BZsxy1WkJxYtkOrVvQ9CgQLSmsvR8Du9Kc51Xht3+/C19wEtO6w+jG4
3Is8pj+PSuL0LvCDkVyC8MQRZjHKlA3uYlwQsT6yiPtCQb4YYunQhriPFpG0HsDJ
Ha6EUz9rf7us3nm9fc4FvK1Fww3aX66qjnMugaA/OzqiPuTfXn7021Bye9HUeBeu
dnEH2OFzHQQcSBLHAPDtmrh5DEPMWvaR9dMMLVXdkKJHNU26U5iiynp3DwNrQrHr
YVuTCSz6/FdYYPIfIxlgbywZKZlIS81/Oa4q0IwN96Yu3cDIZuo7r+N6H64ZI76s
93RY3Qf8Lecn1zhSU11npr8vRGh+xwWahPMpqRjExJAoKzha/+WVbRTfACLtMIGx
YEUODbLGGWR3m3yNq0ybXZZVMnPeqG8TErVcZ5t8XIA+xAPeHCo/9eGh4PqAZ7Ys
6oXyNjYUgPtlXEpBboS5aVmUx3Ye9MdvCmsroNRr3p/WGCaCrzMWprDR38IaHopW
Yi7xoP6Gn8kaNxjWxZLIT7+xr0R7lKL5tc7vCDYHp1WxaV56fDlrCpUzUdb58rch
NEhvzhhClIGc+RYsn52wmlLMuaVALlgBfpst4DnhptZDjPMxLM9ENbns1COVYMsz
cnta7JyCLyuhKFC1BxKW9M56jyxhyvK/rIdZlBLyYrEQYGqdLPvD/YtWIPGLWt7B
t9tApp7Jce9ppJnNCD9BheAx09kPcWN2Z2f+ZS4iXjdqDfsg3syXddXtUSwSTkYZ
zgdkSDtAZBfJLJZpSPdevy96UI9MnbdSRjbDBPaABRfQvYohL36k99M5c4cEhfUE
ZLHv/f0/7DUF7wka4JkrXQDicK1geD+YPs+fWcMz3fXfxDXWM85/0zGaGgqiss7h
tJMnT0+Egyty0n0KWWnWph7dUbUd1Iam6F/GB2ehxU8cdvBRmn2U9xqyFhqraQRj
LvLrYwZM4MqTQR0MuveuQJ8bSOWuj/uFoGSUUhk7YUE5qKZhAkfDKM6bmhRgO+AP
amfpfr4yVK/qGd7R30KMByET1hRJeEAJ1bho5Q7Bmi8lIEKU9JbTBV9VErQdzhQy
NNdS4A8N1SwB/PqEYooCTP3/tN2TFc+8INMUPXrK1doS2QoLk//bbVX/RIxoLBjY
YoZblRTkFpjjaf8AjJPlxbhBZ3Ggrr3OF/AHK2hRQzY0L93AJgn9fri4UMAFdY/P
frjR8f/I4em4zGAOKcWklhBKTUtvpMEyIzQ0r2WjvzR96R5yUdzbfn4Hy1M0FDb3
pULm6Za7nnrbzHcQMtP9llIz0yhx4L7mPXAhesrtCOshiw/kFtre0ycpOnnGkPLD
QaIfpNNXr3DIgi0HGq9EQlFF/f3bZpKQ2Cpful2XvOxehhJ4/xzijCqJy9Qfo1hY
2ue8T9EWA6P0lUEs0R5UrqDKepZBg5Ml50UGEZG7jl7lU5fe5+d/0mwjlzyK1Dho
UDJRYpCwAL6iHl0IjGJXhJI8VZbydHjP2Ide8N3u57Av1DjZl1LDdoko/AhHJ/oM
Fte4e40LNUSnkpUsgOP1PzqXZNqnZJN2TKuv36GOifiQPowVqc5m3N1eMRaozMEx
qUopYhYHxewPACfttGBdQ4WDLFb8Z4qlWyVJ/Rqc1AJXcsCGe8Vy8rcdpw36tbmd
W5Iqx4vhUxqb9n08QumhLRknj9AgAx2u82GfOPTSvXwzeGHKDOKKuDuyq1C+1BGG
q/Da0UmZbhyLsxoD0BD+7ViP3ve6IhneoIUYeHp2G5kQuAyIGNiJVLzxffss+Z2a
CuJuCZay1INKYMMKfd/8gwpxHxEfB0H7rnoB0iuns1l0aH6D05PtUAjHq3sFth1L
LuHH2Pw56dfr7dX/9GbhILa5JIR4GpMNglPHlf1b2wAkDm+uMp2tnCpvF3xFneId
RefYuJpBjcGKY8FyocExis5JBVszivBKrHsX39FGEpaOciwEEI07wAaBcmpkrf3l
MMUya4DO7rzc1g9JwIF7YYZsaWeQww3BWyK3na0YBJvOsYR8VP9mrKVVkWpoZD4V
/Ji+QBAtgGjXDLX+qKoXg9URW1omuy1M/OZ7LqLfdN3oXwJO/u6w+OgcvTQgJSJe
FgJysXZETO0VN8QPvlntTrNTPzlL0vtB+BWZSRLsZKSkwrPxwWZPR/LrMycwhzlp
BqZsWpCzJqdN+HT7C0RPphF5v55MXBK5x+dkIR4kKI6u4LULQ/3Zf0I4VEKgDuOu
PD/FEFbunbski/1cVlWwFFZQBD1CO+VyjDzx1zjUF3/DNym5ioCdAlQnJ+J7NTMZ
Ud4amT/RX3SJ+zE3MR9rJvC+FWkG/z5FCSjYHF0IJWgAEOemZDfiQnGwe7BRsHyI
I4QskK9Agy61rbZxGgRgrG+Ng/ksZlj2HMwvVvd5pOX7dgM/VrVaj0zHbkPGaPGT
kvy2hFfD3PhoLZTbkMwAO4bJ63BCspxMbL/yciGqrOLwdfXdVBZLyp6PueeDMKdr
bejyiQBVR7RTlWKm2ApsG/GsyVyRuH3UxCch9VCxJCeHy41HAXo3ZnMSYbgXM4Gi
ZIN+9asl5mqXcBbmFI0iix50cNJCMce8JuzuUq6il5JtoEf5jcQhJjMHhoaFm8+V
85rY+qqdBxpFA5bDIZH3m8lyahS1tI/jGxqtdheTO7fimSFu3Smjx4NWFaoh9+aB
rHg0VlhJmB3SnsPRT4HmbtyzsBn7vaUSRpi7Jshv5OSffEAg93nVeG3WZz0HMfK3
+0/ARHkHwGV0INV1RwFhP9Mg9qg5gVTL0WTpXAlHc69fN6wOj6EXGPFelh9Ikj6Z
5NB1rbqIyxyUuu5vh5KtLN6f1K9x3lF8vQlWVDKds7mYNtmjeEN8BKIcjQbNCLmG
kZj+idOiN45DWyCm9hjKY4V1oi+fkpqi9v5tIjn7GHlcTXcSHXq9oywNEJ5jXsHm
0ueeakeoNX3DRGzgdTSDmgevfYO2atuQGNN5KrRfPhb5pHux7rjsJMbKKLRAtczu
lQOaowH5UzzNXO4XMRTpe5JzML7lLGW3fLiAb0wY63umm38rkgHNQk99NWG/wqH8
WMBmTdEDYcUTDUkEuv7vNFhF4UHTP4X2Ij3DQyTk3NjrtnTqKq1Q7WTEpVqngcTN
xS0G8MDBU6oXDtjzOQ4Bre9Ode5ZsdJ0kZEhHyjP0nQ5R4BDexPUWD4BHvpmvIWw
0t0Lcbi2ZacW0QzfHtDalOPQ1rD8TZ2WgI/G+VsQjlXSiyfW112yJ9nTXIPVVlyt
99/p+535/YV+42Huec+EyEtTGs+UAuA4hbzHv68g0Lf2vUZpOdiTtfVT3hndWMcq
lFwAn4duYqmm5TZ19gFgK8d3HegWOqpcPUci41MvgB5QAF2en/xvZ0/4Zaid+y9i
oZD/U8ZzQW60a0KvK5Szf5aXINChV3I39u3AqgGUKurWhcSmxWnEG8Lf90tMqnfO
8FP5eVAj6u1St1IgL1V8YzCyw7BD8TeeT8hQXl2tBL0xf/nrjq7O+E2EJIILdBCG
5wFNc/X8RXTfzUFKFU5PgJBSv//9jlvz758Buagv5qXHdYrNPfJbCmEELmb0jknj
jcIkcoWgje04kI/ViOw127BI1kNO6l5APXyyMURJHmqa/L4+zniszI9ADlLv/oCZ
EHBS16JfFh2YQFbjUeF8OmJiYKCQqIZEXn9f0KTE6C84l6akHr7QGUnb2eauWtqM
GNJjmvIF87yUnksJkV3jCuJ7OxpYF8uW5U9nm1G2NVT33jvBiu1t2EBUvBbWspD7
CyvFI0ODcDsuYOuOFNv/2LIu+YfdlH+g4HawdJiwgbQ61YOtRyHLrayjEkB9FM7+
SAPFdF4h0HNKr5PyFCE+UjEWNOYOitbPOSR+ZOAEPUqGWLEnv5xB3xCzZue8rwA7
DNDN8XxSVcMBnvWsgvUyefHINmykMkov8OayftWLKJMDV6rkvJ66VIslZcC1rUgw
wa7bQN/pbcpNbwQiFYdXAdhooqG0humnCXco3jPpYol06dEJm46xwNiIiVENL8Hu
NY9tzaxqmMtaE8wpX3VLf4sMN5lAYAXIU3IXcQTsBJdGBf0yDEQaBPfaQRrBUZ0J
QH+k4vWeatUcgjhYj9LI+4mGoqlQQ5Cl3fXcbvI27tjiCcoPWgBGMNJ1/pYqa6Qh
Icy7k1bRKQSC+Ti5lsTcEUnU26hqfp7UrZ1FNm3TuInp+qebNPhLSxUy7uUrR8Wq
sxc+mYs0fuoBFVOrkrQDGf1TD7WWs0xU2XCFdDrjeeqnQ7hO2mqd5S0wmXmAYOme
5EOymtbBpNCCDYGN0iiT0jmStFTM4jyESKqfKe1qsasr/Yj7TG37LOymqglHez0P
egqEiJqi/40WsHG9fiUa4zd6bCiES7eSsHWXqnbmQx9chyEgWznpAw6c+RwFG9DP
YqC2qUXJ9ZJL+qVYSvZaWN5HRp3+icjBBXuOzOKcsiBcnCICpUp4QOI5RNkTE5nD
j5Rf5Qd6QVofeaflPzPlZbpTMDHeLqkDEI0WQHKj6ioOHjCmLbXqMZLb3lBvxKli
Qol6nWIU8x+i9UgnyFB3Vhyo7AUBI3vPCV3fKxJEwjYvosSRI3Li7mW4yRWOESNK
0WlYD3pFeWe+G3ooBrBjOmWNXI6Z8Xy0BgM/H97wNWfBwVlQOoN0KVSbQsaMEwUB
wLRh699senTaOg/NjPKW0mRO596HORrFXTHnNF13DihL9ULoUSiu0rnORY+dH6eQ
JnK+eeMsQQ75UOmMly43r1cfMqoBgny96oAy47GwgEwsMKKUvJ0xLzdfXulkSUIm
SxxkvGzSxWP7Pgq9bsJWrqS8WsVWNp5vXMDIEzrkKjqVwwHbg5VeIrFRVTbO2gsv
jEeEA0MEml11n6LC0zqkz93K+aJB5K0nXHAKbplnvSmAVnh70q7lpvLKYf2AtVXs
Unnw1OWCOzxNX/chHLYYiPzjC+SrmI00yQunjZCYI0iCmIqWpNGEqTMthjZTsD6b
tztF7Sugb6MYDek4O3pXJRlg63NiLzlf6Z06R6c8iHcv6tetPkQpsX/24aPUHpcv
dBVqcw8SLHNeYrdB4T1Vo4mL6x5WrU6gu5r65cuhQ0v8GgGL1P1robxSmxCY+7sh
l8Q+3hFzcj1sWycOR0bgfXn+HqejP2DVG3fkhZMLKWeJUuzMB30ZOm0ZjlMBFKNh
gZ0UtzInDX1tzrkMj/ZVG3NiAIF0iOngOH3Zjti7IlrtGFK9MHKsP3ApHHt90Pvj
fsyQLMUBGI21MQylsrxxeE1qGPktp2BOZkTYgUcCvAunqz+N7HdNLDG2DgEwgby1
9RqDOmj2ggkdZFKCQo8UJBsMFXODx15Wgi2EhruSBGyAb0XIG/NlhE8ArwQgwLLh
d/vC5gi8g0F+79auGGs7e4pYHUXiN7VOiBjY69u8FDxPVI9risYmJi/7fFwYGYfo
slApQ5ONR2E9+TnpREbFTWCupYWpwglRRu6wpMXWkQw2i5L1uykAz43ndhyfJv6/
gWWXaTwb+qdBIvaFhq6890T6vbcpzUw54PUxhd+nuYIvO7txQekGAKqQrF8cQc8j
kKtrq8xhbohBGzr1C+IvG/Nh3Y5Fx9iiy+7M/FLD8/va9e8vpMscYXzdhXI/SDrD
UF+hO9pXfVkoSZbND0tCaKLagV+gcFTx5jfcnKUlKHJXDTz+4o+ehx0tmExLnwUt
uR/esRe9xPWAsMHJuqh25HTV+3bapm5V6nhqn+MZuMjZJM0HgeQFnXYJ5NG5+htm
hpeokqXeKQqWF11nubBkS4E+AsEaXox3+CtpbIUzU5uienRpy2z5xujs4Dw8jx09
bife9XJAX8J7aif8U2rUvWkKycUecK1fMIvYSDr5OlS2tsH8cKn8uUop/orlaYBF
MZjsxhtidyGqCmNQFAkvtphT142YFK8z90mz5/eL2Iw8PNCNakDYzFsE3ok4pxpl
IC3+j/e1ywzDu1BgTIzlCmaKsxRCDe+c2PxbTiWqg2qxZNC4NdTlPZVVRy/DtlFP
XT8WagUV8tjbllMbR3SrW3N082R4iSYygGcJ5MJvdOlUXRRRZh6yf/Nt8ia9kMGw
+AyWM/8IBKQGvCcYyR+z3JqD30PptrvC0pfqQh8nR5/gDW/ur17zuUNBk4NYSJ/W
vDHhcA8Mi3VOUI/PvjYuohD5xNJyMxuAvuA+6g/PegKQfZD7b61l4xaMEaTQHdLb
WVljeYCxUPUlifUQrXViE4sgLXPTi7cyTqoW4vXfNAEIMncU4TaguWvt1xtpS00Q
LDO6XtuM6Naewduztf+FZ7kNsjS3hORIABsHDfFLqASrJi5NIHQg3fFeR+Gdy86h
irybpWlxJZBVmj49LKwcNa6oVUe0jG50Uz47qOvhnp9xcqCMErPKSuPWU5mn5qBY
1LLzEZvajhlQtltEQmyJTF2KGwPFVl3Kdh+AXztYq78E9cXR5kaVkecrHjvTfUjf
uS31OeTClFpmTtZFZYwnyZlZqtXPufYTQd5ZDMYF0E15XdDQQfaZVWcyB2Xf5BUC
w11dJ1iKWNvKXTtgJJyt7KkoD++Gw9U7dird54cNqQ1+7QTw/jmG7o08iLP/uT9p
GdmbwT8tdINUy57OgpmokXEgFhi7SltqDeZM4FsSqpH23KCH5UDyQz5XzsEzr/Rr
UEds7FKrblhZcvbCrLQNEWtv/wEMm3SI7MVvnSbvTNs788a0P2Mx2d/b7bwyDUaO
YJLFW13n40NRsi1Gq2wltxOm2xqHLrE6PAaK+fIemeAFGIC+qYXiTVmIy8HUK5P6
/zEmjJtS2ffheplNJntiTrBMe4QBzxernkUIUd8E+39gpcHGghETsfrXcnBZSXnD
ZK/2j8N2oSTh2a830eZLr2TvAzZYO/GxZhBlXDP/C7BmhUAw4bal4KVsMqGBqcNP
GwE2/xLH3/JcGUxHq08hbtBqWc97qj9VSxwqjYnWSPSyMm4cIpvAMM5vP7JjlGax
CXhSIbeDuxLd9U7ePfqqclFPMKLe9NweISH+f3q3xdnhbc8/1ZlARfMB3jyARB6e
KEUg2dNSY67KbmZxMItpxrjFD+l77L5ShzIZFGRYDDfA1OZJLfqVabZfzo2n/hX0
Hencg/M3g+fye9UgtC8qbgo5K951yezCnumIYDxjlr9EknAhjcJ5/V2Hw08mKLmY
ivLeBIOuZEF3j9il/cI+OM3gnq3gyUGGli+Mb8SDmS5SOEH6Cx8rNK71SZARhwv9
6Aauc8vqqiuA8i5kXiTzRGn9K6pGYJswTNNz2UFXoxfwgz2fqUaHVTR1q9RRWpWc
id5R4p8v5Dwhi63tqb6QrT/2ONmfUrVNF73K7GTp63QO2+7IKF/iWVwTKxVG5WHo
wosD+W1TBda8X5jxdYGLr2Tme8y2lu95Ay3/Ns1ru13vPQg/1ctsx4zatERRQwxi
bRrJ92tO7XGLXmY+ZFu9J64xpjUEqtVLYuheloFYKpq5ptz5KnkAnBSNuM39wVuz
KNB5YiWBeZI8XGDxFSQMmuPpsTFhQQRgn1mbTcVLAgP5ogar2YKtKVcOubIGQT7y
XNilRmqOFsmE3LGCblb4qgrvHps+vDuDxNabwC1zftr5qepPW0CRoDgBurcPmixh
7bHnyv+Pz04KTGazlfGFFeYCvECaPxr4jlN34BsB6FktTuUcuAM2FcazlFmyjD8M
+QagBVBGvZIqudkzSWhwRjwXvEtsNZHi+QywsMwn6zSgKW1XPcXhHGDah3ejasO6
G3IVFd3Od3Mjfq1xhgiWLp7lb2AbYRe1BQA/arMipFYD7eogMppJSJdyH8QCpqW5
HYdDIxttiqRj8GpDiX3Qs6K9sIW/HBWfAU748YQ6JmALRXoSHMEjyqbCT1QSbAly
CT1ZiD6D1Usm2Qa09TOrmXJmEgedIB957xj0J0n/fn+R9HevNtpVez8v3+pYqamd
4rln8Y+3SRif1nYvaXUy169+esqXzDuheDbZeZLQzWRepZwX6qAVY0RE+KP+3LaR
2/+aSe3JDuIVjPNQac/mrOAaA3VFmvkaGq++jBL1ZGxt8id7xGXON+FdYP18woHL
JD5aHoPgIVoIetai68ASk0A3LjdH1+g9aQwKGvmJXlAcPtp7tkAoyfrC36EMFqIW
nwQoy3Pb1yo2qXeIWMZiHTIjXoYJqi8aA/NYALaUYjIiJPLRL3ackVCEwO2uh7lM
nxw2J971AkcP/JPVQzt2QzGgz38wIrcW7jZ6GaAMEk1RqH3pGRQOHOPbGZG/YPds
tstYqylwaUqfott1kNfZBhd+gczEJqpVnyu+WsA/E+oOFcRL1HwpvgkEVebL6C47
ZjQycfmx81sJyp5hr8wkhryk/KBWhvQa2snvlmILebS2rQlvvRzxSuj3NK707VHN
MFPq/uVNkxe1bBNQZXhpFtE+05B/6qO3C86FZ++lG/+ysJOxf33dF2dK6fvDbJHO
B9aVtS1GwL7axPaG3wfG9XU8xTWzxvCkiKNjQP3wnX3UOKucRg4kJjau60df5zyU
0i1IDYoWhe6+Iz9oW2qLFCSPW6IBJlbb7wJtIm4GLrEZisZ/F9KSms3ezaGIfyZu
FbuLQYkW4xz6olarJNf36RZhfGT0YCnXu6iOIXErRAZ+ObZiy4FwonO4SCLTmUzK
ZnMoJr4DW8sDm2k0EJ6y0WY5hv7m4wBqQkiNuPx24bu7ByWajHUZOjHUXNsWwX82
6D6+cJotoymQOvAFzjx2pnU+upiX6o5eJGg5+ka3h82/ddJ1hS+nwRlP6zTfoVFL
bk/X1gsFIPZNjZyncbO9b+salP4/bO3jSKk8rfbu4WN2+3YdBEEIpaJ7i6JmcOvi
MnBunBZbA0h+SX46M3rM9nR0PEOcQJmVc3RfFMM9cyPBF1oWghSPEC65dLS/b0vB
KpcRj9YAEJOkCPpfx8hz4yeB4tuU9T9vfjdvQUT2ZbMzxiN/0+XsK5DHAQRu1u8S
JHyUjF506A72T76tUum8pGVp86u3R4SN8k/qudeZw2t9LBZWASCoqwrAvj++9Ckf
0IskAMf6EjpeJIsDoMpTdC6hW7VfFrsxDz11SJgKZNWlP5TEFhDHAvgly6k7eom2
U2rrrDpNfayLdZMHq9FMgyb/NkMefYq7QMzglhITUFTu6qq9PIX159I/26mtF4jP
xgU1O1KTZupeV3AP/wd5eRiGZjwB8DCxfjNQ0o8sv/Kqd1bc4cOwMMInbnZ2iI4w
ZgzKGmqjvWLs4J+ezw8KgHjkVYGYDd3XhRX6OcO2Cbt/l2e4oSL4Qd2oZJKYVN+L
JRBSXPnMahwpmtSCs0HXGHFkQvx+n8y0mfNthXjYXTLFuHjT4PXlISxb4aFZlQGZ
z5+FsCc0am4l9zIJhPWiBq8rbw3snAL7bpBSuTn4D2gGu11HHJJToYdcsj7PV2Ib
i3RCtlvsbU/+j4Um4NGvkG5YCC7wxmGhcyv0a8Zk9HPdk9/eGN+G5F8EirO8S0F4
TGNxX4d5CJhTKcudkkegufzxfXfIzHVX2BMKgrqY8IQ3v3eTNgLTfaq4JOVU5o7e
p+D22mr8lHXlO5bPf0CTDqzluiUxNd/iOjKOVKIuyDK5Jb3j3d20rf5hJjofZnvL
knJV5fE7UQwUDjiI711abE3xn5qwnRyHSs4R7wHBbCXKUpGiwyIIUtCxgSVaKoGf
AcsuGMcy7oJNI2/D/qGGv8u96dlPHngZp+kPk6TiuJ8Ix/ciYE0dvW51FO5kvpz1
carXqq43jOeSmxfA1OAz5OoitcEwdMaP89NJgs06kkhA2Pq6JDKrwcfqw/GMxkFL
itfQz7vKT3BfyXa5v5x9VdGtaRhkyte79kMSBtQ1/vIQ3Sb6tYpsRZ7hTiFaXMqw
fxxQttOJov8WxapfKd9FsplXCSrW/AsavtGWlhAxDeYU4q0++p965AMiWqunVKkx
8VK/cc0/dFAIlIzXvEaNI/lUPLpYkrt5IofexKrKHT2t6uz2ERtYurx4V7uS3i0Y
b7d48ti8P6X4q01pBdNRG+pTUKh8PbzhVKBylRo+Qu7iwhmezTNKY3spdJ+tpTVp
jOir8KNk/v31QPswQFWEq3AOzU4nt6qPzZ06VYzIk3v43d3jRkkBHpC5V7CxSTLg
7gLU3KfLzvzAQkP/lf+AJ0uGI0L9KTGoh/9mBPJgq9l1TabBA5DgWbrEevx6eYDj
G3f0G+jEC13JpAIGUtYnODi1CBez4IHdDimBkWeTPB8kbHD9ITd10JWI+BF0pneP
X9duiOCcN/I6OVfXqF5DF/PK9smbSVJMMrOUAmsLnVIxvR5c165lEUiHhqSpcnG9
SE6eD/AiC/ZCQv9FzpodM9zEA8MuiyOSWs3ItymnNShGyME6vo5hfjs/Mc8AKDER
9e24FR/J9QDg9aJjbJn9cIvc8crPyXfWDjrkgU7ddJ/udG8aGtCEaXO/LPtmTDh9
e6s1VDhcaP6BRepJxta3+Q5YAE7p4B+c6gSvBKNTJKBSQYDShZFhm5sZaCJMxSAv
M6mX88cvmMXbMW24oISv8Dt8cQb0qVA7wW1Xcuxba1+ifLWD7kPvvHpzADG108n0
gfbVtSa5mqR0jLEfCw6wSEZOVi0lznIV8Sf7+LJ22dexChCvdEQAxvKkTpqPpBSD
Fh8yDQf0upkSI0Bt38tmTFXelu79n8q7npfUw1d6vzvH/jgw0XPAX/ePlrHDHvNV
7o0e7eOq6m6fUP3lgGZA+FML4F9NgmYR+yhhm3hxS9aqWf3f2P06mzZoKwyRm3Us
su91YY5sJGbVoad8WVYcSHiz+/sX/aYWTAaTe1LEuPMEgCe4GEvcaQENI4lKSrL8
2MbFCSVCcTJFAxXqWDiYO87ZcD7CkyF0Btqic1WJiTAnHWUcdgP8ZZQpgGzyl2tI
FuKLcpbayYDcB5qRITDjucAezS5cCX/DHMhKIReeQP8Ssf9KXh5qeXLAiMI68ee4
jsSaIwqKQsDzyM870DALbw2fxY5COS9c2lGZBe0qAE1C4YSUyJRioRaVv2PVEvWu
FGFt8QCWuNVMl8z70Y9ujNOSF3b++v/xxloVS2oR81FqWZI2Nw4GYVQSUa/ekQoG
S4DJsVVAgbhAAl6Fs/rf/qLYZ+SpeXdrx94WGVUaYj44BeZNzVTluu8AKwrgciuB
zAXPGouuhmAfpkZnba0gXwLY75nYY5wKaeR/12Gw3ZXMzpc+rOucT4hcoV1zAlWc
RNURseLMYvg6cUNlpjA9KYhKqB1JXtcLJv4YhXixc3b0Bx+xrOsPjkDzl5DBZYwI
zk2YoZOMdQJLSm626lg8bMiciknGnTsjNKn5g/RPfRriQ0NGzLBWYlPI/yVGmtI4
uaZd0yvsM4fsDqn5msfX2V9Y+0I/x8u77kH1czVreZtk2gG3Zq+NSkaKAKKdPKPP
AbWZWsgGWOoGyk95NmhiivfvqywwtRmrHGx3/bLDRQyfpyBkjcT9Ifc33bAlC0ZZ
djvGqulOqK6mOh6d735NsxCqqkf9fZJL5O7nWcELZCXueWdKTnnZmOb1NFBKorhK
SQObTyuSCF3z/Ed4Tthk4Ko+TQoRIHuWShbjjdFYG2u7gvwqmQxNJel33YUhR1VA
Hwgppl5YaA4DaDBV8cEqmwJ+0q++EM8dKBMs5LR8T7wE745oKqQbhBbPNTQSxhEj
B/P2YKp5Go8DKQSZy34NryNEaE2xY2lLxp15SglG7zbfeJN5gzD7oj35Z2oiRBy2
XHouldBs8zroc6oQlO53kqlcMNMGJupU2Z/+XWNZQkUZ3YaB8yMFiHD0mMYeaOMT
Vak+ix4OrixUyVypyYbno7OmygHR3EVyHkpzFoI59FiQeZaO/6NIregHwkCPZXOL
O9Er/GfGvYZNgFBfjrrjCuysm97K13pmcU8aMvaL9tfZeoSo5bJD1EezWhC9+rCx
lxc87q3iGabMFd853Wp3C62TeCHJPaBhUzOREDLkOok67elgReb1VNZcZ+Vtb6AY
/mLrFEtdGVWvY/K3Z3IaU/jfdx2qt94mVsUncblkS/urf06GCWnR/MDwNE3HdL26
DrPilwdfdJrEVzQujC4MWtLlpYgHzFGNtxnD9dAXf2NODZI+AGoW4hR52GNzggGi
jGapNUMYuNZeDjbatUxt4EaGuvFhQ27vVpdGWv4yTKz24Hc38+oMrprLZoax2wlb
/bUaRIsW/JsumR1nzba9iiLuCFpCiokH4pYYZf70iexjZzR5BkB3E1cvcq5p2ZJo
hiym81rrvjOOzINquAGkPVTixVx/YodQ4Eh1R4Lw9kQ1bX/enCcfAu63YPYjEGlU
oxBooc2DMNFgLqRgi7+cIqKT1OqwK8aIcNvjdS9arbXYRo+3SZZ2sOJCfpXpLPoa
uZr/1+aFMnTmDlkfK7dDkKNHbjAIRRV5ONkUiDa6goObehHF6es8B0ASFQrVY9OL
6SphaSqoklXctTnNIhAX1mdf3RooFVRBy5I6TOc0mIGSmQBNzum+yRrCzKFY4iwZ
FbPXNdim3eqZVy0v/dZpBGQnj6IwJA1+SyaVH7JdVMj3ZJyn3aLRmNFxBciaPGUK
gNe1ZwJI/AJKJwlmvTOkTvIpfdAPgX71+uK2YwnJhFgDliCUZk9A5C8ewYfla7/p
B2LmoY6Og1qmQHLfPigukybqe4RH5uAmxxa7x8YL8lhdjI/rpcvG1X+yJlNAhP9F
LY4ol3O4WQkh49Nlxlz2e34DzrC990d4vc4vsA56jKLRrUfKNY5DzuK1Ce5nOmtl
UQAlWMdTDz0sqvlcNIubrLlzexeQI7TeiEhQ8v3lCTTm8Pbu3vezcnfh97NdVIHr
QipJKV56XaPBGFTSKr5xh8ufROkiHSov6TFz1b4NZW/xk+0AXpGNmZdRzAON+/0I
C/l2QCavOWsDNmmLXjwYp1hapZXYzeOYo/aLdIMukuwWPqKuRwJ+UG0hwZP+6BoD
JjcvvaXbNvDOws56dhPkCxxNWeAYoh20sMDUNxL/AyyJzuPmp+k3mlGy5zBNVG5o
6lnfDex1G0Kv1d8SXj2EaQwdmO0UXF1YZiKy8BM1yeMC0vXpLA+rcRbBrXSjYLYI
ycD5bPBK4QtBCJB/e522S604IxaYLwkv/FpqDQOVWlmWQf2JFWRlLYydoI9wsR+N
d+zjfbKdRZUgAJWXHaXg/bAUcI3GFl2HgnfELgUNrzLYvO46grxYBAwHxSFBMTkb
YMyhQ8adMNCe8jB9HcBMovIkjTRlEQEHANjWVxicMn083ONQAJR+tHXxtmHAadJB
Fwm9Kf98yIH9hasRybnReCy/ov+o8sYUJBmXbeGk4e/REk+Sppua1sTLNpyAzYiU
PlL7GH5MNu1k7iTLWr3UkA2wEVui0vX92ILIeqFxKkTPHjoBT2W31waItIemCRq8
so6lFaueIoNVs/62w98ZBNkwNySuA2JcUOrH8S2zDsU3i2fnZ9skb5v38Dks0NCe
6hfQjtJ/5nwwjUuUhqJF9umSurEXbVpz4zMXB25EhjYqX2mpkDO87/Lz2uVd82fB
qWMPlVBcYSp/944MFlGq1Js6XF5QLQ/LnlKKUWY4sbwthYfgCthXMIxh8S1MFTuu
3hbDqR7oTn8MlNIemH9FmpSie7cupvVfoZwhSP0DrcwKbcu+hs41So/2pbyY+3Oe
GoMshbJXwU7bfylNJeFCxeFpR9wvPtZ7L2UmnlrB6r7a1H/mnlK5ILrtlr8X2ntq
5wOKHahVd9EkVSXqh9Xzz3tYXTJtj7tSwBcIsoPL0L4sU3qazZqPxFHiDz/zmYjA
ES+GXMuUhmvCcqiEvb9Q1Omcb+hcONZwyW5JN4wn62XD8a62eJuWWalvvQkC2G81
iD9d3RPSvxjEQrkzC8SXDE2JpvtzR74B54WQBae+ab9tBapxax9s1C20DqySlWMZ
+02JkwfiIFJrwrJJE59JAeOgsM7TWsiY52rGZDPu9mIujz5VHVrHvs2SwBxdfWsU
Pm/Um4Qb+eQDmBfCIWuGNp5btiYg2s3OmfiO/C9qRx7u3fQlShlAN0Fr2tD5m53k
h72uM1Yc1t5IoqLiOMQ9tCAN8jTYbPV1E4Bj19Hzf/51Jtfli/sZxwW1Oon7tM3S
iZVr79ynshMSLbj6NdyWbJ+w3tkCtLCskYnpNle+nBNFeS/It6ikGWhZQf0AlG1a
TG96rWdSxxaVFt3O1r+9WvUouvBlleQaEIKvBf8ZvSeqK+bWuNbsmFBm7PP+2xn4
7yYfuKwtkV9FREDXJqWMuI1z7hW95uZXB5wTEnCKnFFZrECNmOqCrKjsxzPCSimM
67dE+uZSGHHK4CX/1nxvz1J8Gb0YpV3hXtAtvnO+ieIDpx65zt4HSIG7N6hWP7AW
3jRw18mncmLPzVE/fp2pJt273yy9eSPnDfOY3ReaZjRAl6QwKf7kblkXJU2sR6AH
XHPFUPBVKyRKaWcHy7FXIsZFFk1lFg1JjNoW+pU6eUl+VB7TFsxx7EPMMyNPA0eu
vuy6O7N28zHRqx+8MlRu0VgNnuYfHh+WzpCIJpaBqz4pvwpblh8XU1AgeF10BVxH
PKL21IhVmXG78kFDQxw+TRla08z7kKo8CUhr8sPkdbxaY6sZO/o9IneaPROx3jNi
FUFGsGIW8R79vNfEU9bF9YLoGnl/H7I0RuOJz4/3q8Ko66ogp/qa2xdCf8nC4LJh
xmmuzcicjpl7rHdEIOEvikf0M6SoLN3Xewq4DYP7WJcMj6hKQwM9s/cGGKMDVhdN
94rzQghUJu1v7dMpD97w6LJ0DGTQZbJZamHufCIra0be83RXkq+rR2O4endmFqEV
H7Xly8L0sFRi7v5A0hH6ZrTDnbdjRtZbD9KlN8iqPddTVBOpFvYgS0JOM/slHfMA
S2gRkOhFt2wxbg5IqNgwGGSt/m1DI+Eb7SeeWrCYduSCkkUXkpSif8yeQ9eCbDKI
K1BnlLLu0krx1YnpLPySHhYfvTAQFgj5LGCYLlf2WmFl2QyYBqOkRD5hLTu8cwY2
n/gA/BKCpg0s+RR1wnn4+dWUrv9fV/KvZpzP2jxn/8HxNsvjue0WOa5UtD3A1t7n
JWbRDVknaY5Homs0wnac3Xx9y1AZSYtUu4tuBKF7mmVOlwtY/jd0gxC0LOC37yRr
uNuayT8yPm3qXP0CgI/iUsxlQHDxc6E5TlLugwTrf1ffxxl5rNl+MRcDtUWm65s9
1Bgja8Lv1XIp8mh9ujo+9Pgblpg/CngokqkXVYEflV7wCFDkTYLZavdqjbI9EnDR
mF2Cq4p1KcwOVLvUbEmf+0yxDixu5Bq2PYVQ7WiJQItwcHkVuTkJuDN3H9kBBMng
+Q7Oac+kR4KbQkkCIHsI6z4c0fTyOfnOWgs0hHJ6BV4fyIpq+AU9raB/iORCVCUS
3uoCqeJ5sVp87T8hSbnItY+NBRzhN3UYyTnFo3/f10i4IrqXNPF5KqgI2ISO3WgU
h+ui9u+akhh99BGRC53GA3IIHLk9zV4ybWSk98NnheyhmrG03kSWHmXWepChWbtL
ouREQV1Txumv7V8MV/KNxS7XZtHxCtZDwSgAmGfGH4d66XtVajb1t4Nz4dELUI0F
EssKti+x9idgDro0DGygjrYV02AfDPetVG671Z/1VN34bqEV21IE95O4/E1M7vKq
f3bUcd2vKmjTQzYFjdbwuRExLRwtI1Fq2SPYY/MzjGpsVAmwTjjWzR5cOMvDDIN0
PL38EhqlwTpRGGx7I3AZJTP2+pNjw8DFRV+TNbUxi7SgiDl6loq3UchOXB7rEaK+
VTKXu5SlHiCKnf5UjGCgwl/XBahQQygwGnTe0pbtXUK0QzmAmxTIpHpCG6rwXO5s
pCVvs0oLM2/OxGeZa1RZD4EC2UBulBKz4WkWppoPZAdcdKVOAg2aazqg1k65yUjE
S2FLNpj54lg2tt2euEik6Hsdna0dCQf+ie0wymQkmEBu36jKbcPasNHvQ1VufGAH
2Me44M/bg8YfacFkbjfgAN5Q/DfYO82X59dvRV8InmrXcb3MTY08B5ViGSvqdmVG
vtFBmsNYd3aRm/tcZgigEv5ZGkA5xPyKJtEhUPjkvqlf/bub9bOIAScyO4Fpwiot
qsBbAse4MyQAQhTIdp/VJWxazd5BEvnuY8hBEseALzhzty4gpgyZVKJfRlj4JuvV
jSyYXgIM+vGCteI+w/ihG1nurLVbW1ewjiA5pOCNNRRRLNHTX/ZLt4ra/tDqooDz
W59OS7MsPSVruHn7ggFMijw7rgKOpTkYStg1J0SlKebYn9QJGRE7aMKMo4oQLo0g
LvSEa00ByryGPgl1Wx9quA5POD2zbhDFBjPcv9EatOAI2hfmC8rVwHHfd5flDGF/
8idzx/rO2/EnpMBhmHDRnyPjH1FO7q/saQTEzB6rkp8vxQ/tGoIz/m0eY9gTwpHL
nwVhHSO4DCtWu58QcYIV4O0CnUpxkoqgTvkGvbibN0+gct9oOkmyepEw3xQ8fb0V
yuftzPFVzsoVclH1xLffHj+MS+D1ZoTXmNFEs9YdkpAalZEkqyFNCQ1P40JvObam
+m9Okg2g3D8y/ttYB06+HAkSaUzKBcl954/98Puty25+zNoTrkOW76HqffOJVY6H
TU9VSQ+TfbWXdRIR2U9GijzCuHdcuoGY+lIPXB9EOPpizFzhTEyAH7UI7pcSYJUu
yqajcBEbMiAKt41I7LM9s62k9SCy6ajMen7udAnZmvyojR/QlMXf9rneZVWVAsxX
BfsXyXNCCPP5TVf91A50ZVstMhU/+qRX9kd/gbs2SAkFzSfKqHoXQI0Ci9h/oO/1
S0S0/m+us7Afo/AwQvC0NPHlTrxIvx/ANaAKNpr/L6ura6KWZJqEfwbVO0VGGVMu
gMHEFfLwdJeGve2Xh4MB1VaLTFh5hF+h2aAwDE8lKo2PMBZxsOUT48w5a8R30pYE
R+O5n3kBddOYILY5fWVU7UsEMEFQG3ZLoP7AhZJwtWRmjBofKExVzrl+hLovs5sX
eoJGvM2kT/p/ZSU/FF2xFv4RHgtF1WOkp63NF3UH6nldQp6MNOA8gDCgSda6APgF
fKoenNrq8/qXo6vZEZFooFN9xx+bsBKAi8x5iI0LmywkyLxUJfWrz/6sD+u2MlnY
R24F9eIjrepfvFoqSEhOHNtudEL+CMV8/sh5nficVz2OOWlOV4jVD8G+LSQ0CGC2
foiRQXeHeeZa08AEoHOqnWysSDZ4w8qgppVm7ThG6mby4y891br6WivZVmq+yGeg
jt7jTOrya/DU2Z/5XCGjto20wqCIKCmXaiy/SK5753uBpEA5EK0mko9eyfCBy5QC
PGq4xIHeeOjKvSVwYldirzhhtTCrKaMQ1PEAiPD2rX2LCzL930uU54Ui64XhfHkY
VtG0ZKmQjdfJtotzhaaB7OgEJZXFuVC4dsq8jKhzT9XhDUuJbjwvxnded5zfeXJP
fh7qBCcXNzep0ANoDvHg87vQ/ClWnJLEhytdyY3KtVv9iZwROLGqI+gTHCLTdFmX
1rVin5uD/388eBfWVPs85rgXhYYpg6ew04wszSJyf7v+DOnk4RlM+ZY2fUK0DYQp
sXHTUiJydChJzFH9qH5KUR2tjS2pGsKyONhB832Br5XIy2PLHjj5n8sJbLWYch3J
HrK7ZAyWoNJrpj/3DG45O38ZItLz8aqC8hwRswKYwBkehuN7b68uEEzKpC0V5SB4
N7Wos6rtdkK8wuXJxRnmKC7ce8vix8pq11aIDU643rcCxaf4bCfKiixir9gwT3Rh
hEpqLEN2Zz0iv2KMfSpuyn3IlDsoNmlkOCfEr3Ayf+TrMODirAH0DsJeuMh2rIUe
2HWwNCMuZRu3dg+9FqKX2FPtjbShE8VdcSda+bISoeyGCkT2gTcrE0wyO9dJip0C
676yP3Zhz+6JercevIKwscvHR62odClD8fN902aIg3kHIYlvPKYNS9xyZK4+6gog
iyH9WRkIYWhMJVu4c7wX+tp8vpT+zYkC0NdXDlqFOxsbGAv5U5DDtJ6n9pHXxUgP
fSD9pOynIt1/IFIN+OAHWsstTGBM3fQ5aZgSEq5m7/Kxkpw8K4HE+yZ3G/5D8E2F
oz3NC5ySvijoYGZYJZxzUnTPsJx6lZisV2ltwrdcaESSS+QxGxW+KBEH+nzgBis3
ODciu0ItH4uc0ModpQielUv66vbqi7lgdesrsIBUrxlcgiAYz0JGuncnYFa+PoSL
QusKmIS2ZShcROhNDX0UJRr1zPQdRGMFSnCG34VdV4cFuyekPfGngALhqI1FLxjM
38CeSCvmMUg9PnmUYyAOu7tchvdbXKynTYp9KREILPBofFm4/5AKpaBE+vn2FagZ
bv3vi7OItLeJzLU/G5LxocVHJIn/5+/kgBfG3ekwIXNXLnD8ATnR1W0Zd8egSiI5
+Zt3c87SXAWdbfMGv/EHvszFjNxF2nnH5QR158Ma30RTB9d4yAxkRTllqZv1cIv+
YvxaHefI+pF8AWxrMEvP1QIAhQl3/pebR+NNaYZ4HsmAH0cdCqYWUPUgi0h1FJuQ
Kzk4At0l1+mRc7nMGrhyVT6EEbeNSdtYAN+I0uZP0CU/0lkAqLNfHbVVlY9kD/jJ
9pnXM+wrcmG2+NemcBqImi9uIsVOWLrzaXeVTZIGq5uR+VHutTk5Xgn6UiFWGnMr
YoTIP++hTfLU/uPGrbUjCo3M3IhjoLXH3ErZZb1T+Z1XGxZDGY8y7o9SvQpg/jFE
52wwnK5/LNq13wY0+/xhmJoaZmfaLd2xb4qah3HZ71UinfelPyyDcOUSV8nuZqqA
wRrSgOz+0HZJJvnmA8pohdAcRFDyneYov8jqd5CpxDLO+2lfO+pl7HLVDirzwa/1
gmqRelI/JzzmLKOFGofgw92v8o9wKaJ05F/CSKL1SvcnNnlezkxA/2znGobI8pAt
y9BtRQom0hbFbYt1fxPyNXUkiMCPl/zlyYULtJIXr0sAFniA8cqbZ4Kko1HaFGsu
hoIWws0hYlUo787ler7UxGJ4HF2Z2n+eoCWAuQyX0oYENB+Gy3RCG0QhkJsYCsKK
jkpQCcNeGBZ2BK5ich48OHz30d+JusPn8DPuYTBi9LkGmFld25ypaoQvSL2RhwTQ
uo7seLTRUsxmu1+gu29reJl8RXfXy4sgB9RuY+vUWbVGqVo7QZH2huH9zG0xYSEA
yJxZjaF+uVoUTga56acuNl6T48N8ls6e9Cn+I4leva6/dnn6afNVCakQeoVtj7Y2
x2lpMrTQzk7luGFp42ueGNDg4YVvaOhUtYQizsmIyYZFsgivViOt6nh5N8F139cW
t0wjGeeQUKoPHRkKobm9AnDrkU73eCcVQ+Dk/pexVxEDU7zNGvowzj6jQFAF0NEk
XcLV6Ry0YpwZHqT+9okeyb/yma6jQSQGNNKYysBzdVDlP81RMXtmGKM9nySkCpBn
hzDrtjXpFqV0mD1rvW7lLy/SaaxyFd4kOhtHy8p8sl2EoB99xIt9ydDBpu6fexoD
SFAxgN3eJA9jVSU969eft/43rkh1lshSJ3UQtA04JT4xCRWjLI5bWy6dgZTc60nQ
+7ycGIvz4iMvBXvsB+GYwDJGIzCuxbDrD+7+CuAdgB4/ooQWltSAtjPZCPetVoCf
7Hl6oNebNFtibgcMTg3ZT9fpTeAzZb99uwww6lLEbLUkROXF2+b8dXSamA/5Eget
HKgRV8pEGybdc3KAvzlS9J9dur4UIMvrF38JLPwsNXTD/HCwLb5cY0iZZ+lWJ4JY
S+DMb9sm7FL1t9ip7nfiFmboUo+/JeJ4gHu4HZhwn+B9GooIyGq4S6jSvHFgl94t
+Dfs20JWEE94j99gtG/5By7GobxEHqIWu+larpCuRsIAxZ3AnQxJEXrECuwtbS9u
VylWkn4zKu57yammgELvR47polsgQNZ40DvKLAgXl2O2lHcg6yatg/T8UMVhpV0J
Nqr/sUOViboW8Q5MYu/q8VpEwshncVlV32S0cwD+f+A9hNVeXkD0iE3lsyQ6mtWe
IRPLAv6EQTrcQhINQ/ueD0yBAqyFj01YeOlE+Z5LtIV56bJnC1FHd74vR22QLx/O
LYl8mqVxL6yXduAJTiv84SfILKuFT8IW69TqkXSqJnTNv0BhnGkHrxx8W3PhtSL4
CwOWd7AZ7oGKH/KWZ8ffNnNoJ7vTN/Mrzpky/BspoMDdpb4csS85oOrZiPq+Xj1I
+CrCXuTuQnz4enOJ+IYIjOt+DMK6YM/DiTTdBT44YCSA50UiqL643M/5ZKiGw/qd
PC5+V7m/GO+0qWK8lIE/HwHIM9qU9nwD1gfVWUaqpACGhcZ+2IIFy1OsZudsYJdW
70VWUZ+F0ijl/EsPukKKp/qsId75ALCJAPegdcgkLq3/xksEJRYwjJsVqUwptWay
oHY/4FhvLGAW9qMqRcdU+VympEzHi/kFmKJIbJ41vUY+a8YcRtEuG+CYpoG9E6jL
5peNTC+2LoZSeSfTJ4hon1iUkFK5kA/jOlxVrLOQnYEZLKN8myq6g7Vn3lsYRO6R
aDqMN29H+t4pt+rmKLSXK/ga1pYvxcJ9IPkXaOHdf5Is6hGIDsqZoMYrVoV2MPB4
Z1jfDm4dxyDiScbKdpBqhr3wvMcdOpHwOELNnWXzJTF+Jw8ellKGjX0QzK5HLzZJ
Ylrs1tpWz1J86A9pq2CJHnXLzLFoc2WY1aHOK1h0TBwj+G05MvdDFidh1JG/aspX
SmjGA0b3HvMSYyDh2dcYNLwlYke4Ctzy/idnjQzJpWJTvktfe/mKf8bMDBFB7KTb
hAAdJF4U3rvzAj0fNns2tonpaPVtGjX8Y04BXasQVA5bDx+I6bPzW3fRWPvGc/qy
bPTCOpT5TY+rorEimV/vqF9OCfDNAImiyOXcLzQiNS4ePuvGDNP6TpGYmC615eFZ
vz1yh8TsU1l90Q3DuZX+OouFp49hrhHVoaJnCa3dMvkgYzrtOOGVDn8W6X8HaA5t
IkFADm+J6cW+n2qE1MNO5v1nSaLYS5krPVqDhgv9KYR+gljaFytFCQsu/pyBOPs4
hDEz/zRLwShQ49FVMdLLo70jutAieii8sP33Yog6woQqETiZjwmpbzhPxwpz1cQ8
ozLXxYxi5km2Y1XxAn2eW3IORWKR9I9k6bL6Rmf9m1Qs8qFLQGokd0IzdwF5TdpW
6kqNbl/Y5Kq/WeLsXQY4ZdTN29q5V198C8PRQ71L2h8e4WpKnX3bnRoCEYoviV2d
79/vhIw7hiOPetz0t9ZnD71PkrjU4w1y9NlPa78oL1iSCbRuTKtxi97zWHxctw4S
fzhuqIVKHnZ0J6CQ4+px3DsCgEbytn7Iha9ZW3FUsLmLAv/fpQts6hokOu3u6qrd
q0mztg1gsreIpdnHMhAorV2YVafPA73CsnJJfZ9QXfZDC+GgfNK81xdMdIqv9O7N
EApR6Pq5E9cs3swUDdN8KmKpkHiTeX3RSLucH029PzDRMUTJBYGwhTp6xwWUdlzd
P1voypLsMkDidDg2jacQkrt93qBrztORFbG7Kcefh6V12GuDSQmfXIt9iWpED84T
J7YAP2p+I9lRXNvFIBxihb4/5B7iRatwC6w6OI1B/JWr+0LW6+wtMRbcD5QdGFHA
VLe5dXfeinypk1TaBRqTdrWAUWNp1+Y7D066jSUNt/jp+RNH9eYCLPoLuyhVLuCG
mMGPJl93ybIhZbpULssrAMpMXMlZivuNi8hj6jLQ9K2p1wsLNk/D4v9vsykPXIrO
ltpgTKhWxfv6h2eUMu2UimMttG/YCWZcTSDllhbAesb/ZnsM5bx+yJud0Ua3xYuG
t9jsI/24zG5T1gqIvHwHJ+Lqjr2GpdvRc0Zbw6BdtS/197/ibccDV1LuaQ6cHawp
ulmVmrvoPuI6+/XlLxXul7OzWXQ9hyvTS+EHpP2Lp6bUmyUCwzmU2TD894/wiLnn
rCZ5mHSoqTx6PvPy+4JgM6JSETiOukFonM4R1Atofj1d6mMsqs+WFMDR23Us6CMu
f5PfIrcvFhYUM/JdOSOfcHPxemf7mldvL0c7UzQu8h2xlIXRzaTGwTJ9L5VEO2S/
66C2hGgPxRCJ8pY2oeNHF4U1Mw5pTEK2EnUWLU2MShx2z/mktt9O5XmjjiCHV/Nl
+y9O4cMEOMpAiYfTa9Y0syTYVo2+gd4R0CTqXoggsRXgIAYiFBSH1EUyomol3rr3
uz/FEPG1KTCMAxahdMYsvoTqevH620HObdqKXA6jpQ5DrflIbhl3T5p+n/OkwBzf
KPA7tZlsnQ42JQBruy7AlpSjKPUmHIWbQxsaye49hMYfJTLrDeVDrj84NRrJiCYM
Fy8q2SpLbA4yaQ+vQh1yye7CnWmsHEyxKGNtBMWdnkW+ORWTUh6Dq9QzG6UhqQx3
XnIhee4f6B8g6b5rg/hmqnikMCASTtsslWQxHb+HoXN2Enczes1J0vLx2GsFTzXG
tMOaE3kXFb7UhUN17BGP9uREjkt6yDSUh36gza7bUkGTQYnR61ybfJnzCdtq1yFC
hWPLujm89KfY9Fut6nBGkHfoAKerx1UhuolO2+GBsCVwWjsN6o9/lvpTAvBFxdPP
6w5PHGmqv6+kNTwCHVhcWwOQshExYrxKFtGEHomm1WRUHtxo4D/fr7CQU8hpzYjd
DD6juXplZn5fYCwJjZ9SA551/2dWZD3N7+DRMZAje4HbtOogE6xU3xiSBhpt5YmU
c2QSVehlf9jzPPZ7RgXzROpMURsSPvnSc5oJrFjBSI5X7oweko48iqMKgrWGwHNK
F8A8r58wfuQxyuq88Y4FfjlHiWxGzt8F4reGnSBeIaI2SvIUiOc/j1Cxetg3z1JM
fNDbjk7WwlITI4pZh3eJE5Dvab8ijT5O+/8djLzvkSLbAg27tNK/E+T/WJY5NVX+
Xn+ZqaLWfqTwqXiksac05gNFrIzGpcrTLr8WuLh3QQpoe/b3ebJgIhCEf3rTheUe
8Ee5w6fpEjw+UDXwxP/EfPJy3h7YtitryXUYzXOrfeu7cdLpC/ol1Y9bLahEHgX2
6V86Zu5yuuzvV9GhXcVocoJjegdeYgKdl26+UOO9D3Wq29UDzFdyHV24a0thv7G0
hiLpntYtT4NZVgAcVgKn5oQH0MEPviv8hfx5KNds3kt4tKLhB+BoeBJatJXJgyXJ
RgIWUACqh1hACOQR17QkUDPedrdLdz8A3ZizueSuQHsq0wm66Ctn+lbVp+H5Gv/V
aaq25uSmUrZvFX3+lDL2Ky9hvrEzMI3ACERXWQVhpHIXvX5ox2RZxJez/nJ9TPg9
+qOYTgIpjvo21o+UF8VyT3wm38+LsBqzpn8ZvguEYKtmCI4fz5v9JzzvH6pn6aNN
UQ3avPBAmHJwK2FPW9UdkBE52weFg9khec4gUk8+PkybcGmuCNn7R30posmSGGFd
pvS41pAoWw4ZhC+InO/IfGIwmC+o3smevU1/GICae9FHzZQtjCAubDRIrJKqo/Tq
Gn1aQAzMMLYHuwpLflZRKQVCgaQL4El4drsE3BQJQCtKNqAnJVecrxsIzWsjxXYz
y3SL2UF9pm1Lji23EAgZnDpUIuX21hmlMzcwvMAgOPbk9BqI1tEYfiq1wuTF10l7
YpDgGFs0ipffBsLNreFjKB+TMweY1zNuIAAheiqVuY13p027w0TfiD8WodahS/oC
T3UYoy9nOLmgK5HA/nHgPNTGmza4bAH95OWStfp4GtP7edzNoLH+Z+45rtMnRNzZ
I1Z6IG184vqisL0zdx9e4TJEl02TbRQMLs0yFEoyCgtEQWqvTGFlwXTArPeehmt1
+F5fafbt1zSQaI4pM7bN/zh1cD1adxrl7vCmxux+sHWPR6UKJINrz674YBCqyOG8
ugxFHNLXpGFlxXfTI31fSekhukHzMtXsVVoBl2giXbpYFXhkQGILKsIRqiEM3qCR
AxanWU2tznMdTu2oS20CAHkj30mFCJmjZkmGpnQVfTS6GDLyOgUrXLS2OEaVvN5h
BxccAowdGaYv4bvc8WIZtVLuExWf9Y89bx+ChJab+4TRZaDTfiwcadh8HpXykB5z
1JeyXdbhkGTZLwfcaQE1NwkCYOZtaIOoga4yVm7eKK7a3tSs0xa+Ng6EQlQbBqCl
7U4GkQJ+ii7ogIDBtzn4F2dt9MNDc4HsggAgEQB21YqcQrmqRPYC/S57q6VO2avD
cZvQ/832JUWmvH/wJOH2tLxrjO/oWyWP/66VLa7X3KEhLCzZLHEcH9ufG3/tHsn2
o0F727i6/Ql5m2bQwJZMjhCb90DHCGTt7qoCKgRYciaLwoo1X01vLSPHDpvEKsLS
DxnFYclIwy3S2B328Bt5tPJuWmG2KE2o7yNt4I6327rKbp7KyNPZ8Xzug2Z1Kmna
1NcK85Zq6/sQsP0MrMIeLUGE8N9WmaN9uoZIEdL3VewvQpMcSUHQnl8u5Uxx4A8F
CYAdFDSoYx6nUxyCqwc5XMPgxrC+blIBW/I7bLJWB2KiHcREqw8BoZRvyFiFTOh/
zPpI77N8VXoZe1HeJ5RQ6awXtzT+5Zr6ZSv6/I1GtA0rxxm94UIHRGOMfFJMCrDj
UEQJZcOx8l2wihwMmfhrGxWSvRyx6j8482bIQeKh30u4IZVZc5ArXNyWoH7yUMIj
BlqkMkJogiiEGdkIqSlotW4MoeYWr+XPfWMTceICxMh3ILL/wmxjFz9femPlItUf
wGR7ZzHhlWwp3wFcF0PS+hif+PAuLtURAp71XpHphPdsLuWtfgjo64pfOtdXwvX2
g+bt6/22VDVsTX1ouNuXXESxv3DHH91C5SpbLut72WVgyPQHAGa1YHWwzy08WgHN
ng1rB3JAO5c36PbLPzAU5/78Co1v0QUkeSgbfmpQQVDhO1YcJJMpMAjR+eFYXUMD
2MFtofR++04E+QfjGjzCYVyArITHt5SRoEGj8Pu4CX/d0hH60Kx8z5CYw48ira4K
o7Z89MGBBQxUHu8MV/bfn6zSaEU8cmG/MbHQ8AN9HrGvcwB/tsjCqYrteOGZ+0y8
CrAWoMs4UDo4m6COk+yTsrnsI2aSx+I4GNfmz94Apk4Li0//N1Uk92DvyA+8b/Jg
gZ0DsyuC9l4b0HPmzdGGM9obPOYnhOEKGfgtQfsO3oUeKJXHWIk2dH/2a5l2vodd
HbSkwrw/nY2sM3XbWmhBgiw0eycGyj2YOy4ZYf1NyDNFz6gTFPpNJEVMQrJxV7uo
+64pz+hnVtqhQKSDcH2JKnKTF2tpFxpOA3JZB6mdnDaS342CnqBFLmCTd2whAkp3
caQnUdxQPKE4KB77nH5aSHriy8Cy33K5Vo9XBuY+Wg5yyKz5m4drktxLrpRmnHDK
3QLx6Mj2z4vIhCOyqy4mrcPl4WqwMzW7An9bDUxLooIzr5T2sHURgur8K2ChOmcv
nuUUQuwMfsgmY9s5vK2z39yjctc9DDYiWOiU2jXPBpIny9i2o3DiryFSLNJt0Dze
4o14CZTQf/UgUwvZuG1BWeqNqb9P08yCZla6abM8IClfGsp4Lm5W3hMT8nfsIo6h
Nc7/IivdZcKdvM7isqu6qogMssc6+YwcHcX5Uh66qMuTgvvFH8rFvVLLtxB8lbEH
NxUC2+et6hLJV0o7MfkCvQe0RRkutN0Dp530VMERUTbf+fnZ5zHqQyCljJ6r/7JD
d/8uo0NPWFgev9Uq4T6Lkd8zj3ToHc3wziIfIlnJXvf9Vu0YfjAMizZo3165cQnm
uXBJb/6A9vvwZGNbUemFyxu16gqTkDEKK/pIjwCa7iFl58OV1G4dySDtFjQr8Lg/
VJMOq2hJzW7Xkf7vwLet0i5jEhB9mnU4ADXI0XzfkLjhlthw72QP2sDyNr9LB2Jk
VeV8tBk/i4/LM2WS1VR33wMm6oNRTx6VPzG6ernjoRmX3F4LuQ0Faxt33n5vMoq2
zQbprltr8jZg2PEJE/Xbe0kSzl51ekjJ3yAL3EADVXTMMvN79l2uLpVylhhgywmF
O6K2Hy3DYEfdBQbVuZS9YMRi9ZbFHm6MbBiDcalMdLx5vqbUS3zgeEatuBh3jd9W
eOnXsJA4cGBu1roV4NXwtiN/Krka0bqSbAnxlzRFyoR84VwuWgV7PBrWal79/nl8
p2wktZQR4sC1Y01zxv3dccZUH5ufCeqWGEzy0zz7/fb48HIvEhSxEgupaVvBvocN
QqI6wr96qymtyJcc6HgWndgatRZDCjozo6p0sXuqKlHUjDcesmeM8AdK9ZLvpoM1
HOtJVB3nPCShcvj3XB83/7oAnF1z0lDK5wUZHyBPAf7GkVD3ITDrQku5VYjDyR/0
1Dq5RkZMwkx0ZjtfYNG6fUeXVGLSvp4sAjloGGL5QwKJL/KPi2ZuXKlNbIbsPvRS
29SuRXpIHT3PChTqDQtdSWiId1QEcuECfTb1JN4NM8gdVveXKMfef9q+jFFEJB5C
gNGJQZKrVvakwuEdhNSO3cMm1qc4RNWpnSjfG+qE8YwRo6a7PUUrzsabEujaSM6E
mhQJIzK1mPGvpcXfYvYckGOkBycnHGe3Yohg0gHq4dUyqzu0ghLvV4+R/EDx6Axe
kTSFsZINOreyFGYxFkqpJXF3YzNj14V34ZO0OmK8SegFWguB0Oy4RNytDd4EID5Y
hfghKB/eLgU0Yq0ufAnc3XZ9C6B9TABDCQVBRNpxufPtuOxlzEx+DNeN14HUrBAx
qW8PcZ49cV7vjLPtC0rI7j1G1woFYBZwnpNiqlavMRYi/7MtyRhFcu8cAGaK1Mcl
Vt/ND9YLvF2kHU7lA4GcRlm0wUEXmXWHjJByKmSJVBxWbphF2wg6y1K0JQZTqi8W
2foM2pJrJedD9I6nkMSgMoE9Dj1aMs4+I4z9j4pzcAHre5/Z4/dm5LY3ItBXRYn9
EFNTacB1cAeVj/YFv0auP23pYYNB71AvECllx0XCEEqiKZ39uzkvxumsV4y+Yb3C
kEGAveZtEVcpwzX7d30gQCf9Z/etByTQtp8kQcasyrW5wmNTZolXnD+IYiBaqurC
+h7YPZHqi9MWINvKuA8I1IyoT+vhxYyLo4ovyBhASpNmArSoZBECnA46OERaH3BD
MD6Jb18bUfB7cbaXz2XK/7FWUa9Rb3kN5OsbZ0tv6LgH4Ik91K8xiQWp5C2MzKTS
p8VfMV/eEPoyt70D5WlitaXqd944kBQ/yp2TsZaL6iGA200iR03iqpgbcz+Zr9SC
iNElV33RlcJECUX/PKlxX5jaAIT8Mt1NmiB/TEb1WI3vMgC+hkfFVK5DvEb9uQ3b
Mr53VLVaH62BtuE0HIaIYdQJ2U9/aZktOR7dwVpRa9w4AIB06LL7RhB0nMwQ9I7R
tXwA9nyLUYQP7JGJj5pBCSh1V6Xew2t+S2I6pv9snWu/jRTg63pkhsEtJwZPDIoq
Hh7fR8I7KC0+tP/myN7LU0/h68OgnaBhG+zJEbjtadrUfetQ86cRyij6vw/QIZAV
88b1LKibecbEmCLE7srmA5UdHv4Hy9X+elMVTP2OLsoTDB9T/4FLf6yDZmWwEOLJ
x1fSTBXyQnqxHIRY/KDiSSTXSVyyNtvBPo9tzZ8e8kI9oRxNLPIaNWR6J1yIUHRK
dDEV5D6t9gdDsKCGLQrjHuFVufFR6osN891Pd4aFhlTaokAFJQ2SP2KEWD4sTck1
sEvuLRBuJ7L8UyMNTe+4UQmiKjFPXG0oC8AYjXjTYkTxE3JhjY4gp1tVy362ueLT
5B7lYxb1UiAZ3hIUmpbCuKmoo32Qsa6ojD/9lvrzp2ZGX92n1/fTw83+/6Cy8lHX
3Az7LdU/Oi+21W4thyIYq9n+mPaZCWxNuxuy0MRMl25iJiQZmFMTz0+BT0raXfm3
q9/jmHawWXEWgVm+KUr5yhp2Yb6zrtOa4ql9/m9gq/YC+HxrlC6fR9D74CHAAUK0
sPccDx7hlbv2h3nyjVRzHFAiUzsHfMxowMXJAiwVcIBZgrcbyzYWakaEk9UxXRP6
gZtJqkdQDfx2Zp3k5HkRW0QkaG0hRJMtZ6rQrvBhG4SFoUHw7QmTnh4hyzoa4B0Q
adm5xSbBeEB7VEm4k+jxUhOa4R2MHDyH9va2yTUuvFyERKItG36u1i0KDAhiwKcP
w8a6dLWPtNWAh2rSnS8PMire/gRlE3+9iEYsHqFcsAQfFyy2JUnu0Bslbyuxdb1a
G0Y1kEwkD45CKQxaQGDleP3fVI483zDhdqtiBR3U7G2WXM02Cm9K9hUSQwk5znm1
5UkOgsOR1c4IPph7VOwK7tqLTeBWCSYQg2LR6CL2yesMusmV/mlSyv64l9/Sqenk
7+8w/R6Fc1ZAY4PWm9Dpqv15r+/1v28abVeTCVTPJggQSNEvDfl/NjKaHwL43zev
dHhWiuvYVQBkPHVpVBs8fGCDQWntWY1oBn2yeyGfWnp1yr0pi6bF0u5XwkXew0ml
31mZdToPT+9/rY1xC2e2nWAc8rsW3r9mvafDDTbeMKhc+c0nPAqxmabOcDK93rzZ
8qaT3vfE4Zf/Vw8bvQpf7OOwydw7GfDc1c6Cu+yvJjGlLOOnHDR2MXvRJtpsIcQt
w5wcM723+K3HSxQE94Dl8McL0OUqlq11mMEgvzR+FprhEMLXbbuCs+7cba7zMEtR
MZg7ks11WvEMrJIPAjqMkkN/YGXWYsAJhqvNCm1IeJ5FxAb8u3kH1xWcNTQyGtvh
gz2/RJwsBc9+TX807VvIGEaWcv2LZMKkTHphtlOfMkMFUsPPXXhvibqPcBm0wayR
RGrUWUjDtLest/WURf4M6us3VukIzcC3/hhDHqbJ7cfU8hNNPfsTG5GnsqEPUkV9
JK163kWn9AygwhmlxgBHjYg5Wf424cXkS+mkR54Z7TvafHWp1PvTUPqI23sf+OT4
s2SnK194gKlEcB0DTQmd9bge3Ra1C+C7lo/9pPl0J07fOGmGc5FNu0x1pHr97Tr5
RXPL17K6xaR+YjzWmnF9fBxLenKY8GBqE1209QSY/Rhb7UrrdpObPKOPn2jfA1Rm
X1jjjIsU+E6GFvN1q25uw7QysbRpcbUz006K6qddM0YhkKnHiRgtmhlz2li8zl4c
dANfvwf3PovS7Fd7T2uswpZRFAWnHffWw5uP+W8I7KYgl1soyxSP+vvWmmZMrILM
hV3Dk1GS5dkz1UVSra74b5nbPRc7BuU2hijzAoWdrww3Bfnz5anBRYx+sv+H8dX9
ZBMkkQK0rRr0rj1HA3ky19Re1ZuOsW40ON+gmDnV7+G+fXD344Xmup3MkkR5T9Ww
1cOmv6GREDVH/mAJXiMsO5W3mDjnCIXmaPFZOlaky34IDU42f6Mv9QT64JgKR39u
qeCP5DTBzIZzsDHZlmqCW1aDNEXpGokHlnwWzwZqMSnMOqiCvVbAJknliWMtHmRG
n1+mHWjxKyGenl1Tc0m7fZGyo37GkspVwZxNSzawI92gDRHGQPfMqyLCAm9BIHS+
0Kb+sBU/aJkLQBCAieJUA5bjI8ZEGrxqHnX6ifDpd+x2CfM658dGALVSF/5/IX5B
V51Rc95a0PvwKLE7iWPRuV0LgdyJls3lxKLgkbJza8Dnb7AwkT/JMT++UtvIlS6Z
DLIdJxBLuTdJ1ms+QX5cwdp8kJiKYYEOwYZiMxU6oxXzME3/94d3uo08qHpHuxkq
rW65bxDJYzr8jRNwYN1UGB1OjTUTebH3iRRlzrCjOcVBkE4OHYcIjUm9QWsgaKAn
yFDLe0cbvZRPj067QUadH/BOlgLNbiLtwiEoPOzoqTPUSBXXY15zwKmJRRPlzJsr
QI8Jj//m3kuKiBSreffApbBUBIMtvAfQlGQfCAHqcQPL+CAvo1Wo5+Nqs/raMXZ7
ICZRmp9zh5wM85LKAvOGSci8Lh80begDLUYB2ZpohDxhApA4kPyT4+PmYSz3roZo
zqo/aKTUmf1YUbMSaK44CpCWVJV7VKdEK4tNxRSfvPDdZgf9rZstqkLqszU+b72K
BBzJd+71qBe8lsALsaa+nHoFIgsukrSR2AmFhwu/zmnc7yFm0Cr9hCsnsQV6w4q5
CrNm9sffWU386rDyTyW9XLrtTRXm0bDHS/OmzfPPCVRyst6FPF/Z1Ienm9JkqNNn
mzyAXtnyFMk7oi8QuH1uKhpQh7ZNVoIiANlEq1zZGQZ4TLtRZ8KIT8yjLE4ZC09l
Wxb6GWNUj6CzJ6V4b/TxNjx7IA3bW2NigvFCBnNVq6YOgxw3IS6s3g0KwwRiqBq/
tqP9ZdE53fmkZy0PP1Py2yDf87horI0yURQvup8QxXUs71du1+PplCRt9aTAr9Rz
rrxepkgTt8FwRFGIYz6IKwqfBCem0TrNgvbP0cicBI3ECherolTmUsISrL4h+yrq
26PBNOEWUpgHH0iN+uQ4ecEVlBjcjZ1/v/o+kfDlU2BBNtCpzLD6opHunulAIMV9
EodpduW/clkgabeYi2ew9oKKbcCEj9as65P7pH4Q4CtD2k55MPNYYJ2oHTwevMRT
DlC20r7Ug9PAHtzc8lhF9QNvlIYL6RPnFlh/dQJegwYGzFhN+6WfkcPToKq87jQ7
DZtgfovkX5+pczFU8j9EtfeiuhdgFXczwPFp2AMmGi+fwrerI4tugIL3MQ/EkyGN
tVGb7N8ct5Sle6HfHJEBCmJ1jFMVZx23GFQRMPrqirBbvdi4Qwi7eL0k/X5IY876
neUPTOh3NuMJ+C+bzbpA9i76yWP/933cI1AJh2SYGB72MpHVnUyMZ9XG9LsseA2F
nq73uB66E26Kppt/KOZk488MGXYIOfc+besSSkqhHbjavwAurACCSHSH10Q7Y+KR
6ID6eUSJjY9P/DD9u7PjHzRHIGmnUpRqC8PkvUlA/OzoNfv/y51SEXeohLxfk0xr
t1dWhSzf9x0POdtte8V4y0DaONNMsg8x8AbnJZl3ffT2SPO71l2Bs2BnR69tGox5
gqo+vhyYS8U0Cwq2ufwnxmnxDBroMRhAYzljxUF4ULZT3f9K8I6f9RV7wEjy22fQ
sAliOm25wXx7KhPaYZGI70uJyYrWL3pGYYZ21qRidx08+3wODSuuZJCqXl4W+1U3
w3h/Ya9TkgbXcac48R1l1x7kYr3hef4ephKiZop63IrQI2jwG0QpDxSz9pwHcjVD
uu0Ej6sMd0s+uVZXtmxFVxGhZTPOSr0AioJU0x3F94r98UMmPz59raohzEe6wzXi
F4sYfBKgzvq6U6MmNBUVs1wLBlK//vhPSWzFz6nKHKPtiPaxTNr2xJl3u9lfpe3j
TK5wxgcVn3x+2VWSnkA2fbFVc6VabsVfrIjrzsKjZs4oakkd56xc9F21ByhfVV2M
fIT5ArT3MJnAzK1DpSISPpXVbs0higKjzFt4xp+gtg0CHgflb9ef3+56qH9GuloS
qjJ0mFOm4xUZ3TeL1iJvNxT+Wky9Wc1qx+TWPfj4SIK239t9sIGXv+gacsQt7/OL
BhY5rvqkV95WaUeE2BgOWSSEqgidnlA95tYx52v6NWOvkg8fA/O3qEX27ULNo4Ch
saGYrsehN7QjZE3cIKPRpEB9puwZcd3STEyvZBa/CZIMq55M0R0H6jYD0aAu6+JA
VZd1py608oadoOthvDNh7j0SWfqZVg4MBRQwrdrbK+OW1P65IwOH5W8WNWKCYBdF
r3IG8JEC5JotS8qPZDsry+oUh9Nggnv7DADUMSKn3K8H0i/oAj8yAAcCGANnoJP3
Z3WdP2nditSJ0AdIyTVkJcjXzkoOhEnONaAxPKp8nIA0FL5U++FnKxv1bpesMSGd
+i5vAlaDBW8I+TcUp8vwnk90Br5LxPnrCgbBY3+B+6gxqHpnGL2X6VVdT96qc4mk
0RYuGZVZCreJZUV7Fzr3QHfB1fyDIBLSgS03M5cDGmCdWebPN1sHIcC+nb/XlXWY
ePeT1DKK4SKz5DLwhTjyETa9hCfkeu5NVe0nuQ2QqmQXMmbGJi1n25zFazmGiwHb
op27gRyackO0REWEda1crEch4ZIFgDdjVucrp8ZOsbvR5uqIY1ViC1eA4evRzvcb
sOnBRV9TyCkCK8JwdIDVkihW2R/XCXcXO9+kZEbxYPgv+5NV8hhMo6ozsplwxdgG
fsd8OR/UsWHndNgoiTDcxQa4hWUPztN1LkGTt8m04wyZvaP2q0gJKwkMoOFs4WXa
i2SIyDEsUHl+xOkX9aekzawyh6w23sjzt81LWCQQ4SYLH0bCYG1f9MEjhU5rl+m1
wrJRhES8kKNynHtQMlEFlBbglf4T833V7BB3hrTGC++FGoQgeFyDH0bkQS3ZHQHp
XGt+msrS0RM2QNZuxFBU1QKFGao3uKLg57S1o3JQv+HQYAKH3v2apXJVFOJbNf+H
9Eoy7DMXYq1rn7zM8TaeylmdNqAzKmkV9oq8dH99Mrpjvfmc840H7p+n/HPYRoHK
cdrUdBEcE3XLBzdJwFfgpzs466AktjZ68u+dHIYx8nhU+z1CZlUGGiQMvGwi3vV+
ikaUt+LHdm0XYlB1FCbstB275PYTy55XPEW9JfJPl+YMwYwUVSh7QnCiurEk3fW/
x61FAcSFi10+KCQyvpTZKmaW6A5UfSEqVlfh7RXSyUczdYht4W/YwLOpFZzIZleq
cOiZLpJhprdF4QrC5QNmKQ9VWPnQx/rVhfAbfvI2Lun+0whezZSXdG8/+3U4H283
p27TK/C3+8xgKe8XXLrbKdYnJJPTym2YTyTR3KAsZC3arpwisAueQ9OA0twY7HGG
vmySPNXzzakBxAqDwEOVhBMWdeNASy2VYvV8aUkm2kCQhfQwx3OWnFx5lHZOFi3L
zspLWRKolg9+ZrIFU0sfTQ3vqKxABgm2Ooru8aLO5zJc1w1ogozA83WCkKEsZ74h
9riAqJkHXJShYciq03Jg3b4XXBehsf7rohdZcI2Od87SzPmsPWxCbCkL8Qqk1MCk
WYlWgXpnXhqxKimcvlAMAZxInf3kcdbpcEqzvmReHj0c2iB+vN04LGbuMMoBxP32
07CZYPgv4zo955eV5XI0pkW4QjC4nEu3Y2L2xtHi/8jCPUwExPpeDUGxxNJAfaaY
jTUny34JKwzTuIm9vrPQk8ysp4a1vSSwEWNmdMD6tGZko3X0ZbZ5f7vI3MMMOckw
C4rPKFWaCkYnYzQVzoqtGfYk0TrYPq3rvcg9A6CIbJf+vKUZ/VMzVzEOT7CG/nOo
8RPbVgpDFX+Ox2TtQ+DOl2YL+m6o3lxqkmkiweEQyPu/+yIirofQOzzbso30W9g2
YoZjXt/c3/ahCJgUjJbSYd/Xz8RReer5WKePM3yD11TsLFJGZ98FTgsOJ+ShZMd8
yoXviA5VIiIyTFFy7ItNp6YYlWTw4YEh8Spndsyl2Y+2IKcmXGTrmy37Ob8cCXkq
v46+B835X5zdhkATh29bFkhQZx6JpRXWLQnSDtia4xIXsOzsB/Kiuu/FoA8RPQ7b
1Js/H0bxjVVFHCk1s6hpH62o4WUqGInJoJQMBWlDlw7o/Rf1b1wLu2ium+TnXZnj
kL1gzKSWf+cNeglmHo2VnYWjvEBTsOMDbITdqJqhqXZ37dS5/KuQ7r2olUSrBUQr
KUQoNpApx1FqlvrnpwsLWJTkbCnDruSIS9vLjhcW5s27UKavXMe/F7oqbg2Qv/7Y
MruziqOK92/fgY/dKR3TvvogB1NCwTsl5CaagnB74H9qytp5wPkJKKnx42QCTvgM
MI+2d6aMpPaKinTndlGIIPh1BtrRk6mgHwEsUs5A2Aat8yAU5KCRj/oNfhZwvrrI
6pgK8h/lLz5OkvINdbtfkTLk+FcEOvY3gOQxdO7L22lYXht13GqsBNiK4m+9Wy2w
2dJOg8DYPdrZKLBapaI56TYrNqKsQQD0XzzYq49kZmx7dtEkt++QutVd98WfvZW6
QZqt8rvGnfItQ5Z8f9nv9PEcseR1Z64u353/GqVds1oMs8nZrcwXn20x5XHlH59J
KS5ZgGg6x3YHZwThcEWdPS1Zs0zKtwB7xlYdpO7LH0rkLJiUxPqIY6HhhqR31gYB
YTnD1JzvTELfVR55QnxcQrXflh6sxGb405M8E2YmUjn6Kh10wU7qth3Wwiz49CJA
1kQXSNVd/0F0r/vC5s/2GRkzQ/3maZJtlgkMl5GEs2tfMUcXWUSqMQIDbM/9iBYB
aOPAxXE4DIghW+4qVFDBkz2dvbN8vrZiKFA+sxj2SsfoAmRVBgfP5RoPc3j9ywCE
8C+gPYy9ld3L+zx+XNsaySZh1TxRbdkO8/K9yG8CfvkWUgrZCrUwhf9FgOTfe6Rn
woQW0RrKJPm8NfcqY9S8P8OewOasauuIXwgbhPkeiXGxKCQEWpy+EgROkm9QmNNf
7OBsr8rPVU7VU2FNwti/oN6Hz47sAjriO90+D3U+Cw0SjQzZS5RmBKZ8iycK+LY8
ERUi24oM5hA68HTNg6Nak14lyzLHcIT35TA1gGcQmSIhyqCobYOapX+3pRTx8TfE
ZLSO71t75Wlo7oWF940zyfPyyf37N1IJaXXH7GZ94EJKX1BfGzbSlXc4yrPnMEVm
gJA+GAriVGaWODstg/pgZ2MZ8ueMkJZsdw4b9DAWZz0BesMaNfpoitPorQHZErIz
lK6rmR7z3m1acIAvKFbQj5Dc2ABwXsDroSgCoMhoqAiSPoCrP4alysFX+6SDxJRW
B1Fdxv8q3cVrWOGgS4HYz3QWQ6DBZI9YG/H16xupYJGSq0IWNI0L50zjpGF1h1Tq
zL+kx91T55N5SSPs+g30iunxLMNVIRJhoPxtDa+T3D/bZr0OST/XGdiRscr7RFk5
zHdOdg28GO2vZ4jBI+gKBiMX6cMN85cOoMAQueOjMvQIcfaMr0u3ZKUStt/lIjKA
lrPm/yrVJ81VsELb0kvELikFdzLsFUJL0amMnoea4mGQsumgfpZUUenAW8TG6wP4
OQjFCeLTMwH2GnBQYJFu85RrKkC/JSy8ZogF7Wo6pHc6PIyZRZxtIBCtyX8dJhS4
kBXQtrrQH2br1dxTwzqi3oRM/5DXaxs2dGhQnXw9uzKwVTEGxNdk08+4GbQmkuj+
r2eNgHRee66tcn8FKgMc7a5iRnea4Ls6/6PSpwDACogUolDBGlPZkJIdaxA2IRG7
+zthu7SAZxoc6sQMKJXouM30iVr2/7AILneSIXMdBsuTuC7qF9PLXBDn5qvDCm/q
fYntMpkf6atbKlqe4zZhUJLqjyfU+8bZMnqOyMOq4wCpAMT+Im4BRpmnZowXaW72
L/PyEjhsEnXO2G9JPv22/RS6Ue2CWcsK5OGJpng7SMEh1EN0w2tNbQv1oQqyK1Kt
dOIsBPC2UKHii/WAF0j1SC8UaXeL43M3cUPCHo+e7PqEBsen24PXF3+oJl8tIJXy
4S39bGsOmnzknWqzpK1zdR4AWOhDfdJFD+Ua8T1vLDPmH7Pnu6LXlgP/TewKtPqn
RZH9oGfUks64Lc5JB2Phf26CmzoDLsCZvc6qnU4judCFwgZSfskSzSIWzJno1XXO
G0Q8BPVxOPnSbaFr2DrAj1b0d1UIC67udlKO8BKcm61ZFkHkHAs+XYbaAmWsaUq2
kdNUdEMNoBq+52c2ovZRAsPwd/ghB/5PHJJOAC7SGJBq8JJEUBOsUQcnDmHyCWaQ
+XNHOsDpOL4Z6wAxOHGBuvoAwX6psE52qj/FwBjXZ40+/4INlCG4T40uzUiQRGsJ
Y8KVGFqodVanDl2eLJMs1teOqIbbJn1roi7o4HE5WB+lWMgbW3B3NR8JowFNy4iT
C4tSqQV7dPbxP8/fY9eppB+ANxBjTfxhk+A96WsHsFavvmmuUQZ24dRSXn+beoXd
gmdL5UFANmiCKyIuEhTUe+jRUpzFgwcN9b7B/1bviWxhQFAFrnjtc9fnSvF3gWai
Nciq257fhseyDSbbAa10nN1lH03SzFH7oQgaXmOW2cu6xjHCD9bpRAA+krmP3MSh
3zz6zymdeSZA1tipbsyDSB/HrZHm/sPzdgjhAxyA48CW3l3lzmLPxPKfUWe+LTZz
KOstIsskxFy9QKiHzZJ/LTqTSn2MDyxWww7m2k6CQW8+g+qJxeo7tJ5m9+b+BWRy
wm5KMa1K0xIWvqRrhwSfd3rwA747JQR+CCWsDpvWtZ375zKlPKUkapPr2zklj0Xu
iW91/LMQBxnXIa3EffobF4ZvhrgUt8KZvpA3QztjOEJLPJJP5wO+fZKgcOKMDJZ9
Ta6NX2nemLmLQ2JeeU5NeLpfXpqHA6yw9JW2WD45m+/u7aDe56iLM64lx+p9vbr+
yBySPg9NlvRhZ+TIhHzOfs3PWjJiKCLMjsJb0HInUUVF073iUbLhpb3X47YgbZ+c
N4pkfmqAvp2rLRFJGnPwJXU3FpX0NAJ009kYNX+aMXbSdopj9E6688x1ytj1FF+4
P3YeQAX8eeiIggPnAnchhxvDx+ldCTY/331deYouw6f9v02qwEtQm7NmU0F/qkEe
lNQegKDdWnh6hx586cTNuNUoxfZOl6BYyYgzaQre148yzkvxuxNiXGCgAtow+eUL
HpWIZQjjHaGQFSEhhlZotua2h26myn+yTsZBdBNFnbfQRYzFXIiCbAxctQqbsCIx
ZkQuy/zoApNJRRIR09CIYzuo2Lzd6ykCW5O1sTen4tpa53BCwikKWxAvL+bIoY1i
R5V+2xoIc5/6gR0gCbh4bHLYA4W4acTIXWY9TUjlbhmEMhc4m4c/gjOJQIIvwwv8
2SrvgN/xn+rP7FXKTTVQajdEKbxIcyDQx1kKuUqV7S0nbtXjubHWPrsyEg/05B9r
A5bvh5Wr1m/eoh3e0pzvdwH0QQym4Ar8F3kna+J3iS3grIaETs75rAnGL1GhEcg8
TgfV8BaLoDV7GlIgsCj1bZMI4OMG9Il3NsXRePoQgor0gKxozi8OfCagok3qPW/Z
ChjHM5648cBOjXV+e+hYymTz6yrkguQjTxbvuSK+ZaU8+epr94f1OOTDIZaOLkrX
xsRwytnR+HoDxg27V0YIcoe4rya/x6j5GSc7jq5TZc4YKpAn4y5VWiKrhT9X9sjJ
Ish0dTmG0X+1jVfVoLQ2UtG/IlfBcbFlP489jY/AM6CUd4Ne4eiK4Jeqhuw79slx
7IGkmHyPC+SAGITBh0GmF9cv6/7GEbqtasvZD+ThFxAcUGEcKmRxqzVi+4t2nhbI
VDFLi8Foz3AiRtoomm0jBAEMnHsLL2tigsUSE8hYtPgr+iJ0OiTLRx2VvBl3xmo+
GjI5efisdrpxAFqYJW3lZ5VYOo7RBY+lxnhqoI5M81M+OXn60UbtZ8CtCC0Nn1Sc
x2sPjzYZSmXXQaMkekjgz0OJgt9VAUOV3SkITtpANNvjSkubbAVYfK2qwNz076AB
9z3H0GtaS1NhuBDn+QxdDLK04pq/GebLkRyvqLgzfh0bduiRQsPc8dzxWGM2lpvP
+9Qy6dTswKmtZlK9rp1v22DtVsjMfWv0+C2R40TLl8sMCpbAshxqE0HeeLvMy0G2
OunbgNf+HcDTICVUMyuDk8oHei3Noka5+I2zUXKcgNWnXq9s21REJlYvffv6XQfV
ka3ucJjOYUMl6wfeuoc7UDyDlhUa8n6QTY2z1SiR0Yzs5TB7MMqN6We1IlzfUR3p
Tq2tbtUzQG8Q7GZw7oCcqGQfB1lpJcXe1Ea3FTzkxc4ZqFduzil+BlT36Og92eng
J3+dBDy/KYtIrFwYLWHC8VXN+vGeGOJDYok8V5WY+XzdZPkkyrecOxrHhUZFEk02
upO/KDLLbiBt86E/5xMvY+7NCDI7cDPRSE/qdtv2uAruvuRtomgJXSyEeCuzx88J
y59ByMy5x8n9pgmQDHZNkT1y2ul/co9iPAp2ade3BUUaFFN86+N2nsWFMy+baD4s
08gWlNMp6e8HK+jHD2w5adWL9Lrx2CqC4EnkwKnF6k7JrcmwTWBXkPEAcynEYerv
LRTExTnEBohf1GMQ9b11SJah8DUoYp9gEancVppZsJ268xbOzSkpdCvZrf7xwwhy
1V+Gb0vdfwE3O6uDWkTE98UvrlnO9mytnQze/tfK+dd76cQZWHkPprqXiGPTTDV/
zATvlHF2W+gAm5fGmYPBhbbNrEmqUTHUQLEOIPq8RH8D+SpGxRiepx9SKFxBTx8Q
DcmQk9xS+hgPri0Sbei3iP+Z6xblF66+uVGTv17OO27CfCf28BX2foMdL5QhOCcX
OCefbkaVkf9bT8e8RqaQtsaTz9ek2gvHg9/pcJnsPlMAmut1UqRc7wlMH9Wfp42I
biLy+2UK3E12RMuvSt/p5mjR2K38V4oNUzomtPaOyvh0oVAnliYWpMrA8um7Bp+9
xI0O8cZAqhEA5brjEL3pDkbRqjl5X7q4oLAbvwDasrdQztGNAZ1oJ+anu2UHym9z
1LckQw9aLRHoKtv5ni7A57/BVmyp6CL8rKaIpIkXjQaGrsn/gIeuyc68GjBqdZ3m
JhE5rfUR4y6AN+ti4y2+6q1qSEw1BANNmy8N/ib586zNcJzkRVI/jJsD3/Ojq0ra
8+foMNcVpcxWNwc2qqZkg9/LZ5oCh7Hfj1ADMY07xkVAixUd/2Rm+OljI75LKYKj
wokHVdVOGCNPubFsqojgOp0aoe1n9U3+h/zT6k8UIW0NZqd1anpkgA09kiHbAX56
5PMxYdsXbwJM7NAHkKIb43rhxux+vsWJ0kqEEc86899oeKl2pZV0yh2QyPwj7twL
hbxuNbeGLgTaLbH4xKOth/lLHVT3Fsqgnyy+ieMaODLRv9pu1ukMkzkpqOH9CSm0
oPJz8zJDMR5t2m18MlkGZERYZzu4X1nn0QrjzYOPK9W/EpGLka0fHufvqSmsbPfS
7GE1TxYKzoryFmpQ2A6d1eogdyli/0nOwRXQ2YJlP8Avetj/jhAQGgbWZ+AYHwWm
r/9gA3jBJ8sTAYjlHF25P62kTB5SBts16pJLhmh8wuUnWeDl+yHUf+wA4d6kqEM7
tsuCmQul+AQH1wSP7bT5NYui0vTzZLSEoTQqysQDKE8dJOfS5AHLB1YAQ4p/+cdd
j51v44zCttDBZywbXDyb+RGYPOeKF9JheIc06iY3tv/eWR6Roaz2rTAt1IL7i4zF
UKytJHmZ1tiHh8tG8BaL7YfTjwjbVj6w6xTJXhmQMHQKRnlknTNSenOvgO30wsJm
IRpqefqrrgtNIPxqPmBtooIQnGLhSBVpfhNrZhm6YH1qsM1aDzP5PYThIyqH0IHl
rbO+RJNbS/m22KFeA0uMqBtE/Q8LRMrKKtm6qjTVhnBjGNo+SkLZd9tRNqwSWKWA
5zSLjpQwjnh3SHWDIEQcB08gkweWo5qpy4i4v77kv+4l0PIt4tIxzSj/STjGemAi
dSLm9SPi6xjaE+K40QZfruxMnAdM7+10hUavQS5ZpRGM5qkORt+WFPvAW6o5V333
YPYe+MCZEWcnuJ5lH32awiyMvujV3pMNDLUIvAFPCX7zviMal9387IoMsMcwm933
udAnThVxJByKzwOmOMQ/xDGHsiYNeM2HHGr5tD4hsV/Z0jYpqOFxNxKFGvraK61c
55elMViuoDzFqVIBv7oSLrFeOO12h+5LxB0qpXrN7E1HGCBVAsL+nXQF1Tzys+Mq
XooIQQ5K7CsZgU5c9VSHI/xE6nM3vnm+XMRX9U1H8a4NGoy2MyGJXhECoAMDaPLf
9IzSTRxZhPmYCyIZ7x1WyWuGEFBfS712eWDl6s5vW+4vW+jCWd0rEl3nXaoHPRVG
I2UWQYFwLUel59nVpBMBLh8GH05HWoPa31WFVGml8/nFMYjSIEijc81pZBiFitu2
6MjW142Q7DvAp2PcjclDYrTNPyHpDMtlq4dQul29+23MatCB2bePNO0idL56tOjh
lv/+SPPVZukvVXeiek9iZrFUh6M3bAp/xQ6uExa41vlYm2gQOVnEjEk+vBRUTl7t
VLTsIj1mdC9IAa6Un+XSOcQvQLNP37eJNGDGnUBxGu5IN3Hzl5ao7u+b1FT0RrXx
GhzSy9rCS70rvx1FK318D/x2IhmmjtCS9g52evxP3Dnv8M9zpj4XNEJVzkowZqEb
gzIYBdDHzFZ/4ArOCntUiMJHcivYVs76qIs8A3Vm+dONNw8zK3FQ3oQ/GNLW1RhS
2AiuvXcdrJS9uFxRu/cCGkvpjCNnzcEl2jmjrxY+24Z6JMT3HUOLSYEeiA7zpmsb
7JgvDOOWHhlQGKyPqZ6c4kmUXypDLniX3mlVJwMSC36Sn1KDMgfi4LQtGz0ZP2M6
dRSLxc86HwjWXzMfKaCBD0Bgr3NryqXD6cyY9gpObUmVoo7GfUIDapEakVnl3GGy
1zxMKy6NSoSqeCobGSvdrYBIlHFy7HCm1c9ZtMaxvCBh8A32Z3tM53HyrjaXAn1Y
wB+9yjpMXJnd30eb1jkMR4ledFKtl/6S2AhXPKonhRAd836UBKsE8kOY8yVxB7n2
SEfyZaWYCTeiD/QvN6iK1OoBVejdP/cQyC6FC7XvGCCEwKuFbNKNPLS0hi6IL0MH
WVy9nfVGsfkz48ZzVrke8hY5tIeaCWw/ZwbWgvxsMdwEnh3qeoMjDFHTqvMoBktD
ewGqT4Rx+gro+uhxSCHFGK1rX8YLlkSupmFaldKa0FIvvQb4FFp4ZQL890rob7uB
MUrbH3X7C12jn4fQ9FTHYK+kJRNQfbKFu3jEYnkHlMJIRIcbUtG7hUl374T4SDnB
XAD+FTYWmzjchEo+Fw098fj0NESSckpidSqzKUxYlrxuBPxMPNKUAQ7/6Nt8FI5D
4B5N44T0ul7EeNjtxwx0db4B5q4kAaFpepN9r4ZrXTEjM5OdEZkTIjSrtxnlhknu
F5EMwNJuj7TxjtlN2stQ0uBzh95UXnL6pQY5MKY7sdB/Cn4JyQRf5VoLHv5w3I4S
/aIZWnNwL4S/33UYS/WvhMYzA4ZNxCz/CWSUZNG+Pc5TZS3gRPDf7z3UHwFFHLFK
1/V+QfQtR6UVFnD42GMWpcWTPPxvXDW5YsunDu9e6cVammS60tvcpgXqZx8O6whg
MyA4qx/+eVdPBkajuHWGqw/Ii1cDs/vvJ0Wv372VabYG0rPl9yoXPBACrGc3wG4i
AeD3kMXf0jwYadmvIrqJTZq8V5J4bB5wbLFdaw8xhfXj+qVDjl2xpI/g3j1cfdgG
3azq7S6uzIuHGwiC1FDPKB7j+9wzESarO256xpzv3Rcdq9qQ7lEJvhEAc4P6rtsi
Fdlt8dbjV8A9B+G47EYDPiorUPRJ1xqoxuVIndEknaMWdPPlyHeM6lg9PDcmhMy0
KHrW/Nija+TJEkH0FjIEAwMLBJnRpr41Geh4cUCB64SaMW1hA6c5uT7eo72DPT5X
N64X2vvR4c+0S0umTLEYfPpnkaNWshIJlR2L3hD3JgBhuFzbrc+nw6QWe54j+Oau
WSIyUV+oSpkaaWP0psMrvGJTbeH1bAvgPUN6AgHQf668ghpLn7tZu6D1aWfzAaxR
k81bzJnlXzKywUz3+P+QvGnXxQ08UbBGMW7LCw8ZNfAeEUChamgAviX5kahx+VFC
wUI0jZqsjGFzj3PjAwhybyHeODuoL7llPO+mUytQITV6fSGTPPQPjKA9AyP4eXow
H3mG4RWeGcdpazN4hBeE+eqdhEQQ2p8fW4TIY//7UiSy0ZV2jedZv4oLu3ezlMd9
fmCwpw47vXbfr8aOdUpF+2L2CT4ounKBGFQWaAA2xgLKJNgKAhIPkwGQaQukkN/1
wpvx8GZumE7OUXG2S/US3z3TdeYrmBENsMVUx6hMyGuAmKixh1CKqY/05gRlbZei
oRtQSriKMrhZ8Up9uYEwKbnhtrA0T+yV5VnywmFKS9QB48hrBtyI/3l5/M/AdFhU
6T3UDqV5BcNxdznVpbfCjwOXddrS6IlOJn+M37zWFvyZ/m7BdjgD6Dul1j0yFjkp
g7RjEEoFjhiQ5TVf4r0GoqO7/Gtpeq+hncvkAVEqgE1UtgNzwg+WayINV83VnoDF
uv9WvBHmk530K5CasrZaHbgnwkTUJiHgQpRBh+5Rj4BtTZGmusbwJLlOarZB0Hey
FxmiruX825wZixArp7nau7XiCAvyco9pfuOg+vZGVYB2nSRntPK9tADQgL9wqz7L
sJOJf2UgbhxnTeEoAR/YPobvYuEfDg0xJmRArXtKIbPHqjkhD/e6GvOafc4HIjoQ
Taa2C+9vhnaf/1VpBvkQZ/o0uSSm6OLzPJyLQRgD2XoWb6XiG+AY2PynTu+e1sLv
gAvBKJlcbQ278sKByOf3aeCTc80OQDZHKyf1HyutnRkdh73yter3v62/iKCRKHDt
7tIBj45VxekzelVeZVeGUwINWl4akhb7onwfW5xnSM+cog1rVtqjX84owtJaDWMc
buv/DGImmt2x5JBjLV5MfhSIc/tzNXcrs1TuK0ukozE9xU/bwC7bxYFbb+h8Ca2e
adG5g2TiN+Z40Z6UrxngPTtJCT2+IyRICk+xfOcpFYlk2lNO6DXEmoTVW6iok3O8
4VVLJ/WCzzVkdYZpjni3Z7A7Ww29wp3SMATAiYJrk7xjkiXlxr1K0nPYr1fGSCDE
hZ94WLMsBAx0EHGxs4CnpeKJNnZmbz7vAfpeRJrHlWrEjP2CD0XvuH7REPu1PLDf
VBENQcGQJq3/4cqrnW9vVLzlwSOwJ6RBuTvw6xI4/yRWahj8uiCu781FGOY7o4UQ
1iKRot9MBBHePLODjQjX+y4AtW6KPDpCTe/SXhPqN/8JQSlsZayM+r1pfCtlBWGY
dvhCcI8zBxYFJnTI45fXAHpgVMSaFGydHjZV9ZLpCpym9VD++dysCfs6EYGMv965
N8CUiaOmo+sWEc7MORnsPX88VYZxj5ljqcEZ3rgXTKxG9Ru99Pf/GcRMmogyio3y
LbZgU8rEY7jTqWtw3kN7s3sSORMNPHemtvV9Wka3NCDLo0DZGdjNDReqd4L5dgn8
9Tzrn319M2GrI4cpSZfe1rgqTC9sdty+sHa1fU5G8UrDMZD4APCUoKmAFzCzML5c
Cr/FnPS/ZuiyR3d4BzHb1487lajTGA33QCRrXV5kabW71ZoLMQRemGnTHLyAr+4w
wERvArr8f+cRQXe7CTu/rxZUYKweNV9On87FYFbcGyTjGOzKu8Gp9LQSYevM3QHe
dUKyP8R9RW7Y8F+f+b+4yIm/DuhHW0R/HBLjiPPd7vXAcbwBaj+EvU7iKYvs54xb
+Ebx4f0ed923+EELXD92JglGz+eNQwzFuXjYKaWHHn3v45b0LTM6aMtmDEDb169b
ZNK2z2dYhzn6hK6wI65SXON051wPlLSB+uhUAkvGotosr00/VvBfRMgQNdSyByoR
JlIzttddgGdW7aXaGkNNzKJoHw79xM26Ee/8JeDbtlJRSH5KipRsp6qGuMCuIg4X
t26LxNYOJScjH25t/nL3tpXD8gjpWs6a2vUcivOi40N5gAqBUJU0pte5jCcMLAX7
BEvZOovM1E8ROqre8gUL0rp7avI1OVhTku3D5njAWQXz+K6GNpXqABom6hkARKJc
S8hnP89EVlVBrl3K6nfRIPl23JaZSag86CLebgMT4y3zT6zec7fqM2wGKdG79a0x
Af/E5JanJlvB8Qpp4Zgld8pWwjgKSMxdaPGQseVIX2dC0tkx59+a4DD+cz7DTUJP
iMLAqkzcIpm8bBhZZeyaaXFXWrdW9a4/+17TsP47ru67nJEAAioxtCNS5n7+3mKI
GVQznGoPbI1RK7Tqj7YX7gqNlVqZ4cmmRFaTV29ts2t3zN3axyc9O3wOk3/vlZL5

//pragma protect end_data_block
//pragma protect digest_block
B62571qNJ6JFLQtRhnZ8q9RZwo0=
//pragma protect end_digest_block
//pragma protect end_protected
