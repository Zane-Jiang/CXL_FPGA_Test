// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bSPKXOkKJCwiWN/jPZ0boVZHILpyq0ZfAquRDvMmGkugXNUv9WObX40IvaRl
he688+SjFWuz1/3AdC5lnhF0FtSH+zr638j4EerA8U7Q35u9VY+Ulpni/OFr
V7BgX74w7gvF5lmmB/5PNpnS1cKtG3cUsKbh2oPd/3tHtF0NyTOt8+rDoDe0
6QPuQXlaeooQpdABeeVd/mYLGusKawZVxdCRCiB+4yPOAgJV3+mhI2xd3ma2
dDf+sqAjpX+d+bTVCdMc2rJZDcfkvTaFDOUYq4wvoRHO+8usXH9hZavx7uOx
PL7BWNFnb+Y7QZ162v+GnbgnDlUfytrOWnzlubIwrg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gJpNbU26aHO7uMX9Yn5OcMtwq2o1CQvENUZqDq9FeoeY8qK/e9POOgcq4mVA
TioSRsMWS+bNctlkfWLk4T5xLaGA4sIq5Kj5r28pkcIwUwkW752WUY+iOWIR
Lygq59MuOXiL1LWxumdl1jH3GNPFaAU9k1v1XVAhjRYEqD5mFQAASQZP8G+d
tmNSa9Txd6DngB47WJihF5jwUb88X8r/wWZNsV+Hux3Hwv7IyDcuwGFJG5ao
NJjWWbdwDPE2gb4MwzrvjMs2XBXjjkRrRKchNQd4V+7+us8Spmf7zh4akKV2
a0ALL92Omg8wFz0qLVpy+2m690avqjRyrxqysnkYHA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rnI9LS8pt2MycuWNTvq04b59Xzd3C4JFFqFnGlpV/qGe+kf3yk97baqgDix7
kLYISdazpIqBj653xKF7+5M+8cfKZTCvqXL86i2v0vVN4xkQkYhNdD3q1UBs
1LsPmqWTVtBcJ8bxcSDsIkA3LHYAfEpahdIMT+l5FpnqFbCDgbW2k0xdwvxJ
O9PNbMtymjNlJ1Uz70/udXdo8d0v8v7q8OLFQlOyiT3yjX75ZbYNH/zDEACz
2oHJ+U8tuiJlMyJVLeJNt5gTzcg/nP93BPyi4cXVlOYTRGs9ixbFZ8cdxBrD
p53Uj0vM97C4zSM1wJ3ZOwhfwdHgm7ZrReb5Sx6Kzw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
V1M0FaKbbehYedQ52UQ9Hpxk4hmiakWK7Wah9O4Tr0LnOJbKpAxswe/wx/9S
qu8qfOkO2KBcaetaXg1yfZCIwUmkjxBwfP5i2mVAAIYY3L2YNMgq4E2ggN0t
WPYQVpfIN6qfdOHQ0s3z8Za0RnvWSrfIDO4Wrn4SsnC5wseQulg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
D3zXsHs14+cVEEzw+pXl6bC1/KKth2QnI/r964UxTSD7bvvJDi8CQ/DykC6d
b/8HZh+v0lXPuDhTio8muGpaEaJD8ciMkk0DTmIoHohGjJ5CR+Drhs4/5eS2
TTl1EVmyX5+b8ddWWFPqAkLQ6jNGS+flo3CROt8TbpLu9uAzDA4OqXIquUsH
FWk9XF6vuieCjY15cZ19D7tZfkoBIRO0QdHcT3wxu0cTj6e2pLKNpwBNttNw
KWAiub2gmk5ETB4+Frwv8EzUPcqhgd4KTMr79zDLexfVEE/cTUDRm8PurRdV
9UYtacbPXcrd58EpWrLEbqj7Xub/TKRedCJ99Q7j3CqmwVm5jVzFqPouwGWZ
EB8aj5dkhy9RMjvzv/2lKQDKMUkiU9x07idrMWpoRElYWrN97+sqFtTptGuY
+eHaf66f9MtIF2sYHUQ5DNUnDxK+blo6S97uStda5t2O/YJMjqsP6cj85Nic
K7/oQvg4CnjaQ9sb32zqKvBF+C6/mnyo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y2q/wDo+Dp8E/GTQ+b+UhcTxNn+fRBDS/So8FjbXVUW/kCQXMUkqR/NDYZRY
nVClnk9lf0WqWSq+m3Qk3ELyiXQw4Ywoya6QiVEsyBNhwF5ffDyJE/NgNWSk
UdanUKrOWr3/1aekl3hZtBal6xhnHcQtuveAaxlQUuL6D8zvRJg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QNrVcRIecJ8EqQG5Xc+GrspMOH3TMZqWNAIIdt0dMe2E+GnkQX1qALJvpAXZ
s4HR8PDcYGgfh+C+s7G/Inf++1YcU8k4sar12BTWvAyPi6frb3AU5bqzVPqs
jffF3zBQU0QRNFk0IsPV2dYw8KnLvxm4XHbhF+29R8qz+cLYnMo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14560)
`pragma protect data_block
RodhxSpVqznfjK+qWlxAxn0MLfPBBCkWj4iDw/+Ue6jr2asj9r3/zI4Dxbaq
ShMUwH4//XTfEduWdmON2SwQlG7JLs3GJ1WT/eYyW3WIGx7YBTh6iII4mMqH
0CSQnj8eAdauBvL12n3+US+HZXAZbj24ELst3qPLYcrnVeYegQCBsf0H9oKR
faa1BTpFakNcUcgRODo9jw3DY9Il9KQ3K/Odq1yS113OTkqSfuY0W9AY5Hzo
d0Iy7Vp871DGc/1uAG417uKlsETJiuzxtGuXnBptW1llIBynjR9aeWxSSDwe
3Z04kZEyISkXC35Aq+T7avrqf+MIeD6bOA7SIyOBMQKUKuk6QYS1dObjyneI
uoaE7Oi8aUtIe7eR/lho4CvWw+DTe2m1gIqVp2xpyvEA7a2UO0S/oD5Dymik
zHmziIZ2RSre7QzRk6TvfEXUjpFKtoG2gMey5Pod1BZJ8qLaXsBnDEb6msZO
P0d7hqybHYNpf3jiaCdIuySZlg/n7Pa3+aUl5k7zzlv31B7cwj8wleImV7vt
dkKEwL+B0z28b03gfXXnnZmDxgJ4qy4OrbRt3MxvsVL4AVE/diI1zcBSae9q
gSB7qWgCxH2HvCknHsXRE8CUNFgO4xIYplbGTVGHbzzBiP4MN+NOGJhYI6dq
wb7mNf+bMkEZsEydNQj5eSI7PZmtG1BU8/bA+6q2b0LqJISChEX/zh8405Ac
WAI+gxxLiQDuoKbC82FL+J6M20dZELC+ppbJFLMV29bYen7hO1J71B1pMC85
qOsTA/dx7lvstQYIL2mB8Kas7zPlERvuTxqhjFBNOmWE+kAyhz7V7mDdzOy+
q6u0dtnQvOeKjXz1GxP00R4h7S9Y8DjmYUWzC+sZfBM0z6855bVji7w+LuAF
4jlUOCMr1MSr5Fe5ybER6jm9eBXCLhFo/wHj9j2rtaT2UnhBlwWHbqgtTBcU
FLFJaxjrtiXuMz+7YgrB2p1jdE8zaXLxVlkk+cS1zrI56CBdIPg7sfko5nc4
8QAkjXrZXBrCs5fU0NPTnU4oPuO7XqWYst9JRL5AkUSlp3t5LoGAq4Vw4N4x
c5ooSPhW7QCEJuvvUEQwrBJ3yAxdn50U9Ei9yh1J+XIzA/zfcD8P0KBI2lQi
Y6MpAgKINDrfzod369f2ZQpu0ydhYidUn/X/kk1i4EvKHINKnkjJrotO6QL8
RSrjLsYHWIU01mnIMMxt9SafDcrJDLVZI6N3c8UMFiozsAI3GhewCZDnZrC3
QUnfkhHYbD5sO9uOX+on8+H8kuW/TyqLKHuKRG38NnUyqxAJlhmCphTWxvc7
98/2yC4RU7JLjI4WVbiiA6HMR1F8omafooEEeiU/aKf+Jd3nTv+rbxvWS56d
uO7TzbXGnei8psR5NtbmXdhqkc2rCJA03w+gVfFlMlCU6Y54fO1FoEOFexK1
04t10w7ePkn8xbEkNZ6BJVpo942Zkegrmn3xeYYH79iUQqikzXbE9/qhvryI
pkp2CSraiN5xKGjRdsgKlRTAQ/xZP4dcCxLCJAOrkmLSuQATXEzD/P2ZkB6u
o8Rm7QJncIdMIt9JdW2ncOzYBXC9eiuhCShZEyLHKvMEG+B5FJj2O3xS639k
w9By3My8W9FlQF12y7pbxHHPJpFGSGFoS4jKkTDZS+qSqSpvSqkcHgMU5//E
L7tmLj1E/g9iaZ3eeJA1kY2VoryT2t5qKzf8SiTYUIQlnCp0USSkk+aw+nkN
3tBHV/RoAG7Q46b/GD1BZvmmvwMV7+hr6FjeyJ5SZLd9PjI3bya+WmZAWBxl
5whFxNZuxCqn1YNNu2be17QIc37vE1zP9SSbmEV+JfnVmIcen3OWpPgJ/pU2
O3ruVpu5ft3jfaU1u409VvyBT5Aj1k01M1u/8I7vzYmLeA1njZDmq9h0TbsA
q8ihwj1FM830bQfk3tbPqwYAEXREWBUQeNYBuMuTjFC5woSlc1kTpfjrTkP0
uA2vgkRQp5MRrgqp+AOAgJmK9Tifr/y6s99AKLTdDBdwS47HSkQuFueJGbkj
S0G+WsXtfpuD7aXzlwfVzRs8MkDZDA0I3QN0e+penojBRxfo1GFCc2xbwhR1
FpeXJJgO8bFObaHHXbHQ+CtG7QL5gMYYypqLNUOGiHKsdYRm9/opiMyGQrDi
adrrzS4xgGqbQXX5Pz/YANfuZcScrotPdjBwA4O8aj+FdfcDkd1LQoIT75Hr
jOSifGEFK7akv8PoCQBkBkD1tvyW6PrYO3jWbjSy6rLyKL3OGfV4B4mNyCZR
PdptINFlnlalqiTQ7nJsZwWd2WlukDMk4UDqAgrGOvpJmjX0opGkSRnDUZ+s
oHqY2Rr1j5aaEg9Vt+6NGsSXPq4dXpVAFjLOZWbtA5YzRfSEJcVSTmHmPBbc
uo3Xk4VIXaYwDcW1KdGU6W6A4W0OWXfZYeF69eSp0j1RRR3adN0BwEbGCf1N
EHkfKg5hTVpZ7rcU0mVYSCdxW6CFh30lIo20VKRA1kunxuF9/Ilx/UjgNXjH
vT5gSHhNATuF3xh2SjGO1UD6r8aUBzFtpGHkVBbOScemzC/OIIoYT8OWcO40
5nWYU6DWveHAWjx1Hx6si5UNylgzfjLFCC3yJkpOKxemaPyUqOB6kWV0+IV4
PEqKboVflnJARwHK9weyBJfWh2obVan3ehpcCeOHe8BqbZdJMTIOIAFHK+GL
H0io/UngdruNn7ziTYlumceomkO/8t7kstf4cJv8McEhg4u3W6JdtzOMIeWA
BmdwCxwXOShKGbGsHYAZURO+6wREn8puKiQVng2hXU7SlYtKfnTr1Mxm6scl
SMQE0JXsRuM6RsaPcK7OfWYYvkokarM1ZJ9nB8f+YSTN2esVuYp2cEXHxmmj
4pkET05b3MITJyD5CZw7Vv0LBNuHf6FdBLN9NMZOOY6vnD8OtKRuoo3hrhJK
x8K2DU2jFoSIedazTY8/aau/2ehzQ+6mo9R40NoJBfxoemIO44npVZf884JG
3fF26s4uIhAi+fCskS/2NprMlqbPCMQSO9qfpFMnXbeQUO6lKc035cRvGRP+
O5Y/di1SE47nNrh3PuuFBFhr+CiJ9jZNSkaj4SLa/iZnTD2VEhMBGfnAcoDO
LXwiWrxgmv6Cii7a4cN6zHbNW/6Sd+DpCmK9jIwDdyhTCYRuGzOZ17jEP9Hw
MU0sbTe5uJ7GOHEmQL/016faMnnbSdmj4yCT8EnSvn3qD4W2KtJgE3Kiinds
l9SxCUzI4LqqlYsCw71gHs7N1BJumGUY+/NZKcCm2OBp2zX0ytflca8trzIr
6J8oTYi+u1xpKCJBCcuLDhKoSwx8CnsTrq2zxOCRA5HxuH8RxS5uIeXBPUiA
nC1NnYxhXqXgioz5H9QNY1Ukg5s9GstU9FHvOCTrn20Bn3mFh4uG31Gk99h7
w1Am6cl0daTl1DaZd/tMSJBBXAIRn0AoK/344ktkPOEgpCYgXKVczFpws4jr
1GTXusMw5zlWIMOrTqqwlstzZZzYNQwkV7pLMrxNQxCmM0lE+fnkQSvqZcK6
36B2SqDxRfL3bA+Y9huN7xfNAOhK9g/Iw3h9J8dizjtpqT1gpebdwLGy5TZn
4EFw6VVuA02oXqUSs8jfHfit7nB5USZfSDyGiCRcEArjxZfouMtgyoRQHBgQ
bgH4pey2NZL18vLWhaHL1aHPdpVpj6r0hFEYUbJvEaHBIHjrauM1IVQsLZ0W
4YfRXrwoEIzuAuyDvyhhmFDqlRHlS9TvvH1Eajcib5aYR50WH9GEYhM00beX
e4xrusz2ckrVFp3yMB1NBYgCNxSPOjPH1PwTbUObDHTAkNH8aiaLeAgVbIte
cVgw+mr8L4Zi6x4fDs+TrCvwrCJA1UEVi+cCDHKKNuN/RA0qeGl8VXMpvQ31
J3DJIZshCKzj6/TSW3RVVpb1zuSh/BT8FVrdHLrj+w7UWvvyKwXwfUjWkS+g
C+MMzA6WMn8nULJjMUMn1ySeGqK58mvvpagjrNIRTUdBReief8HMO7QW+Pie
9QBJPujjuZWKeMzBcOomek9ZMJFuL5C69+wkj4mhE63DgkzSBXQ+IES2ZcKZ
a/2RSsDdfQUljCGc4QzkbBjqZAYQCJ1Ytkp/mRWm3HzDUpzXPa5m/3doTAb5
vzx+7J4cvDEOxrdoLDLbLeXhRBS2Kx3XVLgbWcm7NrQapQx4jI9z1nTWMtMn
/Ry8+wG8QuTelj7ETgQ/qlEVJN+Wbozu1RrHxaDWbHRnU0qptuqZ9/elZW4i
/Ln+kibG60lbR91bMhwxnkuwF23OcVG60i2sIcenjxAOdwvMCRTJLHOcDneZ
FQcWZvLrHwa8AG8vK2tM+DG3v+s7Ujg9266Kag03oG+ruh1gaWH4RLQFtLpt
Rs9p9k9Ad6iat5l+AKzmVdOKmf3ab2nSK0QmuUKMTqZURV8bl69tR26XWTB9
bDGyQayL15WzRJFTvRwGQu9U5GGqqZuEaaUKtjF/4Ng8ua1a0AacYjvaqf0+
pGGLrKFNVt8PbVAfBQWLeNQnNXdTRncGAC8T5u6tQSGbhZRh7U8Qcg566Ie8
C8EO1LILp4YaA3d+zot5dKLeFQ+OLdsvN1wRU+HhnUaJA8Eqr878Z4f8q/ZN
1FeQMlHtXNnYaqZU/DSu2RF8gKvI/vtnBz/tdF1jUkapRth96ZbQDJoWa/8/
XqdicvDTC8eZ3c9c0e6rc1gNMxqyyhTP6noLuqP8QyGK92laRxGF+wHIOAqs
f/PHyRF42rUvz6pVKMm/flbyuv6vjnN0AZNFagSvJpnRGnoQnX+wykOhdK4a
UjQ1MhvqL2d0x3anv5wk0TPhByj2ybhjDtZwKTSo+udMFp5yCUiVhP8zKTof
tz8wfYm7uxu6VkWlOsf6xw4sJ2CyQhaxKnENGEekMoj1OSpQh9eijvjs5vH6
aCwYZGD1SP0YMwUw5r5Kt3ee7YJqdzQTgFbBXPkq9HVKfR5qV/OegcoKiipd
0CEzgAZQacPDE7PSBUCOhpeASeNP7dquk3qhDobeykEsuY2WKw4SCD8E1upo
RVCoeVD9LTU5eBRQ/+6nlAcIwvPjZM0vXD8ptISwgTVJRxwp7NZsHZ6bx2Er
PGVjK/bgerGgTc0GnzB4nldsWYSt3XZl7WgOsYZCtjyGp/y63HDwoNT7BrS6
3XfO1+dlX68dQqFOdIsBISf6fZBjYmk5G700X8k3teyqZUUqDHReHE4lt/yb
9lcM81iW+XuYg7xeWTlxZWgZTiwRl91iDoEYXtKCf8NNEohkektIf7eh1MHG
Lr77SH0XdDhVZoov/+BrSd+zW6oyAPJEtlmngvdvCUwimZ3/ESeIpN55PN3R
iJYmP3ZBFtHKMbrreRF+kDY6B/OTZQ5up+FfjqsNMtKB1e3NP7stOKllzhUk
dl/cU1AVma+lsEpPHuqVqlIYM0xJvtqS0AwG8tYQR7HsAqbdHiv3QLZO+Zz8
F9ydQKyza8XaVoyNGft9nmhFNO2sk/ZjFlnLXXu4lWPAUshMqutMrHhYrFXV
T4by3TbjvEW2SB7RxO4BWFrIXcsMLacAmul04vn31AiBX7ZYdDm2KZArVUcw
8OIo6pKgAlZcoMZ30IbzaAFOUSqn2MQA2DqKG/jlmlJ+RptVHfm7igBFEaWg
t+TqGksh64Gitn4dht/lE0h2kBotyr/Z//rwDkgh3v68rIQkAPciHZow4Wel
IcI6Sl95qGt1xN2dVLzQKTaqeo6s5i+QobVE6wr2MtZLUFhTI3a/ZMn4grtZ
73A8/nV1QW+AP0XP98576KVNcsazjNszH2+7TMgYQB6nTrKEULKVA5o28kom
uMa4nsBUuzJWCt4Y7AwxzI5fgPBTVTWT3wdnhl5uFJhqJ4zTJTnO/aTXnjds
DIMlKFTPV7WVcQMvkcV7nRLsIVRHYFtHebcGV7IuMr3h9tXhvnwOj9nutZhT
9SD+yavVj2G2znMYdJiliV1jl3r/73k9FmDDKBaPJVmY49cSG1YcAZuKBn97
q6Bqs/gsOpb/0L8HJFWHMUFUHa1R8etRVLX/Ax9oGBxMPDtBkV3aXCObbZTz
fC6onNlSBHag1ab/rQc/u2wvBOLxdCEiw/X6fALrIcgxgseOE11NvXq4PLrj
KPdIchPq5woNHyzoQeZb+gPhKx5h15IEa9oxYqX/H/rN+n8h0yVinw0yP2Ir
swge1NTUJvC3xIArMWL5bGZU4nNDCITI6uuSCjztHzlXu6gewjTl14E3gl8N
RM1r7vfQLicsuOZTfp4pslvCpvpKA/lwllZuQig8hTHTPAZ/NaCQlMXgsMHH
7nPx19qytYfu92eKaWBtJq2qj2M49qi4gMaZPRKsYY18a9hQ9OtFUlRb0x1e
uGD/oygf6eC6wHZhmAgMTxWx/abOTw4/qGkqUsSsxgv4M9wlFYsF+ioT85Hc
RvXrHagbaS0tuBmlESDGCDEjtGE9fdunFDY0Z/m74ZkkjiNzQRZLubAjTwif
722YrIDfdcFbgCONWow8S1XloHR/BybtuBu2qHVPrEAnYNuI6KWGBzgbINzI
DGNiDCLiR7seahxkkTEve+OxGd1ijOndAR02GKwHlSDdp/m2TF6oYe6qZ5ek
YGu97TrfIg2uw4D9FGySwzB0HXsvwKUrlo2kuUcc0ocz+kQiFquuiMUCOoQt
fLPrP+GF5qpDZQfkT0SG4C8fG5TM3eRyZ7XnfoqTCvDHzrTSpcUqIQPLsYzG
uNhretGTkQ58XzZIjmTs529W5I2AYt+IeF4cKbcpdP5oFDXElmkNGonJh2L2
eUUWfI8ZsR5tdLgIpZTWspVcBlR/Ii2EUjpE6AjXjgb3rDdOY6CDiIHCFKmA
+vifN01uY9H98V3HzmSeFmNjnWnc6ZEh3K7jHY4efMFcng4gC6yTLPh7AZzs
2Q0urIAOceoeyhkwYMlgm1sOnpAN14da2BykhrxyaIhHRQdf8wAIY6AHhYmt
k8kgklis2WmIME+TGJvRWntjZHFmC7DDw/Huy2FMkbE8MOYrq43eLhorDhqk
ff8icIqAyTAmvs1sqZGfQaUU7pWpkBHRIrBN9By4dnqDiNeVe8/yzxLuMV8n
WcwPw5S0aorZ4Cwr/rxOcfTz2kUSO2pdZYAZbctKiFoVF41G1/JFiZa+KVdJ
mGkTj6nviulraVIbyivuLW0yUa9zEzlKwOU3NJgEdzr0DUug9Vyw3SRVzBGP
dUw+m/vUWTU0ifkpkPTUV246FHcgRNkGeI34vIxXtqVO4CsFXDtXVGcr7ttB
8Qgr4fF+HXm/fAWdCiaOo7u+aDHSvml5EXRLM3OJbcXRHMxVRnP/abCs5qVh
ABt0cQYQulErTqqeEfjzuwg48dzbfeHfg8zBdiRMXIj303Jz2M/7iGkcJtlP
y6JPNK6X4L5zLAoUtgkJ6h2oyeq0+apA+g9e95ukA3qIZcVgkK/PE7Sd7m90
zjKMczk1PV1keYRiDqrv/WsgNdUJcATxaikDiz6bWCXMWmdUFJ33+PTJWo22
H93uZJr7GDcSrMMve5kHpEyfZqKyekEMy9T/60UkPzkRAFVFiaweWOUjz/io
p2gtPKtAV15gUqx22ds1i3q2d16MAU9ls5+iHG4yctPY1AN1M23lywyDJ5Xi
8l7jORQ91mK33TQnNIt2p6k/ZPRirrrUvPCGpsK1uIH0iC1a0tLpJaVxR0fo
8kJv+MbTkFRJuXQqfKzcpcvqs8ny74ajz8HKSyN8Dato91KqxdDiUC+FGB/K
SanXc4kK2lEjs+RGb3zAv3hr1sHbHpdeyOvSojEPHmYf4frN1M6IBAJdGxU+
o/urxvheJVyW6MUJGo2ZVaXsFRHQI+e3DedqRbektyA+o5CgFBJd/KWVqsO6
mBCX7dgLe1BAaAwCDfb7kSSFazUkzBLBtg5tpI3qxN6sBA/+hvGBMvGUP+XG
iOX4Z0qQpzQhVj68EDe4lMGzpBKD0V241h6AYPCRGI2s3b6RM6O/n/94tu6M
v2GCXoE7JdHQiVZAqAcwkYm+dOLC1bBHMiQOj+2UGTW2gK0EC2yU1CEd7iHK
xIl9jxi87939sw8CsE3SX3x0Gbaf9gmF3TP/c0Wn6ZCpnSdWuRPEk+7ejvL/
d9m3CsOQFFlrlaBMujB2rhwPhJOAsW9iSzd6D35Iqqzv1xuNsRRaxtWF/6Wk
eTrIUWKcA2S5Z4gXGcTHo21/4B6/ofcKkCBR7X8cXxzkz4iknv4z8E2UEH/6
28PMB1TVLUPB6unDOo8AJ1PWrL6Vn0ja+AVrgMTh94lXw2N9nrOrUiLlfJ6Q
9RzTJIssc0YUjZxFieabBpyJbxaJBQ1SnJJdJuy9hK7PuzMBGY+OIl1Az2bX
sBSzTzN5pKIqAr+IUo3sQ6e9nTKOaR0kmRDZ2oNLWbjS47Ox0nP2FbAdCMky
jk3lChJdsAVY0f8v0WLfVcrYdxXZnIp5Dos2BNnd7jIwWRiiV36sRSdJexLj
favHsfg0PwemsQd6ZitOe9EhrfEWKcnkC8fnblocbwTd7UVbyX9g0Pgn3vVo
4Juh8WtbSKKt2fgNxqQjW4eU43THBARdSQNejl4Erg5W15TBjIWFmKVnVD6I
F7eezIU8EJGYgZccCPpHrvzDhIofUYYpXC99eb4Wzz/+YDMNSeHVuXDXtuFX
dvN7SiDCXT8AHynZPSFZk+GlswEMahwtEHQbTqCBD0lprU38c6RgILRINVj6
FyhtL6VCYLGJwshYU4XZSwy9fuz0GnzLwzEgXdIHi9Ny6O4ODU7dnmfkf3oE
dj1uYZWRMwp6aMixTTVg3ycpzmrYzVJgiwmoeaDO3VpU1F9KW9308DcQYLmg
XYddBf55QIH/qpxXxrAckVVXftL4DiC7CwH1R/Mb5+/M0G5QZ5ZU4J+Rkau3
otHMy8RhJVRXUDsed17oUyxdaIfUGOmmB3mY7r45F0XwQ28pJa69qOu4caII
yaH0QMx2/Cvd6AUOtAZmsApdfxNyrYaCvx1vYTiFTB7kI7AB8HBM4z09hLVB
zOSSXg9F5iZwUUZZdu5P8/zTwVsa87EcbX6Av3ml6iB7KwHgiAwCstawAwHk
w/kxf9QfVfiVDt5/44qpM+/ybysVv5PECdSYudfY8NvEOyu+rUIM0Hf0qrQP
JpdzxW/NsrfbIcZJYftCRcGbQhv9TH+MUmBBKWVAEjaftiIlsNdvQzXrtgvJ
FVndDk9nRqs2TfPxE2sak/VosxxJLj4mbqi/kQrdFByOHSF0UetyBbPnQOVD
Bzss6bdggZNkI/x9JTjknRnwstso4dvKUEh0se1scLPPlFLNQSBL0aNNt8PI
OgAUnXeQwzHVMyQtDH1ZClZg1NRWipahM8FqQXCSTJML+6QMtAjenrRfUQh3
rze4t8gUxpb0rDc1CLx9WSIFFBOAD5UOeVzK/BaHjoepNvcNEGSHugXrKZOY
v6ifQDWghsE0wxQDnGwZAqpcDS1iAy3CtNwzjKi313FymZpvQRbdrt7QOU3X
lPP0FedA7tAmkCf/NmTUPK1otTEoOOUZK1VEgHTJRr8AkOWRLajp7aMFC93m
dZkRqdIOLVQA4OejznnxcV63UTTKbdNulvhLVx7CF01nz+SWiL4OCYQrsio2
VBZ2BhXPJ4naeLW9z88rpkL3RMJDzc+awgJUbbClpFpq30hWL+/mvkTPt84K
buvaU0S/gobjdp5VL+pHel/Hs6uhrreDeLtJrzwveXvG9PA6Z2/mOvYGT2Df
vDT3LjWfGhMpaueAvTxonKPL4Jysp5HezXfYMtme5Fd5E8wijzeqVEyoYaTg
+XR1Oyb0UIbvYtkzI4ZvHyp0sgcddHDrv4rUsIIgI+UEuNg90YsSdQsL5tQE
USkeMwOg7j+CgEpfToOtvZs0A+kn/K7wqvsS/VmPnHbP8Jp6X8tnQ+2u3vVy
74r6HhQdxrGGZi9qAIOltXnJMLTIS7z0a+Dto+nqsBvuRBQ4enfeD6lzVxap
gQlp5J9XIMK6HcfnrPEJuHSAAAGC8wmro/x6iNRCIL5Ix/yEhsqETRkuBPuQ
1yDpn6uXhg3ri6hB8w/tzH86jhmbU1bzPcwa7iQNN0OYqpaxaWkCY+PwR1Ev
ntMHzVOUOsWtMT3bfdVFFv/jSoRP3LB+Zp9loeSRZElxGYugXbkh9ka5oak7
uKWm5gYgaFrHNPT+y5t8Vl+gt5QLpKW5O5okillWTrycpacEJgM2Wm8pLNxA
bXM1dS5VN0eSKkh1mDx2yhMzagUcUb1q86L53cbhrvPuh7djc07mTNYdfPXd
6MxRU2+Zm8mTM3Li+UIsApb1QlYPshNt6q5KJAx9AS1rYclQLhbErTtcpoM9
C1Kec5mFDVtqK2OZvGpNB2c9qi/MZwnuA7kbRt878hH/EN8kmVIyfCPKvcSB
qLXD9FJxJuKUJGZD4qfOnlEu9bg+OhuF+dlcXkrIF7mP/wj5TVDCaIIMWfI8
jpy3YTJp77oZYb3i40MQJYcYP66etE3iU85fnVm0nP7Zs6E1axtG9lG5n33n
6g6chg/PTPjgL5H2PghFEddZAjcs1mqSbe/McQePZWoslamgeC6p1oMv7qkB
Y+p+51p0TIeoZThd9dXETJNIgooZ6V5KBdJxBxjZfU/oXPXFAJeKZNefz2an
nfIXGR3Wl9ELSaM+K7Db4YBIk9JKSsIxwNMNelLqsZkyy2Heh/ZLpcm+WaDH
Nw2VBRdRbQrG13shoLYRKdmO4JQ3zdF9P7OLYo2KX//5dZO2Nej4GiI7mgMj
H73zIGFJ8V/0eRyqQOdxjUhkVmUE4qEvixEXyuyw374n5v9SE9jsROOHl60Z
WHr3ZTDSyHu+8BDc/pmZBeodmC/arwgAm9/VKx3ut+Au2qqwS4Yt/x4gT9Lk
ujqA1vNtDTLLbvgA/OqgmGtp2zCb16ZWjfEdhBk6em6rHqztQ2+mV5WBtWRM
mbbTCVhX+xaqZ3Ob44Z34b4bRZ801GxEOdpwFtr3I57q/0+wv/Op0MH0+U7s
wOk5OUoPlzZH00o4zeJ32K46Pw+9FDXuyUcg9wkz9Qy4GxtfGT1tXMOEiBk+
5PFm5r9Yy4UNomXhaczQ2Ui43VaM6frJ5zFcsPRX2kg2vTE+JiZFHn6mYr+5
BzhbGVhQ/feOS9mopCGQjoLvrpeuP8/dVOxw4bOYE/SYPgG/J1lnn66dq1tv
9z0fwsN5xJN3BXBaucqg86Eb6gJWmH2MU1VHCr+1EX4HSZEFvthk3x2GITiV
ScL8JAfUfOfEH2mRxmPSYWsVJTPJnUfsmdBf7tcR7uAg0XLQJMeikOnTe/Vs
ZVMQ03MCfQaJEfJPbLYaErcD9u20ZygxzJ7PXnWGGftmMRwWXIjiKHv6QNae
EAtIm6GG+w4VpaQbgfjOgOPhsQITYPkROOnU07PzuT3XRGSkdbhxpp4WhBWT
J6gVw2UYDNGVaSlBOCrm0NZjBs5l8s3rf/eiwNWgp5rZoBDMNygeSHgfHJM+
iDkcYaY95Bg/E6PWV869E3W4g/X5KI4OZ/MGSCjrr1ksHjPrKSCKjRDlER/a
0Yu8tLVEuwrPSOG6vrz3c3MWcIByW5EtFe0IhojmreBPxTnjmCLMZEL5rdxq
HhkNN1+xZui0gZ3QLxkLPl1hDig+FJxK4d4oEeYriqHHhgHZyVtRPyNVouFo
koZbeWEWy3m9lhGldJ/XQqjA1RIK3Ebp0QUO4T5BfK8dz4nRErk9YWn8BkIr
JbjLVveDHQXIBT/hJwMTCWSonGmu+v4hlLtRJVLGlFT5cb63LydCaVxbZcPq
IwyG9RFVP/T9XqV6lDvZ5XChemtnkQXrEISsrJpNFWp6+O/RCER6vR75hf3C
GuwEu0YUx9WKO2ktGK0A8PdjEkdC41JAtiDyBVoVC7/IOaPnXpRWN3pskT5y
k+ueO/3D9uioIQM/a/iRsEc6MfDYlaxo4Kk6kFqhGR4sKJoboCy7yy7Jf4kS
k2YThXZy9/j6/WbNabxeHY4nyunnug61LD3x5VFP247E3mkzVw+L98hJTcVD
/+OA5hayetjflbXBjOAKrH9quTstyq7oSJaYx1GV94FagD11ZpVqaMvvNuas
HqHMgUvi+Gg8hL6E0Zao8ZtT9d6jFZUtL+3/D8UjdrATzL0WiGyy/eJ+4XA/
oPEdHH0Lo5aFkW0RGMXtfmahDMa7DpZpULkCUtw2LWpmyOBlzvBRbwK6h5FT
7AuR3dhqUriPm4432CRmTGPe5JwnDObjSfutUiwPrraIVKGcpBcO8u7cCMdP
R1Mrle5Gu/hCAnaGrgKFc2XjcuHdq7Na9fgzW7z6Lt0wdmEfJkOBetbOgZ3c
IepxK1cMH+8LqUC5wMh90vHEp/NPAu3q132E/azsCElmu+2BbXpMsIxCZNiT
MTPIqskHhqf+1VnPDpa192BCWCWUeR6uVrm1FMR42bIuAZ+XaCF4xjxVDFv6
/BVs4UVUYDMIWYR+ZH2CFdro0+/qxobescHRakBTz0ionBkYR937pAGP8Vi9
cJd5OG6QpQKnaR87F1JbOg8+5AiPK7VpQsSp3h3YH4BI9dzjnawo17KAu06+
eszy04IFrSo1p4yPWjg2hk4HqZykknyS0Fi86t9O/fU3km7yyi9ur6xv3g9m
wTTJzI3Kztm4Iy6iIuupeWjifVYoDWxE25OAyvlWr/v7ONCyOvPGSrIWzMyU
r1JUNMwy38M7bVOk3SgvEw6FdRxRVIOc259wpwAznsZ2UjagaT50P9cpMDvD
OYDJNb6FEc6YCymp/rU0GTwY+VpazD3VyReBmFE9jW+Mi9eygqyaeQ9VWLum
dYPDZyM9XohqFP5ZCcmosktsgNQ03uY2/0BzCDranBTIi2GVaC3OU2G7edwh
ECE4JInPGDQuYbZF9Q02QE+Bc4dxklSvZZNNew7Q2LbRq8ELSpOlxqIz0rWA
wySW3sY+h597R/rgQ7vT0Iy+gV+Hsl43i3c2p4xs7CX7INOCRHSGnbYizJoi
jlp2Eo59/SqCKgRPoauSmjLCt2qpcZnFIZU+ESm5ANcXDiCRfyfUCG+hoWlF
4KHfOtyOdEIAwWI6p7ui+zrOccljYbVQeQKkS1N+/HbWgCtl/ghFW2XCy093
AUVgBsTIKE3dU3TgVytuUVC+4fXm+MgsmZifm0NjUfQ3dINwTlyGZQni6tJp
i/g8KXpzY/ICY9jJjDEZn+A/v8HtlNAZ54iUchKJ9NwjuTbsnquUPE4q6fOA
GAHpJvR/HLmFrbv5HzeHMU2F4xaJgAa49dh52jmt+BgjUKgudVsrXdvJFz4e
JNERGQC3LDcKQJ9SSo6OKCRd0L5tO2cfKGF1GywPVFNbpBcrdE9wk0Xvh2n5
6Vt0uv9eS4GXB5vnYi1mlmTiF833iR1sol6OKslTfiU//NkYYjm0kiTIg14W
iN3vGhcX7gCmU58UWzjveV3Ca42gUMVQhkY885HWw117elW7QSe7iwMyGLq1
Vk+DYqHOJXLGOK/rFvbfhheM8PB6ljEXrLw3+ur/XvINCn3lrcCK/usXOJkt
rO/jCbNbhtttkzrx9tyFMt3r0Hky2zLZf8TtFXsWRLrftwsqt3/w7GVrO5Wp
BHXeiZNlwucxa4+RmIbvLg/d0F6IrYNKqfRTDUixW/rkBxu336vGS/I1BMgI
qN6qz+s2xThI8IytZ8HbUx6r1tI+KlN11xYYIP4XICCbl1QcOdpfG05jYffp
1XjfUXg90Xev7RJpCFLbJaqSuR3iAkQIiIIAF5IqY4eQJw1UX9anr4KrzsWS
kGpSUmLsE3fw91ZWsbQrHaTRAC5/Bk7j7Kw6033M90zLT4EUE3FfDMfhheg5
/RBFet5BctRBX4GuUm+wKjjWk0SdRotAQfslZyZmwRyDKxI8OfGwbJ2XAnIA
9lbEdqBUQx4tF/7uxENorT/qXZrE+Jy/Nf/AiOH9EHmRSalDUBPvvRXNAF5O
/7lXvuritdDIIO14b4ahou/tk15vFNteU1cFVYlz4tNUNtDjobVdzEu1Qg1i
pcxPnDUWTIQOTj9+W4rs1h8o0rTxPz8Y5dClYrNyp8cq+j1QPZxWaw/9rw8s
zwDaJoFvN6Q6cDgVSgBYT6FJ9zoos2miaqJigOARQKuoek1017EuZfEZkmQC
gi8MeZG9w9pS77Zn30iTSkqq8I6Ey9ujgB99pGjMsRJutfI/FHE7jNWSymM1
ff3dGTy3WL6z0EzbiQl0tCEvq3hSkCpim3CuxpCALQX2nGWxxVT3O2KnBJ+p
NBqRZ4N5MEmfJ6O0H90PG+p/fl4rSjoQpTt4UpWp+84gY87SeWq7nXGKnWWO
UzZjbin+c/xCN6DqSvYEVbN3j+QVJQYqYnWmHZtQmPFsxdUX8lOIHClUqRSH
K5jMjalJ2iwneTrGoixWUWHjb63sGqniSRRbBKFrjJ9k9jlzx2ULULvxNudO
ZpStLMmqB42krg9EKQ60SGdd7PcKEs6uRfMKMoYjTJCB/xn/iqDvtgd5ZN6D
U4fkS8n9MsFGRVIx96kY0q3eCa84mSqLFGaGz2OfDUZ7/NciiDuSytASuMyG
foPmz9ODUHPqALggapxFGsnyBePjApV7KgahDeGRH/z0u+JlSAG+thSKCrWl
QaVEhuUPned6Nr2nFJxBloah7NTeeme5xK6tQN07L4aKIFg0SDr9G94NhqLS
5tArRwCC5nCaLKZYAhINHxYj6Wvv/N6jz4Z0g2FGm9IkYsovaMmGvqtG+raz
/fW0/WCNzaUmJ+QlMmLRLuystGD2NTYvmy9PcTl8Fxae975SfWhU/65dpVHP
roERmqo3ZzUq/XXJEV11zdkrdGMmddfThNnzAJ5LDLkwTioDbfOxEWs7UVyw
tt9e1ZcVVpJmrE7yAhbHpo9kBWbCceihYasjKL7yX3arBF3zTjQwiHAkqr4p
PPmo6DPOsvRFk7K5cqQ5q033Ly07E5kT5GweYIORBt04A76txU+7Mf8J/+EC
s1XvQzXL8J/i+V3pyQBgzSAaW5HpBZ3Qhr7S0TNkYdffV3zMv2l8C9fiE4vo
iV8YbJ+Kr0jltoTjBpNy8KA1hAi4wloGqajXU43gJnBfz46puQO7ilaTS6Ja
Xvm2m41FSIY4jnSCGNzMGcM3y1Kf/9j6qVHmcQxOxDZF6CFo44VrN2DJHi6o
p1Q4UW2f8K14ebzi84/8UoGAouJa5ttUYana3rtQmUljjkyEhMIH927qldMv
ZVO60oseSjWfnkrMQQgZfrnLd3Q/odW5at2h/GRH3G71TJcRUKROD1eHfhXo
i6ZtZN76RrOf+hLOacnkAXmJ6mXJnyAzkJcdZjGM1UQ7mUovKzFLLQY+CRMK
C+cTxS1TBD2UcoxwPx/xGoqKJcd9y/k4RPf80cpuLMfHi1G1e6abtXJzjuuw
2+nTQjrJ3FKt0laZEE4Mt1sQM02P61jBFboBAn0s56FNs3gLW5xe605pL3aQ
qJasHKp9KeuQyTnLpb9vmKNX+NTVK8nDbOYyLMUTqsZcwHFOVIHdYRwHoy01
rEcc852JYTmoDjrkOpzDA9vLrE0g/peYsbODbXg1Sy/GWwv9c0epAyYSEtXr
ZFZs5l2aFLOL7S9VFDXBApyzvDf7qUtQGUtToOIw0EqGj2OUfGNZAlRW7Q2E
37z9fIkiCBMqLL6q0f9pxWRQrZzlk+ix9CSyHkSoXJ+1zyXO7lV/BiU6fZr3
eMbD17HNKwt3JNIJiUWf3va49+A+tEF1ZYDqqDR9Q+xGXfoO4DD+dmQtruTF
rQ6BfieXH+eM2cI1/4wR5EJ5fZ+lD+zk8FRTdDZD8XqSNwtQKTh30amRYg/I
y2efK/RvwUzTVX35ggZ5WyVmvKp/2JVllw9MCTwdMR1Xu41o8wi0B03E21G7
Oy/PSnCOgY8Uo2TqY+xX7Qsay7Wn62inwofdG3BAOZnegAeD+B1dHiEeJV7m
FOeC+vH5BKaM+yI2oawZdI4KHk90CQZgbOl4ogygGeP1woDNYCuEV999/e61
qr/u9CVatgQf6ajCb+5C6l3lvdrRSA9zDZYUJqxWFY+uTsleEReh+guNao6d
pXjQxd3Xy7952Z6ubIurrRataih1w4aPCWzsIPPY+pSHCuQQTXr+QsiHfBMG
/vDE+yymD3EP4RtikrWw9meu3sig/GLoeQ/ZOK367yAzqlOMEHEZt2upD4vh
TFsc71o02QE4ehKphKUjR9S4THtiu2He494cjfZ+pbqyD9nrnYhfmpjBVwdV
No4VLnEvWySh+wlEngEhtka598yQQoOCJFminLdEQqv0AjQ1D5Hy9oPEpTos
iXY0xOoVK0e2OcQoe01aZV/NggVP34JfpTMQ/sFK2HTgqQO+NpY7QwC8cOOb
8GmEdEn0vuZxGv9teNu/+fXftm6dkzTWJdj0hKhAz0Ul1+ibetj08thmfCwT
ZZpxz3U/OgBiB4Q3ftT8/aDUDFbnP2A1ZPJskXvzoplNYx6sIJfw2ObIdov5
5x07LRiI3Mg+1PZ/fIg8BnauQIZ0mjvHIcsMSnJhAuwusvHWz17BAf+Lck9S
0+I2K8r4i2LSzi8dm1wYRWCeuNHw8SL0emt4Mn2gwNZHp6paXE0DlGCgNe6N
wsri0nm136w3IWvSqoj/UywnBxzq6641hNYDBjGQ96zbmM38f/NFuJpaCuOu
XPJRZCpwy0LdAhRzSQWxRgdkzwowAsEoZkxVPkeEmKhI51GfWoEYRZV1Yxjs
bC6LX+FY+C+8YBlNEBi+luY+cvgZXjCIfo4E3P6QHoO08bN73jExdHlK9lN5
mYhrRKU8SnVNOklWUK9PpwOtNQJX1C9UqH39nMxC8EkrZnjfNAvNsvf7n0Oz
/P4PyWZRHJFSyGc0X86XkEXKU8vu0wSlIkqKutKNdeJRYTkdEGZSkVEkUsqM
0iZSDoOCeQPATtFgQyFa/zrWMXOUJvvUxWaWMgUlTtAjpWsc/lV4G92Ve/0k
K9usl8v6ouzfe8nGl2rfa4XG6hSFvmloEVwZwPfaOcSV6NW5TUBM8+74UA66
FACRT4y5dQ/R12Ok2W3z7knI6kvTndnexnoByfqbjQMVnNDRXPNrA8qwWUCz
MXWgYt6yoouFxOGYD5KK5e8U0g/9wvM84x5ow9zbU0G+umq680iIfL2xFeCf
pWB+NVmlL9bmaQ+IKfz0eE77/aye3PABzcKxmMEpaJQM+8+/UqABxhQAAY9G
rBb8gHR0FEwvE4GMUjj1LC31h0hLUnXdXP9Fz2ChD8hK9sSAgTg8OSxh6VsK
8jFg7Gy2HGrjX80ZXxHYqP3mf+B2XTOcCgxc6HTXc8r8lWvKLAuDhC+PxxKW
tAgbO6xoLuAn+tSaaN0XTrxuueKz7xAl7eibRCe4Xapn9sp8oergnQCU6Z6J
7WGXaEMSxkganT9jfMZvOWGtiIA6eqpqPggV76S35PqpoPKzsgHhzTkTKAhI
GwKtwAOYiCJYv3qhA7+IHBD4aAwwTPxjaq30ebKVOOJEBrMR5DftNwtJ0VWy
p1T/PAtq5fOPec8Tv1ucBRcuXtVCE9Cs4tzbM9gGgFFQ8edVhN6Ou63xygZx
aySs0byz02rJu5jT0/G6p+OcbLntf+BAZ2eWyz71scWagxtL+LWqvwVviW6S
Knf3D0J635ms9XdoOCFdrWr19yAn87lrrJlXQ2B5l4uNs4szr1Nf3rfsTqdX
gPk0j3IFgavRGYHaFd7NwpEfPta+uOVdMvZB/bcYEgVC5E5ytjCUydLSjlIx
LPc1ugwtRZR4I+moAZu1cIQ/K7zXeucY2OH+ZlESUxqPZmR0b4Mop/LOgzXg
dhiFC/UzH0wijbEzPO234HpEMoh+Do1joN6e92vhc507X2q6UNyOEoxcqDO6
Nafo7MMqGQ19tQJZ+VDG5eGgJ8z77/u/qWfaR7A5MUTo/ZgAPNebtjeAZEjK
UUu1Xekn2RtTGDlfTctlY8h+yzDHMNsVI9zKcfFpQRAvhr5FQRmOh0jG8dFV
LAe18jQfHuuCg9fRUu3u3UkwimiPPJqnJriW4cX4IW/bQ6bjk/n8I+gvzUpu
TF6hK0fEGsqPRH9JBjVIuycazpOI+eqETeGkcu0ecOS5fO26I8p6IZFmXqWs
GAPQZkksH9nQszE/WdakYJuYLw+KfKvmIgRkiAEv2Yb35/AJXdwhY179nN67
P1srngkgD/0i2cIju+0VtROClEtohc4xxpsdIK0TG4AQhEoBl2bfpe+1LSoJ
lnTDu/zIxU706R7m7w70fCBkb7hO0s56UbnTjk7pq1EOMcBHCe/K86DYF29L
/d4F/zO+phSu3hIF2kZ5OleasI10danddBJ/Z6hWFsBcjkiO262H34nHJ+ig
OW/jlAQqkNJYCPBvLHb0mlxlBI5puexJD/y2B3lzeZ9fCk81xtfTWIihSZ/r
BtlCY57KgtDeROjQeWVFLDXG7RBoYw4V6eNp9ROQLWVikTaJwtzb1h351D7S
cCsPX5XDlSabiIeylCt1+tdv6YYCQiYXWbucHc+eUjwWOv7W1ziNja+36BSH
npF8CRKfxeR2qCwQ4ypnTw/OZIPcxSnVxyozTyqH0x7rNASqJKUXW/JQ5N6s
lE0imHwFXUg/TrRBXoooJYFGprT+FN1O597VRXych02GzMmvDR0iuh7ajRmq
gV2MSjf7WhA4VVZgz/8RkbgMYHxfucmJ404U7Koy+ax8B4K3DpmaG+dVJ2UB
zPqcC/SZzJyZ5z8wUcdGJH95+j8TxPprmHqDfb4b7w6IIJA5qQduMQT15+F9
Oy8vi2aPTMHF6L1qReLovx5+5mWvXrfTVtkXeV9bFP6scSv6KfL36ZRh1ytc
EqPEUsDhV0m4h1iJ9dA0rdIsEQlZ3HQjt2xXFbuKNUSZ2BdQpWZVIlSSSyfL
6hjIhu7/2zAya8OSlwVhMZ1YEPNP791Krx6vNu8Fcxn0zkIfbr2RQRS3e/8M
jV/tO/OXSSd184xxWTobvEdJCa5/WUOqnGXd/Sa0XJEwIRwsCzdYXpw4c6hr
bEKsPYFYDV+7r3DLQhHZhD+D7DIapzDv8CDhjp/0US+nd/+Jwqdv74cHqMEE
dl1WSwx5UFiAICEjzs1P8HUqibNkwFAoyUNKGJvZvFbeKdfueG2iRcx5838Z
VU2phSiG+winnzU1dniR1Ly6UGrnoPm67MhV/dF7e2UAeMvvPHA1yZ4390rk
OsnxNS5K9W9pkH/EJ/BCQQc/ZWNcXJG78lZ/DPR6qKASVehG1jqG4dqCbNkm
CMM/bDMDMEKVz/MCjJZd8niaeNR1qFHu41orf69FnR0/zwt4bYUvppEqzyv0
h4KZm0I1jteT+qSThnhV/UFrd/7omCWSROWm8vbTJ14HgX+Slzjxz4rClXR6
3kqrQLJ4C8gbbjQ5MD/lWEPEH7HnrzNtRtFDc29BDWtpbyF5RYrBpAOel8YH
gwlPH9hTYJ1yMbP0R4HCSvPYqDL3BkhEMQ==

`pragma protect end_protected
