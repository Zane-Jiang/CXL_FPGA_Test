// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eA1goy+PJUfyGs2vyOlJMwlDGwe1qIBmN6GbSS0QsmGr1kp8Qwy+qjuoV/Il
J6nRbjWPPR5YEOQbvwloixYx6wu01TfSdW2CHoi0r2ONYHm2s2F2fb2LBxu3
lNrvR7QvbRmmsy2XY9RzaReNXTDuL5CW7ASlfacYpAusygJPmNFtOrABMxGR
R4TebwNfcMUa50ePaZq1ECoyn1rKVnjGyg6sVFWK0R71xqtc0fti2k8cMUoN
xrqXI/YMG8tQqJmEhifeY69HGkoo11O5EoRx5Z7meK+OnmLsR3EHRBqBKOpI
jSyp1jjTb02O5LBUzdTwkn3I3oz39KIs2jgpERDylg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZFnL45FnmHUdFoiPKKUYJCjw1Y52YjemwZG1kuBCt7ebU7/0ut/oV+SwRDRU
HQTJA792bkhDavOPEYC6lwChGpcnSq2f1nAb/Ur1NiJLFpyFlgCIS8HaWsMn
wxGKXn/kcgQwwaFVasMX3NcEu+rssXmXh8zM25yzr9E66k7Iek18MfBihRJn
kEgaaL+2YFXOzxklci4eEYtEcIUL8TL3NAI/BVbKJjthobfWENu4aleFVeIw
uZg+BG+Z00VwNKGLEXtsnL306JgsOYZ2QfTaDxnek/JM92AGuWppB2fIumm8
XkGTbudKTkJa5b2ePOA4shh/JDHmzba6LRsJWtUa5g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RRYns+3Rnje1M6TbgijlsrS3wuvtNIO7132nSYAOp16t/LVqkuLM9CPOu+BB
/+CgB3IV+R3/sFHZwebCt6bXWtm4j8D2DlF73AGeortum3c7RlEcvt+fuYN8
A2EAbYQspHnkHrzXzfATSTSJEB2SHp/2QoSmZudtFWIcCcQgxX9uth68Fv+a
RSmzBjbIEvaB9CmThAC5FCCX9MlZkH02wC4JKFQ1GlkC19ltbTdMiiDaFBkm
HjR4xM7by+inBH3fH+DF6Ol4q11c4Eoxw3ovRbqFb5zOyu+5NChwuKwlk+i4
tqIQPUzuLe6FYQK1RLByL5rDx6XkKaSUrGxrvVFafQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p68bg4JW92Zq6g+JoQMA6bbstF64yWm8gxfFUpDooY87XWE7iMpr5PuaBfTI
wpUw5izfCOPvhMEUB87Hf9JuDjdVFrMRCEvJ2FSEBPyiHXxHo0t//Iu57bBx
b7BcXWgLCezrQKsa/dw5borUraop7k1hQjyca1nkBOKeTMgO+pc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
RCqpe/nKxhhcr/MleK4VEKjcsyX4kqeV1I9Slfqe2qsMfK9i0dtWzWXp60x0
d5d+10jd7eZlaNhlumTpwXxe2v6fVeutjW5Ljt3zV0oqGoUiNC81WmG4jsQL
0OqzvabeAbHq3VevJ9iB1QhK2dElkZhaSGoKQIaxAfx75hcqXEZm6ojXFLsx
QfuTrZPwAS1lTPcoRWbkZNVrjMEjPgpucPGaBf2HX9QUJkFUqzJ5KGwz1bKD
AxXMxSxzJqOgzys90qWVUsVFlY3PTL8wneTf/XdiE7s9pO57jHuww6EhAOrI
D7vx0Xwbkak9kXa2KgyYEkcqQ3piEs1iTs/GZWD6UP8IOBGV9DYIm48tABxb
sk43opOyh3wfRTNvai9aVpJQjdT1uZNxR4/Ubcf9KVURUeWnjZgOKcAAv0ki
lzM1w9wizSAB0ce8avL/ecm7LAUfyF46iF2sadWatk28wc3aAcr6kgPMB4C8
YIw1IMUVu5LFfnfD0kKEgAkNmC+ariYI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tIgFoFKybdi36dScWwROL20JQTbhHhgLyfJjqufTr12FfQb/CpPosIj7e8wh
/Fu/ibpRH66cVXOI/i7bwhgIKoGk11xvQBjaCY4Oj88Qqf25lby0MUpVuav/
VySufs0PC9MJLVdMhDiSpfzJRKMRKoaK+406kwuQalwV/yWObVE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SsKXKrX5NMWYwiMfGPvy74ga0Itdd3rb5bmN3vrQk2lNa3dPvmBEcNwakWZN
+nFp+bzjAcLtIIdenVmbAmTBWdIX8m3VjAId8nmepDy7psDoAc8sgF55hpaj
QbSeVMAbw9+HuIfV9l07ZFYLCzC3wtQvJLa3lgMEhDs2Z2Ve+vk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8784)
`pragma protect data_block
4yo4suyeHCNeeZT4tpTrQTPrTxUy17nzcnr8f+O4g3A7CjAvV6QyJvOYamWD
EgMOSkrL8yIHwTs0YfGXfUocwKCCTNsSlsxzFplT8iAqfN/ik0vMlDxapG6r
hhiWw6zLfkwvEqgaaAhz7z7kHHhfch2FkwJ8CCBl+MWZB7QcCyZ+PHs4frQ0
8cpU9Hz1mE/ZpDwt6KN2rMhkMG/RJj0sdISc2rOoQERjxHvbhwXVwAPRVgp3
O6H4GABd2DYIdkzqS71dvbw+0/YPAS+ZK+eG++bIkTxygJBWT81xU4dsZNY0
nA42xLx1cEo2RZppvtZ/Djq63+kuz1yNf3yMHW7ZF0E0FawYVWlUnJZDqLt9
t7677w8mUkRT/9EY5ikgb36kZ42qE8G0IJoWzEGLb3Tn94OI4S71v13l3rfH
YnhNE5n7pk/aglp016cYAIo5LvbB/+Ne5Bwyo9HdEdoAKxVcP0IOoQ1Tu6Ib
9LUL++sgkb1nGC7hoEXQ3ls8CqtNWyWbPPa8FjibzTdIfi06WxQ1GsWbvV5S
hMXja7s3FH9yLqRSiqA4onQlqlAbnvClb1gbEh1mT3cpHpAFKwwo5gQL+t1L
iOqMAcF1mub+zHElW/XdtUbvq8tLxKnng10SBjExStiY+mA7F+ArG70yQYpZ
MtMZfxgu4sCBIWUI1EIe2en2XyxuRz57b69cVUnFCFZA0Uqr2o1GKJeUt4FU
5N+IKoOnt0PlF/ytDc2AshOJgnnJjtxxYUl8CsyYlLj9nfxTpzX6qc7pWOka
pt12dSjVj5CvJ6djegJRBwH+RXNbUVvzlbxmHEuVFpi+PC768buNHMo3Wqx4
nTdpKHxI41jt1oSPtPRzNHbJiySPA7p5tdyrtMlC5Dx4AFx2ZNr0oJjnNo2m
VB/70RisPplASo0GIFC98Y0F3fBt3UzCHxMDslS9qszYxUpanS0tHfaV8Yn5
qO/fZax6smP7DKSViiVelhBKsDNOmatiJ9AF+XUvz0OQLMGy0tlAoj0JcVkb
N7b9CscANPC01UkBSrS64IMapqE1RbuNXtVoeNkNkpR80muEQQi+LadUxprv
T78NZQz+EMeDjOn4j7Hcmr556D48a5kDjJ5RKRy8W6p5iphmflrdAdBJIQb/
43GxgZmdykce1k27DVUCH+4evA+jPaImyjEyNsBcVR7l+z8GLSNZsP2xk6/j
2Wx+lm9txqK44k/mM+W9keSc3NZpKAnHEI4ddSUkh3Bl9D7t3RyCy7iHdHwl
f4vqJm7blMwaMQOfWz+P69Csoqg6N6XxCk3ieIowzhshtD83JgIqmSztEo8u
PcwgOMjb4/zTEn8vLmOBQj1x3x5Z3IFWqKR9Kwk4iD5mszzWgmf06+SAlXAP
01V05iY9DoLA6C34muBT48XSuabM5ZMPVK+/+C/oTh0fDq5HN3idrE7+8foQ
Hr7wU115ldQe2lSBAILVtzt6EkJyMIuS/XlfwUN2SxwzmFZwVkMLa8fC1yYt
YGwI7StXVThuJOJd3WAEuhGuRsL7F5dwgiIiEexz/2DvG++oq+zfJXl0byAK
3G/pY5LAY4+Mim0cBkHiBDH63EmkiNWYYcDrYDMqQWWQo2SK+Ny458QQPvnI
arOYQQVmtzxDoRm4oUgzOXs2wR700ygTQmTNjt1XqBaWB4h91aGE0cSYRVvB
OijQGcHFeStBWZdXI1uBSLYW1tcUV08ydorQ8f9rrshUnUuskAVZhkHm+New
YSeL9jVleEqNGCH0X9UW/t/5Ux1G1YqodlxXJySP06ijl9xkc+VWldzpHljm
mobuL4xnan3mz1GNDwYB4Kg/EP4nzvrlAWvlHe8FLlMvR0MopmoRk/WHipHc
SrfsXMqPlQ5SIQPS5kg6HMDFRCN2JphS/Ty2S2kgsMIyMBwNG21ISruEvvE+
Ri3gv1Tx5B+roNzdNWsRKNIjCwdqyjoj5lXzrJizj1He4c80fyH5OHl0g1hp
4o47QulnzLtCEBu2fe/cuwQIqM3V/punU5INkaP8DJwCSqBU4nYzZbTgv6n2
UT+1FsqZRKKiwmEeNOoOxJpfGPz99dtFm606aNBFWoHQ4e8lbQLO+SG11ESy
j8hIsnnOfF2o9+4zwyqzEHc9maLJl6uCYxBo3ryhGZKifBfMAmEOBvwWmt70
fsjoIrFPUP3sP3gDo+PKjBvdU6IGZMjG9hzHlBNY358RqIPtJYO9wEl4RH2D
vpWjgMV30+bgWi1axFXWpYswTuDR3lJT9EExsh6mfjU6LJCCzRGph9GmY3mN
gUhM8SMgQs0y63YCvptM8z7p0jDcOUjF4/f2lIEPszVeY25pvfo9yHlCMGMQ
n75PsPtwm4wu1LCJ0Bi6HmG6k1m9SEP5N3TeQl+IY7DhYkx+6AoELl7M2cfv
t5VSFzky1xI5cezCBqm7ztyXcio55XnG9NdzjmpgVPa14/1vEkssNhYw3ebA
oDJ5xrAWRubZ3Qzt2c9nW2VuNKOjX0eJe3fbc3D98KwNQUSck+LZnsvxInQU
AITtjziCnowi/G8ypYJwLJdgnyJ1zdFlqs/Hn02Tc/W6cirSSfvwzIoIpiAR
TwGI8CBqIGkxhyTehOXyLJzHKLVEMQ3dMNqQ33edc4ybco+ykJ7/TDMvxkQE
D/d3kL72VNTgoNQmLGSuN5q1e9kZZ9TiZU0SmUg0ST02kB7LLK1G6LxJZi0x
00BdvPma6HpTBF9nDbWYnWe7oehS0tEmSKnK1WFBfWeW2m8lcUEpEOKfcdQb
6MctkGmsbpHziINpZ7F178em10DEv1mHYGjct448Gk9WMiXpT7DmjTnEmhzD
+qG0IsoKr0KXdtT4DobvWj1K0AAhTvVtQOf2He2I/RC9lfOsqVG6HHR/s++w
aWU2wkdSJF+neatGT6RZ8E3QgTNS2escRUDIrIbTGtvN913cbbEfHK80YYRK
dLjil+Kr4rG7+Gz+t/oCYMkAhQQTVwgm9qk3LdRYvKwIvFXFUPA3l75iJI66
oSGTJGRsHyqu9FiULXRusuJ3sKGs1oOgI9oQZFwWA4krKcQUkig3BGc15TxD
cbeI2nGrL7AraAJD2DbT8nsUjxZnPGskwdPBJ75Nldrk0CSxxDuLzYJYyexq
BRNhDOQq34RwsMlNt787vmzj2UBOjincOihPQIMg85UczP9x4nnp41F6JNMa
ibakLfYyP9h7IKSqjIPi0+kyEra9YThg98Pi3zp6+qZE9FNcRwgMuGPXvMgQ
vkJGno+bgNBPnM4g3X241s6bEs/Mb+qxIZdV1ZzKGm1xAnhsogb7Phr2lVX5
32F35GsUYPEBURrearBEOmQdF2FiNMg46SoyUz3dlFa7bzhWUotaa8NDKHGt
5p3l7lYwtESibPQS7226w0oma2gMzXeD5z3HFG2egUZ1GyAk/ApVFUQaRTZl
t02wu+8OBJJ4DDgArtr+kGqnUHeN19fQs7sFRqy+94fFaP2gZ/tKreDH8oYs
XElYUzipJB7pWUS/0jJqD0zMA5dUF5T+LMD5UaVGzRaYzm0+4PZJ2723CglF
z0FXFZ05n8zRRbbx5E1wppVA90gzubjSfMAeDOZsrCXb6DChm2LGw9wq/MNo
J/xZ2O8lPtcm8S35SqzarkO92/UyDTmoSTmG/v6mR+9tJ/fn/JhmwrbiKJqk
VYMJ16M8fkZdLi1bgNXTX6kvS1sSGaQHf8l+2/a02U1BBMbIyP9tReV8I+Hk
aNdTKqQ5SpYQoXDlA/gi3E+/2dzmBFt/KBNdBcDlP3+r/WbjawKMK86WZGn2
GEKvKJTv27QBUL5teEWg8+3Pmg4rHcJ0L4pq+S559N20R67ex4e5QeukJROR
4a8w2NIAEfsC7xzJAsHDtOePr1qBE7bj9bMZENnQuxpyCcUgoNHV8lNJEg03
9+A2jAO7GFnCaQO5fRVpFsmlxQ24kOihLXg+JcwiWQ10XLlFb1QlgJ/iS3dN
Q50xWCDPqIpKQInfMYzdwwJpOyoZit71Y0hwO72rvJJ3CKb6smWJKQ7TzXL7
cM9hHFCJkJnchF1y4Q7aC8q/7RHCuQEtzvn1Bj+ERmLDJ8v8KSunfoZGmSQR
D1zG7FhS6NF7scm5Ven3EWUzAatVZLswFjZo2PZEoTNVgiGrVOSa3aT7pPfo
hFdigVxdoMZWnfgrVxfFdSt+bNH/SlMkzl1SsdtB1aasiYrGu+2lumoKfuKo
LYFH7AOucMbfuqpmfqQSWrrI+YPcgQMoc4K3A36IXhyagpPB8fYncGr9GEGU
O6c5xSf398uGXFnV5IxpUW5symHFBmk8CXFCMXkSLMAi3BQ9huJ4R5FrxoOK
oC5SyzL3RBJq0DcdQIAN4RVTfLJxw5vlVw6bbIXJIhhQEddg5D35sWDPmp9k
sPNFVatkn9qOKHkJWiwwPut74jNQz5gRrIVul0d0x/1EK+G+Hz3iOpnkbb1A
i7YkNxg3MYPecOehQBv2NBCE+QrFScLiaa836+AxIg0fTiXVrMgHIw5WIJwI
sbIehZ4r6yy2NjOjtDcY8pCSH0ndwOpkHBXfeKwDxTuKBN8a9cpWIqg8f5Ll
4Mvg/JZl4krh+o+LUXESauOvUmrzVkCWew7ZuFT5Tf3jWlugLyDD1OMnXSvl
92Vt/UDpv/OhcjQ8y2Q8nuhVtpkuTb59dv0CRpXIt9dg93VhGLcQp3PbuqU0
70drkC7dmJOoFREfnKAiQPx/50jFhLUQihLpqR70Q9z4Tlhal05VgxK/UGC3
dCsw7ASjiWC+wmZ65elgGQAFbubmeXAlaAn3Qy1N85x8eyH0zlvCZFFY3Pxs
Q38JF/gTq+9NK2kjfx1sEMuU6oOesAoWbg2lraf/ez7J6b8xwcN9LnKvEOV+
7VvVERz5a7/+hpW+Pjcx1LBuwqnbP7mCcm1ib8Ix874zEmQGq5tH1G4jKKJb
e01KawxFvIgHLSIl8SQWIL8iCHZz3iiHgsDcqR1xa3TmnFJEq5/6F5ISkxm2
980lzfpecyc5rj+C5XGPqy/t0dU1taLvavNM1VS0zUoWrdbMOCDoudp19TJi
KZ0Is12uumBKoURAFPlbsEBxzL2t6CyloEbZQPFjWKcp9JTxfvs8j+1HY07l
Eg2gNdrMFYlcd/kam9NYKUG8Z1+Mi40k5LyYL7Ae4oXYU9WnERmJkqn1e2HX
MUuUyjK7vHhiQPndUrE90ldilAwt8XeNkbaLLP/RIxrEINFyZJWS804wKYyj
2o4W//ic+n6ar63DzSq4BycYhvZXpXxtMbzSh0J8UquF2zCY++2idQdl3BPc
TJqbBj9rrgwmOFxqLR1d/vmScxGJ+MwlXKPfRutbkYGuZy61rTESd4KgOb6/
LiCr9yJqrewYHkqLukDdqsdMaoO/mUF3MAw3/WhYK370AiCsq0jIsRoZsLTi
Xn9BcK8h0pPIbf3RLS2EdhYMLSHbrgoQ6hEuliUkfnxkpEkvDW3CVNn72Cub
v6gs62BPgSUsm70pPLvv5xbRld07C93j5g8cPezdAyN364JVnjKL6fn4Vhbs
V3MGuB8bTeWKvyvU7+9lUlSQgF+oRDmd5gLTlqo4oVS08v+TwNQXBeXdVj5s
Rs6wUvkPHpxGF532T9DE5YYkzehwh8PrZC74PHj9oBFSAeoETHWhnS5IZ39P
Csrt3GPMuBAPihxO2HsJZX9pIjmYyWLrduOsFGkMqOD21oK0GfvotqMIJpou
VAa/4k3FjX5kqCFRneixy4MkEZzCmQCzn3l7Pps/qSMypUZfliEnnU7INvwD
Z7Dl4K/ex/YQFUPS+8WMGCHWTyvrFHZsAyeriBBTdxfMapivabNMrwED75Ev
zQb8wVnIuJrrt8tWDy8MpokrIzppl+TH3LuXDuIx+tWCoHmVPlfjyyZ8iD1z
qFl+maLgLOaxYwqxW20aqWoKm78TIVfj032uaz/1M2M0cMDcWiHuGHEMeXIw
+xdACLr1E9OEQ4G/ytsVPQBjdNDtbHWbHtLPhUtgKn3XzaZavlZSYA5IAAaF
Hs6uR+Eip9l8f5CbxDt+i/zy/KhuN/opOnYSWYJEXyFU0NcihPVfbw5qVeiU
Ju0jlKnJZndPOyMgS1VOP6qRbc6uqGiBKUPAHYlIjPrfzvrhOKQMH0QJMfWF
9eSoCfiWPhQp7ZmULHOMT03oTwiDqvsrgUMJupS5QgmqosCMoIHBNJMAuZVj
w/qkXYySsiOPJK6hkdlMLtDI1MzVjsouVkrYmZozrxbRffUVeglC1Ro1QCYW
qPiJtt8eoaJqbWyx/SlCFFbyGJQFQdn2T0aBOh5Y+MYHT6NyqepQTjhk7EYG
pZyCDNALCBtWTkCEusvFmex7sB9dNO7NVUOQNWGv5EKVmnx6uQw6c8573Ffw
TKLkz4gUKc/IeDCvJMx0Gk+ZS++tGOroN3Mv0vDlP0Smf2Cypebjq3SVFy2z
tN4pXT/oih03MoyjsnGwX6WVelkZ/i3pX/ao4sJBNU9e/NKAfEOjaJ1+FwY6
9hdB7LoBl3jaJI98Xc4rvMk3B30YqnjNDNmw0iz3a7AModZp7lQ69Qb3KyWs
oF6SpxC+gvf8eBIiUrXUIV0WDoCGY43VVwrrVtu6CXStPNHwPspnDU8vLnaI
Cn1y0LE8TOMi7xgX/D3hOs52Gyi7oNJoBcb8n0ubGAEdHSvXJBkm1OUjN1i/
BEyted0OMy45zpLY8/g+nX/XXy9a2Kiehh88StHYTlZBGNP4JEOYKQKM8dH6
JrVVs4nWCiqkk3qfqIZ3giI8kDSfOwTGCO+CfNLigLRclquqRURnIVJdaqha
z8Txdoadc6Kp52ds4/thDFaq1qd29cD9GVTL4FcxgaS9DBZq3X+jnjAFAp/o
Gzzpo012uzTMO8BLX9iPRTFKPgxclualLY/EeYSFGvvd0QNVSP2ikMqchxFq
D0yEsIYQw+JR3I0WGn9ZbfQl4uFj6DR0Fv3pTg27W4QeXyKeQOIovH7y/LoY
tCBA5mw3EQSPxz/r9fGBklgygiK645H9pNhiHMsWHjBCRiw023DcoYcKfuv6
KLkHWT9nDi8jq+TAA80hr+5jZ7p9sqjDXNaVocH4ulZzS7irwNJoTun5+XM8
/neEEGnBO5qw2uznllb3xxHATIWn5h6quwhFB9bZMgEuSagqc5byJw6VsW7Z
KY1mf5HZ/gslsViwpidpPkG4JHfjCnm7D7y7EBDFjmT/JyWrdYkdamg1W3kB
uVotjg3qp5u3zl7htW6tiO3X76JSrApex0ppYnos6HNESflQFEvDUofxWmR8
QLrCqOzXmQDPJBuCzSHGXu4sOn+QifsUm5VfJD8E86X+t+3bsosLpJLUEcZV
guQf2i21lKfqngYm0Rl0UTSuKeXVq3cdvsCm6u7tptSF2Ex+fYJa5CFcnwu0
z+oGvMUY1JHAdHY8hlmOOFALtYwW8yUwzt15FTfL5Bmwn27G5xrdEXkrypQq
gU/bUXYjuddFuNqvTjcxCKWdGWltdmg92jY3wb5ez7GPzQuIrmyOfaN9O4Xu
dREbTXY4VK9gVvKHgcOmRNpV5DB57MoXLXK90lTkuWjb4hjOKQcWyhtmVin2
RxeBCss2kiWvvjxFeAxr5DIybY4o6A25vOqGMqAVftRa5AP9SyE0MD1eBG9M
FFlG1BNihsM0RP+V/m8RQPN02tke1RNamuIE3D3mygEQsV6Orq2L7cq7dKPu
kdaM+c9VZiSSM2ein5dUSB6iwJ5honI73R59YrPyZ0/BXZNT3hRPmC9/bXM+
oJodWcC6eT6vGqC55yamuWqtOsHENh0BFwGmqLLgBkYjU6XhzY6ewn0nPZgJ
55tKwkl5wtCRxUS4MsJ50rVW/zPGEikqWDtFCZWTjKxINPYfe//bwd0epz/b
fcT4sJfPJDRiSj3XuYM2kYW9DvV5u1Msf0U9xMIIpq9z/Qz7Boscj3gaqXny
YPZ9tboiWPkdCKAngbYV+Uun1UB7oWtXbUme+vlNcAcyE+R15aPgtBHbrkul
lLsMKIwulDI6QupWExoBB7srl348H2FvKh4vbYoHE2zDEmLzBoluKc/Pz2oB
ENbmXH69nVmYfSobCiv9vBRkHTzJHvSt9Fgu9YOjGTwxfvG2Mtr5vgYsdLN1
OxGysi1ZsoEX3+0/Cp8AbkJUZpLWnNvTq/1PKbHKZZEjnNHX1GK4jg9QNWNy
fo3aOhxDPd3YhDHttqjBQT03L2VLJU/mlfxF4ga2bdbYdIQSRpkCYcm4ZDdG
RMAghTQNmLib4CYGXi2GcnLjqksOQA4avf6ARbAT3lwsAbITwkM+8LDzDP3E
e2rbwV97oQ7g/75dga1Z/Yzm3AQ5v8Muk+Tc3fli5r36H9XrcilYiAeLSvYN
BiSu/pF/ewA4R520nBqNFP4aMuudVI8aE9CTkl1GOccJnBhShydtuURfgflT
vE9lCYFBfcQ+yn9mFyhkMpZ6AgfpYCW9rMzjhYGyhQ1PQq+lwObJ+El6P2ZX
20cigoMFF9gaf05laFzZ7rAgJrnRUtyyeeiYVvEu+hJ5LEgOESWEMhVraQxV
EXwktD+jA4i9WrpyKyoyeKCc2pB7b0oC++Xg5QRl6rpTYuDCIlgvTo3sMnUg
FhG+Oyj9imbjbhLzhYYKJOqLzHkAzLkh3sYyT0zEvxzfQ6hVc1hd3yVThBle
An22A3rMZQTkfyl+WYQnWj5WmYG8tUCNhC44uXrCDKabp39ZEqzx0ZYm81dq
JwklsbnPxD2dm/UZT0YniAqjdX4NorlBKUOUB1gYzX6xialFxjdOVMUf7oWu
Hri8nAdNKmMTO9JuJhm4lzUWLnFoe91gEidGMap1MRPrFZkSyaVwuTkzjz9h
vrnehm8/3DX5kfJ8DBalLmez0bIJpWHhjultPZziDi1a8zExq9gLtHiQDZps
LjcU3lOcRdcBd4t1OxcTJpdRL4jQfvRE/Yu+7czw/NiXsjYAh6okqsrmDzmg
Bxu6zU6vxhgMoe3nk60V0ad4/38USonG6BUUb9nVcYX35gzmc3swhfyCl7RF
FCQiYcOb81IQnycADBhjxKJi34nTOtiIsyT6fqH/fVnL6NYoPDBlEyhMibjo
rPLMxiv9jyWVu5a5YkAV8acwNp11/4lR3+LFFFhxD25Z2rDH8J4fbZCU8Arl
F6OLtStUiZR0Ks1AB/Br/le1WVaG3FKIiroFnEvKXiCwCwBzucNhtejnvWpt
D3StBI2s7RTBLa6biRuxdpBPVWDHcVNvxS1W/k/4zNRYcVq3Mm6ndo3s+8En
1NIsvBtDqTJ/FvnOLvQWNOzivkl/9GsjJw7JhD5PU732cCHa4a0UuCOHpHoR
lxceWvK8yPsp4iYounnF+oLNboG2sKamJtKgjdOY/JRkgFPp/wFScQZF84mK
w3Oa8ynFrV41F+W5ABDOugG/zOuz0QAukqb6BxTvDu5zre8jqxSLvoVgRUpn
Vp5uUX/tXFXGkVL5Q+bxUZMzLkEPbt84KYiLMmpGgjPHPECSE1ZoTSiWq385
QGeQekIlDKNpt0jCIGBOZOKKZAFJmsTR6PGONQZjfUNVSs+JGJR9Ht3ZVGUR
JsIfahjotaVj262fotLc72Gfd8kvDYEShhssWl9aPom1uXv0BB/hwFoSn6Gw
BC2p0iHm3pM/dAGhrXDaJEQA+g1g/9fSM/O31auXH+1OGV+KunaDUnfv100O
5BfKvOKTdJLDrYgfooUMDr/kYWlrYetzwnMVnvVR7+tN6hT4r62cfxnm3ZNl
YXyCv2ldTuDDl5LnSaaJCZTNuHioZKkWboep/4lUdMxxB3rZ9uAV/Q5qrQ5o
RUB7bcnKE/fwK2W03aPirejQ89UgS8WSbPKp0nB9qvYKDuD26WfeYEiHx2j0
eAHZZWkScGSin6NJaz01JfrrXPnMvllVRfb/staHmgH995y15H6qP534CkW5
sJecqv02OVzxprBYV+n4joPOpz8btwBGQ6JE+4BGMZ5voV6DuVFEdpUeeSNu
878k7ihvbxjodR+VYWfvVvcfoMmKbhionfOEvHYOgs0H+JkphcA4RS9rooOn
wTGekNuX/zFBSJyRACHZFFrOIv7yWbYrQ+W7R5kHYbjD7F3GptIT1g7AkH/L
l4xMqDBuIAZ88vbt1aUJ9rzklmhb+4icmxUeEngOJV8IS45tDKihK0b1qmmg
Fm840Kj/6vMyW/DGUePRZ+w84RKKNN9SNeO24Rwnt/mwGtehVEr8XX8xfYrV
/vSf70x6d2IGF0oA0I1mvefl0AE9imhFmGatfkg2agGFJZrms1Qubyd5addW
RKGcnFw3mlZCXCb0gJb4NB5NFsndlx8LfHYVMmjsA75ZjIwGtV3CvgPVC+DP
+lecXPnseX+frEq6iLS6sQMvpT6qW6SZZ8KZuU+T5ruxHfcec6mMu3CF98Ab
qq/RZ2vlzP24BeCpH56mZFhzoBoMQU8b591lxnIUr+EVcaYcs+QGKOy6Uym5
cBuXleoPL+NwWEq6MTWYopB7usep1Uh7A4LjXNSGvePKva3cnF2Ue4r0jX32
jCNp57OV5OW12M7qtidjjQWi+L5tLM6Uk5KcWo6YE+LWqLRutqu5gZ+chXrx
sLvFqY6viAoiEgACZ4KvKZUc+JTlOBaBQVk6F14orJgnEgdzLF8bwwBkUEIJ
EWYIGBcAWmIO2VSfJlTywU0nTSfCXutbyMr7x75ydWCirlmXE/KaEe8B6/CW
eDHpL0zEoOI7FTR9Pg08JUycULR7TYpe8woZs0gpisMttkKVjhvRnvIrcoHG
5ikaTsw6g2sCiAUe/rHz/FhEHp9jhKA9raEw1I82kvBzAcpS7tPAiweYmri+
Xe86Fr5K94KBIMbh27RwnPJE5tJIY2rTwopyhBhy1M7bHNY06tpx0FhaXMkW
TvZbH7a2ooJB7jvPmO2rjV+6ZlC/TN+jQf6zSPzfmp9rsen/jMQ4QKMcXasP
p8KGR2snOgFpGRdcKifpcKKNZJMcosSeOFzinDax+qjuGdmpbij2M2Nq2n3W
CtvsbKZzYDxOy6WyIWQyNQHFLhmlzhK5QgwCio9D33QGAlGHM6lpo2PUlIxq
1qPoVNIYiVQGTUssBT7RgHypYRuEcpEkFd/ZJMWpk5xFIUntmnlVupj07ZxA
MJlJoN1QiL0VPtIHmC7sn8HiPwgNVjYo/ICryFGa8v7DSeZbSQJuLx6PHjgb
97yciaaBYwrW2bZMqo/HP0vB6uC6YnYJcVj2NC04DL9eEC28GsuVRPPHpYQ+
KChzIcPu6So8MhDaTn3I9xr29/MVyVo2dofB8RKnLemfg5TDtfhSpYLpLpLG
dFtJH0+6buTsVRiCNLcyWIaMuKUCNsmMOCQTK+9Jas2ThV1eIz1U5M33Q2pp
CVFsTFJXNI9jHuw+q2wI3jW4uKQoJJpnW8HUTC2rvHevx49VjFvaGVdTVlvN
ZrpGwndaSX93YQFq7UxARELnJtWRvFlkc8mk+cCjLtvS9sFLWogQY7pnHaiB
cQJ4W6YbTt5rOVc0GeGQVu7UbjhQcR3SLGJVItFwv1W1iRMeuqgYp2BaHNao
IaWpknlNCSiJaL7qpiMdXdMZLp18DrLWfAr67awIWyNtXIpvPuFha7ljH8nN
hBrQzHhzgEMA/nkug8Hfqbrsa57A9UN8WvxUoh6LciohKvBtFfVflngPPWB2
YgqYNZuGQ9YvSDi3jSyRC+6OuFpPkMjrv82Dx5hcWpHVnhxsGi2UO6s3NJ/6
Nq68ope0v1Tu

`pragma protect end_protected
