// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xEqnDHApM3/KiFWMsKBHoHswWZQ53byGSydbJgto6T8faGRiPeqVHJZzMT9N
+7DjXBlE7xtuGC7h9/56JHA6Q4Kr5VS2WoL3At27r9McqegDiTxDPZYxOdHm
cfrF/s2wrC/Mk3fXmk9fdzq6dMnVCgmrYmL09KtIz/LULsK6TIyWSc81oNRw
Al7PZJNLkEaY6V8xvN5xSrNnNEWJOXewEEzRCLF4TLE15Jn16tclPWOOgFpp
3Fd0EyItq3b5C4WTDDdKDVOgZF34UZMQNtg/G0BBf66FEz8UhXneBdwC9SEh
jltZ4Wgz0+or0BRp/koqZDPxJttsn44IqxdNwfUfhA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m2gUzBffi+t8wH4lTe7we0NtwhpRX1rtMui84CHqrOcEzjUqH7OLcoB2yEZa
7VIUA44kfd2ri7wBePqla+DDmaAfLKXwwuWCrwt0eWmZbFP/r6LGRL1Wvp6P
E/jhjV0VMaPY54N8qkcr7KmpWi2jtvI9+8pZrSgN/zpLH2R8pPe3EOKbvZEN
mOQSec92FW7PSbqaW73cAE8rIfjm+d+eT1j4SIAS+z06GCeEzF6tT2BaLvQx
W7FX7bij732R6WhMH2S97VTDquRFTQwYGCJtHhhx7VYjyhGGzsLFCsltfvfo
DRTvK5+rkJkGl66q0r7ZjtUP3D3R8kKykLURCDJCDw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BaVdnJxgPzTSOaROqid54Oh9bWghA47etCTNloUn1ggcgrJoUOI8bP1M6ya4
Oa5Bta2i2SwF+kslLGxtvBN9BiXxpX9WGkiNfSXt+vXt/hz6Sb+QWVWcv7//
DKHKQZjJ2f3oGH3Y3Gzrs/y4WqHWsh6hXUVSNOS6HLgyeCV3uuOba4BLzw3H
gQHVv/Ksh5dvyMjHHzY0x9/yVUvnvYe7FzpO4y1F397JC9xGBQAGM5LVgj6a
JslDlbeMZjtenQ/6h5QsH6w/XiA9uTXxVG1+OTRVgpGeNKo3vAM2cmxhUzUr
03hSIdbCmneO9T67438jyCIvy+kwM7DkrO/eLYPd8A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D9gn7eu1i+KjodQPtc6s2osbwk6KAlHEbdi7XJ71ydpC+b+IZrZ7BhanGQTw
m0i67cwUk9wU/b6bk2m5x2dK5ElLHHF7HQtuna6+v2jvNw2oF+YLvkAuc56f
ye32XcPs4y2feEx5oRQyMrEXTftksQNWOzVpwrJyo2I5QlbaBM8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AcSIvsJvIl1YAdQd63QZmhS1r8nFP/+xaHbHx6qJYze/acU3qDkVZq0ktYAS
vF93imcrsWQpqlWAtBfy+I5/TzAZPb2S5XVDvloUtfJFgl6iSkcp0op1/EWI
fZEH6UNKvjILp2IlskiaVRvPgi6rkort6kNvpsai9Eg+yhIxvHYSTZRqZ1tv
A7bSj5aaTXdDRnpqXPQxjk3h3sHytwJJv+ZwuxISxIxK1P+E0v3d0Obr2lch
+QQSLvsqAuFvLTKnf5XwVxbvTkuP3iI1aKN9bRlmARYcEVv7vptFZ/uI+s5w
1ZvtfN5AZv97XX3nTg8YLJPIajiGXNOmNZ/k9yZ/VsIGoBA84jOuOOoB8K1F
Q804sT463F5rz7aSihj/nbV8kph6ck2TqAkY+EMs7zkaY/Egd3vNN2xGiden
vFqih0PIgJsoUimwJhgUyqvQVVTVvoTSTb35fSo4GS1eS+ImZaEQKDZRRwUo
4MWAsqRUHpgN5o7P23fgi1PSIXFL4OzT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
M3iJ8vrO6XFqSrx08pBulgP9kC7+cPrX85pGr0YBQd57Q1JnEk2jzNp6QSLH
kbacSjE8vXRwCTr8ho0NySZWPorXmiZUBcMiajSVz0aKht6ZpD3PLMHmvLm8
rUN604LQO/lx4Uy1WLeo3BdDzz4EysBGSJ6r8A+Sayn3tzhCVgE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DTpy0+TXTgUihlqIYx31stcT0tTo1FqtW0yn8u0d4vUsKvkcNlm2JPt9Nocs
v2TMl5+UPHHfPkIGoobGytfFFQ09ItjPAxbccmnR6kRLJ0Z8ROb4nyaAOu9m
eHrXL8x7gMweJRn1DXUkOL0z6OP8n6YT2upZH9gyBvkkCZ44dlU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 144800)
`pragma protect data_block
z6xySlpL9o+UpM0jxiSLZSKAN9FwlCkCPY9U/ujXHmBbZ8yyHkmhAwOeY72i
Urbm69uxkZg+xc6SuGFnaHH4sUwZcAJIXsvmaq/WfITeBIOXHLK3aD/aoiyj
ITO34h/ylfRdmud9Spw9NlGC43wT4SXmYznyizruiJi5P6hqBeKltXbNDdJX
KWiO+GLXiaIlYLf5dZVasPwmfN62N3RzTvRcX3r/FuIjYhOwVAK5wuFndtBk
zqjZ1sKkrzhz+xGjqhX+D8DX2OM9dbHw0k554oDOtCj2dE8YrrYWYQ08+br9
YZd3NfQKf9iTl/tYJAbILNStR4vbl3qaymFf2p1OQtsZhV8GAMADgX9AxSbb
7YLKWbUBouRJWWOCqu+71blD8bLpZ4LtMB69AcSplzPPUyjjVeH2LCJaYUxe
zlxQcERcfNVlKDhuUlfSiLFK+ijmS3CCcSF97JIbdRPRx6E6dPRba8X96Szr
RmO1Vy+GjgbWgkmKJXzOV1wP25oXtWl2jgssMBmsQKYmAd9+//EOM0G5NVlG
9Wl/XGW6oU/9bxs6nscYtEZ5ROu19XjFda/PXTVb1J4Ju5u05y6R/7OXa2l/
+4dG/fKDGhKyQda1+OAmC+4x2gAbW92d9TIvX5BMAzAmBRJ08wiXbeKMJ3D0
e51WHGYEx8mSkqmJc5b/Jhq3gryA94szjNuo64sCJERRY4ZB1T2G89pTHV3d
s4sbwlEpoUkI3t3UHRCzwy0+cCwyAj2C2IcButPusyY9rCxJ1oqxr4KmAFO4
+cGFrTgRjb0dW7umrB2vVWuD+yy15JdZ2Om/1A2woDvOwXWSFd3Qn1HC050l
onl05mj2SyFulRAkZMwPtpDmvnxm49AjOQwND7Ot4CoKzkNvVBNWARCN/9SG
MqnUW6J3X6kQ3QmmVzI5VTTBHDoldUgs3pvdWVHLFYLOFJTlJ5+pkHfSlfgQ
N0DOjtbJZOFUvY3OhiQKCjXgS1S/D0HVz5GG9fkr1KWdpy1o3BlRuH+R92oo
XWXancVi9vzGRG27Sa3ZEic+sCkgxlgNI2DRathbMG1CIJAf9lwMzz5GtehM
D7xdrznRVKQNxxSZ84QzVGzjqTZ9ULL1JWvfyWlnR8KQhU8uq/pQYmcACygF
VNKHSnpfTtBehB3h51wTkeUijCjEVHXmYMTrzmOCTbOe8XSUnp2pZ8NBQTI6
ldg8ROdN3l8cVT+hfOFJERO+6AzJiDk1rG2hS38oX8VpskO7n/RpVJkKgbtS
FAcDpMGdB03a55uLxefxDA2kRNGdtHBBBNnwrVncKhX5sEDPzbxO6Mu9Ql0u
pcHocQP78eZoMS0yukXY56YMx3Be6Wgv12GS1UtBhSgX4BHieu6Njt6Jjr3r
4swPiwis8Ype/sSl0WiItNFMYGsifdFb95bV0MihHCzbW78fXr+2Gypz2k0L
7ugbsH81/5dt/hR8krmTBUSLhwg4M1xlgaswKeBV6Bm3jBiMa3SpAKi3LdT+
zRIV0d5zbI94JJOxpLNc9w1fh0EeSkHh9pNnENppuLcxq3Q+uSpAC9EUEg6w
IFLgDbHG4cjiqmbElw9IOmqDlxs8Ssb8v8gwfgzRrxC+YbfXvBcVzzvlEGxF
KjWa6HocS/grQ8KoRZ2CPpDwY8eRHeObe8xbEzmgTWJssVLU3MHr8D8YQrJP
v9ICyeQ35zT3rxo2906g1CEaYOnWgZPVvl5Fx/vLuvzK4A9BkUM18MLkGx8i
vKc0NOaa5t9OJ2bqI/jfRCchZBSJ5Ul0i1DFQDjVNLg51ixtz22uIBh8OWmO
aEKZYVmZyz+laPkXZU9gl7HYJq0LSVPj28Y+ZCaGsbvnxZHSnRDWceeoF0rM
YxlpHbxxhmLkPMqrYqrOpQT2O0uF8mF++drz+J/BbmRjny/n4WGHTBd8WVtG
uNLI/zek4UyKmDjCWzSGn108fXJZVw6rqSWG7BsI3hXIr4u+pWSm2t2SfEOj
HiFORLlcLsUQtFKCJwMYDTO7hIzi6RYkeDp57SemN4AQRt6lbPOvNhs0eWuG
+2PZVw3ewBvmOTbjYzAhdIblZ3U9Ih9skdbD/TkkE5MmB8pYeqqIzuksrrd2
/8Y5aiZr3jWDthr/E+KLOi6+6/AUKUm1ojhTJOxrgj9ZpzvV/D3pwUfghbhf
7GfPkFBfNkE1tY5IFP+Hnp7CwJrthqdai3ABS+Cvzm/d2PnmKCGVyRWUJBsa
kiqdixHsu/YTmJDWXfRIzOD1BHNpDBXyuffL26YQRiCdizzEbAzk3gug+KEY
NWXmDs2cT/L/vpOB2ly0QP2vdkSBYv8oyOBvsaCSNT0KP2RUIop3wLAdjfAQ
To8IiC86VhZBIYYTFaG3YsaOmbc/Eqk560gHzsn3qMgK5g8kh5xWlaC/V/yQ
3vtE1aMScmQHUxnsSmq3Vdg3wTGgdoqRCHhhcPOummXwBJSqtq0Dr3M4KHvt
JHyr4mj0d5t8kceL5/i8hJU1v4QkDqFzNE9Tc7kkzu6U4k2tvImxgDUJatPe
CwG9MY8Z4mOu8ahYnyhMPNiV93PLsV1a8xtyHVCCgqI1GPJArtayBMZSP+w6
I5nwKkSUGtgD9cAhJvHmWFQhDZVsSsgQOf3h59R+La8txwmdy+cZTndz5K1L
17m57LrSuz8v+0wT2v9L/egnx0tMGAOAIwgt4cTrehoTcPCWk/WgEoKvbbJl
6aTjJ/NKgM802i6OQl8t7hcmbknv37P9Iq6/a2aBJN7mzPO5FTGUWlhDMaMK
hrDiHK2KMIdV/8S4z9xKxHRWEUjM3NgQePw+Kl/KirOyPHyge+Je3FcFtMg9
F0ZiA8dKnRdjOMK+x//mgBT0bzZ66gDgYVjjKCgxTLxU0TDGpmHC2Lmu6Cye
Eq4trJT5nCFPBbZmJhdsFu2YOtWljPv5OnFM/M+SDHnxQLPvcPRRv+g8dTy0
x04NRDSCzB933hqrVTTHl2uGkF9arqQ2uTiROEINXXc8+ksaW++mqAcZtFiR
XDJ/tOBPQoLFpfqSlUmFCMVmdVjeBJ0knWRsdYK6mHGwYehRGmqbTOnIyc9e
5PTa+VwdvJhPzcx01KlyiUwREm2OjkHuMhVUUqXmKQRiihzgP/yHjQPgjzj6
NtnwbWNH59qtM1cqGx0u/iUMutu9/BQNYDXmmeuvtN4paYkF/xu0FGdtfqvT
9bOMLKVIvzvIkMFqoAbv8gM8u8ymt2Q5cMVXQcZBr/wsZlA2lJyxkIZ/jtmp
lXA3+c0LBlnLtAkDgeh0nQJOpvK9gpKwkwZ70h4S6VOxdNpndJuVTR4UFPJO
c8V7CsS+buTa2oFcvvglsuMSdeU4n3ASNZHcsvlee8vkqZ79b3NrfmqFiVQR
QpvM9P3KYl5FFRWyT8+QpGdUjqSc2ezPaMAf/UUdo3OwcSI4RZ2shlVicSI1
o3sX6bCTclM6V12K3sDysLtkUWzfUm7d+9UZ9qyqYUDc7+70lEoS15/rr9kR
te2DmxM/iyaNySoYG7Y7kpANxJZ4ftejlqz69j4DWrQE4Z57+ciE7IKbP/5b
T5BEKqK2rECXi5iHNZfsIv6naYmNoQ1BUX7dXI08DVy9Ub1EFs0KNEgtyTp3
/8WMlUFj+Sj49vxdcFuAAjxZh0qejKf67VI7iqnPESuyZxuNFI3j0sgo6CcA
KVXvBl96fVOk/nVfBjGakgHLOxgFQhFvFn8PVBDN40xHSIpz+hk3KAt6IuU+
C4vt46NGEVyXsY4pfg5gqStaxNktsY41IjafMtIxZTh68L7n5SVMaUWXnj/c
yKorbhygMqgSBIYS+F/aN4avRicjRvk+Bqx9nY2QR5kYwMWbYstBxqwoP5s9
MSt1ZN1hr/vV/adyJpl9Y0BxbxFyZnuYCL17tQX/pARdiSxhWCxfJEMfigYu
I5JOT5JQ9CBoVEMs+fDfB/anTb+KV0v+DgJB6/YY1e5ycY5TyyimFhr6vhxR
R4DbJubtFVHVRRVDSVW6fWdh3B5Auv3nZmjQOI7ynOS92DdXeL5KWobmxnfB
O41ye81hMrfAhq5xEtTki7+2iWu9N+LAXpFns8LiDiww20GaOgNz4JSeIIa8
CrDm1G8L3DMOfqti9zaAVupClHsVYOFMnJatOpXLLY8BiXVCPU1p/955wleG
0a0/HmwJWmnTxXBNWta59hJf6OHtjX9Zk2fqUaKXaHe2G4VFjkmgDFSHSKnV
5p0d7V+p11uv1vigxVv965GgMjxf545EFwGuRKk+7YH3yxXPqRckYbXj32RX
DHDAn+m8dl09TpJKScwDbsUlUzGoAgCs43tC8f9F6agSrK5OXB0b/ZnlJ7l1
S+tp8uHRQP12yeiPXSX4l8oe7ZaEatQt8qHkn4P5PBwm3ZZvhWGc9IGMOBjp
MBVNEvn4C0cPS97KzECogUh2yU4Zzb3X86cCt8CyyNCx585EBp9XcVUtksle
L/3TjXT+Qx+bdCU20fG0jaJrzXcevGtwKzFf7W0R08lWNmMPsX/sw2ptjQlI
MvlwdCA4oa2ITMCO/FUk7dZ6fVMOzxunsfAXbFRhAFFRyab49wLzIeGL3SU7
vsSYk/vF859wt9dumFIziMpTy5n4Km5k/wzR3pvplUzooe4BaOrw/fKEGYMv
oeeh62nDNOVUpD+2oTha4qzUVwE+nJTuhY5w7sb3aB/SbXSA0EqRa+61GZ9c
krW4RH4UANyDBOa0jWdZLWyIbuQ5HVmMK93JJYUJj9Vq16+PtSIPS/OCJXIa
oIoNzNAAjBf6vhgO2gGYexapN8meQa0Mxm0oom2klHnTadKvchwr/ArrBpf5
six5XamV3C1iW1jzKGA/qpSMY7t4G3R1FIOYkojTJQJEnYy8Yrf2et0sQv2M
wc7X3izAKCFKYqCr1kyJQH0QsbeDnYsVjw0vc9xBc0W8P4Fz+PhubaiPICYS
hoLrCPf0ZKgUkiCDoR1mnvXC75/L4N54H24+ho6vgj2jydTG7Gyjpr8cJO0g
0SKXOWFnUvof1VQncgVrsAZfTTnwZN5jjPW2Zwv6BtAZ2Ryc1nZ3M0qoujZl
GcsxssALdSkL5ySOi0c6UwfFAjxuxi0BLGIMVW1Z/1Oh3OHgCWH7fnIad7GZ
Y9146SPuFjjKA2nnlNpnkZUi2cAVagp+5urQ7k+UDAzqQ/kdPjFEqLyVwj9G
PRWq3qaSQI5Cn3Dtlv4letsCAffEXjrnv/BykvIbEzC6bVfsp/xHuutY6kQf
F3iYAot6vS/Gbhb60E7zxa5lMz0vGAwzpIffH6hMPpojhiqYmCTVs/yujOlB
1bfceFODA26aTNe7u2t8wcK2hTrt+1IIdkZTvVKgOECKpmJBHez62MvCct0q
j2x858vbufO8IwmSTr2yNyb+C3a2A/WVCpVGXl1d7al43fJ7EdFPqlZR9L5y
1+CD3ts5RlTexCviOqmWueGhs/ib571KvxIY3ozKrx2JEKmNBVSMIKWWKoT2
BEmW4g8x7CwCdaW6ouEkRBkgLixHk2fUdUr4emGzO23w7hYMggwfjpPjHoDS
S1Tp0prbIbt1NLfX3RcJTXx6H07+sUbbuY1PwM4vspTcshdAxa97vlgE0Rc6
eXthKKrHvrL1a1+eKBmy2nElsQupQiAdpSU0lNT42NX7SFYxn1CGFztFSLcw
xUruzKFBMVs6sNThUfF6CLKdjRhMtEiWe1delENZShJ5ny2ZsPST9Rd8aEw0
lyPMGEzQvYCLk3sSWmRX5K5BzrHmUNJr4VeDwK7mJI17sJZR7iCAelvXOr+K
ZVlN0MkZvUSVfma4h30AUIAqLgm0PWamXOqNC3XkrFG/hESidHYlQfjDzOoC
cNnkVKcF2DrkbX1ERK4f+8SaHI8goxQvZzvidVNv8i13dTXqX1tQCmp50wqb
UmCTWseyuZ+Qetg9v7vFSkXLgxYRz9VZuUM9chSQo4LxArydR8XN4OjI9jY9
01XohCK88dGCgWwpcr3pQJ8TidPJyEYy5tBdYmmQmCrO4ZlxI0ZcYLQt3Vsa
3Yp+VgQn5sUPYuanCEP8m5w5NtLTT+1/f9jdmW2LHbJsjjcr8dB5ksP26mDQ
tnyhThYOh7tgJsM08PSS1TVovn6JtuEX08zga2rXp1Cp454EWFmZvhy6nv8s
AKUID3nGzXQEYu1PCspN0b6r0IsYU/t9hDtiEv+p1HVMKoX1oYY7T7elmIxn
O5ku1AWa1fiqBGPeKZ4QzL3uXeKNOBNkkj6R9JwMYqxSe7rwIBj/cQe8Eg9S
W+c+rwU0pHlz4fKdNdegB53Y+ErYFtxxr8xSGOEEAWJfPXZ5x4F8eIEr4YcC
bXQ5MBkVQ+I4X0zAyTkqNq9HKlK9YCJ7s9z8zPRSwHn90Dt59rnmyXfbcg2U
kzvGvLV7Ks5+L/or0iiXmnfAZKKuPfEJsIoyWJw692djBAf3hltsLTnashYH
8VmWFh2kMWyWPcs5ge+CgoNTULJO3E2gNixkHw26T4OA8zc9qtYAGNxQ1/2+
J/dlL7sdR+mwM+11m+RHicfxjZjy1SfG8PDDln3WN5bLGoFEg03gVJiLPoxb
qEWmQybWK2MKA+BgNIQe8X+qKIPEbjQGA1Gz4PNorcaBRpp2uq2WxBBaCgXw
zEkFSAVSyUDBEX9jt9BQPxgXh1R2qiS6q5WnG7iP1Sp0MgO2szPq6OK2dtrA
A0y+yEbCSdoS763x1onZ5nq+XFR+Jl/rEmSBbN3Ur+syh+zI6LqPsMLcKTv+
kJHiqem/WvKH2mvtNpoR8v1D/wRKPPZCcFsmoElLpL7GGat3B47RIOyuQOkz
wzb1eY3XneLdQA2kft0NeFc/ZfQ3oHmLdkRUzbciQLR7Qvhgna7Qn7jAcoyy
a7ckdwSGFPNZisZTUElxoxAqW0980zottlKmAI1stE9+LKvTHxwbAAmvvMWr
2RgTF+8lkeEidnusn9dsYYGciQ9VdHf++NWXInpyjv5FDmfRRadBK4FUM+cn
+t9f3VNGScSRSHiRv37j76L12EucFFl4gcIcty/QKJiMqZ/K6NNuhdgVpf0z
ze390HHSmrSkmaha34iXdN+VdVlb5GPMVaaQGcHjk7kEJIto2i6HfNM3ho6Y
4t4Vmr3saFPSry/X1zf4Oh0SLBM5QPSg2m7qoCQeoJAoYlmEb0lVSJi+OORF
y3cQELTcL/NWTJuncaddCe6EZZM2/JZ9H+VmbOOLYnr+x3hnaIuIJE/F1SxO
ehfvLnXZjL/87ul+W1Ecl9E12tJ6ewhWV9RqeZUmXpfGfDMxcB9e+m9dKcC5
g/PTRr+nZOy+nOa7ECodQesn3r3PPZ6M/XnmfMrWt2EG6LkfhDlxiSgOSLtr
A0eyI8PRdE21XxnjU89vBOCykJaHg/I5yOE1K1IQjiH17dew8VQnPtBHs+PI
CItZtaL9jTQvpvLeo6M3cbduyeBs4QJFPilETiRnWIF7NYpEXApufd9SGSxO
Xdv+JHZR+NVZWt5Ll8IJDbKMn+j4UybrDWtCoq+t692FBzJFiHGWYw5GBObp
yZfHCw7ZDNn/IuYvMVQT8F5BBcKSlAmNQE2i7Br8he9HZJ6JfAIHBHtqq4zN
JiX3VCY6/QzZMtQVnhbCeNnB2K0vqK6MvZF06XWMRRuN0Wji1VImKM5qOpTh
6fab/kCRa/jINixSoJ8KtK+wzquzgGQX6SwCBmFiMFMdx5EVMhgY1z1KKhtF
LXp3ge/X+SQi7jYqVC5hd23BY39g46gr79rWROrcZxNUyJ8OgEII7eFgckXX
1dgF58iOoaOuwPWG4iTUxcHAPMBwx2q2uf3LOcxDLqKOC+69DST9iggeLT1J
43OUWArFK7ezVxkGwDwUt4XBss9lpltutfLyNolGBX+7p9f1U83mONDkh6/c
qosVXwzFeltKprAG2F9QwNuWq1Vx26OZBZUoxFTUDtUHBOW4bmAiw5rPetIb
SqxCD06yOryIRP2hMDwHCDSnthR6tI2ogsy3XB+5BsaLV4TOkXbCkmAnfdRP
bHp2z+nbQqsytNB9N6oRs1JpCqRUzk92fKl62117rZBdtqo40oAENqDJVWjn
9wA8AHGKD6tz+fnCF+3hkzaCw0REvyyLvHh0OMXxq9eipXfz55diwOWhRDRg
PejGmNzUufjsrMH0o/6zLl/AMPCskwgK4T7/H/T6X7JbCummWBnc+orZmpHI
vqPD85KetQzwJ1/lWvzezu1KizsrcNzYhOACIr2U6e8CozkxU1RHJ07ESuUw
yX4XD+ZcP0pxtZHgWNozVEBfC2pVlgRmqzcumS97fMR0cmPKjQGqMeRruAAB
94MAFEASYhyJN++R8mQbbJ5ZJIJqg1jh6MikGZHOxl+98iFHrl84PLS2ixCC
kWy2c8WZnrP6Zd6pD/OzrEv43r524URC7KzXOXqPTcTOFMSw2pcmUSedNXsy
bfb2Zl9B/g7oU8uYJ2CV/K6WA5FNFGCO0X7HUb5IXebYYcvE95z7iO59apTN
nOPhFOZcPqnxmEMnh198UBURf83E+QDukG9e2ugtz5HPjUB54SumHZ7elxf9
WZUfVpDRz6vG1x8BF+2aKfqILD7/xOGwRrP/OiiDaXR5pWlnXgaGFxJu2ieL
hhHliVsECwMrJNMt70laWEu0DcOWj115W6P1VqnLSTHJ1p7QIhh1LuBm7gU9
Jeey5OMyk1Axu9qmVkzTZI2vL9JY2Ok84/3jNVijpmb5z0utpaLoTpyJCEyw
gdiplDDAHMbgFlO6bd1TOUlt/OKGXk7nhtJh7KZAC7BiwdRoqZACANnKgguT
fXie47hT0RddlBD0u93RnLpxYrNA7vqahuz3W65803AmYHuMw+FzjpH5JJcW
2Abeuze8o0AAmMAf6NXeeGa0AclHX5HsUWhSQr6tE/eRhMQo/slBBQXD4NCu
NNpbzT4CzCnwJzN0yR9gyAtsCKMSn/WRePayDRIUAkMJIRIVJzNfMLGrg3gP
01fRu8p6kNgizViTPJtLRmjnqBrAVpXrMkgFMbUnFmyJe7fgo/9/EQkRepb4
RmlbUGDgx8Ji3N63gMN7TzAzIWj4i8WoBwgJFs0iL5wbanGtVbgBCyDvaY76
mwgPC8yDoW3TdLU337OiDv56xMj+5HHXBr85ZHseF5YQ1JJ1q/1kiTpaiUV1
dI/8M3BhFs6sSTSj2ujlwK6RuiI+wLJ9glVDEBcZfY27U41CG42831Q4iB6v
sPeHrb14ENpTF32kD//ZaBXpAp7MNmSAqIvp978IyyQ1y+HliBfeMUXtNvz3
u/BuMfiF4DzPXSrefUYb0B+qWAclO+rZ0iUdknTFwzv2WL1LcGX+LWaa6D8x
WPYaxWDNTgVzw5dAVeYzqtjc0xizq9lVB1/16c795cVr/XM3J/ElSA8GjtqE
T0cy+//nGS+Ob1K1+RjVapX6m0uIbqT4BCptoIUbTaE0Brd7RKJawCYb/Kf+
6Z/qjDxu8M2Jc1++d6vjZwq8GgiV67MQDGCEq+dZY66LiDiOZLB67p5JIO0b
HO7blms+Kqw2Alr6jh9OuDRPbofjkNounQ0HKfGXwJvhJTr9UPvQpg+1kfHz
EYbGN7Tmqf1kmCGN938UjdYWHRFENO7uVlqGd3A17nBb5uqkdlWF9IMgVuJI
gZfVKY4hNp/5rW8/4+dRHO9yk/u3GMwi8Dbn3Pb7rln6LHhAIxlvd8OR/ui8
DZNlG16VmclDvNEkrThlT6ehs3CC1r67Odev28pfr93Ej0xmaGd5OmEOhI3l
770UISHtT+veKpmAZEp0S8rBr+PwcLbL5TOiCH9CAwsO5M27KmV17ECubGeB
+HSgnZO+nn1WGyPtuZZxJmVZoBeOr7AUqxxXbccuXx8UW7SV6G21SIja30/t
owDFrWXtTAzfKW/CKUjIgXqjA/IrnLfPu/6U6LWqMZ5psJ/lCuBX95HQjhda
H2I7mjHHkH9tNAa8tP1zlFPyqe2ZW4cG27V/qS4aCukmF54fMpeUOSp42pxu
tMi3mwL+D2PO7dzXMdxQfN394qb/pyMmwcmkWVkHc1nWOpQw03vqTB++NshF
gFY7YVjsw7zHT6QiUMFOt8DUvpp1iY2J9XRSqdEtuR/ZezG1iq+aoAGSwpdx
LE995PCHel8CXH8o5yvbvjNPBUSius/tKH6yrZFFPn8HEor2a4QrTirB40yu
8yZtQGwANlaoU1FO1nPmfuFOoF7X+0YSv+zTclwyF/hUUY5uuMN58LkB3bLk
0ce7jEHRY/Pfc597ymOGuMIYfMXZrF4lqe7euzqpcWPBgI+TYEHmOLAKWW4x
+Qw217yQeC5e4hwAC125Z2Fyi6rZJ/dn3BgnMjt4DBMopJGK34UzrSCqruCF
jhkV3Z3FKDr0l72Ayp3Ef170l2fICdOm8vZqyZ7HFKhBJP15ppZoK9e8aEgu
OR5XEAL8LcS8b3oMAuygMYjKdNWpQhWRV2q8eSdpP9sp/ZAka3ocp8Q6g/56
pHfh785gZ6a3vD5nVZjM0n+M/++tlMjYU/jQCpuDvoGO2RwuKCn6qUQtSOCU
eOtUSXhFiT2w//s5v3AMORou/obA/bfOA5+bXfqYr81w6iKt6JpCKWzSbAtB
LBMpLLCuYjBPfCotNxcsReDJ6TD6sWVnvlGztOQAzvAdYq66XS100SnIbHLF
e5OSgoTe5wSMW+T1J810PnBDS5eBmbDJsij4xZovw8jxo/6/8wA5ZUCQTJUN
YnuGs9qu9LlUsmrqIzkokVmdyP1elxunZ83FKf+7Rx53Xx6UEk3/KL4IbRPe
BHglGoZRt1p4XNpDn1sd9rIyUYxit0Vqu7bMQUoboZsti+yPIJfT7LXJXG21
t3ygNgd640ylgWFi8HHWjRRs5vAtehzAXf3wKQET+nPxLSzbIYnuzbEReIOS
H8CIrVxhvMeCTcosA3BDd2CtZBNAv+gj87rLiuTKsk4l6XtKXpYQtJuKvJoP
oTcDeOAdtfgNy5H7CxFKhjTczsUjfnqWIF4zU2eP7BsGUy1J1znbg/5MitFZ
0X0dc4DlwtoSqtWQ91S+fCl2+tMl6dieA5JPWVWcIJUpDtV+fx1yeJyiOS8x
569TxPfV57fAm7uaMxw36TtkWmkco4IqOguNPU0z8JXG37oVxOtjhrkkl1vQ
wLjpv6BkPYVsG5TUck0oUMJLJqyeOMlojqP3dkAZQUaYej/4eLsbEQFKDDPf
RVkLDto7g+stO3BukZmfnHtuCmHuUlp0gXvrP2AUjXJMSo3+/BY9YiBZVOas
D6BuTU9vUmVNYlmWsNcuzackGX+wM45Y+16u6supZC+pxw4gmm4e+WUy9r9E
n8t98rS1m96zgYzwVbSYJ4eGnxAyDpWo/BbZo4ZmBXDB8bICUBmQqgOsHQ/g
aDzBDJkYA8mN7lvAzChWZVkmq5yurx8kbnrtRu+xC2dCr4oeK04xdyDMsAsC
NZViKPhNbNaQiCSWEkicR2YtNVQCEN0HLbop4UkLnXFF6pow74Hy/XHDay4M
TILQZadX3XJ6YDc1X3Kx0MOzCUXgjs7piEK/pk1eF+w5SLLXjvF43We92irk
viegzjt0mGrondnD4j8zhCfiCZG8Cb01C6JkQU9SYSEpnCzvh3LRe3NWK4di
l/eZcIRq//eSpmyXVi6oOKR+JOLRAqXDZUR7PS/OqnQwxck6vtuadsi8UOVN
zM4lHF5efHanPoGjVsM+hy5cVJDcvGdTdonyOR+eio/zVh4+urfgWz2ThU1M
OnJFpNHcrx0fOjUzD7PmbQ5QvMeQozbwbiIEKZrfCiQHSN9KeN5QoUCKm2H4
eO2nXge5xuL44HR46jnp6EFjwAI5bPeyE7ygi33VRI2ZZvN/IlMqDFToLOeX
yFIyXuQ0uBqC5VR+mzwdutK5tRx4QBsI06sERL7r5TpRekzJLMLqkS3LgPJU
SO0S764yeVcED8iw26mIzJZSVXWNPSPYfVXzPtJRsx7alONa5w2sJEkhqLQv
Rn5GL8o3qt7GKC0iD5GPJOokKF3Nct3go5AhQMiwzuEvC2cwzF51za3QW1VO
1JmEF6x0ZtohfeYFU7R/tiedUftHT6UIfbR3Tge5OSUEzJw8iRIACRB2yIx4
+EUvjySbRSHYD0u3wNgJAONGS0dtoRNgp2HpgneEjh9juOdDU/C7lFTOfHUx
TcTS8C65ohxbtYLICFeQS9p63JvhWYwaCMqQnaMu0sjSxovuMt7dtri1ybvG
To+2xPy4uZKPbSqRyoGV1DeQ+WYYp24fMfpRpDScYKyYmwO2AKq+X50YY/32
NkwLj+5CneSBWzfRISh3AuaMSmUZBR+xbTyD6IdUoSkvmFSsAQwcPyck3SgN
C/CB3HFJ4CB3a7fd6YPtubypt2yAaN/HTpKvN4a7+wI5WZATiSt5EGMMYrK0
8FoHuvSTmoP6NogiwjHzVdiJviPRbR8XVFkz1Nfjkfki7BzgLaQKXKUOriLi
N4gm2lI8D5XBpFmGlOwk5Kwb5jFk8FKzh7vwmyXRQnfCDDueTQNKG2fa2sfp
62kb1mneSvjMbevRKnvDad89G3i2vlytivVpHAPnyn1/0gs67obSU5C67Bd0
xCyZQfp7+UDp7nDAyHBcHnMVTMeY3pC05fRV2+o3yXAXcUwJw1m/KJtafZ75
qlrKX+a6bzzJuUiXzxPeR80j+rt14IJdy+/u9XZvOEDF9vJ3dlqDi4mAiFkE
coGMUJU9NuOeZAgNbF9HcPXZE2clTwxlCZXtcUFq8Wq9EhCiY6wgBUX4c6yX
MaUXK7hWh+K3OXAJbn0JieIMppQKYfisGlwZ8xld6qGDzDTZHpgPPEnDrHxI
U6yv4GDwPg2x74CxFrLO0d6TX1k2xst2vIB3Rxiy5iixFyUdfqD51Kbz9CXF
q8XGFyPMGMKarSQZQAClNr4LqBzcD7I8h3PEfFTHPOwE3VwaEe78o+MS4CQX
yMHCNNryE4Xg7i7wzUO8wPxhwXoKxOq/n0kn2tCHTvTT36h+dZ3JP5W5nlqk
uRCJb3LB3Qe9aM4V0UJRQ1cvZ2WfK9waIHFVB0McvOffSfrb85glvbz6j8Op
hNZwIUYescO4g4vgvXQBGCreuFbmfD62xVxtDXXVHckN08PL0WAZyjnbEUmw
eQ19QVO1mNJkWiTFVZhK8cu3o8Su6IZU8bAoLrqLOHn/N0joFrn3mX+rcvAr
dNYVk01v8r/1bVa66Hr54xtqyiC7SP8Jj2py37nfCmue9FSZQVLbJUSbl+EI
BIyLkHJTM1eLbPY7qkLNM1c+gEV/xTjbU9IBd3/veKbyOk/KGHYkyWXftus7
F3fQjGNuCJGv+tzsfs8xuO8xe60i5L3pjMoF05Xrw/d4MlMG9lSkAFNnRw0q
PhLrAZ4Z2/0xpfGLZFhGfSMQAMkCROdnIGkv+w4eOq1lTz7aMJ7nOWcZx81S
4L6/D+v/deFc0aINOTfoZSUh1olDOYt/qCoNzsYTb98hu2ALgJZEBGhF3E/1
tfT2aP9xKfz6lJlxRq35aB80rKWwrobHl5j4jx5oZQV+n4PNSK3P15nisFNQ
0AFBVC+5S6/CbB+sDXJJGSuRUzjtOi5i2HM2tj+w+7I30JmCxTx2X8q1P8I6
IbxdchkXpxND8BzQUoKVQR7M+ZZCFLdreY5qhTCMxthYiAIpD9e3Au43XHgA
kAFZMvPol6astuRi6FXT1YG5jHovGpDFkEeFE3I7Ac4wHzWRuC8CpJ/y0cSQ
irXBMSpeV8pgBlpdfshYLzEOpn+RpI5EDweF0HRa3aLeqmPXMyi/rVD7cIUM
VFETyfxZlInMMyBHDD4piY6LaUhsphY3gd1tFXj6UKDQ0XhcdGUN8LQMTHAG
EoHWqY2TXZGOhIjIwsCCKLtl0js7q0QE62CQx03yYGvTXfirYwXG//c6NNyy
uTFnKUeETbHoliv3aBQvmkaGIa07MAVs4kMkXKJv7h1sphpNal06PPIIW4N1
Dy1GywAh17XmcJpdY2pCi2a7z7fv686FAZPOlqy0lw0isHK2wOG0AxA/28EC
P49lqFxiaVwBYt7M2k8kl1hIen9Wqu5cmGCaZh+ntbOfVZ2nN9NEKOmQOPrj
yi+qsXKSWLXkmDXKYd3loT6lpB/rcq4H3Sioq9INpSnWP+Mm8vyBBsNu6Oo1
fcDiWIErakjyX6ILo9fxRp0zcXpo43mFpJ1ImpDu/jFz8TMjAgTzXd/KqxHM
dIBWrKqY/7wD/zKB6kWYLdV8022dtwlpALqOb6P4xxG8PLyFkgS9pLdguODI
4ttkwtP0uxyF0URieF1jjD8o4cbzyB2oS2NDHvUBfwrEZnbV20IjfvhY+kJ4
bOb4lYUkhTR+wxfe0rklEHoivF3jfOmKrivc9lT8Q7Hmit09ZbFfCoKISAL1
grhUJuqOQfV9viaH7XQtEMWsNzOWWWlMdujWULfuSM78svnlQH59GxFAYcDS
dcUEBS+pd/rVwJGQAvzw6GJKr1eXmSO1aEhnzcKvCWVwnZ5jrBdQli1O5e7S
om+nrCLuY2lVGMioHMG0hTLHITU2efFPhThytab3kGiXGA6J/ytWMKfHVrMz
HOqUp+2mzPEIX0asY/UGj1ON9+D0BZJ/ST20aa+6jOJJkFPPJTiAzVzKQdpb
8UBbda+QnrnWaJRXwiLym/5C+lk5g8SSzzJWxTWBCUvd8ifgPDsVFYJc7fkd
xgbBEMsr1spv+cAVbVPy5J+ugEc9j/iiMPhr1DxQBungAUBNLEgRhsZ3iIX4
En7+8cBspy8wIPwzT5FqdW+HO+xJJOxtDQRyT1oe65Rzs7lnVjoS7GJVVDWv
qXHu/4c2YdvnD+aMHIKBXMoiDWXUO6VWuqdJU2C+6WoI1IhWS1Opl07XYaU4
IxQ0wxYG04YdAxquDLOJ3+MFi2dvSvOprRMMqLNcb1ITELJd8Wa+Q8XpMjOo
oKvuPN+tndwJMTRqIgviwli3nS6vbIdZUPFyDGYdYNfrrPbsDQQ+DKiKIBkg
woC766nalgvdPnHDjm+tZW4v8aFyR3UGKqQZqBsQ8GdnChU4ovSEycwkAwht
jyZYWcBiml5xSiO+UsxBmO215XtUx44EQiOUCSdNI0/p3LMjjALFPFYCP9FS
RyFZr592ADF135oVA1yObpkF3N0lAK0+IGTbtCcwZfxYOP8IERUad190x0Uf
bSfS81WXrHpWE+gjbaDfpWRs0YaYnHNOFuEW29pGiXCdtsQJujkN77wQd2aN
SAMaN7WUbXEqBgjiEOeLEm4bZ6SuB7SlWTWSYMTiirsNj4yQf4UjlMK+LHHt
lrsRwN6Gp+S6Tsh3LUm5a1Is3WVMdE9gO9U1D1jUj/jJ0kUF1x/tm6EXKbfB
0ZUsjjWbOMTBvztUgqY/NuWmr9NmzTUFtoGILsYDvBraLOSF27OSvpa8S+Le
8m0B8/o73hKO3cfQO8bD4U0b8NxRpJ8fjcuvM+zAUgXIKWvZY96zHg9NHICV
jupIcTrCVVbyZtI44PpOz3IOhiQU/4UlcJm9S6sHcxoCFt9mC+haf2pFJYcq
RqSxiIQwiRCSZ3lxy07yuAKbsfmfG45vjCb6gx+97Vv7Jf8EC5pcuFqWMbhg
5ZDZ6SV0la5Cb3jR0SuBpabYOWqhq5sfLJ9WVFGyCJxhEu9saPsoJRIPit+4
ByA6yZy1+riQ6rGQpn92SSswCVuV/eRTG4VhW6W6Lo1E475glLZuSCvkYvIE
GWzigfq4W72afP2dLu9MnJrVRlSvibCKOkm9qqxBxF/uD9cvyDLlLu2/AfEe
3XZJqD3hDtM2r0hxBs7aviS/9TPj/akXNRA3lFTJiQiEPlG/L8N+oNxHULI9
8NafV/lQxv1uIEWYYtsRKdXJV4/9OpVWXJIyMSiszUQNNqvW0Q1PrLO1MeLH
yVQOVal8B1zL6Z5yqkvv2vUyyoH9Z0yQCwEhfG4talVEF1EJp+lv+ey/vRyF
sQzHYga6Rlg41s6gN8JJy2cRYhtpK34Z9OidBa5NyVPC/S5MXyK+jQkbRcCj
8v0rrcDqwAtL8fWzHYOspIM8mBW4Cw+Z3ZVtKIkZgGMqOXa31bwFGVwTbU6c
fz9Cg1SafxbC2uPH81DKCzK5+00TBZvoBeR7tBHOAZxdhEN2Xx+ucdAn1a3j
UFE4Z9m5T9MRNBB2YTIekUBQd04F5Sx619k+GkX35aM/ewQQXbxX0svVx7F6
j48qGEPYsnnE+IxDWSyTTyd2CyTlX/kbVM3oXd/MND3mOFTgJBjWYC/n9IZy
KhLnQ9TIDK0Zn5z6NXtPx4fXIjOrVY642KPQXHRveCtGG25sG6F4cbUS1MBx
3ccFnx9593qGgPApOTRwKvAxwVhTswq9fQS3CY/j4QUTJ/1BEbh+XPDZAXw7
GnJIPdUyChqQNkSIQgj3UprHEyF97qIAh0Jj5Q5Uoz7f8Y8x9XeyoR7GgITZ
mzVkTsp7gxhhEGiBIqKGQxgqI43RWLX/+G/B0ZEUgzgUtHawqa131CkFSMkG
Qi3dU4rUgyhQgbZER01M+YXlU7xLeOiTUL8MnmSRbkSrK3nDF3gIKOHv8lDW
VyfNtFpGSSWd4yHu1IEGvHpvNnYLjBzW1EmIL9Dug/Hg+DKLXXmzMxeQPxV8
6dXUm5YYh8nH0QlCniLZLcRybfApKQtd1Onjo8/waz4KikxdVmGOD+EdIJgB
dmu+xNQUJ0JMNK57j9jB1pJPaQXZq3oyyqv388QCotlqeHAdQa36pwyFFlRo
KMxQHA+RlwrS77PlGLCcgkP4v4oBd+GRwCnQ+h3SMdg38KPYjTiwKqdY+jYZ
LTBKGh7K3hUDbezUa5d6mSl3ecrlKPHevU7IBQc70X+DV1YBbRjXtYg4WjVX
mjdVscL4S0TIOsslGCsnW5bTG/HuIakJGtI41XD+6yayWn+yHLvrCm+Fmykj
p6Cu3+Elizk1yCikEIlNIa84TKnWsVRaJX0ByOkBEyDh35E6AeptK/2V7/Eh
CB/aHkKFE2LtIl81gYINa+nVIYfc882neb9x41aCvo4mwVX8/XzCgeXihNi0
/lEr58VdwP4j88PnWKoVUg5clrKXkuFOo7vVJfYln/cVbe7R1H+NOjWA62Kb
CpRKaC/3RDXaftqOnLaQO1P+4SH9F4/z3Yat68YFmVGZZ9arM3DmVeH8fqmq
OkuQbsqYoV1xOyjTcoSTv5n446Z97DV4dHlHzJ7fIW3phYwxQlCcLLoKRqC8
EsvZuwUMIr+JmtvbL1/LgeiJCu+qqIk7QF46xfaKZZtnuJqRKJIyCSUYo9zk
fHyivty2DlKezF8qOxTDhee2MObiTJ/+PrIVLg51uW+xg9zujFoAfl1BMa8U
IBfSxJEjIxUFaEdmB4HVmozMD8lvQskes5vtf4r3an1FdIF/JPkOo428Q4gH
pm6PiE9E4NVJntMtC4RgBbbUAn1bjj2lC9nQ4sTWxy3Vbhkyj/HRmaQ6xWcj
+z3bwChh+ge+OkMGAgLgcSUzB7ZdANDMoJEE9mZDySexiJwuA/ohkPNp/Fn6
Isow476rKU59mClSSUEgcfUTZDNkCh1xO8jS2WV+gcK4GVtBj8mwSEri71rw
dlW+NFzEDAYVpQD7ftHFMZdDSQdnCbCDjwX239PRRTNekO0LxCoC/HPNeQI4
oO04+/pK/suimzF3dKr+6AkiARUWeR72/3eacamjsVQTMvAdqDRPVBODKGfo
0T2A8BmQNK8O7KZkw6oRf7vK6GMz/1ykK2qlvuwSW+zfQlQcNgv/L7k+4680
lli+zMAHPLNPYXLDK8KxsCwmoSPacQhcyroxl+LC9EuxOVFkj0w/SQThROFm
pEUOXDDJnRBcE6TOdUGU1HguohjXd9eSeMFqQ3e4g5HYoE275GTsJ8Ow0h4Q
d6tw8w1NJTeOlTlMUh8/O07rQUfJFsjXmNjA97bQSGeaEyldaMTJ1n4aGiSo
R5wadUiWlCPiootQ3Ln3u4wosjdLBPsLcD7kEJR0Y47OUud/xM+OQBTUUHoo
NjiVcleOAwkgElENAb6fw9aLDQjdxkbALclGz1xK1k4AJL10B+8KF6W7S+iK
I6GgFZ9gYzLfRqSTvMCBdEP2KDR3kVpD+6Iygqn+wthYNzj+Ieh67Qm9cuuo
ok/rHSpL7rZJQhMlnL1ZzufolhCQ78z4nqZml+ti3WoV9cVXG9Lu/l9qs53s
ddrMVleb4wSJdyJjCJe9JrdbSZEggfh/MZvudU6caGSsxoqb3J8XVE3dIQHN
0PIzxX81cIKBXS9jS5WmnlAi2fgzvLJ05vjfOAzNPCkv7eH8bb/OcMRJq+Oi
0cyCcmTSKpONTg1jwS5F2fNyI/f6VxU15gQDX021qnR41ZSrssxgSQCHXGBX
PTuNUw+Rwv56xAgt/+Fm2mDMZqqlTJeBoH2KrwSnZlrkwxExFVQPlZqQzkgO
wU8pKXdT+hX2wQUJRf2ZtXE5Pq/CHdFKrAm83ZJ3G63BM2aQBQgW/RXeFp4X
LYbVkZxjuaxN2kehMTYuSZtNZXs1B5CSyA6CB4KCviOFOG/QhEHfSk+429Py
VPEywYE51JprRfU/w4D4lCAkuIBo1yzVtH4k0cPSAC/pXjztOhG4tUUbjCeJ
SZDuiRJ3hPEKlY5wXwmUkeGvVCGJ/F+oMbOlQp4sc9Kpt7ufsOTm8rrC3NSo
kZTnvb6GxpDbLHrby51Z63M8a01mxPKXJj1jrRw61PDMc7ELW2ujDtHiCqxn
Er3qdPU2sfJ9O9Q+TY4oD5On0kqHO7SRp5T3LlSX3eP+6mHYxzgcv6HHLqSQ
OQn4+yk4K29jPZ1+3JFkH03o//PlGK8poKQ54U5MEL0DczVMIi/VF56x1ejP
QroK4H7MiPhlvBjVi0D1dicbRqd0HbzxsJEpquSKdyeuHabQ6UeM2Dr6SS42
EB4wWM0cfeKY+XKIwwCW9P1/fpjtyWZJJlwJ2y/A85D+sZYkJZWE9B+KvaNo
VNmfRBNeN8pZwULMOHr2beToGcndy7cmMFKhbv8Ev3nGKiocUtqmeJRbYlzD
OoBkp9xM9/YK+ZkbAVsbl6lmszNc2CijVCssV2cjTlROGFjT1KU7o+OkTwno
CNwaGbEecIz8BMib9QkW0ZbjeA9Zyb/blUzpJNDvbZ4y/eA7CAjzUNQZCP6X
rMrmUMVcwCJIqcp6/2b9QUmvgox+8Ln3dNsBWXo3vHENm8dwjQFOFtUPSoJw
IQ6J+Qy5DkghBIv+zdvTjl6bXwQ67DxFXS7w5Daq9rTub47+SRPAKTFzXbZn
FVTpopX5ib6nU7yPcsHCldt4tqAsFSabyGlcXbJjRgYG+grnxyrm1PQkOvuK
5x5o0hbE5zPW4uZ96CZ2MVXiqYfJHyuDvbG9Ihyhnhi6ZVo5Iqe+hykO2v3L
tifskiCBtlgJIAHEtM+ddOUxbu0pVNlTo/TpVTTvQ+Y3rXGp/iwt2TDtwjey
1n6/QnwibB+eGNsv6KkIoHfK9+ssKHQLYcm5X2Zbywaw4+11tCjG/GEMpNYV
gpJPzv1VO87V07uDyxnUyLmDfGbukyr+Qdn8sFK5ndQQW2CaTFSRUXHu7Us/
Qj2d0ahZLRNm2Zgm2CkP31PKBWqVsx1QtDqhVYzbI78vPjaJCXCC/sG9/d7w
s8l07Y8bdbgH1q5GZfR5umiQBsZlGlVbPOJSR3+nGvUPjqlAeRlfTBz/6qOB
avPTMjmOU7q76ME4sMGHXBnokPDaiBqwU7nGgc1+2+aEaMN37nGUUHYoEHZZ
uA5/1OaacpImRHRNNNGAGrkA/pOCP0x7vBckkoTnhWEMpJKr6llfEGrRU3kn
HX0y6nT1szNsi2QjbdRL1RWbCxxbcsAezIAWVDiWawZlLxXlPeZT3R3vWIse
ci2tzi5ReflnPAVoPTNGpWsKFuEwiCtv2E+C5drSMfZ/zhZ/zpiXMq0b9DTX
r2BuOg56JSgjcJlLU+rJDK+sevn8ExB6DfCOsOHHsCNetsvYq6qTsNkHRhw1
F9Jbr0/ak4x5rxErokSeRdPOL028C8ve0co+8G/wDn4YkPOtbX0Hr3AHRbyZ
Zj11H3BvHrLzdzmpoZvt24KTILjXKWJ0b4Lymbix7BFUCjzfo1fXBvnMZvN9
cSN4LqdwnMMauegW4E/SEVnHC762XYddOqPKEL73nqF0maXxSP6zix0LGwmp
pGDFBrecd4qBpr5/vW9m8LKPzI7Rl4cc7SgPt36LggAsQTp6sjd8S4ETqKFl
x7zoYV7bPrnR76bNUBPUVQAsgxR+FxbTvi1OllY+yNHQgOj8VAdJoJp0hsLR
cG/002GJgAyxaG6p1A5ZPdN5hOkmcMnHTjuVw60TsUu1i3C46Af6Zgm7k5Pc
otRgPFfgPokleNVJbbaQXPDE8gEZCCdfIHzDXx+RK1I8kAfnDs0Wh0vhhVD/
hVFKys4xOsIjyNGezFTe7wafJcmWn5GCyW8qYQVu6+y7dN40iTxiQsfk1GnK
qTfEzr/EgyWwdt87DPipkwSdHlnLZgsSaDiN+o3Pl+Sf1uOZJac4z7Gf/oye
BnYTKawSv8xkKwKph4EiGPCe0Txn6p7G3+F664Iy3SKZV5MmPFgzKQFuRTQg
u5KWvyZQjuhOUExEenoGnjAKZbbM9r7JvSBeFy3kIJYUH566zkuAi4HxjmWn
nHXVvWf6hdN8wXXDoJlQqL9a1L+U7h5ckecM+hVYcmvQ359QBAr+2kVIvufk
obmbw+0lbON+0EgwkaQDOt8oCSP7CR1Ieb2npT2XcUu+MizZtBCYoIqmMfTf
cIBIHoRRQ9HAHYRIuMUGeRBDBhzphZtCa/q5Ej+fHiF5WA0Wsdw5nCUOre1P
rFwP7+DZ2z+Aqqtxl2pLOvidO30HJ5f9YMoSQnMWarP1mW383zum4lCcrQMa
4UmtIRXZL7qeR6rJUWgeZeJ857uITt6IZb2+HYdW+zT7YBViJodb9IAR4g1r
Pp8lW3KUWuLAhensdBrUG2mdTna6ixd8TIWQ0XczneDFfxwoQ2EXh+A8jdVO
sK/DBrG+MuXksJzGOw7GlBStryDItiXLmJp5oWl2+5Y5/cxYZ6SqXEKO2bLM
kxFLJl0pn3CP93kGgImUP275+NzrT/XU9LvXOfZ074ZwEG0n3SdhjKw4azVE
7kkGkFIZXwlLKNw6gkdF7RYLC3yIXAywwZcWe4j0GD4V3gbURr48AyaPgMUo
IhYprvKjuUrFA2kIdFFKuZC6zCW0/ERknoaztq/tja61KVQBZH41EdUZUIsy
YL6PZXmOpglG5FoI2FKjoAUonWuYD+ZHVggeOXzMTf8/6UShpCOok/eHMzmY
jkoWFF5Z3icAfwhfZPfMc5ZhefevoCDsbWUqk0nELao2KTFFieoU0k7z8bEV
FBOLwOLTKUVH2qIBWKtRVU3ThFD93Q1zz5t0vNBXbA76b/EobV3xPdDjnBBd
VBDRBDpyZdFpHAky0ADAXTgv/ZV/jm+UXekRzOeym20DXhChcGIHcmTGETqF
yaRk8liYVNUp1Xh5Ocjd6cuw47FGcm/AKRedpDUHiOFcM6k2hcNi4hQjiFPo
fbmxZjT/AiyeuVddXEwLpptLplrCm758KUfYhy43HJQiImGgsptwGth7n+rv
GfwUPchh6HVuZQGSn4IhMCxYQdewOFCBtl393ysB9KNobRyaVJvR14dJT0l7
dBOQduxTo0FXM7Yq7R4Oc1loLI0awQ7rL0ve7VCCNMiFlFSU6wSR3/URg/bF
OT9AWgBjG4sglcpQ29qSkM/+yX8Isd857R5l0GTjj0pjJM0zpglmSwli1oyW
ptLG65U13mS3/CVSt3tSaOgsr2LCjh9+Npw27NZVd69hzLxMRBMtaux34Sux
q1UOkQwv00AcRzOA12fdZkYw15070MlZgm2SaKiFqVt4bUuRaXLZdsFfnKQ5
F0vN15Yf8NdVHWfgEAbR0rUaqdl+kzOH8G+dIwvUf2iN2erFDE18ItRvxW3f
T6PTFxYNHYdSPwJshizeVehWdoTfjmgowxrN3oWLFNyksygalmEiR0UrxnAy
YSAG1PMB3Glo3a9JwF+4k+vahHCyliyj4ciMq9YCvJizrVGVGwYeF/VEqAVu
kiG/nWUydYIT4Y7yEgAOGQJlA9HqsmuQxPDCwD0OdNvuz7j9knrLF+fV1BYp
Lj4fVVph0iwOH01aYmQbhpmaN6kZV0rNi8PR2EUmhZFiFRSCbkTD8N4UE8DX
7SrmddzHBrZjBoJLFk5j/S5sUthg5DkZVEmXBVjlkpruAmR6vSPKEFuv6jN1
KhMxupzI7v9RiaVdwrXV/ZbASxSKxWdchkarORHcq4qh3pj8tRUIO0SOQF+Z
5vjVIv/FOsA3rQxnrtGCeoBE/xiF4sQzTuJdHm3Bw47owR2+QUdK2LCd2bdc
a8wWQPk0+xZvNK+M4PLuR6RKTBe8hQ+I+vO8pcVeUBH1tgUtrwukVBQXYlua
vzUAG6pYZ0o6w/6j+jPk59SYPHjLbmyepo1mqAzSe7wWuHxerT85QNRJKA8+
4e0Lh3MspWlREo3yUKTwGuG1+Vb/cfO9FYqT79rh+e8LmjO6U9TRpTi1Fxvl
IzmH7VNtZMU04TlU/+W6sydKt8gx1PRfxR7H+58WY665gd553btN/VKXfTx0
O2OsAvMtq9KgsrEmdX/hBolNNmjiOnekQUdaRBPfJhpTEbP+8DPdkXlZKibR
2awGHIS2cTQh5XXdQtrZMD3dr8YDeLjTrS/g88RcQpBREeoinuiC3Prkq09W
zQZx8UMbtlB9Ig/4FqY73AkMudbWOwZphSwi4ud6c/fkBdZUNYXVTrOfR5sS
i3wfkbi9s57kRmSgDUEq4K7UZy433ZVE+y6zd+ZEIDwqQGZDk4xBBH1lrw6D
KiuLrV8BggaHKc6+t92IdY5pDK1EH9fixF53tVI/KmH+JyqSMYSY37m3FaAx
PUS4bGAG3tbfIXttWfzbdsq6Z9BZtyCvPjBlBZTS5Kt9kLg9qZOVCD4sFfve
cjNMCW1PEMZW9BMoFDmDRchnELfV7Kn2HJU1Co1y801p2txeLgtt1rqr8BCg
iWpGmP3KpbuHYjmstpOAnJlYdoNKMRh4qxS9XAey0N91UL1JlWKBIuDPlQOc
7etduxy5eQjSTbL4p9ZShicKwR+0haPizHgjCjJSlw2NEQ3vIYnh2cU1kJGV
YLtk14IDti8Y/HALO+cEwX6SJi8X5GYecFbCcWZoGtomShUthrzi10mEyak7
3avoiB5sYmF/ncJzEDC/ZQJxZSaNoBU9fLjeznSaU+eko/oCpvh2AZYBKeG0
3xbihdEHaXGly5Aq44jZRNSp9a/9VXJec3xu2nwkuWjsPvWrMuZKiQqjqBz6
rsJeg09lpyvBD1A2v+3iiyIfG46LYQwjjI90BRPD21TUftPIXOCsE4Ms+AF4
XB9cgP+o674//E4Fpk85hegKGHHOZvadMuCu/eB/tMkv5ScaZdXmWKqDUmjp
FvfpbkrEVGYw5/XliCRP+aTILtAv8lPBQtYU7jSD3QmcfuPEQcp5NWrS3f2r
QViWMkUVLlk+ErqgboKXdQBG0gZcQwO+6D/SaZKr8VP7hDxGgbcLg5sCCUJn
MUPjWZcYlcS5BFXCpLNxCYcCOshP6kE/Cjd+pQBTupJLQIVSjfGTQBZ9UjJC
Xa1lTmv44vVJT0O753w8kgRz3FneHmHJP3rc+bI0grvkPLcAvN0o4aqygUQo
f1Z7BdZNHQ6soQTDov10ZpoeECQIfIqpKPKoFIgs6f9fZBgF5qpEeFiR/heP
KpgbwA66s5q8o+c7ySAyhES2GFDmJJBY+2hjzBvO+UsxycWih4TmmiQJN7IF
MvU7G5uKMUu/CZA8CXYnH3ECzPCP4h911ZJ7aEIAZGe9Q6lGHaWgAptpLktY
1uN7O9Ukt0wkhiw4CJIow84L+LheRaST5oLKDUpR5EIfYBlDFG3afOxlT5by
slmUz8l8Wh7YbqbI4nsI+sbhR88r6oolejsSd+uGMT77Z9XdKjpSpr31MMH5
D7twOVBtPQlj/YwzwXmxh4xQar5xqlHoAgYCiqukKghDisaooCw44jMwPxKZ
ox7pUwZz+xg4tIXlcw22NuZpenSA9LuNyxiPGY1CPDC0bWZRe+TiY6bpru6h
Kil4e3XfjnV5jVfErUfkU+atzAU+ZNGSDfBr7Vlv2t6sUd9EMggSwJnhaAqx
KC11OgI6XgsBdI1dxrEbCRCWfviIZU70vCFwVGhn/zgop7Hs8Yh7tWFUcgMy
qEm0kQMqhOdOg2MCjb3+wSAfFnus4HoqkxsfjT+VCz6rZJKF7Ny9uYPjxkSq
BuKK2tE/kN8Vbzd8IsKgy6h+JJwNK6LlXTQzQqeYgAnhm9PB9TXpV5VxbOyK
bJSbokCrWQLbOx5Ocy6yDWRqVNO4SXxlx1fofUeUKXBP0r2PqkuQtaxAhw3f
bb7HV/A9wsJnbgQ16TLOCxUwYkOTEnIcElaQjdVTEHSMMOjmukx3NXf9qHos
yz9SeLGHoHvkJRvgFP+/RIwu39JgMqIAodLndNxKGdr/noFr2XYwAk/ykoai
9qGTv9dmHUDmbRoFsvcBrqz5HIYqMfVhTDrkexFp6/x5jRfmKj6Li3Fk/Wpr
Y6FmNPOWOaZ02LpkFR4BZkervE/0+/v3bHllqgfcSYE9+jAsjsXa+IOpFOH5
pwZcjwnaW2TPDBkm6QMPPtWiVBXssJ5+RCSkvP8FPO99rnHzXaLvGgH5uViq
I2uaxhUhBNHpkRteQC0zsp6vXQqmHMKNUTv+u+ZoBIFTdI7/hSxmkQTK14wM
zHHuUoEpzYO0GlKXO0c19WXd7/X0KEbfVB41qcflWVURmXWiwdGTyPgKvntn
lhBlDBm1iUufp5VydJph3UjExkBEyZFzQe+QF0cjKTLj3pF/6utW1+gEJUMB
P7s9BWzrx50k0KRbpdlthee7ny/9cENOIVZPIk+nUR+OGSp+8WimrUyv89Dn
SjOL5lYn984AU9av/y/cPJpi+pJzsC53JXHkJlVV0eDTjcLmJtmUCS3cIpiH
BJKge1NUxOF8TKIXJzitUUw1jGktvtJCPo3m6gvP9WQcGoOloiWQ0axflQEh
m/P+IxEg4StOP3jMinPNpNcBJNC+oDydPhLyHl/XozjzS+fsVQXTgs5cGYM0
/EW9tC9rc/vOEQ6wTf1xdLZF9bjZb+fkkWm6dbczyOJyqBaAGmG37aOdduNU
NKUgnv3/ZQjMyRJFGJ7YPVpZPrOYtLyYsNrPjYeFkeKZS7Is1dQ0nDgb2anF
mwO57b2Tlb1pr0rPlmYS4euZHhaVhsz0rIQs5IH+k+p3Fq2A0WUW2V3oxmtl
LNDTRkjxhSjKoza8I91N31pwX2U3Z+ESLl1O14pnby3X/BAb7CuTJSmo7G6b
HdTMNiFVBNIodFHAJiYETWR8s870o0A2G0CFy/zxymXv0q/z+WFdXrbcOIFn
uqm0UUd/04NUPGslIhZnWkdX5UA9eIrair0AkVrd/NZzx1le9vNkDs46Bd9A
KvroYpvbkbXHsFMGs2Sjpx9fboWybDCFFTRDRBqy3OihVt7WsS7kr1TJ5Lns
vcQlvEQ1BEm0AxqWzWI858rD6UMjPg6RLRlCsAGFgeJ7M5RyVlUIoAY0Jk9g
FDN8p2M2whooZCnS0rRml/fWbsssBrbTluH3k1VytkI6/szFh+QkdqpSenM4
X+DfO8w3fRI/1niIWctQGQqmPrxDGg78EzIyImllfv9kIQ82BKAdCvsUSyRW
033C/emcfyXWjdS1EZMd3yxZWwNATajTuoXbPQHONTbCfy7AFW4nUQjcItku
5n9J9L0EbXJhKK/bqO2umGiHa+oJ0DuAnNiFHIK8RjdmQPr3DjTRWptmF/LZ
wLOsXC7cUtPPnyjNYQ3TBuzcYzdSwzgC4F+LHSz8D4zIoukEK7X7m0vR4iOw
AuC8eRCuBLu2CI26kzr4qe2YwMJ40hPOzY44I7AXrin9py+SUJxb8AZcLuWC
t7FlXUbnlfYpjjYOU31uKQDIWuVpVx1JME/ue3pRN2cezWIFJ82+/1F3ilQU
ePVmKaF2lUV6fx5Ntx1eWjwiwDry1mSOpr/1eYMVX1HArYyGVg7QGexxfT0Y
ZNVVOy7e6l+ZLVz5uuZF0oPaC4/Lj6G+IMbOdG7sTrgt+RTdrf1rttcc6pNb
ASrXvB7ZKHH6wQIZPYhdu5YdXmRGgcHkQ0IwVhTdfuu/OVzkJHuQkZrCVRR6
kUP/gyEFMfHj1CVTGeXYW82WzI7OCzn7lvwcKp5OECDG8sooEplRPdaN98d6
hPNXem/mMBNRr5QjoVVALQiQ3L/NcnPHLcRotgrwAATVPP7Cdgl5HbkWM2ND
hpuonEtF0+Z5Mgf5xnCpmAuv8oJsZIrIpESP3OOziqHWFp2G/CSEL2bdSgqX
RoINwAnxPdu0pZ57CISn3fHoXP6iK1phc0Kf4Sk8uEqFhcj1/ip77q/2R6fR
UNfaVUJJs5/j1j3hPJ+4IU9isq35nyMnQ+AeCcW1VtWimPri0Q7osu+7tPbo
oxOhhMvZjtQDyQfNS7POufQbaqz/QBqkSQ2RY52K7F386Y4/0Xcap2wis7JI
vVgdLoLyhbvEAUcCaykxitdozoImFPTMPBn3UHQ8qcGj+45WXIhe/cza2o5E
ZSnSrBXO4UZGrsG/Fwpn5m4mQL2vYQB4Qn+jh0Vxt9Loh7G/3fGXknEAhq6U
zAHhsZMS2b5uxrIgUDxxOoe6cfn7pVBCnHDflrrdDHeV5gRZb/0t4sYPjJfA
Jp48EWDMM/0eu7FWw7Csa1RWmnLBfhB6k4BZ4rMyWkJJNG7mzIcVEIhU46Cu
WHwmSbbhWn/YWWQ4qD44tgOzGd+/LVaDAI0gAJn+QH8URKLm7V27gKtpJxVk
J6lxF+ZfoCuKsxVuHPL7jqEQwcK4dR/fvdTx/t5KV1eyhN+ZP5WnqsggBibP
kxvgnMP83rs0WQ4KlO/ut3GMnryZ0eE74TujJZ1byBUtZ/Esjrxj2lU6HWDG
A96S3ECL+E+B1HZr9A9kdnlvqo+v+qpC0I2TkHAiN/Omd2qI4Kif1bLF0x+a
ugBOeEq9N8dvEPeJjTOHzYvfTJWLy+mpE2aICHTMCQEjGovrfrQg1C/1l6gC
iC9DmZbarnJVaFe8zRMdnMN+WwlSajRo+s+riNcIMY0smdxpFIQWlmTyT2GG
GbRZQV3R1W/6Url9uMDLPUXDBBUutG79euJBA69+wU/VpLIHOZ2F51AhRw3+
dGcy5eNb19ELSrbLb3RdPxhBwcaKuACbYsTqzkxSSJDEdUKRlcYHZJQvRtPo
Iv59r+fkYRU5tPvpFIVLnF1sjPVHXF2MIjFR6GCJhripEsVpkeTacagOA+yP
1F5pQVbwOHhTe5Ak287lpNrV34uMpdtd9uDH3MJpZnsOuvy7ei1unjSjS9va
3iyAg6qqtjHsSX+ARf+cLOftLw0mo1ACqIv7piAlG2QSxthq2ARMMpYrrWxo
t+/DACuCCzJs//aA6hFcC6+d8w7b8Op1VzVL5KorVNBi5EU5RMuRIdTF1bSn
uIVQBlCBpmA9HMkuXZMMhxhMFli7XcVxXiN8n/cRWA6sLHHOXTj2rnCxq2ON
6GjP0rbkxQ/lIQr3rT62wJLErYxwEw8HKBeVaWot4v7mRIOkVzahy9cP0JmD
Id4c8b1W8H3GgVkPpk01tdh+OKFlkkyXtAJfsHtZQ1O9yAOQl8kRXCupemd3
hTmAm6YSfIcVisSwg5xIZdJYLublcPuf5qe2pabJWZyNfaFoCOlVMG1r7Txd
sVErE/XFOaabjulElr5lg/gyu9uI6zvyZXgzYlrmUu8i6cXOYzJ3G040ubGs
DDAK7mDhfWFMZd6YktMDl6jIdgK73Mclt0sTiGbDbdVPAZCBRUA7OfNryJLr
MSOa7BWX5uwbIpJ18JpCwjy567t9dtPXfJDqiV+RcyzxZ6GhQMqWq6FRhfvB
/SxSgABKlweWn5earvYeoNQ7pLsDmZeiYM5NsLUAM30Y7hD/imo1Y6wgR4KI
0JtPKYskRNWrIvIJCzvdP8mjVwV0Adyyn8rI477aMtRTD6ixrusBeJ1PyhzI
WujyAfa52j/5iv+loEdb2JlgYbc6Rtme0WHWhnyzEnp3emt8xQBfYRX6ub8i
iIisn8IwwcxOtvmnwg1w2trpvoU2CRscacvhob3eTlssk10rQVE/MLBPwY3O
R4zyhD7U0xLBKdq1E715TrAfR5YTCj8Qb4zgXkpEKgTOEGFgEqoV3X2TykXI
dGoMdl/tSio6lr6dY3wU8FrGDOR7vVsU4yy70BoiCfCiZMHFtyNRhwNedNrR
6zw/xK0dEWjcypejrvDeXxR4d+I1+SVy7QnYo38rlZBxdCsvjOouZrxY5gpc
bGb7G6M8X6FwM/jwDhGj84R52xZg1a6h3S2JLxmpOJZPOJJHbhfM/PClA1tJ
/4SzNjDWjHKrKTt8yHqC3K5cbjukLSQ5X/3VCvJcQfgvTYUm4mdamzvu86k2
ig28XbILuFmOioMc1NM+suXZj68t2ni7lQb6rVvdccgiQQB/4q2CDXWRyUJB
uPQhQu324T3qF8i24eJUDbTotWSqVZvsuSXiStk6CId4wcqlW9hGOqjFmOP7
zKVZPYsXBpfwnI5qkD8OCZnvsLnyQgK0qKAx5QWtinTIHuIveC0pL3B1QcqY
7mC0pMrj/Ty5kzvqW9OR0C2g4EB8LxElxzw1KCdMyfIQKYmgcWkn63/dY4Yz
FYzh98bTWyi37ApcwhqM4ZgX0W2Hdb4/yB2Y5s+Eky19/Vn61RNfyAyLxp0m
2qiXMYz+7ASTv2M/tDy6ZV9KXBytObfSj5WKZU1t8xihJuiCmy/Q/0c+dyRn
wu8YoJoI/Ga8X5zBacA08aGkayofuaIUF16q6PgHtyAAN1MxHj3+1Xd23paF
iJ+pcr4FXaZLTnnCUzK5EMFSiXa91a4FTUhsc0ee1djsCezVPVqCLmqt61yo
vpWBtN0y2FnQ8cAhZ8pzHPlLQbuYYu9GjoZOypZ5jvwgYlUDiq0tILbjxB5i
w0GuXa35akKeNrGSM5uDG0UiPes/wDN9oBbkcChJZc5/MJEWRTXOSCwy0+p+
VPc97OZXZNO+sKhiNA/baLHAzR8wj1/4K8gNP/wS6n1AVS/SzObIdActxeLw
ZzP0bsToOdiXRO8/s+9BDiVfjKXF8HU4AM6DSZ3TtoZV8Msd4EtxVj/dq1QT
BAhhEpufmnOwvO1YYQ1BSvJfZLb0tRW+iP862py33Wyvyz80g9CGGqRZjsn2
9n5AepfxRqjTxb8eOCqfIvGwlSsIoY1PdF8smThNrv2FKm4QRix5MCgZye8D
KTTRRXwEhMKOeNEiZdpJVEU9PqTidDnkK50oetZ774HfGml5izkNCAkHPKlW
S+j1FnkBtPa86BY+zxCwkixWWjXlUDUjyZqcx1t9c/C+JWMtkqHiwR5E3JPY
VRyihHzU9nqdCJUQjJH/YHFFI/a3YFPr9PdX0fNjoStkhrJAdevkUPkoVkYK
zqknKd65adjvlTaxMZKoRIDU9UTlRoCiGPe5LexsRO4svE9Z/5lpJdmTFIf6
mBT1kzT5+FiCNaGwk+5swdVY3AfEWESXjuq959YCVvazg1puPuDn+6OhzOEA
9WTdsWhiFqr8GC67ncrQwIUWGLKZXq+L/L35Pye2/u0HN09reEZbsSo+oB0O
JNWcQp7hXGKJTtaG4ryjJH1tipy7plBPbxsb+r8fgRj+IB/tIgEZSM87xx5c
2nJxjANEnHHSSwUrcXxc2rLbxLi8xU95+afQffzj74eAOP7HM3O9gvV2OsPZ
Jn4UFnnu9Z75/F1085KSkuZ0Vx/MDL3Lx9HYxh8fqt4YmtbUs8JvHCrTipts
y78zUyvh5DElV7qU+97R4veeuQGhL9QyKAYwavHAc2tvrs9Vm00NMy120xi7
GYZ2L8JtKg9Yem4IonREqlmjWDuul+KIzPAOaFUWzVTEob5EP5Fi9NA2V1Su
R5kyT+VXdvRucw3hrkuv8B/uBC5frWr8JNIz+twsbmprr60P9Nk1fJgNdgOI
fV0Xd7vHy0HQp11iAP6pia4C2hmrtXB5RB/J6FhlMS6G1/jzxb5xWLok1QWi
i7iLwuho83T8N2lNXC2RoTHH8RejfOVkEahGP0Z7QANbcPzeUknuGnY8lRrH
7YPsDu0MzmxLRjz0KufCmR5Rl8mTMfrbW4Sur7JrSz4qV6V/BOaadesFZyx4
6LpunWJWma1nOLLK+oglWmwICsDD7n4Zwm6AtlYhVlBQJnfIO0mZdB60nghB
RMtRsjekGvdGU3pBaFulKcmPWoFv95d6eHnB04Azb/YWJaRbLKcSbsLuRN4W
kB5hMDWTqduNmr4FUrccagG72tjd2X9xjQQFMIOykbA/EFdUe28p/6jRlZve
DCwc6pUVKAvFJAWGARIaEfMVLx1XXnS6CyljK/SAwRyn4W8yc9mehMFKmxLY
SOVt96vt6IgmBXl66gFiwi+i3H18RNLAoAA1tqdoKygNfuCShBWmr2BX4jML
oDc/irtZPwmZFg42vW5Wzlcask9nIzO3SAub/D8TbrYcJWp8+qnk37ijq57E
7eogDV7ihxDpMegYne915h9O1XgYtbxKtE7GWxg36Ssx3deqIVgx0UTK9s84
qvGEuUEBso33hT/gUPBZ08dOUmtepUpaV6alNY3FCkFrMpUOaQYx0fFaKhNx
apW07CMmEglNVZAk7ZtcqSJwwvPurA9fMfuMSuHoMvrd5OzuGBEqcwrbIT9+
wD0IrJCV9a2F7cYVTCYp2hOG5aHzJOUin/rGveue2YrEASxnTxqE4iUML/1p
yAP1ibvsIVIR33tTfCztbjZhm+6M52hPpL8GeGd+fpWmhU0/iTh5RzVJm64n
BdBr+niRlHl0JDKUx0y9AKSXCUBdCIr6IebODanmMVtMDa5p39w+jAPWsFz+
4BTRjPDnDOkVvW8xc3d5fBaxVfUrjaKRoLty7nXqWchsFT1JHzX2SFOfhNHD
48B2V0b6RIgr57l2DU+lcCRtV2pAGbW+9O5GCQg+P3COrVbvv295J9DDKdYK
6eWS4QzfgFD+I9DCnrBKH1IKWV3qU1ubPOPqB+YMyL5cG8rGPxKXrDKyrh/7
Hv28A35dAs3RLnlh/HRCFB5VotLd9cQbaxHMrQX3xlEMTj+xUVFN1qoyIKTs
cKqLNOfc6yhXSi5Edrvga/Y8CF0eDRByp4jqwNiSdQB7TJcH+yi1E+yYsSua
TZX1i2vJlHmCQ00Yu2n/WshF+jr9ieTm+CyYAqpcokxhhDOF7H6iFq5fYSiw
SYwgdouLDJpai9LqR4QBcWWtxEipwb3wwVcQKcsS5Ck451TR1n9oAbqnKr6i
ZhrAqCf57jerb/ULdUNjrnBR3nkA8/RGO6hobFV+b/pPRjkSfKCjjxDpwB2K
6e7ms2utm4ZotNRq9JNwK4jl4rIpVb9Y4/oyornK0LB/ifwwzCp2Lk5u9yfg
PuTcAmgiAWpmdA5PDGM3ryAHupP4/Yvv6Pnzk8pJ4ahcU9kraDS3LOz7LlA9
yeq5uq/HerLUMJyyqJqyoO51faUsmKoOHtw5J6g9fGx69W6sHgEux+S+trS1
WbB0oDGfGcF48PZIJwhXCSjNJdHr6kcAshfvnmEXMRzsWXJoF9jXOEKDXtJI
iqwbv2jAqNQdu0h0p1q8HQKXxeDWPoIcDCkBXwXJtgaIoI8gbgHOswQPl0kN
DWHWnGvmfuMcoN+tLk6x5SOfCwdH6mpxmdQztBG/Me1aJZfi+j4uRSrBKXrW
1HSzYqckxaFXx8W3QKvFR6fp/J6qA6m+TPEslnoJr8jcFpeh7D7KVp+1jH5m
CS+uuuYbsBhicW5DGtdYwhnK2ePBuuHSwkByaLnsKkjpLN4zWWKRCnA94JmQ
HNeWzlYbyxpSILmIuDfUfiWmGNv1lQ1ANKpPCWt0a6rc4iWM8rGSgNtF47J6
gNajH+s1yhnr3rI36jnloVfafzLDGHQPj7gy/ub0jtouvSkJILsAU2TZDqLj
pt6umtSUozbJExDsRkBm2z27mBFWMpexVuJfVsenSkGby+T6IOd4eOK1Q0ve
f7ciD/WSVc03tnsIaJAhmaEK09mZmNmS0bDlgm9nCOfsiHPJkQrG9W3z+V90
lE3mt1i+qF8r0wNxmvUp7kF3pH9hhrxTpeVPB4M7ZWOTMwyGSaL2h5afae6H
Ke3N1lunqZROg8pK1cNNiCQXDeVz63ciVcaOKk52fjmYkWSuuXOVbSWa79+R
7N5D8Zn39KrNzx9PmthZRMoIPLR7QiMlir9nSIPqaW3ptxmuM2T0U5gm2c7V
8qtuOa8HF/UxO9COzIEhiGGN4OFzYGOVdkhmSaD0TRXIhJGIfphv9IJfUkzF
3vk8aMEoaZAbfU+d1k8wOgcC1KL12tU0t9ZAbevdB0namtFLCTyQ04fyi5eX
OHCBmbooNtlxOGxSQr6FiMx+7bZ2yug5PlzT+UuTf/loV16bjnfOrYMKSdKW
pHGpNfvWb99eK9tgpOQqazC7jFxUot8BM8GtA0Xh2qMECm3hSYlldUmW5NqC
DQagE1Y8tZQ4idxEVqptpPW2Jrhorwer6ZyFkr7AA2jEM5esCuQkLZueCFWb
KKQRh25+jU1kQb9TAkxI9qk6IvN+tbgKeBTd6xtIX++hisO0DtScWgshGyvC
bY5HpgmwHge6DX3aVF5FU3uD6565x3MXOz4ko7sJP/8gjKB/xEGCpjb5tJwr
IrTzEwWis+XqP950WaRrWRjNDqVQ1eR7tSfbiAM0oJSCRhMDnqC/wFWiE/MC
DUZfI3CKW0cpUEB8YyYRxwhE0FsiCO8IDKBJyalCQQBwqpFQkQBr5le2je3d
9LwBdQmlPNgtQtKMQE/JsgWLv2MI5uGlvSG42JtuzoYACW/i0Y8qpmf8ZtZi
sGF5ZA8XJ0HnkZ8cAS137KB6LOA5M3IWTVu/iXVusevWsNiZuMA1Y0McAe5t
3xW6FiKWpr9hM8bFf/XNBp6eXbmlWPx15zETDlvVekVNFx6YXoAaoR6+sOV8
zQnT/jQ/OX7GVvrLSbcPkMMm934KQA22SuLdEgR/Zn/vO6F2R9I1ohnKT30e
cPvXbt6/kXgq3Bpwo4+uW8ZdkfY4s1SdOdu0KVS9BkmznkWQW8qoYkmAkLXv
b0BA7jaTgointImIG9cT9PnTdGwcdbZwp3sHeH/NmeV7SN8DKIOLsDI/y1hD
4B8+Me2byaKzqxttLg/z6ViZw/S2kA4SpMrYBspSJv3FyQvNEZ9PXIWzCRR6
daa71eZv1MwVeFxYm1lwcPFlIqZL0fy/eUd7eHKG2qY9mXASh4oYHv3USzcd
OVM3F2278FYBGTvj5JaG7XuKnXQbjtR9Kiaz4inmOJfz9CfwfxG0qlV5zFHV
baVH5vvzgNaVQyXYUmMLSQ8Dfot24YmZehYFPiGr94zygyRqEnFj0nofdgUL
k1FVWhBeNQBmfPlKsuBFJ7vnpno40I40VR3FV1LX+cz89bDJGcYDmpaW9TPl
ygwuSoc1/m6yjMo+X9png9BZbSpEF/aKS7MrxEE694A8A4aDTr+AfyLSUXgN
SGARbkno63Pb09TfDm5CokJ3fVjZ/S1nEFLHSkx1GdPjSXnIQvDgrA8qYG2B
U9RhbkHGZfriePN11YKs2522wBzi6IPN3nt9+znnUxVYd4AYtMIs3falRcRK
GDZibLUDVszdP7dlgt93oCM3HUaySXXOuYNPIIa0NlWgCdnRF/ylWS/W0pA3
2me7H2AkDfkLOsjrNxP8wS11X3quC+G7vAWymkDAyBT466/eb18pIdqCAZk2
L20qhTj3iulrejwMGsT8vfXBRlu+Mmx4pRRXmMs4nUdJ1rKoPZfMfYO+xPfd
i7TCcsfRwCtwsIqgxqBudreG4SUBk2BvFQo8jQDKnTWCB88MN6TVAZRMlkz9
5QiCuhu/phUNHxVo4Oecj77iBA43L9qDzQR1sfb7CuB9Ww5hyEszJTrbALTI
moGtELaX7QZU+FYl1EKuXt+l9EH9MXOqszQmEWIOT1c6OKfXerJCIL4TJKSk
g4FBMy3LmKyDMaa9BMWIJdIcGne1fN3GW/LlyhMZtgJxe1D2PpYj5uf17L/b
J0cwgG91vpNKk1aIEelEh4Q9EbCAgKJBmBB6YanSqFCI1d2dXy44dffOYqvP
R35FHFueut/SvBxlhzVSNZOLORJASKmwAArICR6SqStU6nQ+d1IkP1SMa9wX
JHfoBnm0+RvMRg7JNWLg9493CBhEMcc0V60aiq0RndslTTKZxHELeb8nyJvK
EBqNnfJFX9RHwRmBTebM56HmYZBtaxF+zcb9LkAsCtNAsvUOg3vtm5ywQuVt
eYNDORY05cXD+r5B1GmKe5YtV0fkI8sieqWfNM4Ym4xWfT6jCYBXDnbqvu/6
40EGDZsveY+6V0qQ0hpCJFlboEZPjgm5wu9+Yef/r662+yFv9cj5Bz5fReiH
EmkI/EOlmX+Jy75moVKW4ZNcDrSHsKKNagS6NDY3Xdl42LGDgH4v3C/vXpkL
11SK3ZkzFkODWDWTzzARbUXDQxDnPh1DvuO5T5/errqOBJdI1f92eUsXVpjk
BK7dBBUNZo6/q/1OgUvWODlKOOQ3uws7QnwD8vT1AU9gRiKy00c6WFItvIwN
ai8wcMt2gGsxef7FKlhO8wGjKBh+zagC1+hgFr4H/X+fAr1gOt4ut2TAmuZu
DYgvpfZH9q4QVmOfHGGXyMibUnltbSGq/WJDfvPEhpYfYOoq2VJQRyuL56M/
m1PFhn9SvcXAr96I5zrajEIcvcBTF5N8Xe+5KNq8rPZlXf20cq50m6+6qKym
ZD/ru+XFbBu30iES4J04qrFsJ7ViEDhcoLmSFrBS5hZG8sgrkdglJax8t7qj
9Crs6gGfP2ofK4gTT/138s88sfJe7NpfOKBjeG/t6ZcwGMBjPdZDj4+cm6vH
ah7p/e1Ko01cqq0H48hQ0pjrNwOSkeyP+I/eNVPnQ8kTU5Xs7yZ5XGFUicOf
ivAsXeEgQdFql73Ywaosr98p0G1Ag2fWIcQvN1ptPG9PIsMNjRoiFXDAVntq
VItIjeLl+VSa22GceC2eBbDotrT8ARmNYYlqMoevWI9WdcXRBqkjp7XBzPGh
4D0rp/PbpiaQmSqfE4vRTBeiR9yoo/n5txeCi2NuxUqsgF9AznQHl9nm6J9H
vXLxLbCx7gh/dexjK35PmnoRs05b6rCvpxgh4z44shseSde1u2iA4GQK2dnY
t9K33pLOZ/J3YxUQPrurrnwftz7GF5QjhNIU38QR1qk5U+aojMOtu+/Z9Zsr
wMHTtxpNgTbI+Cm4vsDOkRqeZuyRiGHW0VSRkY5GlZoV3CVkCS30BboEOmd2
ruxlmYtF76Zx+fN8p4UfPmzVPV3HTqpbOYnee4PjNctz6ihcMr3FRZleyavG
GqfMKOUnlnd2AJMBLhjJg5sIObpvwyaFtZ3bnoh+FCRtZl2A/6bvsUxVdyIf
FJ7u8lqxkxYkX/ivF+swc5GUl7MRCmblz93mwI5dEATqkDjWG7UaDFWp4aWi
2JBiRqrpFzi8YFpkdwNrxEp1wyuDbnZe6WmxxbVKxr5W0FlMcGJaaGziKsBk
b4jKlxL6SCQkrsZgZyohFuzqdqvI08ztM6rmufkDlmXxLOMaHj4vWSwWhGme
Tz1W/om8hHTs5SN2BfMO9d0YSUmhZSpFiTLytScBz0c34MeTRneUwsGUNTHW
3ieGB8m5jUWC8v5nosc1EnlWv3liNRSrwAyZFyCYpaOh2TrMZtQlRjnMf4OB
JyXfNCPjub+Nz1o33LhUD5zVhup+nGfuIGrowTtxGenGpy6+TRhB3eCYWFjT
4b+PGXdoB0yMaXHcURY7yYUQZOrabpZouIDITeV4YnWyr26qzSKg0j1RYqxm
TANJLeo6LOnBCdDu1aQ4unVukLpHRioiBVD4z1doHjzi9vOEwz0SMaJANX+/
EPgwF0IOpyMkPOdk1bmGGl3qCPBsCmqt2QWxvjTxZPmkgB0LY14kRwkvJuw3
hcYy1L9aKFI3H1vsGA2dks7Y215CBjXS5xRKS0pMpMAFIWPuzKLb3pa/m4C1
fpJzXdaIHiIfqbgvV+rnQWoyUjJQc4IKq5K2UCtqjvJ3Vtq/JGKx8EE6mkGH
Csb6rNBOYXkuomQmreWfCsTHDsApx7Zjgge4UXjfZoWuGbQLMpRgDI1760nm
/RFm765ZFhsFNEc7oIH/xTj5FyQc+gchxHloImlKv21fHsWVxOelOJ0jGluT
TNL41mvABi9fr4CVMQ2qcATltybZC30IYUx7J4klFKiufyv0sL+QAbOZ0TfK
OyCHU3fphVRxuVIbFW7f9T3rDvFNwkN9+gk9sLRItmQtKJSNRQbES0rpWxMc
IBC39DlCEFabY3lod3MaRf7LL2qHm5YGn/7Gt2yM9zAVFMm1JZOWlBTAeQXK
lUjx2ME/7UGaG+1M6SGTN05tmgANNTneRkzddxqBg+5EJE0W1SxYnxUtq1f3
N3uzBkowWdOiUxKE3Mw4NS7+9fpGj2BivU4GJFoObWOW43hXXNOQiKKo+ifF
SFQaI6TYiUrLFKt1kRJ4Xgb2owHrKh2soPquNQxaiqVPLZgDpI0adPtnhy8G
f9vN9hRNWZXkNlw/8UtbihWO96xD4YUDTkHHGzn2o4L/V6LR66L0BkXSPMiI
YmNLoTQcklv2DN3yqL7nJtSnSz+1AG2tMfDpY5Kz2F3rDY9HbjzlylHx2cat
smHH6V1ERXyPEU0Md++JvQi1Gbng+YLTzqG1VZjywRkzlmiLL0KVXigSu8o8
JZH2hLmppDjh2knSncXd/82N3j/sSUyOAL3+0ki/2NGAnpQndWNpUBb+Pug1
/bmxz6uklha54n9sDi4i/eu67P6mLWK+naPzsOD4vjaC7Can8l8Fhwz0lbL5
GiPx83UhT3g50CdziTF8KvYLEjSGy6KfjFmEaUGwUgkeP4lWU20tp+ni4A3Z
5uaz/pO8UBaSzDMuPFv9e2KQZhWvD0lUwlCBmYFEhJPIBbDJJvtLsYJmPnnI
/bXcOrVrlvHz3fTa/5k3QG2xF4Sodw6fqbywpxVNAyc13psx1XvBCqT4R/lb
FIqUGYE77jhF9+nOQSNpyLhtn61E/PD7jVVsewzfvOEI1nsJzb+7f0rOF/T8
4vsO7gTPz/wH0ciwcg1do5ohezICZKumKNms24VQE9CCJ5JsLfR+0npXbPw6
nkO/UAOoHsf8ztmQmC6MEHTg/09D79dFr0CZ3gO5ZHZqaktQtNv5+LmGOnph
t20OOUdQDmeFnpnnI/+4JC5u0vmqXBswH75ekHsXJlMATkO4jHI5Se3nFXAY
5Hj4kAuQNe98wy0WmGAN3MmoGJRXm1WQzFRrpde22S+x78Sw55thqP51bIZ2
P1hVdWwrKgfhSAoUlDNRquJ+kWlV8bnQtFh0d9wlzNoaVMMCXHLh5d++3ook
IAbf8ulAnocmKBSwGdD3FUMt7CkZb4CoGl/V1afFmtvkCzD2sSb9UlAPRmX9
TjQPGDiOY5GWfHV32l2s6Fy3DzLb5kHgn9cOY9hvuJrpF/v2x85k3Cq3ReVo
6j3Qo/jlGjtzoP3q8t+Qk32TJR0I+aX+ptoqj7UUypmPvAnv9YPgfup/xmbc
jYVn653ctPWp1tYrZcnOeH9zriY3S2lO21w+X2sRGWNxlnjMFaoM6z6csXss
XLudg9wFF4eNZNiiUjg0tLJwBQOLHPEcVPzKcCLf2gYT8p3XCIoLCT9iJqiv
K03JAZ7SAmhOxLPJBIkCkxCMPX0Un1Rw5XtWHpBx18zwX/+95s65DhFCMGTp
V4I9hz8c1zGxi/VgSV1SHuGDnVIun05QlhBFjdueQ+kozTCjyJRRSFWw6q3x
t1RvsUde20f97ifY7pctkj8XJSuS6HkI2iN/XJzQ4AWBT+eyXTYLBkSyr8m8
+l836Luf69Tg/Bv98/38wrV2Y6nGaWiWnjwjcCHPktk7NnIRk+XpERmcLQAI
JJLpNiJGTW2rG6v3b1pqyhmWjHQcL/P8GQ10LekCmOY3FlMryZAhjSCuoeTj
Qu6pRf9gNwHyuxQUmYihvcdVGvmycnX4GwB9bFa7x3oaA4+jGOKPT76uSCCE
t4oevbCdXq1MyXXuP24jHunUFD6aguLvEnbnqC1kGfidwDMRb8vsxvcTf+gz
sDCvd3utV0Jpz5lQt2A5UOeOcUe5BEmYgC7hdwJXLv+ZcSPmGmKN+tHn4/pK
9EGsr+/xv0Sm0iNhnxIhiwyXDieoQRd/AcA8JqOE8wfArFfliO3hjflIOdWL
5X8uJ/its5Ok3RYPTD9uKtlGqUv4Q2CWzjRB2WKgTsRHpPXY0O91Idvpfm79
XMUcVqiWjFAmCyjDjVX3nZTCF+nB2Ohu8O2y2huldBDMIVz7Ln83MT3lUi8a
VoRk84GpoqJ9jL8t9MbNz9sAU17c+YyUQ+66XVO5XPbVq3YXAdJXT56cBuzP
S/ub6+ykhbyx2CxP/rLoh2JpIr6qbW16N5QCFGht6iRu37tGMKhnoABfV4CU
6IAF9xQJx6gNn30NfXIuuYM1OZDxSKpG/prigt6y1PgjhlGGSNEFtz6TGEOD
Y52p6t1tqHfUvp6JRE2VXBn6zfRykFFbDKjPUJjOgVtcRjqa5AOdttUFDnOO
ddFVuyUkQyzbi4Mn5YdYeBMJ27lAfuAx8Z8KXkW6B9YF9u2yqHgUGIebmLzP
/3jfnmYzNTp5ocVJe58bH7LPCePTCz7jJOAsnWhimIYcNbChVose5tunlGZX
tvrF+WyzFRqYpdnC4EfoCEjLC/alg9R/nSbYtLlIe6rj7n9cxmrRrjYvccvv
orowM/f21ARehAcG5vb5e3tBS6k7pdGWIWjn/SZmYSRqVN/BbCUOjQnKk22U
pXTyt2jY5n3Bm5EMJPQL3SqsXrl4h58K0Atn9k5u4bmOvcp/2+xkNhsEFMWs
UFL9O94/VbkXyb19YPlHn5AHb4FCLvqVqsDMbSHwIEmCsGcRY7htnW4QEcdR
irjHAWrJmpWjYZpuQlnXyHZJ4c4cx+9FCIAXQHkOyLhRqZFYcU0JpDVXBfC7
mb8wi5rQtk7KJD4U28MFl2HFSOqXrFj78FKwu6toiedQ0T//DaY0h91cOk0p
8f59cKMa8le2W2oxyEyPZvEb9Yk+nI0HZbY2lgruWzhvF/Ly8eHQjTMVteyc
/On+kBBmw6u/fXCzlTwG76Pta0iU6ecXJasVjq7jLBuzasSbE14JrDGcEVue
7bHxa+K8Rdx8HkhP3rCILg8TvbXIXRk38F4gvenVYmRjJYaDIoTuPrlYzR5Z
ahoV0KBPoBcVlMRy7bCYJNTgh1mwTVRakcCjOXESbgHP608tjdwGL6EjX1zj
QP93m5I0i/tsZyny4yvg6jD3FPfoJ5pmEPYt9JyWLqZYL4iNGvKwtvCd5APY
PPLibs8lQYZarF4uSWyPqs4m2B1F8wKqCGKCGwIp1oxztDRlt+5JsIi7tshs
DvQGU633g0pba85mzw5AyeWjzGOnrSQteZas+21NeH0hg+BEfUTw/KHqC3/E
Vx4+N1CLPte/+dPsbzv/hjCHMId9uq+l/d146so0bN/cdpn92GtheQ+4nCzj
ZCRirvO5L7OeculqzVQNa9OGAO5fKxTwdUAn+SSmaKQF6UZYftQ+z2idP42y
u6BtTVgwrjDOnwLUa86sJQNRFbeEzXphIziLxTIOu3F0wTfvYEpPn+6RRKd7
Q4RwjobZOqIsB8pf5zsTSnZOCcdWbyCcb6b4omrg/NSVdZSx7iSSyxHx/a8v
knjrjMC3mW2saYHu37C6z3Qvs8iKTd8sBu0OPvrbUroPhcXg1pHrxkRVdcMZ
l6mp9LGkfHaEoGEeP5sV0vIExFpcJ4xwj1sX0MiCytkn1qJKNdy2bVuOqHDq
1QlM+WXKSifYhO+VY2Qhgm5PWAXTGeXj3Ti57g8jbdEayG9kT08OiHYh3VRm
r8HNfD6CYFHvBV3VFfBg15LGONcU5rqvJY6xRZNIMpw8SaYL+ZBRazN8t6mC
9UB8oaIOVKlhvfPxeBwXkBf1s4IcakUYQEbcy7rb4b1sP2CH/e0FoU9n8U5V
l8YXTA+f8eRFtNcrUCHyuZ2UQFcKR5VCRYezwriBHid5FnsPM2FPGvfuKTMV
9psMFp3Bl7jxINCngt6mc44+zPqW2hsO+Frh+e51FWKblsTTF6NFsxnvy3cU
JfPAeQ31xKx0HfzhqNRK9I53k1hVZc8FzwsoOZU4R0jiDIF0+wPDCHJv4b4z
QeBx4BEmi1LAS6kPYRqgrGnVSlsxMX2tnZ8YVKvUp17c/VhIl7YAZj8nf3pt
/xdrOeSb49TSDkNFLIcDtU6e0wzqDo1dQcgJNu7QrovFOS9o8t+7ClKZ4rue
Gf7eJRhNl4L4lynDID0tYyvrHIawHDGiEoelTa+zgPMz3Rm7w7GVnOpg+0h2
p/4B5QO0asSSMVZpI2iS/Ei3QI+PZ2qTS+yqyLe+6/PfQH2SHZ1EGVOIQCfo
zDAR+MPeo5RS3X7+ZeRyt+Tl2rtEmH6wQALWib8uDPx+242CyH9jKExgk9hL
7ru03CoSebCUDEC8lP9LkLvD4Xx27MMEjoY+Rf8wiu7LhkpeCO+aYgaG4Bdf
/w2M24RgWhe3TRdQhuGWPiCLDIZawm9tGL/cgVr67FWVe8zJGqOWj+fac8Kf
n71HJ242m3WE07ndUAVW0B+NDMpk04/vk+Sh+MSCtwsTaMHjxfV0kQ0wNhLB
Lb9qO/FHblWcsCRAHKPbJSmnPmqNbiiMNCSwJnmweGHDim6XzCuOSJ3M4Kkr
SET2ROtPkY5lGQch6UrBcvw+SBXFlOUscWQCcqJsiDmmwOt0GOKBoILDr5Vq
b+GdKEBMQIkE56YXsUoOjQv5FWDQdkKogwx3fnkBT7cqyhCLEDUegihUZtyE
a1IxcgEHR40n1IviS3AJCG5xUTTOoxZKl5PRCWO3irbK1+8qYQwlrXf/bDTY
Tq08g6Sw7OMUloKKaSx416C73whnkzpkFMN8QneBScPfcT9a/pbEluDs6nNi
KRakTE5hdjj+QGQozjb2AscdzUHgMAMbojgyKVWHqopKr00HA2AvnOJklPaT
X8kkp1iARL9426yFRNATxVcC7+i4cbX1H3zbaHbAT/Ae09VLxHC+Z9dQZ/ks
BcPiv8DB9NasGU7Dh2LP29nla2GvsBtltDQ59P7og8S2O8rm4w0h4VC23Wqs
15LAwoS5MQXhhCny4FABpi5CqGxL9Ve2JP3iLOAAlM0+Nu3MZySTifOcPgbL
rl9/wfH32vuU9+4jF5TORbyYnnFzkxx5eoBwtIjKvKo4S5GuKv7zNber0qK9
T6+88dKA9m5aOUGKw2OtAc4M3EVLD+HtY7RK9GYvM415cB8hEdeHz65c+OtN
P8qkWQFZ7Uw8tZ5Cuqz/S2h3h1sMSgt0+972hM/f8wRTWybF0c05VTFP9rf+
scQ111rZpa1GsG6DDqkgS44+M17Fo7LFkx24HKWU+3Ip2xonLY2sFiK5Qcrd
xJQRV9rzljpE0Lu5zKelENcH/qEKTZB9BhyG0B2pnVq3l0DMcnARKrmtOpdr
BpvAiVfd+iwo3hxcr1WytMyOqewePCprezlaq6FXlGvhBVUmfoTQVOr3A1n8
eVfAiZuC/VQHxBAHbtXyXbaaVKexyfQ5x4KtWe7jBw4CvGx5Pyd2D205359D
8L3jMj6HqM3L4UsTrVHCcDOyYD2DvB3iHcnHDVii03nX6E9gb4VuV0nzCct3
sbU9LTcb11zHBgthvNaQqoCnMFLQvwLnam4ALfsH4WeZW1OzsVPtPj6Fd4ga
KxE9jJVuvrTEFSFeOotI6AbziotStDmDuOqdlc3BZlpM/kvYImizm0FyUKnh
WkMEzp9XY3cM9IPHVg92fEI5zYVdK5p0/xaZHXdVhCqlhsCDbmLkLCM6S+SA
Fteg49TyySgRoYJ1HidDquFat/vexZlB0SIz5EiUMl//rA4OPy1GbweeTjAs
oF+LE76ZaF+LNKSRc4U4nCOkSyEyHm0DukgHnQEfgsK1vr+fjONpWNyiSqiI
xBpHtiRo7KMQi76zjkshebXGhCvFcjgw7tFO9zOTO/pWiOJSUdkHw4K9tkS2
Jp1Oi4uA/fcKti6+Mu+lGhU2GG+ERBrmOjBncmniZExjKTaq3t+nT/oSCPLH
abjOuatxFFPcOIvm4RYyH4PaLjSRlmupSmxu2S/O/l69XPRqDqdIc0b7srNY
u1sZNZQmKEoo0KlYdW1O04AKygRVboPgMInzIdmlF/2pMCyfisJ8NaIpg9S3
pOWNyFARYmGYVVgGKNdshI4J2iM9OHWWiF5adfdQQiEQ+TkBloBpTe6o0/ZU
5byt7md9gPl391s2Anrfzg/oXQ3ZWyvUtU5Aj5Ihk0MFLC66r+pYLNJqjnOy
zzZj/PXxfHv1bq5o7w04AI1k61zNqU8r+fXHzfb3VgZSmQRYr2BUzZovGPxu
cTq7+aJrI0LWlcniq6vPoOQPgs1rCKY0xq+mK7m/YSPcLbv0eqtTpJW4T8z3
8l4nSacICC1hLXd87dlLmoZqY7A5l2T3UmVdG3qTn81QjEfYxrhyJf1WwH3f
RSRu/rYgld06GTlOlZ47Mz1gVnJ2gny4b+ZvShPUHD/b+yHpfDY3AM1v75Ps
aBq+LW1jzQ4cqi/wmyVAFlwkhlcj84yMUxhqQ1z1r4kedPJuahBftEJP7kDV
peNrwtLJe0lo/rD9BHmKsG773JhBIDiAIP9VScidtlvCsPxweWXtP6zURZKG
f79ZaYXRmGB6YyYPck5hfWvzIk3WZBS8ir/646wbQ1EGP2CfnhnvMxu++tpC
PgKJUXAIImKnTmx+lBSCnqJdXIV4P4O7PdnaWQKiozmfpHpRnJNT1NtAsh3j
eXZ5G2uKDQbLzHn8iZdVKzhUWEcOOtMXo3NIVrKsMNOUf2N9vCl24WKLoKSr
zaEI0uBj08yFcM037raq8QXg3J0l77+u1lV2z4LlAuV6e95phO91VjBAkoq3
wnQoOvJVOLqyRynRPO/wmijFwN0HPugqKUJdAtIEvJtdhsK/ekozucQlgeKX
0K/1r+SIInjBcL2t0PuFv45NEB30sajR7mSSU+F+2YPI2nvb+CJ5h++ihLj7
oBoRPkvXcTYaacZk1QQgp2Ien4e+a4ehTn7SjjyGA5Elj9ksfV+1rSIIONsr
8EzIGG+OB27r5MQoCgZBl0vNpf8laZEA0ApCTrgNDD9bTolMBCPHb9sXQivZ
32av+69qqPGMObJ6iVk26D77hsqOMTxPOQ2LHCkPPGRMMkKqbeMI27kG2Nj2
Jb0RHaDawr+3/dkH1m3XZ9Lkv7SCTeO9aRfjSg/oWnZ3DkTZT2dZEw2Gi4Qu
OF2TwciHO1WuBK/us1g8RtUm3sPaw35GFAgMtVUj/Tf6Ha6w/PWOd7P6x4eq
5NDhu8i9rFKtDwWq1D11+5Wbu4dd1ym6jvtYSDLVLevW/4S05tilQeYcaU0t
LoLZ3rTntWBwymu7PJwUBvy5nWOWpK/mUKMsMEOa6fgQlOsIfOZboSJHiN9l
sHa1mJIek7Z5ozxnQUPcm+pkFRRN9PswOCYFkhvI0KgzjQFYR1Oj2DAVeRp5
bDAJDT0cN773trc6BcjrW1VXNic+8VYuYvKUXT6Th99p4YZamttiBYSsGuoo
DTVTPeANeTUAOS4g/ZTR/0HeubW4vcvPg/V9vkZd98rjMVYIZnrTj3gBCbvR
llIVwgsFPligaCLwK/qSrSbDgcM6EgTFUg25K7LGnyn8JAqRP/7JbFY+vZ6q
gt8XugMxrPW4yU6LR+TYsIk29bVarMgivA29VhRI7BqqcDUqOlXDQmyyQ40x
9IVJ/SOj4F5GXz6WxulKzXTuDGDH9ew3F1+9KO1zFwEWBe7rXw1Qd8RMsXil
7yGiaBi6CSzEKivJzboMC41KoyrpQXZjBH7WdMkIKb05o0m1b/Z+t0tSEFkN
zFv9B1j331bVmdAqMXSBcpIU9x4KaAEc3F9m+VnmqfmfLb57alfcDPt7RiVm
Vt+07qm7GaaprUxokOWjqJNiKn0WOXfUu7h+xwUGM8sLyImWysrZiQdOhtzk
lCE7lnn3rMl9VGvuUmFXLaQToa/9xpRFR4JCzQZKZjPmwC8XZRyKUUTQB0gg
RPJtlkFsSFuieGoVe9acuWA+TMXg2VtNpND9rDjE8gJUR472TRl5ZbvWd+Uh
0OOgk8jcn16SVVvCskThL0FJ+e7rY/7tCFvdwHa4uoUm6yWIV+r80VMk6lOR
7K5XgU3Q+wwmKFW3JtzPj7G9ojrGqhVWPi0l2MAUojLCqeTE995YZtc+yWMS
CxJJnIMNf1Q9GO4n78KNrq/ch8KYhb+50swFmh/Uo2suiwioFGrkytUsdZw+
HScPlg0N/J9M/+PI4BP3otflytJfGoFS+RqRFPeIqRoBhFN8sSvxvfLMgKYv
Flf82hvrlOy7au1k5jFQjCgakqG9s40k9nMHBuvQA0rFdlR7wiXZ50cfwJSB
8D3ovAvU+Mi06aX3/9YsmRpIJfIsHQsP5ScIRytb2kIq0wLztNNVvuUOYzQv
5OzbQ8xf/W7kRY09Y8XCE9AnpEKsOvdCEfLzEsvkajd3ZKahYKvsChsz2D2n
q68jSdUDQHMJy/wK4IQfsX4hZXh/1aRkJ2D/y70y12ZB3tUfc3zdoKXDFCvQ
aEv4GSGW0vfoXTWf3uOkIx9lTCthYwQvbb3Gs+Z4xtq7LLgchGigyFu350Bi
PxGFyUabRIKIr/VtF6+0pWmGnXdRhb4WPKZiFUUolbh7uVFv0WpyGjgTPUju
c6EC5Rwy7Ax/DfxyySeG0kcZVtsPNbHV1ehWFFIR/qc3akMlBkSMr9tHOQZt
ltBeOCn9GeUdqWbxqTxsXjUFuEYlcQUdRk/w6HLvyvhp2qdr4BzCx1QqO5Wa
jCQn5j+gju/qp2LS1+ruu5vd4EYtGU0hM0zWqgwz4mMJlQMzTwIWKVRXvoVd
CINTSfHtn/x1Nl6o+SY+zdagoFg+JcVep04QZmBSfkjRHNUKW96VhZpAncm2
IF+sB4sZQQMd5vGvDZeykakUnBdgn1K31CArqknLX02ceOADiSM+NlEaEZJE
oB59zdU7uiFdtTToHpeis3CkRrS3xIUhLFg9nFmyt9PxI0cMEh7cejzGc6xI
XQShV6d5V/mNxsHWFufu5wRpU5FhyEZlacOa1K0eYB7z3h7uhE49RvDRGlJm
iTEdM7lO/48yqMFmmc4Zpzo1C4u4lEv1/cnB7l4TykksZ/NJygfJLfFBTk38
YaPNLol2xfmXQUmjiQrHXIl05LUfEtiRdy4HJl2paXtMjU6GTbhuX8mcOHOW
ge3CFxyu/Q69MYPqMrvG9NDULUDj0elTc+7T5Ko9zRZEjXJYIrvAQ58TZFs4
O87flnTOAWKjJPH7nByz4CSDTBcABW9xIW27CDiJPH29fy6RQletu+4e5bIO
IRj6Q2b4JwzfbsAGuv+y/TfZc2T19DIw5VPy579335jTOKYGX9NdfsgYMOZG
ZggIj8SgX0YtNgmzChM1YT6zn2c1G/tixIxrChf4slPF2tYBzSn6g32Y3uho
09aify9ogPgDI3tLNxd37zdZ76gByNaCAMzQGent38sPEY/t9ITDm+Cj1Jq0
StuFF/L+yP07LPU9J9BVtltB9JxNMskOH41+0Uor214183eK6x2KmlmKX62C
0zyuKoN3UugsJfGS+c5oJsncaJEkPYhxeXGe13X83LXW+GiECNjguaEkK1/E
1tSwelrJwoLicMAHJd3YSH1gmJKCPcZGciBXAVVcSk+IL8MA8bnuJ7Jq0uEO
NhiNEb3a/K/3Hb/cNJPRiqevD+Qe20Trdamuex/PKCU0TGwhRDK1jgBF7iIB
P32H0km7pNtqNjB00BQdXNoUwGvrMdlxluWNQ8j44zmTEdxgcboxrlZ/zjpA
J0MNGImKesZ0gmqVbBmjor5Kf5v/UZASifGvxitMg34V+DmthGt5dADFx8ie
L6BA3h68vVqnlN+JSH8/UiIbR9Xm8RlwKrDLNcoCyV6wZX9L/gKElRl+ZgH7
QJo9RW1MZ63yXhHqNpQh/fYMxRZbXCZ0tnNcVuAVlc59iN2d0GCWdLnoyN6C
O7gZAtn8tX0s14ipXLhusCzYGoGcqs6BNb8dfoXzMrigEzRfXuFBQlaA5mkB
GncC4EDrZqzLCSoDH8qZyqYNhrk5hcJLG/fcGqfyMysZmN64oa/N64xF3Hyq
UZJo3YDBsm825zO5npoasf/woNFY/vfuR4DUJyhfVISRSRASF/LVbJpWgh9v
rbXcuA/nOSchthLYrcu7Q1JjDVLJh3WmOLL7F2Y5+j/r06eTWF+8TqZws6iN
Nt0xS6cI+GKZIGb1UeJF7kxLSRK5OtYSp1EYXkC9Vq7GXximffCZqcvrMHJw
/9rIpV/XgFkHQ3iV8Zxj8jvKcENQhQN4TprISRe8lTvsMFZ8CK1/Q7CiwARk
0tHUPO/Rq+113CFBEMCPZCQ/6yQTOHIJhwPsoZY2pM6EapdDEF2CoH9hV8ED
uN54KZcFd/2RBXY+q9XmnOH07Ico5pVo9RSiiPqARVYcG6zk0+dhxmLop6Mu
fbABOeXU95Z6GsFtab4ScXz8fKv5PViB1I1fSjXsvoeYs2JeJO9j61ZrpDsl
FwEgebygagUy9NPaPiwiFTFyDmF8AFFBRX9ica7bU3pcm/hEFT0FMR+j4zpC
POhGre5VG1epf2KISNR6N0pKnoAtZJFb3vgP1Ozil8xZ42ND5P1WppWZFuBS
1rtyFTdjWi/PuPk1DIF/2Wiyfjer6h3R+R3zD0uVcNEbvCc8Cfsh1Ykiz94Y
kcMJ/ZLoRRxFqnfL6eSOrZlm10HRCMywEy6z8a62yDZLx/Nbjf8CYm3yUqrP
RAegZi/dor3KVuEK1/AQSewRHBX3YLW7kWPgBooYb/mvXf+LKfP3O4zxN8kl
npZ+qAgq/F3ULyrGULLg7z1O2dWxZk9YKGLG9FHYoKPS3r9GeBnm46Ui7ANX
erwi1R8IBDCbDYNN/bddCCQwANFvCGSSkz982i8MqFs/4pBsgJmcotpRsBDE
5zO+6Fw6F62RGne9KcmLVZNA2ah4+cX9ILr9xcRqDhAroLEO0zAgKOJPZrZR
SPqJaAg3Wot94LdploYCBvdkhvQN5JgCDfg8CR/AgvVXhk3ssX8X4ZoGz65I
canW3oqlSgCwcrmBXc9deScgB4gauF3gMFk8Lb8kAYehDJgZucv2rrFZjj3W
52fsio++o7xIwNpIJz8YZTEJUYlhrF50d1+klal+s6aKhelGyq7TphjKNbUl
hGX15ZlOcgzem9eynvflj2xkvg5KmkLFP+gvVne8TreQg41xHgDuLgzZxv6n
P+IrZ7ntQVQwet/qOk7+ukAmM7vGpVw/iNLefSHJIZW5QvJWu5Lhillc60oK
xGRIEPiYnTAVtjMo1odFB3TtFtG8DQC4dkPeH8xfAAJBK8ri8kLwJK6xfYfu
k76F1TheZ9nLr2XNAK+15HvCZ34U6QswLNrHD9MHsw4tVhszgFV09SlxqIyY
XI9m+eHEZM2e76J2aQD802G5Gkc36qKOWv5+13Ff3zdiXjwTa/dgxdzS7AXT
8dJ9h1cmSIsD1IYZFP57UI7wLg6XwDqE8MHTK7NS5Shdtzvh7ygpGeomOSgj
RNmoUa1jv8nEFVMI+GxDmpT8DVP+pimg4CRaJ2fIFNMB1X5hphGiMO8zhNY4
Gg7e3CMO/fsj4qzy7qI6jPJTDsm8grB471dViJkGbVOKBkQy7MHvnm1W72f8
lT2trGzScXW+vfIMzhpILQjMC6LQZsk9zM5lJjnsslzOWbFFNxV2nmN708oq
IIfBHRf3FsmTB2Y0bUkQ2gTOxntyj127J7oYiqQqHTFv5+2WF7o+kuWxRwIY
p1ryKeaCbqZJGKhvxN4gquBR/UGOKi1iWrg/mGM9/VowsHhFAjRtsIMpRfVQ
uvuPbSB2BbGgEQZ0glOOyobXlC36fb478wxOdFCBeFzvkPz0bBX4YtMQ/b1Z
kTOup633wPbAiIrZ3J8+kBov8hqFWRNbsIiyBozX03Zspc9mKbOKXY98P1Cf
/nj46QQCjFtrqlqPn+bkVCS8Vdo84dr3Es+bk7WJq+l7sGj8c7kHq0mKqEAT
4KVLXnH1pk48x/0C9lU+mRM75tZqpBI8RnH/bHnFxI8zq0uejQeNr1GBSiUF
UWdE8WlqEbpRVCMerzBjMKaXPQrLW2/j1BFYsKk+X8VF0uh2lSDpwWIr3YGp
2keYwbh3jIfvcmdwBLRcpqeyosCDZ9z4OWMO1VckYBdtaY4zRA/QK9mlqf5D
5d1bAA8JF9vzAibCnrpPQs3ChRhYSkqnE6YvNozHR2XmRG8CoYYGtJ1hw8Ro
odZjerJrku5nYpNcdZZKmgJ4bR+8Gy65j82m0SEB1OKd8ZRI0BZ6mDRqBA71
5AbvF65rKH/RE3wcuZh8MQrS/J8I5kU3aH0wgUy8ajyZJ3198sT9p3SpeQiB
Plzoypn1+vC9w+0coJsiEXkOzo2neNadkp6nhKbUdKfmDlUwRlvD9EyL42AG
JWWa19kIH86ER2lvXKqr/ppH1/OCGSKvrd92L/HDI+Abe8sY8LnzIOyfFYcG
OFcqFfxDnAtHSCKfvgNdMR7VOwn5KTP0dRlivwuZ8wXm5AIBM3xgyIy5+e/x
SglvPlLpVk27vi94VXZi/eI+9MVch8NCbX7bh7f38I+Ux0kEscMVsS5DE6qy
Wr9Z1V9cpK2//Vt08aUt3iVSFBFJhK4/EJsHplWoLdI4jXnhw29/lTcFk8OW
nPfNorjhzORqH7aMyjZIGjanF3hOrdu5DLp55Ky1FEgRLqRxcA7w/wLiW8ab
Ov3vsRuwdpW2Sam/bdedIWtnPNMyP2KU/e1uAt5Pt0xJKQ0vxtqXHYxXBsJn
SaI/RbDmtPHKQFQnicEPfYY+qEPbWmRNDbKI6drbVL3iiugfIWb7CQmgqEfD
AtuEVtp6iRUpkiJpPBmWHo4hos0USp2nbRIIpEjCaVwKEti5ZHlRT/BqlZ6v
ofhgKLGfTzkR74M/pg0A7ANrqXLO9dBVKWzqurZ7stRj4H/PbAAQ8SlL02ta
JBib4lY4N0exEvX96DYpw33ALhZfhXGUMg52Z8D+7UsrpfSHQ3EmEPGcp6lo
WM1nJCTmO/mVuoJ+PkUD4fmi/eplxdN3dbLGDnx5WWYE9uYmAm3ChDd6PUzu
tasz1/QyDtM6plxhvp9kW0vdLCdE5u/UfAfW+UG+Qe+22jea9XgHNxbqHoB1
V5JMs0B4Hc935VxFVuI6Kt0I8dJJOfTD1nbtGwvWWnzQe7wL8gYAknHyTK1D
2qHa/KZ7sifcWncfivql3xyPMsDZWutOJrAoiEQfcQUl4t8IloTygck8qjmB
eqCPuHgS1Nz43bJD0Lza1yz6OuRHY/1p4MzJ4NNJlaXrzPuy+I+ZCRlQEP5m
YyCISAibxNbVX16m8GarBhmVAtvi1/IbEU2lTA7FDPr0mQnKs7gpboYXr5l6
n8uILYpN1NjXB3f+8HeiTOG3Wdvf692NfIFVrsuztjoLFzR+KQ/+9P6cgig/
2GxUIjcARzKvXdCSgNwsQWgBd7Xrabk8yQ77yrkp60CZHiwhj78jSto3Pncr
6WgxIKrd+xvJuiExPCgHNBj799WD9bEqWNmzRsuy03boD2IfF7EJEYxSbR92
OvwrM9Xzdv64BQiaA8UVXJovNm2Hws/SXLpqp45v/SJHBfhz5c3rOqsDqvew
o29i5DlgNpO/UJqMVV+qsDsGagB/dxXbg7DgUUoII5MdCUJDWX9a8zIWrO6z
EHdEYwAPLG1dBD50S3iQDtEwiwqon/H53iAEwnTy9xleKYlPJfFtogc+0MwY
7HY+0AxeBjve1UmLwerJ9jmVQVHGJz7V5iBKad6W+yWiD4n3oEZmoNCvdigD
kbl4BPlNqxANk6rTlKOgY4/mubXT5TPmpC/jgpG6usarxuBSGJsT56e55Tju
V2yLB/yfhSHev94JHbXQFMiE8LTvA4SaJUgUSIH9wu7pWDL7V2P81aRiXoPH
/3EtRxROZZVNSm0VHK1eQVBWApQkCZqpu5V346DmHsjMyVxrSQxPPOvm1BeZ
HlbDouqKp4bFFCgELacqsofagjMsfYLK2VNB4j76WrRNaI0itWuIeQqBTqIH
rUBn/SKVWXcwLBMq73dVZhVwlCa5xxP+PFMVdzWXfkQ29Bl+Kk3N4Uevfdnt
1kDKsOr0lulT/esBObbvNlL5l0BT7znIjfh+cNj1VwUgGbOhef2xG1fx04TM
1o8EnkdvGwfBQTAoOmKmj6VMK0tGXZdKc0va92o9e2GnmAkM5WIWpQ1bhd72
ZLtIqpRWb1CrYWnuN4/+8yoIBI+2gfbD9jsnr5fHHCbLxdUJ7xfcghfeb4XJ
EHxcnqZcWlQh7OQmjRan9Ge/dY7kWvgr+5RtSdx/ArY8ZiSdCVf9b4JnKRJz
9DqwfOiLj3yB/CLYcVioP1djcNNtbKykQ8CWm4TV93QWYNadA/FxrUbHHz0R
+PLi0ALulrfKCoFWQQCoMVaYnUhPfrnj6oJCjNZ7GTahtgSyWi03oA9Dudx5
w7N8psk4ZV6yJKl8ckZOn1KslsEs+eBhwJRQNIH76MB6IP5weL+XnhEy5sD0
AdVmdLiywuvquez2bhsZ1tQx0td2ty0Dg2J8whf5uhf0r7fMySDu2bK2cLV+
cs0f5ak1OcFLQvXqdTWRoguzt/knA5qjbkvxo1DrZHHGgO2Nr+8C7hoYbcFe
ytMARHu35ZGzNJ6R/tMxbriyJWXXrY0gl0vLHj+F0GNBMZJnXMzn4f8OGJs/
fjRUVeAZZyt/32XxtBX66MyIKebKFrimxZEWl07WhRpXCOrIiL8B3JWW6K3i
MXAxP+pNcdF/NkAp0jTYXCHQjXDx5RaAccgP/7rhfYBYTn7cWEo8l13sa/MX
DDaWZmmY1flVJethheGOxddKSHCrhAugRWBga473wf8t6yasqCAOwENmEfdo
fAv9s4QkUHMFPNEj1iZbkRZ7qXLubFX5w5uqG/nt66c9joOLtADVh9rYsTNp
iuHJSxGJRBBZiSlCwOwlNq2hLksfYRZ3dZ/2Z37s0Z8QvaupCPKs9tAUc/2A
sTdKRjP8gwy+LPzJkaKoqvuWI82TNQRBUkrC+bg/a5AkUZ4Rqpuh2kC/HUV3
skwnnYytlchlFwiWQTGzsXhn4adpsJm914HPtNbLxB6uDbVQ+TvqakC0DiiG
eOT6ES9pJDcy5eJvRGb5FnjETY8RDrgTes2AJM+Dl24UiWCZ9r8vTTKPPd7Q
lonzI+HKTCIjHgKBxf1Rp6Fgij+fDEvYGG+Emre8cklWYIqt4m9EbNldE44g
tQUH40o23mDeCensySILd6hVVC2abUi5LVgyD0+MCr0zbvT88QU6+NKnAKrL
DwJdPUGrwSM6P4ktyEwsAJjZkhWsdXkH4kVrhCVJ8SXo9QBwqFO92Cgtj/iP
lWV+4qUvoVe1HGU1qiotc2b83wvWmDwa3oE/76U3Vkn9atYLg24LdijaAQCo
6Uuzgv+wHT1GJsXj5ZrLlvaoEyOwmRZrhZpQdai/BvRtoRUJ6pmoYJXRUdvL
pRbq/9EKLJvnmUeAzhwIGPX9YLtbp+9NaOiQ5x0AxWxo05FwK/uKFtRFQa5i
dkf7xumkiij2DivXDD1GMmIkuJz3G0sHhrj+xpIf7ps3Lapt46erhx1nh7aL
q/IMKDpvGyVAyhubX/9TlnxacYFQ181yv/pPudZpjONfyC4crzIi2ysgnux3
4b9uapLEq7uvHgq0j5T5I+GPGB+mTsaNqbFTBOKdNNgbxZ3P27jVXKtGjbFq
ofA9EehFYeRnemjON088d3Ksox0ozqNKk0bOnK0y4yNbciPqEPW3QDD5mSEX
dvu263wGd2a7TKJnZoezNjLnpOV0d/TygBzp5YMhRoL1rpJfOF0afK0Drt5n
HF9SjrMPgfdzFKP1mQJLQpq8Y6P0amSYb2KVSKWOkphqJbvzQjnLTI8A3jf8
IVO0EJFn6YrCYO12Dv3hi3XAbC3kvlYlsFcYj0N42+bdzEGc4jPIXo3VJDQH
ol9yb9o44RZzpoY+05gnh2Uvqp/m6L8Q70jNdVyZgwfAD8Jox+k6NRM8pTYh
xaq5aLjjMwmYiDqvy8eYewLZxR0oygTTPvZdxZmApIzEqXAnpV2P5btumjV/
+78Wys5AVveEOIoebpdrwJkmpMSY5xQsHTyxEUmmAVjMLwRIzPrNxgyoRBNJ
0MrWCMXyPcprgG1kNmxGFlAUus6UqmQAOkpDp3fJ/npJn4Yyb6oXCeMyHKG0
3r03QO2dqb0OAcYw2YhKuV8NlZ6f6C+61D8C7ONdenxyRyFUiEyj09WL2IvI
r9wB9Cm2mFtcx0NSineYUOfVYeiQ3ZumNOzUfl5rYN1uMPpRv7G+HVMt7rAI
bEx9WRFg8RU9nVtjhrd0t1F091ET05AVyvUNFkumKiGqZ6DBVM/W0yLwp5WS
ynA28pN2sISFT5KCxwb4NoPVkmniPCD1/gYuPvbBtPLTmmeZ/fB/gPSOSWeJ
NtS2Ql/Khu/JX7MO922iMYyP80Xq00NUB/dEgGSIEsRrAG8Bvj+rNN7m7FK4
IXVMlrMk5xc4l6gCne/mGlXWLV/shVv/NxwDvqvdUk/woNnat/lhbHClz0nt
OSsFZKcWolwC4knkK8woPHwdVQpL0bXFdiVGuGymjN6dM3EJBaee9nDQLdL7
9nCmqQEmXOGxRD0zPEDILsrtm0y0pyYUUTAssFYQpqrr84PqbqGP4NG+g0rB
tAFSHOoDnyaAjxRpN/q7unO4a+Utj/y8SG5AMYh9BdnrITtR8NbfgkLS/Gvx
Rs0sGRk0ad2U8l8e9/RLNIodyYw0JgvjHZ+5x83URGmsZFQ8tt3nXFE889NH
pg1DsmKw5Or1A4b8ULEDmzHDj0VETH17mhCUtWinzLzWXnpUPGvLmOGG+EB/
AmRLstLC3CD74woKuzJvyBvm5eyYXiwJEUZtEYHIeYaRFRvnolSZpmA6owLA
0PFJiaSv4oxhhTuvv2mm81ONweH55+QlowzpTRyYmi4aAXxGMPbXGqS4sQnJ
/c21V2Nf50f4MOFVUBrs3uFQZ2hikPYP4EEh0fTxrEaFLsGBcRODJbRuwpWV
mBfwSb9++ccyfM6TWksYakv29z3zx2joRNAQQkBUNYRuJNDz+Bcn1WaH0Ici
HUJSZYZMOIxl10Ic6eguNhD3GfzmAmZbtjPtjR5lfrmVX5XLD6u7vyO8qizW
AQQA7xuQzLg0/Kxvb9KMqwEiiZMLiqWHPvVVymmVq1Wik3oxdYxOtW2apuPV
rgYwOhHk9DmZ6YjYPAR90/AY22d7xcM3g9JnaaVEMLCivR1Dx+XC4zmzEHvr
zK8jjtA6+LI7hVG8Cy2x4CI+AgkwPYgYEGJRsnhbhIYaLcyQTbRK8LEYIf8s
Ru5nGl3a+0NNfaZ4Q1ENNXFROBQy01QFSEhj4r/3Yx55CLnyZqowtwNFwLFD
4Fow6bGOC1kT2f8qQzdtEspQYOjTKLcQ7XxfJUqMsZM5jSk/0ZihPNkimFMb
WAKnSuCimNU5XRzbD6pbv3y7SvlAOezkeW6YL9JGpjQgAsyJlJEi3meoHOZH
GNuW73gW+qSIvd03CUmU/3zqYbqxrGXBmji5Bdft/oNF5S3DdnJhuxcdLEPO
Kr3DTgSMbNEo8Dbbl2/eanha5vYpb0LY17tCF+DzZ1X622vGqVTANaOAeZ09
VqLpM5+OD+SQYfLHJTi05IBLipT4je6nLRc2OPCxPhlU4Rvn8o0Mctz8HwAa
UIhAhvVnDVuLaNkeyVQw2XWxSX3IXFfRgpO/uHmvQrFchQ2RxlRIHZs2pafb
WnPJHIv6OpW383E6XJtPccGpULqc5RNg4HzjztBDyKIOakuePxMVtveqnot8
NZgVpvh0K7foR3hNRhmPAE5e4zwfhfjpRY9+n7S3MCktiLj1UGr0bSENy6Zd
cF8oGPzEqv715tXktETVdS7erBvvBZ9f/F9Ffk2fqx6vTyqsOJOdEwDFWnDx
QxQJHOWWkcQw56qxt6rrWvYj3YHdd+BVhwRMq31fx5frZ7ZW/AgROzw4kAno
XIddQ8fYgFSZr51tVXe0z7w5ByLulqmpwkvzqPiKKf7t/SAOhsvzRuuWDjnX
f0wDpnKLLC+AN64ikFDag/R7wlLpf/zNiln6TI6Cp2wg9RXhm5128SSgbYSc
SDukkl0IYbsz9Y0Y706ddz9TarIyFiCBTV7/viNUjWzvXWFojokKBMryFyjL
b/U+vamKUx150qF4SuATDQX2jMPM3cNYNWWVuliyoes/cvtkoVQvkcm+OU51
G5j36Nn0/RBWWTQJ1JFi8JLy/A4hD4xgAYSM1Jhrz709NwErlAuaeXqsLCQV
4OaIRmZ8JILodk8sBFYib/RxKkYX+ix/OUmCchkSekspzJefTi0EkakWNLxt
e3V26xgKgY/UBuXS/YvopXQuvomUkyJRXK9FAaaa36P4/F/StV9UZwc+BYGK
ApJ8eJuHwggdXaM+6/7UbDB5IxB2g7E4vLBNfcpW2vyxQhp5nrTVa7WTCgri
S88GiO7Xr6pgxV76PGKuSFWy8FMlT8zUuz+yz/pn+qJafqkMcixTTvL66l8Q
9VhuraXOUOJkGMs2+48qh/GZzxeb9rXGd81b36e2jNVBNa/2UaqpYC7nxGlL
UPrDRtRhL4G9qGxtf1YSUM5uob5HsiWBaBm1NXCezhTSi1Wa1HyGfVkKQ8XT
J4TVWBnmx95+5dz7NoVlmpd73G0wutqRUlk73+fFkWdOeDYkJLZXG/WKfC9E
Rwr5QeVs5//MT9IAQdRUyz4+V5Nfljra8P8XXnJ4GizVUq6NvXbzQgJ89PJ3
AEmv1il+4Y+chBJRTpmlxPkt5oEZcSAP8wmXyg14/PDLjdvDH6UGO3I/X8va
J22gYGV/JTYxyBu2OZx4SbIlej+7HsAnTKQ/oKppQUf6TPYnVQvW3acO2F3d
42Y2zW+D3hPnYSc/9AXZpI6rtwfoGFfBjRaPA6DnNGPIEWeLTNBTaimrudU+
5txcBHSL+VVUXhMNgJPcgqFAGYESjTT3wtkqd8fVhD2qSfFPhpwun3Y+URY2
36VNSjxOq+/Yupk07JKN8fisbeCxgveayVRMCqJwlVigIZ/FoQa2s25M0pll
/PM98JbTCtFRBmQrWEtYshQX4g8klffxMnGV1JbGiJBh/POKBhvSIwnIES3X
fEshzHuttRaFqUwVy+n/ALuCPVYgHcKaK31AlKDzM5ZdHTm6NdI3Vaij9JXP
9hd2cazIdzY9MaZLj+MLWU5erTgRhNMQoawHfLxOohf4e7eZC/BL7ssevl9r
SYla5yfxTX/VaEfkWXon7nMS8aPnwYv4WeTUSWjtS4fbFOMIqkj7LT7RY9S/
jzpOrSeLDL+9jICTEvcZ+755WFJcPKh3uq/voshJvkNkAW01WQSQW2f9lG5e
2LXrcRf9KNGUeeicES1eqZIRCkAEklLnoBSuUkpY+9mGC2lL54P7S9v8OTmR
LboD/Ovm2jECVuGwGrwHDdnfZy7Z6ogOlPKOG2k/HCUw+zK3Br1iLL7OFg2M
CYxvN6jeY2743GlzLbw4m0FNZgwLDFbKZN1BqfI11g+PYR8Tobai/+V0jzu9
7ozu6U9vMUr4uefviMZis64wzQJqvI/4pKTyG+qvcGShTKQxNh2euQtUxNAk
fdIOFR6b8qH9myLq/06x1WFVI/uXsS87MCr2g82rBm8i08bop5tDvyfGBLWd
Uzlv1fN2TZctU+7M+QDsz6u88NM5xzJuupOohUEhL0ddo8YcrA2DLC0sMklY
h6UImKXU5oeAMNk46V+MHJFI1clO9uqp1bzOWYrADE+iOzyBIrqmy7iOPVed
CyfmA01Lk3WwrgjMCz9rYKKHHrNE+ehLeWETtSLdC4NfR3j0vuaYPQxZ8KIF
HWvZG3RUGKuASdeuBMIYMsWdEWP0HR2z062mEuUszKaEttdeU6PkZ97f2U+Q
Tey2L3ArAxwzpbL/Xnw6i21Bmq8sTvrxPu3tg2uj/nNEiLrbbTiaInVbjvA5
S9dx/17YFAwpxLAhXRnNYul101oB5e8DOXAu2oO5Xjo83DJvzOw8RqhQJGPa
LUWq/GWfN+Xh8gcX3PeghA9Wn5DVsoCYAvCO3QqY8UJA8qT3cgOfWp0SEWei
N7AjJ4JeiLVNaba19PhVuXM3/XQIToieNvZUxeeBuNQ/O1gDJoZscyOk/FF4
EIc2EgfzQcdDVARXTn4vl+u33ahvcmW6UbuO61b59X8aat0UsjccgDM9uaBi
ys7M0v8jlKM5LjRcdTk33dlE8kyq28Po1QDVMfWR80BdygWCLmFkEtGJOj5f
Kv+3AjdszMrkLsoVtcB6KMN83elXmQ02+PXS+8gYQ1fRb6ZlkYk1ubDZys+9
7MWpivunqZcRqjYX1186HrtrBrx3Xt4+J9tFyVfwerGd2xPC+LmbLA6O7AIb
Vf8VI+U1b4IOTyWrVAS906Q4teYv+XDr11YlTuJhRAIAqpZfMvfrSR4PEfYP
ne5vRBdYWpIjk7VY1ffgS4p732xvECB5TxRI21VF4+Z2aF2iBM86DPgMgU7T
ZAhAnhMHD3kYKtYwce7xZUqjwhFSVKLLS+ws8Hvy+w54GbNh2PvpKZPMyrox
sb7pyXaCYcELikkaqaLImduHRc7UOvOJbC+z5jwnsUsZoIjbQN6sPtYtVfET
OdSRpyXyXFIgVQUt61VH8xGwt4RTSxVXCR7ZTWLXKnAU3BN83XrHHfEztcVo
kf9/ZOzO1tWEc5k9umUGa/wTXjEML+Cfoc9EBbOKK05VRfC17ETfnH50hljH
RVhh585BRbBDa26vTsi0mSkiyZhWRABBknJQIPC94sgM1ZMdzRFlG6VLLATW
ag1o2ZbwX2Lo3t4ueAVYBo0yAXvmos+gliRSYicj3t8QLRPNLFm04uuydh6q
VVypr8FwZAKPeDDUDUdR7x2M3BEaApbSi92Cjy78aRYIy8XzQNgMMJcpZjFj
vLYPlefHSPnCN5li8b2K2zMTVZCTJ2ACTtKaos9HgzQXYT7ZDVUnhPqBQb1M
kRxNr1L9TFEomytHBy0aXEJ1sJH8n0XnDVeVt7lUBvkIwAmqeycD30J1BIyK
h1n0swdwrfjrUPI7OK/8G4OY1fzP+BA1JbhKW1GhE9TUmNuHfxRDtkzQtvyp
SQZAzCyW26vJwNDrDUJm7DAmx5vwYekEvwWsy2KOW53oHBXtHr8iibLjk+C0
KZwLF0X59qjLbDXa7VA7sd2OVXJ6jHbwLMSUQjtDUjHBYbHwiEQ8RqDvm7K5
riYGLUKeDaoYwMgxbd7IPkOtwwxj3erdIwfvyqg4yoQ8E9ChTJFEs7fj80Jw
tiWilcnLObGfUSR8vkmNqSoA91crPudW3WSAyTherl2vJ0gZgpVqTDA8L2gW
9TCTr98Ani8KRDxU96JdBsuYjB2tIjmjga7CFA8j+elUN6qWS7Tu+qPYuYQR
BA8V1u1dsoEiHJkwP8m7MKHVy0ozJJ3qW3CRNTHFpoP/hLORaZG3BlQtBEln
YzoEAzJZAy3setFd7lEIbJrotd9qzXTCuS0svh0qhVcBLkab1XqO3M6xSEfm
TOOVqrjrQ1eQ8hXzSd+cslIAnUsV4qEcUtwfmmXu2rDZvtutcCfHp3qaoLRa
M713GScz4I0AzcCjGjmugGU6sVvtDk9IWqNzSmfz8t87S94GlP5inHY1vrUk
ODQUNgHVxzohCwCxvYZaRjjm5PnoybHXgWNx4JnySvlZHi/CVOlSAEgGntU9
a91OEd9frjSbMoe6fvgXz8LMkyVkbURfSYmh+NaZohMDgaRjd1QPAM40bf1h
xQ7Vw7oXbFDxLuyBnrnVyk6mR6fSs075hS6TebqhH5birF/693N1rbcMUfhY
uAfflBdw6/oN0868Olb/JW9GkdtsWvRc/av0wn8Hh556uN7JQmyG0f36vY3T
jxEJ2OB/ZCq8NY4/KotuKM1ixeqqC58AiWxrULmTzHJ8H/CPqxWV2lUXu7j1
c2wb0gr/NEzNFDeRiZkZp53tl6U3vItM6wITSORH2Rly6w3e3xq2voTCuvMQ
8gOD4RWy12Ccib74Glon9iNSd2Tz5RhHLb4YtVnmEznbtZ7sgV3jP9LuZT/O
tMhfNRXndJQIl6RdulKn54RHDAbjnZ2qaPNet9QvHBKk5SDjP8WySxRNrDP7
ZZAg+dtyRU80kOffakNRudAxjsYwnuX6sadWQeDwYBcq13Ksv9fVDibHNBJG
Ii33vuDIoIJ8gLvbe+h8rb+oRIYb/HUpx4SKqbz9GeoBeKyd1ijECx0riDPL
Iw4a1pQseeH1vYdXwuHYId3LLNW61utBI6tvEheyvePq8s2Z/WLGZvEJTWH5
u907dsp3mwB+lgHq7B8OCtMIvcwo/TwzYhAPH3NIr0WkfjBdDMikFRNEA0Gc
8Ic+iGUEGQVwoqBOtpqMsrTEOBCO8Dxz2wat4LLyo+IBjt30+FAt+Ttr0Tpz
YtI74ntR6u7reOOlLo+T1BgS+v/Q4bb+szc6at7YuYCH2AbztjVEOYhaqSg4
DvHSjh5ixY1ToG8/EtPjxQVSI+SziFuQxHYWsfn/8xtDa9amcMNgQmmxL8fz
J4uBz9YT2+IDPX7cCTPEYISTwnhoqO96KPQ/t3RPIef2tsTT0od1/gbYOFco
zftahciSHeIDacHdRaHLdF1+GM8OiqyNdDOZxQwLCwqJZ4CfwsuiNGjW8n/c
obU02ffw2CezvgOI/C087C9JvxM6QskO+lPnikB+1nihKbGcGvSwzOKA5ntP
IDfzwnOQeIOg1UuBLipFzd1+cY1SM/JrvX4ZOfwJxkp13dcJ5pOpaiBLOU9W
g3ToI/KirpQ/5NTsLQZndmENveqGw9vvAgW6kqI8vuD8cfGlsiL3zuU5cFMY
P7xwZWXx1isapByukfnf9ZI9OuHQeJGui2FYrBEgGxkemqMEuI9uhI3iZH2A
cOoKJhFjRtDnbhYGwEGkTcunzOIi/shs94rimldlLAG+emZaYzqOcxYMR8jm
i796rEDpIHTdlIUw/K29jrdW8nj7o8Vu21uO1MzhbKHRkguvAw4kd3Dfnmy2
PFQNoDZY823obWD0u6kNgCcUqxxRtyHqtTA3HtY3NpMqLkmS/h3BtblgCCZk
vJzzAHUZaWpvfPk2UNXnUk4Lin6OBds9918p0WMurlPB6mJN3KNp/JalihLb
1PaxPtFg39Oe0knYzzqFc5KiZ7Jic4Try1ig5ZhUB4Wuook6E/9wc/WaJPk2
EgBJ42QHCCGyjEA5LeVy5IFTAcWdk2Lk/E4KdiCs8J5uKQafI5eSiRPHv/BD
qganOHQrNwaw+DY8x9JnZmubolXuL9N0JZW91UPdcYg5nU/PO/IIv0tSsGBm
Lwsw498DbPFlqtNElu3rxI7bmbSuyXAX1SBpiaRXarcgrnfbmYpgSt8FkH7u
GylWItojK87WLv0Tl91qsJXBrvbSJyVNkSTDN257VMXyUg/3XfJ0stlSmwH7
ePQSqcnaJenlqtE50yztBzygOUgEc7YwURP+38/XnTDLthAKc9skjVW0o2fW
KIr3fRfREKEPkTdX/0k5kpyz10qI0HyXK8qAnwtRtWqGVb+bVmcqR3NpSdl4
G+fX+Avn52lhuJD25hfE2Du4jQd58NfOJyU14TZKfjHiX0EFGK1gVsqxdmDp
Wry3yjDgQqkyw+JFHLa2a15xEUz8OEsB5FqXY11LnEoqimL1ebzxqtk4Yo23
9s0UZX3ZYw67/jPyRqlD/PqBCsFTTI/xKpidGtVmmIBagbD4N1vSqXcrmlMk
09CBwPI4bqfVVDOTMnBdcSsCW72pbX26vrxHEwnjZ4hCKwdbjF6LWQUH0W1o
/M6OMHmIlWwcYFF5M3fU6uYdqyiMzUabASq49X56f7UCAq0FrJKal8i8AI1t
xZf99/3jsKEqFKfjEp+WuzIdCUbsJzEKdXJIvqBX/XLL0hRt8vZ+3BxPOWE/
OEhKXRg2VI9pvK4WRHcJKFg+zayPYpCySgrg6i3th4oMgQts9QlcO9sV5/1K
peLirQKOkgy9sSnQKNUcGsMibmYe6UrEfqGk/RTF2fDGrcWO7pyvqtElISOT
v1exTwgQ+myRbWsNpJ0iIv8IHty6s2rO+7OhZS2ktFzfSrJjdUBwzEH+FbOT
c55WZyB+fmvXvHo7BYWyI5o2zjPQ4aXH64WXcKsXUaqXh+zeMdhf5U1DvWKR
8n/DHWCl5vxvjtnwLucP2mnDC12DOT+p5bl0Obj4yD6Vmt6T1IthNEsJ/ued
wl691NuW+mhghYMpSJuFfxC14YK7IWaL7U0oaqRuGPb1GJmNjSj+w3WXXN/Y
4wP8nl2hyNR99GQxBc5TN2ptRpP1Hev3VwXZCUD3eskTX6oyxQ4dWetKVM+o
doWXqW94PLcX7au8QPr89J1dWiy4Dc7lQVi7TNiezElH+oRyd5/lYmtcKqYf
EAFKZTv99b3vLh37RZ8sOX3GH8eUwhB0H2E5pur/MmLebKyW2B4dj/cDj2Lm
N0r3HlVNsWpXdUXYtGsQbqV8/BctedFsz+Q8SutCPSFq5vJcw2AAtlF1Sf/6
3s+0hBWZfe6e/jDECF5Nzv9tRUh2GYD7mB9FpA/TNYvOiIKQH/JOF4XttaAj
CppbWvw+gvoCd10fOo6uj3pSqyY0Q4XDBkGdQ3dBpZwsAbDsK1DYsACS60vV
vx/XJOkWWO2jONw7jC7YabUEamqzezVnVmfnPvAhk+gAovPNpAkx29vwgE6h
r+luhKecq8xY2J+8QC7V1egdEFi5q8znJ80+q5umbHZIE06UwHWqy2LrQVqt
AdKTTtDvfI8Xd49ezsRWyM8/q0yjOJ4GjwQzg0MlqhYnYQpIK9B9muA7dTH+
ZeyD7TeCwdYrkDPOtgmTCk24ML6dFKqGH+8K+8AT8f3g6yaG/P1qpx9GoKO/
gjSXB/n6tNEFxou2hvISYcCJL7JS949oFBcV6oqwVwR9AX8PClqdX2yg3ZCm
nVdxfdSfcofubHWT6RLhIdVFyOT/ZxsGDHjGr3xlarIejDBmpqhyT9Cc5LUn
GBSuuGEKOmUf3LNNnHXtPKGASZya/yCL35n76TyynTzQRaUkSWldXBoBjpou
v9SxvCWXATVdsPqYD8g/6zULCOkUAW2LAMR2gUYMUnImoCGQKCLSQGWq20OO
IkYZYBwX984X4myaiT0XEb1fLnnwi7k4wFBdVLvb+V/0/yS/1wxW7X4TJHF6
TMtB5NfdjpDwmpMKIzrk27/gw5nHTR/7vmvM9yyeaCKIAz1UlWyUCLyDzdvT
eVxFz11AXAnu22GHBMvZn8XqoXmc73m26qQnOTWa7bRzLkAq0lei0Y8TqB65
qBQWtN7htqLfgwjK+W4x+ZzlFT94m9Y0RHl3tugGi+c/Cd8YzdlTe1UWtlir
IjTJVZaCU60mshwjHn2eYEjdbdENPnyXhTZo3IZ3hO/QJItpS0wHCoxrcK/e
13U1QEu4yA8djvwpksMIhYu0s6PwfjukSoOnFlb0xwhPoS/ojYQtcEqRcL+q
HStfcHNRJNOHPsxJHibL8yxUlMZsLW4r1YxVRttqfSBsb/6FGN+nmykx+RW8
IDgLk6F7AinSX0Gt7yowLKJC0v35/pLZqCsAHZArC4s/Pa37ol293aoEJG+q
D2XxeqrH90vHE6S9Xz+6NOAddY2kd9Ebihk/brz0PgpF8441Y3P7I6XLwM67
5gIQ8DOLbi/YaCGpea7uLDlpVfe13X+7e7RzULplSnR7qsTaEEEhEE28lDMS
N2JnQj90DP+DDDMwAQMrwMegRK+tiRVJg9Kx/qJrbKCz5E7zoJrB4QcZKlpC
wSkj8R762zipBgpuqLsrvE1K5t0SrVupkIj3w/1Eaom9z2xYycx/wlJW89Ko
raU5xB/rJ1dz4f42yzOVLwjG/2lZFP6Ddu1HBOdoxtTqWvOfQDiLnvqTTs60
lbrIYEPx2rbk8ilcp/Ulh9VlpKxZRbsuMLCh5Q5gJ1BpdI7TrmGyuoK264YQ
X/4ElasjVW+BS61gigRe+IuQ8WMv8ZqrJKbQlvfQlcjakW3JOzFKb47MoCIV
zJUJJUJurQegcCDCOe87/jnnZ1JAQ2hrBxPU8OVNO/vKh2WvJ5mTRZ3bzzVM
jXxYeWg+2+4DZ5HVAVbe2jdzRhJLdZmUHhXIMLsojxdcWWNjLIvbmeDlq7aY
q+pOsnAsDJYH+pFTNx/xLi4PX5Ku+2yLgXd/2btgfETPvtoog47AdNQpwvp3
UetUhok/0y5u6BozSn/ltAx/cJQL4sSAMGlT0DCl76s6UJfvZeqezbNe6uyG
3H5LvIU9+1Xj1oW5rVw6gmdBrj2BE3xb/X2rj5PIQvTUK27hosZYowLBbqFD
OfAWIVqZ6+W3ToT9JYO7vjGf4CD5snrsRk0fKEVNUYERs3VgEj7ewJ7UZO8k
kZtVmOzilX0Fyvvsw9Pf7wdaT4zi8/996pfJmR+USXMcw/pmEphqwUq4SyBn
/FhWbRwB4FOqgrKeBgnSzuKQf7WhZWAJW8kPA4u3CI7X+X5jScv5uLAsq8eq
NTgImELAej1+VVtmQu/aH4JHg/RH40rY7MvOaVAQz5nZ5iFAoNtdhj8S099Q
F21c3imasCEBXJpji6J1mwZbT6gnM/x9Sp/ur9wxWwaxFXGdn604H8dJEX1l
cu6h10LtSS0atrxI4RUIblZtrGGTqQU4sra6/STLUUokMCT3ui0bKo8Z4dwV
6cgLNlDyix9ACA73x9aGbLsgpS8aCkhIL31mHETEg4YdMkjBf0SMWVYrbtgw
efberAaYt8uLaIRZ3wM8dvLnOIHpvQWQjYaZIUWJDVZlvddRXFu62Paf0kri
hW+UFrr9qlsLNIW7xcXF/YkGnc0CCtXATSMVDQdsy8mWmrM9gj1DrbnVHd78
y44MrCrn7q6VnHrdoAjXUiDqexotCkyvU/1fOT5ifW6yrivVbxB5sdpgA/yl
/Qthl+ZzlBd62CVpTxFbkBtLGkws4MwUGyVNLm9HjOLn1Z0WV7kbhUP1Nh6D
Pc7Y6Erec5iRW93CmXI6myJsHktv9hLfKyG3CDflrZHx64OGpi6mVAbTjkNn
qFWQq87Mrv2xLEMSoCjDBk69SlKzkRkX6Gq8z3giCzAro3d9V5yYprI22FjA
jwpDs6yN4OIGkUPY3eoXpfecTmjDVsm8zTcqq4pydJKFT/XVe3OgTjPeYFgc
1cCYW5JcqQB66X5weaFYr/xTAWcm/Kb5DyjRze/Yrdd7nO4pV2iH38eRPt/W
Yj5/1JYbBROOYZuX+wTasteaSzlPgbDHuhhrBWKKiLbDQLUzKrsdsq//CjRM
1riIlP/OaIfmxry8b01m/ywdm5NsYfyHifbMk0iHF9Fwn31Qgs28M2WzNQNs
EY0Vpcj1cll+hAHEu6OKczDv7SKvrIXfgXhbu0k0w5x6+os2ts8lw8rhpYQX
yV4//W4knEOpZUMOSqdJUiYb7Ku0lk1rRt3BY9POcZyHuQzu0qbXyFTFTJH3
U3nhiUThPIYCPdGb/z2X0UPNe8RG8MHrMl/DjEfJKgeuaXD7KPkHqVeDIz+E
mTp+Vb09RKN8nH+aQMti1fkra7QvthvkEgyQRcqi5K4OjazyoLRvWdhSO0IF
40F+oBOiU/rnhd13TC9tetxirB+Kle0E2gGSI7IW+DBJeGTtYmFvtEwo6ucA
ucHxGap5OHYBnt/aHhv70uWR81ZHGwKMUXHaGmDLFxYqX8DoGqQHWBjr2L3h
rtChrSYIXQXGLIQKxphxIj/cos/pOF/EgEVBJBvMXKCF+JA3NXDfJoMA0eIH
7Cp0x6QxF7fyp5ItIJX6oVkm8tsr/YJM/tZ9YhF6VkrZEYmqeDu2H5QW23Kv
zLVi+lWdFvOZoAKXXxXLUTZfOeCYF2rxTdhvTPD6M0PqNsRCVaRNyIpRiXHb
drt7UZcLCxSAJcq4xhgVn4cTnfMbxKUHevI7sFC9g6N2x5aguCLs/ID840sY
z7MsWz7m/LP2eiL4bxglHoHQJF3SKGp8h0sJQhpwZYt4x24Dxlz1k95MM4A/
0YTJqI79sb0zHPPgpkYQ3Vi5MxcFVdKknCQz6H1oyGkRbxU3ooyHb+i1J5nh
bqGb/ZmI3241o8YE7CsGX9iT1zamVpDZoCy/PPAslB88QDyNam1entDb5dgz
/cKN2d9b87pnRFUd2RPE9YkS4MB+KjH9yoApdeCV5RhNg10eErS5+BC1gloT
SQniOkKMZo1PjWi8eN9VZPhmuJOMnPfhadW/h7Ld7RG5s6EjOkySx94I2lWy
YD8rz+JuDKsVLZIG8y7KdqgVu/ChBRKAru4mtRQmyUjTTs5dBKx5TLNGKyXp
FY7eSZBlkeUfdoVQpxgW8EKJFtiN/2Fm35AV/smh4/TQrB/ybf5edFlC3pzo
+Vk8YXStonFYRUfaKoAR+P45jAzbuJIdoNZ0DXQC0XNHw6/7xoSztTazYZJY
iqzkzznyymVKVQq0bohEy9yCtZo6bzW33WRR4smy9gry5VBmzUgO4g+3zVPX
O60acpAOsNeaPc2pXcJHLP8GEB3A1BmNHbjEwWgkcDoF5LODN7e82csmvTIC
GhFiYCDbj1M/w/fNAs7d7BPhQXMwdBYmRRPsoDwWqcMBwE3MapXwY4HNU8vx
jQAqTdP4xOnXO0Akb7x8QAPHPu1gKMWIwfp1KOhUIx1MhCHFvNwlJq/YUQw8
8oG0xHOeQVZ5jZ5sPrF7dVQEmQFVyQSScX2ZD21XN41PqMo3/N8CNgpvMd+/
hhf93rqy9LZRPRMR5ZxcaCJxej8zIRm4ZEO+ucgeSWx5aYDq1KmN8gSxMrNX
xkxezZQFtsA4Fau5yKiqLMF9Fg2JS2lfMdjmnF2YzmVeIgd0xi5C0DwLJ4bI
Mxlvzfyk5FNKPWv9J9mfg+sR60AAlh3YfJ0+BQ/YCY/0UAjjIVYd26CyWHRp
9KSI6hAAeTBhhdZ2RzCvB3GU9TH6tefK4MtPLq98pUkmgr9uDVkmj75NrKwl
lyrXLZZVP33bcy+S7xbYpQGkrfxKFP0ZN7ajKUDYEOn8uoUM56peAa/G1fIU
pDDt3WLK6K1mSayspm1uuAfa7VrHKQEbBmNZjNtkMrZyE8oiqh8DI0HrxXhs
xHIB5769sqejQAjjfGxT73GKs6d/d8IZAbfQKvRoRmVo7rmPs4xjoKDLB2/e
mLLNCp9pilmQMav4wZo2EmudT41YHRZqs0s7pe9HVNydVnVfT9jQXQyMhjqP
mvUrQXj6EfKPK8MQBhHu+Nwnc7bnux5oeTzWhQUHIcoWSEFfiBzt6G42PTcy
KTxriBik3Ll7an5HyCd29eV+bZqGBTWrFLxMvkRCyaxBnkjambt9llLu76yr
tjs+A6SC5rO1NTndHA1N02K5WWD86q+jYQCwGwJruv9HSSAmS3XPkX+SJMlH
LWPD8YH6nTvqNea7o9trr2kHSOkNzkfmt0hnXvXkdBCCmstF6BSbSSjejf8f
vKIQHzfh3n5gWgKrPDpySY18jZeZRk1FkBgPymYkMfVcw09eSpYhx+sat17I
exyDdIw9ugXpXqegVGEDSUUH/8BpcaOKaORzZftrbpH4sLUWWLniKqakPwhR
4LUfmg31onbBw3d79/GyPfRpJc9yj0vacjMtZlGqGEGKy+ozxsdfRldo5mVY
YhvU+ftnN1ZYP9ZxbmKP/enmn2U0svg+pEp3VGT6nk+t/H44ePDlEdqPrTH/
4ovKbU3d6R24fbaxs0zs00ik6oToS8ewdnwmnZ8Y/xDZBgvaGwomR7RGVOcS
Bi0pesP4iefSRmi/9hBlxSFKsS5m3t6q2MbzoPBKnLroLFCtgxyP6gwwrcCg
4FfDamC1WHBkq+AtjReArDBGx1ye1KXYQWMyoobb1q37qmGCY8F2xHAfPlS2
2ORBkHycDeVI13xlSMLuc+q78xhoxOhzCiVwEJb95EOZmYP52v/IyyZ5IJOC
Wt2vPCsejAF+OetF8gy57y5MTZCFYD431IsO2fsctBMJh/OPtmCqoXUNyXqf
deej86tUzpIm2cR/2SNnCQkSgC0dpQNwFNTu47GSINlSJhydJU6tuYpVTHtW
DeELBaLR3rqAamWITtns++1ycq6PAlMRkHKjDqO05k7IJaKS9oGVpcYMvn9P
xdEQ8STaCY253R+rmzEzUT3ZySonytU+QR446Pz0vOr1DEYtdtBJuyMMdLyl
9dU+z6L8/8EPI511dTpJxfsleDS7b1qkGTqPz+K7HAc3QRHtcjnuK3izIkcw
X1p8KK8cr4Zz68Oo20pAGMic45afZJzszm/O+LH/wtt8bxXsMfOi1NRF80Cc
/Rf6NVIlDqwWEia97Xn6IiN8f554RuDfVAVj5gQabHQbFLVwaE+vhTvjLGKJ
42t1wB119YKU6P071Wdc8WkJ05gvlzkzEGt0MWPHuv+VLCeanh+Dps7x+pEB
SOZh3EttU1dmaAZ7P7pizKdw6GqAhdmQwoQEGNO84vK3/2u0qkgiWtR/HAUF
0V/aNq72M/oijvbUCrabRUS3+mCb/NgxoSGFvmSgr5o1AB/EbO1Rjh8UeUcF
QC19bRMZhLSvETBCT3sKCixXUNSw05Mr/FBxt/ZRIUiUQRRIaVkG81o9T1p1
uvTO+donQfDdi9V9oaodcK9tzwSA8T+ieT1QSa++NUQd4Jso5X72I/C3JrwM
bQYx5FLkAPWtrMP84YY+s4UEsC/WARtQnhz4c0ujzO830Mc19SWZt4Byl2+j
iLc/3EvYzafpmyyKPUwdNlNlwhNaVvPklBYM3TXr9t+A5Fb9sAfvcSaPRpPO
6ttGiCQc0mFn909N2QIWBGnRXcBRzn4Yj3kFGggSNpJ5BevEgUecG4cvTk9P
FAxvDpGY+JqEam40vZBnQZCvDCuOahMyoHWiZ4GNrdotRNV9YmcL9Tq/VNRA
8H3zfXmcXbT1iy++UER4lw4ID2PJKvelwryF5DcLc/jId2LfX/4Ff8m4ec0a
vsBvwBkOINiPTyqM8BmFevtADbmDE86+38mkL5vYbxNGobX5FTJaiGai2hvk
2QIYvTNx547wRkVuluZt6junlIU8tVQMtNqJBYdzo2ifAvUEwHabRyyf/YOb
4BDymAh35v2jD0XRkhrWupuVTCjV/7/5E6X7rYW9qnvf6aByQW/Fs7s86kEk
hKn+j7u9VelkTOhEAlBnCbuP4G+Eh38cr6QwQypyXLIpbM3qniB2+D8W+8HB
OJv9I8yrXMTAKV40+zXWMBbaNT7yPw9BNL9fPIuIGUi8rDOYnoAY/yVOa9yU
sqbYrqi9o+XlWwIz0hMfYD4vgImP6jBEXufjJSafqC2JAUVNqLLCl7ltR1qf
Kh1GOsCUDhuiKs8nEswdBxDzJVRIQkNqIdmeWSXP1QKhLPz0hjunFgQ2I4v9
e5+Aj1hiFip+nR2mKV2/duBAsR04H2+Djoh5RdKms67AP//tmRDvgT7OWjJe
Invyg8PN1H2SmNJEGiyMufSX2rn7NTbjhX2zwQGhQC2orp6+HGQ1VAWJPT7B
yUASoUjiHQ+2KODOJKofqi3/rj8Ay7zP49dmi/a9yyXlIlfpUiNzNnsdSBrr
RpPUH50599azZa9ZPCDrVjq+PH1zA3woXmipiTSF+vF5ic1R7AzhK+u3KnnA
3eQpjwamzLYGYB7B7+IUyIS8rzVNqNzOSwHJG1SNyeuU5RhoPKkgsK2oQeX2
IJDEaHQ2afuiPq4AA5oNK0ltC1eS85znTSr69tuUGFZoLUFSX6odEfCwxw+l
sYjr4PnkkrEJ3n2krzbhRK7p6brEfK6IQkIhoKzbCkSeNa/RPuyk8RRVIa7h
YwKiBC6CphMEpOVPc5kGMnx2FXLE1WuE5AGY6HfWnks0zPcycdvj52QHNV1v
fwzlIkxeHRKSKIA2axy+Xon/LkYkep5A5VrqR+Yp2rd7RR5n9OILUZaeczBK
MGjuYZrPsZZ09POCeVohZosbP6aNgjox8ttprTYJWjOoP+7R3icTK176Oo+h
HvWO6lYjUsLrCW+SPd8P3F6ZL/XTG1hMulFvnE3peSJorAJexBb6Bz3XJvrR
AtjRY/ArmC4KbPSb/RL4PhYsEhDtyy4hH/8kSzO0OsRJ509EXZK++iU5Qvc0
KWVxjTNiIa2V7qIulbTa+QFkbMs+dzjk2gSZEeQXjJAA2+7aG8xHc5kaYXCx
m40SGWZ0Hmz1jfF/fN3gZAlRPPwAVYDE9Ts9KDZ64Pnthh3/3FbDR3Q13utE
sf2hTwmP8K3oO8O7W0yCRCKK0/GDa7dbx3iLurs2Wce0F8Y5jb3t8l4KcRmj
lUhhUr3PK24+CqthV5ZxWoDunKNP1HLLmBP50iL3CJlSPM/KDWpy/C++/tK7
xnyiTcKnqWUtxL93iDZ6pf/f6OX707t8P9z7wSiGoao4+xN8iJPBKAZaql92
FUgNpB9cW1yxyrw1LSE5JYlK1luRs+4ASK10GU9eMOblmMxKkG5sGiw92JNZ
cFcsI3W3UPDc58cKP631rRLmqEZv+JUIxBNiVXQ7Mc0RqiGJzJm1rGn2fUOx
XzSH1OT9CXSJW5db9ccCC38jYh5Y3avO1q+loHhQHeAm+Vlas1E0Bf8HR87K
lKwzNIhcTIzDjqob9OVmJrscp39YzcAv2Oir4B+3Z2AQDOIoLlM9zMA/xekx
k1RzjEyZ6OJZDiK0nWGQX10nPcdV8z3ac3XQJqWvhyGchZ/PTb6TrgbqcKwt
KHmxzXGMNOe+FM6zKJLqgsVe2P/SFw8cXKk1AsMWaNjOiucdO26bJq6909Mb
D8YDQpyiCzvDamZqb0NKszJ+5r/PCONrdzyu98W0f1+0kXgokBDB1f7teG5w
FPoo+DPPo5r5zdPzTpQ/hc/KoiydxIvc24P0fpImiE3tyltyh5V91H1yPf/b
m6BvQKGqv56FjMJUCIRTKRyqjNKjK786iwSWcwpzeDvkzRtwAFEyweMj1sxN
dAllm2KvZzvjF8I1bD1Q5nTvTxhNhNuVbcP0H6/V6FVJ3DjfkgOmyqN5M5ZP
+MmVRKmVUZzGnlxU1piuCfbT5TNfWL6HyYFW6vDGe5m67h7kuxqfwIeapGZj
uB9p2KTjajslStQRQnnqnufwIA8YOUzKdaq1UAHIqSF5KimYXfQ08/KH+Rsx
laVA5AF0Ma6FuF5YqV27FUgSJA/3WkyhlOaXBx4YabErrx21+Idvq3sorhyh
ijLg9bakUXwJ8M+y/Dd2x65wB8uvsWP9pKFLpE1BfbdNk0+gRO0vlJkL1sJf
sU3MalXuv0M7jA28XJfwmq4SpsEHdPmq0fW0IdOAvJZwJ8W3fgON9MGFSHxQ
AmRL/NRe+OmZ/0P73H0O5u5ReWIUIJGCLufrX2vGm2QopNhq+0BIxlJIvgZy
AOF8sLMBtkohIL7jG8+6gn/xD6/Ig3Tvjhy+EGYVwnGgX6mVPcTZuWju36Y5
TCkfzXycJCK79xvnhd8uc0c3lq2soiGFEALx8VCbZI1OXn0EuYqzhjeLP+j3
CExny9LJM3T8skuzJWVJOXk2lp0apJR+Ye8Rh6PizdDXL9MRs6m5vmAHLucG
5MwimXQj5CrqQd4v48f0069u9b1g/aTMJNxhqe8aUHLtCiy5UrETUoi4RaOW
vQ1bSWhkabZp1aDhGXGEUBwt+lqSDhEhOy/xd8T3TOihuiZ+jb4A5hGJXY12
OgzU8Q+5Etwf2183xvziJS1G7U8A+j1bNALU40Y8/5w/6VK69XYZ8zIjcoUa
ygvMgLEsYPmuQMT+dN6sM/x21G5O7C1WzNo6OI5mPpWdCNzgJbEa4NXiKI1B
cUPv5hC7Qt1BmC/zhgA8jFlmH82EgOvFDwC1RRTmfLHxDZYz366Vsr6E8Mmx
s3vGqU8xgG+CgloE0G/hK+tRsokQBl5rMA5Rjbg41Nc96FTOwmbojQIdy+iA
hw9JnmAFKbZiQZqvA5n2/j6HnWa1FibFg+6T+GOojkb95Q5VlbwOs5/LHOqB
60HDmBA0yDjef7j5EQ8AhsZhi7IG/rEhP7q9AyqrMGRbbw9tzhioBHAORrU8
YBgg4WKuHvwiNkaBH0Cy1JNYXIshiPtkDj5TUEfXs2FLG2i7w/P6TqmggzOY
fng1cqDDPqTDrJlvjL1htrS42aJTUonJy0wO42gPh2d2/a9kFm5v5FdU9+PU
frFM7vgb7B5dtzL1hbzF9fhCLWG6k0+v1zup+da7I5hUssPSPkBAtG4HAB/5
P8To18ZGIx6CUST73sJ7HmIvAZ/ez7yt5CJyO7emKoo49llKi21kgMHymF9g
Opm10S+Oh2Vegq8/JSlgJ+8rnvJ7DQXCkFqQr7olf2elYOFcs6LgX6xikU2Z
SqNwexw4usfouYIQ5w2G/MukZGYhVqTtltPvnW6dogtFLa5BpMqdkMVzhvXS
XwWS/kghfVv2v59xqTo3FLtAlcAhkVAkRAwR/H4a5ertWoG9ulBh2ne59UBE
IP7+hW6H38K2+UQFBm72bkaGE9vxV6m6RR6TIQra348+OxKJ/QB4V1pWny9X
fL7a2dVGIbCm2/MbUCBOD0/gmXKrDiH/ripUfxEYRQ2eGXbQbkzPRRSctQ8U
1RT250wjJTKLc3m6zSFKFAkmQxTwezDu+nmX4YBV/mqXkJZRl9hPsZeoZ5Z1
Sa6diSXfE+Sc+Onn+WXeLLdWhc01cKmpRbcGUEfRB4erE0fWNYnX0kNga8zL
pWCTsgO7uaNZJ40ti7/VfkT3RmVw20/l3Ap5uM2DACpWIR4TNiyvoxAJDdx1
GMV4ABRjD9F4EFs8ZzkrTFX0/WraYwXv12WtXYNTqPJBrZ7iBuuMxN0rCCKI
udpI6SjoEC7DAMD5PP0kpDhhQjlw92XxpJs7wTtZXZ5Pk4UnYvynR2+o08DX
YzoosajAPLbUrQtvdKzSmmdH+VskdCJC4Zdyc0uaN1gHtqdgHDGOibFG52l7
SPxqVusFYY388T0T+2rz2Qydy8WCsQgRJQyPUWfzWx1L/gu2jeeXc8g7Dq2q
6pRnFe0ylpIIdAZ4fjKLePz+eMPRRHNZ+OFu56wf+FMdqre6PJJTD2ThSXLF
ViohufiAI/rONRYLfJr6Cn806OTBrdKp+dkEERYg/uDZ8o/AaP+KlJIpRb2V
KjliWJkfLV35Wgq7hr3sgfSUoCijOhrv7FizHvHQwm7PD20lyEaVuog10BYD
yGTbSeOakVXfJnw/vpkWxmMKGrjN8EXC3bTk0PYURvLWXqRjbKTREsfzgFNd
Gw0tntL94SakVHNn2RMyvQNfHQITW9IsXIjHZre6dpzV5CqCneKFNYwzh3xe
AJ0uNrKmaEhqoViolfwDDOYrNuyjkA5e52vBwIUTZAm4ynL+IHuBfeJz3Bju
NJnN0A4mzlomxr3324mNg1p8h7Mz3VQDvwn2xUe+FQsaQG/m6742683pYh5G
dLRmo7gDR+CvYwjKSVtaINkP0Z12WfFeLVL+h49Rm4mVxsBV1KNOBBmuF0VH
gACO0ECjWjeBDnkoyeCyExP8u+71UGr2JelEP40hWT/FgUzGm4ZcjwoCEvLX
6BMHqhRhlCoEicvVkmn1Nontfd89IItEkTOV9DZXbH991OKFRzaUI1u3p09y
bJ2RGRVAtKiiV3obv0dUgnvfW+N4RXMHo3siXcKmfEZRbiOQCzUZhxseZrgI
G6zuGmw9c0pRLQ3+IlB3cdMdZ9nKh6l12MojaBk/bY5DS9Mey6O1dGcQergR
Z/Z0WIR6oI0P8bpuLqQzlyF7P/5F0d9hifxzIXh6jTKq6mCRUwrjwuSiA/NZ
9fDiW/jcDBjJ6fcREeoPyWawtYv+nB19smv8Atdm1BLI8KErP0gkexN8Ooqp
RkZSEMoqLpohCwzjzzIknN7kCHXvaZtpJ8BeHTsNg1ta7MkSohGHdM80kmaF
tUpQsG9GK/I6a6iU1Z9Ij7TRTO9kyV4CzCFXT64ies2yV0v0adeNrLGXDHp7
QyzMjU2IibgkhrkVhqjv2qtPc/Rn5SUVSQZdN1dZ2Rrpyq6VtiGOwhPm0Jc4
rmOH1/9GKdkl/ujXKK/bWAoyvl1NB72fSNQ69sK40cfQU3sa+c2nD0npvVtI
G9Vo+yICZp+WeF0IbVBgk5u9eJbcREdV2TTTsbiMjngneZWlJ9dZunvIEhYo
iGM4Wls1Dsxi/Mm7r+J4vSDodAiIvk6Hngn9baDxXY4UrgudkrOA+PfbTCfT
ojUzDlSaGIRO4tx2POQJ+0qgLjUWw6RB9Hk2ub43oZ2/gHe7Mpl9iE4+5UDr
AlRGKWxh72fbbVwECqACdMCqlsbMeZovrLusR3t8lNMpEVBJ5h/psNVJvb/l
hjb0ARkrKBhaRiDkAmT5Syubna4ZJA1mdQucdrdjZ02ZkedYjJHbiEtcyJGH
/23GR/XuE3MczKQxOSwjxhWSTrusWM/BwNl90WxIxSDGGH8cj88wWIz8SIPv
V+XbuGSwlAD+2fd++iOkTC0oGcGhtPMxR+b1UM49qTksNrpuh09xjXxaPplZ
8Cu7ldYoYdT9JTlfrU8gAIIvULYul/d9jRq3pt+GJhBN/gFtNA7eEkv+ulwU
NW5ejl0GPfg5zazVo83GNtFWFsNUrB2k0NjxjZjl7hD22jzeGOLIT1IK+0dx
MsLt/Q1kOF+DImzvpQRjzbt2NHwMMgD9GU6gT1y0D1WLJuseQC6wqThxX0/M
b9Q9YZk9pJwJ6QCDMPN5Hy2/PVgJAqIC+Nnza4szUmlsAoFRByro99WTXyrR
ou8ecNyrcSXA46q7gDBboVm1nNl9WmDvY2AHGzMJfaitGoF10Pd4B+ZfTKHq
s9SWiusFpxD+WOXFJJR8COjhIEptRtwv+J2Uehg1vANWwylfN9RyWvTnMjZ9
DELJddEIWI3kIQivL3EdbB+gWJjvI9tgqYL8vsNmxmM4VEEbDMpWciMPZQdD
IGv//3rQ/t5uGY+nVkBOjxX2Mu37dxwLHLqVgLv6T0deFTfFFhdEiDORAMDg
rLu/Q/dJh3x/be4KiVtj5StsZ5JPx8m9WvmAche3XhKOReIE/RLOP+kkfXXz
9IrRV14m/zjb7CmUpPI3pwQ0UaTQ3d2Ga8khaZ7fWRKORDWv+4D3z6V7Jl11
ZLv2s5S9JsxIdVxtrCE6V9ijjJbIQjnWKcTHAq8fcC+OeaxYdtCxhVhqf171
I9HFHaWdxAn3Qm9KDQzl04k/dPkQjzmfLMEkrZHmf4wbgPDgPQUcVFCwxzEn
dyO7eiX96khVuTdm706UVkWATi6gcjdxzBlmkmglMqwtDXaOgrL0/b4KUYDn
zMVS1/hcmf14Rqu+JzehAPzzauopV5uNBoZk3p5kEhvlqTzqun3yDA4feI8k
7mh5hdeCcc/P1k/6QMDMQHqhi50ZJ5xxQERR8tEk6IgJnb1h6N1LaF4PkbUt
WR/Lc1HngEbAJsP/sDySGpZ0x9BMWJ2lQA47rIv87QUWgiQLsYezGyla+cLO
z5Unv+NTNzZCjzdhyAlhB1gNyhQfM8/EboIga5NN04u7fi1HPbQvYsSlvyq4
X/yQ/9MnWBXIvQxnyD5ay5yKeLzNsPPrFXTk5VhxU9bXPR/w7vehs1cJixd0
xHXnTYhNWLzKKBjcVlGXPb3VI44jgqIzqiCUNie7L43G87cw8Z1CCljq3uqQ
9Dp0vzKGjSKuIRJhJOsWdXmJABtfOXJuR99fKUBDFOCS6XTFyCySPMZTXFaK
Rfp3OhuvA09zSFVVeRRtYcKTDMhOX6v4LRiwZIP8VqSw5poGcJ52jOSuFWff
/2tMfBU6Y5E2T8HK4LCuHx73GyP5HyqV+hHQRLJywJ5kv0ssVb/oEvNjlbXA
mlvDsKoRrRh+vFcSGDDCU+5nm1aSRcuJnVGOL6pfSSktPl0PC5WtCUAhuMRs
O+zLRnR4thxOEcb8UbJ0QhIv2dLNQYQjd/QuvtmFjTdODjy681rUUfdNBfwm
IizPr2isIoJcTQMpDgIpU0/JXY8emNZlYOac3Bq+ZpZ5Cvlshz3lN0++c65A
FAtFpzlqpIGBBd8Z9rVLQ8vJ6ZEdkE3l8jnV/IAd0HSw8i00jrBDf+RcZbiq
Mttso6IYVy0l2C9zvzbJvarg6gALqhEkLtHRxs4+MzbaW5s94jY8re0nL8hg
lEfDe9o8hmbbTxILcSqaCteCJwwyF2AGSsKuyOQlEzJHHTNYlAXiX3cXFAi/
AJhV7B09ljXMY4dDCP7UAyq5g3Flkc5h7zV/5cV9ifY1ejiLQ1dKF+Q2S0y0
k2pPCYGnjdqsoApOnvQmL3nMZUar1jZnPHz7eet3Uh+Roz/lLjV+V+9+uDKB
kuKC14DhJ2/gyF0x9Arcz9+Gre7EZo0uYRY7vcBHPyn3kPfZ+w0nEqfGJhGB
5aZsyrIkFJ3JHaSUtTDqremjyfe8n1q2RhrSNE7zVaKlZCG17C+RfTFxRjFI
w4dXVB6rMxFs1Jrg1M1kvqTaKXaMUuMxrTUJDX6L9Pxden5eJyeScE0iPBLG
1HVKnMHavzX6fJX72y6v67Lt3flfy9tuG0s1cHchhrlaa17PKNpeS1hd+t5v
AwXGhVOFQx2R9SAUQRASCssvLr5cXEYIbUB9AjHaXtz7mhDQFoK9Oz6isAfI
VBlpDGihYEDwbjsSDD9X2b4XGMWZutgMjWuiHzAVDMSVMR51uWzKYsPG2NRc
MBvZp3AZZaZJylIuZ1JU+21dYjGFm2qGm1W1hLNPlibMGata5uKTgM7NGi/2
Tt4+xDXyKxKQzGVYC0adCx/CW4tbC9YIwwFfQTo78Wwv6GW4DxoOEyqX53a9
BmSmDbXae91T7dhac212fGUhyDcdX+cp4jtwGiHZ8q5z48qzPtn4vGR2Oc1P
3dBQ8pr5Sq9Jq7bXxqm+WrQo/NMu/C+oXTEOAEIfBGW6PWvBPD+OD9aelFAo
PS+ZAfVU2NpXLp31EJOr1KRLGaVzl43q0rYtBR/Ppz94QaoQZX4fn/f+OsNU
CUBRKOndqYuTfESHPeqcfBzvA/Tw9tySerqW9yIeL0lJYWCsqTB/H1TcT13F
1wNJkHnzYnTBtjtKRqIzZrEqbP5qwdtabCXMWeTSUWMo0B0GQ4AecYa60B6J
D8OsLWdLEpbUBwtFHYdiwlgAelEzQY0eIqv6Na3re/tb+1t14CHg+wjh+kNu
rx9q4+ovVvoH9FU89t4NuGTw33lk5O3CPXO1l5AoFlcqB/5RWVT0hRst57PK
z7rrKIAMf4TzyLx5GJL6Wz5feZd4XTyNxFTJu0bP31jzOeHjlSS8iLDZyE4Q
SPRKHrNB1v6KvwU6xCUXqQ87Hh3mxGdElsx5eNi2wfterJO8X/gzNbHWE6Sm
ddbT+WUM9DAl2+5IMhBozh58FKJsiICLFYu1jK+xlSAhoo8eZRtNwW9AWSdc
3xwRAzguLz52tAOgbzDOdP3UqT57jpmiC/5BieGPmjb4mopZXTdRIQH/qy1Y
F3mz/dLASZ6HTCLrzDTJSsGaQYVC8C0mnxiZMLLgL/YnzIwM6Pif9WSaLvGU
SmXB6ALAdWgG+5Tjz2xUXDWJwTUoJi6hl970jsDgCk+ON627FUtC6VhkJPtJ
E/kQvcEJKvJhxppvZeGpb22cu6rFPey6PxLExQH+1J+nm0JCOYUL55bMRZtl
duXqrqPPQKLEfLWmm2SEFry/Fs9EZBNYOG4uiltQdhDnxlobQUHxHxvpnoxV
8y8zYZ85LY0ujJtcp7LgdIXYjso1xydLINLDDg2lPL1GOFB+LabcCFuC34O4
Lgq3coTFIWIIv+qTP8yYbijn04rI1GOjRPbV/8ilo+OvPMyUvhLRCp6RBF6d
oO2mQvlQjsztkTpNem4PXGe9eTZDmwcO1vM16+o/O3lZTfX68dYh1QBfDDam
xndUFNFvITyQOAf6zV5W46lykUyksenJukk/JZo89yWhidpjSRRst7F8+Utj
8CjSwoeyTu50Gb/dEJWYKTMfuB+Bc3VVYJ1BklPm2vuJZ0TdYQxf5p+zWnwF
ZtPLEZTLs5hOiU7vDSjqoZtV7S2FQTKGS76ZS8gzfo1Dkt2a7wHf1JC9ylwG
0FhyESjulhx72J6kT/jplseZSf7yOEB3W1YmO1nzoBeyy6lXXau8E6CdmeN3
bhkIXnnudY37HKhw4M2/HJPhpLjYj0vZ4UE4XBXuF+KE2vySA8uzJ/wdHow/
1+cL5z2DuFGdWKikHvJOZ3MYvr9IcWGIFYxDHqsDCAxieMrulXcXuKhqJXci
EpzKvaxrDQS8hYbvf8GRISfJ+r/MJS5ot5NNZa9dQWjSJLwYue7AioEQE+sA
co/e7p7GN12Kml1yNNGL/K+GtqihCfjXWwtS9T1mlti3fdT5YLBE4SwDfDZA
C/bdUvxIsubZVNUf4w9a4NRx/A1oVqHm82wrSfXd4EOhCp9rQepT8aVrCHip
COMHJQeBKYViIpRBjnOEG0+fImQUGm2ZjCtifollry3d77KK9Wy4uz7wnBA3
GYkLtJkEgww7NFOYz+pLk9ayrvhafQnVjhFfbVv0XYfr6uFQ8hsbrFDkSqmT
zy0ALipwAG/A2SKvZ4v8l0T6eVo5SrxfILrj7fN5SMzv2nHI2sN8CY1B1zgJ
KFaII/uRL9ch+zWBq9ieChMbS3E5VfOQvtI2uZEBcoRP4YzG9wP/sn4Aqnfo
WRF1qgJzIAmQq2057bxdw1hypM1HGJ+Eb12nRh7f2FZAFCT6CzoIMNi96m6d
Bo8Pz9634jM7qdNSTpxRBOv1+aTdedDfybGMabLs7/3UsomlBZYBp6kCA5ja
vSzTJstaZ/qvlh2ACDbkmIJac7WB9pHocyswEUua5e/IWiOa0jp1LS8YcmVS
v+NTD2fDvCYvWDB7+aqPXhswkqvBLREQ28v4zdN7xHHvPrNLCXWJf/ZaOWx0
IcpHknvzrH88UNLkMiK//nAL8Y3sn2HWXG+J+m74cfMAMJS8otfjIzrKPfxG
WB3zSMj9h7KYwA0KyZYxMFY3rpxPoLGymgXvh/dsrJJaGNE3Q/u2BIo8djJO
o1K4prC4S7PiKJqmlbrpVR82sXW5AhG7zqST8B4GaMPChFGUuinC19VOjn3/
OB4PkKQ2XTHnFQe0rfS/2IuLUSH+mq/aHUH/qlSKaJU61ZA3yxBKfYgqstx1
rMpUwqipiCMFb8LNkGxOR7e/1BMhcYNGEL7eJIuN45otnwI/LM2wxDITCK+X
De050CAW3iykvm91R7JfNjonj4RQ/f04cc7sE/vBSLCMf4q9qk2rvt7Nbri7
O3x8Si68F6rDX/iq+MDviZ8qVIRXuWr1PhcHDhrK/QBeri2aBZX8+QfUhDTs
7LFHod5pjEpjxGeBdkwATxT7s/fzoaQRcoWyYYeskqfbgdu2c4pbPxBWuSbe
VDtbp9GlHjgFvYBO8ToDi0j8uAmGQU5RNoRbe+dUa6+oWXRpaz44w7O3lOsS
8Ir9AJEBvaIVFsGXVkJ3EuL3ebcj4WA80ydZHyTxDGs+YmYsuqBdR2OB76s9
1VI/9+ZE+hrO3FnCUOH0zi/IaqEmjOXzaSQaNUCnGVaowPEVhy5w+YLQElr7
sIm/TZGcu3fJGue8OT9MQv/+mm973rI0m2TA5m4zoFnoWs53f7zxVAuaSXFR
9ktDk/d85LOwrK3SZltTjqxRINlStvHPNxyEHev3y5QM5vEnd9jlcCBkBwWg
l2xrwX3JImKu5UXikpCfoYTkQPCE5WEf1Ju3gz2r+4cz3DmSIZzpahyXmcN5
89/OScAPUW8R1usccA6o81LeUNc255rWgNnxdbFbPzDUewt07D9NVod3RM+Q
o1xg79YFVo7R61fcv86ntDYSf2zmJ/GRM3nQHgPWAIZ9Dg3GnipkUT9iBJHd
txoqciOxPa9uVEqX1UHDf5Q5GTRLzXEUX0Gj84GIIn3H76ipff7hIlEePng8
j/C8x3jtzdsFYtowq9Xx0YOkMSbzjA2Y1e94glt0+qtn9Njk4DNelFDZhuGh
RmPJb4Za7zU6LGnzyTA2VIGpswFA8eOqqjrtP88wIfPbGTcPOSVP8z1m71Ou
FXIO1Iv9iEbEo7VgnF0XpZm12jY5lO0XWcHrmLLp1poqRAj365tpBjLWGcDm
TN38p41JHLs/+thdybk5BFfPz2hBk1Cfk7GWjhuaVVMi5/JKwQQgZa9A0kUf
DgFHtK5kWP2idm1pJooUiImZoA4mtlmeb1d7KesuRjcLn4XZfuC2nYX5iWwH
y/wrJzJxvEoDV1s3zD0GXa2A3blPcwPyB9otfMBEGAkwYRmJolayUbR1gEqz
wQekARutpVugXSY3Fj8gSYj3mGQvgneuBKHi/u5JepG0FPsEvbcnxO75GEXP
pdueG55hplT4+nNzfyyXNw8rblJCskGTzGVfIDeGYuqZqHv/M82+HG+eHTTK
+TDvL0MEVGD4pu3Q7lgOpGY1r2IeARn3PObSRvMhwGTvLzjXPCsU7V53dETt
M90s9qImnO352dn23E2BpKfv3RWFA+uihm5GeGiwOIA7ZfPQK7xdphoGcv+f
SN9L2rBcSPhringJWUU9zB3lP9X9nxfxu3zVhl32SHaFiWSCJGP4vbTgjSHq
5wQt2fWLzbG2ChkAGj9wfr38EYrXFMQKk5kh3lqZCaYdSrqpaVnbmOAbQt3u
LukcZFBUWXvAw8sjsXl4kMKPHlJB58zLIoM6+oaAgSxga1/+fTsiVi3lWvb9
7UjGuJW3USP7GvJ7UwCMg8Dc35oUJ9cxBZwQ4tZ7A8pdn/j+EI2t3KnEjecc
fr6TufZwaRTNy/z3C0Q+9yOvCrCOQ/WfZkO6Vunmac6pEmiOymEV+TvcMOsC
wZk+4HnwQoZzm0nHukpRgM5E9Sqgw5U9MPNE/OhF9oRpdaV0QZKjqEWxHRP2
nS6aEfotZ5kPKuBmoOnyfnmdZyDEIBsX78eFhL8/vcUxPlHwset7i2CaYe1B
ajCpnXLitiXubOToEnZzyABpIZ17OybHEiw6eFcJc7v2wBjQx++IehbLEifB
DdhzspSIF259ZzeWDmW5PNis7Eo1ZlR1y+PTGKgZQUmoJKKgVINMm/8i0lrk
+jXUR4il87UJUKQ4rK250S3BZZBK0awi2yW8gojK9ZTUu2mQwfBweRUSgG9R
4ClZQVFiKt5eu6dpZ/yy3Q8bvm0ICfbNnMU+EoN53Cm0PBR01Y7kSkCgePSY
v+jiYbIAyN6YrHq0rDDlrQGvNvDKhVgx9EAGE8Tas3X1RBgW1JHOsBPNBdML
9XPaauufAXbHLwFlS3X1eZCQCelIHp3d5ymAnPMN/wENBQx3K1UuxTXSdoA4
b+8rCMjH34lQcjj8plr+s1z5QM9z3kOtmAsHwny9nCBMAOB9iG8+QEXRBwAE
kYnV+NoumAN77JkiwZFhT9W7ucjXm5NkA7XZ9BpCblMAqpdWFB6BBCw2UNp5
Anqm+3+qkPos9j1IvLcjPsAmYP/4iXM4sH4aVw6jKRyrsSWui3dj8mDsW72E
3qoqloWOfuNK0MWrLcYABz9UsuY++poO8nCVv9JukVAS6UDnuRLk/JSBsxBu
+0PKHw+UKcKDl3s6CjuVgYDgG9Gtgz0Ri1A6klkrJpAzBkFwtQg6fwl7crQk
GXflXZ5rGxn9J+ydRFKbs6MKznmB4+w+V3dcFkep+OaEf0luMJg0JqWkFVhk
lQA6v1XrI3F7BJx5LW94CGYjqF5roAcezAXuswhwrrQMZctanrzNi0vFLy8+
X6w6gAovOehZngqglAjRe2ZrDVCqhroeCHP/Qqaf2VkbnudTPA1qIYkeYoJn
nCs9nNsxmdGW/xBhsvKFICCeLUXJxniQ1nZWB3HFyy6vApeiSyDVL3c352vt
yYstyTjMf9a0HEiqSSo86HuSyhxFnEYu1qs+6DRMlFdWxLT3oGZnisaINYez
C9kbMbD8xC85ILv/VbA4JiLCsJHatyhYCbDio8biABLP2W4nttbA7SANtcPg
lWqGIC9iJjo9O/wCeTe8iypiHYhqfnXsNJ+8RQQM6TbtlR4MwkvxpB47l7qp
36er+dAc9m36lbOmGsdgcPbDV8z60t5oPcVLrRYvDgXUS1iQBlyAXaras8nO
aJpxm0ZKG8FpMA05NS7SbvMXdKfru+dfVMLC29cmQSk6ogXqNPMf8UOfsxYv
UurcjpsOptDdX0nhl5HjF98xaQpmLP2Wye/qFDxUVIi2Z5kurwzWMQLPWxw3
HMVgYYsBE0WSvKvDFU532Vz3zwTDMWWUcOBSTLWKDl9q6BNBQDjmrLU1OP51
6Uwt5or7orRadIQQBxIxFD1EgfZzlR5i6dKBS3dOu37ouCHFB1guHmN4cvy8
lOsVrEI62ySSMfwKN8tvqI7cz+qPt11GgFZJdRQ1ouKAxbx8JZi/NhArvkyn
fRJ6nc5OxdaNojuRj3A/7w6K8mc/Y4th6FvIy+lBCtMBr/MieuCYbmsJA+7O
TrWkUQ7NWH6waDx5wIwmwyNJ/uN8GTZZzoUEi2klhdKEFxf4EnRYUNirAbgC
zyYZjCDjhKsdSD67gphuIdtVtoIBi3N2BKBoKw/kOv8tK2UTel0C/ajfCKsC
yaVAtHXB+8bwQA6MY1oTYYiP0xs5epz7kgaiTUQrvs8IBQx0vxaKnu42Pmno
OkfbiQ2plmYgNZkGIRsSJuLmR0uhm/dCM6ZG8bb9KNRi5Zdek7UEEW1CTmuF
U+UxFrPRWSabdijhxIC3bJHQ6Fp+cqJ730Eoi5LwP1mqt8MKwyE8KKPhWzML
KEwuYbr0P2VvBx2cUBWccUFvHfR4oJsrO7R2GTwhpw07mu/PpDiheIG4FJPW
8y2Ad2zGlauc/meDzxA2tXnHD8G0UvNByl4vfjIUV4C28h5OHPVj+oQlwFof
mg0CYAM6e4V2ko11az8sl2acNpLqEtS1pfb8+nJHobCDR3rzh5ZHjfBU9X28
zV6/r7DQx4I5pFlRFZk5gTHXYL0vL4TjSakJR5F4Ow8RpuzPQgYKc+6/ZAh4
tyFxX1lUHZG6xr6fS31PhXgiMy7lgnXNnMR1lN9dktbjG6Cf5YcTfymu0saB
9JZFcLgpn1s+C+UaX7YX45TMmt7ucemNYNYmtuhGYvhn/PXAwrjmbDIJgFXt
ysSUSlVH0sIU3+JYonLmCFOOcplJKuKyaM22bSzRDzGBwDKMFUrAZPv3fQLp
AvOO64zMlcCblUe4qvB7RXqZeCvPq7LeexOTaeuVmSrf/Rwv1VdMyjWs7NK6
r0jZzOJTZEzJBFM02R1epDUd+pdOQk9WajmI01oz0eCgytYC59oey9K3nklH
GYgsLLgq59gkwrrbONyIvDBAl4SvTGm+UzbXSYD/yoDX7SxLGNqUq/oAZGrQ
1dfAzrvgRVOHi4MJuqCzmPJ8oihanAwWP32L5BS1YL73obAWJxd6Wlk7QsRV
GHR+wAq6py6C0H9OhzEK/8Z/6YoZHYlaphbwNofuFtwb3+WaAb6Iv1xRNoAE
E3VWm2jM785kzQr9ncPif9dAcO4yKLQRbYPyqek0Jz9NAFRLBO5QtTEEfqhn
xlnLcLh+PQmTS0lz6+ZMFPhlr9bNmP6BA9Edcmt2TKr0x1jEzmxG2bZzbnj0
kCf4QWCP16nEkWNFgf3FuviM8ug3amsqsfJHA0TirMeoSglwtlKi7OQQvmi5
zs/HSijS8ntz20RZYVuYiZ6Z32LM9bBA9KQK+tgHL7BuLCLz77gnw7d1GqeO
RTrL4M9E/4j6ZbvAvK/mU0WmWSj4THdYgNzaaUJ0MBJ/Y0MVHsnTBzAP7r6K
SfWAdnjrbkw6j1Rlq6AHEoPdEBTTUNt+icZy752gwDyr1lmBIq4ORQn3UE6U
W1ddQGaCA8TORy6D6wQWJrLGaBzWsgB+eGLKjBhI9vIV0jxuL/lkIDV4Klk0
P3Ki4yFCCroALa5SREPsBRTZrxEy4bnAT2NYh5wNR8OFkTaFfLgF2geh/GcU
L61oJ13TNMwjtO056gD9zZxPBHqYcyRieSLS00TW9Ni0QWl7J7JyiyDbyG7P
02S30f6Cdo/qkyz+9u+tovkxsczNNNy1f82fNJtsg+rRC1D0GdGzFsSePJvJ
93ZGTCE/E95Q6uAI2BlfO5WEQl+PhAG2N5lWehyOSl0DArFdmWagthjxa0Da
NNhz9RR9iB/NGyyoKIB0QlIesFbx+XkzCINw7Gvd4EZBPjJhHJ2Sj47RgWZg
5MEhb+fA55PLQKmvXxyNpkHmTMlKHlKFq+CAckEFIWMu91Lzv6ym4akN+SPE
JTpuvEKD3FrVb2+ZykNNFX1WdITLibCtTciHKsu1miOd5BrJpSzNUKHJK/tL
ShPLPLskdgQDkegzNSRtHtDtcs0t5l1F+4OUUUNVSNrPiG9ZnNnGj7wyA6mZ
Cai9YYi2CtUONZ3KzWzMeTt5WBO0RnFVKLoWuKUMr2v6P7lr/6TJ075S/Ig+
BnzXyxXM/+x6r3FS2pe5v8yUyAzE010RgsZJlWxF4xwX+Y74XTEJJXavv7kK
ASgkVOyX/s4J6Orv7k70uIDyh7mM6jSCLHWWAUJPzhuZ1Mqy+yuXSY6XnYZM
ZVnkFLM7IXHLhHbDEy53x5y61CI6zMPKueVbbWAQz86AqIXgYvgCFlLtMfgh
Jem4R4Ba+aOjkTh+OryTYnk+W68LjVf0VFEGwuROZJ2nIGZnP3oD8InyGi0l
l23+KkifX9sf8Kapz9urxnTcMZzUTXZuSkeiWe+7QC2OUGGpl5aWxUERvclJ
h9jE+t2vywzRV7CmYRtofdr3r6Q2dXIl/A/SviNE3H5gLzIPzVcNSAqBH8VQ
98MHvfO2d9SWh5MgfNXXpsHoPPCEJ0nSIHPqRrycWUZymQaV58o4llL0ofAZ
yCC1+HMG4CenafyR+bRXP3f69QaZuzascTw03RkR0GP0gqO9Atko91J/lQkU
Z0TpkSc5nLC3SCarep1ZXhz89G6TMSgsD8h+AuwvP1vny08QbErVGLYSGqHB
ZKGbeA7dItdjIQ4/n2VTnWifh/m9k/EzNFJMy7mbmATYG+r5/WaKt/CflzRU
di/kkHLstT9obqx4aSMLetduaktyegKeJayDBlbDHDaHbBuQ+2b6xYz0CXYj
HHT3G2Ed3OMHvry/gE1BESSz9bhQGvfkugjl4BTS3Qc1llFDQ4uFfjr+F7om
KPta2kv33DvxCl+WxOkbe0s5YzLg82juW8RVGHOH9GBHzwcnEoNbij7+0yZk
bgOOLMA2gedr5SaBiAAhuaDr1kXIbu1GZYSc4xq6FVUTgUTnqstAk9Ua/Dt9
W6jJlr76dxSI8Q1dmsSQ0yKpqnGaWsPOCvDR/pLGnA+oZqXCnlfgIcviTp89
x3VOG7wHDQG5j4NZwnXAtCtpujMFPsvJEkG1sUuTHaDpEidiAuA8TM3KEz8E
wJiNQxobCc0BpuhVPTLDNPTqA5IjKRqzY7nKBQNIdRsJh54F0/ArkhW+vIWM
urGulKo1JURVIQG5OcEx4PJyChMclklr3ulHB3jCPVLfIiTex3xllaayqu36
bl6/lmYtJcTyiicknRqbi7gUjNrD609A+437WznrlIOgFsyoI0oraDjfQaTr
6wbZC0N8gFF04xjjp0pdfMMElJ7fFBRP3aH+po+pOndWUQiZS3ySbYhzEUqZ
sG+on84nzLiUP6RT6EeoGdqJ8NPE/ZPLOM9qm6/7RG7n7C5ewuf19fuuUMXB
hn3/o9lwihSSBp1j/0Ur0yEhW+V10jE9V5DNOjueN3OJaPQxIVI/N85nK/YX
pZo+trwq+8LJ+5US4zXe6DesZ8moXa5hwFfvaGPM3W77r7PR9vE4K42gC3/c
OIzn8U6NKBQ0ikilmjNKDpuqEspMf96mLDEUqtUzjS7bZKaSCOZqeTfgN5Qc
O5mRszE0hIcXswvy7mdUV2/4YTojwX1wH6pPYBBFwfxQIVXzNZZTHUAPAsBB
p7L+OFSfwaii8V4DBxwE8CRuojIsBfEn9tjwMSCq1IjbqwhSKISpkveC1RYK
0Sjr3yZ/B8LBD8t2ymXj7SvWnijmhJE3+0KS5ozlI+w4wJpheEhVkMGFlfpm
wbqGy+45l0K9mUNxM6IoiaMU0/EyNPQ68l+9fAmqWaF9z/pBN5YahznWrb3x
UgLz0WXhnSeEsP+wRPKEUsSPwjFd/VOFDtjgCbF2bpCxcI8ne3ijw09fFBh6
i5krLVk/FZmyBK3CsEphXGHeR3EIU8qLNuwSfpazPOIx4M3aQb8LALZ1QysS
6PANqzMo1gJnl6HPf6WNBtBai2km420Aw3rMKxggctWEoFFRQOb5T9BKWnt6
UHFINdxVUXb1aswYUc9s8X2/Tu14As3Gy0YE2H91260n1/HfkDbPmCJ/gwC0
FF0PNNuSas6XQri2WHVOURa3TPqZ6cEmM4TbRfQ85yd6fjycBSMFFL+6jTLP
1eB5TwCcvX3BXkWjT4r+MRtqO0dXVpwmMwRPC3de/1W5kV8oIEfDedSkVzx6
dJpB5omi++SuH2t4SNz6xiX54nCfStDv1IP4cwIE5b7fr6HQVLIz3kZgE5YG
ux5p7Zbn5VXPTTyjM9Pu86MjA/XkVNJHAX9s5SiurYuP3ER5j5BavA9om9Qa
WCyDF1y2yDNuw+OReDUOiyWcq9hSqACkvrZgeqx9raWadiXgr8/GgqNxYIWB
mALHnb2IYrPELKpRgIVBMz1Mo0SWTNtCFLPfY0vHse8qgosjyheuvNlTvzFR
0SMg4HuXBamN3PrZHT1Oso3HYQUUF5AVVNETjzYzcgcifDqknUWMJabooQ2c
qw6woc5fmwOoDGyZSBy0tuVIhsqEMwbYk5di4fD81sFATRhnB/wAaMJgwhYH
mcw18nmjW8UoIal9eAOkeizxiFekM4R+kccdmpCbv5BlEMzKgQEy7+fw4iwb
UOvq2Jm3FcgEI4MH06CpsyAzrqjgy8aFqXeWnqw332wghRXDgSR5rjx/+TSz
kU1bM0Za1dZ+zFwCVvRIR4PJ0Zj/vuTb8JL58jgowE3UTV0XBVDBI3czG7FP
+L1HZg3P0mtITCaWZenUypvrIerrCAG/lsgBx0dBZr5JQd/iRmWa9xqGn4CW
XGgkzuvopIN8uiCZLshfRmTYNcw2ZCslz0UvdZodht2O7fFFlIhGHaeln9Xw
GJg8EFMI9xD+YFxOl6oSLnBBjLLDVI+mHuWlBtjPzuHuFv/IJfytKZIkBfwj
8oRz2bHcLSLvVVcIDz6LXkuMQojnoTm9mm6XzZnjvXq03rJbT3oF9I3qdvUq
mK9X2cTEQ2Vtegd+WWFHfU8NwwhNidBptXtzTw+eaTZ5vYMYX1qiR1WYqbb4
iqQyinol/itUFhox/keUAj4GbvUohhzLcqA/Wqj3iQkew3kUcOIUaiNURC1E
46TjVv/hw/c6lBMox+j6ucPueHdqrZ7x2gl5WVxuKN49KaAULiO4BlNIfw5z
I+YPdI+pEVABgVH+xYnXidsU99d5Bw0+jIIdMBkmp01FtSwrlUNGzS6bly8s
kMUkgvuV+o1RtpF/nx0MuzhVuCI2PvKGwMaTeLLYw0qlH4A88Gs1cjAFuIK+
YRrUUWZnNgDOXhHLLEHAhAc9C+WFai6IrNEEXj/CnZ2yJt/KQODzEiSlsLDM
F4ZFJK1zOtn4jTlNTOHrhxDEdxyNAHsKVWkq/FV3BfiptriC+7f3lbpOE2KA
KaouwmXCOc48QIGDve0sJChR+MYyd8EzvsWU0Z2jihIYGAZPjgGqksThRZzM
fbgMhjoaANSNS7daNv+9MG+niX/RuJhxToWoUUsr158EOeyiBU3X2DgCXMV2
9ELsJogVN0KHkPhpZMAzAbRNDuyWrvHH6g877ZZ5Qw40Jsd1xVrW2ccjodkJ
8GUJf4UVHqNS2cWILi372xw7VWPaW+N1zBx0+Om4Wtyro5HGTbpaIk4fMX6q
hIpLOl1Evv9bsojZJFkNqmXnENftHmS2x7VVTl6Dm+euBhIX9p9hhGKy2DTa
HPw4QjIXBDTu43c2/SuoUErFFrmsDw+b/47gq+2P6qhKZTw8pwwv3n9n8yb2
lHdBwYLMkf3QmDuUPF2GpcbgslGA+gK/H4qf54k1IfspglaXXxByyt7ja4XV
cReImRlNKcL9u+MbzDGVAaYdESMZICj95/84pKgTM+2Imy0A00TeZmVJ6+tu
wlyDbESoL05JuqAz6ZseHNMx6j1SpxLtVQbboSI6Aqq81Qs6tFtzqg4Ptj1m
n78vlux1CsaayaQcxGszJLF6TS9XSzt8I9VZb7bUt6NMECFXnwYIuT21UgFb
2s/QthDWgARc+Uh7S2RpVHs2Un4I7Ezkkk6O/QKTN4Sf9vg2ubFSwKylnnez
RA7qg7reGjg3KrtrYhby8VVCGC/hz3MZsQ9VCbVUbTcg5piZ1olyE5XVjiC+
w9VJkE9FLxZl+05f020CuL5fKhZSt9xDrMfk1rn8jk6AFuoO96L2fNe7tXoq
YoOMTvI3k9NXEnCye3cKsosYcsuYRc6Rgq9dCIf+lel6AyvLDoUtB8h7t3LI
oR7/f7ZKyFMSMVQWLSHddbt54KTOnraV5MWSwo0mp3KVyUGoZas71KaxCP3t
ekh/xuWRJJZUGY+h+9FXWqe4LCVzuXBPTT+GM/a3Wx+L2d0VjAHL/eda4wGG
+9adCT2NBinFYtoVNxhD/0ZtRPG/qgWiwnWLczJLG1HYBSH4F0atc9VFkQzF
/co3ERWRREJnDYqO8qt9hIK3GBKhigzyA8m/HD8qKgBLIpY5LymBVdYhIxQj
5f9F9zpIzke2vIOmr1lRA/k7DPwwzHScjtj7AczM1vHD8VrW75U4JJcwbuA+
dM9A/RL6AM5HqSv/tMAmH3rMuurhzvG9tA+gk/fPos2nrElmWDBKiLAn/GGV
dTMyzST/wACWYXmrM+aKr3Yp9GbIJiPXCiAtntyAyCDbSxOjmVOw/ZOrTLQ5
OOzWD12mJQRWjOz94VMKrTki1VoIBXaKiLoGoqXTxN0DrJgENgJHhcwR3QKV
1g0t6nc9KvB8/C3wib3Nbjtrmbe/pgy8RGTxulhtwg52dP0eJWmxaD7qyEvq
VweGObU72h00uh8vqbZVouYUuQHdf1SMPV95++BB1dr11+Dw/zcnaB/DFU8o
f3bsGap7QuoHD7wkAO2e4z6LCUdRAsNaIa+gxfLsGoNGbKaAEHT08+RBhABG
0gm4NlDC25UPMguEFU62k1/ab7oRdP9EjFgaaN9vQzJR69fNw3ZBrCcOOdcR
0vPuWqZ+vl8GeCSSSvDGR2d33dw4DrJ6i3YwSyjghrRjjGqa3ensWJ7SgX7q
vvg6yKGVN7Dn6O0J+A1W9oZisIHf/XvFsWgbml3LaUfpgE6fuWW2rqocmtPF
T2wi51O86TF1ni0n+wWD4UTBm6csqUMS0RzQwKD8dgqcarQSXtJ1c747LDPv
yhTm+3OlsM1nzTAkTXnu2KwC684xuWUlBbai7RSOSsiriR0+CrMKcnCyKWVI
KUUiC3EyD/I3Z/pXhSSn55OSnYfCpwcqt+0wOIf7unFN1zBqoiUq6IKiL+NT
r9qRIk1YAUF9fxos2JyZ3I5IDwR8rAKWy81sLe2K9KR1JdhFXEXgtCtYhxsY
id/SHGDkdTb601P/9qqc62JdL4pnk4suUX11OS7GLIXpomiwshkgNDLfqG9Z
07BZDbNjuvAJAo0utBgfS0Z7+BvRD9J/6t8li/D1gciM1A6SBS05KMjiVNXM
XjmWAGB+ZJHB9gqrbUaiDD5piqrAmnQ1ClDz/f6yhvQjwud1yv2r8Q0H4eyQ
lFwFsPIpomK6XYnAR2XvQo5cCaEOvSnPLSrbqCXwiav+/avtVeA7CnRuR2Ms
84Wj176hU9O4vFekkAIsl20nHLbyhXCkNJjm49GRdEPBplS/G/iaNCiYNYg4
3NffEfIs6SqN/6KY6ZZchh/03jn+fr0v/Aak8DWRgJzqVvKhjVblsvEIlON4
abavru7dLLShlphrEM21XsSHlTlNkOLi8yuUmQF1t2IkdUBdIXoZlmTZoG7Z
wxtvvMJ3RtGUk6FPb88YpkOQDcvqKNtaj77ijWS9s43MaMyn/Hl3fP3u80ZU
wbpbyudOIqootNoqEt7BsLY1zxFwQ4ZEgazqdP27cX1JByq/XwWOM0N0m29R
KM+Jp4cKeFHNLAfR8BzPrI/UYHc7rLZBt/XeDLJIQikcD4f4pyyD2wmH9eNb
6Pwe9fRQBU4DYHeXYDWyhOWkazSCSyZlN3s4BhqVGaX8v3i2wFXjVE6dwH5u
v+4SnYb2MHPcID/bKEyfl0x4MfSmz1R4O1rNVh8b0iORaJI302L1Vo1nO9ad
F82VA48uh56iIN2nZmjAL8QVJ6AUhdyR+QJKd0LAhpsGLwDzAAd0JGgEDfFN
hR0c7oZ9vrv7N5RhTzqhyCsrWvYSNlzGX1gnQo7jdWPI6vOnVDz+kF/M5V1a
RwzzuZL7vGGv6A3wXzIzJM1fRO8kHIW3pBCiwyKY2oyYboVU4vkTvn9Z1HRw
3xU+WhGhk25d4KtVrdhx0Xc0GvdkRkjEZeDysVPOHIlKxpJoRT7PaYfUBINB
A3Si2wxhLnF4PRqTHBKZKA8WZjlQMojYU1DPGP0H883G1ZOUriU3ORa0jhDM
o44koEiCmVz1V4vC3726+L5tiu4Ox4fu6mF2kgJbZfVkHjUlFD88RGsB4PBT
TbYI/OrzVKNPkDwh37Kelnqig1hIkV6faD1evPdkI+h6yNxCwv2hDWNRRcDo
b6DyYItPoisY0znHVGVTxv6QYgAh1w7/jYPqRz8xciLX75kPea6ZZXGAT9W3
Bs13mmTUVpvPD4iB4aWgLJRCnFbSk9IpvEGd19TERKoiaLsbDk9j5ufHdNvg
2KaTod3ORz04iVnq4Unhg6/pjQi3bqzt+VaqT7Mhebde1C4Oj1jvGRCLX+pT
VlImz9BwmZo2ieYNbZk7HVvx53K1EsWe7NJYvOADqM1eRVLf5HNIpP1O+yOs
WGtxt6oa0JB+c2p2n/mYmZ17IYeual2eMEcADRmaqp4Ul9wIpQQ+xEzu4MLE
lcu64U1JY2UL1JCHENP3q2wvodfl00mUIzKBB38KPshW49c9LmBzyWJiidXw
SsuRDwijXp0fEjMlKMWIMWwTaDrIvD3qK0OgLS2Fx7Mt1kxzTJoP6qdYre66
+8XvziyB+kL/PcGl3qH6Fsjj5h8JXtjowuX8MeDXC3yjdyGl4a7ORILGucTW
idkWTeenpcLF0Cq05k3KL8MQlBmj/GGroePLoCE50ThJVvxobmXgVbonrWl6
i2O6atgHiGWpvNKH4mefK2e0FZY+vn0OJvdjJnn5WrxJnYe8s9oXdNPH30xY
JFZizFzBAw359phjjeP31kmNW232rnfeYpuXSGyq6cZkPl3lPU68RvX5TkyD
3XLN0bIO1vGMUVwpbHgkjtt/IdJoVw5I667Y16eSEkLBS/m+tP4KsXT8Txdr
n3oN7lIMk/3k0NVKwWV6qpOpiUNmOevAgD7ypOjpqcKZqb9ODdDdOzEN95hv
zvrdLc7D39hJJjdmChmu4CkDuJxeZwQqKAXshAaWBmMbM2658y+n/rshCi1C
1bO5H6NUmVR6WD8tM3k4OHj+Cavs7pcc59gIsJAWqLqR9Avp5eKxcaeQ9feH
AvUzhaHnyJJ0dPWF2GhnfMXi9rOmfQ508bOCSNZqPxEqCdHgmJdHH3HsBefX
FzY/pcJHjIWkfhUVX1TPCINzjFbN9m/TMJk/BN+oqg4mPuYT8AiHN7rl3szk
WLIUKsrQozC8Han+PjopdFLYSEVqCJtrSPMQ79+6QBG3Ik8kF7f62TRDD1u4
yexdfvcZIgYBqXdfNu9fFGuzAnNX5oTwBTiFSkprrZUxBgoQipeyi6NNw9LO
AqKGeyItjUgr37pHfIHuHwFDn0LYpDVVurbh3/EwIeJzSS2ecrhD9WgUyWSO
0n0jdT2GNxh9qm8gyCRT6nC0LNKUpTTi5kDz1vJbRCUtYmzKacluHGHiUaMV
wn3rOBXJlHuEbWEEROqE2DgOklkT7gzT8d13PFooWBIOqhQuwTmq+4y9bmsW
PTdXm+OvYaBvqz4gyaoqk0dry8u54kCGHcEwBNnlIbe/iaibmQNzzhfLw2tK
FQpIbbUsfNMGKzzfHAx9PZRUXMP9Y8ftgRb4g9yV2Bhg/IyRhXpbT/gJGwh6
nwPwaBmCY+053+q4ifX9Cr8qJHTU+qME6xbbbqUXhIng+81Xb07fc3LcI5g0
ia8RY85mTo5urB1yF8y9TR9qVQBJhXW1Dx2qR35iVP4G9pqy/z29N/ZrS41G
kauV1jhsrAI76BJ2zPC9nwR0kxmOmuwam7bbg4voc6ENrn3LDhqUeUl+ltMM
h8+723aFrUrtQZlzljrZe1EyCFIr95/BKMA97oL3xp8KriHcFnTgkLUqiGSk
EFAnPyOAXO09gvdWikth75MrqFTRpF7AaX0rE1say5ukXPsKvpggxIfRRhki
mLhJmePUKilmes2CAnPn41N8Ztztz/HpOLChRNsAPdZ/JTmT97suuTXvdpan
OWfIEpUaiB1tNhX3byRCTswpicaYE8YFmplpa+0pHQnegIOK3qfOMwGINoPz
5T4QFoIrgyiyzHnXpzJ79MMx/cRy3rdpMn8C27ks5lEn+SgA0c2rH9o6O8+7
BIpETWG9ZViQRjWx6BEP4CeTu0S3tJ3/6hOH6r8iTwEtcADaLT6S+c9NDzgt
7ZILMk+/8XQzGDwe24VSWWpZm/Vd9NueWiuN/ZKwY/3utghCxpI+av4Wz32b
5Bz4jZ62e3+X8Du1nB33IkqkOB85kWbxH2GnVJuDQK9oB196O5QNK2PExnMV
a7U5vRBkA4rJ94m/e0tdJz19fk1HaoY0GyAAvkK3CwyjBwfc2KvsSAUsmHmw
1CAqNpqFszgJCGwxpfU6Y3Fy2ry2taIYSRzVaqGikvJ/Sc11KTCCyJUeQZcE
1AyKL1Zip9a0ZQFKFctecuUe4KUe5i/wR7Rzutd0BGdH+GUwinSMyw9oyVl2
CnlsOXoxcB6sgMvpNcQP2nrrKM9pHV6oFAPJq2SbB9vVoGiVaWZW3wtYcgQm
atjGsDW21R6mFWyDEL6zew4RHF2LlKttzoEC7mhlKuGopxYB5glEYDzEeN7L
lt5jrgL0fxBFmJuaiDynbsjAO4jJYI8bLQxAIe6RGFLsIUb6tkYT68ZGut/V
HHt4V7O0+yS9PTqi3OCq4PpQb3TvdSiPtnWrnGg1naAwAGSGvC7RyCnLuecU
0euyCz7cWHMWU151Dh0DpomQIzm3Pub4u6HkM9LA0YHhVqXEYqdh1PMh1t6K
nrv5zcC09xqVcYJ6xtA2QC3raVVMeH/dWWSmgfaK59J3ZniOAazP6sasK46h
W1YN4l9FNs+ecOrDeEVRo3yx4Wy1Drlwvl12FZunh9xQkoxF76mWCS0qJybU
bHvdD9lda1Vbg0a189G9dKuzMM0FI2kaPDzlxgEKxxNJ/5pH6yfvcm74no4n
xjteGWaFa3bUkTaxkhQYlWZuwrp5H8lBmQVCzrY+aILgz8ZWxnTD3nYf5nUc
D9j6C3fMFw5a96gdj/k5ueRW/kzl2jvR54xurRU7kStfkZG/qo1PqaT+LfdD
3FiA9nAe4XYym6ylBhbz3CPFfa1NCFZhgbsxofrC0FMq+CHJ/C3MYa4CXbgc
bo+uvvQ5WTJuEEDAzogY5b1YnmPbztGS02JsQ18R9rtLqFBR1ASBJSWJh18o
P/Ti3sOg0wZsH9Di8Ub3hqFhqRUmDfKQZEjoI6KegKWjgeG0sPrKLIRzBfa/
f5hDZkGAQFavDYyMYRfDRWEm7WRMgcmq0HcLOLEWKyCp9VcoWTeVx5zMUo01
8sHuC1mCpfjT7In81D73dQdBCtGzVOZy9qfTe5akeklbbP6LWL7k3fR+mQqp
UXSBmXCcItM+fXXMErTpND+dsCshjibtNjdCh+B+l9hXKxeyn+F+hQWckJ5a
xCOfP9fiquvaIb0H6Uuq9kTFaQ/hudIWQuWOCU/j9gpE1+qyrkYztD/6t/dz
8SNopoQ/pgxLOob9NQi5v16LuvtxE0MGc7f59BZFHB8JqL2PP1Qtgho6zyLh
SFpjJAnJdsnhEH0ZuOs2OD5pNT7cMLyQ6nYrZvPrtikYoW15ekrncUoblHFE
yfhTVfRCiu59of+xhC6WlWQX5tZg7e45ueyXN518pK0q+SqmsyfpMVlFALlZ
5U7ZtYxaQ5nckIjhl3xEwb2FTALNVnGKRquyt+a3pFmNFWUXdbIIjAF6epwH
PP1O8VaeIyX7wC4W9flWhtpZ3MzWn2+hhTuntVMk4v4VcwCMQF5B44RQFks2
0UZV1JhjOOT6fr0lMstUm8wH7wvnoWyLI7hypfQTacemyCBVrlo2HQeKMrix
TnbL7M80XZdGDqH5pAZzo/HeV0Ks+r2VDNuPlkv0M7NRf/g7zjDFfJA8NqoA
VYqdo1MjmIaZ5LmWaQdzJGm5UYg5SuHbwqJx+0dBLLrABs25ulsZjDisMvoh
1Zozc6ydYViZDlmsl29UirWLPoI9LdTO21fLHPS3f2STp9ub6d+xNWCOfooN
+PmYehyk4x7usUbI0SXd2JlbREgCHku9xhH+MahJk5mycLLClf7NZJeI0laE
oarsppEAdv5+aze68XJCyZMfOjSrvOmB5oM6222Mc7CkzZSLWbitEqpc4OTD
jGaOLH5X+GeY5xGDbiO8ZJCIB8eJ0eVKS7RhI81fGd81UhjTCnGtGR5bl7A2
vLvaNcLgzGJJdzb5M7IOvqTA1QaBB8sdwGQ28q1z33BoTkRErVq9m27tU/90
q2FTPmMSgIqawjYfupt7nt1SrL6atpA2rh1Ec9FRf/ogmyJaS/XK9GmIHu2Y
aSEj0wfSrfD1sREfYYALcx4sJHweW2LjHFP16C2NCvzOt1yDiij61JoqKWZK
tOiiJGon8l9ZbJL3AIMm7XVY/WyRMXOEZm/KYITaGmm1r1fd9vAJnZcqXmGp
V2eIlfgfLq1N9WPeBBNBPRcrho6OkpP4jPAWqqSWZbbKAH/e2cbrLi5BDvhM
rLQvKYvR7QVjLaXWYT7MhK8lgjqc5Pk2TV+Rk2qTJ0ZLCzrbSeSP4IP2E80W
JX6WZ/x/omQT2nBJlBOkvnb/o5g6FjcZhcIrIbZowTxepP1EjnHH4NB1J1MT
6E9+mKA9He4vxCEnbYRj+NCwnnaSsoYhFzbu5hLdOaTwNPjAX+2bGujAl4As
tBvUzWjMrj8nJOweWN2lkRXjiGrtVe2ZYC6DLT+a/nh/0ASIMfXcCo/zY6pV
/b7qMjtXWpt+qlaQ5efwVg9LApE70wc+EVZLVPZ++VZBaO6Dbdn5NNidwedn
rQrtXNSTx6IcBl21JurJbyEoDH1k1cv0ZA1rrrht9LRwPKegD37JYETdtwG9
oGCvByWLxUgryMIlT0RXkvqtCn35elzaEegb4euoDuxd5cRJpEJwnJHkCxlH
pQ2v4aOXsJTNPfjxKqDofckt5t/K3O0b2R0iKdfy8Dvnch4TiLrqquN7bfle
uU27/rQvXDvzl4SZ1uvkml4rIhP+xAScfX+ItAcgLLY9ktNTyWC3JUvmKAr3
+0P2kOFLRQZKGYjUSs9yI/bJWT2cbLIfsrz+IejZ6atGPRmrPgG6T+odZYiG
03+Qh7KZ4I1hGq9Jb8dxMFyw3v3qZyVuiOilA/DkLydqe3sLmvOui54Kl2NH
M3W3Z+5+9IIh+kf8IrBq9V8I9geoPUfF5qWJd/encDzvhKIBA7Yc+FwWJWkU
QiKPw3YCU9+FwZxiCJxJ70CGDJG07mejNnPq6+FEqdEMMylyT4PXia1Xo/L0
sdhozgkRD960dhpkdkwbR5nz+m9c2WzpUWDTXgYYbmYg64sxDRWNVBiEJmyT
Bt/eebn0OHtJNgqfWkACGeCESlZ+1o5wmLyAWEfiW8cBeR38KZkhfTBYJeXp
/GE3UjUdW/TofNky8CJw1aM7cLpVpigs3fNLUlNYvjYOjYXmDwWQslkUq1Kc
KxqrwjIZdmphEkta48G+Mf9zIsf8Poib4iP34gcmJJcu4mOjC0lF2MTdtqjN
1nVVzii8snq1nh90AK6xVJF68y6NX516xnn2U/GzFqvms7rtcudtO6u2K+A3
UxXL5SxxKtLrsVAjDCvZ8bOPSmsc7ZIJ4NmSkLHU9nVO0O6iKq+M6RLud86Q
4kpYaCEw0xFyBt4E9/3hmL5OQMtaujf8c6bFn/g7BKnd1/xhhnbFr6kzmety
1r978Sf5XtV6qTuKKi0DRl1Cw4PKvZJyLwjJzEWXqnuWhcH/Iac3eM+IqpMS
g0RQQDUCwvWbioOH09hZRcTTWoOFjee9QztNG5Tf0TJ5uy7GOVmUGtwXl9Kj
f484zvvFQAgRGwStJ00lugUkvtXzFTT3EU79liEKanmv37c78tx9EvS3nIgC
RQCd51Fr9XZDgV3O7z73QpECIHDUG/ydROhy9GCfqIB2SGMn8J/onJRQD0RP
WM3BvvvdbJEI2Dz+rKScUkzyo4CI8ty+naIrwScLQRFgXKMGGu0hRUmZVjOP
IAnBouwxnWqKFXroCt3JIDMEbU5sWbjH17gZCgAXWjeirLgppemKDdeHG5RI
l+bkhKmxpMF7P4JVcMUHm9lXf1rXruiJcJUw0+8iN2Gi8Xo3IknpaeUhenqo
r8yTazMFF5CX+6WCyA7GGX38p9ITS+NG6Q5tnM/oUm/xJEMk9qdKsTdtODFJ
W5Dv/Z8otAf3RHX/YLztEWBby1YoZzwDyZ8ypeAbZArJ7zyLHh45fYCB79iI
G79Gb2HBfjmy2yo4tB1qcH/t9SncElHo92Uus113tV3NuWMrpU55g2pVwE4F
fcPZwXo41vslby9KA4rV6nlFBYhZX1myZQZ3wW5WTeK+QCcgUI5MAXzDH0/8
fTlTrCFIwETn9syQAbe80UXfP/LvX08n0ivoXmxa2PLg8JskKjryMREsfPBf
OehMV8LLMeBbfSv4VbYQ/INuQS+Z6fPrxWQGO5YKQ1P7ffyFRSEzNPOHM8Ld
gIm2T6Fd/CO9wa6QmhrhEc4K5ENz62gMU/McxzfKbgp9T/HetFO9+qnG2L+Y
57axC/UahS/tgTe1inTpF4L4Dc/q3UwUzZb4XQgtahr5OL3v48hT0J+yo0RA
QH+BV7gkKizjw2aADYYclw9CTNsNaNaa+KvzfZhASJzZb6m5xYejftSMvpXF
Y/L/RFEQUcwinDokUPx7eZULqvaVsxgKUVxkAIP8xm2XP40tZsw+F0m1/Y5f
0X6zcRBNKoXT9rFgem3NpOq+z4dS5Fv3e6N56p/kHRZK7nqi6+7KMy8a8fcK
n9mVQUWIdNxRnhsiik+DJsN2zCO6m5JF8Cz0cgWRttUTKqkL/ZOcjEv/9H9G
pPyMlvGmIGy4yLn2rXX45rgMMhaqkZ74ZGmQRCRSKPAQiZzTnRMI4SeK0KyN
yj0VZ7ESIBThbAuPiBKAeUQqHzY9Q8TV0QAHXHzOxiMNpHJCE7425n+uVx4J
dUwbcMr5oYPn/VV9XcYdUQ49adwWU+YbLbOrWVLQR/z4bnX4MDRoxilOH4XR
ywewV9K7ztHk7HxRD8CSjb3qFwQVBLQFIZWCq1xgt307uOO3GWawpnXb7GMV
cGdag1T3v17yrqiMPpyHB6raaaPufzKjLrwYC7yB57/dcghZKxetEB8jQBWM
2Ay84CAiBuXPuS+7M4yFYb3Kee1RFnB/JXnCBkpn0JIuse0F+ctvZZ86SlzV
HcjL4olWZXvpu2NAeIZhWOy8fIYcFTbLjz7FQqtJCdmS7nyEGdH8kdZ3G7Vf
5fLX3SyBYZPazLYEt++66q5vg1P04i2+dvv9ncF8PjvMMOQuDufHGMAtj1Qp
MzuzoRmiGrARCWkEyS5cbh2ZYx8BXaaFti9rVbPgnKqKAOJRMzhaTXjXFewn
pvLIsuTobHGdk6lAO1eYGBzx+3ig1J77QcrAsuJKi3zkKZVEcpcRLLHt3fWf
mfPOqnKr9v0j+cZl2Q3o02EjJuwAzgpCLxcAsr809k186rGmCC3vxBfICwbL
5ro7qJN9zKiNOwLhGvXqZL9ezNtf7LRSjBrMES9ECI6ELO6cmfs7GUpD23Nv
fs5Gsp/cJszrIb8bx0y7ZCy9Vh+xT7AaOL1arfNWE9nj1y1BTagbFRTRi38r
900k4P2VbEw8iRzRLRTgrkXtmAvA1yQoXmfPrCBGjzCGLVOW43RC4MUw7vIe
OioC6779mpF5lI1pkJZ6ceowW4QXtuH0c4wGb90D9Qrk2UWOU3Mox/xj6Jy7
fdW4q+AC9bva+bFol+44hFoV+mDL6Pqeg6CQhsFefFTCsvu+JEutaKeO4s/4
pf6h/fXasq/BlajPq/rYlvZ4AAEy4r83clOaofM+Nt8ZmHZj5PFJbrU7W9cV
Bore+fXuLctcGdbmfCRA/2N361DgRTXi+2atZWCweYGK/7uzrblo4QsTp+gT
yHOa8IFT1Tabls6TeB8nW5es2esNGqspNHMJcEUMXjealLBMbgQq1mbPp+JP
6g2+vSpQUS1U8Yn4Grd1gvWEUx15OXxW3Jx3t0YgCtBrrhzVVmY77qbbjfXw
Iq4TF+sDP6crkxpNv0MVXyAXhYEbvI9M1DjZRKlWXHZ3ug3odGuyVcpNGjGA
LNmSyDWj9JUXuFbv07n6z/e0LK5Pns4cIfIljfAC/2DIAOhZbs1vLEZ9z6z0
PdnZrz9Qcvw/K8s2j+6XoXhmOukVCOvdRoL/UejMUqhIttsBCYlpst+dL7iI
NyHK78zUIK/bULmrUsi3Ch0VtkJ0FLjQbiNfhA335d7qAf4hhiSFDdBDtHkq
QFA0A/MSh6kLcsnN7BN42kAwNscdOdFY32FP129xYJ4jbObcek7yOmrxByra
yiNEYX9e0+JNNB3eqkQAvMjBP9C0xeCrXWSTlj3p0vHg6+i9Aie5WL1BNRLH
g6LpDMz/cA2jO3l9Pal9OCWin83rr+R5f8OhceowL5zKFqhWel7m+/niEAoa
9YpKX/K1//aHT2Xfgjq57+HYKJS9yboor3fwNMmEuJqEdNcnnFoIjbTMXP+m
a4Wz7+aAGaTnJgJ7ST3IOxdNo3vNHBdXlNHnkKCyLTsMbBmV4puMy8mZ+uhQ
m5wCohBbkToVQj96TqUpdfQSUvw+XMWmLSLU70SQKbGV2nDT80g68DQbY9lI
ku+XJoeFYGwHEJXD1r8JIUzyoFIUos74eIQziO0CYyTzVOHbYCcBkQpbmVDs
ed47X11x/padHYws2vq1g4l61KXg9vQEqMyLWhuhf8QWeKi3JRHqBf3ceiIN
FMejERRj6nOlbFwA2RcR8JuGxlPdUqDTswWXFSBVto5MxEPKToMfrhGhvJkj
jSwsf0zGMemTCiHSvRsNiqVwpW/mLTujj7iu7hGLcK71AO3tBtwJ1fFjyWjQ
iTcSujVBof5C4iqo7YAxDHFUQV5XW9HWleJO0xrlrusJ/pxSpLU/VSXNUbuE
QXC2hcpxlXYsl13TpC0/PG+jCLSrm1Xd9gNAM5MGdcB2c9ND3PBVRye297wH
zJrux0LullQ7S4QCRBp5OuVdHzlnevQ7DvnaWqEvKLx28S0SB+oEO1I6tu/B
2x7A3WPX+bxzQoy1q6F4LcFGAuHrxXbZKAgWUAky/DG7V2nyO5RRCz04Skq6
l+5sfgpEuzMkNloTvKKSA71CxEyyhgiXPKa2LXrD9rKGkq75h7A2vn9DJ0W6
i2Tme8aYLZj+FCFoKk49ZC9AEnhKcK8YVQ1s9qK8rC2bPTI9pKvjezI42BvM
ZZLIPJWWhmeaAyLGsRzYtHCy3qCB5mmZVZR5irrQJKG7jHcuMsmsOWU3TMj6
kM9jsVJjLnI8gaRVC68rNjHwour0ilWzzxTkW/7XuB0BbAxjn8Fkxbnh+HJ6
WFLycLCZHJa7ilz5fYk9MNffyMREj9iLKN3h5qcYyTwY6Z7l0a51vmNpSwPZ
KX5AcmgST1HCqnVG4zvfrIoHxHYShhBhDilianYxQXDzH4g+hB5xVXG7ga/R
D90EHstf7XXQFEVRRx76X1cDi044Zr/EVeT9GN3vDVCPoR9LbbezkCSze3ow
iSxrKfPI3YXdbH0k/zZVjCi/ihdmTtoIhU+gqFx+czxF9VdTI1YJT0efw6WT
5/rLJuHLiMg5/PRMg2OzJdcMr9i4051nq8FnYBLbM9kEdQqeD0mG4GJXO3mS
98U1i42qYfee/a8FMYin/DscH9z6nt/HA24Xn6Fa+9Ghsfr+EFvq0xVXr8FH
J1vXn58taKfulfVX2vnvJH0L5ZCxIz0QDGdtU/wsj5uySZpND3tfc0NyiN6+
pdn0NzsNc4pXqDfb1K64P38sYlmy7jTROgFVOV18alnAuUUoSF6sbzwzT2hq
9ub7KzkVkRbjw49Sl0paOLIf9GUmsc2ApFTrjtv8bObs8W3tAaKBEep2MraP
WQftKeRe5/ooBfzHXMNfAVPxJX/rDnIVZyQto52FkqMHORS+WwjEJd344F3T
yVwvTrdZu7b0esokiSzaN5/u44q5mlm93jOUJ8lEne82zNft+Zgab1zKkU8g
11Akd7Sql4OZLTq00jqk1MPSvYMxtRQCdj5y5mpfQC6nSlJlrEKyBiTokU1S
YUXKr9XQs9P6/Pedf4hPqty2wfWMZwudRJtdVml5h75zjqwWuhCWO4+LVUyt
3gctf0jPEgYXEbvhTWAUL/6Mo5WBGtlAUwyri0XwwVmKFCNV0aFFpmsRhMea
EVoq2M+TOIVrFWioslnTBhQin+Ru81umcn4Tzdx1Lcou92FkqgjGKqo0HHuq
htpZyg3QQ+ptf3BZZzmg0016imCUnRg+LYrSawDCnFb0lfNkZ9Tk0jyFe6EV
0FmYqhBA2LMxwMwUTb0SZ6AZjStggII1tTcT70o8ebBStzSdT9D+FVpe1y9O
vb2woY6kc8NSz3hQJ3CX9Gf03lyqOP/39V1laUTm1UXmS8yWRwvXJ4MDpYau
fDHq+xo18NJuP4NoadzpLTtPyb0R2aiIbR4TqQM5AYTpFZ9WqpN8zuR91XOR
3WfldyxQ8A6hh+tUNo6oKH+axTSxaudLIzEurq8JlwJR4yvGaYpDGVFob2fe
giVDDQysEml5xo5I5PnJ4OzV7MRnUJZIV+ssTYKG1oidjWZsG0d2oXTFVQKl
o+05NovuGBbTm2PcoTg/qydmkpCj3ztTKFqWxvOOTRY3YEz6XInGoDsPZPMx
dbDX/vWZyFRnPsEzEk395OURnDX/GJgyAlNnQ/n679XdI9V/ZGNb5FR7gEp/
PVCzaIvnayIfXmFTjMwR2PHIx9SsdxfOwK29en+PlN804zOFkouodcE9fr/r
c5PZyCk3uRVddA3p2G/jXWLWBYFvWMJtieFAEEB1D+dAXizfS8Ht7o0qRv71
z2kRiQEQLtNy7lXiyX7xQxQZBFedXU3TcSkAXwSS7mB07lIiXaPYHbSpEJap
XqHli1dd9CDX0LwiD+qMYHgkgfD9CviTjPq25kkbXbJ/5zWfnNPtd25/phGf
vFEADap+31wODFlYoPDyQ1ioNGjj+kvzJMPcmiGrb9wlFP2Kgs2j71C5jgmZ
+23QlTQy8O76++u9fTuPXjgVtWM6BMTeXDbynVizjcznHdF8vmSwXTn58Hzo
Vj6zZG47/7Dp6kQm7YVPBl0UXO9yRzHmVcpxZj3VIp83+MkjvMW8N3d3sHTn
Lp4MNEqPJogY2eHLMBsobg7/YSrCB6ciFIg9hgRehOnLrwSN6zHuKaXxeQNy
bxou8cuHWuxyKHuA3IKgwnb5vMc5wzvvPQ4cAkK0XC4a3JBk0kjZY0QSVvGw
Vp3bEwDpcrUE9ttiH9polV5z4N0blDNBrL0pCYO54G0f0gq+AZA3y337SWMb
74/uDSeWz9DOi0LFuBGEMlkM2H6bpDT2n+KIciB2W6Ah8yXVzmQqdICQfnqa
ckMtfYKktzBeA6YzcE4FV5KUJbSIA1VtFBR/a08Ff+C34g1KVJrs42y0Iax7
ahGanwEcaMmVW36J3aH7Sysx8oNInAnSVML0DxRgFDTG21YYlOsX6yVHa5ud
j8s14WTxdVdORYLwtiHZMIIlgo2bC7eAkMDX7naiXuh9ZrljpUHdQ0+8oWu5
IBn9B72N4tDfwhK26sdioFGwTHr7wJIEalTvXhhC5y/M/3i5KrbWEb3JGeSg
8SeVBukJcIIB6WpGY5lyM64SCKTdMHR7OjXYTj943SLxqHw1DWn+GrCN1VX9
2QbiR0ZWraLIzDq6qJtE6ouE6bUbDx5EtGFiMCkO8JbizAPFZGKmHeFLIXIe
3DjdXSKCxyqus4dn6FShTd6Ef10vnzK39zGGnXNC9+zg368nCkehdA3nKZl3
0eBXMZn7c/F5+OAaa+lMvm88DsGcz57IC72vOETei14overwTlGZ8Pqhk9r4
PCtHj2qtxVTzYQIhZlox6BXIYc5fVnsnaHqwGG5a7x4VmOsgx3mOGma4FEnj
pXB+IxACcyC4vtRqXe6IlywzHAApqDG/poFXwWOOROgAehzWjzKSBV1+aXeJ
HPNpEznn/3PoqNSw4W6ZIxXQyBmtiQiebCwekHWto3wAhyFfRTJ8LQjoUkjX
zU9KAqImAakyXafgUV5ZwOHOWNL0fSYhHx4tGg39ACnoPDKJdmxuXhl7Z2EB
Rv2sqSkaL1Gz4Y6KfnO19OEEMQQE6MuVrULvBOML7C7sV9UIcxPA1Hpfsulg
E9qJ/FOM4rb5gn/G7HVdeaE2uMWg64SjPT9v7SZfyrf/ocWxuU7FpVEmtuCh
djm4ycQj0oMevo8ECcmyGgWwAMdkpbpI7atAvjVzGi32sm+4OUL4J797LajL
Yw3vUlRl0orvMiFbSZ0013mxq31RxsQjop0ITWi/chC9NebT5ujozweVbbi5
BhJZtLcGdaqCh8n4I3s8zgcpZcKkVsJxqExm3TAM79anPQUpsFjsQZSAIaNa
b7Gz9/ucQXNtZpTx20ihAadp+62VKAVEBVt3oaDhIJtxW7my+upCddt0wuTP
s4UcheO472OjpteGG7+2TqNYwUznl8xD6KQaBDet6rJXQ5wkocbPY1ftsI+T
KADyxLFKbj1CNRr5LqBwvxTcIeAUPcHf6TSxPPo3cmLuoYRZzYJs2qCeaGWD
Bssr/SX2AZn1uKsua5kp3QLua6vdtneANQoaAFYlN/Jm6ItGR1x5fwy1mIFR
N2w47bfVxlNtePUmpViEhAO83Qhm8zDvxgkUsDYShrYyMUj8l59Rvc7larn2
D7Ql8mKttkR/ODkcuofYy0lypsudbewXB4ROqSI+BVoSuldJYkgFwaIdCO/2
edGKe3Cxu+D1TsN+RXjHmFsy7g7ttuSOpZiuJufjpnNdsxmkh8kIDq1rhz7Y
LFvrogeD95RXLdwuZKBGiOlA236qzmuMLxJhTrZFPMNTtLXU81V9bxUH9XU/
sooAIVqVAYJZFI67F9y2bzbSUrraY2RpwIO2WsN+PyQar4CYVgocDGEYC3Wy
8xSioPX2FLMNYD6e8pZv5eLr/bg6vKmKy85c2ybtg6DDvYcscqgClmrlCD0D
ZY4sLdRVfR4QWZR/ht8yvHAabR19IhcTY6PfxDbMK6/l7wF3rGw7WWK41SQ4
+H1Goc4OVpxyiZ+yYFL8TMjncOhhryNCnvfhLvPnollUiDVpCq7ek7iwqCrv
TAY82547TYLNtzv9uRN4PAkeb1PSB5iLKiUJ+4N5a9sH/EWGJ+mikl6A59nS
TP4hAL1EdpPK7HZB4W1aGfQdhzuu8QEQs4LK87VRtxg4seZt11+SouPIWMP+
iRVeIgDqeEUszE/pzorPQMO1YWvVQsxgMwV9qTEZL41K+1dgBce5uxf8nbwO
J+pRnxMCTJ9Asdat/44KMzmtJMLATaQ3To7iHNWWbtyDpwDuzI5+SVZlbBEa
NuQNGo+tioylIosLtXCmptqCuEcPe+e7IUa6I+6pGl3TTzxHea6S5eUhCtiV
GjWV8Vsb5JG9/hG/+EJMB/dH7oB1hHWjOKTQggWSABq4zHYvGuLM3KuAB7Hi
ps6SakOFJyOa3v0Cj1TYG5xooMR9nniWURbSkV4+IAzrWRVhofcC4PmWgUbm
INpe9VnKWsHQVPJs7UbLexBEwdLdHC+SGqgeMGzlJD+HlGqboFeLLp+olXp5
bmd8yoJjOqxh8K2Trbwn9RUvuk8Dj8ZE6MxYaqfY70CwYkL4g9Bi+qwXWc5D
QQGnfxC9JBqWuduqRO6Z5YZl/Mz6kDJrWUk8q3h55oxtADrD/ps2XaGqXNke
yxlG29OeqfypPoYrQ0oOlqQxPnHH8zsnc+M1rLWTtQsuUA92ig4jpXWhHx5t
7OMfExWnazhahS4MrIag+FD3mNUDMhwunRLzI+K+BzotSlkDVfy93/pw/Rro
+hXPYckiPF3eZdx40BC08IuTc6owkBlku9uxSOFjumpDoFSGXGIFedPoFqMW
Qts935h48x6l5WHhqciFILCeiZ/BYhLvD61Um2FJWKicXEQsHpfreKtyTP+4
Q1xCPaBCpvcVi0TlZwj5dFW3hvPGaQtnwJG4HPVCB59aiN2QCSncAkeOeg4J
VgGyVMv9zWandXX0IbQjZLePbnEvtBc01s6bR+TEJE2crEqNKjvkPC86cWEj
mlQKIzB+P+mekLD1Om3IQHGXi8X2bUjwxvrgxxLENBoIKmsmD5sA6C8cJDbR
GGySLcy+RzAknMBRE4LX/Xp75YGMenO0FTv7i1G7D4oGldD+B/V/BlNTZyrS
MKCJuqQDgF0uNrNl/tJjcDn08YPuYxcLME4szc6JtGiAQmxAq2ghbDg0DJew
6uDwSt2fJaIHdj/hxOBH/Sbf1xAeZ8Wr7O98o1BDCikvkfeBRH/Cfno/H5QI
PejZcMOeyJZhl+0UvuQ08p1xp6dsJ+yXtFQRUHXy0/E74urC7fTpJBUvI4Am
qR8yK1EA4oILgjKG+j7kFIThsJEJJozoDxFCaER2YI9XimJX/QchUYMosQTv
LKMCAbYL5Zw4xMR7YdLt/cSATX6bSr3pKzR6VRryz3xm7CnHVN8g3i+6wrZ/
dL0F95GMySED54SzUKSkQVkc+kLOrVzwOyAY8klGzy7Vg+uPxoThqRTI6mnn
wLn/Ss10YWOlnOPLShjcggQbcgVe5+KPBrI1uPRndMRLseSFCD+GI9ZQTKPD
VS8qtPOc24veoll7abRmWQeNPNjOrZl+BvaJFzIFdTv0FG5gWrj7UU8xKYJp
ch7YjzVlehUdbb1UslSixYQr5IdWn2fE9FAiDjXJox3/qwucw8xs0wCWI/aU
M/Sapy8u/RAdGGQy5NXuO9g5jyPWJxfR/4I8g/D36sNg647EdGXA3Wm19fUC
bmftHpEiCm3tiUB7Lben2Rnq7NpDMcUB83UthRn0ZZXPSyyoLLibrl6Xqxu4
+OUgfCir/SkB246UJp5GGd3FuQOWm6BWO8U5fR0OhHuRUGJku6Fo+7xRY3dp
E9Y8n6KateBpPXDei8AHAFgeAoHtqpusv9IaZzBOucwC2w1tuIWSsvIZU1n8
XoJ6ZXRCRUM2VFP7Jtn4XwQMtM0944YEeMv3tY5J3l9ENY99LFKGo8yXVb/j
bLAC/dUpe9/mKOP6+kPvvAI5HdriX8egof0CE13HDMvX/7LDmdm9h3m7D2fO
hdZV/TLQhM0JQCGVE8C3CCnfuoGQrxmQXdUPCX+eld0c/nJ3Eymbfdp4J3lT
z14jM2ojwC8rzB/KWLapS7ZW/p+eKhLwDLvhObDY3KlzXsJ7f0whLywU1ho7
PpZvRggWVAtv41ADgmmjnHWMRIaDfpsBtp3klMgAGtTYPTSdLxqc6Jf9GGgr
6j9wjZXIWSu2OH9pc8/vmDC/SYoTkhxOYBBaRMdO6IdzEH2rnzBXJINFBIBw
9g+Yp9GjiXHqleIDGAXLcdrHvrvsch0IJQUB60vmNU5KbwW/cMsCsyPLu22a
zZbfHXdloYpHfy7Yglj6955ZUzne70VeJmq1AlbvScY+x2wUBq5zu7Rj5dM0
RDX8W8IR/yUd0WrTYYWNJezwRXHwz1VZmwlNQmQ3pPU2dXJw4o/cMFSlgJQJ
4gRnhyX19NOR26W28xj9DUkKXRzyrnYJ3RPBNbouEBk4UOvHC/hm+gWGDuor
yU5wutPQp1ZB7TuAYo0v5XQyIJPb/q4lSetVydc54U6X4tVprsBMMejFJWok
ACeplHF0kSbV2EdBEn3qm5MIrKwLgZEYlHoQW3Nk5gyfThEdXj5M+yRVbD6x
RQNzyfoWGtj/YdlDZp/40ZZ7HebjWGvESErSskjsCU6mGWqySkshPVD1xQzl
ORYWQbtgkYuAjOSfMr0fVcllGGTdyUNESV6zVL4XT7ih2Oq64c1kh4CEMdGt
gQPhodWruBBcYepSXos9ZrE6Mt4E2Ok0sJ4fAMYIup64wi18d3PW86pk3mmT
fRYsvjEDo+9NdMvd+9h8D+mpk59J9Mv34GUoAO1IttbwJYjfKU/F/MOeCtp+
wbJWYJloc8vsbm1MYBEo8SXsZ5ih0XW9pSGm7/9t6T4FPpWTAOewVuZDpePy
XjEz3x9QqNrEQuP4mnyuXOg5f82pBO/4VGmZYZwfMEelVoTXjKYnu4RcqdFn
gDDyTvUb3m/5tSsqoieKzDuXUV0JnlFcWb0ZWAOF7oxm9PCD2HGaGEnLgU6k
CQHZrlyRSmH1jLPw7JNjllpsjLWZ6izc0qLgXZURhik65EK3yBFmH4svSsLa
Vc2sDGqGygB7CYofzA5CgPkPF0OGmb3eVCLiSbqMt7TSUdpn4akPE/dFR/LP
wyUh3oj/Z/3dh0aPn8BlVaALycEhoCDDsFQNtxvDgvjdj3lspQGGkel24Nx7
CRSOfr29lBEDJ7ScncRYLAk2opiV8f+i9Qpj9mamKw6C71UyI8dgB9aTuukG
nKG84VMzwkZo+hVgzyPUI01uKPsp2FkqSWxrGm2ggwR2QOFrTuxT+HLsWMQf
CYxbFU0XrUkA2QYwYP+pIWOdkhTFusiwsK5xjAIiqTqYoSW5F0/uOYOfxqwn
XBdUFOF2mmue3u9dRm9o+2ogmDvCjxZgdaJN7IhN061dmDBxkehgh4/rItdc
RKFSjUbtd+Y2LbMmBTroeUiIqS5S3XAu0CTtMET6wuPhY7rw9pUey2w3MptR
o537PHcW0CHj4g61H1IxtexrQr72Ld9ES7Jmza8Xyhv69knY+KZBhUJJ8fRH
rA62O/00DcgI57PxKPPic/9bwHtK4XZgpxxJi/ZQHJ5vEXo/uaFnaH+bEyEv
STJLcfVeNcn3N2+0DLnw88fd64LqOcjLe+sHL9LcgIecyl5puyOUiniROapx
C/L6T7Jamnlw6VGq/jtGKXt5CgMWpNd38EH/YMbo4YBUH5AuOp0JoUqUYc0V
0h+/fjYZMgVxtm6OhNOLs8irohksrOS0UyGHE2ta4EsGpvB43YyYvbXEkm20
1SBhr4IsCx8Wcx538V9vJWZaA/GOqu0u7DCOhsV6KCx64gET1ThNcjqYenvp
7gXn91n3PHjRYa8jAa5LEHbH361i2yjfPW2LzPev3aI6iKGeG6RxHJpGXKd9
zHuk7pEvJUOdbgCu5YCqJwR5Rkw8HkqpZwCZe0IyPU9TDR9JqJdUPRaUKizq
9nL0THBgEZpDAJXAal9F3WwlE7eqLSyPxAnY89xSdhsE3LVoRjGoCR3WcsFl
pkH0FYxyGNY8piDvPNPSPhMohF4cwYMd8FVngvkRp2DvNbuTQN+Y3KvW2DKF
nP1IPahn1CYt1/cDKhJ9nH9IV/t66EmBe6m8CQQ9AUBRhXJSBogoy92sG2l+
QiCfM49vYat0eROwawrZRv6rLt2pJ5vayxmUjUVz1BlZMgNYUKj5s/ttQ/h2
c1GOk0bSHKej2lBrXuXnGNFIrSXkKkBonr0JNHfnG1oz2dmAe25KpcToZZzd
WyCLoBSRL5i9hfgT3CMlkw4mUT9a3pgct3NLtWmX5nGo5FmTGpPSoDxkPzHJ
ehJxZRoMAWFeSSvCK0mpeIzne8i8Xx8gGjcOWS+WH0La2QP6FoQhBzIYEQ6E
PHEE+LGHz9P1GiEZOlE7Lk0z8hOuYJHhzjC35gQ+IXV9wyzrB+rjszydIs/T
gTW1hrD//+g0s5DWH0L6U7dfJt24RzsVotzjkDmtd14ec2mWRN/sVwqrTzj8
I+Q7O6CraW7m6+IeI1L6F47lm8hKe4Kkh0xq9FilKmqa4RJsmQ4S1Eb6Sw1M
9eSBfqTfxhS2aByKkSOVkc1yRTG707wwFCpxjqc52rqoQhHahv4Cu+7fWYMV
tUeMHWwb6TB9Mxr+kcKgzeLlJjEfIjAF4IQ+ryvZ9QSgtZpusqqsiC8quVOE
HScdD4C0E27JEzjtvFUiNKpvBuBFS0b/K04I+gj+hXwEwNx1ntv7uWdMIRHv
e/LKWi//zpT2cQ3mdEVZUYUZ5JRZIugdmx6D557M1yDM+KSGKnDhHlWVK3Ei
1TcpMO7okib5G4XVSul51B0YMTnUtCQXqfy2QpraP3CexwpeDe7sr2DIRX9o
IXW8qO+klghuqBS8nSZLgmDeEx3JOZAVdPiE0YJmoHu4It7w/saFjZye11S5
pkCDnjWLZjx704aBvmhaoZNj3kY8jun1+u3bF6vsOQGepAbb2+k7BDl9vgAt
zf9zhEzMEK4Qa1iG/OtiPR6T1xH4axYxGp/CjJOhtGHZUKiaKWWzXoZ9QO+U
4iYXVB2TC3wQ+AgwxRPTefhVrTKr7HeO7mIMUUaiYlzGHuge/8k/XzPAdotq
ZhoAk8R7zzPurndB702UJj+9vjtynxyuk53v2LGHKjooKEGD6KDQmhDjFr6R
reaQDttPxxGAP9LWtovjgBp45g2LzLrL3xDkZfpP5nJErKEURBypFWYIErL7
tHLhXTPvhr+GeAVHgHz/BtBQ5fu8K/f9nmI6P2YadnDlBwpKsmnb6c4kYlay
yGK7PqRB5X98RK59ratt35BZANGSliNYJs4ZAhVlnHbhJdcis01nK24969fy
1L/TKN3IaKESgObgpYWC0ljdcpAXEvPXtjdc0Rs81Syqad+UdnEXvgB4CyTW
KsiN0bYCSQGZVmsPg1Hh9SeIcU5+QiZ0M4n8QPqVIEVGPaRV14bEIv2mZrPB
mZMkAw0xuxbcoAM2dgC1w44ZujscCpIZpzSkkcRHZlgpj+1n5fGSc/g2A5rh
k86Xb8DiYrW/+G+9Dq2nZBnBXpiSfYQFhiO6xEgoSzkcfhT9EhtYpcBDzlfE
jp4DyZmOE2ysU++B1XMzg0yuiiU09FJHRzeaRIKTMlTA+BNIgJnk6bXSaKfK
EnrcQ0vcOWHz/T/1AyOYDDn0gLdlezSkfc8himHJWDDEwBOpUdGb9R3MwHQI
cUzRZJZ0ZqiXwwz99lrGmr/rL2Gl4wmDd34/arehTpm6lRJ71XgVbZocBZo6
kIYo6z9cjEFCjr6G5SkZVEUhWgs6494OU7J/Y7x5tmpyKY5qmd5aNJ5IQXiy
ICVSGBO5zSPDHelpsjh3PxVi9y3DfH7InGizizc9U9G6NM/AMlnWryGkyJN6
O2uWGxQRx1Iu8axM+F48v8EzXEnqKC3aiTliy5ONcBWHLEXID5fIA8baq1/U
t1UQ84OwXh+si8/y3te1iw4vKJBtULCFKuE/D5Zg9+svVtX2sX0AkNVspQGc
bZlt4o2onAshwDcHFUnzTgNCeAcFWxVeFoL/XwFaZ1GuJllZ5EzCxtsTKXgV
Ah+ia459HabnFfxQDfeb70iJrxW66nVhsIk5HJXf+0+SChItgVHUaKzaffbn
xKFnAASp2+fvQZWDY/4b2xLbsg3aO7EhfgtRfhHWiyyu9E/Olg/2JdTBYp3/
6hv4n/bAt3f+eYXXeN/n/tiY+TAHobf0cJ4gOHscsLk6N9DQQeq9SpC19lym
CvtbGJ499UMFstH7X+OFGSYLN/UhZKmQF2pLXEeNImFwcXeI7m8sPlR3eJ6N
O08WePpMrPnLIWqY4oUx5yx7y02my8TFEQ9XFfd42MRUcyG6+qjAWcGY3NKZ
sdhvuFEFWnL99+qsbuUdqVoMBqmfZKdY2KvQwM97HG8e+jPiO+UlHu7f2qBT
HxydAFQinAVZIUtineP5uOwGUpzaZm5D0K1KCUdwfs6Jl996lsvOvujIgF+q
wiyg6GuiAyaSIVG1P3RkV8Cz7Gmuyo5VarTpToYT6vmQqRf3AD+8N3esdydd
2Sk2hxyjIH/kA9pcNzzyXB4HbXBShrIF+ACCemdYsYUbyKPRGD9fWeNu1Orb
F39ctyh1gReZbNKoboo5LAsthCzm7bMfPMHO2iRKDERRXOVKhfaCMSlN7IUK
XpdTDjtmBkSvmvzNViEthalwraooirdxjtntO09zbkJAsESTozHVSVOJNkP4
yfW75IpLwJXHCzeYxogRwssVBDW/GFXYj7928TfL6frdMaKpkTT0/pvB0ZZC
z9QBjnf5Z6IGwmuEttFQci1KPMqW4/0Wz52/1HUvlT7IWKWFrq+GSIBf91wE
uVW3W63z3pgYMclWDMoOy/BjiRruCVxQKmXYm+jBPpF0ZwjLgWYuBXkTfAxN
uPRM6BMIOE/bFIeYr+Owz//ucP5O98svZmtHI+OJjtRB4StNvIEFSEkScSkd
68B3mBr/9UDOyNnBNFW4tvpIu/7p57Qdec4+Kxnkn0r7ZBUmDGA47LpOczje
ZFeNQVCO7jtA93zYFnKNakk10jSWelPZjiiy6ysTIj+MdfVRY/95QWGKPjoQ
inHy0bHeweyHezLUdaIyQiLlZ9Nuokr4kaqmlv+T+aO8RXtu4WYYZ3mw1omX
q9zXzRz5v48wLhlL8gm01iMrJ5G4MW5awJC7O6WuJJX3BwF2y8As72pCkfsU
m1Q6e2bf4b4QcmL1bRwewlpXHX2kZP/Ht2skouFtBhtzsW43IwOz/N/Tm1lc
IxLcKVs1EvbTCOS0T7u1GNYMfH/JOXSkaqWqCnlmFJzJwr7B0GNXHwa4fRbA
sVB9m0E4CVzmLRpqE/0EyfKk5f2Ltdzb4oSsJC9BKevYw0/yeu6X+32b7bbW
lxkuRJ/uBhpcALic2ZpSTQxWMQ9fOy5VgwOhORyrsbnytIddvMI5m8cGatMH
SPlYXNpfDwrPj+iu6TgRriHkXBsggs7bGAu5j/kvADZlKWg/GtAFvSopQ0kJ
wzkvbIzkL2IRnDohr94zHkgfoLM2O6TfPSTni+zIGDhV5oTjUfyhnxPhnbSy
jDPvYKJTnls5gg23BFz1sEXpp6XkLo0QeCxiT+OHc1gy398AC9AlersgM/2N
0wW+zMLCEvDDuIOFsqC53JeZIH5K6VeLhp+PdW+1FWpS7zq6hh6Jujceu+pB
wdOCH2OtbGE9nlrCAloU6XAVChtCq2Flr9KaEwI1RLVKpYVvR7Jk23iNIfbq
r0tOcwr0usIxIo8p4q72KfSxszNKt/8bWBmK5lyAPUSlTxmEpKjEhw+97lF6
XUQ1rU7b23r1OFAi4xP5yfy1AHXTSWguYCVG++ij/g5Xg8mHT5PAemvydTLc
2fpAY0lobowViPeHxp6zfP/y0wC7aeRIS/OZwXih3E6BVQGE053qo6sIpX91
Zmm96BFZS2BjGQpaL4p+9zq2s8cEuqUHoT0E/QlQgdcisjIaKziQnKzUl3aL
c3GmU0ZIOxUNJjeqNBxsZen50aGW/C3XODF+MBy1P/IuGKLhWB/V2NKpq9tk
17gx0SeH6WjZyP3HT0OjlcGcaMu1rXcq6cdOtsgl1JSVUkZAk035sn5RGhlA
3P+UqfXWUuhSJ48orTKG9qBMakgDr2YHa4ifQvvUEnNA3+0eemjTmczrW72B
yyQ3/tuPfXMO5uqPs7SPw62QqKBlnO0TxR8l8PDl1aSRU3zd9Ov3G8EICbtn
0YdNuteF91DVgPX6DPNoa5SYVpcTGIQtD8sh+b6E6RmMnVlZnlTQeiXhFdUy
6ZiM8/LJ+uxP12Ng58AeHaTkzq1Pta0HWO8UQWREBql/NgIfTONVWnCVMUns
WhE4cjRmi7sIevu0UoGq4A+Rke+siIYrrcXasm/p4z2UQ7lCr27bNQSx1CPV
OLy0Qq5Xct/EdrmPNf73qp1rFAX/vs3GXbJ4pIgyTHHsYQ4iplGiLFYnn9dh
pShdceoAZp7C+SAgsEaeaeKcgfL83c8xK82iRyHNX/z5fch1EngEr4oryWdl
W2gASCBNuj4kgbzO7B085ZAF8Dxzw/2YqS+CmNR4GphWERb7wV3y9EcjkIvn
cicgmxXNYjj89J95QO+5Kw0xAVZH437fr3JU6rqT0v+qoXKTKlWEJsVtfvrf
IEc72JuP137TKy/7lBHkkn8cJeqYrDUkGggPMF5bJuD29XWzROY3jAEsMGHk
sInWiwvs4UH0PuoGYVeAjYR6oSodeaFRCbINWYFchRuWHrLQhxfn4ey8k3he
YUtlI/Vl9gOHJrB6ci0e3rF+csDoCrx+/xT0Mkr8BREida8VdOsAyLV4yAz4
/XSrj2G0yvrwSEZ9x+fWDOaEcDZpciIQ+tQZ0Ka0mHNsKgjof3aYzfkMhzAg
UPV/X61srkadfM7RZ9t4tQqQngFc1hzvReBOY0lajkEH7r6K4vKgJKSJd7KE
FNOxxYQGW/0qS8UdF1oqrezRN3KLrOh6pdJyXFYcQsU1a3M5wsdGMkQyK2LP
BfCr1AR4D4qZpLzdKt8j9TObJPwbQJG/XlgeXgQfaGft/yWAcuElLPaX2H1W
eyFLmh3ReBsFS4fxvKJNFo7I4pN1XdP4a2wpgLTO/qg7RUs3UlDu4yPZTyiE
aQj6XTV4qehhZBKSei9xFz5heXuGtVxHYQl9Xbm9kBc1GNZG/n1ACn6eu9ty
3Yrqu/E+j6HTLgGhcSLqTgnV8RZ+0ebbu4Yyt+xW6PImHBuA38DRHfHID17b
TlmZjMwvXeRWE6x0uBmXVH3g6TsLuS/pMMBmz5uXUP07v0mkGf42KjM1Aj1D
ijsZVGpUm7wtxz0FaZZWVHO1SVuU7w1kRaJWhKE/2Nri0P0T7QIR9eUQBicT
GVoLOg64PIs/78fFr0sbgyGyxk0SwXHZm7ziVJvUiPJhqddVe5KfjbA2Lto5
THy2LdiT/0nVK+dhWnIbKiK7fJv5zW2IOGD72aSgLfJYa2FYqB6pWBWz1zAz
lLcprSyNCDKBDgmXVSmmuJpedB3dHd1G+EBjOSBbPjN0OSC5sDtlY4jLp2NP
OlceZ5WRh6tYsdAHWYlF1TXbY3zbV7kNGFgzyv7MfAzvM7h+0yRY2I0dVRw+
vL1Ptt00COriefx3Tmb4l3hJqzA3qaxd2ORa8sykdatKYgzu1iDcqti5xGAT
owawhvBXpnyhFeO9KieLeu/GQhb4r7U4C99w2osrlTw6Pk8AWRVr1KJSdL3j
gQ300fl84I1Pogt2PFtP5ZqJPKYgnq79VFNwmG3rKhaPVur0fJ6bqZgNvZOd
IpI0BR1ehuhRAnGp/iWE6Qt3u+Q10zS5c8TG/Y2dA53iAgtiwlKH7HPuU8j0
eF2hREZnT8CO9zQjXnScZtsDG+Wjp7dC8xZOcjslbGfaNX7Etyt0FcOE5g/S
2vaacz+s2bYa/DJ2Z0eO/0xzkbJzVrNeetypNPY3l/ZL/APTskkU73gMe7aZ
YTDpRXhgH0PVl25Y5vFUkKC9/DkYde7nf1nxc1a7KhcFuzA0rAOhNCllcv8F
q8bPnw/CK1b1zuXmhFIx6PMWM2wV7gf/JIUVKuJLt3ENF9A8sZJeEov4kxUZ
qc6IHIgexi1YlYPACykPw37oLZTpe87TC6dpXXFr7/kY37E8jZtTXi1tmZak
wMHhjBGBapDU9cxaDvk3NOTZeCbVLqNed/CQHdNJa7Mn3dQ3iGZQYJWCU+et
KqGCVVWOTyhmEG8mtWCYNDpZhwJQbnUoIj0RmGHLN3ki0r1PLisDm1A5KvxK
C+R86HYEALJkS/uyoPO4bT7H64Kwy+L0JtkUShWZ4kwZvX5jQuolx5hwO9RY
wZZJdrtMYWbSp5VSrDIO+FGLAxYuEKd5NVG79bsO+ODnMolzNBCCGw8Polry
joDbZwHeiEZ8F7q/6rA2sQlde1Z2ZUDqO24kl71JHJjUHT4XBrPloDP7quY2
ZkRaHwh5VZyViMc9y5U4v+uM33f/6I5yRtLy9efosSI/FqmzvFsgH8iiTIx/
FHSxqYVxpckypmkKnXLxAhlETNoX0a+Hipa3Xk6wAIw1LrXqpkH6aAniWvAn
qLKb+FrXW+xsKMRCkP9OCnY0eQQPzGSmp4J8V5XcOOdpk9+ArxlZI0puI+mC
r0Ov3oYQUjWKKX1ihbavW7rneifnlDhj0KhaAEESPk2qzufvQ+IMxnU3GGJo
paA7REuNN0ykpoHX2WXFHzU/FhfdBN6N+xENknc2oyeKZm9YCj+hQU7kpwBe
mXZBVdYkpwiYp+56YYYSNlbAQTQScniwZ2OtwhHuGIkI59A118Wf8392njzC
ElivN/G/nhogYFF9GU1YS4Msq7SHjblAoRbeU3qbRadQ5KlyemuJLsT7kZZz
HfBo7Gdomb+Gs39bDFBYOWLDt756ONhsUT+toDiHh19I5j18Ab2/mBzDx1n3
H8O0xY50Gn/HXbHTDqzpHFn/6/u+q8zptHeOuXn/1+7sM1Az8gyLVgDGhAwk
xSrcdDNYu2BgA32InXiUT6F4AJqObHIjz/nS2l/mLTk/GQyQpxf+BprdaBZ6
LWirlSzQndosdzJp9yAMOEFG6YapzIr1whW2RRZ/JNx0t2kPtb6C3fyouVtV
Mx7y7cjUYh1/l/yX1PBvtDYhyZ09JYvWRggQNIdGiyIB9ye0dLLwjXX86RDy
XBuzOEhV3kT7fHdaScN4Nx4UM+Z+1PyrCasdzhvt+aa1ij0T9eefTDv/U/0j
IHUKsYr8jdhERBTVHg8h1iCBi3JpaYemTY3kuzGigZ9MDdLJCZ7fImXMA1Pp
UkIVQMz5gYEBd7vkJMmXn2apVhkJsVOIimPZql67otN7ti+bSiS3yEAjdJAF
RGcuV02bPT4g2bKFKuGux16O/5tVqsntiMLBvlP2QglthQjsonHABR0/lXBR
kpxwTEyEvvtelMn7F6JVUBkr0u2YlZEX28cVTbvQ+3hqf8r2YWmcJPDTvKmw
KmwKwrmurd1ohMFvm1qAAyF72qRbhth2W/CWlH9/N+ie8c3sGhQg8O757e8e
GmwKXMquc5Jk22l+WfViFC6qhw/2oSZgAxXvxE7E9WizENH/U9/77F7m/Gvz
p/hBQdKlYcEEC7EvASpy5Atczrx7BSmpk+tY6jyoZS+GZH1rUmj8WnCw31X4
XLZcgJC5KR5uXegl7o7b0z0cV0yDipCNG/mGoroVo2xDhezPzjlUGT2TfwMf
PNgI/GBrNhW7aJbnhBeOuw29AFEXbJUV4q5c3d+6dija9NRQwIYTgnE1bfLD
yiHiOCWQbFqDmbW77H8TN3iZKL2euFkgHbu590WcVQKNCVmZFYl04/40lwRQ
24jiXEeffBDP+FbTkg123Jpy/+m+JDn6inry2hk++LIv5f1PW2TCAfB26mz8
qDvo/l2QHGESuD3L6dLCsZot5KERyh569+x+d7Ff7fixmHUOVieAVekq7Qxb
9woiUqNb2vBRm9HyeTtpR9y16Pw07FNg3tIezPLtNEVir5AzNSmeINPtztfF
K+R5lXNp7lU+6jO4q2qJk6YVpRd5gglTGIoPWnvNJhz2H4LMlYsuW4A1+7Jg
TJjP1vj93Vc4ydnLdM4DZ3gkRcVRr+OxYoDXQ08moR0zHQM1XLdnBvlsFLgx
oewvLj0aXTl2Eai9uyDw2YkTJcqRgNkl7jVrb/V8F4OPk1MRLc6jr3JR3f9p
dtnDov3x99MufcGeiwmd4Kju57MosEkYLGR8d9vuO3DJUgVvsg0vbzyng7M4
BGs6VmeksScXNVTomxhXqceqIWV88GtwwpvZabKNkT2As346NaK30qwSblWy
cxNQ4Em+PbCvq4cnMJSd2oQrCQzhdRBHg+TRI0YsEh0ogbOCLCRUJdol6wjg
YfZ+F/DW8HxereO2azPDzzv97lk6vMNjF3P1k2mZlmmE0t2KGDbIkzPnWg9V
NIW92SAbN0b9HfWdotSiQ29TNrSY1jSg+sRJy6w5Qnb+Dt/xgxTgNC1xjc50
lYPzu9TCJa1DAqT8E4fN/LAvFHTDmQnKIX1cyh2YnjT78Ua/I63nw0pPbJbP
KPMzLUYHWfR7wmqfkVCRmQBZkTqg0XB9rKfdiqCD/T4o6RWHdkSZWgK/vycW
3WoVqaqtNynCOJ+eAsHPAe3tvaRR+V0RwLLrz6IpzR4dC8dZVCJA6lZBkUef
H0n1MzVfgLpaY5Gbg9ysrOmrqHqOCwlxw7wE91xFDLwyvXmD6MDLIXAuQ0On
TASBkk89nrkyVpxvD6igT5OotXTQs0fVv3zRvx+PxSDdytGL/eWMmAzKkL43
k/ueJ8O/nK+CGXoZ7oTeBJKHjTMQTPbWbJh+ZrXRCwEh8rRQxfnDEiSqbkGF
Vo8dJaJuXK28EAZf23GHYIgx3EkULwCfUIqVGC9jvo3mlazANVYJWkQM6icy
IJdtgX/h8o+eRV24lYelr2oyOp7dTNlSrXA7d72XJsenakeZmxf79vAfbOoB
N+/9yAzDEEtmCBcxTb5H8K/I6/M8qYMtzBXjNlfHE1jkNBdNhMX8XA/vAoiD
q4SGnDoiftCTKxtCst49DUZu/QqYsUZybe3MHrMdxuU5vwIVgCBYdwRTS1hr
8Hq6hKJSn4FBO0CXTXtttPnI6PIc4C1Q4I6lh90omKpbOsLVgxr7y8hSafup
Gr0b8/PgSyiDL4sAlt3AZSQhjqSexBXkWmsKjSroN9ddOv8oWH5iZYqspaj6
b+VJg03kDHKW4fNVsCXvMFXzYlRGxV6nJbAAUJqXTNeZW94tMaiegqcVOcxO
usbnKow5w8ynWcHRJjtu8cDTU43kGj7dITyw8XEChIKiKvFm5qLOTYOka+eg
qO6XkToua8mTGiQprqz1Q/zbVXG616R9ljYVVRq6NpaoLIyViR+uSl5tZhYg
UMOyNI8R528a2h2nW+9PDo9gvGvL5CLY3MvZyfrjhnE7IIRskxmj0JsiYjL7
CbITCKGns3O2ZQbEz+PrWQzWYHP+gxS0w8pcwmX3d3GmGDA4VpHE1ZhH1qWq
mRa3IkHpT7X3MRrhzlKnFoxyw3roh4l93HxaEZ1C3ya7QkS/4014ohUghmtw
wSkYkCt7ttTcJd9cUtypAel8jb38cYR1orU6sIWEUGIktJl7XwMfBoo00gwC
HOtnJzSaUeh9BvMEZf0faT/amspmPBadvF+pwGbVzRh6dvYth/d0UxCBH+9G
pUYwhbP4/dtlyKWFFTO9ImKj9488e8U6e4oAF0oi3gIfYfHBXlPtOKb0szUp
bKAv3UYo1vWJHad5M0/Zpu6/dwoQdAXVUd9z7pHohly+rQoOsSL2T1m5pSNU
MIVCXWbA26JCCSNbvCi17UFRK72lwwml08Ph0StHAPLSXJ6ZVOB/3y5zwI50
F5kxaxDo11A5zmo3caVy2/qJH8fanoqnsbhl7cIYeOh64ub3pyijIM9Hixn4
sOWF14/vrwworNschIj+CHbVhBo1vbJDcJlP0qnK5xkniLFbxtUk6GKB8tNE
yzjUxatfur6DIqPLd2MAtLo8WZWflPJTZdCv3wQ5XLb+fFCr2KhzwYUuTlcB
hryISZUWv19+s3j3ntO/XpRUW6z70BGhDO/l5Hw9adqtR1UGEMlVoEePpBej
0YSH9woFqaMtlcMwZswZqDSEu+KT21j52vCLd3Ux/alzvt9lHKWKwyqkYW5y
Z+rnPpldRBQ9YoDSYseqzwYRTQ1VHtOkr9uc+kZ9XAIUooa7E3+HGkdsG6D5
m4I/fs22CU6210FcrocrR+ij3MAJHItuIoUxkGLilnDh/aI7009SiwVKXixK
XNfmI5TLxs4HEpkWJ49sJoR/VI6CogpUJMBql4mWtTLpbmF14Ey9HF2ON0ZL
NvSw+5sw4TSWF3cQd3Eq0EtxM5erorF5smbTg1BnM9aFcA3kkNKtU2jU3j/K
jHgINzNergTJJBmlM//vw95w9iQ34MLNG8Vm221vgewOCokvlDKJx63pGWg+
zU3sANqDenlgDt8NB+dKX90e6B+dAqczUSR19L2udrsacW1iN1PZkjVg85IO
QkNz7wHbrSwmLbGx3R+li5JuORVHJhHkRZBQdo/xlBdBOBVgW4mSPeLYEC7L
WI2YWWBQsLd6hvhtBXFsKdlhetYgQRdRVvOEIhXtQWuL0jzPt/Nbr+DLV7Ah
/1V5yhEkkpUzE59rZ57JUV6y8uvyzEqXNxKGj+ihLa6VB77EmitCuMTWHJ99
gut49lLaT8gewEOTpS/oJpxpg+WlwSLpugJqS6MpDG9umzQ956Mp+j7ycU/+
aBr4UPbOdMcITolNaRxNI+FkMQ1PUDlA7g+aeR+BtG/dUtNQfTLtEU+sh/dw
kBKv1Llzlqfjp+byEx4YdZiQzg0nxdR8wRt4+x3kAzzWoB5gai+kGXgexACz
eKlilSqgwjDa90kP5o6+9+HwbrJLd3Giu3KsrjucbNVcE8xz1xESXwsK6RwM
i+YrqIExpwDboE28XjHSXLGJR1wi2v+SUVjBZyxKDnKKyBq2bqBcyOADmpKx
tq9dFY+f+Yr/3/tsaseWSqw0WmoSXQhC10MBT5tjf9lfAEzvVNJ6w9ncCVjD
dIHpBiTFr2KCe0JI9slYmJpM29zZw5wbnh8E7MUN57fRlllgs2og8aOztRf0
hKlrFd30skm6MoJJsOLPbFOTwL8ePv0AMGEgSSq5fN/eVcqvwB+DeXXc/4q6
yEdFd0yke5TIqcyWCRjucnpI8UQuhw0ALc/81vX7kvQ3oqyG1sfHYSB1RGoN
F4ABKzyi8J34oPetRdnsYEVFm+ah4G2xa9vyqiMoQx0zcvMVsvQCINvcvKYX
ohwshbME1l4/sEWeozXRRLMxlXW7T7PiwJIF1jSEiRqxGwgMVa0pBJ50gXiM
rX3Fz8m920JyYWGA3/IkzwDL13G6GF4ab8NayvxsuDqjb+eqQTXSZQ+cbMUH
VYmNZjqvQDlET583mVVkOx5oWIH42XhqpFjBtFKMu5/jK0uoMWwVQNvTv7p9
qym0b95zLQEiMitRXiOlXt2OPZWwc8xulSFh5xiDRLF8lfp7lZ71hyZbc4sK
qU4d9N5xaDefNXEbiWz8sjcoHXcAHXF0gd/+BRNaze03k6iCl/nxMGTVP/c3
dhZ4KyHaznIj0EYzfhRz88tfmB+5GqeW8gAF2dwtOQhjcB4wVYfsgE/R7psu
mhvK12RAJs44LdZ2jq4iHli4hPcsRBtYMzHQXOh3+4Op3oVO6M29PU6VHDSg
yl0lU1uUJ2B2NrGOAy/GYjjR6Up6K0wM5YehNapIx0qsAmgYKItuPUtu700l
nmFOS/0CUxJnaawbk/lBkhNZsgq43BL0UJ8oS7xs3Rd3UYyr7YpBhdxurKbY
BFv/60B5xR/Kzl4BakhFisfd0GddHpMXzBzljefWtyjVdGDIJk58E3C7YUhN
zeJweXtWqHFhc5BMzJEeV6/+ZB4HIPyEa0MPzss+u9NXu0CEdvCIue99pgyB
EUKzAbF/uwcce8NwgBLUMle5g96Tl9cESPJMx7kY1dEmsAeuFDL7HHziR+xB
IFxksFVZJ4kMLFRKjTYQTuSO3/ZBpUPhcxBeD3OdfAzPA3MEGiuuz4bOBoiA
nFgz4aa9lQAXrmpfJH1FnFQx0xjrQ45GetTyiFL88E4a64sZP5/DSdcbdduf
RWbpqILUDwoJSwns7QznqhhzcKC8/Aq1PqCziyo+Bpntt5msfxsxkiJGC4+n
cpNk7jws79BXetgaTONl6maAOWpnDqAyXclMLxrgtjVvBUrXwUmm+LsCXonv
yCwXRT2izymeyS92uzl9eKUSYdUJRcW6ewGSleEyrx83Mu+AF8tx94kDlI54
4ZuACWl0RxPQRAlKeiSmM5+EtClON/aVOpNiRA12Bzer5m9QgfWxFTPBMAP6
YnAdCJpc/TH22cjVx8F5P+mesiaXp/mFqBI6bzvmJ6ARTtMPsmOXn/RiPTKq
NOoMyncDth39QEPCaPcodwCRsEsEEnPMIp0fwwDHJZNClu2ur41MwXH/uhmc
CbizQ3G82q/1P+TxacUgSH++rbjQL6lNqG6OCz6mZU7cThYdNdYKEB8G4xGd
1FpdgYR9X04rJqd7LFCJ+i1V+MFWbPGREyIoZOAYSWcz+OmWUeThOY0x7+C0
yxYa0ViZPhhYlinrJv/O/DMgN1IXaNL1XRfyPYsIVvkXfHdhV+KBYD7hUzEV
f3Gb9rmimNtgZZ/ETQg/w1gvrn/pw4DZH0axVfGGqoh/ZWAHScRgBf1ktF9E
0lQ1PBNLiwrqhBuz5Zr4PkG9bVrcwRBgYjDYNNN8Al8askMYmJsyF7zTZl6U
AkLt1CA7ocxGBcPat8vsYlV41ztI0ge72WCWNBJ6qtSuBAfpnpGHwuwTBA/5
rBbpB5f6aP8fzgJvBdA10sLKxbnS7QtqMJYnTdNjHKmR88sLFMXNPr3y/hq2
LRDeHdrPjxyBO+mKj1ziguT2oQSY8JZINrDFxHedYntLguvLDgRqGLvDjyV1
bDbSZ24AnR/FIGEmv1P79Cn4uSK85gtvcWlA+PgWHdWaVwdebHyF+rLg/yjK
fALmtsOBVCpZs05FJ9eDEC148HuIwrG62aWr37Ky/D4dsELOQQ/CkPxTrl+X
u2UnxuXEHatilqACAW8fMB6FVoFOthpT4+HmKCmVDkgPIzf4ZDft6/AQ3tZO
dDuTdIkvUks4aaod+zcvZRgXNMAnK7CliWEylkkRY0R7nRQs+o3BdojB1Uzg
D5EF2apfBU5YA2f0Dm8r81e6oyonSqLVCDl+5cnlaffVvTlRFVziP5Wi2qEd
PbUnzKvzun0jp6pAMiGlFQW4EF6P2iWT2fSQlrE7n1O2h4S19+BsnAUwPFLR
//N9lIANPzj+uq0wn+oN6Tl50A01DWrKO2kfbQybSadDH67GK15Z7PsJwOj6
YFwOF8UV5PBjtwSKq6tu9PACFaX6YQQlO4WI4DECCw4QCUidK9OlV2JkjzZG
G1ySMty5ZborpGs5cCX4B3OJVQ49QH/BiobjicbGm+9zYC/af0R/Z9aOiHfm
+c3NW9nP0MYJY1YFB4+NvN5JiBdRXf88siA5BR2HR3DzdAHRMGA90v3am+9k
/z1eiomdFUc+bii4g+E+3BQFpIxOFmC+6tn77yT12APjbzaWuWrsCJyIoxUX
WvpIwiJrmlQXJ7nn4stc5jrwksNkV/DPSOQ716QNx3BZ2JmJxizkp5+jQ+06
vTVz744JQDjuox4OAgOinhdj+MyginPfwYszVveqKf/ypkcFnB6Mv22f3+GD
QyxPTbTzehVzvMuLTs8lD4d83l0bZSUGLXYFXo2icMHj3JmvIodxBM2gHnId
IQVSFCShmJ/cd3i84fsSkdZTTl+7jI409JrU9tnnZYjdX8oxhfQkxBS57Z7b
/rJFgAaaj6yzG7/VrvTfkevcVCAu1s9OTwnGfkSQ4bGxarINWDVEve2x2BBQ
hE/2ep+Z7xJXlU4b3tMbYfDVAA3+fioD0B8+Jdo56sn0pJD/yirA+fCJ0HPi
fCVpLTgOg1OLjVFhpqDFD9iRMFtgxH53PplFfMYJMGtws7Iz0qUYNgIEsq77
fkZXlBScqb7Ga1cZCXgEZkaAWe4V8o5TVXRWtzSlwSd6knlSIQe8vCyRcvcs
jM2uuIoukv5llrpQwyTab+XIDV/jCnpwCXE4S/6dnt/b8m3K6qyOQG3ZvbGu
ZiRK6XMmzyZplxCrO/Mc7r5slwBflX6lnQSrvb009nYk70VydeMmaTaKuPTG
L1tvBSAEYy50Q8IJOzIvQJteRGVyzoU5LON+HOczpZaGcPUeViufQDr4tbWS
3yVhUv3m6GBGguafYLQN5gud5wwj8WtoIxnZk2dPLTRlJzM3WjXlHVvRNu4+
aX/q2fUwMPjicOf5YIiWHq+mXkB+q4WcGkYVPCSQfOdJZH69YP8g0xAPPAtS
86BqgTtwWSqvXtPAE7TmtkQ4HcrzKM0xpZLpZ26YjbEoTYkg13diLnK+zvWX
N6mkeAk3rxzyGjqHIYovNFvptAUxrekmQgniUUFO37imnT7uy/n6fKrzWZ25
G8E7rpVRHPXSUDe2BPLMeTTfs0zPeHssKr7rqwEk65zo8zg8p1YEin6+AHfM
OVc5F7MZDCqakjusQVeKTP4WeBfbgAHYNIv/Uw0vHF4kmJ6GYmDD9+dzISw6
+Bi+ljuwm1ZLS1mcS5d9c7h1pSqAZSrQGNsNoF2K9fWSRD+WaxBSBSzIKrUR
JfLPkpAQlbsrh3rC4EueWeJkn1hf3K9czxV/1kMb981lTgRtLJwTRIn8zcxZ
eGi4upcNVdAVpVlrFxBRXI3Agn21p6kf2Hqaq5CR4DY5mWlZhZ6EnnBZLMXb
kiJ7s3LbbOkk4XXR+SsRsIJQePkrEmmXGVD8n4Yx0nT2SMFHzhtqQXJHuoic
peJMJSl2GlfaG/VeujvOweQoGKCctf7ZFt27s+stPvYHD9a4bN4qadj/Qna3
0Msgg2vPcpbKwOS4ynOfjlkm9nXEx1LA6D2vBHVPGac8FB+EUSGT22oNHS8g
TiPhf7pkuPnEvREfMeIMdxpy1yCRX21aK0qp1MUXNkWgL22AjIthZbd30y37
n97imIog7OMxFALJHUBvcUWo85sOEaeZSHrcFKOwW38E6+GDqlB6k1xtxTMH
7R2+pqVzfOaQpr+OAoFBLa+PlYQABDKVdR4slx0fGj649dlKg7PBRCGWBA7B
oW25oq+ZEpJ5ir1G9Wc69Q/38eNrtfjIcxl26RfpAI7gqPAtWwRBvyzsUc6S
aix0bXKd3QPd9sVxMEkZ5wScWW5GX0mkroipGSw0pp+C0dJ4acx9TY7m0Qjp
sNvjQgyXIEzJ0QkYiM0gQdx+4nALWkEV/uAH8DUJ51pL7pcmITOlWXpKyibP
gdkJWiIO4Si+yPF22XV52+2n/bYXzzJIaz3GrCYmfACWG6JiWXGoIBkJXEMa
lGOObdJJHRX9I5skPo7OqEbcQgjAuFgECZvK4u9igNHpzt/RaZxaD4Rpf0A7
QHuSud6IIIwCgiaNk3/j3den73eu9PHsOxXZhK9zRN5C0M4mMnM9wN59wK04
TWdXB+pq5X2ZPdBjiIEI6FfPmo+kYTY3dfwL7cucg5yQuoQZrwXRdeH9Es4T
tLdK2ye34wpFOfs2LD16GQATqNODJ0ZYi+Zl1ZvesQDOUxVzVgReGxQhWbbJ
v+4whOlBzjOTxkNLsjnl4wqBEbft/qWzMPvBAx0ie+eA1d0ICcCsChFGeOnP
Weox06/JSqW7pM4TPMMNP5OB0RYYYuzFSZWhQh85w46d+MtIPNX4M7qZl/IT
mOG/FjNJzPDu8KzuukqJ+j1Q/XpfDkd9tjcLWQ3oK42JK1hwBd5d6KVso7H7
XELaKMShRfNQfATvlxhEBVdRNSrlCuW7KQxq18a/5e7sCUoPxsOC5e7ODceO
DbzgJCwsuFfuAkfMf49frjLlfKVhwcdW3x1JXLiR4FZt2hE0ebElF3QPEtBv
5QZJ+xm6dUrueCbReyzsgjiyf3R2cnu3QCv7/cNbJUeGyTHEwVr+qfZ9xI7U
TypLQwsgMArY2k0WZpj85waZFUTQd8ZwvUA1z4M+mJWYgIQrqcefwuu3VUyy
BZzJBLW9RNVtl+Y2JCwG+DIGNAGbhqM5uBXhFBnfi46SGueb2B7tHI2SybBs
EN3y9dYLw7irTjtcRCmpKQ49H+4atttwfPJZG1v9FnzilVSjdonNo/N8VOUD
rnvp8CGKrdLI093MJMkXSqbubQFscAf75WnP+Qo2m0kVGzQIUrIzFzA80LMc
MFADAxfc2kt9dIY8ZWTdD055/00icc+voflxsAzzylYCfb3KRaFUYo5BOAGB
IYZptuhxhsGHYIxSctFi9vyEyMPyLBVUsZPIpY/QJkOMNU1Ju1MPJ0L0TArx
Wyox4qV6m0z13WAfd8tcKkkP9YBMM6lJAYhgkpyBVRVtfzo2KlVftIg0ByOu
8Wuyf9LgqMlQuqOWLgT02cKOn5RpX4rdYfzfnfxxLXkgwfnvYQmoDWuhwUfb
65r3V5vxEn05BI82/pjXIv6OinFp7aXSe5zUr4AD0lQwOVRhAMZFYQmgPcVg
IcP96UpehWX+lbC7iXhNID13QScAtygAFwqInhg418cCiXw7F7DVsfva+Txg
Rb24UpYjXXE4NY8cTSfEYtXasjRKG2xnhyIE84QrbLEEiXFMJIxGI75oCpbu
2iZi6ukPuTz3itTmsaQXDoOc8KpP4gjkAJJzNrQPenKnifpxvz0q8F0iT0ht
oyEMtn4Onhm+A0Dj27PXMROZz8JoIYytUOKLujHvENz0ZTxYQEWYjdkz4jlz
d/jZ/zc0lW6jkf4ZPEfA+Dt9kL0LUzcq8g9wlOfENUUcQVQhadIxMYIgbxWu
n8AaYVa/zm6kIjylvHcvY52oEhw8jc6tnbnSg/NCuDVkORWlwLXTd+WCucEB
cpFGtMVubXUTWVLq7ib8cVYjR9oe16XhgC3GbX5wZU6WpC2/mt58Jvg3fxOa
/eZ53L7wt3wAeFbzlYXw/HNzPKH131drVVQT9RPiB1ui/xa4WMUpG+wHsCoz
B4PU1TXeLk52wnOGoJHCLkXmXbSbhCvraDwWEGIcHxseyuoRzWdMOuBWz1rY
YN/pRDeBV6lNmTVEck1C/BLe8wUzoZHSM4jHu9gViffJ8OAyywC/oDqD8uUa
0F2SuNL0dtV3+iweecibicda0z7FHKToeZHqehfcU2oHtxQ+3sadKYk83nh3
1J088JK+4eBtXSNeEufghePsWGDxgnPMjK8fylkq4oZzhVIpZbBjNBc363WY
Arof9oLtJ7bGVFpWmnmJvAsalXY8QiulaL1WEdjXw+jJUwkCGLN0FwBieqwQ
t4tRulWc9DCEa+NcbKgKoSuSMkiRObYB67zu6tB89gKZp75VqirKYUIEFbCW
sYeHDW/D8Imaj2UWIavAvYzMo7bwjPGvHomXa5WD7M5hXaLnuHBEApr9RzI1
2CfCMzpZvzagF9ieJ0agYjhUM72cgVS/rOAZi5lcO6cR5O97qpS0qfOLfXUa
NRyg9CPnRog9N14F9Q3f2TE+jt2Fz0YmoDQ40g2kM2iyPmqzGYuWwTSaOwJD
OraPfOOQU2Kb7x2R5sqD4KdU4rQhLyZ4CXyXLh2/PaDFqXHNu0+jaTa6tUcD
iBP2uQ8L+2S16+iU6hLLlI/f/DNGXpktNT8ZFzJvGiBRnkIxdWScKTYsrlDg
NJCgYP56xVWJbhs3SfmjTMl1cc6wOzeuPfiXwODvVnTo4u0t2ie7UhHildbI
bNitceBc5hurtHdeKdwVYTMxwbJZHKnZ/ZX3cBq0SNbkPRp89Cfhzq0hC7J+
puGEHnqHPPtLW1UCR1FOMO038nx5bba/9hTDsmgEaTuQYGlftDNrTnG3rpiA
7arHewaLUJr5E0704gBjb31ubv8yjalFKnLOHiJrqN1ARFUTohUW5GKKu4Y5
XJr3U0XwiCw6+TaqK05W4STZTMGoQBFAG9sqxZeomYi22OYTz5TLuzIdNsrj
jnSzDnWE5qbxAzDvTtblmsNz9uFsQl/0d57NeyWPNf7hvwWuaw48zCXiogqA
nWQPG8BGf1iGvG0TY3wOxOgMxrPSZhMLfLvvu1zvcCasm7A2qFVoExh5eH9U
43qRzmprgmNTfiaJsfeSEK5jUcp7OQix2uHUZN9qMuOYcZWnGG5vQFWhZmjF
zuU5s4tTTJqJFO8UEk2M/8fW/9wrWJqvocNV7cYVneVQebwAOE3w7BUWkc3M
skeMBCEUjGZsnRIGqQNHqwYg1xCEOPt+E9U2CMRB9p98Rn3Vzo9IcL6ZRbXZ
3FBmxbrjmYFCMnfYyEjKtcXTYH8Y+jNyGTBqKzWtgyqmiE+5iTFO+73CuC4E
6j68O1dShBOtKZrAzmUC/COoL/tkvyR+PFicY3adjzXSpnMN+KmbPj0wpzaV
8SJBJL4xuIaHtkytqJRgEFmyq7ioxdBztz0C5LognI4uq1Jx4X9WRK2c8rIX
iLKGyPS1x2lL6PIsCABaWHW01CQwnMBB5JWZoSwdZ/TrulSC65+NweukPatS
TZ2F9eYSyPFB5N5xhj6ZSVQl+QowIZWK/5OWP409oRxyC8Eq/iJ3nooTn5xq
p9DMx1agDOb16zhd7cVb/nBFVPk3i6fsWPv7/b3A0joEguoYJPCT/Bd6w8Bf
pAdxenabYzTXY0CFfXxRmxVZdn8QcKBB2LK2kdGOOL858MB7qNKDClKfvaIi
Wmlv0f9bUg4YH7LDJWH9Hz421yiZxoQGRU5YyxG+bQMD7wzOgTxTloRglX1i
u+wNGn0QffjR0Dxt7yl2JHYhAnZXCj4vF/XmXOmnQzJmBuCp7QuskewKOc8F
fFNisQrdJ45O3XymixR06Vo79kUzQpv/fU84c9w7LNP/FluZVdotn9x925gV
0/XerLwnAg6PPtLeHbIoNIzn1UHsgCiQwumC1LwsIoDP+leXkqtvnRs/xFoL
Abbf6lrSUt7BPQoLAjZVps9tROcUJdFnNS42izh0h8m8k6YF9IcgotyhFCM1
HnY0B+otk6ef02IrTiBN0ic9Kh6lMnatc48NYRjsz2GRTOllbIGzVAx98vac
NT1uazxFy46yGdRC2Ek7ZJZwKc4M2uNtiTjvPVU0PwMzTRbgiYo3UJS7S51V
HMEfrbQlSRbSfZbTYiOLU/1oIfbTKNCunJyWxpecvyml6RVXMhbOP3vxoaq4
VuP5CuVRen3nauvg0GzRh3OyQobewiYNV7GAV9Keb1Sf2xWYNvLS7dUSteVu
adcY6o62Hp2+5x4bdc1h4HLDzruWFwSlsmmx2XDft9wnWymXpsjpK65fqJmm
glbOlySu1NbnUBNuKSKypShsQX0HmN5hS8gUh9m8pgEhMhL/3AuxG6oqsjvD
d0lUrQTsNL65bsi787lLipZmh6r2r15uqsN5+jdPHS0YyNqvj1e7gbncTOFI
vZ0QH/zr3sewnFSniGb5imI3WLH+UH3knwt3jq/UKW/a0gyaKnmwHSPLhwP7
2LtnxzFvUURg0lQs9TxoDSbWPv8jKuNoM+9W6SPf4NFEMZNHepHaKVYW6h9b
W05uLJVSLTVUrrUgj+zrwZQTx4digGJFyidN2UBUdiTMNdVMtGmaj+FW9rIn
NGbs8HxC9Plsl+9KmatVT9fx7TAoIq8cWHNSAgSnHyMNBSpkXgERZLhFKhGH
mZxL9ooZKGU8NbTF8veRCrRgguj1ty9qcDor/0EPwAFccd1bWGjO67/DbbEb
2XNhwTtHpaS2iIUii7xpAn96u22k95uo3+DsHYyl8MRYQ66A873Y3luw5K9w
wpJtEih8Jzi1+JYnsesVn2EkLlDwM8mYZJWe3ZbGHmu2E2EIU5nfjgp9iDYy
ysqDnMHYj1K6SFPq1zR2mpqAW87VVdK63ic08iXk7a7PEgz20hVnLTz8V1Iz
zGMQ8yLBBj8pSCLMX3f2VAnsT6dVkVEG9ApBlyzQFr/U3y9f+cuNFhSTjENU
pj+TkZNo2Ft5zPnwxRIcKQvnZsScNSCyIHqcq0z2+mtsBy/sjvPbm9pIw0Qz
EjXeYbnFivUr/TZDRGCW89nnZ1ghG3/Hip0nc8BjON7jeAHCIhvY0jcRDT+b
RxZVZgJhsxrQZRa275+gaBLshlKs4qeDhwctpoz7aTEpwEsm/RK0v7e8ZfWP
1bpHfmPUirtezzOR6HgHce8eMRpABfsSxoaOTLlSJ3QxZ4Nw6NEhqvdgDVax
394FVDazHW4TgG337QSDlI34kzkj/uVspHYqbxcKHElLDX6EteCmffcZORUV
Qc4Z2OcKtqno+8DaWdLE5vrIfqwEtW8W2tL13b7S6zMiegLrVNLthDOPYM0I
+jYRYanYHnO9+TnypKFjUmK3CQC+SxUXRNQvuqN7GoQcWxU7IDiKbNX9eAYZ
e1od4+T0nfytqj8prvwKBps94T/g8OY0DIOCivOyrX5wR8evyAJU892jytBX
cV8DB5aRygQSG99be/K/jdALMpcXwqhwNwU4+Tx/X8+XAASkek3yEf5kmLer
6USfNOe7IIGyALj/YAAUS52VjX2T99wXVoQ2PGA1DiDPl15FJ8dFHpYRICwY
H5bzB8Jq3wvJw1Vpizm2D8gZJ9XqBPM6u0FqnjXeYnvrL86spFBqQgPp5qxu
cEDkJ58rWqzs/6v3h6r69oRH2i6qdjjQmwYGJjMjzaRHadT3YfVKlKQTHG6g
OOt/NEyi3WRMwd5j4iyHi/EgQs23MY3G4FJ6jcAJVJ8h02UIc9PMPoFr2+i2
2FLttwrGOl85bxvb3SJVAfhrKDtgqgIe4js9CsShc4RVARGlcBKksO4clUDN
NqagBgxf9GlyHB59tWvNM+lzeB/unmE4gQX2SbX7Dl5Banl8y3CR+wfhObOA
jD0xT+y5VSqXOPu0yA05u/W78QbGREr5IPUlBYd/uvosYDcgOVAX2cCtxcGT
4Zp2Sk91VfO6GL7zQ9PfkDbgjVUPYI9iFOgF70lwovpMXuF4HZx8uWKCydyY
jA8+FqF7ZycUNXLvlGucMV+X7RNH4SKa9kovpEH8p1OBtOEElCbDLjPyYglu
qxXN7aun2F+SiJ0EANfG07jBM6ByuAeED4ACz/1Vw4OiAQCvZeXAkiF2T8Zh
FaFeaSRukB2tpALVrv+Hx2NbhSXyqVtv+mXJ3ThhkioYpMtaarg3Jm/s+B8S
Qj/7wAcgUGEhG8k8SPL7duvPwNhiDmgr+9eU3orsTV9bf3GQ0gT1+zOfvgqi
d8ptirG5MsUe4f/Ezx8fElh8CfaF9W1skBxj8vtdtb1Hk7B6iHo7FCTiVo3F
3s9EZCwv9HpLdn/GRLcztwZ9ulX73nk95VFhFjNW+9P5olNoWeo6CpCAQgVg
aUe0RKrg41K7XrW7z8jr5OBLhaqJtg4NtASPgOPqXC8SHuBVDWgFBTVqjYK7
dJ1b8JvGD0FjoBqMGS5vGkMmzMw0fP78q7zu1JHcq7Y8nAdSvnXstISnogsr
Gy6Ienkr40bTiw/TF9kAA1QllrU5sP36FaT7JPDyd7nQlk1T7lk1FpSW7Xt6
ilIRH0IXhOld7oDHTy1kJfDs+23XmLoBsmhT0HQ9FZeLSxoF0MGRrQZCqh9X
M9yVcwa5kqldGvtnz1q8m4IEsTalwE1KZwl6DNTfNOTaHLNT+HH7FkYglLwV
UsTxD0rPzCO5RMSuoy168lBascFlUYA0TEYj5omDzHeOD/ldGqDz/GSRbL69
FQhC29FzCnAwTividaONa3QrtBUDsyfXoPiIHU8xpQeqzmKlHBNk2QemKEqG
raxeuCc5YZz1P/RnTeJMM5Ie2GyORDiTVJRbo6381AUxESWVyk+vvUnDW8PG
InbMMeuODC3K/qIzve0RvlcZ/Pb41KhHKzRnNwbP2RLlBcNAwjEpaSGYetiY
aWNKFA5Vjd3pPtkEfuT4jz+HruUqx4HbAvINaL91h+1WqjqQo62A5QMFmS1W
bhWa29SqOla/b+sq8f8Lrc1XO3XGZDIbwl8oerfh5NmFjBJoJxEOdiYpSEdH
jJ6oxi4pr6CAO9qEQvLPltAqvx29bBEgVQttsMNEv7a3+CnCRMGVibIphhFO
UqB8nE6LXdRUk0Fm/KauTVTXeXdffCMLkPpgWlMpf/qHIYuVrgE6Uke7uQAd
MGwMA2fJEkezs9HmeGVUgrK09qc8/boFAJQKgFdrMc4Nda6mWJUX2PBXmVz+
CgZGfULUKGL8uly9PNWPxueqGfYvR06v67sR6nhNIHqkheR8RdTvf5yxQr25
GnVkPqSdRwx3XjTOoiTBIusETknbn8KgjTWwcMEiQ5sgrbyptX87ul/sTLyy
BIFl7pcAXNUs+a8846qxQ79YRc6SCBIQurvrtZ4Q/IsbP0+oXvkF6n9GNAty
9aWB9UG+bDwB+loaI/O5m4eBSh91an+tbyDIwb+v+YH8oXCOP39ETYNpNWFS
j5AJnw3QZfHhRe2Qg3Xp9WWgXOym5CYjaYa4zOtWbPV758WHnkl/CYASqeNZ
TBItLLKulNG3ZhgbX2Ic68Ix7W0otk4uzbKxtmPBw94srtFHlm7rRoEW7fbH
nDij+awttORGvqGVaSNRIxee6BtB883uG2n5V1Ows/HEJZ9Sgvt6BuTiKlrN
vU2obcpyt+SjuzgHi/z8iWJK6e39X7lduPQgKTpWGfGkZ2U3EFTAQovkQNqy
gP/b6dAfiuWmxS9bBNiD70dF1pp8umjeZSKm5CGkL9IJWL/9pP4OCKz72S4i
WU9bjgAmAedj4CEuKlPhbKjF8nWdpzwhW1/VAtYKWtMXEJ4iBas+KHn0E8s9
lp+NIU0TE9c8cHNR+k3cDrAUKdISFDiVIvL7IPg6uwBPHVW5xJoG11zZR7pM
6rCTOqZw4/OedOxkTWX9eJpr196lhrFcUeVniZYYYF7woHJCcx43sX5Fy983
4dT669KrZxtRuFVW23dBNEPHk9s8SjLVLRJjUcWMcpVSyzksdJX88yMVgE+r
9B+B1BCliH6YWggFPPHT8q0YDuIXujTjczqpo+NGdMp0IIdVS31Fgfaj9fTM
xD7SdDO3eNlLoDj2L6fcWAZUUZDGkPySnMcnnE1itais0rjsE1//rv6Om8f7
TIrhYE2pCYDdWRxxtQHOdp1ArekjyffFyJXujiG4MWSoRr6vYpDfKWbouiZx
PJFrW/JvZRg/TRY96bUVlhOWD7tjVSkz2OWwsdkxE5Ky0OAcZ5yqfYVSrAHr
qn88dcySQ3pBkTidMF33iTCuyaWzOZi2CzxaH16jxxuIxUHMNT3esw20eLL2
L0kKziCd7ZZtoiAxvEJvT+ehSvGTC0hBRvArWf/504oUE87oSWxD3I0Rsx6C
WRajMJf7seTcU3ETMJ4NRGohy1Pq4/aXAXqv1DV8cRI7J6eKT8LB4BEtNIm8
PjvtHIPui2p2sxWUWRtp9anE+q+pohd8rqNLF+3Qo9I+ql+u4CVkI/Pm4Ya7
AFABhUV5fOTzEdHAWBSBdDXHHVBlOWyFvNiODcg0M0gZCeQ0fLsYcPdzOX8f
FFekspmhts8kFpT/pbX0lvusW7KlaVTN8WN5t595HspAyliSPeMBvqfh3wx4
RsrGQf+kb9+JaYXlCU7nNCp7xY7hwLlMyVFj/OB1uAXlWwDxV+fSC6XFjpzE
aP1n/SY0b7IwV80pXay7oTVAIco157WDa7TWJDvSCKLaZzlmo8J3mpoKc7/3
QjJFNf4gIkQX7Wbpe56zED1HHPJvqAXGWQ/WyrCYd5sg/Ou0rrudlSDlTVip
XHKsxHV9msxNxpEcqkRRXtA8jrrifPTtRczEVPS/7fPTFyGhOf47UxmQAZqI
D4lxXnO2dce5HCmAW+Q8eVXtfbSf0OOJXshQe9nAOc1p49W4KEW1rUEbIsGs
6TcTo3AeGu7sYhqm4gGMytNqCmmyl0vXVjesEGP5+JDmoya99hEp2xRbWSuD
QWzx3vUOewS5Z/WFQqQdagKQJHbFsN8MmHcQDJsI1zmFpFPhugHKBIHhrI3+
IxQR9PCw4G8bFHzQ7qbnXX2ZA4jc/Np6ojRYDkal2FYdPhr3+qxu/c1LxP67
KCgl2XmNkZ5ABkvokoOk3sQ5x72K56AdlLaQ7qk8mIS1mWOCPy0YRaleL6zF
FQqN8inU7N1uaNXqwsuOckqn6SXSFT942jv4uvrYq3Jyn0JGL+RXwE5Gti5F
MMjsla4jIB3daGqzCMm35xUcoEhlHR0ba/S1FZj6PGuq5/d0unpPrf1HK6yc
xsQ+lGsrOq4yzDVPzXmT6l9oZb1aXKJLKBzalYLzPOSrlsKZt3gIud2jDFLN
FjFVcl1N6Y62UtsyfilFyUqBqWTFXmjbMzu2jzzwH2mcN9/jySULmThxHChR
8CVzCKmsVMYLaB0iI8iY6+g15azneMwQH/NM0pGpzJQ+ateQqDnVZX/jHi8u
L7+CFVbo5FH7DVuF90seHm367WOy0UIUxrOBlmnN+aIkIe24L93qQkZKXSfK
2AtsRJzEoztj5MFzHOCf1ff+QYZjY+XppzYaaY5f127AdQwI3sHK37S/U9xv
hu/8/+ZjdXy0aluW917Pf62EHHK2QY+Wky3rRnNnMO7/dhZCrbDnhCDBplri
453n5IOpIA/AxXZb91bbi4SCTU7h6syzbOqcmUzwMl9+xzA63ICDgB99uVp4
XjjSENBm59drl1xxYwUtqCftkwR5wLXE5kw/WGwn3JUl1IY06EdEdjYTnJ04
+YCPXcNWdEHdJCyPo92ZOjVnxvLB5BvVs9En8kkRHTm8sB4aop+t+7l8a2EA
6y7ylA9B2Knej2x6PCPw5xHIvCaFAiSJwqTN+nbHiKnY25Nv6iOxQioC62Mt
lb+rrNnwq8cK/jGdFRwjMuZ+0sl/eHO9yaQs6zhXCN9Qj8u3SQDKoNBP/xoM
vobDwo/JnRYkfBh6A/oHxc17o9QOpAgK3ASVG/XB4WjIgH/FvbrFkoXRmrBW
hnv+golEaqVwahdNEbdatMCFdyrAXqdfDauiyaqcrSY5eyKQ2dbjT+m389u8
RwGKJ07/b50HX7EUoR2mIRP1ko1o6Xe1fE6QZpp6GgY8EAAniS1O7qYvYV9R
DmoF9PjMsCsj6NKN9vd2bOt4MNeRWDBE6qNlrnl7paa4Z1OBOyRZK6E8m24N
277QF8D9aquNjTqrv9w/3oKmzRcy6vgGxXby2c4xsdflOZyXEMD/Km6h0JxX
4/nPfFTL7mPRMAvdZNETLx7yvhF4qG7z7BSJYmElTxWnqiLoR9o+dsqcsowt
sE7LXbY6KjJCy1RVyUM33/qNzaHJbEs1aQYBqOg1MIWBAud6kfRPehNO6CvF
6uQ9QBH3HRHN7ZGbxy5S2mhp1bg9rR9U1A0kUTi9HlkPXogmLW7gcRCY3EKt
cAKU01pDaI3Ub0BABUcFQtvMLcOGgUPo31D3hjNa8XnBmznmww0PiNB4IhsK
ZSyYm/CY3U2JPrdbuZm3VjtomoVwqBohbDc3JAS3RF+JHkaZncoUirozps2o
lFe9ZRYqdRIojB9kRqxOxpriqc8rO+HFyaGGJxzZrBpabIzZH3FUwLsRvbN9
xw7KRz//c9Y+l+cpV2B+f4IbCKkMYdv3/HkZH5qFVO28NP/DK9AwBMewF+SM
qAQ6wroxlFtDtMnvJRKbBAad1lD9t03WfmRM/8Ddn12HHzrpxkrWyIL1in41
WGYI4m3Y2DsHad3UziJTz21ug0sckeM9fS9T0DL2P0Q1shM1dLurBTZH8OXY
0dNdazBzqVaQIvwbQFB/EG01IBNYIrAfEtDhCYb0yB5pNCGVCih9g/54jBJR
rIUC/v43sJCPYOA79wcdu6CSE8alXoUZGOkTqnYRgdrFZe5u/lARAT+vbu9U
ObCglOm3npIrC4j5X/vjIKAycsCVnByVpGQxCb8gTy0hRn78j6k0v1AQXRlR
uKX0znDCnCnx9OXSBhZg5//pGmIyaN/FNxMIuHNdd6mc1ft5yzpMtSX9/FAX
0l5A56mH/OwU6srp121suMmalcslvQPMcBAp9tJfYVUYbeJu+TUAggTp+IfF
jG0oQwwNwW8EdecqBxwLLC8BNDD7NAuvEZ9gKKJeMczbwGm1nG+gzZL43HRe
126FySmX1eEVTTVOIS0LkrnCb/gHpE3evUvfraHqIv/N0a9JuPdIAxIqnYQd
Rml/F6n8wCS1zHzR1r8RyoEtFyFQpSGu4cQ0VkCQt2E9rBYQwz5MQNMt/U6C
56g0ZFWARoq8jtX/lnvNDD8y957vmyaHwN+BWMKoNPvdG17tbLGl0m/Vjzrr
2nrsIuTK0pg6XAha2Pz1+r9/zUy7dFDO4izriTtdX+cpSlLWYS0xkjW4Rwwn
KCLpvV53CXMT4LFO2NYV6BP02+VqolVY5VMtHCAQcibW4uab4vBLGydPnL5N
hBxkwIkDFZRzRvYwf1fhjzQMra959uK9C1HGmUC5sr4TTyhgbAkwkvG4oAt2
pBlFbxHn7SZYZTGcKJUXShQ2vfZbR5yAyIutX4iISp1By1M6dTBs97lTqO3T
UhRAuLaHktBNNrvKa4apdjsmmjxxdglU8cSIxKc0A+a3fJTvRS+1dBKSQMQU
XBleoVSZjfRaIBZn/yZ5idgbFaUvvH204H/m6FUdYTfoUcRE9QZbPShT2tdd
Ac6G3cF3ZkgLjUmndHv1qu2guGWvScjI2Co22ooYEBHFffDy34qYhkddRuyl
2cE7Z2jNFuZ7pOJX9VeEzW0/t29h1Bo0V35bzG2z2r35m7MUr79g3kma43GA
t1Y0ngGnY6YxoMGLijiLPMBxr5mbT9S2IdlNWi1ZkyuxmZn4ZIRf+G6b6eHd
WAyv4GkP4GUr7Bv+PtokVfNU7wdWwDp64D3Q3o5PS0VNVujrskgyeG/08Hzl
qPtCd8pvdmk7UtU9kGU4y91oAedQ6i10wFSKPB5Ih0xWYB/fkoKQpiLsOhdM
YytTfTSW6+W0q9DwhyskKGWN+pHZKRTERcwYwHCOYDAoo3uBhl2rqYlwVpGh
Ulpergd9IRRoGssRINXOe5REGVTyb5k/qIMzWPTm4Co3+u9aJ+i3IkA2Gr5P
4IsD4/EM/qGZZBYvk1Ze1hc0PLURnaikXT+78VKWrcsW7SUfwywtPusvy7Yk
5IlKBubFp52b/V826Aag/wyIQlL3oH//WntgWEh8kDU+sWR1JZpdRakLz1Ye
uZ+PW/jbaUx2taIt/CMA5Zxzr7b2G0lUnzcCYQLVWmI/FSrf8pgztrTbWADt
6IQYVdnvwK/TDGkA2O/NK+47afpg7VRI/qJKUvkBi80Vm4+Mf++67g0lVc0f
YLOMc8hsaolX/b93MWXNzdMt8/R+uoMFmHbS2HRKBaxveMptoQQqfmdeW9NQ
4P6rOwB3wrS+fQNR498tITarE+hpBwJ0MNUonEQDyA6wZQoUZ1+Hf5LKTSGy
6OZqAuFdG3KReCJIG8GzZzpNp5DOydcg9nm4kyp/t+V6yfb2YJs91iMASW2v
qyBpfcejh2M0zZrIt9QcYWeyP/+Oxw9pyAnAuMO/UN8OguF86galxqfKHHiU
O5wELe8Dl+q87jkJ3r9n68LjprXAIrdXfeVCfTxlaZr+njbV1f44HoApI+XE
ycIgWvaT7XGr6rfZ0TYndF8e21aJoa78IXUpV0jyzYBG24AdrE8AxHl+so4Q
OdHtbp2Mehw4+AuOpySAIJI7p8Tjbv8TVpJIIPYKdN2UVStqjj9qEZG4Bl4k
Z5zQnwSMShIpefP8DPf78q5HGBHAvYo5m5MWrr9shm9WLeghj10R2wVt0NJh
0Aif5/3LN/ppYUCuaq9kL4weU7/um8DXWdreQyMSsqIhjIOkzzMEBiB6p8/e
t/aH/pQPS+wJV7qomtmaAQU71vkEMVpTUIjIGKuexMIfHhyAWdoE0igbrNfM
N46CNqDo7M5fGGOEFKeNO3OO4ns4iTG34VDvhP/dZfbidwymvSH8DgYaWqoZ
9v2BlYRoCDULlpk4bMt7Lxl8e1YDwQHWm3WPTNHOVykU04JBIrP8Nbgm0D0p
2kCFytn4p3VXsrWW3eiLvzbg/NR4or7Omd09S9IC6wnRClft0E4WmTfpom+n
TX+6t/9a3PZLoBnChOgxdjwVc50Q/gAM+axX7eRablBw1nBrF3Pzm9OkUgXC
ugXPBTsGnQimeTa06CHwSwQcAw7CUTDyOgIxS/VpAs3viinijl+S5ZdMJvl8
NMpwO5RVgUGdii5OPoPVRZC2ThrtEh5CP1MOyMZy7mFzQJoG9rw9pHvJeQZY
4f47huyPMOp118erUEFNgd5mPlzdRqDf70XDDu+TIlFQ67y6uzeGn/8FpBTE
yDbVJtH92/3b/2s9kCaR3HVEsK78gPZtQJXnCmv3b4YLGKzPvRvbtBFwaLd3
J1AI9fAyYtZOcCuOa/3j4RF3oZBJy4ZQa5enaR+Ip2qBVJwS6vs2GGn8BUhk
BHIavv+xqvj1UnYyU1DsEo/JGnZUXFEdtg/j4vFge3qBw6nKiE0bGmHkJz2J
8jszKTDmYXtDEyoEM2BiJ+9YWC7L3CrmK72Sf9YpOei4rqFqDjwGwlWPHAWZ
n1ywL3y1PA3k9QtqAepdGWbblhZf5j4U8L28gZr6c9hc8YOxj7fUSj6tVWqb
Db/WCAEIvjYo2bLiUrKHfBG1V8e52Vxwx1NOawLL/UxHWZAvQWEGnFtaEXmd
Iqqq/luLATF3r2jKfaKQoP5/i4Gnb2M5GqGnFJX1fOyFcOoFdxYEJum9SVFe
ZzkGtk1vrl1XMA6wlmhlv/kVI/DK2ho2W0XWIzIFmO4Y7Jx7japW/NC2T2mT
KeH5UOQM9WcXy5tMHkWjoyHTV6UoUY5djRuxREKPyr6Kj97jv5Auqjis8bLG
hKVcuMdL1ek8qmzmKVLPTod4SaFjTiY6bGEO/ke0rCfLotzXSY5nSvas7nGH
XQHfZM9cZuSyzm9DnG5S4/g3lU7L2CQ2raGxcO+7EHkcESkGzaR4Oe84fya7
YxMdG49TL/oV3g2wdA4QRPLKwWqG5+lzqpYIOwuStVqsxsvKLHEQsvH6R5is
fC6A6NJMXqDJzGu/5CtYHkxNjJtwJnHmgwLyIro5ADJG53oPaMpblgI7k5wr
9IQfO2ZHhjNtqIE6QliS3JlFTRdZq5tFaC7QzmhRlfOGq9MlMGj8zyXTpFGq
uJVIIJhDB2Me797Y7ZdVYohkqIgHWk565mwVsel1fDyyxXtkpdDDM53M7fDl
aYTGHuyWiernlQ2Fb5IEjMNBCE7bxk10BdPVWNtthLc9MdatBYV0ATh6fz/W
jJcDYUtRsdtqF4yB1JkYOmdPvYVBUcLw4IKV61WUXfOkLq2xdVicKgB0g5tF
lUR8dYEqKzLdVboaE9U5wlEquNvr8qV1AxQyKFfMqwhKAFKiMgrDWITfgjhw
yNT8vTHh14J2C1zEolYK/8z3Q4EL4AM9jzx02gvwuH2d9+HTxIA/h7E+Jn/S
D/6MpnyVulDGaSgooDGLUmwOmDXuY8adnJqOk2pgbYy8kK/tf5e1bpYu+xzV
1l47zNJiOZy+cFjqj8HfT8sA59yturaZXqPin51HpOMv0MuxhwZrY1x+r4k9
GRYfWs8yGSI+ZgyCIfyOogF0Li9Bt8fEX1XPgsVYzAR13lplRVKUBueGjjP3
ekIqiNPx+NG+w60jphX9wV2xpU44ZHEV4nBY04CPk5UwZ2PObwXjyVhlfxjl
ea24PWHGc6v7HKIgWKtr67nFHfimDjp0lkwvK/iV+fE5LVxxDQQPgAeqD6IU
EEi69H08bWr8evbfnTgBgehF+qh40Kp+eJQxzup6IPaTIRaxv/LNWICEY2pi
9rv7mn0kBAUraweCMusO3nPTBxe6FhNGt+uRRGnvoUNXJ3V7Mc7tGZDPdMxT
oprz6cQSCOWe/zsdSqQtcEaoR310sqyZ+JRaT7mLeLwKVJIzCC3EYBLKPJ4Y
RPFwwGVg234Jo5r35kxCdCFTgT9OnYiInIkn9EyUJf9zWLs5o/oCuaorpKE4
M/nkKmnCF38Wlzuy5J2RWlglIGsKPdPdU1MQ3chJpVHoNEOq+whbcXQROAW/
7zd/ptCzOcp65MBfqSbk1qZDa/8Jz7NeuvfdTT1vcjL3vvXOUF9eupbTiGTC
9VtWJN3jPTNGX6BH6pzLZZmwMYpqPpjlqeGKrNZCNq0cWNzLOb97KLG5buZh
nb+gvUmgRYutlaxqQqq0Z2LnZ0ntej8qWn78Ac/h1DWhbi9Ho6RM+0hNVOXo
IMtA0dmk9OgT7yXJ8Pwt4qhNvy6QvRPB9eml+IuLIgvXQpmO+Lm+YkP0b9iD
hD1+yQsqvUvqiMjFie1E4jY8EuQ27hTvMfkXQT/NkD96VZCIIa/V2aLgDOnQ
LiPyhb1PMkvo5q1Ay/SKURDMyDtkCOgtrD1agg6qoJcrvMki15HR++VFwE1/
G55bGS92KiXgmyZVKIwFu6599Vi53APOen1m2IZ9r5Pn40Va6nZ7O5n4bVK5
7YZC/efY23kw4CnzmF00EGRmxzOytqV9vEYAsdJEU5WzQrAOU/hCSCSlXQVH
q3m6fxx8CzXaYhGlft1gEEWbO+KTaWl8z1TJ/mkRBAX8NknknNo+9tn5nlqE
tix8pdANdNZfT1LctLOApb2NlUh7P+EmIeAPf2Y78DpvyvnKRFG46OahINvS
xmXfm6Mn/+STmekd462ZHDnEs2825Ops6G14i2CMzEFxFXEudISe+lsJ4Ce1
Wctds0rFbn9RkQRHfT4eGSzSXsSTtQtqxonIpirM0gFGgqF9hFqEbUVaqLHO
oOPesf6BlMkXOkZiTEKevfydYF59tQIH9zU+U+hCoPR6REYhb3N2ScoM2vRt
ZJI/Q36kQpuUux6Zz64TZdlkhJ/ftsjvcYR8/CLearGOpN/untc7k/p0WlH6
SMn2uEPiKzhRVSKvwdNCrBQwOcUREIgb65CKvJ5uxCL8V5o4NA0MbPrAUJ1L
c2rRyi4mQYweSfvo4te6zl+NlZIV5QK//OshrJ2CwK/ihG8kZAlwFyog6HCw
3ufGBzLB6c/9rr3a8ueCV0Z+UcmsPTUt8WOOOWLb2KerOHOamYLFmg045Pyj
0vA7pKtHRwVaIaMisbPMAwL5/r2aldXdLUNeOINflsWLvPd5eKCbKOM7xgFy
PIVJ1d8TT1H4NjL6M8NqFgvoPVgxOIL9WHB80L4/Lbsh46cJIuFvNcGtRQli
Dxm9JcmQ0mTVqxq2Gip3i2L9iMpcEVNVQOFZ6Dh4E66SQODgEDnZqyQ6EsL4
6si3RIv/qHyub/KJP9KABr1ksLJFiMgjNVi1Do3LuqXt1dOzEwytkj1Najar
RasURVfJ+gPacedPDvSU3RWQ8yAOSuOUxWHpjIBE2v81NoDtO/AYIxOkSVwa
3BuEviDox8N8i7BmR2v/88zXBteTIzGgBG7G/aqG5kXCjqWcBrORKeF+FC5F
ZvIBpDU/0lClrl8ARytdU8ZdfXMGT94j93kPrBbcm/ibki20fX8nrkP8hHwK
/Ag8EQ2Zrq8+0XIPuQKrxKLHDVqzIXtYiAmJytPPsyctvDhz4phaFUl3IsEp
5D7NZv82JJhDZG4nz2OPCIXIjXPt353FtWELaSKWoqvsqgQjrNZ7CSBQT2QH
ISiiPdZoOjmbnUOltxOiX/rCcfj0xaf4OgodusF3bB+cUAiLAtd1+oXBQyyh
wuvf4XqHbR1qeCReTou9fG2Eq78Z86J6MOkCTq0t2fAi/8CrltUSnWerEJKV
buKeAAhwdENFYeARt7lMb0mjSE/G0rFVx1NszPydbkJdqyXF4v75cJT/nldg
FaTgtFoS7CloVQFi1K40rYdmlS9AWTXPOgnNXpqmh39tiLt8wFxWQ+E77Uio
SHy/k732SxaB0/Du/Men5YPi5otnqNzNX777amWEuU5rdvzyOqr0M9ZpjR8h
5FM/Nb903NCwTH7/zEQh4ArG0sND2aDqAVoOpQuVfo7MzbgJJUd9BaAHCFJF
2btCxJzL+PFERP+UumUj7a9drXknDMXY7huYH86I2NxgtMnebUNpu9nKrJj9
D0z+Pkd9LTTNrramWCIEX1HMFPgOPmZuvi5jup5UO+8QvcRkTJIlyyMJTQ7g
CrbflkaKhpbqy+WMf7juwLsoH5nNzDMWdOfxPiqYJOIVjZf64x2WhVWYohbH
WdjElb/5XuZLP2Ic/4TFXAyApfCkfdk+Ov4laYgbHp1QWahWNivFMhUyLsJQ
uNPk1RVlq/QDSy5syE29o9JfQXolHsRUJKTB5L8Me0VLkG6VQUK9P5U38/yL
BhCgI87v6TwC3b6g7WoRtDJ5akhzieU4XcqFW1xbjgHenBnbBRv9h+zUP7m9
b1boxkMS5VnwHoH3EZgKOMgClrzaTcgx+cUlhgDJ5SjDaVW637dwrNUSUX3Y
LnZE1AqXdJdSSUL43i0lYQtOCwkfYg4rDikB/3slKarROmDFAeWoVUgmeM6y
h5xLSWlSBPHbqj/SrDDQe/urc5zpMG9mppJjdw8w9rcFq1kn+Zq46gXS/But
z0VBnXDDOzHWLZWB7VkhvuD7cLa2wL34WGHIzlMGL/qlhH9i1e9xhyr9fMzP
NF43TI+EH9l47ZislAIWFSsxH5X4GCcAmATi7Csye/Bl+ez8ghjtnyyv+7JJ
chV8ys4ftrs7ovegJmw3Cb3C2BeuPkHYKG0AbTASwMHg/0iohkxr96CGOUiB
fDdMRJsNYJL04R6cjcalU4jRQloWe8xntpZeqfbxjMzKdlGi+LhI3WLUm9Sk
wwhQm37btV1ZRro19zduEsCvLptYCAKfyNJ4LpwCFbkzOXdAB8uhWIcYLS0r
DQ3/lz29OV3JDHE8BeepRpTA9dWXnYNZZWGoYlbrxy6vMMZUWR2bIOeVihY8
JXJhaxS5gSTd6qxCYxxX78cFhleUR3QwBzd0iGdX5HELMEyGyhCRhSvhDdMc
0DnFBFf5ugbmZFZbevn2UH+cLXwsgIrGf8t7MgahOd4Pf24XqxKr2xG33kfF
F5SpppCvBjAs+L6CItYkPO4tqNVSNt5UmrG7RWH4eHdL4gyQcYbPK8Y+DVfm
P8oIsmCiJtdrfiZphw7XxxJf0UpiZq+K3E2TTNJMpftn/3L2hVRKJ5h3gPzx
OMolnRMX6NuTdbLBlIlZ5ypVlL/Fc/POjuwPH9aTAXJcSuLCJdxNqdzsp7U6
9Ptk7u8eGRKgXk+yaZgmDSbpAAulpKTJZnn6zVHboeKLi5f5T9VbnO4NTG/E
l5Y1mYB0ZSZPYrOlZ0a2b85H8CtxhIZjoO2h3RP89L7q6+Z6nVpqMzAfnsGJ
RZIOkUl68+tkO302tAmFwkGSa2MuXATUpWs+KqEe/2vlWMrh0e+gQj+KjjOh
kXpjbcoUadJUi8ZBrgf6u/C7PsBX06VP1RKyrjcUhDoBJHjJgvG0ydSrqEnE
4oTRPzkor3omaMWyreyq6j5jz0PYR44HtkyxPUwig9dCcsRwpt6dfltvE/yD
nwJeBjOvSu56p7QQ+fhuaoPU1XJMyHFoSLFegFr1lvvowKTWHGTVEbiCqbhM
lI/CXoyChlsL4Ht100p/xtpchrBMqxkA/tFNSOy0cwHbmBSiGy/1tEINh8BZ
9TTYqTrZwHNIsBm4o0W7goBcQaM5JjvcwQZpAnSGrORYTrPqEEqE33uIExHL
W+P6VMUiNPuRXlf2FZnWK8IR01XC4xcKOObILDS2cChCsHAsDGnf4ykSDjGQ
Aj7rJVDJyzH3mOzyqhL4ZhqM0dBZo0yL1Fn4e5Dma4JLtFtlh17xFkbBClEz
DszcHRuqxea5y/NAy6rOSDztdl3hLAqEyMfvX5DTuMzWc9JCJ+FBfd/t4Lik
2Vjuub0db7NWEijA8utLtEK8tyAd5J1qghuPdKi+Cergv35Abk0Y/XE7KD5o
0qcfPjgagM60y14pb22kFqrq5xASip7LlhseWzaCK5IiH/qvtxNYJY8NAuRb
jgmeh08fIINTTgsmBlt50U5iJIVJwT3X287cmQX3ts51VMX0CzcMknmLQ5sV
oYygE5SAqK/xRcYSiKh19cmrs5SgLazlalB4plXFJbWWdz4C/tqoKB20aGx/
XCyNIn92Q5PDBoVQfIItVahSSxsfkF9QcrOzmyIdXkeYz/0jZKKMHs98/YLE
jEIKY+OCBXi+iIxy+8wYwSOCDwI0EBhXDKSULfhMCtfz2+UH/BqnQoQnT3PY
ZQx43oAX4H1UqgzqODg0ciNmTslG9acmNVH7Uao41IHhEeBYYBZouKQUx5sG
ZvmncM0MqrHqMPeHT6fNQWt2WvDzjavkA79QNClmgS7uztNbklkYix75XkDN
8kIIZgH4Tr9WSZgQL9ucQbxhpIzlUXfqD+vgLzLMRo2Dx0M9usS5kI/uhhnU
0URkX+yHSkBo+UGdWJ5pwsNm4s2VTutAvLzxsNFK4jCH4mmu5q2i1w4urLUD
N/YsOMw+Ba/mglnEqevSBFhVzRWKSKdAoklwbxvPL3WYGFGXOumtyBvWJrG8
d6hXEJJbDOu28vSSN2bjC3r0GBZNFNk05rFQ268Plg70YNV5h2/tE/DGdxnL
TeyzS/q/K99A8Bic4f2kQsVyk3N83uTPw0A9dthZQWXHitbAzc1uirN+NbOe
wsMhVGoD8gycaoL2jOBx4q7GTRcAy3mz/7jmXaGMUP/ac+Kb6GMPkXlLnkTM
fQqAJ8yNcMfkmLPqbbs0BZOfxpE1LOsYp5Z3lqC77BRfPIgMd73otrFnonvl
mgeJyzKzmVp0dApLsqVadOxQo2oOSYpfmaJqYaZERBPCY8uGpdDwNECVGzba
/n6l9M14ot3gWEO8kDzXwgJ7zq0ERvXjhNB8xJPQcT36fmG9gFTHXjvEBaHr
TpRVr4inT9YDz/qzwkKfMX792MRykUNqcukAZJrO/5kkfQUJ00xAOAzDJR54
LBOCtFRfE++3M8sQjRuK2JSSrWk8ZqogXGsiMWc7e2duIYAMgJnUxROavfU6
+Y9TAoc6JyC3Apqx8bd7gTfHJC/i/UogDYHO0NQ3g6t3ZfgEz2A3lBgSTzqc
6yn+fq4CK3XlJKXMzj7DjJIRvisOp8nQJNP4yOaVEUq11XnqBchWskfsxSuP
Bve+OocmBQgu+40uBIfr7aN4XjGd/nFxEiLrtxl994qGLFOa/7wWV02qe1DB
vfGto4tk6sHsiX8at1vOrsuwQyPRY77OgFbz0HKobip9apXUspXNgzbYZqpF
F7rzijccyxDLXjEYSI24Wz1eZBdaWQW5vSEVkIvLbTZTDtyXbaFl02bdPV35
B4zK1xy9xQ4cDdWNWrDJII8aXYCl78WIZiVSY8nsIlHIa84Aqod3yN0n+GEM
CCatQLwbSjuxJ1YDzDd6XtzyehSnZwAqeFuBLsGwCnF1taDTPIj0u3xfR9BH
lSYyxlugyYwxdtByWesI+/HAExPEvKnoA4p6wkJCRukU3GUZ+8E3zJt8DiVk
kyirGwuSJ3tYAThIk5k9p2s6+L/KyFPvz8wsNUMpeqKO+7AQoLy3mwLh/LXD
mA5ci3OSIyd4sL6WPscUHLFKEzPnQkSCpxrPGPxvwZkPgYUQSLCvV6ODVjmS
zZWduzYZ1um3tyl109WD8N/T3mPV9l6mj5PEgQO+pp4zFLUtnL+J1fLYUO6H
AuiPRoLFQXVSken24+Sl2k0IX50CiBlOXIdjyVQ30hkQyCF3zTXa1vuXVtSE
c7CzLNilSZ5J1EV2Q4sWCrnlcanA3Z8124Lg0sjrgi6lYwZhjpGJF+nyij17
gXx03t7A+aOR+6kfTcVhn3BQs7kN7r1CvmfHtVgjsTQqhMuvRdHwqX+b/K8h
SozccHOhqYpX/05VwVfxmeKVtxM3wRpoAxRqab2M+l+vKpEw9TEUw5gs/EV8
dh/D3ZMbt6yuo1zbf37abHhqbeV+/Pw8eku/vfC4ziomtjxTs5Y7gyI096m+
3+v/ZbXmrXEhgzfSUn9kOVHsaPx6UQa3kJvMSldC6EAiwWxVExBTfTFd2uEW
P7QUk+sYT12Pg+PSbaHOZK71Tw52IgJMLb+iPO7J/Ns6H7b5prBes48IlZGG
vKXCa1XGdzye4v2n57VgY+PH/nfKZhEgxc5jQ8xHrs6/A2PXQVBMpOgoXgF2
Wbjp1OHhf1y93H4dQRwWb3b34mpXJXmmuGf3iKNDbfHGsKfLlkyJMm52sYKw
P6d4r4041kb+mB5PqoIT6q7GzptFdwG22tVxb+9V9lNevgn3vmcpm1thlMjz
tIUQh5oPb2d5nhuHCW9kK+hMx770STQxdIJCY84lAMb0CoRSHlPZy22jAWa1
jF8LwBCXPS/bBXAkJdE6DF29EvBbVcKiXcGLuhTs5pRIFuXO7s2G69+u5F1n
3aY+WWJ63kW8zljkKvlUGnCnySUNmAh7EO8PtSD+cGNElugvpUkQbNpwDFV6
edKdYd8UUUBPSqIYUdcNTGRgIApUGBfHEmD5FL+Ourve4yCAVpxp7Xm96Wqa
vHe5erLK2feJoou2o8m7m3DhVAmUDnkyITYCl6D+i7wzB0Ue07BWgBuh5yyL
Iq7KfiraBwUrTsJFkyf3iSVFGBinDpmZFvgDvzPBCNrTSHOJXptH5oocMdcr
QQPn9Gf5NN6HNWX8pt0F4dXd4cQ8fDPGl8xPZurLZb22QNiH5dz/Kh3PgVNu
AlluFzUR5WJrGzyqvzzzyRKC0adZzDRwx5YLNpw/GEYLRjItPNXM11pk3Rf+
0eRDXSgEPAV3HGL5DEF9fJbCeY7S4Cxl1Cpe1dVz3CKzrPq5BbMZ1dfLqi7P
ymNbxklSdpVuyY0YMeSYVsFvdM86q/Gsf8L9pbwKYaSPEzsuwj19Yg8be2t+
gnEKbHqh41xKyZhuKRVHMD+HueV+0yOUEmvM5dNFZWtdU1HAq19xla2B2Jw0
kB6wxggOZ9BoCSa0Y9Z/6akb5yvklhg6zNhZEBuzf5ZLnG/y9DaKJs+5GEFL
yBBs6Gytk5n8cNb3QVReMv2ShVxIb4N60GvohO7clHMph35cbA9uJlyPehEJ
+GWCvS5GDGupSYqShHmsIOFIQNl15f4KVmhgWZtc8CemVOoSUNtxDx89v+eq
xSyA1pVt4l0QvdE7tTshVX+6QHwBb09roblMJGnGPbx270MWxM6xTNIsdq8R
gcSG4PMEQafwfFlFe4JE50sIYCj/rsgp45VyYNFXfHJebs5D3kY2hvmLU/Es
qyZWA2yZMK15JluV3jxrztWDOmm0vqpP0TgTlwBFSQDfxsMq+lgiH/4CwVIQ
RRpSOhtKXzHc5M1DHmaL1N/NbgPi/gz6oU8vN6bq8om9gu2/tvLokJq7K3zD
xS0YvhPrM8ghyOarF/Mt7OxWerJdQT+kPr76kJ9qdq5f1V2OXUyoYpAlMtVP
MPEFN1Xxl0dPgTKIu1nxrRBsZK3Ga5y/2N0NUnWu4itAGQC3bFg/LlZ4BuS6
xbuzYtgXxTcuhP3jOsbSUrbjrtu1GotZ4SQRMWnaD9ZzuwiSVjDL8zbp6mGN
KFtP7ZSsbF1D+1hk7K0Y661W7Z6MZElhIDSDyhCoYnMaj9knmAFnJLLRBFCJ
9K2OImEPwuaG6lklVWuJyBD15n7eTISIadmpBQQUuegrS0KrJBbOAjS2wjgL
DmeSK/kFou00YyQFXfLxnqFHGIU4wVCUQOhWAvJg6icsmfe5gGXja+8Y4LnN
PlF9LoK+vcK+RAHMkRwe3kMP86/L529oCQUf6o8c9rod3Pb/4b7/OhuCe9KN
WFMP6ZLvPLKSH2u9ZTv08/kL1nSI343Plyl4ZlH+mNjuqMW81aj6L/wbdB25
M21mNY8iw8lIOs4jXvN2MENMykLc7q2NUQ9zTJjkTYgejePZV8UnBp6TTXuj
iaw3Cg9iCvl93lPpDCGk93ayViC8ZNTbQgwyRZUnuqOP2U/KPAeu+AMGpnw2
euEyLTzHOS2ns/gGVSww8FM3BNf+AD1PA9Nssml4z3+cq9adF5D7jF5mEoAN
prQgpbEhVraICbmxQMmF5hm8KovMpddxMDVtA1WERztaiRMHGqXI70ys16oj
rpGIJRCV+9nczv6mUWX7l3ol+H8k1XeAAncLSztK3rNj7HWTY4KSTvjSbvB/
GuX5KIdbmh42vbYgLtRtzOZBqV5u7GXw5TNCCt4lGeL9ij+AhDsi2sPxTQD3
hLCAvCA4WGqdY0ul6o0ib7aku1cVdR/n9J4UKs9lsb4Bllixb+5Ws+DMO1UF
lTR0B6hFR5sR2Stbaovb1qA/FFPf+JF42LLuzksUxvnfMqD+O7HJUJ0yjroa
LKl5j7aD9LDQ3EQkT9Bn+Qe+89MLcJe+m3tMxeiUwtWQqN8qvoimvlolikLU
Fo4w3C3S2TaYTi+6LtAoVfktKtmSl+NNoV4t6ZlA1utHJEX+a+pasF42IA/E
b1AUCV63RvbLicw1iiv0U1HLaKi1XCn+ZceYwA92pYzRfNNo4b+3a2FsXA18
ulmRaRAi5/YA4gq6y9AWpbMMAorha1ljH1rIAVqgfMJGXZVDv/xeyMNITS3H
yv0pp/OW9ATxcKj4Q2IE7oXo1SoXrJDIMawh73asSUPdc5BhWx85Bc4viaAI
YhVCAN4qif/hgq4BNJ3uWVO9Jk1ZuR/kd2qLcT0JQWj1Y5fMFIhvAL4/fe3w
y8kiheJZOlsIQJV+RI6nk50tkPXPpSmkFMyP59MJy2AGT7YVRT1wgLPhxRFZ
DD7I0jYhGF1p3fY8pwY25TzfDJb4aJk72mwLknfoOENDbdTahKB7i0LmpUVK
hzC885BUvNfRdc5Doioo2u5zlD0XKaA5RqLL6zucsD8nrkp3RHmQBj5RxwFq
aWu81NpZmulXn3gwT5lfHpmQai0FGCjT+xV8e4aHi1pY/nQIuf+gNgsI+JbG
SDHsMqhVTeTkf2+hBbr2Em4iTMnW/j6OBWUxWdfn7AIM6zUzgQL7fMr+gi6y
sWzmwVWM9X5IaPAfioZCUxN4kjez1EtUxoQ78o8WvpDyIk6mpAg9W5i+3/gI
Bb1hg1G1zolxRVa68lV1j+i/9Y0XtLRs/lDzWf+BxPkemitADFnmkkworSH/
atbE+YMUBXDnqTBLxOLM2Qz+SJFtlQC4aISbP2/JH9q+I97iXJt4ioFDuWZa
OKVjN8d6hcZJ1KdIn5zyh+wfNA6Jj4GksYfAB4+F1Cz2AS8aGLLJxtr+h23P
GPdqh2Rk8C7hEbetS/TSRUHmM/zux8CfOq323bClMbMpklzojPgMeBb/QcWW
qtDT5842rUKaW6rEEopoX7RWoUkgJk8zmEZuKXOEMONXPoUqlViST+J4uUEz
yFSnaLjPwc+yiKKERlCrp1WqwEeeqcUZ2veHYy8BRNE6oRfGNHqsZV5f7wx/
ogCSM5gDQtMxuisPxtU760yz06pbSmaJR15zl7kEEeeEUyLdFkTPP/q5feeL
auW5ca31DhHbbETJKdjbt2fMmOcSKTfKnR7sLr40AWtke8M1R0s9/bdfBKc/
pIKos5XBm/30Zc95f7KK/0DnyxiBZjt9t5NrFaCp+eHBT6e7A9ML+BXvUmub
hH+pwpEdPb7zX6RP49pusfSw5zW/q8Tn4AC27cGl0/nLRLXrOwFA6AhxYkXC
GYtBJoMG4MOH9mL7RYY6qLpvSBX4kvJ/D43a6aHmzHBUCu7Krsk0SifrllRe
wT8Tr6V045Zli7/Vgx7cjGp2r3weHFJstA2fX6vurHThkZr1hTNIWX+0GFdf
qAwJhMNKMe38ciKlJQIYsRcqJVe5pjbdC7dXom+NGmhdl06TRuCYPAuIW/tQ
XsvkXzzTx7W/5+TmX0aeQhAG9DnYkwTc0RURIJFudKAU9BITpYUzaNoDVxrB
sJIoegbG01TOJp2hYeeOBQKGKnNmqEjIUTn+D7jt0pBBeEJ/XAwjAx+5B5gR
9RwL47QomY+Zvw4ZYRUTXrN7svTTFBB5cjwCXN6ik/QY4WLDiGAW0UhnYgkD
0b0fn6JredpbTRglJiyXAEt24eZDAqbOBZ0Y/6Jbz5IhZChFzEs6whOh/wTu
1jVRDlW4qQttLOUtY2o7I+t4wLaQdiCRu7VsJUL9dy4lDPohxFOm13ZloOX/
p44jAdic01i8mlcCnK7V6G1xJ/1xqSXgWrVYzU9gihmt9IGzSgIkU4FfYMix
iobQXq1oIzacFY9zKFM3ebMAFIpxGcRpjAj3n9oBUsVwEi++9S0r/kAl4INP
g3n1r2vKU7TzWGDWNwN9qkxn37nsamepfkEQmwp2T1d/lqit8JDnk1SOz03m
o+kcfRSbW+Vt1P1qJ4UtutMGD58klGfS8CrqOU2oWUeOFH+FqSmJSpe4nWrL
2IFZkhdSY+W5Vvrqzx4fsWRNsBgTTlfG8R8ImbLD4TcSTM1JK/nbnVFJE5fb
28utENm3WEvh/KHeUYjhc4fpdrEI8stlbioOnNi9eeVO7Xi17699KMjWB6Kl
UL/JdDSZLdrCwVoeBPfVCVcmA/fmdRa31I6soZW6LO9zVPtdv4NkecNyS8QZ
cf/1eB26Dn9+4E+4xrB2QyGjPy6Zhj+ed2TWkvPm+VMecYga8TRuzZhV8elF
GAEo0JanAG4cztawzOb2UMIMQdOYglGAk+gSZO7MSjOeiP5eFbsBhL9O8KGV
pChipiZtil5MFlLtGux6qieJrDfJpd1NVZe4btmZ/NytwtaWtUJIIZonUcIE
ssuUbOG4F4cG8u7qL/7TtShDtNANKExQKRH890fEcuO0JZBGUJRl+eYODzfT
fUqfw6L6ssW8M/qIjPYK+nLtJfY9DEogu8eIcQaps+dwZ0sNQm9vexer+Zjk
POyZF+xT562vs/dk4Z0pVdtG7NVr7tzmZABZx+n7tRnELk42ulUIVL8DDc+R
Rd0PBa9uLzbJmuom9rHtZogq/WXyTJiCan66uuA3Hin3L0Ez09m4Xrsie7fi
Ykyn3t9xHrVBZHd2ngUGh1A8oZ+xIMuJ2ULEFLV+wu/zNn6VIfAKhtJUqUex
UDvnR1f/zueOHyPpfmcnqER8ZOwFUwXtswItRdVuCfIMwswcTPV6ANN/6Wf2
AZd9LBLsPzqI1tpAMieqoho9vBWaXiVdMD1gla5tXy3RWy6qLhDkUDfMAafw
c1QS5Ugf5HzJMSSSDYRPm9OO8O6ZeQ+1NbDpcBf8XX3qf/xe2rSdmT0HoAAz
20DzoY9hKMyTaqDTNB5FOhQjIMjrzKUslyp+jfhoxrcb1n/Nqehpt4W0bSXD
eEG2DbV/n484/LeLvnn0s1IFWrghp3fn86cnnrLHUkTAD18l44EnSk16yqdp
/APWcgvlCWoKeMrVnVjdlhctrBJRCQf9aOP6uEd4r1CgTD9uSiv6tJufnRsu
Dj4LT0PDN4UMwPi9xK2ZtvtLPVJhU0lwAcEEXis9LyjIaXMEe7S23HZ3eEnX
RRGVImiqXjbTjWBWimPbyaeyj1JI8FpCkRirm0sr1pVgxNG64T2vzhf0+97g
yiOicAR+sDDmsUQk+4HSDwqhNp+q1Ibm5wJyslMCaQvqfNh2clDN8dl3s+7c
6BVbVRB1mH/oGWZDeLAR230HkkPTsxVProsFPqQHNI+7PA5bdL5tyG7ky9m6
9hlKNDCEQ44CSbPpbB2U0TerPX898wIXH3zPNTaXris4n0M92xBhqrwQPyxv
VNwjapu5PlOj47LcQVkboKt3ZKyjugpIRRJ7EAA3opsLDnjw96rnDYx+pOnw
y3drQD/aXCq5gphbojGgcm78GYb24pzIqCdPVUpDW43wYA647mgcutqZKbj2
eZYoQcviRRxcpxwW8SHzmoSw/6WFbCyJLeepvlcg0c6+eFK+ftv+88dpqgbF
EVqvIR9oIbZN2BzvSH37oy44+5qgXFapZDJXChI078mSTzT01o/RzlTHjGE8
pBV9pNiIFQmt/bYGpxTZ3aL574XBX4+7kDfR/f0SmPylXPMSavWZm/A0mYNL
0935ueuF9Q1+fuEftTOx+j38EPFPCA+hjMuXCiZPA96uTG5i9TXAuROMvZnq
hTteOYA9ofgYdWoGHJOF/oGscJoMJWjWmmfiKPKMZn2yI6+fbO2DwAAEpsjb
ZmkM9rmX1O6xt8xtUw35V3he8kCmJZOcpwlZ098NS3vOYIzrVckSJEEWR55d
nCMCvX7+mrMT8Le7hf5H3LJxEuTOb7pnt1Jbr8C2yXthUhsj9Ce0GOgkBmsx
ded4NHoo6KJV5hORwzcaM/IMCeLpb+wGiPsl71HBhJiGK6Wo6bYgPIC3jQob
Uqm+gNqgCD3CFq4amBZTT4HU53VdSSBnXJKKQmYp4QxTC2Ut+M+rDzA8BXrm
JrY11deuD2bacMq33ZF5qiDQblDHXPfFNrO4EqtltGX5YxVmVllm3B9WcXPl
GHW4fo3rlpV1HqGFx6TWNow6HEf+CsARwwg6S7WgE1zSFjc4Bz7hjNEstU19
1QEu9Ebt86RvSTpVjsXF5YLXmxmUxD3pR+Vum3+bnic+r6i93T7geGH3s8zt
H56ZmXkmqIUACHr4rYzMKPHQkzTuSDrBy3MaBrAh6gaRnoMWUlRAuWtPxsYY
zR1TzRXc72uG3wVM/E1/f9alv2D6DUGJfsdNxYmUm4FCzq8Dw0kRHebG36U2
WD4ff7nI/En9Mvbx07FflyBVfIw1mUCHCPD0SCp0UeFG59DJJkTjf3ae5C4o
hz5Ac7zOOKVkkCVcJZq9l7tliv09fofW53b5jFmUQeO5j+JYfi9DWY1epR28
4zEI5AyRM3mLGaDm7dTMFmQbHSoJ98kjVsCIbl5q1hZ/4MIhJ4yVA9n5oszm
LTLa2mw7uKhv98UAoJk3UCG3dFPpQbk1Dzn7p2cIbrgclQnYa4pxAHUtx3GM
h4+4Z9fGtwmvR7LbL4n4T/z0DgMafY2+hsLoM8i9XbExTQC5k8aNK8MOHE1U
hdxvWJ3zSmzcn/Fk+vje/FbZ/kUK1bJIi5BSprCzJGxP1JbK+Bz/zCBiutTy
1Gsty9a8HtWhSux9MItx/Dz4jmTPTEsVXQwM24p+lJT7fsxTSKuNR7DfsSzF
xcbrcgEy7jdhfCtbJNXkPvnMYCuOuMIECQqVFIWKxNFh2UlWWxxD3JNon195
J+z+KQchcLJ3ri1+RYsyJiQH3/ldZUl6qiH7QZqVbc6lTCZbPkY2oUC7ILn3
Bd8OGecvTwRSpSLCZJ9/61NvspV5E0t13VU2GaKkAACx/tCJAAemmlY0k4ei
cLI2Uizk66K0AaRHcTxQ2W8oQZbjaWUcXJ2ROnFmwmS92RIgCPMa5uNo/AZC
OOWY3PPC+kEJRHP37EZYCTLqOxEPU/PCpKPfkW1N8D398ZBpbEmqh/WAGA6J
iZo3HT1b+QyPzNxijFZH/qZJELSNwI99cRGT9dz2qX1ZHsXdg9CDUw25t1z4
rcgPDBaqQYZbPNtTcXvC0WmgcXixzg10YvPb7NgN0xCccH5ijEMTNl0JHanr
PKKGM6zBgCKh1JW+dTCqX76Pp0mMg6wG7D+DETICS2qIyNxIR+DSMp5jM5n4
R7xq0Wynq1JyPPnYcX7QZ36FAlfdZ7uzGiOvJWZkEjp+/s/T+y2ohnZfSG7z
q0MbYMsfKFmsru1+XoX9Rf/DKX/B2UHLWy7ByWmTctjgYD4eukLz27k3WNf0
V4iEBZLIBu3SkR7NcTZfmH3mM9S6nIoU4Wdg3dS8WrDel7DVh15YrdlBwIgS
z7/zmbfQdaj/2RMB5ZEE55mQrQoDe/RD/gLo4A9f/FDJ3RXiQdIDSdRZKTaX
OqRx/M4AM7SKyxvK49DDkEvhRGhOW3+tVayjX5MDhsEw4T06oJ4mQiK9hwca
mDRt1WdhJ9SbYilbT7O6QxgNuko7bxMyn7gxP5banlEPRiUeKwN+u9rBbSba
VZqppWlKh2+PBsf0CvqsjMFOZK6s31VOadS6I2t/vsA1v+csApIj+jZ3TPOa
mQ7DzanRtU7mr1VfgRv5tn/621dIaFxSAaRi6LumlIE8neVey2O6J4sWrU6z
NzvR4KmxNhU42/rGdvMRMuWgWViRlZBtZLavJqdJ/9aASa0TjVj0CimZ17aF
IsKmKg76LQUt/BCH/kydn9sZLa2h925+7S0bQuU8Npzy4vZ5+Aa9c1XwDF9q
CQC0sl+BmpOFXw4KJdK8gD4nuGJn00t4rPBtFovdT52E3RbOyLxlYQJVNdR6
PJtqt//6ojcQONwIW2iE9iqnyk+sf6dhc3hjWYERurVKXU5Xulh0S1sahRon
iVTIYTKJAWrOUCre8MiPvTBOWBfiPLPJLFdkMpcqGm2Zu5SWZD3UwYw1rQIA
CoihWM/QGAqpibWAUkCMvBI3Quj1JLQ/hW9v6YXJ/US5DWeg9oW1yWpjZg+K
JInnLaWb79Jnl98W577KTsnuZfdFj6jgZKHC5ar6mJbYav2MKzkSPEZKg1HL
uzQwS8AZKZV734kr9wRqRuhi6BqIGwm6Jwl2q9qzBVIwZ2mtJFJDShDp6bSQ
FulcmuMXTzCVmxw/zILZAvOmksW4emjDRGrojAuYPug/CdIaSc9lKgwFWMjr
zg/Z1aro3M31rhb3opko7p/1lz5w7aFuzkIHpUtRYiXfipDc6vY+LS9E1TtN
1EpIfPP9JJXLrycKZ9EqPwD7wFO3be+1we4lM6LD0n5Hcn5NahEUOlc1DtZ3
3SqYLk2txOtV8rzpTmDOmqZRfi51Pq33ERB1XE7zHzxB6ONDIUg5/d1Gu5mT
L1cA7HjBU0xR4pzACC4/LDhkFqmbHIVxvuDVZ6gsnREqPqwws5IBXXWyaTsO
EO+SU/l+5QBdxYbULrmHlYumvBL9v8U5Tn3Ze0Nf/U0diTxqh6L0rhUdQjB3
1HgHnTfz6E6ipdMb3bg1c8xBpRiVGmQN753T5VzVukmtPCY3XR6sbG806eDv
3p8D4f6qxFBf4yxuU8w0Op+a8R33P8PsqSlzVzZncv0n+vMcrDygBtAER2Z4
3oyX6qqAFxQaHqGRkjjY8Nk6ut+ucOfkE8h9cdrpIbtaN9E0HPmUxpWs0R+e
Sh4s6X1JI5ULrv+vUuKOCELtkg2SGOQinuQlVYL9nknMVZ4LuemlnMor3dQr
Zv2Gnklpzr/BZ9Yv5YFAIN07txcR+3LMxbo1uB7mamWKLVPZ7nhjwUJdOPHZ
O5tsoPrFIpa/xYUuPLj/3SX7Q66sFsY6bXqoXUkW7HOwtRdKTy6n3ECPqRtM
ob+h8gMBe1Ji5HpqC57RYBzO6LNmWai3wR9e5a+pAMioYAQUp8BI8Hvi+qqG
eiNCI3NitQAiOta8vww+gyxk5XrxIv7BvdrHuZBF0FcYi8qykB0/YnePNxUF
V98rBbvO9fd/IZ6M+DfyXf8nWM61CtLczq3x/KSOqJtKokZQqekSdJKflxOx
m86uU/LoHh5SrKHIZMxWCJuOrfmFAVd3wSxzNkGNJ+FqhfuAGycq4eu4icIu
Z+9n0e5TNdESOTR6/MQKXU/F+5fcTps8qy9aSRW6c/SWVpbMw1TSYTTsRTZX
cQcpzIZMm6RsOc1vdg1ZzEW2QnksDZyCaMZ7iNVX+Od3WHHc4eSLSKCsh/vm
L+m0XZgke2gAgflafH8Z6dvwaoVnqUQ8+yoXyVa/UqbP2JbOjxxHMwPcojVZ
Y+PyL6HQLGH0BVnK2hxYYWVpX4rEQfhGXcMVqg28+vYRqALR598jtuWvOeQx
9Ck0CPlopEuVdFwM1jVZNyG4TD9jyzAOnQVBR9go7NHAEWP4mTZx3Sp90xGe
x2py1GBpP5qTtqsQR2WOxPoqPBy+iGIjPSsZ+MI5smJvk/UhPjZpKTnl0h7g
0Osa7M1nPKTxwrFvrUHhIcbr2VEw1B2qjlwzo4LxikPY5lWw625tFxyfvHZp
N4Y6Eu1JTN4J7cMKEVErt5btjRmDXixxbloj3fHSX9X5bFLfbLKm+NOHviRz
Pe3UnM+kkMTOeVNDaXPzZuQw9o9SSwSMXXB0YrCH46xjzAWoh+nnwpUMbyCG
cVjvRrblIOkSnfKEByKcaNSVnp/wkh8WslFa6FP0WTL+EehWSu7uS6f2D4Nc
3d6jMzrqpyABTnelScv0WfHcwR+Kba52FGC762Yks9BJ3J6+lnBdlPZiRS7I
ZSLg93QNJEZikjHpb19M+xzjM2IqQKp+0ZRem15BqAhbI62xLC+83Eo58otM
1rwvhSeFs+1sIacljr9Q5YLuaZVOQ+w52cR91uDhYpAOdCMCHXNUnd1wrY0l
TLfMah1ex4FBOzeW79G4ZPHYPFWXbU38o6NxVw91dLrWfbTxdQPJqjb1nbWP
yIzml57hzENpGE5ZJFqZOr+rQsPOhQT0adRvDG1hNTnS887GlwtZWIQDiQ5m
A3Y43guc3wfyoFH9zx7ScGCa80M10rP1fOwKtYLjPaKBhZMrNtlOHwcOl06U
hmS3Y6rx0XBWjouAQd23SZ6Fl2z2ofbVMYc+noq67QBSuFyACf4GTeRli3Nb
RLQe38PSPcaKMMsNUgGSOrxM9GQ9JvwNUXFt9Cq1BDAE40Rw68fbZYcGe/K4
b/bDzCGokiG/2Dyky8RyYBRY6ksjNBeNqo3/gZ1xaZ8LRk+0KRZxigU0iDU5
WPZ2ekPGx+PTsJDI5K8dGlLgoosz5i+BTd78lmtI2qG5yoRr9fv2C+Hfgabg
Mxbb5HoUdugVrYHmXXCaK8pqaCMeUJDpo2SODvjgWLEV8U1Wxwa66IfIKxO5
+8ZcjWrZ6fMF/fUCKvbrxxCZl5ZaKVYyBqvvvq7Dmbsob3lSNKEhlZGe8zZa
4nVNfB5hxNFxeyuL5XkzzPf2Ev6Dz1lf88EozDBg9E0e/Jh6r84YK0mZwaiM
/w3QULm4rRvpaHIcSTXxh04fAy37eW4mx3iCjXDQV7XoNm6P9c1TrMXc5sbE
To0kDM698+K7M1YsLjdZ2tVN/SujiguIwiQpPq97wftMFD3uKsGZH5EUIkRo
AvmwEqSvguDrim1S/MpZoRDR/Z10m06dn43omF+1J7B8dKE0ur4wHSg4WK1q
pZsPoSViU/52Jwd+uNVp17D992yG20d16BvleScnifwONZLISPrCMPEPcf3n
9JKBEyneDwH1FZzSwkKa/dZfD8H4C5fpjBjyE8idap0DpiWLFLkQFIMzX/gE
F43KxSweXy78dreRKWv9HuHIDG5aUizvOogLZNSk/jEmz9jXh2MoNYKpY4r6
Y0xOv2Qs8LBn/t5doIxHLuclQ6h6pZh2QHyfdlkoZ1d3AvKVzD02A8zWOsMV
iybf48fmxnRNdKSUemkxM0yBscUMstqkSGyuQnUX4n82N7g/q32vjSmB1HBq
fYDqMSRVcDUMET/8VvweNQWBStx5FhKiwqPHBlCMPxY8oeSPYP7uvZDY0OkK
NGiYmrnQ9gSYjLUamyx7NGIhPK3xhpQoGboOv5Wgh9Y3zDVg35E+j4TLj7IP
OwxSYb8f3kMZ+1yEJ7d9p4YivRPyo6JMgJRMSVw9FakR3Al7V/99uJs6iyRG
plWq3mGTqMwlaKxwLV86l0uUIHqh++Bbn6ZJFHn8uPaZv+Gkyp577Uwg2bsz
IkY6OVBkyXXJBPGQ7Bds8yS81M0HKJNZKFCBObzlshyFugkvleu8FSZH04nx
OA2jVEK+eMzt+g92PNILQtvNeCVzO/no6snn34ZRJWEC11dmRCQpHMqrv0fC
2trm7WYKnxiPSHDO8zUFM9onhmUrzK9mFpqOJTcunqSIIc5QAQc1AVYd37XW
bxE+X9rRk0w5F8hgss/PJWbcLzZ2xQHnVfMLzZck6Li9x3wvo9jkcuDFRwtL
uRq7DqFi/JGTOKY1gDr3bbZ1eXG2POLp3w1xKfMc7IrAhYfi+HVsrcvhTh2i
ml3bD4HrQSNVtNDBisIp1vZoK9kpWghh84eS9Px8WkW2acIonikKPGaZG1Bu
vZYP4Q3YQvjZtL7z/J7cJTb9sUn0Tpk8ePdsjl8rodt0poRlQMqCjckXHL1L
WwcMgVxX8WIm4bxF6Sg6dvS9uiEA+bqH6w0wJ/PCa1r8wLWcZuTavbFt9zvq
gjIos2CydfSuhy2sYG3AG3l56Dfjz3H3QUgHrLY9q5ryl7A9RPYJJ20b6NAR
bw4DvbvU9kGnQZqguQUa3xMNfLxUzdcwdkx5lR1b4ZhualaiK7EI9928PtiN
NM2Ks7sc8uo8oVyr16QHMIpkd9FxebxD7kx0xI8fbh9dA99N6KkDQZtJYi20
zKmx1taad8HNbw7DGd1ux9106vd26s9EaK+PCm8ZPnzgJGXsy3qNbYbEPSgk
Gld+G5BeOc5XuZYVg5uLlVoe/bGtqSBneoo6+hpQV+Qpw+mPgVu4J7SUMvhg
XK4rkiq8D5oRcZyUBNEb25NTrEfzd79kNuHZltRiFSE/fxtRYGozSLp5HMUJ
UM94NRmqvH/jAC0GAzJv13J4op42fLPyW3uyqHxBomQo1lfjswJuaZDgVT64
cco9xO37QLBwnoYwGjPrBpjLTQvv0AilzmlKSbN4aJD5gXQE7vVSq79cZq9b
bEiQaMZfFvSKMnTg3yMLW3un7HQtgvzlqbdH+FE4kCzjTI2Y6qDfGUXQ+V0q
w1n655nQJU3Q9a8JsGgPOVvUzskoDlkgjZq6Zuw1u8GI3vYMyuU5LKDsMX4s
ukBAJqEQ+DAC0XjsRwOUq/JRgYhnbzod4T+RatLn34s3pgTzo6MiKf2+fk35
/shgyVFVrpxvAur81qpDhn77QUYbVQq0Xg//WESQ24IYuJV7B6ZLaHdH6D5G
0DzwFjON0daVR4yBeNXgnwIwdwKY3h+uAJdNOh3jDunhH89KcXZWnJ7aGVAs
vYmMMcMIeQ6QId83kw4SDah4Ri0HLKUxJ7cQPIlSLPm7cjKB5hZmKavGUYfK
GvQZV0p0Mlc4bUH8bX9Cd5Ka8y4Rvh0RkuOVyeWp35GJhPTjYI8an+1h1OO5
IyF2HZyIWeIb6yGk9doVFYk1P0Hzcx/zuMmHG4gJvDVYUQo6mvcZ05uvqhkZ
FzdWDTJTJ1PUUpSXGX1S+C25g+B8oyualGcEas0MWEKNa2hLG3vP8losdPXi
4t9Ham2Uvi/+V0tKEAvS55RziBisRtNLF1t0SGVSQFniSzTErYYnrTtlBiNq
RZ2nW4JHQ7SFFGTQ2Ir1FN4Pni39VYG0yej1yXBYPL/xgk8veFgXornDIQ/G
904C5Peoc67FcARnKtYFXBRvQ/W2sqP1OMYmsyq9ao0NSzVw50YPpQ1ByUDq
XDsPPAJB/2I+F3qL6VP8t8DkI7MOEwR54WHGPtcD4Y+B/Ef9KwN4IQJzatmN
gBP6t3URXD1byR1bXHQAr4hkfCvpJ4gi6b3RsOpJ3BvsPZ7u76Kq4trAIOZ5
Uqj17I294riiHOlEfabj7YlLeJXNoeiKark/4jF5eLRcE8+7QuyRUpcm/M7+
UF4NrJy4asRVTYYC0L53xmjlm4m6wrIA09gbki7A9C5Ai9Of+xtfGHWbBm1e
doSmlqqZL+XjQ81SavV3YP0KnXE+DRghHXAbzd38Zu+xmXuU+WfRtxxYey91
6V+h5zjZqwZI8qSazMLhSmgH9itmdj64NLTw8w6uFX1hSIf1np6kgdZ4+Yjb
41f7Jd6+VX0eVuO2kVsD7plbyhfvdxKmlOxD/9kHWKvdCiJnto4+/hn+eGGb
MqyKMQ/jbA2QTiWMt5Eh5/qk+NY9mOjvgxBVoV6W/IiT0Nr+OfjsNIvYHMkB
Oqg+SDHjRvhcTqX+LYaHkyHjlWR5N+o6l0Zr28uPaNI2Uo6wHDMy3X3Cel4f
gzrZjWM92E6y6iEx9l6LLNU/6v6dQGf69OXw7gCoCbTbT3v91bI8+m3uCl2N
z2/quLqjTXOuCVgInGLt4UbykLjrYKqT+xQwjqvMWlxkd6dm/IVa198XBNOz
gYp2xUh/U50ERofaeTyDp4aWJnyHabZqSmNhack+3/CjcyNptDKouD0EDu0S
CIUsQeBfw4gzSU5xC2IoZje738KmjugkYIUSGahkQElCYBrdwKmIEAlLjC9J
G5RgJE5VgajewcRRk9nK+s/YqA6A/9tlUJj4bLgZNEzlrbooo3QKACYSXhlg
hWktanQlhEKLhlqsL9NJpTWoGgyiJsTjSIbzNlfuJy+O0RE+ovjZXZXKF8gV
DfhLeUuzuYV5Q5oqV6Ck3cj2nkknsojZ+tVq3znpTy4osO0aNxoFJ8pYHVAv
NsgG7/kIA24KEL+BS+SVZ349VjHbVTfa0/QAAcCTFU+CQFRZHgA3yyWrItFI
VaNhhCkHvKopKDOKPoS1efqBjPJNpOqCDFzuNz97yKjh/rSheooYay4J0LeQ
ACjY5NktYGtl72XKi0R+eHtnxccz574tUC9cGAqQgFL7jMEJ/w0De8mio2LL
1lYabzdw0ouDjK8Vht4pDEA3cKSmPHyPmnbs7K6GRoAfy5nXunelYtYlOoPz
NkNxgtJ+wc4ONvZ8Poi9r95bm6P/zwKeCNPPRXXoHIZMqLVtCUClriDcV9lw
0KdSBBldaf8kxdyWKifMv7BIG0Jj0+AorcFXmdd9K0IMVLjyKz5T28IrcJST
D89R6RwT/RoQe6hcLj5PoLlAsJpNYqUrBwyS3zOT+bHuDNYMRZCrD2d5idnF
ujOxZ/O227iAW9JPtPEyMROezxrAQVSHc8NSo2v7xPQrOicMIaiNkmRRz1Hh
euuZJOPI10lHrvGBlWXqp9x6S+DDVA3ILklUFBy2VUeOXzNjdSs4nWBiAQAi
7rUvRSGlwNsdLK3YwPDvte3WjGS7xfwboxFlvsu/soXk3GG6riKrivTDSCuC
T2CxGIzsLhAP1xMHz8amgAFHplcf81szkAjGfDtzEc7fX3fNU+nf8P7sPmP3
JHmynrqtMbrR1VAcJLymhtZQKTzSm+fleY8C6DYvJEKb8a0LCtevUMJBYCdQ
YHn3NQozhDdKBYc+LrP3F/LGen7z6k/RdSQbEBWK/GBlaqCed9RwFH3nx8hV
xieLtB3Ba7Eavygt1reh2GwDtu0Rh2ttFEDxxDp3Yhgc/TvtzOeEl6OgKywZ
OXwXJicmmfgj7RskQpXjlzcuTGsZxZqZJhvrTQ+0f9u9zfeMrsaaTSj924Cz
SZx9WUwi+ajuVBCqNJRJtyJgx+mfrW59o1B8vwc0anFM89Pf8Ah1ze4n0YZQ
RTr6CS+cxfR3YtRW8W+szxG9MnxloR9Exh8dCkDLsHBlhmz5ufxXRAmbPGOS
RI57/UzqQinw1h8aiJk7aWGNoLtosFe6oMw73qR/0ukHqfClib4MzXG3QMB2
jAIAC9AqyqKYItrGMigvsZ3Wz3feqyiOl7e3UtbjVD/kXPfD7qr4dfuBl31W
QKU4Vux1YRdffE/7q8tdzCmNHHfcvHGP6ZMryJ+vfyLIQ+w+qbTWFCbrjssd
laky/+kjn5xAyLd1URW+Te780fLrXJNJSK5W98zD66zjeo69A5Ff+3b8+Wau
dkh1Lnz6x+tPBCzlidEKDKoyPuCrp/ke/VsN0AHdax0JvbYV1qaB7fc4oGII
EDq9gVP0gfCQsFtuNoxzatxonijF6cE3FZL0earMQj9sayasqzcdp5CABUAA
BxD6hEh+01lXiSqdmGbSPTe5Or+5lzBKanb4rMgRXVuB4gxxmq2vxA/l1baG
ejD/DaSGrY+2w9EKQz5KGN7DABGBYy31owp8+uT+0s0PgX21+CxY3qZHhnfN
EBVxkHg9mjT0BDJk480N+xc60iNcvbvkM5hwcK4JgducfIdcTIQsd4NUdEV9
kqUHeLYX+c818QWQMccj9bJtfG1GbUuKVtu5c6z6ABxFzoqzI8Gfq+aLhwnn
xxuxiDZxUMqpADRb1J9i8VPmo97JiSbaOn8MJXy+B2+0EFdKqumYS3+jvCpU
VvOzLB3X5/BkwQ6aiQTZ4Z3lRyncG+Qgm7D/MluGBU4GVXnVFEQCEBlJywM1
qAr8SCzN77AxfY6F22cz4iEmXfYXFDoVSynO3YHVF6EdST52eSVKzVifVuvS
+IC0/1VE1d3dfAvLYcdFrTDouMak9RRW6BcCcUZ9T/Il1LmovMmt4VvP6bJC
MjgI8soCXEP6f0pIfzBQrilqdPK5FO9kP+FORqL0JQpH8sJRv+gYiF98fLNn
VmlBwjZtt++iSYbQpSPtFKduJaff2iAKTreoOHPlrkOva0GtZdFC38hYYVI/
0agVVAzEXLBlCxoy0jaxfdPyZPNSYLSjbDH82zaiu5REgiR/qYABjBB+UzFC
Nsyna19gIc42Dk5v53oXgyWnoC+vXR4QNwuQK4JgLAORsgclpBSw4LYJESGI
1qxkJO664CjKmWaOb1bzNrHABr2/nDCWik9y6U/JT9DEMrvmd1MS/afL+RCy
ycCnaTmMgxyfJRfwcEb3yUySH1/DKAjf4ah+8+dSnOnhXT7unI71phN3AgHc
YZdn66k4/Oxgnsnl8QxlF7kRq5SQITD6JoW/EdcI0Ty/h5MxftQbh+GrLxHi
0kGHfRiKAq6vAiwdZZA1gGIfnV8F4/HQ8JE8Nn9XOlkyLwwEzgqjJy5up44Q
O/qqvFcXkLWZhNO2lW481Ib84yP0euyQGOTdmicWx0cuMAQiYOPbsoI+4sjr
qEgp2OULnN/YgqNT0pHrj6fbsn+A4FTtRYdPT+ManfZnqCSDVyz+HBwXAq3G
lK9LnRaXDKNHIW9Vj0RVbmDAuUDsp8HsmQkOb/DIlSuyboIRYJK+8H4Xap9z
jMBq3hWmM6C6PbADpObSPx6crF6KI4WFPlyGILLGRCnrNm0RzY6XjB3WheR9
HgMq1F5kisHUB420HvjfkpKkpZdC6UduDrAW78IWI2qfLmKzCUMbI9Op13ct
u1oBCwpf/9m/z6gMsRJKn//HtBsK8wn16hxjwJbFcg7PogT0VH2GvCIOaVHn
kSkXJ9Q0/J1/OVpVnb0mDf0rSSifWRZ2m1OJ6HLGAKn58BFXZaoHp2H79fuP
pGT6MH3SFlYQsmOge4jzvvXpV0E+NKgtLdXuUWWYbbtp/VtW85DrZ0zSmrPN
Fl/cfj5fSy6VbgGlhsc6uuBhaPjwlqIMj0Tc+vmz4DrZhYs0fZVsRgYtlGgX
MYTFjnPLAAl855Z70XVjYxX28T8NCJwi9GV/sAeZSS7M4shtOWH4zKNO2Kzk
AP7OOp4kW6HwWvGM154m9P26RHJUpgb+zS1GimgN8vX5VFekPin3tAxeG71n
RWeHtSTWkaIt3AVumswks8Hwtnuo4tiJsALHjq9XZfYo/kIWpNdO1KUdVROp
SZunHlLWQIc4N+5h8+NlFfwtcjjlN1l/wrrVhxpxtpuOyV08LMf8GHlDOOw7
kfsoCkjjZq3yVazLwr4Wf9etu2Bo+VJPCyD/8y0N/8+vAZUbuohgjPGr2VcX
LfkQV0cjkeVnD3lgYLJ2zx0GRT8tIpQkfWchNl7NEPTtqUM+h/B4vf6znZZg
kWN5czOSY08WV4a/wbVvk2WOGAgM2/6KUra4JJ/6bCykkRiM78O2yrwYns9r
CfvQ3GMHr33GrVgECOojYAUA/l8qVtbArK8h/QMy/3WFicFuj3yPdNScdW3z
Syn/JkIdk+yo8P+UYlMrLgiLCQb40dBbhqlBH3v0FceuY0AftJ7iAm/WSvxL
HJOK+wICHibquVqLYqcAcOo3MPcKpWtxa69qQnkC4bZ9vMnD2lm+1cgAFQHc
rrZiKBcD+2yedoeJ5eFGC2J4L1GWO2gk0apXZ7OkuXg2EIv02MUYidk5SX2q
rej6gpnaJbTa/XbQsUegE8INiFig7SRFz2BvXxzn37zTI5c1NEEXmTgCk34f
YA8o8Hk/LE4dH50xiCjtruaPpm00y2mKcv5mdK4oAedqVOEXERixsMJvq/tY
PdFQ0O03jzPBbrLALSFGyP2YdEUZRDJY3aTDD/kPIu/W/rVXZoRmUgO0SUlo
db6bCWlV8NMQgg3F2oVXDlOuMEu+iMyTQkMYzH6HczxoNMak7xr50GF6jooC
NjFyfpiBKpi0kfpC5eGRmuk4aZ2eJ6UhDNKU439LS2/MhALva2E1EmjpKqf2
aUH7pYLNa3Vu6ne93Qo2AmmOVymEhoY7u8e3QDARgwWFTtfuQtBHmQeBbCcv
6fmJA6VyVhP0U5y+CYwuzrD/iSuHqc5onr/4smcICjJV0BEUVOR5cyZv9Fza
Fb4oVab2g9Y28EZ61LL8K7ZB6M/MKTXpXUjqaF287mZCZZtDvUOwDpyUuA0y
8Yhq/EY9ZoTQkXOH27OphQHA6oUq6Wggdco0vCt4K4rfa4tZMXWmEI8YjaWS
5WnQvNsLAYaTFEYQLxSGXpnWUl4MCg2sECLb3swab9sYMRU5UPloIs19JaCo
J45eX/qrNbnD/HJEJ7L1rj32ONAmJGmvaYPb+4oaBQz2VveDNrSZrNMf1Qtn
aX0KCejvmOrZ8sTNRenjbaq7BICHsBJ3p26cekvEWv+9d4hlaUOpByoFq8+f
DhlXYEiNGmIts/Fzuivt3oMi9FPG8Vs+kibOsCrwM2j2Lo0vDiqeFQyAxTRQ
uOuwcenlVJxIBgtbvWLIzSWgu9vGGa1/Y4XWLhPcGYiLYZ4jk4Q70E2H54qO
NrLafeztk8SUvwZhcMA8KvLGcHF6FbUgTAeX+/F7rAply842QOUJ3wMk/IVb
QZKsByOoL4up/cWaV5hLyeLG/3tTJ+0q9+CKJP1jwOanwGHyQx88PJsae5rf
bc8zvWLVqN2Cz68X1enKxiPywMIu2Hu1EPD2ZCqwuMOklgiDiyBwnw2hhNmZ
Rui+39ndKce3Yk9RK/IYDj6uknDoAYLKDqMLcaHk8MvU0Qi3wzlX9hh+1vQy
gkwlINyJwpTii72qoyE56ktnEf8HlyXfic+e3+Znp3LAVYZMjVNDDqvRs65G
/Qa7jzz173BOdpDeowfcaw6vV1QI2STtuYVvlHgpoOXsyciEGmFDkb37c1dU
LKMuDeS0yMu4mXZ8HyXp0HXV7bELzURfdTMbsl54nhgh/A3oX4Ak2wZL+Cnb
bO6xpZu/u5uEBvui1153VAfJfuoymo3G/dD9f0KPcdsyl87H1011aRfrELTP
aC+4Hsfr7JJe+yNl8LPqQmp9Eg3+MP50pnxNwiXAVbTgURUSJ0qXneCUrraP
GB/oaJLfGUyCajZ8ce62MX5oDfPwBKvsIBZgXhy3JBwBbiwVxnxSYCzkoMWw
AoTUT5TtH/rjcerzAMNFYPNWMv4OO8SDH/qLnDkFrGDzM/4g+x8LqRodN6lO
nYiqj3o4+r8luckl7vTK+CI9OQM+J0HUbJtRtF7598cfNMd9B35v3V8IhKxI
1IpYc+OJynaCJiFN7xWhRaKmbL46nEFJI+kKZhZj1otJhRg/f6AxFe+JRWDT
HCe3edcgvAqVRzucNX5FWSyN89cAP88EgfjtfhbK6/DweW/7bgU16fJZZULJ
Lr9jMsigQYqi6NBMCrWRsUqVU/iz9Bu97Ze3jd13CJb3v6wWXQORLj1KMAIB
i9n4zouvxc1cS7r0RyXwQTXAoj96no0gw+IR2sewnIsMz/eBCJzqCgCvu5Pu
RVfjdnjXX1vXr98Aqd+HheWAa6Hzr/vwtMaGtN8Cv0mh2deNWofQ3Jme1Buf
ZHRnxqUNcfo4q3EP5KHHTYTOLZrkg7Jpf9dUDVdjbWbMZhTP2WzjLBvqqtXI
EA385huqHBI6k0ai2wpQRZRosKRFxDjnSuSIgBXk/KMBCbsS86o0aFn1Gmlh
b+LzbDTR9pL+xhNSyHFlM4Qh6wJ0tFAFYkJJhwyAi1Ev0f34kRSU5asJr916
OD1pafEqaH21fpaSqy8l3kxrgdMTEGj5n0rw6gBNe/9gRxwrSh924f5OUGjB
Ts0us8wFsdc6A1JOoWuv8Jm3zFOj9Xt1G601KrO0oHx1nWkXY0uBHiyu3cb1
jJEpiyDDJslkVN40ntY9kkXBqQHY1HMJ0/jsNhPsfKGmwAauZ8w7R1J+oH6x
zFRAZT7iLuekQYONvTQFzB/3A+L/eCMj9+PiaAVnvFjoTtwkojXLmyoNJ2wc
wCNbtKv2rC0ZENxLhAqJBEvqDaVry3l3wBATEncxzSWoUgAe5Tg2tJBPeW7x
HQ7OYd5dskZcnyryeD0eau+jxeeJYrgZeVYjQNqD1YiypfQ842t7s5kBc+Lt
bUndzY+4F8LcrESs+kjDiT95g9k7Lg+i6hN3Ony2VA1kQZe/BJk9GexEWULZ
NQZrqLA9+Yayozg1WVwEfxc7oyO7yiXAE9upc1RX9XMKwUiiI1jH+B1YRRRa
x1accZkFKlUh2y9BaJ6tRNuu3H8N+hwhJwWidTP4W7ufxc2ZMZLTmTZuv377
45lGeViT9gzllVepBQ6cry8aJusoqm8X3cAyZRUBpEWUWV+hLY0laJoFGQH1
rajg2rEfsuLjCPoCqS1zhXFAaNi32HglNE+KHZPG5sVrXRQ+z8kUH+1pAVmv
hEY33XNhuSG4uRBP6XN8HsM43e/J1YXiKEEqAi9W3zBVIyzOcIEz8lTs2Lw6
ofAD1N4iX5R7IGgjQljJ3HITgBIPB5euBIoPJpN+Laowq/pPA9uXwXAIIZEV
YCn2phxqr5MXH2VF5gIxUP+I5sOaxd2K7OkfFK6U4DE12cAp3ANkyclNXXBM
LuYRaU2eb9AzO1ujXrsSHTIas8DS13F8bMoD+hoQFAhuIWYj3nQW7P8Jeo0x
dyuhhQG3BAAEX/RGIXkfd2GURmAeAKVdASf3kuSZu3SirdAX19vJ3o0Xi2/v
OM4+8JTjCtRPdCZ3qvkLNNeIhMuEklT/5ZEKkLS0/gB4xktErc65YSJjWEoa
ccoF8rsBruz8XiOMKgo7gYbFmDrDjG067ahKW3+9Uhab5Fu5vdi/m0aDqhNE
DkrOkuBteivL4ztvCACTbJhT3QkNHVIY7VIGcB+cJyemiVDM356i9k8vkg28
zKRwRiTTQ5Xn2wJtsSf/sWQEyEH0gv1zTOmWvDjk8NcpWQ/A9hNL7FtjhFz4
8F6qiP20xKmbeyM11/asTY/0fLGS9RM3dwrz895FeV2ZYxJ5oG1FAPubEPyu
MabSG4JlaO5fJ0xCxNsUQ2ewx47BErsym+VsN9RjRK+kddzBBGsAZVJsn6Lp
NV+vQZxoUUKa9JbmAYLvYRonrPLiYdYfnXuEaKocdA9xUH3uxjNv0rJd/JyL
lxaV5M1i3Nw7k2d6vbCZET/1AfrO0j7ll/Ile09QxsHa4tLfBj8/kPNGR8EQ
xDHsHax9JoVB3syXNevd6sX6lL0mUjILxUILfmX78k0ySipxAd+kuHExjEen
fGt1kKB6S8HH9475+fSJf20l13sDXDxU+le+AvSP6di2Gn8/9F4KuMVnSYnb
rsfAgyH1tyUZNZ9Ijka8CPl/OB9ZvHmn3MbXf+jZZ9Czk/qlK3Y9iKBdQeiM
XkexqoDyN6U6FMJkKqgVLlts+hypb7mSBRy9jOiJevgzyp7qClFBQkWcWClZ
NYH9IbutnfjI1vcFkksUWGVKk69FXqp7gDUFQFLdrPGALShwryxYF5ORRkNS
wFo+vid/khfQkFLRBtszDQJsBF6dBJXF4UytbdiGCpXk3ZIwAJoLKxaRHk3A
rG/lOF+C8vCELhl7tyN7Iy7u6BCuokcCshIKklaFxTmbTHdDM7VDo2go+JqE
ysKd5a9wP/W33E01bXBHmeBWuXTtmoNrXEUfFejMF33hQamsQtNJZa3IDdBS
l/6LBwbPsHBUouE5C4Hkkhp2P1KMk0eD1TbD4i0/upeD16H+W8/UtmevQPro
gVI8bIN5G7KwSWT9xzmO/wCUlPnIxfjOg/Mm+vNAPAcOjMJHsTKj2wIq+A6N
biE/rLr0GfYCnYtBY9xiOBNPOYd0PzfKyaeb15Gf/srU0HFtEXETa7V6iENQ
YhIBX75GZba7DWm5daN3/ADBXfz4FjSgMr+dEGaefExw06taJQw2QTGkyrNk
qeuR7lhrsKM1AOB4SMBmRDWPzIjtm4rk82FD2B+W8gz0SGrpMC+FMrb97PCH
OuAG4zkmzaxO4EmN0TmXwv6V4Yy5I0RmVlPG1o6YwM1qwN9LF4pAyr5rT0/W
Q5VkmHqUO6qGIHYnj640JgclHi12LgTjlkT6/chnoiDoVMhdBCw+eDqsJU9/
63BkVRQg3HHCpNjWxyuqqdatL0iu2DggqjVVf1TTyNt3ohleYdT/UDKfKaoC
s8wK4XjnvQbquD25uwVTsRiCk01CAaPos2oOPN9xFdY9SDZl0LnJP+oBbYrm
i4qNvSifpwTludP7W2ItnzZfdheu12zci//u++djMN/6VwIpKv8ccGb9Kixq
5drLqLmp3OLhoRDxinppi8EwR+tBzMuVPUOywVnKOYew0+zW1KxEY0iRVL09
k36drVmwR4kOnAdDow+ZGZLXpbQp3u69OpbZKhOQj1VVnbMEdfw2ua++DGVO
/dPgjTlwQpav3DeIBlILRuWvuuQhWny70umnbfrzEld13sUofdGl5ExNkr++
3BYF6Me/vl+OuGEXM3nl8JMzXg3YtUIL36FHTEXPxvBS0KY0H4azgB8G6n0g
3ADRvYx5UrAHHyRM7N8AYScrbIJ532k+kUFcA7og8Qf6Q6SZqb+FetTz2kD0
EeV+HPu7zf0iKN4EY++yRju28IsEo/pIo6f+fw5aBzpC2s6GqJ2ZltHGBaKh
Oj0qCHD7wSnGvktxSs5RKfJm6AcyFTFeqjQmyceEgb8Jkl6jC8GK1dvyMdea
mxXF5+wL51Vxgfgl+b53JjtTEvFJGDhD+AKlltAi/4BOfyPpAb9dkFMUGHVr
E0mtyIL9ZgeLdJcQEFDKcDFOWhn6VqVxb8u5Ar2rTsX4ydcLhQ3IUCvhyGSb
wKnbxA8waj/Xfz3dA8Mi2AY82bgNeDu7w3koeuyWNomv5Hp6d/B8OecHxFfQ
a7a9Dxo3JZg2ZAGGuyYf3XJV5AGFZF/SvhPYCvpolIjh9ie4Z8GJSUfrZCAS
zs0R4J3rGy7WQ4ZC2790MhykYFOPka/vFZTWmma9mptqfiECd/dMlq6yPYsP
V2OIU3wF01FrGjrQpgNo+2Xuqtj5z5aZ5aenAPL5X52UgJh8RwSYwdIGkB7b
hrrzOhWtptG28I9H3xeMQip5tXCZx4KQXepWJiBB7HzS/AzhvlcneDgQAgZg
Eo5bHmdF+yWstx9cs8IW8o8/RtCEcwp/WedtzjaLE2rz8Z3zFy5umX8L4Vx+
UpnVYwSOjAvTioa6Gb7ltKgSsW8XwkmZQSdnC6hFK8iblWxN2reryEIGrmxO
gfpW0e8ZbVpcdv6jz7XKKPf2XHaw/qnFETtcB6Y/iNV+rYwM63+A+qnHkAGy
C/fejEOH3kdg0riqT1tVVHgH4OIzQfr+Q45f+TQXriYz34ehQCbh8P1bY3em
yv0PF7LQ5Q47UzCmD8AGwLjfvemmgqHqnCFOIbr/asXlQMmpYNtPMw1L8cEi
oiUzj0QxVxSQHKfjknHjYMQExELd7vwSftmnIBjGmEuB6DhAz0HTC0g/RiER
l9YxQFsl2o/8AGhMXeLi12/AARG/sJuwkMDk+bALs9lEQ8kKAO0kxLy9RAN1
pfthDPCP4EAyxZXqzhEWQ6qwYpbQS1k3S5BpAzAIRvAuqGNS+vlxbeE2dqOo
ZQ4pRajYdsiGjhlvKBYv/gwrm9Ahu7s/yeqkd/cPtMMHj73Nd6RDzbLuwASn
kW6oSqn3qdZpoXKL75z8lC2YGF8DbKEjH5ANPdsahYR8Mc1izjMhdiFoYhBS
jLcYOT5bOTpyyTHK9KTidxtpJOO4FwtKJzaKvhMFS74LCj+rUQtHey6xGZh/
PRz/snO+XlkLUzqPPyFVe0yeDz0nClq9xNzcRfJpbWvGDQ+Rme+JlSLYL/PL
ksRb2Cv14aJYjJghN/aPHxjb4XtVlBFL/dBpweg6XaavBbBpNwqSX2z8h17C
10AWybqrbLRu7Hy8yQXSeg1Cnx/RoAfm534KNnDHb1Y7+ZeeJrp1ZCHiGSMn
Ii9ix3sXTaX98Enx1OKhKq03S9/GBHWaNGr1uJZTAklDOQqG7I6tej9/EHO1
MmBF+nwDI+ZHcpkT4olB8rH15kuo7pMVLfZIUIkq9yOdfx2EBqTtyVSIJHDn
2ZeAKTdqLvuNjnyKOleT6t7+kPMHYe03W+4+M1Ep5XaOCWM6Ytp/WATrBWCf
UXXMZH+ga+piHbFp0VU2IXRZqdQixoQmeGchc/S4q+t4JFgr910asa0rVxMC
DbdGREFQ0dETGTEyFrbq+ok/WWB/Cb8PQfdpVm5DglRfOw7vTPE2nfYqAb4n
bvkYfIO4D3wh8LwfD50pv4G4ov5lFPgTOqAydEVgzM+ghi0ScFQTgiThqe7F
RbliBs5Y97W84bavxroFWK4aBcimBvne9/39ltWgPWJCk3EZgMjEGzp0yLH3
KjchhV4KkG62GNT1zEbge+PJvUSd4raC5X5MPYEjvnw3kz6s1yuqdU6/9yaB
FSjp/2Z2UMl7BTEWRU+xSwNXhV5dyo1xPcM2aXC/rM1iRXWjb/dvaes9wExr
EmmDkOZgS+HwANdwFTGBOcF6u9r7fK7fvKHk+ism8ONiIKbWDnXKXqpVNmZC
88t/BsAMzfGwB64jNrjmZWfk3FOmJtCx4pB6Dxo4I3+vtQUzRX/1OopStTVC
a+sLeim0IFpr7Gssv/k6+/pHMSv9c0w+K5wLcjJQOgcDEidLMrUMMfQFItlu
8htSudPu9ZoNgyEpNUNcXIjzUJC+swBIJ/6gDHB4RV5AMrH8knp+u6DsKxxU
WxS/evY98PMgfCp4R1I9WzaVqNtVDe+xOVu3uxRnb2p+4jSJBgiY2NVAmcYS
rthjH+UiL9lwGpIM9hRTX18vGWcpMhYkXw9Ez5ltfyHqbJ/lXbRKjVZc8ygF
4zoOGbV13KghqroNlHmx7fdGoyOCuMuxinqhJKWkaQSCK4FqMO9GNxLJMcUb
F/bk2vtDDBnMO0V7cb7+C3QLAPpjFx82qWPhN1hTENrMM+MaqDJCunMMvTyQ
i4Qw2ZueFo5FJDRzXEnHrSZPFIDeR4gkRPxeRAlsHCgI4DpQxnjg8UCdWa73
Xf4CUc2efXmNpTjDzOMJCdMs8JdBfjl1CjcIQtdn0eawC3aqmOsRcQ+tIP6h
Sh5l90VMI+St2t6a7vemAk9ELS5ys7SKsL+RWmOS+BbgA48SDXXo+2Sc5Ch9
24RUfvAqsjD88qQ93REMvpR4jsYDc9Q/GjTRKhKRK/7LO777d0Y/FhHV/L4R
1+JPD/OwAGKr7T4ZQI0SsEsP8UH0mr8riXUXU2k91l3frCf3dV22htLWhaCv
7tfEh6TWu/aEDKbO4OcOz0cc46dOZ53G5IcurIAtK3ixA/ntIC4qKOsENzQO
FgDy43dGq/HVyfdPBHLtVUg7oN470AHLnagHkFCrtROs+QSXlm35cn77Auq8
h9jmE7CfUZDN/yui7UlPlLqrZxhXQkMBY90ZmENv4fXmDFTwYBemyDIDM+aa
re85AVMhGqW5IAmt/GydmIv9QHockuldzMWNwOlF4fhrNzal/yuEl9ieRfgD
NAmaZkd3oFHPsI4K11DytCD6a/0KpGkChgknNxL0wafavyDkHne5Fk+OsDly
cbF7DdcUCvCJyCZKb9pye67+RNIRFCmMN9sS9zKoXWVik5m/+MAoHodZkR5i
JJYJ+vi9xmTpTUQoG5ZpZ8bO9/Yae/OqiNIC6HVyB+6Ouq672/NMlDm0njh0
BjErTLQtSwiGHs9ejarY78Lhl5h5LOOtBmMfy27a4qVxyIpFigKZXZ1Y+7G8
/UimYKGgWhoa9lFiuXXwYVKpuWuTq7kEKpBi7zKLtP2Ca5Lg+KDapq9LsBWS
jhoN5/8ULm2EwhhCTCgpPCUakCxbvVhPlGutCRTGMtCofOYlY+jU97tRy0wQ
s/h5S0XiiDAoSybfa5x3XzvZ6X0s0msjNSAx3D8SQB0a1+3Tp7J+svAVANwt
POg1pMDAzpRE/eun+GLaX71xU295XeNkw8PfZeqbmJFWEYpHc7kcoNSxzD/0
Ymv6WEAwFm+F0jvjB+tn/BQM8dTADMgZytw9haVmn7ySQ/zU1N61ym+0r96S
7QhC7KbLDPwIDqbeIkQy5JMUZSD/mT21ve35XMzwYDUi8ji0MIDq4CRyE6Yh
0y7jEylku9/mRhnmyOEKczFWWVxkxAZPSqy2I5Ih1us5ZqLLvZm0THLPgO62
c2YrQowUYHtQi6G5lO7lOxjDlk4tUocOfesbrMc9VnrKOjNon6paX3RvqWNW
7WbrN3ImRJEe8/5s6S1JMVe/Vf8qPoVSRfflANYYDHmcksxuvQX4AAW8rt3G
2YOsOsCTpVQt6AR50NESzKbYHJcj+MBcM7I4Uy6rYa2BYXzqdHh1DLxhOU8H
2TzuRmlZ3ywGvnloVClFeHaz6qD2ql92eFs1flY0BICGFL7es5JRyjwuEHmA
17LGnR1P3EF5cSt9cA7uYRgnpKloC4y3TRlN+bqwN61Rt9epvPEQGib0F+ql
ymRlVf74OBxFXdkNlyPvuHpqUNAFiYupA/h9RP+f4qXAGBJdm50/c6+IVd2E
sXPnc67Mk3Jh5eHYBe9i0q4cass08LIoHXRc3lc6tc7SgVKr2Ppz8SXbMGFZ
W5Z6aQPB4RU2u4haKjnjQ3lbWAp6AkuibyGtvddZg7zWZkWtMNIqaj4xbxJj
E+mgTTBmTX3RSc5TO42Dt4jJ1+k2K2tVPRC6xNqpZQQ9fF0zrEehUi8IlHIv
sJ3V4+qv/yTkwTB2XkA8rX9w2UjjCMkacO0p6msTS685il9fvTLfdTftsJJv
JN1DRXVfeMO6nw4+FoKP1WUG+cEdEKp2kf1liDAEFerivLCqcQH1mHmTblJ/
W57G571CxjBSs3UY2UKGShPoxCGnKvzLXexQN2CpM92EULMHts7g01Hg5JSS
FnPwGlpko9vsKRoOWfoRyh7hshcFaGuj+Ri0rJAd26Rjn3sfu/YWG1tgiE/R
Btj4W2MG2BOtgxokJKClEKcUEk8/UDdwQLsJLNzBmwfvAsYM4dGZH3H6rc9Q
t2K8COnRnu2G4yIaQiPVBIAsLOQgrNPJq4YaynXHJ8+Wj7cvjcPfJJAiPPMw
1f8gQDP3b222f6L0zOaWRJn58JMsty9n6v+c15BEZBs7wAIAA4k3uyK/Vc4Y
DEcO5IQBpklsUyt1FRJI/sT4VMYItolc3q4adO3AC53SOIWxeHy600GYBMCr
5re1X3DgdRAVAmEqkLR+8xB6jCDTd5S/LkP1NaYrZFDtzaUzwdiTS/Ryeghb
j3iCCbunUb/cBIuQY0yeFBV6NxUei59O9H2cJmY1dlQzo5iI834KxKtPY1P4
k2S7SpllfZKh5SegeQPWTCX+7YkR0+W2TEjmvqh4O/+EIK0wWTfUfBdWIei/
HPr/Pf6Fy9rJ5xc6Pgd61yFOjnB5i0MFFxSB7KJQv4GXZ/wWBCwXqlkXp5Td
J+REXxZGlxfSpYgeuw4u/iUN+qHi2b6bMB0kuRgjaurQVlJuQjPN0LQVaPGB
IOkMLEeA5pG+VqDkPQECfcXaixL9DgJ09ae9ZmDVZfA6bQiBkLor2Oh9Q9ki
GfgISPJWBNwUnwUpC9S4555zZT3IRgXHaWPljEb32wO9iaYR/wHdhmMevOUP
BP01yEX+FMQePqkV6JED1TRgZ887Iukqts8htwlh3HNlOlq5lYbfiWj1lQJZ
9gm0hdtdqLzgB+HSKXlGqpdFr1GXVdea7x8idCZiU12axgF2elszPGqtsDB7
+1085Elf1H7DNN3bwWWWd69xmUcOvw+KFW20PGJUtDziW6CSD/2OQoIp7dPv
ab5xAFYmHrUwtccr0mzbCjBZa7W5IL7qCBIzof8Vza9kJx7VBGZTQDoKiwA2
pjdlov3S3bt+ni0if3nrlOZyrvONE4OAPK0Suo9BFMNN8O1nHrSwPfgkPbUh
uQRWM58yPThQs/bNJCwmlcUzMG47ssdBukCumD2g9CpeM7MYeQfpEAk/w1cL
3cJKO9cHOhf3/4MTFIabu+L0F8460+k0H4OPrnY3wNQKbtwf6zUMN23T7vyz
J7lfYNCLFS4fOBIlj2vJIQZdbe/05/vzOAsbahgwmDf0Szi3+9AHzo5dkWMv
jzNOx9HTXuGDzA+dQiSwAzyntflH+P3P5zuvDJmk1bu3HCfsEPbN6dW0sZoE
ACEIG69eW0bTpt5ZI4aFA10vhCTxh41enn5FOq6Hc1YWABJ2I2nDwt61LNHl
qQKh7H/0sNPKqjWF4cQ6vsz+eln+jo9WaGzDuRlDje3/sKjkRdkkbYRCnv0z
56AJ1j/i0EThj7zpjQFAbvSsXDFpNP3UWGeMoXPU2r/owUo4az7qStrgxjF9
oh+xZTBCUdQXdZqBAXUnNhMwN7Qyh+uBCd31Z7lU6TOYmZVE1+eKs6hBhYNd
Dt6f4U5WkGdeXajFdKErJX3dWVmeWcFQHpLxfLqlBYRQptah0ObVdd3l0+Vf
ykZ7D9ExAjVUP8/f2o+QMuBpDNANn0X4wU71t1jkF5jJDai3/K6o7pBq5Fs7
0BSz8oToGVr+XqJcUJB2OlewlHGIrqhLcTVj29xoP6LGxvrF7NfpsOIgQGQE
gMeG3U5QUXs6VwjpPozaNpqDsH9JytNC5M76fgmRTSSPx6paeCZc4d9Ik3hf
aq4DKXXTZUXW7DTPg2mGE04AZDLvq9vHjdRtsBnZzHW5uvkSREe3OoztxwLd
4EOh9/6LuYocFzNpg4hFb5hzwnSd9mmhDLLAiOUa00udVvBGSfDizgkoa/Oz
WoXq3BvVJ2N77vPjFJq6JqHWXr7LLsX12dDmqAmWa48cLbgQppFwRUJy8FAz
jITxtKsHiJIONlPFFpnShoBvQDFDa4UyEiyaYba0BtVySJW3i8E1hx94CnhX
EHJeQhtTrroo3S11YDzjFNI635JicToVvCvz60T7v3MHM8WFR1BVdWu33XkQ
39jNI6ba8mxkSKNor/gXFOUcCJQLZgzrG+OC81XgFM18SjowbEAJMjAP4h3u
gLWNbEPHtUYKZSY6AMGc61DRy0SgP70XdmN6Cn01ssEA7BpbAMc+CcZXj9DH
jhUjeL5kUd+7dfI7RvHqXKOxKUUDYcoriVw5gqKepjlfsKp/H0eBKRpzzRRR
qYqw34xJSp+MLM4Sk4hx2sGE7mvg1vNr3aJoN6PNMjO0Kd5FGgSry1B1OTTx
4nuhS7N3DnVKStcao3Fr8LXGKlK7M1xfFwUhw6+uLjbo/lubP/b1f+eBHAng
wATx+17ALupbSTAiJEqUQBxgMsNdSfIpEarKkFc5i5VeNI0sonK/EwcxCNBM
4A9n/IS+KGJ4c7cbcg34oN214e7nwvvlEqF48D+in8oRRf8OCk6AnPQ8rFO3
OyyE88HaYoZa+PDVa0cH11l9oZz0PRx7BJeMfq8OBLMw8Jy3bEBsQ5QqRJRB
ucijFkEL9v3tZqldR3JpBIPtIvNkvdwRklSe8lb/hGL2ThlNOMCHOQD1XD5l
ZyR0nnnD6MFa0pKOKqjOtXGcYDjieXryPeg//MflAL51h5Z3H+g8FhbR+JiF
ilLa6nLhX8HB1J61R/8f29EGKjcloYxzhZCqXGa9i2I8SSYg3VKouMoLXA4Z
duumPqn5lTLQ1sZGH/0fW6gz7t5qLKtC11Cy8xq5ABo6nVeNebmqAsOY9ocf
hkJ+p5CaxIvmNHkxYpIFDG9orkKptlpLP/btLlLqYBCSgNQ8PYL88zgHH+WQ
mTu4f+CLOtNiF+nMtehw7nJqQ6MXrO8SBR2kFmJCPc0OLIMoXQ9twZyhUlrn
yZ0BsbouX6MQSk7xgpc2jG0FJpPiQPQzqihvafM8sugP1jG2Kjf98YyXrDcL
dB7JvfLrwsLnIH6sU+haan4b3fGDiu9A1rqLJq2pCDDCuQCC7L9LYRmlCyjp
8WFZskHmHtsUv0zUodGZ7yBbK7oqHyHOIL/yhPQ15RSoLZiCN0XIJKLMM5vI
gcJ7bOGCwmOwgo9oae56P2yeO5mcWOv/cFGldTwji88+iYmywZqG02y7hSLr
r7FpnxSN0B+LCKuAypeNpskruiz+S42toWWGBfKaywqdnRNoivSVJJjB24BD
fgUEM4DDr2gyeXTr2bmTAhhima+j+Dm7XpH/9xq6YOL2OhNed6DldM23D9Sc
xl0ip2lnUtUcgVsszG4uA2nqZzIuwQpGxeldN1Of1eUEfGq1+PBlcMYqmr6I
CpZmz+Agu79crsl8w/U9CqlAbI64EBuIrVAEinKC2qm8za0Ie1I1H0loerri
bdXQJ/gaA4tDMx/HlhgWBci68p5YtzpuBcui06bsFNbWbw4gcMxsxrbTJMjb
r2CEhlN3JZtDiNkHmmZx1FyjaodUEz7quLjnsWmAoGGYX4SyVdF+bJcXW5Lb
8cfh8b3TgEuDxTGFKb3Z6214TH2BSxVMYbrw75Z4MdhYKGaFhUr12tRb9nVC
ZppOiP0c8UD/zpEujoNE9Y7gJkAeu+8s/1WAwg95+4OGU9fO2MbUjbs3u9DP
WurnLWB4Cvf01glM2THiR83JbMTfuKMh9S6zs73II7nbbBv30ztLhpk0IkaR
bXxhjpyYCjSVBFxo4mtG7o5O5jn3iyHA2Bz+7rSSZUHU8DP+Y5wXhC2D8MZR
2tZVu6L4g7dctoulNY4yqBpiOHzswrRiI6v+ZLEkIy0Dm8h3mTLQXZxlfw/8
YmvRcwm+tRrAMyw01wID4qPx98CYBnHtCtLQDkYOMBVP3B2xGsM9MtA1OraS
f46q0cNrVNNZcUD47Ujd2lKJ0llR9tEAS/l93LEHWB89blb/mbImDuvdd7o8
HHbhYYso2gZcGDU9haLAZH+2+ghAmp+dCdE5AYaoN5JI7wwn9voYIoT72b/B
/W57uhG/dCH5NqX6qXrVR4vq8OGRpgbp2Y9CwZR5EZGqwI8awvdn14AEdQet
1oVCqUf3BN/ZQAShzInb9zbP3Z1Cp019mshTrDgB94GnFRoQn92alroQ48KB
0j8JZ2A/83UVLs8LP9B10R3y9K483WKSKepBUj2KzJjh2P4VhdIO0SCr2VT+
VpH1tXvj8cq79aN0TJaOAF3V7BrhJBdvRXA5M//JcbWLZmOR0ynxBNbG84gY
CQOLcUpFsrjD5+JLNR4U/OlP4Jo3qJe8ECux/3IlQiAJNHaXie+Fi4VDn5YK
8Mxn4kJnvdabCbghTrKv/QRVd1Mm5er8GXpoBMnvrVjKM2Tf7W2WJsMRUSca
oMH05kL2Q00yJkRlwTw8ZbiS3sbzbTkmQcfXYxu1RyHEvi1jKlumoRzDaAww
Wws/D//1afC26oIVH+J+xRqCET5bzfdPjSDatq14bZPUe8NXJ+cq86bS/UoS
ShAWduRnYti4q3bEy5qKTfea4SJMS3DmLxi6ITxfixvTmwoZ4IzO9w0/DuM2
xKZwCFwZMAoWAWCTRUAotsoTlRj83Y+5TbtxDVVbyfmoFtrMK6yf4IcxmRzJ
K39FIDq7fpChggPmdTR3emISN2EoUoQ/IpV55EjlPZpQM2BWWsD+6zkJ1iBq
GIPUr74m5cyJiLdBQwFFKjRVWdtjiTgiX2Vv4eJc1G4iFGIw98fUv4B67sE7
Xt3xsgfTsg4JzEdaUb89tvc5FuhVsWS/vXeRRZ/2t9GLuJh/o/igrltrADne
EO4bTu1qmBgwEMEjBoHBkw+pbjNsntFjug+BUjgQHRSQpiybgfqt2hYLl20n
2PPfyyE6VWcbTxtFQyb2kZYDwvP8XhKzldcKUvUAtSr+PT0Tc+SMJDBiFUko
7Yffm64EVSfDg0LvKOcgWGd85FlxwJ4ezJ2/p5Kwp7UF9p8rHRM6wZS5v54f
z4iprRseenD2Y9iELSazR7EMnWWFE1Cv3LbeO7Sb569TGRR+m/oTGpo9uSem
hhKDvtC0Ln/i31XKVWKCXaHHfNY8HAsHr1kNBbeqx5YYr737ng/kZ/q3Hfcz
2PV9/HEvrOP6nY/Muq6HQBOwHoW6WvdsZcrEj33W631Mo3Gvaqt2uPd+ODVl
/nK9KFMbF6F0rX3W7DHQLDk3CbBojPnpEA+yxT6smvTO29u1FViOK8+EoLlk
4zk8/ybR4kgjObKkqg2bMCVw+HLb9qtgneKI2DboJEK8Jnbu8Au83svC5AWv
N4QOgxFdt+8qo/jYrcE7iLvNsaow0yt14DSlez+eegW6mCEs+LeFdzmaEkHD
DgjFzhdReMdO9Tior4mBCUxs7ylbFBm99ZGu6gGafReJ7FiLs7cCT5leJNTR
tujJoMh4LUta5hzhVZVr3HetQZEGjmYZpcxr1PM1vlOejpSKN4szDFuAsro7
T/eH/vhPlWIuzz+1XR4RvwGoNcFpfqpLeR+NSem9kT53sVcon7SzE7FObluJ
KRk6AZcmNdBX/8PNrOlm9ekEiJOpSCxMtyULzRjoA+I2EqApspE24+pZqEUs
OCwWkIG5M/dAm5cgcrapxcpfQeRRtpuKRgOQe4+qdOVnzsnh7WU5WwGrmJRX
siupv4Otsb2DWOrjMi1Udgcgo/ns3v3suTrmFpCY3SpZaon4Bbp5PcdkcrCi
l8DMwv9Y4QxsC+zV9D1FBNDGxsPKG3xJGrFfK25CAkqWRm1GuqMaDegmcaDu
Z1ELaXLEmMzA5Fv2YAq7ENhXiGOpeT83WP5mEqynVMi+b96JORFpUqni0OiC
xv1NzTS+FVbEbAn+ft5J1h9psML77zbSmRSuiUjMC3E71MsfNs7OVx8quPne
0s21Cq3F5ofuA6ZJqssKCuWBoHMW9SrJdxcsuFxtFnrWxDtRiImmquSHY+E3
nx0WOWGff0dWPiqc8zDckrP8xJ369222K1SGUGMB0UI3+mIwkQzBfYLbUOgX
TR9yS+PPqFTwe3E8L5o0aSYLzyY3220eNrDIUuhFq0x0/oVewsSqsE4NVXWI
Dg+sNIT72t0NuNsMjIlAzwp0unLn9oISDf+Swd0guxPv4UZclSyjISlcLw7y
1aRqhyyOPGF+2s+M2CscoIziyfWvSKTxUY8xvpGCvfC+AYnnsayXoAi3UBMz
WTQVMx8GD9ddqFD62zufSCevOjGQIvQsVAp6r7GtU4ftQppyy3cfqRwywY6R
aKRCxuBMZwNshp3IIC9At0Ovt+JiU+wlavMPBYHz8wqLLCPSiBfWM1i1N1rl
M2+AD+N2U0XmVImynrJXRyq4TFSO3pFlDY726rWYtLIBKNQgO2CBrcAszuhT
fidnKTII5Oqtvk7xalV5T85g42bRcRVKfPejiekXPYY8qC6OnWcwL/V5UCu7
VeC2cltzzqgnrIdXfLoOiDWPd+EJYty1UGe/8cKCjh1wN/OQj3TW5Hqi8pQ4
UwiUsdcelcNpZ66zWJ3F2jN/vEILMaqko362Q2w2RCLDdI2URU+ZgaAWj3SW
2hxpW+4v4fLUCe7iJaPeH7vpw11VslkPGKc7cp4Am7wHR+tWNZeUThx9hoQf
/FDW+94F5Jx1dacQ1MlKGNJBaLaouS7NjOIzEkvBddNoq80KVYmwZAfKR7tX
VdXezawtXisc6PBT4eY42jTvudcmjCZjO3I4MBDeOyBzN85iY3hoUxt0UPIR
17ojp85IIG+xSbuyVjfKwz2/dRMz2J/ydoZmoZlRUc0Uj2kyFjfT+Ohnoo61
7IzLnlm59thRQ80ScwTmD6gAQPLRlrsAhMkuB+furgRFMZlC7VweVq2tsY7l
95NglSSuCOwvE0ZXLorFzbx8mcF1PXI8UW7wFg5oreLH1WuJfzd7OjXCisAG
/dszVR0L/LI1t0kGOsP11EfZMaTtqxFs4KzdKTtYGnWNoaL7qXOHihtal2Qo
8n3sU1v95uQ8iWgjxhzyglTHATQrZ0tYE17gUPi0MAr3VjXx75VqG/KTwDuW
QNbvXvTdAjQVwLYo7itue7Rrq6Nzlz8CgxenIsND2uXCGO1RuNWrZUcPEPH2
ZKTH4MK9QK5OzapPX8wYXrKEjgMkz1wCyiOResrtoP/2pHDawSuQIyR7r8nL
/yBlIf8DPvVo81xm1kwF/3D06FvltmT4DFsIGOvp/z7scHuXTpZLScZa7QwV
OnHvUTCkgNe8wkh+0725XDNtRd7PwkpFDGJtgVO5AU7hFSeZh95+8iCZRHW6
5K7P0I81KvYr0tFFfwhX7Q/qimZt9Enudi3SnRzhmRWGGKS1vfmwdnnBoTMU
nzMZCIvYkGUENkNCo30EhYOY7Z0lMuBaZJ+ImSWbtXVit0gi6/GsDlUY9Ry9
EHQOJg3NS2a2+C3cjitHCaQtp36GozM0+Fk0d5Z3cxH13Me2hEBkdqgjmmy4
mbZXB97tE3JkZuLyB0GGcuc5JogdNtZjD2QW0eD2VIu/K4RAHFMl+D3EHW/f
Npgk/qlYvJasM2leU1dX1WuYhRZZbXHmjG04z7xIBnpZ9FPwWCygV8UJK0/D
xGkIZEy3QZp4PTx1X0viGEGYskiEtrBKWPtQ8GuWJRaLiHYdp9xzj1xUel/5
zDBsxDN3bhG2lAd9swsRUSAHJhQ2KouGyPC9a/jHBk4/0CEzVoTTcl+UjwPV
vW7ZP3p/U3L0pgMstzmiZ58sCM25xSr2jqoI2fSpAWDY8+FN7ROiRiVG9AkS
O2bBI2XI0FkHdw8zNHeBydAneqJYFy2CN5lrawTQkFsLKBzGqIfZjviPk1x8
7yYKM5+XyR4jovjUdNqPs8ws4O8lg4yPuw6sfQQhMYDyh+lUJfzf6czQkGxs
Ku5Ad2507hIQ2zm34ucsStm7pTlYUM+MnGhlbtVeYErWyZTLWX8e4F4VWyrA
Mtf7ZN7kAe0E9zVo5NvyDaYaO0aZTiopn4VaM3MF0GCbNw5kVjhi/QUn8XDm
5z9TiHLPmKq7PiEPnGnczIp9qpN/grVwRO7Ih51Ty/49GkmnKRpWelcyQdtU
yehPbxuV/eFh90hVzhD381+Z7Pi1yZc7fwYHy1Pq7s+Vz7kEEV3cd8CEYGeN
EP+wfMb6nWl8Rwk62atf7T6pqaPVnh03a9udz4UZ53wRYtTvXRpNLOaLUkI6
RkQNuVIkMR1gIWdsrPO8QZJwp7LF5GkuovhPAXV6YpCbwTInXhpcDaelu/sX
pSMPs0EuovUKNpO6O5Dtz3RRzP2AJpHn0BPfs+9aux4XRr2EICh+Z+e1mXBK
Fr5rwQI0xoeZo9n7rKZSk+qpDtsbHStsK/rirBMJHxkgCFASOGr486cbRC6L
eMIYwgHyGUNHuzW4tGPH9OHx1WCp77A7tvW7GQYgv1p5AAUHwo8XpzPDq1Tn
DiCFetXwZ2EpP/xHks+7APH0y1JfQ1aXCkSY/MkA6NBI0gVDe5EEiHSTXG2j
YiXkembr56Le1NfV5kn4jCbST6Q66FhofmysLgFoEqzDUWT1nGZyj39Myne4
w/dH5/IAK3D1dSuiCb7GBfQagL6IqXFtSoQqee0P4lIKVn6JbJi5IuekyEKh
iHolSbMF1biKCWa68ZwnC5oE3N3Xnwy95cwYVlv4LvajcqtkVseT1cJ/w3qD
kCmfKz8lOUeM+X8VvdM9tRMl58MKwnPUVbHOnhuQdxbyHvWzN7Gobvt2iSar
CE8vmum9sBWVk9r2yV+zsWishLxenWFuZ9/4b9BX2qp/N7Q9AeGAjIexuTRE
GB7lhyoETL3Kr7Xg0QwKyYO9bllIgwoSV8YMozTdMkuyUye8THmctjddHkTX
/K1JPiZQ2BM2XXJEnAzG1Zh7KwQ0zt1ghrtX1Q6AdOIPRaS9oedRSnyLTl2C
MQUmhw4MJ1HdSV7UNgcPLmjVRthc3qGan1qJI1Yfmp9rowlrwhLN4HzYem2A
vatG6evVABCA05SbyCvEj4U0jzUJc4+mPyumFNIDyUpv6mqu5YgozC7kpKpV
EId+HdkDhnKnvGWtxswYdNG190VIvK/j8/jNxH2qfUrBcUHLjtI9h0Jvz7MZ
6wzR5fI7CDmnHfc3ocxX0MEfUyQJ+VHCiuP36di3doxiOKyGAKwOTDcvvbTU
fitHWkkSh+9eF1lnPRiHp+gY4SWCw+aIeRJFi6oTWtzF5yGCCqHHwWyjLGTx
zN1FyW/DLY4AQuWx30xHZK3VLv3sjRtCQlBqPGFfa15v4lbinw6n/xLRUwNw
rYcXI9aq4Zp88NmqqkSAMgBPM+vtQuHMrNFlI/fz2OpRAlWLu4T3Imco90vv
yJuj79RwG5X4eS/4ID+nySlUh2xC13V0XNW/77xOiI/2ltNrpx4d5/FZBX8x
2wjyvlKlGpttCnj+CBNkTvArR5D5aT0yQy09CAd72VXtEfKD94aTbfqdINbx
svUt4IHgyFtKyx+RqejIFCCjopr1HA2LveRKal6GT6Q2Shk9twWVfKsZaKky
WdDIHXfw7Lzp+MI0s9e6ULKUOxenqEiJIZSN12l/HToz71LRVFm8P/LRczGR
bGH07V8p1/VBmvl3NJJKx8VezpyxC9iZ+vw8c+TqH5dfXMQw1TH900bwehsJ
TqM9+5AVZcK2GPRgktY/rIU/DlojE9DzFw6+JLOchUQNY9KJRxSZBXCimRZC
wMwET8GnQCYorFNFRu+3Ee+Dv6fy1KO+EULOcVT1tXGeYgJkzyX0vQW0WHCp
DaSUUiViw78V0qXPuEyN+4yd8ukL7nKaVyihgABxDpT+8pNEw41y2h1sxhVX
g6AwoA2qIl+nNyG0cGwzY0U3yNxYpdWWUKzm+H4PTxrx0u642hS4HjGWFV+h
Eu559W9l4GzQtiAWXztYTNwXp+ocTHf5gDSlZ50BDcyPl/KRUKfcYSK2TTfI
KboosJItlXREgzst5YwhDex5+L+S+mx3yGLPXFW2TvQaeFDq9IlydDGY/qaT
M+FsZPI2W22/h3gu+ZPq+b/1cKijrE0j5s+9JZXq3jLsxLNCAf/BWugVPqOV
/vfW8zY0augsxvRhTjZv6nMbs5DfNNZ8ccAv+3gt8mK/mVNUC3twlFjUB3xV
wNE4eHQAFsLsl1XcYxUuDJRAbUchK/mrreFg9twQ82AwMcGdMmZhtc0N2imK
J3soAL59xdiricyf7mZs1HiT7EvOQOPl/m7BYL65Sr96FZpsIEoM+bzId9u1
fiZdPOwzfbUh9LdI/L1HpIF1gaY4MiTHbFLrQk0InOKcxA7N5HUNKa/jU9zz
LigqLACQvwD6iWSNAIpqZJLj0nXmqZsSIxtgn6nIBMfLYAAmnFWEoWg3qhqy
1uSlvA0TqVS5NuyIB89oPfY4YOin7gSjQm0L9CguAMe9avcR85GJoXoRjVbZ
Fhkeyc9aErElKOmYhGbB1Syw7ZGQ3aYbxvSR5hl4vu1Pts9+t/kjElgBzszz
W0x1/iztvcd2Pho//lTan3QZ2ZEA5I+G7LgYUWtS1ZfEIoC4r61jTOhJ/jWO
vhlxU8IQWWyxTPJeoHkbE2qxi0HFCN6uXmL0UMp0sW61NbIpkfGuitQ1EYel
RBwiBYTdMy4xFSpmL8AtT2nmRbNXHbP1Cnvh2VvxoA41krj0hhzC2mfvYXCt
sfFvQoAz72tqUvWT1Q14FiD+1l58jnEdFKuxLvod8lnSBClXrlWMvasFfxua
j8YHT2eS+CUhJMTZHdF62AKdwZ0+gU7xD1ZYzHkMs3FHMuMYCrLenYQe23v2
vHCbLRhA0myD73iVq9bPTZbqL5ArHa7gRgo9SNqhpURVZ9gARBVMaZaOMhHq
p2sqp5pRhGSJCizju6W9mLzZK9vZjVv6OgiuoaIfw4OIn0dskp0HjiyH76xI
bTLkG0DnEjtUBx79lTQ7G9zPZZFVcWt9CIVJruTZOXf4tD3uUjMEbCaCMGkt
ZbN57duv1GZTUOsG50x3U5hUaQ6PzNoZBoT7CKxH/RMuOXgGdWgEu1oXVbdx
q/L1AhwjPQfJS8MUs45vqwcm5mpNKIgUShjD7N8ioH2CfGK631WrZi1bnD5B
fhji7xzKKfKfE8imKcwQhIpMegFdec+zGNPOnXrsCzNLMtve34Y7mZ+BbMHn
iP/17DLvaMNAyQrx3Wvoq6vvvatu9K7N+GdvJW8V4vLyc1/T2BexdVp4R63o
y3FT86sESaFP5tiW6w0yo6sSJrxpwUOPo1nFIaNMWdtzRk0a/bRKpk9GbJfS
6mm7j16OH8EBjlZ0uiJafHjUWn9XWIHz1WcLSLkWgy1pBEYOii2fcv7/Modk
nWBL7OwnSKFlcw64fEr9qAf09aM4QVrgG/LCzYoAf+dDK8mk34ltzzHteZkB
AhtYYODIbhn90z830gkjY8J8IOm68bWNpw/X1oHO9sabN4snqs8eBo13XaUw
yPIL/rHGOLbDxyWEXsmg6Xf5QE3MgmORmW9HLx74fymiuWWDfPjzqO5AMtsn
xCISp37LLRh3VagwQPuIAuRRAqkRN8BBUeRhxNO5u5+VI/J5e7wJcTNGhYZh
3AgW4RUivJw5vl86CVR57Ad71pwZq9IvakotxTAgtlN1fwknFA5Yqj1btr6U
OP+gldks4P4KyuhtagvH2qAqtNH5oCIAJg5HBqOxLT51jZfaeQxjm36HXwGt
tIQ+FHMwfTrotMiCUTm8h9nw2wnHmfD9/9uHnNkmw1ul9tqjfRIO+oLDMNJp
dH1MXNXtTMaVbOSrCOUsl+gVlT3BVH4gW2VInT9rfGSP/Z6QbaFvh4OT0v8H
QzNb7KhzFnl9skDMiKpo4Rq4602YYoFsQFJlPBXp/EzeSKdVmsUlzZbDPwZQ
GkIVQGHBSie9P09tSZBG9XAU7sESj1yyLO1ZhoVyVqn8BBwUfZTXDJ1dcwEi
zxZYCTUSqwgEvmYBcexB/RvEJMvnB7Bf82PktbynB8HlXnrcbM3UXcNuK+ia
ZafsyB/X4yIif+RNwHqHzV9vbt9b/4MH8xuVK7V2Cpa1ieofKFpZxhHUPENj
tQfNlD7C8rG3KxDrkWxEiY66cRrfNRPxzTxQkAl0hAecZ8oIX1rN0+c1p44u
W1X1n3Ur5l3rXiXu9YKP/ZsI9NpgnDBcKW+2Wk01qR7x8cvjwf9gXwGAQDYh
+lJrmdsf0xgnnIHdqS9ZKasnAY5N0ZmvjnqGXzCOrwku0+xDhYUVAvRS7v1V
j1vDv9x8Uw2HtB4mUmXjAKi4bzDdb0xeumyIyLxYhfqr3B5CFNMtZB9oL105
B+/faTQVrX1WQEcP3hYnmxFcHYRPvSZc8vzqmSahdDRg41yzaZlMTmIuL1je
Xr1V0w5trdkuG8xQ9DVmY8/KkSIsWOdp0I8r+OcGxYlVMwNmiWu7hvLyn7Z/
RTthrjPQF/3X8kBnvaXqovFc2UjTd1X9ZUMBzh/WW7bXQekRtaWIiBOuDPUe
aXKRD7gU2SUfGgge5gL2HCok3HKH7wNyXi8XPvQl+Hzo1SaLZHedzWUzZ1Qt
aljhJzmDImxwkptOxKelShBxIwDx2AXrA1WVfS43y5F2vL9FGp/K9GrRVV4k
1AfUDxeg59eigIJvPcgMrztiKfy5gbyKqjwCT6Li9Uw8rTrjyCRBI3JIlrkk
Tu+ABV+oDS5wpp8Kb3YlKaHtz/bofW4/ddypiHoWAdzVjNDpStxLPfWVTedM
zAWUvXhnZ85ehf5qGo/3YO/Zl56vgFcyVh12JOZSrGwvW1VRuozDd4rAjnxj
mmt89Ausz1GmKYEXj6GzJdqk9BFD02indntLpPMm7+RoZ0EwByte5dOpXyse
eP1PC4nArNUV06AkHknOcfQoyC0S53vAbd3x8PngP7a6e3thI+hGRvzxj4uR
wtp6nTOkuwCFfJIkS1hNchFlxedPCml/EnXxLmj3eh1oYdreh/HuFdJWfNkQ
lhiauzRI6Dfl2HUm8o8S2jUGxPq50ZayUm4hE/QCOvsZkRlQzLrnmJ8GcqT3
3kH/DmZRgUdoMJB6rZhu/BJVVNeapQtNogN2e7MI6QUb9IgR/lxknSEXW6YO
XUXj3t84PDiyL8pvLzqiiT8+eganBSwaK6MnJHCN2Y3nGfXeZwbxgO2snJPi
fMTKHjk3jREaqk7cMhOp3vIq8BrDNJETBb3FmHvwSzDszua2qHdHskm6BoED
3E/XWg9CUfGAVAJ85+ibPvBjBcr7/gFRUlrr0nho7pDTFK2yaHOVzCWVwgrw
ztI4U+w6gdHFXXP+g6X+Ed/XR7AG2MlzoKpyRkKYm17hrHNy/Np+AeDWlzwu
Hho+1itBFHssPlycr0MRcQugunFRUkZESvrXiJWH1+4kXA3GvOW8RTDbNA0e
+aQH24MFtY7b5lq7ULUMQ+EU7AksyIOMYcZRmSiZCyGmMt897yisBFqqhNPh
uRQ7grDqLjb0fTsqOSz01e64mbzNej3wBBDM2G7h3MY1XtpmKHI/ZqXpg/Oy
3nBs0RhmqMLgcvOmVZDYESgdLwYyjIZj0HDocJT7MpxnF5XdRA1wuktEV64f
V4uahRFJAIv8enFOgkn063iMMykE6TZaCmDE8LrsSfliBjHplDveh8Q5/E1y
+YIyiu8VQ2g27Y4IPhM+Ysb4Cg/uS+2PPtvuuu01V8RT0BUumlDp+8AdIS4a
cqonZ7Q1PG4qJHxcenbfPfwxloc7IWVDSiKH9AmBC9hCIYf9p5DvGI4HaWbg
8o66NHfpBe+imy8H62PHE+Xk1CEg0c6LxNRE3Dfkog0rP7/4lFJGyQkPekPz
D7VuJaygB2TyYTS96Q1Apw1Lu2sh5oH5oB3RsDancKJcRBQnMTp2ZlCpAwId
a3J2yTJHeAJu0nQtxWKcwwDYuJiRd91F7yDXDeuUWVUlrbvHukvLNBANtvui
9tAjKWimhpQv6gqYmnhwagZ7KfHU5gNikiGdQefUiD4K8gkNIkH/f7XUSHkZ
jCOmbetIMg9hIRAC3GpaSGsWTZh5kyEWuaJ/YLkmamutbQtcyl7DdjDJQEMh
mbSdfXUvRpUjQUe5qVkYgRtiSmT4qxeq8oeI0mTUOGrwNzLPC8hMn7ntRPNh
6za/nG/I5zfm3Uyu7v8NSyERcMt15t1HoGRqdeWUAFzQewhRTj2+kgzCbWxP
9F8yjlmt7BvkNPDmatZk7vPWQ57EFZ45OVL+0Dixhehgc5l0mSeT9f6IAJPV
T6/gCU34L6SOoAU7rGG6gx4alVzNyhRi6kxY5lAIsDvpjRwxeOBBXxdNHcZt
pZ0iu2If9ww50xKKXOjcr0l77786w2wyAIsamH9QfKtAPlUl6S5zlpFSBSij
vce4kRGiWIENfjN239oF0uVf6l9piTG9rqwS+mI0gd9DMrLxQQCTeeqdtz5s
aVCtuuHtvZVTd6bhEZLePVLUNAwt0Itf4tKnl8WPfSyh15VEwGxncrLEapUt
QuyBOx09nxTuPd//Hqd429WoGHMzKoA1Y2oL1Z6B5dYjydvlnvaBZqorOVfJ
ovhs7rKqwWxCvgOn+tyNokizahXqICb3sMpD+pU2IuxMaOIFLReym33zSfaw
PkGvTaJtqqKKBTipuaTxN1H495oyOOUFQcjmjB95oSdbTNgLlCPFMWFf39nc
2j8VoMS3mXDwe6akhrnGVW29l0Y3FSmdfJgA5M/aUpIPgQW0Ap8vYVJWWGJZ
VORXZtXo0ZdJiJGjvuhqH3AhQP/nAR0BauN+Ug33FyqLUMZB0cRSaIMexcQd
iEblmPJlqbld1pwJ0ajjb4hbmn+fvAASMhzwaK3nY24XhjLcDiXYxtnCeeOA
a1s6eyMl3/nODWrlWm1kJ7fYj0OxBeFDP/TLzTnU9WIw8PCCQJFWzFMxAyXL
aIGwxDWBv7fQJ8I4lZx0yLFIrfx8VeVTkrxiuWlikH84Y/4mRD3CJkH/V0n+
4GOwN6oQuz/fAfdt5d4ZOKtKh9y9kyqCIkWsLiJEQUOt2ZshJ+sEM63+zRz+
0wr0NRH1dYJxkd9oORQJUq+uTIbjcB3ZXHm9wJ+0G6Sqqd9e5TY/6YvykMUZ
d6D2TgbBfvSNzvkX299NSbuAprqazAjmEShxI+aBqsO8qgsvuLVcG6pYRKk2
2vEGi/LlMg0oiDWreDlpKrYdPe3xyRiJ+9qGi01YVYmnOh38R487nDp+v0QO
NnIHMb8UFzd0jmEKXXVZHYG7o/BbCj6Nme52HpRsym1SZ4Rq/lkc2uiv6qZX
r67rXl55stv0olsRr+nBio289/ZImVekIhfzaEhhmHU+ZDMSJRktd1iC+ZK0
B4p4Gi9nEHaxcDYE14jPXO4jx7JhHF61PWrQOC2XHKqRQukMUJUWCByc4KyW
uEM0U2JppfvpWBQU0eGsgz5aOEYe2SCA9dXPtnUFDVg+rkXysV4lA8DPJQNE
EpBmD8aNe13KIeCrXkQ4v2iHeqQRmrZ/W/HHJRvvkALJlg5NfHFgwXcNtCm7
j1vCL/a1KOjB1yzeEyLMbS0mi3KpjkcJGdEG9nuGrc4E83ofmf1/vVvRx+D6
u2Q0gm2WrYLVxJtVcGxddrKeAAWE3fNgg9kzJY8OeFLdT6X+AEQORS9ZhR85
1uggIE4dR7itaDW+wLfITk2H6xbyDmHWMkSZGjRBfMGm2nzus55MWzCYvRzw
Qholzw/kxPBGel2Tp/KQO7tmFDp7DXBioA+gonLNclkd76IIxMI+o5KW5yqe
w6xvAJkx3UCVZtGKDSRzvHvV5SaFqRgVnRLoQq0UjuDPTAyt89JGLN9gRmc/
FV/VqKtIotE/prlASj0MZpZPJ2WiFqMGN17LEF0GuauxhmgF8MhOdAdgLdZM
jjmveFYgYTB0MMSyb421zl9LVQhDo1/CDVsGkXLG/mVLNmCPxGuQa72M+eaa
eKhx34s4W4D4PVKzOnMS+A87j6gvvf5/j+ed053Nb50nWzs6qpDneIQ5+DQk
vM8mkZenCbesfl4SEFaEOEZWV2d1d9keJC1ifsKg+VzHLXyviWima11Y7Hhg
41c/OQsYnHo7uL9/sPzGQ/tlKI0D8GEtJpyM2lo960LgQW9TBBZ1mX1UfzKH
P1EVzPI1/+d6hD3+I9nSBYmd6pbA932bHL5bj002fuPO6JprjMmSz4wJQeo5
nLNKBTt2OtC3sOev4jCAmQAn0ZZSsAYSP0ss4ZhQVnMYkFLxb3JlgHFaC2K0
CA/oL9ECequVqrWGb+q6U4/v62h9Ezkk7lhGCvUOospJR9n2v/H6Ix90ZAGp
gS12KcB63Lz58FYUikJU71xIQURVQ2Gb2oZ/wvDmSHVNl7wI/1jcStIDJssp
zkxNXQquKj2vpsycQyemtyd5MS8tq9JWhqXwFvlDrRelQRv7/7o5jdHdd87E
KNxyNjwZ1c11dSqSc/Lqumj431EA0s0DbGTiNL3ImftJ62DI2qK665rrEidy
NAVRziuFvfchMsoa5SXGE8uCv+ruEQSndEeVYnPysl3YCq5DzynOmQen0+cV
Nw1VESZ4na84exAY/QD60J3/u36Kytaczm13YtmfX9IdVP396dciWMnIXSco
2BwV3WHLSO4js41GNH1xjmoUEAoClgfH5HU7cL3/bEL3WrKIgKX4TbvhxxPX
Ofi1f2xO2HxejisojNrNHPo3wZJoDpOW/YHR7ujPEBbXgZ21QKnru1zayc8S
aZGnopYu+CPUOGSUfQG+14lN0RR4AJutkNzTDW5ia71TwI7D5/mNvGF89skL
k9i88GUa6ig77OxATzWSMlL8zhCzFx/5yodd7/twJBsVN9sQsQCkOj7SHLAL
ZD1YQWuZzxZ1dcCwunQCBlIvpMoShpFMZBa7djMBEPZcBGLMSxdDhQTpd+xs
uypl6X7BZF2un3NiQ2Tf5NayxgrvkmoUsr/IZLRm5eYJS1nwtdNW2Vjlf4Nx
eNexlCyJ2CV4KA2XgvrAqnuo0Hv0rw+lJTkNSE5p/nnGvZmi3l7YB9pBZ2CA
SYjyQtW4xvS0MyS0V51ofHzyRcYKASxwrljm9lL02wmqy7T+MNEv0bs9AKx1
W++R+Ls3nfozx8cO4ijo6OOn/9I5cXi3I8MhTUO54203fxIT5+r/IAljr4MR
CkWEqc71gGR73tezGdJ8blTOO8JUcnI3UT1H1FBKXnceqy4VGeqfOrWHDZIF
BEYHlYMQrnubft/gvm16yfq8Qj361ng0J4ezidbxnTsWhXUDJDpHdbSNpwAQ
yGykoqO8YodfymXp7uRXSXfvsECmP2kY9KUj+T2cRGVlaHTU0gj3QGR389f8
z24wOzGIdsIq/7HtAHLzkS2tXtnn/piVoIuje90shF8/PybOZHDX6sdmVuyw
5N5idyTP2A3XbRvLJh4wUS7oIB/oCVRQmI07LSywsWieGfCyMDdtl5cVTjCl
OnABwiCy4XmwTWpEh2VtH6sQb9D5BUb7ByI6w9dBf0HPf7UcJxmuSf66eeN5
4C8fVi4HI/z7t2uUner8s81BY/wq4SB/hclcbCnI8aw6b7U7qriM1PJfNF0+
frhH3wXETSDYkyUK6BMKdpKdIMtG8aaQFRuexEFPnuI8N1lcE1c1N5YnuUhk
qLnHdYv7C+Bz3q84rKxPPjKlAxLhVgU0+K8cXG5nRzBLO+HM1g8tmgLvwlOq
OHxWySmMKedo94XBX52PvA764BOl7QWiQBd+zWmg/JqJZnwwwpUMW1MPA4nV
gwnE29YgnUq7v9Fa2oJC2PyrI7yLpp9GsUsBCFe9TDOkHlkxH8joAOYrcYSx
v2OT8sPXi3tgdVG3IttyeAV/cGoo0IrrkLgESg4TzypWmajYZT51fK4QXPaF
qTrfXBbAbxLRQNIm35iUyAyOHVklfHGuMN3CdVPsYJ9JypXwLkQwp+W+stPt
lqpLJT+iHxddqdBKU/0NtuVgrf0+kBy6KbKSJhH3HQwlxxv6AuZHWDpP4+8R
GRMDbtediE2IeE482iZHUIc1mq5RR+rlxxjCWMKcZGYrWMQCQSq7+4JoEEMh
rTMUJI5U5r2Ei/KP9PXKtM98srLbo1tPOKGyMh/BshYQkdMmnMcIDYkBkvR3
PUmabMRtptfVnUm5gUBp7ml3BHe0eHS2BBFaVGU29KRkF3fstBcnIk2k1LIm
oHZZLXAvwpbXhIUtonbWeNt/PNZztzdO/uSlJBZlfHgmFvdl4SHm/aC79mCL
PxsUPZA0nB9ffGqi7ioUwj+j9Zk5CLrJoBandt6NYZGzaSnanGmRHzxc+OBT
+2h2hqrBYFVqbdSMFQ0KIfhhaf5jw1yoHztWZ2WmCU88MGILqx03Hy46D0id
NyMzA6XOq9diVN8PHFZfg8LGNk9o/vKBjXGlnJR9KLbkwTwWQOfIqMH3lxpb
ce5xyuAx/bJpbUroRRzPU4OzNLTEvPV5OATAiQwXdZ6XYqQgh/vstFEXeNdF
3RKpol3BimyFx5CBj+RVFSEXAVFjNO8CjhTk9oshDV/dMscVtKL2W0NXiELW
/yHxlsVv0OAvybBjlhw0/+OrYU/MqfEwQmTdsQvfqb46DQdb4IMy7bo+hDG+
VkA+qU4HBNJJB2X3th4fz3nXEbUXMazkaKggzmJmWCTd/F8tvSmhcCnj9+IS
aNO+1L0osk3vDV/KVd/0jS3OHgsODeX8iIHKr+uf41c7mMGkZsWOpJ8tgNij
xcG77wpYf5g2z+/lNui68SIy0dMjgk0cCbe3uIdqCqeamsGkzzwncy22cXEO
+10yHhRyAMU8SybDCFsFLW/ELm1fA0u1UyQZ5YJ8ZaB+LgFBznhPjjjCg/k2
zyQDGx18f2+g5BbGaEi2G73OYNAPGkYKDwxuv1COXbPrgDLqs4O00WAlKUEV
Igyh29RSKGxp/pQhx9CWmJwt307Rids53hKhOuptlDZomB1O/p61iHQMLeV3
Kg2XZTyiBuqtYZxmKI7+LyGLvJ2dIufeaPsH2hC99vJz8mwkjNy75OgT1gwP
VQNqmAGC5DfDuaSTgV0d0IcHImLRhhr/JYDf27fsNUAPxrWppNb3opxcg2dV
Rl25djloV4vg1uDVAt9b0AhObV4W6r42yqYYyH/H5p5GGaErZCeu3LwUgVwO
x89FYybNYN71IXa0QJ8Mvoccpv7NQ06xNDgkaEeyxqBRQFn5TaUtW+jprF/+
UbThZ/o0AR4sV30Awldt0bhhAPWDyn1LlJJZ+8dOb1OsmQUvJxoRv8/pZMUy
/URh36QzKmXP/d6h6F1UtBSxave/x/5+qy7yVFHIuaAGunP8BcPDxgRXXzus
NGuxa6ADiK+ojXvCgB9YauaTJlXlaBzH4R/hntSsB/MqvjWUMRP0L1Y7ldS2
oRZre6aCHyEKeKTZdtWPFqoMLVy92Hz0Zjx5gXV2pwDnNjOoo/rOKYhjtskn
zDWjCriJTNEodMv4/gCMb5kYfawuc7cAMVNHKt0Q2hrUN8wAKyRp5tNtsFkj
Df8ACxNUiAoNHR6aK7cMdbee1YFLdXQtKoC4epeorKUaneBxdlL1t2U2ZcCj
/VmxfHR4sfHbtOF1oODko/d2e2sqx4ip5qu20z7FlcW7SSABIacx2M7VVxQp
js4pnAdV5ZDv7/QOR7uAu99bqGGzqOA0k8saJopxYffFo0Ii1mvQmgs+QWYY
xuD1AB/gM+Kc6F0oSr5Mwb8rm9X7GlbE5ZY24dixZCxbI/7CmEjnVCBncHhQ
kwtJmR7K+TQGIoZ3RhimHKv9Q8tPCkFLPU3WAmPtgnn2tHnTR7n+TEJrDbiJ
N7SuNzTfixz6ZaoJPTdppj+tkfesCaA/gEVmvgHvIYkkPSvPZTzDTaG2TJsd
McUY33Ry8m9oxdZ+/WRkQfiyB/TAC05D+448xIYO3qspss9OAXt0J20e1FuF
gHZSnGK8V8+wU4FdH3PveINmPDpVxt7Zr+90vkuzpBCM43QS2e16tMokpYgW
EXzJMHiMIOTT5fyOTu6uIA/+ViJEwZ4jy3R+ccH9HBizjGc6jgZkkB+C8qJU
FWgbKRd8CexaVDZqHjphTb56/oCcetGpnulz3Pj0TXJtq0TH9iI0j07aPUUE
cCjx9FdUWHbyZHSU8tZbY8edfXkLZuT2xna59c+wyqTZt/2kk5tFGHHXRFjt
Hu4WtmPO5fgAx5UJA6dFnDJEvGRpR3sEboNX9G+xWNr7V3O9Hqodm/xjhfLZ
rLKLpqa4qEiE6/3rgyjgQV1R2J2UYzg9tb8YX7cFLiRL4iBIofkybdgy3+o2
gl7erjM4Pku1QOXZkG2aZxJYQUiza2X3PypBBOp7O3or4yKyt1KYcvQrrUpi
KThEj/TMh62odfYQVV0EjIQujbC7Y0PFbJk6/RKFgvvUG8ArmLkeOWSaw1MS
dtOOTiBX9LwUSol6M1Z6U/d7wv022QFaoWy6kST5jSRug6UhINt/frcke+ca
NubitzVpH/q0AhCH0ilETx44XVregGK0+lCFSFCf1YM/m43cFOenKK/smQHc
8+myzxFdnXiD9BAGj9b7U238w7jaMdD2Yr2/BoDyQDVvfhD/kB3HywQ+7bi/
g3kemYpJdpAccQBC9V97ZX8D+w0wUUdr9yEphQdrxf+8pC9aSkQozAahyeof
SZuplGj7s+0vra2wqjd7hByDhlN1EN2w/R2I2wMGatByUft6AcWfqA27M4ZT
wE2yMCgS5K5FhpwSdxXWuHT1kv/Xs0xCBZqsfSKGykB/eB5ER0tqE7mJjBcz
2wRbvyge1zvg+32etKRX79kqd4Aa1AyARLzL+e3OiNJIUG7IrZsUFg6lzFLF
/gELlbHz3jAVwLUqocIb7dJxpS6vvMJxDuo7FuTT1KA54SAg7DK0vDKdLuYP
6XBC8UghiNQow9H/ph0cbQD8yrTVaMcGoIW4QuGWcShXmuxCFdcgaV4X/kt5
ipfzri9Cdlzjmluq6rSHsX409Ee53hwfA/6yLjwnIrXUdLrWnG4P806xvqLi
z8fRXAPSh7lI+OtEFb/Mi/uqBm5PzNUXSKngTxSmZUObvBfmZNt32Iwb7h7b
jRoJjTT1g9XXgzMW/RKN/twk2C3mt7j3AJWykFhMvpz7yK4e5R0/NarnaoCf
FQkfLYCbKbEoQ6BE3le8rT1MXadn4OU6DYmgH2KW8ZSRfHPx9Gfi143ejlnU
zBu46f4WGYIU2iJNx8fPoj0a17gqT9Umq3LyAbw4Zv4H5xBRMBklFSePUuat
9nRU5l6lq0Vux+1T6x9J2P9vMVn8cg3ZFavV8fHZ8D/0wTls+QIJx3imNHdo
M9j/2DE8lxyLKkFZGCBa+Rh7phO6YnRkhJq1VQPEiCJ2lh+//UY3hqczJwZV
eoI2/u1hXHjeiREXI3Wn4RvO3N3KKVf7u9fxVCmgyJ0OBTGInMkMArv0TRJ7
A4jbYBKTeO9rS+f9UBBSnwns0MOwFonGFVBcS7j1+3QTh0Ztz+z5dFkJtyS5
oheXw4yoD12auO0FGqhNnW4hv+H+HYVYxgNwqpXWXBlkrHfe15Bue6WKgLQH
CVJzPn8KP9qWb/DgL6LZsL8ceyuPGQ7KoNvTNSleza4fT+c1i/pefqeSQxHx
eSL+kNtO+kpvYRSN/D2AW9cpWh+/s6OLKqtM6AnDr1BFjqtNRiCy0spd9I/8
3X6l8IJ71+CxL7WZYGQLsR5XiUoHWef0EiSxKqI2DCxV9xyoG3G6Ntg3QsGd
nQCfG0A3/m0cxl3wXh8q1jkeq1emPNtLRmvOm00xfoGAPAar22HfM1eJxSha
JofABz0uO0Q37bynrA36S98F9xAwpXmzN48FJEXux9Hqz0m4RdJNOOXuSrb9
bcHZDPml4yaqDvpUPFcQZKfAwTd7SADy6U+b690GjtC+fY05ddDLmopDpfgI
kLJxRFnN4VW/MRTpWplbk3ApD1Ih4OXae1bO9s6wjORIBpzdSILkParOZqL7
wfO3ESUA25qA6VHAKFGwwkjUqAVbeK4asjK56+33SM3wmHVjaPC5iGLnDN0+
EqBwq3ZEeKe5Ye5bMcIbvadgNQXETmCpdKmQIKFsI2zEYv1SYccJAN2dWHao
4h1clESpXe2/DVXOkfzQZp0dTyTRkkwiw3OWbufI9BtSUMilAeLTKEbVpj4b
o8tLOyo464EPKuVN46wrVENhhvVdtm+SlxcRGCuhwJE136v44kXmktIZdHAv
2yYbTNonDsnROj+OhQf8G70PQ9Qs8hOZBr5A9WXkPMwlx8EAQW/jK8fEIxVy
U5EVTPTmh6GE6Dje+RdcIznqUqKHiF7wRdM5/DueBf0t0zWhasSlvB0Je06g
SzJ5q6fWLzSvmvF2cRrtuyXI79ePa0zPsA36PQBlwQ7OvTO73NvR6qmzscr8
yRdkcQVYaBk7LQ+6NAuYmk6mu+j3t5w1vBPQFj8hEbzYfEUBFwrw33RqgOqT
+S1s2bl15/1Nc95P9a5jkgmwGsBPZ9ekEhshaT7iHqhIii9NF63okmW8kLi6
xx3dlAVFB1o1dloAtGARVriDmbyQald316IcFgfE8cI5twWFcTGh89TRA/xQ
jINyByNHG7sYJOYFMIhvOMYkFRxdrGOB721KOgWRjpQAlR3Xr3urU2t+sV2l
oy0KsdYyZQQ5ctaAWLMQbgPIzIFCn7voXj0ppgk62HL1MvV66uztID8pV246
PwYVhA4nt0vL0Jv7BCiXMGOms8cMqKEn56YOYyV4nFY28rRuwgXF0U8No5Xu
iBLXxUwYC5s905FeBT+9I+2OyAOsk4Uw/JAMpBlnnMn9WIOSD7dEYHXGnRmU
F4hq8QqEADFGjBmzs25AXJ9qewrwsSLfxhGy2VrqJarcMqkaky+B0EmCbIhM
DZmrXZ3+nAChC0x8D7HvdSr79UT0CuD8yuRS8rrx7PCcfTNy0CAtG9JrZZXb
ayDTTbckTOZ61nSmev3xErxdymWCeq/EAnyavJAKZePgacDsCtsA5b1pbClN
nr5gnNJexVXdta/xrh4QpkEmy2rVotDRkwNYVht5NtLLnHDF33VwFcbOWZLJ
fCFes9/GrHZG2xV9MV1VYJKup6wJG1/bvNFGFKxSt4HQiQLWLI+NWQh+6tJE
M2i8+11xivPHVCmyPmdWSeW/IFrT9soaQ3LStY+8LHk2puihdu9JuINzgXa0
jLmCUEaaCrLhvJQeajkJnNuV2paracJr1yN736jec9cMm/QW6u0mSXZOY66+
rHDSIpVyJQOvANEHb4upT1dYsNNbCfdw5Kd28cH8jcNyLrw6S7BRSNlk9Bti
mw3nAxDLaXdDRT2cUpASfCxpinZ/Qwci+4GG0ACDCiEJkYp+bb7z5ytlhFQK
H10Jt93VBY3nUe5WwmYgb3n1O4BIn/roYH5m+lXeBrHHAFwmq2dW1EPq5xDF
LWelVdN32IQy/lgR234OvaLcr8Gp/QCEZq5qn68/jtnBTIuAAYUvGx+TFkSh
sRXqW7dXIHEntU8yowxxqmwPOvGmBJfb45MBYPBQuADpqEAElke+tLQdO1bL
hlcxAyQ/YwrBu96ufb/dhu7gE3+krIOzipQP4eXROcNF1MpgSgrWnLKt5gLJ
iEdfT7BDwhLJpfFI7RrTQogjMhV+Iolo2MIG4ftyO6WJ6Rbk77ZU8QhLyjeH
EP1cxB16BMmjARBmI8TP6MCFB9K0F8WTVa1lQWwZszGpXj081PT2mbuONF3s
HjPJqgmG0mfRpLa4TofeYdIBMMdXD3cjxa+BEtxis912QC05NxJsDz3ZKiXy
xE9bilfebkfHV5wXpe8YbPbW8rGS/04maAE/rs8nlxLah2V+AGMVBqlxYYSx
eg7SnjpCnnMSHvisatE3xAmTlp/d8RLDiErX3NY8lE4VVouYqQHeRPT5bbpe
5sHgJQuWbMlqBwY5t2se//DUXWsTOXZTjCv8FjNfSYdxvE6QndZCZpeTnuLV
kWoV1HDmuUNRg7vkHyDawSc1es4lbPsd/TyBBt+c9m7TH0vRjoRHAY1a8V1E
LhFuH59LGioU6wUyCv2UJBdxvNyGhMm3sM3ICrafug/XJlsNUGFC/lfuYvEx
uXoh54Ol8S8ADr+076yTMipfcaba20pQSmbeWKEfgyH7MBg9dpRXRfOc6hdP
TtKX+BXjfPdQB4daRKFlXO+EeehGpIlH1ycqhYypDUl3tvcVbT5wct0pk7Mx
+NiOnl545SUTzrhBJFbFh5i0j9d3FvlTB9No2GVO1p9DY8NAJqPw/C2h/5/w
YLuL55frq93p3RKAsdKOrfu01+nDp3nQ4kUGEr4yEkDTFTevKlkj0+UwhNzw
shjpEairrinb/6rzh5zGbRjMa0gZG2y/9f1lOcbAxC1mhhSNsMkmEOv9Y0lC
htHgDHVjSsRl1OEQ0a1ifNyjU6QsEPSQXvsHCxteoU+R/OADP2brrYuODBrJ
bjggdka39fpUQUrInOaUjmdyHr48JD23JxfQR3V9oZZholdzVTtEGutlPnPd
gL3Fothfxc2VColaI+4Lqzhvfg+NLOXkKi0dSjaVMREJsqA=

`pragma protect end_protected
