// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
T6DfxHC/ynOS65fZbEb+AugtAhcFZ+rNq9RQFBpriKaDtHTpbSF0jfBamXUv
wWGcu3YBIVdqRyL8Z72t7yt8ghWZwlo9LrA1S17KyhnXwgTjwfg0eS1LI24V
P5h4vCANhcheIyvTJAMsef0KrpO6lekJ56CwpEJHf9YelD5cvVC9Hck+cXwl
j5FBqrvvbfDu5NIjJ7vg23iYUZDl3Xqsv/JbtAdG7PuPSa9scWvVhNUVHM6b
jffCBBBmlBKdRSPXvFbZZ3ffXtUtheBPSGjwClgSO4imxfGvR+O+6v9F61lH
PPoHmr+8rlJEdXoAgJPX4viUdZuuhp47B09EK8kQ0A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WNOioioA46o0iMHHSHcMMjZ1I8ldukvBcKEAVs46RL11/LjRMlwGBmjXgnaG
RMBqQPXvPyZuBZqjP/iUT3bF25FMt2oF95EdvF9VfZ/eHN+z+aKlQjup9raf
xomNLeYBpW/LrCeeM2Lu9Mya5KYkEFXCpumF3K5Cb771CUhllN0EQPUN2Tmh
EBfqApkaK7Cv6VhgWIqkP5/bXnXsSe4Y8x7NRdVVVRtCeX98mzetb/mLEKB3
Xai2l9plvVh8q+bVjBhxbKCURxSWHyA528RTYba2rLgbcJ3960C8YkQfwnM1
503zGfiguXzMn8jSEDpjS4gB1Zc2RZKM8YmRocDKSw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
POAErXSP/yEEDna8V3ORiIN5EfZGfCP2q+RoAGmxtGLYApagZgl6VyRejIyD
JkjODzCWISKFHAEzIqEWLBhMkIhMwKfieJ/QEoKT7/ogX6234dK65XsYy7vM
x1ZqsUmx4neJsAjpx00dQI/uSppVzfoWtVwLMzkpmIDRTIaPvX0nx/M059/8
S0skoVOsylmaDbsUkQAzD4n3MlJ52WdaI/kLQ584QYkgYjnoGcHqHa/N908w
FkUy/krSXppSsd+D2AEiPp277zjOOkrfFrCHabyEHPpwAdNZ7mQs/adJ2m8P
x/8cxMt0Ou1vGLsTA2ZmqLxXZksnxBqwl3Kkw644aQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QXHCbWO7WHxNOZh0XLZH7pOqMUpKU29AOQH79p2LwUZXQHpWQRLGB+YTqppL
e9ej5WbDQj8vjw1Vn3OtpLykVaDa0DX4rlMP2TnvWtuTS93zTFtuPkzWmliD
51XydqNWcrXDv68V5MkFmkzQ7KKA3Qxr3SiZslm7sD7+mGXXp58=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
S0JoHK6APL9hmdbvoTEGCacxLKaJTnYhDb5+leP3nUD9xsioj5cqcNGIahBz
T2aqFhNZF2mfEw7RXu1uEipjYjvXqQ3nxhbqrRel0REFD6Qz677lHUwsy/Ci
Zc1XWzaYfzkezqH9lVOWhQEv6oGeGPMqIXzLt9DME6Jbwgw+MwENh/0v+ULs
7EO3yOmCUn/ZM2G8FbU2WdE7wg5tBsyMQqVX3arx6lcEzZ1mA3Ia7y3uGoT/
wo2w15B1bFgVhSBDIrW9S2SIDYgi+bH2mTqzDPwbIuZnDFJIWDRZHzmWzqAw
AWRWVYBG4InYmPYIuCxVR/suhdicKRnoeqCzY/WH6wBMH/MmsgwwVYf+Uyf2
Yu7hPDrtX8BNu0/wMCFpYlyJxLOWhgDiJpbqhjj1UrVi6fUXUQ9JqDOFK6QZ
mjrVXvh3nnilZ/3HrugL5wJTGPfYy53t21VXMGlNv9b+DCDhO9ipSHb5bS24
ArfrkijJjyuoLzX+rOrop2IkfDiySisk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TsVkvcrzpZ70/1eYaQdPUDIsmlnR7CDChidpiZQXst59dirls+xoDMaXB47i
EReBFaqW6XCz6IiIm6T8pdE5v2/RLDkMpvotR/cYUj0rlNkHmzkk03GTUtXf
nqUNLdDXZXDYItnjD0KsNcvj7W5lf075ImRbxCHLq0KI1yjn9oQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ezSdtA1KcejPxepF+EBVzFaPGtQg+oysRyfFfrpZEJg2MzJk6vxrql8egexe
icRD+p0eIRaQh4bMoVHVlRv0wLsLqDfSA1v/gnAK10qOHy0Mi1vGWjA8Y3DQ
CVftggwjGsZnb4OgEVFvOTal1NM0FU0aYGuRwP8xna2LbCJhppw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1968)
`pragma protect data_block
DU+18iWxq0n/YtjxiJqYoeTU5mKb7220UPnVYzIAcshYtf4lwD5S4iO9YUKX
UojQ7oHSRRjvkyIczc/p2K9pa5yCB/PYcdjdWD8d0M46LL6X1OdxWsE2ekz1
Qe5fDIHORPrsMiF8NbRoI4sZsGloKdpFLycyn9FCAAo+dZSFtdZqXWkXz2eL
2OU2Gn9oFkkeKBZoc630rktw/53AHfNKbworvGSF+3+7iUi18OptiuadkhPh
vRvoulobECSCbwT7GAVhgVffNCjdXAaR6ESuShNWqBmBBI7nl+FfwD8t61TN
bZowy7uPjBicaQHqvNcXON1jSoTOTKc4ugPx+Mn2TmMJFMYSKVe2t2C9lx9q
LnSO/idLf1oqHUlN+8+567luqx7uZx2XfK+vCzc9ril8UKsr41Magxqgg115
/z+GzY1ULm23oXz8R6DDE5NlUJdsaFdipSDloV0YyUbFPvcwem5PnC58y9SP
6nXf5Paz+3NeyqQIOIX39rYOTFQxthllRDWV/oMQaCFOhgvumJ598t/kTL94
11mAuyraxH/+FBQ8HwNJsUSdWZVDmvpqayGyC+0dXxoUkInetiJCHowx5dv/
OHFqRq0viy1qA0qN0FlSBYJyo9NRKzpNRN9eAB3KZxILiIv+GtO+cykqjkNI
Fuy/Gah1Ze9+9W6TFacHcVras2fmiS9grpbtUjUJ9QYg8+eCc6Ux2RRIgWVQ
ISybezZz9DK8YYmOx884YBZSSRDlnRQI6YJ0Yg+X6eXy2+r4jkWoqu4uV314
zJYvk057A3jcdApviAXGZUy2pcPuazeO75T2NyEG1Zi09iKjvUOAE2mRKTHo
jWJWW66Gw2gpPbkgmqWWVRsweZL4gHhe6kaE6BuWBfSSrRPLoM0uXuo5GFEx
rHJwMvJOmVL+0ZWpVotMeWOgoxUBj+NiMZqZ7j70BX0Zw4o6MLTFxsAmyF/r
JYdx0vFSKKfD4rNpaYnf+xf/7bOpby1GKXix816WdjXl6+n784luhNGHzUX/
63bj23yK2HoTJlFBkZmoPE5p88QOFDYGEU/Hrk4EaKMCBsJoY36EJuQKSAU3
FH6WCbsifAN96yxjvYYoJDRxWrY6/CxPuCmsuGQUZDm6/Hze+75v0AXtQAfH
vzN8HpUfGYBDuE2is5ea+1PMAfWIsioaaRgDPxxxHW2jaAUGUIXnpDe3hzxl
7Sa0yj6+5ivNdr7Pd/K6T7AsBPbIKv6TFOdLjrtxpYegebn4xvwB5GZvOD54
CNeFSRZ4/dgMpDCKxa9IJAEsdwXxiYsHOLlSb6FSsrSguZEoJnrPPfHVpkyZ
RvkTCi4v8KsqcXNgI5LfBmTA7kiLey3Du8hPeFlcZ1LdDjYNxoburEM3ci76
siIAS/MOERbtFLcYciJ2Z8XZYxnO8eX5yaI60Bhezm1oP29qqKRNAKsSvdkS
AFtThGIDO6FuHo9EyvK3A6lcVUiPGWPFF7I3gxICbjYKMsKQA3xWbSsCHIE0
ByebbYaGb+b6gK7lo3aLIToyO8VFNLxyFChjOVrgu2GblZiQmAPfI/usvAt4
6QHQijNjS5761RBKiTw0T8gRKPRvZ8Y5QB4ySfTAf1AbuHF7aUV55EJT8igk
tSMq0UhNb11E5Wo18/QyiwPj7pX6ypAPc3vGy56xkMnxrXWU1Y4kEjMLEGYp
uePyhbLrBL/cE1/Kta49XKE19tcW+Jk0OhMbPxfjTuo2vXKqfZG8cPfljpWR
f+Fsw08+kH26vucPst1aF0W19T0JpYmfV4y6bnwQ82ZQpiHB4F71qEzeOZat
0wxE7jeHx1Yl/Z8nR2wBBrc7Cv7LacGOI9ICJ0t9UXV4V+loOJPA1U0Jngyb
a5eAjJoTzIP15xwVamR2BsUK8UZ3zg6FrqJFDiqgE/2b5OAsg2+IK0DTIXQ6
r+AER0bhs2CPuCEYZwxPLaRFYsCJsP/C0XAYZPbQKYKb0iIsTWlNNfO0v4X7
pfaVCTOGLVt3cSFJ6l2Pjcb2dkzKp1SFLFagkrv9svosg1hu54B5PA186i3h
Gd6EHPdQMGOUhAR3/5oq60vFPcdkQdlB8AEobMBJBVV3QQ1Mc+2i0FYg4w0l
fjVsRs0i9mJXvjU3vJlI1DL7ZUEkKIYVLENibHTYAfDBUYbOp4p8vlDtHiIQ
M4MsO9z8FKpHbaQZCiCbg7O/F2YFCQXMzL9xbWqZhjZKNO+CigXgyRLq1Ulg
RMjmVVTJMZcGnz01Js0ZBVmrpShed2VCHwGvl6wY3qsdxwUqacm1ymPFFJ7V
r/LUpXDkyQMTM++w2/zJCOBsgM1ZFvQBhidSAejxGbYUIof+wZwrkx2JLbXY
Kwli5EVu6NHQc1rM8GJ06AvFWs7dQeACL42Ljkp/PfQi1sH4sPeaegb8ZzaE
8IGk2zhVsc38JXYaVc0OmclGj2PRRMsVyjUI8hVrlZhNZO/ibCiASkrKx4fC
V0G7MXUH5vLfcPAcw3uKMi7L4Onvn6OqLrC/bX79v6GUSP2eMcAywpscaPGo
2OOKiqbGj7yJCAtLvDt90+rydU7O3OmArQWxZTs4ylyCCHpl9dj+KrujgPna
G+DJwjKVbdMaoxDq8PwODUg7UPM2h95b9bRU/WDfaFOp

`pragma protect end_protected
