// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
KHX29i/vUSVOJe6t+EXMPP6SrR3Hj/e6DqeKc9y2oP2bdjfj5ioxyt+Qo7kukxGE
+E3Haq2NpY5cFM2mlzwkmPF5XjB6gRXBon9h8yliEBzpQzK1b1C7QbXTOxRatlTN
80HOicKnRbD2l24E5xVCFlAw//JY32RtOqoumA56Az0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 13008 )
`pragma protect data_block
IAnwxo96b+5Pa5v2d4QzL4qcGMrSDswWULMXyYjgZo68J8Fvj1W/wzhqeEsdEMUc
QMCkRBAYEhdsMM0zUmM/bgwpEpII1g3pv4ejlrLoZ6ajA3wZlpHi73/pWVJog7+2
/RZKc9tVoaDLCmfzM1gwP45U0RU/yRLRD2UzSMSM4cK7PgKaz5zQLVab0IDLlLMa
UaJ7hZRp3UqF44Ou63g/TYtGS3n2TPf7alMHRxRc3tSrzOGmAifZT5zQF5cESliY
BGUekDDi6sMXJbp0asWtboAy5spSklqp+30VdK/vy4kpAJ8KVQhP/c2IMR11xA/4
cj7GgWt4/oPTFu0+j4frt2NCiB9Ac8NIQitc61RM014ugNLlv9tIIvpcdZxF12jF
i7+s0nIrkaCDaWZAd1g6nM0XvulZ/o+TmsuXeny2BY3ilEMwW1FG/xexjR0zSL9r
XnHhnyo5GaNnUBTPLgNVxVvFO4l7ld/s4CVJuXG3Ymqar+Cick0cUC/+TZTVwS1Q
8b4vjlSKrkGQX6EcOuWzsihkApvouRqS3XUpCHmKNVt6wpIdiXxn3ijwET7swoH6
Yw5PlEY+PBCH7ybSFJL6QnGUaH5rmfzyYewRv46UPyNsTB85WX8BuKFS/tGyKA83
rXjbgSeTdLbyPZsVZqi1uMqT/DcmeYBKGlw/So4quk+tqDcGToPfXt66EzabLLJ7
x5DJvhf4/y1PRZ+cCly9mPOtS3n1LRVHwSo9pcU3NqHPPMOQDXT8nuDSfzOiX8R5
+j1rPcTe5dKw8BxwqI4KCoEfyZcKkT/l29FbSGkoqqfLGB+2N8W4B4xojRD8eqd7
q1FQ7lFi0pU7mUrxrbhZF5UBNzEctMCKKCdMlS39uReZkuXCWGCZ2sVjmqT5oEIQ
AuqRBYsO5hbnE0TpPnyRrB+5siMTexY8FVzxFSAaWKKO8JWpG+6TWm2AardCnkSQ
iloL2/5lWw+LGh202+Rwrk5ZELODD7lEW7pF4kZ43YreG0ZD+21erAnn8Ev7eZ6o
8q8NOysPkXK/xlVbQdZsipPfrJkqv1ycxTGgknz/Kimo/JY/ja93WP7HaXPI0z8F
zRc1l02LRQ14nda7SxkNs3zzAwBp3qxMMAnG9FZGLjD5FD3H9knliiMlqMAPk2Xe
qVMfXSGj/mBfE37ghiH95uMHFF9qe+4mqBdOcQIFYUoULNBAWXdBn70jeWZDzOzG
L88CypkkiR9OghZrVZ9uVaIkcyb+PCVq24NjyUSHaqt48xN4JSZnpEiOuqNO184T
xFGdbX1WUZbpojqFSbMiKwFqEWjCEC6AK8g8VbWkASTfuswIfiq08DvcPeyfEEz/
b3ANphJGLyaH1TctwxAEKga/OB5dvLg77Z2gO2Q8AVkbOLayDA9bgxzHdzGJtCZd
aWcCZty2KCiGK9mmas85qrZT4z0uMv2ub0SyrnikHwvw2DGflv1hzZbLcMmfBqBE
GwE5lyJwkUyVf0rg9McQnh6pGS6NayiNgyIEVRhEE0bSTE6z7DiZbgTFOAO33qhy
GNUuzOa4PYBV780IBgXFXEAqnfzD5bliE7iXcycIVN+HAb87RVnb9paMaPWCEwxk
UP844vd21LFfj60wXRPJufik7vx1VtW3afnx+V5IVcfWKUbRXR4fVD6DD94aGj90
iQJ2yk8D1osJaGgBtmArd/8JXt5A53hAdhPvTD7rSTYwkP4Z80pVICfKkc9P9v3C
nqusopEzQed3LiFkKu8A/MKQ6dxfzRmh80ehK11s402r+UrSSe7kW7FqC1TQHjyR
edR71vE5sXv9x+xo8eiAEC4NXREP5zCX1f/Pm15Fnqkw7kJpclhXY3hoDeYNpOF/
pwk1ALwpn6HIlTeF676dq3CBl04DoNuOXyClHpV9fthDtRD0l/07zmqbK0xwR4Pv
4aAbZ0PHCEuXNOe8honHOIDDdFTv1SYzie525aZ2qTlWmwMuv4dQ/aQ3RTEZif8M
EizsIKnUntA+gRk6fYuhXPfp4Pus61zj9bm90Eb5ehFbb4PkAh2gpNU4GmZXFR0u
e8M/GUoNhH54XX7Fu99alT2LGn1pTl1W8swhdWtgxdvKfxfabQV1MNyYaVpbdaeW
IHEZzQmRwFZLgiQ1boI+eXPsokwi0/HUQatXB30VAmJV2yuKLhzbTsA1UkIDGhKa
VGbaj0s/JUlPnWRdfARSiSg4DYIeueuBttifp1JVyMenZjCA9LsD1JJiwywV+ECH
JfLwfPF09LPL7fer5XkTdheduZz9tcqgEobOvyAqRllG2m4PznrIW5mE2Ii6LhG8
Vms6lMOSr6GahASuMDC26HSl/0tXrQzsVAb5OsnG3z+RPaKC3/HWY8e9AZSlLnvl
lZOJI1NipEPRQzWwjgVNHKzQojDXUiMZDcKk/Si9IocE7aGJTDtkCGXH/c9RQ2R6
qP3fTDCk9exKGKPnGrTpnzJfibr+uHUsD6PQJctNuI42lmrj3GvXnhgeR2x+xM1X
8DING2MNSHe5Uv1Wd4oV+33Eb5cqsl/7eCavy+VAxUSNMAMURuBbpavMsVxXVA9F
N+zzwAeo5+Pox0BpSAV980DzyRa4Vk5TMoyVMudoYUY5N9C6leQbZd/LJNFNDkWF
6ID4DrMbhwxKzrpXoQgl003zGYOySb8xjbJMKBRXYlD6NADWfrC1nTDyJztEQ1E5
E+q6u5PLXhKI5c8rLTejtS2TzZwu4WptBvSlP0iSeWf1j8PXASPoHPXZ/Ns2ptIx
TMnuIAd3CnQzkLcreWQqi6ssiALM7mHOSQOEmaRYj9A9bbEQDDS6GPKMjfCRKJZC
D9eaOGByZmsDZQlR0xJwMw/d2HhL7L4DTQW2fjJweOHqxistap6EMv4WjYt67eB0
ID8gIp8gIyshbJZvv6rJE9vpo9hyTXzTrsAfzJ0HZnLe8fKVmAHyJHgbUeNLV+Hm
dM9xrYl15xZ9RxhEjGQUQ2u3spzKB589IkYW9D+jytQmYYPE8JNkrxh7FHaZZDVN
h2OKnDfEAR2XTt1rvzkeSYxFYm8o08sqqCWfPe7LB/oweG+uEzKNCEqBQPZEoA30
IzBBrGrUbK7+ukcdBwByNeb8eIitub26mZHqrItb8IG9IpX9BgthDY96iGZbDpbo
0muyxNDtfDDVAIO+lWaLIIRmFuTyD0JXartMmABU3yYfz0PrOZ7c7ILcaRPUcUV8
RI6emN8W1oUToaNfLYQEMkuugIdhgpFpklmGaukb4Li0hT72No4y+cLPoG8bM+Sb
i7hZmkIQPeddTfORJYyAtS2yMgdFnSYDtwnEqGneJHzViu5ISqX997XBE6b3qoxB
FjXS5ZxjhsU8nMrdMPv9IPX5QCM05u4HarKCn4qjCbCpPcguNj8F9GCaaaeZBs3L
af+5qFtTrgsaapl0Psd+63twvwnemnQMUN5SGyrPb+KNPRRPGVXB7R/yNCpeQgcX
vv8yTrNxLkGNqkBCdOZUAOYLBCNHR+HRhufPbkwNz9Sup0ny5gS5SUmGwdtW6OiK
EO0Jw9KffA36w4jr1uwgdridRpeAhm4kWfbOuXRaZO71eOV9AHCDjTd8pEapMpzt
0rt/TKUx1rQ7eKNi2+Pl4zziNVe+EMkkO09oI+UPU0FMw5FMqkUMmgHrKMSuQiDI
+68ExeelZxLIZcLAGBPhGx3ZLrfgrr1Oi0tTzt7mybL7LPcsdfX/dcLqh1MbMKGJ
92sXVIlo2GUQpeGGFn3HhWFEJdbFAUVf72UcjMCNckzXUbzcAjDzlcDonCv0dz7V
WYLzWrSYBy1eBBvNn+PMJYPrLh1vHmsbV0xDuf1M75OgNNLWBowUMqOKHB1p49Zy
SlbsRCzWj7JnU/Yrur+tek7KOVPIfMpo8oYHZBWAajk1xr8XcJjg1KGR6Bk+ETpU
5L9BbovdjaF/os5mMnYmUSUn55nlFa2Q29nSbnTG3xkaV00/m60C8ebU6JvU14Wk
IVX8TXLGduM73mjdBOpjbLlQNGdyBhe/v1YfYU77G+jyEes37JGtDthsAZi/XtL0
r1X3fLfbOQmUnDOS/lc+GyN3etS+TnFRaut+52FXUqL8DUtGzLRYk/stawfzZfMW
AlYsY5CV30IkSTZM2R758WqTGzXoCz2uVZSemPvBO+HmNMIQpC5WOVnqnxHtkhBk
0EAEvP1U3KyF0ksCUR6nX5M4ti8VUEdqJ9hcD+iIt3wkb7LgyQ5pf+P1+JM1Z047
w6u4BB6T/YiRLEYzVz/VHy0Vbab2mKnnUDf4MEHtJgjhEmX/YIJ+lWYLc7G8HdfH
/azpasn7/I4HqpajzCl0biYQvPeJDLEzuTq3fmlisZCK+idVOxCYImgvD5KlTKBg
nARcEgi85VlC2Sxarmn/RE5E4EnRA7MrCO+XL7buEURrIlzVV6koN2tks3rIEyxp
4m03wKOCItERUN+96Bmsa/aRIYRYO2ZRYIEI8F1wO4EoMlYfDqVFZzorLkzmbPfr
RBMsrJw21SjR/MUKV9Mh6pePFqiXh9iDD3Uenjnt8H8pHA9USxhp99Nony9GngIZ
FYVSo/YKx4DQYX9WP6vwffm1NTkQG4B1ogRbtkd0/YYXcIAnxOKiRaXpEqLEWo41
OkT1VQTqsUntSxKC6k6jYJbX1iL9zfD1y1AUv+5CNeMGhX5HSNFEyvlqMiDcW2/e
RYbsk0c7eRF18Zd9Uxd95dhBDLGSz5ZtOT6m9P2CEJjd0goWqOZZP8OuEDLV+jhJ
v4sl0DipQfcVGkmkzLE0cXMpz1ABZyqksOXkYRQdx7wFFUIJJwpFyo7XSGqFx6Pj
wMV6ylswRZXHqktfif4potKlnazwNIR2zpRv+7JaG5qNDDPxpmE/5BPgRqiJ+9Cv
pQwlfUpVDwvlMHLdhOXWGXeyduu4FlNMrCQQN9lLzjTsAWaz452zgb95tmK9dpBQ
Xdh9ZpoZK27o4bw79/zNEjTqjnXcRTMepnjST7ICNMhzwOedVD35kmsbJ2+qeiyT
b+gMyuPU8rYA47rBUWF5sO0LRjUeXeNx3PkxMzxswPhMFL1Wz8hu8GoTZ2uPs07U
RWGthZ6Aj7aTddnvEz9ghBVOHYyVJ+HwyAx5syD4jO1oPI724CXDM7s+awPTHP6P
VyXpxvO+lZTHAR90CIVThq1fw6pcXlHoDQ3vs6MH2Bzq1rAG7gwKY0lsVDGUwgiQ
3biF/OwYiX0THUJvqOvWvgGxqV+0i78PZkGggRnWIgdkv30zLjfPPxn/V/rZzk2i
1OiIQF4hGhHfMmWVgxVrq7RgO2WbnMA5/xmwMbSgd171imSGncFmYgszniRayyML
W6ZwOysii1Iws8Dh7aRpALMArkb2Ldeqiun5MtcT+xs+p2BVvIB22hnI62wpCRMy
wlRbRX0N6xrqxT3BCW9dbLd3mjBa2mbEKSyr6JZalZU9J85w4Pm6E4C+Tk/ZaVk1
CAqKBxeUicpOKQ/nN0+vta+HtCeO7iKWYrv6Ym1TFEvQ+4IusPxCp2syWLTcRjRH
wK/LYQfkQ1z1fVbEGRLn2Fl2OYC0nsfdjmLBOhegifuXLnSJq1/N/9IKx9Skmm3Y
9/+lFraihDU9a371Hh2w5K9i+60agYJbjaX8gAgNUsZiA5+uWVUxm5DBgF55iEsh
ueuVrI42L+ZjLTgOmDJGtIPv2TuRJTyXd62Be4hr9OpSiWggwZycxuxxvOjuFnz5
VBLZhdr6EO04YcquETuUj03Pm+DYG7V5w6w+rw59IT/wHxY6Wwf5aCv0L4kiSu7p
OKwpXTIjKnUpi4tamKDqhTMqxpvLxdXziA3U09+NFBX5Y2I8+9UbSfjeeNLUOTyo
gVOvHJKIrR7N/9hKymsRi3eveECwSiEnLzXMej55amRYBzvXfT123jDR+lBtV7rL
vxk/aMgke38NQBaZ3CpsQzmG/kdUyYzgjm+VWPXWT08oQNpOBk9J2g/C/rDIuIJw
eu0yTd1FCTQKltMTq8nfBeqPXRItYdXYseNzghpin/U+vF+Lik4ncCsQew0h0a/L
2/AIWOuK7+cSAqTbroddrPUo3In8UEX3dScfyMUnpzwtpcXfNB60jAFv8TScw6xF
GF9v2oz24pXOxFnN9Enax/ehg6pLT84Sb3VJFybRE2cLgWa5YJqAdZ6xd4lDJJZH
cngFv8S9IIWCRpZKtPyTOVPd+0ibWPAAt/ArbWq5RwhbmaCEOPt/jhyKiq5kWQL1
xs+jvyoA/KLxbbnIdYyZ+hB+RGFxlDO16ErbB8XpY3FqmB78NT1s0PgLVt7zUJ0R
MLR2p29qV0nt/K9EFA32XvwqtMlS/almF80qL9WdFLA8WsOWpi14PeE8X8eHRkOY
k20GaeXmlOP7fhaXHlJbxkCRGRNk/B3QCTzaHEf94xQl3OdnRPGluTq6RkHIGlIw
HrbvDJYjbg5osqD92fsZxk7bCPXqGaIikRHoiy+goBuEgY6FsE381cVUc16fskSY
PgrXrtbpbkF7tBpHJG0ZjgKCxjYdy10IeT4/aqrKZZC/w3opMl3SnQaSPHV5XNyd
w/o3XE9CweRs8Vfhq7VLNAnp/8SX8FgR1nVqMp8AAWC3dyYNzPLJB4+ZsgHYojbQ
TqFlSLGpPuUOMoGQcmu91HmjiVP/OBNA/wWdUj9k+Eq69bvCu+o4kObWaCIieeVZ
wyWXD/ysIkKux991Hp+VgJpiPNn4z76VrbcSDoEZqsrD0lolGt/NheiklShv6oOh
3qded7Fpy1+ZZjjfZYkAObPBIfPzO4CU0r4wqIGdOQIAoKOyGR//e4/XkdchIJYt
4cEhGdN3SF0RvyxERU9hANjqYU5VrzEUgIrqttvwDbvcPNZ+4cjoK5Bx/E00HY3X
EUh2HYqax4ubeo3AXL80t1Rkf4OZs4xeVzBDldQW1vaRpxGEmOLAXM1nZMs2Nka5
/plZxHfm4r/QOlq0Fc0i0XOdOftgYfViEIUerzk1W1ZcNFoIKs1IoShJKtPDz09I
3vganZ79qipXa9rRIYypuyoc1/TH+AGTBNEVEQNL/xNNmWo7cOPTQn7hNKaO/oc+
nxmNjEQE0Gtm5CHUl/sjaUenBwv22FKceo3ocJ8nszcrsoUemzBJeBm4zn7/vigY
002dezCE1OxYcwKqOKNb/dcrjIor0bTOv/Ch0vpSEV02jJ1sfVU7gqfg2S9w2Kxw
MHAWBrZsHdr89D03esfthkU+FDFt22JaJu1coGai8hBlaUyd4hQ6kM5/Bb5LycEZ
//pUGl+A0LSEnC5mB4SGXTLtigLtONEq2PD2rm1hZy+cznamnvdjthKhc7nHSjkz
y7f/qxJ9x58xXEujeRqG/ChXk/HR09lhlKZDE0/BxsEMoIi0BUFMnmDt6igiZ8gq
zIPJ5SZghamCfp5b8L/xDjhF4AwdAFDR6845SkY0oZ8tUZGXYEKg3gGRgjoL2/27
wIpTdj1VIwiSFfg3OurRIxin7ZDF8jqrmJyYn+HqPplvLG+mi3/Yoep3+ifXI79b
tDtyJIjNx6ZPEDMLPCTfScicnXjKRPqXF9gcIEZGYivQPO+fAEQD4IwaVNiYucV2
KQurxgeS/WRR4bgYCgp9fzRo0p3aNZjtpQHbLPfK9LN1O4vbJ1Zi8DMfhjRnYwEs
unpVolQMaJZSfEPXWEX8Au2WddVaxk/rEN3DqEDIy6BgH7BBtxYSx2YNFlOZuZeD
Hujdz0YyU+iDyNOBxlIGwNBw45+jiIeB0XxMiB6hoHyQLLdUa8tYb8n0A3KNEc3k
R5wLusyWojJO19yBsrynt19E41GvFyZ3k6wPDSTQbicKr7wFN3tTV6JIAmRPMDNg
G3pfuaOhaspzhasJ2MjCNr0wBnKZIKW9xXSHH633gfpDnX5fWB3ul1D/nRoVeiQc
yNaX7hqwpbhqANV1gFJKk5Yax3u04n8+0J2fb3fhRs9pTGWVOeJL1pd5DEzwiXEH
rV5tKp9EJN/HxwJGXHOlLd6JQ0+/FPuVXI1FTnw6HVAty1xXH0UdPs9jsfFMRJas
a8z6VeFrU8i5lcIiCTTmapFubl9v/WPp2URA3cDXCHqnWK061LxDMW44T5fu5SlR
tS9nQVOGt36zNlG3Wi/r4aKHm8ULBwyE7VxhzSoCtfb5/71Tem/ZmDNA5rP925ww
rdQhzE0LnVgCUJByYTxqqnHtk910g/RqGCk+XYa2qrbQEDQ1wpsgs+Z9dIbVyzz3
hhwgZIaPzWW1CLaZqd430kfa7eq6xa9HVQUbO0yFemWHszgQBQEa2s+v22gwPCrt
PCkqZbtS6cc0wUQwytVzg3TQcPUaWXvFOdpuATc8vbztz1bhCih81bc7PA2OLzV6
UFdP+1Liu3OWLlkZCu1Fu/ICJ4Rc12/S+IZlBLrctYtJkDigrXx+wRRtAPO/MgBT
2hRLmUovskyIdmEMqTvO9Ium7QzAeIuI2xlT9yTuRu4UKLZZnah2Jc0uKhCHdpvI
pEPrSl/hm9WlDRRiHUE0eyrtyj0bGNAWj+LtYcOncTfcKoviSq57Z8purNy6cksA
Mxv+jgZ7J5tzWbDqCVxv3iMT/ehSLhsU3tQqFr3YtiB4ZOoqkAsdjLEuvXdgnopQ
//ugBmq2s05NmnpL8+YLWeztZyKGjA2vLrMY/MoBc6Q0cmwlV+ZTxeYznub7KD4i
oRKKNT4ZQBVsaoRTVrLWSt911mIqnj6eiKCMVaZcyUB3FnBtm2MtmYOWiQpD4lew
CYmxqlP2dNjowUf0jWaNVKyLKDL9IM6BQKO3Pf7FGTibIsDIkbZh0lAq32F5DIRk
VgRPYBvOIZy9BmthRVtYJmLMC5lXyKiazOoI8f7h+MGxyZi4zxFKjWyBc+Mf3M1w
ystBR/UX0eqDZgEIbOYd99R1UlmqwTJZtBJ8NFQTSonWOU83UtJ4uAj6V0gn4Fq/
FbxSEx58C4/ispx3vcZ5ayZyhIhFdWUHt71zcvjJbFQ3IhXgYNapZIRP6n0ofdG4
1HBuaTFPGx0sQCPwvkIrvhqF6PR8oJgqIIXyTMLUrNriF/tOo9i/5O2jAPxRlZcM
3YEL8yvYxsGrqxF0bfv4hOKjEotOXYs6w3L9vR0JGm92DSvhRXNAW1l0dPe1+w8B
+APCwCDi17E7Yh2WZxUW9QY2E2gFKlapKs1JLqiMdEuvBClemaKW6AIRw9NYMbZc
aTgSOEdNtjOuovn7CN/OGTMKLyzHjNqgiarDt6FTKr3wOsdJlg2k7je7zbUjz2H7
qlKfmyAGHognxI3MkPznVxD9GSQif+RWiBAbXicjcC7C9XERzbI0aZOfRJj/yhjy
AuX8Hp0hKaeCUlCmfoaI0XeFKKMPwuxS3Q57/690b/B/am2FISLGzZyha20octfD
qGJQhzCMyBzn0fU4pZjc5AtdgQkFcyV7WsS3AMVzZdV2kGnJPaP77/9Tzea0f/0g
L/owk38nPPKx/bE1YHDCinuD0ALJ0xEb2e3f7FjrctRpSCPLI0fp7f6jm5rWOWzE
/qqrm6RFyULKJbyDucOcm/TE9qavfUatxI3x1S3QOXXSYy5/yZbu76gTNSMLiO2x
UWbF2HqYd9+BeiP4p5agO7+FoBQg0dBKv0y4z1yy3QB5azhaZBzBCu1QVMMeGdvm
KTtqLnSwlcGkZImKvBC12XuLOjU1abyidEPSfjGlcOwE4Fo3YwBzGcWObxZvwqB1
xX1u6xhbFpXADI2ZDz36mAnTtWTPoByKEE4yl0U3W3q32tBIJjFMcVl730jgustp
K581oXFaQ6yYmvZrPmEwqnQXpAK4LS0WKXHIrWrU4VPOIfIaM29f07GlWCtlHGkS
1k697/SJEoxcM3OYpkq0Y5QL/VSyNs6IYGbnUBjUsE/I+4eIPBbl6AG3axO+LrAp
TIyl6wYEQM6VXft4UYsSi+7E2uIoK0+ylYXHgET5yiQCEEPjiOgcLuiNu3+R42H6
TE20HrEVTPe6DYVvinzOKYohC2ZUaWwsui3Vil5RS6hW1YKBX/HcqRGGWP0GBHCA
B3sXmZ3TkDldxbT8989Vq8LVjkRroWGJXH57K4Ueru4Juw6gyRozGsu5v7oyt5Jj
bJX0Kp/gfwYWROr/YG7SmWtA3sj6WcqOLQ0FbvsNjjw6EgkOQDCIM2ECe3JAjMks
RaXFhhycvq5FrqSY6IRY+HKLpsPbW98S9SdEKgUf3X6x0kEmOhmDeGAfoVG4hS1f
xXV3f74UTeHTjY0z4Ipw4kZQcT0HsVlT13AZhxI0zTtenlrU0KLzaU14aimkR/51
cruQMt+ntFdxTL1eIAxlewkW+ft6Ztmm90eXDyKe7Yy2+44ablQ7GnZEyjJ8Nc9o
/oedc3HT9RsTk/ubCV7st7tsqeVbnCSlaAKaUpm7uWlVdBUFJcqgsitx/jR4IFTp
1Hw3jT8ZGELD3pOi+LqdT0LaDoDA7zFJZUsGpg0xaf+vABMbfDVNCvn8BtqnjA82
jjxVU5EeQiPqF1zPS32/FwKoJ6B/OO3XMZ18K6H7nO7Kga6n85/atEwhUTIVRnse
7+DAIkMH3WDj0OLiUhxVtkRjGGf4JwJ4OKYzNw1LH/8IAPEP5VZbcqpl4zRav/4x
s8YxuQ9dS9+lBKnX2dXJ1k7jwkke2QwFvdOT8c2CTqjDnBlWbYCH6UyERBR3IhG4
6No+xZILoH8G2GZViSRow39rYMnE9cy13e5QCScod42uyVqOpKtNvdqeyPwpNOTi
pzJ/ADLTErXelk+vPPenwS0AXHqelQ4lSSNJUhDtw/C1WrGj8qj8ynnYpksKjGdB
fuxDKf5gXefqF3Klqhim173KykjnVbJnoiS7Hj9A9MJQwZz3+UYT0pgxFyVJmhlU
itGn794w6ja0NKvy480C2pDvjacI/vdjiCUT4LgnbYmG2t00pgy4kc7O10iJt5kd
jLiR6381nrmSrClULa5NyTV1dKSK29mju/sMGkPspU8ApAqNmkBoQSf/7Xl1JIyG
Yyk2tE1z7ur2bJAIP5krAA4RB4Yx7YkyQDbDKpPXLt9ZKCJRUQ+QrCXHOAZBvfxw
k2qM6WMbQ0uznod8bnpX2dcUck+KVkNOhc5/kauicBbbn9n334sIVKJ/35BdFpDH
3BFVcfXQd4uSdEH+zcWSitaXExTX/DLNK35x/7eJopbFUd9g5hXZsLWrtH8FZgNi
IYACc6Vj0z91uLtlZ34K5/wo6maVF/jUlDrtRV27L23rpoDgGWekkjKKaI2v71DZ
bUhsvA1vPEVrYVFePsCYe8zLRmAiL8Th4ITerpsTZTq8UZDIAd5j4bRDmbvDoUyc
qFei3YH7DCeuSNpLPrkoAsHiQKO5DH97BrdtUfRkVFk7IZ4BFYc68AVT1DSVJptT
ShdWzXhQhoK9Y5hDWUfqaF3W+r+YgiyrY2iXXLF+EhK72pjSKbp2k7T1dBphyjle
HyxdYnbExKsCNvBT6IHgELiwvb4yGV/jZPE75wBBdZ6iRJvj02EY1o5XPXIEeqND
junQ77TI6CgUCkB9Mf8tV6hknLzn7U4rjtsxlDsL+o4ZDe+6B4Tk5KV8OQQFMTiR
bG6xSttbBi3T02FB6A+LNZCd/1Lkg/uKEu+94hrUSeCvDSY0ZgOl5Gpd4I1/LbXa
/2dEt2be7oMRcwmKTy6HH5slw7C+FBWj9jJxavJWkOPpK3HUnChatzkT7HLh3V6a
6wHCywxO4nQt098yUBhx27LTzxILWE/wUjGWQHV9iNDyaeYsg0XLj1TbOg2Woh94
uL6bk24orUo+qCpu/LCJ3TpmDCrQ7rwzAlTmGo6t1kT1G8Q9mQuXwjsX+7hWI9wr
lfPvLx1fNq42G2Da9NV0t351KMPzhVbe9+P6P60sAFQeEWmw7V0ClY4aJyGHvR8N
RjQ1nd5BiHfjLl1OhUjI5X2cKw4c/EBzT9TATP1OIDuYzE1zqNhwLlC6+AA72IbM
Mn0UHtdOwC8b3/plpUTv/3Xe+Uhs2UYesbxpg1981TrCVrhLnnMeLuRBO8OLnd1A
JRTyU+ryRBgUnRXWP7RyxuQzIyfO6FNqgZBuRKLXI8p4kK9U6Wun//PJkOaYSIf5
liOO6qRFkanq9eDlwN8XPWqFZK/p5eMGmLKowYA7S5pAJc/Bbh1JnmUCqZaAmkxH
mUpng3M0h1gSgZPxYQ+3AWNZHaOWSOv1ak0PcslXGJeXeT2o28AxZzAYKHDQJScN
MlH3n7epROkaG/xqZD6IJ9eD++7OGHrNBNYH74HQu92uHTut/d96halaklwBzs/o
7DWY/cKVIBLr6nsvhyF3JF3QYivAf/1v+SOVLrNCpx51bf91XmKDMDDIG3ghGJpZ
Ih8p+nr6DVfkHuXm8BgnfqgxgWC3rxxCHiUnNEgPe89HV22OH6fLi1DWR0tsGvg/
1uzeKZVKNPuokj47gyzMTqVoTyMXRt1xQyqO/mTCn0Dmnzm6+0s9P7vgkscs5GXV
fa6rAh6gfgyiKvY/Uiu8KhPKS5I6g39leWrWB4pVFW2wKivckNdu5BR7jikt68t4
kfQIbleKYdKhUprubEFZrpO+EMqMxxLcbNm3k0V4IIWqjToqa9Sen244exXoD3XJ
ovxKaCm+suLGS1wCyg3+7Pwj6jr5Pr9zP86oZBodQbneLntr+hU3HMq9EvNJ4KAW
Y/p6Z/QYAOKoO7Y+ulkD+R04WcD9D9Nk0Xy8jQDXphHqFxXgdVLVCdZnsloihgM6
o4TeA7t/tPRImeEr9ugqoP3916KSgw4IXJVJ4Qzh4eKSS9FtOVIHSjHGaqltp6a7
2FAX6cpfScAWPO5bsbkb8pxVlim19t3nI63eeEjN5EV74F9B6pqCdbZLOiYow9fX
c23HocYklq60fAH4MQS2ViHaSEh5klRThaY1qVO25ecmieqoqdCVdHrdLDuvPm8I
LLAUVU3sjyb2IX0ZfHn3zUqYHaii1wWUExzMYogHti89Gu+c0GDsmSToJ3q6btYi
3PfqcRb4wmJsDtIjTLXRIinIHdIg9Jt05BbIHbqaSlWDVgtpTOMj11fdtt2M+6qP
vxLabUOUMjJ9N82W/NKdUlDbk/lvXVhoNDTGbnbtTQZrZqaRZZ5geLBf195yhEuN
kOwbBRyKDQ9AQli35KNa6b828l48J8w7vi1ydxaZlIBzYJ4qZFQuUjsKXs2tJkoK
Vbr+3rlJviBzEFK9zV073dPf7L+fhInZPg/T+oGJQ7j1DHzqft2Zbs5aC2tdxp7c
7wqY2y4iS1/VxDRbz8UbryV6HZswuRMcDo33N8ciTNTYUVHn14wh3C5ZSrbKLzBR
KkaK1UqjllYA/ahIvXqG1EAdz3juFuubx29ZW2tHCa6/4vtBIa78slLz+ftwF3UI
Jequ9LpmJxa1ZXe9u7LOMDBs2+1TgQMMNfRoKmern1dIsHDVrXM/v0p5hxAwVsSQ
1VoKMWejsVeBLULi/VLEnGSbtG7d0ZcZ89R3Ln+xmtQz6fSflQxvUJGTDJDqURqB
FqdikLygGRgoN7E0aCyCnVB5F5aFdLqSpCF7Stp8q0b6Ww7Ca9qakr2IudpOnyBK
zfASiidXYPscY49UczY4jXx/ILSIDFWP1TkugkK5Qmu0rX4XnuT7l0dX7Ru/oQzK
ZLATTP5Vcz8SEE0ddyqiiZWiO9fVl5ewte56FecsiWY1ZP/6K8JpGThy789CcgOw
Vl/GityNCOgvDTIxjosIrkzzzIGf4ijDhESmf5VxPv0PGEN2ZrwCYpn81MIIiggP
uYFvQopnlSTYy3arAqb65cMjdR3uKG9zQLmmE63weH4kh7Cb2fbzDOgxSJILktB1
SMVr9DZgg3kwO0aVVsqquc7+mWX0IiyrnGNucRaLoh5KU5Q6i89a0hHb7+rgam+J
R7ZMp/ieLnLCsWdDSPeQNfWYB0x7y46v1y7E0F7j4KDG6iwqsyJsR+G9ytJVG0N1
6OPiaumZVoGeMrS08W05xC+q15YOD5wThR9lxF2WzRUWnynz4i4U+0N24KgxCd1D
exv4ZmnwrjJykApFrJ0wDL4qUd2zDU/kBHNVR7vxdF0jRV+w5PT1WfbrhjfgIrj4
z/QnKGUwpJCGQ8aykGn/78xR9YIJ9ZzQhILlKqy+PJVeeFhDUoqMbFBBmYMCPnDw
YBSCzUiDJLqPtrNvj8Bu7v8ij8qjg4F4Xz8sRNv7b8g7DUa/9kc7NfPAe9E1Xxmf
zX1VnuRjIqsLGuDnTGmy8SLSQzwxo8gEFLVSS5iKii7ZDjOMJnxRSR0tJdPM0Pr8
Ef1HT5i9EzDjHn7d+17fCKh2H8bpCijMiVQuVLwO3bbkD5WpQwHcP6wAaMRcgdYH
vbekVtFiEvF2sovcmqppzS8eSkN6Patm1+0H95oFXtYvh8oPshoWCg4E5BLYsId7
61bz6Gt9Ip0xMI3SpsdwfBmn5N7fjPTD8tTfWkMK1qJSwFYxqbQblamEDEwIOgXm
+7ScFk30G+BD+/u3W3hpn0sFlCxKLmhhA1qBF+0gCNO68DjnM++fKp2V6Ttv8NL3
etrlI7zH1LVpJHqy3YjLZ75j7fSXXxpbwwukdq0RuCH8R4AjjVcHyRWb0rTvknIv
MF/iCWr71RsP8L+QbjQfkDRhw4W3L7rllBqE31zk9RhaZ3+LnMl2Na3fFPQVXRyn
K5TEiutT+ukGfHXbLdRyCmgmHTBca6YPLiqT1UupxeW+wzgFonqW4DpUAtk4scqu
IqTbRfc4GUS+RU7T0yTnZAhZ1OQus9FYOlmb4jFRxG+QZEXaAY/BaQqlRwLWqEs8
kilFcjyhAf/SghIdrJe1rASSv070KqOp3k6Yd5gebOX1gIPB8QCRoPi1/BdUywDd
fLO5JEbfvxzMkYXYpoMLfkND3/z3+fOrspQeUwHvxeRDX7E+3+NacfofWUKYmg2p
CRC5oGn/weq34m5lDIraeMC5vy3w9z3dNUISG7GnA0wJktiQ9vxg2wNaYPXqyirB
JuQBTC/5WIrLINXo0BYjXQ0/8/neHEq//rmWIKQwgplekqcUZ47Itza3xGj1w+YQ
lCNuLkRxPmUFTaPDYjlXRx1fHkevznF3HrYnd7Re2OjI4PlegcK1VHotbIB/7OJP
kitQ+sPNeEjV3SeuVs/+CcOPViu0mqtfq193CSnkb498JMrpJRU1981t33OS1WIi
G3cPPGy5PSKGb59NZTwTIh16cAu57ufvpHleh8UCqWyJyLnIldLA5M64MuTA752i
nVD0R3NfM8rHUjhvrwteYxpHoDx3b1Q6c6KQlQDnCskFnv6K5C/g+b12VMYfQUva
WU83PNWLKK0HJvgBybD8lv0Evf8wWbuHrHhukMwM16ds79kKJngpPEgfthnUlwRV
A9rDQeV5evzA6SUpP7eQO7u/7CC+skmYwgGWi1PEy5heOPUDbdtYllbo5TLPh67G
vevRAdCghbHNLWULHTqfRavCEA8DhA1S4Z/lbTBA/kmZZ5wQfj+S4XGo55zJGk+y
97I4MhquiIc5k78yyHN6HnJHAjdfxb1QNWTeoEpMA2WnRKslrqJJnNIJkOPsiOaA
cIaLntLKFq6pKxbjM59sidjOta+Jp6xaPZf889Rfz5og+XHN4PNvT7WW3l22a2Zd
y5OnZ5k3r7j1kEGNP2HUXoMo49tEdu/GWt2acLPvIPm/hFoS7WM8J+F9E8qsX/XT
swnIy8++s1E/CSDFprnbkA8GV252SNPcc3G1xwL7LCEwNawV474MFXgXFOtZenOE
xl7eJ6U8EEmXM393bYF2kUzXNgLca/K/KegLmiAIWn+X7EzM9EUfrZRSjTltg+nc
X0wuCYCONkUqbHtCezE4pYidwCAAdamlo61H+pAZFizrVB7OzhrvZj/sU/pQdb4g
l0+2vbBgT6m9iVFrDwC8CpF9j/MwAi0aFp4Gt8lb4PlhzrcEJBlW5c9puH7QjjW5
esM4NYy+1Z14i7yjcVb4Je6ZCcpRynansF0X/6IkZyGx2mpYCixDqGs7K5vG2FlL
OPXR7We0i6Hr7rObbnNbgXvKkbJAC+udPVCFwLtWlWiKfAhGNHKtjXUN9gwcNa5V
vWVcdygtezCfBCwj8Gu5Aaxcfv2SQrF59jL/k0CZ5aQNs1zOgT4bi7OluL/RS6Lu
bZ93jSXron+QNJxYWuTgXhDr7Yipc7lgtBPX9DJ5KV8Spu0K1cmPCOSBserGGpBn
a45e3yMqlSxdIAzu0k0lP9bt4ik/SzKKAPFGjR/B1Iq6JtOJi9j+b0JcxfJ2A2sS
S2+1KjJbFM5NNURprzqDtc5EwwKAeiNXea6SLKUAXGIwHKpDoLbU+mTc2sSwYB39
nz2DyTGn3DOcsJtfQh38l97JeZ3MuNL814Hi9V8eo+xS7Cxs3DrzIzBgOt3m/n6C
uX9OxCx/M5DMHWHLMz8aFcKaaulveT7vFqhUyD7SnZpyJba5Rnqbq2yzqXylWPlK
n8mmYwTaygaxoWewz9iKXkLQ+llYHzIOUJmyArg4VRKj+k29pPxkkjyD+bQfUCBp
zOPe+6iiFzzY9e/H1ymQsPFasJFnKGxiicxcL615NqlVfbj4e3mud7gwb296r/qV
K0DY7chlw54znbvzsrWF3hDv8JUnypdoC6F3T9KBDCC++erTShStC1Sy9yOsOki2
u886CYFCpsAx4nDfILNNFJbycSqSEAB1jETuIWEHcF63V1CXFK5VSXmBP0Vhv+2a
tXyhDr78wQILeqA8RdpqWo+iPr2vulWobpd2yjOlgt6NxZbJSAb4XsGGe83XWjn/
qSBm9jhXbn3lJjDdDOuovby98WcGCxiTdOpAULziU6rTcX3liXmFSP+XMOAB4JXY
0ClupAGDMDKVQXPAt49T3O66XSRfgk9ExbtfUB7J2lvsZ0ZGvcvg0yYaodKsp84e
SeUgdgB0IML2fKfBdB/OqR18u7s2BgpFZYJ4VVdz7zsFKJx88EtPFSqfXejDpPQc
vCw1y285XDRw3g64yClyFV9Jt83A8kU1WMGprk2jRYHqJQRBUNggfDqO2YM//I0Q
fpVnRCKFJejOtZQQilRhHEEL5ptevrXD8Rm/guz36OPzibRLU0dt3eM6Nszb5MwJ
X76o/Mroety1L4/CLwpDh0snLFe3yfpv+YYTcEs3PVesvwSsSG/h2BBNmVPEab25
P9Awm/go6gcUFlIyWeujPvbQnDWPMgZmkzq3MTFQ7iHYmQOio5McPaaTFu73qfmn
SQ88U+wcl0X1qufI2JfYTqO2znCfIZJw4foZRicDs8Zo5+uIMS6IAq4edlFnj1d9
jD50Fl1DEpGu5XBBEvKGVD84kXWj3Ej6+lUbvEJHM2MpVOh0N1EEFaUTmEyOYlh1
cfpbMNFDGQdeJtcwoE8e7nUqlw9mvSoasJt+Jkrs4XercHuqK43RUl8G2bYgqvaA

`pragma protect end_protected
