`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
kgZAwkb0CJkF+Ts1NZpun+S9XKA3oZHvYFceRoRUaqerBnRqjpny2zBfJdOG2gBv
88P1wplIne8gKJpntEFvi/IXNGWTx2GKN9YhZ0l5ooms2SUi8SS1vVdOjsApwPYn
KbMymEXwUXgJgiRcEmEUHOysEQgtv++hCEgrelnQ0t4=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6000), data_block
+2ROVMB3+1ZW2oXzcZfg4JoUaRn9Sq5gEzGmuHFHY3i954rrtZQLfI3zJITnZkgk
6M5GXEEkTAMWjoSob23i+SNZJdEZWWiXE+0zK5CWJRDvU3rZjOdUgdYlBBd7+TFf
YbadhjFH4SFGNh5lgudQM+6+Yihf1v/t3cU4MNNwO1niEssMXhOr2OAeGtd1FySR
zEPyuljZFgFo8n6dmyBCII79HmVfdZCNvb+QjvFn62AvnISzWkBYDo1V9JBpCcK+
SQxkZT+41UMOFbA6bydZN1inA5h3GS3oxEVhU7z4RpWU7msLFEI37af8R7GT4oCt
14RY09wFFdUOmqs9BL0ANGDLfeEZBmU4iC5QYN2TfXH/aEIYqUBnqzRhEwTMAE4J
vxXF8xtWoV4gVYFiCYIVcIhIJxd0JrVvGHmU6+JbIthSaW77ezBaJ2jWYEwQBV5n
R35FueuH0rX58mjlLEs0j4APrCxa5Mx+PkgkRaqwa4fQq7+HGrpReK2465Up+WEm
a2MDOx50I+fviESpmumx7vNvWWAwkEKpM8JmHKG3PLfx4HVCW+gOXhcv6KbS48nA
o2rh3amVGpDfmWkbv68nCkOH347c3UOv5UNVt57bn7wncE04Lww2wl6oPRUOPw5Q
USwGYwCYFcgCAvyc8cILHU7PdfY3hVZCEA0Rj27UQWcUoymKteANgHgth0vfUyhX
C2165LcmLsBQsuUOoXvgMwv2IdwR5OmmpbZ0o9MavxqvAdWYAmw2KKeo5vwfSKYr
J3otGdaqTJXgusQ+q+zx+DZ32MAdwIlbaUiPv6CGotNOxNXX0XI1sQkhxNj31o/g
mozfM9m5otaf9XQpdSQ2ctLF0aX/IoSxMTUghvOv/0OjbrZ2kr77Kkb/kT1mfts4
v6lQo16mrvOKuapiJN324oWwXC8GJcjVm4kLxHoYqJr7p9JrosCmR3+2l17rZnW+
0A+As+uS8UAx06QJV4QEwytszeXEXfnPuj4JyB2O4uQ8aybN++KIaxxBZ6fRYahK
HgASPH7V31zeKP5mBh52bbnugOPaEzVZJj8ZBkzCOy6N3lxj1nO9o6WxZ1iWgbkF
ufpz0hasoqP4BKzggv4dbiuY8l/VHD7wKOhdOa45FFM6WTVXzdZX4J2YofuZhPty
WsJCkPkIJ4wpmh13UdC6dIYfZxZ4yJIcZ5eEdcd7z4Sa+6YZUjQoRfurHO1CObHs
Nk732ku7yLbTUeiD9d7SMwrrGnzoBGy2vfjFUuF/KSJ31JICChnwJS934ACEdWZn
Dlje+mppc14vjCf/VaepaYD+XHBZ9qL84L0thHO6lnFUZFfIHp/2c2onvSpVYdYX
auZ69cZAv48HhGcPW+vMygrFIhWjhoPcBtIRwIxDFTtfxlJqhVqFjS7/GHwuezVt
5fy/jq2s6zPRY2exG0XKRkvK6PI3bb2Bj6GY7YSjQ72fjbM/jZKZw2ziiV4qlAVZ
EgoRVvsofHFg22DLV0LWa2W9tIHoxhWp5dspkCYYKRLzcYlBMDfW36y1U6rDifcv
P2pbwsxyW251FtSXBZlvDkSXcsdeUTyUuaZhpHtqmF3TKbv7GrDxD7M/GHuwmlys
XSvIvVvtd3TTrSz1IF/6SpCG6WQhBdXiLmBom6r6qGfcigreOWGs+MhuMVZumsMW
Nj9u91qz83MzXgEIBB9lFx5WTUg8F7VgD+rg4Oj4+/+mAaD12eEynUbKtzde9Ooa
BIgtXeyaCilURKaPcgamJHuoP5apALSu2Xpj78b3/oLwjg2GU7eb5xhPBoEqMlFq
h37EEtFabOaYBGzVMOQ/QfywqXEHmNLBwAtHRyC2/Khdnm7/WpSQxYn43dQdEEwy
3JDVGbP3Cwryj1TSreXhqUuLpZNMNeTaszGL4YuKrnZzotpEz8D1BWwnDIZ6vb8s
/EO1hsFE+HXTlHleLMHjwNgHn2DIkvpQUhvLp4gJBUWQyxWeiVWOxbb1SIUGl1LN
uk3AQs4DzEnOlqZMfQ6/KLB8u3OQgrc28YQBc7NoOaL+Dz4iE7LuDFEelauIBBlp
+Z8YD5y+7d9cDdy43PJokDTW8BcWGp6/NBQYoBoh8YvXBiMJ56cihVewlXGTsniQ
af4VqAf3/qoXIBUaboNtS+DYT0s0SIe1qwXq8/1jtSTPB9hnUSG+CIBkCivVad1f
wQ0+9Vy8+zr+io6Dpo4iYo/lkdrX0ubzr2ZLPMfE6gDKr5Ryq32cjGur9sgfjQYh
Fu3wUeG1KS1UIiz86UakJC05WnZNgD87e+xkIw651lnfuEitH5LQYPaK+nm8L/p3
SiW8Ylz8tWHDFSQvO+D7/jpw+EWNoKU0j99EiHHdhePTCPZULHcVUEVlt6/b60sF
mZgUfqfeUiWuaWOCO42YZTGMpm6KUL3YzQGZ9kF2SJchP35cB95aBLbshBR3WKnp
was254Aw4SdIGPde0NbPG2EFj+uRxCH43Cdu6EOmwexRmo1O87SD6UrGq70jUtdD
magkVp+2ZaBrfwWkvnstUczEtdBUojzV4THN9jIOcbeP43ul4caZvZDTUKIRUJIq
xdESrgxvkiMMtAV+KMfn1a+D/Rd55cdx4yAyuISdG1oTvILEf6G5gdcLP2MDE+hP
U6XDyDIkKH1hw25t2YqGvtCxp9FCtHwZ3kvjPyWl+1iTe6OYh2B6NsUHlkpfpC5D
md3/ThGsprUphUhtEgUHLIMuMT1Kv4gSV/yL84ddckf/Xf6b/v5TMFuoErUPAgb3
zDWL61wg8QXRaqR+DxLLQs36L8WJ7y7YpefpROfqFhf7koxS6w8m2xFZApa5kDhI
9ZFLD4B9u/TKUYcsv5F9LdsQw2DHfNnLgd+bw7F6VCV0haNyDNtGZkXWLxyYDvuZ
TqTryG4y5c6j8y5G9GxXXDf9uu9dne8MPD8cVZfI1/ISWrYNkmh8YNZrR1bz9hLj
BonsaRFyC0sNaayGTKc7kcF+8yG5Ke7zZxQ/i6smThzLb7jLIXBrKthwuV9EUZVd
wTq5T+RhQbCUlAjEuU1/l2tZ8jhKgK0gReTaPuLYudSG7QbBR454/GBonLluJFpt
HihtCqL3QZE7msEUHldVQTHIvDTeGvJEcGGQbKyYd+hZbXmwrZKBDg7q7uTHCixO
FuIBM1EROSD0OrXYVQz4qcXK5orFnZgtwN736Sf/WhyXiQ7ySEOXKQ2JKoSg44Jn
FTryACde1N1tvAUXOgkqNYGlO/92u1P2kdDXMPXe+c21l86JP4bpJQnQSgU/E9J4
D2cTm+3wQ9EC5IQPlSngA4xdVVPt5i/95yV/VbgzNDe0ds2aBSaQhEuwMMLF+nN2
2pWGSNLevPMzwaVyvXMA9sIh3CYqgZMid94499gFn5Ni35hTsKk0DmC7UDqFMLNm
Tdeb5CwQsfK/i5KoqptoVF+ehRHw7GVOHWadprg/o8qFSJV3gxIyVbRhtqhK7X7z
H7C9eoStbOYWxYX6G1gUn8fhfAKHL8wTslxw8JUwRevquoRXyyk2sHjU58zOb9Rw
P9aEPyetzTsEVSZqXu6loJAvi8kFIIIxpZ7czM0+VlUxlQtEsLW6D/v6RokCvkaC
rkeFdr/G9Oy8kX5mWvhgvisyUDt5YD3xVZt4XCjEAGBMoeYhpBXbaamhQftWbRut
E2q3NULFCbGa/p+UbouHa7Bdpuk+X0CnTIpDY+3t89icLgjTsC9IeYIK0zjF++Cq
Kl379+B938vOa0pjfFzn8quhB68SsdMsSpzBLf9ldABWA4OhioNmDDcxxIm9ganX
usQ99YZI24NUmhzo0UPEN7U0QxTXnmtOGvM/3a228eS6B8zFwADdCbneGOVMmGvC
hc+yPaw4uzsV7ZOCazPmTC3FldrF+y3UJdz3vH3pZAjG7JQaiYWXagbIIi2jgKh6
uwKfd+tfpnKgEIUKCy/7k5GXerD7nizE2N0zu/zTGAS3510lMN2REzYLwf7zM4+g
/JUMKGrR3jaa8D5yuyXo5C2yZG3eHjNfONiQOA0eCBrNv5Ax/uWH7sL7o+Jnl429
l3aQyvFI3s8py8Lw9KCVpD2MQwZTnTz1oZ8IW08oyG6Gd/lTuQyrNZJZqbVqhI25
TIGsSBWCPT+uvrGf141elUjUDP0qZ6Glh3Dvkyw0/sIKmnBk9tnO9Ut6WBgV2lOV
R6r4xpYbO/sYeeqxMke207zTI8A5vD64TzZb9ENHT/aETLAgkdlUyav5CleUyF+B
j1cl51a/GwyYt+/BVZ2JPRsjL+lyPJ9Yd/T/B39MKYovJZaYA+CKS/2arhycx3pD
T4n5Ii18r2wq0na4GLRGx7Nkp1QOOFrR8BX76Uih3GZIInrjZP98YLt7TWr8lEOr
JYl7Avga6dVFHN0m7FJ7iR1Lp21+15sr39HRn7TWvLZdPpBp1x65eVLcffrMiJD/
/Afr1bTkay7dzU/9CjOPIRzDQL9nWc1IslRKqs65Y7cgu4lra27FT4ecKUC6RPMi
IUwYqthnFd4XMC3VB/P01B3a0Rr11FCl2BiInUBpGsPjJPDztG/CM715SvK7aonH
40WuIyWlC5GiIH0eSbpoz2m09h12/g8Tczphl4BVFux4RKL3OV0fYEcjg8e1NaQq
AoYylwnEeytgdvibsN2sOjr83vVHdHmIYTO9CWzxJgY4BP8/1+dfWCtL+gJ5zpnm
ZC9uYZ7ekNs3pDNKxQf93/ebjpIGnF6k/uT9w3A4JGDfxVjVU/1VooGZ6zDFRV+Z
CBA+yXOW5QC5c8FP1sae6dkVeLgiJB4TbPuRxrQF3U1CtPz8BhADt0XnE+iAsFGp
spxDTCkVBWPCP65FlpHqkB1UPwUNiLL9WR+p860mM/QcMAZlmWiDnzJ+Qtk7ue6D
CNgKhte0L11bA05MrMpuc3tO3sEZP8uzwUo3z38KuaFtrujTU+u38ze2f9XGiSJG
yQ0Lm+JJc06KuZTxkZ0Sol/R4T5jYD2A3+ii+zg3DmZvwKPdnGVZBlUX1KL0wgwa
z/5i+Uyp4MrJo63o5GEQAIVDWEaH3Xb2lXW+ntrOzKkn2hpwmHwt6ryxYiLGCN/A
SW5CgVjBRePo04z5az3Q5+oAWsT7HgpyYK7NldEWUUN9gvlYSymtgDGTNv26OwIl
636GFCSYlqVtY0x5se6pnfzarIE4ggGwU2EE6f6wMVEo0lm7YmskpgAfFBNvh7xW
8e0LAyn3oV8LoRbl0gN9vmtCtMSXjE9vHXE2a2IR10+0jr9FmSHEMarDLNKVrbaW
tqQ7wfz0rbZlH+S9u1w+lfMWVTiwYKUsORP9MR1IRqLC4reIQputvnzKAcr3UkCB
9ZzjTuynB+Xf6rFaEPGmfy9Nx6ecInh4q6N3NJ7t3qBhVK0bu/DCvrhWvVCqeyFD
dYYdQ/+MEO65shlZgnISg7EP0jNuhUpmQf+bO2tw7skIjmOBIQp40bJZkUG7q4Bf
H6eOiMmxAR0LrxSlELJBnVNQWgo3Ne+0Uh5zwl41oXdw/JOF8uJPtFFBjB5bdju6
3f+U0pbd/qxIX0Fklq417PAug5eubmnz1/lJZv0T57MisygY99PfbY8h6dgDdOCd
kbcIqqAlI06SB8kUh0UhKUAGApMQ82N4KxEpuknp0bej0NkOqXE9LJnESypS8Zel
TJDgB3BwFz+ulzNyvC2+8FL5My2SvLwlerP7gCSLmmOcXwAMNB1GFGqcvDR6vflE
BcPyULjWVmNHyMYHBmw3NNfwP/hHuojMoBnLUK7aEWYmI3NSUjquvL+UDzIzBZ2H
gAEETS8Aq7LWqMTercyA6vnsz4ujKk+sMKP8fLTdSh09ccM/QHqq3iosKCpZVkhB
ZKa/NtuZjhRqWC7KfTwgiOZ6QVz/34VsnCKw1uQ8Rj5RdXPoae0SOD/lLv7kmkpC
HgzMeraKZvHIfYN5/6fjVF7pd665dqojPohU+r44zxeC0bNWy/sIYfweBCSnksTH
QIPGFtoUwY/uHNj+RLbpZyQF8YMTuvnQJTC4htlD61PEF//Jk70sjEBd9sUb4bnn
xE1kRGn25z/E9D+V1lf+8LY5e//1T3DSoIcN3xFSZnzjXDU7JisN8YKIdcLOQYo7
zWr8L8/s4CMF2rd/4SMcgwiATXNUjuIjFQtqFqeXoqgbIJBoI2PiPvD/CxdKPFuK
ylAHdrDIFls2kdMQhDUEBQhXfZoz9G5s2GeA4mXI+d2mNREY/RD7aicmJcqwgxGr
TR3iO33DrAXJv5LxVO4/9weXhCpcjnhVs46R++xb91SOU6uHLmsx/rwvg+rwtsuQ
FWQ2yhQK68Wct+fHPa/2mzCu15Oa/T94YdywmER1tHjKp5TsgiqunmdfXo6lMOFX
P/Hfk4eu2TyZb/VYtpe749e9HVKWV78v4BYVLappd1pz5BQ2uKd/zM5ZpVVaRBZ8
jHl0/oWxT/F0l2jruGYm/ykjp4eWAxv2b0te3JOdXQrRFYGg4GLRd64VpbfXRx51
NsHhdvMCDLqFppKkhffLr/MhPPg3hte+xB7U9xpWSVs7f0HB5uM19i3dkw8pPPoJ
Q3edhouoxinuezJj3Kaq0SnG1TCdTvFwM1hnsXICc3wFNPWxUJ2FDs08PC5/oHGP
aedAh0yvz0v0Fp7aqz85CdRpGwnzHY71JHJaFfEfyXMMJ7kNvffCXa1bNn2AqWLF
+yvtfhbccP1YbZIiLdwpD4fkUmt1AhmgZvrb/UkPi2t7PlY0Yf2Bda7ct5npMSBO
cEiLxvC2y7ObkcLS/EhOhM6J624ESoPEPrDckqnhPx/djVZoNkH1QVn5uGm2iybH
yuQMFis+p5FgE6e+V4wUeIRpWGNSl5iA9itvl42ulb46bH9vBp+2joNVsSHFB5xN
DFcfoRR1NhZYU+zLjB+AD/Tdhj8IpYl6VYkw8j8m28J69FlqIe9PuRR/IxkaoGMK
r6KZTFoAL5tNb+Y7PELClatantZ4NO4Mc1WmNbhawrunythz5DyceOcCQnty1Vye
OIfOoI72/H4lgVTpWEoZ5RLW5/7dwKsb7C+BNdNiWAv3szcGrkRkk0e3DBi9TAqg
pYVIxSXvTA/dNderNW9xTOI18tYJtQlACbkN4oj9qPBwHFdS61DtRGMH+zO8wE52
X96LafhT2913qKXXa3woTP4euZBzv4yrItrD/QqCnKSTyXzEcEs4yMO7Byr2npPr
pGJlno59y2tt5X/t3+4wXPpClDSM1Z84Op0AL6fgtRSMYEj74W/jdy0lhtdWPJxF
PCdsESWz3SRJKMihKBTw3uEGw2WUDHS7kkwKeb7L1Zj9IJfLpIQs7xN42AMuMp58
WKI5iDIvc0EpNnx+bHvOAEHQZt4plaEgJn8dmG4TOwwJ44CN/1uAOXSp4G47Nj1V
Oy53JYpc/+NJkCAHjifu86V3DCco3rwegIS8PVMZ2nTz4a5ARDYCLKDMgbZyh9sx
c47ekknU3rd4dLAB+5RTov9FUcO8TTXPBPjKV5VAhOAOiHbIoIRg6aClXolvk4iu
ziGQS5EUXziDwTgWOjbB7lOsFyJHckz4Dtmu48FZUqlc7sbeqPoSUE2dOoysk5BW
uKhoTeNM8IU7dDv3ToDXWJQoXCAgrEFVpglza4XclWYDAqXRQbm9ZGdNLDr1dM6V
3dDapbfD3TvHGqN2Ty/mDrdXO8Z5rqyTBpEZYCAKgaBYGLmXuEUgUcsTjzSUQHVn
t+Lx5yqFQokKYHK0hj21Fj7mEACBvZMxgthQLt3IHTkQHhbb+qKQxwvXYZnPs4bK
GIB2Ind1NJiC9UsGmpQjXXMjj9gwy5uYZMBnlf/cXte/D4WiyM7J8Kw6mkolGGYF
GZPoUR44itQg0VpDQe8/E16B/Jnfd13GF4o1GAXhhdIyOYAweMYNWodksz+ny8xV
HD/FiInEAHau0Js6kKKOypuNwqPL8oP39kgNiBTpYujPUoHO44HheOSuGhwWQM2v
Cp18acZ0xs9lLzzJq/kKeAaJ+CfdVdmFIBs2ZGm9BiuhakmiTA9u4MpcyrV5fRbH
`pragma protect end_protected
