// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
x3X/fP88JNj2f7rUrXJQ9QwP8XbxphCggXg/OsUx0wHBfIw+I1stPyahkIhV
SyFeE9Nw8wgb0uRr1NJdGhQqjESKAageWT4LRJbnx2T/Ecp9Z4fFvkkNnPDE
PJ6SmrSpYx+NKkpDlb3n0twC32+imULUtjVERf6xNAo9D5rE6Lcaempv4MTD
1llTwaM1HpYVIHfjnvxfzm/5RtLV1gj/jdTT3SAxPePNrgvMdFpRFjWq0cjq
ZMkwvnba40yYzk4kbGanO1uMUzwnm+SgVi6lOhiPMTNLCyI47+N88zVfB5W4
GiAcCEk18yHc+4LW8UMQPi9BAbtavRBpEfPKNGr6NQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
az4YYJHm2hL9KKKEhspWMbpAYI1c521c8sdEBoG/qtXBSJNJQVAh8QKnM5d/
kgx3vaRd5+Vwo80cLJ1Zi9uDUQ5JGhz0qlOwymlFa3jZfW5ziAi7ucfEBKMn
oGCLgCk1th+9TlLwR68rhB6YpXHaOCKfeprgRLuohp+60DB6Xn3+v2y8exXd
LUMhSUvWVQXAl7ffsMc8Jsrv7iPc8R2N5Kuq3O+Uu2VuHw070I5pTHeUEQVn
umyohI+goFiWLqRoDaX38HsOfaKtQUHcd5pGCl/+hW/6s2hMw2Djp/B8FbLA
CxWo3eSSwW+z58rKp47I5jHkX0wFIN9AV9GUw/M6dA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ljsh8NQOa6NzwdlTn6FTLnuEweBpSsRdO38wxsTrk5c9/iFJ45g1ozv+SnDl
j3zVQQ7RxfsZimvRnh3ZJ289EOYvPK9yUke+GEaRRpYe4OWOFxSVX5SU/ZTi
s3sTnoDplOSP6mT7VGBb9d9yX9l7n6oLBLGyqUNH4XntAZiGXmbk7JYM04ql
TZj2XqWcmZHrY6rYZ1fEHzoDTuwI4LO8NA4HzNJ4p0l19d2MkcPoWm2YpBnu
j8rSmFr/OB7U1A72i92GQjWGo1Ow70H3eTSPhWqQXakl0Inzv6BP69UBK/dV
7niUW+fqMSl3fnl/y66aYbdd/vQ7hNV6zUYUQHRJug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sTdfZZf1FrAipnKaGudt+/FGJlpjg3cn0YVnsCGDqOrodcYMEYFzVTzJTRSA
D69rm/igX62UTI2CvtpwErl5Z3sFO0NwanhQF0EiG7C1+5F0mpSnFlvPphP7
PjfDmImUs+snRZ5xj89ObT+4DMvZ4i3T6WvOktpIktflJdo3oPQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Se320FPiaRo4dEcnNdfPbabjerm30LnpbjliyAxtMUaTEFoTEPpUXiqGN3FZ
pPMIarhVerSZbzYhhN40aW011FK9OEgiHHsRskS3ak2OHlsNmpTHTH/CKti/
Hj0FKmjJdsfhaY5rJhC8Pg84SdZTDwZgWB6CxvCuDSU1lkmcF74Dld1ViyQQ
gE5Xqi3OZIMcOuklgklqh5m2FQLy8DlWP+tDb0VeS1B/LXEzePy5ZgiPL6cn
brDaE551CJbUnSpJHb3Zj6vFBZnQjwrifdpnKr/xtLeOLYdQEG0s3LCRsrlx
5HeUqxq8NjJywa/yWUhkLKjk38LJCuA8n5msWlrTsalVr7LTb3G4V70xmQOi
YOAuHlIEvRy6c67wJ2aVSZUFI0TS9vCyaKbKclr1Z6SjBR42yq6S7Qe2EYQ/
vhhGY+/NDQmY1vHYbbADas6bCw0N3Q9LmWOcwc4EboI8QD9cbhTLo1u2iXvU
8c2cV4OC/sZ/nsW8OPWoCZvX9dW2KCcN


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gx2fLVg48wvb2fdl8QzodpILTrgoKYVT7JRNUr7GF55sj63SFNfJIzwXhb5b
5XAgCvcJ8XnrQHBn0TluKE5BMpWwdUzxjTBDLjxuF79gxlUn98WFZUh04agr
GwDksv5VHsRH5ejBb1uF1MzAllWAV9d5NU5v9pF2w+4a9wGy0kE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JsCvKuoI3N0Q1+HV0jlnJqv7z1wZryVuhzE40JREq/5YPbNVRZITAKDqp+jP
upDauqyAsEggdfTQemjS0u82MwazZM2IkTR/K1ATA7FY4e0zW6kqeFJcSK7k
gXzBk0cFsF2cH3IJenrFkWMSbyYmaTGrVz+VfmsijxX0h6FL2vU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 79776)
`pragma protect data_block
bGlIeJlQJu5MUQBkSamX1kI0fz4l3eBcmXDvCdxHbcghxBfmBBDZ0ZH97a9c
0eIsErP8m4SjQNmMIq45FxHu0YpEWvqjbr2pE8vawS67zrgva4x+om2AnMih
zYMDosZEtXvlbQ7mmAKtcZ9F1hSXp50BBW0+lRFwfqctgNjb1k1tM5g/wA3g
PydvOUFXi8wJNXD2af2KUHvb5vaAUJiDoC2jZjZdA8whK4HiyCVb+Lo7lfRC
YzPBWDrMQn4nL/UBkD4zcxJwQSlvcFaWx+wZQG2B7DUwSQn0+lGZUrdzsEs3
227Lhk3GUdxPGOsRR9+0HS/gZkP1laOByXB1y0PXgA2jHo7jyd4nmxs+wP4u
x9uK9N9A7cjEEJznKos1dY+c4Vp3Htisf18/w7F+pyFEznHL4g3QH7018aaz
mQG59fZxR+ePgSViNGPSYY3O3ycaZycArPca//7j/DGtupq6eKpCaxCkMnUl
Z07VRt0iqEGjMdHNmd8hMILi9qE2O9YJm5g001jZ28/ELcv1IHq5H3Rg62up
Gvw3A+eEyc2SaqFD5kvZnFjOSYVrG2eN3ZvslVok5d3sfho1n23SzhKPMar7
juer/tceb0sx6adUYgXsIujAY1io6/dJUi4pJc/+q/vgeTVW/OnN80+oFw1H
LEL+k0grvn8XiyVIN74iR2uX48ospFIxRoX9bP2B2dBk5W4cCZnUIkFWLGr4
B3Tu+1YKCdL+YSNXSB9EjruRi6xWtTCrUceLot5/6WjXC8BcPO2iERki6U5x
jj5mzonTmbA1KBl7Sn+CzH4g3AUkMzurUzbLCwDxMd7txgrze0u/0xoS3QGp
oJZbRhgT/wDlZAw22TkPk6iHJC9fRE3J95IuDx2lT8PjnEkLzE3xkg9VLJed
l4zE72gOD9GVbUY/GeSp0p2xdXp7GsTA6873DLrTJ3DeNvk5W2/+izrZbatw
Ox3Qmu2CNkZus4DqRkVKL4n1lZPp+petb4RQsltb1Can99OaaCvXtt38nVP+
EvCxFd4+0aAdaNLap5Wnr7JLWNnkg4Ud+EDIDUBhn1vv5Gh5GY8ebzqeWhpy
AZ+Cc/SRdU6/KtW3VtST3r4NaDsBCc6D+4KGiVOTiqhEEXxk7g5/aI9Hspfk
CZyT34zj/C+p5jlllO1huIgVnmaDQQnzQrAjy0F2Odm+Wz2DoX8RHHMmVs6R
1lUPG2lPnUtPdWEYhenXOH1nRznQ/J9MDRqYfJP9u1HIXcxIb9Wk+Kzb2WLX
UVSgVCAg5n9LurUIyv/3Dt6puWPVJxGR33dIDTxGSJNQxBNAJw0yM1rVfRc6
fLL8+UZxCnNCzZFAa6fIyoGvnDzR5XpgVFuN38vRnoFChrD7unWUCx76qAYC
+lSmzrGL/fsvpu3s0Slas1jLxSsTw602JAt+ohIJkr8WVIvsPmPTPdZXD/z+
QmRrfZtSdD3lN4pAt8Gz2ZtknQbFbOfqdXOXdWebt/5c37sD1IQc1+Go4bGY
9TxJCKxnPyxNQQ6QqYl+vIQuImdKkr6jPLEu2dhOg4mkfsAzBuAaRCmIbLZ8
UOl8sTplV3xk2wSEisKw7Pcty3yBLI2r/kNBfubz73Cm53PiuGrPmeTYmLJm
gY12n67T6+XhEHbe1ZknAIt25CmUzipvmB0DK5/mDyOlCJBmiEeBmlJ0M7Z1
Qg3RjsARP8Bzmd7jWqnGd/06Sv3MQ3AxRMjQ3LtYAHb4F4sKqC3IsIZTf8jM
T0tbtF7wkwmQhZDoQu9JTKohKCwq+Y2yuNR9XheX1wBCiCYKLy/rdkvuBhtY
w9sDuqepCK7fyUpjObp3ulZmdz2en1gegUcZBGj2bcWJHOB0hAQ3j3jlAt8N
d4Ruxv6qVURQHq5buMWEbbjlPPgJZjCO8+f4qDVScSvPHqtJjn1BVvLkPabr
jPdyTjvQFH0HM5wLNBLG0v9KJoPW/PkLebT19RcdLajMNj01/RSKRstVae+J
jwTaU+Omhjx3CKvwDcz+YoeV3DUWZF/qnhaQggppYh0EpJIANv+ib53xPT/n
0U+4WaTwlMiU2D00bh1kw+vdoypQ+iexVYNlsHMXnW4GBIrGTrJffk2z6c8h
aIHog9VUWOBcCjCxczRdyLp4VqLcin4uI4dpk6pjwEiMDfS35ikWbcZUl1Hh
fDcBNweR2nL3n5tWh99OD5q6EcSHxEGBPvpbMa8Lx6QRoC1q2hg/pLe/Y+xL
DFUMJqEqzYr/9exQcCw1oDNeuOima5qV1Y/aNZS1/sW9AwpRYOoMTk3dVIJ8
FBqaUKlrD0fbzqSYAQgrzwkWy2kvKXA708AQO4lQlni0VOM/bQSdbMpR+OgM
86ZHXAXbhKDyxwPxAm28djrn66pmfWPXJDaFSvZtuVf5mQjM3mADM8MWaHKz
fWL7eFKPx1U43fOC6U9dzudnnhdv/IQvLO48fKM6g/qJwYYJmHDO/vpw7KZ5
rBGGwATceNhKpjTzC2V7bIRE4cThvRRxsQ+KhR3bgOSRrhoc+tE7+8ugyN5k
rbr30O7k6+kXw0+jDlq5CIMnAhWx7E+DLhzz7UXcVf4GRmsXBd7ph1x8tgCB
aWmjEi69w7P0wmcZLIdGlS6ngO6Mf5RU7esDeF+0tld/9KwH+DUKg4YJ+1RM
XGBB6U1QdEUCFSzmubE17JsVQltJKHHhtL2fXoPy7CkRj2Iqm6W6TX6Mmnpy
eaTX1kk289bVmhxdsqqpUBY7HDyL16I8MGEeR/m8/sM4mqwIxH0pNVdKpe0n
/4ixeirsTj2LrgvZY2VwrQBHDPhNFAy7dRjLfcOnLELTgeA96B81IMVPWVP5
7WXUbnq36FIwwuhzbebE8HgtEFRUEHfmpBCfJ8p7YrMslFhnKDEXnmESvi2r
56LXR6ACD8eOUtn1bY8XmbJbA0sv5DfcOFOthb885Ig/jY8RPgvywszPWZv0
pt3y464UmWKG58igHx8zcOR2plsDeW6E4pNGAMQm/+qHDLAHH758Y97U51zm
hTrKstbP/9uMKA8FhE2TA//38bQC8mZa1ZQz52vdqsq9EBR7uRvgVsqvhqrZ
7A+ncbUxH45nOSVZdTW90e3IN8nbCAGbkYB56AvZP4FA9Aw7EohIkJ0Zhdcc
F0OvQJu51YDXEgrsxyn0IAxrm+FbmuGPagUrv0NpghQF/EdF3bVszEqiTV1O
AkVIMPPxezFutmWGUR2SzJyDd8rzfHh6KxF++V6ZXNozMBUsmElY6ZdkiCEb
VcFhcC5lFwH9HWh0kIWkrNyrWkejhTd7NNIMSTQOX95g3rqIqIuCzjSEyqlz
s2unxnPW/04xUrdAr241edUHavqkh6vDbvd7MCx2KRBLDjV7HW2iZeWn255I
9uNq4xmwLVNsUFi+e1t8EBTo6yZe3gC/qqzQSLpu/wCZQRNcT3olgRSzkZpq
N3f/uUjyY8AKkWGs+CCGzhD4hUpgW3anOb3Ae/1aEOnDpg99hQvJXB3y4GI0
uNT7X5bOVKBocjLZqxBHDderrnRQRhiufkAJP9Ra9bpkiDjdQKB2ua0Ybk5W
7PKEzyvJhVbHfOUCYZZnu8RN5ETNn2QuVpcos+qEzKYaQz/ivYfY38vVyW9B
QhspzLiWe3/a0jTl2Lza4ePvoXwDraP8ULiGLE9zWdoZmArP3KyUzEXhafaQ
eAI4gnDbgex1xGGqr/vToNeA1gn3GZZu+AYYu0HGF0ty3AyKgplcK25wcAoe
nCo5UasvwurNuVcrglU3AY2SUW+fGHqxrE5/dNJ7Qu9aPDXWrwU+cf3jcMR5
xLHkhtOfEdbSNH6BgUYnkGbmlp6khMC0pFXJt0XIsFvokCgkuMePEH4ks53u
RcN0uiaAqr6nR8dvgH5ap8NRUByklTCN7UW3NQcW4N0JowfBNHn8IHiOzALJ
W4XN3KlyxJw5ho+qBpe3JRJDiukj25OyjKIICyk3qiS/gMGXp5ODlo+OjtRv
j/HTQIqRb+RDZZkwtTV1EMP4syfhap9SRmkvyOKxDawYnnlyxYqpxMGt0veR
rx5oclZbsRjppFY9/g4R1vQZmAlawO186bGMN9O3bO8J4gEi/OdtlrPjw0iH
70bBzZY9T/6P7r8NhduM9/8Psk9n9M+oVJZLK5pSk8qKQx8GMx3joMI060Ow
XLXV6yEUGxBrgtTV0XXPTFDxShyAxYQvJtwpL48A9RLOyOzBBaBvqFLXkmTL
zkJ+oiQ9XaRKNlInFC6Y/GBUoIJcCctiY5tQrtQb3vFHvdvL+/dIBC7mkqQ+
EU5jKN68RZoTQF+gD0MAt8RHF4v7CYb+/cd17MIQPnmDXc4qcAbD7ajGsNCn
ELbRh7yPCBi+iMsdbsoocGi1tlEsvisq/6+77vkgtZHB2xqmIhXBYl3cUPuJ
idACD7peN5arA0fUTo/gysoeC3QN4WpWPeAvTMbfxxsABLnaDhPVstQdS6zt
noWxGJxyJqU60GEhiBRkfkRhnfJRa4/VmhEOGhtIbgD7INVodOXNvg5FCyLZ
2dxWq+yBkGZ9MRbLW4D5oaHdA1hRW/CZ1KX1+PrnaPfYmgq2HcFvsQuCXCna
0g4ByETXA7bBl+CGM1sEJYbh/+O/CapvoZA5nygD1TE/7tty25LaydpekVnS
amCCT104oe+heedYxPZpDluXEpG28Z1yJvMvenJ32EZw9GI+PKMZF2LAMlf5
h3RE/aT7Q+GZ3Jp6kfbFsb/N7+5stwWBKRrrqexcLwUTQuPhxtFviHgWFdmH
kz3rkdmb/SAphpVY/pQYoPaaQjx5CQS60wJnRYX38VMIh3W9OejsOSYknJ31
nW3GMRDczO/oxemdTlZfd6wW6E740kqSUMvmVXYwSoAyFK8ZDtrFhlj1lBh+
hjoYU5/CpLDzAVKq0BW8fvbscSTe01jad1lwmMB/DkB3q3yKgitLvWYoK8uQ
xl/qlsFkFB5qI66a0rJsuO2BWswbcLloVSonr6geZlQYLHaSXrAL9pYNZhoi
kLtYCIzkG+5TYHEwIzBtoFUanyv8LKx8xL5WgdKCvbRKDpRjepNx8FPRiU+P
9/4Eqi6ob9vt05wnpqtgLyPXXc35mI1ELl/y5y49AW3JDpW9R+Lg/LXyVqho
3IOHhv/KNHF6pHhVhrh8OJaaoJMQwuwBq2Q1v+R7Kb5NGPAI/9UsO+QKUQ8q
cx2wBlCPxz9jTq8GqTE+T4wz1OhgOkkTYKCuB6grlkM6TRMVCp6I6lymq3FG
sw7BCuYzRxnIHMgwRKdNn/XKInsZNskJCtMCxM1FMctSOlBedqSAywvg+JyY
nRyBLxEcIweL8tS32To3HuZnpyFkTSPnTLbUP0Q9BOlvAG1Xi90AxIxqVvWS
9cPC+ViVY4FomGOJsHMeXvdoKeBfzATp7jp5ejNaDCkJ/QRXhLLSwuBo9ISt
2C0sHAukt0lgfudWh2iG/d2I/ESGjEUNYo+q7K5osEBuJrHBjElh5i4nfihE
CH/p/i+1yAFUuvsUOQ6e4YWcILCP+Vb2UP0UNViKovppbcfCJg12YeTxkWM3
Jdi/elOtWrQifeBXFk4ME4PyO5fbaMZtHGhADFG0rqYBaaJrRtWt7waHqoq0
HVD2uYzQRjLB8iQxRWdyN2vTLyOapAo1iz4z0zI48F8rXLCuY7bsOdbv7Cmw
Grdab2kcKwzlPyo3VHm1/36HHMfQWrslTIVp7Io8gj1fz7NB40NdCB4bUPsv
3hBowFQlACy1Zu71keEXz4yj0O0lILYX46co8BNbHg8gkD5E6erMWQk7opXe
QYvtqfs0UmFiveh0RxihKgaDXt//GQc5VrSq9R7eGUXT3xB0sbMdVQrcw44b
Fn++60RqZOkZFklntEeQE+f+LjDzuvo8kmVFieIm8uSBgnSgZslaBGaGzcfZ
IaAJyIC4zcyE4tJPamjLIe+0d3B49bKzsgebguYCX15JuUHNXnGomoRs5irG
Zc19rEIbQrYKwZnHGAqzjp/Cau3mlCN7SO6h7XofiY/edAe5xeTUP4efGmGL
ANYquJil1yQ7xZtnxXRXucK+0MP2rmJxcGDEfN37UFMMDhmHxUQPG69ifJle
Un476YiGN2uHwJp7HzddB5yZiSXJzvTYzKf9otyz5Ak/LptAq/YsX1WjhqSp
txq3sb1aUTPk0wiszsFMuQ5GJOuPjFeV07DV2jy7rD0HI+CywkRXyDu49bc9
/QqHbNjupsCn4AzMxejnZLujdLTYadTc0YTEdajC28hGJZP5QQ7QdWu3TgwI
ZcWUPuf6skpLrwUWFD30H5knR5CHWStfKHp7dOE/qtHty8Ms4MPdoeFKtheo
qZAS+nyLG4cxVDfixFkLWcsbfsMIWmokW2IuWGZvzX3/09RewO8OThI+eIJ/
flalu3lApq40GM+okZoWYW2y/816HqM5H0LoayjgzwsUrCoYyUqJOGs0mUYb
VSAgvFeA7AtGXLO4dzx3KtwTgacH5QC6aDxH6ogLh0NiydqQE+FLFM6qWQJh
WxLFP6+7Ca4J+mGlxN3in9xfIGYV1gboUcnzEoB9FW0cdY0jgO3nsR1w/Gls
mwFFiFBFmxbp6MSJnzPux5koxD134Qesou+92WjKHX9GTZPV7NCDo8IKXQiu
mMYUpvKSh2yDbw8Omh6K1CbFZiF2SZW/ls5O8hHMlZN+xBP5xTZQSmdrbSFR
8n3QIdp0fuPq8tAZm+4B3kYWdgT/AJ5zBKDFR8cS6/ap9IAcV5rj/HasL19X
JI8AJHIdfHnmcHW2Ld93j2QQ4Cuve5wcvImjUpplpJ5Nj5iH7VBIbjEEkveT
uh8l9WsPKBRuAvcO9/qaMn16UjeNlhfegCENJ2cOCuzDw85mpKTZXTN8TQ9x
qVntHrk19P69ZaHKkwrWxY0NZJcLizE9ceaeZivPKA+Pj+MRJWFAmalM1GA1
BbRDcXhB2PWIoxSW9eYigEMvO8OjQmoEGGFEIQPEW3sSyL9krF/NYK4W3xot
etntlEWWMyxEioyvSZPdhVMXhWzGTtF1zl6YB3PjGZBwC1x56Hrwts1zQ84X
RQVAZtuA06iIGkuEsRxwkgnu6QmXU2iu3ESiHWvRoLdiZ4cprqQyT9R3IelJ
L3rdlSOxv8xwhUrFj6LMrg8B7ztKEPobZIpf/9MKr6Ojt6BxeyL1kDtbIc+W
RgbH99qca6xa+7zNL4ALrS+ZLdRqwRSlFvCK6fSgNbB+JLJC5SfRjTdtY0S5
XV31xfad75CxV4lOCrMNVAWn9+DmK2g3eCiXbJQoPj5GZNkzHYFx7GT+Xm7S
deFVeYvlrDHGGsthbmzoW8s+zngzUBeFvtszDJMoXp0D6EEvWOlLLDVdzHgC
Mo7J8WZ2aKFqTNIZ1EQlxlWcXmu4Xkg/gcM04pWCNAx9pvjmr2fAO9DsuQU4
gYydusvhOUFfrKVQxQQB1XYKk6dkvHsX9FxOujR+VShKcpMtNV4JUC4V6qbw
6lagJHz7nWUjlM/+DSHZiO1hOc3ku32tUbNYDS4rBUjXiAcivuU6PxAZnDAa
zdcJAQ3DCnwlVK0jdHySlFPMtxMyQ7wvBhTcdktgcYBm4hwh9P+mIKJjPpHr
TeDBzL8DoycdlfnRPRAVqF8amk/jDo8M7Dyrlk+blEOOpbp+Skd//XZj56yA
SWZGPX4+bPKqpNPXqaC7SNgbaAjiuTtd0OIr9CtJFYcnoNp5u4IUh6C9lMAD
72tL8hxm8kLlL+vIF+7iWuvdSRrueFYr4yeJMNq3P1wYG93gZfw+2KwBG6vc
hqNMLKzC1yuKoXdMe5cCl/sYJGj7PQbPC6pXNYVa6UCh7PqkXQS21ScRmBZe
tnbdn0xzzgbd3E8nPmNkm4j7fHtikrQ4gKNXDFxJaOpEektxLtEgZwQbwco6
5Yr2B56LNzY1/HfhZW7a5N70mP70QEn9HtX8LzILrq2Q6kJyzZAcUFS03t9m
3g+LQssTfEX5a3SEBTWnOOPqvzuYoVzeaKs/kR+LFWGnVfwf3Cn33BFrYRrT
iaRlBn2nUQXeWJl6rkwkbPRqZ4uLo9HGDs4ASw/uKEcnCetN1Xel/aOaC9dn
vuNM9sts2mwq5x54ip9td4AX1g+FvNkWh0SOsy5pYmZjnG4S/XK9uEWgIpNe
YDYc+y7wbPwlNGNcInGqWr2cmMBM6SC2u+iUzG14b4S/9I82pjNccnZ0zNp9
LYx2e78MZgjnx7iHQHFkTWNmpoEJ2zMK143+J0WFj8HRfXeAQ7U9HMugpopC
WFVZDxAMDpK6l4sILryoVuAeQ2Ma6eBrPrw8lPkChaMWcUxG6uJPMOr0lUi/
OJxHLHmQeiaVqG28bvNDcbHB06xyKH42MOBxy9AyE9RMqVBdQfmswyTdI0sK
gSDnmHxqx7C+PTTu2AizXZvMpNY8tLvI8Pz2CJ4My0u4c0DpZ7wJUoVVDWjq
+TQpoDQVEnbZw/Df6W87SkqROBd+IK2iQ5BwSyLroW7er5M0EsLG7NA7K4O1
rvyVlaF+NfySXBZxYdHjVqhApOzc6EAJP5BazV4wFGOo/LUIrolpBLop5Bsi
nE+HnpOcKHtirJV7lswtZkn/4J1U3sJK9dmzsvcmRLdlfjDHL7fNyhG4PLqi
mTIhGT0GIU3s6vSRg0Wa1HTlKqv0x2Gj/CXvZHiRoQ++1Mm1FRzanu/F0d8J
gdGrEb5FqAzIP0s6A3vwU0yyoPeCzKR/qwb5Ob8BCBiVvhj2IJvRV7jhI/DO
Bk4/maVufyaZcyQZ9BlwVcVSo25oy8x5pgMhgP7TErSsHPeNWo3OWgxW4KNq
EF2VbotK/VHvgd6NzgEM4wvgfhf0o9tqyhg31XLUJHs5CPxH4EcMFXpkcbBU
4AY66OuTiLzi08gFJbsNgTB9NOc0WJMSE4mwceCkLfWtCNuczoUb9XoBIG5g
ih3Vxe/NalrPxJGMEz6rwA/oJUZ3yJH0stUHYoaIhl8n9bSRp8GSz5XH73PJ
eKKRhBTRtqTuKBXCM/GLhlvLOXAHUzv2jretxl7pWAli9lZxBxrCGyMv7VpJ
4m96/uvIz6D0Hab3XAKmSXvWELVK0ZAttS1ABwyrXmX65NKvmlWtwW91UrYw
Mq/1ime2yo1D2L+/W2E0aN9WAw6GE53xmcLyz2CQmNJcMpGrboUCJZNlUt4G
9AWliFH1763Q/fMBiJcwI4JPpcehO/9EMWsosjWnqcKV4MHjMicM8QgRfbge
4grR8W8cvEoQTTRsWX/cR4TOlR6alzRectrgf2BsLn1DnAex76sbHo61ekhw
rsbyjiuu6CzZPjX8GtkO13dr9Cpo2yyyXT0Kr0aV3xIq6nCK8425C2yYhfZK
YngLFI3Pj9LTRvrbA+nSsinVs71bX+OvdjyaJS+woqqYV4aupxBddLJZfRX7
GMDjEvvmMISrr/yga3O0n3oCD9IsIZDn61zsbY9CHVd6K/DLHiZLFxVZocCG
7wramk/1VSCCvvpeZYNU6XmElHyLqmNDGka6WAuI/ZXr5Efp3s21bp4visw7
ka3jwW9ZYBWA2vWnWJoIsPgZY6mq2NUL2e5ZcZHqmB4ZXNZ7M4+kmBZk87ld
JPaRDe+Mw4HKaauzAVjVgd38mH2WbhHx/gSvIgpqQgE+fEzBhyR35705fQWc
GEKJhXe0LHdpalOZUEmwsbEEetA0iD7TkfOB0zd9fOp0A1AOwnVMA9/FYWHG
Ecd25tSOVzcgtBsziZzGuAmKypGt/YDoSdfZG1x5O7R5xfp2LvrgDsd6cduS
WoMbfHxy4YKtDDmg1J/650xo1kKXdP16fpytUBFFj9DudQDDWyWlzMVd4Z62
/p6smT1brdyerXXHZsgfVbYqUwsen3NRFuFsXhcZrY0YkPb+u+1gum6NwFvy
akbaFX8yUJTvmPYIiqVQeVLxJMPRdjnS+TvfeZmNCVoJWhCQkh6XvY2Jxm+E
KZIDXmaZdNS5/c1iFJYvEzT7O/BXuOVAFnSAySYJutp0T/RXEYrfDhUJvaBM
1h/Z5ppuvYiam122bWZQhy16ZHGSpMpxNrfx4z9FoAinX830xsfnPlqw6imL
twuSM4wLYithXymb9i+itfArhrYW/OdG/luD+tqGTNAN4jvB7mJNQDL7jRbe
qwVqhCMx+2o8LgaA7Y6rNtcZ8JLT2442LhBLNnbF1I2sYY+tFr/3DWuKuloZ
TtfzNNk5z8MEQHWfQygSnjscrq+DNdJNzBobxb6X8mFHJ0Mg1V0D+giOrSjw
gSeFgIOsPOIkqP7eRjVbx5zllrAze44fN+YDub1r4IbH22fiB7CWNqqZ+2NE
HNNyZ4SzEfHJEKnmsiKwY2ZWC2QMb8wihjHozzRYuSIjwqTUO9M4zzzjEQKK
fLF2GlwWynHbQRhWTSV8kb2N858e/8oIrVW8zrU85QHP+yQC2LAyZ3a4RxrK
mfB89j263kuLE67/hOXBNMpOSlfF8WtN2PpQZwVt2yrKXGaUGkpYXrJrClBV
b4BFxcxTmxffS2CQr8fiH2oRUMaReHBLDrT5n2uwvqArz0/Elnl9IcJwkMaV
hxX/LrmmKLqE0QEmMs4bix9m2snjTqLimptncV2QrPohU1f2gRMt7zb5A6AG
oIQ09Xn7Y5fbNSBB4lPOr5edKspD0mYwBebLTAd/tZ+p3bOat5BF0gc+Mv2Z
cX2E/s3/nYSOfnlcNgvKzeeDimOMe1eKyupcDr+hPt58H6wrKoqlciqZscNo
SlsGPUY/LAjEtFbB2SO4YPuxHV+qJWhiYz6QBjujUB+EMAjcasjJdE25HZ+c
Y2RWDKaW6IUOeiCHwlIEWvpeGJCJMoLu0Jk6A9heVy26Wx2FF4tNvpw6stz5
9KyBYgOb+QJxAbu0AXhPa0NAl2pz1IzZUL3rMtSLRlUUbkHttW3lzwslgQUp
uehXcPxEtBrYiVw6piCP56BBE2dv27r5AXfRYNFgawKUabeGi9Giz/kHcjfC
UMT+dwWTTgDBJ+ZeAVjjfl9gCZr4jppEPB1FuU37zf5k/cC6NTVeJhHa0liQ
WIIVnfOf34D5K/fCmo2UDGIlcJ9EKtla8R0v2+zbv49GoITm6JUyoALyRc7K
efYUIY3/5JnUy7JeDXIk5zer5I3gDlve61wdMxAU5mHIFY6zfUi3519rScAt
pMIMaK11nkZmSIJqTGAWWPVbHLtRJ+HaNBy5CqjnIVZ6Wqceb6mD+ZjVsOVT
mP0XDdBi8QM4IzRL+MXoCQBREM1j1caFAuuUB7uE9jPZHLzSRuzenpALVaDW
tMFAM7ILzSKKHaDKVMQ8cZRvOjCSlHt8N3Xj4X2Qqvp1EqYGp949U0mprbLJ
2TUGT0G6DXOE9PEEKk8O7bmUplLXs4isEJadj7aWI1XoltkX7/B5mSc9htno
+5wPtiqkLYIUDXm1kDrTU0d3E8ex/2eSBaSnjVuL2B8AOii69XFhBb2R9My2
GrzSoILZpLgu5iZArwGVAK8UCSvKAqTuS5KTJ61GSJHg4Tn/LpL3H//EdFdp
HRFsRw32zOZ1cFoPOJPukD8mFAxcQfXUpk3soIF+DZ1AmhCbrPZZghJHcGsA
UBDN8GvFEteL8Ny4rvMJv2UeVXx5OwEkaU2lKtpFP2ysLdTGpTm5eXBT19Nt
oku1uxCivQ9fAWaNTWFaS0NVsGNV/Bh+axMxcpkmQsG9i2SYf+NaDeM1C8Y8
3l6e2wyT5bwfwSRh6VIwcfaYdlfETa01763q77+FaWKqFcIQ5VIdq4JFH/C9
s20hT4SdoKuC8XPGDrpi3GkNqgCeeiVQoBgwjiviHLXpoQfv/8iUeFbYekyt
imDhjV8PnraaTAbsGwQ1tYErNbudrb7CPH1tUXULqirEZrmZzGrNxEl6MQgd
J8rZkjnnkh4tD2pNVu+IHyP4wIV3OIdTf7mAezukJY2AVhL12AwkvbKdk6Zx
9JYTboLn2A+grRjiT6+CXm3HW3iEUxs6T5RsmM5DRckPxmM4O9q01m9o1Gs5
mvwNXFlxkBNscP2jE/IQEmVRQpd1a2+MGuo4nhYvuZhcPLpUFAf3ZaHHaqDc
+wBS5nO6xqDnANYFbVg2OLW/nEgkwFSnOyfDywVLry8Gx7h8Jk+emgpGgmSp
kWN2w6mArjruhKbE8JFvgM9UF1CnKrygKIOXJR+dZfjtezK7RDbMMXWf8+vn
5AgnMN7Fm+YDmKuFfYWqNXDak8YGuq94Qu6aDecYEtc5qyxatY+5ZYmLjB59
nPGD3uKbCtcVWLfJUpmTzNqTAPXUxCGgnVxmKvCKK7lYKVYbkqIlBOwcAFBK
Y0WW7hyDop1hF3slSLMT8HUYNnBrZegwW25KAcYRdbyhcj5fRrMKZkyCSTdG
ADFG5FLU33zj8n2D5prZFRX3LmFpasZ49c/vt+E68Uf7c3KmkOnNTh2BFhuP
Uz62us+Lyd6/XtjM2w8gvABsTEO4ctbfTXzIQyadJqN4wdICtmbiAxA+Jv2f
XQoqCDkmsP5CnE2fAXMOxqnquWUAs59GQki0HJ5IF5M/wjIEDIU6srIv/0z1
BgVAJTi9eHZcHa0+2SCaVMAU4ugJxMYn8L0hfFEyIt6gdJmLuY53eysCKDoa
2AgefyQ9h65+CDsryv5V6ZaHDDT4a2UnIzpVJN8jg7U906o/HAmaJw9WhdCT
sIuTwwCvAYWS7qRfzmvrnCEcTFLu1/vvHF2nxuYvbfvbgZe2S58r9v35BNoa
d4fwPaezYuOw2vYjkYinhIcClUSdKhQVoJvVL5l9mee0Y5lW9fVKgLO0Zy76
6//QgS6iIWCFchlbL3HaXoVTlHpRghVVyV4E3F9JHcisVmwfQAE+d5ZR61e4
mmWu8cRzMt8lKoAGuZbsey8qXogelcdDxuK4DbVYFWvj73Pkevr5adgQpI4f
Dj0ytOWMzZMaOq7KQxbf0bkf2zKbgPEHyORjI3GI5LV2CLzVU6UBKPXu/803
AwTiHBdgaUVTx1H626+TnAI+3FdJCVI83E8Jg+ZhXhdharRq6uermGA3Z0ZQ
2yK6+Q9LDty5IyjCrLSDsqSpd4T8V3QUQDUbSKUXaOtvLfMg4QpTTMios0rB
FhXtHL2NTp6wwgd7oMbtclpjIR+qWRm6KhhaPHQXM2+rL0mQP1SOanVrM0Va
x9F9S61egOdn5QJU6s+3lxGmh+w/YSpyi6krPxhaR4ldwV9pp6slLi/atHr/
OK7RDhSLGAXvEhQbAbI57+aHe7Wc57lRUmllRGu83r6lQAqzqy1mEEetAFcF
ZJqD5Kf9E/9uDw1/37uJ4ZmOyKuCB+sAf1FPBrVWdlyvrQZISLvJoE+cG5qH
igshvW6Sf20rbJgXVp9bBFJzXqcUuA09mE4yItGIc6CcWSKA67GFKUoWFe6b
yZdS8LUzzfA5wsaLR1IVZgqA0X75cJ4wiu8ns+phdk/8aEIiisCVCmapKIoo
RTcD8AHx/+jYQgnLHTxtX+xEkVB6VSySoEyKMRZJbyOilvh0TAeFIKH/CSqK
b8WAp0qR8SlOSEM+3GduR9zEsS+UE2d9eYgP8cMdAz3BkUW2e0ei2EtKePvd
kVERfE24lcH2FdsMND0TtoKu6fKPOi9QfgzXI5u+aFEeyfSb8ASNeJLFUAQP
6N9dF9xaATID+wjCzCziKks7gT0wJDQjy2VGh4RSOrpdK/aibQnFGBRgPdV4
rmF893Yhxd91D6IytKB9ItTEZ32+46bQwTtS6S8rqI9JVzDa+wSZUGaHRNI7
ld76VSr5HEpKlqfdY2XA3ae3jqtBIP5mTVYHBdYS1ItclQaeTxzhpZQPDuLn
R+yF6Q+/WXXC6UL6mn4cfG5JtRZxPT5HluZlvhjzuxx9lSPxaaNAUeM6XlTe
sOMubAJE0+pvs2DeykiqMrpGmCDt8SPFHav4cCUKfvcZ+g15xI5hpC5nE1pt
mWcFXT1tdf5+vd90CAW1butahLuQObqL/WFsQUip03a7yYNU5TfE3Ge1XdK2
m08zH6Be9AajWKW2qEXTHrWu2VXufPnslhDT0vJTOESIh+h8zmss6nQt8s/9
qXfLjBkC7L503wWBXtrLMjvarV+tupf1iKU2kUq6VD1ZwpPSymRYLw8kgsnV
FdOhJge5D4prisAtUiWXlnisX6LODm00VaXZ9VrTr2BfhRg9ZVdcUVcl7PAl
2ZAXzl1pB6QjnvNTStuVKBg5RNZdiI5UzPkd3KGXh4kJiAKxQBAC9ouDW6vq
OGpDvOfN4iY7h+ZwNQus/d7IqheoO/edD6VN57bz3+gXEPxaMYZww7spBjh1
MYd7Nd6iyI3y0d+DG+erJ4gDhvlebRVbR6BKAhDfBmg2+QtRuUjILZBAXs/r
/dMaceDXb+60ZHaUcCUi/5SS7mz90eA/4w4v/G9n482Qyb8sfZ+BAa0OusVa
uN8i95W0DnDUObFZq5K43eEleXgcFgF5wyw+r/oOW3TOkHucJOPd8Ikz+Dk5
nTmJpbssJ3A+B+JT+qJBwj85/nbi5rQZUouK0thcW9Okt9GSWsH/HcWT79Hb
nzkq6/ehBZmz5BMpmEnI8WEDbzPhFNllcvfXWpIbqtYpyCDcsXNOgiv5ZxKH
mSISeW+eFdFHmCmrq3eoudhN0CzbxAXSkAk2OT9dUooDGn/HUR2Oru8Sssmb
GGRtATURJRP5F0zhSN1nAF1sJqSnxbzLOBw8L2WndTOJ2R/PnRYMuLay5g9Y
KNdAmu7au6490T6ho8hbaLbnYvlXoa05NLmJxl4c/HMP6JhpzPZaTHUH/+Gi
1dKPXiFntsR0asTp3lJZbTN09UQMNme/q+KcU2PTr2quuJRk2BiwAjdi0rIl
cZid0sEU9x/bRheHINI/anw8WCHDPqhKqeZhYLylfCZn02kwncH78bt0ZuXH
bI4ZIddRc8djxzpoaltlI0DbdsaC5Xd5//FUuD6U8GOjk/FCZYMxvQyC5GUG
VRAcMeZOXkFxxj4Gs1hSaSt2s06gPilSehseBeo6Oy/UHcH33PeQPQfmQe0k
kf1w9I2v62Z2CDBKvyBI3WQDNuIRuj3n0+F6XEwmE9heZ9EgFVk8TXoSxlMe
lffIAhiEpl5yMjStycVXVNMFZBeQtroiKPCPfmVEferLGNlHhIqmCByXX+b6
UwMb4wu7yI97pITGtyvuiUekRdtDfEQXL0x5f8L/7VIVJACOp86e3/4FI/su
ZlSOvHCM19XCgV3JUtB6nJlKl+lhhGnZABvGCKo/K0e363dvhCjuCgP7GWy1
OjbrI1mHcfI1z+qFmXUN2EqevcLgwDJFDN88PfGhRe6yXIlPlBBiQo9DNq/N
+xcszxIR1qhWS38+YvmyYNUgEgw4lOs8EyaNfVzrD38bQ/nRf/WcTiPmGJVZ
kajwIJKzb05szQrxe+V5Fy7Ow74H5MJq5hq36njKlztaTbx2CnQL3pMioP0/
cBetH1oRoRsv/HWXCPIV1QeujA2E04ar19byfCra6PYU/lgIsjJS+zpakUfw
/cOtjE+ruinekpQqQg2ZCgNmDpbFdVF17RDpsO0lKYN55hr5cLzYIqeXF2JD
0kwGfJZ4N89H0Nl5Ror3DhNeR6RnvvcIw4vtLJrrmWbK9NQrA+UE9Ki/sU7E
RhhGfAXlFi27icyJOgXwcYZEpPSQJrFKVDe0wiJSEZ4RBaWj6t7xu7e29F46
27PtJhrH+ipe5t87YzMDHAtijxey8KDymQCjwTz/VJjaLm8T90xlZPXthZpR
lz3SywVlLQNiz1YmRlEl6tfxXzSKd0Mh06xRQuVMDCAEwIxd013+BMBSXJad
bEexQnyy0I6yBoTrSmAIiPoAvtNL4qDoZLr0Mf51yiGRmgyIipCqwK70M1MH
SVMBFLuVTJTCNSi5armUFJpwoKyfyjVpYooieuOrRu99yqkgiaJYtVREbYLY
ZSm0cPkM46KeMkKfzikwM4SImJ9ivh+eOyAwtV6G7DfV4zIHLAPVgos3/7nt
vIRRoJcjw7Q26851O6v4dqRdPQY1swx6DpWtfQdcg6s7+Tp5JjDiL/wIojq8
6FK4wust17gQQaFFONgDP2QyZuf+oMv11XY7sW+OHMjrOrJmCDXTe/mI7tQH
r/pmFBvQftKr8TthF2LRB/CiAYTc3EY7XGNqIoH0Dzq+90irKCqJgKxVOmog
+nxZOjFjCRj0udHQHWrjKDzrroZAVYXrv5i53H34ZAq43JKC1KFfbHi1h88s
FMb/cRQqgRvnZApiZiV6HfJt0QyovQVcsOZfFsPUUEV4ULFeH9rXRkPD8Y6t
5N52U62tV5z1aptCMzymHuvT1WWI4W3DLuDJr5Fp5CS/yBtVewSJ1ibxGERE
2tegjelhjtufA3gh1DmmJm7oQHPfrzYEaofIftU3eTtWasNK3wRjJKrpyFFh
YzDeEr6GcWQ62DcKV23LbW79FbmPzGRxOXbZIn0QscmC88PTDlFiXHrmHF6O
odC1IVxj/C/LcA8cpdr+2NssAp2emgjSqd6uGTUYd5KAqOx4E6esZTXyqyXm
H/Kb/E/SGjvFnK/g/aJInsrtDHw0v2fwMeEcCzi3qcwFVoP3BIRN+Be1STSz
p2mqehCDWqhcl2JvvOBfhmiAxU12joLfJn+buF20V+3ZNsYxArDWUIv2aKy/
DOhem8kG/ogTSpEshxizIQTH9WC0S2dkG87s9EVYrqroMZqRMO0T1LX/kPx5
MI0UhimSCDAIQ262vxiKjVze9bIyj03+p74/FV2o07T9lhWT+x9lK/XWXRRY
nB+tGJyeOZyuzkX674B9ECmDN0N+q51TqUn8fZguYgzc5sxvNowkUFruZCgC
7kBjSzf5KlGTOIrrrg+wANveRp3q+K5fEkAqeys3YdYzgVKwx+KMad4f5M1J
M8c6RAGAsXbwLvfYaTE2+rxmNJzy+2nCLbSf53AnMohDQZc/nzaypda/zMK7
Yz3GqZG//v3Vf2ZwM7MgZIpIxh40POgUVuYSHZJ1+pdGAxQBAdHI9qOW0S06
mTscVRL04BFhVXHgLNSKG6wPijRhoQURYKNnUVYAVTHrZSfRk2y7In2p/AV8
2ZsXiRdlq0buLdHT/lFK1BNH7qwzGoTP12/NPMSI69kbBEhNjQexgNzOrzRN
fVejo/wI0dyMQCp9/7+TEIruclq2K0V2ldSJ1hPXvr6GzDxMn585pgqwLQCc
whIY7KL8j8pYztsxqvxtBdAy2kBeqUkhWrQkIGPTocAztcOQ2vRBEQtmXgLp
rg6RHPqgKt4XkgVETEKuglIrqKJ5WESvkl2qK56jyMx19HU4wfDG1aOKYStm
54Izahz/wt7Y97BB/ndhW4t5hznrySVa3s/qv0/l2ZXh4uVMYi97VyvgOkzM
Q7WpgFDsZ+TxfTGlhX7uZAyXQHJwPtdx5M5s2Mv8/+0wejCnBm2zam9E+8Vp
DeWownI7BSkXUOlZtiP76dfT7fa+qSZpdtEmep+uKkmNHBTxoCZmqGA3ZDR3
Fsd7Kl1UAlHaFH9zbPI2NVS8CAv9mo8XlMrs/yNkHv43TYuj9qZtwZDQG3vv
z2j5psHaqCJjp+raVAimgpkgTeFxm3mxJg8KwuMHfhC2KmE0B3rR1dsZL4N9
xTGS2Tybe6zPWeZsbh0wH7xLGI3kd8rx0QvTqtmWHD9gEV9PT8BlMF1dF4EQ
Av/uDggLaWMipiDdqwPhpQfSxPssbKZk46UhYWsqpW2VTLDqFAUxHIYSTSjY
QWX0uUtc+XYMr91+VoIterjzx/8re636+eSc1A4HbPMPfmaRYz1AwoF05WYh
A+11onZBEJBegFP0LtgQA2qieS3yxrCRLsQicHHy6JUGzMmIyAQODSq0J4AZ
zAvGu/8R0Czy+KJ4s1eGHFq1jjnkQskKxWztPb37HmOpX6nFYU2y6hfJN2XB
gQ+Q5S+u50kIrnxXuZ5pFyFfIGu0XC029E9oZxF1XPzCV2O1wiqj4PvY19+O
3qwckIiiQG+ATGcmcuKrQGKqxMF+uSiggKq2TRAzDYgSKDZJDsCdXkBR7Gg1
lM738ARs9fpDCmIiQEcxkP5JVHUrXl4jIbsih/ta/VaTSP6esUAGhVlfbxVu
UnUEDweCv+kscsQguWGxZk8SOzAz0RLDaLYyyyhT/V1Jxna0jMOFtt2lNAEg
VcntBPtc/wuF2OwSSuHVl4s2aRjd3wEIZwaCxNGmh3iYvNEIpK1RPgiVZMoU
k5QnurZVsGJ2J3z037zgX3seOpTVz4gamiizAU9NTPGq6IqjdnLAGN3uqu6T
CrLBWp43ZM7zJ4gWSNZACiCzzgfnm0+XvPtUvwK+oIwLNY7BBgEDKeBqNrR+
kfoq8j9ZC6BCwWgiqgerunqdZgbw4IbrEgZ4RrCq+h4smGuhWcdSxkQoeP1e
Kun3zPb2zvvj5LIniXePIh6v9Rl0R+tt7svCdkmGkSWH3WhlhnMw5OrSnUkT
ppHPwEKhNxgzllB4QPjNTUWksPhRR6EAAzrDfuh/XAx8ks62Si0DoUZbOLHg
EFDjM9Wuxeo5Dai+Bdop/6iE3JxHvqTN4FqCITwzaYtd6P8Ll51KCRGi8UOm
dQ7BZkIyukY630XnXZGfHjPiiJe2/Xe04dS9u4Ihw+d8jdAPZs3GL2TzutXg
NDDrwQouheg3RUR6n4hZodZDjue0pWDp83esraijMnfUZTJwvsXRRzKMg/0I
2HOzdcbJIsd3uyHl+QtfevtD05YZD3J8vJk4Br0y2SCB+lbGR9rn8Lzcs7LM
rZC1RGxCj0l85XB0kJPd3LcDrJ8fvyemWVMev4Sg5iOj58GNaux+9X7UUDsP
y8SHGi7Ak0uXX96HRqKiYjz5B/L8yY/y4VchrDye1ut/2pkxBG64Cbq26nBW
fz+WT+OO4CuKjli3wJE6cnYX8LpD3pUtgMmZOX0RM7g4kfLA+ergPoEjbYVx
AcpLpcb1HKyojMPQ7KEm25z1c+gyTRcIzeacxunWe/7R9BpXudpC4rYK8bbQ
QAlsFSM6cXJyDOGTRrDiQK8KyAkrtynJ57MU5u4cESfvJ88nePj9bmS445fz
lpMUWiy/ZVtBzOOIHX3vJA0zY909mjcOT7GYjdvMDiwOfE7Ln9zeWQ3jgLEw
pO9kIkUWLy1d2VEg3+V4z0bOfMo6YIgsC/hSTeOpxZ/CJawfTtVpiebGlaMf
6lZWQyufNjeqFLwS1GceVf6efEwB3W3JQVZ2XEJPqPkUDz+Irhvgtln55OGb
JimUI2OaZMmJM74q58AgswaotU3imy8Xy8e3VTd8jtW30KGMeZNnH9+hi0nd
jadvO2RhGBVB3aw826yrmGTynYAeVYFw55qbOKilk+ynp7WRPjhe+2/8EHHi
hHeO61gwmobXddZSS27hHWbt8+NeMbn2G0WlSBsEqCSXI6Ugwrpbq0Xlijq9
8TNkFqu7dD7JIOFHPuprWIa9qTGu45Sn2z3n98xTmDU2bow63IAleiLHy5kn
ahRENY4PY2w3PUUw1AjS86hq3DsdZRNjJoTbo458w2UBIXizkpHZrVCGBug0
4lsyRMExPdNMFEqGKm2BaQrSXphc4+BKJDGW0UJd5rxsTtdrB59jWkIatbaf
wdrPs73p5GeshM+q/BDBnM7DXM5bcYG/oIGl5Bza/OyLbmxyZcrc6OIwHBQd
o84z7qmU/GCcrYAuOTF8LA6TnNH/6fLUB3sef+HK5qdRfx6P2pHNpWFwlza5
Bt+oVlrkOQquzVCk6PD8hA7P2JMuRdGQ5lPxE1y06CLgS4ccnsTq/W2lqIY0
rlvhzl2GdyC6oNITefFGOKgE7rsTGg4bfayqH94XX0AV46b2CKlQwNa9+RK6
GHo71LNwWS8+6GBbQPqQVrkXJfxRfIX/8J7yheoFkQS0tHL70coXHEjP2vm1
FBCEEQheZv/sHZA9vr9tPjWNFTyYAzznBE1tTJBbTTTWdXut7zdsOhTdcM23
WkUjyzct2q6DHYY25KO/KW1CyjooIahTafxVMCkPlL6Uy8h/leYLuAv75HZo
NuEHuXGPTEcef5caHtXKJsOgI7mgomVxYxj/QvzEko1D3Vgqrip4k8VEStmC
mOHlNs0tBfiWpfxAmP+6xzY+8hbhABmd/C2Wf40DC0cWfTrYdIc4iaheqr8d
WAGZs0k0NRuMyrJ5uztQGw9ijZUl/CrspPLG3T7j4BiE0ZmWnpRH26sk+0Cw
XNXoNllBHYhmGMUNyl0jH9EZADpny0tqK8HIxPvPWcdI6VJjYSvaVeVDVzge
OgTK7MA0PcBNocycYUVVouObmWJSl0bxs160QgrS9CkKG3hNnuOxWAkD+EYJ
mRI5skbrsvDecvJmvQ/d0ykCtwbEwvR8Zw/8uPtaVCjnnW2EWiij4JnqaIKa
2AxN+E4xe+ihqEVIyBZ1OIE20ZAtn8Biy/SXsf3abKSkjdkMXJDO7PYthllz
pPOS5RC5FOTC2ODVTltVhAc6X+NhTkZ4mTxH99fBFn3a2YpbCtta31hzmyJj
h1cDWOwKgPJKsJJbs1kAl++iVNzzbNQEm1qZDh8Cb1acEfdMtJ1+Vh17lOvJ
RHV5/l2GFQblYWORpIRAwXKilqnlUjwCAWOfuTD+I6+GIaTZiA+ex200QOQe
4U7C82iVYRiiQ5fhKOhEQhq3VBXMyV96hqcK5MCI47eRCyamxmOZ4SAoAtpb
00r9zu6huJLPi2HY+8vmCCYwmG4vT7EF1l8mWTY63qTU0hZLjGp08diEdb8b
aXpyq/PHlqwP9jpMokd5HN+pMrZ3BAcP2m1IbUblXwv9LSY9VFEVG6YBJ6e6
YuJEz/86nva/DEo+cvLFVSQlyK4SCZL9XBHV6FLzl5XVFtd9a5DYqGQBGkUg
pPnYJbmDaFzZwd0yY6xrKMFhDITF9TZikbpRTnh+b9KQysHU/HRWrA13EzWj
ta5PFGtNtvIcrfGEKg1DWWan6rcFw0yxl7BiPC6HaOnppKsDIYVJi2C6axCv
aSyKdOBPZY1ivpDfWyCSJAVDMcoeCIHv0FqUcOXWnn71oa18mChnmNuzxlR5
Nt9LHCrCig+VutzmN8S9xXx/X2i1e/2OKaiADr/mFXtbCdPkPRp7jMw9rdks
SDlezBNLgfhR5dxQLM4/3Nzv5Wnb6n7KHwUw3WixEhOXjcwI+MDNQBwWr/G3
p3P+vzVoyWhl7j+Q85w9uDXwDGPBCz38yGZEwH9vLC/CruCtDyEH4ByuzZki
oYhbLfNIBmgBBw3oFmueA2oa0PuQMRzLJcAS+zcaThsY4zxXjz9cjQJuZ5zO
JivPtQUwQx/kbeqKklWrAfS1duFiwMPo7hlGAYTbnY6FIAbOcUkiMxqWqHJJ
D326gqx0E6JvJYeaK0Uy+mvqPxr7cNEx5UpkNvpjc2xBnGOd0291bIgC4EHN
j5xy+qTATFFHq2IZL3AHQd05o19U0MCt427gl8iAIIslfL4mEntxPHSDV/U5
0d+26E2ZUSOrRHhKFEOFhxPJghqSX9ZED2wKlVN444hUGwtzXxZ/GFTRf9/y
uivKLCnfxZ9QpvZSDq13jicJNosaEizm1GmzLTh2MfzCfC/MedhyvKk1VyA0
Nv6f4A4pYQ8MMGXof9lMpCBoF0YbIshfPG5W6j8/J9HvK/wssXpwrBWk2jhW
vqxtb9PcewzfcKLGgyOtbVa2D2pJJaI3kM99VD3KsXnD44BuKdNmnkrWFk11
BkaF0tv1/waEsvn7654JUbLd8GLKaUGLlkkcmLtT/0rGNvWmV7zLTMN3BuPa
48x/mPZ1wi+rLDp1oAWCdTsKZdvxaJwd9tNNPSZ8LyD5s8qGDhPYZzytl1b/
O1s/OXlqACrfmP55vwDTqT4UkN4ybEOHsO9AZbh9zWQY41NBAbryPZC51SgF
B5ZkC8mwg3wAXwhaAVmaEVLrm/2D+YVZdqFzB5jEvqcsDpTIGlkv0twxVXFx
PgH9W0bVvEPs5jMMvae8oJGFh/p2GQY9mpGiuqKDRyjuk6FzsgFh4fHwUR0B
d5/p7Q+DlLRGMw9K9A4poj0dXEDS+r9NYANXllydZJ3P2ckSFDPSv8z2yEaF
ZyHvt+MutXjZIAjyFm6LGVJKNYO171vAcWUUg7APp4CV77iBKBPZt2F395va
F1f+x2BpJ4KL32WMpF6ulWs26P3KVnWyssJ7l3Wjdi8JX1ZRr7S6OLJUt81c
FPZL22joLiCcUc/L6Bkm7c9qV0kd3jEY0UNdGHHGRwKtSmM0r2Snlk1uFNXo
489F9x783aDJeqOFnqs6V/eROSLJ4IXrtT54xxG5s0uEzvBOYlMd3xqoYZU+
wDtSWPqaOTQiryjNn2c+YCUIsLGdj6d2vW7qvnDeUvxzhwraR7ZSpj34RoVl
gH7IFdgZF67cD6vQoc8X7ft28zadP1UULxO/vG4uiQ7dg7Yclus0ozzHtPLv
a9zFxUOMYMnrjDUwJBVGEbFRg1i3O5Zo940udWdv+fCjUmu7dRSok2lUkfTL
rqgn7zOtZKPHaS3mqCpPDPuyHgHfEs33C5/sLISZYR/XxjccBs5aciVA9EtQ
tMQNtl4aJ36aEPAlo7N/FT7l8VEk9nEB87IFZUrXSIgrJaPmZR4hyIr71d9m
lcsPXs2KEnJedS9py8shl/iOMF0u8ospmprSWt5IRzyeRrPw47P4+kayQ+6W
3LpvVLVDWakghpirZzA8yt8L7OEoEdc/mWIucysMDGXiz33r61GlJHd8HYNh
/5vizueJMOM0BZQy92+MIoLC2UttWLmZwSn+//PjQDsND7U/T+Iw8qPuOgCS
cji51xdl+3FZmGshcjhCoLmpIyzNzNp29INtattLYf92X88fok9SmcB0X305
Dv2zRVavzUk81YeptGfM4SG+eMjQaDrpEGnBkhqMlyfq2lOoG5WMBf0wf1rv
lY8lqaTPNiwWo2sW3SaAJeufZMOVa/hxOF0g8VOV0ufb0FtVu+55fVUzhDHd
1oHIXT31qfjhW8yGroR9XPb5FO+g8QluQmcAiFoUXXEUtYcRXhEw199wnfGu
h9vIY/02JecMuUbFbrvprn8sMwWj8z30COF3/icL43AzkX37aBOpkr8Zm/K6
2zifK2tBAC+nUeKuc8jLKHclU7GOYdJ0NMYgPTxK19/AqKNORBmH3KGHgal/
pnie8VUO6sT12CZefhynGcAJYATGwt6GKy60HKRKccaGs1e1+e1sMUJLuKKI
Jdnk6vMj69jdc+fxLM7FIRKsy+FqAP1JnFF+ZgTaJkkQdKEP96F84CZACIS9
BKiewoHJ8zj8o88xZ6no5+QGxnuznZrL8JInPvQ03Q/v7EyGBf/Hdxxf4luW
jFSbWqYr+Icc1foWGW8qrHkmnDJKLleXUe6roj29Oc/4qperDyOxYXFpUtbq
7jrJ60pUp4KSTmoCZ1ypowAvaNOVeseju9epnGEHqhl/PJ3SoHKWRStOsFr1
gZJZapnONbhp5IAFIwUPZxoH5kRJgeby++gwp9uoBeOWCOgft8lLPykwCVp3
1VqVqv5rxg9O4Gy/1FInfBzlAynWWq6pnAcYEvoFKhF6056snX5utzuLLU5d
40Z95sWrnHj1roMMZAI4ftywR2lI+xSBceWHqIowjvIxDJWwTXYtz7gtjBVR
gPGU5U4U7BJQq6gsjWIntdDDEbneGR9zQGXyLHm9n67H+u1O2Liwh3R67/6o
vJIKq5iRmYtRmTJDIH7ZwG1Tf5m62BRQ3kc1uXMll/zfk6bB1OupUhOJzNpx
2ehPA/2G3kXUCl4kQuceB2eiSywHvzMk77kH22oM4C0gwfH+WYFI1HKJUset
TmdgCEFiLNZcVUwHemLwuwYOSAliBLR7nRf2jjhEX/ZMlFRm0cFSNxh/JLox
3Zp+5SaPhmrxFeiJoJcHn5BaDqt1XRJnV6DdP3KoU/yP8JFCa3YkBek2zWv/
22i3RgI4anyc3lqNTVym8IRR1gJ+Yg9avFht+k8BjJv3wPbvvc34GiLOBO9e
KQa+tgP6JzEfIeZC7HBXNO6DqpN9Jc1rKZTvO6yl3gYJzrd9ncO88tk+qpaT
tTFHkqFjKP7lzjXlTf/pjRetyTUOne2WGH5joIvuYfstjYgHm/KRXBBpCXz5
YjHQaKunB4yq44CT3GCID/aLXskj4fWh/2G/YmTDQ9jUR8426x6x+j4uE3lw
nRj7Z6TV/BXg8C7Celf/2UFoCLbPYmL+SZfHsEYpiDlOt53jZ9tn1t4Y6JPb
kJ6m6JvWkgE3MvI7sDzyYJgm5j1NJwZHvmVUNg5MFRYLw3F6rp07AcTtDrer
AHAachOfMfKVZ8rAnmUPlCfz6USNB0QhXksE5CI4Iw1CwI/0j7doQbO2a8DS
HpxPiEMLE/X8iypSew84IQchOgXkvf2HXv/wQpG7uozzUjD9i82fTFsOByi1
A77o3Z8ZZ/PEOpT4QgtFfVthp6rwkdI2rQSNZtkmmr45hjjj0/97+JoTqxXu
ZMb4zTrHQnKhGCC6zswAgL46xXETIh1kUlZZ41OgvFi97XaBeJtIKdGr6UQZ
Ryw7/h5ENy4XMkPvI0BIrkvkoLscVqJ9Bj9mloQz/jTC4qzzxS6l3i6mdC/A
EqdYUg9hIeR8BzaBjZ4TEOsmLmVzbcd6jof6lrgyP6uQzK4W3572bcTh1gkd
AbokjQ9r94DNnK+OAslNnJ3EI9r7HBartnBqvdnZxUPPmu//i9wb9lZvHYXB
CaAeAV5VR13dUOa2thK5yefpLon0wAtVwMDoHCa+ctY/TWkaoatqxZQ6mIcU
/TWB/TipMQVTv6pp5tjqR35Ib898wa8kjQSF9/cQuxdcbzIDei1uSRTXSjW8
+3cZVB6b+7j6T0XaeveQL32ildkQua0sDf24Ha/pkP59ZY97NZdSTOfQ8nd/
mjY12FRRqa3KEA/loggTX39ozuNdFCZ1DcpkFB8nscIR7yGr/TtwyjcOUe1X
EB/zaZ9axF/b3F3x2TSgOlickArkvxrgsQXXkVX7Zw3HiYxSEB/72zPqeSS2
7IKkVQrF35NYpJtQeDb1XTk8R3TdomFfSUMn/dWsWtOc9kEFi0YNWNGkJ5tF
ehhH9ZXfhWJ51P8TgqcdNCR8F3eUCoayfcARJeCJiMNIa/PdKmrOCN12tLEA
PT+wNwwFHi7sMzi/67fvLK75LBK3FZq4z3rkuEZk8byqp1HWU50tFPyS21dO
6ulaDKn8pyOZXTz4epGyiXVNYJQ7tapoPPr+ZSUrAqjYJV67EkUBnYuP0W9g
vdxcVOaxiv9BfWiQy6CyJP8i4zVrs1wDnwk2GXntehlpJ1hTsZ9dUGmf5M+1
9AZmtyJlbq6HI1tYsDMzkhwGuNp9wxdZxWfSCD42fbCrtiBKqVFGLUaoS5pc
s+nh/QPad+oJWbvJ7dKkzlIDAEwJFEtAITzmfNgmpWWpVyAqeCbIt+Bl5X9T
aWRgw2X7kWHgP19kKgLC/uSESyub4Ks7M5ZsccB3QwfPSAUkwDFSyVbnQ7aw
e9y9xpLXq4Ufj4yuUe89P4ODKM0fGiBtZHIgGeW4kQlCXhKwJFuH1rE0gVM1
EyTrgxQJmLqqfyICcule1gu7/KiXCXE3uFq9Dth35KfE3+rTlhOKasAiEhOp
aMwCneac6XD3AtAGLoytoCDiEg+TWEPbgdmWRxHNirt/CYsiCkHqu0ZEpOD5
BMJYgcp9xM5qjuV1i/85gAweG72F3C4PsY5wRQ2SABgA4KvsZOv0TWJ1uNm9
vHFxL3sSFXcSky7D4yq12bNpXKR2ouSARCkV0nOI4SNxPxQXCEete4KOVoQQ
+nVCW1AhIC2eSVNyJdt3loseEDhjhjgriWBvT4Gq2n7Bv+Jm0xVRGZl2rBPY
tm5DWzuXNDB+lqQ76H/GoElhdeVUlz520Q5/m4Ochk2t02tsQqQ6ZDGCuCqI
BHmyDHWJ9BYV3uUc8r6P7ZXMaEYpDdl8nFwEsqJ9AYXDd7zapqaQ5JYJAiB0
2JLCPS7kPBQf1R3K+M+xDNMVMs9j4ibiaFiVn2hL0yYknsQUecDHB9Alc9/W
fGhZmw7gU+iG9VQ7Xz8qDvf7iaOL3FsrcyxZ+iQPT9BGb2dMIByULXLAG+Bs
X34kNBmO7YLu01lfj9xcuhlZFwNEKtie1DYPUV1dq63hd/GEAQKJb/SLHoxI
sjpR/7QUJ8HsAKACjq470gcwWEY0R0oWVKwFvszue7h0dxcywQ91Dh8oKpk8
Eeyvqyh/x+XSzp2BfG9SitNLc3962AKho6Lykgnsf+Osb94sq+V2HqmBBjAR
GtfxL3U6eWaRF6Ub0Ovw5IzvElcLGhSoUt+jWWQ+Jo7pGX2/NZ8O8RPcyeB6
LoXD1QFvR9NyFH9NJGT299yKAX/c+84C05JF4UH99XmPqY0po+P7r79OhnfJ
EIjzvGsiplsz7baYvi+WamW7IO8XPtAd0BO3IkvDkWbJouAIoOMwMKDQgDkU
RNr2rPqhOzGBZuGGuSONkDUQCDcOOjQMLC4IOxg2RuYWFGoAmJ9QRfF0Qaa3
8Vjw2VgsBDkAjx5NiKzBwFCkGddzhHNlZVfh1n29aQam0oIz29HLL4pWrfaB
6bagbZpuQlIo6+OPYC86ZXVfABQl/JW7LdSXXnf5JLp08fEQPRO8cr6vVzAh
Fa4wIkZTJ9nmPK/yAq2kwKUoVNCcEnLCubF0aT3KKm5xt1ZGZbE7Kql4RXvo
xEwRehhCcPFQCR2CbzRYLYthzaA5/JAutULn8ruHbycuJg6K+hdfPRqse6U8
PUK/mG0VPzAPqu2rnBo448JCVh+940LcHk+2NwVEXVeCmSJNPDW031EQ7uFj
aSx0o7p9di6P0JLLks6cAqIHPXWWPn9nPrsML8kqwf6AdRhg7abaL3qmoBAq
fxsnDsaEK0Zw1xSV0mwnh/ht0myRwW0XeXGM2ll9xJhXzD1+KQiMi/xQ3ZH+
2V8E43E+3ipxzWhhb+fypCEsDt9Zn00ooDUZB1dzi7PRNRK4J3LADxMym1rz
TR+c3hY4W4OLCCoM0uSi2cbFtnJRbTfmJo4ew/7zTUMdJcs25Pv34KgkwVwZ
2tMdExrgVc49KvqU03iSbLRQWpLFvxXJX6/3gzWJiyoCVl41Q/WbImUFWxRc
DusTDPpoGVDnAM+HAnVoVXLog1bbHhULF7iSNbKq57lSWJggViWAidBCpSJh
CE42CaHvhKBRWHhRKlcQB6a5AyHJyW/2YcpGEJZHwKd3GnT6qxDkFl81jUEK
HN59ee/4yaU/9Y2xRj7UQvLd4cMJLRm7Sqy9bvUWgXPfT8aoUZFyrHp1rXD4
0fx9N0og0yicVPPTV1UxN/UTONFl8XdvwwI59NtJVk3865s31UzQwdbs8RH+
qmETFJF8M/l8QofyFxBLFsheaH8SWDBL70WEStBiITZpb0ahfEWFcHsFKbP7
D7SuiLY6Mcz1k9tJBJPq9pn2LV6GQXTSXcE07lo2TVL2Y3r4h10frSgbLqF1
k0NoHKbEeEdtJ0u8KoSk02V7DgJZIWcT42pUs7kMqWvZpiRVDFT3RJ6DnNS7
PCHT6wuXJ8EmI4CDeztRVCCrR6ocJ83lI2AIgRb0jZL6WugvJd/hWkQe6QNT
3HXrEqXWGHLJao5yHGkXwgPn4/S6xyWs+rn95XwzSE6GD8w+kpOz4vCYCNER
q+dRelcScGw7vAl+u4dWKThz0s92ZTc3yS9FQO6jttySH7l1Z8u6J8D9Bvkm
xJtqgpkeg6xTYL3J85KI0RrfAmhn95F1nNFjHIob8aQoZgYVS7vOIseEAxGz
+xy5a79IGRaMJD2Guvh8cP2sgPFqT3sWIFsXBGkFzZndIezNuxd/dCP8Yfp8
qsDbkuCioK4FRPAGTxHNyHQNbkRHL785vqGxc4Hm6ZN8QpYqw43XudSZ2RQ3
Ro4QaRuhWQ78bBsxFcAV8CqG+4BggwVZCDJwpLrtuJ66XyD7duEGxCB9tmYY
SGOW54hl4owTIMy8Uu3/BxjLE66hzlYcwrptmSh87Arc1C971sF5XaWtulca
LTt70f8PvL20Al6vzyPaiwXnOnOo1ToQHzAM0ZtkOlNOdWW8dgRuYbTKamsH
/bQNvy2WsSTkpas8cWgJTvO3qJPK6QxSQmT3ERdryDOv+BYttixEMSFSoYxO
3G5i9teChdxlbvn8J0A9aTQoX5E7HM3CN0SB3ZhtJ8y2R+zbkpTRx8mQNzoJ
60MNqwwg2L8sj6ZAYJvltm9kim8/5DgA3jFT7L4IONzVKzVctEuCDgs7WQpF
oV2SoPzkdoQCESqK3kjK6OCa16lNbcXU40coNLHN2sEHGi9rOWoAm+JKlpc7
yj0fbj5/04uGYIuizRiHEHorWVoQA7+ahErRIl0NstnaeM+QbGPoHCa9cPex
xDd/Os3/ToABKJL/smdepCh0SJzeK3R4dogdLI4o99DVF+TuvY4Yi4drvMEu
sOAnnExAnN4DZdELGdBgR1cfhUt01JGgNkx+gKOOyUtuzca43CXaSTnaC1m9
bbCD15fo3Iw64F+AtkHAVSpB5WLgR7jxrZGclfO50uhtTZ2NPdaa1liGv4Rh
s2mgucJhKh2++NFBxGThv/upoWVArVZgSboKtMXAph6skmjCbQ7InXGQyE/F
5DYKVY/RAY4ulq5ZgBX4oUo/zTxaNc00yYSaqQNQz+W+u3a/KgFUlaEDLJCS
yf+kP8VJHf+xR3fHQ/KrnQeuN4JLYvpOeVtIzBIgKzEq/kIPhMF2RJHFE3q/
4vLArJz1+s4RUMaOcAi04R411w3blAGgHNJ/QL8Y1/Yc3TZ/FLe45Inb2hZT
AL59W7dURXmqp9EMgiwOKWgOHQXe5jj7DZhmtfZrV3xHu6bV/+Gyz5G8jgPm
s5btGUk3g2Y1MX5gdDn5tGEOnMUXL+f83tMyTFQ2+XZeyBlwuWgm2fmVqt8h
ST6udVEy4XE4NKA/wxHcWKL7VWIp6AwtDppjLQ6hZRKvX63rijcZ4zPoVlmq
HjwW08kP3xs8HvrbF+72YJw9eBFBQqgvACMNDXCbVQ4kjDZb2VZMXPiKcg6z
JT7BzX+kf0PBTCrDwqk6PxGdRWBhPqXbCiJWllKuj/ItgHLmGROUDmjn7phy
+APFqWtmhwljol6WS2W494irpR9FQSl1M/lje6I3JiDOrl+7MqbKFNKgIRFg
bS8AQS7NtiL77r8tiOuCHezmFeVBn9spsHWossPnEFbTCAqQVhgS70k4Whh0
C2e/8HsaQz/s7Vhepg2OzYc4yBUTxnp2AMpf9iY0Bbe3Ot0X5R9ZcnIcNTgt
RGbxDQWLTiPWlIJLZwK1Qyq+33Rb7ntK2MSBtYE+murgyUtbgG/s9KtOXq5O
6aEewNU8cupWmUy1e1K3r1qOIXCRlVXTdKVfDuh8OLMeo3ccZeQf+J+iHP8S
+Yw1ikoSg6C1W16WJP+JYzccxZXrGzrBOpEL4dD/7KtQ5fZ8GkagokNclb3f
QyNFQL6IV89jvfXFR+qDph1nOuJYG1zYW9iBoZFSoL4cXMXoGFe72NjUolre
e9BUZ65AWLXyjB91N1HmiCh2n24krd/ee8SdhYXYvKgkXUCe5xunPC/HT3D/
uf67QEEQ2vpDdMZDL9RjwHl/3NcqzNEFtHpSbuQJt1gaGNq3nz7Go3nGy7Ay
nfkV9YkYS+Yt7Xbu+tL3OZDNlsLr6vJqJPk5fcna8OJhwhDJkNtMoCCuHPuB
BSZ4xOnevCQmBCtd+lAHNg4osB9ReNCls+7wYYtaV2pOxUFF30H3yNwMhMRg
si7gzK4K74QC1HddwsGuzs/otNvvu67SqT2xECW0kzoisP+LDnyxjjcpMocW
LOWmudDrSxAvPVAe+UYMKHKo6CQL8ZSbIj/2DUF4jiOXhH8FZ1wXX+aWuNFk
6x2jUc7z8xd54Q9d65JBpLMalzmdUeYIcd1eCTogvpzcFeAgdYRENU2kO1TG
8mkXc63YswUxycQtYybjIFvD4O7Bq4BtEBPSy4uVFm8h7W+w2Lnb1zJ4SmiT
sOnJb1QuA+j7mFtJVajOI1Aebl1QyVxD5MwoN+L4SSHoKbRslUx9y/kdNVc8
Up9t8PAMZeKXDY7rfSeaAbNq7N2KLGIP+kU5FN88Wy+8nNMntR7LKyCvFQdK
bkjsKR6oXugymNbE0385eU4TFkryI+8u/K/W5gWrlgHK8NqDuwaNcc8WnDjY
2WyEbCirLNEKQb8TddbL0KySO3kdo6cHF7BWnY2eE1yBp/6yYy/0pKbZUtCf
sijUaWUG84gEBzRaGDogVm2ss9Tf0ReyDAK4NG6vwUvML0of4eFm7TvgaHB7
4aV+2tLeJdt5bGLgdvOJqZiiQYY7cTcJ+/ziuW+O6egxcx2GnaooXMFV66W9
X0TP/OoyWnqhWhr2sqIZwkNIk0fO6685HGTHp8qZXzTxnT9gNvcZObu3SgJH
gmHoo4TbARVM5CXUU6jl7dmqdQ3LypRHzIU2UAe+iDwkPgmhwEfxyeDL5pQ4
a/EVaVBJiVkVdWTQnE78rNH2+q649X5xHPqXFj/3Bs4TcI2PrfDo3eTYmqIp
wpSxHqn6z8Hk5QMZHFUpAYovFkoiwOrRqrLjfd7QFa1cA022zbT0dRbxIrWx
8CJ2SlmeJ7d2YRWiqS+5J43JF6ceTpruRrieFvci5rdMVdzCNq1BN+3R9ISw
vTpoHial5oSmGFSVjZvAf2QNVuPOyj+LEUR1YepEeJwxd92cWFNzgM3Ti9mF
FY18X7Cg0VH1dKdkn2Hyrhpj0OYojwaNvfatfRKVyAy06YA5hD0QMTReUtZk
tZw31RdapFAKrein9M992IzjTL1V+ITOsHEbVRBO2TT33UBvu3AI8yLICPgP
fZeT0uG2QI7bhMBv+RJGg28P/RWeq3zatQq3NfJrCE3VamDzeP0NR8Ucq61U
snCJYm80pH03uTX2XxoWfexyn7WUBjpTFT3lEi8plKabjHxC1zqCD7J5bV79
J07D2F+TxwHGW8c8mmq3TGEQcD4XXvqGhSdijoivTulGZ3c7Cc5rIL5N8845
WVM2aTPvJS617WnX4jlzw4miRfL2vEcV0k41gREiUhXhAdV/y7xm/G07O9Fy
PQoG35PEZwM1mgqkEig3sIGmSWstyxdrjl00QZmTjWi0MEVKsLnQxoudw0Tg
2r+nMEC+zBjWkGc+F3zkaEJUn4ESwVCaaEfMR8XDP7jwuAPOYbF5wbbRs+2R
us6ifygc+EdWOIP90iGgoSfYyUUP+XLX+ea6ttN/E7eZxV56DOofzlhsG6YJ
NVwmS4en3hke+jbURtwqsic1SbVGZkjY+awV+Je8ruOOcRlsKSBQpaNLQeAU
0sqIKGL5d70736cHZzmDuaY++MkeinmJVnBlclZN1dCsJLG18LU5mj62OA4w
TZzUl+TBEiKiA2dK/QI1nYCnoUv28OSjn39i8VFZc+ypKZlQaQSOW1PcFxFw
/MfQazDJomifpiZICSJfVZwc+t0n2NI7ijr0W7W4V9bfOZ5bTgHkGxzkOQ/H
wq2AIODqKGyaYYG0vqi4YudXgFxtBX5/pZz+IqMPyer1eihW+vwdbJp9XGyn
qJjvMAoGpx4on2U2bRg243SotoncMVkRWGhYQZwdxwhWjzwj8Ygzn0kpVgWJ
fFqMc4/VD0cCkpU+FAu/SiZUkKUDloRPHBBfBYG7UE75W2eHC786H+8hUsN2
yt8169dzLMIxQbXRj3XL8FGQt0plbwH2WcKphXmX18fyjObB1nsC1GwRbvOx
3Yv18PHsmJ943VpoVat+4WOirSevZ2iTLILSw8tO4DnUw122eS92XAKItjiG
HmiP2rc/dV3GmqtgdUJO3O+Z5/vSrQQNzPUSxayCwHegfPRnPc92I2JsSlGs
wViXPWDqDwwYeMuClzuMid6O7EIjRwjPt6tfS/4r4enq4yzRORhJX0FXdeqG
3fXyhWoU/xYF/qT3+h637jNtHYFasJHlxqjruAun3OrFfcG1s0Mt9RjowXNA
RmDPwVjZcxtEkIdEY2f0BpWmxRK7J0IGvSb1Elku0YAck1zvgZTaa9Qmsu8N
HrDSs2hCzN89GE39OQ90WfsvoslP0Enhv2j9NKeKaFof0pmKy7+8jHi9ZP9h
rzY7tOyZmB5hnRQBDWUBUrFahwxa8yx334KZZFicWr/Y3x2X0wuuSR2SqPLQ
Dwkoj+AjnkIHOzsit1ZnDEeeAPjSPQUWkQZ4bEBZSLMQfwzAocZedPG9b2Hy
Xejw0yTdl96wdXGhqejYBI7Ce41sffjfqfTbYVVekyF6Tv1NupOG+8zcHPO9
TsksJcPFQsvlmzk9Kv5s5zk8QGz1je+4A5hJPPKyrRN2/HoOkVgCtefOIPNw
HxxJVCZFofUUDsVlCLCmHH8k+8cKeu/0lB8BfXHlM95irzQS8DU0KddEzmiZ
aT+0ReTohSqGbPnVZrcOMAuM4uJHUZab+qXHizH9Oyn0K9C021WlNB4aWFn5
xrArASl+yqqspTAmsGvooKkZRB+pXOwrMaoKZQi4XWJCtMQ0QI3EGRAqf9iS
hhMTjZmId43BCWX+CmPMBqKTsJ1CiCUsHPwvQi+ukLHc3Xjw/NZ/g9cWJsEi
fuWETtvd27iN9+qhhJVqFy7jubfGafQBJqPBFWzh0irTdqnAe/vsc57i549P
yQQl9FdqSk5pqL5OvCXfxdDdr5S0zndnBAMO2Kh+c8PMw47iqZqIVFvL+4xg
yYIX/prcSinlBq5+cBl9TYK+n5Xtn6rtwRAtW3j9d1uoCm+Cr17PmFd1Wb7n
aOkX5GLT4kUEbQWw9QotNuC8Nj6ELgvZ5fBmk3fY7AGZr9rDCJhf/yL6XoSx
H9MnVgQTj8gkjG19rdWhxSm0qJd+QfmMcUaEAGgn8H9hp8/WwvwglkfLBgN/
uNQdn7nskAA3jrjmVKAirhGvS3oSRX/hjBxf7iSn5dk40F7cQJVUDAesjrJR
BFqd20eP4wL1wHnWDJJDg41N8EotLgwHkeOaGiJNUjaR/A0LWtC1SEMhiJ5o
xgKZDQKhXW+2hlh8kTEdBlbDOv9/kH4EWJJu47kDPQXlcHu9tN+8g2pPLPvZ
IaRjsRfbY14QivtBpR6FrCMSfSNK8Hw+PHMfd/JXevrMXXbxkYsGI6gjX5/6
K0jDjp/tcFQ24SdprYFdOKnwMuG+BeLYMXv6ZuQVcnw/oDpHq8/MdVu4dNcQ
fgSqa12W9ZsjIcApr9Ekfsg9DqcnnHrWZmsv/b31lTO/bzBI11vgD5Ikrte4
7vvUFZ4ZD9Mff9vrWhwiAVOtoIGXm3g6p4Jq7uPtFEuRYWXIEOXr68Tr7Aa5
kIfuo2knJBhE6T2rWZn85R30GsD3I1y4bcYn/AQNcDWpQIShfebCIdy7i/Xg
8tIek6T9QvX1HzPCs5sHw5SSIY5m9QksCjYs9DsCagzWxBH9Gt6tSt1+EPsU
u81DLUb61nePn3HYPi4kybW1Ddzp2G7CG/uqq883WZS0ekfAatjzQFOlm/3X
MrzJJ9cHWroKhn+IXq9CuCzTvCAc3OHUxG1K9rbhheVmb3cxfaYIesm4hLsh
uAbNBmOoHycMvU9h0Gt69JnjoQbccWsa81PLKsptvP7Mj5Aioxe7uiQ6EDaQ
1T4on95ogmrGBSt3iByk2VVy61RcB3PqgSIQ7w2+kuIFVPZ/7bFqqZNK7Ac+
vNDKosOC2JU3/Hb28qFEofCb3YktlXbEd8O0Gs/9b0cMVbWOuv4K8XfzZpsJ
mOTp35/85dLq/t0uXd8nzQ1MbhTItPi1VXovEJKlzDzLGQ8EWSNCMy0zkSAm
A2PIIBwVQVOZtAXp0qVhggF1LLhobQfzhfSFb76earxKA/gd2sOqlXvTy2w3
/q0iYfruo6KPFQB3H+ai0MGHqX7ALGMQu92MgdFCcH1x91yVfSGgbCSo2cC+
ciyLoclpg4ljFqr3bW4lywpXdZ6JfWhuATw1LS663HNPc++Evoe7Oq66GYKV
ucJZWmJj6FvP+GzXxyDHYiVl9xoaLegFrghga66F/zczp8sFW0gRfrpMYO9O
0Emy4TGDbeZYaWL2wQewbX/L891SZZGQPmgdAC5LwiyYkZZB2CdbAf1jdZxg
Udob/EdrYL3C1t0QYWqridjtnFdDVoTGIap/Xu1ooIjw5DDfgJGICB8XyMcV
i3K9Jj5OsCmkrbgKnw/mUi78vSx04faW+vD1/sHuCugf+SMYZT/WFGc7VfUi
LvXjPA6oK2PoG65bsKpgUqE4XFCfxDgzvxk1ffXDRCv8/GCPAJtV11vKLGta
NNDH7WQ+OkZDpgzp3ZCZqnAxlleYt/9VM52UjKWC7k1QAUAD7j0lmbOClhv3
qyy73Ez9ObTe8SYscWi8/BV7kM9e9zW3losmhFHsypfOptd1/3DxviDXNIfa
bDBvtAs8jiMXjkQ/gJ+QID+prVhZWg3TiR05pMQ9MhLSjVbUfebEbiy6BusT
RckRXSjPV/xQ7aPSBZWex4OJ2XyKnx4R2XfguDqxemP0is1NcZBkxg43cDX8
NW9Kdeh1Y2XVvfPWrPYNe+XtZyUgnMrqbD3oyaIBdKBUDZxMhMT16VXkvO8a
mQB0d5QP4GJ0xS6l7cz/x1pNzF6L8FWiLKk3U7vr1HTJakrRAGCbaL28XRA9
WGvvdKYymVXsREEI4BxmnqTsziwUAa7pSMONxd5ch9+28DixcBcX6ZNDjkDX
Xhl28TVLoyu98Ldi01mLLGVGTdRZx29XGr+qReKJ4/agYvQnhrQlsmeIvTpV
khWEG3o5liuPn+IZKQScg0Hua57spX5cLb0yq3fdApfN4RWwt3ImM/hbhtbm
ufoAo+gbh+w52Yg2uU47icE0GHxOuJ3HHbUWi0o/xvixbQWPXEKyJSomEFER
wOXf+ttRUaZUlYMOF+JFntUAV4VJJgjLoluLaOoZhyBTwYo6NyH2qWakWvZA
y098GBDpQOkMEvmXBq5El2EE9F8EvmULdgI10qUtQ9He+z2D2uWyqIumMNWz
Ydwre3a239OjlwC5K3rB+pHEskC0Kf8w9hCJoD0X4RxQAu+AI25cY892dluq
jDPmWe+coTsmyqBnDC6h1ofDbO+wLVgJdYxAx0G1La+0lwAAFB+1rmbcUyAL
Kh8C4gOsuDO9AcqF1MnzrvNXo1lgoYp2XvO3l6H06+JfmOnCVqdjhb893tB7
gxZ0+ODYRlG/3O9ohZ540z5iB3feapqrgO/19l/DFTzIGNkm1waG9x+Vbbzx
GgQk2Dm4fTwlFtdv5MkTNvvWkBP2YHDYaREofsrbH2rxE/DnmV3DXMJHXN6M
Ysq1UQCK4CPeyhN2c6nypZgT7SKoxltmQJkYLjWql5NcuI8zVfQYfqVjT7Ul
LtOcWzITSXpDOkdn7eb8bBrhgRa03I//Bs5abYwB3eL5rGFKW8b409JAT7i3
UTQA3Vo/8+4LTwFTANMLzGA0bd49An4G8fLLydarYJA6F1uyN516z9OnbvSr
k1x5WKm2V0eNcuNkKKpYwjnTg+Gik/NYVy696YkvfJawPTU65HvGjGSnEuvx
a2kj7TIg3HTtaCWIeweAySNfzIO4BhNztnUi7r0ZoC1gt+NeRDq2RRPHwCEH
dLNLkhChO93KQ+nwHMoVxnuQZUg5KAnMnHUyik6Y1cM2ZzqUaK9cEnBG2nZk
clX7SycarY6S+1B2RzjqVzselE/69+Sx8l3TFoYwjJ4/0Qttfh4yL0QoWHb5
TKpgDi4VuO+hwdpGpZizBGvkiwbPrDo6stwTsCtV1ao/11vMBiFLhAuaFB3I
fJiBXIrPeFoS5qAdv6L88GmB8rp4B7HSBz/VAHUAP0ct8XTAuew7HiGFZ7DT
nTG4F0dNY3cozH8fAUgZI18lpDRRcfeQvZ89Tf5M/mXeCB2uxzOZUm5XDbhK
eQQa8MZCg+HOWzuy+RJnVB1GNAM7Ca6KFN/qasZ98wlJhavHoWAED5Mv9KY5
vy459pPinCWJTfZf/U0DweRRAi2ToMcRD9wr3/ZZgiuM0CSPkQCHOALZ9cbV
jTp/i4n99BWJiL0jKYyMNMh7Hc5CvISwl6EW0a8IdLobsLEV/DyF5zxhxccG
YLLvdGX8sNAen4QHxdpOfRU8JaA+EAXSzLNumcg09U6gEL4nELyqdUXrloLO
25+JAzCYse68K2rqE8jusuicWHwYJJ5qZ2jmXH68fzcKdlPbygQdYZUz7Dn5
rFbzQWSzH/xl3DxGwc3D00jzKVvOvG99QnMgGRe5MF+0GD/H7t5upocQsJUL
eQGvwkxFHQBcanc5Cy4SwQewF+503nWEWiO59czviTiOnzdHgqCr0zLTjera
x6UKzRLGeL0xH93Z4rOlry/bCxWWvzhbma5KygV4OU26uvtH5a9rXLHm1qcc
WRZQEx1QgnrYL8PUmNMaXlw3n1k/VsMVQVYjVZXIfyDkO5Kc6LXcS58Pon7q
HrgGBx5uw+dzLfazeggutCwsCVzFvpi3PaJ09+oYt6Cc0Zyym1ZuwzBdS1Qa
kRyyDAU9oo60nBPc4xD8Osc/ALcERS5cBXHAErlUWL3V+t2r2e2SAPDRHzXE
dxh2YMziE6trpmRgNqLdnOwDwntnJLdJRZyfmOm3HaMni65giJSeqPio/eL+
w1PTz+uIUeb3mojnZbU2o5xgT/pPDm+/ezFhWqviT3pW+Gjog1S6p5W/uW0l
XS9gPP5YjPX3i0ixyHNCJpsnELge0wXnKsc9emT/tAtNQcctag/b1HqK/R9X
JXtj5d8sszOV63vZ3IxXR1KB+ilpxWJOilEzq34JwkC8849AZkLr74690btm
Nk7Mxndotghs65EdhQEjhY2TVs4+/iMoxSRs+p9usgj9m9Om9x6E1olHIfAx
J05T66FiGpdoA/ZmISBYUKfgtQyBBAQB2r3gV4a8IS7AyvrMJv4yKVPhd11B
sNIsZ3VEdUXdVp6UCG9SsMIbN4VqeE5Ae3iM/lCHdJkDT/M1VINFbaW8WwGF
sGRQ1D7VOBCpmiMOqk5UpWXSsIZsTTdT5HM2gtk3ho0cPohLtyVwDCxY5fLV
bj/SogCPSfgIv3fXv7bVeEnSXciYr3ZNQUJIShqEBm8KL59qsmiG3rVjC3JJ
kbGrwTyII0nARoWX5oYPcMiuJlH+0m19CGHvU8bstroqTTUi9t6aJIdHAZEQ
qOUYkoI1O6HJXshMGuON4l3gmy2i1Ngo4DqjFodlBwoOWdijk0iBkTlJMO0z
ysbSqLt7PjbdxFj1QOS/btOQcIe6my4eSsdpJVB2vt9qgo+wP95l3pdGqzAN
C3//TIiGpicZO0VrDMxqlaI6OucsaeSbr67Dujoz2KAaPZF3L/nT4HrxEeM+
V8Yhba/Eyu0wMF6Des10rXq1s2JqLYlTelCCXVda3gWkX16djmynnGLxFuq8
cBw3qoX+S8pwGNPzvPs0jAl7KjNnR5Ae/EnvdRF9lZNDiHuds0fx+fvHkWCa
KTpUysE5ETvFUe2AG0yXxjfONhdPI54iF0aM9zb1JMATqUNdsEUymX4LrVG5
7mLmpo43GhsaPJPi8Yu8JuXrYTTSBvd/uPcMv0DFv/SC1RH/pfCdD7VW8CsQ
Tu5wftjdCMZqbOwD9QXqLBy+wqSwyuL7y3Whi/VSX/vHPtTWj7vNk2OVm6Ry
YT1hOrVdQYdUC7EZkhxqti224kwAnIt2V0bG28xj/huK53ZVqbxJkphnYHgd
X+aN/SSiVUrWVN2tvOiCjGkYh+Q5l3pqAkpLLsBv9Cas2OozRjhioSrVVxlK
kNy1NJLI78hzezfxxOwb+VXB639GwuSwamY+a13qwmtci6ZRQD/XdQnGFfBi
juvUaYYxkvpLI9rwFZ3tVYIt3yrCY9d5eHpasvWJuCwVW/BOobRlqWI/sqKb
2TcuQK/LjP7b72EYC0P7AEzJx7QpULGM/LanSw44miyVahQBIPtdlrfaoewP
wszYFInew6sW06PNxH5Ybm8/9n6/SACq3CN8SDKijw0avXcIL02fBTt1ZQ+R
AfUs+l2wjA/J9AtSptvYB+7tJ4ia5mxGW4gM7c44s6+DkmC8eXSF2Iam/r1c
1moadScLFHg8SWjaiN/xnC+UOo62HTlx8AKtndTy3BFT0g46e+ai/luAIqu3
oePTYwu86Y3r4bwBOwmL4IHppfKGFZuP04RR5Fz2Rh2fHvlSTCmwOooWvrg3
UjFeRCl3aO3iPPdKeh2zKC+SNYG3om40fFkDWwIYvgDaUlPAhjcHbnBsoZeh
WvCJ3XxsZtWIXqn3mvc5kHsfXSduVT6ZccHaIlWN5USWeSsxF+U4SGDBjTXT
36IwegB4Z25nl4i4yCwt0HE5uxW8lK1JXdJtFEuiC42LwWv96eDgAxhDtFPA
M/o+5JGy2nJdj4HVR/9oLGY75X8NLcXahZEYlZUt0hKneD+v9LFw8361f/Z5
5cPvDQweTMF7jAuybjNNaeG3C/+lyabBZFib37f9yz6K3ipCrWTIE2VQSrql
Jv0sKnaM4QYauutXlk6ffcYkm/15gpF3rjrylr5+W4PPIgsTkpKdaqLQjcQf
TLSeOS3Ly2z6r6Fi8weU+hVGWnW2bhhhKlHSV4Z8jPIvxNWU+XiJOnddlRco
K0eoi3cKRxAgx08R/ceH4mK5+j5OKYRQTIgn+XN4O8dmOePTUebZDsXK31oS
sGjrmBWUAAsMJ1eAVPYo3jN9wnC+LtTUwqxD+FpBAsmrFYjJTwOCMeAyiP++
4BEREeDPk2kq3YpBs3vZv/efAQZ2hPIKaRDMUj4Fxje5zmGMram8rd4HrSKy
FdATniS25pEQxtRvEdaP0DGOk/PkI7NL4KDkxbLjem4DbekybPTOu+uhg2W7
aoV2CSK1jT+Tkg68w82Rivv2wMWUhVho5e6gaSjj2+neCDdnNdRCBJkEaKlA
oWNIVqbzuYkN8jkBz9TX8htaNs78ef4OmSyNK5n2fVjdFloasfor8cPdM3WA
OBpXxgi0h8xwwL/gCN/MIskJn1dKtuE3p83vnn1nUeouXHL+0Yhz6ElJITYs
BrTxgvprrrHssHnpQ3JxsNqaoTMlMrRIy3OhencjGFgAImi5yOHBW5jd9+/v
G1KxSSoU+CKX+76K6Hp+IH97+PLoKCtKXG2ROgj3IUt5nXRL4+isQT8B2zyA
qywtqz5WtuBEAC9hDycNX4/Zs3RZBHeZfviKEh+4JXN+T0bhJKnJA2lYTJvv
8ryILL2AyIysrWtwiNMKSX696SG8XsKNhGm1TTeoUGqbFoRO1KU8a++Dfnno
CB+Fu+efwC3PO8MBYWdxHh5EChEc3R5yHQpF53+5NfXLAJ/eMAzCT+9s2/Is
FWwdN+F32j/aYfVzIAqxZBsYdqJ2f+ZzwuXT/6TuKu+Ehv7XFV9SRXGQArZh
R9dGBNpIUdK5C4OJ1UvXiuZ4JmPu0l6PYl94k6EbcHWlX95iumM+QSxduPAY
P4DvmpFlP+AYMtGZoi9QldN6dZmNvp8toNKgGWBgTOD5vJxWw5m8zCtHPvWV
cbJA0ZW1yQN0fXk09qD4cgwn2HBpHV0tglZKZwvviFMhOGGJ0AfmTRnLzvhH
KfXniPDFxxDVljsm3nXzXFt2fK23k79FH2v8BK60IAXYoReQzB3gIIv88qe6
D7oetAiuyEGj1rE/PTjH515RK8rQpEgwFY3gDrKbY1zhCKq+TU7zlmQRyfau
lTMPiISJEqsQRszy5W79uyUMwf7SSTyrHOm8lKAYtWeJIXfmISZcCjNUeADo
/GD3MSeh9tVB5+hJP7WU/LQEyxPUGN1h0QMQblXUQukRLSlHABUm8gUXVbec
xaQzLOlUQEq44sxZDmLaZ1IBjHK8vqgI+TesJwmxngh4pHvxMipUKTIaTK3z
xC7E8IwW7gTMsmYqRNmRS/FaC4GyPIMOot1mf4eKosgCumRrO1rdAdHAhC2x
aQHrvd/kZI4gm7nUb9DqvdEXm2+VM8l+oTt1DWLQSEC0zmc9oTuVcCAUH30E
rU9g7jMNi0pPX7/tLnIYxLIR29Y5nICeHs7QVkz158kx0vCBF2OpSbIUfRfr
HnGAje+ZTc2e4r7r9ZrvVs/jL9rJbvIgiyb/9a7BYcRwOFIBxQ53XzHu/Nli
X4U1Xj/NJbMmioWPkhreoGOdOj2O2R4mOYWUyO7AgF/3FIxm3d87SdwlVuwk
ipZnS1xzOME3u0SFlLPO4OUsWmK15hGGHb2hupIy86V2rq5Hg5noTiVtuXxo
TZbt0GDr5r3yP57j3KmqNM2Qc+lIIySsTzxQrRtfmElBymoquUtHzJdHfq++
r5RsTncqp+alHXWEhqkKe1ZCMb2HEXaygIDfigQxHLz4nXq7gwvhDgoCblA3
CedgsX/Sj8JZRVf5rUuf1QeE0x28sH5kOELNSRQvv2U9NcTTF1LqoVLOb0a8
j94sJjDIsqm6DAPTZ1hJQRb/AeoYFjjcl6Ai2oGulDwsGWksG5uvhdZ2Um+U
AXBqPnBjBVtoc32r687W/6SiWFWwL0UqNZTgJeQagGMSg/0vYg/RMssr+iAH
joSanzhtPxOCCyMPaaE+D2fRAYOdAlqRwywR+7z4oiLVCZgztvLIVkpIgA+k
C60aeu6FCMmdphJVFY+OjGaPgCAdVdqBoYPyslub0CuTUXYTUVlhVsQ63SdL
+TDcFVPBR56OTSjNfkfGqej5lTOol6cAUG2aphxq0tvsahKVTAv8JquzQHnu
fdkpM0ODsSHXEJYGlgyESITEpN6jnvftHst9DSl+KS/9NbW+j1uNTijY9dh0
txG3q9tC+mG7UvjvoBhSYOsrOux71BvR+Y8PUe+YZIe/Mt7xWXh0XuqxJJtp
tyAZjeXYDrvJHD4P97h9BIHYRkmmke3SalnnlgaO3K6DhrGID4wzByz4zZTw
FVt9/hY+Fu0XRPA9NVvTyysWp2Er0OtFvBAveZfEKSMrvH4sBRxXtNYISyuK
t+gqfrBErJeeV82I0hSjdPn+hk7seWgmLtr5m+FcE5B1upZF3o+Sboz8HDoJ
jUJapsb8LmgUz7sX64QhREowKhY7QCYiF4BXMgEYeJh/8Rfpiz+op4/xc9lK
FNUdqe7tsUp3kPYu0koCStRdo4qZvRNRPytORjrk5XSdcZhJ+No/KbBtH+YG
eicLxn+7WCuHs/+EbRPt6ReoLLOq1iqoETnTpS2O8QPAryjV9gMIUQX1R6Pr
eju1UyH3FyirapMUl4D+HlA0LLFukBEkr8V0tEvp47dG9s3gB+qx/a7UTwEh
aiR/6tEYDM9Agm6HzjJi62CLIef3btH/IRYlT0aLZotz4ou+tDRPtIYkzFGM
NjshgSUpbKuJ5JtnS15FwpB8xkt8y11DZ6Aslgo1b673bIrCzzF3UFvYUP2C
/wRW6bDF/29NZqgwUwkEvQCBhGBKOuXtBD9IAB4nli3OUSDubYlRjSeeE5Tp
085R/k6wyYz99Zrly0nAnW5hYwVxkhWLBDDLRzuRYw1lgmKzf1XXYZi8i9Pb
aMOK+0Fx3RccvTBgEqFKLpTySKptwWtqFrOH6VaFlOnkm/4Ejx/wXI7QrDEH
tzAvmsHpp64C3HbskpMTmZnC7TD1dg2kwsJaH0yRfCpdpDKwxyB2J/SzgwkN
/LseYXkgY2/vQmZDzvu3SpTZCHPdPEDg39+aT3oPz46EfOk6S0UfTbbJ2w1L
W8oOGPc5JP+HMuiYOUayAs6NxE39BlOnvyByj1G98S/CAgJtjEqTxmTmX1mm
/YPTd4l8REKYGY+6vNOGn8BvzBRRQ0eDV5pwgXL8aMC6c9iLGUG8FQr88iSt
Mn61Z+2WCNGeyO9yyoX9kM/EKOwi4QJXm368ciBqrn8lA352f5ADzUtmdnR7
3OVuokfErztC70F8iQA/w84vCoBWN0EkLdhP3bS7Nwp7PWpX9sb9b3341h8E
5nBnfapNek4xfL+UuvDOt/tH01AVx57k/GWqzRK3/KnooYhkchTT8dz1DP10
pcwIwwoIfu9aZpSAx3GkcaL8m1WcI25LgshTA+e3iRH+n9na16+RtsqTOKTZ
CD4xnyvkxqGVCn4OmvJ00+7cNNn7HpRa14xHYXScwQPApn/2F2uVNC+i5d8s
zV91bmnZ/RMKRvxLW91RbtYreMUp6LAJz2i5EJ0fP+1xIq1lWAKMZJvNfY00
2qUj+gIJmOuq8mq3FkT/MS8jPVAyfs6dApoSq9qFR1I062AVOOz8RJs0+WJ7
dmakSu3l5rzNmBuAUPVbw0iQmbbpo0P6mw6I7Jl2s2oj+ewPrJRCWYIfK0h1
9bvCgtrgY3vd+N1ydCEPp6QB9mEb1x5imcIcKxfCzomGJIKyIqoNfCt7mGza
+VJLWVlWkUoUw7da3ZbFUWmnE2tl+utSWGDJHMPgNGi0XmExnAA+q+iGjAbx
Gg6HEpk63b9/BMo5YwbiOtvIwtiO8y5dIA3q98rtIsA9LKi5vHtlZFVokb77
OGKBS8eG/G52C4oudlxIOrWji4glNMYXXasXfHv6jvlgCO6FruZv6hxMEwuu
aViwJfvTlWY3L3J4T2q/bIYEfANZAWPtIPu5CfKmPN4FoOiq9VauHeXrrn+g
qqJXYlYZVL/gOCVNIQiFQuUuLgnmpDzvA0ehWwSggoC7tzNPJ0xFDGIG3jyr
8FDX8gKXk+fBw6dTeKLZLKGeBscC7lcgPFzEyV3XDkW997eTw1i3yRbP8sqQ
BAB8x29Ptnj/9QCYAwyb011JvChq+sRB00kGwvLDDaeCF+10id2VRZWvqjZ3
bHoq5BrMdZnEkPTRMZHTIlfmCrRIUC6w81HMGCFv7oz58K+qg9NUMALSbneZ
MaPu2XJiB2U/g7Cc7RPpILyi7+pEAS+03huNXCuZdPrz5SkvSA3ZTL3kUW+s
TqQm0sIp0OOxd/OcUKxRFe2ZrvPMg+zgNk1942gGud+5iJZWbWPoGadFpsn0
HFSy4KE60RHhqtYIUYzO0BcJje+hjWJdw3j061bWLPtTZCku2vXwbKPW+uEb
eNz/8w42VIz8MG09mRmfeAa6Os2+NzePKxbqb0tszj0IgnHgpXsBZoVZ+IFC
vlBO6NYNEbJ1na0uFGE5sNodNZgyYRzKZxk1lCfOn+ESQRISnquay6C2xy11
jMAFchZrOVlWtLWCkS3bIwIpinNWzO7tqVtPTb7h8es7dgJLN5Q0xGf3H9YV
b/KzMZ18DK8nxT8vI4Q8sF0XKujO7EDjnMSeHCFVia0yQLT1VFkFfcjyHgcs
d/TP8s3o7D/T7KvD0Y1ZtI8OJFxIthM6q3Ck834mU9OIO2ygg7A8fcYLJ2/J
6JX3oFxLekQUumU090L7Bm4v0SVFmPywNmNbKs+u0L3GUf69KaZHQeqnsM4u
clqHCkcvTE49eNpopXCAVyZGBTt4lz4YYgvRzBDE85lBkXZhvKRjRe/aI15g
N7wqMYXuV+uqfObBjhurgmXsq+HAEssOJxxuL56dV911zwgSqpjfehDn+eiK
joR1RXru5S+84T00xvMcKAltXXDKihLbVIeXK9hMzcxpBluWjHNSlKsei+4c
KXlj4Cj4hK1w/HJMPH8W4jYgPC9ChVYhuZQ9UBcdowEugfak5QZaeJhD0grp
NY1DMzjS2pwP1vx2xe3/S4XqR8qBi0aQhROVYTzwa66riSFPr5z5Ijk03eU6
JLfhwRMlwG3MemLN/JHM1qnBUakrKLG4B4zt7sMldxxAlThUYFie4zh+JXAA
X9HW3A1mh8y2T8ZIkT7X+CYdIm2iv6HaAGgRxwV1jQ6dfq2da+WiGrEvTK+k
gyV9qoWv84IkMTGLOswqD7O3bvWSVx9rJLJ119B5lLrO6a+kS4go1vvKXU7S
Hs5SQD1Nm344oJ0qitjAXfhkpVjfMZwwpngeuqKQZhO5IpqQdaGjNPGc2CIy
sUiTNvSTjvpw5lqGZWxdtwjvSjwi7VPvQdT2/rnalfo6Q/bSQUMNEKAUUoAm
nwwocBOJOc5lR7mkHFJ27xVPsP0hncJHLcIYj9bvHQgyX5RhGe+eI2lKYq67
7QW+4zlnqxfRnruciXcUtiEN4Uh6nrWZBrBxf+2vxJMq2vQFakR1QGWLiIwZ
uzdnffrOY9XRMTZf9HT2NekWrEHx3bEYwdrB+czU5ScY//BZXrdgv38DIbIK
aYdJNHTq/ONKxnbLSLDNN7hUtQ5fOgDtcP/NeRTPzREuwU8Ty/hDxiLFYHEB
X45drQN6ahP/ZjvShLPLCjWaav+gd6YXkTMbMnPJNSFhuqQg7c6RY0aJLDKr
f6GoGLOsC1CCW+aJRMDimadnjngPVAKlfV6FT0wDWONuJPTNwo0NF2qUW1v8
KC9yT/yGB3ZtBPAk5ND4SyfIKpszMwEm69bOk4KihUjg3Xs4Gdxmr0bLQsdP
+N4DCc3KjAoJnW5tQuf187ozd4CQzm6MpwMYKfRNglJrcgo4e+AwvMSgG1cG
V5ELYuQTJw3UqeCNAqBTdRSTmXTiZ2t27Y3t1ZreyoqCBFTN9DL/Hd1adUqK
OJXN+9xRxpswAUJZKkuxdE6K2T0bjVynvfgeOK0T7CaNb0m4erhLVcX1OGwm
l1mCzWlaYIXGQeVSrP5u+V9OLqEtrkK34guc3Aj/BWn+jXpZOZ8+yysIgntv
2ld557A+m7vNembEDvoj2dyamThsO70eq1GgpZkadX+v2dKOUliNLwvTnlJy
4zhmmTDVCJ7/Q1b8v2zxQxXIpVVsoNxDUP04zP8Qvw0DG+yFo+Utv/32m+Vt
t3b1yR5WcXHVEZlWQShRtasVYPPxGGuJ3padBVFwltJ2AAkoJYYTBS2MxwsB
mn+gP/80XZbzUFo4Yih750ovzrTzR5iq0FC6jkw+3TidVHy5S/ulGtCGjg3r
E+OVCunoMAUkVJYx5di/SbzAnEWwiqpqSbK1ALj5GszvtLXX/UYDW5QiF3AB
wJb/+y/HrTJXd3LBM9erG8SAhR/BZ5wWqOBCvZFMrXqFa58sxu/8tyEL0Xb/
SIGLy5aCbAkegze8Kza5IdVkVZeQl0ny33Xq4HQt4XHckFBlQy1EvPQyTF/n
Oi0LuFIO5lw52RiZb61F64j7MOEZobt0CDMZ8qmlhKMiur/urm8YEwpwoeyC
RnIK+duEPm88D42CqtF06WVGT12P8JMbIklUX9lGx7gNBksh+sCbg8YE8nIf
Qnbk4b4vGRGpHlabbL0H2vGcnOmFxqjqfmoeAv766QCp4OQAB84Tn0tWkdwQ
ISj7XK1UmQSpdSrK2iyQXm4MLvfWTBMiUO3jiQKbLiJ7nymDfvH8mw65uSyo
Bv9DvL/5aXL31/ws2KEbysxhA/ejsRxCT/zH9o/hYuffd+X0P1PFdu5tPo6h
o1QYatAqkO0PjXmEROwcCaRo/02Xqef651o8R7dWajykxS2Bg0Z1QjTf0h6/
h3O3FMsVypz0SnfWFqdSVpKYc1Xdxmqru+Gnap7+suV1fmpD3iz1ukUsalhL
G3/9y1vWIWYHnLkHKejWorsCJ8pmgnEtveZxVhNRdn9DAsXRvZluyXLFG2Us
9TMQYZula3PN4b85eBr9cJ51FOsOriMBRFp1B3Xoi+bHWvTsYKFiR6NFGK/o
1hHeBhg9XB0BHuDL7FYwyeMv2hxgRWrKTdOPtjuAhEWnx6ETNqvNwX4f2xGv
JKL8M4n6dzzV/7mHZ12gQH0keObSADITf6mBZ3hh+3i2+PTHnZQ2bqCdaEqU
GxxVzd4T50+NiYNCROE9LlW7+/9Apt7rQhYuwe68gJDlQjYb11LT2N9joqtX
XlqeNTVQkl+0jcMgCW+/Q94Kc6pLFU5/BZ8m1JJJNyNIVx0esrOUoSE+gPVm
lpKQ74De6Ljo5/Ft623iAgK3yi957MQ5YsA+uzUAUzqA9uRGWdSKBlHlQs34
Sxxb6UC2ISXf+GlM1pXPmgXHAs/GhwlHx3UaT8Yo1phvjQ9B8w0+wEGfAb4m
/RBeNx37U42XvkXTy5Q4Mbm7hYHZJOELJX6FVwe3czCuqVBUSbw3jm2LPdvg
gVtK4U0wltn0BuXgM1lg1GcUnnIwxzWdx/SEQJUkdrjYRvIcUaI5wEFGWNZH
a2TURRAW75W+PmnTSuqCAZiLsE79mopViOSpt7LWRG/a6HTvggw8tMsqEv+l
ztG8GSLfG+ayOcFk5S2MsZ0SoiRyb3EoirbvddImJueJO31F1iE3iO/qoP/2
+yLzIb1gafLfn9Vjh1/Mvkj1D20E4uDxIjScoqoXXqDB8lv7Csl3d1sGJfzw
avb7xom5xnLL1g7B1CPfUCMqrHc6lTzEiIf3MuJ+4EbMduataItYj2te+USW
LuUAmdCQcIiI3lhlXfUq7GiBfCkc5iUlXjjRQDS2CwehJndIY1MvB02atIPw
/nyAFuhcXhBsPHEQZOt+f2nkwjHu6k/ELbrA+eHXqu/Y+ZM65BrwgMaxm/rn
fjL0o4eexgnpLVO+07YlZ4ur8RN5CvfR3yHa+LTUW1otVxH61qhYLvcAfHV7
ppMbcP1L8Afniqhc9TvJMm09L6I0bL9kox95G0YoTyKiuJ3gcFASAgXP5PET
VNEKK8VHt/19Cu6PtS1sFO27acc9cmPWnNeyiH6Pw1WDi5oZ4j9xfJh1lUv/
FnSJ8UCL4KYdon7qx+Eain43AQ5tjBmJYgnnJPOA/iEXdQAIVNRmnQfoYR6N
6FU6HC/up39tA83JddZCLpRQdTYjEmRd6a7y2/XwOdrE1lnpIXfHtlDRbmrl
+sk9WlHr+eDmbaZwCxU0xIyioM8ZtOSLX+8ghIXta9yywIzSmQumwA1qnYRe
zsBHwKXChP8SlGEpS4X7vy8tpI3OJuyCuOKXCsh3UhXOSVTimTX7OL5LJWxk
OrGCWGgnMJU56NslDZhU5Smgy2lTizOK/dzZdrvJyaUHXMfT7W/RhxP2MeJ/
adu9Hrrw0358/nee9wD3XFZ2UkRflVlFaydJ8xCJiRHV8I9eeN4tK92FqqCT
nvUj0bqQryhzRLPsfJ9jyvOo/u4Uc6zecZf9kCv1Zx/na2kOaUFx5NMvOpSe
KB57AL1gyAE1vy3d0gGeBMVVx6zHFo9Yn2ZvmoPx0GK9HHsmayqWQmzkwCTn
ohBjnfRzahixrakXDeyGw1JafUG9hsJMGtOlc5PpLG2q+q2Nh9oYWpryH8K5
Atv6UplN1s/xwAGkiLwajgeqb2ClpSzNMlc/OXw2xmZ+4sq41YlPhe7n797G
Wm/YsjlUCGeygteg4IA5r5RbkomxCsEXLx+e3ibTjETlbYjvTfvSGvm+KJd2
IQqOa6un8MIo9Wsr18UsNKhKS+bqmoyaFnohDAjP6sNiiwAv25Soe6nPNQZH
/XyXDjBEmFza17K8AmvD5GaUnI20HMjczg4u8hzCnFYZ6S5Hc4gPOKR07gXg
ArEy+LKVjDgQbYFP7zzuycmzl+vrYdrAqlAks/J28JDN4569Mik4o/DyqsPc
qBK4CQZEXyqHpyejeG9z/7qKAM2Af4/s3ZjV9aZVSqVQWQwjOnhHm0/iQ7lN
mpNQBzQiG5aIRTcJUD1K0u4Bm2Xx6c1yGVeSkPRSX77M955YUBDwmbEoz3Z2
xcp/s5ig33IWav9zYDkHYAQMs1KCwoY4lASqZgltoPnHWJpPrfmwf4/V5kXa
yW6IV6QxZ7elj9PfXJKyVQ663AITCtjm4g0C7gg5mXmQUiCWa+hKwAIuiCHs
PJaIWX5WWCrDwoUaNlwrk4cXKLamz9oDdkuyQNBxmztFVE3/KGyjd3FSdtgt
xG9KiHBov1PYWWEvDHVj2D2Z9E/XBLxtyEhZy4prXWeO1MQjStgbrQvD8sED
qOxABwu9cc4Liy2sQKFaFH8dfu4jGskEW/q57xk0b9ThsLOaSOGDWwge4rtL
eN/ZcIRTmqKpA+G6N41/oO7XPlBrgOD05z4w5lRAfjpWbqgBCXCb7EFgllEG
ATPXIXJC0XGgRPosEj+VGluzZhv9ruSnGU5wXykL0SaiMjAIbD/h54nvloRu
RO8un6TCmL/jBxoGSwDzGDvXhtwajn58PikzZhI6Zrx+f4FP3nER6x+bZeZ6
eAq1aYFoOC/hiPcJxsOoVLfNMm16UdYlWBxZNECmjvfK04IiZwbMe5a7jYQX
YQ8X8/isVmWleOKrmoofQv3cYpi7ka84eQLGXvCnSyRC7F8oWX4qFET5D101
T/d3JeWzBUy+n6b8JD696mkGheEIUho8mxDm52gGO4ABiDXx0d2lg8S3wuzg
74qMm+SCqnl1CuozwL0ZB2XwhZavXFxtsEm8lCDaHjKKqnTE9WFB8VAYWNzu
491tRhTah78MYajMI1UCIrzh2P44qnkG5OSa9KT9nh1W7+r6JQ0d5MJFuniD
/N1Eo0XwNj5x4NL6fofYhmUtBnADrIfFlVoX+2zz4OSWSOcp46x3LSP6+RdL
wMADf6gQ0Q/Kezjq9o6rEhlV/VkbuyBYudmGUO8S51Et1qW/yijaWd61p9/Z
wn01P+n+F97cCZM+fJlegA4APqsjcmtAahcFMDN+VbRBkZ7Do/m+T7EjmwSi
fUekgXoDtInfdN/M2pj8udRi7VYQdLJOGUXFNW5Oom3eIS6MDcTMmSIbkvyp
Z+HcRlWX4EJ3oJ59GU03O60x3Ei5ie2/TpZxG+DSZ2hJbAYbirPvsFbEuikB
YMrvuec+hFquBkRFys+FRX9TYF7DI6/Mdl/tYCe8SzZS2HmBHAcKH42ctT2/
KR96A99AgLIJqjjEeRGCq3H8ortwNpKVSrfkav5579myc96jlut2xm0yuASL
Jts3xo4VjQQZ3GZZZjYcxo8CUTU2+iEqVyCMNkLM6hgH6RYsT2nAt+wj3NQl
KI8bjIeXZAoi+a7/C1t1cNNh5tdVJMTOcE6tAVvI/UJngk3xYRZ2Wl61i1F4
N6q4xksmJoCeM04Ln5YUuHJhRqQ34QLFzWRy6uj5w/W+6ASbgqte26V2Q1Tz
YlEr7lsg0xM9iKbpk2B1Uofg1RE9Zmfu/LQTOHxAaTi/hlvFKvGxdm0+oM0w
u3CGv8P2pWNUR0p1NPcLsL0+CIQc6ZC/Thxx0q/X9fXB5uNnk87DtrHRI4Wn
mBjqKm3DQd37QE3ZEEca1v0+fH9tMjlUrNNbCdujgn+p/PE2zbzPiWoGCt0p
AEPRNEpS/T6KeA9cZ3ODwJwA8I8dPLLx4E/CR1dY6x/GmNi3ZbyxLcOboXck
lRdmj8WZHXsdPczCfHZPsgpDGC+tDdmSZPfS32z/bjVgT4dl5A2cNthCUBuw
WFGpX4NMDo68yKIwmTauB8ZtZuwgLTGT47GOyFBUnU3c5baycO69cWGJVFqX
eqErWu3g8ZC0FhybdT4NilaGWE+5/ZFoQ/CLha4s17rAQi364b7VbT9ED5jz
jf/m5G2KLBtbvAC1arGExQ7NJE15gCe5L2fcHAPVviEn8YEIuTuATa7aayqr
Ax7ROSvTRYaob47+RrdF7+7EvOA4KlcTLjYlTV37K3Tc26KKcuQSiNhY3xwU
nWT/sZF3jIaO+5fdO35XECiOJgaGhJEp0VWqGkFnvay/erllBBYyQDlQIFnq
q3YorC1ozlCvFQ1kReAZWvQobqaZIY92yKZfZssehFGi9fRTfFPnZyAuILPJ
4f73K0GtWINph8Lute7M9x2RzSHWfsn1LAacjqmArom3rWgaf/oxJNTngNUt
7ZsK+ShPkNCXkTCuAlFvztMdsaLtbj0WyuFMXaqfk2zbUOkAK+i26ZxMcJr9
UwhvbW5wHQJrnl7gmLMSxHa3sHPPYpQvbj3GRzaxckc28wjpwz35kl8EUq4o
5M8tlqpqeMENDohnlnD4hDxJWpMsHIYO/XDPFWcI3F4fT6e56Al7ofzcBnxJ
0cG+dbUHGCe/cAiAk9CmHq0zNTTKdssokRHspUypfRj6P3iY2q5CnWM4MEO7
Z1BDz4bPucqbF+F18V1DHaKWMaGx03dIM9l1F/onGcmm8fUJ3ttOvEmgLdhW
IbX1dD/pCQPuC0z+z/x3YC1ziWRmJdEGrhWQJsWCBk/CwVTxbptqWNNWo8ea
hv+o/IKNIi6zySSf+ZVbMaNHZIwqrcOQyNrmAPqrvmUZ04nGWAylnln633l9
KNHKMNMmWk1HGOMdkmhZPDyi6V/ETOKgqrzlx/Zc/8w12UdEqt7ezuh7z9Rw
TuGb1oLRrsR/GMh31oV2cH9wU0eMLG96XZ/AxwGcW1jXVA/qh8ARX31mkVE7
Yyu838IViw1PoeYWcQfLjBu1aIiLmigQGbtaHi0wApq2vPwK+wOBW+vqfqjC
cFaGPfByIsXuY6mG6ApvpMgms8m0uQFgJqZppCUTCMJC7nd/pla5p06vVTKG
9MYeVsiVpD2K/oQZWF6nce6rycm7uzxZJeH9yjFNY+FtOQ5S0TbbGUqOxHpY
lo2LRdG7M466dW3GRvQC7jSExoptENDr2rbvdJHHeHN6kH1AgI8p0XHVOcQ9
tO/T+qSVMZnkgjg+DFLAL78zl1Ra9uZVCtMoUvvhpW2DsknoB/5oVrSM/gpr
/uKVRMboKIHMtFg0QPlzh/7l+o/sQ0Or4vVBzUA85vqTaX1sX7zvz4IDuuul
U2Odun8SbZHlYXTeBbuZN+VSQisq7Unp+sv316C+0C256KGdCuEnCB3Eojtq
s674Y+jW9bvGKOJf2vFw04l8NfJc5l/EhtNvyLPNG7+oQjKj7bN44uK+rRLD
7CZHmOWW1V/OQah8OQ2F5nyotW33v85Slwjab/SUi+iuCoeoIDh25oTo7VCP
/7wjM9Jr5YMoTsit2h4M0Rez4lyx7eH8SotpziCPt9+LjxeBGEnNCQa6PmKt
PZjP/qz6+PLocasvYWBmaaobKcBuKVjP9RH2zXe/KdnO41fWYhJPFPE8BZAm
KL2gnHgfjxOgvj3GUbC3oa/4hj6hU3su7fzV5yWUHHEOtCgR4kSZ2G8IBwvm
dz+Yud6BeXngqZoNhsmJPasGOVJsaBXmpbusrECkY2Ki1YeAw+nZEQG/VhX9
+u4D4v/o6/HzU/z2ue1Ua+d0+ZQKJ1e4PKtD/i364+vT8A3FqChTaT5bTTFk
GJwHCfbqXK4dDALBP42MB+e+8f9Pf4rMhdOmy23RRiOkhee6RjaJ0ZZPRXsM
CK8CPdmnG4CWgiMNkzreckQhnyTs5stPWOjB4zM2vhN2xOhrCsIFMVQ//8zw
5DY1aQc/+46OHeI+sDBLRdZjOpLxRvTzspCbtxSIs/fNIJ0vXwZPDWgVKrR1
cWG/KSIUSVs6xsZnAKCBZxbFTz5hHshLCTeAuiikDSqVGEUFo+Aav2o4tnSv
LceVKrGACEaQzCmPQ0vFJtgONoHXyOBRKWLACSG1Pm7oI0efX8kXroq1Qvt+
HiG2bE99mFdisrU2qRVqBBh4i8c9S3on7UzzW3UpnW1ZpOJehNF+Bp+9gFgT
oABGl8IlzNgxWwoP8PbOzXunGDGOsc4GObBAPvC+b1FjIoQ4GgqDj4rEhyO3
CSHXnv9ZVTrqXn3+v2p8+MteU0l98wVkBZEsp/4O1JepOilwSEVKRmoEVh0r
iQ3YoAzfJhchhZwcbX9Pj70GvBGAMsUy0oxL8xU98EPgrdhvf9Z/ZjbeToGR
66hQoK4/0j7GA5XZBzPv0MpWDg+CRM5W3yJF4fYIUafrc/Kit3lWnjUxjCFA
JV+C5PN1fvabbaRtSVB2WoD3NPCG65XNMSV92Ev9uaFRu6jUiuPBZ7CwUEOV
3dOX3US5xVt2EYYoI53ytyKYcIoJ0ZGkp7rxjBAlFjx4lLZwlVtTWj38P1Sq
EYMq/puU4UhABTPagqd9tid4y9hylp2Bf8GvkMQy/vQDZkVPrw+/zmoJ9/3C
3sjsyxd+4CKU5wVxXYOc6zZV3JhY40CWS6+HsiBl+r1gJ1yDrvVsj8rAlnJB
Nik2izKQ1dcaE780zVEw6I4Y5pu2NdeCGoVgoHwfu4VJ4ZiyjDPvaUqovQ0S
7/jeO4xugKTBUcaUJFC7Lyw+Ij/jC19/AY+fazGNhegvLi4UsSQJWzP+GcyH
apKAcmeksQyGqxindWrp6ZKLEfvRsCSlikB7Sco/yfXRIWU4i1miaAAFZl3V
001rIqjeWIIJNKLyTbmvp0jqkM6mwbbN1/jK3aeTA3C+9wyOafdmvKehkpDN
8LhwzIldsyw+Hb/bicF5KzL/PZv49gv1By83qV+K9bH/r3QPzB1jtGFfPFUG
3Qr2M/TTc35+Sg3bfnPASbA2ZD+RTuoXKF9JWfp34d7/jKiA3UHPZSAOPS9e
o8l1AQ7UpGDw6IstFTSE3hachCmB6EdIdY0BbR/YPoysxq9VimP0C6y/yRl9
gJR05Xd/UXrwCRuLspH3yUmpsD3tVsweebIjZYoK2t/ySB6a58NrMGIOj/3C
3aufQ733oZYnqTcYOOt+L21ToSy7Oty4BiOR1hFxT9ux8kMoeZs1no07Yhtd
IPgQBP3y12uBJNmKOEAEZDFFYnimRE4SEwFYHgdev2KSEJcxpVSBtH+dzHWT
oezrddrqmpfDiuatEUW8uAj0RcSFUTNSWf6Whq45tC8a4/UpqaEpcIeHj9zg
qkfgcMEJzvPmutpNKAqEcl6AcLnfLXVRevm/GEh8CGA/73pZ9Sm08qlqNpQG
Xu3yHDslvjJOiePZh4iJCuVT1wFz0Ui5zrivrt2sfAzOwHIvdLnZ5lwa0GNW
N3JM8/nTHPBy+/NYVaiEYSdwJUH+0EzANxYVAXB2OTAmJBy67FIyRk9kyniL
avM8cDHkbrjR3R/g8KBa+RpGowXIsWV1xXzZ3CYY9bsfDmfaWvxVjCgVvo0J
f8mZMFPGN2fxg5qwgcWB65M85PJAMtmdu/8NCbFr5C/MgYYCFCr7clb7Zprn
au9xrZxXYwDKwh54CrgrVmH+wL+cZ5dqZrO6yJ32of5dxM5DNccvo/gUlWrh
LcYk4+tVXB7E/iSFeVED/bOKDqwyAtj917s4/MJzebFy0hAZXXV9IEJ3Rfy/
+6ETGnTNxwwViP654UxTWao9V2ea+TvGIgwrLdw+28HfuQoWtpiSTtGdpYlh
+7S8Mio0AvRTLh9hYuZhjFEYZ/0rU41/8WNgvaMXSLsfrqwFc37O7GXD7fDx
aoC5u3TukLKfUp9Pwe1hJ5TwW9Z5N3kUTj+Bma8zFVoO47j5r7fOSjVsziXw
wo7RvzQDCBSMDhJbYJ4zwHqPSbT0BI00y3GxwTmgOwWYs09RcDL9/fjfKV5H
y+y7xZXmXnq3auV+xPNJ3omdrX9YlEFbwjYyrtxM0VoB0/ba6uDMzyqeieS5
EVSPL193Q7D1xduCUCkioc5aYawoOltrpnA9FR1Wu3+BgzLjzL37iQnDbApE
PkuPd2ik8LSS54APaYvdTC/5MWNPthBqAbiGwYJztK5MVRN0lkHNWiPC17IY
921qhq+8tDqmXPbRLQGEu10fyNcHAzrJ++9/19f4/gX0oS96GKL11uMK+u9f
MdwR8lzi7UQgGpZ5WsEIZnw9GE/XFYycSo/folsOkljD6KTpWCsuo41bMh5k
zYZM73W3e2JGR/LsmqcHI3gLONWNC8L26GYIu6xOPFDbVrFKJux48Hh30ptF
2zNHWceUqMlUqXU/+CANbq7xTeo6OI6YQ8lVE/2oa4jUM2sPYMSAZDVNCwuH
oyNsHEt90gk6XEgI+BsMSuHR7rPssBj5rmqeul83vip3paMEA+sSPgrzeOoO
xfSAsmUCDniIiBp6vNcjwwlPWggOec9KoVkFHzaLA/FLlZ/RnW9/XFJX1KLJ
UMen7IAlJTNdkVFBRawGRXOIXmzLUTnmnSTJRdTHnHaIqL4YnR1Xtu9Fxt0y
XxzUU1JSZUSuHuJBwBnRLOdkLTsjgkODxKtr/pHWcCrXX5iUmtu0G8LiDaki
kyaJYSUgNUHhZBjBKwV99eTK5S4erWowyJVCBEda6Qt5RPktaxoZRj353nSs
SBau1DUMN77ZUdJ9RUvXL593XgY2pl+StVMqvVuFshLTDRqKv/pgjs8pVRLc
5C903lU2WhnTZgGtTwojKuC3i+30n+SX8XfIQt1b0rOd2jcPxxYBX5Ud1mad
Ed44fGMXOB/CSkR9Rw1FliXHZh2VcbJV2TJasVu9MYpNa3NBVJkvFthwMxFA
FVNQgttmyYPtqkt4iOROlPoRnX1zKazAAIeIlDeZW3VYiKBJSzonWTDTbDt7
Uwz9KGFsuQNVmPMtRjYnY3Oo5G+r0pdeGKR2+HUmbbwm8Dyvp/j2Nszfkar/
4DOj7WuWAFcY/CgnSMarIgJfX7cDMgaEwiIxKbOmtcr6Ss3bpk8nEfIg2MKU
MBJvQiwP3pxZ9UHbw8Ds8CNiMjo1Ddvvi9dKYO+nM638WU+OQ1alM8Pk4JlI
vPbp8CxuciTQ0yVvVdsUnGL8lBdOa7X65wrp2SZMJRivyrojOiV1P5pRMRa+
33lFa4ajfKT22KhMmnF+gZ92RLlce38x6tjsDntoIWM2tfZWLXt6HAhcxJ9k
dDQsEXZvpLc/OT5MyNpKHoygfYdJ2XdLYncrXbbR9f394y5/P31byzKcCPuK
kNO/zrTb7fjLJJZUans6G4BItz3/WmQMiUZBccU1tS1nSp9K3vCHYqVOwaR3
PG/GYmBxBeIzDFj7pwQJ4dplf5gv1HfA9U2LVmvm3/sONFJu+yOftio6Jpz6
G776wBCI7xX6fcuWH1xqbFDeM2JiWuU0NEIqhXH2kwNWUU/38r0oAJj/LbBO
CRfWhTMT54SjmRmyXiziMHKpP8Ac4nvuIWhAmnFNpa1t8RPRCc2FTP/UDa3s
EWR+8H9lFBz37jiy5S0+iNN6OZLG29wuEPXnAUTlJsuv1rodfUsUktnkko7o
6Ijv/NxZN2eh6I3wIJZ255cWI9kIr8SXKMJ7KGJqm3Ubg87T+E0+YFVqFTJF
6kOqb4A4vFldv4M8lcI+DeHN2dGDfF1vm3Bxr8zV71vDxz/2Qed/snuHeyv5
ldHxzjYyrPguLHyfqLzOfJ+piYUYmkyzTnU/V2o99T+3zPA/pXe9XZYaryQB
Z4ZsnOk2FLbWTXSUOHjocGaR7uLpM/b0xOxg/Z0WSgQxKHdNHgoEnIxMceTY
yu6fqI4JxlrAbk/yKrhMYAXYRcJtKV7cimNPpCKiC2+piARJYqXWEtMfnPvN
dQ27/j+jzEr3wS1j+gTYwV+m7abIKt/RBig9W3ioMruLSnQrqq8LVgU+zMjh
ibLSnacoyadF87cZRE28ikKMpUd2b0f72P3xOzUKPxJ0RN2HCg6r+KFBU5bP
xaAwQSbQvQBu1tsQZIvl5/lsn8/RznNygwA7lEbrFUT0yoREkwzNla5vDKhK
ZQL1DRjIPH7GZdTNjj0q7U/uFUFy5LtNQqdPtLyq82XzYc4lrDTnBYFGx2Cj
ZHbguUzd6JtX8mkC1NBP02IXbdMQss3iA2crlGq0M27aY4aTHVIYa26zgA4T
ifytFr53pnAuJphONYWmdfr4B71cdMd80pbimYBSu4RO0bvJoAMjQH3C2Psy
Py6P3mCJ4wHuK+Q+QfGhDXdOBDQKiniMhpWyVCrXPOTPxjU7GfX1dMmlXDXX
6wDzeDm2eVvxFG9GN96h6S+ocHH0snEuTkGHAy3bl2EidYGU70cqWgw0D0cP
wRYaHX8PxiSMGpfWOp68OBsRexXJ7KGcLcF2Zjhj6lwRipYHTV+UcSkSPiuO
Yq8PQRBgr/SRKx4g92lCcIvbhRNCMn3iMNekK+nck4XAsdOjJhnTZzOJA5ZX
VUbslOhmDSwIoE6QXnFuerrvNcuqOQccbbx+trbdm6vnJoBvtTo3dqbRsx8+
A/KnAn+a+KRvqD4/BE5HjCKwqBaoE0/0X0ueJtDkrWs1lxj0bPMnlk8MulZA
d/4l9rWberGr09ZLFO3WOPnyMLVfeqsTJgL1UTClRVtE1e/N48i45Oiz/onp
kqjDq8FGdcfASE33662JKrxfjJQvp79atlHv5Gj8bx9gk015Nuluirumw/6u
pjzDFvG3pkA8xf1TwzLO2xKwpmMaxe17n8G2DdNSsXvDeUHDIibLoV5lbU8u
qPKF+8eXl3qLLp6G8Bq4MrV9k+B+OrYD3qybQD3Xg3OC4/KSOB8hfYtjkWAI
5ruSWj5VZbM+5DBgvxOcye0q8zk1O6F39JYikMgQLHOB9qdE5XMKLmyR3gK3
fOs50E1KTznrSkPLV6OjCo+E0OnJ8GC4+vUZOcBgyBEsza6HWxIrXU7Ypyr+
bLwEnTl2+swkslMv8mFOEzrlNCW2hymsSYel8rsHTTOuR1lQC40Bs94gQ9hH
8nioDrGo3h3Fsfgx92XLT/ubuSV9O2A4MzgHa/N8PPcRi4bxYgXfxOqlgB89
rXAM8gMUuAxEJsYBNrPnr0+J3Kf+Cqt3sAG/C+tbd8lsRYfgwY5EezCyfENw
2eV/v0nWm2Ycs/DscX0QbCGhOD5OL2Fw5zffoeDm7PW3PkVb/BZQvgaAxdBS
OmxT4gqqIz7UJ1Cg5FeDuNRW0I9oivzZt5bGWioKGg0MwUfuZInWYzqVm99v
1H6wMnn+Mg2Ahr23SicBNnc8gb93uwL9/wu8X74OjhkrBsv6hcO9Adq5l0bq
aJbSA/DxnWXoYcbLqwelwYQgXhS6WZ3NS123CoCFGx2Wz1d804B1NSDKxHZi
UgRzbEasFPMFi7S1+M2QbZpanPTPz85SGWiX9LR72nMBLVzV5UtnPsSFvmDh
QN3BbXPZGDiiDjoqhg4teySk5VYl4Be7+ZqI0apvHgxb7flE+IlOimSn9ZR8
9rWnRN809x18ogBOTyWb/1Xmns+d/ywt/dDR8LkPcKnOs11sRmUMqvvXNMuI
ckmV+JMRWIR0euJjvF/qblOWBW3pGoPUoKOsdXaYxd3p0NKljzYR0c+ec4me
w2Mwad80PDbFQxoz8CXt1iOK3nylmIZv78o5y3/7Gfb5dKTQJjzT2Ch09ybY
Z/KjoWKRXkVW0nOha7yMNjs0UYKZhuscQsaa/pUa0zzgi/Lpm/yVYeOj0enB
6Vf7TfeK1+Cqm76EUjW9zEg+TctBqaPWtA9aJ+rX8rJQY1T1yjOX3UE51i2P
+WgmTtF3fYLZIXs9Dal/OhhuA2SzFuKn8Y7MizrOyQJ0TNe0w/pvoJlTvvds
pypBBxygyKmkLtYQPlSHhE/23LoXojkmJ70mNlkMxdWffkR4sH2UNVAjJ/G2
gwAJSCn/TY74zkD2f6/HMAt9puSRXTCaQbs7yP1PVgxhu2I5kJ9usfDEcV5E
mkwEUD+UCTDcNv0kn2iF6SDl/G5AheVyMJ+XmRFSUiSjZZjiygF7UtXAPsq0
jtPZOnWib/qQFgZSjxs54DieH1dBa0rLfNWFAq357Mr++bojOKfmyxZturma
Pt7WvcvuCsggmgxZdEpp42cnhNXbL0DGUD8koUfdbYQmgQW9kP7eMmjAq+q3
GqMSV8fQlYMV/yWtGbCzuSXmfk6pGhlju9CMDKsaSRoRedJQN0Iu9oPBv+1J
hDvvUGzD7fd3sAGY0YKox+hYpTv69TCwL2wGEBz1tlHwDpntCaCEk++rAyKT
4xxOMO4cNefYiJWRxBF24w4j7COXW+IdJNFIUJI9IPvCGkNyxC00TbZeSUcr
gHWTsc+VgQ4gnhF5s9ELocB5OC1RIMYpbfi15qeafesKu6dPA+QIjVpqkUwg
MDDN/SfWnbgXyAAUo5PIjzV/HszdwaL+bM4v9RzHFRs+TxrCQVM7Jyghr2UC
n2cpg567t40+4+tMpEg8UIIkZlIhCuasgUBtoGAjN0kDe1f7/etd+q3l7xq6
g5rX4EUhK3ysv8X7Ac2FRtNrpPJvFSFugItrZEkMJifTYAJBazSLPB3+oNc6
m5SSxMzBhs57BmQ0QWX2vdXx/GSMKmavk2lJmyC5B2jl/Jg5BaCYws9BKvMS
XMPR2tV7WJxPASixVqUBN2+hTv6FV8jOkUq/QAXjJ3qqDoKtS8xJrFMuB3bD
yLOcgc7AffocJq1B0KEJELn3FzPCp4gntI3txhEZZ6rfSxnulBacGxB57bxf
NcyYWsicokgwsus2wj0MZapWRGKNXRkMDzP86z1Qf8cjr8JFQ0Ri6XcBjlFB
FZWNRJ6qgrN6KYUlHYUJUmHi23RoXlmInl5XOPcQ0L3+54sNrXnAR/wIIqKo
BH5amseLsLLCkVzj1OclyQoRqQ3oGUUQNvYAT4rQeYGpM8S63td/jLJplGNj
/sPTKPI/ihrzoAgcdlvmGXgeRIHuUql4CL89QKqc7S4pd4cCta4ejEyg/xnJ
t12Ze/+Q/UlM8gLFuLUtNRAcBK2uOwl6WaHOkflIS8fFQOiAFtO45H+F7V9j
HvZ07di5JVMJ1M6XN+7VYISHQb0skwHzGJo2dvn6bQ0EphgCfPKa4Li6z3ll
QJeM3io8f0yMFyfkBqt/SwElnv23GWlcHx3ecxw1Kzh5NhhhLUoR10Z/9pqE
+5fP9v+i/k2+U/5ns3c04Xq102unIcizT2Fv+K1M275+MLPhZ9L2S0w4b65Q
VdJ9TtzqXaAqk4pcBuq3ffcKb/itZ17F9PQdcJ1dt3xDq/AQGm82PygMySxl
fV3v75r+xx+6W0keyfjQ5BKFF38LYD1K2b0iummRh5rcVuLAB1L93CLGfnYz
vdo3d02wba8/4H8uSIO6E3uOeBb9pqLII2BkFvC4GmBovRrZp0VEFKZqXpNN
mdib8Bo1Tc8spcM0HGEj2gRXgdgercrsmPoL6XDLOyIa+kEWZkCU//sDgsNi
Ivgbu1XqxjYxiQy0QMmcw/aUg9uD2UHWeU1CYRKLSJFoyu1MV/X0nZgmZaFy
YjMAONAg7f34ZGITA9im6iJ1i9SyvZIgJhND+QLEc3/8eo3MfAG4d8JAgaKs
LuETdS7C9QM5UHCj+hqz9NllD/rtMm3HfsTeRv7DTbL2ZEg0T3yNm8NYCTiu
s3MRyfzs4oItPv+YryFfETNkpuKCQWgjqN2KEzKzHlqxW5pymPTQw7w8acH2
jfnogvp0ux+fZpK6qgWWzo14sxy/gYwdIJExZ3qzXNcfP95BTasfP2Lt8szv
PlR5cJCnUjWNo7k9wPeH9BNgSir87LD/qHTCMmmquaxlGoiLhvushqekVvLi
ZJPVJ92wqKc34ebbzlGGY9R5ROEVyh0DZusnYE/GtS60c/V2Al8+Jy6RCkLR
PzkAhxlRjXKSqugdqswdD9SVNZqu2LcL9P1yjtxovxNZ0YbdrT0zJ53dcuDz
y2GyZxXY8op42TCH3sjGG/a+UBkqudXSD9dv9x3wkTHNjh52cCV3mkIu/QKl
Y+DblOC+cQM6JV45GDuY8+lAHj7MHNCNhzxEL9OafdupxUPBVdo79NRIbNck
DwLypNq0Shu7EwDtZEauNk5iFx8VadPogaCi8g7ZsT4b+RXhB68hg6awzNJV
q1VR0VT3fUbV8FYHzAhdV1Q+m1tCXEp5rrcevHjGTCrrjBkojoCa8cKbSzDg
UHobH7x9HxNQtbFseK7KfYpsQQFPM3LBNBGkAhrqwS98V1hjicS2OsO6r3t+
pd4bYt12+mtaQBG45dBPfkYB3oHOEbEczDsA/4q1TFR7ZI2FdSgkxPt8YOee
Df8AtTMWRCQAL81XkpQpdnpJB7ZPXzv53B+CMhMGQhR0uBpPWDthSJVuwbg9
OwejYbkwSUY2ulKZjFY2djvYtmkUptU1moHlmqSbKbKS+hkIGIB9ldo7XR8w
uVyC8AC0JQ208Jg2XDlZ0aBlyTbrQy5azL5bEf6bV0bLkbDrTmhIhqyxLJx2
RUSOfotU1NAX/0dLObFuehcFx4pV+Js/UsZM+9QjGgqmZrz+cDze+//VEnK7
Z2n6zCiDsIYf7b08N311FvtDCgXDzDmf8qdtC/zAzMf13TLv+FQ65iZsyEfO
FEOjhSCNpqFgbSuyBZEMbVXsw0B/DTx5T33vfRtedOO+qvA+kFK39ooCPqd/
O66CA1nAPUv3I+Qq99qio26jLCdjNzsmuZIU0XN5U0r3NsMXsx2wN5tT0Kl2
2P7vT43TmnE7IVufGZPwzcuREGGT4lTMCSAnRBjiofKKKSq7I6zt2XmlbQqW
R28YaYejw33FC87u9JNnOv9QOg58d7btCK3YzbZfXpLhElh1rPhHt8MiJFEd
ytOfIYyAA+FqekjCFvDe84ADpi7rCr3PdAKzB/zrFn0Xa6/7XQaLVVbz7JTB
xJHhNtAzXCTU8bkuSbblD2CNlfbQ5QHV/UC94xnyzPntb9JlxjSsjUtz4l96
eT0P9vFUbXJnnUdf8M4fKyabRD+taQeorhCmar4aqewsa+p35f8YkgePi9BT
ME+3oHnxAwu73btwoOlhoeAcfN8NWRqgPl7HyjPc366me/5ro0nFJvcFLMoF
KHJh2APl4zHSmo29R5q/OU0PbR1q41P9FB0TQbhYmbrzLddVI91UmDsReSM+
KF7P318tgNeRp0ueyA3phzUzVRb6FcBLjyhNhrF+9ZbAxVkJ0395hE/7NUJ/
DxBabG8NO0rUmWxXBZ/MqjI1aAsEgwAdXpNRmgFXb8HLWIjW0nLezxtxXBqf
b+oRuwVtCTAutZ3FQo8s0DycrZCDEPv2UZdXYGvdlj7cEB05jzp8h1XRRFk3
Askeuvko+LcHGlMBEwb70uxQfpjBOhumTBsp7VVLzXNX3spn3WvHE/QAMpaK
zIZ4EsJRKpQMUx+whKENXgkRWKN/S+z0gkKhScTH2FlwIde5OzTnDDVLYhK/
houbv1LtzH1afef9E0lnsovpjY/Wc8MYFX04muOdUJCDRfWBXETxuQLYQO+q
pnl3LjL49xi3UTahQXhzclidPOe+ENvmH6FepmSa3gCgzAdfFOgHaImNAKOy
NGYd2z1FP+8ytqkBwKENwmh0FZtHDaQVtzU/9hSoS4GeGyRNn+6oX9xCj5gv
Dzk33u9sTz+fwxX1cdC36G7abc8ExHFFsuRlCKJWZTQiCF2IV3GLh0PJ8Cjv
Boxn9ppv+sZZlD9xhOYRSzMdQGn4XiSqR18kzbyu9a4p4mA/JgM3KaZDzMUj
UkGZhZ8ehvrUAMgzNpyeLDvPSJnb5Og4tX0SGyMvEZ4/JX1cC01gASyEeySf
ciB6qsPWVTkhbUX3H5uVkrUouka+sqy6k5hORjm2U4eN6zPKWfUpJi2VyD8I
ZBvG8TSDHRU6ktD8uz3qcvOBb6ntNS4XWNtp4t3+dgfNGMjMpIR+tCKJw3SI
nmXkx454VxHg/EE5lU72i5nua4gUo6V7RoP6O9h+QYAANbSq0bj2LPm+4L0d
nZPRrOJcVtLUDeQayIwI0z2e02wxC1RGsJ4JLI+20ZlePMtfbRLagiGtYCC9
fIUcXZbJ4OAt2KdyyRZWgcQy0Fg4lzYjALUHTURz8h4mfl87LqVFKkpTLcOg
1LY6OWhtP6bK1ba2e8Rw+AYQgrF9n9vuR9/Wujmsbxa44n8Lq4FwmF5Zl2ef
n6KyXP6vnzloyuphb3b8cWy7fiJLKoMYPG9upUyeU4uqrCvB24evLx+sPy+0
LB0pViTWKCsC9s+i/xoEYOVH/FYY/1AK8WbSqkXr7p1xeBDsu+Wo+7AWGmq1
BAfuMK012bl/hokw71jOR6eW9AKG+xSQqQWTUd4S0AkVPn81qWYv5CLTnqxq
IJycDFRwaFJ5RypIp7QFF9zQfLMhbKG2hGegxu6M726XLI1pWpU5QkJbqg30
o9bpw8jcVP48woTeVhZc9F6FDgN2efLOMQ3cfTTbOEoJKsJkxeidHNPl6qxN
5R+2zX7crar+ydl6gWmkxKxYG7o9DzVy3dCYBhPA6r5DrsVneHVytZ/pxV2a
V/iiz6Ci1mDVkuQez83fkerh74PYj6vIbXke4QurcVv0VrsKC4NA+kUFzlWJ
r3Ju9uvUBB0nb/l39cZrBwLKRMUyPXaV1jyoRdZShKioKCFx4Nf67fBpeBDc
OOMVKx297b/KrBtIIHGAkKaNgiNmGgYaI1xjJV4mAiCBo4oSiAAz3ANcQRMy
AqbfT0obeivUWRRNqvjkt7xWAGwEktc9wdfa4v27hchaEngKr/hHFN2RLM5U
oXoH4nXGUWON5sw6vJhl+j4Q9wcf75uI/+GvjKG3CooIJ6KAlzhdoCAmPY9C
Bn73531fYNsoGi1/VZRB2MZl2sLAMNYeeopo2DDq7Zut5soihSH9Vo3jX1ju
5PJFPVsd6s/RJLpn3gHld4zmVPaXBecQA6vCERwaV3xpPqI+r3EmG8G8dctc
6bjeAb1Td3E9EueZPXkN2h71qavxQnfnzDBetzX9yguNVS3SDT9iqeAeTgqa
q/q2BMidz5hGYcRrGaTuXMFQLxw4r/nOBmWWWlpNAAcq4Yj60qYePMZEdYSv
WeRJi66PTuToOiuAaUlu88YDPmdSUmnO9dCX44ZmXzHy5qaL3Hrb6vupMwzh
wRnoeMe2nhdRswgg3DiwsffQD7XZ86oSP4tYaC5E/M+9pnwALPXCUhKgkf8U
QyaeG8aDKDnnkJpNnv5etWTLczpJJXfa1EqnYo7AoxK9jDNQDpF+jQUywerV
NUaeCvRIzrslLh5h15wkrlsfRC0HhpQw15+6o1aH0UT9J4TUriJEA/tYh0GJ
t8R1Wh8OEJaIiBmma9YNN0EFReirj2RYJxT24zl8vDxWXJr1GbkVCiUXwxf6
TXMbTiQ/d1SA6G08uaUQ0RxnHkk9iyv3GCp8hc+9vULErrLR6/5DSmtVuJOp
xVlggn/8ah+vRrHS5dBJgPel9mbudIloa1elgfbRZAGZ53YeLva+8bgY82Zm
IdJCJ51sW8Zpu8s3bqC98Ho95VL0Cqy4Qqc4AbZRwM0zkoxoepgtki3nDmAI
LUN+xjWHzs6VdGVvGYAPK8McFumdeziQlQ0rL9U0d4glFP/bj4/NzSF+McJI
7GlhGAuR5oQLjznVTvEPP6SyHMcKhpgRYO7onkwm9Tb1lBvqohpbugkyW4qZ
uZiJuLgrUmr5745rl1ysTJqZORdeeE/jL6Zf3ZJ9nyAJgCn8kzGFav6BCrLJ
7rVfb/g4vsyjRf901g0EmfFCTLp2XW8mznQOjVFhc4DdaObM/nhhuJwDetP4
c4shLuGeOzzu/tE8PxapGcRVct9RS51jmEp+rT9Gt5oidJxUgn9FM2nFp8gR
Nhq6PotvouLg+8XVqkCFhl0p2ct1gDCbxJfGKVZKcFMdXSmYb88ox9CW+1mw
YMfCu/+t9v4fFH7ao7eY05GPYOQTwIZvMQcfrQMABobtQHyUHr+eMUEaFrr4
AOrFo2nKoX8mMBExBCiCbSZyoYwb3yRF2Xtow7aifdqs58D2YguTrN7SAtHT
U40Pu3hVBoj8mxGOgFqpeCcUikvyjtI0TeUNRRWGL6/fb60H0v732zABOvRo
EU0MPoAIH4VrrX6o12yz082D/leknYcLcEQh6vP+3JgnDRfO70a9+RzivkX/
3VIg1aqo2oeJO50Uysyl3qXQRpnD+Rh0RhTKTfKLsd7ZzUeHnc1yN6Iddl0A
Yo8jpFznNSz4iJnLlzCaJBZRZ1fLjt86H0jcp2WRAXpfYykchFXzfn+itTwm
NeTMP4BGB78fpLjmN+/oTQ0bfXgINcgr29QGNU31pxDE4SRFQ1ctD/+EQKtI
8RvM3aaYIiK2/H7egXFG/1GnPkGatChHIwbfQPiGID0cq9/sP9913MUMGtfw
ahcBG/2MHyjHvlBuWjG3h2IzNtLcylP608EVDVUNMnPPe0Z2R2r86DViIP04
kpyUhMITeEqjBfHlpu1L7N06YrYYEA4mydY02PZ2/NYLDWUGiXTStHwcSV+s
onGcVTOQs7J6yXKWqPk/kaEvDnHDq+2HxyFSMVn75Dp+nrYrosfMorIwhYun
GbXZfFVOnfNjK/PGtQ94s9XgqvFaXVMzAyiA6JZeRv4rvfUISeoGnE32MzsY
FaVi6CUCBbeK447B/BsWVZXBoIHkmmHcx8lFEOY367t9Sdmj3XpWeM/bb4z2
55gG0pn1dI7gwuarHr5UoEjTGIl/PWp1C9t1Zf/XTAcL7SclIM4EFhFGRqfv
rVsA59TXvXQ+LIKg1Phdvs0cSdNsvhwwfzfgVy8LNCVak/S/PuxmVgELa0EB
pBIJVrxfX30vC60JDTVCgy/Xq4Bd/g4P8iMOsWSXS0LAiTocqMLBg880inUj
q+jU8eg/T+/ReRTZwyO6UAw8ruAlcKdCUrRyQQN/lY90UJwlU2+6IQcGsUMe
Jp/BjlB5dvR8eDvcmLA8crurEegvc3DR0SbrC4syhjbhLCMCVbfNUA76qChf
Buul6ZfdJ1rawMJUwGZGw3+KFrgRnTK9T3SeFQKVZ4lCs4KADxWQEBxnPFkY
0+ENr1eD1LtxeBGYM48aDAoBYx0k5EHw4jN115K0uvtCx/haR3UnhXeuAYzV
9CpowXJUdEFBDW/PBt0to9KHQ1oorsCNZsd2I3S5chxrq3aANf8bWwhBDdL+
gf+Hjl5uQoNFFuO5Hz+sZi6zmThdwKzFnxPhccvsnHQ45eTV1vKmO5FkadRc
hek77If/k30Y0pTsooEUk+7/Ol2cH2OgzTL4kyD88SMBzMfIwZozRxrLu1Lo
vnT99WhjLZLubW2G+O7GpCSZOZxkdZgRB+UCZyxyTWXH+uz2oXFUV6p+plUy
PU6QTUMCBm2u4RiMj7dqbaymKNsw/HXqExRtP5iFTleiliVgCcIzjEeqS/s+
NOhW+U9PKzo42VRnXwMusVTYVdDB2pWzlQityN4NrVrWptQb2LiAgH2hLRhK
5bnTukjhDj16X+STTKVagXBBznyIwY+x6z5jQZ0uvXm0gDkrOcy/At1Nhsma
9lvHLsKyd40S5OjWtZ6F+Z51abImjE5efc+sWgLhk+hFiYWUAdpDAsxLTtex
wKZG9+KRBFRaU3HbSElNkeq6Y4w+xNYxcrM4EUK/8wmPgor3T9AdkVa3DcVX
9RaSW06CMz/nQY61CJdd9C2iqXhH268KWv26EhOGF9XC3b1lKVsaajKBCYz0
bOGBB/A8C/tTj7bGCsHLUTzyF+wQfAYiIb7j4Ip3h9MMuGEBw7B5Qb3dqu1V
056JXbEiTk75Mj939rqKAXVE35zcVbFlYHCk7SaPdAMRlB0hqC+WNfpu2J0k
9zSYSBUT+kEK8By7nY6wFdoj+xt8iivv1rqunaDZhA5IPV2eaktVwaRuzmfT
hayYL1OfCpek5sb7lwiqSH/K9ZbTeFo5o5CuYqfkvUb5f6pgCPYkOexeF1KN
+t7xxdISSJymtalMIRmEJP8NXZTZaMX2gfGkMZdStVRz7hr6sIR4D8XDcFUS
EtOCNxzsgnRJS9UgHtkh82hJvbe6WCU+X8qTuh+YaTOTcXtzue8gFCiw5/1C
Ur7uxQVnmNRsGDcO+bgGXJvU9PHLU/84KsLtBgfs+hLKPhluJ2w2kt6rQdQh
8z/753YRUwlTqeqIcsVSgl3UTjccq2SRIxJZSV9UVXeBNq6CcEaJFHSlYEO4
KIuKupf5RXOsd6DZjIO9ZJTMHOQQZQZqMH6xrsySrtpoBZCKQLnl343ZWiJ/
zuzU6i0ZH2eYrAP6mhV028bne9zbiovTynQ8Cvh0B6uLigSWaPCSuVJXa8eF
3u8eXrpcAvKN4XElfIz89XUyzYFgiqkuDQFTj94WGr0Oh3/nj7m46ztqCY3r
90bMlHF3otlBjIYnfJjOJWhJuH+kivWkW0vfXyzUEv8v3gvtz4GVGRGiYi9h
y4EKfDmlPohAEktr7Dhz1IxW1TIkEsqjyFjU6IGBkKWRrJGhg9Te8IY9GG3g
DQVtcVheM3sC6/QrsHZ9xisgAugMjZkCKDiHAXo6dLqk+I0gYjpzkCcU5Rpp
yUt3II/mcXnzUPoDhVYx06LENAlWFaHODWLYDQLWWR4KvLRqhQssl16aPB0N
S32AgRTV08+SmTZr+T2Fycm6yv+H8XKxsyls/ZLzdCeuM4oMHm6suTt1lF/Q
5GDrKuhxzhtHf5BjChCTaAACYPaog1ktg+iUWknhhrKHbDLmMHTBWw6XvfHK
qBxN48sEJFMQbD/eXZjK0brTM3cTtuWLfMpPM8GDEZeCyrEscUvGblrnA2oO
z6Az4uCtah27J2yR0AAmRRKTWzSWisIYnW3SdkFU/q4bMEQMLnqJBjPWmwtG
Y4v2gO2WWAYCL8xORl4GJDpBIcxyfz6NKcl0OtTuLwdQc6idVy2N/QD7Pqm1
Nltamh+fcrxJdtOBRhhv2TXFlM/srF1NfIHqZHi4jJLMPpob5J2zkme2zZJS
0Ja6TN2l4RY4Rd+AZ5d0UxdnAbbfvtcMogW6LEe+/Z5VhnaQhgMBUqFao7u+
CqIGhsyUJi+QtmpMrIEPca2bWAnvBThupMudSNNHfAGRhejcHzjS495bIDpP
sdkMYrAOK/vluT9V35lnkxy6UUbBuBKNH+0E2JxDUnj9lIw+tepOFZ/HNhCO
JW8QixkoP/eCGNsAi/i4oT/SNLrq4L26AdNGt2g8UsjBEvZpVt9jYbjIxVDr
FWJdcjBcXY+Q4kRasJ9e/dsajrbBvyWb2MiewyreGqRgF+vZMlJB5X+lG6nL
NBj1yuNUkGUlG4Dn4mbCzeb3BBRnqgoDFoP2ygA2iZehcUGG6DicFBtGwzd3
+mIjTArcb85o83bTCAaJPYQcEXLDRqPG6WHfPzJnFjM7rx9Gf3/nVFNmxA1z
7emLT12mEjgEapj2k+A5tMcfN1o9KZ76dalRyqpBeiyrQGhISROKLjXk0QLo
Uzb9Z/AHdRJ0YqJU1GwRfnGR1/yjrQdpzYeO5AxrpmeW8Gms4OSUdbvk0vy3
adcrsLVVMO23kLhtBH4j/dkg/qow57+A/XBy54Urcgbp49YKRzzi3mY2GltE
mVTcg8a5g5NIBH5AH9Irzo2t7zCGOGjeRe9nE9yfw0RcjJfSHhsebMbnWDsh
LUQWh/3+Jc9ChTIsVkB13GNILVTIGAnpOHfGdJyj8k38gcWDf5drk7sUI5Ji
RZHMd/ziAVnmnyJiUG8DbtpCaAacEynniN9SfURL0AYJEpJZ671/BK3EbjLD
nqwnvRozq9nUOZIHXiOg1Z9imm04OPG1k4K4Ty9L6WcZ9xvBrwGgxjuV2seR
5S5XaiTu1kYMgnFdfA0x4uLVNV6yZ/M3r/ETGPViZgxJZi/DMCNVJtv7MboY
pfjGXLF5ZKDzL+KF3tJhTG9Hb+3idjfQLoCTmI63oeaxj+y/Z84wwhPuTJ2v
OK2ENHTVDVwPepe72dJl00Ps4KHc1fXiT0Ur3PvbGF0COAGp3RPlQSzixTb9
7kXsQr8CJ1AKERA1CvtWBOFwefLlNLmpAlF74y/8MSAZEwTiVEVbMy+IvcuA
haqVSPMRQekpG4TnCmCFs70u25GliL+ooTWeEfzSCyk+9GXfec0dZMq5w4IP
SIABxZo9ymIJ+osDq3QCd9qyIZEnituB69JXDmALUBMfgra9tN7ej3jdTeqp
fijrBs3X+vP6z2Y8O3WIKfAHuMl/qcsOyVLicHtbUd5+aEDc8Ox+5dKH8qsT
+mHJI2J03TQo8/kq/RqxvyzRSC7ljHJDemTCoQqpHcF/XxV/bDPUuXL/YzSo
hKxESWjjBj5diiIp1fkzEzSU5yH8T4yADIuK8DFXyOl6PT8AnXLnXHC2Yn4X
OuEsaEZZAXyGsAmm1zlAl3y/rG07egYL7UqhwSqbvfyJNv7VJ736FJlkQpja
dEIAVZpm5I10sYQRAssK931mYoRtRhA29E8AdG0ORboJJ4m9aNmxt1t8KcJ3
goGfz85Bv1U0ICLbg49bJTmi+KCRwn9+M3+bcAgb4FAv9Odp35RYLXPXOJPg
Gbe8JV0wMTkbWHBRVN0Zj7CeRe6IHR6NBPKCAZr2XXVw+yw0CEdqlf27o2SE
WTbxUmT3+SYhv6TcJ3YLBmH3sBkUJjHhnYalHdMTeIgzeq40GMvkZjCZj6pB
88w6g0RZJuwbxV1BAUgxkhJpeX/1A03/J6LiNwVItt1ovyrtoKJ7LQY8CNYE
sJUdMo5BaDcecZ969V80ANVyjtJSec0fWlc/eL31a1Zc0DhpCA7Y16DiBpeh
7W4XLAV4oZMMQjjrkak5+GCsqXrlY0tT01SItbv3DxwgJIRu3rmjfocKn/r/
wYKZuWJV9Xlww3lwA+UNca2O6JjP4sXNdwrgnm2Ya/ioAc6+n3qNQWpo4V1C
5B9DccyBVn+bng6cmhqq4PzMQmFyD0+0/pa12h7/veCOmAfLHaUo1DUNJMfK
JgJzMvWr5LFXXYg5lFIy+9J+q/01iQE3cPr0WCe629Yau+yx0dbukhw2OiuC
8Jnqw5oo7BI3rsrenQC/55DoZDk4zPFAsiuUaBv6SQzPEikhfHTXgw6CgYQb
mK9ZVaYAXUEyZnZRQZqRVtFgYDfkXQqincYwchsWUNb1DQpYskeO0w9+BaoC
Ss051wpkNjYcWe+y/Wi8XBg9l51k2EEp8OpayGvIepl6xrxSr/6aNPJtSDYT
1py1+0DXqElPCq7atRsslxo2HAuetsczJ7OXVtzgw7bxVE3SGX0tN2i9yJh+
bESQiVbI8w2ewAebQF8+Z0W81GRekjwpqxxnmRy6YmkCL5SWJnDiOOtVORRp
xgVcGEzQzalDhufpYnAX67ga9hfeBvRh1F+PwKQ8AjT09cSGMPXAhyefNrdq
aHrA/vTNN4bS+/PcgPrhUSX8P5bP0MSRmX/BBs1tejtNDwOh6b7DF/Po/LQX
73WIcFqiGQa7DSpIcpoQh1Fp5QsQlDlV8LhjhnxvabE1RDDCuuDhHV5zdZhi
2NYAzqlPsB+J1eB1hZ1CNrtHFzvaL2hllwJgvoDt9e6mG8PMFb2BFxbgQhHG
e8c/xtzR+0i8qg15fSGcQsp/W2kGyjtpezxGFYwRR161a+ZUwphMSJvjAKu8
bvQJUSgY3+Umr9i94/pAmtlpTsK+EZjMwJiiitit8ly7gvwednXpXQbGQqR8
73+wnRFmzxlB/t0SsUL4hoJMalCatSgNy0rCHNxjNV4PpC9vVP4ygMhbMosd
BKAZmYlA4zHC1TBZLom/kF1CryfspswoLekYiJrhYDIYrFF4XRQ4YJa0a+5z
5hi6OHeAvJ9WHzISE+i32rkMn2ifKsPKdzMVFfLwLcF0Ubvdod2av+W7qyju
DOe6I6cnmQHhcK4koVmASA02GGyQG4JKiJiTopMZH1YvUpLDNv+JOee+lGhd
5J8a4A0cTUfRiWHNeMBxfqWwtU1hsH2iUhOJE0ya9RZUhwqlt/0i5Oad5ilB
mKgB2NdaAKcYPd+0aYt5Il7WMs2iKAqdNCBItMRwTlIYA70208ZvpzZ+GrOP
QLP+78OYErtXAgUzoh5NvD18zs+N+ix5asxZ764oUSRzwScRTL5qQtUaLbOK
hu//xZ3WzeDPL1fAxlZddaa181f9Y8BQ7jUQ5NF2L0Oy99uRZNd8CSiYFUWG
FiaXHXJjkkx99Mza0avF8odOexaTm7JxfXQRg24vSXNhpzo9iq+CqRgQAiE/
/3nIIF31dBuNQEJWDri8IpDPmbWnZTz6gcjRrwGl1MaJwTy/en5vjdTyhL27
iXtIjZd0oCPQx46uvq29ASCPl1sKamEDwlSBmU1pXl0lNn5FyQoB6eHPtZEv
1+9gI28nDeoBGi/rzgbxnHHAsNwlwRIDzgcW1N38uLb6dOZS2conHiQaHeU7
BYwB6fcWiy5VqwlMLWW+mN4try9V3F2PTc6PszgEraqcpopWnr2x7Q2oFqS9
+HtAOrdw5g28nbdiOK+N5vbzQole4a5SsYjEs5APLWGBJTqmh6n1EPLRnSha
WIl5GS+aluvrqVNcTf6YdR2io/+6k95m7aByedS0EgR7eJwcJYQmkoBDMxEv
jcU50Mud6CbF6qrVgEwHnzXY6Bhnm3xBr/1V4mJg53vV+YsLLa9TLMs4Q7/l
aiUOOwibxgDusHx8DxbULuQkP8ZRGRnGycy/Q3yx0LY+2IDRlgJ336bWb9gK
u5KRE9qchVihttFOavzvYMB043F19TG0n9RC5scmb6JUQvCale8iaHpyEQzj
aEVLNcIaojWEBv481/caWkTsC1i75uP2C8LNcJQ+fqtPut4mxRSvt+ytZFsS
2MRD5mNQK3kYtQaY7ZRvBBzVqnQW3+9Sx8iMhKUydB20N0rE32szE8N048po
OHi8BHCgMS27mxzbeGK7ekoQC3/TKwJhsFgVOJiKNdR4VFwi4YP+PmmFV07i
HpnijtLDUmoMDSQn87i1JOsS7dXF3oRDzwE21pbrO8ne5YT5RKKelIv1mGoS
9GaFCe+Y48nfiW/cIqQx8MUOUjxVhlS6NyQV6nZGH1xYnTjvGlSMkjenamNj
GAv+tl6oI+pNHE8tetqwGBJYYBHFuWm4pbvyE0d37IKev759L5pIlCl0p5D6
FNd/YfwlD7eUKhd7VKbL4UgXZxNL4lalMG2qSqLXhHSUmVjcuHS4f2e+1a09
a+HlGmNiQEHMQqcqTYcJxdqcGC7/WAqflg3OcpDrRt0I1oSfSYg1O1xcjZkj
TVi+cNGVMTvQ/N8e4QGRlA7o9G+nAc7C9UcS4AVQLRll+cpJA7e3RHJUjS1q
BeBDsLJ3b+u0eqIIHjTddHl/i2WioKyrseNahtfSc9PCGBVsiistdxVT5INC
fr/FuVjdBaqEMv1halPSfHaWttAUjARR43FStOxAaQjx2O9xMZawQA7mwNJK
aufO4+ZC40Lp8J5XXGLrZFmHeI2gVJi3+UP+ZT4HvsQMS3R4biIiEEsfzRnA
jkDM395TtZeOugHJJebYXWZgDviMXn5kxSKOhyb3TkppozVMftj46m88nZtK
d7DunYWxDdAqpzrToUJCWBScfS1SmKx7HSuRx/phlTpn+hdZB0Nb289Vs3Mb
mEPIly8ARbxawxvDCGb0mxYzokEw8eeR+5NtmWEBLJDvi5hcfV3ZxT9YLCyr
xhNkIf3YYs7sk/RloqosSpPyuEUWF4wtiBN/Uj0SAcW9792w0QL3MLgU/ZcS
LN20bbruihA6Jh5SDcfZ4Td0C1+yc9fAgsqy4LarKsbByBzDiXBb4nQu3Pir
jvYle3wH17rgwyzeUy2/TTrghY40B7A0PNP8rGjaQNyBLUv1OtV+HHTCl3Mz
GuNlQDswdji1ASWC2nlAaDnNM+Ma0Z+ZOZmqI3s2q79bkmVwaM+RCf32kVYM
3ZOCFtZkPDCMW6jACd4kXhM1Jq8gN+DYfmVPFKIT4IciFhxmGNEp0+SPbc1N
ThDR16bC5tYDe93/enn/GiV4x7eSC2pTdxZIYBsawQRn64KYC7EGd6YoM+K0
kYJ/x86abIW5iRvX9Iyq5gfO7HgYrc9k0J6ecQriUWg9iFPnXdHvJL0pp/pw
XP1vgzaPD1gFjx6VNbDWBQYvXWIgkze8r6UQxL5fzRM57kgZSQoz8yfs/PKx
jwfiU9yLx/NZ/ZgDtPkR8qoRfDijuKf2VjbfpZFb7kSypqQhtzO51vI+VSia
5dygdKE5sFP/5qHo508M/K268Ns86BKi+LNiscz3VvMFLyz6/ibv2avHYxze
yk5NVObpc7Uq95EflgXe6jiLSxZW/I+NBKlIaipKnyKEZkrjyIcpN72oLDrX
EPfesqUJDP6yP2T09H+Ui+c7M9P2H4NK9c+IgxvsExZtJJ56zoJ4Oz/ecRzK
2pMzk2gYPE+MTYfmdXwe9zTqLwM5TUcnzTby5WPXGipbbsJmmXn2qfj1h91R
vIJdPVVN6Kx6oOeK8UoA4Hw15yb4qA5S+bH7r6EveRU1eMtUu0m1uQOkJRWC
Je9ZRuLjjp7HJsM3U2ZwtMxrgT7gXKDrMB28zrA675rH/gn5MTA0II9nv0jG
ix0qgUfbIARK8Ga5bD7hbzXunZcUTZLEb8y/KqJiQ/dKYMc7jcKqwS1yK3dE
IfmdYhCGEAD7mPe4t4y4T4IR5xCBRqdpGDASR38UKw5AQlN21oqfWt7bZ7gL
PUmnoB9LneL1GzU1LltsPs9GBF41z8f9GtSeWKT0Mpgbse8eUQWcGJCMGm7X
3UKqPRCuUxbuoPOjuvr5qmil77/ry5rbUeMfreusuO4Rs4FGG/tCowInRb3o
4qUbeXQ4T0lCOvSEKH9H9Ec+N/yiH88RjlZ5mtqe4985gEBG+ko5Z8wSd8Hh
5wZlG7D9quXtsY0bo3OECqV/D6f8O02KdlRVKItl61yo52tpSczq1PsDPPUK
zqTJjIYLkdvHWGLiF5up2qTYJ+Ke2uV5xnCtE8xwuM3aeKQUyMz6vxIo8oY6
KDbF1Svd4XpsdLIHnxRmp0IluS0vFFvQRF5rjPOVB+svAw43o9JTCL5LkwE5
Eup8DsinFGUCngViGYRlnAzVtzBic2lwuC4ZmastPE22u3PWIusePrLVe2eD
JD4Kw/eZq6Kx3Yg7CG4SrjDmDFg+pxFHiZSxrzTBhbwlNTazwuy7XQX6Ah41
mMNYJSFO3ww0nPbJ0shyQmy0oRlxI8mTtjN8MEl9KPreK0qdpTWt157DoIxZ
uQ3FkNE5mUxNEZv5nvRuVfnj2pCErmHrCHfIVNRMLeGGSNwib8pQgh5XnV56
plon8bGrweQJNf5j3N41Dpncl7mBshT0JPCBhGj3ElsGzvy3BI99oBBvW+Z1
IWCL6cpNJ4dvCK4GUB+QwpwBgPFh8NAoQlLM113oFPkk5r1kK4xysauv1vNQ
MTqlgfdCFfJbrFYCXqcyH7/Q+K5gd0oRC4qxIT+kaUfvCsvFkUPGReIj0hTG
jc2Av2tIdVbQr2NhYvPzUWaaxj1EH2MNFtk52mR6+gPDPI5taxuO3eXmqzhg
ARy7boSYTIOPn9e0+LXmEs48A9mTxemiG/iXYcKL7MfTbiqe6lLfkyTkIi44
zxr8ckxIJxUIFF0xp9rEuj+OMiPI9GSaY/fMvtNJJgqkeq95MUhUzst9vVSP
udS6qHKh9rk4rVcVa4szqqKXzt086BoFQcApOq9kKKnyinjiNIDN64qukK9g
lebId/zFRQ9GBTJ75R4RbRuagPyUcVUiX+hdQkpxnGSd5sJ23fqL4RRGXi9D
UmEdfD/S/AyU2wOe3pqWJ1/L6uU5u9a/sJSMAf/AhmMeTy/bPc3cZAbg+bDJ
DGlePfsEw2xZwbm0Zy0g76of1hI1mXT3EXwQCY43kk4e1lsTTLCmftzT7+59
ruReTPzUsZxOMSJ8SLn4gdAr7VuaicyrpawYgF4sqqH1+c1VQThd1Jp529uA
oDXLYVQXVaoPrubioLVCHDVC6nLSdRBfP/S215KNlaEqmu46qo+XKJJ+izxX
AUGMmsqQJzrV4/OUco3nqfPZxdoGNc8QB9YsbFBsRrxmcoSd+vDDvb0F3M68
ghBYkyP+6bAx9AylQR0ZX9h9FdKAbdfc3iLLKxmyZYueomsjFdAWHDM3acyH
zVi6x4DnLRiqYPIPppNGj/STsxb6QmsAAcYX8btpg1U1pR2uQ/G/+Pwvj3vn
ABTtMkaaFH+lNcyM5GKrpgM7D42LldIMUs7VI0Zju9ilfL1pE5te32dN66ti
oPAG71rcgxm8k4mQrI4zASPBUMCJtF8FGbagDOoe8bp571Ps1AcU4aquNfVh
IczXJKgRJxNNppKPTa83iqF06rh296USedwoZCsrYUI6CuxRQrN/n+7dYFhk
5IoH6mtL4AnjZNOzB+0dZHF3DQJ4i38heibdD2c3AKt6PMRvlLVicfhKUtGg
j1Iu5AuLYaklMGgO/hYheSMqNPp62uQV+pCZcYvO68xlEcuXzOoocXm3BuQ7
c7Fum4dfjfZwqudsrHpxpFT0kxASon2OvMef0Y4etwPE0oat1/bIWnWGKmQi
OiXGd5heMqMz/BcsF82I2rAPhhm7p3bb/wsGF3DCScECHcLZaHshzQ8gvrCd
s+zurxyNe/8M4KKUuWJkSD893CIXwNIUXrcEwaVcl5QLZ1PkjANRhbzijW4K
yUw0pCDjN2wa1aeFFALXVfPB6j1I8AWOA0U/nUkJesIGbHG7krMebrsGHuwy
n4/E/gs6x6XXxTSpXNj91suWCccUuXgT65rDUQd8qK4eh28bOOsjhKesMHfE
Ady0X4kzM/6CvHWriqGcXzopIbpcNsCwyjeII5efKj/5YWhAA6eRVK/DlNov
51sCoMaX8iC5i1kyu2hxlFqH/el/pyt7iU6R5xz4CtWI0gmdA9P//b9HEScp
nHunzf3wF2GqHYKq+fQQ7YJxYzRgD05I9wE8S4yfhSPLda59/BzF4vwZ/RFt
RIfUyqABIAlgtM13SIngMduedk5tRygoaqoskbPmkKKFvs2kwReLLaVl8H1Y
hkF4WDWM3jWcf9uWdHRwD+y+FGlZJQMHqAoWMuXI+vVgu4OrMNj7o8VfvZ8D
zqYCfBiOlQgV6xZNKPbJrwxzuekFkrQ7ZePvp+s4sIIG0flUVUmr99G3vdTp
x/Xf4AEejfCdlL/qiHj6iQFBsgQmhc4xttjxQk8yqFv14HQiWncPMlrTwgQq
8uzIKgac0wQWjZFdOFoK7zprYtNi/mXx0NxZXADMK50tpJf3XWmYBnl5v9A3
fmZvN01l3ISeLC1S5an9rTNIQ/xwZRyG+XQZHjc6n0kNgp1ZYx7qnqPSGz0b
v0InD2CFTqgfk+xiI+VdyyoJop9O1GKXKHTi7b/bdsVY1Iq+DCq+3ig2eQvn
YC13d0vRTQOCjigW9yqFrQQf+e4s5whrCztOFHwtjTKqM7em8+kaHWPwywjf
MEXCqcKkh9PnngHPbDAiu1WkPlRiy5GyVsIxfLX9a8qroueFAqL8Wq2mEEaF
oUTVdoT3ybFdxoYSM+6kElksMKMQldSZYyEn/C876uQRCcc76aOhcL0MVnF4
4PBaYbz3ziEz/4SIPB8t9QVLlFjraEEM0OrHDNzqkfqBaxQHl7bv0Vf5mqRM
locRCt+8tf4DnsveZ+PukMSQtHdYu6+XEzuRuNIbFlCpqlk3EgNm6PJT9eUO
g+bfMnJbMC1Ob7NYi3HINPwoQIU936elh+eFnjvN+IGD7D6VtMhHUFLnxM1U
WlHuRJCbuAAtnZ4W+LMjeTaVfg2A+YJBxnK6vz65QmMkPW1Qkyn9NzB+sOr8
/lbU8YXL8mgcs59XvWRq/vkPegYeGI5+Z3JzV4gF3orUnzz5L4tDcDIuycV9
d3FOz+zm24iSL+IUtsm9+R/sjKhPqswQM7RF8VEYth/RyacZi2iWnGR9gddG
VYax0yQFQXeQzn0iXOoY2BM1Fh//6PO577JId2M9Jtv4FM/Tk/+qIByQzVfY
IZJBInZpmLAgi1nYg14y84HDdsAqznTORGhPqcbNIULNnjC+jyvuwVQcu8v+
oQNpPrH1h+PzWaMbCueXHx8yb2zCBN9sIHchww82b2G/9x172ULvsFf8vimT
9xcazGdv9kDbJxbDMsIxinlE4YYFvXYyoQytFjxE93gMNaOxF9bfXK7+vEwJ
hyYeDPm6zgHD7/R/UtUIquKtiSbKWFL1yg0rDsecTBfbTz9tYXRd9nBN+zg/
ddNrIWXXBN3MbbqrY8y27LGvIpI+2gNbpyabqc/AB4inol1V9leVXJUf4iqV
cAesefL4Cgh6DG2sx41nJXX/NMGOpUqu9h9SRd+cGOEROERjZmMD0VGRJT2Q
STD/nqm3ftWOi5kXTZoPK9HTpl+cwzCax9jhLdFQaUcg+RNkTTjI0t1d9p/p
lQlAJ7qvmqkg0Vnc2uoRVndjn1fXvQOC3E2xJlIefRNRPlCfG3N74EUW74YH
AB8w9FeMWfUisK1VQWHfMs8XqrQZlIQs9oYpUl8yE6cUc7fQXC9hYqjV9fhw
kWWIcL/dUpWs+GtU/HSUdu+gcT91F1t2hXT4I05s98oFpEPMppSb8li38ecv
kQoA6+ycIjfdQoKGeDLT/CV5MPW5svc+QKZtNnRiovG1eR1a4uLcxII5O3Dy
VsfqjlGjnPWqgcVvWqFP04r1bV65iVLJHup11rtAdBQ9SI9AbDrFzcOpnCZ0
yUW5LshWYZARpZJYDFgyrbTfma/n7Fdpbbz8hfTZjW5j4vCwAoP/hSb2fK/3
bKydw406moDLMoFRBlcgt4BjaCeLkpgkvvh41deASVXe8MwK4n+s8tY7Y68p
u0ebxCjZ0gafoIIB8GQF8LIEostH9sJTy+Fvzqml/jKgFkss9xafB4GJNpQ2
ZQtw+Y+9hUUfyXHgeLc64LO/exCDB+NoT6Sj3nHiUBRf+pBcra6EAYHEnj4f
hgwXF5mgeZLVSLmBBOTkO10Toy/ni0MnVXmtWVLcUV0xBnyBApWGQ/kjXFuU
xnL/dPltZDM5VH9g5UN0QxUcptovJrqYnVWqL4YmfJU2ijbHkTh7wzG3lGFO
YgHYTCzx1zJyrPr9xb53X2w5w2EVCgayhMCk7djNlJX7f6yuSxSzVQz34es+
pR5GPv7ycTQwoOc/BTSBXe6rwvj9tJKRPL40nJfBpvUVGQIwOb1uqJQ1jq5J
A4c5kwsoiZ6k8fW9YJdccoBH8rX4rqytk8KDrB4lp5cNfgcMG26xIj31t22p
wKVEGbR8BjHqDkdaWtRb1aTSk7hHPC2NtU+MYg5IKEOtCLsyb0yKd+LvGtsz
CAttRi4NYJDnFBLKHVTIfByc/nhV6Iq14ooSAtPIj22G6L/CtUk7AEX3qr/e
BQA/scLinn18asCdGqfsKdkoKcLt0sC1waMIGihPnnEny/vPLGPqvunN5oEz
4ERo8safFwylbw3bzOJijQVE1AytTeLkJlV2QGIy2CYZKW0s6USV2zF5FgtX
6aAUBMjTEDSSQ1gpFfedhcR3F3Qr0hUBEvg4HbgkyKWyAcx4x9u27KoAsj6V
Hn80b5SFWQMlyMOgmxXw2YWfQMVcNf4Pwx4bF6/k1vO+EyeHOWDzRrUehCM0
n7SiAUkATcqRzvsEonIEIqcoemimtA9M0KXVriSecAL7c5a2adh6Yo8w7Nbc
mSD7yb/ZmB2jVCjada9NFJ1uk0QpldLYc//AYtFWAuZr7CTw4/u8kds9TDmx
gJocycqjRfJx/ltf9S+AN72xF6qsZ3YHzlITeqAoLPMtYdukfyTn0Puy4MPK
3M9Q7eCzRfAoIahNPNMw/u0NGw+0uFCt6EHMnHfIUULUCh6dc+dxJd7wtUDh
FR/Dxuag6s0ju5Aa8McEWLVnBpNwslS+gEH3sUkBBDrZTn0FJQASLXBcd9ZN
/A6KLBeomyHPkqVqkX9lV6dDfvv11JS9OxVRpou/WhYJGo3ipah+mRc2hGac
KxWXHxwHZegBqLynQIyuKef60ykgXcal9TkuEQZll2WmMT/rFqr7IIRzUZdD
6+QOUS/IknaUkagSOxyrrwoktrCtLi1tprQDRohEr+3y/kbgdptR1ln3ln3m
+gQcR9cAEUIRt6oz2roLqDxJ3Rp27I6CypUdR/tSUomkJwFm9InaSQXZH3WO
4YwcMKAklUQOvcSQNELgIsV+eSS6wAcFYf1DfYUBn56JB9QbA7EnUUTuqFeL
wKsl+H40TITdB52iNzQ6LzhM0/hfPiW27zJpdKnREPLODzULuElXwoUHqHcD
dtkzcfiSL3stapNb3RL6iPQqyo9/R7r/aMcqmfTSL3hL8s2s6/9f0rEVhHwc
hqSEaDl/ESouxPRGnWqaYE3tUt7Qtf4PLYZij1Ze48bstjCP2A8awwZTZZa+
5TaysWT8O+gaJvrMMhxd44okZN5yDcH0N5c4LcEM494TCHsTTNibiMxmuRjB
dlotmlTOAW7ZycrVWv9c8p5Nh6LbnHCuHVuP4ZluoxOvP6zDYTUaJQejCk6W
XhcMaAF8jPwXHuO4gHjzgY6d+pr/3rhUr9+BJ+rj9Uu/FgI8lkmmbJZ5MwTF
Ci598rUYfMbUGxj70+OcZy5QnlJkmi95Dd+TCnY9UnqnPG6IgCbJiWhKUlNr
qGQcDtshzrPHSuPv439MGmYX4jNULxg379jsC3er9fkOPhYUZFSM+luRhJi3
lgWfJNYGgJEaHtyLv+kEH6Vd60JtQWGGFoeqzorje7Fx8NSSVNHnB5FdTwwm
bpIOGkBwHMFDTuDyGcPJSm6jjAytkTeRYf2DfE1olVZ+txF6xdf9FH4c9Sfo
qqXgn8sWhrRdMk0OodWQWbTc1rWXKxNsjyPKNqn9pHMgsNV2BPHXX4Xm6f4R
gFF0T8dMMTMlsnoarh9d4Jw1JqPpke2Y1HE7kSj+Vh0QuoZrzKq0rTH3XLaS
7B7elXofBSfrhM3qPrVxkt6KrFAM99oIm07+D8veprEyTCxnl1BqlpDKZetX
4NJdjG2+SnqIoXh6Eeyum1IQbJPIbvCzBFy0mywVzpmvYX+ehXc04q4WHmIu
K21IGCeybHh8X6UbfHoStG2yE7Vph2pQpyIh/aFw3NNPhxZ4rhx86NmM2keW
6AkynrLdytSjMsSblC/O3Z40bmteyd/7esRc9zNk8N2gr+hWUqkAolh57xPr
84K/Jypror6PahcDflcOg6UV+IAP3YGSO5ec2N6RrgjKbP8u+SSYxqAnn8LL
/Sz/TDR4lJnWxzlHvsyRmH6V+egCwzbZ4X25M8kEboDgJPg9cDndrx9tW7Gs
qdi1QUC0Ef8yaye3DIW1JmWCdgNqkkkLPBC1rNGBtYIhW6Bx9IvHE/+ORCLP
O1vEb+Gcc+Wzd7TFg8TU3p0QnkDxeOepC4kClLA2eu5tFYAbVpDM+hUhwa7i
q6rp8Pwd11LGTka7BUdTcLW1Wiitr3/dpX0veKEXBHmFgHOtkuvMlP/mwQNf
pPF9KJj2whUzlwkM7ej8lBPhEl356g6KltAlhaw+IiI9D5xBT22rusDDpc9B
6sW4U4jZlkv3t+mSasjb3Mp/13sFWjperbK/NN5CTuNgA6T7pEKQ/nEChnWf
4dCPMnKxLIy/mfz68aSc/dXN7GqjqEu4I2WLpuHJevyc6fu5JHM+T/zqbKMZ
QBSLf6QhbJsGoRGQx2+nJXDfv+m+pLqmGeeDMzxX++3m8vN8JTjLI/2SO39c
3gDb3idqzmkIaj6qBytn99arkidSEJczZxxzziN6sCHz6N73u4bYhX6RiQdH
SeC8EnnAr8zsMp7yy0ulVY/NdnH/7qAY0W9m7BoZJRfizWTOag+dXXEHxjq3
Go+9mqCC3XmglKoiiAS/cj1nUu96DaV2MqIIyXIQQvauRCLIVddqJJihxB84
uXYUtVRo8aoOSRkoS9VHWUAaEjHcJx/DC/dKqvhAvjX9n7odN0nFIxhqtKiQ
XUfmc0eO6Jo4RvwCQnfBc4zydZh6WTMd4uPkX0KtD0ABNxf7HkvCl/2d6ue/
bpvS3OrE5NZi3RvCUkPmCA7e96a/A378KVl+NmcT/YkV4o8lxHvsdZ6KDEH9
7BMAP53RSW+tWclavkQUge6vrH93xrtRiBVDG8bJMSkmNPHZGwhtzZ3h7C37
WEHMzsJcfxA4N87lCQLUlbNrAvzI9AzZv7Cmg0PQcp6lUImynZ8vFZTWS/7A
x/lvUqzveE5txX5TIpgqP3ENh1O0uZ6KAEJFG23Olqi2aa28g7ck4WMWFXO3
UZs/cdIrcFFQj9HCbhr1vPh5ednhTTSXXPOd5K56913QvZyW7GE9YHdPiQXR
ibouVD14nQbhJRnxxc8kHFGoia8rLCLhf3JiX0IinfamKC24Op7/IEbHjs0n
n/aOHRxEP9VP1rA055k/pR/Xpsmc8TDviUPCSdqOaT5m8HWu2XDkUGTht0R3
NS0aTlE2Gfn08oV8aOvY2WKoMAmBRzwmm6AcDBinkRha1kQpmiPSo0n/mhQ2
eDkoRhcFhHbE3E/4p42bCp3xfLYdBOPCHfsaLi+ziMFzwtX0bVzdGoz8/+lj
B2HMpTBU4T5nu0/jFrdmA8pbeKrl0v2/YiobdWUhl7MFdJqgsAcBp36c1F1a
g4jyF/Aqw269yH97N5qopLPLDbc1UrJjU3rzRDh+hzKg6ZdUeo75xEhf/W70
0dhCFr13GGnS5p3P1ZUDLqcUBUBw1/U4O0QohurE/qdZFfFIuETQNGzWdEdU
JhFSNzR7zq46vk8E4wc9mW0fQsO+ayE8K+hXlbxS4uQEQBoPnMu81qVqhtUT
8GD/GSPvgVscDf3jGVGWluNES/zA7BpauESRxDRXDzNlI2M4jz5f9Kevsgp8
U8Cb0LsmiqPnxjCEE4fovIe/CoAMQLd3fpQYFJeOolFWIixaYY02gYxUAc3y
on5v+2Oew/DG4cPbtJVCaypF8i3mhjYqyP4RIlKRlMwX5m/7sAzEdtW8mZ0w
pwUFhtjXg0sebBy4R5dLE2TJhkt5lsPIaPiGJzK2UOvxtX++SzPAoPtiyiUF
P64JYVcqxitOuCNh7VVV1Us40FGW0jLS6H7AArrFTmd5yMZaJKrZcWRU/BCu
LP5FB2Qd/Sa3Fkpps6i29S7IEccaG3Ld6DqHWQ8B8ABaBEmR3HzUtklUHjQI
qW2Z99bxl9pFk7oM0zQ4o3D9m2IEFf5N5pbYO7VBg1NX6c0L9WkSLKUrKekw
HIjtORB+PNGk2mUb7/FwR76d27oTSKpkSVEZ2E79l/JYeVInzsL0h1yQg7sN
V5xcdMmJo/TJVYxlt5VhcxuO7kKktL4yrX1HPRVFQS3dDYFy4D+Uf5DHU25s
b5LseMqxaZVoc3Z8HGLU4EBjeNtjuZ3+s0EG14LE1cgdmUHoEF090JNuM7/n
YU3zetT2d71yT/1G7HVjFsu/JCPL81v+VnbO7bQ7qrzs0T9h0nEcdr9EioO5
GA0JMb/bVyE5x83yfe4LKaKbXDZmzdlAzAojwMptESijN0zT9587ygKp2h/I
wU5mjPUHSZ5HB5N3tKamMP39ixaYU699r22KUctb2hryQZNZdw/u7Wb4zkKQ
BIEr8dT712tCV4d/NI75nSZjj6pFk3C1ZBs1x01zsAVteTORUQihVMunA5Nf
R4WGSeXFNaMyOxz9PrMmapohshTVxTgEFMbpn3MofoYsDrQ3X8QhjcJTb9PD
9BZCTEWZV5lPlunzVDd0YwrUfARkYbFQf+9SdhF94CtG+I8Tsl7MW3YPPAyu
WM1Y9HMK1Nr3NBVKCsfAPIJNfGCi1ZyQjcTGK39LKNVzlMRtWWpW4oic5IbG
2wSxLeRmSOG1SdzfJhw4wIago+0pQ33XXva+n68ksFDmO//q9/BMA9m7mLbq
t1rxM3hqO0ahl/Jxf+dlukKs9zpeSgiBlrDXIH7Gr11xL/Sn/1cfBsdki0Gu
ttgEZf0ZSYtgjvj0K+azqZToC7coCUjfBvl/49vrshv+Py9630mFI+sXrqyp
YzClHWYETH16zJllMsoQAniOpy5LTzAo6SetXmWJXSImm3WrJF5CkkSSFjBl
98qOJBXQj0LhcvfxQchg+JIQR+Uue/xNblkMQpD6DiCex51HjwEHQ0X03ml6
bMKbnw8IuS1Zj/ZpF4sGUXdpFU15j4t1PuIuiOKbaYruM0lxtb1uwtoxXPXR
eLjVBKqj9fSeOtp99pkk1eG/Brx+52QgXGfqxnCdiC50FiO72Mgl2Kod5UMQ
/v+9+mGZMp3+/I10coP4xGMnl+QsuKaAWSBwx3BtzFNtTm8ik3ZqUekT8y4h
Lwe4VwRiL5khZPhiul4t/Yzk4mkT5gZiwia7r6ICltHVWitUB06zoVvlODtX
q8svtaxXt+32H8BA1sGs2agM6T+aSeusUpRQpGASYAZNDPpBkqYhOXVMhOXa
KQ1vHBD+FUM4Axek0G9UtKyrxm+Lz246ZeX9VGfbHIqVeeBWc9MWiHLCSgAI
eTVAlz3Jb33W6nKEVPXEFQsNrYLmeXyYHoLzjaalM5UI3XPh+kRc3O877ex3
wYKbb7NMRtXIOHczDwW2Z6EF/vVyVRIXYR72dlYuz07HZoUSYfE0e7BhyU48
xaTwsSj+BexpnQWKD0zQkJI06hQcSb0Lann4SSHAegWVjpEaLY8KALoBgo5B
Q6Pj8LcrZhaH0BMR2uT+1snmOIN2GkSz4kSd9x/UldPGiADnIVArC+8lJHv1
cc9yk9gCTwEuaYWCcCK+ubACE0OgubdJnrw6fcIgCTqVgdpzeKYoBwxM47wO
WHbr0zaCz51b5tgTb8fT97O3dha03HzhvZ2NctJQRF45RxoAtUt6NfY+t/M4
IfTdK5FoaWyeTJuVXc6mCFFARAevgLkurA2YXFWB9TAr4gTruKVxjSkfCHdg
zhv5c9LU4IVcmdpckTT9mGYnJMug26olTil6YCQdmKOw9H1gupsFNK8yXbwx
0QTXlV+82tJzYHzaKpvcoBvYngmOMF1mx+PK7PQtBr1J4CCjVZDdgBIYxqH+
TNWznQTlJwOzatLv4EC1it8wzPkT3qW+JZq4RYVH+szd4ErUaV4bgu2ZLIzx
6jJ/uJCk2chG7dNbXAexygVkv+m24rZ+c1/dAhsjR7d4qywLmyMzvAqrXkEU
j94ldner5EPYLmZFxhBe99Zw5kwPz/LndTE+jcYJZ2uH47wKWEKzB3NnBrDz
IoSShCk1l4en5ODO5mGe+aegivhOdSOK3MUhM/tzQ8rbMKbHc1pb3sBOwhTQ
2I7gkMfwmSxGGYUwJ4Xe8UpYX/S1IIdvqujbv2+FS9uCXTH6lvaqVF6dj2X/
hWHh8MiAM2vv//XpZLwMekrJqgMsCq9vNEXFHY1rxn1Dsp/8wkzEe8dmzIJO
9P84O7meMMcYLrtEsE6UIA4k6ypEGjBCNVjTeG7a7/bffD5EIdiFhSyJ68/l
qlk1SxyOVxlV/9HNCS7GVs6Z24H0BtaD4r6/UzcDn48JC2QxpbMAPgNiMRIO
5PlvI2+yy4hNWjXlrQPWm2fNoH4ftAj3US6/AiNDEQOEd0Y2a+6gpaGb87RS
JIBGjdqWHbIlhxVW0EvKE2Ukq+63/pJ9peh7g176UlYPqJljbwSZuhh9TlRH
PByhtQhimZ6xmeCHyJe5LopgsCFbpKed+S9e53m2DsR3ZGA+PhUMDXzpO9ch
+klCp3JGj+M+CTymTs/SemneEyrZs5K1yhfmfCtNjLIL1OMlflhmamMZQuxY
+Z6GKRp3dSNK9E7nTvL/zIIUGnelTSAPbsB7c0hCyPPk+dUYPObTuky4areR
Zt76eRSrTJhs9GkhCvINlEzF0sYbFai+P6Lwhg2/dXpXc/VYOjZOjM2rmIbm
qTS0Ob3aSFhjwcxVojiw3LUPduxNsf4pq1CCTQ7cles4P+mLKREnUJssFtPb
oJ9IRUSwGzJW7CtHyQvejmz0YOKtEMU4zVHWtEVBx3v/+XjEYvCj6xWHUgsL
6b6wxM7aiHW6DD4JvBqYBYuMyKHaPf+GSudVyLGHyln1AGj0dJXpB5JonGnD
d9t2cmiKBr+UYTU4LcJiN1n/D8m2lyIflV8tsYQaDhwLU2SyRx/5Fgx+d1m5
JcHIkcJykreOnXwtp75k+/tNaL/zrgTKwTvNFiI8kJTcV8nZ0pF4rNLk24mW
7zHWDaC67hDlr/70oayU0mK3gw+i2pSgiU6psc27FfLilK740bH0RST6phFp
nBNHynoBZxBycHeUjzgc74FVZjWJ3sWePv1fTw0noEv+tTzwc/QrCrC+V1nI
uOoKhDPigO/mLuYUQEK39wvsc5GxQTxagFzANGQ99L6BjUrHaNwrs5sxW12k
9FDExaC5OENgdFp3wP45azYtNNnApyd1TPT73IeOmEu7JymuHadka9sqwKqC
OZAxP/NvklgF1z63vxuD0P5HrON27wmNB5VOWtpjQgULW/XZ3ixleJj2FdZB
U/OdIrw18eH/TN/sPEK/jj2JIKpYYQaKXh39O9W6L3ndUsyuBILf9oq0l3EB
FXo3LeeYmh1n2PweG1JirQnjZFX9i+kKMu4HXtF76lQgV6LB0W6P6uI2yZdJ
FXJCw9liek13wXd2WOPRDwhuacSUsfisjq7C0SDJpwjiEhURffik2azArVP1
1J8p0jPfyOLtodDABA/nKz/6JH6kAnG//oYOJmhptBzIkCrLX8yjXahUtp0B
KyWV70zAKWgKPbCO1eLwxL0XoQM5Oqm3YaO8LksLpzQtsS2qGdAFMPqioG1G
bHs8rH/Y/xcNpnHRtAQ/JOEUFCBh3j2fjVwFUmI1RcZmeuhLqS6gByd8PaIB
tYf4+wsIOj8VnfQteMpsCge0BG7+yLM1rQI1VLGc0P+WyZV/y29Oe/vLOdJo
nxcoLJJaogdGUc4ID+m/bwN7E++zRnbo7wcqN7wIRinY0euVw55mjIqfcxzU
VofpQjtfvVrZzpMMd/BnrGGPqjYLHpN3Exm9iytdotQmwX2Klw1/J/nbH23r
CCzwFO6Kw8fHPHx877UjjDUh5KJG9AlYAG4K9c8FhyRe0ldOmSAA5RjoBSV5
m1OV1SI3rY5yMT+TG9Abj+TlKUQczGU8/6O4V93WdJ1pvDI7/7j9UrUgR84/
DHbxaNHjnLPNvp1q+NH340Co7E6+wnfmWLbogQaeslXFyeKED4bus6v0FtcA
ly7pxClJACyVzWttA0IjDr4BrFIwYKmCGvXDvBoB/eBM9U4KPJ3niN6cyBAX
5BRA2ndcljJHbmWNf1AkIXBuwxftszGjshUGWr0KdDCe+WYoPTYtNMxei1QJ
6R5Gsa1E1D/oU9aahfw9VOR712sXDaIp7RCWjvFNTeR9/T3wD1hAK/ms5i/v
PGj2LLEnVEdKDah8uvdw7PYTOCWL7CNKgInxXcuv3mg+tjciJZqv0HU7QxCC
kIbJVoHGZ7Su5+EhpNf+YSqOdYafl5msJ1I6tmbuAeIZz9tW49zuatjAdP4m
eBdYWsv2HB7jiN7bXMhc7YOLplmPLxI486sfmBSCoujPk66U9PfU9u+YdLgB
djg9QufQ5Qf1rTgs8RXKkASaFbBBzoPYK71StvunOmi0LowjcjlnLbY+aikA
Gpb2rD+JzODeuTE8VbPkQcRk31xoJoTB25jHQlBiVaZvuVB0QZW9CyNTPEG1
YPwroU7D24g3eTECUJQXUBk2/khN4h7yJ4qxKHlyCTmjLGjO9/zvS5iTW0LT
RZCHjrioNL6VhDsMMvC3kAamo3nQo1TUFrkNwiziLXDrwe3yzSI+0BTIh/M0
g4IlFCIXfqGdL2Crn7jHoc7WopcbdOwMynKNR7seIEin+UhaH33QbaXDax6h
Bc0S9m17XgGUKe0GN//Cqmr/2EvQ8aK+rDACmDO6Mcnyd5H2bTbhwWtfnPzH
vvrVDOtyglBqP9u5a8Cz8jXjJQJbhayvgLEwegnsFEYNHT+Y+594UbLp0r8G
9EfXu4fcJuAFa0SkWoMC2TXfrq3eht15J0Aszkmt2SMfoOFB0wZoP8QHn4Ro
+5bm9NsaqD5H9KjcRFwtxhNkqIufV/wYuIbkzZTp+WFY/fF7YAEeR/RUsih8
/GPZaK3kyk7SK76dbaUG9StQITBoYIrWVfvKgcvuNpY9tV2EzuZOulB536Ov
mcSXRncqGWmmRE6NbukTkIvG/uNqYdExllbwDxXc7Zd6CWEN0X7pca5FrhPX
DXcKsFAM5JWlcR8Zx/4sxQ1tBEGFDH5uJ3tTvDT0g3tZJbLAW4ywsJ1wzGEx
KYg7b+XHFDlCaM/uWPZ9hFqdGG8qysx1KYHhXvd2ho4ygH02Tou7mQJfo5z6
3iUE+k72GezzUNcHaFY3gUzPKZLU64ozCG4EWYaYtwvLLVFBQwfcYNUlA92V
D+qg5AvwKjvlpQ59QMnrGqTny6Qb7wGLN4afgkWmDeH3NLL73hie1Lzo6sTl
fqUN9m1t91XhQsSk4agQ5vP3iQsjgS+Vc7lcZhGUC7VTvGS1rIYHBPSmczMJ
Mw1uW5kyGeFoU6HJow2ISgs4z7yZ+dUSME6l5Egi6p2HLveStVYvgni/TWD0
OVpAlkZvZM5DspnhtfjGO4V9Epzt6XAqIfsbmO7KVCsa6zhR3jyrBJIXrk/2
mTVFZBzlDnx+XCFxv3d/dQ05FG0/DmwP8VSEedsiCmWbOXUlE7WgqQPJuzj1
EvoTAvm6Ln8x53ETE46Er7iuTEwJTDip4bJcGrmpFY39z6oZP6CCY77sJPhq
uCyMDyhZTZLSktLo4aK9Sijj+wgRmfBzcYWRuaTS51DMsYVUqB4YsnFJtuTx
T+JiESIQzRcyFXGRmJpTYYE01B3T30HELYRNp6ad0RqKrqI3cF6oqrjmdNm6
VWQBETHlDg2VIX/v4CHtENQpvb1RhpujLBOu0frysc5FvAdBnuE0HpdFROMx
MCVB8e7/+Rvk0eCN9nvS5/9cHt/nTh6kkdh03ixhZM8893m4DtUU9MlGXkFO
4D+9jDSKgj0olG2zvY7nocpn9JfHC5238LQN5QdZtKiG2fCbJDsu4HwRgbZA
060mM/dsDEit1ZllCDCHjKJ+t8cIxyPLG+o8aeaKcu4Cd20/onuNZbXi6Fnf
yOQHjT6HodvS4S+jCoVXLzMBaX90CaG4bwbxXPezm7PaP/jIUxTzTNVwFJ71
X/TL2F5WIZY1FzBsRrpkNoBG5QBlzgcf48GO1sDZWYJepY9IB6xlu5jLrKEf
e63B8IlF38gXwYEBiDTEeEZ3xwHFZr0JOiEGj/+JrvT4QlkPZ21z1T2OpAov
7eG2Pn0b4eyrmMsSNeg/k1flZaTpKAAZOeLSQJkeDRmEckg2l1gxhioK7bhp
SHWQUrDc/dJuY9uRYz4jwB6lk31MlV+HMl9Yya1Z2B6+gj5yjMVBSMyJynOs
3okL7WiBIF/w0UncHAr4sc6reVAQxHA/VsNesSCtmmiiCb5jTCzUoq8UGsiD
vHaIkkVlR1LlfSZyQ5+jJLNE93LDYvvJrbASbVk+9dJyQKh338FDcgreKQd3
Qm3ISlSUT7nr39a9BYVhhKu2SFaSWG27pd93Eotzolu1T8ooXXHNH1tE9aYr
DxRiI4Wd94Leaqm7h+STHWdOKvWdY/JppQgexVOsdvQTnihhzvbbHNVPJyJ2
Rc1AMS+2Wmhrv60zrO+bNPy/XasoasIEL5ogHlT1aIVa3Mi92l6P0Y86T65J
gSB5c/JImKZyj/0MYDWhVrwM77kCnjQvKHzDIS6/FxeAuuTuwDrPHSXAPwFO
onnnSxJePLd4fuh+tEZcMyp4o2IN8eqdx+Ez0REKSBzzeRFP7P5GlShBqk2K
wNSlIs74HzzWjrI1Aacx2ufnF2EvXYN52EN/MG6nASdCu+PlIvBVUXXkxKRz
u6ZlAOJ1Nf+th18JOMxAynM75lGHYsL0e9/8sEEBVZvBbUq/VOhbsdDOsHc9
k7vmcWsXiWwJxoQTYrXaM2F8/FE8pvFYHEt4cZ1qkkfBRBhKUBcD2KrhxoA0
sfvcf02yJXlDB8beAe+ApwiCMj3jQNAOqhHLxm+AMKEEeZvrnVHBkd+9zAJD
RIoTIu7oUFzPP2nwcEE7CE5ksI9hGgU6Da1apT0aPX0Jtvwn72GJRrYUzBnd
wHEhfcpLbI8uradcELL1zX5yfQpOxCyxU9HkmHv1wjEhNb2bxJfJYvL459tU
yvZ9XgdhCBqcnTflkYSyOZohpQo0gQmD94FhsL2Rst41UW611xNM538r0ddV
bkHOJuvlB83brFtwhkUXr0/Rp8ZGM5TcJQdYRabsxLgooDMecTQj0DAHVxg8
1NejjvTC2FXCa6qRE+yeo4sDzMVRiEneL+QrHx2SywsG259BFjDRKSDJXaJP
ii6fNSineiQRQ4tD5PPer14+BWgfBuFEfUxyBRPpYUbH/zurwJe3WWSvcg6p
GPzmvzsVOaWNm9h5084YLadNb80ap1CdckVu7fXUj2Cm5pk5haF2Goc/97Sy
y0thkedTe4lrXpbcihkLrNK7L9MfNRKyC4L0U6ybavfeZ2z5DRZp0NOXJkt0
MCyyiurGAfR2ovqgNP67iXdPhRfJIYGDn0xBcchdZyPvR1dBvMxu3WbxwYh/
q83QAvHJxRQjyJ2524Er/50PcOKiLDErTgfecEPjQODsvcbKxOcm2Lb+lT6z
uDUsprtEfvsmVLEfIpkCfYP3qmo/SNTxT7iNbB8wjrhR2BKTs3XVeV8XQb9f
vgGpSzw8qgSXmRZ4OIq6UlGz2hgYTneSlQ5vv9hEBlHm7A7DmRQP6dvOTLN9
dFUJshfkCwoBAwid4TUGt19q60CU/MGhbUMemIJdroLawZEhgZgsiJKIUWmH
H4HfGKc2CQCKfaNCSOA+BPF6Hh5WpaWshO31bLl/6S0fl7lzsWKOHiXLXWzW
UsOyg9bJUKShe1FLPQnYIFNL/NmixUM18/GLUh1yoaNr35PErJuCZgzUtsaT
oPrr6PWwv3H7+Z7i++tBO9g9ebxncBNvMONvkJaFGbk1hd0OmKcO4ZjkSCWi
OQT60gdQvDyTstLkjC+OcosJIV0mAyBVCEE1+bfaddlwe+804UkMkS5tbj1o
qBHj1tCgYD9AoAm7HC76Lz2+DIyaTXa5wKHLHw2PZj5lWL8Z3vG92WN7Mxkw
1ASm5oUZT6yuEfh5u5FwYNhAzhIu8aDjYWy12KU7pdKaGIv9hGsxWBh2wt0T
mvJabwia1P6gAZ0gJE+ThiVmYgNOqUzeMuHln3/xtXTupXSjGvcFnDbz8r80
3rIWW6vsFw2AE2qfruFbOvnvGdQBFWJgPTbXYfKPMmTRr3+DFenEi+CkqYl/
/5LipWxkgpaO2IBpvw7eusmfF1OhfYxuDHb1n5/MhgvnysQFfrFvaVrK8wbK
4jvKwomuJ8vCaJ9wzlllLsslbYtXurIOkvrMHB8Dwwu13zmEvlwWVXpdgFvr
0/v8qiSu20ui20k/1eJ9jGNpgnXZ3qQon1CCUQu/SHYbvQtDTuhwBKZGp9vH
cOjjoLSjdOc4GcQ+v8E/BRFo9qQmMhZEiE0QXcNKf8Z1aLGgaQkT3unkLQe4
5w4vkoI2HKsrTh027G4yrhy0Yh1YJK+O+Xy35sjurgTi7m0EiYKmwOQhRL8w
eRW3nei+FR13SPTWxDhpZ6Z+9lPqt+T3HfsQrOEexIH0IVR6qcScEqH3/NxQ
HM6qygSTr6PdZWHf8yAEZwqNCni8FTm9rbmxlW4cQYIqW/mHAPMpHFOzJNFA
DzskQSz1gpoBR/mVHQ3mbmzRSPsheVgJOXJcsm5wxN+uJ+gKvDZCfWPgK1gl
x1go/0CweLG/NG2eLpLkj4W1IwUhRkLkXXcNdk6ShPRjKTCXamGzONgFysIU
eAAatBs6qBx03VZoNjM65Rx08PB87VRbAf2M4QhmdUvnYeZ7RpSqB2eOgGMu
u8ifBuVJdJzWq2cIU6ELYiuuPCnsDWMC+/cgpgCeOHb7slYIsQfLEquxhlr2
RHpW3Da8o5FQiiiqGUumW+gUJX7Pk/IssBwRdCKmjN1mOBqQO1i58qnS8mLs
LO8QyyesukhGbhN18vseiVp8nHheiQpYGW7fvGKFY1HYBzcVaWydnROPvdYC
pi3wTKa2fl0p39vcdk2oRB71Niv0OGjUFC212tJHujHjcvHmGbUWJIiThn6r
ipVvqt1FP0/BpKL2h/Yx6iSmntutVQj9SrE7QE27z+ax8RGgbyIO1osR/Ulx
gR2W6zUbAc20bHH3zAWptm1XXX7pMBsKp4vK5SNTd/3uJ44Hrz2AVxePod1S
6RhsbPqFiQsa/j8ZSTu4LX4aT27cr5SVQ/jB7t/540igzEM9PI/z5vJq20Sz
Xk6fsKi7WNQZlVEv1kq6gELKovbhiw7+jBXkopIoqna0mAmrlNpboQv8kKJZ
/njC80cBxvRioISBLEEz5zJds18xfFqM0Fk1goqjN3dG8olOBDgTa9zM63+z
lnRMhwEF/oBeqbOJT+S6fvO2oAkHIE/9RBNo2EyleYgv+zD8PH+rw2ox67T+
aUJDpb0E2tyxxk0au/xQFB2v9gtjcdKtNvaJL5CkSpcQmCtPItAdSi8ohRxv
p4bRetJ/CDkcdewyqxAE95dFFqkIhPaJitgysigf3MEEVbxJFcalxnwAPwL5
aspTFH6RhwZrlFQu1RYDT3ORuoM3yDHEZxjUx43keCgOXTpoWRahs1q49+y+
THoJOPNSQR+SGjwvWjQ+j5YCOZ73xWm4hXxububhEeZ8DOuoFoelqKo2NJVQ
IYvZUf5YiSAl8RSRfQZbDtsoOlmScuowWxuRfohP5aL6Assz17Y/Rcjjv3tU
d8j2rrKFxmfGvPn46z9KSjz071nEZi9L9NTqRX6JoWYvhphiT4KoeeAef7vT
vW+AB/F4fr8B0Nne0BjQv53+wioVqt5WwF3kkaSVZ5FAykGNOf6huSQFSkWx
oPKZg5KO34dEFwG+pRYbFAeGYbQ8ojDRT1q1nsctUQlcVoP5g3DVtky2uQT3
GFWWnJFg1sIIaaeWqoSzyRBfkY//w1D195FHJ9fWiaRonelekg8Mpz1ASYkB
aQzDqw+wbzZxQ+4+AROuXMfsvCxT4yaxDxyhPhFJnZ59RmIJXLiroainYunC
T2/rNKw7hAmPbp818rKgbvyzAhX9OyN8DK+aI5y72rU/z5vs43EV1GqPq/Xu
rvKGtwZg2pKw4jK4rsUqbQbJdv54r76A6GwPYnd2IuvBfYH1888tPWNSVM0Z
vKBU4DWrWchMbGY+ABAoxT6Z3CAlfzvqW7R+E9ktS9J52VFqGM3dHut+AGjZ
7r9BZAUByOT2KAsaAIUPZFMLAPZ9IaU3RxXMlfGZPQSoAXsQ8hSfn8SfZWTU
3QcCb5d1Jl138U/NP6txbloqGCUBpjSzRH5Zz59Yd33DwPw1WinHpHZvt8zm
tvC1fqFrDl4l3+X1tywODeQ2u3uDWAqLjB1aAxHugBlfB9eVeYC2/kbSrf2y
wNjr54EAS2jUfzjXoMXsMotUXQ4eW4aCL5UWS24WCcI0GooTRN57Y8uR00Pq
oVoeaSdLz6rxrZm0kAKVeuEeEG+/qqvF6i6ZJdMs01T9MENQu7ZwWma2vIH8
cpto/oorujAI8sANvVtlmmP9G5ygEdYK67j42Fc8IvgI74KicbuDRSSDDlhc
YiUkHoLUaNDaPwLCenpwEecdyr4+VHmaIyQAw3T+VqLHSKC6wAQWpqN8ShDC
Lkg6Is2WCutoDsvuG5qQF4gZ4MmBWOJYYj+I9t6R4F1c1xRyC0m9vg38Uwu4
gVdcZs4IhEzmdl6Q/sx0lldKsoXBlPrHGgUo+UdmIzbAojuOc7jHQdAc7oDa
5T4xvGwUDZVOwQfc1myaBPx1oiyeVsv4N+4Nm5eaaB4i0XlUeOJv0lIZnunC
mZH+xuV3xeorPkoWDtZ3WYWOzIz9QV1YEoxkEf+GKnBNLtLwKRWO1NB1eQ2b
Pz8YXgO6d6atoT85Srjd0ivbm2rB9n/aju7174uKzlaO/uhmkMFRz81Bbt5g
H66nEiDnuEZ0BkGVuFIhG6eXbWhFcQoygYzcZNxjHo7U+9Rh0CRO3ctWCfpa
J4pca5+jCC4HJKpE+Z4FzPDO6qWga0Kx+nrxGV/qKNVDShGPRmfsOrP2EFVZ
3iNZX5CfUv3qnY98CxAHMQd3uotVD8+yOzeHa61BVTduRoeekLunC5XvZ9u5
k7TOZmcO8gJi6wUhDlpRsvh0VX8PbYz249m35kfvSF7al2p5rRfUR1KOEpP3
L5cD+ZYa9AVvOocxyQjI5orkhBbIUh8JMEGz9hGVILI3s0vKT1qcunhSqCny
ZX6hXt3O4q4RkFtCp2fXwHiY9F7ghmuRBKeZJrfG/l7kUEtYFA+gZexJTgQq
9frercZTxyPmyT1FVc6VezWspL9Lno8BCGEet0HXQjYnOgO/kDfZULyqPNOC
GOlKTm3C4GmMhzYV1tmgfwAm/XSzuRahvtinZ4ETaEmYMaDsoHn+SV3YFi67
bV9jjqZmwoJxRgeuK1wGreUH3DLYoKff2HmIdGTf6yNrNYJX9j2XuX5WWz02
/UXXWnrwe8hsMsFPQyL8HiXwxlD/IXgyMuXxRga90/nuvW/MeH5Jxnc63Xxe
ELtZgHMzrEzH6wOCu7cLqeEdSTu+cRb/5kQ1xq32vRj4cD4cuk8y6N8A8Qz/
wJgKePj0bU6Jf8iQPPEZZBZVCM2SRndTBZKvhirW+B+wF0iMG4/LHSLkJNSV
hnhWAyrBtlO4tUb66eAl+U/qQ9TOBcLSTtpEv4j7XLlInN40sZGffeVyMrQR
43wpg3rZ0rR4lamnIJ1wwYlxQxohplznq7d/5nOcLexdkyIYOiN7zlqNhsdA
Qp45MJMPM2DDlYix8ppSdKvw0VT/YfzOJIhd3twC/z82Sx2VxqdJPFT7ocKx
3EUYFVvo/fQx61/iMcat3Pp5t061y21UTi2+WpUwnxJvwb7C9NP+lWbG5aOH
phVJFEccwHWCu5kjOOSKApqNrU/SwSyaX9klcLqJhg/p6anx5cwD7KPpzAvR
v7Ysf8W+9eepdupjZKITx0BOeVCFfx65Ogze3V3rZ63qKQ4ua7/rflRcnkq5
IVP+X3QmWOs2IxAMKTkggmtfwtVRQSs5QyfenhkJCa+PjyQsLxi6haKfMkwY
NR0G7324mOESJLDq93EZng5MX3aLUv0Iy6qPp6kx9jiy4jk65bfha5o55Wmo
d+TCw30XPXRLfQIAQGkrUylkD5+FnzBzkmppDa54MZ674JbLNgSFX8sDJ1wK
79GHRLnVS+cSMTdlUnv+BgrEOvM8LiVrEVeTpZB5GCcGx9h+rZshHeX4pBU4
Nid8JmZnddGVUqq6IoPozjHz8F1b2Ylq8suNH5CuOUUD6NCtC+NglhoKQM/c
QCLzebsTTF4wXwhQL3Z2UiNWxcmbJ0EacqC/dub3+EnxO7q8WPYhWG5wXXkP
AaFIDnhalrAt3d11xKIdV5uKd+6sKOcgTJC63oPb2Tm2oIv9bYs5gFFp0Gih
Ul5N7SrrZjTSUEBAZUx1VVVFaITTOlRIUNoUW0FPYoSI1Bj7dp/I66jJ44s2
rLeLJgVYRYaxSDtHfCa/YC1CVPaENylbZZxLzdI+tU6CGLKO68KfOnNiez0W
qcdh9tbSqTjujuvn9+ucYzGof/7Qg3Gs90XyRNCyZmvKrWW0oyFtjFijk+BQ
heicdeKZYdGhwcuNSLSp2EX7jVXx6rAluYYc3/PmvYqwy8AEoqL8oPMlWxe2
cATV4dGXPefQGmuB3Jrf04J6WADiSLW/THIWBRITcLXrBkj51pAPopX7L/cm
OMSJD3dL8/V8BvgjkQDNc85uNPaXSx/fX9dnObAxCkDAvf7eQXEQG7bRkY2w
vVp6NRez542EcyViPKr2Xt7SkZbH0LnxDNtOw7P4bVUT/GSGJKjTIBkChUQR
CdaldaVuqvNJvQIomlfR4+A6DVd87+IpJ7+6WYE8QzUZKcjsUyCcto80htMH
dGrvs9nGmTEsTGlkjD7R+22MCK7HoTms/5e9wB9weL9NxKFW/3AFxCOEC72e
YkVyOpa56ZC1HO9+Vdv+kmJPT54kG5Hd1JcYu/77D4Z7othrpOBVjFKYHNsg
obmVyvv2LQercNnoi8zKjDKAx9oRLhHmyb3c66OSZGpgBMZUqDX8EMoHfSLI
9d1jUMlXoEoL12rSpGp9lHNDHKehT2jHwn+rVnuZaQnYQWvPDZA/wfn430gw
ZbgUORRBVmGyoNQ2z/DH8v41lsZVTxuf3uHS+En0odNX5GbgPYmFswFLn+yk
rLf6mkiA48vlo0jNkDZdK/7QV/iLdZqQ4K/LV9sSw5F5eJ6Vsuf66o1nAmsZ
Rgy3RX7CuApR/3sZLWKyWbIAtRMkMCvXG3YpaSu8N0cxnUmux8RSiijek2as
YJmgyyPQb/+Q2wF7sQ3g9wZzd7/UsV2z/YF43sjbmVIy8YKEsGQ5kzcUH9wJ
ZPv5O5lNaZr67WzY961acelmZPOdje0q1YyqIaJL5Ru7CvSiLYAA47UoU03b
4Pq0E15ohDrmJQzpIW4zb/YHrxvP5weudvAeup4leDt5Mfmt8y4ktKXE2F+z
QMJFl0v/lIrgewQ/ztw8Nmo8QX4df+2MDscPyUOtuoXRka+diZxjwqdZ2PZT
LozUiNtpXX4KXr/sBqYPik0sYyo3Iacx1UB8/+n8ASPPpuag08w3IlohZhBl
9qZVKYjV6u2tX1enjBS69J+/CLRwXP4JBZjjyIPfgU1ESgxIXNkncD8BuYl8
7QUksvNJcgkrN0w8bMHa6RNtJSexoRG4duvjfGZZlrCoacTjsaGBYwx0Hf8y
4/5d7lhfNx6RHBUXQhUK43t1YM4yxp/B0vtyz2X8gFcrQN7nnS+Re/50hjoK
IfGslbkiFDsod4WG2SjhkUD/KGryBdMaIODDeC7hda61adaOItwejlSFFory
KXB/tQXhN6+AIHUtmQC60SFMdbmVbmI5vv5/sXq6AYQj+1VrZxRwkdoPk1ek
YTmUvh88W9+0J4qNMsb40XpRyaSOkRyYb/4G9jm+NEI9D5YoGmQ0Y9cKIvwh
Ko3JQ4G2HMo7WSRbz2lVQr+cayExhBYNw3mDDrm2q0VqQk2pfXLsBnDy6YNM
NODYiTD87aAbN3nOjAsdLucE7vT7jiFdND5d1NHRmLmWoYfdJecNKkQrM30a
zGUvjg1qGojDLRd7THvrv/sL0YxLXleX85Jp61k2jGtsih1daTFWYdECFG0q
XxbI+NLhJLxTLYg2FS2IT87nSpz8KsCYQg86oY98KwQ5bJavPpHCnF+Jb7zz
757yqFGW47eWF78ODeNyFRLoV6iDjro6o2A1UHdZBPw/dyV436ndspAbnECZ
MDU8Z3Zin9o03+mLcf+wUNmthaDX9xJEVYY+dVwEdpnYdWALMlFwByXbr1/d
dPpPJXMgD7bH1qZnzeo52EAP1IR5m/q0Qk5si3Tw08i66aGnDm4oDblXMuo2
X8S9/cgYCrSUwKuJhF15C8aQXCxOsrq7hhwEIPPBee0cidZgZZjGsRNDAeBK
GSm8tGoq/kOFs1WRIFRQGhiFm38uDZOvb0+PiblB6CEW2Z6Bk7qaaDKDBXv1
opW57pnQM/CIB3QDg4tJ4M8nff5Z/2Zm6s2xoh432tMTi/n0jf9DxtvDn1XR
LoL39sb+PLrmHodYeSMjT6Q5a3T0XWIsvsOyKF+XSsdycOxQm+cuVf4hmzKu
7AOqhbTxdLrL5x7JTrkB/RQ4PqJLkbXNKJuQrYx3RK9a09h9LcJDkP6VVGw9
HiTt4Hj8wnVx96koOr+5H18tER5LZwV/6rOKLQ44zSfsBKR+5jk29vhtXi7V
8d1MmP66G40BqSviFTj7P+f0vT9vXe0ZDs3umlw78oiAJ6vUDbL25DaeSg5m
XMLrFNTCdTU077LIrf/jRtMVkDawntFr8Wsm0tgBlwUMSGmpJXjrJi/cMzc4
Xm9x6o3xBi89AnG0OmY1d+dZCJfSlF+L+EX9P3gKFhLRyhq2o1/ZqRYp3AIz
QSx+EdGBNaOaR+Z3cFjCyxJLzJWKLs28kWuKXKkEzR4vCctOQZLcP2kjZJg8
X4RCzRaL9rZCUPfJmIqzWCAwnO7tO7OMq3dkx9398NlwFDWn1xZaj3bQkCOo
np2aXBGRuniNsqBeFsU9Ta8319YzRXTjVbqxrfzfCe/ZE0YMllNfMkm0KY7f
WIWWNlbCxenb0M3KJOf/aPXAd8WzAbL97cHLq8gBrt8+pui9pVfqAkQVxgMj
XiV+hSvD+lLkkf+Z31Hy6JoNNBoFVUxqCP5uq0lRXNtdbmyH5hj77P3lfX8X
XFniHQFN4oAmHu7Y6gUaEL4i11lsvBBEJv9quIzWQC0wasg4ieG9IvAleanC
kdCMWWv7g5PL+b7jQ6vdPA4fB0yWI+V8bf637p1lisiER3XxxYajg99+N6yl
mqc3shG1iahsnShXSlUnGg0uRycNOuziYxegDoEbgc8wiDAiPtJGT2jdnnO8
GEHQ/gwpwDhH3emiXrHE7dVmtJDB9oiL+Qg+vFEa6H6ydRfckCi7rt3b/kpM
rBCYIWpXWPJoNdjlZx+SLBGoUG+rBGgEekmPtLnEZbF7rBl83uDP+7soKyvF
YS2I0ZpveCAYhN45b4P/chOb7UHPieOdNA6HIgyoJP+HyNlC++zUKQXp2EF/
cPqUNM51HywNuKuFWfOFFd0Y14E2/9knNFiJVo5YPCHYii7ne9MHU1uBxwQF
Qb5TpedWbWSo4sfLBXiWgx3KyT3Qq0H2KBQPVIWBWr2pZrnPwZT1L/rrSm+I
TbxYpaxBAYLkkALQE7yH6d0vlimryM8dVQTGOhe5CC6+WnuXLO+thyl1uIbT
jZgpmGFsW89gp70jh+/r37sApUuCAIft08X3yi/hHcmyuThFBGCHiYJt24pX
pVId0L0RPyml77wUQN73a8F/o24vs/yHMqnL3rc/eVJRROeTIue2BF7jDogd
dUu2pLGiYH3bPv2GZ9wk+QcxepYnN8HLSPRMl/hRXA82X79ULnVEE/vNESLL
IEcEivBkBxVmj6R1t1jyQbIap0oFN55a966SHCQLs33tlIwTgeZ2M4rmZUR0
6lUHsJl5D6zcxD2Vrv9GsmAfM+jBSYdsORXbe+OwP8NBlEqchpz7dugk2n+0
t1yKJwSmX+TTZju7qvlsh3NhWfmmlTNkACNpqSrMlJW1pAwCoVo6wHpOSDxi
SpL/73KYgE1Bdw/K1KK9g5okmJQNPkzwUHuI4LaN83qlnaIq1vCdpgd24sU/
zQDW/8sPgXZjkfb+aDAaF0x1/jC2e/v1mZNZ+hi6mxYoAJxaDPbw/LmUU7rj
DbrJKzGmfTw4BLQ6+sqXufsnt8DkZjVYVs9zv98ClgT395/t1SV5/27Fve8t
/EQ5iaKaEC9IOSHaeOD/UcuDBjQ4XgcW88ysVxcpr9OEg9JZPBA0MDXIuUzA
y6V6zeu9qHQq+hPF1481A+O/m0qJx/NWgCU9HOip4Rg0NCu2prl48qIkTR0y
IRbpchwNuxqkzQwcGIvT3EBA3z9sUTU+JsXT/ewcgRB7X5T8/mdwKEDIfT6k
5OQhva2YsIl/uM1s8NSzan8Uxw+yRvt12NfHAKSK5yJz63tCjSewSXdDkE+m
gKM0J9JoHyxlJYw1KXwoKopLCuIZKEOf0Tx4RprEUIhdytoZfjfvcyZ+wrwe
TAzNKKh1nGIuJDyBoHg3EobWNLEIb/nl2cr09v0o4vbWtu8pkrU4MG2aYoZi
ynT+WbUeXTFkfjytqX6aFmiIhDkrjKQlGFGYnqNOAsPIqC9G1oDOgBD/o/qV
1VCP0uI2Ammaui+nojopTnv94/6jgcRjnDkcYyuHCFPD5YNVlnCEfmafjind
HPVVKPU5DiHWbdW5IEtrydOwfAAj19Zobi/3F7QAKitowfezw1sWPjn+F6b6
MS/tPWslhvUEFRidv6JfcV8d4dnGKhW25DCkWbEv9VQeo8+fpFuu2W5WxMez
kxzIRMDGJUoJZSrGQ02SaopWl/25DwPoTtYngVzTY5wW+eFJRr37Xf8AIdoe
7THofJXccb+NxwsiiCPuJ9z3rI0gQo+Bf0QyvFGLpZHO1M9zUIRo4fMS0OYI
7J97gSaoYpTwDuVhGFg+SU+yYLbGshGef8lgRn+qow6+AJ0AyXJ+e+4l5NIH
XWvFQ4VUCQL4jyPEa9QMb0qF+uLGUnUzeQBgDLnNNMHJm2Tr1GtOD/w5xpIj
u7tg7L02oiDR1e0d6U8m1RnLnAiR990lR6N1C3S9Y+O5MvaB2rNtZhsJHSeB
LKQvFodeXFXSfhrK/pJVRDmSmgi5VW0z0Y+6e5tn80XDrVyWtWd4S3ljqA+r
ELmYI2XqrNC2SorvytODydYPBkdkOlA3jVm4XNEo8KkFqQ1mRmKNJvYvouM3
9VUkwOy/vKDeJy2OlK6Lf/+WkcBSRBIHwhI8tDfgSJHui13m9v2aP8qZhlbR
ar9GnOsbIqIBu49oigwGU5soYxNlZdMWp/5s2XIpDteu7rdEPvoUPbTsMG5l
hU2BMKgn7r9UMtzJ3dJXN6w5BJLQlkynvQQuHVepA+f0y5wX/bhNNcNS2PM3
EuuokWg1IVPIibltIiRN3u0/GNkvQAWhjgDVGCsxRJWdFb3egzlU3JMTV8/A
DZjnKINPFBeVLYt82+9Ia7cFYbFaVzy9JSuWQ54coNujtcGImK3z5Uv5oSnh
0RHZGy0FG+wLZy6lAMK+lVhpandNd06I085lj7etLbL7N08lcwnXR5l2ZBCN
bmZMS7JSQKgZiHUvPd4q77lDnp3+dnP9niGI0bTHjsBxC5HRp+WtfpV70Y/w
jHnPRWO0XWBTgj2pbkGsJIyPQbR0s666qdsPjIaA0yXI18LG56s2Gow0LpBl
O3LoYS9AZ3b7Ych5yGEJFbnTGXcCplnmcFswVt+0TDM70t32BBHdREM2/8ns
Q6oV3wSISZ1EFbE6+PkkDtSd/jz8h5U1Y4FWzuGvpLjd+dD4iNEUXiV05eer
uOnr1C1czChw9HzIrTA6hy5KcJ/99+AySu5dNlOYR93yDRVQTcEJcAaPOnjW
EpNkpyzVmz7Q9yM5wz/3KTxnVsMybNmkYSKyy/E/ASBDILlnpgdeiCE6B04T
KyQSlqiiMPQIhotTCCrmQInCf/8yuLrIznZ1MY6Z7Ub3+IgiXkK5re/lGB4L
5DzqzvJIHAYlONiuAw3Gh7LkzYJ2PSP5a/VJiVyoUr3PT+MkN4FmADycPxjA
faKIlIv4qAD3OpwSaeH+prADS2B52Hshchj1/sSz/VQQBsn+hP4uJSBXLSHU
j4zg2yhnwvEQvdZzujzQ/OM/U8/FtHoIl3SLuaAqY2yf9qLePVTU1Us4rP3T
baEH77tPBHDlVxKBlasI5/4qPNWiAXhXY4ZiZmHcjwXNoyeFmhppksiLX7hF
yaps+/Pp9LnqLP3qFXDKzKPoQkg1ZqyM48IwzMjwrqkfcjwZVnxJ/0Fv4yPi
3Whb1l91ph/L6vc0GDnQCn+F2IwoTmwQGNvH/aNcxc7Ry44aODVRAYO2l+NE
kjG8vLAvVxZct8YH+dhuTZJfx5mRSh0zW9vCVJoDKxh+ZITPYKMmyGhJtTlY
a4dUMhUdJFDPexPK+meNgBr3Kx+8g0qdkAtMUmKybNr+I39xE1BVfH21kExc
zVXyd3wJX9fknsCf92R7DZR9XaIqTbzFj22fUE9WvV3gL1V301qHxTYUZieW
62VhJfvbruGb/Ly7t0AXVLDPolnsSrZQdd9Cppl0v2vNDO4yG9e0CQAmqbXf
7LjFeSOzkdemnkGKMBD3lPf1kktfiT0M5JvcYkr+a6V+KJMxlJc5zbp8D3pU
xlwUshGlaDduOYVw0vGaE/8QLXmd+XiLrox4RkXbk69VXGVbjKodYPe+eVB4
+EjuLTEQJdN1ee4br9suo1rwvNbMh1CI89sOBikPJQ7tdqep793IMlO9hurE
zB5FY31JQF+pacOaSNGfwgUctSNNbWGhvxQGvqdtSg10Enca7Az6e77jZ2iW
Blp2lky2FT+PdaL2bvp9VExEt8pyt6vXMiuH5TB6Fg5sqkD/jRIYulzeeui6
CTt9tVAwGdHDaS/eBfNifdMn2E6UzIF37HBG7NpwrhPHETZfHKTzr+n0FXpS
iXg0KgRjtXL4soLYMHtW41opgYVRXn57kg3GKc8xCCU03Ig0ICx0Ds932vRJ
AIUEDIerfP16e2JiVCAZiF4WJNlbLJGZunN7MIzI9w88uMdAor3gBKYDQ2Kg
ZnAQW+XgkuLUV5IPLf5hMEjib8vThooMtd732VX0kzpfVsZj6+aQjtAx4usS
lisiQsVrarf/lRgGan1uLYqcK7qKMGt1Q/AZ/G7LBcntA582wUCwHP8aD2xs
NuMilLmOrEuqyP2/6baPsCDSRARKISLPW8lb9fP+sjNpfa0Dlm9F4oz40LMq
mSYTCChAyjz1PMhXztk6+S1DKcgh23wqcGPmuUSrPRgs44GxHPuBuGkxHBKd
0qrfV9GuMa4InPPeEwU6mkZoPq7MDddv0dDU1oD54NDv91WLFa34Xc2TdUla
a5Akje3VymAEgLda3bjRENgYl47iJZvs08AZZB99fSahCnnF8mg1czz6xzrQ
u4Qyr/h7TfSeDxHknNEyM8Q/HoVRZ9VQRgyrN6Ecoa80OjhH7pEDE0336qkb
NZyddKz0SWSI8QX9GV66fwXWjzxzL3bOwiG7c3TG3cImKBr1L8yl9e+7pOI3
p0pe27z37PD0rmFgzSgeY6qy6KJCG3/5nd8qtYvBkwD2eaeN5SWujOTo6lU4
+rMJiKx6GsqTjnUHIxUzygsw0kdpTEwmi7S9Kx6AMf8fC5ILXhQMKhnQxDG3
iIoCAvmu7sejonzhhNJ8lisZr9N+etvfOBIKn4t244BKX0elrFKydOkgEIEZ
2qkcVZf8sDaKbv+YpiolhcXXP6nAjJBMboQxWYJ4Pv3SD5CtzbBJi7ORrvZx
QvOqTvpjbRYSlEPdL5vvQFYG7rgi40gA+349r7rRZQO/pSadkMH5sQY0R64S
D8VzxJHVIBhjYkG7iLWdY8AmLNTaIe7Wbr+ODW7q7hELFYG9WIH3R286D+3u
kAP5NLy7GAkVR1JexKt/PbE61SGEh2DTJEKw9J0QbdPds1g+51jv8ylBMpZi
KpIl+vsu4egXEQe8OozwjVXehye8z9jv6EWKoHXF0kZoQfjK88B5nWlSBncU
+yg73Y10oGftVX+WLjck3m3EFLFQ6PyJuAYEiYAY7BizLoTVzeAagBrJkIrc
7fTwomB5FrTkkgXtJz7zuA+Hyf0C8M9Js3FDcUFBIBlj1TClofJOe+y3M5MO
N7hwSWsnTZZJZr7XDTcDHCW5JCK9LHdHrBKrAl8SHrghHScJgkX+Q0sv3eC0
Mcl1/w9AvzQvLXuL/RPGE37IvKZHRNVuqbuKxNXZ/smkqyS7rq78TzdsYzN6
Rd/wsffUGMVYMz0hJ+qKg4c9i5cLffAbiQlkpr5et1ZlJ8uQvVtDzCTmwFTu
yNJCy03CpAQOFKDl/PQtzcQlrY48Ycva5UJeW+USU3d+ArB2BId5AcLpn6nS
i9lJhQ+RmPSDOBt955/RTFmZl6lwYonr3L0WQo1Dg10r7i+TgJvRtpFyhNMc
Wzmbay0kfKNqoL6VfOF/c+yHjy6AA0Pv0JGgQQ6m3satmzk+oUdGxlFL0xyv
v+RQdV3LmfUUII/R3Kp5TybygB4BFZ5e8l2J7PAymRbmF7LKS9HqRujqFi5k
wIrJEG0i8MDdg2Fmfe8q3GUcBptiJEUbAZq5i1pLx0wd6V8DdlV0jyopnRKg
ZRFHOw6AG8rX9f/WgjrvvzJPhdvuzm2fhPrzORcTD01EdNDWcmUrJCSoEW8t
1VOjGvAC1/Ne5ZJ1jytb5RwpIa2zX2hsLqzvSADQrzAAgAbS92FPZefxP/Hp
m3IIC6CFCbKKsU2Ptkxa8eMisjhHDDphgAcduiqT+tITt9hUdQDCkR4H8jFJ
kZ2EMkROc1nds+XGLGz5w3vD97UaVOtCvFVzG0MNRYuFkATPaC14ouF5GQg+
R5heqgW84MaWeuJ9MoA/yBe6xvrY2y00V+cGlmeSQEwrmhudB8QcNc6w/B4Y
6YlXwDtXJ1EvlgfO+O3ifrXaofjD/q6ONtNmWX5LqPh+nMgGfDF7ub0uvVbo
GjgVAl96DaYPTL87K/bXsskxquXha4KtRu17J7lMc7T3e+gF4wy/w4Rd1wJ6
pjHVUoIIk3fnGqYZNiF3GiHC0RxjfsT9qp7II8vGvY6/dGfsP6CVlvcG9rWR
wxUxFcdQOIdX06lxn/Yvb3zUlIRqSIUaSS9KgvX3/ILSS3xFQG3v9t7HbTxi
jiYab5ZPm4Nxxm8yPb+c/S5mw6p1grNcOP6oT4MdGl1Tsv6SYObP7I0sreNI
ModFWW5hphiH3+Dxc0PeYlYT2c7tOmgEVn+e9UdWofmXaaY5D1bJeu20aAwr
LAAnd14AmLXQOjVVtszwx63RC27GHT5fxu+PnOOkFKcEY7SyJa7w7AIW7JcM
dEC8YKS39pnKaretuCn6i1aAFQznkSea+wne8Yw8ewKedvVJsV5QsnYl2q4T
z0JdOLe+Kl1IaSDBNFyTw9sdeOfejsPcmucuSH5E3/vZaWHBhP7bY6/OJW5t
1o8NmtXBAaqSWtudnl1mLgKWoPujUePEi4oknRyanLUS6DZqPdsOqC7HzcjI
mBYt0k05Ps2K6U4HltFBsxTE8uQ8hq4vgnrIPFiCyAScg9QDpm+9aHE/gPYP
URdLWKpZ6VBijmfSUxgrCEWMecoFHzVepdrv5i+F97A28z0cnt+iGhM7egtQ
fZWi0ysDaICspPpbKEpbqd3Utk1SMUu4GpLW5pkYmySrdD+YbfA13hFplRSI
GOXdIlCtyLeZXnC0/tQ6Cyssq97nezWq9t0pSjNm21OjI+q33r7LMlI8Sh0z
ApvVd/mEZzqr20bdNjdyoL63Hr0nKvVDm5aTIzkUKx89tYC/IU49wUPawpi2
vmf+ko7N6lMLUEz1ObKMNtiPsrsBFS4yuVEIxaMIPbCM45pcBeGa1YtIa6IH
5Rz+GA1MOqT9ycnCMOoJz3APAxUFIS7Y0XFUVqsXM/NGYluV+3JgzjVdVdR9
h07SAT8fJljLKxFxe1ydTyOQFcTds7AD1g6wN/tbfL0pL6EKCq6ISaD8U87w
tPopeZw3umkpF4DeK5IhJAb0aji2xS6ZHcyKmkIiDHSc+k2znXIIqblJbNn4
thEYKkqWCtbIZwOsPhQXu6Dywd3eLJYs5868yi0mRbS0TDT1Tb/B3WO1KxoK
QuOMy9c0V5us2qQB1y0i+5RFNS/DLkg4MHK+2saL2Hxxf81wS9Ufl+FB/bgN
5HKJOraolQM+4jADhT7/nBthhm1hAWWlvIlXpWvkULIJYF0+bmwtNAHQSvZu
k+CmPvlZ7rfmwuRugVncb8UPlSBOS4e1z8DwzJPy1+J91Fn+0iQVLxpMY+ud
mojFnwW4j7WgLMreWILz/kehzlLqwx9MTTxGL+0EqgZe5NS8ROGNml4uvxJK
bI2GzVTvt1bnu3uY6yuhESYQAqZfcnumdgbFP1SLIX75T0At8naKhDzTGRe/
2FJe2PZqqOFKgK6Q66k7OL8V8q6XWZLx2Ok60WbTeHgKip/CGrBIgmaZTK8b
JPz6hVeKbfMOcgFR4ftTVX6/HjhdDLcRjtPUgCtAOfM+4519o68orLXyIHnH
GCH9g7COKdYBkxXAu1S1jZk191b1mNYuGZcA9Ls+OZ5/3wvOQbCxCmvdI3jc
/MjMSH6Kxxi+CGs2RQTgqcf3V1Jp7kMEMBp/z7ufeMxi7b0CsCiBtcy0Fxd6
EXSufecmI/Hi5gjKllpIOVooIcQWFiXNtaMBL4WTkTEuKXcas1bBdEu8jIEP
qtrUZOjLGAGWhSqBU4HHF8VZTbAie7BMu88KrWmzaJloaO6bLzsGJJo+pJkY
x0rJV0uZ6BeChSG1nFN/F9tl63cGu6x/9vrAiWSUCjK/ME7okTTcw5GPZpB/
z+++dMfF/+IORG7JMmGeWsJTtCcLHHB0BE4HIDx2IOLyq1iMP68Yr8DEB7tW
zS3yTuUVtL7j6itvooR6UiToalWBCUaNIq/9yY2+YW/tMOtyydYWFiTT74WX
M+4W80NlcsoGtAqZIMJWDOf++75bcOzfrDKZfyXW0NOIcZh/BayGRu4KAwAX
4G+aA2Fyb88UErsNcQzFjV/w1gOzDb4gccfCuBmENrzyJ6of2TrcR9d1rrR2
OZvBLCuAxNd0Zj52HcARVeR/kmMLiQ5r5Cs0UaJ5NJvFv+vpVy6qnIXMlhh+
+0tlcy9A9c9UD34/eoqYOpbOC0soit/65koTAmeq5NYpDv/NucxbN4bAJdMl
hL71KWURabBBVOtxecWFWt3mk84g9oFihx1PK6cFCWrz2V2XIHFrm2MnDCkC
2qxQt6H2a1C4beUArdy9+BsvX0sBAuAUcG57xz23hsLPkYo+8Ri3FM2YRz3Y
YUNFpFKaDGpYNucuXxCYIbaJBXWZ/G3Ed1DI5TTOP3ioDjtimIBhk0F5Xz0P
v5EcxAiqziRwCpB+TkIpD6KcshKZAe2TumL+SA1Zh1nc4y9T0wPpwEKgij9C
h7ukRQdZwymyBuIDJDAFVTABvusd3NktuTxoeWxD19d1H+jLxgeoTyBiDmoJ
oIG1yU4gOAdR9OoLHtHFqTGcvs5H2d7Qfo+ZB42GnCSXnZcbWOX6Jpub+Hdj
M0JZ+6Z4mGpm+pPKE5+c3Xns+LuO2ueBVtQsUqvlpBhGe6R2YxoZKT213Qpu
fCyiHSGryXubnfGepw4xSSbUwz5e7IhBikZ/x16kMKnyYcqCtKK0Z03wHrQ4
UbwAe8g14i/bPMAWHcxjySgzAK+CpvhbkMmXeO3Jm7agHNW8HhNjNJ4TvZ1Z
8oWf6256YQ4itC6C7b4N+tpeeUHr4HWBLvhYWR4MKMFX2D70TIN8OI8V0czY
hkdTvfz8iESNVAM0cZJkwb0qCP771vG93+4rfpCrxzoQolH5AdwbnUCDe5Iy
VcCNmFKP92UC5lxptSjGWwMMr85D0UyqDYCHcdBFhnPICSZdsFrk2awX3rFg
uNOP0wzKwVULAh6PL2d2TZ171ulUz/ZSDvzzWXawHJ53qUW4IOVtzXVcMofl
0gsofm1U19ZuSj9QOeLNiVZeNlWHg65zXwHz0qax65zulKqRNWs3gSHsrHfN
nBWsSUTPIuYbzEF1OA5mJlq3eAD9+mArUTgMD7KukQz952YMi6R2Q2TpUHxB
EF+Mliuv6+07GHpHOxKyMEfSlBm32DDED0Idto0/ere/DA0LSpHfKLCPf8Ay
eX7bPG7YhCfl8lKq5gLhiGcuLbGvne5C5xo8AZqlezvoCYO5y/XEvbEbdK6e
9WQC+r81/nXI0rAv/pzLEUWiTA14pPg06H/u5ou1/CPVLlVmR9Ap8qJ1e0Si
ObDFCGwJXSE+aTAGUuh2dEXEMI7Ab8WvKpGzb6qdCwrFl+QKof7TWmEsYTUv
JjkP7/ry40hpnV6H9fG8YCrG0Xk/gXMaqNIpFYhh7bgYkcBqvh5NlNgPkZLe
lS+hPZrNtSb9uVWx6pQrQMzGmxfCq5+hTf/BFtwb3qoJNz/wVyxGLZMb/0o+
3QVaCGNWzlFZEnKaj7FWeZnERy87bCxMZkosEyl/Gv5rd7Qgx/FlaCl0R9KE
cPZuGV1S5RNEhMvAeBe0Hma8lvqFhkgD/Z4pCWk+86jDSUP4g0wQDslEG2V6
ItgcWHh3+GYEv8MBbCb6mQpTVFvPFT3k5Fra26n251DTu7HNImMDWs4TBM5U
XBE8Z5fjpQw1lHbo5vHHJxwoUBPo05GiyDlwMNxsPDf3f6msPgUrwesKUilq
afOn/HPNdvuUxhkeNSDta6wrCA2sOrE8kdTPH+DFu/E0mbrRSrYFsWY3bwbQ
nUQ2/bK/acosTyjZrqwoaBL72epBcDX0X8ZpGzJoS9mNmVg8Xa9RhbWWYZLA
215iLe0iIUEpq4FJ77BTR+GOu010SM9hNUXLLzAbScCVNmeDHqtgl4mXj9fK
lspI0TJrd9j51E5t254h0w8MPv8+jSW+0mBn3CKxKtNwou2WKg0hYy+FdNxz
XLo8e/UhiT9AYAVo4hwS8cCp0cW35gquPJ1TK9Q7QGbeyqpigOBv9NJKbq+s
pIHnZZdHIxyZvVT5b1keDCToef9BHi57B3mn5PCbwzlkukZ7IVTMoBVGCzYY
iQ+DUVgyWuy2npd2yvL0/W8tRBsYHGF0VLoW0kAl0G1mWu1KACl8c562Wj9k
wzeLpi6LTWm1gr2X6TQkaC/3mzggXkiTTjewClANfZOX9SazHzaJnrhahWCg
XTaxS9av3dzZ6brc0E2Y4HkbfAxnloetOWNYbXqnkwC9I8wd77GrxwcvkdEN
8gtwP1BakiZtJb7JmmfnjRxEBFV5vNLdR+shtuaij1L4dVET+iZgA4a2jkSe
j/gCHMMKvZ8IjImc0M6M0w2zJOTcaIPYuwfuTfM1EIaQYHjg9u8fv0czFjs0
kEUrv507VmuNgKWZVPAkRkghdDch+X8q0aKRjivKFZaIXfcEH3wmaBmFhp2l
Lf0Sn+K8JNE0LAgCDs5km+bYpm/4qhsxNEcH3kYcYIVdvwwcQrmyqAnsKNDI
GagJxFThx8kQSeaeibJOuOCDO92nFL0wHd3M4KFIfV+Eq+EC1GeJgZU4oPo6
YEqzDEtvRzyRQpzsXpWM0GmnnsOmfnvAZ56ADx/rQB2DEAIfWyCGcfl7y3ak
pyS97DGG265NJDGC+3BeHqSNhTK6iqzkUEs3+Nr0DsVSf6HFysovQyijoQHs
dSHrJSDeCsvfBnCGtIyVPqmwkxsGAau11NTScSpzfZMTsiLDWIeUDkLtfBMd
gUbZpVQr+TNC3/uhV/NajFk52+W0LMfiMbQG0+7qut+iY1MRSY9kWWs0e0Mq
f/sSyzQqb0BfDUi7f6ZTi0d+RRenZ+cNg8xeWCZHA+K/BIgbSWowRxj4HIBW
ujZXBh/XR15mNxEBaMP3IR9jF89Jj2UiuROYEQtUtx/noymQHLTSfknOzc06
Wz2TOk0ORzQKU54JdgN+ryiv6DYXzYKYqGjdZYvT0z0ufKbZAwBmw4arq/22
TDl8vXH3QpkVz09b8DJPMDWfCa4+6cFiZRcvyWzAgEzNO+Gtuw0vPcHr632L
NLiTxVrRBLahkQh0AxdDykMh5GNO4l7T+h8SOKVOVHzcq+AC

`pragma protect end_protected
