// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BUc+jrIkvmilKaSEZAL0sVBHwkRkwo6ltJCWxUg6IX8n3sOGuVnoIpjJvH5Z
41j+qqO7+AsPECIc8xqYmuV7+Rf2AOdxUoWWYVkV63ka5+jv+mXZrNGCKvmS
jVlIk2R3A9i/npzqyh8NDfQXyD6KdGwQ+Qi8OHmaIL9lXe4AUxH41+ySUyDs
+eaZCnzWaLBgE84KMLHbkVm4eLhT28QYbNRHWsUveIadrN+Mg9xn+P8bfZeC
e9S0ekff5fjl0jv7fCEoWltKCzPVT3+5DH/f5dGTmBBczkSESnqnTb3ycQHB
WDg30wajZXSUwsxPmAoRzo+OwxjYeBY0ql90G3JHYw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HXbHWnc1RDPC2y/RFShw6IrIsKDqXIdQlhvm0RcuytDobI/PsNPw8QuvCwi1
VgFru7y9T4r6V9OSEhUDf8c8+afq6SNbLS3QQOZWXSuAAqWElMw0tE+8wmFy
0K7U3Q0tdprtM5BAwv5g0095iDrxfASZtX9fkN/nW6vgrWjTdXGnm4vpZtjS
bYFO/ZvFvDHxhWakj5UGL88PbVJMYKH3A0w36ugcuGLqSlwONVsDjU048YnH
IP/ca7tWqFiyyHL3Cj8dpWp4BD3lajOFAkRUdVrVpky6lxgXuB1ibr5Xb+pG
KeyKLKqiMahgQtYkDofcXIfrqF+j8xNTi1orVeWm6g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Elp4uS8w4+MPYlXxtAPd7ueQSxNWw63xifdzQ2RRFAreUsw4OIZEJqSzLXWR
fiCmyIXSEIcpeLgPyu8jww+FYZvCeQRh8lFmaNnq2BTUl5sflXJN5PXysPPm
W7xaYFGiyoGP7PtBHjhk2zI9PhnjC/rs+JOUtSVfi1/vlVSlshNwGgjY/bjt
uUqU+AbbQGoOJ9/duBnTMVcX9OtWx2+8tEpyltPnJPcquwAR8oo5AxVeldQJ
+jXgCdG1CG/umQ6rHJ/UkOLr05gKmp3nqpzkgaUjcjyo4wPu8JH3ERw3kRIi
eJe/NrHaBtjMOErtvtonG1t/JJlp02AabGheVw78NA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VxVMhHs/oeHM2+Bin9Vc0B3b5PHAdAOyM81+hG7hwu7nMRB6XrJkBgUFIacn
B8b5O5GXwqkj1Ps6lemqdiYL/YauYMSObLfcEpQyHCBXZZ0feul9LmfGfVU2
7PktJAKzYOVtwtLUvKHLLZ90CvTMtul5DS6L+37C+fkqdlCZ83I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jvMJEbXX5E3DFiF46i1JRDwX/UwhwWh7DpVhG5YE8DeuXPJQiXijqqPjZ2xj
Pl7y2PgIcNLQXJ+mO3L3oAoGSEvNOoKq7Cgh3Lh+LNB2tJZQSeufIlJ+3kJg
PxpUa8DAsvsOH5oIOBMz0KKdYVSj0HPCsxhZZubg0yp0imUZ+BniaqojsydR
ATiswbSss2kHCxA7LX5EaiMxYG25kJGRKhnWXfFz9kbtID4xxZZqlrO9YbG6
1LkNwdhH/iWPfjxzx7v3Tg1MA/m1zm4XrSjnDQeP3wqINEacIbLjcpruzbPG
LNxYaeDGKE1sqf/7NcFopmqi+txoakWqro5lmeHJEtvqj5IUtWC6Sb0OSKHY
IWJFx3ohAqr6LD23jNY9XNTjOjOPw57rbbP+CP2u2eeQvqB0DpfTXSwj89qf
CLJuvkfOTZsBze3PcT7EXl3I1LvPrWjMpOfoXq2G8zzdLIUxe/JMy2kp2bep
nCwUxAHkHQv75ovKBIfASTT8vaeUz+0U


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RJNacRcxfJsiSM3SVGkkyd/YJ8vCtwzVItyiX9vm3ogIKvsLQdSKl8ffzi+B
niTcCnhonVzg7Nmgdhj+WlCV4MH6FedQBt74HBgoQB53MoGqC/RBjFNn3reQ
b7xNqZRUB16o8D9EOpGm4Bx2GhDuM8tNvi3z8P0/fdR4VAsuTtY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i05kLZDbGE3LsFF8VCZuMrOa8L/VUkVRay859RKO0JRpHwKuvlO0sur4C/e9
daJ15vZGISnWeCX5YYPpZbzOFcoGmhtbB5krGcF3LmLu5N2sVorGWfSZ6JP5
4amrMCyzTBRvhkyE8bqHP5gikF4ZqNn/YFd4tApotRuJsZzeWM0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8880)
`pragma protect data_block
xJdFTD4+nSOO9E+PHWEZt8aaLRDB6M6FQ2v8g5oraAe6SCrUvrnRhmmRWk5b
bmHiOZ6/EVWxuup8ZExJtp0vVcQH0e5GKUC1qnPH/YFbxbkJeA5xqAj5AYjY
hbaC3F2qnIZswl1b1cHH4OSL1r/8ZpZC7/+AyIU9tkeDewXi4PsREYiaV95I
1otW9EnVQObHNYWHJfGeeCj1Sh0+TiJyKXPwXHd6+FOGZ5POB6jPDio2bUva
YEQPTlL9nfQdaRdwBfXdyr8vlp2JIKySbEsynBe39DnprrRdPwVuzuOEsaT3
AP/ekKoareHH5TkP4uygS92VMfVoOP/b1G6cyfcvUoh5alzf0j87MhFuPKsD
JXSEUA9Lj7NBJbSwLGB8khMm0HuQzjIUfLUGd4b5zpXN3vWMgFdjJsXeOxT1
o65Z3mdrRdE1ixuWWcKOZd+o0JFaxqVxzRkMFBEjL0eIYrCgb1WcFr6GMilV
N053CMMI/6ZyJSkY5n88Bd/p+MH3Gt5y8xfsnoFrpTNwqIH0goSywABCs6BB
6v6Rt7NPHlafLCE/UUBJ8WYNKsrrAUoqKZcGDOXUKQgdL/KjmDtPkOpBfjCD
nwDIxIHUi1wv3aLJI9DHwJVsT8J0CgPTiaq/PkRdcI31+9Aj4b9ZXbbOHQtW
cOLJtaAiR0EdIRc7Fu49P1lVZtPjpIND1D+K78fgnNsw/Sw2xUUpiROn9HAa
uBPqc5xtnGy5r6BN43wZogb3+rfqSykIU6bjScy+eMRxau2RWCpJQXbOrmg6
oLzsef5zDyqgTMDji+2UGdlRpAbIdPl5TqVP38PnbucY/qA5A6bspQA/TuKw
gZhq/IBZQ4KY04GC1BuuPW3XH/A9mKyuYQ+zRhJ8KfozRVZo0oE8t7IlURL0
BWJKUBlKi7G3BuHDFrriPH+WXjA2FQTCyYx4c9WEnFvhdF8qTjwgODlsr3zX
1FmYRZktzCcF3LnIP96H9FTjkTkDvAEcioS/+I7aYTAIkxznLMMjN6gL/R8j
l/fISiH5VxbqLse84cvESS0xLQqUyIlaUUWrI9/6xrTrOTQlID0V4/yK6NQe
tYiZS8Vclgf6639xxV5DbLz6NkO6bdA4+ovUvwlnlwchvuJvpy+AiiBlN2cC
NSobJEK4YADTx6/KrE7H4mR2oy9RZ1AxyeVLu6tw3KJlK+jy7Zak5cRZlLFv
wqgHZN5A/2tBLuUoYQkny9pBO6POXfZMJoCLPlg9kcAW67ojbvY5TZCAQ7jc
Wdvx50SoDS/0M/r5kp1S68efLX67CAua+RXxkexEPiIfwZOqQM4QduWEV5Q9
6a8DSxDvJUd/JVfHN2n5swMcRVBKsEVzHx4EU9PlJ/MxQlsS8jrrb9hn4Q3I
+sB1JqoPvemjL1kDSaq99NvLJyH9TIxx5FCjKUs5ule+E/sAAXZcWbzorelo
1XXuBGpz7cEVQ3vnzmn/MuDBSBC59ncBClyYLLlyl00eBch/zeSeo9j0vr5r
dhnNAiCYQcNL8sVx/LuTq3E/A9R6MtywWM55Q2LFw9DDnYKjNAjArMTLuAXT
gRb1963S195f1JFHVYRu3b0i/X6pyLrQIefPhOm+Jn9vcZOGBXQ8O4gyOPZv
QfzejlMQcXVmvu+U3ZYlA5nvShYAJn5TyM9IjiuLR6oc2OI9Efo9fJrsDwgm
9Xt67vb5zi+w2Nrz5txHzFtn7TDe2mZdiZmVmrDqvZ8jm3FEeMQeVdf3l7o9
g0zlIv9LehzdQvjm3Ik9v3YQFGu6ktXqkcPkUfdo/5y3yBOZPXko6ZKK6/UW
M8fNlSjhoWHIP1oTLqpol6mD03UYChA3+BcgbVTNhlzvNz8uCML0pnGz3kYV
Ipe/lmo0bfS9OzBL8gpGYSk96PANAhEKGsyrpNeSPRhOV5O7Nx0rbE4Y2YPN
UQ9QqbcxL242/vDCMFewWU969dq3IL05uskeVd6qiOZ1Xi83RDznxoaEBxgb
Z0WMV3XkviozbSlT0E7pyGtWrpD9wqVM1lJOSBdUN9Hr8UdpveyHqGxr6nx0
lKDrtJIvQhpXnsMvOw5y62L4owMc0sPI10bcPQcs1eRhIUUQpu4K/UIq0maY
6JtqrryF24eZ2LsbZ4C5R6d8CSZfxX3hznfa0u/ktaR4selD77xKNO9eKuwu
Mxy4TB/W1kKFjtat+5TOV6U6O5QCnr7enqHokkzR6uoMIGHK1x+MfydSu66K
6JEBYqx6UEcHXsN+yIRi0n1OySxZmKtHfhkp4maM2PFRTIcl0c4o8P9MkIN/
cGA8TuHr+B4irlO9BpBTEilnkMrrc45Dx6T/EVlyMlqYI04Wl/RoMtuxYJUE
nQgE2t2crR+Jyrfwz5y5KDDhmjxP/uRWe+PvArDLADcpgbOm61xjBu2MWr7D
aprgFor3Ph5r6YbUUazHnCtAJShgymGmXIU41XWxQJAwC2UonNArysqeCR89
M0Ndnff9GRlYJ0PEhptNjHZ5rEFQ78orzPdd5NSLS0xIBzn7+UBB18PZ1QuT
VJxobiTBGLULDq5tMJSwlzonkHN+P3LqGB2x7kwLVF8nbKnu+Hr/p+aTQo8o
eIjcK+NXbkAENu7YFWlopROBDBZeFwLvrHYwrnsAmjPPvSlrqEIeTqhI03bH
cNgDj2qtKEEQxu2vK4074IcNOG+aKCYVSbuliMiChSkPAYZTayJyEW3KXicy
PG1fCTko30HC0PTJVenEhZnoJ0B4OFw0VWC+vzWby830iuIaJPR0HFE1xkya
+Amc4kyltmUxkgVe+47RlzhN9DD+t7Hn4WDc0BeXMcKIX3PrtF9ggurcsJSa
H24zILjNtNFzEW2IaZb1jm/kykZtB3aij2fXrHvNyi83WZwr51ukFmcrgleK
AHhu1hUhPzRBV4bZM6FvW287W2g6pdaQdoIG6J6CdKbAHeWvvkjLdlc0J+wg
mQRlTfaGfPAsGCKy/PNPVjIvxOwy+NkKPBc4eeAF76EO7CBf3c6Z3naj+zLE
X4Vh+5BDBkniQAWDnvi5BX8u9xKajVoWn/qto4AJzJ7vVSJfSkqbdw5qyjgV
rMwWb+bLcXtPSGtLjn4ntgiG31eXaexitwEWddWOno/AuiV4HJ+QqCeIBNgQ
LpPnrdgF8lif24SMLz/9jWYgKg3lTgKetwQM7ALzlgORpckHteW5zR5k5AUr
jBdBQ3/JsQCwlCbKX5tLhLPvt5ssOrjZZem23kLldyyn4KBea7dojvpOjWuk
BO00KIAVZaEEf52OvBCsJHXUZlJmWWFek2Ur4DqesezjqO0JcMserUrcwiv/
qOQCOoQZmJPYtDVZCVyXctKeVUvq7k5M0ZG7/FYE3zo1rio6WGh6TKxGg36r
oP0tXWJOhThPYXFNYA9kk0FsD5qTa7460sZbrIlOpDMWzPzZlUtJUOGgYK5G
xN0hFJhsEWZh2YQpBicRmOtmXDVAiplgeW6d1yz8bkRzU4q6r1yUJUYd2mY2
d/+Yyuuowf4eG8N9f4cYcmQxabWZyBZwlEosoVOzQL9Se9jyZsddWk/KdjC8
fcf0UmmZbgrIHyuVGteXWLF5bZ84x6GTcuKeg9HkDmKqPlXBYDTVvxouw/Bv
tmk9eE9p9/M2UxKNzg10YFldXZ2/4WcVsxTbS+LtR9TydHHhLSQzrqMFxJQ/
jtbcfPYCpOjHkwfb58lsJhuvtwun3eLyXrS7VBFuK+Z8C6C02W7F6Oi0zO2r
bdSdNHB6xhmMnZt4sz8UMYSALbcG+Jj8lFhf/hK5HDZcdoLyfgV6ZRPANesk
9rt1tSNHZNnl7fjWFx/KRbL6+JUVrVeMoOP5XTB8cO0J3EwpIO0tFY0D5D9X
SY71pYTVtnb0zmyu4x0f875aRoGZOYyX/TT+pjOF5B4YDAbsbKlEu1G7lP1t
jxTclQw0Z85LTIYdh8cc43Ii8UbtDUzYM3hZfsWN3LdIfIKvitOM53RY6W6v
HRDyss3WBZuktfhhAriELhdpohc6hZ/pbOHG8nSbjGGf9bRp8ntSjjtso4ap
kZ6C/e8lOa8olt1DQ3fXN7RmVXtiZX9/7RIRjfUu5gUcWSpMVtz+P7uYq5IJ
nfeWTdUkHlW88JLvgWHzSt+nFs6lYbh/tgAMjAs54sEqOjplDk7F/leO7JkF
0DuHiq7FVaZE2hTkmsFMf7pJLK8fC/j2OX3DXHy/u9XV1TQHh9aR5Gx2IiwW
0c5a455M2lGBYTDFubD7Yb5c/baE5eoezu268TXNwgmN+1ZRa1xeoFmRe13l
EagRkR59PmX+qWmVOVt5S5DQYi6WlLWHFtDGBC8svuGmEs6TMpKHEeBG40Rs
ZC1Tp797rQ+juo0kLv1PatO+r35LcQ4gxnatfxxZy4eHfE3G4CxiKzcgG83m
pdWNzmgbyfTqqbd/Si+kzNYfd6ZFORrmj8eFKO6Cc1DqU3q1aYQrcbv3EvB5
2PzPwK+je4klQK1qC1udCdgoQmEzcRN/JehD1mZq05uQRxJk7iXmZHbdBy5m
UYuBo6DoPy+l5AsQBBWq266DQd7eQ59ExdJLmt93UHXo7SgQsg8hXlIWd/Yv
Yb6+p/MvN0xIDWNS6/keCzjBLkNs/ewhdMOxxYUjiDWQx6tSMtpb2zgac+S3
vkApnJ6jb4O2w8+tRSZ1c8sx/q2fBFqiaKQZFPC4uFf1ROybtPV6CyQ6jVOs
XV8mqAqTYfih7n2Sl0DtVvaqKVuR8oX/UH+kAZEj+W1nNe/xIgjTp3fCMqrO
wEsPNIpD1jtU3SWTRhbTFA241EjbxFRDssOHTDCeNKV48RNGL2Cvijo8TS53
hHH2wlg1P+XOnCrPDzkpOUjgmNBR93Zdo8g0zzovZZODz2pLUZpeG+czjskr
WSOobfQh5cQ6Xx7VjFsOVi7dWlCIDJBJ4yLMr+oaQZ0V4tE73xFlHkm7VkS4
pFXf409xEuF+olMgX0vJNRF+6yGaZNYGv6JHdwiRZKaM2npTaR+09YBu3wCe
PP0929bUQGL0sxjimc90WvE6ucRoQapMu1kYIMiHjDBn87VCWoBQyORA/wAM
SK7vA6p3S5OqldIKndthBEux0eLNJD/SDBVfi94e/cBrQ8I2i6klJoDXG3Z7
W3ASZ2U49OdlU45U26PWuq555uWQ2PbFRwBbIbB8dllKRd2kFwNi/ay5EV6Y
Ma7MM9e2htWvzNI9qDL3up4rrauC3VhKt6p6TCXEhMcoDSq3Fh9UqgmR9OhW
mzc6UKhaCuDS3LMaJgPUxI5NrKsr8Ca2UZpHFdeubrMAablsMSzFXW376dV1
scMDevrqM7OAEakCX0Wv1NKNBMxBwkHgkyPT85WhwqrzIjwR8A9e9NynFJ7E
ePhlKEbwOObKbPBkeaYMSAo2zEajBJ96PjgEahKHAlb3gPQ5OOBKQSgNUf2S
KRbHsoH2hYHAcMoir91RtTMP5BqNUIjCR3cbGaszRnKXI2wIJUbNXz8DT4i2
lcPly6SKfJc3XfdG7MIU55lWIprKgzGiIZCfbUA4867HdoIfLedfvTp8Jkt/
/UTElEIafEE07aY83d0+XaX0cH/ZEZInpXNakjchqgvz0+Spy2AlshxVGaeZ
ayfEe9hUQC8v83Po5VPNSt5hJsGSV+K3cNixqCxb/sM/fCrnBQnbUiJAJqXo
JF1iMCqfnTsBJ+peag6e2AcR0Sx/I0jibqshwUW7EKtR/CyNhtqN8miD//BE
HW3uxGXZcFjLcPX5h2teIJME6eJWXOuhfQnmmYzpkVT9H6/Exq+rkJ0syTwz
ztSH9sVyu/PHC3Ov+s/Kecjz2d1+GyJwE39d3pmMpkuq7qguuHvWdIo8jr4c
sS1KVm4EwSqayeh4fYvIM52yoBh64xAAwsqsPCFHkhy/VxD6qztATDnBbCnS
x/gRycRvAjnxWqUrSBLjqjg2RgeMHwO1/FP/JNRsokdicKIFXS0uEOGo+Qgn
rwRolWBam72tvoFX1E9vw4+WmkY8axUifhD/7QVFZSNAXMAkI24XAit9yWEY
KPpF0jXJofkV2eFRvMW1RHPDbAgnavNzbj1Tl+2aQtoMj4E2r5ju2yeUuLF3
z+/rTtxeftDcIRnnbyGEOnqbfJzlqJH4V2PWYdSfd6IGXMg20hgjd/Ay7NqH
ArjOWr45Bf8NnnRDNfxQ1yVenICDcQ6YRlC2kN6CwGXOh/5FRot4LuvrnVVS
fji5362QcgURiALvwhs5ONHNV4g8LiKdlJJF0jfVvekbQyNo27SGXgi/BEO/
E0xZ3qZ+FKDnSeWct3pCBC0So3kRSdRIRn6ynciGDz0awJ3i//YKTRlcicwB
jtuNFliYhRgQONu3VUHTA/d12PJv9rszTBVhejatceqWilpn2BAKpZsSLzKo
B2RIxIYsFaTVMs0TOBOLcZaLf88qqYkyG825k8Q/XqU5U+yDJB6hAkWR9S4x
iVvhoXpJU5Dkz6stgZih3DPi8E90Z/hwLQF0JM0zLyZL2GY+YSbNVJYCUGbI
K67GE3mm8cl6SVi9jrujlwQAEHo5AQwrdBbPugYd7u3VFeMEgM5Xh/+eRKbY
SeckEyV+Ww7HfWp4tYVA/x3n1bAZK4dK/rgAKjSFispA/v/uwaABTm7SQqsm
1nPsAXfMgH/SY9Mq7kVSkYOJrZWRhO4RCf98Yka35zj4y49NuZPlGu+yJFfy
dIKZvShHFBJVWWHejTFIPm+hIVuH2IjaErSV6Tp4zXqXoH2LppuNfUCyMLEw
OYr1bMXhICgiIHm6PgAsQh/NP4qCqgLBNYYIf4lBdqwjLme/+xdiGIaVJaLA
noncMeZ2ENTcyuksNQwxpCDWj8S1OCZQviFrTYm6HutQjl9kAjbsGKOiGySb
MEBG+8YXY4qJK0/hXs7lvMlxMusoDl/Gor38eSbjSKsh9kuh0NexDdOeRz7e
SoSJ9WEciwFiKkMs48vr+lXP9v95iWCTAFmSn+2L/4ZpabeOxrbHhshx8RHq
ztm09fmzj49iiJzxWLLge7ATOaEZicHpqGqKOvHsp58Vs0A0FuSnSQ/GI5Hg
mobsNNZ/J3vjmsTO0JZG3SZhy5Ifc4XuZ2279YS7i6ejvv8uXvjN4AfIZKsD
wMMVu+aDO0zKLZgq0CqSB2s2dBSDEr0PcxjOqoICOBhe5JP0wvjQqvxlvSP3
7ZfPUveW69DR8mYiKqHy0gxvT3pUb5w0G1vIOqWoNVmGmwHdikHrP7Uq/w03
EfINvTbM2mvmUKTIaaQao5hzmrjM9OcoIttkqc43y0mKP5eTAsRrbQvRWg6r
l/Jn25pchL8Hzg4HkAhah2DtOmB2t6titS5WZCGNrrcYC47+qv9ulFoB+dy/
NNuYoXbT/jaIZRd69FIgNMwjY6enfg8PgKMG6yR9C0SzWLblJSIupbrivMqD
45bzj9rjgs656yuOF+A00zXuD1YzXR0mFPuJnqjPPcBkEHOi5mjkTi8SFU40
lk7nidNmn5TbvZraOstQSbNTSD90ImJALV/eyUo+lx1+NYvmrHr5FpKEA3Qy
w2YiXafWx7fx//AOTgcKFEKERmcdyDxD3YZ1cmI9D9u2CovIm0MYn0dl1ZD2
qMNz7nSjEI4OPZxUlu+Q3Dlj6c2zlQriDchhct5s8S1GITQMQeCBhmybYZxF
0v+eiGZj9NoexWmdl0ebEIXjlvXMQ/ibcYZPx5A372RKvyFGX6YF1/oH/4rl
ydJBndPidYSIrpsGzRk5hFUkPvmCdC4Z6e3Hp8v2I/s0ja7FaDp3QJA/Pw66
SUAuJX8Tj2ijkLL0/VLsuLKUUfEZI/raiElL+3pePtdx6ALiqWTL9V1OdsQE
W+8jfcConI2UHLP/cI4ePtaazWgKz4sdI35O7iN1Cfvnakd0Q/dkDfjQU4+V
gHAhFKWR4HiLRnJLbvb1AdqARLZUzdUT4bpjTH0oiImC4ETmu3O/bziTbvwH
a4mUd5Tn9g6hlL6qXV97B6tvTBVrQDCTI50e7OflyXTtrsyZRJVR0na64fNV
bjqKUejKJhkfdTaMDO/uEzeM6HVef9mxAylPCr1UBTSKRi0M6pEo9M1V99uL
VBv8iIk9wr9p3jGtUJtQUx0GZg1J3ZNUQyI1U5f8lbu27cKLqLBQSD3GkWnC
rdrHs1QazOLvJRKDC7HfM3tiWyEfcS4WjSaVf5jrrLSk7x93UdDumUkvtNmT
mcgER5pe2zOcc7iLtUPVdQxArOU+9e9XLQjVge687LpItIfhqxNuI5hcGrWM
RYXydNvX+mY4agG51UwcCMG7HeD4DSH0WZIJ4X+z2sWdup9RweSXJsy3xmDo
SqqV13C8aSDw2/QPrTiczOOhtSkEF/PaD1dxlfC05/IYfp4UIcVJlYGNaz+n
66zGbb2UbdygNp5fVRyXFNgMXGtwfNyxiaRE7I8blhaPWhSSbvJKdFPXnZ41
Wq6UV9vomwf2dOscAVhOdcpIu8T+ldC9PHx3NdRlUKyTzRSARfszrcMieJ4U
OoJM66cbkbJjrhlknLl4DXeeqlQjzKa617zYePg75WOCva8K4FZlFFCeuLxd
+tji5Ag68BOFOMZOohN1eTabOEauusc9cq5fkmCl7XFoQxBVDmoiCcOY9P6W
VgjfQp9RmMGcWKYraRZdrVFRzdzozthQvOvDhy1kKa95D/gxFz48RAnEt7H9
5dV3Jrurvn5KuwCZ2FFxXhuFXTDZzF042rtruCGdR38MaLc6CcAGE28nlQ1D
gzJ+sEUg+W0XE2hCwsNbUcWqcJt40O9Q6Wk2c75++0XtnUyNcT19GyNBGSKx
5w+Z8OkkLaLDaYGj0/KOQC5Ibs/HkxFgBOhxunI0Qw64RroMI+vf8L9BRWHs
BUhInNQyU2CErfttIINfks3n8Vfq6/i76EY1mErxU4eu8N2INpE0cLWtpaYk
4DGLsTtUo+mNQO91wXxeD8/bKqj4qvVGl3K6Yj0dZdOMnf/3xZEh4HWQolUA
H4854sc1sRPSlqKPpwG+oQulvQjYy0eGmJj7nOBjGxXUFGJxzD+zMlCTzM7I
O47vm53v5+2amdUFgB+EOKJH6xWkM2qSCVkWrjVpOfOhUCFuoHlCMqA2EPBx
+KYQW8MlQ0ZOpQsNfnryRGBIK94vwt6qGuYFxqGbo2CQtUrW4TQi6qf86mZa
ODU7pVF71+YNEpb7+sW4Ovv/UAjmn3Pr8/tDVhpBHNm+scW2KjcNH5MhBLTV
WdfkvUB5I6gS0Vmb87vlPyeOSh4VbjoD2IT9VI2u3rOCTCjjcF2V58eUyTLH
Vw5sriE8t44TOoHinCfL/jf1lHqvAZzjy5BBi2gR2U/olEC7U7BlW+SDy6SG
NfKr8mpESEJjWyYbE2QjPCsNoWYCCiwqw4dxIVo87oDfm19mW7TJONZS5Vjf
limxzvM8AE+ALUGUkInMzHElV+Itwc1eI/sSJJ3lZEJa3kQofbdfWGQKFmwk
CIVerSyNAi+m/SbruQ8yKDyZk+RobanJ7ZCEBNCI48waeAk1rPKc/c3QeL36
+oqFPr+rfoVYLmthrf9/eqQ8GQkHlOkD4gFcE3PU8W1PdNhMwEGUjxtbkX+m
yKp+qiE5hGS3eV6yCDVvLNe8hjPl3Sb8zeQuvMLlcjSvz80DrDKhEQ1H02Jc
T8KXqiRgWkWkCzQwQxE80ZPp/USJUwhwg90qPoygJpjAeunWJ6WHVS+d9cpa
bZFAb13mmyDM/Q/G5VrRVU85kYkWRNFd2Cn1fe9yJ6IO2wpowmh7p1yFmD0G
cpQ2v8kDeGSkpr0mby06yNts+UrKBB4LCOaTIkU8pQ/YuDUicmnjAGo4F1Yf
Dh58XG6bqnRg0FDGFk9f8kjAKEtlOF6j9Mfvgi3cgIizhcpWgQj7R1XyPCRJ
i2EHkOdIq6aDaLsnTlmqjudmcyVJDsisQ1tN58WVM5jBDhIualcFbdFDgYL1
UbEecI8iA8cp1muESBckGlO7YTgs1DX2x+wjSI6Kc0jCF/o0lQm5k4gVWGBU
o83PkCJHvtBFX2NYC1ZEA3LjNoNfu/Z5bSpmHi3vH0KFshOFmtpuGRDDZQny
Uw88LkOJIIaiNSaigfjdgiilfy4nyNn1CCxLxluEuLMQqWgAWxT4OclkkN9e
mqG35bH8Pkq87s4E2YlLFEs1zNZCG8CA20/l6KnX7oPMpLaU+WlJJFbwuuxD
7dI5AtoVQO98QW9rblGMTlldAdXicdxbnJuK13pm3HmeNuQIIDTr+rUfXPGK
jp0UdyvUGMBrtUOlABczWy3B04pl30lSSW/N+6RWyXCLpRpwYwNpegSmpqWu
yo3SgzVWQ5LAbBO4LApPGqd65PfiPuqL63yAV1zaucHS4eeYiFUeAGcd8V4X
UFKfPx6/P+6XjMmlUv4ymAUQw/vH6weB82SrK7OIw/UNAt/kch+aP6xMzYIc
QFv0FGGavAmUqkeBriYUgAY2OHL3ZRB5w055Fx+7r63avk0vhJ2B+4yf1Zbt
9GqcbLtLSUCqi7X+kO54rV/VQZ2sIpWak0nIjt5+FFNy+n8O6h+JHE/BWQNY
1zXIBu9JQulwL3cgGfKmE3PUeW/PazwMZnmm/C7DO8QWVm3NjP7FJ5y7oZo2
JDaEVt0Wy2EsZrgV0gWfNo4w7RVtIKFgcVVsTx6zcEZ5z8R0nWmOUkST97fV
OaDrhL9uGJ+pp8wWLYdGZo/PqAZR5NP7+6uRIePoFuR4ov6QPBLxqXNtgzb1
AMt0PEBzdcf0fRvqCCyM7fI7BHDbWi0FcON8j9IYfrQTmMScTKnrSp3cKE4k
MY6NRGWJsXdc8AwoRF6HlXjlSk+orrtbr4wmXZ4HhKxFhLqN+zWvWcDrARRV
/2PIfYYfh0UPF0GbokbOS2L/FicwdPyQ/KG6TEltH79sP1kBLrSPCL/3h3LW
UvnzdmjcZoUt1IIu+E+JAPfwy+j74OjblTRLM/vJl+7RG8XtsdJCEabmsJFw
b4gcwWcHt5qkWJxdq8uRbhoZXT6T8LviISfNI7QX+Z/FKsys/xvA/y0xH8wA
IjZaSlvJ0I7suGoAHwcs+G0YHDXSYlatGUkreymZU/Ypo8oqlIk4U0JjLpX9
S7QSuDMeF75kg26eJTnEaLtAS8LQCmrqm873BmQpyv2Fl3qvDxaByzwNXeqh
ZEJDxK7MXBk7IigXl+3YtKoE7q5xHc4t6jWPPRNVD/OhTIRZQ7DGj7GNVYXm
qRa1p2H8hmYXh+HIr+shrhdzS8IfTjqrIFdRO1mDSBhkHlekmMCu3XtVvhM1
jzwd/swJedUBaWRrvlHSkf3s0AJWbBSrpR7y5yYse2fBFWs5MEfVpSuDpF24
JHkhN6W9aMR/ixah8zVAIjrvAsC9G7CSRpimgcHDNP8UPv//PJIokPW5sAqT
jg3Wpl91Bm188Cvek2a6oXRFZfIUcOr0Yy9ZHF7zrypcDXi7e/NB03kfj6Xj
IXqCBfdB2NkKq5Ck+c+mSSi/P5x/oD5lBtXJbHf+a1doecHnJaxWCqmIgYCp
cuBsj7sV5nHdZt8vFK4snGLJdrjYPbFHvGlcNNuCRL0VHkFeHmjxeQWVoM6i
Ke1DgPLOodP9R9pnI5VlRdHYavemDIcAcMRAV+Ryzg5dB7QMznVuVp+aFd+v
Wtr76/QAEZDqK6BE8Y7/QHCtEIZWGSTWvxXP31Rdt7LGUoSSBAEEShT6RBJv
QD2hQi4a/nSd+iIVnwF872ckxxVa8WPGNt9OiFg5VGQSUaYSai/RghXqAV6O
1cxdxo9wdyhCDjstMlTKWNdgx0kLsOc0v/PjE+KZ6etjwDd9w/HRJvTfjHRN
YiyxRx8iY0U1mdSbP64vkjmbRxSpnziPKr2tS+cCE8zm28/pt6n0XZGk7t4v
wdnOIGqd8mCCbARqpBRT

`pragma protect end_protected
