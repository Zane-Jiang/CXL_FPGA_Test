// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
XunNq/rR4kS7A6+/aDHoI0H++cbjneCSo0EVm4WwbwBKqEkw5mBZMOD0QCcw0cMJ
fkex4zqWVpAtNmdJbU9l5w8JFABOrMMuxxtnRx1gae+LFq8UH0ZpG89cOujK+URI
/eiySuQ5mb1wUq8idKdqyY+Y+FitI3uqxbKXH5rFCMei6azIzhwEtg==
//pragma protect end_key_block
//pragma protect digest_block
MRun0+7SYVGqklrxo0nQcZViNb8=
//pragma protect end_digest_block
//pragma protect data_block
K5QFZ2lbpk1B7L9ieKXJvY3UKg3iuaPtH/I38+5pRdFDGQExra/58JkZPbV8OvM4
G2IqB7O6JVxVeUvDewrC3/hFjzo4QVDLxhMHnoP2ypGRYs5jQkfYY5dyP2cFqte9
F5AWVyYU0xfvt6/kSLUvBKiH9PomSyXhRhPgM7wworD21yzNC94HGwnPQRTQsGWM
gtxkj6Xwc/GGsvEU1IdhpKrD0t3hoFCfeaUimqFeuDcm37krkKAgc4vIHOdG8M8l
A1WpbsxTBpGMPMsTTcKNW6pzVB18p0QGgBuTR1eolZlbkSLpg8NvYk7f7BK/M2zd
oc/zJzg9zTGD4UFVYAeI7x6M1CQtMMR09DMF0wEZ1UBBfB25CMIhVZCNPgZ+MZs7
PTdcHuUtGWL4Y6FnT85zLN8heXwPGWLkfqPq5ATXbWJLvBHt0pJ+Vuh+bjchim8D
koxUtiDk5oGXYGBxcPaQHl+l/mGsKQnzAquKjH8s50zMvdEQKoy4KI3jD6OYBxnf
clW/CW3eWfM/AQa95hZI38RNvEOb229Z/cmOXUzTt0HimU+8DxchROnmEYA9GoMO
jCsZACfzXwb/4Bz+VO5BlUnwrQ0mxt7dCsThN3PtdXfDk+8vfn4/BLBA3oNMEcfd
jk9tUTf4WXjzldFE7vrbLcl7uqDtnM2S7Jvz0i8abL6z6AzPfM+F8mIRD7yKj8zj
fgLZGT61nh/JVcHR59h2tLSzqz8Li7tEypOouhVsAsYK6xozKvuj4d4WmtlZ+Szn
oW1XwvvAmuRCez2tMTdTIKkdzWBVGKc20bD8wjCbz0CdWlraiy6nQFkD710W0oSE
VIIDMxvHhiSPlmku+r6phPwHQ4tqfypLVa72YophvofHVy0Kjo2U7BSGvNQmAYdF
D6cxPOFG96pBVTSS4hVgS94XbmBuFwg5phXC4yhuPBpSWIZPJSbVvtEglxsw7RbC
BiXeLuFtoKKipOrbwkKxpuK3Fa2XKtMUEEIMT/Vn/VvZlI11PuDxJgk80vR+9OB/
HSIZn7+bRihhTvd3x6pukYttkF36MyCmWoCgdHNR91FJxC3K7BsXMdmUkgLh1xN5
Xh9SFoq8m2bYRvBQZEXaNHkYqzc8GGdzS00QBJ2dOLvO+HECWY//JMLWZblBPgCp
88NUQcaJUSg6LiTFWtvwCbjL6eOmz/QgAGNN8aOe1C1PNWH6AK5v4CQ5HnsNAbyT
9m6mKbrKPPy7nnc8cC4NCPO0cU/Zmp+sfPrkf0Abv6RWq3aKytRCkmLcp/sdCrGc
LhD9I71lYaMirWuLbv7txSAJ13yDrHr6VyElp3zy5nQpwprWwvoap6Fat8Cx7NNg
0fifXvkbdmlZXLRDGYQGk219xo8Nww5qOg7k6M2YgzDRSrXswH9zy3HXO/IUnan0
1p+c83VL/cgHwsBSPo6DjggK4ajE8q/vel3kLCLH/MRtVv0wM5oQgjhlBFbiVpkc
QGV9hCAH2KH1rIB+pyVdw5pMlVKIi2q03B5tS84prnpgunro1AbzyDTGizyy3szS
N1JIwveeVFyFRdm/ozdnmxjXCkpyuzso616UJVbDux7gHpAog5AjF90gxrQHr2a+
WLqn1Uxq1nUwIjVpPA6fUgMxVFBvWRjhkpA+zZ0qb4CtHfHvun8dY048/tbKeTQz
OAdADspbZ0lT6P7nt6pwFq0kD4O/d3jUToiNJcXY5xsVQrOW0dFaH5xLVM1KFNis
fy7lr77Gotv3Le3s5pLAc4v78bpn3Se0mY1XhOZNKzzx4a575+iV0OxnMQSiQsyF
DS7syiyR3Xdm+yEknfgQ+zWEy3+PnkQFuXoGuEidSe53xIMxSd6GBymvHzlbIIfY
HMlhELpKMT6j62oTeQtKneLeoRsmdTYz9aSLDLGf1RT8zkxkkbAaM6CQxf9qst+M
Uv4qsytwj9mjwG49SU/W5GUEnvKx98GbGhJH4ZyhfPiDMZGXZtZlOuMrfLg++Ieo
eGjiIItuQ4K/mRtGwFZEhR0Q6vFJWQ3Y1vprSgugPvrd/MljeeEpOKC8cTWXLY/k
PXePlavOD9cO+WXZ1Uc0XbwtnBrRJGW7/bZAw4H0bC5PPdNvCy+iM6sq4Tz4q+8T
T5w531xAddMzBZVaD+KB81XZ5/4Rl+VB4p72IFeaQQw6MbJqKNg2T/8kGL2Q3aJ6
WqS6mc4Pcmah8fiCQKL1nW2ps8csOvPP/bG1PA/xZ4cxtAuSTxnCRW+nYr+yF8dN
Z9sxzaHAVYH3GArO40QUlXdUiw7sTci/tn1zhO5BIZYGo02gh0vHbmU+YDDvJihb
EJbxJxhKRD0j/RzSxeog6z3qI8JLINdtAWbGEdwyD9NlgEyAvVVZtnvPioW9F15p
7sskwyLrxc4NaDJ/LjFkWydUsDgpsKloXF7ijzOzrOMxvD8uLKsgjKiMbL0ycS3u
2IocpkSASkXvsqY2FTRTk0+mXqtU9xK9cpYPTSK0+rzRuEfOFUlocNs0NvnoQuHz
31S8sQv6Kn3vQ8F6sMiVusCfwxa8KH6as5Ys5oSEYSDC3SrSz0Tb+RAWf/3EQIau
G8BfcPlB7WvGOch9tf9X1z+rFXo0OSIhtHZhale982nln2bLPRb9ca4mrOtbcjUv
FNyZ+7uKGRm8M6+T9/5kqRAl8gK9GTCwAqWJyUEcqYGYC8U0NJqodcD877cUNtEZ
dEiqsyK5ySq9AvA+E0nOe541e+0YQX09w8tDO37DcUVFTw3ZRVysnRVEzd1vSwNg
jCvxK5VBxlfeSa2rXGos/1N06gGH4DS44MQDTMHhIT4sAcDppNV8eUd82q9Kr58e
p1li2XRjWpXZoMS9pRvSjVeca5QBcUjQFE43lU+TWE/VHzrucEOkM6NVCDKLba5Z
SHiuNfB1uCjnVVhNZQCHPt0VA8zyerFXqA5Vx72u0mAZFKzQxqM4lGmpBao9QzBu
gyjCst3E3rnzsHZ8/4azEm4q1XMkiFB5EGNjca5j83irCjrpTskYFFRvvcIIHCDF
1+6SNY+l2A4bsLdV7wrsr2S3qg3bWO/KG9llNGk+krZC7Dpnf2oPV04vJj/La6YK
mHkm87gdB3u3l9GkJ8gE2ntbOiI0Wx60hLrb1aE/e8R3kyhfZT/1gaEKXJo4ff/n
FCt5qSo5tUoEIpS4pKmeZ3Kezn67ni9R/YDx/k/qzA27rIgUMtPB4FPwR2V34ZeL
/MIgqrtJAlkO1HfiGvWt/ZifZLIU7XV6JPcJpiOHcwmmPzKvrifjk9wWhfb/8dy1
Y9jatp0wbAbK231YOjiyhTlKKNwr7Darlo+vrd+sKJOGCmL0Bc/xqUPjckbv+gpF
qeUxcO1/Xga6T6Ggvnyuvxs6S7WKF/LiJRO3FItcLQiwn8gfW3ZxMzMnZlNYk1pY
dlkBtCDCrlHsUBcPH2+/QAdQtTKApvkq+p44YZFNm8Ia+TuQDLZdbOZZi9iDQkDy
J5ie5DZrdxk/JcxEgSZAbuXxKVljry8gh6dZzlReuVTXzLOPiDf6ejr884KZYZeE
UjwM2/D5z4NY2vYs8wgJoXU08+LaMWdOUtQDbst9kNSRpiSNQYyNXzQwRTUcLYxa
EC2L4QKrLkIZIQocRSD5lcodz3sHf3jQ7NI28UJIu+NZkUdL+OckUOvqegpUgPVF
L+0of3E6A2Q74R251mK9HMoI6PE/jUXjH+w5Xbg08c3u8j1W3/maxZUmGPrPeEK8
7OiYuGKwnXBwxRWPsL8ErAIbsi4r27plf2GfIGuQJfjyVTU6VEgBvnipUprJYjyB
2YEPxVJqLE03m5OTo4UTy4sVNeKmBjUbIbcLCDIMIxdXgaU1hYlHIvjKfJs+UBwp
tJJ28kI4KjBa3SMd+6bHWc4rM8rm+JoDQJMOnXDKjGMw1xjI95w8mxcHERELtU6W
VIcRpUjfgCi8+1sbZBnZBqO5oZv7f6KeNNlLb4pBNY5fZgFzbQu78hi95LsGN9ux
Wo4KiqOFPpQaiOso0lSNCYwgCaX0+zBuopYq6Lqpn0Um+tA4qQfvGDggyBaFxJO9
BKlM5SRl777O2CS5h78CZvuwY7M+igZir5iG+QL1XfQVBBahob5RjQ2+4keoYEru
GsabJB9LZwBlCB4WB+zfjzfsKohCVDC33kRLJzQNPYdz9s4M2fZhzEwI+fGcx3Ev
gXNGJH21Y/2vRN9fyViar4mllioXCoFT5/BYCH2+phx2AOQn6u41FeygF//GvHn/
LD11vzAxHhmxi4JiXyDhZB5pzmcFZKm8y0IZRuuo6Mm1BgYm/bQlrGjdBa+YGY9d
6uqdCXAK1JBqZRr6yd59zdW6SqPyTKhPbmXyslFmSNpo/l8zaBC3k9/3FaiXceKT
dZ76K+X9r9LTIzpchvugINmSbN1EcMLk4JVor/67HyQDwDmy511ogGOfEuBdEXvl
YCXie9xTEPbhU2SCoUi1H7Fk1ZAYLcMs+vylY3kjrYUheLIZlXRmFatM9eAulAb3
Dm18uQRQEInWqFD0L23lfzyf8n2dPZ/tfjtRyXaiS8cAx37BnBG35IS7RypnA1T4
KalrMGMr8c8y3PVSob6wkalGmrStIj9cmPpWGnNrpIpqpbyq5ORe5Jk9rnwFebbm
0dtfgmwXMoQsiR9qWrd2CghsL0IiVvpT6C8Rbiry9LdTTdJFFGVS358TtU0eFqBT
/sCCDONWy9inSD4pFMJPgWHPij2eIFyJVqvcj60gvSMvmSv4EDJ2A3YG5awKhyLU
IUygB85uhidcc4c6dsAoVUSNmHLtZYIqJ0fHAGUrtU63TVDDQ1ZFq+elZv9ccEqX
MOJFIRzql7ZeqKMzY4hFZ1hPqkDIajLuGj6FuTZh2DxRoH7dkNcksKKOxoOgkFws
jnc85sPHBaS0qoWYiNq9x55vll5rtzWMxIBLks+tbdhQLbnPKfpG1D/Y7hJogH4W
gjFJn3JvcWHyJCR5jHJEEw7aJbjkp/PlW13PeZdDXUsnwVVFZxxR+bySm9we0YGf
gl+QPRGKXfPnjOFUOVVA4MT1X2r4WXbMGZ9DXnn7DDJBYOy6Uj5eAUxDuOo7vtYC
lY53PpOKU4/xkGrEeu3ZAc5kTWApiFR4J+O0tcqSzTByD5IRHRbxMdNAkwR7wlT/
e9cI5n4aUlfNOmNsPXCKCcEQdY2zJ1pbELtqUcN2+55taYnc6O1K/VQBqeEkwgAY
ZjJa/YzLnEIhdb7Bh5YU8W5LN8LgXXgCGKMOWnGmCybvd3Ei1fHzmqX0kfYy5Cb/
GVMAh2dBiFm1RuvP+PU6yk1mXhMcmgqRVpVgVLWWh3o+nfODUbMTo88lXwIKk7dM
U3dl7Mtepe+HtTd4m+GAl1xDJKxprIft4Co0/aV8S7s046mfpA1j4E0MzHLxgOqe
dcbHg23xr5DK0dwkd/M+L2bKw1IMf81JU53ws6acdLXP+WeupIq4PLfxcdTWefVj
5a+JvJVTmeeQPtzZZtHRhvzoiKMT+zr2DgxR9ZdPL5nM195hBnv5qWD50PZF5nUE
hcJxfSy71V84CoPfEu031FGGPxKHDsexas+0S68oRiXQwCxUDbJCRTlDLy2+Bd+C
oobWDVcBRcLcLurixy/iU+vepryqMRWByNGk3KjvVLSA37+qAZwI8R1lH6670cq7
ojU7Zjm5nLb++/YMQN4E4+4rfS8wVJxDXq/QTasqtiKRtkGT7sD1WvWHlu2Mw1+n
ICzSKyql6GHyR7SWbcbm6RYm9ednvNpwJ4Riw/CaHR04vhE9cim8H5tSvm+xrKun
s8MukNySuOd9HfkvhbhkrnBDq0m1Ku7xH4qxutI7ABN5boQhZUOwN4CAUHYkEtXc
tYZFNUA5m3DxfuUcFG0+llwF1zjJJQ4rpig2xYLvvvhvvRVZzcy0NthUKm2PBLPx
Sjwzcrnn5cnszGdu183NQDgC+XsDhvXNZFo/JSBqeM7SFiPlWhQ+qZcei2HnsXTy
EEo+IRGVaJYwxgTucepZ+A7kAlr0a2EGgfBTBz2PSOy4TO1NlOBQPMcaMuNfT7gw
Bpxubccvmp2J6FhSA+eq7FvGQ8HpWt2+mW2n5Gfk9RN3c801r9XppgXS2+HJr5bs
RlC8RQrbPIKXmwCgevYHJkw6ETuaf1oFvI8NugAXN14ivKt7sXCWNRRl4M0HJ8C2
oO8B+bNjEut0vBavsPK4wOxcWFyYiH7R6Q3KsLRrBdtT9bznt/jF44QILOw0zlWn
S7v059CvoJnZaK1sYAhEijXF4ol/gIcE9IHY4k+c/WY9Wu/PLQ5Pt06lnIG5/YLA
sAL0RmhHi3kF3w7+2++c95n0IjLLvNxgZO8DlcQadZcgzLi1GG4KKp+KcOHaqkkp
9hCJvdIWrGcP98anxs7ycV+ASTU+xMLZpbk7gGH9//IozkYiQs6DwcR656mjub7v
/CHzL5Ql1PHieOR24RHdOALGXQT+P7BknbRLZVf6pwOlkz0oqUO0jbmpmakUzq0N
apcU/+8xvsaf940G7t8yuWnVDbt799fiK87aXCCZxr4nEBPmD9JnvYuljBZrN7Ux
Szya/oAmWrvJvvjLDsec6GBNn3RCmFFgFWazQfDFn2f3uVm/uiM1ovGhG4B6ErMh
O2NFhzS+FaArzRnMdpSBfGFC+58hpQwuuQJ2/0oznlwjXAo3FURh6sNWNjkbfIDD
HRhVn7Zkgmx9QQBJdxXapCRF1dvlWKxW0Ubyj0oDia6f3CBVNAyqDEIvpwMfp6Id
U9NY+ZxSGZDELF5nX1lZnXbXsqTY36HYQFFMSH07HTjOzF/xHTuEMuQes1M1y12W
5hFwvWBPSn6RJF3KrnNuzgi72fZGbF3mRCnYabMPxzMO31tZopk6o3PZlXB0v5vF
XT1e8bSOS240S4uLIUCgiEUiMtLcCrysyqMnHfozj0qDBFWeXtLAKdwgkZs9/v9V
P2P0Z5RmXZXGPNtPYqED2+8cKVR0LW5Hya/LR3kmO4nCVAGPWwZ6sJYE+qdhGGzl
gX4hpY5OZQt/NjO4WpY8lJSoQUEMNajfYoqlxSQYx/sawTMq5g4UcbgC6QZD/pFK
s5JdegfUt6NPeB4wYVrFHBWRvjTF13XtoD+EMteMRAOGs6QR8B8haxPH+IGlwfr0
UIl1u20vNLWqWdiZ6C65Jj7iA3o87ulktlj2u8WwTJMr2iCmKwxR40IPVuOqwxr9
gwRQmcKrAx4aQp+CCW9eMasQjjGMD4rEuNzKQ1kxb0Zynsf87uKK63MIsxLIiIOd
cjgzperYmb8ceNB6Um/8XF2SbWmJlSezMTt10une9s2QX9blF+h4dcBYCTLkow0v
i0fq1W9Kfo8k9wNkGIAjHZ7fV26kkMoctA1ujBrGS7bEZ1yV6JXRrAVrHYINjEuZ
lWrf2C87mOixhcFtDsaPvCgeb3SmtxhcXDw9tjP7WgiMzrjXyaWjl03Lologinv1
nLU575ird3CQ6GHCQAl+OuFe1W+yXDDyZ2oREy8fXGwjXecUxsF9xnqvGK5PuZ34
SodsFxKaeRACT2ceUzbqthspZjFh6Rc0hao4H3WraYNxrE/AQ8zOFZZV1gdlD10/
cYj9j2L8pNEeIALHhweA6VLNzsK1MEIE0xuW5Bo6nGtJ4z4CkuSsQy90KQcj1vIS
gQ+CSgpMOeUdBKj91xEP2toKWtCJMEhaLHMxzBFVQmJmaG5lNsxmuF6+F9bF1to7
mUVRwOX2lK1BBhIEqkH682Ci+zMGiQuvBGMSizaOjNqO52vFsqw9mTkehDQorTbl
GDpIh+RQjyci/lje2Kno11ARqKXufCxrOvnfosSLlb6t0zfmmOYYYWGK6b8Fbedf
HadkHbgFDTKofUgp3rv+aF3s5/cJFj28cBUb9CfZJm8k6CROmFHm7zcQiHuZ8Aky
W6oqVzWavcqs/hF3XRvlIazxiuoVKP3sEOLhl3VRmmhRM3vW5TTE90gQrNjGhH08
MPx+4LCgrQfKQmZSfgAS2hHnJ9Dy8FpRV3WGGmc09j0EB/xjnbFsbLKpYpmW3OWu
90lf8NrnDiwuFdKu8nxHPCqmFqJoF15mF4KPaYu1eJzyTyVKWcaqVPSkCETFkaFy
gh8sA1GGAJ7qs76MiAqTqp2DZAyCchWENAqX/eOT1nuO6e5mDu0OMaG0PaOZ8l09
F4b5nkIY00TUKqcPMGxgecM5Rt8NWchDNEzK6yq2owlrovF+KvMhn/r6X7aRv5iu
Ubs10hFcHnBvyZyK2YvF4yc+Nq5uPzsaVsrtC1oGrnzazL7JJOD2OkoE0G7gXv/M
+qliXHd2+l1kehoR+BdMOAyJWdJxrm+AJgSc1ReHm4+M9Zno/dOsOSRK1LsfXMnC
APmSirvnBjuIyI8/a8v+BYtHeUGi1GcaS1zpsC0pG0QyUWNXKyGS4keXXAAO6Nly
i7l+Tl1wpBPw8heyGbrUgJCZdxWt7E4ECwgffw8lZsL2o71t1Qbc1ywbYP8Y8eXv
m5NYJiKjiKaJK/X6Sn2JDE4T/Ku8wQPfgHB11NkBLR5ysqHASLc0LTm4T+gNFKQt
p4Mbfr8vCUGG2dcumiHXr3nfYVWvb+49bYO9/l8uYYSSwV+EET0wkYILuhonAj9/
vkDEca24tMFpyYxa2EZ5BCPsHV47tZPr5rio1es0bLBsMTUpb0Vwzb4VybM0bUgV
gXVvPF7bQ310INb1dwsZ5XG2Y796bMxF2RaFBzpT+YN+B3hMYRkG/Dh20ByUq7VL
s5jz9M1omgWTBo+0AvrjJmvatzfs8hzqwW5nIiCdC/T2rqn5QuYWcI5dZUi/+8i2
al3xqsfZkP+snpDn9fEkhhpxDXX7oqWmChb0gnKH3RD1KpHZ69iz7vJ3WZyPcl4E
qS0bIPxhlJ/++fYnaKoK+/0dN2yizFAPYRXPJ88nEv5Ng8phCI++cEOunlWsHQhW
sLmRnW1zG7uvzR8AQ0AbT76eZqnSjj9QFv0c2KqEAatDRdLVt+0weTkksQAy5l0b
mrLnNiE9HO+yLOsCsU3Zl5A8wZAUSesU3yXIjRZ5gj+OkV4ly9Pq0N4jMmkK7xJI
+h2hUJxa+wFps9MLQQTXowrCPzyiiYGtyKTojKdvm0NJ15pKAWfsOGN15zrZ4W7O
xvkdG2O4pwUBiM61k6tFfV+4R7So5GKlrDI25Fj2Qs4nIw6H2SfCYPHXjwxQMphg
TlWXLNc47cUpw/DizuDagSrSwaBJic3xM+qj+s146SqLxgj7uL6UW5qFZ3oySAox
v28Pv5A3rra/eCTSQcknXUMeV8LehxMrtsHRKPCbLxo+kPOv0UEfYgMruFZakHLM
ulSUKDduC3v8u6BdKhlQ4xZ4OherGSj9oH+m8dFPjuhBLllwRtVJVY4ltzAZqZzW
y7ILymj+VljYDtzrQcyecrPg/AbeQmYSA8DMw3J4UBIIwwAio5uNskKKLE5orjVN
gUuLHhMWychHyPqG84V+kh7breMpO45hGNZWS/OUlKD3LZ5l6g3/waJAiPKEg8LF
YvHo6iaobdTzl8Sk+gbnyQIzwFIjKi59xmkLKx91IYTOqHmkMA7Mbb3QuWkT5FY2
LU14dr5hzG+31KjcUmuAbIQtE5p0CdXHExJ36Ir5nQKapwXO3Cd7BawdmOkgo5Mp
B+7KBZkpPuS1tvCt2+1uji5Zw1PxisJj5vQt0+2GlNq1gs9Xhtqkga5F3lQj5dMC
h+7OdEX9Ye2oC9YE27p8orTOfuARYxFpzHBXEQ7H0lEAa5Gok++GhPGOfA1E5jpI
3cZ34vph7+AmXTLyhRhG6IvEwl3eZGLzKgfXWoM+1tLQipDJTdT7oZaqa2QRKtrp
5qUsIhCSf8zzGUBbaZWU4srLa1lMJqKRmVg1OXl+KdIb3mTimic/cEGWDaB1ybmr
q4M08Cw2B2EuNYhTTOBsUYmN8es8LNliDaPcTPj/u5V2gaOj/ok9ySNiFILeNVBu
IkG23+la3yNJ45cXs9SyMd1tPrk5OoyD3Er1sWYnrmPktbSDhfdfS3GVMFlvrnNJ
dPYab2eJIkTnePdK8sxdz7Cx23NeWfhxXDURrz9yLlx1xIa33Mnq73n1/Wk0aKjV
PU6as8bSORNjN0epZry8ux+3YZV1rSeLHe+TWSpzRID9UgH9Ht6K6H7sctzYhHFD
DY4guAGFlA0IyViItpCO2EaHk76tmStmcuaplEazMnPkg5YPPgshE9XzXjTL9L71
NfGjzd/C/uEo31FMWSuXv/HtBT3OXgNqUQmSNb8O2epCfQ0T+Qy1rwx91W2uGmAV
kncCfp/PGyIWJzSIlo6M0ctWy/xQaD4vT/SSZjCy4yKrSLzTZlf4J/hbk6FE5iuf
Tr0w+fCp/wgUdgVz6A0RCqydAXfK96feqv99QcdF/a91JSASaid2v2O72lr/GhkM
Qy/Y5xdCJ7uPJkiW5+1d4Ebn2CcvwAnpHb8gYDvEW9qFrPNFbvWGeXgJw9BsF8wD
6Mm51e6Ny5xMCiUEfpd2NAW1JWf8KFN68c1rmYO0fqGrRX+agEddbnXGrD8eeNbx
MwTUMZoOEEwSOkJ1z1sbtVUZnfjKctGKLUIShtzys1aSGUSa6exiEBtJzEkkWKbY
432rL2HP2SNgQ/T3QJ+lkLmJfICaLKXw+QZWgsL1vXL0xq8pNr/F8y1Ogc7OGBdr
jHizear8S1j91WPFeWzYmONWkZZgUCM8LT/J0IabtX5D7uD/CcxMgsrq/gXuFB47
h4jmzN8WEaaKIEg56gynq9N/nEgaFoCM79MiugwZlv9e/tdtYPVV8IGDs5fDhHpD
xQxRqXkZ4PsgwdgwOqaQWbEC8Wyus++fGNkgzlW47WbCVBpJMA86Dn04+086Q9Tl
I+CtcC/V8J6WoZZbulEpqAzZqwmT7GNZ94qNBGf+BWpvgNSQOjy/9voAgsTagKU2
WyLsBvH+yt+Aqmy3vLxVJ2eluYlBIFJqyu8AiMZhH89T8N93WCuwIwKGKeD7XfjG
pMiHvxFcpyEu/64X2koxgEFD9tTd/xQlAtKIoYdA2kqlx8REhDLLRadV4/N3FGgs
U4B4l5fncuXeXQPcHMXy751JDbeJ4mhoeLLSRLhcsqZ5vEPphyG+WEtMbwfLxksm
REwymkj/PwUsduL9a6zqzFkS0ImO18KIA81qEFr0Ai84hjxEbSr8dOsaF1RhgPH1
4z6lX43o7UZMAlEg69PIrtAHmU0xR4yO0hYki8YtyyPOvpK/CIDnj60aPemqHlUf
vDTImETCzzH2PiPVPv12Gg23LTyjgB2qKhzwWsI0VosYCOcvrdSaCNQbosKGYQ1E
IHC3WUoXSNgYwxK/tx1YSYhv2kw+a7WKtTHm+dXP7XUp7qViO36uXIHyWivhVdJ4
qDZvOJqC8sw/6Xp3p0Vdzm1nh8Z0WFBzez/z5ebi3XmDDwbqaEzvrNtHbhrJuzrQ
l7m/YJl/PiTK5oIMX01VNAOS9qCET2qGVv7vy6ZE3Eja3YejUagfKVyBntBj+g/N
O5ME0UtKAJgXX5XcgyIzrAxWmc3yfT2iVAfRhLks/dOY2LApd1mHkvaKHEnDSAlN
tppq8RHxzADLcqkGalPuSzNvWmKyZ4JNyeRi2HllRskDVUf0Ic6EOM6kIJchwBWZ
I5hag6tFVBrfaqTQVBB7h+HsNBR3paiF3BPwvxdY57ZNE4lreqDfFxi+yz4DUyv6
uR6hij3865FpiXnxmMHopxiTLNjdNRks/7LG8VFlKg87y/7TEkMjaC9vOmIZMCGZ
bvVUuQd9eKNpa3BzBxAKXMkhDDhms5B4U3CB9vHV4q5Bq0nCPLaDEjDMkDtVtxbg
18FL9KJ3KER9qqHg2ofJcY0oVQvqDR8njZPZFWJnR1PcMxeD3ROMSzoigHFO+Ier
Tw62RNrfzMAgC8qOTJh8eMBpRt16GIjEzqJZaXyrBzetnQhMYwyPHGdvHZG3DcTc
hl+FZG5UZnO1gxdENeK5CZHel7lJh6uMTg3aJBgSx1fMebyZX+6bPdNloGpzRovN
5tN9R6PEU4Qhfb+8VVru5v6/edCn25xIBzzq1KHB8UdDd/uBTqfvrL+qDEluQAWg
18/j7ordCv7Klu0VC+gDkck4kwOBxDuspq2en8WiURJW/qOICUPHv74UcuhrJQ+i
ApVGtPE/lcvbCVHWXabX6JIYYQfkW9l+T40RK32EPWc3zzQFSWvnUZ05fqd0zKFx
8d1fNNCaH6Bj/rLYij19OrWGpRy/DkWmu+eDBlRVmzHP96fpsgVzH9mg5LoY8toe
MEny5JCoh1tvipxgpxBZvU882v02M/ftxJtQ+PF1LQ7s9BqCZPSHSFfyE2gzDezy
KtPAsPNEYvzy6j5o9nGLJfTCVGGzxqe8Ql0Nbak3F1l+8zaoz9wFJI7wlZneLksH
Cy6mQM9mXcRgujSYQQvDMz25cATfD0P3IUji+NxHSIHOf6iyUsP3MH1Yl9i6Vst5
5ayYvs6ybSiRPNg57ROBRXyS6aUnkToG8HGKEzGID0ciWpi4mytryWcF4DkSeXOB
SfJK59hBlN8VzTUpOJcGeOej7/jyRWDlAwmv+hyeaz27XAUk/dEFIfsFWm8PaswB
/fPHlIrKZvWkkFeIdjyyeLLJnuJGk5OYnfk6HhKr+S/YqL04PxTbHRKJcHWn2TdW
M2sz2/SuP3NSeOH/a893AhmNWdIn8gr/KY/wmZWjYzGd1FEPrmIc/UBGR3qJDFsb
YXCxRqKEuOwA6IeY1aBvzlkvgcHleJJ9E7mtR3LuFoR8ud+GakqcgaEfuBfSTO4v
5pP1WWbvJQ0HXFFm8WIT+ZbzC+pRu+YdneUfMxMI1z+nsG1KJsYyA3RQks1Amgma
Bjp85X7SAo5/Wimc+BQPt5veKo1AHDv0BmhUKcpEkS+kByuqmacGODjgu67rPZ15
EmKRpI4JKvduJt54ySAF6YYZBKWN+zNsSAaYnE41KPuJcNJx+ofVmedfIsafSyY7
m2Woou6RKi/eBHaRaWRaDapqka3ePS5+pvJDVmC6G33HkNWx3zv8bxrh5Ha+BQQP
cO8PYgynWQy7Q5MCz9tpzgsXZYuSB1GjzLVCU4TEWpeAsMd7foPUfusgMawJbCs+
gJ1qLAP9uwHEnepLKpfkA9pUrII3lSh7rr34nBrjkkZZ+NhtIq+8ozdGG/J8MCFC
OAoTc/T/fPsuBKWLLCUi2rSnqjILbiq7OmiMX8bHPoHDm3OdMV5pOjLLZhi94+6w
3L/KjCzx+WFgwV/WXspMDPNsL0rDkKjKyQERiOSSKf9hLDdjhl7zYLt457zCtoPV
ocMSNwgefK4lWAgpNmmtHpkPgpooTFb6Lr6TCSoNTrlYmdswuRnjgv47sxeVMNhD
OZqLH3L81dUhuGukHrsUsNGWHF6lGhuZSWWZIRaavMiq2eZi0byBVIeSWnLETCD0
Z5cPePxuSVN+KEZ++7g2ds8RJyZ9BV4y+xXfUs1C5k0LNTKpfaqRFeLGgJrXU2fr
3rOhpPB6DxpW/9lG1XebjNiIyEY26K6ohUNlBJkT7bPx8YVE/7fmoURglycd3xjx
dfYtDDjxQr+wg0Adgz3Vm4nHpCPtdXD7rBMpK62X49EHybrsxOZg8iAcJgxH5lvA
KFj2j3ngM9iOYThZDnoGGQDKa9C/dOkNXK6DCU9Ix4+SVjRjMWyzdIR7rHrAZb05
+pP+tEIU3rK2Gd22cVKOJefsb+FL20NhBNJs/3cSDmA68iAts7TqdSfFKi2TAXMi
6Xo/xg0koCOa77S6fUw3UfWcIa6nRosdOEl1UjH4MJmjAQ5jQ26CaJ0CA2AiIrfx
YaubNey1sy1dDFn3Z5ghuIXR4o1kxhkNcMEYwleVB3AQCh63j2/eqgmZEe/FSk1/
MX8C88CuFO0+ruEqwVUEbXv3t4yy1rvawEjVAJB8Sk8YslwkSueEF4d4cQHweFVi
bhlKv+Tw5TpU9KTYtt/orjZ792f16iOALiQeSWkDlEFeb0qT2yRA0YgEaJGE2vNj
Gmd+nhdJqr1iEyTRD5f7rKMZN8SFDJU5M8B1PDAQhZBizEaxx5Kpk4QrN0G+UVow
wggXITJ9dZcV6+qgSFZVeKKRQvjurOZCpxnr1x/2zenY2ukO3VxCJEuLYCTCKq9Y
OjTIHj9iAKtfGh3968Ud1mx/pyOTsUL2Nbif2ZZQVTklKBHuAibFSERbc0DHFnD4
mQsMyGMHq0+bDCfKm22y8AICEE9Bc72j4x+X/zTT4eqovU4hdIMotrLAUCF6/9Fg
LKeEVPE0AKGyxgqgorL6YCxqnTui0wbUK3fS7qPGRXu8iQheVnB0Y7PGpqXW9X9E
EBHdA4nOUWIYggCHTgLDESBNDaV/kO2waI1DuWb7X3JlOikGDIZO4o0gt9nwaKdP
zh/00KSFU9qQTTHbUlrZxdzMai+HkUbdZccD5gDTGx70eI/n9LDwdmfz212Lslwb
O8oFDjPNXpytU4NI6WCU+02HJ7DsDHQDSt4sZFHf1I9EhhW7PvGStN7FIguc/Ess
YlzNnV01Edz+8+wgKRD2QfrTURUM5ot4znAXvArbKuDBsDULw7y6I+qnOJnG3SI/
9WOQLJB4/0ng31uXjVdhHsFkYvsDP4FLNQB+5xDBuydNryRuYCtc65gF+q0hYrwm
9GquDQ/PAXEuoXBZXK1nmRjm4lfmCVTEHfAE8uU+p4cxWBf01sg59M1P4ycuhyEJ
5jbLKsbFJd1qUvld0wtAFvxXAVt/8HYLk2BUpLz0BCMAHlOyWlOSJ7pPWAqFxkQe
pA66drESu8cX9RFJHfU+EeBtCA32WPGNK9b6Ja05uZwdfA80XHs39e1Vpef+/gew
G/ntg1qeXoJLkbYT9dXPLIMfWhpyfxo98qHmLKj/nnOHGcm2s+GmxgnSscEivFVq
ipAmvT5mUw8D0I+Xjhz9OPYc/SxbRpkwGOQpueLsk9veO6s/S6z3csskY3Q+iVhK
/QMx9MZonzqoWTGZrS3qyOM/Ind1gA5ub/B3Ftfni2qZyAKI52NzQVrvzPiD7yLH
94Di80e3iU43bEp6FwKVjCxj89CRYPy+CnpPphb3+f2wp6JIKc9AF2qR8bQVy6Cn
jYG4xyDu1QCXS2bvlRrnOFxbwqKMtEyJpP6JLRSfYVvbnk2VPuni5qFcfgva5XoJ
5uAHtMW9vt6UZPhUKw8fSJYudxpB7RfFNvdrvG7VJ1MjoEGxNC1/RlBGJbmlPLrO
BaXIU5xoE7Ppu6sXxSgvNs0eW0ck/F4405iRTFVFCUYjiXM/Yk8KFqH5zRHNdANO
hVjsahunuQ1U8er5AvIWaV86bKMR43ebEgKKB9z0R0t7IaFynHzJ0eHXM/puhB5M
5gw0GUnY6MAHhbg82d/BtJWdx3W4x1Dm+MffP4nZzceceXGAw4C1HM5wwdEb7NHR
WjL1m1UZeBh0wcAa8GAdVX12FwGbDUVihPqLCEmvOy9VojFkpp1x8YjPVpZVDxp2
8Ip2wlsoH+HtufqTF8x1M5uiUFEBdBe1kWOkb6fFIzmsZXP4uV/PQEE8wocXU3O4
3QyUEyxugpayTWYbVy515VgKsE7E3qha9rhfaVeB4IwgohY/iOE/3byqb5cC8ktJ
vlyrODUo97fBeQhBua0UnaBdLsTPBP2rFUn4e8tak8d9iTied3C61XnazzSSFNxi
3lspt51foZu3BstZZSAXICCd6TNgbn/XBwVv3e/XhM7FxTsX2JxHj7GMTz8PfvEe
ftW0ZuuKPwH+3grcbGtjVrqMqjnpmIaQQJtZsrZ6coUUrpiGaa5d4pBk+C+xJKLO
m2mWX7niH4hiDYFcLCVOqaN/QlPj1TUuczhQYIb2PwYxMP3Q9Q2EGg0ZbRJPx++W
2t0EQaVNvfGjQNt0HTP2VYDhmLshBKexYrXby3vRuSFji9zVYJHH9l1/8lKmsh/t
ESWOlnEOyLQe9NcIIUncl43bMkythY3PQqM3BaLkp1LINMN5xrM95RqSjiCyKDRg
nEzk42qIkie2nwp3za90liGIcQxYAtCIteLnNs23Au2HyC8UPYCgFuibIBVYpuCn
BWyLdO55u6vMxl5wa6qLDqisPgquhzZHkvcAJ2flmTNHBvVMXrmwgYQE7mpkB895
rj2ceSq5QFGDq8/S8wpN/ZIauj7catkuO+aYkLnuti0+RTMYUt/tCBDVicynLwu5
URthemChmfwnhfFSwUDhn7jJm1QO5/+cH5in+v6B5ue5Jw+jBEkOIuR4c2Pxr5xe
yelv1/Pmyx8z1O+/bChsNlZ56W+DxmzyqhppE9mq4a7+1eByVN57PzguI/ZNwt2e
Lu2OALsvuEcei5lb9pHfWz3UOk0mhj5oTJ1Rk8MycXTSxDSrl+eiNuZmObC0wP6Q
zIC/lVT2w/ftYUFwQk6JkXXD9KCJFRJxz2INSx8rZKYfXNFxOZb9SAnA4xYGbnY5
HXFMUHtIW4NG6csIequJQzPhW7YIY+xKDxMdyDKGs7JX+mFfhNanTQLhUqgbro/I
fGaV0KRbUxWO2DDBMdu8xEDGQT4FI/aOr7jJ7xfv8yd3zTOFhuyEhu+YaMbjOy5d
wxOS+J+QFfIbc69ySsSDfIsyCXlnWXVd5t5cSQnXqNmppGhuWlarzEPHHWOXjjg6
nJ5h2ViS1/pm7IMtb0E+5rWmUqdewYnhJv4RtyAdw/TzykuIjkLZ3yPSaMDuple0
S2+EZXELoKTffqd3AvnmgeW7wBDmwY0TD7j/2mZrau/6VIZUF+Ck/kexjsYBW6Ah
6xSrYpcjl3BZbie/Id0qUEO3SLcr/2tpWq8wDMVtBTmihD3RzHZHXsNXjyZmWMUJ
N/w0MrXCZBGJmej2D1bc86C3oeQP8U6A7kINsEI3kQsjhdmUDiEc6birpXrjorer
RpbfdAXDiJao1TgJBJkH2p/nJe6d9DlLx6RnG67gO7ap8tljdkB+qiSh60OAslw5
byB9oHtOx+ZC1OrQN/Rj2TGWOPiMws1F04RLY5nT/uOxs5pTFh41lmYsVz2prQxu
5hGO5pcr2ALaLpMSXz52IPkvaWEr4MFMORFxboIwUx/8Rn9jUDLcZp44Bo9Z1Eul
FPXXwty9Kn6RXwsOBGc06zMLMHjJT32q+NXZ1ZjMUE44jqTTyeDQpK4nVkxIKsO7
PuQB2KNFoQA4U1/SqYKLogBZrThmcqoydLcA963zeyYc1bo9y9m015VZjbH7n3fM
tsgQYFEEBQCE4fUXWgICAOUQG8W7Q8pUEJeSUcrMaF659bKfp7cc+4GeYqZ3VEzD
AlH/CvuV92P9dnGj8zdqnX8RaTA05g8ULIF8RIvkfUiO7HS+ei7LU0yd5obnk5+v
xsdfGnlUGIXH21SBZwNU71UhUeIWD40wD+gkk6aFPg3Jfd/E02+D8nkj9X0s3AsL
9jWKAs7f1kQbe58DEpLti15iyR0iJ52xpFokrH52X3Co6SsAURkSYREL4DlE0fUV
9Z5x1DTMQ9KLaJDOhWqlO765V1dDrGbHdHVQsXqO+O9IP5PGhfLk+hwdKBfeELle
6qIH6Q17lcdKSTToMbui3GcWV3K955+bnc5cDoGaE8+RG/oaq84+MFaMhyd53mwS
l6XPfwEIBFHlAo1D2sbxkCnIvb9tiYLzN2oIhwQO4dKPlHz+IcE4igXwicdPXaO0
bHCxO9JGd3KEMLxI4GvBKhNYlkk7sIzEJlFfV+HFHaeBSSXE56zyeczriu0DMErP
yN/ZBI7HjbYRdFpVYlbr2pCuWiNCCFSemeEaYjRS6Nw+t7u+9HTfw/EhtRUXWE0J
RMSeBBrZpuQ2GS/43nBcfwWw0q7BqFuzjLquW4jIYvYIH/CtsSvE+OTdJOO/pwKt
NSb27EEp4AVPyRc+qz+WJvY1WJ+gGIHKATJ5B75mQzIwgwmhYav7GgEruUCY5VUJ
ewceEg6Zb121dX6myZ1Kb7M+yFfVT1iNGe+2uip9Kf7A/ByemrqZYLZ+ShS5vAtw
6sQvP/4F2Jb4B44xAQhGbHbSGT85G/BOPXk4FjG74LA0iCorLd72VtN0h9FK2Jbh
rP8MGSO6NwMoszkeVi24APDNsp9LjEFnzfIKcUrMXBPcK22E27j+HG0keZoGcpnO
UK3E311oJruUXQ3zLwRjbseHlF0rntSYZ4sgdNFrJsN6ZIMOQvCbjX00471hRPIq
I0rQQ0ZNgtYWKKcZOTWIEIKvyINLOVMAIOXrzwcRuXgioN/x5OSxxmjN2Q7Cinla
J0FIvWhE+BBp+ToSD7hBhP3G3CaAgjk8KfiRAkNtFckD/hs+l4fqC1JRvSm0AXkd
buDtRNKC8yUzwEuxG/J9DdcNGyuZ2fLnFFrjw1CUXiGGoapnofWWCuTCAtAmhsUX
LUmBqIV1uxPSgW4hXJzrHfOXayUGNHoVdABcxJ1+nHdmtTHi0XMO0SUEGEtwqEAV
0kGdowbtIZXvceNVaNI1qbf5g3wutCEl2zKN+r2A84/qHg3PI3kfE23wotkPK1Mu
RthNXvHz/gQp5KikUAlkxj6fq+9yeBGC+L1efawWO1DHiQaUOGrHnKJyrC1Np1a9
v8B1LNuz/WXP8/nwYLPYrN+bmKQZbg4CHGxE3BYz4FTgnfDZPJOaqMgupFfC/A0j
HBGq2YH3ZR6rxvE+OLgJh5HA3PLYl2qoCGCFgNKHAfGy1apUe20TJ76nnC7+i0s/
HuSjzlOEJ1fnGA3hBDg0x/kNGqXEwLNe5x9eI/uxbVnSx/xh7Wm1TX8zprFN+cIa
jyx79JKt15FKtEFr+qiNlw7b5vIncw85sAlJp3s/YJ+HasRDGh6wS0fl2eRQYooh
m5A8LErdA3AbBqD6v4QgbXKPA+3UeQ9NzljsW/48by+3+al+ySk1QLN0RL4cg1Q2
NRBA/cRYijsDZu8Ul1kgMN1pdx78CAdxOUS+krH7bOVUQqQc0Lb61hM8WaF3O/tM
7aERuRO9SLz0gd3FZYz5isfZomLNMwkSCrBuECokL0yJovE3ig1K20lJ4QABYDq1
PO9LozVfOLHBVGwVJfBTBXO/XM8jRZcoHjnloejJsyAxXPq8ymzJTmBGEEQiaEeT
APF2JXSBIFVv00c3mW/FBiycY8sXtYk7yXF3Jj5nhApn6k7xovdvTtjOe2pKcc33
zu/4GzMB3cR6kbMwhXnTQ0I0A6Z85Kpwv79sVzqt4cXhdyKNY2rID5pmzN5fwqgA
PLh/stMpPH5Av3iyK7vrWmKV549gLntjVWrt6iu2eTzDxEWEPuOq0Hj/rdpJl2Uz
E4RpCPcDVNXsg3gVvCq3kt/XENBpQ4OT+2gNcgKYV5j6roU5zefZp+lxUn1+3YY8
dOAeqCu42NzHp/t2wU3QkbgA4N0oUjXQEzMIOjc19FOq+6udEUZi3wZ5jtoCR2c2
oxdtki2IpWvX1rH9RN4/q5NAEBwlcVwP2Zbnx4rZ1sVLy/Ck9LSV7qn2dMENBZtl
PVhMDKBj6IJc5+MgIRSZkvlE8Ry9hbmEpQUwLs60XaEQ1XHPpMhyF1uQhZYRJFos
T9fcOBYHEMgqEdgZOFhw0B8LMgQNBVyA6mNIeg8zwUOx7ea4fITTFOvW0HEVoz2E
XnC7eZIyweO0ElLUdNOOS4IFdgfv+69AL3AsGSRmy67InFJUivY4bpKvs/MkVB+g
IM2WQLorf028DCSzZFKm9oe6Ve3QrZ85ZHjur/7RkS+sgLmf3Ec7/psPdqNw3Zk2
vG7c7imcdkV5gZsWWfNke3WnlyH7cu2gcSrZJUmoxkdFsKIY8qsvyJAasA5KubgI
NMEUDni9FwSk+uQAlgX2D4ZtG7+JHW9oWEKkQfAZsB8m5HFt32oMtYPcS8qXg36z
GWEwWM2QJlsBwhTHTEaPKjCLYhh0UtVKVwV1YEzy/0HU+CM7A7VioxZaEBKuYL+9
rgBJLaAmRjXmB/zsHi+M5LgKx06CSuz24SjVGge5WLTmUgMBbc33TqQ2Ys4s41hm
B1Ex+oVHoy2t6VNw6MAmNUW0suciFojYo9KvjDJtENVaDEzTjcMlPdxG0z2gS5BK
MQ1xRypU9klgkypiIbw0o6dqwgL5vZuurEDYkl2SCzdz83Zk0QdDyvRxdLxxvORa
lv7Y7xcJKTTDl0BZGSmu1nW1TRbSSbvWjkmN2LG5vezhklFr2EGAs2ra4HIZiwun
QWHLcyUCHoer9GXVh9lT7WV0bZ2UCQLWhuRWwEElotng/G+Elv61L+P+0hdWKnkQ
pMbfBGf5Ei8oWT3iOLaVxnB3vCFcRctM4lz4VA53A0mIhkKh4lSDbzz351cLQQkg
mt0jNQYS83HIAFVRNFT+7uHUOSLJ4BBd+2NYkdwJTUA8bG1DPFvpD1KZ3q77Uy9V
Y5i0eUsd3+u5xT7evTO5bou4WR4tqXIG+RCvS+B/lHp15EN7bUEZ9cOJYn+JVgni
AwxHSw+L8Qc7BurYKKSdY/WTK7b6P4jytbnIL3ZbQbGUqJG/hNRWwkahOj3vmojB
Rq04zrqDGj586xzDO9g9m+7J5wO5H0Nb3xG/odTVifM9q8Gvspmonvvc13sfWKlb
4pMDgR/2uS4H1IzdxUVkB4DcW/CBpV7VUbPTYIkyalzSvfWRrNpwO8W1lPRqAeRq
7cGmQ+QSO2eNzxG0yIVcSi/g1ClkHG9zCbgRZpUpTmDAsRhwIk3r5ooCFKokJ1Vl
0HhVEfmahf2RVwnOH5QZLoLqeToyhWFuvTIkpKeh9f4TS+mhkalWLedKSDglf7Cy
FAExe+aO+MqBmw1kfTQtgmJMyQgs0BaojefoJdsA14tUvbAT+qGS8AAmpNgm5Yl5
cwvjGszVtzYk4x3IKc8rO1xfVqvah/odTh4QmQILXDKVrEuHLzsdgsUolMxv/iL6
AIoTfA8u10Dc5PS5Jb+xBPRB1rBCPkHyehlwgnWg9OiYqlc6t1/QFsL7yrOMkNc9
rPPnK0nKnzPxmiu5AK6Dx55hR0dM1qOOb5ogxE1Il5OmVYKNtdid2kdRwUpTB5pA
KbY1A9+sS9iUaMEk/umkZW+RE14XwYwYQTvWCaDZeTCVeUxhy3JtRJCstYCwgHn7
oaJRn+UJlL1eLUtFJ22yAdR/XRm0VayWcoblgEaLqRWih3LQNsub2UBPOHeg3meq
L1iunQFgnKV+TDJqgU8p/5iSMoXjXRVMigKbWwMSeOdA6xyz9Gb8S85tQBc9kBMG
xKngPzml7G869pPCC8PmmF+izhjKILXq83jUbHzrn2xu9rOiVyYdWJQQrmxi7BsV
JGPwT8ZE2dAn0/pRd5qsWz6I4kN/g2ysE5I0T7qp7JKvyauXS9T8M3cjaiF9A5kt
EcxKuGDbkOdp1QG+Eu6RghcABO0KcQES8XEP/BS//0QLYNVHvWKfw7Y7tlrTFbF6
ycyTKOe68oqqdEaSZUAoc39WRqD0JztBaf3f+9U89cpmbkAzpUTdiuVNdoLWdgDw
Kawb57vl51N1rY3mG+VGf1T8i9Nnyvs8obZn3gYdm5DdYhzrqe/7ESIFI/xVOFDX
FI+v/LB6SBn6/A4FvGtGWWFWXL2gTl92VKy8yQ2IPwmTFVRdIE4424ppM7XkfLvM
L08XxDm5lvXdwOJA+eJRYk78dVZhNdi5plwlLZ9VyUSs6MWnv6koPq4LMyxIGp/X
AGzApp7xDn71mT5ZWMGEZ0UDtJ5YpoTW7DeHPi5DJkuuJ20tvSVlqVApBmg8klrp
S2x98M5+MdL1UiPmBwt/gHtZk06quWAxJ8tmL4kSF4VaW4dGdAEyrtKMVcMkTRpY
AxDGdMm2eCTC2LHh8SALR6WXb6idxvLfyTEJ3fuT/IU3Rl0cZTOoML0VYOOc1UwW
Y0Kq0GH2IG8DAeX6WL8scIsh5INFlsToopuvU7F2oNF0koM7yT/QkwW31XU2YMoI
2viPqFsIfvDMJ9pTb4Cxkg0VCGmGdS5hVPAFAwnxYGzuNNoPJhZdPpbCLCsXEKC4
Pa3ezgFp93BHGTSzKTGnj9GdkaPdgOMyshBRwSbNfIc2v9S8Pa6S27cJi59c5Y+Z
L/GcXhIeBiyCukhZjizWPiKDCG/0BCjD5XJXzVDOPyoR8tvRnom9eKFUkjvdO3Ou
+W1/Z+pt4jcOh8WtflcFZbM1W/DR+BrGYs8E4C/znZwuYSQQ+//K2fL6nV8MUbws
7LOGs8pibuGqw+EB8HOg4x1M1Q+wiA7mFp7Gswe8HlmQwXrgnjtuK0FKlIIGXBro
Dvx9qYbyL3cvAf1m0OjZNOg0yH9UA3YssEfuEqYEnxn+nxYKpC/0wlww3F4lG/9O
1+0v3N2OABavgCDqa0jSWWsFwzRUAw2TZteOCmMSz5G7SyjYmQ5zz7++0gQsqS0J
IemyNMzK4BhTqnlQEnkKz9Pan+IH42BWoETL0MO5enhM3V67AMwW/cfg50NklOb0
Sz9Nx6XmYfApKP/a86aXaEhI4ckk8Agw7AIopogzzQL31opQl5eEKGsxzXBjqUS5
lc20B/2LWFmT53SAvod1Exd1C0AapPA5YITkyZX4ZSguitqAfRdcnZfVSkMG/Ctj
ci9KWlGuU4kBbYwn5BgI4QD24RI1trHe0jn0LhY89gtsmo9PElibcLN3QBIuxkjg
ZzHEFrj/ebWywIG4KVPGRI7LNdUAVELUf6BufUoBy8/k3pIi4aLFe0Y0RlhMdbHQ
6famFCRSPCmcy0SxQ6Q8u0n/jTZvIVOJ1at/2es2TDww/EQODBH5t0p+r9dr6U7R
SLza2P6Vec/qccNVGinuAsUoRuxO+LIQq7SIa2s/pjaAAk45Kd38kJWFgBVHhKu4
OfMVEfuL1b2Ty9cPeVfMGHmmpzNh5/gwXDM3J9a6LeBQJh4K0JPoiIwsxC7EQ7MW
lyZ1GumPUBIx53KsD9gf/ESrcQG9p2Xgrg5qbr0pTukZ4xzTG6Tzwt21wzHnLXf9
gOlILqkqND1FJCf5HFIiKTzXq8tBfjMesdfl9Lb6fhnd1o6hdRY9jzI8ICuLSgxC
mXvQ2ZiaKPtwYiXSwEqDQdFcmNdMsjHamaaD8fkGdXTDFn2QTjwQgaRPjJzRYTB6
7sxvpgMXnmJfTfvVXNv2g7bnv1PSgRfLBY5jXpz7iXDd+aXmr0hhzkL15UaKqLnw
gUUyUD5sYSe9mkK91d19eC55n5kNNc7q8dr+tFBwwbilKh+uG0EewshaWg1bYgAW
b8lyon81MwzsK+QxTCYQcRYJH/hok36AaPZBp/VC0Y6abarn0oaX24uxnkqyASqv
6AhhHZ+fwLTpiUFHgVDEqndKO348AyVsggTpNR/JI2raOyoCp79zwkteh2ZslEaB
Vnxi6brszENIi2Yl97JivmrkiV9LpLXBULn1Tb1h/hBr4/sZ4IXzsXri+ETG6PLQ
5Xiin9CHCkJsTAZ+RTSIv3YcDPie8XeoGmk+B4dcAXMMNmJTRV986mz6YpR4HAJ4
oAFO1kng+7qrF5JkUpHJqITyhh2wZrfT3VFYDB+h05OEsDjJmJEiyowHDQMrZHYu
zLzB1SoAayA/xy3Iv0s5rJdl/lblu1vxxGgP69xxj5Ht9lzw0Fipy/1i0kmFU+/b
zHzwKZvZH3IcOERbWuTbFuBtnMtiiiKWRhkGAPqxwgFKcRUDrM/ikMlekFu7BmzE
fYzxGPxnVmDN4/S+weFFdIHwDXnxVDq+v7xiXuJMLkPuemeXvGrMu/JM/m5tH/vv
jaod9yzs3tycignLWt9PwRv/0yNKTnJDB32p3iUvneCl1SML1OHitZq8bltJphB5
2WQSMm1+Qfu8s3pTf8jOZEFiW6zPxBUjckETREJhhYzhcy3/zZ9WXGdWxBejpz3g
VgVqqrmyBCocKCzBTBYrsZqkeEzjRLLmtjvfHdLB8AiCrryzVK31G/jTB7Aw6iSJ
mWmHtWZLwLMpIwxzhFFeUbiWzTHh4TAN5TrIrdQJwE8Fzuj3lmlCRXBRQQDtIcaT
TwYf0bjTT9Od0qQFLe3h++e0isXPwhjwOeRJYAGFsXn+0IU/qpbSq/jTeB/XHWqD
aoW/3P+iqz6GnIXwY/bevjiGd8YjzYjEx08ev9zPI1yRXfUkg+6i9RYMo59w0A2p
SQXgspv6XBk6h9KWbTja3dCdjl/TGozJxCXAs1Xc9oVt/Hr/KHsirurmgf9b8mGV
n4c2x0ApBWWxYWMn3NZOIL92TJ9g6ITghBmZ027C7fohpDDg7JCFl/V//XsLwTuA
U0Vvkzupkh+f+1zpEbC+Sjxaik0rqq8O0WBFGC91V9hzn8pSeUloP/NXEL98kmWs
93edM0V2EL2/3rt3/qOqjUBJLcl54FpxSzo9M1dYkZYKw5fnkTuBpSi4VwT79+xb
5HRmwupL2c2LgARrz97djvXd0ktXL5qk3Gmj/zzaRauc5PN4NZIb0jGTPKeaKduN
cM4MBsLVVgNI8nyqPU8Q/TqvArWblq/o7JpDM3huhMEaZn2F2bKbGHn8MhE0zEkU
9EPuELEhCXv99tn5P7RAsCv19wdjsy24+Ujqe10wAlj2Vtg1EuJGqX0TfDIWateH
TOdIurpSWP3JVH5Z1Hk4Um3MssJQco3daLUoDMOXDQfnhr8osFfN7nwpvHShDKHE
vtLhqOcT0D0I7R6+JQ/0Du7jT49XwBd8yEKM5qnb7okqfje8AyiOh7U1j8Ry6HpK
0EXoWHhnbh2re7Tkbn6VVIfDQ6YJkCw1jB17ER6Q3yqEPABZElfFzbnviLytvo5L
0/1XAnA3hU6oeyHpf0vlLCo6yxEFvsGxM2YSYoREzD3sgUSMwkK08OrK3r5mfGqK
5PkvFdibNF4ucLubeT47k35tRElEcW/vOWWUqMY4oT9lNxYAguN6VLyB4HIh/o8L
dPuJkDSVrShxBmRez+6jJeY2z4nOSjiXKTkBPnW7McXjrLMg4ClinKfVhzZX2JBy
COghSUqnHaQk7pgetSPHFCnwuHgpHHVUz7WfXvrMsLMeBxHwqUdlWoLIsIwQ/W7w
TGR7QXSCE4lBrTzeLpRhq1JqFHXLj+9fWog+hRd9ZzQ9OYYUCBUiuBn1Ar3RA9/x
mT9kHtNqsnMhxQuD7i8Kvd4Sj4tjDdV1eJNkQY4gq1TaVT92Shbz6z9ryVC+aVMc
m4eyi9qyfEHkqjyufPn7fGXXOa8clh9Ar4IEYoY7nlCAeEr1uN0Ks9jh5PARKpDO
1vdildyPVR+XcNyW7m4NKwUrDc+5r96ZWyjgIIhjZhG80mF2HXMel2MMw9bmC48b
fQyXNeDdb6I8ey3DnKs+Rlb0SryoxlifFB3mFbs60GeTswdhlDxj8ecVqGjlWCfT
yI/v2JER5Nv1O5OkC/ci2y9mlcfGD0RnEWQH2+ekda3iJ1EC1e10/LUR+f43aAA5
r1NYBr/LBlOwzqtR9XeZlkWksmnJXkTyQaQW6PSWYNlbL2RHqQ0Q9Z/CydVSSU5z
j2AnZu83QcTc0nRuFlhp/RxJNhXphJO7F7wUZ+uVHLegFn0l3jEHtgToho2IvMh7
7yxLuFspYXVnNYRdV8TQ1puQCFL4ECrv/PVYoABz/8p47QWGF/aYtN9+u4o1kU/u
9Ew4sA9eaaK7bjLCpeiPrV5OGTmv9PkICU+HnkD8eY+e5TamF45D8/n1uoVbjrft
W9r5cc2z4YoDfgGv0NwFPcOQAzSEBWVOeWX9Hl+gLNEb0emF0kaMCBr4q2+x1zT0
Xz0IF7JQBWiv8iVNXhSp7En1OYtOOQ9WDsnJHAbFp+CsqisKOlAucMpHvNTB4xTL
R4kVeRgUq5qJjJQjpxf8jSl5VGmzUMXVsqfsFND97DYrRXftA52i2CBZs32z1Vbb
K2qx4abTKV1fG6WwIjjMwBa5apCSGsu9Ct76Q6V8ZXBoI9CS5M5SwHZB6WUpg/ZW
n3Rq/eDxAOA4CBvgtGHSMkxMQrT+AvXN5XXAp59UBFlBOqeGLNMbliyhqpn2IhJC
iGJKOhwnBRzB/n/FK07bSiu235jbAB01nrbL4dvsK7S058z3TAIVzCCLQ3h2khNG
DP5n3aFPKgkRWWAvMSjqLXtgKL6mnXNTzuW/ULyvKIvaNQNjRTdNAqr9qJ6NaU6b
q5F0Cbt1+vWy7q/uV0iu9RxI0JkhFemCDDoGO9vKX90Ryvv771KdOCRt040z75k4
bK+AyeWevuGZ63R2aW5LlEagkfX+UhMGHyabrWva7OPSAAqQynSpcJC7ywAQtaRo
qiLRxo7QGO/hbCDoMbwzrjWN6bqQCFELrVY5Mejr6iOpfPIFDGc4E98/G+Ld+xmI
NM1weoDJqZKVrV4gyJ7Hcs2WJXw6uJMMKfOX5eOF48Xfu+W6vG1G9bqp8o3ExWs0
sGxHbFXXsQD+l/KSHVowiU6ZNHTKmKYE2rYAw3jfmfR5s9cdSc6Ik6iRpV7aw1xC
+VGonQWie9HiD/y058TmPoVeI8P7D8OJSEZh4o7GpbgOCM/PbrN3WFHVxGYlWVh6
EeelgexkLCvu4i2GY0i6Uh4hYhIm7JZnxDhf7T13X7It4Q0dEZFO7h6KlNQoM26M
yoIohN9i6shV6FSoekoIk7rdMk557bomHpann1JdwCQBYzknaCLoq2yb3z3NKz1o
u3/k+BSUTUz8IEYJ5bTO7dXv/EVPz8rNgRbwxYNB+zkSQTQtEpRwuNjlU9QIyf71
CAS9bLmXQ73NvRQs/BW3vM8PiQtNN5M5YaD7ayD3fvyEDSX+cl0m49+AalAEDzNY
NqTsmbCfwAr5LJ/uY2s+Lgk8AEHcjEWwtHZBkJjmncOnBP6x3t6JmHT7wC+UxvvZ
VLBhn2hzS7C3+k+XVw5WvF8JJvYzV6p4gOxPbFBzMwFn1IejFsE+pH7VYKHXkFRF
jcQ15VKpf37DqJYFrWixUJacQm7qcZNlSzL+ltz71m51B2bz/h2b5LHu/elnHXPz
+G5EqW5b7ovgZUjPWdX2Ch4Yfnx8mB47BfLsELt0nLqHijNLNZaFNyO1jH+SIxSw
s9BWvFvqbO14+khBeNmcG8hB83g0lRQiEB6zhEfRHuY/eQYc1v9Z9Rt84F7gIN4r
GmZFsddjng8cg3dBqeNGP3ovU1Kenu+qRRT/rcutl3GJJtO4+FgGGoGU3qEJNKvX
bKErP1qEURRzUCir3f4gVUU6Sl5kL6Orgo0ya22wEViMdfdCy5CcEgU4uxoUZzHF
B6GU0OwIh4CzXH6+BTxp+Vql3K2mT37RFhEsCrxIA5dF0NXHatOcFl8nDqPECxSF
8d2lJoO4ZE46vjRoCxgmKA0gVyBzf7uoiLo3BY/gqTWycoiOg74tuZTBdXnlKl60
dOaqH9YHgYBRNLSq73hOUc0KM+V8vOMAMS0h9qRuc5oh0PXYCE/7NlYBmexfFz0y
UaWNTbMwKMbcUAiwNigd/xka5ZhKMgZlVFE07Pa9kPYNCLaxpOz1wVNGKoH/orha
BkyOLY0c41gvxNuaG7aCYbZLt5NHHLPcGkGmAL5zRcjo+OwnO3RqOnODAw/cbPF9
sDARUiICnAe5HkLX3SlNlg29QloeO443nzPD1MJ5yyldlNZ1yDUOW/8X9N0Howsk
NVEMNiiHmIzKTqXfyOKACzu234znWYg6aFxjfu4nfd7/PYmxKHbeGqyV5fyN4JxO
fWM6kdOD2PWDbwl+3paxLnRk/tDDH71/LAy0CZIIwl64fzP7WxrxqMmJU0okxOGY
aa/FJaOBzALB1umAXm16jyFpaUvz6DN8+lMi7URLMdOYBZBOq11/UJc4x702Ts0H
1HJN8GX79Fe7JhC313DrD360/Stxk1RyhG9MRsZ68YR5Enfg7xYm3MmjDj+s1DhD
fG1uwLqf7FqMpW3zZamDj7ioPATBycXl3bkYkk0rVM80eMk+pnVqUHz/DoHbLhTM
hYcuZ3xlUzO5MVfGugEb18dE2ibsQtoqo4I/S9USKkXKwZpz6ZWlAn6T3K6W4k+b
HOz8K7U9ETkkmx6K5h+5EPhEABXu+vSBOkJmk7q7DhMUs3o8duNvlWUCS4E13bJS
CaoMMKNJmSCDswVXpKIKbjUOqMQhYx0Uf01zvHwteoqSx6FK3xJn/CbCt5Hz8HBG
/l2uoBKSYmSeHkI++x5zzUuJh6x1QKfPu5s/FaN9Rgk8TsQDONxwoLwlaHxGQIRV
93v89JFVeJ6hnhrgI/imMS+4ODAbljGUHrZDLgY4HNBJIocRNG9l1TOOtAz4pDON
5y3CmEpnwgXR0g3CoVXo/KQNjL2mZtWsou35ooXIpskvwmfVOde4Xx57Jy/iM4GO
OKVNIPNL+yG74Ofg38c/zDoHRin141ZMhAWiSH3ZMACuqczjNBeqEY6gLEFUhusZ
nnt4DZv26oA2ISTS16gwsbdhqNDS7fmIesSnN/LTp8HYM+Jt1aayfvFu6LOCalth
8TjSWwGWskywqka2r3s9Dp5KRebR70UK9Lu1oI4vCkCbI5DH5BD1RHY7xsLZhZTe
7VL7I8lekvJcb/xZ7VNja3l1FvYN3KkSiGzL/39Zl7v6jmqvQcMaOkZUQfK8bW6j
vOokBpEEF93QdtNqtVvEBgRlGMDLruvar3KW4/+DNQc3/VHvNrMX2daDy7vQO7Kg
apOrlf7ql4jz+KignDAMCT9euu7k1QdQVY2eK6aZNR1yNIPA+aS84VZH43kHtvsv
SJqEMX+wblYQjGFL8pzYp6m4tKJbxpeeQFl4FVIMp/23ebecPww5tV1s6pjGkcbb
WjyxQbE5LqKZxAYt3iGPvmDo79pQ1hLaKzIYRkxzcr+Ybc6YPVhVKpbf0lBFYz9f
GjZsvoYKylHcrjZ4//zrwr5FIvN0/ALAKfanxy5YVyXez5pOMxDTIdxv8k7hAPcZ
26feBPHZ4gm0glFNLlWQ17qChfQjVALvOcfBs5McgT4v92phvgGQXgkP8aszkUZs
NYWCg4qKf92PNLzftk8vD7f6mrD1hhF5k94RmCuEicaYAk6MoJj2Su64Xt5svBVa
SK/o1bM90H54r0F83tc3/Ezog3cI6mmUrHBXuk5Emvc4QMMfGkApAf/OJKUQS1Va
z2BKH0OudIfZ1Zc5K8AOA81tyxxemg5OcXoc9ozcGxbzVqJdP/tbXxjS9Pv0rGIv
dgltopQNuGksKCawtqW4Sr7tx5CR4aQ/RF93uZGozwA/7cg7tW/fbplfiTH7xEOj
Lqi0vMwRhuIup9ekY6V7TTFn6wHoCH08EtsmJ4gDYZXc9GRRu6WnnuTOeDuSATPc
5Y3iHnQ18vtEg7ivDLzRukM2BVZ3z7CpZ+IWGwlNTS+OfT1v2uHIZ5N4tSp8hicI
UOuTnrOuTFNaWR7NRBAbpFboWUQqFky4xmlv7vHqVx/ZGXWhr7rUe8ZTW1IP9t98
kYE5foZWIsRVRya9+40gKugRk/nV1W+HW5DxnaSkkvF+4SEfdT2wkxy3ia5x6s2g
mBDwDQWdaxws4DINLQFp837jOBJceXzyx/wIf1Q2q0mhEMwxp33D+olZdoEdlBWB
CiYJ4Xd9oKHqXbJ5R6//pPDVKZ4wEmdQAcJRnpm5vuReAkPrSlD4alrLRiMCRqdl
xlwdDd7kon8EBEgLDk79OlMcAcUWuaHCVciawbkkAanpOf8Sbf8MVJ1igco7zHot
hQ5dKNluftSyTqzjSIjXX6SkTFQ5iZrP/3mGV11KKJdmA6IHBtEYT18uSnVc7e1l
t+3cd6POAkVu4C/9kpcv6+xe4ZIWtp++p1qIM/f4m+pRdGoHQ5g9H/shSCDMqYA7
u20BB9bTZ3JVwmb/LJqQL0eBuryzjHb/isvJZYdsSrKPjQ8FO0lGfJL0N3+M8eI4
sozKzsVfbf2mRLRXelQqITZIt6YzS2m/S2/JXvwj546fxTbyjx8WRkylpaczHzc5
aeYQguFOtT12MLKRCEcVOShJbmRu/S8GBNYifzAYSLODz55j0IqrekBfNe+bKBNa
k7oAopLBECGtOtrr0xZtuJrdQdxqprsiywb+JEIWIW8hPfImKjOa+RDDjhrYdyIN
Mq6mDgRZWba7vsJ/0AObh8nIdZqsbRFMh41fuNdNusHx2CHxTxrUvMA/q/gUTFlg
A6BuqVdRmb9kmya7k0Iv2DjDO3LonJ1tNI8ufS/Vh1j+VH81ElKgaSLW7r/0mnJW
Azy/jOLdqStE4hHkjnsoB8JK0rjbplmQd7o7PPuN8LnP+OhFwlU0kTy/7UBYAEaE
8f+oT2l0hJebvYc8toa5H86vCq+BorY1H5XYoQP/o3b67B+GIPlvQ3A998dGormW
aE5EEVAhz4DcJls4IXGfk5qpATnPTveTHVR0rLUSPo0W17PoOAQC85TK0/cOm85i
mbrciAaCj8LYzG7V+S6S6f78RN2fp/GdH1YhWeuSDG+9W8UtNfE1gHRrbH6cCdFU
geUrZZyEtmMps2yLQMeAhxmukgTH4fjeFgcM6Bqtyp009vPE+CuZKw0YIeJRxnmr
0LJDMriEBWS1o5lK3/edmXFtKJPq05tqM5PX2KVqAoXd5nTXBf8eWAxnQVsWJuLf
Ay8YUtcjI0g+9zayYw8avrufbFeYjPHjAo0ShMxPW34l1DcR6ULhrleGgwVo/fMb
VQ4bBxUpAptPtyz6SFItvbjz8/3ZbtIPHQ7U2I4t6qkhT2q8jJlOfA07XzuNeB3O
3udyYj4qzPd9sSOhQSRnwZD89TJ9M57VpcE5zJTwW4VJ5vOZGcZZQ243JzN5kIfO
K2Azqmv0Uxd9OEptNSZsTQBC6C5ozj5eU73aernYoTErfLHOINeT6Gxq0GT/Kp40
zIxRJgXBZ32CeMoB8GRDrbB4x14uKwCKEVvNcGSW5C0t4fdHHbiJXmAt8hcyezCs
9TQ/+OLX5AhkbLR8SOqGVYmH9lmlSpJyFXhotVgcjKTTTte6y40rq7U8VGGbkNcz
rxuklMZKdYkFFI+ghvhPn0ps1gp64COehwb9y3Ffq3d1HKW5JN4bI1PzNIGVOszd
uUb7D1KBjY/C3ZI/C3yDF/lERVnPpawmBLaiIthu8ltxNTbKGneifKnmuo/SUs8q
wn5CQbWWlOA/J/0uxnk88gE9VC2zJXvhtjbIYQugzavWR+Jl5BCX+8nVLMVIxjKR
chAS82rdbGqEK+ia+hkwAWisTpJjpdk0BsgZKQW0y6DvGCnn0cUHsw1gKcJhJrcZ
GZPqlVsCMW5c/NeTERDTpCz5KzsE5v+0wG/BDDOjHjB5MZe42vAOjrUQybintXoV
XLVey+pSOUWZt5WCFa1T3N14JDMPBWiccnOGJ1GStm/nBVRlk9j2XkUYWFWZbrsa
f9Bz2KGsTZWVlt4p2ZzXy7fMo87OuFRo4DrX3imjMTsBc1yDd+6NqKRPQMH58UY2
1BrKQ73zgnFT0SaGe2RgwZTOuZEE+EC7s8qkhFMOZjhtzQxeS2kHq3DNFDA0U13x
t4ilE2/o2XvWQgivC5hbzrUBG5MAkfkImXMiLmZZgNLyQNW9WNvlGJmRxho7w767
2v+2HzcU/padvhQEPH/h7eNa7Y0rOkAh4W4c8syGTY80Yecx489vOaWO2//54Ee6
w3JqWEEBFmeDCUKT4BTDv7eFgdjsAI+hyPgOjcf8rxpZrl5nATvitjZX/5jTG9tt
n32Cv/HpKI+MQUwYHQl3ljgug5vuww062cwsecZ8TA5FeoxTIIDi/guFx7cahvbg
UFtLyowOZX6k/VrYGBvyseybXUHveUY4TXMpIgKx0pxdpDcGdSqlbBnZZoxHclZk
Bq3BMNNb4p4b0NUaangfkFN2O/GzFNemtgTw4hCKMW8f9T7URevIX6zFYFW/l8XP
P9niVrHTYpzmAn96HA1sPM0evzoytJHeWSEzxV2F18LjLpkFEjfMDB0Nai0GlMdI
dY0szvM9qkwJBG42gCWS6P3PrmEizfMNqlNUaAiXhe3OUGBbNOxD5Jd5HEI+7w1M
JOqzIMfAjtBqhGOAhx338GWUnHsOuDeXFnYslC8nRpGbPvQ8LFfReqDp3gp+QQvk
ZpNE9/NZRVzzIN0xNAdSCokHNbqzUhvnz/16dzwq3998fNquLhuREr61r67VFC+U
vGoJpEy17qClTJm0lLCeBOt2CrAj/Ge+QgGQe2qK0iBGk9dLvv59ozAkQV9D/DdC
vIpe3pDZFF3m58cl4SPJpxBcc8ow9MK99hAATkaFRaiDUH9GG6JlVsmcgF0TGVwH
QKYlHHQLRlWNswJiFilLCl0NoVtIdXewK3YxVz7rYQgWFQKDJ/XQYQk4+MAqz9ZD
zkf8eeTJ6HdRJ0Z3TF7P0L7ZhsrHF15mHKD59lpTRK0NMxouO24mb7wyWhEmRiwA
sjo7025jkY7s0dAPiEUyCpHcfK5kT4JN36zRVu7G+Zpwe+bzhg8vpeJmN2BN/VJs
7U99WEqG6IIR/yrsZMXm4QamXNM0A1oawq7fBrZRW4PCYUlbZ4SIq5Kl+GbAewrA
aUmwUXlCEow+xpPYEES0D07OC/HiFuf0AN12+ADS/G/7g00jKztH4wUJfq2iqCZI
IrlxNzzNxTMi4JFys1pftsIZn9lwHrRNX8X6fYs5iIjIzbfRwodqrjQda3ZPxcor
hPCF0kOvPbNyWpyszCCrW2lT0rjXpmRFCDMWULcBqN7F7vi0Kgd2vov0wLlKHpqh
aEbD9vppfSV00QMTUDKfkZXQvzB3G486MyzTxRuK+IsVJcK3PcK7yCrjBwl1XM4z
zXldphr/YOyDA/cJrEvvp4TnSLnlnHivQ1r/xgnp1kJrOIw4n4JwoS+rT44mxpdm
PbkZzIS2u/5Au9ocnuT5emiRD5hg/Qwp9CwTgECnKwJCENoMD2Fjap5wcs5AKgEt
g5ASwmtKvwHuZJhlPT5L92m3gFCHjUvH0jKzAzrHS28HvfFZm8Sm1rC5dBZ+VYl5
G2q1t2tkJ050GafdYQFro3MuqlRnck2SGXHUtSZZotkBbgdoAZ1W0TujipQWVhcL
7IY0itOcouRBrNzRA2z2ehq8Db2MTLxwtTdRqf4ioKRvxpW2QyZswPMQwMjZsAox
bw2FS5KstUVtnMLE+I6erjrGxUNh5yn9frqx8z5SWrSK4Txpq5zrZUQG+NDukcwF
KWbzZGlgnJmh0UWOLlZPDcWy2EXT6X4D6hE4rFcyB5zbep/KyqfnXaN63wTqniq8
9pFmlShAXHw4chWL4M3fqU9rRB/skULWtDnpI8wpIYDXCtHD83+eYJipqspJOHdm
8AMrZSr7IVkypBFabU76hFq2m3rBJnzb2rWBcQ3mcixmuFUG4jOkGaI+i02R3mj6
WNeB5TNPxdHv7kZWmEMZVqbmI9bey3YQfZBYqlegFmE5DlV4OyxLq1oDCAvWkvKr
iWE8LpbuIMEfisc7xK6Ib8WrE+6CccP5YfyvL34ZENMfLugkNUP1EEHMM4TMUeXM
45mgxZn4g4tT+iuQuFbOykhNZml9eUJT1hDbS7U8Sk1ikB/qsSbqKv7hbxYU5OLY
HDXL966uVoKHy5InC42V/o9Dwelo9cpKcNhNCn+BZJFl9UD9TbaGE3xkE70CY/hL
KuBqLHoaPHMq5sVcS5KSzJzubnvvKGYVGe7smkc0anOzz725OwtRiPKfLSrfpjbz
HysE/dWSWWHouRBnmOUK4R/eDJiWuZS/FQggbSjxpRFPeXYOfwHstUNXgSVJI9ov
mPCfplIovrdo8YBwIZPuUW2q5rHT684BopTXpRF/vgmD3heVo1KqWAn0a7Nnv7r7
axL3ysp7co7UllteM2RTvRPwjo768kIFJXXbuWeQun1DZgimxLsWIqm6pWqeiSq8
SBvfPIoCK+t+1wuTLvz/TEnMUQeR7M5pYXT1hbAsj8iy7FsE/mTkVfyhYMwBkBYf
Ft4Rs6yozvtLOVaRnDmDd9U5Te+Jzq7Oi421Uab5ohI6NAJuNr7QHbKU4v6ca7AK
nqWU+iRKF5lQIIPU4wQYk35vMipmtlvUkYAUeJfyRFKHcSdY+2+9sN92LM3ODVBc
80u2jZJdZ4SHJzMQMUKkLfh8e4Z9g5FsiZIo3TTHvns9+LtrKXj1Q/26ssKm6qe6
mcKiX32hFTbDur80lvmsDU1/82GLXMIDDVtXl5ObQbPy4vfirXPprytSS1i6+81J
GLHWjRuRW7TFWUYdxKpEwbi9e2GycvR7Ugj3aYSv7uC92NnRzSPNyn1N0mz5hGxp
EfkKQkrzIzJnwNfYTy9V8F2F1eQN0Vvh/R0qJBCtoj9l+4Opiswy+baSOa55U9K/
kX3pF4yGQ3aZPn958xpncPKKBfsxpaatzc7A/A1e5XnK8cG8vN4t3zMkcpnDfxt2
SzvG2jxG8M3UC+6kL+Wmo34zAMOLMAXWpCV/wT3yZ/oIR+PcsySgL13HiADE65Jv
nrn2juohcbeoVYITXEDJfGAUyEYCRhiM0X1qHi5tc2jRtbwbcVswKhwqH1QT53cj
DmUHgkCDHERjSbavKm/dYHizly/SeQeHlr82O4iXevPoCfUp4kf1gvuUh90eag9P
P0TAP4m3BDrSiCw/DaPJcNgPUKFnsAUzmOgsrOBozIMcfVKgTWv/XMNATEAn8hSH
vinxSQzNcPr3kPpxYHj7f86WKVd2FJbSMNo9IU06/QRPv5tGgxMbY0XT8c3wlhpA
zMVBYZLFfisEAQpm7t71jv1oRWwBHugwBnSwJSJBP97ibR9QQ/9+n4d6J4XRZuUy
CIl+1Y0M6EV2HRy6cM/TTTVYdqX3GcMaJJGMR4lT9LU=
//pragma protect end_data_block
//pragma protect digest_block
6EjRo8FJnKLysaVGxVH16+QMg10=
//pragma protect end_digest_block
//pragma protect end_protected
