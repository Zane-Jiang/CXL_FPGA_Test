// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Yq2eDr//VMAmgg7IkI0FiFJ0r/3VpJqRqIRIiZLj9SE+6tJIfa8znT/KaeknEy4s
21jrVR2waJYuh/fokaVKEznyBDbEVELRUoPlcs8e46c/6JwOR7LFfYw0c10xLMGA
tcPnVu4sTdokPBidk57KLo7nNHJmmpdAq3ehEVTfz8vDRqYw5e6pRQ==
//pragma protect end_key_block
//pragma protect digest_block
3OIUoLzWJUD7ueY8cU7gDFEALEQ=
//pragma protect end_digest_block
//pragma protect data_block
9Pt5P3GVHxhLU/Us7PUWEbJL6NpB+I1lkJYlkDd8Mah94t7a5zE9hiekojxyMxy9
0nR9UVDKCm2vaN7EEOqD5cwhZGcVF/sAHra00zwhoe9PLv2Oyn/nICLXF0gfY2XT
GzNEuVfvnP9LxB/NpgluptjZ3B1wSZim1GkTH47iyISWzN6d286bPFZJCrHiq2wB
2jdCApmDZCEbkup5C3gCHkBO+Rv9uqrF2XjkxhzQfYDiBIFBn+UE+D/9Qf7mNkhB
t7I1iP14FeDSCj3aeF3hsopngzZRG8e8ck0Irb4YZzgEBuaEBIFVETBO8GCZeUUB
ogx5VnZByEcbQ21uF5V1YeZnUU7hxA+ZDkGSxq0PH9aNO/Q7frUARx3xodeeXPv8
dilEkJw8MNaks7KXHjFqyjyM22FZFS0D5LwXhbQvUiFRG6N4qs4b1lWN7Omm//BC
KUgE6NsGU38Ve7bHdaUnDRiH9vlWGWBUYXylJHPXy/JkBzdPmy/dxSKlYvBmVCMz
WTZIK/VFGfc7g4F14dGh4HEw+92w12CGvuKrJPKF8pwMPjjgWwGesqLDqRGHtsCp
Fet9o3oCniQvVGo2aViOpC6GQLvpjYCTwRJP2b6ufKO3KvZORe+frsGJNxAZ5PFT
o2ambTv3r+wEnSN4rhdMG/2aNUT8t3XPv6DH7DpIHRkd8tCUdln4BfkCPPiXwq7t
fRy8ZqSUyiKHjhqnvftAKXL8p+JShyoCfbfTPCObjMeZWOa/3rbCXxMiaUjzO0xD
8YwCcLi6xgVNIgXnG4P6fdszgrKPvsvrfuMpJDW+SG67mHxY7cWOYBldbAh5FoVP
bwQ3O19qcx42kiMocwhI2FD3T4AkLRDSN+WK5IzM7zr2pZ/4aZvkQltZdfMFuWpw
jvEDLGMW+8kgd7RUolvBS5whPClBpVAVmVbCUaDrU2JrUNuFJLPK4iemSYDaHe9t
7EuPM9lTnMLQ+2cw1cV+XZfDqpZD2P2/7Kk9NFrBmrJocDOeXifEeGetavJuRhvC
/5C8BVmgUTVCWVw/zGFKsz67tQ4ct6ggN5aHik0DBCs8bfGv9Uapso3C2m1IwWIm
d7nQEgFHT5TkjY5QvXYGbldSs2xFxvJZN4NKLfXiPrPF3WAaxg1v3/fo0gbgWaGU
MXKnF1iR7Qah4ECQGzMtQ3AtpSei4y9xEerAUw8XNQgUuDDUqiNBbwji+DhNJ+pd
H1EaHOsR4VrnN8fIIpMirlmPSpMMVGLYMyZnz0Q4uJuCfYhoxYGJBiD3/xynCkMS
UJL+AMTRVrgTLu4rnllksHZmhK3PIP/vf5r/u7JPUjV5NP3KYxxc3HqzwPnzGjvx
is76WPlrD8KWKZ3n7WLqDoaWsymJ2pnkZlwqGCIk3r0i0Ps3BAMJBKviEFyVh54S
JxAYMA4JxhcbHuPcN2VxISd7JhmzwUBzwQpCb1kucHw8zPTCnpiJ9Ooc5pzz9wQE
2xdvLvcYF6U6eXcQ6xmx+qPq10Po3Y5sl/giDbR2APe8CfSLWLRQBbzvrbeI97/e
bnlwZuNYjxi03NTC5Ujd7mCUdOzdRVPUvSpK781Okp7f4kcbGf1FAzSNrbaeL3nl
QtPhm4utKL1okEV8PbdlPg/qnozsVoiGAnA2I2m/NoTw010aN7ruODNudHArhg/D
AeeJJnrM0tDIwt7EHV5PeuBJldjK/Wfq7qqbDOnpfcJTduFfdjA3NHtl3+U9rv/N
6PXao6ib5A8rN0zYfGVXldeCDhje1gqb4/fJPWOZ2wD3/At/fg61DJsj328OyYNs
xBoEKtTv5xju4bRQKnHYm90d7p9Q+sZ1bzvjEewIxY2rfvP/9aHVo1jPyqTMjemp
rc4Bx/iWi3Fcf5kuLTZDD12FUNdrepSWqAv/fmYRVoqL7jwLOqdeq4n3EnQtBkGB
9XBKGf7yqCruScj7rgGOiCi0B0jwwqpmtF+WePZ4tZ0wB35v9RMvkeu3GkqppIqe
GOcidJZ6hxPPARz8jwAfPfKLh+9i4E2c3av4cv/bpSYX9UPALiiWww/FoUBdehzn
2+gwjac58oksWC6a7L0gdcYB826RZQzlxqPfNdJUgRa5U9hKS4P+LTT27doMI/X1
+6QXQ2Po6aJi6TA5A32oZ3U+0B2+j+t67CDO1E7v+yJ6vv9/8m7lrLK24e1lbpfu
2VfHGs2xC/p7nhuwWV6JoGGsd/qLXBb2wL57NeOUawLG+BFFyD8C56BWCiw3D2xI
c6OLzn+3ebxMxKn3h1AfLTO0Xx2ggimfZcsX4ESSBGj85WtSMMoSu34L/i3ToBEu
qRgDlu+8xLOU+502QIyuYXobk5hs0pSLaD3BAquu2q0wjzrMI11SbYbNZKLiU/R+
d7jzPMXOXzN5wpmbbgrI84DHX+qApmXPEN+Lg79FAlPRqTdSJJk3MPXsZiznYOAL
rfbTY73m9GzJBS5C5eLL1D9dUw4UgcZUNzhZIj7pGrAt8aSRhh/zXp1gCrfnlcUT
PTXjPoip84ow2hIqp0WXchO87vuwruEL3BH5czh9Owc8IEnmSRK5katP4eS3O6Ha
rsXkvOYAMs444BWSDNe/7RoVWtjNBQm9LWhawMKub4IcWDnGwnn6nXCPKvOGIk3h
V6wX3rGyiQ/Eb0zlPe4RyRvZXD1roSuAsZ0XpPpxAobDut76F86Pfl71iIKcfPqf
RYS84KEyFkNICgHIai3EFNOt2p1zpMgcogf8Lh4h2Pe/nIpd8byOUKFug1qL2gPJ
bUq0ylxnDniXANAXEf5CfQgteY6rqkC8lvrmht4BEJubtTef1Be6rDz0ecHV9dI7
7vfU2d61ovVUVeVc637PU5Fi/eTk//cziY6G6+QXNGCMWV9hDMnE8CF5dXm/xvGm
mpaTXt+i+nbhhy3Ldy7sYWcedxkfOUyRyhWoYxEPgf4vdSW+01saZQ1Liy+b9ny4
cxN7AZTuTYXysUoDQfvOU2/7I+gYTIs0vgw6kO5wgpqOa4f7Clv8v86hWMUAEdNe
SwCQlZspiFJdMWrwuwb3/sNabDYWyP9ycS8zcgynRL1igFZKpFOkS8dEUhH5lc7b
UUgMolHXzcu0cMugWIjsAg46ex5QKd/+r5Izmh9Xfv9y1SJgPM9/ZXAi/MoJSR2A
Nn5Pt4sDewsP1FbVJeeokoHGzcrUo/cnr/wwM035A4wOlkLY6JHC7sVYD03EK8l+
U7vRqIAj5on1QHhapTpvRjx0xfe3CKLZ5uhTO1flDjZVRiHNpThVyoBeh5Lz9D7r
Zr96RpZ375+hgWpOSAFunkmOohoZKlUpo3WlRUu3yT7VdPz8ncZ0zbfh8KQQcJGi
uT+KAKuVlws0nrWD9H7cfpG/lAskpXoPleWU6xRErpQXJEJd+786sMziIMJeNLsE
hxZa99LNN9LMmfrnjNZhkNpOhGTOCrbxmN9ftZbWmh4DGNh0iV9yy6euLP7OsJbx
vEdaPyYn1coc0+Bd4M1qeAOzunvlGXKPWdcfiwhPfGHvD0Mu9QqL64aH2r+DZf+N
p4hIsJo43CpQeyxUbuxGPsjfllVEDZQYb0AGgA/34JbSj9mL1KS+fqdRImVAnKWi
LW7yPJl0OYZPdU/nlvReJ3n0RFLax5ygitRLHP9EhstHYvNAQbDBPxgZO33XAO4K
q2pvZfg+2t2PnpFArpf2ygj6vf1Z1zL6a/St/5K43aVlZoU39k7vXgMNuVel2fhS
Hjd/xnZ2n7M7cpSN6Je9nc3pIwllA1yKGTGnld2CQMbzeR8k4rAoVYLv4WS/Lz1A
nsjwf8uQMAj+W/kowtbmb5puC6LHxdYukOBlH99ie31mdMr4xUzPQHpGlCckCKve
m3F53fEiNDHImM9xNg4BbZ0+aTiEiy7C9zMTIRkkJRQ3fKl+JJ/+pyKh+8qCunud
CiNSF52TugXID+FpLB9UMFFY2kG9tIgkghblQBjaQvHLbKnTMVhjCixrvI/8hKdD
q1tWNUFLYzAxjjy4DBQ22U0Xddk0N8eyY8NxiqVuz0CvTJ5reBBNeGpbqoUZnyvv
r3vMLNMN1w/8axjQfdHk2JtyaqayiOGEvXdpFsCbro7dZ0u7WT4rZxXCNcjy5w97
zmoXcmKjY7J0iaepIVWD5xE5cNCmvGaeLNo0nZKoMzvc1R3VFkCh1ENX6YWNLZED
ke/jlDTtUJuXTZFSF7t7S0yOtqIrlKShFbzJlV83BrMipMzKbYcbYtQx2Kt59rRW
HSpWKYpoG3ykHZQhEB7k1YP/MKrd3KZusAeKStgu9Dst4hUuL5f36EyUxUjzAKhO
2nXzC4pW6rJrUno8VaNHMLuP2yFUcZ/NiNhodUItHJdoDeipfafb48NejDg5wxrV
WEbUX9BUAUy5GlQ5X5jpcG6YOaW0hrDmybdBvo4K94EyZQpZGHQSfoJeUiiin6S5
KtvdXCjUSzO31Y6QhQ0KueyXRMZBEgFxA/8rkn51+HeUl7jhnT006/nEjkKKn8Sz
0w6fy1BmoFV57lO7d8kI96/AP9bY8hYtxL3uZyQP1ro7m14HYgwBMVP4dkchJhsq
SIUqSig5oa2aNKb6dx0SiqXdpSgHtlzo6HEFoEXZJ4WaEt5kYUaidIy+qTegxn1O
WnMYjwWXhxeklhJmFroFjaA33cDzslsCusldBXK1dPezApds1KvHet7SEDsiteQ4
/awo4CIF8gu20xHnZkjB3xp/lkZAB/PdUVEqEfI8uyRW23t1QjvOj3BlofCSyXwi
KxP6a6pH/DSiLy4bcgCrCTS8lB3GtycMrpQuso7jCC3Qna9XqmHhVCx7G6NREDUo
s1S09NRRalyyFwNdU/BKEjrrBu+d619g7+8dfD60ocU4oSqgZ7cMF/bx+7A04iYG
gEoT8CWaa01ODhZSt3Ssa//nEzbgFH/SX4fBhsDdC0WRZLumXMfxN3VINtW9ps4J
Ns88elr+JXt+TXHoKhaBonv9CpqIkH4mH1sWwSZVCo5iTy+kfjqYeHA1jR+kELqD
yhy94NTLPEiSQhdiZc6gDiK6hIs7HsI9NJiR9ZP5e4rjZpTD17XNpv4xkosZHcDB
ovO2chtXofkSR1s2GYcc6krsLjTymfkQVmtjjElz/b0eu5VOU7PpiUf3OjDUr7bL
X4iYOSDBX90Wm8Cpz5p/maK7dVlZPH0eKZfBld5wJQng4b1i28K4xPnXPgmZ6vsV
XQqW+a1+xzQsLSuJBNnKSW12SKGqNt9GCPeToHyrK14KZN9v/3saOB+GsRWmcpz1
tW5aUyiwUUNnJK1FCDuB9TUnCowpQsnijdRF9xKXwOTpEsSpTbSGUfI5yJsGTqK8
iB3DdfIgilKm4v2r4jBp+Q5C3nbGQ0sEGqx/yg2fVEATi+QxY1bF9Z9ZSirSkTyW
IWAP2UVVAz2A6rUFSM9s6kqPkzfYHyI1cPqzB1FUSEBWBbhzdtkny7Uek9gTGR95
KrnzN0XYAy3JKKtcS/b6IabHQXbSN8Rywa2kmqfWk8JoztUv+KrH6u9NEn+creDm
vj1uS4l9TvczpDckbmQZ9ZZu5KIdwrsmJpoE0P4tu9y/tbOg9usa+1Og+dxiPEB+
K/46ZS9G1SNY0Ra2f7HoGzKmjE/l1TLQME/2bnJp/fHblH58Gwi0g3QzYCJMdjAq
kimFxhab4OvMvn/462oykeTfDNYNIJxZfamzUfn78UccJCu1JCBVWx2kSgbgKyHr
8rUOGzO8fYsmWw+SVWIfxspCwzhhQNTH2Yt/iXfMtJRoEze9Bdqzimxyn4XBz7io
YBz5DQ09aawbYK2ygdPx/MXwu0zj5+cRTG+yn1A0Xtgd09PPDZyGWAREblNbvV7P
XJMuGnFrRjeipCLLhC2WT7+7xqdy8UeGgAk/azshf8omlGHHrzB6NI6CSPXbqHrM
Ri+qROhoI0awUbI9A36O24wdOXCShJOFmPBGFIYEYrI6PJh4lcuRwNeEwWdcPGjG
y65MHdmgzOdTLQ/O9agvNnhxEWvOSEL2n+fJB4Y2WXGNAssl5KGvaK8xzeEDpX4V
Y7eVTx345T0+4jsaCgVrv7IawRMplnQUn+VI1PD9HuSkYQbqjVkbSQgY/GdVhuvX
J5zhm6tIx4ib5/Cbamc5aPrh/BZ5d/sroh5iz4pIY5TrBJDkABNcL9SBk2TNGQ30
K3toWHUm+wuGHugwIm5yjnxXe/3jlEyVMHfLBu+2wTPo16M51BHVqQ6ZpidhHJR1
5B8s4RXzLndJNIOXlPdZSGmI765mBOga2LXZPttckvCjST80eoIQ1w3n1RiGV2Cj
C0nDZ6JSMzisEcIyOjrZvScKOFuKANSVZDsMkplhwCR5J7zxg8hMo6/eT0KuuTdP
E+qvbuUGucuUzsEspqMHNHYrLU3uCfcFg+yLLKTuTmRCi/F+dnHPODBLz4j8nOQS
z9XNF/j7ANtFykBc9bW9NrDU1V5szTCfCFvmW7m7nEH5p7VeA2DwKBe6yxgwLylE
4I7PMqsOO2JsuChgGfmzjU0nfC1mEQggTlycEbzgvjKvXTTFQMth+nSdblQPiMh0
SvruDq2hL4hq2D70B0zeyuYdCNXSDMGKtbzIueEUvugSgaA9145/dRcJiIJvVZEl
ihQZsJ/9lLjof+3VsPR3tqN2WCwqr1UTjCyPfGrFomyRTvFB2k+YA6oZilEsyaF7
7OHlIdy8NcP1QSud0pjE+lkDLScztMp3Qh60x0viCQvSaJ9yOacPzAw0/sMZPoaK
2eSzqrM8mEFtuOI3NS82yvjTDW929pYGn7avESAeNkROjhIfcks9oJYRbPRO7gDM
u7bzw3NXXHg5gaQ00LEMrUDmayzPoY5HsbxT5kFSTDpBG59RFrjaN19T37jzYSOz
5z6aw2NzAh0ZvNG3NJitXO44EaDZv61ifPIyNfbgbYhzaKzgQY7GACrtO0WbsoLc
Mq0euUExK50/fjKzcV6QejDxUiuI7xm/E5mMNZBBhKJxE8YgX5kzpdoQ+DnLW+h2
LH5MMflOK0nCnqlDsJb1i8n9mXxoSO5mQFwJ4BJ+Boz/FbudD0pzXSVVIPXCc9m0
DRvrF2ZYvykdc1ILf3fNAM0i5gNMmgmATnqxjpqx07ymBP2ROzLalxn7NAIG7BRX
ZdwPAaL+mZkqC777gADh/vVw3I4oEA5qT2zh7Uz/MFiiR2ZM+gPWK0iDLYsQmNvM
m/nT07Y1mlt6E+AnGddB2hohuuu8SyAjOxS4XiqGqvZmFVYxraeIZBtU0ZeW+5w8
piHuu7XSqD43q+80+QZAdVLPnRz2i5gGJw4oyMiOnmUpk2j2f1ej2ed2MvAXTV9u
ByeeS+TSr4ckpIJPdpgGYSsjnqhZJejYPyh7HaelDaaU1WkHaqQbFsq/jSxqWV9e
+5cdNzLwotJaL8uDfl4XsvAkg5+pkXMSAAyeA+MwqU9Bwe6iLgFMxGANNH2eeTsH
m8MjUHpnmospaMO6ahoXr78j8DIBtZcr55eyciwS6AXe6NptguRKcgaA+aFp4C0G
nUX4fmNFtPTq7UmsWnQDClM7SrnsGv2tURGa3RGiC/oBAH226Er9JiK5tSznSCZM
ECkSbpEIxg0bjR1yvrSM3bTSZ8c6MKxKi614h+g44HMFIrKi4Qqzww7AvU6+46JG
8f7ZFHiqOo5OzmsSDiFWuboSIwacc13aVHDtgzJLk1WllkuneEY6ALG3geNYPClB
tM/O5UYtl2X7x+3kFDFkb9I5GPOfZgYXvZaCOKxpWk9PuJOK1JERhmyLyQFCjBjb
LD8vBUC291R0RKeYooto2FE2csIH0wGN8HFIGwlToHYGCVLMW4L2Uz3CNATndYsG
QBKqn8Pe3utik2rJ1El9aqE8ZseXJL0yy+fd7ssNLkYPX+HwFBJy4hXCpZKk+Bj8
w7+VlF96b0ONscY8+B2BPYAwi7hL/G/tbjCIxwRhA/wxpYLsqCaWT4UrQAefOy5T
xFcO0tWdVwEbtwdvk6EM8FY8EOOtjhkB9KKw9/l0k/H4vGMvLyBPfXdTbc81kBjV
blK7IBT6g/PTeJP3fPfpQZVjMN3VjBX0QQuqzpQn7kMx6ROEdjugDNduzd4s0sts
7MLqP7MO7YbVMuQHV94vLzG+94f9WFAt3NNkOEqR2nl1fvyQj1D8rBWhwvDE5q3s
8JjGhQ2qG/ig/QYpaXDDExrFb5DrUGYZW4fI2aE6nWy1ayGm0wIIwLm7KMERR6Cz
daT5nj7lbN/KdRKpVpG/luQAbw+BGNIiGVlVH5w4ZLFBT4K+DhlA4mwHaXTRfAln
C+cEDh3luYnkD9WfDPGJtOJAM98EdT8kXyRzUURavSusZNEtjBSUB9rq0t8PEqQq
t7U6wxPRXfPpTq+PCQBs9zrie50rr2kvEJBUR4K4VWpeHz6qxETqwAcJSv6ucdIk
ZKeMxQCnyBHn9kdDYnKu8XE6OJ4a4KNVFIzIfUoq9AW5+CBKp9bru442ogwUPMU2
DPkioCuhH2WqNF4MF12TKn3yqkX1fW9XCscPQo3fXo4hfhJZ3ChHbp0Le0SGTuWe
yRQVf8T2xgP1b3MD6IbVWgpaL94IRM30DMs2K4jwJMqDBn+iJr/HFKqN1q3yCL1S
ZKPRT3WrvHD7Uhepy7gzPWdeFwCVQmHLBn0TCUI7WwNfbETdUItOZFcpXvAgnJQT
VtK1QGAW+ineBNnjsWScdKG39zIF++pMUKdwhiytXc8dhI52LRmROQNV+422TOH9
Az2LbPBu8t+50clyjj9GiVRYrqm4wlbdkTR5uaQggzbZeqcfN97MMQM0k5q186xH
LXgzH7Kat4/7/Bna4Lf0dhZdXh1juJx3ekmuhYQTyd6plBrc9Js1eWiS95EO0n27
8KgjzPK1hIjanCoOkkDiSPPmCEpYRTFi7xskWmSL5hus2m5zb9W+gDrBJzfNXDDS
106egUYREbz1/GUDRalfyGZTEqF9O0tzEfx3wuNLXjf1CBGUgSvzQdb28Ywo0yLx
KaixWPMZMiOITxsjcVCrjMgLY+5mB2OPdCwcoOg/TCgTK8FqLLuijUZE45OxuTOz
0XD0YXfNrJ57lUsjnvJEom0dD7jKg6SNBuMmWHAQqlfFu7O411uTzlVvSowjoRDG
qgiTJsIpXOZrY5aeUhbVLHPAX8xbvZ9vxddjrhyZvNABcS1czReF3v0shEeQ2ypZ
obGCSnl3dqRKQvikj9WVZRb3FcioAZYvXpaICgCuC/tXWNp39DpqmWA8bub6ukVF
T7pYXCpGz3ZYDV4sqOCrpvWfisv/nJop5wXNkL2+hW9lHdY8ZYCIvxgmI9mjiOIl
uvvqwwsFPPfsX+wUOAIne8Pws7DSVyqiuoiN/H7NPazgkephR8m8oIdJnAyJI2MN
hhpn5IV6txzeesob9AYYHxA2F+HWaxu/G3eIBpb5T6+6Zy4OOCsOz4nUk1S3h4wf
BzD00s0vFifBkqmiPCZezGLQJzmCX1T4/CZHvrpKjql96E8O6Z/ltA/tStfdxOOi
J/sqMHnC7eKJfOnOGCUqipql4ZYKvT1z+P9UGPq5i8RVMxDkOIQVOAq1N4/U/8wk
KNXPpzcBdJ8ITzeVA/7DT4/7DpzJe0zRbou3bDt41KJx3bkj/4pX9G6LriiotHOc
GwO5s0pIfAMTLHNYawUInsJ119wndCJNSsN5bSkXyiBe5OYNM6YYCjy2QeVk2U06
IlYsZwHGWs+XL7Wko9HfBY9QZISJSwGBz4x2iKRTmBmLd8CBCyj5ib00N06f+Ry6
DRY4xgGlcu3D3wvvMrKaBtTZdtVv81wSDvCR6EzHxdpgMdFEQbOPOVuVKwEfr/BW
zaH0DBm0myp1ZtgsCm7jV6l3Xa0kNA+kwrH53QEHPkJQ34W80WlkXtC5iJeB8Hhx
uaOPZjYI7oniqaQmB1H9WgmbMKtg+Bk77jC7KnheSF07j1+FV3kP+vAw9sptceka
fGZnZAeIYCF4D78goFzcLzOPY85nyaJRaH+MFEgC3GWcxjoHfvuSlwtzwmPFYsRo
OuRVAah1qDmgKeAuXKKrwLw+qw6QBGckRhPa2z73y+OhIgmB138Pc3/Sk03oVOqi
TkhAAJZ5d0Cot4eZhZiO3cs4hIMgRcXvtEy0QkDCF6CzjTrgYA2sjXxlrQiYi38r
yhmjT6Bz6EFx1lCC8RgIoSoef5Pexe4tCn69IMdbZXZtryjWZ2EZXwVpbYjU+OaP
DUwmsfyFwAiNi94+iDqjPqYaFdiZ+Cb+qBXupEz01Y4fMDWAvq7b8AAu7G2DjKgG
/5/K4RajbcOFwr/tBj1qxosCAvI8G7H2MSrUccuUi0sf/6gMpSKrObzQoj2REQUt
WfEFr/q1ad4D4I4UdVvh3CYEOmfCWuI4Y4DnsTvEgEJ6t9+qkFEfenDUpY23NtsP
bAxv4R/NS7aABc1ywUUa0ayenxhMLZS8XICfvJGfA1wWNjPbZwoRQzq2iTYmVne6
/MTJUgnHLgdVjSCqD8lHD+LYkmvRMZhyjqUJyqBRiKXPNm+JdvtFrz7CD1hRicXT
oiX3py15/E5xzktoOM+VN/XlFylgRUM8ydW9u9ohkCZP6Dxvtx69EyBylWL5xBS1
gP2d+R2O6f9veLakRZQlYaLpwaEqLIWzb9iXO0M0y/N0KYzmkuUP3uowDq0flM6N
c8ibeloK1y1gI/bBBau/bOkXA2Y9cnyM0p5dQub1/vRk7ldwLYr+gBCwGtCUVEWF
L25msAvvBGOk8OKE7N867PQhG0f6rl5g1VEeOuHNf3rPwAybLFPBvamtHHl0ENYU
6r4C5GASp/7lM4pE1ayvBiSh3cGTZvr+YLrHPbJ9W1eO3ndd2SMbLfSs5IdoKqbC
P+O91QRr19FwnQbDeSydpVpR+C6bvK7dcsp52opf9w2HDz9nFNfqeotTmqTcShzs
8C+Hw8uuuGgm5t9VYraNVjLIavZGEd/fscUM5FGJT79slmxCZtTPje+NPHCgNp7O
vO2tG8+2OouXvTNgJHEQWVPpgLz53yaxiIHCqefoedxtnlKT6DVk6ovpJycFqwzP
YW9+bfWefTFC4xp98hVDUFAfb9UJjN14YB8LFn9Uwc4PF2SIVadi6Xhz+14Emysj
1mXGiM5S9uL++g+ZKiW61LLBZi+ujZ9iM75kKKIeeB70QpOmRrj4fS3F8Ix5WyzM
wrD+GuLxB5pNhUXrdJYjAeM1U/JmUmsb3nMwicZJxhLr9vXpF2otW2cccSdTX6cP
UIivNnKK2g5Sgc+PttNZV/dVLoOq7kbN2xY/v8HYhvmvuj2auNCMfY6SosEb8zEV
wk6zDaek1TnLscZqp2XNrpee3f92CQJt/OBz0gcLsbJq4248PZFA7+1Y2mVmdSRs
CM2jF+B67Hb+hwXPvhE/Butf65XREWwBlQV9xyqAGgbyxWwHeGK2DMjHFLQad8Pk
ya2n55hmlvNvnJ36yfRYJQy/Fn/uHoqR2g2IkMddiaZu5HFb2Fifg92Z5D3v+4E/
mxCzTnA9XZK9P9zpGcYvk5T8yDHKzz6KvTnR8L99kwguehgoYmmMBHfycvGVkzZE
AFLX+bhpZTnNN7qJ2sRWVU5DZCLlZNbbB2/+o8w+Q+bHEhY1aNayeAfWcRNyjiQJ
qpQkWJXXX9qDwWOfKt0a7ToXfIsiDpmb8QM/U4AyR7cLH37hW4CHpMUKBNDHFBVN
tT1ekwEGbsJbKzVPzg0lN2vcOPrfL8FwPhCoHbRPcVMn1dGT4NV7T6V+n92eTi7I
cMu90zWY0sARjGzdmiCDXp3c2IKYBVOAwvRvbEAcGFyDVIX+l12z2ni5drpA0QQ/
7MRholQWYpojBWPs7aD2/ELK6VZgTS/Qun6EEdLSxZZClX+eYnr78J9lpee9jHVS

//pragma protect end_data_block
//pragma protect digest_block
Ky+II28PPWnbqbtyd/tGtBvbo3Q=
//pragma protect end_digest_block
//pragma protect end_protected
