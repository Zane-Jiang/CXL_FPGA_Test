// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
sjOPnmyp9qS1M6lybJy2UXOIFMdv1e8b5IWf9l1qpc0dR2GOdj5K1cnWs2GTDpIVF3tew86Clelx
bC26SjCu4/KvHXuqi6hPVqVuvD3Hz5NFxnqrp84zL93dJqjJ9Goc9FCvnWd8EbrnfffUwapuv7g+
P8Qr8gbVK12bL6V6eE2HVgBRH4nYaf7k2skXpI/HwB6iiOjXfBi3pOXMpQn+8j3wbWPJ+G1l0cB2
0/aEw1JQa2zBur3by0NEt9SZPX1CvCcxPx+2y/HTVdusfF6/M+zKn3Amxp1G7uZTkyZW4EUkRuAg
FBvJN9fRJoz/S3h4fBRKXgJqY7+FeiT9p91zeA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 76880)
Rpq0xUCXwhb+2KrG3wptenjo8SS5rNHwZVxygI5aGQHJtJ0iRQFwLnkmI4gXirJcldpOcyfDtP/a
Y8HS5WgGBEsd92DZCMl1q0c7jNCxPNlcdBt5KMnBdWUwO3Ywy6vtr7AOyCIJIN3iVWJZHpCOLm4n
eSw2/mybHUohKYjVmVJF/Kw3SOENclOJ0yts3Vhd2jHZ/eo8kkaTvzJYx/QHe5PSeeMBT4zI1i9v
Fg/cep9BrGYeK3U0NfDaocAAg+n6olIbCtJ+I5qA809ZDGAbvdi7HK8L4F5lDolC+NSyHRupqpud
BsA1rA5OOxoZqKjiqN51+feBBC4F9C4fUB/lpXMJJnR86jJ5wTulqg5GqO0WCG48wFQfWXhQPPGy
tBy/gC82bpOVJwYaawakDRULglSmiZcZm1VcN5vsu0WzGUzFVsC6rUwTH7RlLQWi2b32Fq9HkHjt
fZIX/e1rX72C5GvmZ97sqTmpFrCLPnF/0QBJMUzo4+UeWKRtMDnZi9LH3w0h3yAtvyL1+QtPTdvM
90MoxW75OsvUBCk5suz25wEbsAAdxoQac+mqYNvw3l6DkVh67Z5TbDx2edBSbSdtlqVmZNHQq3r0
1DYZ1BqcbZQ3kQ9juoHBvDEMd68kCPtXZN/a9rg1GG4MWR0LxtV7PqNpxcgRjnI19kHtwngBEPfB
09SWYYPea70uITa+XU+H1vAmbmtgYSFOdiYXk2cE48stWCwBQtx2SPeL+Fz7zcjsTAZc1qTASULy
enVJDymzA94KrXO2WuVQg6Z3H0WbaRyAshc2fD38Z5/3z6Ml2GevhIJimIzcdpa8bupX72OWBk3P
2ssg4Om5/PhRu8RW4UHBAsFAK7v+PHd1bxSM5yYSxFfyRo5EzMJbhygELyLmhGjPTQPZNfCxXexL
Js6sC/TQlWHqsEattKEN/TBHCFFV59qB3IYQBKJPacgWFzQ2o9mpkrKZRS2sUx/46wk6V38mSa9v
Ee6/6phatMqzV70SCmO4EUUfA4d3IcUo83dYKPE7kzuEf1gz4MS6e9vGEJgvxIn513WIuy70wmnH
wO2qtqmpjLSqp7UUnxSmlFyRrvP0QRG4U3VQqytrYgxFcjUzeIptAhd1nCkObwE67dA77RyD7ZMr
P4tZjEVkWP8yqQJw0+nrqYaOqAOs02fTrwreaFCUy91WzwjjTKgpwMiOphUhWJAYL7YgDW3yJ40q
CG0grkmfxeF/jIGV2RJAd7Rm6wj5d8LOnQQVzGFYh3QmnX21VwGuU2xqCshrEeGBHOL/HnBpuj8f
2a/JX9m+gh95g50X28vge5jlpyIMi9/txwIVw1IPzEhVCttVoDsI83EAob/cXDJjw9cSmjTsJcFu
WoxiMTy4fU/4qzMGcdwmxIEKGp6XkoHZtyp8zNwyLf8MrVT42A9SkG7APTtzWwszC30Ah+z53VKN
o4QX839uY5x16jgwjOeYlgyZG+zcbIIGZd1qnGmkaxMTEQtqck9M4bcJlEK8VxGwg1yunE/Wqq12
/9/NhD4x/hkVMrbmec9kB2vpiz6TIu5nw9JGvaWAzFMUm44Y2iP6z3DTPVTJS1XnO+LqYmMSj2HH
TgVgbrV1qL4qWeBnySm0TJbFqOBVas8DxQ3D+SXAxg/xCF6Kxa6yn8l2jEQiMSP3pVcibZ8og/3T
/V9WafnimO9Vb947xWWBzmgHBspbROi+ePfqDnX65Qn7b5IAtaElGQgapXuwuohE1IAHbNxO4tiT
zSydJhVTgnFrJbAVqWRoB9GqZRKjX3HJ0Ay9eCacJTyiUEGLxMG9QXvnhbM9gvUdT69ce/bSDQF+
TYoVuq67BdUXt+4fwh7pAtFkL/P7EgGMAvt9MzC8DJNzpQ5qVsVYmgffy1xvj+4M0JD0wKm9EiqQ
S88hLBmUTpjYqOSMKNcWY2y1B/0u8Y4gJM5Ve/fVm/VvpyafbyqwogcMJZfS3QiOOMOhmsMSE2g1
1+d8dYD42H09rDzaG52jY+YTDITGRlesKsjKZ157s0gCHtOqgsutsC4WtOZ9vBXa6YuPEpasGAc9
t3551Fel9qxehSJ0kjmKVhS7cFFN9q/RtP+qOQHtRzp5c291nHCW5jwXjuy5oZOCOE45u+F6R5LE
opDE1gTn5Az9dktSrvCHbLBE1E/bsMXYq4XfpOeefLNaOzFy3iWzACb/RFE/2FsF2lUiIm6xoOXH
ur4z9uWSMwXhKKsI3AROy9Pj3mEJGITiNVxq7F3XL9dsRx9/PjiW14TUCBTCVh5Vglc1v7sF21xC
ysNV5Y3547/2WxSYk/vhbZqlWrW3ekYVa/1HPjbxhL6W+1xcHsCaJixf1uBtBKuRKCQdfs7mDvpC
hLD0c9s/uDYUPoKWQER8lCAtGdze0qAf9bgWEcP3bKFDWE5DbpvBs/djvcoWvFMxOE9ogHJU2TMB
hNwrHa4vo6eTOY2H1C8ubINjkt+gzB3SBrLONrXS1IEFmaqFe1SBjRVDX19+gYEZPWYSVEYK34Fi
SA7tT4ZacK7Po0zlsbwkhhIVn+7forOreJNMGpK1//2Ml0Icc3MBwsnDBhp7u6TyXIfIi9EkpDxN
z4/7G/uy9Vm3/0Zea0xHrnh14/bkpq9X75FGxWNthQx3jSwzIp/Zdi5opN6Jshcj/u1JhWcUUcJq
2dAh38sRf+K1bOjWtdbj7GjvHbQ1BbyZgXqQbNB9drFsnqdAeZX84584i19v/Rszy+xJP4vvXYU9
xK8L5TVevS7Vglqh+/HSHyGC8AoEHkX3qKEo6ecMEfc0B+C3KwQIZEKCmSQVDVfhk20ExeIXrxuz
DnmeYoFAqYhe0/qWNx4Gk+C4KFp8m11zX9TJGtJVyik/PiUPI31HKTtqIsO9eh0xq2lesnOjkouN
P92ZbDLL4kwzHVi/HflL1QjQDtDip+tIzWwUfhfau76e4VuhG1plNt2GhdN6fWdBnS/Ggov4p+gn
INyhEiDH+nWMwjrm8yjhX4tnGn4F9A4go6ZGDfpyHwWYm7eHAbrAXttc6lzEQxzh7dPpImzhyF0W
3fSH6IOu5pKCVmwEGsahhqi+yyelyL5EwTMGupwVnpQ4EbcX1KSyO8NTCoOvZNsz5DCwtPoQ85M2
yD1neNBkxZSlDGtoji9cI0SSRDuvLkWLzdAe20aTymx36+twDJ3m+YJOcUklmmwacbm/+cXA2jXV
nHmc2FTVTZTeSzM/BkQCcL+ugPU/JhX1Fuj7gSrUfuFbePsqSzWO0ELh7KVubAW6D8AvzCq13Vud
BCLUCyi+7ioW7C+c0hT+2HzKhxyYEUis2RqucGqjNH2/N1BaWCF0Rq6jbkbNd92KZPXzUm1X5gun
k9Wad/XBvrdnrLRZGdcgDNiMkD7O8lLCzazJOhch+4bXqRARsNBde5j/mh+sriUEpEm52Xg/9Jtk
eQWL1vasKp/fxFQH2K74VxnPEo5z0BId41+h+g+MCt2JSj9S0hn4DbSjM7Ns5b9aT2NjuCpuYAZL
lNvVh30VmOPJ0fbShEjlfzQ7O3hrGmjNp+UJeWX3xlq0wT3kinQd9W3/P5mwO2RwnpF1K5f1VBbA
rXI0AEmUPs3N6D8QsJpB7KEwFH044L7YDv84H5t4Ov7cQhyLxtwiBwN7UU5Gee/LRYPvjC9vT09g
nIVyRg2DYH5os0kaqSdnk5gz0zigTFncSjpA6SqCKqzkX/Ke1afpf9m7byzKM5VcWOc+8F/Oi/QW
QYdvgOO6xI26as9aJjTiDjIBViGNSR8KOhDascNh5G7iBYrjckp6T6iL4MkxLGF98r8Ol9UfiTZC
aV8FoyU3FTYNG3lzPigUXWoGiW/6bxAeZCGyKY1c/XV/+g73Ol90F3wmh/K6I+ziunQYufXfuNdV
/wVGB9l9glPBBbqExUhnJ8ve5FgCkSfDSQdFUqSik9+U1JdxJQ1Z0xIDXuxEaNJZ/ujsS/KHBpVS
rsPeEan4O5DlI0E8QZOtWcPF26GMQnboqebMNYyYqBC4lkJYYNor7fGKhhs0a/LWGvL/cL1nhr+l
01jYNdRlzg0N4BaPA6bKrED3sJ3ef6VHjawecnTRsrnu2omr3DJYAL1e5r0emOWfLjvdbjHMTHJd
3uDJuNLELU8PuNHpr8bXN1nHnoamepYwCbqs+57Yxm7pC2TfHHPcW6Lk9np/23pEqtXWKcd19tk2
qO60lXY6k1FF82Y4r+r7+bYlgXoFbikhb87I3E5y2ShKeQKFqW1NSepMSJiMXQVLEvo7JFToWxlw
xtyh6UKD/PGHMpu+w/CaqYZeHZHpcwZAQJoCOzQy8i9HMfhZdzzQ0Ia6Ep2/oRN795RMwe54abPT
78kh9BI+qTCNYD8rvuYJZhRFr9Gk08mFo+q7GHRZ+Nchs0nqWV0GE4XkNeuu4jbXV1XR2mkxBmsw
dAsTAEmIUSDCenYJeOgTjIVoqVa1CffOy68cWbokT83v0yzgohrvNhrdnCkyMNKs/Fx9XO/6HSOQ
AjZKucxmQUkXRlO4AdiqMBIl42OIOF1yoTkiAJWKMX1yzPjTs4Vahb9n+C+thhH/H4jCrOYULnPt
vin/y82ajwGJJZoKuvmMJ7nbMKlLII9+DeXh5hJWV8LbNUoFF4iojT98KrkrCv74F7jTOeb/g4k/
ijL1jJAi/ZMlO4qwlhI5DCBlvLDs0Vk18dHQSinIXWSN8qHXD/aXBwVGZdh/Gxns/t2icIJVpUY+
42/A2YvwaN2MyFJwsXq89SUSv6cg//6gn3SV0ADXq+N7p3RdlzJmcK0z2nfDx7ISC7VzTTLFnL/9
Nc8o0BjqEgg3p/U/xL3+3IvYbUmC9y3k7tzuG4MNnayGsmzmfmACMhpXQ3mOsPLeDyKDxGT2v+Mc
acH7FMHXGGuqg5WXERyeYFoZQe+QaoVN0xplX9PIwqF3wk9CsKUlz/RVzzHS9BggT9SJok0tXq6y
1FUE++Q3QBD7gRHE0eemmGHFA9p1CBQsfw9WCkymtvB2fuv3Zhfg0iMboE4BW/Kbun+yGH06YQe8
G9Uu7HRQsgxfYyB4fvrW5bepBlAMTaRTPMRSG/JnIEjL7nxgBVmHhRhIyFrpXmCnhXaK5ImsepgP
LxrBpj14/cOY0E6E2ZdvJ/b8ItLjbxBsVojuh9IeyNqItiroal4AjbG8jXpONXaVqn9pt7U0b8Nm
zzzx34xGnisSZ0fggHzRKBHc67rFgzgy65hiS9W4T8P8a77qmIjXzWkRFTG+BlXA+rK55u+nwlBi
Nwc+FZoBqlcEtilpmqactYb0HXPcwEW6gIARzoiYnRMAxEtyHiF+KytIjw27dSq1L/XJlQ7kPj3Z
evVGJsWkn3HF6Cn/sqHKBA38ChBAf4r/46/gdZlGpO5raFg0Q+r6mtfqZRLI8ImmXlLLVhZxJvRX
TFZ1H7GU5x8LAX1n3PBX6JGOpMSuEEJLcYodFHp23bcMonGm8A12Fg8nNIy2dgVbVqHYBVpxqDUb
tVJFF8OM8mg8hftwRB2vMhXL7NX3TccZmiMrAxKpdBzpNcGHUYs0/Q2LpT4TfxPrX1ykUIm6Tsnt
TlzMAnk3MibQzbnbG5XMW7g8bZgZ9cYavEWT2Xktf5E8OyJDn9cpr93/6HRzQ+eYc7ckyaB65gL5
HhF4Ug5E/D+7wEwbQzMMTlcDKfqyEszC1EPy1WYCx+wwPzVLatKHyrK9Upntg/y5vqrPfziZDwUm
gkE70vdd0+45cs4KAHm5rR9HnCHnxOJGMkiA/Z85tzeFgumbTdbRljbCRNoAImjtSUvW4oFeJNgQ
nDCiI6Sy7RvMvPjP3tYw40JHQNEni5ISMPtBMcFosXV4Ko4ZwU9RGcpKGL2VzS+Djrjr73Ja3lcz
5Ldexhv/uLGye3mc9HotNkNl53B7E+JbF1gHpo3oLqRNE+9flPUZXj/q6JAC2Atvun/DlsQKw3T6
e2zytLSvUUKUbVWY/B/C4K2riQ7NSOLbJDJlmOE+gBK/6tasRGn2ivOsi8wD+GAxpswOpbaIetAt
k1LU8q5mz+FnywfZnJb6mgD5aZAsrxWUcFBYgtbRKiIr3ZUxMfPBRgWjECDh/smkMNs+gyT/2zk/
rFgF5hV2Qe2aQuOnd0Vbqc/0wIthjjriwlmc0xl3nzkm210rHBTmZ6jnz+c7RkoP4aXNOrJ+dqLO
Zs/pK6KL5flj2Q/ECrPe0J+hNSG6Cx6HcMST1KRwd/JSM1NAy7nHPrWTTrBYe0WefIbTS/mxPnQ2
DMRTKZF0cfZWr4OdcFKQljMar1z0NpwURVcU2BKM1SNHwpTNhItZNb3iI/vUAGg46dbT5yY0buWU
uudY8yYP0Op/k5k0ij73U1g4zyfjGvmT/8MIF6qmZMsdyMT0Oq7JNSSV3w1u9Q7xkcj2wal5b7oy
wG9OGFt4XjrJTYenPTlB4p4D/N39CUWil2O8D6G2AdbzXpQVx6uGwdDypAuV3CrW+05vXziQ6hRv
JcCIJuha3/eoTXC0bBjtPCKeC8uYzZ+FxxMVOFI2Ntb+yO3fSpo13U7GtlR+uTgAIyMnRTQYOKbf
2XTgmxcXFXau4L3ASEe37wJ7bC77xN+medfixu0VALpgewVuQYjIdaklo3d1kp/P7W4nEsTW3cX0
n8cXwTEnzQ/hPAcUCaONkJmP3POboryeIo7YWGqTDYvy26T+zIPf54DnzYcy718wKzBw+j/ah9Iz
5AjiRl2rDdhbhFEdsm8TUcfBl32qqv1tUZzOjFfEKQDP7tKLQqJjSiYaf6dSzhOTSRaMbKTrEPWD
ama1ferM8WpD3LMheP71EdVmvpsNfTpxtlzrJLpn59YG7w2SAPUeI5ZKPC7jxGOzeWybYvJ6Neje
1wP81ljsQa96K/Lk0UcPhNRhK9hGGJPPzJjF/2xr2/h228PaUUpRUnEdaNduWFVSz+VCEFjS8L9z
XCsD9qNJT7IWcI35Tvi24L8dMmS8m4lAqQnlAKPJEwrNKw3sQqljg19CTSuSTa8Y5M0o1L/DuX98
HWg84TfOv7e8/glzbN6PEZ+oGefCy1xkGbEmAZHOEW2dPfJTUc2eJbbsMtvWI5Zo+ff14BrGyZYG
IhMy5aLRRXPh4P/Qyp1MLVdP8wEji48xowT+CJXhpwoS6sbQEUnNSSJgc+08ow+EvMJ/Clh62x8X
nFGdE77pqKb9O4orB7Z4dYRe/nw9aa/SfDgiEnZjEpd6KAsi+zu3bM4lDXHBGHhZIdPs0ewskVzD
Gr3cTWXGa22DPNuT9+Z+QKi6WHuN4s0RjDPvU29f38KkB8eC9UEgOqIzf43gEqUNqK0pOnhudms9
GVfIJD0uZjsLlk0cIKNEo/4QSizq391n+4aPToY+m2REMQxo7kA3NpKfzAIA4nijaPCrhHqJSQxj
PopVB4qfrEd+1GwxXuLvYWoduRBxOL0ZmG+D+0qyM3Q+MVbyfuWWrpRemKEnWWJLqEwTaWRhVtlP
mlRY+n87czWNPlMoaJLF+2zyQiZjhYI/Y/b550OUpI1f5v/YQI+GNsbrie5P5Avr7hJebKCKeSdK
jmAxzrnFR1sYxcPVgQSjZgDmd25rbfvBVuhvHrJjumkYF1kFPVmTeTxvUCprEnOstYZwqBjFqF3C
K/fcMigf4pam83UBNfA8jhX0sU9nvYKrmB5yZrJnqFcSBubmK7g8ukAnB3V+zoOoHqZ5Lo8UUygv
VGitlPJYgq4kVjTDt3/v1Hn8J0fu7IOw/Z5T98fVIHC2VNpOsWlROH1X7JbjiTgmu69MlUEuhaPt
hz4HXniK1jAlWxzzC5exqM+AmxrheCc4QgOl7CE95EEEgY4NTXwZOifgO9svyxDrPqp9tbfX7NJ0
r9TIKwtdnrN3Dr0fsjD+ESsULnQwM4gkSXtMyd8p4/J4wBzdGU2EbfQ/4mUuz4YegcGdU2xkPWyQ
aV/z31Kt1pGdEthLh17b/3Jbr3h3XICsf7tFs75+OTNafcpxUt/4BswuCt0XVh4JrNxSLCDcSTMc
WzGNrfsiRaXHhBkVINcgwAPtSizEv57uJJI/iKsJJrqVnXT43qRizVQHpnvkJOCWrFf8AMzk1a4Z
bQ8dWmPGq/jEfvxXeKbfKcg7WlSW+73lUZJsn9qB0hRqNB19i+MUFvQqhqx2sLIR1eLKLqpHfOkK
hf1ta3SFN4Yn9OAW1DBBoM/O5SZQPgmLNGG9FZnGTGQ8eod8oeS/DTLXTTTT8bCyFal0hSs2qNfl
i5QoYu8JFpAD3+ZEtbj6teNyPuJ7n8+s0LUcAuL2Mc7JDWIvgA4QDL5j2uAj2n+SgY2aaTs+I0vN
r5/wY2vLm4kC0mjif8m4QNXfdMVc79DZPhEiGsisP+3tpuT/FOo87fPJqWhmW3lhyagIgkbRKYtK
Qfeiq5JfqHG4CwB7+0ra753cfqskE1RluexahaXhw7gcleJiBPk0/oze1NybLCvCdcsFgO/fqN97
yVWH1wUvWN6EDuLHaojGJQ6r2malX0uL7g5UPr+BF+ZlZ+77sPQzqN3RGCtgoNUdn5i4/BakapDs
zm0on6rXeLlikM/AnJsip/1xSV5xTUoGMlc/Ai9z6xstZGySDaMkREv8+CoI0Fv1i5syL70Rnj1d
quRrmaZy96wfRDFvpVzfllLUgNs2/4lwOLJjRlJ5GmcfaGb66+vIUvwW2WWsLGFNFhL1KpnXKQwf
Ep0wwFB/i39GgqggbB97XoCXxL2bPHd6K3+Yd6HFG0i5mnKGgchHxKvwFCFUSTW5cJGuslv+BQ0g
CPkhNA/LebvR906RQ8CjHWeQ1JGX8iM7M+kKcfoZ0upLm6iNb3YLQpvTIgwRzpaRfFOYjQz1WK5w
uA3+NG/kCg0kS4TOBAdrDn3mmAS65oXYjz3uEKami+LDat332v6+VIsASjBJ9I4+G/WGpXkCsNR5
PtarzVZj++RX83Q/SYVXZQXG3JCoeW4RB8wsbS5WKFRz4KkYILxDlpWiw1kq+0tYSfW0ob5BsuH0
ke+TmuFZC2TFQHbLxop36dpcxMp9T3fPi0QFKN3QYUstJ7iYw5YB56A0UBEZe66rOMR6PfZwYtN6
gnqm5IzcgTpoDLRm6oYpSdY74Pp3utSocfVbqfRnp4I+N9HcggCBgS6pJNr75GLIRPl9hEpCCJuy
XeCuO4r6y4fy0Bnvev1LQPkGJ83HdFVxKg6ER1GK4maL7EGfTiYbLJeW5iDk9xQAKwyNn8blslwj
zg4VqBVhNPr80a6VmS0RkoTIPkYuXueoz9pE12+Qr4Qx1Dw2PTi8frB+PjQWNSEbk2p4Er3i5AeF
DpeIfd0tDHfH74hHlK+9Cnnbkq4ynoqCW4nNOmu5fjqS1HiSpzCjr5GIKbcskiyZdUUjk312p/3g
OAzGS/cruY8iKMz6IQr56ITS30yGdnifaikEgBeOenN5D4fhR+RorEEUhR2HOJCAQkbO7KvO68Lp
wC5UuXHD44fVIfGZvAG81la1csskksH+R2Tzd8/3iuFZOWpit6ehB6o17RW3ww80KRVHdUitbj+6
0B7egXtbJI4Y5SVThnsgLSFQs1J1CeLlmgFVPiKyEH+6Oo6IubXRF0GQwQE+UHhCGLUI+jD0zj9k
Se4s+2w6VsLdwlddSJTZ2xbmpdPER30D2yAY/OtE5BUQM8QnVCxPHXu4qYWzf/QZqRkELK4iBTQc
fa1iqL+/a6tGKJXUHE4S0YArfgZtFQYh7u2Q8Wb0BczVx1z1NiOiFot1g+PU8pp5KghhgUdHQaM0
A0GBX/0IY8NN+AOLqZpckalrMOi+VwJcM4C3dGbi1I+JlF2DvUi/DktItUPUm0W/mgoJdI1aH/6N
AbkCzKoDhwKZV0czqZOnWA4pfz6eX3qvCmcwGJ6T7T7rWoo+iVIVTfsNgIdzDUrxRwA3Jihmo/gV
SX31TlxkUd8p/kSUeLjGrqnXxrYu4sOyyp2aLfkSOXF2R6GmfeuL+I8+SrhaDObZoEOiuRnHH+Wc
z4DxKPgbRV4F1enl71o0nkSvh+gebmJjyfvbI1BhOGPKEmlu6ST3OnOE4fhbHDxzrD+h/JQOlYIt
Xn3mGoXuHvZFFArjndHlTsXVaHJv/DfCKp6iapmHywVQu6ziSJ2NJNf1yDx8O8cL3PeLX9m9pdlJ
1CoU/E4v7oSMpQypiahzmU9R/04CXBAybCw9UhGF5UkjN24bfZm12hM9x/bLHjk836+2UVl6cab6
33o3k/Y4rxsb6Sd9kvhxAL3aUjVSGWwJuBYZZR+TDd2mGG39gu1mjDgMU5dPldj5MJ50mOuRLYFs
EUJB2pfqob1iO87zec1R7dTrkNrCPINfpvxKc0jMBOteCNqYxQYe/45SEiXjaYoMhkrvvjW/ydKm
J9o23X1+o1XiUjxNa9dKuG++o4iLoX/E5Bsf1o7jNYB/rcZgLwMnvA+klJCW2+rbfn5uvoQZ/1HZ
BZjfTuPHrp5EoRENwWaLK/kHWEzNlMfbDh6jWsHTz7Ey/thaQ/EduoeSbCHrqWSFFXCsKZndT/Vj
UQERf9xYkejom+3rD8ifg7YG9Ay51ahKx7q7oBuQ+PR3CKAGCE8PUo9njHZVVP1XWUpPLQS+XpIH
7EeyAQwtiEhqfhsZ+xZfb1L27YjUtVwwEy6vxgajPaD+9vfA4Dj2TjatzAJoL7dzaRebY5/Bq0hA
90gkmQjGxTGgBnwAuUVPc5d58v2W6lvrygfWJPnoXMEIjAgE5psoiJgRdNr159OBV9V1c0kj6/g1
u9iVdmDfTWLFEFAzahPAywibaqJy+fZJvwnq4KVKA+up7n3u7l2txUVOQMQWj8XoGOESXgnXohCd
rSfY2yMpn1QQ7qj3I0LaD/O+ejz4mgkFjLfzg4L3wxpFyst2NEXh0dB10m9jFLa2+8Rbz3gHY1Sr
rubw9uMwH9FUUYEOde3dNrOyhZd7bI6tg+h55UBdx/r3NUZD8kfhtPxSc8WGh6bTMmvAJeDDwRUJ
zRMlz5QJVDo5bRnr7OlCJxJHQNBpPQ9oC7/DDNXMGsbadEiGzR4yLlg2OKPJM8zW2bHCWhksSNsO
EfRpADX+UyKVObR4N4vJCVaQhrfubikNge26KfQoWcP7EBJDXP8dbtpkMX5YMDAywAMdcKS1j/P7
d7OdRh3+s8JE4ZffUfsrN+y7kcCf+Nev64bPOrpdUlCCX/TcEuF+N/qgbXTCq7dEAVcPx19zOmsa
rwEg97JqVptK41YPgx/1jpLTcnJLJsXxr885urcwaS0x3Ge/EKeJf3QspyRxHRSh1rIPbBCgg8Ru
QuThNFXZanfNMWzvZSXkMLXgD0xK0RRityJxX81TQYqffdzdbfphzIbJL/tX9KASFT5bk4Ag1QNJ
ZMfzJ+GzGb6ngCuQ07ZaFxOlB89xHw+uBWTdFYLZHtL4/Zi2/DwcZh2ucyw3zVA8YEP89cquW66B
nWeoUeDsLtoc6KekcU5L4rUoW98Fz/0SPrqvPz96BJoTHk/R3iK7AJaKuCwpZfuA9LiNn+ijpD7N
JD0wWIfcRRyS6gnEnNOrgbc51bzfZFHq022mvQhOs7CrfEz3B1lWUr139ZN4cIYJF3rhNJdFMVad
Ine4HNLKT8taLanbgIwDeUKaTR94lrBIV7Hd9Fk3s8Rhp9iyf8QtdMVCXoNP73XPtfbZ2TTQInFm
3pwhfOdq8wNK/7OmW47sKR4yo8J5KEpSr5xSijIezCb+v/PdNhKLQXmlmAqGdBz1nnJgOctUY4b4
L8j6yd/N8ZUN3c0WkTVyw2eb9Jn7h+J9ItyzUYKFNA18N4Zc4qeM28BmKaNe2futv3gph1kA3t8X
b0Y5KaC4P120Tgdvc3w8tC/x9KcI81YqdNTojk5QvAxr6VmAKyqnA6H1oGN3JMzGuXzQlpCKxhYo
pgK/K+2S1Na93UBzj7DWqsgSfZol+zu6mIGMPRjTJ344gOl+E46qk9fA1dTmyn56Lg3whm58UQRz
NEZbzc/rfdjwjEVQTe5y6wI+qI3iFSzVNqXIpMjIFHK81plCbdG4/qKAYrvv009DdHGoHWgXGOWD
QK6F+XF0XwxZt4U0hqvrNVPBZL8zOYXvKE0xd5d7hnnMDFhBNSFVa6K/S5R0K9KXnIfZGaTQqK3e
Y3j2JAuzvq++On7EpT0PLeZZcqHDsP5zqUAw542b1jWdD016QEQGxydIgZUacVihPsXjbFFeHUwj
4TKAJIn6v7ZUGAATyGZky/8uvHpbQ5TYzirhw1nOSQP31T5vt0iazrW07NLLDlAaEwZ7FwASwnwP
wKQehgrjCCGGzPzLt+3o9hN7wlBDwQp185bSb2kFtgWipYKRzqMXCdIkBfB8BTiDIpNvxc3GtUNR
bmoEosnfDGvVKNSwpuuObuQ7+aq2dlPj6buLninWKjSDzNF9b6ATjm6QJVT69Gys+W9xHBQQ9kF4
oYA+BPz5fAtJPHVZi37x5gB6JV3mwRracHCFFV83+8DxrSeWxYMwceBPvhnaTwid9oBhMjx2tlxq
xhEjoCOoyO/6IQUOAQM6wzQyUphUXbMuXlPB25lGOAN4CRD1sl9ATdDR3zpYlHZR4Krq3qQ9srgv
mOi1KV0f+3ZVvvpPG4XAEpvnXgsGFBMhrnuvX+dN2EsNWypM9uxeVEP1Fm3nMS82rMfPoXzcnqOj
t2doArSwrCa4WVetLSSKHl889NpiLZ25mXeAqWvsk9hMOuPUKmS485JTxFDP3DcLRKtnq/xaBh3z
o14AnRXngFZsQwP+GnbuwpU8dRtxin+RXzLypiZLbgkHyswgv+AMip82IKSEE4G5qOXUC3Nl0Nk/
58T/Vc6xvSJAOSHDgpZXE9pbkMTYoPHOJU/q9cPuZlwItIaXrgIAMxVYdCrYfsGe8xx0TMQkatb2
tlSU/aCtNMUQx7Cd0+yvQhTmCuj2QDx39BCyyvyWYoMEPikoi3YkJtVSuxoTdmFUp8I0AoYhndep
kui9NBxrnmSc6/XLsxZ/7Ifn4FFpPdritzUBBmG12t4tnJK2VyZQrNbQTG5ozBJZsYmY2w4gyxi4
lk/Y/MVPmLG3yXHbzn9nYAvxilQo+cNqxdbAlzdj7elZ/QgR5rdNU7bdAo5k3yFXIVez3d87q28j
15aoS7TO+1c8YpTzuckJkpDOIRg1SD0zkGOpLlOGg64ymr22pQXJq+lA+SVcgaqQtRYE55uw7an+
+brG3zQ3BaxjYCzkpJ/wVgR0BvYe+q5WxYnNlQ12WktIsezI51OI/BJH7adnC8Pukota/+O1/JSr
X1l54ZA4ca0juxCcwCGO26WoX4ass2FRVyRoNKK53WD7xxPAa+NTaYTkqptFkQmjlrAzYxsTuTyt
0v6tXGKhEpr5DPiGssYLXlDyMziHraz7htmnXdQWAwJrOwNTCNE7zANtLqwDpd3XEDlmAWTC/R1z
729s7DR6XNsh3xtbdjiMaHDVyQMLnk9i2T6Bd7HRBhP9UrjkWNwF7vaJGMWTUw9XEK8qkzTvTa85
KDfD+LhWfryJpBfgHDO+8XJNvGma1w9wMZZFvASRNjyr0GmyZqvPM1Tx37p23YowZk/zXJmYxoy4
ISrnBVjALOQxtqbvg92yRPjqx8w45wlju37CpRyTSwl1Euf27LWPsOnJAH5LGrDwkbhdbeO5ZUAP
ZMU7lmROYFxA1qV7VDM+z4YXxD9+DAVZcl/Rl2U8ZdPu+d9O3XIHTDqRSP9fc2CBXVeXUKLzaJzP
I6tVwexnFti7eIxvIxKpuounD4+n5KgtM8JpuBwpuj7RMoX3NuDN+TD44UxYq3/WLll/1aINXUUn
yj87eoeGyQNMaaC+mKr6Zv7h16hy57eo2GUplcGU9vDYQrF1VZ3nmY/jSAXXOVco1hou4VXO1Zw2
WAp605uvkfaEqjjtj53Yc/FPcw56fnQALqkTp+Gpq58H1Q0CpeBWo0EpSb0YnDtfNzzFMEuV6NRH
XKoE2LUBKjaGMyXEZejGg4bMz9K4OyBc8q/f23Bnd9LMrVMQ1a17lgr6dkfgsO21IDl1a7KQIEqO
g/+MGgWWCGWuIgSSDAwjS9jJiHkKwEvTNj0bnQVCPVnwEXgl0F4kxvrsEat6/9/2vyYfvFounQNG
2ZwQg/kxDGOH7aTntAJ7zW82aT6kByFxNFry5NS6K/LlzbQbmE1FzUe3Bg6HDgqUrO0ZQyXyZoUI
ZnUJYMTcEsq6IH1HcKd7oHArVOrzMEIkOkxDe5KPtLT9GM+gAm5Nzmv05LZUc4HTbmPUhdT2vrSl
1PTPYflyFkmqveUoS/+cS19CfcV+74UBaQFb0O189tSYt9SB/xVFR4sTucnkjPvsqb2DYf8dlmDE
WhtNvflS/G8gDNMLGUlTJeyI20nBdF4IeEXdV2z8DcUL5iiXTw6EF3UWlURzyoU+o2z6AjPvrRAA
/4hlnZoQ/tWQAIX99nqV6eCOrJxBxqzLHwSGPMNdNLep+WPk7YhGKz8sUUqr2cF8a7YLFnNjDce+
XSQnuO/rZ7S2LXWXiy7VRMb8afSyRxGCkJCKseTfzEkV3+wrJdYVk9+tyL15G7qXcayt5fx9oT3y
LhqpW5oRrjLwmFxLG6n+i6a5Px7dsDNkowg3/+zSPLKqZsowyDFMfzH3317cFxnRnnnOxefZpVZB
N4UG6M1cgl1GalzePEV5HCsXQW2ldWjstvIXIh3yvQRCcsqioaXmPH4BKEsyMaDSUS+CxZyDueNB
Dv8jP5NNk+6dVmy7aA8XOUN4PNP5MHILYVtg2dcFjMDt6prf0X1jlo8SPNHeEgX76Wgv7b4x3H/H
QWKUGgzZ+gCHeEVlzs4tVWCOnW6ktC1yubZ6IfB7WG8chZ8ShynFP0QzesmijyXDIbUKYPx3XkxC
z39sqQzTCChGFnE26ZYaUypqbNPIF+5ueTy3xUR2r73KTc7HiT6BUPgslmH/J4ntj/s3OPtWTX7x
aRSMpiENub/v7gx2kUEvWqf5BLWSNAgOLYe1sdi7LywZtbVBglJtpYvRf5jXMIF1XMik0DlCai0J
crBo7hw3/H/QIhynLZYsoBSW2G2siSBqfIfDylCEXE5rZUMqvP1V8L/7xSsecZ08p6Bj5mBDRCzu
Fmvvv35ccVPnkyMnoHjm/W685fmchKrE/JSGpo8n9+/p0HTDL5uuRd4Csxn5F4IuFYDYiYoAOlno
WDIH0Yo7xlUjlODvR48nQriX3WP8EGPRwY61l57uo9kkxVZQnlyiWqzl8XM6Nx2gWGietmT/v4UD
HoouUruzX1rdcGQUayWKPMQv/zBxsU+lGS2pLxl8NgMQ3VIMhV99MCqGvLeInkSrszKHlViey3FG
a/ewVkVJTTk4jEe7zuomBIh9Tcdtu8AwXeOPME5vOxbJjJBRZg+hI7uW1EOY091xfWwSY6+5mcw5
k0xZEEZBek4fKRV7Hs08AmE0QC5BD0oxaoBtSVcTvia7VW+Kd4YCick8k5AqNStJnv4+UWtyqAQr
edogmb6hhhe7VzSg1dKEGX3XjJQaCBXoc4MCN2zaz6+DvGFjl1doLZjv5VFmFn3Y//DgM+sUGIa8
yQN0Tx0Os0yneQwTPu3hqVL4JgW8rMFf2qNMX+p55WJm2IeeUFrMy82aM40wqI/gGwLlCh3vhPRJ
xxSg+U/T7sUxLdftyD5dIk3seYP81io6GJnXRnbN8SypN0WTSJD5yvZTygae5Qv55QPZDOTb/MgW
x4LMs7+YCBIqMNdDD2MyBmxhsy6BblxTOB3+jwJufXKCCSGzDN3pdIkyBcQ6ScSYewcjhkxf9Sab
YOPUDZqb4hgX5o76MJiH/e5remkBAB+21N+mrR9CBVC5ehG6fNd1iH7CEGMhThrSu6M8RmLbx7uJ
vjbzrvztrQFnREag9y8bTojQa/hIueatAhKx//s0w/q4oGelR+zzYc4O1wbD/xk8RBveZzjtdY00
crZXc0+A8KSPUxOyUr9Nlx94In4aUIqzkNS4ORUzlCwRZGWUAhXpAmFLYvFh1wfKktg96jKcCBJa
6a5UxadwngKaXSXXR3dVYDR/15xTIi0V7pVgl1eX1KquftQm9iwqhLLYMJ0IwF56iPBdgM2kK2bz
1YVv98J3cDsrqNCHIKlYfEEaE8elwmZpuN1Clyp7VsR959JCZbt9NFnH77fenhxZLY/xLaQER+mu
eqgvb6XBvOccD7kicC2zT+TIuot8VEl1dWR5sTtJEcvyO8vv1pWuqVpKsZns6O1yiToaxiA8mjdm
ufbAs7v1UJl2R5WnEGsw4ZsS79g0fPNQvR4zgGVmLPAJyiUknS6MbVCshh6FaSVV69C1S5EIRjA2
4shp9pDtfJ64wnZe4hRAxEkORFaT9ifZTc19ZVrVt9THB0RFDfBRMyndCvR44+j8JxO5fbn3ChrQ
R33qP6ana7fAmQ4Blo3D2Wa6N3V911D9ZvMQDk3k9Br5QNnSQFp1t1HJPv4NO+YB3mJmiMuM6byj
8td5lSbVvEt9GnaBMLF70KUmLRuk11X6KBiT1I5BiwN/XbmdYlzi8d/4plM/7YmH06vJojS4RxDI
Mh45/U7OoynKeshM3Qya+nmXcBHOd1/3nEpnKqRLUAqHH0z+xtppj7ottdPtY5+5CSTgOgNzqPdC
7UYmGnq58CmZFlg+29dGNJosTmGainDnhpD1BbqCJQmhLC2qe6w8GUVy8JaHGOvWslPIduih+Trk
SXd14u0+585b4aW8zfmDjhNRmkgtKC4JLfDaUd2/RuRKCRIDa1VbukweAWLwUBJdJDusdifvGjOJ
wv7Vt1SIk82JCat14yPnrjnW5CLnXw7UiWpAAsaxdth2isqnVrVVYicGMZes5U41RZkZE9O6ADyd
xVcvW5HNL9uE/0UgN3Zh5rcvV7QkE8XN7cFuYRNlllusN7b8HvViOrkc3/KtpFO8O7JeFpxNtdv0
tObIO2gkzppEE1s+5H6xYYGM3vhj3G3aQJS1R7D5eH+i4m/TBkCUOfF1j1Y4B6jAIafiABB397+m
H/qYR6F1JthQUyMh+5nHIFd1z3XMxFeNqPfF+Tg4FB/IEBdBvXEeCnaoIrFiLIVQurvYvaSOHaBE
X21aaz+MTkqFYol1xR8Kqc+AAgezT//LCX4OQIXJwAukctKGumZTVQr1EVERVvn31RTt/UYP/UW/
cAvZFX3E3dI+Mexb/nRE1d5bLpTWU50sLb3n/SAOy2xtpGYr4l8Np5cVeVEC+jozxL2lTkiOb4Q+
TL9gD5uqPftzSjPcUWRmMhAouRIwm3u3V8hRn7kuBUo9au8XYeYvGfH4kc+uudFqIsuI1jG0+M3i
GWuNeyBwQHkThG1gtIq4zqVmMejSBxBQIGXGIqVgfkbf7iPI/9NrhwGE0mzbM6fTubbcYUoYhnkm
UsGjdrgfB7/+fLit//BpMJWm68wzlXZYnxM6jYXEA6AcQlICxT1nv26AhgdUqxpkHC+iZxZJVa9G
sxlrdl6mdnb6QAR0vN/eBfjSAbjjMVpvKgRx79aXJyb4egil5+IaohKdqoIGU6y8/nI+YodlTlzH
ZC7yDsJ68CSFxFvyrR6zUIg0qP3Hpa/DKkoHeEGnejb7J1r6ZvUkFQSlLXfyXKXidrmHJbcNcfMS
X8q7GVWfCb2vLfsbJIkct3l/NPEqeyBwEmZSU8G/D1r7WSK1q6tiACyyvqXzpXyun/PIfZ9DFTIh
Yb9kWKRpgm95KYRJ2WZ9Gm8mcjgHLs06NvpTTGHdoDoUH2Loe3HzZUHISco5asfSqZSwX0tMPjts
nLRjlsnDujPb/pO7PXiIIue8hSi9sojdHoG+Dbf2MeWGXoOMrZln9lRKRjEUiQnH0+orrtYy7sxo
LCuLNqSwxtg3AHuZ5dOuNk+oi3SxQIxJAe0PnFyq77eEREOoQ2YnewuFCwi6iB8nKOw2EQsGDUr3
t1SjJ7usVv3LzpeyVAVT0wHUqoA0UMmt9GQnqpO7/tTiEn62uB66j6/C1dm+vmoLZwzG84H8WwhP
aCipOaU4t/Vw2QDeHqGtZgoNM6amTWoHWl0pnX4icYToEmaATW9suwdPtezYeCFqwgXxHwJhoLCP
kB9+6DtIICsR6KKY+Y55jfVp/M7S3LvOe+85oCpAhHmt20xc0NGKBjr7pKqlseVce42K0p/hWc5O
qCj604kogh09t7f20lc2JLY00CTgtX/aLB/MUAVhU10mLjHbrIr9jq5MGJ/B8nN9sRuqUn7Wf7+V
yeyqN79bCB69zDOdBLEmE77llGMptbO2rfDEq+BROz2FgYfiFIvmLtITPCqR02ElKtCOxR8iTNaK
TlTOy7T9Y/2eW7tVDZa0Ow8tQRGQyvWxCjTZY5k5LMB6cjrTpdSMnejiFApM4/+CWA1XdkKR+3LC
XygX38N+JdpB6EuD2jw5Ga27OdkpXOqMVyLlFkdOrgSbeU2Xh3p4QekD526bMV/2Sn6UKZ/2fvfm
8tGibX0V0Vmoz6+Kq3X8Cwgw0kJ3ajjFQ8fVo0c2f6nXFpC+G3Vp8UsefXQPNMk9fc1PBHBsK0GW
g+TMP83G45RkxUlKr3n7mXyFj0D2RrIP/un9Hq/+X+qSMVPs6bWxDs1vZxKzPly1JU/HdlbZPE1q
JzFNyfS7rBlzgAaNNRFvdMvbezExFgB7Awq9ZuTCML4pJ8kag2Ax7raE6NKlg9tbFPvW/xPbrn/U
E3KXOMIMhFi7oBUXKUkQrZmYdXEyqg/GXaX+nOyveTutkWtpy/bfCZGT9Nr1+s7yeG/8nHIxE9zp
x2b3HotUENRw+gk9NaLVzVqyKTgaufW79VOfO2v3xjTlY2kya3aL4u6g8mIEcABa6CAIIgUpRI66
TEIjRteCytxBU08Q1iYR5cbVUYgA0q6BgIWS0ByVuTDsPbdJuA1BTaFHfg9/dUEU6tyo0wkCFSoZ
3/jl1tQGpkRMfrFDpnzInIPe3tg+hgFC8IoA2mSMXxy9GjUrVWlpUKW5i93KpqBHPBpEnNtk5aj7
6w0GdBn/Bkyqq/KG0BIAlOTZ3LlIVfEjDQFHXFVKkOG5q03dlOYixDBcdbXkkk6gO7HSJj/2s97V
e5mROncBnW3W86pLxn8COB9SICvt2s8KW1BHkJnqDPLlAFbbDwftNYej3P7WGSkDJlm6HjrzpJ2n
vnS0hBW4wSer7l5wY1A4hxViyshzWHHbFtOYQx2czt76vfml4Eb0IZyKbpO3bXnfLWKApDYWDLXW
zDp1IJkfNoQ5Nbu5kGD9JHZlfBoSxqw5aId8ErLxsid0SxFNTggsBNRSE6Z8IDHyKB7JD06/dn4Q
BnvckNtVPkv4jNhFQrtDzQDqxIF+vMIQuBH1uvfG2ud4dy5jo300v99sRHiCves6rh3snKK9S7Hc
yrPawZEaDu5ZrtgulAjSlhBAcM11PuS01TAb4BDNKgoOF3xxZu/V33gbEs3j1wg7mYN3aVNnzasF
PhUityAF8c2/DIoGGV6zyBzaLIc9leGcvdOCIW+gGPXvAi2Zrj/sE4RfIuMfgq9oW04ftiXhy6nj
Hg4y6OSJIuGQP6okcMROQf9VnXfOCHJZqENz7YrpXk7f+SIOBtZjV/mJLiPB6ZuhSTZWcoDI7CFC
IGXegelglfQrIN57JjTHFNINg58Kzlptdr9NHDLk40ZjpXqgtCpEvzoFcm7vYjk841Achp9FywZA
iJzVJyMgQIYiTYjiS2olyZc+2IgbZ7f42xt0yjCbYo2E8D/TQ3FOQcC8SoQ27uY1fwajh/ElJkPz
pgO/6HoPlBU7Vbdei8Qe/Wte99WC3SukDVaW5LGdUwt5XpFDjLRwCOwu64FTuSMXGPL4MJhIyFt9
y+Q+tNgTPbR1GeFrvEBmphm8XZxw4pOWNccSIMUXy5F6ZJPpZ8JCEwWobQIvVkpg2zGIXWgvDDxQ
Oj+LAwD4fbXVgcICXkEPa8FvwnuakMB8NSbzMrVv3ecAVhnjSI529pa/cxyne6gBBA+rRoJwz0zX
2NU4Z4oDRTcmVIjzMMfxgnl5wigF3jUXS5o0me/5b+xlDzurn3UaCQKNtXymeRIqBmyIktbcmTfO
za/1ozAjBA9acruJK/2v/z1HmGKLjllO9aRd8ChHsuIBVqFYAsnMmydRCi+5SCphKH5KZGzlTY59
/WxmOnZEjpHfUMMrt4qO+lT3PsmsuXn4JVpX/TNyYnRkleXWC53B9PdCeFvocDhOtE6cL1WQ6S5m
OrEOYn6fsE5Ker7CovCHtlEp0vDhVtMKKo5e5ENi/2aQqubNy1zYTqPQhp0qusLCvY/nU0F4fU7U
xpxtJInSGYsT+S9FmGLWIc+tXxj6itEWbPffVCyzlkHg1GkhSkpAjDUVFpnv4nqyk+/2TBeNKQbE
AOe1AFEzwykL/CrbDbc1R14NmC1+Lr61CGg5ZES36y1HGcfvQM/FWedDLYrBDlyaqZSCl3wIw4kM
pYBqUi5STxbEuubGan9v9c1JPq2w+2rpXrEUCgTUDE2+GB9kMZyj2FXwXDMHGqCYiC3IbF6VZ/Zg
b53BcaAg/iqXPefrdrHrRwFezI6glejdCgzZWtq5mA5UkE75IXDgJHN9kLOLDSgcfqh3V61LK+f3
dyZOnI5betkG2p5AvKPPv4XyhyarD8MuXxPA6sRqZsw0qVsysBD9dDeYx+7BmydE+yl2jyNnD7ob
AQKrtT0HQ7pjnOV4z4QYNemd214vZtglBeGyhdj0hQtzsq9CfEg6fN3+lWelmy1SZNya/VRxYEwc
8mJZ1nw6+cBhpumqvILdprJ/hLmzr0UxNMcCrCeBzTiyh862aCu8EDo0+gj0lenCElDWD8mvHZEm
QbheGFkDojTYMN8L0aRodMJ4g4CZDy5VAllXOYi3z9Cf6Zej9A8kunuhRJuCdfqANIFT1WfCwL4a
7OcBsaNI9/CVCVZiWweK/TeelnQIck3TzWDBPgsXjW1D5PFvXI5UlsBDPI5O03gKDIvYnS7FYEOY
qS1Pu2RRSpWScIe7ow5K6bJMa5NgMJVzMn/WiC0bZAAzQi+n9INiVds+KWXXVnfQHPPmP/4nc0Yz
X29twwQTVBP/Q5j1ZHczqQNRbl0lkP93A/5Iz7zvU+0M0lvlnY0BpRVXSFc2IVBhn7F5WeoxBzTp
DGUp6xsBRIkFdQSXmrEBLNu5iq+DC1sjLsNsDgE+mBdSCxTAPBfh1Ma89TJ4o5be7Ii83SH1yTwH
wEQf9fn1Lt1JZi7iuB0NCCi0KABDxkzOfeurujiQ628/dlDsFXzJ0LtUsqvOX8K7veIIivXEjf+j
g2tMIWggDQ5cgnjKureVQRbXEIMy6MNBLo4AQis1JwkbPB482QUsnQ2rt4VR3dK7Iuds4Btv89sJ
YxlXMEdqyYEIVdmqRgvaNHPVk/qsjUQS2rLsvin6YVOb0z0pnAkVXoGg6oJNFKbQhDo4DMZBkrmM
2MddpDqFxMfkYBHCJFgFaK5npYUpwrd9+JTgO9T3yufAcB10FWUcpCWQv0w1BN324Wf6gDNVuL7t
QNm4CLmDvfZ3269rKTfJXbUuniKQu21et4BAgaeGY2KsmTExy86rGWdX021sBK6EvAM4IfeP6GXH
98tZqM7THpnbJlRORjieQS/FDKfuzWDyASnNCt1z5eg9Q6idEkx3pcyNNoZfcHl7Tl1BPlU27mze
a3qqlC0AxHg/O5IKbRYnG3T7LzF/XmmzMZtM9LfhrgRm9eT5m7gwqZ4jTvxR/oboKxnz6mMZzzzc
OlOp8qKQJs7PBXbvNU1pEYiCW3zYUY3Hm3GOB8Z0Yv5jF18AZ8iAX26mUpcvJZCuCcO4TeuCasfk
JQgTYXxch/kiPZ9w3X+ZoDXmvv96Qjep6QX4FfrCZ2tKuB8Wi4jpYSDi63P3PajXO1N4ofi8aa7H
TGWQj5Dv8LsUCS34IEX9/Pe9tdgjyXfpDD+Tgd2EaErMMSuPNQlZ9+Ll5KMSX3B4hVabQz4DBoDE
PPu9jSQ81qAd9ZCvAz3qdwLtBdkWAH2xXtmGOpZSQvSN5nd7CrCopw0i5A8RzSfEUAwF2QnST4d/
Iiz+QT7a08bo0rSX1oNL5krT9S18uVFY88wXZ43U6YLS/FJ23/CSIr57lsYwaO68Zr6pAWRIp4zQ
9bCjtEdwouJcvaq7ian8u87rYgQwk6hhv0NXQLEF+daHr4gb30G+P+nebfYOKH5RcfscfW1CybWW
XWTkWpU20N9Ncdcnb6+ztHZZsvvQvz7svbi8fCDef9lrSXSWknCTt95TI78p0tMvH0H6hhbOY/Yh
p8BvJamAlua0lkokS6Qv6W6vD/ZYgeeF3j7FKYloaudqRiCsHdS2j/hsiJlACNw25V3YpjXvPrLD
nDLUXMG05arzhdNgRQP3Q4TkpEAB7QWybjfOgtKIyYANOebupbdf2vyf9lRAMHddeFN+opHuZCm5
YzbhRuegwl+lVVWm6ei6l+clmHwBfTXgV7pWVKyAJcWr7hci3DHMrel5RM+yxbwHA0pOheCiaceE
gAUmpLUucYiQ2i1mlKwFYTRgWharyJdo44F2J3+dJIy+Qi/nh6aEgH0aNq1Ii3Y8+oeqmrVHLorS
t0UvVrQD48O1NEGHedL+Yf4Kwe3AoyrPxEmAUxQWOfJtrsR9L8UhsI08xAHGUBzXonAFV3pFDedv
IixQk751Y0/pZSfR5/UqjE8WxLtoSKzvK7Im2VEuwPyWoumw7Et8y7Lpqxkpqdad38nvt/Rh5b5e
H3xI57BR6OHqrXGrTT6DBcyRLmCooFlaLswOuhDTqlrWHaV/TZnTAd3L6h1y3apvn+icNII+j9B4
cVLTnCWKe/iWGbd9UjWmAbY34u/QDuy/Brt7SNkDG61ASoizHf7tgH9cQBBVJI47ahk8nHqM12HD
oY90RKE4tPOtOUGVAMwusejPt4j93qUtLxRBpF31c/ybcKOHyHXfTOFzmIg1ifYm5G7lSbYrAS6R
0wViYcUe2B12yS5bLoCdIDnnOsO9Yl6/rKK8ZwCDtcQsILJZOlGqMHEWue/xq+F+v/4WhlvvsbCC
z3Bso7UZZ0fVks2hTYRu18TjIzkagXu+SO4O06cFHdI8L491HHsoA/8qvCXSfTdgL9HrO9is/PMD
2Vxk8KAItUvYNXrKK2/VM+h0+KKYyFvpn56AbGjX1fcpJWRTvDtOSVfTaIBFirhEy+8DqZuC165p
bWFN7MxWqLXukM4T7vt2bhVy1hfcIs4LxJTQjKE6kn6wSpywTCMB1XbxWOsC+FYyglse0dUQB8Al
FgjOTkrQVn2AnpFyO2+cB6IOgkhs+Aukj/7b43LlOedTtDr864y7PSJ1FUVgiq60Yu0W7ZypqwQE
bu+NPavGf3pMMYsMXbAM3wHD9ljRCjUAGPne1QOGj1ngRskG+m1B9oJuIbtEr94nZscSMg8Ro8f/
aZiFzQWnz4pIE2Q1Ao4ODvw0cf+iEkHQfbUQ9j+AA7cADYi+cZogpvoxFghMavkxwgJb7w5A1b9C
sz/uyNQLrXSQfNlMLLHvr09GWWSUWMfLoUkyi3eNhKaatNdGsf08GTPDjW/Ny6Zuz8L+TEkq3wol
zqpfA7qjxoPzrCunABe9evGvLbnOn0gf1azkFMNLFPtmqfp8pD7odjLwbGKL1a2T9uhZqZS3WaBk
phRrPnJEiuKiwgcwIQ2vqM3lBPZrT0wv7KpiX0qkTwbglzxivGoeBHVnTaAtZNg97q3R4Ed2a93g
+54myHVMHZG2/nghyjTQ4dT3TKjpqMft1onJIhqnHLcctUc8ysvgl87YPMDBidunm/OhFd9qNl92
OljMD63XftqU0apcDj+AKX9IF0w+sd5A3zth+uxPH06+S4f30d8LPTc9RacDZET6Tv6TCQTlPZ/x
Lh4JJoBdwdUlSbpxls2l/AogciW+hwG0EfeYXxltfFG/CX/P7IDjwaB6m9XPKOPEWOKRBmVXDM61
dm7twtNsCpBuWP1cHoczvPe6bxELD1n+jw6bOZBjsMc6o68MafnzJ947QtTMH9PjQ6IxrfnBdGSc
5DBSi8LExPC8kZtUuXMcxLMr9oenOVMshz/EClyb5aQ1b7mXOVGxHJD05XHhg3Q0RtxNmHO3ydiC
TfpVcftCXiquMQ4qjYImcEo4jofXtitg1gINyovTzlNpL2fcfP8c9TAg4zh4Ckil5y9SL/Nbin1M
Yp0rDLJw+2og1XCmwN7J40TXdMdVy0upzFH/odN6xkktNGTyq1BbQleJ7/VdkiNThuzQUx2whgKe
53vO4A1gEFwqY6QLrh7+tHGpjv8npaoT5ajnL/bhbU8z5UTvKOB5MJ/3wDxmXBVrLdLCJTMvMylu
TyBHVSuJyRxzLWiEthfiLtJ3KQBqNPx1lSSVYv1xdconPHLQq42efprToTtM5hTHZUUx2DcIABVy
SDq6vTCHbU655qBtcR47OsqqSoE9xdAL8/ZVXRhwgGAZO+sUDVUTzOKy/zVvDY8orl6PFxMT4g91
+kJl3ZMWEKB3J5kWcllb8pd9p9K+fWwtTn8Ssi9D83XvJDoDNDmfeJjCR7eC6fpXxbHGMVFvJ7SY
ALoPeY3CD1fiDpur0chGhzm9+d3lf6gOsUHuFQb9jwF+2kN/J8Z/RuHjdhxf4zg7ahFzrpzQkUvf
TUdykkkRo7QZiTRCSw3/bm+f0ol94mwchFIEv1kEVYfwk4mTmUSAz8bWCrfgZtDLYsnvMcJVbS+R
RDu/PI1VBoAcxdaInI5UqDNt45NQVfG2TKugty2ELIreD77UgcewoRXYVo/Aw/1cY7gw2XpY1UYk
iq9eKu30swRCYYkubX8s4yvVz2t++tVERRMqbbOkal0dCtvGpYOE+k8ZCRjqRnhZmTjZJulUefIr
vpT7h5D0hJBILmmmhISyxV0wNcUt7Cy4org3WCLK+O3y0xtLhsIAN7XI/yhSHFvLz41yEgImRhu7
XiML3DvkEwENqn16JN5fYyc7qQPmWrQt0ONYkbpSA6IuU+8b5PvOUnr0RJPhokAKtN0vBPzFnM1x
H1uoWD9WjYEPwhisakmaBB8zkA02ziThHvKs52M+BBHLdGmTzyrfigVGzKfMW49OQPQr35Hd1DdV
STvn3ky4jf/tpAcPKjZ7S3JMh4LGMM+KYKpiyzc1PFRwU1kYpsNuILUKjR3mpDh+n35yb93qbsfr
fNr+XheboUITtEr8/VwMr3P31U6p3yhS7PipBCYgGTntse1B8PW89pX6XM6rYC4bKhAkM57umi+f
Idp7Dw3eWwRNnBjCunWFeYP7RNf+wumYB1itf6VnOfmFvmUjwD4it2KqtZmwIYKNzXLhEh4l72L3
xeivMexKPNUBupGr2ylcL8cgApTfQOZ93Rqx/oHzrGbU+lY9yeZJm5Kz4LBcessBMwXHTDPd7Sca
6TJDzmsJj+u3C4CDi2JcxtXHBiN6lvE3zaoQ3DhepPJOdI3NTgksTueT8lAS/TQ2cJTpWdi7JKLy
xsGly+FQeQTVJP9ssHMA6hghghM0FPs9aMcay6B17Y2g+FIcMhJ2WmJmWXMM1xZqQnsYrC9Ct5Qp
AdX27kwNKE5qHoibI/da2j+i9FrnTdAsSBfbhOqRo8YL1uwNkiLL9h+7IJ5k2LyNpNHiGYkBfjdc
3E1mRUpljDK2mOeSvCfsISJeKGVisrERrcFIhkO0DoROKT1331Z4nJOfZF8co5iO+u8F6yHOEEOB
N0UMiDZfXEDl3GfukUNSDrDkZB4uNIk6c3wZj62U/lVjAM/3hxhM0K/HpkjOwIZlSlSI36x95DEf
tQ3xg+XA6OWbhhWlvDjXtZWOmUuIuEVtTW76Lj0tYUL9LipDdlJj2kk/lp7VOZHTtKqdaUA63CGg
gKOKkEM9oFQvnTa7d9gZAOmkTlRnIfYmwZkYoGUCScXB6u1LsmYHKOe+9uEytZfJgzIDbNPHg0Yo
+PyjcAfSCWpwszCGIZTBLBeDlgDxCzPfHOTpniRdKkZFIUHWRe28t61Hu9YMVQvu7pqqdhSwt+cU
89RhO7xcM5eMw5uI7MjDvc8juVjP0/mzzCOTfHcP1a8QgvYlS/74BJSElIsFQk2G4LLestEPh6Fq
GVtL9/pN5MjinlLZODKeeydLaBCyURdW0tY0RiwG6srIbtKuNB0HGzjaOeP3HQeu3FdD8wnyZAZp
Qad0e8PtaG6GfNwVtHAkWLm1bA3q8G/Kt6KVzbJ1fzp+BzxRJmO9BvmCwkyrxdozB911cX6yD4zb
ZqDT0sCT92G9wCdqw732QKy7RKhJGGdxNysLf3GSDO91JH6xbcHuXjgHjsMa4qec/eUIv1C8i1Kv
oktviEzhIEkzLV5KLy0x+eEDOXBIJfgUhL5e6hTa90bzudgs/t9+AY3pWc5AnrHbAv1z3eVLnVLT
JvWzWbbYQGK0QFhMn5g0s3Ol3tZOoqwFNCu8IMGPTTXLuwx3BZdms87B7O3cNbfel/0zWeJfbs/N
R0Amgc6q1Ob6SzCAeZrYpdf+lZvhetuvNL5Ht5T+FLNMjfYJxHwKVMoCh3etHAyIqv+DxFZwj7ft
U6CoKW3hwLpDUvjHWX0ia4IghJimT1cgvt7zDKYmmF3kQ0fzSbjPSUuKQ/B8hDnwriuZdC9btG43
fE/OYEN6VV3ceiTMP8AyVre34JbK6Ht8I877qkYK2454NN1+mbYWTePHGrnNAEaNN5PdjzLTug89
cHsXlKtfH/mhfzkcHGc6NJQXkLhPii5uHolRDPDQUv7A99vxIWcpMaSmn0pJZDEUOoXXveYa4Srs
l8rb6XljG5JZd/zj5K18bQE8uyyf9JMLOuT4HOJiuF0Est8j1NTLOADDxEetQcHO1UdqYoY5IKij
Hn7qglpoCIQqjaTnilxQXTvKWKv2T85weTG6a6ZhjwSnzhVJQbYWiwl3ldDPSM8n4R7FhXvA/Jrs
CyQMU2bSrZNO12Rl3skmQXy4rgva2XbW2qLcefWGsvs8b8h6HCcJNCWqSPn1CPoWHp6LRi7ONby+
0fkPYyLu5MYb2l4KAtscxFckC/3UJjF/n9q7HPxJfQdBdx9x6vaNzgQ4+C0eHkj9n2v5lW7aARER
wE0fIdmHko/Gp2axnBKCcPkOHthhnhFWEsPvPDdCRJXTnKXKAshUCdKRECNqz+Uf9sYzodWUV4I8
LaMkuUo3dEhjbK3MLaIpIJyreaBK7wkC+Kc2f9dYbpcfvQAeGTsu5YkztvVaPvWp0vBDVsIV8GGh
dAmTZzUkhSR7GgeXK6VcqycBR/OsQMH5wd3Npvt6+HnQnvGBRup/FOTjcH07lmVLSwEfObdxH/pq
8Rjefjf4DUSKD9GvKJDsEABDF6u3Tp28IxOubwAONArCGCx0ZNQQbV/3y8u4PFame8gjVB6XCOfB
v1VbABzabFNyF7e+Cg5Qr+yKDb6IdNo1FiRDduAAc5LDZpH2sHyvhzvTXuI7HsUjiH64548qnA2M
icBoL07CIYIpEN5gBgLeBWwjV2Hmb0svr30nY1KwjgPp3x0LeLateL7MSPVzC30lJLIYvSoBf09j
gg7dOaavX5NR+7288Ax7kw2mJmEaWXcBtFmLJyKWXufZSWVeQ4MS05DEGeA9lmnywU7W1alXiIoK
u+apWbthD3I0rJ3fKqOJFEdeUPS0xxzKvhK/ekXKMOh4k/NzPl/CFSqkM1/5f1WFVaq+j/s24tLK
7rcFangllngfISaMs1y4JtKfBWJd/Fj0HTPFEDSBEuy/dp9/S1WhZIlfjUY+p61L3pBV4yHkeuUN
wMXHM2Ii5/A6ixmOJgw1ilM9FxS/Z7rClJnW481oNItV9mDatesn8w1pe9ANbawXL6KkJmT63dUe
JZfVceVO7ArRe/OoVMDKu2fx1P4N5EuJ+ahOliVQuFdbV4UElsZ/AvZTmXlWwGCoP8i5VaINM2+z
joSlnbvofrSrhPcPsnLw1sY8qMB+EXFsV4MrFBgt7++J1+3e9ayiusnCJIydM92GZwJCfUZWrodN
VcoRYNFQe1y+OyPax7C5k6L+ffeFehbLqVC4fo8BL35dLJToJ46sAitkYVppMSJuzXknfyenTrdM
CK02HtzzL57msl2tTruNU65CfoHmfF5VkN372QPYaCGp+Q1t7S1eSMJmTLCPC60/zWgzMS5kOPCn
uWWIElOjWJPRflEpZn1/yc9tWYs2yYzy4vQa6619rKKxU/Yu3tMcowHbiN0Bx9jn1p6s2nXkdqUC
wkaCsAUfjhRbLULCxoJedcWx49NCf0dPSf6UxZyQ3SoqYjL94I1GWQMyHKTo0JJIKJJpDuE7UIav
byWWhs4vb/J59jyOZ4i1PgR4328b0AlIMxfnRUv96OilSQvWOchc4icB3RWNYmOTNMf71lzly3KR
ZSRkT9WSLYyOw9qgPxCltt3XIKw08TUC5ZxJgAiCmE5iFwUljSzDPa2eqQYUrcrxXhW0akCWIk0+
evaAXvUGhgGW34e97fZ5lmL1KncthKGlXNEq+hxEpjtrsECLBKsw+10aAxFUUp1mkpLDQ2yKl/bF
WbtuA1Bnw9izGjZZBH0XMIJ2o2n55Owie+b2ax/ToxfCFMor/42KaGZHDL4SaWqRFlCN+MLuuz09
VujG/I5+lgaGohk/HhtpiYwAgRReAVCVqLMCCSu8DMfqnnXDuOoRTppV9cY1cUfEE7Kpbdd12P3U
gaOGOzIu53Tks60tfL8xWgclIqjNc8XpbzFKgKW2Myt1s3jsVp2FBhKIKKLCMJkY8hz1KIelxJou
7RQijuz6RiKd+w4RsDu1tv5q431uRCHE8H3Hc/37bA5Iv++I4FEDJ7VTj9rEGF7+Vibne3G07v29
vU5nj3IYC04th/cqDoiW3Oxv3OrS32GFDg9EkupbsA/93N8wKt/VdlldmXuh7E7vQzJ1EZNMVDPi
Q02r8FgjU7j0ndHqvC0WgzkuS41TUqJ4LC/Wz5cmRWveNjKeKA6MRfQXWmuw/tLz6HTglRA58YZU
nXGZYircEfRfIBljmldGFR7y/FSLekOKD7f1/CZHJNZqFeEoJmcBSc+3mLOS+V3ehh5e/3rqEuDS
MDoQKJ+tuIATnwqxloeHIVTKbvx1ZwDu97mM9PvaSBojhF8bpAgDtIohoP5YSJ2rhM90pDtLnMYQ
M9xHA/C2Z5W91rKUfGgyTOC2PKNatUjgYENlgUXKJdVy6wcaLLmVlk43tNskKeHpSYSMOIVHejim
YxF6T/JIQhW0E4aM1abZC0gVaDMr91S86Hg5+lrbqPxQBAs7D054uY49iAMUUb3wy7fmux4KPy1+
C9Ku4KMdLf026HX3VUo60JYccL9oiLWx0SrcI4/dda8AMmhJq2cftA/GD3+frrpU6UA79mdbw40T
Xukik8pIN0amc1GpXWL/ZpTwYM8qgqNhlrdRpusyUls+XfGacNwMZRx/iQwBw/cditsbEQ9TUWWS
E7riq96VdlDPX4nouB5CzmqsI7zE4kIhnD2bVhn2rOOCeO/AmpKe0O6O2zYSMfVNGXwtWw4H3y1E
N/BR375kbMQ2v+y947iV/oa40djLuYEV4NeHiLJuDEKO5HP/4OE4ogIBhmJBJBQAECcCCubCClmZ
i3oY/3eNRPV+tz+0c9JLMhkaDwwMHAveSjJ4Q03Lwxdq71RBc9nvinCD0ORJUx7+PfF/ieEMDrAS
9rUqaaC29GAdiQ53oEx2+eLCDE9KEtXf76Rm7sL3lNPt+Kv5mS/D8P7TIvlPls9Cjym7/i0xNec9
RozC9cH28Dk5KqlD7tFHef9jD6YMu9oRmGxeBtWxoYu3AZdzvSStzPjSCqsrMRmENF7PhmoHVxlp
TWwgfDVpwsKW9nBrk4O7Mmy+w4MJjlCpRvh6Mm1Y+nn05KpoYx++f1l9ZzSZJaAdAUiKM1HfAh+e
Czt2swjnRoLKYudcsuP/A69zLmouIKYLgWwoFVGgLEW7rzO/J0YSzVshGe0KIZJ4T2Pq2uHofmqd
NxQ9bS4NKqLw2OjH3B16vNqqSKvqlmVFaZwPDOwlRujm0nsmMH9nWzlu1mz/a3eNM6rcT91aqNuW
rqqZ4M6SeZaoyw4KriqEcGNvb4xwoiBGFC2WrBReU1ML5z34LBqJNnlwSCegYq8vP5ip0K/+obGb
A9TY0uVsBWz6vMJe59Tgoa0/2ZbrTJXai8Uxkj3DgZGgzirpNEQyL05ZzuNDUQiSrww0MzO6NKMJ
dFQHiBg+DkJl1VphT4UIn5pE7akYkKtEIp2jUbTpgRXx6AizSdEZerk8VjRKevU30COEMqJSd0XB
kQFtM8ziotNmoQexlbNvA1Uti3+ANt3SVftqRPmyO9AAQa/p0o0IsKDi45MVEPgIU9ujeK8DpiC5
IYzXPsukxIZBWWFbFGle1Ai3lj2Q9OIrLaEHJPJFbcBfpNLCsyf5+khi0LijFVBGja4Lglc0w2RV
DAC5LameWrlx5/rLUe+fF++uEEx1BD/gW1b7wiJFR+xe963YJGXY0asXWhnZlmZk04HvoA8yiOcE
lnIxPRMqTCKWj6tYjdzDtCWZ00fyvXBBnqZDBl2FFhH9DydG+XLwnAEIOvloFoM10VZAxjKUvy7y
mHLVyPIRq9HfxVOjL/VIlfn9Ll+jiayahOVZLBpbJMj946RIQ1QPfSrSo3/6mgC4Z3UqBum+9ATF
eyWc0bwZTQUGzPShxpzEJ+qeKmx5kGIVwWy74y2LyrXDdGuGJ/BkzwJ37Wg+nzPjBqtO8RefmiLm
HBQ0VVlooc/VIYFVlnRhRtmaLrPQG+L8vXIChWxfss3viiCyDYKkElwt7en1CPUvsuuYvYyebNrB
9fK31P9CuwI0KevzwcA92rTUIOAoCz8HKnq/4D8wvD9NRP/dZnsk+7T6XLZ1xrdp0Tx+iwyENSWk
c2CmuY7FbuZbtBUT61L2TKXnCyXEtTM9TFK+E0wDBTfAwqhtEJiwoo1BSnm5NNaOri7UI6VhyJ4j
FuquZXak7Mw9IRaekMuPxIKYsB73T9tQyQseYSOVMQg9ZDWjKOgHvNc1jTc4CfYOEpBmuUYjm/1T
86D/jJphFw042xCbGYDt+jBV8G8DUYbMGsxT/ClveclgN/k3cIti9OL65sjTsoPf8GJYtwWS6b0B
9+McKBkhZzknMY1IuKmil5uiDcJu3sq4c3NcYfOIEgvMzwnrjnKatWh6zBrGa7y6aR+42k77SzQ6
A/lbz7N0vwcoOgHiG+gc/UkeJJp+ahFkTU+QBwDseQEn+PFTSXoLVdBOX3CNBGP8rpvvXn8CC7vU
lWohPuiGMnEcqhEYBVl3EMO/WEfUPObDOPbPBLD5Ytc4C/r9P1rT6s4n3JQf6q7EexxyJ5bzMK2/
X/3wT5SuDR7+R6HuN+9nl38d9GDZUXpVsV0PBGMyWcg2ozvxC+SB5DcAEepbrCBZIbYAXuFwMA9q
0TeGeHsk/WYA8ESmZcKQ/+bnDXwXHV7jEDiaZH+s/h8VoEtLmijhVLvFJkDeL/7PGP8oCGmFr/1F
wpxZgQsEiBVITNTcMbNj19jE36kvAjIAlljmiFDlg9Gc9RatQiLaY2LsePZJbVDRr9xx0JYwr14L
PoAuWzNss/CYnbvrMhgiOvvKv/QXJO9H5UfeQkkYnzvH9/JV+1fTP+pC+d5s4AuRlKfT69sh+yY+
KW7EygyAIROepnFgox+y0hMO6KIDTJ5TSRfA5ftWT0HknOAu4QVDymeD+EWfGn3lUwELACWhJWIX
EgFdWPUcGht7MWA8vEMepxzRyYSc8mbTRmsip/lg60oVdfk6QtoPbCFLu3IILC8ZFH0naR2Y/Z85
irh6LI7GBZSgUln4HP9hcj6HHh98/VaC4fryIG5s11yWKYOiSVY1CvX78iICuYBBcn+oxRIjU9jT
mrXHZAXlcB1hU5D7ORST4+iPZnsfdwGwIvNoHIpApXbhw5x8fvX8Clwh9PsEDDKCCNx1/RkVv1t1
Yb7hxhzw2ZNpRNFlVP/UsX8e8RAPnfzfIFlYc3UV4eTGa8Bks+ljYDOly0VrK9SrE31QQCdxuXNK
ljdk2+7MixmDEx6gXSKvdHPxXcEStezScOEXvBYsN/T7mzHCgPmiX/+HJaE6HpVYvJbPFiz6iXdv
Uy3bc5Ro0n41iMJ2PzqJ5+VwrJewsDrhVig8ZG990PTCTuWnVui1UrVv2pFZo3vU6joIufZ9eE6k
9DFgWfXKva5LcowV8YffAd1/9A2V0rziD0IQeweyiA1pIy59GqLPQeL8aBWTYApB7gFzxderuoGa
Spyuq5iGSxIcua7zj28ChBG+2SN/nr3pYj5LiN+nWdPi2ZJDkvql4Sc6m5bU7bkD/zdQi+YvgT3m
bSYxkw8XmPYxNveSWcdvgUbEoco/wDQ4FwmMjIjVtslJHPlgy9tPJ0dRvdA/GfW0jGEeciBUqbQ+
ef2qhyIo0uHdXj1GBK96Yq9uRkB1mNS6YtSu9XHz+vf5V3evpfCt/3X0sj3ATuRKj/JCEoRLTsny
lkf0w0Id9yCNMZqKkRVKbpKBVKnnXuK+lAduCNF8MGEQvhj6BUgv1N3V3AkO0/ZL3YjZLa9BqSy9
GMKq70v3okE/eBsMA3OOXukJq2y2b9sXO9qUp8tG2yuJv66qDCoeSFIzR8Nxwx0Cr+wRJPRbWAT2
gxlgQcfpIUtvZP5LxBh2cqRtjuGS5zJjM9yVdtIHqsGco2LKKbFk/6/OO3/dBm3SIG1HgjAZxCBS
LSuls7X7D7vf+gxOy1C7otyK64R+JxSsiVYB8jtzBnobjfz4U4YbCp8AQXdHHbtJ84JtlFxg6zb+
J2h0j2pBlo5pCPIzrK9/O65ypkEXumxFnzTguIWAShBr44NeXCEJ++2z2Hdp7j9IlD8iQSgixb8y
hen5+kFMhSR7TlZD9MXu1OxNGbnVJonwUG0hOdT2ADoJjPzdHHypLp4klBBCN6enh3yBV/nNWCHm
IMHTL9ykln9w+KmSJNFacM+YXQzJAPSymyH9tzHT09gAneAZ3n8AgoRjm5IQg4kd5mw2jbHwuxcF
Hy3WL+hWbkIOxGSklGnUM8ik29Jv70fCKviBC//560xSvf4BaesgO3tnNTe+4KPI2ibw3kfNdVJp
Em2YN3W5Wkh4sTXCq8vTqChpbM7XPmA/fakSSkjpLRdkpFunp0ZXlKTf/mLcy+aJvES0ZPq/+M/L
OPJTDxuzWjHK1hYaXcejPdNbhIvmKDAww5GUKekX6x4VU0B7wBMLMTqlml5KPpUqFh8ZWP0rIGn6
lIC223tnqSVoP9vQ/DtviHuoMKh4gINbjygr+pFMTJpmgxGRJag5eKx5wwG9gFotBpyKgxukVct+
6yshZeptVctoIMd/46MBuMWVszGshZA7iPUzHaPN3XVdO3lL6BQ3ElaFhTBJRtz6rp7OA+kFRhTl
KY7UPnItfUTbkbWQVAYgYkTFtL3UCVMOD3k32JzAmFTw+Evph8PWkChhE1Er5a52yKccx0guimaf
1McFlGFUo4VrtTo+epcDWYaEy43d5r8iHl4GR3mOequCcVL5b20r5AwMN6YtI14h9Paza7PfJ7iz
DlUZNR2hjbj8vMRMttWVns9fjqfIoC78MmsD+NsrGlgtWG5gp+8iYmhVyATcn8SzKxCLA5UnRRFK
/IYAcHsKpE9e15J0SjvfdUbU4yhdRPLgHz85SeewdwLcD779KeydISBcNtfCNgURpjjEZt9BhnRd
FtPqsYlFo8ZUCG24SZC3/qr0h01iZPNO5rYBoCiVnmGF1g2kc5ZDtiF8bQ4Sp9nD7bsrvD4ifIWY
6kIWLTiFpIS78BUeHwnrxGa+S40oyDXnNLq/UUMvS0lPQipRofAHTCxTigVWLhtepiH98pU46x6O
/qLUGlGm+d5zErnWMe4oC7ZG5vT5N7pB66cJYneCnrxMjlymJg2Iu9pj1BUVdIGfkB2hNu9RhkvO
0Ub3yFKCAs1ZX0iW5a0xJka3aXnD/q9xV/zOfco7smiUL9ZPcS6rUhvMfC1K5m86tNlBddu9EYKz
HILCOAMfjqTMYXeBVv58RCyToWKpYLjiCoKcq4ifEsxqmCPnz/fqInTluL5U/XCIH9ltUcxZPOXh
YL7Gw4aGZhoc4dnapElWBTOssj61+kg98ZXkxBHAZfuOwlpHatYMfeF7ZzQnmEauC2jE9H9ehjgY
77XWbiEHYrrs8ijYBmU2e5nG3aNk1WiBtvywMX1Ng88tb+R9kzs3VlIBD6rfRQ6pTZQmM1cYRUFV
zBiOIVpmDjDr3f4sDlbBi1H2vtmZkZ76tSkR1t18JDul6CjY0IIk9AE128/d967Iiij03iTtX2RJ
obJpXknZtNxRzM6jriQVaYhskwlNG5RbJWZedwiuri0FZkxqsyqQQOMWlzvzqL4nLoNPSqKLJmM3
F4f6b5SXoGRlNguUq+PwCcV4ZADvctwkew9dqvYCmwUTSSyPawO1S3OdWX2rMPCAQLvE6SQzK36O
pAKztBTnE0n5lnOiTDBT4IGqLUF8nrFBt+Urdi9Ip2WCsVxZIN3zx9tJ/fqAo7wyXwg7WdQHMcxj
OFcg9NXWi6zLhHkjsWhKhae/RWoUGjgDAuPohwXDZT+C8Nh42FdeB+x44fWpzOahakfC+h1hsf2Q
ET4IoHf25pIZ0ZMCpCHgahnwLdOI8CPyZxXekXXoSLM0AXFnxPOPvzB9s+AgV7guKHbe8KRo1raH
peZCTrpYIp2oXDM9STlrFALcW6sEozdIfGBQsC2PdF6jQwdY454EGld7fChqSIDvsNqU1OOpfuQC
CdDyhBBStRet+kkwJnglBTTiXgAUQD9s+HI81x+GzNZhFRgotGaIJmlzV1Iq1O+PmrHuqzcXFil4
EYhjLOWYhSHL7vS8W6E2rCjaE7f9SYU7JXc1SXHIxJ35nl3x0ydG4Z16/med90i73mpIKfD8ft6D
zUW9j9bF2iQn59zfbrtVOndAPCPRHjVGoHPZ0XXesWixlO/Cz++ZPvOLEgeeuS9YJYf7gaS3T+Vs
WB04tMQzE0CjjXKFWXVqnT4JHRtf/DduiSThddgEPKL3sNc1pdi/BEWsdC4FOjhbweYKtnwGwmZN
Phw/fNiXKNEq8RIHgDlzXigdlzqGh0G1+6mcFr356uSDm1pSCW0+8EGoxTsTvPZ7FlHhoLWBjLe9
rZcHym2GriMPsxC30RfeLS19XHJiWQE8F5hi1BgOkoy2KrbRN5BYdELeGFhWH2S/XfzFnaOZk852
HUJuXpAc70+L18uVBP96GrYhQLwHSAtf/p3XQLp2V6UYQZtcohQQdcOFOfvZ3csD2+rrdlsbeTm9
5Cy9BZQfy0b5IfPM1rTbs/MiZcWKhvk7D0mT0y/oRZc9IEgVn5SGZHVx3cJtL5Sa0oxn6MiHWLJU
f6sJw4zEzLdHosvX7HxCiaNCU0Tig8NURVtRo+16Yvv2OG3InmV6fdV4ilBzIHLvoPYP9MZhYAD6
9nWjeUWbvlN6afTiVEmv+yZCg8PvHajzctjZIna3pYY17k5ywmtoET/7idk+vK/OlOWd9eTmF12y
weOcHOKUrCCDP8vz0+3yTZu/nAEI9Y7e8TT5ZNhlgSRj8+MgDzyQdmncx9+QvWiRv4axsQgRhvwA
rbHYXzXzvoiGhYa0GfcNxd8SSl5liCx2I633b3NIRqLPwRvkkcxcRhkjKf8H8YVD4LTWT1/jpHCR
VKqoHIWHJndcoE5J/6/udgJDvY/M+JcztNma0eklDkg3jNC3FYmRN3W1KmpEOcRJpEYViiyCpW9x
3NIeSHnkTZBBDRrO5HQhTxyMpcdgQGxfvrKVLBtgt6jHjoY4dld1h0zgBYCjVSPynAWa4KhjnkcT
FoEvLlJWpDghpzFFrxwu5qxX6Ss3KgeebBjGHCI7217b+IaH79RkBfvsUzs4H0cefladYXE8glog
dmIobML13jR6rZcdzwYQG7Mi802Yq546gRnxcySY+2lHBFa/38xO5fMv/jtSV8gqzGO597lNTAuL
inhCiqei1neeA3zxlFsQz/z3kcFvCFbg+GZYgIuJ1nBg75S+MOeE8g1fspgctnE9CzRFjIGUJ+YK
lM/5798L0gLpbebSr+gPHWVlKtbztqDoWB5+CuGD8Ep+i/25vvrjc62ZNvOB18BntxolRvjyxhDs
leNxH3ASaZdxbs0eBQULrGOwN5hZai/jSJkG4iKuX/HXnwYrS+SGM4Ij6+zD5NgTSkklAQW1p8hw
HOQhMaXTW+vNwVd8uo7O9GO9qXyhccYOF7OvvXBOkk1aApM4YrHA8fj0IuLGNlOaW7ma+jNChZtb
Kgf/Wa1Xl30NsmcRFj49zEoywr4XisuXDO4gWPDCrJamFJc2zkvdltwwlonj+S74zCgfsURmFki0
rI89iV+krZWym21fC8p2Q4vAKVjjhqudI28ku3k8+XRHyACnUycw/L4GmyX0uUUNLrXQ88w3Xsou
o5eXink57C6Q57UFjON+uhxKtdiu5Iff2Nf1RRt0NkNdgiWTZi204VoZObvyr8DJqp/hLRCHVo/E
k9PZQD9wzMegwTzLUwcUWZEwU/HDcZ+ZVHEJ5j/SIPvybrtUkyWFjNQzV5Z9koU9hXFMhJSeWDMz
nTFY38zMpPKuoWNc/RmnZ9PtxYPlTSukbk73Qch/CJyCVcUFEgCs2vNZWxgDHW8x1Mxlwx4wHv0t
ed19fayNwJqTeFvn0TVWmlMJuIW3kU6E+C7yLlFel3rn8OuS9jvzgbQmPDDfiIq2MnRuTuUpaDnt
tIqTISiqqkQcRIYrMnCePDmhqPlGeZexhPk1oXk9uxb47PFSreQDw3itL0LTA9sp9vWHtFRsFlbQ
nBqI1sONVPeavGpRwtowM+Yojz5Uo1QZOp6TtrBCoyTsY6CIRwf55j2VQpviTZT0oNbcldVuhv4p
0Lgg1WMpvEFpVnBPSzH5R2bcMzDTNfnUxrahrTovZIc+U/3U/IpJ3FVhVcLE11zVIXekrB1aB+j7
u4IBQ4VWH8Dlg5DPqDsDemF9G8dI5vNfr/eKhc9Y3gLOt/npzVDX4fTuQqGRT6lOYpF07aFNUQom
cIHVEcLYtbKF2pjxUo742Y/+gZLNp3Ymjpa4shkwN2CYlw4ISmNDD35U43Zg0nh/xjWXHxNSn7fF
sSHRTFLO+Lurgim+BsIYpgijp0HL5F+mmhM6CtWYC4AhAN7oSsQKDcv8XTX3qyl5zDVOoEug2Npz
SlTv+paaJ5tHA9ldaHTO+2BiCtuLaVvWgPjfF7qORjkBmkkU4zoocitdPErogVcVx9oKJBVOZ7j8
XZeF8qdDzsg8Qg93ZtvKJ8auZut45QHUv6Bi8PutAX3G4ERMVkuPAXWEouwR9XXNKPuJ8NlPhgcu
Hs2zLce8n18wZGAGvnS5VohCM4CCr/jh/QJnt4x7Zzzha6P5xCEQfxFBJfZB7Nuazbmk5tMbgl37
eWcsRfsbCSmksvj9C4k/2HCl3cJs7DBMqU2xgrkL4A59ErB1+7OYXR2kdmmWimCcSXg4rOqXmiJB
6LdGkP7od1OHVfAga39uh5O/tBplNiAVju9lyTQFLjKcI3dxCxEOiclkNCux2bFdwI+jktdlfdso
T0/06gDiKFVXlHBA3GLrTXh8pi3plQNABsjqkr54s6HxLEFge0Z1ParuHFLuXFzF4vadd2PJvSUU
7YTEXD51XB/+H/+VNTdeCuecme0y5Y91h9UT/OjQpOdFOQCAtvZF/SPj3W/MFoRx1vxtzdODLyAr
0mHGmWWnPFla/KbtFendylHQ8sH5dQm+uP7eCWwVuPUAhO37DfYLsT3JJDF0BAMtoC0Sjy8ZkKmK
pHmdTqy+MitTMg+NE2hmgDPk20l5n5o7Yh7uXEr1Kap8PgsDuJDz7CF7ZEFe4Sj5YQkDlcO5iQRK
VvuhR7AIwGaGXxsfXR6j1dLQpjQwrxvC0vxHRbWtWPdRLcUNd+gyPT1GGx+Zbmf480ty+GncBx80
GT8uwqZe8nu/KERs9hnaBV4oBuIpeteSiF8B00fVwsakkTgIPXx/5JGDUlAfGVmFf3auFHBdy4iG
b5pB5pC8CRePazOFQQsjaKMwloUXcXafyCKoj2aHz2Ku490qzw7bSnXa4+92GTV3x303BVHGhIFV
3pRDOFfSvPUFzwFOXZOIqaU4sP0NznGfuzewZSURHSrCI8VR0hcWlcWNRB7XTyphThHqBusbNVsZ
RX58yyMI+gx92IYeXcapRwquJ7UOomoYHCAuvIhE0W2TobUqsZvvx34J5J3v05rUpVOyhM+tuZIx
SweTy15UC8MUXCC3RpFbuBHxDUWvApMujc1VOxZELgV9Gw/fVT42FM4ds3T5FCKbc0mGbx50La29
rS6ZeOPLQi6fmlIqoHYurUvictmILBsJXYWYLhOhxSnvGSl1oVfJWD8tesJxGC2oQ3LNmlgQMQ2o
CDY5b6Tc39nxAkDwqMaFCQHACObbWLVcOxKr0LnoLhMf4fFotaG8cWLkI/CIKqQLp1uRWl71QXvc
u2CjybEeVBak3GARyrYWf/nPtntulYdkTQS8a5OlujkLcCp2S99sl+apaEJcaBFNo4rZla86hK8l
TmzkwhOmO5fc3GvsNkf4qw7N1TneerY/Dd4WO6ka6ISoJOe7xgOSXE80IkhU+io48bbhtuiUWUlZ
Ebpi/M4z/mPgxjLAl+2QcePmIhehMa0lV0Mg8BTWuWwNJ/jJ6hoBur5D9efSmSkp4qruv1hL3PFL
tRixfSi1O90xhnDvrhQE5ty1UkKlRoAEtUPyg2WRAttuFtaS+kq6DvpusEQsQVuZAdhQKwjQDjDH
aswhib7sRx04ZW0nDJEyycFI+H7K8j4p8VgpBibGQOX+d+3VZ5MDdwTgCws5JkRMP/r2I9mZIUbb
Xqu2rnogM32rm5c/S2601Aw8AHLBLyzxO3ZMGmfXv4DXG6f8zf8FWaGZitqV5Jd/k4AD5iSBiQYI
4U9vMDR4THIP3RO155gYR7duXbvN89oAEChr847YftiF3r1NjPwAXuiNU8beNZzUr2V7Ow6REVaD
t2WLe+isWgb50B6TI4sh7rcZNBK/+QFbbwrOzEfpzjJv2zSAJ31ZxHPKIKigAstERA1DHq/X+2Zb
qtKzVOyJHOBPEFhSlBwC7ggOIjhvirlO6BYys7n+acsGwj1s+uOL6Fe7qL8HofjdbiEcnYzS3tAg
WfjBHOaz6AINH1X8YoA3J37dSCRHGiB9O0R/S0sUCB9jze1ZxruIoxbpJNm9UfwjRsBwLMBK2PJ5
qhiYreuCtY5shiEL4UC4A8KPWsykRiwXMyMeaXKOTLYMIii5kyCTnfWMyml2y8dJu0Mz0fY2jLLE
K26z3EnrUh1XyWhitHp1yRy/MDd46pb9K1PAjwk2WG074SMzKqfDrqqMW/RqZRAIVq6kYbCR6zZL
NqwWGco0be4/g+YYZVLylzR9ylfk8MDG53EGbQ1aXNtpiH4QEy07QSGKO4J2ekZjw7pKEvM3IziU
d+/eC92sFx2ud/j7sl+KMbzcLPjQe5UkIo8Uk1NCX5Mo5ztcwwrjt39/dn35C2EWKBV0zY5fGRN4
BQHVEZhnAwycUG3fECU/NO+55G+ZKXigct6sO1wArBLuW3lQnaxfsF01i8H2x4939A2Z1WhVcJ3I
crgshfTseDiNZ+CXaRVxAHqYobjfBfpyALxsINV128GCcM9aJM9m60+9+sh9dbIyqmFaAQNdHUq8
il3U6kocV1hWNvR1eD1DSj4KY8G2l0gNvXlgTbZVI4KLRSMTd+6ZE2C/lhYkJetk3BRRdcHU1RzQ
tt+PAJBjReqoEZgONS+rq619TmRqDnRqWjA9MEv7a+pbu2v+w14vHiQWgGhntuvqdeOaYbIYmfV/
SEoW1vlcfq3oyIRrlXvnYFWs5Gaar2fxy0fdp7bjvHFJ/FqswB5Xaqoicy2uRyhftkaEWHGpuNet
O7apdTAJUkkGQs7qoH654TlNpvr50eaHi0nJBvLPk1BuDhhHa6PMO3B/ElGDT2JePud9bZeD3uys
PDFWroqAGgnLCDNgmbIZBwvpjIlcBtvqIryBInXTcJ7hFbD+rGe8cFbHS+CXY7gea0Yqu5vZ5NWN
9a+EIZbWL33CnZ24GRuB6URYX1TKebP8PKcRspgZk3cQnMz8unJ/Agv2cSM5ysz70ezeCDmp68n7
xSJ6bYhE9Wf0Ml6HQqk6mQOn/CajpMG3UCtwXMu0x+i1tmm8PLPblZGkIUaiDLEDMKNrldwUvvFg
6QXxxMD3jI7GTtv6XZXPjNbRyAOkhx/wWhtvqkG1AF2S7bDjXtwhQo+k9KJ3ZgcIQpZbJJu/79BO
o33netxmfULC7aMv2tMVgk6S3eNm5D3wbGj7JLsqoM9SLHoKVPN4gNqnRgEkMc8K6HEO0Y3R5aU4
ozXoAb09IhmGbge+GoZnymKFVfYgd2CwoGwVxuVyx+aYagODKUuNDfMZ1qPZzYYpBmXn/1vDofxw
TMpbsDLJGfjCwKnvPTvOQXyS4vDmMjcrplCTHOXOtKrn7pIPqxNlZr7s/27sNJAdG5K4Aibpp+2P
b/sS2qwAP+G8hOD6nMbD5o7qQgG0cziG6w6011PIENy3G/ZGO7lDQ+MbMMmVgRn1jVap7SS/YC7R
6nkVvZMPASHM0GGmaVW+FybnQ1E7fd/XzDIqyYQo6QNtnGgI5AUguoZYbNObyCAYS+wsWOQ0aSv3
Owqi8rPh6KNM1ley6vvc36t5QK+WmC8IMG3esTc3MvyzdTmWm3SKABQYfiYxD1W3FhY483dANu0Q
ilOs4XrsSmjzcG9WSF3QGBG8wJhkTVky9rcx0Qyt05ViK+uQ582HPeX3hZGgCIFWQ0j0zSR2xcVn
SU/fckOtNnhBVhVUNqjD9T/dfF10ML9eHEyF1663mCWGt0p6k9wEOF+szxPLL8etzM9l2g3vE+2P
qXZVDBl1rXcCIBQNsPVKHuKiL6hgb0iFx1DLQxnukUB6sjx6aCepjD7sK770dPtM+e/gWRXQAVll
DqcmjGfcUbUvZDcZRMfJDfjquR9PiMlQJk8g1HZ54q25nFzYpqIkKPwafduMViEy8CTZkQZmvN3m
02mhD/PsAeSfS81x8OX1sdYswX+I5Vhj1TmnJ3xjjM+k4rPAji66OFKRlVxuSAdUhjFBjFw545fK
CiAeDsvaA55l0plj83wxWk6Z7zjZqouw9j0BefmN9PFKRbBgokzw3HYhyizHrZZ+hNzP4RracSsB
TleuPtK38zk7oUz/NcTTydUuwEcP1XJBXpuErDo8HVbj8CVoprWn94ZrU6SZtv+luJxndeFh+/A6
MOxp6p5KfJtxY8U/QxIrfN4i/q/2CdP8jAGxUc4YsHw8AgrJWvF2oC6Nbct915Dbhs1CArI6HAiQ
ggXsdfrT0emH+z2SiIStN82ezpQs72z5CpPDPmGUuQcrF6o9ZOWdHAdq5AOmWdH1qBSiRehzAizo
JuGkNhQEHnLwTCtKAfGBi0wYMslFTc/xONKn//wqSqKinxzVohGIBXx2UPb2zjKexwE4A5yrvsBe
3tdZTlh+znz1NXVMOBEsacuuMUJ88gRfasILEFacXf8pQKmFekoJN70nNN99q5BBoLUKQl8rERq4
QNu62WPo24tcCMpCsLlDkehP71UotK+65jEqNZqtNS34QL+i49xTkqw5lb9u0LrOFzpd/2B9KnlQ
9/DNZMQEkinwIB8poofoHnQwINQmd9HqXmo0aDAXkcq7CVTUfIOvJUv2OeihBU1lyInvyRNMMdXV
m4SH1TsPXY3dEvrQJ7QvYDh1F5xsY0DYGt2oNKtPkVT+CmQmAvPJ7A5MOTT+guX/iurWKKiXE1uc
KsObiyDHSELLWYK+FCP2I4cJL4j3w5/h8QOIHJ2OapNByhhxARWZ8+mP6MPBInAvjaS65uemA5Mw
ZOCshCJ7zL+qkvPhBmBADp+I/qYsJA64llTgrY424Y4bTcChoo9ApUjbSYBhRoVtxuvpwXhaHiJj
HpFtYtz2vsJErmLXpNDAh1jJ9jWSFS1otadpgmXTPMxbnqabX0yUm8GfN1qu2IVMurukQ801EDRB
JHpjZcGAlp6sxbdhHFSv0+w8x3+EXPZ13uFT4eSPB5vcxJUHwX/MmJKpsaKYjjlYcPN0h7V7b+6n
t/SIxSr1zEqc9kUb6sJE9IXqkFjjqTPai1rWTn4+0d0DSGSR+m5SB8N1eIBlzkhyA7hMmfCyP3GI
TN1ZhM/xht5T+ztOT85VWVJeOi3oEdBIjpTGkTUXS5q4YFD0BVgT5k2pQGa8vtDkuDyMX+pbs4zG
6sqzFRVBdfkymYdOctjkn+3/j3k7IOvdRpSflZlXZ5rIV4kpK0oENjE5b+E3/DPITVzcNCwfufGs
Pj5KZskyW4T0wr+UGQVxcSVC+UbQTU/NNYz48dD+9VAXR7VmIfzfOKooZm/M1Qc+bxloY/fEpI29
7jW0fe7W7RkTuIV3Mku6g/DWVdh+cXva24vQ3l1AsJOddQo2gFaVRl+g4AbaY2868ojQdfU5mmtC
aQFCfW1Btq2rFJ9416IFlldXzUKufRkFd9rexslHQmymwdlVGWC4VoNauM8TvFv0DweVRh02S0Oj
aM19axTedgB7JoFqWnKrKIuyKP0VddW8RqWB/jbEPR8Uhez52D+zjUvZhccDlIsyY+R9b1EsKDDA
83TfnHTzBpdKSF8xhQFua3y5C1yIPzqhP+WisM6rg4efaPqJH5xPajrTO2lU6WVMML+U0BVNmswG
CO2lzl+pNik54RKzaW3wt0DOqpduz8L3YUI2nMHo2FXcGc+IvX0Lt8h1Gn5W2gVUfAP12rNOwS98
jmQy7EjNT+AGJ8h9SWNSzEA8tatr1IfwBcuEVtuoGwRH+wqUa+xmEuieGXb2kWJcvwTBPV3FumVH
iHlJqP+AKNDD6hqHQYzXBH4uDYn+hmMW7BmFdqR8H1cx6MqzWNQvia07ynt0oTJK9ckRz9yEgm6R
aPwGNsiFeU6WGwpuiwwl9Q6QFzvaf7Y83D5E95hVSmzNyxaocFSGaV0exhltPYeow1c84WES/F1f
SrVz0QsD7NRSH8WRdzJrSfK/OZnXBjS8z+ioSkHVz37p7abkgcVwDaMb6LOlGawmyiIiPLKkEfOJ
PSt4u0DKlTZ7966r+KZwlY74KdFgYqZ6xxWHal6JtWh8Gd+kck4hwR+jVczXTA9B7A71FG0rSLF3
BuZ/H1sqtLDroQCzvwqTujXOYFsgUdCyWfwgHb2m/y555BPqmUWzg7NJ4y1yyuqDbI8CFB9kCVzj
OXDcps2P2n7ktPzK3gFJRT2kO8kAj96rSZVpDTpwwCWPMeHfIhCno4Bt1o0kQxV0nGyJMDW/0GI4
yh9uU2NYKaYXevWy4p+I+N+RuS3w8UquAIsk3rhIo/P5c8tjHUQiOaymW+Og35YZ5JIz0yHAgccC
hG12SyeBNfonql0qeUwWYskkIqR5b5sO6Y2TW8tgIobMyhTRcpgEVYIP1OH6/YZ8spnf8l7Cc2VN
9sGwwDicdo8qw5T5p4u9rstqZs1FBfroy79P+tsNsatUQ8GnLYJ7AmyZ/Hk/tk4iN76lXwVXhV0Z
d/d3wY33gx7ZIMLMRb1iWPfsXMnPas5VAZQ53rBsX8tDQVSIGcwvi6hAHzkzMvPT8f7fjxmzPz7G
U/ISmYaNprj0HgD+AAGAY7RbwJO6OfS/G0g+k8UbuTKLmd3hhVEwHL+HfNQAwmkZbUzZ19t1EvxF
kBEVgK/aYbMRbUuGRZaodHQlvGUAPdHUA5c+vVjldtWJFcns1N5ZSOhVlG84j/kyaJybNEBtTHvI
nCigo3+W3hoQPaOJZ7FNsjcmmUEkwEpcLCWZuVJtDvVWLILXd0HBV5UqygJtOZJbwdFSVN2idocH
482QQZO4TJmrWbdu1rDHxMeeVT9aF15LBRHnU2Xunu1hCWizW/rcw19i/qV4pl7tjj9tiMJy5t6/
NqI4YJEWzQKy6RnFV1bOrJST6Thsda/FsbYsGcU7SU0ORc+uNNYHYI3Lpm5lpuNey2nIgwbCrbTg
KmJUcrZdZESea9rWhFVMAHGFmsKILQ5LSPTkzRH3u1zgF7R5wbmnsP+8okWURVdq0RSQx+xOse6b
T97+Xp8Z5UGCQV9B7bway836cwnCWBAN8CQAl3ZQIowAC9iVtyGicaM1Z2Biet+j5Wrl9n/jIJwC
0i3kLUkl72MFXPkJ2VSuNqnnBttw8GY5vwOt1MgH1Kf2tCquJ9aMfkbHABo3sUtUspeg0uOWXetY
WX7qc1PCETGbZHCqlqcRtSe9g9GEko6DTVKmNGcvE71UiYKgbmEwL88wdT1RwiT49sj4LpA8sjYO
RTjCCdaQne6bXNbUzo/97CNdEIVh9fCpLkELs38G7MXUfo+UmOqiiKWsbRCClAGV4L6j9gP4QcKh
UZaulj0FW/482FXhUguFk2b6G8SQ3gQGlvut74BE8v0XsOwITytkz6b0ZOduRJ5vlXXYaJW8A9kK
gBxQGgQcIOKjlK0qc00yC2VL33JQ2cfsa5YEj9wFSf5tfo3m3Cwws5oFax0gkcGUhMF8EEYZDeai
49AWBhy7psvGLS5OTthEZhcv+ihweusvwMnNDqwdLkfCmpIewDJivHKFZhQ5s10wi8Ivs99FWTA8
AWzEzhgnfui/SS/lpXyQBHS0Im2pNseY3x6fA8WOBGDctFFGH0JjwkLeOylVnCxjH8dUZ6bSjivy
NyAIiVaFgcQkQWM0V3jFQbedzeAgj0IRRaZvNwPPnimqW8B6/lNlwLiX3BIzybrdrVK/5B+jmRNR
V66gSycW3wU1LhAgNdRXva53fZtWnAbD9y53kEzHNjLlUYuthVzG82F1isgNkTsXxFoJwJw9xuha
wsPMlXZIdpE//nMSe66JZRpfkVyASwpw9XKd8CSJGMPYILLA3GT+KPAzGzJbkFu8DeKDHsI7UrFJ
4U8TZvLC9dqkxSuHYOiJTH8ZYL5IOrrweYYuF58IruXPCEZNxbuBgaD5Vvhk5pGdjT9+fwsVqFgZ
ZQfMgbC8lIS3XW2pxD8ljhpEn3+sjTN8NCusaZ8yLwPPxaefSAp0qVdXnDoKEH2B2gn7Ea/Zq11a
ohZIj0+EZW56KmQCoCGUiwHWW0MyCMPaa3N+8BLMgJT+IVWIyycG5rE/nV0+ASNi49kJcqiVTYpH
tatVL8av8YpoFuwvrgT6SWNWRCfpio/R/Cre5H6SHZuMtcUs3ukj420cMCOSYtYZSflJQxtn6IBl
jUf7Rcg95rPT3jchrRex8fSoOmzuwQ4JhJt+G0TUAsZSgZHBThwY7d9Qg2/FErUwZmWT3mU3ZNH6
/TTrPvBE4D6kAa2Ac0t+ii0RsBUJGc3UKQIwePbEV27EV7Ygb/iC+TeSBHIRvMCVlnRwO2nbuv8O
jAtqbx+OTO/LZ0EKdZ6QbT2GQcotYWfbyzxP6akjHSLIbjJw99wzrFlDDOZJ4drBjn/QBgEf5BA8
Ivt+XqWgHmtDEn3qOOieSyy8B1NYXqYvNN9abRuhbVFNbbkS7rm6hNEUQVe0D25rsHwaxRKwAwKU
gDLPHpoIFtWteUpwnoIahNnt6SqNGfTmaJQo/mrSf52gVf7YJohPxSt+yIvuF2eCQ1jBqxafll8G
vcRPZgcyqzzDDwhPoiJyWZdiL4MkeWLnHzYys7WBJlFE5UpwoXhW+JNSPCm1O5S0L4K6GTZMZtnn
uWd/8JuYUqKJnHmFABCqDC7GVGPtrBbBC0/QRkJcRAafTMIUjaGt9XoLZqt1PrHL9EEGkDBOKG7J
9fcXuYhIfET3YnG64k4alRsvjRGFv59HL1nrpj+L43tqoxoVz+sXiyggOXBq4ZahH3zu8gfLOrHK
WWCz+nlqD99ZyDz+OouQZxOFV6J25Q/PUp4hX4L9+iomQDmx749gh9peT3bfB32VOQBJb0hsEs8/
020yFfJvt9OfjxAKSbvyattP3kkYQqFX+j1lrvfcnRLfkJfoPJyuLZLMeOzAVd4j4jgJuDWprcBo
Vw2UeoKkxSYGgCaUQkwRT/cKoBkQDXMo4rFz/SYIIHkBv3kbh3JnjSGzg6SlOVRuzfc93Ntm56xs
xxRm0Br5k/n0Ea3YzDdAIP6bc5yWJtRM1SKACVaTE/OI/kuMe0PVxSpPuNLjvnUbK7VsByBhf0LQ
/x8n2PTOzdzXdafu+gQkdqVOEsGA2LIngsvZoXWPMMd/+Ltw45riSRi5VtcIUx4FgAu+x/FOkDmu
COywDfpkNQym4z3u2wVJXghz8k04j8gduJW1dOyi7337bSt8/njeSN83kNSJU2zXGvmDoSGRCsmY
QGBB5pdggDlsqLEwL/9lOs/mbrXMDSkv4Uh2oUItAiA0HY8IeXDRm6hND9SSBxJuAn+48D0TQhOx
tEMCu164oZ4YUhqLAi6wDNds4hWgFx6uGSKwfss4JEiS1ttjDoL/AY2L/NIYmxbMDww9qaYIBOyL
7dUk4Id32IlQ1McUSw/VG4SE3KFmVQUWYdOFvq0nXdEXBkRoIT8Qh1qUeh+U4FYdSqLRvSC3i0Um
apebE5WT17/wcurX8UIG/w3Fe5vxQnPjwq5fsV8Ya4ImEYD+CrtUcDyB/OBqVozsU7vfz6hLXzKE
BGOmQQ7I0nix6tISuKOw+7zLJlD+CCJEzVKvuOWp3n5YqjLqga00jyj/YIQhSSD1BXEi1tLMKgaF
p1mHAr0GqcAgeDvxikZTcfx6Bzi4D0y3sm2thUaffxLRgZYSGrJU6v7zi/t04b6plvKaFsioVhnK
50Ccf9IzHJnDNBkXNoxSISJsEatiDj7pcf0t2nPKHoGigaTLeBe/OSAeazvT2VkfatySdYPXWNGx
mEyYVgcfUn+jeoYzPGvFm4xi5z1bqpeuWoQ9Jjs319w34nnrhGwSTX/WiX1Z/WCQbFLHpjOAaRq3
HGzJ2BQJVaTuIhM3aR+J7uiP7TjjZ4sbR4y8YU/0Ic7eNoMGEZkEazyhx4NpKlWmcF2jHJq1bVnK
58yz8Xt8+qp36WSjn1+DADPNE/Z4mTQ15K+Hbo18IdNZ6WbnOCVdSyY3CEAL84PENVlAgMvkVNyU
8bV5NhXV3vdJlUN7Vgsdm4Edstu2+elQKjp6Czm4znjdkb+lv4YEDCRVOTqzDYUkm+LoLOHAbJKv
NLPy6Fz3RavLkyfnOQyNyXMOz57GVR725pEnzu/vF2rQ/fhs+7Uyt7iIqJgKB0KUdy8OBPbEKZaO
R1bf6eWx8M/IQYOtdlHkZiNnPp4i88da1xVtL8ZdHr3S0yMNR8BobS6XhTbt334T35ve/gKrxn82
Ky94WPTklGwNOngjd3VixPsrke8MRWrjWpWHe6DS+EFPhRAjUeJjiYqV3S0tfgkRNP8vKgfbTQP5
YXV4BKdlfOApUzH3mTVDYSYW8QddkKByzcI+S9DurPvxuS2o755dytT2szOe74LI0qBlwOqrJMd7
uptVGlvBlhtV8Vjkt/jjOgSRNw+IXi7RPmpucrfGzeYhJNqnq28M1VXiz/A3Co6wS8+a/qPOg2Bm
e3cK82/qsdSihYXY9bT7hz49w7i1usAxSBh6y/vyY3voPy1teb1cOjOJh4q/dZRaRB+t03jQi69l
MQF2rh+i+5SI557v5+VPXTU+oRKgIEPoMJqB/KY9bhuDZmobfaj6J3QfxDLTuSJ576hNHoM4kT+n
JULAKjsy94eYZMDOuXxnf1omhOavLx2y9xziq9ED0WhViua1WwjVBJo+MzJQNrY1PUo5uv+kLEFh
enZApzNBPpORl9LvZM5el1urBCZPj08TarBJ7TK/IfliRji7sDSx0X/RCnKR5+u8+SdLAyJApx8j
jBK0/71FT2rM0B8ZHbp5bNRAPLCXhSHvvjcINbWxVakoPUK6NAy/JRTnsT0j+kJc17GtUJxn2ICR
Xi5flLItiWF8JocnPT2rdoNea9x4tstB7UBlOBiWHKh5v0/CVcAK9nuzlRnbit5EjgmMGnmAvgZy
rlvdZXf3uVbgj2CDneNpJ8NOIChmDH9jbl3rhFDAakwp0oSVlXlReDmgF7qgBAcbsvNxf3o1bv++
Qig/MtmZLt9Ns+voztQ6NEZNMVh4mdzMOJUV9KPNQtCnHzT5OYFKVYVvLlP1ZpLcLjCaxrdkhXbS
I440Ag33Ko6fGf0aOHztIaz4GuGwW1vyqEM0T5FF+xS2x77cn0MDOsqgRHsaxT/6LWfzFEg7rRCR
jm599AGMq18UlRgzOUAzoP3UYBCMtT9O2+HmxXi8TZIM67LgppesLYrLl53KzWSWdmxGuLm66AAL
8uIJtjoqAg6q9wRnd4HDCdst0pEtbQdcw31VJ+Lg0PB4QfRnt4ZawX0Cayhccqi90ZVv5ln3NkFj
dZV7Xcky8aD04s9FYKm2UWbE0BhdAe7Q4T5dgJEVDM6gn7cpAPXgL3XXo+ePCzZL1MGH1gMZfgQI
XbPDUEa0M1ftdu/v6Z8ZWpdPUW9cFwern4sdEvfS9mhAPJ4xCvyJdGx0KNbhY0nYL4amv5ui8t59
fd6mXeflShWhtONwAK556UZsQj/U4/HGUtafU989jAbfwnrzl5p5ycig4EOn9wBs4++2MIh3sCuC
lWlRpSEnZHsr1cxxL2CNyqGEQDVAVnhLihGVRJjOlwusPEDMFce3OG6OA/Nyiz+uvHLfqYr+Oi2J
xDOWSTcjXK0mnoBRr+0fF/XjpRhvS2OuxHi7t0kXosLIT1yT8WocxVSfiQ62DJ27HeOk1XE88cLQ
FRd4dT+dkRleyEGiJ6fzHvlGUIGq85ZrSc5fUDzLhTmH0VwBdwURKUuLFh0qDLm9dKDd9mekkWB4
lQMgElRwrbOsdD+u+9I6DYgryrngwzOzZv8rj8bJONb8anLm1QVCQMBPoCRX4BBw5OM2vYtkrpzR
5uOjq+soVrjhwKj1/MDDMvE7YtvMp9r47ibKBFdoVExqzsQACdx20gKTgW8s1Gsk6U9q/0CvrfCK
hTe9U+gpS2fu7339TLzg7/nOiAmsoJ5ff87wRWorIT07GWCBB+Cjt6FE6MefSRPk7B0IYwaDpHeO
asexrdfSXgha+xqnQwixrxpPNMJUu89OLkf+pimuchulmgSNuqokuu2CNcRphuplWWhTcAF6pEfQ
goe+L8RqE3Gu992rD+4O1pM8204huP0+N0Z9plHspgMYhf23pNosq7/hw7YYKD0dXHnE4hWg1kKH
8DBUAi4Yrb+TaMh/9AUoygkxsBnCsMDp63xr7cHClLqJrQ9xkw4rwzIeMCRF/sPDFFGVdRS/eFsB
0M2vpYt1XNfc+f5rKblChfPxlm9XhlJJPOtPg4CcdQQxtG5t2WRwvdDEDW2e5cdsUid3IqdujdBf
9y877/oYkzY460Emlp9IANzSys9MMF1KmCP1dBX/W/sB7hCEpPV1lS6D9HFv/Zv9yW8wTyyW781d
DWerUMFWsKyB6cJ7oCIV2tBjK+ZXDNJpqNsc/Sw84FSIMcGNRE3z61V1Vd3+9Nj63PIcFdl+ZvjK
NexRTuAgFDU9Qh/CE76KsEK3d6lVw7lpva7bJL1g9MqX8uZj5LwwyEKVQFMbABZv2RUyRslMiDsK
OEPSQt/IjlgrGowppzjXKJ2fnCOJWI8JPpVUyRohQmEUUaBLT102kr7ot3RsSk13OeIdl5nWsxZy
PSUgZ+X5E0UNE5aY0NfniF6PD3D6XOZ0bZMIAMJH8zCpLgt4GTJL/n/omBXWy24Neo/WXF3a6c0w
QbvCUoDlzNxj+M4gRIlNiRV0t5/S7yhHwZjMjao2kQhlPhyaiO83kkoFM94sDXRQ1iYTnCfKP4lI
3RY1txsQ/IFll8gTsmkKbryP0m6K2XN00Hy3fOeU7gXbgSc0hqogc+voOQ5iPXHZG117gOKi8gw7
BwoDh0QUfF8LqkHU3T0BjxoN4J+KcOFD0AwtGHT9zAX8ypjtAD3KryrxdSRhTvxehM5BSWllbGuI
4+IAzGS8P8XiV3OtP/Fcr9u8G99Ekd0GUhjSKjC46MAAgiuq5ojgkeOaiTU0C9MuztISvil+OZhB
ZeofpV+X2ViBdJ6Es3oOZJFFbtiufofsvjUY7sUZNcrrVwSBkz9g1u20QVD+KiRVf19FC9yKh0QG
S8VHgNZ3f6nMNS4BWeiCn0z9djxV8CbnhMFlclRzKo8c7/rxgwMk2ac8UgaMsah4rG/59qV8BqMp
g1pXilfT3WkMly3I+N4+5Ao28K2qtiQ7khHUZTd3CmggNItsehqC3mEPRapPm8dVcr+V5efnRS6J
H21Hw7Lkycyhqt5wwqEJVB6bMOnHnOcaXzGwUvkletBTQoMIfmSVF7wMepSqrHho94omxfogtYJ/
TNUQvnwzg2fwDFroI1D+aEJ4YJlSodPUBQreghT5u+lYBWnb+gA5TOX/68+zzc4nf6gqyukKUTSQ
I1KkgCIBSfekjLtRjdcBmS8etWjf9piIMhcGmGj/oGZUWnDVTAY8DF14lweGzRB7FlcEQvKNPUWS
EYxA+eE5CoSrkEhGW+KuqYd2dTjfzhmNARz0C2RehKMHJnqkTQseqOtDvh8+NZkfy4ghw71ODCVT
ISledhbn6Mn+RmM2HGdog43AVy3PWgI8HcHd7uxkSzdwPe0saPj9qZ8PJFmiNk+8uJSKYdLQ2I+6
Qm+JhndTEceR8uVIUks/pSnKPkeEPg8p8g2sR4l6JvO7YPyhJa+4qiehwGAgIhdmF8YrlOpFfzHc
EU/z/P4RH1Y/kPwUrggg9nrP/G5q2v9kbolD88Z3yl+BS1B781mI4HwkJACO2MBpeb7hieg5XraF
+Ka4qyHAqJxAR0xKa30Dtchs/PCaOcSKWOPNQxcmfPc0B6T5g87I1BDdtiXQuJGswMRd01cIhieb
kv/V8DD91MhBFlDXRs+niqyTgYMlla3a5YRrU/AQETsXRwgGlzJdS92DeEQalrIGZVpY2cvR8EYH
qnL4Ytk2XdbO0onqXCenVoaqMsT69UN29cokKV1O+il5tFJuRxZSWHMwuRgxrKyZOd8Nt/qrXM0R
xtHX94GdlNMPUDP0uptpFETwkc5XM+hRiVvHtXTmGPz/Tmlq5BzgAzoGn5Mm7UXSD75KQbk+/8GA
jFYKH7uZsII8w7txFiSbY6KMOeBSFy7dw7wZ32JXPQKgm9NcZl0SYzWdcBGXpCqzAsKsBPZMnNx0
AVmS11XQ6HOjFSVYBKcPL+84gL/jd+25mUB+rbvvlZKh7/ytt3faADsjgsqmwMCN2+CdqTH121RP
g7XSTPmo8yxl2eu68HmOD4ijgq/aVN730YBlPqszb7NaNI95BMILSf60hzA7xduuhF1g/LlIzBiS
OXLE9wlKxUGiLYEEEc9ieihXBTojyWZH6aArOg+NbmrI4R6F6aecdnXTR4D0+JY3JNdjGY1Q1A0I
yHZvvKtjitophcnZkBV9BWH1gq2Pui4o78l27md7/XvnH71wAXi/Rzfdu5u5F5seRJwU9NTlNn7W
pG/HLj9bfb7R6PSCqGRSZGrREdViJkzD2aYDFxYWu0GWsfxO6jsOBBaEFI8wsiIbKpL+9NY2xsam
oZ56/0V+wJQI8yLU+Ty9r45ovb5OYMfmwzqh7zB6OsbmtTkRX0oCyAsYqyssCxJc+e0pLyKtAA2d
qNMbovGwsgwrMKyIsBnmox+qoUWxUqVyvvTh4SWFb7Xnv2fcsi+vXie5qPPUdhReB/oZmMqQ24K5
YUEC6BmN+/g03xwSjhvEbs3QKoEeV9Sw9yepMQytyGs3XlVvHHCcxNrhfPB3PI3RcxDBtWtOF3A7
5Woyehzqsw1o/Q1bzOIbPmAaAOzklKO8CtYn4JZ7I07/ZKZkv9WYAKGdKL3rzoJZbpfBzRSTmc2p
ZnYafOENk6zKUYvUkyrIj0yz+YXIVD8Imw3OBtXQ78C7VR6PefPBOoTQe1itv426+gKjCiAXz71D
01TE5HLSwS3kI5lqAsu7IlUyKhHyuDUhdyhirMD/fhcUo5NFTNlzXdyiWpe5ygpHTn9/Xc76OFIH
Rh3DdrSEgE/thFL7AnYG/th2F5WM+jLxWP0i+gfcBzKcGJ9RXJMz01kWrLQGLj7olZ+u433BgMxM
6HLC6vZaY20BKOHR6qZi2maw3yT44QVPKUEdk8uRvt3KNz5KFyakgMRAjjxYXZT9bqjT0Jb51O9w
YTvPAtMMJsWlL81dY5bRduv0PyEGWxwW9a3LqxViZlXiF/WimO7eyvURNYPy4spJxql1mmCYvUka
TfytnXVOLEOiVCwSPE0L5uzpz9pbC/qh9U1UwTHIb4SsQljwZl/ZVzY6RnN2wFNbsuLfw3CT7LxS
AFGxOK6fJgwLtO+/zrlSlHNIkXqI6041QkjbKmF5kQSXIElW7Dfm55xQR4dJ3WHb1HaKXs+NdkFV
wpy7nRZ1tWPOdcvwyvRYBbFWfe/DMLvaBizudxI9GAb/qbuI2YO9tj/68o4IUAdVhSyoo4piOHw0
0BTLPfm7nXn4b/nv/OU7DR6tbSjtOzo4rAuVEPp8qsLJR+3l7DvCBv5YBBbqcljaK6fHXkFGab+1
rMmmgr2c19bA4KT/yIaMlE0s99zrD4mavMx+upZQb4HwYMDLsKYGksviMNRiiKVtV7UN7Hq4YsqA
6GVa+/9qSwsehC5/4QFLKGZ7J/Ctu2ETQ5S2RJWo2BGdGmcr5Kzspc7d4Y/wMPx8WhbaAlMKBgVT
pNXJLq4ajZ9l1YCEGYcddy4K/PyYZW06PS9XysmsbdX3sqJoWNq2xCUlXTALIuTuTYQidcgMnhqo
RuwYEXk5cuZlTr2XcxSv9+uxKTau0EMoKCdbIhiAf9kyJFE1RkfhyEy0gMO2edio5mshsQmRS6la
caA/I5gGMAbT4j+8AphbIeO1pm8IajvpHXX4jygAzIPPi2SM2XfL5GHmBH4QWfwh8jKubfmUy5m0
eE5Llq+l/5jsBgo3OX9JkzPgmKgwbytptYKUxmvatF+DIbGwJ6MV/se0GDLnHUOux999uj7OUYI6
bAZ9Mpx6avPzrgFLrZZGh4+e4WRRg3TbUIaYJC5stFXJpruuhejnS1V6rK9XL6eRmHu8br9LJqT3
wLBMMGxOtmq9N/gD+ntlLJSRxiMWRIp8qfoiD86yus2kfm6htMbxAq/70M+jAeiZyjQNCkUeWpRC
HurHQUgs2uHPAG5j8cvDeDaY3w3s4oWp/ZzWsg8AwKzMB80uSdmluTHvOAderIeO2j6vqf5s68Ei
3jQUZr1rBhDD0eeZ9PzbJTgG+YcD3ina6ut5rnlYqdkwG45tSvkTBM3LzBZL0tPen7q9/v+7J85U
Mv1hOWZ5GjFVhyw4st8nIW3BI9nSrfM11H+z2uEfmqlaCUlOgATKveO1LZJ4P+8fL9IXGU+pisiy
agJI94UZjhJye6L2W23T7t6xKQ/aQGEloPYRZ8U9DH1IlQ3JAWosjyf27Dxkcma9f4hzaDVEl4EB
moAtdA6MN29sx0tDPcxWk8pU/72Yd+nSpTE7qXVzH3hg/YopLArp2NH/UOvQcX57VXUO/idv1pkn
+6nwTLhjReC17TuY0Wdc1jadS+VjVZGavlQlgo6J8jN7aSjU+HcbyGxzbMl6RYRAAZLvQm3WMZYE
xdijY54ZC/pqZgoKrcuMvLVfwdjsvyDCcLaFT+rvymw2HV2XIfP/GFQH5wHBBZKkUYECR3ZzDYFB
lIcgnbOJ/wZTT0i3M4rKp+w/km7bAiLj2tvke/qIq7RRdPtS1c9O88myuUJa4/2AaikyhpX+D9WY
DPab1FCfdVC4mCowxItzZS0TcNrpaUfNqdFPdR/ieIpbrE6qhLy43hu0lD1XGfJtJjziMVPWiUUq
kpFjlpWc5bm7V7nD4LQqLh1hUGeWHyk6MjWDXLoczQcIoP4WJ6ibi+O8wLzqOF3aBLQDc22YX2AS
JPNs4Grfu8Ur/IAALsO4khLfgkgUTJ7cX8HkKa2r/uRGa5Nl4p3ewVSH0u3XM9hCkH2fKcSkh1xd
FM4NYXYZ2uuCVj5TeRIwpVi+UpmPk8zLj6G5tag4L/TPQWdEYFcfByNXnwKXl14NBUxbteVb67bq
dklr51I2gbxAybxFqFLSJMdHuKMgF7b8rIVRl3NWHg3gyM3DDfXnt5xVCWi0tmdi8m73rUb/T6r+
6V+WrX5jZWpspyxDWmTzVmwnFFlfaYq+0WrP1ucNLbbXhDjSFFgsa7GOGmzns3emdkaNIgtRtoFr
pGHAorKpZHgBWFigq2mjXkZRxMmWsiijxSQmR4nE3DbrFmQtXU+aSzb3e23dEpfdnDg11XYrOk75
JvdXc6xaA84JUUPb7+3zDDj5RodahIGW8yI+3cIR92KI34CDtndBTTxi0KqztFBEt2WxnW+DtJBT
K/5mg9GTUASwgnuGMcWx/OXRODtJVwOrOvGrDnCo02o3B5ldH2DLQX2sChHr/czWmRZbJryYxzPB
xCpSCkjylbfvPgJc6esqpzPpLinByk/tPWvyo7byiufZEzNCY9wPo0iV92CNzSSHd+qF7Wtqv1n/
n0P765BVg4khGm6ZgRDuRLvAPq0LbQOXt7sAjYKXftBWv2lDXGv5ggacWeDTR96r9PrpR4vd5yX8
JTKwZsTzF6bZuhebRwqL3Bj5p0yf8U5s0naG3GZlLHYq5qyxxelcfF/CrrieP6UBO/CrqM6FXKR2
gku94v8LVod37L+IbgCL4PNSOMdZd/Dsq4gFqk6DoWFXlBOqQ1SrmTR2my89QzEdYwzmkL++xAmN
MDiMUSId+sSzeqSK/Wz5Q5e8qubUZB3cGDzsJands0Gc+p/sZ21VqRAfVaMVZdYVaWPUS7npdjGR
ZOwsOue1pdtT//k6qJ5bsh2xW+cXNIDNQ8p/c6GNpocf8+n+TTD/xO8qfe6EKzv1gPPnS8oL1YBi
7gkpU4Km9FLXQABmpDkWjydBX2OmXRy0diWHTLpH4lK03/CFaWvYRzT3pm9AIUNRMuwfUBY5STuf
6hRzET967mPaEuGBsL7VmiB5p8958q2e/D+ObN2o1MLb6wYn8YK1TmXDP5tQS0u+cyPDQLsQ1+UT
p99b+BAC3shk8JrD7ghMLDwzQ3kXllGZOVHYxfnpB2YZ4wwW2QzAf/vRr/X+h9vWd0ULDwx0tdV9
MeqQFc69wsNJLvHlp3h3572b6snl96iBlZXdz5NmCKh27PW5WU3Q1vYAIeSIGeND5RLg5wufJcnF
nwPQSYBMWzcic8H8E00fwUd5fLzH74veKABpDSfDO32FKJ8FbVUnSkzu3WE/+6tL41h4mQ3kJ/vd
O/MQVLpzWZ3SCdNDZAvUDVcO/BGROwOF+c0KA3mwbOdS9Co/mYvmeujFtP89H3ktZZuV6AtI7Nrw
VwIg/qBw29bsjnOrjGqT0GqBfeAgFXvzEzlMa1qpx6egSNQmMBpeddpwB4myQ4PlFbF+yZ+AetXh
vQKWxi8v2HL3q3+GM/Fkdn5iTE08+MnMHBqnskmFZ4gwKl5CEeFKlaNHLp6c2H7yWtMKhdORRAWg
0I1CEjCdUHCwK47zJ9HoZ7XWv+P55jfUKiggB8dGW/924JOv9KcT/oTMH7l8U3PtyF/GC7kI0Vr0
3G+3ZBdxjbeRexj4WtlTTFpXT2xLvvbUGy/Lcz3sDdhx8jdc/6+vbZOfHgCNdzQdjPHp2Tz4mDbQ
wGJvzrh+J3qWXb9Vuw4etqCx3iSuS1bb0SRLiNTYO3KI1CySJvQ/7/9ZtiQzvgxcylL9bR8OHkoN
RZGvrm1itP1/As+t2g+qT6SBc19CNIbmPbwTHvpMqSY1uUgAHHG9Z4q7JCuYvuNWPO95c4gDVjNw
m02dwRQhdw8Cziv1cyhauk+p2eJz16KGzLNvjARabKN6XKZlAcUQKr8z1He1bEvZgW26yleFadkN
9tcsd8MEIFwKSB18qWS0PWftDU7yad7igW/hQWl9A5YMBTCe4dn7Za9M6LI5Aj3dScYVingtVv3z
bRn+sUoV7Tww7SHJApcGPN0Qad5+TOVPYkqvJBg+5mSHcY/v3A6rq+DFAsjzPXxXvMcNhjZuX19I
HiQHb8mzMZzk356Jh3XzAZ5et7zaRK7DQLpo8KXzUGHQvnFqI3TBzE00QqraxM0gn04JpzYveUs0
HfjchsS/ivz82Ox5PXpdeMmJU43+1AWscg3P6VtMI7Orv6K/yDiyKa+KrQEOLyRuXCP/63wQCh8R
aH7usPDmbyr56kvHKSSqHQcFNUQ0+rLScEAONdYP+NkFeBWrzO0UUddd29X4xdDS9/D1zFLlYybB
q5xeUYZzEZEKbsnsXjM6u1g2g6qgx+Sgw4U7b9iEc9p46KbSPAIcSi1z94GEFakdMJ6fvIJ1mFT1
roADaf5EbCeCkuh1rRCGd+QnGNTKPbv7KFGeZ0SsuBoCiTaGAiyR5aMdp55UDVCREEr9leKUkYmW
hevcArsloKc2O39tJofDRZDtTdmGUqBK2ZD+GmqQgv7dy5QmVyJxg0xpWtmLvm7TahZbY+4WgV3j
87Ck4+NL4YvtraqZ0Pazta1wm7ogz5UTyX55falWnpTNGansTW/cG+zI9Liy5Ks02QAK7498cWjC
SbZ8lZXoz5KlrIuG17doXZSmv6FS+8pOku2Fq18qnaWL9FONu9sCSQxT3yktkrTvZ27i4wlc7KDp
XMss/8jCmafBxyD/xcASRIULY8osv84DCKUXjE09zZAB1gj7PQVoibu4QcCejvhuuaIr04M10qyW
VgUmA0ChTzkts+ZlMvUCO9PzBqOeUJMpeaubbdg4sNDUETgEpnzdiwcWq7Y7E76bo51ks9UfEjZE
7ejnZen9TEpdp4aOr1Bu5+fA3zrlNU+fiq0jyfxrUPthxWeBgWBC93zbyL+K/UBAsRBZwKOIkciG
A0A2SguJ0GOqXamTW3REaDEdmH6/LTcity3EjrdlCyMq6uhirMWv6jGBEQf2pEmHorsbHcS2CUpk
xNPNqtcmE9SJuSBVm3ky8+CJXSMbwDdBQtG2UXBTgV268D/25yB4FAWuSd/h0h5XFO5I6nRz5KYq
NavOVGeUXqqTh6i6oFIN2mTLL5m5Om37zxuyBFmTwD9l53pf9Oq7RaPLnPH3fMiIPwnE9l51yhdN
ixWSV8SQJH1Z1sGXiV9OG7Rf5h9JWMCqhIQ8C0ue9uQwQdBa5YOyGGJ2p+h5xKqQexBSEzJAoai8
sdCzln5FYl0nxOsjbRL8iy8gBICgnbPcy3gYuA4EZ503U7NWydmzvEK/f5FWG8SoJkVDI7q1CnLz
rRz7/51mCzwMpCpHrlZdExgwJu27ayXebdbXo9yBlMqjEj/tkk272UqiyjO4y1Ny7ad534yr4JwS
M//kOXb1IIOuhJQ+/4TKBW7tt+GEOobAPL97EpCjI4e/8/mq0N/BM4cpX/w+Mn+i0hnNT8nqqBz6
ixJgsgbw0r8biWM1pqkPb5ePVQmatb0+fSpJq8tLr9JjMlBQ2dFToA5uuCstOpUdRA3OMCs9cGOY
tT2xsmg61aOvOhjZul9vrTQ67U7t55l38IleVZvMCbKo7Z63A2QpqLDLBD2azaBJSvd7M9fkWULC
BVcAlXjYbjoloH2179aYSzOI+D0KxokDqG7npQ4cRPBvRXlFULUvdZuovwCT+aw4MxghO2gWbMHU
QZdlDGiF9ABvS1dl0XwQPztNtMLW/fKHp6gD6CL7SBPt4hmwQDIG/ebUT8+ZUk7lwjVVTE5dkoN+
PLCO/bIFjgKRIRQ/jNR48gxdq2cwCmsFrSsrd01ygkmiTGv96VEfRpia8P/EuxCCZx+ubMZAedQf
F12uGw82c2F2+kTKwvaykgXj9aIt7C4z6qqjk3Oo9JWi2strYo3Wmge2A/x27zEjQTAn1DyRFohx
ntcByLCBIcEYdBq+durPjlaEiOll5AvyWLxuIUAzmCkzvkgXXpU96mgMc5Noh9T+BvuwVfbXTbCb
quinNPQO3cUTTXdYP2NnlgdO8nbMWvQNiDqarMg/i+cnJewmZsOkWGB/yLpiq41+e1O9M3lPH5n4
+JXVvHN481LRe/jX2EK/+AYbp0IpMx/o7MKrdqIROzTIFWhb6mncYM7/D76/jFyYWcxmwSCa8mSR
5n16FXcpV6SXZAcwsMjt3cDqcZr4QwRGTquwBKnf26oklnIRLdEpozFwsrzyuUxBppQPO411PIc1
BH9lNnydL0dbXtwbVgxszmsn79Q/ANKz2vmZpRG63Nc+S7wyxBso0b4MXaik4AX9TtbJyE+WG1sp
lTj8YGWi+dpx2w0Po6cCUtjXL1baAOserHq1AWWt90uULCpWizGBivC+84jYnm7SwKmsB5YmNHjC
nNo7vtezXeTzpHTBhDnVhntZuooi6kDWErtKD7Uc1KhFO3JSsQAYslNWXANbiwPELg42Kgw2My4K
WDO0IETFzqYNP3btODet5c9SrF32PiYe2nRZLsyMlkciMIYz75FQQxTtoat7EZVfBqYsPNOFhT0f
zRD8dox88N1IgKPgeE5CmK00x9JF51UDc9b0vLDi0miiAGoKzWaOQ4gsK1StikADPFaznq6EjVPf
ME7y1NnKWne0IZ1FEi0l+mdLy86UTukeXUocjiVBuWi6kX0OpLVmf1chiZB9y62L/ADoZZ8n7FeX
SlBcCC5/EM+gpSRvJnj1KxG0StteMeEPawarZce0sQQmKG/ywzd02CeN7FcNy+iGMTClOh4CRPpL
cAgPHEHH5X6IJRf4gW7d8zspEV5On3nRraBezZBkNUi1JaOq3WdW2nnowcLr8c8SSqNTApoX0Afw
glpGbyv6TJu8fMRniSiYaB9d1Gc+GsQT1KlIeHkV0wcZ7+8Yyv5/KfNONxEgE2+817rTSRCLZ3fD
OnYHJTZcrNWvObHlmvoxdNZLizIimzmsaIMq5G4xYP01Sw/o/SXLSedUjoVvtjmoVouRzpe/+3Wt
6eql6K8ok6DGlJn8mY4+oi/lWGMhc7/2KoGuToP30hbHwqZOBMy9t/jVJlP5o4vzgRVF+LVGZ7n2
HUa4jVj05l6W3mQEbVmP1frEK1RXMlF5cYXbmbUd9s398Dux3lTZWotWqRIZ3Ob+W8dQWDofKqMW
tjSjJpXMru4W3rruq5UVyrvTjQGyR3f/fVH1IxuIFiRVwDzRgUELqnv5OBMPIIzbZId/Ix3MPIe9
HiaoMrP47F+Y0DRObtOItjWYBesu7/jrwLHd2O/W3q+cwsgPAnJZs+TOHkOaQOVOZWYPvx1aQeuG
Aakk1VQ2/dtCJCmT8Q38O261zEHkhQ9DPoyrXeEPfd74BxC63whJPBBW56IvY+m2HjxDybrfCyLy
mZA6xEr8dO71xWDwEVwZ/TrA7qDPUGoxQ2tSeWV62HPkBrEEzsHH2h6KfwFCGMoYlmliTUNXkHtW
818e3Rjh6X54k7AnWkFFREnsrbJtS2VxjnyFWF0RhLWZ2sq3O7RLD2JfF0De6nDjNCE7POcGoutj
+MZaByBwzh1Rd8FN5qrHpzesNWmoSFk5fE+M4V/DFVy/tY897Jr7cjVUb8MSka8G8RUwq2juzzwU
ByN3eR0dELdC3or2fXvO7m/dRkNIrvJxEb9XiEh1hAF6rPsDuWv7KLtv8l8gAQyqSS+RPADvo4v6
K9c/8H5y3RPaqEK1eMlRZyNXnjavvFtM11LeaWc/rA6oeZw6mckZQvz5GoMYNkJnShTiYARXY9bX
5QaEvr8MfWuHmqBQr6cZQgQnl+Q1YCGgz0aL2It938d8npggnIlwhe0PlagUe1MqfI8IZM74Yrcl
KxK6HkBkdYTFXzPaU0KSh+dHidIawocjMF9oya8rOBMzzNNJmnXAfCpY827+Xf9qyIIh+/7nkdXW
So/DDvv2svW/xQqJStaL4z/oN8fUGxGH5IT6Hlg3AQj1Ybd8vMz3ii9Z8oc2Ts+Rxlf+yfwBZU8I
ajFvfhXuo/ZZs9P9FnSBAl4N1aedLq3SAbgk9Wmw/jbS4Suukqr84xt/MFGRPXvM4bvmgl89JJDF
Ppu7PVaKm9FJVRsZDwF62w6MclBwqz/I87hWkQa7ppjwSpyHKSKqeP72Q4B8QQZnoAK0SM3rWy3Z
05ALspWkAHtrGlcqcyguuWbMnlMWfLjeKzAOIcDbH8XaB/lgf4zlvKKrkbXTH6TAt8wtzbrFyTbL
ByO7+4mev4zTW6Bekw3yLP2ozHqG7m3fmhqeTHWOi+vbm+rIfn7sTKGIIj8feGP36MudjiIiogLP
qe1bkg/wWPEEYmPqs6FyqD8ss6NWpM4XCHolbgo5NEKCByDx/mpmhR/NnA6CdusdIk8rEEaJyDI0
2YapjP3Oki6Iv9JoPoCe0SfO8I7kVSBK2+ojN7t2gqtRkmAlrtlwf01G2ZtT1gJuBu6ThN7EjMnC
9Ig39Vpi0fHIbvr4LdOe/+3C40gG4OILxUWAijwXWXXdGy4l6cc0MhPTl12TI7KFDM/ZzNhq2QuQ
pplNB20WE0SVtozqPXn16AS+2ABZ6rmk/DbkxC9HrbiKXbgY+cJ+n7qlsP0z0y/A8w7CnbEWRl2W
F8z7gU9gdQp4xwYTeZYbfB1lYH+DxnaJiUQcdB1jKxwwPt7X3bhUtwylDsHm4hktCEFjKHx7NKwX
o1NlDF5AKIFe9Zl3s3h+1Utrrq7q1c/Rg+KJnm9JveFq2L8+dVkdLe/iDL6QavUDfyFFtbn8Qqo8
4CXSbKMi0Q/MOVemg7hNvNXZ0Gp23g5qzyXnSTmbom8mQvukDHiK4ojXvDDVyDhKdXzkHIJSHO1D
G4JbaNdQ1VnXYWTS8hG4d4RIEYxvw8rZrT3nQvcTqx9dTysQL2dvE1C0XF94mDH5qpZk7Bgkfqld
/Qu6AJOnM0jwXf4NydTcaG4IF0VUIw89iQFjWJqMvjVz462rr7gbFmfuPb+iaVWT6gvBfV7CqAxI
ISCrWkQxeiyUYWaxQG6WVu1IEZSHnv8/rSYqiNdhqApZRUnCuRB4/X4IwrzTR4KdXWfzHPV09hAY
fWnA1NOA7UmO/FoG/6AnQEf9typiBn31Q75NMYbdVtoTE0mu36PPg106xP2m31vqNoCSSkhASk0N
VO9D6uWZ/ncT1PZZqwKxJwcZPC/d/db9s3unE6O1UgI2j7Y4nE2MckxrPjy9zhA3c5mIH/aRSXAq
pq41iL6BJxHkmuJeF6RCDu7cVll/7lo4fY5E9UnDwvmZFLZ7VwlxtbDAUVZP8lgIys5J589EUOlS
rHrxjDy6581xER8RIrpnftjIoP8HWzCzyHRRFBYU7qTwR6tuWS2bA9pqStBmXicW3hxXQVClXMIQ
vH/UnCbboY2+dEpM4tKvBa62kwcoQB9sUeHD66VVaz3MZ5rVevoj29g9zHzL0zDXGHyF1eWpLmlb
4Z8+rzklsjXHhO63DE7UZ2E9QH/liMNLSVkjvYcJrP/4rwV/KhtgOlfmrhrjePPuQxOQDY/W7SUJ
ZphbWCDlmsvxsv7i5DZZnMWILnC9tqSBLaDvNE0czgI5M4WvTNGAjDyluAKCU8kb/rPywG2ot3rm
PBruV0mCpDNGxf3H2Gn3TPP3QCMA438Z5gXt8oit5wVore5oxdK3QyvCMeSWRHtJFB58QaYsH5tK
3K+7DZUFd3iVPacGUtAc9seg1IPkUOfypPoefHAXcypkbNbQpwCYU4edi8t3vFMIchCVU5t5yPK+
NIg7hGilTRarGGTR4rcuvrqgFJ6l6JdTWuoPlZPmdgG2yU4/28U5UoDJ+MOlH9QdwuKj6Qs7XGcy
JAapo41WPSjRiaSkuUEw/bVrPSiz94rsU8uZXaMFtGyuXaBVbNAUe/kV8IXSZMBUzJ854mPkBgag
T/cv5Q8LtqyOtpS82CP9X4SVXWtBxpExYCVpqRyGgxkyItIoQ2IMsYce460eUr9qN96ADVOCc79Z
yCEYAcQ+TvzPQ9LvFMmXHFX+E+k5X3kPzHIxDAxERGTDUDI5WskLlgxwHMk/cvC0hcifIkx3XUmF
hQuGRuAwfoHHOo2fOBvIJC3Qse5VUosSfMA7qhTz9gUi5QnfgH97Kw7oprnGOR5FfnMiEzOA00ZR
dR487BsIxPHJmQ1ZY4WRlSzIJ5iT8MLmAcyg8vWmMD/QkdBWbCOd51AeE+aVPScVUYvLGumzWiEa
LpaVYrNgbz2xAYKDVDZ5TFZjP+ORO7l5Rd+fPo4xwEbdnUX/aXnsM/7zHreCN9uXJjSLHQ65k2Gm
6m2UhSES8xsbatuVXll1eiT7/ACoxzTJXgBMD3VmmVWSd3czT6GtLAYI3YyYEQETiIrDpshyXEGP
eMq+dqhOOThUWF9OahmwVnKbeEcQc5avqmwPAzw7taQ/bALFKqoW9tEe+U7wLKoUiOKPqS27fvlZ
l3QuzxLYZaC8ZxGgvFVp+3Ef1m3Uf7P7Oq5sUzy5B0tHMZ/EJoHL5lhiIeYlgKyj0LOgl70o/s3H
lU2TCOoha3f4BicuvpvT82HtSFP2j6O6ZV8RhYpsRzcycum6cftZKh41SHXv0pv8bBMHlCvPPNu8
1G+yDV37FtrTXlP7dtYTbMYG+XYAJEDmS6Bllp0tGZi4nVifAr08t2kcYs0sQpVKLAbiCPCBiTvx
MX/cqFEYdcze1Ar4DwQxlmmn5pTMCASfehje0Wg8Q4hME/TomOz9XUOjuuZlnIKOLim3wifbi7NH
Wfzh+vHWAaS+y3oS+rPMUmvx4EzoXcO2igQ9+TbSZX/fYA6tOn40SNHL6jpQ2DsvTGhzSQEnZXH8
f5GwehiOf/t7Uk4DR4O2kFnCmNDu7+xd8P8eiRt9hqnrnf8Anw8XkA11flnx3zjNnwNs3pXnsWcd
VXD5W4+7lj/DxIeqxI05qPkQ7wPJWfLuWzsgWXNFdWvO5LG5Qc7eHAP9xQOscfAi24ZHKOuA4vDa
u/0cYQvMSeQWDz1BGDNLEiH9CugXGrYycEev//CkJJW02v8fAJ5uBPujgdUisKzdRM17wyw/tPh3
YvhQBvE2WCGhoPxv1QrRJQi5GoyLtJ7EgKhP2y4EXEE+vLXcRYdbsrDGWg4+NEVTSqu9AeDwHxbf
r0hbRZpvD7r40OtjETA/rpy6QsoHJE+wY9+m35Ve9evhz0oVhJP6179V6mcagwbmBZ8jak2lDdKe
B7dEzw+hCyO9NhsPUG0TWDF5JJyEVk+NbWlkyXg3aqU9uGADUsBayw8VPmV3//v24uLguhQA3Nkk
tyQIptBe0g24LO3VKthGnczd/5GSsU5APOISFAF73Xt2GEVfpotJwA8fsKEEz3qGtXikIzwhJhhL
0lRGen0CglvEoOgqDzMa0iF2+CtyGpudUwoIVZZvEYDGNsUret2e3YZGHRhmCW7V/ojzln65n8O3
Cihhf8cuQw4sWvK2BYWgdC9N/F4cHEB92kGYWlf51R1KxPRg7qPQuLhSNQnSSpSIckMohSxjSUu+
/C2+TaJtpS8ySLsFuA0325mukkedfmvCona4hyN0EurcBl+G3hlUCT6hoq1UMLQG10FZupl04c8n
Fxrevr9QWPhaldjbSQ438uvHFR4DzgPFl3G30mQWqlP3s0vz8LvL79wu60O9qemc1m9iGtxJ4z/U
GHt/dkcoHqrNCM2FUQ/N8tmgleQZNO1pnOyF7zDvsW+xsv8cmJNeef8rDKapwIy6XMefP0BLeYUZ
mLIoOoS1WdJnBfjSCfpzoeSRo4kxJlBiAxOmacTXNSXyxR2a3df2IbJqN2+R9ZttP98VGFdqjJ8Y
Fnp+YlaY6lthYDJ9bsY4WxJBf2du0cO++i/1V1BSi8ZHjOY0dsadbTv62WYO/U1eWcjkCuhg+HX2
1Z01LcOEwumI2dp1O/X+K27+AiXRKIa3POHtIPUHoLvZWOktOsRj18pi4AAa3j9OEYdV/zK4bAkm
EpkUzRPWpfQbT+sVUASq21KX09xwZ8wRpzfXt3Fag4lnWAmEyDV7hklZioWsSTB0AIf4V3ZLLMRl
5PW4EWjApV58yNnVPJ43GtDf7OVz80dbaaz8eyKKBnWSFxanSsBmwvwtI17DMJ9DmYtRJpCRoaqn
+X3T0LlXNLuHZsiFMl2JiQ5MkR9PTrxUIlwx9gfvltpUJdaGxERoANlhzRdGR1UCRVVr439xAqJ7
Mt2dMhDBd7zq0KrVaSg/xRGF16f6MdrciNaiUhtSrbaWCZvv13Fv34cec3zkNV6ohjHPH8agBJez
tvTCeepvhhaba9DMtCgp5VciTwyluer79UIhCnhGDfC9YuGL0oYseZPjzyWjuI6osWiq4bYeAYAk
JkcD5ekmnHCbYMDyb4DSqAwm8B5yS+VTDdyRgI2LqKlDnPsK/UTGVNjsizsQ8w9ylEitiwW8nJKr
T7itbAJ42pCK80Z9VIWWcAlG58vnyOM7sTXvqFXFWEK7w7ihndl2uAHevuc7UoStSGDHMmRfwpmq
RKKS9xIpaqpIKkiOnkoaXXseZ+YBGcwEaddNvTC7p/QVi9phJcJ7MmuPOCTwr7n3j2LydKL85wVG
nIWJSy9vKY8Wb7yVJdUVe1bQCVA3aZ9gnCEOkDPetJCpqWdzaEyX2IKr9RQ4jZQC39Zf4VqoDQNC
nZIVAJiBkqbylEIqTJuo8ieHjOo/nt0B8CeAW9rILZZvn45dlEF8TN9rmITSzJ9SmqNW63ni/tL0
/pS8acFYvFuDfurbRWPM4i2c30IhqEBQLOAkuZcqZ4XEDxpVT4hhaiY4vLbvBQ/+OUez2jd/iBQU
ADwaNUDWPCb/4tcGi1oNqrijOIupYnnBTR2yK8aI4AjPuO9WMEElAhlp5Qg1jeH8Pm+cTzrNkUB+
7Mw9Q1AIeU/yPYrJrbliihreK9Vvz1NxsobNgfRxkCKMOJPNpQ9EGLv36+ufIMv9IzS9V/x7L/dP
4R4EpQg58D42m66OmWEBuSRQdSQc+BAwxn79415O5Vwy/Gl/qQ+/SMtG95mWONGYbIq90Aw+9m4F
9o8KKfRWZChJ9gAcSVEhQsqEx1tLXNpL8ZGz8suTfaFXuw4wMYLLQx1EOSTRY4TeRJtK/mLbMNeJ
wqcC4/1jmNYf+rlHvtrrn76bmbaqzkIm3NoQNJ6OgS70rYvrifua5YrKpQf/9EuEHj4doA5KuQnL
noD5FUuI+yQEqQj3gXtAg/7IiyhGmSuAq9pJPp0YtLgAziu7ZwWEG4GQRLQdAaT0GyyoZmLOtRKt
WLpuzR/VrD+vVYF7i918SWS3Z6K6kAAonSeg5Ii6RfqeYWcLiprGBUCMjHqZ/Bv2cfr0NHRrfYvx
AGPxR6rlOOM02QehyhYv7VG39DPkp2uG6+nUJ3fHZhPX9dbieRrInvz/tat/SjJnsT8QfNhViYso
/H7pjPxFu3acIIuNO868rl99yFnA8iWR9tE47LXlmvR49G0tWtbDdIxWkRUMz0dzH6jzr4q/PrW4
fpdpbq/jpRRoqhwelN7+wl/feWUXKvCPJCWKoGrlUEhz1bAnbO6BZ1Cr6blM4aIyCZqhGmJOfgd/
EpWiMTSjDevBkUcyVNdJwW5l0kA6vBdu6O741MqVBC/b3YkEBhyEl4t0fiZpVUCGeMoH8n9xU7Ox
//YK+h5XenEJbEVRnIvaqOw0EAhKU1883Hgvleh/UFn4FkpNgwTwkYBgaPv6tj43AnOBDizURSnA
bYciRZgivgMpm+6T4trcgdr7v8CWg5hOLkwq/vSkT53Fl4gEGVKDhDOQjTMraKbkuPxraGbMmsdD
O950lKw3DMfHpaN7rXIkVYFuN3+f7XUNPZak3mpPwgkfgFBE/oA9rf59wJwdz2rzk//Ga2/RuxEd
nCTj8DGRbYuiPqwu3IxpSGxq+mJF16zHkE0Jrw11yrpihT46ubcLaHn2BzhPVkd4qULJaGlQvA9B
kk7A2jMuHzhx0E7MmnLVWSIID/1Oh7D/dre3A6fPyrmRrZMgsXc5+thBhg1kWo47Viuvcb9MA5GP
whOt1BL89xWy9yQdbKL6Z9QcoBAcWVjTLWuDZuSkxjbkw/Um74obf7zDuO06BUri36qTgpHa7qgC
qQzKQAUPs4L7qPLgyOcMPK+E96YzBa+06SpKdH79PGZ8Zp6e7AAJESBqbvbujHNrVLfcgap4GvZy
g/VBW23p7pGnSgLL6Xihm1wbXZirTPP0eg/TNM/S9guu1m1GeCvba318WNeRMOp2no8eSfNqSGlt
iv6NogIPHE+KHrYlf12+uzoh4Wy9l6/ID4S8H/0JzPRxVfk9+hBqs3mcNhHBpePRyA5VbkCU16rc
UDUo6WZ2r+pnlJS/ycyFIarIrTeIfnT83yx4woX7MZNOSDz6p3e9LzskkVzGrcPQSq2Dk/J0NGlh
d7xiAFXXS3aXkkMLgbp90KUMllb9qtWJdNNc19VUpJUQADdnw4YGOlboeDdQBRkvc0UMWR03U3hc
Bs72qFPRWf8aAvcEwpy97rm/GKibVR8Zajw9JnDhjkl2DG2Vqk1ToWyqXm+ugAV4t+DZgNoM999H
xDvJG4X9/aR3M0INECfs2IxMCqMgh1jJp4TUCdSrhCWjqFiNkn7x3BA/Ow5+LQ8gObn0APiar89p
1KXkybbeCm/DWFIGbQYeF8r8nLeLC05POgKOscLjGsW2pxDC6s9D7GudmotoQdHu7c5FV/RmeN2x
73flfHtMxl+dA9odXQrFuyOtc6G9rZ/TPb8I7mw4S7o7tTVyD19SnXecT+6cZJKp/4mTzgqtORQT
0ukBXBOWNpNCmXGJUg5cnGtSKuANPaoyEv+Qz+2254avpK9pymVLOuC14wSIuk1wR2phYRuU83Eb
UzL94F6s0i/OlhiZ1ab1pi4kUmzwhahWKQ2rwH4WqAPDCk4lacgLK8LKeUFxHiSR8wOOG02Ti10v
upL8/iO7lB8lYjCY27pGtfzF0RMM99GoCGBb9Ro2YIV8d5Pwd4iSKCOoY3N/1A1WdxHazbMWYeKb
NcfIfdVVZI/knJuxGlKxj8fIpzsYR9gtLgseYm1Ya/UT+l7uvLZshrg+LQkqbXhpRE0cBEA5FXuh
VjBk4ALvnYy5sEcWm208SP9L7jfRMbWd1+Uk0513/nOIrwbov/fQL0fN+u7MpmUM93Z+9pq9B3rf
xhAAilTKc4IziH2ssQhoTcafRETfI5aWvm1duKaHzCkDk6dts71XzBJ9rKSoHViAKn4iqUgT/FKH
fPTcAtHc57OaZ4172329t030XsLR1HWERSS1kyX3ujnFwmW9jDBythjMj3UI5rdizF4f1+cs3iP2
9+K5FINtc3ECq1C4F+CF4hcr0G8POr9ghjmFU3cYzYhnp8FT+hX1W+T04knK4VYTT0CQksmDRu8I
onDa1tWADb51ZOWgTGpgM/cT7PgDjfDglHeJUXc4ljibGKsy/A+BTw9+E9CEgnnTZIMX5rBLU0BQ
dvhezM1FeQz1oR5BHUcFf/Ugtn4vEq/WpXud5uvHMvk14LDQrH4eg3/8r0e+fYiBOn+HmEtpz1/3
Wls++RIc5kMZcG1EtOuQm92TqLNNYJld3DuTupHoHjSc3LzTW7SvmNE+M1Ho53hrr5nRO0K0v15e
EqedcTXeKfneLQM1WmU1aM520eom9dE2qWu+6ieG2Iom1/0fz8AWyMJf7bBztsWbUQQ2VTkof1tQ
Q1oyY0kdntW3mWJfFZenEmVdGo+cocQl+6u8/rgmE+3l5hbKZ3MWUiaViFGzjtcxBAAfQ7xCH7B+
Beb5KwY8/guL5+d028G7Axt1O2T7CL3dSE5a6Cgmi2TwTN1Gi5r6jDeusXgmJCMo4rBm6+VzugTp
r49mCm974E864Ec4o6RxSV99ml6xzQminpICplX7xda5x5qpeVGmJE11RzfctUA++TM1nyPgROUf
fgh0tb4fDVwDMS8Tzdo3aZ7PQSjasrMNBsU3n/TwLTUualLODiLweiSNNoUaeJgI4dA9Bi89XwwY
ofDh5G0hqy+xgnWmNZ8+9WKLhZUAm6LOFRVIqnkjJsJqF5zOhW6UeDTeRhdBFsq22WUXRj1Tvv2F
nhw5XaGCMZNB0+TVCux0BQuhbqjtsrUBjvCkl0/emRNlZt72+hs57+h5rz6ggkBcW7WkYmw5GfbU
lJAtwTgkmkej9jH55ufOI8GJlQa2HXhAXtUktU5RQKNWslHqMixcW8+EXk4KifGSVFht5+XeJ4kT
LFfls+MFFqKNO9shk1aN4BJVtOSf3tgNSqV99Eqs3RN3lr8nqR42ICKEUM4ERhFmXnyweJvKjSiX
eTL5eGG2gkPrm31VacU3vGpM+dwZ3sSbhSYcrpB01prpoiP0RJoCTIR8HFD8k3x+OlijqEmzCyaS
6poBzhMt8o+u2kXz5YPusiCdnoXbBx7I0omK2iTnAaE4FpD9Nkc5TMQp/UUW6geYjBnyLPiVHWvV
CNKWu3hlcPw9o8Gt0aGypsKU6agPxcQLI/6jwI+J6fevWDJyKz2qGmD0DA8x/fD7b3wzGk0G20J0
6Gx+/JNJ+PdOiwDsihnMCnxmNRBrdV1LJXfC62ETTFSRoul3Sx6syT6HQ+Ll+KrdlK9iMmOmc8uQ
wpZorPibHM8GAdMo28cLOY4OrSx6PcPD1q0+Wfm3qTwgE9pO+DhoZLtMuSDiu7kPRNzoYGZiRjUi
6ffHkvFNGrQ8TEHlpBKlgASBufNKQG6xJiZu4quiyW4G6XHv9IzF0UeRqDOyrEkYFUd8/N4lULNd
oTe01Od2rS38d2uTDumA6DhYLDp1Bl+damenTSNn8tGnRG3vgg8v8Ibc761ASugFECFOynxwJ8rd
jraMNb1iEQeqHyv0cmbAxiIIysy10XmvP9nE/sjguD92W25WpSkr3Kh7kMp5e9R3SfIMt9Uo+Cqg
Az/e4ZQvrq12CdSsoIl5agj6hq65zVJ5cw4zkIXrxatYDwpHIj0ac+TAsqo1z3mIKljlBK63Cwva
+sMusqA1qFUjtmJD55j/2EMvl1Mw2lsNS7EKMl0MMQOyn+4oJKvW9QYlqVWmt3DbM7yFM+1LhdAi
k1WmRqql/IktHBLery6+MVkvcORIz8F+p45GtZ/cMpzQoeWn37sYo1bFc9xMA8wcwRhFkIkkpSYB
EgHahZ79o5Z4+LlXrDX+JAoeKoKSDB0tLx1vf7ELzSqUPtRqWCSFmunwDN980z4oz/HYQqPsCr0X
QkvlxaEGfMjRHkWWMWDzXgu4fUmlaCxPxC/Fd7uF72EYrU7GHPEL0ntk7ERWWgtWK5+IMrboVU6z
CSe42H6+tEZp5vWOo34I0XlLPEXHbPEfxkWRGIe+aYWSFd0sWv53QAvFepJw73prLWOjWYHIuUJZ
COPNrWFgaZRaBS8ChdOrXW4z7cExRwI1YqN9Ze4Oabr2V0ZZzSGWMjyUNNGEv4/jRipz64fML7PN
kN6sm+LVmvcnsfS9SyBePfWkP3l47z/IXOY80lpI5WbyRu7bMxIMZwlIEdv3eIcrjlwvWDruWMyH
jBU3WhfWayw7Fyt/cc608O7YgGYEhVZb43SBhdNQq/jthoWp1f+DEKg2FTT65ByOKEsDlMOkxMBf
IJRe7Je1mXC+dHrzTfpz7RuhNmAZu0aKjcwTLK1Tztl/S5TXB04Fb85Qmh6MTbhueafVCKjnYt00
RHLqJl95N50fEv7fNQHm5u4jN82Oar4QNlF0VAmowh+je4b0mehOEz+O2y49fCXwUgOyxMFF6x6/
TYtrXOIPo1mXAuuuI1bMDYbfH/6ZMb+HNvvg83sKD951RnE/VWPowh0t4YLEvfaRWlrUv60L89F3
dTwuoZisgqKD4EV5IeJ6xThTH6dHmfLblRbkRzGlJYa2nRr7Kolo1i98QC6UrsjqIt3wGRCy9+PN
LyzfTta6a7CdX7cZ4d9yM+KE/15Oc2Bpk9LnP0YudmdNgWp0DJA3Hz6MMnQgF/ufsVD+DSzESEqZ
p2czq7Uw48L7b1/IwvePl0PueHmRIEmHehyaS71iwYYzIzAREi6EPd/T4u1WV0rTUimK/8vxPXbT
DBhHKANKeZzQKMgOjg467jJ8QhDtXatFUGIOCkUl4a3ADU9BqqEF6XtbWOaukrg+4uP6wpOpb7LL
XV0dRBgQdCf58xoqZwjLgZP+/QMkUEgzYnj/TH5BPdRuX1UvAsmw8mvCCP9H6DNOJ6657JyOjDIb
MeA3Kv0v2jwoixbD/6+ihGtFWJFARWYsbZ/8+6CsW0N7fLQKWAfAEuvCSnCbvCS4A3QACLRb87RN
FWRrz/Tb9n3ginEnxIa3O0ZjOQ7jH1ulXd228JOvT/m/53n4juplbMOajDCM6lNEfrUbTNwaJJqn
NAzO80ELLp1/OEKeOLy0lu2EaxXg4+GTu739Kd40yCIi06/XsM49xqDYpQAyEEJv1wBuJ492h8dj
IjIafAb+CUEFQRgiahG6qpM+uTHSN7kA+5WBYGTMgZ/fGqOGzN7Kf2g9HNRQOBdymUMBgMVCKHBO
qSaKH/66ZmqniWRL9NYlO4+TVTOlQ9wht9RfN0Vc4zU/XMReGvtZW44FGsexUwHXkzG+xx1O192U
iZD1zQDT3SKcv3VHINTQTXOTvJuT9GucrimJU3b3AzLjf8PwXDc3p47tqpzxNEzMkvBhjeHk7a+X
q8acHNuhW5IRVLkelzHt1KH2E2YiS7p9sLcMPt5xLsPhamItQe7ZCpD/7bfyebcV8x06fhBGGft7
SofVPJWuKugjtwCheDLIq1hcZRyMWvHRUfkVrqQI6G2wKugCnp1rSHnbHLiE5tVLvl4FZYaqJdyQ
Q3/E/zSBsaLzenpTBDnT5cHLgzbCIGRqbjt7qddj58Xxs2PslOwCl5OKiI2XlXeCtdEbMBilEzZ0
qv+k4/qE5d0nKiB7dk0aVXlJnDTswvAX66Z9bBWANjWSJgnVf8SvLNUiKKcfO4rsVzbj4T43r2ml
/UgliwjjIKN0yBsIjirjgkdIYDQPMKccvtG8DZG8oBZp+Ptms2XaICn8go7LtvooJOliNOAciU4E
mtI9PgYp61tmdEsgRrqz+t/7+W2m7oCxJ/CySrNktCjS5rxvIVrqglCN3043dJIJ/j1cGoBKBiWa
YlDyG02TwGr6zRv4ogAqjEEf4+sz3E9s7xhhd7AGz8GXYlnvueIZFJeg1BkRjg6EmjUtcuDThHgv
BCmMfV0tjLQIz/5eeDrX1xpIYX6TwbHdHw6Q6wSHBWuykMYobfC1q26giQjrrEOzyBrL11vdaHxJ
EVgO6n/NFd4B1bkgwuTT/ombFKUaVFtUFRJqcTznmoLni3KsQwBwrMIT9IeXWLmFFJqhly5g+GK/
NU2Ia/TGNWCAWhyEfC6cQ8RQ/r1pXZBZ9KDbeC519O5pLdUyo55ufgCwqahfRKSqhO2iYW3NG8lj
O1Hi4J2FiGkSd3ZGp3xH/kaajo7ZJmthu6yigdbgeMykPlJl4M46+F+Uog58TwB40Y9y9VGK3lpa
8wtE3wCriLWfuGrHzVHx7ctaO8HeXXqXf2sTg+GDh6OXGXVL3YwcCSIlfN24bqbcWoT+RUlx7sRn
+gShjrOHCLjkKI/FEMYMepY6y3nwImwkXFDOVgkSvkwalP9k7lNekeAtCgIya6vdNGcMHLsAGoeS
IM/jYOKv5iwzTbPJdF4xl7Nyyl+DIwwisQEw2yfdkzQi2oLXYHtws6W3/Z2abZybP8Z5mDxYzwWq
FE4I6QQzD0fjA9pjGzH329TJ9PSpIEI/5lhABqNVvqU01s2zQPehwIzXS3Tt4wwEPQShR54t8bYT
fDxGropqTIfXW9lSxfyoTqCBokQoaoQpaOKVbC5Pnbe1LxvDvBjIEYLrWuL6WoaxnlFRP8K1pTNS
3eqIOfTDuMlcIoEF1lzxWHr3NA4d2VoPHAWb+o5mZacCxxzw9yXBiZgQGa0LHCKttsEBW54LvHdr
wtefHslPIf4YJxInsWI984fmmR3b3rZmmBQYtQ2EyjoaTYj3vCiJ9eAGlj8FYbzJn9sU86lchK+g
AHCd9XgZVlOsCtr22FwHOASfw4fcuhWiObIYgH+Xh5S9p6JhaR8lfnsZONrQ6EwuFGdYC/wEax1g
MfLilhPWvCoWH+6XiiGtBu2HpdiG7CeSX3oWJkLHHkXi1UWMK751k8gv0DbGAGtXiFyRcGQ/c6pG
a3vacY5/6fEUL94BFI2pPpHmFVTprQ25xDYD1FYo2CEWGPiov7tzzwMDm8BVhhgKbLZG19d/o4EK
lHkcrZG/ib1E9CGPsVKpQeOiS3GEUF+3+4Ow2vcrEbD7XAWmJC0+Co5vV/2Ue5/8WBbCyVHPt5JT
PpYN7s5hItbRt8jHH4y39jh1qLhsd3IP4Cw1lVIB0PHURVXdkr9bAyfqXqraZgN8XmQbzv9eOAqv
1EDQAaC0/pPRY4tbGjnVHc7NnidvTunI1YaT0Ds6Xw0nrtz1iVBN1y0vbv8Wx1lH0kXrbhpkaUOw
uTfRVVCzXAPPMnrmJwwwFWdKR1XTiaUnY6Mx67ACBj36HtNFV2uATlm4LcSGee2LAlywfRHLln/X
ukRk8XOihLae19yIWD7l66tbmau+4WPHMzxDKqnmmBxFU1etQ7kulYUz6pbvXWnCCfwjFR82bIQW
3lDIQI+Gvjaw0YXVuqQBsz/zAd4FCJaOLkhrSXc8McoHXclM8tNDXBRI8MQl3AtUZc5bidgEet8h
e5V2j/z/aAQHYbiF5iqWEKIwSaifA/XQjrzIvHmNc0qfjWUVdOLWQrXc/lwBmhkGRJWtPtt47839
wFqp4ieu2nJyr8dyI6kyj2vuAUngJaOeO2YQlwL1B6x7AQIdrzV1ro1lXK0mnyTYFW5M+Q0sfkFG
O0+ETXJ8QxZ/+gO06ffUbCNHIMAdLRbDjRlslRGr2bpce1fmaM/pvUhKwc9z8OKrOylyBalNaA0C
iYRB9NRiyuHaue2PQtmVqxG0vkQhy6idbSUsaioC6In89VG0WkXt2zsNKz5rOJfb4rpsLg+2cLpx
BWv/+seEGYSfjRo63tOFr2/QgOkEmXTSTP2e4URgX36stnUsQqWJbI/wfdtHhPCISjgDV/aKpiKA
nNCpQT/QS5f5MEB6xkGgcYZ/SOHz74zdk5Pvr+iHqjg6Jih8EF4sPq88fEvujieg+PL3hDLSBSE2
c3VboeYN/BYwaCZCqZDt+t0C9a1qE+GQOJooGP3UxfMQ4+uFVlUWyg0HFfAc+R0pOQksyiQIq99d
x0DDWA3d8iVPuSlj1104eOh2vP/jgljd6Iy1DLw99Cyl1z43Kr8RVYbdUIf2pEERQjcCcCWj/HVK
59W0LvGbFffBkWWV1/ylerWfUuc7aIz6k3TgCC6Tg02QU9fE3XfMjjRt5UdP6NDeW/HuSus5a0eo
b1dCPH4u5odHkWbD9ecye771Ann+dUA7+g50qW/17f6UMkHyX4FexWUEoBIgTSECli+GVRoo56nu
JHx+0ri+N0JblRSpYf9TW9NPUJt6zf4LECJYk/Rh5A5XKw/PNyes8YCBswNQ7+9VI+CBQ2fIlw9C
VhUFdX9JL8+fMPkOUzRk/FoTVxcEaascYRkGAI9zXfaNuHaf/4z41t1h2bMaNiFSQW7jLWOwmldQ
IIPq31ZVtgb29igNlDkdMRus41nU7ySnpOrvfRxceJoN1s6KSGWERAvC0sEJtzqeusoGHSGBX4Uu
dq1X/P5NgPdWQrABNCIMnxZhcL5ewMOFnFkS8pxw/o5t+i/qtvHsKbfsIAEbQRnzS6SFct7oWNg6
+Ld+NaKYDIP9qTCXUQR3G3WKySWASVGOadjBuU4eMmO292r68nHpiz1gZ2rkdyF2ujFSb2LfqIPP
CA2nNzIf3aF5/KETl7Dtz23HD3PsPVIYm8u3Ymw1sEkCfdp3hRhMLBse1iDe2jUqKPW00XNIJlnt
Uiol600AGml+COZImv4vcAP3GXQQbiCNXnXuldMxiMj7qfUgdQdouRwZU1hubFS0nlr7skQLa2lb
Ctll8RXLRtnXwMzL4rziwlx5M7S2ptxwShnvYhClovmJrtJ8C9JZCb6nhNdBTTUEBFsCm6F+ixFQ
42cSDyETUjaDqvMfrXtngwjVmEjW1NwRhQArT2VuOvmZNQRayMj2XuzAv4BUtVVhZ1e7CU1va26O
oZ3mAaslDJU1y//t3JkLXI4VBBc+MLQcaouF92ADtX+oB7muxRGQo+1JB/9OCA7bQi2UHCRgOued
5YlSmMAVzwa/APcMlfzJ8+gZLUBuASvuaRJj40fmdq/M/P5fxQBiXp7fV0xulDeVcHXjC1N50ri1
nNGabTy0hh9aqQvRq2jW1j4N5QKeTBEt74ugVZoi5/b5fdOJI209l/DcAaGgSEDlMOBhotMtP1RN
v9tDznxqYxSCXAlQF+l1kI8LEYbPKKzQpvc2qQev93CR0BkV7EjXznuHh+y5L1YKf4FLrTIBfHfj
Tm4ML2kiZ2S8FnV6RanW40FWri1pBkBnuEQhIcqpDHdf02YM5cOmdyTXm89e4okyNtl6LgxeXBTh
kUwBio7vCoCgwJHFtBhduWgxQCfb4CXql/Wpe/2mnKEBzTkF9wk7scpOoigq9oiMqCVfZXNDKIfC
ihNfgj3CvwTt5l5Z/ZDqnGwzfPbX7FJFGi1Vq4Hu8W44PUcqa33sr9Tj2GKrmqT7M9hmfZ6E6n96
lNzaFkn2RzOGYUGtLeqTFl0UzcmcaF/hCv/+SLs9jjzt1Hts8p/crpOr4YuwXQXIy8YdcNr3e1yg
bMtgmf2ylLFn4QFpRQ5Yxd59ccdkgvlorj7HHq/zn4MbEUeP7VBQuGnU3Er1Wixs70de7UVS9hQh
fQjT/rg7zoj0bQWBpva1trOKRNDMEQ2vbsJxmJSNFPX1pi3hVvbYN6SkqLs6LHhq2P7ZtzjQWTYq
ti+g8Qcz700ztktrj3k9VoSHpPlVxSMoldjImg7YioK9HW3qfPqYm8Iy5+zxADbdngbIxIYGerVq
aEsuxMwFeiX/aU49d7kkXQI1CAcpBUAFZN6kCkZYDGHvvdxo3GQzxBqFrPqVpz+XTCefZzijROLq
kUYWP3gyAY1skj2zvCtXts2lSgjvKuVuveD3lTb8PEYC36uiAOaGvuFn45bkaeLBGjmybtMpAY6B
xIW83IqoanTUbBWuG8LeELhaEilpk4Ni12panB73z2LGPNAomCvC/5V1woH7NnTORWV0Fe+ai3K5
dWcuTRZukZcR70lWukWbW4gvaAzBhHrMadyXgNjbX51i1qANMk0RivzxDtktJ0KzXRxAycdSzJKG
i9CURnq+4QfabZqxsvrCQCWC1Job8QKmTUYrrFBHH53O49GOI5UQHl/xgnDqvnYyhJH62JA0X2fc
CL5oLbDIvi4Ssk/sQe2RYwvklX31yzkOUoHh4wKfOnRRbVln2GXw8RX/YuNxX76RJ4ls0mCp0+Ps
hMHoLMb08xWLDdAysWkvC65xHLx26VBIXuIMHOn55cAM7v7OKp7tkzmSqKRlJa7FzS+arVAwwzqT
ykprM787XR75eRfNxxQdrM03wKBGJG0w53IPgZ+ZUFoCZazPvR9HzXCaSC2oFuhuQ0vQEq5EAkDj
TcwtOFFN4FBaNnzfb1zKdBiad9awsUZz8HVRNqVLiAj2F2XDS7g0kJXvchEHyvBqOo6mRtloPYoY
X8mZTAmafCPaSHQlwG4gAFtE9T4SFsxgmXW0tp8P5o/0+TQSoaz07EWsl0n/IzwalwI2EZ6yEzLm
cW8Q333dVRvnAhdqu4w19U9z0spjK/vc3zxOZt8L+Wq8nFEmX+hjnMA/t1MGUI6W9/TQ6E4dsx7R
KnZtkn1kogZxg7elKtqxmWu6xeXzNjZOo4786mzkI2FNF0bPUHZ/EoiMuFfo+qeS4ZyjT7uwHAw6
0HRELWGuP2mb2SZvl776cA7dvX+sWpj1bqCuYgulVN7tGOlCa18gzV77Ipy0GLCpYef/mAHz4C2R
qpSefePb9dSp7oFRZgLdKqyUkkCrKrvs5omEcVOjSMl3vS7ZOJXREvQNj8zIGHcVkb5Y7o0Yt/kr
KurX21McMFgeP0UreqMPsTqRUOsjtqskn7H9lwetsKghSMr7oHLwkg+JNiHywej7jMuhXXt02i0J
H2/FQFF1+1kiCEi3H2pR/unLBMebEttopVECMHrZ7lxovuD0SUp4dkAENSRj+P3ZiWAgMn+secCb
8UlucP52HHDwbA/4A0TD/tH5N/v9T9vrXHWH7C+EWSTzRCvHq0FybABgk3BXxqA1WuVdicodaaNJ
RJHPn1E1fQ7tY24mjlIKUisvV1jP+hEN8seVDAc5qiIH6zk5WfbrXYXg6AwCD3yB8dYPDKqnPMSb
9+yQXHWnQloR6W6OVhWUzLx7VsvrUpXCfyd5F0LE6FaQhLSW3+E1+9s1uDzdhwsBCQz/nCkVWZKy
t4NVahC00VLqqpL+XMsbvZlD/Gvk3t+LGQcKhaLY8V04PWvS8ftO2eBsenysUXhlxvPq0JypiL6K
jD64NhZTDl2ZsEO98T+ECeyfixm8fwaBxPxhcec9sYAa5/7B67SZzgXd9XUK6rI/GLXuaAgXuHSJ
5d6bAS0k0OmDBcyO4kpNtCYn13Td/gTvOLZocFPozlUSmlSgO2Q/QaoEaDkMrZqMmXdxA9i26zXG
HSN8b3zixhxtkkjvq9VfMVtQQ2U5usG24SO7Gtilf1XSxjyVeZ0JaWsPhDzX9zKYxxCqTFbs3Ol1
/Yz7clDX8OGaIEY07uhBHgLyz38bS90GA0GLcJEMERtTDn69xUbR9NgJ63DwTBbrqEM0/JmC8Ldv
wFG05/PSZ2u3EDtHCqJPN3m/tvIrEehhaBJNeRSjgqd2Tl8gNAkUpCNuR+qRL96zsHqGcGF+5btA
T0ldMBG0UZxDMDvJS/Xvg/jBu0yKUHHHOj8LB0P25gdrF2z/+wCfqllAhkuwSIQZgNsqArJtYdMs
u77nAnqliuAiw9JdpILgXSKfgICCERDz95Xp6uVeihRGKR4/TdReSHNB8seX12seo7Q6rLKViZTI
G1d/ylFT0dqNvbmf/bhwP196LDAf1rRyiHVynB2RlS3ia2eUSW6nLhjnPPJFIyp6CIVK7jmMsBIT
m5HbN0phSeXYAasMLv8ECNXSAWguLxrk4UDQSchwcxztUCtm/GzZtQ1SkNYmSnx0ZzYfKdheBnvO
PX+yXNOCvbz7gTCbo0EUhNgnCQbgok0PB0Byg42cjsigAeq2NShbM4WjrKqgC+RJalI6VNcb8pIq
tVqERZqw9ccKSA+L1WgrovIhL6r/+cGNUu68WuGX4vI5xEurwJoGhwdwK0OKoLOLPdND+affMrk7
JFZ6n4r752zvca1M/5VQHakbHvdADczWONIFDFUr91iTUUiIfKv1WL0qLLPJk9Regpw6ga5pMw8o
AilseDyu+oXLJ2xgkiGHmUo54iJt/MiV4IDWBOq8FPFrJNE5/ZAah3+40wLmwPO/G/oVqbROkMzb
o4LEMEv/OSzAzhhnYQrYzloFQa+bt1g1c7Wk7yWJuULOME+vuMBBcTzn9eMjynypUGueSq6Ve56z
eZElbof+D5MhVfeBoi/VspIGvnywVpkRNCl1X57hp8bYLd+aqMhXCDMSeK8FnbH5Xv9ov0qD1lhZ
go/GVgQWPTuxfy7C6oT/Z0Mt10L4Ae2WI6gBXq2exrEz9GYWm6SRXillUEW7CfF6tuhslvzslkw4
bXoJQT1BKtnAXlIhlM06MsvWEEYiHcVSVfbDXXbPGxOjNkWrxBrvOOmeh8kJE3FtR6VAPL2SdRzh
NFMxzkKM94RA+wnOlvmZp2tC9LBUtRBpj/9K258OvQKyqbymbcq19Erfu5hv+zmuEEPmlDjJkblS
atwLAUxQEP6942KU863ckLs+KLe+rgC6PxOmXvHRCKUy0Rf7MKxnvy3HPPUZZJLYh28621GAJPQL
KtajfH2bkVv7iIIXGLhWIGigi9X+tUbklJGfeLi1pAaN4Tl5n34D57FtzgpGwKF9Lu12H3G0p9cu
xA2ErJmA/XEiOqHM6JEoSVNSTse1GEs0A3NSeDgWCqCxHXSi7lCD6WaKG2/Yur5gM1MuPLd3Vr6K
ueRwnSICzmYRmU2lmaijf5ZNnP0nEDN6zmLNc4vTyADPI2RsfTNqB6El+93e5j2GcDdBaUAtFym1
RTpo7D3kTkrtU/BXPx/n6mYSC2WRLyPe1OabNbIol5HJTHt4JphFjoR0Se5PfqAEMWbZzakn6TME
RVixApwDV71/jFVEyBfDWa/Sl2J/dOQbTz45cCPYHafjvfc+4Q5gIM4kgeBOG3Pe0Ovy9B9zRIJ8
K8DIQ7Ly0BrlVNgKMIHCn5AEDbB36H8w6RDcySDj1Pksus/NNlj4qwEwOvN+3QbS4blWVIafxN2W
A5lsku5lX1nETHiMU0oE4Zz71DQ2E3A2h1mOTnQzJGHanXJnZNJcHkHJ8WTbSu6kkJc3c2slHsgR
PoAmygjg1Ffr8ENHTycsNOJlsYg36ESlwKqsAiWGs4jJCVQnUflrpfSIkCc9qI5Kli1QADdgxBWy
PRXTzZY+am2MLA4hdDXDDr0hLeGQqPZM4aTMY7rpoz3aI3hO8l6dtVcLta198ZraE43pbJfCYvwX
tUvGTh6kT9T67IDKzC0hkGaiLOfQbp3qCss+W0c/HKHfPSHlEgoXy1a8Hgz84n54wgjX6qgi67Zd
wLs9Bp644bn7N9X+1KXsMPYEyzvjrKkUd6JewfhvjrH5DeDqEs3/BjMAlPkyBq+UnNfLx2LGvYW2
zaezqZlauARvF1+ObMiCXwFLsEMQY1IUhKrpE7bWrfOlMR5um9UOLW3oNwVFLh6kYJGz3GKIeVQE
4Emj/GWMUmAmCef0Kyq/dYZ6Dh86QIGoVRW1tsEKq6hBnmKlfsrquiwuv449azeVQioS8PbK52QR
HQnDhQ8/E6ZTVudv5F3nnXzq5oG8AK0/rgM9elOb+OeMpHAsKmpfm0K7lfTCAjY+h1wCW217+y3/
44dq8SNRb4VkcHUGopk0SYkYmADORFo4Pf8MB7IU0LY7Rwuy9PerCV1Or5PdK4KV1ogwafwTPhmc
snqMzI1sUA0Uik36j+9iLdzJJPj0n3vp6M1ayuAospQalEt15Q7ueMZn7S8bG8SHkj2um/KzOsa6
NfOQe9ddClOuLflh9W+NtPCATpkelFMKezG/0JCJ08qcQxAnaAMulRMHgiPV5hLbF5Oni600kMwe
+kh/1oclj44A5lbMPM8HVXO+AY08hHs3+9TrCIS1N9FGy8f1YbatM1n+BFXa/p9sCaWfwIsDNLW5
VQhCIVxplzX4Zmn5smfXUMxO+7W4ghLxYUJ1V5jyecheM7z15ecNagyCGnZwZqw6A8chf2TFJDxr
b462eOAdzMi5sPLmed+AhZb6Ns9YMuqQhUJYMFlM+Qw8Q5NMw9x5iA/M0B08hBbzmbGcshZP0/ur
KzKv4gL28Ep60ykjRynmp2A+LHN+uayH5suqry8j/F3EWMlqXqL1IPHdlPVOzcj+mgM71wkF7fm6
LhJ4dJ0wAgNcWghSrOTCeif9VEtmrmUOOgqfWD5Yxu75AUgtU+/YEr699MCSoaEQXzRVTEbFiuNO
4zc2uk17ds7EiUxQaZbKVm9vADOYrp1w75iz5n0RtSW+FVJyVLkEedsE0MMwY5VKYfMoF67n6Lw7
YR3LA0SNrzImwvxago47xAOfx/Ja3GKlvrVomASKH439aoYPkQtCmKbA8X2kCmpG1f3a52D2LuPk
8qpydG84Wa7cY4rCnT0rjEdLkuS4aawYiAnpmOFsHCS3kZp8JN6ezrEBAiDvJtuv43spWSOQGApX
dFURfpXvIWOCTlkKWGMb1rPusZT4rRKiDQtkxVd4OJhtBpQ/e89iviOcyIIVttffGd0sCEf3FYDO
H2TZqKEqxKnVPLqo2x7h+EMvaCxLm5vfLcH1XlazoynWvXce6Iu4iT8vB/ir7T9I1MTNHpDCWAID
CgmmQhan3tmN8NvGWxQ1HgP1O36lyTT1Y2xjn4Is+159Ifa5sfUe3IlkVb0vVO6mjOvnDCFVFJ66
mgfb2BS7DVcCIaIP/lcX9Bt8OpA49Y5kvugJYCDBO6jVh9vNnYq9cVR1pu5UOoobwEwBJUkRQRNX
BIBKP3XP5lbaE7hvpDiXO1efZDnCPh/xkxMmCmpjpJgYbmEnt3FQuSeOEMZksYaWDDFMBrJqANIa
J6PwjdzKWzYvvT2HUKLpdOiRGhPXHyF0oc4imZt61EYzvtDOmMYnH6UKrzeNHPW4T5Z348pFyQIA
db9sDCsB5qJMQ/fD7G9EjBoIAIg4pab8m/LjCCEPEuti5PZrTvRReHSGZCUbw0aJVf1U/7fA1yGm
DX3ZrRqyChA9U5hYJ/3wOKv8obqtZwinFgx2NeQgZbjk1LcI2PoSfVtybP+sUf05ZtBV6lZjhUzI
Gi/lC4904FPlf1Od/d/Z5VMLENzjntKRNMFb7dvNBkgMk+i7bDkVyiOcmrDt57PCQ0Fq6xyEKms+
vEG49MbEX0LiZc8azuUj7JrRIxT4xFVnMeTkEiEJptgntEbAD0h4lEznOfG/6yU24HhbTSJbBtq3
GvPw8j126gvdaUucGnpY+5wFZyNpHqOXt/pb9vLdaUlA/MirYl5Bb3EyKC7c04gwJ10i22u58CIo
wI4y9mXjQCafm3R1qhguamuBDzB6bd73VBce0HJ+54SYzqtAiwbZSl3ZGYtxVFyjoNnuPP6eML9e
NNHF0i/VfFpQLpDyvASc4QTy2CsB22GhHUGBs84Uz9jECZZqEhUc+gFkj/u4dwPTxlhKeZMmg6vC
gJecdZjdfEoZaEblT9P7YlVr8N8KZH24CpaXh+JUQ58QzCzhl6f629t9Fx9YrxE8vq102q9YDogm
9lXNDMNmrLlWvzCR/cZs3jLYXOoul2cODKSP436bH4DSKw9RIuZxaC6Mp+3tPts536v3n/DYQy6J
458Ks9SG9k2UJKLVeOWYby+yN6F4oITQMZaGbCbfTry3u9BxMq+jlBIWT0CAFg5ZfqyxV+jLWiHB
WdleM3UTIi6IyGDtGlvTjIwDLQc0aV0xOlKNMQWuFRHt8bUl6XZDrSFMNOOEcKOUSOFibCcCj0sc
JPEfqEEM55wbPUKrRpiLKC42e0M8nymuTeQgf211OARGGzuI16pICkGgHcpbnUtYO+KeMSdUWZOd
JCQL5Ip3Ar6ai12Qy9YGuCaDj9fdZYlCYdhr7kWwkl5ArTm6P2Pg/YiVaIbRhoum3pSUW4yefq+l
UafiF76s2SMwfFonZKrgmsLudvH2+YeXt6xuNJGBApC+Rd028RL05VA7Dc9UXZX4C9imFQBMWcTA
weKEF2M9mT3LLKg8MX3jV9sPi9TYsECKKeUO/KZcKFPK+/wL6Hcz8zLx1Xpx5EBkaQ9IxEheeul/
YuaXdmLx8pRvJVkEckaS5QZvjkR57vV9qvw3RcMcT/xyZ+1lj72N/H9+RCsKmTXd6irZY0kLKJXZ
Jc3kdiSlqZXi+0UsGsxAdsjkbqvwFzWo8XvhlIrOqioLjxsW8tOcNXkTjmuh0WcDxupAC2PMLiJa
TXWMaOVHyGNyQ3eAs4DZuIRaqLwtUY/HUvR+Lpfigs/3X2Lk/KNSWzhtIVAKCovoBComBqlVNP50
4MI5OBb9/KXqqtPNAmKncMVGIFcPh6osblcxkBpzneWqCw5CY+ykSwFN+jtko5CIWpULl42i/D+/
KyXXkTJOPCtZXloX/3s06kz0x5A1AhXx4EWYDn6bOX+G72+nBrXKjYKr0L59sCe88WS5738BTqjK
jGAP7OJOYpu3HAMIvs5aUYlPOZydVxhEXd8T2EyorfAIxKPrTaq9kWiOAo17erDS3ZyXLc5LpLg7
ydZtlovkbGpe1jWREV9Jr5vZsLxObzWhR5cROQYQvmvqLjJeAwVIwPd5TRosdQRI7Md4Vyn4jLEl
5Vh8k6MsMZhXqyZL7Sx8eyjRALYm48c0BI+n60K768wyeN/IlvN8xEQS0ptvrMQWf8AvE7MuixvV
2V2qnmER53vaLhnZOXoedNjzgYQURE49tny0kVg7Tjkz3Mvu8F9ycvATq0IvpVRg+gp0570NNCci
KtHSM7/o2NamCpgaDQnAMBPgE1OqxKfZT/Pz7UPmHSmQZoszKihiMUlpS4OeB4K1Krt0lbr43ipb
QDm60VM+sAMj3UAj4PS/MMwPQww54f3FajXBueZ0k14ykKFBvvrmFnaQ+EmlFPMSULGlSXvzwgvN
SizUJAsJ/Lv+46g2LLN+sPZT0mzrHeBqotUkkiHB499iICpRYIWkwOef9onCdjBkzj1JyeyWrb5o
8nnFJ9lgyFQahAkBrD9gvuw61PN4p/XVJBUxhvlC6VH+Nyt964mykxnkAz/JKi1iayJ7DiVS2mzw
/0zL06AmQukwp95jMrvDZzQm0BFT7UTnTQXWPCQun+rxYgcnHUxJGLqjCCTJuaG7nHCTHr0E62P5
vOw1ZoTFdbxdp+JvU2hS3eK+BMuplGU+WL+kqVJYuAvTRHDwynn+kduYDJTrcau6dv/osgVp51wN
7MLGd3UagpIw7AGWRThbksNhnw7zLaJLXABTOFXKlujDz9UW3fuDZa2ihnUU9T5/pliGkNwD1/kv
mLlCnmZpg35bZdhJXw/mU1s7zi1J/jRt1Qu5tQyQkLK3ReKSYhoCxVvv2FC3aJbCITzqdY1TV2Px
zCYczhZyfwK240gXLoWydhIMJkOpkernGcybQwRB928Cy5MfRabr5ZJ4bMxOQmgFpqkrVYoz2jud
f3fk4UIOXaX/BpFahRNFoZaU3HVjGZiep0bWFKUCqgEMy1FP8g9pL/Lra1wFbj6ITMu/a+ucovXd
rEQMHP41Wwsi9KH8rK9vMWenu/ICtZWRjdeQMJvwQ7A3DlYxP9KS14PtFWFXlLdXaF3/yO5eDJ07
3UgBlDeQ4JSNMlSp8Cy6v0+2gVC72+CLq1n5vbqnqgo37hQ5/BH8KZSVrrNEIIh3znm2lB51WjIv
poet1JAusXbXBozPRvr7zvTUkTvBs5BaxycuGR5WlF0MTdKLP8EeMgbwzO5gJ3GGFMR4jXG8/S58
SsE4TN6cq7RH1SydUJ3sKv89/EvUHIILx2aT55aCoPXqi4lt8TqpIuYVOKCt4yb59++6MxJ9J7SY
eHtYzqWWZPcYsO4IoGEMFEhMVs1xrf8SLh6Nb6rAI6eF5In1q+u0Yds144e78jNVSplidh/PsGHI
3Pa5uqabTXSiLs7V+1n4inoAzsUvykC8lIEb0aLiB4sUUTWJJdERzrJhkOQwjth43U8TJtlR9xel
bRHh6THnVsGHJYojyQWuL3oZD62cOAupHHfHNmT54ggpfLXaEBRwF/FW3Iq8B2dhesXwBF6WEZVc
wBwF6eazPho18LAziGEOTbPesIrJAhBgn3xMQsNj7AoLf15TqiANz+GqHXHZw8rcYJ0qQs0DBLCK
BeT/AO2ByK6Jx4d0cC3o2sqYodWrahrHutGW+lHah0jm7GGGGXWEMtxuyP6gNRatntekGreNwOC8
Rl8H3UxhbFyL6cs4wKyednE/keNh2PX1VfYhV5B0r7J5kSoSbkCAuDP2ATb+F7/9ukAaULJOZ18v
X7ugec7Nd6VMqff0OQbmhGV8b76OyBMLQuS8PmRJD/aEM+LULfWd+ocqQgMEY+9v2b4OEPhuihZl
tNpTlytn2tGu4sxi50Ekpzn586hBqiKS3ZtgcXcYDUGoZN7jeS/RnhrmyiPMxdReqjzLRG6U93hR
KpwH7/Bl/xDbOjo5J0Y5LwvAx5UPbTrAvki1lBecL4UehAedNo75aNIjpf8riDA103orqMlVyAFL
S/VhHchVTUUbdT14G2/Dy5kuCj68WR5zzXanpPw9zV4AO1CnaEO3ugcPVfu895yyHZeMdch7sFje
udRsfzjZxl6nzyHl1Sk2IdBKtJq8X463tGVNOyFUtoaRnrUoipWJhC9hlciR24dis9Kl1xwAenFR
XB2w5lP94sig6XBdFGo5KenEg9oGTezHgYJPcy8B3s9y5BxDa4r8nHnl3LMcFF9wbUFrsoN4x1nO
uHa86nXNJZNyqUMNrWSLWuBSf2uSytDeBuhRY5FMi/np7hos3xlh1ZWnw5cXkKWktlKKHy3/PnvT
R/2pvbU0wOPYvki7+VNiW8w7bv/x4V5W7/PGY14AU+WduTdT1BW3MAE93Z3S10UCmVat1logVsPq
DVWPpzDAQden0Ouqf0mQmgITvNGDUPqXwdfBCLSRT4VVCH5WOw2FEIvVeeUfkI4jA672pAExLr0o
9TyccFMng4wWDE+Pu0mEHzMHroYqvJkaeDe3EqjEC9cw4+bH3iop4f/9C2eYaJ1AB0UITaI8N8A3
1LSkWY5YKk53DY+TNk/xKd4itVFaxQpOoTkgGMF0n9bwCu9LAql6XdmRIdWfpvF2M6aGAv8Tfqxt
UC+PvBk8F1uIxR6UnGScRoMVn/YQJ1YSJ2Jhoo+2n/9SaOULcEwYi2UjtY0X5R3GoenBePg06AAe
gYYPPrQQPHv5bLkljZExPzMDEoT71BNTZ0vodwBGS5bVmERr+VOtJaw2VFfjYmCXxm0ggtXjredt
eL+3kiuoPt6J726jGgJr0LCabHJk9iiG/NYgVh87ZMV6/FCK2ftPTyXyd5MRx3HS2qWrOvZdgSi0
dxL9di41/WYx2YKnxmqRiQ8ewrg1Azm5/Wc+GHkozXSK6QhH5zrY72HjBzhMM3bZYTC2W8gSLXcc
1UiY3Lelv17k2NW943q9xKMpqmdI5FYpt16I/dJ6FARGhXHDZfA4vVQBoDKyEeRuy2uJNncf10I1
rxyM7WgkJrL7Fp7t0397kLznx95f+W6yA+7MCquWD5E6fY07jSJ6RawYk7J637Ylp48dQkxLfJma
ZH3XxUjKr0LtcHyRgdncG2HOGVCV3UcOItwNilXCK5vb7g3StvL5hlrbYwZImwV55c7wk0n2P4+0
M7Hht/WMMtIrB6ti53yAMrRf07W3kq3ppFp/HkGyVY+yqfhhzn+ZSjHfnf+GWSJThL4ggng2mu9j
hLzBd7M1cKevEncqETHYNGGIAqNziZzQQsHLDEk268xllUnhsBTuMdRWNriH7C4E6MBcRDOkrKaW
iV1jfkpokSBMa/1mgzI6wYdOQ01AR5OJbyZFckukcobME5UiOSPDdUQt2ycaMhArnsYuL1suHUtw
3ETGtyR8bKjUXadKUw1zSM8iUDRiNLbTvCBURzWRLnW4esQhP9Y8YnuPjztKlQRqOiM+NqrwdxJp
x5AEZXj9s9kT5ltE8SI/rPI8uPD4ALl32/h8x8D6mD9Wc71ZmZqdiY6Wsh+S4vcQ1lfDbxu82qUi
Z8MIuF1qpIaS4lWRZFx3g40//zJPrxu9fwd7mHHbjp9nmyoWqNrkfdHc6ki5swF7IOLVoDltyUt1
cbE6L0La9mD6zBUde7RmdBjHH4N6t2uZ2vS4ZnHCKnysDK8C5XmjFlwXJECHOfh1G4YfPq1Wpedq
/Z2RttDe+zaJt360g/W4XqZKpuKPoXVAoYGrd2GTQSNuAUV+sSMmuf5ZHmhGoLL6F/kIeiZU92uS
BnKgx0hMTqlO0jXAtfMQuVeqtDojEwaexauC71aUPhxzi+bvDg3mwYIx7p2P5xVSzZgZgS3h70Ui
uL9CRsId1a4vsuRTiiC46YHWUSVMaOvD9SLzPoreX3db8xTrodAH77oRB+BwjPEFjPZVwfaEJqP9
b5MrGxVVSOqWG+VvXdmVd2J814rbN/BibMKMpZ71/Ewom2URxJ49n+BRBkfTU7dQS4wY+98Rotbn
YmjrPXmR9Irp24S65SFeY/GvPTf9FpzYrd7aMgItFJwUTIQUfpja1KLCwU+rXzLEJUsJz/DNqmIE
hgDUReX/ZFc9O1jVCRwtJdUF+C6dmiTE7eqU6Cgljya2KZiY+/jANgdGTQdnUkZuK0H6KxdwjuYI
ENb6tOPiyzDyZ1UO3Z/ehXWjnoWgk1yc/PDmHgwsvu5xFyHPZss5d3qnQhXItK3qxG2LBtp+xVmV
X/as+zIx+lRblZDoR0doh/XtJrGNQhB9mbNLEDbfOXBZnn5041YmzJzj4w8QN3gbDftBe3goQXnq
XhToTdg5UGbzwMGK52W1E3F73PqE4y927QEjKY5DH3SKSRfHOrCJ5R+BTimtuIqKgyY0cwY8RCbj
foLmeGkqJKRFaz9u8akRkdsj+NW2cAMNAqJBorWVq3xjDjoWwOpGw+XNGsnCL0BfbmzZD8uVg8/k
vk/DoyTE4YIjoz0KrqK0cujwEk/hI8qG+7RMaGBTINVuoScmK3fX7XuhkJ13LWL5uSmGllqPZLSR
AmWD0Y8DM/daAh2VOOtfFUcyPwsl5nx4KIvmt35El2WYfaKJ/6vi0mRjJ4Z9IT36okOS6/6LxLd3
cwsJ0EHFC4AJrGfgo0kE3Xgw4+j5vyB8zNMDUIXbHoVIaZiZgCdduXpzS7TB5Jc4vpi9qRV0HP8J
Nm0kKh2pJ3DTUul6HfJYTVYznR9MhqfojforkE5nSedWdxLqNUMPyAHm7TLvuTnX7yPwAd4S8qbZ
dlagr/JfIpgc7k+EWh1+0xMAy4LeTvK4O84AGl+jYqvZXCvH+oy23ghz2EskNU6ulK+d1bm5TaPy
C4gAs31xa+U0ez/Up6PRwy/euULVT/tOt7qwKMop+ZKHz1qMbh6o4BaRLoIpE+GxakgN5npTWL21
ZmAjuZp/fyBWW9drO+ptM/+uzIX4tvR+LVWQfYiW04cGOX4v9+ZZnDct/xMhXGHwKIAKnJPrrwlN
jGnnjJuW54Q5QWCpKmgbBvgnlaGarIfEmcNcqs6a2ubSvILA76HpxudJNmZ3P/kUnRrL7ENgl9G8
xJ1ZJq59ivKVuKxu04HzaiC7Sjz1S+KaeFkF/60OkfTtg+gzUONYjzESk5ZhpJTztgJZ64tbqhZ3
qgUaqGaoSlo4V1kIpnxzX7Cm7NK2HT/PNDl9pxnYVH3/fxdPzvtr5Pygjq4gnL6JT1orWXLNCbOR
dlpNXCdhw2+4nLrGHhR0v2ojicWRzr+G+2IqZTdVQBzC6+pL/UrVuF+jGDo7lWbx/WYMojKjX7B0
igvTEyXKJLoMZBuAbtsxJH7x77Y+IXT20QeprhXj5/98Tz7dm3uivi0LxgSrjIDsmy7NwzNWdNwk
vLKNTfhVnP/F4YrfRC0sjsnd7q7ypOuYhryLpMTiNOUKZ8zpg8v1cSV9etXiQY+mRKJyC0LV1/bK
hwMxWuqGNSntJPP0Lf0z4CXybtHVy9B3sMtfRJPmTByEmGnsCKrc6Gd8kFjFaa58TlyV4zK5JF6t
WzGk1sFHPCiim9fLayLf6+0PqahFOeN7b++3Z+ug+UaHMkxZwpQAiqYR98KgRxx9FkiGigjglA2k
XYkCMeUhwb5OaAR5s+xzjcPQmZF7mHCahZxokr9KIjWonUX3RcdtgwyD+TDUjWrMDNxqapKfhtQm
j7m++OhSithuTAJT0cIgC3GX1VSmFUZPp4fXUdvgDSbv4tT0Du7F3NcY7Hn+zmvcbsEmRFKIku8k
m4+G2UrrAujR8JRveb2em/MtXMwB2MBRDDLGP61QVn28Kt+Pvbjrm2XQknyk8iGSnJ7hHs84h4CX
lXhGT1mf9RzvSHlXWgFSEisCEu/W2I3/hTWHYnjJPnNQpGL4baWMO4FPb/yHeLu5q/8kVVagVVbG
JXFjC/eUQuURQvJJB+AJYy5L5hEu4kLY0ikt0An3Ri42vHfQ9I++gepSqzoAv33jxlaLjfkLM6Xo
1Exh65XrjbPpwyWtxy5com53OtOsWWm5YisaTz7+KODga9F1BenGa/Gj7AmTqWMCr9ymtqX4rW86
fUmtotBPHJSUV7zLB4+3ypyLLicu9Iqw7B6qUiXGnjrVrUU/BHCfxuXQD2twNtXkhlT4IV7nr4tf
3GyoU4HWnpn8OwX5vxtkyh12ERjLcr5bnvJioOLTFhXLWhjhQyKQgG+LfpNhvyWmKQeqcIylOVto
aH3lpm/punF7g3BgEknFZY+D2QiotzYZ+HXRvaB72nhFKmU/Z2KEGMHB6Ry7vM4k50REbAYN0l1i
wFCdBoEv+okP8ziOtfehlpdNPs84jTgRhoz0bH1E7AKC4J2f0YBK375lowwX+l2jmxMVe94o8hOy
ewj16A8gsAJYklBMl44i9MYBkkLpUggWCCP0R1D3Hfod8B3c2s/JXs/+l6NLzSNiYDae++oSTK4P
e09jW/Ee4NBMVfEeRFeqNguQBUEgI2aBDmhgyflyCTqI8YBD7qSobxDa7QDPl3QwgUd5SmpwssjF
BQ11mse+AN/Lw/YCAcxzmapkMbVrcCQIWowR/Yzfw5rVuUwEaCEts6/5CWwb4YBeAmQcuyKbHT5U
IWaFC5WFW7nwEIZB66gF0zEo38sR+DhN5XqKBJ0a54anFkU+h9A/YeG1GZEo9MtD9mXmRi6s2uSJ
E61K2LLwqLyomoH/+I8plowcs0lQcpUS3o4tJlN2mF8ph60FGYl/Mi0bWYrDqzxdn+EmfR+D8osm
zx0M+fx7qVZV5PPZU8qiUGpZz/YNpeDPm/MXHNuqg/pPKckwU/r+31AZLAgeTR4UcLYU3pXLwhlL
F6cbZBR5IzEUEcVZWUK2xtrTkKLkq9Pcg+0Hn5y6q8XxXOQBP5vn5hPsH337aE/hXoffTPyRXBFr
VeryiNZobgOrZX018auP/J8bi2yU9BvTdFXRPH+POaP/7doC2ATeA07EiS478GS6RBPifChU9kR8
kI2n2CFqnu4z6rVwpQEopEG3QIPl78P2PHysi1QDGebKOVlYJC858rlXgTq5+y8HQnVxm1pbS9OY
KKAvJOpB+hGvKKr59NL4la11Fr+WyJkgueyK0qd1uBUSAUztQEzQ/Av6rRT1AKti4EVLCRM3qh/v
KiiFRR7t8Ust0kzdSwnfm9+NNmI8gwIVNdWpRmH4Vk7Mx+OIwMyAOA50oBO3LAcU/x7x9CaPnpbK
LzbcvQ/sw2OjOL9ANiQe8D+sBQf7qIdXzcibvnlkXkIL9Q5XIAxZdlMDW9p9trMifXIHiSTK5b44
9l3HbyBRh05IHCw5C7c/QpU7zLLueS+LRzKWoqxEKwdclDRtpq4TuyKl0ONe0fIzzsBsFkQq4CP3
7aj/uLoUgiBEY+1sdSiA9OuyZITm5zS+HUvg5axc1giwNNFJj/nSe2kgNTiqhcQ7BQso55kCzc+q
o0VJrUbQp8hU4WMR8PHZMlZfSpZwRQJrIiPF3AKr58S+7f88DM2Xx2fW4VwZG3XXIMh5SgqL9htp
uOH30JecmFGKNja/AJvqCPYDW+iw4pZW195eNt0GuVgBiWJpGN40p+prFEKDvAuw694UDNMpWQJX
VU33BIPntij2zo9LUsAItLYNBcCitBPV0LFzJtXoEeP6sSGq0SuxvTTxKhhw9B87fHbRdj+FiFDi
vOkjZPn5Ogi7EMrdTS2PXnIqTmJf45Snyp4cxRuZDrUkYuaIoLVU/p4qCK1dVcG447aS5UtbHr2+
8VPYT+Ho7KPRk1qwBUIGdQ1tUtqdevL7CdipFcGuPPIlNSzqq+BNJi292Rxfk3FgZ+kwqEThL0y5
PRSQWdKVfqbmMsZFMBw4QpY6YUVZpyg6uRkEpxfdU1GPsi4twMdHImq2KRD9Anryv685bhc8upFt
1uUYuGUwl4eUv9Y4x+TpqnBMyM4obybbCD4aV+uAfB8snu7LKiL/m6xpK2K9ioD20err6pdkm+In
iLUfR7xQt9HQGhBuSs1nhQM0/xZ5pFth/6hVXEDdAAbo/1hMb4uyMi2XJP3riEAxwP85e2pYn0uV
BZr2KgXrxc81aewUvZXf2DZQ30v0kT24Ao1cp1zf50KdQvAw76dOjX1LrJh4iftLBGiymyJUMVxr
PC3l+I7hPWXlBTNHp6Ungqd2naPm3/weQLnr2QJQ2iWmk3kIeKXTo/L34afrRBdXAtpTFxP/c5gi
qnuVNstvJ/sm9LXqiwXwoBVOAxCxU4+0D2JYUw9C7wbyrgX87nEYHuW41adrD9cguD+XWR9/3F2N
jAZZtoKa1xZh672blAxiTZrINg4BNfc0p7y04NZMlxuVZeAoeaf5Zgfn3n//HW8TaDu9IRVHLDiL
2rC5vXlHu+OHYSh1kxQ2jG+Im7VyD3Ge5y6S1kJfQixSvu5rI8cIv8svWh6e/9G9328uwrpP18pX
Vzl5T7rUOfy7vgMuZvzafWbTt0BwgBasxHv9+KNH+RHblLtlMF+tAbefrCT2sUXZLvBFKKc8UIpI
zLTA4xxetU2mBbac7Am63iq873zarRky1PaDoHW4TH/2gM79WJUv7QQnjv6QJjbcX0lJm9b0IceO
i680TJNl965SdNMKDIZiBnI8A0hz/SkBa9SRwOJESw8pYQqyXaRTzM4D0Vr8dAFBlqU8mnxThOP1
9GiJ9VKwHBRos+Slt4qXvikImYLQzHMkgUVh9z2IjaZxO+16aP00dW8a4wIlMTQFXTwso8OVnmhP
2mRAsssCnB89KoM3cUrbW+4As+MQsn/y40u1HaH1Kb9en0O0YcfasvYtOqZg94453hhv47UAk5Xy
8BMvGnXPOqeqHzdbnLWDigX0AUZUH6Mzrnszws14DtlEJwL90cnPnA1e5/5pelhzpwBRj9R8rvY6
PJWeIOhHkR7asJPsYDYyC3an9bI8thIGhU7+Nj1Oo3NW63v+tJ7VVZVk5j9RJPJUIA9vtTkSZOmv
Si1aU8MjEBtSzhSPz2Rne4MTpKu0v/tVJDdKsytcpgmHjhyAJKBdNF3JFB4EAVsJ/uUOpEBNKjjB
6cl1soj0hAk8zTd0hHcaW6/C2wO4n9VBeNrFkUbQFC7JQZ36wOocSn+DPgnBAsE/COR5+/L63swi
A5B8odsUaKTsRRSgH9OVhw8tE8qnF+ylUOdhP9uK1g0KvsatfcMNXwXP+bVSCF8dCm9uxrz5AcJo
H06cz7hhQ5j1+HWgKle2u82xMG0cP9c/49GCGtqv7DRElUsGT6fE0ZzJ3LiZEubOweos+16QSyl1
rxPOFsAdkhS4xHiN9IsOresJxuCDbaFbH0yPZlYcI/bKmQ8aBuUxR9mvcjioOddfP7t48B0UhjBF
gf4wITk8XNhaCjj5zcmOlmJE+rHyn2aNpdSFGNftqT3VZojmhmKkyt5aEnEyhZEfyd3dTBygXn/M
Sf2xQl5j/eGzc0E3UiwinI+Vb84P2rLibt0O9qQThFcPIPre1KjgvG5DSStOmNN41E36Twp7PXKR
0nPHbITd8Q8PUXcjgx4YTMYiuIx2d0ehhhdL1h7G1fLojMRi1CAF8KF+f4OZ4g6Qqk2dadXxC083
lxQGiOyMPLNJJOOCJnr4Tz7dxaRKX2/ytF7kNOh8Y3Zbcj9WAeZpJir/3xIa4KshcFXKbGJ5Tw5+
NBWtWxSUDzTmBEOirPPea5Lq2uM7kji/P0Rkm5CqfMTWrWgClqXS9qTGwJwuqNuPwfwYMNGgmX49
sHfOyiR+ZV5Udq0N7i91YLyTjKL6YBaxNTqzFCkEUK6xjHJkszMX5WnHI1WvoSMBkBK3iEtQW8ko
3mAJLfXCqg/gxvDvLamJRVG6KQZDz50FQGzzLN8J5w8zfVanSAvc4bWnJmiqyPWcU8e6EgMuIWUm
ZlXoEGh0FCI+rsnopL2W7pU1t4tSTlr7fQYk1KAQ6JIvX1Z5/FKQ4owwNmFC6hdUBUMXLyOTzcHG
Rdare3nohPKdrvdO0KnZpNCi08A5ULzNHjM/qaU2IAdLmJxBBk9OVp3nAx9GlFKEr8NXmK6m4LXU
waIfHW5txzZu9MAjNuC0yyQYDvU/MGcKvQII37iJlyWLYKI9oJSw3fRcrOfZdcWPBkOi5BOvZV9j
o2jUbPaGzL5fto2mW5j8jxs/aSiAFP7SCG4Hz0AVxUlZz03/ZjBwzKuugdNO/qBGzlwcVsdkAgIt
bb136UpEQ+kS7NdASXq4DeofosLdbTbPbBtshXg97ufKSnYNLCv2oOHwuTIBOnZGs1Sp1q+dlEvn
pKJFQykvNIqDCet2x6waFRKpS/7HZG6fXxx4qoMObkwCDvNGiczdBVon7Qhy2LU9TyELElX7lmyp
iKcvMNZ1Z2aOJFixW+CiJooZ/W9kO+AHiO4T3jfulWkwes2JyXkXcgdpWp+EmSsE5ZqYBkQJHrp5
VHmeINUePviCXDZAy4dyXHN1zJgrv5rzoBpT78KX6j96qdlBXQ8bBA+YtvGsXBc69HsQIKC6Y21g
6qi2QJzaaTpBaAa/LWArBJlcP5AGylM5gsvgRrh10XE3/y/XAdf3Gu78xFaNIbb6fXeFOFgLPw5g
h2HAWXGbYvfcKI64TCq8XDazFGLdWQXdJWn0PIYhO34F8xYstcGBywPDdfBJ4uWJKTxoSkfwKjpC
rq2UHG38ip2QA6S+zlYXWLfrImzMpdUjwk6exWrR0WB/ibWPJoGtEj9pICxS/TnHYmzoa338os7J
oRA1KyoeRCEAMHR6VIMnv37suSAZq6Jy02mMU3Opgn62yfuNmtggaDnLNVlqoa7a5LQ7jJXyjGce
oEfptR3oBIiKu45gS70AZnOHP0fWYGpC6mDetF4Kiy7O9+p1zeJ5COH4xsSQrUawDQ+CmURWgzKl
yOyTak/jZZsm1zDQE2bFUPqoG/yBxvEIsav7iNPNvHkj7ZSWs9WAlfUPtXc4W4sMW52tJke2YDA0
1jnR/fNXxyTEw2O1zMeUP1HxIaESKjyhUAarCPA1TxjjM5rE357gR7FqWNf7b+jp4Sq9SC+bPKyA
DmEQIZ8wQR/CgHuaZqbIPhfM1VnTMgyxAv1AZ0XSalo4GdqmEUirmO5Ls4hpxQ2KSz3tpTNCn/BU
ZOdz5OqDB5HBV8V4/mCfNbajvFwPaGpYspHpROqeucREXPqE9mmQmOq01dRJ8XlnSNjzSi0UFAQ1
9IHzZ3cB3eR2nFYLvPazp5vRDcWjV9/y7qtBxGdW6ZJWDYr14pnNI29eJfmPdFULGNyP6euCSBLh
RRiSKa47b7UjUMtbd3hRv3Z5SRXEoTWL9+GV0xRjv1TaXXnqTWhKFHF9n6EUYHtsSJAXFIlZW5eE
58V/NhOZ6MSCJUplOk1sfLEPgBilS4BzP7hhPVM1bWudTCbkjbuF45A441kUK5tnkEUT9teK08H0
O71yjDU0m/i02CbYmAXf4K/MXbXJxfcJKeFxsTVC6c39oXR6Ed5rvC9sO+tD+A4PWWBPvCgSmno2
bL5jkhPc+rcI2ujyhNFL9bs3g7kAr38bCbgFfWIrRQ4MQebTLdzd7fA6ED6lsaWDLfa+dbPJC63C
nSrvOCQn/ucw8MWbu65UHv+y3bEJTS9andWUhOIlFMqjoz7eIShXtxsXRjjiAinmwmUCpe8QO5Ko
z898P3jhIRZO41JggbCLKFV+/Pt9hQtdxvcpwPF/LhlvnIhysjv2gupbhCy+203qSM3LwXmprD+x
6jpU2X1oxa/EqBCvB6ik8DQdoHbfkf4nJuWxB7ptxSpOSb4FF1/SaXiif7v8Yeyu/319YZhKfjLm
RPJoljxEaXSo6GcUPv1lb6Nk0dJPm+WzybHcmtKRtACh5DudUmWF1bFRAdQBzLGT6ZwqrnXqXf5u
Aed0mUyHNLgWrrMMpiF8ijLwAQ9dRQWxlGkFv9fXzwWe7tU03SVZaErjeh4GJmV+LzLNYj3NxDrO
nKXtuxvghTHWRqSOh+X+w38K5582HV3/OvbZWYewTR9Zw5qAB+UQFWU727xH7wpeLb8tlpS/gPDY
hDaZHXUm2p3oTsDSeasHrdgX/yXGHwvyWOUS6WV7fSylndFZwE9/XfDEW8GmvCW5Zjo6+BtFKRsA
thKMEM8was0OWKgEIm3sxwCW38OVtwWgK0wP4prHXy9HcSKnjBEuOu1X0TODrIuDKfVMQQ3H+YjE
JHfFfkFkieCXclgEzjTy6oDZOL5HhzgoflInducF7NmrbUbQvP6scheeiNGnZm5qzZlRplgYEwzJ
0qmN2NPDii+kGAg5J4uUh85rny4rqxF7YuopKye+JVy/DEYWdEuuo/FQLk9Z+AxqZMobPXuYC0gh
xNoF3Mvy7TSJpZYNPXGH6+dZhaDR5h8BWUKAnMxbUe9XDg0ZTVtVmCkRZAS7yCBS8ccYOA2NrVzO
kXIBAPMWd5jf48sV2AT5N9PJw5b7s97b3ouUtXQaJG35TzpcS3b7JDo6ifDAnKvyXtiWX/R4lSWO
VHLhs6WoWgZWUgWXr6AdClXBg+tSuhru7cvYGPibkralB0XXH8lEv7rXxW7aRSXjXWs/HmA9SAQk
l8/UaJEQtado7utVHwAGY0Qr0Xxu2LOU/uqjELtvAGFBYQx++/TMpvmmWvn7Yv6A1O0/cYTkgmxf
CV6gKA5shnNIbvH/cudxMUr/sLMVaXBawi2uWHKJh+L3jtb98sh3U6NtDIvTo1JcTfZDNNsrH1Yk
sBjrrDeUPYFoMvK/eC6WMaBzVm+7WD+Jw62Nqj0HnXFa4+e6AZzdWcq3pfc+qbwr/ppBoFKSSd4n
9sFOHUT9LuVfOIo1gk/Muwvggzd/qczcR8S0pQyY9W2p1G7AF+AwGCGD7fc/dIwL/qaZJOApa2Qz
PBFA1sWmpGKkcHEp1rYyJ4ic3MmUa51KuYwpIJ30Qwe2mnRB7N2LlaAXNd26yV+LUvsJiD8xxtOw
ktW6jT1hirJgFtACxDXQuUQ1GToDf0yh++jEHahW2dzyhow1qqBjcIYMsxV77VEL33Rtl/+a2AEL
Fk+ldSCyOf+hk1M+WVuUzGv1Apydz5b4XQ88eWw/auPhb5pmbRKZQeywHxdVJn8WEhIfCI/u43S6
agCTMq6Bq2ogbcJXiqEZ9UaJo1l//xr6hAbSjkqOzkSifXN4D8w+mOLG1puKIKn14WLMIcKqDA8a
4eNH+Po0xYu/BSwdr4k7mgdKVs4ecK63XKUYDF4YTKBuFKuqCyCWedxDZPfMzXk4st/LfsQa+MAm
SOA1xkm8QKeMvLiozA95ku9JZfsyI+er/6eWP3gziKlQRunQZBE59NUfrHDuKpGouSG5Qcs5NSet
KISRju8vHvPfEjmWjII+zJkMx5L5iSNGVHoEp8t47NLt796bVtU8zS+nTPShm3PRB9ndPuHGakdn
8N1X6UaJ7I8VRK/tc+eplUVJeGSjLH50/wXuFOhpAaRd9KrVSNF1NoXGZeX4n8iPji4GSRvh+hZO
KpLzapJwV5WQ0SslX8nnjJURMY+mLcULSbzxNHchvqrOwcdxgn772sp53XVYG/BlK4b406uS9+EZ
zUww41QysMsmFpMn5eATv3S4hLnt69F7fEqwVMFrufHowpwRUZfmSWfAOsZlRsIM98Vs/DQP5Q16
+jFo6onrfjdD/+vhtslcyCCdw6DAH80G1q/YO7N/uicS6XRrYH8t9vPWpvzoFmkZfj9nGnxCYUp5
z62yGrtNW3xsRbpK2FChdIWThyZbuMDwz6AaFynj7FLlXfxmaOMgZIqXr7fpCN7I9EbIiCcWU5u0
X7/FacdC/9lYxZ60nZxmH1BtSZGKL61C/9hm+VevmPkkQgriJo4o6EAGdWVZFhQ8dP9dcSBWQUVM
YkXqoEK6dd769xe75vdOl98Yr8jVTTbdPDMZV7iA4rRcubEEVYWef31Ziow1zxkdV9kKL4E0oLPw
ZN7RWzZpx28fNcw44I2wVS/Z5BqGhSAY/h8N5loO0oZkEUaW9zCMBIaxk24DGXcctlR4xocZ487X
/SoerZlJXX9tRGNuQL9MjnPsSzFotWQthMaW4fw0bD7sIUL1s9lGN55cEjd1YMsn2WtW/4gKNQLJ
6s8X8nsKKK0SPZtGDgzijA3bK+WPkYeDwpCvT4H8Hygdq6KvBmftePVgjINQvIAR5F0w3kc0Qiu1
gZ1TKWv86y/Fpo+PN8dW8NkWFNTHTJKpMKfNqKcqKs1oqAyOUj0ATvfIy5bTUiC+12LFExbipib1
6WkYSaTKiBan0LIb3MHZqEM9R9cvKtWoBEWKMWJaJCURNGxHvV2wDRSBE4B3BgonCjQPMwsuwQZN
j5CrXs5I8D1LZO62YptskkrxgvKRclX8H7gXqcV1wWvuvr/x9pYG9z31uN02fzB1bBKuuZcsKZdr
2XzjXvwuGOl6mAKDfd4AfsEkMy73Ti15KGRQ/U+osrwTHNtLdwmnZYn40MWqOYWmPXbHIa6cXUud
poLwPCNKnnqxOpNsuCe8ih+I6IJAhAGv3NmapqWtxsvlIbSjXaqTkFs+TSKU9DAgH90v9I/YAPFf
Ymx3HL3/ZvTt6EWMW9VYjTbLsvE3SNzdZS/x39VDGAgMKUhWytwYcxELVl+0Mcqx7LfvtkMVmJTO
xems5LS9xz9KxKTxLpdtkpOPAoZCHn7OOKK2Vo5XjePfq1znugVrbgwth0mdmQqiOmfhg9JONnlZ
I9K31AtOJ/EOGWUgDxNVpYQm/30e+d6dstvH70F5YrA00v3wE0TkbBNKCL1HfhhaD1nuWoJjj1c4
QdMWXx59akT5pnFRawnw5VQEGMh4DHgQcES1NSOGJudo0KhqbzMmUvQ9yBYudtAmcDsSfijSGKBT
CvCkyjJvWMa7e5plgMTLP2D1326q9ntaZO9IPS/J8Wnb50Twz15sNSpha+Oc2wIGKWkxiwRf7yC2
Ez2n4FSMEgogpCANN2QfXMLNkG6NiSxbhqCxl8chOr1nc9LhXTzOtNotvPJoKVNafmYNCBxrzgMg
DxjOFOEl9L9Qf5wMQ4pFKzbzC9X03HsKvVdVvoZWISS3oqkO5mw8zpAn7AmIeKRaL5XoXENrG6yc
KsWUBxkdQ3yb7VM8xFS+Ru7SbBgZHZHumP/Ia86UArpyd6RFVHHA1SfpZ7+iHMGSqytpJzuXZA+F
y4Pg2PgEbr+QnWH/5VaAhxda1eLqfrFNbU94vZ+F9SRItQKn1ElG9qSZdzXoqLdgQzIbjFWvAur0
2ztxt12CFOHL0snfUeBLGO2jUOGzK7BolU+f+2hYQdDeY6/H1CR4LCengYZ+IRnWU3gSqJkCckJb
rsU77nmqmMm7P905UgfaUONNy44pTEeq0i9Jyr7FEp/MQDMJzDQv+lgCG7ZwfEMWx7oEOs5RI2xx
q4ScSjE+Bu9Pjpk+MztMePMk+Yv/TWg9K0+KI1nf5b4rSjHG0QIDL3MGis3849vWvLjYeBFBNYWn
mgKzRs1CymwPJdMDC7ELBUoBsiNAIUckDj/fOIONImr6TQNxhRCzEs43rlDBZeVLwvEt/CrPEs0P
3Nuyk7OuzspgIEz5bXPls0GX01qQ8H2A2PSNuD26lGjb4XYNw9F1ib1yiVho3+hwdXcyUCedIkby
XTh/acdb9XrbBIbNMd1TzJ7PA3oKt5cHtQfAcSdIhjxDmjKBsYVZvdbcKXXK/grOdMytZrieQHAs
j3GkOy/1XJrw7Nr1XbEiPBoEEnqB4I2+ydQdqn6NnVocLeM9rLjivMmzIgS8Eh6Q6J7mA2EMPVIk
JYJYX0bJXFYfcTZeh8sx31teGYSXRN498//bGAxKXY8hxdOqMaBafE+P1TR2FEOIkvmeVVeQemLJ
NR49RQ0XfaKXh3X2+oH6hgA+qB8IHOrB7RdbHc7WK3rVM7/H6BhlY+KxHmndLSDaH6nnTgzPvI9J
YayZE2Syy1Ec6BfbmKHHv18XX0RK48V9TXvcL8BWc0H9O1313c1Jt1sJddeerlg9kXCpNqj481Fm
K2UuE7Y0/sUx0+F5W4i+Zy/1tY/NM42DvKi/p6nzX89xBH1h+kQB9d7NZBDQRp1e6fegJXhvYIlf
8EAjIrFyeYcFZEm0KqIOmvT68HWhhdXghC5gaIE7lrwh828aIxkzqZngCBXm0mvCGidD3XEFL1qF
CyeqYGeOHByYlW63zUacOTeeVeOv+OkdkcxXKLwOxV+W6xW5kj/LP6oxzqHDaNSgnGCveCX3ipK/
vyEHBd/G2LptQgujVEwp8bgD4SSklwJiMb+kiUZYe7Ka58b95/f4jyEHtOEInTxcxF9n0BILkBvI
XtenC1bgqPOcOqi46n7zbuCjFp5NlDz75nV5xzs4gsebQ54mshr4Ow0UJ/VSfGmyjsBasGgzLJQw
SFPujWhYohUnC7LjcLCHp4yMNAoTpfMi/+ujF51M98S3qBQioydxQxAGMyAT6k1bg9pgnNcrCMUT
spX3qEGcryZYHHpW2N3i/lOuiWqjsGA0Vk+l8ZqGC+wYbHsJz1Oy+RqyBrSNLNKvI7E8oRyUWpDw
1nT9f+85U1S+Wx76Pfg161IcEX7r7GAV0iiTlgVEV4Cm4dA/4zTGsjlYr3g5ZZkhpr9kA1IvCqzd
UIDmYpepP+tRc+DU/ZQAd/qAHs/BBQrNEU0VgVeJoUnPZxb+DbzJGTKJVAlK4olYmq7boIUr7h9z
gp/OkXNb6OnQWcvkhO2EPmVO3836V/+Rl+4QNMpHGrysEuL4edNKKxWTpyxqooZkwS3jdpbKkjOf
fNd1Wnb9RDEO7FMuxrm9Kq7N/yjmV4ANEoflPGkCwFwHCZ3LTCl/6y9lK5wt2raUPCgZSvUTQdB0
BogDQr8sa+bwBUTLRYmI39OeZPASR1cLNUcNDTN0Tpp5tjNiV5j4j50B5VbGEKT6I/Pr/SZhjsFP
Q4WqysCvj9shnqERu6eqzR7iNtxjbc/NB90WkXyNwRo0sS+LLEbWg0yIIRqJWZjlkuH7THRzbQkE
ibc1NpIO1ExX2sNRd+qR7TjaVMsaCyh5+YlEhZAdvK8wo+PI8RFXMSXShw2pS7v85ULNnnqEkmfr
eh66LqTrcnw1kEM7xyOFhc97DUk4t5ylPPExw/X8cjHs0p9bg0cSrqQk0LsS1juYDrUjhkMfV8DA
sok0j35R1uZxf4Z15RY/5Owx9rbf3Hr4ak/npA9nl61Qd+J/NGZM41nQDzLUhZRAnAeat2QqEAHz
dzWdnPyObc00P8QG6W6pLAGNPnTAzTICVi5whysPQgwEU1bv1teiADTtwoPlRxXP0zb2E4t/IwxB
iwj+tPltd/BLXIUw6qDWhUhwzM0yIinwxSYVw2/6YLgUt/5QmvGXcZN6tTwbDpR/qQZxu9zJ9jTY
a581mL3z0LX3MPm+yh18epEqQqKlgQFvygs3t7CkcDBBl5wMmpnPAo22LmbavA7cTpv4dDH+WgnK
de2SfJD7wYsntWD1IDjUWn2NqD9W2y1xlIk1JQ9VXy46AWFDfPHcU+OfMWZakXXUnsFmgs8EKijv
MdyYhaMvbDDz0Qi1axeiW3ihsxyfdzm1+zgeRKCtuitUDM1yoXyCopb0BXXHBmtft1J2sqrFW/Bs
EzJ7jfhQ/bqlQy/E3ghc3bnSk2Vv69UfPFUh/PtDBzNUaB1P8oAQjVKro1WEVUKRLvjHos9Z5y8i
NmHwWeOruxN/Y81JYgInWopDk+oIZ1cQjca0MrtUUEdYVFxVoM/rBWdjE8Ou4RAW+vlTRduyJvjT
mNuhUeNBcJiA9RAX4OhNMzNYuW6FUWE+UU8zZ9OjqerzWCXa+9WvdpV2ep9x3bhL/wR23hZf12uy
gw3b5V8LFsTq3rwJLakk0RoTBD2kUDSkWgKEAcdhit+c3e/KM56FMZBfImJgqxKLzee+gMUQoP8W
/mmXOqZm3vtVArd5JGbq7mFCYXns9v4DAFasnAo+trhmkSZswGpca/ksaE9SXQPYqmX54fY9O0Ns
wYEYVH3c0kklBTJBYy9/RIw9FTMTtZcyi/QMZqJDulvNNWXmPeZLZLaL0BgOzT9rhvhO9ugcmLzt
zcnE0rs2gkXjaHeXLVeIgXbAgKwtPYlBhPxbDsvqyb2138mZiHBb3TPH0LUa6c05PX18ehb87XUq
vmZBTZN4jjM9owrZWafYrOi/T5sd+fcav+RXUI/cHvNUHfuV7BsqO4sw3u5Of2qvXX82cn5c4ToO
OgdZ7BVO/SI52wCJHknhDRAhRirAUFjQhfKHEsooKVGNzAmEEZgV7qUAK3EIyCUEKg430IH7BEwt
zSasqJ5vMEyCXVrxvbV30AuBv3N+phDWTV50o/vTpWWLvsQgyxu7IeQ42XXPmu6LLLpU1l/z6bsW
FDzPxv5IosA0DZiCi+pJ+GoQaXph1RS+pMx12m7GKumniwcjXCT96X5cNz8K1O2b5YuIU79ekNZ/
2uJNNXOK/0FeYW7REJo6L9VpCMzWhRiq4JLKIBPtRK+7I4gWXJisP2e3I3rrnGY+yIykqG5FmaFV
hDLImvSVwONeLHH6tbyHwdd+GpTyXhDywyEiDJsnnOLjpTG9eD/tLmawNJ7nCv+aJsGAW+OvTWfJ
DZ3fdA2oRsfEcyfWBmGJuVZ9xaTs30sXeNRWOUlvlYxqSUhHXE0InLq/oXLEW2zW9RnFX8zYCmrx
fe296Lo+3RWJuVPNo535Ndwwu1H/74hDNQnSVx8IUiklIHkGKiciyjFJVAodFslzkBDF0cawoBbb
/2lofpbRJH6j/9ehDpiB6WB9/Xvl76hY4l7sNcM8in6zJEWeoFVDDvA8Vtf+uV5ohrm/ZRtGCBW8
9zzaJ3agXZUXW+jA3YGLvFQkRfkJZ4Xd15qCPktNbVlHrVWw95rbj9385ZmXDWu4KKtQJTTTmQiX
+CvvL7pqZby2T/281HtgnTwR3UOVArbecOLBuNSWecfyTm56cFfbrzcd0tnP071RrNH08GYvv8vh
6u50v10Py6JSqqHBxEqpKux2xlBfb2XRry5aw4luIZsz6hXFhlEF9y7igx3X2fepLfZBfvYjSZLb
h3gUQdMjZOJs2TiVNGbmDIlFCUVYbGWnPOvGzyPn/sgPZEXgaTH9a5T6HFtS7WhOV4gfN6ejt4jv
/0J0J53JgJbTanbgjFi05bEyAC2+Wv2MqdHy39FWEKSLZcECua9qYqotCAGDRFsdsrjRHNAQPzhv
yHSrp6reYucYFFjBk5ZsZIWDNr84pO3bkW6XYZ+b57k3EqVYZ0tN9nmLWwjZk/E2FzZaE10bFL+r
enyps10MozfNs+TzSyhx1ppae9cfIvpdDABtasqVRqXw/VHi8M4zPxtnharhdaztc2zzd6IPjo9M
t3jMgWaq4w2PVH9J8Zq0Yr1JTNA2pscHQ0yUyhrLOh+GLo95kHPLLBV3Ah66hQq1XdT1AK3VTrEV
chrz6SvoHpoume+adtzwr80kYtaVNsrR7iYTKssg8svztDW0xSwaue+4+FCbSXQIIAY9tiNGjxrm
z8HHG9fClNfztErJe81efinyYVZd5vZW6ICqh+IR7L7wNt2gR1Zxad/voV6oUUFLB3r4wrFTPz7U
g6PuyeBrKo8lEHAt/g9l4C3Eexvu2qJsU+ovg5WoBj/9s437gepwHqTKgRPIpgXELbJ8vjgF9erU
NdRGvjpgwpIY77iE5b1kkDzRjXya4kEaTXbC0OP6xnoasNxFKJ9Mz60AdPsOm2yOOl/qdL90e1XY
xK7XIwRkOKmAelwop0mgrVLRf6Oj9ECilgiYZl+P9C95bJWhTJJbQoYdx5rUuWWp5jhRJpMJRTBP
rKtg+iFsv0ej7VlfsdZP1x3NJpw/fevLOGw7qFQh1l3pd5AQLTqu38v8CElXWF0KCz+gkHtauQcJ
dn9FdfgBQaQxvZkAeYGBTmB0s649bgUNrflPp3KOnO+ROcUg6ffIkMPi9p867kJwJAmYpNg9+kDR
0rbA9GcZ5WaDqaJyX3tvTAfjjp7XM+2HBQ2g3mnm+/U+BTmFaL1n1c6zZYxXmMGvcjW1oN0/tIC3
Rk+S9OFBsX+yviD58oVvfcHm3YRk+41vN8y3qKPQmSj+3M3sfJTFjItdHb6a3JOdoH1ZVqnEMNha
/7oE72Y5g462Yvg0IDSQp+usk/AP+vbZLDl1wlESeCdpUoS5OEwIzoHHbWIb3aX3p6WRd7Y1S7II
joz11ZN3NaV2hEXLuZ/s4SHv4PzZ0GJdMLdTH3OLo4b2r7V4Wpxee6Yqbc68ok8u0L70optVa2/m
jPBI7JVRGo9eBHIaRwee8aMDHvHoOl4MEmnMF8FAuNkQ++wPi38df9vyXF9xCxpj0sHRybTqtAFZ
XJcpXET8amJydwI4cNNTFwu87FCwrzBjhXR87IE+816LyDYYdgcSZgPYRrbZg6e4QlyqgqNLMIaQ
ZY9h3SR0Zjr3foBs0K6ElLPre8wBvrXW9mzN2jLJm5TzRP5MYzuN3naYEeMgOC5R2aK+4c/tN4RF
qKULCVm2PmFSmzug0epaTK5mlorXtem+fSVDXMZzl0YVkLyMjquewazI+SjvgfeKqWXqsxN6T+25
suZqMUEbfoYLwSOES5uyT0Yk1vJCv/WbrbwTWjpTKXiWdWqPXdMwdTFL8xLZ3hioy05QakWa5JjR
2xZAFLH/CCb2A4lnPs+qrBMrNWuLEAkobeU/swEg/M76QhZAhZscHQ9H/4J8tv1IbmCd2/4EQtSY
F6E69sZxHyYeFoM0wwEwtKJgg34z3OJ2HpMlowXfMoG22t+bKmeIEwAJngSdwhB0YZmuJ6Zs6Czn
I17U7SIOjWTA3Ee0rFd4DHgoeVfs0mtp+64ryBQUhHFz4G97OZmQtWe63ROPD9HQLWnFsZ3OyvBs
/OzRoZLwc+iOfdj++7SKC65/aqAZRPeVIncpo2VoKF5jQEgLvGHuMy+fDJQ=
`pragma protect end_protected
