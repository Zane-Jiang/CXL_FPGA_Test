// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Oxgzh5vOAHGMn6bd9AsDYNIJyCK5nOicDFl+x7CMQ82Ei9ia1+ncHkSIR5iXxbHi
mJAq4Be/O2mHWLBQ72sRJBh/n9CjgT7s1dkfQaOtacwk1cMg+cBlfyMxRMJm4eSx
RBj4nqIori+q2ELlPffRPkbwgA/bmy9R0oP4XSimqBQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 25728 )
`pragma protect data_block
pRGRDnND9DMbA4/vcdoB2LsMb7kCESNoFRjchGe4phjHHwmKsw0H5U+I9fqYKlK7
ipumd2UJ7BQcp6AqcWQuyCrEorHJ+3D8KS554yC2k6CnM39nLCon8gMEC7vqXr2Z
V1q4pxxHzDs1DO9e3dHNOeB4ZjGF5eIwOWl+Ysj5M+w7dAACSQHN9omYyxZh2JgV
4jMtjr7yTL7J4YbOTCR2Bv0RfI4qs6bWk0esoMBZRhmuDnxPLbc3kCtPK1wkAp+c
1cwl6u3/5DxnxZqoWfpNX0eRjln/k76PyyB325iK0UE1HFsHysBlGZJ2RyEPhR9d
XHh5qH5055D3b/lzz/eEb2sMIpydEx7ohvqTlE0JLink8bO9PF1Ok/HjPfpMa7QK
1HXRoOok8ZbSOUP0FseTua1G54i/MVnGhbs2+dLsXohvkDJczs4ofIdGdoDk4eL0
junV6H2Q61lAo9ug5GsCy5PWV031FxdNT3ydpeo/4z7VHG+KNYoFIabOxmJHWEpV
d9zYwf2n8tWYgRHC7OxLogf9EnXA/G1rCO58pj6RFPkkIcvm+CNCthDYD2ZoBDCx
ry8sgQ0QZWkan5mNdOCk7u/kevQ7gtN3uqYxs5VYP2zPkRw0UbR0mTMSt9CUP6oJ
HPjVqbtV5iaLgVl3Zl2VuPcom86IgstywO/18YHJKjdqSQwyjsFO3PWYe1IHICyy
tdxsNrrcTkMOmeuRJqS6Q5+cARme9d+DaRWUpb08s4D4tcqoAG8TSqg7AOiHMxPS
ZuY1KK7WOzMpCOBvSbxnko85KGTaYqk8ftUC5DCKKDWVqArky9KWzD6M9rxOO5EL
zU0+zSfVh+hUMQo0wn9IrwMRjiYBWqLzY8MQ2myLH+cw5wpa1rf2Ujk/i/XsEYko
VOM3bM+KMdByub8LcVih+yQu9JfNwpf5/FEvErsTjjWce5m6Wh4kESbghr7SVjlZ
3mtlynHCK4bbBlwNJY2NehT8tgJ/J6KqGW6/3b2IqAByqEsxJLSl8J7yO8uMBoLi
nc6CAAw7M8YVlDjQtJIZ1izqCB0cRWcl3Zhp7nPF+2pVWJSgV1EEHr0dK2gSv+rs
hGHz95QTdlMKCOQz46lP5+7Thb+3bGWK0/yvYMeBshe9SZjGzG5EHhlxsNqs2JEp
YQox4rtkUsJphRgElDNek1a/62akDfEf0aJYUacp1mjstq/6ud3VCG4rUzFWOSrG
d/69dZhC32uUSE3hYfbOHF01L9ojWOg747uydkzFr9zskjw+S6wIWpMhxl4LMnPD
NtMtTrHRAXdsxWQZDMVKzwN7HD+DclAVTPThwZ42/C9G/Yg5U+v+OeP3elIo/AMW
UCVviXgOAeooTT8jCfxHsAwATG/3f//GeFiYRGwwST2CrOAM/TfPPDSidXhot9az
auHOSoO2GSj3ATbT57cpKXYEmTKfOXPLn1Hy8iohhYTzEb1ojB5F1o4vh4EHBmKV
oesIll+oX5M5PnS8xWLWmjIMXz89pQZ2pmiYfd0Uf7JJtpXV42OYozvP3vrkCfNI
jkOyvrd482CANFnLuKD8qg4Nc0qqUDxf0leizl+PrnRiOTQeDOrvUSB6uJGChP8+
05fCgviUStOutt5Qp57WWme3wYheRfhlc/1LMQQ9mn9jcsXJ0mjdnn25kAM06QEK
tq+z07G317xw0+IMewsaEG3yKnT2DyfPnOWrt63q+wiCs01gLnIS2BvGZ/1+etlo
qad2stw8e4ztSM7OEXukTx4M/D+QcTqq/rbFS9FfFqC0aGpWOw23UQRuvriL2MqY
eAMJVeIxR+PBdYwx9B6AAiI0RhmbL1bH3Rk6Atpv7ZG204N7kv3OtWRXMOdqqyvF
KeZliZ20yJvHAY/mhpKIC3E485bEf1j7MtoRTD3YCiZa0GbF4+IP+22RkkV5xnWb
PaC771ZsapTPU+Ur+VtZcOcWIsI0tJktiuh86WxRye2AY9r9T91kPr5MnlRpqKZu
Fg7UyvbsVVFW4VMaTcEkfTwxm8h8KNPlqAUtyBT7cVJ9WOS63umgCXkskNyNQtBG
pJxE2RURifrMocPt+0KGJLih8ASC7Rq8kXgbQOdTmE3ICY9LE52keSaS5yonbig9
QZ81BbjJ/1Pn5l3eQE4fAX4L2GIDlPbbYTo/n+piu53MS2oexcaIK6DbDvm2F5Oy
SE2aQbqFHGuRr+905BjvD+q2AxVNhowkRfHqjWBdNFbPYAFckKrm82Fs2rMpN3M6
jX2qfzqkd5k40x/qKhfm9DTokbguZEuSaeHGLYxGA6g6MgljfzvFpOpl7GKkf1qG
mrOpBzSWDy6nR7l99LzzhCDrvAkfII2NW4ISTPuavcktX02qI7GSXnDGiWVgB8RC
0tKZ5JOOZLoO+R58aXj1HTQs6eX6dhazMaO+JKun/Viicezj/Pw0m3B4X6JwcUtB
0iy/fc2DLOdAzUBhHA3g4oCBgx7VIX4Q5Yn3juUO0ws9id4DuFRM7ZfPrIoLf5g1
21Iwz7yNntsRZcQHQsX6y5rWAO0u7nl7wNUtg2sQzm7Gk7tlwWojfqUl2+fvOqZK
hMXX1TPSmLclHON/uZbW9BQap/uWTRF183A0liyaUzWpdIZVdDzah1SQJO6su491
JsWYF11LV6IT9WRgTAI3FSgkQlXsF88cyzx/gxM6OqBS4B4BqB09Qy1aMdzFKb0x
naEFIdWZWDB2yHyADi+eRRelEka2jxsiMPJZjxXNlXnqGbTpQ4XXzmCKAnoE+ACH
lxMy1UtKBpxkXg31/0KSU2MOKZDy96wcwGl2EoEmxfAB037PTmGD/2CL3r2dmXNV
xV2ky6J51Sl7kanY/6gDRAhhSHwe99+fOjtPjPRcL1TbfsYMV19ZVzEmFf7JULM/
t/6EqkVCMSbgEliID24u/Hsdp+d61I1hE42U5izhAh1gdvfprPINhebTGdeWZsHD
dp6QRN/YfY0oGevEwAHiu8todufw1aXHABFbncr7lcwp+IYlGBPPd9HGhP66Fq7F
mXbwKoEhBWGoD3UdwT6BCOXLFBqtcDRZWF6Mlph5GjCaTlzvImZe1dM0WN1/J3oL
xCWGOmEMPgVWQLp/WSjW+E6Ktz5pj8AeQjrOrfe9G2LXcxqbrhqsSP5qNVl21jBQ
hav1ks8kEeMGKMyn63BqVwLhoHTB8W0h9mRo/xaZVP3gU+oMlN3HaKUQRfXN5e/s
buSOLFa947YRyyvfpN8xay2WVFPZfInMr2Kg9NYA+AtxFMwrQL6iv02hPBM9RzNU
cIwvjn4wk9seNwI1+0B4IM7S36WdxtmbN9NwMXEtbKx/3Nol1lU2FHgk24+wJDk6
MoB5ONistz65w9iMX28N1xhe/ov2xxkKs4FUCvfW/gBrDNYdzgPg4Mic2Z+S0CoR
SorcurCudQnOxePhL6zWxanH6+vPraqgWnxBMJ/sffzAQWDeVu4xNaWDuGZHDou7
NRAspqFYkLrQZ07knAm/CP5b5NSDS+/JWhatu4U4m7MdoqlIGbzpucrMwilChnph
1gckzFJ0evX/qz9Hy118M9Q+8y8OOeA3XMGhTTHLGBzleMuEFSPgEyyCYKStB8Bb
NfFUjCtCpcU5JZVY7CiLxo8LQYvxpjwhvVFnUeyhg+1YAyABMIt/FpQsBxn4NzEN
m2vVwplkAa8CKjtw7VC12EA71HHDDAEid/jMws443cvkulDJgWehu2x+ygkjAut/
m7qHYaHHHO9y4mk2S+GZLgZVLXlCbmeObX4pNqPp9+2i5Tla8IP1yckNXY/SEtif
L7HanJdsy+URkG75LLmUwpkvDpx2BWEcZSLGWxP1q6OTyIBiIuUdvdrBiAG+gghC
LYnaREqAK3Dw1wMMw1lCeI7upz2nT98I8fagosqJ0+0SbTL1OyAGV07EiyMRRzMr
4q8CJQhYWtI6lgXUk5apGB8Jv9Ut6rPkaeojdznE9ZQrDcEAJNOCHSaFrOGimZt7
YWMJtqx+H6OlkyOrz5GvncH7jK+QYEGetQt81cW7thJIhI2BY4xxJJ15dLxV/K3Z
dUKmEt7S7j7NPCm70e5hM2jfoxU4y7kR3rUofujyoejXDsHfw4lyoonq/I72cMfF
jJiqXnipl6c5NmV9Em8zvJhsQe0up9ynafneTK7YdDrlmsw0HnlyYaCPbSvww9MJ
hajj7c+ZllbEAXDu+Wfs24TPyF5VHO+51vHSUi7S8VT5+LtYqHaHG+tP3LG4CNI5
8ENMfUGpF9eTrsKfJcvk/Zr2+/Tl2zXdDpHUD5vQq5mbft1BaZ+d4A1YnqTLZOQd
P9DAePUluIC26OQkewOmcQORKTfH5UI2x96sQx0jooGCfXBzdF9wuDe7Yh4qCkJO
ujP8JOeb6TUrqSvDHQQqtvDYFJrKtYsMAoF8T7ilkzr9IaqI9wUKaV2Z17ff9Yrz
C+2ydhUZq9VyDO+Wa5bqcxjsrAsl2Lm6Mxgp5s3+w3L9+tW6HlTft3MOqwJ+Hzw9
SXBsRuOBGqYu/g5f1YrKU+TgqsuVTNn1mu/Hx3IHOTRlqCVC34On35QZggt6USFu
qGty1lA8Y344vfQUDM8PuBNyx7sZgpJfj8gNFH0/YdmjEXpuFWl7hUqZCPM6B6b0
caEo8ArT/kbKoUmqH/+7/l1Wkq1WknOqpMi72hsq3nevPnIjz8i/1cSKIYFUkfPn
CZgZ/qEAZ2t70UvQRWDb75UE2+x/mLfwWn9i8w5woHYhiSbyPb5MCpJX5aVSO+hW
0JI18pN1sLXJa97RVTqC43+yheeyetd3yzziTLlhnUN5aXrzQu6uMxfxm9Ohf4Ng
Kkw63dqIbxYyJWuiuRvocGf8MVbWpsew4t8UI12O32P0XQrC/BKsIRn52XY0XzAc
bljIDmSvSUyy9hTfArpormKywEAPoEJDu4GeWQj/mWjg0f5STyLVyiE99MvikN82
vduqklGVTVVEFvKgO6CngZytI6eutlYfgo1Iob08fOb7hz/tlBCwri9R/cdE96Zm
6sHaNj+s3zIByrldoGIcDI+0pEw6yFuCSAE8/PuJp+hLGjS8LGdocipp18glRgl3
fe0i7DkHp90mX13Tg/CqiqW/P2++DZgN6Jn9vcImAv1CLN0W+1ooytyqk9r/BJdU
RK2Pgau9OPl3svHUmzKu2Q0Oy5r7bCvhoO9LOHUbX1va78+ptLAo19XeGXFbxyc1
p6rjWn5DyF42fqVDPiLpIOd6YwIzlO/OKrZCUwNEhzi2suZun1JVgB6oLkNsVTfm
ESbqgYgBa333l07hy8lEuzp4dR2wNMgEjAOqANVuIhFbfrYCIFW/Y5KWDFvL528j
bz7Z2L3jCli58U2YQS6Ttc21gTqenm/9ZrYAU4hqSH75rorBV9+lYCeK1AGvCp5W
k20alQHnolMSiM6oAppM90voMUoaj58Yizr7Ta7yJ2eWC+ITQCvfCwqwQiG20+ZN
y7AV7Up+rOxJyZfCijHy+QGELcCON+qydY/E21+yz9OnxZujhr36+XoP4jUQr6dX
4waRDX/26+Gbkg7mV9gXcqNIHhnV877tykEpjRLwuOSXSuvPyoxkz097pVlJfn8p
Ik2tyWwYDMFf/gpiRar6FTVuv7sc8cza0PJYNER+kgeQiVdOuQm0YXfD9Dd5gsxw
Dg4kq09jx/YuSg1fqv2YSSEQz9y3jj5FZl1wJEfXo1oDrTt4EzavkijneQXdDu96
X6HSkCsQYIp/qw7O+mtOVdQk2Ou4kIhu0CNr/F5uKL1nSWr7nBVMiK/lLNd/ivEG
QTTiLAF1QEKzQeyEgMtkwuzsQ6lPpM7zxBTlrkd/aFsYfvSBAaNzFrJjKI8a1sl5
gSUpY8RcwX//qX4xatz23+7CEkGrIHIySFYpTVfQa7IU3CLBAvWMw903OJDdYJKA
EER8bkGz/z0ts9UQpRYfwX9hodlT/neSKqZi+UcvI9e1h9baauTf2dCYvs2I1cCn
kNj1ORWivmsbKYzFZW1cXjelkCBICS3Nqm/zdovr4AHWyvh6d/7K8WHink04Pbr5
qkxbEnUnpgjOWhp8IOkQBFg0rpCsnyMEQcRqmyDEMzFKXfe5FpwCoEFthCScO1js
m5EDEXLYyTWJ13vZSDH61RGD29jmhyUIl2QhBN+Jo2hNGBPV/2Ix9jBOIhAhyybp
4WOAwAy9Z/5thwtfgsD4lpoqmU8/JfdqbR5wzheOHrhD2X4+ldMx4K9sqBf0Yvv5
Pyf6E/PmZ5bQXXn01Rj8+sa5Pbu5U1LeAsiCVTEBKn94pf7T9WRqDlPmuElacbZ9
F+wbXuJE2TLpw+4uHgPkFi0/EBza1V79AyrsS/inKl5yBhtGQSZQWIGJTPwLF0Pb
g0KsD2lzbLcFLU/FgncpGf0ZqdLPehvQJDjGtTF2qcQk3pKLR3diEjVuIryZ1LzP
S/oj7BBlM+Re1SfNRJjV6lHI8HeZwIezLXHdBwhnXtNpuxeOo/Hkf705Wo9H8e1r
hhOMZGCA/sGvi81wqlpfXgCSNtF22Yn9mfsqKFlidGPX6UZC803AOk4wssZrgeAX
tBuIJ17lsUEt0YwchwB9Rd3iqW479GfIEseClXauTGLpWV9WJKeMjUD3Cx9kCQ3U
ERPFRc6NXsejS1RZC1m0YALUjrP1pmNMPEXzCIsuFm6xAlDvDLJD4esVpctJFaRr
jspQG6m+qVByu+RsAldrEN4ixAXP3nG+CUZNVSl4d0VpOfCnx+5yMr2zomX9y77u
pSCNYXtYui2MQGNdp8l1J7YxfKPn65WDFqbZ1kXIHD/05wfnMulXZ3scjz2Lkf48
zCjfxCeQ0RhDFbDP8ySB4KCjGYNefYYXmUdLvqkKLsp6jRMg44Z6M+51fePNiUkI
aMHKvR/OuF9Xz4s0AiEyw10ZMQQdo7bjtqWvYZwMokKUYAiG+ZZGGzYh1dQplLpZ
Kv75FVVwmrOhHWvgj0a4IcbdjcUx2Tjf89i1A6rgvPUNvziKApYtWTh/eKW7LhKw
JSIKscEiOb05OtRf+UvrVsg4W6iwaWg7QBhKHpaAG5UgjCspK8wspY01IWl6+eeG
SCDrUgricgKJEqMy2iLwC7Hr2sDM0BKAFqUuTMWppxZEne+L0zrgxQjIvYUty105
T2r1/V3gMiIADlzN6sVliYsdGP86sN0tyuxOvL0ueeZB+1vLX/uCbyWa2uzJmVfT
XiJy+ZodGBzWHJSTUOqPz9URc2NCfL5aBvG8azKZXcRenMf8srVeaiMcgDPpysCe
seniSC42rsrhQgdLRUtCH+Nui2zDzXKQe7BdN+bIZRg5mwD7bPY+shxH6Ya641vn
RkrUslhEPCpfk+ZW+y4JLKUd6yRzDkvVZBmbVEaEtcEImnDTQGmbxAi6PxM/F+4A
lIVtLLnQnifFqO1pFX2V6uG++1JyIv5JAOiNrmeCVSB04Te3CF/9nWwuUbQT64rU
JlTr2xtw5GaaEI6KTqMreh87WypTKS6vwTf5nO4fzANubjkL/rWeoNhgGjS1RzOU
sEmhejkHBtDn81GA0zSaeocFJs7rvd2J2MGBYL48o7fndteRqEHDvME2FRGE3hLK
s3+D7oAnjx4xNkPiHwHPZMUqQPoAbwi44vNCQoDYPgEQguxB1xyiVvu7iAoi4TY/
vQwRgV2pA9Nl77iIjEjhWZ3m09js/1gmjHPyopGofxyFUql96L+2qyQC30UIchTl
A+ciZMloxF1UE4CmirrExAZ6XuKXFA6qLI4KUG3jBxMTUgFO2L0eyYCxwhYunmTc
4mSrPUYYbc6Dv/ULu33xTUuiOSnaV529u4oCXXzlK68YfQwqaED9oQJpnnQmVCcX
HQX1ptverzoV7FhxDbp5XAOxKrPRc6nGANqxuyoLrTEkPmcEPmW691aeZSrY0P/r
qfy9ojRGsZVSZLVAHAp/VM62zYD/edqXm0MY1Nipe6eUvtWnb9D3WTzJThS21ij2
SGp+hGdIrWfrF1knl5K1U/nohXWRkzhccSub2etgrlv2FDG7Y3wNcCuiAZnEXsJI
a9P8AP+kfkxrH/7c5xGV14bUrtFKP8kQk609+k7zYMNS2tRSFk52alUP/qCwEH5i
0Uo0QjDv/ytnlpwfxSoZU4ntIzlVMwDGX8FoDjY5ryjtZ1QRqUAnFnOf97dyMt/w
p9LQfY5qljrhsrrWGngr6VCuU0vE8T/cNxlk1Mu5H89NodfTixchiVDROq38udxj
aWShgG5UqFRya8OWhs0KYFDNX1hBenF7jg2VS3Ek8KBTxrfx7e4fktMmM12shPBJ
tprdsItjz7zrzZkrRmE12zvyOYtvNBcx87amhNyoq8wykBx29ClgusTibCTeIiqv
zNOiwsFxdqFS7TlJJOROC6w72o1hIFlic61hIbPUOJMe9i813xAm1TN0jLSO7GcC
vHstwR+4X31St4TTTVStDLxP86hpvEG5iJfeJ+8hBALtYwq81lWLpuHhGQKqSZk5
xeXm/l5LDwPsFOgSu1eT6bLyYGAMh/nBn5iMjCq7IjsaVWfxWSVna77H1OSA3nl8
FZ/J2BcJsBDLHY2R6Z4PE0ZZQ1RI3N8IzGWhw1kh1/5zpMuHRQXnIkaEH6A4trVL
dJDEipVDBgt4Z5UKdV8yym8swnBL5q1BOW0nC40S702u0ieRoLCnGXbkXaXHAJNq
RoGAjYffK30z09GQsPeXvBznN1B55gBLO0O3Fqtq/iBJEQtP7YQzR/Z6NKoMGXla
VLQVnkoxSdCaWQzqI0nA+cXLlica94wLI+EaDZ+L9W3tPd8mR7K4sz5InOMk4102
2pqXC8ZjONbCGk4b3whY2y9Rq3Ii/fQni7KZprWMXFLj0VjETOcek/fBppIBxqSz
Lz4JfDYCFPkq2cZl+q22zSW5wRDbhFLs0nbKd6K0FCA8Dcu49TTpr97iJT2j5N5e
G8kzMRKflnigaWlt116nqjXgRliYDOr5iLah774xoYMgkIb53ag9Mddwuwiwp76/
E9wov9BjkovJkOXX1824fF4EMcFGT+Ga7oMqerTwGel2fqKB0kZpLjOfJP+a9gqq
qLnEEMODTD6yB1fqXMgyC1dzswjaX2Hc3pIEjY15hnNmffnoTKqzdwy0Vb35OGgY
6hVGvp0RRB67DGLDqH/GZibyF7g9xRjXWTEGCVlhwOVlHWTsLc94RvOGVaEB+Bar
gj6DPaSOn/xilrYQhxyR6LaF9bzYAr4kagq5BNRWDCw6dc4m8bgnwF8a+qruydtP
SduwxCu4UN049lGdJ4xUpcC5twHUdSQsGr9nE+tvkuFU5ZZ8SmyVzyI2SOD6uaEy
lWVcEXBt0lQtiLUcUahIP1IDsR8nHimVFjVKgmwXlkKrk22IY9TtffTLPHC2KOMT
5pg+a8mFJwlept/LcDhw/teH0WZgNVnLXO4Z30ngrJXSuYw7avM2lCUzk44gHFUL
Sa/Z3Ln6Y9qBAXC/rY1f8V2QJizqC8wjozg3GsRAy7zlE7yetHvYIPPX80HtrtZs
fBNSqJnhBtwAsYzbQ98tH+z2VNQqAnHLdsqbT/O7e0SIjvIPAWIjC7hMYs+M7Bwx
9fDLUoiWfCaQks7n0RyW75vHLkI3FIbFBby4Emh1sAm+Qq3INkcZbDA7hpBkAc3K
BZHfqj8AcozezZhEnt7vaXITxFTCL7j27MxrGBrXavoBP8za4/HvTNFySpPnr2kD
/JySo7AeaJq/Kn36UY+TAOPCnfvFP0kl6YQqhopB4IJ+7ssI2TsrxZzoKGhCAMyS
lDu6okNObPa/uSGQ4LjCammczc44+91kFMdb/uOjFvYHp4u6VZD5BO/0+PHUDdAF
OqBlQLmxNoLpCt6o5kpntjlVCFdZpJtMmYRzOgHkJ0L34zDR1taRzymUU+vA7KhP
GTlvifhjtmiq2S016KUES1p+jewU/swcLX2dSyiCAAbVV7F8VFH114tx71qB8ZoN
PpOruGOn2XfVnBAGRu7rzFMVwPmKAUZUjEh3Yov2+8DlfcOQVUsRzZYS+rBjip+m
N21adhWY9g9viCuVH16G2GE+cEJz73qj67GSct01EENUkZM+4yZWJ8BybNydQ8lL
qY0BFlqrhMybanBn2+nrKKkRa0HmBUITUx6Cr/aB6xknpLjHlRykLdayI/KZcqfw
pFzDkPBwuPSGXggSYDWd2mARA/lQ4h7oH2+kQZzWiDoiOFRtr/j9rtEdR2t3fv0s
LjmdfPg8cOY2S3Cp/QEiHKqG6E1HucI2sDQla2MmNWCvNVG/owl+YO3nkAmeAivf
BiDCF76GZQplCrOcqIgtl+OQYw7uubd1CzoPjcVdPGlCDN9nWoleHSSbaoQsxAJk
i6cXtpj4n5bhn8WiJ3/pMALo+8bEGz5+bb+XxKopva2NbgEqe5I0mo6yJIMR1C6U
ZGcb5Ma/Lc7SzR3OiZkTiU5MjURnmHC/9FNR3VgG3AOKOlBRVn1MtUvbShLMfmTD
rHLFHrhcJ5fcgS0wTmQFRzTrxPMJWzgJA21p2gjRzv6mB9Xb1d9DjA7e5gwxOUJO
f6B8vBrCikilSi8IZQkIyJ3N5eqGOWiPq9aD2B6T9yuoi0ilDjNdjvQGKEbWqOwI
QToqaN23PqZs54WI156xDFY3PMlUg4/f/U8wrccigXbPwD4LwSbrXjXEj24gjtoM
Oj2jNmmYeyCg7HmEVw0vd39xIVCs+IZl6JXTfgNT/Ok92l4oraXGidiPFdG1fFi/
5oFsmGVL3NFa265uPusBNM3gS7pOMoMv+ZY41AOcvx8iTZ9UCwz2nFbnvPPDDz0n
8f7P4RY32RpRldq2sokqirMJvXuJQARdOzw/Mic7j6e0kKiXt2Y5n7fY6vp29nc3
TWvZ3bKi+C+Npx/0Ea8o9Z0eGw/pY/AIcCStuxZ+KAS8vls+BseWQIT6FpMtdFEB
6kqrCj15TKIYuFtzTlyyGylcQH9vyHc5qumu3DSprFpVVJ9l4NGkybBVQSHDDqRY
tl32uDs9EANp8U623AL0QpN3iUxBq79SqY6jm3hj8Qv1UYXqD54tT68rAyR7qveS
Ub63XcHmYsnxGL9TEEl/TAyX2y3LHQl9DS8/gT9fQcy01IvR7DvYOUDBU8xpGIdX
Ti3MWbmULRK4XTrUG9VtokW32ddgZxg++YtJX0XNOPgj/SSuSV0sEOyrFOju4M9y
BpvGoPASWtkFyzP4JyYsPvmMV+AqTHfJVcnYJn5w+2jY+exrqGno+vpWAWIfG6Ds
teKR64Q/nU+fxWXmWGjiglNfxvJlK1aC4EmOj0NOdhEKUDDhnmA/lIW3HG0XC0Xi
CO81N4sOuYagCpxHsPQ90cWxZAxAL8le1p1Tm+/XH8NQzAZ7nnyD5D+qu/vnnMEJ
99FVeERP+4pCkFBujmgnp0exjyu/pIcmRdXkRFcvw23/LMiVWpu8wLkBOY4dZIm8
gnF42BrHzLDOzbh9Jsqz4iwDSMMJOipp8k9L1OAm5JKvWFALnYlBA3PMXlnmFLtQ
S44RJ4LTnLxq1venavcF3wJwrlfvzjx5rrHVTl+atMEs3Hhcmt2IFLAVY+hYO81x
6QRgnEjDLsl+q2VZ0Jam0ohZG6DJv7kUvlapFmZbSVH9Hw0PlvfYHYFeItqyfhkX
e3JRzbmMPuqWBLayzm7GlJsFciAxZe2c74TsDmcYNHtZcTM7v/GtNKIUUrsbtp89
mCQQXC2pOb2r1/uSYoh7RqWgZXMTXfTP6wwXYYsD+bfukqtsSID4rrH3t1jwBNUr
h/zpiUTELHl8PX9ShIHrfgfKqgfCQnOaKu1SI3UBK3ycWoMk2ykdKf9yUqgpd3rC
iIgiC0iSn9+opV3D4MQ4NZzYv9ZON4hIGugT98jOSJk09k0mPie41NshjHJkoPKl
vdr1dlX7LL0Cxj0H04A51IlVLvH2tGd3ZONraNpv8j73n6WgOAka2GhQ7xMqQ1DQ
U8wgn7b4pUFokfFRJ+XYm4MA/12ZevCwVOpc6vfk6PiDDYwBtMYpOl8zTZpgJOgF
VkdDCDVsQs7/ZHQNPodFBuOricbcwrLd0wY9gb546XNoxHLUlfW/S+zmTEZZ4ha8
Egh9PlmNl3LfwQOhcJhY0kmVQP/XO+HnM9Vq+lwy0TKCJqMEmhOw1QYHTFLBuq+Z
PupF8L7n7iWbZV5BsG+f63hPe0M6upl112mLENHR2lm1B+Gv9QGRy+CU4NLK5Ihg
a6aGC47Zg9Vuy0eyxTiTeFlqtMbFFugZRgjSOo15pYBxeSt/7kvXftDyYUZJPLhw
4xD1tDcLj0QduYEJmZqOJQ5KAt+xCOEc3vCQvdMeICPcYa9PGpL8zQsOAwGYgCU7
X5shufVfVn0Oa4t2y4WriHnYKTdrhalC1HdMEBWbfZIJ896u6cT75SpLYqkHxrPH
2WetcSJGXFhfLZmkemxkVK4zKnYErYl7PfCZtuYz/ghHEOfcXGYJj3wRvTb0Iklg
NEIZCBBNSrh0VcmIipD+pOtRJr4TFxBaIz/+UDzoxmGUj8x+3Bivqxes3id70yng
RbjrWprBY0CPJPRq8t0l/ckv0ridbsapTAsHbPm7BhisY4pzO/LuCxeMOFcWoQDS
54PjfO3W4PpG8w8py8dew+bVFWLi8MLtn9tKUBHotuMhWSpNf1E5nfAykfSVXQ2a
mWIhNaQwBhvgz9OsLJchU+PMl23vG81KlS7NtqhPDUrnj3IkfT6/+rL9Uh5XH8xE
f+g4v1LjXe5WRtgR+lnT+mwXKoIXgbMrZLSWYk6FIPWPW8KjjAitee9UhIlQfX0I
CyE2VtnGtUHLen/9ekwmy0jcaSQlKHno5QI62bOD1hdgey5V4RJ8n2axXP7dvEHu
eZsMiqhcnBRERNLbSPHEWvIh5KpbUyj2UoJLZHKimNZoR0rdeKbRuM6ICIXnTcUv
ep8zhVCxrbtujet6T4O8SA+46DzyvArgijcFQdXfDWj71PYGfpsjCPHxYYen3RoF
sJpca1A+XuIuQSQxZgvJ695wsEhZTGXg3HQZbDPQ+WmKYzDAzYoqHsk4jL+161DT
N+aPCfEkRvk/ypCCdvzEcEaRNojmPteU76g+9z9xtJkcO3fEyQFA167WHWSR4DHR
8vsEAObjkspRzrr1ddfzSrAIB+8h/RLxOlACnP1/JqZ2TKzd9+CnsN+9lX/LOGPz
sFbMuJSA1X8vaGXPnkS9kyRtFW7Nsvr6RvukuL7GR4yJcuVwVC0VTk+4pzdn35F8
Tjd1uNRf57/+kZqRmWschbr9mnyxyJ5v28Wwxwf35tUAxYHy4TSXIphSRX7jNPbB
rH/zFaf/IGivLxXsPgxngOWbSv/QHZE+2VyHrk9KcJYoxI2xXKFuNerq/jcPAugA
fk9/lKKjVkj0Q2XogWHCbLm5F8EFvi7ssje8CzZRLm9Q2yOQVgKiECJPFOw+0l6S
/alhhQvcPtzVfRc4E3efZAoVzX+IWatpwrU5kJKskzGAxn7PP86Eo0VDRfxxJsck
NUytH7vqIvEH1bGvgjf/9R/GrzH2EdfWU/Q7KBFsYlR/yElDJ2aIBhfkedMZRyMG
aSadfBTAN0xeUUFKnE2aIxtw4NsHU/lf7GTBOOf4jGfR2fkl4CWDXO3pfn2sEUnM
gqmbBrzy/1o9/BanCj6U3eH6ukHf8BFY6D8fe83HkSmxUK4hEK91KAVAubuK9GU5
mq+lrvbeMAOjZ522P2kWknUN6kNR1Nejk44J3z5mJDX/5LD4o2cETnxdWWdmDfQu
kKNbojzQRLsxiPuA3OzUa06tmkrwI0AF7kiqJFPg4XnMTGol7A23X3do2tBKU30X
VqGxC87nXA/Kqg6lIfmTkHqq2rVzZ4kifzzQNwfQGGfahKG9NLb2uLMxiYaPxK2h
zXQMXTfsu3Tg7zhvoV2Ia8QpnrsRzTTcHdZzgIJWrRCI251JRW8ABP+p8HrGLl9m
yo6wyBiqVmgGRP2CQ3joKEpDXH5odL44pn5llzYj91O3yI3YEQe/P7iKC0cwEofb
mqFV8BTd9q2xbRVqQY+LL2iLyUOuFam4Mt7zPnsXGfTH53Uc+9qJkmGbgVWR124M
fEobWDxp46MKs3jnHqI+w3b/j6eAa7OYEM6u2b8nlrX4syZvtrcWAz9f5cHCfFhu
J1HS5Vv0BmNbkh6q8qRaLyI9H+Z/QGU8SrwjdOGaPrYfz7uHcIMXQ6zYbhuvMfXS
YPE/rNx10hFHQrDrtvxXHr9jPiVxTl0/82aBfyq7X9DbbRYJN07EdWDBkdx2q37f
PDjo3oRtk/rtjrwxrSmJjX84/FOgLxj/ojvpDjR3yTsUEahr4reKVabW40aVOZKH
/BRTVFmMFSAvii6GA0AdC8Xx2AYlercBdcR0ZUHXICkWwAU+zYuV9N+5WdMGQh4c
tgkBIP/zLtXxZyE65cv1voJJnpum5gMkGWPaTRru+5sT0RSbcm63EIBouZ+cJa7g
kCcFXDYqiedz//7PYbeRUxd7tQOoD1BBYgiK/rq6El2uROIvWRJx5QHoS2Za8tTi
K8zT1VfDa/Hr6KkFdmgCvfy64wMtMyhPwP3MCWc+yT1PkwbL11lF4luAM7f/dhpf
UySr8HxmOltEtqYUbwX8MeT4Mi+q9MX+B90+Ii6usKGDI1xNFlB90x7nsuK15HjW
rcoGFddiad0OXVCbZtlZUu75qr3lYQDgs96QWZkHbYeOXn6N0Li8t3NXeaJ11GTf
9JeF/3ldwm6unMAAkhwlkWOzoIiBke7Mli2IiYXLZDXAZWjthYIAOxmuJDOCWGd6
fD85h8dPrjtav6/A98wCMFfJfemffMbse5rGljfLQuK4yVSns5cb4Hv+AZJspImD
yy6pAAEjYjwb8bBGCECZ5b5IlJ5iKkINvVUeh51jJ+QUx6FjDCxD+isSv+TTOCm+
yGvXr3TVI5c8lIl+omak/b4MTD4n/dzbtV5k/x36hw0Hrpahyhwru9oSOtT1N5Or
z19rYL7zX0MZPIy6ssrM1AkBqaMjnsp7PQhgXImoulgbICnvdzZhLel8bcaiM/So
LybYCjz3jA5kwfQvghjnQ8lAQkbAVaXGnuhmeZKnrVrCccjOeleCnKHUE6Ca2w6L
TFHGmm1k918s89lGxjlLA3N9pM+Te+NA+7rJcvmkuQpWya4E8bX2wEPX4JyBIQWp
Z0vBzLOsFdttdJxjl3ufYJx0OIYdPxdqSH0LFUAZZmlDF/dTUTweE6NNL3M3baKG
iOyF1X6/7BN6tSCMLbpLpm+Ld/tVrUk2xz72jyvyyvEwPHltuTrac52ms3NSJJza
kHHMYHWkUoSg84SeoWOfUsHpsvZhBkGnCMP9mmD4jOZsrm0z+MldtfxM8FG798zv
3sIuM4ZcKqviachYqQscrC9bIffxGrmz58N5hk8VGCZXXy/w+BTpkJIBKUAGl7OB
7Z60bXoBwiHLbF4ruMyfakKz3pTsmunm7ACwAZpNu036ijv0DCCsUmRV95gmqbqr
mCq4hsS6a8IHbiMIs0njmF4Re9i6oDtD+CtQVhm2VlPWFywKJ0Mv5bHkR1j0hQOg
2SmESa3KtiVBaRUlNhb2iBWIfJj2Qbtx3buBNaMcdYAFpVbtDsIS1Cny1RPoth1l
MsmyjONyPGYQLA2pOdpXO8M4tOVdeq4lWNhF8+ZvGZ19p9OhHVaKcjwjxMsFptYv
dv+lofFMPUDiXER3mSdxzvYUzmcEUyxa72b2UaKn/VDfSTgElPmifYmF+HYY1Q8i
25h8FNvKk2CNRf7Q9ryIk9TVRHUlve3ZtgN3EALXeFvAjUXcbVDUmx7keZ6M2LeT
DaZ9GJqc0L39Y+1m0jg44NTKj6A5hxY/dX6YVGrjZy2+BhSC+wnKmkjsgyLD823o
F2iseYP6sfVhL93UW8HRgUPZXjbSRb+NSYkDGMm+sm1myjwrSD7nTIseie+Td+66
HtFuFiaEkIUbmCycvjuFpX3FqjJtr15muLkP0Y+LCKY6g0lcvDrCr5Wt0TDkZjhn
zRu/2arStz3MOfK989vOQ6phLSXvMxSoS5JbiBtv17QpRG0qqUGm95DcCnEEANrg
8D2R1FPw0h1CvUxdJq0eg/+YqsoNCezgNZ8FCfwFsxr4ROeNWIn8wOmK1T2/6soB
egDOEPYek/7elhRpfOuBuqTQ0vpZQAHXs24PDwsv89w0IFYEuuwEoiEZqOuymQst
WVBmVBuR6NWI790gxudliF2/nz1l/FqNHhrFj+dmxWSzLr6uU6wlgWWiXEjE2Clq
0/fqBKY7LSLZD8kxlfz5CbVQQ+YjbouxRWSIdLlvANpux1YeXAaDwsCn4TQp0CIZ
YELQLqJlTSUH5KicsfATAorYSyQUDWsKeXFhDNHVRRp+LXME+X+Va44BtwPY1LhZ
XVZxnpeQbt/5dZnTKk0npgGDmvGBGuyCAaInPrU4glR6Fe6shji8B5i1sFTnDpNG
CsNEZ0BRf0Y1gECOHss87loZ11DShvhVMGGSGqlGGpHxEqdplhwKFqNrneDZT2dN
0xPmBn0Ua2PQEiz+FlDR0mKZXU4MfiLmLRW8L6lED2vOvf7V15cdLmNOBUrssyN2
QAD+/hhPUJfYGdwRmbenj8PhLno5nHo1PUjGLCnk2ptFzPgGNfDXdplG04s0j6UA
NQPaIMmJVBXYwTtZZJMXek8W/VVAg53Gf4QdVs5eK9AzWOsfe0tvqwLidA1kNHMY
RehYb6Xefp1OB15JZ5qrA/tpp5U3NezBoxRo9+dwRy8WIU5d22+DplBBdcEkhqY8
5aT9Ws8R+OdlBePSa/bp1bQZhsYg7Q28UqUYzCL3g1SecsSuR18Tjar7qVMpSnIi
8dTrya5kZZpMAr5gzq2o3Aawse0zAxk8mCmExuahzYeDsONhreMxZ1qdzzbQJ4s7
fx0BshtvZZ/klnxbJv1DD74DLtniybd2uepRDkPFbVPOaQzfWY5Pr0AlKjwGMYR2
KKeahiyZI5gxHGn4wYrKESZqklGPQd5JhDLHylW4lwoq3rH/qW5hBTEhjwXgWAV3
1F5s9yiLcRWYN09wSYaxB7ophMMj9gRLPUs5T964DskKvvdmUdwWBhQLD1m0g4W/
2aWpIvux2ULaqPoCoX/21gt4dDYOh5MQnnBG1ZD+Hd84qR9iYPeSC3wz1wtZJibY
00zYwm+ekM8U0/OxDixG3VvWg4aPWxMzifeA8dOKDzHJx7mW0286JK5dk5qt6gna
I3XTrGTfFzNhzx9Np1lHdk2xYIzreghiG4jtBGiENqjwdgjd0GOhLXkutVGagsXw
jXcrpBLw+jUGIWRsU7AO89xsB59iCis5rIt8WH6SuCUMTZiGsN2ZltqLn4mTIBiX
aOFv2adw7vBmTDcC9MD4y4eTQVbHRPUo8TwGA86Rn0eCrmXqULWOtaAAxCDo1nHS
hJ1a7XQIx+ybMY9RiMLARhg5ZJokQX+VjDQ4YbAjYkSOXkpca2ZMtLg4ZiobUsG+
7BIV4EUE0eQ9vVr1VNw82zqetoZ/v61vy3mKKhkKIjOg2qefyypm4OERo7c+M5RO
t16IkjhAXbwG4vx/Mov5KkR77RXhMQyBNJ8Gy3lL3gTQ6TIxq93Q4qFRYEO3Ubz8
XvSEY1LQsiOqItpOrc9VfxSmOKXN+e8w1S3MhaB/vNuf5g7aJj7hsxZ8DOucVRBI
RPWCFupvdqW31J+Pun7IZptrLcozBTOAnRL8HNwwu9+cEDPb2d8r3zCD6MHy7pOp
Ucco024j9i7A3BJXQfr3n0hwqR+VPW1KzBA+AXaJ+zUrnZe7Y/yUYz9Ahm8aNmDP
hJ/7qUq7FA97tcDf+5YyQExAy++/QKZlXkbBogSa6MsHnwgr/wA3Ip+hvTRAU3um
xMXu7mrZ3Z8OPbqo1WyRf6UeFTWOtfCYU72syiveYIbkwWePr/lOtFMD3sDytiRi
wWd3DSUmRXpshunrpsYE8ek6VinAhnAcsqRvBsDhqabHt+HUf0DQ9ECNgJR1iWS1
RX3oqvK3Vd2u2EOJCGX7nlOW/IzZcGP25TpPAxt14qDhD0Oo4BH+JgDtQ8szrusY
7Re6qMs4BC8P2XmsKZmHzt16iVixJWDUsgj/g1E4pG7t8+kmKLtr979WV+s1PgKc
Q8e7it8gTZY6XR3eN9CQsxWIiup0a3mm3Ez0yapfZPD2iThndZ/gAsxWy90qc7Lc
2/ZOVrxX0foatRkb2+C/+gXjNGfeSm0IXCRP5sdpHqE19DaTqHeOeuSj++Fd1GXR
kNt3mpG107LmeKg2aSTyuldLm3xw9qWMdEaqBHYmj3XMrOspwa2QTFydWI4nd6xL
Uuhl19Epv53woAtq575WwJoz63vV3Tw11/EfgiJkN21j4pszqZnrgFcUQeZA9zjM
m+xAKe463uB7r4MuniLlaZRzKScDilSbKrxJuNwNUNpYAOOeW4r2y+lGoBFm+cQh
O7Z5uES2m8O0PL/wJZjT0y/DYFB0wvaBNvDFyTHvz0UbU8UEBKhh4uMRCsRS7ZXu
lJcByJugZfvyUds/bKf8unCKMcqvZFpTWkKaJgJJr2q580nV6Czm3IJ6A0jSQO4D
yskoiFGFGAdibpG0QTjXcuWXY0MRof0/6VzDRw2DHCeBDI5sBy3Luo4mW8AS/sY4
sUf8WRd2yMTSJqbV9ofRZbtWEd2Y6xIbBVRX/WWyngv0j9bZfVFC2xzm62gcsvCd
ZHzppNn5Gv8GszpzML/qPur5BgouIusbwUWr0f1IOv0PJp7Hqc+lD6KcSclvVVR1
sckyHy768IBxaQm8vcSUNFaRkxfqPpd2AcBceBge/PLCmrsmee1Yx1iQhYbmg0DE
KVOfVeUtpCzmP/8I2FYqO8u+luiPqqs857AYSfaMof7sJw+TsbODRbGhHduP/MP2
EDXwkQxBXlVgLzVthMZsrtGKnDIUY8NdEvWBQpi7jD/YAqVIAA4wzZZNTpm5gao+
1M/B+DgDQ97Bxs/x+e7UKunvOiZAyBJvQMoN4oPlgsXlK2WwA3gUCBQzhu9xb48E
WVQQm2UVBDVTDM1QA+zF+MpHQu/of6W8gEwEJnnKBytCwQXoSF7awxraV6azLTYU
o2Z+Q3uSacLlLA+QRXq2u+SLDoxh7l8WYWuGicTav81+lLduIl0WRRBFcKB+CW4M
eycHjbnTPjoNajz/4N7gUn55W1LniMuUkFuQDYNdTI2e7isdBkLHFPu4/aXfEnsj
MBWaifJ8hHeUNCBDMOSwEhjooI/B8EaSbSyDtyDe7duRQj1ZsVMRqrtK0URtRgue
gFs5L0eV/RlSUPoqSCq9/7kwHtQ/fnonbX5yJGViyMoGjFmdK2eog8GwRGIr6kPD
VE28Olmu9J0hSggJp5yVlZjhvy11QIjUqxanZFOdQifXJPg3CsHvys+u0j+JIqBD
35BBEQ77yvq1qb9q+mw5Na813t7Eq4WcuDXL7WKEhh/afstjdxP52J52qs7tUMQQ
LaYlOha3KpqSPpDuVEY3uJd6M65kvqQ6jXfVoRKyffVtVr+Kl3zTXDFiUUZz8B6A
wl8lMCWW5z48APp0xkfBcTzuqwp148HdVukot+qHuSPRPqoYV9jybxYsoa+H0T74
ttjiMhb8D1zxUjwuiDKPpZ6zbtOtfHIdDnuajH525G32bzcyfkOw5CiqbMkRj66Y
wyUbsTmIx7+oLTAKKIUn5kWDjBMLEfFzcQsJfEwFi81K8G4g1UDxfKqPin8H/Qbp
N7hz1Iyiamle8UNR7uraV4SHxidx1CvfFs58rMr//Lou7LnBwIQyOASh0svqQOg2
0a4FwzNkMeMkN2bugxSunjP1PEit2jK1emhkSlpNGPgcaO3V/Pa4s66jAp7EKidx
ResC1m8wjmin6eDJ65dpYbpvjQkHjUPZupkG7kruY9MV1+diUWdLuc8tKMaiiIfA
9a7VeApM0UEc245H224ztojqGHsiHwg414sYVzenOE6juEJAw5RKH2Rl5HtHU/3f
OBCcwZBokWKa8vfIxZU3jBnREmEOmlK9eGeWQ7crTbrF4BgB3/OmX46frrhhYBwt
zxkBS6eNtU+imcCxxOZ7No5mVvWLYffoX77fCEo4jYS//plWN9IjCbI/TKTfa7ta
KNxjND5hlEy720rzzSIReixy+RusqlYRqLciyKThLR2N3uPMxkJ9+psYqnLWQqAk
C9CdHPACVPT6a0G57MEEfad9F3UxBASMbzy30PpXGhHbN7pCxoUpX5/Cja00KinJ
9hm9gdXN2MS/BUk2Y3rnUKeJaFGjYUgCUS4mu2OPKJZcBSGebKIKVYPr+6+L5Sz0
JLtU0k43drF3TFrbUaTn7L3jO4g+9HH7GrNjtKUaRVWugBIPRQiGYZV6bHnUw3z5
B5z942kIZ/GO/GxvGyagab76omWXhmaKP/7m0AE2asv53nLFDYZR7OqrbCAiByV4
aOfYUCUC7Xzy9F/VCZyhYMB1hauJu7HP8QiVS8YaNfy1Obuey50dKYtDEiq+KHqH
BdHoGqMQunHeB7eX/i0PNfK8wk4KFvcW213ezTRHdhiHsSdBwuv1DiTJDInnHSwB
DUdkhMoaOYQme3HFvKtQFr1JzpNhOKGo6xBmypnOoryRKaRkDl4y6aqqaW/b3Xpy
blXWXhFH0L7kkbjKaF/IAT+AaqNBi7fhQ8kuFg+VqBzXCKF+1jzLtACEjWtt82TV
rPU+O90tFu4zPfGNENXMKUBcoxgfP8p2OQM3y1tkW7Pef+3yyO2J8wjiu8VYU49e
7oBbnkVRdSkEZzRn3SqqEe2/hbtUHc0gRDd8qf6h0C6v8RT39HKYDFi1SHzOKb0/
UmHYM5ftAS9B+4sfLcLsxsi4E+aG48XqFvFrC9tVxqoxrV4bFIH2VVFn+P9/sgj3
XSB21Dar8tg3fwWNEuoY8Ltef8G/5gxTkmIyDwsF77Lg8xPoMcOPwalE4fRskDUV
clSXdzVKsrsAa3lIri5IwICnFBYPYQxL0AYSZi1RP7s7wqvxnLDFNikaWO3SSAFa
aUkNJ4UrlrkTH7W3gfinJwRTPochOteZ/Y+XJIso09Bmip14Ael+/HuwHlh+Xj03
x/Jb/B7ybHoX0QiYAv9V2A3IDNbNfO20yWJd2y8EfutfRQJ76H9MOSXcZU+oWL3j
Wa3AXWq3CT4mBf495r4X5QdfmKZEUfHTBARDx8NjkzW70Rk68mwwg5GXVCU3muH6
zODfHIxezNHA4xWmvjPFsplhAmnKPav4k/6wexlwmxeZArrjDy1Eu/5In3JYYrtY
BzCWJqPOgBQG4ov3YrMfsLhSyFKRP6nJfHXN6Kv43GiizuWyUKqJLW0t1iMgx3Oi
KD9i6JYLdI0N9e2zbnRpjUY4yQDLlAD3WD1Gbtns7u4egUHbIZP0WaNSNUkrD3n/
G/CIuXXlJfRIkMMdxhzJv77bWCRcUbOyWi/4pYDFubjPcwVE/9puKKrYxr3N8JhL
yMfcukI9exTr6ysie0HVpTCdp1FCcvkft7oXvPymFXFe4xJNuJathAD6sX2eA3DH
fgyTKsvltvPh6Buu+Gk26Dhqx5+g9WmZpPUN/HvXsd+07Qo9WHS27JKwWmAvRZ+0
An9XnXKHd89/tyxD5g15PdnhzI8mxnwg1qfS3oC1a+CJlXHIxOo6IuZiUwU8jQRq
e43oOKrhYsW+md13uxSEVI7bt4GmRJOWuhu7dZX0VprZE/cgL1SB2PGHA+s3nH4z
gV8ZC+Z/Bnqhd98Uysaw+DXz/H/zdoeg42NZlQJLE+QwEstO+0DAdIKZNAjgIC6p
xnCoLN9JSa54fsNFyKgxLHFgoiRImh8m26YUBieI/EyvgibBonFMAmE9B1P2Rqym
YT8jmeACQMx3ouzWF2cyBNTF9a/avUfT8W1BxTHBHMO3IdBDiPC1Vz8+rYV633WT
VsByxsULmw9DsovKc39t78jvL25kZmJS5YmspRdpnTReYG1733vwqlEu4lGUA8FT
fdJa+zFE8FQ+Us37e9JtZeADsGJgwbRJAkCYAypWgRyARPKY9UWfCmSnJw+1Q13t
t9N8gAMaudFxA9Hs7UJA0ESe8RSBXapxMeeTx3gfZ1F2p5bgQR4E4JRe+URRNLFP
U338R0qE1+msq6uj4QVumT4WFZVNTdcgdtT0QOmEo/6atZ0BMiLm8XvEAYsIudSN
yOF+KOzIOZdqkXjcApGaF/pDYhtNcQAUCP9Jp3vcvZvLxZprm8ROASSuuVa2Mgpy
DBEV77enHKTeTABsRVGX4SXVBjHH64t88kuBtH5lPTsiAbYy2BxycLJ72UOxtrLz
/xjdAUSrftqrhzf/zt2yxiiMDEqFGn4ukbcxU95/HLundyXMJ6vWqgt7qG49VbVa
xuxio3NjVOAzUXYUk8yToi33KOMxwe8nu92Tlt4saJgoNmnaBmylt+oWs0lfN9Eu
5+HJqWo09wDaTkl3BGHA+PjPDkE6AgWVOY1rsV0SjNLuxaO1JvjuQvwAQBwXscdn
ipsjHjOq37zs7ARnflz0tHf3xBy+S1zEMbQB8e4YZlpT8PKOu70buEfRSr3Bcfnd
/AykxiYL90bnX6A2eMd2lNl/pgnfddGPjRyRTa3z9QjcUQe79kvDUJ0XP+aqdXOJ
FbSRdydVPc1OYgU7grxFZNoIdDdepAI4iaZQryayapt4zCipGlDb53AT9WyE09BB
a5wO3S77o0HyOBP/7IxMN5480zHPM6eD+PWEsPEtHTye+jq9neo5zSXyWmwzkjHU
loo91Th+bmh5VO7CtaiUfnzUAM5AyEbyXPyDIhja/13HRi6rJDjd7nhyJpg9xOA1
alepSe+4mcQ43JG1ltb0uCXgd+vRU82mrX8LIlEQIRwUJ+0XNzBEOUdaD7OnIenJ
xVtEWEg1tZ7kW8AVXiR8Zgs61hUNE8/jTyxtXI5FlaVlgqNmC81+LNPdm+7zt8ZP
QnUbAyEYlK0MVU1GUpSJkwcMemO8XoGULf4A8rtJmhgBIN0+JWLBIPg40XHQZdmy
RnEYZ6m16lAo98Iz0flO2nQb4ig+DYowDkrMZecVzyxV9jMsf/hvDKrj7bcfX1Dk
Vee/r7AiQ+FreuFDgPQCXzCvXduju5F3ucHTO2FWQuTMI2SrPZdr3A0mOukCxo8o
eHO6szq0AvqdfdeHP3BHGreL/PyOwUvT9tQLSOIdzxpjNO6zRCg8HQLHe0iTnmAD
BX9KCXnSl6oeIzAGuJH01en+EqFST4iCTIKoYF6CQGRw0jdpt3kxuNiPGomWTcqz
t7Vroovd28chCPHe21E6v85IwadVp3wslzqsO2e73EQP7m5tXcVAnYGbzS+R9yW2
/uPUkHaqs1d7wsYtoW0N3SCvEYMa0Znoyur/4koX3iN+MrMV6IHOaUNOqwoCMOt2
OsdxNABksAcuM1r20+C3yqiLpopzXz4x+vHexnvFpbnFurhxIiNg7j7ySvKdK/xs
uh9oRsCLE+vWknVu1vMj+SBUyCi+TFCzAb+oI/fD/sqS3mDO4geXFrBBbKlrSoLk
F7X42ppvkDy/4/7yXNTZBJ0+LvDt3ABrewRe1UTc2iPdD2nuTQf7M8TvV7lJcH4/
V4K/IDFfxw8GdZco28OKkJr+WhF8Z1p7tUMTebadK8IkZdeEtXM5AFF3/5zRO5bP
g5Fzwqz13xzGsNQ0S9YYs9gAbHUpW9mVHCYr1mwUhx+eOgZKMaAxT2sxxU1IYPY/
PrLp1ByI6KJwK0YwQzelmtvZlZLt9sbvyFxr0sVDapgKwoIfWGqlkwZpYv6g+VTN
Ou3tfhTiQq+By0g4hoiu8T0ZO7VluPLQNdYhu3zI+4vnAOxnVM0qFiMMvRDnGR4g
AhoA2r2Zu0Wi+FCBVSeWVLRPpp9EisxkhzVwLYfH9HYq1txkvEZd/ym7jWhyVkJI
q9g8lTWUqxL59mDbHU4ivHXUWGelTZ+GsaL5kV4/hEyE+jBdql2HbCQgKVe/s9xA
z4ILLb6NoE0vCqyy2NMaM7pmAfZi0cYUJvc4kx6dRYgQovOqM6jgtRI5W9bp0OIG
tkfdJjukQCYW/npjWDTBXDjKk3LILdU6Ls/cKmRuCr+MKU0tQartF4JW4I5O92Nw
VYK9VET2jGsi9Yt9fLRxoHgLwFi5gcho4pXIuTwGRG1iCKmxxQrZBtM4yuK1IHaD
OKBtZU6iZTnHfKl+1SW5Bkhmg9WX+vXUttzprMP5i331fEVjrJco05oM0FBLP+oc
N+i9uwRLTtS31gjbzkqvAyqItFw+rS24YCecUneSeBahzFIPiViS2o5EsuYpL54G
cZ/Ngdu3d4i9bJ4rslVx8NtAVOztSpCvfwwGlXc1fQq2zB639sqc4VQO2e0ilk8y
QblCuidrseswpyEesVJCO120OeXhFA9G/ZJ+Y8PIQL5R9BuoREfs1T/UGlUsZ9zs
mBto3CpwxMpRiM9Fsl3CjC3jn+QS6FAx/nmcDXtAJLyISyC6ZLsqzuYsf1t0Wdgh
7RZnj8wudPnAwR+KV1ONv+QaNAenH5Yo+BZ7812bMiH9RYoq6NOZ6sUqbIop8/Mg
n9BWDOnQMcJcXz3cbMr3ozke1jdi3o66MYmg/NYuBl/W2Qc3qBcDGPbFvVAA2C3A
hAMg4y3mMF7qa4QmOli8fcFjyny+B6I8o/HpqC0QLLLRHf/ISdV/ylo0pY2QR+zq
04cmB13tnQHtZ9Kdezac7IjJ/8AO3c9aMSz3SYw9lOJVNntyBdst3gz3z6NoqZgS
Vx3JdPhokC/uVBMQkxPT45SVUEIL/sVB8F9FzuxmYKU4Jy72JFtgFhUt8nozwkWx
nfX/q/BfLOAkrhtCDI5k4iEz/ZKlluyG3Wt1xZIsUCw0gGJuV9xL/pPWwT7Hcbxu
HZ7EzfYZXeYztnVHLSEQpqno3VngXrJG4vAAmuRjeV+u8ulKHYh/HjtcTBk+EShQ
KJosTbHolDlfzG7glYdXJ/iSszWqEF5Y6TyVzlU+T6tz7Q1SQ0NY9qIN0qlxuEKu
cMMOyH4d3KKA6qf0swzTUylbKVSqnK1gnxGguUilOmywzPWpBxGKzSC07VsKyCnv
abh6LBFG6e37/xJPhWWQDRdxUygqw2naKtSJhhsTqyGhVUmd+upbom9880rk5ooM
HCYuMLNcCuK07l+solxHmM0YDS3rnjIZTz/cxIph0c1hdYQVBq4RyIt2FoL/bEX4
dNIdHAaKonuw1XNchseCBOwa2789+iWjl4kxZIPYetL+fxLFhZ3mwepL2yXcQMDk
/0jQ6m3ysJmnJmnrqjc1oFiIFBkyCgHRK29GNdxnoAx7WlYxpW+AXwllWfN6fHCo
cF7RtW2C8WxmbVFJDYzZyY56WMuYIRTWm0zLS1vqVygeN36PWODL/ijviO7+GS66
aapGQQdKceZKFEySHYQpyIXxAM/vSjjF7+a6SmR8UhlhvdbKKqk7HodTopJHnkQr
RJVvBYDxOjvOPTujtpZ0rpxreti6mdIHUsG1greF5yU2P1a/tjZIhronlUOoT5jH
Te11hR44eeiz/nF1kfQGN0Bn8Na8ISDoZaAcnsjWREqOKyzWdBSxXUU4sLSLpGSR
M8yR5K4KEFornBqTRLFLG3COkNuKYlX9wJ4eQWxS1ceyFeKhLadVFp/Gf74ayv4j
0yX3s9xOMhUfzloLSl+dB4s2eMLugo0hixoXLPwco5hgv9mcZGmf3kNC8G5+Nr6g
zqgDMgAsdMO0+o/Iwxi2jxRVV6XcpvoEub36/C7ejYBWoxaSFk01L1w0l+4xpJMp
kpBwkHUg17OGZK17PWVSumHMR43bM9IAkwgCftwn5qRY/AAuSAroP7LZxa5GsvxJ
PGU4B0BTLPdCHNFkBxHaSYCZkTtdtZINc4k6bDeiWyh3QpGHqNlUNfd78Ieh3EGk
bqU0U5+MBQ50gnj8N17G9eEMOiXU4TDFhKZDNY+hi5q8HcxF5LXsyN4lwDmAJMiL
MEcvS0/IR35cw2f+5NYnSe7t73lXTNWbiwQKehytCvEZ1+I7EZPnyYhWF3/poMhs
eKNbD8fBBf3qWcX0TYFUMmWJ9WaWzzwEBC7pigg4xPyHmDeVyeyycM5LHfTqpNl2
Ncfsb/eGMsR1Hyiqk3KvXgZJBUprNwNNdpjG/Mt6gkAaokkqWDPlczWaEj7vJRHe
mBSFyviHnC8SR6KKjQ3ej7MPrU7BH0ahlXWFxfQpul7JDrH9YhK4C2jcaE5v1nDl
y8QHc+ifpiRYAVGI80q/SoOpaaGG0OiOch6R0C2tA9YYhn1Aw3kHdp6nxfGmU8eH
pwmPL/VZU01JUB0a6R29jAJFwblAozJwz1G8dwm77bs4/GAFQtf56WjbxEH9j19/
VBkywPv6znmH70tsmS1YQqW7q8nmVuy3hKiKrAObvmjuqmPDipu+Wv0g5CXbM8d3
rXCvtnlnDPlYvfiLQQK4alE0VpjLpCvHBNd5JYunhHNJ82PRRkF/F55pFN0FeQ5I
/dt7QbWkvx8vF1UmpASt3YmJy2wmAqKrKAIiiWeLCSoxgO3SroVRC08wKQnTFsJu
v+CqtEw7xifdXzafAR0GPINJ8tQNR3UlqQByiULMARJPWcva+6JoWBO4J+3prdzk
vsSE9nsP8HXyE9xZV5Y0Fz1hixMqcpQhCcTAXYOedmkSt65BGyWdWjGz79Rj6iJS
Kc357ddCd6WcFQoNANQhoACn6WMZF0uKZBzujCf2PRi1rhYXvmr1zZ3H9w60RdOJ
rzh/Xhn6md9WL7rWJp0wQyxGMeKuUEdMVkWhL+0Otmp/g82LDwIhFyPDdaD7isQa
iduRzjgb35zDT5UXTc9QjzXbtXzh3uUdwxFdoW7GpHA7VnHyyOCfz+FUKWdfyns1
4ya2ocn77rgk+5rBpl++tgKtQZwqT8vQNNNmZnyTvjr7b5KGOZmJytmgPn4p5vAd
KFwTwnStI8U+Za1WO8AH1j6GuxmFNX1wtLpK3KxjitDktNOQHG/bcy6AeterSBdv
WmgQfUJ5LtTVnD73U2Iq5Qa52p4g1tSE5sv0zqmzhAypA+oqEBHlla2F3LMk0UMt
kn6Na0YkkNYxisXe22/K1ZDn2xQBmoiF7UiWkelTro94DF9FTY2nFj/pk4X9PvvV
HqcX4epdSJE17oM7sLMb11gvbO/5KrEZX7vGWius7noe647/YNZphC6K3Ih5y+A8
WXSQAQSyRzP5ZeHqC/sveZmVjY9V/BePYigdJ3UmB89U+FuO9h1/B0FUS2vwyv8p
L4ogPhT9YwawjTjW70q3YLydrcI+Wn2LDc0fRhYqMiwPfRGeuOldm87SEBTrvI7X
nsh3untv92w4PW61qv9HPmi7kd9yZNJvlN7CVeMAHN5YCdFbWeEubhs/UNy5tCGC
b4dvpUj3l0CLqKQN4s1LRFd2D9+nHbvh2rLzvdpA1UnodOaMfZrBDd4edycKnIRt
gNhiiYZqdFX+U0lNy6FxeSFPjG8jI1Oy4zPvdqIkmOCdw4rP0P18bN6u5BljOrzp
NV9gmDeV7KBOgP9oVGP3nZYJn8KZ71hCL3vv/44s5va8w2XARIB2/qtYEwY6PxXn
WZy5IwiYWApPTXYRcTA+SfAgOo9plCIfbwKiuwYZtsNaiFsoFb5a4yPrl+JYa18O
ulxoV7GjZ+GjLRtcR/ssVwYalb+TQoqfOEyQ9j5TF5tIbOqxLm+h1QfI8HhEnLsh
CItQCQ3FcSWB3dVRaSknj6c73It6B3JhhvVxdxMs03zTduh+AlO5prsjcolhT/lg
Yss/VkwlYnwTbH8Mq6mzBL7fmcjJBhMX7zoXRy49Ym7xnoc4424CQQ4L2QNZhGKT
Fm1UzpsIAvWoN7M7RWU9T9P4kYi0u1XPbd3DgllnM/r+OtDF6alrNRsb4MyHZ7tz
h2ipILiZSM+DozUgjUxNrRjMjRs+cGePxzCvL/2nOnJbyS2W/mavPAB2kiybk43P
1Y+Iof8gubQucz2CeFCARIh/5GXXs0OSi3TZYyMJW0n5Ka00Ll/4kOjnFvcEpTQG
HIGfl5GurTGvLyMc1pv/d+M3QdL8FKC2+sgugGBckuph+j/y03giZRODF4c5IXjp
nBRAkxshW97Ay5hhtGX42eXwboyZrYYM/I7f3q9XaIR+6NnJTa1qDDazsHHYricp
1enz1GsmOCtX3RJl6NbZdFLZI88IJGfH9WXwmEYvHhFzrh6Nm1bSOrlM21U4r//O
I7BMBZv+NjtGVV2v9R38mGv8veyNbBwJ1nbQkXPaGryI4C+8oLCjuRZ0IJ8FFYcU
XCWl8vvc8kn2/Et4c+TFsyeWmlLWag0TGMRh7N1RJ0wKHw3JYCE5v2GN2cuzia6D
1Mi0kgYGUrmWzfAaPgKQ4elev9zwXge0eChVb+Y3jLE3aCCLuZ0hKAqN4WN3WEO+
DTsl6qn+sVmNlA+fn4Ai8gzfXC92AubnNX6kAWMV226fo2nYSmvnHlEq+0Cg46Yh
4svM320Qd7cXzmy1fBs96B0shbU4sr+Q+9gCZ4bjzQXXS5KUAKuVLKo9qnkRTm/H
HULCXLO4mkHqFRP81G9fGPVM7O8znmzLPBRNbkhctPjj/S+epzaMqXrNaDPjs2hX
gvrKmvmpX1mFVpU/onLd3hN+4gdyuSftQj6Ylr3bLjF6G0eR26IfsCJSsQIFZ5tK
yGa6lUNXJ/wtHXK3sJcaR+TWcPo3/LWDFJ7bgmndnCkRFVOBIObsjXhi1IK8BRux
IMcI8S/BejWSlRwMWwE7ZbIJRNEuaDCUCzyZg7xqfyQ+Q4VqmO1+PXRlKI7ROStg
q2H1EFiWkFRvpt2+M/Cjevz7crwePnwq29Wi2kRQhno85oEDstdFgPBtzDSrroA4
91pXvau5DFUaz9p1TMN1iocdYNf7oOAryQjy0lIwDy/ajXifeEe8aNgMBchj5FSe
DtsSZ/4e8K5wxM369B/BmSCoh0jnPfXpDY7GY1Z7OxmENNwSa+yPeqxCDQlboCHW
716yAS+kA6qV6+OkWaHDs5U/f8RD+4vpiGqkxR6dBzDCqlfvzBUyrBO8mhwfhO5C
RayjMvjUFzf+hDfZkrkvW4/DkYfdvZA6bZEvuvOM1jHxz3hsnTCrhUcO2ZShwmsP
9J4MtxLaLqQ81C02XYrknDwXFCvGLu0wv1N3C3v+vEEi6kz5CDbnTdnLGQ29VUwh
Yx0q+iniyaF0DI6+GPU+gQ9ZKt5G9AXBceLSuL9LV1GO/dvzch3Bbljf2momim0c
eeNbh6hppt+xIK0DnnWT7LVCOGVcbww1OOlQozURFBtwSZxQyO8+SeV4Uv5cFA+R
4COw4qtwR/OOVxZgonMQqYleZ8W/Ke7WN5iqZZNGDNvpa4xbN5tbJtG7ys9TuKe8
t0qzli8lM7Qbm+RWgVc5O/4FZ8uo3LkN7AmxQO+ypdqrXQ2qyk5XRBRI+L8UFXjo
uORQasvfAvz6li1FBW2BaDcIVnY+rTkVgBnPEtGs3IBbhrJvidrqCSomxutjPKS+
K4cT2Lwz/3wxBnJVUN91lyOQn4Cj3mYjBdRdvZDCguVCguBlRWOWIKEaoSZMylaR
At/jb2hrIUjnaxCcuyPsm6TOJeO/wkNZpLkvtPdNo7AMHlgrroY+EGemc7B2Ckf7
VmyT+730RiFy8C2oz0eB6kELjMR1zRCltEbT8pl0kTdev3EyxwvDf9U2jS/I6VO+
CW4gES5DSxks8soeW+IFv4trFbHhKHXH9qrpvkGiWpr/LmYC2v8bVqmwieXDnFz+
/nanC9x6lSZBV4nR2oXbSIqVlFZjqNgmmqQyJLmeLDEW44iP0STp+YFXiCtVoyLC
YeXppuTmohtDoQ2N0wSX81nEwg2DzHPJfPXqv2Zo5bzFZD9xfPCoaZOI5HgBDd4q
i8yeybXZY91/1ec9uuhZZ6ygLJYOMt0hvhBEtyemm78YZ5YxQJkThWBh2JDIDu4D
G1vSL+6OYwlbNjzYf7wG+qhi+aOK8abnAy0552UcuT9DUn+V3XyALg1xnYfs6RO8
C8rNOFfBp1IwFcAB062sQTfn8OCozoOJCfGF1VXOLW4RuBvkHNerO2vnLsL/Ac1z
6ihHQ2bYEY7XjzHe/mvMfHjQePMBInFZ0iH4EQK8EZm6Nc+04TwijnLNf6+V70Qy
VZGkN52f1XEZ+BjO0qV7udtfIGN2z94fnHEgpzbHe7sKsakyKY7f8y9SA5JF1uh/
99jJ/HjDjKeCZnIrQWwoEtfvUZGHaYneWzkcrxEbHt0YmkelGFSwsMmxv9JEb13h
WZEoNF8du4kuvClv8B+C1GAMfP4bgv/n9mRBmcm3t8EpkbhUgNqcfeBCXN2AG8PH
2IspvjC2ZmtjKCBMCvewSGtmynKGnkDgkf6vz3Pa1gW7xfu6nfPk9fRwMHoAsHht
wi4csqM0tW2yCfaTnTKxcLdwEi5xdOxoIurzzZcNDpMx3pxpH/h3dMrxwCB4HNIC
mQYTziR+uwyl6SRY5cnUlTW1eX7k/e+4iN/WVAGZGrT4quavF7cfhrUNSaOXIJK4
gpLRFKcf76AVhhP16suVtOgy7Z65HyQ2Q/mPVhmR+rjJy5+3QYXygydOnEkQwqbq
luPRF1O9Rz6yEBOWMgoepnSKmImSf6UuMOF0UCKsljU3PfrSZnrRvpYODNcmTjqp
CotuTMesZvnLC6rHmHKJAD5xh5cL4ZKD/oY5t2r9vXN2kKwQVkrqaS132SlKuUOO
WtxRZ1meOHw24xelJ+TX4Wh4zBPJ4Suh5AFu2M329DBb2iCUwd0joecCxTphd2RO
nEhAAm5Z3tvhXiU5RP43hSDXq6tbr6VuxF3RViI2s/qSDepGPYzhNP51w55wfHxc
msxA9FXSQISsnUl5at71Ma5dPZA1GJS67+RfKcZPGTAodsByRqi3M7POrpmvrpdb
0ACtLarSNMrM+lxaEFJNABc0xy8pFUYPIp1JqLIuVfeJbijOoNyQEmHfM4x7Wwr+
B6NAKzeaLDimsTVcSzU0yPRjuDeNRsXiUpU9wh8y16X4Dbyr5ps42MgCNkz3ZVXN
+VqxdfYrRShW+lZp108bgvX+prKix3J+rqGrLCRcxP4Mi0r2K6i3j9lwk67yFRMq
aOJmahtBVS6vsB+CNjwnC37Hz+8IhRR2m6nApgxJrf9K8O8oaHvlf8yq+PE4qrUB
EqaAfcasmQzMtOx74mMVI6LLzNhui8XEAZRhs18RB27rbV5UnPGrWyecKMOi+gY0
O/YrjcRaOXxLcLtlcJeVUJA6maoZKo3Agoefsyy0PlDQTMAeK4BoMlspZbNLlPYJ
pa3YrK9TKQxoKPkmZVam0TaDkX19xKoDQELqC2wZApZ4otkLn3rAbAq5sXO7CaM7
5uANUd7HB/92mkDIYJz2WnHpDiw05HyxfJ8/Sr6Vp9gUFPlDQSxh2G8ov1E0gZhi
PW8bIIdt9wL0UKW6FmWshIhtWcku8E3Pop5k5OhY10SOiSr87CPFqv5Uq1+jBpJ/
cdsOcQg9dUJq4EBIdlP2n2j+oMy+7pygE85zqknsYyvwtyrYWScF/QI+tXHPple7
/06ojyQ5ndlcYDNCjrggS8RjeRLhdNyygWnj/QAM7Btyual4u4VvESG9YdN0bE7/
lKF2OCa71lH3cGJm4yLzCZ2a7b4gn6Eb8Pn724iJIk+wfKKb+b+fhYg0It/uDPwo
yXqv1gSSPzHChvphFYCWvSUHVbf0ajCY33OE97vIdii+te+1bbfaKwZjGeZdr5Cw
LfO+jnlr4Vfs9rj3N0b5qc8jr6QSWBzruUhQXEQaMPLF1sOVQmj/chWY7b+Is7aI
nVpVYvuKuZVzn5Zcv4vI9T9lVz5/XZqcQKUeNV6BgfyJOU3Dw259Vw/FjHR1YtRQ
ISA5QV+q9yhqEIqrG5U4zKfksFPr4wsvTfumyspt0ZGKSWeqN2lLsWNs0ZfB7G8H
BH8/aKxqZjqvyljRH1tYPy77niGquuQQD/6DQVl3fm6UKtqLGHJz1AvGTSF/1CPB
ES75OmHLmhy60y2jE4gzOH5MBNhDN0bqzV+ulLLF/LA8NztNsoQ8JQirEzaAJeJI
gUED1FfdWIR6wPjmERzYHseuyW0zD7enVaF2Z3zG5innZ6RkLe62u62SPuDq7vFV
AyhIbB/Hj5kYc2FK/0K8u3i383a5a0roqvhtJ9BwuEEloWf4C3iTBjlbOkSuKGZQ
H1aWRDCSyF/P35VMY0e0wuopaH1I8OI0AFIWE4Oy9czmw2tpJOiMZpiFyGufveVx
eV39sLufpjDg9pM3vgSy1n7DgrUuP8yQaNrrVtp8xlRqxN5UhuwsEW7Qw3YxJtgy
mgwDQ6hVFrmypFWbw0MohK7+Dj1CTuXU51lUJkFnPseELboeRCo10a8cMgpTpExX
L8UxWeAzcVhh0rw5ar2Lc1q0iyyE7dnWFoQThkSz1QH3EnHEvd1TlFpbPCdQNpi9
SbN0YlgOWIyMmgG8X51p5c2TFiS/enDckIgAkRZJlpbjEACq4FfWtGq5ozHMuRRV
CY3hjfCaEgv3yy5BbM7GiagwOcfbqZs/+2T4WpDnIps4xvVqFI8F4GwAOBRkxdru
4PJPD7jlx+vH7tUTu7pmcS0lAL8FbVHDPhxHxK5psMo6q6oYjT54y6v9raiKPdSZ
Zn29SVoiRvcq7ndrtbdJB7evapulfNC3oTONEmE+Wy3k7vyhiAAzm00yDnI3rYYJ
A6IDhgDhJ21fgGI6YEVpQj41XCW4BkELseS64f7aQEBCe5r9r1LVmSwgyW/ffP/B
UXl74HmrSiO+xwL7Hr/9URVyaD5kg3knyJVe0aU53W7h1WApiTwmPK3GyPFDkcRu
Z2Dab9OHPGDxeMyNgREBoKaoxmjm4WFHMRBRg4o3sRBJMe7rbIdCg6PkRj4fK0Ey
VSjpNC4twUZ4sHQVuoML7D4Vq3rBZwUH4J54SO85U91Jhrdb9k3gd34ufzwo6I3/
nCWbkttCvOivegYK2chNAa7aLpP/21dv92GCL0g7J1HhFTjKLcyce5mPMuQXDAGj
myF2YDhEZQVXhAga+FMyK3C/SfB/BEihpmkNUpnabC8AxUIucjBemoMyBEz2QpvJ
Kgjlo7mo65e1/q7soVgiV2u9j2mNpwUCxWXNp7zr+roO/G2KAvXoWtcdOAdjIXub
0VDtr9YRL3QF1vzMFoTouP5vabbuo1ukWoVP2akxLodesClWFvC/u0uP4/oYrRlp
Os1ever8R5N5N5k4YzFTOZzueGOPxel911IpjEJfD4EbpeeN7si1OBz4zCtBsiRD
zSMP1b99bRnr31Rz18q9jOfxTNJEiUQDDyIf48WJ06VGF9FrdHDwEGoF+Cu7S0tz
ctEN5G0grFtnxEqP/p9SE3oboS+ryXGzd2irO5BlitrwqyhCJejKFpy7B5Trkrp+
luQ2uPkyZSFtX3EPRAClBvZ0D6hu0GSmgJSaVJ0MIj3lihrlEaQaJ2k8t6oOakQR
iNMeCy/zPgC03R7hgf5hIhbFdZHEKnplJ1Lm7HPsSyKB8lbsbel+oAChoFrmVM6/
hWL+Q0gW+2TqvoJ/jF2TJ3Y1/qHZdSLf/Fy/GJFmyar4xaDFAE/wJqgJyDiyc5jb
Pp8pi5+4GehzciuGeSaaQpcmoKPGMDQ9UHy2xkczUxelbzMvnF8i0zKd5giPFcSv
u21GVNuBzOIeWxNUckuM/fL+QmZY5Vq34G6cr4Bg9hiwYw2uKToRgMBZsdif1yUJ
dZdU/AYXwYx6I+H/qaALN7I5AVQOZKw7774uOrnR1sZtirPVKzWZWMNTQ2ZqsgtJ
ShPGEcwrnhuT1bONidlm+CSiuV3LySox9hhvfmtqMVKnjBv5jiLPao1dYs8CTd6r
tDYFtDn4C2HE2H+32YUDUl3gnaqs/y+Lh8wtz5H+fFANxcjniKNxP85Dvddm1mju
q38luY0uJ96fmfmRsmzUPg5mqfX/UzsZOYA0e31vdLktPuJfWIzOzVnE2IPzF/Jv
EspWvIrvusdbb4QU206plq7Wn2LU/QOfX1QYN2/MAkB53skTcGKUZfuKpIh48+bR
IOMQVT58hDobSK3iRBbyH7X7ND5f0AZ+pxThawKjOFgN2cA9hQFMMimTm+pMUQ3o
xC1r3dKz2+rBdfDaMpf4U6cq7dHQlCVPLuyNeMYwlgV4KQyuShjCUlGhhaFWcPd1
y5zKpPqfg0EI8+J7gan6nFHa4wnoUlApX4CICAs6vU/xtlODeuDNErXDxB+kDnbP
XRDYqXm0l3Zre1l5mMlt+szUTaPv38Hl74ezwHxiYzfBwIHvs0uch1j0wb4aFIw1
TvyU0Hk00BYr1gHO7YhkVfG4wLv9GolWkraUhcdCyJjEN3J5vcwTz7I+qZFmhnF4
t81/S9t+LGRfpJg2mXxsBnnpkjoIVoQGJLEDqxpLBSfoBXW59dHJqdJpccpxcoUs

`pragma protect end_protected
