// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RxcNfV6thp74RIBH6Sfg7qUazkENsLZF/iGqrUbCuHOvYXpSYVw0VXa0d68q
Z+Nm5/lJco5tRvev/FZxDrBYHjxqY7jPWmehsZii4vb58cLOlWnjLL2S+3Hz
uL+4XkxAnATzyIfPLvWrkV/B77oQmEs4eHt5XoNvqENeJgR9c0wjX+UBJrz1
zbhCDxNkS3I6BT+wh4WxTY1xzu90WbGbHp+JVopuLu1IkJ+nka0LdRZto0hv
IbavlyQaupgLEToPKDqAuJP6dRRf4MmBKSudA+Dt7kPxkbyp9Vcn+t00kZM/
DTbuNpsLMELcd1vL1+qOKEIYih9Dt/PFbn377fE56A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AokOB2s1T9AeQX6DdL2BxoeSnjbdPgnRwm6lVd5j8has3xefHOpz+X+yO6MP
/9Ypk4OdXFbAbAFYvjVeuxZHL9y/eVyuZ0wAEnkzPlkp/sdQ9/oTKZW7eOpj
CAB5mYvqMzHclkEp/LoiN88Q+iTt+yQkTLlrxxfMWE1QrAJq4T5hcd7skw6Q
lvblZq/qJxUYdTbzdL2pV8tQRNoCIw/IfZtSFkUCD4SxSamqvAXQwRSZqdcP
iSgL0KNvsrH64DZSE8a2UN808AYMYL4WtP3bAil06CPgfb7UPj7CzOfRxUn1
kW9VnpGBRMEwSlTtRASyoRUzHwGIcvC8r6XNluEESQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Vc46J4FB0ozVT/UhMXZYbyoDNB+J3t+A9tb6lpK5KPXGrfNRohZIWFUFzeRI
V1zM02cfdgLDEivnxtcJ8UGyujtZROLKcAEJbzFXvFN7Pz/tJ/D0In0Lkure
PFjzXeuFqhfkL81qnQWSM4H0oHl0FzBDK5IhI9PqaVgr1St3LsZ4zNZFgpXv
rcZP0aMqKgH8wuGq2Fcgn/Wxgw3rvuPh/Niqvc3iE7CnoGpm7ksXDWp3sKcQ
LY31x6g/34wbWHUaj9kj7KfbEzE0T/7CyjYgpo9kbpnwz6FWE7X1L7hlt6K3
/3Lg/cHp3+p6GouZm5p8vRSVIBCf7bv0OBqEtow0FQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d6nwEH8v44t6pCsbRXFWljWuDj9ZuJSD4Qx0okzOPlSPUhwrRLHPcbvT270g
fTxXt1mS8Kj2wdbxMeE89t1x1H2E/k4DQ/TE+JsqxyoduI8otqfQ4fh01DYM
vVVIsTsdYkE7MRHhKxTZx7+AeZSEjEogaLlwE2SNQoUVqw1PIO4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yDGkHXcRSEaH+so8H5nnV8fO6pScgIXCAizEW71Yg+9D3vl8UVHgfx5AD46b
t7pFy0KNgqRwcDo0mlyMAX/K5IL7cLe+MWttllMUS5ui5i4y91KQOqt+2pIa
2KqwGXzEGmnt4zLpQXO4NjqFoa2atmNzx9trx89lG9OXb7T8ThxypDUM8Ijt
VlgWjYFS5T54eCHmPZkEo06maB4bO37Drde6AmPYCJb5ivyNB4NT8Zi2biDo
I0BUzY1hpcqrCUoyDAQ9jHzgYYzAuQfUtnd9oB+A+PNtiijjq2knenwa22mj
/v7YsRboa7vF/hFfYg11DwwQezxoDlreHzrylSiilRnl9XNTWP+c8XY18nM4
SVpeLMgeBysi/pQs3JOrGl6dT1uFVrfi7U7H0fv87MdyxF+7nS1ldxerTdYT
unVaBAJD6ihQXycHycgnkhKNQC1OVDHPHlVGrOR5SnSdNQp4n3tX1p7ee09b
PdLoqNAeU6K9QOK8s6OkQshS9lJtT/M5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NJMQr4Z6CWkUOvBx8qS9C1S8TXJsveqtA9oaT9ozGCqxlQ7/WyhcoZ5OCXHR
93K1rAxycy6ry6rqf6yCufmM7pRWTGMSVX8+Tcbw/u/LijwNfj9Vrl9HXZUG
bWq7XXRIXP7G9GGeG82kvIdPZ+tif9rKHeW5VbAkxTO3y5NAvTk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DFLORUgi/QQzyxYOhMcdLAUlgCiU6N/FDeUe9a4TcQ/Lw0hyrzxz9pKPZYfu
cqkdqni5znbfyJIr9UmDLsAigI8Tb2uYDmM93unvCWzgK8oi+N0Mo5uQ0nyi
b3SJY3DR1dbUGMO7Qr3Sk1g4kPAt3p06LFy2XugCe8oSlkYykZs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8544)
`pragma protect data_block
gPcBhJ3FAkPnANb5kpy97rCv4hhBxMbvB3vRSCGlzLzsPwVTUtVU9mL9jl1f
C/l5GqxoNDRkoOBDk1LVeNGGE1xTjIsxRSVrD58rpb75eQ/gFjGpWjFLnfSq
g0CdD3uowaNmCeaHyXyddeBW2jE6Qw5gTqk5lRV+K4zIZUWoTok5fl3D5YJd
CJelOkCw8Q9QyZdXwgvWA+ec+Eeir+iOD32ANEA1iQb0rl+569PNCDUG+EFq
mNn4ilodzAsPGDrRdrAM4mubm2DPMJZOsMGyOCU4xcmbl4UT5winc64fNMDK
1hTDcoi1q0c2mxy/98AFHR3p4Pk71/klow4Qoi0rzVB62MJVKICAx5rEXdu6
fWl+Wlv2AwQNPsJqFJqC+/jfUwBhRDlHFp9VD6Wj6kpNvukWwvOK/2r2yzbk
axYMbu1jpcEQ2aK0MJzRvDlu0Et0ZJ5sU67/2I8GG983JcpEeVorY5lC5nq3
G/mkRxbLxFJJgCV7Pqufms5ApDCKKpmiYT4LlUO4Fti0lT81BfP7/yX2NIen
z8VmiY3o1VvoSnfYCW+PW0CjaCfXFd4bRmvZsWfq3pj0UZpfo0Lom5KZK3m1
0OwGCmMc0OlBDp+09lemiUc/kKWA16QeGSPTwA+JTKfBrLC7WWgieDwfzdh4
2ITWJeff/ULPctMzboUYuN/GW88cqebtXVnOrCyYWAHSQf+RxlxqkQyZLyZj
xq5RZ5SokMRl+Cz0RuTcoeeFzKuB8G27TwtnVIsOa3gs5LcjmZd3gYKKCI14
k/EySTGrHhlRUhqeSzHyMUhf4g0G17+hR0hZPIM8/IpsN0ICZgfF5BoXdxQG
hj7yka2qSS19aYDgYJQxP1+mtkA+RmWolxWIia9xBzKPewv2nXIMoGAYiUCx
eA7m1oLmunMYXPnFHvwZESyGBetUgFb4IW7vtZaEdTtiapyecTh7qFJ22z5P
El/4/k+sLnfEvyMvS+BchyLgQRS45sQYGJlB0rlUVhM1vdSRn7KgNFAu8V3z
VHbPaof01qPolJViSVDFjdvfZSoF3XaZwvLlI9gWeBa3RDiaPW1cen00MFs4
fCnOee9mYHSKe7ACDGNYxFNisU6vf+vJTcpY4dNnXgw0h+ZiKAB4f3O6BHEs
hUv297bW1tqazBV3iMEQO4bxdrToBWQB1O49oRBaA+R5I838TNe0m7UMjl8z
5443BXERajtdiW3V5skNrItR0OaAzlbycxh/BZ4zn9Q4r6pNynaIidFTTy/M
/f8fNEQGgYALgpSyuO/NDWXQjY6P11/wS9AVyxhhOVwWimo+PdjmWo4TXtri
sCm+Ll84PQaxMcSHRDk9UJ7z4m7/0ZJ+HYMACPHinOxYBhL2J7Qi01tXHXNl
RKWmPtipTtnl6p5oJj0t8rAIj+8D5ydqBqL9MD/BwAbjTH1U7D8fBp3vdZ8u
Q4N/qyWUF8Nunz4XpIObKNlsUDRFwnScvFH71bOOLWTTQKTzMhJeWQa6hrqL
QFe1TQziVfDC4o9/yumz43ekIQGSsjzMKmgREnbB3w8eRsbzrMiyQsD1yBpF
NPXA6VZ7b5kTH9KnkhO2/VzFcGMtjaXKqOuxp4mKKHHA+0AYiCEUEaFA+Lhi
0rQwn73s35Jd78xvcbJ+sx3CXVM9SSbCbVMSdx6oO/10Y2mDcWXeq9PZWfFU
93tSDxmqUXbrFbL7OflPI4PH+16hDaY3TKusJq/Fxkp6AVoRtA7xDTvaGtC/
MT2IODwKHiAjuvbe0W0rAjo7AgU/yzEFeW37hLDtlJLGEhihyUtPIpqmVkR4
yqox5GN/ySRghQ6jrY9VGWPpesYztXa3C6c2K/PXgml1fU847M0F0xJ8Gcbi
oOf3f/erV1ZltPjE+tvbv+hmN2hmF1oEvypLWrke1jDvtg7EHBKDB+y+db1X
jlipaJnk7JfTeBFJKdb0fvOQ3PKWJWaozhXsaNVPjb2+4N7/ri8FAerYstwP
mQhr1pqC2eW+KG7VlP8M5kCksTyyX1Lh8EJFVsgqJE1IoUSiAhAeeu4iqLjL
zc0JJkqUd+9Q3lzVvdI3XVuWMEinmFh58jCxozQlHNETWeudTUUi2Pxz1Nvf
jldCIo1Naa7lczwbtPuRY4lUe+IQPhjTw7KY8PJLj/Qhc0A9jDilaJxyM/a0
zui+yZxwoc40tOuFIectgVXrDGo9KKEZE8W4pXhsKMYoXc2yKNW7pkwyc+0M
dsHe5gWPcGckynDg2bPTiMG930qu2mLMMhKazsW7yXLMyXgHKy5LGJ1YrA6q
cSi5PpxWoGvmbbMlqaHvGJXTpE813tkRY2SuFbmjJ2uo2Dk6/GYazLVE8k0c
Meu882MhI/ZJI302OhKi1xcP24axmjrpdii3OxST5GGfjxhTQtJ4Y092EVk6
gHxLigEFZ3dKHD/yhCHfPTuEjbiqp9zzYV15r22nllMFoNWrWsnah9hK8lB7
I9XA6O7xoUL4ZAv5l/0Qf2lXi8Mej4ujORbxOSJ8lf0kL2FfQ67kpRVzG7SE
+DrfNliIvFj/X8OsbYgUnAWdGHsWesm3nv7caSYKnegkRTfvYSqfO709u/cM
EQIc6ZytkaQOGzD2nO2uFQA7ZEuGC8rDQflxo/DUDoZCsyTzmeuUVLXPsNTc
oAsx1oGkrtA35FP9lYOPKXyGZySg336bd63JPkLI+TcvcPoIIvzMXk0rSL4g
dmSUSxieKk7JVnoFlH9zE+WPvBgGrkqoixBwXpTNiDw9wZCJk+ytbk0UMsSt
Wp0ZvFzBZFBfwEiYeiXNpaa2PVCphLaDCeE3HbNxWeGGOfbeLFd+CWz+lUyo
kMSrEf+LDBRfBfrxirK5HQXPILJ0qYfFtwbBzEh6WBM2DjaB9VmZJcmlLBW8
oV+533oQgHorABkj0CUvRzeEu0CVrtc3OnFumlwx1wmr17Rhmrqb5KSQCK1z
4cYdlTENYGjMr6brrSfH/ThgeCBANjHqEu+kiBmQ+atox+XgTZX+9u+JmLLe
LdnEe1ZnrDOLmdsMEvqv5i1HLWr4srV3GgGq6TW75kaXGQR9sZ5/cj+HQOut
TCF9rbe/OFi7x9OznY+Yjlb5QgRveJl5Kz/R0mgSqlhptEudCXsEjjjWzADH
oDtC2AIj+7sGrc4IUhqfqYksIILbLbB5imp0ilMsjlM1EYCZilrZDMWcyTXE
yLzHgml2Nbn6YfQ32uAQEQlczl9Is8Lv6SWZC/QSEWad5UiDydsPMP2YOqet
HjW2PtlEt9kOxz4GDJC+GppX7dLgLtoDVDVThvYAygX3rbg2x1ZXnLBfwcgu
e7ag4psYkGzRsYpFZD0n1ZJtwXxXethhbzvRKvhOU7eKYpkVuPdJyxO4LX7z
ReFWXcEoX6aqF80ZnTQljsql+3aBweIyjamY1EyRFRgcFgEJ8a/N9Wi9RBXV
rv2wMF7ymT9OrbmtHRjaO/3jaIpG4O8vV8/5P2yX+y9Z/hDkipiOksfMd00P
VANzef+5pYy7PxX59w78r4mdC0VqRF1Ntpmo1pe/DMSyVDyKnaq8eKutvCO7
Fmg6dtndVWufAGsjHQkx5jMILJD/kYSbPRKuPELHwgkSGMbaO1Z/AmWybCDh
ri01Pv21V/HkEUmB7Ini5LTdy9ETdrDiT9N9hIFyrUhWlRMQgNpxllqsISAR
zxSTlVsDDlwKhWJ8jgMzaZN8QsSTJwwhfKAdIMwhkq6d2/LNAVpSiVKczqvL
NT6jPQMo6qwwfj0/QI3WeMcLuP2R1vAylXsjNZMAt1o+KcN35lD0h2zJEJSA
X66mQOiW2cx+cNFr8n1RmxQiPd/31J4S2RYlVXdAjxG/q6lELdg2ehnJfE7l
8R1zW0ih87p8a/LeZ6YDPvYsRcrLMlQYsQY59iYzHg0OIxXad5mPtlera+jC
grzwTy0PAp4w70vNqTcWWlEByrlrNNG2IuI2r6VlOMQtbRCsUadxKXI3cFIu
jGKcumJ1QnqJl1n7GRGc7Gjq/b3d1Ms38+++K55tZncodO1SkG4ls+V26jG8
Yko7fYhbB8ELWCGWAGXrDU4EwisQK8xudcryLyj9gOm71JaFDZDKGpFNVB7W
r08li/ioRX0qWru8oDOZ5g4OL4rLqJWXRvQZoKQgY5daRczRvDtfRbobtUIg
Ihv9kvkI2K5fEaPPzPWPaDa4P+JCoJNvnX8wcsLKJMJAxz/eXPseNuucl7UR
rM2gMnl/0MJuCHIpHOOdyuy71mumiBsxIeBql31QMoV3d/RP8tbnKUrFP712
Wl5FBU2EiRVNvOFq8FNn9GSxhPQhnKQe5ahn12fFPFmuwmWsMClQA06Kw5GY
tnRgMMmkmQih/6XyKq5MRpyNFKDNYBlFq9Bi2ss1AVnAmS1zB32s4qnMUKSV
VPkMc91OBJJRtgg297dEKyNFaqGS3xf0J3ko61rX/wAaoC8moLqi/gJ0Cc78
KKc93BTQaHr1nUIXcpXBIVDLzvaAl14RAgk6QalPiMKTGxmw0CRT+lOnVsls
9+qJWRsP3HfxI2l0zFEx/GQ6/nkfrOdjtrrjvzXGJpVofyihGMrPr69/J27W
/xqzrLq90zV4qN+TtFH4Jq/F+JV7Qr0Rd60A48zReR+ZDR1FeA9/jxF3xmHq
EHuuLFNe450HcExX+XqFBQH+pYVb3LUxH56/7oRazZ+yiPp0cYjrj2ICE1ea
IYE9XQP0yp8FgAliFBxcJvKCqbFR1SXHUSvcQU2d0PT+zEBiYE2EMnXXBODN
q14qmOngLvwr0xNWs6e3QZdz3H57KuSGZpXGlfbN9ohJ8aYyOnGQ9RYy7t4H
LyFl3aha6oRPFzKFzy8Yg8ycJ8WCAsWqp/JJr0GTwNBVzsUVOFqyHNvRogdH
jgWqSg6QwOmmM04fBvZ74bl/OOo/ofzvM45sr0wrN9x3ae7VsvVODLiiS3bA
ZrSdxhWGSfggNdzfuZdUdqLoLRwyaKvCNwzFoqYte3NPIJULRk6q8zc/GN/i
uoZsPie1xet0/BEyzu/nmc0Eohpe9bP9jMTJ9+YC1soyHE3SK2Oz0Ur6Dy/f
Lo6GaOpuBZ9DOqsi8+6B66DM0EzS5SdBSwTZlnfY8f0tTzTgGHBI1emLA4l0
Hp1UY80+pqsC1A4zNlbwK0Rvc96zY6U7bZBLCDJHYm+oARbO8n45h+b7ggMj
txTsAA2AygL8hZwYqpr8cR13fFhcQF5VmkOzvdQg+NhF4ywbFtju5CMbojIv
rHbJMFfi9kUplnIyLNZlf984U6ajJsu47csyuQ1NyP152/p1HSHPIiffd/NH
CBAHzIZV2j+ni2NKDUXMXqefyJUa90s8z/cVjnf+NSHAR5REkW9EYqQ0Axzi
SBBy7FUuyTQFT0UYIu7jqBnzApM4G3oPC1QjAT2V60udpPhhltHApTAf3Q+7
ylhhVZSl1e9clt3fGZTW95yvhZobRUzEz/osgoso9jTpK/2Fh8ajFwz4qKHr
/xltsf48Yk+4Te+Ty2x7haQKYd7yDKQzTSxCXU9FwwA23AAaAHd9Wdx2TEBh
tXiGh0xblx9A7T72Ooeg8hlUlTaDjrr/+lDfNDpNqKJMgvY5y9jOno1bZdxe
UK9yY03RdyRiwwZvGMVqxc/OSanSZAywth4dq7WkSrnuTL7AHDoE/GGjJ1tx
x27x28ecyo5tBkT5g2Sib6ZJmga0/zr90jq0LCgXcoNWt7pNvLksQyE6fQwS
uW1wiLryTox+6dDCIzmyP6+yqA8JPEcWezlsrOdj29Pjp9uSmWFukAlEtpBq
4MEQNthDSfx8M/nIl8W49ukop+Z+pyzd2mfUgcyOaVzmhUF90rso2vrKjTej
EX2wSAStztBWOlokEDSJG5phF1mLup/Owrf5lh0lvLsOtR85J3mpjKSfSZa6
TdOWRVo81ZOT3YTckbDgK3Pfs6NsqyGyNTUl1R8q/j4Xo0iC7YhPQic6dQwX
142hn1sukLA6eI2gf7zCTZy0UiwET2SKH/QFjZTGzhliK8eX4XEJewGOTWE+
FwbGptnVGKSR0QOLDAHZkgTflYsR2Xq5VmJvMw+aNSBpcngs6SuciR3Gxx53
Q05QCFdjsd0/o2IEuv/rWKXN5IOu1V2TbCs08QNbwkp7mR6TEnfpU6KoROn+
hQeyKwfyemzjNu2YKqtKTEXk+cq/B54ywsuPq81qIrHofCSyrM7tsCDqcodv
oC0LzoZOEWOwDGrY5DQEuaLCrmWMrgmtJjT8zIgd5VOPSAVVd9+4X2Y97AIk
q3H6Ziuz2L07884xmuCUOilDcQYDQ1Cu1VbweRcY4hjv8R7P0Gn5+M8NA2/3
Uu11KzXbZTQV4Z2ZGp3rGtKalUhy0fzEU6WYQFQaAdDxlLFteuuKFOE8iOH1
R4gUPYUoWIHINVp5sUFNtrQQMH0UE8Rbi2Bls88OJp0ThBFWXRjZIjX/psPz
mlU1Lz53KwVx1yaO/TPE0KbgbIAn5c4V26K4yU89PeybioVHH29JGCg3Oo7k
7Zx6bEyKqz0+lfw7GZPHIXUXswriIe9LZnGba/KsX+JUugCLc+RuWcvsEeLP
FSDt6ofNK85OuDyrU4MoBFXxuCE726nsE0Z/hBNv6OG30MqYBUYdykcJyO7X
/p/fN1bE9pks1yJmN/VKNdLUPdEgSerg6ZLDPR0UnL8egqIiL3i5Ah7/v7kg
ss6WWFJVQ+rnpfi8Jgi5l7+MhuU+wwFVwdMHXaMM6+wwFC9sSlmO2UYrepn+
7NVRRwfH4BQWhzYMLQjfVvG3l7sCnnpKWL9EahUUY8Iggff6f+jgIxX3dGJI
VlmifJuLodLQG8DN5SvHSQoeO1muzR/beTZXHeOx8jylIcus3CnC39GF9xt7
JO+HWZMb1JiF4UQr2vz1psaXrMXCtdMabLiOeGmZHRnjlOlWoVOhUT7mVldn
9TIEDAdEBQ+TniSMG5kCT5A9e+0kPYjJzYrQM3UYVgumECs8ReHVuyJlhVGM
boSHT28vBooqOh/2sD/8qAkunKb4Nu+6gC1VRZTR/mgcGFPpSimP753o/mhS
8e5XYMh4gYb8FOV+Hq829gQFrupGCfuczU22Wk+Dk8Fhy8CSaL7FB/TXW2EI
tOoyT5pSS/O3TrZL4QbT+n9ggEdtM2ojvML9wdE984CgYo5H0uTNs0xiWVfj
i5bzUTd8obktofIK/G3wGOND9vbzf8OG119rGqPNJ00ZABAJNBHwpGYkefA8
AXp+7hTCmSgYGbV2L7qBN3h0TcO9ygFmLJBlB7OSRcZOcxgQYE7Lp8gifew3
gmW3BJrLtP8bBFFH5NVl12/qs7E6JN+A6T9ScEbciRw/MNITGiz86Pbq7Rwc
bcvu2g3WMmgRFWHeHtgPRchY96JJ5kM1qvmw94HFrpmX6PcFXa7/ltTYGfa+
VXeruGxRbLTlHkVdV4s4C4RQv93Fu4YvfEUfD0SBuHU53VXct9TrX5CzJHYR
NFe/0U1Qp4MwiSkHsBFjXm4tqBsdcUwWYLOzNYf8kTGv1X1ScZYSAzMnidHW
1POL8EmjwHCsRhG0ePks1ANylEXw84oKvVehwwWdCvT440VQB9u+Xr7+v14i
SvSbrOZircaXS9JGqjd3dDdPy00SLwZSSjTMMnaWDMB0y5gaPi2+kXhkcFJy
2QlTRCk8B54tFEgDzLWIre8JLVa8kb3Zeu6wP5fPLroFVgYGbgYruh+EgPGn
u7X9ugA7TdAChQTeyEoPXWpJWuFFe02F0DAMO3Z7voeYVH5pA9tM71UDCLVk
egEQY8PR2iRIYsgDvRIjgIWY9zecRAQ6kavvDnywycoxGGL9DLPmvVRnaRa1
LJsUg3FHpkJQGw8OUA0XIey5DupRNtjeyz8wgqGwVTOuRtY11bZ1/TFgvp2k
l9qvk2Ej0u8Ath0KPtM3lZVWAIrNK/pHn361YknwfqH2UVLyHcWT443yn8vW
LjW4itS3Hih7TOzx1X3ah4RazyUsreojJhvpWCDWaVEDgEA0wYhRqr26dfuJ
Cr92vUX6KV1/nJxJfrX+CikGQgER/Qbvm+YWY7zcFu3xo5jy/J3/K1HhByYp
n8wG0Sm7rzdwYUCGk5jq5Xa+EDz/43MDOORQsznSF2VDxgkzsZEoH76Ob592
CNSAQNDepAJwGXHGxkvz4UFNwoi34Ek9VhSXPSUVDVAK9rCt6JwSMU/GVWM3
xugCjXCy7rI1s95r4QFA5l3Nx49DtaCBQBaNqdnRo1ls3zvbE5terIQVqd7d
u8IvVAjO7Yge55wMdKoWrqv5b/ONJUrgu7YqD1pj6cmUvOfkZV1hbVgQrdY8
IhkOn2NhvtdRkUvi+8bR+6bU4EUkYJtFsKTroLrcBPegMKCNBTrf1gtuGVh7
lILhU2v09xxyncCZXLdCY2XMvKN6fR7gpsQ9vfCptGKmXyYAlhHCwGoKCEoO
iOtlLicqumqqFkHRJr8IsKb8zvM1Rq7MU/+xvTR8Cgmi7WXKOomiKRGehowm
T5mKhl7pcfYjiN1NrJMQmtbufGGbg2oJWoxTHWiYj1HodVcj1WKVwrxko48D
akqaIkiw2GFAO8Gqq7uKVJ78kx1FATFoW0OVrhixeldivHUMnDSNk4JVTQyq
yhfKEeeAPEgAZi+5BytSlgdTLL2p1ay8icZNaw7KYj0d7vFEZF7f+VsX4dyV
S60NP7QL+UdUNQmqLidAB5rP1MgRC51Mj8+SAKn4ooEqFvJ99FUZvgdq3YEt
yavACtGztTNOJmw1+wFrkNk08w/YoNOgpMi23oaExHjtKW9rWZMyFk4MgY/E
2InWniqtULCFDhf6ShWIiBuqweMt3q9p/U48mVxr/A9tpFLvSkzB9DD52cyh
pA9HotwkS094XUrvJkeWo8PwGyioX32qhxkjHvK2tn6P466f0XHxqmymXNmz
+Op0VH6ipYTWUzutX1beJwU3F6Ycn+5qk4l/MXLdeicTEkV87nvEOTZfdKDt
g5MFd191n4qCwoX8RGkKdyk1UD3q112T2DwH/SKtb7e4+b884qSmqPoxWh72
jq4Kdn7rlqHjZzn7HX6MYpbBumkHpeYf2m6+01GIkmeOR811fr5fiRDEmQel
XXMvaaehbYdZmZh+LnhsSDzAGbe0fD+PPwB3iJGyKU9wWmudseWpJaHbxw5F
EKmofeuwU1BJGOWlfYxOgNedE6df/Hz/O5zZ7BiCyZ6M/BmapYOdeQrYcfoY
mhtWJbwAJ1IqHaSqStReV0fsY4QyYV22Ehg/O43dVeJ9I74b2Yb67wC16tay
KDhdvacBXfFAthsnBR32diH3ilNg27Ivu3KasNE7dFgByW+e3TAhiHbSbzDq
RkAVcYAJjbB3Lj7OriEqarFIbfjhqB7Dv8WYQMZt5ESy0aKB14P45mZojKUe
gE4YCoXW8hQS9B8mdgkiUB0DVLZMSRwIu/aWYsz+435mCRVUWVY/pd/iEnXU
Dt2jqzou6iRXWRGryeFHZeNnvoLA1t6jHmZMMSfPb+Zx+uvYq1kmX50jZLy1
TUpaKyKDMg5ywndya+KsQlhNk2zzOFex+ayxdPU++TUqlymVDyNO+TfG2i/j
jaTloTZmBvAedD9dtTmTaUW6k8R+bmNDr1DqDwhngjH256FOiFgVtSSLZYkn
MEKIaa/q6YXVcCq1VbeLeXHuT20/kuf+Fq0ErNeGxQkuEUZf6vmrHDVkwxUp
fJlB5+80hobqrOouABf+VWW31HuEKDJmL+OY46MwUjXQz2ddhvAHx+krfWAf
su4ZGOF0V8gWIh3eT1otlHPRE2qKVabyA3IrtB5R+U1bo77qmoluPDowU3DE
bTuWOnqkRX6zuvqqkjIFG94klmLeF9xs+vIgm8HTkhtgLymQagoK7be87bhZ
wWo5788GmGLhBxE3rsCW92nQ+nu2e0Sfzhq2yK5TSsAPfRZks2Z3FT50J4Ic
s39DmMiYOrhSXnSgtVTjyXBhmV/0qZb5OpO5KzU4V+soI4kF7s/vFeSVLrCo
EVYl2RIKElSl9QWLtB7Luo2EyT6521bjuPjqkYJ81UpWPkUjrrtQS4LHhYD5
dxQ43JrzXLstkH45A8G5lykjhhKYNUFoWpKJvvpnWvpsnjuU/EN3LkxfiQzx
LYctxowaO79/mJ2byxafaee9XjcNm3LMJT+fLrsk5Uoc2z6mVBLlCPeuiI3p
6XGd4NNzovW5nX0N1ZxCHnTgJCCWH7jdJbW4SkNJlGLFh0R+Cvec0miwwEtn
pKT5kYgqQgzmBdahxAb8Edo9Er3ZXYvPRtpX5ODysJBEJgsINa4j29akIop7
UneWpwIOuNtqu50Cws7YDhNrVbZOKIPr56pHxAEktML+ly2q/rjWmc8iPKIA
QZGyuIjC2h57+gHx8TzwBjOgG8wAUn70R39ti9WiI4DhWXKh1H5WcVug3Tu+
ypHFe3hKQRqroxJFquv42+C8ranI5TuALE4N/aAja8yBJi0Sa0SHAcsuZR9J
wYIzIODbzUomTju3P94mbm2DUX6iurMSO0QruRITG1V/0ePi2+f3E9CgSPXb
Dph03Mhy2/OUFxYF0jIknEJ34qINVD4+RuaiemYmMgUsHtYZWdNT5wGdF9wU
y08SzxX1kWGdll+iMnxoitIppBG9XuZzfryPL10yfI4XEuXQJIEVc3EKovJE
+WaLo4dOeQx58S2Q8d26ZOZmljLRLHBbpUJlCC84pGXv3+tkP8CIG0Japqek
tPvy90NwDns9SU/f5bTH61PyIuFWIfZJJyF7FB+S+vXoJd0/oKEJbRT109nI
E7CdhUqEFKTQajoy7LzVtBdOua9bwZBqyhuqhTwq+j3TyaXbTORcKwglmyF0
59vNftMM+g+WBIKzMOO/03LQlVK0PKlYox4/d+svZEiMgJBxqAxZlMrAuTsz
eGWOymwD3QdQ4nxhIEhz90xm0hcyyFjxHy7ZR5wreqk1EskPQrPVJ/ItdNss
NWa4Hv0TZGr9Elo2vM9cej9Eoo2LiDzZe8GPKj9vW/SkXf5x4fqdGGC5KKKe
wvRhfPLCxoLcbIAuQLrAq9uHwVCs8gqH6sp1npAulp3UbGKF/cvaqZAR0Upd
GD2tnJ6yZb2tX47hR3bjD6f+jNQSCak9c/iOh0UleVxKO1wxKUCN/hWKTdyI
F48t5V+4w3+rHSaj5Z/bnett3ydsR127nr0VFmZxlJ6cfgx9+PRHONHUX6J2
4aaAicty4QLCK4tGaTTaZW9/t/kJhE7V4h9QPPJdwBEmqtx79RVFmNaD0YWS
Px/BrAK0DN9MjJ4mmJsdspVzUnmSxJIlt034SHpXvdRrq02LdSDgmKrsBVxA
Nx+T6wiVrFXT5K9GpJKNUashvJk/eU/+56c/VDJViD09FdKALVgJqEI5mQKi
WaH2CSgk4sIiUDb4RgkRr/wSWrT91QUyk+wYdEY2qXNI4Qp05XpD

`pragma protect end_protected
