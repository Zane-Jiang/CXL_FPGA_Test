`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
ZOpvGaKJTdFOSWPn8LZT7YRqXh7uV5VYeq8lpMLOzfJ//F+EOgmy+FMlO57xVYY1
iNhjuR+tV+fURaDyiwnaReWMOho2MmzfHWJ9VdRwfqXbUx8KQsjGJGVU3VdHMYlU
s6u2sLv52NBi+pVUOkWJ9jTvVOkvrya+pl49FT1Dj74=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 32368), data_block
8QAe1KrV+jSwOiC9COxs7+TNXzbDR67U5GJzzeeCWblS4JLrD+LFpyi+iyAjYOFm
pcBUq2dh07MKNeYHbr++IfvRn+B/ikaHktC/iIre4m7J052+IUAEAglVxCxrrqhM
BhetsYpatauhxXVTDtuqBbJ7p8Q3GBEwnapHJHCG8INfeHG3yPuW/BejUt6N86sA
TBa9MA5LkOyh/STb5Ua1NIj0Pfxtek2PDMyEJYGmgZDqJCxG3qCVAyWmfQTYLaoX
whkW/PS6+zaswmuV9ns6pBmhsy34lkjje+/7BHUekqHGnIT14g+Jw0u7VifnDQGj
af6y0fMJm9gRA3PjEMmV5ZUVljQGS5tPe/H5vIMwjyM/NdISS8DSNi+ejLibNgyg
oTK0uKk8eGca17hSZeDEDhZcxMZ2zCSzlIwK+DWhP51CBYFzCrbOsFDgST/oUde3
qTFIK/eZR1HAyXEvnIpOHadSPpAsRwTdUEoD2Xp/63RwxeNycssIrXF8XyfJvGeN
grwV9mCOf2eGK1U4ZbXARsKA6oOSFSjdSGJdoLiRxSrAF5B6SFtLtFZF9RbmjNfv
Uw/c7YStw5OjBbULunp1XazXo6gwQaftK6qfmRT86GzfyLgQ6L3K2Pf8yRqk+2mm
CKtR22hjwhQ/nhGp2F+pLmX9jpeSENaNbt9PzEmQFEeBt4GFhW16/1viJZozyrTY
W3IjtGjqujFuHbuU9iWzyt9AhmZC0vcYBo3+LlvPgkJGM/RCAYvx0iwC2EKWVMzE
2yiuoNh2nVJoWleMK4Z0aHUSI6KHkWPJNVV5lNGxlrSOa7UuwtPyFAwnRXkN3M6c
CdnZv2gomyZqgJmcYQX7+kiSnov35YGqHxC1Xa5oZpzYVlsthzRejFr/JQ6sr669
LwLX/0xjJw6xC4GkkerX4kmNghNk+HU3YkAYqElywjON9jMZYxqG2D30QIS2atKS
u2bhOkosUiHHNV2i6LQD40hj9/dBV2ixyEX0BrI92+/8OG7T+u7RodBuOXUP8nwJ
MNpsEER0Qm6l1aLSi8WUZ3dkIphHzxFb2iOyseoSfZZsfVjrqyDjCeubvVhi/xyG
SbqjYX7lxy1z2XWuiWUrN+C8ab9BKU5C2DTIMiHMYiwkBd/XwMWHNwa629KzS7CT
aD1u9qwtUx5dsHan7HkfNGzP8+t0AeUH9B+Qzbt0UUA+CyhymW1iVcf8FkUmLFTZ
CQoa+MJ4q6W1l1nPwADb1S7xGkUBT21hmWTQGkohpnnpk7fv3u41FsW8oV9U3T8D
3Rf/1twHfnBzopCziZMb6X5P89SWjT9YEqDnbSNeDgffAXhtYTcvp6ryerF1k+6/
wY35FfoGSSLYFE+DXHjOXKo5MNf6kKispqX2r11n68nouH/rCFoPwggKDVrM5D3+
epB882oMvnViifldWhf/0nhelP9eTE6RuijKC87HxSNtx/DqMb9yk4qGOHobp5VQ
CzW9yvxRXdKkzmeh7RYugaQ1xyBy7NDFoEKpvT+VI/ZAXcSSuqO4Aeq/19ItXIv/
SNbi/pzO0MQ1gMN5eLujJafru5P8rQ8ClIh2ZQTqkidivkP2oXGymW0DEKtW9pr0
KQDLNrPrEDydD7H1oVcIFqmhKLNjHXMApRK3yrBTpGa6vy/O48rnWi2pmoaiy4Xk
WuZKPHtJkVZGq5Y66NG0gWu6qcmVyW13FW9ufNkfeUz+SYh3cprSqY740NqiIm57
sLOU/vHgrQbLj/oNyw61FAzbhog24ZVAOCGKzPITtQWu6AWAx6lt2iWfQSJD5xwu
FC+xc++twIcsGwGAG7NIFemaTLbP9azqssJnGs7qz2/vXOIeI8jVOGnnlSL0nJmx
UqTn48+XvlrzC9sujZ4Kch90lWSBL6XpcgJ+4jUzYKNAvGu44k01ka5evXuVpG0+
S1esAdACBlWYtJUaeM5lIxkrIs8+7gjP4P/1KUVz/gMOOH/LsCY369svLdP+0TaQ
4+eSiyWqR0blOWB76DoVsawNVDgB2W4JPcTVhYTztcEckXlmKItIgeQOgZ+W0xEp
muGTRqqlLfgugqC7+Tjm3VceKeZRe+UCNOszFmrmMDJvkN08CsyjhwV4JHoqbsZT
nXIqvyl5W9BZZNItSHoSX26tdJcCCX4VFvaCv3f8ejkN07m479A6yjnPkn052Zmz
z1nVShZKHzKuq2TeL4GrI/4PPa68UBmGHbUtXPpKQY5dJ+1BmqGmUViSj1btyrY7
K6mp5AcPTVbU1sxsTjIxFGv2nbnNkLdsZnOxy7f9FG1br6vzfoT4Ouh8JJ5AJHPJ
s+ZejRBZrPIy5bski1wlvk7aY75Ssvt1xFW8BGsrk7GDS1QqsqNGLdkoBZ4Tw7DY
kMLJfP+r/tIG1k7p60Pbi5GSEebcyngwyw42CxTyxMrs4eNN92rGcHtXMj9FIgWs
KZVNuSCUynizM12XFCFUmgFMdhdqn0zUQSX059/j5nIGfiHggVJFDXYhYhoc2CrI
cYiixD1dEAgz8PaDK8gRNRO9RpErPxkQ1XApmX22nzifnU4ahzopSY8hNcXIUlJf
R/3qWqDiiuVQMs//AohiKR/CwQmIOohmluY1To8eUu/7PV+rdZGuZRqPLi8YkCFZ
k6zK4YOuM8jW/QTPf1i12Ab03XFF2Q/oav/Q94U37H0sOjkrlCLYml0AnlIs5Ge7
7VyrW9wzNZJI6uCLM6ZTbHK1BsJxDq5BnafJgVLugPwij5ldvFhTalNa1bmkyK1S
lLDRX4ALCS0JXYgjwS+bU2oO0yAkmhyg0IY3EMvjvxYDbBWtfj2TM56xbEvflHyI
5hagU99hlAi7tO+K+IR4p6D7CD35+O1s+Pz5eWqW9xChK7hXSDJuWUVsnuPzwfUb
5AUtkzIqqeJAs+eNS5pVP0U1l6h6tCDcU1YSqxXn4LIYqx1UnorUlMw1nn1urdIX
EEzZ0hW1WGLdSLm53rmpFn0ayRd0V5GoO94sOat9Ho9OcdJvGKPVQaJ9FNmpva9k
GvAvKgm2m3sz9HDYamao2/gpmveSuAgdQB8oeOdoOFXACiZMnK/KYjKz8UGOkDhW
aQS18CIuThTBNSDhIrIv/renxaIx54DiX9gni/dmNmUNzG9dHrqAe5ZVslNZ8OFB
z87AmlRQyG/5FQ3p8L26ASCVplfMr3WH2Dpudwfa7NfiCOuqtEGRzhzszPLU1MSc
67TpW5LRui0WTjgrEegomeuW8a888JeD/VY5QSQpaAgPQQux6J5EBMpvV7qGSZ5t
kmyvTjrwRqgtTZpHpjntM7Qso3Ai4aPLT/Y+Nu7ztBW71gZwKl9Pw+ciupVoY8m1
q+f7Mu3J5lCBIHdaANWsbBFXyOKgIgQmwaVi/gFPFFXB9+zVqol6OINCqU7fWQY6
+FHyjveHHRAA3iNrKAPQpLnNL9FsGen8JLkWC2z+MCC16LMaCyUR5gLMxtWK56UW
5kR2GYnX4o8D+VJ9rDKC8Ok0UIWVWAWnvbWZ5HAlg3qIUNh8YSVDdMcgBP6dVpBE
dAPqhoGeOi3o4fUoik4s4gth6yMl876bCZv5cPG8QdRKY9bGT0njWkjQNPvFj9sq
YHcc9UUtoygUpVgvmC4lT6W3R/xL/x2xcvnxAFeuwGaDE00K5ZmxamHSfYkpr7Oz
lKfvlWCKCyWsZ4mQGmKHmFZmO8L/5Mzo+/tQdIx5AEiTah3ZsSSt2WOZ+NCgffhC
Cp9pfi5gg4xvSuSrA7Ho8FxWxKplMo5Y73utwXDyfA4d5NZQboaNqVlr5us2X8gD
Ze08ZTrcDKMWVmGa1FA1PAuHL0Rs76aTXznM3KKH6qRB8J6SSZVwB7AsaywlC+RN
Wh9FglvVO5XehNLzSDYY6QhxrlKUbXjmCMAjnju1oE7M/Kb6Y6iF2e9gM96mfcYD
tMuA1bpBs1H87R8f3zkdkiO4IwgE2BjpiVW7FxHnD+slX2V6QiB+hluEgsuC9xCD
p3oilGusosBrZT9D0W2Chd4qYEZbqElS2MB1BNevRSiW4y+Xfy6z2cQw8fX9JErg
kgXlFBt2Bj/aCSzYGYx/nXw95E+pFE6udGu70E0s2aAjCBPjxKMaH5aCNGUwcdqc
GoK0GlO1urpxp+1nIfp3q8YV2UrJZD1QUra0QLiDOJjRa5CpdZgAX7z9WRFfQi6U
jKmKNXqit/08D3+JtyNRRrvdKlIWJZQHD307zg88lkfYes9CykqNee33/JD17aFh
xWfxW2V6+9X9xZjTqCZQ/WhHx7nT0oHipUqa+QnoEAlAvHpcLfhLPLznNbXX590Q
xBniW/hIqJd9cThv1cYyb5OmACY8dRRz6rZ0VXVJkv1hyZ1+Sy+zAZDEMogvN8zm
70iJWqfmXFHtRJ2vPxbrU8hzyRjL/GR/TJmhfDoKfrxQQKpnWXm58KxUFzGOiGFA
+LRXFouv4X02VG9/2Owgdffsj0MiEIBQnYpwyiY2kekzG8kFX+dC/XNQNXPEcncV
ZwoAJYN/9hrwTwWeQJElGBpE/q3hlbGOjzkAEcaj87LeepKwfKB20xT/q0h7afvu
oSjpUfsSfmntxS51GitQRBYMkCUf2yaLu6Hp1qZWsHD0EQIN7uYqsBXFkAs1CWCS
pfqCPwBPKuoTcPlQoK95waVB1aD203TVNu2vsYwxnm6Y/kuQK8AlGKAoVvGDTsLP
dqETGWjDMx5FrNZitUCr3IOoNESEuZjmHLNnq/bFf1+ZsJF2/qLxF1hijcx44ndO
Zv/w5Yzss0/+5rklO9ZKSERQavPTrdxHqv5lM67ipfpJo63KghbW/HnDf+8TZFjX
TF1emkEtYkzGGhRYLnz4HmGIGAvYbQnZaIv+d328LFX5NsNIxHe3DOzqU4LXnRNG
M4ss8Zw9TFOaRSZX4ppSS42INyTtKrXBUopFuhcXeCtkgtSh7zSE0yJB2HflkyhY
pCmvLdgp2Q5uKggY+PMVSgQdSecpWYDDexG3LJ3zQ9M/KDcYKkbcZ/wkptMyHKno
tbEBO4wvt9O73twi12FX50DrDDOZzXP/aJ15ZqvIpYVN/WmutbdgzZ88Vq8+ke/d
TJih0xqjuiVHCNeb4Z7KtlWuO8dHY2dclu0kTN5p1z8txdP/07EoPWNTi2RlJSxW
1Cb2UJvUL4TJBBweR8GO3F1gfVxAfcApa3bpDzVOcMjOeU+dLeQJFaT3YTs6FHOu
y6rZ63PJ9r59Bhpa0cdovNhCJpgic/F6xjVyJyjWiEdQRt3bGUKXCtoaLAul1vCg
ClbKWPHM6W1U2TF/DQDnYPn6WLFbzUfathUuQhzKjOmFh7nSyaHh9+EXOD7bvRDS
fZEZv6a87kCvd/t/mYZEMOPMuI6QAlf0XB+UmHHnUNobc/bC0gOmNF8CntIAwUEn
U8lULsOBe/pWttx8UunG+fX+u5NcN6gJ2JkV0hIux3aONqQ+QttV+yb2ekhzg+lV
IR3Dj6tpqYFBlSgtbYvuTpSwc4TnnTBdTpIuMd6XZFBLbbw2rI3gAaZrOj6Vwtf+
mzn7eWJ//qSnrI/xpg5GyNElE8FZaZafQa5OXj3SEZKgdnvKTjOfCwWj9SYIjA2/
ErFhsn22Pl2/f7F6llJ4L1hJFvDd9b7Iubdu3+ru1N/ZAj1C2fW22iMXSekQ/MCf
mQTeZse0TrvTg87YBYtGDrmwr7orfSLNWdA2/WtXmNsr+Ji320KasPCIHxH72PBX
4XJnAct6WpOtmw+sya9qLhixqZL/rypJAcJARdPqfr68be/0DYTExWjij3TmJwYC
f2iDcAX/UqwsTBpaEZ2X+0dB/5UD+jTBUZsVsO4IdXi221ihxc1pm9z85Dun1F8p
auWrUNTBlrXXnglIvUt5h/332fUTQUvVI+k84JBxCNJ7/NEeowekb6PHaH3W/DWX
XWpJHCgiQVI6bngSOR/hVKDQL2p9SU+QLuxE7jZk2+WY+7AEVK17c+VX9zwyMWEO
me3FsSvjYoA77l0bVLi0b0k2iYpOJKPg8XNQlJiBDK06ZyirzP153+TXugtN2w1H
sHsJeH9IP4uV3wd/bJMhVYhebmG2ZfJQWwNaXraYZ26otugLsjyjP+CuSJiwWFrk
98LpQjHfVf/gL3lZZuqRaaxr5+vb4D4f5rptRBT4fuveMf31/qUnxJltvh1wUIia
a82Ck128XKIM4vLwc0Pgm9+PWdAOChhqo1j8eqeeHmutr3M9ZadX/5fIP7E66jMv
45LJHW3eS39AdGT1zX8p9YuMdB0YJPav7qfQexA/sq3SLh4GAfZNS3PmTEKe9ZLy
l11yh2I1khK7mnHITMcDBWBeSmhJ3gYEuSVNJSKE8+cLpUCppcXOoEIoMzVwNMGJ
lNRxgcwOtMh9+UwHJu3q3ANer24lUx8Te9bFzDpsXOpVrME/YsKjEkexa74t9GHN
/8iOl2g8Yz5BooErTP6mNJ4Te8nCNRQSDblizDaQRQdz96kzyzVFj/iYJGDqvlhU
gCXGjSTDDrdgdrVV/LvGycVs9SwiYs1Na0z9DNuaIgajfb3ioX4vQMIyWJXSw6vT
Ui98GCcIdj9hpoe+rLv5iFuJEd1LIZfDSAUev56QY7BQCCwQlesnSB4RUZYHQEPk
S6yhMtqQgggI60CVZglEM4u/08Wf/PRlkHGkH/ndnNeYnGCpvskVQtsqe6aAOuIH
FLOi8Gw3tdTwG8SRZauqpb7JDZ3aweBf3+XhwAAfBNf62/RlFyi7jpJviDhvZSPH
WUvHv1+5mJmwZz1BDoUZ0EF5eHd9ruX393689GZgtsn0N+YdSYs+BLekm2mmcxX6
XP0Rx1eUl/pRBgNyeGE2mYaLiu8Qk65arDCMDLWYwyvDG0zz70QNooIgENtFY0Pa
TBgEcJkH2wd5NMEtOLBO5V6C0assJL/To4ik7oaP0ByRq7I83ZP1UuKvPHCWZbFO
YxYlEwjtzmIreQXFKNHqQJTzVyImX6S4zLJ8a7n/byafJAWsjCTbTpRbFhNxRS1K
15pq1E97WwVyyKgREu5bV/+xrJkY4O4wX4jn2ZtqnAlWy6Jvu4eVlQdpQldOftYF
uE9i0Qrp+5OAIl1S1Lvcnjw6tirzDjjw+y0KyytkSk5bD1zgHcMtODNUkdvKvmxO
i5roZiK9wxBGVOdqJAXXFzMy8fNIw+7G+g5ekzzCbmc+ZOcRYFbSzeWii6F7hKEy
5ZwYDoOPYjABPyi2Myk0aOZClL64Ja9qI0PuffvW6jctx2WRj1XTIjjbd2/6VFrq
Qd529iy1ScOO7gLepmtEDqbg5bN59Ean4YWvZdgHbJhqqWkqLDTnOB5mnOZvydCM
0kNIGFpnUay8X6p+EJ4MCEWZSLEBYPCWegCTMxsyehaVsfln1hXG2+iyDGhEmQEd
+fVITX4NNBOQLw28FArfk2qTGd1g5uyuG16IJX1WMFZ/gDyEz4WDqFenNoBPSOUi
vyM0TynhQJTgXFiP3Lcjrp3YX6vPFu28q8OmwjXecuLigSGLl2j3DBsWARzlmba8
BzaDAy2XvxxD/3wB48npDHwRFqNaLrYVL8liaLtpu/hU7QHaTHjROdDfhaiG6Tmv
P2tNu7iZElt0m4Zpp2ZegFQABqJ2pY09ERi4wiQHYMvyHKIy7ZeVZkrvXDge4kXT
yRFN9B0mKCywoVZ9NhhTGwenrqZH9HgsdKxqxksfJSqin8LwOziu1EIT9T00Eui0
ixZk3EdD3Fpe5YLTdxX9sl4zE7EulOSyhj//sSm+PMEvrUlF5/c4NU/jEtyWv8mO
iquWObWOLr0UGBlGMnKa0OJJA01eRT8LhaP/C7TnNcGYUQkqfKzTlvT0g9weqJJ2
HE3FtXFyJTp62phYcE5BUmy+LgiTJJBe3HQSICDaCPiapJPKdSwHPyzRHyJKYIAs
PgCjQWdSJ/BtOBW5WmdjiyJ6imNskE4HcVsdWTj2vLroHmn63VpdlSsAf3cvwnjE
IslH79Kd8xf4g8a+wEU6IZUG4SBL9Uxnptt1DXHeSUIRC38FmZ4Nj8XqDcPs8OVh
QIoUcyH1iZf7FlYgXQI3mW4YA/XE5XAXkkLweFTVKRfPPTHQyhUHb/VvxfLge1z9
+Ycgfb2rDh8I25uQQDyMKxZXb+mjUOhxu1z3fRjER4G19o0YRmgI+Cax9z9RGogP
lHZRbu0ecfq2JYPiEQM71Qx4V992uxk4SVX6+nXQSFwBXMxmYwGao3ptE3qHJ9N2
Lf9UOa6IcZn+vfFZIjl/WFNOKTZFYdz8EUdstCCdnAUTSMOueRAu0564X4kh0Os0
a/GUikhF2OxsVJSzapv5fKMlJGu/ctgEILC3KF8oP8HGye4Ismb60f3NrBrWkQPU
Ef55nGLB3HAiDf9hnFBtJCHAac7qPjZrGnTjti/xJfdQE9BxD2jQ3LUImpSbdLrC
/tu2VO6Yib9unLWGt3vz5Y2kJq0jJcOW1nyq0acE/4Fp+3+EnBOSAVbGRUFkXBl0
WrQkLAwbPJFj/EVMuFF1ruPnb9b7Nk3iuaNxm682TYUwKxrjj2MrT2R23awv/y0q
C/RkYfFiMf9Z1TxziOAjR6Wxj2WSlQE5FU2Xp/kErZS/zC19cH96u9LnTKSk0xmZ
W3ZQJtL5f1NTVILJuPxqu+u34G16QKRtdthS1Ly06YmvVLMpvkKJvo3ufvB/TK0X
NVsKpdpjyBv94ukFFUAMUghPngUA/MqyTo+uNSYQI030y+lt/nGQHm3Wk0oqJLLF
M7s2Yh3fWKhre17BCV5labJmK40lHSBCTTN8mOFQFz5/FGs9bo37uFR06Gci8hx/
ESR4SIssLlkqzXjunwOkM0hyCwwj8tUN94Spq7rqvWp9PBrK8bU909gPtjGOXlzU
nCrm3B2bFVCfGsNXbb+SMNQV2SJBeYnUMH7uGSluGPYdUXeskQbt/rElqwq+axdv
Swx/RdbHQFO+TmmGaeZJyDqi5/BfvYSZWiu6yF/3T0j67LYSiXLGFaVbzbF7QEl0
zLdkIbQB+nx0MHqyUTVN5Wo0ab23G4FnyTHUYFrEuRWM21fuuWAkdZuElYdLFYme
fMVhdWoK3Xj4AYjumkuV2bMAkgVMLCpn2ifckJ+KkSKj/kV9eeQAGAuGmS4LlgGx
xY00DxcSlgaRblNKnQkd8aSVIEF6hoW0JiIBZUUlytgKs9cHg/FkxDADqx45gD8X
6gxa9DU7XOlyjcNI1HyvK6ajHoYgAH6LaBtpogD441efDIgJltKZuUi6zN9bdiXR
YAGTwY4ryYpVH0ftFQSjkcrAtvtDsvas6cmKq22oaAqUePXu6/RoDoTDZwW6ahQS
TLjaZ+ytgwC6oM/QoIkXN3yKH6y6MNHNNK76Y2ohidcAwKs3H5ago4MCgCFwg72/
TmsVzHi56jn0f+8+O87buB8dImrmiZMa6U7OLR5plqAMA7dtxM2DLTuW4oPUqunI
T9J22sw+1mpzN4aynv6zTW+foKNLdUvlN7qalOhRMwqsPEug41JYX7aXwsH4VgGm
1yv5G4Q2UDI1dciVO232yFkPhYrigx5llwGnPQr+7ZRh06uCP53/PGVAxBqhI/1E
LC4YYNQYYdd9L4ZVySlr7g4wG4scyDSNl5Tx/OtFkZF/VJ47O+njKZSkcpJdytIQ
VK4jad80p5VgsJLop58ZZTCcyBelulGz51Okpuhfb25X7cIMfvtRtI0VFakxRPlF
JImudACmvpBPTeu41bYN7WecYUhPwq5v3dLV/liQf3AejoXtUWi3Kb5qhI+Jp5oW
6/mVh1qae6X0Q9X+e7ux4oGB+m1ehRMcvS24dOgQFSSJFoT+biGKA1eW3t4s91i5
Nh7e+7sx8SgY7QFDFa/YBfYClIHXfS8YvbH+ATVZUw5G5do9Kt14jnRKQ0rw+6C0
C4I4FUbq/7uYQKi6srNl30FrroxaujtYBsjQCDmwcMycCem0cF7zQKmXVvEfghMv
5gA0l3WARdjQ3qkmsATloPZUjp7wQ3DC37riIL6609ZlXhjApvI8ioVtuJGbyVbL
bassBkd9UIL3r840x4Cl9u6gNyWpLXciHrXazarClkD4TrCKFV2RIZWShk9nT4ED
1HUd8sSmjF/CJt0Ztm4txMToGiHykxJUuFbU+5UdFlLtTVzwDV8iGT8k5IG8tA5w
Mi6EYiXV1bnY+KETl0mc3T6cGpCdnSW4+Wfegl6s0Ah4Yd3H4tyieEHytUShlihL
PoeNWH6M9Ed31Sf0XcqmM8wkkBZ2ExvqQVgmv6R+t9lx29fjMr3ciGhwyXRUsivE
8L9jay5NrlZcUYdZ5kXN8EXmHDTjaRp/agqQsunwmt4pioDk3w+1h4K0dN0VJN/J
1WC+AYiOinz042QaNBC5J5o0I+5Xca97ecqI47yEzQ2CWBzVqv3iP5mWeoTXfchG
s1REmIQw/6wFoIGM+tc2LeA2orzkc6sD26VZzv4pXcrI2FpqGJcMltqp52IGG9kJ
DG142VUs9g4y3T4P8RLmTwLawlaFWBciyDqNvnzJqbXHij26SY24TTwhjQ6beAFF
JOCnEOxDHyS0tE5Yd9nfq9tMqq6/2aMwnkuKUKerQpJDDLf8XY20KPiprya6d9j3
aSA72XwHArh6Kr4oH/sYiF4URL9rADSZ8GepnGWx6jQ+uRvXj8Z30yMvNTQ8kZ/K
IqP4B80DmG3ex3NwZwNfD5s5p9lIlJt2aVVoSg6Z+iahTn3pBTmqpscXypX+Xk9n
paGTDARGRltq8aUTE0IvxFMF33khl48rjpWAcpwV42uvcDZEioW4NxJ+Bm2rzi2V
buaYOxkdq3g7+rYsbmGKBW7jEd1ezLuFg69slvAG0LJkNiJplIKFsIizDWeTD88j
XDp710CQLHPwCIgjhFfCHQwx9nxHoFDEbvuwPWPcLQAeyI5HzFvmt5mHOYBZd6YU
6/2Rjq89MR/v5fkBVGWrf3T1OQ5lvIQkLmlWpuMwFV81FtzCowG4zdsKrGEtvGF4
Sk9zrlFZ9byp1n95r9tg3zo5STatj5YLcWo3tjtAHsgH+0sWp1IY9rzd1I12Kw1q
nLm0ZdGOrdIEMu+9U6uQR6SpcOaNFhw1kVn74V67fYP2wWx+mn77EEo8tGFi8yrf
Hl/PNcWb5zsjGaazr8HTn6VDTFJEJIZcOQaZgExd3dzgY6pAqkrtLmpOQ8y48II6
eoOS1Hy5sQ4memJ9JddVqf6ppTCLl9/1eRVPkaMFOWDBR0IEiO3iNKYTsxdJtX47
jzvXfryHHAdyTnnz9E8JpwBIUTZRiJkoBM7cepif+sCOtHKU2aHO9OIJLb5sgnRw
DIumLj6oaSAr6Q8LbtSOGDLLyOaSRIRABAppt7V+mHTJTefFWAdO0zs6TO7UI7zn
P4D3uUU5SPmX/4c+LE3M55G1CnGnimJqqnAiyXhWXweQJRlvALkLfQYOwkYMCdj7
RM6cCs9cOyjfgHvZOcS1MycYExa4DhKjRSQNyFCO2Jf51cljFz4XC1auebDFzzA3
0/zUwMAG8VfhKjhWvSJoDy8K0oBNe+vg/l5Jh185+DDdxnQt8pz/Jrs4oguCaR/E
6XEndH2MwY1zu3tVKshaYR3wI/QfIxn0OZ8a9FqUgiD2MOx/NGvh8Zlww+fbb+y5
lbgAeXO9xTfuyowLuFpN0UH9Y+7TSyAyVKPtQgm1gBGskN1GYTuNva2osYGWcWFb
cFD1KI/ICH7kL6dr/7vFgg4NO445ZRzCBscXqzUHvEMdFfolmdhbqQ0WAoJH5icD
n9JRnSmD57sFPVCxiQAsc84uDhDmYsyYL0kBvutPbScq25kVNmQq/eC8dMY72VCm
TaXpazaxK1iv+EorvDF+ENSumFrCB8dwIOE2pEkRfazoYs4YhUSKBjNO3kHuRWER
lD5szkiDZ0cbEp3U3QVpbAfSXh5vMAii2Qnhsgy1uWRKIuPbqPr9907p3qvERFDM
RO1kihefbl0+1YM/iyEOUH8V8o4Pyp92/dfd7oSmotNPLvGsnyyq22fzcWw62+kb
D3ITOMzHvOd8Xbe+Ouepyhjfg5YP5U0DHfcfZSm0kwQY0na2UelQjRBEF8/NYifB
H/GZxiWGCJkLP2mLrzjA6v4aG4BU91MmnhQnJxKw7ZLhdp+IWEDeMtzpyaylogno
R7fDgNQDDvBKiz47SFhNwGj4EotmLPLWHNhRDmkwpkYZUczgsrRHtOhFlyBqWg9M
JLoBHSnboSlysXoiGrl8RYmCL6kpy3qiJ+g0vBF05uo4eAFh967vddN7pHoXBmi1
TokLuhkCtJ2HI4bqroPUDCWw0vfJ8O+QnJw6MuBPLF6b1owGFo13mBro/YhafhYA
MrLXrSYnJrMl3O/oqQyVasfVsHi81nYAwCMtPm2+N9G86pOSaFWBEq3Vniib5a/t
BbljpZ5jf473f2sst8Ir0MemGQQ7Kakb6qUxvQtNeBVkKNhlBv1sNNq1YpIWAm8Q
FTbs2dlgcp8E7bEzPPa2B6/r8WVjOyX0eaywZbDicFypS9nhaB9cc2Cc4YGJPilV
iNvjK2IVnH9lbazVU3dAfrMtxeouQ2YOkxXaMKJaWBDHj3BtrOBPTl6ASJse0gtI
0nZhFek6E9YbPPRVf+4C0EQNrEQuJ2KxprYm3cEEfvEtw+AEbKv8HPtMK6Vzv15N
AXqU62G/fVdHz/nfObnIYI3he00MI4jAohHQYGMPwT6o4FZYOwHKvLL8BC5pVJ0M
gWrqw2D0vEEPmu+U7KMqYIFp2L58YE5RZo23XSNejzQBNLLgVrMC9sYccms1i3bk
xDeBo6c4Tj0t1IzCFtm0KIun7HbTHlKaZisGGrKk4yfmCXsbE7+U4sxOs5LQcY3r
unSsT070RqMFxPd16tkoJp5pTcAzOTC4ROC1xWrgLLdrXoklwG3ShnUPFWEhakEI
NOSf8TJJXAoPx0KbUDoq4j2aHNouvtN+DLQUvcuHj4OZ0HTKOaH0rlInPUMX01Ao
rnGfbhXaD9yH2PzQkVZqo5e3V0MAnDffqgPleIuLQEcWLmvG/i2bBmRTSYJxFNpg
YD9xre1srOJFzj7e8yx7S2JrWXlMIJlzktwFh/IztZ+DqzaL5dHW6CD+iAV3u+zV
IRLB5UVG0Q/6p1GgNBE2ZWY0qpZ/eNIBBBsJzQGzyvQE7ZQ99PqkYv9qCFEi6oau
rT1wOCBnM/iifVjlQy5QWC6W5ww94YFnNm41udestHSwyGrZqKf5XiT/ai62Tfyl
Y9JAIHKTDtQshfEa2RfbbhQLRO2gvEXlOl9WQiAtcAy+Mv/tq9xvym8o6rAYFWvX
USgVQLkVuD4xvqB0ZaaHqmOyOFIixPIw36WtkjEcuBhNAcwQpYH7yp+7Nt7yroHe
1JXyc6kXFzUwUtMHgpOGurt1gWMh0q/uf2D6Nvrqlr7+skpyfl5RaqBGxciIDPLn
cgxs9IG6SRUaGdawiLg83BLcQIuPBufXPt0Um6hE9XJXp1XTe0/H1DDuBTgH+ruw
b2yyiR9wIdp0Gn9hQuyeWUYWH6UDUzEwbrEU4dA0Dskwe+AlESrddGMaZ9rDci1o
eEFOT9K/eCJ3QSyThBaX9AaSsI5YKNdOr3fGZHRc3tLJLuKEetVUw3LEVfZ+miHP
cIUq3t/6qe5reMqZAoie2pAuxbRQMhBzRfPBp4zolPZF+xDsvDxmlKJ26zhAaX11
Di3v4SZAa0yjxUyUhFOa7l/JHVBpbD/AWsFNeSOa84KjyYAbkJVG4kaGzMDGHkuL
PEVVrWwKF+gViOf9T4wUQR8CI8/zA/Dr29fLR7GzonYw6i+AzLqpk3J0UKkHQXsw
v4AB7m7H7p9g5Ft4eZZ9wATiEW8io5x0z8Td20DXAUAMdBioG2N5sFrluMh+arhL
evJpysGBFckGt/HHouHzplwQxuTZD6a0hJofx2QdHd+l1HLNF57O+b4O5uXpIhH2
EO/rgLlm9nUuBNIGhDCaoKYeU9jGWXvt9lbjodnAmQRlMAqWx+JASv7kWQOiWU2M
o80TIq0azCm5aS6Qana6gAwRKW5vSbTOt9a/UOdiBPDGjQuLocpQmE1C2zRc3pTk
oe43YW73YB8Ey92oEzYXRv2PUJnqKIal5TfYEbq9OQPJ47FBJReivEE2pAoLaSWP
rS2KR17ZDGccTg7fMhiL9Rp0edmENyw5IaJldKKp7YFT7N9xc4IqUsjbWWZKVy5z
C/GiU5/FDGOqmkORY4viZL98ygxLO2mF3U704Uw5VMMzK/tW0HaRGlZH1hVk1bCq
NQqJdUZmiOMQ6HHb7MZKlPnSuAfbOkMHLI63ntrMtx+2wgz+mUVYM33pOxsseXPq
8Xew6sz7sMEQPdnBnx99XHKcjUwb3UoWWcctQ4EaF9tpa6F9gpIJ3KPCAfL1LUpf
OzQJElkbvL3G4SvZPDlyFLfJSJ2wYO21IJO9zPRbAeAmxjtd9IH1kQjnw0dOVIhj
u3PJwONYKm24wjO6wVJG8ENRHFPylZ1V/rIhRYjNphQnGVFu+wgFKHZeIz0F+LkP
x3Vb21YjCiwOYk045ds+ceByW9gdkmIFULW4C5rPFa87h6DfzGbjnVyxc9gto4s2
/aJuvzSVMGZnB2B1Ru/CIx5MZFpEmQawyTH8tlpS2eDr6RZlazDNSM6MvFpJ6227
c0JKx3ANhAn8+f+t5Wstw+6jsCfuIUbBdMVi2EVQrBxsv1/Rjq4qmFSzVSXdVzQ1
+FF4BLPzyxGa5QPsPAqvEGUTwyj2piREjB8KL3kI2nOx/lVKgQ4q+h3VVutDXjwe
i4LGycOqhXmusybwqxBIpNavuIbRcbH+YtKMp9mltR/+tJbV8uoAg8BmHL2zMFMf
v6gEkEPdCYZa11BPv2zWrHSvfEHmqIJ7tYfOLkPo7sEmCHNWkTYi5ZD84BAX+ny1
nx9iVdefi3S00cMtdiihHhVIN5oCYrgkwWIBpr6Y3kEvHlMSKuuT3o7F6odw6SaD
QMwkBdM6EF8M3vkycJ04Hx8MtSU5y03zV9IO1oRPmlouISw+Z1gOdJX9DFoFNkVY
k+sx899+91bTGsZU/LqD9OiamXg+Hg3RlN4/KJFfuas/8ZhknZJHldwpMS3WNcf9
y0I1atmxL0s6HBxUAziFQ+/3IuS4ydlCwlrlKrwj9EHVwkMc6NweyzBrXO7bgxak
GDqkRqQf6mHeNOQhnlHmvCZjk54Mqg7G9GZfTk2TRyW5N6EmfNnwYRjRqjUvUNsA
aB6dwVeHN2xsVtv3cJdFz84aJYCHKLTZWEyzMjHOlJHaIAvtxmCdg2h7XMhg0qeL
DCS2xEzNp1E5SZaYF/RtQjhWrhCe3YDqyW/M8K51JYsVP9XZ0UnAUWTbE+KcEBGq
BgANv+02bHjHzBsyZSSHNgldY1DaWsoBEGBjiSQq3FkzEZvI6s5PRa3nnQZ2r94z
i+8k8ay1O33yIoyUuqB3koVJtHZB9z0xuEv9/aktP2TFn2MPpOrPk9rEY/K3lJjQ
1BSdI5aP2/tnXH87LU0GK9gpdF4GaRTGNfelNkJT3xXTPCAQ60yHG/0nH7wnLdrG
Rq9/6J7PN4KhPD40w/27J27l5UEeUA0hie5fv2uhIU/sN03jqPSzKC/oATeuBfoy
LOx0RxykOYq2vRCkQQYP9jIeuRR0jw3OMvNUyai7CEeQUhTHibmL7nyhTTeIvjlW
6gBkukHZjkd4iPOQUILiOpdTA4REd2IZmA89hnIkvBfh1Q34Mb6+XW7AHzTWltzH
7GSo3N0zR/hxduq7gOD4N3lq1iCMOklZrdRB8WYXkDWQiunuGnVkQqv3fmpYACXI
OP5RikYjr0vVgernF/nQW438U4pScdTKQPrlAf75WPt77sL0DLSNjcqckoqOYNM1
IMmVsZM2sNs0ay4c1UX/PbHp3Q21Dq+op+flO3b3BThcVLvOx3SlK82wsA5by3X3
E2ht8kayPqXmCFUbKpT/udC2XRuZXcHrxTTt4V0vPzXrPbeFk6xjU2jboCvLxOA3
tjYLTw8jmF5gXJo1mgE5R5zEbxLZouTFCG+ZQH8Hc4j7qbGZxSuVV8OszUKQ3L3L
zk+fkffWi9/OB6zHwOsi8viX2KRpYYGiPioRN0PZFI/1RKKEPcYDWH7cWQG9uXog
qftnGsDJg7H7f+A2fCUGkdlhwCoD/URuoZG39YUY7LzW/2fwfVDw4JIyTEPAsanA
7SuAnruBokX75300FDTS/iamu7SyHMNpo/cy5pfRTadSkkLfaKGJge2HErh22+rG
Vmb/CD1d7NTan8oRWjzG1NvqBtkeahydvzM9HEHO5P9/Gch8IlcgIv4lBHd5ouRS
KS+gr+YKaDyach8lYh20J/Afvoxs7aBS4l+lzKsiG1zaCAV4Kfchv3h9RbTCff0E
7Nl+Wa5CbcsyqUXGzDbaAtF47AUsf4YSXL+h/mr/GUTZ0s0OhJBLiGVGfId3LwD9
99z0DjZK2FLnaaAnjmaGqkXLuUlnDeMHJCHQCFZTlEIsC++wYo0gSo1ECxBqbplF
kxlrUuWp2T4I9TsZb+aAbIAAi3oWOZwC/FJOtcx3SszynI12o/lESj7+YQ2dETul
RXveMuN9Yto1Y0tPaEpKY9nTYFJVkZXJWYDzImfR7P6dvGfe28DrlYo6r14En4SA
Gsy/qGGpTwFhnPPOJPRX4pVpi5eHtf8SKbolFw10Vghrjsco620Fi8nYL6N4tKnd
uomsQfU8xRyWDf0J4mVLPWNf8cZljTRH6WhfkbEx4t13WnlM2EVE8AQy2u0xhYe3
rEXtKLcnqieqNf1a7LhAUTczt0pKsWNdrVt2Lm+l9j28jC5kQPSDvTqSPU2FU7Bi
Lhw9ADQICM3GDC2teie8gTCmWsyuJ7jY1vGvJIqK4zDMzgp4kLClJ3agB4LCTCfK
zocWEn5llQsuvQO6GCPF4UqXoHkY3l9ov06UPOMOR/oRcqRBc9i7IIVgSpfkA8Os
34J91afhpmiUS3cz1wgxMj60crmeupIixLktvIq8wJFjvy3LveAAugt0dKOVozyo
pFfmg2zp4lJ8AerAKVh0ZokmL+H8ctKyZSKU9F/hFCBCyOamSDqvLC3BY7VOur4M
aqq29ry3kRJVP9bXwG9W6IzRrAD5i5Aln7dtqVUsjqu2mOGWsG7Geg13Fj0+skPJ
pV3SjejpeEf8pFXVm5xlmsvKbFQ6BQfVantySUXPRSet9bnzy2NT2/SxXt0Ry7FD
2Nrt3Zfkz8v098gjQzV46zdAPkZWj7u9g7Aq2vK3pA7wg0kaWMPDauh0Jch36Kxx
2wUJrgOQe/8Kp/a17cN3ZeL096hy/SvpEVdToq4H5TB0jGzzP+MaTT3fSRs7gFGb
VOeKpYKnoLnkW8G/pUkI6x61/HolOdwcrSugBV+5iP2dwvCi3KPHWAY5i27sJGd/
lwWyIxHWAVrpMLxOpknpCoBvbCOQ3qmneT1Kw6q/NgGV3wEAIYfrlBl4f+oEwxlN
yFhUEcMRa8Joh6vCiYX46QuVk05OEe+RMeha94Ci5gL56MxmkWLYS6clzZkRHQt6
H17NOA9vjjpfIAFJ/r4SXrU7R7KkGQE+Ih9T8nYQMjuulg4WOgydSXgv75abe32B
HTa/VJaGCz05xfTosBkn3PiKNsK0ZdnC+ag70eyWT4l+GGCvVO3VZBoH0AiRF3Ac
qgDiCL36152+yKzRI0r2pB4lZkxuPMQmWRH8cfivomNk3C6kNU/enxdIHjcfexy9
TEIO20boudFNyHt5SaZ3/k3tqon2foQxpvvSymee4lTqdi3u5x0OUeHJouJA5ZlR
msvLZuWc2mH8ZO32B6pcP3vBTWbk3XbrPzO8ZOkFjlMiIgKaE8naI3pFzny+8lbj
+zi96gHG1kCJskaGC9/O/REyj1l3T3Q85t3ip10XwT6wUi5KjQXaZHzk1+TUd7+P
d3YIn+NwKC/NFi+tKzb/26cVuARV7uKyA7qju3yJbNRc/Hu+gFleyvAbjmnpmWRt
acZHSVFlpBJSCV6zyxS6RQ8L7MEW/tt9lcENReZrDFus1w4+wkvAW8wis8XS+Qd4
wHqnCfNFCdCutD9w5RF+2dsId2SkWqon6x4aJ3eSVVleWNRTxRIA0f8xS4Q8t8PH
eSCjn/mmeQGOTu6Nq8CvKlGTNhLLQO6VWvYHxWbDKaIAfCHXMlDWQb/8ObmwuqSf
xynGbZGP7Cg9qicFK8Q/P8TsPbZL5vC9IaBgWe8dhDwmQk3t/sOfaXsLyzInJ6Mu
xal+JlmDXyQ+GQIzxf9zeJZZtDx5AsxvDEx0NtPc2+nM329BFwz1QjRSvsvZFxwg
TZlJted2XdHexNZejbomYo6nZU3jmuOrYIYXFTublAQ/9iQlveAsvwz1HKbLcE34
RqPGG1xUwD+uORzCf0HIzWiPfVWtFHyZE9gdXXVKh7kIK8/wHyzDyzksIFyN2BZS
2HiYNkDiF4OHTbInMKiyYd5iY56rOtt0wniYv/r44+RD19KZEBQL9+VEwE2GWfwZ
Wc2pDRiV7wuE3iSb0wdY+lN4O23c8CewYYzgGQ+daK3SEl5zWlLOM8o69WIWNh/x
vFCU8sWszQiUpwo1Z44PKi+w+FN7BM7FxVvSVdztmX33yvpX1a0LFIPLtuV1euoy
NbsM50x6WDl1MaFfnf8uBbBIwsV6RnmqrFw+XCwuaBaBEIrnkQz560tCMmozuSfJ
F4Tggh6i1UhN0G1YFXqYjpJJskyIBLHUkL3toOP9ln7KJc7ePHIWecT3NEW/LM85
Dd5+hj5OSEJLHTyDdhCvVUKHO78z7JFDMwUVGQDKQfhHrRKao7nFnkfj1c28HeBC
ETzvDOCdkFnRtfEVYDMQRmTMi7cFJaAW7hrCLrmi6ZF9o4cTrwfSD/TBCvryag2w
hqgjj87zl2LbIZyX18cUNvtTW4HShNKngBhsePkoU1fBAF3alDgrzMwWgYYN8Y98
8wPdYDr/l3rQMh+YUQHvCv7RCv/IvSIGHgHFV9Upuo8qMHpwHadExoh/2CccoTnc
wnFKCk9XclIDuAAramUa/wJ8pziHxSSYkD38tRdYDnDsxnyKsMy1SlTt0Xo4qL4o
9Y4HNdFJQ1GCpVUmN8wTff68P2//dxtIuTapvBI8IHqYJc0xK4ebIzqd/btazuXk
JigVdr/6bHeSvmm1lC3FeFFKmlSuE88OOo+AUxyr9mUEAX7wisbOSxcYB6FfpXkr
LaUi7L2lnUtSL2SmHcyX6PMpuld5IEqBnQvjlMVTonZpp/JeJoEjaJSyf6yDnZ05
VEbIHWsnmquhfx86ILBs3RYj5W2/Ot95/V9+K+ZagMBdJV+BZCVTwbHqSBQ73AX1
++Cfu0R2jlKDHD7/8EzklKo1cM61taWc9r0CYGRbzRH1HMhHDboDj0l4ucsV3L6e
qsEMiTopr0n1h5XA4+t5ZQHZgpgIXEwav5hy0oS0AoSYU7w3xYFCvz6RWG9X27Im
opl/eip6cExqLqRuRxzosrFLE2kx4hxlAIdgWw/dhLeT+tKXfkswGlXVUC1k5iaV
f5qUMlSBARUD3z6RocUVPr25VMpjYxU+cwXBZnygVBLo/dPwPX0vcBTVpgOWhHEl
fRIFAK5yMEbFaCGkbjYTe7DZZUV2Wf9bWyefKkmDyOXHbDyvpHaf5V6bbeyGWGk3
SeAdTmScOMGrKRmBN+iJheaRBPGBtTftx8we5/new6Rbm5W0xiqGZN2144pISpJ6
7fB5frKTEcad/I3RALD5gq0lb86vgA9YOC3hfrGETlYSEiPUoTdsHdHDJIMm3qh0
jTPWeoW3FHI1Hf/CojPCencqWjgFtTeS5npNM/pqVY6wGAhr+uJqRUBj2osSQuov
PYNH/Iui0+pokyE/8Cezh6SR+Vl24+5fw5d6e4NpOAqTI1z30Cvr2Z1eHEp2XwO0
A1BnmcD4dAW/DgiT1cYR8hH5GSnRNpppf6/FPVmxRgy8bg5O9wkObBO9tZQ7hhr9
lF++hP9S4PCcY2tk6kYMSpIaUCW8Zl7nFG4WxP9zcQvbr+zgq/R9OhQMaoVNMHZU
s49XCQq4d7d7uJ8uhfFFLbgVvq8EODkp4L2OnmY5BuLou/uexBUidTdj6BLFyFCm
w0VrBtby22s5oM7RJpQB6XEzG5Ti4l92419eiaTwcGLC4IYTp5ejrsItjPbL5Ei/
9iVdzYms8kXPoczQCzzRaxVgLiCJKv8RwS92U4bDNRrsK2fcr4dtZve7dFcMZDoc
6gc+yZGqtrZSmV5E8SqSME6kd8uOL2rxJim9nfl//ci2Gs0/EKcDhjvlzyk3aX6T
K0hCTzBOZIsH+oapSxsxRCL6Tre/IQnTW66gkdBaBdbpVk0hy21BKAd1VDHh7mus
1eE07RFKG/fAKu1SNNP/VwE1jhdbI6mJf97Z62y6vyxyLeb9suXQShfrMSn7+1Rd
fGQvsh3zzj+jB9s4v21SY4K79UoGKDlW3Nf3x79Tsm5IYk8otijFzCGQLyqdf3rk
m/1NEzvrPjxCKK6zS7t+0mNSePYrIi1dan1Kc1WxY6LcsKdYrcBhbDCXXHNd4VuB
TLsWYCVP8pfv8HgWYkDheqq9YJ8OUYBkKt0Q8IILPm3JxqIMS9J8+dbBDDSNMk2u
WkVKRAABbZyjrZsJ3mKyntA6wriVSGcW33fD7zrbFNVEJ4lKywbFsotMjFRGFm+T
MWL+5oLxV5WioEIZ3EMKPZL73uUXfvkWZefk2VSig4gnj2e260bSyph9CLoIdLe5
dhnGs8jJkH/v3TXdEhD67tHXvcNNb+SgC2cSpFwqOvFJJsvPCGfQgGU1tIE5ce1Y
IpL31rz+/QT/qW3MFHb0YLxxA4zuTzPQYCxX9lHpqR2iMWJlGgvsyRJI0dztyosn
+h9uvTRf2xnk5dGaBr1GrcchiHmQNkFVGOexOyT/bYEEl0hSJB+zoqbpsAm5GuWP
5tWikak4u4EN0ofNAnM2ZyNuQVTWotgAkAP+1x6ujuapLeqyM3UsXmycJ1iZH50M
lbnxYUN/AFN2csm8kIFv5UtGB9K8tCIP0L5PyO0tG3oFtm7VGdHSIYat1ZpwdIts
YCUUNIfc2QOaBm/TXhFmhA7eA0arzE2XcW31gbXSDrnysIqyuij1oJnx8CeCPgb2
pR5lGVI7H86UxtRfdIhvjdbR1+ZKKktdnndPWXi+gTk/qigC1S0LE9ZXttvRcvrC
VsW0Ea+eiciCx8p8WrSuZxTXXvKhoIG2YAgikkoy/ZPl8DpGvicv8TAsoqy4sI3l
wn6h+WbGRKW6JFwOZlUEhFEz+upwhbeEgLih/hn8jMX5KO8/0KNvVRkmLBp+b5cp
BZdEfsqdLgoa9inyZZyNHE0y8mVwJuXWot1gIxXy3+48AoORO8jKRi6VcB6Y85L7
FmtaoPEQslvkaLMrZIkFoqvONTQRgMwg8ra/4H59X3NqnpOPk0orpR9lpcpz+K2w
K6jtLxgoSLuK5FVcWS3gg4knwZ8Z4bKtnM+7dfghYJan5z/JZpR1FdeklaS6/nd+
lsPphG/tsFgid0LNMdnojVXCGTLz7LeT1KzsaZoiTvBgXWb+gbJm1tzoQzH7C6mL
1skcn5gYUbiMgHdam2nnNdkn6fG4QCDrFC6gkf3coXprpyXIeMhbbPVe6j5R4Wu3
70U82qK83ADK5fo49GL/Q7xF+tyCKwDOylccdOSu2l3dugsxdkjBV6gz173NTLxk
AQCnuzTsrxtB+rizkgjBxE7obtQtW2xQQ6TA2fzbDFC7HpweHLyRFrO8LpdXC7x9
gcO6u8bsV7NC+BSl6FJnQ8V7aXa6Xr7WAPGYe3h44R4WEOhxoc32hWtLpukTtaXb
YZvm0lYs1rxXOPzRy96OtI4hhz8t+lpVYZ+bYAqttdg38R80Lzu6GJgdck1loQhK
VMcVf00yK+7hnwSnbXbb2oNSGN4I1pRnkOEvVFck67ElloyqtuIXFT8StsrQpbdv
DdKCcqpOcBuNcI1aqRokfCfZzesThQnrfiPJnwG3dImbb/UTXZdX++oXovyQcxC6
krsw7UlzJ3IezQDVwnqy5pDaQRjpAliCZWFpAmRa5E22nKqq7XE52XHbLddnpk++
tnLgJYeyOHByGeRcHaFpvOdUpKzN5D5F3eDTgL8PU7uucBJV9VHqk/cGnbrUWzZ4
Rd1hOD8TY+X2+8AjlrnQ1azHky8qK4Pqg2jnwuI0uSqdrgdHSn097U0yWxdvnEYt
K9DO0Qdhq39DuySBEjUGNaGcw+NGnorY7PQbKv1ns964xAAF7K3kmoM04ZDhRNy4
Qc8yxWiwokcDfEgML8yNvW0+qBgh+hTGyHdwezWm/5U+8w02Y9/e9IZUzlr7gdx6
f0/DU1Ow1VDXaWUmGb0VqfLOk0/RmNW3jPwQ7AMDMoZDvb1w2TwDkHOdCgHkbmNj
XZUJu/pUt3tF43OZDoDji7UFT1H0cnoGIyNjBBnmNi7C8JQzLEt7Zyx4TX4uYYxh
tx212oHPXVcnEMxhfiZSLVRFAKjHKtzX+RumQc2v3yy3BOySondUTr7JFdY+gCAq
YA/disVXD9X8Ljxsix+YfG5c2mXv4y60tGqYvWaABMakrclJcKTu6jQUBO9fu8NS
yZGgWiHgM5JTwTtas5wzpQXcc7WYLEH8ldXqj2S00OyCHCizwofMlZjgKqiGqvgC
vfePkbNXPmLeV2FSXyNKiUahjhtgv5MS4Ussn8v1ynJLDW5rw1V3KN8gCb6bd7o5
UOKNWyOeEe23OSjXjhQXfaBV9xPe0hGFSCNSGOTHC3gjHFk2CsfA0mceaVayMz16
vH7lba9rfym1+loVUcndjGZWJcFQLpvLcEowW9qk1xZOeCoy8y9tVR/6KWNGGQPI
UnQBHWCBwm//Ht0rCC1opzTIfElMa9kDLBRJClRFohYIklvEg+JjiTXFjrrRFNnk
5yBMgd36FfFhfor5xldJ+7r16567PaYGq7vzaKneWIz41L6VFIjfhxJBUrQG8NCC
gemhM7i3FXsvQ5gnEVzQ/ezGLT6omuRSC2j+hFnu39sNLteKPxln6ktcMKhA7UlQ
1zzL5TLzo7SnqSgiTXseBLrwXNHTk5QdnUjYLmOHub+LKbzxy4KME4oiXBIX0FnK
5rjgbMQoYqfi7wCibteKHWsCOzV2MOTBPXbgOCcY5uA028SQIQ8eSmxo93EhTCyK
DG2dIOSSe6SpUNJ0ziJ9Eb5UJnKaAb8UXew1rvcVkAYRniD8NOziIcIBLN7qg/lA
qi9tajCQG4zwnOsbinHoww5qX38/hyYAj9o251yto2DZvwtIYUr0mrjP4XMpFeuz
GGwrzhfJrGX8S2pePolW2z/iQjuEdqBrx/tH0QuZsJpJ9y92Qt+WZziYmHsraWnV
S4CqQLZgIgnCTuQvaULNdYPjS2NCoRr2IBBrS8TGz3upTtJAEgJJClsM4UAVusFf
aEllwr4ZArcHNJMRc+1Y/WmN4QnCgwtILsFnHUDuC2P43S3Q1dlbRUIhkVvSPiI+
6m3rTfZCYaSe0zv9H4X7J5vchPMJUkQaEHonBP7IR9xGjJp9CiXeenKceQTJX4JI
Wa6NE0dcBKz853OFcGaZ+WMDlaeviVnvgijqaLa5RaPdzSwi3T+6VwhdAqRgikHF
LFos+UNyfjBAJNz8w/lXVRlvPbv3Bgmb2gTWukm9iScT/DAGinB4lo8fEITmSuCG
oOq4uMMIwCQiz5XhdDkslu0RDwgBzB9TKyFfiVjfM2TC7HznHOf2j5y/mUpvKcBP
foOaT4klPmx647HpvMkwze2iMu4miRLDBmyfkXRE9gWaa2F7F60B0g/N3UOkv4D1
oQ9r3NVCZa9Q/Q1vepql+vQjfWunRqwntMYs9t/Y9pANZOdtmyOIrpsIAyK40hp/
ey6Ot60Yiji4QUUksaduFFAPJgRMB684Cd/Lr5/0AZ8VuOFrieNxroCv6uGBVuNX
2z271XISxQeBM5dW0snesSorWSB+jO67AhKZ8FKxZXH5/7hsyQa73G9Tv6gMfuvT
i5j48T44UsGPBIURrUU9zo5EnDiNLxRJ6lgcKp6+GjBclldPEkO9qoJwXrl7C7Qr
zU0hPjvLWbbqJPbH2o9ZTeIuuVz6xr+iYkw2odPQ3R5Zz5B5JWerpKtGERdyvb8X
kMnwInEz3OcajCqzk8px8lArKHWDiFYoRRonlW81mhyEl6Q9amPikiNrgEmQ8g/i
2t9MUg2fygc8Rmp1e3fSJWXzGy3tkZ2uK8qJrZftc8xqN39fDcCW0Hp7clxVVpYs
pjEErG1OEJ5GHD09D3tirVOiGmIPRH93nXygSojshyrtF4tAOdF61Sd2pN7rlqT3
D0JJEcN31DrJkNYJsapcT18chUuNkXqUB88+/SgoVDJM015mNifTTLylTcNwsQLb
00mcDdZIzXSp/rUnsvX+L0sykOJVwtMBK4tGunHVAJAinc+8I46W4rEAgNFI12tb
mmhGgFjbWY1RLrl07VLe5H2dPKuXQHLVzxWQyRiqPIA//tcBLY39ouqizYKdkwrU
K3ln0vwB3V3vN0Bt3UoWpB1BFbQ1lh4wlUQGz0v2+R8ApZyDkQ2ASDvGpnUuOquE
eP4wi5g/ufGyVH3SzKS+xj3Zvyrkxr1y5wvXU3JrN4eZRzsoVhitGL1FSY2mxils
FbcEhezhm2eztTsy+y3uCR9TcGdg++T+rboNbmEbRugu5ZaiKxzje0kmRDtkcL/m
2tqI5xlMvncj4OPE88hO5FtOtpjORB1m+FcHjot2XHliitF30V6XBNdOtfNDS6qJ
miwY4jNaiCt2q8nKrkkrHcjGi3BXa7KQhvH3zahtznbIcSiN+74Gvdr0BmUis7S8
q5yWs5278K6i++wBKi3mr/eemszfLIMfiRLe7uJcNLgGC58FkbGX2ohhRgGJ7zVO
ylsKMUlQMWapOreerhZvMavN9o4j8u2KJ927LyzbRW52+j95/uyTSnWH76VWCNSO
HykhTragWynm8jBAc6BQCFvfMTv2Hn3jiWu3MqdMKzzwvnu7I/4rekeI7PXI1wmH
I0ICoB/GEEPVDbHPF4tSV3IPhBId0cesLr7zkV0OU54pCcrhV5pobeNh54XdnoOl
Pjug405UQSKo+7IhKaU1rMInq7PecHIRY03wuE72j6xvcLonaykLnLXY4Q5QF1Zi
pHd9o8LSbvqQ4fMOIPu7LBiNfVua1V8nXa9R0Mlw5CpVGLHpactE4wY1B+HnPXZO
uaaUUktHiSawCla4ULIV22z5LZBnjS2TiH0Cpyy9XO6ejtxp5xYvUVlRa9tQVmsi
6Mfa/BvTDs59j34fjmk9UZcN3nt91k9hxRCUdsFmjkw1UGneSfILB/3P5XFvesx/
5Ac9Q3UlLQoLmPXJcj4A/VMWE4ttOgtFFCE+ZtMZFjYrSFJsvbpweOb9ehUH828P
/jDTrRo5B+KgJrwBWncARDcCyAeo8Ze6LAu2fXh6X2AiGSbopYmjdYLoafll+pxh
Mptyt5V2YGw6nbn+r1y7BzG/oCWXkUGpIk9zI3NB1LDFWY1lRlQFsf/T+ePWW2+3
FyuZZcs05Y6eLglVDdgX+Bi3K5E7pryBNYMmHjkn/eClAIRAfWhj4Tr5wUv1RSua
TpDZTb2UgwEEBmDns3sY9JLDRIR5G6HcXZ8PX7GS++0ckVySdn67bwomDEtefcsZ
Z9pg0xQzd65vHrU9tfebsY1J+qQP8xVe/RsshM2bTF7RG5KHQuoiZkZzgKmF0X5L
ihrcs8HybsKWkolAAH6XXtcFpTRCRsgQI1+9IDYxx0BW/3qldEy1D2HYzv15PWhI
nU7dmA6rnO9ush+K2jt0cSguOxatuNbUgTzTp9iwOMuQQw57Pwb/BtedjQQVicqM
V/oB+bddzSawAuyZjkKNIv2ozfWwhDqR5Qv8o8Qc5GAC3XKVwOr/6y9S6Tc+ofED
fIJj4VNeWJVKITEHcAb5eMRDtgJ5E8bJYt/mGJNhvKRHgckveG7JGdgAGjQEPfdi
YkrfIPLhBVrO4nCI35HPaOdmQ3bZCBhKs3yJo5PB4FGhm4O7bNpgfeMhZrQEPVtH
V1NxAI/FMTQ8+Y5vNTWMpSMTcxcq+QvoQFYeCAXYAMzex5DpTQvqNzxgrVZ+6ztZ
f4Nsns3how8J79eESy0I5FVqJ+XTKr64sgSlHrkhfJ4d8hRRWLDd/I6xgkykdhVW
lZPxERU9nxPIXR0LJSW2zjcGUOATzcY0/Wh1t5NY9iwBnTKttR91twf1NRTVrvRI
e5k5nmHTaZodVTAaJ8c3wr0XiOIg3p3qmvXDIwThI61Zltb2qwVUFZWcUaJIxmQs
705jZLQjjxOvqYjxpdyVTBFb5GmlUX8171+B9kS2jaqiGD6rHAtQ/FWbLNeTPOu9
TClnRQVKruYFnSpd04FzOlijxVwUPqRrjrZH2PQCXhvCHQWYWQ4L8VgQh8dTJnir
il0WORXweIGf0Ae3J+XflGlU/SsbJHioX7Vr1eWnjRZnZlWc2fBryGSwi4uqESiN
mxn508PuiNkGXc2q+AVt35EJl/SwXq5+xlwx3A11WaF2TBg/ypWmIXda/V9U4l/S
/XheLT0UVVwOB4l5e91hzlLMmWNAd2R9qhxIFodTqO2rZQLBubCIQNPjY4Q45a4b
lmRt4yjzM3l9PEMtSx1iRdVlmf3FJpKvyFrchu662Ghzh5MhUuHm5hUaPTkKd5GN
saWmDqu0GTKNNqzypApOR0HYwx+yPMkAdm8Ow5FZ7SmGUn4A3pqztbUeUJKlZFLB
l6SgkHVNIrR70xrRgQk2eO+I428yMIlnqQF535wnx/lP2T5MlwoghHgMQeKMAHXT
ErAeD2QkWn99z1vCpwuuEQy4kPr8HUQUGDC4G4s+TlAAaEdF7PAcOhgHMCQzNOcj
sIpskb5wZb1HZx1Q4ONwFqGH5dhxvabwJod9uRLN9OYwSSo3WODnSEjpxDjzMx0L
xDRM6TbxAXxLm6OGkxFjllWTHBUU25HtCwb7k1E/1HSzs/eoU5XRXH8HnbO6H/KU
4YVpics8Cb90kqHgu5cCcb91CTYxF3gOB/E/Hh2OPUkYLtjcKMzYQUN2kB0rOa2p
by3QjJKRiC3DZb36LURo9yTcGVxnC2P5EaGLTAApRRjp8/e0mCD2LUNxarar/e5B
Z/qJByMSTXcEiKTR5qOlRBc0jiaxEUlgk6ArZnxwXttkdHiIAQZBphW9YlYRsWJp
64mHR+yz8KYmBO6jHAGuG0hNu8C/OXwVgLO3xGB/wNTNJOqY6D6vM6UcHiJZq8Ni
xMOZAQ4hHGssZmvUlLWUnMN3vGfdrOMFywmEAGDF+BwNYr4SMk/y231hxDJ97NCE
hdo7SrChsRvd35U68cMWirXax77w2oUxnBezc3lYj2/oU6mBbx5nwV4cAT1XiwzP
sVZfS7OwdWTQWTWQS72dWgYN6h4NxaCKjfEE+DqUKvR7eXVPPgmtuvmCd9PbEAYG
yMN9lJlseAyFZtx90TWxFj221Qr21J6OLQ/tLrKHjkKTPZ/cxT1/hBJxKaLE3J5r
W0mmzWJF/1rmK+ZizocgLG121oN37t49qy4QLWp+bH2TjAtnN2RcWbRmlWS9JzJ5
e3hTm6PeeLHPNwX8pOpUvthLAAB1SKxyWJdLktBjv3lyirYpI5AyGms2jjbBPWjE
ES9UQwcpiC11yn14yp82mOkEZO2Gu1vDH5JMTzDGljrFSDvdzh51uGPdxqxEb6wC
sIZHtJA8mPA6yCUv4MT8IV80S+96ipRS6CX+LhMWxw2LnnEsYJtnSjLBIdZlbJln
Ey0V+jxQ8y7BrF4LNLBvwEmpZ5485JkcVIAOXTrtkG6I1+p7FwGOzF4ve6WMkiWe
K6INSEmbANGv/VgeTUjMNuw9H8wzFv2BrY1+PgiORhrjsNn7rivHlpL0GrrtJ27j
stzKKmPfIngExjZQG6L5qLRSPFUbtvyuIyf+Mi+RoAjKcN3EbRD238CbH+pE+yrq
vRUl3agvvA7MhVLhSxAyG2hFJmPoNAHX7/q4o/Hsx32Hnb+OVaH4psplpeSe6r26
Up/EU0qlljN+5JLODLt3OFdPPKo5rO+EW/i4zzXBhdYP5pHyyk6C9Ds2yONlqBzp
qE1T7HlbcNX8RSfSyTe38x9k+SOJGC4uGNxlvUw6tC8wun3RYfDbvzD/vsYME2/t
ur+34q4kNozRJRQ1dQkkTQwQ0Aof0Pd3+ibdU+esfT8B5EqZddf4bwfVo8rpkMIB
EvkrEAIWtw2lf90IlsrmS+aMbGu2tZ/CSbXHLHstpdwbaMx4c6k0f/yDcxTJ3InH
4RW2HlGmMM09tE0y281EQ0FyvH0op8ItEcs355KajFoETMryKbEJC+gCRqKYWFJ/
Lh/hjwXWcQ9oR4u+ld4FuyOYRjgjtZun27Riw6shp9hNYckqar2bUBAMi8+zcUkn
h28RjacVPlfxX9x8qMqfEX18MRUcv4z9kgXE+hRQpIKkYeBCZBwz+zxjgHozvnXI
7f32NeH6G7Z+JmBVaM7lu+CMEi+NUhk5JoBODgmtVlB6f5zLBGAUnJPISeqU8mF8
94n4H23uYHMvsbMRzBF3OapfF4AiLjWsfFcqp11nWVzNIYU9Hi3ThuCe/jeIBCBR
l4EkWtKjXt/CliI9L4gNyOdrYXXvcg4CEu7iecG+zWHFEnd+NgTDycpTu4eubz8d
n+cGptKqGZtS6RYpfz42vovYPfvFkglFwNVxiwAaCkFWEsNRNfdy31VQFo1ZMGid
b3jiSyh2mq0uI0FH6nCCj3LLK+O6Ff35tz/M+VPiAk9CDo4v7+cGBoquE/U2MPoQ
h8RTeY58e8Z3XNaeWpD7zt/SZOr+NQNbnIb+TcR4UFHyQKVc+wBZnASXTf7yIL9O
st6a7LyFmnPd9vYiuRmxF/jxR2p6tmQv+JmRyc/ufXG/9hF8aQ83mMNawomuywEm
U9THXG0WvQniJJhMd8K8UkmXyLnwZylSsVBiSbuuu8Plsse9pgaaKUugmzwqzs2a
nzd+e3GoMy1wJ0PaeXWNftqPagVWSYqsf4G+Sfu0sjHQDqJ48tb8SfqmS9MpeLGt
TsnjgXHtxCqO41zVHn41YzvIq78cfiVsGRkNjSEcBzL5NiBXVvKg5Me4DIbdKHzY
6/rjQt2t7H6sXlKbdEeBbxDyk3qZWR0dEJgnZnixj0Sc7MgpWQCT0uNX1Nzopa43
7caXfHape0JgKBUwMbPmK2cAIykWUaV4XUfSXj7BkQkGeF2JoWbTJk5f8r0nCeMk
oVjScILiGJTDLZtTbJtj1Tx9jZgj8HHUSwKYqMjwIADphOBtCLJt0p3vbImlmsrF
FxN7kRCcXa3Y8iTMrVR+scpB3LqjlnX7fZDWmzZ/aDRAbswamKKxIG0aEk9wJRI4
SnnJ3c961H8zrFwxtzcu4XP5lM6noZN5oOOV0xDt3W7nFLsnOEHDDtc93KAxuGat
UulpzwcWte3OZvnj4lNZUKZavvVVl5Cs7q1n3q8ijzfIo7/1Lr1F1ShjbnEXpU65
+iFEVW8lzBIP4xOBkSsgFFgjdQdPabSxyahgpXtjgl5wK1QKCocdwDjj+VCNgM6Q
kNyrkxviFlAp5ynfXkf2ZgjqZO5Abtzyp7IfC/5FusC572vZwKHiRra46Xdmux+V
Pkh6190F/8kM+/SPWT8UZi8h5FL9CoST/0ASY0uwr0UlSgUORZ9sIFu+o8x4ckex
ySKfby5gODGEPtaK3KLGG0d5dYMUZIyudZCiGhho0Y9/QP15e0Pv9wCx6AGpw1/M
jbUjqgLJ9zC2Rc9C95avKdGOVA5m2Id+JzvuaLO3mQtgBO+mvvrWf427suFSVZli
XzlcwOV700iHfRxdkU/jMG3X6iYk9YsH7PSCuKqa4SookLdXlb2pny9w8tnpMBYY
yggaCLDyM4D/NBLgDhfccN45yxj78i6r3pNaWGLYzOa51p5JmXm+wXmdMP9oKlnm
5a/4wQ5h4abxcs1bMSXc/BhuPjuZw3FdbXU1fd8zjK8MSYqCNJub7CWOGgQ/SweO
X8NEfLco4/vX8bpg6WtH11AB4mgFfDUzpGRudqemRpn/sJPgX0VcFer+Xm6rlQKT
oKCzqeDfuSsa8QRUTvXWiETT0HVbDhKEphYogJQ1ERMvRMbbdu8ZlJzF2Vlb1wrG
i6zv2xzwDB/UBW4qTjDEgt/CkNXYhEZqrYolVYO2f5Xv+TlwXMw4frpKfV8MEgkl
ojUKhE8xslvVHnp/GhEg80AUtam7IN4+MlOLovFrFtWfOvH1BIZ3/EiDnPgb2buL
AHb8UY1rqZ1IW2Tbq07nvjYPFVtv2SqvOYo0xIk3NBW3TRrrdJ7JEK0cJ1osURvY
ohajGUwmhXO/51Vyp6b+DsQE0jsPgXC7/CgGzkVcBTOAninDFrjwhBWOZddk6bUa
JfrvhlnWlPZiwGOAcDN0ZqW+y9fdg3MByuneFF2AUwEUUkeBWGSjBiCgmNxa5Uol
TBpl1sfESKhhL3y77G8AygUKND15I8RG2ue02Lb51LhSjiHJHZL0J9xI5c3kOTT8
Exs7w2lkGudnI4bDP9CPaMwI8d5ym/HVJOUe+srwMC5W9IEj9ZAkUdfihle7uK03
rLbNePktDDxr1jvNLGjx8ta9ZKYLL2XRBFS8dHpCM7v1mW6ZvHf0YEEJRhkLNFnI
5nr7aUEpipoDstoebrXI4FNa1t4qI+Pa5rKeJjoJTD/4UY0EkKxxHAgvgkTgcL09
4bgPI0klBxP+3FN8sT38VUyrYsGo2++aQimGppSL3YyFw3CIm2XFeUjSdp5DIW8H
KoZ4zqPjiMMCD2+l8LgmHW9ziDXxqrb//uxA9ELDxrafd3rjc1muWvzw+SdslYrq
OHVCL1wN9qWKAjyDewLV9DbSIeHufwrCPBV5DfB2mxthQCVXoIGGGIQ3uw1P58QQ
b1f/T3MsH5ZOiaL9rVGXIMfxOnqWIX+xlDVkmbyESNMitwzeNb0AAu0saD2AFIig
SFucMZBG3sw/CrhXCnc7AOdIYGaIvfHECqDpWzyDVHuxxSFlVjLskQIxLZqGn2J+
SNslu3l4/rCfmfivCURwOjpNktVH0B/kujenVz9/B1Bn0PV+1cEdauNhDjLiAkJn
BWB2y7BprdagNak5tKEt+qiyNw5SncUXNkBC0qZ3ZOmswt2QMPAe7IFWuCe3WreJ
UP4/Mo7N2PxyYQi+hrhWSvL6Bq/ceuf7tezkH7eP6PvmnTivqHvT72+TMKpkKczZ
OW3GQ/3tsJ/TQvgUkogP48AnlPr/80/Pm6wkxqOxaUQTJhqySDo5nUIAA+oanpSB
4OCkx6gC71+ucY6QEJAcLxTp5OX/kbC/4w4jdaz3+S5IfvtbxEc7pHRbRXFBDYo+
WGpKTn+8XihGY5P0SFF+fBxtlVhAr4JxPyaWx0cASb6d8CcK/VEayejGTUWf/Cd5
0eCNjsVKYuhPH3j3VvXkDwMLL5E7vvX9XWY+wC3sZDzjQpHthTg6SdWISVPHZUaO
GrIudHwfiMWa7Xo/Zc0zxkUPNdwz8FxtRyz68GIoLkD9/cECo0eD/lyXM1lWRYB2
z9WwpZIXBWbwjvKFYB9Ww59ikgsTaYQqRtKRR8F3tL1DBd8YeY7bH0sc106kk2B7
LhIOqwgRM9OfGE+q1KzZmD9RkKPfKWeMvKMIHpoAa8kddQnELN9ksn5qOYFYTPac
v2QhrZryB+vj1MJ5YUZyNE8zSeddrulCP6n9r99cxLoFJ0uvKpFKgbQsRTTgsEwb
uMiDACqU8UMxUltUHFtnOEbZwU3qXRdWRlh07zojMJLsFAU66RLaRYRwLwvCJcPn
czlwL8jkIzjA2DgtPSUF1S02LW/vv9PpnOandH+oiX0CvwLW8BRWkNg9uOChdw71
1os1kZ7AsidWho16xJ1w6fNOxkH6M5TJJtrQlRn7owyXmjjB8j3/mV1DhONMq3ge
FvzIfvlCa5pZA4J0tBFUyYsKYpAwyJQW6kRX4LmPWEK0FKuhEYW+Obaafff2JBh6
TPxsv/+Mb6VNFtbqD1++1klwVXHcbtRfd7c4IJm8n0xWBVJKYhFBTGB2vOCgnPEi
VGxiDEVGJwNxiVArKSQjNtdjoWAQweSgbleQRy01xa+GiQ7/FAG25Dpjw3S2b91d
ARpdZAR8xFy45xQhy/jJCQPlMH3S9StUatcEIkW9vjhQ4+k34a1fS1wx7vT1B7g3
aAvHcHWyyk9TGkyaEwAkNxabNhQqWiqK3HQdbiDrXus6Fly/WFz3IEl6a0DdOjfQ
2nHeslBLEKrU4T2H+VLpUUlRVKCMovLhWW123wmkeH3YarJs03FB88A0DfKJve4V
fjAhdqUSF+CdHiMhEgYGK7TmJ9WtzJh/0UUXda0QpqDRuxjj7xGZnTQtdGHHHuP5
HcMiUA5+orS+Pwq4xqcrVF1q9yB2R3DHhvuZLpjjLR8G+z9N5pe+elNBFX/CmQyA
GOAsM+JnIo6Ku/f2oDSGy1680vAyBjkP6XPYyWduGH3590R3pxef49R4mnc7UJGs
pknKc88K+cMr221pXgVm4Is3fDSmtnXhuxoHjhvolQ1hsfJ75ROEi4MSAOdWpHzL
5gjMNAYobW+f/O83hsYQ9gr9qz5Z6NnskZ6iOu1fICXruxLxXjj7W37MXPcO1kK+
pKhv93akmhyL1A140BI37biOPZhm9/5rFoIsX2wVMHnDi931FmQfFxuTpZIe/1D+
QSwKmUrsfE0OdsOIOYo51rbKDeJwIK1JkG9Q1x16NlvyqK8JCinryEBbNUxalTP6
v5fBTkgWoXDB442i10rdqOnZpRWDvRpEndIFMmGU6yHs89CM6VUmBFGs0hpwVJ7J
Coxi6eKHhPHFDaZHhOl6Zpf1AslRFQu38WHHE2NX8CT7Ds0umhCL/g/qwAQMbBuJ
pckuyzKrJ57WI8MyD+vccNPWbiVQJt9j9jKECVRQLFbW6MsU20fOg/jd8Oatb2DZ
5BqS0J3ryKAkJsLRSA4l09oJxmz/6mTznbuZi/rE2xppumvmNZCNqOp96nIVdjKH
BBI/fXAZ4I7fvBEcVWmyXLiaMpXaUfP51TbPWeH2oFuFqzIjOvJQnf0w9FXLnoID
Y3awTUHxxIDmERFGq1xMo7SHtRO5yL1OzC2A4QiPYxT+/uYRFFbLBs15WIvr9GqK
A2p8U214z7/OxiubcuNMdG2XdXTS9zy9E8kboBjPe7FI9Zr30NlIj9p7EWOs6tng
Muu5F0N7+HaFD/R4Kb+yH/9SAqb+DgVeqZNLWJmInezC8eUczRKR/ItufW11WK2R
NbpkAAb19Wn9tTcDYcvAh4jbHOjzW7edmqS+fnXLFDDKdX9CbXzhovnmPwiEw8nE
WXZGSkvVvmZmMMo3sbY60ipC9IbobJRbfa3uQNke/gpYYPwklZ1SzQtgM/Cf2PP3
hr5byGfhgmZ/1bkf6VesoN/bA0N+AtPTiYjugrvJ7OBh9oA8rCB3hcA4S4qPqV2R
4RiTyMMdGLGnRB07FLuWRepfMzB0Cgc8fsZZGI9tQYsIhGJ9hkqif2cmapeE6ckw
oQXrsJcFU3PxofVNMqVLwbFo9uObFF4MUely/0DpITmqdQAn3vR8bCZNJHwx4cma
whrlIKEfc+nlcwz77hZehrGSzZu7ootlAgLgbcdwzPmwNSMAEbqpS7bfmu1TcwCY
kZGjBAu1pP9yHGdm7HysQB7+u89VuXeCu+gbzUx2CJw3MYKINHksq1GW3nruSLzZ
CjVlK518nLUiw/1GVxiJd1ysMBbR9r4XX5FEnT3ov3d+TkJ7umO9Y32iufYuXbRG
2wUyPHP7Kuk/3IxwV7hdtfZQA0LHcbeLtnYTsWJTIXWzw4ODu3ejQw1sYDSJCKTs
c6X4gAy9SYkChUYcMfH58KBR8GLEd5yHqWej13qwxcI/oRdUEnyVhVtRXiXqgd8S
7PoSHfjjubeSPh286maSu3CkvtsGFyH/Cis48GFH5R18jGONlj1ZmHrIu7i5M8nx
2FWrReWzgbD8L8jIcYg3XA02xeP6oZ+uG6wkVOO629/u5CkUWiLNKrY1EFrGV1oT
HOKmU2S8UpdewJnQkaPU8NDcetuiQcvJUVI3nRHdvljD7xW5X6R4VGZeNffc+OTV
50k1PH5Ph2DQBPnTiMZ11hueYEWzW8vy/8z5pI9AFgrADLs8nh/8SLr0YBRCilqc
6jSzzDA0codsSYD1vLKAjcNp2mNwBu8Q9zrCSpyE2KVNudX3U5IXzw4dM3Ezx8FV
61XbqOMrySfgd4izkkgLZ/vBR1PsMmC7i9AkSXTLksUaR+Q2xFmRSzI1KR0/Z1eB
cv7UoaUatlw/2kVNm7KJzoMhK32VteGPDLXSwdwqJS3EKxV2kpK5S+0vxPJWBO+J
4VWCXyvkkZLMTF8QvPxMzusId0XdHpr/sraqVQE5MrKH2EKCeNMn/o/CB7cCHRNJ
fiwsQIEAseJxQU2BKFJQ3anYpDo5hquXS+/pcZ7UK5DTWunaBg5EQCi/2CqK5UZI
419SIAnV+9aXvHDqx426qDu9TSnZSzHe4N9c2GpKSjG3MGI/CXR2wl149n63NiOb
Y7TDsrjut4dGYKyeRVQejVRx5DEAV+/CK6lbFlw9xgw5JQJPUA4JbYThou4EpsIS
2bxcA3p26TjEO9/DlhojR2Qa6EQEaze47o3+nUJR7ajLkhyjSYx6qmmlbRe3PGl7
4gzepOU0y1DT2Id+mfuJQIiPRg6NxXhCZNXwHfdb20Y0C8YVEp/kEN3DqmanSk78
KexOMJmLqeGMlQuzXxUhs1TvbrWEe7fuB41XyeKdTU3Uem/s1JhGYnpQBfuz2Mfn
NkL8BA0LDZ696bc2TGHYlmakllBdfxJB/CErDwS715KYVw1Py+gIJJnz8DpgVpyI
/2c0CRFoqaeHOh/ETRqKZWNBfrSyFEuDJsO/hYg33zg493UqCVcSKYsfQ4xFZwW7
JcHYUNogX0pOV/V2OR1ghSPVJe5dET0OQqvmoKl1wVfKOhQzygu9k7MkE6a8Z29G
i8MKtanvEbhR13Lnp6OVizc7w6j3l39kweRsKReB8EDD4MFKkWUOYgFhUqK1JBOr
p5Ay01JU8hzM2s1xMrjV2RccQs/PdwQIyzA3b/mykB/i7OHbQt1uU2YTc9r3HaWs
uw6xH1zjjgT4Fw8WrNUNJouftVDdDb11OTWISZGNYo5+zyGm/LgqkVMmP3xHL812
g0PSyUaTJQayFQITwWpOmKuk5W7kGl1m/xq6DJBpZ04BP7n+6Y7T3o0gKoBhLGzm
VxNrYLaist8RTZp5X4hsq3zqkSyxAaS8RHHz+lT9pmDQpokh4wjg2atq3B9g7Gmi
aMn/deKVwDGnJeBnOE7NF24y+Wn7oqQ3+IYrmO1FBzgV1f4kKiTbIh5Vg31Zyl05
pfPzawMcdJR2aItqOM5D/bqJfo5SlEx96PRHQdqrfXejqEvp4ydd1OZv5PtHyP9v
UrOc3V2pP/yWJGdOiyhuWcbtEydKB8yD5vHDor8HSGN4FikSG178gSPUpFzRD79z
Bc2QcOw7sD1h6S9ualbpU7vFDct/GO0fw2IPwXzVnu1612n582JAdMhhQD9NnGoz
AlNFjVLCsddyzyut/T6s0WKQAKdbmWbR2Zr7wY8qT6KN6yo2vnC6hL1bkt2pCpZV
lfqDEGPWpk8sfs6ynI5/f3yAecSiamPY951fSxYwlm1eJThbCdOECLJVZe8pg7fd
1N7fbGD1I/WuMIPJNbWPS+pz6IOkANpH1dZj+RzysWqin2nPU8N3GsI2GcY/jGcJ
RTMTgW+dMCjVx43tG1Y7a2P+iu57D1yUmKoeymEbtHyxHyY+lDG/M2eG6LJtrg0p
tkuhlFJBM7IXCR9p4fgP62GsyDBCl8rkk9LW9QsiLA85LIbFafPUS7GVq/xVstPv
9ga6MG6yRBbJ+ALoShJLSY4pd30UhR4GI3xNWNbMtj2h6tXcZn1oBapinVMvkgN+
WXt6TpM7xXt6SdIx6/8JpQdcDzC7aoeNvBReg1EjbIVPe17dhj0aOp6g9gzfYdpQ
jIZE+o81UeWSMWLB/GxT4CsBOjee+HE7KIe49Sva0EWZbsPGaxS9nb+UCnkgQ28a
hSvH2QDiMIowqwuD18c28emAaDlzcqKBfaPwhPWIBdy5RyDZ7sf6TyTldivcLP1q
fkwR2Cb0jhKQnjxKH4iaSqjxWX8fOxST7gJdQGT1jhjX53h/TgaT5PTJomYEJryz
Q8WmlW42U/KqABQsPorkLTMPH9qLVD3f0lBfi4kyr4TR/xhU07JUiTU/8/8unaw5
TU8viO5kLYDFc/7+yJdvLqzM7N1ViO+uYJx7JF0s+REf+jE2iza8ZjhzGM5wRpj4
huDCi2wIHLm/ulqnAxl0mTPdoUMFrQRox6r7P1wI8wAphUp7IV3oisMNVU+T7/Il
o5h6Fz1FjBsbp9ZQgecmfZIlgX0SuHk4qtNwo9e0W3ncnQVJuGaL6ZmGb35/WuzL
3SdCpoHMEKCcXxhwK/FgJR2KCmxVcPj3JWEClJcm1V+6OBfVFJmeS2FrcaVaRTT2
VSmYkol6NB5qBo0LYLm3767mEeq3MFw9SDC87JrVpkGpHxahGYYXwZbGCCh1c+OY
cVJe176sewKAV5zO6cV9Ak+J9xxkuN35ycAu6PwJ+UsCrGL1PMorPQoJUJF5JA4M
5wQD6f0iUlHwUAj6MPXtK/WGvaUhkRmVbPDDj7ioK7ofyd9g85hMGRA4p4Sox050
+OkGkK9pp2m4EcpIMtqCjgK40foDhr5wrPEhHJfvftZ7PNOU4OETlbkoQverxvJC
5soJkyd7duZPFwPPPeUYONAqaiHHIuJna3biQkPVrsPB1d1pobhueP41BAkF3KFq
AZnwBcMGc7g33Eb5fGbVekaongbMh11/x4HjSjh1hPGEuCu4i3Iy+0k/yymDtuhD
dt81fwvXvJo8zwFAvHsae0jv82pMNqPZ/zkXYdvqHvwou8iaFnTyYtUHab+F/4EU
AOjZhJI1KTC17G+OnN58W0LP/FLZwapgg1y0S29wtwGYDlK5XrWRY+HfnFe7U5LF
lPCeQjCg6p3wDyeRdlXh4lhD3hVrOHv83CaVJwceS2t3wPm6Y5dVqnxdI6S7osWA
qJiMTjUNWsy1tBUtSNads4hSo+IcoW3jKq4pXypWQDI06OYjIJ41SqZitcavcH/W
Ym6TjAAKqwoI1cZwKv1Pi2ZUVoiTrJ8DkVtO1nuQNXQZhx8u85QaRlVhhA8HvCZh
BIY1wZ+ZWfDyeKd4LYU7p7nRsGFwKv/Qby+4liSD56+suU3exsL6wF9CJznuNz63
tsZ7j6sc5BHv102bSvhkpuz3gvHKO/EAckumX4+saHPrSZ/4S/0jNboUgCRgdHMp
HoQZ5qkJ+5ChZTMw2Vx70q4+L8BsvmDJq1V8uKe9DWgo4VpJkVf9cXBbf7KgRDvY
JJkPsgOGaR9iA4LefcPYBJe7zAvrg+kIauvhTqp1tJIItAY5vRQlq9ZUJ8tIDZOE
6n/+3lxotHyukbaaV0gdssi1Fb8SUxiuGfMSlXMG8V9AkBPN0fxLvcYQfLEt18x7
BE7bWEgaCcfE/Qqw5GoSHsGcG/+X6c8wkzwn/WUF0wMYNRs5UeNY3fN6L+SQj3jE
gf99MyPa43KAYx79n0ak46iF1fb6BoThmzGChkkthQCbEw/X/K6IbXLJSgs0DDwo
2VH4yIOY5bBTXFcNaMjs4HLNZEBwe2RvANinCfVDOFdd5F7MyxF+niqcnR5nnVW6
t/91IctTqUi6PWKCnLf8IlBYrEtMqVnlKQcNGq7LETR6/dVCCOTECiTQUENPHHwz
YWY45W5Giagm9BorbVnPT7WWbzNxYAFx6DnGX7qa0T8Fz//v/vg6FdYvlcHlbC8k
6thBx1udo+BuSOi/KAdw96QPzxo4kX41EjVTyiB2iYgVw+KngBPV0ODL2ujUv6xz
w9LKiEyx2OXU1Zt7j6NTnoLPyYVy1FjbgaWR59Xv06z+7umTvDubMWSGv2w8UCpd
zcZFzpzEAlilqI4rTLLD3JGmv523WtxDCTHk7Tl55NFpll79oQpA89tNYJFMhI7J
vcBUzG4vEg4OpsLeqVw41wV9PMFJGKsiSZBbTO5/FWzuAi5cQaH6qAthn560bEvX
1yGIQtCOkfoKSQHBOhRk3qX4YyNQMUrZhUFOyRE7l+g44UnVcHVVp/jl70Ha6xQL
VW2xmQqyhNZybg8ARd/237lrhbgoUMTt6qoUiTJka6gu2gZmGQ0k3qvWzw6l+THB
2bVtr7C3K8/8ztgzJZFuYHc5HVjPkGCpVeRWfYKGzH6nYGCiJUd9tbnc3M2VNggV
FVDwacfUiD/4lIejE3i1MhCXu4MF9GXioyIz6xNRyF8Omz4Loy3ZBlhEAO5ro1h7
lzArqTwOTvu0I5JXlvo8GgY6Fp3OcUXF7BAplVHY9zcNQT65Scgm8A1F20P0Iuri
tpymWgbne3TrAGhM7wbHjPgHrUss46u9TQ7c6Ldr9c+DtTeD5aOzyRobqRescaPH
y/+SrYyTNAvGNxK9oVmv6Ia+9BMHMCGNxEW4ck2E8i9EYoZH/EgT+DGL0Z0daY0t
6wU5+wc1cDnNxS/S3PuP/b9v5Cx6Jf3hXqOZcWuI6rDoxE5EbIIfC9iy0J3V/Zm7
41PsCs8NSxhL0p8ZYSuhbvW0jFjp3AGrigZFdvkZRRZQTiEAU4eiXRUtsNgjU/ni
eZ6FgKKdf4jxeBpNK9Ca5fLbaRthuP1amQZ+AVaQcHB3ahCO/66CDAg+XT7DK2rb
cBAWyUBfcNryUSsIdbhTBl1bXskiLD9QoMHJhPIS+b0JC7p6V5r4LBxm7cnQ6QdU
VuSOZnJWXq0bZ4d5qjKX+NXx0nyAN73JK6+CxMZy53W1oMEe/2Vpg/COrHvILsM0
SdbJoseTy08F+vtlf0LEJfYcjq2a+4qMRCISaeNdIEcqL7cdtfmwIyyfR3FiWcP9
8groWcCUYfoa4VrAX1ENgSyEVzzBfIqgIuDmAFPQLpTRZSZkyWxJFIxIiN24FddN
I631rGtuitQyqequATkHnZyb7mzW3rd5GPBiwuyUuH83mAnU5nMCy0nZmuwwAbaW
8qmQ4VrXG9Uznkn0Uw+9JfPoRFy02sUU4aKJCC/gKCUuOZ5L02hPKwsdSuPyBBZ4
SsNtzxOUsvvg3j2pJZqcvhl9VcxisbE9eRY8fywhl/S5yMjxarj104k0l54IbHZw
OIbznurDzjmSaYtuPlgqwxpxJPtfySI+TXGbPr7dTKckQqTtMetpHSzFCbT8tTJh
woQADJe9b9MdVqFiBnVVnC82PGGzkeZ7e15TRszyiScUPYTQjrCwD/Uxxn/EIZcJ
gpzeVqhFe0ETaqq8yjQ0JgL8FMgHnMVqkYyg72wT7gMaXWogSiIzWleg6SgkCZhp
O/m4RiVzUEvemx8kAGEImmowpjtYZ3c08YOSxC6U+jn+xzseooyCcwmNM+CEtASw
cJCwVUlo+n2yc0+qvX+H3tYEr+oWOEzTElzcHHORqL2GHWCasa07ghzsx+TAT++n
3GQD9n0NTvgRJZg//o/oGPDcRj6MnS9N8X3lYltp7DRY4FhZuYd6SAPfm4WjGjjX
fPixJ941jUXEhXwIjO1gA1NCEzQZgAF8RZc5rd+TBa3aqPkG1vkBaBp/acd6UChU
eCDduEZHbyVbD39VyPTv5H1L4N/BVUM3/I6O2KF9gi/BZPNq+asgapTvgm8WSLv3
7Nuh8o58MsR6O/BtQWhqAYVv35EPben5BRXwupszjwnPzFAXAo9g72xAB+lFy0JE
SyZB5Eb+np36BYr9bJVRPCZI7J+eGxPnPt2AfKEdMbtZoaTx5sN2g9Q9z9sma737
LsHAgvQaHPZ9C7vWBheG28KS1Q7liM41ShQqWk6WnvBPbTfbi3rte7/lnbQZySg4
WFK0gaz+6DVpeAy+UktfdK/XtiIkTSjBVVAlKQQ1wBs9D1+FI9tdOmdccgRHhZUI
6e5VuL0I71x2M0N0c+gChED/Ox7bBUImQAjN26+FXvl8ljN5WGeHYAtCuTeSZ23d
9/LxhedzrvuAZuIXAiQmi6vJ2xQJijVMzlqkshAD2hYhitX3iN7rPrBwGx4dWbxa
6kEIqehkcJ0IfwcPFxnr3DXEHYUM9Pqp/eZLU7y97UxM6zXopmvnM5V0zsbFhs9O
+3WwEtObdNkszuM/t/ROEYYva5WCJCRbkbpcMr0wXFA8Cu7BINT4bfhJnq36NRRH
tw6EoTXAs+qf+HF21U7M8dYcyEl/JUckN7zqWRPZ2+MKRom4Ms+jhv37glMWWkA9
jY1G/vH3kaFLrvjPQAZXbKvRQBOywHjCZHIAkCpMtq596clz1fetNdCafdhW/GnG
OURMXedO9vKu3DD2RR8cBaNJF0LQUfFSH1GWJ14qLoy2R7KQxRtUUjv5YhdOQYnf
Ws7nPK6BPE0U08nTX8PfCMHV3+Bc7J2xjyniAYymws2idFws5bj9Jx1PFjSIONNE
tsb7b/YV9vKW+e5dLVZBs04F+XuF3ZcQNTHJxKRyjwB9FE8ZrEY2tfU8vrB1X8dl
QLG2kL0rsUAXmH8iJE4wXeG6fRSEOR2qRU3K4oORxJRzGTPK+KXnAb9bS2tX/Hsx
yNcIDkUv2SPwIM9s77DTUkpHu+WW4c1k1vaq8AG5wi0jN2ZwbuG2E/nfHio0qr/j
0+GBb+cPdHzj2Xf6d9gGdM4r1vvveToO9SBvj5zJM8qUAjxr48QgfqygO614iWn4
2MrXG8fUpKQe7lZeark7m423KxZNMb1uI3x8dk1Yl2n5EexManllwBvQhT8SUW3E
yhOfQyjdsAGvsn/5TRtTAaSKwVEO/X0FYxVK05ix54FsjOPNSFJeF7wpTcR2gbYh
hXAP1atlps4zr6vfpJ2uqdurjk+Rcy2/O7z9qVy0u8VA2JC+2i5UXiRAptdMQFlL
w35kS9fcWB93Az7J+ivxSa2Xl3v8v51GLFfK5HmA6Gb6CEfN0Ypd7SiAfJRZ8J8R
epWw5Ffe2P8qYP/jTmjsEAR2JEQCGAx4xqtx0fBgBse9v+sbvCOT1+TxzQLQJaVn
kN9FHWY5bVvTDCKCqB1Qi+ofHrRAfIh75d8XS8GMjRJC/94z0ESYOTx5UOPa24lF
KewMFxMZnQU/GexEo21vW8gs5k8s5AMe0OQtD40QeZmIIEHj2JGKHDCD4lKTxol+
n7NapW7HhQO4nDZv4KSU0pWQU+0HXOxObvLKRff5se6ZH8GseGmmpf3Ra7eKMUUI
pVQQTmQafgmGrYbTm66+kuqu74YbNpcltrF/L92QFzJl0ehfWWytzFHO4NscR1WJ
v6qpb3q45LuEdqihuRBfu0bszVOLRo4q301l1eyvIJZ9nzUhCHxwxsDUxVgGdKSb
/AVAUpUzze7CYsQrzJnt+rOghp/ChF3OZxGYRWCNuMPb4p0xuNIr3ogiJm2pawaS
8NTnKlpx5LyN3y5iDA524EuFTmVQrWUzs8CdBNVWzDhZ84mdYpjYfZHJ3FCy/BoE
czSLOT39Rk/A/VtE04JcMR8JDuCPGt4/qn85ug3E19gQfDBb249leXc+SzyPOMFI
oar1HxuxaUm44tZKJQR6cL60x6r+HzErBsK/fdWLEvEua4IECQ/BpP8CPA1freZE
2m59zNWLVRBxeOLxvODj7JGO8NfL3UbLrYRAn8W4rU9SvoiRa6IomaFi3LDnZ8rY
Tw/z4881gVU6PyqKf/gqzoC7Cu4FlRQjoatFu+eZeRbO6bR10vBhFi3Ko9ka81u4
6jb2qQIz4JLZp1kH8dU5mbz1P6AKK0hmna6gukn2SwpZthunBXvJ8gkCshODpn/w
gTPh9pyxlwC7RcGLNj3hqaDqugTMs21AAQSV0RXsXZaG5p6px76223kAbb8mfn6G
Kco2KigNgPb3UtA7ox44MDIPMxagynUuYJ98c7YYBxh0BLQfohZseg91W0jRiFCY
5WGYOc1fR32vsgD40pR14hYzNM2avaJENNzVJc99vEsSescMi2uq1H/JfaCceXQ9
21q4u7zabRxJnOeufUWmMYXZh53vKE4j4QNcLfezNnLFsouh4EGYAds5yHbPDhWZ
P3WBnzHJWMUeNvqLM7eezvFtuE59l68If+184Sb9+w37RzD+C4pbnH2vfQ7VzNyD
5+uE+XyhcScAhZ0YCWM5Lm0THWZpojZMETGgAvgtHQLv2xKLT0QsCrO4xdBttYOd
ROUKbYFOS0mfTZmBMprTOz61z01RGt+T1FZMT315ZrNLuCWHA0O4t54WK9keUKHn
ScqJuuNlzJN39eBkTGcGyx9LAmNHmvqBbG56Mx6usBMItP5GnGrbzZ/cevOAzVQg
kLjKuap+n0yji/PbhtJ1HiXjCwrSE8kxVrqUcvy8uDikEmQv7c5U+NBTk/CL6NMw
o/FgL6ypKQn9jNHCNnje08b8RmHIufS8eKCfhMABMlWfnaQXQW5edKmmcZnAsxeY
d+JCsWwnpOpnHQSohsbhOiJOp/ywQjZ1ZV5l1jnkcBvr2uHa3lRktYiHG28x8kP9
vieyFsXYn7dCQ6b0MlvF1ouFey2QBK+VQr6auYS2MY+ChEFu1O4PkLldnf8txRJY
NhHbxkbx/Fj4wcHytHu2MiHWDNeTZWEUZvmWAb28WOjITpDM4+BP3+MVzVghm+zE
OMj3PchU7rZ8qr85XaysD52/UWtxE0Yf3FPFWzssFC9uQuPVxVjwe5iPFu6ufz3D
izvdzNDWwtSxAg5jCFKbS2JuAEgA1FywUGI6UMpMWIlWm0mH2iGSXIU2s9WWPCXt
tMlys9uUJKRMvQGZZmFu4ockIflXkokBijG7XdERPRziP/tR9GnH1ebTb3Ci2sGx
rHMSAak+omjFC6pkkHiuYO4AeawCSWjtrA1btDTR1WWFKhHdxDzhVhIA2nm91685
C1tSGnCpQfvLRf0oy3eTvrpyf2GQdNfQ+RrWXq2JYbQi8gUSwQpZCvXDCEOxHwoi
i/VFWYQOuJrhznCuK/zHLRNMi/tGfHsjBjklAW2qDBOPyjpisZmIUJ9GkVHyUA90
Jxgk2Y32+ucqXXusss0P/ZnQ+sL4lZzT9E7+EZ7e+cObg8zZbgJl1RmfFkVs6ObO
uoPJbGfgMRufBA5I66AQsvjKoAnRig2uC9ddl7KcMoWPktbbnYUKP5v4FyPmP7dS
QEiLbx6pBvPAiY9IYTErNQ==
`pragma protect end_protected
