// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
WCNZy7sj8zMEBgqnCD3sHWAyVAQa68A1DI3fBsEULjYpl3gC+qymxIhddhOj5y3x
zrnBFvlPEewitlUwEJf3CCcHpya9FpioEMSvNaXPUeXbOkttIO4kC1PUz7P7nw8l
8MhuwfGJeRN9MU+HHWPxNQ/QOBr/RrbL8pORSqr8JSk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 21936 )
`pragma protect data_block
MBifc9SKcM/aSbVc4koEflSyl0F7UBz6PiWIj0gjzxV5jkMJTvY/eNO14HKsRnUR
K79Wv8M3Wqdj4rAuX2+LjviZfEuRuNtXv/CYbu+sRgDSnOnSyWoNI94UJQ9FcjvG
nCNR+gFlBStgFSq4ndWY2GVQvfLt/aI2CvLmCmqTwmXzh+n6jRBwDkmDwvN0cZtt
lzg4a3pWYiky1qMfEXRqj25xEPFSxSHMwQAbiaBmMOTo3WzHtJK6aeFUQeE4J23t
Rx4I9k+Y3f+wb22L0PQo170Aw9q87Po2bh8dQ1ntGHcPYCFePoplX2sx8NuDXdPi
exD+PTJvY/DGgvD5wySvfc8IdP6u7nMuhaC3Vvk78hNZUb6a1Z9JnDnL2iULghg8
kAUVkZYaV5je8cJg6CNG7jX/E6BVDXrNENlkJ862R0FRD5XwivE8vQux5qdPegkH
MyPXmNlAi9Ur4i+Za6cjB2bK/g6c1432SbMAwpxv5bqOyWuquVEnMU7EAGgtGqvX
aQNm1LVvonGtlxPyd7i6JR87lICyS6XNmS5KGPM2qya9n4ThHyeSZIvcXP6LmfPW
5BEBBkV74RmeJjUJTjgfPR+U+joyBXjtoPxNTSOZOasPaJpx5ACXRLCbzHGeS0Co
vj0zmC+RGyL7+xTM5qedsdF6g+A2c/iAcUj59WjWy+Iyi+52y/SBNF7WiWHIlTjC
37AVANizKP0O7sUjtrlZI15CNsrfWtqmRpEBkVig64Em9N3b6SQEztnMTGCrhrrV
qlZekAQO0RYSYVXOSnzv3LELN0PzTX0lebiCuMDiFTX7nLJqYU1NivlwC5Mz8hgD
hgcv/NfbCGlCsRdQGvTmpWnnbV4oR67hFwa1EpF0bJb6IPCDoyQJW9IhWJ9MujCw
iBJSSemloaSjuNSmqYxTukTUDujrileN+LCOW6fVUZPOYEn1zkhAeePWh0RSfuGw
wqitTUaXWBDwCx3ZNASrD+7ZPkonLTrkBJet3ycda0HxVCDihSCqaY22bjDq0rq2
NxG8kd2qcNDOaaqFTDnsl4QBm74wDW421Md/LACbRs4632oNuonZ/R7YKTe5L+ox
hlzeitvcF751fVRrQODU66pvjTv7rfwGx3ubESSh489vmtGqodMX9DNBOxrWGERk
FSsH6RwVttPFHFUvlxtXoKq/ipcCmCHap2nj++0Omc8pvUuEJxrUnYGXi0FPPdyZ
648YRHMUvyppszHq5VPEOTWDPZK3A3ZuFgo/wbadtl7pRC15Lf28uAY9DGVXe9+3
t3KCmXYNA87x+/R3UNROoI5R2XAOEhPJERBKGEUGZiriQ2Fnf+dm3+KMFvT2EW3K
kmMtBFr1+2acHUnV9ZY8jfxAniYkYgz4qUiqLoVmppEtTWL3ymd68IcBWCBNRO7L
jGdEn0S2ErCvnmUs9bKWFDaj9GJEysMY8WThRcd8mx/dRMgWorhvQz9Q030eDoQy
ez9npDEveQ2nmLx4UPvgaAf+EHxvWQUScjI4AhrOIffqwKlYP7KXNa4C8rpaPWLX
gfT9KMZ7mhsFitdeh1jm1dyHSAcExx0dCm9ITDSVBwDstJ5bN3kf66FvZjTqnPTv
9qPklU1kX7tbbkfaZUGZ/b5Huop6ZaDuG1BgLfL5XUYr7HFq2sMWbOnzO7uDe0uP
qYYZNUlzpvbib4bmEwN4fDcTRiqKSy0iwO88OOvWGVAlUif8lTZ7pAizRVHsabun
xcYX51KL90miw+9PV35Pne8xCwoU/GXCMHPK9Od0/sn3lEhSkd2pGRxX4yLXEBUZ
PH97rbaDBidMmy0DuRpbuQtmgg9u/rUv4ZDz/6SbwvdZ3oFPr9lfqXSHcNi6i2OP
t1I5aoIttfloQljvmKYJP6UyWrbHYuqPMFQ4V3d8QKTNETFLMqnf9a+M+qQPAHxQ
JnQMTlvbPoM84LbB4ncDF4oW19XuvsaQ/XfoWKsnspnhzBcrdLijMcqhDMIVEFVS
A34V+/heWTmcXwzwR4eltZoiEhLJ4LUegiAy4OC8qjK1bQC07yrrFYy/V1V6Dsiv
K3NvmTCc+M38RaA4fpG6P0JzS5DkifLI4sLApDGs+jJy4GkTPXmj/i08dil9TuIP
EFxFdEmKIFIyDTqsYghwRQxYwnpElow3T4ksKVKIXZlZS3ug4ICk8+f3hR3ApBkH
nBW0fs+iuMmYvlobcWscFXsC4Y3BOJFGPwlCsIOAxROp0F1Eo4+dFyvESOTWpdPo
tiwSaPsGh7rdDO3Q9tuXFm8o25mkZAEzmG2tGhoGmw3IMc3UHvi0x4lX2l9VexS/
EyYujOmvw2be8TsV+nID6hIevGzYHTMw8W4afJkCK3v78vMd+vVnlupyxoOp0DYr
kOEwp5N5EqGzCNHj5T4wBkT9dn0YuLHOwlemI32BwamVdnBuBsQX4ke67zDV18+9
Bp2GoqaeDI3cQIGPZFIabhMjjrWyjHHS/9VM1L3pO2lwFGeX8MhTrGqDa1ZUlTVx
Ix/s1vJUZohv+D8Rz8SIxYHQzim+xZgFZ00lkeESrooVECImgbeMBkbaH9LdUFjt
UpkKE2gM2/ct2Z0WeN5YrtKl4Bt2WFcvMDtjzFXvKKbYqC4BaQcdpDG7YTkQkbUf
8kHQQamAZA63n3uXaGr2oVsk1ucbU2Lqg02ZI5wpByCl8np9u672HgpH6+IeEnD9
9n++aVeDCaSVkTJg+V4it5kRam0CDHBH1FztlbIjeXMVGrGVOOqWyCZyk6ANfl6D
c9q3mkx5MJKwV7jUn72jXB84bP+N1exdhbL8QOo/RZE/9yLlFs5tG6dgnIhkL3by
Ivd9sk1Gm70yZxxh42yFCmo0fElo3njZtrrycrJVeRoCLmVaOQIHaypvPCnfUKtj
i0ORT8Qy02nVAiAIppUVYNSntEVsXofUjbWzaAMSUyWyeRRwTWOTlLTYcLbA5WH4
uewAB1TlDJ1YCyrZItqea/5fYVRfA4ItjolbUeOp7Jljc8k0rkdVdTPYxNfHMtzx
YdCn+Vn9T+QvRN5IeO8ayMJpOjQX7nZv0fRJHVHtLqcUGXKebvTkFuW+fQk+xD3X
ug86gyQ13QOQIiozy7gzuSoa5sQ+C/+kCK6SQehwSLSH5+RfkQ+qrXcG/Qw02qCk
0wnLnlYpYQT4ZSUUWJF+A/5nvEbd3hSkX8QRLA7p/feCVad/kDR0dHyM+f3sXVej
2DGwb+pRB5MYP1UXgMKe6v8qr+XQEbV4joLcJEWtvKeW9fOrNv2/teoNazhjhwlu
YvSLAJAORsmqqYG0iIlfagKzxFNmG/dSRGKp+PqL8CuttHgTstJEZ80QnHFrgE1a
bJl+8ydjm1eO8jR9mgj0O7vSnHujpmhPDq2wmDuSpnmm51kO3vOXE9UygcIV/PDM
ck4wCTZDz4xjr/Pd3VrjYTkPnDo/C8EBW2b/8jklZiCO1DAVs9Rg2vpTw3KzeQxL
0SaQNdn1I0IOEOYSTz2BC496g4Uk3mNNxJLHRMYaQ5+yXqRSfMu/V+v9hvE98CKc
sec/KkmoxwkAQEtMZNd78Du21ZF29WgpRg3EEUjltEBbkpJIoc6jU6zC5vP4n8jN
BTCYh1Tpr1qFn005O1E9TSVLQS2m7Bz4PBtViNLTd5FjtO4NjYhMiAhDM3ADwKwY
sTmpb329qexpT63SgF24vjEBPYQ+vonguUUFIRITtnNWePD2poUdddkBm0MFSA1M
vcc6KxvynoIe/T00HECkMw3Tmg0ZIW3XtOgZKX6YemIMhn1rI1y93FW70gX4JOl4
puBntJmnxEwkCstg61cGxmz4bQAwe3qtZd+Zd6BBTwfEOD4X/FEVRUNJNCU3HX6+
Z1HmFqVAjL6QZ97jxpKxb70efBfKtednJ+A2TSIQ12xQZ/l4i4ccqU/9BcsJrNxB
h9y5tpvJku8FTAxbDmXNspsSTiM132+9W1F10jwSaHFcWg4srkvYspdJeRbRMABk
FDIgSvTmWIH8sunzVGrCndjJcVUAHnAvvVrKh74ZUoZXLEKybQcRwf+a3xup8y2f
AZSSHW55UH3a3ddfVSNPwF1zqRrmyLqWAFfj+sXxPciPkk3pNjMOGIPiRBISHcmr
kJ9vP0VRbfBVDmrrcFdDlP+p+/f7dId2cxomZXKSVbfvKHF/aYbbzuZekb7XlWd4
sGBuX7uLrtNoqgA0rOBhoizDauTJYecmCsgEsSlS8jXH7WKTXIppJDNe0ccX8EMQ
LPw1x5vZwFP7pIHVJox7cpOAPRA0oY/8YrR5yH2M4UyYYVJlBPtWvVvWFoJ585AD
1n1jX7XYB9gT5aGVHRPQoFAVepP127QKopRij29u4Unh/6g9VVUxmz0fimVaNNjz
+DptkxZ/F9rF7cBX7kLZ2j32CCwTpca4ehGsjdXafNcnGNfldk8yAbOe56tAW4u5
fuBAffWjhcRdY2ztKLmtHIhhTRGMYosaV+tgfzuyTezSdZcUxPcZ+5sppE8eE7te
xxHoXm1o/31fIUkWAh0cTDX+KetLagRyoBNPxpccDlAlCUoJXK6mXVVjHA7DBDk1
teWw7ilCizhbkHRwQehJPZp1i/ll3ZzPOB5Ol75FWDdj3rfCqS4mgzFwdVZF8TzK
ST78RBQEExN2VMk8/ZcSnGWD+3rsFR5RDaTgo5r0oVeWWr6ZRZLxYBjed5s8hQia
0e8tuQ9kuJxUlEq6819uPNI08uGsTxtE2Xl6Qv+8NcZqHNpJz2VRTH4k88i0DliW
Bp7oEMWNagxFeXr5/BE2LzdZcvP2M15IcokOjXaZi49Tgb5msvjl+fePPDnrxfRw
NK5dxjma+r9JiYE3AIqDn0Pmy3kvKYnrfOSinB8HdStOwK14F3aZQtjXSqtp+27I
98nWeI6gzU6DMu4vyaLJbVgIp5LuuQVdG9Pjfu0cxE/5dPWK25H8PLO9ZBDhcaQl
OpJxAE5Ik/YuHs31VzCeUYEZE4R+PFZgM+1i/gj8DR6RQgTIsdnHChk3LPFE3120
nS92aaQtpvU4SmXl3iSw4ntNszcXq27aELaYAnDONlpo1CHVNo1HldQxdXGFhnh1
HsROkF4R+LYAsJYE/eEyzOteeRdf7F12uaPV78gPQqe6EH7lSFvBBQ1G2Xi4M0VE
rVK54aT+oY7xcFLtk7aMgGsLe6jg7trLr3QuZ2wPmqs8QlkkJeTxFU5ehTcLTTEC
dchOY19w+6Yq2mnfXD1GfO/hbb+5jSr48rcx7Xspkc/NmwUjjAvoj6avp2BuOn1D
GehWcZMmFB/drWo1zvcKURw74/jN/WpSdBPypuFJ96RNXYDoHSUCsqG711Aonj3S
x5CG1HD6Pv3IfZzD4osYyj9CBP/pFpLPXYrMbLfM63JPfYl4eoq7oK165fQP4y73
jnWuIu4W7bOyDaR15GSLvUACzhXXEhQSgy+eG7lm9h7BRQzLu4aWFNcCMrKf9gHi
QQIZqS5Cv1V6OvSZF+ca9rzVYBhantLAFV9kP5KXYnGxSWwvUF0yRkAtmwNpA4wW
AtUoDHlqYTZ0/fpYlUK2gCdazuWoea4QCzI5bl+k+rbledR4Ycr9aDhKyHYe8I5m
oCmaLDlf1YRw7vRmdMq1kKN08ZEfKORh59AfIi4GfEHCH3juoy2h///mkomS5j/Y
f4uvDDwUxINf5CreaVt+G3Chv7VFGCnJCl33CD+crfbpcWCBvBMswdr9uqc1opLv
iz1R5ILWaHaDdXSXvbv7kDBMtgdGVdm/jvaCY0qxURzhb9WKAUMANsxlVD5bjcCo
iaYLhwaXaV6aBWwG3czZ6NvXbk/Y1/56AvtFuKGnsg8lwW6xsawkI4fp5pU+GKXu
L2qO/q/roDAhfI2byI8MviiE11oSBOKAPCP9Cky/hCDAJtWHNlC4ISWnlmwCHRWO
U3dzzm5vGF6TflcnU9pdk02QfyPFxTCxNBQyzwdO+vhVl6k8jnGvcC+Pdmp/oHTF
0zHnMJ8weerUWFTv6Gz3b58s9A2FcVtqvD11nuIxZfCXbesnx0NynSRq2OJ2gAmM
tvW3aTn/tcOEpO0KCvN3G7fNs/tqLfGvYSyiW/pLcCS4QBcFJyAcwvLjq5o4Ez1X
AKNi23Rz7L7F4o4Fh73fFrau6uqyntuxsg5QtentTxFPgFdV/okqI8l6BBy1PwXq
Vo0lnZEmSrwXrxX/h9y5iY2vESCUaPRwJv5BoLL5g4qEeR3TOOIMBEnSD+jNdOlo
dMSJZXanxY/tCJAMWyWS55+HxjEO+wKdBtz7pAaPbyW+kpP8+GpQMVB2sFtvjRt9
2Y6yf5Zj9rouW8PEzF5rX+LFWEhbsOhWb/yLlbC8k4K6WZa3HZRvZQueQ6Pt3W6s
TP5yRfByA4EM80LpHYUPTlLHUkTdKn9YpswwBhaoGI1fdqkAf7ftpqrlUNF+4I22
ih9QjEYgPCb1gqCYiOfQqHY+xlrQJtW9UuvOkWznyN3GjWySIHf4ncYhjb2QhkJP
BTzU4/8LCkVGyf5vvSiLj3x7IL5Q8n8arMymFsZBMudTgDuXn1zi062slHCVSF8Y
Mw27yiO6Bp+7o9Om9leXgbdRLW1TDtifJE7QRMZKXkYEbFp6vzDm5JCspRigWtRd
6TnRUGbYsSSZmcEmlKY41oo5ZKjMMMk6S8FzXs4yefpqEztCgXMECI+2vMluM9xt
0JdVkYq58m9Bqt9fMKpT8zbZYWE7yiY35n4IKKtgt6ThKndX8tKOmYD7Apj45Ib4
KLYT5bg3WCKkzCMbZe//OqgIoTv2CIq3W8PSwmCVhTbxAe6smvVhwuNBV4LTmjCj
GOu+RfhZQHA/e0WieUO4SIoij1mQ+HRU1BDoVGwAtudunGDsL2mvTg0atRsWgSvv
oBXoHXjf7V+L5c8hoxosrUCnz8IZ8ICdfpHvHvQ3/puI3CMF1ChjNIWq7J/Bqo54
lvs6spBhyzsbm4uksiLJZd2DPtyulTDbDHdQc9MY1HkXa58j5E3DogkR4Grvnjzb
9cMKvyxUZEBIz/9zodvwA5AQdThypAmIllY+0Pw8J6JEWkeD71hTD9lJ4GB36V2D
nDBr1acTYMw0DIUenYTLOENcNwGtTYyni/rzzLPmJUoxCHQxhDWvglr7tvuXCuap
Zwt1nhRESOmXu5J5qvG/FkYDpCL74rRx9OhRqMHwfnbDMduw/Gntq/q2axpluMCf
a9J+bfKOgnBr2E8WcSGwD7+C9+EAOBCkY0qp5Z9M3T7TtHB016Ow0ypX0z3fSQ8G
eyIdOZnszf8OR/u6nlD0uWvN1fg4oFeS6DJyNZjwEbevK3FjUnqYDQpGwLxiocHt
0SxE4MtLcG4weIcDibkxidt/JwjQj4eKSD0Cl657AHzZtPR4z8GwwOZmvA+xpcoA
gQZfqurG245WJWVhxmVN14ygeuJ1jSTJCJZ7tgBsypuneXo14uVGY3ES26HX0p4o
CMs8NVJ1B+HjrOs/w5q/mu7+jWySDYYf/sw2kQJKTdCiGJVFovLFH3Y3QmBV3U5A
4m+mlzDpDKJ+ymLqmlwo0Uo/6mLb06vfBiBRgnP45//sgvaxJ3oaGKoomRgSixqb
662UILv6IBVWiW7fmDzDNig4jO3Tdsb4aqHGHW6CwiokMOZAF6tTu3lR9OgwXrXN
XUqIh754dNkiUZCfVwK7ubRwSwJzHcAPfX84Tku/v2u+5hQ8N6A8M3vo+vvUqp2m
99puSfvvPG0HSHgC2oK4gppSJdLPTt1TVQi+NEuAPO2pnOiByrrPJNqwezflsYDt
J9tGikKQLgY7dRhJ5Ig4Hni06CI8R0NPtLq+bMt5N0ASSsd3eveQQEYhLfKfLdVx
6xexM2LcGMMdKwvkNs66c2BIRS2cV4XHiHriUcfhUvgi5a1Kv60PoXRN51YcSp9O
6pje69S7D/UMAKll0ZE2yaW5yOUoAPM9L7Gz7R+qYblKEsKsGHP7hhg2N4+94H9L
61D2Ryvi4Q67aOtCX4SiMlQOL3LnMsSIVYXw1EGFhKcV44EVB+5h8AinR22KClkv
/YjZNlgdyYwbX4VCmkhMwTkvQFu4LHJCxTyghQITEJCAhx9Ud0BRcYfaFt12yEl+
SGQ5tAvyuPG24U0K4KoZaRWEiEMe0qaB1Cm6QilUHPJKHBTD4UTfPWNZIItDlPVa
bdzB0TGFno1LjdRKGgX08UU0Pb24C/w3SuShMCTgV2Ef0qb2uZbaQTgnQ8LuD0zh
onX2hKuDlKEUyk9IeCd0JrU9/kkYWCN5xOJsfB0MhQrsNfguksHIL1uaAizHpnhO
Rl6yVIeyVpbRRkPMTy6WGJehzcBXMRKE/43eztvm1oYm9XhaicJ/wk9a7bwsWZwo
JqBqRdsO82b/gl9A0gOD3oZzh7DPs1zZ04KdaAvwcIezWCoLhgo93NU0GqAXOyIK
2DupD9WmF5CWcYOmfzDksxNWS3MWDSrMOkQ2lGOWkOG3Wf3VvrMep1VbCw9RMoI8
9K3IbUqCqrLGgPc9Ylo7hw/auE1+IQ3M4AXR1bKDKxkNUkB6VgDw30McdH/oivNN
lDh/7+IPMmfpX5MSFa1eIE+nZqatjHt+Ig4vwMtc2Froj57ki0sRVemRGPsfUiOx
4BZQA6I+RX+w9V7bKwKcTVECq4yPR5QozUWnvgPfFo/P0yW1g0mlyerBb2Kp7aIb
shCIyV0W+GU8XJ8gIS4f6cSSQz4Lyc4CaO1ALUStTcSa9JVjrFtREGCsKIO8W4N6
gBMdTtumeBEIMk9qumVc4Ll3wTLjBZPn6RYqkIrlQWRN0EXIot1mmfVfrWgeThGP
mjY03NjRJ6/qw4NFHXi+B7iw2WXkn7wMTzhx4ZKJdvyIHhdd2/IiyOHYQxUQOv7s
xYAFDhuxW7ZzqltnGERYiEBUvzbKvZcxn3rJ0dBA0cug+9FdSpqARansM7xiQE3O
XrCpnKFy2oWEmYeKlS7Z6i6WBF5YejEGu4r4cU38SLX2kiRvYv2oIHv1yih6WfUa
VGNDRi+zAv3DKPxp972B4th7O38qEJHRGHx2/P1IGETswZfy/mq2+f5vlGTGazWr
fcVPLc5r2+/m/Vb8T2AQ9TekJY2j2qvFVsHtxDJkJRqqyqnNu+CmTd2kYwR2t/F7
Qxr/3RKWejR9iue/RBWughyZx/rlcuehCCWHZ6t6MnlnI8jjrSCAaYwxcEM96Vz4
n3KhgYKcEkK+dItBvhH1GQiQriaIyQtu0TDE1E49ADsV6E5Bf2zsEozirRDUniam
KnZAOFyCNnvibjp4pX5PN5lBoG//lEhri0p7/2HYtgJDgOyoxxdbnmJQZ5YWL4zT
8Y/ESISanms41cshyt+nJ9TG576wVAO+1wumaOuqVoNip+Esfdqrhn4oWFf84sWC
vYXorE44f1cT2W1IXUno97D99YH1/0lx08NBqZIpyniVBhn+7Ia3Dr999oDowKUT
Hj6qb3q+8olArh4FtLWTqd1VdZmZkoldCb7/0VoiAoONX0VXaniei0RNMjz8+Z8D
Q4xtLZl2rS60gacLFxik+PduIG/iw9PKB8ify+0kZ/sJlVy2YqYBz4Pef+S3Y5Sr
nEd8I6KeUESAE5GosciqWO3rwCOdQCrT9vgVXHhO5g2viOqEbsmUUQHHmZHAhCD3
jLbGsyGaW+O3Bw29Ide9chdwYRIlETDa3u7C/OTG9GDD5TyIGiZYSlL7VgTWIrqI
DYlnD4L0rj9TehacOxCU7c1Qd9dvjypXyFTn0df4c9h7KCxUKxvY/RbU8X1qBeZl
C2MVcxhX8ArWjOTz3wMVLQEgT8YSInPU2ivsvr+0V++qmi4ai5dT3VUIRRqbxduv
/JL7xK7ZLvaJiyeWJdaL42N8V1RdDjxkxlAOjmj/OUq6ZpL74kbFjaOS+Zlk9Ipr
kYkQA5E1G42fJQ8szLDMmorfJHWql94ANXPIfsPexOhNkTFFtQFw6NQuOrPchBXY
VQ3GAyWU9WhAH3Egmn1ap+LqcvixxITftHMV2JISLR4c7Xl3rf7QAXcBny6M0TDW
l7194vPe/ALFPWVe19mTpbt4B8ZZi8zWtoSvMi70U7NlAOQLdG45SgOR/0LrxeTS
XyBq+pgGqLGuGzG0y0fnrJga1qkUr2NwU4JXOOfvUh3qRwlEdFsa3vR0j25nhJGA
vSdoltRxOnh5j8l+abzj4apo+W6YG3yLs0r+13NYOofAXXfCEV7wVBlMwgBARu0e
9N70iXwdswA28zTnuUCAqZYqohhegeYmQ3LaO1jaojgSxUbDSOwjnpnQfFoelE4P
3c9Mn0WHw3WfawCcxfmfXucc8Uab54gmKjxTr4AjazOxQPWe1prVz7tlARFHIrFw
Nlmo6obzchgCvBnGnNB0En6GglvQTm3YJPpHMQtEMmlb9KGE9b6d2Dgs+9RO3A4x
PU2IyPaqgQYVCJQK1FGkeOVjUhBesGv9ofqs+dPuavUJIrMWnDGeCAuHDCocbWy0
X99ZsNOeZqEg3aTdBAnDb/qT06nqPYYgK16WNnj/k++j+5Uv0QlgE7Ta0bvE6gUD
Tl8onQJ1FyjTQQlkf33k6AACMFtwZMwElzw4uHNqTompoz1SI8euZgyi6xKhDwvo
ozJ/E3JXHnZoXZciZu8Q4KDKvxBzGs7pu58PCS1cB2i6y+ILkwTRIIcG53bxRM7R
H/lf+kF2E9UsLmhBISaClNU+hmNhZeLE7g+PHABrqRWOhCqAeR+kzLqnpByPVxZ6
ukuX21UxUCceMwhouSx/IVflo7hnXB8GFyf0OAG+f7RVlhJMcElmh0IGe435W3Ok
gZOXNW9oS+BwQjJBwWVPQ+siEj88G/wiDCh7IT/EhKwe6r8ywD+mfvRQyQpiOAht
ICdWOF1EehP76XWWQM76FZqGzHNQ1IJx5piBgRD2x/ChXQ6wbSMxsWDWp5dS6gzL
nGs+PlIDORoyDnqUnKCv320jZV25yxJSJ2N3P3sr8LHuGKNM955v0Tn+U3O3bUDC
M2dReovG56L4GW7FQHpPqspH5DdhtSdih9kLc84hjUVJmkgITxzMaAuJD/pGg//g
26DW8+Q8UDtouqMCqQOD9a1KXQrqEevKrcgu7lAoz4KallnUfwlUupTnEKyrkrCC
DQVSyPwsxajQGVpMjhK2htGTeyn4CwYhWSOxDZPn3CrauALiJZK2Cf4LGGkk23YN
8JNCHdEzkUg4glScy9eoB5xwRkW/hk5nJsHX8zU+mB6MHMLBLdIssw2ZM6nKvndi
fV8IfMstn1ply+tHPFmXKpvhe9VhDYVtFhfLRcHI3iKg9czPUzyPRtIEkMhBRZMt
CkTzaombNx1Xsv3V+fr6vsoeu7UkIEo1sOgx2KmrZgvNEUFT5lgeeIF2lVwj6ZFy
w9IfIWr5nju8oy3TOli83NfW4rrJiAK+H28VtMAQ41puS3s0HVKrgQvvNTE1y3LV
eO9dqKZkNry4zO0tp8s+dCO9JssuuZMzQRvgoDb89khXUQgPwx6oYNZ/bFmJhHSn
gHtReI10V+gwuR28QmoAkShUntBMJuseymF5tFlXmtJW47ZrMs29n6O+/gT7DR7U
TRTYZQ8SjSHhUhebOTjm3r9ilNrLlSPT8Hqk0lmFQhoHulVtnjlCDG9x+98TYEkz
hBmVECJ1Jw5kr8nmzQAXafdUnnHOtpCyO120zCkGi8DwcUfIhx9+Im61BT8ZTDWf
4gUXEEQ05bzhVPUH/3kpD0cC4bh0uqCW/tJS6QMqVOlkRbHB/eZJY0gYqnhXpVj6
jV7my5aX6osef9X+TpwH0OB6XvT1TZR/aOBkfwj89UycXpifimtrLvHfjoQ00f7Z
msRfh0PyU7O4ELrBGrgl8HJh5T2jBBtMPYI5FKM+nUaZ1q78dxhwpSHhAAA6V/xi
X9I7zh/MMgY9Z2vxV8cnXNMR8ZcG+sDE9k8/6f9alniY7KeBcRO2A/TZbd9DPQo5
v1SBW8L/Oq/D0PEFxbPsFlH4XoFRIiKJKgAeOe13CtMP2XnZ3ZuExHEmMWeJs5IY
meehdU9YjjUZibvGH42Rya5CcciT+CuS4TS4a3feZhO/7WKrz8L32MELY0glDBum
0MyKdFqTpD17R8Y6LeN92rUYRQJIETHMV5D1Sg/dK/E/M5DMa/AiZSNPLbhWGRt6
rlSsYF+N/NcMdvNQCWzjEq/cT0VXE9zfWAgDcyAc4yFoZY5/L50i4dYGGMP1aV3q
NmeXoKhewVb6gHIXaadvwCCkK9yTvSI2FVz8OeclsB6g78dPFfsIWgUibEy9pdvV
5ef0Fp3qIc6a1givtRCmPN3IVQXm2mnsyteE3tdv+/a9ooH7/3aEpNH3KhKUrBot
J5qEqKBrjscixhO6/lber9UrjseIwFKPMWo250H7Hfu36hBuXRqOj6q2BOCQj+KI
Kxb+mXlQodhDm/Bw/0XF8Rf9O9xBFZWzeUwpJNx6Bf9dsM9OnX7uF3rZB/J6yMlw
OpFCLhXgdkqgBVO2E09KT6v36fyxdfY9WyZohJyBFl+OQsxcfj+qynYhsiQbyWLs
oOErgcOjVdiCIDE92cqUX06iD/SwUmvE1LasuuDs1KViJvddeIfI8jTGNZPIZUPP
zi+r4UePYlECkP2J1R8EDxvSCXdfJFs3dpDlq+eeNByCJUPdNtZS2mCqK6wb5nMp
If4w0NThth/6RO169A/mq7GQuwyc6m+nQ/ur2DDp2jxcXQmA9A7bO7YZ+VnutJsw
OcwlOy/bYLRR5CFPXeeivyoxtPni1hGHSxAJV8tHszM9//fdMwsK2MhE9W74Y0Ch
186XB1VkqYMSvMEt9b0dn8vV7l2UjTvA9kKBy042lqT1g/Rrl1P8kq0gb6y9EJck
D5Ug4WJ3EKUI4Ml8TPFsFRfWvUrnHoOiZEcQguzAPwBFHb2mS37c/EHd4HDr6b9L
JAXeuMA1MGhXj12hiBpyaxTaRqkZyKrz45AncxEJz/njHwZYfftfRq273JT4iGxt
8FGX3Hltnv5p8gOUFx4RnrGO7kbmYKV5S5hjH4ls/7yuNU/JBzUS3tCQ+PNt/dMn
8svraJA8jBgnYLzZ/8cz8HPTrI683iNwRn0I//IJd5M1WdvE3fgjjMM2ktRIQ8Dk
uxFGADiBFLyQbuznWJPJe9vFuJQcOvHdBZNooiUvtNW6YgjgSty3XzCgZMpu4CB7
dlBcFZCtxH8dq/rJnnYlbuKfEgIJj61xKVfZUEBldRvdyq2Ifn4D4mfcNxs7sW/N
MRylE9rzWUBTVUraiVP0N8z7FJiIkQLw9+Z24KEc8i42EV6qdgdl+cT7+V6zEK5N
pLPbH4vmLOQ2TYbmLmuc3f4sOfUnT2pap4W5UTNBuZ+51Icik//bdL+2pH93VHRd
v0yLku8fJALb+EP9yJoqe5wdv41xf7w2jX0Qrti5cP+hxOWCyXdh8N2DHMZCj+hU
sHPNILjN9XAcUI8FKLy8FGRw1BYtvn5R5ypyxkmT1XKkBqE2YglGCTWHk735sG2r
gRHkp+nN3NO0X95zupGl3HvThrX4oDJLVskhmgDd/WCjmrjen/xb0oI2npVNENLV
iq4bxfHn0w/3gwqHSc2A7CgiTxQppSiE2N5o2dZ+ScFytC6L/Pg9mJI5pq9d2LRB
4PxCiaQSdfVXBQtaJIdJWWij4pJERuNon/H69ggx6sGUvg1i4RyRTnaecDDT7gZD
i1ZR2ohWjDabsPyFVJtO4AFdPmbpcWlt5hey70WlpOVoKq53p+68hQxlcv4tSNhD
86/fLayXf2XlmUudtvtmqfFE5XiKrd8sMLqg1aQ+8irSwPn+i9naRkzQ5Lo3+ir1
q5Wggmg3QdvaQdm/0R5lQBf0QT41qXfcKzkSYrkaHkZ/PPpppd40oVmXxPewex7v
HvRZ5/+iek5bQZjBelCeDTohWNUyw4wCbwLHAuGb6REa6i6LK6hp9OQuKOOSlnxe
rBTv60CCHXA4mFrq0sig0f1HEo47958EMFd0uhg6xbzIcT0hOCHhYXzm7XhIXvPU
201GVNfR2sDR1gpJamu7P7dlHIDlqGH1iZU+4cBmH59Or2ZNjsgJJMCWmYG1SLTa
0/BmSkicBz5OmCMZdnSQuMzWU7uzLsHxCaAnFJxX00UnwYM1eCwrSV7YOtr5UmoO
NBB9lcwyYSWOxgwHStqvgeu9Bx1XCZTlrJbeWzYvTPvkh2AlSF9qcvgGf5FNWMmx
9CQdMUh3xZjx8hDjEzfZtGYKd4nmPrP4W6gUAepFTuWYhjTPLQU3pHW2N4MHPlij
ZpOFuxe2z0ssSimeOn1s7Ugnl76VWbAyZKdaOB3PBKHYK9MnHWOknF4fBanH/QB9
5+P9aPRp0uh5Km2L/Q9YlnPj3vv3RvgkUSyNdke1/ODZ5GTF0AZY7mw2YWegM5b3
3aJDCcX+4pyg0wsUGVR1s8DpzP42w3gVam3hct8nJ5WrnsqGAD3TgofoynfdYkmt
jL4U6wBWLpnoNT7Dw1c5A3pc7oh+tbxYxC8RTg0HTy6w5MtOzAp1O4too9DOXQOu
gLkYdSiEF57wbvhv3bDHSMLucC+jjDiwE8xnxmuwaQJT3BVUmOIMZjxkbRvTA15n
iVk6OIzz8gELKunI8RAVeCL7yDfeJF2uztO+RljUfHgPvyY6GvrrqlyLQMxUdOTU
lslZT6OBQE9uoHXPZinyeiscpwdP0S2QsPRyc96djb0mPZL8DvAzAc2fpm/KQWbx
pDv1x4Kz5DY+ZUweRZQoSEz26Fa6I3u40o0+Z4+AQ2jnm9KUHIrArm3dn3Hwf/Rc
3ipBSpvl8Xta7qtJJmjWgmEGl/2CUyCzzEmX/Z6uprvoXwLk+fYtMBYn/3uMfdrE
11JcBivJs0aKaCaLc1TcP1Gw5Msjdhx4y83nUVRYt+h9MB7jOcGoe8vY45XcFMao
pc54xNsdwNFKazr1NGteymmbx55+6v08fr6y9gbhNF+sheMCWpVMPHjXu5BiR6O9
GhYxz7XBuELqWS+fGVYS10Jq77jVKSeKTD8DEL25YH12v5hmF4YK8r0qjxQ+6o97
V4qvNeCD15NdZo65rOWyG9z8sUXr+ZLYrcaKKPWnErZu+htP6YSXmx4Xk9t16LNX
k3x1XsPYtkIghnFPlTiFB8Xixjzl6TqqZmU48FcfG/rnuxGqwCkktE6VxTSGwKMU
4ONb3F8iJB1VfYNu3IFyyAZyht9NGqcaeAGpY5WvCHFPhm+UvGEBHPM6vE3LJukt
VA6NJMe8SEJr02SE81VonasB1QPIH47d35hkKVU897dPhsFMWpP+w4kuITWPCZqp
oz7O50J2ny8hxbNyXKxlbonNpHl9YZOKCFRo/ek8v5ZAhUez5WqrKiSlQ+phGafH
SLb51NEx8pO2Ezf1Eusl2gbdR76bcymjmJoIy+C0HcDmCWKhzMLXvHDP8MEMJNT1
zNOzDOm196w5A7NE+MHOLrDDo64jpdtgr5BGM4i5FnqEMZHRUm7GLLcztpi9TQmw
CW8cwx0UC1GSpJ4Iwauge72BXNpe+uOpDPsOrXNgY9usgdLRAl5WGEy7erxb0DX5
twvrc0/rEzsac8YMQp2q4OTxG/L6GL1W7z6bLCX+m8/Xtc09cpe6BEmfmBbjDrWI
iLjoN2R7dKBlVoswmIrIDzvnxRWJagaiAfk29kimHfFCTgYv4QJy6NQILLWz0mAA
VtVccuzacV2w6PqEPYLH706ABBO+rFIPMLWVDM10PwOk4NMVoGkTcM9I8ZUTuTx9
5cMEKcgqi6LQdlgbT7NQahX7j3I0/2XXl2+rs2DGaygn/wHZueGQOXapv6uzG4y7
eEUoImeUFgsdLjVgxQyMeVyGCPhcU0wF6mfbxixvvPIt/l0281SyTujEHGk0nnrQ
i0rCwcsDQVoZQezlMOs4ZK9vhYD0NOLksuuIcQg/1MBu7R+UAvbngsKNT9Q4cheZ
fNVVwwP4tN7Dyh8TUBxFxojFj4sADr82B6enVFCnPIYlO3MoUBCpV82dzUf7YX+g
deTgUj2Y5gji7RxU7L6Ad+nZBkZpKfTFmhykRYLqrByT5WCOTBKoYW45tcmSTh/H
eGeOi8hC9RF3sapIG4ZboRg18CXzQUgpstlrhp83wroDNMDYrOk3itUIvlS2CnuR
lzuxae5Oe1SajU5rNaRbTV7LIIqAitT3hIp9scJd7YcRRaSCxw9gSHcU8fju2V8E
JVNTRAZMjyCfybjWNPMTFx0U4zYbICrZQTqmY0WEkc9rCCBYL/XTPI65nRdYS4mL
IkRESuqT/gaCmfIBJCyYQWPX8Jqjxm3nJjN2IzVL4pz5+BbwKymxBgQHfgUc6uVE
+Ija0BN9omSd8DUyXEU28KmwAwQshngtVrb+JceIUEY/4WcDRNtdMuDJLldT10pF
ZHuicAhCTBd5IQnIDER4s+vIZPhTDwQUL82jG+EdiBhiJtRMtUPWLJWJvN0Lp6Qh
QJANP54ZxFz/tWcBfG2QL6Dep11tQ6p8rDC+ZeBIPukWqbZijqbxeXidUmZaYNba
mCmr4vWr8WycDHIL4kR9ELLrpHK3CC52qTGOtMV2ytc3KzaZIU+6ObOS9mNCwbBW
V8aeZCVUGidPxRXa+1HZASE+cHPOY8WxpTFIzKaRp93RqtGod9LIZCJiEomfFrx/
35MqU0RTJjqaxSMWL5S24gs2szsbpDabvQR1rtf0QGF8SxvlVKMQSFJpJwnrM7Eh
OSECvaLeqrS1pZykRZP2GIUBIQKKiWA9EafUG/tz3JkX9IZOOuqw5vSif26GKlTX
WlOmd8iCYzKLLY0o0c/exfSulb6ktJWmVe//amIUMB4UrzK1As2aGTsGpsQSC97h
n4Lh/7un27lWlhm9zMbRuhSmaIayLJP/zy6gGIX6QwjetrxVveU4WtjogQM+0II7
spBCiWxeuhKf6ZrgUWl0zOaKXhBa/tVMmS4l6Eacg+5m7skxDebzY5SpMowDkLX9
YhOXtiVa5vNU4MOELXCOlhSsBOYjTgvQ7QaFA0a2s1Vnu3rVlOoEnxqtWb75YuLs
0fn0q897B87jtDbLSfhUjywHX7bIj1ChSIFAM3q7qkwXEu4aU1My/Jhcx0JrqzlA
zSolC8IFO/G40bcXeswURzYmfwha4OBIMWwooioDt9cYIxn0+vnoT0HCmyi9qzMq
8B7vwVCZXuL5/gfMwgjD2/R2oFXxNHIn7KC+ANOhUiDTCtKPCmSOHv8zrQLL6Zlu
Lm00R90hZ0Q9W1wjPEWB8zymnduDBZ4QUVeO043iPs/YRo2PepDiDbFNh9DfemmN
b2kpzhmMtXF6Ms/jvcBJTQ04RWr8FJC24dKUyIy++XMq4jN5zhFExL92aJc1UJ1U
o0dV3LgFB66Xr8406QYL7spJn+HnWlQTxg/VPRoZa5RyWvl4r+jfTD6qEag2+2v4
TlDgTE7+c1ccosYXIVZkjOuh8QqTw514kWvFaLUAk/ldsYBWFhMAa0wvqAR7654O
WDCDoyISEotBaIc2YWtVmGHl9TDihrd5IKBIXonizDPDHlGAJKDag8MwAQO/Brgn
il1/KzlV2RlJtGZA4en3YYYUMyC1MDBvlQgLBBGBM3GVBekhidkp209H5ravLlls
SL+3JrTSS3FQv4xw3bfD7WEHBPe2k9O2DiKm4hOwq2KfTyDg2VOF+Rb2sIfjkCJ6
sNMqrH5dW/mNHG1BQNmpantUHz/+UQjmdoDUbuE+i3yx6MkmRyqQKhc/DzHaefwB
jT0HuPe8Oj3fUA4cGZUUje2394KORfAXGOzfeK+3gK0BxTG3CL51Pzfwa7adQwji
IukHxoIXI1rUgU/iazp0+ddUSqJ/RK+Xkfmqaq4w1QAnGWOu6G6xPX5FAEQQM4JC
rlZKycj2RFb2otGtzEGtzs4dp2dqJNxGL12HP6Iys8RcHLElMg0HDpEQ6nGyXs98
t+qBGrLdrnVkN+x4Ulh2VWypeYgye+6/liytTNsWtnMduD0oVrWTEC09XPMzN92x
L03EQtgaicarWMXmuTduV+8w/99pKBZBcwuBckvxFxfsgy7Kzr8fZlg5zb6ujPmJ
lDITtOPIU5xatXPlyEeor+/0sTzDGkn0KIoqoytdviJ0QBLJNdjw0ZZJbchhdngf
7Z1nb+Ofkcl5DEZjufWVAKpsc0iT1z7sCjZ3lINWnOd7aQBrC4rmLf9a7qDKMn6j
PdKdW098/4b3O61v9Gcj3h6e3zN/Exjvsf33LycpB7DF6WlpW1tf6KmmjFztOcdh
p32ItfJYhfMLPYs7QkTPtu1pZj69yS8vmF5PMkbEFaS124p/ZDswmX4hG7PVOndS
nRgX8woA47SboZVq61aS1Ni8syzjpOuB/vgLyMTvgUF1GU/rGPF1En58j8DGpAtn
lMVbpwIaw/WqJ43CcmBaRBhjfI/fH/R2EmwzakX3sofKOJyUdeY/HI/ffvSkyNlv
C01U6/mxSmN6sV7z7P8JLFjmMgMUV79WArgGCa39ffPgfdy+5JWC5yLJZFnsub3z
jeF2Am/Ea9i94/mKsULPG82ngz/+rlBtQUTQ8PGDaWU8f0J6lvZ0e5C5IK3fPbPM
7XY2kElIWICk+GtITSIjVdugBDCN8OiTiQGR4RAO9kalMYlMGRLK9rNh+ed6b8ES
zzw1jPLhC3tzPLaBzrVwoVszgbkSnRtTvH6i94WrPzUqwDbaR5O6H+6lmHLxqd59
SC5HOSIqxHw17KY71e7HmzB2Cq/gIzkSgqGzUkp8TV4YggZxKKOM6PY0BBV1jTzg
GpeyxJDKOZ5QY/HrgdEI3DovFqXYNVCvF5g/OFPCKxI5LglfNS83IUrWdNBLrBFE
V5v0KHz4+ny/sGEDtVOj+ekbU0IAehTu/ZEJ4tthkCn+AFD3x9miGKiYwVcmLV15
bZEoWM7qqj3UaZnL9HuOXJr7fA9qwSG0kCgsKrGV04xOsHYqrSzjXOc0EFjSPm/w
cRizpDd4kReORYxFYMgoULW2yhcWoEEiquSfKEHbNLPJBw+0WrjKonmOEV3A6o4f
8dsXTgPXAXLDIyp8vf28n3YRUspeN0fXePMGf7rna6PDlKsRqO/vuZ/sCBcgf8WK
cRk/d6/djoWzjRX/J7ps8iHJuyMPteGYgvE78qxRlthSzJs2DVEDBt0FWZgoYtJ9
ayL0QEy0wiBcnk9lLga8YAm2+lZfZMinHw8LhMcZjJRIuVLBr/m5WH4JQBbRnruQ
c4zpDl4TtRr1wdlGo5fU85Kf8xc/ejUWuirRmo2GmgCHBLDeloKEyBbmXdR0WvWf
yo//ZWwCvHU4SIXmd0+63D/ZMh19fJcByYsRROtGB5HneCNoIvgDKFOLlVdheALN
7OTs1zZzsNxqVm8Z3jY7BamLjRuTSmn/AjQ60VrzagxPkmjtksLctcnvWo3aLN1o
DNNBtZ6Ihh4ctePQ9ZUK5i9SVV+/5zwY0AgwTCDQ5IiIkBDaDMU5q2IdMBdC0mUA
k01t/QZu8PEYlYBl4NzoaAd8GAnhh+pnZz8i2+U9QSLVzg6suwbsnSLKaUij8Dx3
/T4hjbBht6xKpfxm5ZIN+jb/poBoZkSTTZylUkl0fZ1LzxKHlefdy22Fne9T8Ryr
6p4c+r0qlFWGxUHLD/W1FYgsdNeoTlqAPqrQc70iK7YNu1HwtV8AuVtw9o6VzfJW
mF6k/HviWTXOBy5y8mrXGC3ELyyDgf6PqT1dK/zza8JpvqfiEhd/Vo6NvvjEuQhu
cYmbLgaxnX+wlezE8nw+YdCyCtcvbxWhVH7S3aNfKOyii5xbo6LmoShJmYHTFPTR
hSsslYfmwrdyy94X4r/UoyPeTIX5onM84KXLkpDojFTeXPJpf0hyCkI+cCRJuNbH
L3f3/aE1aheIReEnaMHQ5xRzBHOUjJn2lCPyhVORZ8mBD2yST22xARiszHrDCOKZ
PlHhv/e7dHrY3nbQR74vCXx8uQNRvJHQCG0yeWvw0MqQ7kr8k6t7tvSmZ1GcaTkx
gXCBNt0xffFawz8/jWZBVMCYmicNUpm1joI7covwbPS9ZSfP6qta9fwguurPBcHI
xm+yW709ZHZoFoOAtAdqqzqGaZ3BHPytgkB5Q683uXQoI99AkOuewqwQRLO82dzt
ZMnED790uqtNi5BS7dLP0+T5FxdDcws9qVpbFtLPdrwIZ9rdc0g7qb9z9nyepwgL
CA5r+ID55FRMuTyxBHlH1taY3n794vJVGaNk+e+rCuTIMD3sypgfPggRvlImigjy
Cb2zxYgB9EPwOFzl50aSG0kN3uvFgrPGKpNcJW0uFzQBXeYYxpWpd91+xP8X2RH2
Z8QNEiodsoMx1ZVxWstdfxL89J2pjnKKkPj14S2wdX3Z3wJyGcXGiB+/1Etjhyvg
N79Wjg0hMQCFNwIb4i0rG/CzddFDnvixPXT53OBI17FzRmueWqCOharhmBU8hdgy
hamg6SjiHNQgi3PsE0Pcesx+1TEic0aRt6wgQYPN7th+wk97Ro8OOil6blJK+CL/
Qypd4BceobKOd3fHSsruinnYYEidlazC5c0OvNqUn4L8f2lvP2guq98xOnXE7P4R
FnN5jmpRydjafkOWFjWIrghMlUj4OOQqJaylyM+Twv13OUSI5nd/f2igVNngP55p
2k1AB2dEmyLucHA+mvn1maPp5IlF+j4AL6JzGbz87YqG0a8bqASqn2iZeXJ2HckT
8QR5tCHRLWW8TX/0YrsRcocYKBXj98V2o2Bdr72Zs78ZCCp2f8YDWnJlozdFYMCD
NaWSTRb599E12luvKeK6p8CDv3YVQbE+vb9I3yKFl9WdgbLP6fZFJQ2PeW4q3Kvf
IcAplJSL2Fwy15nb4eQ/LOs8BW0j/MLAVulvNB8hKxxEL7ZFmiVmCmb4uVWuya/U
NGCYaE6Q4REIX8gLH1QcPwWrjixUjmHJONN7rZBQC1uNxRq6zmTqU6vjj25XTOVw
+wrShogUkk6LavHzI6A9j6xCBu9R/DTfoX3QTiG+BO9jhUsOQM0QUuRgyTe2gSHn
zq5KV2JiuRE0Y7VpEgMzKnMVwyVfzeaNlFGoCnrlRl7YNkwR+SwMIcj+bGRkXidV
eWYmrvYC+iMqdki/epcNL9rOQLQa0T5R9C0uzlsmhAQA0A1HcjGEV3Xpvx9ZX+NQ
52VmTYbnCqLHyR2MP79nY0znFt7xEj2AKB9aQ2UW/LZIIDm6SZZ9fetZn2sEd1EZ
7XctPbTIGH2UKv78alwbv1DBw1J9RjM1zT7UJfMOfv0k1xVtCkd18+f5kwi+JcvT
Xek/EcUVF8iPSpEwC4dHY/k4JTGFuuBefedkbXC3AGCsHL9VaSuNQOXj+QNeLqzz
Sz/LO6sGp8G/hobXJODXvSz+PH8S7cjqo3JdIa3uxMWwaEvQ9xYc2xlj17P2/sIu
zNtwG/tzpqiQwJeKE10I7A5htDG56mDf6AHDXoFKIylXzsq06ltfuGXigiQggCbn
VSAKzzMXwIuNQuT6+EjDNOSTwvrE2OQffDFtReFctfp6F11aT/dpvWaln4P+2sUD
Sv8JmY3OtGjyhsrAHYG3kZKBNfmFfUhGvBjfoxIH62xzZsY5iHlM0xtdseH+/nQ4
XAzSxZRB3YhT48cax72zEre0jvz2QibL1H0yHO89YMaCjhC8Y8WsdYFkLc3QFO3P
N9YJ0C1zUfdDQugkLHfvDg9Du4gyzcf6LMy8DxF4wveuEzp8uHHS2pbXKzhG0VDF
vDZ+RQQcPyMIXgHYsQdMoIJBNymmqARuDVoQnsVhvCo/tjFUQLRWpYZRHpS9v83O
5F8yKYTTP6mJuqU64Ts0DY45FBjn5dB4Sqs8sx5rcMtuQqMC1/sY6ge5rG+3WOHS
yr89yNtYN7pK9hJt9/tOvSi9S4VnkG60KsGK2vseWdADcj6vJZUqNMid6Y7M6TWJ
ws5nmvBgyg68Dcd8FrPp+ufD0o+RAge0SdiJuBeasAeU2HDjrrBnP2kH7lKCBpZK
gqfQPPgAQ0S3gIGw9GZfTy2lzl9vaw//6ql8+xWid03pmNW7HqAVUhtJUHkbTCpR
KPOrBeKlheA6lUiSSRiyM2SkjFHGPfN2ZCdu3WClXSeRj0zFVIKI16ZF4n+h1xXE
ybsT3TUFpk2QVOdzbWConjhQNTa33UC/xUoBleY2IWXOX39lYc3ENFDLrn87OEDR
3D5eEOO79hJcL0E0RIes08sa99zbQA+CxRYOA0pgXE8gSit0qssFib3CCL8WpzmL
oPNI2eNJGXLvJxdGvFyUT7w+XayXF5uPomRpDo4hvmJARV+WK1/szKZrhpmCnwPt
uR30iF5cllosrInDU8na2gSXwslu8N3LJoHNsuRODWOJ4gbcLN91LOCILce850uD
l2C9h3eI+5GcuxPl40kVRg9sVQMuQQreZDcj4P925Bd7w8KGmKithnOgBg6m6Ltp
zA6ViEnbd1An8ecVTqYVHAKmEAmnKV2Xumu5HZkgSUS5/EtPiBCXBUz0uaiuFbod
x9L63cySza0uLwF5KOHp5UE53Bjn3Lj6l/NV+3AjWMnWjss5q8KwHUiJ0OXF3pza
iwR0nZ+BbPGU6TlXsdj5yk9fuWcF9Llqs7/HANGgRetxqsK8QOMbWPWMlTsNMW7d
gjx1OnXnMvCMU1AjGbFLJAm77Trv38aUoUhr83tHfkoe87cJiuNF5IRK1LTzyfFS
s176slWzPx6c3i94Bjn6HmOAspKYiVJQY2OS/j4CyJBs/IFCPbrySYpJI2QjBfNc
qj3npvgMakj25tdkm4pgcjv9N/m2H69NTvMdEwAlMKGwwBRqdWU9KH+use0V4Obz
GMuL1yDKpeypRScow34G0WexbKTWuXakSg3puVPj13cmOLoljApDc7JcgLZeJuRK
uOq/bdn5144fYTD7z/dq+rWNcu/8lHIASjULHtIlAJcXMWNe2o9mbO+H6QfFei/g
mx+U2X55ZWBngSXEvlfql6VAasj/31UzjYJsSmvr8duiVHTcxJa6PulSUc0e0BJ7
SokRU4eIWiI13YkQNnqrRFSQjA1iq7pTEJ5FoVidmXHsHYBeiNHTF7jXgPLssj8M
8PgyJQoHGnJpQubXXH0fSZ4eX6Q8/pRcOe/RSy1G2evGFZXS2zKVWv16jc6LPhAs
kdyXXQnJz75J49IP7k4fAg6NXS57j+FmExRK3KHnF/tZsAFuKZCEcsFsQ7jepu6n
YL8X1L2StPXaLGJmx8bnr4DCpYfW3lXh0STuVh0hhSo/tgHoAogZ12EGqMbgOb0u
Z7qrbr4+UbH2z8P3UK6q8QAy8i3cdXiRyRHnrITiiwJiaOS16wBM8QZFU94Y2w8i
8/8SN6+nTE4CZrL8ozWO4AQBefa0Z4PP54vQd7Z059+zWlTEJ4vzzE3OVkHCPyhe
LS1n7GvrNpJp7sI4283aPaYLLILGSlLlHfa0+HEWYSa0TbVzwHCFlTJZ1rGQF38e
Tct8Uipdq8zcC/gxjHnKMI7DEyeLqQQXWQiyVwpGoB1ipAoXuc0lndE643ex2fb1
CSTu/VdmjCIVQ1eMjzVVaIAGZJdKq3OwDWpP5r+kOiNse7NQs8ZXvWiGnd7cFLbV
mBZCQDwt8R7TmZGMiC3JfrmFbWa3Dngx/Tg3jN++z5O+UDmAxyMI8xeKutZOesNq
ybp6OFxrCEk2zmMRhmZcWYY02RvM79l9W/mDAnr8ZgCd1iiJm6Vo9j1NZ3Y+jYMK
NG7xt07v5eseZS5J2QxviPIlyESxkALCsIHluPC32ksmvCgvveMc+LzJi9+55bXm
t2LdmX5VXKr7U2njEGKUIjrZoe/2KZ8TpoBW6caIbgpelvAkLGXcixkccKwXQ1Gs
jWKO+92gaB5/uEGlw59a8vCVi7ejlSpspMFmt6DfkbisrRM1YtkCkmgxmx85+5u9
synnbqc63zsl2o97oFEMZ14j5XRHUr+QciVMPsYNcFYFiUn7v4yoA/j9EBH8Kfcu
UYODzfnrz/FNpRWs8Pxso/hYhKybwmRyOCMgW+W1y7d6NDRUhZ/nOmUCDQpe78r8
NrR2jrAOqw4HMQaeOYHCFB3aMM5iqRQeW4JUT2kqJx7tPreureKZtLw7y23zmGGy
dVPqaMOa4MqNtEn4kimK9XdOvMXeaYr+O1LRpgEg/nlwI/HBHV+rRV88/2yFLRFS
xAzoy0nAcEXO+SNuQuNNbwaZ6o07Hm5pXS7bZZ15hGPcmc/tVqwX9N9p4hTybsTA
0P8jI5KRdUvrba6lWVv/i0eC68383D7gW2/jXOLPk9tMAMwFIR7vQ1sGBXDrL5mu
SnC5f0QSfLZWDWmp2Cqo8fhUZMWyLGB2gAIOUz7oSmSo4ZyAu8ktOX4/9E+ImdQo
cj+tvZQdnynELp/2NT18BOPE3ssTplOrBFge8f2FJN+adgyAqSYVll4B/pvc7cQu
EPupeQkDTvLH9LFumnFOzy2Mrsyd3avHAn8KNyrLWxwC01muUDy63z25h8QkFQmc
A68udkxdx5MerTZfiyYuh9Y40ATyTQbtLq9y7iCQYtSXhE7yXeM0vjHXiDKRzPTF
m3udR9MzM1Ydwckfxv4ARpUqExBimbrXBfujO+T0qtPwurcFiA2i6TQmz5nuY0lz
z38bDBtUVdkZeOV7DllBCg2OWkApoIi1e+C2TZ0iMiHZOHTVH9OW/eGKpavA6nJc
rHWn6QCQKl1HxiLc0Z+q1P7wMmK/svFdOX7OgRciIc12dx+tZ5PRf6+XQ5ysDwR4
5uqDV45Cfc8gozh/McQuoN65NfSbEm7uQa+b+YpJKUC5zDcGr9M/CbFZHkjnNgtC
wNvJqzw2vTnObmcewb+nXQ9/S7zMsdNiaF6q/EFV0yyyfARLB/UJnawPIeh5V25o
0sBdW3txNczxSRlsTeo0YyFz82KbAEK1XKG+AV1oKwy58JOwypgRKQr9GkiyNcZl
QAY6ZMYjCKLTP9zXKFkrVIZGDytE4ot30vQiNgTz3Qv4loSRkm0oxhApccwr0iVg
ah/Wb6fRMebvNtu3wnVEx0OqJ9KUZGfkIW8cOOXPzvZFZfunxcN0K7QY99Ws73GW
r1H691+DHB1ky9UmsmaqQ5nbbnYMj3OCP8gRdXtffinJWl/1FuehEPDUsoEoar2f
y7rc9IrBA+ay5fK5Dl3tF2/VcQvp8nCkfOwaG5LqntGKHhphUL4pCHiwVEcASZ97
AZ6oCVSOApfbkrVc+GST4bJ1XcKclskfgw4Ep7az5asZ+J1UR+WzAhUSEelA/j0T
6N1zUbBXSMy9Yu1Aw8rJZSM/x2rgGylSKBJY/n3YBeib4ng3tnXmCStE/YclUqQP
gKuPz67i6i1/8aC7wTMKK1OADGheWe1mi9xC73BPwclzQLhUBDWEjf/agUeaHqey
Lx/AZktF8cU+2moQ71cKcqZwgIwa5El/eI3KrwMcEmZWLNBSWAfcB5suxjA/FDpF
nbMw0zvZazPeVm1eK1/tnRTMv6qIbwNBmi27Djl3kzCTZLvhUnQGPmeg0HZiMJOD
89cRmAJvjvZfB3oOyZfq7Ofq1+c2abXxYpWHhoze94lRx5zB5TQzBYH2nMyWqTHm
F5yaks10M83udQrvtMw1G1e4pfPNTxRo/kZwpn8C51Rc/O5t23hWON6xPCazaHxX
QfW2AJDMay4QRrnGHlIDgnxSXmGgtvR5cJqRV3yQZMdFTvJj2Gyi3RP9xPS4+sAw
R3M6Vn8NoAo9WP7/DcdNWYdQNwxdbWAKVgg9zcdPvOqWZSJBryzhokmdh1dc3iky
rZ+2EGmlnF0iYXlR+AEZvZAo+aMeAPfIhYfTtAxhmJGEWNPaJ1RGpo4VR1OCDQ03
451pVaUO68Bn1HRV8WjSQ4/L65xw/B/lGDw0Rgj8hfwbSO0rMlxfjLDm8GH1HLIM
N5ifIbXy2H1F+BP2XuII4CH1HLvl5WVEUZgUevCDdDNrpDTEWJVL51g3JD91+zdX
wgGcmTsYwowSIBuBtZ89neFa5bwNlO/AqmAQMn+2zNphfQqtD6b5b8UNuRzylv0Z
7ZUwpSRl0yHuwhpO/vxihfm+tOCykldXEh14HSgshPqbR00ay20CgCGv30DgAXdx
ib9xEH4i6wXMxpvRkYE5J+oT4iAMq8fynbmE9UvCFQWfEuaRJ9gqAQJclWTX8gCQ
vF6ip7+5ge1+t7cqHQ4gfxRMwgYTRwGEa7beN0dbDLaM/ueu/JEtsyfEkKVbRRpo
Gp894ugV7t4LCI2gg6AzeblJG1/OoRfrVgYbFWhryjJrzVnafPSlmW29EVvfv8KG
jXxof0jbnilfIZkLK7eZ4g+7L0epjzt1PpFbSfF1CEs4hOpGpDnfRsj2EwbZkX9o
/+QwwYZeOCNgBT5SIDV3BZdpes5HKxWrurg8f75SATTFTHQivQuzhEzb5P7T+hW0
HMbZLs8JxTMznM6g8avOMQe3ohoPgKd9pQ9PX6pHvj5UP3vKTrTDVK1cZtJvgxfD
50J6s8XqfHq/SHrVe32Rr9ojHscu+4cMBwGHnbwLT10fbmLs3qAcUUN9GbWicP9x
nv7NJ/hgnTUCeNPs2DEBjd+9YdvMt4uR7uXLBXME3WxELx+8n7YIT476ao1gGw4x
nOdqffmV/XTB4+co8LAvPHhzDfSdkkpxWTbd4rrNycY5bD7ep1efxRVyVgGphtv5
NKu9pCibt/JLj6eQQP6bqRgm345IUKgesQJrjPTL6X5YW4hqGzjz8GTv0Df5s118
v9BkO7C1NT+7ioOF7HaQjlwonRKNGbkoYfzeVa8H48qQXydI2etyy6tEUUTvc+w7
C/LzzlBemmj0sNdDcEDMc0FjUHfDAavu63fVAl+mEcJ0VEsPS6EVGCiHPshH2RGl
ezBXft01Q5uap3GARJe2QcIcCLkrN2NnoIaC5skBwGVe3u1rpJD0pxXNWa7XNply
kB+8UJCfTpRGvxwW9UOsmuUTpe45coAmOly61GAIkKOHK3t1xEFczQotKkwWa/OZ
E2AJ+fHhfqg32HKkf2Ux3//ERpr8To9u8Fgjd2rhmzUduEpeNV4Mnj43E9gGyiTm
zIG1xLEPMPbbsIW2MWq6jAtZxhfD/ayP4NY77JkaacnzA4iw3LWqKjV3DmqJbh8I
NJZIeEkeCsYhngIr8W4cQ8iKiUsje1rbcAv3Caoz07gblWbbLWCrw7bzg1mL9LFY
cg8jhaiStwcH3m+ExnyNAZLYrSsLijbe6MZY0rMCTwpmc4zy9ETBprsDBu9TIrF1
0Qk3MP2+7e25hEnTmURw7hEEMQ8gzWe4GJuGMcJFDt595nM0+1mimIaHRtYAU+xK
xseLddq2Hz+2xKZk0QrXN39DuW/Ie0MSADXExluD/3TbVd1hVKtMxAd+BN+jqnDh
y/+NKxNM0R+PUK+ZpUOCYVmZYG1bJU3EEKrf8YooVaG5xIS4xxr3OSbqm6y6UY3G
sChylOef9RPxepNvQ2f+U3ET9hZAkeGVpIxpqaI549BG8bLfRynMP2U2SVcvn/GJ
2u8opS1ZTAiBlyG2Yug3ucFfVO29llBupzwiXDjwuGTy1y3ULp8Y/LcnmjyWvuyA
sKLRycccTgTFw9VZi15aTwRQkCYP8A9vECR3Vx/3TyUfQ7FUpLAZdF01NmL+Uk3f
x4ORr/i0Jb5hBA8LtmcJ2AtrADGtaAziSTi6873XNFZdXlQGuglSqYxDmjOy0nIO
+1ArLbFPZbNryMyigA1AITkbdITgYPIPa/mjHnvyZzMfT9k/o4By+tYQ3KDu+1vj
SD1KS0uhuemMu4XYmaQE1YGXoKA6tTiGvYae/esJ4VJe+rJdDAEkJ6fm9WaF3xHc
Ky0kE04F+SjZwakpU7ovBgbopMd/CEN/mFnLEkhxojwrvFldWv3tdND87yo6mslc
RJXA7gvv1UpmfLAZztgS7845E197pS78MIzgQp8EKLH+CbaDj9Qdgr+m1XeH8HhM
6md1bDvm9eeX49gGV4cHn/3h0SMH8VSXTugxh2UTEHjU+3OzwJYSH+DjlQN4m2it
zz+Vf5rCCLocxJJlaQWgEXO+9AXvqKNyzuDvLMp/DC188CLHdaIxw9VHqD6nbEJA
Dm+1cvvDFZOppdvmxpN+sMasJJ1VKQMth3Ng3xqhsXysD8Suq4RF9Fnd+Wr5HOPw
oqoNCRMin/flsLdlH1S0UbDXUEKTzlkcAqyAQWzDCczgruwcdc0rg69qaRK8NFjg
0BAXykaweG8jgmc/j0pH8KStM+ehn5OWnwFdAAY+dRqPZD70KHhsDEWcQFaZleoB
z1N+9ZziTF6dMkcOj9NxfVeJ5h3y9hZZxdYe4fB/sTkwzRF/eCB8z8XGkWG8SmXv
Vsytn3KyqqcTaYNUEF788eFnsbUTDiSRLq/ot0tJVy8bi7S2m1jRb5p5FcOuXvO5
x/KWpf3Byj0J2Sqi/B1eE1jAAbqTpt8FZ5x5+TR3ipyfXWEMB0nmQsetBDMhLy5/
KQ1//lcL91ex6a1OZznBKft0On400NtsC3WhPzszpvnzcf2q6FQifKljzY7xrJ08
9kNVZE55B9yDYwH9D5nYoQS+w4OnOPDjhU4IwBpi1V8xpNpBPV96qIrUSMjh+2Jr
DON3LtVuP+EoOKtGuVPCLy5OKpAcEXUb6PtyOm8tflfojYsFs6vmhCAnPKQ9D9zB
zW9ijmPNidXSC55UlRvzJciXR2H1KxkXhWd8HWT02xUBoYtd1TxV/9qO7vVpVCW9
1rShWx/EGscK25VpNtc4FcFKXNOlj2Nso5QiE63LkwmkfbdcV2zm3a1blaBSKpya
TEOO5TedeqO9Y4B2ME3Ns8+v75VueD8I0ItOnyRZCHHwdesludPjRRbg1CLtEQUl
zIUiOrEZndCtznhogQQWlpcjmLLg4lYxKRAU39kBO5Mgv8DDuZbnEHTuy2ioaU7j
6GWjKdjPvvSPE9kjMmtKUMei2viq9SCw2ACjsJEqV4HC4+SPvDczLbBGnLO15QxY
hmvvyJyQWZP51A0C+pbwkVhqfSKu1gPevDWvNLWn5EGYE4pPMSRMxI6fxRoWDmVJ
cR6l4DABizBOHG1ylI3TgtiPqDjxiA6pZSXxuMpXUtDpnLpI1v1EFBsHt58yuHcW
6ciF8JrHj811Hbg7zvHZdm2iuUUPeGXbOPA0LvjXVeHre/hlNLZol2FoGHbTK58S
VfWdoVqtFIhtC+1v8axj9Qqq3Ci13WQUzbIqF/S9jOmzQap0hYiJ9C9dYuAcs8wT
Q+UN003XytlFdPZi0be3yH00rHFiDCln/RJ3mlEoikJt15q5DIQa3pecUy/2QS77
inK9XD4NreDQLSIf6cS0QBajd8fF46+3vUVb7AsezXP96R1ViFlIpJChVIYO513d

`pragma protect end_protected
