// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
iKKX/BZJX08ZVnmdtSRgfWooUbetI6xFTLUcQVWjV59uyecRQezej9sNgBj0jpyRsfEfhq9bnEfK
SumBtrJ0RV6wscc+JaPvyJ2H0Ri44JbkVPaun63CsqA2U96SbyGS4di2ts13J4PXq2kADmOfzNYV
1mQeDYr0YUVY0pw76iGprELlM0MKWv9+8xWh+uHgGvDNV3wGK3iDSNeZ6vkne90dnU8InZMEdxNj
f6YZcI7AbMugOpIp+R/QtBs/iGuNuNxIx1+bMFJduwnv+0U5CXSsDfe4MV6owWGs9i0etP60eBNb
SxCJoUgdVa1GqZEHdRkKKphEyg2y4jbhQovE4A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22736)
4cqn/jqCxFUQhSkxlOhPmQyxDCY1wInM5ps/HygWFzRj9hoUzPdWbTHExcJRLd7MehiQRZgw/FSR
+RKlY65gig4hk1TBu2GvulF3YIkkidNd6epnAIzm0tCx8Dibm9cXyWOPrLjvpSK3RaUZO/gQyI0H
bpT4TDix0nFRhq5tV1fXZgSeENJfAQ2kVlH2MupPYNc8604NwETep/vdpOzfvAvlzNbyNj7m3fzO
0ENUTXe0k9IpBUnyqEONeEK/q2VkqYAYehK+Pz0koPumYo4IWRVh25SoIqE98gW7tYzZt+2h4RgN
x0PESWbYYgdvUGzYnwd66J8dlDw3AZoG8GvYGmBpm4/XlsTX0RRI7j9HPCmozDLZQbx5OfXpFd0i
GB89J0wlnmEKIOS85uDYanhuBunk800bpUkSCRdEW9R0fRNimGStsH88qfD2UDVHXhJn+hapydUC
Z2OlFw5To7t6AtAW4xtbZZSjoO58I42aV9lRyg7LzW3Jo3tOD7upahs9HJpzIKHY8fCrRl9GzWjq
oHEeVJW+e0c+jVX0q3habOUKWkwWRzAxUseAnLejgasSWTYQUX5RCFQjm3k8zEJFhFJ7EueSwYEU
5eCda/dhQN0zMu5F/dA/CbPefXMB9aeHIFDeDhnQ90sR1B1I2n2Pvhr4T4sbdxreQhaEGEEZwJs/
ZR3LC02xRtm2ZDY4eaASulTChC/pe04t9ymXvLH2/p3hXeJD67b08WCEa03WOU9W/Ra+r3aMGN2u
m2SMD9JokT4f3cxlVAbgoygjqaStNxCNu4GOjMujuS6bV/vLyrdXWqCvw9hFqq2yJ56bAXOfjmtv
D/RSuRbjrNuLv5qDaITQSVWA7rJOeCAdAnpl8mgxZ9Tw8sytI8E82znri8vPVEuS7ywMQsJIB88v
D9Z60AlUuOqpuMocYsx2BQlBP1Q3YRiK0ixDT1payNqAOt4Wh8w68hXQMfL0h1NcYiy5FXqjQztp
o4ywlvjXnEBzDUgc4Ifyk8Bn/cFWqUQ535eyo0eVmuZMmfzhogiiTy3nvwn26FniIez6Zah/cxJA
KZ8Dk3hxoddIfSv2YvHr7FmNeqTByVRwPJJshJ+ZRnoGn3axlukTcODkVIONXE6N1aZe5Vm9V0MJ
NCtsUPny5am9ocLHiysbgiQTXdr0nIx8XYaiYwWjjMx9c/FXJq8I8hnU7y4PvU2ILRfqa7ISTGaT
8fh9dK8MOrPU/OToGvpJmE3jclcFZ0r01yvd3yxvq49cEhi/ekrl2mTN6ZbmtFtRiD3PA5BJejdr
VILPhi9uqFbQC1ISRjqibsh8jF6dAiGsOMAAHkkmG8a7FGPEo2FSmHYzGnaOURCB5+SK6Flw3/CD
s67Qwtu4SIXJ0p5s/5UfNm/3nOkgDelldYUhZsw1rFZ2kLOIb2Ila1D4cdMy0nnZUpv71xQF4WKs
rhM8vgQPr6W/4Zcc+xHgOWpC/C/FdqGkUttSt6+rkQad3dDOoaLKAtOB9dqrFd4VmA7ahxxc6R9e
m2KTvKqZGquZRLdQTuLCeBQoZgNaSUgS3uQ8i+z8eAJHhjbnAfc2mWlbPSgzUssCY2cSWs51c8Z0
Dia1AtTCM9GFa4Mzz7s6+5ZXImJkmB7NAoQFF2G2Nbw171bUgTJewJPHY+3fDnhctiY7gvZL7TYb
jIWnxMebzBYRqaqo52hen1HyeC+RXnE46Ch2muX0XFQWlscdXTvzTLpnBPJm4bNLxYN1pGV0ZftX
Rux5Dkr/pTdR630xOHz0kR0hHwuXMp0xciNwQH7xogxTKde8Ycqu0KW2bBTP0UxPtpNOctcbXD/1
iGx3/obGREw0D4C1gOwUfyaPlXNZL2adQWAC1L2jYaITca+muJEcItPiNYwchKWlUTn0CjQFZNuF
66R6wgNs/8gVrJeq5rtRXYHTmiOdHfN5NQWyiEVFV1Y/QPOD1eSMF4S+pwNE51dEhS1Dg8OHM+Wz
Zt4d025j7hmRZWLZBKBQan4qns419l3e/Y1ylz30bhzCUuzapTrFzdxW6l10+c8JOBC1kBSLKDL8
A8G4z6V6jwc6XKjm85v3BQVr8GpTsL/MhYL/aeABmtUBQohyFF9QxljwXgKc+wEXaCztAhfXGrpn
AojX7BoWRCgJNDUrKHJshfIKsT6LqwJrQU62jhxYRNiyqT9pk8IUgYTd6RTAZE9mo+pfCLb3PSyd
pEKqlTaf5roEjKwMi8bNiU3FUnaH7gJeDY1gWKsnpTFLoNQyJf9MW1Ve6ghU08w9Ugqn0FrQSWxB
iYrv9PFal52DWQlhp+OuwAGNewCE/9kGZRw0SISLEaMjhewaDzRVNEO8iAtD2N/pSPT9xMIdsJ8N
8k/7S+pn3eXyCL8DMcJmWDo/sk5C1AiolxK5QHJRBlopCnxDyhYy5pc8dI7wJ469ZqlKOUAiIc8z
lHgbyV3s+ULQpY7SlWjFFuEJFpTIKF4/5d594kkXZH28yMfLQOgz6ffwHpE/YyQ2w3aWYeSdGpxx
JJiPbuCCjfXt9Nn6zAOCOO6QhWAwXxXQU+b14jaZMg/sozDiCTzCZN1fmoE12tT6ETMhcSBZSB5F
rC/fkMGltLIdF1+CEPfxQnOOHucnr0uzSQ6h0cw/RryfUGuMh7aKPLACzmsrcVkRkpg2qmJBk1qG
BnwLCdUl10ik+5qbOGg03uU+f8BXa3g8D1uFf/5HDBYyaIB8mvHusNB7yGq8GVfHV+nsC93CtjEu
1oR8E2O1rsTv30fRNP0YPGHark/qVP3zLwB2sJfRadcg7UxMuMETAADbw0YzaDfGMWszIjaUw08M
tU/yfc0ERuorFv+biEO/Kg4FRmF/QL/VyHLdJ1h1svROGB8f22IrcDxdgZeEgZGuEfP1MD244bLL
XbfoLOvUxYmkeUPZUn82f051lXfYeHNMkqQQGK5aRXEGW8oNCMJ+ZujswOjCMFNeTbUm9TIb+ElI
PgrCxVcirPT3bsdj+xNaCWQgWxDmtEITOhEtXLVglQxkTaVgyDty8jMk8ZWba10kkr8dekVs0h2Q
iU53Dmt8w3sY7ImM9Qfgtt5zfhldwyNmeOM/3XN4PksSzcAMH8PA6h/nTMzg5XpKhO0A60NPoM+m
aRhYxeDLcYC4owuprTmDSgi5lMCQ+3kHcopu2FGlX2u1fqgwARTDsCjmQwzA4vSmgwwf3cVnRvZ2
Qblz80sTGA/EOcHiPU53LccrLsN6YCb3ZOc5SO4t9HstW8y3BG+Eww/b3LptM9mwig+7fP82N4UZ
0/CDLoyfyQnxFTM9szwyxE4TA7NsFh+3Zp34izYRtW0Lcw6cWz/dKCoYQAcRnxKmfnOPkuiJYQuo
YaigK807wW4mHMP5Zp7pXYnmh/7JFBMl1gcptoWZxzXBmhEBbjD0LCYemYHENvydTN686mUWJj8k
7E+jG2xpmhtOcQlNg3Jd8ONUpXlfI4O3lKJFuJvf+bVT65bGHWmltdmQeUU5RGHE6I+ZnpKJh4mn
iI12ujaZlR7DrbLfsKSd/gygWJsDMfLjNNPFahDPamRE3OVFVsUY6iDDo0bYtH/SgfzgoAVvVbaq
HE+5x7FFKl5dF7jA4QvBG9l8lRCUURH3le2iK4+MmJs9YDuBwdMNuxB0RYbd9+IIdGU/yQraoqOZ
HZ/+ToLiSa4WN9zJbJjFeOWycDT1B/+BX8x2hSoB7/5i3NztWT91IwwVWH21aMN5By5FIy5Rv6Oy
RvqBLOAoPEkZnWKaK2t/rZEc8WBrZGpFsD1n6GsjOf3EPOZdmu0zUTEG3L7eL79PYwjJYdeILhno
wK/s7DACGd2Crx/erAWAKYDw97yyCGDDcZ0icVsCGDIAanEigwKeeuVosX9664p6VDiV1nbHt9Ab
sxVTS0bTdzqarXlmShJgnOKfvMeVcuR+XJOv/vBb8g99a38xrugEOdXfJKSG4vbJqNMachW5XSkP
+rsPWlEE/Ukflel4HIrGGvHin2PYObYvll8QSo3trhLsqvytBAIhdqNcnRvHOfttmqQ49o0QOQKJ
BW7KeOsh6TxXCvL4Az4amO/Gg2NUsTiIUExQ24S7tpYa0dgTT+H+Am7o+QILNkTm9GGnd/j9o3rn
X6hD4mPhuw+97G1N1w67qpIsCI2kw2VMcyIp+i0ZRglcrNBv+KXatw+z10RD2Jsj6GY/7MHa6lTh
mNMfMkNMltRjsb75FomB8lv3BGSIsYfw+BdiySc7xkOHQoQLewk1+vAxHjeNmiH03DWErHEVCokw
fmR0Bwrfgj6iXH7sGrF21IsjgJeWr3P/YHcp1jonWk0aWIktZaXAhwX5bd2F2fBFSADcIyve1/xr
A5R6zwQiEmWnW44KRLZQf6WQXXRHuBE/LctnkOOSjVBPimCMiUHWjVe7kN33SyuYvvVv7gjP03kd
l6ACkTe7ylE33rr2o4ZUEMV5J5LeI65vA1pVGSfpEmmOKi3r8ZBrDW40MdvGzSie3hBQbVZZeOt5
4FZCdm3pFwCCQmVWJh/1UVHcj23HJn58JrkOrX7OMRA+l7HIV4raSfqpB6+eUOlux+DrfuFlZx9S
0xvGw0h6/fkhlMyANsO5ZWi+PhwQaNuFgKjnklYPfxN5qeAz4lJ7VsU/vzK5uNj3kDLU6GvP82Ge
l5KvxAsBtgn45R/CvOqPJu4wPalXOOgwKGZFowiWZZ6dxXjhdejhlsHHKbrli1CEDKfPn5eL+ELV
FRRXuelHIYNCdNvlsXRGpwLWenzpRcQIHI1PS9N9kyLfx1L5ZZuJU1DQWbI5CNk/TkyNY+GRMHE7
KHw5WxbQbCdjB2tIuZv7CslfSDWFG1PnOTAVtAifYTwygaUfxxERZuB8plL/IRfIzhQpU1gfOVgK
U++DqZbvVbx4OMSBc6wetE+9mTldg1s8G/KjpmLM3VkBeDYz+gU+qvLLfh7zTDZGhtS7k0AddeqN
7t1iRUe8D6LIFmEZh9E3DgOlGpYlca/TVBblXxTuPGCV6o3v5ZPDcvLpz4i7WgCskAsMlwUtATAG
wlfk0HSp+BgCallGYC5VdqHMelkxjnpaYZ99ZAf5/PRKUz2IHDqTeF4v4ut7djcG5+c4l+VGCyFH
mJ0qgEopj251NcdQq4DvQcwBf8qg1tY2RvPNZPBiPm+3Wmi+F4NaSLbEiMo1F0YsrL5w21keUwBT
Fis8yyssggMx5S4a8Z9IihFOnH2paENDQPV42JL5Ac196ah8xdSPAYQfz3nP6zNBUeHQA6X2Y0+X
kO+7tYsu4MnpsP3Q07APdBas20S5g4JaRdJanKUMwKqFw8hX+YCdWmUTjlNs9kZABip00DuF8X5s
CfIVkYj296qDyF7SswJNgmUaP6toJGHcwig4WxMVhpyQPqj48npU/aJxLYwPuGfylKgSIkS+uJ2o
QVlJRwbUXDeEbT2eLUAf7eKIOWLcJoM0Zbvxl1aMbRdK4YuQMqgPSjvUc/dDyF4+dfMvmdDVsoTj
AnXJrFGYXH8D9YWn3KZapLryOWzNkL1MSTKF0z05b2EOPkwrK3OkeA2j2dPQqBC2rUwkOcrriWh5
iNiRPU67X0q0OSJXY4Utmn+cL6ZBt3szkoQpfmFVC3WuAQJqJH4piVb7Nbl1U9cW1d7Nw2mrG/g6
wQEjIVnC2+AyyisvOxfn+YuHz8+giAqVHtkOqH2GFEZz6Ss6mC0U8Bf/kZ+30aW2uqzDu0PNmJET
0DkLk2e+iLvlH38+6RGwYkxSlu8daovshoCfBVuNESE0rqHtGHHcIW9BBTiYc8ZiyrwQsgHccMHP
1ZJ4A2dD49fjmjytwYtSL7fH4X9q4KI6f1b/MlNpIIc1s15oEC+zTdj6ea5ZezB5At9vTEFtWY85
6Sg7NLKHkd4FFjNYv58K3CbUOodo66xxG3CmhqpvwekIwKEjD9MTWDO4GKVGqYvjGeHUU5hzJw/Z
BYdA+kvKlcpwp5KmzfiaB6nnV62dxUHO1gt4nJkv2R8icgqa/d8YobvBBl2SE8VkGquFeMWHZwDd
RQJp12vh4L7MfGWrW8kvd9D/I2IiBriJJM6bi6/d/uGHUeZ+NSXUz+p5u1StrcTsbCljExCPDZ5o
RFxOcNOw+2RcVcyqurJ1T5FHOdhYF57gl6CHwtGO9e0B+Z2AhHpTDZPOsBE4spX0OeugywgcKb0O
FhkRNrpdha10CxDuknkly/gXMLx8LVH07vhyEfS9tcS/gvPp/tSILORRhVHPNpX7u7qOvgHh+uMh
lMa31UPusY+ZqLAcGDm3jvxe+/8mIm7axG8HwODRkGMUi3u9NE/teZ6xYTI5AxtNVkym+Y+FPbGh
HDsrjqIETcp1FbWwYS0E+h5HYa9qY5ZWlW+NGZZSnXSBJUOzT5OIeB3eams38uy26iH6N+dLdjbX
Po4kNZ91bcjSnaq+0g3lYhNpD2lteDil2UU9EFeTX9HNLreYvH/0dwvYUMHtG2wSBeTmRr/mImWW
5xu0w+CwruWPoDgo5pRHAHz7SVEqYDIaw2ucWXUtSDVuAt3VINe+UW2RBYWuLQ+oCti2VW0kQind
WA7Vp3Q/GujdRV4GKWm8uGh8PP0kPtjpSZBAhGs+m8r1wXvP1P4ARG41wfA7zscrkyM7bDAW6Ar6
yBmGhBGbNxwFD0fNadHEZangwzK4IEEZ5hdp/LFEag1S2NigYrYKi1kalxpTKW7NYZjUZ0prNcDf
gT1zawMV70Q/AFtpJxFP19ZtVYdIyEakQe44UmNhConCSqTu8ntfN8DEtgEC4rgPj0wZwiQxvO6w
1Kq4vHDLjPtpGst9TqTE4/rmB4lfe0RvB+qfr49u7ohiYXQDddI67j+uJzlWct5WERQkWEzU89+K
7xTd4WfCR3eH13ZtAVNMwv07JHAHnGbNAjzIp/hsR8i6sYwEhIu9gFS0EbyVTZdzcmiOyrQymzF3
ZeJFbMnn1aiLpM4lPnKMyt+k92o8KW77LLhd1gjeTkHRWKNn8N9NA3b53Mj1fTEQMyn2ksm4i1NL
oR9UCCChtrCIuZ6AyDvQRaH7CEc3Lz5MpSpiyMV1o2GPqzQKw+KBkBaLpTuEd52XQ5OCNIytBV/o
6oLCGSjgGHA4JD+qYWL8d+6aIiLWdVm+ytl8SiPdmz9Pa4WlMjp6wS0b4NnhXsz1y+00IbjOS8sj
rOMGbZamqjd6pwZ7uTabodgfOmnaumM16Jxs/TsZLyZyerpDA1E7idbdhF9JgcxZSqOIhgV01HRd
BANW7JMdTmSeTbx/3St3duJKYRqSe7H96iGJGAltL9fzpjTrdad5YZYnUOKP/tgrSgLkP4qrNJWh
WwF5OL9fF15Bv/miBn2QCiBIJTemwL027BuaM/1skO6iQwEFXr8nJVQZNWgmwnhdRwMxKyxcCqlZ
+L+Z5/PMVUGrC0BuOOw2kr8ZvignoVSkX5pKcpUDh49TtZlOSyOGltJarEo51VbTTQHAGqh35tP8
FWdh1zvb/QWZAlSZ//tQWy/tc9kxlyAiW8BbAntNFrXucpb2QxXygH4LZlNC0avtLU6QEyy1q7cs
Pjn16wkFl7pEEG41gL4JbotlfGskG30x297rZhSSLx29f+zx0KEK8CW7gJXY9+bX9cRVhKrTZGt/
RwMuLI7I5Gp5QSaVsJrdZaY+dY9Qrq/M1BRMhsF+6tkLD3QNvDF2Tn3VveQ56i6dhWURQbLkChgd
gWQxMs+M7lhga4VzkqCpZEgWo6ERvz/hyo8hrwcu6C90ML2CQIyu7MqHD4nmDNKbCBEbLi0EEMlP
jgIziSZTUuCm0jagC47BHYgcDSIrWN4Q7HShA0LbNmuCEFxQGhcRZXqd+IemunLEwafdyVkKVkaO
rvwkSh8mj+S99OyHAG8FFe97ksXvW/TMzGdiYRWTcScob2QtawSqoWpTzxqC3yIwsDSnbG7Vljfe
zRFIT5uhw0xe+wVpdN+5ZQTp5O3AK34X5mP9IsCKX6U0ouj3VH4tMTDIOI4uSIE5j14y2la/Jd7I
KpohB+oZqnP+yZhbtRvasV+UQo0DI+Kgd8bVgiS7CxN65w9mRSN5Rf4d7BB4Qg8wY1VLF219t7VP
Gf5tsxzUKdX+iUdfUcGwVUB0ZBFp3+1Y+ivnCl1ER0EgQoD54QPB1mhMmPsqYYVVIVeYIfHW7Cat
/YeoDP0DfKzExJ2QOle9l+GuYmrIuhI8Jm5H1o+z6Z/czXRi3CI/ngGvTqrhu9Ses1fYELQpdqsx
3JCRfhAOZq3DBetDAfI5dpRO07sTxx4c8KWx5MfBb2n6wuX3kyT55sDlJjYLZJl4bhLmZSJbRfT9
p7Jy624oLr8AZdazcWS1M8QRn8MNLqIb1WdOp+eTSaOimPdIIhgKCPwdBLNS/FR8irFGVIAzU4e9
Xf2MFfmQSrmV9KP6txL9da1AlEde2d2anHuhUr2U9VCt0ZUzGKVVxGFq+PYzMb6RikF/B19fPSVK
EUUjo2NB+YFWAoRGAVeQkJMycoN6YmCgvWeKrvMj5EUfQ8zETxmlikBcFIqqwkNq9QKYMQE2fzxO
5N2VZWC3bMQNtx5OzdkUvePXN2/HY/Y9VjXKf8d26QqGG14ZUy9qN3y56LNeXg+iyh7ZMjtK1GkU
TQ/eWE7NtL13uffNiDcpgh2KmiBw2cTW+RYuQXmNJ04GSTziY0F7qM6nrvCWC3liwjTVQgiw3uYc
D43lEI1q261/R4kl9M8Ye3wTdI9HOvDZtF3a5ofTHamS+OYmA+HqNpoK/JabLoPwqQJl9zIYAnyS
j4vyEAL4lzmjAg6TCrRN0O/he2G/wnrnVVLrzgBLdzoEKOLFmyyS/1x8tjlgDhfN0/QuAdnfnQyV
prLpTtE0cxYxhlir2MOeQOG4JNo0U3FfItkBrIxkJEwcEo5v54+SLSBc08PQFzw43gVOmV3B650D
8sDd8biSdjUqLcB7u11lTQYPdFKiUOH3+BtU8UgT+Nhwe3bTcey5Xo7N2Sj0TIuCeykcwxxnCW20
EoluJp1NpfuJhRofoYVDTpW8rpPg2qR82ppwEl6OZHe2PECYRImSF76sBvvRZ43fP9UaiIcr5jch
B9dO/2Sdj8Lbx3+0qVyJTD0Cuv1PQc3bmrIRwIt6dPVmzM3gB5C/l23JHy+Jn7bYQLRYKzPSf2SL
LEs/5PxicCQc94ZM+MDAQrsiMPRkFJEfmxVIJ8H2xbT6j/xTZyR2qHaeuzF4LvwRdbQjq6uEwz6s
WucTDEwoWGBIHaHnXucDu4alJpC81nRK3HKV07tBm635njYbPR19xByWtBdrStDu2lPqcBemvDqh
iwM6tzcDyWtf2DqkRZas10SaRa5L/BhX+oJGM+h07SN/gsPJX1ak7jhq+fewWkKcg91ngmdvywJ7
xPM8pnd6+WpuAHM6s7oHkK1T4Qu5AUwB8w1vB3xBzwM287b2riKPD/wybnayq6Hxn+qMydQbCwRr
p7VFas3Kg2dSwv49F18+O+CpF58O8GNTMk8dZ3XX/s3Gdn4nFerof1k73FnvcVFCp6APsQAxwIJW
mf/j3r6I9LYT5oAjqUAn7QsLT7VeEqG3lPWnNMM8dOB/x6X3JuD2nr0deVNx0lUaB8yLipSxLk23
ev2x55WOJPMmPknVgihXS0Z796bGFUnfzWlbb7AyB/sAsrAgCcYE2hqGS5c6fWuZlREF0X5MqeMm
GQN8ZkrcsH8Ynyp/UukLzWOe/E7OOia3Nsx3dVlKmYdj6m2bNX265bvstng96XAfEqGelYlonXN0
6EqH6yJHZXj02PcUr2rO77PVYM+MlcjIIPvLc634XFd4YdSg+3F8mVU72Gfqoy7JrsUN+Dsx8q9w
8mZJojGXmmYkC3xoqyv1KI/tMQPIdLle97GlQOSj6AGop/fu0EHhmIxdqvEy+89J5hAvo9wnl0Eb
Eg47eAzaV23WuL4cY7ZL3udvvvoHbHltp3komkjanXkjgn+nMIvXY5LjMJtRPLKm/DDlqWdeX2rZ
7jb/Nxfhnf5EniBpaZZFbNGrNDAUyplxZ+DtTvtdaJ8A4F27Mv7O8pqFAKAF5b2EbkpUe2Z2Mq/X
0SCRJWa+p5VVv6h+++TKywsptquLn2uXFJjYbJScd6s5i+00xB4mgucHamLZt1mvQk2vRsBs6qYD
VOvzMEABQNRt/p9TfnlMIoQTQPmw5ijGOFy+5Nd70u0+eDIHwKBKncYdYEZdnREF7JWiXRedLgJ0
MUuofYeIbkV83DVmJWqF1XeFTmPRKfeyGxaCyDkWdUDGf3GJGJcr+gGD8meNd5dPSJr4Co9NzLag
VnVZsTL9z/ZaNtUmwaeVeP8H4x/cvyxRvpHgzYay7IXIS25Bx+t7wM5afs2HryKtBGbRG9sOXrWL
CuoTs/VUBt3rHgWom6c4JJ/jR9I2/H634cKwY6sOdswAVmLCbNEFDDFk7L87OowA/oUEc0/o9pYT
I2rD8m7eDxB1wf/9aTIp1MOshFBr3i3x3/NXwAjNuZsh1JbM5Uc7AXHXlgw7QgVSmF2oDYM1sLgL
acUYk8ZTaPAzXE24eLr/LXrYVsNkOfz9Yleaw3wTWjkwwJWOYy+kvXuTsgJVQEL3y/DdLM4gJOnQ
5lM4qBl4nRqcbJmwT1GnTJM4lOCc4CeQVbh3sA3XKFrN2laTYDeasJhb0r0J4sbY0zvr9lWnKY03
qisAAwwImO4/J9hHo3f9q2qOgx51yvfNhj07vbW+Jez8fpK3XuS9gDsGOxu5VM1BOkJZSCVyYyrd
a+ZIo+/zgDfpzLVa6x0s80NCP+M9dECLQ+k9bmvH0qTrke0YZO8pklFEUkzI6UNeE9BqaJfOjcYU
aimxL+f84kWLDRiWT4RsRiPHTrqw73Wyz/U+pFP6KIY80vgEt+jKBgq5nbD0ZBzTq36eWIcF30Qp
6AHRnVy5/qZRK/baIKJrFd2+nksxoKUht/shksy7O6J5zK1avPa/tDXJcyN/XK9AGF/M6ng0YiwZ
CTM3oYCUfhQC/SSDOnvulbur7xaTrGIZqEGJ7a+lNfoeKlg8sl51kKLifZF05iBZFzDsVnChzz6w
pQjiIODSezO2DpGwXcgc5SUJYQABtZ2LSwW6P1EQssz/A0CTJelcClpUgyjL8JzN5stqgVFhH0oR
LlNMfFCJH1yQOtHFIeuZHlQrPZL4VS7zsoyPx7qLw26f4LeXZ1QcM4GAgz2KcdSTtCBud6muFrib
dTabevGAQJoMNXduyKdPm4HwkFN44gohAXufNQdu6Yc1mgn5OdrKl6xFYywHI5hrZrYVg4ILWgu1
gmTsUSJPKiBaM+R+KmgPU7Nx8yHtRoqfbrTZCoa3GbkrxQ/a+gBqK89W5CtLGnZkOpecR/KzxY7M
fp9ZtyIyggR5pNYWC+yPzyGDqhWcmNdzI/qHg3TmlxWz4GOteHmdir32obUyv0A2cu+13NIkUQfQ
u/4U2eKejHvGO5yRTNzVipmD6FePAc/wwKOnZmes12UkddW16UNyP941aHubwoXuGTv9+1ozhXL7
xX7avolOuFyysjabtXZOhQozIEWxabiLlRMKsRd7D2PJnhiaH4qlF0gRlRNmyrGg1PTFvxVfpIqO
gNzd4iaFO5wUz0ZLel5qL3ER9t58873ZRsmEqskR4T/FhTdBho5grt9S1Pc6oGsTBqvLDVye/xom
qnv0LNs85N6jTwK/4A3HkLPkLaTn9/x3Bn9/XzO4CasEf4ihzmQDmybwOWHfPznTl4J2NtSkKmVP
c9K9NBuZdpqGWTHRlDbzGYC/pq4wrUKbL/oeIjgWLOK1hqmjAvYEvIWxQkjQs4yYpuZHUTmCn9Ma
opRDDeoeEna0BxaIwg6hrnhm3PTIHdZQ0W37oGA80ETJpi+G7GJV+E4Vp/O9kUc+1gDlM8GlvAfF
oCNShBY50sPFxuXLmfup2UydygitJ2ENghaJa8VZHNfhGTz39d5pN/EIsjLaDDnxkloHHDK99g9Z
65Dkf1i1PGwxBknmzwQiMBmv6shwtnW/MCH+bFIIz3tttxkkcdO2OPu2qutCGFdrhiEWF17EoUAG
D5POYLcr8Yu8ftj75WBmGMYXIR/HAHfsxQ+IbEDrd/BEXwJNob3frQtIWUHwl1sUcdHAG1RMD546
cnpspQF4BTUWndL8VJKbAuRiOD9SeqNFnUBJuHEamAROYH9W/PxjIW1ZMOXMxx7y/4Ee+MWNxz8n
w854ghf3E0EzfWo1OOZtU0NDjMeNZ4AaBjHSvvEhtaA1q1/oFx1MrQAzYUvX0H4aNJNwo9bn6zeP
KQwsLvWEULlplViYxbMgjAGoHtntwIfV8L/MdYuSy6sFjgk60Z48hoNrzHIiXXsvQw3f2OwYGKNj
mZ+zl4ZcJxRwUjmuAxIo1PWYmKm5UEodaN5jH0QcDLVO8YQifhueUe7YhbvrzYbARE2bzyZyS7TG
kidjXyyeF2e5kY22jyejBEWUjeezHkqjo70GdN6embc9CugCWaLJ8zevKzBJL0YuOlcZZaOAyXaV
epjCmmUZf7RzvlznD8kMdf3BopRgm/5ttX+gQiErgpl1u8p8dD4pNAUDTZ7QXouA9BtjPuOPhspw
KR46jsPvdqdEvr6O04teJS2yVuC+HMvQfKdfKB9y8l7RVUmoUQQ2F5OO/n8jl36Vxsznn6o4FDvB
IUSPpeDzDdWwDlHReM0jU4IzRKNKYA/wQ7YzWdB5ZwvBV9RL7kyBeGQriLx9ZoJLoe675F57F6Iq
Egii0hdeR5J8WWHahJE0emXzlU1kXYxwnw4X+Pf+lr14OC1C+2tU9LfSEwU1WTEUNCaxPnNgwkIY
DAi5Ltsa752oxN+rm0r9ZeC+fzWFwR46/hugn0SBAVH8ZKZnLXvq/I1fCzRU2gcD1FicedDqsQ70
07Ag3wxipGz1Htq8StNjSZJsT377Mh2lyjOzXmjeh37dk+kzA5RmmDQsnlR6oWJbQ/4CXoMMDYDp
nZculG58tjlyAcAtqBe0tppKv7lp3NvnN69LaY8Xg7q/oelkqgMg4HgE6XjzvFBUBur1MQHYZqik
W1ATfgq9MKRMtLDJ2Ju8ttPAmGTjzoQws7dTIggfxuI3rQNoxOAZ6q9QWTnnpQMyMyzypm/39Mmc
GMHWTYxg9KIyOS08IZD1T3JZdOYuBqdlG5sWNI0LYu/KXsmUDjrk2D2ycJz2XucZxSXxxYtW3dIe
ppIPzLZ5rHuBYAOMCqX34wb35TrtSY22huzVxrH9pOXd7mOm9XwW8yw6exSH3ClSwZzhETmjpFWc
/YoIjIwc8xG4AhQz/gwrMwC2p1jtoTtj86/PfOOp6W7xU84hZR8efs8OC6GLhtAANcnMt1EY5h+K
S4lhlps2vWmJjZ5AW4eSiXNF2k5oJTZNWBruafhMfoBCRVPO4w+gMwXoplMH+1EwGzZSFykAENA7
S50sy/l6m5ObdMFlB1YcayS7ydDeKEYzBjE9WfCAQXWsoZdKqTBHLDZPj3G5kRkbzA3cbS7KxsTc
c/Tm9fVlxXXyIs/jaUMvG1/peKxzy7136eVl0IjN3b6XKSnYAPZyXYzBS6J48q+mcwlLzIgEDeVK
bBzzCPF9hRikDuHVxp/+iTIR13+uZ1rkHpPMmxXG9mgExyQmWnq0v4ZTbvaG5yV1bS88d9aK8pHF
wRqF4dzR+L/4CvB+etSGMelPhaUmKCcCqDpIg3pwVyUWlxmVZTF4MYqn21tPJkia1d5gsBj+2D6c
sk2mUO5ib5d1Z5MZD7FleHxutYOvSq1TXN80vlmn5h+kl1rvV8u1kNSPRBXHv4/4MxbckvTbrcpI
JAtTdHIh4tgGtkBcIWySLQXHQMr1zgKEXDEEzGHx27eQvsaghFx1Da2Hw4iJcfZJYKpvbOEA4+rm
K5pverfW/Ik1BR7isHDyP+lQ/kMCDWhsgehwgf3mtCjqDG+wnLMfoWAF2kfx1XCqjMWWttbGjmGb
DLdICJIFwddznjt6UdAiOcA6De0MvVUVIODLbcsHrZBphx62jqQGQ5a40yXEzkv1vhriDAWaHqPh
JfvulbhvxWNKmOS/I8jkHBCO+cZcsiXcrB5nwdJMLyq0GB/6CptWJ1Cr8lmMq753YIoj/PklPetj
wi3rRJxzoDH3o/BRyfejomZJ+fRoLNG3X6NZa5sMRTmma+V2wW78yLxnykWK/nR+jBXMD7+O+/RV
nSrKrpQv0gCNXyChPv9+IU3tfHlY5Gtum4VtXrFQvtFCTAE6MnG+tPbnGXgneOzyHMk3QLB3O8Km
pomhQ+eT8RPYI+keTIPQlOXgkeFvEsg+XlIbVJ71h1M3PF1I9Ewz3+XB+nN2nVbyi3gx3RbrcGio
+UDn9JlQIyRXJ+wli8TD2O1MN1I2kJx2gO539oAIV31cxWih25I9ynvbblnT46sT/b8SlMszBpcW
MoX8EHpY2Jd9xif/KZ/1OiOifLd/aL6o8LZN44OTAUx+A7eFo96OjxVJ3IvaVnDoQegrK8M2oYtK
56nohGS48mZq+41bptWoH0aj2hzzQBByM9POWmclOHmrYGfovKB6QmWF/+TuIYz0jWSF3ggEjP7p
HTIzQBv0wdnhHq4Go4+NFeOpQhZ+yYUT9m8iC7DoJ0pZFYkK/2GR/IXiBoW5fj/lCuOnO2nysTp4
7zylzxMwlBd9jYo5pWvtYewm+1oGZ7Eig4QXWHtfzrbuIp75ALRue6haxZGOQYtCOyHVj/6J3Vd2
1noAjWwhbEJ38YvEEBxeS1MMHN/1gBxO9aMKVTftiZQcTdzqTJj6ckPkXtP7XBMTe10N1bYZzivI
tATEugRhxksSUquG0HMniAjpmlnpyAHgiRwwusjNn/eqb2osgDSwOdULRH7JOB/UTMC01WYB7cKv
2u86dcEI1DLzA8VsWMamR+B0yceQ13tBuOOQFPMhyuL4xrtEF91I1kVXXuXHail3D2gR/vS6eXOk
Hzg6pgT1XwIaLYScCLUa3eJjrxVjjDcSy5k6RE/QrRlV+uia/QpZ67EdhvL7VZHnCSPt7RpNb4ZN
8jzo/TOPBhEq85UuUJQUZJG2XvmSSIiFivTYsFitBnL78lzd2k2wNIj7EXEHq9EYWlyxHGUOWE5y
vGyNiHwFcx/gfNwi5V33/+piMmjGWm6PT+T3jjiTTWDmqXnS7e5S63ukz10/49Dgr0bsOTaUej9u
C/YwVb/M765P0YFjtXVqNrKi31CnV9Si4wvRuI8WhfhJFXqur0wRLQuKpvY1aoGOIWT66xJamwLH
N5lmI/tb2hEuq+DnxZ1Qe22SUjVawgF5GmhiGolL7WqTmxOIJNrIMyNMHYeaX8bU5i4Cp4KMV5wV
HKCtZUAlWRQgJHKskryym4kz5i58eBwx4gSL8adDsEhlOAMB78UD3Nif6KzDWAG2QDaVtHYYuvuA
Wwkj5TMnNfcJETxVU8AqhiGaogDK19x6pEUzJ/SlZV4AkqSMqzINhCqUc/BT4qi9yFxOpDx8Iild
KUHu3A2FEwt27vMEs8fWjp2Oz9h9E5KCtqacPvXuiEccm9pWJYlr/y8Ndpx2+xSP+w1LP8Jw9vo8
7IB2mgpOIsL3alWabt9avN58j+SaGBrrJKvPZmQN62BHG6/x+0il0Om6Xc+kkHRMv1X5Aub0lKo2
k/HDu2fHtkJk5gtVcuDzCdPm2kVMcCGYimLt1TrpOdVPOutscGvXF+0ok2HA92UMgKyF0Xaew6+s
Bx9UqHu5lrGuVYEwsGyE04g5gSdVsMNrlwbe5Zfg+0WshYyVFBV4s4VTluQHHy50cN/T30yzz15d
WsmyDDtNeZeXCNPOvu/gpJnS56RJDHeTktWdrp4+U6keuNlaAYbzfUZDuYDMiOpYZMTSmTkIorVj
il13FuG16Fpqt9cRt9Kv3yyuTpRkuDCz6htvu/EhPer2E0QKWu3lyamqc5NLaCm7HijkDRGKC7LO
sq1mkfccZLYUEyoCIRKsGXGTl9I5Tgx94XO3Mdi2Q5ec+4afflheEK9huyT9DwNl/f5D3LNKDim0
t9nDkNIIg0GAiO744hyg0CWlnPPfPCIPLdMM+6+QozlIjhWUzbzNsgQeiL7mVxu3lH07HVpGZQ2N
nq27HsFsqyFfVfCPfc87Ru/JMAGT8Eh8WDw5xjGcyMuui1hN+3bORQ+3wEgLU/5oZECsrFuRVB5Q
Tram3mQAUA7xsmsvTuBT2NyezAA9rb2kWwIzDfhd+I2yh/DI3V0Rxhc0Hl322ao+sYrfA7tlp7Pn
Q1RiiEb8EL/Q/8yRAGQCNwsP5dpkOLRiyQKsMUt94j3Ad42bKqaZJOfJsE1YU295S/SI/rkL5Ax7
Ru4nVzGwCJXn1aG+aWcnBsOmsQTSFI+hvru/4Msjc1QLpJJuFE+oC1h4PPcePxqrTHcHFdrD/EYO
wTpKh99SDwNgKCr1jy8wpnKEMOXtNO6qssIb/fnXhtf5ItqWt2/Ofrr2TvS72ICJsrnHDffOnIIC
Zu3LVmGqaqibnUI/hRzdPBdcdDCL8p0MxL+paKASNqUuJzwEsOGDZOCO4ke2XdFYG9gvqHm/0Gka
6twxKjvWRs2vlxmtkdVv16o/mK3vpXo4AWDQGSP5i+rfhhiDWGE0sHNtKq3UZwlZHeH7FCqRql78
YcyMXGR7zmBI50kSM7a1sGKnGpyJZmTW8hrQOG+ubY7YPRJjiCy920jcw2Mvfs9aXWW4a3x61hMC
ysAn0rPb/J9/5yTJrfUBW7VQJ5yhuj8zWL5aZrO6kfpFdw630oNvy+Drqh/ewdWjDCw/iELTaY5U
T1I8EiWfdGFj8fH50MeAEiUMx7Gqi+Bvn+KKJlwfewVfHLV99bqKjZgaCjcew++5rmZ2s87RQhoH
/VXT8Bpg6vbJM/xV44Jc0hgY5aRDVaWAy3mliQtPWp9fcb/XBAtefeGwLT5f3Q7LjvKEh65MJ0bO
XN0YCn83bVU1px1zjVyhAJ3y1kH7j303SbCaMpZmQENYm3tgasTRLQSWakfIjeRFyV5FXOx8JWdq
Dtxw3Y3qBcuNu3R1xXaZnmYyZVtnDMD2BsmKXR9Fy1HG8ZPQ3fVTdmJ561Kl308cIGrOG6C6vt2/
gv6fSbX4EdmbwQi8AtXXeYOdcTKhN5LHdc8SfOEEzpDhtHG17TRvWX2p3MdywEddmlxs1HtmV9x3
iApe1WvzAm2cuE0B4R4uWtmW61/oKAnG6K4r2OWa01LcxKmtIb5i/991JRW5QZd3R+Sak+0PuiOh
TrFHMs9a22IfcgRYXcApgdC4LciLcTXbLeRPZ6MMiOCJwYtFj6zZqYdjdF04JXd3vGqrPvmlWamc
13B7wkhw1AYLMq7E8ySibI4Q4TKnCiH89w0z4dZNeO+oPLA31JSvWdhZwNpOIOoFKVlSd5Qoeddb
BHmMDAB8PNpw23/NJDKvuXQtFsSCgoxxia651MnKzu6X8y3k1u7qPTMWOlZ8oKGVH9l8fkbE/P0N
gTABP0TehtmjCPlaHYbGKcLJpYzuuD2K1bk88bmjTLdYdeHCGwcvSiZ0Jbx85XupnSsQUTk6ti9B
7a/AbcZ+UsCxnD2GpLEsUFLlWh+wWTpfEtUDvntPi68tLG9IA/e6WuM900weP9glJOruHbuZHT3H
TbkgNvwiy7trtHXR++24AQlxZQhlD9Z4TLbAjjzkSNWxifkRlDFEIdpiVRy1WTx+I4gXIasJ0KXC
U76d0vF6el4RAp+TAj7S/DYtp0BYyWJMfxcv738KByrXLXBft3zEVBO2dqVcXraMa39fI78pI6Wr
G6DvND5XCfK47sAMxesxWHNItAl/0NGKGujey4DoyTwYNTX/PssPUWmZNYnq3n2lzorN0IffKNKt
j/sdmpIiMILKaq93vSZB3bwplcvkitI3ES5WVGn0wPvT9f9I3bPd8sdHajfXJlir1kkJelXcoWpH
WAz9LD8GsdqDaV1MlSM49KwZi0OtITKTFx1IkQ08dFCLBXzan2pEAdL0YUVjJX8EqwmiRQezj/BH
Z/Il06Mab9ruo3GvYsyDyzY9Z/auo1Lb+jCbCy/b1GlBG+YXDdtr/J3fCBfq7XzxhExK8iSz3adi
YnvPsMLgGfLVPf8m+EQtRxN+2zmGc/N+p27YhnvCtaoL7IwltoCyMM8yJY480d0bKZBzxGwuDS/W
fkBcVKkCa5Q+kDVGVf22Tp5+oLwBC3sVLwhv23k1EWsAdwzn+Gdlr9nSr2GNZw0gaUm6MKoO8z/0
tWu9pROCGBKfMnt6rAqJsvhFgfiOHMe1629WjwEObanpLekTijCJ2tADBIa/mq59Mbe1Q6et8Li7
o4lMtaD1XhAm3Sm4D653POxAWfJ+vIb1GuY/Li/Zpvnjdpdh7y+/sm6we99JKybO0xizdHGAhxX2
XUnR5NiZFz7n8szcKFNqrhuFe96fNIwzRwscgtBVgYGYOxZaNXd9m2TGhkk7M5gNkHisbh0v8nLo
UmH7N39KpIcFHNWIRUKx5SvDMJ6JntjMCQomo4+N2mI5od5fQPSKxMY77TZtob+xPWpcXn/IAIbZ
BK1tIv9YYWISLqeVkTpw7THsST5Vw4F5J05QRQpOGMPuGdfIIgFFl4K/l7aCqVNUJCpQSAyiiHC4
3MWCWMrs3Xz/c87x++mfNzndT4ENTAKcApvp9tZKyduytN5y/n/xAzlIhH/Xbunz1Jb+dSiJ//1M
sGK9DRBUdcbsbOajVfWgEkxJW3ESYvZWaysqk2vAaJQ7EIlie6YqsGrH6vtT0D6SvMuUPqj7qT3x
0h1CQ4neKEDTD26ovOznDdXMKDcPOaGmHhbXoJoleAZO4nwJEw4QkOOqfYD3TX3bVPZhifrtp4OK
3udW/qlc6i9wK6ZtC+K2mAW/Jrv9pHXwzxeOulRdFlIfVOoPYOy7hR6LXwlUfYPgREkdhgDoDKZc
2s1bpHl//7sZqdUt8n9CieoBHvNqENEZqqKIgt8bj/1dTYqaFcgx7wbwz1JVE3xfF6SSlJccIV0N
W02exhOfHZAkqC9WMtIlncqOtWzuQ4GLWr6c11Zdin5ogyAp22UN14StjmN10+1m4FYMWv+dcQ7c
6IE3u+c2P0tHum8b2Tv5pGgKQ2AVluoBapGCNX9100xBOmI1vMG9bccrtsqNcNcGxMvONX0RFdMU
EooEJvkGA4mSFNBeCX25bgIIBaqqYOE+dxBOMbapussFIE5QwAaJmdRghuRW93eZpbXDfOq4Ww9p
Ak/+WJeJ8ZoeJvfIYhWdrpt8iPwswFQeJCvjaYQvk+GM9lK1y0ehaHO1MEbeYDluFJO4bAOmGfwr
uw75LOq+2Gi15VNzJtHsHI3boUWMvorHevRLYVrtqm5Lt1MP3B1l0uS5BpTNri+2WC9zbBMMY+nS
vrjutewdhh7kWjgMevy+lHYf4VxiaCI+UsLlS3YlYmrM3mz0GFZIGf6oyXErkSu2IUivhqXl2sTy
uWcys+slKoQt0ScdXQsCVV3fgB30dNipTHOvWDjo+MR+wXLVwWGtvUERh9QqaCZjbRYsMDTK0I6Z
U3PXcJdqnNtKpVYwfgraAPBOvqrUiA1gq+Ehb1WtOLC3BK4Kf2+OYOBSN/ztR/mE1z9nguZ302ql
LCBW3bJsEnhYhUoLKz9azRN6clxCpM4HzlWXnx+deaNi5QG35gVo6nM01V74aknAYDYkapFzjsDK
BRuWGKaSPntd48yXLatNnTcfVg1r0D18HXCK2bnsAOIFtVznAwYWGL/GYGUDv1EFBG3wFTIAhw/N
fsg9AUXwZGKhYqD958XuMA1hAqXyDZu0E0kc4Ze84Yv82SJqhX5bkDeECyiamrVGcRsox5AEQ86Z
ymn0kt9JtRcPAR/AC2G5yZ7VxLu51aMaGrxFUDxRJ2VkkHkokgbvz7c0MuUwgpjdoi7g/NaiPumo
6paykZxp23VWp2r5z/zIbOpPgRp6atBbmvG+Xr4hH6JB/y27x/cIBy+TD2WsSL50hFxwyHz0EjyR
jArkeZHuLeOSU70q1BwtJJqAISUODukcVj80t+bu/LWNxMASxC8lRS2tJbG27Fotz0J6x/9nBYMt
NkbPvmDusIJBRGL8bcE6P3fyV5TNkACIrg9MXg5hdi4EPApEeB1jPR2gTsk0vDwgdi/Utl983ubN
s8no/xFwaP66Flk6YFsfxF8eQC28ww+x2Av8G74CTn/qmIJ3gGNAU8PusgPElD52DoWC/IuM9ShE
U+LmhTZYzeyXkT0KctbOrb83tDGQ7eB2YkBdsukVqODy0FxAu0nGKUrn2s5Khu4cNHhYWYbO7x3y
BV7xsbUHZIeSdEy0laMspX5OTCwoxCrRURZmlwqZUjzhBm4O8wFkyVPocuPUdFoWky39vBVb53ko
mU2QFJxAFQ9AUbcMG9KjUCr7KpcJK1MfRScjoB7sTuaoz1krGv2anPdygCkdMYp45ZuGKegoDTp9
d+mos6Hju8kt3LYjcDXTfxl6We537FZ7JYHUdBSWzhVzQBZyD0HxuDLGlc8a1Tht6eEHaj5xs+Q4
EADv9ZwIpLN/Uy9evcbBNGW6lbszfAQwxDBmP/PY4QbWLPZU+MTkpDwEwLuVMddhE0/uFdBEfNMa
og0q0tChOQotKfo8LXc7GPaKqD6cIIWkOUNPi+POD20PNrXCKyv3WD8U2eaYN/wEyOu3im45Pk58
5jBvAM3CDXbOPqtNTw/ZKfsv2XMvRolExIB0EUU2SBJKPpV56eP5kx9uByePPUjwODqqL6BcTFqt
QiMcmHQxxGWXN45GeWyjZkbDodfQrAziYtA+gRIBTi8ds9FISJgtCTh5bZ+rVyDwJAAOR32dhfaQ
KT33ia6je8xSRMkM6q7KdAtn7NSNrP9ykoo1yrM3hHWpw1fV7NcxpJE9CoHkE4TKZJSb/GUJSrlU
2oROTkOb1j0Cr4MZix3182KRhBkM7hLH2wTywf972hdsmaTkcF2Ht57H3EzCv7tQud8wehFrqamS
Gj1Z46VvI2Jll3YnC4QdrAgkSGnDNK8whEPA+luXCpT7zwcK6yHUj6EKYgNac2XVqxAqO755Q8l5
9JIBujvyb7rp70sbgBsDT59wUHstBD98f/aOPQpfLeHCE0UXAi8T6e8Z2LPyRr/AcO6MxWN6mXhr
CpACrwDBPRRpHNEibOBWQaKw9B4CoG9bhOqxD/WzdzoSHUbrQZmnWPb6SF26My9dc8J8cNPSSBcV
uUTQ/9vE2z8cbHmPMN5QF0hcDXZfKPMyqSykI/Mugs7EgAjiAsLfQHWzZ1pESiwm944V3P7J5f4w
aQgw7HnK/dlVHF33UcvEKKCDza8IHj+wBUKc1iVigY/tit282O+OmPlsHvuKGq76FCCQeQTYy1XV
lIfF731wBOdfD+RaCFCgsivdqdgrVzSYU7GgloZJlxsF7tmi03AwRKzmcplmh6hRoU2Hrs8guH2h
oPYhgjofGybY/KYeVNtd4xuzW/CmpdxRIQEI5F5x3aCX3F36CEheXEyacFC7LvuB5y9c+R9Lg1vy
zyeFLNe1mOC+EmKPpN+RYeSOjNW+eRk/sMtmI3DsAnitKvH5q0uU/CdfHlLyzI/MLb+qbhV9HTOn
lUGOR1xuXhFBHsLKYK95RZtz86nMBQYOu6Qa+wuHwm3vHnuvAGhUR7fYczc0iIr51tEEmyUaCjZW
Qjfu0BeU/oXou8ILpfg/5h+vLiULhum67ULGyKDfvDpck/MVVskCYq3R+EALAhmxctYO0T592GLQ
MyzAyfV1ns8mR3+wai72YKtrCEZu48siWMTm9Cm6rSI4Vq643nvuwMF1imG9aXPBy6Egwud+PPpD
EEb+Y0F9VKyAWRrSqudUgiXxmSwTdvsbx0aS1Lg3D9MpwGA1sPYpEPsTduHe4CkJuyzhozdS2/3Z
pRtA5QDhr1S/8YPwFpWczMjbaVY0/AX5VbjNxum2L0bW4l6Dl42iCglvi4XRxGXiXaO3NVSEWMy7
GM9Co3d2sBozP9VWJAxIfNxmOnegUg5mg8OoriArQ7XF2IVUlSuW9cnDEGqtxX6fnWFY38C9TMfH
RyMHXiNadLXwqgsvV8rdPAQnNugJ7RB/tC8wVVsk2w/RB7CldqhxILa3U0bCqExbvMCVytIm+lSH
ba4nkbnQPW1L52UDQFqOGi15x6Poy1yNNAAgBNpapCUVa4el2/NIrzSKK6rvNi9nH++wLYSy5Bda
y5M8bF4Zo3ryCVx/BwibKpPYdoK2+JUGVAjh3GfGhaegL3v56J9vL/zlB3VYeeEEzK2edGXXUuqU
QSXpaQlDbgI79y5KyOkNTqHnHdAaup/rWx3VC4RZUqEruStrKKSZb8KpdgndqCoUL7hz6Dj5Ncsr
NeULzorDMmKJIkEnGH9uCB+M/YPrEsjYBjdYb/36tY7FtLl4Fz7734TudmXPfjpM11uZOytP8RBc
G+1te5sfgndPySqPE+W11A+8tPoV8NxH47RllI7kvicy3DWzzyPZx5C+n+vNnmJEKQRuUwWLU54g
SuFUnReOA7Ri2s4cOSmf3TV6Qut/bywiFS+Qr6UwSP8VzesE5hWza0Tg1THYM55HcCiZUcvwB8Ss
x9dVaFjXNc2dDpMLXwD0DoJlfXuWn8mE0f8Kfn5c3phtXMkJAiGzxCfBo8b7vnc7zj2oaSPJUowr
iECvtgBgzMrkRnOymSKX6j1Asn61Wr6xKeu9rz1oQBijH87sIhlSEGofZo7YqxGHA9az5NnWBH+1
b18f3CDbEXMACNx7T3ZhmHpZu+i6l4H3sqgwLS9r/xpnxiVx2lVMC3OIts+E830Lygbr8F8CXAJh
lvEnDDN10qy5PIkgO+mX1XRRtLDlsDjv00/CPt6YQloLu8xeNP+u52j4LGy4TJBF372De11jimHc
HC81jwaaFgIxEn1pAqV71N/G99jV+St/Iizjao/x3Pu8J7uGelyGAfSsqJGXP6oidIXJAvAcqGdJ
akVYKq+UjQKTimCR18Ax5xquicNV4F4MqOrkcocu8D/auHCjX9ShqgMFuFjg6dPioMHnImIOhAb7
GEV9S2Jc9fAJfdeQUG8IV5HrK66lX8BHsg9cHkUsK94JGKEP+itmR93lZpmDAB15EePn+1zBpfI+
+dO/g52hG36sg/g2CEkRjX7DC5wPq1rBuhv0PNDybQ0RnGDOXA9TK5EgmPpLMM9jcRsebYPYyjSh
inh7tankMBvdRqzm6KltLlMXYgfyjqdOelL2ws+JhWU6KR9oAaifHl74NOb/pVcNcc0fUEQaVa1H
pjq9DT5oSVK9+pG/rsR8dUvb4lzQyRtP9puQU2Qy8CkJ+bEJFebfKH2PtJRsXrEPCOn0YakuI/L7
B6yh65dqiBICVJ2M9gWmUKZ3vHEjRI07l674uT1CFlAPS2t0SA8XJs96L7RNMnWzjPga9Tw+/on0
9E+PKMPiDJrNlWjK6ndnfGFv/CKLOnwu7V56B5LMZnT4VBruXdvCKNoltCIQSt1efNuykCV+EFsH
FTfZ1xwWV7/Ft3o9SB5KKqkxx2NtLEE3wka1tvwCVKUP+Jmdh1fEUkpEkLbTiFA7LAVbelT6MdhA
N2FNzbbrsb8opHXtDsTeLCiJhN7YUaEJFruh/aP4G3L6vKgl8E+Tn51uGnXT8Fd/bUa5nl0WrgRV
Wpe2g3x3NjUBPL841UsJF16hMzwthNuL9loyYM8Z2vIdPAQ8oELde+1ZAOCFcfUDzNTxtRk3N7EE
HD7S96/ToXopI4mxA85+2VSwZ0Y33Sm1KOA93rkAZTL7iSmvWN2opOefyGeEzSpPdqVkipVSBQuU
L7oZOGB0qK4kyPVNQh3OprqT7DXJXZrFymkuBOYdb3eFTEDSkl+t21FuGAlbz5KDTnUUEvp3A/AK
GgAvbfc3vukSdtKCIVYF9SEKgmBw3HRVXq8Bt49U3yIVqB0Onv7wFmZFp/kF8n9kaSu2BnPaMbfF
ypj2t2O/I2X0lLyfo359//JihdMrWbuDeF0/fn0ev0OWZoBbu6wdmRFzyapl+pGFBqn3+40V766F
K9u/McR6rucq+a2VkRG+mMI8Hm1j6PN8wDkSNj5VSv4D+21bFzMEXZ5nAIXRWzpMXsE6fOO7Q5Vw
vTRXp+NyfESZqipz7ORtQZOlhKeLy2JnHkVHI+G6Q1UEDirwljMag091sCkzvnFz8tSlcuNDxCE3
xSP+QnZzUNro+aVqKMcw9vyNJssjlQG+p8GC6X2q9h5ZA3jZzq4espSMi0Qqpikz+m+aMKFG2MCC
qnI5npY5EN0U87HV8M+RGVrbiyDr49WOxpfUuQUuqszRh5sIHNdrQtq2r1gWvyxp2hsWVEoWPa3v
gtP4SVLCqttLOe5pQDlqro6j80E0JtTSwl1Qavbfna3sscdBsvEJbIiVxEesJ5wldAhLYDpW67M0
nb4+d6lSoeriCM8rZnoc8lPmZOlwiNmPKsiqLF0djOnGKFrv4P9hQc3dA0vd55UYto+64QZDk2o2
2nIT2wuc5qVVfS51XnJ5SvIO38le0qkq0D0XE67P1WizbOs+odFnKPikrpbkvoMYxgu1Bnkk+krM
+lu0QUlJeAhNfKUTJ13/xz1rI2LlqsKTiaEdmwvGGx5AUQp2mXLD2eOsD4tEiVY5q/do6M587JxC
tGFeyth3mI/HSClIgedoqEr2RkZSW1zS3dVdeJHrTVNTFOrl7FZTAHNExhDia7jLLNX4b5qLX4fQ
37dz/vabux93GsEHF7PxbTmDTqPEDEnA7Z5CFSMQnaxmFUcPoX0jr+YaN3L18957VxSNMv1YJahI
vIrSLuUaiZVTJddgAKGT5KGEFs/yVUKtsSYmk2MKrcW3MCrT7w2Y352xOd+yqjCTS42BJ5iChMJ+
PoRUTTFqa6g32MHND/AN+R8Tax032o68rzoiGn1RkBnChbjkDL9tqg3l3zqJQui9C3RlRXCN5oHT
nmdRQ78Pm8o2lMODz/NNHpjyjEZp0Ws+7xQ7/mtRhz0RVw5Jfu7Z/X84HMIEBfT8E0i1qNkaTP2/
vCoHLCS2/nQMDbctSMchZht4h8qNoTMY8KRLPAOKdmcEOP/dbJN2F/vB3pCcQ2xFEYAaHKxFKMMF
Zb0zcxeLEmb+DvJcvx8eIdbH02mH8Dr9SVQYfV02QpFI9MrLn23DdWOAcLcOLh1EoyiQsiq5cyRP
Y9ltK0N/4EYsTXXEiASAn07N5mo/2E8Zdx06estFlqRyVHigWSBYDCwxieEnBz+gBzvqsoHXcoDb
WddF8QDWRGOybPP+xDgE7WYq/GeLLmafTxDWF4adqTQ1FL/JYKKrX0W2VlBZeI7Ok2MgppIIWdEz
WagnjBZ/emBqUwMNu6dU7PIPILGOOtXdXsyfe1gpJ5/rn7k4LbPm1oEP/CpwnYcHh0zi+K/z58L+
El4WhfV5FGxZd2iK5xP0YZarIaLWou2+co78qayNSW1AJJH1Bx5enfiQxWKQjjFpfOaylVtJI0k2
TRgaCWsQYGGeaklGqoRXFGqh4cXgj9B/OnzRDS9kR4KRfGEGgEWgEbwArr2NRMGtvxXQBr0r68LP
eDrOK6pWmoYTNZiHFFuz4B2o8fqx8Xq61QiJG3lr44LtkyT7RrGqyk3oJtj0JMNaDVWamFaaZOWP
YqzopqbTDBGJoz6YO/PQL2kB18DVrbfT+MbI23gbsExIl87yeVPl5YxU5ajSG4NkabeXkf3Rsk7c
iebhV0bD5UbV9SPyxM7OUVbRdS12bUhpg8Tf18lApBtWgV68swZmDmF0nxK/9b6buhalmI2CGsDH
C+9hnb/NGUngZvR2+Ls+m5B5h4WqgUF1St9sr4aLc71fk/uakupfCjWwW2I+Mj14TqjNsKbmNvQP
QZ80Qw8h48b9oIo5DOt+GiaQAQQLJbxjRhCBmjwpU14fH3qLJI/VSOvoR6nqLmYPTDV6bsuPaj/o
WMEwDOpyO1xynh+XsIqMab5O3MtU2Ut+EWoWUt4f8NmoUVHJ5YNEOPX1Od+s6H7WKDXiAONZmpiE
my7CCKkAE+mzKLqqVNSq5HskvNYJ0WxirN9lISlYYOEl9ut8M9cbyGN5Q0zSeXXFJEf/V0f1q5kl
s844uCT9dedkasQW0IHe6Uh2x+xQD93WgFQOqRcFXxtwLpR0azx2SGphdBKnX24xdPE1UqZFMb+7
0QufGfVHm9zJtIWGqVWvJESkDcoXgnCBimRY7G4oimPiPx/FQQm0EqSaWMmeXjDTCCommQanmRVc
WQ8FZwVsx0azbr+iL7OZlTjs9FPaTMklJDB+tTqmYP1qWxmZtl2vxaTlKaacCwzRTZtJ3S6bKuKx
Ck/bp27XDA7uEoIN2s/H00xWAMJ2zYtFsdtjs+5t65IbC+IisAb8SF2P1PI7vGoElUMBHWg6DbA6
ph0CUMSnaTjD2Uq6aZ4FU5hP2HjkW2n38YW3kZiIlB75HjjXVjur07Unl31ipAHzu1qbYRSaolFk
JBYQrM4x3/E+pssphhLNGH6p0MS4yd0eCU6gULkFn5U7xRtVndwgF/l9F6k8U/jypWlbbd+2+fBm
6rDrhfSzRHr+AaaZV0hB/YRfjcMvfyPDPVLLcoZMHoXzlfclGsaH5x0bQY7vijaQHbw676szVznf
AFSIY9V551nGnjaM7G5WAERv4M0eTjPTKrqSR0LLE+4v0OlQEP8G91qlyMKccEBMWDls2Apw/SGf
VwPv2bPhaU6LEfp2Q2XCddD/p/YWA/U0mV0y+TqM5SIPvHr4kIPMTR3fSMsiJud/3YeAvZ9NHKRe
VQPtPQnPogb7rLww5YpbgQ3lUfeyfhMhkT2XzGamBv9y6CYiRmlW2BWBY6MrDYXFJ5P5q4WWgUBc
xuE1v3oloJdi3+o8UFB4g3rB6edF/qSMXEctjHEPTGpe7D2+6Dl2BZJJNHMiFYIx3tg6TfgCmtLe
KPfRJAhn7tdP+YpmwUGecISH2h0ib0i9+TMpScli5eHPQqKqE2AQL28t25eX7MeEMqVeRt9v8hJ0
IUsFFMK4IqgTriZ5SpJL0dDFHKKD4UT5MmDdZP2QqqLJizSwFdSskdcYSu5yTjUva9vbBVAtnv5k
Jv9AbYHa8a30B4dLwzxK6dKOL6aw8A5J1ZYuKKrbWS7omEna8ZXI4dzcglVwp2agbdsx8kFq/3Qx
AU4RWhNfKAeyv2FME5EovbncWvnyaEcQrZSV+BY+x4B/mruZgTzFqalBlVBNEnzxC7l1nC3TyOWc
gvIVu2ld/gbzALtmW59xWNEbVn4Eqc8lWNLb57YcWdhcawKIvQA3BNZGCkwOMiUZLgte/cTMPESl
R8PZrVfpYneMERRlYQ5g2Wxj1nNC2Bg+7E2woAKD2p6z9JXSCLzbdUqbTaXXFJPzkLwvWYkdn9yq
Xh0p/mPD2d4ypRwI6CnwDtBaz5m2U28X/NR+Lj5ab0WzYw9yvGFzYGUrWCqq9koIIvRW9umb47qW
0s8CLNAMsPl0aYz5U9NHSXKprZc3yDiQ+D+R8YOqyCEliUPKcOJzpV+z9zmAstW8BKrqWOC1Wia5
oYrjkLevWhOhiJkdZ/S7aZ1KDdYcqHsLryDdV35qo+SaplHoBLmepHs8VOoVy0wK/lhi7F1bMZ7M
2Kq/fG78e1jErTBIHRYuzgrOeuN1ysOaRTdD11aXCorw59Y/TvxkJ1DRU7IilJ2ZKpPHDGCLygZe
PSbjC37Z6oxTWSzplq/Oxzv4b3cT06MHOHsRH4k4JfT0WnCDfFWVN1sYo6iS+GXLheHj0Qw4zgVP
oiUH08mzGKNgCGT0PKbaoljzj72CrQpHqbnoakkXQOaXLSUX8DMjQjjON6NeAS6fSCDVF2aucXUq
PoZeu9HYrUA1bNP3ySjA/q5HXsA6fydy+SghmGUrz+EXSzbL6251Hq9GzYVRa3D2nlcaPLGAH4DV
qFGg5uS37WmYFlLzVgTf4TDyO6xZd9qzWyzqaFWGjpJC82+5B45DnBnMu1W6xbaXQToef0X7T4La
VgZvWAd5gLJnsvOSUowDq9Mr9Isuu5hcy+GzEQohIVELE45Cpxi+FJG7tUlC1FOpkcZNQhV7WrHJ
+Ht3a14BfS17GqoamIYDrzzg4Mrc4lKjj3qEdHvkN2BF8Y+tGQkl6TNta+QFZKgbNSGb1LKqGCym
0AOhyfv6moCpenTP48ECO70M0lwSRz79cx0+Uh82aSl0Fq/RVIdC6A0AGIo2d55Qc/KZNLgGP4Qd
XWMk+QZsRX2mryb4bN4L71nOyPygc2OeOpYDhvMtx7QoaAwhQtWXKycuiKHLhbvxfe6Kp6+HjaXB
rc3qoHmVas7Ylp8BMQvFizLR30Lchd+190hxbe9KhL1+3kBMzsUH9ebEdUmUwsbluGo7QMEiQjjh
7X3uHJUF7+SSnXYL084bLZs5RK5zPbLccsBj2EjtHpmxQoeYCkCjQpjFR5L3bT71CRCPM1x/vTuM
0sd5wvUVoXAmRl0usc6uT8XsG7+Uh0XwMgaJ0p6EUzdAFLsiTmFG8X2kg5e4A0ptrYal+qgLSxsa
wzXhWTaAC33trcIQ3EEfz4BQ2GtWL0DpyhTmK2Re+AbR5nAKAKUrg7ILdolj1LnQLKbo8v7qDZWP
OJVkuMkhY0SgaiCp+8zGVKBMWkwkiQn8zP5BaX+snWzozJ8NnhwvrrEjdvY1U+Cp/u7IU4NlZitR
iN+wk/kD6Gk+/Q+e/C+E4JN1EzUT9oxTP2qnO4z3GTznLmSVRiH4exZxA7D4sPlruKa69gCXGiSd
hJaa9dFR7ttkjt9mhpuqNioORzYu9IZoYPwR8QOEe6y/5FxZzspo9gnOw2yoARToydUCFlX4VCxC
9x/Wq9QwamHVdo1ZydYnJT13xXxcPscMYJWCb9NISmOBFCK7W9cPVCa62lhmsdysT/I3LBxwLLKn
9vkgHIg70DCOJ6+3MGoBoUS29qxvFXqOewoVLTMU0tCM0xnn+DpAyk2XBJx+C+fOObF0EgiXS2QH
Zx9E3yQfb6DoIsQqtWktfWh8DJMAdEWjlhyId0dRBblf+HdENV3Xwx5jhxNtvrJ7naCEqKUwBCYr
RcyGN3ZfRohs555r4KmFKiKTQ1QMzjd5XbVVOD5oQlxxBnP1R5fDN7ERf3G1VuSlqKSVapGtMeGh
2ycM4CMxfL4XcXiJiXLzM6dWxqthqOa/R555v0c9678xazG/lC/NwRODywpoSe5JHxjdm8bPaHH2
jc8Gn0eEIvNSYCSwRAX3pii5FTHGFhB67TGBGY8CImhV+Yt4Rqe//UO8A2cPYIYysQrM6d3Ggpfa
8K7tBATaG5e+YnpnKP+hE1/JChZKtRUy30YXjFsLt+/PtNpn0GnstYZGDYxf38GpJotTUJWYs7yr
WzbQMSGJIhOuWfmF3KWWxVqUfqahidNXsN+Y94Dx5BcI4eayg+9VmiYTm0/DKNQySvLETUor3rmz
MLl4z/VH9Zgf5ksz9YqA0/ZBvn96sM/v8wEhn7yyK1KKkU7mX6I/mv5ed4ffYhtvvd6RiKheu+ro
tYjuGkt4NtJZX7ldCOJuBXnKHo0MKvn4wtzbyptuiW/iySwMXhdv2a/MGCebY0J7eZ74yVY3LFeC
WjQqUaHmI/nOjWuwi039PdClNx22hPQJ5CivNJy5Y7Kuayqh2n9vODi6jpAyBPgHOKu5FjYzomVa
1vlkJygS6g40av/1f/oVGMk2MUEWTp8HWrQICuhNyMGz6e/ew9EY4vfZTs1OkstN6Bzi0srHgm9f
pUnZfcKk228EYZ7SRiCu1uGgouFzgYxMTt5pUCk4RaqaGhZZjcwqAojCfBBI2+gd6JuokCyHabhn
cfOY2ij5Nv1tbGZ5SCcuLZ8r2qXGjt7v8oGcNNnqLinMGRYETE89LbtQSCoA4viZuThbnvYZXB2F
skP+dLorOiXW5ZTBqwzh5b4YwtlEepiLZH12Cp2D2TfWy05sxR1SgRfvLEC8UNpumNEHuu6t8G8/
9EZJOpRPwUlwcFA1IasqQs4Ws0s5oxpLQIW1vYQU8Pfg7km3pn4wBXNpo6dwpBuyyq07H4BeQ7WM
PMdCeMQGZf84cWisMW2zlZ0I9smFClhC9ZaOj7DsQl1WCTYiKoJO7yCxN2JsieMu51g1sxlmnHU8
/wYhHlVoeNyEVB/efS34d7JejZ3DRGTzXdqry4e19zp99Ch3zFkaDL2OzGI/kKBZkZwAfsVclZ3N
GeOSdPaJah9qzzhOhRuwAv2Q9UBJ2ePTtaIB0lFh08xNsokj4ioKpkVoyN1KxSkpmnYTkmzAhmZI
0ja3bC/ZxXyDoofy0k++z8JZB9wVvR2HO73W4H3z4NanuACrsm7Mn3/8OfFdhh7fj1YURnpG8F8z
o/kpTKhPYUJBksVFwNrRFORQy19vAgmqufG796yeii0FgAH70HOIM4f4+M2pRqrRWy8=
`pragma protect end_protected
