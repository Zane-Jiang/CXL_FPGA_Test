// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
wQFcEd+068OBuTk46Ft7xdOyrBiRkIJC40kB/kAA0S1tBNi+x2gMht/JSUZeVqSe
3SK/Zgj3sn5n42GoxkaN1tVqqNjoEh4m5SRWPXx22AgRlonn+Y9ahYAav0nbudw8
QIbn3SpfykmekG55mkQRxk9bZ7M+uA8CHGwXuZnAX6Y=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7824 )
`pragma protect data_block
J5GtAoA7X09AeFTO9isJHd/lMAJutAcrh+z4Fh/bFeehcMpOFnrsnEHAr7Zc9d4N
oxsA8MXsRrRMccvDOZLuU9r8l7FXYBeUHvKEP/LF84STUgBkjJ/Frp+AbO9cvUAG
7AB5YXg+swLSqFcOWG6s6Fv7MmZvxn7PIFZVYPp/3mIGeVnIG64QN7AzyeQ7KSZ+
JiDKA53ip46P7vz0Jya4uepCUjJzAVKsTo2y65onkSPA3GFZxP3QQui0ZiIUg44x
6u0B9cp99Yqm1YBRYWAmp1EM9l7LInOBjwMo+vwAWy9VogLn27xx6/WFgk9n6vd0
UMCdu2b5aPinqiLxyGtwtfzlZpfdOA4uU6EVmJ90hv26OYeYcbJI7iyODrjXxJSk
PO2NrUztvcTfvruO1tNAuTPQ28ZB8xfHtINvBig101pPX6h+Si6asEkj+yvhY/ln
P8HCYf74KyhtqnD0eJhk6GDDsOZUtooZMo0IFX/chKcqzHwgf1E7JK8/iaSL63Ir
K45sy/DKIv3/ZPfaJCgHssfBOaIFzLTvMHvk/U0iYsjmRN+oSZwQt/7lQ7jO1kBs
Ei3MH8DH0GA6VwKl8WQMopihCV/i4J2rlj71HdFqC0AvIN4WwV13dhd8vLGlNEpU
SsqJyGaZSw8BcWr0wLpCc/vymGqHC7ZW8cCKdXry9+ilcJdAhIiz0gylAR0H6mnB
5PD3+77neozuJcjnL5+WwVr/bSVC3hoCBgNFsAdrxoh3a4ikt8BXjd0bPnfnUppx
gcDkji6x/ty8VgsxovGszfuBkyGi2KIl4fcpgkXWyOv6Mk21ZKrZBdJ6MkF/LH2I
Y2KHE507k5HrAQcMefkYHMmkSHC8v70E41vCTu3qNE9EIdMuUUPUDkMGg/BgxTxB
CfacYycYmt7a1JHDieSF9jkNrfo4Uc4iJ6L2ZnqH4sVEyRGRMHKytzM8CTFpnuBr
sSeK0+o5ZLZ3qWkr28wg4Na9t35Jkt+9FfSvLTwhfpYsUxdl3CTxK3E1Rn+V9OeR
sPbEiCd5z/l9Sk2u4w3BWPj8GGuq1xm2Z/DJTW+nFn52n6XdMVAmP1OHgR3KQHnN
oGF27o/Abvd9sC6FbkfI574Ub7R/wuqZfoyWNKR35UvBNLOwnTdsTubWzaScjFqz
8jYrV3ybfjo//qxgI/V7HMlUaoKamJ5gTlibu9lN7GrVougGo/4NASnSZLWFrzrn
tFRD/JV0zkiPwjgEr3SUssIyJPM2S2Hcj/rbNAYoYte6IB+OdvUS149tbdLY/vwO
/dvcrfo8zraG03yoq85PhaIaHCRlQr0tttwhDR7bPS6aqd1kLb/fni/TUJ4e16uK
qG0XuSeN5UuDM3COEgOwM6znXljFMZOhXH4sOVemaUtJS0SDwgSS1lTxhFeYG8l7
+3acmwK6uhNrv7m2DjT/CP8+3XZYij3SkXSMsz+2j2kXIENVTzIlCTngXBfU6WDx
3KWCwH5CCBToY6A88gonVqqP9Hoec2uA/hnRXFnG7Xy6Fd9Q/g5HxVhRiU65bQKH
bSEWdEbXh4+26bxlW1OpsFZSQXwpxbz/mMq9Z6FITbS8I9KTPPUbnnpQWQBLWiH6
YIdB7ACgyWhuGzcKYq9/iu3cPp1pd0RZIdEW2JunSDL3oZXOokPXwMBwdWYbA+5/
5yxfgEPoluSdxbdVuEmKw0oG3kziaFxf9bCzJ3Hp3qawCG1Xeh0TuDhXc+0XULFi
Mwrm6N9Zlf5EIp/Xoy/RwPbxU1dMwgXhE5/FcmaFeXEQvFSD3SnEXKVyyN/KSrwI
5iY3tPR6qrDR5MwQLilbZ59F6oP5M2dklpC80BqiNslBFWXftWVx9AOEL1x+JtZ4
DiVOcJYKb8bOiCU8YXm5ykSgLyxWKblt0l4mAfJouvw0RYNgSNe4IZaWeCUb6WzH
79qLGx9OYZHr6fbh2aOeVeTXlAbXa+vcI0CurlVqQdPLIrj+kmrHnX2VsHk2j0AK
dFV7frAIkrOrqoAkLgb0dx8/34siOVsv2SPkPTJAj5iEuatpsqctar8K+Yyuv494
swQVx1EoJy8uSMaIpmi/z5jObEyi7NZQXtld0wuCfrjTwJ87umtc6YYAS8wrPhke
pdJpLRt8tc6hM4mlDXIQdZA7cU5/7556g4yLS4YmDmFFOplKAHgIOZmZeEb4SxLr
kxhVSSiZ/GoX60MIsc11rsS0omXbN6e5tEtMXwOA/QNdbdzLL4tCLVBZz8lFzQDD
xNYJOIMn885U0f8iCmD6G8iyhWYh9bchyvFYTKM+JzpQ1QH1UFj/2wDbh3Fo4JS0
xI9PfJIWLF76ufeSUezZyE+6D6GMDiN+UiqDqSs9gRZXy9DJGHiZ/Qrv7Xhj8vKK
kajV3UDJWn3F9aIS0/Vk/RIcpjNWP9s8z7rZ/ffzNNd2iuldYCBaK0DHw/TVkhRJ
CJCAQs7DJvIlY1Je58QekpYQ6zuggXFrwaIradyB4YEDkx9cbJ1o0Ofo5cRXTJsP
BwPelnW54tkPqIk2hOYFIQZ2GNst0lJA7X4Nsnd7vrbl3IEQk7Z4DCEZMyduyUhU
bqpQgLlN2N7JfEk/yTvaUdyWQUJ/y8/48YnzYmLR6Ofc2PIBjxD+wi+ui1NUp5Jn
mKvIfg7+pbueugsecEyEZFFpj/+vmKCIrt7/fscfQih9S2//kxdtXbI+x17hu2He
cZccernkm3Il87DO6mQ7gpSCD58uh5XrLGHUZZ3jafvbR9E8lK2jQaD9c2WGcyS1
F8SvEqyAg6bmlvzFEHcaCwXn9RD5uVO3TsbulhbcLeTpktlSh/bw2jrG6XM9ImoV
5HeOAlJnnD6l7eltvqJfIhaWukWYOqf32uLiMJV5pZTxRlnqsltzJ86T/8qf3VzE
bmAtfIGzovxBPkUfNxCDhz5ZIWiyqirUHKhF1T2yZ4yQQyMD9xwp8aYOiPVtWKII
lT3HwRGd9i3qizsSFpAz0gYXmKzP+/HY1CimbOAtMBx4XKKOAn1dnbqD56OZEGWg
q45eX7wkXSSTY7q5G+1t0TO5jJOkK+4TGZW0O0cSsmMotAD3HtVMYQ06QV7nc1S6
VQCZ1PElKnE5p2btVfKN8hxQ/2SQTPzOcGUC8qcGzc4tUNcugXy5Pid8nZ2/Dluw
W7cuaS5QDqDtYIv5G87HSpHhybUB9E99CWQ1loicp3/ExN7OE30RQRjsWoeDOGBe
unIZnToLV9tPVnzG4w0nKEWOAR5PzctF3moRViR7NRg9FN+PpfpR7Z5o0wNTBsnd
L9baLb5zEmlPE0c23McOu31Zv/84Iu/68ugLegqW+a4t35eFfIPNRLmc07kcfDKx
be1oO9BF3YXuVl26IGnRcSqkfyBC0GNb230VDCJqrqnRhSNKH8NNgVTIAYqlIaPy
HaAGdoD3GwYa8qbnQnfAwWGPxq72mspa3Rrm9gclbW3lvcGufItfjNio1l4s+ma7
Ha5ifXpTs8h1CIEVgMadxBUjwEV0rgihZCh7k9BUnVpHZqAbi6cgJdVx5Uk4LKI4
eeQBALx3XmXBtLTGeRU8L8zmCPOyW3yzewZwNEoxyRSwxjlrtOAdDHQgVD/2zvYj
UmRtb4uCCxKu87zHFYKaa99LMFTvUy2Ve+clYVwhJ9RP0zjwa2c0idgAk4VZfDks
+GYYrVdZT7+U00Bx7hrHLMoni/Nh6wwtxq70ziZLmCD29YCQSWzRH8OU0ge61I8D
JNLXK0lzH7xWVIyIU2lAaGuQPa1dY70ZZ1kpMN0+qpsl+DPh4DH8wyI9F6y0HNqa
mBDHvuMSIjLdQUYoRDe/pUh1EcYeSL5OoeUdJQQiIi9qVQN/Nc1g5EexS4yXPs7x
UfXbiZOcli8e1UTEd6mlPLvpltKWBjvA9bsZGcBPTWUZZGVw9f9VPZ57094GU5pj
OOoRBSb4tu7iGGtTi2ynrEu7rS6k8lHjwUycKGBqwN+SH/tdbSAR4YoIpB0MuQE9
Xmngjd2XI9B+vehRgmoNKOzkIXfko795m53TFBrOiyfgNle+XXmQ6HSEuu6VUeR4
CgLsysDe8OD3SL8h3P2N54RyZLRQXP6VxLkB7P8fs+Cl+4uzz0aqe+8yOiaAqjbY
SuL6qKR7Nl8FSJRweU2/FCeM2BswrsD36Hw9MMFNk7X1IS2MLheM17kUtG4BjoP9
UrnooPdfyDMRXyxWWFmN23n5L8kaQND7Iu7y82i1p3PS8eTbg1R52bXGjg4+96+G
qWDJa45nJflfTBpk+Cp+coEVI/Fmh8oImPgB2Pyr9pbBV56bsV9oODwoStr/nq8e
LM+VG+KXGVb3t2+oH4R9Cm1EgZU2XGZFNQcpVNskG49fNAa0Dy7Sx2sRcAMlQ8DJ
kHhPORufEH1eaa7rn0WFUD3kv3jE/lSWH11ql5MwPQW4iBAWw23Xj77R5MyKEzg/
3s4FHYZleKQydLCiORtRoIODIWOcVqQs0FCgGOEa1i1szt182vxvnA9LFWXddFUc
xegDT4r2bJqo+tyi4wCadKwe+WEWthZIUBH1kAsqdcd2e89++sbs1jxImmti5ZG1
Riwao3WfvYqLj6KoXB2d3W+Tmmt2y2ril3BQo4EF7a/LaN4sgoeeO34rPiFds54Q
5T1BP5Stsf2awgh7kB99ts7GEZ3YA6Tf9eE9sC2lXl9mPwKQKZY4/7kEfT7kGsFV
AjYotmg4fwA8ZdN+BNVcaXvOZexdnX23EefLYhq84afcujQWpKdABMtwin0YPlXT
0oEGaR0l4V5B6iQbnbahAPoUp9L4QDOXUlqqerFJ4Jqwv9k3ahUraZ7ruRZqGkdh
pVjaYx66RuBir7UHEKQKsa3FMnE0Saitdon1Q7hG2C/uoTrLwxnk3unSmcfjs8Nf
+j2u+/tIWaAmysiCxd3hGt5ONY8YkZKA7GLuL4d3KeGQY0v54TDVJx0qgPjZFLsG
w1cKJDI+UDmDuvM9qv+43jzf1FOP8KrJXi7pg3aAx84HAtfMMjhVYWVZtUslE/nW
BRQMhpbXG7iNR1FVZ6vM6YhfNxEWHqt6sZzHOjG9+fcNUEZAO7tsd3RoKD69zT37
SvK2EOm0qaYKIdpKhvZxDrPzc2/sVut26hKb/AaiiAD0CxuDPcf8Rss9FrQSt1eU
GqODDAI1T4zR29OuM54eyIEPdo+pVz7SJVJ2X0N6n4GtJyA8e9gYfk15L+Szr0dz
71TSqIAgI1CsYDxTpxJwr7EeJNJZnFKi//TMjMl9OCR/cwBfKCH3Dp2sS6oecZFX
xY/aXmVAY6UBheSA9Cqb/ygO6jQxViCknc2+WObpwrhDYwpiuauha8vrE+eoQoqV
ku1bdVGIHX/vF7CVH6Us+Bs5lSnKfEGe174Rrze2IjTq7P2FmlkYMu0nQY/7uiyd
F3q27XGxiMWyyvUCTPP5oXQmR85gQd3FIEeaQKv2q0Rsd8f/HWC4z36x4sYxK3Ou
W727V66vVo1XszF+U9qqWDvUxAVE3M28TloNB7RbneV7sXXABDmwXTZGV1Vzr6PZ
cXj6PwdwAyMfmGlOrU28UG1qnzoU/MRWmN67Du105JXSQ/l97i6MaaSzWqWzcKOR
/C5R4R+ml5IbD+fX/ERMgW8jqHpWZXakCM3bn5PvENm0OwJdtol8lzxUlxVcqbYr
nKXSTqKGAWXrAEHh/GQNDgfRpogz0R4OCc/PzKP7qBz24W3dSHh9cPlNYUPCwYPz
qiXz+gKZEBrtOCMab7NVARML8l7RCznHiWMsychqCEqQFFxaV0YB2sGff3u0LDJP
DJXSrO6leFT8h2bIiT4hrsLf+J5yFBvqTx9s6bvdhETpv5SMut3cdw/OC+wTwDgQ
gBbhOlhZrBO71Re/VytvF+hjflLE4kS2ldTVVpeivmCqTCHAXIYQDu55Y0urvkH3
mvS5deRh2fLL05NanuI7z8ZAZ9MRz7czw9j37cgWjyGrwug7kkqzIKYVQZaQqh5O
EVrj4lXC9D051fF7ql0gwh9/YqI68NB+LJUi1aKBb8cR9Qo/7E0aujSXnpGoc//n
tGVIL9Frp4/HgN/DGSj+VtsZElGxmsb/VNmc827pwpqSkyprqjqm0HCJLDbpKp6w
vpyMZ5x5rVrlcZLjGc0qfFU57zwsVy+BQunf6yJ4iQPIllHu8mCDr/3Tds+eTljM
GJzkpe2kL6vaaLLkVfdMcpzLC9lpDQ0cGiIZvssIwXCxerYrtnAOLzS3yna4UJ/F
Ecr2pN4KWpniOGidwO1RymtVrba8FmlUIfMJDYSCaKGqrAERZalNYb6qlVhsHqSl
a+CzmfGb7dVIiSbhsuVDhHvOZ4h7vXYUdFZuLrVOhmXQZQMvFoHaDDfSyxnLchVF
Tir5/2ezO2FDQEcz2NUzqpHCw+cKphAoLG83juQSplcEjZkqRLY/EiGoIS/uhiDc
TY4l3VQBUHMuSIGLdX6dWc1+66LwNPwimP2vdH0F/S3atVh9XInhdtpOw8U9PZfB
PhTi4qDN3mINcaw4HYuHI5r8TjB86nNx8fb9ZTeiu1cD8CZa7cl1HvpexBtObEaA
N6wzPN62q3O/WCZZs5d05Yt5ZWcnKTh+f5Z6cC0Z6wfGmp88mTxxSt/cENFTDSn4
P79DHYDYmpKgagn94Dvj7rbi1XVxxytAV0mWn+Eekl7RFeIbpXCafTCSKY9JwjfY
Z92nf6LocP9S6hHdTMMt4b2UZMtFswP89xwvg/aPun/QOMSsw2JA5TpUQtBgz663
et9sZChp+Z4uCKFq0umT/1md4tQuvQZZ86Q4VygWQXv4fN5UNXT4kMghg7apu3Q7
QZe/73CKq/3HZdvnIwgtiTJ0W1Jp1sTWmDkhm2brWY+FdBt+Jq5po4KlJb5gdlGy
oeLW/AOfi/eJeflGSCXBTSwsaRlxBsh4jPnatZctSLsFRndA2JkfdjXlLjD01tdX
xRWxTgA8HYgQifz+zT2+TPbNxt3fN6GAtQYZOpdRZHEOYVehUHuF9ApdJlPJ9/uf
UkZHN6o/BzJyxSQWLMdTR4LvRsu671L8S+AahLjcLhigVXVsV7X/FynJs0FKiZCp
qLj+PD0xmqzKptsb4W7bByC/h1jW415EEAotxz+gYEGAf4kbZjtcvIOz9VHE6Z1n
AmjPzAkfI+RBPKxbvOS6Xnobw6s28pPvSImuP6mB/983/uXcYYCOins5xjWFrso5
mDIVZPXzJzZrbrqCmAsD8g7iNzOAEarYtcWTmbi+n+AnDBQO8Ex2bEbnXFCIM3yn
WuSpjcmp1FO5C4wXnrK/jQef2eeGh9Faa3cYaL4cyWVaSlasOnVUHLAH5gwT9d6F
+/jDK7Zi8Hdj0TbiOkWUUIKrDryYSS+5ZfH6x5RH58UvV1xYX3C4thS9ssJRub6d
Kr69rrAn2aoLDl228M+04Fl0zSFzXBLVrSxGvJlUwOTXodG9EvCEnipcRo2vcfyh
zwS52U4okTjHNo1v9DalLMPrWfX8EJ+D5uE+oCTaH2jhKirhYiClthaTLGek4lcg
5axN+knxUDyAUNY25LsjPmnfALduWVh2SJb8rUJSLifCCZgYX0Hk7kuzOL+UsXII
pKPkDvbEX3mwehE57GMQ1v72URQdJu+9cG3mylNyswaaF9Wfe0m4HLR95F+IMtv5
wDhs4wj9MOuxP84Yf7C92jjGP84Qs5idnjEnuPYfGKqgzV11VAtQZqvQCtR93jDC
EV6dWK2qIRn+mLS+EXYgKuiIRcXcLo8oy6EEqaZ7ytqSSIsEv/vORAtlBJy0SaAZ
FVFSbHnYrW1S0m8/E/pV05kPgHJF0iFh3t2YlbnQO4HS8WS4jA6wpmHr5fI8yFUe
ZE8EGKhkKTGRA4SDSaWcXZ2f/T+qRhjFGx7v8AddJOTRUtgzXm8vL8BSYfMLKFy6
lJ2s1ox7BDTlYxvJCjsEKW2UqcSENnax0yCeaez/BmgujbyM5BhR497gipJ3XKVF
Rg4QFJMVycOn6cP+Pl22fvr4bOSf+5uZ0Hx2edPsDvzwMvK4RCZ8P/j3OVCMCSHC
WC7Dyzp/lmwy5LhDDb0untK7JBnAhMq5W1ZDodtihYYKMk/3/v82iPis3Q6tbJy9
Yx3lxANPNEngqs+0wER47wMtuQUTEpVlGIuXnuLRLpbxEW4KJ+SyBJz/mbyaTJzC
KyI25VMgIqJlhA3YtyV2OlETerUY/qI6ROj38eEFB467zCbcmfRPLzyDwtqgh65Y
o0mRA+B4lZGsaxBvHd931TfolyLUvBl8h9SPO3X2gQTdMTTIlbUoWYpwIMr5jlE2
Dz+W0OiW568Jl8CiFsH2hrcZtK32nexADbHswwgjqb8yDcMVUxBTVhtqxuerkUhT
C6xkzTSGb42pcnaGl14hHzdW8Jk10/ciTFeyJmYr0KN2G0rODQepSsd75BdhO7bo
Gw9kHtGuuH+LJCe20XFYd8EuYAjZIrmtuy0exc5bHqYtFC+MpTKVoa8RXqNWn4Um
rNri5wY36gHFpYXAY41elEjumcqeh/CFH+SWjYsakQVpmYDVBN4ah54DWMa0gqp/
Sx2fkbO7oPZPpxrIDM24FQv9/TsI3QjG2aX73S5gio3iwy5EbaXhudHZZdi438LJ
NduoOZjHcM49vBg5/TCTUiyWjmhbKI7eVBfWXfr8JEmeqDWCDO9bz4jElSr7VkAu
Ghbj1Igof0XOxDI0pA+Z9fGaCbg+WpvH43ds4WvaGnpArnt18XbR2GNZVmpFkfDm
UpTeFCiPjHKOCAKI0fO1CpfWybPRLwEcG5UpVQnChJIJn9I3qIzJMBhM3ETeFq+o
3xmI7LJxTn2k6VtDgq25GNAalCP8wP9U5UycLZ/Kk5TO1ZGhh+Kip6cHugPCSLo6
Ip+qJ+/LTek4X2jkEkMxjvnM8jQ2KRmqG7rJFotKU7uweAlFKUegPLraS9Xl3uGf
Qmn0zN8VrmbVRVQ9AXs+UsX8fstBAxJAS3It7DH/6LzhKkZo/h+cOnruib2iXZZ8
vFfe9lsW2u3Frqaao/ws5uyIBUfdStWePE40Ybfx2i8Cz+S7buf1BCU1jm4gSrhd
/5W2VfubM8/jURhrM0GB0j/mWa+pRZm6ohQ5Uv8+sL4nX0QvXeOhzTJypRU2Cy30
D0dKCui9fgcy+1jm4DVL3+TRZBzmOc/etpwfO+guMxrQc4O7L3qhu1KmdEt1+gqY
Jd1RxS7qwUvzsXgIuw/AlG1LuW3svWY4IJHUciREuVykFBVyPTBPxy8YABHy7HP8
TZB/zvlx9+Ewv8HzvAB0D7CWlaY+UVi3nxVOy/fsj6UnYDNNGz7A6Kv3dN0zY9fF
vniXiRM3qXXMLdoQseaS73Wopkr2WvUaFsPjpmXTFCin88e4TyAzuEq6ywHYvs16
7mnl7z2LN1SBIgjGF4G+Tg9QYer+JPrRzB2sPzMWc+TQU4qyfpSq0UI1x+fGzjRC
BS4rkEblENmmhE318jE4aJ3Q0Oayk+NQJuHLo45qCgHjYSZ2Py32BHx176bgKWPY
nNqzVlWe5DTC1+oS92LjLssDIILIxLknZJGJKRV8IN7m+tOrW1tV+yeGYMdptLn6
IO8eku6f1rcMmxJKhcnFIHLCM4JkxB8CWH+cqdfqZZpTK7kCQ3mRQt4V50dkmfs0
RKQQDgs+ncPJuSSfJq9HLkG6bTD9tyoGxr1TENPVYBzLqEz32776Ll5PtcYAbjZg
dhMdajjHzGOiWZHBWh7uHJLyrg044uLdVx5oCAyLm/+p14ormz0WjjfppsaMnUic
3SAyfz0Js/gjeCGP0/nlJMpC4k5qZxKS0auTjTIX7T6IQieaRu+IC1Jyz88TPziT
q+T1hZ99M1xqa+jF6ufoAvovbImJIcckrjVStcdJp4TJ64nuNxH9NAq3tDMInyMq
GbClA6p1W2bpIG7nbzlr+FZaY4aVzUnhmlfle1vs0/iWjpFLEgs9Us97/6wxb5HB
8OlN2i2uzzaahtWaULbfD0RZL9tovOCmK9obuMzMtdzkTG2TbCBuJuMD2ybkKXY/
0MGyvdoJBigLMsaDpR0H9f7h+X5StG7tU4ZBPttWmbA2GSAFMzUMa2Ff0WGOOR8z
pPEtf65JBtbj8m1K2RNSKZljKDCq4ZpMWnFkpRyel71rADL26G5k2HY/01Nknd2J
xyziZBiMSmMHzuLQtbiOgetWF1CowlKAACmUc8UP8EffoMF/0ub0IAfd83HpfgCa
oxN3S6rtDT0pllHhcvYOPogELPVkKJwugX7V+WHdKD+N2k7IHyoeQG5/N9tOFwQX
TAaUD+Mg7VOsOk4LKaYJg42IDzb6aDtLtVZxG4F78TEhu/9+lVI/ywl5c3ZiE9V+
fzYp2f12gbMkWKGTd/OhJ7mtvWwk1hWe9iYV73rLH1cPa9QfZ3pRHdvbsNI8Egvf
QLCw7Byb5OcVOGKb8W91erTlAA9WvC6lWq/Ttagkx1oqMdwWg/n39xHqhqWx1VGK

`pragma protect end_protected
