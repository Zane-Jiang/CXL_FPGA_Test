// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
lqhkigpOM50Ngg+x6f7oZviWzuGI0Tw/SDZsPJbLsSBmWSxUePx5IwYcJ6i3L/eN
V4EVuOG7EagKQStnVZqowwASjrVLPBeTTuNejXnWh2lQa8mhOEX/LNNrlYdHvwN0
ZRrjO1g2m0QXxonByqZ6vWji/hPG5iddqDnqHOectB2VgClh+a+e6g==
//pragma protect end_key_block
//pragma protect digest_block
fk6FJb3CiD4pPnD8jSbfCzIySM8=
//pragma protect end_digest_block
//pragma protect data_block
ccnNpZURWQzmO4/cViGbnkF/DWJQfU9JXZJ+41LBJPJzVxDXEF3JhMCMxHVt1xQy
5Doa1aAztgxxiJ+Krl+ZITffZhrhiXkpnS28nbp6J8ipjtsi5UHrFKLE5xg5GS7r
PfQm0gXF0H9TvG6OwgwSSdiiO6tc++HD4Yu0Sho4ARMipdbdE6MN3x3k9gxl85Db
kUsOPTmRtzYgcV0E12c0xQi9TsUp0mowYUOazVXQ8yuKfc0yX9LfiQ3hunGulLAE
cT+zPQ1eHg0AWcVVFixkdvA2cR9C1PnaIxARZJMffpJRoW62L2JtSbJVwPmIC2/Q
IxtHxmc62daxUQTl50rZ0VZk1RMdglANhyr26NPhlNuWdJv1U8dRhWspP4INnZYb
cpyn8pDI/Tsm42K5+qSkBjNqqrzFaRnk0RQqDfGTPjSxEaSNPXcQa2jSlm3NFxMo
JUsT1YP/QIr0iaFI6PLYHEQSK2gCN8sEnCno4e0sXxmCPXfUCf0It68kXbhhlZDF
zdYag35cKufpMXt4R8/WZILCkUG6bUfP174xnUWCA8Ao4+GJL8wwS7IlCiko+26r
X0Jk3M/OJvcRkCixVVFcp/5EF70RflGpF7mxeGuZ4mfPwjLt8To0rItDRoOvLgj7
0MjkIjGr6whMhin3E8X1A9v7OY62H3kfn9s5cXQT6ZkUDA4yXjBjNKA8JKihoEmc
2zkmGmdb9qxXKd0PAFnbK/Q3UQ9CBeeRsL3k+9k8RcYbFVFM+sy9hI9+9yRSy0cq
W0+egZDeCfEuVCiKqyfKIbQiB/STB28c8vTm3zxvDSKTLTlUA41swbaDJVx7Me0A
XxFFzLnN/k+c7W7BLtVJ4QrZtpqgKdqExzGzuvYyS5y6WQ8F4cTfUtIw8QnuhDUT
EMKoWoQxbdY6wh+StYXwDePMGxccC0DS06J5U78tSOKrAbFp4GSFPQlC95723Sny
UfIfPdjeUtlLiIfxpnePMsZEy17GMxp1OUUCjTQfJrH/qokgSLRNlJR8iQES1Jje
kBWEMPZI9B7g0f/xiFnCWiB1dvMHEvuiHwc1HNztDR1p1wiu/6oMjR0cbih7hQU+
26dlF9XzodB3U9RildMVA5F6CTS7knQRUsHo84W79jNCAMjyr23SNxUvyUGRheOu
UQR9jDNbyk40z/FPSmYOYSrBB8n+VhHv7V0A3GiE+t8Nj2XYwnXwZJkDUjEjRB3C
RUNdUDaI+09MtOvUayFJIXgbsOcEp3keFeIME6WYcMUEQ9z1YhfVvm+YpIsxbrFD
yD8OJLhPUvJnZ5eCmbx1P//EKTUCAsPD4QPeOo/DjKulbIljQnPOEXM68gEu84y0
I/RLbnKCsWB5REJ7Hrj1/Eb+grWEDhQE8hAzszPEh7vMmVqDN4Ab0Gnx9XgPlH8L
1loOQKe+ouckH8XHj6o5pRzn9FXWqxfvP7F4rLgKxnuSMXxSZ8F30BRnEp4+bo2a
VbTgm2sxEHRA+flAWap5vYfkZeF1n1zbZBWnVisa3RYOj2BaggtCuxkMFm2W9sF7
XgqKaodV1aqsXpWWCspIAUKtXF291se7kD2fvuNF2IEgUtCpiR6ijv6+twrPNTTb
YVcUNF+5DNAq9uc7dV2ITYIIMb6UuZODplv3nOc2gBgVPknHgsqqYg1bW4MKHQdl
AMdh/TxbPsuyl+XflcyOLdgMhAyxIdId8cqTR1j/LCo3I5lW6ZnrBi2kN0eJMAvz
q0JRRbxpiHxKVAWRZYvDLI8FuhuzDux11F4E3ONAElsuCPM4s145NUDQJknoGEjZ
bRaVojCjN0KjZCy07W0r/fCp2sgs5Nc4QZG2bOdCEoGUUF/+akG0/8IzjqMiBSq0
0JPqu56dxUCK1rlQJgu1yUQ8ZTaSYTgUMpiipUWM3MaMXR4s5LU/NBXrbjCCalfn
7I1SO8hhq/VB33ON5VXmLyOfHe7bTQ+aWO0zpfYl9FTrUA5tYjaPSDkd3C/INREj
R+RpoaSVJZTofIC45Yhjxbg6KI7nku+uP7REKPIX8L/6655qIewYtmNLK5naNxGn
c7zMdwac4NXRF6iWvUixSaLKoyppU5zuo42bZXXO8mAbDFziP6GHsJqJkT8+d5jH
HikXlMb9yO1AaisYF+WXWB3DJsI0Z5CZLscJZtuihzfWzm/cw0pTqJjYpMF2jpyJ
0ucn1IlijZtCuqz4nlbYAvoXpQyLhVDB0OOVZPBPfeGj/2tUgzbddKyT8jiN9ikr
Zo3Day1A6LymaBVeWvxrEdKHtb0nE6jDmss7HVHqr0w4QvgzYvdhxlnNTblKkIaO
lRzGV4Bceoi+GXAr8gCVnQD1dJu5VgS3cSQT9OUxbcXbBaoMPxWAAl6UHb1OrnJD
U/QGx2d7KWzv4Jnb8NPG7lsziDxwvA37UaeM7MmI6s1IzX182ALS3/lBytFBxWP9
rMolO2otVWYTGfISceawUQrNGi131b8KhSLsF8vK8fdmFJWTMBrz19dHoXShVg3z
vzR9R/ltQCUaD2zkMIngiQEjwrVzPr8Reh/9h3ndDCo1jHvcYt/EejwRrLy0evHQ
jgm9W+IjWJEfcyq+ZCd3kqK6PU84+n32cHQUr+CLfJh6TYrKOREi1xsuayH/SWXq
kPWZxA/c7iFj09FyU+VdE4NdG9LTj+gAUqDUfAyiuI5Tew7IiUZ6GIihbsumTwbN
DQskjm4AsleixinCXNcNI1K5k1H5GX/SCogm74BeOi+p1Ef/DhfU2BYrX6UWuxvQ
Bdznljgic/wWbWr9kCEi9DVT2GxOKjIz3qMPh3J4YKsNg3ccCIY5UtWv5z1JKkTI
86/gtpXRm25F0gBN/4ep302lvy9c3ahUZzw3lqUozFA9+xwb/usrUBMFGk4rbn/O
QySBALUmxPfdKaEE1ghZ/BPFnQ3aK7vNAl/NN7+ADjzQCi96+NeiWFgBKzhRUFgx
hKnyVqVdD7Nka9l3mEB2S6zExgUZE1P6uv0gj6Lvsuh2G65u6oI2i8VTLN3mdCYx
fPL1w9DWE0FDDZOR83nycrIhhOxxgPfIpOO/BbQKjAaik+tMd9b1DtVPP/pQyQpM
npBtbh3WSrBGIQt4x+PkHDZye2mMEU6xVik6Jg31m+YiX/2dJZkMSDgiHmEhz9Ji
UlvAhvTSHMYztzXqNVbHHCfBZtOyq3PC85BZZ95I7jlFfyct6TqcSYWr9HjAlZrB
Su6gSZsSoJLS3AK+PSwvGQbsUFBQPc3UN8mMUZCkkoyCvZbYdCrnshT3WhFXqo83
ypGjqi9iT79e5MiX0l77JVNJ3QsJXneFq01RZyzv90p/sg1MpIrcE/CpnE/ZqjFq
0fqXTBK6pKRHIAWA7Wpc80Y4lv5wq3nulYp6figVObOzIWR5arcRK9PiQXCEuZ2N
i/VoLsSCxt3rj75L9hTeR+wlBg2DKd7HrjE/hlGQGcEXN9VMjrF+TVtz3oTKo2zI
5rTQCndxOEBR7EnnrbXR1r714XpogdB9nKa+LStHALT238TreohxjOVuw7jMiEt3
QhUE0jbygYLmpgWzPkpmf2dIiJce0/1ujyIfsIDA9szwUoi5YiGhNjUKDFmkqsEw
ZXZQGR0eu+o3XM7LyrPoudd5xMRffWCpuXeMK1Khyr+NgO46acSok84WtMeyofE0
kzuQx0YD/+/L0Mdhu6F0ce5hRCmSzOFLE5MYO4k4qqmHbCxl4tRe9mbgj7IyuQ6H
PH6/Wh/z0m9/rGySps9jUAdI9npnn65DsSVgH3ajYVBo5L7BwgKppyOhQD5DVARZ
0VWIwswx+h6T3SIDgSp6SRgFEak55Ugc6zwlYM2hj7WbT62a5v2rLdj8VVy7JgZq
Gv6XJ1k40zKz7KsO/DAZk9IY4DTPtoGpPrIFgCGD0oCgPaYHvU7/QWS9EywVghYJ
tqSpDRJ6tOva55t2ypFTF/uAQb5YHk6EoigkQp+ZqWbUsEkA1+sa02QDon+ij8RK
rerEiCHyXty1xGrD83VSnph1EoPkvmTj1XepaGxAbZY2t1gKLWkTWUo5rRG8nZnT
lm9vUy5QE7Am+/VXAled4Vkj6tioIhAyYbSug049kFPn9QBEidh3s/xpE0Tbju4M
Bh1QRYWmzOt1YHjmJfOmKooHKEusQGv2mNuIeWQUhO9tVV+aJiTyBvxkLPJK+9NH
y2sAelAmL7id++MRH2BeUMeCeU0hcjhgFKdk7GMg9mdLnD6giLE0uN3tux2R3o02
0KMzmNrcEi1qiVXBM2Lz+cOVgMjQXevNKQTpX1pmg6+buBHhGD4EcDcCY2BybNvB
izS2vQrVyumN+bRG1UgfifeN0TSg5qys3Nrd59GrCj8ZMW6F+nhPuxaF7ZhoSZUg
B3zP97YM2RJ53pdOtXCacrow6HsXBcWD8lkvifvcV26wQuDpAvnLs+48RUuiuLYU
h7B5i0AeAaNZDOrHtoXGAFc9LuKn1G0mRqLKK3NPaxjM0VIghkwulajvodaQKyEH
+Wbq1KyWZ+eLRacG6FOq59lC4ULxwT3633gr/Vvr1zg8211JgAVGvse84c43YU+K
MfOCn5wU/FW0qD2/vK9Q/XLKctW0jm5gFoypXPco7z1pMQgYAjJPG+Dj09hcLGoh
lAdVlpBvfA5urR2x+zwY1nrBHO2YXkWKYbs8fnI+Obk7D9FGysIMaTF2sEyh2Z0p
fsVASe5soHtF4i4OQXCGCEI0HVpB+UHiB83RrCFAPPob/XDSE+d5N+wGxjutr3w+
WWs56SdkZPt9tcXAIeQ9qBCCoFXpL3LWqlzE7Cdas/MJ8TaJKj7iCKLyVHuXsM9e
FenPqncgPmmzUT+7Q0GwWCCxURz+ERQ5k+xfJ7u+L5pT/6cK8AvC6/TiCa0pWNFF
aNtYx53iZdW0GBlnmJt1s7gBuEMsThD3Yht5sFUJsbR8dS8VYoO4vjHW7pLA9k8n
fyXlDKxjcJDRU0jMzIxLG1y6M9i5jstIKPNffudwXG4/n9Xl5uzvZ8/Y1v1w47qT
SXbzMRCZ+sqcT8GvstYnaW8ywLVz8hySI1vKendBhYBbDvW4B3u1PgPNIVQ1EJjA
pBgWXOxo3LsBYpNU8su5Sa2W/JA7GBrLJmciD3pi2ygg7Ufjxwt71ZM4xRHZZPYh
tFXgW2uxNckgSHrcizxr2QVw6AfYT7auW94CH/a1gyXxB/c1LHjf5xJAoCZTcrp7
mYX2DZlueC7h7cswPWg3WIXUx7d0srrMWJh1eEZAMVV3OYERg/+OBpy63+ecq6Q8
ZvdPEM2GgFHdTx8oxCxX6Gp4cqrrht2ByoNb7xC9nY/ySR0+/+r2gPHSLwgT61PZ
qeuBpLwAiowZg52Yuf7/aYqd4ezCMTvPRDzZTRUDDUnMtIBaLIcf8Fgju/pBUWj2
OwUxix/NRjzWNzCu5dNtxOnF8ynWmtycUIsbG1t9Qn+Q3Dgfguf5c2hSOgpD7dXo
q/QF7vAnFS7a3jnvebmbZzPZ5n11G5cSYeP87A42NJvsiywRSWWzMc15iI2mgGyp
NVJKFJxXc/P3nqYCdr+BTbeHGey32QS/En98zhWuV6Ilhnk8Rk2twVbXnzt7IN+g
Nc9m01bSFcCIKzNICbRsAXlYtp33E9aY1/jWbFQGA8Qi/K9XrbPfSR6anjsrspil
OdBH3I7B4kzjFlL7CCl9mmrgKrVPagPkvgWqGx4Z5lH1A4jOc7p0H7FJ2peqFueH
hCKDWnl2bSlCR4PD1/Q0y4h4OGUWuTcZSjnXx7Xqpu4P6z2ozQMp3IndRGgMpw3m
OtDP4ItnkGocbi0uSbZ/SrsGBql+qENNTEF0HOk1+DjwDFUBwVZuxYj0c6s6g03Z
CE3rq/LDabTsKY+LpghRxdJDqu9fvPGRljMNwZNtHt8NUgBtUuIryjEKZ0HS5dcK
qBUejXqW49VrMrcl1ODCx3j0j6RKRy6dHbIDk+vydrKalEO1nA7mrVFru6Y2Oul9
zw/ecb18fUdQI28pC6Y6LY1nJrz797/0pTgv0EBJN3xTR1H9cMR8PCDUIrUrw7em
5CUoKKoPHPe1vsG1QQXMmQ1N/qNxX9M5HEZokAXfKmx56wIRf/jFitIj2X/T/HQD
yyvThwE+cxi3QdymM6YgYBU442HXq4PjnNkpwxAsi4qMy+21CoVoJdKcvxFH5iJO
SfRrBQETDupcx9A1x0ZFf377U+A0yN4G9SePq5YdAJ58LKuzarZX0C7bMj0xT2GQ
SdXf0CdV8C/6x0nsCdM2X/O+8QHGdx+ZYTUtWJ/X/dgB+LExbrZpP5jgmrm8ZPhd
LmeCYQet2jSL1nu/ssoIIlTVU3dnDBHTIRopdpLw0CXH92f1j3AKhXScMG2FLq2f
quQpTNMxlbfOAJO/YkTG4y2s4a1xT3Tlv8QSUgod2BEGi8YbgmWS7Aa221E5+bx+
tFWciaaS/5cv2sr+yyZy2CDaT0BZnWWONDD0TEEzisjQ5pc+EVIOZB//gwouGaxq
VHdYBoqH7zm6RQON3/6I+beVrH9oG6e8jJo8mCEodqiURYVTuAAjGsv1/hzP2ixk
qV4h0gxxN6HAKqEN9nS8BR52d7AyvKCkOibY8p6xj0Mnd5dICdozn3yN5+2GIOUG
dzrbSzXSS3bcSan8bc1duWFnkyetugTDVyHrJtBgCrlqgeNFpKOr4o0bhnD7lQNc
xAbMVUZZZvUz/p/jr/MmrrG8oKiaQOwdz0gkU6zL4CujPNY5MA1xqWTooJVjR8pU
DIIDvCF4QZ52er0LmZauJPPY4tTdfoWYBZF9fwW/0avwzvJQZkRoWzgIRYCjN3RG
X5N8npa3IsZEMLtg7lCtc/JdlbLALDdzoiBOLvDznxs/L3LcKlUOzxUvVcE8MIOH
Z1YODFnW1CkDMgegrUnKHCsFjw5MB03NeoxeuWUsPenq0mH2JLxGTh2zsSdZiFbC
GmRnBuj3iBWOA13Cm3fSl7ENk5JlWScsTR+nHd2UNoq/nTJv/Zcw6Oob6Fif3xNp
iLlmRGPG/Y/ZVIZR580EP94/5hRyk+WXztXLoDLQAi5LkVnJi7nBU95QQ9MayXTs
oT1TKIlaDkOf6XRy481+ny3t4mjeJmKweVUd/vlpYg7NRLGnk9Ybrh1DotgK9jWJ
KTaOOR3OlClajaK6e6eL1BPL5/+wGxmjMu6U1QTPn5vJqxFAiC24FTRs9eozo2lG
3UswHii1x/sbNrtSrXr571KJwLRrsDySiJU3AT0cCJkMhQaIRRxkV+tVzA48zMT8
RxyUi3gh6L3kBBcSx6PwPRAfs9V7Cc7ZoiDbt4WxIUjuGZl7dTkgwZIMylpyQCut
O2VhZynBsEiohC8FWYWpUYhDvguAALnqF/3kU/e2HarX42agOQWeAFuWoAFUevAa
JDFKfIB9mIlfuGTuY7fGWQQrzmmvq89jGUV2WNH1ZDG/H0p4qsQo39ASN2dDVmIL
eg8HprXYkoK49UpUpuxp6EsJalMXzbB8t7qFm6ZxzfmEl9a9jeshKsYszMPey/tS
7c3OteN3DHDqpsBuI6NZPE6EQA4GlVC8Xri3IqwzQp3LOYjbf5XAMcpwm3U7dkul
6vLM83eyANgqlplNtUqka0xgHzzsf+4SaXZJurWUUqhGN+8m2bw1jgvdsKvYBBtr
j9sA0jPZiL7xx8LbHzwxrNPycnb1s8mVXndcLo2OlfZxGK3jz/5yQYZuWp0IeZ82
kgZXR3TCI7vlJRM5Dw47sqZybiz1snbB7SgWWINuoxKbIpC4/KWXCKVp7F6UyXsB
fPUB8Dii9vSmyjTvyC0WVUkPl8C8+68O8j3rkJCLpMF47MOMCm5n9bhuruu3duk/
I12htxW6cJ6CjsUTIb6hqGF8ZVEZs0CIQcMf/HcAQ5QiNJ4IE0n6+H9O2Xi8y6d6
3/+e63IaYf3YeTI7NNYY5mw1t8mCsiwzleumQ8ne6u5vOOzn1CGBcNYOdYKEFKx7
wCGUTZ54Nik4sRm05v8jZ2d3aLXgbxBlhH+RGVYwij0lsMOGaFeRlaxDDde5Zfqc
wjoAZgF0356Uaiom3ghS5+bCP+AGEB7gm4TsPbMbIT3AK1IMVjuV4HOrx0qY2nBf
KF+mFdYVn7P8TG1xvvnEVLtRNc03jXBcT+io+sAC0WCvZLyQK5ojBDx+aMJlEOH+
Gi3RZGd0mmYOrpeTxOSWaCAd7GLNJy9F6+xbuPPulRVI8KRoh1RFdCjLPEBGyhKb
yky4+7SrS1cbeXO7PIp1AAx6XgtcJcqwKWBvwa623x1gg0EZnje5II/fl5T33Kr6
k60qzNRX1KMpYPzo1rJmdhSQfzpLaAT7Il+lVjxmBpbwK3DVVEkAmO39RvUUyUkv
kucjk+7Ql7rDFOJaMObcjBgwAhYZ7KASdtQPSbk6bKBD0fPHKLTl2vGBKxr2ogcn
61FqODFZT5wbjm00H0LfMO11A/xGEI7J2QAeynzTQThY0Fia0cYSB0vIxi2l7u/T
Ql97GreXicDwiAbnZNf/EzTlSOTCE8vxRJw/g7HynqYJXVjgsd1YiiXSZKYW33Kh
ccRuqUOd9SczUZCMOKgG3ZmBSOxufCREtoQGjndnx7y0eKEgKB0XdUsnfHXtFS+6
ybC7vk6y+24QXRm1B3EzXS0DMNJc432ZZ+y0I8hWI6eaIWeUe84R+ssfbbCYOHlC
lEJ2B5XN27F8pW5LmWUCxT8Z/FP8OWqkG4rpcZiH1tBOoo9Zm4Er8P/KHz3Ebz7x
GCtFCBRP1+UGXL63QC3o5Wdfj3lCSlkbvbOqVxKGgQ3NDIJq+HWytz2ozsre9GKq
Mu1nMMYVEzhQB1vR4sCoNdijXR3e4aY7bYnaJuoGwolA3tGAWS199TqEof20OBEq
8Q8lZ0VCJvy2YGFAlLtHnN4vE1syP0/RnGfGixwwH8EbXSJses0/MKjcS9MehJ87
8zsuWODjlRCCjsMic1IL8aCo4xZBga+95xlm59+onC0f4wysrmq3M8TLM6aqiV5x
KON9uvmuAVfNMHosUUvxCEkMJW9WLhAETC3pY5zrkSPps7fkGo6nXJLtLnhuuAUZ
HrPd8ODGSgEOa2K4vTNlsvIZZzLR9IIK3EqgxOETb+WxDnmQ6+FnkfFQdO8MONig
loks6GYHJBdsiOxxJ1O56FYh27ZPglriPXkDPk7d5MlkAG6vDhuqyeWKTVPyDnYO
MT/YBmSUkAVCXvNXx4vnRnFnsu4QskCITbbMOxyX+SofcdbO1lymSpVyi3ZiqelR
Cuw9GQnFyA19IBobNlfhc3QV1kwpYTpVjwYbiCnRucl59csQ1iGn3pFDDN5ULZBB
/5+Gtdr4hPwvCS6kiBYSjIPEVYFEby3JdqcaZ38Z+ZG4YE0GSIIVJoJxchprgzzT
qzHctiLpmUlIyjrUI1VXie8R9jAeKj11GL7fT70SDYD7eMLRHM8426+u3WzTXJ02
eqs7j1658uhvZ0OlCkPIy7pZtJN8HRy8oWkXn3vvPh+4NguhN72cdCG+2rgk3yRv
RpZGSlNWUTSCte6Kt7PntDTK2tz01cOMdEcquRJl7JSgCi0WIObZ2WvE9MWAyiVf
AcEXS9KTnTk7SUb1uFPwUgRVtjnhNDgWE8D/TB32K6JMwQg7l0z1p9J63t2jZoTm
GUCqrJrplh3kipbOSkEx2mCE91bCucOrdVMOstYXB+gPFH1whzdmYfWSKvb4Ht2l
3hm9CJ1vM+gOe2w/qUQODNTzNmG3zjtywrVuoli7tLY=
//pragma protect end_data_block
//pragma protect digest_block
yJtQ3j4Vd3Uova6nOwcKQgeq3aY=
//pragma protect end_digest_block
//pragma protect end_protected
