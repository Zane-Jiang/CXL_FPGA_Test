// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
smKbd3EiVdrvhmCzoanzd6n3xBRc0dGqxekYVAKdKAbdf088+eLiGSpKgUN+
59wet7z6yjADml2PYa65Hyqs2Xb+zV/4xeOiFoKmesoeiYbsb8ntOHg4sQCO
8kUVABujHxN6ozMTeDhdazhmg7Bh71uQvGETQnabSNB/y//iyy89jw5YOE8C
R60UTSwg4i6zv78mE2xynAhY7JhSxJOhwoEvHs+mLR2RT9BmG71ExtQO5ogo
NKgzgGUGuqx2YY/P5RW3/HDeVzHZ9RdlPJdC7vAJBraQ/APXg3Ab0qa5CTyW
JX5YREaHk3vQy3lQB8SVFyCB5koesfju6SRyn3dFwQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dY3/CTPfxr3HbCNGrJwMDjWP595ICIzQ0oCDNEBKyG1MtqTT3m0R8QtPBCkn
ZE4jj1ZsEM5a+KRzQdy+7LCiccwwxwk6i7SQBsbL154ovmvGjud/eoINT+lN
xT/FuUkTQtjzLuSO49SXSepZ7IoGHW769AqoRL1q87/1ntg9zHDijHPOvZqa
Xn2x7MF2M28tb5Kuaz8dkJYN5Oz7FQkM+eoXNwshhZvHXyxcEot6p1N8s/wP
RgCAvRTrn2kt59cqXBCaIbPdEhxpwWEqTGKa85n/Fc5GwURfmliG8p9ER19Z
ct1oEWyTLDVK9Lohib34FGd56KlPvoRxrfnctwFZLQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H9yE1BmfE6YV4fbpR5SNNz/7fiwugf8UvQfMcaw5PskyiGIAo/7ubhcRCz/4
hOnaZnAv1VkuKCBnvdk6sAAG7lGTzvVgOamURXZwkEks5Sy0EJsZBSnlR5uK
yzEVYRSg2GNE9qi2iJOlTWIK48wWWOA+h1GuwHiVmtzXB5ZcyRvHb1gDftDy
Ww8ibwX9vgMH9ApJKUX2lGb1b3vpooIsyxcezbqbPXb3bcn6tgjTd6Sxat77
7RDk/aW2irduKnCAJ3PL3le3f6Z4nMBPsCLPIYR7ExYYg5WFugrErUfXQicb
Kw8YCBnz3S4iQtYNh8A2It0FNjY2Fco/vWll4rjbRA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jCwBlbrufHKpw8G3lyf9TLWZpCX/NyA5PlGxR3NoyJ/pTGS+h+px1qYwUcxK
LZr4Sszl4qsyc67twJAeqjBrk4Vi0mE7sZgU/rhc6BDDo53gIMsmS3xyg+WX
mnTazZLTxy0nElOpvDySGO7S8ALIMGzFpZJV8BBTJrci9TvexDM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kTZ023OusHbvrtdOvmMdDfoz9wxeMSt8cwFKvucTgKwPjHFh0H0L0j0vOQX7
I3YUng5+plVZ8Jb4UJAr+ffRODiU6zvke/zUfW3+ZDfsHgUKCMJf6VDJo2Xt
aEM3dJwt67DjP6znsOElny+P3rYCJJ65pfGdV18I7z9lEoTW2iI8YzMKHNvE
JajhuDozKoyPFxCygfSgSTlicySNZucwKruVS79lfrkHxghXqcY45vPdS7qX
obOnwp4VPZAgb5IWDzjYJogl0dUjgkjVnX/OJTpileOm4syykZN6qfUcdAoD
dUqP7fQqOCNNqZvUa2v+ubd/BddwJR0fDD3ckiiA8E0ii7GYh2y6VifjVnA+
EDYgvf+iTnRcm9sLmLujs5Daj8889SeMlntQ4rV6Qd0kaNoM/Z6RT82MZmwY
9bOeHyWO+4EBVgqxbjMNW9ymKu1aGpH6wqymALpGasLeIhSHq0nw+2LHhD86
x6LvyqLUhkkvdq0la2hIkhr5azuDzlas


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A3cbbjW0HDdqrQklFHToltPaxSC05TUvs2iuyhbaJtheddxDCi7qBR2PxuDf
TXRo/Bq/ZZThco3PnyX9q0bAzKGWqmh0ImNVibyv6rbzzxWSBtQKV5+oEWW3
Gcgfmq7htjIu0ap971euQNjrOg6+XYnV829xAgvuTQR2RrdwSlY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
due9ejEhFYUwPhSoJsCz+golJn5LHq/bUdF2yleRyp1LNL2dXVHNiPqkGBWe
HN/CmFZxonUm4aXG172pARKYb5BvswHGRmxHcZcHJvpZbySjRhFgPtF71ZuC
0ly9PGebYwByjdroy2d0XzhAE7jJhOKyWGRvuClDxwvs9nWMfYE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13072)
`pragma protect data_block
WY1C+cQ+p8C6UbX+4wRTge7+T8IOYZty6yq3I6xZCV5Badw8R0ubfrn9Vpgy
JDA/9JEp3DKiz7tzlkDvPNL8ETcNN3cG4q4qryvAjBurM/Qh332vaS+EyDt0
jPRdY5a1bxvMbOTulIcG9dq/7JJr0vT19Www/w/F3KeYLIVDh8h0y20sKBZG
b7Ofii6uNRM0nZ/QWfEsBdhzO7M6CWoTxJFPoZ80G8wxwt2+bH3JZIH9LziW
RDfxxTISd1Zj9HFd7nwUpROjHWOCX+3HHscI29p9bcUAewWU9J/3tJqZiZkI
DxpvpeRvWUnWlndkS2iqlRJXYWrSgI/uA25CsFWxvU/IAwTEY1cYmW8b+LI5
H2wkvzz6kmKGNo1HJwKfMxV00IrUROsTkoUJEk0j+oGjl8Ab3HnNvcVsCAyZ
QmpE+vzZUtB7jPZpQ6rZxVio5jNmoEMzVwQ5Mka6XANjHA5GJtuAjhfrr/t7
b0wuYXvkSdx2qlsAm0q2gOyYmKAJ/4+uYLHFbWsZRbYWft62BrCfbWypeLTD
V49VWSyMXPRhS+SqJWRxiAU9ZONzraj+Tr4LcLmBWa/1rZO7A1Vl/gAv42wA
hDM+XzXverhnQ4SOJ3u3Y8nxHpwpvXICGPutibukBZNYiG2yA5nIcWZ1S8tK
R/S896aYqNpTjBdCYDRlNdWwipXJyy0cxuwsAOmGhYyzBNzzF2S9MXFbG5MF
X5NsTqUicV+o+ZFEQf2SyBmwekA1UyGf4pshvGIPZbrlH6gbCvafjxayslcN
pKJa9nqnqdXuJT5gZ+tOG2yauzgfELktniXC8kyv1lFYyJcJtrL3EoSSLmHn
Fgh1dI5t6WfABcbpiZga/Kx10z452WA8hNAskNCdBsuK1bx4bOzmcF0xvQLP
Wd3QQkQCoseRLC3H1gBvKbYKPPphWVi317cgBZxRXnRHvqChztQzzxDFjX0X
GvJTr+LdgnpXJO+GXD4frR6tqb+QbnIKvOfWRjcr+gmdmIavUl/MJFaTemrB
KVF6fo9jlwc58o806EM1wKe94rPaE2YXAHKnE1uds23Zt/k28eTE+u1frrx7
3OFxCjru7bjdu8A5tkI3hSgIkIoTBxNg/T9vwLf3ylZmciVTuCWTDS6jhPil
n4sob5P1PsahYxHrQA6d7Tewnw83LSrgl5knNX406rMbbDgw1YJ/AoJmbPPm
Q41t4GslTWzfwLVMbBmuwCXMTlLK0vm9OelWBkMXFl+gB5HvF50JYUn2wmx1
yrVCdIJvPwuV6m+Cdec6OOhwJI7wRhCbDocRnzt9YyUESAfkej8ORX3u/e6c
v2diuvlOkxIRoZ+mmeKoNvprGbSNMGlirvVrt+sZLoo3ywHvMOiUIlSiz69J
9K9lbIZG8+sYqSsJ/kYjxxsCKHnPa7tRHLNr2pK8QtvgkSZkAuUni+JJsddh
Zq9PYPmbE8MiPjh1J7X1xQwUwEJLnDmIu782ZVXi5DbyuARe6ybtdA0NZSYS
2X/gqoM5+/Ia/jZ4/mokDM6Z+FrxNuA7R2Es6JlDva1UOk2Pcvs7wVVzVKYx
Zg0NcWlO64SKafpPr2GcRhHRd7sCMJQMuwsllH0Z1TLJZ0p6UB3Rg4ZTO16q
Qh8DmyTmod/82KJztR0yEiKof8t07k82COmNGZ/anOPO7n57R8mUAACqz2pz
Bsxgjkzrell9Fq1eA7meeeYpl6jBGrPedWVnn2nuvAVjpMytjc8hOsXNGj4g
HSe9HfDakueJACjbGz6mUCURTnRUhsxgF8qe816mBn1thaqgmFAwlgZjDswH
mZmqdWFP73cI1ZOd0asYPlRej8OQM/z3CpaXCJ2/ET+P8DcHn7NbUDXyTG+X
oi4VNEmm6ppjbMuVgj2gulP9BXC0lK/aMWHyoIzokWXCJNw/LwRZlawGqY8n
ECdaLJ4CwfYKcfJoy7eBpKfqawogdnXKz/g57Ac2Nfrlwy4j9hgZzRJa6JDU
jFNXE1Gsp7ZC1UmCnxiZU8HqAedF1hGRyLEc2znrI+xRDKwH487SM2jFi6Wj
P7LqfIKCRjUhe/PjQL2VGvrlMlNn4fND4Zi+64S3TkDrjDj9BprLVIaJmgcL
7mrBYabWRfMR+pPF9/nFarajjplYurN5eL/NhGnqVsl35w02EaASXbsFk01a
yEMLktlnh2ft6zcqTdS4d8h18mH+RIIHwKKUfoHd+aobAcbmsg71woNDWXsw
ynOhp5swBFPoEr2Yi/xhc62TCyxIM8qEcNyx46R25GT7jYaTn/fxz7k1CDPC
FDOCTu+AwvNb2iPa72jg/p9uoXPHngY62YZcwx556W2Wb1IYHuEVrOrDqikX
g/zl9F8ynECyzxOoURKp1DHKi6anRFig+LeUmdVuDKCZBc3kkuP8BpVE1LKb
FLcybhUuXTka26ePxLl/hUmS0rvYtBnMUI8dv7n3jtwIbnCryo5C7NsR34+y
ey81v91sp+Boswt/+EfxjGkTbAthWdPelo51muB2cAoTeC1C7Zq0TWm6+1zo
LQ8x1YzvCPs9ZYmV6m4wQe7PLT1gHt2f57pTTeJgdLrcp05dCXSKeTWkjZh0
VloLicb8HTMvAXex8RRh20fl90TsjmAIHK+zidwVUPBbNfkvn5gaVZ66q0mE
jVmk/SlkIirYy1jJoTuABKAaPMnocxYI4MsMT0lsWqKqhSybI0GdhOGZGQ3j
CflxVJ7PHZeA/0DHq5QOXYO6w3V/p7kCvZzjyj7a0HqGWzgOuoFhrrlipZ9F
+M8I+sfHUGK8eLPhn3w4gu4eqF7jTxpFOxLacBC+x9rs5CIrA3QoOhbMltlI
SE64W8/FSZFaVPKmeTd/+6cyYpFvD0yrGbKOG4xAw6+oXwTXuFwNzYsNSqfM
iTL/BGXGt6dn5f9xFrAOKIeN/dWbGnIYWsiclPVgADvjiSVr85j0sQE/Gp2g
WbQgwLOzoOuldTof6saw/CzAo6NxUBh/JnheCpa1/ZVWPfXXXN79G6ObQD5w
Jy0dq3oCb97bZFZYWZEB1SUN7RJeBlyZpVCEq7MHeEzAl1OtzOCD3kWrqPmg
X6xwuXHwvIa121WdVUqkD54qPqT9v7yqaTRDnLWdSngvhBQaPoWkVB0OT75t
iDQzpbiYW7W1rJxSvs6B/1t0QtMB3z1rxmZKTpi4/IG2+PPrfXfr5ZsfUJDf
SKeYcKhmEApNYZ76fGQWwzQxZmEcLsdARzk/+BbgYv+0zIoeibzfS7vRQ2Nf
L9i6VDJ5SkevraTUYp9nJWgKisNX2pqJG6GGE1P/8agN6EqP3UmGdSB5aEc9
jDAKHzYF9x49kGnz3/glJgrazR52SG75Spnx/3BYqbNhr97vToMZGZZCwOY+
QmzhZEXM7+toVxLM8NCRHVzLCfDUhR29Ua/VNW02SE1YB6k8fZfPAMsF+QWa
nPj3ctl5kFhAmG3Xy907PcN3zDANmQ9Ts9Jw6MsXr8PgEMWOSd3X1LMGNMCK
W4sHLQ+yrA3UfdUReopYL5ShyB35yFUDBxjUIEWMSBL7tCWqz65VT/qHJhLV
E+wQnZF07HN77LF7TlLfk2dDXbPbkBI1FYBms9AXbZdH/oauAwV8sFdozxDM
vX1zcyEB6JMJ9oGxslVySU2pUtOHlV5ialKaI6N0sOqQIIXTx7bOdUCQVQkO
EGz8/1dlGOVJJH1hEbgQKu7TAEE2dC0dfDCpwGcHq9QOb0Kfral6hdnI+pX+
UNZBiNFobS/EKZXgRkWnY1lLPyH7tarNpq3e+tbvtNp28LwQSsiKiU+uGx5K
3qT2Gm8emD1jzKTO2hor0j5i4aODQpcHOtYLyCrDD5UfZSxKE03hGb+IhMEG
RD0lqZRk/ADpI4AcJx0NbljwBuKlk4Dsu7odZxJzPwOncPJ1OpovrTV0zF9o
YFuz+Ec829ZSH0t/IePQSmw+2irWQWBncYMrLxWtpcsTjYK2Ikaljfj/LBCW
7f1gFMtNh9eqBE+rDjT8CmIHEPfeM0Lq/fYrsyzG66/gYKl5g+fLechncd/S
Z/wu1aZYrZrSgZ2prxaKP0YHFGs1z8lFpCBwOek9uxDKRrBdaLRGi8wZGKOk
boYEpLBU2KF98eAJFLI6tMzMOtT2Ud66TwpkgQkSwYZWFwbELrjVA90zdM36
nkWApIHMktkLFu0bnx8YuB8RU74B0UzI3/2z4rK508I8E/csbLtqQLqiUzTj
Ci5uckNxRQEKlkVnlcZNhtL25OD2mlHqHvw24N9r8ubEJvGISBJjx6AlDAV3
Uc2rJWRnSHGiueMTwHpDiyohV7e3UgOrPb43OF+1mmbI+db0s4IZKNSAio9N
iFyav3paTNYppcpzgxOnqclt+QSnuoEGXJQfe04Ey2Z1M+mGj6pcn9PVlVpg
F+wDTqnzY0pAmCwZvVm4uFAFbzzwc3DeUj0kh96+QFE9ppCOUgGp9QJ2n5ca
VONyQ6aHWGUD+6c6IDVAGgRLXcFUpYkbqcR1oivW6ko8d/dqW8xsXI9X8ECn
ViEIJrgmbd0duJPV9dchK5DSmF1xR52W2O3Zvkk8QhvF4q0nkH1+X2/qE9dz
TgdQiFmy2k+XxQhW+P+Ebe+6NpWon2VENwLzEvtVGgyqpxYB/8rkcQs0VilZ
06MuB9iH4E0DV4uQ2N0NGzc1sl3w234lbrc3/Z0/ujxgl5MqSKzenligh3Lf
pwBMPn8Ou55pYZH0pHCxiKEBd2N4JDn83VA0A/uBIKK69sY2JCHogAMoZRYP
8sTc3nzCY4E3ir6QfyrZaM9dMlKy5iq9KgGlcT//VkeS/wYXdsGedg0SShDb
nM76IA3eMHOMqA2LzcYOrQ+sH8bu3NUIBF4rAVzW00jigEAbiw7i+39D42Ww
3hngRmbY6JZVS1dy4DBKlhsETc/qeqxtnD69Len96lwc0+L6/rsD86Rs6Sxy
rcj35wXpY6EVpR7dr/1jgUn82bScuslMmcbpjKONQTO3HCYybASwZK99sjBe
IktaJ7GAHN6tYAmp5RfDnF79vQZYXK1rHG3mBIaPyavg46h9YQnaVjL4mdV0
vMGJVEqbV2NlqHYHJ9eX1jwWYZs9ZzVrLG1z6TqZIDGwdDpfIWd8eLclafV5
5zdiVlSUQUveITNxo4vPq0qY1WcSBdVbLoyhecbgBGYxcMBMv23uXTe6Hg5R
ukokM7QRaQsibQXSkDWwqcqfpCzi+iz88bEA6+OX4m0nBh5aQ8cqB8QYT3qH
XpskjvQQdng8Z5Or7V1tBj7uEWYADX3i42gM6vfhHE4Qc9HA9F8fZwKBLWmn
9AtnEzru/1CkI3G03Gt4ryk92ChysR6OVdGTeFeDVmdxUtCR1fM3iri01FDX
ZEJkfZrDANQL1+LJJQ8zRLPBlsyomw6NBO5OdC29KahErlvr806qEokO+y2l
fBTQQGaPxZeC1Ehf8XFutUL6Ch41ObbhNlblbcOHwNby5kxbN+ovirhsz2dL
ES4pjDCbhZwG5mZqGBz7DbOLWto7j3pZt71FfqBkL80x9w+run76F5V7ZKYc
voHp/z3XZX2+Jo7DWis/cIX0vuC3Lf1ZWdU/0SkKTnbuj16lAjS+T/WMtRLg
Lbcv3jtNFz8SMTGdGPlbSfTKc2nJpM34sBrSngc9MUFYUKeM3/rc61nuyAD4
NGUnChH9K+T9+dgdRZ9hgtJG5ORA250VOYLo03feYZ/ivUW3TR/pN5oCRn2x
jdkcFKO4DOBwgIDcfsQCDSlufYI4SHU/wGbs3T7WE9IbYfAruShVMlIqXx9O
sDHR9nlJTmWJHdMiVL9MyAJ8iZT94JiUkGsMdi8cBReAeNFA/kqY6NjpPHUU
bgPgmzZQ9uj40RBqV61P5nh2t0s4iE9D+NFeqE60pj2ompfIG/ZhMMZdimhl
+8mrBKrRqWt/ma0qcsw0kNZU3ZK6Bf25hC4ekrB3Zs5z1eJE/nPR3VT9e+Up
iM6aXhchLmJ3UEebbCDxGUcvzQ9KVd6C2V6Fl8suQ0POIPgCjzumiaCt8IC8
e3UISwyNul8fhPM8wfYkuouJM7vb1cisWey3b+J1KXo5Cd+qz764/EhAD0Qu
I2TdseuQJalN/7eA5AGtiNlJsMkR6w+Wc+V05kygLVXgiH5Ei32ghN99vMkk
2oEXD0bKgUhfX604Zzn/oFe0NxTUcCBaNRSmLEnhA+OYWn64YStsCxAi6+y6
MNpuegeqj3txNEy2kbi96s5XTqTAx3YXMwGHMuR8KM67c8kOu2AKJvAXyr4L
75o1m9HlSRF1mUvkvpbDDYwhauR6jFWvXAV2gMZeLH6k0CrmWyMmmqvkbtyq
YDbaW6ec1I96JSje372v62cuL5O9qp3Q5qG7402hNEgrgdZ4UE1eEBXAoMSU
4ihobCDRwrZCEqREiRU4cPd9gFcTQks0355wvUwC7o5h/67gnHAtLbXsBruC
ECZkZsh3bKk6RfAl2EMv6b9Idy78BtnH/JZoLfz3FnP6tTGqCPdkkzdL9/me
t7WfZLBgLhNx3e3CG8pekjrAKkXMxCXuZo2I2Vf77lqul/D2sxUhGxs+G9pa
1p5bvJeZhVGV77/mb5nLF/JIGPI4EA+0g2UMzS2O7v0bFFiW8FS+DPZPzy/q
a/3Q0UbZcQAcHFDXyeB/VYHgO8W/Sgyk7SqvH9Dm0etM6BWyJzHYhmgkQ8vQ
wH1TRp7KgWVY1cEFbN6hugL8LB4YpVU2jIQIEh/cyRrYYjnKIr7pO0u0egNj
mVutWy5+GjDXBmqW4enbR5U1fpnTT1IYcMi7PBZXLKH42KN9fzfXjK9PlYQV
6yXmhC/cAMpE9qJUITMK1+4E3S+wmEXKB3w0ppXGX4dn9C7pGXsgUN1ggE0B
g8HrNSh7BlUhWFiOK3cGsCaBedddg2pK5PaGsU+WhOZR0HbBDjJNVODJdao7
BjP1Q3U77IGUzNKqCRJxGba0Qwk14iGP+sDeTYVVDiEMmqdwYmRIxNzrKtXm
72C8KfJYMPuJERLCUNrK2xNXoxFaOuSOxeu2g/B0d1CLMrRbykyaXUcpp3rP
oC0MI+NGl7EFu1ka5ndtd5jcnnSe1/ztbJLnD/Cnp8NM+oYyk2lTmspOiwMw
7/GjzPpefAReLQjsIY2r5L6BoPll0u+W8ttTW5Ju8PkO9v4fQD65mMj9F2A+
tVeuN9eP5AF9K3v9GyE79lFfB6DY9mAVu8QfKQf7eJQQyh/w43OB8Uwt8Qch
Ex4saOuj2m7YQ3hXnhN+H30aC8thzqOCUrUCiYy2GCTPcHIVwAXjqFLpcEWL
+kLpZgU6IxdTQWG3bGVlHSDBL+efY7JqK259SsvNo3ge8N3/Z0t/6Ma+Wm7v
qmYdIEaz4VSailVSwOj+6xB+NMJ+/nAEJDYL3v7fbCLivEo2sRK4GssDb2fw
Q3IUv25fteXwlaO8V1DhZHAUAyH9i6d1AnN70yHh9SHQdf7JBnO9f7KCtdEa
zjo44gz2B9qBpz7FmBJK7YkmB5jqd2oV4p1WT5mi08Mt5nh1CXuQap48eSSl
KSnQgSopsz7ICxrtkuXn3LLCSV+yymwb2PMDIElgbJsuOzmswwtvlFAPNSqM
jQxAZDsjj3B8Nfzdrq0Vz1TT7XbJVJ69Pu9G0EhaeOm/51oz2sTc/MHApgff
GRRqFKDPGSNnnE4vy0uPYMSXsRox9/N9MGkc8PI1xG28ZC7UHlllkB6I4vBd
6IUVIrpTE9TxRAMhg7afhhqy/pouhGpGs+MMek7M09C6hoEq2TM3gnswHOMS
Ma8h6zugXq087Xulj81YaHkC89FGYqCexK80yXFQ/0FftJdXum5YcPibr5Cf
1Sy1Z/NJNJtEpUp3BRyxUFrwVo69S+kQY2tXRSpe4pA7QQYcLE/+yy4fsX6S
d5AznwfRrErb/DbpwivKQOsOUVX4tD3AkrxihAMlWMKEtkA0uZTwVehxIP4d
S+W8SrdNtGMhQEeLQCVwH/xGytGNgmLLrEmmtTp8m6FLWwjIwagD/0llGdjM
yBVqKs3UrEtpJNAgOQNCFqeutiRoO4KZybJEt99aHL3y2o2JGeLvhwO5qN+z
KHmx22P7il9IRXsFc3hoRTxCcS9Twg2FMYyH5ZD09LF5IM0l1Ffv0IYB019f
8JTj0vBGTxeADVCS0la2aHpAslgtwO1vtcvGmpawap7d6k13j1Hz+bDOBvqb
rRzIVoyV0M3/ruBWojZr0y03E8+Mb7goh51Dntwd/TC8nUjeSp8eZuBJkwBH
0IpWJSIN3q913R9tM6GWOS7Co/Ho+vjhv24ApeAap28uxLJqd9QZGXsKrOVC
HTuc587QNul45N0FBUUXTeNlqzRQbpfQazHbEMglqy5kSohiCVZQj6qEdnn0
s2/KnYJKlm9HD2F0pzcO3OHNBcm66BOcGe4IR17N3PA48SsNILG0pq4F1AVz
T2juhoYPooyPy0ef75ZhvsSUd3y1zFfNccF7F7z1nFAh4TRt3hWpvzblQCjj
BTglbc1BlaKyt6kr/2zIQpEMzp9sLZBIKMdxR4UEGgSL9EU5Q4NDeKXyWszk
K8u5yQXp9qlSQV/kBBZnTdEnGUAqtnMGYjs6HIv/XXdvhqr+9LtkZQSPYiQs
fDnWbFWo3dWNDZ9MR5BwWzQpEHuCmZo/sGuLjhzZX8iWejm4Ebxf+KFk7OsC
tkF6pSBK3p1NgzRzTlgSUyOJ06hp/2nq+6DpfvS5Sda/Rjg0DFaWE63gDQQZ
AXFhXb82VJWpeCGIvOb/g9spIBqWhR72nnmZN3yNdpwB4Z/vbT6U0N1ItnPY
i+/5YbyQX8KH/rsk1GgzxOdmilcp9hNBEVN4cX+qY+/fepExEkmjO8NRNHar
SfsW5zbG09UsC/rcNryne1zydf1i3V+SqPdS2L3l6FmcdWLNql/PBUsOsqzl
RKue/0Qrn96ChOVSEkUWUNgJ9YzQ36NJfR+K4pn4WdpTnx5g0r1gu48ORfW8
0mgp6LaDVv8lT0ahzFl5mX8vC2qMNXglRzj1LI4MLsbLR3qfu99qg2SEhFOD
UKTw7EUGTmvnnr3Of/fbzgxWdDNHTM2vV8m0sGfkrUzqgZtfgsT9hAgNw/xK
aR1Q6VcueY0M8ClGf9Ip+J2Kqj1d/wZVoyXD4jhKCEQmqVIJ3DXh3ys8ifSA
2/0peNuQ31TlHtH3VIZ+NfUwPFcS15uOSBX7nWvWjVFohBdVdK5FhegsrvEo
uxdIwRIT0tD9qn0NDq3XSSoyuMFrD2CRI7lC/fGCszY4Ol+xUaCI/eE1q2M/
yhoMyyNGulBv6Z7DzAmwGWOvpAl5mLPwnKyVIfC+BPOsgRwTQuVJB9f37vwF
1xYpsiQEZM0tqksZoYqAS+2OcxQfBtXp24063QdglKpK9W71IHpt6xtNQo5N
MOJlpNGzbZKIW+b2qWMSyvEaN2x82cE7Kz7V7qlViVeGWMwmskpstzigBEE4
bWzD0A+kRH2H9M12kOpFKw0KJshsT5huMocZ+4EKNGGDHNpVpSKKYr6qjFr3
7mGYeya5CoZNTdhkZ/He4Y2gg44WF+pD5opOhgMorV54EOxDaQc52klLYfcl
rj8w5f84PdenG2bLfgLzZC0tEui1W3KRPWbgimi9BGgTH0HGkb0qDBKwvFe+
6dxul1TpZsFgg3BxGgJp/1F/o/Of3r/PtjnO+Y4T5uefGtuHMD8SSkgr/KtV
Hs8p/oceodAyK6aj4BV7x/y4nq0RzVqDSHlSlw+mGzWNSL6J/RyVksVi+7d5
XS66PoFgVWsNtRsr9o+40Pt8JLIl77ziH3OifPO/ZRaLjLnYzqkIIYoNCcP4
SzTFOHnKgRwTSpOk1/PdqimXacq/N/pmJAYg1W/McyosXhistjYlKf98Ytun
6LNDSupZG3zRTL9M7i3i3JhEXAq1OjvN6JihPyUMwurIvepwVTOh9zMPwPXP
a6bR1OUO8lsZV7/co7WfZOSjqoZJGb+z+idXQPGTvD7EIbkxl7ABonl6UXOV
sJJunfLcp9uoUQsohknjmyYtLWo+TQCT5BJmfZwGUAnWJ8I5z+Aa34X1Lmcl
JJXUZhILv23oNtk2Q1seYtGDHzjJYoK37fXoLcKCrAdxRjbkWHnFrfCxDG3g
OxO0szD7DR79Fx6F/Uirq0Mjk0+j6uhklcGAkH4sw4ldbMSM4vntodPInvi1
+zu87pLSPoe7eQziv1CH7jGGOvHftk6F5nFbgeduflkSFOfz/OYy8z9eITe/
17jAIs3BLAoZB9DRknLeWJYwA5APxfm1b25dfCoiZCbOb7uSKGpIC1YRUOCj
XESe0mkH/yid06bZKbmzEKb+PQqUbUVty0cMRRhEUzdGi2euO306KsvcL4kk
CoOQuDu8vwJIiIWjvpn5EtkJSV/hKJ2Tb6RjwHS9UoSiIMbZEQaFtOkWMXY4
5WZJtrZP9V8Par/MlKJmM6ouSDyBgKklR+6rHsFJDSzuVZRxoi/GwUned90Y
reUykagzUJwKAWc1tbMnqICi0nxiL+zAH/JjxRupYZWZHhgomLnQ/lGIf7ur
5k8aG7YMx+6ziDPCpykhybznWIlj8hVcByj1OGlr0a6TAFQ4/6yqWWPAqTQZ
lwe1A4H0Ez5qH4Y8R8Yp98CqRRHB5DJUUFkt+SFpUVrB7pmdrTPQRiaGi8HG
Kyy2+7lS5zfRhfvzwiYp19QucGGtFh5pVeKNo/UBvIt4HJ1zwmjUqGmiQu2B
VykUOjOjCb2BBcJjmy7Du3Y8sx/N6/oGDILmfIRNcLvqbh1PQcc56IQikYqh
ATE/8eyU2oG85rB1FHSGKGoQiT0xmlFL0CI/vOekVPed3fhrggA2ES608K+w
YTPSpKSLnLAcjK5xkx9OFHdqM8GsrIMCScvGWMDkRE5rq70whpIJ2P2IKpyb
9kxjjrc5BuXGouUNpTD7Qheex9mCCHLWx86I4oKzuBWpb6aIrGn8ibLFU2tV
+L+z1UjUKrW+y+cjB/K/I32SSII1/VvMHgVfenjpb0njxNKpMxCeHEaX3spx
sOon4X52TV4i0exY4y54HS6vqRltNpxfDBqNGpgKyLl4sERMgNGQYPg8q/Ba
BS3cdDbyc4TdJQqkOxt2RRMaZ3fct0XcmtFSN4aKgAsB0BcJBxttjx9mtzSt
zWNdkj+IxGUTocEz+DLmABDVWXgcHLZBlHcSYgvTcB+AbcnX4snb11CmR/9I
fzYdMiuG4CBJUkESNDQRkRqWFlQdou0GO0MDtIJMPk0xdD24wrWk+THpHahY
LA83igdXNqd/YrwIxXxPKhNPTjl14Ewf+cG+zHBOIeEnAFEUTuMNhOJ6jdLY
NZovYZuDCqMwUc0GsRZRJmTIq/kLECJ94Iv9gEju1dC1A/dnzDm8o+Ip8cPW
4+YVYOdYcENkYKZvkL0pNJfWQX5SWkH/Eof/Zk0LgaWg51hDGJBa1Ka1cx/H
LIJIWkSC1DbhbXtBzdGKnR4ArPoJfSR8Y77JsOJyP6QIJ6+VBjpVbq/t8+Fw
e4JfqpxklxUvBDtqiX18rIRwcH+Lf7KCbT6A1LpHbETH/pnuXJf8rTiYU1RB
MF3q6eEWsCE4zP0QlDiFgwz5NIePsPGRVjl3jfxSnjpvtIuCBr/bK4fHl/N3
RHfQSy+lNzHEy/R9z24Crpu9qqYnJei/XwZoV4eHVFu7mlnrdPY85hJZzSvP
GW3mCwmEUzIOV++ZebFxKw9Hn0IZvlKRfgiIS8L3FVhd6lO4OsZNuXJwRbg2
G3nbF9z/jnTupuTZ2nxnDp1FrSNJ1G3noDpiNffbHigPL8iVueI5NacEPqUl
ajsrTEFZ05kJ6WC69TlzXPRnzzp8bGRnO/L1Tja0+laryXNmXl5uw0BvEvcu
TR1uqhgtkLfU6E5wg8iLupjL4xt4ApFbqRen6g5hxZNQ0WU/IG8JNxsiOifQ
koGXMqOoxAezoIPD26FhyH9y0jpswfAA+t4JXXIN1NfmtRND2xNCPrDy6DkV
Oum1IEvi/ntWxJyya7EPSppDQfNlLI851ENZbp0UuA7m+dDfgTVU51Pp24bx
XY7NmW1JJDBYdC0MHivXZYqPsba3AaX/PCNEtW/olf5L6D7CccQBK5cbh6YN
it9myZ29dnJKIZDS2vVMDyy4puopMAX4FkjHGgKyXH6cPWzgVosnorgxdbwD
b5S1PuK7pZl6H+zmvZMST3qArVPxjwzxOoqsmPYBEqDXkY4+xDmz4IXUc2lq
mkBvBjPxA8bjHH2+FF7ULdOR/PwZZwnzvdYylyg9qNhNHiykCQ/PESFwX5Aj
wC3lm7UBYkN8seMrGJPqhffghzGJ41TlXa+YPIUeDRrneaaozMsVeXxbuABl
Z+OMSv/XCKk2GlRky+Wcx+VcU+Svyx8oxPT2c5v8eWNeog/XZEuwzEzQcOo5
GpuYBaJUVmHv9mIKNK3nTnrEooKuUJ/FTYnkZ1vbRcP8bGkO2oAZNkJgG4Mg
0Pk4CoYrtDT0+m4LppWs0Z+b09vDJnXRxYczzbbj00ijlARSZl4sZi92SmG4
BCnfZQ78pLFu217hhc/yvR7Rnm7kO2Ys1hgnOP/fAk1uQU0TieMb8T0bN/Qq
MuUObKCI93Ih5wkDWO9ErnzjaE16FwPNMEfgXWPMabLfHWq5HCVIzcPeQ9hH
1aiZlIu34Y+TTTKDQPce6Rbb+AUo5SXVpCleZbtGLIhe2MF3LLmIEhgkD0fv
qU5gSuhe0Zy4X1aVYh6CkCvfGIk0sv2CUfqgTWaNouF9f7HfZCfgrrbzsifz
OeBscu1TbUR1gaPRpoB2EeMIf7fPkOzIpnS7WF2boe+yPAmkjUAfAPbK6RCd
cTYGL8qZN+GanIynz3c9Iw/sVLQhslbZyymT7CQmVSB4Rxj3NwVQR5ieLeOv
5uDn3jkMA+G/QBMJtDJ1qNEI+zJf8QYCBJvxhS/dGZWr7NbH1yvqMTsE81aj
gIaq2iOHGLywLN1ymVwM96WHqH1XFcqxPz9E4aFO2Ye/S7Azhxz0XljPsnjW
KqDTy7kaIKRA11nCQ08nfM3MCibQJyb9rGB8t2cy2x9EHgF/srN3V/Lbg3xS
nz2AFvBS95TTYaQHWU09dY9WQNYZ5vDbYomdzrvc0w1AEsyORJkQbC8oz1cW
Jg/HGwun9xsuDv3wwydzDQKMKZDS3Wlhmbr1pv+KbT5eD5Da4C/LYgn44SVu
kv6YFR1+gx9xkKi8Fs63pu7hCAHgbtxpBA6JYxQ2nfEHMqiuf1i8j7lwh7VQ
/ueFLkH0YaPOWRoNaolAcXVHpDKDlcuYZnZmCQUui9G1sNt8Vvn55+viC3rR
zKhMPv3TNbuaDeyrlqTIkR9fyZhrHoQFCpVe+kJFpn32zahHSDUO1EdPca9l
J5HGXhbovcG4UT9xh7iMa5sJCUpJdbHmL1WIA3EutzkODCAne69N7lVQvTaF
R06Axmhbp5vUbjIg8Zrv//RPlHGLH2Ed2TkG0dvQDrwVNf4UK7CXEAfC2cWC
DY7Cq2Z+edjYfjb4OKnZSWXiuHLkwYnzhGZ6BfI/OyuSPE33ynVTi/twshZe
C5FPOvulKyIk0KtVn36E3T77AnJI68vTKTLl/MvnZDRpaJdUTWUahCXZrrKJ
ZHhpupbuLh2j/Zh+0uzCHw+D9UlshgMtwXmMP6BbLM3BkaIP9+vzuCUYoVaP
6XmkrNZdTKu5NOxzpuoZSaTlaIUqNXp5PmxlWg+GTJPXVNb5KER9KykOjOej
qTBHKAU+AT5m5CJe1dGPRxefDgDOg+8cSPDzJ2vIE0fZt39xnwwpa58yRHq/
3uNaz9sTgR+rJyQfaqrL6z5eWOq/OSaSSHTlSgeytcqPwtBu4OS3jQ3SrWs0
HlxHElOI1/1GjfeL0HyURFQqKdWZjRWlUf023EY7/JjVekROisod8+rpLVbY
C2bbtMcom22XtXZXrS4NKMfJUyktJsEsnJYb0RSALRsiFO/nRRtrcIY0J39+
s42ClssaVBx6fTfEk66O6zt8P2X9/N52faieI21k5BBgDkCwcQSosLWKt/fK
LARgXGTJXxoEMKLLCCMQOWU4HjrW0STUXtEbyNnJMgk6dMtdclmqxJWliSty
2eLCW2nz1n9SnQCKNeF39HN8VKn0A53+f2AUL/pzRI8thpEjsoWXC3Isz6xz
TZDtZmn2gdZcHQk+0/gsaOJ0hfhVHuQ7TViASioxRAsB2jQNE4PNl3GkYY9B
xe70wBGfSccQX+mFG8Rbxbq9WFRXa/rD++RE93plYXJdHpRfMccf/leWS0Df
XtKJsYLovieaIgjAPmlUcC8IZv1qfLn42UkN0ZR7C+tzRpKTl0tcB79D8uXY
bDUTcYWT3oDoFQf0M0GYIVSShJshlDdqVsO2OavV7GQ3LfCLffduSD4rpTXm
bGWABj+wgNfED1+a4Ax1/tArUmU3nTujyHhdH0OCqaJlYFTCXtLTYohMdxNr
eHzArNOPWBEq4e5Klamu6y/YvdWVmsFeUOQAbW2MdZ/zBboo9fFk5QoR1heu
nTDFam85wuCPIyHl+qKice5ZBuNCILbnxfxqrWn+/2pzSNFOpx4YeexPZkZU
beL+arT2Ai88GC/o+VJmsmp0MWh/f167BC8y6Hg1rv911dzBDMQdWy/q8GEK
oRMc4yRzCuVL8DGebgGoFouuxaifm9jOjDNM298DtLPlzTeAtDA2D/dXsUza
LiVSqLuN0ufr/jopP+ON10tPFKEagx7ld3pFRW1rko8PN+ou/GB8byAbAivN
UCD4cxVZyWsm8sj2UYsyLWpMSUnuc10BTBLInBOeHpoQaK81ja5XZwju6Uf0
GegXbe4XdrfSsEgaMOku5RmK8vYlXy9eihoblxvTHxleQMk15+2EVFknOdKq
GDQwuFxZyaKG0WZnyDnLR1KVMMgy+yC3t9vj+9DAqzBNCrGlBGAjJpNRpjTS
6gLHzjKxala29BTiAPz/H/2tX5U+wxGdD0vSDYgt1TJrbTbaHaaEgvWFcsQb
XwkTht8X4jZEqFIJtAKyfebIPZrN8YKlfFQ4NzdkmDe8N+O97VSnodLKCDoY
W+LvOx+GtjmRDRSZ+I4BXwoASmivQhFY/XTG1h4VNX6byN3nFdwRnTphh8D9
x74bAuFj+yZbZ4HnqEXy6GRiHD/w5onFb1syXr8gQ1t203xn4xC3o+HF8Vls
swEJrFl7hqRkwo1Om7O//JaxduF+GN8OHPFnWIApOZt/ruKqxGkOwN+I2BrT
YsnSy8nMd/u2nBQUX9nTfuTGqIoGQfEJlxmV3E/gLFC/C4B01IgkF9WxFJAQ
l5sd+gb5FXUpTZlqUowQNibZ3RDgzZjtanTwokhlyGWnjqgbW2XyIR28DLU6
cJ36uHE2TvoPI8DkJb39L69IKj12X0vjgiYukzM0UQuA+IVQPN4KzcOg6Zt9
eROjWbtxJh+kwYO4W2h8V/my9F6XF3INcqMcRCQTvqEudK8XchhJ/r2n3U0I
ESTz1uEFcM3i69s1WhKszi2tc5gCrmPPzyZrCZAtmVAvoe7RzcUkrWbsXbTU
ctQwTcUcJV9JQyQFm81/JSNsnN4LyXRDrq//ijFZzzVQ5lKHs7BmoPBrcDCd
tKzCSfYbiigyuynpc5VavptpbDQGkzX4454wW8N/412m7UHImDraVmhVk53f
rhd6jmzgyv1fVSNPkSlW+dqwC57cwICrRn8oZuqpDyG46y48BGlJOWn6AqEs
QujzuHpIhlElouJMoNl3osfLoQDWD5y8hS7X/jA4TGQ2L4a/MeptgaufDl7i
5dn3GtPdpdE10FXjt8zzwVldA79tUUCJFuYCO9hWY1HmDYXs4FJfXiHK3W8g
9ADg2vppnhIY54IQRgcFpyEK7ut1Fp1D8zEzWj8rspZlaxVgFeFJjqB51u3n
KplH6yhnoydoj/JHnplkbVMbyqk5M8t1Nb9Y7StAjDc4sVkjdqK3q7GT/vKI
acTzyqf5vDDu0dfdPb2Lc6/i8WoVmhCM58sT/Doi9BpjLdELZZBPhGyKm2fz
b2c+6AnX6Y4mfolgdqfdGJvtEF5wYZeXlRvIsLnKqrlVRztBmezMk54SBQZI
r+YAlGoM0FoMk6O/Eh8uTlvP2hgdRqvAJpqVemnJ/w4lK5aFdJ3M7GRE2+16
hJgtXRckd+AnvTnx+5WX0dxPz4rdrOiprp25pU0p9WzkwQhVSujaZgJxvxMm
HzXUcV8xDqgSESO7uF/2GEjrbXM+RfI4LuoMVA8nYwjZmS9NAynJhdN+Zuf9
4LQYQGxGwSutp5M6BsvElVWsrTVGJgo5emtu+McZUGf4+DUzpHa6/9xpQJ8D
RQxLiYqdqPBz78uC+YvSwW0wdL3y2TJCBZOI+k+KYoFbI+at5m5djddClj1Z
9dMYbl7MWNyjQDrl8ExIgzlDYtflQG7nRncZa6qgc0DV10he6T8+DCEudM1s
AIZCULKgnHhjUCmBMOMgZdINj4Pt0tLRUqjT7Ak09me2M9ZW4scK5I2oSIkI
WhLCkNdo530XG9vcd5WQ5jSUD4/+Vd1TcPXoCbCFlchoTqE8QyoElDhrBfD1
f5DzQsQAy2iLYy8AZMimp3kD11kUZlYWMZSJNQQQA0bdMZTKWZjn4g03Gc/l
2MYVPsH8kPJKJO3Xo7Gh1nnfeDKI9CApjGU33Mp/gqh4dsbqs3AasIMfJ/oS
uPAznJ8fZ+LPYJ7Kb3aZ4X0utHcSjs12dNN2UVf3ZOhvgp6s2k2V9CEu30TL
c64l+ir5kAu7KvwAzAyHEPyZRnQGAe1N8cC2F8coNltMvFDAe6tbwJGBD7F8
HtqOy8RzzAwjdUvrTETRzfXT742GtUUGdPFYu3hoZAZy3E4OeoQCIVwqpyvY
GGQCFAhdrQHBeaGMRBHYZ/DXWXldqiFdc/gs1g3MRFwOrbZwqZMu0+cyxLCY
Hf+uxMDuKXodX7+sqN+SnQ4FAGtB0Toz5OAbPslUEQs4nNOo8QfhrqsHVyH5
WOOHtyRb6hDFAzCOcum1FjTRVJnyK7rFhZ6whH8SRFPgBXY/0YyUhDaiOWKv
EZeHYXeS9FhPSWxuIY1h2DW5nSS7IlnSS8RXOXAyGFub/FJSsqx+uX0XQ/eV
/AQpQNDBaFNXZpujZp5YjdAYEe99euNt1Y1tA21QLVNt2BzaO6xyf0ZT7vSr
GWk2rkuwZvt4kTTaeBn2gC/XnAVpzZZP8xa8GJCUZvsPR5dyfjnWk7eg9A0j
ssngZV858mHahHUZE+tDEv4XEim9IaPVHPp79LvxDPrS1Jm/+JyXXKz7517h
Rrz/5TN3/onHie7bRoSg+1pRJl+pRSZ+uRZfbXiMVdJQOaMFA/4VTxYdfXhZ
1EmFtBi9AgOic0HrgzMqSoFz/nzSsclu+VR0hS0Lp9AvJqUljxCC6qH8u8lN
4Ro1EUgI8PXegHu3I/ZIvwSWP3zPQwCZ22VOJz1Luqhkcmi4MYNO6ql5Fu6L
bIL0DArcIqJBvjdlhD4QRy+SucBLgA==

`pragma protect end_protected
