// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VMT1E17EJvA3IcuO7DCK98HBtksQQAVUYunD7HXUkciArOZ1md+Sy7yrS396
XxWa/24VV9V3rrodF59u+g1yInJx15xuQUO0KTgIupI6+NlBu3Nx6W0dWHu6
Y/+kTyxa1Xwfn7jBam29JGsZuw4kOUCcX3E9r98D//wAD1QKFtsjCRMxCcNd
xvAV01Y1mkjfSGeWPqgUYbBc54kJamd/QGtA82qiAgZ4mAoNUw6uagWIIKUy
1kuc6JdrRXg+7pw5JlVS7H8GexQoQb3IMq8WTasAEXIvjhY83y8VAnIffbXR
sdg3DsOJ0denB6kqhz4vzHpkBYDoVbDZBspQN0OrwQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h/jSIiIMYk2sFEF5Or/so0q47kHZ3ev9xMYPAu3vb8yuxfHZIjckV4vQ6sjr
5IsxVVWhjl6JPcnLo5raFUHoz7rGjRUeFyJCMtQGHYGCzhWUrjbbXA8Rh37z
kCZb6eTsZGcHJ8Pj/ALlkITymxeSZ7C1KRtH9GwLL2oWtMan3b5mluqtKD6q
HVLBReTh8L/0gHVwO0eJ+58j9E8i+gDwJEaXlFlL3/YkRrkM6WS2vvYv7I0v
40/OppbvYqzmY4bkXCSwbiIUSlipSZO9TuTwVlKkvNyK0Z7jL8jp6mafM7rU
/4wp5jyypFl4YVNtPp6HE2yJF9hTdJv+RsOvVooZcA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n/Idi2a9tA2nqmjLW63JKIzHk93B6xiwy3Y6sihYl/fqXTtwGIC8b13Z+up4
xAzqCYOoBMA4/5eLPbDvSdq4BjSlN6+sTFZ+9M7PnYaAYJtlrbW+5MeOgjaV
G4Rn1U7zxfvg05sTfQPc/r1Y/hrdVnPBPnHG+Of2F0BRjl2GjCxjUny8vja4
CcXFfsoW0e60XG2Us6GhZxV8J20uEjuaLVBgdW87mt99uvIgD6NfN8GpdDnO
UMSBBD/2rNHlrCTwKT3XwiKJN0J8pTWAB31zX+O8qtuwv+/YwMv4he7xATy8
eZXSpXG1iLyO5a7B9+G1XG0lkZGK9hbYiVpZ1n0pqw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hoR2kWVbrTgA8lCkpL2cavgGJGhRvS2ax2CMdCVDkNCIMcu8+DlXCCG8fSXQ
OQ8PWpw+K2JYQ/6M3Fya3Y7vfHJlIwBCv4oMPsX0jKv4qIh+tCvi4Choh6Gb
duzpCcMjxx+vEQZ/rEICJZxmnBbTgHGFVjQJOBnMZ8VoLbNaNdk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mc3hpnAuTDLPGAxkHFhGG8PnBMvH2rRVOpBfcGpcQF9FIiv1Uk4HWSyNNePa
36mP5T7kW27O6/kPtg4Ju8iOxPrANnr4JOc4WuHua3aDQtP8XTQ60CS1QpiF
3EQ7g+qbst2oCaLIpQn3NU3Yb+v5zNuWBLspxDBjkDF2dDk/ChkoTpRFknAX
53Z1aO5V8ZpyA8Wk7XLmGk4VnJCGq30W03j5RstcIgqiNvIak78YDoOepgbz
n2JWw/ECRuXwJtHbh8t6QqoYYssAKWw3dmrG5o8KGvquTxzkkHVwNajNs1Aj
2c7qpsB4KjBMiYJMSLSEqkGrNiQoUNcp2yGFvl2Rb/7YX7pdrFqob/JyZUaq
d2Y/OiGCVHzn98WH8I3aH3QKrE7NVk3/s+893rJyuhark/Celm0a0gyjy1+x
c3qLbjtuGyXBD3KG2xDMkzoML0iQ31cQSm7KOFuFHUZsxi4nwmenDwwBGCcg
UldKFWNEnQHWm/xoQbLBlozevGMMisWJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uTKn27iFXghUAGS34RI27MVDold8JGupl4bMgdyhT6qic02G7CRqX20ihxvZ
SRU5JgNzCnLNo4zl/hT8YsPIBZyGUSr4ieqzTg71Iy6Q38G6g/uKiylSzacQ
DcYZTGZR3EqX7eh3jDJDRijzwr2aoueQGl7vMeb6B+Bid4LFkJg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D9feILx4N8X9e6QkDGYFkg/9hlxCiC2JuTciP4ml/F3fYyIOQCESvTgqm0Gu
2IClqbk9cTpsy8Ue2ZZfpHUon4vwGMG1/Km/VdWgrf0rh0FlkiaMkBFO3dBb
EoVb874Y54pldEq1JwylrJjYxFnag1IPcBz2wzUkB6OYBxJQJvk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21472)
`pragma protect data_block
beORQfYjuqe8OEfZFy4374Fda5kUg4W+OgPcja4y9zd+KkKLejWC6MoXHvET
CJwlPD4UEUw0Zrtrz2I2tU6fa9MaHM+xlJqiAslmqqT7y4lfcmUg2gYOmgzi
kSuvPce2QTUKhGOgneZcfECsZhFW/T27n+NAhdZAb4eAsoIRpzxnClCMOQK/
yqoCT4Uq0pGZUvTMcXFV8i2i4Z9oBDRlKFOZ9yPPbZHb04+wo/7BXI03a9F7
0bqx3YNNQ5CsDfsDG66Kwmrs1t3p2OYK7AfKFLKgaWernOlz/gbln+RktjLe
DX1CVqBvsyeYwqbveJAQYXDpsJ4RqtxuryRnTzKXEo8wQKC+BHAcHLYT+a+k
53f29rviQxNa6rOjzrKsII69GyqDxZZ5TdHv55rRmX5rmO1VQAtvPnwnZYa6
bPyrulY76SI+3+WdRUyDRjRTB3cydDHN3hazII3SOyyS56pDA0tmJyQ8pITL
mNGfxRS6P5Qy/vJfPjQ+woZA6w9px7GLF7ctG2nx+AWwvz35veCNZRksEuwY
QAaYEguRHbCAsIlwdxPcA2abvhIbhCHGrSdr7V0OGwK6fycSzBLLAXDNEQUY
B+T3pgYrzFxfRSnE1vMJ3jW7Lszf1YAoi/2kbHSTWwSc4DJpEbZwBvYgHc+W
QeoN+fuUTmj1OsWWjYnXiP//xZ0tkKrsLy2i6tsrWXq3nHUalrQIJmLbgnZk
YpWK8VoaLszPNNBl8bRK7tA7KiriR9alQE9aLhY7PioPfLna4UFrqn9f7Hut
mdFTFJ0MGTLO6KkAMUPSdpOaqy6dqdYXm8tQnBRYf90eWIJM7m8bDJdKzqsp
fgHHMz30EzHvT3V1pL2Z4LdAtSsA3tmRAX04ZowkdtwPPIAVkuy5ti8/3ciA
n6sUC+9M2Yl1ei1z6ci3851DwbJlfh2PhczVufNXvJbbXeQmoiw8S26mnw7u
rRTcBM92GXtWPe3UhwiuuJ3t7FHcVfEhtVJR/ORZotyzgfjomsxi0poRaKQB
9Wn531VYYhb/9NZH2sO16JY4obH060jNeIR9IYUeoz7Kg/+14G8fV+j/p79c
yPSe+YEj9kbJmtCNP9cNBhEdIe0aI9B2a5hZKXgTQDAq1KeVT6ZX7gqD7zbA
10SXzBCMJ6TzEo8OGB0BLZJ6rl0FPgwYyZAXrFis2kux0TdPBYOlYKVBd6XP
WPhVbz7U/NiYGl0fAALiWVOFycdiQ3rQvqrEsFPfBfBbWCs/KgenlKNEmlRu
CvAvNi0L1gBeZ5Dsc/fqB3rYjg+njzBPX3UIjXZ7CAe84Ux1BoH1tvCS9gwB
Qy798gF1BylZSwk2xpmglPVN9/tI3XK59X/nSP6qzGeFK3YyWz+vslbdegdY
6R5orH0uCRejwbnIbh9brWCOcLMZlOkMyeU6UL1xa3hy/kKa+G3q7OaZ9nX/
Eo390i+m8iodgFFp8CoMf2YzZltG51696h0iQXvRsFLLIx3CrzPocw2Wk7oE
7dZ5AXE1mRaKSZs9zlL3Hjv/kN5dg+VWluSEXPF9YjjdwZte/+DolEysCYwp
MLNCq1t1JgSR45lumrikONXxjKAnNbhHQ3dgEHv2yupyXyH1l+VCsYj9zBgI
k5O+KHni9PHJURCmAmZEM7VbNxnlWIZHcYiYpBHqRsRcKmGE98s+fcYpW7pu
nd3Ii/1YsJk0refGnqQqWbNJ5S+LVFFlgG60NxvjYaxcg5YoXrys1nzsDJwV
kyyZ7rS/HKpZ+tivZ703GSYbBwS4/iTwnL107piaX21bZzwSk08HtfHQfvIl
+OkoEL6sHJteCcqAZ9n/1iPW7wxv/RYyQ6MNauDmfVZku2iJsWLMKZDPhhZ/
2Ubt/AQiOE2By2/Rb6eXfD7XdwKtiRKSCqIYb2ePyCPnReQRMk9zEOopOmqX
fzymgWrVPRYt/El19XBs5R5h7l1pKrYFMfGb4HaL6lmND/APt4rkjWoMZAwt
rT6QpzZDudGzOb9xD2oP+c0DxqxlQjaTI+WhJVvqpUXmgJg8m5LVomULrx9M
53jKBmlBYm8aitqT6Y5NfXDSX3ddflAEhPxB9N8ZkUVh3xg++TmTH7jf/8YX
2G627s8gFqer3Y2VSXEs3ZRL0/NCuDqER5okV3qwu21omdDdT4F+pJWzkxlB
Dy2Ypmj9EPbJuMFCt7Raun1O1lHx9oAMPpQp1uhZNx8Gl6PHAjH98gxGYT84
Ga0jW1zvr1Wrng8jb8JJfv2ynTU3o6yekR/+4ZxqdUj69WIs+JCgTpyzxB59
ZnmuK/ZCL7ZcM0U7xk+3Hf1ojvSSpJKAATYNshlAYCRxSy0l7OB/nOQy0RTn
nmti+4RLZf8e4RLPp4qVS9QQDcN+cdEJnh7d6h+dneTBxo0jC8D/+cL7rI9/
uWzJaLTzDkztn+cveZgWEQer9UcgDG2KIq+f+QxcGmXjYuY3phM6YxwEYxQC
bDg3GZ1F5RBKnkggEW5M/H3D2VoyyAkfTd4/Sd9V3aKDby89uHwi4W0VgRk4
tvN+V2VqckH0RwZO+8p3T41i8I7nkbUbbeedtq6gow2r7yj0Di4OF13HTOkx
BuRCJkulP5EYbxGbGrOJRXLPJbSdM9kKgim4lN2tZsuxzji2GIQXHhkbwjgL
3lhGY7HTlUb4TvagQtZo08FPArNx++2l+rSwiMAvKTf2ZLROZ2UXRlCooIxu
qikViUJDE/k96/TmKqD+sTCZvMlhPs4JfxtloZAKgXweUATDlW6GWO1qMK6H
Nn+N/D0D+VRIUO+0Xvj4Fgl9DtS86qO1fTSugtq1nJ1N9r+U0KeZVmS6Mhi7
TiASeqDcQzDFMQZUn9xlnBp0IIITjv9ETy3g9/p5E6PnQuh9mZvSuL2HoYgD
hG42jGklxWR7KFfFrnHZHN/Il1Sd48hkL6oDSnCUNPxyFgG+y3svhqllUIWA
Q+ifuabO47BXVAB/1oz7uGSYDX8c6CyQAnAKXTw6RrJa2K6pfkzBeDg5eVpD
Ymhb0FiXcsZ+gxX++o8l0xfqtuYcKe1EK91lz4wIpoPLzfpgLhML+AqXWYaH
E5ou8eQcqIFag+TDTlj6/BsYTE58Dw278oodlqk9t45eSDRYxHOUBrjQkCDH
BXxka176lF0yhJxmRs34j/qLX10E2fPn8meahGyxcx3LxIlkR+k6yDbSzxH5
n9Llk6nwk5Vo1tOwFHvV91SlfYLszJHc6j5FhDn/Nj6HZpVEEqEanXRpgHHA
cASvSolrL6HtKOIdfQuBAL6akQEAeAa/Zd7CuyvNG7u89eY6r7l6nBliHqaN
S6OQeMtCxfXUmrziyzVKVRZmtY5OqwB56bZYvQc8rNwv9edPHA4Kfea+aXOL
Nloowkf4sKYmN0uPPvw+mFkN4oCgTF+xE5k1nHUsNrkUavgWHumCIvOeV+mS
xwPCsY/fvipgPUPvd/e/kJ+UtUPo9LgwgGl6A2cRIixixOzff/Nd3d5ul8ge
6STrqOvIh2/H/sxU4X8+xFjHkaR48PWYdFIU/5p48MUbMu/Rl7CFErc2o0Dn
CLnx2hHg81fKrtVE1TlutdGWuRV24CBKq6/s07XxH9GGnjNBvI7bY2YBR5BZ
nMjtuz65x9B8QBcjjlIwM+pfu4rfmA0R4UH4WAiHOxVNM+YVADBdeA1+ajXN
/mUjLbcVw6s9o1BYTAI9f2NVXnTJjdkgs/QMMhKUbAjxtvWe8S7ddqSW7X+q
n87JEemJBtNRbwMf/34LoSyn8pT0MzMx76fv0g3nM6yEme6BKhzoIWeGA0Nq
cEHSRpaWA0q0tegE8V+1symQNeD4RGdk3g2EdbkNdDcmWSPnV5TL72yT9sKA
c4Cj8OQn/z+UdfRt70t2bK0ge4NmuCBPBuYHqXWni2Ih3atIhQgG8J1iy/jy
fwohRZxU9KTV758jFZZf+rAQ/pdHbd55qWDVWuwzfTIAARpRQitIWw/1ErlH
nGghYcuz16Q9iaff9SmgxcfkbQndVr+HjHVVYbJ1P+AyaE45fgeDnGWf4xtB
A0BOv8Wfhi4hOVz91Jfjo3HzO4TKLGNWPzAHZTTSekZDTNb6DUVN4G4vCByZ
Uy5h6pV9utpuDuQgpcedQV5rcwbGfEyni9RrwUeGHBkhI7npS9uXRnpF3lUn
TqbGcKGIYIin7s9ubgSB1M+MgS2wjkSVka5qd6aFLhbnmooSNqJiWElpSI/G
b5mvv28yTrnmzv9MgdmHe8QXwELfBH2fYmERA5gmqCaz2k2xg/ixI7n6q8Mq
MmDstooKiovQqqSRG4UZoOY+9NlTx855vUUWEvnUS0JAPorxr5luO9aBUt0S
Qxt+Q8mLYYoGP4lrbMBNKHVoLxaO8W5UmJdmXjagmEoKRYQ+v5vbgCDZBSSt
OEWeBr1rzVdb74k2tXZVXy5mx8Kx7JzisENHdhUhUHRIkDSM4Jk38vZUkjU/
bTgiMrfBXRKfH7mKStxJDm/Vu/NR3MuQxGlcogdhvX/JMj53hqIHCtTsijUu
AfnOLGpez3iTxRwzGUBwAOvdkWVyPtiHqIv6oC6OhnC8PzQxh7nVzFa8LN7c
o7/c+5mx2HdU2gSyvS0DLpf5zal5u8cJoXZo/E03bwCLaevayLPyWh2iw2hQ
xa4/Q7t4f8L8VXBy3qyXAJSblyCsLZIikwZt4cgVtAMh3jawZW3CkKkDzJZs
fl40Na4jascfLlN8yFGsjWsvyNR5ai0nXHtetMqnRF6+ksW66QUVnGh6YZAx
JdBN70K4PAKZqiMLF9oe+BOBu0cAJcSPoluVoN+3GOLxjAsBO+au8i8IJUAv
9yZyDvFNdaKMoJIGB/Baq483aq+U6d1TGxNJiNEyqTnlh8DATtvWpd7bq0aV
BidNp7IfiXlejzq7LvtZkG++Ucq+VhH3aZOzyY9d7Ub9EX2qJ7ZONbzNheY8
e19orFHkd559FOZUKCEYi7+jPJ9aFPqOKQzKbTx+34R0funGgqJVs46EpYUD
xf8aNh+iIUR0t6wxYT+zdriihclwCtLvY8qwKLwx+Ova3Z+oeL4O4G15h7q/
RFAwxflS4KPWvtZMk0VcPENzN8L+wxDQJOB4zFeJf9QTimA/SGMPSVwGGyF7
T0Obagbrd7iniLTQ1oyh/nW6JP1sMIwG4FK7yErG0nkq/efnyUhLIz/z21BZ
x/SWdmjo5KDt3J8SdcEQFEYQjaxPLWz0u/c6wRWOXacH3nIfMQV+kpF+iLJM
0XEeH/bUA+X/2ePXropuXtuhJi4taWOfWFE1EC/3ONmSMO/WlYHZHeEW1Fu9
p5gjksT6hZ1vHJk3ku6TZ2ZoHyaEYzRMrjTyEmV/UajET9hFbpACzU7oM13S
Xmgla3tofVP5XaASAyBVuspH9VNpwnkvUwM1hYNyeLa8DgCBBBtWgtOAg6tp
RJgNH7A/Fkmm4mMCITieti/NfRVkQ6bfyu5qpTAutqPJdFm1V5QGcEH63pp+
8k0j0w5EaqcQJleiswyfRyzVPM04xYKBd/y29KdbLPJe2BeJoKclpa488rIm
n/0XIi/AKrsszTPAaovUC9eqcKwGFIAUmRh83dIAYKOAr/0NRNCXlj7BlkIN
YCQ50QBe1n2KjG6Wv1ATKqVYyXd8nJCz94XEUL8MPGc1feedNBE2hV3py9T+
2cQYWeurB3cFNVjU5QKY6jhkmoQL09frBcaFODWkbWhaAiXwQ5nFhKEm0xMr
rBRR91pi2Px4ceOhDvrxdMyZhBLnwm8yD8zXLRybZVsY1LDEeMZWffFZQEhq
bkI87We6D3uGrMrQVWSL3ag38cXWU6hetWmv7xSODSirY54jHZmstMFP7fOB
3XycReUHZPxUA512Fg0Lxppiky6xvYF3JAgsDGJShT/QvMfoMQTXd0ky05lX
4USBlbuUH61j26pKMyz3nrkNEEVA8YpNswf9Y68TUXyjhartZissm3eNi/a5
cX1jcEnEnatYMM+DkQdS+tL0gDSuBAe7nAc80Yp9t17romeSQiRu9uvHT6Tm
G3QvI3cBZOpjLTSW+l4c1IlXBc5e5YGAI0RYY6i/cSXHgc/T+nfb6DCfHZoc
AhDRmvRFT+KDr/Kj/0RGgfNF0WDhJEvOJrkPkMHJfshdOM72THa/Nu5SRoSE
vru6+IaaKbLqLfbt6xC+zec2el+/+2w0+5ur09GmLRdtTbmFkf6tZX9exs8c
1KZej4J4smNO1H1hTnlmQQCKnlf27qzm+kdYLMsq+zbkcVVz71HI5W6RbkbN
wwMF0N3n4+QSM+cxxahO79NCnFZImgXSL/i9qo2p01MPkiCFb5Mx46y+gSrX
ZmNx32BmphtVnsEq4gGjykMpxj8mBoB2dqksC10v5lrA00z0gtQscL+s1gXJ
HCSCHDIkusTm7cftOhBoi0g/Q5+ds8oqiCyocNy6Ekf5nPOtJcNEnRoa80mb
xBvHF453mKsM5U5JF++RDGPmSwY+cGYLvc247h0IwyrLNZ6LhAqOjiCx4Uj/
iZaicnGGWvFdOMZJQDVr0pFDCrHoxIetONX/FjNoZh7I0//2m0DyEOvZw5OF
zUfOj2TiZH9PV5DwavlEazUdCFvdmP1/VJeg0gtmoYh/cXRMFdSE0oK0l9C1
MYd0HAupBQBaC6C3sdwF86qmQdES4R+yk3zHxKpck4v1xzN+zMSxyasb1mjC
zUXuy9nuxiW4W1JQpVyQ8haALqJn7K7kN0uRs2IobESKJz7Qa74Tsblr++6I
4xY77InesRKRTWbcj1XmIqXPXjazYGqHNwn/BH6zBm2fDOP5Oj3/Zl/V11wF
iPS7WvklsqZI7MP4wq3JtYzzphh3gW0KxpwA6HYsburygZ7TugfrnqbPC1PH
6+fBuWz7SCC0WBESgd8fi4Fu/Frn1WrbhLl3lQ/SuCdO+Q55bTic4SsWBzLT
yQiDdhNAuZ9/07w8RvPR5hZbhRXRPDH+leFRPxdYkgK7MYcwjkRW8nfSfkn5
PKOctLMjgwVJmVQffW47v7AxQvtwpZUkRA/hwMTayi7dy39Sl5C10aGmdHtX
n6IYofrJGun0oS8HvVP578ur90Zd8/5LFEy2R24BZ8LkX8YkgvjKDGvzmX2G
BgZVND9AOZifFm3qqlmh0tqfvg1YySosM1V143iLHzXtVff3vr0t/SgIvhHM
rCHF70Z4T+J1tJJywkDYs6HHtOjTw9Ot4qloI303GuwvrJGhLyrGfvL/t+he
RsS4vQZ+JBjAd6T20eqLCTQqdnr2im4a0uXlfD/df1HrueAiahMyr7mSdAUd
rYUfzghqdFuIdvcU3eqoe1ZWzjaJmDriH16o0FrCG8O21F4Lnw/AyXfxKpcL
7ubESAOGGs/NZzmzBXlBqSvxmcv1eeyo6ffYv3f56PUxFAieMXEMNiNeBDbR
/mIK9DwOwW+2+7s9UxtslzkC4Euj7aLiYYNpdLDX7mmPpCcncaIsyBjoDvQi
XErctQQdnjw75AeQ+hiGappIVdrMOAfcojBB7GAMcXSCr3ytRD+D6J7StvcU
18YhIzPzkovGbcy2ztgpals+i2GlGzaDIp1K+WQih5uPUZut5U/shZcZBp4F
ra3vwlEQhZbkEnc0H3uA33Td4+xGgS0vUvwLOpapdmLU7HbHSVIJlWJ7Al1V
8Ejl++TR3q3DLGdndsaMOEHjOe7YN37y7YwT2igyyvFXSQf137ZywshPFezb
taDoLg4veTCPMaz9wlNqauYfKAV/GZ8KCK48PH51lobt3GNcH7mkx146q7pX
YysFLk+GcP3rYZ2za6tgrjsSmOzIC7D2NYb+QChVZKanHS5W8ex7FfZL2m8k
Fn+QPJXx3SlqRACErvVAUJ2K6K/kQ0JZM/q4ohFOQx5jAlkdwfemUWoamt7K
5wkiRV+Vbb3JdK3SWrAIgA9FaMzgVWUiEZBBEhM+sQSdYFUXHIHFyPTjhIJ3
B1nR9Vtrmz5DRmYUWMCPQuZYHlInXOOHBwsVn5rPzwWpt4ypkF0PBa3knAxc
ppE+1UI5qkMgCiFkk9KD05/eMS0USxGV5feozmAARrK2HNGIFoounPZudYEH
NLXOQ7YXNBzM63xNceoWp3s3ZXqJZX+6lgaEqjvRHa2S1QKEVhnGiGTvgTOb
UsmaxfEtknST3uiXd3gWoIBvugDMotdQqx0du6fZJTa2ldyJyBvX1AX5CfmM
9ZBjlXgDRO82qhgmK8qbyWcatzt4+KbhrfvB7JVOV+BvvBbckfmMU61dG3lQ
FDOpGl2Oh7PnS2TsGu1awoknDWJANF64EcoCwaaPA4rlMopK3CaXOV2mQh3/
pqQf+GgnrJkFC8vWzKgrm1r/o3Conw/BCr9tD1WNyzYEQT2Bnq0KjPtPXTBj
gbc9F60b04yVRSKASDFy+uF8Z/Nkffsdogiyg4x3dRuGAp/yJOkvG+ow/Hrq
6Ycy3XvS7k1xQ6E22I0uzPy+Rfqt8OKU/4P2oFumDSSM4ppTc1qnN6LPWYKV
F5GwFLWu36br2EVzfkYq7RwOKHsRTVuqCCOKGUxqzYLWJkC3ojPtLC3GcFxt
unNO6yZkvS9NWUqjDl9iteV1J/Lmqe3YKF7HsPTygx0ArIU69IVSrbh/ML2B
X8CjPWf3eSz929cInnPkMmArrBuXxc+8uz7GphvuSmNXgj1+hdLmnQKaXmhD
dp9s6n2Z/gUQgDRhMpQrz8vJOlmiTrngJ8agTsuaD4n05mU9cBCRwda624IM
BmIAmuql43eBhGEXhP9bEAqWTSpyv+oVI4800noTyzhR8/MEX5ap9IObc4L5
7fWVCrEiAUerp1+Q+Kv6kClFZiYmC1ivmMn4eA6gP8ae171OeLn0hjWX45P0
vndroJVvPqGo/9ygGpCXFL6Dpiz1CMu+FzDO/zp0l8L9DY8V+CNEdVdDU1r7
0C22C9HhQ8GkqoVztQQjAdijBtHlCRumCaTmJr3SNw8IALqx4d4qZra9P9eb
FnAeP74za297UMmqri1W/pV0X+5ZHDKcXUvWxpHLX5FA81ChQYDWhOEa4Mvr
s498miSqUUjLpLE250OevWE96slVheNrWqi+99g7m9bhVD+pX0I/eAg5WkJc
cvOkzL1H1z6KoO1zdkPDVjTF8v/RX153g4fsQBSGr6WBNvSDWJLreyp701lL
gN7/gCntcs7WW0+de/DH9JOvPt2Qkhp0PU4JPphmReuPqYj8CLTqH8ff/3p3
ZIZz6bMMysOdcD/mxm8lv9p/xmniW9q7mmc9T+AANNVH3FpA1qVuAAy+PAXd
NLrYrnHeGu2dd12mdyiPQn+AKmvajnGvgNlXqDv8pf+HPv1iMyj4ZwL+0xvp
BguPypQ0SqUuOSrnS7abApNOv6BKGwGtvwoReolJjqluzHQFUfydPQx7r03b
agg9XKez4yeaBjEnuAfproK8IZAywiFkJD+pXQ/E5a22U11IVyYthV0rSWFv
pVUKRH+lZOG78Tmox+pNTOOwKCoIFbG6n6/iH7P1KI5Nsp9TZAJrh/1AQLYH
jBkAAVaB76VGy9JdsC6YhY4izv898ELRgEmoY/Lo0dPcoW2kYpuFy/EQVEGk
LmpkJkdxrgsbcyUZV9Y7DINdqM1lKVWgvk0P/HKT7QzS/+1SlEReR3t3ryL+
14OsyfvunW6DTlKc7RotrW3M7Fj2KJxTbvJMa2B76XTuaCsT1o65pQfqmfLi
/z6MVe7jcA0F22cRnWiiI39JaZ/xqE1mS8r5gWuOuWRsJh912qR/Z0InjIPY
MtLYYB1KpSWCfpxVFXXErjaVMU/v2Qb6p+5Qs2e2Anu4VI68R3y3fBULi3CG
p45nGUZQsb2mVVBeOxcT+eiAQGIzFwTWRsdesEPkHAEnMeI8ik4OESlq7ssQ
9nhQJcQArzCu9xkjRLXR1OPP/PooNID/+75RB8rMvUYiT+DWzqo+5e027ZTV
IuDOoadfAsw3Y0Sphw12qAtJxm3JlRjjr8VLAreg9+gMzZE3kHE8tItcFoen
7YrT1Aj+vHEuV1L/5OaRpnK6pwevALBZM7zJw2vjzEhc2OnCvxAiNzDEJRbV
l22K1xXEqM3juao9Tt1eFSHDWCkSG8gp4LM84hqwvDSlvS18vGAeRmJ6hbPY
ReTx+VtPGWnigi0f8sjGgQtuEsJFZtTJDvhoyLAtLJLTurYjx9/Gpvece2PW
fGemA8o9VOQDXiudb5wy2AYVrrD+cq+4HdlSh5mbcCCBKy6Mh/LUCIddj87F
3QPC1F+dpU/cadZEhzfgioGx3zdLoZ7S28kM63P9a6EBK6bRBlGANvsXn+oJ
GoHKn1pFnjXxlR4vUu+lheFkueqvdG4eqQ8LnzgzsZxlIwiPuRr86ZASJur4
lb31xnKOamQVHQNuEid+79qYfr7qdK082KVycxu3uRUth25VH2dmx8F4gAEb
MpB7QWNgocwlgzByg3MHH29Xw/kDZe8AED74h56djspJGL/avwtX5Dveru5K
4z/C13RRV7jy02FDZYZp20ofEWrK9LKt0fEsooa1JumejA48VnvM5tCAA5s9
u9kp1mfmFC3m31W12T2JjSvKzKvPnuME0xjzVFYyR5V1SCwGGS2PvFy7vDsK
yT/eWM8nvsRmdZ91ISoAYyZMvPgVi6EliVSgqS/r9hlclfz1079wQxk1WqYu
dx0QsvnRee4TlRmdNj9SyNxP3w0zKlxiiLVsOHRsbbwrdmvyjf/U+CrpKmpG
EYORV5KkSj0chHBE7MQ9d3R3GRGAPZa813ZwhhkSFNUL9136lesUDyRyKbP2
+K6qMvqB6a0YBW8JH4EHq2hYi7H1JubjoZrQJpJgJ9V+qZyESp6nYBXutoSW
utw1tESaVbutFl4JopccjkAf1PGX4WzXOeALvoFO0JxvnaRN9fgWHxU1SfWD
1Ap5w8eNQ8KBHnb/IP6k7CV/bLZyLSyPvirA3iuTnQHaGm71Kv97rWKPcfRO
ejc0fh88NxhQCO1tqEANKGj32RzulG0PNgHUAUcg+/2eY4pkj/cplIj3GAUM
VY7p4dk3GS3c8wlJouhiK4LnGtxJEUyaOLhNgjas4pzzHx6/g4Rg7tcd+KYS
FBGeOGDDp1TETGVeycCJf0YhL5SlZR3Ey+8NQPrbg9C6hcXAhZKqt1WJSwTB
S6UFFUhE9CBpcsMStg2C6FNhKFvf7ZqDZgO8mo3rs0tGgtO8y9RNGPr9YGlW
8v5EL5M6RsILRHD+Acl6KMAkr+QFHX7EuHBWLBS6B5l7b8iH1nMawvPtZO0s
lnr+xPZw+uroOnGd/tMwtmGPg6T60+bXFJwaHhPww3SdOdon5VC09++IhUl4
RSTcxIzH6DXAp/Az+MNbeHKVeB990BVt+6O343rG+F/w74ryNKbD6677dJ4K
6bXZDpN857+HkbYwXVik6hvIdsP0eFbdyNtKCoFKxt+Apyspin0EoymPILJw
uW3//YFTwxjYhfqeFAp0NphcVC6Qvm0wXANUEc7E9hJgRKD7d73J3oegNz02
EzZCN8X9k5GvJpzm9wpbZJywNgKQPH/g04d7/C/0J1tVTCZqy8H2KWWnUaPf
vRBXSddYeKBXN8s0VOBsTWuOetd+LZqjnsZdgfZD2PPOErj1bVLZHyfO/KcE
tCI2UoGyHgF2cs/cFKOK9Yl4UhMCaOPYVySCoq5N2Uer3zgmhM8GEJpRzCBO
bsiieQF2T7j9Eb6J3fb27Gf0ehnzSz4XMZErwLkuobgwKqVktQeo1fJpsosi
EJt8hW1b0f36581KEWEHARWFBtKq4LcJRz1Y35GRW8mzgWLtXzDHeVPe7kR8
9CA0UYpRn5UxTD7Ys+szMSS3pLkDs1fvW2GAqGIoWvhgqerPlT2mkxJMt3Lb
PHqIdDbxf0H/cqnV+njWzvNK3m4zDx04E/FoS87BsJwCwoGWksyDfa4pYScb
rxaXytMUbzjedqkpIAZHklQUihFK0i5R4Asr6gOtNKEQoQt/cpTmQ1Nfj0/r
6fOGNj9KVzOs+pgJ1INCmXnaygSbybq4sQIuISsOxTtIXk9BnqY4By8hGqfv
gfRC08tKI1fA8dBNNN+uIxG6mjAuPet3u5ez9Gx/ad1dvw7+NdYl49BTbKtJ
+tsZBIAFpqvxduAOsB8z51+cGQIyIcek7jRa0P026g6OUVE7YYlyvxH9ZwFC
VFVh1btqO21TUmMMzNy+mSVCmVZZiRBd9z4J9yoFpDp55tVZCo9gSFr1XSmQ
G/l+JBQ4SWQruTdDXsOagerzaHs5u1QU/iEAooZbaQlXJrfxl8vaPNM61k8h
mlvKo5hhgiwrxAK4tp06ETEHli7ZUwvFuabpaAVcmIQYjmTBL3kbc6bt5uTo
OC0Sd3sXl6deswC0CP0hNkoALU6LaTNwXASAPv/Y/yykHl7dbdxRDIu/xmZc
wVEZuL06iWTMYFOX92S9CdMu/fT1D7czhtsXooYRFzLrgZ9QQUHHa/XWwYCo
NN/2fQOcVjBDpE3LZD5ccYvXU/CI0TjNWW34JLPKq0AvGDO62H+GvbwygO/8
HjCSeNh5BdaGd39695OM7I5YSD5J7GIEZEq6oEg5uSRKswlYQgE3uHKMK6uL
5xP1dJ0Fu9Ffr4yPnnweJqjsdzxv8uHeG1HJiHQYbxBZ7xt0jhhGTPR8KUkd
ckuY7L628H8MbFaNvuDEWO/E4xHZ3dpzz77MzQ0Ajgj1zXnrLRWRfUpcRy9B
0qSKwvNcfro2RKtSP378ULvE6ERhYPb4mCDF/zgsQDdh4UDIsN3t6qAlp3oK
QhDnTlqcrbbQ7rMymH779RDa+FJgTzOszKFuXZKKTznOqGA3crALAhQXzb1Y
S2Ekz2v5nZ/eEg8eOlJrDraLbYHsaN1guRULp4L6KEPgW7RfnMN/CrFnjY/5
n01dKVwsTi0bdWzKOJB7ltEHrtlcxEBDEorX7eL4cJBu1SrTaOnqp/2BPOLN
NGeSjaZYC7l0W7OoAXna9Be4uDlgbvz0zD787+8GUlT0p/JxX9geXypmWCrj
uof/rTHbXzeWAIbfmZV+Hj7QCrknFOOHWJWJUmooAP419HCWoGRUGgoQsVMW
0mY9EQu4+1OnsePTvKkp8eFQuLxxIefs4e1zM4dY3hLWP2MrCYIY6xCmt/jS
umuOB2UJYhvWwB0feOxV5bNsOpT/OpQw91tDRyIKlJO0oq5m6XvLvn+rUyfq
4OG0mWt14oBAFok8vf2PeJOR28JBucdwChj/XenIR7wIdOEQYmvj2EZAFO9/
a+tpDIFh0Ig+i5s9Kzp3f6D7tL0DgfD7/Rp1EnniAeH8IGxiws76e8zts121
Jg0lr5+1I2jZWkPmuIsfNAym45t/q0rmRXdR9dfYZcgi3or4DmeToPyQ/J6B
AN37BNuFInw2DIxfBJF4TPbP+jugwX3jnbPS1qS6CfzpW+/LyDjUvG4t/geI
IjOk14Js6gy6aB7lzf3fwTePO3fA1CwqADJSHAj/tvYPZkBMheJz4MIf4HkI
MfXF45nORSaof3pQaIv4NSKVcFVT7i4LNTv4HEvZCcX0ERRM3Cvan8lPDN/u
FFr8KXIBr0lKr6cfA8tm/rDZE7t/2riMZFgpsL4JGM1hnd5pv3TW0PZpf6aV
8vhwjvMHZWmWgrnHhZcmk2G2IQ9Hm2saEPMIuMpKBKu6d8ZqkcPArNNbgyS6
ID4lz1zvmSxtfkKjVte80Xcp2jCUzTbHwkTIv8nZTgxSngTj8tFLAAp+Qiuy
fNQmgZ9Q5MjXVGYtcjFHOIEr32lOf/rsYY5Kk1l2X+fHwhqK0r5QpnSmebxf
mNb1u5o2B+tckA0+0J1D+T9i/UYfqXd75L8p97cuuzFecmOqgf5WPDqlynIv
Q8nBXdFFDpPk4DZq81XMHHZPI7d1C5QC8Kj+GsAHbTEBTkDrvy+0aUAuHtPW
3zQnAu6arCNFBYw5bSpVHes7Iuqba/uY3zDaxsO9a5Cj2Mr2FgYzYO2J0ZUU
ZAls+s6w1HLLfcPS38bV+3tbWKt3so6e/W83oSGUvfZDEklkSrH1th/VMyOa
CwnvpRH1RFqkwtdbpNwvVgufwtnzDscxbgziIUajJ+u+ujdqxKl7C8HIZ5kD
uJcLoy8OuRCAK+4qlaW/AMM4U0IFsynY4cbBqA86hBH0sTJ524APFu0uE4GT
LTuCvZY2lQGgzGfi5bBKhz80AHZhIFSJETUe+mtS4WOe0i/gdO/2cG7vwmzU
+K1kpaAPmAaMuawN+ROHoSfLonJHjADC1trZA5B7HgKyG84RyJc4fxysNDS8
RT0UzQBBxx3g20DLkDMIki1k2XxX04tPONrdBPjegATxWeyvZjfEJMMJlKgO
iwRiIjvQmwHLndnETS8JKDrFdmib111SuoZViL3WMIas8mbTQ7zH1OguU100
J1iuKqP5q/KNci7b6w5O2C6zHEGcjdMQiqhG6p+xv8uvexdXQvk8fhlLtt8G
B7k3kZfu4JaXdVNYXqTdWbKwIy18gmbNCr8LUf4D72Tf2xDsBheDgi23P+Vc
Ui4/PKD4gXHMIy0lC0nStIM1TmdL0so+nvZkJjODvqw524uvuhwJAXo68SgU
QLiqVHu1sT93fHmzmgGPNcfmIWH6AFz1hGJmP0aBVP2SyrkPUBILF+NaNLUa
Jtr1V5YkVqPcCHYqBJC5MNZgR5y0nXW21B3SR60RnQshe+gZGkD3Y5IDVFQ2
yPd9m7dgxoeAQap8rgp+EBNtv1s6mtuVvPuSqx/8HbOc6orfKRYuNnUhxHNU
4jP3T3Wmizlx0IsCLd9ejW4JDaazLIwm2m3I83eLDFGj/VpoF7dMWRzXiN8F
Sw5je3GokCXtDsN3y76Zh0rbBT34MKxZmKhjVXO7CJC7UZPojNYSLaDGfAHV
bPyXfPsyjXzhuvZCzheo2wdVKy3ZOki9Nhb2SHRhOf/LMCN47VBOafJl7Tx7
+JWto01qmE6EoSkjmZWoZqO/HUnRc59a1xQxzk+Af/AAjrOZZ8KC/jGFXJEb
Es481jjNZ3GOHRvN5jztGiRHhc3LtXDFODfUG1pxS9j2epAttqQoAuZNXI+m
XWlAopOxDxtkioLLMJB6Zhe4eH8p5XGOXMgVkjC6CY2+unk0ZtmTtMTcBmnZ
2o/f4L5rK069HMyVerDN0Ei5WnCLIO7dP+z/8SIMFD963rUq2Iww0Bv21iWa
AFbbXeeWc7N8KOmRkaqqF+aKxl15M7iBSx3z+OfjpFJ0pu+DXlSz6xLeQ1PU
Fs8J4NtAjamO5/xQQciDT8EeseYqESyhYpIq0ni3M/XW2iMdRC2HkhAj2flk
z1wH98a22fyRN5GRVeQOFC+XZxEF1aEH8+yoNgWsjcaR77WS/Qx8VuCh0GnV
Bn4J+8F6yPHgMnDlL06qFcXD9fGkis7Uzq2/fyaqawIxbI9z1YuprSeVt319
VwsM5uhPGFP/jC26BgcyLflc6kgevSDQORk41mvqxD3kHAHq8jbTFTstVMoP
gntEwsIMgxgM5OJRctDemNp69QakjOEgynOBhCshNUHNeFN0K7rZ6hJaCPsA
oGGzld7M17VTEveQSMBAvuTsAu1q7GeEvDVnt6qq87lMzDZzqWsGGHg3+RxA
TvLnJ6TB835qPJSDAc2GOW/f/RxiGTfgYFBwGkAXT7w0w9gNXlGU5jF5M8Ro
bfQGr3EJJGcZ5oua4bqY7C9vXsb04/mZXmvB0c6TPsqtNVP7hDnLQLZh21r3
N1xpiLxWt7JSkIBS9EP4NIbi3bdyu7TdLMV3LK/qe5MWf1qYfYtzqHhey2Ue
+Ly5qkylpmAZqy0tNlV25FObKiuBvBlbOsBxv8BH9HC25vjKkf48HDAPwIMa
mUhga6vu4QOIMoz8O8c+y/K+x0IDCpQc706wRvOU+9dX02gohi4sBWmLoPKg
quAPPGiq1K/J4Mqp2LYGrZbP50/adQH/KcEg67zFBdbAyqcUh0CsWVqZTEC8
bdn+varp/J7Oc/PeguiU/OeH/39v5fzXIeJPBjXxrcyWbIMK7CFHB91zwsuw
Gdn8s5O1UuXbk6RRcxoPLsZsOXCrGssQS6NSQU8N2WQ8DL7z+Ckqa2OE3hyy
QU4nwuv1tUtoCLG7ZHPmxxIOfFqIUVj/zGbbnboRGa0NAAYbZ179XV5FA+wO
OQrWjJwHORUa0UFQSr7ngFnpnKh9S6WlydXznmpxKn8a/SPyTspvrF49/HBU
hXPeK9D/jvxnPLp7MzNIUz4XSvWcH5ZMEd40w2+Qksqbjn45osVF2fMGOcHp
NJreHagmJXlSfxaKWkGrVGaQv+kEDFzB4QZv85jj3PJIV336XUq+vudw/HW7
CukPiroy9ZOtgOHRde7BM87rPOSdDBQoupUcAxU5OW5SUn4lbli9SoRAAoVp
uUcrcpz5IJJxyvu8UHu3kCJSq0atuPccDVl9+O8j74Fqsg1wcvfUHg4soZcF
VSwWTF30gG6tbEuZNQ8s2xkbaBxP0f9IJWwWNOSa+9BlmbbzZQG46IB6TbrI
XaVtNZwRGKOE0iJVQ72bE7WUwdrp3ulVO7ytLYx2iqDRMlT4CC3cp2TFUVQT
Cm8gGmCMvCfMqY2bb8B2TCESSorAiEOzy8FGx9VNy4KmCbzyrsbzwaB5xcVA
3TjT3EWzSLspTJ/CKw498KR4J1fXmMN39xn9JGw5MDwhfuxdAJVBjR0Vjddi
tmEl0IRaWMMad5u62YwhKKDmQpH58P7IPutl4pedPBEME3IN0vn7upseTza5
XfPCOnLJsKCMYt/MG385VsFP+9I83jpfDWqdYEBC5cJxTeX69rVgjHRruS5q
BqmvHYQ6IpplngtWrZ+5JZngDyGQzpErUKdBvA6LrTcLxhSrefBPb0Gkvj/7
6K61RYiaA07dlGKr7ALYYK4xa7+4KnkFzcHNNHJdzPEPJdwMf5o97giYVt6z
418nOSooj66HadxobXiX1l9UHWAoyYYfrVW6WycJeGf61AO3yBqkhJ95FaQp
FiPJ1lXkgMgVZX/FGF2tUnc3lZA5aaEjtg2GenuWDUI1nPzTYWCIiLR7wvC1
QFhNKwmx0hF027jpX2J37e3OBVXlt8jmdwXFcIzMw0Lv8x/J2aju5314MtWn
goq+uwu0cKmLb+rgyM38XEJSMr+E62UHE+ea+dBGZfpQhQEL8cZYkodKKvDq
HiQQukdiVUpLB3Ou7Y6TcxqNf7tyWZj9dviLDxanpAjkeUdTSKFOx0Dql/vh
EICQsl2u9FH7Ueyu0QiVNEHqShsVTaOAcoUtrc1+LILQ8gWPZbNKmOnPYu2O
7GdxxbXqidGTWGQDXqyBoNnymlOhtw/SWqH6AA0B293ZN9dHKxlMXlsxnmy2
WRrCszmedJWcsaDMydyiDNHr+Zfst8uMFm8nHS3GbSLICFpL3RqxeVUHDusp
MMZGe1ypwrpCjW8Y/PMTSkQyCEx45Px946OkZq0Txfd4H7CkUQoD+oYsuzhZ
PbqfxtMPsg1XQucvX9xWlkaHN2SbtFDOLUc/uyf25kOSi2Ol3XuozbOQ46xD
2GJ4OnQYmELSl8MXhHkIAfURjlGhuxXaZg1ZPYHqTpEnRNRwD9X1gdsVKY6Q
KoG9UgSvifapQ3YEdrIRS1+HoSJKLRCJ35d4lMr05O751iin9Lrgt70Pr1jp
7pe816p28INYJEHh1zwnICgxNghjbalf1m1QlUMudKk6qr1A52bbsBYAsb5/
pjlT/EzoufhKiO0jSeX9Kux9AFaB2GJwAobjZaPf2gBuGEOLmOtkWa6pkRxF
snMPfreNgZcdY8r0oIyBdTIbEztObdpG5SvENOBbjuiltH2U75+ldn9K+bvD
0+Y2XEOe/DfKrXg4G9hHKZdgqWOMBwKwluIeTuwjJgeUIWa1k/dJffAL8fIX
mA0glUtvPDtvKxI+emglq84vVJAiWXgD5EsRrc2NSK4xFGaoU8gk49WlIQQU
BFgnegmuKsdtN8kuRL8K9mXnsfP/Ppm+UXVHKmkw8YAywoctkSTNOnp69QIx
VxW1E1GzQly0lySt60X7tmZHuNhPY+5zIYzXv2a0I5OpYHLS+nrF4NpeLWYU
4/EDg2tYGuJ2BlNlueAs1c5GciycE7h+i7g5F1mHc0HcoLUdg9wgOVXE48HK
04rAHe0IAvypfsylrskiTpjlVoTd9C1c99iXXgBf/W540eSkXtkbQfSsvV7h
MLuZ2uC77Z+7vVOQcPO1fGF6D5eNkqcpr2IihILOfIMhNHk36ifqxWleXLTr
Gw7aoeOKb4uech2XwDVSlnnxuMdbGlMcSn5qR0endl72wzgkLUb3TCTtyfnE
ZRynvHbNQhkHjRWmv0cyTP8wBfhZOnaI1fhnSj57D5uwRKDjm/l1xA2l+A9s
K5YQ2ovQ4mqJ7lBhI7giDPvc/GNxVR4AQOgmKyQDIBEUKN8pcJ1BH5vmX6C2
FUIXOQ2zAyB4DVZ1LwpAw46ebo7tFOvAewroHAMFwCHvbeHJ9BEU/bNU/PX3
sYHGt0dGFPTi790bHZxH1RFOdFeK7lpfbv4DRPTfrt62GHodoPOie7ms/g4N
L+pDw+ZBUbYN/w75Vbju2R/gvcYLQeaus74wM9GuPv1XGdkakeKMtnak232Q
6oPcMteJnAEorhSgN91OW8WdA35vYc7TxI2dZPXqjgi9e1yTZgjtTkpsUfXq
LyHYE4IhWpLVZ2ctbUwKc83uqEx60XlRmbwf+RiuHF+q0FJK047iTT+3m3Un
2llE4GFj3qx9lI5f0H3s2KwMVcdMgI4Mhxq8oNV/mx3Ks3OvIOcq1IpRpujk
1sZwNL9SkOmnxVxozlKVF1URtkTOxNtO57xlTd2wETPCcbavmFOINGPvj/aD
VlIeOB5bWZiaY3R5uzt+D6dM+4fNwRzmTWaw0uEnEnh6Jg/pwtgNj/8Q1Vl7
a7HU/O2rimVPCuhLQpn7Rg1+4pEaPKsUPf+vz4beFSTInnRRC7E5PPYHO9yp
JQo7NTYduhxAfVmWgTR8k7LNTW0LqcKtqLa+mq+4xzecyZjv6K85pXHSB2He
4J5KocQNBQzy/E0JpbgS52mVUPbdERCy0CeSbrqH8g3ayPyL7iEmL9sIzR4P
NwMjFRJ11vwZekdQM5+fJNh35H6pKbDtmxV8CbQ8CoP9CbECSvcftpljD/I/
0o4ZDX9jxlBjVksZwvHj5sUMXF9N3I7liyL6iJqqhovjMgB3mZScH9n1DL1Q
axuUtFQiESN8Q3uA95a0OG79bW7mRx1sX2UU2AHG7wuI0r0ngd1021vhkPVX
GU0MQcuZOQvWZx/m+z1OKfAE5oWyi50Llx9dFyoA6FzyVE3NG1QPueiP+Q8q
2Gtz34fz7cdOdcmLOm5yQB9PE2IfDZM+UFh95Iy4X1XxMRhipVyyt4+4g3gw
uwcos2YD7Gg+H/ZlWM3q2WX6ZYqG35dXwUh7Hk4qXe8dnl5b67OSVRhOsAcB
nUvxxIdZsqjsxpF3YFMveQQ2Gv7PfJEeK0L/f6pKy2F1DHTdM6VqOlbDmz3m
AH9Y2U2nIqZZms5vTa6FiwjBQBggwozu8ghxeFJ/XxvAF+lGuQFR04W6M4P8
Z/++e391Mdf5qtR994BL0Fivnoc2rwxPHVNiCeHp/GJxGg3AfRZmhjrcx2lv
fJmNvT8gCRtA4uFqFyrhfwocLoQMqLJ3EurFRlV9QKN1zGMikBfzCv5UGLJG
+vneajklTBmnUcafbKItpWzq310/TURYgCDoJEXH25qEytG0y5wXOGBXSbut
D+Iz9NXRyyTd/K9pk2NfqsVNZLSlRdoHnhiB3LZQJh0FTvCaD+eI25Si20OE
Yph2cIOQd0YWHjGHXCkB4CLufJLhaE/qyxtLYQY2nhOazK/VGaw8sIsIfJQP
Ovx56RtsZdBkBMVylhNdzkbKxZ/nvmaD/t9GLclKrDzn+piQb6Dt0VE+NKAj
JwbaAQtBYnun/1Hf3bfs6X33wno4Y8fBgspcU1Le5VvQJMZVwhabzHTyZc4W
U4iz0aHBr6Lev0Yyl8h7pZ+38tOi80i9/pnT7Uft7v2ak3g9JlWNySYkZ+h4
Oms5wnenGqpJhc4Em6B5Ig+lu5MVdQOg+6DttGjiKx5W3SExUNByuVFpgPwa
uetsuOggvmoCfGYDslcc1WDnFvmoi2Vva8LNU44i5QuyeQKrtC8W+QYi6RZX
1VAVXPE2j+SII+rXZS5THhF+pdtWfzSEgo68+GnyqCRtPooAL6yyuMk51ICI
wCmzgbdKg5m7vIz9QLuSEKKSniv9qHkCBBJzToZxDt5FV0nFJdEat8CqLiR1
TYhWpuqon3YzSUJH3KeZ2VqeIQGoBxk+DCRcu5nL8I5BVjW2dxuvX4ozP5J0
PzzWrK3grEh5JXXfOlJ8cF03t/CO69Inn+O/PBueqmVRRmo7uMZ6QxEVxxwm
tvXj04ArGaetcqmQ8LXFKtPH0ZmWQSbF5T59DgbIrkTFA9qOGyQaZHVMQqIR
+twAR3lQhffTliUP69oDgrjiBOBIv004T/bxCV5YlrQEP4CMcGwFRl0hvEM/
fXcjst5AIgMGMPwa0dx6q70LKJtnU7RNqjRr0FLFimMJnJUKnSu7lvrqzb8v
LDtaqenWbO7VBcLIq+XNNGYoR+dkuI02cIhePhGHGwwXvmFpP/sDyyuJUb9P
AMOwc6yeNfp/yPL+Wy853aP4HduE8sxZ5JEMh17ZYfr1cfFMv/eEqcu4Vuxo
DAit0TeB6LstInO1xliAwGjV6yNLXFXtElZDzBfIvco7kU9njvo3Rhuxlz72
gPHFK++FQXW5d4H5i9YAbJtgS+WD6R1VkdnXgRRDGFyn+50rboiUkx7HAZn/
m7xEtYYc7vmb4hrxcfnjxHuXTMIZHcdY06ya7DQcHc6YQZz7pxZsoGAghPPh
Wgd93WtC52uRJkfXqs1jRbLywqkqoENSBVdLnT8rurwaa1MV+M5vqWg84p0V
Hj44xHpKZ0AJVVNT0Vvk0dqbg44Qsig3OBXJxotdNHXFpZ4yia1CftrLgckT
kX0jxkUUBpZBhLHXsLbSLWdK6mxUgoFvEcLhW5pJe9NhiK472Eyy/rEyxK/4
w5lI+OvwgnUxLllvIPryp6wUsCpbC/R4kzXVYobIURQ6E56GwRoEmEDe8mKH
2ODE7Wrput5DCopTpVfr7UvpjMl8LgK3XNMCmUS8IbD8+9r40FqdFc99E3Ah
EfnCnOJcMuWHu5nT8JPbgK/n6p0XUf9jHK/O/BShx7uoFc9T0f8HHqiyarCf
HPphuMIZg/KKd40wJrEUpDHJTiNVRGB/yQsdm+TBAGo8YPVwbWRvwa1h/VST
jBRoHfrpP0136ItyogzMPGBAw5jTe3fjOe1vSaqjJ6AWLdaBsJi5WpNwRFpp
pjU43A5XZqEct1UCAgwMybcIRr4X1lufLrhrmOnVO+atN3bT+h9Fw5Nvont9
opAb3GvNqtIhrBwv0BNgkzxdZczKhBlaX2W09YfL+RE1KbGSt5f3R6mWH7fO
3YEYvQUfCkZfgRUD5t17VpJrZyc/HmSV2FKUaxTBOC0Iq5nlcPoUQaqLbrDk
D1uXbFw7DIBwmwG4sB4KAA29zBTWuWpVgri6lNGoIq9z6n0crjdHLSXzZq8x
78R9rm2gwxrRVYz9ZuChwB/iZ6j1CENKQ5NUhd1mCygofPtbTY7m81Fg4khZ
NwdsuWh/KFsaH/Ec4zcZ2LQikyH549araqyGfb+oJatAh0m2FBWdNX+jgUrV
Ttwu2//4GdOrzHKq6xs2O3oH1Z+0GPQrwEJNky+t3f0/ZvDeTcq0YtdxcU6v
Nxgn3HKf8eiPH1E4sdNmc9QBcbciY01hqJBTyPB7RYzw80QKBrF5pOWLPgBE
Zol8vf/Ozf1c+Nhvcnflb+4fQrYpGAe8mxLWobLwPXH7R/IHy4f9u28nvs3o
cJd3IYZ7rSSmbq2b4V9yzWzLSdc7eeT3ASje0jK4e+7wovBXXXfHh63AgzZl
O5kxC4dH/J0g4offJcVJ+MdY1hVwsUUgYW0/N6S7NrPMWIKzxMjqtA0GHIoa
SBdF4FAfpJMwXaBZVKazfdbZDhv1sfsYsHLdgySZ0VMDfc9yLgszeTmUz8Md
dUXYLmj1BZYypzeGN+qnIiXlyv7rdCQZPH0ukCCjKAOQhf48fBuJNCM8hdCD
f2FYPTwMhnN7wSh/UGZyEeZVPmEipkrZx1aOHhQ231+9Bt/mz9mtCGIDyqE0
x1z+kWo96rtmnmC04sdqMynCljraFnpcYwQLz9tLiIpMCFrlPSlFR5k63eJN
P7JxjFISeDAhHu1MJcTTbKxPjAsCTgEZvCwsePQ2jdDZQ4KyEfv9jrNOOnF6
ZKjL0Y4QcmMhFAyjOwPbDooNgbqe4cVIY3pPVLLi3vSBA/Q6jvIbKSFYASDd
FoyPUkt4/Jid/AyoOJIxvK81kqlBvgsF0F9kMyFqVs70vgfHDw4sJaGF5zWI
d9fPU7tTzm5dBhI8u6spYLW/sSmKA08oSkEHI6PYxmqj90Ns5Ni+sLPwJHQp
FHVLvMRtK3u87yAUIKWO5S7fZH+0zNvELjTbSqKkUKpsl/dDwbPl8zjsyWzr
RxXOjnbbfrUWdvlrdLA3Jcinqi1c9gziX2cgeouI/3JVf6b2n6aWx6aKV7Ft
/B7pz6v6qIe6po5x/qjSgTSBhQrujts19qhU8xDd7Lsfln43WpaPT1Lyekgr
W7KoEJfG5cWLOpeNdMMaYzxNGiErTcTHTeqGbMBwoWb0zDyRvnkRJByUth2z
66GcFa59PYBYk5BikGYzDEzFLPGMOAzh5Qvfz3rPiRo2l26Xpl8YsbCfIA30
2NhW/Oc8C5UxwnLclg/cJd2YjCu/Z/amgZxDFp5irYTpXdWaS0wSJbz0KdB3
/rcXQ8+X9qnXURjS3VDf4PNlYnAkvF0kGyf0/mPe0lB8lrY7qls1dhLbQZBr
+58kWk/uib2NznBZx0i/Ob1+M+uqnDg7oKKX4CIPFzNF2EnbHbDfOfX7aKsm
fCPzDqikSIRoEollHpu1vgDhswb6gExfdLACH3Sj+nAKLCHmSHk/LX4S9WKD
hinGwQsOfhfiZ8XGSdYKq/GqNnCHD15ZHekc9pGRdgiEmWJUfzGHaNpM1b7d
W3QWsTCA6A3jGa79gRt3VXJiiYpPsD6ZpeOHdRAX4oSB56WutL8wd+FHcx2j
Mno+k+MnB6oc/SwVZjVRbvjBvT+W88Milo4VKO7Rg1/B40R456bqcwk3Xoeb
ppR6z1GB+cIWgBFyL0SEOFccsMOT0hcq1O6KzSd+vXLlbic+1VG5gLR8rmFC
LLS4MSGt12mzO0gUf9E1e4CwnRxdY7VQ75CwiAYOvHF1usiQrDtEDmcppAM5
b38YsZW6Jo8nYwulANNtk9yAIKzy8lMMkP0KgaH2ykTakn4ZT26JL9KSkURj
TpkvkmB9QPl3ahMmclv3aywMjy0538HymfSJkourUFecauUpQCW8FarYmaj8
CFnnG2wcB64SAmM9VGZciP4sjeIv2pCD9R5tDkau4JYwD6DXG0l6ekSxx2hh
Q63vJdKAHMQe4AscaH7hQysQ9hiLi/wnWlfQY6QDldF75p8b4ridCDcpxFgc
zkBan8hHRhFi78RePx1GlRp7tcdu8fRKRjH6wofVxaNYa/AgktF2OH/8HMpX
9WTAOlkm5hh7ESoR4MgWOqNn3+TyXJOO4tXKxpPkeHbY0m8HCfbgQAjgSt5s
G5//1tHBirwEuFzIJ3Lt54qivtD1ehxCoJ/4eYj1FqxWs6sJ73BfnDX5gHkU
SOvOjqvVrCXmH/znER+xWWwkB6Np+yhh7ldfpa+5+iFSmcUJyYc65x0lr2xW
h1N9TOQ2CIM7xmVoVAR6Sy15IYgIQIqDwr7K5k1e3EpcrwVqfm+madXLzJzN
DazxzM8QgPqNoi43Vd40nw3muyLGrhiWomneizPGHJR7GIReJNE52ZMXpSzQ
QhsB/pbUGN3tcSurGetFWlS6yLFVDgnB2f4W379zWobRMuUK9/91WPfXTwMX
dEji5af+7ZdRPYfcWqr5m4t5ZKpC0EYck6raNGTiG+qgLeJoNshIrdEIFduV
n642inm5vWsQxO4r+VUUkGRcbUFnWjyp0t7OoOupQAhkyR6O6d7RFAAl4FOm
aGkXN9W1vrlWkaTM9FOBqDjcNSOOoKIe5pKW21L7z0DYUSqt83gKZXkDy/J+
QTozPSys/pn2glLcEmOsmEsGUqQuRClxATNlIfTpRlG8CT8++1jHEjdTLaiW
z5ux+PA8WNr8C47/g5usZDUEAC+QIzBZNEfzzR8JI7NWUaTLcDkdhm10kXo6
gqYVv3NenU36tXeJ3XURUDQT1h3AhnwSw/ymeK/ks4WIRK1suCCCW5sChcz/
3PS+W9c8w30VUoxsWIAswgGPieMxR9bfrXc8Yc9aLKEPygITpxzGMjLObk1J
NCYJ48NoXdpsSsQdhSLrVcGFZPdQKRxO9K0wuAluwCju3oXvgvsZ0yryMIe2
6b43zP0qRpRDg7dA7yJWEy0XT4M+Pqa+xxUYjjSnOurxfDU0tbjgELYLSUKV
etQnq555GKZqx9OBVIoRObpg8WfEA1VGg5Xs+6PmKJhrsfH5hEYZwvhUPtdj
eHs7GzGLF3egxiXrNGofX6Kem9uCbHFJl/CrIv9OQ0skL317gQW/xepWFJRV
eT36ngKBV8H/p36582mIKQiRDzgW6HuOcHrOpXu0Ye794JXhEidRA/1NWHMz
lkj4wh9y2O19EWp6EpT6VyJaIMxNDW74mxcZZPbbri+0Wzz9MwPMkEEdLn6N
O0p6Qne0hjTG5DzRXaXG5TVtX5MnF8byke83sswdhVgEO3HHCcTSQp7FEqfw
iaVOPX7uWDoLXhCCfLCxxJLZnrpmA0dCBCaJHxQEwJUWy+ajj1rIMbEDdQ2u
m65YUTNb7usiGOa4SXYOj4bVL8LzUlw0bRwWSwjdsC1SJ4VJ0HkZOMbp23U2
jek9zGyDfWJb+N6v8x4wyehFIt4IZU1CH83Yqyo8gm7qeqb2iITWAgHBwTKO
r/S5FQUs2NQ0s799EUq/n2YDD9/HFeQ50ke3sV+I6DgZTzPE7FTG+miMUjCF
+5rwOTgGVb4p30nHQFlMI/5D4w4kDROw1h0Y6W0UVVIzWfem0ZDxqcqJ3cUF
GZfnstUSzkq7Xdj3zUdfCgF9E2PvQoo5CM9My/Y1+5HJswDBSzJRGjgQuYJQ
5RnHrdL8rAJrYwfRfz81WPKQrOFm74jqQUo6dbpK1/KliRsAKoTxv5sC9pdI
3kyEx3xAFlTBDOHBwhIfpvsfBn/AUeuEuAuPd8TFYgriemdbkvTeaEfrG9O8
J+Xun49zhB/dcuq2tXg5mVET2iKLJc4XDWfKyyg+CHHfWOYeD9ZXVVdjja7t
IriDnV9yXfa0cFfVFycrHZFImSJ+xxvXDWY9Mm4eaU0ydRZb5Hj+E9YeBIRu
8KHGKo7hKwUONKWXvT9SUfzG2vasEVFUAw3mFIGEOkNOBXa+cyEvRzf3x5zd
PeZBUBA6bR5geZAMmHIEzc5JOZMhtxryY4CgAT9VvMwVlRbGOzgTyZiVHRmf
sGPvCxT/gkLb0V3dwp7hwRMr97B6cRye/shHAKmLw2cbPJ+83SjDomJPPm9p
Mm8Z8n1rnGDhrd1qsrsHlgEWY5x6tI+Aj+3jABzy1qhSfjfqWunWKHwdKJVt
NPSMp980AEZzyPb9N0yhp9XRr35F1kp/bIyhOATXCz/GZWN7d8MmJScRe64t
a+KL/JJmzxpV74e7qy9G8mC9CVbRkP/zVrF9/XRo1m2kA2UiHa5P5YxbBIOV
jdlwUqu0LjUWldRLO7e4Lx1FK8IJQZb9jx5KkxTqWj4Vyc7d6RW8G8sVnRTJ
VwkygIr8ooX5VljEW3HWHyUDCMGGRoSt3jMMPiU25Xh9ohiBDd1Hlzg/E3cN
osEXy0LL9HOgYJOb80HvFBfbWrawVVdBZCwnvFHLV4esUWbMCDlKc5fbAue+
tfEK+aOluH7wQXOqkTDSHOIVYnbOw/BuiAYnwWpZPCiPHNvi4klh0Gf/6v9v
BaMkOjSjbK2lSCxrqabN1isuknYgm7wCN5kpJPqOnDMUWci6+2A5Zrnz91Hi
pW1L7h8wJhVv9aNdboOlCgCKNKasLXf4IE3jQTU6dLJNJu+oCa6kQDZLAhbu
v2PDuIKpqOb36Vrv4aYD9NWlpXnmr/IlbGcu+rae2N/FP9ziMlB5esDVvL+q
3W9at9GqMfqLn0QVbFAa6VTtwAdhDgk75XoKP7taaARhFr4BKwKdlHrbI1s8
oPWkQFLDxzBfAZwAYmEZ8sfbtUtcwdZQBthQKmWrQlyWfOeOs0sHVPv8Fepj
yWS/9hI4LqEEZ8DEr/kgYY/Itpbv3121uDwZBOa8+GHbIwzyFTIrIW2hUReH
HFAuwhVrKbiPwM9vdRIaCIiJ6D8yr++XBy1Dv4IYR95kvvwPPBiOHZpLoML/
B5FxR2z7lukY6C/gILEsLhEHbVU7zR+OprGeI90PLZBdhYGArsxy9G1z+gdF
XGoDGKn5DqkP9/+jvYIdgqb7y0cjWVc93NKOHVrasTx7bL9dFVEHxTaIJH/F
8ad6UKii3tzj7jHrAWVH2jINI5Up5ff9JE95t8B6V+aalz3FzldIf7zY9q5l
3D9UmkwkBzhDFSWV0gM+hlplmxBPBhwoGkdrJJHjei9RMxGktiecEOx8PSaA
G4rhfvgvGGwSeu7mCX/CRCJy0vOMHyxpHGFlC+B4hlyqWKGx5leUxyDIWt8e
1ZTuihxsRwrlOXP98pKLwuyYRGI91xUn1w/S+Txcs20+gAbvgi9VCQmoldD2
bQfcUf6CJKOQ1tgK5OlZPcu1z58UJI7K50/g30y01Mt6/qtLEyJQNbmNGU2/
yZNBVxHNJeavbEWyIWAs8OxjIj1aLpq2gGcwx/hdWp1e+UUFu60udgbPPiEi
YpQoHsiIh6Pj8mM5GoZIvZMP1UCWlpPtNAH5m2yFea3ksI93PxBRWF/JK8RN
BoBaL8AvMly0ltiFWfXoO15mS67Z54xEjfb0cWGAqQy0TBvpg5rOgOvlGEw5
udS1LO1AO2QqYg6Au8qdBp4HnsvCZFNFWyRh5JPSyO7p8OB/lRVo+YCAyK+G
j1mX154QmeWOZbglGUnQuqWvO4Hf1nO3+WhcQ6n+0OWYEquiRQvpt2vWKlES
JA4K2SU4cE1Hy5dMocfsxs2E0K2Sbv5ywTDkxfQHCG+AjyuAmHMHYIXEUWZ+
IzIPq03j1+/TCgLCihWbk8GDZj5N3YETLtlq3CdpPpeZIVgkda49TrHVrf45
aB6KOD1E7/ay1wsLcFQVsm4xHpCYbLN0IwHVRTpOwrazK0eygtbmvCG2WLnu
ZsgspkjBWHnZ/m3XKYcNGKC8K53crSz7xIuyAl8u2p220TBj62gfswukuico
jeHalqsuLc/PGAC2uiI33T3Bi8uQ7JqZ0dk3/L0X4YcYbCfwuj0Aju1Uq8RU
PYXgJEg3ARaQmR5BUwnhEeRnGDlB5/Pdq0fHr3BKrReyET3onUhzol0HdId3
EIfC5Tnh3AACb2Z8IoXnripb3oWKQCjXKU+zxpR8AF16XugPr+xSH32eFqV8
tLMNeMGFg8aK60rGdJuxFnZGtD/6CnoPCBQ5GI9Ny/AwtN1aqrr8thCJlgBI
DZFEiXXsfgByZbWPlJs+Q4ylcTIAXRrx6uyk5n6x3fFVZxF74AbscnlesYmQ
8DjP87PrA3B5uzzO1LoOPrQW4xb4gHSRyrcacmGn4YUVavDruaCoDbj/ptr7
LpanLZ1SMqYBuQ5Z5S9HG6lGyulKYuwvEDzR/cnptXa6y2bnxjsbmPo2eA6k
NppMpYwmTP+5sReoWatlrWsXd4lYizVSRmHrAaFJ+3beGMbIAbLedCJRpQ7F
EHdBIal6T/VxEceSO4TbV4AJtv1GBd+xVRrmjy4bqLKfF8/EcwJiy/RzbWyD
DFJ6+B5pOt1ZaEYnlW+ro097Awwg2gjgQRSMY0+bpwQiWwpAMMg3EuIxiPZ8
fU2TTG6gd3KG0SUgkXFTeu+smXvFPY4MW8N8x4Hdcp3kP+Rf1rCFVUfAOKSd
wfLxtCudq8/fDbdcLkYEBOMmswqkQw73ToL6zI0WuZH5T1J9l8PjRiHr/ANJ
ubGxu7E4bRekwVBn0A2dF88B9y37wJWhRgwOgHLp8VvRaoVwUGuqabzo/3ol
6Vq73+8HZX6vJqQ7FGYLlDBZJX3hUalMQdaVq1AapYz7z7aRGseWJQKz/C9P
Ez8HM9U+av5MTPC9RVTXhvyc382hapzu9ARiOI3vB7zL//YJY+eimaJKustc
fFZl8IGwnjCCFvuU8JltYitDSzD7cDKBusxBoc4vqKHDlf2ULji+YzPkEvlJ
/8U+SLNj9IwWGXwRQ0gK/d3g/dZibUtJlsj3ER3VsGFGbksfsCAa11kJeYep
GFpM2AmN52mMJLdPzHnLZ1EF1OyvdKL77NfH0yjT9M/gYJ8jc3oZ20uVsnrN
+NKjJtSC3afTOuQwhM07P8ynt10ejqALZMO33rurr5LFrrKhhB3nFLAOPkbG
XBkLRH6L6wY4Xufh1h2SV2++5ksjsvIXNWuW1emhl+2a3PpuSmmyHHXnm3Bd
PvQuGvRHw1Y/xPZhUfvO1/hujdRIBfM7C3MFt2Wl4vxllvdhGTt9MdVxPcKz
q30hDMBx6w==

`pragma protect end_protected
