// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RKR4YYYb84FqMcS2mh+s9070lnXXOTrzaqJIJk38hGNGc0Br/q6SpmHMgDBc
erbBPTrzXAXXyswgWE0MJ/qsrqFtwbYJVjOUjIkt8Kl3zd+hhB72BKEbbvIm
zK2qlKivQKC+oZp8CGae6q831YePSXuvTZo9j1SMuxJ4h0zNw1yD1ApAc+x9
yRaCN2SmMg47emALIUY4mHTG9VNMUJW3M0knBzSaGvSIF/otsqDmo6Gj8xo/
l4eFp3OnlmL3zo+LRrIJv/Ghs6xrloCDkzPDDVyhakKwdEbniuFl2SopdZHO
ZhOLtfyDyWDqwV3vzDPNQ9sZ+YQM1s4yqPrNL2KOxw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C85aGeG26pP10RsDuKvJ1cKY5p1x4fJyj/wAVguEoSIsLisZ0JLj6p8YkG5t
MzP2Z0tKDrv+bp5gT8bzggE7wCIdQTTDHIq22K98RAZeB51pnOltZFMfA8R+
dbkzQDbc1T5kEeGsrJ4vuowS46eBwJEN5iM2NNlUnjluYyxKaQEdJezEMtqG
y85O5N4tdHI/30JvuUNQirElUitQNaGYLu45cibw1mI1q8T3s2jwrdY/fLqT
xtOB9CYmcgM5Ead5FxDBRziRY5IX7u9SuJAKuTMsDJHibL0NUAh4LCsSO4Tr
FXmI5nEm7/TFWWVUeYgyRJnMZcCk+/gey3bP33l+SA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ula+zOEzHvARvbxfnmnSZt4FyCQb6L9qNBLGrbqZSU3bbfLDYUKhDw9gpNDj
QFFtJVjdFU0N2myQLf+YYASjPwK0LhAJGiiG3ROkSn72cS/zQW5+kK/GrT3G
FB8OQvxGqSKv3/NavcXDVGsouNLf2Gewb7EemQAYlVo35aJ/uGTRD08fIZMJ
SkG6xM9rsocI0APCRt3lC+dseXV9gaCLtZ3onf7bc6g82oZ8+MiJdfGPMl4z
u5Mg/B1OWPI83/1jCi9D0ePsGieFCfxbs9wo8UP5Go+O05G5Ru9FtY3s5Uzq
8rDcjHj9+vS6jL/hfhMLmzmbAVQZZhuUipV5Fb/iFg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LqVfIIW1w0Br552FlJSLsL3n+Z1ZzKw2YLYOGHJHvbrogV4x08vQ8NvNSWmc
vsoFtsXV0go0fvHE4zRpfJMrTqZg6l0VfjVXSU907gXRQKJBr4PlM/c3F/DF
KFOpNjaKM5FA4eMICVLkF2MGgwNqCFiDctJsTN7NqX/910Fy0xc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nvEYwGqqzxmzhjQqM/reVNTQcTvgtpcXXGtHrcFXNSLbgTa4wEiNiWTlvA/G
060FeZdeWMK2GlCa/u3A4sNpC7W8Vk2GkbBXAObdkVEIBd78ag5Hzw/BzyuI
UP/IZX+IUd9ioU7ZkVwhKZ4TcDLTuI/NhDNHh3mnsJLAiEPgokETL9Nycx0g
ntzbeOJd7VdWJJiOJQXNEt8cCakXPKkQFsbMqj0skvFA9LrKQbv+wNBGOs28
X9y8QTquccwNPHcTCDIt2JlEblqP8t1u/4P+gevby0BqnnxxDLKLQe6aFc0g
tab6BGuDDHvGqva/fMwSV44WmW6Kd7nyZMPgxBhsApae+WR3xZ46EJ5JHoU8
FgSP51a0cns+FwA4aaPN9BqjjXQmUgt/OxDv4JhQV+azpdErHsJtmoHUuoyx
gA51UIPCsrfxGLEJuW+nxXcoeR9MAFp7leJMagyR5qSqK4LFozrpyE+7ZJTr
N7To3iw1wCiqJXeW+OLq5TW2wlkbdieV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RzOl+fcWBMqbjD0WiFJ8njP2hcJkEQMkoPypjvi9QKGe3URhdLRS/9i84Ev5
wOc0slXa7sZb2i9MXUgoQ5i+uZaBhFM6//8zbiR9PQ69PqqpddWEEPMeWo6o
tBZeot6oDJCJ9ljFuDVBoanNtHgSlh1UgGt2lBfL4AFb/bBgn4Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a1Tes36H3SkWz8uqW467r023MmmSxsGVa5SlIQR7Ay8gd6ytX+W7eEWTpH8a
ommeS34646+ZObrCI59Gj95AU8YM2PDDdveA7JIx6wY1dmaDRGevfbzA2zyQ
v7GY2dUzonlQrFmvlk1RwO2MWwWk5+XxQcCXzhEdyW6/MErbEJ8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11792)
`pragma protect data_block
rnJ2/JzQje8WhUwcwCZ8ayyDbyRzUSKQdEx2dK8mMwJmgCjwKJUMS9UXBlI8
l+rvoI+v5ACQLTzhzGsdvD07m0YGn84I8KSfGKLWGrlar6/BEZaFLeE3w0ZV
DYUwFI2+QFFO6RIZoGjGBHn0pIMFdIdVeFjjRueONvil4WyX7tgyAx8X+Bl0
otyn0XEWPkOEfYe9FgLhHa66Vg+hunVhzNwn+l6bBV1tlQB33SqcKScTsOui
WTJqZF1Ey6KDYx1ALIUxrxj3yJui01TewFgxHN0j8alLDdYb8YwIZzb6OVDo
CFGZVR8eutIVb3i5fzeO8/sVlshDpUEmIa7Xr/A3NCfxG+9mQw+/0Agls1eF
yP10O7MSZGxzGpSS4Bvzm6xMXOUm99GMF4DNfbcOImPYpgIy7VbeYc7OCHY4
R+X9kKnZBfLIdsSI66DDJc9b12dsumjhrcszoKPg51lk6z4e152GqMXtb84o
9+fG5/ff5b+J6ltpdxdBHMwxRL2npztHqa+WUA3k2D5iGpRTgROEL53JnO0x
g9RpYc8EUrCQJDYxJd9VTgyVCd5B2P2CfWUeL3Cw30YzMG8tv8w1JCgzQo03
rANtnOYpy8Wub+wj6R8xS4irEFXqTREcjo9R30wGT0CWVyJl6LamU7WhAt1q
7/AP1K82qMPGHZB01l7brj1NGWhN42E03fORLHi9kNa2sqKuhMVmSekrusQl
Y+HoaRlkGtiUKBU5vSu5YgBaCttnMH5phcm2eKydCZh+9Dds0NCESY3vAPjs
piLtF0039E+qZXXuq2IAnFJ2ig5hd0ik6n/SIq1pjzWYpNt/94y6lJBRbtXI
mENZvEBI8Sq2jpkam43eptR8DLU3ky77zzlL3FmAL9UEAjNsG/rzo/J7OwoM
2x4qYEbmkZ6nobAHiTCIbL+zhHP4/RPtWcM1zdTjCeTw/P7ZS/1b9cfHVmP/
Cs6jQhohLqCn2nQBEkFLlUv79TrVqf0AxgvOcJCcwK48O+S6A3EXGJ5l9s1r
FK+zkffzyu9M1fl6vgvOB+VqVq35gPiXenVbilBQC13tV3T8+ZtNJ8E3W73G
qdr5ELninouBpb/PqPRoVmnRi3twWG+RBW5GN6pIWV8dJjjAXHMtYv4CTdXR
83uOUFFzl6cxAqEAtXvmcyaLkEZI7/VjFms5q63AMw96cl/Kfjbkjk7F2dHG
26o5hpFmwiAvJTu2r7IK7AQVEZpJqxADVqpzWBPeo5UX9Jnt0xW3z9tv0OiK
sAvjhE9TBu2jf146lH3knR3psJemhGDZ0Xcx7xML8+zoUR93MzPVSw/cWt1D
OLSAJLCYtVFC/QFk8/QoUO942VL5dUBFD5Akg0+pCW2Ty9t9UYKMs+hhMm26
0BHHPL0cKCXNwCmoNDidUfeaIXNAiDrzeeyUw6rrjAoR+oR6GAZRk3BP48I8
6/UZmMxGd8pc67JEMu7nUIrt9omev0oU0ruODP7/5AGvvvNqNtKBwRQbLO3H
2lB6ALbnuCafoktKgH4aVuKIV4QCc0AeukKCL4Kt+qagpfnI5w+S2WiGgGjo
2Da3YgsNoaoa5QE790hpNk+oayO9PLQqD+7Se0n/1i2dhmu9WPmSoAOZ6lCc
ptzAM0dvqJ3FcxCl/9o66zEmsOmv1vA4bgl4LqVk6OZqIpDrtXeoWk5vz3BL
4dn/1xw9cWfVQv89mkSZCcVj3tI3lj5mwgOzQykvknURMS3nFaJOtigj7UNm
qYFUPnx69APDkqUafKdYGZiQPVPQ0YmWU9L83Y3gz+ff6mhSDc5ZfUtLL43o
Hrrh9pfUNaN/So7vZq2L28P3cUMhAU/XiwKGAukOKghaxxdZtu80ZKrUaAuP
9X3SlzJxigprNjaiCPVPmNzTorNk8cF7cvUhYEtg7Nmih4XurqKvmPc3xpI4
dBYzdQzIoiLxNNTLbFG8l8DL90p0Tb2M1ZErQkME2mKoQ/0lY+YlOsOZzKl4
TB1BBXKYYnIcmLgLLyF9td/Ivs8dXz0M+qlIyma0kRpGyEwUmoniYUayItG3
daxj2b2rPEfOvH3l7BafoAavEqEkHE15YJZdHVJoLU0vIc3vIPtvxT48gdtk
h+EV1/iNpwSmJXsMQf408B/6ATLcU9zs4/1AoJ/5oPFInsk2d8lOBMlRjTa8
92WOOjr0SpAFsE+75TSuBxUnxRBQTkek9hkVxyogt1QAUroLrKL8mqSJS2zT
0TpRw9G9rixoWpOeNRHkEBxgdMiB5WRGIHiY9Fsl1Po9ZZK8xtjCTPiPoUc5
ae08sjaE04s+DNVhYtBPd2GXuDnwxK0LN4/selaG20ugLXGyGTVaaHnwn6NI
NMq4vBYWjQHDe/l75cdDQAsEuD3wvRwxl816ma3+ouV3bD5/nfA9RL1nOZDS
nd3prZh2XZS/vijlPXDN6M2KkZd9v1WKUqLjgStQabTRZhMOZnf4X23I2Eaf
L4dHKVSnvwFzwgfiHA4Iw4iHrbiUgM224V7eHWP/JW3sKN7W9Muwr4ty0wHb
V4eKcYrbwX0z78sxWnOyedDKBMVC8/EomrOgaCUEQcE6ZXdSMHGQ4LOcTlOS
LOAN9rtqF3HzBXgUsDwc4cmNf4qh4VxQrQgNfnHdoPeEikrmd4qKQeK5kp9h
klazHRKWulMMweRkMQI2vaMUH6JMnxeG12VFteyD4t6lPU++/aOXLyUEDZHc
g4H+feJfrsj7nj+wkRjdP/abTDe21/KjebH+2nmXCMIVfS1LoGJPQ7z87zMp
9FkQcXJ+lNjJGq6AHILkocCGotTEgv8cf/3WglLWlHTdynTD7AUOfiKqrZkx
+EdyygLO2rplRc7DwwRJLqYc5H4mBLvdJEToGJY5HPxXBp/Y2GsaJZswuIuD
xM6hF13jkGmP8kVTRmt8s4KMJUM0gUqdJdPw7tMOr2WGFuiT06JldDAlYbz8
u9tZ1v0M4mKHsZPrmg6lAmZfPEmcoF7m210KSITqJyui/1IXu46/OzREHK87
+RneHnazSxEcR71dHW8T39dqjaZPs7p5SzPZAuWiqbh26WD2ZYvGqlJ/l6I0
HHThNNh2iQKRAwyHIcCAWmvf2GIu/MIWVPQC0hxdq1JK9EP45LTOrsbfRl4o
SWu+xXCEVLgr2DMiKQg4tYRGM8Efnv94pQb150ko5zJOzh/t3t2nmeo2zj6B
80UwplawEqT/T6RQdY8V+f+XNXeSLj0Q/u4SGRErePBV8DDqsA/LlHiIK6Vg
kNyS1CaHygvReTaym6GlUmwOelpfza7Dlpoq5cOU5z0bbgvBTlkkB1gBZG1x
KZgBlQ0e+jr7xp2kV3CQQsFfTbmryG8SrPj81HEl6JSSHQgk9WYKBSOhacBh
mf+Q/hZWQb5oR0xL06UhX2leBT7KK+w2blfK6e1wtuUC35ck454csV1eVqYe
81/6qR6idPEWkPu+W3TOOzkvtzMxp0qbx8ON0waGerUMxZ39uewVyFH0e/vt
Rdla2rm/zs5pchVqtmMru4NiwJJ4o3IrmGJHlJc2FoMJUayMwuw/x9C+gXsr
umECIhF4PcxtRdAjY7FsBOFmq4CbxPzgJvFgzEGra9M35XN83pcAUyq1s6rP
EBM8x9XBzruVPw8p4Wkl/2mIqw06JcB4lNXnx/xFKNCyKL5KuY4UGtuBFdrP
7TI98cx/s4yDF2oN4kymSxNAns7YFSH+jHSMf21+VmlkSJA+beI96civfn1+
yfcPSxf/+Ch8ccbP68JHNeeUhCQDc/564wnMstLDopdLguN/TO4/aw2YxEig
OElmiU1t1IDSyw4RRL0BvAWuhraQidcN6SexPRLc0wRWwGHFRghBPgtfRR/h
/PD9IFSvmxwVs8i4pj39OgLRcOO4fwnPOKelH4cp/6AkzCIpeNSfxtO+wdkO
WdRlwGtsD/dJo/97Y6Cjv7wZWeP7FspuX45cw8ozvIcqb9ZTohG9PKnvhwom
09Qh+wReweHkLirU+Zx820wWVTrXLy5RdZB5HbPm+5lLs0/+IuR7hBnkR3l/
ahPvJb+/iNxPjavvOhksqaQ63PJqSQwJpW6pko7oPvMR95l3MvuoTIEEsiwp
rFnN6ZhjPHJjb0uF/DY24yvBtZ9TwU+7VJGWo+qAnao9pBks7vjyOy1UxNaz
2IsUJlGAhOwN+cNBjtn05DKfI9uCaQ1YmkOfPJHDtKWOFPve8wkntQGUMTP/
gnASmaQGd1qhV63ZKnZa5TZtL/4sXbYTd+ntgLKYLbfIDXVh/XdG33WfW1Ll
toMoHXwijrJThvLVSoIy5g+e7jwgM2nqIOGyvvOjuTqLJcO0Ptx8ZtEkAS4o
sLMKiOI60TUTNCFNk6lnh0YKa+4K6BcT83mj31fZUSpI1whU+qcrI18yAiuG
Eivk1E3zDoYFzh8FPQzzESRp3DKzXacB9m76jw533qz2uG5JfiCZlVtRt8Eg
XJTtSbFqMlVctkPXK1lEjoDX3oKz/M7I7+B/+4pgSQHcnqCGDT6HpGwcNSEI
oZdeNeT8WLnISjUTOXDnLg7rm79gj3OgkX0EH3SXvP4k9AnDIFh0BfS1Tv/J
bqDVezhVHRsNyKppkJV9BtXsePVzngl6RqZMZTjgA+FjhBepzYM3JgSvmAqR
JIYh/UlQGVl89mGbIjgneu8jO7rTzF9e0HldVLuiSzZdHLgngrcgUxGN1fgp
/9BNkC8l7ylyBofTZHrwqq6ZM2XrG9XBQwmxmGY0z33thHLJyPBVAQVnCzdZ
GTxUw8vxP58Iwi11msRkEJSYNTgS+fTuwoLorNgaXqVHUVtb9s4mDRV78nw2
ChbHa6yHu1csHpcwUCR82fRakPmCRud7WWnzklHg/T4HcgdQrO1eCxqMOCCm
9cwYaAAltLVo1rDVJp7+p1mdwt/5YHphYkmeVeFBONNFT7Bw/N9VLQwm4f2K
EN172dTA9hx9/RJLA12un6pvBcVoIuDk4eqo6GXwRhzM8mfxVz7f4JtKloeN
2eg+Kn2naHc0x9dBQSob5dca42iwJ2K+7ESz2lpxgpaO5Gamg8TkZGj4VPOT
7yS3U7/gEBInz3nXsCSLe+gZD5q1Qzj6BODAD2adYh9BfwOxXfYqf8e9qMui
2IGzHXQnEMEzWbXiMnL2uNrFGOQoXiX5ufgXkhVrNMIUupLJaHgHrTvrVyja
zqH3+9tsSY4GwtJJqzwBwPsYhrhtxeE4fyXPYnE/0Ug0I+ajr+lIGP6/bioM
7VK0j9QRbIOvUcgXhC2F94H1T81v8GnagiMahyXlH2hoVdXENPiT+TYVBFj4
VUYASwtnZqe4JamCzN7McNlMEoXv7gdiJ18mth1LtNsMu0Al1yuhnQCwfEHA
n409A4/HuoAG2uZNC+6+/hv7DmA1zJurFd3hdVkVNXm/7nWLjImwB665nHJp
txIWUD5H/ugntHuF0867FyySpK2AIKvSDyndNgJT/vpQIoVq4dGqtRj8MbBp
IqXgmNRr4u83+3UxUty29C7c66HnI8groHwLhRT9oZgBx3/K4U4upH14WZYJ
UVF98XsLk/B5j+3Bkjo9CnucewVJ8utWmo1oEDloLjorPbwL2lvTxLmEGGbC
dDMSK9EErOrjB5d5jcp7Hn6uKE2WMVu/bcvHm3zs3/G5lQdfgGMBq2ak0Iet
6bwYDNCwe3SHaKFljXzeAHMfZXWNjAS8CEQMzM4CQ2QfhVFXw3uOZ+x1ZDXL
BEOugaGAb7qFNrjoho/zhbDdO79ngjg/GxFDaVXZQmZfZ0K2xPqwD+aqu1eE
moTynes6/0WbJbEfiFMMi8bFvm3wOzqJh6+f2IRmNeeLKYow1uy8vuKauE3l
X065r3W7+hmBB0XsdiZNQVD6zLkojhowIa7xz+00UMhlolHuuiDuXSfhgvas
H6KURll51kJvsb/i5MIJgQNkKjDg2VmG9d10JVsyl+fVOseOmM0ng87wqOPI
VjO71Z50vDDtUoKN2lWcRbsNqnsK4qrsd/Ky3L6D1KPznkyB1i+FRgzb016J
CPU6/yeWuAyfLyhJMFV8+xPQcwv4HfmlZ+KAK7zJvP6q/E23R8cfPGf28oO2
IeK4AGbNccesIamuEX5uoo40KMOXgEooRzM8JN2QbjpbjYalt2gDudBZaAFJ
xC57qYtxXMFY1AK0jd8DgwVrCELl6tiSUUa7jrZrI9wKFjcZ7OGUiMlw31lm
hbCwN8CgJ79IDnJiJRLX3YUvCYyI/b+64zB3WqmW6f6GOJOQxecnzxVxiIGJ
EN4glYGZZFWECoXPrxSE92HPm3SpNUf5oHcjwt8ys41HQ0+iXCk6lwyQObAt
jobh3LqOFIaTk8pGso5eTm7Bui76wBFvba+gbYKWEvX/6V7OjUa88NtTy9YY
oM5jUFSAz+h32ghv+50ohKhZZmbOZ4YJaF2uegcEN5656QJdNk59nwmtzDHj
vVFDNbsy38AiHjUiLO0IHNqR68/XQKvkHca6qfU8sNlh84fgy0HlEbUf/HVc
5NatT4t2QtFh45do/rCSvahYbZk5CdaFQGedOOqOTLET9kvDVjH40H2fLqjM
R6Te7RQ0tENC8HpWFUjS/tYkQjdyrIneyJGF/1enzGfADwunhs/4DIdfar5b
QFkD9YTiQgC5qMcl2s/5KMBdQuelTpE47sl+H5SU3kigPso+dEtmdytyKqGI
eL56FseK98tG3ctcIbEZaHshd2aAaN6XVXKl7RydNjLvXha5FbdCf5rYNavu
iVvUGuO9ljpThy3eozQOa1lJwaCFF7orW3Pcb/sLNetpf3p5NLIqM1zsISk5
IhOTpoGy6ymy6WNgi76yyqiYMDJjO6jyX3tl/rCmLodGPoeVZjkU/qJfAI2W
8xxT4hBVQhjPkWecjApFutl0Y9zJ+SRcPx1Q+nOXJ390GtBqT+PqxEXOwG1G
O2fPvTANb4RNr+v1nA/0x8Mic4LOr4oIcnUQ8rml1zazvWHVai7qn6hMVDcu
NeIqUOJ+LFRsJ09aygl0U1IeIIVecwTX6ZcVNQhms7C4f809ocEiCkATipig
nSwmtCp19f6iP1kDiYN+Ny2pTkEb7jyYuxQkLlNDw76FB2HhrOkRcg0FNKg8
8JyrRQcbRQ4w8svA7NduNhxRrw7FOQ3HSVk6dPaZmU+zGu3boanFoussaQYJ
10dmCnagcHpl8034V5kYCX3zMjTbFf1D1AosMyfcaQCwcCNLMSGIbxbABNz1
+DtyP02lp7eV5FBUXEP4Ieg82DNuINy76FAhdO/qk0EkmZUDEvyovwddDNgr
H4solR/p9oBo4RwPgG9/ocyX54QLYWVNVVoPCULSlSrjh4KlVq5UJtHh4/Sp
Hcb5u9rK9gCBCDtw8YbnbuXw6pE7RRCRKo/0SNW/i/blO9DBt7ItDFjyKuHa
zpeXXxsjlVRvTibHNG2iEx6jivxoJ4/rduLVzEel2viZpP6r/RBsBUlrVmJg
VCZC+YKFDlEWwsyS8tQyLe7JSGOgD8XylrkPJpwA6OLc7Rtk3/VmX27f5ehL
aT4KLYRY40SIGvYPX+98Km4qJNF8UQA5t+R0NExYsZahNbbm2wfpw5ZVWCe1
mjjehAMtnvZjsHUhiDisPRmHmKr2MYPvlYWXsnPkdpVthLoyVT/7n7hxDrRH
3pnO6Y9BYFK1Q4adhWs0AcyIRAmWS3mXNek8gmnxLqZf0ApwheVGsneHB0DI
YmgV2R2XBqXs63/smWX9hfuqiDuK+JpUFHdbslhTXkNAkUJuWqNqWLMtxpJX
/fftlsya/0Uk9D1lS7LldToSM+WE9QjpqX/3hgiqcpkDcppGkm3an+/6bIgQ
WJ6l/ejaGRgb6wRLT9olcrAo679NzfQ+c+Vxb7SQafnfouKL6iGnAUTiFTWl
/QmXLX8p9VHhdAMx3tfgjmf1ihjFLxN2weT4iTARuS57ThGdgxIunNcH9o7a
eKXsoH9tc6+icZTLQiWmp7m5QDOxGA+q3gd11P54gAC4BaRaJgGO3mkc2QhA
rRFi6B02qk2BuHegf9b4yezcyo7yMP7fcpZ6iWOzR9ew5Ke8KlQgDTyEsY+V
gqtBCxlevfWak/sP9rZt4RrhK1bm+c+6U+gJ3ISj2UMwmoJOX8Quk6DikvWr
wJ6I3cxwYna6HAdLUmjQOtjUPfPrhExa3iveNp44ANnqm30h0rezVsppipLL
MURJor/dXy9oMXpDb7ggkzgX/5S1qAn/bOp6dMGNs81OSU+fPmpg4P0nXk82
kf3Jg3xI8XGFCpJjpSQDrizy22gv63xHF9BVcVC3Y1qr8l4RPvtSGP91f4hz
rny1HeEHkfZpsoNxYw+4Kw92K3qgfK3UwChNQXv6CIPjaRuiUU5zO8VowgWo
q/BksVCsvikfpCFf0XMxnBzloDjz7QlLBcHHe/EyrULzEj7nCCV7Zse5Up5o
ECvOVnlt9ai+tu+NhXN03iOdo41vVUhBwf1Cf6vFhfWHpY6SleZzXWK4Ll+7
up2jCcNfCBn1ozitdoi8Z4H/G+oWnY3d0aVLsDanSPwog1t7MCyGfXdZe3Ld
TFwxInMQwvLhSJ2CCDkHb+BDtvR0KNweuZJ00L81mqPN99koCav0NorAlK/r
FrTZjnpxiIb88EMPI1lhhcFiOjmHkIU/kixODe/ZIAQ/fyJLycvWSObWdJjZ
u9EYzDSYHncIcgi5ACR9irv04pWLQIqlB8MkR5lh8/h7Ifo4MFTG2hKsyQ9X
cUXTp2MIelzWMjOCJQixQriPJKPRrmKLi4Eg+lfk7REbqGr0wFQ0AIsWEpIW
G+e8CXGj0wwEudxn79oXjg11htmnkkVMnB99vsMqDuXQKXgs/LFFkh4x6C3d
2zRwAikV/k8vMdW1YY1n2yYjWeo5UhLXDAFVsxjklpeG6Q1tdyYq2BJCMEXR
CKQfW0x7mtHwRlAcvHYKonGCxf63AVzVJ9H7R+JLPfBganT30lXHojageWma
r95y+uaZZuZqKs/NXz3JZ5rQA5H0gijSvNXb3Ebw8YFlkUCf4wplqlKJihzV
ZSm3fzP8c1M2sAnG3TGkpL8HBkwsktBFnRxmmT9a+jdXC9PoTTuMfP9trmvK
JpjBxR1KUXtG61bMIfBZsvHLoo7ccgBtDYrlwmgbKSVygxvNjodnK3eEhNbv
UgrZlNxnXeG2v7TKdBVZr2d6/enlzn0/gphEtVKHXaAtNSe4f0vhBKdz2WCn
JwEOu5own2K9txGeqHbue8QyERZR6o6rqwWwoe69XFcuZb9J92mNiI+l+2wc
7QRR6JiGwqE02x+KsdKjxzRB5IzerLDXS6AISRsFOvzVSYiFAc8L+uPRAYEB
0WC2gx3wwIo0cWtKpSoK79/F2BY6Ttg/sb/b2EkKl65/e6Kdc+H2rjxbvlbD
e+COosS29CwKBtQthmuXpcMUXef/3lOwz0pFgjbAJUmFtQ3/pdbvlRtvevrc
rL+8SeKdcArkFMzrMVEi4CYnJSju/DGSqxwUbf2HfdOY/TdZTN3Su1yOSvYT
PwDImf4YSQWFbFZOS8LKv4w3gnCQBm+Bhpj0FfXXNax3VkhnKa17PfkZsw6S
wXjIdt/2XoQeyJNM1OqoJK4jeSINWutRhQk+sAzFimeuwvk/8T9bz04ErMdi
dfLXrjFK8othBmQmYR2H1frYUJKThYPetCTTyBBG2CbjDH2wLOaWOIYSursy
5tERG6TePXgHYr9osjnpjzWLiOESYx0e3yxbnCh+g0JH2DJ5jqmLfFukecu8
Dm+zhaMMl6PHAH+8Jd4Mgjo83GvLbkyw7CVmAADgF2kHDt53XUENd+p077PP
jQT1TchTReN+PnIDF7vgwQOhQXEjyPHilvKLvXedPfHZ2SSD4fxsqRUMm76/
WbkxebRQpZMstHVYbcpiMC6LcOb40QEAGrxhQWk2NPkgBHO/8rdDHMRyku9v
eVIUafqWUercY64XI9sE0AMrOXYG0v9dortBEhm3i8gd61DbC6ZH9wFBUi1z
bR0pA+ac6f8oqzaeaQzKoHXOsVt32CMo+CQN7zg5iicYdiqNlrsJ3xeOEdDb
pEuGbu+UbnBOSaUnXLWzJOxTLPDQJDYpUtvx1SLasmhWC7ilF0mmVs/Xa18f
uCJtP9Bq/rTOaULeFK0s/N/MLDjwnoFz6nhXafmh1tEwSwZ5jLRG15dUESQf
RfMwHSn9RrGZ4R93ZgsKCRZdk5SXrEDg2UYtNjba1QG+cjVCpbmFKDtHpJCw
ogmPEUblO5FnU3t0hmJIZA+RQrZBJOi8y/JB6agGwu3DpPD8YTTpoh4b5Uqh
pcq41fF6Lmnc+vp4TH4q0sCpLGuEqr6sdH/CvDh8hTGGQukqHlKCCxh4PgrO
WmvdNTsAif7uWfU1yBwJDsUhlWqJgdDRWrL45cbMLHp37pZkoAn9hXwh2LRi
buJVgr0do7kJtoNemS253Wnemu9YipQDqcSGHdRta2qbLhML2z548JFI8dsU
QHR8VuegGNg26pASvkpJYg1DbTUrzUJpedZ0r6BkZkmD+V8BvHAPPWIVMFUD
I5EDwai/Oje18jkVTw86wSA/EhjE15f0tJZ9jfrh0KVla79ixJB4sRAFnFHv
hq/s1nIIkIAsAI3At4Ww1s1zNvLdlXPzx0D6NEN6nIMu1xfvS7s9tV89lByg
sGfNSj9BuVddAofZlxt9yJq6LzDN11A25+m2ijeqY609os80v8f0mPYWJxvB
hc0+QQ+4uTZhF1KPwa3O7fanfCDYbtU2QNX/0e4+ccUTcVeAvfEe7UVSJuOM
zQ7jeAkyJDE+AyeBjIX/9b3YIVY1Te01y8qlCyHMvwZBccRGUr7Sh5217/q1
WojpHZkNnftDm0PZ7fvIIKndbtc+TyAncfq7xtFHKjjeVznmOtdCQM4yb/eP
BPmUJYSkFxKIu4fmDk1vonrnAnY+tjgZ3Be8QKQpUCpKt+A7dtmf/ghlQmMe
1YN/pVKU/lsD/0KPSzcVPnCoPzkj0JYaLavdd35T8iaUtMK+wi2qA0X0+GXK
FvthTnPjMse/1soVLaGRjB+qGBw7Y2I2yEe3rbdbwCsI+KW6io1/A9YkKA1G
5/jaeAcHRF0PcO8qJXBK7R0TWCtd/aNtCGqn6Z9UbiNr/M95gUMO3iWPHF+y
BJ5UOVGehWvWrSDQP76NFb0hF6QbTZyWIgpzNg3d7M1RVD6TOHoQi9vdWqOK
kyohvqPfRsi3Ds1eWHiU0RiBJhRGpPrGSYnDMtOU/VhB8/zH8U4DuBFteuzb
MNQPtqEYbB62VZvwQ5nrxRTB//yZNtoDX7CHt2Mep+AIK4GrHnHZP95pfiTv
24l2GM7BTrFWv1oQ2qPQPVQuV1DakaPjL8eO6xq0nGfC95qxfXs0lzyGrsc7
SGUP8P5Q+Coy9GeLh2EWGwdTd0KKLtBsJtldevZ0kp7U2hNvqqCiXDJWzpB5
mcVb9LFmcavqEJA0lPIiJ834EXxlRASd0xVKKao0V5ZPk1LqVH2jdPH3mbDD
CiZocBtGdxBAJGNAT44M8egNsngBDR8Yiu5w2Dhi1NugT8jzNSSyV+LWj+ON
fjahOt52M+BoeqyT5V1VEL/ZssHmzLksnJC6zJQl4fIY2vpYnPpvZ3CA7LMm
OPokyCVWEGpMtv5Dy9+Os3RXEAPy6b9ojVtCb2+vCr7mDq2U1BXPya6Vy0JA
2frnpbCP74FVCMVq1jBL9J6sszElF6S7beWkw+JccoCfYfXvHKs0VLxgCixE
cu+SJ3c0sa2TIyaNDhteGEABcPjShwSqLOvwRlyr65qSBoqDzakib7Cqbm2i
qW9fqmnx/hGkOt12pZjB8rveTLqQPBihaYRdvGqlDoVqJ4Cfj9gLLqo1aEWT
dMveR/tDGW2xFigRY1u0PTigJetkM40Hy4igg6JR2rkHtGi6etDVbgr2oZOG
t2NyfLYIkLOd0jQDevrJ9bmsy8PKkjDlUypZ4ocsbUvmf9kE/XBuJFTn+HS6
3FCbBm9P4PQgXr6nae3rtxUXTU5xPdsB7pwpWEYvQyVrCQSCdBqNr4uARhJR
yNAkm5QCFmogz9XwySd7psUpHJnB8h2UJnN6IZwk4xkETY7jNxHwNDnNQcgG
RpMFlhIlXTZMthpbTJDoNqrwvx1Lq237q8QbF+py4tQlHVTvm3sL8w4nQ/ro
IgMEGpr0BbAJ9QAgnGkauGze/nOdObMR3Hp9DhehImeVsynNHv1aQK+OuLdl
KE/ulCvASpQd3TYvB5cMcEmH2Ty4VG29HXRLRDbrt3Manr8yQC/Bk0JwzJcA
Brv9Mpsok66U0/DTktnatkekkd09//jaMU5wM0Z5hm3kjSUblEHtcdecyaRz
Sxh2tr3/UrWYzDzdiQn1XAwpOF/vt5uYgGTqGN+VibfVAZ4EU5wGX85PeUWN
qXnlajrr6RMgY4ccbKv+VFtY2s4/iE5+oAASRKohHhYxJ8bhjMmiMr1ZhnkH
QRso5xvKeFtDosrx2Bsh3LNLctGtrHREIHbUAJp9flvZtdmw9pAeSRRfmTm2
uPBfpyJ10Bxi7En/cI1Bwbu4BkwWL+qNrANbkd5SDziKBfD0FBr8SG0volFL
vCcP5m+R5YvO95Q5Kv8HkzgCk6bYs6i8sJrdYAjIqpI+6F1OhtflgUX/LTWo
4hrSF2CtHPhQJv2lDe+6ST/9W9IIqT97J/epyCBX3fswZqFm5IzD8cqvtyHx
dnUkCeuNjp5mv4GjKPAlR149fqWu+wjvoPqxu6ETKAOwKDzPE4JHgv6NBbMs
bHgCMPO5S6yLmV8x/Q+T+9LNgOO3SrsulvfwgXxnZWheVnrx1mZxMBv8hQ2R
rwgStvJYnSH3z6qwVD2thJZGPIfX2H1lrdiQ9bfjuH/hMZ5BLizanOxDxBvJ
y0CjCHqYava1oTTqZtInkAfwJvVbPl9M+vOFsoEPNY5g6RgwoDuMfiTyGmo5
I1iMQIzgPHjFq2SgABznNkMD7weBicqa/2P4IiiaaXA3/T1+oyZK+71CRieb
8f7A7XOYZhqZf92lT0VRWclpq7+SLjU1E2VNw3WelhNPxBcarrVJoseiNbDG
QXRRxctbOHcQI+5CuwQM4yDO6BHoqoWMXS9bBArYvBrZwv4TooAeGXhrXh8I
WAcHtOBYtYbDmkXlvX9swOkZI+fOdBKScQoxTSxE1l89E2cN6LhoGMu8t5bs
zpwX4vp+0eWB+UvU6nzxWSKkbDT9Hz6GV+7pUxeXFfNqrFcWEaAncvXogsVv
Gqo00yQyovqIE9v0f3cJDM3iXGLFOQMoyO5bcUlV7bWCCreo7DSWlj9kWJ7w
CvNqYKVd3tsVR5sc2gG+ddQuusWLArCn02zgy4sbUsHI/z1yANPS51R9+qRI
2bWBv1FKu7QYzyOWcsIGZqvdXQS/mnvXyb7Yd5wzqaJArAQltlYq9CFe793H
UUbd3NZB0GkEs5NDhIVgIlUgqEBQh4kwY/cjTBUFNa8wlgPUohq5bStvXGPa
ry7391UqDAoWFahzSpxWs9Xb+E97bYhsySPpTNMT7RaZeaTFWYv3eTizeHAk
crHiQmwovIq878HbnO9otI1Q/k2zANN7JyjIunDBJAMsKZqO4bRlB65Z47eM
H1pUp6MRhFY9/F+oVG6WTlsw3j4iG3r/j+6EO6MK5EUdJJKNtSZEqIJgySxj
SpdYrVLY5YdaacQgDhKBbrKfygxHRjD3pEQBjcfnEpIiaDfB9xgm2pBbGReA
bZuhnd66N0p6Lw33wjJTPx3b2CCz/HrqEYxj6fZI3dZ2oJLFYm9JE7bdcJSc
xb1jF2mtFQQZ+N8YmIzSMaXJID3CMZWtOv8cCgODukjIMPxuMNCRk0QlVKiM
M2uOvMrpIdQq6UeZPCo2ILd5VOXUe4Hi7ea/NQsLHjZZXsCUEHVP7uxjd2sd
kPwXOKlZYdjZG8RqYVRYmYaXIgl1egSM2jZXtTrVqUc8D8NWg0jLwiAj6bOt
8uyAmLMf9rIiRm0IqHttOBEJl3WC+VCWzJJYZbG00WSfQ8IkRX31mbiOkMQt
nQisZb4LZg+0EZye80NGwgSl5DcilenGpu7zQV8V9W/46uWiCK/mzSwv1KiS
Z1qW3EbTN8EO9/U3Olt6lke8ZNpvs+Oo/PxROwJpTOTEX53jeWMY5l6BaKUy
3Mg4gVNpq70/pjoIgC/5fuynJ/l49fid+rNuTPtknnbOEuu0bir7d3TY79Nt
4ni8kj9p+rPeBypoihA58MvSiAh2CrE+Q7DjZ3G3kho1ffdULusnroRwFtPy
5da7QbOkVw/so+ejSk52jzXROBbtnuFVJ6f/quOYMivBFkYzDPz5SBHL3SCL
Z9ICy0zZ4GvvoxWIXwiJpMkdP2Ysly8q8/VIjfkbI8/KqEMeYvzgEE5yjVl+
iFEQOFU4EcYf8jt4N8wDGqVcdP2EraN95aF2h2xjHHtZUtUBji3WApEt0+f+
2r1StLAurhgPm0jk5vssBcugVnOrt0UlB5PsiEdFQJ5uw1eBbkoZBLtDy1s1
eoTOZmHHlURVo59NYdXiOH6b3mtVUSr9SEEEs9aE1SdSY3O+BSYOafIO9zXx
oZa2rWLnq4VNlpkXwvWIDS3V5amuG4cjGSE+C3uATZffzBHPkVcgq2L3LQ31
UzzgOngTTx0IH57OQsi3AsnqmQW5vB55nl+PPzaC+1yJDYb4G0LEPaq5/24C
Tpla8vqyWO70mXBHLRAxWsoU11L2tCPTWve4u5tdeAmD10wud40tkt2Kx5E3
hHYchrAuLU+WtGN0k7zC4yhfmKU5jTYldIs3REbluy0BwMUnzsTrpm/5JrHi
sXwsXm7z0PsLNWw2WOSokrbJ8ECMnkOXaG4LrqHcooLV9zp5dKDVY4HeuwDp
yqVyi/Ni+G71FGmZTCh/fNqNmjzfICzV6cRBb8xgd9LKADXr9ADzT3T3hzEB
P3GXzZzz8C3lJs95IAQS8mjQ62ndNXtebjGsF62py+QiYma+3mlLJDghj+uQ
XdPkLtcPjC8zb8GNlDKfMT/gd2M0D+znzDPDMI94Y7aP0g6IcMXc/oR7P7ib
fXkm919KQp1EI2nrdoMVjscLft7d08R/52DDoXPyY/I5QHxdiyC4ywDPTmpx
ZEGMdRoBv0ZELlD56UBOWfyq1j0rSbkbhZzKI645O5dJzd2XIQCFrnSmKdgk
MdysaFc+N1ogLBvAF2++3OBpvH6roaXO/iBAlpCvoF26ru/Pq9pYZrCTSQQ/
SXzmEJCnaXp0NT/AU7Hts+wrhYrsbnU17oMd0XLKLK+YUKLyET9IHDMA/0Pt
bMlmqTAVpu2509WoA545y8Ro+sbUC5FUaYonMCzwch0dlpiup9CaldAPbtVK
ZQpdgDhRuFi93kw7JW6VAWTszriFjzIshmJ3E8fdFSC2l5CfA9Am/zb/HG11
r6gUBAdrABhoXjIvQDpIe/INST0t8/tNL38euFFR+lT2tlfzqUJns1I7dgMs
3ddlSq4rZWPkV+dn3hy7wVIsLayhbMXZsFMTYLjBobJZDuNvdVPP6q1aVYy0
GzeWVGIhwRKviTiKrJ/WncNqcp4KEbw39m1rpWlvBKoCyxO/wmnntiDLbUM0
b7dRQ8MuhE9HEsAAztl+ez9IeUpFMLqK/RU/TfZdD5fboJQYDz+4cio58rq7
jkAm9q90P8212DimQpVedJsU53ktRLhy2L35wFYstD0GPFUEAZBMzoAUuOaH
rE4eoewg9x0GfXvNATQuTeMUnZ1Jqa52PdA7VEMCDilI7hxkvCM1cMXoz+Wn
bGM=

`pragma protect end_protected
