`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
b6AO678Yl9EUskPorRYvIxSINp4UWjiDp72SE5WYgekc56rlYS7S/2MGp5ZH4VpM
sQwsLxE/QskUUuqqQ/9AITpyJaCqtQ5KAl6m8sxmjLusWlz274pSz7tLmnatiP2o
upbBWdRrXDzN6xHkMqXhLdSAvhBhVBK7ZIyrw8BZInE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6224), data_block
ijOrq4Mry5FPa1QWIORMTJcFR6Ty0+DcLlMAs8hJ+CRIUb489YoPpZTOO+gkrc9D
pvtHzti3hjj/MzLIV3vvfDGtdnQT8hzGPfqaZRMOHuAL3PgO3h8dckKgISUxw70j
zttDG99qpyd4+k8ZNAGL8orLx4kF7Kw9gVo4wIO/0LKm4VBMwktInMqtXC2TPiVO
jyXOPdEDc4gD3QOOzG/E1Tq80L9YgaRvrVh7cPBGtdAPVpxTEUiROWQaPwuB9JVq
xpmduWDbBAcv8DdyMGc2s8dK4+QHfUIqvu3bpHafYNCPL7JWATSdPbHUaj7Baa1s
6SKcax5IN0DO1SnBLV2d6N92s9INDh+cDe+KcHVKmPSVkeuCzymmTRdTKG66868t
l4sV/Af/VfdV1ZZkjYunWtuI8+xSt60kwg8hZGp9OuAUdQpAk7ZQ6cAd7bZuliNx
Wk1HQtSdLHDA/39ILTtVt9XBWn6q33zQf3ndeXPWqgI05CTVBE+fs2Zi0QvIIgHY
v7Z+0nKqwZDZPFwiQEzJsBqUOFROUhZBTGo9I8R0PM5o7eL1FW1fTJIckncfe7+z
fEb8Cyk+4oq0EA0EuIw4XluFpcEkO9LPz2vvAZg/0tG8Eiy8Pk4z3DO3GK0EpgKg
jlSkwp5cbFqHuWywXQnivwiLsq3ydaYKe98tjc4QFp9knmLax+gQvjZczWTcYNtO
UdaqdnE5avIYrzXwhX2Kha+rFe2sMCr28oyj8Rk8CPxQgzcQ4MrTIFHxNHKt9vpK
/bhShEfBwE2CnGOinXpDRIG5qkygGyjzvVUR1LlzccsrtbO3n5PaaYsEzq3bSApP
YC/5fNuvBejqKSb7ztlQOQfAppZP1nRw+lDJLiymCylPmFgt+8goTiYufQoMoIKH
KmLSSRgWBkC/Tl1nLvq4KhbiyfSiSWMs2XqS3vUElOQioEFgllXH46EFurJntwcu
CPznuC9qPYY3Jj7EmgJx06rOJNE1DTWzjhU+4Yvakhq5JnxIEk4N3NmIOuuD2U6k
Kpua5qVCMtZWRZ+8QBX0UGo6lxtjoVwAHaiasPiV9I2upf2iVHEItN+0EtxnC5M/
ZocCbw+a5VSj8L9RoxBOh2RCipm+uk4j0PTORB70xkLfU33IRWX2rrlM+pGThVCB
r0UwxfOcPnfWWAV3778/NUUPocXsaStAbMFmEHryyDGoEV71kCQXA4rWmsa/qOGd
Pz7DNnIGtmmOhbCP0fhtTVbz2oW6xWjUjrTllr9+2nF5WBkt/0MCf9QQveh87g9H
zcDsYIUfdvsUj47GYq4+3aYzrRir5sjSyGXBDHxICGlLnQ6KASb5orOTY2oL0SuG
lRkFK7+MCMvklZHWDlSjjTwL/ly/4H+iFmpykXPfNYuQUHwSwPO2sgGyCOiCg66t
DAh+wZClnRUNCRrTx7XtnI00/YsiZkqaiCADpFXyQ2+zB/Qz3g6Y5CqAOe5UiQYT
SMJ4JM4Eoiw6fOkTjRi2pCRgllwOud85VcIs24T7NfuI8svhOh9YrKEAts0nHCZo
E3gj8xx0t4YHdHtLvJloGgR3gxfGqbPGPdIkaOIU920lpTQNABoVXmTCaiUfP+oe
O0oiLSvjRXRU+Bex8VuZv1miO7WJ1r0VLZnMC6H3EeRu175ji8kN1N+5DipSRmeP
elNbvYHmSr25KYsI5x9ihVL8s9DuHhHfcJtSjT4wJAUUma70fbwcHQLDavT9F627
rwISbvObliYl/GU+wDHkSst8clnwexZCsiPtmyLEUnAZ39wbqQhgkLWnfN3tTRX/
zwEybCGKbBcbgXAxHN8aBjG7cFJaTwfURcSjCygLQfaERpWafE86r/0cB2TLyqLi
s1tcn0tNbg1HvHskvjLMvPUKgQeqNs6uYPAJNdp/nk+zirp4KCLqy4dEchj/oKm0
aEo6vrRvheRaaeVZLZ4rEILfMeiR+CitDFvw+jUbJLNADy2CMOG23fkcqFT65b7G
rvaUDCfo/NxiQeAeMG3qNxbFpz9n0KNXU2ZfHrZvXH9JVJfuEFul2vPYqGWwm/bZ
DcU+5iTklxD6iW4ZmL4Vp9d5V0GVAunuhqePFRoY76E4Ov8qGKV7Ppq9+jroqmZH
6PoG2W18gFHR/53IEg4RRgxPbjUyw/x+8nhESJh4p+kjHhv19QJZpdWZQ+vTbeaj
sSCYKbt2EeQPFwG4RO4gbAVTNiBAfDvd3c3vyzMBQ+wNhtP9Mqpai5x8yfxH2mfV
SU8rrlXI8tOCUPw/IzeVXx8xnv1x0SsfvsMH1EkaWTs6LqszeSgKdXmmY32m74u/
4g0Z0WV6bUdvI5o9ZiPo8PoV7PJXXMGZzHA3MY/MeTcjOAcLegry45o5WahSBO0S
jD4TjFloSux9RpuZVYWHw7HL2EjYFKQ1u5+RGTH6hksaLsNQA6z5N7SyTN7ADn4I
ArixeK6NzduAsH/FeiHCRDytOTjYVrlVcwlDwiNCDfNMpWrNUNHiMtZwWR2sVaMv
cWzLRF3pWvC1Bu13Szj1ECNby9rKRfeTd9zJBMEdRiIv2fJL3gg3TKDs/ChrnoS6
gyz4RMzM9Zg5Xy3UnVrFEoa9iXNJDdpGFBn0PeNp8tst6+wV17FEX+lXWBwO9KAz
a7/wIx0fHnM/v/HvOEutBwJjPZ7ukEnRyAbkPgKChy0+GnOetYtUZlSWspN6Race
cOIh+e/qCtoG8L6Iq4dmcUEFQHr+zLDaCFwv1l2MLXR/92wvWBsw/Pjitjr23OYM
JSecub3ApplOBcTY49I+w7O7ThyN+tnJL1Uv3IctCHCzw6L/MoAO1SL7lgw4BL7t
6C2ZLBAsu7w9h7j+E3JMXpFa+jeL+/YYD85UZ+hxSKmsiUD+0c5bMjwzJB7t2UHC
4pWYKXqvobBNxFlnZxvuPdQ/o+UE73vLK2jHoOIyw5XQ6C6Du2vFauulyS/OqlYc
TU7y0SodNnQ2qWpyqYnrjd3v9W7dUZwlnTek01KsvKOP2mFcvyv/d7Kic8jljprP
T0IOZGULLYUllDrRON6GK4/HK2HBxWt3lDSRcrHj78UEqHStWstLbRlGAocpCnIm
Qaozgq7XPYj81EJ29KJDVvkUTnIxUtgOLOqabIXvUhK6jJsc25vDRhNGVsB5UFXd
RBpdqmC1bUcGlRhSs/fDDTyRmb7aClKJq/31Cl2/lyvd4+LEpHf2iHMn14nSx073
4nj5UI8MWYecAIJXVN1Jzi5CdimAxMkLT0+E5DaiQ6HDm/kuRB98Jg/8QTn7T4Je
+ETPX9X7b+hdqKmaGnhb+2SopsESgcPSX/jz88HOw/zFjWXBg41m8afCMFVB0HFn
KZ70MjP0r0tc2e+4HMQjY/k3seBviTa4dfs6GJhANVN8yK6uAJs00uB1LQSPNzVI
S4MXgZJL0lFyK1abgJkU8Jm0appdMUXx+5YN/pRUPbhCh1ucdasD5je5SoJO31Uo
AAC8r/SO8ylqMyndq2Rknf7QbSdltiVDcbVo4RICoI3il2rihH85bvaMCOuvR9ls
1btvlCNSNVuRRCZ/25eFSugY+7C0kqPnlBntD4TuCGuQAJKR6WneMXl613a68QjA
lCkRlxoBzWfgZ3Zs6nHl94QpXmbFBmCVc2WEfIwAR9aLKfAUnveIbAlj2tV0M2fB
P70i3hYxO3t/H7rwquH4fXF/mtlraMfUg3r52Zl3VjoKVMRl3ef561YENRfCHCcH
LsRQfxI5j6Yd9I1lQEu8avGlyGESbO26qG/g88Nmfo08xyeK17sRNFX9ZWeKsg5F
XygWnmUAJxKJN9IbFJIO2w4YrvGIU3XO4MMjeQ5ygyY+OBVK1zlconaeABkI3qFF
5JnARa3WKT/stTE1OfpxlJcfWg0FSfeoebtA8OctWY6XKpDGwkjBmLgenrhV6n1N
BkfglKj6qrBddYmvJdyGCHylO0fbrqCmqXrYkps3OcHiY6HceKHJyb2DxAgR6A22
LDwWrKmb/DQb4MEks+30oabCODbQCQ25ikRB4/bIPZ+SAzHJxhG01byGX+LDfZlR
vb/T/w3ogOanXXXZ6FbAO+EljhHRRPbBSG1HOAgCGPQxeyM3VIhk85NHC5/LY3n+
p9sbUtfjJEUYBKqqf2Do0JFNeLE+jK/QDIkfamsBpb82c6eWMXm/fWFo7n2+S2Bw
TsZWUpM4TjOmW6GX1NGO1aLZE7S6ld0nU7lsbAKe0t5fxOx9EBggcCCIgEkU7f97
FkRcjmcmB6Hko0FxHc8mSRlHz2AJSnSmdx12OmoJd0VH0j33ikCpt3KnJtlUTJPy
rtFIeutPGFet8XK2xPhsBR6wZNKC7lK+fqfQpPzaxXGgghwdzCsjUqqKCBbDdY+R
AeGJfX1TMzHpaGdnurBtcs9y/qrzFKPADegkNxuH+YpOyXJMTQRO7tv4Y13+i5jW
LIXYzk1NklmZpUla6Ay8mVcKrBkaVatZE2O7lxErB8YQY2AEkFGj+EreHce1dxOo
yNBYI2YH9LrjoC/wwzQUQT8XjO4g4PpTUkdviEfRxSY7BFNQTuLv9rXOPIPcnLit
MC+LwER9peZ2+EJQTj3Pxitmy0UagjwjEIAUQWuGqAdtFyNYCQ42TsUR0DlrBdUq
d7w79ijDReyPIXl1lQGsRY9jXKxGXisgyU4p6E7/HBjrVw1gMaU+HqcrV/wK4H8i
hgxwY3U9JPmKc1YCC63lwGCcRGeiolgihbaUONOC6W5v4lmbygI/DoFj+TPt77ox
aROGU2XCsUAEHvyMZDtgHbFixEznwZo4BIF6ty7655n/kMkB2311RPnHxo6WiKU5
qcty+W3vaiHZy9YYmEBNc+lAaPjKbmZZyW0uJOHXYw1GAt1KbC4zZS650BLUAHpa
f9dlTpHYIwqg+LSAxJnUS8Ye9rWyDnzRw73r1h1hnmUonMD0nrcLq494/JIpbMCM
1x3YkG6i9l50Hp0VQ1WYSX5p3zj8uVadDRbNXJB/fFzpivzMCVqUAAjv1JbHqYdo
wCUWJSnhLxjb5fLUXgpXgVNzgk/v33fJwcj/nnhiSwC6Bx0Eln3+2Oi1nDFB9kWe
6A404fm7OwPMKaSPh7ZiGVkQYzfh0d0MmepDY681IuHuNTiVrAulwf7D9/cfqTjT
+Q/C/f873D4dLPwEbHcE0eAGTHRfEV1hyLMyPo7IdmHe9xG5rDryrTPaS7EVsFZG
A7YGv8wQMXCD8zgLXmf8Ku+khazrvEI35eUQqS9bleW/q7DGHSpIaExRuY+j9Qqi
L0YdM1XaJMCmxbb55V3LuglQoWCrGify5P8y5WzGqbnQjaGK4ky2pmNOUU3HeKCY
oGD7JnN6Xo93TtCxGa+y1b95Lr8pNLeRtjVqGM+BWFkGP3cSPzCZlFBSfMjhTO0t
ylekfeclQia0uLvYDa07j87HmubifyTUQmJ2zCvXAjCeIU5zhVbOOjzrKN2yTERp
lVn4RAiqa8Ja3err84ymhbX2wFpnri5UG+RC7PZkBhJg+hnHr9eVFKUk4e1mJ7ND
iLzkWEuwTO9irtN9KlvBODv5jq8xpNPNtXSesCq5wrgj4qtRKHA1a+ZOW+LOtfmD
eP+DwW32viTmSP2VmkQi20h1FMwWjHKJMasQ+8TmAqN+ycy5sneRcs5DjxwdI6IE
QdH14Ds7gWqlEuLkSJSGhwoIsaQCCBEC8Mzi51BG6xAeIuwl0/tepulnOHxn1gQL
7QmO45sgek7NVkLQJYnQJ3Jv6kFopap8IU7yUs6PZLtupnH7Q79k/X0er/0jn/RK
qv6p8hLnPArXhQVi76x89yK2ylmqk1LE5rEsChO30/lIQD/M46oTW3CBUJenSETI
9W4zlIqAM3mMV64sFFaMQ4Rz91JOZO4AsU92mvC0BQzumwsZVNq4W0kQOHRi6jRz
TPPdMSthgEIa12lhZO8ygjN1FjYNSQRMy1mYm+ow8a1PpySaVe21cC9dASCpCF7T
CtJiGngJp9BBYKQFZIIa4lJsjLDQTNzqa8/Qd2i7f8vhCa//a6lrXD4eWNaox4DM
vkLsWXhktVvWsADC4d4Fv+lUDw+oYTI6+G576mKjdIM+rAtAbhUlb8OsCygmKI9q
VMh0jjvofHlkT7KYbNxZ5WN0ZBbFP57BsLxyXV2f3u4/wH9yrJEtql/icwbVkGZ1
UCJN/AmYK4qOqkd6/sok87hkMjxvTk4dGhlWukzLghLLBrTy3vgzgQplWeIvvClm
vfQG2RVRUUpGVfQpP6guMSMX/D1Wa5ymAzLQE9o7WWvKpXqh2j3kvokNVueGhgQ2
4LJ/emD8Xk3HgK1vSxhnNHAxn0zFJ0yPR9A1xGNQ3WIaiLG5sgofAfs6rhBDLHHr
5USv8bVCiXNLzoXnSK5Cjw+GGBWwAJoEOAoTpfVtMkVZT/ndwD2THC2ZB5gQndPr
FUH0sANMiZXueIQikLcxumW6vIdBQZlN6fn2ga/jj24h0CUYp3ltL93bZ7ZFgoST
szqT4fmxEL1jyTIjdH8V/Nz4WOeyhyDPHeIUa9Gy07bP9VLbq4K5wwYalAXnwi+8
qp2ESX12CR8sjIB45Fdw0Gj7e5EhGp7hlxqjV4yC0VGv9y+Jggej7n46N4r/z+50
DGOJMUpUcaPH7a+fdItQt2+p2jjind1b7ZwY+qlF4BuTNqjSxDS61C/8yyl8dqtO
X1+uXE11CTHKM+9Bs/usq9V7o5e/v1wUpYOc1i8kVv0hzHicVlGCLbhKHIKmKay0
Wl3PfypO3EKb8DBGfzgwIFwMVU8lHpwEwn2lP7XiLPemjGlQTkpt9vU2ZSyb90XT
a7VKKL5Rg26cwogfCyGB82QSVkDlp6A6FOenCa0/HT0Zvmk03v178yJfeV9vaYMi
FKBGODMwVUR2Ly8nM1kFLWJYpoaYkPqxgCnvObnyJzVwtIlpcBDEHiC0eEZOBy+z
aC6sNAmBxHK/HQPYQifwl1APH6HSPyq+oOOxSYva4HwF/7YQq6uB86Kue7hWJud7
IlPqoJoAQbakn9+FfzHAAIjSyLXMQesbD74uMqgBmkSCSx1AHBT97nSxn2ch2G9y
TeHTy/oWEqAxT5DUIqTaWTjgbkje5HWzNgqY7vPstWrsRdxmopjFewHhe6xcesbQ
gO6c2QkvNuYXvasB1pMWaq+79ClvF4U32XvFQGNetyCJFtYB2fWKa305JN+1vhPX
aG1U7Nktq/tmZo0RzP20+skiIFrU/OmEufVZt7luW4Tm8ab7a3HM+w/p0AGpmJZQ
tvmBnjNHjFBMyxhfHbYy2JVE8D9HZvdIQn93xO2yb2BEKxWZY/4lM1IBLJYd2CM1
0wRL2MCQm6j3bDNAEDIfiE3kyKcjpAYQvN1scjkjvxRfayCJ7xU2l3dWe/2Ee0AU
CYZVXwSm4/YYQA6HoOjqxlgiXJs1QXbnoZc1Ky17grnmGTlnuFbl4ykueKoQciq/
qRDUXmhGH3yY+U6aN7eZgO+USXD4xBpQIG1zWHGg07tZtlSFAeVaBZihkWokaCrv
A24Glmxb+kcq53upoR80C0C6HqhLNisTsuOSWkht/Z3w2fcDXbICaG+xESORxTI3
uVVv8QzfaDjltvVjlep16j0jYLa6Sj/sSvy4Vm3jPm2c6iXB8POWhbaGMrwKQMbV
a2H6vHBEorJJzN/iXVJ6W4HI43pqssncpXer/PnEKUnnn9xCgyTo1N6NjqK38gvU
7lyO9GH2mKSc4LAcvW3NiBPLSpmvKtKQhfvckKMrz4YLFE/c8Jz5B+MK1gAecFqB
Y72EsPSfF/wueLEOBXmpqYjJ9HF8uVikuS4cYtNs+eEKZQg4qGYIsrDbihIZow2v
o/HyNAuuPzqLORLm6soSc5iTIjhrddWscpA28gnbkQV8ahYZthP7kTQ8k3bxHsba
8nP8JhhuNYrQauvgnh5SdF+FPg9tHcXDLb48RuodX42jREXs2EQdAHdeSlydfaHk
X/M3CZxOccy78ccKyhMT6YKhZP7tLRGrpyLlcaRPdD3bp+ABUwx28wzF/tl3677s
CPC/Ic8hoEtNeGgditJ7aE3hBo1uGLJASRSbCOlOXso3GGpushGdTNPztEqbRbnV
qp5/0CWNtdb00DkesdGl9pImkHcJjrse2PuiA4yUDJAlf/1XeHTr9kG9GVucbILi
jNczEBP3D3/RcfCdNHW72PXQTqb4vnw8x6j96RsyQXzSI5OpViptwOtryL7C3S+O
b0jmT863WVewXCwHRc6CS5jgPVE1wzA6P3LZxC9Rsf8sR6Y1Wqqn7TXGvhd+YvSA
LoQauXXJ0eTyxTko/X1/nHKcKXB2B3xsNJpVzoHnfV4=
`pragma protect end_protected
