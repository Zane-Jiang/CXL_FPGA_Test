// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RpLxJlOXgZMJVolzCR3NGkB7tsEG4ALUXpOTxsTT6GRntXNhi4y3gGn96Jrd
WJHO+KEmvEQwrfFnSKMBQgMuaJl/CnVHKbhKtqJkH9eXejWfGawGgAwOfzHW
4KJqnNjQZIABQ5GNne7dwERdofNpO+6dxjQA6awMJTXtt8lIWXnpDyyisawI
oLYop70nb/sqX+dWtNPP08adj19lSfkk5XKZ4rXBUdOizlaOeobZAm2cdpUe
H/hrDrNXECp31jU2LIy3/iqqyfCRuRgjXMS8KUvOBEZKSWInLiF2S867gWUO
wFNrMdU3Kow5Iy16OPipjX5tZG/BK+e/Fa7upitl4g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YABhHms7zztW6Jdps4EbkoG0kEcQ9egsQF8mwM9nq748jeefPjEScmas6ZDJ
oUPReGkcAs/rZMJ/yL9+YdwY4Fd66Qz0yL4mRbuz5dvbia2Jwnog4JEVA7ry
5pWjILq5T06zBPaYajhHfWCeY+JWrqG9wnzLfYDaggP8RyjDEsRH4s8g9kKr
uaVtxINDvmNgA8Tj3deiH2rOuPiWbU4/sdCnqxTzLhweIYo3PRfWFnUoKetj
XRZyRU9pIaWuK04b/0dnAu/IyD9Z8wF8rgl9U6+7Tik6M0uunbGpUwXZ+3C4
yoOuXs4ocOe9Q826aAMzPuh1BOkA+t/zKUnCD+4STw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lk8JLNrcd2shQ1oozqWfsEkbn668v3Xwus4h/ORYPr3kEJQqmjUEzIHLG0Wp
ZMhvI9JaIrZi4iRU1xXVsotIoXao5H1ZoXaBFKL+65WcOqrFxcZEm/skbjhS
chb9d4s04tK8OWHswJU7ae3J4jGlumKeOwPrzcXWugYFOgFmwlFUK3v2KYkb
ei+Ld9HrFd+n8ggxdRyJq1IQ+s73PKc4A011Z4pEZ5vAPRPuts6crU4IY4Jn
cIQ+smzYa4oaHKXednO68RfJZ3IfpGpZIT0tO0FZCG+DcAeoubsL5/5mvayZ
QhuEaqB4C4sVqEWmeSunrBf/S12aCsVYwX47i7JuXw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mZr3AJnx9eCgIEImXCSYHkiJRi3CSHWU9Kdgk7SOf67RJ36iJSOxbf1kCK94
IyVaxX9fV8ThNLhyMhDmI48DluXfUemlohFxu9VGpB4e/n39Shzzhy3thERu
jafTDFGgwfjBpfAeYD3unF9PGfi7QRI0EWYaECNqpXIRopsXiGo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
CnwSNXv6fExsaZjKyOBTPvvRdvCpQZC5dj2yfloR+tIZOJpmO4AEQqwzpa2s
aZwUgI15t6E6k1VDUDcFxhKHdW7bHyxMK4slc91QI6P9DqSQVRlngnaL7dka
c/I247THFiwrSYgQop4ihcAjSaQ4fDj7JhdNP+PV9NucKWtOJAVp9QPvwlSO
UxtisagcgRCGKU3iCE1DSf5oAHhI5tMngTw2guY9LzLSIvfKNGoL1Ve/wKal
nxhbvLz4u15S440YlBRc5F1gq8tbftJvT6vtiDEOiTbpj9JLm9KhfgsFMDs2
je85BS2FZyCuSzpxOeSqeLosrVj0/HeDbJoIShgoDPurPyO2uyIMa4JYV4DE
MDqSEAZjdOk0fS/lIiF23i4aCO9+tsyQtiLOSZynECyIGk+Xgh9ibLt7Oecu
zGaKryhtwwaDwyAKniNGlzkxFjvukGYe9wuWeKLSRBvmE1CdbZ5HvvpoNI3U
uWki3etlj8FUEbd1y+bDNwy3TozkMel3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tTDWE/woCLfOGGYoYt5JFtsNrfCwyPs3Pdhx7ep9NedGx2DYsAgTTTYEK8dT
uI9+6w6KXA/1qMUt3APEFqBHqpg+8y6Xqd2/bCcyuAQBCd/j65hBizL0SbtR
pxjBOF4VUUNcP4JnTAKn8TbWWLOO6w0ml6FegVE443wPvluuUEU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rwI1Zb5MMcsmZIK6ieEqwc0qeQl7IRA+xykBdYfnt/8De/hMBPHzl4eYXxYD
eW/zi55oarGiJopiupfAkxWYmY/zYyFArwgTQ9xU/RS6jk1CkIt6be8TATdx
Cs858TBfWnt/Snv8XQa32qcB7YYmZmdbPY8hXh6kEp/STKXfCC4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31216)
`pragma protect data_block
IkyNBMZU84rSv+/DRFUfBUBuytQNt943Sz+0TOYLMHt0aoSM0/xnTSuw2Z97
2VutBjdlEUdId4M76z3nZUeDx6R16Dkk+durjy9vBfcU4k+HpWUNx1rdOUR3
3P+PSBfPOb+wN5HvjmG4ywxfFszXsOqtl5j3UkdN8EMspUd5K1x+VTy8HmOc
jdaNMVodX/AcMd4lZKsfv9rrzEXnX721Oyrjf5LxqgzS/A+JFa6OSw5ck/Mc
9fcwHXIpWhbLharQ5uawwebgJNEhSfe5ux1XbJR4HOcUiyafg+K1DSFRgQZr
DH0wLOQcf6oeNLbkY+g4LxFwLJeDZBNh0Ves27SpH61wobWfDxGqIRT3T5pd
ZdC7IiPp0gFuZSbrBs8DGenBTvyhVg1Ye6dRoYU5vjoVm48UyWjY/vxvGjEG
fC0acVqZmi7nAl6PkCNrGxSYc4qIhtvyMrdXSgw2kGQM8oy8gR/f6p+seGCa
CsZTOMWIyaKkSrk9Ba9+w6uNQGJyqUrCLTpoxc+fFWThexRih5gM9RZXeh4e
kuUXDJr/hJtMyQm4CF3oB2j1V3n1h58a6SZegiJPgOIlGvHFmloRiRAkH5fO
/4WrUPr47zVByy8bUMBr+fnQjsZZcpjGB7FfrvYjjl9/JhUAE3WpgIDy8d2V
fSH0Edn8++d1ELFs7RS11vzQZg75H7csqdDXnZHjl0mZaRFrgczoR70OnKe7
Sfgu8HwHcHH9ZoUiq/R4KwNx4lfLsCfsd7XvdC+UIxjNuqEMLKqoAB3ccQCv
0PcZbKXmQSEmSr1kDCTbIE7Osz9Bgpq/voNj+f5CZ+dP9VXNDKoPCbxXh2nj
rrKyy8kFH+A/zIMig6ihFy7O50VtU3rRb7E9VrmOwV9Uu6vvjHD4SJBrBgpg
SI/Icezy57ABLFJYxIf4UhzWZ+dZssBipUMd4VQlipDfkOb/ioZLHue1Re7a
3jj2w6hEZoIvuyiQsw0jat9t2Xayo6VS94NfiXUaWKYkVQPv4/RFK8nmeiLK
QydmswYGCwJfQaTuTew/Q7dSuPPKSF+13oplD3NDt9jz7f5CQF3Ud9WVgQHH
Ajh6BHLuik4QUQr//UJnDa8mEMyONNR+QVuAYszLQmls3+U8sNeC7I7fTywZ
C3sBa1pxWH9bBdS3e2vYhWkIapEyX3kIcVVjRG4SPW6ud1yIIpSOU2mENKzt
Sed+Pj8t5uMmRurn1hnYKLfL5lwmy2J26Ezg9bZxZXD7SBm98vO2sn216rIu
LUxpj5hBE+JJuPezAh1QsLl6DQSlP2cEYLp4JfygK8cuokKNMGzUIIoiH/vO
1dazte9IArZUhPw8my81bqoJn4RHYromTbGrIbhrw/e9oR9FDELC2cdsAw/G
Tyyuf1k/yBeeUK5ASiN4EnFkAvniCd8ubNGILH/Yxlz1OngGTBUH9Sma92sn
J5pAhrid18H4L+O5lwxQ/tj5VRpmGZqUWKb0CqYimAzI3lDEqiVDOxCfoKuZ
uJViR8OWBKgz4kT0zWVblWkg2fgYwQJoq8kC6h8s5kGCNk28fJp6VqPygbI1
JxaABXuuHjRl5d9QkVA7SHPdi0rSNSIRrBbGtw9qDRKUp+szbaEpEKrH9HXL
auUA+EcH7nnmlIRtlKozKKd/gf4LU6IAaWNoWCd/A/ttxTDu0KXAJ/JjQfC7
cv6sPpIb5fmrvxUTvbSwMt6k6ntYTVz4qpMwD5W/mwGCNndkMlK7Sg7IeErN
BM7iie1ZxlYfPcAiSXHnANr5QRhvd2sbm9VCmcZ/u+e4tCrKbGceJfDoj3se
aeykG25OK2QHLCj4YrSDBze5C+3OHH2vlvi/hJeZoP8TVWpbUW572K6mbKKS
VxTXwuWscKCHdV8U7Hc5YLTO3wdo7hKo7dpg/1RxnDKBcLJtjLAM4lXsUl24
spcBZAm9zbh0fCJUI1Q47MUdc81h5aMRZA4FBYjDc+MDTcmq6QXogCmxrd2P
bMyKp2o+sIeeJEWoF/rSlfQP8WJB8kLaLhR9fHFOaTbcPI8mvGuURdaKCuNo
kKivpbZasaQweWCFFF8y4KABimdl3pf8bhdPY5VZd89HcDaeQA1w2RWffeps
q7jzhabu4L5GYR7rqiU3SMkJZglfhiCWHNRV2IJa1dhJLeAkb/JKDY2Z0iEk
HOeJin2mP0dEleq1DU/p6o6+uvHvWdZpxlvop1N0/SzK8Bt9GCse1AAoBIRq
2FCkyultz3KgRU1OHQQgEPmgA2oV962YkKYrE6GjETj4YGouxcfcMl0b70vw
cAocu+yCdRzhWHc/9/c1c4ASPR7gf1jZbck1scfXjrzWqAivvIRhOagWf5jb
ztBc976wTcS/3Eyiq8YuL8VJhhHFEOY+H/+tmDOeHyFMuRCjTL9ZMgVPx3lQ
E2SuXh2Il1CafgT+5ddsdFy4LxZR/TT/hxW8Q9yivrczqhApCrM/8gFlrTJs
WX5ySJk0uuutY+zML8Xo7HiEcxn7or3Et19Dzc3qVfVNRME3vf7KqXYk/EPp
fO2JdJ9QzYwLDEHB/6AMGYj0rVVQbRRH4/YbcwFFarSk3HU8ZL70zAGdNvsY
cyUboRvyr+RfWxfoIQPUW0aInorDzRLlnqJHVz5kEza84wJdjcieWkMwmwtg
5JsruneBIYgI0gcnSHCQL7RQmroes/SJvZSMD5OAvYFtm0jY5AFA34Zz0WGi
arl9DQHIys2mSeWynqBjEqt+YMmBZ1itHBqYAax0VEFOH383e5kCKDHCcnmv
tOhOyDW3veZbaEK1Gxh0dgh/37XZ4f4if7YT82KUHwjmx5F+M/r+JU/P6byk
gURM93LoWnQbuGgljaDglbEkkCY6NzbtX7ofjXL+zJIpmXLyCG5b+UUJixVK
l61LGsYTKnwFxpAxk2w1WE+5tkJ7iIByN4IUFyGjvzMWQWpsCjaBGd5rvgwe
cbopxqAHpGGpzAUEBqzQNsmhJ1Oi8lpI/OjMULnPYEnSHqCU9t2uiC6VRgmR
jYEB3L8OyHvk/gcR1FOzub1Eurl/znNmG0ccf3WKZNmroB04TOs8HupwBugt
SH/cyt2usY0l0qhat/oQfHWRGdli9g4W5/7MykLx/TjYya4DgrartGbR6Key
78kVne6W0nZERoQFSTuUCU1jbu2YTBc9hlQQdeGIKecJbn0SPKasTkbg+FRG
wwR00EXc5xv/Y+a37dQderXIEn8c3FrCYjRlFaAJXBqK9tENShu0IXhNWbkw
8qRuMNMWOtV2G35DA2nXiF7+/wfEHUnrSDTFPZKnMlwXRg1EVRpzI3nJNIkT
QLLu9ly2+6qZ0IY1qaKbriVz2l51bKBhSLfqOLIi9QSwVDNIMNyMX+CVaiSW
Unkzq5GL0ECpuX2PsIrzhTK3HGQhfq4zMxH2BfxUwu6+ryBmLfDJMh4+WNiu
GGKTXCFEs5b1UGyPRgvb5HUTNdmjOv2VsPi5W7X4qy8qrEt0KPrGJ8rKZ6oM
n5fWCf8wMlzbhe3oqXCYK1DW+CUf6fKrgmwhT6y2ISvukBtgkxJeGPgHsLtP
fGRhMA9nQFbiVdz+Kv9wsAWTJ8AUbAZJ/Dv3ksCK+zLQUKD59mOzv+J2ntsN
H71n0IuJoE5gPYV7NkszPYm/t3CI4+4NNdWQoymVKg/TxxSvpOglZOrIEsvs
xGwi1BWW18UnKIoC413qBm1k9k15arSyRtiNLR1i02dI9LsnFOviaDK3197H
+ql8GVoByVozygpZA16/sPbc36JpRM3ehWqp1xD/fpEinku4XRg1ahriy7lK
eqHH9z59MtWytuSavwqCybaqwBGOldQzEQ+kgkMQuDIaPRg3gxBlkAE35ECz
7nnhNtBUmiqNgZXj8ECseNm9aWi4mk/jKaAR0jmodUhpthZeaZwyvnSkVK7M
Qz1tkWOKg/85FmSIuMm/5Lw/F3/Bu6cUAE67pBdQYQ8nZiyX3pS4KuX0Csgp
zb5vKighFO6uIYz0Y79I6+5/vffBX+D+fQtiLCAgz9siaqA2PahtIq1AnOrv
BZiYAej6GAfFl78zo6D2m+VYT5g38tXIGcmlXlx0BVMMApR6w2Pv45vkr9bx
Lm2ZWPB0RRuek3CJ3K+yerbKvhVJ7y5oiV2Bg+njKNAsoZZhXHR7xnBPLKDU
jIVX+ttznrlWJ3eLX54Gk0z3KsonYOt0TPnza3juvvirv8FPVMyIze4Il37e
mES6Va5lAFVwsun93vWnxcMnt+a+NJ8+aGp7IC9cAMVDP2VeGZsZuSagvNin
JJUoassZA9V1i4P/SKD3yjQQ5hktIwqAf6ClcxXyqRNVk2ptI468J8CiOEut
eUs4F7dgXx4QCsPHsgz0/856srEI6kTebJUev0dIMv2LfxilqBK/lqPTC+iK
M0QBhYg4tX7iZylN/Sc02tdIY5B5FAEp915/zuwCJqvMYnYYGT6kqfgH2nNh
EW4WSVllQcsYv03muXkoRS9P7NZEK2kcr+qI6M5YemX6flq2ATABU8ToD87K
qJkfZCOuFKRqR+nmHlN+eay43G/OXzN6nuoLcEZLn3O0NSFiuHYBJlsMw7SM
OmW0DiakXo8LxgwkgMi2dpxEwS/JHTFQeMDD+P29VI351NVD7DVG+ftjmCEK
8zlh/HIxAiFbpcoKzUk3aJJZFLiNZI8VSFvlF3281wI1pqphVJzbFLgguTk6
ZQc55FH2OeG41MTdbLeHbvFyVv+8Qbkmf0yzaNna4+zXfjBkuDt1I+gZmoOr
HShlPxiRAoVAZRIQwp5IN/GWRFjROzwZYdFg/hoj9X8e9lPzT5ow0rMDdlTn
ussq2kXLAPrea3pU6d+XT4jslIbjE98dSc7dXhuw5dP1usDxSSKqyYraEtvr
eDhoeXhXbKWv6Dbm+JDLGICVPzEgigdDVrt82ahwwAU3ENXq1B657Jlw7wLD
28O2q31FPlcK/criCCC4G2FhomoERn3McJaYU10oVfX6Aer0xNKT9bI+Q5Lr
TFzyrFlSosh9RP4Q+vlPikVCIDiaFfAXudNrR9mMQYYfdWmdNenixBHW04qT
GNBNZCNPgFI5MV7qvdGadEnu+dXYwZs3f9Un9or/3YMlqFYJN3aeVjS+W0h8
ymLoUUBlJm2S/FE+++sUxxppS4mouA9AviB7UWYURPqstJTVVsm2y7czB2re
wvfix97vwP5pBTxxu2oUk4b49Z6igJrAHSV7EC3EX8CvM9fQDgF3bhcdsQca
vU0K0Tsz0lM4K7G2UnRMSM2qsSbLjmPAr9ml7nMKJMvnlpBR0ubrwQASv510
TERslHe2/NkTeSCYiHnyYWapRxbhz1J+zyX6/mszF0YbWLDzPMohLWPwjJVw
/unu9rQq9GeWneuYfILffkNYEnTsUFIbQQWb/uQw8iI5BckdJSNgv6j3/fdG
nj2+dIsc+rBZ6Tq4UYwPaSW//yIc8U3YRyz05zFggthDaVaoTQzkMwR1toye
jcSbCVy4to4XSek5ZphMpbyNcvwhPRZva6neKf/8sd5VCfvUPRu1XySZuQBD
hCfWkvSIHWaxvadOC3O2ybxThsroPpt0XETlF8o1uKV1QOuTFQx3WnwbHRaG
wcbp0mhl/dx/SuyUdUZPBQXHXmvk9QKjedprFwKLxYB1huQeHP88F/zdo3eH
dOD4zvMLyP5n2jObPTgw11Q+WNSqx0uDllg9OWvVx3Ig/BLKzj047bPhxn+v
2+crdqCZh94xH02XMroE5OoeJfZoQBBp0+B3P6CQk3CBK6dbiMwe7YnGe5jG
qcuCEy6jq4qQbUTzt33ZVr/0H9RzoSWylyYU/c+p+9f6bWdVwpSgwuQOXjeA
8YqYANjoMXjS+pB2m0COm15F7FIAE+nraxhcrJ/d+1aDhM1hEPxA/PHtwei1
CmqfWM1UBbP1B3b5wqdRPaySAe12H90ltOvhmLe+8qvMVZp2LLlTYVQJPBpE
/o/G4f83KFaLjgzpCydAHWME4IXH49nuU8drzKg52ZJMGbnNCmLcfvBhLtf9
iFrXglEzSIph0OnFgcGXQZL3Fbn2tWxF7vPA4ncY47JmV7ascGgTpa0VL9JJ
wd6y+sskDOvCjLq5Gj0s0VfjEUxJNCForOgwqNUpxvDm69oCtQ9VgqakL9yc
oV2DNIKcbMPQFsD81MlFuJMNhHkWVo53zDkrcrC/zp45ysGbVmYjMHcYqUp/
XYw+aHAcdnuAptZG+1p4GnHfaFLeKmM3PPka164lIfTzhYXRoYCxu1LETP1Z
wBS862y4Yxu2p0ytUjF6pUyIMmUWTK8KQ0fOsjf1IjNShmZruKhr43Z+XN+o
FbDPTk49ZLDrrT3Yk7noUWWIGClDbBiLvPqz/ZLdQdKCrPGxrDhXnTjU7bMS
Rw84rxfri4XlZXJyyLIjIgVEj9yyzzniYe8g7uRXTEeZ/4HFsG4JfjmShg91
P59KbFvIokFP4zsqpAZ+1UbWishk6OTkIq9sUKTNujI3azs1ZBoct+RK46xl
92QsgoAZA2KUxLslpLW7fQO/WFJiIpOxXV+hFW/9w+FdeYLO11o4/Mas7k1d
ljC/WUgVmgHQdBZOmIvsUGnFR7XwD2L9emH47DK/SutPZe0+cxKkVomHbo96
igVCHKxpeUOjsIQKlAFaEU0sjiWj3OV2rXfDWoThiyCzsrz8uV2NXpcTQLzU
tJPfXWwiwRzbZzm048i3o0vM/MjhBzTXoRNNmhsBPayjf8/AxjDUg+6981nM
IXzxwjIgRAjzvST6C3U2K6mTLUxHuwvMejUdNIdYxUkkn4RJzH+Rn1ZdfhcT
hW91HnPqZ+wM2d9P2iRSAtLjjJRgi64XbLlCmNAHoaOsl0K5QQfD2Y7mWjBX
m1/QELwWEDyzyhRRrwe5vxRF/y6B8rcv8A/17wO9rSNrqz1SxgB35t+pKhAd
G5tdQkC90VptxhyePYkA5mirsGtKmNhLMbrByD0s6hqz8gtsyXPHfbhBUciH
iRkRkPYi/j4jPsCDThJ0Ae+0dhPM+c0sFH8bfqATZMizb4A2lIMfchzTRB2Q
oIVKiM8uFIK5/R0bgnPfuj+wYFSSfhnaPhzHGrZK+esgkHtEHsaGEdVpdhAy
HAbu/igeSAnqiTyqLoYLF7BS2sOt8vgzHy2R/vog90YT5y5ey9Iu/IIzdmFN
gIlfw+xxQavoXMk7bkqT9GG4UeQ9s54jq0nxLVEgsA91QZpvcwqXvU6U/oRp
DtgdnKv7GgBsM3XnHGobVh+Xf9FAN/8AQEXorqM1lXeE5akAnRGY/f5+JAzg
sWRKAT7XbXXldlxNCC9gIt7w6b4ayFW3br1usEVRTYsJa/yOCIG4fzcFVHCF
/xhC7ii5TxK6CP+3H+3YSOTOvt7HYL6ofVlH/d2udEHKYDFjP80nx3teCIZX
uIvTEw9Mte0m7WWqA/fx3kCqGJ7cR00DinkmyMDobNm2wLwaKMhA4H5N51fG
A88gKUJ4elHPAUHaxjbCfAU/h2BVi/eqO1gBFrctDokaVRyy4y9j0Bf5Vysq
s9MqJZcCRqGspeKeo2tnGID07cFwlttjaM1z8A2EugJRK30zDP8Uix3C3YWA
rin7iQsshnTdgKkwqa0StwoYHmitE3lRP/rBAjmIaJtsh0SsVlJ6XPelpt7S
zNBr3yh2QFK/9ciReQfGRh2yZkHZuKxqBH9YGdiVbNfU46DSyHGrjN9HhQ1l
SCBA5k88ZSLhMbjl9PmjgpHs3AukFza+OmHzoFKR7ORWuqrrGt5x+zodbXry
9nBglA9pa3RQtkShQbwIGEWrIIKV1mw45b1f00s2LnoXg6u5gjQlTvz5hOga
EiPidGk5lYFDV+8io4tSdPMmLAUiq1oItN7K825JKjwryBoO3Hl/zPZZ58fZ
X7MH6RPNQmZoL5ujtiNU+5so2guN9ixdh2H2UTfp0ccnVE6IFDKIOu85NMRp
OAGJquSaiNgnBxQrcdRiNBo5U7Uk3Jdqql0t7CpNQjib7scQQQ5kaQuNAIqN
w7CFsQKrzxY3fPLww04p8tKgxKqoKIU0nLkWlERDwos7FAjUaBysmQl4HFPh
oK0zSsKPCS8v0IYHsGKNvfDjnvLjQpcX7dpg9KVnEt5jt4RGpuk3ur73E5yZ
RFiAGKlma20yuQhIustXtW3noqg8NU6GfBYld1izUk5B38P/rU88U93F/i1J
qbDQ0YRX5SMsSdi3rNfbZ4eQbuuJDAGY6rC1Ebdz06nxvZEBMPcVf+19I2MT
gCSPgl5qfh+jDAAzGO1YVujB5LLZuMawTwoOTn0Dv+aZxkvFc/mpCg+HPH/S
ftPyq4a4EAG1eadZX5GMwlSUgOf5OiQotlCXOt1vSfM5VTI8gm3UKrZiMfCP
/CTEvjZQpy7dLl6YBj9xUV+t0I9tgoKztADz4HvDI3HvK9VDny+qi8qcBdr4
/duaMFYuKw2HZF+OiBwKpj9YOgHo+78I+qL5qWqsu2kWkk6zihRrJVbAjtwT
hoTyN+5l02crc7UNcRRHfE9DpeVrRHijcUV+h5DR2jWzi3mvojFigMwD5a1z
VyC7Z7/yp/FzwjsJS7lcwBDZ9oS4LbobAdjyss+p16Ibf8QZzcTs3hjiriPS
tGottGVc2PspI6NkwEkLbr5xcacWp8GZ9btX27e2IUeuB6+evoHo4wsX5m4I
riaiZH9ER53Qbdkh+TzI/wVjf1Nu4GecTMjj8AMxdLDL/bl7JcWx2/yXKHpH
aBzjC7MUxAKr11qBwslVRJF5vSdr7e4D34KPUFqt9KxGi5/F4wyc98Q2aVi8
ZgxLhi3gMk3G3UTOZgH8kh4th4Bpr60QQfNSswalBXi3M3xTzSndtXv7ZEWU
3B8H8Dttt6pR1Ej/6+NYCM2vTO6tgGdF1wKP2H9Up8IqIvQL05NkEjg/s7DP
iVRQirwGUehvjBwQaTeJK6LDHyKrjCmog2GsPwzysJuLepp34QRyV0GA4Xfs
PONwBMPQr/oJh3rTLD2q8q9tCC3HxhHjtgiEAyKIQptCJHISdnfetsnKPOkD
OIH2A6xzc6fSzNaaL4GMpSlUfMxxwntd0LUEtPzgCOQIu9DQSX/pFh5vWqY8
/wm+QOb+DpSyhho1/aFktLlbDcbOBntIPmm10Xebfzlv+Lt2TQuslJBleAn6
TaNkFqg9rtRkMuGq2L/zWCW+8UPYtLlIrSOB2mPQCCJMSKJ1UEvdlnFEgj/W
BoRtB8xlbZtVH/FBifn+oBP6XA+n3ib+dNaWJ5bNLipkp29xEUs/WVBoiPyM
1utDLmPyDx1mQ2d8ZdGuwoF/TsZ9ukX6khEH4x5nc7JmO7gpFjfmwE09E5Fg
ywHVZqmWHj1D1giHS6C+1cz0HTZbX1lIKktealI024IG3ftVVT8edBshou8O
W/WyJ9tvxoLo4IjfBmvvYUCv7Wf4Czq0Y0/QDN9KMJtEJy8KwZ4dyDuESLNM
uVOuulzDc6zR+t7YoSf+696fub7LwXFcBScgo2/7KbU3RUBC7jnDGWsdwp98
k1r+egCEPe3fGUlYCKQ3XQ7VgFqQsQC3wOe7jA3jeB9NzDx9tTalEoPpDTyv
uJyZX5fJXDH1kDARBcRvYYaO/acUD9KBHv9JP7RA19fLTvItsc73MGQvJu0c
In7u7gAcq3BdHbnMr36TUUme/zKA6CsJwuBizHJ3jFE9OyUnS1HpQGWf0AsK
9DUirbEYva4i6wo+fudnd5LAeanGMtysf1sEZtXneg1LCr4Ac26EQqwKbD/5
2UTUIV2YHFnRWnX2mIX79xpn/wYDC/PSmb9mOWrde40yOhzo99dVY2veuHRZ
Fi8zgmK7gC56ix+M3mzEUNu95GxKOy8dOqH7BAP51wAsAK1G6J2Uei+EKFZv
Nk6b4kTlsphNg42DtNK5xxlm1oMlhbaecpNu6+/S/8YNN3+/6Oa8cWq5BZvU
VoHB+7fXpcJ2D8XxUh67dDsADv0T+hAzgs+UverHJ4RddJ9/bxK08zF8NZ7L
3IkbYw/cJwjOJoIlD9GAQUJktAgVhOCyzl5ynYnYMt3k6T4y/NIQ01lEnEok
wW0RC6pAjwsZDaUg4AgkrjFxG0GLesL9P8vh1HF4oPGYxGMhz+uBLqdC7K14
EfXReKGC+7LOEhxzDxci54klBae3zeAwQD2SZDV/PKBkOnXCyrBaEbAZM4fw
LWVclefgO0UZz6/xNCms5fTaZxjecytanmnig4NG6svc2OmR+I7NEQm4p7sI
af9ozeuGgR1e6WZp/eoTF6uTbc8dOzF74u+DTrbsbc21BvGjsCaBlUkds997
VgoHOPDj9uyNZLVVcKI5frEwjtEiWF/6XOaD27PTuDgDmCb6YkSHnxfkGnHh
XDCHradRP2okEioQn34sW+44LdDGJq/55DdLhI7Mjm2n1xulp7ZMsvlkUj47
YEkaMSFdAsdB1vBI5G65/OF0xXX8xD8Jn1mKyoEXwxjRcLDDJHBCSn6uLiky
ycDh5Cv8Yofb/YbWFT1PkbgzTQLs7lyvzBFlg+K1lKfr7IrHeRTvN8nE0VL5
XzY+FBk5nkwyssRVPx1pUG9F8Ht9nULKURG+NuolGVTkplpxwKslCYaxS9Pq
/6ZQISV5EkcRso3HnC1xpmC7Sgs38gaxWGraOcUwsas9qrjdi8Q2QOB9VIgl
NlOyXwMlAEs7hv7pF8v/hEG9RavFP0/as/dFoReCe6XJydUmrFROqwyRg7N0
Iop/oY8NcWfQBzw72AQg0o+jbpVlIM+PT/JQywkqSYMLtyHzUJPEk/kXfAZ+
9CNx/88z3QtingUYCpm6+Vu3pu6TTsffp0ieoLlixX/lii+Bt4XilOemhEPe
lWIy83EX9L/wpIToST6MYRYIJD5ZSdORNwcCWquADiC5uL+9cOuwpVjYPhCN
qJoKfrLESl+is+Tm0rNVsY4NgcMrzxFG8o30jOzVG5QwzYKBPT3VNgU6FiEn
lE1ADesiJfK6hJX+uinN24309D7B10LtQx7DRqUqeCqhpMZQfbm8KK+9PXU1
2/jL2+SPlmi5jjN5n8aJuEIGPGTZTX3HMZYTO/Zg5DLTHVv8BvdJir6vfiH8
Ij1OOm4jwuct6mZdn+uBfCwGfBklLZCdP9j5ii+jxxfdFTE+Jo/wowhslmtP
Qx+dKJabnttamUAJegqb7vEhd4wjwp7Bg4SulJlhO7GFUWLLqI7GGNYCZE0I
Dvt4oZT1OUr2f1qGCfB8lgal/Fs8Vw98QZ/7mMsZpxhAdN9BNhWAhRivGcwY
sopPQGzEN3X3dfKGC17An9jq3RXvYIaktqJh3iOeEVQPUDgGf1HbfSLQ9L2B
y1GqwvCUl87kEVQDCQccL4vkT97jDCvtlo+iTzfrOoNt+zZwZq8VsRMTDswb
DgfOTZZhTrargdWylVBArDG/hEDbGRxepyKH832BoVV12QLF0EUNkr3oAuFo
nuZ+aOWsdhjSjeeKHl3lhcx1qvzIeOjHTDiXQG9W0gr8N0dG8eCAeF/7lWIT
AuzosM794sK23Ef4+7XMwBGXWFmnk7fmHAFXnl2SkX4SufjaTHkUbyA/LuUU
sH8jZQTqgeveHU06eKQE9DcEZ2tniD2CFvM1rlrvj0mD8DSEKn8zVUTqcKGZ
EsGrTevNgkLmG7Hae53Q37bp6w4mspsOtvnVY+z4EcYyFFxfJxBVQBYdi43F
Ykt2aX4pE2leztpGUwpL0OvgIQmdJu5ZAeeRYUnnbDsqouvUrYKGrQymsgze
ngn9dHBSydGUKF88zNjWgOuDpLb8PAuQSp2m/U03xgMDjsWbT66UgToUzXZM
F+goYW1q3ExGckBQzbvjtayOFo3o/TEzFkXJAZIkAPIxI6vNm2z7wsbL+Lrr
YWVNq62RtLDlFiW38ASh/YoXmqKkzyaU/JMOzRTechRTs2rHZRLQPxqZZki8
OV0mPZyJGCWwjFZcD4LugOudv7/KYyjaAkyipjFh3sXUcHfhd8kR45szfYgV
vANwzJhVPcZbY/01nEaquKvkMM0o7Yw+SWKZlUVWXzO1IRAUnoganow0A9jZ
5F19fJ4u7NYhgQ7lSdrnQHVGeZlrjP5fniKoAYu2yGJiHq09jKpspDgNXMvZ
koDbSuoLVd+zPNvVRe+G9FrYryufageNgOKkMfo+K/mv2Z3Zyz6lGFNrK0+1
CEZDX5/E19vQQ56fGKbnA5Df5TA4LWDIAR/RmTl28YLaFaZadtyCu9kIQqur
RHE5zD4XH5LW58DIEUHbnsU8TYFepOsET0sDwYQ84Y8M2eN5wFjzSziNH9TK
1rE0Owhc0/4kvSzGS8dEBTQFjnMNARGLgw54mBY69ZqMq9BGh+FyY99ehT+9
tcuJpO1UrzNBd3NDEwLmUmYCrLuRhsssLFVjobXsNLvVDei9ErwfOyX3Lsh6
1gjW8eSQ77xOz906XgZ/PZLlUkRT6oDNikcipAZb821w1GeGonGO4mrgzR7R
MIZehpbUc636YdYAa9y5HwGH9tOpwnCiCYt1Hb2V/9aCoEj34KGCtqy6Sfgh
eDrrSjr3X3fHF+pB1U3rnJCxGujZEKVLpqOJMJpgZTlq4S6hfat+jeYOKpGp
/5kU48G3jmigAXQ+3DOB/VV29ewb4doSfaH4LTvKJfibQWbSsnrlKBQXl5eU
Mcbyeh6/zlAO2WJD/w65tnyEz3grIMyofWe78117xLSHRYYaQ28fshFCRDD7
MSsijSjD6Jh41GJtG3D3gFEoAkaqkcw21BKzAkSxhrKYKuIjAOjCIp5RJTIo
l1ckfjWdoaqwJhuUbSp6O6pBCHJWOvz3VwaiS0ZJIA8hHS2aNbqFGFFV1C7O
nxzZjk36WDuMe8+JoLFin0usyOsSWCxs3xqPE4s8AsXFPebgyB7ZnDK/yBva
QnRq6pGV06hzXEjBz2HpaHrweJkV59RZDa0O2B4GEMsK7WUXb4aVMMEcIXCA
tVqvACAoCcYRQHavAQabxyUgqchJg8jtWW82NwRRDFUTWqz3cEN9f3LRA4KT
bV95K7mr0flCnk0Fz7e8MZCQLj0yfajLWm97PT0wT5kuD+qMQXVC5gP10tYJ
0E2L9hFHIkEUdYQNb49LGQEbU5wUvDoXKhjSuZlqkJs6m7hKgpXxCho//CF+
sJYO1Nga02qhyox2YI979+OGwvxgtfX5D05P6YmpThhsbDcnB6ZFDR5hBezW
sETWEnX/2f4qTDAaeWMXXnXhkcvtuUdtQ0M6I3mMJ2ooYHoswczH+Nyx9XX/
3mB1ojIYJbuDrhXGKmH69elbQECj0KyHbeG2YWw+jz/ZJynm7wc3M4eglP5X
/0Lndj6VA3vE70ENoZU9nIo3EGRAhDDWu7+Tpi6XimsfhlravC+11G4TKowB
4xnY/nuuR1k7tR90nh6DVZmTgp6uYKEhOBYQRIs43haHMQv8xzuqM/gp4Nqc
LL2DPeSTGY+VVckLflpcL3BH4nCtmls0CyRXKX1vlkzcf5lU8LK2Pz9gMsBo
PVIrgaYFTFOyrLIum9LbyzvLi0UPlcdq7FOKGcNgzhVBMWB9nN/6EVFqAM+0
x+CRjq+M5lwp4oqyRJRoe5QsWOQmO7mLgoOyy1Aun84rZhTF/6I3NPsxCSUr
MJ0mvC9Cfl4Hs+y8vjjcLZXl2iXu1uvMTN6MiU8mr8pV/5AjlbvBoG/UlIkC
ZJvl9ksLir/+lFALHN7R5i2GawN9rUzmunwiKO85BHXYxHuQ19ZB/QRVVJTf
mDWcWEdaf0OI9iYw1ac90A+Fp7/1lQKq4vaBsJj91IqLyNG81/vEUBcV9B8Z
eqGWhjnL8QWmvdZaYokfO+Ip9+OF2cSb3opceC9zlpurvtxyfw3PrfGallxK
wDMBDTq2/8YHFCLvrGYwLzbZaM+l8Uo7dHnW5axvSSd5BjAMr5DOQ3MGwFPv
dj+ZcLZRHSkBbKxluzMG8PWUPsPEJOJztsD9Awv5ettnrn+oxTU4NZL96fXp
T2RdVe77nB0dma2Aunmlgpc8VVkoWk6DEPLONKgWdIbCYuiEP1Jn1WzOkZNV
ROxWWw2vu8vfhjM7hYIuwopIwSu8oZsiXL8GKqAnhFkIlU55O2loT9ZBS9f7
Zi5rpWnZRzWv+5hrZHDOukakXj4F+Qk4/1F35+vMG+wNLfq95/Rn16ntA0mJ
QnCRtdL/9WNe5z6KZDFX80rnp72Q9XevVwnKnfw8aUV//1OLmDfWNJ+bY+Hx
Q01adATbjoRGMNgRT41FL9iWAM2AemiwAw7Lp2r+NY9IrMW8D4aB8MWMlMVd
vr9E6frMnUbIxycOl5r0sSXyG5rGc9xL4lZKQYpV6WoWCq0bKGWjXf9HvtB3
jxuZ2OynJ3TJ7cFTEi40lTA1EOlOVauSYme/zWtaMMDj3w3G4skqPSDEFTEm
uz7kySuEdZTyjxPhQ8jMM3n+1F5n4z3+CqvZStaEHCg2v7Tj6Z15aim4xw9w
+q1vj+dsK1RAJRTIpugIqBDpODpbmpf2xNRvYSlhnHay7vb9ZO+51aLcBdNX
6WSeYmOr5ClO3EUontD+FBQxwr3ognbgOXpwSB0ceN5mpSspq2SHY6uXpK/L
/Y8ow5SJi9CpaWtJlZ+P5Hd+CdD3wZEcRAJtSflEn6OtkhKiOQnHMR7r16ru
V10whwCUnHSYySPCKrqqf5tei9Jh6xD665f8G8wTaFJmIaV1ckt54LRdXdQq
nwqVQLYckgzuJpqHuHmISx5d+fYksQPR4rcMEmv7fWLXd/tt3kJCmcnDD0M0
+tnjN64/H/alTtLTlAs9bOrWgR/Oi+TEoh8xRisXN00qmq/XhW4nAvyvLxk4
97Wp0iYBr7BiXt/G9++6DyTt18UUcwPEszbqm43Qo23mK7pSjhawnomkwglH
cBxvpBOecvcrOREbNuN7Ddtu/cJaJKS/cBBQELKH41RW2XRtKVPtVYL8iFmF
tGAeLlBWxMrhC0P4Sovx5ghM2ML0baLSnGXsYvumX9Us+6zCeQn4F8/pSSUo
WezHY+UFr9t1CTbHKOt+/BMoUYIGayO2sKBs2f3XaHnDcmhO33EZyjm1b9Sf
PmAXKCv9CBazIC0HuPxg8QX8McePtl3L/RksXqbHduV0OPIAtHxA5apbVFVn
/zDxb79GI81K+LT0mOXsJS0RwSyzOzDr9Nw1tIvxvS1zm6UEPslqofmHnZNx
4BCBuAHvUWpbNI5u1o1gyOG/68d7AAIXyS0qf/GsriIG2V8TlwW1819X4igO
BiApfgtPUrV9rfKZh9njVRvGVePCJmPhCpdVK9gImVX1YqChkPiKdayuZo/y
8BvAAFLY21jfl3o8jlsRtKcHzmkDfBx7AZ+cFk1UUh6fwF455PKjLcder2hF
8tGI9l6enl3ErcpcHjNTfpRTWnRZh+6CMUvjamcw+17OTP0F6E39pEwvFfXT
kitBr5Gn+JGaSM+IPz9mrIaFLEPWi3C/zZwlc1E+vBWnisBXJyagbgPR4Srj
zdOAsgy5cT7UwcRX73lfb3x3wlvOMaiRiDDtMFi1oGmJhyasKPBPzpxgAi0f
hBK/f5mgcUCBQM8uXtFAGZiBz03GSGcqU5CZ5RHUei5HIZ8Xyc8G/yPuvHkq
UN9xMYE+jZgpENf7+aq/3H3KnrHDYLGDmlZsjpduh0yT83B9BTze0vHTSQsD
ryRAb8qPnN2mjt2h+e5dgK+uYOTXc5tfU1TOF9roY4URVPfkE0QLgI+1d/FG
moLVkGOIITFrLfO6zNmd4rAdJXv5fgpQ841Ek9+GhQgZ/f5bx/Gk2etUOhHS
gCHYtYRbJr1Fw7NruWBNzXpBRVMano1gYMUSIobPPIEw+qEDfOu8yCEslOfQ
E52JcyEoTEpC3iCTkGK8JcypngohwnMPBmxg9yosXSY54D4BeQTLVwjMPstJ
qy10Rx6jlcMGfHgt69QAQHoCx63tZSulCywlMYRQxLdBZmVAMOTnx4A5SHgH
yRBVAVjTS+lXEwTGN7GJl/WOf6leuYOgjpMYZ4BdvofzElD08uU6N9UyFOkr
UlWabpUP3ifUXx9veCVkvNJe3qO1sV47SUXnlUTOUR3Aef9dgKxTHasPPb/9
D2mVwP53hwESeD7sy5IZgg5myyAv5LWzOnOXPWVmTVmCmgGXXM6GAzK3OP06
80c3xufGXpXGWJTRypaHWhlUHhKn3qq4anTSFEHZY3yU8Uo0pHzdxf+XiDG5
5C5gyJ7m/5rxKIyygVXz0594SIM0BTFpO6bwDYB0WchY+5Qw9P4VoEaNYOj2
EhUdNv59rr1f/GO4Ov2TmP424hB+jl0OLB4lWHZS4zNCT9ArqYq756lLGZm3
jqJuIDeZ4//xb5Yq8PiawvWQ+QN1Dlvf4hV5oCn3OSySZpHvnnGTLc4VUsZf
n6Fvb9ISlPJY9JhMlPsG6wTHgGaNx2NHi4hZpELYKQ2b8/+dVY3wC4C4IPdh
Pz9ZItv53fW0B2pHHm5E39hdpgCnVA4OPW/er9OthBxaCvXEJXO3/fh5N0/b
ANZzLUCaTprH0zvZNTTR9GAwg46etKT0Unh6AYvI8AjkSmJuKi6QUrU1SrAz
a/a8pCZhzVPLdiEDsn+OOMjQ0xCu5V3Agcslox6us5x6Uve97DS1EftyLHU8
3+SvytMQcHnecDKqlo89HAojTA/UzqDi/DiuKF1h9w1fGXNJW9X8RvVL+hIF
KSkSrPqJ+hYQonTaq267Tg+GA6RrdNTGJn7FTHn+Cse3KMeMblge7TOWuLDN
fVnW9jbnaGzUqsY99KQ3PJHGKBwsOSUNagvjOkAe/IQh9nxIJG18qQ+/dq3P
1IxO8LPQSCSp4cCEDuMEQdvSS95cef+JIbOJ4wrT8T3jLUl+FOM9oCM14mzz
41qJzflRdTZ2EkAmzemZry0M5zWu9MyFKWs6JnnLYjNC6jfx+agOjVuh9qlZ
c4KkOel8t4dJYF99XAWyAC26HqBJCWvPj4aFpKeHGbXdp9T4xahHid5HW6Er
hz+G+qOGUgAp25GoR0bjuAL1keUo3N42AevBWM+wzBoPrGl8v824anFg5jaT
Cs+b+YgedugG8zeBexU1NVg8YMmA/OTVdfSq5IfsgAM5kK6hTqug/Yx+Gq+G
ddLKfBPHUjX95OFsnCAc2nHFDdczXMsaJcwXsS7hO9lqT8byTFxxsxFxeK1k
Vx+/DB7wvMsc6zOHg6bEnX52pRxoxOhWFp1uz9wCyma63er+yqDiY2IZlh78
e22GwF8yxe3g2XuKtfCtyBl0K/yA0m+jehflDO3Yq9aCbHMk+9+hRsFL7YtL
BsNQdWSJt/WLtuX7qrZG/Giq8uBwGgsbM1ltLxxAupnNM88uy0JrKr6nfYex
hgd2CbTSZYvuyHdv0w08YR7V36FnuAypkg/A9Gl66h6+1sDvTkiMZnTDPOyF
BEX8wRJ0CxTz7iHQfasjdeYvbesucUJ7EWvQvd0H7xpD3+bY56v3VpBHk+oK
3QlCLpo57nEdg3xwcMaH17EKJUBmnncR1AjicZhV+rIHW2cee4hEQiQqxAGJ
XC+nDTxe6lDIV0SCK3NWRdKvwaS4I9srYVU4FXTG7blAsJ6j+3tvg/wQ/Jbs
8Puq+0lCBlXbJHtAHtE/IIXzT7reaxGFta000yzTvBaogyFHVaQURCB+BR+U
Ziuug1ZwmU6K6tgEqtSt2HJRxAfcSLO0mUp7Kuz7XaCFxzjPGYmeUowVxB8s
hY2GEXvNwe9TFv6J/uL69kfNARBX4zb3P39AFsEWEMFzRCX+EuInJntxgMLg
AJcu2xGkSzKTd9uYusoNUWxKvrznTNPFyLTx+/U8dpxwJuyU3ph1q0dNERzG
vdniGRnStrrxYgi+15ts02WIz0xxTddAf7T1YULMlJeXc2+aB65Y8p3Tw2Sw
7Et+Q50eojdnRY9w99/tED7/BeCsbs2Wvt9EtNhYHNmmZnPjQEHbE5ImtXq8
NwniUNl5AH3SsNPjusj2FPSzZienMUK2Kk5224shOb8d6lPG1qW/1H991s4p
Er01YwmhvOHf/RKtTDhDpg5MBISpLlz0pYBYb0cFnRYkpuXqaVRIhr4SXigJ
DC8W7WsWxzQ4MIoI9rFAeAc9TQROq48d8F5i4li/uQ8On+pAWS1cy39ky2jr
4uoKj0mJSM0TmaWPOaPLK5+wZS0+veNyDJNY7vZ5NzasiJNBzD4bFxNNCpBs
7tRzrldRkTXIWMK1ua0uRfebyiL6zC34dLCwrRoe8ZXLHFOkYqx/MVAkIy+p
m7sPVp1GotQmDDlhvNdMexDcCbJqg9yMo+YmCqTQUGmj6DyFJ4iQbYDXOwYh
4sEotLwzL0zjS9DMrmO4ZncYnQShEscf/X9OGaWx/1eMfr2BDHDVQLvrKX/Z
6XV3UGrpx8TMbb6GkFEZsIdBUcVHMcunmUK3rjYa2LSrHOFp4czBy2r9y9ZI
CjjoYRgjjiyr7fMPIMPTg1+LgcDEij6+s3Bpi4l4gd0/8oslQ6161IQHaohc
HrAP4NZaDI67GJZjjwVatsl7445EDbDyQ/GNx48lKwZ7RYaVkxC4whnH8Qqc
LxOaI6/b6unP6L7ca2dlJuODokkCeYZ74ZHSIq4cfkJ2X+t6SGJTngqWu2Yb
EnO4VCX9ifhGEOxVo2QVtT7j8/0qt7oAEjCDPQRh9PsTBLVVL4UQb+t/vkDz
dMqO0e0R76agfMBrfzvAyLJ4+5gYj32gAYi8IxWzQrNCt0Me6DDAM/dgMMZp
aEBEt7ehesaXKcsxdniWXAzMO7V85Tk30M5h/y5zNi8FoniyrHdLkwldI4VD
tJ2CMxvHIkZFXjV6po/omZACugI1rxXWUF9Lxzj84dMNkspcajUXXGcKjbYe
p6bluxaOAMBqOE5OIo+PbiijTgiC5UQkLm29W2Zls9YxJ7N3VDIex5iOEVQ9
RSkfU4lLiBOmMRqeLRJk+URvB2L5BC4Bgmv7d2dGf4GJIV2YTsfZDsSXxI3f
kG2oXY5z9FCAsIZ2SncTb1WwMm51/XuL7m8fJzoUVnN6iisO7leMf8bmJ3bL
tuo4Ix4G+cGeXp/sbb3dsRigGfQRYpYK1hYDHj3pDulLROixxdUXB4gc1zzD
WZiFuF6dasMH5XLX49bU86csF39/n3hZW2kYLTjZ12/TXVL3pI0lVPeI4Srj
U2ME408pUbbHooZYBpLKqq5WS2Cin9riu0wkwnPXF761ENQ3EXj+1Mh/FGpC
SC6JD7tV+qG0XvHkLQDSNdkMulbFbVacpdbo0rYMehL4ZfpcLbp5wX3gCu1G
cF/6pE20PoOqAsSpimHE6sHO+SXjJddwUUix6hF9v4hqFNBWoM3V5Snq6dgd
uIee9DWe+6Jeodp7eHkeOb6qdt7jeX62wcs//SdRM4/fg2zk6XXsGvYSDfH8
Vur8h5GM9VD1MFR9ZsXHFxiNdXBdGU3cIKZ7SRcLhAyX3xIHdnXBGw7bbtP+
v6eHXld2OIIeqeUcwj174CikDctPoyX0w8/tnnvIUqEMUgoTA77LYgxgQQ8c
/bKuafR32Mc3DPtUpn7BfPH86v2LR9dJTElCGknNuSXwOfyDb+uqIdAxrcYk
uHusnHVRza6PmwljMwLwQf967oXNq8EOJQwNi1mW88oFzaii9+/CEZZ+CVlq
eQYVX3tTVIUNeq/gdNyktCKVjHAxFUkY0hyYU+4fGEnVoPZGEZWbaHiK/D8M
XsWHO0N0af+rvPRr1ftOz2W4NCRL4H0OiR0ha8y82aNvNYuaiNikp9/akD9b
bvtaBpdYlhARwrJbzlxY/6a/qKvs1rey06mL4zbi3LypTxMh5TC7PzqPcZbW
dp4NoN4aI4z4i0zvuN8HdtyZBQGHHdGGSFgT+M5sYatakp//WOwFPsee83VA
UgA8amvjKb1RBIU82YeoieHoA9NrEWi/dBEbx3ikOBlmKDieaqcMiXozg40Z
s0iZHo5IrI8as9afHbF5lz8DXWYsbshtq79ILwYtO9IEsahTNyomVekmUHIj
RBzQa/hMWgLzyUF4Tc0F7PJ2gJtS/h1qb52KgeIQFT8VZYpi5CFPq/kEbIEn
q0iP6fCXu4tiWYsAc9s6QtsJoR1a+f1lt5wNOCD1b1QWaUofNeczUqqdbiSJ
2S8wBWZAOw4S9nOPqvec+OfNj/EvVfMIWcXbEtSmwapcUpRQSMnjI2hi/UL0
2LS0vrhKDZcHJgz+ZSvLNdKT+zQ7o80tBrRLkiYwfXyfvSlNl2zBafUHNXIA
In7GgGTeQ6xQOnZt0mlFEvpALDjRBpVDjlmwzroB6jqcYA4gC89ibRrH8JOH
rchAs3DyyQa6svdC9i4E9+aZLLlhpusR42E0I7NGyJpSNTPKwKVLzQocrcKp
FNATTpo8c6NNuYHkmwDPfBmzUqYk4KgkJnbPqi7BUBGWAM6MXKmEf5O7zkU1
oOvz+V3+yAjR52a5ESgXn3l+q/7W6RBtaEEfJmqOqFHVOw4FtX5DiSzbIeln
BbiSQKfakcOOpEHeZayLXemFXOeEBHhWd4/x0UWC/9kYwKWTkFooRWQgnjDD
Y9ERk+DAVYjsnTLfmQfPNlBLAqDj0KS72TyQBK0oQl2YyusVmR2SG3FPvLvj
zRzZzBFVLFiyrp+JlbrBRkywIVfQVv+9jNDEesg9aRuIa+7EGS0/OK7bj9Yr
eEyan4gFGrb3gH+ShAykSLTE+IddGmaa1khyPNVI99jvvEUDgMgT1gtGWlgn
0XJHv74n4Q25Z0fbVKkY3OsgKiZkejgDQtpd/cN659Zutkbgf1RLwyF+ZJFY
SbkTrmU/gY0L2u/9DgaR/KsYvtsQBQ84MkGVvCdlUXXHptLtpuDdXuYgOuCx
u+qjNjdSkAfuQKyQyKD6WPALdVZbsqkJZpUsUNfUEinKagIF4/U/G3C8Zp6w
3nteD9Z9bto5yCZIDX5DVW6JXrySmNHYYFiYVFt6/ShQ4/QfgG0XBVRfT0jA
WpnxbfO2unRmU0+kh5oeUFzVlwRuVo/ohUbxELdUpooCdV1TQH07AJMjJwLf
cAuETAolEpk7UvUAKCFm4rEzLW/NrsVEbJ7nYISCl8hC0BAyzWHAnZBzmVCS
I5lYy4U7Z0aHLr37Gz4Q/iu7Q9pzCFbMkoADbGS9HaFB9e/dXXSiBfvvMqVe
JQpoHjl2//LbKwtw+kKlKw/XRf7lME2RU3v78+jrAhrCrp5mDd5E/FMH86Jr
sQkCPoMjaLkOkzST0e9ZDKlDnpxEUqOmC/Y7/p1jJ8rbNu3FKQDAH9C8KOVM
8oMV1l8qM2BoRRzkFrNS0R27a+7XapgsB4wTSE0CGFwK8mQgeiOb9Kzwa88y
fn1xQjEqMS/30Wd0KkODVL486NiZTiKEBA9SIBL0OtPswvAghYPtCabw+vz/
BCTKZY9STinmIRo3G6S/qOOzOHDn8om4Nx3UxL3askbhxUe++O8kygC2cyXi
eXBP0TScSWRhn3eGHIFHxJd/87oZvxRiF21BwWlHEvRZfYGiG4Kk2MfoOhTn
J4cg4/LoIWEcDEnKZG2u/TPbgXL/DOOG72r4CYMteIg1HfrtH5ZsG7ukf1ai
6AnzHCyZvzRdbmlqiSgBewkV/DZXTXu+cEX7RtYOHRDhI7dK6nIswr1feVbQ
mF1uJEtlxUjGbaSMgKn137sMXKC16iW+JonGbIfG/dZPp12Him0BI7IqjCBK
HEyyie7n0aMaXQnk0p3QVjNxqQCXhw/QHVY1T4K2ciaWe0/c/Vk17CqflguG
LGDlZf55qC/yVyZORDusGD38rZQ4q5K0Va0t1mRh+HdB8a6sEtFluYONKGjK
IQEKkNanFKT+5sidzWhesGV5sTfDl7I47Ej4buirrMCWNjIr/Pqkic0Pnxi7
3WpP5BC2jPKpqFHO8lJJAxPFnXd86Tl/lWt9Ji+jCWoz8nmVTHWKFPu3kQKq
hCLoGSzHjG1tZIIfdCLPNu/t4ab2KpRv4PszcjjEGFdB7VEexqoOby8UreHM
6+FJN/CytkYD8FN2tbUHxgWzqbtr89IQ539n9os6mGyG7OE1Nd7Uf8g8T1GQ
mbt15SLPzgvgZsDiRiI/3Hc6PdUP/y/L3Z2igES63TtAHSDh5EZ6ajLCvY9c
VOv2+W6tZslpqm2dQROudvGM38hjYswqBkzybkw8xiBpBQRp/BSKWV3WI9jI
04IZegqorRSBT0gasjalj6kudAQVDLvG1JqBJBDQ6oRr8Peqy3Oauh0PGkmh
LFeIf5psBSeUQVnaCDVZbxu6si7YoX2aY8JNrrJ9jD3Lhslwz8o4cjk1zJVp
/RF+bEBLnN+l4gbiOyRoL7He/zf8Qej5kLC8P2unxHCJfJfAPsvMX8dVecB5
0rB7vGq+2Aaa7q8jJKsrTmmbc97zQ/sWb4z5OqQ5kbPF2jGMX1X7v3bBQnzC
CRrnNxVuIezCL6KNlhTXG0jzNn9wZU6TfdVlMVyxdT3s01YomMGHiiFr8KJT
Xp4+6smdJOMKye7jp1F8d7dXtxLzr8lDHb+x3BASdhTeqqUkTpNQbbtzoNRp
r1MoiZJ4sn2ywdhpDKoAnZHMPTuO1ggQDyKj1dmQOHJgpF3wWC20C6cCN7L6
0LeP1ZGsVAnD1U//9RwZKnlxvkWZuAWFjkF6ZKVXkpiXEt3QByOxMqXPzTQ/
vq1lqVQHve0Tg/agC05Q+eoEI5SL36hjVExgnBPQd/Ss06I/IC7+tJwvtAh9
1uWLR0sQZkxxPQ/1HsXWnYsi8NkSgK8hHfAanAc3lj2QAMgTE3rS/46Cqca3
b/axdNhmvUwt6ChdY34h09AU2gS17cv93Mu9coe2yORb4tRObbVFxXUauH2M
xmONbUlEv3LpPIEEQZI8GzE60LW/Fq75oth+6u8GKWoLyRdmlMEPcZuuEKhm
gjaPioJcA9OoP5e2LuHWzN0Rd2II+0IbKEq8dZiIu+U7EeXxi7+N5CoxtGEz
q0MpErN8rtYqjh0iI7YeQoLAct+SVFcvT81rKrp/WKke56dO225aEGT6NSDT
vbMOJDBs+h5KiNaqGOcjN0L6CsrSag/e8CArQ0+YepEUbDrBMbOErLVADDWl
KzOlQiWAAWrWFK2B/Nn0AnzK+w8WRIiNuTKgHtJA3cRs1Iv088Qo6qdZWkot
22CErKugFQrdgDDHjZkZ7xfjxlV53cS5Mcr0SGPQ5EOrU8/gybMEQLhQhIGF
m4GApZOQTDL00mgkMvcnaNV8QzuKssRWZpFFQ2DHfDFwy4Hd/uyjcOfHaX6I
Aj/ROI0U409PFghQ2FcGW6AYf1l+z1Qal0pOKnQb+UFS4la+W8dI3LvEusOI
VrbXRkUQ61lGlEBtVNUSqom1We1Silh5QTkj4iUcYj++eCeaLHoKFiHHcDfT
HGvnSwpR1YPj3FL4DCDSdbcawsk0VL5G3+qxBted3GGEdeWCckYcT0u3sv0G
jBCdb9WjEhdddQFuiSB2OUiUwW8czL+oE+GEEG+wmPz4i4KV5qRgY2mTQ3sL
igmna8vd9ABruRfAxZhKDp2IpU0GuaaYBvtKOFw2jP+vTXy7N5v3pPEi/4zZ
m0Iesa9lJOCDeJAVpTbm/gWoDmh1Tk0q9GAwH01iYbZOUMzTBSQtitEdo7J7
jD3cOASFarjMEl/YU1NC/KpwJeyHP7g1aMXNlt3x6gyn/XMKtuj+iw7ztMH/
1Gd/KUNQEvctDFtWR0ZYHNrbMYpY5Kb8PrERjRbnvSpvlZWLcbEryT/9yc5m
RcmtqhRfBFXAM1g7TYKQ67UlkoTJ/MscyOS0rBQ5nKQcE+Kqe15nU+lwltGq
3o28/55tE87GvuCHjotgxtl0LIBYpbt4NE3xf70CyC6A/AdPO44J3YhJKkwH
ZPSxsOVPjsdX+L4fiW7AyBaGugOPlN26/J3/3lwxH/7tUcKj6Iw5Ug6fUIC/
QG/ifLwRB5qQhRpq9OzcBeLadqRcnn/aI69RKn1sGzz5jQtTStKXy9EgI0OU
VB4Vb67qRR29zedXjpFltgULcAjzkW8I4eqjYouabfx+/2oYvYNzaLenLQUe
Gxj8eDh2AkGqkrqH0ddDSO3fWoz039j53eL5YCv3EO0yAeYr5JLlkBWQeJkO
K4c+dpCCHKOCdFGeGWQkEnKmYOseJaOOp37QEayWGXv7j3HFZQ9c/cJ9NROk
zZ3LrhysdIkNmgxkLIrCmChpKNqcFThkg2mDUrySVbPQbuSxmAIg4OYhrZ6O
QmSKU218yKr5ObSRMC7wfvbelAH1uNUu0Vi5xZKhfUKPS9l2Q/2P/nUOf4rj
AVQ6fQwqR3GMz1iohkU289eXRQ85HDcWvbjkhaDjisUWjfk6sUrYlMUGmYMl
4hV3eEjcjya4f7wIvOiAt5cxbC3RpVahmHN1a7mQf2YbRAbclp0wv3suRqda
pgGrgZ2mt7SB2n+S5VRMq+ybsed2PbuihoD4ElR4IB2g7zP4/qGroTQzKjIz
Y/mEyi8LzP7gLG3SHubq5AkEbalj6S5ZXBHkQKQO6avWvDPvQwBcR5nYORZ9
YhhUSANxkMRAcdug1BIkm+pXO1mzx/A9OHXgOXHQDPVKA69dP6meqfyBV5wP
x2joLlrqC+iTluBwc5qyGRO9rFB5xcGw2993lL5rl4WzeXWxftEE6B6OgbJP
YemAuoBHgDPGiLIB/eQD9qnuhWuis3j8kqh6k54EITXIk6dUq8gAOBroijED
Fq6huZ4vBi5AHX172PGSnOzXzIFqsOehbs7TBrY66bVwOVDr9YL27REJ/yta
HOHdVndmExeqBppNdiNLpMCVm4UCOpx0wYUAE+wRxnq6yfn7wL5dhVSK53G/
pRhqLf2nrl7SeyexkPaOkAiw8y91EiptY3C1At7lBgkojGygQaPyjVD08ng5
ZWExDKiaA5l1wU8KiBtgXripDoCnh7iHFR/meYhT3zlX1c3Q2KJAFLDL/vPB
xIhfu+DNtYEm64i+qta9qlHDE+0lsLpQMOtI+caiLzidoLILKISwmWyeat0N
3hHYYfGJDPxNzxihRorYpQG3kYIHSaBaOLGOuahHsfHFHOO6qoKHKBvCkYcT
GEMhVhwN2EcLpiq3XY6DQAi9Uuh+GTF6LSPQjetl3zbjFl5ORZ5laUAXjwqw
Xyg5iv/OLQYxfu4IjoACMtiCLa63hzECNU7LO7GV45cystqC+63tOE7oFXy+
2i9YNTosGhHHxl3grcJ+Nn2/BLhZGqOVvGTs515BcUbFZPYe004omE+ORnuN
KA3bo9CsYYUVGHTFBMJDjPW75g//5KiOjfwAgcJwVii+yrYxkpuDujDXe9dv
vhRacCxB4YjaD5v7RZbB13AkVYLxeucSPHr4eA5KkgRtV+sfIndmQEtQKbEy
ehvVDfc8ZANsdUYsDhi2rU0g5/on4pMYY5dgWRl/F9Z4rsG5WvFVfkwEX3BN
I1/ukFKzlJllCbp51euP/m1RvyvOODxK2yctqojz0PwwlJsMJzbuYTFSxP1Y
nN/N4Ig75rgoUOfuihar9fb1jd9+6l2QPVC7NiBHO6WN9FvDrCMBEdNjCXSJ
v6BU0S2ZgmaP1lNehvUGvKSkvp+oZvP90tOAeouHsH5PmwYGsu3oDnazMoQc
vfQPdtNhDtz/nbdRfSX7x9LDBMUSvphUXQIVdi6eJ/Qr5RL8875CotGPsTyR
FIidVmJ131nWOvF4CBEnj3LeNAOqxdqoB56xQvq6wgqG1Fr1S+TC5iUXREIs
lwUCHXErZGV0Uxb7USiIdj7WluEXI5BsDxOBdsx+TMXXp0Zn0+Xu9/tL8ryz
Fy60+PF9/JOj3og0lvX9R91C3KF3PKpOok4O2RsQ3F3ye7qOzciZrJlR5BCV
y313IOhQcr4RAeOCye8hUBtl4Hu+vboOWABB6hn6a5SNWAulBO+uLtDPqWhG
uVGrtZN0G6Ihm6jlaDfsrBMI45Z/rvdTJF5faUCL6P//wDScPNpz4RlhRiwM
3KpB80EFxEbuucVDLe3fJkcPSKjVxvqn9dDpCAe/SRRQMUbOjuF8EtmRbipM
TS5XraqcH6cAVfzOFbSXECQzxWrljloDsDY4HRgeuhL88ls6r0gjFrt+MBzO
Bkzrr5ZWo4VYTcnhLFihDnau2noCLBs7I5IuhdUePw8dZGdaJtb6sZXlffg3
GpiTELonDmThS2UdSM/SNiDRvBJKrsYX7w+82OogL508XIzqClaHMi2wJUnl
cRCt2QjD102q7xWskEZsmaBnm85v2EdFZAN1vhGt+bzHQmGsvuxgZqIh4gVa
XXEqGmi9OrfYbV55n2EdT64vnPATmaBDD9Rtrdwye1mYebLiRsIDl20HThLA
7Jfc93ghveRhntmzfgbO0apFqBqadadCLX39XNwBsFQ2duxQgoEAZzbJYOs2
2jzJsFvCQ7p4oyiwksTQmzZdepTwIkjiTWzbQO2lyKUG96XM94com2Q64Nqq
wHcLSlUZb/4yreB91H1JbbvMk4O7u+ZMmivZW/XdJBziE3UdoWpvLutRymMW
MOnT3x3J957Q9QnWyJRPHt96F4uQfRWw4rhagdH5QfjttKaWb5tgBDojsj8S
LyC8PBtirDTcgUjIv9DPoWNPMZKPA+WoZ/97r86Sz3yot3iJqf8/pa24ynDP
bEH82KbkYvlbF1yHRdqxfnMnYmuugwbS7rCVLTNDr4BWjfSU/GtiUR29uxvK
59IijQn0KYmbebstyD+Ad5yhJvFRuI6sv3zhthRIvehS5A6d/5IRPltChdlY
gDchp0iVt/3HBFbFTOOZp4D4dTMzl30XmrKKX8AkZdRYUxldJJ+ITOvfcExJ
xORXjcgYo4eM9G6/i4AXh2NZ2xGxvvrDf5OVIFyF8mLEO3m+sB7hU56w0/cT
riB61UXx6VzVeR5f/qGS+MZwy1LPyfG0ZdX3rNCgSYwXPUSzoQl1Q0KOfOVX
73HwZo5xBdLtvZ6b9AHAnHIS6D7y5bv6aRwAsdIhUk0m2VPxOEcPH5uLp2bh
mrWxbcdlEOd9QQozX4YFRp+GWd5zXkfhPkeCaDJEPeyO8d5cEuGAvYAxTALS
uZoCXI97M+03evrBgukVNe4e0tTrlZmIeMHKSzn1ug4L7LGywk+wvQwWsZRX
a0YUgi0iLr0VUwK8KJGkOnTJKsGwJvQK7G8oaxhcfTH/OqD8bHnHcRRcHs/L
X687gBYUvUfXDGd8detL6DxnPGD80OptA541In3KfsBeB1Pp2dpLlEQ8afJl
XSfinGH558ladwfB3lmfeFAsPrXg1hC6Oq0RudRXRHhhkSCBsm1lmDW8+VYR
mH9WFF8uKuJjRUKyMMCmdyQao2vEJFPkFPC/FlvYFC2B4ggOgU6aEYxQZmJ2
S8YM/eSKh3YUvKaGo0pHSthMWYbVSlY/fLtHUlhyjyNI6pybO0yAfqVbWkZ1
cy6GJd1a1owa/LGuO0a8rXNRWehEGs1IxHHmh5Q5GDqYcvbZnNTw/REAqVPk
/L/tClnmjQ3MyKLVOkEAnmLNcsRV4w0grJeBCIg5F4NeSpw+AlqUgf6A3MA1
hTigpWP207NPEGLxSa+yTaiNtyvyTbmewLHhgoDSMACWPm61xJkpktljx6zO
NaVriD9C2Yq30ien6anN3aHBsOPqG8T18PeQEL5mmAwhFlcZxigG/zB38mEX
xA+IBkLlZKhEBJ2R08QywpFydU8DtSyxtJMvPLD+5vaVBydAjtHwBdbcTUQO
ZBILUr1s6FgQkvUxTgO3W3L2ERnBFu2t4mQM0BDW+kIEaLOyHixYD7g9/4+p
QnuEmdPJ3MTa7ilFFqhpjgDlz7VLWp0eLO1EIYTFSPcahjmYRxGN9sovkI70
wxeJbt+hQf/XVOerZL0hmQKBCrCR4GOadPFLzmMJ5DhjgXnX144NwqLIESip
4RsglV7BDvI4ieCOU3Wxhrw8EJS1PAfMsaHaLq9Ev69xGWBxsgpl0OfAcJnZ
lmfNQ4jxCh3/jwBSJgQtm9EyhtJ+1OxFk5+qdpp15I9mBAGj7XMnE7XFXbGi
rLMyPSgREmBDam+3woSty8+brI+5NMbpB+0Z+7X2xsQ3YEPXspAEpoz4TPuy
8KO+GAFixAw/USQt95Qxbv85hsk1tyfO0Ueqduo7p6sG3cMuqI3jHr1OOsuI
Sj21bfrktdKqlD5+4z5LRJ+txxJrx9pqATR67MmpPuQd7LdomtOT5LUPpP4R
Bd8UceK/okL0UGg4lbPxjW0X3BGfdhD4zQ2G+t16Oc4gZX7WWzefp1REvCNK
SdhrvsSeojmhQYnatcu0z5UrRrJEnSQ5twk51HVtl/DCM1QP0r8qW0OlwN0q
2L/UhCJTTchH7YCz32MPhw/3Al3WFgqLryc4lgv+RhjMbQmeO+3U0gZLJedJ
CwF3N9IVHbCOp9qUuCXcrEVFO0LRBB0QZsup3ne9m0XFNLGeuWNYzgn7uERQ
Z41L/KreQrt7gP3pkPVvw6sw8RMkl2YWsxwC2zlybqPfx8A5MoZ5Xzt0tIaC
0m6m4dqnTzsdpHvRlO8Xyqdl/+PLzBCCTFBlmlPMJf7MGga7/mmTCZ4f9RmW
p2Xez37dgD8zQw0VOKlTG1jUTCqgYXf3pzKAblGY/TGWWzEiSw4OHAzqB3iS
sH/0+XqNUy0JCgkR+FpdrZy01Z7Y/N/3zD7quGmKH8hFO6P0O6wp5tfKsRzG
vSqR13VamgrIUJSZeMV4Yoo1NTPIQFZMrSZ1qSx/tkDwci/0Qx8lgJaMntrY
FBOl7bpdoW1xb/jvzgH3amz6+HSCAjhssqd+RyBhLFrt1+mTPio6/dUl8hJX
wm8aUjflyUrykZmXIzFnsap9BiV/WPEjU9N5f60OBaCfR3nZ3xrXwaTgYVqZ
n+teJ60+f6ACYvfwHiUbtc/vebT8sgff1XVzvgCW+KW0d4hoFVKDUDBAx4QL
RdoSJ1/RppBqYo46HoirRtjieUiilSBWLucaymhIpw9Vqbv44OZGwpdMFL8r
UpucG3pYE2WcTzpT9P5L1JUnaMP7KMYMpN2xaeKFeXWg2rmyeIze5V8hF0n+
Eudw4RCf66aW0fH974gzGXaYPl4/8SCwXYj1XB0L+gfY/twiiR+Zde0vX4p0
u8C3D7PAoBu5CNcifC+ggxsUjBNBCGkNwfrqc1exiZRy49Hj+dD4mIAXjz37
3qU8nNbCkL9kk4ukW2tIyI0xTq5u0n2JoQ/hbim0vaHqe3Lg0Z9FNjnlYkIO
nj7piml5CMrkxLueZNCvyKsCsT+uG3pn2FCOc6a2h6AXluO5MPRTrWXPDcAO
2rp/ombMRTRLKV87++I1VQKoRTpX95HPFycnLcAQm0XhmUb0PGl5+2Oijpwh
bJ+NAilx10dHAGaORLCyR8MlOT5iU7nvmTfo7FgUIJ4KsPUXY9O0xdnYAx89
sXZYg8d57QdrTukqiDckkHWs4RrO1RUaRNXm0Jz2EvcQa0cGEunJ+li/u6vt
hw3ciAOiTLAZ8rpLgKat0k0v9I/zIzLm5PBERCk1sQIKnIyHIhJW5dA7C7sf
2viPkAIKZQz+khwvJFwL8+h+GHHAtCCQO2xzqqDKwbbHz4i0V3p2alPOjujv
83VxhIKtejuta4hUxu7LvJoHGbS4FODDuf6+EOHdCmVoQIlFYvg314CKm/XP
Kr27wQYm4KTv5RKsA4bLCPKamS1WyFPfO0B+QOFBCLBlY6se3pb2tqSGCLdt
QLbVFCRVq1j44mbK6S1ujKKHnjJPlOEH/VaZkJMRwn3giuL19o2GP4wSxSX3
vpXdL3IqB9j2w1ibpPzTypT3nMD5fKDPhn8btxkPItg7T7Nb1xwW/PEuVwTa
/tLl5zcZ8JmaBJ9jQZRUd69e5sQaSUjy9HlIVRHmNcwFa1gt0bUhF9x/c1zY
L7xGDBM9+FH/LONZoIfxK0q4+mxQNgaPv9Qg0gHFEArQB713xEs7dKpcOzYa
sJ8EqxHPxRMjS0z2+MWWjuBREuEGrIjm48EwCxDTXqgMcX1CKdSST5Hrz8Z+
oR/0Bx2g5+/+yYMWQruVzbc4jg58mjiqs6zMWZb6pARHvg4oE40b9Q2ZyGNB
NtJH1GlgLmSSCfiqnCCXausqudNBVIVxCCgoJ8J0xmuavqHCcAYZkS2J6XtL
qcMBZzQB8W8eyymm2UhvLl4BFQJRR6QxTnZW6wWaq1WgIsOGDwYnl+JRU/P4
HR6gtYXu1iq5e7SVZpQDcWceCw5BdYHoYihc+xooiX5b1LjWhDL/pEEIr85d
iGsXOzWYpkHqIbfqQsQq3zj/5h8WsYIhxmvjYo3eD9wWDsdC77LyMWFjKOgh
ClB2mEvWIQ5Hq6uQmjOkv2b5B4etclTwwHUglJw+vDOT7YuaBjb6f1ECtM64
ekEnANzorjNbT0FIPHIhsOrXMCBPEAbWEIwGAyy/5SX4LyZIaN4HdTLYFcd9
uqS4iafX7s1oWIOTTOAwBpkKO8jbp9MZ1R9L3Q6hw5d9BOkVMXLTQPYGGZHu
L/YFuHfY3NyVOOFylbX6QVteUoi9tBHkFaEA26r54sgHtvZq0RUiUM489JB0
4RbmCr6MQyup+qaQbwuAj2aKkwQVB6mGlRKCeZrxfrIpUJt4ci9BrNWBmicT
R6Pl1nCSDrdNkk9JlxC6teAGb2npJt2pk4APmdAoUxVBgNCyIwmwGDpkAMFT
R3x9/a4Fm2T9coXy/0Em4a98OO1NGnwqSW5J+v+/geV9mUPHn+srcsinICsQ
zFDzt9xS2MQyJ3E1xsvRjrxV3pyJsJBjIwzTMFf1+bEvebfVfymxeBJoEFcc
xeHgdP8APbIwtpsEfCqfyHQzP34wmoZ0NBEeGTwkv/QaPG1HlJ4Cwcoi9tS2
ARgnfpJpeSnNJYylwdocVUCnnRD1kaeMChDaRRWa4/1OcC1E5jzJJC0ugRec
UC10fSrc4Vti3FllIlkP1mPnbYj/yooSlhqIpKE6U8iG+AJHUu3hnudNqcYN
ty+35C3id/Gv9aQLuxfcjg9pJIY77LqKrVMpS6VTWi1GZVYHbkbz5J2BYuEg
WI59HhftuX1j42QnrT9JC0rmVt6Dmz7nPd/DdyNEeh1MJw3OJw0QkM3711mF
1FbS7+YLBc1H73+Lxyu8emsKrL2nxqgXsq4zUU4Wa6aMrp5y+ilgEdMIoCB6
NFZCTtvNuvb4rMCIWcDWCDlMk4iMUTR0CQB4klG5WzeglXI7unOnN3FvKGzW
mOlAgETeIrzebDowHfZcaxusk9dMhOsLOtgLCWa9xplk9VbjP6t6q92BDpGk
CItDxYVN8jK6QUMbk3BdsA67775yQShbAxfgJwNUaBMciDuSE7HN7YEwxlIt
QpDKz/8FYNGrCf4aupfOe2TI99G7QbZ7VKli8EyCMgG1uSPIHWW1btgxZeqE
wiVn4oW/Gyn+DfrHvh9QMKcm+DKxN0HwfVtt6BBMAF9e21nXz9KUa2R6K9g/
WsVQff61mU+Lhpy61bmyVf00dUR0ETu7XF5FbrBaO9o4pcD5c92jUdN0kqpd
6KohkjaTYVlYZeufzRn9ubvTe75MvXGm9oa9wq/9+bvh/N5BgWVD9/mTH8y9
2Ir9Zs+wcL8k3AnosgrjDQnQ2SpTMwTd//DkgNqDgVKmOFWZySLevIIQS2oc
3nH9yym84vLpU8xbROJ6ytxQaF1CrKCXnjsatmoLCmYz+pdLEbuYusDl5Jiw
mlZNS3eqRze2h4tVEjBtjkP2LMt5mBhIwn9VmoLXsjIm9fWKQB5HKdqCU6Ez
pF6pnvU/XnY1T1MEho5qzfw4tcYyyZnRvEButpMKQAgdBt++pwVqxBkSVKS9
iGRZ6LUJDDI1A78tGpoy2D5+7FxET/vX5nuLi3wEzEmyrkE3HmjTJKL5dpQ/
6220fAAtwfzF3sZvWkjFvkIiUe/U0lemp2zM6EF3POjX1V4Hp2CilW0O2uQS
neoGmAylnUY5Mfon+0+z4xA+lwZB1ezng1G4S57Of/R5zhE3gBlu7Xt0AGH+
TBsvsh+humTBY8+jhH1DA8Q9pUvHzjWP2MYmQgzIEzyjj+y2L/m/Gs1umk47
8uoxAKUFm39BzOdCjfnMTeUTyq/RdjjkVtFk/m1S9b7Hw2H4zqrOEArG98+g
7O1Rso/NmOyUnyEukhfDveY4cnDG7h9XDykUm6VNYNyZnfbt4f4n1x7hWT2e
6b2xzdQtVzEsGva1AEgkvsqzo0C0gDd/wFM74F2ELWL6Mh1SHfO43wdRbwHd
1CXw6sWgtR1D9DLr8EsbJt+27ytj0M4szZpIDpggXgdsl7S6qslmVi36BnkW
KqpN5/0iOah+djhKBpe8QPxbGQwn8DixDeNjL8GK0GwMMiCObLg6UhT2xVp4
fbqmwaUMrurqdyinyyZTkdcihpmpQcbUSRzijcxYP8QmMDiaZdyYhlg4aW7C
mNJ4FRs4kzfiI6o3lQQlv38YXmuWZIfG/1af7rLQU+7MMWmGeJFWQZbhNVqo
KJmMmWb1gIX1sUremqZDs4RXkBFSs3aeTLmi3/bzSorCAkeEfyV4DRnunjBs
ro+i3mGqiw+qtIkJPaUlGBkt7JHnHRnv/0JeyT4pDCmTMeSq4Zjj9+P6Jl/R
zEX0boc4h3/1W4YOR0qiEgAPZTWkgrdQLfL52WBsyVwAvANiTHcowVz0g5aW
1xxhCzsax4oKk5zI4Gvb02+GxZCmLiWcWhDLKYpoLQtfD4CCcmQ2Ai7PUMvx
ae7Rz4fGGmzcC0EL9MgJSDxcIb4bINMNMAXJ8vDRfM2z1+dh4ypcNFTR3Ago
7ujSz5e37G3+Hn5xv2bgKHTIm5j+hFSnRpDlEyXYEqNVbOUuCpFO1PbJLAJn
chjgiOKfA7j+7yFSI2xg1tMioKBrvzwoAfjB5aGfqVilqZMaeygiUCfLx/Ph
3uVWdNysBvI2ndgGYJn0z6T4hfGkvjNrwuAa1KNZ7PfcB+pjhWT1AFg6axxA
0IAmIyg8YdfjrzG4BHGy2NaSwHf23ZL1u02wysVdryJZOSEXu8vBa74pyySU
a+7PUVyOCgEAJ6io4sHzq3gxkA2b1pmHsK6xjlHxS/IgdtjqAfaZYYTEK5gn
uZOhDX7UF6k+8o1abJodauvWJOmyY8FETJIOH6D974MJ1zK1hA4zn0NrGvbb
DWD7+AtxDh8V0dg20CNPXWPB9bWYpNGrREoVQmh6dMZp5PcLLmmE2TU8Do0O
+QIdLSoZynrmaq5JAVn/AU5+r3zfk/DrczGUDgUkLAyPMTRsnMMeZuu9TQmC
bJZ1rs3PYL5ujlS7gayXGYqtglCuEtdanoJYTRLgVgFhR/+zMBxdemxs0K+z
hkxTxMj3mgf32n8qX02/1WEY1XGZ35TxZp0USr6MBw4Bo6GcWD8vSqwp7Fj/
OpZdhXKnS0i/1QNZ7x9+mwYMrFcDiqA1NYW126WORC0itENQ7ohbOkSSt4KU
v/Yqka5eNm4/HG5wssN4EYTMPgOzW/FzQs1Lsn6sEE3fMLNhUikgpzfib7p8
4uajIYTuwEQLvt6Mz5jC6wOZy3s7gJe2QAo8o8k1h5EyJCKoVSn8RpZNor8W
8hJ/vvsBXXeL5PDy+RndYWNk9rKfNc7Xz96UsOvwpqf+4PJ89vxj0qAcmjkM
mG/ATxP/wwaEkLo7N8cVbykwY9y41So4p/XYjiodGY9oyFUxkmhk9qATfyWA
fpYxN21D52nMaitY6KFkBTSTrAk30rU3c6nXNS4Q1AMFwPJfMMBOynW1teko
Z0gJbFY6QBi0GmoH4ZdhDKVwdEycKnL1kRxxGEQT78jS1TRp1AtfXDqai2+n
BMeN8nNjs3oQccOQI7OazmaRIVFgYN+Korv/Q1zBbTN9egLWlNyYYogUJ1iB
9sE3hHwmoh43nM2/fwdyCyKjcCMTLbN+9RHTk1bwvciste5QEQ0w60hqRVxl
wgw6JEehQwWIXJNS4AaxuxB/zb413UGWV3ZY9433Zq3QoSfX4g2LKVYUIW0I
L0YEpJhTm6G8OjewUylfKby8LxuetVZF1BMDYMh5IHfUyNx5dfAyuKvxan95
rE9MQWjih2mP9miGnHX1goSMrTIMQbe8JP/zUBME4rfnPy8/uKERF/jFwfC5
lJXCluHuylLVXbe8vqjaddm50VSPCWxHq0Da3aBiunQkjA+2G7Zmth+qd+iD
VTF7w6Hbh4W5SYnkzvAC+7xNTqG6auTJ5gb86hPmrIW/J0D6R1KNCO3U3jTG
2O15ik5YDqE80BOa529oHlT/yKqstnW1VCeB3WI2AA+WgDOfNzN77pV6LJ2Q
PIWfCUZBvkqOuCTBJh7uDy6Ha9RusUYH8xSMGNGLqJpr0yX7Z+rMTkOlNHeE
/+e2aB/4frF2njtjZukgUfzzOI1AVSMtPqQLgRRdS7UjjBoLtjX9q4wuhnzw
JoSRjXBGb5R41VwBqgxYDP9OiG6e6Pt2Js3V/HyTg6YnXFGI5UTNBmoP1LBv
DgcPNoTMSC0LBZXi1b6r5TYqAAFXY1mCvocL83BOhl3gQQp/Yh9l/kgSlRCV
jaSdUtH70qAXYsxs5hT9NDW6pFtCLDCKAn/YNU5Ym5DZhI8vaCEIDTtI280D
CJOhWxLhQMXauJiR6PfltM2GSPgDr3JhzwlT3QB7roEf2V6vylpjGKxycvG7
lrcko6CtElbUZddc4OnSdTTcNoMWeENvWCw6a/U2gjpCnNG4Sz3zSul+ft8Y
mZEtfmFPeElHHoenMAhzrdcym6c0E7gspHcfp2qO/gSI4CI7ydkS32IXbLUD
FTr982WkJql8rFlbo6v1sL1Grrxj7yz5E15DW1cA5c8aHgLOM87Kj7r3AfkX
aYFu94gsjiQenUAA+Lc5XSUrgZiRVwZ9dGZKrAHwonP1rvUKD5tWtu+SI3dK
1xs0vDk2r2TtP0cWvBba+Oem5lLSh0CDshN6n2hu5zCetAaYJxuy3D80OXZJ
cXhKygkbnkMWQzKZ7RK54ep/a7ZNfJzyK9HO1uvlagPfGuLBu7cy0OkV5gw6
lPX6jzv3kcX24XxTCkirsKaUtCwP147qnH1FVmPF5YrcCbwoMXatmXbumuKM
dH2mhrbq5HsLpVlbIt9HuB9fkOq3MqyzNTfJY5fgaxbrHhR7OHIdb0U0+QsB
odY1n3S40cVf1BRNiDNiVYw8XsTyPGOgzbyOw7wIs9GaW3tEsVK0fg8AsK5X
1nXYqr0/L06o5gTY6k/Y0jnZU0TylcQcqhreynkkEFS8ReJO9tyHkWbcefZk
VEqVuKmEAPOXN8v3bRPj0UCHpeZ88UtWBxJcWX+AXbmNpTrnOJnwO3IkxcD7
jUV856pNF3RPSVyCFFpzwMk5WeDpcPKo3uXIVI2b2m0hZPkoY6kym5NKgxgj
zTUKK9X6Tyg8+ofp+cXvjuMIVCi0ce1e0cIZEI4IG0W7cHoYNpeLVQrM39Jf
wZtcja+SrKXP/83vs4s3eOCTJiMf3KEvxvY74ea3JJJDeYKjP426frEiwGav
lpXvNtDMPDYZVJuV2aaF0F7nkPw5Kstpx091ugrPlLYSMFSMxdJOzhmcGzKf
KnQsRS3hzGXnz+Tm/uwYHzTI3mOSzapkeAP2exqOSJnhhSd8uCTEh/kkkEGx
7tv90ufCsa/+KjcdVtUVsq4w7fzm666zu97pZ73yDzJZyyRZ64gb4nMnCxfy
ClkTkUef3z48BexmHQoPsJHzhsCu4nO+XFLRQGxFPthyg8QQoT7ZWGkabVlv
yg/VbAE1h7hlaJjsP0LOfPGlxDs4Bre2xiXpIhC1DJ58Jl2Uid2mWPXNtU65
bzIGU5cHy+d/dkXcal8zM/WCRVh93ppDRBjTFWIn8RhNdM1ldyKWQQdHJCeR
+HcHGC9gWRYaJqDvmAtKmiyMPKVFNSagLtdCIsWp57ym37UVuZrSqs153Gen
5177elYQgAi/RzKCWMpZ8iIAACeJaUTpF1AHlbyhnrocQZ880cfwvqtwlGpu
Uun9Knlo0ifP3bXeucFikXgvYZPZCPXEVbjp2XtgpoAeqhqqVgj2enBpP6LR
Kh5GZjmgrUFldDQvijY5UufdzSr+Em/WGGgdSm8uxsaUAKEjGy1Uu3MaxtWU
GVMF14gf28qipm3zwBbT/oyqL8mB1DZKyG91JT+odyER3+yk8V1FOVSN5MdY
0/d1RA7uYZ9O24ZWMV2MRZ6xlMK3domQuct4+3BicLmmQ+eAAVXVPCNxF4MC
Fp4wewtUctMYDEUwjY8dXkOsgOww6anMN2ygWjdeBHQyQpxXJfz6JEHYwlWl
gXax4RZzeiq6vEhvDuxL09FukkqqV5uLZIuhuvPjP7vgKdy8jYieVzFkyXLw
LjySOsOyLym2MQXS4sQuh+kpws9FHgCq9Kh0pyIF+Zu+NUdDBk3tBN0WdvNs
Ee/LLF7eMdQMPHA4v5HzXFFLC6WbfVESib+ATYq9z85VMHYUvge9SMvN/XfE
2a/eqrR4/7X4zMPBaje5W8kxo1hJG1hj7XDZg1Bckz78X2tl/e/zsctbKOHI
06JOAxjhy+5WYnHdZAoLO62ypp4RvkLyr8wD0DMgojAWLOXJnfMPaCk1ODEE
7gIYEzIKMgfl1kPrUzyKJDVrnf7jEq44RK3zi11gu7xVjjbZNbbf/RGvXQl6
P4+prCrWBpVMBhh+GMWOFSohBPE1nxisO24QjAMhUBPKk0iT4YOl6Nibe8+j
ai9kv0f6zcXAk59H5AhPGRtaT3+NaUaA2+MWZvx4j0xoqZ2EBGkd1bDTpvXF
uwZrZkmuO0si1hFWNsGjRCbGfuoCd689LIe9hpUlC4GLD9PUAKTRvZgAzhBQ
5zBrkePxZ3I2sVDP79mviUaUwABrgHkhJ/sB3HAKQsgSyf5/xVlONbjjeBf5
sEE62Twf3c3GkKJv/s4FpkDuhHvF+w5Bxi1XL7uNYbqJB+rYiEFLzX2YrRMF
sraOGrCjVD5V4ci/2VDM6TgbQc8UjpAe+Uj0dwNqKBTKC7scjTlsbpnT8wtf
0U/ZWeypKQWryUPjSx9+stzLhdnrA5aC8OxcwtBKSY4YuDc/jLKP9Bh4s652
gYiYcr/CMSatY1NBXlAV/6gMsB5PS+owhU1meXlb0ar0GoNqTgu8TMdQ6eqV
DXqrSAAdhFQ2/RlrJqJ2uUUUkhsxLeT/C4TM5pUcLPeI/UbXAyxx12bdxZCC
bPEpbaCLssdth3SDtVsW7YbYEZy4PYwr0EXaDCwvliuU5E2WnVojDbKLca6p
DINkQn0HiHCmC2E4ZgtPg66mvQl2s4K2nYc9XdMHuek4BrDTdtI1EhO0crLC
Ghj22ULcXRI+ZNNFbECk/8QTdIyRn3/sY+1OWq1mURS2OsObkMf1iCE8VfaO
RiNqpkA9oawVW3J7/hs7p09wgDd5JQlsYnZz8iPiyaa8LvTNvsYrBFd8Bx3s
Un+GVmtXkiZ/gHQ8iSU3hday6mFN7yDhgoOjM9NiNJL1aG+KFYrmcF42rZfS
SC8ETLk30TmAac91xL5F2t5IoC/fYHanSZP+mx+QoTgZjE1HWHp/weXIZ+g6
sKf7mRpdIGuH4nQLuhsgA7ujzc5/4yiTOzcbm4NNlYcasKKMsEg3TqY/roJe
2FgXFmUDTxPPRrwrNIsrsX380Yzh2RCdSQGggz8OVghAQxOKia6Vm36f4xms
6oMOVP+OQ5LPoWqJVIY4HVOJrgMSXT7NjQ+KFuaZi+XQhNqWpgXBmlT4fMZt
KrEP9sK+XegaH+1Q5CxZU29Zqev8/JGKCj4ZQXt+1FDkk5WzFqr7yEuhX7Yz
k639u/Hcokh2CKTXMkZFMDn52GOXnbACUcEsTV0CVZTfWCpNNRM0d2EqqBX9
DzWim3TXPI1Qq6clVaFl+T7h0NwWUE0w6wi8LzX++aZsceO04iGqsokz0BDT
/noqZsQ154l+86v5JP9dkjTxahsIsugMYNTKW6vBbMy+NG+6yQ4kwaN4W2WF
qZFj1hfhuQdJTwPcis8kNS+84c+yTcEyEgFXT6GXIl8cxVhoTXl9o1+0puGN
rBXWFxVDPAxNavzFQUBfigvuLV2n4N4wGcAC2KNEzcjYcjLjkvqtzq50cruH
74ShBSsPqD8mdYpE5DQI2B8t2C9nGfDzCb12IBYRar0nUXwQYa9F8Zi02N+E
Lm19JiB+QMMQJ9rCTMKUKbAMMgKZ2Ar0YfwEZBLlZCK9DpbhWAeGRy+YV7gH
XQXmu/SvmKsYV5P8914uxJPfDA0iXU/VxJC87LrSS6LO5hjzZhqPSz/55nHM
wZOquw8w9IpZp5vumtFvaEb6ZcWXiUh0EaNU6qJSEwh1BJgSVS/x4Ai8s0/6
7G485zjMxJIj23cuagYl5Q+6yD6LPF9WfzLSc7zDCJHYFmIPrfQTF2+VzYtn
vAT/Tv06wzpjv/2h9DSB6dX5FYiLrMpcVK8bnHMWzE050z85VbMPVLCIJ5Ff
jZGvldQzTZmp1Llbj9ULtN8LCgni2E25NzVZnD+G0Bz7gKNmc1GuvmeSnEsO
fkjZHZzoZdCz5uNlj0ICaQurpMhmjuUI7rTFzEUB2rk871Jly1Pr7AASzx03
ehKD89P/Xcqt/s5ZsRBBqBpY7bQqGrUBngYu4ADnFqdB9kNdwitU0BsFzzeI
OTBLplFN69uy1K3nDq2z60GO6WpxDr51pGBQJfIZDNcS6s/K5qP6tb8aPvJv
Kqm4AYtyT52KmU4C7AGdfYAOX5nQb4ii03U7U1jDnZYYgn+EH4qJ/y/QXm7w
ENCR9wfgR/8YF7Gh6QEN92iXN33v14qo08iL0LXgm3cH22ldKRYGY6v0At6r
MxQaLiGA+mogyYaEjl3YO297StcihVgW/yPl+zRV01SmngfxmhyEasKJhe9+
uZUvPnRoGR7IPQn+/Mr2noVkS8t379n12ChZ5svW4HjZXrHRwt8C8rcQrwWJ
slM02o400fdWuNlHlxH7kO4U2A16Zn1rH+728NZgTa4SkIiLSWXeQY1yF1Bi
4IogslYm2Jqv+gkHoMK60kNS3E5SzStFOSpV+O/02b/6qZs8QjK8hpT5ujTi
z377AKLrb+v8IqQTpyldnkqaa1EojyCQSAmCcxKUrEUPrfBACAvBXXQ2Bn6r
nvjQsWJeAYp2s8LVe1KAhFoRmhw21xCFaxabwo4OHJA/2oIrpwRxBjKBtbzz
ZtBv2i9m91k6obnYNSOSEvs6g/k9HeHsgqylhjsJit4bXZ4u7q0Rry7Y/jsa
CC4/31GemqL6v0tJpX+MNdhSyIqJaSTbnwP5f+bxRMbZNzg9IM1QhkUo/zB8
cbIboRsu3iP8wohls6ldHz4MI/KRWnoQ4eZ2BJowfpKmWH6pkkJuisT7kSgP
/RA9BsKGPYbXsfEOJqUZgkInmgfgy52odpBhUAYhpXRaSHjC91FCfvffwPHL
6OvXAedcGU+kXPH8TztlRXKwYVU0xBUz96V1ymKMJ+fQjHoKv5LYNEmuXEbD
LBNeKcwhhjWzYyRdJdGhJbtSNiQaBETPbth7OoBEDLznOCJM5Dah3qfpfF3J
N9w6D1kPxcgCPERV/w8nRAzpL6KT5lahRbxIGHYmolBTxzlH3FlemJAvgbdZ
WYvEOoU4ozG5HquGJ9tK6XSEYh1OELHyTv2hmvB8Mmjk6afen6KOm+2rMjK7
kNzt1N+osf+4O1eg5f8vZNFLz/TW8P6g5Khc2weEzZOD1pqhdl0sPyJgPD9U
NTtx1+UsAcwJ8HCCLqxDD0zRvQcKMsDwE+MoQiFh2qOeiD5AK0VTp3JQIhOc
xeoov6cGLYg/RZb3rHWc3GReDcFJMQxFGMY9kb1utF8or2eWfZ/dtGQnMyG1
b59k0FSNSgnrO44NLKAbczXZ7F2RAMgtIfcIamFZ7ER8KLj5bcU0EsuI6kDj
NIApQKGo7Ph9stJCX1BcYH6m4mrorl+r/BWC6gy5SZJzOgmtZeP1Q/AK7ayL
+s5qRZtXZBh6JeVFabLIqDEIeLowedHmMuJ8nGBC+DswM77WJSvZPgnH9Ewq
7G50GjqdRcAE0ZqCAkxCsH0cBX+BkHqaYz9e8YY9swubBVE29Ki7QT4aEMq3
mKYjebPRRQCC6x1cXZdsP5WUrJtR/IIYA1JxLY0EpSyc3NnNI/vSMIEBW1xL
4TDQPhD6wtDnHsFeSKH2X4oAzMj+Vafa7ztmNCWgcwAcDfSyblJSUmEpsIR8
AmLgwfCH4wVgb/MVkhPzbo3eOmwlNcQNtfvPTv9f8yOFuV1ojmQd/oBaY7FR
Ex8rai/Z8X92utuOyH31VsW3RlPtbmglsmDWKryxvsR4XoxGybVg5xkoASc9
61BxRWzmMSv2oS35O9ifBtAGHZvwQNeXRubBzSPlDAwNZkWPwxQF4xNaGF8A
07N40wGkheh5YWwTnjvJh7e3I5YBFLTqouvztfvdM0GHHHbouNIVDUs6WTEf
Eit3F+KhK/qVr36Z5EXDZU9EwsPF+IUek9cR/p5wJLsreBs2DI+bgGz4MBk0
1aZtqMNInX+rQkkRgLGN3CiOQlLAZQKh5rOfhhky8rwhMw55aEQ6SEQh91/v
gkq6WoKDwaIPQmfBnZ4FPZKvduDPeGvY0wiCbblXs6sAmtJP+L7HVvHf4Xae
RKXHqrSGGDxOlNQnzaN/VFGpcAUU5FtOEkfSuLd4HwCbf6JlZh5bSt0jfB3b
Fd6L2w9cwyOpxU5NRHXLw5cEwG80jyWwmFxGeJaGg3A7zDB4Ud3S0IkKjj0g
imrZ+SoWJeWktQbscnBCieg+3Ljujz3ueplflwLC4REspSrJUvPOx3j98Inr
6cFlOCU5Gtg4EAaw+rHsMo3abgWvrSrgngAt59reZtMKGAiTxK9obEe1W8BK
TPD5VTlzdap9o76oxQKWzqrd8ohIOYP4H55YnPG7jkFkhn/D8w9NdohC6Xpj
rZsSlY0hf+AfOxQfEIrD9By6Uole99cIDwPCEIYFNQedkD6a/OEppGthGSZ/
mQ1ZEzYcgLucJUrJMCzD8fv1SuI+9Rv4umkMtRNtDv0cVZ4jDmZJSOtaek3e
XbYdQWV9Cnv5zeVQhaL+BSyww5Pl/9y0euFtqyHIRyK9Z6JF4tjiv8m7fuvj
qoH/AiGlK0N3vYZWlIgR1S/R1pHQj3L/rXnl5WoBg3qHcRqvseB5dTWHeRTH
5b/XkAI3yXlVRc0HLwA6pmh5fHXfLq27Uzz8FdEEaaivmlkCArensLhsC32A
2Ju9jcifkW/bW/KDIutviaGbd3fVaXbEBejNGR6/TNBeuyOhvHGwju5uKR0l
l5nMPCMOK7QMOj8xpgIMy2rOoev+HZT38httpWJF1Vh/xwjEJWTCCJ+XepVd
mjAhPG6pnvE6Fb1x4uemuetMnxg553msE2UB9kay2nFfJyVC1X2xv8zgTIob
JyuEB5U7GelQsO4FaLZEWzxTrbfYiBTbSo6cAOmzATRqFx+ygJt1l4Wf6QfJ
gB9wQJeSNYqDYUAY9c0ngn8oMojczGrH2AD5c/KNSeiTegQhSZrFvX0fkG5D
pZt3iDk7nYa9vn00MIx+0u5MQzUZiyz60d9XyW7G2Q+062fKoLmRSM/W9zzC
hoIN8GIN/NcSMtRfFtrWyDihaRQBMPTsiGjXJUFi+im3DPZurHgZIKKmfZUu
o/oMDIP0lo85jtvUA256nG7qlgaubyZ7JoK4YhKk91s4g1sWrri1MJ4FarYz
j0JFYw0iM9GS2Hi/aQNfnKVSSLc3oBOcQjLlqgzkBu2WMJYpTmvM/M6P2sOB
XhJxP0/rvWdc//dk1MsqaQddiMj1lojLgmrq3wPRsw==

`pragma protect end_protected
