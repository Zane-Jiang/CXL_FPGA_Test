// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GGB3SYJze20f0NPlu7idsbzsacssnski5zhpA+C29sYiXjuScWeIkco2WjuS
Q0oR/aniOalJ0tMx8cH4MeCIPSPay6WDcuqCDp4lp/wlUpKa6vJHiwZN0JWM
cyaZvi/gK4JFRVOSkp1gvNhz1WRsX4vBdB9pukvKd7hW6EtNVHFjePyuIChk
xdCoKRbfDAo5qJw6JQSHl+XjUdqgUMCmY0BLPoHVdKUblK4HkJllA1oebc6q
QshdohefM91LOCy1fuiN3cu6bVhvPkaGWoI22UGVEDpoKrE/WUbrbSxHJeyS
WZ0XwHRWvvbn3UHmWD6XZvurdsBQMW/Wi/oKy79s6g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
quNo5oMZtQ5vvoIokNsqYBt5aVho0kxRfQrE1ouLf038o5qhBwGHa5b6+OHi
Sm0cpttm/wy+d//IYzAxeGCXzt3Vc66vdiyQ/9lbHBZOSkapg0chF21FqHJg
fZXPpdJG50ovBSBM4jfHzh8zuJZFPQ0qtCgTWIuve6FQ62JLQt09LpXOcyX8
tzl3RWYbomSZgnG2TgvklOAvvyYK7ERoGsCms82m63qan/RWPrqSVoZkqXPO
rJNl7iY4gY7OtEtYbcTGTHga7pJB2hofditwqNADDAGmInRhhV53myavndSs
wZS60NWa1i3BJgWyELtjrIRtN2PxN1RspsWjlHDcTw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NcCV7ixVT8LT1vYQe3GYAW1lmzIGr/b7eTYm6U9liRr3nA/Z3kKuN68yg6IT
C9wnW6P9CnA56l5IIjZ5PclWQsFYB4YsHSWYGUXCXx49Q7uqm1q9YI33kMBm
6Ko/2DTrAH+kYAU+C0HwPZ7cZZ6lr9fxYURJjzWSpdMFcWgaTjjN35hjG52X
05JOD4uF4soDToRrAcUYQDcdcbLev4G0hqVccZqGif9Hk0pd7671da/I3FOl
/pSGH25wfKajHPGdh7u2ySGurTmfLZfM/dvm1ISdEXgRkyxdqgMjtLaIaEsr
9KRSZDaSwEVVAUIXUYJVIyZUKJVP/Nfy6ktLD3doKA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MN1Eo9yg1NoeD4R4MF8YuKbGEK9udqKmZc670WE7cRCaYr/DT46uAYraWLwH
Kgz0bNLt7B/fXfnZwqT1uXOSijukOlzpd6bvarob6avf17C7Ien3WwpSlgRI
LpfE0l7A1mdMkXPJ6PjQUg8iUkob3wXQBEBnDQcDPY1o3inqDtE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Xv8YmqSVMDOY34EPFL2H1pvQO746bbgEX0VNFeh5z7dEWnz/IIRAuqO3kihX
gQozSJLfLZOuesXRSLD5EVPgcmGH34C9CNzAsZv0e4SA25tTgJRLxudjnrkQ
t8xs1sPgvzKABEkrmXio8BKSEdYrNt4fkM+lN6oC2zAI6um4hH9que2JuSRw
DBR9tRgXjPBL52b/Lk2Lp1UEeTfmlgiTQnTAIA73HslWGoisTRQgrCrN0gzo
Skb3H1KT8B5WUy8jQIhMnv35fOh26Gi1e2TEQj2RX5IRKRfaIgGRQNWV5z5m
oMHY/rw9r1Khbt+7bNsn24kuz7elMMVBA+Le5Se4jfEQTmkA4t60jjBNMChQ
72mFw20+fUH/4FXq5jd7cFkmDlmyN0xHj27M4uskgH7tLQ5ufKcJFhDFBNXe
mRBhpGmlc0YH803KFNSldWmaS8l3gh/8nb99sMmUuww4+ICwpikZtC2sUUlU
JLD6XY8u8kSti42nLLguSVxm+M0zu47N


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P/A5lLUhwRBRmSMR4dx7yQ+FbhfIO/yq+S0jFiFioeNuO1y5PFWhCeR+MGPC
rAPwWd2MHPo8AFlD3Hvdif6QNRGFt1+IkOKTUBs7mxwKaelwo2bmFQtb7FZo
74tDMGFd5eneha9AfT67up7ng9mxMomsn84NrJic+sFXneUGuLw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
N6K988U9l6s7qpQslyx6tOw3aPeV+y5QT4BvY0ul/W14A+oM9/o5pCSFEcIV
F/JuAGbxNMAn8AQD13HW02vWdA25elxM5EsQk2/GMTROZw6axOdJxvY9Go7z
4jmzVYOEZdrWR5IqUNUOs6w815ALKfYgscoANymyCI+tGN4yHAY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28656)
`pragma protect data_block
SagQGjBjPolbixrbaRwQk8pkbJZK4zLenueM6DKmgqx9ifcSNMBzOPMhJeTK
87egeGpiV9ruStBKVLboEodwbDpQDThuqgoCsJ+RWUcVzGCPenQ+YJDvn8Iw
Pv7MjzMNM53MqMO57ZIL/uOHTemq1owpAS8p5UcBg/4wTQOJ6gpG0BfKNO0u
viQwbBswLifMJbIHeBk4+yoKbVzR99facCzzjBeR0+XvgJAtUYbp9jNHiSll
xNPCmkl2asCfNaf473UZHyO1f7X7dZShUOuZLy5lFnXiluBczx2aZvMKLXlG
St2WbHj+apNXJY51iyONS6hYPGD15Cf8tqvgl0sRjnAb11ESSPeWR392QH6B
dXBGT6G72zZFoTu/nPyyMlCxWMX0m4V7KqJW18i/Yw1H1Fk4MjcOwSLOMzih
5JwX7XKb11n/eYoQMQedhDBvX29PdTpt7or55zlvXG4YKx3QiKatJxGgW16y
sKDK4YXdCsz+yPltJ7HhHGVmhlilO/F5wSvLJWNKtK8XITkeDUwO9Fjy0bb6
eWJcAnpBUUaAjE/9mm5KvPZ8ZbNzEch93zXJhQYv8qkOCJ0xFnxRvWntulfA
0Blo7QavD4hUqbkZRrDrbH+wm5igcErLpH8J5BwJEUxM8suONPKPBZTpjk88
VVusqvDQuwGJ9KH2FJe0MBvCoOe7wY7Gms26a1JvEwcSotqXKCBZysIi7FoV
dt+BFGJpzfu0m/s8lQqcMQGC3vWtlbDrQ5uDA+8uY+cpcAYFXNnXCfFuPfSN
38/eJJhww12FRU88NHdDiVVP7+WVF4a9fu5zDaWQlN4wWDN1xaMgci1u87pX
JUfNueq+zBMWYDlsrcJTXyRIV/npF23fUngN64PAhcEeztg7b+q3Iau6THeB
dA/dJlzg6DZv0NlnfB5qBnajuWozABLc042XWCwu/Znic81VRCqXfGHZlDZQ
CuohbYqHaIK+/8YEqAycd/9PkvFItGmCY12DalaFrCNE5P+Tgl3nVUMLXx+9
pLoIrz2WN4BYGQmhn6/lXPdJ+K53750JX9h4egbNjKL2k1LQpNdsS8L+No4E
G2Eub31YzuaqxmANfo+YLIUHh4J5+jV2bwTGl6YL/eO9xiLmjYvp3gPJRzwj
Fcq7TgNXXfpzWRekWdzzJqs3Nhx5o3SWPXsLvWckDUd8zQK6v3NwUf+5NgdS
oi3LUOPpyBv0SFkvebUinZ1A63J2unYI4n/fR+zxyRbqA7dMOu7eqEKrL3Lb
71oGG1zPaLGaq+mdf6qj+AQtBhajC8/MhOfOaI9Eu35LHHrDcSzuxpBhNNa0
3H6Mzp3IBvA2KlaKKwPY0FaQsL3xRRgb0FeKTV6wN8Pn90VYbyYvpPRvOdow
uXE/zNTZIp+B5goI2WT+JL91qlDXXl/jBMEBtuEq/ge2E4C8K4DF2jSBbYsR
LlledY4B+CSNblOFACjkYL2oP+mLYeI/8IT8oHilQSIDwT9RBXcwbufX95P2
sG7NQSlB4PV6jOkdhAk4y6Pa1dfimisLmlJnWwpYQxQ10E54LVbTWC1dlEhe
quH9Ewqz3DojqaU5jsWaVNwBk/dEX4GLySDjEPooFSh5xXq40omIEZVavtQB
Tg5xfI8lFtzkGx19szXaOaDYFpqtP/IywkYOQAQxZ/w99aYrMYMjqvcOrdUG
z475cpaCMp43YNAFVn0bUsVwv5yuEivW19I5OZOCLwH6ts8sVTsirYkWixhs
aHGgfcIUkzE7A+OlwUfvA42iorSjqAp1jKkGMBQmEymhOIWZqhE24wxBTKxW
Pa3eUmbaoLBy2WZgHnSbft+7SyjMtJg6z5l93UrokX+S9uCXg5yE4QFCuUj3
YE8FfOaeN2ReKb/9KkApsTwTGF4tPsqvcX7SgLuIiMXMvOFut9fjRD7yw9vB
vmqhftBKyRLWWH/9YJN4O0rmQUiNB4na3cjSXW/hindJMk/bfxPugcS9S6Fa
ZGtsFBBzWWJEWbJNZRx93R3aKWIWWfH7vDJz7fwbHaFKP8yi6387JV0D5zEl
TAp/RprAlPzenB6rU63L5aXrM2jj6X2FNPeoSwZrMseOobwn8IZhjRDGueGj
u9WByXKQpXhVLDykkEx+CQoh5HngZg3YpFgMVDD56tRDfkuX/MyXkqvbR0HV
HuzGJvC55Xzjp2/3fKBkNPfUTukl25+A/aHCVuAYZ6LdycmFZITJZIY9mdHF
16nf/9xWzocn7A7+Yi/unQzV0DuCNm3LjUPxU930gemlJojrT+KT7h1EsdPq
ZJSrKYs5Lz5Nl7Gj9N2RdFQpebtFmeeU7f75R9nPwLmr1eVJZal/HKUpKj0a
NcMlUIApouSAr49w1G43VaA32N+IAVT+6h15jd5R5rpxb83CInPr6kEsk9v+
lrP/mdkUYVnU79dzHcWcpRe9DvETYZ5ZMi2vv4BydUy/HjsGZVyHupsyEodM
OcrWrYUvtxkQe3UlkRSzdfPw1sP27dZ6G7EDWlMu0lt5xPD1UkkKGlSul8Uc
tzeNMJCbOpTA3j/IYwZJNpo8hVv2vT2WlimSYdT06V1+L6X8W4dtpyF3mhBl
MjpZQKYLhKCgHN8iQg7cDBxflDulw/eK/TEpqz9StiGitpmITtw0VNZxPAsm
bbzGt9crgnAx4AjmmRWKXR8stEpqsp8umF31J+kAuaY9SN5csZ4YqpaWknDq
KluLe1EMh6mWZwvBH8roRK45fk4cPfROsN2HTVnruTjy8nBvvJim4v9TGan/
9rAYv7wfy/O8yWOWT+N5cCZ2UzmVkLnNA/+I/siSdnM9/i7WzC+ad42mrTKp
nTZPsrnb2yVSJfcRy5qVS+z/8PaO8WToNiN+Yz61X81jl0sbwY44v3RQGPLW
Pp8X4NKMvestqPEkNM/piE53bYgAsCmbXaA5KJKgmKwTqVMfceWDzxV41Fua
uPwk44/+sy5OZSHXvem8T9EB6X9KLSxfaCMXbH+2zfaubQFiFHF19xn7bzke
RM99EeAtpbqs+siWi9olE8AaQs0qseD/BljboqeHE2pvSee3iq85SrEzlEFZ
d7x8Jq74ho2VOBkFOp3kqY09zLKPW/R9avwvh7dOEEmzPG8VTf+7OXwWI9tR
/S0ymPtdEqr2tKoeiHKTFlR4QzWx2nNU3MYJ8Gh6PIYzN9jsBeabHMSvHcnK
LvkbIN9BjKJboCQj8AXE7efq4iuqYP+k1ZNZ0/tU18BZuep61/hAb3Um8nmD
LgsB3zPwvxZNPVoVv2qPK+1IjhSH6/rcritnYR9v8oDm+cxsTcoBkDDEK8C9
5wqvsE5hw54SXTX4va9T0QBNPWY0CDeT/VtpZJyP9AcOd6whgRl7eFpojxff
ES3hI7vy2EMVXjj7RkEav7hqn7cMAt7/Lz116IiiIsNBq4p6m9KwQy3ozDkN
zEIBII06JzuzOxpJC/jZpCOzZNCRQ+gZy1ffnohG9O94DD+SQd73Wh13YgHl
/f6dN8FiDMv/oXKLrGdZd4Bj2UanzFvdGT3xGHW3gxOI2ZTQhDhflPQXWtmo
a3UL281q5OnWfxKJMYu1FDIZj+j/tis3CLhzY/EpgNCTmKfNbAYDPxAVT+8J
0Xlua0ZQHexzb3olj7M4T/A7XjfEPhHdjF8WtdQteyFGR2V4/Fdsq+wMDGdZ
0o9A6aE76UxhQA/9rVzi+xHPYbdtAUoZ5vbgJxitwVx3OX3vu7U4XXMHCZc2
k7zJL2UCNXXW0+5V1vL+/o1vcTTVvg2jLjthXmtMfiwmJXKQ3T6f5ISTZjgX
qsiFl3vpu9yFzCIKZ6r0thzHPAhT6ANOkaekd3n++nXzR2sDzoQwdj8QZphH
o4oVTWN2X/iiGYq1BPhcCk+3vY6g/ZryJkmZ3he46JuRvEjhvAod6lqhpOXl
31RUcqKG9hXFTeYsT7hMH0ATTWHjN2lmP4iFwycTStV5SdDgfTPHkPjVAJ9L
yanA6eT+iuZNPP8xnLmWEsb3cc/WxyKC8Su/Zc9xnjx2xu8DEaaEEce8Zt3s
30t1ERQnoIh7nFsjqnFMMqro3askaa0kPhtnjzhtwATWkO6skw+T7IR/m2M5
/gMzk8dJWZ/D2s/kmy+RKdf+T6E7UbglN0oepwYb1N/EBt9NUuJVyV4wtgrf
V7FcaytqFm0YXQ5FMti0txvD9b6Q+n95o9ka93ApLE6csJ6jW1L2ZSuznFsg
2ThzNiJ5k5h1Cb05XGQudqboiwCKjId4NUIUv7qYWf9jgoXpgoWrC63o0Sjm
syAG5VNdIxaToa5iko4ez7r0mcSX5LUUVKg6dUMeBuAEj0OTi8A3/+vPnMc1
oE9y034G6ssnJQV1RLyl/sRjopMTAtag5KMgz3X9NRZQj7hyRkCY0iKq0sv7
2RDhWVShlYlszxkWvNvgJ8aBBEvQXFS5j2WVzkiW5oS5LzvdNrn/BQ87VFra
cfwdkXoePE7KDwtBkqg/TthUj6pV69dFikkKs98/+3cTyGlKbbFY9i2/id1A
NeTkVelZm4U+psE2NTmzdS2pn0SMv92ok0gKkFtKMqwYpscXZzowh4J+wyUX
h2qyBzWUAaexhAAgEaeuRreJXQSBbzahvIenoMtGL8vTRdgPqWKBN8OKjPHO
fW15mzuwAiiWYzK9n4LXa99prFofsip3mxI7Y2RutXPzYuLDAow5QFbR9ikt
C7CMrWB9zxWnVmzy48d+r2a0KpIr/Xge9RPhCpO56jgQ0uhl6b9T3/SJ+Baf
eE/5VhdiTHRHKVQ8w9kNw54TeqyV8d8uehfTXjZhAQhE087sXJuRP9RnhwZh
PN7iLh0Wosb5AaYQpJPutbrQ3KVBabQY2UptnxDEDBtoN5sFwwwyG3i+Vomu
WhyFB+qlSAgOjtuIJ6K9FVpwcm0mBIrpIqr3+aceIj/mHzXvpKk2yJ3nVhWp
li5PKcVX8Gjhhlmzl5ulHu6/VmAXhRakJzTgqKEFotieEavzESamgzRzaPaY
zkDSywtolMqVuWaCdwrkzQNu3ZUTa9QojSUA76TsFodnebgJb+nxk8l6Bclq
V2tf8sivtt9xVNlQos7RYYJLWrMAA/kFLEI8Kw+I7aCA7zrzF1IZ0yTER+KQ
ooYQ5dXIuGUaDjvFZg6hH/k8H2mWlX5ZULbO/51m1FLydRzo1zsO8JuyU0F3
J9P4O3hSS9j0LHUVjcgppVbUV+EPgSBeeX0C6aSbQFymIZMleRUnHcG5HuGl
0J5UUFtyABEdARGI/CGf8tS8d85+ouKVzC/Hh1xybOCLCaQOUANjfrQdWAk2
2FkwiiQyG0r1AB+wVuiUBJHdDRusZ3/kQzi5qAgxlpzDPnDGEeNAL06pG4iT
CwZYvmhevRsy0L1vFuLoYyhNwYx02Kd3/8V7OlJQ1G7lG/C7Zkg2auHzNHH0
OB+Gze9QHf8etxwLeXCJoy70eVoaKgtpYbMQihaQwBaNCLYoOW3sxa97vkY2
DN6XgRrTVQJ6qnxOcxJFfPlMbpf8cMXtsvU1jt/TUx2IO4D2ttpC8ioLDjhk
UNLcbRnV72KYLaEPX/ziySH2Depoo9884k2+SS1wiKLUi6uSkb5s3DgNyYP5
Y/DH/ZzfBW2Y/uwNVdggFPl7Zo8oiZXzxHD0qU56hWtoRDA6i0V6cuqyYRnT
847KXJb3IoP0yDD4HKl5FQVnGOmWKP2rtIGAVz9xmwIebgetU9LZBONj0FIZ
n+JwBoHgdaCIh2YJ0ug9E9phwZ/nEM4YEt0ZahN1qFPt3QyTIuFqqqS9fPno
PnKag2bwgjDSZbNktJE8AXAWqn9LfV4/P6zIz75QWwzbTk4vXmDLMErin+Ih
mhPdm2Ed2GF+OAJigc6/TND/s4zMI26LzndvdfTKuj4ldDtE6OYYXoKl0+t1
TeP/0U1yQqb4j43r8VpiP5f4plAsRoWK2Dh1/it6GySOqLo5G4iMvpAwx91t
TQuJmoOwIWuKNKuWQ/3L3ahNhUdjwkdvLmxSHtmkBmiYrmprzsPwAlsvwgCB
yg8svBOr5w2WmYL3XcTj5BW2r4zmM1vezeTceatyKZJrq/STlD0FTWMnrWQR
LcA04CJyp5D4W95xO5Kscow18CrXAfeB18qC4n1OlpKc8aKmC3qu0rLsLdyz
X0kr0lsn+FuCd9LrZycFuaet2hsM8n08/akPJtr1imaSB2SKSVWvnlgOn5qT
lLxRMsVA22lSpWyswvmxwXoL/KyG1m6WtLYaiQm83z+586tnG7wfRUogaarq
YKEjwKF51sp5yAN543zSBENZ8By6WTAys+HamjE4oJ9vWn/V34MJQlIcKZoV
r+3N2fesJV1wpR9gfeaUgwrWfjcLXSaWfwLnnQZfKY1FQtKsUAgKq/1paECQ
4RsWphgT5/xBG6bXOzrkCa99rXo4aEmqLOGdGlkNq7322x0CYB5WlIMQt8PJ
I1ayziQiBPI7eXOK69RMDAcas+maJQYKz3sLLXkTQK/Ruqx9VBTp8QH0vKCF
Gd9UWhz7h9w6UArzl/DQ6HNhrsnayta3F+gvYEU9SyPuPI16kZ5U+zSjVQxb
PLKc+ppHp8ktq/kojpriHln4NXROXQkiyFSTfb4yXbULon+CtsVh6Ti83X8Q
BmvJnVbIs2Nn/Ui9U5f8r/kUPc8PlWQukNjx8dqFODwDPgmYa1aO+axQig5G
hcnKkTkaltmAT5NC1YcCYHRH46b3jdGa26CZJU8Q3HAqoT2Bvnlga3SB1Wg2
SbAPTewRUwkQXpujTUkg7rC0/EXBT6/22BIz4SAUdLU4qG8H33rM8y0IA/J8
RCTsSajE/7JdBliv33YdpGXqGIC84StQsiRtLjVavqoF8iC9TRl+TlLcFhhA
R+kFIkfT8ctv1zIcDnbrsNPw0iwM/RTkqG0S14H0LBq30PkjyRZxEws+Z8cY
9tYNCmwi8hPT66ih1ggWK+D6AklrHQQxZtuUmkPqCFrImCRQaQ3Ej9TFSDQw
uM9E3TRzVFXFYPnGj0K9ZobPT8IxCqoOakrIZ+wMLpZ0txtfU0lzjoGbQIq1
9ko5ip42yodoiD7ITzr9WSFnN00IDvZn7bzgzppDoChxL0rLlEBYOEs6E6c6
dCE6r3OleS4mZp+WYau/gjs/8A8HZeqWUf9m8SbCbX3OQX6vj2PymfY4FRI2
o/eok/Tk4Mz4dIz3soMUNuVUhgo6AS8zN6bpYy+S6U6dRbtteBrwyrUePDvp
nDU+o99GAxyDZikCSQb/0EEvZ7ms4N3Lo25HKugS6HYTojmUEQwmoRnJ+kVh
pFUueyMmpc6KWRgpA8XB0jDbqd0Q5QknsxO8H3yWBGp/NIx1gEwu0G7RSHlp
1ZQ4OREZD3R7VVmyD0HWXBo4EUWo/xsT7puZxgq66DFdD1KE+L91eP/Usf9f
qvE1KqFVtBfgsKJeYtdBFxJPU3jaZ/g50MH6AXnkzE6GM6bsTaanFKDQiul+
WZbplJKpdI/s0vYMvOxFPGPRyPSFBIhGvLhlVQR3Pd5SQ4VldA4lxXKv+5uS
3nIaPHh7FV8RdncPz8BdqgKwqHljtkbP+DjePXGNzPFDFZ1jzmnhhcUSReh2
nMPrBVjiXiD6Lha5iBMXxj1yKHxPb+15gJbE48Zk2+5dmL/RNeMp8a519IUg
7EGX5+5u0amQKEocfOvVCM5P/hmkwTk8KmxREuxTk0rEMGA7oHh11JdkTXNx
i3oKt5gVtLksr1CJxNnlEwW/WBcHAnPs5/b4RHZXOVXYJqSKiyFdufgmUbs8
eFBqr+AX5QIXxfFBhcOp/HraWLH/d1EjAmmI4lNbsjNMkA0BsmCp3/VKL/1Z
rpjMXyjLZpB3mVrDw6vAo6K8cAVSs604mOoHKbvsRUiqbiimdf45WBh0z/qz
vtFdkLEzfIaustf+WbKU+o8JWk2/k1ygW1vbhwcqxBI8tjfJwjqYsPvU3SEg
xlGBrBdf8pomLmXM9M/kafqf2jZHndKjfi19A84YQyuYhi5JLAKPienLJDkL
pgKJ1u7VFZGzJ9nG6URyYuvJm64oI7eIRc3YMTD7MGYKMKSL4AYjra7n7V2J
hWNSwnTskWasNDbiJj/OT94/MIRg0IheihkUBNm2TuBhVnV12TMAphFtNMje
jYnyfMwqMvw0ZFN6Dz9ELhDHV1OWbUn0tU2mbzTqEeo51ya/ky7FNRT3U4yy
lkjQz8qmxPMSv5xzqMQjFLU4Bs/dlsCiMtZKl/cpZ8kJMdu632XahsZKvmEo
+46zwW/3/JabkgVDrQwHg7sFUSKAm+qY2lOjJy52XS7aLr9OZfXpQyr+4bc1
d8A0MW/OJQQoqYUbLUqCL4t/TvOwir/KzTifUOZNwMMMAbfIfYMLmKaM7ZCG
LMQ9IIlcdxHR1j5TbMD/bbCfQHlxmCbkAmjY3khzV1NSdn99zKz3RDKklT9D
vLeq7QSbywJVLNVZBtZwD/NE8fpLtp5d6oGnGPRmbAq/Dy2mf2zO8jmqtAd6
V+WyKXxBdb2RaQa73o8SURnwVBcZ9Ofpxm9ArkFjVR8GMF0gMlGau9k3Djds
DtXFKtHv7gk9NO7nMJOg+Q4LtoYxeyQUD9ThxqJgaPLaUn7RIvqnV8dcWS7d
Hb6OufE6JG3b3xS8nVYKhMElfnXDXck2b7ZuhXGhVJYOXRorl7V+SXOKzFC2
xUokvHbW3fr22m3Ng9RsZxp2jk04apbG87YpVx3hdhoakQ1Nzu3Gkzl1McBy
cMsM0ycsClvDkW9tjnQzQd+v8ARGczL/DaKXeedFRM/iJGQFdMv8IZofhX8m
4Q71ypxrHP01XI+cqQmhax90xuSnNCV9OXLtqdLQw02dxEP4yLAGq5MsIvWL
i3TuHUjcuYXpp8QH3k93BBS5y+/dHjGENR3b275f0IZozj/A/XDurZP2H290
bFFhySGBN+fRMWEfoEmpp4Vbyh15UgfKtq6MTm4lRU/dE3UlvyxTwM0vdAzL
AqTsqQjkH+ndaNiTt8bFuei+oVDbO6LXd4Yau8ZtBWBDeyd2j0Ro4ecPu/WI
xWG+PI67/ILVo2igBvLSyqXZZThKFdUZ428e5XqBjOwtnR1hHlrm990/R4ka
K2MOGgqd+hF85NYTxmffK/r9l8jvIuQlb7qghCrfmrEsQEo/J0alfFc7R6/c
tE2K75pu6xPy/2klzL+Ru4yYHGjEd4FDef3GjNVGrU8HP5vuKHdYCauZ6tiP
/vWPBBJPH4w9PFL4MrkrsCqEsTYIlgUXhXXo1Y59hX6I37KtXCDFdmzZBBCS
fcb0iQzT4VIoBSKFTr2+dcIy7f05/q+P6DnyeckRhzcokgbEWZVBN8qu7yvd
rlymdVPQqKEx1oeYmEqIfnmPVi5Ng6dy3LOmcSQDo+wSod7oXd0SOe56jPUU
5bB1agXopF+SJw4C1hSh0/OtcJSuATMjTbSaq1ZOYw2bYSFDfVdpEZ6tX3vf
eoEnkNmx+k6hdG9rm4vTKrKK5OC2DyeQPIi1vqh3H4XxyYMusGMDYFu1eJY2
xGwP6dgB4zLeb06ONxZk9JB/2Fh5G1L2i8kB2rbSrNHoKLflFvLc4XgpR6Tw
GZ2vqNyqQuTgaTSbR/HTgu2sUUbj6xRaDqaKFz2YKikLZNo9FVZH3QeIGpeJ
4wcS6IHB/5KUo54gbFkur7UZK4HjZRZoDF4Z8OezUcvDDLp8q54026hJsSpU
eRladqI7tlnH4EGqOVdBlQx0vNjAYyNQJoMN4cu3Eqf85DuGbJsDRp6eNqrO
66/ul0CVu4zkkLDop+6jkSBAHXXr6/qbvMIyScAIqJqVxH8Hx4vd4UYskkQT
1vncMueQo6FAgWPOFziKBOnouHidzzqYqz1b+wtvm+QQbiYAtsyKQwWFPGgY
3CMY8mUjTfZ5O/F/oTKfOliu3JMQ6b/J2cZ9ZhnmsvY7jjmLcm2cMxuxmv/C
0jEC79eTCiTT8/HqJaKLxBFOTgZSSgrDUU1UP+F91QEEsh99UxBcitSAm2tr
Wcw48L2rLMffpqlOwWYjJo8S0ZajwENsiWEhFIAONaQ54TLwvRs4scOsyscn
drsxoaIXMyr11OVbkQaEcdTRu8erhQ5GhgEhvqY1iQKtLYfyU3gO/TlnjAUc
Z7m70LnNX5Gu4iz0FvHahXzFL0jIXgmW/pXDQ7zdi4lt4YyO3RZeEZa0VVMg
dIGfDl11K6iHKoSZlRJuZkSoMIkqDd8Und5MeU6c+2YJVby7Z0g0vjOc1MFw
fGBpUcqli5IlM/9VHmyd1PRxljSYbfwOqjptLU7NbmLtv4ThGcv0t/91Z9zg
hLtZ9oCBn9inzi+SJST8v/ICCKIHEgXNZfRyz1e3wwPEVcIFZJVm8+J4TySc
oYucLGNR2Y6oYRAW1TP0uGuCUYZrajIuxrd3HXa81AnKOUtpRNpBR82lxU7J
C23pPkdnwUxyri3iNxQP6cM6sg3+2+mPWlRmuyh5il1gLOE97aH820OejH75
Lj7J7fEqRv/NVl/BRVOg7WXAgeoAR6yQp2+ezM/InoTvK9uPMwyOBOshI9rI
yYKZFq9N8US3y79bw7MsKfHWef+o8wqybkWAh/b3aKEAZnCtGsk8X1roptsV
Qwy60mUFjVX5JY7uzyQIXbjLx5otUusj2I2qDEmKoqQ9SHu8dHK4a+4VeghB
bOXVFrQfeLdJtjSgaI7bEMiVtiTCXxeB0+TBmo5ssWfNwE6u+sHJNBoOVn6u
DrBvM7Cqvc0HE/wA9Ur9qrcswXuUYvTfLCVgGTkPcINaOiJFqfWIpkbuOak1
6AWvHFhx9Yg2l/eRyHWDOr3q1KsLRLWj+y/I0G2EjTmAzpac8cp4RSZn2noQ
/1btMdF08gWf5b6d9W5blz7smcdsz2xGz4bh9avfz+f5rhSy7j/1IB4AwoAK
eEp+cqe7KMA23bwPGXJ8cBYTA4vIB2Xnw/zOcVeHQvVDIgvVm3dwBM+2vh3C
kQ4jCCXu9hcq/jM7JMu+vIoskvUnC/r6eeSdniaqDMMZ/xzHWclVmpQ40TH+
lUzvQI5A98KWHEOOmmRdCqfSgAUpdaSRO4PFu2E2/3bFJMYRNIi3xfrF2mPt
4QySdgOJs+DC1pfkqj7dBq8VgdEbf3JpvHUVZYvyibP6qTzHLMWIIxdUAah/
wLlzzDzpXMhFLsi8hkbiBCC4ogYJHw98KhNXD0zgYOi7DrlA+pPOU+Gk1UAB
jLKLDIRD8NtyGq4Zo43bbByXxPdz2DZ7EP7h5QNpMibhBacdvZuZM9O+WWha
NIWFyqOj1RsRel1a5hJK3ONY8CXI+BUf3w00RBOD1IJhe18iZnnEvAuz9Sv0
TW5ce1GAry/ZU3VrUBCpt0iXvhVkvRbQUHzYh1rel/nb92TVWDJMY06lZ+IT
Jm4403puV4qwE3eK7YmmKFZNO7fzzFPVVvnG/wyxOqL5VX0bsNw8C2+odiU2
FFLBaN7KHN9V/a7bGc4Om0sIiozY4uZrY5JeayoQxqwMusdj8MLoqIr6+MdW
gwFc7UdigOEA/XjlOEq6xcxMhiVo8Z1djLE5sOFXvvDB32HE2KO2W3ua09CL
ZvzOyc+dAfL1iHdSe02n37zfyi5tO2a2f/fIsUqDRVCTkSaHgSupw7QJ4HW/
5FJGT+DvYq3YBDipahPCx2ouiQ1foxa6F2WVZSYKOAMLT+koiznntVnEVcD1
0c6aecWoDwois9HlkV+pQ+CzSl0VXJG9GNmu4eQcTspGN0dzzIdwUP/10UPo
h8+8caUnJF8Ehrx0uqo/ed0jORxNwY+zh+S7hXST08+XiIb3LWChYX7L/15+
oiB5rlvC26TR3ItqeNv05MkM4ITGeagGsSDpdBoH8pzTphem01EZ/QRGvanR
kHtQEKRvM343CgWLp1+vDUnUORfy/p/2RObkNy+ahNjWHAENTAJLkKhUS6Tz
Npaj7QF6PDkmGg8SsS1ofd8m0tFkurAQ0eCRlEsbp2bTHTZDR9gtcP935s5H
vbOVjtt4DppKCmZTuBerCVQJMMkq7vMzJOSLM35zZfy61lzqss0d9cGL/st7
KysV16ZPV8tXzUztnZhGqQ4poXcKfBf/XxyWT1g5KtvcWGYpoL1eoXOwrlgw
XitAPF0fNgeEsEAjnCtFCUIzN5Uolhk9Jz3hWNES3uoxRp/t9s/kSA1zBuLG
PriDDQdeKcdrI6Zvef98XKEJD/DGFEytaqXjZ/vjysJRh7BI07NRuCuCBc5d
G7UnMEOm+cbuZGnO3AHwUrhocHnh7x63CDiFJuhneTsND0Pt1j6f3AqhalKd
lsGqyCQ5lpd4Bzhqqxi6G571/lLa/B1nr+NBdCG7GEtXLXcOewvXSRGSmHk/
+zVzj6PoYV/pPsBh1Si8jOQkttgEtOuezMPm8uaHeR5L0jmP/bmnBL49DnE2
szfRU9lcbfNRk1A1nfEzfQ9Ic0TJ7JXMGXE2YsBCYloEmlaBdmPi8XkMxzdS
/PT8S+tOEIgUjUaG9xH3P1eeiw5dYCNtH1/EIILc2hu7GN6H2UGc6FUrhhBY
OcuX6CRwaYeJVLGavGqUwo55YK2RR95elz5kLWT73asQZliojVI+x7reKeu/
hmLf8q1yyoFgMPCvgTs+3GklNqyWpSUGZ4wrVWlDIlol77MfCRd/pVzuAdJe
g3Ga2H37OnJYCXJZlNszZw8IgntLR/KLoq/1FyHKX4Q1m4tqLXoatGy4w9ME
noUvJLcnkgajXjEwZWj+p8FRamPaMAIIg72l9l+A3FztRV6oRxjXCibdlBVv
5b+E7Cv7eUSoI8ES3oJZCvkUfpxn81K+kihCvLOahAUdixeQ1AnhYl8RE3kz
naOuWFQZTa5xhCQcXfz+RzFy7efTk/DQ5tKluFgstAVvR2s0B9iyjn7YcL00
Zer2XAzJTP3Q09ghYBU1W5keseQHECWr5J/RWjM68aSsWXqHWXoqskcpcbh7
dxRYeiMQD581eHG/LT1zY5IMFiNRvOlFfrRCVFOb6CmcDq+jIauIMJrDeWzK
Hz22MKi9oXFDDPhHNvsjJS4ClW1aOHpej9nwHYg1T0ciJQ7Og55Ick3KPfh3
8crbL0pCJF6s44YocVMQDGhpDPTlU/ZBCR0Pq5xDq2Fickfr6Z9jo41a8Z2D
m8LsSIbeg8TcG0yKEJyjojSD/dNve2RvpBT9Wq3fNW1QeHAu9MUoTHcStq2Z
VzFM8l4nB5KCWeut+yGVqlgmGdkb+pD2AAAl1982qLZhbqDmm/Kh3JFnrYO9
cSHE4t17rPpLO9nAVKoTnQ86ApsX/Mu30i/l1uwXSOb/ugWtbI4nYnGxAUbN
56uemHrbwQUh8CvO7DDIUiRQI2KJa5iEnUMHR9yEuowBSgMeEKS7aRWGRIv+
i4VQOUF1OI3b6lVYSXzv/jwmbgh1jaIn0KXeK5U7rpIGIssA7IymQj85n+nu
xAPUenvoV4atzCjxRNgYSUtkjn9WT/wi+xqGIP5nJ4ur39ksRWJZORdQfhnS
ParW5hL5dZnzML062cUDPxcBi+BV3p7uk+mjqWFIELr+j+h0OaIZWkNEjFCR
ydlHnagMGa4rYArXQE1RlsEd9i++DDB+kqU8RMb6JEJe9XHWrUX+zWJp1Gd2
Vz+wwUsg/4gwyp4Oxk5yUp7TlI32tX/vx5HSL+L8m1PjvZy46H+kKKiazy/s
hjuED8afBURhUTgTfsQp7b9dizKtzjNkcZBgFeFEiuYxzBkLvUWBCofxKnpf
fqdDbjoEV0eREI79K+JDhKuvjhT5kyXD7X/5VqtJLXeYeFpKzX88PC1k4rnJ
MrEz/BqQmsY+RTedqZq2lrCMEAOLtcQgYj/Tjh8hAhUwZ9KJr4iV5mDfBMpK
AMCnAAep+DDf4D9xbU4Uq7i2KMzDtJpFVlS5x8TgdHbbaNH+4KED9v+itJ3Q
Bf0FnxP/NFteY65nfKIOWuiLHP1r5cBQS2k0kipGJsc/Y7dSGvJ8CkFHukOa
h6he31HWOpgbZxH8pA1+jQEf0sNU/ZO5AoIRUagMtLCyqZJ6gHongdQjVAcH
Oi4uwybYE2PykRV92WJgfvju7nPnrR9eCoaGdKeB7zjqQEwJ89uOOti7VtM8
wlw6PpdmOOSm53V871+vGeSBGwuFb4ZKIwAQZGiLAS0rkxFES2wUxAn0OsPv
Q8vRQTOuDlYBnEfUcSrEQJ4bltl+5ov6axd5uJkfwyTNrYOPTkv9EsdTyLyV
X2tES+dcoHArFndbEs1Pjk0wDcS+aqbPi9mTy0PW2yeyItUzfjlefB+cos9G
io9t8MCWmoD9SZLri4of2Lx22kJhIYk0if+HZ9m9hiL7pDGczoIcWxyNMkH6
0pkdt/KiLe3CchIlsaxjO7cqjpOqMM4ebxzMl9jD2ZgEEQgolpa83KoCB5QU
/+PLzW91Ow9Ev9czKdicjQCeJnqi0zQVGCjMVzxVw50P3LmqpYQV28kGk03b
0eSgjN1o8ADhAzgodSR0ih7MwKjow4KqGNwh+FMlewTk9xJXZlVXC9+wbwAz
b7vAegcCeI022l6T8jydVzJS182LGki+uUZU6IRvmwWEI/FGVNenUbeL0U9n
XEZ/V4EVmfFSuWqs7OHtGnt2Al31lczVgwNowyebGAiUyCRRWM5/SbsTl2cc
rQVa+uo4Xgpc3XkZUXnBCmNRx+Y9eBvVhrQ8BZCRLQ7eMMtft2pO4knIhdtV
39NfauhOfQvHTx6RmswPoD+TND1m2iBmHUHDsjN8kUdQHgNemcbv/HLaygM2
0yHAOpnTf46sH61IDgVApCHskbTSgVVVo6R18r591VzGIS3TwLp3gA1O934N
xwz5+WteC5q7wuSBW4IEFu/ukou3ihNB0SUs/HO8+WULbYGlsrE8zK8UuvDj
UaEuMakvpAFnwgvjVcMCg+bWFyRJoFbgaP/rkb4RslRQgQnUzhyl8DwcAqGK
sitt3F39qzInd75hOFDwigeZYR5Stbf0IohTgpTFFNinEJKoaa3n8l/U3Dst
Ofx27xQ7xv9YA50GeeLc+lBsKciel0VP92F+GTVlCsTShjVRhPXW9FGcFWdl
fvTyri2Q16f4X22c191gwSqYEFKeFAlkruB42mWmkrD/3YFY6KfSbVgz62Yd
kePZ8fI32GEGm9zt285HA4tduyprXwqQ2bXFOHbG/i53Y7Xdm4mEqgqqf4Ha
kiWBisy1kJsvDx7V0ZtTXF0vDD1ZYnod8dMNTt+YQQ9OxBTAEc0yTA/dejGh
wFHBfcW5yg3+hlTFir66VZ0z86HhZ+kiAYJ1izmHOBp/X3Lm4/W8O/jUz0Ux
y8yuH26OzYnnZbFxZ2iPWqIQKjsKJigPtf1S22XY0eTPojMfNI4ClcieN/65
DW7hMcAOTD7TVn4CctPDyqKLzvZRk3K93Q/4RgEJgeLcZ4/xwyKdmVxyVlmH
x9UTQVGxImDYNUuHeKTZz6g+SEoU9+NVLbsuBgsbM50Nbxwp/HVHzR3WWPdF
nffeWOVHbq17n0sjirJ6B9B9ctDYSNf+eUKZ2LM6ebVP2d2LhhMQfgMZo27d
pDdsE87iYoHyM5Cd9vfO84xFa1K1nfufWhwDC7ICED9rQHniVvXdro9asiPe
MHuxIMtGRkd6qALUqnBcur9Q8hyH6hmsMJNHH9OnV0rmbVFqWMIvbZuvlw11
z/oQxb52fNLOBfydgDN3o3DtEQHEDmh+oEsszkSM2F7PK6iMk9BgY+S3ZuZA
JC1EC50tBpD519SOWC+bUgjmdhUV6WDY0Zpkmb2ya6ptgJNIh1kaPuO3iKAe
LovaQaFjGfg1JJAVWedF434ljDmOfaZhwTDpLY707+qGnl8ABp3M4wLDRO7g
HTXBpUowA/845zqpSB4MGbxe8/3YnTSkrW5H50zEW9z+NGh6Enueiq8xtbIq
qqyWMKPGjrIMapbrbnV/vIptewB1iiI/Kffce2Wr1EviMMjlGwNwNiTJG8eC
phdH8uzgkdVK8W6MN5j/okWO/NunwV6XAalahjc22m6N7YiumBpfWk12yek0
e0fUei2tqcVHN7oWEMSze6WnzxXCG/1lUa1vANlZL8D0Pu+xS6WiVcUqd6xd
SwiKfrwqlDCuU3bS3IHfnEiu7P6RhAZj6X9PqjMUCzjO3DiYre00V9vm3J1W
u8XR2CJ8tFj4l9ZRDy5sVBA3HvV0yb3XUuS0P6yeAd1d7R5GyllalGRQlPCw
yNe45qCMuLw4lvfCSzBTuIyTkIKuu+attw5H7IyJV5TTeDOogT0nHrZleV1V
mWH7+5i1/u3/Xsu0Y2jji3FZL5C9BKhkrYO7EbC0oSVxUg1IYj+Jb4etnMGy
K5X/ChlvI5zALLUQ+OooAD83o4Gu6r6fb1AnQAuL/KX0StUyWvDxZDxTy1Cs
GZkBh+ru/p7826MbLoZLmUV7XJHtO/jkGaMhtzG19EiJHthL6OcS4B2yvR57
56TNYprOBQjAUjM48Z1MO+MKGP6tLSgq5RvTXRp7/6CM/cN1b/SpBqPA/nRI
iccV1m/fhZG2ARZd6JYkzmHLj19YKuiYbud96oyll23spYAYeGiY6SkpvFSF
7dn02kT2WTYZqQCPlFgFxQErkUnAJ42AjSW5wRux6zVxMWTUFHTt//Y5mCQJ
hE5kGFFXceFYJf/vZ36edEYZc7unsj8b3QnG251cv8JX/qbU81bmizSqeZpt
0cwYMl1Fngo9qlOzfZWfTU9vRNHZ0w9b4U5ZDMTjhAiZNu5KchCVbBtK4zOJ
dd9VW1DlI7MiHbZMWUpOXfvmgra23uOrE/z+dE2yK0FYZlJyLG5zgkdFSvO5
qHBlNbebY7A6rzQDEC/Fq7POePwQNKad7hpUOjzWo3muIFllG8WBXkzPQ81g
T3C3MWyXtibLQZ7qw+Zb4LIXMxMjpT4IZImt8oEoypwbox9IBNzAcHAVbE9K
Cvwixdt1vktMdN98vxtgi5xsJYS9Mqbm5CHv2jfneERpJH6xdSurSVWuAJgk
ak+eTtQmH9811Mlu+Ouh0hhTc862EEcX4GoZ49pBVoxYnNtFA8heo8yL3/+v
StppEdGLDzFRvDBhVToUj8ViJeyni+MW8beDPG/E9wkfabcK9Zvu5r1quQMn
/WQclhl7dyqZEHudMkrWaPP5SeHiHkwgxeCXU4Gsjq91ahePJFPn52gF5RBG
5X/ROvCYtM5JWC12Ys+i8J0UzDwso1dsy6j+e9Cvq0FHGPx3hTap6uBzU7zO
s7EfeBRLv6xS3phd7WU2BkJBM/xo0seZ4oEmjpwyMiGYQT2jAUEMlPBvOi7a
nDUYORtPQ9SAUxy2GUtdqXG4oPsjOuGY/B5K9C+x/sPUfsc664tDj6HVc8fL
2uFT9TGA8rrJvP2Hp0LadSigoyDJgD1XyrtKEondv/8r4rlNF6T6q1mezo3W
SpRj3nOJ5I81fKjHsGMeNhabKnUMlopRDDtD4iawMCei+VIupnnCMEbYF4LX
d/lA5x172Y7MT2J26PA8B27jDvCUymyMBYBo/AZ7uJzMONTpwplauz4AcZje
XM8481RpcmjgdFFjL00HJQl5o/KB90Ipq2t8gVxUnNHAwja5AJ/oqcRnFI8u
ccGwCG+rz0txa8wGVm1XbINTrH4bNUuIkI3gqM3sm5TGfO7xhvmRK59Z8qXo
NQ4elO9I757dWtXc8i5YlyL6DckdvJNFgzD1ZCRrIyvK9uHI83XpFM9KMFwf
OoIY+lOsrj6sLTg9vkimrTJdyJH6iDnCKMA8WgARCLQhXm/BmfZDqueTGHPk
obpNRjL7c5EOcBxiTJdiMGMdR1vAvS9Q7AcQIyIPp0hURyUrkLZfOSyPb42G
2XBEc4SQhGN9HR4aoak4Yo4sM6493oXeNtZ47QubV1v5nGkCgDaPHt5rO/Qv
okYU+s03gpsDatXfcMc8IqF/IgTCSrOke2v2wgxicWaH3iTQ/afloweRFQyW
jXWqufJQe23J1Qc51CmG10NulqKFkz0TD1MhtF7JYK48aAut4LopJN/egNDU
Qz1bSggI1Xmv+2NJcdlkVgvfIeGMDOphxMX7bxnXGpJo84EFPmFr+Auoge5T
cOxICku/rpJ5YzQ0QOZq+BSYwfPTGY2Vnn5XykmUIm7Aofj077LRyDSnHnJ+
LXOcwgLYCkF60i8eWmA8U8O1ebCx5gYiy3T6Xix9O8mNTuL66BOMotrIRBKR
DQQlg42oirHqvS+M+5/WCTyD8n3zxXLiism9Ypd5KWBHzCjuu2ZP+ZpKbj05
ge3SStYVS6c/IwnPRBk91Q4bScsmdtqDY4/7aJklsPxMiF0DlW2N10bH6yWW
1Fb+rTqJOfseuA5IDhBWq2hf5LYqYDu/0qc5iBTY6UrJ4ghqEP6gTGw6K6Wi
cY0lRmm93q73tLgjOhIfJMOjAUED0DYkq+OpO+QylqFBpQwu2k/J42jq9Ovs
+p+R5Ro2+sluCIuSXKdcDWMEf5ZAAO0s8u5RNL9NX5T5qEJy3FWyG7weLYNm
9/fqyx6LICS0PJkXSjOJZq08jREBV7vYSQMV+byOE3TD6VizbtGv5HLY2dnz
eW565RpmqIqZU548qsjuiopDYNWoUpXYdrf6N8+34xTe5rqQvXumzpxUR5Hu
Gx3o3q+UrxvBh+k5YwukgRL+Z/DAcwC49c1b9Oc93vzey59hGFf6emx88qL2
1XUcUvPA8q26xZbxORqsJTr9Zo3rsJLhfCklr37q0HmKxsVbv2TmIDpFyZKh
5trBepkWDCZAGm28lRyQp/Sxb4y0cJVH0S7Y04t1eQ5J5JlOl+NsaIzoSkFj
cmRk8U8sUMEGbJHD4Tn92DCd6bcHpLaQaQhQJ0tvPOLcnLxaYi8vq/Z20II6
IYGhTbMhaBux1lO7I1BuLg9A2ywfDlrdySayYa159UB0lIDiflsDZxR3siuP
Uz2rvQy+/CrsBA/kGLBfAqIkEHNQ8JyzVibSbB/A0aHF6zRUNbr/oXlwu4Mu
CyiJX28y5yF4hdlDh7CNuqtR7xrzciUpKVlXsxZJPtfrbhjI5HggsHnsvMIy
0qDvggwwfpR0o6CVX2BFwrrdekBn37LM3eDLRQJF5HUuDMgJrNPm6XGZp51B
8RGw4t9NHptZLGzfULJoFZ8c2TCZFUBIH1b/2gvqEDG0gxZABCYznQ9RrYq/
0ReZcsThkxEoiHGGFEo1Sd7p2dXpbPx1Oo9DMts1PfnlSlgUIJzsGcLqsKnE
l4QXsrCG4wbRkua+53baqAK91WTBqGlpENOBpoHP70hYLNeLLO2w1NP0gUV5
0gnS5XCHywy03OZ+PCh/jL/wsB8tp1YKQ75jj7D3B31ym5Ae7XObLpx7KdLC
uzQcGkCWCrffLHCOxn7CRQHS1Y9j4tBVrYTa/DXJ91Om6WMP2bpJdtXkzGaN
U3a6R10yo0fAWOMhXpZXtEDk1cHldQG98zCXjyS+R2EqSkXMEJauWnDz9jYL
tW9G3ldn8X9yC6gLSkTMdJIBI2pM8ge5fYZgDViWzScwKejzXOJ5W4N+G5qV
XIX9RzanSPYuDvY9QyfSLAHytxv2dQMuGJr9grNGFv7oVIVvEFgVTEE2UC86
4mW2g7Zy3mb/lHbJTwLjFrMctzHRfN9BYBKdlBiXN7WPYzfURZBMEOve5VUE
BCWl9V0x/iP9/qlHUzJ0bo1fbqoOsbwU6oqLgQLZggqC+8FP3jsII3Nk8wFx
Ap7bwXn2joWdgbgR8uVKDO6XDChA787Bp0r99CyylTarxDtjYBGURb+CK96e
KFUA8ADsKFFPaffpODokOEPWIjF2bYx7QQ4YkkjsEGjx8RD9blL7U/nlrmd0
pHHGpUYXqXp/4Olk5lYdmFU4uPRLqe2U6Wi7paPuXTrkeiydJ0pPabVed8EN
I4uPxiDOm3mYwBBt/3RUlR2vdHTaw1g1NZTov48Q7x55yJ3BbSAn77TKBQZe
oYejZ6PK5CFqj7cuOXzbbHp4uYlFrVe8jvZTmdKbZac9LxSXyeTJsAo5+oOd
oIOHU7DAMyOM2QMwUE6qVloV8e1Xv484XwGQnq1SL3JT2YC79qYwRE/zPUlr
jHgE/MSql/4wNN8/YFtny/D0qsY37Q9gtkOSEkBfYM961XebFwuW9INHR8jt
jmaroS1zg1q90h1lB78cqe6iRVILdeR0qUDHw9yX+gp0Bzt5o7Z8/FCWOFCI
3s0gLasdFwhw09j9ZH3xz/IgXwJ9cTPV+7fPabJUwpqWBMqO1hQTE7PjjanD
Ti/7V/+rTRaMbAtIpciKYmNy3dba+LaIwW1/6szauf5NswGy3yjdkkYdwkM+
40Fhv8yz20KpOz2kDt4a9k79e3E2VVxoUIOTIxovkAfrwQ8+KgTbx+5aZFre
h8zMj3PUzY12Yz/9jzCay7eXwSjtIEArsIKn+WuABPcMIsreB/1SuIMUmEzj
XdYxIoZ4Rpxpna6qzkGaCTMR9aDVgetMhw9em+ADLbUVpfBTUKoaxv3th16P
MR1018poNoddQKgVGQSgI5V92fP3kxo+2hcyJeTWeL84yVHp5lLSHmyf80Mv
rSXoGG86429V73To5/sJCxOqUzheUrWyblQ5v7XHpI72fGbDFcSDcnS7lrC1
176Eszug224bFwZHoUSsdH5OsEybv7YB2pXG5ppVvom7rr7Ej6i8twG/br/1
SazbwxgWXiZY2ECXnemIdNIQaiTqA4Ab5frqUlz3UMKHlQCvp8t72CNgOXH7
HZjz2qT2tLCNpsN/NpBDZJ7JmQVZVsEqAh1SMsq6gPsPWtz1WdoxQ+UWnaKn
SZZR1t86dg7JM0jTs2Yah319q3+q/CrkN9YrieRmdbfj6QbyPopHE5uvJPox
dz9njQDNaPdFcijVekA+s2FzkuWrjSzAC4VPqCZzsoWiXrcw/MPK5+lD4Xnh
XbsZl3idd3McabCBkQsxe0/yGl52TOqz8jYI2LYPiLMLUo9Rn3DP1O/UFbjP
X7yIOSBO2x6PN259ECVD6PzrmzfG12JWgjKj0J5GrBx0ubdiMcq18Zx3N21n
4/QUO7WGqZ+wPFSFZygTYbVvqwVKavv6oyUqCy9Hdo+B4JLhpt3EO475xCoO
TwXnMBMZLMRXrrqC0HZeuwGylsczq9lzCSoor7D31qof+SU3uOEyriY1hnd2
V24YhDvrZjY5RFV/RoZRS8tQhF36UMujDMLwkpfy7T0zrjpnKjG1U0mLHFtA
cOX9uwcVh7JDWJac68q0c7E8NiZ/7ymZO86wM/iAuGpe0RvBOMfjYgw4Cki7
DG0mqyVy9YDnUrwhbfHtA4o+cOTrYPGEsE9yiEeUYQXB+z7YI6qxjB4wxeTU
t3my2LCkbV0mI0AQ8REHm1cH6+qmLHSfJilSw70YiB2yVh0gIDfxpC+qVnts
ceyrBx4Gymb5bJMhIYFKqPx6qFWASd5OndVqV0EnnL7XjQniI3QWQwMmi2Tc
DiNytxsrxNNkrp+SWXE99rpSP8wYvoacm9dOTdU4VhRoL+l/1afkkvUwALM5
FwJx7sxdlrP5p3lLIzdrKwgeruD4xDGNWsJrtHa+4jh10WQFj/wiBSME0/en
ZCiBGzHm1/XhXjBWd45KUcjoi9CXKQdXYQeSAu7ThdPyKnwsmkxr+avEKBW1
64jxH2I20ruYJ/BqT1MIhBRcYcJt8sTiyo5dbTaxI4nmKnTzbNDbETirgb6x
iMxrsYs772HgJLT8WyMGYP10Si9iCzvJhpKalo1Oe+d82VaxRQKyG6uRLIZU
YZbMhbhYcLBVba/XcrN92kiWrdOa93GmX6Z531bgFOglEtT53Pvmu+nfjhNY
2rNqnY2dBP4/oF5o7C9rgcXJW6W92XdJ3C/R2TZD0g5eiT+EBQHLqqKpuK68
nWLVMmHeyXD+tN9V4Yj2pLSzf5omN+AdIR8jLwKuz4Yo7gRt/59uCdYs9rIf
7f9TFyoa0PQ7PtW7cdoPDUbAeFLPKrlrdQHO48TXeKV3W1WavAXO39Jyjm01
UySKTwmFjKT2oqv06u4+V0MwJVqjTJ/FL/EEZCb5QIv2NbX0wBQQ+TlzvKSJ
Y5E93hQfcHzKN/lsjACgBSf1qJyctEAXrBW5Im2zxLnyKyy7xQzNjtY9M+4a
2S87DMByRej2cvo3od9jlpnLVksh/iQ+rAPCkBp7sBXcdYivSqXlTIrQ7wh7
rzS+b1P1lSx3qWvk8hNpahISnUWuyTYLGwVaVF6LunwkpXkJ4vfGYTaJzlSs
7sVyPkCV7VA7c0yEFMVYCmDAIXFLPMGBf/mStq4XanRhs+PAPbM9Do3dtE3E
aGWWGos6Kdiy0goM/TERCCBQZBjdVN3mYQshnOZYQJFbp/BRQ5niJWL8n1kv
2erkk+AoSSIXszgB6gbzJ43s4hu/V94FgNdOWAuOiCELxjuUMMc2UHbLg7mz
7BZVoJUV8LEL2sCaCUJydelPwZj4G6Ou2TU01F2DNZQVJV0C0VrEeApSBu+9
0qTqQHvNx/WCOWsj15Nhhn7GPrS/aPUdJozTJGD5sdJK44sQSwA3n0Uom8da
JV4NDDdQJAWZBZCf02vXOR5FufO6bXybQlrdD10I6vXGh82A+qy7QxQ/ONSE
/BfK3SHWjzZnlWy1Itw7rsQSW8Iy0+fd59DbNtcBI3IWXFYZdNeTNm8oPN4w
toJHE+ZtI/qML4cIUgpOEZXMJ7KhjZeRfNL6jjInx+ELG8LXXLcdkNGjgkjO
TV0tmHUQ95M2jqfHGSR7wp42+ACW2YlUfQhTfiZE84p4lyG3coSoR4e4jxuQ
CqtnPwZ10vDoK3+SpULorZ0a9nTipiW8dCHl7tAnzPnphujQjFnTBpGPlxXN
ac+TWqrO/wZ9zrB9pNduux4kcRhcxWk2hc4aDWaVx62728BjBcOnTU1hQyxa
EeFDlDpdDqahOs1hBvYIvUTnI7uRTcVfRjVVWfgj5TdWj/gRYUT4JWHNTFiA
Icambv78cVslXxC6wcyGdfH5AxNQVG67NO+5S3mCn6D9NROVt36+H/9703a4
+9pYf5QqCY5hGRCbhU3NHeCZYW0s3As1goGM6okj2o5n2EKlzSODp7/hSoUG
39OHeFIoXZCZBsblNrNee36N20UWzN1B2kL3mx8H/q6m4GRAJl7agAj+vTum
ECJfQnBUZZRDXWeIIUhYRcZNy+7WFrfggIwileIW+atbvqJl81rDXzKtZWIw
FlWNcX1JxVtzHitT3SLYPw4CbXNuzmtik78pi45eXvs6F4cAZvs4RMyWRNOU
UAkVW9A3mcC5En+rwABpyJU1AZoXik050WNJOR//Z/md5DHWh7e6uOziYHvs
BsbWyXsTqx+0gMkMzKnJ2qDxThI+paAthnZEH2MXrImYo9H3uHQ7q8Y0yWgo
dPnB0hpplVMCd7uw6v7wOskAZSkyUNA3klXAvnT83wFLAytuMGeLobDT1QRu
FAh11wcN9OkedyEQWKsOK7+DbYJW9azRo1IRRp7/pCWuVgpFF+OoB2253Q3r
dljVU/4YzoEDfDQbCdiTP5UZ9/tn8smPa0rAyjlYGYqsCdKZV+yVUZEjMr4i
gN29hUS6AnHVQkHSAg182PVKrQHwFFpq92Z/GeybJ5y2EkewopP5MAkYtfbl
9dUL84k0SoAfHf18j6zFc8WTCRJvzEyg1QAquDN4qOsT+j/edS9h051AgqW4
OOEzR953pFlEP7pxY3uSpAPPtqpna8XppAZ0DWExRypdKd6M6cz8lreeBuCT
tXSDunvT2/CiTnhqW2Q8Lv94od7PEFleVDG4qQz10v+GQDf1HK57iYBPEH+c
snvj5Q+Ws3fej0bMYSmvKcyBy0KP/k5psIYgdrg/kw6Dh04qIbumdFfprMGS
1S9urdQxKhpXcqxrz8vyWLSOc+iZM7x4hUeGwZz8VkIWl36YzEoik49AtQJD
i3SsQQjNjav2ZmPB2OCuqe5uXXaoKIwsgIdZaW7gdwLvYOztJ1pZzXhtE6yP
5N0cqVYypslj03CZ9VeBImjBwnZ6IYIqNXHhZatg/3nUhY46De6RnDq6wch4
pAJWILDkaom6QT4Gpbs9GOG0Vs4suO6zm7FKo8+ETvRjGHNXEmsZo++Oefhq
RmAnmGIAh1HvX65/8AU8bOyfWM65/s6+RFVspnmfaMH5ur/+RHUn6ux8WT0x
65XzlQ56lT5e07QwuOLs4FxkHwVBk1OFWdaPKoXE4DV/2BZjMhfHVpLldDUQ
fYj0+y24S/gQo9kV+6jPlF3el9ULISDzGuHAnLGVtZyS1smEk3mk9W2tWop2
8fusWJ7T2MQE7XBGr/R15dj0mVGtJLDXw69ZC7QPVUgatUddq49nbbWRbBQ9
SqaQZc7+ZHsQ+qtfjMxnxPHAMoZce36qMMNLmVx2QEZUBLGGciDq2HTlBSxN
P41qmlNqxvDXhg7VrMmHcCsSb3CkcpLMvWzKiVIhE5NLAC7qhtuQaaZ8M00O
Jcjd2/gbiyBcCV3zSHgF+Xkw18UJFwyiHyzKYz4yZpy/zXkXwCKhgeiJHtUt
84XhHFtQTgHFyXcDdStrwjWsF6BKaRgwCvY062s+BXs1KWqvuoOqLo95eHdK
5exRqGftsEYqE6NK+1Toz7V2STBgmvtP+VeX2X6G7Bta8NmqF7UmYN3luBTc
hoTGEPFb3puimFTlhmkMq0sXFhSfXIQAalKAhUUSmDohHm/Ea589mTPyRAhX
pfMfEbzP+UlJ4iMm3b5WrXXj8FQkVvVY21EYOv9H0BwWhSwYaJNK+9ZmogAO
ZCuwCP30C6FjLsdu3H2kHKtijJgDbkQozjf9UOSBF6i02ngDvyJ3+m7+iptX
vVmpquhf6Wgpp1Wn75bRThjTKLikLz8UolWMSKyrXbVbZst3FCILEx7XAD4a
rCqtBeJpED7wRWRMEWyDabazW+nyxjNi8vIEKgSXaIM7vCN/4CW1VvllugOC
1cM0wG9c3bPHJBoojEVNQa1k0XDEcozGgnEEBVCuMhXWjjHBpDfrALvSSP8Q
3qZiRgYiroVSa5XDunbB/coyEhkjjNvUdXmKeCP6ucKLX7e7nSIra0QXyoEc
bdaH5/lSqXY+/G2gHXs1DxGpAXnfmDSxK1I6jni9Iu6JHDIWthc3PuTpL8KA
8dhFKWl9aMFR1FWMfWAunnMsjX6/SQqdzOaPwmZ2nUZE9YTXpaRfYFhYKxN1
ro34oEwyAQhzMGpWU08GDyDrfiAyBcH/R40aqAW7uE1ZX7Z5Uw192nBvQpMl
wTnGf8gtE+TBhzabFj1d/v+k6g77OdhiUMECfWr/88jby47UlsbAd6GfWXTw
DHFEuoBFbc58F7EfOby5DvDzpP4D5J9Sc+1GwYjrx8P/l6TMFdCKLSAwoD2c
SUiExMWMllViQmPkDMuMUryMjSWf7DI2hz9WOZMsWXI4GYaNSHZrNt1B7Znn
emQ2L4IrGUGZ39hurI5Dpnz8JvfD+pp8b+5GqK41I9/BtFESYzETbUAmeLJE
QZy9B4HzHYWJBFh38vMSBnavEpxFNlgDcEIQi5PWGfgdJLM5UrWsdV60V6g/
MhIk7VQqeO3GJyZ3p4156JtzIBXe/up3l1lQmUa+ErAEDZlfGRHzkS2sDJti
Rgt/UCMjgEyslnbdcheb6qCn8H/2EhFc1dzc3KOsNKtZYiz8Wcuau08gmb/0
HR3Ycih5YcpQLtEfs6kuPZtrQj2Bx37/ZHG+uzkwHndSvDpZVnuHUSjptNc2
Q6Cvr1Cdo2InKMN36+3ZOWRhw5pwANKW2qCiaLCi6ymx3U6xQJTt4DVL+/Me
oBhTSOIbdEbzShrEXqMQiDl9n1GcB9cLcCsDi40mVdPeG6TdXTl8tzydA42p
KfyOGBN2vBpwzzf4JJ3tJNpfUiiFZ1wfD8CGN2FZPUXyH3IM8MxaM3GiVMtJ
E4XrQ3+yb0S9ZRc3DW0KVxGmCxTHQQu7wTAX4XL9jvvzXFuczQG/0EvAJLts
x0vOsK/TVfYbi4cUZgI++vo5A5sk3tIwIUdVMCQKPTuKamKx2YMaSRZX36+Z
0OrgfGIfjzIOYzojCy4oZiUL2LLEwitb8E0lqXb1LCw7g3CUntZgeLa/IuIX
Rz0QMT0/ve/zixaK0/QDbFhOzAZ36He9VzgtTcqr4bMS7nF8DsJFcjCPHAzX
dKsCrDEJTuAc3UAk7a/oaezkyf6XtbF/IUsnrfLSirqjZAF5OZnwmBE27ZVH
P6RQHw1wf4SW4a0rh879YqPxcQTWTNYV1XM84ldK0u3zoTrvOboGzbRUlWAT
7P8l7vBWJ2EeaxmiVRaUh3N0VylgPGIMO0KKnmDIk/mnJy5uvWmFA86MwOb1
RssvUlXcTRJAdtiuLfzPFf+sPtP8b9nXwJJk7/arnIydKghhHVIGUM3BtzY9
2TyiNpfi57wnKXUvw4b8pnPOSEVPoZGv12QFRgHdoQEpeNo5k3KPSrt/5+sB
KfEu3Q1XaYSOGLHARsLlH50cwEOJjp99h3Gi+uLlVJJ3dNmTDILxbuJZLjPh
VYKB54VqBwwyRmdcJGEJ6D2uc9b/zf9HHhPVp9Zjnlgtdd+TCB4+qLKDp+4R
5zJ3z1DCvbiq3j+OFvJ94VqjPTQ/jWsw5h4GLfVYOkfwnA0Mv1lzF83LM+Dg
GRY93fBnd9xyqFilMi4dQPPxAkRB4HJmtwakz6Oz+81Q5KJCxmd0SsEpoIXD
XpLxeBkY7Hvk2DMEc6lsY/W+iElHh2sv61EMmL+2qo86BhRu2/8GYChMix/M
0fCR2mPAlKR37e7eZBDyzwm2Cds/IEaH2Lod7iYyiizseKE5iJLnuFO4p0EG
xNCj3V2TrPgX77WuqooReBBQieRFbrbURSnNoZWXPsHevQCimsmpptjDuFok
YMUonYuWs3NF5MQF4zDDWdaf4QO09pCYeN7MUfCgt7ID5NKD4OEmytyFYt3H
uXYuNVI5M4lxLXlKApUYK/76LpqAf0hfvvv6Dmfw+BWie+OiLMNgI26ErFIl
QsGDreXPsvukv9tbKb0e5NggkA5bIvzyOQp2o34o+8AW2XAnt4993EYUd3wp
FYKl+g8XfNUV6GjYgAjxKqgs9yCimhY4VMHVqNGdZKpsM47HwLRINnxaa0fb
0ECg6Fdg6qexLd7C28qVxNNBHOccZR+i3CxVp3q2NFjUFhBy1jc9cV0DF4b6
RcHJclXKU0yg1tcmvjAqlIfwWKFV5fafJuqhnwnpaCrL/UdVpWcUHahb9+fk
I+Y+Dx8xcPEkQqJAG+UiQi/9glLpc49ruvyg2NFnJ15DhKqzj9uyGCq/w2/q
oqvpzfKPcxlozUKPVJQcxkRdDqYNYEy6ob6gxWGJ0CoyL0btJEnKCJsYo+F3
Z1zCzmHLeNBWGfrfj20K3GcTeLujLsUD/xwCVHvDKRklHrP99JdX5qiorzZi
zPR0rXIdi8MfbDJNRU0evkq19k9yj+/SunodHASa4tW0e+DTx7aL+/K8Ox9i
4F8aKGQv8Q/m9nHUCJpe7dGyVXw8QAyVIRuFZgQPbmm5GSOXusws0RbcWtj5
hgXjmLvSmga8cNv2v5k2HbSMX1n2QBoz66VocDOBxca2Gq9RhJ+f5F7YEJz+
iXleJYb/4TlCtioopZt9TnrL+bH9LRg+ibyyVwPlpFW9J/+H3sWKMtZACMdc
sduLcOC1ChKFobWuklFQKNNHCKOA4jjuFVvH47mw3/ssytTa9EDGRGwgWJYQ
UbO/cydGjRZlNQyqbcCCMDW7Hv6mlXR5vJfojIGFNKm2xtUpg5IB92eFtL7l
pP8jYaimhmZBgrrgSs5GC6F68WPn7QzUIxfmTdOKOwHUlBGJcak5TdAdRfCs
yylNzUluXbqkQo8yLOsYLOdsf8hPQiQ4fHX+QFAPtqaHzY5vz3fqsXlyf276
wg/CJ+Kdh1HPOFIqjMYfZI+G+YNY2VQr+ipqb9uZEofzrLowIaIlJSqaoqO0
CuC2rkCqf4f1EJRcm8I2hr91Zl0Qv1xQl+JZvzk5mxHc/gyfKODtAjAWVftM
8EXvvjyexndrTLUok68Q1Lw+P40ZQDAPJ/4OktDMBU72UuV4pAE6/CldFNIj
XQrkP6nTvI0DIieP+rRtp0A593YpzsWUTj3oigDux3uDNCZ6CIldBJmCMLUT
5A4gqFIzJygcF4AvzzhS3+scYC6diucSLHuqRDJo51SWdvbu7MSDaKbnrBbA
5dC7bvHDotUE67S3SYoEmutbfKD4ryrdUIij/qykRwsnJsVmhxGASLAyq7uC
NK526r+wLnYxagrduqu8kv/p2JqKWkfZysESTjbvWnuRCk5iMRL4UmWpC9dV
V8GbLOyr0FR0yQ2JU0lTV+YzEC+oy9K77bCrte1fTYKNPVQnGYiI9TCcpRyf
aWHAJ/o9aiWgTbT/8y3pYE9BwaXDhTVQhAKOmQRBJ/fxsdFqm9biYobWlwIo
DmcGftFJ8vAcD0PSb3AAxFFnAlnlMV33nKrWTGYlpaOBURSb2dWkpfDwkipJ
ozjFclCyUc3QAtexigiXqiu6DnnyTuJWrmeCwvt4nCNd3aw6/syGaPMEpyqG
h+DgFgnD7c96hug8jX0QTYpv70cJvuTr8pYOGdRPy/FAyoBFfnJWeXQuv3Rj
U3vHoHrtM6uUsxSkJFX9vou9TiIPLkMUseGkPZmtavSu8bEb7btWMbU0ysA+
Kegsi9WDXj75fWXNlpaYKZ+8Bj7xkNKxhPA8GhXrAqZ+4ZsGtIqXNvyL12yn
nDHw30Knfoz7cqnxIXqVd6uT8FR+srL+xZvOFYrK9LfPesUSJD3Du1+Macg9
mK4SbfRPbupOfguNhidIDMxImmilnFikNKNMIkRIofSHBTo9YGcSPY+WFone
XZGS0pQ2m2cmtFOUFRuNnUSJECJ9GNCtbfSgZYReAX0wcWDYIXVoqsCYTDHO
YnwjYJjMfKMZqHdYFEwKETzzKMred9bg9ru9Klm1RmXlL+LCLywrc4Glq5k7
rPFl540ACy2z0M665WlJOqPYeV4ZRABlRTe62JWx6cGX3wGAyMFSy9BA7SXI
PhbT6+3Y2Ordc8C2KnalZwL8KSXUAS8YPZqC4sZu7OoR2tyOxVTLZQIlolx+
AedeD4kL7E2v06btCrXpLpqRH3RlY0xkOQKdSJ2j2G3w3JqO4FUzBHN3IBq9
Q89ct/iOp5fstBkNVFRnz/g9osyQO/MK2seylsk5tTM4zsO8yST90C/0lAA4
lL7NU2Agp5XmwCmpGFoKJbcXHJuwT12/IHB+jSN4Kqlg1HudnffgvFKj5jTk
LMqAtz15GeiLZm+WcGkr4NI6ncU0Tc6yNN/ijXmiigJcjuQGa/a3q9OssjZS
F2mptXU7DjJs6q2FomFm+0WQvIg6Hzdu64fuD5GzqfN0Vw9Cs+88HKzjMkez
UfJ2/6/8uXAzHFl6aSujj+JIzmKUDym13v5eMEZEj0jRflbvFGUEE4qs9iLN
wc9i6mbVdV1izSTgkrP1+0Adg4htToiis/W6FS1Xdx4jGjOr2Xib4uYTga/V
WlWsQpmc+3gisruoUsazJuMntVD23/9irkStnxoexgjxuxGK5q+ohakXUqRY
5asSBcFGP3B62AVXCURsl2+eOoR0h18dHoeLkPpOarUMySvMi9fwhWvBB3uE
GxwX6ON8eSD/dGD+c9ZdOD7dpLxTISD04R0v2Y4/D/Fag1GHQ0Jl01P5c1Rz
fpnyOgKJNhKsL3fvqme5wFKqSlZMTGpcVnRFFGSJbFHvEm8+i/ycXcR7/Hds
+MVnrVBMLaimYdCsNWXF4ozoGWXv6N2lf2qvH4o6e0A395I9AXDVGmWn+eqh
dhc+nKK5lpjeUMj3hq5VbF3EmA0hbO7x0pDL31TBlrX/Q+5dkEdwI/Ks/4Kv
+eSc1YugdQ0PjN8h+5lamyc436+Orq6G6BwJybnSKMopwmbXhrxErmnSwXPA
je4xHoTkbDLtbXcGiuXbCy1J8alm4xCd1tDqzDfS96KtVBlY7m6bqQtstI4b
9FWUzYnDoSrNw8ZF/ZGfsrYZOz8E5k0QG6R2bVHahH25HeiD1e67aWwxYhUk
w3Qx974Akdvu/Duvj6k5OZJbTzdmIPAkwwK2lroF+F0j9T+jAu9u8emTJ1lZ
eJPt6cM6zEgTLjjzCwohQvJA2VO/6GUF/3vqwvo82k6SwluUttcpVaGVFGiJ
rfO2cCs93Ghm8di+x0q11kKfgW8iVwCHp8D9b3nNL8Nut+InKW6ZGo7iHtNm
x+ZVdbs0m8ofGpU2VfAmyotdCvOG/irGLLVqJs9t9qK1Unz72FRMzSNLHO5k
IK6ewbT7QBlq8QDHuGybE3UoSfz7zONXRwQwy8nOOGzCY1P2yfCfHiGll1Wg
Lmn98Qm9CAOVuKpjRrLDvaNfu0ohLRHOuycynVLMrnwJ/R0sT+CBxjUzNLtF
a+aj28adOy1/9fU4oqr+yIOVEz1mb7CEJExs1luOjAYZUx7JpkdGuiUr1QcJ
uLyX7g0ZCfvv/qVFb4u0/L/sMmOikB4bMb8H37eI7cwwKxbseh8MWxNEHSOC
9g2Uyy6xHKfGOpCs+/+oGB8KZGjff/n5SIsGSIy+p/rVoa2/JW+0hGT1jLij
rfvVcGX/+NFhemwJ8CC+WjQuKPY1AdyAvI24+c0QH90d9iuflHYlqlksAFgx
+DyZ6NfgFHiApcoCrlEtGO7PJAgd1W6+1GQXcAKs4+7QjzWBHQRMmyOTXZ1d
sN3zDm17Zj2muiczF+COQxBOXJ2v+JdY5tffLNXxTE/psK3xwwWqDmMLUTDm
5j9VARM/2PLVf/A/aAKFAa6cNslZLEiiXf3C370GSCwTR1moAv7vmsOFs+mr
D/IZDNCVAF6uNEtYKOv60M/G5ObEfo0tLadHiVUg/vJrgo8wxqRFJsYKh9WG
bNqzAdvqwWF8Jqn64VtigRHrZ592Owwl/9oaWmzsNx08ndo0/bK0BssVUxoV
MH3vTyaOnqGe/8DxCcuJGleAymSTCBYKoI7csTS38VCqBE2u0oEuWLYVPpEz
XkvLiKmjerv8suJ2z4WrKierWR66NnNu1d4vt1bNsnpE3CLj1LN6t4Fhss6x
IbBqFZMQzIeWOi9cev4rFWhualkJuBZJJGCB0kcOf39f3UIwKKauhlaAdXOI
Dunn2YYFpETamGEvgJo6BjlRPewPDCcuoXgJ9uI/+Zg4PLkREwm63/4o4rry
uXa7mkUdfiornhS4BHuSqxy78P3nBM0m0WTLWlSUv3JVmloPT9J7g58sJhg0
FnB1faCUYl5w7A2TG+A8JliMhSCLLAeGTwYTPdbbWBYHCf8nVAuOekZepSen
MoBSt4X9j+wKe6C5cIx5XGt3BM6aYdJgNn4ndBJh+DQCjbsQDYoNkBeee8FZ
66S3W1Rsz2DA3e+bHi3ZG2kgAVMX7OQCuzM4xHo5re+FYqqRMCUCGxITC0i9
bvagbbkXy6YL7yijqKcW+ol3VyJREtzMl+dD8wGdV/KEOVAo+TSF2C31CRGa
HtAL4dgkGLF9nOMxo9FIoum87l82HCmqAdjSR/o0Uc5Dsjxyx7REUWJGR1K4
aKwpqHS7ImPueWq11LKMyF/G8zXcmD8MpIq3TC3x0YRPN/U0HHXmuusFRSEc
IvTISWT1rmZTI/AsQD9plpWefnQuEggkBW/2BkSuc07Y9Huz19qBC/ejcRvH
0Sxp8Z/e6UybULeBZwv8sVXyzneMvMfNNHtru5NuURXUGUQgXGIa6pX24c9V
jzXZoltT1oogwDeJyhqTAhEcrO4a9aOhCCYrUg457Kl46dDfYB43nd4LAZCd
dZ40DZGeyEWatCjJAI6fpMJoAad1KbvJLO4GUaQ8y+NzuAfjaOu6lxLsB2HH
zdMZk5Os3G216NeO4tIT4YF2bS54rq/eSYa4chSegvNnJSbXSjSZFwXFA3Lo
2Afcftyj8ikA/p/A7QwPtoLK3VtBVWTT6KG7Zjl8xsOb1PSGdREB5YCvdq8j
aLhlpe1P83QAAeEOY5qM7gmDNITkpkJZM5bAfr1ZRVaoh9BfDEh+aZp5h3YN
YeHIi6znvF7PEpQ+6SZwn02I60/Lv5sF0nfvh5RaNo/v9KG8WlF/FjPr/ImO
x7+MB2hrmAzBEUXvGW4iYnmYXvDMfWyrYYHfNdaB63A/MuoIhe/slgARxUqe
Sd1sxFEoWgU8E0DajWZxSkHBPOr3WeDhqdcWiQdLE0jPY46Evp4hnc699J59
/ZCkjmiG3XNN/88DxgQiO2ZYInbAHPVALNEhIDTUJDaP7Pou5gal4qbvs3sN
pBuNlC07dLjugi4HaIGKUS4Z90tcBRaTj5y3Z+Tzrevt/bTy0VOe/rLLNdB+
rOUKiad9dh+XPFNWQZgAnwhnBCAH+g7cIMsla78wOaUiqF2pnDF7Be318HE0
xoW2vGk52HcEyiE/FlgNz7Ljfg6SwhvJ37V87HH1SlCuW0ywgKDNjnJCORvj
vdMvENKN8JWbBQt51XxUsyBogbB/Ezju3dd8JcEjMh7Xx37AH9u1qkWTd32Q
zhhEXqLvd+q9bt0Ax4N9zh+rMkDe4P60s3Du8a4oN5rQmtjO9EHpRA/jT6qi
5vHqLvy2V2aGpD16oV6ZlNk2tQ7he19cmY78idepCX3ADTT3MTIr7HxYEglc
56lWiczFrzaSAJoe+51jnm+hV3huhH+2noKTi1poA2mW9mtn2CNlSDo8lwnR
4rjkeJ9nmh2qxevQ/6nU8QN06A5xh3trEYr9glltS1wzr0joQMHP5IJz5l5y
EyUOO1oIgf7pUZOR0Lo4WLq9KHkjJ3mmT2vJvUdZh3NKT+071v0nQ3qCRJOi
1/Ij3HUAZKWav8RGQl4ceULI1JNpAWOn7guK8PQ+UeLoYcnyYhrJiBj68mO/
QRctfUMK+Gx+4ZMARwhSMkNXab5cVUp2ZtlRikxlmbeLMDqyhulpstcCAhES
NoozrD6YHDb92oKdPcKc0wYPafgZ8IVvTkDEydrwuoaCEClCukaDvhk/28hj
I798cSjNiTa6eHa3flD/iNdYUJ1QQNMMqvHyNu7/le9UkaU7BtJj3jCOzynx
pFembIBk0ZtoFPVoYND3rP0aMGYeFGjSmSY8pm6hzbT4Fn//STw7CUDpa3vO
lb498cw8n6+dh7731lARbcWsu7zO2iXn8V+HmFhOnCG6xkjgzb/ADjXN6aJC
bljI9e8k6NLk5OrYl7PNWRIIL+YvgkFt1TUkgQH1oDTmhf8uUERN8RJ9e+uI
GkVKwwjEx6pxQfhHHYbY37U8UN7DnjKL11YWWX2usQmP6fMfoUeJJcgLWSig
5IQsNBS/ZSN0JOUqp+8y8fVglETl2E2WElu0rF5gtvSBmOELSM1FKki1Hseu
aEVDW5Oic9Br6KZK9NV7HZlqMFILkgU7YA1tlEWudi2l8sIPvCVTVUs6XrGQ
q6qS6S5Ik6zwCHtA4FY2Xp+VR7iPIBxDWX5FytV9+KZgClGro3oZmZ+tLbYK
C49W/YWJO/8g1PWv0Hbp4jnCkKUjaYL+K5498GQWUa0jm0meZmjUU4oAb2DO
Vj8gwL9kY77aanpKz+3Nqro8JZZJQpwAuMwEQ5wLlvMvOGqF+j5RLZFdEHUc
ScHdRDS/q6JG/lc8MRK5KsGcBJPfZk1v3bujqWiIBd4zPimS+aKB8ba4mwYp
F1+OIGUZVGGE1sd07/auv3r1aPVShUWXuZxXliAjKo8W+oOPt6DrlTatu0Nj
11Kb+Gv2xmMTYp1RKTlwJMcMWxZ0uqIGpuAgPF3D8sTF3nAcY0KhqKGFJ/Qg
8vo6xpTMnNZP/89Zfg8vY+yHudwoJhBhjtNhYkB3Q5pZRrCfPh5PRhIQUn9n
IZNHtBOqXrk/DqR5Kqb+8/pgWcGa30Is6jE85w4IRv3u0bXzOzn6RS3ahMO2
wyKgWJcXD7+TWJ60ZaHHTVR4S8MKdkfBNMWMi2Ojhv8HApfPo/yZbx8fqyfi
fUEelMkXdFzjPZIMbFlGmquhhPXioos/6H6U9KiqHvcZJ67E7B2+8ObpNFmX
/j/gT3TqBe7MBGLfXnEDxOz5E5JzJCsbVL9VvCGK3/10yrMkHBpYBM3rI9tS
rLmUnCLGEqmbt3jj09dxiCZGCECzEV71u6yQWFFky6OjS7lX6zYeqglcpHSK
Bnx9rTgNuoCj8oXfTSsEYxI9lBrbAgUy/hF9rJ37msfZDmM+pfBf6zAAiGJ1
xeIX0AfyUTRwgP8zv3ghdqCBJhHPQS6Ho0HPU78HQ8BnT2eyT7aTDt/+YYNA
Qn3tUFPRmGjF7OqVQ2xcC0CbPCHr1BpQSj94kqM+/au6LjwVwAVu15VcLOIP
VHxwRsZtWr85vpF3Qx+qgFfR2PuaDVR9Toh/1B09Sm/oATu5SB3wRPCx610D
+zEafsRCLKGVvJjmIKQunZ+HMJgewMDwGwTbnVIIZIdEgjdzLGuR0ETqUZJG
AE1QzGRkCj6uVEUtA5VMUT5t17Z8smAcjb0nKMWjmUkb39Ny5E/pfp4pbH+6
NwoowlJkk1e6+n+m+IbsxalqcM888hGBWpQjj2y9GPWZSqyt1Mxm7tDcK6Jq
crX2/flrajC9cx80VRCcOst6MubMCJkbI1Im9wD8yuPfENadPSN/hA5Fr7Nj
7SX3ArFH7AirWVkXZGZYdlh++uAunq8X2Sy1gPHTELPJXvDMvFpy6RBArBWh
IGERVUpK7LDfGR6W6idXtETw8Fyopt4avBxqlUKWFXaLjt6Ygbgmp/b4p2W5
DNuRsxgc/ynCibuAsNtDcfzN/WVGv385Ts+bzD6M0GeQ0T37sGC7So8EKy8K
RmY3L4w6myBDeaoZIeTP5Tk9NSX2iNhDW7Ppwsc4/heK78VLWcu39WkSbPtJ
koIL7Ze0r3TKtEu5OyVJlUgdXgx6hNaxMCpAukAEJsfLseQJffpzk21tsAla
e0nJTdW87bJEoa9vT638wmCsXnngxjEWh9fXAchKubzJBM+6RrfUojfTuZFK
/uMXcMqVc1q4n1HtGLcvo4HEt8OZuH8NJZHPaGnu7a+yLkBzyZnj+1WWjsT5
0+6iFEsjrRfmsPeCIsBVOHajPQVYPIaqBuASMI4FgUxbHB855Fm4S+zWl3cH
tJH36Yyd25R2p/L/uojUyP2z0qyay+5zyscFdXLWefJh/hONxWheZXgH1pDN
A3wAs3/yHEnYdLXXfCIJ9qndXy0WwFg4bE91lLKMrSuzAlt5x2lQOjuaiS1v
+wZJNmw7FYJ28BqAPRC7S4Yk3k0V8ZHwQYuZgFvNWcXVpNm6SEFQWqCaFeKV
7GsOyS7YkL63uA8xeMFPGZueE9nfn/7yYIFUv3CYj0WxuPP3gTvlDDT4n/Mw
bNs3+ZUZdAaaKzxRMOrSKfYzRSwsnVOWCyA/5XU56zVHAMRU16+nNs+pzy0Z
CBMeg2nSuqi3usY9Wuwcvp7qbAvefqMnaEQ/tJkSZtIHdbWdeyckyqC4VB5n
Utr/NjN36MOoBzcFLP1x6aG4A1ycwgzjCtln/aNlS1mX9Tw5D4HXn9E4mbBl
n4GbGc1nhdmD0f5tPYtn9qS2DVw6p3VCjPugRnBB3yAjt4R8xIbVg91KBFp8
UPsujXndYfewMwcrAZOPKpXksAOzHJnoXC8onVgYZD2H1YgoCkx2A/WH8ElY
mriItd765FQbcfEQHI0z6fCAGwHwwUV3e1vGOOj0ocrOQ5WKLOp4avB8xc99
5e+m7lqp+9S9T1aHuHO83bfSXrrM+Bo7U1ep/OU3qWldC3eakckXxx0vfsBn
WYeyTkM9g2RV/fdYE5YYymmBvUyPoM7xDYzdyMVGm7Wgyk0hzn3TawbDFm1a
A6kp3nJSPtKxkjYzkerjIgut6V7KhqUzalEEPW7EA+7UualvEh3SnLuSVf1Q
tnFoHeht55CJKXGcAhV+M3X5eWpvF5kWGggBkthQGs9z/PkTGolvn2hI3elH
IGEe55yk/PQoa/C4QQUQXkRfJvBEGVvkXQVDkAgusd+wmgKr3c2UIrATJgvY
Ni91Oq6ZuyVEfWmoYGsL5c4K5nUMyUpKbW9v0YI855Sy668XnrsTjEW+A9jf
ZDGB8JPO7sJp1F5eRo6sisQeD3dqFEG3fI+4LzDm9uioOWDvqr1hmSWiQ+Ql
awyii+Eweuro8gco1zkKPzsxBxSQpBgAy2bfGcyDW2hnPlYBXiuJ93pGXT6a
ENvJTQForYMGOvDlXkYD/VLZEae3SIvEKURWJjEgvQdTvZ56g4nAxdsmFovQ
SFHfCnF2WPvLN6okjAPOuzsyB0z3M9x6Vk4C7Yfunz3jsgATF8uxhHp5rByn
v1T03b6ZwtRTG7KjX1sEFUIgtoxrAyTvo0twZOVPsjGmlgU/3RPc2KZ3INTe
SidV4mZEXldL4BmVgWphgcfORTcdX/8yFbCI/sdWV2g0P5nnReeJRg+8NLwZ
ZHuWW+LzDNEEVJqEmdY7bwndcxWh0vzib72L01IZdFg4ZzQH9eHa12VMat3A
s3xpOg92orows8YrZXKnwMlxMaQoi/L4DZE5lL4qL3Yd9lMNzeNWjpRo9D1h
i6FOrmhqcR2oVo2RwFNZfW2Snc2aJnXzZM6JnTWhC5wkJNkjGe+cmIutIj5O
KZkibJg6oHlJPF64YfnHPGJ6u9XTC8R/OyDiILz+NwR9qk/suVjXIFdtorNg
pj82lyvak5K3yGnnf0dmNT97m/RnmO2xbqYlYlvYSN7RH/Tu4SH5HVojTinu
m2NVTrPsfbnd/iLTbo3fERVDK0fIOk89plTzISsNd4xSW10XFMFDjeAruvKb
843jjYJUn/hFvs6mPOafiIcYy7lIHJUaDqL97BkVew96a8T3+ptBIZt8sTVA
TKs7viVWLWC2l+8vAzwUnTBPeaosisuiX0FbALkn5w5QpB3ZcHK9DeeMFAbh
I6QRrLBnR2MQ4ZV8wr62eibWOYNfZdH/Q4J9/fTVEN3fCQ5l8CtrUSvlYT0F
V42xuOAxnn8c2Mz1sFZrDKaJMWlTWN953SJ84i685vUla4uBNyv3COHZW1bb
15uAjupsExDxo6vyU5MAoOquxZaKXlchWdI9mu39lE+yGE0wncvmTaeZcLls
sEh2rR9q1TV3jv9yjMNoPD90NqcmqYgAXh94JgMSUsWjMZ5YkPJoDjFdU2Dn
rnuZze/K8vERDzcDoIwzjnKRGwSJhwCk6VH0TXqRZdfHlpFD0fT5xSUELaK7
R4wpsd4U7utGbZMmVx1vv2/e2GJyeeIIB3EpAPD+ddSBNcQeAC1KIQeQCfW2
RESA0/5pHeVuo1XW3p2g7KpAz8f8ORyihTZxD+BcGnKc/OCL671BWoDf+RVT
Tp7iAcwQ6oUis8ZU7VEQS+p/4aaWAXeZhkTyMhZ+cVELqqfEU8E12bEDxFSn
WHz5Pmym8nUNj5gjB4kJ3hlTw7ZwrCK37bpzZ8WOOruWcr97DLV1mfhV+mRZ
qQKK+G7p7U9+OovHHHXgabgbVxkxDT2kIbEOZSuPSaMuYfXPNrf14mmBk4ki
0WmsBY3p3FCnbHTbifK5gXOkB90nba/HbtNyTk+OYcknpLwySytkrnjhmEoO
5GYBeJTuGD3XEFcUQn8GRswRCBC8mB7qINcdg1a/zDxbaptOOyBmoyePm9fS
7Y0X7cVIX3sTuL1So9JVUB8NlnIg0If2zAbyAxu+3o238EKauxKw90nFmZFs
OVDKs9DSj1dQ7RhU4BsgKHqtYgUZc68PmGfFjJe9FrJqPdYseoUWcxhUuvbh
kNIno7U2LEvW31WLOd3BDETnpX2+yWIqCYL61Ypg3byJNRPnRYnoXB5bNVpf
uYV9tZPcl9B9woe1RacawqhqhKsOa22n29EepsYQkQ7sVelm62tGySoxL7ZX
ELU2C/aaBCUKtiYxcP93jy0wXLZqtKBKXCIe8JsJxVj/4CJjomXb6m+uLxxE
66o76VJ9O6qjAZfKlukguSZjHTiaR0p/DDmMCvvj1p517faS5l9Mi+Jl6PAo
x4QAh+/qqGwJ/6rXmmwElrhwuJkU3pFrmtwCP7EVnpePjVk3gqQuj9taOkaO
azrLUi5usDL6LgnP8V7zzhsd9nHrmK2DPzoZ2WpXUIJI1mE1q27j5eeeWOiN
37ZghSIID+lGFY3kABbR2DnoM5ZvX6aAoavqFSro8Yx0Qmkzbgf/YIZm0nbA
EMw2KtRwEDk1xY/NILRwMe5WDR+opyOIm7NRA9XIdfrL4tziySzz6NS3LFKj
etUB93JjzsW1fnVOPknAayPgmuxTOlYIofvxl434rdzTIB434PCi77aKmRaY
D+KnYWZBsya8eIwrjh8ZHlD7aLIX6zgN8ejRtNizfM4DPOV2

`pragma protect end_protected
