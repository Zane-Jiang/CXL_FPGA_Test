// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
j3quCyvnvdEN6QqCoJgCeopNJbMi6UN0QlbhqtVjWBnEw9n0HOyH/cXZNUfYJsTj
US0MAYGJA0dYRzNcG0t9+I6v0bwSN495qa8cCzRFgTHCgGmCFXmQuS46rxDB9g9w
jj6bOBBIcN/jboMGIAVNKydlY/r/Ow0DcUbdrlN4y0aOzqvMpDZLWQ==
//pragma protect end_key_block
//pragma protect digest_block
T56Rjq8Mi70cl9/1a/lQkuL94+c=
//pragma protect end_digest_block
//pragma protect data_block
fAjmwUjkNLoU4cz4xiCVgaYNgEQLWremup3z98uIf1BbmIOZ2Vjy/mE62wOTgLeU
UjLTtLwIC+0Tu/LMtgI/WFiIwICYWkVtYq7SmqRKLThKmud7apCb2POF/WQZ1M6x
C4Ez0kwJmotlDUrJusTUvPaeVuoqpPqLiN1IeGZJ4Pw7UIxK9fEEpD0zMKGuYQ3v
OqyIrEyl2qVmWUK20M3WDNSDcHItIvHoj9ovhIiMD2ychbCgiX9SO2+keM1CXLHw
ibOU3U1XA/WdXj8e4dYeaJbZOfSDBQEh4X+vR7OpQBi3aITfloX/+a4CuMzhwact
/kkmcWLTOavY0tw86/tNSp0MJrje5s0+HdigMRmCRPju4sptm3wUN6QhVpCae2Qk
N10qRvbUjkcUvz+TSKNlExG40SKeYs4Yz0gfzMQiWKcVgaLd35nnY5jDeJikpmau
t6jqGzejF/ohMViG1JEGLqhyWkEArtORCyeJbgwKxb5hmNIRZEwnezMAveppk+2t
UROA37f1aBNOs0JL3fMU5O5Bl82YDEneQUDH0Ksf4B2QaepIeilGArb5OjlKpHU+
yHKd5jmN0TLsmxPHFSy2JQYA75rTWMDurPEedMhnFXxRElEyWPL9RTTF8OB2OjZp
NM1cOhX98dadoF92DCmUkyD17OpfVYixCd80PYJn6HjHzCQ05/RI1/CVL73A6Rm0
UgVfhc20XC7XU1X+7RBoULaT/bSNKip1RTI4z8f3HhCMliz1WwjAq8vQqwcHs8uM
kdsLu+lzetYVyd6E+EBSahGxNIdb0wj0uzu2W3ylLz8B4kAAovNeH+SH22pUQ5ou
BQJD0J5qLAc/VG9QHhSd1G17Ce0yBAtlZ69roOspqunQxlP4poj0RcPlvNL2vDOE
HZWyjV/cSAGDSggL1CrdrbbX2gxUXk+FXy7JDW4gaNDi3E+oB/28DjusG0X4PV4x
RFmhSk51XsibtU4BeKLFghr1poUTeI0g58m9egncXQuo8zowYFdYg6NJUyBebijQ
4AtDRyzM7Pj3g9FoOwlOLBQYI3TqjW/bZOIm0s9ZDH09ct5s3iJLA6STujEmeYNi
wAC9XHpTm8E6jfp/5dmQHaO6Em+T5eA7qmlX9UO83JL3GKN5gpPTqApDi4qXij8R
+WKHO41AnEBhmkE0WtVBLtjVFuCW/yU3fwhehaUUcS2Psy87TvuTUS+lpCh0ahHS
qzDM3J3gNWUnwZLhYJWBptfNbGKlN8Js+dq/WdmVkS/J+vzxba2Ras8PROnFiHVz
fLBj2QO+joPOgg4VsId+fnqfE4ZmRSI1HvAvECKQtTK+s8mAF3+faod4OEDH+8//
750zl6KHMCXHL+/JygMfs/rNnReFcmXLSMddpSiSDurtLtKDt9vIbQHIOexV09Tm
ZaOvLrZElRvFAwOhQpv1PjK7Wb39vl+dSZZwB9G0Bo9UBWiL48UZdIvUQs859jct
3iLA9MxTQs7ra4iZgUhc0ZnLQARApywuntcEdZ9HNoWz0Or6ZoNEJU9kuUXgJepY
cKa90chW0+wr8mT7cd+T/GcnlClJtPlfQQDj3d3fl4gpw3kmICkinvlt4rNrVitp
6aBFRgLS0Ftb/yW3N910JxE96NXDcYg2OQWWGME0haE5ZRqBJluzgPlUeFHNO54u
CjhhDJtrNsES2fASTmvn6cKbRj6x9dfBwweisb+k5rk9emXQFajgwLu8vwn/EMzL
bvugxQ55PWcu2QDYUc3oW1XbHtTVw7YKjKjz25RCeTi9K003C0OSqKiyqzfhuxcp
Uu85bNkqM2aiCChi1zbXrxNVsw7LmKAPsEIwZouYRjVuWcrbPsFJ1zthrN1JNn/S
WeqblFuJobr2w37bWJuqDPEVR2kDpYXX+DEVUxX/xt0mMTc1Ui7sejmnUKW0Zh9t
uZKFx4rcOMnnOuTRoxz0zu5tr01RsafMpbnqMTX1qdBjlv+m8B1XY0RdlZ+RjZJG
lZ4fd863soK4ZIXGJnsatITUPNDkV2cjjk7MzHNdC4cDulvJeuOmHS4hnqqp+CJ9
JD3Zdp3dVGFB5ZSw2nIvtsneu4PaPLBlvfhBq2GemP3uDEUdxgTnTEPvjQu1kzWM
+dU6SILfGu6biO7dW+fu3sHYz6JivzP30ndEO/egb34fKDmmCQ2/9NIi2ClHfrx0
ob/c+UuXDVW6HXE0Lcm2N2U+gQV6CgCCeFJuPE5EeIATOQE3TXQk1P3TP74OZrOG
R5SCWoqdPMVyUYJC8UD6WT1RP5r6LLW0+8eQYxq9iMKhdtx6dpO2wwp6Xmp+p7B0
rEjnvwtONXkKW4uWvMyUqvfAUI1PYhCaYXZCQlffEjTrvH6Wfa6deZpDixlBAQx/
PiofoRf0zfrBVkVGHV7HKeL67hTmXnbqUSNHrJAVrWc8Kjb3QBGbL069DSugNiF3
vK+9RLdxw3QdndNfRha9d7Qvhs7X+KLtogHRBhnSA4YKM+1D79bE1LbWuwQlZ85g
p+e36RbtMMHIIC8D78+ETLgxLAH3TeMPCJd+bWMKfRH390gh1Ifx9S7t+XyNvhHQ
3jfJZFNJh5eVpbxo2Zbe9pA0Owxxe3PTy0Z8CPX5otVwFQNbHjQU6bRlZyViPdvC
K6eSZvFfeeDo8+wmZkjozTqqYsJKfabuPiDEAnqvEa0UxmROHIVWhd1Y0rNWfe9P
vTzOwBvDacqAdYQlTzpnBI29WBp5YYZ5bD3xtZO22oG8zoJXy+I7LnKxIRqftJIK
UGYsl1Us/C6MFXMRfdQEcb1t9PzAw/zchGpAzYVatGtEUmOMSVQ7EgBc5biFrAS6
ziSCBtPb21/++fXQwPxRDA7qxm0OZiSD3N8hhYUTuUTdhw1EYRx/VUYnaZZRKa3Z
Vz1ejNzljqS52y5c+BxDRM2gzmXS0bZoGK0GtLYAPLYvAgggI758QAUDbSluEdwu
ltO9jcB669D3r3Wz/ZADKDOug43ivgVYz3mIVNWMkO/ApEZ/CrRrjvpqztDXUwqo
5BzTU+k1+t4aTXe4QU3Zu8XuzhSXlkSrbPxPzwfB9y/sh7jUErIfbFyNGgVnY6Bn
mqvQu9HkrOjoQYDbt0EhzSF4V/OGZKBU/q/12XIi9T6d/W2vuNQpshUfqKMzoj9a
Ag0Qsh3cCjVAuwpStBdzro0d1d+TJnE55Yac9Jow2Tv+2UohmAqQuk4OjZSatsyN
QQndfnqL9VZUdYW8KZBBsB8srAmCV2LwtFQTHzV1FzP9ENF2zgAVzGPEZJbbykat
t/b03xRw+rW8F7uDDzpFnqyXizUDdWoLRmXvZX7oWBb7I1NizMb1jxvceLw429iC
XDLTlPOCVl0SpTl061lyLyjSu3ekz8Tlm0zluhoiQkc/jALNtt5bXNjumhRJnP+8
nIrpZJgCND/LgJpb0kaUBKdqaxQosw6Esj1BdUpIN+L+bqFu39zWEGkncnk0aeYE
RskEaOa22+6zc3dNzOOhKFxK+PVY0pA64fTK1LLViVAnN8DNlC8FH7SFqLiJxmr+
i5v8hrwmnGMBnTDezyc6QKMbFjICIjKy/VUXwMp0ncN3cSGXi1PeFQsLpNxUc33W
lzJdnHpMMFhJV+93jnS/zqkWvyfp/wFkmYlJV8C+YpUL1us2NTWk4S4sVzSPgO2w
ilDEsDugUrZOd1VwGeul0SpHQEkYRy50H9IOAvDJ4Q7CJa0kSilNHIjGiQmZJLSf
XJQvxXd/p7gFGlpFGFb0EsYIWH/TqDff4HRBnEEzelNtcjL9Zs9z7FR774ZZhkMt
PY9IFBYrlY2RkrqWIYj8Tqg3DnnjMWX512ZGjSLim3bn6iOgS0uurydHeHdYyZ1t
OS9gAp51BLMYQmc0H3fp5orgxI3aizJQf7mHKHJ5MI9/FuSqAhIlJ+cH8tutm0q1
eoz5/dg1kPQgia8e/m2OZvxB3tD6uZR3dJeiGvavVX204sNgiS+o6LxPFRyifV/3
e3x8sxiYQZk682QBj3wbjRhNgtn9gfA7E4MYO5h8wRwNw9ogZ9JWhQsbtlgKUG0i
NNskxiwZknqJplHqAr4xbIacUrPhlRDEXbPtGb5Z097pBoi33FdrYp4KnJ+JfUKo
3c+L0hIjWRkrl1hY4ddQeyEnXE/bXqXLPovf8OsY75yzGF+/GDMG3nfkerUPOKka
DXy/HpCkzXj834KLqmOoQ0ONKW/mg31g66ynM2P61kJ3moy9uHe8N3Gd2J3qrVIT
mb/1z2nF42iMs9afNMYtlJLnqo1Kmr9J1suylo7ZqW5T/spAZZ3D4F/U13B7qyCb
VdTVrFXg8IKMxxFn2lEgucfGrXPmymayD/1iauEvtAEMLMamPx8BoymrbN8bMDPk
bt8duWf/5FakB33TW3LfiTQFCRCqQuz/tq6anvX/cPZuwZbupdVmUbm3uvQr0lxw
3BbH2eR6GeY36Lf8Izug/98TXKKufHKGuX9sTKjqcrO75kfj7Q4n1/wZqwQri8Kd
8O04I36Tt+6EElCfPG8EwMkRawACCxlyFKtchzWXDWfu0d0NtrJ5eveUYAnhg0WY
MMYXSFVRlvUK1ZD1AUgAQzdb95cRXoh5R8RJ4FCT/0wEzGm/U3+GG/V4T7gW2WTE
r93Ai8KwxXX59CTcyEynr9wXVdOhpsEuUNm/OlSf4OVUK+X0ShZ56dGwBbAfhQLv
pAOfBliKoBdslLILKoGEQKGf38/xvzDEj5dmgUwI1ZGjL1+aGfg1oWUER4vi4haR
PrpZzGgO2E+UwWsUQ3L9MOQanAFOTTo3yoa/qOJjffrYFAfAlOWCg+vLr4Kuqzhw
21t/Y9Pn2zzhqs/iTF+25liDX9ElPE9iiDn7UO0Omm51ADgJeKA4KqudA1tC619D
m/Am10z6Ko6NzotQk/we7fnwYDxnuXkUk6c9Ohi8mtbFFX93P2c3lNajsU1YW7la
VWN/1J6+k4kh+pdn5cIo6TDrCunzvr9Wockb5bgQUmX8TW6bmCy5OA/gxve+Ezx/
EDYV0suL9yTdjgz/igBWR/yku3HIMeN2fb2EJWEXTY52AM9mlZTGGdIn6y05J/1L
zM2oPqTC89qBpTFM07joOGQk/ntSx2THd1pgDe+oBCdYSUjOCr5Lpl4Jf4Bo9VUm
da8+hjbGMeyzKQUiR0fM8AQewPCzICbzHg+z/yB92kZ9/fiQo9tM312l3lTCcEYH
xqsBeKu+7bBt3qb2tgLf6vtpxzPdDcirtXNnggmz+8mIjNZPFcE+spOC29QWfp0Y
LK/59wAOSFKXGRylfSE0q70RG8gHQpM4+wecvIbgLtaANHwjN47+HG0OZI0q+btg
MYr/1cDM4M9ZWdlTwugRj7fMMyk4Q0BjXDV8dkRrhch6fZzAPO2E+iBeQiHYjpoA
qkIP68yc+IUis/Kn9wjxLlIQMT7eDz2ZcUAaS32bRiIlfBf4jJjPMFi+DdcU2bDs
Ny0f5byPTpBMPJWDwwrL5Qu+xCThDAm9Bj1eOvFA0W88f0+cs2LZaVM3Joc9LlJ/
a5MnPwepuGMh8Il530h5nj3YhQgu/OF+zWyvFbhu3dw/MOLrQzkS27s9OuNjb+N/
tFSCkZFmZVVdn+bQYnMZSLPvvmsBX5g3QmPJWjhZivF1AkgJLJwQmX3O34GSagqA
PHmlrmDJi2h54BuwmzYvrP7lVtmftQ5vrx+Q/pm5qZObgLx+96lNhK7SLzVJ0D/j
C0OIXbduEqTCWmvBoMDPFxLLX71Gw597oUOb2QG5d1VCRWJgYFkNbzdeqbLVwYej
MylOIM4s6vwkhCb6BHtmZxRuuVO0p0SqRG1y6jfZZoD1MGLpLp34OIlGxCLzFH7i
2x9o7RNREMMePWcru1lVg3EL5hWo1oFnNILlkPGlc6KuVjBPPerJycrAGme/WqEb
j3DVwAdAKau24MzuFM8EzYsh+hy5JuiSOEFARUiSb8xCRSYKRhU7UzI4D9AzhmS1
fBgLOEMUkAIPZucPBY5gdPrUys8LXxvVTPMO8hK/lCOtU+TvvSk85Qb3muuYSzWM
NdeU4X9PrKvUZPpHRT+pkv2iNoatBzX5OjhWQ3hwAqoOZHaVWYs/ousJTijSABKt
yPOJtCfzqs9Xi/8Ejnt8+fFvlcL72RU8rWK0fqXbz6YEz8mbYJWDAElwmB0d1A47
rhotIP4UlgPjs2shIF2IvmG1NIHn/H0hdvQRjjPdWGT0cbej72WpPKmfZuVP8BhY
YrbAV+qeUguuyMoxJhjyWzlAfwje0bzVmsxMTyW1ay7gPBHsYvYgYSwGIBRVzBkL
0ni1KQhYAkN9n7Z5ymxxCpFeK9q5AWWpNJlKnYhS8MqXIladewZp4LHjz6Br6tHx
vEX+mjxPJ4vsmhsz7Q9R4oysPOc/QFkyYrc+T2ZQG1M61B844X+Katfl3CeoOfVa
QDhBpLrfadUOG5hnkgJdShl1xnX4RnkoBqf/cOTSLQ3gC1iM7S3M8NydPPxR6YXe
xcGiI3+zkIKjlA5L5NFBtjCC2HG9Q8oG2vLIewZRKu5NTauy5pSYjlPAhgG471Pg
akhQ+aUBN25FlkYWbizSmIMV7xVNmi763cOP9cMvrC6KjGfMIHCB0WBW/NI0iKoI
nX/+zO4I4yK9VcGpQsOJwsai4taum2qSBzasFYCC5UXmHlNCcr1Maq8AilYC+5aj
kKVqVpNKHCPlithdkg/HY2Cc0mD0abZIiT2KISbz9asFOpxt2XVIgtQmqfjx3/yx
Eu/qiusUXazsQMlHyvsYlnacwvbsVC4nM77C2N7pfQTAR5cy2UEpQyj2PwJ16fGP
Wknli7H0CxaKxEGjlCV1UDksfgGFgsR9yPupNViiUSda2rgOcXist87nYqI3ToWD
9exh2zHSDqmZURs3Jp/iNP6QvMaJN0ollWD9Wy+wyqJ3uj8gV/st53rpM+yCNpfP
tW6G0C19Wns1/N7l6chtQfxXjfSPAFz+YqwZQlcYPnrH0x9re0T4622TY0RBK/2f
2tptJtChpoovdswLWJuJtY3WUJ9jtdqO3onA1Ur4bwdrFDY84Rr0KU9Y0CjTAasq
AS/paHQ3mBg4AYRIw30968V/KZWpSu0GSwiGB4sc7M+7XmYFqWoJRmAcDUTMai09
42mRK6WBC6MOhel3LSqVjJ+SnXiAJbydzNddbWjZFL+7PXSGHO3DNUVcSy9dTqFz
W7zbm4VxLXkGmcc6lsU0eUSZttAUyaYbACXWTrUBT6425IQStSCdvn2skxp1k4pZ
43L4QKN9GwekLTvq+fLrbWtFegDQObw1z5g7Ub7pKDbkGYbk1La0TmUufmNg5iYt
cRJLu4UYD7KYgO2J4Bib0kHjAz2emnylayqWJ4FJ2l6n2NyYz7G3lGmFA7ppqleB
5YEfBLupI8DS6i1xyAw/OoWe+dLr/MmDlCqZIMwjrJH8u+QSiNkr0Y4uqoxG/K4k
BdmB13oevANKrSvJZJXWskA317YSey1tN3ndahFbuPsjXKBjYUTn/HsNeL42MVUM
mNu7AGtaLNj6K1xPpT62wpsuh9AFbTytnPER0cC1hPVL6yNv0C0uevXJYLFpYhT9
J6PhfXdXDmK4aR12l6EYpIL5Sw3qVdl0OhxFPgGaAmaT1EwNZ5c8OahZf4xodKJF
dD0t0zwSY7dH5aqy5Ko++sx0cM7ZwFt8AozDijjMHKz3lvbRjsZS0+GN5wQNaItv
quGpk+BFreYlyfSLKS9yj+Z2QwXKMG21M3q9nnJl6cuDY3RdOMRJhE83VpPwj7qa
zKtuTOAEcL+bF47xfMvj/sa4zWtjRh/aoDxwHQFX94Bb7PgY61zXF8VadI8CkdoV
BRE0Z5pNWlCmQMonEqGu585MEhck6WU52y95W8DWHfZa+Q3JezTH1p75KKY9raj0
ePH2Ekn1Agg52Hb5kFrWoVYPOfg9Ei8xfsRHR/i05FORLCRviX/z8J1sxvWmAfYn
Vx1fP9V35VtaX7evedMvHSIta+2o9c24bTvpvF0JaAfmwMGUWJpm7HaQVVWimCcG
6fEg20oWOrrSYS/OOzQuoI/tfudeJ7j28R3660+cUJcPyQHeavPINDAEhBOntijt
JNxpQKeTnW5LR4zlHPAkFNWE17Pz96E+63ogLTWsCckU+9RTtAVl7Ba/WkkR81T3
gr2nNz13dgFcIRfG2MNuloYbEWJKPQ6BEIGSmVZKHmg7dmCHr4fqmPRH90HO0vW9
PdK59HSGYxmq1mDl4OuhadB2wpAZItwC7xekYZLTEN2Xbx6EkznWaMaRVOLMQdR3
F/Y4siGFmiI/DZsOCsRvkQyDaZzd3bmOxh9QzsnDaa57o6V5F+UV+eiPTZeuFW66
1ezuzjTSm4YEtHOf/Q2+jfcOsispBAIb2Sv4wBTw6XLdVSsh9RA5cx4IllmeMuWu
SADtywaCtZpiQfNFUBYvonuWDustEvbGLAR9tMu2M1WidLPZxs38jaTnR98vsGSl
eMNcGNeOW/4jEwKVr9jIMH9XdqwKi4w3Or337bS94eMHCWfFdaQ/mfzMdqAjFynl
so6wDHfEiAnPVYLxfA1YPGTZoLoH+SlE7ZxeW1G0Sl1gD/39AIu/9UFpzyG4lfWo
g4TfMMvk3k8MuGeuPYlCplE4h0MBR3vnkAxCWGyjXt0nSdIbexOQDYJc53s8ow+v
0YdcVTdHUxngYUv1RS09orWM3A9Q5FU9mjp0XAEhCrROxVC5VmrM//YmpMpyXQKh
ZZKMCdIISYP47suKoSiB5tVcHDOHDdlwfmN3StaahyTW100HLZJmkhnBApw3D99/
BzNEnw6XGhckC45CeofTX1Z9w0+jkGp2zh8lOg7UPFdPW6d9nF8Si6M2gx9+XB5g
h6+vOpJWh6QJGuORBM7KcQF6U0wEwVdIAvdy/iHeQ8knF5m7NMw6TE8QBTjv11If
YAosJstQSEiZ2loYhQIxLECLQwRiHsxZmhCduu5utQ048WcOLz+52B+Qy4YV5OAI
NiaCJ3jnoHuNI8/baIG6nEzjVnpuhMTuXMe/DyTM8SOQ4sgpzh4R/cstoCgM+0gu
5OgX5FUeSWKenOadTzxQ1uzm4g5+gcujRTpS71sTQt5FLYDNUFpBkhLNDNqskVkI
MSludacPFMgogwDy6hG7gpMV22w7o2TUsXN5JgzuIdVk9XkGKgqDljJZ+p9IkQ99
ZsYAkKWqlYAzb+dIKyZ+D53LzrQ3yD7QaqDxLWAhxhaOQyN4E9tQZxxPTbfPsdaC
lEmmqwY0wBCU5lJBElFuQApennKeTUBOwmzCqu0mea0CDFCkjS4tkkNxY8ek1DVB
RU7/05Qc3wBuxPh3K7vUgM0TNUzGvSJdhdGzkqFtUO1mVYDKE5PCBIvfmzLDlcEC
FkomeSFvlEV5hUSO2GfnczbDEKa2q905FUfLl4AZOgMfl7TSw8IKV2OdM//64Eqa
9GTs6uQkohwK2wcrGu+chtslplDfENbCnGfSbH/82vN7WQSGEUqGq5iDTxgv5oe5
SRC4K7+ITkjcr+14QgIdq3ggeNEgTbTlZgRLTS2dSxhILXlsT/Fezn1nbpmWm6eL
lAh817riYqlBbom9BQDNEEGELTW8uAnJ7HJWZmGagf4FkTIMNwznJELwJrUkswEB
BP5QneicTLh3/0g+jpF72CgVSvmimA1isDvFZQWQAZSze53NviuvdpyUlrqmeMyV
gcf3yp6DVN+r9WF/V3xmr35PRyB9DytsWLk85zGCbHJqMRjHSRsigCm+gujvgF4l
0ucXkhaVCACDx3RWuK/xdsm/glAuGC5JjdkPN+RYEhLIDqqzgq6EvErApKO5ksgk
8qf3l++g2tYv7e24skgafAM8k50RRRQi9DniEmuP/nxoM7xwsLrRBl5kHsGCzSBF
6nNAlVncSftv43tijxeyZTGZD6jXEMg4j00YpGACrr1+3BAdKUyyBNpOpMdN42dP
iU3lCbYO0pS0ifjZuSdk9OivtxiiTe4R0dE0Ja04ipUPh7mNX9jzZ+2Y2t0/Sydv
Zo043S5cVQSztvSibMckKEa369dA85iW5BdSwxTnfAyr9lzJPKKwB1H1iyTtPf1N
ZEaa7PxUa4P1RDRbvJl91Bq+Z/N3FvGiCMxTSVaRjvIj56yNTlksGehVvIGE2mUZ
rX80HGYmcaqk11QhR1o2iyuYFVZEn7Jlu73CFLzrxWHxF0l0CHomKcrtlDnHF9W/
NvB1LNAnt4EULnZHj95yEW5MC01CmdYxxQ1ahKYB/rK68MEMoB2y+w5pw5dcmDTR
3ESNSoXARX+/25xns8/2zzhrUnaunn7I8p1JZs9RRH3jwDaGdVL15CJsNzyOXJ1Q
CTdZscYwlDSF+zes2C8LNSzj0BtxrqGkN7Md/VEwnWcB49Fk0CsZRPPfFYmKNiES
w/ZxypUtqznSPfkcwF7MsX2fKrRNFQxf2AmgDF7ah/+bNc6gWVPJYx4mMYv8tmu6
GaYiAx1jgxj0vXuOmdJuxB1VKwIqt4r2RjhIkTfHyTaEcTsc3pqIjKZcy7Zen3F3
7K4buj0TSzrftwJyPbO/oNd9m4FdN/8U5k3Xpnf74PEv2sJB7TJGTmAHsz6nYuc2
LIhLzezKzGTlkgWdIdBDuOkdm1esLNn6eY3mI8sjXMliUZJiE0nvfVkc5QoqcXmA
eV1FS4QcozOrv32DF5HGgue6NSF2AEapXNWLSKG161XNvK8O9Iw+7J7r2xtIMVkN
QaXTaAl/Np8e/1by5UPBiYUD79FmJroaV33VFFrjMhhNFGJqy7ziL5+aRJ/1ZT1g
7Fq97BVHWGX6AeQYls7TIHvlj8EJFDeaJ/OZtEDKbPlzCGewuW0kqZbJgBjHHdHA
HcAgjnyFPQNtBbHJiRx4TLElT8AY9QCh7eQbKJtZf5CuhCSfmzhR46q42RKB0hY9
Bm3enQJfNmjVOfjqwIgDbNiCTwVXeWDrsGA+sIdrhDQqfuoby9/bQ7YYF4a1U4CH
uzYCxtqnLK/N9z8ryw7UEYYMkZUXA/DlaNZ91lkHere8Ue2k50xXLMbPT1LiMyj2
qx3xdwK5WCE6wqvut4ZTHOoZgM0tY7twSdjoYy9si24w76cLxWw4bR8E6sE9cNov
IkZwzfIh0MOIC1FDdGGmAEnC5UaqEQ4qHBg5ZwNPCXpu9viBsJHICPkcT5eB+yFs
7z8WflcL/+7YtXceXerLfnFzwkG7H3j3/2ZuL0EsMp2HbeaDwODxgXefoYDRJQky
c1UDA8h13ZuoVZ5qb95yeFgKorphc4puGEpyyAvgxJzfSvKb4e5OEoHLOFJBbOX7
dDdW63s1qeCBlXvmWccYZkXUY/CRBjBplZSh2OlA1x0HwHv1ZC0QVIeakNZflpmr
bmm+wFKT7GeBttMK3tbpJDaZUtAxoLK/8bKmi8V30R30Txb/+mPmJgqic6b99U3o
6zdCu4fX7O6FmhTC8IfWdXg49FGvw6Re2MbTaXk4umfcO1SAJzD3Gjfe1ddgTy5m
XHrUi65XnDE9eCOYvkaJegvo8uAPO1xceP+nOJWQptbAgVKNG1Ja06uOdm4NiFNv
aiIFq9Q6EwqftoPCxZ38xQpmnj3hG19+CS5aTmym7jloCg6XtjUQyEQxY1/3ZXNt
+lmrAuWP6jzwTyImOMaoGw840Uz5CgHwED7BWeq4brik7MSE30M2e7JcqOkmXtbF
xd+x+BL03pPC5MTTqmpJfdgKd2X2EIkKMKxHrinqxIC6TVQ22XpsX5GGSUV/HpNq
OdZlkWbOUcOeH1DeR2RJHWvDFtLclRh+5XDbGgEdpktZC4GUoqsx/O2QwvKbmbGg
iPoFqY0XFL9XU0bFJ9rHpP+DYPJGroWPk1srom4pkk36nQfcBbrZW71DydNBzzQc
wqHYXwHIsgl+vbqwcA6WNJ2YIRU5XAeUrKcHfAjp5hJtOCcupGYJ5l9eP1cdisL2
y+j8R9Zuw/6Ohf7vU8C3Aas083yhFmfcN+v/bImYBtxbWLTuK3EI3pd1+vNQPRTs
UjBMGH/kaSL6ZA+W8jNtYW/5nxyRnSCJK8QvSPddQkTUVw2U4pbQif4E3C2JK96/
tULrHq0Pg6POQO4DZW13uClE7vVmNd1Wu0t/LildgXA/4FvKQtcHHbAazV00Hcu1
LeGIw1Ssm60sDaLXtGe3d0pPuYKZvTEEOT2l7qWieccJSeicvMWDPwWig4bmhlwc
08segRzm0btmvPk0oO19t6POZYJ29MQnfycWgmdu0u/tLpdHJwKqXH8kiiabX4XU
gYzMYtWjgX8LCpoJetJ/nfvMdkEjZkKpmR0TFpeVmTf9wi+DrZ5xAPEZlZFH9zJl
zlTN6UiGh+zNMC7Gw4vHDMU+awXoG1GzlKitiRwWUs1XlCgdUj/v/ivQur6qf9IB
N+f/H74LNr+1B6lctJbiBrejcTU1YnKjRGi6B3OYlpiBfqwGpKcovm7FbCXp3KR6
Vb/iyRiX6vFb+aQ+s9qqgho3AW1RlY8DNWH/AYcKPruq6qRhYL+7wJp/PPBNwp8e
n4OSCHAnaaaDU9k1prCiAgIhAG4KbKTG8HgmXzf6UQQtA7QyDvOhFyIkaxCtDbzO
+fTkFw4erNutcXkaH9rBfifGOllcCblMAVBXr5cXFo3S2vp2DUnhTi2MSG0kgrhs
EtWbu6qFjHvPBxQKIRVIKDcwRxQKpOdtOulxaOJeGB4GmlZFMftLC6Kf9EhfrOhD
7wpJrrsC0yx5gYrXPORCwQIrgM/fNF9F34nDw/0wyNjzGGpEZXhOh37N481+6QYQ
60iQmXIcDRi8uRWe0aZBxsDJgyFY63zeZ3nRViOi2AV6Vrk1nYkk1Wq7G0hJT+fz
sO9zySU4L7yHydjcBVtsfGyxJLXi/tBbcepuDmogoAYoVpS/CnojEtt7XoxkMRy3
03KahHGP85IkGexBBLw1l4VbcwRhhi0UFuuF7zvOfKOC22l9Y/SFYGtpTPycggjv
BYoRWHjT8ClKQ5u4uS3EaEGe0oIroXTM7EgFgle5QvfriiGTDWqB9QYIYCOJEhGM
aebSE4nQpYF4zOA6q5Ljx/WcR97cn8VcmPPfakr3v7sL95DxFEK3gsWwOoiRo7Gt
PrrrK2lCXcjOBJp+YQ8rJH/CdGgOFmsz0D6HjHRzGeQgb4vIbXs7QYKW7DNu+g0P
cttd/ulBNgCyHGeKEhy1kEeGvekEX/dmFEh1i/dRTK/Cck1yVrPrbQNkEZsVG1dI
5vrE4wIBNhpuMXr1BAsKIHUXuY8FtxWHdAQYGGsLf12azgmmKJYCVHJuuhcavK/R
wiWFgS5qP9VTnCwlHh/4oiM8gnYoO+ICehwQjv3kUl1Dli3Efgt5t9ktLMdUBPqm
POKPwLRHZoqDlDbZYA1SKptjSg00kEdjoo6q/kdpsF2v0Jp1LIczwM3vh0tX/kfY
MSVaxhWNkw654XpFOXW22kLkzZDhqeNJ5SGUv5K44nIjy8tDFJ0sk44a/nRAS5ZU
KJ24mGA9TmvCLwkHPfjWH3KnR6lT21yvvjxOCU7ONq5hkeoJWzFZ32uIbOCgzyOR
x4qEMzS6/TnEC5wuVYDkTX1OycINyQzoJLTbWLzbkvDtuKOwXaJPZ+Exi4taUzs3
x41p/A3egHj79CUbcywFs+Kfe7+mJC06nBUNZ3DTmofwX+OzFigZv6K2ERMrRHJN
gAm2o3Nabc6pzMQxfYRJ2B4swOYU+pZqk2UT4Rkh5LMtTbs+BYXWYT6yxF31dWlh
89scRaxDyB7lskNu+VCDbQiJrkqvFSOX3+0W8a/dWM6jVbrzDVnKOzb5HeEP04kL
0dAnA728u/Dtnk02B0FuCHKSr184KTe3/Iwl/CUzIL/luWRHxYY1AV4oC/DBRuYc
0rpqbOHGSnrzRb351AdPwOeWzLfz53k1SU7+aS0cgJpm5Jv3FA+yd80bpz89OVbx
iZjOJZuJe7NW4FMzva6aRNxDOreedtqwTrL0pPJQRtcqgyg3cm+p2pFUe3hpAdtl
x9HwUOn8V9oO5hYr+vfFiPBaAeSCvrOc5sgY9PkmjHRjqTelgHHQYQKfE3Mt1kmH
QBPPdokhalSjGiMCfA801jnVsrbnBkTs9j7L6s9HPSGR2DvnrOYyRiyuppW81HEr
RTnk9YgBJEGvowE3aVA7wGQVrDpANXzAh6Feqj8Yo8mrrG3Ay0qUbCnKi9hyvROH
6c2CSSGTaVAprWTpF6K4OjkrrnLCVuf0Q6Mh5btzh5uxu1Jpf69JvPuDgXeYOdwb
j2J5iDtS+NL49PM0eIazzMPfy98whkTUP/7CRZJKNPpQBH7HsJ5hg6UJkoaGayXX
EMcxr6pzNyNp+RgMTR43aNxHXy9tbybJevznQI0ulHmDiZqMB+hWleuGp/bV8Osg
UW7lnv2ZpIbSycNbBqTJ7bUu50FXDr6kjCXFoyWYZjg08dGpqM1bc7ENdxxO1nbZ
XDrdplnxtNk5S1ixw0L30PWg6kYEtNHFK2hU/lLuNCVCwVlcpMyNtrTHvR7xHPGe
/N4fQT8kf4ujhrbYoooXolk3iOTq9EWhQGIsyhDcil2MEhD7C8n2NNlb7TaG4mau
AF29fGjr4xdW2HY5Fa3JFIVWd43Ec9/aT7wgQWvW86MsGEBQtOY8vbzfBZPlFWjs
RoTB5Roek5XzQh+Zlr29tjag0vYgan+1k6E6BYCuB9i8OFfbQjEWY8B4d1AMqq8g
JfPfsm9E0jhUfu+F3Q9XfRLn3Y16YKOLaPy4DT5InvNcxB8ZOq+uWvZGT7QnSABz
Bd1NMjnkvkG0f7MwCxgNJZzKRnOTgpXvEDbYRePkcgGl/GxpBoJQdJ6dIJFJcf9j
5F91OJa3ueHaPlqYIbBawhT6ifcHQcJVLEwdOZeaQB0gLQbprZpx/73hkEUxm5+g
nMPv0Db/IqbdMtDUEfVwZ1xhVtERhl8E+QB6jExTtaH8cMbhDU0iaX1JUG7wSliz
+9G/ldy82ZvvvuYxZVPSfiDxfM5z4uQMjhDcYw9W0J8WAIdU/MO1NbMDYixX8rrJ
e/K/3/EAHXcCUAPZLW+ffdi0SXHgCoIVsy3SAtX4bF9py9pxpUBI7HTts3umuQkQ
VPq6vgf0hJAuvJg9eQrPecfTYGB4yedLHuvP5Idf6l0XsGsTqwV4QqQHz0KefrCj
cjTUq035c1EJzhV3PN/0nvmPcJuFSfaRuGUcAnNHQ0Dhec2R/J/5zytbiG+/SJ7S
OPLWYInW7lr549Iez/rDphkq27sKK9SA240J/MNku+Z9oRUYImO5L6U/81cJH1cl
wT3CF1SosbFMx3WVBQTEvLV06sUdqIt9dSUXDJEft1AUApDjSuFVeJx13ScJlaOC
uCTik1uTTkoIDhGqBWe7U/mJfZ0ufg912DAjKWtg+Ot8WqWbC8OrtSryp+LfuWzh
JCeFmYLviPVkICGpceUxTkcCihzU/KmjImpCtQrn1SFqn4oDnxcJMl90dKrDPyiO
Awq8BASjm5ICa18PzbI86szY9u5N1N8yhnb1NFVqIjuDb333uvFFqEs2UvJFJvN3
3CvciKl8J2byhNTaKie3iNJFAsWQz6xKz4mSrOPJGi5eRL9aiqLqRHAAZoc+ZcSX
tUfpKWAxcWI+UUEVLwCrkF+kfww6KU2yHgKUqt35fIRA0m/vdL6Rti26DL4U4wsD
UduZ7FXchzGyyn8aISDFSpuOKraRs6qkKMf3oiMcnjn5P9HxVok22jMjPeEhvaA+
Qbaa9+B4nOi952AGy7d/6uVBAL9JjcjOOFbqz4xzwzVz8Ek7MjPRDEarnt72fjpr
TkMSKVILpmLKNpXtMEImntySGDldtE/VKQEWE95wbG2yL12g8TGwdgtJnHVIGpWf
1a3UTSEGjvmuUTCLlSl4xB53yj+Xe1T27vOfklfFd0SIXzBeFM+TLt65m93MCso5
bNEGipWxVSs2yaDRRHoOxqRzy3ZaB/Ag5PWMmUf8WS2VCkGC4me3Gr91WLCkIb4M
l9yJr2LtLuI7Y+M/OSordU6e+/G6NdfH3wTlnBrZFXGnr0ZmKHEB+P/KoV4jNQw7
a0EOJPWqFEpHI6lEqRSZ+LyhEY9QybhVKADTSXfxdo4uWMhuKSHcl2fxxmnkTY4K
ajzkaQ/wqYBJLIRXOHBS0AIyWwpHcERRhnMtGv8C0YLnZKH+vDiHLSLa4/3SqlBH
TWu1iLV07uy2yhzkD+EtspF/84+m9sj22V+W7pA2BTFBoeqklWFEdzOdR2Zu5ZSW
AVK/ojpH8g1rGrMLxhlI63gotJ3XGHXfrGTvnQHunZHeMm+frwycCKeNzv5yFjW8
WQdHAZE+CKu+3GDDYhd3qA8zUywzeJSfx1TNnZl/f5Yfz98F2t8vyIT5bOlzTl2y
cFzzUWcN3EX8Su7hjhkPSjdvuvLuEfXDbNOpZeRxgg5z/cEunPGM5s7Kae4NbIrI
0f4ppGhp6CSx/KZmcfSwJddqNrYgD0xDwBCDAWhIZ/vRkn8WfMXiI6jKBSW0ieup
xe9PU89vyCRz1NYwRcAxvQt2rXvp3Lymc8dTguaUBoSgSx2UhlR4XT5hROH0GMPh
v4dvAAtGIkmTqbsSQRwUC9/0jb1sVeJWOlOs3Am3hHIHMC1w2hBqj2aNNU4sf54h
onhndrvj3mL5yxRua8HW7VXwQ5+s23b7H6opCO/DrX8kpTdIni5e4Zlafa1RFno6
dOKrZcONGHpcM3xdMG9Lfvw3ALspmhrvi7nN6LTcfaiWs5FBL9THByoXOQia0NfY
2MdKEsBZjPHij2WP5it+ApjB+KadPw0AAIPQZAQun8tnPmNSG94gEJKPzSwVnhRE
E6/rcsfieDxhRC0+2HKEVWrGz0n/fpJKAuRo4RECOW4KANT9UlbdiATeMIqjdP0B
0qk2MlevAfP7wtVIrfwscPyVEEmS7cHhj1q6CEFXt+vWWXU/i/P2VlxIfC6z9trn
LMrVstSis6Z0niygOIeJnwlJdNb6M0UZHfzRCvUHtnod8d3Wr4MeopMzDfukph3u
MLqOSpTO9aKwwTBeMW2Hhsi3M2TS4ffkAb0ZKR3JOK2iqot3L4zceWRKGSmySZpD
8bhY8eMvkdAMmQTu4mH/uNAMJ/Hn7x5KNWUOylUO84oLcizWJRpIlg5lxDGjkcxf
iqhU0Y5zq7/FWNYiPrsdF9AYltj5FtefgCMEOBMIAFkGtqFVFxR2N2rBDAMcUMnO
ihv+XM3tsAXXnfgYLL61Y2M6k096b5gOaTssrveH/Z9FCXdngXmCwiMX8FQTKAXN
Fh/e1WffGcNm58jVDFZv0Hrq9xKmsycu3OMdSNObHJ+I/jV2hU0jgDCZQpQTCu/p
xclvCqylIuiCsF4FeCzYskxwlqd2e0ozANmht034g9Dj3rdIEFzqkBgQKEmzI6z8
fIGSv7hyu+QZojYIbbNLbQvd4WmTbAYXlJdcHsR71z7cqyzJXnrkr+EiuCzFblyo
Hhs5371UKTOTeIrnZsJEYJVm2R1Fa+wcpNmOrzZD3K2dry6TEIKV0HjI5mRX0L22
Lu9OL1pfUS6Qt8yDdmCR2cv4d3uz1ViPTAPaggvkavKqsDQ5d0vipnMNV1XmZNGO
283WrP6zJrXFrMtv+WEc+sgEoP6tyqhWUD1z1vkYR82+6AnKs8hbrkUyeOodVAh+
x480OxEwCMbXqXObFkDD4dZse+LGxJQ8YX43LSRdIdu5Stk/6AbHRg/0ochPlE0n
c2Qk80QLEfPnAp14BHKLI27J14m8F2V7QX3C6+p4RiByQ9S5xlbX6qZNvbevEGiX
opG64Tijsw0Gu1sIYQfvhi8G9AXqOoFbrYs40vSMgKw5QI5AuavmhzH73lXBtFKo
nyOx3o8LoYHtiwAo89dlkoa5zzenvSct65gM2b7WjduPNM8tFakrKiCX7Nt6yC/m
LFIqMJPFleOXTRXOuHqJdkkM4eR1mA28fHZ5wHI7Xk9p31Fdjh2YdLuSZoQ2O4nS
l1DM9R5Poc1ao7syXQG2SqL+XfGXGkm2RPsc2tjWymI3VgP0/SVFY5NPCdCefDzm
SSMSyH9FU/f3MszOwW3D3cW/leGkiqsf6iv3Vq88Q55g/RBPBvODrLr6rvL8t6zD
RqrYigiWK1oi+jFRxFeNx0GWGEI5LIVv7OMGLW2woqvame3p+qmpDYaxrlZwGAsv
w67fxRK3Ts2sDQM+/d+AFromaL9du1ia8p/uJAQgHMqjpbvOfwKBZNis6yLg6Vqj
2FBC0VIKQZqzaq0DhwqxbD2NUH4vk1t4xks4sH1GyppxuLDlWPksIXWbdQAzHxQo
KsaCStvnRMk3+GE/0e+R4xT8x9soOj4YUg417tQj9YkHkvP92D5V1ZX12ovZgFrH
Ta7S/JiSTDwe2snhyBsqhgSd/G9F7E72KfnzxCqoB8EigDhNpm3WhXMYryWkgCIH
qK8OLzOnJcmzGaOndAgwHcd+Qypt8XBE/Op6mdxu57Qqar7ORabQNs239rmyG5xs
O+27CaPoyhn56Zxp5+Pp5RhPsG72e0JNyqfj/KVuB4oizLq97zcuFp0Z1YcciBX4
oNAXKBwNm/7snv+lvozwhNsc26m8DH4ua2vEJsLI2izFSeoUGXsn9+fblOY0nER8
Dy8apI+gYdUHwdqDmJHnQMd6wE80r/LanKzdl8nBbBoPSnXPTVVrZqwqp7mhRlKY
dLj84Tk3OmK6fU19PQ61PqH2UQZRi3dHZERTs+Ed8UC/9nPpbDZLcXB5VOoo0MyU
OVY3sMS6W7gJk7Troxn9h4bEESO2CeCSaIUD29fPxjhxreEaK50hXDZ+IFlIXvcd
PEgfwsJBIRswGvhOYwIY4DQ4kK+cB2k3PlnVfiGWS87fSGkA2MPCU8yc0sT62628
XQXY9RV0vlZfu0WXsIzkta6nzje5HS7v9ru606vVAt6TCwaVJtWcrPBWJTCdFhRd
u4p1tacw2WLOHCd1/V0xqCxJNKzjxPW++LEvUkb20CMHWe1m2h26+VS4a6KW7A2u
EaTExm9O3DESgxjSlcUPFWjKbTsq1g/2L+pI/5xNt6EP/8iOU3r5j7x0UN4JESDg
rq47f213U53+s9myoTW2srFs1jAL0q+QelNgG/civ4gkbERcVlqMwnClF9trum06
534MhsafwsvO9DP+vi+jNHLJ9KFKFKRzZC9C6Jg37CGygBwiXb/0cnZ0MU6cj0gF
nOhWD8tC98PbmRqfIGF/CkkJmUIdeg/Hp+YcBKXBqsN0q8vC3nF/bDQAJbTsV1QW
11nImSBMIBHTlX1kv8UG+pENInKRAFEHOdhjfSHEm8rJe2P6xHOANd5tpEHGjPrP
M2YCvzdm54tss08EMt7pKz/UyADjknQ8lFDjhbqtFWQHc2BpPiEiK5UU1wzS4Yvw
q18cyKSnDYxhHnm4IJOdigGVMWxu1Y2YqPd7cg73CaMbDF3NdPDwD3VA05VqJO69
brMs2+UScbFeUxJiem9I87yw7PVFYx9GTWZjKSEHdwmlLRhr1TB3l1rvRTC1i973
eBsr2UEynyRObVQxe3T2xowcpErgA4CdRTdBMkXhoymt1IPJHqDWIASkt2BnM/MC
uifBgrxwLUy28YvAAu91BqlVpHv1fBhnLNWnu2ORe/K7ifxYCnMXJw9x8pCZZ7L7
kHIR0mapbFmplW/iV1jakQMNshp+6nOFURDBLFGgpHIv//QSkVhlvSSV+IgLg6dm
VwHFVyb6Na+c8WEOKQMm0ry2PRurSZvOTLSW+OSr49yS7lubWHYtaV+T5IHbEYw3
yo5no4UsgREyeT2vi7w6MPb2EBAwzCshMbuS7n4+iF4mn1jjWVTQaeMKVhMUOpAh
C1Ib2MGiyOamByC/lDKxqE3gB2l4JV7YbBVq2t10+HYJoAd1Of9+tjO/8rSo2PDt
m0oOznRR0tFdX++enZ/FFaI8mLHXJUb6giQp/e4clu1lo1mp4s1FBFEoAZIN8lU5
bZSrIrkcsiTnh62zb1ExlOs97/8zTEmBvaDyyEF29UTn4jiVa9juSdUz4CzBJnqJ
8ukv+KoCxvW4okYq2bWeMqRXUcO9/SNabSl6bN0Am5JibQ0RqzeBaPzHGlp5hcAe
eu21YD5Ix1dPjn2QyTM7nScszms4AR4VUdWlPzB29szZiGBD/i5TUdV2gUjunNx5
HT3kmIMqkNS4Gt9J6UdIbObelbHTdJjZZxNPBLYBuHbIw3o7/sHMOgCEE23ZLlI+
uIMP8M+XbFFeWxmHOCFUadp0aDmL825F7+I/PkwIwl3+Q/IcbL8D0ExQEiFLJOKy
V4MI2TM5QnyoaZ/kwdfwtY3IMavwOqtqtbp8nffEwj1pOGyLSWYj6ZAnDp37VSkk
jC1gFfOLGHBoazpwBB11BAew6fBggVUgoDbhbT0XJkJyzhp0LLxlk22dCPyKPE+r
UVhiiDPhBPjofjJmxT0jeXH/Wg94f1KMq+mPL043//1UQLYL+7Q5jCiv2gTKEnd+
giqs70/pj87t2mta4J0Ya9xdCJgLrYWRGTNE2Si1UX5QsaDQoF9UGpXzuZpZQbwT
+McWR5OtWo3+FRO9D0Nd4KpY1O51VmpDImOKfxS6X5Bgb0CNmMAyd9YafjyJt4tC
PxfBF3dVoMvvQ2bKqxQMjHJf1iW8+2TS8/4fzzPqdFLM97CES/yh8Tpf6UCcf+27
FrsDRfNL5eZH0xw5MN5mUQ8lQAM8pMJQOQD+NFuBJue9ZlCXf0O1fxUNykZV5I6V
cD1tbXA2wX6aA6TZtROdyfDzIJmfXXSFHM70xhsF8j/ocV5XTLo7AwZfUJMnVq87
xxvQbQsSTKp+3kBxxIV/jl6TxFG3W33lAXREQVBO/4Au6aMGaNhi2X2bnUIj4S/j
FUQ0OjiQiS5jCoUYcTK0UukHHfCFj+8QtNMg/eVMb5K2PRfPfU/BDRiNF9QX+E7o
GGJm+pyCf9mmZrIDbS+hyirDefkHR52yg8GL5Fe6Vf7pZ7gVl9fA9TDTWhhA3iO6
CY4+QO0V/N3eD4qdHpQ63aqpZoiosbOoZ4Mbxvd/uXXZFmKCPlZVz1eiuzbWSB0Q
YcfKWQ1ufqZ16e/UqlYI+VWLNtQsfV1KxR7ClSkNVF59MLAzE9rpwDFpRFtwvrcX
nYKydE3Qw4ZbqKfww9Ox52fBeIaZ9DSXsdAIZ5p/l3mpgCAma3UY96QDPrJQ/dkn
Xr6OuWmcQl2QTXhWwqkamZ+dPR+MKKVkf0s9WPKU9LCDEsFVx+n1RBMj32QVV3dn
GvKFlH5b5LnS0oHWr6+dwuakKontHYZ/LBDgxVBazCUkc8g/FBF5Z3LOOH1UstVD
dtSOpNaInVo1mXeWVIgG0Vsd6ca6Ko7/pVNJhZI+ian5TYBdld64Fp4MVnTfdXx7
v/p3UNUPsQQqSI0hJsALkPk7HdVq3EpnqkCsuXbFH5p/28R4ey9BUWralR7UK5Yd
dTlB5eDKS4jxyKaRwMCROp2M+VYjpUNLfXDtZKOSleDu0D173Y1X7rGABwZ3dcHv
KfEjct3or4gQ0ORsjHuvgFDRDSBhwYek/mR6Y8qbbhDMy7/EWeOMgHWU8yxkH0dm
ezM7AQYQtomEDRqKLfmhRXh1bxKmOFXP8+b1tH0YeQ38Wh7nzSDQOSn6kOF/3dVx
Gx7DKMmfPHGY5X2Hk/VudU37UQRPd6Th6G2P1QELoDp0Z/OwBPtwmj6l5GS2LD30
UHEhOGUPc7SGmQ+c9fqM/YpQ5KOZ8TeXBETNkrQH+s12XMfKfz/Jt3twGn0Fwavq
ru0Q8KGc3eONl4rD73whRDRjdtsk0nd8yAyb4uCFVciWQ8ZE25Ifan0FjTAkOpu1
mjM5ESs479rIBz9K5stf6UZa8rrtwdHTfTTTd0dtOjmABzR2Cj/3ekXvUmngr1wr
DnV9+MXqbQuQMMh7xVNtrNJhgZWPaS20PDrWRDFtTFMUNuJhq3RsxGZ4pzRq7nEp
N4acHlXli9RrPFfjVMXobf/kTnzibo2NXRjoB3JhNMR9QA9b4nXzVAaGkxHFMEUv
ZweFu5r1zpGqnlrZ8O8HRvg/2YiarpgR6d8uSSEqsFcnvYZsrbngmeW/eQWqBfjE
00o0B/X9Sx/A8pPgcgIGtdc0ZcHCBz0cpQJx5S6uWRdC5clbp5rClZzN9K6yfwdY
RBL/8WCZDjRodJwIBQPSg5eqK1cJLmgqf/rQvmx7hmbNDkbkgfZEkWu7kwxhA45N
GQTfmdSOM94jTmLSM94LXROy9dR2RF0aGronS2EvkYccwMeyLmXGqZEOZKf4QgIb
NIqpvli0xaFsEJLAxXo4kdvbZz97kRIoHvOTGOkTZJmT79gOJYRGWl/qZturaVzl
lH4whFgYYCJC81bPOZ4FtjxO/KHkWRi731hwiK0lE1e67MaDH596Z7z1H9v5ja14
q0ldoQC1i6J/GGjYlit5HD9ujvxZvAIPOQxrz1sXVXmwypOYhbmKpUJXmR/e9o6u
cA/jYqnBaiE3np74JV5XsdABaHZM5+FKUg8drGvWa612KVuOJsUhsS1tHiLLKmng
1nzOFSu9oFCLhMbeu63JdJ1FtWgi8TUr1WUN5sKy9DBKTfjIzW3VzrZ5D1Mvc+Vt
HOAFX5Gmbd/qbAsIymA9YRs9CZfekl7ExBNjX/cpCo7RmXUA7tPj1B/oGjmaJqGB
I9+Tqf2ykhgP29npM1VybQGr3Ht8NsagP3rM3Qxgh6Mtn37oynjiN6vu8G9KDHZL
QxnTaZPubx9KqRletgIKGF33XVBJuWSHlFwzqEneZoH1hrybv+vC2zje/q8tdPuR
Cf7wnLzB3H/X0row/qhBTL4+t8SmxTW8EvndNEe1NpJDwwPiVB/9TKCUesLjpm3E
tE1mqg/BOyhuIWdK66noN4DUGM25OR8kHlDQ9iP2KjAkk4DvlpkKLJA25LsbOPyl
BnZ34TUp8QDtjeRdKJ4nnmNqEcXbUCXR5zKOfkkpNTHpuV3Aguh9XRb9s/IzCJOP
2btBQQ3YBb3Opg9Km3UDJNbNWNfdG4SE3LjFjHl763LslSvLH/9whsYKkjZHH9PF
TZjrV6XV1DI7wznTN+ee085l+FqdV9nnRGCU0CD0xw1dG//cER5L7rxKiS9fD40E
xsVJVTY05anYRdrVnVYuJCZ/zBMD1fGAeQMO0t8NlLb7XdxVEUCvVrNG/HyYH16A
JUyyv8oLk+e5MXuho/vB3TCZeP9vWNIUSpsQbuJAbGod/nlmkxv2Kzxelbw5lYPe
DlzqbVo2oB8859G35Imf8ZoTN5GErFPv+Bmk03SWceN/gABlYEVI4ImXSMYnH9kl
j85WDxjN7HmmZEhjbgggrgdtsDtl3WMmBVHjGPtOZDWcy84MVReFKGLA2/P6BPfC
T2s2fVY1XZbCxEzyOHthfciPpaMIR7m5Dbv/SsoxOv1/+ENsbGdRPrluZFF0AVNZ
CgklmqgHJhNG6k8+QSEfMcUMGFJ+ixkpbLThpDdRpVxH8Q3+I7kjrZkIJXl1Ld5t
Xn/c7pzqTlk6Mwa80IHckwcEpJ8GDq7FB1+PXWaT/xXIOK3Z5r8PvH0AAJ5xjwWj
uTjv5mjG6PguldFLDG+oSffWRfooTYViHWJMvAHvf7j7YoU1E6MXyGXgmwr9iq9+
NWHMwA8Op6+8GtS6n+A9xAcW/mdTQa0ZH5nlgO/2Squ6NoBAi5+0Pfx3qof2MMTH
Kes6MeJqou3wbkRUasWpmhhuzxNZaUe3Cymh3Wn7kMA3SYcwgcPG9G/PylRb56tF
CFjtoCg6GiGP1ENUfhMzPbcN8UH5hiaMOmqns4K+oUWGdkLWFtec5RWUJD5NRwJb
iMf+A3KdYQiuX9exAqUYKUzLQWrbalUtpGxGL/X5HLZxzum6bFB6HrzeizTesCvH
VPmdDJyYXISJx1mRfkEssGzBmwvYqFivLMaWyx0ps6uEPZyFTZCD67Am75apV3Cs
dF/sX0OApF+s4gWbiluiKkXwON71KPccKUNc2cgQsSBXs9Pphiz12rW4nKhL6MLj
jHraTLLGSvsV33y1NzXZv4iCdvh5LDUGsrG1hK7CX386uAT76HQScASoikZU3FP3
iYO3Nwi4w/qS4FtxVkuJWWWr2bUwu2tlPgRtyL98HS7e4MqO7X1kge4h8EHYcveY
sGIvwJM55Gi/ii7Tm2oyjrGfFD75O/SqQ7Snx13B5bTLRN87m9W4/TC2/6BqIArz
H47UhSGxa8Y0phrZcZTiKbiI2sQEgvHpImeyH6084MlC+nyRfakQY4Iyr0dl1vXF
wSj9ZFV7oHO8aOE1bu1Q2N+tqlrLXuR6uJH6ivbKInJ9Kr+NV01u9dsH8ARMeWLF
fzlnWFW0WgHbLSbjZ+cKvc9XJPK+mj6EJEB6nz9QxBzAb4xegoyGLKNnWKBV1ii8
UH5NoFsR8KkM09Fxty07Efj5BbLWrWUT+tTb63RVtgD/reeyuuSbsz4ziR5gs+1S
ZdVE1JcaYn38XUmA3wy+JfF2LTDOEBSbINdI1q3lPqJXHgkMFrSGkgs7ZghSVRDG
MXZkcCrmZkWVQeNLXUEQhhjWOmFtd0z/IBhoBxH+mRB7Gpjp274xpCkyc+Mdf/jo
do9yvNdfZgGwYEiLij3/Ig0Xh4KgEKpytOSgR3JrJmPEn7Z55fMxfGldes0hscZc
CzsbflDFwvPGAHKP+KSR5sLSlyKHcHU1XOIKJNQ9cUOAfVHBJAvVfwkoy8EzRvtj
BSBhGuW0cGgiUvs98ULDOX0iywQ7rqNrkzqaT8MUCfvM997SDrwTx0uiOSo7TXJE
n45oiWc5a5Ypme2jCoIO1TL1rmfimCKUsq3heS+Y1TbROAOJEOOa8QMitwlkGhgX
mGtgVnonvbylfrfi/BKkl7/sjcFFjp6AsaXfCer5t8suvDQAFXjTCaaB2ySfIent
t6OHGLvQ5IBjVjtJvyB4b6OIsS5aIyPxobcNesYgGyScIqNOjpF62MEjcQGgyA2c
SjHk7Zc/Pe2fbN72dZ+dJkawt/jCjS/peX9PbaZ2VqBnj+VzMwg6KTyMht4KjvKD
RnNw11UX5ulbPbESAePVKibKJoquc+i1JAFlMoqJIT3HT9VW+A0esX2DCbjwb3+P
KFOHOUeFijVWoByAr8kH1FYjx0vpvPeG7aGKrFIu12YncrC2RS7lT6+lT/1QRqHh
q9K/U5Nha/vguLhkQMZ6pRRnkAg0q+AsPvJyP1yE0/7drtGbGhV33Ej0UFAPzUZZ
vZ8HIIyAJjmhxX4o8QcbAO32gGVbnCxsB3moMbFIAwJeWUW52uvNaDgbeahkLLub
GlnkFvkLwSbK9kxathHSfWl9P3xGgn4HwtQxasxAkKk0/p0P0NPdV5v6t1VVe2MO
FmOBubSq/rhMOTFARUzl+4GYbgsPeD9CviXkZa9Cf6gw6WgBrdq7ORFChi9QtQIU
Rv6KqO9J4+hI2qDYL4/V9eWosEufjHu5nvJzHrSG08a+dB4HrYInqPc1i57v6Rjr
HnJSXTsOACnKwl+5o9Q6kwzrzVbcH82WoL8wxeBveuU09UeQaxS8UDZb/Zo547RT
VbzMOruQIUmzgumIrw8B8Hjb/fTBr2cNkCVRUPb0T0VFcnDHsunxTSYYza7tHdxF
NZ6fpSNZOGtIVD0vYN2Uz5D6JmFCddmmkgwfBVl/cSq93UgvIafwwuiqKVj4RxUU
ffUnFuTvMKUHkNdFQGsZWXym6AZo/Tu7DMc8S4mwvi/4O3QV7W/kmdsdghVmtOch
q0sETD8/pqf7ot1VB2UlVWDpqMKcMJLtxLFP0JmljHX7vLhlz0FkBi6SlQkyKq50
/ollxyRj+sdLo3VodKV/zvxcvSi4EKvWjaqeXq3t49Y0HO4L29ZfbNhnnZ099fp9
ZlRxkxkiiLEEKt4oHVoYj7o3P4+qH/tdFKcIumIdwqN7hZRmjhomWrM/2SQpJpzj
q+ukzsKQW0JVG/vCrByCUWSxPXjGhw2Qt9uNz2UV0S+dFC+eBYUtXhMmfPQliZhg
cUWnXbU0pKgOgKKnx3zpwfnic3TaS1vHrC5UjD85dTNZr36P2Go2PnC5tCYIoCxz
mWW4XmviGKdNryu7TQ8Ach8Pr78TcN5Zbv6s11OQd1C7JdpdbpGvt5VkzmruI3Wu
tWNFycvHQl2ZLu5LeJ/v/k6/6s10d1GvSc+ry21KuWDW23OwbCYE6Lkb6js44Uvn
z8u40Ld5PWiycagOg+t9xsKnYr6VEFHRUXId2NqapS2mk0DM0jJWkzyFSgrZmal4
fNF8Y8XXdiV88AuY8SKO0XOgRDSUugeqUYLgwLi8DD7CAbNVfDvMWhLkqZaeQyGC
kL/a9l3vRKnWs/VsKIK+nboOsCJcs+afUbgjMTKQ7gTlGJDYY1mX2VIa05k7xP9h
75fPMCE0mA5IcEbJlieyntkkdULiLZTHocetKKnWkym7Y7I8GDPijmni0Abi8q4r
0HYgkYwlAhteZjZIa/LW5Ta47LH1HFRhvNznea/Vhmn4CzvutfMrNWJxMxXJ1Qfq
U8isrEcCjRlPe+jaXd0FZYVUILcNf5l7WNu9+q3xfLIM5jlvNiWYaLLd4MmOkwK7
Jz2tjOVXEKH3ZumI/y8s2DPxCPYgago3seb7X7lTMSrw0TS4aw5VW7a9EdIDLCVd
2WdbVY5YChYWkWQySKpTHpy5Ih2pewCcoqeyqSdogIAgzNf83AwvCRHOktxy5dG7
XDrXQ/tElZij4Bl3P6LHZWkBP4vVI/l2WcYYP/Dsohw4qwItAYR9TcnUnvnwCDn6
jd7rQeQ3vW7vbwJQdso5Sx8KqGcmR2VgTqZAcSNw4iWui7m0ZL/mYZqaFJjD0RWa
pkl3iLgS1UX2sOW5a1oVxWXBW2hzM34BhhiTZlyYJdlwIuEk1uO+ZVdL0G17X1rI
5bi6wfa8K6FDlVWTxqOlIrhnQBhq8NBOxWPpE/lEPaDURBOWIrcsYjytpWo/5+K5
mC/rqVFcYb3W8JiNxyGluiyT53fSsm0++WwF05zw+g64Sk9i5wp4V3NGpu6YNLQY
eG434M2E/aCnJQIiKvk/gfvVegD2jPAi1tsPPAzOJOlSXknVLmg4FxEfJHJ09YYY
Hv+AGih568TkLGHt0FIYuWWPlVvNsW+aaRN4RlXvkjRDkDKxODbVoU4UegQvfOyQ
7fjBI8HuFVD7+nwDrHmMk5BFHlTJhHR6cM3qLAh4FtW/WRR/5Ux6dKBubSwJsINr
8AP8Qbg0Rrx/nukzuvCToG8aALMptURpAlB6TtrhEwNRZQzbQSAODROlAlwgwhVz
BTKGHW0xgmDvdgz242cPkG38sh8JYWGLZDChFfuDUo8KIOH1fKI4C864H2qqxn/g
836rHGIOhmIFEZsNR0l1RgWtfHAIbiNdhU7xIG+6xe74kAVy7b3v+ZmAL9GdCTG5
Cboc6wxKMiMF5FiHGepxJa5y1uWGKVpG0jx+RItS0JohMqnlrayb+QbJ85HmqplQ
wUDw1HxV8oZ25RTb75EBkmyJZWyYMVbrDeyFpR0gZmwA/yWBT3h/ggRmRsQyUjvY
Hvl0ATWZSJ9Kq/uiQQypcirJLCGGPQDZJyhuCwTsbgcByndgepFrfcfyRUgcb6YM
pzDZuNxj5xZHPzu8iEwMTYoGksq1uALbiO7i48Zmj1S1oJ8yqxi90+AjG3TfbRKq
e7Ic64SW2qnp5zb9KKObDyu7z90Dm6nas/9Ya8BhhAhj6Jn8uxoCseU/G5atjuh4
k+iy4J6JSR0AJxNWXNYIFt8Eo4o+9xlQ1OkkVQH45rvcRhnzpeV67kxYMiqAff9W
YfQfHfDGigIcMXVblIzGXVYyoIEm4AJlhPASM2f6BQ+o8RBeyHENGSn/AC4HMIRk
bODfeiGtxMQALYlPDjqRgKm+HB1LqxpU0yr3vaVMSvCdz9n2He8YZhfuG4gJUPoB
R/sK+cobKxqg73jXT/qOd1yzn8yrBBDKlrHXggD3PCx0fMi9TvNwuoXTNqWeyD35
Bxetb34oDS2NnhTT2L+eq5W9UjO6zHOZnovvclS7nBL9TrPhXJaOkfAKj9dewfiz
z4TeGPsokSsSMNPEufKWcItUuHwwxovrjuzjz4ovgE2zJZUanS/35PRE9pftrx1P
WW8GzbqUrJIRwy+hqlwpJCK0ymCkCx1FvWmEZszBWltzAIW/MOpPNFFXqD4zqjc7
/toePC1TKQjzYx7UKLXAo9pqL7/b7tYYkzQrq3p4qBGJvidN4przIs9UZj9imsjn
FjT2N792OqrS+4HQPn8aGuZK8xZdabh30UcPcA4ZUEkyGuwhGt4x3YXYKoU5o75x
G9BD/epJZkn6bO/S0Lg6b/lCwgEKKoFqAzBv/Gb6BYPxW9z8GdY7nY3aOTtVYTuJ
SYk/HgZRtRgTvymZMXXmgykCnFAAfb/92lamDc2ALDA+BMs1r6+F9Jl6385n2dPR
UctOgcIXfGrmMp/g0MAzNTI0/VyXRMoM1rXgtzpdO47Wp0vMeAS0qtuovkM2p9XB
EwPxHzwLR5QjOpriuGaUz68t9X8/KeOKdLY4yiSZK0o/EHjnnbccDm7LvZZEC1Np
2LTiwEPhQstla/IRS3U7/24+lHLsDvT6/TMQe2nHEXzkHm9HFBK0vo6ZBIuq5pqt
SeqQ714f93Zkykf8m59hjpJt8yIbbdEey4co/fDss9vihVWPc7kBMAAkachTkLLj
8p+FtK1HQ5oRwBuq3pmStne4g+x3EcqwifL+r2B7I2RGzyu0+udpeCPl5Sa3zP8Z
mKvBIOj7wDYJqpcig4dnbkjJY41P63fVCP+9ZmKyXVlwtDOWpyvWm3AQdfw76D53
4NteK5QIXMZA4bxX1P75UOUnxMkAVFMHqzbe75OWW+lrFBpT1Rs8kIJLPb60Zkb7
hYnjUAOodGeoAX6beqPV5yWuIFuiMCaxZqmUcpae8WcS1u96bdhfl/uLfeJN3nkV
bpWuxmmzr6Zo/iXFPFChOHaK2x9NAJCqd64yF6UYtQcmY5T2cqQ0eEdZGhoKGgQj
UDJChX6y1/Rf0nrKAox7YHau6tw7jQXs2aqCNEt5NermJiYq+l7nhl1xoiuuvcoV
ktieGv3OqqTu+NRXmLs3ostj2Lf/jB0EGE9ynMyTdxEW52Bubz9AxTl28mv2qX9S
tbUROCkAAoeqPjxJS/GwBEmuqXBmqU+XzCsht9JgsNniTQdI9+zSHTUd5grc56fX
Q4WgAtSWXW+gjw2ANmIK/QGNDu3tK0NtGMZwUHq/jPzBU/V+JYCxBVgX7pNyHPtT
od+DLcnMWjGGV5LsVj7+e/mp0wC3qC++0Sj5BFOZAkYYs9XhTLOIEQOI2fJ9iOnN
mOsR2PabO3CL4bXVoneQ+xRCKdcJB5JALzDscGGrvMN6jb/kFKb5z0IqlFyi1nJp
cx+6GlndCAEVpWpO8uWUS+fji4NuS/OY0oJthV0zmmharbDY6Kpv1waLm3tdS57P
h2wsoM7as6okJwRthW1vtYgBfKucsBpBXDIxt+VvN2C4YO+DV2FuGSzsKx7Wb7iI
tdicBK3nikrh8YA/o8kxzEJ3LvDKE+cIIHPpzEBvOM0N6nuJKcP0Q70bv8oynKFW
Miy91cBi7einnWGR4YxWOy38lG2qB87jmXXwllJ+vBBsPZbHdzfcwK/Vfx63DkCS
UBzDAXl1k6B/nhA7ZMgdvGP2/iaW5VJjD2fJX4Cyn7HIL44Dr7/+RuwgoREfUWkD
u1+A2c9F47cF8fe6HaQJ62t2PlGrYs7QpLQteLk8wn0q3kLL6LdUii+IxBcr4KaE
Y1YLejitaLL97jnC99DEkWSt7pCKrrXt+pTMH1/0RaTJDeBpDVmAjXKw+XMgIkgx
n1sTfgXNuSjiqY+6t7m/UaObTddBXteZ/egvi2E+o7I1NuN0lYf7LjhzW8YCKI3o
fH0V9Ygd1Z36GeUZJfbi9ScoSHnapi26c4vSeTKGc08=
//pragma protect end_data_block
//pragma protect digest_block
FGLK6oXrpQQSi14mLjy/njDY0TI=
//pragma protect end_digest_block
//pragma protect end_protected
