// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iQ6n3DNZbMfA8DsHFsPngq15g+c1AWvX3HQ4tyG+j34o+FFDjNwmeAqZRB2y
54tHPKMMGIO9jwZLCs7/hm1kcaeNet+xpZoo+s7iUQxuinrehYfs9n0YZnjT
U2+h5XpRyi7IjGCQqKD8iMD8LFmjkoIMCAVeb/5mDqMqemDH7nrHW0cO6ina
ggeY3rdKjtUIL1uOC5XTt6SMHlCdlX5hUjlhwhVVb6EJkMGOStDCLcwC3Ygn
Z0F9Hm78hg0oAFA0dfMGdndbjudfBtLkL4qj5XaoVq6kqMC+pQ/8x/zxUOF2
WhYYU68w5qMMQYRag8M0xk+hoHEYorkNaCtcHCMCLw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i76nQTgfRgwZTg7uMVayvUt8oJwXevUARkX5VmKbZ30s0amdP+EgYUfzNBH1
Lk2eH6t6ssrty5S6/8WIuQf1fPtP/DxCVDTC11t/Cuz5J0NwvXa5AG87SPAw
leANlmasnMr30puRsInTwbHp1RCCxuwTOW8R9UrKsFjSkX4CBaO0VKJFk1OP
2uw/XePgHiZzeg2LDYmTY2JfOaOa7pZcF85fh/f8dWRS+GUVh1aGtdBjKOTS
YJGBHx2/3Q8cIG1NXuNckYyXIqW2lLqXXNmipdIKNcjhxHESvqq1oIszsd+u
iPkynWKq0MViSIMjXGOFg4LTtaSlbvuvES29ctuLwA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pgw1zesB9GG9yYF562i+ZDr3/pB88Uze2LsqLEBGKtrznI6oUqIlmSOQTN3g
TVGjsEXoP3ij5TbNqlpqC459aX+lMR9UKJxZwFtRKPKklnPjLcUppEZJWiPd
T9Bf+YNpGZSSiOTOQSWxG0B5jkVbXmEv7VIp6fnTU46pRtLhrFAp78oG1Wtb
Z9VNRr/uafYXICDurlqDVUyZ2pwiFd4HeuSScG0jUg3rictpqCK2qCbdAFGz
h84cH+PrlNeuI7P9sv6HBcMI91i9okeCrarc9RtPDEnigVuv/8/4fTD59UKp
pVRfm3TShqljG+/Ybe9Nnw28yyouSA4fal197Fe9eQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KrOId4D7udg6EGDBXNuBmhbK/35aZNP7djwB95sWuZr2XAYkuwQsuwv+Svr+
ia/v3TdkZjdGfSg4wQm8SR8LPe6UP6ArTeMz79vb32hN8aDvdrmTAyN88ZSe
AoxRzUFEEPxtWY3fXiEW/UUewwaU+cW6lEcwkIV4a6z4p9MudRU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IvSmiotroHH51TrwYXJ9gA7KvsxWdBvHvsKpxSE7N1iILbHI8hfW0KyiTQgO
7bOn5QcRxPCS6o8F9zDthUGBnx0dcubK5JIS1JhRwN87IPV4OJNqQtfvKK/3
zC/g2Ubg4ptWaQvXzWjz3q10P9uj6e54x7EzfSNYDBKQsONk/zqXa4re0pM9
sTNwxBQb+2v01gEVWVikOTJO9HXf5PtiAvs1NWe443lebqbBhwN6hiihH/hb
gnTPnv6mr1qMN/MvUAyBgQ/3fX0w+t68PEWq5SgdGj1JlgIOPMUswEiTar+o
SxBMC2KuTfX14292e10atus+8eYFWOvpFg+S/85IBBoKjIXYH9EdKCYZQZ8O
2A9PJeRjo/MhONqtW06vK9bXmBWrggeurVrL0d4WlyKPnHQVMCOF8IL/gICd
KghRWA/qkS0Jw5j1c+lg0JbwrAeA0UKZrHPV/xPgiCLaddZfNgPiVo7WUH10
012Z9ZvkHDsexV0rhazSNmUGtCm7+jBy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H5YnIXW3rZB+kWfOzObtzl2uRAJU6ED9ZLdsKW8ZaiKlBe2V0JBtY5jo3b0V
kLDJE4YeOmrawODJc+S2Xu93KIsbMM2bIUY7KaLcBzB8Q6WNnWOS0PLMJ01t
51H2YxS4qbKROJgwGdZ0XQrTMCdBCAkm7XpX6/WE4SnfWGgkWDE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ukMDuMh5Y3yqRAUrC82B5TvmsE8vFvmeNaArqGSP2vTFJSXs2geemL3f1d7h
pOqERYWthajrMCFK6/Ujb5yDJU8AtUEhAiP+UFYKJTl6sGGEJ9DdPEZTWhme
npGpAfACox0D/AP1h3CFTcepptUXS/HQp3zI8aPTbWM49XX9E1Y=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 24096)
`pragma protect data_block
6W92RPZdcgZY0rOQo+SYWs4n2WW3t5dpKfFd+KzWhFS6Ko3EaYO59efh4dt4
XQfq2Qx981VJU+9XJL7FiWKHXjOO/53ep/+fAS92lPptu/miYVVtOzw2M15h
Ej6ZDj3CfMb13LlsAREmaQqaVBTgtNPbEQVZCCLnFfH69V21HJzLpaCqVIo2
2b/3xN2zpxMxKM8OrH3ptoMEnFLWdGDEY3bmb45nVG2AOfYSkER4aawb3LCY
uvh5sP9ZIfp1itlc4SBacZtjJoaSz67oLdM1MHg+ZRA/pNYxxQlVFvex5Dh3
ysGaVZIyCn2cufLVi9qxpuyquZYLlDyJI4kPtKTI3cHxP5l+nDj8Te/9mvFy
1EyN4kqGs2eqxPz5q9ZE1G0z/4b/q/7A42vVbzeo8NBU7GEy0+z/1eq4tE9A
sYa88afAwHwyzMl2jIsPnrpykiJLElTT2dK6/XZHiaNNwiDX3x3Gxi7gUAGq
rgwwJWj+sOFTfqBp8GKEhUC3MWcppT0hY/sYMFDQo/wyCQ5p+U/7I+ic7BKY
m9dpBsP4RBPpibk90HskRprRVazy74Z3gSQuHefrFtR6zU0JxcVNlu7wqD8E
bnWOLQXZe+Mof/gpn7cmruJLpy0hndVjZ7T7HOxkBYte19j0UqgneqoODbD2
un8ZGliP9W0CNHEmPD78jZuJivAnXO/05xUOVbUxyjvk17FbccjNdLa6YWPd
53Ab8JgjTKZyUaTnFaY3uHuE+ujY17kI3r8uu9D3CzBLhIBtC8kc2OPArJXr
ZkBod7yHfVsdy//MMv9BJ8oaG1nB86pOLJQVqjbSxgggmF/eKn3/7A7i+1nL
J5Fgx+AtWgaOQi7x5oJj5iwyic392UOKzmT0QdiQn2IONk2/xLOUQhxeFixX
qanhBlWPsmdJ/jnCmYAl5/H2KS1ZK6ZmcpTLUFLV4vcGMhu0aeI1hmOzxIQN
p+suJtK6OveOwOJrRYIIB+iB5ANXObXsG4baV05j2SP+gNvjuEjlX1SLIUjl
L7W3IH4DrsY653tjwjHMz6rUnekEMbHQqU1mVF71qEjvAyvDcubgWtOl1QQ2
hG9vKk3HyT7hV5SmYg13UHEhwGE4bWtuPBUzKz3VVoFGG5XgGQ/Fk/EBLogg
WnlG3apfHc8uqZAixpJSvbb6tlbTHIvo0rQzw//lmJrXCOMz8z+C5m6m4hKs
a4tgpY9n83FoPJ6EAA/zN+faVlomucpGmsIN04R85swIOtRGec8ZtOP8HKVm
Wcm7E75KGOPzrhDn8bA65i0cftXOAj2ncW5JI9XnXET2RP27KqqS4yMTjCy8
+zWyR/Zu8UJup4JzEQKQFyWtAg105R8bWHQDwX+P/IhqaadtQzDtGTjog9Kf
fCSrcpcg8ATlfKw4J/ocX1tuQ3GJlHvsI8mYKCirsSHdGSOTOyZMpfQwVS5Z
CqJhhiQpEHMeZshMnsJ8Ym4y+r0uzoZK1vpzJFq89pJfQA4i14NoGyXJTDex
RR5+ASaM+R+Stq+gsXHBkHcGTrsU39PHMcM6AmkIKEqzcRAphiiPJx2GluZZ
Jg1+Aiq8g+9AOHBdJKuCUPruPBU4HqxmiOhArILjBaxCtd0js+CBVpQqhVkI
WfAQsffOdsE7SypvgOYsaBa1W48u4NKfZnv5DGFOcrRwYdueV+1s42TxWTsW
MEon5T+QAFCQbSbzPgB8D2hAMkZ/3JEW5AJ5MN/sPAApMfgQLjivhG6k+qZG
Mx3TuXaeO7ImkwWuLMoazA0InOviBEfHCF6WG1rOHPlXs59zLyuxEF+NIVsb
kfoy7/qw338xB4z4TkJf1YsocCYIFyZUaD5qzlx1L3AsamlDWBHBlmXSY07y
TSehJK72Whx8XMfY8cmTF72Q2vP3MwYEiJJ6u6bodZyM4v3W5oiwMmEPfua0
oEcmz8yoR/taHKbpfUkQoHNzEWoVbxR5HcIBLB5PDLKAaY5UFo5S5bdrMfXe
Zh/9nyutmXsreIRXTo5DJUlyYVSFCmUZMubsTZtJUZtELRb3KNJWZR8HsRB3
kchoyQJ4IEcM1F6vwnDpdh+L4VFtVkWQkEOtlAfTzU/FdlrwfNbx9ACIvvs3
ZXCbjWb+ZJvNnWk6YwGxBxm84HJjFNJDp0EUVHakSwKaW9Dd6Nmm15+PllFs
AZGBb9WXGK/W3WGJy+N8W+QLSxIa3pS3dIapUASo4nHDC1rGaVqT/n3RlMei
YZz04DIx3X3yHs1kQRUcR93ReBiTs7hsfLvPikzeqbnhq4Tf1kcASsYcYyOq
OnpcXnD1QHJDSDE+f611q8uuwThoENf0gQ9buE6jHuvix3qGlqbqIagPBOpi
I/CPSZRg2I0KwbwWNjczr7WZ3uMpUzcfhxZMyK0mq/mOdC7tqdiL7USEwb6d
/ZgZA94pnA+EZC2w7VMb7g+CkMyn5hB2gO++qjppGHz/QCYW2oGSNd/iSwDa
nNZUZNuEbGSAR5JV+SbRgzWANelr4/OSejigrNUD8xxslxhkUcSPrZ+Uc6Nz
cKBOpOPecFtTDcfHrDzQD6qAnR15twCJ6e2nNn55gGM3fqvw+wFHLvVjASkk
3E8Z2E27cNwJJSqjo3++f0Adcmq7OOBujLSj6GykKy3ZBNvLK+4r5rpGDiOp
XGHPTZSByxEIN+jmfk4FxKtTGpfdxrIu+0ppRKZktY9f0Obkfpa5nqxmFMcr
nnTBLuovWtgnD8OP3n+7qltd9bSuheJ2FI89zL0sVA8Wm9kOz1zODPbPBq08
DURW7ars8cFyDvzs+uIocO7aLIq2N21BNOGW2BuN+IrmQ22NKk1isOvpdj4/
qmmPOoSPY1DzEyHJsEo7QkNNdXHc0QFx+KBwdsl8GIWKWGS9/8x9YZ8iVtAD
/beWXg4E1yphSnKySN0s8xicJsFf5m+mMRb3RgOcEwuhuS8GmrXJPW4mGEdS
suqF+67HJABB3PK2Mfxdda99eLQA5BPThDJ87g885NslJNtgaoDIfjUzq9Wt
qVpVllFVrUIz6/PieQZIeD9R3D9PKT8PhrG7AyVaa7H7M2ISZHEZAkG5LnnS
pARqCL760rvfJesReYZdaHKZwnpaosZqmKHpIotlD2fAb/fIcgKcSHGQfqhF
sLfQTedmPGDKxLZLtN7jl2KxUenT6pWZ6FFPLFS46hIqPjknvpnbSU6R3suO
kTJ74jf5F7Lm9s65D2lGP7fTeAlrG7z4iFAy9S/MCTcjdNJCrqxdiFkddRX0
K80hu73UFrg4F8fN3lcKF23M+Dw+pgKk6lZQwWmuZXniFxVh3nTcuCfvL8tg
xApPf7SHkQrt1X+xFGkzbMGTqWeKEZHEm7/yYmT2/4K0rPvOmH2vJJRkO3RZ
XnAjNMxtli5ekh2tO41moMMgATEPa61B6ZeK83EoPeB2ceuNOqkvWiju8+65
QiXsM5G03PxUDhAQaoPhj63eoRLzX/aM7jIY0ightENsDNp/Pvh4byZqwlUj
yOPfue+OcVxSO9QqAwAHCKcVkGtXvDzGMSlrSX5iPIpoalyPihEFvoxJs0e0
i48BtC2j3iAwyJUiEJ/zC292Yq4U0W87tLkzEe6Ucy6iHMKKVhHoVZ+tg3RP
cONfKvlJo9yAjJQo6Z4REUySKVzz3gL6l+rcFJTGFqcTX1fjDNI6BPVU9hsa
TVcx5tblL71mJuqA2h1qg4y6gKznIOz+4UdE8fTSMQ/pEgsH2A6MDqbfKu5M
fJ/Gueb332tVuJh9TJYXlw/huTmMsdhNhcdCfjZodddG2ACxuV4xAwXNx2Ll
g+OUz/zbs9ij0Uh4sC127xjXeKFOYe7vHdLmvyCmEBK5ZSFzrSK5ZPyBOrwr
hbg39JMmGPqi2IIzBq17Nn8Ov6lhBSj7ezoyrmT0X9nOTmffoXCV9MYcrnPp
1zeQj6wf6cE+CNsMXBNOv+e32VkIYL5pXQEcKeEZDruIGUXTVU2k7RF9dfSd
yjLQ2IaBargohXO83l7ZEDIk79t+iB93cHQb86QZGI3R1Vll25dcLctimDt/
BXnTHkO0mn+oRcmbvc8LNweU+RvkdtHr0Ral7Y1EeStwzJgIirEy9fxXsCMV
7g2QUczENHcJuLNkdCN2MW4+2vCg3nuvlIwb6Je+eWSUC+w6Q5qIznEwqFYT
ik71es+u4tDpnm1SKNrdaRuKuvwymlu/d7pWafUQtRX3dTFcUy5H4N+VoG/x
hw0MkPL/jl6iUVC52RKl6JsBIwdUB29orsCm0Mv7LUvaFTnNy0YBRBYX+9uv
genxuErVlzAXUuepVOhkOmo2RDhD5nqN/TrS55AxcCG27+w5Gl71nHolQ34z
S/TmRh/Av4TTmrAKs6sbq+Sym6SXDidRO/mXkVAHg3cuD9m5YqwwSv4pk0Z4
dLbNemRXjDfw+TWAX2D1AAvmcLjviY00gH1Ql+3A76JUXfX4Nl/quBb0NzZx
t3NmMLXglj6UI2zNYDx/fu20rax6N6w8QEqNfJXJKX/qNNnW9LbEV+ijVlh+
1XJ6gAEOw1fULPTfC0r915cHvc+4Vu0kAHKB+UPZAPmbDIe9arYRdVJ/hcU1
EgneUsdtT0bGGraa223ni3bWYiEgTNr1e3IPYu1Schqw6An4UX8miHxp56hv
Bgc3FR3KleqFpN54RuRjDMnxX+Rdwftf7q/9YKV375CcrwLNuK0U3zO3Reky
Rsy1Jwf63Mc0css3mi0OzbSzntdBIOkBuS2zgDGjT/RMuHbBurM6VJytvi5u
rWRsh0yBCuqtgd/290rI/9hOHvaqIZWfNBJ783ZbDZg3GLvwk4O7MJoWNjhU
fHw3hpAC96rpI4MOQ6/xCaDiolFXbHK11NaSpKxtzgnq0Fe3ONFmXnjJTyp2
TIb5z2aG8pCw47jQJDu0mvo+CWOrS4tNZzc3/MLO4Sgdosdwg/QAs6WteEoP
0Nn+kQCjyUHXkd7lpgNZZ4dW8+BVV8weChQAN3xrdu1R2tHiFz4z4wJkZpfp
5EboYuAe1CZLnPoCFDOHukMBC8QYc5T+XJHcOcB64JihvC6FpOT1PZe9sCAm
10Goma2cZmnKMT2x656qaQPGHNpyC+Bn0PuXlUsIC9C4adcUG+XqTP1Kkruf
pBPwmpTZmRGzi9L+PvOPIKcK6oJgF+1moxmfZ044D7N4qQIyCp4k2PlmaUOH
JyCngZeoTOrj3xe5RkzyF7H35jbMvIoCI4hL/uI9o3d7/k/9f/cH8RZTZui4
M4qkbNRFEy9iez8nDG9TCAbq78SsZV0FJ3zYnf6VRhl34hcJZfSMmgA6BZVH
On7CM6cd8kKzb8uqO9MCFFaLSK2mmMgxm9v2jSkMS8cnUxa+dBfgPvpbKfao
VCGifuNQZ68sLeN74n/1r7FvyJed/qPGXBv4LNhsYVKW4cft1OjPL7S+VwYg
+hlCn1eFYJiq/K9DVBYOzuDo7zy7sszc4XqRXHZcq2Np+VyfNqQ3KqvppmUR
B8AqYkUKVW3ELBDODfRyRZLxA6pSF8ao88G3igMEZ9cIAjeE4zQeU89WPqjV
+SWtYyDqOgXdFc8AN0z+hfBloM9fV2MLoLhipbBuBAOvbJL6VOMIgP9fCM6a
TlGQer4Xi9p68CAnfUw+ujF2jr6+GctBkYVf6hdCH3lc1pGaanOSx6ai6wQQ
ZV/bLbOoEvo7ZZqsBHh6owoSWGhpmOC9N8Dtv9E0KBD3KAnBK3kU8PGBChtI
7n2s3d0m+txjp/BEHDUhCbkULvALL45bt3WM1b71ldxPlEgaKgrPDHE6jvTk
SU28K2TiIga6oMgg7XAaWSV4LyddzZvktDy08Z5XWuEESmvaqz+eHt3e9l+t
1tXXXf3DFo5JL3rnGZU8fx8LE/8LI3NokJiN7GNIiRi2fcn1iwwwkc0W+Fb+
K8FGdxUnWyRbmeS6mFgILOSMIGy5TZ1+1Q+TbLvaQ2jzJjh0Il1r9Bpnbitg
XdcsvVT54ctLsUtimGWS8tWVQq1utueYBoprnCxEPYmT/Y76ILOnftyyrzdL
KS0iMilLgAKQNfIDDrVcAUF5Ol7BEzuU4xkTELea87pLIL/sAfd1BDZZcipN
pjRuJbcVePfLfgDBkRr3YatB+NwKHMWK9+/lDtNdkUOM9febNeJoA0zBZu+p
+1v0OsMVVolJr6OQEcIdxSNuMhYHZIS9jLKz8gZsDDXazuTzmZ6FSQZKXhMy
i/7n/93RZRxstYuTuaYeC4NNFgPe2uUEuHX/UNCuxA/GBjYLAwLdsoADY4C8
gzVkO6QPvzvQJH+9aakJN4fQKeffBVNKtZvUeyiWqMvVnJDyGLhsowdnWD7j
gTI+vzxO3KTEUPfAkTdIa/SbG1YZSYU2ElszAReFM36dczW6/98QLA3x6mKy
uh7uIhZm4tH8F2EF70Rx7HjsXjpQ1nftBgrqCMHwy4b2ZxFvRRYvDVTDuVbU
YRN47BEIBvVJtbZpCvOlJVCgWzemtGxzK4TxEaj8CRgfB1CmMIDr/IdZHNhL
naR9nktKL3a6cOdqSIXhxPGJrm0AVgIZ9TO/DD2siWBI9lXHPnzT4KKHfVOI
fRNtcM61pjsHl0T52gPo+xav9Ubej6k+lOF+ys+lLhY+gphXrJbpCzUryM/F
93ZG/jthVDIoahATEu5MA5XIGap4CoP8Obybcxifpvav408pjWItsZeQURRi
H6ijWFG5r2wEooCYq4FCVkzP6/kYhS2WWXUiImwwmgPwiLIqEDG+wbF2g47F
f/NTmRFgCPG3RKdv0X2tzgbBbwYZre/XAJna5ATXzd5xNQSnkfbE7u/YXrvM
0998M4Vnd/GC4z/1r0fTnUKDIdl4lK1iFyIGDKmtAClktK4z9TtADFYa+7tb
t11TjGL4hq0HCQmOYjTw3LW6VUGQIwvxWoLqjS9xzK3ko/9e6MtpcSPW7weY
T1CfEhoiqyXojA1bthzocj78fPEuzM9NlbVeAj7EwjB6kkKKaTmuXuyblevQ
Kb/483fgWE1k6/iXZEBL0tvc+HVO/iJDj+dgOE/ThqyoWCEyyqA4xiADgXCP
qEo+YB3C9qJzT3kEvmykWLL0FyrFgN6+4euIOayzdyXah/gmWm0hrz1WY+Q7
O4Nbcrh9RxPrmycId8BseB5FjEfbjLylU3PmXzpKKoS+1SgCz57oYLRNH/RB
N0ZTZrkqiToWvRJ8hJ8FUP0U7YNbwDYXZe4h1D9LlCrtrTwKp1g7RRx/khc5
Lmp6ltQVzP9Yb5vG06XqGoHMiNxtgw7pvQTSuyG6SXon38uSnIVWGhvW8AiE
yf+sTIXN0lofqHBIGyoSt2VokVUc0c2qBfgUbZR+PMJ5Aq03axAgXSxeA7PP
j0cdY0UYAdI0xeSg6ogDUdBla1Ww3aVq3QUFQcDaaCC64nlzIcXJmiTtqa0h
T6H/xPm0B6BdadTEEZ7nxqZDAbsoMaNjtr4kgnHA3G9NZ3k1J1YjU3p1ZC9w
0B+ZqYtlBczVpKCV8CGY1uuLbi3/a2b8UVnjuzdOom7cUg2mE3Cypf3+oifX
hRswy0cJt3IeUVLJtftq9GHTLAsW4THxRqWRXmlOwMZptPZrFPQ9PH7XkDgF
qWK5PcjSjANY9NsmoyVzN+5fbLkPlhIcJHj5FjxQgkUQT4SIWZPTvLmITRr2
hs5ApMxLT1qiaozG7+YErzUNpWZIBuOVu9qizfrynIxkLOHOKmidlNnKpXUC
VfUbZqqAkgt1DAvxThjHrZT0CmQVFBJ0w3u6c3bq21G0R8ze1N8qE6RQPLC8
c4o5PGsjUV8SfIkDzmhGhhs2tSXHCPlpIq2bGF7exJkKIVnqDb9K9xYC1Xrr
Zp/cB0QcJ5Swq3AFxLjWr3qObLYB7K00+DGrwBuMfvdnnu9oCZ3UvrtIEXJZ
k4za6V90qn+bAFE9DjBgvbASeZ+f2k1KgJJHRcCpBNMd9ssosfFKYYpQwQQa
/sh+u+rxJ1jVZTvtMgSU2jbZedRTIwcNrmwmy02Njp9tvYH1Pvo4sWH/tBPe
Qctpt1vNAXYWG4xMjvDQBaFeq7R5U/i5ThqTj6loa4NuT4cnvKQhxT6CXCtJ
HmdbGGVFUv2TbYAWjbciAtLhUrbL6jkmScdmqsKX83j+e5F1Yd/0cgpPnYf9
18Qe9N8v5JJH5su0M8+wxWVDW45raw1NVAsyShW9WMLJ8xhYUKYo2bbjG6y6
jhNrCOMQ1bPIB0GeNyJRYerTcjL5Sdy1YD0LpscOAYP2MRwAC1Z61FUfhwcC
r66qvK2mdO5sQlNyAcSmkmEHlkU8XIML6w967gihevM8mD6Nhnh7KrbIYh8m
mHv2PtixiUT7656UB9Rnb7JAKfMUhLsrCdC/FPyYL+9ilQkY1gG5YV7bnLl9
0WdOfB8yMuj882w6Vu8wTnshjs8W+IB5W3IFl3rfa1jHnaelmyK/Y9ovrFKi
chXuIHYb9+/F+8gPMcKkSroLpZEf1xPEOMHGufGRKrkzar93Mzq7SAJSGiWf
Q6lx5pNskifaUifeurAnNfLECTJzJl7bjv6+7W9DG4FY1DagGw/2ysAC85Yz
febMZAYgg+isWdJUFijPj/U4hIDacqaFv8cswdKeBoTlduxzvAubL0kv4UXC
PagQzYTVbmf4/weDN25H/fb25nIJrsde4u3KXqYMebtJVFOwLWm5HbCxMeXk
YUoYiTpBz7BlaDKkvf4TJM8brln7EsPd/8LVylctC7MPZbXX5VAlnoI8LwzY
YZEuQCobLXiT13HikqNm2C11XCMl5lDMd6/qq3jIPZYvFY+X7YQOSi+suLY4
LPOtSQwM+ywDGO0UY5/p0SVCEvTKYJbYwwAxeWBVierewNaIseIynBWZOTaB
OKqWGs7jo5GLrxBXAD5wrLkFbJvkY5PyZw6NSeNOgSOvdP6n9pGZ18P06O8n
eMqKOuBQoiSpulmdUv3k1oSLiIqY+15JG+hdm+6f0RN33XaatpqV+tyX0Kin
b2sGqxeV8/2rePZtWQz5+g1bX1623HNmbGH5fwsPE3xhhBKDHKMadfUR/jv1
AhwaHJG4+XYlhIa1Myd9BLhTKqBKLVQOhW/8A4Cc9dlp43mK8X53+u60cKJC
Vf06H+9iU6JPkpTKXDO2Ne1qS6mevptez8hEXUb4A74eCIOXEoU54UhTrM3Q
rpFGDurmApOnIMdQwKftqrR/YQ2XtqqxNnElzv9SOqlG9sl8KxrPO5HHOCTI
0xXyt44pfPh2PBTIZRv9AWiR7QWHwRND5KMo6n7O48DKe6C2tYrtD0vclcim
bJEY3ys24maBGoaNPMsioGUaBJ2FF23n22F+oXM3JE4PVtSiABdFbjv+Rc+C
TE+kcqZzyrNrSpsWWIhr17PeHHWw+msalvMiIhsTukmCDFscBKNqlGQ/IyLw
sw5/Atbr4kBHSUTpT0fF3QnTz1mYUkMu8c+KXMxsYxq100bVzU9enXWoALpH
9woDRoRROHQAkJpPF0RNElZ51R9QVM++e4QnDGdshpqO6vreSQFRwHqXSBaL
n9lzK1uWkeMrLFxVBs5RqoWASTDfUv7gdclkb8Jv9N7nR9JpbCZkWo0aUZDa
SQ158nlBdRJ4Y43t1Oo51vSMqDOBBawJiWNT6+1h6WWPDSRfp0lI5uP2TWM1
/efnH8qaBFcy/FCHQ7ha3aqG170kLjksbkQfOAIERthr4/mt+uuvLqWemP3T
pnzPYx4UUdh6iz9WXrxQot4NbSww0W07WzLB+RL8+C57cOk2V7r6R69mRFEU
XWHTIuYNxOQMMEkP714biCQH05EtTj356jno7Ney5jLq581dDNrmyKW9TAbf
J3w9BfM7kHG1wSZUu6OUBihbXNn2yE7Z6R1o2ZtFQxnLGkkMHZzt3A/CAgFw
R4dXgkcn4UUnAdGlfk6CXMMMDWr6OYrOwBfgLMgfmf+dyqlkOo+Bg8UuHacH
m9kUEkiVJlBn5x6zd/MUH3N3apyiO3QL/SEOB7LPuaO6HqNTDSfWvEpO9wh5
Fl2xvKi01ZLYmsNQKYlV+72SH36nqkXyLPuUej9XQGJ9d/mTG8BluYWkm78c
TjDNLUEV0f+HsUfPKvb5z0vo8QRs/PcauucWMCp673CzQjDwH+tguJw2ciMJ
Y1Lrma7OwkMoY8hz7YGlA1lewFLUFKwE/D7YkviigAIuGExnT724jX7zV3rw
kYpSvUTwOUV87CGNu648I/n1xf6Mx7krEslhzgFxwJWTKJhbFXIWWhzMN/pD
nefmjqgdidBN+kWFT9yWJWJYJlR1JpCyUa8oK7g3/kRMzS6THzw+gHSGXBEJ
IzjIt6yNHtdc7TRzTxn54dGXEHPDJwvQgSjnaUebnhqnvOU3gPIB6hqzIkSZ
D1ug3sCdZTORA9/gR2xdwudYN6vK2n6x5ry6SyCSMLLc7VF8EHPS49hDgpi0
NxYqr7Xn4wLmIh/GeCUXfUVSDtcU0K2mgbnrDy8SP/93QPH21QS/2AMuAC3D
R6ND4YAKSWqy5ojuGPzP4JVMB1jsnMdJN3d84n1FON250nKTE2icE1kLQBpW
6usJum0/Lm6P+EKJJplNqGO39ISBGpTIZcBNgKr85Oe+FdOPrdu+LJ/W1/tT
AYONhRYNnekB8j8IVeqFBUjOVOirG6eEezHDpH3+ZzDQjQevcE1rfhfPZspF
briCSi7dK2gVelORsk0uZn8TFIsexb3ROr1ebNcNqFPHdgcEAMPt9CdtwXxJ
VpzHZmXs0edBjdRD4lTLqN0u0i2dV3W64e0ugKDII6QfDYaLRu5i5GofTeRF
1n6XPUZBd6nIQTpCyT5m2skcb1wWgKTyuZa9b11R/iw8RHAGNIY9p/D7COpn
FvqiAsqOOsYWPp9WazWtxGcFtcQPsUllTGSrHeKLjOlpCsM94Nr2iNBgVw62
jdBOfMpCPrBKjvdzFBz1Oy8BjyQKs1mLabEHV8U1B+IomJcXY3BtIQNPgBs2
ubcpHR4yToc1HlfaH8eE2EKSIkKR2sr5j+hxSAdJRiv1oFjYcHKXYHnSDlyN
tsCJHQgooh9I8pjwrBitHz4iSOu3JNHE2UFYQ3SeJ5/ZVdVYsZAzZFR2nbkS
0LvE458R3tDwziTkQhsZj3uXR+6GA3qKG1KOxr21euiV6yS0CeLr3V1QQFF2
N1yrex5/wmsANq5hzkFIwVBBX7Obtiu68/SzwyZzsjgtd28VFSgeIduED1VN
NfZNEH+5fLlAa12fyM5gLoOx4CpkxAtf52eZVJPTchIXUlEPvsXB7xLKrxCz
4lHZGf7AfaO+1EBE4Fk5EmnwX/EdhDq1pAwn6COQYffT63ACKMJiiYuaNU/C
JuvsOrIXKEC8utdWNGtljSyrRKQB9M/5mxGp2fjSesj5xADmV1N6g3uioSYi
lTHAUQMvrMmL3Jr86ixfSkTKGJHMAfqfHeEQLEv8XWzvCzr19BtVf679zfTP
lQsU4iQbV+HArghjhZB9ntZziIMjexxU+iX02IWNr75Jt/UBMqB1BJH7S5J7
Tg8eRzFupI7iGvnY4odLfnXY3xfuQBRtmaB313xu6URFB5HLsa9T8RT6GnHU
dY+YuW38fbVnIKUiGw9EclFaZq26fa+9UWA47qdJTMktnaXXhf5OfcBVcKh1
VFm4e1sB6lBsIj4yHTDVtLrugMmYl0JW3lgTNxKprbX6PlQsIIpN/3bfdu6I
C6O4dbs9IM+OdVbSiz4Nbexxm1e5d/uV1m2DgrRpgS0BarkDdLsJwm73VZtb
BcN5TLxER9iB9yDUqAAlJtv1tjZQNn2doebMLftBSWLe5HubdmXKOkML3YJG
GFwtdGd9na4pgEWfGxEWQqRinCaFIChpeAc8djRtCQJe6YH2Qs5bUxtqHeED
c6rmHM+ezJYkrV1ER21i9++90iuBIAV+LEl/+u8Z9TGrQ99S0O3zEeQKeY7v
jLlpM9Z9f5mElsSoB5gyl+nY8Jfb11u4DooesCwip3a/kQZ0kmNcgbLDH6wZ
cVYwAcg1+p6/IdxrlBYVuEdeO+lDVIn+E5/I1R5/pJuTN3WqJicbrEegGOuk
RyHlKAUwcwb07ImXjNHcz830QHzmAA+fAVRK8qI9zJGneLuc9OVICHaBrZjC
SbNu00QVFfeegei4dCws9p6h3t0W5Arj1RlP8qWLsQw22OK4HrdIh/k+Jd58
RfIKInbbsLbZMAPOiYvJf79StF+PcrlNkOibiTURXzDVP0Fiz7qszL23PG0G
uJ7ocVO38ch/XgR/XHh9O1e8c4Ytkgt21xDtIsGLba1ohjqyDjfB3FowUOsD
7ug7OdnJ3n/RcDHL5t2u8h3SbCvOmGvJlIAiWQue8VmGHJq84/knLmIFUiFy
mDQJYWANcUz0oI4hOoXhLRfdWFobMmoUYBAa4G8UpWi2xrJpOGbBIdguA2/e
pW6BGOfHukK3zzgNUDbp6Y71hB0UfhqDV3A/lupXWoc8PCTjSE7SlbIRmcvu
kH+Ig3I/7GhZrQSxs6oGuT8sTzImY4T8s43BnMBXUVk+6a4+9bsXgwUyBCaA
e4xZbIkSw+O4FeDsEfdsEfwQkREUYrHvf3brnJuHHnQ6/QoRajj3YrSrkHPZ
Cjqj1FIePjOupZHFLrJTY4F7PLorcndT/oMxtaDzqMF+n21ulE3r9luh+7CC
F2oMeVO9uuEtYozezJZF9ZXhzNA33NNpEAKn20riPdDf1QuYhUmZBzsS734i
GPKR+qd+5oHPpl/n4DHQucBMjdqhiMO6956+N+rFAIKlqgX0s0saOrn1uboH
p6fCPbgQIGvrlxjYFOqkAjwrhvphZUkXUo2AK43102p4vueNd9hKI6szxVsl
fMbnGPg+DwYMsLFO7BXwEdCIjG4SYyyEZe3OcAOWSfRyfDTs7BU+WS3MwNyJ
5ofzKIgjuUgIDmV9ARFu8dYIOCOeg/EaIUmfDwis9m/QSZ0d9/5ns9PLA/yl
JiBflcrpQsP+YaPYV4UkF4Tfcm36zhiZw2ywPDkAkW6qUOkaREUEZmv5ej9o
KPpVaQOCBUtmVowSSNTI3PVkh2KhKNXMqo8wxpd4GmyoU1cDr+GDzZv534sR
ZvHJVdu9bw7I1jOd0izGAYzvaZ6B3HOgB8CMWIH1va7U591KKe1/oi57fZEF
subvtHsagEvKB+jUIXDuYituF9dDVA6nxs+eaHxLJ3cdd3x2gy8vp+HLrujd
MsIjH9VeaeCj10SIkEcCy+RBqIIkl/rU7Z0fX7jfvCetOHsg1/fSBCFlmy+U
aafZ7TAajNJzdMmMszOe3ha8NkBUIJcl2AoUcCg0IpfF7kMGZ4RYSUh1f3r/
lpoTAwVGgi1ZZAttL9Jq71LG3V0+uNiq76Y2dHphuvH7zFe7twaB1lbNXO0L
d1oRE+DvzohPTs2gKvN/mugu7A6oGe7MSTX2SU/tlzbJf69e3i2RBbBrm8hM
UidB9sga/+YWO2YewSvWRLmfQSlNPW2OKDSsDhhzho04UPammUkWOccIY3Rr
fhdsYoPldDygp9Wy+21AG0JSu/0YZ+e7QM8haHPZVFI2en3UV3Qu71zf2Jn4
vL941omMNjYrmtwI7li6vihlasw3jKeqrrxDX8AlAPRqtJUlrcXEkwGoerze
3y3Tvsf84Md5rOup6jzIzEQZmg0CZZorh7izntf7gjRxBobTqmSHUFuJjq1y
+iLc/sKvgtQ35Li3O6F7GJGHmAoVEhdJmpELF9N1tpF36coRh5/5mBy4ZPZe
TDL5yooV/9J3obV14Fb3UwJYyFrcgReNJ1iBXj8zjwKizBwqzjrOGF3MigS/
vFxUdJ2LgvdAEifaq00gJXIYcpeU7JMJLK5HjurA2QyQJ/L1HhKxbwv8bp2f
w2e+CNYFCucbKBAGhIJsjVjPVt6SM2xgcjxqr2TDznmVP/fM+fsNGKp0V4N1
9SdxXLvrvYDgzeZUSMhnsRrm08eSrS5th+eY2/4x9c9Jlz/DyLbmdQlKxlL6
WgEq4VVtz7iDrA58Lf/afeQm6jSoNblgTMIBQ4sYEBwypu0MGoUlX/H8/wUx
dJEyikCcnFq51k6vUdxG8Pu6g8Sody/RpXIUzzajTvYfwKnMqpfuoEiPsNzq
eyXGi5W0WMVk8vvz/PWFFvCJLEHrKyRQ6MbxQadMhQm5YozkAC1eVeHYub+y
R7LRSEHbniAttb3QEQlSGavvKmZA7ZRWtZrfwXFLl2ST9CtCGWc5WGqYajjv
/72z3tKdCCEYIcX7ybQM//wj/Bo4HRavabdyxv9Vmuip/03KdygOy3dZVxGK
LIp3CrDDfI6kB99BScZAWUhj6YMiGc7dYkfd8YBZ9hAOMzU0DI3H6b4V5duV
AjssDoobWobSlKhYCVG/wm7VO2b9GhNjOM2Dnme+r9KzjflfzHGppKKVNGlz
cKBjc+AHbTnJKKBPSccANs2k0nMVFxx1lpKZ2MdDLAHd8siJ1zuCCRO/SZEM
g3lC3HJN7WpLPTqcmEUOqud/qUwqNTGSI7An6zMG6gNG2e+gWg15V9StjtMZ
a9joqkGcvUtcrDr/9NOvsuCOsVL+7bnta8idbgioRqYauVM3qGbDnjI0Rjvu
zflB45/kn+1wiZUVh57q9VaB04ZrzgooZZbZQOTGYLkno3cunEbAx+CrOeeA
/E0kDddW4UhrKXhZXdfArrP4GHi7cl3jcYLwNZBsipy93SxHmjnlJObrQDqc
MBbGOR4VlBb2+2wKGNNd15PlJ6jnE54qr/J+E/BS/p3/42tXWv/lynHMs1r0
KOKOGmyJHM1VfKRcU3quOPeSNr1tFc/elxmtmluSY39Iw2/E1kF8hzCDlzBt
IF2kmdOweyC1h7J+hayEhfPs9cgVfZTDIpOf9EXNJnDM4z+J6a6mrq6TxlQN
vHEsa8LwtG1f83uWyE45AMNDusikrTueVhQ9F+gbrSmZl7LZit53lvDYI2XL
XbKoUfVkZXJB3p6TBhtt31emXsWBAj1IUyxF9xHguK8dwZ+/gZjbBG9tW3dg
3IPIURMg+tsrXC+m043oRyaLa4ZeMJqI8GipHGOjKIOPOEoQVQDlOpn5cfLh
MedWg5g6CDShV5YDU3cKUKi4XwKrlPOtTjNf43+lckwbwh+D1xti9Bg7koVq
Y7c6BiQNzQTHH5bbcaTVRmBCeDu/kGY7/lIpe3c9Jkeemvg/Ut+0qad/PxGK
h7pSJ1xhBw29k+HtZi9eSA3rmKZEjr2wk1Bv+W7gSOxRAfSqTmopirvJtyHk
f5ONM2Z2T7EEmlSWBCycaIE8CQNmYkulgpB6k7YzmC45f0+hbzVEdyO5jNSg
ffcLKoz81P5yB1uhdiDcwwgdJHIbIZkgciNcx7NGpP80EdoIaPvVQ4cH+eUL
GMQ+eDow8VUedlwz6rbbhTmgI0y6HEBNynRvFLBJJefAYeA3/ZWYcd/nd3Xo
j8RLe9oQeNCu/ye+O+b1Iw+WpVICa1EKB5aEhgjFS5DbFoIn5SGCOz5WY3Fj
Rt2z4kUTJ/ZvIkmTRtbfl3tNsAM3JpqpkX64hqGs3sxzELSrKHCv4AK02Cm9
SOvQSe+qacKECdX9LXsfbkRhPxZJG/BdqsxqHOHAeDu2JCDL9evcY+MNii5f
eugkccBKTRsVfKBmZQXb2sf/87h5C6shgZT7vI3dZvMNZP1WBdv5KivTw2pA
K1YhTFRnYuLF+2WwZrvjxgLvLDpRuUnW2cF42ZU/lyB/XVfDi64bLpalZlH9
cCChlc1q8UcYsmynOV3qJwCbETvgTmu2GTcgkiYTe/+PSW6MVTov6g8NnF5v
CYQM6fPkj091pyjCbS5V4IYYLHNBdUnfTQOnplb6ewA1n+aa/eKTD46R4bOd
otB3BjZXsYkxRz/apkVpE4ZwTkRoAX6m8jR9bmRss6ejBtOrzjcdNWQzhY8E
siqpC4D+JBy6By7o7bBkQ8CSwAhAINBEUGMp/fU40h2QvmPdu00wtgkCLRcV
nkJst7o5IUWqv26yG8xqrIHp3NFrTbPgQ9rPLB8Gs8EYZn8izIoZHiH43B8h
9MnUfYrOB9JSRkFBsCX0o+ikxWs1sdmmn586yLS57f7rp/qSCeGzGGqymyn3
WM7LaFauKk6hj2Nbh+DYswXMoEiFJR02WZ88ATzLhmc0NPA8RmRwHCDirkVw
p/2+h8jCTPmZVDbzr0cnxV6JRoSsYoDdjj+1lkum/AEheK1obKDNfpQee7af
3SLQ6mPXSyoSh13/lRLXnkSaJfE9JBcfvIDLVxQwdDPqTXh9SBl4DwXWr1CM
IU97qOEyXzE0kVf4bn0/uXrTeBd8RooKuvMt8SRM1Lwo/YkVCgyQW7A8g/Nx
0fZpw2P/wpRJGqlwHGgyAPz14DTJsU+EeumRPzBr9Sl+adywtcK16sZ8wa4c
neEUXbreJAKU++ev0Gk58zCD15WYcaFYK5BlIu/aicUS/x/LqQZhefIC6Io/
98On+lZ7g7N6kgEDQ2pZ1xP658NygHcjlu0q62oeR0BSTMaF5U3VTmT3TKuB
5W3riMgp2biYc6J/sm7GFmaMnjI1KYiYLqO9vJHUpAsZxUxYBoBOhBebsAA0
XpeOl6VL3qkYJbZMjVhl5z0J0kp71o70Xn3xeb2v0j2pS9L97WRMkoNahHSy
XlWzoSjcP8raspNqBMbrwHyfyZjvHXXbxU42rJKIlNigKXuDLMbBY6h+XWEi
PRmGbyoHQ785ucQ3FoWo5aBwpkshPrIJZIeMBGo6VhinXIv1SmQ1piIZyhpY
gxs1mWWsFR0K3HdliG00l1Y9HZ0PUCnwZUadhxwyaNw9X0Ax90cBKFcGuygI
J6BG71D5SLytxGBmJFTLjtsJ4WtsjN3lm5fMDy9k75lVbgBun7Xi1yIIqx8P
cQGzv1CND5eqIv+4udJNbU7837AYUZi/idg0pUNTIs8d6Rle1OH9ACJ56JvN
eoIOM9twLaJr6o1o+GbXmFDEEROW+WqTVzVtSZalU28kR4lg/i73s5IAHTTD
9S3EI4gYUsEZPGWzbHUVvRWMtDYfAR/Wraa5dtQM5MhwLvSDE/EnQwPYrm2y
btha+aTRPcog9v4beCRQWN+qfvfwF8EUU4G3ejeuWRYz4WGF5WHV7irRovgb
a0r1EH8nfsYk6tuVH/4ivuAQOY8/joeqyE56vz4v1BXWmuOYnnawYGyYoydu
Yyp+itAug565fKNggdbND38eeFLMEQ9zzAVbr0wENhoW6w/F+fkeK86xOhza
e4Jlj95DnOk5P/WnXrlrri1qqQvrDKxVOCPrQ6f76/gJEnaBlkqw0KX1h6WV
942IIff47bVy5nygSHGo0iD4CH61ztx5plas73/DPT3Ka+hC6KSkMLh9t5aT
uKLlHi5Kbm3wZZ5sCt3yMUlUQAS84YgP80uUqs0H1ILh4FzDe6Z6ZCPB7J6H
tA84MR9MiotAKfH/7i/IZcsZBphuRzHxVgSwwMTvAxW6Cz8mqEmiV2Pf6DjW
c9uSgfC2QHlSryD+W6hQu6srydfK4SLYbbf7Ez85xjkuMMEQBIAYa5V3LW/q
DxkEKcp1iea2asQlVDZ15FwcXL1Ij7AD3K4/KvldjTUFZAZ1euEWG9USPFst
SWb5/pKjEj7c9DVfIapWs1L9wR4KMPFMiAi0ud06hvV4n4kElcRQl/IRerrX
Edw9PIy+4x/JIgUrdBdRQjMR9delYsF7tM/+iOvt6AAoLWoV2OUTJF1MMRsN
QHkyqkaijLZq6rnHqe1imghKXhuvY7Y1kO6GjwrxBpQOUTU4PQ7aXUJ1m737
RnyP7oMBavAt71A9tRN8UKl2DY8108MjTxe9F6cAPzrVgEYICnaP1DL52OGd
VxoH27VACNqsYQlmPvk3/du4H4m/wNm6U7DJ41W/9iqFShGKv0xk18MuvPgw
9IHNs5OyU5/bXQTVE4rZuH3E3rtwNoyvYoYBH6C0CpyNC6Qym1Jxod/bObRK
UO1PetTlJxdYrjSz80ngvR0Huocgxwp6y4DbOb21XPuyH3avn07ISatAg+A0
E/mwQM4H89ei+FmIPUz60506egGlpLSZkzLa+/0bb+WA+OxgIzue/TCuBPKc
57UOykw5uTVoREr7tzS0reI/7LxBiwLTNbu/v5Dg6wLrHZpt8XbvKXMMuvjY
tyOJUo+AFGUpWVH+SsyFM+WzAoGQNqy5q1O5e8wn0xePlEBK37XwD0W6aAzl
kHJnQ4ruZolstxMg9kVri3o21AoeciVz5uDNkW3Ukfay6PGrfjPd6Fr3EhrZ
Trxsjhn3OEmXM669h/jI0YDHxUp9E+FF5kYShBGxu8rzKtxgoSrXaQ9mZFDH
W9XtAq/ze8NIpJbExeLywkK9AosfUzhHNjXYbmGoAb8zkWlvvCNelXpHHtwL
uefGk2tD9gt2EANG2zNboEO3VBAjarGZVKssW4U/wn7Lj+0o6BuQ3PfInVoD
J4vSPv8KdVJRsnoS0lmKFl33xWJIGOlaWYwcDaPUDhj6AJbTfeY13Ahjojso
TbruGmWYC46XdINP3IqwSKQU0GEbXiHjNN4eqB5lJ2xT1SeThFJeLbwVRkly
Wh+EbMp4umOzKiekmcpeNmFyE1gJ1SzhIeRpCwnRezKX4lmauDbUcTz0GAHF
x8UustP8MVeHwXH0k7zyZAvKikxiBKduTwoiLz8chYhDA4W+2/Izj6czd7VY
DOCynRlN3lxT6vZR1qrPvSmyhyVwLklJFMlQ6v9lnknV/W9nvnPThOUF153+
UD+K1jlxAiCFw8LtI85gahHevkVX++yi/csgbZOAxwE0cMikPybnP0k3z2TE
YkdUj8kJ45uHPYvxQi//esYsjZ/5ceK8OZGxvWHiL3n26tvalOTmuLkex75e
3xwcKKBnHVeJEmyMV5IkN3pQgZxMzYwLJmlkPVN/yXumlyJoeRBTfj/Ftttt
LnipOQv5RpUqh7gUJQCbox8Zdw3GGzRSY1CBSt+RN5hantZctUlkpfTZmkbi
TPv1379F4e0hr3Grxm1PeLOqrWHFFRQ5McLJnOysYqiKco4WC5aQ35ke3aBT
wCY+lJ1iFzEWuhY/RSQmHL3Qq+guxGBsBYhycddORwnBuwucmsVnFAHVydYo
ZDivaA7ZhF28POgL03aCIfIg1rskgPQZsMxDzrT5x6kHut87nMjRNIWd3Jcn
MggVMRSxjQ3SM+oF8zRyzxd2oOEWEWQAK1yTfV8hEPhJqchEw4bigIneDM/o
00C4SoeXEM9XJJGfeyS1u5zIRYLzI3pe8bWdV30akEQgChj/DrY2LxB67vG3
wsjk5bWgAXbLon3k/9QbTlcj2xRm34EHw9fK6ZHKRbx9k4XlR0vMXgZuqefr
9eu+PwSRTGA6Pbxm0+GHAp8H7vkhoHHPr+Y+BsYIeRd1HmbDf+sBaUZ2aSzr
9zKx5UXyIfwiWnA67DAgtn3kDfaLmtJ4l3d2x02OX5OMPPwEDyi4Fu1Fp9eQ
oSUt87Cs6PTPktcTqiT/jhuFOI8E/+vmCwGw2D5fuyjExuUngE3OcScyaxoj
kWzTXbDNfBk6q4/OU9c6RmFnOaqPetqoZGd2rGiZsiAzgfwCut/rD6Sp5eEt
bxE4AskZu6kAI3jR3v3tAzYgyclzw6XJEPfppDxbtacjWkopJQQSFSRxWc33
+sAaWKWQPR7SZbMW8fyWPDArxqBI7BLGkktuCAkGVbLuy/LTokyTeS/9ha6j
o1pdMF1azDKRdRmfmcAvX90qz82hQwCFMNk7Oh+Rb8NSYyM6jWsAbugmAQse
f9H30lgral11Kb2juEBgm54WN87e6oYMIZ1oFBahs7P2GhG1ZL02g+gGqIFV
ak+USkoTgrgTF1uOnlbeLBvJjTqGy78NHeB+1eB6dlsX6k4jIJ2/yPHBwPN8
wmqVseW2KaAS0sHCDrfy9bDK1VwgyXQ1Dxx4MAdDObRBk/lBMXtxXH8mBQY5
SUGdcbc75BDEqUgttXNw2/ukbhhwAQrValP01o9DozG89vxox5RJmdrjrrnU
u/6mZ+9dja2Xu1S00gXXa15T8klAPrgjeAxID1Qv3xUNyNHWhdFIGR2p0vQb
L1fdGcb7ExGblwZ63qMVj7tt9YuITpliPBie91LdW5N5t3WwE/fIyafaPe2y
AIUwZIMVfEy/csv2JN5urUkFsEGlT2FHXSsVTCQCT0/lU0+p8+eBmJJ9WEEy
l60vNJ6meCDgE9vXJ2sFEu8yaFnmaN+GcMOm9Kcud4S6RZvWFO7dhlTG9sU0
GxPATiSrAFxOPc0yuenc2qDfw0UEuYUgQPb1b4d1dJbUsGBcQgcEtMoO3gY5
LsB7F1x2QbxG/0rv5Ef8aRsDj4oroczBr17XuBOWmQukHF96+LdNy+m4DHx6
04S2vDue5XXYKZezKbrDqneQzu7YhwHTIUpttmQe6YFNEquHCRbkYUEmRnf/
VLoQ8F4FjEY53mRx91PxYwOcokHWihgeiKOgsidheSuua0iVvt4us3onrY/u
Dgyq4sdh/1NRAGekinbZE35AXI+rNaAlCDCAlPz0M565iQ0/H+8XwkX8OLbJ
/7l7RuclzS5+JozLKYS7qEY0CUODvr/E+tM+sar3Kjo4jTlfNzcbYSq8MHTQ
vmVAGh1CVsqRXWkcEKLy74t0QpYRjqv+uoOKgRIjOo42tc9KTmqmtKZWENm9
3HEc1cKFFJvqpHtmfis7uiB4dsWzYOe6xPMsBBEfk4gVc5MEAy8kZKJ0yV4n
c34HN5qqFlmsAwnztKwcE32BClKbIqwWrzZbVSIMgOqfqU0K013yst3qPqGj
ru6iydkt1//8YFxlXYTjG7fRqDjCHqyBKK0+cZKTJPRV+8gFtExeYAVkjWVK
iiUTR2tmJGMFiXv1lTALx/ld1OAFx1x/1vrfDSFgmJbIKpu6oEdMNUO9uo9B
wAjWPxv1Mer+9eNB+EhonMnrZzzUKmclkx6H7uIkW5kfrZJ6LStFSVRT4ydf
vZ+0LFtVxxGLqEzoPMAcdnrusE+7L5Ra1STFAGmQt8ITNZ1ZqlHDoKo6sl/8
jWS73bNUQTV6Q/vG4sxpVEXz5tm+lkYEgFgKrolw/6JVQz5CYqTgy7itIibT
gQ9fZWSsva0a66Tnn3NPfzQCD1D64CLb7VhJTfo4/wBUASiXVAc+ygEqnX4H
dCEYBex+2EX5YBDcqqjWof7X5ZC1OQTbuR3sJuu/t60pZ5uRV16NftUrYPza
XYNqN8R+hXnEPR/d7pstTeMNga5/OlpwLO5YKsO1vYTd+1KS7mWRBAWZClV5
pd4FDlzRHy3SF3nq9Tu9tI2x4RYutLpKd14Aismw+/AMUAMK7BZoUjjBQ3QW
GOwUN5m6X2yIuluVG0Y5qqSPen2nzjMZl2NQhRDftrRpKbJofFlpshHnpOy1
xzxd92VGVG3C6y2Lczlj7suyXCkaI7fOBaWKw6v+VS+LlabsFMa/Es9GQUOR
FGcLiqyG+GKeKFkfgAjb+BK1TVXUI+kcHBSMnnTbZEAWPKamEkXgATjeHKKt
3FjjFhh00PPBWws/zzGyF/TTAyYJyYsr9EaQX8enY4+um/Ilqd7/niMMJfO3
8wOgvG9W0CgkHFgERthkuD3D9mP8iJ6DGj7h2PniRuFJ+gzuQoKkDCXxumBY
KGoSo/k/cKaOA2AGT7IiZHn3Sbco8+3CDlAM/koEploUn4X4WLpwtuhCne/+
llS1sdBr+p1eHWjHTXcJmPuoskupyg24SQrwgQCWAW5p9IZD3pFnHmJthFWm
W9yHv0PiQD1D2kA+wSPaKhhOQA9/7SA5Lh/Aup7nXbic2y+sUsS+XfFNqUDc
cKgu8z4ZcK8/u/ovLCnpvfySKofkHT/GYIMYFnXeY/T7q7YFWDUQvFZ+ySsZ
8/QlQRH0TwoL56c5rDCYGWAm0NFxEkg2ewI6ily0btVkmxVp/wF66EWzaNue
kgjGru8VDXQkUPpRoiRuiAmwRc8+OLvku3h7y0ACYcP3p/IoTdKbqzu/dQbS
9vqFvC4pciC5h40PzG/3ZiV1L4u5VfMif2Oak/0orPDUQ/MS7FDJIgjKbetG
KVJj06m36bbZidyEppBxaUBoIp8+YkGlwBiU8zyMfW2sl/XuNf7FPw7KOW+9
lPaMX6zN8OPT4+f84NQYrdoIG1xujYmWZtAKkol+JFXTbKZ3BbWHxbAsitx9
AY1geKVD5GEKDkJc1Z7ej9oTm+wm/883s9JpAeXyMpUr44w0b01iEXyEdoaI
VyH60FOY899M5FSgFWA5QG7+31JvO9c6ljT2kz5xDiWYpyiSBRS08yM5IbID
n+GZfDYhPyqkQ8X4fsXsfncjouhZJWcNajYLaAjyZzlFj5uvUd0qfBA5p/Iz
YvYksIiB/KOAHutjX5O2aEevXeKZluDt8X6EeM0TyYwwLxAy/B4wdnyrQrMf
3nkBOpiYdKRHxv77GazLWU3igKMzX4p6F13e7ksR0R6mTuo9z/YpREY3cGhE
ckB3ld2PL2nh2GWW8kRyZIqMH4oJ+U3spr7nc6ILss2TaydszkHgDKbEN5Qg
mstF4KsmIitmb32rooRRQCLsMqI1H+4UPrsMGbcu5K4WXsOAZrFxnl8b+cwh
uxg6U4wsSaJJ6Nv+EPL67UDdycqDlSCNPLlotv3Y52LyHDW1Re2cgmqKJEpN
PnW4bdmi0RVrY77Q7xEcEAa9psojcT63y5ahuNhMemPSY4tP9Xn9KdIXc0N9
VEdesv4dx6LtLyfoNw5vxQIhp3cIn1DGWaYOb/y0Tu59U/YI1HtD87DK2aRs
WKgsG8FpFBnrJ+G+pleItX574S5TYvij2C7YqB59AYQ0ZCW0XboHshtbfERF
NAhF1sciMQIhNZcw4ef4+9FfhqUNhFsR+aLY0OgvgPePnuCXNGlZcxwqd/Ln
Vt/W2QL9ayrT/WICo4XizhRwLnySuZpdBZCJKdhX4sw+38VnB0aKw4YfqC1S
9p/9nBtasXZHNhTq1aBpVm2Tr6ZqtdAv5kkdsNQJiUvhr4V2lRoYnVrDMVEI
cJqZfxjkw89E2SJl+L/GwAw037+V/7PWLHTM91vpfUql1FgHIFSXsjIH+fwt
LPgMNqUMlAHCaKY9d/mVhapwB6+dSiUs4V7V/cg0urP3k5VebN1ji/2K3Z8H
291kPHhcduxv67GFfY/x6R7j4tE7oE/K3p99N5rjWMr+UR/8zhyPfhoP/3N/
Tg0x5GLbNrfA4yr7gd5wh0lVmnCLDhSQ/4GT/5QW8JNWm3Y5a03SMHkydEzM
K+lHK5AkbO8XdMMQXacfeVv6LbjAGXsBkprzP7f/9tyRrmUsMsbvX2nQExxQ
EIh95fWENvORuu00zAHcFomrCyuNECob25nwomBgQkSCVnLc11l1d1HvLB/N
VhV/iZobV08vbDqaluixyvAmsfgq6xyiFEIJfoF+4CTQRyfnfLRv/LG6TI20
CSiJpqrikJQjqshThnyI3Y4JnWdX1IAM/r10q0trdh3xnwfMNmA2I/SzM2cq
EVv2VLOOPMhNT0ao0o3DFmozhK5jxtegI6XeIcnGyfdpWFzr6FIgpBi1PlRT
MfF8WoRGXTwZ5iJOGCDAcLh9Y1Xz+oEvc4MTBk/TTwXE7KjIAzQxmomhIUBO
mEEFTqlzGeDxfC4ks45MfZ1dgt3NDkZFnqUFpLKwAN6ynA/0C83nH0bWLt5H
hgJBxJWE3jsMfwyC5lb2k40suL50xq+4ql6Ag4j9aJ0mR4flh/lmZenfOO05
qeKYhTbvNkxbbeDPpaE+TK79lhrDRARD1YXQ9f5vhElvtsUC7gzxh60/wdnf
EJrP/fRRkIGU+GAuCMm/0K52jLnaim86yKFyBMfxDaXYlOyYSROvevk/pMbm
pi2KrtR3c3q3zvoxwjZBaawxjb650o02S8yvgTpiogzUD2tNnV6Y8Mu2Kmta
UPuRDNV2m4M8bfUFtdIQyomHpcV7Gu5ybtJE8spx0nEq/TAgXtI/YzuQBefK
f6wSlpJlXnxl0DzicB/8775il8PelSJvJsmP8ylR/55mkW8nyMAxsUdWL/oW
SX4MVs3LlmBeEi8Tpss1CN6iejETapaSm310Xigxr7ZnxhjKY9cKYAnPdY+4
6pnFRixUn0dqWARLQyijGEuXxHVADDJuK7nqp34rdBJGPhhVg02hkRshGkNF
vr9lzFIoReswZKPVPuOr7tc0cEUgaUxvlNGrmmLZQE6fRS8XU6xDcjfesoFS
dkyvbhlsWXRfkZ5aeuzGfK/m8W4ekw2akdqlhUeoRTpGRUHNyRX+8JFwxEqN
ZPjIq0oRvRu2nsZIt+qAyOaSjxeYkBymSaM6skQfAG9IKoYPyuFsYxPf+MsP
AeTjpur2W6V9fh6Q3J3KxgWo69eVgv2sHDT80aIZIe6Db4S5oIEAmRZys1sW
cH3mcXxyVKAcomBzUs47QvSiIut6GdoJvthSP0xq5E2x0xV6IYnb0QOi/EWD
ZwhZj6F+F7S8HwYJsmKIm6XIsOAgn95xVfNw83FR7Spk2x2K57iABm/ZgzJ8
Ox1+C4HyBK5NMPvbbhKxwuQgvcMArXojf2+qFSk2qZhUtdmshfE39i/n0P6S
55Zs4B1laTEnXGsZKDYOsy/9NqHw3Dbh9X0rsdOZOOLjbVwi66Il1N4H6hCJ
hbjs5mpnjklcd3yZ4qym6GyDLE0XgA4hRQrWNaQ2mgdlhKf+0kSMGkOMfCvZ
GRXxkzt8ZtDy4IG5NbxOOqnPx9ODOH+Xq7qHGPvPzwoAD4CbCBzeDh52Qna0
UJ+0db/jxB80O50PUR1fNeiTM8i6XrbWkfnPkfk+TGAqr9a0lxVjh2PLLhjK
SbhaurQ3o5qwI6kEXMzcIi0JrWpvCaUgOBcs086PBPLeSHvjbWw8GtD7XeO7
pT/JTDhRFjbzvsv8DSK6SlhsBlSsyZZI23dLwtRGo0EqYbarKrMS/ultLTbC
6wmVlLCH81bYkqlpLyVuNrDdkLU8BjfqR0qAbHHcMBsZXZXmfsGx/cIIBhjy
izUdvE87BCd36W2/eprPm+u0V6dNOFDBqvnMvPM9MY6hdi/tXhWsT2BghtFx
lNRvzzz2InUrPyxwx2179+KT4v+gjQ4Dq+HPkckExYQXJUpnRJaLD02YmsvN
YkYHtDL4d3xQ+0UbaWRexcIe67iZs2CjusvyTTicOYgDaJd9+M7QMLTL6leO
zHKP2g2Rt9MQ2v9KyI5s+IzgPp0JYkeU7i6kI2DCxERyOtACTq9L1D0VYn0F
U9TIY8wHHtXMM1+H6l2eAe0nahda8VFWHRiPCZtup6PArziFgB43v0OXWnrT
l80y+luJbf2U3SqQcMcn+9zo8KMWHor6EBjTiy4c3xIFXOaCQwj9l0CHYQl1
lzEJY5HIn7Se9VoTSHlYiRor4cSBRl4bkyUkTEc1jfVTWmciu3MpgvC3+7G2
SE2dorndwY76n8pLcPw+XZJH7ukE3dh4UcuhJWO49Tc8oDmhCQH1/uB+v6v2
gdXJlXTAynad7WoCQdX2PI7Vw/p61YGlrQWZu8qfrZks/HdM8coym7b0EMip
tue2BXYdAU2L0Qy7wPAPw0L6qIyjGUOaF1cupUKNAXXpl5CPo7vcJ1wZBF07
Cd0+3cd6c8Wk1UMCepIx3o1utVavf0OMueTjUM5mRv0EpJDAI7vVheRndpaB
/Z5nKmLPn6TwINvRChYrBKtkkdPsLK8ooTfx71vJ6CI7ODDQQ5JjxYQxxlM1
AydGdXPac4so2XTpFPpJBN4oMARBdVF+jP2ptZGsExfNtuLA8FWpafnTZZSs
Rc7Vjwe+9ICgngyEIZsXcXdsvKr7WFz/uJldD/oBxgoUwvrs/Yupf5DAvlib
3jGup4+TLaG1tSSWPWbw7mfimg1egK8lTRO+1XtBQmmBigOGIZ+rGTpxFenQ
5/lCg5rGL7dJmAxcLLG5iYgsnd1au53Sbfh9x5L9c4UTQWDMI5sRx9WFHdz9
9HDMcH8ZrYBmg26TVjTd0mkeolWd13FmP8Fxi5sEetOb3cNNaa+d3FBxJ/IL
8yuke2SXn/hoBlaOmE053Gio2zP9Q335JOzWTwFkjqEeC/scKDI9uKfIooyI
w0l5XAHNP1qcjZkFv9LnNCprl3IYLPfLHopzrDmaZHfzJoby8FJ9z431jGiY
LGKABDwTUR6c4pAvoLwTKoM4NgafA46VRG/tN8YfUpKBWdEpx0/kzVQFilvu
+Ng27n2URv+dTLfIYTqp5QFZ5E2Tjy4YDe11jDi6is6FTcEywh2NLSNMj/v0
gNR0KpU5+HNhU3d7ak4Kj9cGOgkOkeAPwVLuRTRmcpBmvLb0hVU8G201s+X1
qHBU/jgmXfJlvJLa6++aCuTdDlXwKFxIMS9/15P2q4+qHe3pdlXGNw+QezX+
Yr0Sl6pFNGum/KgwfEq5noG6nVJlFR025RBfJnB0Qt1qfRGDRxSNuWaTTVWB
wctUrW00S9C5IOoXF7wq/O6441rXx6+ZjyqRPYcDkdiBKbP2dnsxrx+Yh1Da
id7kj62sCAN7yF6JkknY5dRjx6H2WtVK9L3LbpXMvyzlWDtwi4UyM+Fi3xT+
jt/1mI0lD12ece8RRzbCLv/v1HRDdSTNqRxv5CVeCyC0KkmI105OdvsbmmDh
EanTaRvWRMBfYzB21eNbmF4xhV3tfOAtKZnWV95gAha5m35CzRj8kz12bZ1i
OCq+DEd9mg2P/+wnvcR6zohP/qKlWdJ7iVxkk7Nbf4t747r9R90n9M/P4sXg
zwVWKsNJ3khV+WoOcvwvO640lJ5NnqtBDUjjAa3cPR4pgB9HEk7HNY1jdML1
JtUO49lxbLegwDDqY7oJHV4X026+kp+6i5/6r/SUTk+kGgoRHOhyhCKJaTBO
+TpDfQquloR55kzLbK4oOt7qOlhoTL9o5IqfaadpfyZ8UEM0kIXZiJX3LmjV
pZjdgGrT0sKYFhedyLiFLIggH8d0bPGRNNollPr/YgPuu9jGZxbzaPiBKhIY
c0P0z60TFZ/6p2uXOpWoHgdT3gDT5jQ3DCxJh/aoG75OR8vS/hjU4zrx6d2F
zvTEc4AjKs3ikItm7rrP0KRjY+Omcavy7/N3zojlDd9WIEwOM9cAmtCbuBaX
lpXKqpGY5BesDg5/7/4pWX/NjZtjh6rLkQkSSjjFf7MqzPsbeSbAHpv3Xruq
Ba8f7S4XlmXW7pwW3fD4KmSmlo5CXvgIM8fSPN5oiB9dDrvUYJib29CuTH7I
M8WmVgkLaW7uPvaYCKWa8RyYT4hpDxSnYur82eFe3qmRAsrbGqyqWIKLh6oP
uZI9ERKXjpQ+GbADZ4mfus7mtht0LQyggU+3XClQRR9qi360ypZT1qU8WO7K
LN9lxCSCQ7v0T9deKR0z7YIi1Oo+EHnyIC9xcoS4w5eS++ty8L8CACGrAHBH
D6gWG4TvpsyTFswExiEqKkoMXHGi/41lHofkPhJymTzDMKWQmcMKj7NUEJp+
cUpgv3Sxw9Dhjfk6NXVNSynagIeHBObZY4KW41SUuSbKgkZIHy8HtUa3kp5R
nxcNtxHjIQckmjfJMs3zj+0aE/G9tioJeUSeWC59UlzdQhvTog1gdVadsF11
P7LQ/lhiVQN+9ccdv/UHW7UgoQMz1b51WEqkJTK5KVOgz3Rqf1oOwlU3On7F
/nEeYJC4S/JrkGW2BBeHj+ZyfO7nkAKrCNodIdsYIKU/GDCO5RW1INS+GW/x
zLPTbhVmb0cR93OUKAngnZSX6PZSrLgeP8SwY8ASWJj3lz/PFixxMYP0i7vw
gp2NGIxzr7I/eisFEj4NGUutQMmFA0vDdUg+tcz/G7oVbgXO5gPuOBK4Wt09
h7IWoJpdws3G0rwsRhDwlEEdE8xi7i/P85hg5d2pmxHl9HVcC35IC3zMFnzP
s+XXvCBqPogKH7gTTLlm6tWXfTn+ZvGtLOzAZ5K+nxAOhGJelDwBh6aud2Ks
PjC7+DOeElT9o19UCTlHnaZsQhPUE7OSpo6h03zfIr1yo0lELBXbgnJn/Hyo
mcoPzHK8KKa53S37gsdxGBm92f7BBqDCP9eCMInrnefy2h+qKPI8rtScHDE4
drvn3HmfoUpieurxWlBBnivAmanjpkYKVDrKWCOUq0cCaqQX9zGFFrcFX8eM
ufO7aafRngCqMeBDN6PcvBS1YWP7umtSKpEPqss1O5//vMW/ylF//UCHm2xb
SAbc2CkysG2KPxAoKRkBgi3aHbBROfhK6+N/0TwJlSCTcql44+YA05swArcd
cbfFcNV/LTa3GQxB+sVOraOnewvFdXDyo2sO/AC0pzzgxOoo32tgVHzWqI8j
pLcEDwZ6xuIaG9jmrLr6o3Kw+dCWCqATngovFzVUDMuDfpFBQQDRWhvPvvMM
eD8jAERNgctlBUbbVFpglZmVRNXfzKv5YjvAUfqri+lfhQQir/7PYoIev6zx
W6svVr5PAjOejRFBJycjhmIGhic4deLJOCjBmOHbLNFCHuXYNpzoKJNOEKM/
Of1NglEoEsobB+/mxonu+CVCQfrKhe1TXpoUED/BGiFkEkIiFV8CaZ6Lt9yw
ZMqipqEESzVWov5Q5HIc/KbMP1l84o6uC/3bLSeSUf3U72pwxLLbs9NcToL4
EhNugp2RAtYt8JKtD+06EKu1P0lKpANBJ3EhPQfsGQTP1x1oRESkPL3pc3p0
w6JChPIY4uHgNoOr2VCVRkJowI6vKu7juBSVrfea97lzX0dtSsUu6NFtLEne
H55U1gYmhq2onS1DagHU/6OfOVgl+2pVqkhitB/5d/jZxWaV6boh/oDNAjPF
L76H55jd7QrkpxNMkEsmN3ABF8YE2iY674piw8oQC7DGr4fk/YUwnu+zWXBD
kICvLvxfEI5wmmrrHuOt2VEEmKeag1fQ0t450v+wnNpT3pPf83+iqI42S4si
pgrczXVytPj4mlN/lmZAGdD5hnleeJ+hC5LjaGw1Pbp4IfQqEGUGdHaNq55H
RjwgyyXjkiMDc8avPcY7L5DDvonr1C2J6O1hb3BSif/5P86Mxhoj1cl798kA
LB+p7Z4nyMq99t40KwbPkBWPHWHwcfrsApbITCsF295LF2wDJmxue8yH9etY
SYROacYPKLPGEnkz5WGdSkK/rne5svZsbgwS8e1bkHL2qWWzLIiKCaqkPzcO
BmglLGJuPVoEcaaPrJMgiDVZKl5ZcueHmfutJ+tkfwNXizJc31TVNfNFG2wC
iOjVjDOpAsrgcxdlyUd4sI314NRDPFSqXvWaZMIaXI2DqloDGuPYRhkxpQgs
R5bhaIEMOAmVVIMYKU2Yg5g+c9+If+wiXX2H67NoQuwnjygaz5jeu+r+kTVE
yEIdWocllfYXZaviHAe0My2WIy7YHQqFEfuoDmn8r70DlT+Kn2DFy1DMj4Q3
f+J2lIiv62ffCjJbO8jnV+hV03IwsiHznN5wlIGL2xLVj4zWcZcvtbjHct3b
M3X/4qhqjBY3x5dH/1J3921HAvbbv/0JCsuFyum9qPQRIAPzrotTMqJtpVRS
lyFk3bN2WQRlTncu3OzUudbz35h5xloFwtHqwyRyh6jqPlR4473w66pDtQts
NV8pGNJtIi0Y7NpCPPheRKu7bwW6k7LmRJrzu0Xj2+rb3aBs1RZ1ziNCZ6ru
KVDDAdJB8dFA5uJJEMjgH29pEL9j+fm/zN1gXJZ0Z8XBsLrT4dPIbi7aJGFh
5AlTIjH7iSn9gSCfWfpV/W2flp+gCVXmoDeRWazSkIoLf5KVA4DFfXMYmIuC
d8xYgKVk21X18gsngVWwwTtDHnCPLdfFFfjAR3tsg99xnO7GWjNZ3Bq6aXuL
2DF6OQNZnWAHhUhOScaRQivxybzSvDYHwX6DsKlT2giYV9IrQjU0takjsdLs
+anQQpSvq5CWBQdPiLgP9/rh3AC8Rha3np5qcnTRNDisxbZN+JtG8BZ6oGFu
IgT2t37KwhCtfHwCHdm7FsK0NbXorzDchMczRDBr/H815jB5xbn9rXBIrp1n
E4jq81m53emBA6UURcLH99KXO5tTdLl1W9c0khksj8dqiXBnTZWNe9RbI9W1
6bbeMhldmSubjZPrhT423e0IDxAxnlt87or4GN1xLmAA+U1XYqGsNwnNVHPx
C1DFTbzjxOQaDh8qY74/K8GM8EpBGPEnIHiOpmo0K/oVVVtx9Y/L1U8/+JOs
xC8stvP+M+1KnUzmpPDHE/8Ht6UxHPTnBoOap1PktatrhQ3ugmG1QmwpmSWu
9h3DhbjmlUWuErk3EchnPHlyR52IMrcQKfi3IFSKN+eWtD3ey9cNq+35PbBA
00e2uAGq0vlhCSDSRGWaSAUb1qqzUJhz47bl/TjUWsTr+5RUcQ/V1vdEmLyq
S9ihNIk7g5COaMFqG0nlsPFZ3W+ah9mc0CeKfipzBzZV8yivEwZmzoQoko+9
P4ExQWv9KB8g7e91DUC2uErjswQGVzl6rhbydaaiENBKoWKSSpAMohl0jFg1
XiNWStwK/UKpt4SZtNyocj1Je5z5qsSvl4LhqZWR/8Gn9nBdILIa6/cxyu/e
mMOWkjMEdSMeqAdy/D4/tfTWovRWUlUn9I+SZcUGglzq2UQQ2c/Ya/YsMTwR
QIGBNIuXDh1OrOd/a1ilQYaKKqbn9qAwcEw6vKFB57HjhtYeRUqg/SAo5ygT
dWh+1uT3V/ACzHFjhaLf1cxJnpXRenrl9iJGTrdsZsmKA6cDvwmql3+G0/bk
0Fkq2DHV6dYbiw+9tNlHtvSq7bhFQDVpeTp/DB0J38fLEDAFgakQr9s5yGTX
cqAKEDcsrWt6QyN98KrjxNP4bP+hOYK8DAStn9WVmudCv0QvlkiD8s+kb2kP
AmliX3H/TwyqUszkpAY8/OBCMfWUaMGt+TteZrRZheHhuGJY/EIEjyte0IKB
3P1dKxPkiliO7Zaqf5MqUnwAnX+02LCyRCRZ1nImztyV/3tdRk9i1WsRWR5h
fRTCH+ywHR/QrGGEX/PVljw7Z/B7aBuQFqa1PU0JigQxRPK0M9NEYfIJUe0z
adJeIPE03r4Zke6vhBRzCsVZq0k04BztsznWwLuEN5UwZsqixAXPgm8VdFgU
huMC/pzTutkCiZkYPple7d2N9/gJjj6bnILeyklGt+q7P8PwEYe3kchZVEGQ
2M5w05zXVsOIO5PJ32YNwXlnBD6DABXLD8A+j9isEa2NMnSVY1WbZPdUFPmU
cq2Ow5tQvtjUzlI/gCkLl/XCBdY37g9T5zPtJJtfDx/QYjuKXOJ5iSkKRjNM
osE/+25t4jES47e9JWE+ejXyjovDe93vBYgAeFo4UUT4mMmlwIFAPKSjhExk
diu24nDlDdcWC2XaMPdNq3+melS7tdBtuWGTEIxwmbopw93m+NYgk8TONyct
Tbev2xOb2sayVRL48TTz4wSuEf4c/7HYWLEU6B1O82TkzNRagtGKAgFJ00Zk
1tOGOf2AuSuznfSqbVDuBKZdSHnEqSyUtEPG2aJ93LrX7CukFOnP5QJF/rx7
DjZHU8ECiCgCXNUUsI7YFEeqmPYHoqlDlwQqsRKnH7qWxz7Xi1csykQLQ2Q3
cEUz5U7r4ROoQTJZpi6bWiMG6838Pb2HzeSp5bEiWe8dAE8gSu7xr0Vsx3qt
ikdaZrbtlbJQB0vQNR6QoSCSWqF0YUxA5XFNmyVrEYGnmOGU27gRdwndotcs
gtAdG0DKZPtwv93YDzKZ06Rve1eOCVer5LVgFCRuiJoEukfbFHAn2kCFb3Rp
v/kwxejwLVuTmFPDJAu4QVB5Q3pqYep4I4W979Uedj0WuvbH63uczF5LaA4Y
QzrrJ/wlNSzvntunofSYK0vko5GTdZllTRXG4DUoBRlCsse7JaWR3uUZh09V
IXgdk7fBioZXBoWl6dcTEL154Go9NidhX2vFurvhOfxz53Z4C8dPg6ZHqc0Z
sZXWfFygMwxMVIW1ch+pRAf7zZCZvQS/GHqiJxhqiNbb0AYKFvmnBwv6DH6S
0ioJKN4UBpM2yL4QLzh/a4lIl+znb1+4iAT1BNIuE81BUzZd6aefevZvMEGX
1lYaXp5P64JX9+Y/JDejqOoEnSDe/iIh+iOABuFI4ysHmqFzdt7VGmJLpEhJ
H0jWohD3A5uBHKQXTm0IjOMeDJZ24NZS/scVhYIN2YGma8aaVTQqOL0GV+u6
wf+Srf+AB1ismQyovt/eU0YmqO/6RNBPHfqWeK7UE6pwgFSGkYE1QVjTMYjJ
RV53GMtov0uwieL/YU4Mp98ndrdd

`pragma protect end_protected
