// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lbA1IF3xuWPHYYSqLJJbl4UjvKnNRFkiKxxn5hjXCd1pBdfqpsyJjuU2KjdU
3BAqE/ycdMYjn9HrotitpwwGnoCtGmDySYjGtQq28iRdjL8f1phH6wz3iI9S
1DCeyfvQPbwtY/whowFQkrkNO4+K+NdHtOWdJvgwBSTfnhrTmcJHaiQLd68o
dzsNRV4a29bTn/H0pPjGzkG8JeP7WzhnSMZ1KMUizy33JxsJMV5uM0Sd/Z6E
VtbR3sfTjsWpGz6+TM3NVk3Iy88opIeIxmGW1PAMmfFMJVdHMoSp5aL+2oAR
bkjnKdS0om4ObinybBL3YKb/eD4xXXgl4hO1f3aoPA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WBro/OpK9KgYguqzHdXos/OkLwPXgWUmXvQD4Oi65Pfkr9zLgErRu/Sa+RUS
23gaM1zRKW4TygcxbsQm0UfkpyrgqCWxXZgXN23L1ljPRZaegBsELqTousDL
eS9y9fsngFNyWtt7qebFwzEcKgATG/5FQ5xD2cqMTyAlP2ljkTvY9qJJYnBr
tILL9atdlVgKOygD9dWjxmdQUQxe1jddNaTzs1sDsQ38w9G/2Sd6uRwsKga8
wNmCYSE7fZnku07SdhjHgMMO7cjWsjQU7b789tre1BNaX6cqJJ4Nxx0xzHUR
Bxl9ri+u2BcgFdqChSyV3rBEt1dqQ8Aegp/giz1swQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SoJme4CDht2tL2/0k95T/XwVi6tbfSCHO/epAQc3GZFspn1ULJ4NFvLx/Rwt
gfr8OLfnPfKRJWaQXZQl72lTNMgCCr8qA2If4N00yDIOfRQWgR/W54AwAOvK
cph7XliNaO5ESbqyL/dYhlGmyMQ4o4R5ADRriWKXdmbXNCgx5zRj6VbGYeBN
oQl7p/V/xVfwkqIJxcE6HQLa2rpKcSlCtjmymSbT6md8QjF/z4nLesJ+h+fT
HJUNRl7na1i+7MviJFuPpMHd0SlYtsz1AKzRr+cP+1H8YU90LfKLu53O1AOY
R0D69/YZzrAO+I2Clmy25w7RUKf8axch+oSk/pe/OQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TZTndFagQCfHC8W/VTfNW1J+Tu4iaMevET0Deat2gn1Xzp1dnZpRCed3WRc3
gOPXSs7E6sJeWhlZf7AbGY0+RHelkkkZcl0tZAEGLQjdRQoWfiTpWPX3JiSw
wcEfKmd3TyEmbrEXm5FoE8z64YIXrxgV4zHZbIswgku5/rATKAQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eWCX+OpclZLnqL+MGcHb64DwznBHdZXjoZ7wWi4kAdcRc+5xz7iWMmz4E4kX
xRllqPtu64EpxWbc79daEAoSgpBRxm7cHhoQgeWshl+IsFlP/XQVMFsPwMT7
mGKZD/nIBTWZU7Qdlmv3/X5/bo6vdGu0mm7N/aXYK+sKGZwK9HczCiuOE0Bh
Tt0cTaaOxSW5ipHnsKa/B3Dsm7QCdQGlqot77mM2iKimXBQHLRRPKf/qu1In
u02tO5VwvhPm0QoehHFSp+/Fbz1t+u5+x976uxHW8AF+1hxHnp9sTSw/bGfr
gqcNbfgVOHuQgpGZjFdlW8XnT4BaPyRJUlXNN6Hr5ZH79aeuPq7jO81GKXtr
VBS3kTjOUKPDX72Nb2OoZD09/cD0ov1NHnjFtZZeCc9mPxawgxEFAJIRxnw3
aXThFBMyqgislALuQxad+6kHrbRW3fOaDOlapwCX/fXFmeo8We5VGDUCVS2j
MxG8bPMQWTUitJLLoFnWI476nMqxjKKf


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g5IQEPb4KZhXNxCk1Y4ffcPhrT9Ck5VzS0RZw9FuKP22O5dg+3vnglarIoKV
ytQ9ifsmXvjhGgWASLKdqz9RlUTdEsgjb18rwbiSDmnhROt2Tc+24Myx5DI8
bbhDY4Cuy1euZPgvjQUdfnWZ9LaN46AX7fiiFbBoODXljEMBako=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m+JbekS1jlw8kup1GKkTj+tPlz2r/lgo4fv4lf5xGgeArIXRSWyKcKLbgY+O
sZWQpY9AsiE0AyQxzhK3gcdivzEbUVEgsY313yxUPwSrRTRNfym2hIcV9vhr
ZjfEBwLcghz6mAgc04auCrlKQFJZ42zXQjoid9eqjnqeTIhJj8c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7440)
`pragma protect data_block
Tyfy2F2oQLjYj7omP/g8L5I6qcxs9cr6Vyml2LIP1a91lJgIuAZnpbzyKkCi
jAHy2lW72zZk/oKVZw2rmCE/fRBYEOmeIH3znEUSEE7OzvbwQtLS2Nb1KAm2
4Il/9bSrTZX87CWTP6+Zm862WGqoXFCzbeZCjjtW47Wibqc1HH+jbGPHHF2g
UY0RGF84pg+HqdIsgzwivW7hjovYc/SECIf6BwevEnF8UMTQEgyBE04SBWui
qL2OtBQJRTRR1BbLhkxsFFOYYWSCiI05vziKEJkQWNCEcrtdnZmeOZLLN7xY
XkONHS+gHv/6iw8s+/qzdUbHBQsBukgKojgbr0XR4aPgvmXT9carmV6fiqrc
XpCX732r105dcMWUxPGZoZA5mbKwOmILSXoWBK42qSz58YZKW8Dg+Gyjvgpr
2AxtGL0fJgoKEz8jxg7Hsm8x7qcHCuMXrCFplcS2rulWmd3bogHsyYC2Jxg3
Y2wWyaFrsegaYcKtTKK/EwofTsIFNZ9yMJ4xEvTOaFM0Opg6BghPB6e+UOtg
4GWu4jqDVmIBHcgVfevULzXs661pYQ7eXDckaq7BabRzx7r5Anl4R+DA/MYO
4p8DQ5RD2C7iLq4++AXejvBFuypgkKb51QLHkVRu7a1ARrEPrc3akPPv/KUC
1bQe3wkMi3udyMaDHbU4NRiip0D8O/R+lNXVa54fg9F6xpAJicQzZnb1yRr/
k2sbw+u77FbBIogb6ZeVmdJ1J+UkjdFgkyj6Q89V/xlesMjL2TpN7bWDK6yI
U3E3idS4UwTIMh3DznHIwqJe+VR5eMm8o7OoTxVXlM+TEBiTu33jt+G4Fp4n
5qb7w1I9i/nquzLiQ5x9/YEecUr/BRhEHJSTRXVtK6nBpxYeuoYzTi87CsKy
KayPWo2D141bw/LMZH1M/Xos6RV6HdxkHD8wPh/IRGbGc9iuZIFYkzegBCoR
h5vs4qHfSeiDLdiC7IaCCO//knCvQOyUkZZlihIRg69gBSN43iecJBfig4JS
/Lw1LgjtSOcR50bYNvLXShZ/pjO5pgJYdOf+c45XRSkaBSP25zqr2uIk9Fk/
TzpMBO9znHKRVVsoaRR105HXvahiI/TPC+7LkNRV/mz78aSUJAlxgq1Ou6lH
XuGjXlw6VOlaim4E+yGBlmDjE6WwqcnlOnGhdgELT4g9froaZ+pfkTyLmyXU
hND4jHz1bfInQ+JhmybcDfgqBCLWYIiMZiameq8S7n32wZms/3nZj09SWJay
H/Yh38clUijvF7uX+ZOmpWcmwTRuYSZ2xzn0CLsLHcjnu5tJcMM4sxnkvtJR
qwn7jQp3s6R4u63uydPEX9cvYozMXQ1i59wLhqIlteDCFR3fKqLHPcfu+oZ3
76b9lBsHsCJJuIoEPE6F+p3my6Qyu9ckV7kaOFH1Xrd11uQQUu4KaQ8Z9tuU
cel6bkVAG2HxhMqgHQYgSW7YWGxW2GbS7Km3mv1Lchz3/BURRxQam73TcTwc
DKkZW7G8kMkJ+kmbRaivtlrGQnxTJ/bax4RIyzHC2OoeCmQ4UKjPdaFkUdbQ
NaKvmOmH7wyrQ7/rv+bjxvj85kkrf1UG5otMKEQjke8bnurq5trn//a+k6H+
+h6onIwECX2/ADflc/kr4SEsJ7BTqOeD84KhvC5mkwmwI4RDwTZ/91Tt+HXU
+0MSjo4/je9bIougeFyt/m9d90b+FaPH1kU6mZsa8IvRk43z03/k7CGWnpcg
kYgHFs48U2e9bKNDXaN9gv0W4LyLkJoE2786Qlo71bzEiDpV3sdMNpJTS7Ht
0yZi6on5eLlMU80cHxjsvZxZ504nPQIRIHpzkSLUEQySVL/ac/TdCAmozXAP
W0KqVYMUF03+eovdliPSuiXJWjI6PgpDNvcrlyJac0m8Kj46QHDiwq4060ih
8ydvVwXq5+JiQr7n7KeAgy7BaEMhas0qoBee3tcxjtHiKFmabgrbTEbN4sOm
ZMzPNXGLW1J2va1b9UlivYWmmH9dXg542SaG5MvVVoHzaW7BtR4Sw+BB7NKg
MyWraUYNpJqs9dD+ts6C5YCYhha78FjbWIzsiaf6q4a9EmfYjz5qEl5Df6Hv
vuM0wDYc6F8ZfngbJwH/O74XllJJrO7aBJ/aONtvBBV/m2hymNr6X2Y4pd8m
Z8XkqgtWDk/2tKsQ5A9XR6MLd4lwv73KX/c0Z79HAuYgZD/OjNCOOlFfIvgg
criWF41WpKcDyLxcI+kIuDuYyjWk0BHAMxb/9/wu/2NBPS7Ma1eLTcov/Jb6
et0ZBQvlBSlI4tv/U8aC6H4EwOum7oQhBE9FsDjGPbJsvVbsRtqAkvkSf9jR
QQct/ZUfCHkf85bxb3WKOe0inZG4hGMSegWTe5kM90ADYj/xmbbPVDxwtJSN
fn0sSitc4xUFP6hr9anGy/gYogbLPq0ThZqU2cfThrmauW+z54+iXlyQB48h
s8FRDy6KCbQT27e4F/ExxbKgrpU/4NSdGkFkgSwn4ZzmwbA41qlSXqeW4PGz
Yfg1gbuEzmPZpkwZn/t/pDhtdpFAsMLWJM02rU0si+p/JxD2Y1wZz80Goy3r
ux45UkPRHt8Mk+baVC1nqbpA79uZGVxXcfV3oxKNuqOCMyB9wW2azWv4eriI
ihewCZIkHGIbz9F8fF2HibirSIdJseRZTu1jGvXxNDE8PTH/bAA7SIVXxP8Y
18azAvv/O75Rn++dZJ5XcZItpZrNmw+MAmo7bx2GpLdikxSzxy4ZyApREYaD
fuu/W2gKyzK9pUvUmwB+Oy7XbdoNmfbFxkl73/edHOwZ2kn0HM9O5BsYoVPZ
v05B+L1BRiHHAjRC+Jl+vEDXN29o+6r7YOBBdEpMTHy3AFP3hMnRWDPTLrav
25orkk9P90r8fztQ4h2qjeOYn5TAKIj6vA/kjSn5Yj07t7YLRow5zwGpSYma
LTrwKLP70/kN1ZwqVUOVH1t/ykl7bufwerm8jADU4MNi1nHaSwsIAxUQNpKX
rP8Cfdrh55uu+vNnx98APZdiSH12kFD8LrjHLT1K9nOdO2CY6I2uWVVtUS0Q
aqrxicP1c32gTQ5CUtDPN61R2c6vBJ1v5m9sodiIFgGSp3qsLXCYUVPGOa0C
YphB70by7Y9OAt04HHzIgu1Aof7faHDXMpw82IR8naYpaoYdKitFtRclFPQp
df6qU/oBJsmDdB2gibs/CUjjFmcCVBBd7Cns0ffEMocHZtfMpgP9370ZW/KH
smSltCflstaUDltJ9fiZIEy2SEJ0gXMxI49zWqs3Hf3mlHXcWVKrLfRK+Xh+
nDBgb12rxnCWHZXn5h3e5BVBDwLjQ0tyOYtusJ2DFErrgiR92Ejg/a+SE0p1
b+ZpTuKGCCxwtiYFutcNqa3Kx7UvWGQ4zTSiEL8JjP5U3gn3BERWxeWMU8Py
lklGVOuFNSWx3H3/kgiP9IYudoi33cGqajqb09Z0HZ4s5gA0CuQG2DICnZsC
/8QmCy6Ppb4xFeCWo0NSrfc3C40ga9wNlvb2uoMI4jrhzlwI3YiZch/uGPZq
yP6rhqi2js72JAp8LNajep7Yrc94vFxwVGv1//p1IRcVd/2SUOh3CRcomeZn
l4rLrGli2Jffh4mo6zGCnnaon6spQQnz+Gu1t71GfB3IdywVmY6UYdmBE8FS
gmJFePB2mGQdPnQpaay2hnR+7e8bNdCVWOPReOnkdQMH5ap/gGq0wkdQy2zi
HQzjUGJQrm+5r4UDDqQ8bz9kMwRoPLY0carr4M22a6wbu3ZRCpe1uaj6kHQZ
ry4o+we5KnXvLCjNCIx9r0jZKutMA4HdtvAlsIvRVE/jUQv00CId5Mpnr12A
A1KtWPm5YxTkEkEPAfXvH7wMl9K83QGpUXWCoQNKxoY4CuMTB66KWtZd0lEX
iNyWqOQRwdraveuP4Pg2fzVHqL+V+qNBt+UrFdAq+XtdLIzCwXFTY9oZ0i1i
auJ0NUd25jwRF1IuuILutBHE/DLlK7tBbWbmOUIRgkWPIU1BTYQfWHIYVHAm
cqnMXf1dWSAWtZl0wZpWoZq5J/M1ajobuzbe7+9XcKywdpuBVTaGaM6LVCTx
gA/AxKdVu4apQbCxpPTa5wu1/VHrvD5lMHBV/0xnWeTUWdjUlOXGcZ6dItLJ
2W8rW2iu4vHzZab6hoNJfqoWrfMsT3bWHnne0coTFDZ5U5LZsQZjmDMUVF8A
OBrLzmdhWttVh0B1sQCLIjVvDDUB6NhqozxF1wK8uwX9WkWptRDww20fIZ/j
pi1/kDfJlHlxwWnGbknalzw1FNkn32WML2oDN7ouomOadB9LPwDacUmApKir
lpySVf7+vyA10p3BA573s1LVub+X0k7GqaChhQzTd+btzN5l/2hOHyfV92PQ
GVF/nwWWtKkLCIkbr+cSSapBVDiGAVUhrZF5yUPQOBwNXfulcyTsDnNHkAzQ
k8j97uaWld1fdr1cOfPWfKbVtyqZIEvb3I2SxRWKG70Lzeqtdfpvrz4L/k5y
K29hoz8oyzKaTk9jnNAoDJuXWK01n0v3NTl0l/JvRf1hKm/dsY6aBZGPXUvI
IcYzidfs/QNSIDDmQx31svjapy6G6eBDzCY4rb0bEEfNaR2wFaTR+fkQqec8
CNB3mStWGE/ovU2ZMoaElhegSmLZkFnQeHfLCBt7KpbbFTpX1Ihyellnavcj
Xfq/52pN5/ATcFteyOpY7Zb1+1upJEflHYR+9XKH16wNs3Hm4PA2afy/lA4x
lsGscKCUT1qOMmUjvUjwb2wqw0RTI5V1+GvTujgLtA5x7qRMAUY5j0oRDGLc
oCF8OXcMmLO2ihc3sjGDA6lpoDfCvDN5QjcquXErxkgDign5m8t5s+XsoCI+
ewxiTAM5s8Ro6gXHVXEB4MOdZlwjONxas1mMVSF2/e9gjJ/es2Iyjhbh81kI
W3E2ou9/DOPswdAEkR/jP0MF2DA2S7pKR3mwpdFiNRvSYfPGeAZDYjFv0YC5
92UL42XT6OVexWIOsGiCwuEhzK/G3hQBdgqF/LVrhoonphmirHFJiZ/7tLz2
vP6Ub9lRhhrG/To3Jwy4tE9CzSHmeEipG2akigpLfX+pFdXL29onOiJazjvB
vo6RBg7ASI3rYKpMozmsHD3LelBfvALFxgFVy/G4LDv3tk/F8d2bw8H7Gab7
IVfLy8YCfmhYaPpw3X2RBIDBjstzYwaqxLNFi050CvXnsiQPwZqRm+IKI6Jv
E0SClNJ6tf1noR07hvZpVtByzERg/sjiKt1PoA4fM/6j6qz+HgezD1eiJzRb
Xk3OlJ86X+LLeC/gerp7Czyu1uyMJZRbw6dOAXDWLZx6OCS1BhdnC0G0XqaM
DIBm19aBlsPaNcT8XYhyEoPvpWYrIsAahcjng/9nERlMvUJGWLJjKVtvemBs
cT4wkRPcsGfX42qKxRtM50JcVusRrFwnX9ds0tusNjOe2wezeVwrzoj7hAlI
RfiachiMAJ2dqgKg5viq1YfovOUQUTQe7La6TxInBlnZMGLfIQd1Bvj/tnW6
8/o3n/GORn4XtCFXgUcaNlxCBQLHm/y+y491VwJWQvzXpQWkn/BxTCpx+b8C
d7FeJ0iyeuew9ThamwYOlTrjAoE60bCGBKrTCzo5k+ctWRC9dYN4v2sXZu3n
pRHZ7x8K7Nylm4IrP78BLbK/cAj1hILbErDFOf8wPH/j1NtoYsQoU1Tjtx5U
tRz2GwWF25Feb/oTSaNJl5XXL84CXyJf6RHjw0fxGDArHaLOs6DQ2bMx8k7x
QrkKYmvPNFqho/LgZCeIUZi+MbonhNA7f8Ii3ZoVc3UknzlYPrLMvzqJ1Vw5
XqANZrOUoyIP6+OpE/zuQBGQr4BnDfjx94iZfrG59P/ooF7B0FA+X0IbB27j
RGuBMBCk2Lx77ksbpUdogCcrC0eA0o7S5juFPKJoMHxA4JP27ZZKxeuJb7pl
FTg3GFnxtXgpGa1D5QOdaoulHRUbRO/mjvNzE0tgdBQnBl0dEfv4yxwVL1GK
5AOoCU4o/BdrK3/6TDOkWCJbYJ4lnwo6f95I4s2YEFoTQocG3kQA+ksLKPer
2wgVyHzQPuyhcFcqxpflpPZut2Id/EXGeYhOoXy4KJxwCcC6j452I8vIqHOr
WoyTgNelODhAci++eqU2IR1vaAcR00liRn1gknOF4IXCE4ncG4je/Getf5Rt
fGk+b9yUbNCgSJMRgbbNZciG8wMfSbjw1RrQEGEZv3KPQpMYUYib6zYHXoi8
79TT7gBIfLKr31EVIn775BlxiW8O+44361Z5LbT9dBJnEYHe7oloduBHNRyk
gKhsTCWOtoP7WDNETuIN1NgNe5pMuIOL1XR6uCukWq/6uDQn6HHACns732Kq
EIdJ9O+Ky9GPVExwZjoIfbL7GuMsrfUDgs3+aCPpuNQme6jWx66BseE0/uZv
FGFjASD7jyHNTqPZU4SOh9lA/lyGK5Hp9tdKCn1fo9flXAtS2GGZgvZAweOG
H/N0WdnU4916izisQavY3Zg7Hu8sGHIi6M1JTNbwced3VD1q2ZhMlnpX8hP2
KOmGWLP391X4Q379yKQ3TZAItW/oRd1HimpUEVAdCH1AzDmpd6ftNH7Zvzkc
YAetNYStSuP6pwU8c1JP8PVICKJx13CLg8iT+6bOfaZmsQI0kt7TAwnHgVfe
hwIG8ZubFyU062rUkLzNp1wFKR6LhvvjEG/QbUlGcI03sEn8rw/6LYrdrNe1
jwC8Pbgi64S72b97WJiYB8HjUrQ/Np4YBZAcepnWZKPzZEhTlPdInvQ/ugxv
ANuJuwt8cHZikoi1IjanEbkXWQF+UIIhHD18j3Sp/yHLkuII4ShhqO7guq7V
BKyYy+gnm7D9ZdvVRObLx/UvF0XRMy9VzbTJCju6MYNikWv6ntEAYUBuYzKj
BZ91ZjVlCMf9psgfIpGdFVYpysB94/K1L+2dL/+q19CCES//B5M9WY6mNpTh
K/dCH1ls6AnL6e+5OuidkgVqWEVrjiS1k0224EXcih1ZrW7SrC+AuaQXv9O5
BhlMETZetnLAGDaSJn4rh7lvcoOAOUCZbuYVufd4K740Thl6yBlvm7C9Bk+O
l1gQQayAxAWK2xfyGJf4dUIgd4aHip3ICdBI85yRX8kVv6+SECleQKNKzUgw
McyOtGFfdGtZQR31uQN4cuDEOBt4ILvIywF4JisOznqRbEas3xXiZbk9caew
BhX5M/ay39yiVD2N+6N1J/Wk3YzSJF2SEXUCsRHyAFTW2kyz0pxcU1qtsVVm
6pPz0R29oEg7I3t4wE+YbOQqf/Gb6OrkxXXHqLMuV/K6cY5eUUrMQKhoR/lC
S4cf4Qgt91CV+zgJZxp0S8Bt3+1ie9m3bFAsmf2YG8zXtAMSOCoMTR5l00AI
Md2Q/KN/yCmD0+QXRMEB367tFVDK7JlJN13qR9ZT3CbLFyO52RJaMuA+CtLh
8fkxKjfBkQTbonR6cdmEpQDz2J7pGRaFDYkKAnu1si0iil5bfAMTF8rrKrNh
6TS4NPQxv9ttZ1FnILfkMsbJtdBdMr8e4QtGb+lutbxUCsWF0nkppOw+qfHD
sNjp+BfLGOzM33tPg8CaowduwmmuNTKg5jYaALpzS2jQN+ErOPZbUghPLgrV
tdX8xqRmzz7hNYf9fo2K701xNi8jtSTrmkQDQNPpUUCyszEU114rsKuPoE/d
DuaRt8OORtWK5pivBPxxm+1Nnzw9UWUqQk2i5+5r87Z6dZc6IQ6JeLXQXwQy
wddvicWOPI2StmLhQ7OZYJFrdNB78IOiAF1A1fgBdS4ZEKkGvdWNL19bDR/7
NE4CGXvKp7rxdKcku1MKohvpGCCNiCB2VAofkBvCpi7SnBmZxf/U7SKfY8iB
VBsPNn/lFvSYVECO+2kEjf2GoRvFxXePyhSDjtpVIqhge1bAWETROUSi2U/C
N6Dn2PyyytimyzK3q2JmzrIbAF9W5aoTeXUwWu3li/e+TBgclwBn6VrJG7Te
jUV6zIXJbW8Kt9oKA4Ll1vTbeiiJVTIzf1HsjNdOmd9JABCe/K6RX7cwsR56
WMHDQo7nvFf4uQ5ezoEfnZAgeXWSlLD9Tk8vaFcSK/v5FijQAiu3duFQInrm
lVvUgMasJXyZB+4XY8YTExn8jiNXxsLtXgbyO1yKrTd84XtuJCeW2/asnYar
KDoUCe4wSfkW09qfIQJQ8gzTCaCc/BQHD7VVpnbHfdCVVBFCKNBs7zKiJB+H
6SHZWFyyVTLUW4uKhQTEuvOaN44EuP/Jey3V15Zvch/fA7OfezY3bsUErsWD
H8t8C9X4cNkdnxVHstZ1SG6U5qINQ/OdszsCFhw1l6Eynte27HSx7hPHMDBH
t5T1pF61Us42kW/C1+O8kk/TsVxKAcYYMjEFtV+XZtuZ1i7djVZaBECI/xJP
o5huRGEu8PAA445/RO4Wc/4aluIkfj5AgvcErvlUkdSevxXS4G9wA6Ga5ffI
oXfZjgFMA4wUdXbc3OL0xJkOtzxnzzE3TqNxDxkHLUU7BuIuzWkruxHwi9a7
cx4A3pMDML5MhKBUtAbZrpOehFFpe3x8ViLwlkQH26W665obdlQ56eV0P88F
ooxl420zby+xJ+gLzDt+heG7nBqmcQMZGedXB3MyaeR2yxpJiFJx6qGFKs0K
iJGFMgD4eK8B2BzBLXvdW8cOhUPQTJQyXT6R80EKy5R9Y4QhhjTEeaX0tu8x
4pjxHj7kKTBZ0+ErpAXmo9ZLzr10ncpYpCCSRofFWwc75O9LaQba6r/Qt0a3
E2hBW1MLi8jfY0E5ESxnz0eE5vGS8NARSIR4QeNttWIR79JV+74725lE+H+R
7gbwRz33cJhwx4uBPXQP6wqbaYhlRIyOb9GPohLzQX3t58nmwsv9g0Gjgodj
g4SXhNmhmppUNkmurXaw3vKcCW9ZT2n89WzUXMSauAGmkdN7WR+q1Z5aPAzO
RTkDB8JvZD8prEuWoI0FZh3YBzH6REDXwlAkjlji9WLnIXw23JBfRQjb15mT
O6dPq/roK8kanZEhQH48QxpLUVCbc3Ub2eakIDTnbc0k2RuMOJFEyXAbdITW
xyNZgV6i1uNlKpt1rzCPo13Kv4Oz6puGjK2ySgSY9EnP1z2SsDgDLIK8T2VF
MVDZDxbEszj/JKCcl12/sg01ZneYqJSLJXdhJJvojymwXCam8L+6KGs9yJRA
RCi24vZg+gWL05Tal8hD3+7dcTqFcb89MW58uRWseZbfybcYmeiRvSFH7DN/
jcJ4CRRMWzzPAi8Kpna0vKldd5nocdGzzz1va1QX8ELoa5iIf363l1ej7dCc
74LOBj5T2AR8p3DPbLUIIzHnCp2jZiHV6miXyv/BMRpmKlKTiWyx8WPk+ogU
4SaL1onVStVfC1gxjSiJ7Iyg6h0b+XIi/Hh0B/cWmEQSxDRNW3PyfLVE2ICb
l7rXMKZzwySGItjb8fd4tUC44vY4K10qhu2pCLpz68Ii93Wg8bnjQUIRH3ZT
5ggEbS7hXWdyqQi167vD14+M8rZZSEjzDS1QS+vloJ60MIDqSRThnfaaE2oQ
m//lBH4W1NXXa666vGdu0WCTjboormJnXIzl8WHFl7J1wgYP5xhnVaBrdskq
d96IioaJbFYt2qoyeDKfrBCJGsza2h11hZ6d6T3AwUKulIcZf1dLI1lSXwNy
h3/UJjtILfLoeK5+PkEM+MaIRZbPTWC5HForbRf3MwVyFOYpH10p/73biJnC
wR4uZiJdpCi8L5e0uWEihAhmxj3hKATDBbNxfgVy+qkP+9LkDklgJLb5gVJ5
zAvYH7Mf2NpRNQk5owe9ASDWru1l0qV1IlcBrDUzru33C3hWqy9GMR8KcrS6
57j/Zmbv+3nzQJM5jwUFcLbt8zkw7DbBGJ9mJr339cHVdSJQKQCt3a28RB6M
0RDkBSjs/4FdjG1I02G6

`pragma protect end_protected
