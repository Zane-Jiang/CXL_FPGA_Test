`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
L8pFAK3eQ+XZlqvSUYoA+7d17SONfOAbPUsT072fCHhTFnSGQujl94Nw4UbxrOiT
5WlATFJ9nVYT4pEVDacXytCmHK4430+LUl2qmWZpagOvD61bObaPhEbs9CYtCSsg
WiC9x0cNgh5Xo4u69i4RaxzxRzB8g1RBuE4i73tM/hg=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6976), data_block
pHoMp8JrNwngNq/TDtADVctVdrAO44GjnHT8PgfWWOzzrNWce6K9WPUbDYSCi56O
D0RIJ5vLACX1M5Qn4CAx90rd5FhrMrfPH7C0Xok3AmePffXvIVVNJlwUpQ/zj8MK
HAO0nK5FYRR8UWfAyzWlBfO2WgnR0g+kOU4IxMMGysVkW6L9/vqlY9wuJC1kIqjy
7PM7ynBplkj9+YQioTQx6BMJrWNYRppK8PdMLcQUQK59uaMsOXyigczG99xHU6eb
5lDfHNC4XzICmZjVZAqMlt30yyWLX5VjFw+rw6OaWs5Zvc6PTxLaz6yl9wuYiOYo
YUvQA9MYAy/frkQg4Yt2FPauuiSFQMoidCqA1/3Fx1b16wTR8J2I3RLGPQCoLq0o
E59V8zoi0uekTF501OMqGL3d0fx6m9mrFGJCY/Kzk3Fk/jeK/9dGKPYpXDmrZG4J
cLpevYs4gJcJNA29JfZlX+XAsECpD+cBImfltL46McRW7o230jAp9xwWdBW1OSCc
JzdFyNcJbMbGhFICVbduTXAPHzY34M7g5QO+kYPI1erimMCdb9ucQy/3mYbAxIrv
XlFfQ014x3BnDXiuDWD0Cc7Nb6WVd5b/zV8K7zqF6lLTZRuUwk6gcmhhdMaQwUb4
pnqmc6N56C7xa3NTcwmlL5JJ7u06eqYd4Rxd2Q/eEYYKQBKvxonqZXXdxX4vGZEX
oy4ahnFZeB3jIc9nXsJHY4wdZoiWg5I4o7+7Qtu9Md+5WiPpYg7o4uwmP6p/3rzL
So4LHmWozIbT4giqFHuuttQUDh4rrNH4+b/9k0YP7DZffcq9tvVsNMn3ye8hWD47
BurdfsYFduCp/p6nOZBD/wh1FYpcbtFnwRNf99ndC+I2EZ5lAnjooFHN7EL6gEdg
vmTbCiYFII5N2NFJoT2ojZUZXOraK+DSnmHrO78TWbH0IG/U2HcTSZqbMlRnekGw
G+aV9W1bzOPFqKIWiyMwN7+9srFhTOP9G+G2NpFk8rkPEA8cbiw+mmKxDBFkztwi
6kCJ4kovmNeoqZB3zkco3y6lXnZ+YlyBmhbWG1Y5bauEe8caYY8xGDZIrPVMdFCS
S+7Tb1C6AmFWWqNXfIyoBRMaDhs+35k1Koo+7p8z+qNw/sAEYQWPZFtkm8Bjk/fM
ntrbGfafMwNb0SJkz7MQsyJKW93h500BAxWdrXoeUiqoGZZlAN2cd305uM1jOkvX
I+v0245yevahW/Nwg8yMq8HS277EPFsQMWqeYRH0QJeD+kRsAjj/hR4AMJyqKT2a
wbZ6iE/qJgWXCIFISWUrWnDu+qc2OrTDonkyX8UZUlr0IPbrDbsPwtkQ55dAx9dV
H3uKrS9WSFru+/aqUQYaVAk/z+GiQt9pC3/geOeUg9xxroo0OIhAkpHzH6FbmfR8
+x3rMeWgmE1qpuNMLI8f5/Y6Am9FF/W8B4N3HsxOjWwVdaIUb37oxS9henA+0Nt8
1vVq9fGfLZ0GAGc7yvYGNEAyJ4vu4fAcc0YnPFL6rDnGumwSOj0YepTXtbfI8gci
VJ31AisIdhXwZWwIwBOCEr2RNrsrBEcqgOuWZ9Q3bsQT38CWMHNTjTNY8lislU/C
5s9+dU6jFyhTssKZyykihQzEcS+zT+wgXPEHMKPegpeA4ObzrxA75DWuo+FwqNis
E7ZhtppURr/Er6uzLDwNcdwJhSk26RXdAdi+sfJ7go3Icxsl5EMYRE/GbYLkqvnI
yVyCi4VMy+5YyN8/EN3tr5W/aNGgb2ZczjdAlMZlfZujdXDbemfDcEcYGUqet5ia
U8MezNwDN/skYEdfiSjpymWJ+H03w49S6HgTJLo06bKUXCKWjPkFBpkxXvAYi/Kx
7xbcL2W5EJQrHTNibpWAFuzh/qR5v7a15+ePapLrkjzhf3wkjaiQuf82R6Rcq1KF
m+JE31qoC01gJNx4cbUj/KgctUIjBe7MEjg32Xg7FhynJqTdfSeCTZWLDy428ASP
09JmUoiXdpytoCSrzAGP9O9qUNWeiCGhFbGVNhsQ5ypTlxEblrIro6hxHkN/G2i+
24E80fNOWxtDnshXZy3kn1AG7Tg/4L6a8Hc3NIkGc5g9Z0apjDU5KM6nq2txC2qo
hJ6kLu6KEph+g9FkKQWrvATRahansJ1Zss/0/2T+3/OdWRBIjccxlLm9GjM4OYBO
Vz7mRTElzrryfXhmL3Rquk3JqhCd0TpbP51QmfPvmEDM54ayG6rdBpnrfNWy8/D/
c5N7cloWwgZ0RLPB41fBoSzK2P3jcyiTSmEkaeqaeD0Qz+VkBY5RrKBkhloHac+x
YrYJ2FUss8qHS/reYJQyweLWtw5p3DVYyPZmwImnmLKSccuc7J5O5L3D1Egcw/Ot
a/DgE/FnaPgA8MS20Cl5bQjKsIMDOXswkIy5SfnEjI7LtdtS8YR3ObEa4EPDiCMl
8FYefvJDggzSG2Qn1eZEHU/2zlmV0Dmk4W6F1kLzNfoMnjVCooB3WtIHgG3Joxyt
jIQ4dEYYW5XGQZJrl1iviD/dBYFKr5Fzz58y32WQGPXb6zCfOMCgi8L5Q6FnFO8d
kQ08czm4hbqT5REcFLEIE2k/du5PDeR0ZZlWaAcAnRKKtYpun86UiEWVCDmq5gmS
JUxK57tL6RFNKce8ujQd5+pXjJVjr9YGlKc6TODsxzOT0cS6bzVNq8VQb+/pjBc7
IEVNbDwlEJY1FuwjH1gS5NqlT1U3YjMe78dpASVBXayOlY90vEJru2UJXBUUaQJq
ZjDcHXvaVDA/eELSs+Gic24xEWRsKA3lfUatAdc8MtksT2m9cCMkXt/LBS/1uvAr
3tKOZN1+fx4fFGxALiemFcsOJ9PKYOSACK6JUwTw98J3g9BaYvX+8YCxc/sjOr6t
Ptu4sz76JmImvBbFrZAoPAA/jQRqrWXWtDlWO4BdzTe3MLJsGMKTNGfaAAZSfu0U
luoUEDwZSVGdbQZBrWpbvNsyOwZhafpOrnLxJA3rniFFnu8YYWpYs2mIdgJIlRPw
Vv3wB2qYNfiAAL4XjwbrDnHBkdtHBeCZFoXOTIpgB3SAq+b8hBokXcY8ooektsh/
xtMj1RojlEsw7fhyYrHPT0u6JOuPy8TtY8eKbnvkMSuCbKJQmPfUKL2tzCNxC/VY
taVN7oFfCokQ+UubCTb52mVSDLrBCxDL+ZFwCaijANNL1BaF/KU8ZPNL3Kn1A/41
EvnTcAeJGOHJ/FoDhy7tqOYnA+6k8+YyHAMkrWs1LiADgczIef2Hf5Og5fxGlpxM
O91kSfrEWW9snDPVEQZE9mtjoVU/69mDexgrubSmvtJJ4W/N7qC4E1Gnc64X3uRo
Yz9zFyVvUfPsf0QPDh44dU43GOzuw8FCtaENBEzMLwna+Zigd4/d/PqYNzbn21bA
mC2azlVAdS67EVxP3QYalCEqHwh/O1YBCZT0SzzZSNviSbAs2ZeyA4JIw23PJqiG
2whWMqEMWD7n/nd61SeJcLVwtGrMZe9JvMiVw+0U2tV+BNAsIp+Kn9YvNiAcuB9u
EgYns1E/HY+KxbouBwYpTz6qXa3WhyZ9BA7Oz0nHPJbVlOe1fuUnpOCB/dnLTtH3
mJ/in/mHJMU5bmQOLWGIPrarchAt7y+SjIwxhChWn8zH51++/8+xvf/nOr86mzd/
aXMMwi6IocJ+wmSFHd5mEnER7BC18GgRJJN5pMbkuogroy1fRL7fc3nB1kf7Vi9k
lLDgjCVv74jDhlFHe9unRnVaD/w0Uet2IXEzcXrdkpMtxSwfNnrTz3FOyMNXflfd
AybxhX419RRmZlsmFaageP+Z9Y+W2e/Q+uNj9sUGb7rkrwBbeQ9r5NFyAyR6j2BH
qNfiOCtytZ2ivqnsiZL8OBQw/OpyoWkZxMinl63BKHbJFDIsov3PrlR1MykKwN4t
0aHbu78RSe61iMocklsLVMqcwhu4O92NvSZWPG142E2ZuZUYQop3VTSRmnDS6OSS
ghrHW1+gQvtCN2+9H8tophkYF6nUDvNaPf7BJKl9uO4f7KZWRmJ2oHfkhBZGckCi
/HnTHYkAZG0799f2avASAj4vj20/RD4rxp+G+pVmpdpi5+9PbuuVR1uXJwB3vfni
TYxdvU+AVn1F8k3yTykpsE4Z1llhFo+9taKTM9iRyb1gvIPg2C8hmmCZa29WDaS4
lsYaCnlLBdWSiAhnQkNS3HsYXBW6+98c7rIWgntcW67L+vPGcvAxZdREQfAgVxZd
6vSvtuhridU3y7RaSW4NkCI8qYiaGi2y95SWUAtm+wJTBOsuVpBhKhF2kXnB2AOS
m48Xh0Fz7Uy4ZLHejrzMsAF77ezqqgmP021SPDIW3mq97MIt24rnqcwHTgoOQi9X
Yqp58/ilZ3F1Fbb01mzkjL7U3LbNr2kHyYvPUVoVITwza0Td0eLgA3quq7/xWYRx
GFxlPiGSh56FhBfWXUYGHICQOE143gr+JI1GytrXvh3QO+RqsITPTse6Zz1SS9BO
0VEyeKSoEZXyaQvjs7hZzHb6IhbA8n9mp89C/t/kLu/IvoDX+IBCx40TJG9A3vsJ
eD6H3hWBWN4DhF0Iccw/yI24zRwgxSFw22meBZ/dqQATuUCsqikCNE6cGvLBPt2q
e0JOuhOtVpiiHUWf28PqSK0U5HMEnlJU0NkVo+esOlc4Z8MAjU/2d+u4SLcSkElR
wcSP113TEuOpvbaDkRWVuOgjmttl/iIkMS0Z1aZZpK706UN/UgavTuusmiHftI3g
OHt6+1KvLB+xFGDRDEZyDc3n+tgKWOM5KmlROq162kF+yNNV2jlbK3aboFwaWywZ
5y/rjl7AVdQr8qy+1Q4aMxgyVXTDVg23eXdG1Wxt8OOZg9EXfArlg0HnX7TaWaeD
m8Sg8o+aROR8monusGqd/WuNrY3yFikK7KWuvQt8ngaY/PafRy0WbKkHyKcu+LvO
+NrJa0EM8k98XpHBqxRd2dwgUtf4sE50hBq7NpMCvq/AVfYC6BUUraqSa/H6epdL
0FkmfAkIBikPqjwzmdQc+VJMQqTxVI/+1Ek9kv7hLZOCwZt+0r2pLjcEslljZVZY
2FO5Cs5VEbvcXn4DwZuA7HtmWDSgRerYxm9LTJ7MZZ+yI5yjmbitVEJmhq9R1FQ4
EvIXzK83RDKe7FbZJWR6d9/ob6zITsKpo7vSdhc8FgLP5FPwnlhDJwHHn8j3TNgY
viB0A5JErrVNYaKmvr/T6V5PY7Q9utwSgDnEItYi3gpDUitGdTRPcxEPXNJBwWH2
hOVV18710OS1/bRa9cJj52ViPiCsyU2G6ac/ZPkgPhb+8ewI852Su4ICN0QD6ii5
MuoE0js5rkdIY8vpmVT0rxVljEKC0/+1/YRw4Z2+Jvqgb3D3Asi5gh5vupWcNu0B
ccsTRh7E3wPMCyFPhQ9eB8bN9rr+S9CjHlnhdoIwnTzNb5iQNwF4Gpqy+iTDlhDY
WpAjmiJryOBDf7Y4keE/K3tfmjZShg1gQHyooNmZ101T5Ezn5qSY016Lr34S9C+y
4LOPv6j3eHBNUwgpT0HcGeoyF3CzCWhEoSH3pisljUdOzw1IiGKAu1t8P97UbEMR
JPq6/7PNTuQbowxG8MH7WDNdlWvpSp1uHpjlPlvlh0EHjfJWQCNjhxtZIKXiWjiO
yvB8ly+pU197KAev3zgh0Q8r2Us/DIY+8vI7tf1N45MwOWv9GNafT+vvuu6a5/bc
o6rSE0b+Y1suX08Own8tROwhZECPp4OnmKTbCB1hVy0d/KJtpN/FKOExRG45RLao
MUnXwQcvVAf4MWm+5Ta8yUUIwU0Ok2u9oY04XQO0bi6hcxoaZt69KQx8iXkhPszO
6ZN2Gc0U7vpBMDPLUkUFi8rqzBykrdG9K5Dm+rhwosrGAsxqWXCWA/sny8bovXXC
U7lzwRB7PyZkw+jbyEdiDYK/buABc0QWYy7b9cLsAbVBj3H1EQAoBSj9ThFon9zX
p0wVks21KnQfEYKp9tsuO2Q4j/+w74bmNb+I5JCLPooK0Z6YPZ6MYPBOw7gVNz7+
nteDUiI6Qt4feFbrLwMrNbHZnU7M4oTveoxq9G1E6JDCDF1uOAmFE7Zeh8aJmdAd
t3GGqca0rgbBohZCfV97ocIxTtVoAEgPtxJLE/UfAIelc8NcVqKqYD3NUV5CRsVx
M6Hm8pXmlzToTygR8xywjQ0TpqU0nBt+QOOSpZsdGvyBK7alLX0CAgTvjQQawW/D
h9lMVpbV9+0FtGX3UlMvNlW7kKKOLT+SimWSzKthZg1HY1EFXtGSHYdXpErYeiWB
Vq3/tPDoAdIO4LaN41HBaEqJbFkJkY4j5hG11LkimRqKBpsOpjkwgslJGcy4ka2G
XHP8uoe8EW388H+J+DU5RyRsvikTIVvdOuW4JuA/waWdtsrzKdz14TfLarvnHLdy
uk3AoWnEFrMlgZFPsvXKVyvskomXhEETUpx/cI9mv7vmDVNDiJjALsZTvRjZsmLP
jPajcPhfXt36q8Fgo/i55iD+uUg2zoWqNuB+Qelm7GPcb+L05uE0S3Y0OaSSQ9gS
09sxOvqwvgOzbmCBtMGfMIlvw+mEsZf2CpDEwO3BDpR7cf3EogGZ/u+QGA0t9onB
IkBiRW/pE7X4VNrRpKpmC3QswjDAaRMUGEu3P95fAKc39PtA06tdl25uQBcC8gaq
fEQryO9625A9LlSdx3fH6OCPZgjklJrdLWrzUPhB/t+6a4rHRrXNcFGmUy8wZ9sk
opu0/pzaghj/wxz13qd6nkfzN9k7DvroSHAY1Baki30xlofnKs+L86dBmHVI0V6E
cqg3g4phH2Dccf+vxTKzKyEbMX01HI9hPEyK0KcY0KjoNHJaVhPstd7FetnQnaZ3
hSvS+0WVfGBJ+l2fo1yQUoBA0MnuKINUewnM27Wz543/rIUzf96KB2BWrpHvfElG
9XJR5xd3WdscNnDUbQLFSGHxwlMoFRtm3uEY9eOJBBMQNFZlJ65Iz1UvsqheCJr4
uwdTDy8LHpp5ZXBGagvWrifOOyqtocsPcE82WU5XMdk3iTNNH3h0weSxqUmFb8j9
AoLLGV+VqS62uyZQXftBNHFoACZZcWFYdSn++1xJFc7Qb6+DoYCgX3Zc+8oYsoQJ
q4OCyLShJ076BPQVZqRrbSDGHGQwNenLfLHHi/WF5GY6aAFSHiVKXF5GX7WtB0NT
Z1c65MaL2JuQC3vxjsL69SBKTAB+hPvvMmPaLahNoHX6fX7AIV6DYQiH2nLGJYVw
1n2S7ghl/ubUArhAPFcLaRulXbYRWJjVJF3sShp9cXAE/nErMeqGwLtttzeORYxH
5gVTcAu+4R/KOv8128IG+scT19O8pqJyKNTMdl2mdU9yDNdGRMTELtQ49wexfCLv
crdFTXpY0OREm1BEVJ5PVDz++4BCYQl6xti+OFJQaqrJQIuaznXykVT6ku+kQ/R3
ZMvjOZoEUE9pXOr5EddpOckCXPOyImtueuwmQtbJV9QpxD/07J3AKaInvkVqToMq
2MSvX0qwzOGZwyYTSlFfqVOGziREJFUkTxSZmEJVl85UVAGPhtx421NcSrjlxW4J
zduvf2xdKr0A3CzAmeyPoimxDxgQxFi86TDsClZ0h7iBt23tqQvjHyfQbz9uLJ0Z
5Z5AZus8GpIUzdNrx6te8yD3mA+jgZAnx8QofK3m8eDOjwJ9g0twg0BqQhGZ3yD1
0CiAp/KjCkhArSQFW27SKxB1DYtcigHSviuN1krnAyvYKRHYCeEuSqwMlscEOalZ
ihg+pp5fcYmHI+zJErXnvQLKTBw6xOzxIJ2gX6D80GE5ZlwuIc6k/c46BvW1+17c
FI+UQvor25muO4lieLLbq2Tz5YCrW9V9SIpOJa9WOJ6O8xy7trPv8Vc3CGe/hjbH
gkVM69W2/Hn6AX0dND/+C68txWPGe3SXSUjaCw7d5aZYpPS5cg0r9HJ/gyK0GjmK
jS6LDyA1xNk3daqe8/TjAE1zAUO0wI4btynG529lv6gybqr4K9rUzLTjQSC2vq0M
GJ2P3kUutoWTVIViFda9My7DreXyd550Y8SdXf0mtERTdXQVT9neg12sTAZt/QHp
6ZAM8pBT+rkVnXzSUFZlL6A8Kol+f2inLlJI/P6JTLPe5aQrvcZfwHI7fwY2m3nq
IFy+IcKl0j2b/Rx/XzKCzMz04xeVN5QlfsEA8umpmtj40U3Mtxo9z+VYMeBVXZEl
wpn0GRcYFu4Oq7mlvgXnu+cwos9vshOpq1EnHyGogcI266VzMWR5CbMe+ri29qjn
1ctDqGAlNsiQ/u7Lw8Ad3UmMQWzgIO2Xgl6hDJH+nQhhHZHOIkvZHDr7rvzuSIQC
CJw3pKKuqgdzFTGQfqAJPFl+tPejANndwcMrDEw2PT6yGjCwmxo7HEbwbnnNY/TZ
FqzmxroeahaiCz2XCHGzKjEaWDGPJJu2JqesMwEai4362oA1V0iyF6NdU5XnuFaJ
DEnvniXgnoc7e8ZxK/Z1JQ7spp9dgtpNrY1WvmHUeQPmTF8/EebWlS42IUcVIe5m
EKf6oEL0mnnq+xG4sq2UCF3dJiz2rZ2B1S3/eURAkrLiXs9rvCbKYErdRLDe4w5+
DmX8hbIT1kuei6Dx7fIUbt0XGIe/Pt8WaJIh5i9ZtAepqEtkZGWd1Whu0rg4vh3c
Mw99z711+aOJhBgx1JuCsXPqNDDsvzTPi0NNPGegY8jympFwPQbqigusCqCjSnD0
k21hZutls5TZc017ceMfH+R7fhr9hK0NAXErVu44VzLQFQjdolf4tKZyVL1/AmO/
6HVEcyabFYECTP1J6bvg0QB+utoCgxhiLwASJlDwimPZxkSit8S8tZ0842ng9ByL
lpgaDdzEV3BSNAYXUIfiN5ZYGXypOp09TN+6atW5k9hXQISrKQ6z1hu3mo4/0HxZ
n9rp7sfv51VxpjsvyjESkI4mn8ymA69Btot7ILSVa7R+vNDJH4ZRiSxsmzf1hRHP
28e5JU8JHYiR8PdLHVGCM9W/Bxh3rhWLNizB2Mte48OyU0BPWI6JdoYnFUOzq75J
hYu7CYY5fzyWvq0O8XHtkBiLd7+xnDK2z/eMxWGF3rOeYeE2w7hT+ghwYq6Ze5R9
XFv1lacsExHqKYXobay7x2V8OIsuhHiftSej1/T+SHCX2O7meeZAFatGQyi1niQR
e/uvDiU0SQvQQ8bvOwahuST87EO54BLhsFoyrk+QCmKZuqPX2pRhlG6uM8O1HnOy
PS13cR7YG/cqU2aO+3zUAN3kQR1eNLnP+tgDnFuDWDb0mG+qL7bEmNzhXssCNs9R
PjoFKiRAlj8qC+SfIbIWew==
`pragma protect end_protected
