// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HfjFJqDwcWRTswIPq7zHg0fP2ykSiXH/7p0W0XWfptqD3z9nPk+eizy1wjvq
s2YFJqzbKv5HrHyN74+gCXwQIjRFE72FMBeN5eu22EfLugxOpaYmaQCZs6J4
+616g12QG4CVRFd/4s3QYiHBJR6W333oi4HyEbfoaCWgFhT2CNT9WV1My+i/
lad0R+zLsRkfSDkVT/d00h/Nt4uSIUDjqP+AFpXgs6GqJdQ+akjrk7rUf7UT
HYIwQJFlws75g1eCRVAk/yLPNe09CtLXDhQT4UP/FGGAKaMLL9HsNDcVRT3d
Ybb+ow2HEf4ZQzysDvhyXgH4XQo1qOtAa9JELyAdTw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hhQ03o0raqH3hSwNiPgX774KDUmqh/nRTb/5ASYHjG00CsddlyDDgey0iViO
6MQfXzkQ89f4Uh0eYJ5iwoYXDxFMj/JguYJf1/vlNd6wJGmQfcgJHaGkwVHz
GEhi1qEAGBvi10+RkxKiMrFmUWPt+4lRaJtell9JPVrB8yJWmIOYwJcaUMok
BU+SpCso9kkHt7+PaWjDSJwm9hxR81YZXkOkbAhgfbt2klSQmOB7T9/lMi9e
gdZ9J6HAROtWoNbTsP5Issm8lnYCIIfRkT7nsp0A0H2LMthDbusn5cwDgdPI
KTPR1UxeBnDQJ/cI68OvcJ4mF40LUNggq/VeWmqXQw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rAvj5Nsap4Aqi4PIyYBAhRRAveGPEcK+15oMDyqD6ot68Rfk/V4b4yzmNleD
fsT93iVRGVrSSFFvNf+d8lRWZ5PC/Dy9gaWzMhcCvvuryx75NPbrAm+ummxe
+9yfeE3dOmuCNWLlq8G7sH+jdJ3F18NU1E9W1MG69f3BED98gLtoAMrJMFV4
Llh1V0GcSkfz3rkeOnCGec0dctSKo222TYocpporNV3czmR5Ll0y88x3RFix
KhRFvHdGwkDFfQTiSP8LQQepdwX3ZdM1D2sASjD1VcBDMoasSC2MBveIpjMq
FY1r2rF/pyXCz5HAqATXJFSkn0CkbufkNDUNuR6J7A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XWocfTdY76fDFZxuQqlpDWteiV1wFWK4mJoZQ4art8hygKYthkFvYHGn1zY5
bIIxh9C/38RyHj6tK8hnLXFKZlGaM8+zuw95gexOavbRZZh5TnZk0oYHIF39
QVy3NUIT7ysGMa2AeQUhQHmQu3v+JDBkLzzOA6aRFgbxwg2+75A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mAKS2MPc9KdYY93kHeOY9TdIfJ34kVLh7Il3ggg2wrIkv6udIN9G+aRqExCF
9sIch4tcPKHOUOfRQti/YCJ2jZoOekEo3yEB3djCHV5TAhPYeq5E3cMtOxEu
3Nzh9fs9rBpu3Djbj2t11GwYT1HdGObVy6bp9DD20n4cPoc/Oyq5DS+wOSHe
qGE8N+McfcTsO7fta4lkOuSJVCHCt0WFl+gbvT0uGPRulp1D1OLbXKb3R+8u
/uABUrLeqN4enYoRleIYgOrHxWiXCgzzrY4yKLrecjdJWIvEBmhp8uma73J3
QDn5QcFVAkMeBfcgGLwstuE2qi5xwA72hAWp/aJmWMDH9K8BmNvC7HXtqRXc
fJHo1BAqovyLnf11Sd+C3qmGWeeeAr2sqYH/fTCsHEw2YvQXqQ9J0VGnGxd4
pvawGO8AYjMcAGy61ivAcwIGRiTEOQYckrKuPoJR12trbZQzQItCh8V+O1Nu
Wv7fvSCMHygvLZb4mKiRSk7CL+edcQGm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H240bK6tXMu37pn0q7rxuXKy/nbIDpCK0B5d6MR5fO/yhujk6ytgU11U92HJ
uJGunse20y62dVAgRx5P15LllmtVbgNhQRPKiBFzC4Yj8L0NNNO99wENqMZw
KnTd4il8CfUNqzDeIseB9faCM8sQWaDSQ/s/O3k9LPRhllTnJPA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kTNU7mz6xtpLeJybgaqp2+na7q2ybjh+5ijvz3ws3kbE7D9kmn7r5bqfKgB2
6XEU21W9bGJ3BkfJB8JfKPDeLBipgh2aLJBJuI26q3nqNek/dVxQw/jdf2q7
dJAqOzvIKZW5SnX8K1d//Sk/IA3dIFobC7z2DDgUIDNg0NKCY9c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 65472)
`pragma protect data_block
DlUr4KOKZEK7ukP2HYmsEEJrLMVG+tvH7MI4N1KtVjSPxiH1SMMIs0zaePwn
r8R9JOIDMg1s56/QjY5WM+Ye4PIEec6eD3sHdZIPteYhAeAxUiRgn4ytTMaO
u7rdtMUL4lkJ/SjtxZcwpdJfUoe6O1F8C1Gmuw0lLkdmr3gQJD0ZES9eT43t
i0qz7jEW0ullrzjJkfgAmjXCaWyHRxUSL9bgtDjdkzOXXaSCiur2q6U2ncVa
feJfaIpTtxwqSnSM1LcJtwoecpan4+EBjGgXa/FtD7mJ6myibxsK4Wia7/9H
+V48A1+hl0KSfnDuZPgYhGaqlLZHxlGgYqab/We9wIOgHg8fhNmvH/JiM8YM
V68VeoDgsSHnvgARM+lSNgz+b8GWOToCrWCpraHawZBw9uQPieOU8OKgtATA
FAQoE5Y729kHGEPhCOT6pS3yYNrDys5emRzYA7WLF5dAl3O2LtlO6gnq1lFX
SxbgfOrb8ysnV7m9YVEM0MhTRZTv3EUHO+X2i63teaOTvq0wKZ/LFBMyALuR
I9krJ2lk+8KDmvI6D0A2fnjKdD2hjNNXvqywZt/0eznW4InB5j+4dMaVeZSr
xrVTVohvyBhWjiyeYuPYTAxSZdZZD6mS6AlfyH15J3arkrMidaGUaZfCgO2Y
r8Z4Q3FSWC0Ruj+Fx8/QikamoAADI+H9Ps9Jtg+Xzfloo3c7mGYZP903LO6T
ABChHhwRR60H14ejOSN6wypW/1WJooBGrC8Q/VuQIdk4nSSF5IGyMDEnVSMI
V9LaQjEKaIIsw/lfJRQmbt1OhTMGGzZf3iqN0qVRUf1C1+EMNSr97aMEw4zi
9jPm7g1fJcwHxmnR7cHhRwvajHLNNRG/zGs8XnSyDrB/tnVT0wENkhAn+JWL
zrsiKiz1pRThEKUarCXXa9zi20ac0H4q16OVn3FNFfOkzlnDFsL+BsBQby/4
pFp/hofZi1V2pGfxFPs/PFp2P4aS/+hCdbWcGPDcMklp/AhW2RH2IF5m0n0y
cy/9ZSmF3Le8nisQsPSLTQEi2CCIVdMkAnYp3JQShlJ8achvOIkbV+izjOnj
08qxEcQCOoasnFVKWaxb4Nr3kLtGjUBgZU1AYgSGc4pC/sqo7mZ3YbvA+4Dl
mYojSbr2AsBOivedbYg+P9+QCJJ82M+pZKI7XlptJjUYfdGq4Nw8OAbA8KAq
0WeFNL3H/qtn3+Z/Jr9TvkLzjtwyxw+I85UTOMeLEtlw2Bxx6uLEDlkfwrrX
la2vagAsDhmgIaw704xa1eSU2ymaSRUh2IwcaUC8cguIREvM3d53FE41sjb5
h9cFEqe5VsW9lTLCtVOgrft0piO4vRU0ZJ9FBkv3iF6OCenunxJDT5fzVZiU
aPZ3sejv8Z4xDIJk1ZB6eUDyY7Mbcw8+aI7Kb00l8J+9TtUdfqUv9UYl+rb0
5oO6DEhxGTZqbYP0Xf07GBBI80GXU55x4F/ey2Zo2tZe+SZQ3iylsLUeR+4m
e65Xb/gyrEeVMUzXYEUNnq9yu7ZRKCNybtqF9R65mW4tJS+ZjcwLahV9N5NO
p5xR+Teo1DrqTBCQsrwJ9Bjf0iepafRvQwWypQIYMBm5tSPN7NOhyi49iEep
oo7ZsnuxzSjSESfP7UIN0D5WRVXYVrYMHnEXqABCU/Re9AGKWQjxkiK+d2gO
GXF2i1yPhTQCfor2JFZgQDUKzD6jxVrnZDo6LWh/PZlBYdYGKnAxQIar+6x7
JlfbXCbw22Wt0FtkzRuy9GFfXrnoiLHfK6CAx0G65pMZh9BjRGx1uA0fQ68r
0EwzbzoRhyS/kMKStOA8vOqhBthLrN74JNyag0Z0DJ7ySwAMAoEVVWqzj066
jd4nQM82Frcw9J5JzWEoGgrx1cWIyPRrB3JvHYYqYnX41DFWmBxYlZHXieFQ
TDKnko3MwrqetnPzSyGLondN/IdT3+hcWejhX2Q+ynDcwqTHm481fKTpFnqV
o9Ij216YTU8XgPSbf/s34p26SQ48p9GGHbFUuzGQlRXmOQ680UA7FcXFCFyG
/vyrQ5Rfk1TGJS9Orufn/qPPvzN+Yrzjt2p2UEJ4Lisj7xVXtkpwaLtJ7oq1
VJYY/AXUDi4BUPqTgnnk6N2iybjiVOtyvXfXqYe+Panxynu0QPmW8BV8+QU7
2qUtr/WRl5e6bzmDzhCOgZQTJKCbXXdGNpgXsLvixwflG4Enm4YVasTdFm4K
2pM6hAcmnXP2zBEMqDMorx3gFPKhzsj9TrDdfGAiwOZqw/YYKa/ivbBO9Wuz
JfD3fQpNlujbm2HqvTUDLaSYv/WHlCZo8Edi6rGYJtS+dLLcLaOhmYP8WNB9
7kLFCt+ak8IbleMFnWp9oQ/SQ+S3IJLZRurkk5xw5pnWCi0hMrwwv8WVA/0v
rtmL5oqEsckfhH5tekKS3gbVVxH8zamttC4zU4IpVUTYmLchNXPS6G4SEl8t
blQBefN3ooWN7HI4YOQmx6IE5qE97m1M4pys8pwtKW+pzsaIx34KFICABRAd
lEyeLRscV+PIRV9zrGeHOS08A9b/YUVYh9Bbu7Q+4AdoiFklmBoL12JnvbXp
ooHJpuOhuz6ELAH7dHcW2FWl5Hp5H4ypvRCegwSXpyoER8St710KLTh/pdgG
NZxNDrPcWpTF2I6Kp23sA0SVCQDdmHl92pZ5PuO8zzLM9ZdcX9Y+HY3qA5X+
jP1Jbu2I38ZqoAAkCTewwdd0iVVSvqFV7W00qUftZlnkNBQEg2rxNlTAtbEy
9q23+6Gzi+xaJw+Nzy1S1ROKO4//n8leSYwiyV5nlg7Jp7nZX4QV6+3rV21G
V1aMiIlF6IOLHehJFJ80QWG1x3J2vcy4aeayWSrBPltCufw5rL8sUk8JMS79
xCRQQH980rG5WuT/AeGELjdJdsJmXCmomJzD0tSrRK+7XCTE/2OyIiudSS9E
hBidffrhkgjloqQLQJ1yNcnB87RJNtSNXlLKUUZ6lXj0F2a7zM1vjZQx3Jqg
1A6SOs65Dm1OezXUxCB0TFYMcoqCgmGFa3aKro33a1jS2m5+Z4BgJVOtMXC/
NqG7QlytIg4RIUl3Q0sDRAWuv8OniJf3epOiqwqgFZsgMM9RYz8z6fvH+Jpu
MxWtUdPdk9MNxvMMFW0GwuRsZmw2sE7OQ7wexIDNwclMda1CxF2vvsQhSjlj
pvH3ignScTzLlfz946WrgSibSn1YFkHwG9Tr2/Ud6EMwFWQD0ny2Xgxk6bIs
vTNtIIN3lz+AR8HZJe5mcPirTYJQsRZ0qeAyt6uxbe7aHxK3d7zA9or60UG+
vDRpnjvZqQBF+DqAkBrnbboNRQUmaBCLpRpyLpgQkMIvX1i9KJr4Fk+lFOmJ
OuCGgjYqLxtEmqIRBU6Ch+dGMfZFbrfZjde+dxhkjtsFCsAXK6lXV/KgIuoO
j+B+6McvbE/f1Zy83+W2/V5a2VD5s59R+iwGhBn9Rh8qmgZ2Y9j7ttPEshbO
eaF7yxXDeCS9YL2PmnTMp3q/u7VHGThWBU2sWdjcU821gh4H3Fm90Z4JEyvm
lig2bWgf50e9Sl7OzJN2dlsqTvT7Ac3KOzHF225JQLD4axyTgTJmdwc4bl3I
nDtOqrWWhq8lzwK6DoXx6cqSvTa3+DITm1oehbNFRi1Jl+rf8Fr+QomFcsSo
4VKjLjU/1PNOKhbVQWsZdNDkhLgYv5btE+7Y5d/oOp1VWPL3cjX8CK2c2yyW
3Te/ObKLGpvTwKyI/66YwYeadjNZnRfFMq7GLTUn47HOWN+Y5Ynf3YWjuple
ilCe3+8Rg7SoWrOZuNrU8s7Jx85k5MysdTTx81SFjAlo//29lja4bhpChj69
GEOLnycZncufInqBn238ZxakZxn4BEEdFYwa9rJQ4y3YAsxMpM1xHRs31zTU
KJEJdySyL/l6Shlh0VFRVcNtMIiQGJxBz2Yb6dcGfEfj/itsTjYVD22QRL07
qmJdBDjHVlTMHBZhLugMPWc8kjrkGO+KdKNSlpcit+PJKgBUQVfazvl+KPfi
2RC92QkZ8ZVyFMQxVsr3XKjUQ8KAQ+ZKwZc3UwPpTomobwafKw1DWOp0mT1s
wL29QMAzJ609A+SgG4jxyLUk12wOGzkr+fRGs2WtZfAZvO5h0k4iCf6uw66y
Zom/EN0eMsTFwYbIMlJ4yqizQsKTnwEla9mlySGkcQGFLNT+Tk4vCmsHyiL4
A4OgyEsJ5SIa10g6ETf2ksvRbyyq6kTW/6QfGUyRz7Ot7W6SUqD741cTPojT
Sp5Kx0dNsiai7g9er/hXj4ui5IEk82q30yEyON/1Nab8yWLYTmxEVJXcdjTD
1EbrSluTE70Pj1eT7ujxlB2dTRHa1OojqQdrqdOZf9JS0tPhx875TrdYXXqK
zsNcZ846ETaF2ow+kHn9XrJmFge3VMCdTBS05JswDlFX9TcDA7SJLTZi9fY9
DLLT3799ycdRvvBu7HYsE9EmjVEiAf4bHhNhWNFhRxC/lNoQOq5A+saZCDa7
QiVEHjPJ9yljvw7ZmsPQTugPY6JOMvUXX5hzgwVjLg5TKDE9yiDyu4alMY1m
LWQnbbWVWKzOAxFZ9cTroRDYt7Io3nZn5DJVF5vwR4+qjidPU1X967ULp/B6
nbKxl33tWHGlIpn0refdOo/n3znsNMgEudAkYCJEErOKWZX4slrY0f07DpJ+
C2iiQ2Q2tiexA3OMWwANCvEZsQihSpHFXjP4W89mlhXLcElS7YFMbkAtM/hK
zy81Pv5K3QhmWrYZpw58NWqBsVlntVyXiFCPW2WN8Mfn43lBsW9PvFf9MxYO
8rPT5F+2ogrYg9Bb3Xw/PjE582JlQNajAe3Qplk9/CtvvqRtLryeeBD8RH2p
gENY+jpRj8jRgM1KDZkM3Pr9RRL9s1O5iwhN6+vrakgq9myVK4znMmRGLwDU
T8NPXk3SduNP9g/KiYQ9naG7XrxZ2ooES+7FPX+pxRkV6ApfUHOfN5M64DoE
oVlktuToZS5YF1fYwo3xaWauM17H7ArfCXrJ52hrSfW4kLNtsT8Yx78ke8Sq
3eHKAZ+JpPjtKRBbfiTUfeSObt/gKsoFFrsLYGBtL1kkew0bPL9ZEI4K1/zD
p9xiF7W4o4iLuXl2yHW4P5PcnFfG7kMw4SIs/wkJlVpSoX4dGiG2/CkniF66
Kcst6RcB0/FRlb8NZ/2HpnaW9RZnP8EaJToaLrlf/WGlRfUFoglW/EmkLFyw
IL447YXV486b49ZYvz/nf4rY73bwS7iH9H4Bi8z9frb7ht2qVuvaOcJco01+
AyiKck6YqgsD++0bIwrA+16OcGK/xqMMA4FHSY62cbL2Q7YElxRU+i13qCLL
2H9tQvrnPL/+2+fwcW604dimZ5eXJIXe4UOJZMDImDCTpJLnwDCzVIPH5E68
mUv2gAPffjHDC3m+SZ+LDxvLnI5/KU/DUYEcFocubFBaJbpsDTsQX1mKxbHr
H5z2qnBmXDy7WjJV9H7bNZt7xZ0BLsYL6Nuc5PHZ7J0Jr2G2JRdwrSMpISW5
f5rOHklkk87GPNso80V8NqD2+Gol74StLZZe6uBHoSuGqtBz8nQ4wFaxbj85
k+OjxGQHaX6QNoHugZQZleJSel9txSFTP7164GtQafPMRbHzF1xHerN8w2IN
wlB4S2W/UgVBcYs38LoWnJp4wijC2EWKBTDVUTEj/JW+GpHCTQk/8e3ybHd2
NwX9sz4ZqrTQHLZARjJmb5pH0phUre2rsWlXT4gzgswuZW3pllLElKsB53lA
uPaimnri5o2Ulvo2mgb08sfFpWmRbBKN/1kqJsaDpy1dxrcpsJyTzkd1uPb5
rGHBwK1MG1gh1Mda00B7IL1CUoPnyXovaJPpBtgbDyVO8UYonn0Ph/JZLtcB
cWXpKuMSYOWNEXGCC4JE/jGrjp+xz0pbSQNwj3rGukfD/qfRGvcfdYggc0th
VHAaQ1ZPjQSLCCkohIw2Nx07VXJ/D8M+CqwSyqK0V+wxXoZ3Cbz4gOLZH+wN
6gY9q/BNR7eawhXtVfSij9KL0KiVHLlNhIEfBPfYxbXvoFCBh34sfu5xKOIt
ecdgO1VZcM1Z9rLlXnbdIDQYfovRTmHEcNLY1zfBSzyI18kuLqW0mfXsXCHm
Jid1AAae1Mru0S+nDlwvQSAOZhF8dVnrCsrzjReSrfNvIN4mKk3g85SaidzE
y8mQrX5hw66eGqOMllD/uz7NRM3wKAioU+eVa72e3C7JYjpAXn9EhA7QbiY2
9NrvIMcEHY/GCBQ0MBqyFvuyTOmH5WJeUQVcxW38XrALoX7o0/t066FcgqTt
t7tGacooeDSZqaGXqJR1YDIDIa1e87rP0tvDMGY6qzmacCFUx7Mpf2hWc1Jw
5BVQ7GamL1jlQEH4737teEcAXhUVPU/4w0kC/9NKonncHTITFo3Lk2OJDEh8
BgFsCND6hEST+9fhpT/J0r95nGaeO+YQCwxTclHPDj2WeNQLaCBZgRYTbK65
3/DFJIHsor0N59Ro8Q2fdoDJq15w3WpS6R06Zn5OBeaKg2xAdMMZXSTyq2dX
KcNWm2LKCgzf1YSEbXWdXp6N4QNNf3X8BVmAnN0HRfqQNc7jVZ4WVyei8E5H
3MKZCsD1/viOQ06Y3bhPNQi8Vhxt5Hb1/PqtqNZ2weYPXZmA5RD9ygEDEMoM
QdpmqnJVxvx4BRsV1mvgcIScJxVicDS9+ke4V9XuU2m8BZZEuArUZXcEgRRc
CcRxHj6QLoXB7qIztcZcpDd+2gMOB/wAf2Mg7Onk2XeYrhz/mDTckUe4Dkei
gN0HSIlCaCqVCy+dKxNDFxtmLzBXeO6mtEvZyX91SjqLQl/vmqtvVNSJmk4r
llJXmbVo3tcVvP03KX3aCrmRhEp4OClm96yFbzfT87qRsI8SmygDAe6Bc6DT
8PaerWsIX7JZO6JsPe8aZd9k3Kr43IpkX2+RVj5gnDEqebElPVnCP1qBtYuY
7fZpQJGy9dirSraUb8vt9uwQzrkJtin7DS4M5ZtRZ5iwyco4cu4QkRjjot01
kObo73Oc7ZIgvbP7HgDnkAxUPBSS8XCHpYOeIUMRSrv5inCeHFB047WfHiyJ
JmYYlb+1tKDLy5CSROX9ArvXhSLjstvJwQ13a0sPZ7rvLORyJxQAomBcnqar
1IdplOnB5wxA3Yx+e2Zhd6xay1tp4Indi+S27C/gpeIEpGl8Ucs7Oid4KMch
q+C3e0ob9YXB6ztWsHUUar2GwgIXxfD2nNZy8+94dDrllkxN8YCmJY0HBfHT
WaxW8Puzw29qW23UV+lxC8mbHZ/fro7WxueSS4LtpMWVGgkAEWbWvm/OYWRW
VekkWg4S0xSUtu7KDNcEi5+ge5nHI+I+kdGJ7OCVA2ESDzqUYDjMIiEZa4Ia
PtY3paXIp3V9o39CQZKCTTKvpnZih77KuE4TdXKPIv2e3skHzk56OKost6tA
JbqMr2o3LEMeGprbMHWcQch2Vt0MOzJfQyv2yfkoBNCNl9f8mMMlk/RtS/Kk
eU7LmikG8CPcakLE3Y2lhZhQh+i416TkCWYt0XN4fsfnJ8SWmLwBPFJpaUNW
c+TGARoCoDwmDxjqmhFhfr1tHXgwLyJllhVYfs7MzuIil5pKH2PDHyrf/7LX
+WRe8U0OAtAUBUJRbhpsmkFn8N2fHdXWA7YAyehV264unRVMHeYaOzs2Q1uk
y76OmV+PFwKcPCU98Ii7/GGgrN5SO3urxKG6bASxFSF1RUmV26Xx6TIOx+HL
B76A8S1aI7v2nrw3GGUEJV13KZgz44Sk2AwnRJdl5dSSPCZb1ENjJrdxslWu
YwPQX9NQAqsqQbZH868vARlHlOPU6HFqbQ/+Dj+83MjLkzM6eVJ944qbRpzb
RH5Rolc1phkPFcYPGkVNtK6gEutHYRprT6d225pt1+DwcddUddzWD1m3Iqq+
GMSpH0C3NtJiYrHXST1XewyfFryi06+J7l+pWe3zyGo6bu8ltlsD4x7pUeW8
AMvrttr0hTYiJJrADTv526ewN/kAn0LEx0FGoXsdHogHM9h+t3UIJZetJa2F
vqr6UxcIdaWPlZxctEsAgseh0EpWMR+JHIR40O8KhJkOpxFL8izXMdtWvb5B
cIc9siwvUNNboo70/cl95C7K4rGo2siWMWG57cWW9SzZ+z0WVFCdIDaqwsAu
X7o7kahgWUcG8sGVr6z1z+281zj3MGRX8UzCMoOCNpGgKk/MWluq8ROYaDNq
QOmUy+TP25ldesZ/ipZaM/UZ2uwicib/aoCKzZI1h1uBS4zrFq6kFYtcvU40
qWa8fLvRnZbVJzgR55FH2KG/QOxM7XDE1ekAams32OBwE2yfRbZK/89MFlF4
r/wmdAsgKx6xGKNRQvYgjqSKUtWPtC4JppQnDneWoFDsadFKPGYgvi6VHvGM
yaIirCC1ZvseySB87wZaZZyo6zOTnFUi+kgZZr0gU+OvvVDP2ABBLLmAuHX4
/eyKCVemzlfcQvL3k7FPQFdFXh3T1H57OhJfmDDkd3qhwo1A82mh4AvQoeHu
mzZEc3KWlQU6aAATgELQMKQR3ehsfb/+e+COvj01xpsDgosyl+t6A08eumWY
oaz29cHm53Dy6PswGmLvh8PzdyzOoxHvaQKOVO92QlSXerIXjRSGlvEbWCE+
DzI1FSwpQlAT+t0gMyiciQLFDH8ZqNYKCDY2xGWwj0ZuIuvoxqguWRLi8WhY
eYM/kZdwrcG3hLyR5BQmXytX3EzpVR8/hQvEOXYw6Frl9QLflbF/1GLaAE/n
jPT0TuzP1NDdd02LB+SV3rBigGopXJteyIPxMoIt8sTjjJG64JfKXhGVBXCM
NCme2d1lUZCMna60IhSCvBQhEsV9rsz59mv5MKIfnKIXovd2Mjod/K/UBClu
CLUzDBJ/x7Uu/zhlLPVgtDJN0VacvfQxv2zrjzraGynP+enW1VIaJdhJKV65
5W79IummJ4/aAz9YcwnO9L827PeO7NuqFzVwEzy766qps4jiUJzwlOBYHeFz
NwRe9SfnVVUwAJwGPTL/rELHPxeVPAQCDNgegJGL3Lf0Qf5RU5N5++ql4CpK
GPJITBpylmCa9Du3XIFEzEign/h7KFWtBKFXxjwelZn/RMafk/f+gdePZVX9
dRzSh1O/0CeeKR8aJWMSjxA70R0slHv76ESn4TPMAfWUxhADbO5m0rC0cMja
PrAxFDOvPvHYsH8/h0JR8xNOH7AqziXIse9bwT23izjCW5WLvsAu58W5F8E6
QIUnciylOEsOXDubpjQL9uviIzjt3f53A35hNbUCzjEjBrtFACudNAMdrLO6
/LorS2vts4JHznvlVHETeDfpRVJJXlWQkQbb6bCiqNb+OLXt3L1/eXFmiWey
GKNmCWlXF0hs4SKKfK0AHqLOCBNvRCMjDkGqyk3S7QK+Q4EsSSP3yFq+2LVw
NpCWc9HN8SmGKBiwQmthzpl5F7Cb0Uu078Kbj0a9AaCWVBSg6ojpdtNbBdU5
T8QpSds1Y2bMENAuctT9olCgU+cDJnsSe1kIuxdWHUU79lLPmFjY+zEm93RZ
pPjGbeUh4Y/YpyvKwH0qTz2QF47NlN0P3NseC9VLdulNu2UpJKpNZt8ZloyC
95oXUBGzTtmmm6YvsTLIi4zWV9nqI6kAbeuinquFU/dJ91Xhf+n9TcJWUmiW
XgB0hPNLfqBVofPoLQ8RZcvst+qbjMGBjBjfkqs95bsAvPl/eL5LAH+9xrSE
q2FfdAAxbm0RztB8EG5uuSFy3l14g1FShDlWHt0NdXS3Qz8sKkECDE3dQwkS
NBrKMqYZ4RSOFwNnRX3QpZItZWwe2BK0umjFmRgwi/W7ZidUgCBCG5E2YaR0
ql10JeDm7+OC4LEGo1Bq7G0eItR0z/Zgd+hPEWrvaOPwHLrzutOAKQc4fbyx
hyUoQCWsoUMPmHuWL4xhtLc6FiB5J1xX1v+Mh5qbAASRv4s/lfhlZpy6YpTj
X65SRtYFSdvqEnUoOCB67iQBWvGoiofLS6HQXq7cHzIYFSGjdGn6PzWo4GTq
csz8uUryA7/gyg1BqlSHNjhc6Xncv3Rcyw54M6Jzsgs9BNwnmkOFcNKcL4Uj
e3vPdVW9iZ5b18bPtIsKMTw+8TFrcSs5oHNLvmcsHS35w0WL8HZD19go//3f
fiOvbzESKjecJnwtu8304dls0kmahEGVR7vXVVJ3p5Suuog0+4IzGBRUcsTK
1/LquMPrIEAR/1yv4YIvE93bhnqdGbZgb0zS4gqKA/jsGRAjs3La+qUq6bCz
ZJhHh1BFAn5XnxsN9WGEVWumzmQTDa+Erd1MK0wC8Yg0ymz0VA5/DiousXh+
TsLh4jysi5XV/2WNkUpiPfUwTR7Z7P/caMrMxqjexkTe8RaxyT80FB5ZdPPT
ycr3p9SQyviCS4UzyINQOvOh7F+FjDZBAkUfh9On99hT9m97Ue72VfRGY9sh
fcTQkmlWtHWKIutMymRA5l5eTQ3fIkHTWvqh1m7FAmAdHHxVM3K1HFE9uK36
D1IXze1azjsfRzFD0QCzzPTIZxZ9Xb40zFYt9xevpgxv6ZQMHtpxoCWYunsE
c6G6wAu0yj++3tkmF5EjrMqofpBGYj49v7mfnCs5AupA8LvV0iM92nJxD37K
5wPHupus/g8SiOb8WYhQzc+X6U5K84GYT1+namglclqgrfgIyx67Fc+pWeqB
XXT3ujUWgq8E+UVW5Zh921ExM/idwbsznt7CojVz8DdCMHFzHBpR1uIJn4uW
Ols3bNhB9fp0nFLVlRHpoJ64D6q00x9iZEByng57Fw5NUExzwY7d9SpujsB5
Y8Gi0x4NGUP+VSYjmAgdoGGZOJ+Tw6jsXjk5yI5irm7ED2rhTtM8cxvHyMmZ
j0lmW/EdjwX63RVxpG2b6veNokg7ojktYbGPNSeZreULNPF6uIzIzUmkJJlR
/WyvaGX4kmLBLWSRJBu7k4EcThTYQWr4QXISOqlvHS78bq8Jv1ex9rcnsw5O
Mmw0kgSSWXQKmYVbQ3I9yFrIlME8SwVPYMshqvp/tWcFYNTxWR0rEs17XwSm
P7hJXL3Y8JupqD75a6w6W4y510QLgQIfOtvPLOCRSo2jESfvMCH+dFMwNs/+
HaXKy9ACefUqZOPtyqJycQvmkCanOCPWDGowJqCzkU4pwKiRfVCQ/ui5taPH
/dPqNjFJ/MW8O9hSx/uS8XHDjsmNg16w66Z1imfm1Ev6IIXQEhhCpA9Xaup+
fSjizFxl7NeaIwWwjtrr+hiDMnR4RhcEwlwR5WCWushPnLHV/bAdIOE3SBjs
X5D6v0UUt91rAocSruH8XZKVMjoGwYiFSaMFhBIHxAxydX1i2WqN5aa7lOAP
Vs/fI/l6mG4XaTVHQIkEJsivv9MCJTqEWo/UECIS2psbntPyYwF0rlDsMEh7
rxNbgm47R/6Jfr/ZZh9BE4ldkoCkwpkjAbBAJF+C/bzdkZ5kmvlKJuOTFrs+
CWiLWV1rzwj+j/mlFKOfLKtl/JXcdrfUqRsxDtbrrLE34lURlw8nSBDrRRep
ft8suqc4uUMhr93xsrUiBlXmtIg6kApITg7/CE6vNi5d9uXrk1aQXSbS42Vh
2PG34tFNR4FM0ze/o9e9JArKvlbBmU7CRycTVydBdzf1pEkN2GIY3jt7wuzP
NwP0S2pErb3yybAWDYDqWC+ztRieqGHm/qNpKCkF0VhzKpyxHo3FkT+MtLyg
LS44V9uzwIv8G1GUmMKcCRoN0sE941++fMD34vLrnc1hlQUmYQJJSR8Kw6n9
cs2iWmYTgxaBYBYGppiNNmERBk9Hj4A2OTLxcT/mAFWBYnYzmhRq31zl3KMW
X6+108JBa/vQ7z9bIFoBmjVAEoZ9GwEBtrmbPlhUX9vqwi24tUJBAtX438mI
OKCyGM+bz2DvVWT3rPWwwCFLTS1DhtQkPMc94Q2cB8kJibhEcIsvzclPbWfC
rGysKMaL3BUUoxExqtX3tc/mpiKgIgGsT285uedEMsy+hfUr3af1Nwo6OUDZ
PfEWPd1tMjXTcTHJzul4FScapSN8mYtIhyqWU74HxuN0YsM/IsKzbNAiahLK
XeaxNSjr6vqp0p74UMTAe962r96EVe5a5hC9e8p9BH5Y2Hybf9KZk6gMz+/Q
wcdChAqTHn9+kwoQuQyGEQb43/IZG303LfZwHz1NNs0cEAADUcOXN0vUXASe
4ZMCMF7NYCJ3EXwStY+rIvIShllQ9i9DpP5lhIuZ1qteFuFb6fxhv4KYMT7I
/1uB8KTlHjKW1acXpW0OkCi615+T07sxnzuLiqCkY8k48ehfHf6cVbSO2OaW
1IbhZJB3HQw0iJkScIorbrIsU/sGg5EbpV0qozs3EKr7diXYHI6MHZfzUtbG
3WuRNpsPeqOYkxtiZyaBaA4xdcouSOAroZ2JZYhRUwMoUJ0ANbKZAr32UFNa
RUkH28DAszqqjwWGtZrEp3vaW3O/BmSEIg64xCTpnB4kVHH80J3/VzdL2Wk4
ggaDMzfQ09YGBzrPMABJpgpEM8ap98HKOvWOtcSwai/PBGWJ/rod+MAXWOuR
G/DD796LHjVGrwB1uJF9fXR13oeNj848pxhloVXaJuKBdN3y2sDzy2tvZLJ0
ZVdRvFp09OFu4TwgPZj5UsV/Dc5S85NH/Gowe1ijqNHmZcrKcq90qb7qU9/4
c0CE3Blj8UjDvZXaCAx1heEmrgBBy4W5BftqiI+F4xNFZurToJnlfbPxeUKy
Mca3dibDn7IT/x5PNFy0tTtygejvRQu/oFntQcDjrBeFa6loGf6JPvJQk42W
EIysCQxsf4T/EzNYVw1xoEVg92GqfhsiDVGoNq3tThajkwi9Txjko/d1wJ2Z
zi4GYZ8DCY0pZbpBnpvXQOIvM9mgG10QMCj5oXQKHefLBMyU3kgEbGPc1L5h
2Vj75mgf8DQ89fIDFz2vrm4VXjNfqpk2LIQc7B/iJHjTKhh5w0GeKFwlz2X4
LcsUK3t90EZKTuujW2WSsmlK4bcALigsrKTHo3XM/cqG+oDSUnU38UDB7tHb
0YJ4L6GGOjMhUovSQe/IUOOe0fANPom59ZT+NvqqRw/L/XbliqgshE3x3TQN
C6UsaKCvei8hSSaq69rD8S+OBG2i333CQPR32LOjhK/lmEdD5S89Swzk775Y
kNZtDwYu0NirDLB81GE1/S3OLMN2HQVAtLLAeY5g4G5kTY9gqLkRkyYSmssr
gDMkUBDHCv9//l1MgjdYmTm1K1rKdwJcjg9uASkCEsUFeqgAZ1C0FMJKqGn+
vqIGfFtV3YZuNfd+X4xyrjEgPoAoi1+A4J4BegLMnlhirIY5a/m2MzwwNYci
eJj59s5OpGbKGF4ZZmYuYvjxyU3+RxMfQyswdtTt+LYd9Z5jpoptL6gL2XiD
RzHehMhg9R6s5FK7WuztTOFUIj0iXrNPmrWgoCiFmeBjPqvZ4MshQrpvZLLy
DeM+KKyV1hIN8gvS2VW8w4QSBTs5tmF7B2mhl2pwnSbGp4PKrS5O0haBjO/k
FdXp9pnB350TOZ66SbTfnMkNEzLvW+h7wWMZ1Fm/uWYKj+NfwRprQvRdP1va
f6RP44Kyaorj4McucQ4+3ckfM5L8AU0CJzoMnTDzSXUQHQuy7HZNDwHktDmi
gzVSdweG8M3K6LngC7CS1sQC2IzJV6CRUJxIOwn+TYB9B3WkZ7/qO2jUwLGj
j0vYerw+9EKIrupaqljXdIBtFhpRcyo8z1qk0IBJV1t+1GFKQgxI49ux/Dhe
LIKqSgBGz756+lUu47N8ZOtAxLhDhcc2L3Kvq0xd51WEB/EM4eSVcQvkcYON
HzCWUXHGJInzewpNzlLkMqF7Mf4elak2QcnCscuBBN7RM+tS7FLguGF4/wdt
YKENoEZrS8u2vgBjxK5bzL0YNxoI9qZxAPwjIHPXz7Ym53T2Av57Vdc5tYDw
gbuvoIUWwJEZj1//LRZbrB570ggU5nURl0szm/QJtjOjYYkD+24XuyKjvL66
WoHoIBxK8SwahMuvJ8LQCRi9DqVPC6t/rGul8MOHFX0ujv9jToTmO6MaX2Mu
nkXEFOgEb4Nsih5A1Tj4JP/Tvj6TkA2l5tp8jbOMH3U1qI73nVM5Zc03lejD
w/hgZSTIbIXzCX/htO3CReL4dcbq2hjqjkGDhkAPrnsKIq5xZybuxuFu5VmW
8kLCk+9K9cPUZclx5If3kI2odofxJ4PTqUaYSaIKb6/tKuJou//kBr8LVNxK
0z4lVfXq0kE5WHQYSiSNV9KFK6O945MXCJDuHNxbrBZmFHaNNNnyBmaflAep
gb6NXuIpT9e9zcysHSC00TLA7dqFFfl6oVw50uWEiFAYCeB1Jl2jwsQNos0e
cMksdHn7iEojF96N6l8cgTpiyTn//7hZKdG1SJqpkp//PGAogGuiJ+QuowiQ
CEfmjBfShaEGq6WO6fHyHcL6qwkWij//7IZBUHoCj7qiualxC47iu5BWWth+
8J5w8BCc57rB0hP1C6fxpL3WlDhlHLoFcCx0U+vYMlNdHrcryowpozoX6SEe
6yfrT5BGgMCfZv0FY0CB6GhqOxSfPVoggk71tu2hNfdYzlUWEK3icjN95aEI
u4ysThd2HvAbmqxOw3cC3FhfKq/N1p+Ac4dmt/kiSMRu+kR99VSP+ocjhgxL
weLrbc9Kez0mnW2C4Ld5hi7TJa6h7AVRU3X2z8rXmuzUCUA/ZzXUPpaE0CgM
yTLMZltQSds5isIjeT1gvDh1/Rj/hR5trFKBklf7SGUp1Agqi0nIb/41CaGt
J/3TANM0KXSqmvklalpB3BjvQKbqaRAZTs+sTAn68WBnr4C9Ti1akfE603co
kB9VlJ5kbhalmY+X1DsPOO7oATpu9tdhQPj0JOd9ZfLKMPVU21iDAvaxzeoT
N++hpEniQSZYqVv5VRW3edAKc/o1XRAjyY/DNRI0okgHQdpuw1gHrjpQZi8/
qmrfxWTqWRFMrFxdHKZE7xyosM099vIefak4bdYzMoSxASRkqScIPFJqOLZB
MrVDaCeybJ8YTqOPBD9t+Z2tW1Iy+P7F3HnFLpMkaqvVnjln8LxTX6SPqYxi
ee+Sosy8FDaRCQPzahtTIPy8ajf8kier9TMUpBp439LJMYDFlslXPaaNAVcc
kb+5eQ0JnxTjZXXVHieKbftHOM4DRtMCvLLUori7TcrYezi1K+VZMOkUUud4
neYtRNwRoSrnbw7cp9w7FvVSlVaMcekWoOC7MH663skBa3ye3fuhXYr1G17E
zjz3ThwUhm3Dh2yQpE9f8IsmK869UBJidAqOg9EDXm44i1LbStxc4rHr1hAK
lZbrqLcvx1U3z3GGxUsBcausdBIpEAb/q46bWhqTFQbDafeEOpIL7Dc66BOl
YdYRixqExJ1hpHFcaNTHztOmMc09gujeXHlXVmO8G9PHxgO1ogM+rAbT0E93
5DUGqoV/+1SRvFRVY472AzboIjL1E2+Ct++AJIDGJBYsfYszHEcGSoF9pwAH
5ep7fryEinOJfw1Rfb5C+Rbi8aPFq95xhajNiMnmIPaZUkuzu/3EfaigcLhq
FoJn8lxa1i0ddUZwzraeU/8DFJxbzxEZ4Kz2iDhJt30ATsl4D0EEwFeGhXMO
k8FhxGQMIjPct6bRugYA71dvxiNPIx6wnMHDVZqvL8QSj2pLr5Z+z77kNQVV
p1AoSKqQZeDNfkbUcScc+4Q3WpSGjKIOyWgsnTS2aBskvYfnJghsCtaVZH6z
69QMDEJrwFcUhqVp5a4rGyZ8DFaA0XM2P5CktZCnB0r5qMZaGZD3Oog2ZxCj
6KDl54QiazLMhcfN3oZtdFP7lUPTvv4lzcRlf/rWm3MoUIJkxcX1H8qzUc+j
6ZmDeYaX89ZdPQVO4U8mkWZ6syYN4QRPOPIhgVsHsrRKVpMv/cVKjPg5W1H5
Cl0HpgdPWgmCOv+ooD5MlekUjoIdB9oWt6iuX0cPjLdW/bUoGy9Yq04xLJTo
ntI2IWcr5tLUEwfCIYV1AKkjwvGlOAIHQf2TiO6rTHSxh/OGBKwnXAnRFWhV
eKnpEYgitaYsoUm6FY6jCHTIOBxq49jywaK1GcwAyCLdIyjoST1WG+N2Ms+E
1bCHLoEKSamKZX26EIYwwfeKxPXAUKWf+RRWbj5m5PARUdZRYqL/8ocxF9K7
PL1S16T1OnGwQFNRh/5cHfIy3la4SkZ2+sGvT84/KVF0xDeAoD1JWoB6pQDq
uQTxJgl/ANvLIn72tdaKX+a52sPUyvQ4kfvx+dLSjQgOKfDtf+nlwwMJCY55
RuVeKgfIWmFp3xzSbHEE/tqPh5tfyWlENfGQaT166IFMcUytMiRdONpNipX1
s7JDadv5TMePikLF6Uj6zioKnMIHbYKzZivPooCileRpdfIGi2Tpy0N9/v8o
nG7gEwogCFzOybhUyivG56BtMu/hYXN0qKTHrDfCJ6iJOZmGsJHlJVW2DmoE
s7jpY79rlM7r2dPTCSUeb567BNTpGsWbCUS/bFFaNmVQmZQDhYSS556D8wd+
2qbZTfEtWA0N04UsBRMSrqhs6ivUX2VhyCG1BDm/7uIM0o8dw0wmrARNmwo1
3fZROPVdKiQBIy53CaG4H+sg8wePIlUGnOV6ICLSFZe5TvImY8WcEjrF/usE
8ZFtoPgfrHy3I6qo73SN5nsmqSFCPGBzgsGe4bu9JW1VqDES6KcrGrd64hMd
1QrWbBEB2LbuZMNuNRkeOBnUXNMqoGLhBkRD4UgUBZqSLdJ+AKvWu4NKjcIT
ulQmoMmwQKKwtUfBll2aVOg11z62WLMTUOmKGjQsBmtuOpXaGkHEYSkqutMh
++gJR33yMo25jQncvdMb7YDSOduP5fFX+A4ECu6hrR5OYQIABE7Vm0rXHq9K
UFsDxEx7Ktzujo91TbdUEJm5HUpTAoLFFr1hWWVKpDAiimkLlhRYmJNGRsnl
G5EunF1UWytrjH+2J0TtjPGYu+LCqcdGWGbP1qr0/gyD/0T8xOU5611+9yu4
db/Mj1MX52AXhCw7CpVNH5YjvQJAG2gGxE9oPnAih8FJnwo1583+rQEQoVGy
PpWvzk9lKr85A+SltWOjkWvf8rTDcKoYRpx886QmMG83sbFRmG2uaBK42HNm
xlbs2x2Y5zrAmn1J/wP/gKGN9ZdDb8TWQEBMC2LC+IW3BBfYZVOV5i59pZjO
m8E1JFwu4yUuE4lJvM2mcaQP/D+5pv7P+KYU3PvAiwSaxBivN4UMMVTyj6VL
sSTSATMLhrsi8dg+LVXiljhjZmMjWzBCFHR02IhJDBJOAOM1AfLMx2knZWdW
cHK8ndYjL9TGqJ1+JgRp7NdSfw0KIyVmrYRv7NfqlPC6y2WANjM7rB7HD9Dc
qVj6Tbl0IAihRb72KGQ2ERtd4Rehf4OWWVSaKWPNVsLTG31XfSYZNwLLnmM3
pspW39q34NkYu8ifInD2+RDJLdv7ZEarYeZJoPj+NDzu/OW66yMlgHsk+1J7
iXLNBAymJbdSrflrk2FKO8MX85OAZZaCI3De/JOTR83zYwrn001Aha41oG7c
jfDS0g/f8vAVOVIGc9sOJECdSdNuZf2+KuGG4AGdqifkIhl1Jgp15IK81s/M
LgA480MDUgtzpi3rMdp38NZSU3V47tWvo7HllmgcBscQUcFj9CesDvZzAV0p
MQM+AdpZBfMv9rfzgIWLkGMx8nYkHDE5kq1xVAxrOuKb8lDNi9Q7Dp4NnpS/
SncEwzM/K7sw3IAWHW1rAqsMwRpia4YTRjmeV4lfw1hXGwAlOzkoXxAH3vwz
8f3rV4ipkJFxtLU3dn1nkAqgnfXVCtpB55ttqdbyG5mJB2Gki+aeb2rnKNi7
OzoKzeye1lksibHKsvyGpo1hqH6nJhLmArnaveSakc2ON+RAQH/vSICmOTWk
I12xP6bZOs0VUgshOX3B3HZjCEn+ZRSH027RCRV1bKTbppZeK7emwtLu5SXs
/YfizH3po3ES8akyuh5DLV1MCP4Qszy4CgpJWplBYQdZFQQolpkJGqNWXnmw
x/CCVays8qc/JOL4f++rEZdHXUaCzdNogAIzHKkLcEMhS8zQ6/yTsFt5C8ET
AvH/b8kOQQ5P755LLzCIPhFrKzqmHezPYyP8bMYr5XatGWgKKt1vwUFgDPJl
oc0cuS9DtJ6RCuwt+X/ugAoXOOwHOnuiksl/P0z94lKfysvMORXoCPSb0Wt7
LAkhXLmb1OnB29Vj7uK0YN72ZfLu3Qj4H8roeJFpS6xIjDMFn3bHPHZ/9l3g
IdX5XWxx0dS6X4jVkevBdfIV+8fAs9LPGGuh1l6drSFPk4QMAC58DQJkfsHf
4GfzLlNciEvRHCvtss17ftfC4SEa+ol7w5aMsgSCRaV0eYJsegtT1VXkVxTD
jpdk5L/FUKpLhXapsmDKM7Ai1QMJDY2A+rvfDAdd4Msq58fS1xE/4ghp6h6Q
QZ5Z1/q70Omg6BDDJpbOY+6zMEvdERGrpTKCIoAxsO7cAjLkvlwmK8Wm8+vW
jyFPxUxGlAnHOWtuN9P6wZ0ZgC5CKEhSk7IGdLUeszt7pg3Q/7SMyBxX0jRb
bRhEW1/XmOUbwCsj5T4e2ZlizOvXkF0SOUYIS2e/jE4vwOOehgrnbvf3oc1u
8NW9UUFV1VjeE3BovkveMacZYZPU5mwXJ2tLothdbsLO+HUtzvvudFTl0Wwr
smh0f+eFTixegq/c5CVUGCY/h1QhNe6/79SUkKdU3/x13jRAj4IUgdXkbkqI
BI9ghaGijqrHL5bApppvWXacXataVx159y7gBdZo5TJBEclxUGEZCpT3OE42
dHO/jrsqPHRmDU4H4bsVbBkjcJKPgLoC8K92thgADzucFqcP/DOGPSUD2h4C
uwNCCsxlcXxlospgKtngJNh6tN7UbftB2bOTqhZFjbpq0jTPCnMs8afKTrbn
FD225JWzYYm3coglnTxbMXAIw1BeouS1rlKF9OW7uSonrEAhrfhoe/91/GIq
Vhe8BfoUpUnBq2zryCY8MgdcBABCKXnU/Ygr6P7JDytWZVgBCpnaiYzqzBX4
osbeYgI0RxuDQ3di8zcI7p+Qi5YMCzF5wqZlj+I1nRo1GrJKT0QhU7pOMsma
vBgyCJ/nmXF4hDKKH/0gJKODK6SiKh7SkfPopmlZB3ybjaioROvCJZ6/dhQI
wG8abwApRopOGy2/Z3w28T+OooN6ieZ0BuhJlLmjZ5e5rQULc1ml0zbvcgCB
Epxz4zXSyn91rJ12Zbk15NA3mbSdMQKYsrAHjFcycIl9QZ8JiLyA3z5IHmXx
LJRYvs78HqBYJ5ZN+svohyV/I3sVBalmgG0d9oR1IwVlbzN22lJZnriEyAbe
cE5NpIVeq7aqQBkapmTeEldIwlyUP107mp+zh8EsD7cbIC3n/vQs415+XcUv
93hBXn5CvBQl1UJvF23za5oDg/hVV9eubsB1Y9gH9dV/rBEwOuPyxJ24JXob
OtVF/J5d6jrDTUiejO3a7BF/c52Z7u61y4CK/PasxT8SnXnEOJVDq9b8SZ0U
HqVPtvWqwAGv+SJ7Hx+nPw+LoEWcdqY0HGI5QzjJ8yiPd10Ohe1jmrXGS4Lu
clAfwrW1Yr3qPDix5dmZ/7BU22mEXHFPGpLsQkLiZWY2T4MRF1wOODbzPjPw
x7QvEObZDK9Qzr7dXpWtFR85UY6XS9r8S36wKy7Be7A5CQGo3LoDxxth302y
e94dqFhGFv7LK36cZAunrdJA85I6QvWI/hx53dbvtjQ5CpJfRQUpPpzpMgvs
je111Oiio6UtnbkT4c+5OcnpJx7lhlYYhLeAFM82uTFmvWW4huY0ku2qnxXG
yF2Kbzpnr7H4+9CvnnnQ+szUciEZCkxIgDe7mqlN95vx778KGdcPYMDpo5BQ
ridsVRN0xwfVwOC82O1h1jCP3a1Bjyk5Esu4tay6TSsF6PoTn+BbxtXldDcQ
4kVrJz+XQQQLE4JiCwNLx4jYQ56BQu3jQZa9cUtHy+GkZeLQLMhl1H8bwoLc
oFgB1fIZablRRhVSVpIz8zqtiK7OyvshDoaPB98K5bYcSHMORYBY7dc/1g6V
wkZ31UZz224sKSTceKoJ91qhR+gctkhh9XQQp5A4n7ejXLQWqt8WGJbd0BO+
5TvfwDkE0vcaMZUIPhpCMXU4MMIlWBArZR2ClgfovdCPpWdQ/FpolhGFATh5
zIMiAyHLZVpjgJ2Dg9VbSqTfMjmYthPZSNMhMvkeXkBMkZxCj/hlm084cG6x
8veeEKLhDQPyiin++2KAAt5U17u0v+mUvw5Pk71yBgm0gaDexI1lVY+j2NW/
a/EzhoEimU5mPaZkB02LxobNZVtxIDsV0wdFVx7IIsEN8VmqaYTyR5gGQuZw
jR+fhjth5tbYcnUh0mqGi9/o/BO13MLN5p062pJQlbfiVwVl3gVTuaFjidjh
D3fGICvE3uRM/WFZQundBYu3PJEUe3GobHap+xKF6YfruB7XYqbTJz4CqVXp
8QYZef5qbsmXy5JAt7LsuLRvfH43m3qLztaTNPsplhQNY07AyEABlP26QtAc
lAl3TOoTa5GkwE7rZg+RY6DujE72KIndUVL8HaWpQULIKWyIm18uVfZdSYjF
mDHT00g7bilY3AU6L85y7zpFyc7tLKvkJ5Krfv5hwXGiIbTnSrYkGfR8xJyh
Y2wC7JzoVGQJuU5uoC1vT/4vKFK+1BdETTSwivfg3qwzcSSxvJJDoCexCPLl
5ifZbChd2cUgjW/AWBAdnm9cBjb+0OAG235bHCRN/nWjIrkpQHAn/klO874R
iwGRftTFMxVBeTvrxrqCoJX7prfceQhMb+qRLM5W6QKgxm3kDKazjJ1eScsI
7KT0fqIgdkzivrqDlzS5kAQS/+D/tYfw95EzLUwCXscBKEra/toZ0ZiPbhH5
QwZ+sFnFrHeMkJNmm8ind51GP2FDoZ+PhVNCpVSX5wCwBbEbLLmQsuUOaWUQ
9y90/zYjjfWjWv4elvAUrPmpbpDKz3eBCueWgDjVIm05l7CNr/xk5xkpMpjl
9JWYSrTXKzH/mFrd64RTYr9lRIj4EHyuHB5klp1S3JhLm/S7NmKAg7cEmV5Z
+k2vP6+ZTbP11ganjw2V3RFjPHjFeD2w4bIGAaUJZPhPM5Z6N3giweIgeBiC
JDQ/4KI7RPgjTYWXR6OsLGCdt5NQR5GvOLPeK/lFhq04As/I7UdbVWscBghf
pF4PhTsL8zkPj0EJYnnP1FsoXgGSwccieua2cXSps+pT60OMSxv5km9C8IPB
yzSvIA/fMpY9ktjbtmt0uKFlX9tNtMLwmJtyZo5TmKv7e/LAXQ0Z+K35LA3i
+kEszZXWRxAmhwTPGzZBUTeGysJyh9ahWrMX5dwh78t5yiM+cvaCB3sodvb5
N0xAgXoLhqZSrtCZhY8vb3wu7szrPbgyj3ECzavndB49JRCrmnj5e9ZwxmYy
aM0/0g//LMf4QivMBZAmZporwikTnvuv7/O4OKT9MCu7pWCn9kYDTkHz6jH1
iBjT/ON9l34jV3VndT+CPdI+VXak9trb0V5dYI5A3tiQBkRYkcvr1amkxqCe
5gN+My/OFdD64m7JPx80ZroJ7f05+t2nEMXeP0K7g2apMjVO3Y2LM4LGSk+y
kJ3AO7w/i+YWJPEewCbg3n101EqRpGFkyjqzdsYeI/RKc1SX91wNaEYyw21h
Pe7WBcG1OjXmFyP4up198cO/CfO3mJDv2k3/eiTpiHbu/4tirYX+nvYXuoki
4mkBvWHGG88cl9IUmklWq9xIpBdV9fixmVRpmRsgTgeFuakpVzucR7vIb0aF
UDzL9xuCOgwIXjiKohXwe+y67EEYsClgSkt0VyAL9JxCjuYrU1Dze4vNVqCw
0ZmXJx9WhsqSBGW3KKtcYnB0EX0MABBBjumGI0VKYNO/etLYnwO5/6TMLcVJ
byfZdGKony0LEKl+0ZnmqVsVwcb91sMwD9bCDsqPWhU85/XV3WDXUKBz89s5
EsPlwVSpEvh5x09rQfq0nBQXcSNGse0OHaMuHUOCkz9Wt43hNRi9MrGjHqEK
jCYrCq8KBSMq6yF8BmQcY4Gc0H6ca2rbzy++7Iw1rWvm39DIt6BfRSvAKbbH
uzGDntKvt6sPiQQDJYd237QC/Yo9pzvrSv9/zcu+x8FDj7KwA6a6NpyRuXIw
YknwV3cr1EMjxG9YSFWSfC0kbQ9hpC1zFvpMqwn9mDJwub21FBV7gEvjhEcZ
UEoFXqyBgRX9vnxUFVF1nuzXbkceQMRlFXbEo/MJLahvefSB7ExFzXXccwqk
h6c3SLLxs2hRhitnf+2KUZVpFW/wwn46ynPGZ/IxqusHC32gqRotqbvCNVum
E9+V8ZiR0HEv10z8IT/U9Fq2wi2+xCTL6ae2IBBStTWQQUUjPR1HEa3G3vt1
9OuG+gge9eCnC2U0JMxoLOnM87/FTBfQRvq37Ecrx+Ry8CnI+d3eQEeV9Uo4
slCZmyuo8I9swWEVK3QBGQndszNEKmvvEgzjPb4mC7vB1ExVVGZ2OzKnZx2l
eHp4wODjJMR154uHDnF/zgrND2Ma2jm8xyzhGlFm8UxN9+YTxg0w18XWt9AK
uBhxkv9khDXV5zhxcwb3hgojZbr8DwiEUydDcQ6YtEijfgMyeQSb9NRrMtwB
L3zLC417081p8VEux4HTvCAIbS2GR26eJ/F+IGZpYp1SyecFsbN/nI3UEDmt
c9hmp5wV5Vrrlz/yl75gyR/xiFDylIx0m4p0K8jElxW20UvaBzD1yfWj0DP+
Fh73fti7CJBMJWm3FZY2EacXq/PpqOlpgEkeu+TfzkVDmSBL8+pzMejS+Zdn
uGjjRXBZyt1nqK8YZ3JMT/nWegRehoLL5kVArxXwS8rcikd9/Xb4Apk3NYad
D+kfHzS4jSzBCNRPzKW+jLpci2xushZuQaYeGsqHs98lZ/AtXKPNcLOS+e+L
bqqb8/IVtZ8maDpf0y1X+pY5zmFw1oDoL3LirlYGf1Qzz3fP3ooCufkN3KtY
fskJvbYYX5KHRwTxdAopn+dJbmbd1EjMzbeUSB8P41ic6z9kszGTBSIVD87r
gjRYH2muGERvqj5lEPCXMQJuSgOuT1r6v20PZ6woDSgsGwPJRa4EM6y/VOk8
4uH+4oWMkyaeiMKpdn8E1+NXwx97x34ksRUz0wZCs8195ksrshSUD/IRPk6P
GNNkHefYaieRldpO5vNxSR7LKkNZwKEOxZzHu14p2RZ6XhpmsT+FyjI0yMqp
LBik7rvuba7KvGi6ruHAPcM7WdzLrfwRWq8U2PqpT2F1BoBTpH7ws1jd27AL
erpua2LAHwQK4Viwdn6mB5C3BLLLQZxyUPkRGbshDWGPAcZG+Js2YTpmcoug
E7WUE8Ns7CCjVmTucFbmbVEHrF0a8mJSTE1KJUlRldY0dalCoMlC2ZmiG8wW
tgjcVbk/LCkszBThZc7HGT0fL6blbiw4sUXTB+GwaDNtmRyTiVFwbfApxOul
i/tDdZj7RMSH4oAANgIIA+yevLizdzY9QfvVqImTKTVLmznMssUXWR+1pArI
k11dFsK0WJXnjawMdEMhn7BFliZwu5RrBYaMQ5lwx5+HdcxxAIQ6mBXkVQxj
PBC9HzFN0FtCLpSdufLyUf5MA0GngBtEMFkNLty90Qs+pm61A7DJx/Lxfm0a
5EXDuMx6teeiZpmIsD2N4eF5N4F0HajLmY74ETythjmwjfmEceSKIcxO0iwF
3KmH7RP35tq+IlryYfYTEjTXai+DKjIPTWvhCskGXfzgoGDdubT+VMTGvAtg
rjsHAKbAqxWbWupWLtqLp51ycTc5iBa5WV1TwzLnRkMk65VnqiGWNSckldos
xffkAMksrqvqv0FK1YO3Fwf5E+AVknxFw6eR36R5tcyEQxmJwd+izZgsC5vw
25Alw/zp0R5a93hXj+OF3HEB6teAMpGMfWabrS3DlOci9H9AHzzUJQwz2WaP
OYgfbuQPW1mNfmvNcqnSYgE5+rwQon8Qu8yoBC2A2pzDL02gAJYTliQA2q2f
E8lXF4NACodgRz3H4wpH5U8s5cg/5heSzMNnhyKyGVIF+q1eKXEv2k8S2u8F
vs0tRlXRu8TAfIu3p0BkkAILsCpFR8Hy4+KqHnRIB9rWxsvx11A95RBCblCp
8zoS+qyVp0a+yd3RMOwP3iBJxQkE6EwiVIoTRfccvXS90S8mYQ9ISeuFsuH3
xG/kvUvwlJoA0nmdg06YUoDPpu3R0im0bnGxGJcVfRCawFD24jVQ3vGF+L92
Fqf8dYEykNCVUWIMmCdpfEKlqS+g60TnpBtxfayel9Mhu24YyM24qypwsJ69
3zDIZATxK1aqVg+lBjIWGUETWh/ppOY0IOEZaDj2oPDbMmEJT657Jko85UuJ
EpelripwdIS4Crxc8M06wDD/qdFAthYEjWgdT/ktC0gt6lKqXqVwojCxIioq
AkvLEuxEW9ZVCPjY5HWSgcyKsKDF3GK/1kTOBFwUzYyl7SE85/pb/smluQ83
WhTVx8quvhWYf0pBIP0MjUtUOPFeoX17cJQZBQzNlov5hfh1sZ3UD2tucmTp
w7XPBw1arUC7fV/n4EGT6qPDBA9yCIficELtncOBy1MIMdbbXHdZI0F7wPSc
7RYUH5Tdr8IE82PqTPXYJiyhJXITyXtLaeuB2R/vGshfzTIt+nvx1/8uqOzZ
Ld4obWH4b3f9jhR3Ql3h0M497xZpaWJqQHs712zboj0xlJA1pF3rZanbh3bn
JZWhpPBGmq3o4e4lk0uGLaQG3gJ5Z7f/CIwIM7tQBMv2tZijKu112IebNdfR
/huozI8lUVW0pvLWckmjwoYGLpHUn/KFiInnJOWXMKXUE4jdorOoc5WhXRxe
R2PD0r4c+kkrEfipyVAA7nDseRGqHeON87pwNGbLprQkPBYJv0P7UVaAQA2l
8Fx7Ey7cgz1D3Y+bVWvlrFdFiIVvGXPeLfoKYN7he49u8qJSjZje72P3XQwx
WJz7TCxkdUCneFPtddA/uE2nerNOKmjme+hzUB1V/t9qyGavcqXMwLYFq7Ut
BQcwUv5ZbFH4UbMdcI3saBUvI+3PWYybFBvCRzXFGAAvgG34NMWIKd+wnZlI
l+9xKNE2Rn1uosBKR8ijisjMjqvloAWXD7Jh9G8Auq5gYiQhyTsngqEsfrni
mbHpA18LWgGHxp0oFiJKli5SsddYgvtGzwSTZ8TSpQzIcqd4uEDMQ+NyFBoD
kOmn9Tr80e5x55QYaCMU3cUSXHIHOEvXXezdsnksG4oby4/0HTsstG/SGo1b
nuhO/mJFOacF7GpmTxEM0QNg3xdvFwp5EypycUnAvWhy6fvNXvXo1gi7EaYx
J0+5rvl4kBE8gnLkI26KTScfvCUl9nhWKF27roZpxzwMi7xOMLU36PFvCQZp
9XjdVh5X3wYCKur/cCY4B5nFrIlWJXJwgI9pTcRu5R5z0sJHI+TrYPUYVLkW
oA0IrBQB6dtkPuOddTWWNb1OpiKx7EQf6fWbda5g5B+LBHw9AyKqjSYujM1a
3B93H7c7jdzCmsydpd8wdEERdmt/hvQ9R/RF9Zpp4Re9o/4lhBJtknGmEIo8
18aiYSPV+/BhroUODhfWkdu9xaABWthJhDpEUxGFWV6CxvljXxCuyWfrQZPc
59tDNmO3cEujBQ1rYD8mejC6eftH4njjRFq+kE9i+ep/m3lanMbmyjlsFxmJ
aunl++//u4SI2wI1M4H3GFBwlSDo8nkAsySQ1DlU7V61NvxJebfavmisqO/n
nK+vOKAwFdvq61C/xMWVlLSwssfik9/KKl0JaGfnVUUlFyMR+lR1dfhtpg6j
yYlg5f0OcKCwMEukQAi7+OhZ9t2Nbmzsr82LsIp6vH9cwJi7BclAV0Nk3rI/
DWy+uT8SeGCDzB2FP6qwFQUYFcB793W9c6pwi4Jg5UGJF+yZ4UEmudO+XqvP
NNtaxMSSJdxvfWVVGkjSyokrcMYIkSDLJBAlawda1NVnN/j7p2phBkeaWc9P
is93BBHv/S9eLghlGau/XuUCt5UCjStwujxA0tEWXkJxIjwElPPbuXMhW/x1
yC8tMcIiutCCcPYnNua8VD9mgZwhbN11WU2az5ePnrPTcbOf9OKQPetUUBIT
79D1GUTUtlWn2MYy97z/cLNwTbu+scA4C2dvqf84YJZCiTL053BhITNVWQfi
yjr1hr/A/v4xtO/CeWPHeH0E5Hiilj/QlRjdp4CFsev6RwcAOH8gNICHG2mP
0vUfowDKdRc9qwSykRCucUkUp2BVOD4pqSBU1VXtk2eBhmCW2LERE4ITr5sZ
QhcuW+ik1vqs1zSbq5D5pAcwVomV9ovdkFm3+W3gME+jzz97oyg3/Ey4ncBU
F5i1Hz57D0V+fbN389R5zvPhsYLNkr095b+9wuCg/tcu/5P2rQQOU50iiYgX
ON+qKE5FDCXAK7AnXcRQnyTrdF4Loe1U9gFdXmp60H6TK8NIZh4oIwYD1y5J
TzkY3rdG9Ohusau6qIa9l0IGdamI7lQrh7uATb5oXzynTAzyypqyQX50Tcn3
abwvQtZ9dPdVo3jpFjG4dRV+Y2WDdV38uJ0DM5Gjar6qa8lAT8WaiAhz/rod
nj0BIihgmO8CIwM9aJXYlw10MynEFPogZt+GJFJwfIDIfKJ4JGuRfWBDdNn6
sieH/aiDiyzLUkaE0saECETI4WSlIdnp5q22bZzek4yj/WhcTapjy8NLeVaS
HbLiF+xX5xxWZPZuMBzfSce+vDoXAjDauDBl7BqEuSqy0FZC8o1tGcEHmf+l
9kl5AXYA8r3ghKZQQp5yQsRTH5Y3DJfR1UTfHYHmx+WHMnQaqYI+JcN2OQ8R
sUi8v5TNa7XfTzXGUou+45LOr6H8C1O5/VyQ9kR+3c7ShEJQxFXjJUX0tw7r
LLqCKcbUu2fCDKnbBzeFBuAF1uEmYgJ78aya71sSqoUVbBNTG2PXcptkW1NV
r3Rp02BlvKhqgildFHAWPiKZ5MMvCYOyqu64kpqt/jNaTWNXr6M3awK4hXnM
xIIihJHnZXKhUs1cwV9pQHdPNPID1o5lIBVDBmHJaaYFSLp+sheNZtMqW1Ex
vDV3TCcnxpnUfMWae16AHjQf96e19WMFXH3kl/0pzND4MUjclV1ff/HXCVC7
lGKHv/5qXCdyQ7Dqslhjn7MctGKRAe62IG3EbMUZ+JI9ReC9KgV0x0kw+QZW
vQxeBunlqLH9LNb9MRJ4hGkwaCWALdo0c0g9or4/EwR26Ovl+FF+QVmcbviv
WkgN4Bd7mL5wW7/KV/RgoGP/eJs1glYk89X8oZVZnVBMprVBHRqWLp7YIVC3
GMXV1JSElIBxcW3UcpBWcp1rThnKjYCIYhHa6yFiS9xXzfsm6xdHN4FzdnK2
Mw2oyQi09W+KxMirlLXuUZZSDwgFCfpxkmQUc1v3KMHQY7/+5WgYqw5fjszH
w3eiZ9jufwaUGbIoYgYGs6sxyob7fFPMhGN3kQcHx4UFtXV3f5bJKXb0nq8t
85gXDLdyU7kNO5/ae7xBEOOxlH4r4cgIPFwV7OfkX+9190dvMyL42HJDkBSU
RqkKkBia2DU+IAUbReQRB66q4DXvma558NjDC6iqlCptCSXHfyPjOA4Cu4Ba
ND9LZXClC2OfW77JfWpyDVadjLjWX9BI4HdmUskeUGHJEv4ElBJwinvcj5un
fjMDVjnargEk2+qQGMKmBkxfBPXD02YMAlnEAo8vg3iGU9SRlvIoLK+t0qG3
1PGcKOxFbCO8xyPlji61oVSX+A7NCW2SH0ZeT3ZHX5v6BEL4umKh6L1n0Akd
zI4Y5hGOGewKqPcXDHB53b7MNt/25bO0vCR2E9LXZzeytrVywBd5EfD9/Rlr
LMJQTyZ9EwX9FkVZX9v/prtXnz85dcMxn7eLUvEelErZplA6cbrqKfniFr7N
nqEw2EfUhFrASNaL22xb5whf43GsZHx/L9HbUrMntp6/EiZhSKqo7iVliT3U
/4OXIIyN8wg3U3vtivQOikW+OoNOMaK4r8TDCDRJB9WLrNwUHyQizx0YH6Dr
iDce/k+DI8S2OyQUzziEydf47FK4e3/5Bj/RvDzzuHrC7JMa6ZkwjrEeyCs8
bxEDAdqzYP556OTzxPoNzxFiLnX1QdBV6HYX28xeCc9PwG3du+8zsd91zop1
8bjyTfFLD0jLaXDQJ4YDMf8WP47kfMMx7z6+XdsmVdF7zzx8S+BEwooyZB5X
n6W1nk+wHgEF70yOiHxkWqa/5ZiE+fjex+IhPlg6VqOsAQdGK0nNDAzO1nWT
IMeR8mUC661eAJYX+KlWFdplVJdG1miLwRO8Oox//LaBoMmkoatPlbNIArXH
taJgGvfPJTrBnIXGpJoJqZ5gIABOiU2FGEYMvUtPVQvcs03KgnDVirfVUNm0
AxMakOiZmVYhwv0g+vocrp0uwylAbdzAYE7EW+GMoGIWsfRz3PDmnMb8qTOL
+BaCjZByAZ/YHZVLEwjqh4hgTqCTaOFqH317pnZ4+dEBX2oJTi/Y00EDyV4p
+pLODDaz9a8Hhe0eijxQApD90pVwc6vjFxuGiiDqW9I+wled6HnLyiTmD3jD
1elm5XCaEwXR4Uc+Y4WKRolDDfFJlLu9XTN8+rGE2StGEQj/1PLld1ojV2hj
VUOjHsesCqn9KkM+Xi+v++yQconbxm6Ff2cPi/olZc6i5nTVBgF/Q+Emseni
6IPnTW7ANf3occvTGLzlMizrO1FFf9BCmyIwkIWZHjzT7aZBFGa/h2QDSvGm
v9TFs8ikkH5E/ohhBUX7yaP3vU0RJz/e4/pxcDgqa353/DFls25+PyAcDHA0
1gd+8iuhVFWfccOdiXLLl/Tdbo9yQ4NOxn74EARIQ3za9ixqyfLFG6NHZG54
2fzOPUAbOpIf+FupNvluFdTYoVZiquNxF/wpuyaMvuu29ZfyEKq76Rv5Hhri
vCX3iQVPWOVPfdZFoy8R3OG4Bu8MKMorvaygv1syxSG9wENrq3rOBu7WrFXR
LPVdMcQuuYarzbqX5+bUmriiZR40lditV1syf53UYAc5EitDphWS4CbX/bgQ
6E+K+cTyOQRE/Yot2d0xy6XaP3UMnj2kxiRGsL882n5jxczEfJzYCHLY5kHU
2WaKikmOsLm97xJw3hRhgpaQlc/atJmVMqR+Xx9V0p7UlQ19l5vY6lLjDoAq
f8bC6gZyx3uIvUF+7oSeWLSqgOO/ES6ZX3HjgfRkoZ/upF1XWbCB4NdgWQI+
KqBtejSr6YcTECauZzzoyuzpTlv7DPKvNZCg0ejLts0zogOJtaXEPnlCNAim
MD+tytEOdReSo0dkJdJymmh1aN8urFyyNwU6mxQm4rrXA1nAxgrKcKxePXlp
SVskvypDFaQD2tRlmFO1E1y3gthCpDb6W8ZdnAfZ7OiITzvmMES7hxgGjjUl
7V1odKDIuz8rzxIO/3wsGnFTaTRZkXfDnDkt53OPGPEYzW71FA90p1tZau7f
G1JklqsFlWkrGdlLqLwA4mLpoghd9lD7Px9Xjrr+b7hNYlW6ETqIWne/FB/T
QGYmlHXdk4MmAde7ingb0jMOrJPix+wyPON1ayAbehpOzYJG2mHdu/7NPFwR
Nnn3jBGzWALmGATM2Nofbj4bSsLfb30g7Eml+SeblJ3QBuKL1rbJW8PO8zmj
YZoXA0L07pQ6pdlHgsAW0zIX3Mtz9jBEUIrBR5hXHEf97zJI4nlNus7rGLFx
pEDJUW9x2GJd81vcqRzufWvcSlOGcuxqbo7JuaduQTkCYt0GtIfkG4DLT2/R
hygwTfFHpzKLWIA0XEHblCPXV+Ok9qc+Gh/FYHvrVc02sLj6PDjFYnZcEGH3
dCXDE7qOiM9TMfypQXzjYsAUEg1bib3mQT1R+t2rz3Y2phjj6F6Xg+V9hZoa
YY5O/ITGxjJ7A2kFQAhVyps4EYirPdnM+O3x+b2UsNAmfpdM5aC9Tsj3UlsZ
g94/xurCP2Zh0aHut3cjsukE2NWFQgZJYuVAzxIGlKVC0UJxmsEAryxjQO/o
3L1IlBMAlLHaiYgPRG/oIO1prQ+RNzeFiRDNhOHldbg5T4u3V/USadcPnGzh
72rCurmkf1yHu+trqPeHuJwTmbdilcF3gbtw+PZ5DeWC77KFTTw+KnWqn2Zz
0Bxs00GkR0DH3oq8dsano1vgYgoZCKaszrJpYt+bdqOyxp9wXuaRpG1DYdYG
l6Xk58ZMBPyx3qeLTFhiz78htkh7Sn45FLC2rI0dXrMnNxM1C2D9fVrjF7HM
t22idZsoOyf3PduesFfpeM7GCQyAgXNpxZV2qbJFOohS/G9cSIjuy9ebidrI
AK+FUDHB49UKMRDK/PpDhaYomafAFlc+6IrlFEC9JOZz2zCgXx3pd21qStHA
XgGJD/dj6otFNkv1pLq5IX99PJt1W2UzpY+hYl3B8G3E8XC/lZg/qa4T+sM4
VkPxRlifmQYKtHn2HkHsDtgpqUgf7F2FHWMd40WUqrt4Xtey7ql7Vv/YlTaG
nRx/YXX6IP35HwyA8JLUIEmVCFnxE6N354NvNFtd1GAfg4KLQcxkQpms6U1h
ij5Jo05HP34ORsmlx9pBxMJgqA9NzBf2A1kz80YAzTaIDK/UUZ8iun1N1rcP
WEP4fvKRCN1Tr0kuIRJbpb6Cwh8xG68LstgfcN5U0FAnF3aOGQo7bw8qpZUW
g5QRfw3RWSow/SNPj47DLj9v0fVyyBJYfxAmOki1IwZsYndHc1JkM7OUpsbw
eYwAiCCpWGRfVM2CqueNsq8FNFwwpQu5O86J8mpA/nxc2DHE/E/KeDhJ7w72
PoWss1BRDjyW0lclhTxExWrjmwIC3xG2gBMsyxCiCdz0AA9Zzr/RqAopmPBW
ML7NnsiwYf1ATjPfOGERmW8tf+1XnYwdHXEFrs/EyGNple42K7xAb8QU9y0e
u9s+16AMSlEve8mDoP8FGympOd2g0CXiKtbfYbJ9NEMqBWVA3zhXCRMUHoW9
likizvkLwlvzLp/MOzty7WAK6WaWBiW6KQ5P37HRoFHJ6Pni35njCzT1cgCi
BeLTnl+eQFwuOBm7wOHlEGLhbhGb4r46sHW5tydR5zjN6VtD2E13uQrgtbhL
1skzAvZVPYggmjvz6HrqJTr1FdYLECJPmmNsbicuGcCbLKpbdn/QwViWgRT0
lnxyqr94oZ62u1m2/8IoeKqPxCcrQ5czBLtkfleJ+jmkdOoEFgGltrcoEzmv
14yZA923DNH5svo3HItzfp93QxVord1iq+nqp8dgzfQ7o4vDBjLFW9EfjFQE
60UOHIhi6SIsMTO7CXIhXb6tuTVZG4DAGikFbFqSzcO0Rf5T1ga+TbNDTWih
HGuSeVQ8hYogOQlNI8Jp0m2YQX7CebBeOq7OHg/VPOlOjXbH1op81EUf7XQd
g5vwfUfVtx5/zxLmPWA0BnLeM9kmBrM0cwwfHuWQtQ2l8UVWDfBkyBuNosg/
NYLNnDMxa54PIYia/LZVro/FVPwkMLgia+6lY9R+frYOg1uHJEgx3yVXWWSI
xrw6F+eas9QOZ/QxsOA2m3IKnGuFBRVveUDFmSZLnzups36cP8/wkE8uiUVL
TEIRJw/nSWZF6YlaXlNhBkiX60aiHRXAypTuCcs6O//dDzBWi5OxthzLcHAT
pSgZdksSL9dWbXl5xm3turcv73LxQvD6JI3/p2B7wJXvUe7vZQuk4MEssBEJ
ZQnj2APa/kjPYWcELF5gZEY+jE+ERJLHZvTnwho+zyR2INtTzgEVSJ3vNi6N
QzCdcCDaL9rnhQ7xmxuWXGd+Y/BlgwPG6mzvm8G/D+4ag8Z9ha+YRzjFySCX
uKjEaoS6bLNY5C4D7Wi2ZqThxWft/uCQq7YXmDT2gtVT3I0ijJMtwxoqajqs
MZyf5ODO7mFlM+pnGX4q1i73e4jazfe4F30i3Z2iGbs6xd4wSXeeQXDTb4eJ
whF+G6GXNKbbl90IkU6zKq/U0+mLZtLSCayDxR7R+0D89wsdwggSr2qorVj9
eLVEuotAxNCC0WmwRtSRsTgQQRB5xY5PaeDml02KnZ/gawW3eBgYKe+V8Si5
SNbacArZX1Jjoy502ADgY4RXBvFQ5JySrwEN+PZaHjXrzT1WtQEUWqRdkKdg
/O9HyyAfVJY4Qg4lHKZo8HBIjMYB978Dh9o5U5r9fH+QmMSo0dVOT4PB3ent
+w6/d01WKWtJPYDc1IiE7Q+/3bAkvCI5sLE9sJxIdj91A8IPAs8xWyGzarfV
p6q0XiA7h2KRZfjqCZtDS1etZZyoo8D4nkzohk4Et/DE4ZRKooAh+SMYrfVe
EldKIAye4sUbd/tjOyV6RaVGZSK+wua4YZRqcEL5q6sWGheQB93V49XBMaF1
Hb1fNAm9VrmOZuqK9WAvafl+Z6lOgjwxBUF1kBX/sLKEu+3GBYaMJMgWHFai
RAZURWUlulK1Sbt/hqxMhRktoHndJdn66UsCo1DcKs6gzwgtMxJ98oY4MbXQ
fhuhZfwVLF7tzwmJkznjPL0qbe/U2mLXsMjETB4YuuZ4sv+5L5eaMAu8eNEE
9yWsksEAcgGTUEF7/e9BhHDhNUbavPymG/+LVysWOgd9Ta9QKMMJTPKSOezB
oDg2NBr8IYx4PRZQdjA0ragqCSIdJwKejXm5mLQfYcC1NjkrT4oTmtyhQJ24
Ar4WD+4UR31HPGQy6+k5NDpafx9fQgoM72pS0i5RGKeGc2qzl0i1puhwAQfn
vDxDjnc+7+5QgJzp17PtazORV9N9V3SOICCsAzrfFZBDF3o7XVNDNHFM0n2o
8eZz7aYGlX90NAURtFYRYPM+TXG4jYakTri1o5ty/cUPy5foA/7MI3xY3tyD
fsrViwelNYjfzFr3Gh8RTzWytfJ+hfgaIQJ2zOuPZHjWYIpOavfrX6HC6wou
qVTxdPFuMJuv2NagL5nIuKH3WRqroJs/R6qrP4jvpA/bJoNOypCw+ZexU1j7
YTOrQEJy9k8MlQ4h930NcCtVEqb2HN3+zQVd6GwBoI4Tc/gX8MVRUzzkeVPK
/q0roxwtWxOV7Z781VpsEcfGIfNbAz8/x7kK0LOiIJmnXbfK0neiDS+BVu4L
MXpWjGFrQ26O9ZlUTg8+eDvk+RpwVNDwf7D2GVASNbojpdhLfbqoG7skAl/X
LyzQZZoZh3N81wSATvTZyLmeJ63AF/moidHHs/QJK+F0xZ6q6gj3Yuvdijhv
zfBIauX148xrZ5rjY2DVCxDD46maxv4P9KA/6pYchOojdjVvPbyI8QyR5N75
0OC7ViJflp/g77CO0CcpLkJXsjEw5Fiiw2cwIMo93hXkC1zzivcmNqdgfpnx
A+RPGIUg6VfjgpqbzS2eW3Nf10gr6VLiurHbbGhSQsP+kj9ksctK6JBJbdBJ
GhwXU2Ym6HC+WDvoQ5WdPsuU1AFg6qbmAzHI51A2+OAI79yUXBMBPRBEGSbD
Vji6GsCNpIc8nG2Gnu5RJ2Ve7Iv7lHa0b6/qnQaR35L+m/PaGCqqC2wepBf5
3zH4YbSG5AJPib3SHacc+xXXDElSYwy7pMuuJERZtoi97UuvMqgKoIr/Cycb
V3FkMbqO2Nu3nJp9rl4ZGTQGzOknsrvwZIJuSd3G896yov1bjQ+mfdvP/QUM
VUCT4kkjrYXOkaheYuZdbzoZxWYRfQvfTu5ho+3BOY177ZLNqX6poMijbrdc
phqFHAo7RhRFjcBBYDOrt7FRg65vPqaBGYOkH3rfS0FODvLQkjJ/qhIPatnw
iASNh6AuYtkZyIZBJo2xHwXNkqQG7/1PC24WONRwdWldygxXORRnTBohEyvk
183T1wydOO+0vOE5OyIHBpV8oCPNv5R6K6UrwrFgZyyF/vn/LW+NdzYWPHLu
SDk5Mo7Hc3pMC9ZpblGpbv1Kvn0u7BueGtoPck6pHVciuvR6amIvL3fcjUPf
YuK5TZxEyvppi1b4mEE6iqVkpBJqt5UueViSRw68NK6X20iDJtZZ0f3J0YFc
qiEyd8RUO5Jpyy0p7P/w+QAq6RX1Wkf9yl+6MUOZ+f7e0R2404gMUy20jnQH
4jce2yj8hFWPyoD24cFLJ6wBCV7KvJvmTVh3dEuLmg5ZRt7UVIXsyCXm8MNk
Gf5+Y7FHBncrro9dk56E8RLl1H2WC4qszX6tyCrj4y97kcQ3DVqG51+AtluY
7a0AIK0VbmDu7F77Ik+BuhiYuYcBJ8EZ4ZP0g7wkLazj5r6hAp5IkKD1Sdbj
mSBQzHzfJ/TesWOToGRYkiaqsVIyoOlkF1/v0bcuzgzW/Aa7IRPtTouzYCNU
SV1tX7IZK0eqxTuTTdt2v1vdYzjE4vxOvsYnyffcnvftFRqTQy4qgpuHkPao
O2KPcmydXr48EJAhwvaL0mVV+RVqXp5ZO9MoB2/QjbiQ2j/8fg+idcNwJZJR
dMRrAjk/WuIT4jNGa3+uhesiLuJL7PlMQQVZ5IxQNBcIG+9NXuywdJxJkzhE
bov8DAjjXrbuluk3G4XQuYUYxA4EaZkDwX+qslhBzX7+sKpGgFDJDArwi6m9
BpK8w7QK01Kf7Z8A1nBfrEO5FO/dFz1mvNxIKvwfTydvvONZ87HObnfZAElb
9GeZfp5wsUeNLYZ72yKKumsWRs9ROSVj6xxZKsk1hgSPClsD3Oi/WSCcb1so
eYIBLdYmhAF9k514Dn2NgCDlFuGsex87hOTdy75cDGlUECu6zJxE4MBa9Bso
G2QIXK99641+dm77zTe4pgPSRiyqlIofmGn/epw21ctKLjJzl4bw35IYrzZZ
mpQoofwUUqP6ps49denxe5Rrk6mCV149GIS++VM86QwPdD+KDLi2A+AQ+Nx3
jWILoksyCQVgCNp3mgLwofUNqpr0RP1bg1inYXQxKMj4MP+i2c/fRwaWquNx
S2zOUdCG082wE1ZSkocYbVQfK2cr2WQy5DmAnYoYipZMM3bW98yD5ft/KVrU
u1AJ8wqWoDxVqNMO1dyEL+AatrFxLgyANFS1Ki3/AOfEazsl/J1wjclGUUm3
74v6y42Vqdxxt8zY5hVyjL5UQE8p4FlSnROwCLWjM6e0dFvQCI8WsKrh7O/0
nel/1VIuHqz2+vVRlNHENzcSw6L6OyLTDH0Tmzya5uSi1ycXktTcvfjCqXpc
qJJfAPtIg6DvP38UkpC2uuwMLvUZ2T7AedrWZPI2F6NteOiu/WUiiMpOCDKa
hY6E7fWbp2C46Y9vULOT2W+QrUOtOYsUS9bq6nlJ4NDasmBp5DhHGpFJhr7I
Sf/NrDKazH8WACyoCc/WoOWY0Kmx6be7aSJrGdzQbHCgvipYUQV4aGtDVm7o
Jz0WrPn4tp1RBvnWdfsXOlvSWXtkU/ia/Tu4akqMHsGmC7DXK7AOnHPYKrtH
p6D7cpHZE+c7Eu91A6Io55+VFM4ojPFgy6o3V4fmgpjgaQpKj8lDUgyXyr7V
4XaeZEt/SEjSi7DbRcvvjH1gr9DgmzZLEJBJplmFBxfpbVP/GaR5rRUSbwT3
zrAMKncYTsRv2hu+NMOYfHkf4c6SnFRR5EBM5VqzTofScuEaAbrL0P8vNU4Y
L8QaNZRWX3WuQ52QlEsuihZBYbBv7ye8B++5Isxf+YJGfaXpxlKibKnzkH0s
4Ksu7KZBclFIA92AHgBtWFNfn0avlOU25TTfN1w8b0ITwcW0AxRE/pki/Fck
IuhcHwggv5329J8JXQEgf3Ip26L+FZtZ0H8iJszjEh0xC3cukIJ9zbvpbWnd
qlBBRIdWN9E5BYkYClg37z5XN0SURVyEQqlnS8Zd0awCGgn9rvLyiii9ukQW
wsJu5e7F6jKbMlgK/ft+mDfQJXnYQ3PBlF/XKEhPm1KH+FQ49g6wOKfyXtnA
wTdqtQhGbzjraBpTTyNoWZIEY5pAv5+K7JsOYwq/bqrF3DZRY+Ff/yic7wW6
EWWEgc6pJwatoxtgl1k0Z9y6LhG5Km1kfISYkVW81U/45iNunQS+CKfiavWi
4pSNRsVKTyGNJ3wmS7n2IdqQ6IAR9ViVwAdX6PvjsAPRvukwHgn46T6T9BTg
g3mSYey328X9tgt4M56tg4P5ph7XH1f04Yh4u1mGXSNLofDg3jR3DaFlrJwC
Nj56A2DgUBHW+fLmZ71T0cMDJiM2gg2tDHsNzQLenC83S/p/8ox0teTwHt33
HfPUHQu3Ou1wn9brG58cfUjFplc6Hi5yBtke3LKxxlvJbZoFgngOhDTB1FGn
CK9l4T5T2A0UBwC7gpp5nw46hnHmlMbEnf+Q0RsuIa1A6nDiacWbCY2+pasg
JoUOz2zlLeHvVyeK5nDY3Cgo1LmgiiXjut3CsS1LuRxo1BbZ9zCmOYRzqa5N
kKEDIzDLfa3EfWiVklkCb1Ddw31udXFBiAQPutPpyOhyXQJST2VqFE5CyCrZ
XPBCxX3XufVqTOZIOK455TGNwinbQJUs6ySZDYHIdla0nHWjA+foRn6GqQU1
ZzlgTldqA/ZYQWd4q7Z3bl0JCrkGOWSsaAo6SHqMiFnYKsBshAGxFO+R6L4N
tCgcmfeeS4JqCL+TY8iQHdDbjpQZw11tD4N8nzhfaY77JkY91yMHp3jJB0c9
jdVOIDQDHTAcy3zH5RMVw/hmQT47hkUL8wgI3uFob+nWY72LUb6EEwtV3LNv
IhDuYWPJ2cnfLfC5lP4ONwc5d3ofNWyD8jwe0Oi83LRwpkpFaKZCjaUNHm8R
dRcmxw6DTP7gItcvCgqagYXmToVcWqB3gRXdVtc71x7+Ox41qRPNwR4AWiq4
NVvn2GZL1UB7Alc3ri7WSykyhO4OG17vZvpa75svkNxwv/t8cCJMNn0/kob5
e8e8oKaTrA/YsF+nfaM3hF08HyYTFE0tiljtH2yEDEIjEVnm9aDFUrc6f+VQ
r4ojPi+cC72rJwRjsZWYmoIED+uIQHUVxUGxgpHf9HlAlZJk1L9m87xo644m
HjWIfWmImNhuzN3AtWi5kDlBUIpesQEHI4eZM6FADfVqqiCdwXVicdh2vXcp
TCw2gqbzZ2UTQhVYEtdGzP7WGcODS3SSn4lgKGU8CainU/5rJcFeIDMEkjMV
RqLmyqht4fSd8yDo1dGnZqls1xl0AF1saAGfUeUvop+MLcUwjn/XLptDCPpq
kYlZO/IUADsbsnj1xOQS5zku74sAt03MuM1SzhRJ5IbESBxFkyRyYV3/EMbO
f3BPhwtp/w/oobxHDni0M8LZcUMePlGqR60e0oErl03IfzSdf76MvaulkfB0
2Wt5j9so1ij8YYNN2mBFGoktMEanJ02XURNJo6kKO13/4XKhK6lsPAUutkxG
ro6ugdHqYbAiEL8EagXmlRxIMZ/4qMM+TKbCWigaAXpG1bGN1B0VmYltyhXk
iHekBp+thlDFx2HFDtUHUa0w46Sp0fjqvmnxY/c5JvtcX9KFbBj2cgLZjWzo
hu6kooUA6vCH2JvEw0GSPYdMyOEnPem5xc7X2HCFR8aQV3x9H2pjgZ7QiM4a
oHUfnRKeVmfe+5cmYZd4lEHBVVHWdtKbHF1MIg2aUjGDhfN2NwMLll7ylRiN
Z2aBJcAO08xN7HKiYmEdhMvuxlqhl2lJfmbRSdNw3uyktiKgB8Rs0UvT/K1/
uZLdcPxLLqMByHNSqlriw8VTpFgZpcGdOMLGS8VscSt5w4Sv9LCf+tpSEy0f
WmBo5BSn0ps04Tn0CGQCIpDLl1cQMrDGGdqm2fwBszkth83Ds5f7xHcVYzrK
F4aJwRMKvlN7nwxkLDLtA7Oj/QKi4Wtt0VEPIDrgOQW9kBS60zKQ5ctEYYQG
1SxWTVCZkb3KnrooVSF1cnbx9w/uRCS4C1e///kSALtb3tHgFN7I9GN76zdA
gGtnOL9gmbyjzES/HjCZ6tQAWcVdYJeDN1J0u1gFwsI0JFQ4fUJdCU/1eThf
pDbrMzGxQqU1kA34y0vV+wlXcKgzqVbdEAOsA+ohMmSn67ONxdw0cnV6CZsW
mtK+bNwcH9QN6xEhYwacLbfkNGhWpJIy7UXJUq6wtbunnOXykrnfGAT3Wn//
utu4h+c07YE5pYBLd4Dr+wlhE/R+fh4wfkg/dN3min2vdbavIPQRB7m19YXP
s9u3HAcqmqIGZOZH9mie/JlhCAriNwNPe8m8UqzwQyEyOryDRh+HpciOY4UT
1qf+y/hGkPdA6FbxhV0N8sA/BjhFkvna38l5CN/ulxG5MEwo5jDdYVrhZ0HQ
8hcxhM2Bzh0AF3NmbyLsVB3oKNsJOwYTka9uO6XUzJ+GmiMbO4QsSF/rMMcE
c/yEcGu5hLQdWBPntp3ttUUbWzvZjRqGwaAyIxS8CxgvSiWdQMwwOb+YOC5g
zwWXw+lt5D+UNGpgTPaxv05vHSPucOKBHxz3Dj7EAG8huqk3COwJCV6QFNq4
dtI9DA/oZKUi8K/C8KQK754T1+KDyUdJegBzPHCll1nfbboXOx6hNlx9aGGJ
eqDgN5sDpyUJh5i6xaB2t1xlfkMwn2HkRU4dgVLomRWR5lp6tbt8OQi7Uowy
LmFGxthZMYEtWFKTTgu5zos2vQHuXAOQi5f2ByP3i3cIwvjjwRI5bWkZdhdD
e/G0gvBy638TefH1o2pLIw0hBt6i6KPtYkIrPP5Hu2OKuLovE2UVTPBcLTjy
XTwxh+uv5OTZ1H4V6WRYXmcow0DOAuQv1QkKWB2Wu8ln8wweLW/VVSk8DVOK
jdX/+Qaz0Gq0z7NVSknhMm0+4+Nv1DbBDKOvWRZanhrULSUWcL3wtPfnhLXl
37W3aM5Wm0mnobHcMMvrqKskTcksRrwLTuelTUdIYQ7618ygpW2NukjYNymU
B4BTOcJMWx7eP3dzUN5IcM2wha3WmsoKFggsak9LFy2Rg3/LLvX8FiAp5Mqb
grH4/rCAEFE4+QFK4t2pIytQwuZwJRN+slVDC/aUQ+O1+u9Lb6fppTpAjqEm
0j3wSNCg2ka22gth67M9atsUs9oBEdAy9K7WmvsMhprBphHrZ467bHKEujXw
zY6lopR5zMPCQ7tbRToRM2x0lbrXdQbRarkgCqIfERRMgqiVZskWyW4sGy9x
tsXg/n3Q0zhRaPyS/5MSCVUUjf867lU8fAA0ONFxpeXKsctxKUG6kCzFnuVO
1FfHVGSzply0f11NL7jk3yCyq/50I5Wc2CfFTlb8x/Vpd43kzjMMWs39ED0j
d2TaUjOvVjvzrm7KYDopCtwtBDECISwYA1BUk1IPKOFslYu5/AICjOEa7sna
Purk3/KIxUy1CPbDiqt7himgbZ0p0/BQesqTOJo8quXZJwmxeCGIW6hXchFu
GSfwKS+EWmeBJPboKzTf5v60ZNNbG090wNFwA6U7n+SErvv2BCP36EkZrpU2
57vNB5eKiJzlkLB6XJ001kbaLx3kdaHki4Q58le2mwIkp7y+7XtdKrEaiTXC
cTG6zSTyysFMeCq+o0J5YbIHGk2CvJAlVcop5J4ommlsYv9mQ5p2Oxy8vV6g
5nrw5DTB2F+FuPIKyEko5Vr/4l6Sa4uBSIATfwgde/Md+BK0jHv18VQb69BU
PqI2tjdeULZEfbbW1ryzisu6tRwIT21OofdlihkT/DC5dfXqsG3huWoauM0k
UzCogjoyFJCYX5r+HPTRe/1CASyGd2+4Sid2T+ToFH9Wvfn3J2o4+A4I+Se9
UA+Cv4fLg4lRJyKTsqUk0A6VJLlV7cZOxpku1YeuoPeS5ofvAG2DqwOmMo4f
ygHvIfP3MW11yf0sNYxSn4RX4S796YuDPUlP7I5YWfyIS5yO41JTscGZtxdv
M7Zs94l1OZikTnmMP+ivBzTM6wfiacObHm/ljn1qAYT0naTQAmt0sf2/W8qo
gELOMUyjSukiynDKWfXePiFyjTYS2mzjPa4NVmBcc+ikKwmBY8gUg57d+sqD
GNrVebOE1qwGY7BMH8WdoDZb/Te/xm3Q6iC8Jxj+ySf1H1PNSlF+tyo90c1d
XWc2uRXdBqSndwRrerga4QsirN/2+HKQYpcKuAUdrQz4wzVsNByLj7d0LSh2
Yn7ntOEnFoN5nL9ZzG3YDxiZ8RP62/kOx61bYXkWYCJ2AoVVqY2RiyY3CzDg
fF8pWExV0jEL4TRiAI2LzQZq60ZY/qDO9O4xsIeUIqdUI2Gz481Qj4ka0buh
7IGOj+xUMnUYkdEYWQbVEPfh/PBpesO9/7bR2d6R43b53s5hB7mO2xyXadyF
LHj1IQeQ+rEfF+sL5TgoJnSUBiqUvDU5Vfy+YFqq9dLX/7g2Fh8lgVoDXiB1
aKbG3DbUKuYUUlhGCmT3enjygEYvkvnaLZc1ThRysnqPKNUh+j8bluiKhj+G
9S7fQCaZGti49bU94HFZld9XwU9B10uUs5q32VCp1B1DwfPuV9XbZpX4w2cg
xK3v9BWjvenanEC41ZMX14qm4OUHgrtC/v14AWeVjGLSInVbxMoB30MzhQ4N
Z+IuR/Jb55ouwt/NZOoEuqKFiFrCnSwYEAzYuiLgyf+k6P3RvtIktr7ZP0Ja
eeXzKfPccGrc+iItYvVdzYLQO1yp3JjSEY8vlERM44zXlGPEKydNw70oW3Xq
CFAy6TwCWgm7kURPHEdr8X/vyDL85J/8ko15Zixqpw7iIPJlzrwFFUeC8PDL
qbmvTfHn+JEx2o11m5O5SOLCOtrGjitHEFazuyGTPzJWPZC0MYTTYvY7dQMC
aZxfljBCVzJ4dUL9PtVk+2rhHYU0ly8KcIGTnjEJs6TKHcr7emo/z32Te3PC
mbf7fAXhi3I1Jyp5l0KnL62WOeDpC+m5FXIpiAbjByXtaOJAsrkqldjvPeS/
zlxhCoQgrB3J0Y/JiW5e2a6rw5b25IlWwg1N6jxEsEDhoIZsQJmfpoM1kNq2
7laYG1evtTr7tkYQZCfogiq+Pn89rB0ZEHX6pyPLfZBj07UGeNNep/VIsgNR
U0yUKxr7ubVImzSKExB8yhaDz0yBQXdoktZuG76yrfba+bJssyKAwvvPAnXD
fplS09SOh1G8/MXxRmwa212kUi0eyDX1lN/q3gEUuXs/UD81Dvr7j8WhiKXR
J7GAF1/FCReVJU2wH9WtUu7tXxFfoTPuXCdKSG+pfwPi6FBmN8Vw+PTEh9gL
pEH+3plhSzVjyzIINBo+KyYcET9ssqbrLe6Hk8x8pyL6P6NAGZi3ZK5YuKEO
vlLQVbVZ32USMffPr2D+7Epa/K4Qnl38ZF1YSCk1r/SHgOPUmdXmJb2p7aNr
bSikVTdPByN9DtTIhL6Jo0aJ4K8aUoDlq0mCFcfa4ZHRY2Dr6nn6JQQ+PFuq
4L0joR5zCq7CiWIImch5NhtXSETmiaqEggz7uk9uPyTGPSOM1/Qxduexl+ZD
0m+hfJ0qeRBs6GOMFP53CFkqmkbjl50eT+40wB3g6L35HiC/FaIUFpYEJf01
a8XhUlOWA6H3rwWYzvdsVabz5Bqa9AHGAyQTzitiDyDXV8XK47KkHn2IInoy
QLI8PTOIJ5sq/pGm1QQWZfWpEW5JgFMNCx8MhrAU96qwQZf0Sy8/CdUzG9ld
tZNWEBqLsSWwupm9b3XG0JYfDhupgsgu9v5rFp8Gc6fWDGNVwuqPAnZVqYGP
R2ZHU5jNgppH/a9OBvvBZefWt3FWwP3NvTtpBTwWFBiZzUlj3HL2hVJDjuTO
CIFD/gNLN+p7ggcQUzjqRBNZdGooDXbX4Eovxk9JlRJoRN7AS/CzKzSu9UfG
vPf6gXy+chBtqBcjJWR2UHGC/lv/5sa/fSMZ4xqDf6YvbxAW2zvtV3IleAvB
JKUYb6rS3S+05NQkAd1HQGiH67MkdiBRsiFG7/jyqT94VkmVtOb3dIfY51mH
bM4IDMnPqV3RCsa1YgCLXbloSyrnrpDdzs78sfZwGsizDI46ilvrejHP/Se1
MUbwWmgjmjrshrSrKyrxIo+kc+Whub3D7ariXk/402vMO3jFTJMqVdjWxZNm
acALawlTVuu0v7S9yhZ04iAYAbLy9ss0/jY4IYanMXO/uxGel7ezKdaC5XGJ
eCaM70TCfjS4t0m/0JNRpn7VmA4nGXi+HdCujWGfpUPR5LXEvQT3DuwM3Zn4
eBruf1bslv1S1Aqp0GBLrcSr2b5IzPGAqxx3I10tCSG4wpzWEW55836CN4qE
ll5rIfM9+crJ9G2d7mMzT9btKmpw4oHhIDvSt5775YezKwuh11ShE+jYvIpx
FN3EA0Gl+czwvKBXNhiRM817TXFkgE6isDKcXd7NxyZ4VqB3VaHVmUXNw9Qw
9Ujgfx+GSLqrZHNf1kdTM92cMdtuN4w6E0OC52MSHopbx/Ou6Jj/w+8FRrC/
UuhbUvgjkFGtzqvM3mE2zB2f+yXHIhZFPHrh3v/3ZR+tr0QmLED4RjhjNngD
SmK8Z5i4s9r1t4gMEUegw2sbD4Fl0NbWWWkOjSmpB/twooi9T2LeLRov58nH
OlWOJlaXByeeRJ5Rlmx1bazRt+07Wt81+cOIAaAPzdoXvawJGRNyKDnI1wVV
rCSWAZztavEOGWvcHso7qPMv+AdGbZi0Aovx22u9Mt9rpzYhqzzjpVywqRsu
G4AANNNnHcvMO9/vZBVrUWuH23OMQdqu86eunKaCDJjpD/LRWexcpmZHukCO
KG0J7ZFDxJHO2r5KNMrvzjmMNjtX8Ylh9jJZDN9b8iX6262nPELBl6JnbQf/
of/rgcoqv2ai/pLT9bSkO8E/lPYhNahoZAFsMXIzYT8Ag4JWgcMdrkJua6Jo
hVY8WM6Y28gYDYcyyySGVtfHpKAOJ+haiXpeBCwlj4ecZ+f0Co7GXMOn8Yy+
iMn3Ii6jrnK7IS81HGMM23UKyHc1r5+SwYQD1Q+Ql83eJlWimQzTEF0T96lr
Vw6DB1nIiQim8v3mQe1p23xBEmSzf6ZCBnHQ5esl6eVzz5GghJakP5FsxbA+
KyAwDrO8iCvKFR+oX8fOGyPqYFfq43SC/FdW9hho6C7jg6ETFczYa40AbToZ
cZBkaue8SyWMGcoxqZ+BvR+/7Pt7Mgff40/YIkzh2n5piqzwf28MeeDPd6Yc
AliAd4XgKGFS1KA1Lhup3A0LE5xQlMhCh0kj4VBZvsCfQ+odm4QnJ3Xcj4q/
fYrhrJOKuN8dOMw40d7xnC4YpJMZnDX+Z5AEcPRVOjoNh6o//WN4Cj14/Njv
1mrDXfSbxsZe56n1JofUar4H+WaOlk3qDHrAYfp/kxclhMwLIuSuFOZpJ+4W
vvR88NodBKNsLQbkRtTkPIIRnovWgrTlEJf3p3Ha/T9P6v8PmwwDOjezMhGc
CAmzcmGvqE4BJDorHgac2rPvoOp+6vwHEDulx8mx3QgeoGdGNGmpkW5+Od+S
sIdypo8sF2TR/HujfOL2wD1bVS8nTXr+Y8w1Ru35dJ3ABiF9rR8lGg/wyD+P
eUI/MmS8qMLot2O+HQGrllB77EOBWowMXWmDfb+UHEVqKmeDzEjKWMs160CC
HDCLAxm5EwIimQzIhk2gnuAcnwWnyV/ezRBggLC/xD4YJ//szd1A6WjN7hQu
/s3W3EtJSAmXNVTRA3ci7h4jyivmXuWVeXgv+uV/ivY62rqpBeQZoDil/Uvm
DyBPeoUwiPWemgO043Bh+A89hmDL14g3djsX0b5c8cLi3x19pSVXw2p5Ewhh
h2yQ+plGzi29M4z9EarJTAekXVe8V6mbazRffXygrpcJqYEo6yCyZQt5AMJj
TXXkhnzn7q/bFdfYs9LQQUKq9ZOfkc6bJTvjJ0eaO3+GoFRvKpi0px1BxF84
dlkDBOGkTbxO0K66DY0o/Ck/eY8BobscRrmmAzObc18pS3Vd5t9RmfloBN0+
6o6KYgBzXlUibsqGVJbAVN2AnECDRkLWP5prfUwZqn1nAKYU/9oqBwKdXNVU
wGbLHosWOsJd6OWD7CluJHXQuiuo5oTz3nwObGIZDPTwksaCj7ECrLxoVpGA
QqllViWIuPrhlhFiz43UV6KrWaT+OFU0LSfp6Wcb+DYvyGCJV79iz7/4bFHt
kARsxUVwzGFMior8Tsv49PyqpWEPY4w8I7DbMeFAezXsvq+quvtag90ylXKm
ZhNf/EvXvwkyqYF6zXflkVYhUdUFr3rZ5g47C+IzHvv1yB46upoBnirgOP3X
BXIWS8ZxLZPXLcrheEmmHQlB4slTGRAQbnlW+W7dnAJ3Zh01+zWOIbg0DSJo
Fj1DwSUSkt64o4Q0vJxj3ADj/sy1ssrnUgpTHY4TSPKQ0WEd3orcwypVNhp5
bQI8I1fjosCn48b+ZdJEhgemu2He3TiZquNzxMaoVUQMocfxBHqVV937uG3+
bBmf1SPHcV5l0xOiwG48Xz4K+QzY5SZVjoGobMFFAD2GTNmntgGteq5hLaIy
+2ISUUJCHdj2JLnG3oMrIYgs8GcYDwtyqJyvnCL/+P7PdKqD1vYZogUqD11F
wAXybO2opG1YsSUZA6LV8NAFKjUILZM8l303082TFf2+NEzYkuYeF4Fq8V7E
sR8rNjAGkb8zpzwSIPM8tw00g+mlLAL+M1HzqcIvTID5RV6UlcqH401ZbsTU
hO19grruFgMRprsiauAhbBj7HfJJ2dWriXhaB+yWH0NPKVSA4riie9unqhWM
21voMSDR6271Ap0BBym5RQFzyB2p2ufxYrSl2ccvdEQSunktS5fkNDsGzKsu
wC6a7d84jdorfULLsVpVhJMQf5OfgkewLR3aorN8j6iBYSgqAwNABZHtQy8C
SNSlit5YuUzkNJ8T0JtqKJxyDtjYY4pONIQ7sF5zOICgff+cpOBjq1Be2R3q
FxXfAPhUX/fE+TCe52CIkPnzQgJ+d7WP6eSOpscYa7oNtEyc811NTvEdta58
XjDT7LBDjXaZHW5nIMUKwXs6D52F7a5gKEdvEjFrFy96eXwKbcIPvcNwuwoN
MlGN5W1Q7zSzOb+27u3kRtLX2EJxebiF2pzLynmxHJZIitgMpIe81heeD5ox
ZKWNW1DWRdFKOf1+HcVb0pd6Zo8RbP+ERQJVXWS7B3kQS9Qce7jVt/ZyUQzh
yGa/Zvxt2hQdKNz+kGAy5NxuecAGzm6iHZsPACvEKgLetpShjtEi0qGYq4zz
vKLRatYBlS+knAd77nHlNN1PfdT8V6se8C6nHxnkspC7eWiigwGaCY8XvPEo
XdIVmqWk5WLJ2DkJ/vjig3tnP+pO8ORs7BWsL2V7ldMF0kQBeGRmoIlWj9iU
KBQ7QIfjP2sbS2jj9A2ocrpL/i20Zgz3ydemOA3a/NLUbTp1n59Gl8OABg7j
0REyrSmWqQu8lkyA4X7n+KGjIGYXOV1qRaOKj+a7vDcWz1p4DTKMiSgI7qYb
X3wo2AoL1jdVWiCBq1HbEZlNvNi0n+2vXPwa1AWYs8PRckBQHxBzMlihEWNO
IjCA7gqQd4/kqL5EoO+q4LaLo5rT8/8TNGD1o9l89fYvh/0lGqTtv0xY4hxs
yD++plu6oHSbRO9tNx9rwhgg6J2sKYV81g/YSP2S/2jEX92ypN1kLXfTQ6o/
hE5DrzCz3T5DOcn+R9BSDkWeNW9lhJx79+Ur5zoqiI3tbvqmg4y1kkT7zxzU
swvyqKftS4XeShPfuaFDWqzpYO0GbyhbpklxdVgPp8/XhQOIWbNwoqzgV43R
Jg72LyBZ3RlMSdLMtclslQImWPAx4KCWGZI+jH5m4cN/fhaYkVsm62Q+qoKe
ls72qRb3iP7gzq74PpcStlyDN7Y5H4RzRdSBphs145J3xUeaHrXtrSBeFerK
7hxN4QW7RSU+bkShjd7syFk0HPxJSpLWG2tb3LSQs4u9yf0tY3gW16mlYEG7
begQ7zLquIdUwSiuFHXKDb3a2T4CK9PuVCLrN9fcWmoWw2dRAs5R5G9diAVR
hfXmjRKnFK5OODsm2+1EzqkrHWmG3D1nFvAfXNdby3v1VUN6LLFTfR+0ONdU
DUOik29GrDOZCE3yme5PCB7lPqnXXG9S1cv3Z5Fb38cskTmkI8qMfrRW0JMJ
j5GTRUnfNWNqxDKHjstfyTASZzRht6tKmNmtqrsqjQZTIpGuQJVc/h4xKyNF
AYjFIBNRCzX4hOpyrqoQQZbesQmqWxUmxN90PkQb8u86TDMjpMm+K0MBTvMz
HB/sz35yjbrVL8mRF+Fx5DgnUm5SKPRNAkbJphmxYT7L/pTEelzh/iLq6eG+
seArLJC5G3lRhBaThqk+/DxnLk//6iGgxjUV/Qt9KBO0oZHU0qpE4Z4GT5AR
FyYawSnEkpxgLgbiOsuqPUpC9UbsT4ywV+w95DXTXFrAplhY0WhkLJ3Me20Y
zAozCMGB59UtfeWQu1L/NjSBDEGRK/0XT+Sth76osJQAc4VAhNoiFW68KinO
AkI4lWvzM8EjBo2XBO40dlubgZJrgCwMVGZ8KPmOL1HPI5b44ZXrh5ZOZDt/
uHaL/K3Wnt6IvQ4qm6X4XCLgwAIrx6M9buDthSKBGc9huuf3swD2N7rTos8B
lHL0yETDEJu7eYmtyHYB12Mgco7C7VRyhatgBsWJqBwa+ooraFdL6AyWtTen
OqmdtqpcHDbN/l052U4sDkQuYM2n30oGJiR/WeR0uZDCyU357osNDjrjaLfN
tGwja+pkd5U7SZ0fXBorwnRQSXvjiGRk5VXv6f6Rtj6U4sqgip+BsDBhgtx+
9RLVu7IziEgRFnE8b43y8kkgbh6uvom0lTKm4LESO4f7sxdhdyqdNDJCYFRW
LOu6qrMWdUR+3y09sz8i3NunFLVVJKUBEDsAc4qSgORukPbbq1qJ3aHV8Uw6
sZ0DjAKLxN9Odg63KL3A8BOblNwK2Jz7lrjlbCIisJu2pm59MbOPsVj7wu9M
1EFosJrqGFfJ8CKmUV8xpoCuVTRqFgIc7/KRdFauuUyPLw84dMNsts2BQMIo
5JTx3m5zHUIYAX+uSi6O98dUyTHZCR9YQ1R3D24JIIdpk5TjiUx3eLSOJkx+
SWDwxJStOdJE0HMLAdDeoxG/beD6Qvbk6IU3ilusRuV5WstPgkhk1fhWVUNp
UlGLQmlO3E8b6JjkNwhP+wF5kTrhtJjm+LcgYDwnup/5PxPXspoHuATwX98K
NfwBHobxpAtcifk9wIaOvXrfBFofjaGPgukOhXoIwl3Vkv5zQtZl7wwIoCoN
/NQVuSUScAcwtMtrUxMZPTph4Sb0J37J3jKSSXLogR/Joc48D3E8DDJveX3v
2H9d2n0mJzbdgZY5VvhBAzOW/w48fb0afGkkfy1Z/KW1VKUakGMgOzGHnxGl
8UEAInBjU5myKjMArdrXnZPq4UpgRn8ljNYGBA6csfmIXBbS6USgVKCQQ+oi
NKu+m6txzrL4zZpkM2McxYG33qZMxCQrOZ2NxoWTnEvXZ++LGcFh5WgFLveF
3xCpuWJTizPBZiCONEnKbNNjBXUQscGlWebgIQMkXWnCdYbgXtD8gDkTUD5C
X3Szl+dR9hWX2KcaiL4t0U00aG/avjVoTPgxneMb7NRGfqjHwMka8AgoI4JS
TRoKRinDFhmV4wvKj4Nc3afaqTbA06EpJaEEXc7iuDPsUR2hKNil2ebh6Hh4
RbttIBbCe3tGe43BA89r9JtUkGWN54riG5Vg25RCFxxSz7mvzPSrHZgQuQzP
KJAcgPov4/O1qAmpRDa6cEyHBDRFOUON8UsUkKGO9f6fClzXkj0kqxkNZaPX
fYgT+7JZejBvmzF4phYnaWNpqxUnD8TADeCthZKGnDEspU/IebKV19T9lvfw
3ahd7RrYlxDg9gyhxb2RZBD7fhrfkxTTbhgLBYsnTTD6RX57ASjVf8YL4okU
cjlZYHF22WxsbbcvNFncI1zHIE7urLJP81mlzLnkr4NoO6bNPEtbDykfui0f
WCDqfjCSHRua+dO+BsK1Uvp8+ZA4ec1Q9JYO9ck3DYOxo5+zxJ7reDY7EKoE
6Q/ytJhAkmLA/tXB1fmsEg68xh2r5EA14d/c6+3p1zW3XMgWzEypd1x48f/A
MdvggCsY4WxQweczhu7BWdofMLpNmWq59QGUd84+nYFQGKIfd8XN4gaZdfCL
Gg4hUs8NauIS7HerOXtgAHcINmgMdkMnwGOaYkuXDFKSKX0qjKk+ARLzna3j
60Hh41fyh8rhgju2CuVYQ3xVB/wsgVxOSQyYzQwvu+au3wcibBrkOxeR2GtK
9qrpEk1DY1lcnia6QWNABurmFaPdmHjfmIHc4M3T/J6F0MaYuyoSTgn7rI65
Hs5H6NJ+exsDZIfVKDilM0EDft3l/pU2Jf3FFA+c6nIV/fksCsjuwb1wMjEQ
07Qk/C8B4GbETMePEcJ9KaEgZIEJZK13FO5nkc25JY0wd/vnJVpemrD9VsL1
RD3vmacvhDvKWXdO1Hu4zVT1jV1RerUg+Q1ordyrSoV/Uuapv/VfHAR//Vde
v5tbeyIPVjYMIqgVNQMDn+fHEFe90DhqxYNVuDTqh7iWlhGCV3oeEvOx/WYG
AVq1QB4CIFzNtJki3LCRuOhZhw3Z8YHfYWz7/aWlj0ETj1aw5Q9+l3FcXT+9
22lPJiFcsyt96yLqquvgX90uEpdu2QAfZaq4p6dMp2xZjnqJ+dyNQA5AJLQl
TAU4CKAFFuPSlLbK19GeTIVG3FZitwFvQA06O3NiuNA2Qs7ow6qPQQ+9Yzo+
PQ+XkkOODa7XzeoRq0N2jFsgPLVzBty6usRIUQE+Vh5Q3yvgU0pvZPWA70iL
uFHqfWvRWl5yIzPZ8fUUsuD0ep6s8S0bw51DAuvapNnx2VsfCvFajHj5O8Hv
YNcMN4xL/WbvyUnw/GdA3wpcMKmZWaNTXPEw1yRTPQGC0NfHN7mytcKNrm/1
Bq0bog2o19huTmypUhju1WiinUgNQrqPiH2d6lAdbs9HaMeyh3yg+ysWn4kh
0mMoCZXaFmM6TTMyWbCrpj5PCTlNE08YWYmVzkx26sSapa5WyPJmNMwnnNpm
54qn64RmPZveCGhRx//zhfJ6LECJEm1ev7fRnwAFv0wanzjmCKYZ2ycWXt2c
ydUQK7d3ZuivdrCgtxaZ8Q4hS3CaFh1nmuuXmHHgcD7j7ioQD4CMgSOOg25C
uXjBhkSG2NSazvnVd4GlPnJZ631c3ucs52UC5jYWKsbCVI6LGT5JWhIzEeeS
jqrKakkK7ndHf3zebbdkZ9SEpamQrcsq1NbVVUsCUHwZfGblcZ/iuPry7yMo
KN0gzvWHKvQkxlrtUQolWSfdGDuliUi9tMxZsXT10OnXsCTUHAgnwc51QwMh
nrBJ4TQeu3zezeCQQP969SE3fyF2vISvr3VTnHv1Dv+eG2yu575mj8QfPToS
giBj/S5OsmXuI6KP3mDA1nD6uvWg0CNvCYFxtOzWtkAMNyT3PQ/vA/H9T64T
l9xH8a+jkwGaNHBLd5/DdXcXqYHTvikxNscF5m2aGTLts5LQXIUwkyGLmkwX
J6x01OEXLwbfJcFbdwhgkL05Bs41fSW5SBwYuLHvgfbuAniclgKLNty3gGaP
gsqmsW5gEjiD0BqSw9m79h+zB2f6M4cs2TqbnWp63z28Nn3UGyAiZEp/i180
2Mfn1GTHAOpiO2Rtoc2s+zu5PnAGiUf84yBTYnZFTDj2ZmlKIS00qNPEIMKu
yTXT/dLZL4J4TBs3uynxZEDHTB8YVTww5sWMPYJnCNZr4JMzDHKJWqeHFyj3
CANYYcoUhvQD4FO247Iwa3lxbiRZlK3L1LrTVtvM73enbiX6R3cAjBmlXVQQ
y9Duv3ebYPxGZty4HiA8N45LFTpVfAcGXmFn2VeKfyWEwXg1wj0vNfnIH2fN
qXgsrlJbLIDKHeZWLhfYgDobcM7xOO+kAsDb2pF5HlK9ngNEGKP5pTmwcv0X
Coq8Zy/PlyTmW4Rf2ed/2Hsr2DM6DbNPgvQr5hP7DKP03Id8Y5UBS0BliygL
9rswgt0TcBFG8gRZ44c2z5HMCLIgdZELziEnH+yIYc+FBYiPJGq+qVpkIWOC
0xU5JTrSZTETTVSh3wHL2uW2xQ+hEhmT2ZXguRSAsIxp/tClhAUFCh0IG2og
w7F8cID8BVCILxbW/1uVv8GP6j7oipaGcG4Y+3tTxHXs4c5yaWPTr1Syx0Nw
yb8rTfoOEu0HL6dJdfy10XV8sOksy+rok1lssB7c+OALRB5P6wtB14lR7s4/
+41AO6UohFhsFeQpkc8GZ/ZCTv5pphtsCRMgwDc8CEkRhOUITECkXo9+sHp1
eIjBTBXGWT1XIQi3EV1Z/pAOUwlRtyioQmqw7p2qmPjIQGjO/VoLF96Lf9RO
KtUc0Uqu9H8JNzDC8GGrKZU44AJD0CziZBOGWesL5Cw6uiyoArW2ETBduzja
DOu9yPbg4mO/ZSvx2/1xH/LqzKZ9G4f8XMEOxLoaOQ11Ej7wq1kN7qCH2tJQ
8e0bppOkBW+v6ZL9g0YLVKfn988FKHfCUDqpOlNz3rRBHupXIvoAvUTcj1VZ
M9qkc/H4pxqUCpMDJQGPUib9L4b2QcCTPHOkpZC/P9CZs47w8fzQ7gf/YKDs
UWiy0hTb1DWI/szlz+BW96F/YhjINNTli+yg5jS7W+nwuvbYstmnBhiu9TG6
qbx+XEPeenY2oRy07x5rAbari8pkVMek7LCFA88x/Ld/YR6ypghWQsKn6VB2
z/wrJXqm1rIcBEfK7EpDAdJJbQMVbQe0JBuXes5JpMqhGzf53QkdopG89Msk
Ja0WIDU7RjMYiJjDiqL747zcHzNaPu8vTLaVMIPIA2hriHWoCB7XDM3ApPQj
mx7raeuow+RavonN+U6meP7zecwLfSXRoQnAVhFXTaoKlLisVhKDImE81YIv
VXFFml3kxpHxQKPDGDKGf9BnfQzeCC+fBsrEenhbbHI18JWaAKTtRs1W6qk7
LA1j2WbyoiFkgQH1byzzxQU8LemzhJMkSZg92cLEXUqrhtEF37ogldu5LjLj
Glg/0afsqYUlJuEOfLQcXfFlrmF/sw1gS6R6AOoNluwz0IpoIvNV5HOWyABd
ol2gi7jtzDZ4CsdtZPrKnLUkVMisEDP2f5y2w6TndCLCC86rVZtf7WL9p7+P
qufMzIy/cENPc9lBcWDwI5Zl9X8kg6/PpcG/wubgxpkFBR7RbkWnJrz51xZe
Mmz1NJcuG3vtYlxX0wzwqlU4SADPNR2g3fkPFpPp2oNUKLM+i5q1BGOfv0hK
E6eNQ9AV/3FMJpA1TjJIdeo0ILzD3H0wRTTSfOLG+2IvSGZzxyLgmvKt5DQV
q1i1fcO+JVb68LV0erjF937E299FVxUJlsQu3g4wulmfcxmoEM+vWoYn1RJF
B8mQEePPSd1IZ1sQiJBH0EurOgRme/WBj98wMZ8MiQDssZKSCtRvEYkOcOOO
/P2vL4JRcp9Xio+SDXT0saZc+5LU37+GKl60oA9yP6ey0x2pETgU/XWQU/AD
7/1j2tMVsbF+EbWY2SaqCkU2RSH2XiJbobY6o89n6tNXio1/r6uAPxsJYebZ
ypuxAmeX4RmBQcfw0kFm+lru1jiQo69A8EvgikxOYnJ9ix0b/qOgjtqvdXUf
TP+lEU+/+BNM/LBMEw9lIqtc8imL7zX7+tOI7sOOBH+DDDVDMknqUWxDc51M
ManO3QGu1/P4FKzxVX5hR13jnZr/6eYBUQw2vqihEd1BV6Sxcwu76Ys71CIK
ZJS8H+E62iU3THcpeno5UWGuEMA6VbVo5HDGDL0o+mjEStMoPCdFCAssSv5u
SO+gtcXjfv99uXgFM9HBxc81MgqEd7lCxiNwsMnxrrG6ffWIE0C8lh6jcfyF
v8uMq2F57//HoV6hXZ5tZYQ6qPSybATlFmvU4svpYaCnooyRk4R7+AhyRWZm
h6tVD7B+Q+16zHZUm6SEJthH/xMcKEYFgmP6CnTdw8uDuJgnIU785UfDLKil
uyJr7ibBFHbIAU8pRNVXlfrywbJsGW+GAwVWTCBuxruNAIbT3JZbPWW6csTI
uPKfkIi2Rj98StaIdEhZDVa6WgCwHqLDAAPhCwaAZudU6An19l/h23lcrJI8
4i5sd1LINGCQ3JstLDflbcoRxm1IppRIba42Pkz85qxBrL4oh4nPhiKCgLUO
GAZmHvA2jsHgAA5fVtoNlpFuIlqqGisj7lovMee+ouq/po5KN3bMCPW7t/t7
4vg93q10hN2HDm4I0oSaywkJObMhhEGI/EnbsyWUawOwosYDhTMPABoYU3S/
WEoXB22/q+jVhOmUuUFpzH9OR1pnpValbb9wk36ALplXBTwOB2kl6VBe7lYz
YwPkhms0TUKWcx75g6MNdnIor1ayaJ+BjkoJDTZgQvnQ/pz1sqTxkLc/91oN
mLW8hDQJwGctWo+iJlPky3sRTk1nqDwy33A0uQ/6oeVY3vQKE36msXIMoWAF
oam1MyaCba+ZasHocrZaKhql2fhtyzh4E/8nuv4qDgNjNaFOfIheWAZkbmRj
ppR8fBWM93OflYCAsVs7MItjlKVCgSG1rA8T2Fi1NmvVxh0b7K8n6IT2yjiS
U+Nd8ojul1bRRUrE8avzAEcuWTWVxXEnDQ8wRPCQMQKZMo9Q0KBKxR6kCojD
3BS4flnxfFEWNiq+Q6ZmuEmV2VY0/HwriXSSttXDDFimqhA7Zoo4GotVd9O9
8yFWKSJxSbRqm2yimxyk4yOxZMrQvEuCTMq/RAXoTZKOtJP8EW5NndpK+bmi
W6rA+D2pX0+9bveLcin1sgK8UwQ9x6pERVQ8J8GSbgLI7PFMzLekgjXT5uVh
+A3jW3YZywFv+GWRQqm/VaDnw8G9rziv7E4nqH6AxBejFZOFq5JZYzQxSGaS
bFLfDu/xiH5wU9Sl/Jh1Jo7zBEb0GhFqnVCEdFsAOjjFcrLE1SUAy7WuZfwE
ygPxSQuQazI2VVczPfnOxhf1w9WosSM8HS0t4NYhLpAHtLoUo7nNeOfAQdVK
uw8gFkqdJc9AQTflf+1AXzeJCf4qovElmZs8t9WG6mKKc/5zlyfT4RMP+UDU
X6CPEiEBwPJV+Nt8Zpe5X1rwEHpg7LpDOBvrVu5oHD+DyGVDCMaj8hNIS70L
5tBPSVZ3RD1JT23OQXCd291nZ6rqBKY25S7Z9sp3tThtJWiI1s5FZfN8ecC1
WaVCigF59THaLI/LOeLnJGc1IiSY1d7Wt1EpnMpUIsecyDIXU4ABqgDSaRe5
biI0fNlrn+3vpZbZMIJEYf6BrXuPhh9BKBhWH+0PsNDsqZfn1jNOHF6D/IEV
omlW8AiM2vh+xjYTCEA5EFGEBjqkzGAjJy4/+iGArrHPIz/b67lS0Mb39Yx3
eo2YHJmucjzEndoGNsMzOpnkgttFYHT+W6kZB1FJ0yfYCBB0PaItcI6Tyxv+
zQXtG6+M9ePt/6LzspjQKkNSRNuzzohLEqf/2Qi9cA5MROA6E5mOmT3EP3XV
8S+aa/V+Bv0IpUAycKyt8TeQZ05/lTtXS3puwH1TTUtitRXrL4DX4oW2uktg
0OTEoJgy3DOhjyh9MHyWjDL4morKAckdQhX3xNnHSScQhWPEQgQ6swjLh5Qi
R7iEolGQIFnJvAltHOIHVc/Rz/+l+5Esvp1XjomqcgYu/IR7vonxVJETbNjT
r6LTJrLSVbN4gtwqPCI1ITcEh+AX/sGURWpvo8CsALxhkuuX8raY85TfGz14
qQLqcj1MsM2DkqbTBprxx2yugGyeciGLnH49dJkjb7+eusgx/ZPtN83Uhwly
wVnz/3Mb42Bty9pgQPRbbjyQcAdJa1qZGXsoClmscSaDloMxFDLnPyrbRzI7
B/NYaD037rYzbKTJMpIXcCLhxtwAFBqx92crkqu8nVLYARBfKS+U+4amZSYg
BGOrt1SGpJ4/bvFMoYHf8Dy40TNkuqPWE4K6ASF/b58FlY+4zNwMqNMaFNVa
LjfnKY9h9IPMwct4CFvqcoYosPzBcXiJBnxYnAk4tFFYh4Pw1B9tvOPRY/sR
v72c6kXfxNCd0xzqw7cYnulOrDzVsudPumOcoIP7q2n+aGnzSGldUhVAjYNI
sjV04jJ27YjEpEavjjgemVBPVGTiEcZVPLBlZLWephbtK7XE5mWdI2uRqp/n
pcA6M99oEGQMuhIb0dJ2/P6dse4PqB0mywoaE2ewxxlov7R90//vJgdQ7p0V
rCv6dC6UEPF7tW7f85gAIRMXqU2DmzujgU4OBqDdosVOrSmqDftbjs2NjWyC
H0ywrodef1rmdI/WwWv37SCcRUBfEEptC5fbdOGFniiIlYlZiEFCAGNmY7mZ
T9rP+Npbqds/kSiVnW6RY2nAiwE7d0HCeXLYLgBVsSstgYFNEgL8nGJIXX5s
ciKK9/aeVAcoDXxmXS/dvobbbdvAI+i19C1v6bex4qPKZXUOkoLvCfpAlhIJ
EcxhBxyldbUpZTWNBajrjEdvbTfOVplaq+yf8YBT+xJ5movSaoX3c/GGUd5F
BzEJnQqUC8yTYj+6tzi8nKhASzy1hyVMQ2iUHAlERFzzqWLeTbg0JhU2LiVW
2moz+S9ceczFLuIToKTBN6MwpJBj6ewXP6nMTULeu0pw4DiDGOz3gCGyCryZ
ok0eA9oRwSvYKEtVH/haFpRzsOihAIoHL/lb5mG0F6nzqZWG+O2sJecJDBCN
jQ/ukicH4HHja4OlPf0BFIY8/yr1ZLnldHJmAxCiOU924tKqCvvoC01E+X/V
jEEVIs5LGKL/6yeH7id7basBxc0W7dUfBCxD5kZSa0nFqzlTLzJ36PedOauj
SFZiDdzocCh4D28AqKkbriplepYaQYNLI0Yiqm4Jko6bZTI6FF3d5UG2VaVD
H3hrhEn53l0y9WIAYZ3D3AUP4FiFLQS3tmaR1m0pcYUKijS/EnwFinTmeqQE
U+fN+O5VsnZNVXjlEx2/2tOSeQs2LKeHKZ5R6wU6Tp69cSxUTijewFjmmr6L
gpGejZ1rvuAQK52nt1mLtQOTuAkqdOc+n5+mawTuv8uu6JhWe2gfn6e1GW+v
q+kblU8X2ed/z/dxm1NqfkehldYVbXGmUBDDIx0dBoaJ/ybBdmntGJ+Fu5/I
1rxqWEiyzFOTLDX96KTpVTEPTBG0e+Y5MUjNkMGZ8mi+vjuKVtEagbCF9Q5B
aKPImktVuGVexO7rsFwp5/px4izm8PlC/yDUi1OHrFUr6IAZW/yBHzyxn0+g
XMm9tKO0MmYIXRboTovaGuDg/tkOmzSJwe5kpap02HBLpikOLlU6y9TZIxXO
3tU25FM8C9neUEr0J1gnS5qs2xXwkpHDMAyUu3b70JnqvMYogvCGzbIiBR6X
RfXMpIAYnApYdsakkkvJCbKwszY7RJ1gA7shndAHRNIQSVv7v4wM5YDV21wk
9R4B4hrlArTvPZCEN1c01xYrIhNxAHuLmsM1occx6MoqK/4N8ir1xOpA0Vb2
Wdx16D8AAZqTIiSI4ac6PPYq0PZ50Tx5/XZCu29B5HzTOOF9a1ikLmMc4G3y
cQ6SopRK1RRAZNDtIpc947UUKthGOYJaBhqwaR+e19br1ls3PDi9BUyG61hi
zD+NXgo2nUhZXO3f4fhndHOwCCTH5HqdGEMmXG3Q+O/dLxLGySgl7oJ90edC
MMtFN0myMaMaNrBrWtc1AcyimqtMj64sRVajvUXjL7PiWRRCRWirsbi5ZB5B
6MBGxE9IvbEEGsUJuYs9I8Go/k/AijktjYrHefjpD6wrzq9Dv2wBPDuhDUzM
OFCXmsabSaeniJCW5FE2tuXrBfb2jYfsYfeIY4A5tAtmwiqBAjtDPYiNOkfT
Y+ogg7+5utCGQHTvI7QbKDo4ayNzvvw/2sbmHKgBpVtxnXSP1kMyo1eDzrCf
FImnks3veTFr0B/MXVT9WxYFONiPCombpFJpbtFXOFZeQ9ghO4LZ9iAGzfLA
zGULNngXHcrKBYnIpTeN4AOUZSQDC3vBOkOytsNdJP3982gKf3E32AgZGVje
z+c8rSGYemTPvj9Bo/1i+RL3+yT3+fMVXvgG3FLFhYgfCzVg5hc+GvTuUW7m
GTxvaiceunmq3VHKYJEmY5U7aajGrDDGbL1P06FcMZLqWJsTrgUGwYYkeuRt
RzAmPtwcejXSpyY3w+9xScdVTCmZLvha2nrACb2cjO+ZMVtpPEZcJiNBuZy6
BnFdNcBE6fSUIdbLQQbggw5UcNJuY8b7j9xR9fsPUzXS8RAj3tp8ZG313Z7g
nNbBKuX2IbCiFAq+NCspFvR1QZePUakS0H1nNEUubYd9y3W4zzYfBMRW4i8S
G+oQ6NPDCIC1AMY3gxNoCjWNAcXw9RjHVjV38Ok9zVibO7k8UMjad0vt/npb
gJYaRBD3EGNluLSlGwbf1tpD0rckxohyEu71MYAY466VRRI/ABaV+fMmkrtI
r175T5Lk0Ag5PMMum/n4iMjODigw56IMr/1E6MaN4AJJlc+pexBJphNGXbkE
BdQ2+033uo9asXkAj3mc0DdvlyF8a29GbJmgRrwddn+QVI3m8KgrGUT5b9QT
zHR70+xjaPLCXVnMLg0CTpjF/NGeCyw8hArf9V1OWUr43PgQ2bD6TWB1h4IS
E/p98Q+x65jL1FGhtJa3rolpl6sEqbQpFXwhewIMEJvpuqc+FkhRJ6FzZPOT
SS6LFUxC6eS1ZyYqP3g/nq97lg5ZjYNgN0+byEVXApAgSfeo+o9dCtWQQn4A
N3nr4y9GePHUZ+3+rmmmnOkI3sa73tDZZHFGU2uvwSwg+uT2EEMi0xhNFbVw
4qSnqZpbyBNrhG6IgCosVjRh/r4A/6R2/9S9wJtVV6k3UX7LopKHXgOgJSE6
xqQUsvjdOZSFQpnuefsa39Qx/OXhfgILXRnAAKnt9aoC8LI/aA5Onq7n7U+Q
LjId4yoC0W86kqolc06qZwPkVy3+IdadtFAqE1q6Q/RvxfrB05LJOShYK7ze
bMEnVSObqY7ZszLZ4ACOriJ2BBv3503e26SMl4vUSuyHfR9TO83Vk6nCvfrN
95NHBOVAsC/aHm08gC9r1lBXbtg2EdXrpRDlGVFq0QiVzk9UyYS8DYnarIGG
27TvAXskj6hWkni+/cH3JPlpd2BKtolshJSeY2HnLYJbHE87JrP27kSVJGU0
SVFDGe+kqjKR/lWeK8Of3l23tNJN8wnsn8UlMuG1wmq5M0vCVxbqCjOUYtdT
ZqWjb5GbyW26yVzRkhCvOehYYxknXGVqb3laCG9B6W5J5j8lgU+l1feolgxi
xe1UpzLMPs7GYuxgrtU7AMUGiqJmMmJGJXIfFQcgu2uZ5jSRWQ/5+SG4fRMl
CU+xpwK+mNjlFHV4A59lWspJhCJK8qeKi23N+6i7aQgHA2n/tvi52efHku1f
okcQq62BN8/ttbfBCeUu9DO20f6qMhUmjGE+wK5bhZaBHEdSbNFZJBKgGMuP
0JjPi5AZS6G4vlZxUJ+aijCH2t2EI5KQg+pYTlU4rGqZb2zEhFYeI24WR1pO
4dH499y2xg5/UTGsIrx8yv7O0X2uR2TX41/KqeMBF09hzrJ8FajBLfqdEUky
W1o0U8UFlHYMJxNNAWzlY7aIiBI/fNegmekmoUQu8jw/Fu3kgsMHXUKOmwci
Y5/dvc2P4seKY0FTZYrzfuHkeNUF0JJLgylmGdthmlvHHedxi+kk+yHh5RRp
HmYzWjftE1tFHNZ0e6Avz9m9XBlVh/J6jfMlPS2BPsbdzO79TFswzjBrlSMj
MTTlpEpYptUsWJjgSZr6WNC3iTQZ6N5sooKrIXBB1J31FDTMaieY/oJ/gAnz
soUS+znNstFbAHbBIBx0XE3Dvt6ZMSOkWq5NQKxQoTjjILkFeK2ramT3v2Za
vMvwfqab7bEsQ5QWPrt/GXvJ4iq+ga+vjAHcjG1alQyKTTj25BkbEN9FGWav
gdt/mzMgmv3aIo0x4CxnRipTaLGpeTV1v3+UQmPtNqVW6/jJWKwZ4weECC0R
B/CR+YQ8LRuEHZS/qyxCbdvrMPCQPMFnfx7uAqCR7JCps0kRUdeY6SrqRGzZ
VmZQUfDbDs9xcqpVUvTc0MZT10Bha77jwdvRbA8CVitvEA2KfIPU/s08llTm
bHTyvT1VwAVE/I0mxY517j88RacRXPfwW8IqYl8qFpsNvYs5Y1V27XIVZ8Mk
fn7aDyghqbbrEpji2rU9pBtwdbOTrUE9AwA94LTpyDC/ro792DAhDLzkpop2
mOynAGU4nlRpXmVTqC3Y2QxXxD1UGWeiJZyEfig3XD7+++6mAByT7zrLLkQm
aMZi/X5AOHC3uRUl+XNRK8NnRhBfhlwjPRQsLR/rj9iGnG5g9jb1cvfevDFa
+ODzpLPds+e/MJu35M4N3iHV2/VtOpF9CtKtEOzVP3DLD3KCgKKzgaehZehk
eTUaDcHkZs/C4HF7WrJgOoFPqha9cxLghzclq5ns6Hx7mN2HhD5J60mTSe/w
j4aqLH8nNKL8vlEqd1EmDJNVCGURTWRwYGKvcmbn0nIaSE+MQ5ipsBPiH6d2
Kh5mBw6UYT0GuWMVRPifR02SV/fvjUNiY98Y/e6YevIYAsktQpJuRlBhnalr
qK77gtmt/97xydj2qH3FPSKpjr9dZaqpaczAwn6Epw52MrTRiJRFHADban6O
VDdObZ6PyDirLcR65z+lWl44yzS+B7pyIQq82wJfjT3FQNaYar1qB9VaohJI
4bLWTo9oJcW1FST7nQuQdrB2ESccl6CBCgxiVNR6Xik8q06F0qbhrQPkQXif
Tzb8rQVBtr1RVzWHO8/YSma+SdW3weJ/WghDaK30ghlo/vE0X4N8j9Do8iLX
1fp6fDYTyj0Hyt4UbRbAYxpJzdZKjzFPzg7kjE2Fk5ZfJTvgUm+dPKzRvSLm
gfrgxmfo/lL8gxd9XxTi9thfFGK3E9M6aMGzgEgCRh4Eq7raQpknJv0RoGms
LtIwSIAsoqlQ5l5jInY43Pur/t7Xe45QMkHlDFBxXlug3ofVQ/Oj6EUeuhZv
tKAvMsyFupA6VNhTuuImA4I3PyCEi75GUt7lU/OD4T05Koqd1q0GAXhoFL8a
OWFATad1YigcFyznLZ97seIqGoZqtijI6HCwDtjLWsrE724PoY2E1Fr/zxHP
NyLHSBUf2B1HDM/OHpSVq4hCIz0tiUDJs9ZM9O71OFO+vn9+WDlif8kaf0rl
Ni2NNu8v438oUG/f6GzLjr9dGiKaTs8IUEtUKjJiiiXsEBymhJI3JEtCKq9x
2xLnDYhQYv81Yrpt1IRymLSVA24ncDkzdXkBxiNGuHJ2SskRB0wSiGKiOZj1
uaIT6NMLpRZJ0txXGzCN5Qtw2i/jutOnwoD7s7zTb5OCLdN+zE4xgc/awKB+
tP/qGOlOlUqdNiaPiNlWWwBOr2ECu6uN1TlMP0w5bulWO909Mmmq0ekHBsfd
okTYbAF09tnETWCpiMVJGryIHtCYftQ7yC6yPC3h8GJtAOb86AJVUqG2sI/u
SNoBP/vb8280kBWztPyX/7reSsmLrRrP89ItKyBgjHbCitAJhdgbw9tzQAKu
eCzBx5TUmEJNOJQOJtKrzs9Xz1HbpqSPslQeFo9eetjU9IZrsgMmi4HzfN5j
0G+S2srb39GeljrGM/f2GcGQeEkV3jWfqndh6SzeqfL916vmvudiZNpW7VI6
CELF+OarMyvWLRMN9Y+i94E7NNcUkSJjKxd9cHrF0F1V+7hW/3F2nKgUCQxb
AC5nfXUtofxyT9piHJhezJjPDpWC63rl+or0LTWKwQmha3dCAHl3zSnrVPYS
7aEcAvQWM6F5ZGQJ8DZLup3NB2d5RcMK+a54CRB4hwM1LSn7rfmRemGrcWe9
EgeZqhjQO4rxbjbVHTLmACkuzZ/3Fw0eCwCN11LRH3d82x3Q1di1U3Gnj8uT
U4QCU4c5OOvYvrR0PEu2VknhDPMCOedpo43dlOjBYw76Q2ineRQ3iDhU1JTj
8FuXop2vdcEHotgnKnZ67h2Z8JV3EP39uHTSP05FoqqxzB/BAioYZNqXOccT
T8UDofOrm5GcWYzOLj06X+0Iv/HrcpWWUMsi6H8pBbAHVgVScc7C+xNO6+YQ
rAIeEOfAqlBNIaRzjlbP1yVUgVXTbzwsYFidc56HCdEx+9P+F/FFoFEtGawk
brCxn3dxRGvStboBnVhU2b2+wDGkSRMY9rtY+cNpDge7Hr1Ns96fIxDzAc0F
nK24qtC/ovJpiMMOWJbCh6R5Sc/cFA5AI+FPhxS2kMRB8QaR4g63faTNTFug
uUFL3yP4Ka9Q0I1nirJXw8cYbzieosnBea1Dd1XEWyYf5E8SgKCZaGzgHvkz
5xoCeXbfUkHyonnPBPx8S+4rewbEB9VLOd+kmyoVS4q8+99hXGIvNsh3Tepu
CylVpbi3eFOKm7RsfGhef+3AjHmK1tWp6wPGbh6XaahBnNCP9C1RWq4jgPpb
lBgiGBr3zEILOctLzMUIhy56sZmbhhfdS20YxJFga5Vp5JUAXY53M01wGrBc
xCLDJZZfDgPZSZ2xwKaf4/UfqXNIZqr0RWYV9sLn1YqFjAacqo1stP1YdWSl
gzwodB2Cwo4q/QLfUFp3WZQ15fyYuDx1WccrmstI6BPKXDEQgWekp0m/NApK
s+tbOjd9R43mPNiIG/rtYSXPLz4GvHQC8Zl7jbVRUPUVCY/TB/rnKGrDEBec
6mTuqj4t40wy4xZVL4YihhaL4tUXJf02YgcMG2XOt3GDRqW+XnjgGlhebp0i
V/Lk+czGe8Ecqe2OVMDCTYVBvYYXHoDgvd8coSLOkLHRBGw9d71y6rn9sOJW
YoPFoNpLSit/9n5Tmzw04nr3Z8oap5OsXqAu+vwnUDhQXWZAGlBWTlB9myLT
DxyWYQatBjX5zerLxlDw+G5SJj/jQEX0s5nEoCRgvPBV9ceiC8OfFS/17Gxt
rxF3Q97rTl4hH04diJvPkAlAmhjTK4IPxQGtFRgUVi0s+bboUD6szcghIVKG
ejRx9jtio2WSkrw+tOQJfMy/YKNG8dOMMxIUr38kdThWhaW4p8Ciz8WDAAIy
6A8Nf/2ccmkB9KV64iDF0e1RivFJIoUYb3c/Q6WiUDSiAx4njlIOr/oo2ygR
eMeHdHa68gUSDa9CMkjuGrZn3g/Kq2ko+8v35sqEtOG/5D3byDC3yspMAz/W
+3RekvHumrbB3Bhz4amobCsVaDCPo2DHlSyUA6FDK1WYpwWFf5HzfGOKPYQ8
ghP8ANMmTcijeYnADJ3abFW0K6pWJml+MtSbHVUjIN7ANGwB6dZoS/2HEsTn
lqablct0mBQO2OyNTDYOM01v1hQsLXxmwJ8Qp8M9ZCvoQ5bXEf9uk9J3eMak
Kh+io4YdvIdzZai4EewpdrHy81bQQkfq9Ar9PGZbXpcwfDAbOCbAN0BhzTAN
SrXNyr93jJM8fpvm3kLIamT7unu1inVSnI5b59BuD/tiSbVg5UJKUGsUcUI4
9QIPf0AcKsPa5S2sCNaT76jG/KpySiybcnpe1v3O+J0VRW/gaRCiS7cYFErx
F09aIfAQa9zO99hk33abEZXTsWltwg8KR/QTgT3jrov8Sww15vrzdQFDNYTX
9RrXUpsH1mEcJPNyF2rYSoTd9p5Wn8Ag02VeyTh+ya583SDig/IYVc+7fW1l
rX1qJMjOdEKDoLKFFNz0iRVkut3FFWzMu9EbW3CmtQ4C0bMGHPw3wn8A4mUK
c0As2M9u7bN+dru5F7193mWgRAZq3tPIQ7DHaid1S/lxO8D0MCQUmnlbANdm
OPONvDxSGrGi0oOt3Dvd126q1igsIncOycS55NEkyInFFTu93Zaa3dIYkoIR
7N17spgXDGgqwcoO4YtJf0+XzncFsxARMWIIL1SqjQoYo1irgshx9rzpE+b3
H8iXicL2zltKZ2SgvBJ1H5tGFxxKbQQ9Clj99FadVgX07NLgVl9oKIyVaRDn
9qRAwbUBIYV2mxdb1k0jbgKekCma1zK/Je0G2tT9/c1m63SPZs0uKTn12/Mz
K4SFjeL0HECaPKrkuxqjcZqSTOaoYl68aIqhGo3uH+fLn38SwI42i2ARqNiU
iZT0wuEgrQ8RsLALASKAknTbTPe4ZxSsV+OnRc6/EVerZKNDdsjHqpjXjkpO
y8zEOQUDHPy6mm0F+TpHcScyW8UxPfZvX3at5AkL/4cuo9cvazhXkYCh2U9t
fhh9EMwEpCKN9gNsh9yV9qDXDn5tysdM82FTApief9WLwtXFk0fEOtWKRpcl
feNxOLs8kQY3VUxAlkQ1SsQg6cRtLTE22JgwZ0DPfbooGACJHMwVlrsTuL2F
ROCIR0EtWp7BSuj7igEE7pDr+ePD8H36qh1EtKiNGUbaiAZvD9Y5mBJMYk88
3rgIX9uBfiuWRD9uoTCd6dczo9ArlQcyEZ7Ktdd9aQbzu115R9ZB03iu7oHh
zhkKmkV+6n1hQ45ndMz79f34qUOTzQBXaZrnjbgxzv2Bd2U3LzBZ4SdNqIrp
Q6ZeNSbBh22VpHMor0jr2/seQ49kHsUQn0h1PnUy5P4EYxxjItvYxxZEo9ia
x2GnwJRQUsAo3YVrwJxIvx5LcSRgJMvra5i3Rn1hzw4JLlXq61BTaSOJYmmi
SbBIeDeCjTBjeg3GuMJtiaDEA2711X/fgQ9lap1Jr/CgYirVCCQHKJhFnEzN
8oCuwMHIdHQQBbrXlEly18hN32swRI3cVMVfNVKz1HsHtLVAdvhlaP7N1Ugl
4EOBxktDLj0EfpFjGZWc1s/Jfco2+pI682Z8vyso7sUPSdEckyzN8mUCW3qR
aNsJJIvfIWg82hve+952pNx29OLHcutJy2ZPLj4/WzvYGxDc91kBGNhBjcmO
E1D11rNIbLxZ5l7sB4WSXwOmhDZVx/ODISSgWW0CEom5IV7LFFbWh+AWKaiG
J4NEa6DUeV7SSOdP2caKppnqVW0bu+T7YP18MDetAsx9z58rariTvxYDZuvC
HtAYwg1CbPVHN6XWFH0TsrXjMSz6zMiL/7wlSVIhwWBOvuLSneaHItCGSy2G
CyQmeroXnXZwBFvhYBEhDWUHWR0ZBe1KvDKo7N+BR32yz9CqajsoFQd6kKA3
VKj4phW+kMvcFk3i4eSF8/MhMx+7ViSwTtx9n1vGMlLES4n9qdNTRYAR2TZO
Uy0ZSlgF9M+TWaOri9+tONvI4In+ShoaS9wIQeTtE9RuNryyznV16pQt8dmM
p1eUKqR4d1lWG+igtTrEbmtx6YvjGxcRcWAQeVCd5Ni+c60R1qDQBeEoVzbR
cxYWuHx2KINQ2XQmN6VmGxbe1A0wpgeQ/NUggIr7gwlaW+XZDvQ3VKt8dTje
/UfoavcpNDnBHy/QSp5fya+x0svXKgktBQ14QdjXEvJQNHP0n7873bThxaCU
lYQNthxUrhrLi9LD0Z4FKd31qgpCe4MBi/FuuzxuC8QMisuQJmn8yzelc06z
y58J7V78aI6RcoZqjXw49s9CCRyeIMUHcyBO76Tkjick5t6x2ws9DOKWGxia
eN8+AEJNosbQW4f/gNuGh/xSYsaqu4hCoHgp2Ey88AgTqcfeLwi/1xcT7EIW
xe23W7k/OE5s7vJPnJZ+TKI4gZAz6QKVZRWQ5GNP0qIERrEiwefA0eSbVHej
4SikrTJ3imR8jPmHXlwcPno2amwe9naidO6fRzDb8ACLfYAtS+8pMOG1N12R
wiCKAShVHDIu0zhKF52hD3VUx4lx7u1IM0PMaLKcJMqNHvBKD5GWwW5ohrod
uclkiqUfLk2E5NRfWRGT6qr+7cTwUgolFC6WS84TVCUgE+vxKUQIdmKtoSJk
SpTPhRBdfATPq3bysmFanHPyDsWV7ToW9vG9+d0NbQ4HbFcLCFH/fE5f+bVY
l5POYDTpcEpSPW38y7V/zi8YTukDn4wUlSIncgCClwP3+wAPhQMnZxwZZPOZ
pCQhjriabMjR0grBAxYpzOBQTNhPI3bWbkvUGLz+kvABhjYBTp/iXP/pY783
ZA28L5mG9LYjmrlgNXR/pXLAYZ9s+m7aIXzGv44fjFvtOQVR8jcQ3MdtueDw
ENp2oTX0AMgZS+FDVqId62TNJPyAKrr8pIDCVEODEY2+uXDp6qFf0Ff8899/
xNkosLc93mEdK9PnYVytaKrWP6BToB1F0smDVQC5/qPWBnTU/cn12IT4HPb6
YOEienOq2qpHRQExk/HnDKIQzcoEIoORkQCRuldOtaxobn5ByahQtSOeKYdB
g45bf+U5qxEM8aUW+ljWOATPvt9gRCGvVrDzE+S/tqfPouMSuv/wAK2a4OfK
YIDw30iLVTgZ+EjOidSqFOdXfp37JQyTfHDZ/5VpCbtyPAf1AIyxFa2oMKml
IegeJRMjWv7ALhh68hMvXc87wDU5+jPPr/ooWwDu7u0tnezP92hdKI9og8OC
7ynr4aUgWHpiXM+gENPj7Bqa9I5Eygk1Ny7RTLdPMXvoQOv6g51N5+uwPDVX
6rViU68EKkmpg2jghLNbp7x7cF+FAD/YGoCY2i0zZBQHufOo9fXW2eXSlKAM
XrDZsU+JpXuBSXcOPa7bT71HH/ZVbXK5B5F3nUZMOqYUyN1ssIlrwE2P6s3f
htMGUCyhT6Y+iw8wMjbes+AJd5cUvd8VKS1iJ5Gs3Jp2tP0MjJr7s/hBPZ3R
Tv8r+9U7cd1WXiXk7XbBAAAnIN7VlZ5m68WSe4W85yw06/fdHZDxXF9TOI0I
hKA8oFDQvtKl5Eyxb8GQN+djIxR4B97XGBHGQhhGnUQK4GH3JchO4SJIlhM6
g4vodgbDbiGyd3N2n+PWi441y6agpYMXTPal/CcYLZWRuBJV2oU5i6PYtBZg
TCXZJHQnyaPX5xQ4InKjNvRGrNnhpQWTI15KG6iZJKq6zk8GJ7kHDqVMXrUH
Fy4I28KHiChVdsD5YW0eMdH5bGTVXeVp/GRBbgBRCPvkmiHbHmikAuECS1pz
ZEzwcnZRusyMkM5wA+Rm/TJqhM15bJ0Z9UxngrIj0++T5z90F/g2taeZE7fP
04SmJIzPt10WZwyVmp9xN/oyIiHLSm1z0nhlUCEZAOnpu5UYjC/uj67BrC99
CGxtwUshuIsJZEOfYRNBjeUkx4O58/6JYvc2nS18rjQCZHO9wO+CjWoyew8g
DAKZWyxSuk6WSIcqJewdC1U/mJcu6ONPaHagtqyKYqNIkPKmvAX086cHsWhN
aFKpyoefyUYYCdCQKkxT7S/8aW9ip8N5tjeb7QK5eUoOvLdWaoI7oIwPlG5B
XF3d1vsL9CVfSuz0d0z0yDOUwSv9bY2tIHA3fX+nfNPLiXrisr9i0n223CtU
nkeyZUzTJKbwkx3mJZCVDKkXeaOyqwgf+yZJi6Uw90F3gSInPxxZcdTQOTLe
ozL9jclugrqfzsS6NP4AF8AJJLpSAyTRFg17uKMfmX01EIgl3cDSqAgsWPVl
LNzkyQBnH4H0Y1TyJ6c6eOJak9tPPzSYyUTVdIHkWhyvregyOUhMaJbXjG7O
3tZPwZ8TRXNlwOwI8K2+Yas+Ob27yPKIjtnE808huqGhc28c3riUIUzVlZra
p/Hlub0joX5OfS6ZJjGBxakEs3tpW41Hgv3dIkmmWL9Jd1WmcY4ZNho2PxSE
a0d1DQbJ3uVOET5aujLgmTHdGEi1pk4tXx27gIVy0tQWbgUAtSP/52tJOJwk
KXLN1ed3dlzXNMNw4kLwSApVo0INgka7leyg2/129UpCZeFAO8ZlCvJr9tpL
/mVAF1SeyMcs+Z9Hbp9j3+QdivEyqGlqLT3+vZgRrYs9T+SjUoyHg+pTPSbd
p3MDDDrcSAk6lmsRqZDe3GzbS0OOdxCjJ3KKrL2SOuv8XFeWW2vQv5nd48cD
3monJGeuapyE/ywCv2Sl+DkhyVjRV9I/4GP7ZCu5vnZ8PdGN0doMu44yVgUa
nffOEiFV2chjojme43kTxVL9NVpzVUBLh1BOjV/xu1yhDUdozzeseIsgWSpc
H6cnyMEdM1X1lA8MnrgIznhhY1UVuttx1cvnsUI+fG28S1+JiIJM1CL3eEn3
kb7Fz9DSoWwbRgswCurcWOqolMVZM3pWQOCAbRueZs637fL57S6OCL2AIp1i
GVhcA6I6z6cic2Umnch41M3kGse+AcVVCnDhLuT4MG0R66FOWNc/OmpV/5N2
0PkiPIwwc8prrKnjh1nBNTl5MTwzjYmrXh7YBhARgO3Q4jjKF91WtmEts66C
bYy3lBJXVc8Asihr2hlKF3mwIERtu0zDVcXRml+eK6OalIKatL1E0gIxxmPT
uEtMytFabkcwuUXg8y7cWGLBvEYHGsYrkSb+npBAb1e7lm0Zwb3YvcSGt6/c
L5I2ef49xgETnfGb1uOar2qtxu8sAtmjtX7pWW8BAyHxGnOD2g9UDUpZXyjn
SvmytvCK8ouOjNwLnwuxNanfRGfR+Oat+SFqODoam4C/TNmBS+dHKldVKbG/
m77U8RKsThTvzokQ0SIAC72VxubC1ku4q9QK0U72kosAP7MZlZ1eIT7rUjBV
9bDpJEgES6W08MgqEnPKXtxXQmjoR66tmoxO/06nHcbF4EShWj41wVO6ck9F
+C58Az+/V+d8ltA+CgZ7iUGWEmEzk5POS3gfoPgZJk8GAsfm4RT+FxKp3CY3
zRj/3TbEdL5dbSzSbc9YrjfftbqwgDLGMNTAtaNDDPDOfg4m7gbXakQqoyNE
nXaTO3iL0yE05CMM/Eiy9JhQ/TqTd6uFrK1kBfXGzmUxZY6ggnutMJNOeYFR
lRDSInGZrs/MF2/622u33igxWDvULZAu/iyGpm4hz9CLjuYfxnwjhwUJGQOx
JYlsi5Yulcu+HsijN0dnqAzOpG1L94Cag1jtkn9URqHdcJW1Ma+OWeLaZ48R
VaKWpC218BPOmrmXg8tBibdlPaii0TvP8uPui5beIZ4hC0TyUZfuwesY0YH4
5GfxoWF6EW5HqwPVD9dKfJuzBe5oedQC4kx4vsCTurFhFeYA+Z3PAWrs7/ca
eSU6pNmFAdqdwYXEMrZjEkKsTQcUm1UumsfbjTmplu7v5FYqsF1tqt/cI/Xw
MLtVRoRhWlXecnmua06gTkGYBScNLvqAxCmn+lj09sv5E3hRmHXEsfYmS0Bx
0HLp8TLGUTITazRElpkmZ+/FYnGtoOP5DWLBtmthy8oI9HJzqXrC9qW7bRDh
tLkHK/412rzOsUs/HEuGHlHxW/xzb801iavQJWfNDeqYc3S2gcZ5yV46aZz+
SK+ruibclLhZYBWjSAuDdTuLDi2oDZUHzfIIYPtHRBJ7JAqY1x4zHddFgDXd
t3cSLyElai0TsYN9YgmrkONT8/4zO+w9ku+d0ltf1yWFUYyQhSrdxgrifet3
jHK7syMeNcbWQlHvKZeLbEyVwo2AliJXluhebUBB6YvzVHP1cmlrbUQcMUAK
FaiYNZUXG7tTFqaMmgtzIb4m9B39pjmu9MQ+PCaXtgGtv4ec5WlUKUc6rWg1
FfJGUGj2NRaEj/nzoS7wTufgx3cCNrTuA6zs+9BnU7f0FXoF8eJF9RsVc08a
IOg8I9DRj6Xik43GKE7usxuzpf6FQX3VhCthQikELsFcDg6kbP+5Mk+S84zO
Ga4fNop0ibykpEqSd10L7zE38HWGiNMlgxMdHjEJFqUpWcimJH2+5Irqt9SX
baolUkmz75xP922G+HdIT5IffJTLAYxJfKF72zhkkag4jJp+vXU54Snc7snY
2VAksz4AAHnBqHbn+zpMSnOHKOc8f043QTyGSsr0vQ2JaOq3ewt+UF0bUAEX
81TOa9WrP50wL+7v4RjTiG5WNz/mr60SYBBanbS8wljVE7lef9yukNfkNby0
bAaAnuKaxO0QCRKgzzyuDEAHIgGYz/XfET0IHOYp8BlKmYBzckAh6OM7U+Ah
ngLh9KBwaqSlYWQ0FPvEXBVj/4BELJxgdsBR+X55dU6ah+r9E4UY2uMREe2H
d+VnQ/zOjfNfakBy8EoxGyxr0xaK9akmllHKwjLd52vWB+h4XRvm9XOtetle
oINmnhSqlS4EUaAH1DJbTCVudgZ6O5WLYaZW8aaGoenfrCRUAvil2yA+KL82
qdpJyosTHI0Yj5P0Gr0gd9y6ojV3WMZFq2FLyzm5UPVxFYnWAWeRNaXETKGp
7O12VSqSFu5S/MUEvi/cCNtgY6BP/OYnmG0T21qmsPeiR/Wjr9W57qYxFNXS
Da3m+KK7LhMhiW4reLGYW8W/5QChYWl2ZmUIeB2cQAxz0sXmKiWdSE8rDOBz
Oah4hRQ7Q2jfEeXDL4knuHbuu/kq0D5to4D6ufRDywTSU9rXIWrI4PPHQJR8
zLubyr41GEpsZ6iF536f8OBqx/dXNgaejzNiKH8jsg5/MXHzF+q1Jzg9tCtR
SGYIOeQfHVD6aDPTSVlc0FUjx3Upnb/DDaJcZs+IoMvI6deqUS5FZg+eCMYN
KaqJpgurGwzj9B2SeX9xlKbgVS+j0V/eGNn4e3h488ehD0y7WjBEGZRywAxI
bVDa2meZ3vuCpQxxxF/DW769muernuvxfbWMXZcRuS/vm22QiDgmATPc7YLq
hRXZqlqcg2grNypAbiv57cuzmRIhY+Yyyu08kdau+9drBgt98+2JHoktqeMZ
aA68KcpjIhJv2EEYS4up74ZAhRiUdm6GezDARBbPuSdkUe/eT1pS+w+MNWF7
kclbYvMzChxtw3I4Sg3PSFv0dV8rw91qLOdWYsxxqlmKJpWWHAC5i+/NqKap
a3bYjBdKgXhWkpjekZxZrz1wJ7DkjmmrY66ToPjmY5sL53OzpJm/GiNVhtVb
fn5jivSaB4Dz8Pa73ZJeBE3vwRFxqJvSyEi6zHW88V22yoqaPoH2QqoqTzI2
hFDQGamq35/7sjH2nxGLI16gclZ4AKyNHM4O0vpcRSwYxCkX3fuyOlQFJ+zj
XYhaEPDjLZLkxk7JgVKjy59dwWHoqL76XMm+ez7rCHHaIQEGNdw5pBkK0k4t
UOy7n/OphE3mADdJfeuvy52dPIHwlHNjMGik03sLLAt9N6zFwfnsVL/ONcjV
eKOEZIA/UNC3wlao1IEapUZE+Oob1SoE/torVsBWDnkvM1FjPKWol3prIa15
r1YHwZlH38uDdFUBti6ZdtK2A5DZiUNMesX+eGDubZkAPU3g88CQc+DO0fu3
2iEJpTFnK3VAQIe/IDa8DCndkbbwAl088MxgZzLQxwewAOcKY7W4QFdUvNU2
bfbjHzgU8QJ5zRGG2as8MBTjslTq7lNc6Mj+oS3+/RiSROnJoL2kHeLiQmqY
uijpar+p7I/Xc2BkJh2D9JF02YHdoG+lqEx6pF9Ham7fMd7ea44NuP4Jmui4
fsvq/nYyMi/9DBI7ZuGODNaXvf27Mg+kIkq3CN4klQXYWhRHQe82/4/vPzl1
DUCbzoW0ZqNGLKK6XgBc0dMrS58EpnLO5LJ46RuXKBW24wWHuztCQw9VDH3n
om6A5M9EMUEtA3iD7jgUg1Htt/1Sbuq9zq1OBaALInBO0XUpH0V4wzPjdlIe
qmKBAeBRD2u5lIqKy5hLHPFU8RwAGvyDmV/VjWJSmfjp5N4HHflkEdPzfVAV
dvH+5irYosnizhawWKtriVMyni+JfBbA33f2nMPiw2SCT+4va+cWkYaax/Vs
Iq0vbD1gtcbEX2UbETYBSvelJLh40D7tzCNLAsca3CS6wZf0DB9Ks7yvQ6On
zpqBNGojRS4AhC31EE4X/67JbUMi8Wy/xx2CcrgMB2xAdgfs8+bSTYqVFofo
1NM5uu8xSRMbf4pu82qyYahd6arNo3QwecfOo/ukZLTKqBFZ2pH1VdVikHWh
z8sqoxz5mGPYySLeTrMzSnSm+P2sJeTU8lzV9ePi63yrTSLVbmPetIz9o39j
DMb6wYbQXuLvdSGHHoMbKvgZ2ArkecIE1XbyHLiMvVobFf/f1Dc6MRGh82Ho
BtLfEi9FKmqvvJvffJbcYDtyvPUKbLIxyLOOBCpsrT0bglqQoB9rOQ1zumvC
oddADklD43Lanwr202tBDL9+4/Xu5MmG1AZWG/gtZHAG2mZ+QMc+xXKzY4fY
Sph+FrE+NhaGO7fnU9hIjd7tE1Qgdx/sNZDW0+wsboDRKoWypt/UVMnwFvVY
1buG6y1Sp9P6xeooqj7sf4jMZ38IKjQ1g6IxzDMZ53vDzZ1yYA1JESOZ4BSx
7QRvizaKqzbgH6WeM8zc9Xk1DAlquO0AmvKVOEQ9E6gejlQS/nU6B/zqlJIy
24hyslNiDGck8pTpZ1b7yqxJUefE7aoOXGd4ft6gbocfD7x8yJuRYWgwBOrW
OPQfuqTCYmsqDRBuWAjBHOmd6QoyKp4lgfossfNQDHKGcn+Cttn9PhELmvDk
I2kskTuuOUNGG/CjmffySUZ459vNrgvBGZ/NPgGCSOFcWQziBeFyBl1pIe07
dv/cLZNiuyUiaGEBpD6ffHk/By0U8mh5wgQ/mdQyhapQRd/RB+hwKbMmoYT0
hWFrSoXtl98eos07DM70xg9LFeORMPwxVKhST0QWDjMPwB3CgcVmXyZjbZ8/
bvuLw0pGFBFQpTCpGJGZBC+zdN5hbLIuWJHb9Qck79qNMQb/0AB+biZBm5Np
ykfNeBKoRsg8QCJxRdMGrixDoKUVtGO30oWOcSUsZrK0KR9+/dF4iUTgcNOh
aAyOWdPh6LsIX0REy7nypUArtLj4g21bOhR7gclcwK5j2sDt3vyleciQWNEO
x/pZwp2nn8kiOcPNZ1VcKOIlE6iL2qCwf+NAWv+bwvNEuVUPuD31RoeHc2oG
gda2MYSsJp5+cWoO9rX3y8bdDR0zL8p1XvAfbAva/SkRbIFpv1rx3xAJ+w8t
bBP/LtpPTZ+deJNCLV0Ned0Z2MS1qazuGoRJM5LShPcdSt583H0qBb7XecAG
FDaq5xUbFQAjOb2L/xPUNFuopnjy10wgrcHbr56pcH/9piEL3INheIDmmHju
CnyVQuea8uxKC7pOm31entx3JhyODcSeRkrFc3K1sdpXw9k4UGE3uE+59e/b
VdesPfQhYq3sUOSjCQsT+X7a46d3I3XKtZYh7EBBhE8blk1LfjDDa+wDjJRc
vVACpmAk+RKBNCJDn6Rlq0e7mjiroF3asvqOB3nCWNvlhuWNdjloDRlibjsC
bz88hQm4n7txTsPggO1twk3ymQJraQ4u3DqY3porv3oTxComBidDoxmFrw4p
OxSxHGrt4ZOy2i1Yd0cFTNBveo13CIf8H61preQf7bpU5XhrCL/wtCdHMDcA
dHR+sr3Y2UowOTlnpQ86BkRDiGvLl/k6YZovbT2tNVEh0SZclywt4uUj9Vuf
uTduU0yP4C8gdZe9ik6WU5BUufmin2Qj/ErpoYcBD2/DagbcmICTl8LB1BIM
WH7icdiGgYCxIKsBvKOxovM7QnBiaydn9vBl8rhL8EXbqQf6F72zwOt5JGCU
swnTR8aN2RT2q7i5ctMNIiUXa+/NoNQrNpg9nN+TAERy7aX9qQAABLKRgSUc
TTHTUXr3OYK2bbIl91L6i+Dm1J/h3Rd8DHs9h6fXulIrKylAIuM75IumPCl8
LkOJikhMPYbQWcwI0CMzS4qvixu03wLGiNg37M33t+1Esb+bs8Mt49JclcK3
sEm/HCU9GXWDi5gUZ9ABVwcytlYhBw3fkRh8RGqA2WgMX1RAz431AVW0m/Xl
o9KtAODZ16aIK0ZsYxe/9WetYcBydXy84HjWXkO9DTwboeOXVmxfcbUnTyk2
ZDfBgzAwEMW3AbyZTXE4C+eCDgErT4Uql6xNQelbK7/yrET7II8KFLoTFkQk
B5Oznr0Ni+3tKdsOBO3QRXcRFus9xER+jI4UEf+Uzdm0xLkTA4lwwx4VHqUX
qQ9c+QcC0sjftK08PWHbmi8XUHInyp27RvGhYq77EZowcowwShOaZ7UXuKV4
cwyjCr1cjQeKXwzOkokj2QBKpotxx+e1RpHshx5enVtR1tkBjr0orFID7mAG
JaUBShAYdohFyXgfjXUmFGsWnbagauLkRPXya/ywcepjpsRsUvx/z92tq8dE
/e5ALeyN9W81Ya+KvUFkDLcaLHdOqH01+jdNe3uF3em1TsKawZP1/zsHJwjx
R5LKYMIj0L7gV+3dHr2xqakktIDc1EszTDtNbmJiBPGdgGZO5FXsvOXPAVpO
5up+Pp9sE1ppmOqaacBsIZIvfAVL9xttijz7yCzHpWmine3vsvKhdKhdrTl/
qySCaxo84fCr8s1Ua1CJkBKMcryA+KIcbrwETpfgOQAcoTJOjRvqvlJ82s0Q
w2OVpviwUFLGZUftFkp4Qr0LLbrB+9Uhuv+M8XkhANLtlbBXhfG5Ce+Qb0cK
YSMiD0/3kuswfK/sHjojNXckfPqC3mVi8GC/O0bvIgoEJLZvyTO2gOvNFpM7
DV2AlxAbV209XCaqWLSMMp9+xnKyrrgeQJMC6VkskdzKaY3Smenj1oqAh+aO
GVYIrw0YdU3fMQuhyIeTyjNPm/MnmwrYXowxuLQl5S6W3mxefOf58Q/tkSSg
d/1kPv6g8Xy9fpw9Z/vYSXYixyTSQ3usK80II9B4CqOJIQT1RNDbwanJp70a
06n9Qg4EFAyYA4Zk0qa0Eefrrv33BfxGkPiuhFAkLSbGVSp0RWqGIwc/JueI
KAH4VsT1POSKw8BT0SrS5/0sBuIsN8xci5mxn95FSagVNgg4ddP9RayxiyJg
d4jh6xx0EYGwB8P7YJuUAV0GgbgHrW7aYlWBIisQEYkSDcEEc5Y+LYv95/dv
ZiGCtSX+kuzXQfSmN/cy8C3OtS5BPx7vquDiZMezcpu4dli89/wQRoKy8cSd
6DJDFxim2cGHsfI4h4WkTw1wQv25tIWTWeGUX26W3XnG+X+fMNB5Uj2z8FSM
PC0AGS7oH5tGSE12scLzwySAGBNsHxgGSZR5ymu2dWPcjVcmiTh5zK2igMVu
ou40UCDtmbkxoo+0olhsELq+sD9A4KOq9ufRHVQv7xbw5FT3AF4ojG4a62Q6
C4oghTyt2WVUOYCMV+m1s5lfcNuIeIhnRfRb6UWaymEfK5PyhdQB+TCF/Jkw
GiTnI7KZ8q2udBVPfj6IrGPFRG4hGGBQTg1MIhRC6o00uCar42pxCZ0DGzyO
bCZQPh25dyo4sX1AusvGAeFjA6SJvwjtungaohGVGfcH+itzCfNJG4bs0OH/
tTSxSwLdaNdWFtB5zwr6XVGj18B3FSWqVOyd1g5GcPyj4PdDviGThQePDICv
JaWsMuPlzY9pUQxEytcUbA9VEO/xCchGoXlTvZO5FlYB+0DPyjE7ZFmg+e/D
yq4qMM1qZvMQHvqTCX/cHUi9GyqZX/pBNPeklcWZYi+mXklsTyp5J2BgkocY
GiwaOoPFXCyOOd7zkA/qzp3v81spZdR5vQyj0tc/KSsb48srzqYRsNW6kJIu
2HepEu3uhXgWg7Wf4g61ahVjZ7NthDoaFVE7AZUWf8J7WQVnUTh7XoInV0bY
gwlYxSqagABjSNRVZdvz9rADk6MQQqNknCByqauzjxbjVzVth+kHJD6mgQ4B
5AzjWlW50QTEYhw9xSzLSeiXHDFmy6QNuBtnCElqe9DOFPuhdtnYfyzz5eVU
Jm6UXsD/J0TbsRE0RapGhWoCNb7cwfGSJ+2LWNYbzQbtYQEa9mjfcbeh7N3x
zDwmKDM/fo042rbVQSabrSMkqooQiUkMMt5mdQEKCEU/xsM14Z9nvwUP01W9
zUPCvDShPl+TKivMQm0a/ug2AEhU22seaMQNnWopcZU/lk76C0cdMFHiEqC5
5Kh53NrPSyi2va8zPsbTmpvZ5rtv/7NJ2j3uHNzQXk4O+TpUtYr3L9FgYBYL
aGRZdQEDhz91o1dg+5Ne2mz0Gkv0qb27KX3Q7XlM/7H/wcx9SbTCoj7qeoUn
HR3hfKfWB8n2Un4l4Z+FP5ezkjCuQjN848+gWbslm4j8yf3Zpn2vduYtCKv3
8oeUHQ47Zdi1vzf0+y/Rx8I0wzZME+WkTn9d8iaZT9vJvCZesDobplmfn7vN
5L2G/MclZmoZ2kY0uMIeQQjdzDt6VJRW7Uk6V8KWXE4ozqZ+LUg63zW3vWkk
vx05CenvAU9GpH6ADX6bDhsY2pclA+oCwzZvnVIfXqDK4X3Ny8GukUQ0wYQF
uwAWqL+XAau4HYn5C7EiKxRixMDYp7Lo+0Du1OMLlJIC9TOkBDvXAD9NOkg+
RJOKn9JDXI5IeKhlkP4p/DudhpPiilDDNhXMdKh1F09Wo+3kw9d8K059JbF1
tEOsmXt31p4HDJiNVo+DSxE5YRoCa4NyScVrDziuWpmwNGpibIcdRnuyFzB6
4eXVBkbYMe7tFiWntWMzqz7KmlBqh+pawL+DzFjBQ5/KZAAHMlGA3gB36itI
V7Pu7kLBTzCpCYeyh4IahN/36/ZBWhOvX6KieD8CG8fN8cCx1Im229JFCZmb
4u2SEbsfYxyVOEYfA8Yye5HSvG6Ix6SZEh7FakDVK4sc0WZaGqCTymYVEbCh
Z8nx5u/kDnIO7+Sj5p7HRWWVrsn4go1anp0piYFqbHuCZl6zms5XXBg13HUQ
RZepDRgupy7BHY1GP3Sx2DGRnSc+kJkSlhbhRf8YhqCF2ClahL0qRs4sZnal
gB2T7CZOpgSrOV/Onjc6gSqSChD7GD0o6YQFKzUR0GC2Crwgf60W9PzTe67o
1voQ++mgztuGtwc/VDyed/X8GQjgonyfWXeaG1TFQ6bBoTC7LtfmgGVooVkq
I9QdbxDX+v8fYuD+AGj9m1GX7Sf6BagetvPP06XX3bS8Z61HqBiDkAWMG4MP
1WuZV3S5EwvSSDEDTu49uemhdSxNleSgGeY1avFRj03Zvo8uakaBj8Dd7IZG
sDv15T3cCOey8rS0GdDvwCP3PQYSkbQjzg7c3pa28DZe56jrzLrZxxTRKc9t
xbUfJyLn3DcYzXKqzjNWJc2dskjuGjCwTrVJ1nBZ29WeJ1jwiUZHaU4sYzsm
OXSvwmoIqMUm6qQQBZTDeK/Bc3yBvoN2BVbAXek2ec++r4uUfKIyvNJ4ilDl
VxbpqSh+34+6Lr0po4JJzcWEyJdNmCtNee0W3tqF6gIo4X0NqgKhPF30mj5g
LMMf/tj8Zy9xRQDEJMB67GOG0fkMalBfXXmOPuaEGkcF/zoPsJtM+B1nbbZ0
hE7nrq42MM0TwsiNGrVW3UDYa00rKpM/UjZ/S3hOHrC4iTQ/wn2jGK81oWHd
hrMGCHBsFZ6Y6tuPhx6e+A66+4bb6xmawAQrqkZ1WwQanRlCO1a+5fkXZ9AF
zNVCovktqKEpCEn7Ii7yqM+UsZRi9znnO1adrVQ7vU8pxPw8SdFf6h6ztU14
xJhhCWbDIRPgnKuIpV4mwy6o4Q9MAdbpEPY1rMH+H5ZC4rIr8PTQCeDJ5VqA
pfA0/bBGb6Hu/Ow5h8iNtNNVEb8aQD1O7MIlNerHs0kV7H8XW05NMci70a+W
wF+qQX4As/1VTeu+S77OuFhFbWN2wuUFPeTB0fP2bMkmEEILa6cIzj+K5GnC
ymuVtFNMvQZns11+ECjrOlR9mFyu1SwwfL/wzjBgLp+kAgJDEvZ/jlU6ncmn
WMKclaqls2OnO/WZ0ed/xHbNSoApAqyOOpLu3twVJlJqIBSefXTV8lr1wNU8
sjE37RX2lY5kgbTkrdjHfaGGGLzs13EkEX5h5C5iz4me21Xhp7oO7uMZCT3f
QBja4ZHXVafVWm/qLpUH8CyCVLpWo++NBsD2Gk8v29aT6hlOwy7YQW/wWqQN
fRKm7kqWrsMrGVquxxKusrY7ZiuhlB6nlfupPyNWE2xcmuPISZ3xKtJCs7a6
qpqZSudMyIpVYEWfIfugkgxui8dNQRetuzz/QVMcuNxHjZfBXD5umZ7aRlJ5
eNj7xL544czkUDGM0ovbx6wwuJiHIf6Ti5maOQvnWfXhDFLN/pQVgWS8t/Pm
sLJHbW5/vrEsi/ghNW401FiHJEISJQCDiwBPzpuBDRFST0x/0TtYOo0nejWI
fgd9bNZDy+u1pQ+Lia+bPkJVm4UDwcKVHmbgOG78FNj0aK9XUZaoYqfnFYCh
tirLxx2s2lxUFz1ziY4iui1ljaBq+1SO7Tidut4UkpFaEAtgWbJCGG97jeuk
gRU22BmFvrM/yGl14LJfTT8IVVMRp6syd7vIZTpAnedxu/b5VdMwz/x/QbQd
D5QouEri/+mIsD2uKxLxqRmWPYTpVkOHI48tKGLCqt5vMtcsCqNVrwgll2KL
J+p68a4kQQD1SbvWL9TNrz6/W6SPii0oY1zlqruzx4QWJ1Che31hvEUCMLXI
6zw1Qli5+z6HQmdkCxROo/1n0K6au6fnPSYdg2CoKbHamdMkvGhh4s4y1GvV
D0wdan8ubyG4mULn090aIbGIf9vi1ewPCv6dxL7KKnQw4646Ij5wI8VBlsMq
oFYHGnSd6NDQKdOA6FOb4v4XtIBh+3VfMoDpeETvetSAj4BKK7CEIe5u2TCn
F+YTJoi3D4O3hlL/LY+oe2KKmflRLyGsjc2TaY0rRKMz6o+aAjxYHGjIq3ca
5Rq+fksbIhZUiP3Ok1p4CMjCH8B8hAHdXPGcW/f1NLq//0z5ueS1UZ7HH3i1
ty7m1PyyD27+sKM0aQkdGry5bbL/IhnItNKUJtVZCoE+Gwxc56zqsm6MHAiI
+OaKQUknRIKc8V5d3pIXxOM1lKVUS/MwHHMCtJDQUlNxP0PUllkBkt0XKlT0
DrlDQiPIVn60ezuSN++xCiP9++MBZrrGtRfHXUnKJh55r96rIuu71klSdQoR
KucmnV/jmXmIwoSWv54fDi3FW776Y9YRpX2ug/s8CuZihJwpwT+lSoAD27/a
jkDGrnc8aZWhagy+i7i7GMOyjWqKWLaWlXWz/z/4SN5YnQxO0ezR49ZtXRJG
meiYPeLr23ofJyWHXDNcuUkhlIecIvETM2HM0SgtTqAW+wQQFd5ERSPu/QLn
rVHahNSl8Ka82vf4eD9GyOoaHGygqr+qIZLXWv5AfJAoPquKfZs0wH6tCMga
y++U72Iy63FXnYryKo/zb06EXtF+HRvNnEphM7gBs9nOdYns0l2PZdpvv/Ec
EzR+kF7soPl6U2KPxGNeBmal/Dw5mEdgL/6QSf76SiGyI7YWSCwg3Y8Quo1c
O8tal4c/LytC+ntVtAQUSSi5I8vHOUORrch2oIgVZwA86AE4/icX6nHqrpvs
NyOIOt1x1r1KbNxfbzrj15KZtlCAaGhSTu8MuFhLaLoID5AAVcIiH7e0jT2k
jY/jijCDgy0qQt/CTzH08SJn9z9QPRjVdOQ2z9bk++3NLTD/4bovbslqCTnM
7itX89znnNutuJlmYa5SSQJ47e/ppbfi1VfKzJO7+uQxUESXv5qQSCVO22cv
ncZW9dh5S3THNvLqekUis/+YFhg2X0YWYhWi8BwjvygvfoxoeahQGehCcBS+
y3E3A0StXxmgUdvF9ZlMl27jfTZhp9JsM3QHW1PH3+SmsjirC0I4XRTTEJnl
brkyX0rqpAP9d5qDbtt9asWNIrId854j9f38KfUvfJbttWJRyyI8M3vNqZjb
3iddMTpbQ6npUPCrTNvt3zCd71uZ7CuKaRHbYv2T3BAXsRCXsqEDJNtwWinH
6+lbd5wj87flfb+yjcyX1ymUQq0Vi550LO2krrz1McG8fsAlLFZaGLwYcpXv
4P5tjm/gxp+5qUh86BERzCjvdeikKHxApbrqt1q0dWI1/wEHj11oS02UJLkB
j/YjOFWZE/A9FWCUbwkkB3xoykBE3//YHCEiQLbGw+eNZJnCcLRtmRw21Ow3
vSHM4YQRqIYCHCXibOlm10relYrtLBAaJvO6GOHXuorf9ZrOOqhQD+5KFr8l
vASIoT9jn8zfjf1Wkrwxv1UWFM06U6VArnGTnnY/2+RbWEHrUyrgu68/bHRZ
dAQ8Z1ih+eTbGr1wz36TqD33gdZzZzW4a7cNHIn7Z/+ISgidxRMsSGPRqxEY
ebz7AG3dyxxFIFJgt8pcItkHxArcqPD+/q+59sNCAohnGa83laUV+dFduVZL
L3syY+6qjaANziA7oXrFZmGKgFV0bKGpfp2j6taa0WTGcFn3N6gnmp0HChq0
idddmLP4zENJQXi1gXX/3x8VoOHmszdW2yU2BsYeRdFxzu+OvGPREleFCLlr
M9AEaR/pJwDlfk1EKwMaGK66+yudEyGkEDO3VLRi8JUIyI9WzH/FgB3UpzpY
YmbEJkp89VYZY9wvOMZb9IZ8YyqxCNOPH441w2gsQI2bHSiYDbQ5+29W9dHe
2ASsBwKbddAOShRc1W8gHzo+K+1sMqISXytal+Z4Tk4diirPieXeeR9Kl2MP
PKQfNNWNZmpIGXYIOd1JP+W3itP8aMDfmtG+oeIprVn4cZ1TxNDnrd99kPNr
TTM16ggy9cPrsTApBXqsYRmkG4cwGm17UlpSyGxLlvsUaECCWs2zYkRHsEfi
RU0JIkSW3N0xGovGLs0JOHwFWo1LqUY11pMLVzC+tG9slnkniOI95/0b5PO1
MyN6yAPhNNh0+r1yr/e+Pgp/hO8F/h1jXbYSmc1vdYwXYce6QhdftdynFZ+L
JsINaI6MJMZa4mttexrW2LIZQnfpaea8PrXtMDyEfCkpBCBQBhhOmC2PuyxZ
cUAlooNJLvofai9Rq9AXKLMA5EGzXSA9sU88YXVhFDfJNjSgqElprhRMHQ3l
KNtXex7pJFssr6MB0BV2AHwoTMMaGbvk/9c3zF9hNxSW+V4K2hs/Pbi9WO8+
jwpLla4jVAApl0vOKgzzz+elGbNbKm24R3f/ZTk52YPGwGhYDCmnEgc3/zUN
UHyxRUqpz2IfQ0qsDzwLKjbbPYA1jQHd1DUVj8kacLbUFdpmHTizdiiZaC3d
7/stF257tOrXSqmSaFEMD31NwK/wDGSxHopNcrqP6sCmLmzKN8kRWP0i4xXT
/fYqxuTP4Wyjzsr2xakjO3pnjA1oqmQ2RTN9nyCfxLjQOpGbfESHbGXkYcYL
rUOPsvqgo4u8ysswSEUGYepb82+AvTjUAkui9CcMv16C7knDD45zfZ3eRtbP
kiM8WaVaUuIRo2AXe3VEGGG+CxihQSEVXJ13M9gTMo6ArXdYP87P0abLyDk3
qpVkzFtljWA9IOl5mO4am9DlM2J5NRoEejsCcwV1ls6JRB83o3vRkdz1XXmC
3Qcx2kjHbgFDvdxsKBu/3gqn1LXHhUNBmhS3Yx+Z7yzu4XUDGPvpBj26I2ws
G327zFCbRpIl0WoreEVgRe0UGsIzpT/nNT/O2Xb+by9L6hMsYa+o3/LXGrHG
a2/JRVUjz9PFVrj0hQoXRZ4lBrVfyahzObDeyM0KG0D/b4zlg/ckHqw1jnIo
DMv82wfWCDiFRpnREW/KAJo0qu/Uo1KKLrbXPJlCeayikKkae3wpjtUE/zjJ
659sgXL+raHpAk7isI4XC8wL3CUSp+ZqF2SnLlXdQKLERCrHBDoZ5Lg935Zn
NNJ93D1qZXcJo13VCe14ALqfxVqtqIgXkHS6OS2x3p11PRIskF2BD97vqIf5
rz/fKf1eJjkwHh8NELIAJ+HAbeUf83GzEudWdv+m6h6Hfdr/RaewEg9pR7CT
4AlpkIdq6uBYAMed0wzs5+y/A89XjH9VWUASEmLHcyJfTNokkUOu6OITJ/Ce
nKD1VPa+SKWhaf0Aoeg+7QfgAsw4sS9k23gCQl9OaqBk67JtHdANnxO4CAHz
8DmH0e2YU6kBFdZMUd7ttPcfjU3Gu0CdnaxhWtXAcdT1SRg+rqEhpXEAc92U
0GaXPWYY4C8+lKaC1aToRcAKNNZziNBpi6i8fKzfeAyffwUwNoEaguyC26vB
XjP0skiBW25HlRDz2McrXPtHjojrHPrPX3/zZJeBdQBFAWKxQiBklqNjGcdj
GZPMR1QcxtgkXsqm7oGnL9p5TXu0s4EFJbQ2bWYj7HUJSLd31c8xc9qGut3A
aZ6IbYc7WyrlRNGpwShpHCocUst6Sff/bPezhg4W/ZLqLHgcfBARu6OLGu4q
UeZPsD4a/f4ubmx28cZhyQQGtz4T4Nqv5mrt3OnO9B7wNOo1WgD5ShyOxC+k
K16eLQXIoieQwjFV/Gu4kASp3bqib3jhuUSoo+39uPZLtt/FR9Su0yXhWxSk
4+Pi/6oStXpzdZKAn3FH+3zQ9UXCbOiJ+/CnXfREh4DvU6t0JG7FvsCn8Ssj
kGtBsdAf5AL+ML66SlwXE/CUDzd22eCVDPfIrEte03d7+IQndLnou179ABmS
TaHsBfY7Z9AUyqocQn5leV3UUrmnYxhv7mgcgQA1jjZLoXYG238So4w0Vluk
aNKkDo0iG9wAymZyMVBiRhXg2rLD9sJkGU37j8OXR8+HUAVKhZqOj0wV8rrz
GYwNJCMeFAehprZB4i78YH5Oh6q2/OrOqRfK/HEYSwluTjv9jisl+QT0Amb7
NQ3jFUJ3tbYgDQ8jdBuHnh8jFDPnn5fUJk4MmNyDGUcus3O29xU8TwFt91ui
MWnbN8ke7YRw3vWMF8MwdR40m9rarJJNQyd7SvtWVavE/6Y3/Bga2Ti3wUjJ
YuYTwPL648yUGU/b3Y+HyWwX+TYRIZAfppd1E0jPgoDp08jhb/i3WO9jOJ9v
ae52UU0jA6ZuyWJePSxe6JTz8mzYdtFsfzg76Dv+dwpzHlUFWIS1x0aoAjPe
+TN+A/yDRtQ2libKi0UkPKhGzRGcn0Sgmm1YQBRJotFjuFTWO4vrCqEkfigG
OuCPuWj5ftbm9oE5+wwhO2/XpFEwE8GMlonP9X5X53a3Pfzz/USgBZweEN5N
uJ2WDo2gASEdyrFFujzmhJJS6Qp2A3aVv6QBH8hmtwxUoWyqgO/tPuVLiBB8
IPrms2lhuihIMNZoXqduqKpGRxKMHKPip2aBce1WA0OnUn8le4r7K2BQ7RW+
/INHRf3D7WOTwILMtINI/gNU0Jg01X4mUXLSO/dCjbJVQnNc/pYAm3mnPpaR
DLWcnxuUbifUHI+GbO7PmRTn8D0oTDIJXVjJF6CA/yEAfz28mM4Y9eOChlks
ycsEnMYitcKq1o6MgFKz4HbmJfdvZ7a81RkGKNMhUoLabPDi8D2o+GLu1OoU
Q66rae2OjJcBpTt6B2lq6EscbyL5E+cohdj/kanj0b+2+DotQWlZ98TO4lla
h193l1Md2fq0Wr1EyaqxOdr4qXrlVqlgiv21SGwd6db+LBPaW/J+mq8U4G+K
e2z9PXuhJaenuUOUnmlnnAdgR1jKfvF3l4T2E6XUNA17VbbBiPNRhgukn2lw
wDJVA3t6W/H92r6NXHNaFt85OUga59UPWfPJ0Rh6y+oRod/YX59Lme03cLrO
D084PCp3pD/IZExKNHchDJKmm9uQbHKnWtCSGDslcPiLu6TZosMSSGrUKFff
9Jv64hEjp614cdvKQ4Cu/C0KuKfepAYn0NU9ixRBmXjiDaUS2WcLMvFoHZLY
n6sCr/MRdLGQKCzkpFFNOyTYgzgrY+pUvHEYXX3JFfDh6uIErd9RIv/d/KXI
2ued6JdbJ91x67J+baHXIghbavZpR2UAJmCRjcdWb20Ue0u30leiUs5H8WmR
/qknzPLurUJufc086GxSrFVKOPvWf9T10Opu7jiA3H67/9hLJDyvKyFv8+x6
icUumQzhdnxvJZsMs9Q6pbjSic5HdOQ8Nf7MEQndcQrWvPqDVW1MyOBCJqdn
HpbRjO28tMpFX98XwLAS8mDJRDv6Ac3qh2xzQz0R51jmJ1mG/rnrdGukpe1m
Zq8X6/KYUxK6EzKFO7m5QVBtARUkmFFxt9UEq0/U2KoqM0RSGwy+Fwoyktq1
XwwJj2R7oDrFfj7g8CrqDRf9HkciGv3j5MjkIjZbktsgx7Sp5knF9b0XhIRt
hzqti9+jgZYNovp05W6A2367q48Yhk4TmSZtrZ2qo5Xn2EsE8WJZhcg5njTp
mn8korCy/OIM6JcKD+NpdpecHxhAqZ2MgdUnIJ7R/I27is6DtdpI/g5Akkm8
IfVugJYz8aecwX0YOZ3LindEA34KsFCOttDBJ/IvFs8RFUcNCdJwB+4dwzoj
I258jfrFYVS78RNa6xm/hCeyW8BVx2GGnERViRCiXju3OGowLQqi4X5P21xS
28wCTxg1YaIj/rK7cAFrw6YttUoMZXwXpBMV7Zj9dWKy2fHtUF+yoArSyPjr
ytxJd7I0aeEkhEKefuHtmZTqk948akavXesag8ldU2hwVG0G4p4eLBn1q2sU
7l203F20UsOy10TpqoHnXbpi4eBJE2IytBL37CNS1QwlkWWe9KMAwShpcQba
GKrC6iSnzH0RfFLf/snHe4LTyo1EX7w8SsJ3ohfFH7Az+WPs1PhZ+DREhXle
tl0qbqjuR5Au19/Fd058Fdnxvbm4Org6mO5vPwM0VJZ+dbdzVzIUx59YuFAm
bJj3HXCRd8ldjFOiUjC7LtA3dq0nlchMS820z84ZJBfxSRWqz429P/+RvTmw
NeDpH2K9RPU6ofnZJKTdo9b7KAMqkKZrHoABy554xK3x54uVRhiSQWlFCEI/
N3rnW7fStz7Gygr6fFd4noVavDoli+Fy9J4/Mu80IQnOxoazsaNJOz1WhXi2
lgfL6B6edIeP9ksxJIw5auPoASLTx8dBIDPYDT1tz3fX2nyuBeOSuNaVa9Ep
DOx/hV+zsVUzvY4wnswCD8uYq0c4iEhWIO4uh6eVPxbjBbs1chCjHjoGizey
9Zc+fvn+A4rdupGdZGTzlRSeA4SQVl/LjfteVq4tvGpViy1rsmoU1kl8r95f
s1GV9NDG0t8KfTvSUuZQFY+ou1osdkQ2hdNSX+/QMM3KyQ6koIhuypbMXqVK
Q60rZplOwSTDavoQEt50HjoIzjebJLTysiiWLX34lYMldrotDYeKE2MbCaHN
5jOmALdSVg769XGyMUPd+hyJ6m6Fef7/1Rgnjt+uPjQ0m6X5OIWMrge0FPw3
KWms2BpQVtc6s0FrbfuA7EmMzRHO74yCvPojOjdppfItKDjgiBhFSYXra21k
tM82O3OKsZ3i8/Wquux+kA/kzSVTX1i2P7fn6IDHkQdiyfc3+K9INfxHn7GB
xYiPBkNvU+gbTR4b0BJIU56yGRn8QKByRNva3rbK5bD+5LKaAzkxZbfBjrIZ
BdRKL/LWbumb6fSZkgq/go47vX+E6nCwCZnvUpfHBZTcQrNWF7tmOv31wQkj
WWLqxW0OeOyS8KVWhNG6EfUORqa5q/vK5qxo9LBZ+8cFh7c7r6cJasEuZF1R
mCXNedFGvwcngYDgGX+qC5hZllkwJXFolbk3QjOHoGUnQgwFQVlpZKQ4W2qk
A9bgJkUnewGfxEGQYVR2Bi5pUlpTF5sedDTwLJFaQvRnSGdDLFZ3MkaoLZKF
XUVCfthAsy6eg6sQh+UIWzgD/6AClquMDXU181WnqI/TTvLPw4XDCpzo558y
9b6ngkB8MyzopNh26WXQo09bAoQxsSvT99neiB8yPXDzkwi8wR3V3DibKLCU
Bvh1bTFA1M/i68U8LaPh7YOUgpU7CMa1LviMon0+gNjeefAJBct/BVrW2xpP
B7pi8DaWK5cECA7hqM6Hp/Tkz8P2RPxjadJXv5N7ofHInuVGccH3sM8HotsT
dQDuSYd636VrgpfrtYwnu4uYHFYsjkIp+LyGbAyraXFwXsKfgLUnd7nULS51
l8jiaK+Skw7nOUFeR8bgtrWY4tMkaw7VVrka78rxkNKzYZZW8rsqBBbW8/r9
pwnL7ovI1Lu1dtJjT4YmtMjTTkkp65pgAIJ5vmgO8asjhxgSTIWoP202MRq3
QCIXUK0AyqN9AXq/uqISIo/RmCoY+Q8LpmPI/IZBCEtEeAjLZ+10eZrh1jaa
ATiAOCF8bnX8KGyPNHbTmeloQ43YjBwKR5O/JVJH3hadD4LYB0FCxN/uezS4
j/FbhxGhYn91aFfISsX/JOBsTr9cvkG60ffKwixDobPjjoXUqIzIKEkxmD+e
NdqPczGGHEw1hLc9fGCf2d1zVtCDfTjNwdN62oyeXpl1OZSvC+qX6TK+3Q+f
CBUkrPeSRW8Mtk4JMgIUjxRVPntMikiKuEEl6OYLcEmvStqxaX6Be/fYZN52
qJIznqMxZuff5NSMw7kp9o8oov4ZdBuIVEH4Gvh/+QcmCLc55Rk7zD1idWLq
SdiAvh9o+4qyZ5V3Sh41NXEusVFGjDscqJHxHAd0B/r23pCMMa7cWIEfJwgn
G93iobWsj60G7ewt68trqy93PkHV76PHPhg3giw9rseXdDSG9vSRltfMpFwr
V89OEyfx4/ZURH2tIOAMoYag1skzodG5gdrr1shosC2mqALF7oyQMj6f2V8Z
97mf5shGOuWyvb8YeubJGQkLDqzdF4viOGxQD8ITMwLbvgCTHm47JJfssUEW
/ReRDbJB91dmyzxAjI3UUT0XmTIRx9KP3SJKHDa/H6ZhePh+fGHpQVfdUzg3
wEbARBUaD6ur6TxcuEOGvJpNqvCLNrLbpMsqm6NPrbWjWpSUt9Cqv0+OEK7N
DTR7nXSdpVM3TGhlu8/gdsLdQeDC8guzpJRXY1w8w6zZEiG+wmX7yI+ss4nq
UMluT9vaxfx54Dmmj9b/o8hNshoKEQPM7NAZyBKDJ+c5Bqkh4NutKeUpAg88
QpgSp+Lz0l6hSuWsywQGI6pzRMiIzf3wv2Tfm9kNslqbeDbeqBXtyo/t0DjW
+C49FsB1jAEjH2tDyQp+FSqlBBE+SWWRg62QoWcZPK3QxbGOGJzlk4lhq3gM
NZRmZl3DYG+wGn5GN3RqHrNDLiOvLfVM0ChORzqRaNu/hraeaO+BqCSAd9oe
MesrAKJJZPJaw8dSr+Bf70FmfeHtluShL9uY+NnImZdyDhpAtteyKH7Uedez
/iYrxEbc9lt3jTZDX6wGno7/wZ/CGdvq6ocrcScJM10dMPhHpaDLSzZJr1Iy
LfpOYsaCKM0Avq8Bkxy4tGbxaqzLSAio/AwqGnU4ZYN1KHOD7z5ezHFJXzTZ
Whljh3PzY9jD05SMIPpDifIbqtNXItDBlL5lgxbD3VwJRTdvlVx16uK2wb4U
MKztSt4M6jNWKiWdNodkVroW9bc4dvlikci0oyzH8L0C9Z9rDKvNfr1RZptv
ATgpfAqgNZQkC+QBlC/WsIQ7wi2y44Yq3s7+Z/QzcU32A35AgI2S+iU90CZw
kr60u+6AlO+pt5zZ8cTJzwtXTNlzyetVY8huyxkSsU7c948u6xxBnOXWYYRx
Fxx5KbjKe/V/F68s1Z4o7xOCtzEQjmsZsEaWYMxekpSLFqpk0su2u+LfL3oW
mAOK8/vEjKECRqEF5AJmIR/XT+RJCxQxiMRAjWcztz2/TwK2bD79diftdGFh
sCo/18mYU3bb/P7wsg78WLM2VCd1QMVhUjy2MBVjzI+dF8pksFWrBUHsEVf1
EQUizBpA0UOL22G6MUoks8syUNtOGYpW2ql4XegGLGUwWONJYLxywcFgFrfU
EBkKsV24boKfEncD3bYfBl5nlcwA9i/slu/sSIMhy0C1qSHDAdYK/HVitD6C
f7DAnvdCn/7tmUDxBDzErJuNloSLUnbECOSpYJ/73avsO3wrh6cZmJl2zLoy
hKjZDWXNpnarBBncq1DUjOEpkrdZVmCKFUUvINE8aE3e1ky68o+WfAyLl2Ej
nz9dTPuh7OopRckx9hnKkq8ogwd/31FW1WKRLrRLI51kw/EWpSh1Y7FQBuwa
+pNFCQPKqR4CUCYGAkfb7s7MfMGXKaymg889pBn7dEEY2y+S5rGh5dSFo82t
5YoC384SPgW4kSM9uNQG75kkby2u/Tajoky3dJlY1qQ87EJZLYcwHkyfqy4a
3KywuD6NI20aTXG5/xSX0Dar/fVzMcsXfiORCo12eks7jny27u4jsj0rA4FR
aIC3sQ/pAx4hH2jXMf6XnorC37wtb/cbNYMeFkkR58fx82JKJ9xF02XJhME9
5IV+JQhZn3AJMUm6STPE/mJol2VVoMtg5J2FqRSduVINyOOciybiouMLVY3r
izLceWyoMzMKPPuyHFt8AffYK1chkln0AFePKA4P/18B233pWpbiIChIGWkw
S969BS6QxoHiG0lJuOF7PCx8rf2w9eHaRssdoXHiUfA+NuWo1XwznJyfB48n
V+0Ne3uMsSpTD5/y4RQEQjRBR9ZByZ/J6CtDpzttvzG5WfPP3e/UpB1hhKOE
WJL6AQxYlOluZy9T9PgEGTo0b8qZYSk0/re+0LlFgotSw0EjnipOy+4ipO9F
KxmtvXlWcRbxRf7+fe1VtBluIrf3MxRyPmqj7/qQZHKXjGJqabGU5Jm9jEFm
jYeVZwmbw5aPQ0pNzUoJ/urOvnnSwENWLgvvEHb5koATigPQo+yL7BI5NDja
sL5ubztXtfbPUCnK45qN7u5JISuUIFCRJj9iPZgccBpGY6Nb1h6p9aMT+Q3a
RkabHiD4p+UCb2I6fUPYDd5K2bxxwTp1BF67h27LO7NOI5SruS8lC3L3z49z
bK727dJ5LJfgKFLSE6FvW1jxj9Pmxee1AN96VCX2EcPRy0wNfQGrBQuQLx+Y
F1xK4ycdrSH0IAtCGKQdhcBom5hY3ObovvPQbhgVBsKvnkWxpHO0+va8VGQe
i82N2771NKKo3OtEXtCYwtI3Ern9RLlPnU2tH3LtkKxrJb3L5KA5yTz6vPbe
XFbPYXSy0/Qlon8rE5mBKbNmRMG91H3AWmQpy3PHvoYIlrPDoe0WjDViooPH
7Exs/vjjuhCmZBqdhbcKUAv0ZVz5JxvS7Se2EEnfgLC0nqgrJvCLM1usjMEg
c+d4kwILex/NKXWLlZESWhi0dW3CcDlEKRpcTZXl0UckkUHO/BcQrIqLVH7J
KV4YSnZIJ/R6Yt79d3hWN0o6d3itZqt5VOsbz5y91j998cy5Y4VmW1goc25l
LwDPaDDf6VXrHCRYLw35KZYgI/jmQ938YP4A6q8o8vhj43h8eKXHtRe3vnSC
IFUjgg0+DpXhA2Rr2j18hBbV8r7AwpffvsH4KVZKXzFs40ewuueMFEpFPGFY
NDxftbhIMGQiY6rM9ZR0CXdD1gMcJ5I8/9uSvI6h9q6Ws+JF5QRYODehReRC
DnvpQp6QrYMzC2IgBbKW+PlyOC4jkmqtrD5fQpZ4WcsDXaCpDfbuLHi8PMUR
3G1IB7+sBKsz4h55aqsuJ92rZ7NsKyI9Y9CGxrjcAhvPHVwIwRO9oHwuO4Z+
8Pd6BMty389P7rHTD8XEKwGfVdo81bHojd26lp+exeOectmbc0rwLpijjokp
7f5mvQM+8I5jQseiuhwrnekZZ7SVvVG+Ybt3uiKxU4kTnfgclsRZrIt84u0c
RYEQFsWtJPv0cbi4WxqG/kK8zqDGA1qNmsv00+jfFLmj80J7cJimnJNUzr3N
gwYk7MF/30pU9BYiZ+lGB9zf0AjNNHw3WjGYxGFCGjd0JC9LkpD0GGJMTEQB
2MTHk7hRsMOMXZOIvFTRbuL4Igbw8xW3un0b6bIv99R5HM/8yzcMQVAw

`pragma protect end_protected
