// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
IoOOUEqMW8v8/UZ/iXICqZsT9RllVGi+DRZT258PknstrxSiPJlNBOGCMTvuVUo9jfwSw+jtO8dE
w/0KBWOv/3QEE6Dl6m5EvMkfX2YuctEEN0Nqa84+vN/4FCf/X0pCnjuvX3E429O9oT9xwcASXEC/
8G4NWBnGIcnot9cIO0ODYY7xSk5MbzWUNseU5niOLq/xmVBJGbmyedAWwET6HwdniB2CYpxe5C2W
m3b7v2v0bQQ0Yma75PebjHgbsgC2n6dFX2uYHKngCAsr4T5wyPYIwN6rZzGtxxfMAW2bsLmoyYi3
GFktIj8WJZCHPFblp64Lv9Eutb969hkWsonorQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 59792)
Lmnr9Bf8gVtEtITR3f+MOuO+JClqUzmDcqkUJdBF1qINikOlIYa6wL81ycglfUOYpRZNg8UBzLis
5h8M4apnicLdE7FU3ru68q/PoQWO9pgi7fn2c8elExMPhZ60brvC4t3xkAXmlFrtHPeaiUYfULqz
XNmrQYQ6Od2Aq3jGbwRgwyaCeRyMKhsTLOlvow3fccUHCwJwk1N5P+7rgYmGjw0lCDrb8/+LmQlU
3/NeaqIR0Z0tCFBqOlsdsDVnzUD+g1v283rrTrK8jnhsr0T5EYXCyBaKxuqgcq7XZhE3fD6uqiHU
63kprh2Ygce/dIamnI1HO1fHlwjBNoYgHESSm84wFYUCygKtOwu3Syz4rQLplN8foG1mP2c6r+lG
eIPMOxcv7x1gmIvbYiXD7RntPV6R8X8+70thIMgoKOT/HT6yreH04E5DdoDRQQrTCM4MHG2hoIKJ
6xxdtLDMPZSviZcw4XgL0ee2jr1ycwE//wki6wtytY2mJprdt/+m15Kixiy+HEW8jXmcRH9Wvu83
Z7Lzc0ABEPUucI2mvlSks+JWyW6sqr28qhttaiaRDlLjNi/Hr6LwxTgnuiZfGpiABPHKtkUeZO8I
1kn8H2AvNLVkN4ewGjf5hrfRNtIM2Qjsol7IX1XbnU0slVY107h/ntN9WFw/7Oklw4r7twwZRxUj
7pF045AcoHLGVXFdHs/ToqcVLdCoUw0VZn6RBryJ3T+Jot+Mqn3KINaig7kRG/mlQcUm4Ivweyla
H61NNSGV76scUNogYnyl52rgJmaO6XPrKb/7il5sdKKUYuu2c8WKK3STCS1MBuxtTVh7vfbMsR3C
LtczZhcpVdLtFEmozPhgh7czfuSd0u/nPHoWPyiT+gFU2dVId9Cu4CfYU6UMT0L1RNQ1gv93WKJ6
sCEkpLrYiaU/njhGRyJwj5HPkKGFJR9PQLPqBlm6yrfsRNXkEvzMQSaKUAsXVWf6jX70IceloMzf
QodtNHaocfdkIZZnsZIatOS+mLQt6LdKlqvPxugRlVLdCet7Kzttn+ooJe6xWeZpZ+84AXx/FsdF
EGn/5xuJL8HAU5qIZ9K4v9flUewmdcotq7lLVQrexTwANPue2diO00agXiVTfiKu+IvG73+s8ezm
VWXqLHquYKLHBnHgEzP1xf0nx0NLhSJ0+vdk2Pd8tZVW9PSeJPgm7JVgNgIL+WA/Dg5z5MDGXmUj
wRRu7cRCEbRAz0h7fsGuMvmuktGbEueYgk/k1lXisjpDg4+8w/7ceao83ETzZZ0wfigriNm0oxPQ
/oFa74Ez9tgUFuTUSga8B7FNgwAg82roXYCxyuKBUldA9JJtyCx+Pmt4CaFp7Ms6VHxVb6f6dGnF
2C4phmfGnVn5LI0f5lYTjUF1TZXQH0Nm2JdX1c5ChtW3w7JHxNtWI0IIf5NDKTk2MwxSuvC2WDsk
F/DvEfIr+H5Hlv5Ck3LQ3QM7U8e5U4DtO7CTACCjK6P58n31jppvTLveBYCjGqzU9Gzlx57ilED1
dkQU1k8LyanJK/zzO/8YpMVU6MTylRJ//Y3tUlm4UqLtkXFEJ8jGsHPjq1qX8Dq9i4BLp9x7RXkj
f0eLPhfVhifPYG2jTUlUyN1IjHxtzVmyU2pMFFRC/1Mlwedq2Cek5uK0M9UcF/m3XiSOpBcg5SOF
c2g9yr6RVNyb1Jp+tS0mvJCawS5VmPRNZ4jdTuN3iUhLPfus7HFSYVZ8nBeaZ1NjZkiR+HbzI0h2
XpOw4TDjvnuptVW9I7/Pmrv4YxpDRK4h+MNRXWH7XqSwr0l3YVqxJhxy6V2R8L8NxWo3lZ1xmXuq
SQLOhtcib4BGsCqjNvHgwZhg+4xW5j50GAAFvsNbi4evZxeEVTkU5UMmcU8lkooSvBDteE5QT081
UDWorp2ntW+cIC0T63qcRLU44oOLm8vHe+IrYct5/AHeOodhtJavJ4zbO1s6gAk+nsZJT0eFTFsP
2+MbUrxKm16Ajw7TnvlSqk1rsyLKzwxpUuYLHmbr2Fzx7ijD4lufk9w6uNC0P4A34qibPECw9Kcp
NwXNYXBXiA8ze1idbxJgYK8StT7klLExtrVC184doDxqiWkQcJOlJZfXQs97dgR2BBR5N0qE4eQY
QHoMO8WF6I7qUZYsH1oeP+y1/Yk17NeZTgKNTj+SxhfyysEu5LthUIRIOL+vc1/ow5QuExLePVYU
/P0nEm1lszSUJpGBIL1Qzvmb8svXsEFomxCU0fgAuL7AzmtDVmBExrdllzwGtN9IInObDYKS5EUS
6m01Kut04Lql0awDHI5M12mCJB4z9FoiNupkW7v7NWg9tDRIEjeKsOre8IUS24sGSCpc4VWRDYg6
/pO14Jb7dJ3IfD+UkBvr1V3affOaWpwhC+AAiHe64Eio32VeSO4tNKqdNJUglKHSTzTan9S2gaw+
lGmZMxdHND94ERzqr7UF8OZtD2VJEBAUUm5aZ440sAxq8jZ9L0Bn21B3m4ex9unu0Pgpu+07IjED
e4y8G3wnKQPrEvsvBoUDj1V33epJ/5n580SIwsz4DNbBDL+Uykggf7VTpPbudxSbhAns4Z79DUMD
CgT2PNpQuJrZIaQ85NiRZJ9qZ/PlIgb4jBZ29oaTbPGvtB5hl/wLtT6msvmNRsDkxcGtGv3TGk9z
6cPbZPqQh0GLJb2QziNpEJV1ea88XwG+lsNOjkGPB5ZG4BZkt/HMSO6S+trLn3wBvfowcnqe/ERd
X7vmeX0GTC5H07S/tsP2YLw+hJXNcEQO9AKkDV6Yuionbh7BlvInyPjQvAf2nokUZb7gL10Pp2sZ
yxdQUwkeaOpzPvL02UOaQglHxbBaavavtU4mwrZO6cxNel/87v7irTHOs+2ILG5p7GZWUgRw/x8W
Ttv2UUN8Eg8ikB9nvnECaaUfns4rEM370R3SPKHK3gaRscXFUQcFVOjW1jbx3cm6nLt4BGl0fGgE
+6WCMLvEgPnfBGX9oDXjUsSeElyeMDz1IVZeZjQzkCDlJx8ZNKkS7fuAegKSOajr+b3XCT3LJ2SB
qAJ4x92njMgYMw7ojhXKT5Oy66zrebYAWBn0iqXwmw7hqUwaMV3nxSt4gp5CNVdwoawwiWklmbAK
SBLj7/M+kKC0QkHu6i34dvbY8eXWbnyueycc5RMmNUAmCCvGS2nR10X/j5Zr3NwBUzdLnCWoSuh8
FVqM47Hk7ZlkxotxoPoDF5J/mHXuooKeyRTFYOa+9+0UuDl+ShgdeCzWGE4jGrmjGs1+UY7JXSvI
/bST0WsLOKskF3q1DLEcUvAwbYdBbAjJHxj/uuhqRmwsrzDm+s+nlM4+OXxwjEee64H70/v1mBD7
NptgxSWcQtW+ojSS+kx9zVQphSp4hs34lzOC06WWhDrPbhKKquNhDqeqNtX4aRa73KzjeN4KiykM
zl8K9F62zjx3xPsmxDQdNsdZlj3FLjrYi7gRqcuv8llIdahHbI+fk97eC99KAC6lx6UbDRD5x9UO
tpgtoYloP9KGsuIKHdorjjd2NTXQjywJGOdY+iitSz1m5z+vUbFpvfG0CObiaFnzRChXu/nGDEKS
oiu9CY00HbrBg2Ki1r9o6wG18/ctDwMBMxDhakBrVXUapTY4vv+cGhBWe89yfUQ5S5zR/Qoxq//K
6++zMZY0n9CBuWlq9qgxE+dhMO6I/iQKDX48N36DOBNixeA5LFp1xnvbYxXVE6s/zF2mk94EkQiH
XWrGgGUI4sKyynq1OTogXQzGj2qwPaDMczaawJEmcWFh7i432bf1AElRB5d+pK5F/Uk3JrEvFez+
uXTsZVjaxe1RaRe6UnAJWYf/IbsEGFCzrrHyCG7+wi7wiG3y2S1NH0UZm+l5cBsKQiSZ96S+pWsN
OFfAXqX1qqS0lYGd1RWlwSP7J5qXF2TyeuGbTlqkCExMPc6PMjFQ8dkl8wNKXraRX/0hpefF6Fdl
GfQapO2i8sJgB87NsVZHCER8U1Pd2yr8W+Hhc6Qcy/aEndcmFaeayzjiu+qc/Nh0tJVwi9rWcdMR
rR+CY03BLw3yc/CnE/UJBibn5ZlGxHGIHu3MIefwowzCGpjGecE8D+KKdIKkehgKJELjMqxggw05
9SOOrhA8fo7id1pDEADvAbdRayUxZWt9bkSWkE1R+m7DelFn3eGy1V4pb/mhCmU4gXjlACngOQ8d
oVCD3eLA6z/miIPFv77EsUjcZMP/2QRF1L4Iv/TfsErrVL5zW1CDr0FrNlTS1MD6Jtx2ywoX2bAh
LW0xajlAXmoegl31duNJYQBNNj0uFUI/ZJQgjYrJdmTLx/a5H37dLQo4kp3hj6VMWzqxEwzuxTfu
ren09RFa2pdZUOAw5R3EqgWq6CSBYBvEf5bVmowbVYNd7JWBrkJnMwUWZAWVxUEt6Lb6p4H1h45O
KNcfY5Jz+lPqO8qvoJrJHbMXDuc5iTE2wHHe8/q62Qg0115EwZQcH5iMMQ+4leTAjKHdR9MbBWPw
QdiKexQ4JP2sX9Dh+W+ytyoDXakR+MQh6qXM3toP/QZfFONp++Hjht07ZuV6OteJ+0JHehWTwkDI
kg4Oc6dteFikf/Qw6K8c65o/o/CBNe8ESxUfSFVL6/b5U8v3hEX0ZRjqZSC2EK+7UZBDDfSJgrvB
KntyxG/EHwhgHZTtPXwckn8aVu1WL1csZMiK3s8kqtm/EBOqswIpofTno+zWL7MQbz5ktxvePic6
c9DRAzt/mSrRpYHIWAzoSvCjFjOeJbofkRJbcdJZ+LcVYFQ10ESDC06klS3BdFyvE9ea66XOnfVt
goQGxtFFBhjJikHsp7LsW8B1BiwxplIYUMWml2xK6tEXszbUa+E2GyXj+tkQH3WIj5euUohve8YU
jZb+eHfGemQmFe/GuUanhovxhls7hO6lvHkld1NVZN1jDaHaxjXGYuH9W3nsY8a0Jp435LdgVN3c
d5cfnJEIFk3JDKw9vEdGSuZAG7cA+Mx8Rhrd0Cz2RKs1gSdWgsg2yy0yiK+5aVBWrrHC3L0NF6wK
CScA4cgZhnIyogNbeHcvf6+s8xGkD8jophdPXaF/j7Ev0bY8NAOlg2+n/UiFGNmM6h++EBv73j44
cT/Vo/h7uOJ3nqY8s0EBcOP5UQFjQ0CPdkHKKcmvV9BI6MorJ1hbP8FDOza63VxI+6JUWCNgcwo4
uu6rfefVGw1vKybk5vUm5Xc80twq5jL0BHcrJHZp+lOhirLKIx7F6qm6TzSI/dF5A2VARWWyN0W7
fmPrET6lmfaHLG4PN27uwvD7obw13vxqJa4JT/3gp2XDTKFDBaNnZbw065GExmCXiZtcNffyG8Jn
tV//PSze0CR+hR+Xy12i61bsW1eCzcaHa3dd15vo/WjBuedioMA5Vs352YfQSqZeGOFkILNl7lml
zkkf1Ep3zLY0LbY22YuUr5fZzQI6YrGTCi2IRWI2ZNzJdpXDaCUfsqT2QmBvJt3MlUmfHIPYIqKT
db9ZQP1HfMeqNcLZI7JHQjcUPulFkmbuLk3/l7x6s7fOgKOt302emh3HkpvY4HIavEd7sLlJiWZZ
XEwf6r2UfQD8wTcL+TUXBC1kOxWgrNcir0v1SJgj0IsqlUjRsPdMY9xNHtcIdMTmUr+zJcMBfSK7
olIC4UuYmhUdrLQ32L42av/h8aUww4YPLfYEt7Mps2LPXpRhjhQRTHNm9BqQRrMjmnpBVC9vxlaq
TUeNGfNJ2z9AiVcQtqe3BTban9LQWeZcROB49z17cMUhaTst5pT5Qb4sfmbwnOcN2z8CTb1lVXIL
W3X6WPhhzhADJHsNu9dJc86kgm9yT4b+ubv/f9jURgW0RE5VPBV8gn5ZRS/7t1BA4Fm+xM7ZykIX
7f3E2qMlKJCor+p1qVPs7siaughd2kaW1qZ1G39v5bOoEGige3dJquaTamZ89MzMslW+DGSqLM0v
XSfCAhOvUdozgS0xZgz8N7WNGDwswXZoP9GKJjFLN4X4xRiUFNRcIviF+xxCZFKju8szYSreALvU
/yLTQdi6KU5eYbw7IhrkySz7wzGwGRSaEYEz6uYH4Rn8t1N8srMsZrviiJ+HR+R81Wf8jz3Dj1s5
X58Z3qQFnmuWeFFh+S0vmqbmdqSPaFQvQv+CFbXjuJMMgFK0dLxoIKpQf+GYK39tXCLPMM/dLjoY
x5gFcY8Xn8J8Y6xe3MHZG32pFi96v6TMOUwImNJK/m/oJhJFKUgBT6ptC9wQ+Gd5/gHZlqQ+B6xq
cZMfSYDvvo06uT0oWBePf27CsJ3iac+0JaDpDoD14GyV3P+UQUgI+1SScDu+Kwt2bRtG8YUrDtd6
vkU/5hdgiCeDDojfPh7e06/Sf7h6H+/NC+wiSvIIyjwNR82ACOVLwDnkHnpJ4Y/hDzTgI62FDxLf
YubeNLFow3X6LjykSed5mdW7xzAr6n2BEHMV60zfrxldacpQgiMQdyVPgroDQhUXe6GFWyxUYHxo
bHeUfq9NLSABhGKPp7tw5neWhKP8rc5iGXI9fgp2UEd+BEPiVnd9zPD1muZ3n/eHDSrERwJ2KXWz
csSzN5TYwYTlPRPYIv4vHULXFTHJPGEI8qe7JruSBmzDGzUklVzk3HOZKxpbTOo1595scLJUnb6D
0zEIQ0MN68ZCWu0QumFdkQX7X5D7PZ69DVyPM+8bBMVOgFlZEbrTDFiZwn0RzFJWqdJkZuU2tOyE
8f6Uy21gObCKzX2l8mnXahmLCKLZrSAWim8NrL9ewWK3HEPJQBg0tYYupBov9qfvRj7a5iF+OPP/
99ELfNnr19xqjmYxSU9C9vxCjKMKCYrh9bE0gUXfqBeRfNZNJY3/qax6S9r3lyn5zhtPQ6CV0k75
L8lV4gO4ROjWDnhP+L7JfgvGLOARWcUPA/+qjpNpEnpPDBRv0dNMwgfqdJ75qfwcW2hKpmYrlDhz
4Do5MaGgvLJBMnYPyp4qxffd+OJ6sKRh2eJfE0X/11u1ZykLTVLrJw4R5vOMYYLw3YZ4O5IZP+k3
++Me1nwdkEn0ZCh+qg4BMbS19g1bZDPunVDFXkvG9/dhDGw1IdvAmKYjheOVx1BKzVHKqMC4KPaM
oG6cw1aztoFoa7wNY5ngngiW9ZmmGP8WgmX2lq+2MFHLX/WmEn02tgeVjwtkI/oBSniX8gE5VoUR
FDu4AzIzXn5sG9dQtICv+kFTjUnR55Xqj5SsOzWgHwH+0AtzYJo6taasalQQuU5L+wJ3iPDG2faN
6xFXvJa/iag9ojearXR2vwO2vnL6R/TUdF7crfXww1oUySXQhMbDVENqoQn1ltidzOyPu69wQ/g/
LwTw4CExDtQHasNLDEZV41AGOT4ihEgl1146XbfvBj/4XYRrEFSLM4HqlyBzYzT1oX0S8uKv4kuX
R9T0gf10SYu0VTjJQ+QpW/YADd5hnVFWS6ShOgFcsYkJ7C5Yj5nsnAlipyDnIlrU+uC0uQnQQxpD
mu/LQ8EJAeI8V7J6JRUwElFItX15bvbfKLHwG8Nuib74So5yo5eagFv1Xrih2xAqvtYP65YjZTYd
bJQnQKN7IsuonwulyiWtDGiybLZr6CBBTJgjdRYpo40Pae5+A1RL50V8f4E3OVm/uMlW+OFuO8j5
h0PadGWEjV/YziHcPLAsuWnIt4Y0AVUighXyMLG7hNuaYLpEUV011wyApzHVQSz8wdPKg86qlysx
rrdiJ7oHgYRJaYO+vpmnE2Tn8M2ABuFUTRQX9HIxNu7WodyIwOxLW5byx3wJQKPG+egrxq2WEGQY
BL6uRTUttndxBM0nKB+MLi4wqy5+ICw5kUYDYnKZcjsF0k2zlxIk6+fBQhWpFlDY2MYYLHfWcsaa
LsaBEUFZdtxYE47aE0AzKL3VGpuZz+CBUjNNSvnx0Vs3JTt/In21gjPBDj7PIy+C6cOztf8RrFen
R5qn5aECqieiF0MkV04+P1q3awJXTkC8csKhAT23UYwWS/X3a/XFH7A/+7GCGMpYExXgiLeM0tFp
HDS8NkPPpN3FVIQo9Dh1WUf+aqV+vsJENOAiTA+z2hMFPvnxAAk/UuJsndPaq4LbFiXUpd1gdT15
7eMJAJ+uTmeyeX+aJO/uCvVO2XC6XruFISV1xDfgBZYcQO/UZodF0/O9PH0Jki55vT3LZpjFK56q
5oQz+lba0iF9YxNoeLcGRvCTv/iI9m8tFY3Op2sOJ4b86zPoPrQasipl0JImFSIG62vE1XeERFIk
w4z2JdKkAaPzN+v4GpQuRCY7EBbxxnw2l6rwxQKdMVFAe4huWuhbyc66CrRhG9v1kp8Wfj1XK9Yd
Ierd37VtO+gAW/S2APj6g/4TmYV3UGq+yoahQnBH2yWKmLS4PR55s5A8qFweZDse50A6X1eOBiQh
RLy5WvigN6pRSCPsooB1NZ6clPlJq2A1NxguchbhkZbrZ9I0LinlF43oc6qblKSigTT0mCK57Dws
7ZJAGNUn76W2VYFSqRPQUDRBfrjKNrtmGOImWV4Q/fzNOADA/D9FyN0z2HfKwbghGElRiDrUh4Tk
xf7xUtI+qE+XF2jbXrALedlmY5QZoh1xTrpKGcpQUdVZEPKuEoauoCYPnbJYMskOyLFX2PMXVK+c
IGi9nfE5pnviTqd7Ikv+rvgAG1R3C0n1c5gADt4r2cUIISi/n47Ok0erGT3MEMhoDYExHvtfP5o6
356c6laiZbTnStB2t/AVW6oZKY6iaFSOvJJhJK0Kz0xNOMoqy9w9TbGyB52fV+2oamZiQi8ZZRyr
8Ltpg6K0r+NkYmJ4VST7daARnlhPvnoqi9r7Fd1see3eTKWXpSxzFxB6o/b97Ana+z6EyGt0WeHR
k0bu0y1ynGbZqBLoQ5UvMrPKbU/QYzL/6Da+MuhhRwGyZLMxFAawNHH5q7v1uUquXtLDnl4q7qGf
jESIhjqNwFi65xSJ7NvuzZKqHmdeeyTZtnLWvyWrphOJ7NZY/4rfMBQT7s/KiaedQoONm5c3a2Ys
A4v351CFvdj6heQAokkbxBiRk7ErfWuZByhAcn3mBUFE3vtY20URgqtHIOyUPSk/68CYW3Nsf948
Qmo9QgQdBikzPDon8YIZcrIxwsXsBeKj3IFQr1ExVxYlryzzn2gnRhdQSbQDIHCpksc3BjLIYoXz
PNBK83nalDYXmUUxsSL/xcCejHYL8+kfB3urthXj8Mlfdg2P3XUuiPKjw3oCs0GyhRClwFQ9nl8y
0fzSsHQ5B1V077ygoQbKLPy46ek0XNOnPEgtsSsq/taskiWdGwbyYg6vYcrOUIf0C6AZqBXNJc6i
MBpE25xbtbLojeuxZcF3zCPNaWx1rtvOMLTz9kbawsUzBnqY+91Pmz5kqgGqFvLf1sq8zdrW555i
4zRGqZVytw89DobJXdDtIETCV39SulF/iv4fcsfQ2HnaWRWv6Cku+0mvoAqC88lViauZsksFI6z/
x3vtaSo+DKk9k0DQE60V7XQtTxvanauj8qtjpTyVP16Kid/zrdUsG9RKaMHRhGdzcwVFje0Dn1q0
F8RW1/itxFCfsMBmai/6JiEk+k2b980Ts+5Veydvu1BK15H6jVoW/uVxanidxL2FD7dVJI4Yphrr
otjAAMqZC1c7lVy+fCvVuUQTmALUpJzfYwPCyCVqwzotGYMQIR5aPgG9u1i7Cg8EisMEdrgTE2ya
0r3zDXS5ZMqwf8hNSIPtgogdXisFXfPgX3UfCgUcOqBlD1THVBafTiA3DG1pllq6Td1rq9zIO6Gx
jS2pTEj9Df8k3jfW+vuYtVRsd0ano5g5KuWHjUElbMWqm3lVcgxJKon8LcNdq6f3veCWFslHRFDV
P52bcRNqX/iUbFl+B7HpA/ybfaGZU/QE08Xz6NDI7Lb/PO+6vN/N2L5kRUYkRl2wyKHt7WLvcVWs
qkndLbXRckUZNaBzQ+KOzio3Hezvd8KvMZLEHd1WZ0n55zohSEJgkIOaVyu6I5/NFiDaelIZi8Jv
mpqDLd5brJHQyD3x/MMrOEBJ9FUTrI0mL+iv5FtVHngdcHsCCnntSbV2naDGzIu5b+JI0bC2EKaW
5OzxMTZVaojJTmOwAgA7z7QvJjbbKlB6PkZsD0SsfzuxhM7Lg5zaoF7iHVMHutphTSwyjFhQUib4
NynjEgS0B7/2hSyc+WGLVVts9f2icIZpN+iWZd+pjnOvHJhipmoK0kmiEibQ02BEZqUwAq9vLEWt
xW9MNvG1Da/r2hYpLPcC19jawdls789PGQPQ/y2sWETcqSrDdOIEGVWCrlYcWie964Wn7yBwu0eK
gRNaUUj0R3Id82LLJAcwXYJvOBEtJy/Cy/eqkqEwyACARtjefMe8IVCQmxcpWvzk/vnfDMdQRkeE
whtaxurlQdIHWh9XCc1VAXmdUeEKLIyQVGr65pSwDSAIdeOflzPz0rckloY35LbBfTryLFR4tPYk
DuN9+o3jOWh76e41KzC3m3sPTvNDRyUEG4gPlDB8LVBB0LZLB4ndkA6hvmkdZ/KFY2UfybnH0c2S
IKDbeEKbnBXJ0Faz4R2Urv4NW+FC4j0NWlgCx2hGCxxo23hwoyF3dSegntzxLB7sNTAIHTxkcuLQ
67FnvIKKQfpLIakd+UjdN4LZVqUd4uyQ8EylXqnBnlVub6sxxIddbA9tYeqm3zpeQwnsfC6naBus
mWCD3FMkM/NpIbgLCYNfvt2JBn2Ih8eXysm7+xbdg1ZM8NuP+ISVOQ+FhRjBj6jWGVcfaoY5YYhX
XpakI9s8uTUOB5FYFeA4XGLmYPxhZhv4jyBTL+z+NPbJRYAc3xcl3gyPFlzuztwQctC+UvC0QOj3
UjfMMxXDa8hFhVtC7Y4hAiFBir/BX4CNK1POynj1kViHkzKpU4c1xI9iOWh+GzgoUk7YU+kpGVM4
MgWIW5pEUSDuKKJH8wCUGHQK79PPE4cyTsJZWf/xcmbu0dL5eDMcjqFBz+MOncJloo4gJxm6Q8Ci
1VJw7YkcL9PvTA/PJIoO/U0qEPFi1igX3MroCEFnOzlaATRcLeLcynpKh+Usfpw1Ynl0MVmHHMP2
H++sV2fI+IQMJp0RHFQHseN0/pUdZzH81xvxDgANz9sjVC2UZa+HqFjbLk+TTRjgLFiLuzB54qZ9
NmwDEimz5vHl4lX3l9cfRvst0QdS3xC8ud/+poVOT/emYOCt9cSA48/SEC0sX2UOWWhORxVFC5cq
igGI49HiBVkWNvu1nvezCXwi/jV/zm6qBv5LFeFmO7pQaaJFkC4pUOMAIiLXhrOOcAJPMTdK62C4
jVK6w0+4xXTKAGGsAyrvpNxuYqIuWq3g3WqERLPtTFKtwBtDBynSj48PlxbMC8C38OIB5xHT+MQi
S5rnSr1fFtGN9dPeR4unQBPr3M9RdSAhjiVahezkn79d0re5ei8ikwLYczwH/PIHvNZcyG8eMf+n
hrTNTLBBJUgTP5fN4jkNvg23OCkJY+GIuglob2SPJt65jPMc0PZHJtEZo3Qz4HNnasz3fMKOEt8d
pjG4rRd4W2Pjw4Jh7n+w7NZLL6quOMYWLXPhbjTe/ILlE2i9zawyqlevGJ1mQ6RtYV8FQ2cawGen
6WqSTQjjWG2cWl8RbJV32q6l3jHjTv5DAzLoDWwQkS9eW1OaWkcE/0qO+c33o52sJbiaTegdkyZv
1FbbT1JGeib5sl246wmLCeeVx+1cKM2J22r4+58L3Ehgo8yldccT9wdQq4BUJKVdSi+JrncYfhyw
S8CW7WBPWjfjuQS/5/lI9DK5Y5K3wx6kt7F285raxSbuM4Do+luhrpKkovB+uZgvFW8dOgqnPuKN
wy4+2ktE3uOTwOitdSrXyDCIgQnC1SuT/HrOqCUbuuxGV8Et0f+sIY/2xiTuQ8+mboAp1nQJfenU
2YfHGqmvYeIZcMMCBMyDNZxwEL9ixK+2MOqBV16m0x7034Zg3crXvlAoZ7Na7mi45i/efFZ/KbU4
yZdC/athcI8/YdXQNM+kGIfoCy9qhV1zvrt/HiktE0wtZC4ycGoXtOwDzgG69zVsXOItYdEpPmB9
9V1Izv8W95QmlO/htEXRGOz9jiO/TjiLbLXabHFeVNX6qPOPm1fXuOELd/B5UrAWqD4tOsyxz5hP
6m07eehs8OWgXp9xjulW1+FzkqAZQmx532/jQgn9E8X5ZBNDTaM28QrGDN4Gne9NTtUcGiXzwFNQ
B3mJks9F3S6YZka6eBnE5XsiQuEt6D13M84Vl18Oc8SBjMlMp9MkJlWQUNiOcb9wqNCRYjrp7Isq
4JziQlp6yp5OnvP07aX04Q8qO40kWHVmVlB0Xkx38BzA0BgvoF+mGaqvS6P6LUphH/hXb6oDzaIa
TzD9LxziorUCgoBi/jfaX7geyGRHzgV6d6RDDZ1s/CpnLtGFg/uJKJQ264/PXu1CQVOrVHgnroal
m+BBmPQFzj7U/JWMUF8bnA8rA2s3GOzT09w/Jdv99P3d8P9siapsB2GMUrRQFgcu8w/giQig+kMe
QUnczK4PejTRbQHfJeYtd1O7JG4CRf5NfFKRHwpOdkTuvTK6JIjQ/cA7kSSbcKP4lEa59ANq5QSl
vtebjRiCGLxL66bCmtRvOwJCXIt+XCqcYyy3f9jASYp6tV49D6qV28lB5iS1FbRZw2HrTryjbiDs
yX7HTIhopVbZjePRtqjSOAXCbhqADUJ+Jzarpx2y2UUiAEBKmrPANYkAP7Rh780EuummfYqDtWnC
Iu4f0+F8+ubUagrzmm78FP2R5qB8mCo65wPSuvGfH6YIuz0IWqM6OjI/F/ZrKzi5dNzHrC3BqurW
PB5w9Gq8yEEdGrd7uArUNR7K3WlDw50fiJVrCgZ4lMkQB+03E6CbuScziRAgR+JgbUSmDvMbE3Ky
NY2UBX7xRKNMYJUPDtZ7UAbBUydYGkMR2BdfLrFHqUPfwDkuzMnZUzHfoMkUBfiSPP7lWb4T6I1V
Ugu0XBioNQtQk/8hjbNxAxGFeseNOSW+cabk30oXoemXldrf2A3JgOHZ2TjgN+TqFnYWC4FG25eu
u8WYUDfmhzZlimTipN29hU92GBl16g+FE63T4AFLYXIeFdZLsb9I0Uk18v/SoOUrt3Zfsex7Vhrz
vwoQgJ4A8/ktbg8FXmJ4++QFwB4RxPUj2Mx2C2AWGHdKu6hunE0LoN9ymOrkAmfUg1VtmAtbg2AR
Y3BttvhuxWHk82k4Icx6QUJ6gGdgYbyhRGte+JRtFYz2dasjmkFu8Wh5VWCLI8gT7yHfVCYEQc9O
Kp1xDCYe1uuuY2EIgqicZUdfnehoqwh7bQNnTXLFN3KVgs9ej1WeTeMudQKM9vOtIjjOGIToJ02V
fg4GT7CpW/aeOvq1TfmhZNPP8yvAO2uJ+j9t57CUI/h9T3FALgtdswrP7s+fsoR4BmJMv7Okk4++
qJKV8Umzoxxf6pmb8BiKjgZiEsMmRCLwMHcuCBbvFNBJEjnjdYzvYAs1qMKCdk8be0jhY6qVdjIi
F/4HPraqKBqd+DL0Tyz5ZZLjY2WR1NFT8WxDPKyRKaV4yM0qchvomOZHSxxJ/GTikvlCBv+wMSYk
4uMoanDfo2Qt0lnrMcV+AQOMo5e+0XCkrJXkoB2KnI9+e+uhj4bIG1aUirCQz/Q/8+KASXZWwHtp
SzIMASUhNK5GhnwMSvHF5fQZEQKGYybdlQ236ZyX6YPkLhDZMSOzbnwGxKBnB0ay4yBdygjNvraZ
yRHhlBcAyrT5l/0pi688+ODCrKjYr56+bPIqG7TJNBd9JW1vbk0LkOvMOQSmEAWy0RLvXPpG9LGz
0E3M7WWVWMm/vlAQ8bWq4WSOawamrhfc4mmhlMw48z3OE00PGMAvEFEYmwA9r7EGt3BrQSnApR+z
2hzWw4nT8FGM6tIEu/SCUIKbOl0/4wpdVncQ+dix6KRTn5G6byJaIk2o3+9EYru4cwNuPHoFbidD
3LHOl5C6f4Odg12UedC0jo0Othieq5DIMW2Fmu6Kg2lwzEJRRib8Ufaj5IMABEqDsE7M6E7HYxYH
YHsHB90TcTnsd7MQCCF3g0vqbkTazaDqxSvXMgjnW/qSNMtwqWCzsWUX8z0gTiJVUxMkb46iElbZ
o30TX31glDLGAIr7DLBCD1EGXz0p2fCHbrTdA7ZN4P0YRl68Ai8cdLUAAF7sjBn56bmhTGb18iFv
YLtIs2sOicIGMhmkcLREn81XQ9Hta5Dd1IrHUPirdK4Rj7irsXci4k9gknOA6NGoIzcLfbcAXPj5
ElcrCI7h+8H+0iN6GV1VWJBPBV/BfdoixC4Uarc5do/CY7+Qt6/Xo8tg7J2bbtY9B5YvRkKAS7p1
IjqUQiBkac7TVfLfNV5uM9X7ppFwu2BlF1Vq0voFtlef4WdJTP3+MZMRoutgqLlIrIZRfslU0/y+
OJq3YfxfIIYHW8LFN254MyPjr/fhqMAozQSDYOFmamR743IWE2ohkEvgc2XS/HSG3qN70QoUVbB6
qYE40xOY8jFtFqt5xzHJNr4aWzYUNBXkAsUcbOXNzlslXqQODj9fOJ2u5xACL3AVRVpLJxm83e0W
LQXMqDzwMvrgPQJBNNsyM1FiJ1PTEYFCYtdD1JjEUJVx5vElcqkmk30L8Sk9UdS2CoUgoRDTdK98
lFPCFPd5Wn8nsm+1f6pPGDt4c8boxOl+NMa8tzBDOTogZKWCAdfaf5sE16r0m3A6Lgn6IBOQpGlM
pzNVuIcoCVMhZiM7hjECsw2xBtJCW4d4EIV9hnB+jH8F49XiIuRjcC96NSFUBBVtLa61vA4m0rKs
B3c+jLU+XtL66VnFUJrp+GOrsd6JpDpu1iC4a4kpIBJZDEhwYiYa3Y071tLIZx5NdV0Zhb4wWG+5
Y4lGjyYYkGFoM5EW9x6hbEz4mtf4b108grswua/ZDKdRFkJ7K59i5qNiUjJ5/8l9NOytIUrpXrOM
T8LxwyjtRZIHtMeDxaJp5LezfmgdtX9zJ3S0sSP1TFPMcaqlmSpgrLeokT5Np4YERJPF6E/ufk18
J82Px5QiuX2u7VfXCmkREAkiMF0mBjCMfgChBeAGqAUHJcXNF4KoMhHxzhraHWkI/55CwMBCyC5F
tn7chUb1OgKP0SuPi+d+zUeIMPCIQ66psdUWk5tbs8Zlp2b+gduku+eDavMJI2gpRKHFnQmnhbPx
S50X+7K3d7NWYEClxI6FH4wU1w6gfxVTQEnD0/jndi2nJeDFdUBb0UJOe9iPS1Qhdw3o6VnliwUN
Umn0zIswwamT9jwQreO89/8f8b0Tn7Y3U6NyiMNLtP8khqIRx2j88TpEN28R8qKEY6ucyTZHGJrg
TXBJOfUO0SPzt9Bz0h2YWbCixDBlxLJaWmuyi6LD5UzS5j4gfBykUdnEqnIk5GDBlNCBcy/bbczw
au0s+1vY2zJyOnzutsMschhduIUzrAB21YjPcaPDtRpXLHULA09NMEClMMN10DbJkmIozdnPQ1XY
8T1BzYAmqpLQMpmOQkNPTRPUs/fUb1Y7XMYXk8+FwoEtl806qlYEEZiA3UfWsbHJvJvJ8WeE6DPs
fM6wdkQBuq5ihIPuvh24cftpoaBDPSWIyick++Wb16S8H2/IAqfeu0mhi7/HEOa972c1kT678mH7
jvkkARDlGmUBj9oRAZdWBO+yjt2XDKTTXwCKfYTxN9Ei74Ii3/KJBxJYFAPSKDxPbEdDnkLmBA8V
kGjT4Bu079+embTXvQe9TETDN3MyKUVLEQZU9Tl+Sj5rhcHKvLKltUxDtSqbzeeYHaN4pjKHIpNJ
QkpmfQMTAKoQa4QQzoTcuXSzs0mMU9acSiZfX4/kLIUYQtU5R1EWJUtvoHorsXvkS3o4iHZrUZlO
8LczWLH967Cs4MyXGWYcZRfe+h2hsC/u+aEBkpwU2sM6f3sCiaN7VO7iCXNNgdEdyjCRLVbWZ0WS
DLQ3p19dASbqPpR/dUQwHdWtVurIoqEhJfNhIol+zZo2VykAl2S34bp8G/vVSnzu5yCxN/RsMaY5
hO56cFS/VcN8XfVNSaE56TgPfal28W3hgJNDMvITEK/habd83Y4g17lK0wvvu7mdp9+NSdN6be10
0I2WxrYIND0ctNTLXxyinKIyIARQhbC0GOMRUtzsBPqcEyVzdIRLWRHO8E8Mj5BzmgmSpAa/Q7nP
WnLBF7WSg4FUdZdGLZ3xqFZARjLS2rG/K1TLqR1/fegZDkuJmssVhiAcdZHJkLu8hy/Il5v2F+XR
FKj0NxNpjf/rUtmydf2XcW9ogtz2Mdq3oZ2t9WX5K6Ab4gn0MBYc6yqX3vBh6VkUt/WszyI0rUiQ
cIqzLO6XMRHPzRGwhGfo/yVmJxYjeZ2WkWVKIFWZlTN7aCMjg0DgUaVw3uTPdGLbNbt1YExYyDNV
DWnEuhgzmvpDQJte3QCsKd5gPPs0/dX50+TqOSaJje/uEpqzCneagcTjUO7kHjWkMskN6TtcBDT7
UGhoRpq8WR9fekA+CoFzIYIDKTi6d+OvcYwk6dnVDXjt8X310JO2y7AQ9uA5qFAJThSDWsHIgk0Q
ApzImHYQFdwjsqfHSmMfYkjBMpbe9imsNz7UjAYztN03HaYPp88v98sRTpiHEGipZHIwkc2NC3dr
7tOJHJb85C7f1EvOxcUGbKoYH0k5S+pWBpdR8sgUFdjoovJvb3r0ZWBA9rQaSe0NLWL7sRLCJRM0
w/2PhXq/ZN21A6Bl7G9YG1KS1DLj78/ZtdS289c8wkZpO/2KG7A1+czQUUYLvUNY5zKsseyEcuEh
IWZzvSKPkkXzabs4M2K3epiPI512LFIWJrIEjE8OLGU2gDgowK+XjTFEs6i2g1cSxEOUkO666WsZ
xMT8PiuiRUZuDKiYSRY7lW+s7bMUIen9kHSkBRmYDss6kW/IyuTGKSC/dh4yYadMXBW805GwJoeN
MyyG71j2mgUuuVTISD7y4HeNpyRAp7id5zQRUKzX+M0TGA2tFWZzEJcMhBTkK5w5vq56DhXd4u7g
qwXCVZd6MH+2ykaHeV8nT6kyZj70V0AVMunKw6fZ9B2N0+XXcI9xK1sXFf9DBkKnkz+HZhKwb/fP
pSjE8Uczltdyy+gzEpa0eIJ3sTulCD5um3BOUADehck7cN8kbBIQQ7Hqt9Vflg+CvlxFADw8lip4
ESWymBod7QjqNRgFBtc+l+ppqdUwJ+Shr1rwOVgpMrom+oJEY8Y4B7WrD2rz4CQ2b8qYQaRiEIlV
ynY1ODpZ9ff4auDp7mSyt16w5XOxzPoV9gZcbzb89Vp+em+DpEEOtGSsGlY4qcamyK3BSlb9Gtjr
/iudghrDOH8EIyPs8KqEPN1E+L4BWt1BVf1fUkSEiAtPNE3StWXsYZZNwPp4NpURs3m3Lizdcu1P
RUpHZ6vbLaNPQs8U9K5OV7SGsumn3XM/GPo6Fr0VUeu+LFNlhFG8n+qKOI8BgSf9ZdK2ozDTN1nY
WKG3MuhoAT0lrkqjA2lrNLRXTXINCCMKL0bUjpRxhzs1J24Y3vy06KTDCWwxJjfg7X25zcSenh6f
rNrzXtE3yvbxLZQEUoyWYTgQP54x3hhGIsZALap3yQMM6jHdQWl2lxg3GI69atYUJ6c2h1YBSprY
rTILSjCpFgRz8rGWu5zIEJAwHBtT1a43m4zxr/zkmrRLwKALeaRqwcbJdg+3OvDKPY7W+rBMnMBT
XC5YOQOFPjIWMJw/n5rT8wdcYm2+r9PtWfiWSxQ/uVasJqoCK85bkDeFUs2hNfk70wYsy4ecIJ0l
2rhKSJf3mBHOKHtC27Q1GxLNZ00+Lia3FWJWEfJCmLtIlt3X0Sr0G9gRkF+NLOL25YyEYgi8Zy4x
ezyZ9UjjOpTB9ge39IHB5ojXy8mf60ljnH0wyn5C/vGDuv9UAh2s+pDQwpWlQgac62MA/dJtZonA
LwZ07brYatIhuiHz5HcZu4xu9kz1XMnUiBgzhzFRsCK/Asmr5X7+vV+q5v3gJClw4/n350atbNvH
c5sL6cmrRNSociwhy0jvNBNxS/9+eu29FsmqwLMPvgD7YgGnDFNjw9cXPVqhvyT49WSRl+kerjt3
vbbn2MjeZOUNhqQNSTWL1YaheKZQgDw/mGoeioJemHvpyVbZkRDyF3TLlJa0BBIPfy5JwK5Rws5X
jQJRmDcqlI++5WST9sRrx+dsf8Wfy/iykDrPJbP0EGHJoPLrHlDPOzc2+9hVbBixnf/kQji99T1R
UEiEaWzDFrnB67vVvykHKnABKlc2Efx62znaAeI4BmLQ7CwnQX1MTHY5qUKoUvmfPtsVR4oFY0XE
cYjiA+L79tq5gLxlN4p48bKUdqyyjSi/mb5mbgWrT+LGd8JCEvJj3EXXjO9bCrZBtMUvcWusVCke
SdBL8iPCaX06OMz9kakKTnlS5WbHI8/5Rk4bBZVi+CLL8SrRGGznSkh7Jbu9U0zG+ogcdnxf+bon
uzyNl9QO1ASELOgrE+y/IKBj+040Eic20LjATJQ+0Y2AtEagBqfzqXmXLr+Ij48+ibTB7EqxIbAm
RZ7dKJp1MsIuQek4tkUSuHTrD4UUDlXF8RCwxUJt3jxGbn/OMIHltBkY2qVDLnt7BNjc47lf8p9M
+q5Oi4Tu9mgI29SouHlhry5K5ucY2xrM3nEDZNzsq8e3rO4YkDFesJQUrFxGa8dtKGqeZXtS2cI6
X4nqj+FZwI1XW97pi++qE6p11rNJhLeV5DYD9m0o3+nWCaZadyCcVVKrxOxSEaJl6lagTDzog3c3
krGnUMOA3dqVepMHQIXoCN1oUqlIfKUXwnqXXyPdq/QiMovrRmY6lTe/GhlbEagMsgxUcjRyeodf
bSlaudPYIXZ2av/SA9O3v1LgkpSOyJCPYCNJWLltnRMu1/o0kV5QVHDL5s9XTdA0PtUJX6lvX3Zr
W0sTK6PaD3+6s30vnFuRngFTc6UQvcGQiB94P27aDxRaxO1U2bG5sBUoZFpxtQ8s0GAfLVK8H4kp
+8Cq2vYrtIhztJUvu2zCkXqWh339ZiXqJVmXT1dxOPbBkJ2Zj3up12ieY8MlKD1gTXdD33zANs5H
mwUwoKgqwcvZSqtw4Dek1K4JYmMkTS1sK3Jft/n8gUV1EYL7XNLzGnAic5cZtPWNpxY8QfF6r9SV
+hxv7M4GKN1yZL+NxW8SGam5co1ini9EBKX3QcbsIZwUhnwSVlinJIzpWyv+jTbyDhlosKb9hspY
qWEQSelFT9Mlnu/uAYJxEWvgVFQGjH7iLo3SZeETQZc+2T1Ki/v+NOZ+vvGFe2r2W6VnoI1bt+P4
PrGa8NZJV+TXEPs2j0V9HPDLLPAAV3h5nABkjhvUMXmBncOliXSSbBh99KQWc8pyxmDZ0p2eMPAY
5IjmrB0PULXry10q2iBiMKUmaKMYlQd7+KwGNHZ+b8su/ttP1BRujefvZYRn9oo2HtEaSqBvVtvP
fesoztmONKkmm5slZfhBR9jAGCfEn0c/ALBHRnm7WuCNGEIpCCK6O0JCXY1CLl5RnNZ99uheCHMf
vWDjVCX9o+YgGUoodVdZwt6JnHbe9nEripAf66bsxNoOIznnrDIZlGwRof4ObXhzDdX/2ieCN7GK
827BxfLlffAvy6fEaNcoHdiGNwg/U9e2HL5OKGr7E5i3R6rI8+NllEGaAnWqeFK52Qr/Ghxlw/qn
Z9e/4Qzvx4KLFkHTyBlXRQMGYvSuCUFavdj8s4m8r9sz7NseWFKFx+Dc98GjjksmHfG+2FSYLQtx
Hkv/kMzMd+6AiH+N2WctThyr81EmUypm5+Fyk6t1spGw/3ALVoGYqp8F1DNpnSIT53tKx4ZRJ8mC
nfyowL5+5X3t1efujwB7tDqT++Z2K44O10vL4rBKvPbGG1GGn+pxk54F3vj2XEUDKWdG2jKqJNtT
2YnbL7jbBGP+h5/WTxO80eiwlzYGxS8iOzQU/F8bkiPjV5E8S/cqPB5DGOJdbEZ1BvCgz/LK4ab4
yCBCtYDz5893Geu3vImeT3ulNZXJENU/kVx7sJVWA/zf9BjyU4fO8+jhsf6lLIqi7Y9fD1f7dZdj
YsV80JyqVwYYBtjZy9vxosiZhYaZHl4CcZWG8RmNWAAN7joAfkWg+Z584/YBPRDwxER4BYCBTWbW
oi0IrcRj542GXf5+c2No2Up42YGf7LCH1wExXfm7YuX+2EeDa+14j6+YLDxvYv2RPObW7/wbIQIH
McTQrqJJZV3j6w2eFUcPs+tb3625B5Stabnmp1hZw+nb3qbzuY/6QPsiUXWjbgagNpQZJeWr6LGB
HQA+TR9bh1D9TG9E9HbmyLaXZm7MfwXZgxu+fEyKCwsBJ7jnnNz+Xo2EMyU8/bRSOOOGX+0vvhKu
Tk1J7QdzFRq+qEK6SCLSvbi8BzdDK9YBeNQ4+XtP4SZzjLIAtolthWf/RHjj+20GEwKI0swQ8hu2
Rpnjax+V/fkS6dwgRRwsyaJycfQKYlyYXYRvgmTWGlwM6dUCEiuDuRi36BsN1JuOfBwuaNWNqNWH
R0RJS8AvPxqkbBuHX9azLOhnM7MYDQUC6z1UrdeYSfGXLRIyrA27q7dRaZbcKUfl12IQ2UuAyo74
tyTJehaalx/X92EH+X2AjtIElacAw2h8uB3omI3STnpOCDJkF7iiZ0KOIVQg8JWedxLQqrkvpazN
i9byIpS800BJCyHu1EEZ2KRzEgQ6pylzbxT5vTe15POzk8UpH148EOLuHkFAMC1HtIvKqLNT1ty4
MDkqhB2DGKdA4bRqSzqQa2M5iKt3PkEsaGqriXcBMHHkhEjdZFwfU0g5Jl5eXGJvxiL2zuPq37D4
bLWfGy40yKO1TGxdYo/QNEfwQSEdX4qx6BcyLGZDAK0VKbU2jI00MBCWjz1hlne2nSPSRbeBtKQG
OQ7/mnHDLIPv+ks+u+dpzpO3ezYyKgeAMB3RNJBsxYjqyuv3drbYJMEXyjwdFBwNPsmVbmd2kSHO
c56+tWiMDK5zIbil7v2uBZQTKkwaXQl15Rl54gDWrrmVTPpm6Dino26ekEqthUVqDzHWG9G/zTXw
X9SXSZ3n0RvMfk9WlOmNd1JzYvGUtfZWLcZdGAxFSDkmAdHZcwf2po4LQRP3T/dQr+Nv0QvIIVvc
li2yTdTogJnBihPhQ6/GWZfNJ805qVHzmBTA3IiCpN+uOIwirjHVZRnQNAk14PSlwqQu7EAbl1w7
FCqUGy771bp0fgrmEMAWUBc5knokaDhBHqHkJuNL5Ahi8V14KcFPYMDpg6jnpHHBMroZLjick6fI
tDNMyU/aBDr/JNtHTpHNym+6GAf4mRSY0fX4jnvLmugKPRJpoKvh0ZjdwDk5gsu/ZpA6Yz/JFS9h
2M8KiYSUDUjCVW3fiuqo+79xdLJSh6g/QWFmGs1J2wQiYnIWqIyd5Gjf3q9dWkSpech2O6KST4BR
OilXfQmVa7mD70JJ+JUfsAnnD+Zd70z8dxprxYdOQuWOmbYWRrB7po8BOzGyzmBR85FRiyU1sE2X
xdgl4GbNnUTcm/8aqhDB4JwAkn5/YkpVF3Ieq8noQ35RUKglqzdm0SAzrAz+YwBRaMOTtWvbj/h3
1JVRtJ+iA72sFt4WSBrY96Kk+qU3X7/MkB95JM81hCvIMhQxJPhl9NdqnETEZsbiTDweCTXIvNK+
6xkXqKZMSCMEwP6e10MaieGRVMyjH3RBFtZ9cJVL0bc+3F9EHInyy1TfbYN74M+VyWU88675l4tt
fgK1nT/dgS+l++qyongiTcyAkixYEyGh3q5nJGGZgQXx/wsYMBEZ2aQ4TpaZr0YW9kdNpjDs9hpX
JYM+fQIMwuYYLeb46Xk8zeGl1TtAgcQLIVIduBwmTfV68cTFh8f/o9lkQD7zXV0M/yZMCrcpHAtG
GShIIm47/5xxAeNqMa28xwPekHWccxwT7aLQImHYxf6BdleBK7ENgxA8YFMZv7Md+FMXnhj0wN4/
U9047vDgbrNg7HDLFgDb6CnjoAqRUVVvYqsIWRWGbLMey2ri6TGGCSoX99g5TgjbR+CiSdD8Fqje
S2VNoOoLOkqfkFbDv7qkHPWM4wxnU8rd17pWnlvaGLYNsQYy2QMesqkkKSufB4zhStwvB4TBCYm+
Cd8GmwIERAOH98YrJ6bulNaSIw4e51YYcjwDPToTK9JxAnvQyw+6IZ22bBvcW1Un4QXbrJ8wIIm2
nQy4dUywdxhYLc2VT46w0UjcluvwqNbx8AG2VL3oktO/I8mw2egV/dyc0aJLLgGLPSAEyss4n1tV
9qlEbxjP5xXcqJzc5ZJLvj5R2nWQq5kWl2t0TE4ZSy67PcrXHfHoq0dEpPKS6R374BT+m8RUfADi
Ko2rLD3eEmUbur28n+9g15NIxFsDD+m47hlFqSXbLY9RlQUujU8lHalSX+m4EwuTBbkL5eIX4/Do
hF/h4k6uZMEJsZpnCxQ1H12w8beMTDCEdkum44GdVFbHWbb3MV251JP19LqTMLeZ1EPqUMJSbV08
x6JQE7XNdpJ12axd6WqM+fWOzWxLNfAz1B/ww4rm3PKF/OGnnZ2K6Rtip8+jwSpHoxEevS+C4+la
vmlHIYfa5RT1ptcP+enEZWYsGFBT2VRysYOdLmiJem73Gez49pTqOsfiXvKf6tyYbqHCvuQ2wg/m
V3UugEzFd3XcUUdQdsC4nhtISNf0ZdPotLL7pvH318D0GUhqXDSNv+UxobL1/623Ldn7bC+uWJoH
NWcqZURv2v8ORE6Oa0wZSiW0H/NKlr4e2RtzC3u0V/4HYMXhtg7bKd9hA7AnaqDEMBryT4criOmx
4SWJLq6U+0SfqvWy6+MmVWN4TIyM7eL586mOJAyz+6uCpNrYasXppj/8UWfow8LDwkolPrDgy7Fw
fzs8cOt8F928OJJgqKm1RDIh3hP/iEajr9u6Fw7jeb0xJ45E+IbmOzUm8hw0Gvan7YTDXtX2dPOm
0zWE3GFoY6Kr3QFGvyJ04Tcrtd+mZlPPZPpVCy+DoA0YbbjasIpV5N1cD4qbbl9AkhvPFHQ9e1v6
E8rZRqkaRsFVx6YmJKLBY3+NR94qAg51sRTncgDDYxvR952N544cAe5hmB6WoaJ6xzSo6WnvaA3S
A6hlict/Eh8REKrAoqdBXEFnNydsaKCaasqxbaldTXTwXJ2nh1ChPEbxP9HRXrMTpNTdam5td/F8
KHi2V1r+RsbMbnOam6daAhLM+I5zZgQ+9XvbxDzq0uLtwQNM9QNn42xqaq0zC08CT42YlhHms1jO
jp6M5DwMdabjyddfq9Hy+hLEEzzxXgcKeOrJiSuKR6+RbpQ55WuyyLBiVKt+YH50G1bSWKV8Oke5
2WtRpuUoPDpmy01+AxfPN+x5cjbIeDt7283VUmfA/leK0QYX3/CZk23fTX15Nv4fxekUatwSTztr
U7aiEi0SKoQu8pQB0/6OXMnC5FlR2yuWHLbBWjFUDL9lugla2XbIdRdX/UBHsQ5uyV3YaN7AF0Dt
5m68sZsfvhg+3xujwALK+YqRK2qqYl/GIp805tvL8T0+ElvxDqzw3j+5U2rqqjppbBcJJt9tRvRD
36UNRShJ/ykvHH8eQz7BGG6ORNDYxLM8v+A/kKmF6QSkvy+5Nk0580sNkLwi5/iMPQuL3pc7ND6/
P53ZKga93BofUL5G7wCMJb5M/mNnJOIMP8utuuXDtEK7DfAuwK02o7nmz/e8jfvZ3rYRGGvdMNkP
8l1ldc4fKhOCu/N8tysyqBISpdbaQyzEF35TJsvil7xiAvNzixoS/Zljn75B3DgUvUvDJvyQBoRJ
VMqAMSHYW1/51D5baBSvtsT1spu3MK3HvT2jbf5dyHvnpTkAq5alj3jZiBLnBwQzeuahPQ3LqUBJ
TULO3FYa+u6gIwhR6bANU8DLvRBlqvyHG6pHS4bg2cUxwMCUww2xJ/eCb9kYHXXRibhxY104zTfl
rsLA5m/8RBWl0WjnmTORur6IeG47oTB95/GDA1nZ7FWKTvAbbLS4R1L19dvpI6E95GqBXBorFFB8
gIU2yCbxaXBMjcoSjNLbelEB36BBzgTqHldIwd5lS+lFPEJ7rUwkFCJQRrIFS5dBzUYlp1ts16xp
Mgb2ZOvXMDsfqG7ZWx90UIELEh+qmDliOuYwvNq8jcBdQQ2wHQF1raISuwC4q0EJkSm5LMa98otl
xWvRg5xKE9xlKEXWMiGPp6AyBb8h9rZlW0QL78na3chff+5tj4ou7cZg5P/yLflCUFRDptGXrkes
RyYD99Pv+QMLVsI3Ux/IbNtd4x2ng5pnfpRBowUnsmAMzRqyheLPxZoLNpKGH4vYwcL0C8aQaYHC
PG2ybgplj36ERLOCXiQewhRnyOpritpRUXMIVsaBZzWTXXsszFFVD23vwrnaXXd7tGsKUmBWE68o
u7oU+HVV7y0v1KOyftX0XIT2jrfAYOQgpuwenErqQ0AQ+L1pf6JkpguLvWBh6SVeRXXaw5Ltles5
1e6ea1Ac93ADvHIN7FQ+yxKS8d6hAH1uaOjhoiBHD2tlAe/+HYBSxNddhSbuHV8iAjremfOQXK1i
1RBvW3iqZtxZJLoSCfqqrm8G+8zrBcrTufUZ9AkrUoWUjuyj4VjuKNyrYsKeUm/XtXbP+qMLXA2d
uEixurKdDUe9Nm5oe0SZlrD1ynjWSjI6AhzTcay+ENqmf7EpY+pwmRBGA04c5CHH56jlqBTGwkE4
Zfwr8/6hTiSIwWwVUzPoOKc8VRA0alFeYQvHtBr/ZDH7BWXFfNL5q6ta2UgWIiK6Rfz7l5FjCeK3
41BjkZS8vZic/ik/HiKZJeXsnTmoUNovajZzwk4/JY/RcIFl1xAIjFxwTqGenrvcqyBpq0eSyrfL
oBymmnwxIz6Zt/v1LhH+jJmSGA9LhnT/Ld75wg5sH5afuIthwddb+72XE7sqAYGblYrYVLr2S48u
0ZJEBthLRP1x9MfOVeGRCMfysu2oW/l377bEvcII+zkBUAPSiuDZi7dHL+SW+pmsxYHyVT91a+Lj
HyszSFmuZ3fBcC2pH21wTuJjzT2TdKoQaSt8rNtu9ezryRI9+mKMyXvU6JHQuHTgS05FhTj7ULuf
/056ZQk0bhGwIG1j3EEwq2tfv8aH2C9QiNwpvERXkZn2ebl66wPpAIN0x7aUedLQy77x2inEaUXh
FL3PKJsXOeF3F1RTeV3OmpdlOdD4Ccrdfg+hfocJvf2TGiFEtJj/yWumDPuSvhXgEq9tLdPumBv2
5U+R+whjXTFmAOgOt8pJc3JXRNnTQWDW5w2d7dRzx728wLsLwb3wFdvzul4Od7B6Xvfxg8W6Q4ga
movfJv0//RUhkKvu+zoVEHU1YWzA2A37phVDJDLeajf5vWVTLCMsAeyEG+URzctJuUdZv3jhvEo9
4tm9AAz1M32CWzpFN6LqPYs/xhz5e8xYLp4zC88l+mhMn5sQ28Y7wa1twPYs4EvIcyEyP0B8yqhY
Idxc4AHse+MCf6TB/vIKIoH1IGf8ujh2rIcKTjBHFtD9BDUDmIE3Q147OtmiT5A8OgCiHrGW1qDG
ZKYwGCLxVJT9+UfnF8jgqDO+K2eXa1TRhUyv5xLnnG6NL174Am9t+hdkdHPc6rHqsxT38xVg5RyE
u3mmgv9Sqc2YhjC4zCKbHrubRzikEAn2YQGlTW9AIfOp1UWK4irn8FLEm68Lpn/xTraI0QKTHyV1
rsk/DnB2Qzk7YxJA/Fzd2JFn9pjaYOEh3Xaj25cBHWHXVUjFvvwD18xHOE1dH221DpFI3UH1efMO
XRqte77UCuH3i3qiBWQFsMPlGtNBnKI/kJH9Swk++yR10P2o1psJI3YGTXwuxV+csda41FSW1tSF
wlduNU5RJUCrWbNBkcgSPtv+rPiNy1i5Y10GLNx47t9PRO1/rP/0GFwkmgK3ycuk4OHT/4oxW/XV
8QuJ2TY42+Hhc4SyMVdWbxsp+pl0R1EweWiiekZ8CnJIs6REeVsOBrOFwBaegmircQMhJwLLjTgD
6b5B/OoXaQwT7wkD6BaOiM6yQ+jSTdd0JBk9i+JhIwVCjevkCv1iWn7W410pBvvqqi9b2eKuhmWf
AMTFpKQbFFIHEH9Sq5BoeK5YalbnWeqhp7Fysf2/vucy30WAY05+hA9g+LKpwQsg/V4v6HF7nzhE
yYCns8cOQ1RApOp/edQZXGqPM20BFPtCjAaebjrUxmrBpnZ7MPMDLjR+oyK3EYAMF0fK9pXoaEPP
pcAUwFBEprsBmurobbkucDF6pb5YPjoHKyX82ImO8+lyhEsef7NjkkYyxXOyQNY4zeyUJVQRBOYq
aDUhB6AVl0Cx0rpl0pDWJxhTcdX7Pemt8P3HpJOWnO6jO2Hwafu9HkrnxayA/ODXeTY2nSA87yM1
Nb3oYL7VNcAFqGqEedrtexv9HDG3Au8RLhUFiisfhV4f/7YnfQeq9jA9BZ5HWjuVG0MSx50U5ojG
yXyPC7hWiBmV7hy83hpidKYJ3iJ4yxXSz+qfQkLcZA9cO7yEh8e5V1VYlKOo3ETdgj8Yw9ic4+f0
kAcKr/EcQeO/9UHcso7WP0yTfKen7xn2fTx82UVvZayAJ9Sww3bqFsrnmlvwufL9M+yLyV296QAo
95P4kba83zsXqWauLXiJJx3sSHLSFh5T9I+li2tpLz0nk/AJZpiiOrSlZsDB0ikx4+qcp/4TaHzq
zp808BmZY3IndRuFLanAv427ijb+YwXm//xtEEaRqzPYJ4VFWsqLfr4VdEESPuEYud4zOraTCmWq
IUSA569bTR3AOX+rrjGKAH4mSjyIHaTbERCoBAWmd9eklpKKwy2QZvukaX2AxCAMTCmnKaWeD5lO
Qf0VJBFkOv+ZiOR42sj7t9qDSjCKVRW1dIwNFwhpyrZZIK+LbDicXU0WZHjfDiw5lTCqeiA1dQEC
TJ2Z93PxL0lhzyr0l1fBQBclMR5RHrLjGaPK5JpQDeOlBwkuGY770kicmcePV22JrypFh5YKUxjj
q65WNjMlX48RhdMj7dqf6M/+1Eft70E3icY8jI71DwQh6hOSIfmnZo54LbCJX/9DlkDZ6F7rFSO3
R3X3jsU+arHHQZb6P/6LghgtKnpoAVnY3NmkGofv8WHjXg0T1MU6NgGc/xDj5nAujQQpHJz2yoTx
ANkL1hzj+j4EDDw9b6icb0vu0kk7bESBypjXbyrTfSbE8ljVblcNowSojvuo75KOjOfL4bVxPro4
V/yFgQMRt6ainAKWmhPq1u4vXgtcSFGUtz8Tx/1Q14aTCAoL4f/j3OzzoLoyWcArSRmX1ZNvVWw7
2JJl7cj4KQFUfYIX8VtvQD7Pm/IYc0FGijsH+H5D1pHKkIfGS7gEbJ3HzDXIj2A+ZXQg3qvOk4C9
8gfBFE++3qravyG3ILnCc7mO2YktZMDxHk/dc22LkA1jc0NWfdlz8vTpJdGQjw2FPaF+7YsuIYk+
/spHF4Kobm7T+R+jUF1hUXm9SkmGNMaoELr5Het/z083zqdNE+7ILlwcCsky1VMdY/1+eLpM+QC5
DURaeLbhy+ieFP/Scls4WEAdLk+nZDBRMptE7OO4Bn4ANt5GFGKT7AAk0MR5xmhmg8sEFFgGNbel
tAx/H5QKBAG2e02HlAmyjigqGrplDrPzYZWDpinUNlCkluOE7AkVxpDXiglzvk0mu5KMxjEO+35r
KJW9/YCxeAszIAdiEbA25hZdVap+kohPEPGM9O1B6T+DDoU7XIQc6lkdnV1qpkKh104JnuJ6Cp+M
TpjOx/MCcD6JZ8TyToiFkCDnYxWVBEgtR5yTWuFw8C8Tg6pRDl3MK7gIBZ5WYm1se9niqHcs2GeE
Ho0u+uUs1OMOygdB4LO+StBWd8ppwZP8l2JGAbPuZlPNHYU9+EanJEm5xG3+qcodCisBX+CscS5z
olslu00aRYXH5vQ860V7h0cKV9BKfaGp6NJmtT8RakiKcEmUcP2UHInbOHAN2Ygqvo/tfGzFPeeM
sYFshra6rV32CBcr2XBTozQqqKUbP2QgmsCS+J4Q2VW7cvT3Kup0CkwEqrnDbvRAiX0NIPJs2DG4
w+Ba/VnCyCnAyxCaXRsBP8cRT/F2cGC7rwzOimWNZDVKNsuTMlhyFxq6K0XofDsbranQhm8jxAsf
bnfDYisXM4RwuBxGuIu4O5zjdnFJwT3HAu1a9BwjgecnVgi/GDl/pPDlqMJaBJiw171Mc0sYSvdU
aJiqsVLqFrwl9vYv50D51Ke0j11FusWzxRV3ewAKTMduW08pQTrfVm2wB2OvGv9CPlgeLBoVJy2e
Nb8lLZj7f2120/qbdo690nKo9fMCUdWbs8yQIfbbSuQdT/91U9qo/56VECWhpb+BzYIr2Rq4cv4i
Ho2CA8VVrVvzen/6tJHQy0JCNcdzZSc0+oMKgJsUDWRFLJY0hF9Nr/OQCYQzi1xKYKNM+RWPOcRc
GGxqs1NFc9KS6k5qej72FVq2mTA4KvJWteQXqRSOhAGvYrPNivvN3sbymfxuy8ODNYn3Py6Wb3YC
r7UDkLFRrmBs/6wQz+UMNOn4HtvN2m5OaHszfet9uiwFsw51BxbITOv3zxifeihRluHYeK40qblt
2mgYWJMoHShHjxr/1jpDAHpvAFcfnx55Q98/9rVxzWtqoktKyhd15pVRjDx82mEBh2Aqv2BoYV+D
lHQx+J17oCEDQTlans89bM/TDO+XSTadp/4dnrZMWYG7l/8fs9SiAxWOrVTqFiz8u29KYXwrTAIr
xtpwkACyWOSgOgy5vBrBEtl/iuAQcbtDm9EduTJrAzb1B+oYTlVk++ETXI/xgRZldCWrCo3meWZo
2qSmoowEmkbTwcS93G2DCRxjXA0rq0qzgV8arFvG3GB86hSjBCk9sAgwYVgiE2nMqroNYKn+Ehk9
t1lPLh8FbGx2A3HZeb1TJHTd0gmhNBwTGKHtAmM0ywQTDOai4YYC9SfpGB7xs5PbPcybgnz8Njit
g3XHHipUibyldq3prr6d62v6IG4SNnQh35tkW8sD5r9PxdZvFxzywNdcEGE2jFWDIlk75j/DacKU
pBNz3S8cfXeRFfXvNIExhzJT6ZCQ5SaDpxC+yo7nfENYHWOzvPtW4jCso9w8nTSGYBwcVgtA10Ya
gJEX55lNdV0jBGAVkZtz6u6A3wLZ0M24gfcgCFAiqZZRiUZQ9qeJRglUhVrj045Csa+NpvP3fCe9
iUHvuPXZq7ob5D+hSJ+tImLzFlMQaxlncf2HYQrUmxLeTO9vJwr0xJ182gQdPsNqSOkb5qScPreq
Yfq9FOPd9UnmloRSU7LNwJAB6aHLUhuVNyJko8GZZ80/pnVG0RsabXlLE/cRpQ3lP3iv2BoFsOEw
VUelHjeri9SWnW9QJZDTNzQXHGtN2/xHL5EFzMOPXjX0jGsNGnvNg1M8TH8O76NAJZc311dJr6gx
/0p+S1V+QldZew0eb1SpBhCPWQo7lHfn7DpjriOT4gKpAeB3JNacIBbGHgBcFSWK4AhaM+htDn9i
AaXlkQCD+AUzuBRg4Z2X1iIa0uWghfT838ntwWRDtPqLMqhViXn8OhLsIBPFSXSjbt/7Jj9nW4Pe
z6BAiEex+YsY4vEBFzm3N0JZVqSZAfCPeIsVdEJpgPQJ0cZQqrydoaTT6w3P1f/bXnTgIXxxQf0A
7jZpbpVpX9MeOTIHFA4EwvJY5JZXOZtl+FYB//UmBcZZiYBkLVziKxRjiVXl+CxTxkSUiiJQNciK
U4+4YUUC7yM4yC+Z8kmWErt/KcgFEXz+4ANCkTyoeEN+jf1iAyPE8V7t8j6GaE25WCAMcW48I4KI
5VyDeFDNiOiX28wNXMmpbmyZ4W4/7PnN5tWekiwt5bIpbZoJnGmOVJYBmGw2eJN9//xFEBQTJSn+
vyVw2dOtMTDUxPv3hWWhMtUP7Z0AofcQWHOhH/rg55YohOaqQ66BkppudxjIUAlKu8BapiLpsQtm
52oHNIKvkVT6zxlTUsqenfli++6JlNmC18iHTj+3o9kwwTNKmhLJYOS+GSn8Gf9fviDKGZiSK/4l
zzAX/D0VSlpdrk3ax6WXh50F0t0NvSLUE0qXfQzHbbEHLRXIx7esUEImp+ridh9zcI0Kg7BQe9ZC
9aZtRTxFNTkiFF88GuS29bzQutuGfROFi3xwe5Llmx76amaAbifC45cDvARJawxm+SVSNPQPiXio
qaqb+OsezTahT3DMrng2BzWwPvb5wv9i4fj8e5Lu6NspnRkLTwixoI1RX9cqj7E59j0cHXW3u9Cf
XDery1CEk0jDGPrKQiRuFSjPGHUIJUwy+gEUxJ47+uTYYlwcBM5Vk0HrwyaUPu9hukW5FW28Pt5Q
COuA/lcX2YFGZ6dqzBNqCpcwxN5YVbvyHQkyCaPMZsMyMsqizgV17TW9H7Q3Wcnf1uWkHwmiq8Xy
q+EihfRgQVgPk/belOXrqgyfIgTQQpH9bISzFizNqw49Y8fFBHYO/wCEffjHwxmqmTfuNw1XgWf8
3KmDtLArMpJFtCLfG/Hd68eSvckkuqwA81xWHRJYbnEnc3VT627clHOI5Wy5kDUsTNOHag1/07lQ
Ssv5d02Cd7KD9dCDwk2ktfwPss9mKo/eP0aobjOQOE1rgDxgwweDrpuMEQAZpeAne5rklPy5eSKX
wmY7eqnDcj4ZM6LWL3uAG+o4g1ghFh3t74fYAym+7+34d0wuqg+9AXOWrnDVjvjfVXKl+TUmM45j
7G+sY36UxqXE8utYdE6ofuuAjI12GMXpi+lwyPEeGSyEVerOYWZuoiSGb2pQk3NbIuNOUOpze2xo
jGthZiDDUpauLE+FvsArnJQ8n5yDhqnbBpLSdceYPH4ZIOYcekP9jHugLN7oCXWtouirx6AyecUr
u87o0ihnKkP64IZVnKf0JmPHylhOlbrFg5UR1JmzdeiVRn8ePQ5P/rZVtMqHS0OZok/NtWxi3Yia
BRwyQN3XuxHXaEkbo0v3XCIL1eYCR+Z5gnGVg3uEWXF9+gChq4LPwX5DRR52erNW9w3i0jV76wDi
UHkSGdtpTdCBu245t4stHGFnnq16TxZWHpA8Cp7JWKd3Z8Hz+rofqkevkNVY973UgfhkcK/v9PA+
QX7jh2y6eaD47G1uUAx3e+wWKZYuwS1ehUPxtSmKdsoJfAGQKmTfr7CjUlmby/p67urByHnxIggX
z4PKfB3xX8mmaQHpflEpsS2Jm/VndZpMmrl7mTW4PdzGOAUzD/1mM3fUNMkFfSf9rzaMtPsizaMO
4xvz0DJK+aVT7xJCzMGGmdfBPdn6zcdb1AQOxAN7eqACN0wQ/q6m4aPevVn1SbYZo4GXTkAqotTt
Eha94CHxGoFdsyZotzmki1LIkl1ob+9T92kxi1aDp+j3pKgikcAEntq9UTuCHdBy2uH1gVeTTR1Q
jmysdP86ZCqH5AG7zGi1U/NR7Hg+OX6uueafiWYt4JhImKc6IiSRcde2KtKibvPvbmL0P8+7RvkI
Mc6N6C/rQAU+dsApyyPAduzD+zjFwxuX1UjVfQ4hTfo3vFxXrEu+xQfhc77W2tSH1puMv/K5EAlm
n/Bv7jDJo8E+P+D4G54Z25z48HbQlkS3x9Bs4lbCP6im62Qb+RYiLtD4MY++nsYCZYCNPz9HE7sa
bKDTvUI1Kc+i5a/QOyYO6KoHGvbbap1E8yzNWOv9COuE2Xj5/iZs1CX87srkP4sROhvFckztk4bB
lcTwRRYfPjy1K6zoE9m0Wa7+yU9LTOsIZitWmbRBw6YDGuHY3sErxjgNxJ7snWJRKwc5qxXkjDpK
QoaAVA68jiQSZH+9KhLiD1YR0kwCf+QWBBK8y9P0x3LKm1QoyKMDpkjtx3RDQAlfQgSl5IzV7xMr
c7H+t86kyMeKRvXNa54rQ90q+ltTTv3mJ36RVQEXN8DzgvtUPGtLAISxpsBXa+2UZvPCIskO1xW5
eUmn9CWienuHmlg6oSDt+JKdLFyM5DZMmInLxV58f8O3AZD3OfV+dzsdx4SsrQVF6OWLe393/FWk
+sPx0W0uRtA0JJTBTUH3JYrrYEDicOzS+j2d+y2JbcAmztyy9aZFhU72NhmRnExC7GTFf1ZwAkg+
fm+l0PMUmJmZAA8bg6aUstFMkLsYnEcIBCA3WMC9ILQmIIQqqdCyjlzhDmg4J+AngP3SL2sNWm9E
/gEZRHogMl9Ri7Xn2b92LXhWc1p3lAxCbAcFvTrbBfZXETv3IfCxlXaOLYZKVRFbYjZWzp/ek+6i
bBVKP8H/DjA8BgljxGd8fTmPmsxePVIVKlqhoGIfkBDQLeDCKU/pFfltcuPQ9sKqAb4CP7+UlUBg
/ZEUQp3TmOgOq/59w2Pr5h7k2h6CVTcV9VJUnNoRYxL0ns8fEJWneaBnno10xjPq0ShahS0v0pO7
jR7go2CBqgp4R89klUk8HuR6zhvNI8TszwZxQfyhGp1jH8HTQ9efl4lbYAKi8n0HwvOIn3WTiAoX
QiJ3t6VgEuDOQ8CWJWOu0SmpByyy7/e3uUAm5zk0llU0K8Yrst9novFMYdJjrjnaEGSoCXrUg/5t
E0tfOQCNeN/ErBskV06SLR+09N1t3RXReQIby4/Ug4QErWXt3oe66tcoNGc8AYaH0CEFRYDBKOuk
Vsk7Dv7v3EcEvSmNQP8PxRc9SNkr5xWndhU57PPPprmIpMTtVT0khcOu3pjOWG9hvG8sj0ZzeDh8
COesu+iQOh3pTKPEW0gcl+/9b+WsXMy6mv67ojbu0DrfU5S5WLz6Q7JwvXsK/HXNUy9DPw97WNuX
lPNTZmracyU4P1nmjgwSjn5yafZJ3yoy3fSsVrJqR6iqWFKJdadmWmlXKR2/CoVXhCl9bbO+X9u1
w9rpQoeqzJeATPSsANcrJXLEGyb3X09MV95DmtqkVPQa8zWs2amwrvlz9b/jGe02izk2Q5YOKIbV
jF+wH5cYahgrHr6W6VY/DnU6og0ddHkfFAEccq0GkixxK1u0rUw41RjD8KvWWpA8ZCTGoOIeqqIY
u+3/BtbRsiVegpXHFV1CJzfNSL56KgTxVWv4Yw6J8uVFkl7Abxrl7srj8KJLto2PBUqMJyL+TN7l
4vpmsqTitVWWdiDwExOx2kPV1J04VQEco6AQ3JotAMwCBwHOJ9uoDmhif9gVgE9iFm8S+JelaeBf
TEAbxICIXrlXOyJJTG35i8fBmHvpTBj0OokePdE1sVjz61zJu1VkvDQEmyOhPiIpBH6XmgVrgaRm
6oSiH9NPJZPDHGSCySPJvhu95R7DMqQ0KzCVWsXXn8iIiMwXUGFN5XI5u6M+R0XONno4arH9pfej
YL1zjFLXs0XYRWw16ZIqsqRf7CbXSi7eV5DrDtHoQE1ZqBHF/1MtOgXpmjF/lh4UE2fyc4n35zgx
WpegoVgA1QtRI8MpbW9DtIamRKm5glWnejSRy/b6gsaUqURmtg2z643r3krBWIV71kZ40pwRCCw3
F0Igv9iLfFTafEaWHcYlwgdBLd6mOFoswjLjv2Dzh7GDDJHd+MNKUNY1MU+NIJLnDHD4s29KrW2U
U2Y1WCVB0UZCDva/e0O11rOLKDMmopuQEcSN5vr3+5N/erR4txn0cmZMv9jPk4r71UuqL2Ofia0U
LrAUcnP+NNO/I+L2WUXS69aBrkMY13eQm7xz2WUAN6eEGcJT6fbgE/ZvN9mdubyIjXpAGkBrZBoW
1nU2yBn5aAAQXYZQsN5d9xOGH+lmJeVcgNKya3j8jKgvutK9W4cvi7u0gyI1vnQsRt/5YdLOwr/I
4/E3xXyLk//uoAawkSXPG4BpPWBUovd+/OMrtZ/h5R6yAVLf86Ez5qh/qWuS8pLfVhu+D4nqWUSy
2ZrXjkJM5SflwtlI6ptjUHItM29OWQRCY8a/VSqa4pL07hVlWprG6fQTpkbG2a9dao5RWwh/zgsQ
ojYrBGU08S1ch1RY/08UQ7Uj6YmT/hX+qMLST2RCUlS+C1OHp4DvJHFaXlTkvDqqyr2OwcZkWCgy
ksfGce8vMQ4HufYyttY0Ms8OMKJUBBZZ6ujkVe3lAI33x+p64qIF3P901l6gLWw1OOzLIl1IEdFx
rEbc/0fzxJBPEAQPWnyBvnukas7h4rZTsLcA6DJujxEPU8WscLGbHFjGp+EPOXsOsiSEYRZ6yyik
3flYYHV17vSw+7+jeoT4ZnZaXQd2A812DJgLPkySoB9SDwSF/M+9Pk+J3h3aMgpTJyP9TF9QBPgc
1brPToOtgw839SzqPLna89qKvOedUFnatszEWyUrNjpx969mPeW+iUqkwzQ/n6yr9Kfzc6x7egb0
ObQCVYGgj6byVN2KA/gBuGDuP1O2bq3yA6GgbzBWe4V3gSWNNBu9BMydRoBS5ilh4aBhue5XBCGy
x8OjkxLeLPJMtXibEeOyLfRjNZ9xGNNN54xexw1bIeieMdDU9lyStK3tiXU8P/wCnimgjTHmT3zJ
COc2j8mltdR0duc+OLjUmMfgyL2u9I8R5xqVx+3WFMt8MOGOueUcmNcrA/qRVlkHpb258tQe8tCx
OM90QnsVoR8UiWdK5Oyq5gnZH0KTaOnlW85xthydi25yyha2jcovrbeYo2anwzBV8+neab7SMkVr
3U0pvqC2a/pZXObe8RDmLfJ2zujwmxkiCGXxSoSP5ttAiDXIc7mtXvahPGajQLqLtkvK/BIxVNAx
qhaX5AsjUll8ossSBYEMgIYeNSbMepq9zaqlPQ6SxwSx3pHxUDUS8UMtnfjBIi1wcsKNbY7QhIjC
DdiHrU+v4bXGflwOGakvultL7l9Cz3/pj9r73Ne6YMpdG9bViCeUBkSvj7t8ryKiK2MAH0CE9IG7
8J912n43PYA0GvHCVjZ/fN7zu3lsa+vOFM5s8kSVpnN4XdOJYGs6C/r1di4G2BiymS/a5qIG1tE3
XmMunuygpOgmk9V8tpF3nqnz9f3YMrrTidXktedPAg4/5h2Qt0fCGm8wbZ+uVvMx6R5uBJ+3pCk3
ikcvUyH1XwhiHf1fWtnG+X+8dQ15mxCGc1fb+VaA4YCJtJkgC7GaCUwYvXo1Bu2a/CFGEPuX7T84
81IMlRUjY+Gov0DMOXRPKwIyuUAnB0EzzRk/TE/SRVKO7UuYnU+A0SkG/haoP37yvA/BNc/Ed9+A
72FDdSa7wtLj5XpKbsbWHUwY17MrNO/II1z/SxkhbvpyAOGmqCelZ3r4crwrxT0e11dcuWRZOq1b
KVRlVdMUTt1//6YjRAveinGCJymmI7hcT3DTHwzlyrpQQKOyuOBzbPr4X3nZp+duLlpWZaj7KHSl
6Ni+J0pzxtl8TpVjvPnsGaoHNco2VMSH8qi4itI2pcu3DE/3IRMwLqPsYzwDaogKDQyz3TYERnXv
vvdq52SibRIyo49gchlBALPKrPjzDXUrc1v8r9CUP09TV1lVnPUUIiCY7RGrILzSzWIR4dz9336q
EkyG7T4fwGJdswAh3V4HVavuk2gPDvfXrYfh/eDJZKI9/1WB1mi3i1SHiyba4yjk7cKUFOO8SRR8
4d9nAx+3GJW39/HKH8Fd3fQ6r0ff3o8y2Mk63fOszcW8B7yXtjTh7RxnAupJE/YG8m25iiOoeH/8
erIC2JP1pwzgwF5cWjsJ+CL3JaV88wTSu5KmR8pQvfNnGBFRgY+iD7Nf/eDPTxzjGylVCv1vb/ao
QcXrjvKDj/9VvunUuhvXGjL9NlL0ryZzrywTcqqIaQHCjXOoYqOinGhETkcQls3Ro5/oScOGApnL
I9ngNp3uKfnkUkMGhAHxcmYKpS+w1qinWWfDVsuGxrnaua3Wrg/TNb3VbJPkKO1OJUefwOdnJYsi
ex4rMZSnxk6OC2QwM2Z1oGxcpkAQeF0JLMkQWFhVENfnMTWLwa3KIAGVX9L7QILubdpv/Ex9lSKt
dbCat1luH/GBCi88Z96jt25Fv1UF34c3dLTc+HRXxeNwLDJXiStc9CpgqUdGWjzMc/x+ubV0agdw
MZ9ZATsXQzuYZ4nzWj4lA+xsFWgsk0InHTRpx6NIMMztpGzYarmU6E5cVU1PV2doKpJ/b12UJY7y
pGCxGDftGqVUUWS8LkaihIBCTvVhX5EpqeLXuAwMHsMigCZvQCrurADwfULmlBxRwVJgwjC43f3O
2Z0H3atXl7OEE8G/X+sZN3A6w5q9a1sPsWHAsgrnN1cLPyiquX9xhjO4aibkF+IGGNll5ccrU8ff
Br1iVC/Fn+x41/y2cOI/JGmiRQz2ZkuhrmQXUlIaatSjLUoQnTAaA54VAPNMWMNjQjBY0PO1c0Rb
5bF7sfwVlGbyzCN0ZF7GyWroMhDKUj02b6DEJmODaLb8aEGgnooLn7YdRupHgZmrWxrblogv7y9E
v/yrzjtXUBVf2882dA2Iqld3tATmz1rY894+7k7CwuGhfZMhDMRHl9oqjZ6hR6dT43Nfq1ABFUMz
1MAE13awhvxrZpI1tn+BK4hE1cecGdNUpqUbYE1XrPwJtN1cIiO60lb0Q0E4jj6MGgpFs7OWL+P6
YyWXmPMBy0xLj/+t0r64lLrXiuBTNv5k9vYL04ejqu9uwMks9pIPxCVSZs1ewZWhnNZsIxPwIJRw
8AufjpjWgGrvvMnoYjv7oijoe9E9QhaGs5h9qor+MBey8r/+lGg7ZK7QKcrysXj4k2cDtCx7O7OG
E2OQODdKZAjS5SMS/uGflWvpAkTYDh1xmAxgzQQ9fdH/SOhN04OabNQq2X6Sc10eyGA+f6Xqy+Ps
M/vaoAD1vf6TszlvdcYBZUT8V+4UEhzdtaqBV0qBMEoNEj9HcUz/Tc6+EFuknyMOwe14eE4a5QRT
tls23IIf6ogSTeelGYRYgfzfw5J58m9hUTuk+KsxXGlyPdv77M2dpHdfuD5HXrb2xF5iBDngjlkA
Z7zc4/f6+loL5fzEYYaRrwgdXFJ67Sat96qOidIvdoE5AqxyLppwuO6eWSex96djRXcwu2GG4sr+
V+xtoycEaaUYGW+ZJSpgz/AJg1hYVa6O3QRyNpnZH3FQ3AwPAaaDj+QZF5mPynQWzcLOWHclzcG1
WJmn5nXU2gHcg+n+Q98OWYVy85+10Qcx0MF3vA3WhynxUdDrrQFKgTL89aFC/MnfBrBGTdGGxP1r
6zbtU9qKBLUfRBt5/Z66yh5jEFqXk7iABD4w1n3dmZc9mGj2aFcFz5oNLI7m/Q7L2szrYXF3S6Hj
AHOXj3lrKe7+/o6ooP9p4WR+a8pdxoGTwjGmfuu8u92EkmZD8SDU/l1BXbzhTrAmS3yVy1/cqxmc
mOW/Lg1eHLSgguSFlwfe0l1Wu6xaBBdeRD1HZAMSKwjXH15FdDPnYsH37Iy0zP4+R1cyCh25v7fw
Zd0NKWUYgcrxmPwMY9tH7L+y2MvLPUGgljphYUFUMuliISGUP8oQcbGqyfhvy0blEYki7NYCZC/m
IVQZll8ONU1RbJdQR256/1V56Yec3BoVAifHRjxMc19CbQDNA50UtKBflDHSSOEnQHR9FwIDjBSs
UiJuDOyW3vDiuw013jtXsoBnqDwxIRgCUpc4bVHttP4jdI4RaI4Dz1AQnGRYG3YGb9RiRG59eL/s
PmvEdepikBLbMAaCbqxqEldrCC1Wa+aNoDoD3fkGhakc7sTO/bvsMtW4GCE9luVn8dQgISJo+jfx
PWJXY/pqrY0ymd9IclD+ehT0t9eVaQd1SK/wJw3vZXPG7Wz/U2lCQ/YqbjSxnaQyUoZ7rWsMyRV6
WVMZnrWfleaZ+Q5pxp31lqd3amLCxLamUXTJ3PoB404YwgtbzeFhyL449SeBXdnEyXrNa7eT1ZER
Rc0MSG3sas1HkgsUT9iMue2MyacPDceTuQ3V43J9kZWG797+qKqhBevDtqYggzjpbAs5Ps8ltK33
va+YbPYSH5pJzNZaGY2ydbV01brUAdR2WENpZJBjX8a2IOoTUxKdo8+DUq4pIVq1hJ8L/fr2QP+v
2K9cqJmMztcrQSYJqB/UH7TsUGUDlCzXlW40DzY7yclixUVTml6fLL9vDaE8ftzs02YgXJP9aVoP
9j0jIqYpkC5tU+nKv/c1ic6+D22BWp/lr3QRFzBA+3EOd/EAC5htEtYSKBmWMzDX2sudcbJhWlcd
koiWMJzy5bEoZgwYNYGgBi+OXLJzSQiKpnQK+Cx90sxdEaKlKRGwylBQLlW3+QW2sqjCfoisISrs
y8oexl2ri+X24DiHDpGvtMHypjUErEsF444fxB5xlj7bkQQnc22rG2UFD3ecUgG0G5+X2tuDQnv3
CXvGJnYWJI5UBXie3P5YA4MgRHMCRFdZ7hAsYDCLdMz2MbvUhd3I1d15kTpCb2thhJbMl23XZ+nU
1JHLIdi2MVdcBLkKg9G6pQB9btkQct9hPkUv55KtKzXsreqv/nLZGZwhBuD972HBqxvszPEnsD7h
2VSe5yE/hNzkob4hObqlj0gq9xtu11hngzL/nsR1sJ/1j7SbqLAo2Iz2BVM7bhfx0R/SRLS15Bdj
KIGRGVbKnopiCbGIywjIA/cZwdW+hSnewkj86n6nVw86cV2n3yp5g0wOIs8bZ/paSyQs37o5AYRD
oj1LwpIl3ns6SXfNVh8xhZBbAK0Xf/m9T1cU2QbWNo8GJpob5qNavP/2vLCd4CEce+itQas0c8P9
KaYpWMKr+FXL3ibXXwGRXJRBVrYrcrYBO/kF4lU+EX1XlTkZfgum+SY6KAE7kpN+JqU30bkzvWE4
igTLRd9YOeEdVAwPmzb8mhjIbEHWBrpksWgx5ciQJPLc33SBP6VLjYotunEnq85BKMJnxDkmEVB9
+XNCRhiOSdyzIDjlgpsVsPgkmgLo96j0OvX9WBhPb54C5e2Pm6vbhS7JakO+tMyaQjy9fbLmM85Z
kuNzCgB80AuixcZHwnANN1kJM/O9v8A5Q0BIlOdeQoP3FkEoe9qusyIuPpe2cirZZ7fVROd5GjlC
gcCjUCFXlxAQPoux0R/8uJXHvIoMtLt+0Kv5R4l/ODQiJP9VXUBBNr2S0x65jU6gLj1Ro15tdpwC
6kRst3h8hr106f6deO2fgdag55BpCCalgQ71k1Dkvs2d06jOrokA3M6R53F30ElxXAHeaEHA4TMf
gKqfbhxX6YCll/EkMD4PBsQmx5KeBbX69q+v+uK9EkTXOUjv/cVZGC1V0BvFiXLoZQe7xNGtniSS
yc2cKGASuVABUs3DadvdcwuAXQyI4nxOpLeHsvJCRzL2SxR6ENPOl9vUNctbm9UUGhuvEe8l5aER
725EnX3h1RAAEILFwOSzDTVZzK2RDWvKyQNS+UGKy6mBByMTbAYbADP7sft3HAE2yxNlDhxxQe7k
xSruJcQhgeUfEFi9vQDyWeSFdK3wxoGMk9voaQS2xMpVn+XV3Q732KgtOVvsQxNP6yjo2ctGiVE4
AdOaMvSbWHstkyeRcoW1t5wcTwnuPuxcFM6u7TMITtPYKliJXUguYFlKeZ/XL0izaHdjcKHN/XXL
3wbMyxnhPNQs8PgtxoZ5HK5f1BXtrYBmOYAPI/5pXzkPevnSsOa3prQb7/fKkRyhO9WbNvmfxIu+
zNnWTEP8vxtPBRu+RwerqQgSTevxz3DJmuSjMe/OjC64yCKDZiOSK+wSuVqc3IVWStxjEOKR3XlG
n+g0P3QyLf+bsS9BQyIDhTT2k828hrodPOXAd4DiMP6FrmTAhNVvGAS7P7dbwikc6aYOP1F/SUax
NbF2z3hc/WOy+tG0AomCFaTqvqCeGOeS9GKMYyWU6pwKjFH2xr/0quAd+f/rbp9d4sgz28kwSxyf
vUo7oNpVOuue9dYxEJKpEi+hlSyfP55U53EgmagIbkJQC5391xnd3yHIYNM89rAHzWN/92jKtnXI
KrMxlOtQFl8J62cE5NuwEk9UTdKCHaaQpMeYOtNxfdN6fklY91jNSjhjBDYI+8JZZtBGfHEp3+8o
Itg/OKZ/jBeSah+tZgg8q1eBeT9x2iXS5gL5S6czs6ig1ry+IKVqJPJ288B8GCmTxMr7HVXGPWPU
ZUnHRsUkRwd7K5eeKnCLuRgg2XFtuzGYVEzchYFBXhwlkQMI7s5Jfp90q+SfSesCIC9ZU6G4VNOe
Qo+D4B90qzz7yW/Bs82cVW1yi4f6XZIXqBWXE9qaEsQmoUuxvj9Mw6GAiTiAvzEstRjeHIYcH0q4
PCMCjdyvO55e5YZti2/TPDq0eo0di3/QJC2NoVAgPqNlxSfNqoCR0RsEN99fFE3cF0nt51FFG3+I
DMPTLvE2FSGe6vBbflcoBfSKG5DQM5mVdRIy0bOSgl8G60iVsrYL2jcLT4WxhZX2KJZzERVZSmx+
MlDqUG0pugmQerSaO262QBuO2+0aFJwQAG6eFvgdAn2lQQu8gP8EO5fFNKflmj5GBcN7GZkTCPCs
eri2sc+NXFzqVIpFN9iAgt53tEZATll4BndZ45TbgyCDLnkHF/Ed+8vjas6e1VxnMogMzZXgJ6im
ANK0lvqtgCQrJz/JyodsHyu4z/0VcR7kD38qFU40DDZylyquj0VmZBxCa92VSmyEmscf9pRdQjHb
tELpl5GX5tdKHHAPYnWudeDxoiCqzqrlz/Ui7X4EksasqPrPmLT+vKQaHynp7nilIE1/sda/bfKG
UlWM6wNaMWbx2yXoumu1AGuddYU3/Q+ggCGvm+0xC5y7sC05nKR+CGMa0XQWwnZKb3Qmz3S+ZgBw
FwyuEpQRFbs9clARwebbW6QM1fyHU1Pe3nrZRNLn8Y3rRFIUWJr54gu6QXa0CbistQvDa+1ANX3C
AhqjPe0GKEBQHFTXqM1Z4kMvWbxbR1YefC2E1x8D+I6mNa1eiRXJGQYoPOcEI7EEWGjUgLYhMWGT
mXQphQt1cDKYWZB/w+uhbf8LkgMLDKw6JmolxayefCY2aMLh7S/8A+KiPGF3fjwnNRlx3bff3or7
vrVBTTaALT6S3iooJjPxBXHeFOTpJtL5LX0XoP1ZdreiA56Fq+Ieg6r/30tZn9oRN9otxBFJlgUd
PDPnE6ZqZCGW/5Fox5RU72ToPkwtItszsw9mdI7qeG5AqVUVoVgZUivCGisOOWi7wSMFyQrvxsrs
Dq+F1s/ogaPgZxkyZ/Pnlgzji2H6+qursuLc3aOkOGzRY745OuwykHCXVs46KzezPk74toTB/LG/
brJNnzp5q4MsOBYOk99VmavLqAtqURcSNXMj9lb/ttrH+a7TMZWK1NvB2G/Ea7M0vkscMiWjCJOZ
vEt94eo0P6xnzyq3l+7XqbpIjuXOex+InzVKn6bBptQNA1wgCE8KTxZNFMncfB7huplnUDfVrHW1
3YPWgMUn9QVkfLlTQd5amza5tG6noktB1zMRFN/NGEkrT6tjgkxiHUeme+Yp638lC14a60EMElBn
Ts5Mu4Ab3PQyJ9xsUEKnyPmjiH3Yjjm9HhKA2SYxXeXpPYQ9ejUUaAeMOwcG2z0icuw06usx5kC6
zplyng4nsTFESOrqL7MKGFQnE9NEb57jPnqRr+tI7VZnA8Rsgc3hySWcu1pxNPw4QKdxtTYxrM31
osU1neYwuuXBo8TkSlaoLZ4FAshdhc5fKGrLrwZrn2pqpuP3b//1gGtJTr7xI35rgGIaz3/ZKITs
OMzX9Ko7o31bWRiGFuj8C9uCoQgXDJ2DIPED3nO33cksx0EVFtDTdEJs+4AkQt36XQpVX7W6Gdrd
c22d9CTcG6w8HSvzwUcZNKeK1/T+9azNNJUSU0s3UkJwRbxclZ9oqfdSbPmH//mTGADPw4j/0IsO
ZmidIP1/4wy6wvnS7r0KtBCvy+hZ8mMTUG1Rvr+FqxkTamnAKkTewkhgQnNTriC9NZ4oYoBtAXuT
XO6QVkBLHJrc1XPBfseRM+7PcONAfHyY6W2F+BUn8o0aQP22CcIc1uVhidkyvHwZG6G5Lyw3vXgk
bJtz0TYEGK6hvqBJKuHIu2KUgu7pxJLjAfZ2trwfSDdRHPtQy6Q5JM0F4ts3CTbFuHi/THTjVEZq
+84LA95qFIAtvowEvPvZhHm0+y5Vr3HURGWJfkT0fGeTtlckO4U6tWsKQR22yJx1ncyUZh7M2vX0
I2NiR+dyL5SEtcEMAYeYAEExMmABCmmxAW8oYaMqw3Zrh9/o6022c1xFIRGdcXZH5UqVgmB6DFM/
c6jCcec7NBjtRUL4A7Pn/xnBQSzbOicBwGEuyJRVE0RbUs0GV71FaxqfGOLLnMEcGAAm8TcAhkAC
FoluYenZ6ANGBRYcEJsSB5+e2FmzFvgPG6uXjfFrKZiQ1KA/y7qzX8qqkca+XI885GkLury53pN3
KbJt2/dtnkpAObSTde1O8J0pW3mLKlMeNmLL4OVTGNLHbtLxIFDUmO6Tordl12NKUWUHhROe6EW9
u9zEIwszl/EocEI6n5w7SHEBclKP1GoPtgEFX+I6NLl8cJrKeqCfYqGkg+zPb/l7YLs+BvQbnzIX
Z21guDr9nUHsCREpmOEKOM3AAvOxpv/nySgQpqSjrPGvgOG1DgiwA9Gf/yjusF8xsK9MKtrJlFv1
Wk3h+Dboq3uXdOrQAPYqvALFma/gkeIivwE68I7OhfUWUIGJB9TQi3/thd34LqJx4UQB5vC5tYYY
k4FkjfYgL5M0xHPNWas7xUdq9ccftp+fqdVCLJYl2uZzmVmBMBCjB4SpUHk0/XBlM2uK0iA4wmNx
dR3KFjNBukFT0VRl4RrgCQVZDYJR88t62piOYQimjFyZOP/+/dCxG7LabP5OeWOhydmstyzK3V+E
ZaHd057xKMR9/nzdZt5osC0ccY95HEt9E3rKGUF3KP4JEWHG4oPjo43RX+4UqPBj1CauJgGuPdWa
AZKjgs+EQ3LZShRCsA02yeX9KyQU0aDm06sqvwQR6Wx7Pa41NYG39PyrN+91T3KfMWeZ44NzM3E1
2c7mJ/eTtygLSbB+3JOGJkOyw7AJJN+B7ezVqwB5Gpdz9DYGgwLSpF/fUyVB1ZGkiH7pTdE+Mguh
8dbb5YI3zxNevgtr46tMgFC/ETD3HpI0karjU4mgktKou2HD0UFEdgEoctgrnR4hTbiC3ZcYNBZo
TjQLEEAbA4KjkXtYIEkq9pRjQpp6NJMxKyXTDZpQCZAAnG7KeASQGVRic4GA3v9iiPU+5bSCK6X+
BgiiE0HODULIhktoaR0J/8c61ULoIdhq3HJhJcmIdc96J7XJT7M8V4XeQMDUZdWI13IJ+WBRrC0A
v1sOKvYfJV3+tyxWp/OJ60jREEmfrz3DSnbiD+y60uE3aLzL+rv7kO0BOT6HIv3cqjSDQDvihnDA
B3ie7+VGsLKWLsI49C3G5rLs4rhSAtXRpyMIuhqTxtI7HEEDZwSv5cTiXIEMYjURIb8QZQXknOdh
qAycT+oSeMFP37m5/cyP9Or90OshHz5SrwZsUU5FmdT5xXNt50H6vOE3MVHuU/LuCrzcsGpDv8nY
JcNfhvMpy5rNtk5uTI/QdqyP5fc5mC9I7UtQYXlWGCucum52sEeKbCWyVp+xmmQqVk3WwlLq7Rpz
DKXx4nzPKdGSDOSCci77sZQ1c2bJs/7GKy9J+tb8VTBxmuA813znXqPjxy3MdCg/MJTrbwJMgsHN
fcnYqVtc4ao/GhP2WSIiHUq4N32UcL9SwuOwYUVAwSPQz0nlIRafg/gdHku483jTDMWFG+lBq5oq
lW3+QMCwztr2u3UEdPYhHo/FYJlBljPtCEGZGboLUSh5we7WkG6fK96Gzy6iFBAj/TXqZE5qq3cn
ZajV/qDhaGnuw5jtpmBkQiRzMtI+KGoAFH/o5qD8ExpR9G5qqo58e1Ad5GHPHjPUWY0YjitGE2j9
l/3eBqD9IpiamqHMGJID9Rq2TP3Z9zsIY6jvtwjR9MNhq0WiwPrBubATV8VUVIha+IqFBANsN0U9
qJqsUgoCWxSWMOXATm2Nh6sr+50ZMrKJBMNRPIkIJIxRW95x00mVMlrXA/Xc16N+x4Hw0SghOAhN
KcFAXV7qZttqCYDyiDSEubJBGVXJc46IigQsuRcet/NU1bznIb1qfpnyJCrnX2pqt4hVaImfCUKK
ET9DXq2PY6/i5731w7/MRN1v0TQ5VPtM9zeYPoZjoA7wOtZpIV7YVN74O9D9uUIfS8Y3U74l7Ktr
6PzIC6jf+eYw6+CIiw9VwATiOQi1vMEjLpzkZFqCfWP7np0vPYLCNOzzG8LjNDs7FQ1sUqhZ3jpk
eeaRFU2gAHpVGVR3s6eQQgQo6MeNzXobqPAAJ5UbcmEUX8QcZ3WOEv2w3H16yR26BjYF7Sb4/RH9
cooeNUQglG5K4S5P7EoMAuLa8OUngrojK46fMzVXHM+hCXSlTbgG4qGaWTUxUQ7ep8cQ+U19t7M3
C2tVdqa4ezp/p97d8k0C9YaVZBx0Dj9BJGpsXoHl2YgLbiQvx67xOb6cO0mnHKk+ugClMzIzdTrx
hd9KBS4SlXzH22X2qu7hBlktDfow1dRVIahEIAA41VA5KeNgxzYz+S5NU85W7o/vN7iMVygoom4m
9L58Y68kygh/77+dohxfqke04+SbO54F56mRF/mb8hbE0UCi6SX1n+/NAn0Y2Z8QbfSOgracKebY
7XGwA0WRRemdBWUkor43TuOF52/sexujVaTdLYjy97hi3REgNIzxM3sxGQyKzRJzP9YQ+hbGNZA2
W+hQAtQgPmCu3T0ctDlvROrsSS3m3kDuGxXGXBFPaduRmMV888aqPpGuKWpqvagnSB179Nj9aIbu
JxiTd9MsAo/56mBsCOVjVEPaWfGyEc4JiS4YBskj5Zz9+D57lQxZrJ5fwqfDnd5lMUE9W3EXCCo4
JxGeK83Mu8RmdXim9OgFxpH6Kqt0AObix0BeWTeekyENIy0d3SD6rClbFAIf/X0caxd/JiPcsSCy
fyLjXJX7uE8RLt7i7jJnAh3CLLtHmovGJG3aVLgz6Qda9Pf9ByGHC2RWkO6ZiU2NySc/q5dZoidi
Bnqm9JYLXns3EYDtG8LSdb6zulUE5yyVy+9av3wMORtbZU6ji9jlfG9P50Rl0i9Oqw19txYPvLHv
Neq/2FjrN0YyqusoVwbeQaIuUvwd+0cQj5YWKGVzVlAdERFfxGS55EMASzwXTJMhpIwE5tesaP7i
muixcWVZPQQh3grt+cN9QveRd4RKqzXOkqU9hDMXGNNGvR2lOgYb/xYnBtJR+Bmh1u7iXyodK4BJ
alkBca9TxjEtRfEGaE8kzhw2Asus/iKTOoyFEnI9ICp4ppIw3fa4sFjkZc+e+oMl5NjS2DlCNGxY
LyLVfKa2PMimw3B9BUcj8W7bLTGQStAifG4I5v/ld7hxmhVW8X9ENrP9p9T/QY2qfqCR0K7egiVH
LIjpUjYQS98ueCiDv0HObAY42LbhVGcVE+/aBJ4IiM8GWqxVZu0fym1euuMER5lHPgF54rYdk4en
Z8o0CAuWZKyXrDesxk8yX9V8YqQr8qyCS1bfvpijWeh+8gGmlDqUFv8QUR8P+TJh7BALNDV8Qetg
+9mVlKhfhZhOLI/gfvPCp8WHmyE3IKc6pDR8ax0Aocb3G0xYcGuK4YN8D7qP0g8oDep65Pe94Uxm
sg4Su7sWSNTwCCifqnLhvhFCWBfjQ8WlZ7wubufzxJPPtK6OmSD8NxuFwPGV+Rv0pVq/o6Q+YqRr
y+iU7u8HTKnTFF07WLUgMidaPvU2iqvuyXUGQmpzEc9elYzDGW8r3qU+euvcM+rNv4vQnJ3B5C7a
ceaHM6++ic75/mOAFgVXgR0t0KaJHNSrfz6GGfMmD+VBEtGO6EDtcUXWayjz9+EJ1N8sEy7Q7v2C
w4k8vqmPwDydco9oMvZcO0Sh4eHcD12c2eCNAmQqpEQP8zawYaFiSgxBiDDoeJUFotx8Yc8vOz8I
dB2kx2m6wwFwaJr3z/hS+Z1Nxrp1mQ3nrJxZVw31dnBOFqMZaoNu1nSWzfZynJeKF8ASC4h4bRBl
x04lwS7UVmWOVbS+7b+nNaqpAyOlnAKcwyi5tspl1Zzvh25qzDNvSOVQSHNwx5IzKMQ806tNXrhs
+KfXQ0DJ4h7SElHAg76NFW2M0fBlh89rDtSax0SnaVWPVkViGfY4kuCc2iwwJJE7jdE5mOivBO0O
vR/zmwKHLYQJqm6fIMVVxfDBJIq+VTWS3FrNL9poS7rr7oMZmCeUrnaRVep9xm2RbVFGh7qIddeg
clHbexYBSKJSE0VAISsiIILqp1vxqWkPxUanNPkVqdbOmWxuSXX09yfKTO+iupeN7be+fqdkg/eh
fa2imwM5nYjvjk1db7b8FXGysgSV/jssua+HKiurcpbMlnCBMjYcrbBdL/Hbrhh0OxECg0bKZ3RK
p2kIp8LrKYdB3Ryqyd7r+aOhUzqH7hyAZMroQRfoEijbLqMH/1WutTHQQfMMvgrx07oCuZ/FLPDH
qML8HgIq5Fpd+xNw1nm15gATaoFr+cZgZsdBAjnDD2HIePckBhxTRYu9//NS/usM7wAG43pf2Anu
Yvoq6pLwDe8P/z4adiCK8oGTZJzHzQLThtqoYLwY2Cy0i26glTgmcEbRLY2f+Y0FspjifOIsMgoL
b2HjRaAP20piF06RyWskHOhx1NQZ5OEigtS2UzFB9HDvr9ofobhLlAwiXpZUwLGzglxPXySCS/RN
R0fTXUBnwPtpslDsbCzKne0COE2yp5a+dQYlmmn8y8P1wuzg4k7dFTr3+RFCijv901lRTZr83QmK
+pGtqefVTmuevmrRg756T5rB7FAjbHVfZTdGWWjW/ucfNn5HwCQXcHdckxLfmRoGlPskkjlyrltR
YnsmL7wLiHA6ysKz1vPKrh5IN6k6lj7qCcO9rKCFAS08/huH+ZphFoobuOgOloEVENGz6UFv6vnh
GuqFlB83sncDtcfUpLKQfPzfne8/Uqo+5komBTvHMuSMWI9J/FEmpMsBoStfdXcn6Bz7lu0nXC/D
cUfN/Ej4gcPvta7gcglLCwaNss1CBRuUVkg9KW3VzQPFaeqspXHOszTNml+BaNa+/WGOn8gMLlTD
enrs0t2VMACLTJGm67vs0UJ9eQ02AlXVTBMP4PCdJ3dwVEFzoDX1/A8N8otDHd19Er2t8c6Ro/4A
DFwnPXia/bMg6YAq7NydzswlrZ+n7TQNYlSKupAJA1wxGecfe/q5u9zJwrvZri2k9xtzKtlzBZVn
OQjobRQRQl2KPHPHZCc7JPZDdDqIJdMuJMmVwx+3L1VoeXo9xaqiosL54nfAZLOZJN5LpzetNACx
ALb9DJnNCN6Mb8pzpWlISxUoGslycqie4NTQctzcRxUPnNMZrCfE6J8XYOhREvYMdxWNoI6JvsxA
ztU97MeBVrZZOTGe2AXnDB0Cy99amILLJmWJOntcF2zKkC0UqjlV2FAgEajQrJWhEdzC3dbpoPD9
L9UDkUbrK45GMESb9oHnFvg3Lb8hSoWPvg8WmgnaNaIoB9YswEaziIFXltmsUVhiTHTHk1+NCKFx
W08rjFlT/+mrXDvGYGIu/b+37Gj0d+5XE66GOgP+dClPLemOhYNnDV8ukwfyyOHC8fjtPzmo6MfL
4jjfobWJS8TpoAYBTJAVlTHcwMCLlCAPFT3y2ujsYluYQiPg7mzgJXnWZ8xmbzZP1SZulsX83RFU
R8ygUMEitd9V+2Gu8YgCVRPMkD8gF0+1YLi6KGdaRcbpTazWElvL3mEsuLNjom0hGoEPTr7nGDM3
B6q729B4JMHMvNp7l49lte43vFF+pAQ8rGd6qC1sM0YJh/o8ZU33Hh1MQ5V6a+BC6CPKHLdYLTgp
8O+c7qPBNfkb+RTGuJ/et3L5yYHCChEfgG3KAtBqTOqW2fkwXNay3n3RobX33ls17Z+KtnRACxMJ
5XErldzUAyUeCIcSXRq87KIby8TbHhKXGOeBZsez+tfCGs17aABVJewVCcu6M6n1nHbxte6iXqPH
F3+uJVADRRhmmfwXMsxl2zaxmNdlJNgoxAA8HTmqQSS8rxUfYtg0MgF7jrCrs7dsGkRfsMx1TVEr
NAebpucKKEJw0NS3NyymQ2Db09aw3xpJJd9iXQzAX8pebzHF3jswD0NbNGVq8+lmdAPrIg+rhIAV
O9420yPKi3iT24kD5ML447zHkwjlWRR/fVwOpAJ+7o3nzo5UuzWodHv6gud0EYmJIEOUgdpDq+vk
q+dj7TtwFt6avrXlw8kHBRDkd7KVsr37snefaF898ROxLVo2EKJJvmZhIHKGTMmetmJjvJlmPHhh
HRuefe1du7C81R6O63h6idWE9ceH+qjwDzpBEoLlo8xK8aZ7cRRd2yVGNJ4o1Cl3BnEHzgJ45483
zz1OZqP6BAaILDGmtCxzwX2HgbHt6tgCyQY5pc3gMDa5T5VvkZia5TiDKHCRbjxouiT0pf8CXX2O
+lyywK1yKITRbkyNy7YCpdnWuz3Yo2tXPNGHJ19Fg57eckinik+DU7vrygL/QizrnJcuV8B16F0u
p1JGOSch5v3cHArx8iTz/01vuVCvYpUi3hRIftGeRpyMCF1XJAfKHzLaCSVIol2fvqPCDtZI4W9W
u2Hsb0oIMgo+FdbodMjNvht7Q+ji+4nxq2uxCGMoX9o4jJVwyYKgET30BR7T0UBLWKx6i0lUSKkW
fHDeP04/JB4YJp4YEWqtdsS3h9m2XwAP4pa22XD4k9pR68s1skuKOLnUcHYl8ubhopdcfRIxs/RM
f5N0fCUGTvEFoRhDXFAnftjNANayHQb4wBNPc8HV1NzJcFoWnfIHP65OcQpmf54C76b3VSH+S7XI
nafKvyYVKiEumd8kR4PC8+ZuAPVMvOZPeJhLWBDd6tykM60q4vUP9k6sGcKkESzMqjpjI9aEkDAT
t1jPZaUu+Tgw9TYZ29yfZutOcOCAPReTKCGIA9/s8xqf2fo4u3g7rv1G7KEcdr/rGGXPWdoDgtPp
BjF9tQvH8TtAaGyeSCJy34NlS8mLSCvwAjFBunvGYP/D67AkF6pyUYC2Am6hSRBtnIDLBGdg/qxe
p25/l12UmTOlRNtBS5ivP9ML9t2PUvt7Tu6rqzztUu4Prz1YjJ1w+U6neTDyfUjOwje/Oup9po36
b6pFVPlGRdcULd/QVY/Sze8HV6JW9iz72fCi2sON0ZP8DtHE+DkiQp7d7lcJntlj9u1JuHroisYj
hQ6antZ1gXO1DQAA7AZVRK9iLbNuXgq/uibidpOEd6P5PNkFnzAMA3h0UmtPNQnSEvkrkN1PXgud
WCFRqE541z54kAEET/8T2ToTVMrMPwIJ8KqOfUN0RXXSVZ+QuWwkJKu+Jr6ZfFBXF+KiodSPe/Gm
NoZn7S6ZYoAEVme3aBELu4JiGApyKng3f65zN16hoH6tQuUGnFBr0Wulsm/ZfvLnKhk1rJDRjqGR
ZLxgbPEOux9OrrL2C4wQnnl85ILm57MDE73IVzbYY/i00MJjSm2DLzt6eeDKKGAayQ0TW9PufY30
HuvBJ9vHFRLWYY00pfPq8ZECJLTQjbr+nIRKzvqG8kf3W9pf9A9R0Xefb43P6NMp7LngHEP5C7vq
6C1Ic+uwobEBG7Qmx/N82pidwkoWl68uFNfRwGkphEAUfUIM9z1Fu1M6oAaqDC686MMXnb6aW8jv
P/z1zGKHPLlgFdx6Zs1Jdeo9I7jE05RtDY7AblWqBvwx78/8F+CrrD4YkaCE06NKxwF0ZBEGal1q
UunQtHnC/VxROQYoSY/kw7hlmmQau0SQ+mT2JDOI8tMt5dcl2xjRvcApDfJMnF6VMTbjDbm94f+e
HyiUHkxfegftx0nOYnWjGSm+7VepVWwx9Lvjhfct9b5MekEsKg6e89K/MbIcIKy7e3ccb8MTAiCF
T5ikqMcRmgdEBmWpL3kxwfSPieHz5uul3vj8pSj4tAus3VGlFF+vynbMLRubb3Ijgwx++ssIRjvT
YG6PF8IlJ8t+I/DL+obstsC7/BOJyFkoWpApkRsr2CQYxPraoGBjnl6Uh7aSIzzrl0yN2lSvZPO8
e/fczqlYvqdLx5HYHvgWyxMAJKOLXtC6VgGAbfFkZesDyrFuzDO0yhyRLVpnIDnrMuV9gMfHpkNt
LDtZ59e3V5i4L5xpcPqjbQjSeFXXC8lUXMSDjX4J+l23N/tSDto5HX4GoZpTqBLitdlKbpse12Yc
+/xw7mvjjrHYrYwR43mjap3uxGJpqRY9j1L1PrMTktYGjNsNhmiLYXqMtVgcWarXx9ok5EHg7QeO
8TVkIZFAxeHj8UG3OjH/aLpZv7aXl1rQzVo3Z90qr/b7CB+86cbR7iMsEOXSqJ6dYkhGj/ulsk2D
qualPzhF7AhbrVytSMm7sygLQ89PqNYGLp/I8mOd7NsA1s+pDP2ExnD2wV3UA6LcsRRLlK3+PvmU
taO5XSMAqm6nejVDnX0RIbbWy7vfH/qjsOsayK935YRyW2DXSlHQ0ujpBXZUfWIxhLurJtjuKtJu
2ClYoqeOnQu3KGU8Iz8QHrOVhEkoQvJKB+LqoJ/WoZ4AYR6pn/DGNuQA9Jx0x/LH7XAvesBJZ/JH
66C/JJLDjQ7uZcXHIsxnxRWaJe7IAet/02ya6HRf3XGca0UFzfbk7WJ8ofZ8v+le8VTeahoc0GGn
/udi4kHZWRb8hjy1IC6B0b0zLXEr5ASUl+fDDNdmVr2iDO94XuPqhljLzO9C9WfawZxhklArx5bx
0BesbDdCEDVH1BT6u1N96jS8Wav+i8dsVqLVDrUytMdfYcZowheouh/t9nkNxycl98P0NbJygtWI
B3PwEiA9tkF4WEqL5vYhen9f69XS42OQg31tL5duQlJKEYN33hqIIh1rDobXHAKevC8FrIv9L5Yn
vWIwkCQLhPEQpuqVjXsZ+ijlFWIjKNutl7fivZlFD42YHIBLZH9Gx9CTUN8UD/sfuQ36t/FzWJ+i
tJwffKhvAdIaNs9hsq6PrURXR8CU3dEYQJ84mgCZpt/4osmXnvKHxPrsIhGwlNENE19C3uWZt8P5
WGETCFp77QLbW4SC6yUi11VTiypk8zAlekrInni3mJZTUN9AdJRvvBO1DedenbF+1jUWMz+LuWXa
mdXN8PV+IRmqiqAhZvUoUhb2zirUpj2NEQwD5VfyZNOeXvB/PNERcKV5r0E+x9G4TfVfS8c+FmV/
xkJKJpZX7pQ5x2mxTQTHo/F4ts0ElJElI2r9QNFTIQgoE+PG+GCfMUjHuQ146PZGuKOM1lmRGsAc
xQ+YP5l+gcsWmRwZWf9MvSIJZI1ZnpCworFhiDYgvFblVA4geKEJPtcfYE0/Y/rn5GfwY9gKOtRf
S2OaClTrzvcoKFOoeXj1T3Wy8weAslmKYfAjHd1/pDL1DbpF5zOFfiCBpq1jjsVzbfZ96OpRIWWZ
3F9nzoPX0XkeVndqbKRl2FB05ob3ERmB8XOhYo6ZWxS8M4pcfZ4FPEumnCmEphXcQiujtI4tb7/c
eXF9DAN2vcFHSekjj+xlvAeZrnqSlAXCx/oluy2qMcDqbYdCADGmUuiRJk1e7+UA5M+hpc9Uet7s
mXq9JZKcALL30SAM0DXc9lmb4K0bevonRSssdS912sPTDo6VEFsuBez3eK5Nt3LiRLikgnOCyDEE
Fiwm/mjsY62W6AQcscuZ05QzN3TgKMEf3ixnpf64RRbh1GF8k1A1LC1nWJ8T87H+AjsdQlxVABnZ
qlei91ruk8NByU3m1eTJo03rHjaisVO1eC0P0s+snIiOW8K5QTYkfqCy+0KotBTPx5XhEo/cvSMJ
+flh1KnTgqhRQbX7YvI+ljObgY0bgjOB58h4/i5YYrh91aCdb3cGcAEWhKVxKFa8YqA5Cw05d0zL
E/F8jzoSAj071j1qAoP3XNXzMIDQpH5qC4AllLF59FRBn4qe4iwham0I2sQxxD2gFL18fVJgAqYR
sJnVY228N8rtgxCjXawTvqZAviMcG+fnS0556roj0P1npuEzbPfWWz4hho0xKogJWnB979eHinR2
UTx4oGMhaM4gomNEtrwoBLisUW9Yt+6euZ7ti9yaxEC21TfdlZPbxEo3W640KWOdBCgZtN4oe6r5
GWP1y9yjx4hFNh9Jv4UMCSUKNoqRB7yqUM8EgfLvmsS96OLWuQiB1qfpw2ovzbTbjuzyoVKfzmYl
/2Tvbq1+pNdDoT1HUbqVWTFF+l64WopaK1gvjPgkVv62VtZFe37PWXfFkFAHlCnpJCMo/GgUoCC/
dByk07wO722RgQcXn3TbrkhrwNUewF2TBskVhAYzh0LdBDHipPJtrZlWAWJTSPKB7wABxoOUJ0MZ
U3toigGPM4LQHK7J0qFknrKIFIB49iEWHU2HUwCW9Ir/cK6Ed4oKrDAqAGWE1tqYF7W5fye2kzeL
T8Gk+G8Q++zePsPmjQP/8UJw+bSNSOtauSXO9QdTv/vJLR3AQKG0y61pomWC90uGrJu0yfxRGFBS
0RoWm9IDEc86BESWv5kzvK32mo6BDg6drlU33ZtLMYh7x6sPIH8baLdT6N8hoIqBOGUFjtbqVF12
vW9UwMsHMIQXN1wJ6Y9DNSSn7skWRbCBJ98CBQsocvo91ldnWz1i00N6iWmSPsLJHNpcfePhsAME
+5hpEyTCxQfSJ6N297LTan1bCBsOgsgxbFTgDWNue1pvkNuXAh1UrdY2JU0YVxbKTU2tAQArW9fD
3Kin9N8j+ih4RZYhcntdg3P03iUSIetX94qfun/XWIHRd36J6xNdQ6W7a+LEWd0qTciKSbW7JySV
6+jl1GPTu+qCc12teqd8c0Q1ph40XwMwWwZ3sdwlbWw6u3qEPA5/gyBjCdXy37Cu34vZcz6Hf23t
cWC8n3wfK+WGg3pVwZlZ38Sar1LOxfCS/ZJbBqp2/dE0y8qdXJa3HYNyA0XpM2LwAodJF5V6nWZ9
aPsTbgxgt3VEP02xhsfK6436iovO0RzuAETlJuV6aHIRjyOOK9qmbQkpEMsTgA/8tlwm+E7cLpEY
Au3X1HLpPAyzSfGklcjyzmWa7HtLwGVqqzQATRZOIiv/PPNXnBxGD2kVTSJ86s/xa2lHm5WT/eNy
IUGu3YWByZOrW27t72Ofl/H8cwHcTaI/T8Bfj+WFjC497UgG3SdDja9+QQnfZlB61jatDSY3oURf
YUYAIXRWyHlpH4mxZV4zzHPrL0ttJFyOw+RSGC0VashFCl/6LUKOqduRe4kjXI1OnSWNtTS7Oemk
gBYGRsAIm2fcv5bHWTygYZQqeVxbLGf7RZPvqM8dffrwsK5qBHIHHnjzZtTrTkuamuXd477uXpEc
Olcv3O9LmhCT7AIw2vXUD9eh7nS9ixLtOJDg/XRD+LwcFd3UgNy9LfICm9ZqQ1aSS7aNfl7yxx9R
2QRA+j4Al/OrMvJVE406XefjaKyawcw/IANY5fD3W5UfL/ZjOOMMmN+h0ZmBTyh+DrPdvMG5vs2P
mmw4USjFEOL+C5mps3OEQ+Dbr2TXzgAXF/zJTzdMPUB0B50VXN8Y6W3kEiULdaJtUC/bWA4rhkjY
egK2H56Y2I/Pad6sEzqfWR5VYpfO7NPLpK4KHmc9nj6ZRkaTXmIbQpbnl1Pv+x4oeSvoMw136BYk
TSA/KnsSwVbKTXWVruvQ6+n/gF9Ff3iVaJOR7WHR1AlCzQxs9odYEx1qX4eL9ubWAoxZajfkSPuC
MJDMG9prPuEklaHVIPRkWbBpfiboyIGJVMBK2Ig+RB6Qel9YzO47UnVw9f07FWfDBES08IGajzMu
fLhwahrdBU7g/uAynlIkTwXy00ihZ3FcatdGwMU1mFuwl+Wnx6AQxAjekYGlJl2Rbg/hL/OrtsCp
l6QXuvFXbSKCamXBGuNTX12j8BYzZeh3C8p8/SD21IPsjMuIfSoXH/RJLsUfTibciwEv6GjMyCpU
E3O77X4/iVzQKibhGSSbqdKDyuINfJJ8bVGFVqwKhFUJe95mHhW5PDBKKABhmXQOjhXCjjnNySQ8
wBEVGwRaMXmYVij9/MjkZf8/quExdeZfgcGERIeGeOCy/w8mM9YElcz4oln3ng3T6c3XrmXtLsIq
iTB+INXklwHbPKZ000XCesjoerer5xk3PYmAtCgICoTWB5oNJM3TXuDE+Bc/FTSkVUw8ytDD1j/Y
1UZuGWJmVtDNDVHX3G9I2JViYQBNq1zWhSoPBvKvjSrbPpUH0B84px+Kn9xa3/WwzB24KPA0YtIf
OwS+jk3COoWDfhRZKDcjlKlte8PJ+vXzLwQcrjp/yzOL5wYv3aVGGJT5tu5XD0zeAMD4jK2BdeXe
J2HgBOM78n6+UiYStW7m5WG3CA5MHfoPjeuHXUXI3oIwwyEqaH8ZYZc3pPwiWv0UXzJJIPvdtZIW
H5iB0cZo8MGD86VJR1SL9uMnI9IoBoKveNEfeGK9yEqteYAph+L0rddbhpR+byZwSZ9WvwXAR98C
A3/ORQY2JZQ2SNlIkbXGLciXgqisE0y7E3e1frGtoZAXob2+3UvELrTQt4d+UbR8M+2LJmgpOdnY
ZtOjV0qHqFszgfetXTMDSXTMIJtMWUBKuV2CZngSVQB0z2sXHNQ59Sxu4M2F3HzaC8ME2nHq7Dj0
HgP9OjGed+DeKsaxeHFGBcIzSCFh3gwiNV4GMlqsNsPp4kKBNPPdUHb8gQifnHohaRLFuHXQ/pTk
s5mK4mpFHqoVuj5waVHkUooTRSj7gttJgpsaxBjwkTaPhx1yUAvN1kTFkV48XEuv5Td656b3t87E
PGC0s+uVxoeK5O91QQ5C4lzfbZIetugLD/YTABP7OMqLrZ8T/bFolY4BMahqLy4NDqJT6uzmrXCv
m3e+4edRLIgMsdNiqUZNBsHXf8UuELZeT61kuBuWZmzufRiAcysYg7lPpEcRSlKhG7+mzy1gmbZV
GC/QYPfx5mexuqPKOoVDduyBQS3IV32cYmnzJ3wcigtAR27oQHHbnWNtB1/FRZ4lNMyaz6yNJa7I
TCajNC05QTO5DqyB67+RbwWPl1bVinqwZd3ZQX8s7ZxyPYejVQFEmw858H6q8porSLJldGxhN6zF
YBZcCDJ6Uh/M1UTT6p9Lgnn3MKpUW2rERVMRWvmSwWDdnvdPM3l0J+Z6v68I3+5f14UOxK4WcLY1
WTmIYcUPxPWlxl909CEjFvh+FLWchNihOwwG+G8gz+JcgjJOADxOenJ0ebybud4A02GyamwZdDd9
qVP8AIMaPEjkxQVnTmZz1tRy+/y6QSGXwwfpKsX2BukhN4Rj9rC/DHkwwj63QBDBJuaxqwn1EUSU
bRR+ylwxGDJL9IvMt13yj0Rpdz18t/xbss2/BfFpILAGq87+Sj+i9qKhJ3Rn2A29k2w4Obj+nFCY
hgIsVHz/yIVlh4MSuuZp2cY3MRXqxGVTgGREzhRMGw6q7qrR2Dxt0LtuZHDCTg3rV/6pH+j6I2+e
iz+4oSZj5kzfk/btBUHZZs5HlZ+lj01Vdr54jvoOxloNreEm6V6RSbcoj7uQUAJJ/V3PZ/xKGwK4
TQNW/Mv3j4o+BeTUReMyLm2vNtd7T17kqqtXTI6Qdklg1HhdA+mFbVLa3/K6R6vYPuH5LRfa2pkF
iWtuhP1SkDKr+NP3rpbpAlud1duWLBVw4HsKr6GtJe1jKo20IDhokbBUsjerbJ8XfNjcXeYZWYaX
5oZZyY6vDTtElL5BP3dx+75sjlIMpUPY+JcxP9EpHlRF21zr1tUhQjKfDx6QQMMVlMD/IkWFxK40
te0Akx3hvnUQXpu/6RePCUOVDttTniHsaB6ioCEFcMGUoBFRattm9Ro0TbxHBu2Nda7BfzWec0/z
1MQAqFrwTfr7pYyDD74iIUeItRqHmXFsbWXlPUumIz7MAxVuBc3F+QFol3vqHR++D6he96VcyLaG
yJ9kANWXx174OT0ll1ohzIC3qsSq6a/q1Roh/Xkz7CdIWjD+ETsmyHjXJRRKbotS+y7ptvZLOIX9
HNxYkvDRPnw4mcGg4gfRYixewAFXQZQ3bxnxHpI7O8p3VgR+rFmIckwgYvr2X3c67siAXKzHUrW7
5KP9xQKUwO/KUcFTyrRY/aLj7GHFgnDvWSTrtRvi1POgQ4/jrXKTx7RUa8mZgOw5BDgXdR0tfrN9
+6WHE+emMCrM+dyBUqP2/DorW8lL+q35z/kj7NLMLKghh+f+Xn/5g+awzzIu0pkLLjbDV6zntxE6
MTp7/v8sSSROWR8w1wh80V/u9GK6M7ZQTVAceP/6Nsef4mv+pX1TAJPAUSwkPA80mHdd/8k5+j9J
/noQLqMOyrkw2Vvb5ZL9m5JoAUT4/vxUR2TV/ZkA5vm4QKeWM2wdXxS5wZC6vvflkScgCgjd0l+1
GcTesBQdN1qU1btdeJzQhyHqVLhHSGjn5iZMS/oOKGSJHdp+uewVPWJV3wlLulJ0QANauJdVwBZk
ryUig6CNrvZMTgu+G5NKQYueSUaWEvLIS+GIWshTSOqS48H09p93X7ud0v1afGwV+vaxx7njMaEz
VtjJi5Ronco69NAy4FkKLu8RuS34I+Q4BevpY2puKgpZqPUKzAo3+XzRuoHfWODFfMjhexx1mYPG
rXywal8EFA60rGlDZYJhQ+HSJ4fZEe5HiUd0wxBJp0euLOxHsL9GUgk2PXOGJfFI+gD1+UCFgv+d
NWD2Oe18JDgmdyseCp+WrVXWBv/UQzcpXp0XbR5HrAadnsiWNjjZFxKzaXR7OG4p6JS2+ksKzWLC
NS/CzuIcFlcT0Q4RHC01ADzd8tynWxgryZet+sq8h8fuU2R83mnO0kmBcJ4boX+aIDQnV6nxtndY
dRWRtLVhVUfMKcOmt7qC7CiHdxZbqRiOKjjB10o7z2xe9zQ1KSz3hYUNnv4b0y1xEqP97YyXpnQw
KeEG4UMlhBLEEHMW4fvzv3vPrtVq0G5mLo1lcduA2xqUyGEWSC6soug/T3IrBslx9Da7tclu2p/f
k2a0fgwx+WTovrsUq6rgQgToVknZrnw/89rozaSjPf5dBxWJu6bua9bwUr5TL7aFH+ziWcQg/jMv
j0NYn8CPeZ4d8Xz10s5qxHxkP+YsgoydlJuz6bkyzL8j/9QF6slOsZtAW38gDDeIc4lmYaSSnxj9
HfnzkgtkXGDCLe3JFFsJnxIawX/KOcEJ8wtYCWdFemE+iiSdvfqD7ErIg9Y8IPWRNH5qkhIPk6rv
qzIUkaEi7YzHslpdpjma0ExSPtxiJh3IRfWTrotnmfnBWjPNAisxx5Hw35jUUr0fhT16D6AMCURx
DTNWgdN2dTP8HXSZTRkVLZYNJkA+uOzetajA9KFYb/iYQmAX0O2yhS8lW1E95Yf93Ele1l2Ga8FQ
6v3FlkNPFSpYb0Xcn6wpsfCK5mcyu1JUz4qV/RwzP/psFXgggtbFfwbrAaTK6roFMfS72mgjPrUX
ynbgH3K1xM3o9BXEWKLCTmWbeFmAO9DLXHKGdjLnNt95DW0UTS6eUySOv7R1g7eDh/aEAK4NFRr3
Bo3R89KxLU9ut5NOqSaFTWy2BAPtfpRjfyldxmyqI0cZQ3oseHsysznQAjDAUJDMCdsYXCDSDBhA
SaTcUv3FhRKz4UB6aRudLAK5eMm5kuIJpPGw/WEwygk0jhQKYS0b5ewL7+kC4bfeO0tUs6qdcs+8
f1MBS5zyo+MAlL8gNZcr7ocCDsWWXaVl1KWnpbcTPSozew4/mD4IJhamHLuGdSoqNEkGbZgg2DtD
Hi/woPlQtbiNZ3rpSHemHU9NIxK+OAWKrAPHL86rAsn0eM8fk702zFzUDFNhfVkkWG2QoDsGfPYI
ztYtLaIIDEO3AS7l+VTKmIc0LT9G6fzjHMArJ1sarVAXTxU9AJ1xOkOAdPPk0KwJSJi9g47KCwsY
bn1x0A+m/EammoAmeEHX5Iso72Kzlr2vxfu6BXouvd7W+AzYOesMIgHObpC2OyWJHkcTBjCv0BX/
UeCtqlEE3UNLYTFT+XEOjkyE800QcHBDb3BApWY5ST3MqOHRx+ol5vmE6/avSGDWngRiJgpeYlwm
dsgjsKXwl+aJm7yM7cQPTzh1zN2/705jk2Rv7twu3G5cgdLOF03TatSAFaKKJZp+Rlz0H/yVRZKi
QPn3nhqS9gItPPUyRrauqlXbe6rRNloufeVtmY1M/Dw1Nl8W8malHIenwM8V+R5RSic29hCVxd0M
iKCaOviQJhVtSUDPq/GyXymzhNkhxIvvrORrpRKIBtLv7NXB1p6N1lb8UiqORaguDCl1UeyLSkVA
ac2LBbLw8PKr6Do/K4E1EkgR9pjt+/93sp24BD9wn3cpB0kbsZjt+0ay3l0RfLbaGbbpS5ure599
7yX4ZH5LtqJrnPBLm+cGa13gOMnPOYfXT1VNfyOMyCIB/IIXaIuTnQwoiWThiKyo6FomnyzarJjb
iAeNOIPcxe7EeljarZEHaItuBi6h5LonjORPRO27/4+Lm3/vkf3z7NLYWt/2WeuYREDjAmoa0Agc
TGIbjX+nEPzoHTIaQ8cV+IUveYHlckL8blf/fr46nhIhei8ZT/aduDkvDGIOzqyOvKRPrzzrcHCW
Y7GmE0UBkRCBIv7qV587VO67hO1ChxiWBjdX7a6pKWLhQ7jqfkyoMHJIDCqOutRAaIUHyOuOrg6K
rA4JznROAC70GlqLwkIIUhniGTPfgrDISczVYa5bX8xBxPgwYusgsof7fg3JsTkn/6pL/PgAA8Ed
moWa9EvWU3MJvQCAINCJbXtBQUv7+hc98utmXhNP0kfnqXmJT4mM9uhOVQ51Q3tiqKHFGGQshbZb
LjkL6reWq4Cv8yfJix/3Y3Q/qU68CoeUVDW+Z0uAcageoSIJc0ypph4g4c7yZxes7G9ggsug0mUh
G0lNnEjwv+TJo+lHiLvmZGYTxFsXb8nuOvGe28LR1h7nJHgVaydsIUJBBF6jFTT1Yd6XqCCIUniV
2NMTvpKCrE1oJKbsPQthaBWvhiL2rwk4lvznBM03lEsPQoewsAQwpFerEjUyfF1sKPL5V4/caFSB
PAJktDh5LBW8Fh5CALcOxQtpqIfWs8D9wrd7aMB28iXtDkUXr8bs91MP+6gk1nJggg/GyF3JUNJ2
E/H5XDleTJ7ScSq7mij/VqO0rqqLWtYRTOzDcS8rnS1EFo0x493X/FVl48bOc9MueaeemqsDYTKn
37QxNt/eqL83BwhFG4bJt3A2c8jvga+dU0HxKdlhsorn9ApOYNhiQes5gDxCI1/YLNr2po5O6rD5
PA965dTrOj+4H3sCFidtVJhxCEdxwNYJqPgzdco4+zqyba4wo4OSUFyTeNtyD/HF9KRpwCympumZ
MX2bTX6+Utqjlekxk55p9zRdGe7j3afqGgNNkjb2nuHQo15skGRHYu07YXV0LWvCr5t+MxzIF8Vt
SgnfrS4q3WWLKMiXVLejNJECjErOQNu2jaiZ06DaVhJkoT2lDpJe0DBptkOOoJ1/4YH7rjC4WumA
hlNF3Vsb7Y1v8VH1A5FYAeVvCh2t/lnOGJ9MFeSlRwVNohVnaJ0jYKFGls6blyKtPON1ovRnF4Lr
Ywc12mHa/G9rAa2tGVwlxNTlar8IUrrvGoNJWSy/RNebUlUfpU/n3Gioci4KDGZBTtBz1Ofal1Ak
gwsGsgQmWWeYy7z9T9mUN/8h+J+NvIqI3/gdGPGVgRBZcrX4khR0uNm6Zi8gVgymaXYIkVNv2PRt
yDAhSDkPR6jJVgghBiTVqdSK7HrZRuYpqxpvVR07Uh1qxPl8dW87/w0xm+S/1O4m+iFwOvZsPBOZ
rwoYlrgl3/0Mz1G+8dO+F+n+6NtPfBj35qI6OXXC6SxnDn8JOK8F1HMP3OrHXXScqs2yKDQSvoS6
5x6WQ0KqkkGdvCKbaeedRG4XfhEMrKH7yOUU+rhSC9SpH6x9eXfRva9lmnOw35lrGlOHBr+rXmEf
qgXCLQlNU7FPmt3n2xJ2FaeL4VGNYHi8cIHwHbqvLWPZ2zDtb0L/k/cCsm86kMOhHVlnt59vN+6S
4J01XbUWM4u40tuLtggK+EK1plrBG66UQzw0t7mD10x8MT4tEXhOYpgQ9Lx28Jxh1LOt2OM1I+AP
GtZO4t5q2tuDf3x+S21WYIjKF+kJOaaYoWHcXqYgAwqwMR7SKX7So1PSVJiYw/dAjHEVzdJcEBwW
8ITxfEQ58fg90da5NQXvP7QumcxSuG6cEOnw6R3jTJmdkF4c0ZLMQ3gTsks5+JivQAitUu0BDgfC
U8BPiPs5BeIMBDHNNF06R1j+t137w6n+wc71vHpgqe2nCSIvDTpby/egGoN3wrvy2LMs8nhdWRs9
RuxgAxI7KIoSdW3JRss06kT6LScovYHY9544QuBD7YXCcPOQ2Oy3n/dN9Xa4Mt8NJF5Ocdh6qeSK
4Df/yHX0JdADcSKV3exckjsYYCUSExzWkzdLuLL+cEQxdQK8ScfNI/5v9JFlqheFSJ5B7Gvc3hyy
IFMa5GV1vWyONyWRizHThHbVkwIhTQ/dCWJygmiGZqgE91EzuDmbHq7Om9OaVAfSWq5C1q8bI9ow
8d4OtWovc6SPMMILqAJ1ec7oIHHofDsi33+EWpegd9s/zkYsOP6ucsvNwpSKgVCOOBl31R2YNISX
5RIJ9mZHgFfzIevgNsz8GXgmJt9f4j/HhkcQuHwyI3e/UK5PAhExiJW9ErNzFOu7j01Vw7GSVTUn
T3vCtGEpBJuZwLZnDVUSfBwk+u6GbNQYmDbB64AkWg7CvLtaS67LOy0R3rsCkeG1A6vJwCF1tqbx
83G9NxHj4Iyt4rxd61FZ4h31a51m0pD7S7D4enGCI532RUJ5MULUrvfmiLtBlGhDPX5Z4e85tMC7
vq3HrH6I38x0i8MbQEthe9eKnvm3x8WK8xP6NSIQh/kLlzsRFbQ6fxpFH2Ar2L/dDLHvZoep+cab
5AwWPEVJZDqSZRA71bNM5EsAKVob8UsS/jsKvbJ8+n4KKP/1a69nryIDbzOHQ6/ckdhuNX1ydvW9
KGAbUE7QUVzNKS2R7lBYwWvQQdzNF8Xy0nQ2+b6OrBIuqN27Zb78Z83cuaXjZUZMHYWyS6m2YOgo
S6keQffXkCPToJEo/hy4tXwXIsKfoiOqmcqPpPHFh4noFElbuPjBylcLKVYZn+GUCtlo20VlTDqd
26dhtcd9Fz4dgk7SQzsOP9osmVE3NZr/CAYLj+OF+t0m6GPgIWatvijgKLm/tbEAMHAhoB3VRuwU
KsotA7HoUyPoXI+Az4j3LjYlZv8JIyJukTWEn3BSc/yIsibPjqPdzAcV3G+wO8jEAuSugnwt0zqX
OTAwC70oUQdFFWiWJz4uPP3kwqMt0u9/JGTPvjS1kTlzjCWZ88jkiLbN5UDgf58on+SSA7wlNDWd
AuNB4kyRr8bRolgxkowCKV5y1z5qn5v1tawLlMsEk7GrcoqWarKrmgRIN+rqlMxMNLSp96W9VHYZ
6Kfex/703o2wvFB2Ld3c9r/TuSAp6LRNLz7n1yuxt8xdLT07xAI/OPwivdutjEjjE3tG1KrAJJ7j
vG/vocz35dGnXLD+lcih/ZxF+vJDbDD9KqPPWtUDliN6EhaGyZX9yETUGNYiyzAzY93qp0KGYT/L
lyRsfEiHGw5X+G2Z3S5JioFv5rx9zhAIly6ey4o6LqbLFbo3GPONP3F6v/7c87eePjVaor/RPxTD
QlKhZeKdE1UTB0ZI/MbPYztvGsnBS/QM7Lnm3zw8oWVkHEbgJjhivW9l9e+Kwsi5SSGoYmjwsOPs
mWMJkmJCREYtTGjZBeb4Sm9B6xzlSoVpgzHj3MO6PaxQPjo3YYvSeT3himKR0zQGMkGityK5V3qk
Ezg7sZ8ZdaHw66rOpHbwJein886ld8o4Jug12ALETAHbcUVWN79EOstoqjEPpsr5BLgR5FGIa1H0
Av6F4DHyjtw0Uum5NnDcteLIbT3wHbYC7Ry7jDWqCmVBDRyk13vqxCztdO7FcAfKE7LPTatPKfnp
uYHjkCl5pyUcHm/XYsxXtt/cel5UMHVMJbvpKa6pIuo+33VZBYobiVm30p4r/pOxHIBi5VdnY1KM
UpDud7f8VzkCgZRRnmiTUN02q9y+/orrWaimaFXVWTp85NlHQEkkmTEcBHL5hqVwuC+xpjJ6YEE3
4urjczG25/lzWnJW2PNQYY2taeyYW0jc4zMi3OTKJpU2EPLHfdpUjwyNtNMdIoe3PGL+7PmZWA1O
DOu95tExU+jXyA3dGmWsrHqueNqAQgN3BXdpGeLGCfQFrRNHySA2JXonlFgkmtrhsLwzoiX2hEkx
7bNC8xICdvP8mWGr0egpfqMQKAbKiTCXFT5dnaZpvWCkSkjc7FbIEcQSi4+9LUlcROcDUu9ioxR9
AQthhdnXLDSooia+WBgjfutZQ+X67LI8owsE7IeEFZ+GvJjiL59J3n2YrEou5B+dUL4P3rfwokmF
68UlS/f127jLlMCT2jrPcONPNhDLd3gLG795TxhJtYRC7bUel/luYB+vorWzo8Wfy04BEVr+F3q6
8rI122aU4SOcXjHSXK6fwiE5g5Svq3wAoT8bQn30okBxAfQX2Jbbo0o5KYPmgbfDoGrC3JyMCMQI
7RkrPy0xhj+jn3eadvrWhOTcjn3T12DZy2Ox1JpozFw5j7zscS+jQBJsRSKjE3wYNxKJ2blnymC2
DzvW9agRXstxdfmCrA/PlXy89pS8M0joHxLjVcUg0TPeJlAfZwIxBU7IoXKaqGZZjfQ5WrgAorsI
kApcQdrCLcyyEaTAECFaQHWkxHCQedzgh5bHsfxSZVFlnbt1ADqDI73Emns+7JwCQuLRpbhamxL5
YtbVpfnbL97xglRgsdsmFZSVzxRh9P3c5FS/svx/VI0CJVRAy3GSjg2LH9Pcd3sfdtKxs6QnfCdz
yumkAGfD13kuxwcylO3Cu6gXV4Sb34h+IQebIl5VY6GxhBl3UjunZqfFymk6DXbI3/Wqd/HGGWCq
du3JRlvj7KVhmeKsCXLyrnvCFkzgGU895NBUfhhBhlbbQglwrMipkVfDTladnf4eoGq0pQjPcf2Q
CGp7KvGKpmYR05+9zcTDPj3WS1zb+f5IEaTFU3+8FWFQDVniaDKhSNvru7WLOYDqnt7vxPXEBg93
3Gq0XQ2EJ2X5+lK9PGc/QEVcTvEH43dm1oGHXg3YvMSoUfIaYp9KKPFuc93Lsqn+JFsGO5JXEcGC
9ZMjhbfElIo8O29uOeNBh4L4+c7c6uKQIfP9wk82NmuwmdgnRTctY1ZeasPFbx0h3y1ErhJKeYBj
Ly56f7kiQtw6FZD3kcRwOnd9hI3Dfq01YRnCNv2Q0JwX95EU6yta1TNQx3/pgl9rKXOT4ZFPu7p2
Z1P8U1sBdgzq8j2idgWS7EgRlmrUnTFeYu7dT1eWMGrHq4dR8FH+4Xq8fpWWyEHMyw1LXIaJpgjL
nQ6vsHpTa5M4OzD+nFUl83UfhZWM0feV9GXXHlWEC30+xLiLciVhoKmf0AVyuamIAwGRlsczIeHB
3fXF/CeG2APNRaWtaRnWJE67awFbtWt85K5yaZz6Phl0mZkThk34DPBO6SUm+a2AQ87gAgkILsei
xCWFlJ/8EtSDf/vuV8Z3LW26iWSDvi7BcLPRxSP3DTlLfCC23ev5ZlJNxBEotl3rKjku/Zx5FPAW
1KYn5GXAciEZusXjnurGBF/bEmobKaP/CVQcrjdbAkBJjB0xme6Sr11EGzvnXlzicnP74S/WAzKH
dv1PdSGxjFS5Apy9TdWXhfb4YwP/yYjWc4xFvX+eu7Y2zbbkrCgKKxQy1SJQ2KJ0+I5UID9ZT6Dz
akRyMyJnPW17fUrFfO4liXmZweMA6iMGXg5eMYENNGReBwKaXpdZvV7VDAnUyx93MEEoiwwE4/xI
/SPB9V5SjSadRrSRLYvBoDNiBeRTKdX9FrUochK5J1P4v9ZMPx+ejxEBC/okOmzRsGQ+IBQ/R3iI
UOJkw4aGqOVNMxpHg/43yMjsOr0sDTBeC1B/0zHS8dlTVb2y32x627r0P8k4BgfydC2QIiKQUo5h
el5kOwf61FaDIxYEiW/madPhAFFaa+OpvHxBh2ABJX7P9pmuoWfyCYFAjobFEo2PRPvNgNLzSx9u
IPbhlhO7irKzJJCsfsWWtSuKSO7vRjdMGcsgJqMYvD55kd/5RTz7Lhp2YG/gWje0nHwZZ+yjudaU
8S0FNuBY25ml4UsL+AjRdpIK11b0n74L0bqmGXo4sfICBHHdkpA01JOmVCcMBJ+4TUPzsxUuEnjz
NuB3mH8B6fXfmvA4rLlj99stL25ZJjohpEntr/e0rJ392bFnuyKjRC4Fn2CUst5m3PicpQX1S1Tt
bW4d9kZkjESICycS998MouPVVZHvez1Psy+n8pAXxcg6gn0rl0QGj7CzqajnSEZ0h7SNOhWFdnb5
r7TCnPsodEzx8xvTVDETfQ+ux6zYA1McGG49j66uio3KwEnHAx0TbaGphVCOVYY4chk5JwZGEua/
n2UzxpjfhhbUjiPvxHqApVo+r4cy+TFO7XRgiPf6tubbQLdb5tcGSfd61pUMpzzI7Z1Vm3YgOe69
D4YHu8XDJ5JDcOMgMLpbz64H02k4rwp/UXs0JNqGvtfEC5kBefEX0YPfp0cRy7hmgMd0MS0z9mAF
zjWmzCar8zogx4Iy14C5r1f13MzAXVR1/LUFF3dKU5VP4dZKrfbigIQOYzAv660Ppgty6kG0qLmv
ufuWapE43HlGTZaV6wi/+iNJgLmlfW/nYKTrC24dRb8OFp/wt678mazCKMZI99ovHUXM/uNR8Bzv
Wt9nF5949/vM0qDdh6/sUCRKFB56Oozt6PDwaPod1QfOLPSc4JStDSQ7fl1P2Z7DcYnxFjoJzjl1
ki+yzfgrZACgGtRlVEnDa2gxshx+PtWQ2j/X2CZehWFt0bdQziFo9lY195viGrG63wL41lgQSZEo
tYYREiDJK4qSEhvx4tcZ/OvTF7phQVPIoDdNodpE6UT5H6mU9TM05vafMPzo60YHwZHIa35qYBFF
a0D7zl3g5kX2o63f7jz8eDKoYLCV9ptUhCQ7u95MBtgsqlxRzFzLy2csI5koTHtT88753ZlutlO8
LVVN/ApHmzAPntDF6VSyDBi1ZZRKuUvl8o31gt4bLKkbCHPiXayJ3qBHKQ/RUcvSO3XJWtcrKD+t
hBSYN22PTYxgcR2pOejDS/5O0qQU9QxrmdNCJbwL7XVAHVGVYyOYK/y4y7Fbeclmhwz5WFP36LrR
e0wV6NohvYBe1zh88Uw5+h8SNq7coHE57FlA3fKqxbMfU9FoEBGZvh3+803NE0dN78EQOm/V8gxI
HQrRVeXHnQrrTUk7Fy6DGCA59tc2MzaqxYTJPX4amXSPm34k+Nmm2viseYbNlaSo7rf33XT40mOy
Sx/vIhCuLNk/e9/QI6FQsnNPEw9bgCSUiqWVsdS+25z/iRa5ciZ+nMCoGIMH+aLca4QX3t6Ov35F
e8+DXe1gX/QRt9qL/bSWtmPxYYIVhXTyWHtPX1dKh303STiOIX4O+WdNEUh998gruwa6qujT4jid
/D6y0mtBevFj79uT6sLQmeuT674FjRT49R7BE/0kXDEPY0sHEEOScg3dsnnwkPYhn+PtqaDeOnFl
0CBsZG8OLzQ0qOByeTCjii/MO3eEVnK3U6j3NaBfNTI+/ehGvok6chNb2rb2RSTbs98c19Y2yfi8
7r/1lI837Zfbb3+ofH7klxtnPjBniJ2Vyh16bMEbquHY/aknYlyoEQhpp2LxjkYAfwAaX5Wcyv4i
gaOCzkzcSFRR/HK4Ohnr7tMcKkGpa9j2Av9S78URcmZfWGOcRBDVR8v+FENvTCSiiJ5Se5yIsqZ5
5OLuHGp/8xFwL3ywelNb2h416NmVfuNK5V8uvjKJR2QirG9OZ1mAc3Vn1pA8vApSgMjmBdf5sAj7
KdORStf/Krso2qBQjM5ySq9suV+TwGaL4sEhtUu3POh4OBbn+t2GWbEGx2KStH/AMJWclN9qC3XE
wrz3w/8iC+4ctE8fXCuw9lJGAjUpJ3C6YplOVmhzYwp6P3e5dhdOj4HBXVfpR2JHPI8Cl+Lu+8pU
DaUyiBJ5vqv7RRbJ3MvzmDfPK8imbfXll3YB+mtZhWaNWFjopl66nr6i/BPzby9gWU+aTg6877pe
TlzabW/9udgWRsB8Zzs1G8/BDi8f6oDDILxVautGaW70IGeuaUykoxmMiDgMtdssxYJcdohDoV+R
fut9fzpQQPjyDNm0hpwF0W/wUcKABKJ2PwhB/t5yMIlv882ofZ02WGtPlxl0NBhxBxeXp7A8RADu
ySjfHfI89qf0qB91PCOtd8OOHNiUf9Y4uZingdvJA05i54e+7xUvOXySJn+I4KL4UMqVlpYpGgmC
VuSoJuiPtKwAtsK7Wx2SvqpGUIaXNmYvNpbJ0ZK3es2oxsZwPDgIzGwHqpKIPf5r7nAct95wmUAZ
8Seqh9nMwdyACJvNHJWkHHVFWJqRZSyTEE3XHPhXeDrfWycB+zBqPiJbmNKR99nseYQiJdvetL/h
ylRz5gEjyJkJ0Ubldh6AulvOk8NrtwcmSnIg1ObHL78vWqdm9XmMt9iGhYX8ZoXjeb+25aSOP+pP
IktBlsWwCtk0lei7YAsDyuC4bhC6qEyd1LfFh1IJqwbi4kbrST0EQbxGsZD+hlWnyVSCmNRidofJ
0Dtmb2sj0uTjuS4mA6a4BU6JQxKhkLH7greX8TtXGBAPfR/q5vUXWaNZvhuvN8qJzc3erPwLlhPz
2ig8rFgWYxhfFEB9RUgiPG4Efsb0R949aXWYU/kJXfjWwn5XFtypa6wmWKVTnCz3ToMG3p6qUKaa
yw/gEwAugFYQh4edRpVyOa3CEuSx8zuEAm1FzrDOIsJii9yre0ULBNTTLCfbvoAiN9l+3JO9ieuG
9Oe9nX1lEy4KYfCBrLTcTWfIZhzPsiaBkUr7Dq2Hv7CilWcwhTIUztcCbklfVjuPg3P/fqU0aDdz
gOrCu0VjH4Z3Agv3Twsdu0Yo7UNHdPMun0aH5fpi+Osl1So+e2HU5TnlMMCMPtVwIzfqnBA+XoRs
FZkW3UryF0OvpZ6jio3hzUw4owTF+BYv5jCZN0T3Sj4JhNvzmCjZpNda7QNhDlP7ZaOGTM5Daj2g
ilVPKbkQ9xQ1G5oqhkVkP0Y3PXP6ffkzDenr3sCnP3qyUCdmXYIGHu70NLXSISj0XIQxwlUk6W+D
CURWEjhfgmvbJ4bNmzd/KpTdyJ4j/EYrkBQScx9darg6zFf47Ufo47Vh78mSY/0aXnaoIi4HzmhF
Kfa5nqvSOLw4Xol5QJVsa2eygF8rSwMXzoD+P/ng+G1ALVMlGUz/9Y8tFAte0NxCAgbAxpn+9Kl+
pCX/r89I7j4AxxN8g7iXrm8Q3ZaWkHjkV9uKfSWz+e5quaKalBbXXs1UGJZKh/v7bKz/oF7tlOjT
ZDi6zc4guFlV7TxLtgk74TiaoCSQNevxhTjzX+wUO+7pe6vhKDOqrTUcoPBHgtBnI8zH/MBtaCob
nkKtmMOPjm+h/vtJnbNDC+iYD5AodvQxzaKGtY24m/B9O2x+UeGUsqVy1gS+RJfFtF2J2rePqdqf
2ycgRe0Tn34WMKet+9iq27bi7P16cqmT6k/3i52r/KskiyVMKcnQLoRRTBPBdO+6WTA61oAny/VL
KJerPExuNhadn+zQeP5r2ppUUDXmkOvOhfU2Dp+vUjP0DuX+qDjOwD0/aktuJtOIcUm1awy9rV2o
a1qYv6KwAgAW3h0uKO02th3aoC9hkcOtz6dXTF1/C2DGzEvP0F03yYm3S1sZRB60ogqGHQqdnr47
BLDjaWeVJheWrlFKpoNpteHausHD5GRri78YUJfim/zILhjysoF2gNiEOlSOM66lBFpd9biVb0Zp
b5k95yi+XpRYyc6Bb/XOuNUDl3wq/8TMVr/mZSROcW0LzEObcNcy0GRJ3Dzl28lplToxahQqYacZ
+bla72yPMQdvAMTW3onf/Al4vRU0+ZgBZXi4dYLTC8ZLTz56PP2myuiFuADjiTOqZmQ36hbQXVCl
k2ElNklIZUQjesq9jlQ684EW6dirFtW87xht9OsJWJDVA0uF8HTI+yBzyZmxeVkfBk1nOuBbsmwk
sivn4B2ph7dQa2qPCq9yu7Ykth13uZp64n1ZuM3hf0P8W/zlIdhQnrigSBgnZ+fztS+Hiy/oSRVV
Wn9HjturkdNqnuyYAwIgsLE1VPXk2Xt/Rx6sIB2HnjLy3Rx76rRY2M+1bnmUQMl2OXI+Y0XD3elj
Jr31xLAmoDmHwj7zfKrt1u6QWTNPZpgaNiZI6W6+VSPzfeztN3IkZ44dCO3ZOp1byMoItE70NQTz
5AgI4pgUdwsf4EyQeSKNX5Mo3GOwf2QQNVXuvIp2Ul+1cho/Atw5P5UOABK3yoqn9/cFWmmPPWJ4
wyYdqkrA151gJVPtDXhBPVjwOxjU9phO5dD2ECeLhZ/eoF8bbpMwX5yq6y26yezd46ZDphn+VBSb
01wpe6rk9KStwuEljspsTbpjeHvA/DccQOy4WXIvIbrUIlFqhrtbs67iRHXxBjAtVljAk7X09lCF
qfOo7cujs1K2cH2LKoJdCWBj7OKB18gZ/Peir5WHS+OXvI8HuD/N8uUN87LbkaH4nrshPw92qpOo
rwLfjcOHJKw4X3rbGXZkvhgdIzLOMcdINN6jqLNcNLsmk1KoR7YP7U8x5t8B6JHZHMPOhr12jdku
npgnyqoEar+/4TuSfyqaCdBRcBKh1HGgByoHW35cGo2SB6nHBg5YPcSpzoQaDDK7s0Hjt6a2PwkO
xN4fxT2ND786e9q1gTBDvgAnme8EM4Bko3L1IOVBZhJKWyyKxQfWbimLdLiIbvNdSTUZ1kYheJz8
pL9px1gNKtJR8ySrVrQmBEQoml0hI99GIJe84d6+E8VmtTGQ5K1M5Jm1ugqa64zOvFN7QcpAT81f
ud13t/sbRATpvUTZKiThgJ5jdh8GAvWDHIjArCR7ORrAOJKuLhSXs2RqGt/pEAcbex7dtLKFw0WD
8iwAQseNXgDV/JP+peeMBuTjeh2WPhq7SmR8eB1I3yEMr5YrfIxbDRMD1dKi4gnNosMlllY+aqs9
TuBlwUhs0zSZ6nf0ZPEIpmQAExAIqvB/pwcytPzkgMdgbpJNi/WVKfYLb+hD77tHDnkjJmqV4QeU
5n/M5o5TjA14rUwSYluuqVQIWqJLizPWJUPO8zMmuko1gnSMVZtlxqyaN94xOLvGL5iv6UzIhCu9
49AtBt37NIcWtgkZkuoEzz/DG0G8Zs3goOyXwpu1hZq5w81I1sQmayZpfI8KOGCE11C8s2xE5Oa+
erS010Q4i26mSHJB/49db9l7J+9Nu5mha+aHbFHVDqjAKdFRPbskgiynCGeqE+LkjOuf2heL3SV+
L16jA9UUw5/ZC4HRGbVloK0BGzmDJK6393lcw3NgpjH7JZcj1rA3UFgJ5mbD+CyvP5SgKTv9wQAj
BfJQ9kDtvZWV3SNZWNkFZO4qLD5p+LyWu6gYbP7By06NxE6a/aaDr3krHspbn7Dn2Z0MlRAaok08
nHc0ytLb5UJTxwwIUws57XnHS28SB3YPFzz9CHBvX4BT/vS8IMq/FaI42U/NONJhqrV18EoZYVJv
Y0O8EvxMmyP4XTcOVPa9GUY5MpTu51XAXtkhHaps0CExQ/1LfbWh8Ped3PQmj3v8HGFBqtbzJE8G
tEZiRf5n/L/nKz0Ri+ZHJ2L/HteGucZ+mjfDcCzXZ9AcZ2PDuYj7ImQIS3YbogN6xlfM3LGA3jan
AyB6YTP1y7C+VFR42Zt+4RFFdvRTSSLrZuwNiWAQiyJxBgUOwit3Ro1ozNJJ1vnRqpkRADoVR17l
NYSIWacv/cJ22GuJ/5l2UM/NbzzseUxF994bBAog9KUKV+8ItwbQzX7CDiAX48rEZbBZ/LAM9kEA
z5Te7wExxMwk+WKbbCfhJAOxG3dYDrabyYL3T4xt2CZKQAo6jeXIoard2mVqDwBdhL4eLHCnqxnB
Q6VhCG75brnz9rlUXHxYadAV2UYFeDZfeggH5fbEcsDisfRT8cUH68g6OyOssCTjmZP9WQd+H/YI
VVNJH/8SelVNYKXoRiENF83L4fkvlqPjovlVLX701HIYR0HblqEo73mu3mb2Ov9jpxt++ZiB7LRa
m2MVYe3mXpLE4k68RLQfktux5uADN0F3wSdmmoQaXWSMp4NSy2xS1uHOHYvFrr+99Li1jIci/C4E
00hr+KCUNBa3O+FefrzQKTj/Dc0rGsEt1MQ4fuOWcR/Zeew9xgZ7WizO3sSl2aFFeApWcoFoztS0
2m9KANAC9Z34e5rNn1Mn3VlW/CvcMoAt81FNH/g1zoTvgEYzW+b5dBR4NOrerk/hzmSmj0Z3kMeM
HZF08nKNUrKZiuhUIuJMR17m7UGHeoJrtQYmEh5TGeNIbxmRbge8me9pUMqoeNogzy1NwSoVcSHQ
QmuA4g6YXgI2QlzQtReCaZhilzEZJ5BjJQ2FNTPrp/cnfZDh1N4TFsXjtgjXqgOOu7glkNgeojsw
/VoIwmHDV4KG3YZyrP+dPRSY84eoBtrjC1gGU2alw6c7xV+JerfCWLf/FSGDa4QOaGjirVKez+e6
qy86yjsi2NgGbUwzk9Oad6nAB2i8uyOYFNhZwl0UM4Emw0Ehwv3Q623US1ARj6mrTwErq0smX9EV
Niak3UmbBugQz5SbjXLRziW1WzDnM0Aug3Bcc/Ey5c8me6WdMvnYI1TJDoWsYigR7T8CEHT4fvRl
2VcqS8S3WvoYVzrEnNuGSpKV7GRlAOm+PXZmudkF8fTzUGK9PrAiPMQfWwCfJVQW0pFySDYNiTFj
/SJef1fZa6f1BrWER7Q9tDFDVNhfRHrQqtvyBZCYFwPZvyFwgwYynzEh6Tk2/vRWlbwZ4erNBwzu
O/HboXBr5NARGUji4Hef5nMHwLiU4FNnoCKkx6EadZTWGOj5mYvfQwYIC6YhI5uBKyp44B6H+bOC
gj3trqCv0J3qlrO8HZzrzm2iBx1IFt6NKtIX2mfzwg9NUF5cjNdxPaSq1JTMzpJ7QjyZIU3saedV
hb36avoCOmmuZ+1DF7ZjBdVa90YRqJSAWhL8c0ZJ2w0C8WJ3RX7hk3/S7VqmKTjjQsbz7S002vaT
nXkSvRsYQqtRPCi/9OoUTDaZeEwEKOkU8eLneGf1aPibozEPYmqfUFCH+wcq8H+gKtQ/jsWWDCwi
Ljv8u2+YN6QQyZQJn4SbWciwjthMhAagiy6qqwdPUafPbQOw9soIQWTrH4FxHYyXTDjDI16VYuvu
bUG3l+mlgEDhTzJsDsq/SbjD8CiuvvFgaG8C8SYwW6cP9CsfG7B59QlLqilee9+M1raY/whkvECc
davFf6iscNAq/81dDLiwsvOyO6owiTppCZNpF7KMbkf3tSDn4MtzHVICko0/jpKcxz/+Zujy92s3
GJDgODHXDG72ky84U/JZk0JZS4dyrgirhboyzj2WiwJMHrYAKC1/B/w0KAwwX9/tpjk7PekV3YGZ
QDos+ROi96d5iedLYTPfVKHP2SWAWjeRx6R+f6FqhukyP7L7aXgmiPTCN744lsgoMWa1NRp0oH41
T1w0mBrVpbF0i+E4L8BR5MU60thaKYhTXN+FdffCSRf7uf9Uyyi/0CcY4de1fMhIfMtXD9ExTdkf
7HSDa8/FXpsgRBKdCg7tm0bRfKok/9NX8gEShoa4fNXnE0SEkFn7KDnJ+WzpfuAv5Ajy20lwcGOD
n0uZsjPSLK7KXDv4U+/8vq+9fWJNJ2i+TJdH8ETP8lKKhEE6YQ+oSfRPN3e7fFuTGZAlDmtHGiaV
gZ4vPqTT+C/C39cpZNT7ycqUWvNBna0TH5kK1y8DHPKAAMDnQ17q+Rd8jXWtvPOhJfp8riRJMP3a
0ujGopoFGaXEwtfZ/ko1EUDyfFwVGTFv1mJaPbZAomNqUW+j4m9VNHfP1X+SJv8+ZdTkrMEmacO9
wNtrcqGRg6UYidFcK7azOCy9UJAAoWX2SiRcjBb365yf0zTzLdsFYdyKMjWbPixT34kZ1SxgQdHg
iDCRre34niypjmE4dF6zcVyNXL4kFE5yaiChStnZV4Jy9UvpSshGAm5n8aPDJEG/weLkJLW2AFoU
fP1tt+69l5GVnL2UZkOdj7lgVLf7fCn9jhJO4n+Hj96ikVXXSFj9q0cuVvpLbuFw/pfBX+fy/vjI
mkpj4foi9UQ4dDyBPeQKq7iOK29CJwjmMvPU2oURuA90ciRH3yGyvW3YE+EuUD4Uq2vojB8hZC0I
ENnI2zjwBVe93gxNCb2Xjzogg8YGikoKPVgwVzNnhAaSWedRkxql2mRer5r5gMOQoqx2LNZs4itT
0gmEzHYcGLhp666Pgd4cGOJbi0Mt12W3F3nTR1WwN7JACaYGjL7nFFdTWpoGCxYbjJGV3LpFd36/
XkGyul3dsML3iJOC275xtD5bYWvsTF7w7Jyt0W0unoadx3KKbIcVzBbNot8B43dIxtxJ0CEtzRgB
eW6un5jUAzu4vDuFoBZtFK0VS+Wdks5ChgxqNnhsTaFZ3b9RUDMWf++Vo0UrksMyO153ARGoXn9a
RJa6I/62JVnm28de+6oMyXSHb1lQ95CbMDizdBtDhPbEkDhBKqghj2enHMBecbTLGLVUc/M2xHqG
hH5tglvaLvCjXSNtCR7eaj42UliNvvjJFDfWUjrZBAKY78U8z6dfFJdWdMpvwFvITJGzPFlXSP9g
f3avuQQf33BZPSay96jcaJ+f//KCZcIYIlxSWxEtIz9Jeikn8Dn22qVoCoW0rMze8iqODg1+7YaE
AsCRvmLQvosCgQDvilg5CwgD2b1xpjXhAzfB8QZ3ivSfZCBVsxl3wrVaMz1IgBHGj+3gRytEBN1J
Vfp7scshxZrM0EvN36jMXSuo6Kr8QYXvt5Sfpuo2BdTfOOaVAf0nMwSRQX+ubZDstJNmyny+kCOe
LdYnzVyyguPQ7bRB2tmvEy66n4kjiAd0xctXL3YAUDKo5DQhh9QAaKINAndMjTOu9hA8pgpGtV4P
J71QN4TbTGDAwUEZVzwC3WJ2X+Xcxw/bVgJnHQC6Lq61OFUJmI/858xpCPj/ANaX6oO7ip3Sqd1z
X7jF6s4abIN9S65UO/Z0/I3W6ctSZpOb8SywjqhrVFgApSRqWdRtRlA72lKG5F7WQ+7Si/KCRrKv
6/gnr8EnYD7raRDJNkcqeMO1DUdAXcDfYBNcQ1RICXuplwvwQpsnbrQxn5gixbC48A9neg+yZP5K
fDIc0ujfYQ2s8jjp6qp1yX3Iv5jAjjMNUrwPWpk0gmjTLjty4puwtdg7CiryMEMpNeZn74gIEGRw
eR/Liex6T/xMprPBGvLew52MXAKkqUVNnrhlDnsRqtXzoibkaSsk6+BqrFZBnaUobykEu+7ykRu8
58iMY7Q1Kdhdzo2E1llWk4FbQRgGg2CsBum293fa0PuDy68RyZFq2ORe5mGycngfYg7Ow3YWcnhW
Uf9eyrrF0CJ6BrXykTZlN/4NMNF8nOEJk9oRYCawv321pJ22hF0JZnRSF4CRa6uwSs+FdGPSKX9g
IRmfEwEs3XlxvLl4Ucicx55NAK20h7SD7kkuSTCPs6xvVYwEFrfJxCsYprkmdna8iMrwfc7uZftv
ekIivotSsGlgNzwZTLpX3WMMtwHYRQPusABOas7mBlkqezGzYDgwXpRTpIs+pXR0bud7Q7zDkD11
tVAfHlz/GIpF3lHXFvrSLo7Qp1MkLJkwNagrIbfUPTOY2ue1CGpwzHc4VRhF66/VcWusd649aOLy
uOX7u7Csr1rCM5USiPNwBJb9R2tKtWg/Aw+tt2FxrwbDQscsOiWQhpv01BGSTh6aGMIPqoTp0pnZ
V005jVkIJXT/3FH5LyxwBKQ06tDK0Znfk9+QEZ6QD7NpfFdKreiAryrh5nOGSD3cWAj7vSqZESeh
H2b2Cdn53ckWlUi1fQNSUvfCQVKpOyhRE6rmGaqu8MOl7UUmCaE1Ay4IP+XwX2SJnfwL+kG4NANw
gedBvg0yLH+BeRI3qjJeSU4blMyLNrPZLGPNAu74XFQtDRsWLLSs2yFzHBCWOKngUf9n3ceaxpYW
ed0tqM7M/yaD3qQkFMfAwPNqVBZxj/RaeF/FKLE3rKL75mXrI3EHjHRVVRipV7Srx4pCGv3w4Kul
SmLR5cXMj27iGs23VR2VF9xZJL9eNIFf51PhW3PutBRv0JzJHTugcR/8KvOC/TLncxAu7qqi0YO2
mK4HVaNV986RoBzvf7/rYKo66jkfZx64LcAL72/LGDZ1qT6mQyI8dfEB2V/TmRqdoSj2B8/GGjRh
4rVjfhxNBt+VdvZBcluA2uvbfP/y19r9iPLesxUdG7gQ7tzMGJkeOjuvfRloGwbumuMXophtOyIe
QssdqHraMkwTlasmNOcKNypr/VZkklJfwIwdrUHVhZI9TYStCcIdSB3fE/hR0OXeGhIKwlP17bcm
w3FW9whT2js29h/LGPU/pOsXFQvxulYX+gvIbs96TTORDSEVF8wruIYWtW9eiKPOnO1KRZ2JN0zk
8XFx3+1rXaKFN9daQmGE05EHX32VGLG77k5x+9xitJ9kqa5XGuhJUX6y8nsqEVscW27hwtXB2GLa
wkBIt8qEPXaWY5qLFjQ2yqSd/OgmDs0MWHWBR98na4/BnibpvS5Ri5QZXQ2fQx9/UuFsnov7R3l+
9w9ylq+9hb/BARybVUgdXFK0NzcWq14/nO4chOjVxYng8iHL4T4h9q+QMwPedD51B4LDSrr1mP/T
0OxACijMxbueVjB/3AZ2QQ3KA8lzgldUr77wKdOZ1wW+esNzdNzNELptX0MdbbndtR79W5v2/u+B
yOqzQ15y8a12Mgzp5nDHEAxS4OFv0RtTdS2NBfTqm/PpotSpaB02mSRCPfE+fragtswUwPBPUHEU
zZPI08XtCWB/qfJpVIhjygL1DYp/qUqhZe6myZN1ngVfWIJxLVz5UVoR1yObYwrBcCEUcEhjDy5G
EamnjMWGKXaOuWs3KIj1afuLzwaiz++yQSc9QsUyLqWaHinhGjDo1uee4qpZ5CNe2QhpTDzg6RX9
rJsjKKCU3Kg6gO/DMr8iROzAQKuqujO/fO7i2+S/CJggu5Cb1uOVUbNtqbTiIBeiYJGUuzHsKu3B
Zn8evm2RbhGqDJl1W7op56rsxlxo43gIVJcVxo02UQNAtGibugh+VXZBeJVxaTh+PNoEk7U0RJxb
pg58sIm+Aspo91RT7iN1q12oBGB/6z4VD2uYVc+/bWnNq61eMMYt5+NNwmLiisB08FHp+RR7OnQ7
NRPgRCeXjEhLK43E9WJHWBHXju0+J7YrGxo6hatGszqaM1NqYBrvHoK5Ijm+wJRWPoXgZ839uWHW
E2rb4C6qn8VAPk/x8QrX2m9fZvs9im7JpjtqJgTLVii26i2NUeIIynMN6HCl4jkw3FqTNEP4uDip
CGU8J4GjUoGorqKb78pJTJqZeyzYkbnO5stNmIMxYTRA9hm+tucU179paauJH7oDWea/fF7Xkxth
imiToGnfyOU3xwmsnSdViuw+NJQAXP6OL5hnKiMpAl1RIzmE5RijS++nPDbAlpcEDRsvpFEKwllt
IZ93KL7mEi+F7JOwxmJKWjZS5vp4VcHMtjNHl1uBjY5xQ54SdIkYBVgySblLxmw2wO1XjBzAKnqB
elsDLT8UeFVKaCXxQX24YC2GYIQ+p6qFhrSi7p+EXMfCUEpB71bTJyJprhEYHStKUeu/ZKu/E90J
a6Zmn/cx5nSgcHFwx4ivIwgCoSYu5FipdP4ZRtKgPKIRL02W+U1G6lubniUaAw7FBT0/4f0X9z1r
Nu7vwu/00DzVr6WknFjEYgmQU9RfWFbtUje+Tzcp1g17t7ElXAHvlOprRCNOPZlDMT7IvIlWnwcQ
w7gRG/aYw9R8VqgxP5SlbkAIbB2ZvHNf74H6//7h3cMzuQqX5RWdL2H8meeqpaUdJ/T0/bXYZmft
upuM7Uud6d0d5K6jsWrVRSoipMfhTZ+5ASmF2skvOlBYI48jQOsQ0raTfFd9QbxV8win0uKKHBsU
E5fo8sebqnkO/niugdGPooBtfs5VKDTeF0LuuBQGfkve849qGkfBvzzzTEW3Fn5OBPIJkMUTra5X
nlhCAy9V39r+FZm4T6xKbzAp30IgvikNngPi4/+whW1NH0XZ43r6EU7GuXv5Tj3BdAxXRTUFQU0t
uNVGZtE+6hjuB4nuabrUuSn01cmaqWG/47IOKCF0qDNwkmYMW/rkJ2YB423+GwOiheUph56Jo7xJ
MZKPuBhMyf2ZeMVYWJDPP6+GXq8oE2S4oqAEWIt7lMtCnUDaN7mXZ5WaajOksUD5tKlSe8kY0AzJ
/FHEBR6npypjKUHCdhHSwYZl9GRZKxtNB1AFpmUJ/l/mUj7aTG3ijNQ9JjgHkKR2wsrBL//LXTSY
sFu6YtD2Wosg0ExKyRmjHHkVgaDWwx6Rf0Qr1TngIQORUBuTZ2NKYQtx3gBF0F65Ko2VJaOHlmcn
mZn6M0O2VCXv71rretzrx+deXimfuPHK0ZZlWJ66FK6jV/VLzOY0rG7H/UApiaUXiYYSou5DaodP
8E9LSzPQoEcjMaLn04uInRF6fo68apM9yPvZjHPhPZBXuk1RVxCg+RdKoYNs/qysLC7hlTYV+jvF
lrlroHFkEhGyCJ/9m7Sg3w4JTnO1r4ErtSZO3EffHA3kMrMbwWDu7R0aLBw7r4z645DygrqJiv6X
+1C4DN14fz5kt8HgAcluWHJED2RD9qrgUHcMW+i022v8FR6Qxhydcy593RveDrf5L06Szu9QicZs
tYXjt1/z6vcbeaR3R8cX5pks2hM3tYZ/mpk05DLK28VcIL4h5aLxZMQvyJMyMRI2dXY6Y6wkXkSD
AWahMQoVB9DkZI7iz+Un3SB8S9K2H+V3SASzj3nUCZJygogFlsOUlergrWce7wulxDygz1Zc0Iko
SgYCfXoaeoFTCxa3MXGuaPqvtEmOASqkKHzJv701e4jje4XHs0FlrzuxSpCXyZSh6O1OyJREz8UN
8k2X7zeNjkZREhNmQjzUD1D5zaeePyw8olx2hO4rlkn0uHasU3Y9rMdHRfezJvix7utNjOGVIVO/
YwFCbNk/E1iFZ+CCpDdY44RRO7NNa0olDMOEgKmokKUaLKgE532DVwXLGBj03HIqnMjMPVxAXaEf
6Y+gi30XCcg8bKC8CXZE5dv8b6+tbOzNeb98NGIkbTDiGBmRAd1GHwuHwM7OeTcVMb5VDmXVkDpX
dZa6OQVz2V4sHN/HgkpwEWAKP5/nYRsraO07YjauAmrdfmDyACxXSbGDXieaoKNnxeIuAu9QInEb
ucVQ3XAhqu6B6yCqJM7n2vLyyP4t8LVeGneu2uPftVZ7kKcCbE5oFczzQ9jdEwUw2BQaeuTQjnQg
HGlu7OobkwxVCoBSAZjoqG65EUwrDRRhRKI2IDBUL4azGkWhnUVf7gJkdFFyCpABH+3X6cCJKDIS
BmPXIBjUT4fgco1CyR0hwxSSBzITny+G8cZSpoPxrJAP5NHrx0j/3K2+Mo4e/w9VrGdz/mZcBK3X
2CP2FOS4nXIklCBRHSUzZui4XfpZLhDM23pQuU1VDkmm0u2khknGWXsiN/VjdgtVSHJhsOpO4Ix/
DSW8f8HM9Qdh3OIDQWFZhHgK4yH8dadIJ6uAyqLPKatdLh4DCzK4obY8WplkP8rXzBoLE/mTH6lX
H8cvcFk3VHV8hqOrh3Qvbzcg85rps/XEx1H3rWWY1rDCvcVJ0lgEOc8f0i6LWoC/W9MHVThF616O
QpFOU0uv5EJfMeaILPdYItjx8zOdF89yRTPdcrvZihaylrniQ1Y/RKDk7xIsTiX0nRheay+wQofV
n4IvajSXdHGhtD5r1z5qAmJkAA03bDmh6eqnTF2h419+aoDz5MyAZLcool7rO84a0aamjMFNAnZA
+1f87pL5fwwlkSwUJLrP8nUD0ph0+J9/uqDtA8GI060KSaL/VudQTh4+gk24sEhxU5EPz7xQXeSo
ugsY6rrT9OyAM78IMA3W1pxg+JPn7/gD30/V761UhMnIVrSQBjTAmxdECRXIOa7NDMKc3ljUyRvt
aA2TEq7deTe8m7nNsmeS5xAWq2xmslJcARFMeW+dTk8Sx4/jERKkBxddRQxjJcv+OhUiqgsqQ0IK
msRNWMpf5H989Qssi7fbJc4ZVPYknJSc895C/Ycb1CwY7xWuiWgWV/uYgdOQdCEC1G69jprzleNB
LdieScElOyHqhlB0cufPCe+X1M+DULjSSQii1vU7HKLnjWVSqyVJHcE3S9E6LegM0mK03fB2HySw
3v2sX9VMTzLD2wUaoExwPhrZ03J8tik7fuo/mReYPGrIzc2gglA6URK1Aw4SgEnyR+1NKYybEF4C
mAMgc6+A/naj73NGYva3kaJcUubo7TPJRI5RVutCHqSUEtLSCu0YLhv3tS21rvDUyo9lmiThlumu
12iTx5Rd6y4lOTPQ6D4qJEJvO3tNuKwyZ7dkKzMXYAqrEBw3DJ0+mHviWwl+dhcZ9KvUh64IrFqP
Rbkd0RrHrL+3PbrvM7uFvv84zAL6hLch0kpN37tdjOWKo2bgSCj7wh1scqK7ZB2GUOX2nyoG6eQ2
OWH68lXcKepMn5nFxxx3aTg+IacSscGHLNrNW9fLhzVJuZeGYTEeCcVXE4BLJ7ptAlWDpn33PTz4
avf3ihtmGG/jqwihW8aEAEB3ovmBvu4bk7EIfxYUJs1dVM/fHrNttLcjBDuKX8ONgtz/hVhSuN2j
LXTp9obflbXjsbVP9PCi6RUazGH8v2naOL4LUdpFi8HQ7cbkWmjeVNlIqrmRx4wEMKH3wQDnQ+/Y
Gk0vdxuHoZwLOjhMQJRWsO9rlKTgsMNR270/47LQXVWJ0yqPmtno/GqG9swdTg1CEwvukyxdRTiD
a7qMM5LioH1TsbXNzuILJ9/OT+qncsfs0xL1VyqXM06Olr73UafU1O8GXzWXEvtWdgoMdc5ON8A6
hPx4uzJieOZOrnUEpARJvwiOrotVeOVEJpFrkuuqTuWfoJbYN+TTUbyPMthjwbuJg8pi12jlsevH
TdyHiPS9arg9CZqk1aI0AmuvvMZtvXybZsA6prDqjjvt49LEXCXa/BkrYGe95wop4Hyi0JzGN17i
KCG8VGNXFJLNKoSiIaNSbFBYfmwc/J17YzNATvsOFLrReB63JUbMNr0UL/rOnBb58TtSjg+Jscfm
LNTsyxKpTEqYvLuRF61cbZWuvxhjzQ3fKVzA+hTLvQf3EfXtK8xUa4tDEBHhBRXjH3wr+n/0Ravd
38ODtBB9YfAkF/gVqb2eqbchv9GGvjDkUPFlq9XQpmLKBbBhj4l4RTrJ4obBeuGAwRKyfspH4Q15
eCZeAajPavcnf0/2mBwfzXgVZF7irvLng5NrIyI+qGxKvJ7uVQQ7h3dMKygyrAnxf9q8yfsJzNzo
WqM9eLlQyTN2IhssrVCKRRQ9zHYDdJcYq6jCYj7I1zXhQwi1WvsN0M5tziPPhPCxmMpqeDhY4GRn
0MDn5HoLWkQa3i773AcTgHmUjKkTWcAbzHZSRffT77QRtF/HP/XN2Mp+orwapayC5OKXNfaC+6Qa
sqUFnPRsS4YO+1GkRJnZ9YZqfQ9kD3nVLq/heM2AsCfnaPG/ByoHMVtquoF4UAfnFryhAXs+d3fh
QrW/0ZS5hcMYIF4UEr01jh193ZwBn96nng6oWzDMSruJ1ZBAr3y85afQNdW3MyrMSITexuAT4iNv
9cFC8layvRcWFy2uzFOQSd0fm7YYS9HcZ8Lx6ZKn3VS1Gm6fh/PcwyfBNPgNP15SWv3vK+zA4wA=
`pragma protect end_protected
