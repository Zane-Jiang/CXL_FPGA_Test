// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Z/BvjoSdYnWlNDci4qKyj+RrjysFD2ScuWd782rYweifqmmgPuN2raKGVRTn
c63/SX4wwFDO0DRp/GSE6tDE4AhCUyYWdyaTFzVroklS4P/bZv9xD90B6gM+
JS89jz0ZqZb+T4ET5uSKApMMSULriAagVCC1WKVK/D5/YSko+W17sjHTiVaC
OC+GTPkJxGUAAmly/6wnQr8Qm5dlwIZGX0fvJHVQ7aaEMVbg1S/h/vYOql2P
BOphnFsA7x8yObzz0csr7Cxs3KYc6kgetEYRxBAaucp4a+IG1brzUMjYEPgx
3Z/LWoWI0M4JDPfJyJ68dyIaomtBotXZbisTkkBlmQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qeg7f432vs6nDImIVELyOfWwrmS5iw/r1gttvstueBUQEEU4bzAOpQhy6c1d
FSpOs/1RBVrCydV4rFEe09Plm4gTRjkSPV/31UXzzREoMOjY55SJq0gw9YLL
Yjvuk9s4JWrRot+sYTD6NJDjbspRHAEU4EXZ0VOLGjd6cY9k6q/wbndZwbiy
VvgiACjrWs/3FqSqr/QO/zBt6YD5yrpSwK5V7sYUNeKdkE1HK2RenmsZiuvE
B2AtIRQzcuhx/SdyK0y9FwdtV9YDRsGER17SjLCQ5CPo6MUpJTfyh9tZQ8OB
fslojEAwGEb15fkKOmoYw/KNzBWtnHc9XORytX3v7w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AbShzWsH2tpHw3Whg9K0HHocjDxwfgvNFS75YphtBdX5hJ3gUC5Io5FecrJP
xvPsZRaNsOT54melLjq9dzFySNgP5yITdiih7FAUJN+2Ha9Kwp98qskBSlUs
TkN5zrJNOSkfPeDjZ+Ydfxfstu8YO92WQIo+P1L8qY0ePb1LjCqL4g64H5vY
MSk3RkAnnVSvZVi83O1B8Qk3zUgY/4ZvqBXxjExKtq48OLCl3l0EWbr8Ub6O
iVoEaydTxNE1szhFj0hBbMRI+X9EFBrwRCDlPDjZgaaU1QyQ10nbdHqpFmwY
7Ba8khhArW2zx7SSII7/nREApe6lNT/+Km415/XooA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fdnIS2p/IkZDzBZqW5gLVfXQuHJDM35s33UWtQxpO8NVOpOL2UWFxX1Rkynr
ztQzdD4cY2+bM25+X7/MxTDhKRnw1XGd5ugMHv+4SWynQsYChFuY9866UNBa
m9IhKldYRkRRWqW0mkx6nj4j1+tSqsVxj7b+xfLjmxriz2nNL3w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
I9O8grU/w0lAXc15zZ75qXZ153zl+voP3KUEzNydugHpcXwJBJNrSi3zzohW
IjJAcCHaMOWDPnMqqOhk1mP8OLNktN/xVwqNd8CF5PrORdPJoDP7hy7tKrnV
jidpFew8mpY66osTsqhMFuvcOkcOpKbG7fnaI/WBvLclRipYQam7FjTwzB06
wIgX237gLjgoRWJbG45YsGeEHojwjjKqk/kTEiRnN3YTlPRjvqndOLjPRJXa
UcPFCv6ClStHAqxEMNegvDQYmax/zAhcAh3wqm4nrcFDtQVmUJO+t7aSF5/a
yrHZmNVJMFw9sR+Y5QUhHhLeZFw2Whjd9fQJ0KqqwaUNdRoBlC55mfg2bohb
YsfcZ/qiGsCs9wo31mmbZL8Ay1jfBq9pvoVnhQzXZpyFEHVIp4V26C3UJDQl
fDBxOxTug2bqWa10C7Q5Fe31Tp4JNZSLXZgDpexjZFnme4cHhZWhyC4K8iI+
ibZQZOtN3rIRRquhegqyhKRnedikRJoP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nglNHdkmMqWBzlG32nYTxL+gGTC5RLs8iEkgo1KIWsZxzn0QRlkbtsdlDLwG
gQLwIvynesS2D/Ufv3sI9pWMKkmZRG1oFFdi2BL2q6k23bFLQlxQtj6M2Sn+
A/ON2ny93ycIbaU5Op3i/lMaEYfXPike2NF3Jf8rB917G4lf4uY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qf1+fIBaE3iXkBOwYVMAmna6/ZsnAo3Cp98LsnH89KEcfFeS2/kOpVtrBPnD
YTvfY9ZXX9RWM8HK+DQXFNM84jY4XjvI1KqMGKM4mKmPGJvuwBjB0CDuZWYl
SnJTVkc/od/G8fURTjZCCS0/aifXSCyYO4ZaJbiqjAtZxcWRD3I=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6896)
`pragma protect data_block
sL4yKFDSGfhmEZd/UpqqQaxdNkM8n3NCt+w1VwmsfXRCufAkW+kBqpWCh6iw
Uvwnq19HCBANG7qMJDRB8+8JtFaIRt4POJYahMUdECDhswxa0Wqs6TRepkZM
5/9SvES99SfRcOZzdSK9uvx9T1v4CNd4Ixhb/mYaGp9L71CFR2CQc0jqCpSz
gRWaqmRN4/SPFvENEcsTosccx1kwOtVnaAPm7Sw4UimuFmHp0c/NsED41G6Y
l5etf3F3Uxt5hQZ7LEqTPM6C2CEUm8Hzm8MnzWQyWy7ApKLLFTRMcrJHbLg5
GdIXcqAQC9rzXjyE3wiQqWXxAzqypT23E2Ys+QPXeX32/Y53YgOBnZDSVdGi
+Lk2uTtOrkuFdETaKkMfuy1igIPYS3/miaPLTY1SqeM0jYAi4Fg8D4+vPRP9
4fDe2WklZRtcvsS6aPtKIdqbiIZiZA2yZWzCQN1Hei9C9bGGZwhduI3ISkLL
WMHVfjj9kXSuHZjLu6h/NFKkohnR0W+bKUDc+b/XVMW3hvUyFSm1f7XUd2N8
f5d6irHFiXyRmRNcBP1fHhRBcTvc7qgGi2dgN88MlI0hrhs6RIalh2TAQqR9
Taovmn2TuN9JjvJ/rQ1iYr9H8ZByTNFFMqucU0QYVvG+6gNrCxMyX9MSj/m5
uqicwTt1upf54UwmEYLw8VUFY6bgkTMLBYCqX4boW0crGQiwuZHzRavzYCJo
QrNdWk9jK0DxSz7PQyyXpK/qhI2wf36WAu8txbk10HY1xLNCWdh9E78NV+9j
qnjUfiZEfIL5fjCAYQ07/JhDxE/d1W9BoeaSgIWc3F8j/AKCRPRGqfqT/M4E
0Be5cDyBUZsuvplsdGZHusnH6ef4wTQbXjN6B34o2OqtllEEtSMk7wM5ZJQR
KTvKF1iRSy0kghaWU8VHSoF5nG6bYWZv1HSHDIws1+0xAREN41OgcRhLp7qQ
Nwd+ri3iEsa7D52464NSgvG1udWPHZwCCWWZPzkYwMvh8AApEfIDm1P+tl5g
Bj2B9WWZu/RMKS9FkfiN8JWfpaoAu80tfS/vUvdqdIlOw3Q5+AXlW1XVHO+b
1V5n0AOCOBD8I/eTVsdGpivQEqNAHc2xgcIPHGyk1L6rvyuGTQ5pBR+oUkZr
dDrwOzYTKAgmAXaxsfFmXHrqj0wTeeZkBUqEo6S5nR9d7XZI8ki6uOn55+tD
3Th+irb2/6t2DddseDrDOdV8B3E3GQZ704tcEboRVfr4pekMjJFHKrCgKTAx
40Oh8946sY0C9TYNLvvAuZdTfo51Ctp4ptIUK1PR/0cIlKuujx36phciSapY
AA5Gj0scBylE2zEJEeHspw+umDisqix1m/I6UFrMBoP62VU7agUMvylBG9TC
0ipilA9DDpwpdXC9SkrTzhkQZpd3jtX67k7emEh644OrDYz2F+sb+U4EZHyM
BqiD6i45qb895K+BRrHpXKAg/IfnYLqJpr1Nbz+0VeCtNUvY8bstW5Aj7Ws8
zi/kucDTrHh4yDUX0KXpI1X/k+2KpsxB5aykLWYagM01tZp9MioF4c23ZdXf
GiV7+ZOMzc52lvTIqpDrSP0Pd6On7apYzkRbf9Lr2YsH+wtZYRVbyKwqQX58
VGYlIMFh4dy3PoG1CUCjKsFsIcKV4EMfQvcmXYAIWPl8ln/adEds6sybvI8+
bqBle1c+K4dqTpBm/oMSgwIkiUKUf7aOy61UFSkpcjoLDRjz9HPPOzfYbJXF
8XNIUiQz9kIXDbj+d3tXR/gf46f7riMDlHEe+cad+BqHHLSg7Qgs678an6lH
uFAdy/c5W/8YGpupLqOR4TvwLyKUmrqf/O+10DuuDoOWRIa/4b4uPOrFW+5x
IQroo08Mzy3C2vAI6g63q59N1xdTj5xrSz43ISG+ZbzkmC1oJTfv3fRKYoK9
5iWIVMdFkmodU5r2+ApznPnb8J0FqqS/zTlDDzEdpwjeeILcCI7bRo30Nz/W
Bujbc+uFqiRU8CDGNc1j8XH3+biRNf0UdJOT6BlX58hDSZX4/OSoZewnfUJs
U59VWqgNZ4nTH6yqNQN1PGcakv/Fn144Cx/sI/ay4QZyAqX1UGr60s+mL+wi
jZWTBlIVCc3Xjv93AULK+8XVqsPum3qALsxMCWTsnodZmGHeEFrL/dQlYJ+R
OTqyhtXYD9Piwbrg1cKLBgLDPKbqEfmH1OA8FHfUZacIKfQWObZehU7seIQZ
sEo0Ueqhn+4Qr3qEd4ToDPmhLjsLpc/Ts28urMU2yyASB5LwUWZ0TitIhB+S
+8sf8E4Q4BGXSun9JW2JWstLh0MZV1XIjCLdozYZyNoRhMNzcouOI5PTCufd
bDb6p2IMZtswPXktO56WSkVKBs/8cp8apwGtDg/+6uNxWRD2ef2zGX9e7lJr
1QhAsO+NK7FGuLoJ8Nnlgz59RHAG0bDp6gixMWOUe0pkk7rGVKVhFM9sgN0l
mqDwjYen4W3nAyBtpv2lx/ss1ltzRAjp/nRHYLuBrCNrtMtKSmUCCQtLgigH
jXhIm5+MfSNJKQpMR8JgnBLiAygJODmPHE/INsVrXLS/dUUG9zEl1S8bVKtV
+S+oz2II+mMzyAyxjBqRsW+ZHM2DZ4cmQrPVNuJa9LKoWnvuGdXIpTBxTOPD
420yzak/zwFdtGXyH8qCaLLws3HUzR19BEKuKOoAYkSxIly0UHoxvikAwHut
JGGfwgS43w72lPOC9UZunrp4DZ0naxqdjF7EU1a3wQn5U2g3GTaXaJeEeDuE
hxKD7z3Kr0bdCPJJqh816OiCUdACZ34gfjG9Q92vOjrfGNofxnocXxKLt9xl
HV0w/hn4MLkpWUwwgMQ8HHZN3TG+v2rkmUTR/3+3P+xZpfhc74t6oJ40KAf8
nE2NvrZi8dowZD0yWkJ0knwmv42Oa9YsKB0Zas61NgR8YDxRpUye231d9MU3
5kzW5iPpkseoUA0SFQ1OX7e4oi3vdo6/tFd5q9EJb6TJ6qz4OlD09hGZTUUg
NnbKs/phO6a0dp6Fjcz4e9naZFtuP6O8l0YYB6E1DRnLQwbu0BT1T3jD3w0O
H7bNfeBtEEu/uzRqaJWB/EsszypnvlTXjWch5h8/uYXy1Bl2i3GK3Qzx2yQJ
bwkvOh+wGhfJRdRZxhlB4y8CCgItb/vx8yYZuD8tdfJykqx5G2OzTtYWN6ec
bGs/WTodcTLjVv4ZmnIAX4RCnOHKKMxkjfZPCybnbOCaOB7fj5JaHkSDMZq1
rRpI/Ta7lEFbvDDefEAxSPj6HcnK2JWKqoqR8sU6bABTADOf5Qc8mwDuHVcx
zALK//ZR/zg7FVEVQOdIs987AH894SiD9L75DHox2+7bH7+AgsD7vp4tHV5Y
ugigPpdnPLkCuyvyF4s9S8mzDSmq9E2nWY5cIwmeXNQzgVeqOwXu5AkJLpy+
poaOvImxX0tvf3wYyfxm1ConVhHISCAfUgHuNqfU09xE9Z88swQSDHb4O/2J
pzNSzM2sIBf55Gsu1xFXFhzG+wSf7ZHFmP0FdR/aLIskvVvva6nvdw3Viqg8
CFdhoAxKWjEtVLq/Gst3Vjj2SInFdL8yznlPWV0AfWJ/gi2z9KPTGmwCMiCN
LwmmSpoDphmvtGvxPV4p/nJ+fdPPH7etVuGh9vHvXIWBxWPjrAbErQGuxhP3
7lkR4IccnqO4xpqg3lFYXBeMT1ER1qC8hKOWVachPU2aa9IkEg7YZ8LeqzDd
teTZuy+8iaelfWxhJpPOQ5MIc0DCOgdmTbScZ09EQ+0LpyImAsoTHrDFVbwY
jr4+Q6YGvWcWJwRuA17U893kY+YdO3C0+aSE3P+B2G5YSA9BHQ4hWauthOAM
Oo9qb/nvGPoH/OoCIdFhjPilEqGVQxKM1zIGfVp3tid5mBjmlg1nF3iR8DYr
LDqYJxPgUxrWzJ+2SFaDym+5xUDwRijFYRUOJA/VKERuJonuRQ9WucPZF237
9+v8CA4WBd/6zmEA4nbc8/+pjqxz6HRaf//Ws5nb79+54IXE+bDJlgr65i8q
Gt+leBL0SdHR3nb/INATFj8/YAHH2wbDPqKgzNAfLEnMiqCJfp4w6/2wFB8J
IxI/amI3uLdXRIE+gKqnjGnKtvk7ANH6iMXb/PipLLJkuM1OR9nVvSmnVvQ3
5yHzvvYMSffq0qAXFsd7dWYTRjCpdz4mypN+1Kg+Y0YxrCjQJTjgFblmb2n7
lvy59W3yj7s340eAYFgG5RD8TukdwTHqWClJ+1tRU+5vYi7W9Lqmv4GJEXqI
4FXAwImAtL3pMIqz0mX7BiOnnxBgdVZP3NaqLFYoQs0d13hbj/e8QziRwZFq
TuLbcoLkXMGVAUg96iBFl545moaN3KPCQ9ZCxY5YjtHhmRb3tyjDYVHOrbwf
GwrE83vynFUigEXyVC0mzrW0tKGgKZTuPdP4uL5AOgvAbTk/gwtyDYCk5ogS
NQTuBGL71kBgR8HLegpj7L15lKYvsdpqdm5lfWlx0fB5TQKYkfVYFyiyAOiM
YVGG3VeKMQa1Ef0uR0NaitoUq0LH0yr9W/awpO10BwEozyGDSBMjvn1aAqcY
TDEc1S2ZUFMhlxNlgi0XTdDsNuqnk48Gdwvdb63Xej1xM0fhbTrOgR9s2AUA
Jm1p01DniHAlTCc2P9TA87MMnRrLLNeZba9ZmnwQUAw+z7i6pEpXpVaCrY2s
o7Mas40MDC2Iu4P41knDcH8DoCIlMF64z0IuoU3SPRsvuGYAuSiABu+adCyf
TxgAE6zjsbBiCTYmlrKYQhU4oY4MyF42LPg0o+WFU8Zt0BXx7pGL4EjWUDdG
nhI3yuvMhjrwiDX+HLHoZnkL35ERxXUksXWYihwgIk8B3l/cGTEbPhRRFN8H
8xkFXW3sQiXIFxL63EiP7kjBf2yljSkwj5QgntP5tptFo0Xh1yOy5dnyjejj
KS2H2JTbrJCw68EXMI99JlhcRynouMVxoAe1pEZT/+KZljjDedldUn5VQWeV
5ydKFdCSnlP6EXiTpPzeDPaDWKEtxS5DuGtNqkBa/qcDtqJTMD8cYHCyeb+6
9ZHbza62Kagxn7DXA85V3Q5oi2aYxT83Mcb9+fjJiiDvjpAWS/zUcDSfPsvU
/bhEHEE0g/VgHvwgh35Su1Af/82hbYz7UNUC9rYd2O1QAyeJlUxVvKdTHWky
YkEYZA3gkPNQumSPn3G8ijz9L9gHjQUs4yq6U/ATavjrHulF0DcuXrqK8MmP
vVcsnEXD9hHx4aIEB3wU9r25imS5wyMhvfzh4VdaUwWGCQbS3prT5PCP8UyO
qtZQgs0jxW2Y8VMl3mO4bJW2aH275X/0q/gsGARB+LJ4alHtqPMs4Sjr05JX
14X2Fo3ux3/i0Umhxti/mTHPrBLRkrw6pKHSwyhLJrE8PaQwyndI57LZ0SbL
gvypippN5/dYGV7CIfbzfgQ09znKYJQ7J8FuaiN2dJUy/gGB/Q3MQTFObcmf
LqWAmi524iZSvVWeyI7J1u5jTPvipOsNDJwnsQF0DCpXQbbV1fHs022bhRtm
QuB/+RdPo0jgX+3Z+zT+ZlR6qRDiDNIf8MSeF8WJbQEaVg7EkcGX0L73N8hf
qy6yFhnJk86oER3qikHm05GHGDDxUsOICQx/yMzlyGt2IrntVXmGvAHbXI/a
zxLzzOkmPcv6DooRzKTSM08U9EKcvpX/Hty3KCexFDDXLfBv6hWiAoufsDcy
soRYmDmcMzwVyIMhpe+qQsiGlbCXEvrKvmDUPSkl4hKYoL3Eg4vdushbKhpd
MYgZVRmCA4SdPsA+C9lVZM/sZQUAikg0eY02UY2PfrOWjBh9t2g2dbCuihke
Xm2omtI7Wd3lROiuMkiKGJ49SUittNhDYAMPlkYsjtic/Xdz4mKO+GdTtXg0
EFu8JgYCh0fv+FCK2XmFeOAN33unFWZA94+pm7I3ct7dxKmxYVa0qmvF8P1z
QmXOisozL9N6ctKrQKS7ydFhfTtGHi+EC8MX+OaO/xDeqvVRgPArN0CU7HLA
u09IO4a0NyzdFRjLJSrRyRtpxfd0h+bs4xe8IBlFZg8uHTfOO1xMfAYsCV74
p4jxsYHOk9dNNXEguRtJozZpR1jqxOPNcbkd89bdV8yWbKiMo8+81ObxzPk4
abIgkQhBVbnu737QkJuHc6oowFWQpBYkXEMEauXgeRKsffF9TgizJOc0TlxU
yUUVxApYmCi5JyELV/7GAdKFLaJd2YJ8BibkBTULiRYkMz9CYgTXDTwHumqB
I7/oB2i9pH4wpZJ7GhV0bsVFT08rTcgBjrieaIZKkor0S2KLErlWvO0wsaue
x1I90O+rsET0JJdAaYCzCaH7FypXhlDh0SykJk00tlaQjdZgsg27WVcnByQh
XvYLa1hZJHbur8iCnAXfyhatWbk4DwnkGwhTb8HD+PBE4D0FM+sz6cuZfkaj
wUiSFi3Ebiy7jFD5dwnQPjvCSDebbgWX2LgyUagsgkl0s6DcnA5UH5PPlg+Z
y1THL4XB6uSo7B7qjOvHhcW/OqaahNYv5AmyMW2Lm8XKnO3M7lbd88g7APZh
iqHcwHpIsupl+r6y2SCN5Uxn8G+PEs30fhhu03OnE8G4XotIR9orvbv0mYGX
ZWXmhPs/TOemJbrkoZ9+2CDTWIPCZmSy2wvGA8dXAqLn/Jzd8nUytBpvlDuB
H82Ja2cKfw+HFcnq/xoHnUcsT5G7kyjm6Web3uR4671WgrsE3sQYkZCWXFXt
bQRiHybvldPWOeBHXIQqaozqG/R4bblraj6MZ5n0tE2hDE7Xheb5VIBLy4Dx
TilP+fmQTXtHbQWup81i092LkcKSFmod0ulW+qXP8LCqk8EpmtM1gsVJqHM7
tPjPyWdpNsV7YP0fLeVs1NxrXIsQI7J4nSLCvO2wBQRYyDCSldmuRg2Tr/pA
MUc5komJellInQG7ulAY3VlOPvC5BnXeWmvbkYij+bB7ZEiT+4Upd1dE5wOU
SDX2C/scQLprh+kmaBDNK7Z/tZmN6FFmrd/O8IEByqqWxNy3b5EPjMLoqyFH
4CcMsK4d+VQxJAhEZWNiaTNDsi0wfHa+1qPsn58TTrteyBYD3V5p2Uyl9kBE
gnjWJ0SEJZiso5AjF4UiP8AHZdmeihdSoCRMdSyhj0TG1eygGgWZ6b4aLXZh
rDK8f6WHVn0idXpyNHQ15nhqg9G3BttAzqZx1F2i5hHyhOALJKYd1B1P/3NT
pfuxZtmCqVRg0B0iiEntIFsiddA1vnsJ/1bafqZ5ei0xoeQ4PTbzHUCmzwOV
2SQNQJz1B4fwugQLVDJg2qdnhFhn7QMPsGsyaJoj74RQwWePzJYdymjtaRTZ
ZnnIq8vurrmu9t1KOF2GVvQhis2ZgCILR47pztpN+9qZBkXwG43vKXkWDcY/
u1FKGIiM3QgTnWLX0GKc5AMPrNnGXBMw4pqF2RcWPfcJ1z4LNdrBQ3eOPs9R
WoVmQV4PNS521wWsGPA/BVLmekA07/3ZevrcDY0X2aVXJ+MmY38Ru4Y4CwhR
cyJjmWemWfUgMNTZqK1pA5R06K8Ukp91k9IPQYaP+goqFyqe2gwsvdVPmhlL
C9n6TflFvyrcVNM4n2tGYFJiC1vqrqP5D8BICPp2ghANey92Y3fxmqNX3rS4
u078z1Iiyc4j6WT1awlyofmA50Qj94Pqad42Br7W7T7lGLRuUeIq9C6rmMm/
/q/FeedxH6TtgGzZSqCKVifnAwuzHuygzKfR4BW81guDBVwTSaOgDgV1gXDQ
btoiIDOL2f2HeotPLHMbpPSiuCHHLGISyWtGVowKrFyJ4bdftHyCqXGbMif6
OdDaPr9c0eUT5cdeomOS/P65GkO+KigdKt8InOLEWpMh2w4c3ZOOr33haeYn
aHR5rfoH8W5twG5WxvHrUuNRxONPl9nc5A64jEntPZYAuD2uHzsRz4c/5HHN
EA2c144kV7+P0E78HRU4YfXf8JUurytoefHVlk3Trj+gpVmz37rN5P3zzsiL
XXEx9M8i3KFrMAFMjEaXmO2D8VaydE9tB9wWQipRydhBlNkKESSf3R30Ip3h
0b9GzdVTsqz/7hYgELs/92VWmBcW/QkN+59kEET7BLXlpsWAC3yxG+8RM0mn
EYM0unRT7RjoL2lCbyW/s2ty5dbkxewVv04GKLRTpslZ5FBYtRZ8ce2o7NgM
MsfA8kN3eHCLYJK+VmTCoYC2JiTtiIVWULgjxt+FbiGFGV8Pvjqd0YcojNzY
WiCcClEumgQzb1BGf5L14voYJP1fNJ6JWjzLFJmVVvB6k+mcHoVdLMkfTlTV
aeEqKa+K4YZwXGNpbZ4YxLUSh1xjyjNjiO4DneVP9EQFem3exco9WlGDrj4C
OwSkxlll5rnvFvVESA3SGYx0vHCaC3W52QPiY/TAmQh3Roe2vaiOpipxofYG
N7vjX33J2CpKr9jsezj9qI7KlvK/I3vyiMh6LhFL1eOGeTFtm8L3Pms1/dEJ
El+6M+gTQPAdhgUxirK1OcdlssSnCpqrORJ+YFe0Fp+fwt2am8r3JhvY+jeU
zLcNP8Hlh06Qmc7rbzqK+B8/MdOVLC+Spi0oR4OBvikGlw+9wgP/SHssxXYr
vLuVGWB1B+D6918GjvqNEK2OzCXm/hOZHJvBUz1hClvyEBBB4fs/mF9FLOmL
Q3B1Nbn1lx+600xqhunYDdygEamLuZ9/0qr2W5duri/iuyEiReKB0my3J7wM
4qU+fYsEaEFk3w/96ITk5sUqS79aoBl222YR7KghsA+VtSkCkwAnuEFZ35RI
uMSwJVrsrL6EVCv0imz2Q7OqwjwMaFR4/kTC+85UP8IKQsZ0qK6YO4D21jLa
5Mv86tI3xk3a1dl4ZemfwSg0KStF6LaZ6I9Du2NKBTlW06izw/VYLpoeQdQ+
MmgzYXTPVh/qbSoJEqTNnogmCzljFSReKWa7dpif6HWKqdAFrRK7WU2qV42s
SveoZG8XGe0ntkXZBPqRo4TdV4BXP4Ri/zWlL8sy09JLL1q9fAWzOtXtkAmC
3ajUqXH6BRYcfcSMc0dE8sfKwyXimWhKUvpBnZUjBuKntf821vJFajEsZ81X
91NH4V0I0bkF6ghexbp8j8VmaV7vwWbCbS3NqeiDyZL0IbmQ9BWP52Zju75O
ukuqeUISKuiZ+W9QdEroZ1pjHh/Kreh/dnyHlAnWkSJZmAtMSeuGVZnHVOX6
qNt74kNtl8vst/A=

`pragma protect end_protected
