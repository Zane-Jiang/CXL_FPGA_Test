// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
jXKKVyZfmPkpdJHRtTnbq+hzaYfKiIiIHXQCG4aNNVGP9DakNWtgPWvf6rPCyJJs
M+qEwBW9SaiSqzx5qT5fEXoReCiEh98h9//U7aFZPfDvwaDeW5hEqS4AxZFCNd49
UKxvWElG7AZadUhwzMAwOe1iLFPP1f4H91ECY6pqxqQzJ6UKCLN64w==
//pragma protect end_key_block
//pragma protect digest_block
FABPjB4hv1LFmBZSc/6vs1vo2Lc=
//pragma protect end_digest_block
//pragma protect data_block
HcCuTFdfvOw1i8Gf39GxlCVUT4rH7RVfeDLmoQjYJpLPwRwBPoyio9TkSKYvK0AU
/sl8rStNZbAesdMppF8c+bq98hJd8Z4qhsmp+9lPFEXnIYR+bTSklqWd96dLMakk
iBV3w/a8NyXsaP4bsAuWeJPN0kdIMavX2qR2PeVBMZBOK/hqmZPORnylQfY8N+rO
dAKJ7QnmizKC3wymDAMnxz0GWFEo2oFMsK0OTiotoQ5M3Sxw4VFQ/XxFDK9MNETs
zVQi8IZtMktm6LovmRw9Y8bxFv5jlUN9/xZGJ0hiv/aBnPA3FKgeCq6IE60Q4Sdj
d0YSDvEMjiHeDabu2egJJCqrdeMupndSstOfcWyi2hYnUcfBHC9nHamm4KIZ1o4q
Y6mTcnFtENXWouHAY19OvTisbDB+C+bn5KHt9Is4BvsbCwa0wJZ2QgNrE8iplkfA
jLMPXiq00+QSgTdzV4jyc95LehkFaBKBvLsHGaGyxzqYR1GI82gYpOHzjt+7mVL8
wqkVZVj0hnglDGjtBJ2Jw32klH2h3W3ftrGURJY/9lvLI4TuEQ/BTIw2K1EjN4JT
iFYzKU6ShnruHSydpwLTGG++Yls+sEIFMrCLxigx2DT6xN3R7FdUgWNwG32a+Qh2
lhrvuz+IL3GOqFvpKCAeAELDUvQBLccO2vkfqs2l1Z7cgWjX/eGk4kOTncHjcW5Z
1KQD9QWs2pzYVREV1+KFY0xjrHmNJaJMaSjdNvGiDiKGrdVPtinXyD4Sz5RHHAMa
y62kSQ0+zWzlEGY7/0pFAvB657V2DPoq/rBZb5DPwGnPdbF/1/zgRdZpQ+sqFdMt
qyg5L+t4w9G+/chJ+gvSuGYXu34RKBSBX9svGCBOlQcdqqZoUoF3Hfk3GdyNi5Po
YUNQhGhZTYx9s4lMD2J5RMljweSt1sCnbyJKAiBs9GwdLgueO7ApulZOx4ik+I1e
mLUXlYObjJZEJeH23Jz43BBFatuSotKF8IyNYmqMV7/rlpS/MwSLnICx6p0u9+5y
vUkXxLIHQ/m3+DHfVqSJn1AMNRTdb2zePbU1IU9rTKHDijYgp0urxBYE+/rHLMU1
fyr1sEEyPhdhl+jYkHsoboIhlqBPOZ79Zuh4ckiP3C/RxXHZt4HiMYkv3QzmT6W/
5mX+OSiTfHwGgFWEjNRqDBz0lWZJYLppc6D+Lo0ISgygLToILi1QERZIj3XQDIyI
vLDXfdSasqlaF3SqiNbfgJTgq5JSsGzAGzuvIJHaJq2pLGDZAq94wGx7pOEv5CVR
F36wT0QjRCk3aU3gvMoN6bZHDMPNCLlmFqheoYBYiiG/0kgNccehkBfkwZU/kVrQ
axlOPBkPXJ22NLfr/jGTS53yjmhHruVm2MV0zONl26mUvdCGJi7xaC6O95aB7OTR
E01852Xd1/O7M8Fp+9ZnvfaK1Loga6ofACOA0Jj3g/TijAcn72k8jixYplqirN1W
6za26gjcS8K6QX1kdOIuaPdaY/FSjkkW2sIO/ux/dIvi0Uu9fGOL3KnnyJRcJase
Xhrv+OW6kTIdEkxpZ/f5/oLJ5Caeopc/0qE35eX4HTkczmt5cOJzEGxz3hg2ZOXO
tAale+ARFYC/7RYyok6zFdNbHzbEHPJj2pcEb5FWsE/bYpZFaWHCkfbD00BDXjr6
K2WfDOqQvumAMaAh/cUIBVLab0LyyCfE0F6tf9r9Pf2XlPJqPiB3WbY18vlc3dfh
1RppzCq3lFxcNUebL3zJEuenddGbGaPA4OeHCzGioEBWKoyj5BC58rzQK3DhcHY+
g0njR61T02nlk2hp/UozwD1y38qTNIRCiIWccVVf1ynQhwmy10U5cAMprKQlS30m
NBXa+gKAxWDyJHBCnJTIamJd3kJD3ITA+wxNVyqBRXgKjbsFO6mJWNPiy9tMMYvO
ENrLU0rTUjQeSkMq580zAb2NbrVheBDk2o00Nd3akm+eIpKVA/TLMRNpGH9ERu1j
pu0qfbXA5UZpfh1kTSu6m7mb1oIDlmB02aYpDgUTQoJnlk1nenkGa9dSGlKXN4Ds
79NeGaHQGaoqfGx701B/HdwrayTSaiGr1DVxnCmIoYXe6QJXpLJjzV0Kt9KxHl19
KQUG9TIRBk97vhodL3/Mt97TANqD+l1eI1HFt4g0x68au7ErgcnYfJ1Sn7m/DTYI
6WqMVhTrRMkz/Y9JqIMRN/oB9xrlUJQmuJLb4UxEhtUozanZDIlVZOchBO6fxXAw
AY1w2ZgQNI67E3yqqaG4jPrhxGpRyueblp79Bei/h+M5wZk3++e6N8510Po4qRwJ
/lfdWExaZ2lmhPJV4CgBSnU/AorqiZyeKYr/1B21nAg1HLsw1eGVgUg7CgBc106O
kwAMbXZfKPSfILsC32ADliKCSK3970GM4slAgjIkehKMQpP7F3KE+zw8LKdHjpf5
e84Q682//KaKweT8PRgL1FA8Bq3dVwwPWV13/6OZpU0axkV6LH7QDoYIang9f+Ti
+sZtL7tR7sIohaBdEs9SdykLp0w2KP9KoLma1+FPgxjHRDAfpWrL5uHBHZK+zMCw
MJusItMIVyeFe/Ffu19dJn+1Dpya7uu5Wlbd/p30tDA+yR5npjquHgEfgG71+dLV
iStlJZn0xJdNRa5AyRPCFdcnLJ8BluW3EdeFqhRR2Ri75ob/CBc+oYzlgjItyJeO
ST50dsKdbl0r/aUrWwGprGqSYicleo7AuQQA3jDjEn7d7sOSFVR0Zy/op5ds3E9n
xpMg2XCCEjuTSPc858fxSX3GFgGHO8OD5/y52vBkG/I1Tt7ZN+JKgVx+eq44ouRS
Vco8a73mEaZaLaQ+Goj6KHfshXs8T0bo35lytSysHklTXrp//Kj/MjLVekGH40aK
qKDtp8brjb1PR3kPONUdAgkmCB1OH7jGxgN5FJp40XPvIZI/A8P3KwByR1TCxUtr
eOBm26VMHiAl6pNYbNCUiqvJQwgFVIufQJDeLZgnWsCOO1yMFeHIV+7NhJz6tWdI
Cn9cMhqGC1jyxQuduod/NrUUAtHgGxw0Uh7KQoC3ITtdNKnjO5PUWa8xeJfC0nOe
qTud3RPCf3vSzoLe/+aXRIpCkU1ZfU36ux3Sb7oK9mGAzH5XJY74BDLMM+bI3PaX
BYseOFEBOuW9g1sFp7SHKMXTXj6u2/Mdwpe4oP7BRALebbejbFys/dFoPo/8JS/D
T77JAIMftj2d5uUzwClHEyV/lOJC/I2x9ooQcA353sOv8A/MGHlHXYIYC4JeJtcz
9uDCFaEhYl8JFsS5Tvsx7xpaVRzj0My9+W0NiFup3fX2fUBXo7ZkCCJYTq62U8Dy
kZiLDTPUN2W3EAxYH1saNH/q/cs9AgbFT3NzjleuGX5OgyqUdIBEaFEIeMCsyk5I
4bIFARIlQkxey2LeRzxTlHozBU0p76u0oOFZ5IyFfpPKr7YlZKb6wITWHArdQvra
oOhax6TMkW0xcQKc0tcuwSiHiy7t+dsH1b1j81SRQfZMR402Qni1yot9B54uDbGA
hGQZ5iRByTYFCR2/0hwcVEiI6tP3/cDuICz5ypvJLFPHFOUdkqwR5hHKIESUXM7F
77s2N5o/aBAujzbeDYxJFrvNsxylI8AWMAAzMqrWm8KtbXPyAtGoBuEG7DDzmkVQ
Azl4QY72kJp4/fOyHabPPios73NgfzoA0RRSD0N6o9yukmzIpbHr5+Fl9F6G4yJn
0Nvc7d8t2BUgbyDqT6vkGVJ5fCYmQRT5IDjD0hKoMoWcIdUUBtCnTJNPjEGWgr1n
mNSzRq25bwF4SiMRcN6moqD0UMxYydnOKDUw05/5WH3SmExzSmO68oySLTu5zXfw
dZDM3iiw7L+U4Bp4F7vT1Ks6NRxP4obKBpghVe44smZxt6vN/bgGyC9t3aS+KSqg
fGDZDriSsVIohLB3FyOM8/ZjZBYLq64KWM1VAgl72G+2LLKdMUc34H177FfnNi5U
7pAfJjfl4lMbvpVEKe21egwr4lzkm0oougRgYsM/pP1dr25S8h8etCB/VT0SmwDw
q83CeD/3bFf3559s5UV0ObcZLuAwifbdcgR8HuBUGzcmCtOu3J018BS13EfylO+g
J5mX5pZSHkAC7gpCeDbGAJXFdaj2buqReqnXUAh1gwriiRY/szEdLQK9zEA7iQDX
Zh91a+Yq+ZgpjuPANMRA1Rg5/aXsfZ6IeUAy/l5X7S7Ow/s6R2AICguyRBfUqfsX
TgFF4bB4i4f74JXVKwL5egOcuQ+nloZo141HiEcItg7NDf/7eeEtSQBD1zwztzWz
xP1CeTC//JZs7xHk6SAWqLmc05FTH48jLJxJE5d+fSc6vcQK48NiYsakkKbzj86+
ITBRFYUpWnVf5y9NEGgmXvsdMKnCoigXH5ylS6vhtDJXe/vlNb0dgAfzhv/k2vym
pXFg/44lWOtXs1C6XaoJEso9ybDp5AQ1e8EOefX112O6b4CFr68LjjW2C7q8cxmk
+bm5Fcw+iS74cuCKmuSNx80HBGQ2kYFBdBfph7hBCM12zmuZGG1cu2TZk1rtRvfS
xqwrIzfOxjAcR6xwbsq+GuZZrp2gM2IfsniCCX0nezPX4Vl+wPPv/gT+tnz10htX
xqbjw+0XeZjFFFZSIVtZF94ZQdNHUuLR9KBSTTkUhlUjNlq7oqAQPo0Z72C72xW7
D0bpcZXjRtjvmQYO8boywPpGF8VTtJWaxNMWMN5Dz4gYn8t8K/1JzIVwiw+ehXah
rHZr3mWHSsdcg2sEo9mfcbOUBrRc3tIp+q5E3KfD1yVZJLnmg8kkifhs5z1kW8sK
17ptyz+TXPdK/aeQY+E4HX68SxrwicJgdjvMBksuh+7ZO+zpwoTFaCIIFGxF+0Ua
dUg+llj7v36ajwOMQ3Gl7S/MiAyzx4yKQpvAUTXmuaZj8q+2xavZlnH+adMlbWSs
cHJqcfrHj0US1klDMs1Wfo8NANWhmbQeJC1v4D4rwJhNnKs8uhKknHI+CdkK/94p
bruSiSVIhCUqsVtgtzO5g9IXu/an7MPMMgJSukFmmXCDwT8oCFwkh7uUSMFT4dMp
Qe089tfPPp4Q3otNu0oAXQZg9L2Hr0tg3UZM4xd8SfbvlL84T8/oTxrGxsbipLtZ
llMjXi1Kq9Ih3LBFr2I/3YsznK/Cm/kvMyHYwUC3ozVPUp/YoZB36TjyaK1VqLod
0Uib29qwghwOWa/8jt2EHHcaO7N/+iffxNVq2Ko4zuxHplOYbNbA3Tl6J3ObsnQB
0jZ4Q/JZ2uRFewA7o8hDPJa3cMW03jT3/KoSX4Faj+iA97VDzDML7gDltVbUhiB4
CzXI5MTyUR0jx0nmwnwQT2FS7b/mRjK+FXxySCQ2TremqwoSN965dqaTOmFwH8GP
QGAYLQ1y+0yYxfv6HiHioPkAVx6SK3sb7jxjlwwwARx9oOr9PzTUq6fnx4PJRYqQ
t1rvTh1CwjVv5G0wQGcRbuufH4P0OfbQJuCeQfVQNin2VqJK/NjUxw5nl1itSX1v
SobgtxLTzCajHF15zu+Vcl/F0Pw9ivMm4QltqWgHx4ltXeBje3nSqwVU6tQKmDHV
1Vcq11gUdQaMSXupTLWFTX+ACM/NWH1ZkklRkB5FCpYfIEb68tHXx0/D3xiqrPow
xTY7QZag+7tWsfguZVA0QBR03CbwT4FpFzBcGQIPus0jNjil9eBuLEJ2A6MMKs3S
noAJuiZeNV3/dmM+QIhIe2gVZdPOD/V0/iMnmXInYZQYQyf/rJMOlGbeAeyQnesg
+dhU6W+h2WuAiKPfWp1JKflWrO4v3PdMeV5O4Hlk1GYSKqncJ7ueZxuPTij9hSB8
96yG2OiESoZztvE4yQFFCGG8qp4MH7yFKnSm/QfJWcirakQa3tgw3ST8bDluC76Y
XcH7Fl3fpLb5Q6m8ZBgT8SS+h5H7/OyTuEpS3fuzO084Es5l3FF1bZrZuTfS/Sj4
4M4+eEBrJ4byh8cLqY+dzw5d8l8AsCEx3i+ld/3ZVmnUnaXVYe9oKy/lA9viZLGL
4ELOWF7gQn4GAXmNx+31lhpIdIJoEOovSilJr8TRPJwSpHL/qrhYDtTSyrxPSvkF
ywTzE8fvR4Oe0BjPpbEs4mfofZo7KU17s1qLrm39WuundT8S6xTyt6ApeIZvTdRY
fjUOOwx8M4UIk0iNYQyVuDZSlvj8FO5JpHlrk5+10Cr+XwcCwzMYw+aYvbEuv0eW
wt45fYQsu5ugG0XOgX9keXZ7wlNs0Sd/l2+pipg+xubZ9r3I6xlctN/qC28xUg10
bfQGjMZA2vxm3dFP2aQ1wTvLIQow6L/tH9KfK+VXwIh1E6ATiA4D+8wUM7WZmu3y
4dTL/6oog4T0ohFZDo/bed76rm9jROtAfOHLaTlz+fta31Clsl70dXFjvq8fq7x8
6dIKWgwbexCsC67sc0qWzbJHYgf/GpsvsMwRQsKURqEpcxzwpBQvl4kV76hNL2D1
8vGICyDUDFe6YrQCDpJUOiWJuQ/t/gW92haxHZfanMmBAoXz+QYH7VqU3JXTSe/q
aQWAaoMgVepWBmnxj2rDfyn+hO2od1n0/BeSEkxgcfubjykIl8x8FHQPz8P9jw+f
mcmPIltaoMYaeVBCsjKQiJt8ERujebTAiHi/H33eEE7TPTDBp2EB7nYRUtcnjk91
g2FtIXNaDkSIzKmseIDqslurnLc6yiBc9zbwewDGZSKL1BpU3v/Lfg8esoATt2GP
jFyMf5O0py03rbLcp/BaKa2iw/w+dpqv0KkDNhahrwRTt9kMPjXDv74xqGD74WqC
1oXeSj7pTAKcg0nBoUr08v65i2AT30HIFpioQ+V6Y8+Xj3L4EyCm0VY0vxx0vDo7
5I6Bk+e8c/gaouhTaXUfrIs09Snreqdm4AWLb4SdsKhdx3M8vUAlNbFYax9NTQK/
13pEZGo4S8paH3wRokfx5z3fmyB+sBr3gOUGCG8wX+R2AFGWlO8eZxiX/WlR4Ear
m02tVLiLSVWldCT3l0uK5SohDwYtzj/Xd8fAqdIT46Ls/RH0wbaz7iwlVkmc20io
4RGhTSNNUu5vSp6FxuAezUjqJJF83494EcaTAK61y17mX/xhYCsYbERoujFT1UBi
PvECrx7sOFiKFCMSIJdxhIyhdQwRQR5WNAXcylkoPr9/K8mYuka/IcUZ/3wl1iIm
kqfjYDE6m9lJmM7HYFDoIvdRHRUyWqCg/e8olgw8GyaUsPe3UBbWTH8iz+qkcUgu
M50CbDcMSSo4b72y9hilPElC5KgFg0NqtYkJ117qupC2vj7yDn7oABgKSG7pAAaB
a8STjbPHMRQU7GfsFGEDAJBP5SJleopK2K6vCcl7bafM2SocLXE15Wwyjj9TsLim
sPNVMelF71Nc1dk+mKuje0E+J4KqPo5ATSXAY1b2ww1TQ1T6Snx/+788ogJJaNbQ
m973pvYcUGBI9wz3Fm1xCytu9yUoyOB7N161vHxXslzlg/xnHbKm7/1NAEqlzsoz
PgaSB1hDpVlzmAtDOqr6EsDv6NonUYdeBxp8qnemKeauWG4ARmXncSPBDQokWw8G
Q+mnsPqjNmbgkntbRqFhczjIfB7QO6Am/KW5wNt6bkD3l172OGT2SxaaFzhYQpz6
VdvgAzxpUsSoDiH0PlVIWX17rnnEcC6/QfffD16N86svFazZb4jmm06klZ8+KdwC
L/qQC94VFN9ds3ruKeoQG8uPMkqSj3vI+OCaesVKmxbmNS63NoXVoDkY+LjFztnT
ZWUcUJt16yiqUHDgfKuIO/GyySbjig4aCXbylSbcgk3piag2l+KQdl054GenioH1
AXeg6k7HAjDUJGEktpzLi6KEwWvgI3J24ZwauZ8SQKuM3MP96bgiAdGAl0JzuUAW
xC+ImsKYVADX9UP9jABzMOHsOh/uIMIw/FXa5Bi5/TMbD2XytTW584oWeyJuNk5A
sL58myUHrQsgrlCVF2NchVu0B9a7IkupAdDDXhCuNq6YPh9mJDozBzdwIoEPKbjJ
Hc5eDjW8Z3piJL6X1F8uo9Ba9er2aTfq4NMJmGLM808vVu7x4XLrJD0eQrSk42Ce
eAq26tGwzJlpzILBR0oW+Wfx5ejdBPXC/LJ0Z7A8N0r3/0tMujP5CaAtqgzCliJY
BlAibJOb1N7n+XD8AWC72BkKCBhA7Rfcw10hRizdHEcx1jWOWbFZ0JNXO7wbwzEp
0JYxRJsgTXGJI12PeaTfOQ==
//pragma protect end_data_block
//pragma protect digest_block
IzK8m7V0J3zZvqBmIClGJp5zSFg=
//pragma protect end_digest_block
//pragma protect end_protected
