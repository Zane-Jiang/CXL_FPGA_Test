// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
jETY11Buyerdyk2TdEzndrWQHbPQ+tdRpd7SOmIEyyDKL0ykKJxkdzpzCblzLQTAxrZ8mVexIpI2
sitaVeFTiFyPUfPQCKfazBizs1I6Og9kb9QIDT0QClcXdTNGZ1chinfWxlkZV54zrA1AIhJIBQB6
apgnfywPHrdamgfwguRSYDPiSEtJk+anpu0yfAbch9AIpcHPwzrKW/v+gr8UUQkD06yL8EnSETEV
IVrAucnu56x9U2vRpQit08hGEoo5rs7lkbsVtX7Q6QWkT0ko7k6gg6nLM7YdHR6Dxgm8bHhgjZG9
GwiKmFfXKk70Hb3aOum5YRxNSOk6jxbZ4ZHePQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8464)
pP0mvXFow2r6AjRxYjkxe1kHvKuRuPHQyG5GTdCbYwwhV9hDi/3bqrt8jdETtHenqCopd10ENykO
cD9l566OQ9J7pe3UJg6j8O/Ii1t7jWn5RqePIRppPqssbrAuxAgdWz6ihhiZ8i7PXMJYycVhSOqq
II2xn8PKtpFjhL1/RB748Y2yfBiGtuPqwjNKRxKitgcBtWUd/WqgM5TOA5v0HuP6T7w7oQV6sZqc
XU92NoQNw4YlSppz54Ies+Kw0hGrFtOM7ZjBjPXnq4WM1iEi+f1vqJWr+qEGKBZvEGoZv1Lz+hLS
gNNE549S4SjXb0lAerHUaMmP3eAWqkvwSO5/q7NfigGZAGLTMOt1VONWHKB07w3myoevxD/MpKiN
S3WFI7w2PJol5CuWdkiDl4Jd7UtSg57kFajAcbK8Zpu/4GpXuG2CbiWxbafvAJfReizbXoh9aYMX
LOhSSlqWnWBcL0dJrRjHLoP3nueb5SSWR1lHumDO2rfPTWwSXKHJr8Mrw4pgovkGXpsT/d3QYlqm
qAxbFeqCNyWeH+1MWLtZKby39Hw0AeYW73XGFua1kGfO3NiQrPUMbpHIiIJW9HGnbIHk6y7vxqxQ
ZyirNXMEKw7xnF5vplq3AD5+3CVzH7XgoiNVyBnO5oXqMzWAg+N6477ZWLFIhJR6wQ6LkG1hFTnp
B/ErdiJJJpemjtp/Ms15MmUU1V0PNO+kxZLbzKC3d6V9a/vfhmXnFEwyxcCP4pRlVi04RG8NqQvl
I6Xnx151NsHxlV7y/C+EolnHG5D2sovF8hrOfNpfSiFOfePvki1whg56W+CpFKInsfe4SFodpheq
GVcoQieKDQakHh5hAtKAuavb4TVm3zGUInwi1B1MAEEkDE/GORD3lAzBTar4ExuHENIp4og2ncWL
6ZBZ2y6IwgCc8mIZ2NFkc4jYaa3RE9vFNnH6BH/1MEe/SSScUd+TfVC2xz/F7I3JAsCIStM/Rpwl
9v7UgrBsh1KgRN6gP7Iavzy/BSboDLEi7Rw2tUDsceq5I4dLvF8tRlbZLQMVhNFb8EB3siK6L6cw
ym6gvnaUihQM9t7pqnONEqC1kx1HHcdsSO56vpm8SbD8k7Rfun8P/aKoNEU3GMpd/ms+I83wAEtL
ykF82ZOHxqoQokLFiGHj505jiAXbJz91cfHEcKkMl8GzejUE4DLWZPiB77pTZC36ZOL5SaUNouw2
YoSfAxu+GmAheXRj1Ot/BLYDNF5W1B22AIo6mxnA7fTJfYKrokw2OrTMsNuvc/R+2TtdIpMk5DYW
SG9kUAje4oHdUb+uBc5aNdjIcVNndw+J9n9Nhv1QaeAqSbUVUlnETYrKB9iexc2eqtDu4ATzxJCD
VYpRlOPJ9CRHyqa7p+QqXxQ9dOpcipcCydpKm3Km+bIs9ef4vdLnvAJJYSUAUF3uqHaNQeaFgRZt
Whi1iOs9Bf5SLigzccowiLAgkrFte5YAZCg3h8xxPqp2W1/xPST6YYKbEgN733y1aEDFX0S067rV
L5UA6tU+z/FCGlfG6tUWO5TuyiveAiqqubpAONdDppf/jVe/Fc1TXfAqXRc468ieWBwUIJRmWA9E
QVHTooIZRQDlhvVbSkEt7AtXT2nuHSER6a2tKYDF+NLdwsfF5T72TkWTGEpWMRO2sZcQbzLYYhIO
w7YIGmspVJXZg6ESfQf64c8vUPByINW1cDv8eTb1qhdKxiFzBjj77tDrR6qxO0dZ1l1JssuppOKs
+5/VtoiIo9j3/58Zgj5Gh5+6fjYG9LWu5WTAgWrHx8fvE8LUxNbGIRxzEP6xEMCEl/nCT5XzouxY
2MAQNoGZle38k9jtWuvUCqq7KlVyJ3pmRztoOuwLHFLqdwO81xHDpo4KWWuwPy45QBOa9dzPpogW
O0NZw5gMCiRFp/g5YAPMwJ1P08apeBPdL1vlWrY+FpiMCPay7izTuHUW5PUkD+7yrn/LvuLTZy6U
h97B/WlVCLSVG7h3CAKDJPvRaCAu/l2uLbuYBDrfx5ynLaMMURoE5IllatElyT4KEQ1Ezum7ryFG
bcxyNVYcgqd+urAo0U559vPWqQbKI4vLg3z52f20t0h1dMrRcP3I+v1AnV6Obk8SV1qqeuTetTTJ
KRw6BgFvYfbL5+TSyR93S+BtIUC8Z1xnIiSC9vgH/hFTcXBPKvLLMVchVryKMfqT/LkIsLpO4kps
w26jlbfZq2cvEVxJ/rfiUwCSry3Oprnw1MIEDR9ukti7j7iwg7LRcytriMXvQXasSYlj1+6XXU7v
JScmJYdlsGYBVikZXaXtE5QlIySBTjaX5mbzGaHvZc7GFwKsSUV5ALz/afRJMVHd+KaTBhB9eMwn
Y2zSVNalL78cZKzY1yOnqatomMHMAiCmFjHGysrAG6twEFRDaCq0/pvy0jRACtveiP2+jfyNrEDb
7+j+q7fG7jenTLnLM8L+OC0WBf9aXx8LB/9jnIxUftLaU6yj2FWStRKuCun0+WZNGKIVGf4qiKkq
MooMvT3vHLOZhWT7v1puOcSSjWMJtSQRDawQ7FztzxLU4qKHKwdVX76zCssF8ZXJxJ1DfaWGfsgp
81ciPezjLI7o228RXNV60l3Ybou9qYHyOu56CnqwoAUm7ngvyqJOsc1iqBFlf7szIwiANms1YGD4
s07Kt8fiDr1IorM6V9mQUC1hbEkGuV9genOCvyP1CzjgUSGiL5n3+mDbKAw2ywI0snMBlS6+RcJo
9Kwh0HBYaM12NaT5/6DzdJSu9/WNvzWr4j2e2XuiFlWtdb4sxQ+e3BckID3XNEZhLHt8E/0arrGE
K53PcyNRbpx4ukyjfoIoFPd56GyPT40b0GuJGebmynPdd7uHFyD8HzTkpJdxgPccDOGns0iYlHO5
IOJx5qzddiEfB/4tFGzVTlMCB6XTPIAfcO3cW5BYhrcJ0eBrXDXeRYABgG+cVvYL5MF8qyGDl4Qj
bdCqBVoBdiymdqpRabjyNb90vPB3goJiyaVVwlLYszpfCgIQWwfu9I86EGjCSQVX4H7WpEqhDNug
jgL6zvxBo0EbknO/FWLjNxTwxDt4m+86SeYm8zWcRPKwLGQUzoyBCGXXk51ALbIqV913Tl6fRRf+
mmTp7BlbWoONCrogPzVk+ezOrIJZxgKALFMThAPE/g0HVV29kGuFmMbKCXIiizXNEkGp+G1DSjHa
UbdBNNIdoRF5Ou4J0eoxg5iJ+p4vxWkQ11Kwu9zR1P4tziOc7TAzaFBUvli27Vo2+twfSMlVk6wY
x7oi87ggz+HYLd6ZPk3sRgoGxJxLr079ukAQtVS1Be6udjPRoHVqQKxHtyTwNphdXb7yLdI/jWST
liD5zEteLPJzoUXHCJxSANdi+PoJDCJLtDDnDSfyhupgefRBt6m701g024+H9wM79Qn6mJIH6Ber
AhLt9xazVb2kgceJ28SwpfPhol2lmmkqtekdtrFR3AXMsUxoRgoBoZwUKs8AoRG+XLn2FifandUP
mivphAyiytN7XzzU6yiKfLJUJxA8zT4O4bBuoojdZt9vEZ6gJeAXjwU12tCGGvAMUZV1I6fj4l+7
To5eZ6eqkexg5GywmMtuEj15Fi+3fFRkXVGoBEANU5sTZbTl9KhZLxG4RdDSn+m9CjkCLC9yVPZ5
3yithTwasB8fLLh+RuU1MbxRbFyoDxASPFcgipC7pOVg91QGJ+NBBAQC3jV5bznbtibNTZMJ8YBZ
BOMKVut2YjrBrahCXV/Juqu6Mchbz6F/MdBS0fzwmDpLZgeSKjvjdynBumuinpD2vOHX83zjNVga
79iOwTbm/Daysvgl8GFOVL2Q0dIc8Ut22mZqMd9IsTsBZdyElDzwcLHrS+hqBBkIMIh4Z3tORwdp
+JvsQx/oTqoi28bMpiQc2vEJnWbKGWCszS4Mu/zZBWT+F1GpFULTgrvAn8oqUiwTVbIRvxFKL4wv
flNQNXeRB+fciAzzyBDOTcbKhr/IbVsDkxOh+l1t9cn3Izrzd+ElMYTGHzKofFKYeknoPPfgFee0
TuxWT6lRQDTk+FgO6e9JLFh0i+sNCxsHZApcxqHZmIPUe4gcBcwkgguAA0m0DRYu7+QaF/tK6wdl
Vtdkr9H5O4eoJP1okG5wcD4clCAWYqOaqBwGaQhaRRM9L1BDarLfE2/nmgcgkSs1M2ByjPEJd9lk
jctiSZPa0/AtZD4ChhMeEnZ3/RgyJpDSDR2EHSvYi2ixmF560hZehaxT7vIsonlxsl7KD7Suc12X
bXehQCA8EiNw3ecCE5Z1+4r2I7WG4DjlAFghgq2meo+lfBz3Ekji3Pd9COnAfI07OHV+krKDtuPv
wBNOjre8JGG++5FsfzyO+fHvIfMrj3mO/6pnLhYNb7AMj7ko/eIrxt3F96JZorgqFazzEJQ1LV86
G/Fb4PAXN7ZCrtBAcoTX02ac5pqBW7fHSclZHTRF86H6fzjNgAdfFtZzkcBUckfeU5ZLx61iOMDd
E2b4hWPJ108yG7QwQDsby8XTTWQC2fOj2CqWhZ8NikualeV372Uw8sFhOvEK/TWSMh/UAppXNs67
01X2QSKlMgdTWliS6W1p/pDHzKnXc1dP/me3nYxYoemWoTWwCrBBR+5l4BJpBFqzfMIw7oSWiiJX
l68hYsn/8+fYUrVHFjGbks2hellY8Pwn2xrw5ztviIInbhxwOxXq/EBhZI+LTAjZz9F2VAizk4ik
l4EO03obj4hbtVXyG23r3O0anQ5B+ANtydB9ejM7HuJtNlUtShOLqDeZZSvbL3GAfhzZvkUIJjcr
C+kz3gyQopGRxBOKajRwnNUFusCzuFaKdkWJQCBaQXLUbrRjt4eM2rQWQMrctWfmXKKKdyNo1idp
crUlbyIF9gskf9ZB9IB0xgeS1SbrI/yKJWvn9PsphSFqjJRrzlYteQRGnmmCShJDGdKVpEX2KKFq
sSchzfLsojSqBEjb7mciKWtLn0u101Ssf7sKehgHXaTkeFMozKPAawl3VfEvs9mo15ayndqe8wYP
FfGdH2mxq4Ea5/ENhHWn4hLV0DqJl9mB4+7CnLb2LfxS5R/kZXHOpnNK+4ZdLPIkVx0QS4NTej5x
lAsF/9B2DdeAVN0mICiJI0+fr5jZ8cs5cKR5Sn5Sj6q1u7xhFglS9Ghu1pvafmhkb7JWylvOK5Ge
XLyVbONe1eSfcAVQuFArSeGzby7ten8HcIiS5SLixsAxDhYkEQlOyLDpLa5jC5r+h6XdmX6JYsJz
Cv1lP8JoQtEgKKDUJd+nzRao7ScLAUpJo42/Iz9wKFZOu6ba/VncFQ1D1JhFBsLy44vcO2BHDK2u
womL/ftb7EisBPCVbIVzZ9zZFVxkBILKYZVTF1/DfTwnbTFsOe9YzBdU09GzWgSkAN1iW4HF3lt0
qCW+g+/h5PSr//yLC9pwhkcRWP0bnXazIi94dbkXPFDBphebTXhFwrIjGBv4HxX3Pd6In+j0Egbd
SnTYEsGRRdXORpOyio7RxHesNJ5dkaqHSHhm9x6Gy/KpEEEHvCSiVO3a8XbAdIEXpRBQUipxOB/E
ZkbRbSd6kzfNd3+EKMgV5vsblINhCyla8U9DHUIXQ/VHBJ6wOB6l8zWH6wVmyHOGP1d09mdpu8CG
IjE0XtVP6gT7qKHRq87HPHO/W4DX1KsbCP3SmwSYLj12KvUp8V0l3IhYzRIoxEsbL+oQGgO5DHhD
ciR9qEBFT8X/PcOK72Nig6/J8BN9WAcSnZ+dDfOwEkfshyNIaHTjTdohhCGNvZPl/2Q/kPipGoaP
SK9ZB+xFBKUuBlaYa5oNMVhwt/L5ymfGa9okGQd5RLwO0W1Qu2vtkwu6CzAaJPgvejCf4JRwhnjn
G0cF1eaF6NedxsheywF8WKGtssecCqXQWJ2/++3XETbyXVuVf8bGPjWBcopGXzJOeN7Un9LqRyp1
W0HCXYDkrk8IYqtWyyWLgRpv0dNTRELr47c4xFWNlN30dboFYSa0qEzyLgrodFmbAE+vS2ehLRPf
J57GZyCJXkLBOhfHNDG7xukJWUy3eOPYefAwD3ZazWS/NcQMSmO/kKHvI6BBkprWsWm/qDyAxHwk
r7xSnaYSUVIS9/0RO+cMoX6qIfAPnzG+461rYQhdFbDCws7W3hrM8WEvB44t6vJ/Uh/g2IP3cNZh
fTl8UGiDHTG0jrs5yuzQmkUBUIqUd/i2TrkoDFbhEV4ryxDJaQHYA6JIyG+F7T7j99FvKLZXZQSO
6i5u0pI6oQhM6ri3SAk7t9XZtOdEXzcmdH9AAi9F/cz7B0Hnp4LwG2TDQaqnGDH4dBcVALOyMdFM
Cs2tblixLmc/cCobxi/WYJ46Peu2S9C5KVaBmAUb/00smg8BR/GYQxsWg6yF7iUirvnAsepOvdJB
2sP6tPSIdNDADT0fhVnO5XLF4RL2LfussLIFK0r1D7EDOoaHff0JlHEmRZNtIFiOXizO7iK7cbcv
mv2gr1drjNBG/KFeMiLU3vTiNQOYB22IppDswKSWOf6ohiZM0Y56SX+egYhaNdhQYeG7ItjW47T9
vOaodDRGWGbMw9OkEMlwB0jgK/HafyZIfoQHiLV8PhxT2WrK2DdtwB97cDx0amQsbpIwkojT+vFe
SNl3it+STrL6aeOnXWLS9g5JgqqAyZDDPczQPn2P9yE73ISGTcBxgLzefYQauGq8B5kae/vgqjfw
XB+gkj3LBOP+7+lFqrOc7Tq3Djns0WOfpkedQbJJ67ZzvPZPKEYbxOYZSXs4a012yZzVOTbsWh2B
BFgiKMWWCutBvFRj3YHShNnJphI7Dwygst8LedXcAPRsRjRWCiRIVTD05iMwzZ/pkk5Vhi/ycnAz
NcNzhzkfVg5WSOcjPjNTAmOyw59MVX8Sl3bm+y1bryes+YW5rIX8qOiPgPV8hJXK/hU5UHGRBICV
A7XA8d0VKsRkr7vCunOyqDbeiwdqZwXKc0JHy0PQl9mYUDn7b4q6OLTdhVMvX3xrdSm9y+yvpvBL
C/yvXLsh7JnEY1if9hFP7v8r93suCSX6c4zuIRw2tCdHAoxcjhHR1ItLUTunb7AOPCr+HNeLBdaG
yLr64Oi8IoeiAUCtpVCif1rO+CgbaBp2IGjs4cZUKQSBaLXMFcL85d/mZP2Rd50IqUT0Pg9rUkW8
bKKLamxgX+MB5w/QTKVF/A1bZQuxPV93bTmlSdC6tRr3tLRZao2rAHTivt3QgxDO0ngu6iBDfTLD
I4/db2qgLPPPPJBhw6DaGbd6WJc9l7oWHKpWhINg82hnYyKbY8ySmj32GAdD94bV+/PAbHRzMisd
az1keKG2/dyii9a2T6G/LgupAOpW3q8noD2+Ec74JJQth1+9ZepiFZZD17CUv2ZzcNXl+5GFzhTv
gZ9GAf1CXQtPwXYjg69kQxpgpB+uun4/QDGQWrWYhH4SLSNk79Vgqbw41FTpWfAuS2eGl0LwStAn
OwRxZavcFeptfM4cAdJBaH6G7uIyVIlCu5/3dW1rJiX1UVbFdWpnVn3nvswmz9K7pnHQHgQuZBgv
t2/TPm1tabZsYx32xPi+o0fbqDNlzx0SY109gtELuC5KQcucdHZFt80rNtz4zKnSYd5GYZ/4yCgj
WW2e6xORYVQ4ugINrFQAX2h8xzuA6gCom3BIn3MDdnUAqCgtGPO7rgAqrJrrnguvnKaRDVLuoLI7
yC9PWFIx2JedU5KGtXdVhVPMRRC5bU83zrwJid7dfJCJJ1mHD84BmqbS3kSv3tW3wL8F3MJAc7N5
fMgPwY61Y+VqiTQ/cb4bb3hUOHYEkRT57lW82EgUggwapPtVKSOp+ZmUUX84bIWuwtKvO8nWQ0qI
YD2KZcQvu847AOyK9kYmMKueoNjITEetpDBSMAL5iYboF31/PMFcjNLgfZl3k4ECm0shazw5gsfF
YD/t8GUN0qnuIZIx/DdN38Y6w0XnfrBSVqEXZw2HWFf9zq/EAQIeuN7BUPg6syew47onVOXzjrRo
eP768LsRU1CSqONt/taRSAhjHux+zL0SMKwqjTC0+Hwz5lQrrmYL3PiMEas54N5sMckvVdggztci
JJ/tQhknrbO/gBlMnjbdB0WuZWe2KW0MWNetkZFG4Hr5mtQQ8NDVn/jxYXots9NRKt3dvcyES+1u
GWr7quzwhAF4O8JvQLRICePeRLOmCqis5Fgd9lgg6c/jJzvYw8KD982aqdwu/ZaU5tysbWAgIFvH
MTEu+zeKdO9IrEWyHPKAXgkI3+XjaRMrXcMUeeMMoGJ9Z1+lx80AA0AYldMU/mWBbCoQufOw/rTQ
kkn5VHwJW+Y60SmpIxl73nARolgANVfWk6UjEwfpbZQe3caGs6dClnlWI1NupOSLlZfsBteqwmPM
jJenl2G67H2HEgE60xu6ow2Dy9OiXsHa8uu7fI79UWezp18so+B5zYB1wQGc6SeAcnKithgQqOvH
7XPiDWcKz6Y/hALXwolCYSk7U2v5yJQgPbF5kbx/HCNmY5pin+fA+nQX4ccRtdKfuqKNSJT55LB/
hPB5oanyWXND43Vqb7+yIm5i74jlkqgiYELyYoV0GsLSNl7nULL/Y9Jc7zo/j5ikjZrLNJh51/4X
1rL95h34LOXD9gOCSJTKXoAz+wqkIiZAYftTqbPx//phsEZQGeebkj5rLEyjFmxPHptD22BSCO6A
l4IF8L9GFjkZdXmXxQzp4qNkUjpGhAKrG+LC6VDmC3QGl//x/r68wMf6QLmU8qbVaWCJ62sKxsvC
ozonCt4H1WNDBfL8zJirLGcxOjK16/ytFDcC6K0vX+hJ9GUXKOXXGfQHyvhhdeOKO1RE068PlbOi
oX1m5Tb3Ba9sMxMxHvmUQM6O05gu7WoQ5+XiXDmi7WC4q9K6MUOkgHJKkjVvi+AqvTLTd1O7UdEB
ZMMDE28/OV36gFQMFfQz+JkM+EbvyBhdmZYON5LMMlg0zswWT1pU9bGfndq2sv4aS2hbL501Xt7C
xQriP2Gir0B/C+m0gFSVidlhKvEJ0pjJKQmuHkwglE+Hj/phivU6eqO1dDwYaeoagAEHa2x3quWb
vUG8bjmuMYShBiKpNSiJDPFexYbeXot4X/rt6wSRkbzAS9v8zjGTZTunvxiKuZAiIRrSnOVGfgLr
BBqScrairLZBOFSZPBAKPX/onwu+i2gvMLsPc6Kd/f+sjXmvAXiUdOt2mCIri2TR6SSphAcPAMjt
z3kBiHOlAh5Z1SMxANNrbEoeMvLxeRh5qr3PJah0rQ6RTcZ7hsRNbEH9cx7UfSvsKJTKbZfQbVuj
m3FMBkF8P6/pUvOibMM9JYxagZOb4wvPv/WhX+nr6stapCcbtFdWrRb8HvXKPJOz7UCL/UiMTVom
KBH/4W9WgkoOV38KqmmE7Lz+H7bjQyot1HWtLyKYF0wkzF9c4Dk/sWIkYxd8+BGfIhhrVYRH+zeH
12HH0D6pJHEojwW3u1WpcvoDpWHGKjS+bcsehJlpXXgpARUXF3nHPEuFdqY/4xjoTfHHyQLMlU46
SqTABpPdwZDtqqYTznI30f5VF8dwvK2q4UODR09Ib8yLAAgv1OC4XLpzq4e9mvRMM+YAQXGovrqh
yH0BvOkBFAMa+oTJMfo+T9zgeHh4U0cqgU3vZrHj+uYdQ8PlbDlU/SV69afWsxb7YHzbnSCzQmN9
SxXCkBxGUe155mP5ZIjOIORwMih+y0Nn56vOKGB4GcZLXaHU9QU6w7TbrjEzDbiU/LycR3yiT5i/
YrBfCA9UKgLHXMW07B5WRDNVPb3jjQvtgIhpOJFvoa137AywnvtmMXIxYQ5vVLIeLsGA8JiyyjXV
pTNXzXD7/3qu+0v1vbKwmaIMed+2qeRHUF9kn+hncC6Elx0yQjfkAKT8HHktShr8ShVZTiyX1THJ
sOpfG43rOXEvmXBlLbKeQMLdR8l2R8xAcTPR+rcs46PFEAzZ67r6ALoQJY7/TvNfWJ+Wqg2iLbCR
bZ9hwMzGzOQELoeZnRLhCyzEQznOuOMVJHP3hghz+6LBGeIR2jiHlQcbCOMK9NATjcjaZGD6YgF5
8OA5dyBixe/ZkoMS0l7Wi6UfKlEzHyx2z1meJqFcwzb2fu72pnSMvp29Z/DKBg6Yg55YECBASKeG
buPNlBqHOR8WOjxHTU3QC8TkZks+a6rdvItcmMFrM91MrSrxupjRgGkPvprde83FYiyXFZb1PRtF
iY/Xfwl2xmWnpJ/q1K1e754YLUokWSq5NYKrFdYw32DWZVtKKCCOX35A4+WbGhbe79D5IevPy4NV
9DaoPpyNub3jW4gvw44U92+vJmsZLwvdkAGjrim/M7xfn+Mkkrc+bAxnJYCQ5Zso/67XkV2Ywz3d
2M86LIZOkw6rBUnOqHOmt7G6UNWH+OEOYuzUmn3fZefeCMDbcc2zmgJ5Ycg3ylfm+O4Y1QVY3zxB
QTv9E7+Prr5aYoUfk/Q054pVBwV1+SOt8C9jnacPcVPIlpYyzRSFC3TGUu1RztdXRWmBB25r8irL
drTpgWEdj9p6mcxJwI2s+rmisQ1DBgaqj/V44LMQ1TvqlN33R2v9ySLXwENBjsMpcpO1Nkfwt75y
iuIiNG5DBTCZeyNEDOXTtdzdsTyrETOA8N0n8qHjPdsVe2bmiYN1pUGC9+KqtrRxf9V1/Q5YSDLm
lg2izv/KYNIAumqSjnOpWaeTCMyINWfhIJBSnisigYQcixCcxTO2dYP/pRgLu8fZZ1ZhfNrtcip0
yJQhjtb4IhV5FEZokrDv9xVTFwKNNIr70bi06fc1MkWqMvArtk5+ackwpl/oOAPD1LYkNqCBU6XK
5wRTGvXe8xg6SGljfYHrWNInArEP/bcPBio6ACgKu4Yi72wWdVO0VmfR88ryU0LJTpUkWJSkZePu
k7JCaohwgRPXTg9awaZ8rR6uthSowdZWuCk80tyy+nFiIQDmfnjw3xQPvvMTuDXEjhXQR/HbKEbw
HMdzK79tDyyNrjLKJXYTZZUFfOHzlz4Cj37Jxk+NtDVtvXzfelmMSAKZJYsuW2wKKJSlHgruVsDI
xCh8dHKdtsanH4E7ameltZyr26psy8FpwkauY2CyMvkl63Oj7TQegmC+1bPLuuioByXRYsy0iGq/
luM9XzS/Tn9hWX8nC3PpdUbL5RuI6G0+Kou2CzYMHMo7yQ/EB22LvB1IWmZE89RR6STmctuhHDBm
r4n+JhcWQpALpXrG7JSqBs2tt60n8O5/0hmwmePpfVG4lIQDtiURwJMds5x1BM0FOBK4gpWgu36t
ToAuCrqIyBY/C+LozYh8TrTKLTsvhp0Whrn3Cg==
`pragma protect end_protected
