`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
DxpIj5aFIBlFLTBJT5EcTlKABA3q60l3t6OpeXN9C5bFTwtTO5rj226qx1yxBJvw
0g2fjWMKpnfBPNTXx2lRCi7XDwpNbnSVTSJTRQNDeELUGrn72/i9FgpcOmGfuRMX
9WvE28Hbrcwkn4blSO+83wwxAy+34A12lPKZW4wCCFM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8624), data_block
fTy9zNdXijiw5xI+m1NAxgK4YPklGfFN8usLRuECvnAqQX30h1twB0Y5HiSIC1Rt
iia/BmfvwkwAu+FHuxJTanz6oDsgymxNQsat64uf5DahZxZXGfPFBiOz9Smc9CJC
7HBl81vtb/R959zdmhF/DWSB7R+I3jiJBOBEyYYrTFYZ3UHRqTyvN5y0tDPUIS68
UGlEZ3EKV1fIk323s15AwVXRgC0IZJ97HSHXurScWOWWImRfPgAB22s1Qh8hU/yz
Z24syY7rW5ExGw78ogtJp5YEQyPO8nEsyTJXmJyTnleA+dyPLXVTg/ShpfGchCTw
t0u3v91Y1/zHlrwSI2IZvRn42wSsXM4ZbZ9mHcissyN2rFkMpzxuGcbXjSoKSQwL
l9vzFN5mC0dp+Gar70Y1yAgCSyhjcOqZpYRwUamFAsOZYcSje4qffpRQM4p3WgWL
Qgv8TurrklPjy9jJ5H8UrtM21pMcQctQF2wnICYtEcAEmKknf4pIBmjqdGTY89dQ
xZNPHAshG/GpeCknWCfTcHbc8N0h/Emy+l75l3nyJxnbG/LPXnjy9XwMUMDOoHJp
pYHmjPexgXhcz5A41VWF42WO4jRtx7BskRBjDZuLi/VZmkCP0B35xsouCtHSKgCQ
qbk2hH7AdIOxNH0AZZL8yd5vJpiAUtZA2aINHTuyRbZ00URxhvPfHrEz+V6Hs3sW
jGXewMmb6I3qud9EYNEIxzm4ZK739INb+vzBnvtvKWs/Yzhc9dpMcw1mti1C3H7L
KKHcDkEPibfmEmADXoH9GQq42SUrL5diLAsUAbCgCYQpyakIP+1kZA/3K+tGsUI8
SzwSod/PT7mEbdR4OxcOhb9YFEHCvxGXN41jwx7+Nwv3DNPdAY/cIBimWnIVFZPB
QGfetvnDT+McjqGppjN4Jqaz3au/bZaesDBmb+pvOJeiNkY2Oy2+GylQiRE7Htg1
aUlW9K1rHtLFOfw7lGA2MnLLmTh6fycbqQfVUNhUcvpDbsrTZDXPJXLyMJoIT9Tk
o79Erb3tCVi4/JL/GqfH6NWnAawL6BTWHxbvJ3y91mh7MXs5j3pzYEuF3I2wVvUs
E/DnKwtY/KkaGkdNQ2OpadbxDKQtWER1fD/Vnj9V1QkqHoH6hhzlrwwvgM93hEsd
e5nVAWK7z7OtOZqQxtVCBZMbQFXIfS9bRQ6ugxTKQ6wLAlP5gharmS43j2OyQpqX
GQOWf4cZekIa7cpfN5lAhstcMAfOh+BckWgY+XZd5tnEgnbqLCiOfkUOs2DNN+4M
5w4y0jxlTDa4mBKrNxtYJ4eK+ZZJjlgjwtMJoiqh2pTYbJn10Tn9HCjriDpHs/kf
WF0eM4N0g9a2c2uKaOuz3T92WILkSRATQ8qAaISIBDslTe8fT4rCBBEspjoft/bD
9VQ9HcCZFJh91tcnDPoqvkJ+xmNuPi+ya5HXh8JoN0/8cWcUABqu0DLh09BhoC+y
eD4NKw8zKgr3p2vZ0MutGk51Zl+8JLr0ABMqeiaFyYU06pVSNAmagvH5pJuib/qh
Va+tIxSxP9OuxMpKXbmQgcNL9JZw+tpYJjyPlW0zmyzfBNrUNsBDrd8XFmCc6OQa
v+clukGGOd5BxRJNbWk/iTN8dXlziBm3MkZt3dLEAnoeYIGTd7cY5SL6jwyZsxks
+aDL+xox4QQUMnYdaLhk95eutG7+b8uGvTPRw4SMEk+QaAewiPt+uoez0kN+7VEu
ArxQ7kcM2WkIoTOHRCNG0jsufQhjcTind4t75ltcpAT8FBUzeJyQNsVfbTafy2I8
uHrWkU9bJqP5ahVEyQ10Y+DxvAkuR6AFfHU4APUqLHdka/IvAHZ3Lylzf2ZM391q
GFNSk7+Su3tq3RX7nPAypS+NS6V0EEbnArx69Qhd8LRtKyInSPGnhgc77D8E0DAf
2haMIzaraTLoPaW8hB5xTGACm8KIS3KEThcIJy5A7AY8jMsObTB2S0ayfwOzbRPK
7ad/cCyWrm/6qbvwto7mxSdYq4zYkDUkzKPvlUSuH5uq1A71eEdl+IQrT2uE5GLA
iP8PobXBwWvQT8BPAWVXWTRytVqC+uyIegi0N0JOYnrCpDC5DaLv9MutYDN78PbF
513pawwFCTo+YfKcqqD33u8uaSvfV8DkhlHMBMC9C1+0Z2/7Of8BV0QSYiq1n05G
QdwcqD6pYkHx0JOL5Vm3DWQVlOzKqB/bGLggG0ma/hHcq4urc+SNzLyjjcqy8Bx4
aib8co5aH9brpLIMuaQ0xsEONRIj5yuDG0d4gUXGqmLbi9wTvqVxPG1KjXoVK6yt
JmeX3/nrv4yC9YMwrh4KvYJcXKEf2f0pclfR/aoMEDRPLAjQWuarcEDbq0h3qGMJ
MDyvf68TGJh+ba6Ol0MmHqh0VSiwrOzWeI3LKCFTG4VUQCNlvLAeC9xofdNNe1/Q
rYhEvsNqfy7AVJJPIdrn//R2z5Iwz8JpsyfFBgBERWuiR0M8kwQ9mDZ4jL7iD1xP
/YYI0h30fpzGaRf8S6AgS42Jw+z2frYY9vBhtiShHWOqM/3KEisIRFZ01gclST7s
YJ3XhxREqAt1Yr4m8y1FzdYqhWbP1UZvNQ+j7MoQUS+kBE96JOPO29+OY2ifFqVF
Pgb8PjyRSBK32Y8nsghTqDFluVjbiS/LpJ9mWmfwC+gd8xIzL321LMHgdf34UFPe
flEr9YGnt2MeQcFoJHgjOtiNLZzq7ZeElxC5q224UrtXolo5n1WMw0LtvRzYg6I9
FyP1gjsIUt8uO66eNR4Boz82+sNvHB+0btlXAPNOKw48+1vhx9E9lG072ScJNhSJ
yTA26vitJpZO4WtjUu7e6qPxpmz3tGGyh6esvFD1w5mHphKny0o8uaPc4S0vjcsy
y/0y9MNHCeVDRP4j0sNZ9W7IWPsRTB5p5qS+NiOMJMFJuGRvPC0ZTXOEHJQbYrFF
no1LRUSApxO10nowXIXmz064qfF+freD4Ck2xrBk7mGwaHk7LeaglPK5KdxPt0C4
EIdcCyZrUuVLiABkDKjJqM0SRvtMGiW8CkqVfY2aMd/hQ/4Fxyh9cPyaXUqMuDcG
fd9varR2916g58/y3e5j2i2xHkYVDsJ+HmfC6aCIv1eKDNG6IkoZitmGxVIZ/p6V
53S8rZjJ1/nSwnmkhHXQ8vwG+JEf9XG+7XeZvDQaQVBUn/p06m3Bpr4yCDJRtTVq
HjGkz66icyMkYxWrM+e4sXsCau1XDL4qVbM/ZZ+hQeEtfB2HVKD2pqyP/H5LFAw4
Ivjnskohszahaf2CUtyI8dbcyEPfRsfTL90WbTTwqyZcPhSmvJAMOX5qU6VIaMg0
HMJYoUP3hsz759G4SXpnLszujwljd9UmvGlmQUtDkr4i/WmHJjzM8HaitII9M1or
3JAgGdlzx8+L/PTaKbDhQUAAGF1FMxPG0Q6Emjkn1CGrz1CMMh7SfdAK2UDPt64S
IZQO0Z1ZUpibQQyjAl3YaBdR3lrsnSNYCSr9JKZBV9tYgtIJmbZLMfS8zA4oUvce
4v+z3Em9noebeLpSgBbJ5fb3bYBszcwmDT4NRjKFsDruPmTWpRcL+762xR4sI6Sr
NMcfYt7sqx25Yj65cJSxnuoHS4caCuXrBJp9xAQKLbj5Esm+Mqh1oAqsswm/TiMS
NpoM8fOPbyqJea82c2lhtUawIEIAmojYha9LyZqXTxUh1qONEBOOI6VVD2i/t4vb
QIByTnet3OuTTOyfucKsNe7d9sVQ5n2D6WTOwNHQ5zJk/kX1VY4bqrsmNIpLSVJz
0JcTOut/Z1Ms4SwQa1fDGMvQMlLneZw3CtrShjhByczs+G9oCQjcpyQoCF8MzgvE
LqY9LQCMsAjUdZXnCnyXAD/RarDH80gx5M9OnVEeu3MzpN4HlBpNnMvb6gFh9eP3
8VwFkTjRHE6l3C3vjjFAtnKzO+h5JjN9/25ABfxF04sj/irDL+f9ooHl48NyWEtD
OufN1wPwSgAPdCAFU5REgzEtJk6ucpMn/hs7Rli4pKzh9JMVnCTWIaqOzCC9a8In
nJhfmPqRCotX9IvXnKxAahKwWUw9CNlhwzyRGx7VLbJI2dxT2JnfY//nPQ4VfN9J
NDkjrp7r/+Lf9KuGeytSBwP1Z1qkU1JAEz4uEk3HtOUyvfhirOqvBp4i8BeST2Gv
dcFjgvupZUdOjGYlsBsWmeAhFRWQl+7uzCa1ud+eAuBZfQCDCJ7Tb5rd4GD2X/pe
nxzSQhwGSYM4CpIE5oJABxiXcFoygiBmnAz1Tb23lBPelmQ9t3GhYMB70l4pJUDv
DDdmhVXadlhfFec0ZTOPTeJTZB2OoTTtC4TeKYziQYW+mucdAMuJNlUxHSTz9qx4
zosFJ16YvcD+0a74n4hpbpnbXJEjvMy560Etv4xhZvmSZrD8b7FZ3vck1ntMJ78u
qIHoaulUH74Xpfgb39rGoxPYoC5gBrKtkBTvTlneyQBPN3XLC72xXze55CqSePz0
F4S8Sn1ouqYWtGoIEX3IYYEAkTpE8QDN/utxQb1bBLNyUp8XqHIwi3nZdJ+AEX13
c2g0wEMboYTP+PbBZ9hWpxJeQLpOoE6XQGX/KPpU7OkSpNuVbiF8hEKUznU89Bpi
7nVG2aCYTChfummivwI+0lZmNBmnCWJ8u8KOnq5pd6HkzCCTJQav9rpMY0NF8xMF
vsckFxiIndbG8GDRVF+RhCV3mDh9tTxNcEVermz5IyRMhAq26rjcy9z1a5Q50pVf
carm423WdC6Lg//jrum1cXRxy3ufV9WmZyTXVXYhhvDcIHWSxk8TTuMrEomY+KnE
evpZvgb07GVZTAWmEqIIXWVglYYAnPq7PHELaZ6kChkTmlt91Zi7pG/tvRyrPRis
J9Re1BZC+vRGKm5b/DmCgYeipJ1RK5Z6tMPZus4ygxtGNLGJJXaPiC9s7i2eiAi/
5BIpyTzuxSbaXnqds4LGz1LYZjtlFHkDPTN5aFoxhkZbA5HNfK3A+Bwf5OtP1bU4
zBJRPq6WAxZriWwWZeuN0DifbRNctL6XI8AcDnaJYcNVLA/WnxtRZAnkMYgIub5H
qZkhyENZbGBvklxnYNKkXfixMcsZ2u9lm/ZFNDbQlYBUjLPnUURs9FqALjF/VeR7
HQv3WGWOuBAwemQ1MeUtwn1gS3td67R2+x6S36LiopMmg+8OsbWhOCh1yCt+Vz6v
uuVSTNJHx3CHg+7xux8SRlejeeoDj4RDs2NxRYviKmaiUpQmTbQNi6+vQLgAq/60
XFPZpb/CC3Ysja7u4lZLUx5PRRruNiku7h5CROFBbVNVf9bCxVCRjA6C0GEXSDBi
ZVkJ8McWbCp0etB9E7Lofq61t5V950HiNq5PXaPE+azaSiH3z9NRswPA865cVLtQ
h8DDaZWQM9h+K+826pB206Dh7zLke+5ry3sh/ba51gKKMZtz8QkpbxxejArFXQDr
1Uv2THyDEusJMVGmko3SIFpVxwYiW0ElIbx/z2hB54WMY/X1Rul5p9fseW1M3fc/
eWxyvQ25DJBH7BsoizpRsuc46HV+78HHJ0jKxD4PlOma/QCWVRtvnoz15XQfi8L4
ZuTYHjBSN1miruTNMvhBKAwK7zg/Gz8YG5JD3HRtxdA0W3jDwrxB64iMz6beRLC1
UOIXHnSDNVbc5T+uaMfchSi8XHqaVyN5oLW6TS0CcFGvsYgYWAKFK5QVXAF4pSDw
MwMp+SFbTTxH1eRih44oJdvPF6tpsNuOI0e1BX+pJ6+M145hHxjZnRTw1Umf4SdJ
0hNaEuPL0zebrXU4Pq3P2w9/zF8vR+aYXegWdBdCRJ6gY4Nj58n7AKj+PwyuHn27
1OooKQZkiWYghPu1veTF39D6ezLZ+MBn/tCFZG6sn367WwOMf0KFJAktMEADxW1+
Rks7DzaPIO3bfTr0KcgEUZYfsZJqXF37wZvtuVo8zTq87tpNHgusXywmivpgGQQZ
cTxRucbYnJWaS5SgpLeudMD3EiACi3r6u3CtG/UJWwDGgocOHgRnYjApr7A/Hu3y
tbkT1ahsd1Q5kUVMpwiD5Hpj79LWK/9VhjbA/TY+EV6gKRLLmgNrqyUaOwI1nLHf
celMYZJJsD/AFHRrvyPrCeFMNGu/bdugSi9wKvR28j4fbHwIFVAjIghQqHhUW7l2
9rtvR/5wBl3r2oyhuSIxSWzMVGburjAUnqeGfjJou9OA3P9E1taIx3czjDO64+EZ
X7oVkAfl0NDqGssDkp1FBSywx9KcTn9rCvNzWt7pf8Cm8Nk82gq3jSwccWqTdFfe
X5PdfNhv14+DF+UfEHojMTG7NwE9m9mtzEjoG4LCDvVrkfQX74S7URXTjpcXpzC0
MaC1moWmdVXrCpjDbtxXPjBG6e4yzPEZbRqHyak1ArgpgaZdfNGPuvZI+tPIeFH6
lRfrLlcbB9cigHatnV2fbppZVG+Dczasl3rwXpLaF2QqQnqfTKK4V1Op3ePJXDjQ
6WcLqvxQ/OtzcxOHq2dKUwCVm3uDttsHEjeDgPcSKKk6HGHFYXhW5W6QQ67N2mBr
s0hsByS3UGW11BVIuGZCfYQnPKRxwPKfR5yarmaZ0V18FzFgrAnCJs96oAp8jXJm
1ym4EdlO3Ow4HLtYIVONFlbHLJXGBRwERhTmXot90LpgEkj2TN4Qwfvlo0ptREQG
+TX5XLdAUEbiIIPFup+XlokSge7/6vj1q5UfuMKC9LbXpcSX/jOgGcExpOH2d42l
bD9H1DFLHelfJU3r5Q8rXlhhjlvPfoNgN31wWXmbEVXE9RvemnmMAv89cLLrJMRc
gJOeOhwY8qfjPRcPvRachVDvxY3gY+TL5Nr9TOD6bSmBe/BgJNT1cds32Hat+mco
wARdT4cO04aqWVXWAlCTjyfkDo2K+j2WbNUH79JdIaHIVVenXLDv2MFzQmvoXCxf
Dgjr/7VRN5ILTtfH+W5upr4fLRrtqgrhQLslE/DO8587kGds+ZYGZ7DZPiQWmkuR
vUcow+iopXWy6tZDnhsTCtdCtbQMwdFhQCJdhxE6WquLcZbAiVZ87dUSUYBrB9oU
wa/ENx4wMPXZOiBKkuPv+5AoM6Uo1dzP11NF/23CTSEL550yywda4A+lQ1klpW5L
h/JtNnmN8PFbNeWSSUpqslZbJTZu4EllMVE2epwa+kknUQvXcudpkavqencSsqJF
WFaj0WzBfCqJYO+KhdSs1I71ASbPRxqF0XMmPwhSFgFa3K2Xs5jJ4iWxRM14LRAv
5gAVt0mIHNb2LAHFrNQ0kRMGNoAYOYBONpanizrCw1zxwsWfaD7DMSMF/UUdJYc4
ICk/SBbY8QPTpgEDw8y0oCGLmOoEdnKUuwpW08QL5k7o+usvwPLgytQqXN18htYw
pExYcS1A3i0XjUCMpCtRH45DPyzWs0WgeilL/HUXznp6sqlpetggB9CSMPVDj5Kf
vq1L0d9ZeC/PCMkPj0lo5FQygkjkjSpKC5ZSD3kj8eJ+phS2AYHDFa2Gi/UPMnq+
fd1/U8XBVd8+pCQloGj0Ugr40ZoqyGPJ9AG51kxKEfD0TU5hKEOLHwFgEfsRjnib
VHsmosIC1viiOett2mdsRJNFSIwqwgHlM8AQKkxFk/bH8wvh/mCVRX+A/CrRGCF4
6A85RP1kP9quGTCxXg2t4VgdPuQ1sxQm4z1bEzcHxIPJFdNW9bQ0H6BfSYgCFyqE
RpA1HfH69gKRI2og81jFPax8wS4fSOk1bhI77u16JZUo5l30R9u9kC66U+/rbDhR
gtHZPoM2HZaoJo6VN00Xgg5UhC89hlcK/O7ce6gqxHD0pqpW4SgViEx2JtTWocMq
9Wpisgr8fSw52Qe3fI7psvIaecobohRk9aTxoXKO52WhQDwYisi7M0Z1fmn/lMi9
6AayQdui89HyCNPXeIQ4nJzisFultnJJC3rdF28MF1kv6SuzjotjlQbUy6KXAs/N
WWJm3ZCwHMXnc7Wf/hCfaBpm4r5mX/U0kfoySKGjMkojW1fqUyqB6yYL1jAVjiXx
hotWYlEaefZoRosldB/L6ismmZtbZd1fvQ1tHMxiD/a/w7EFvpCOPavLtMZXcnJU
zAWEMKYcBS8ZKqOlUKTL7xcBQhUtKYJy2rYVrby67tNjE6SoctDy0XD8NwtpK5r2
WuFtAsgU9+wE5Q+DCxJbWB+YDGmcNeCXLOvtGg/U18bvf4gFNRG0PlQlUMOgNA24
FvmUQUe19rHSvNMFbiGcI6LBYTDhu8byQeXVka7QXzbEN4ibagLjbv3gF11cwoDf
V7zmqeGclhtOKWgyTBsUaCiMUNG/RB/q6hxEPQvnX4I7DoN5v7iJwK+NGIQcUe1g
FJTBtAvZ9Gr/sggkn8cpAkp0eb9bMil/Sc9442bqbclsaOKpll1WHDSxVJfOuJ7g
BroQXy/o0VXCt00/bj7ZjBC5pn1/buFgxxM/ZkNuctT1tbT/WvZjCVbaVyoaDbgm
5aVbwLQZHOwXd2GSlFRbSFl/BRUOVNufNx5ihCpiwAAI7cAOkfWXtJqTVunrP8pR
4C/90XO9ii3YyqlXNCsHQ0z3w2/rawBrk5RIwysx1PcWFdSnQ9aeVVB20ab6uXT9
VSuoYcETSOx9XiaMFpE6PpatX0rwaqDRDbplCLuIm1gnROcerDkSTuggYTK2SfZC
054ApNEmvmLYLipFiOXhnfjrqfDE0rC59b21ipqVEY7PvSeOfXbyIq8pS025VUSf
rF80aY0v/HDG22YI1529KQsLo2BUg3bvpQm5AmT9DKFPKioTJBu7wwIOh35S1iZL
KD0bbxfyyObPLshhVuk1gpis7KR8wl3WVXRb5GE5Xhd/iefDucDGofClvC6F+O6t
eZqmBXuC3NJHw3uhOWyPBPw5VfiD/oipPCcL1+T3gL6fRsNYetGseuSRiExXrz4L
DbJctWVqe9VHJNQllKJPGo9WTFy4kFom6u0hzPW4JFNVAjxowHHEeQR1EF5KbenP
P2m81A/kvhMQ4bw4Hk2awEqawfD+auv6zYLTdyyXqgumTqhLRD3cLXRW5lFWMBs9
RjfzJ12ZukGGI2pPJpZ/cH6dRhfYlcbGHwy3llKg/8IbZucGmVAgZShqqAx5f+/1
Zf9oPDjpaDhN5vrlwD69yK4vZd3U8FLNGCO9RRx1TVqCY4adP+RRlIvXmttJA9e3
ZbrUD/D771yAGSSi6CwbSvr3fspENkfSfyzBxSFGJ4guWwKxRJX3fY1ld89ShraR
mfyNbazdR9L109vSUX4wZv1NjMtd3u52QdCD3thIspN6z+q57j26/WGV9te/fs9u
NhkspywjYPLtA+B/q/gWO23XtcpLdS4q7mAl1uGkhhKsrG1YW6c7mYlM+Y+0QRrk
GeLzPkYlnyRIwGOfJ4LshJM5hKjVVYMv1KQmPlE5JaIcnnuQl2dMNH2RvY+XXZPn
Kh1I2SgPOyD55OLLY2Chwo5ORvYWt5FGajeEcGMCz9RdJ0ReVeH4WuVeFJ8sY5Dr
LOcNC8l5LdjaLmL3duSkKyC7XlRm+cUv1WlZWPTJKlsgFp2rGr6n/LBGUXe1kP/7
gqecfsZL4c1ee0gGHYxUG2wYNrwhnDUinFow80VesHhIAEI5ur43Mui0QXrJt+kg
ztJ3TS6fRq93QXIR1SotTEXZ6B+DVP/XBArBguze5sq4salkxyr03SaokTMcJdrU
Bh1IWF8ynGO5Tf4hzN9ghwiIwTlP4itymJjW5GGfOyXxLPFxsX+CJaaIdn2DFaha
YwDRlg0ys+v13kOSb1XnUQ7r0MQv47BdVjx2CayF/WpuTP7dz0JwwqfsAVCKYD2Q
dJIkDXymBKXIryBiLo3Y3/VEA8EhtR5krOiNV9S6bWGYOrnFHPio6+tURPddA9q1
gYnpIM3OYs2l1scl9/pv4La2Q7xAWiC+AQp54oWQ3s9bQ0pJJa1NBreHiWYhapXC
90pTnlC0PkjanviEoWVP5AcquXw1W0cPRgtqb6VO5Uwzv7Fv41Tdl/eF5rIDey0n
T1TIsuQduRX/FyY0WlVoiOJTacx84H3D9L0F3KCGIjCx3TEGDFywdRs9J9xTfzMm
Ekoo1xJPxBKYVb4T/ig/3yNXUOQqNEthmw6RcvnXJxQ1DKYuEfH1iyDw/CeUPwHw
FXxSqA1foa63w2v/Ujop/cghSD9/vTD6SramRulCyxR27OTyWkFPV41Ps0NgpfXq
r3HEklzL0cHMT/+MfYvjDvO6VTn2W86RdqBILrKPTKBIAO8bruBR7JmPJluMgfG3
0eNVcIvQbu737I7+9UVW/E9l0+Bi3NBHu9AxYaQIRiIXZSNUjk1EMfIuBjmgbaXA
wzX37W63OoNUpHGyNOnDH7c2TfhxmivTqjrPqQ5bi+xf3gwUM2eF3H6eYCtPeGvq
amb/UrpWBEhaJ5yByIpQHUekpYtkURRYVi+l0bFy/Wo2e7gKigLXdAxM3JSJrZq7
QHP9PYkqdFTSvXhTskZJOCAhcHKN4i7s/iHk165RgxlgYZNUgVf9KjLGq6cZAYMh
YzaN4SxDBtPsOZXGjnONnQ7oyTKIYI3uMLWNQA9pZkKxVsuJu/1K+Rw2B9b2GXxF
SWSMW0Tj0bwArCTJ0t/YP3s1kzWA0mj/DKKDXmzdhEElTpezjGPGWe6xgWutOQBo
oUs9kkJvu1f3i8MnHpUeoM7AuKA3Fgw89HBYrsU2w95M20zVIKdfzZhH3B9b8FGL
NzF8Dbih5sFb5HEmQkuBi13/tF2Hifs+lDDiQrALLSM7sVsn+6wO78AqhmAFaUbl
j2qZZ/djrNbr66Pgq3C1cZLTt6YoM6St8K3JI+CEzrl6AoBEK/NObhIPWjzvLRCh
8iPACS8ZAMY+CaXTk9u1gYMAo49srfJw9qiykNimJrnPA22JZTuUssB5gFz+VbNR
Nxl1WfuIokmJ+YD+twBU57EBUEOELwJvQPUmT2XiisEswtRx6AB8VLjsdawehms4
6XfFifi+esRojqyhqxZx/VyUiQyIIHZLGxhmxFn4EfXj7LjPLb46RJA1CXPkF7ae
cS86qJdLC9q/4se7O67P1ioq2GG0fWDwgac3Fu48hHfWYYrCeQ84E/ggLx6PpCIQ
yQxJEfB2lSX8r2BAM/5Le6AgXBGJI3nN7fU+me8eY2rogSv3txO26nm5A3a8pOOh
zSBzLQDswIU3eyMDk/LOfpAeova+nJliTzTrpIc5hRsMg68hUihU1W0zvXgS6VHp
n1dQeE1QDA1dO5wsxJVfE3HXnz50zWtWwuyfMfZRMevkGq8MCUnPkWnQYftCAMpr
PkZ1rBunacUWEdJ0EVsNR+9kr2IvXemgMSLpkZJLv3NjhEsf8lgJQ00onZVHYx4S
Iz+higwMJo80cotQ4FjgaKfClPSyCQI5SkV1jceIBD1ukvO50ppo/vdp9jTirxB9
tpdQYnK9Sy53SU0B7DVzkBPwNm3vFPDu76fH/PUg1xatYjzJ+786kf/yqUbsVFJD
+6L8owU8zvO2Bh5YAqVB6VKSngUqU3Ys9RnVYQzS7TQ=
`pragma protect end_protected
