// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
LFAYE5xyTPLAbuop2Av91RXl92kb02LtQmR7LnvHar2RLkFQ6RmLXJFZfGZ5FbHp
P+zNK5dtKA2SL/Od42XaiJkU/bb6C7n4zR4FJHGOLYLmDZK2ow2cOhtU7ADRsNYe
97UQATpKzfgv1/ciIoWcXYxQ7ie7+2GGrzM8at7RyKs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9536 )
`pragma protect data_block
Ir9RcQv6uXUvs78iOQCbjpA/vFxthw2tRQTqCSGamIkbstzNghUFBOeR4e9T2HEq
IqRNr4HSzAw8c9SV6FUUJk8UFFdOSNHn6/3J4jQDl3EfJPpCiRnQzPD1qEtLGV1/
D30MtIC+1BOiadTbkDbDgGSFLJ13SzpnuqIEHXbBDExpCnaBkU+KMfqiJCqguBRl
L3Ipmdg9Eu2z9vgi4UtQJtvE52ZRBMBMIso9+4XaSYoGRKHDRHfCxOhy/8R8yfwt
wf7G5O5Gn0qtd9Dz8+UNQEM17sm18LfDYhxT6wZL+//EGGUPnB9gyxz5+GdOWJWB
vOZQv1q+tQUXxeNLLpMaZ1yQn0qYZSkJZF++o52eyW42hcSKlM1NE2fKZ4v1TYIy
/evHj76T1hA68CVxtYI6BagGtN+r3dOQopOoPKPYQ6qHKcv7TY7eHunEKacEiNfz
GcPV0oeKiI294AVr+jKln75L1imYUdhVbqhlJJnwyJaT9YQGLfSRIp8rpfvmdJV5
hYywrWtlXx04yuqqLzuEO7mUU2U+urnuMYC2xzP8fzZa5eJ6LhYGeTHDNnb8XQRT
9ZB5NNp7sV1nje4XaBdkljjf8lIkdoMy3de8CKxkcZzkyW4GD8vtdfP3PR1fxpsa
zWJdBF0ybUKPK08tZFqjjQLBukds3XOb/nmWvYG0685V1BBnf2KKVaSdezJ/ml9N
eoQBhf5qlrfBhkQLZZwtFgulZoB4yzWtIMoYwPFZhwCPsCTWo9FUUUokFUQwJt2B
yfHdU0bD4ShLi+gxzM1GvXO5hgoZCVn5fPPVIgGNMnPIXs6ch7BF0mwe8f35yIBk
L31LnPRoLT+FmkpJ7zetwtQ3ZTIsDn7WvmgRaKdFMLj04irjAQJBQSzIW36z6N1M
Q/AYEM4I8n7i6iPTMwP5iaagHSeeVNbvFp6IQ/7yHbMtLXNxSo3TgzTS7jt953EO
4zBBhLgj/L/DQQQ59gYLcAteLvyk0ScThKsyQlZidStZk2QWw870oW2q5+tT0Sd3
9j80kyLNTg3oYdO1av0r4fqiDTTIp0YuLWflAYszapXlSQar14hIJpVDJk0g3ErK
wqgM1fVVuDSwRmDe97U8ZbRebqVvjgvYorzjau69b/AaY8D6F4rRNVII0vtPVxGR
XtaJ8wUWYqhwTvvINolXE+pSvn8jPGfJmcKwJ7FEX0jyM2hk/8BWTO5FZFirRSIM
wf+zpt+SR/XfH62TzSZRrUVWctqTkBlQye6qec8uIuKYbJJmOFWlsTMYNOXmtQfZ
jumuLnEuEd6EUJEdW4rBy8Q5RVJMdUYEUWtnid9jX7o1eXVsntXyJnmVOr9iwG9m
8cQMLPTDtskmcwaHm61GZx/ZuTI9mxoMbes2UPRhoH1EOVQ4bVp1EMmclneDr8wn
zZGhtwd5tMxT7GGuePPXbl1TjtOxsm8bHUtjvhqgzb75Jsqh3tlye6U7/zWBjzZl
LuEI9rY4yuVYC2d6nh45OiScyTHQcxo30PYv4Z3loOilEJ3xMF2prI39Gcx8MdzT
aopKuAD3yd2s9EKX2Oxg+wJRzvnQkvPJclEx+jrxF8B3iRUBB9R04gFSgT0D3vpQ
EJtiqaZIEfTzIGs7IC+O3RVQlN4hhbTnWY6v3W+rK8ZjgUt/qDEOsJyJYaEYjp4F
/JZlqB/NYu/4PjvLXDInBVB/1Gw6j8Nx5BLcjo5eVyJAC6sMEYlepAWLhTAUncTJ
wy/kGk4HuHyOUkpT7CfyLgXps3yiVmMhNr/Za7SI3/uY/4BexnVMe9zQzPqe/EBf
IfVKivMupclfrs6Qv0GMFRWA3W5CJWH0lhb5gg8JQtfkgus0g0Wk0X88z5zjnmDt
S3cIEyfXVA0ZOTTPDjVqq7Lg1cU5RaA8R39gx/vnN33cR38rufcDxZwKH0CLmKhs
+Cg7PM9Q6MIJ5rpBEox8yTQPNkzq/Pss2uBZQDiz+x+aMOa75Zk1xOErhMlAQqU8
WJbgSxeBQiPJPIWGnjSorJSCWk/gUOcoHZvAXGhNt+cZFEqVR3VyXxhISTl0XR/n
UM72kOWc5BQJVB9glqBjTuTZAtnKxHMr9h963rGZdC3x6ODiVESHeugobjnl1cjX
J5aAigB7rpLs6ST4HaUqCdpl7s0S0rDPrCKfGMc+vTh8I7+mywgHv04VwlMlm6sZ
8zGGor0MnWqubhJxOjBFiaayzO0YiMBejS1MnPXSdydhc95IUVyX7cw6pQT7VI++
CKgdnCmyOLZr+Xr9GCI+qaUvqcVrkdAxgC0DDE74i+NnKdX9M159Loq0WavEff03
QD7TVwklC8sSUW8QAoG0NnDkdBwgM4sXc30bgbdJrJipuMqLgnQoQQhQ+iFpyIQz
FrK/WygSbUADBj6tNGGWMuaakkTB6Fu6F/aqbQp4dtnhUs4mJ6ztq8OVOLEEOL73
/lkn30m5teYNo6Ha3slRti8mfwfKmB33rTKPim73REZto2dHvCFG+nGLDnLQVc4h
SjRvS+Eh2LClRCR3YwLGDALYK/JbMMUqBJIBCaCFnvnR2KOg9gJjeTJstTx/aPZD
P51jhHDO8YZ4Cqg6BogMDJf24FLW1d/fSsyb3bOGR2tow1MuLOW7Bb9krSJBzamT
pNg4PDAE90DvftLU26lGOCleiocXzFbSuHXgY6yYjj3I8bbwLZKEHiugXTLYCspQ
CagFhWB06tNVmT3Nken/xI5zhyALRH74L8xNXRKZTDSRdgL6IlfKrogqrBPB7oeK
32KThP1UbhasN4lNQf5AKhKwe9Q6GucXPb9XebdVq9JiMP9O00IA4iF+I2iasblv
0XYZs28iNQWYzpH/Is6Wub3Ur1LTF4uI+NN2YWlwHU0mv1MIMyXBDoSZk99Ih90/
3KxiDJSEAx103gQoZvPQfyHqqSi/qi1NK7DqfDwrUiJ/yz8zQortG4c1gq2qviPw
/dnT3F4Xth5/cEjLGED5gXBYdYQywoyDSWRPfxzrOlo+ouYHoyBLrGHtZ/cqK906
n2QaZKEfd3/03uzHTiQLkNgSYYNenD69OGRJ91Nevsfh6BaoOlgjdBviBUCsanG3
CBWJprBkLN9rmd9iV96F/EixAKTehK6KnG5UrlVtpc1tP3/CEBmbku64CuetFq6P
xfKGz1StjRFFtDHOpTh7GelK9+c8Ru8sCyx0n32KgQFrDJOW7wHy6+uQp2f0eFWS
cuPSpTU2wyL0vfd86pYAF8xVA3uVI4mrV5y4JiqPW4o6tnI6Qs9XzwznG0QtClz8
r3w24Fmtvs2GEvUjWuCJkeoIDGvRkb5qOz6+IyMua74brwu3krJvKfsXapsSUcFX
MPhNkXUme5EPJRFqJI7PBa34Jcz4mrV/D4kNwC+88IfaqgLepQmUQAvb4TuyQ+JC
Pnmda0/dibd9bV3jBxLC2y7P2Lm5EEYMqfletByW9UvmN2W04d2w+QrAhytAE8Fe
EktvPSV50dFK7J5CvtUkvbOqO+hdK9QU1E5eYSR25dGj20a3Vdevo0n4chjZ55Ni
HAfbD9of1cv95HjGt5DOY3wWNnaWhKycIDScWpOvtliPVc8JHVaP2dI1V2qIAOjX
mX13NnPPGf8EfP4yN/Z2zfr67ePd0SI+JcJAuT2NCcsbly1ZF20cSgirNI/evIFQ
1Y8u/p421n1eo7upviHbTKHIC6vDP315z/RD72xDfHzGkTzr/VxgU2EdpvVf2frw
QE4jd4uJhGqN3A0s29qT/zBuOwI3X/DHasbtSuGQx2o9RUwzCmnrhnnHarav4psp
ULzpJ1ck9vih2fZXKuENvqmTrdwaoRQz/9WT2kvfh1j0E5ESgrKBc9E7Kl8u2YzT
BpRSdHfDeO+VAQW+eCLuxD7xkYSftWo7Bter9EoGUOVjqwDBUQVznWx51I/5AQpU
9jnoIR5j5ERgOU1Ol1mmdLu/EJ3mYlnP7HHbHaKR/Jq3dBUj1kY5g1xI39k265+3
Vj/vU94ICMlQWcP0G+GwmASGg0ayjconUsG7yc1gdrnLlC7k9A7DZTqHx7YA97DB
aa/YNisdjmHNTNS9lG1WmLKSIS1QbyfdDJoIhZKiRk/sUKj402Ropd+geN/LzbBG
jiRGOJyyC11aL5XAv3/15lBaayKUiVZEjJNGZeLnSoXXzkY4PdR6JQTqUTvzWKwZ
v+lN/SchYJ2/ZtbJCljaPcoZBozMHiz3/aBgA53dnRB/iYZeZQq+sxrNwN8geZ1k
Kx9j+XaU/4JkI/82GGpwZuAALC5xBrj0oQ0qcWIrv9hx9dNdthhYOH51K5y/q0VH
TAdl1f2fbdGDndOcvaIcsuvLf7SU4uUxxT/WnBeOPU/NcgIAPjHn/kj6WX7/sChX
iLD4RSi9q185NFCIS1d75ov2bmgWit1MgpO+bDIl3v0tz50xnFKENjYq/eQYrv3T
X6wOVTdkXPgLJXBaAoTepFEIJei5g33e8v8UuiWHpG6sxjx7JwFQPJoS31HijqDh
w7ihN6JG27gEtCes+a+sUTscqqUYlVYQ9GxB19WBop5Vr+c/prIuE/rNN+UEYTmI
UuMbu6dB/MIeK7XdPdNFrAyK8x9jBkDHwjFt23AAjTF7ClHtmY+goChIil1rkVt8
bGMp38t/wCTnCBaZ3H1EZEGikQQDxTuvVskAY1Snu4YCy3eK0NqSLy3YAl5Hv8AD
3G8hY4HgAtq5iHYC1ulAclyBV/t9gWd/KYZl66jpeoxHwymdDg6TSiGQefvO1aQw
D8mP405Cvtw8iJU2fGc+a0APMafAFQNAjjDsjA+SA+4hRVZpDpMxL/5QSReVQ52O
TeCHjSjYQLCKrES+uRnEGgCVwdhrk/2dtnsuyi1CQMTGZ765yvXLhIcWBXx/wQJR
Dn3Qy/J1EfaAmCODQX+8l4H04HGX/0AWMG2bTA8hsPqwWt7NHjn44pAwP7jASKOt
Nlc6Of+SeAtGU76qD8U/0ZoPN4mS08HraNIOxAS8BC4kai9wn9ROKvY7dyJsehC0
A8930EGeM+6JlzUt6vPgS7Uatz7pD0FIiU0Ct54ohu61m/4+Y0YAJN4kwAOc3jGk
k3XtNYLofmNaskApbnV4bsbiHzdctV6ZnigSaVkb3HHP070YaNNCU6ocYyjG0lWH
IZ5H7hIgynydteWVQyY8rdUP1Ea7BTVINBTdimQv0GTeWFO4dD9NVEDL9Nt13Jpz
/hopRAlB0wbGzmL7cldqPUqPHUHuIZAWo317VWiiv1ezMNM5HO8L0Q+hXMwrl7L+
9Liuq3lvc1ScExMRt0vh82BJHvVriQ2sbezfFdkyHuaZX6QhVTDeOv6QMzlxL9Hd
iRgva7ABOEP/hanmvS97UOcckXW7yPhIcLUbXHIVUWPwNBF+wpRaRfrSa1vfo8sx
KUl0xbyXHJWW6FFH1iYnseaok5UwAeHLnVCWa/blDLQyGfY/XfwG2lRbp/QK5mUA
IL/ff6mP/nHB1kWz1lkWRdtZ30f4J3ALQj0kk67xcW/HtpPQeYE2hEe0XgVlgEkh
c+OU3q2wU9LlXeIEJHyFDzlfPHiazUiiMkChDiMTLU9nl1r9ryQl/WUD+Ohzd5SU
dAfNFuNjrgtYSLUxb3mdUdKnuCrcU1Dd9u3zobpjtjQmSuUndHrwdK+P++gpjWaz
eV9nq3PnTyTC6VTG/bhdMLNmFt4IDQsR3I5e/C8diuFdtwdX/prCXr3IiMAWc3zs
DqvYh6erREejD7mE48Vo6PMVgUlPsIBFd9vPRFULgZAh13yTpSyRFfPp+oBZ15jC
cY7HMsDdakj7n6K0oPOMCYSfEJK+M6vHxAZA28cSuv1aLY9IX5Q08qWLBoAPLkJQ
ZWZ34JMIpJaz784T7qVarZU3q4ZNzIjhfSGtCBAUeagMu31CBcvars0jzfa7cCMB
vl8Q9bAeZ/h8tLx0eREcQceP3qe2QWOShrgmTyCnLT/LH7ZmDJWBKT0wokbLpbo8
WkOxllKCvLMSz5IS4nA8iFN3NyrdrHOFpqw9FA8c5+r0UTKdp/k5dCTIYGzTAnK5
30zQaToYvXy4L5BqjstbnAN5UvHl1TWlAfG1uNSHTeZ/EYKZCoHTvRjrmrUR1C6h
eSIEG6a+CxVm+ePnCWt823s1xyZODFZPgDerncSO96x1qdpoJs5gAzR1vpsB0T2A
3zMQhouGMZ0mMGNHtgxBmeZcsuBcrpN1vij4nRhTn6y+HTu8wjdnHy7GHYxcRYil
Ir5m588GFrLHwPbir+odjlg35K9GgjhxIRsYKW15yUDy6kLG68tOg/hf9wMN7tZn
9A4kLaSuJxtIpzTqtxwGdxCkaal3XlUR8TjLcMfmWIFT1u6W38fe4stFOGO7cxi9
cpJC3U2hhesKjMr3uKkxbRuiqSqxmJkmTUM39lu1/ZUZYEkI2hBKjlsyqzW76KFq
8Gozy2mjjwVUTgu1VuL0RVOvmFZ+Qb4tVzi6zZlJbs1J+7CJHgBdHW9THAztLqL+
58KcDCOq2cFGqzTsRW7NG5dAtr9ENBgb1tZsao9qVCrEBdtaBj73HaYSo8O7YpVS
aGl3bUAHDOpebFvrUufbK6bS/iLBe0V4qAB3FV3eFC9TVSJqFmc3cLmDA3SeRxnm
xDlirzgd58E0J+GeXWwe8/SAk8/NanJzMAtefu3Pkf/VKiOJq3oG6Qaxr2mVrZVE
K2CTHCGqIMHPEO5Fz1Iphkrheo/BU+mf5VNQkJa6obV+1g2JZFFcmRFlqdyZLH0M
bVRHDm5FiKps4fJoQMPqAVwdy0/c6v1iqCw9kra4c712QVRFlG7L0qzcmgGPh9OI
/+jF3rmOd0/5lu+JvSdfxO0dG+xf9VP0dzIW/SZcuwAV6/GlFE9O9AOLJCFlSXrb
3JlqESASEIfLA1WmrU9qD1aES9BfU99oiA8BFKQJS1TdvN9zcP9G5bSpUEqGj+my
0WrvApZ/vd1aqmOOoWilwjFpUIWQUCIw4xIWAK4f7gxUDNUpesFpPRqdyCKiWMkK
PRPvVl2/RYc95GKRHKVQ3U+w95Vi4YLzStavpZlq8piy6ypg7mcVLyXRrJILzoxL
IDHDHcKChgeXeuyFSJL/rg4c8IwsrADxFo2V2mhKNtczKI0P5+xE+Oer2pIatljL
Cb71XH7QKEwHNeuraM78tnEFzsBW/89xJLZQ572IIPMyOaiTUGEkehosJHbJCHeP
vImqxBbvg274My9xwH9uuJeVr1QDWCpsOperrpKQTnU7bWsaPxPutODFL9dmml5u
f6RDIyCvOCCFeWjnf1bpzSIh5Iro2wWoENuHZ9jVWzQrtEHsM3O5PZW6p4zQ6Wpx
7VbKxRditg7CZ+/sXUU0JyZX92fBtlYlsO4P6FaxQ1zRC43T5oh8uGjo6V8MY/a6
Wqm9bOLuURfqrL8OIfVNHEPVnJSVrlz7TM/+w9gQaqOo7ctnHmU4w9QGNyG9ssxG
LfApPAEgFcEkkypTyKd2VWfAJUU4b7E+juM6PVVWdGtqKthF4P2YvAdQaCGPJaJu
Mipuw7IyxTlWIJZOEJIujmOTuCa9ueKkDymKllUXOvp7bZSbfQsLArqxZwmg1Gzw
EEN7lfAmRGEhljCXktamh8HB14/dQYLSwtSMoDfVrtU4jK2StJJw8iqbkEE9Fdh/
tkp4XJpGtYkmHgn2Jn60ntWeqCjVSCOp716iIYtvSkk289652Bfb/V4GDHG2JpVK
Vl2fl1PYCV1UausEa2HCECZV4JLEchVYN+7/DkBgrn09eZK5oYlxtRhSCqkSlzsh
vfypuRt8jwEN8rkydxNZYbt47LAE5vqCQfzvY18Zq4sqsKSHuctbvOuqDRnIz6cT
GxGpmJ/d3tIwNOYw6EwU3gmpuCRPuH2miYycv14vFc4HmB5fG4rCdkuAsJcg93XS
irduDVDJZODRUypWYwEbYlHY5Nwfg6cXp4ozPOnMAS2ZI8fgcuMm6YCBrpHLMNmZ
gIilzKTDWPhKXCin1dHT/Xh/JGSW6oYxebuCh82EQSYdh2B4A/UCzFksX2eRtNhf
wVJMJdE7EfMwWKfaBV3lZcqgNjaYazjC+cmhJOKeNtti6/ccOvwP/PBHOLsJ88ml
0zJXlTo6dV6TRZvEA+ZPDgx9rgL2pY42nmxWsCDjH8MDQpxSA1+oVQUmIQ2F0Syq
WD+byoCW8gdAhmrxETYswDK8AtCQHYGqyB3uqkvn28HcKDC21F1v+hWVavgV6jk2
g8/uwjqiP2D2Muz4XfMgZCCpN4RegMaoIDAS8IfrudmPXX1aNvzPM2dwPFF0u8Nj
gQrKqjEzBoOo0ndEVGQ0t+xJ2kTgH5F4TqCEkHwVFdG42i/tpqDSs7W04FZCZljw
Rf9/h5TUpg8GDMwkTxDm1SPS5FyWDCpXb1S/7gAdRFRs8Bu8hCj2NZ4XTCYZPwUg
BPBS+fRb+QQISkgb+mdLO7r/iSg6RRMvnDHR9yeAmaznpVFxzipx1V0D/0IWYiJr
+U+YJ818AercZWGAxqw8RBq3kplNqYXCCFNkmWR4bTDkiyQptlZYZF/GJOS3fu90
KCVKt3RrigCL5JHKQxYb+L9DPurRRWPWeK2pZ0gFlDJrpnjXUeJjtVLcTa2m1vtc
Z6pEAgerMj/2plp9GeUjFsqZ9EQHiJ43p6CI4j6FmFuhIsvi5oZO08pVLnPxOy05
bscxWGB2pRYhoT4JgNctfxQhvQ51kk2IxiwA0Ds2XMuQobKIF3sFdrKzllogKaK/
UvFRDL9ZAsYhP15nQ5AJP3KBFpIgd7/0Fvj+rR7zGgdHNT55K7MeXYAK7MBs0TJM
in+esry+BXiN119zw9LxYy8CDZsQ4dOxXYnK3B6glJ7vNS7iGRrEXFurJoJbi4q4
9rEEYjrbrdAbJgKqMyVJkoIjijHKrhxMqxx4NGI4/J+r6kjwwRFM2zlYhu5HBLVy
t1gK5qSjsvmldBbdiIj3Sn828BfJ9Ng5obz7tnN2lBQ2Yjc38RgGjTEaapW0RcQp
/LBuiUpbtm9ku+dGyMocBOb1555qpl2naGzJ08f+r2cE5MDHukCX3075x9gG5OQU
6+QHQdSZGOwWH/5uPBlsUnjE98Td3zbZZq4XkUq2jVyrhVs1RDxFk1IC0SyBkYr7
O5xGA6ofT0gIpAgD7tsa9b3wpfWtShgkko47H9RBleUfZdFvEt+tZ2F4VqRFWta8
TI3d/hUveoU3u81svGLgtH9Nh4nIlud5Dgz3pYXi0RahwgVHS0wRDFYPCzie1T32
fmjfufwXnhAgnqREfDXyAm9TXy4r+Y+y2BJ5/I9AeyTTBL9N3/23GdaQBRRW77h+
/oJnvAwHJb/cQOcxRTePWTtR/ymX5B6ddzFunrdwsmDdgZGkdEJ9JVNYlc+rHDuQ
T+XVtV0w0973HnGa/61tRN7gTgRn78YNDre0X1hcoNez2pClHF4pp0OKovY4C+/j
xRwHPA7O64RXd8RWqoUuWzYRSSBFJDNa3TnLg83x6J2OtdWxSjE1qE9YEIyHLrIA
yi06zwJzVPIMLyO7vLBgL5zbw9RRuPAj1mm5lF0zC5x5Iv033DPqvz85RHp5Z1Jo
M5gA2Bbv80PNiTt2f5XLa3FfO9HZxAgCsrw5t9jQd2RClDZM8ljeiNjYrT3zx093
8CWTed1dVLJtVNEAyOUh9kKTa7L0e7e7rGA766CWwcQF/v3n+cxAhB7Ma2Gdfrz0
3AB8K4/WvtkP7Ork9a+PM1aA0tKac/xoA49XZXSgTys/v8fae8skQKZ3CoJ4avxj
R6JKmtRVuYok0W7yAnhlUwCGUe0AlQp5o2SiaQiIxxLI1da1R/nIZtIqz5JPwAab
H23LopxvHwHfTXUApo9pxZ7OzsDiU9N7S5TWtny6iASh7SRU4ZbuCIib7M5Vu97D
tFcjhOmk0fTT4aEOtp41o76vB/iQ04uXu5FeYXW6lPlDi2smgtnssYacIC8127Mv
OG1zDZ/giRXwVtydyb7hXa5ZWVNpMppShQADfwgpJxC3iooHktWzVLTYJAouAR2X
zxuJGPyO8YaU05pZFOVBbGCyYQkykut6kqrfeVFDEu0vk1Jko3+FJZg7/OQV+U62
ZhVsYpZeCyH+uTXjZrj93DNnY2a3gq6suANLdu3vUyarXioSpy93bDV37fbEFNpY
5VgVWJaIumG8/flI7ntp0WJUnGEFqv00t8YO7zF1NrSCDqXWUrXdHuRPjN2TDHWo
A5pmJdNCtJ2M3Vy7XF3d2zInHSwWh57AHYYl1OfU7TKO+JK5NsMSyYqjRovwtsnI
tQBouxVsdrjEklvrzOv4ZzoLO0dprqbG490bNwdF/CEuaAUp/9exa4dj0TCz9oUs
bUy/8vzZTeXfynFaX0CjiIyXYb/cU+XmsmJ3UhB1UPbw1FFgqIRkWt7++SXPQWbl
CyCQpleU8zhFjyzeti1KtYeVRThDcbqrH0oTx8iqRZarP1p8vwfAqmPMJjOgG6xd
6GCw6PGNnUqkC+QezKqVm/ioDogAUZKVddWIC7aCJggQjcV8hFNYBu0FVhfaEEls
kEBRG+6eHRseJWgV5C6aqSdlzfSVYLukN9G1Ox1KlCQ7wWw/JHxJSJ+K6bm9YRVA
/YlMxGLECUzePrqS+6JQFHHqhhchGktU4dDOk+0tK03Y6XSXmdrGnHVVAKh4sjBO
sZTdJ4kBSvJNiTrXfB3noC9Uj8/zZ0U9IW8AWSl+tvVUaTeJOfAr5e4vpPFx/U3F
9BU9SX1C6h9PYvevmk3l2FE6s3J+tJc9dA5/7NXGfdBIww8QJT2b4TsB/Wlgymr3
C+v6whtoWN+eYVz4ngC2CqhCD68Yjk5LPvRNljD50w/z9pccmKoWDxm9Ugvfa/FY
dcnqWwtbdUux8M0k2xpawdmFLNdyofNi3qr8fsDlo/pQmrBs6fAZ7NrK65YVd1VD
MD/XsfcY6IW7x841uN3g5CluqZRnSv0YdkzIfN4BNWc1Qg4qfsnEuOySeO+dymkL
KNLvxqIV+qd/V0BYg/NlKD/2THW00hdwqG/QjaVbogGBrEC4WujwlUrT8+kR5rmw
2yx/3dBKrL1uHFtaIy2compI3MCQDira+TdVeF+eeb6+/aVRm4UcqctPY0rVXK+E
gIqg9OtfVsbWvnH6E6qSUY9JpN4omFBD7qM3X41CyPup2pdmCjyUSFrid1FZU3P3
4HMp+B4y8dSBvf/RaW8CjKk52s+u1jpQun9q3Ak5aGqqg6l9B2iKvXrgnldKW/O0
Zu70q44RrLogTys08fi7lPqiud1v/K0uo8bHqAJLasnaihRvoVg9TXOcDDDUKCPl
QM3YXOfZDKZ6eZtR4FJhgTY2P42UisrKN34/8qaUJzN6VFpmR69xvkgSfzASfcir
RsF1OqFK+ecOVVsmPiHxfZP6Wg4tXmxUyQRT4cUk51xIn6eQycqv5g9tFzMeFAtY
+M+XDUGsGr+4veILxa+gcvvRuTPyZdfyXKGlRI61vz7EcDfVH5B+1uBSI+4oqP+a
7O8scRlxk2tjyYDqRY1779LGOBOcRb/BhyIauyCdtQYN+JU8JFrgrfoDYvhDK+YS
/zmP5cfI0nRl3pqZbhytY/QRqI/pESsyvVeSb9GOo2ayksDNLRnjgtXGerezrLFc
noVnCeJY1UhQj5IlxKKftPW+VsGRjPh80CDEbXGAuzFd0V0lhYQr2+DWzMYhxIyX
OjvQARpvPv6E/AhNAEcB8TIHkiypRjoCEYs0Dd2F7R8ZhKhn+5hUBT0I5LfVIbPT
FHgpuOhMCLaUo6/FC/8RDnqhD0aEqoyYd+gEAgSi24W1QscnCIpaSGXnsf26RtYE
3YpV5EVJaRQr5f/RflCvpyXCU9MOzQXYurb646twOqnNVk2qTF51+PT7PgP0Ol4M
e2ZT1CKQUsI7fP0BnuuEOeIElwNt0gUjjiarhakx9XjwmnSlKQKZtHhsd8az7UZF
JvSDz9NvkozT5XitrQ8A75W7H/+1cPocDvGg/huBAqRUrKrr+Hk5LS4a0C9ryRVm
LML82YMdBQ79ZmxsIBV49LuldjHlQQA+z3L6zFaF4uqXDRArnlHB07ZstjXXCMHx
hfrxP6I8Gmvphr8hnw+4t0oq/bGbtLs6K2ZtULQtRaf6doKvs5h97J2ieOwrfSOv
Nl4/fmFtt7g39dqXa8nAPyY+zEIkbV1Zc2rt8UsWqyEGcEag4+a2+OKuD/DBecBg
g8W1KKoh6/h7Fz85XEkhj/LkOVTZFU5BbXZ03vx3kqkfijEcHsO9bnC89vDDnfTa
ptnRvuParlgHiCPo4GF/A5zpI/c5oiFvkf1+GmqmPhK06CZgEeHBu8bqE6EFuAd/
yf/M6V+Z4L57AwriIzvYqtwXA1D/U/LuxgD7W5N0GBz7r4qC47XZyW5D6Exhz0nh
TuwtSZJhCk8QQ+0U/WFNJ+2Am+GVtgCqwukl/cXcfuwGu2iVs8dnZs1wG4tk9P1Z
Uyslg8QFm2DsbzXF84x9doOYSja/g5Iv+98eaIXNjlV8/yNBjjPZKyrDRKYQnDnS
00UYrReGiBQk1m1/E4O5Ypr0OQeBN2cW4y63hSTy0x7BAL2Ci+RX9X7z/qtfb1pX
DaagsmHq/pqDqLYq0GwjS/9bFSreheGoVWuPHoMfdr4nRACkmw3SPkgcWjJ/wSAD
tBKpCOk8yADyNRyBxCddzXbpLvYOjp8+Dp3tH9G+FTMdwiinrs9d4xUCAktYaE8C
nu/TWZLAn0RH7nt449aijZ+qrysN7cSDjQZTZOxax6U=

`pragma protect end_protected
