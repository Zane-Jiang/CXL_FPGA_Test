// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
FpxP5CdlL87VFnNeJ0JTfDCRXETQk9owhnNAXeubM1E725oi3YbPtVEHw9vIESdA
8FHASAPfV/FPRoMOBSmjaOBdGzplDr27uR1ThSMNDxqqNnS1orbb1rfi8e3A94/q
UiRm/+SlDzGy2i/EVl/o7pkY5wuylHMUvQ/itlVu2Fc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
JehfJ2mqSrPK6X1T0Ru2QWPmmjJgTxrXs9hWpeeP8ISY/9pK87b4RND/g/NWslwk
0rNQsgxScJoLd3OOizxNzmSG20SUtWec5H2NsXCO/IzUvk3xofqf6rorxHWiySw/
f37HpL2qsdvZ3UiiFuq5p1ZbpSoG67PctzD1lC8R7+HhxO6eE7wJaQo8YLUyHj1u
97/P4zjxEyyD2vNVIKKINuh4GD/CpXCjiab1VpTfe6QO+9rR1ajktVwg1tDRjbmd
LtByXoSyT9LMiyNKWb5iIdmbiTxogtK7Rn+8EsdnYP6J1UpUeMTqPv4ES9U8Zwpy
iUhaByf/LnEKaCvIJbt6FjzDlY6+FV9pmnaIacfQ6af7SmAUy02AjRLrg0WSVv94
EyFvKRo2YRLalWkQE3INjIdXvJGa5geiiAvDhsEkHzpf1q3Y12rRb6RLSO2BkBIU
roUIbP2ZVcIeY9ZvlfoCnLrUD3+BErW+WNEUNWFRDAgXgP5/RKahtle0OF+FaCrJ
NEwd6J84ZIC5jmxc+h6BtRlszPcu7GZVJ1goA4qOzFdSkNymC6zndXJLbG5Iq9P3
trqVUOhk0sm0PIaLAZAK11c0chNwTHe8c7iQrEMlNwgYRMpOv1qLDM+hVBnPpteO
4k7LXCjbwZtE9TaM3sCP5ZkY5WlLtjj06lNhN0qIvALUa+0M0JU/OPqt9fFbaFXI
EjyL+ln+NxcWoTAegdc4FRJXBkkAoXy60zWFci01qfSq21M8jYiUB3TLdRkH0DBX
iM6dGoV9HLBkM+4dRoANVqoNuyTu7M/vpnTBLU+iAtGNwfRnjulfypLLfmGaB4cL
Mgevy+Vl4CmBjQJSuXNki7EMrC92pe+xPZzSYAHdYrPxXhFdB4pdAWsoCdh44zHx
9H8EfN2k9gylmSKq7ovEUINx/q52B+ab6Xnd8oxJukGo4aZZAVQTj5quIl3HOCUe
Z86ersilLRHFd+09nzMIKRxOZcw6LX5fNAAlD1XCvOh7s/MV3iSmJxn8eJhNRa6V
wFUBVZ1HUsZJ3iJWvk5F+Sp4y4d0zjdtfd4oMigTmrc7xNtZBPiKCokv6ijRmfwM
qNtUCPTzN8zvXnR8/SxgnEmRe1G8GVEdD1Ph8JS50YStFrh8QyyqMrnvpIxHkxBH
53GcuWuDvuFasrLdnvsLJiP68Xv9fZFrjNwC2OPu5tylWdFgHi+4CFj39VQHxSce
wNmS+hDKbHDH4T4tnYQUS5/xVVnOIicRFN2JC4ew5p+YZlJoC5LYzBXwBRNcoYIt
kJvwPOS3sNBYA/j5BMrAzqJxuisg9QvbH3vDwpCj+BDc/uvbl+LzoLBkHXDKsIdP
WTbRx7Z5/3sk38zG6/OyNpH8IFxrHQMlmByeRCtgPlIbP3lh65FqZiJ/IeBBiLLZ
znfSXg/8cVS6FtCuaKRPSNtVQsI1TZZYymiYFGeRDCRAJx3NkVTFPg20aNrHtF7h
GlLYGIcrig0xEsLj/19Fx7zPcq9ISIujf0VKhS6YGwZKEWBIjDzdSHwFBZxbBqld
/gFxTwHMTOU1z3/8mpxkm3Me80b06qjuM9hu3PfzE2SNd/TkRICF4/vufH/1t4m3
wW1GuWwIoLhn96M1Gof6CxpKfOl64cQaHqpI699HAWPeKJNQgXYsTKxk1JfbbkUy
I+jzMX4ZCrddrCVPPegTX970EDBK6TZFRw7rWVSAxBuvso1EHd2SjajQDMTYWH04
Vo544/Jov+wL6ekphM7mg7FcKxKL6LIb+NDvcMaLFvEv+WTf1BfStc4sK3a/i4sq
7dz5KD/nAgdwzV0ogY0pSjJDQSpVsafjbu2LYvR4B8mQ7R7mPkincWz/zOjQQA8x
kLGvSO6r0bplQPGsIA8AQxSaJuk3kpWr1An9R10VBDcMH86QfbfZWWM9wU+6rlEX
7ZQHOj4pRjciFcwstjGyqwZpiYfmuN5i4rTtt/J/Xrv0No9QK0BvsgCoa6twUFzO
W42rmYfgSjVvaAdX7RhWPr7xG3vWOTRABMtb91tuFi8Jt/IUPBVKeh/Yzylk3x3q
Dui/ykwqF1AJBj0C36k7p6QKBSMhIvK9aCBcdZj0v8X5T1MjsAzc/dnE43gEJs17
9O8Up8x501WeEuQuobvAq9ViJEK8dXAWKdd+FNJZVw5akzq768z2yT6r5C1ej90d
+SdB8uAyU7uf4rmbXnBFVxr5zeaxxfhCvMeLWd8eIYhx3uA0Xz3E36LwavoRoAib
MxtnLjqRfzPzoRnsn07Gj+WxU88SJlGE/J6o/q4ALbop7V+kqyl0Rk+wU4uD9uQq
r+wKt7yxfa5XpyRFbCONGDd4PdKuq61H09vuIxm+mgbbDsS0+y4RJwfbZ6DMDGsj
S39yQ3gKrEjKJSdkGsO6ZxkE93sRU3TZ9KP0wGE/ikV8IVZ8NZn5ccPXg0a3RGRB
oB7B/q4Rhk7aivO9HOtwnCpSzt9pDY3/T5bK2vLqm1jF7IGP2KA1W+cnB4fMs77J
No7EEMrAFg13+qsFxDL3V0h/+isTPHBzxHmWRoCUdDHeHebHRWEsRvojRuq0OwTH
a0GaGTrgBa4o6ViGfyv7DGH4yzy7YGexUPbZdlrBuNxIxg9wUE5LHNuvt4Oa/6gT
RnjaVGbCmlp5fsxivdbaNVtXiNzMSCd7l9iG+jvImz3xb/Ume9WurQrszSxzeMS1
DsMjoMfyNgOB0j1oa/ID9UiXMgg9W0U1nPNfOkvz7t3kMe0tXNd67YYB/tAnPy1P
2qF9spLt3OfJbrl642QqnrKTZHVUwdHgdJM++1kdsxLxE7cIO900p3yM1CxBNuQ2
M6oU3svHtjNbcUAM/EooTeyV/b9uGaxNk3EEA4BwucfteZgW9tW0QmnusCp6U9LJ
vqcYSS2lsbaqfkgvby1jAp/5R2H7v2ry5dhjEVHAd3OEHkNYdUj+o7nmE2j963ZM
At/tecKa4uAbsMWvrqIOEdZQ/7akbRdtYqDFiBItIQ1QfZYMrfBk9gJeGjDAIiMk
+u2bEJin1EiyYiFEX0+ZezippVs2LvpugOdn3lBrUrD12JwwIlS3hkXTowVJmzpF
KHUFV6ReekfDhwyLPJzwkRAqqk8WSt9OWeJRmNNfWKbm1WYe8srGfh/bBzCFz80/
4xh6g42UJKDwXDM+EyfccmMJaylF/f2ibHLzy7F2jlU7IQkaFv4IOk3o7vUG3WzN
lvRZMqV/6FXGq1jVVVSrM7H6Vz7SuROKxbh5u18GtHQu9KBFde6nT7WyfWIT4TS1
cVSFVdlzMppi7fCkzDdL87RT5KZgLlTPMWw5dp22ivvuwtHDL7KBGb2cOk1+3zyY
OeGCiyaQTNa5xm2G5ooTGlalDCS/XGjGm+Od3R+tWbRhED7F4hJZr0kh0dHM9IcB
QTC0r33kVkXN4r8FxX7xgNYJWqfKidoW/L6iCM8hqXV7t/5aJ7hIascZ+27JGbnk
0CFe9ieB2p4exoTX5Av9i83sjwEK1GnchX5Pzt+2t0Lai2XqXMe4U/D3F4QiRcW0
r8zuyBh2G4pINGWBtkWSA5do+p7h7TMg5g0E4pbAe+45fJ/TFNm9JWsMtjIJI3BD
WnhqwCJpeZ8UAr8XAZktc0OSzFGG0riDORiq8yBjaMt4PwKE/uGjyeDGFAypx0NE
yGZHY8pL9c3Quh+frsrWTcrN8ZeX5RoL/6ZV3CPCq6z8mFYeJ2z5dQUTbPr3hUVo
9y38w4O5Gc7NNlXeuKib8w+4H0EY2DgVjGbzFsbtWjoDNriXnobFaXmSL3WJ9GBY
5dY10uobH1I6+2y8mX6V8AUAR5xa2TBuoIQ4on4KX9yWQK8Qmvlw4hUrPpfBXxpq
ID7KaD65n+uU2ARX2oB9pLPn5SBKDIYXzLJyI84HpEcCTwAZpcnAsQSWiIIl8pHP
spkS7HoO6jizv6jYAB4GgsHC9XwjVKIF3qctcNwtNUJxQnLGtClFKG6xpNbvxIEL
+k43MtjitG3zDOP+gdue3bChMf6mPY8DEDp2NGXH8kaPQRUp0sHQw8THiqnMvaqJ
1qo3+MgaiQnVpVyMYR3MlxV3G56mS5hivATIBfOHxJVd5lgXAflkhQ/YOSK5KDSn
gX5XLdFmI+RJ5ATFew/tMJJTmV48bSERCsKRlR3W9ehU92JHynFPixa7g6WQKjg6
DDPsEXjV4TRMk0epPeLfi9TckGdRLwXHCjVhKi+IUKXXIXX7pfG9lNzj4R4boaMQ
MUdb0P7DAdT8h/qpiBBYjAzDBN6kK0h/Px5UfN7i1yXfrSSytPDMttUKe5qSTHw0
uOzwf6czZyr2N246AjBvZAHe4Oj+kliBBdG7X5+n0uA+gKmLshymI/9F6U37OR2I
+155S2JEpy//5uBCauJ1ZfgJiyH2hhLcsjjLXuuwmFefcdtnc+YqTbdqCd019NOv
ZZMDRcREJ35Ve32wTmd2oVtjO+LbqVUv0k4VOOoYUR7kIXB7I1v/EQEq9N0pE+Ok
WbOHIwmH4Pknq/yoNXekU53Eghg4hTg/5qUWKTnCB6vUPdkd9QRrD1PUGL6LbVsg
FeZZmxziXOBN6PtlwO+i3o6rnKx3kUx2Mv0+hhqvVVWBjIvjpInVQ8TrhfUNLkxJ
KUYE76Qv7lkpauvY5gk7XPl/9Uk/UYuZD0M6OtCxRyfAnaSDCfppmCCKeMRQVW2i
MXFoGvojyjICOy+qi+fJQTn549kJI7Hxg52i32EjKABmvU5WWA66PeEHawSIj4rw
T6w8gc+q8UKSrWo2t6qnIMxJLW5NvyVjTnDYtorvzq/13AIohMm97oCBSs/KqTlO
cXedPOc527W2SqcLjZK8sG29BJUE0EEqYgsoBKiQiyjMs5Kx5A75MMxLw+8KlVij
JPGp8kqGt5qgOGDiqL0idPE5EqB3wK55u4JlW0Yw8l5qnjYuQCfRkSWmeDazpStB
AeR+mnUeubBnH++xQ0JLd/F0sr5r1p22LJJ+cpkDGA9FZL2E3dnLZpVrtV6Zz2Kt
hlwYf4GZY4b37YI2VTvdaewn87qp7bbPdRh2PPDCJYukga7MSUtDe+kUpUzE7ta5
Z88g8KYmX/o/eq5hPqDSEeh2zACq+aPQDi7le1RPFO9iYqmNlEIdbbzkwJldYa9o
rTb1AJ6gSBqgRZaw8Q2USj/ihcxwCwsZHD26flW+wwpY8pymrxjdtssKQQWnwAnX
kU9Gcbd+v3jzFNyDtR/dQggS3QPfD+3xtoKJgTmU4zT7MVH0Fz7CgCwobDkMgm1d
VM7qC9RJYDyHjB27mUDjAHVukvi+ePXNNtrueWP6Y12yrodPcXAOAvMafsOYauMS
5MHDDIdkKgrl1gFvnQiF9D4dWOxGghpAZp9FqqM6l0SYdetHSnsZaIwcYUhITIFm
iDkN0HgoXxb89N+Im2C8SZv1cr3Xw/kX0yMZrBRLut6U+2D+ygGPCq0xXqNVkVre
lWlsfhFWNxjKydfreEuq/Ob6SZVvFXLIknY2xdKG0HH3bMob81dm72mk2yLTXij+
EoYwAbo3UjYFChOaU14KsZo+Ue8VBhygYU7miPeG34A7ILhJgYQfbJM3yCcjk9Vz
5f2A/cwQ47ewdKMPFphxoPIJX7HXT9aw0E5oso+X+Ia8+oyA/UhjYE92tVI4qgwL
XCsjIJAgK1UbotzWGaOoSg0ZRbNTs/dC+pvZX2zu4tM3yCNCzKuOEB0xazJm3F+A
ASwn3jhQ5RbsCXlM+mqFNQ3IcMmu1eB8S1k/hG57uTtoT8/fHBxAje9JEPmGNKDt
qEoar1svsTmMgz7I8h+bpkFuChk1nPtvTkOmehmilev34y4j1Y32Q12aAFAzcYrd
5kOGune+tUWF1YA30EjVQ7ZfC+P4ySxAwqJOJl18GXcftP/3Xl8jYxmmtR13KUaP
lTfXa9DrSXMAF2cUK5sgpcQNaju01yWn8ucpRkGM1QLOuydW4VzJoGQgFXn4DcCs
AfxkX8tIxvcs5Suz/Nr8Wkh8JxWzG8B1AKS+ntNHgpTsNwMQiJQGluokvSp9uD4V
7VQVPGmukf4ghJVHaH422PLHwI6of9QtUcv9+qp3j5CYXSdoaZRsq1n3mnt6YHjd
1LOPKEHr/fLYA6/mg0P0RGw3WVfFeUDvc7qyU1jz9mYOnYa6zOompGVLY0Sx4B/c
2beDa9IQ8BSaC1Qt0ccZub5r6fjXfTsU84WKKP1i95ipK3nrxExoiMipwjQxuqi9
KmxZxQbDzZbySRqn16+SIiKNfRJE3ONgcu3O9CUiF6gYGnuBTfGkbdy5IZphL2Uv
fGR3WbreMVYt9WveRibHyAqJOymz5wGy2Cv04GpWfdSZzypvGTmyAgYkR5KeDxjm
GOh4ICaeu5UCqlSMm35JC5uzz9hR8F5oIT3R6/idWE6i1dvuOdzO1LIOqE/Enku1
mi7QJ3OW8pFt0FEiViz57jV/PjXH06ODko30yKiPXpYEvmNlcAO0nna1r4zXgDni
C0ntX2EzI60Bm5Ui6hMFMfA/B9aWnVWql4ad/fK8Flg21d+MJf5PZpjQz1CSgSPf
Y8QF7uG3YAgMXKqryHv/NA13ADbZFaBVNNv3XqvtCM2ogXOAqVjhP783RSEZ7qVP
60jxOM6uAED6mPGYXbRw0nH6zKWJ/b9CVDto7/ZTRN9gQg18nO72TrzKB5LZ8zNE
MZuIcuOdGsSqInUOlERAK2/PaReAoTGfBImYYXCpf9CbdH8cpz11hfrubxBNCxjO
tacTcMTwr0uS3bfgUJykvBFC/CLYWWlDMj6V2bDDghfg6kzZDCBMUrDWlf3DQ/iu
NwOrOpB3GbcaITdFclyqgH2w0yzx2/KdYAF5kz5rN2M2J4ob3rYbP+kgPiGZxvyp
g4B7JBBfy7ZCxTD+qS8wOX8vD8YRXcfPPY+Ww/RIKpOcntkteCRCMEORjGmQk8vJ
0B5yoNOV0/fIdhtf9uILa4NwrtSjidqTscbbdJ86jtiz5yoCbI6cwF64IvQD5ERP
kJb51/gB2wqFRm0zhGs18LSTYiFji3sWlWGfHhYCxNrtbucjEHX2HiXIPL2fgVrO
0RtVe4i6DbZkjAhGx4pM1SccVT82XiS2MZT/gDxYmG3mnu8QPlyV3zFXoyuFy8O8
aGxBh0M6zD411bcYlixZiHM7TK8IUSmOPY/jptl8WVd+pjpqDEdsIea5AfGeEZmG
FUe9Ec9d1FDuGkYrvcNaEcAJzM8/ToHcR4iNnURuxSsP7/7ZBHFWYXbh5eTUcSpQ
kvX21ITQSirISwFcl/znT7wJAXJfKLYIWMU+LVrycXJSwDqi3kqpMBXMfzMP8RfU
g0GeEp2NN/IhFK6u6ZJoR1wBMKRT7QBy1LLE90MymqMYzE8AQ6O8opHskiBBSwZT
MajQ3PjdrVIXSyjH9WVFHh/Ast6PXd9qGZkHN3fNVsTWklUgXvuaeF19Acgq/dWC
hqcFKyZpIrfi0ge3I6YxCcXnHzol0Pe/a0but0CG0matcXOjoHNQIZAzmCN52EYZ
733Ef0pzouq2p0H0LzmVpqNmUBa4xw1ZrMDlpBxyJ7rTVB8AnwMHBr+08p2KsIX/
fUwvnT5AHHHzk6wpzqZGA4N1+oYGFMubOJGOEZjXugsyfZRc/L1M/0r0AQZFSKOr
pJUtf92o5l1snVrec8ZzH3boYXIZfWUuWVYI0VgKevLwvlSyDRcXvZVYPzCatG2t
Cs4RbcdBnZButXWP1k+H0S7rvZPLBTkPg7ptJAnt79CmNvs6ity9xC/rozpHw3nY
vEC5+Z+rkfwU+tja+vHigqIJFHInYE+j95KICfx0AygDVer0k51CebOJg6FtvJOd
f3I4MEEyU/RPY/sAXCjHQBDdyuY+0WiHM18SyNiQb21CaBdy6XgvMyWVMH/Me3/p
ucM3wjmpPUERkVvtpSzLh1snTfPObqcw9UmDHjfbJ67VFfcw/cfQoGsgJ6uZDbhP
8t8ba/QviwpTsQrMKbujleWQEvHcV+3RUWRXlMtkKWFNSQLgi/dTYovlzDkFMqin
ocrkih7GTyDqa51lhbT+eE3baozu9DENaadoDinTe+WXpjO6Km2SuwXzvKVe+Bdi
fQ9QcQ27ma3cjwq0kcB33SBVk5SRcPslAdaBEXdVBp7TsFwwAtRiw2WryDygfPMt
tvtz7co1Zbm17anVJ0Ty2CIp3PxKZLWgjTXp7xI1gtf3BDIDobxjn0+CeW2Gh1uK
gqMblMS66N9zEWGhgDpC7Iwz49aDmgwk2xrxw5vY6kqUOgU4IE96QkCYbfc4E7KM
I9pQtUvIgujaM+H1729elIgKI33s03VxzRP9K4TLPiq0UQF+o97Nx+A29+5ot92n
2k+j9i6ZmyjzT/+ElID7a3uWVa/hY/U2ATV3DtrA0wXOuhCnGTeeV3A10YmBe2aq
QlND3oL3JWCeuqYc/5VB+72xThH+y9yz/jCYZGR1eQPZxWLI3smkrXcAqCxjbYP/
2zLc9NVDVj7fWjSu+6vuuxX6b/ri4LlHnYqBFZSsDzO2k64bZGvNRHndu5iS9Mut
Fwe6K8Tl3rLj+4dHv4X0jkZY6qAkEd+FpreijI6/sKTKuxrcFGLUeSgrBkq1vuGs
cN3Z4Dqyn2n/HqSM05/stgmc8ly9I5apK3+Kv+gEyspJG6BPQqz9DIA0ExrZq2NS
JvJSSeoHHgd2eurIb/Xnbkbbashrjd3VGES2zTAMX9cD0SFha22jGlhZhaaxP8De
46zRU2WsWvWk5XmpOe0I6PCcV7sVzEXC/ruP9UYhwdvjj4jjmNDuYGybpvZXuCIU
HK43fjhc8tR0Cj4mxfcBfgS/WicAfZzP/KMg7ZD5YfsuJ52wVbRs6EvnEtfUIG5k
fZ9yMJ/0pe7f+EOb1rmdIIUqrIIjAmygUbth2Dp14w7xpUgNJkShewwXUKiDOmx9
n9QCJn3Nmqae4rf1o43baThxMRW2QNPgt9cvuLa34tlSNoa0cCHc7mTqIUPtV74R
9186zlfQIyISYJDtqzgEP+LndYfIqUx+s9vMuan6Xvg3x5r1leAD+ykaGSnZAgBd
aBJA31QiUpf8o4b+cWpPHW4Q2rgbaHqqsq7bOkFL1F4VpKE3iV1zDRWaUZlDuX4w
Po4gOL+L/7EcbAd1gkA35Upa5GqVBAfslb445RmxBzRqAhJ5m9Xj34MExsbSpOFC
XiGnpMpz6JuJws4UrpX51Lmx4ybCKoaWhb3Jg638a6jUtaW+aRd0BFPEULZ/1but
ejcbxbPWOivo0N//HIa52E5prDhpEhBT8FtluY/MT5o7Da/Cl3TvuFcW9pKVp/Kg
zYmmOnUit4nWA6Eu9sZ9aq0gsgESqNBcVX6ShLGLXCvl08tQ9l4UxcGGiUTd36Dl
eaeSaWoCdnPuvDBYzRZ+oumscMPwVaUvzWOX+Apm4DtY4M0iSa+hHlFYxcekgDMF
60Y9YKcsvcpDpUXXcRvLcXX2Pyxm6duKZiKVv4X7qTsE3haPk7fjsA6yCk3xC//A
TohtA94zApUnnamLAzLC9G2vLY0fUokjMklyomU9ZywRBKTEOy3z6iG8zKpPo3xk
xi/vvSKlfTuToCiUWw0Rjj2GA5RFPBDEMSAXkOjH4+wns6wWuW5Nnxe9UsFsWiIX
d8CpUhqD6B3DlJ95ywDbyKYB6AjBc7CmQF27vbknBASo5I80Xk3WsJUS6QlD83lY
dD0c+p8Cp5i5NqRG+WfQc4/80veoc5wf38xsRy43RuQvhoEYcegslGrDym4SVFdk
rSrR6qiKa/CcKFqyLf2dxcyumx6RhJp08cNcvIxwq7jM/YA2JYh2mMB4iFkYFCt/
bP5U3ResiHqmcpnEVqsSIyLHzg302+WIe93xvjpEp90s/zx8QoZYckpHowNLifHQ
3AF1hh6ynwW6QWkObiB6OzvNJx+Jw/l6hwa5KwUTw38i3LDFf+x09uOWRwdPIU/6
YQAAiqNWzAACVWNONWuHDokb97R6KnTf4NJiS2SFIuddElg5XayTOm+TFSdM25KB
VvYAERxEIhmfjVU+BiqT+neEe5aE/02LvRVyPIPuz1bOZSpsJIlRG9rLCK58sQ2o
+fjFE4Z5bEWPxKbQao8VciUIC+z52uQIgt+n1Jn2wuHORAfc0uVkOYNEoOTiFFSt
Sy4ZiISS0xVSHLyTLdPfx7q2OSlaw6/Rp5EkNSI2yRoCJT2JIZeV16naNdLHUnhg
oPlHWBFY+yA9zLx4KKIGiGznypRg8Un65F5iFafMiD6bw4pEFuTPxIN4tR02KrLt
+D8+/S7n5byzsxhcGUWzhizV8kZE+5oU2FLNPV3TiILhppaHq8MzPdzoF19VJleX
PJgnDuxBoR0V3CnlUTmLtCJtQavDikxEOrhRqSUN19AW0zOsF6gZjSvHD8uztgpV
dk0SH1HPDBJRoKcSfIK46Ys9tbuPd/PyXmNV9hBo7AiWr/e8g0zATgM1kaHVFXnj
gdEIdsFvVWXfNYX9TB+2g8TsMzC4+ixs235zSkMzULbJU2bC5ao3n78YDcnyAAYj
/VNyP2+705BcgMfguGVWXDvi9CQOQgytUE68RLjE2HQWHLiWdej4pxfRaCuE19ZX
El/p6LggKSEVbk/3g+yXhBHhQrzsGD4WVBq8DQGTeiIHn9EDMz++Cj4hiZnGp5ad
TwTOQIFqc226gp0vTc3FcC3o9N7ji4xI62U1fzVIAIQLb8WHB4kyv6Y55p/cSi0+
59MsDZ4/J+kIwg+MA7pFNwUzcZErQS6SZh732F+/xI5hmISMgKfBTw8h5wDpOhJp
mZh6TOVF7hB25+hAFsstdE7c3Xo9LQhR4QR4YjqmuVc7IQKRnbCmYqodWC2iANCj
5Kap0IiQEVqyC8SRumnO4zVfvuaIMxgPDAfHPbd4v7fkPCyz3u8M7K3a4pO8tMhy
ITWQtslDU7fYwrUoS9u+gWK/2eHMZROg2CQwaZ0e62x6ckwKSapx4G2EQfZZZAGO
duk+Lheh39L8tSTxg88iDhdKP+rgHC57ScN2gFcr6HxVT82Z1gouazMsNuxjeiyA
cHckdZUTJmdjzHv02TZWDqs+u48YZWO6bgSLljIKzVPmT6uGJNdJCmvHGAmNDKM6
Iqz3CEXCesgqHd4kJxvS9n2DFWzLZb7LCu5ypwrW13t5vy9CFCaXrR2HrubibYd9
KNTATV0tp7bm7tDGXOf5cm8/7olCUICyC/YkeIBM0gJ0Cxr3HOj9jeg28m3Vkq5Y
bhjjIZyL2IBlOG21m/iS2XezokL7Fn1ChSNXvlvFJtlQwg69B9sWaO5ou7grdfRS
NqkUHaMubdBL+/yf1augc2psjGJVtYMRQ+6RjaduIDpiELOwxTyPBswqYVuEm0UN

`pragma protect end_protected
