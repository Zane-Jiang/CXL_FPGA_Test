// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
vJ7aYA1F26okYODO491p7vyt4W5OGEnQ2uHDrgEJNmnEMjK3iGXSpdVF1BFNs7DJ
HGZb+csXD+21C82LOW0ku8Qe8hUm1D0X68ERtvdjrFe/WhhaoNQoZQgZ2RMOu1yl
Ss5twokVlMmkgAzthOCQLVq3Yj5xaqBCWLdmzb9CeSo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
SvV8rdF0s0pcXow8ogax4MQ8sEr6+a+7prA2CDQbOQp1uKLXPDmOxvp0HnOWYrhk
+pBZArh8+gh3k9NJTX9HvHI/HrE8hL38kb7peGUuzpX+ngCVc8MO5lml8K9qZcs3
9ksZrdvLWP/MXE8KxZDcABdLj6USxRKkD5cvWuaZ4X9yHufDA534HXOspA0fJJ5B
bHA8fuokUjdHeIPJrO/pWk+JnhFcpODWBA7IKWfQ373wrnY+T1DkkyduKrOj+ws6
wib8cxDoqlfESTItUQvWA0aM0o6/0eIZWnxEW14PP+tICPK1XoBmqe7Y6uunuMUK
ejzZOCL1ifYWRzqFFdq7CZOfnI9KtVaRIRSybkVfgXTERuYef12Wur4AfZrNYafs
PRKPx3He97x/uS7DIXticlEiFilaFZ2Qyacq4uQYAj13SYkwvpxYtFnYlXK2pgYF
Flh9gwQkOe15oTPRXjCRsleSMI/Ju8SJPFR2p75SGJ94ZNCRmx4Oib06EmuZ9nko
FY+wSr4NPE4m1PQQKYc5wO8sbSTa8tDw/KH+EjopH6Hl09LmMVEspNXWuuvWR//O
cqM9G3/1/97EaGqTWd87wZw5/a2/Pvf8tzw1E9FefmAFi4mThP69DavJhLknJJV7
L8474d0TQXXDr61SIrquLSkgWK8vLizVYEwc/vpiOY53f/qjK1tGHYCyoJ4iZe87
xMi/rquOBcqchKEmkmJYTeYCUQlHhqGweuSm6YjtUY+Rz2s7eyfKmL5a/I5WwNfY
e1+s/miM5RFdeoBM+l6wVp3ucSLY+leTOfoOgZmoUndmZ/HaVNFevUchuEaRNW01
tbYtBeOxnmUUAy8SooQKy7Bd8oebcyVvvR3fVbrrsDFURzbg8mXaxyIK23R1timT
RM4sqXzM1joZ0LuUGSFvyaS0g8Awz9PFrzRkVbbJYGD+N2JhzOMgV7AgjUwAwacu
eH2lejUCWiIlSdY8/BmLN7AYBlQ5yGQak33h+oFGkBLSRswukBrK94jdw0kP45R0
91dB8860hLMrIf5oxK6zTHn92Wxe0J0QMiT35uDfVEqWMsbhdF8cowgyuPwpQIYb
WWN3qLLzPv5HDbyk30Q53tJWE855ZwcpxcCS7PULMgaxDJG7q0hRZCxCtW1wdvq3
i05fbuou/Z11vuDwY4zEjGNl1DlVswYoFtwNFgQKDlPX8mpy9WhH55mQBWOmeC5n
yeW6a8SSC6cElsmLYylq/gvn3ZDv3Y+Blb+m2Y1vWKno/NSJb7l3ilDDFzjwS9s3
9F71CozwxlJWD6KMAC/amEN4y3us+TZ5+dlNeZg+i2Z/PZtnpRpzsXfmLY47tFMe
wyzv1e3msZBp/lhejEeTjWggmITXb5Yl7rmcxvVTktodLSVYRZPa3miJl1DWh7b6
LzzSuirYhOOkI/pCXYnIKSqzh3y44wnCdZblGOEfeB1hRlUvSVNLD5VqvHNhiRFm
AAm66fFi0E/s8KIcgNM3HQq8w36E83gRWEu8GxNZUrvMrFnFKIYXfxUFFnGkFOhs
zVBszo4CU5t0q0DqS8L0kUIKt3kGrDxUBlDjPMDMQ1UDaCY6jrEL/oKzAawHR6BX
fjZsyrUjf/sGIdlmVFJPqIoFHvmKDoEJUg5ycaiXy4+pOsG1K3t1gu1CP2/4snnS
px96R0efi1z9VdBwUKEZ465s/K0fdiOiEx4NaCrFH8t7VnZTutP+a6Dmc9Kk13Kr
cQB+DtCDpwNUezpq074TYC3QvI4IFr2FQKZiOqdELdGsU8u1hA5BlZI+NFdWPr0z
TZrgsOEGzmZDJuxe8vYbUwrb6sZ4iNB0u0uX1TVjCl75YtXMTL24H/krHMoki4+0
0zumb6Gg28O8WAYzsbzO5j+lG364WG/sCi/EBJtgp69Gm22PEgSjMqDQVF0IpgP1
DztoXQaPkcB/uxbJowXZ9Bdx9hXsIOgHwWKxgpuKouNt5PIygTX0PH/PSYi0AiBY
jE9Dgyxcmxp6JP2liVmNOWW+TkWUSJl4vdCyCgEhnZAwFkygQX4eCEXt7YFFntxv
avtb+HuRNu3CBZO1qsQX+qWH0eRcxHGOgBHsNr6aszNFw3IM8I9VD1anz5o66Vkk
NUH/+3aLnVIubfjrEoLKJBq0x4aAO/M+mDH/xzjFAOtQuL0qTUNZg85hpIvZ396c
DkIqoIwoTIrAnGcCWhBG4k6cr1oynUjD8yaJxfyWzBHgDnPAmOCQ3wNTrhOwjCFk
urLwfpsCq5QcQfVPJkBjIIcu45fX/SXI7axQuceA31Mz8rTrkjgp/Uo5DzAWwY2D
ITmnaq58VgKGFv7Rj4j2zxfaWYGxNI7eW162gx6lFRlb7J4TonPf+24Pd1ddWKKE
UkatfoDDN5wkah9KSpI3Z7LbU6ShHNjLu9PItcGYkz6RLCTqI9+ccLl9HqFQfZXA
0jdxNpLY9Hbc2ypvAFs8lge/BpCtdGoVCgmTw5ydaA9mjGfHtIcAb0AaCbbho7nL
SvwbMx+9hV0I1xzxgetAWErN1Yz2vxysLFm0gDaS6uNlw3YPMPY51Rp93hzA09Sa
1+dNe5I4BWvnXwBta1+zyP7VGZGjeqNn+32i6phlp8bDF938jdOdZ4q8mwOk12r+
U3lnc1DZXsvjQRM3DxDCeNZZt1Crqy/2E3fbuGqdwfXarMXHIna6dhbXnrEKTUBo
JS9uvnbTIf9TxyLehIqliFOCtk4DB3vC2vZrqxP7mWEBwyS8BqaF0giuJFwGA72q
tZYNiobJopXc097NF7D3DvFqKR0568oQ7vi+9aYGrjiDb5/X4U/4Tn+JIzThcvZ9
wx+NgbhXHLdipHFei9c9zsaocFReuDk1dbTqLivcK0X6M5KChJo7lNnNMrq7AtBj
D99HTwmGVJLSVLeCpiYP/7atunH3oDQVM+uuqW3FrYsj4GAz0MNIG3u7QhGUW4DA
alaoBJH0Zr/Pb3jAkd6I9j1PmK1a1sYyXMRn7s9DLFRd+5mro+C5pKR3xPEy2Tq+
qLV3SjzaH9PSm20Zl197fkT71v5vmT0XDIn87Go5W89Sjw5ovB6frFb7Tcci01Rl
d6X9p25MWzskecwn/tIOrfs4GQ3owweW/m/X77P8z6RjGwy0mf076qBmYQhwZukL
WB/5uRDlHDXDYMXphxCBK3Rwm3hdzRrbTo2q++RHFPljz0hP/0gJmlwxdrP2v/om
sXPw61MwkNzPpk+qVGyq/OjcT7TxPHWeBWTOZjTjTSdSrjx5w3mXDW/nNEK5Fpy4
pFkotPJYGzSOL0O8us2PvYdqTuIDIg0U4DlDZy2yQlYf2dipui1nZxMMyVzvp0N5
Vjr5EysgjivFVlwf+59JZnTFzzRL0zVfdHqpY6j/laqomXFdDKkjY9L4sls/ML+R
O37pDYqxIue/wg8+vkfL9YHwFE246aQSlPhPTvczgpXEjR7hos2ByCkAh59insR1
q+msF8izAYqchfkV7hNLNf2epZFYo74C8GNOf0GYqM2wKpTH3pI7CclWcISWrPea
5pVIlT6PphSVr6EKnioYBHo0is1e3aT0bYJArphOPsoPZE6ja4kBohU+oW+Wcjzv
hr0se/R19b7qz3/F9+o2fYo0KyunGAE4s1KGLEsmw9x2ZHQ0Mzk/d7noIe7kJTdP
Lge/TVgIXkQoFiOqbUYgYF59Jm9zFhR8Bg26mZTe98iz6yb8XwobN4t1tT3gXaRD
NpaMAcPuZM7ZXt449lZtXIDk/ErYiv5Q9FMMRE5KiI9aEt+UGCW3qg0wB6C5jUaN
n/NjyDbBFpJo5Jxtv+5v5NK8Qi+Yq+9Kwj5RSG3o/B5MNjs/StK4njA9VOIs6dYc
77qbZopBaxGy66iQLf4l/YBOB20ohrWRhemsgGNnoMzqDQf5YgmFwH6otnpHZJSE
lpkHgVrqNOpz9MSF4hn4P1jnoqpvoQG0bApZQc5sRkcvtbDX+blIpkdamw7OTd28
GFYrj/bNNZyLoaiSAHRMy5+ZWamQ6XdoQqXRd9MmMZJ+d2H6LGY7W3Z2alpgHgT4
+fg8mSf1B7SSk43qn9yyomYXkr3cPWa3q6LuB/W8lHukRP+6OrFJXIPF6eZnOrT4
bx3rrSLyVcDQI7JZjMwwlCn6wb4lAcC6zD171JKu5bg3Y1VYG2IIlGtXCGzEJ+MN
nDzTe8U6Z2K+/omeFTaKbFYWpKRzqLsWWnn+lmsxT8tEkxn6MLeVlSEuZ23dnaiQ
AgzOiF3p7c/351Fqq5neQM/PpJhAp0dKrnfWIlzfHxswisdMYwwF8J9e4UKbkkR2
efBYop36JWCqjuGv69Lg+Tm1LeY2smsxVWO4y4FdW/fCqtXqcLlUFgztqVvONo4W
67z+nW/4vG3u+jfHcG10Cp4r7CUzoTtM2pYBcsUwy1FiDMk6t3KmInVRkpc8fAqe
eFLaxjKwx+OW8Q8BKh4rChTGxZNIx+MvU4o440/2ha5etUTd6F/N4dcdmtFe+OYK
naqS0ITgMHn/GmMs14wYstirHTpBVvcfOB41UPAu8zAaVaHEZI9TYRBccjBVolex
ie6sNUHCZ4MXF9ZJ2csN22eY9emKFpqJI8D9v6JhHtjBaqQ8Ucah8yDm+5fnY1aG
+X+9ZmDsw7L/5jo+OSrDMDJbtoLSANdF833uH9ogL6W10yOg3wUUMvgyaq2pG2c0
gzjEtfsnfW6C3iEVyHxtHPSbf03DQzsgNJ2XQNdQIfOV4TGQoJ+8Vjw+tEW6Nfqm
yonzp0Kxhdx4Dxpj/QM1rGqZUvO9mVuUWF9ULFwW3pYSoNY1WO7Ih9RLNuBGY3lq
tDrg+3UltE5G6BybuNeS1ofC0ozORi8LZYgCrs0ijQP+bYdyn+6uCxyokf/Gf0W6
lAOpvNPPf+OOD0qoW6lb8z66GpT9P8A/XmxIKXe1yqQbFX7sZkVOxbfaF+sftwWr
MRllPqt4n8YertQV1PuBzX1wRIONX4yRn/sZAS/gJUfPcLwVA+jIo2xP5LZrg0UI
Z3SkhYT5xyy9/DPr8K6buvtUr+hUNdtS88od74yWVyuquKLxGDHhzu6epbPVtdz4
YkxmEixTHIbngxZ+PYcQFZAZP5N9lPEDICtnzEAmqw68pkHpkAfJoiKkWwqvnTV9
lHHN8RZOCvSk0+k1aEjCAPFDqKcT1dyU6ixpAGn7cIJPDNePeVf/sUXtp5dTxnyC
FFZqCNdn7g/ilT/4Vdu0fxUVANIshfPPP2GrXl6RGs0xBLAMyhlEb6sfmODysoUU
0rh38j3wwxfFGrnzAK9S9tEeqzd1E3Ojgod5RAueNu/a4e+/2C7PjxWfsdLoIfnN
ParPyfcxwcPUu4iuat9P7L/mWcHsuZsMjxUhVf0pSAFimuvH3UQpNp8zZG1a476r
CpFBZR7EXIuZLc/eWKNbrZukbzxs6XG75UX/U8tA6LXN3EexA8DbhiBORLLLNYcm
v2H/7v7ge3AlpFiZdurD2DqauXMggSR2+Op8T3Y9nm0jm8WOIT+MosHeHdbF79u1
I5w8cZx0/EvkNxQSBIlBNfSuSmzlT/0yHSMcp8KWb6Uaeqmfz6SzN+FwkAjJpg5y
mEPpo+npkzIE/LowACuIissiONcZjAl18YTJgkTPRPvgsspvpXtTrO71s3EdF+DK
AEVyRmxdDvMpYmZUQf+KTLlsn65gamE7roRi/9yxrQxFoQZF1gMkzi+x1gtCqKFd
bfqkHAQNVxmXmnOgWV7sV2pJ3SGS6WfxlvCWPRGERuNwBRxJHFcdLgzheTkxuqkK
5BiUx7NqFXNR2LPERCNjlxT+4+uVsIAPlDSp8YL7lN3o8X7g9lyUY2uXSkSezOGR
i5VLZxQzNoWNFmKCEygpKPmUhgxnWM600Z+/TZaDk6UhnvgJHZjzrPN+jq4LKYHA
sW49X/ZbcdBrczkOtdP6ACGqhMTRALrlOv2LLBbzZcxzfMkBN2JQBoGLztIe6HNo
PPrGpNSRyhasl+qkGbmtvfOlVemo8m3utFXBUkFAiNw9NMqzt1j89qBI9ecZ9nyq
gK4Xvewc12UDghmUiJ1D0EJ2qPCnrfswrIZy2cRd9xDiwSbFIOfRVmp6fAs8gNI5
8KCSt4H1KLPiJvT0vfRYMdL7w3TF0u7kSAcBVZVWDVJLeKHtl/APp5FA+S0nGnUe
zzYPF2+IkVRRpfqSu2039I12xySLl8IVXC7lakULrr4TN9vJ50n7rdlx+670iJww
nw24LUN6gErWOJQ7PatpKDUU7LR7C4QUYO85DqwmaTjqQE/sztZkmvuxHwoLgsrp
N7NLotMezzpikU2jTm2kckZIG9tfaxjsCP4+hwfs0thCeTZR0kXzjm9QzkNExJ5U
++Si5plHmb6O7FyGqLAz/u3nZ42DHpa958L+TLWUK/T5Byzf26a9Xu5pRE9PCWPu
M1s7O6UWVdVByhlt+eRVeMMuRPb16ASaM0VXZwZSnZt2NozQLzcKKFBxnJ9V8m/J
BvnhaABYmAU1V7JzGSoA2ujJqH4TwqJtZ6OebfQRJUcojyiTGejET1oZ9Y+Ywt3z
jYmk05E4bcc4n4ibxvTTCEvYXSleHZZSq29v59DJoce4JEHjSHIPGJdydedTAG+/
sHtuFkaVLD6gWjSwz9VLvrWKqZh9BsfHKL5rqvAEb/oXSppQma9ZqdvxbwIfZa7n
Nkimk6H4FK8l6g9oSDNPe6MjClmYErDbfdr9l9R9NTysN7BGILgcV+k+4mqzz+RQ
QXj5E5N+I3hxnn073+sms1Hi7oBRiUAOpzGYqjfgoGjW8hALKmtum+WWY/A9y7AO
OxUfhBnF2JJBBq9KvDYNYQMm4USYPMnPFBktkER+3gNeA9H3zFpMchkW9XqFixA+
zAymizQPF4gsDsrVff+vGix+TPBsKZFjFR6w4ugnuJn9QPggg771yEp+/ktGfDWv
uXtThvybZ8aEPP8+U7vCYeDUMf5IvVlav4nmd+jSzAvOmfF9CsmOYsE6jX3g/7Jp
V5DpB5HomhM1xjKRqpF7CWn87rrzc9urNn+tBu5TCMOvVgIGXshEPfFvp/2gzmXi
M6JClG1A+9gAlW4WAoatKEehj1ascPvxhyIfX/l0r+sK2K1hCZBGSW4KhjRs2vf0
NBagt73/Mu9FbYzPD3ieokSthghIHxim8ePPf0ujPHbZWcpYb/+/eJ1H0xdvLzca
i4T/KckxWLSE1DzuU05rFID57LF+HheToXcAt8TgfVo6Ov3VGkt6NIthY9b39UIl
LvtYmdTj9nf8IrmCn02A4gT6c+Qoarff840gtYk0ExbZYcPEPD4LjYC0GFjkDWT4
LiHw7ZlSdHrYuBhntpZEYzg0uNVus1Z5c4wAZD9rb17GS6E3CgCoeg1Y+is55+uY
KyyYlpOXjWV8e4foV21rDHHzxU15mgmib+dEHxVX3VgbvywQ29BYjlt8fo5GE5y1
NmQjWF+P+vZu4fTWBH56WN2sgaSeVrNN/aY4AUrLnn3dZYta+lAR+qD7sy33SakX
Zq3z5PerPhgLzzV6DUzXn/6z4/QLBK4a67orGuJPyAmV1w6X6ppamsUNwMA101K2
GqS5jRpU8Hlxf2Cg/Q2R3AaYyvJAk6zQjELJU+3DMHd4nvIBKW76dl4a8P0c4a6j
AK2lR+Ibl9xg5UI7P77OlcpzGPd6lVwcKGNJrj3OkP0LWTd4HPVhyyMVIY0ym8y3
H0zLYVeSxCn7mSqD0pdTX6UwkiACANc+lrUG0ZurnoVVDz7TU25VJgExi5d46Xn2
50gk9/FDmgF8XClicVt/qeB2YHXKmVtgexe45BV1+Zp/NRimj8pcMl5GBNyOCw+n
it9c/IUzq9eGkrz9OTxYureBGLE8fzOCbFQ2vBEoKZIpyc3mv0ZBXV0xSKpsrABd
Aewis3auB9u8qTnA2J3l8t18BCFhXzXZHU7Qi4YUAa6w0PxuLIfFR7x+1JmwKBrg
kBdl0gy38Dl0qCOjnRfQx6EEC9qcYc8eXEqNeg1m210Xa7l5PT2SaU4wKVoV2x9D
DD1dvYFgkyTOixVS/EgH54/uhVFj9oKl5f6UST/unXQjgnhd2gECr903tFa01vJI
gYzo1yU1r/FWXHDdvv3lMTrGaL5ErnXxgCtTpCVI8Zgoma4Z+u5+uXSSB46fWEbg
i+CSFCKTqtI3daUFj/kja/pf08ryTot1n3CLTHIT8v56GFJDwyS0g28DbF+8WNUj
TzgSPB1E1WlBT9HgUvx0kuS0ZahuohXQ9o7tpKiYLej7EgQBwJaFA3QQz0+X6U2Q
t4pkB8HdGrdbQVslFZAevflScFvuyLYT2sEe3qyBBFcugSbF2GtbhX6wlWrBSEIn
/sq+cKvNPNiYrN+WJZ/xn1mMHnA6+yPSk26eDZYC2LQ3lkrPp2L22zIu++2q1LeC
7j2uUmgrp5M301c15pHGn9G+K3zYByWEWkn0csuz/AQQ8O6OsqghxsOpMZEZ5kuR
RCQS9VbRC2PLvzFDkddVEukDTasBw+1LxhzigmFKcWfrd7XiIWtxbfUMFHTUfgdx
y9kk6vf5AOICa8pPj3xPcahHl7PINfeP2GwK7JSHIH+xR+xYyjVYfw/KOiXUqU27
LrlijYhxwUqSSk4qZnYfHZdFGeS5CbbQZg+9eyFp98s+pSH2vzBLYfdY7FzUQHNi
r9Vpqv9g504hXxo3nNOm7AJ5P222RduXFuhrIDy5aayqhI370cCoBJOpf3A2893O
EuuJQh2T6eSU4HaUIk5gy4nBmc7rTfIz7YN23EOeyCvd9TB3Zn2BS0oiOAuQvPS4
X1MWgC00JxKrOMuavrfluBBMLsHbLjsWElauDZ5XkJ2qiu4hQtFtLBVxeFaU/d5b
T/1FPRKtc+KZLPhhrk2zVewGzk1VI3F/jkzNJCgH5WdQZ3QFwCmVc7ZRcDJ/q53O
gGA7XraVl6RwgPupXr+EddRs0sJSFvYjft/cqrVTpoyNVGCt9XuCC/MwbZEnqJuc
w7xRtn95KbQSN3jTVmcP/FplbtTI2GwLiBq/6+cNCmM0Lqs/XU4dAIn69+yvDkHm
dxmhS+7rRwsiOOPNX+hfoA7gU3tideTLKW1PngdmOuNkfwkwOFQKq0BtWlgtAphq
Z8KKRaFxRyGBxzc06BNgw26+LuYPq9iEf8l2x23LliFvc+/kQu/pHGepz4+bTHNA
fLn44ZDlHpIRdB0PmjwrxbKYyGszpvCzu4yrUj0CLu2bG++dJHuDif4QHZNeQ6We
FEPuzCiOcwWhgAmuisI7car8IdWbF9k1tYAhQEQxhKKdiNUJC407U7uIBDZZ/1e9
dw93rtNDVqa+UkuLYS4b3ihQXwFYajvquyeCsZVq5CY9bDRbH6DxHOaN8aC0PdZm
sO0gZmNMTeRg0689Vc017YjDomdAXbMM96Sl+3mgG2Sq25kaydaS8oyv+Vry0I/P
NmzadDyLkqGyV6tGcerUKsuFnXUrzNdDyplTaFpw9DN/Hp9ncajdQgq9mwDwC3xt
YS09RuHj/0+nuXA7VcUch5M3Q5EAyAcuQ7kMMET0YwXJxlRkyeZGWyQEwfHJy0k1
THi/uilQNQbvv23CcGxpJwDd1DLPTkxh3YgyLtgkCTSemtA630ZNmEkSsQShkP6r
eQn5QmtuTWG91DrI5qiuGh7oH4MYZtRRkQiwjoxXOjyNocJsKJSS4E56MQcjTh9p
K6c7yCGAIWVoxDAksoOk9DKH3p4Raf0cUnM2Rqy+QpheZ4800ek0uKKiS4NSgmgM
4bpV75IzZxm499RENBy7DZJiH7NoxKLHFipV1V7HOXIRVwO5SYM83I0zIdylZWdH
biriQ5ll8tanQxx4++G9eW/5IohAgUnoVdCtKbZxiLAPWBToaLApVtKuOJkw2FH8
/pALYcKYhwihB62ssWhVVoqZ2Q27owDHgW4TMAlYblZNDcajDsmAHaNDT8u52LTZ
F3B+3kBbFc7Ik/hMdWeEB+/2LG82msPGItyuw9Z+fTWe4Ep/4BYcpJa/rwHtBHHG
B/XBu0DzKWqcp/7h9JJaNi+b4YWCtzjhXN691aSMXsxKfYlAuokZE7V/v2pbuEhh
/YmzLRSgnrb4DyllgA/0USdsu6XOFS7PFLcTt9pdBWEdeeuJsgB0EqHev6QySQ98
IkDzKSibIP9seK5WjZN1gyA+0cvoUwQEdBTGlXrFSS7C5X0qNczMKp3uyr9CYUTG
pELPkumlwJ09KxwvTn1ybgeXS//JfekQhDnLstSom7qQaSA+CTFe7XYxOdHIetlU
+8VuDiJUXWELETkl34PRKbI03DBv3z+eRT8/3UBmVF9+XbyuQBuahjNrjMtoIAPh
pGtxoBfhVT3WMTz04ITp2hb2huODwNnShLH1xvgsqgX+I6KT5ekT/ZdVvdSPqUsG
jS47Jq6APTVAYsMV3qGdMRtQ1h+odaNokvrBgm5U9anotrmusbbsnHE1mANxYC2C
TxWsfqWj7LxjG2NanxxNPd4eMHAohPUx52fhd//U6ga4n7jXiQz/PyhExE7IwG7S
akfl1es9aikweT+sSTfa6cc/cvCEh+lm5Hi49zh+aTvfUnAUkAl+1vnReqLVVGmn
YRZQzPnWnWnfsITJLdS20jU1VYrRVoGxZNuhiNVFCG4+xfbWsw1Hatzrcziwnaz6
TI8CEYDQ7ww7wGXeroBLhTp+fLzq7mfpwhEIYt/NIzVdcuOpa4cte57JQ2w9+u7D
DLO+secaO7aYmVmtgeqrY8xbx8imrGhCmYAxZl7l/fEZYRZVoZhrjTtrXQ9hyNPb
Ry63J9SzxRuiGNleLuqjNkkfspoSiHJGiN+uQKZRxw+Uhx8Ne25HMsCzoi+86MoU
lOCHCgXyfMAVwos0jJHlbzQ2/TDLR1dHnuKZAh6mifv61hTD8WLI9iew0VnZtZVm
OhYS9Jnu5bFUl5uUcs/WQdIM5MDb5rx8kcL8N9A5kgOKQNxRr0YDrSOPe4rgd9AK
ew8huF9a0JvF6bZ61WanmKHA28emJuCYgVfr5Qf2v7POeTfDOFpqtBaJygwyMnri
OYLbqRltcn3DYX8aS2nf3Nsnt0u1V4GhTILA6uHFuUu5Cu2isT9Jxen2fwljF5iz
EKQEQgUfH3SYdwzIWnQu01AZV1085Lsi3cH6w8GbrIQ+tSOhPu+cxckexPpoDgHO
STVutivepVFsUSCg0giblTYnthgvREGLHYuL7M27OQs7GdV/6M/iRvscJRKEOlDM
x87csvMkE+h6rCejS6j5zA3SV9DyrmKinYwvBh/VREleDNvhNhQUWdHWON9U5A3q
t0xPM7nPB6O8KqEzVzeKFN72sm8+XeZ8Oad5zo1vmAoENM5SfQq9XU0DCqo1kPQ3

`pragma protect end_protected
