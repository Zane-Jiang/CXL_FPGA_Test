// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MjTaLWdW2Zfz30FnjtGpz9jqD5Wr47bmHW+In/ep4NE562RaVgfzdVCH3iMu
DxH3r8K+B6UBKKNiVQnKmJydegyWFzP6QFDlpDVqd6EcW8bmuQub7S00Eqol
4ssT8wvMZxbO4nZEihHEW4NEPvgkk9B+/EaUt1c3t7Tjb8mZajZH6aHvse5D
QPZ8RjcXwNZuGBehjFc/Pfe+4mdH12I2nM4+RfvPELeT3xpxWuquP2OttPCO
JEH3Bx91mYgSI/YyEcfXwUgG0LAp8VWP5KMtAv5f+dJB4zNvqNZUH1Kx7Uoz
0wInKhAdhPwaZhWLsmf0InoBfyABOcdFvUBamqRjfA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AX2aWDyuBdqJO0VU4/XqSdG8zy8J/pU3S9L8ID0aEfuAVwtL2QnFaWebjh2W
tnrkKOpmkMLuIKidftWDMLr8uHuadM4OoITzfAn6ixjwJVQVNcP3yB89vYNk
iujqHD3tAOD0YxVK8dtWl/wIzfOjChhJ6hma8/SjEtQds3xlJ+OndJMZf5c+
pXO7lplG7sza9ts9fndcYAejPbWzwzfNlr005JIL9D08iNocOBjQ0T+YiwUM
HsETytQMCqsqVGBpZFkPcah/txiaWmJAwJD++riwpM2+uY154AobAdoBQ2RA
0BOjkyZ+6fYd/dq+72KdzT5pc5E51MPDHgH6sgMHvg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJAy2/87iBOPrly7TTfMovtZSEj6b6i0fHSxCkIgQqb7zW5xT7juO+LanmCB
2+U2TNURJJAvuokE6vbJeXBQuJkmDmdp+YtGwtichaQPJU3jlwA1ZGTj2v9o
ZZaJ4pBgeDPVuU/RFkEeOEqDeLVZnm7fEeO0NY+Uru6h34QYmVaaNbc7o6iZ
yjKLswK8M7SvKcu66b/ro40B0fo9oVbEhwK99WGeLWrWYaYQ4k1S/zv/AFYo
86f6RRSIjyS4Mv4AW4FHaK8nUjjbPEQoS+adg9eFEg0UJ7l/JxIZib7pb0O4
IeB0L59Yy1SRzh3LkvXmJZArvNNGEahBleEbaagbxQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IqTPzqcU7u8GCPDTHfS2oNy0+13AV7GI0fxMfSaC6Yi2ouze/O8sLIlXJJHX
FJ2xBwqbmt8jPyJugYO58hVl39QCzH1/PDK10Olib7yiP1RNAfPCkBRgWrDs
7BTO94dpF0t+UwiVBAXIsbYa2jYNS65EQEGTYQx+645rHH6doaA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LN/fG9P4y+u7NTcQ7+5V40KrhYm1mfXfOzW7fjWbMFok6SxuH7732h8m/cgB
nXrYI7h/DnJWf8S8UrP3wUXSiF+A6ANUacSGeuXjtnSvM2QyE1ZG+SkfJcSv
7v0nwFyay2IiaH+x3dth1DfCge2oIfQ7rqd0CW8sNwNCfaVDydNZZgvpLF/B
tIA5tJOhovsah+obU7HrSnWOYZftnQggNHltWGDwqy12ThOApPMca33hzkI+
6Rn6OqlkgdaUE9DXxvDOI/VLoockUYfXmtY3TmtUoVX5FGpzrIaGRulqp6RC
eszNK69/jQ/jdxHslYLXjrFF/KsY2iMb/cu8RxWDKffzmorY4troVjr+lG0r
riktdMK8T2cf/7LXk04okNKc6s+HqUqcP5lYwXKAQUKH0S9VP2++WwIrLxqR
rR6WbfoYcOJviJxWvXBDaCpnPJkMrRAW08t9GqmJKjxx76CiW1eNFhm48/Py
OjLbwBDz2frgD2QmdddfvdA2rIzBqrbP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oe2Rgue9r/gtMmNDxtB8JEJCyne8nFbwU2KI2EqNzEfc8B9uNmE3g3Co70Wz
R2Ji9nKbZmX8HjPX8yxv1IDsz/RhQ/Pfcn8xftcfO7I+qn7js92vJisoY5Wk
Y+gOU2m/btEtHHadb3BhlcSBkNriRvvcE2bXwF9VBXx9MxMkkBs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sB+mrstvM+eSJLyf8SBZBJhEgY5sH/pR2kHClU6eDSjtb0TSNZCPGJuZaDB0
VWXkYyDDoY+x/UnXFmdIKjzqznDpY47bGZHcfWkmwy8vNejFV81jPJ4pnKHX
p4Jq0eBxJJeU6hfWq9n+FZ3L3MX/Z+PkIRHXDjGvHnC1s0TWzHw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4064)
`pragma protect data_block
98/i7vmpattMTHxr/9Acvi6AsYPa0XjORWK1XEGj285L6w9kUp30g53RjBYT
TPBXtVZmNAlxEq01NVmeQIUqAO7bfuG+hrkUkUCAcBtJCQwOBfq67Rmk8FJc
v9ymuuAGznqt4YvQtKYslGFVNoCs0RDDareRoFGYGX23pyVF3H4kRNhQS2GO
ixGOw//tIVE/7LvuT9ahjJxclLCyD0DJQouO4jRcxnP4V/ldj3IWCqnFjXJ0
CYs8kZCxb0mR8ZBGSTsf3ncXrLL/54G+MWep7AJuJjNQ0rQwI4JrVZZNS8+6
dO2TP3lM2HYxX0R8xSlJPF7fC0krst+DBf8VS0Eg6bbtyBKgOQcEzHMO3qJP
EBwLmFuhJjmjWpTAnwp7kFndvh17atcHjMaT4M+EKDclvLUbS1UUOfwIFkW5
+HaJR5ePlipGzKmOhOZGNIjhwGx7V/GlixxC7EzyuMYoGWFgSync820Fq7Xb
RxyHevo0KPcS5xfaGdH7CgXQrFhLfmEr+UHc+xSC2a4v4+pmtPkYo2TiPhY2
xvsAriqyUi1/rKWb1Y0Gcn1kqk90ylxnLp9moqUR3oibbEBKDqjdy6FSSgqf
X1KepsxuQqoqGgjTUS/IVOYR027FWrzcRRZ6rb5WTKpDCzARaRetMuJdavv6
VY/fc6fNj3YZMkopBojPm3N9Pl6E/d4OfW3+0ijFUQUn009Q6y9vNRW137nx
maKNZhoVptJjoF/ptT1/w7KWzu6FNAPg3SGD030fuQWRO/4AeeKZNgfjLFd3
aggdNfNAp0VZLbUIBPpFbSUHFNxk6CnjorsLxWLxaOq9wIy0uP7VQtTWBjgO
UzFK89ku4IyR5E4Gcq0Pw1RRoIvJ3gv+egr99zWebzLkXKPIq9mYm9HpCiEg
Rl5szYN0lMgeu5lG95zPUOKMJ0OlA9yuNesDpcMRZn2r6AOVBkl8HfsdJWlh
cBzd2CBDwKzSE7XTAPjHAoJ9OMBJGBQ5I19vr/+LuzsX63OnefEde+g25I7R
qYRh/NWB1R791xrL9Yq7qEGkhDEHgzucjx9GF/ovso8jPL3G3LEP15yMruMG
kpg55JCWlr2zr/uPlLn/xYXI7uRnmlp7Cymg5tC0wo2H4/WwnZkAWmxW8AxT
3n0V4ibqRxZHU4TDHxsCPYpRJhMP3lST4L7xKfZmZeMMNr0ZpGTW7fdqwnrz
HHwCm1aBknn4pFDsM0st+DjstBZIdB3hKYDt26UmbsHHicP0D1G3Asc2aYJL
6n3KH8fTJxpy4vW7aOmKQf7AxnKkxd396VfcvVBmt0zhv8OrLzPXW2fmpsv4
5naU8fqaZWWBFqy0GVeWsGZLaKb9Nxi/sgJtD1LwdMnk/jIPHmPXn4oz8EWR
alorL2DnwbUurN1iqD3rHlXMxKkMEqdpS6LoJykK4gbz19ibHovVy9/Utc+W
yRZkv0fgmAEidOzp33QmhwboYXTr2yRzceeWAxADlG8PPqGtiE1Jqpjg3vhh
LdkIgrJXFdC1Ks7qTtkjWGOQ86e2AuViXb3MtD0hQhJjFBMuEJbkaF+fF8m9
v1B9DnRyBJ7BjTLiKJkDWBXnnUDpIt/B5zWzEcs4PI6GE2HTvUZJVLDfrvRE
VKBJ2S27k+qkCOyNpyMjJXs2gSlksM1RpIOEkmLC9pdyGmuN+lZrir8Qvx1v
G4qkGp7SXtHU4K+HqL05vcVIOWF7AULlEqfX3m4GEBjlw1pQNT7KTm8F/fiy
GQuLEZzxDeYB+hOdBHa1qje/pjclrlzsNldVmAJEHulkkm0IrxDQRVwI7x0A
JUc/6b0OJTtCjYMZeFXPbTt0/+vFay5mU1wV20u3IXUaKUbu+fMxnqkEDg2P
BznGxmhOuv/XpkXFaYasrpH8L1RnDFBxgeLerpr+yNDd2olfLs/5FxqGAuVk
TzeQlcnUbYbV8+n7oBkbtDxmXNqgk+tHJOWH/fCZx0ISaVMqUa/3PxBe+mEP
lauvo3IMWPJCYEPtfVXTeEtohdR5xJu0Y+MwRbEgIRgacs0PJlW2lzGVUZqQ
2aqCh5kNTW5CLUVm03JCytRtj+B+1ef6EUWxToPb6zUg4Ufa6oNNvmqNrEHC
tCs6dNsIeBYf/V7MjnALNftNh7KgXZiBpePrtNqeuiM3kSKJASC7AM8v12Zg
+0rj/pxv9JhcD1RhKTNYPhq7utmuUF31UGxAZ6w9BX5vz5cmp/208Db5L7XL
2VVAu5EAw5nBtW+QsCrUKYQslBAWmOPSEMGxxt0atWAaVy2L4hotJIcdsrbn
Qszs21V7NFaNeboqnpOYaE69COLTWXTHCJRrZ2yCRwUgF7odMoU/jpKtqBqu
g631EhqiaSksjI9MbaqCyMXfLvTk4BZZyPtz19S/P7sJ6rkJ85EpIrEJj4bs
2nTWXRUqYMmwAWH8fBQ3SNlwP8jUgMMEGRPw+oCUseZltKX+KWeb8wZPRquq
uXb/RqjujvjDWkC4SgqxagqvvJ1iohHzK/7SmikeLoEWOKFyeGJnogK0gVqY
y6z6kfwt5wXqeGLaA/+hOquM4Zrq1eETzvtJn2RTZ/B6EjLghHoz6umkpspe
AkA42lZHnNN99+cAb+tOCTikhDsoH/L1LLbOz/mgC71rsB+bBS7Ifs1iDd6K
rSqJaOdS0EfolK7xkn1172HAobBCMPf+9Be66eI+0JvXU980X6h7R3pVLivO
2G+zhJDfTJnZW9rCvkNP0reZnsiKs5VMfHiv7OBpDdKHfc8C/NFeu3hfHKKZ
ptl2PAZKbSxYqj4okRFNsEHj5RrkQVxBR3FbL2SwRhHxhomCC4/qQkhWOZIP
blOGlkpIAN+vLEup53fKyPZ9u8xaLstNwMBrtCI2eXZdNRah/8itlUErg7ai
MfL1aeGlSPBx6Lzetf128zgsBwcYvjc8EEn+APWUOfDMfyj/dVMqy/VOK+TD
Di/NoPC096MM6VfJGugigAhciOcdKpSDl+0kXsSeWfCpBvoqMHHYN/uHDgFX
hIrgX39NVAPiZREXNRiy9xSXGvBfnGyyNXyJNikilk+Lb9wStLQrN07wk7O+
O1U63eGe3XxdpTz+XRzCGz5C/oFMmN8hTb43qFrArVZBmgF7vLiPK8fYUskR
/tg51PHimKszDREgh5Ybv2m6KxUTyq7cgJy4PM46VwCvlUnTwToDXx6vMV/H
qjy+AKONlnP5HIsYlGV9Itnv2Z/X2IizprVvHn2ORliGJictCmwgR9I7kwoM
62o3HQ5AwfjrhaB59/MUaho+aIN7PMcGtFRqXeGXcAmYH+tcvmWUFO+LeQBK
N2DaHjxTQskU/OWv/+0i0YZvuQG2mxZ0Pj6faJ4JtvVYbOjbPmcg3lcCGVVJ
CrsuKuX8x3iyYB4AnEvWOnR2uuHSavpXGeETP4HLaQdH4EkZedKtmWteTRwI
QB9IHl3ieErZeG12PA+MIOK5u8KTguanoOZra7ps+RUlhqjtoKep7XqXD4yy
q+/ZfCIetzU5khFsVuRWPiU7u/K57WPVVO6bOru/z6TdlEd1sYYvHJDpVRQX
InyafU8vkBC5tVv/GqUQTYseE//pJeNXclLtVPVbg/2tYXmHWnDbtsJ+qMTS
awQ7w/h+qkT9Fcq4NSTktUSye5hYOM3rfrojqWKioKFCHdqz0SG3Ooib5aaM
qgkUVfot/PJEOpH92LIV8MJSKQ5TjhFu6dpO80jarppGI+LEJ29apb5euQ4u
ZREmRdEPaXbrEH/cfRHXFNbbBaQWcNXoedxlz5C+8GXhotOJxo0TniYl+8kA
TKYRJ2lgo0XMrz3JVt6G6cd/Y0/n9mEpopkCu6ezXAjnsO/lC0mjbsuK1iAa
OTyxHuevREVsRfHZINteGAHEqd8M88VQTVpDgCJxhmfqSjAO+bqa9kZnh7Bg
LQIUL2VJNqrAqzGlxvbYon+tao9CdqgW9uU2qn0l1YmDFvjG4HubsU5irtEB
HYd8AOrKzhp9SvI1KzHb8+bM6QX0pMK+GL3B4+QOedTp3TcDID9nfTLHSVCq
QyCMVluppCgAGh/RQgpEP15hJBvkNfB6/FGTxDAE+OKpd3aT06Ez/26qmSF5
TNv/+KlRy0FYmPhSUHbA76cJDI4Gxyv4PcugRICpDgRJKa/pMo06HJbn4ytp
e4FC0L5rVAz5oV9sckwIk2HDS6XfW0zmSZdznGs93hR0dvizHBve0XxU4usO
/hDPXtnGP3jFAEM+aWUOY/Rh6p/DzdcL0W6bQii23YVRdwbfET7FzGJrQV2e
ziXZlARYDQsZgi42dpihxH05hz7h317MRZpQR/UmvnrvDaMR8aDLAEMzMzt/
geESiSzis2ShJtXA+CTQCjZ/yM6/3KF92nFTlu2T5fc+lXXhLOgpfY3wjLxJ
l0UlZN70KQaFUWM2RotHAP4uNiKMkUjRivoXgDZl4XA5d5f9eJ2+qlp7xKPD
IUPeeXLv8FkcV4e9h94ttk1841pBk8QzOqIxtx4szP21sQ8NDrvXkA+mo2S1
MCRJswhn5j7+xLXRD18NY9xSNoUl7uwqR/GGGYvBnY9aPU9lvb/2uRDN6OyJ
c+2IR71YDh1orTlHFSDL6nmJGSEqLyIzVY9rtCiuItaPm509gEN/2snO+n02
BCWCSwdnxofwAhljF0yfRAzFthS+nVU9Mndf1tYRviX4JJ1GD6J1TsMz7fQe
voYQhh+9X97n60q/uYStZieaGJ58iaHAuHDujA81vSHIXgaBIyN5bdx3wLdW
58ChVBh+YvsVjFtPbiRRCM44Jmk08vI6DWCBDHI9JltQUb0+3vxmAUW/4NVH
4AwO42Hc7coZv7g9JLdrhq9ZuxX5hYiOYRydn1nD1CsAi9j+yhtaUakEXFPT
hdZsE7teHy9g+AewoTUeMxVIaOanvyR4xPD41585fNWiF+B1FP4SjHN+AxpB
6BV9OAbRKB7O1jsQaBo2z/7WYx7q2277KeWN8+orhoPzp1RL61pgcieKk4xp
2tzzx1LYGKmWdfIOtNBJ7ax7bUeTZ7mqc0FaQ20qUhLDmOTjq5bes8J5a/fk
MGVknTB3sRc06CqhX5dYEhsh2mBkmXgtVERvrHavZ8pykI0k/630JR4Vwyq9
wzZzLkqbpv+56pibQNxMkGvq32ejBWftTZZRtN/0OEYhdZuGNUyVlIGL87Yr
1QgZP4+Wz7IXdzDvRTOsqfxDjk4whG92LSszpxNEnsQ/Z5OmgYFqPjCnvpvH
BkLRtWiKtzqzg9AG5+C5g1imZ/cSfMSvBuTT/1VP0FqOUNN5afhCcOCXmWgA
pfHZFe8OxzQfIlJKCSxZffhYU1bdUlWonZcjeYAG5vpQwG3/qUGRYvShH95q
2rr3/fwv2D14vOeSX3jn1/s6bnnKnZZm4Ju924xgaFNca04J4BijivkIYDEo
dDqyG8r42OZUoGIBLAA=

`pragma protect end_protected
