// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
aayd5uchpIbfEtwbXKKKp3iOE1m4ekC/mDtkl1NoBmmSCh/3qaJqNpg4o2CFEdOB72o8WqwYlmE7
Wt+dltmWT6GuuYwvvAZArWGTvjtQDpH/JICnR3/nMgZ44fvljIjMMBuTkK4g2Irg+upd9smAHlUE
a1Gu49cBs4i3f6aewoUxcQfMkusRndelicPXIeXIKOKrlKFpXuNj+NOsRAwJE5MKvArhlzulDwwD
Qp3jJJ+wvv7j6wLhRNZcN+1fDN3k2HQzEdLMxSN0JUsTxhkWXlT9E3sxu1JpBYEyZwqusXEuofmT
68z9xY2yCTf51IAfvfPZC1K5A8C7zqqQ1A7DxQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 50208)
tIm+M6gs08cOfOivLtXfNpeGvcsEoPkfctvrY1fwGamn8ezlwQo2V7b11GGuCRR8FpHo0cjHnZGy
GKBpjXOg2jCYgED7YsyMIgnCCjbCY31dBBZl0fH0/YpwzIlxs92S2+8h+VX21eeSUkAO3dfRqQ07
mKBCv0Tj/ApZI5MGmsjtSfdmoQuPjXTBnkO/6rACihdTlVv5El2570d5qBCEKdx+V7Iw9umIHLyk
csx6ePfEHyqx6J1vdCpN5BPocXsrpteSsPvQRdhtDluNAxnoc3fDmTzu3jjaPw6igU2/1xNbx+TF
5Aqzmn09ZRPf8wiJTaUhtJOhZN8Kq2BdQoGVLhiDcL0jlEz6Q8iCcH/tzBazJY7AIlBtM+CUS2V5
2EbqddbevnryFxIdGA425igs8SlqrPBLaSJAZmO1LWuCPlgQ6QscfCWLZLQ32TaobIgtEesEv66V
xHONVWsAPfkGWkNMZAXg15lkW55T+ABtQAp6p95bIIZbSyS4HX705+Jksrgv7aevaEWX21Ejx68h
TzGpwfNEcmWCNwN3k5bQfwdWT4xOYFkegeS2dRcBgz71wd06GIVjt/eWOWlbWMEEDsFa5xtDWVc+
Pkmv3d0PQmcx3tkkwVWZKU2FaAhm2HvRDRWx5VUUCcGHVTa61PVz1tMrr42/ZIkauFUuE/BQUcqm
61IgszYC/nfYBvCo/6GucogfR15UK5gi+9Iqp2o0/HbfB/nC10XUhqj2dQmMBYC0pm6JsGkRtpJG
HHiZcks/jneT1nsK2cO/wxlROBcE/ie2DT0+vqI5i7nM+uN8g0WmrMtqnsQwRtC7Ow+qKRpy46vf
KLSIz9YxjVELfoQSHlifhq8g45MfLpVdT7x+jFhyrMz2rgHysFzHu4FqqCa0DYlpoAn1PlivtwNC
jJ69WtDjnvwsx2YtDvbzggf7Vw+S30iONyorHg2/jQ1UBZhUfgMYlAXlRi8DeZHiDmZZ6z/iHDmE
dIVvzasIHt15BXsPAytZoMefsgLJ9HXvtPrPehaWsWvBQkIf94Z3H6Rs5fG8Qnj728g9KTL2OVAd
RsFIP+LN6Oy+ICUN/rMhoX+8J4M0FjIUNgddmAHOR/m9yNaqDmJo0FP+nBkdmqi8eSHzg9RMUnJX
PHOkhN7+qj4pHC8nRoxYz9tyVLZjXQsEknITD5Vjt2muuYHJVqOe5dnLGs2V/uRtJ6sRb5GOaYrI
T73n8vXrvt+QwNx3JtyHGVvKfMZKtoKtq0RZ4RTJng82Glg+glAKRXkW/H3/LXjTYALUnzAAVjVR
fKxV0UgOZprPWkIQKhI22FQs9+sdEr2ZpgwisQ5WPg7aGfKkqKOwmA+1aCGXAn0G+SMDvfFTQCJp
uX06h3jDWS/lYpzKsYjlYhAhx3HDJrG8IDWideDPI6sYItozmnFern/oTCfWqeoxSQaL7JTDV5RA
A3kBpaGcKW2UA2XmfRjY91tekCJOiBhrKx3SB2bY+Ei1V+iiwciATRc44aGCAaBo/ccKXI8w4VWv
DyLu7KSjgN6vl5MXdo/T4gOcK9PiSU+/3Vricr+uAEpfVJd5ZBGh+LUWMT2tEgoK0VDNGjQOWgiV
4drWHXSjc/BXIS/U4nMbrBt7c4HKpaXcLpfJA35dTdDbiTamfyhildMFTUrshHnwgd7fHdswnzmo
AHQn9i1Ot3hcjtJwX9/40Taiw+2DrvP3krNrouxxSkUP1WfTOdBDQL/pNLOXwTmQudN0EnNm0QTE
13kl9YqYj1s6RfFbX5nVBVp1grsMFbzqYgottu8OI5NBgjaDN8adQ1DGUy29qTobHGPQrHmBV4GL
iKcn+PVEwbp5KU4TFLeBhZvR1W79ImMucBMp7Pk0f5F76bS0McXe3MqHYog5ClXHaPJveFfBnf6+
dDhSEB53quAqQkLIQNfYM+q7XE6xS3t78xzjhB3uaWjammy5A5mOPPxpeUbvGnrCJ+tkHTkPPpkL
ZXubxuYwnb9rhcm/BiVX2Vwq23AaqH0hH01MfqseeuEOwnqCj8XN8JArSmYf7yK1MOvkp/6+i3HY
FBrLj29VCSqPyPiiF7aHp01MRO3xIHC3TcJyqZtMjJ+LethI1idpvkKbBc+LmHGCPzkkmRvkHrtO
LL2PYz5cnhR6SvKw6pi3KB4bJg3LWdh7lyLj5AUdbJZT5gBtyE2/MH+n2ws+tMDtDU/t0NoYFM0a
rA7y+doqX/D6mLi0EWIoW9gFqx9Z3x35/JsNjeZxK0bWZjGBFukSVuxgCRTKfzkEu/+ybL5AFqAi
hIoyCLVyUWahjkD66RWVk4a6JRHuYw7P0qTM7+r7Du2twdeWIXS1fBvHCS1TQOie1aBXy+2qoP1H
7KIRzDgVQvx3+Qd9Uu+1HSnAe2+MGYFP6Wzn6uCDlhXj8ZAQRvmnIUtOLFjhWGvtn9tB5ADhkyne
rS29xFj4UxH8OhcuJ0Tfp5UVzb+sZN+I0/hGDmNVCMGmclR0AByObez04QOzpi+ypmqy21AZJ+pL
xSljUHujUYy09fPNKSf+M3AJG39ewtrdK9FX+aPANlWhtYIbKmwPlo7+HdsayFyNjStDshEnj7J/
Eg5rcCr3SM65QNQDtpZ5gbDbRDC3u2L11E2zsLRUcw5aVPTKNittSy0oZIpe/Mkg0nhQK3x2H45r
hHia+7ZW5QzNmLxRfCLDDMTITQD/ZOD78etq12iwxfx84KigcLh4jATgxqJWQkfGWk0LFc4J/5WG
uVoSp7dSDtTbJArHHUXhdKCr1zjDLo2YTm6g6Ydh5gBsK+geGDLObqsQXy91LF1BIFNv2ibcvKU+
dxm8s1KDvFVjIXCfPhtI7fv9c5MKgRMNvFyPm9rLaOqMSn2E1ZH2ixkX9LIHOw0A+Nkr7nY4zQAf
w130+idPEf0mGUut2NCsmNS4qqVi2r2FszLbTVP3RdgYjYoqyWAJv9153m/3tc6viFoqZGsESeLg
B9w9kyBhL7eDerlNXBSNSxvt3n/iGv1xavFvtdtqkGlRWQu+g6seZv53XwJs2iM9eftMnDUQ/QZi
LVX5Hf6RSl3aD/qkZS6o3LyO+jJ29Aj51904RAljZMdl8MeEEMTMRgrEOfhIE5d/Oa2QhXK7TOUG
A49BCRPBati1w1yfgwdEjdvo7jGDQUlnmsmLmVg9a2SMbEnGqG/4LFVhCsum24XaSxYeIWQc2EcK
ZYVgqQWcWEfJuCIdpgtshPElzTxwICBp5Am4cgJw0vkH97zmq+VVbYAxklxaxWhaNuxr2AXQiu0Z
jQe3QttJPXMMxr1u6UfH8m/YJ+shxgGmGuMsAavJXq1RQ0niRIdUZ908rHv8LD21ZSSXrlaEiiU/
S0EjcuIRWbaQOqA/5WENRUMaJxzqhhirEsHQOfarleRVRVVlZOgMqJu0VaHd5YfEPaGZydG0v+oL
X52Qas4zyj/f4zpp9aVG4k7IV8CML4NYVSHZhhS4D4td8c8aaB2tmVCWAjm/pMcJk+WwuL7Coz6L
UdlWqOvdHE/BKwoN+SWM2GWO06xc7Zig3tCvfezgTznRYi1cm45hvLHEoD4GxhHOE2we/JkzjiZl
7foxz11bHFuON/bLD0JPIJFiaNpib7DIWhHCCy0apeoVELgjOFA1jtn0szZpSvvem0fHmQ+mDK97
Z9c9+aq7tac4tiRvn9HVar00KRvQBqDArIOXT6Rn+buqHu0o8wXaSqWPYKycem1W8MCiu18gesa1
FOaRdRwnbXf6nyVLJiBw3YJa72pc3EIDS2PajhH1amdpbHuHvUm/71c1djOkiLAWXXqScQ1YhFM6
7+zTA2y/1iUIicZyi/pI6vxPYeDiJ5bzV0xWkk+3+yK+Ih1gse2bR45qPCjLLF7RZSZKQHpmx/4/
hclzoA5/GFvDbQAfGSmpXhA2xxOMMrbBpdSRbfQ12D3aQyZ7YewWs6YxqQ+cbChxDfl0VC72RIzV
3H+VjMDWzl2+e87jVlWlgdVAOOggMPJdHCHQSrv7KDiS37PoEEXF8kp1dxkJkCKAvjf0LKqqt/oX
KLFCl/vVTg8K3HlPup/j6ex0go2vYNw5m36x5i21oEOIqKr3k7XsyO+HAkzu7Hj5mNB/ZqQqtuU4
S+IIJeqbWeBsx8EnyKn69DRWzH9c2qrJqgHIYTQ6i7nAMavJNF///tRrEAGBCKUrrup3lXYkWwI9
isZEe9YN7ffyzfQXhku8FrBxEHXK6+YoR6p7kL2+YkwjEKzzrQcAi09jTKNCGecDryqv/7yE328p
+NWRyJe5WmHlrtqGTa1aQ0I3pVFjjMwS0a5KkG5IM2/0oiC8kmPVA3Fv6efcvvv+ycg39D6gceab
NGVLVY9DS1fO1xFOxk0TUiyZgeKNiyaZHC2HWJrjU32VBpuL+Kf/fKeRyhr07fOI79h13DDfrnkv
TX2PXnY7PnqBfoVY4E2knW5bT2/51w9vSOMWe1HA4lABPh2Fmi3ThrA2vsUNP8+WYt2meVRm3f2U
LfLt4LicLYGV20gE5LCOzwiryEwW12Y/udCR1qDbNNARYazulTs6k55FGMLmMbDpX91fBUifb0m/
R58vXMwpZZvKGHeEUxxmyFnesjXi4i4j9cxzsifA9Wxj4gvUyd5teiP2z5r4RNKm5Zi1b7WyHHxE
SYb/QDBuHq96lV/euVgsQ6fz1xAn9Y9V9Y9wTgM4MnyDQIKHvnBZUvB860BQ2S4QqD8/3AFEglY/
OjznjJUbgghKm/TQy/7/xWATPdeX1pdE6KJWMKIxS40f3I4KOgdeocnUMGK5/PIDND7PQZFJfRhq
ccqjELk6ZonDsHfdIVRnIu8zBwAKfrYtrZjS98j+ajk1dOTfh+djTT5Jx/C1EJu1MzCqlVkIpODT
yXMHVd2TJ9sMdiFEPJFa5H/syklbtegJQljCzOYGq2dF78HYF5RDTK4ifr6KD/lB6CM8NZcEWF89
Y77nBENOSbl//EhidtB3U36mzkOBkZmgyxE/BXkosZAU5w12SwVAHFIitB7oBZ6e8plEDOJ+a8Ks
p3QKwjvQ+/xpMy/2XJKCneEvjLG3TIG8ADO0XCcXzpYt9L68qncoAOEZJ2URSKCg861OH9ZIyxpj
6AhFFRCVlOwLiWa4xCI19y45I6FQ6t+VnLN8xtVVFU3DnanUg95glNS74piL2GoAah6STgC5FvAJ
deLz4fBGIUqBWj8eYYFICsleFfUNb0dX9rpafRXpXo2itYFV9UgsXQi3RsYJv/WK9/UFSO+mxfff
5AlWU2K3BX/WnNNJdq8j+BBs5TnbIdxEAdDX/q5ZxVb2j+wXu5wgPIRC6iQEPhZ7PdkzOE/0wlyU
HIDlY38yfBApC19lyLvVNQxQuaX+xyTcGFVtHOo43qpWlrOV20wiLtLlKIJznUwHld0uXGPVMXA0
JjVO747RQPhcA+JJ6Xz4FJN94Fxt5L3yWFyLbbx5MTwlFRm/l5u37kZzZswgcDqmwsV6WWMhsEVp
RU9P/Pi7Az7sCFIF37a+cfSPSpVrxdGkxNalcSG0hHY2RdvQXfuBbc6THTWMRE72dICy+Jwq1vhf
LvqTgytRkfwIUH7ES03yNDgFYsfcWx2kfyrmKrgLine1JnHRezqCEaVZVzHvJqpLXKYUhSk58uIq
HGRbda3mH25VNOYcbPslZByo1oxIseoLVoFJ08gRDRSaCts68R99Rj0iv8STS87tFTUNfm/GuX9C
wUEmX0LalSy9WCslFs2BFJTs9HLacmpPlApEV5gKLVDkobqb2JOLMtNBMU490zVL2BVAKxdHyF62
fDQq72ujfbhICgI7S/CORJELOs3n81a5Yl6s3qv7cco0A/ojotpPI+rF9m6Is1JUC04YpgW848bw
R+7hOv/2gW2BJ8ckHEbY1u2yuFNBjN/qQz2jLhM+bHISIcTzY7sUBtuWF3PfZhor/ziB8nNJz2MS
VuiUkWZVN+x09XZ1vk1FRhgUpgjHSn6+tlLNafPV/5my+UobYnEIgHJQeLpC3muOtCbNtpAWaeND
0S6qlazeybYmI6wiQ4IMZ+8kAwVZ4nDSurBYIZdsi6xCXulQKDn/0NJtaRYju+zWhSY/VAI+ScYd
xC/zRq+68O2EQi8i5ZDw17Efjr/riG62AiocZU7tEeD60MbcWlybK6W52l/Hu4XBskdLdx26jxO8
7+W0B35RkVgSmdRinHakO5cAoby+MfEVaOR1Y16IqNd7grMG0m+85qkQpDDV9VUHc11UJ9FFryPI
eyo8ILnZlFHSk6i+ulXH4uPm4BtODX9hIYFs7XznAoVguES2npudBjS5bmv9fdQ1VCQH4fjCbUoR
/giJt122+LQo0hSx11SogLyn19I3H24LA+yIaCfbhZRC5ZFLAxd979FF6cwDUC+c8ut+dGjN6N9a
g4t7/J7wv3MaJTpm78AwzUEIt8BV7/jAMLD4kJx86P3AsuRoW4gwbBlpbkV6Yf1+TK7DQpKF2qR5
00FyYHFaCz1tuC+J9waso/lUxdwgW9zPIADNHiH+tXlgUD7lO8psCXpyKgR+sQCfSHITdW0x3a4h
bMYjF3T6jsUBqMm6g83fZmBmTCm5sHh6AUtnSZ5NzphzFkOV05Q2LlzWUUwwtgoiBNtKjilHWfK+
VZ8uKRGti3Owxpjo76lSMPsUnd8We6RGz3gudo55e7ToIWDvfoDzoS8ha1i3Qp5cs+66+SPC3fRK
+irCd+yjZFF4ROJzaYWmVPLgUrNC1u1h5QxJsJpeGWs8zT2eEQ5DvIGURfIxFz9/59XOA5F66XC6
M8qQvMeh3M7EVnjSIbXGDKMAk0T37jQkM/w4L4DQ4fSYzxf9kq9X3u9ilmHrCk5dqwNn5AOVrfQn
u4sFRF+nLrD+gH2wMNsmxCb7aTtjffprTRyq/4UJY9MFC3M5F78gPeNH3d7WDlDpL9guJGBDG0QI
CfXIgHebnPbEbdgqSDDomjFVK6w3ksjm1dWUYNQwd6us+lzfWbtJOzxj3bCG1KbGvO6F8CI5xd+9
U5zN2ek5U8M4ALqCJejp4+4h+k3szCkKqQTTh2ijr+EkR91fQb4SqANMQJI3UteVJO9agD5uaXFA
19OxBCxtlczZ5JMSMXF1O7dmpAINTaV/gjAhbIkmjELWrgsZZOhEuoAqg+Va18s9eRqDJl6IHVYE
5eCbSfKHVMQgD91ZW0WiLX/aa8bknk2ejfvwiuwws5yc9SEvNNtkXFeAAl9L/PwIRiia+RwrHq1u
kMLnXCo/RkBtiBEp8gxMPdC0Ymkq0fQCS8uDHH919ZLO2L0DqBSX5sLMkIVANqpiTALP3gP5eXZp
qS5zyC1/LUVartaPHZLMUjAwWXqi1UY7k9CdLc0DyACe0iyFxUItMHDWWEJYDiheuT7J6i5ODBPD
k/eg6mARjuieBgBIY7aYAb16t7FKcxxeNJBZuJ5JE4k/yk77dMYBLoZvwDcJ+Igoa173nfGopiAB
YbrcPNh7PDoV95PVG6vXz9Jc34kGWBYcmc1hZjlZTkz2VOSW4N32C87zPdt4qJbLNcdBcgzgN51+
MBWBRra7W4El5rSMT46eL6VRkx/wCzURxtAYeiLo67n6GZuFHYcdQCJ868guO4vJC3NO4f2rMKBY
IaP3B878qyWUnXA+PjRmmYlPrRREj3sX+NCO5Kjoq2bwatMZ5oGPZ3PN1SA5CYcNxKrayQOIP3Ji
0iNUb0E3pSAx66mQ9fQagc33KX+2qHOliVZQnJEHVF4pD5K9SljiPYnefTKHQ0Fd1jvOzMmILEK3
C+7X3xmpnA/AGw9JRXkFkwCuJoV69c7eFJD8O+BwyWz1dH/7pC1EjD2NfFwJpziQIlRqDBsDq8Nh
s06QvDmOLmcRmFCfKkgZQms5T5eIPEBfxtKRnfzwbZYoRwvhiGw8G3xKbruHWhnTgvkdIKXtdIN5
3EnZkEaXZBo7KQqYSHsQAHlJcGStf9yc8IegrWBP+Q/3xFkXCyeFqBd+hK4henKguJjWESlCIzH0
VSGMuS2JgAkr4plR1KMbzq7wmL3ygtE3cxtk0gkSVlnKccJkMK8PVZb3m1gAjD84W7MNApgnP6V3
J6JXht5wiS2yfxqjlBjQ3V+v5Psa2cpM+4643H+wdqAM8SrWU0r37i9SJzN49LZ0MH/tLwV9Kcm6
giW0M7hsz3wdRUR51vrPskt4Hi1X0OTGCQKgGLCjEi92YECyUtzq/5yfwyuq24byeFEksEv0ONSM
axwa19ZeTIzn/vraUmnYTvxKuUIN6uRN9EAVInxhK9EyKSPwwFUcG1nBlhqcao95cbpoY35L9oa6
SxC2hnCCwtjTBXyCocN7UZnFrbc66xzkIC7yFO493qMc7B2zUvdffevAV2+492cmSbqs9NvtSLgE
MvWiYWOlIix7eQa/9Q1xCylZnokwgI7+ru/1iH0wZzoLeVikBqvD/V+18eZU/xe/siYp4BvYlrvb
gGx8a8NFS+pdAaWPhYde9Jknkq3nClCLJbQKaPsPXCuXDvQyOYYfId3uXFwPcBPLkVQgIOT9f6sN
NC3rru9VEcITQ4OQbb4S+1hre1GwKBYGv32cpk7vHyVEc7UPyogcnBySMzb6TteXD7I9ulcwrRsw
a1L9Q8QzZudiHvBUV1cIcTGqZU5riVbl9DpIsrRQjnvQsAlLjaN1dn9iK60ezoWdyjonQueVWxhs
RKEK9EHoIvSvvJF+PNRzwW7f4sX7zGgk6rEQOsOqi41ZdYbLEWH6RlnCTIQlxZPNIzXIsMCK/Lxg
cqO3yS9q4kBNTXD23vWCwt5okg6v4gv4eGJG8laE2bx65Wi7ImDlpwlxVmVnZdxoqB6KucZ+tCDp
jnmlJWFeCvo+bMRlZdQGHbviLW0Xtxk6UHDxnaasD0uUQFayFMBuDDgh/7fje5tR+DGF+V6L9XiM
I04sprrtQwN8PoAZFcpBzRuf816wINriAuWj6uG9H3Nx8E+Xz0uOCw1cSozUB4mVJgdP8SuKwRvL
6bftwth/beYDp8i8vIMboqibLV8obyrd44TkRbK3WxBNeWZWq172LCilV3eRKpLjhqS0NgbcFz+0
gXjY+DDvAMvToBh4Dd5nLhFB6hfaJ2ZAhZaSIsqdFLmC9HqG9iWVCAETvP6Gxgc67HL3cZ1eyTjU
GTGMkaYb5DMbV5svk3cHV66Tdg/JBHWqqfCbOtnqPP13qxv5ABvk9fczfKTJCpZ7UXwSE/H02uZr
NJaN2t4J5WF+jDGhSfIN/abGzoeIvl7evTT94ytlbQdXV9wzo/zMa5tHIc41bWGb7yWYwFoILRqE
Hr0OtRNVih31+UnZ3Uyjl3hywwP1k4JOBFEDoa1/+XfV17BRgubDO++mCljs8pmVOdlKPiG+Eoxe
AE/CQFIcteMkpgZWwz0Rg4IsQwQwKXnl0KD8pYrwaKXfkMX2U5klpORLuYf2oHVOsK9Sc7knPzZT
hR+sw29Lthpuwan44Zu1G/Ml1hjanQyNyOhjsH+NbmC56E8mhGS1lxvG+cEImg4rayKaaxh+Epiv
UKSwmsZWx8Bg/SYaELYFDJOdisECQSBksr8w4ZkYEzbKWWKqzMIgMFEPiNgkK9tBXD2hXUYRxsat
BWhdZrwXbVoY3RwTMiJEEn+NTYoi6Rx/Gb8W6Kjq9XSLBvSo0Bfwe+QxWoN/WjImj7nvvOw8QCOr
FICIxvOr173rsi8qfpMrierRkXnQK5sMcPTxf4QpOzmkBucCvZuAgfgWptS7sIwUu0U7oP87HqPz
ITRCysTcJVPEIP5B52Rgsw/CxXYgO69NsrY2w7vy65U2n0poBImxFFrPzyENlf8L1eZox6RHVG8r
Ecbh8RLbbTVn75cYVLIGYTaW+lBpUt999XEo1U82v5+lItSgdCJWByCxc7Pmg0/6N4rGyqu6AhbJ
gAip53WmyoycBOQbrpBCrby/eybZ61LUToapV6VQ+hpjZFFpyA22lRphdQNVhNFBckyXXJLmGeh4
ipVYYCGUaxXOoa+LyzkmldyvzbXOs4M4BuG/LIVI+AajOp5K6AyYB0XHUVb5SLvWIlzO+Qa+C6Oi
3ejaZwoc73ch02DPQVEmgdrfaKe+RdxO/8xBlDp7sjmWq6tE9WuQNmKwNkLXbUiesSEgJTah6pLe
/YY2yZhgKXTOAlDhr51OQVatPdiBc1hH39A3RtBkkSr/FY3IBSunociAfg912f7g8fCgYpY65avV
UpdDQeLoqOWUyyLaqWWcgj9g702sr1pDyuD+nlW9Laso1doWhzBAYi0MXrdmBanP7GH2GnpKl1yt
2yjOCP+FhL7fQzEL7Q7FDSUxBTvAznLUGMLVCstwh+H3to4AK7O344aTqCtCxK1uYfpBWqG3PMFl
wyjUByyNpOJlbB2oJqhPLyzfijbqlyjzWtqHBaN06Ti5tVlCxtjZLKGTamH/mfMTNcfWXDlWs15W
6qkbtVJZCMn6o02kBEFuq8Y7UzhMGxr/pAhBjTjZoDwqWWf6JUWf7xS1CxHOqQbgRoKWElZ+7Q+U
pO8Ej7wXqngxaoJ2NHcWwTlJO78V2G3p2x8G6u+QfWllNaLTSw3tBuU3TItoHQwWrgl9j56l1x/P
WrARVFooDvCK64Heo09XJVVGBIKYe3MZM49/GSHVWI1k/IJI1aN8B7d2NTxtYEam2HDAJhDuI1yJ
6gMdSl6aeUinZKX/VsVjciGtyYd850X5imcJnk7NI9WDtsYB+V+7+P+lFjLQR/XZQJmRNKBYPwM+
SAkcuEEuoTmjWCoxPjE4n55rwCNGXww1J6/w5fMnGgRv6dQ5T1JHTlTPnZRGe23JG531Dg2MMmvE
Fk+cxyFm/70Mac7xcIifdUgcXu6cMznzAUqfCkxmT5pHMg7SmZxMqfQ1IV/d1Q95rnoDD06j9LQe
WTUmXE1CbRwcHXy8axnMtA0TGmUMh/j3rPaUn5Eubu/PmQxN7G62ZiP9BjPXwClvT+MDvfiBtyHc
NAU938+MLTAxYnR0w9xPPyzHcJxz60SpxBk81wrtvPLcyJNmubzlo0adzp2PVgcYVujPx71cao9h
04gQvqC98vSooL9rONrT52yJ9Lic+f4TWaEBjiY9qaPBKLcpObx8kZS94IU9Zbxs24lqOb9DzwNb
xRQOTLCLPGeVQvskILF88mYubZTw+Y/nCxn08rfU/cnDD+Q8tMAtvg0wUcqeWbquJp6K1ROLMhp+
QPOP8VXT3vBN7YBlht/1wKyjLVoEFluODVMScipHQmsdZZT43PJbKKu5fUIFJe44JHimSQ+r2frN
TjUFc0CXEy+npFFAkzPd7d7douBwOR5CuWqfv2KIhdQf3MZBR3l0jdirb0bjR1gvh9oIcZxbLFdN
ZntdXdPv3bvsox3zTwLekYAjtxU6Y+Xg7oFa7ZW6R60TVcKBFiBEIhiDkM2AnHgzFhc+fweXygkX
+1HuDMxcIC1eBTJtdSXYgITe+MXAuPBdgQdFbghzVmLUNAGzqEzcLluE8vTnsP9+oiqCgbifcMvp
QYUpDGSsyzPAJ7n3rKCxy9vzFVTHG0IowNEJDEsERCy3kLBcyTX+yueJqzAD9FXs6PPPuwwPxV+Z
piLMSadVZ4Q01XGMlZC56+U/gX55x6HBSxNXTTHy8ueaRbzcJo0fJRFnovFMXhmogZBo1jrG7tQ9
W8NqzllWFR573hwhOprJky5c2wvi/9vnu9Ayk5YXTEsFbXqtTfabgutAIFNhjydxMrXqx/XbG/vH
NGfZYyu4ZwN+x2bjTa/+wXQmTQym2FuzoH4BHGGm4Z23W0or09cHQ0x7GxY/da7vEsxdhicDc0KD
YI/t+l8S8JcD5dgbgF7ZVMB+kLTBN/YGGNDd72cPLO65KEYpxm7yFhBcdoXUd0oNuspGs2RlL5Nf
+mV2gUfYztlXARJwSNRwPxy7HsG6/fXRGNUrHSQwv3eq8CosJM8gaGqpH/II9tvsWcXGf/S1y5jC
UtqDXEoUcZM20euLyULNsOxf/1XKASYFBwzk9E0GVavHYue3oO7bdMFtFTWhWbsVcvIC2NTWhFv3
KDuYO2e4aW/FBQhMIaKHzZEL+oXKPaqr1mD2/vQTxc1VfEnu3C6B9+TdJlaV1bZ4qFIo/Rm49b+m
wcWUGilZPz4UKVPkrvrO32v9Z1TLR/TjHZRY2DJWi70rgMc/6fwKVe6E9n50sIGPCyY2SRKa7UVi
pNlj7JiSt46OhbEPUD5u1tKNytoMhvYlQA1LrSgfDCnjboPkswLN9VK2wzSIhowAVTT/5FLQHXUE
RNU1QrQJrUdEiKGMvY7YbXnCmSndPprcJcYXXUO4On86bV9pwVwaYUcdymuCE+qds/zZwr7VMAQP
MmokDizYxs4thYP5EC6EpbqGGDr74/G3xBzu6OTngo93471AEseHJzbhmBK0Ih+SrYafDQDa6AB3
mcDaJb0W3rJ4HrqOjIAEZWaZIRKG8x7KcrEG8xA/oQyx0jsHgQypZHRt8b3VbFsZRvY1lUkUXsdV
cEZd8TyVzD0xZYWtns1bUFqjo8ugzv0VOCd1FX+iv0fo6cWtO1xQQMl3pg7A5gS5JRrSC3sddYLc
o8muYJjI9ovvelSV4m4hBEDXxfTc+Bhfkk7D3UE9sx2oen71Lsnudu5118vFHB31TRa+n0Dl0bwQ
eF5DMlTaDCviHixklJmkMqKOHEu8vhrazrQ4y3dcPi8hyyZOYroOOsG9k+bBCwCffxnjCtY8ZoY8
uKMwAVRybdMLsknZ4VWlo+k1w6uIL/JoRVgo5HX2y3DnCG4rpiXaSNdutGWocfFo4kKTrVFkToD4
g6QIsXDsccKYwbgSh5EciHHAyW7CFovo8Af+OvKKCMdAA7DQf6GRcpKaGMMtG8gamzIcWCsXMLEh
QdAJfJSF9cO4FaRB9h3uWikFpImqTruu4/dGn3bpyNgGOQyEcB0horesqJSnvISzoMl44r60SSmD
wUVoPg6POfU9VMcL7uva/MvR0NZvbNOCkTsWMCkNv00KamTE+IQKL9WCdV83PSEcCjSGyFAiV2/A
hXuCk4snGqUJ3ElSFNfDTvxz5Fe7SP1GpId3lK2uG+6WWm9B74+6s9BGjtEPBqORZijEBVLcF1Z+
GLB/l1uYULbKmAZ/ntuyfwFFwVgPH28HTW/5zfcwYtS/N7KpwJYMW+vb8b7gWZtyBAkolpPIQw9i
9tMcc213sa4BVMBTdmZA91nGRoJDN7xUR2zC3RkNm0gg5zgDjwE0Od2Cy0y8SFtJ5aj4DJI9BTdI
73/Cq7ORqA1sr4ItSrBoj3TGXeVIHiy4kvKfRSyfZOeKBz076vKdv36xzeUE/9VifCM7M6YvW/Nm
wRtCAUz/cI20BkKWa3GIKFA5upQLTMQQRb/0zv0o/zVhjBUvU8feq7hIac34jP9n9BjAkP2IfnFp
04F/Pw9jkFP0xscJFXSjatoXM7VQk7/Nwbkz/IXhZ8VNmpcvc0xWT9mxTBjeQi6maIB9HWp8CTb1
AEjqzdArvAdIVMpZXkxdvfLtcDZbYxjLSJEJfJ1IedZDR23hyC3M2O4qE4t7Pq3rxHjTIqjcgaEj
vRuzp46cEnrlSqyZRJurDdudeLv5HZf6V/l2Pv6rXhMGORYW2kUsBQk1HEUEtCSx6qJ51AkV8Roy
MVWZ7j9m0mEwXwWuQzAejT6zGF3nCHF8HIavZvXMuV59+B/+GT3CaNeXjZKE0wAabxg9tslECBZ/
Lkvz6I98BwotZMyV37kYv02cvc3hLvVUkVvtbrilScUaJwQW80lWrCXdA24VGn2XAgNmB90aDR4j
anc39vXD8ZZ7U0a9Uw8Qx9vDBg/kTqEeEjnSyunlfPlSkH9sSbVFgY6xAYi0R5d8GSpiSAECpvcC
b1OtjDuwddFksOpGWVWesXyqD4EKNq/aUvIsVh2a3PXpl6ClaU0g7QbXi43cW/vIwFaLlLtNxT9m
lG+xa1jjcapEJTLZgh+5YZGnRWWHRw7jk86DlqnCe9BzP0WtZIS7JF958w8mFceTPSJl0HGHw8Y3
U/3vIhxnrTklciZjm/p/LZ4YIgp0gDBPUYU4RHWh9luIZXIA6sOCxw+KtmLnZ3VKT0nseBn8KG7R
Ue8lwNNWTx9NgGrAf+zj8J7iYD59QS7jT9ElBAVZkqlSNVaYjUaxPLIR56ijYluOGFm51tQZ/BgU
c+VSfPri1df2mXKVtrNvVk75XIUt7eIjCbkpptdaOHDwuuigIKZlmpu0gNj3hb8kJ9nRPrwmoUWd
MX4GZLTW8t9PZLL1tEYnlc3mwqfgHlJmmiTgRBVWy+WP04bSFx66NPB8Q9iHSzejBPT33WuAggQp
TbVRn2+BgkBBc7Blb05do5uordjn9+I78/Lr2Ov4GyVfrXQGjPwy/cu6JCFGV22FTX/MeNh9H2M2
RVDzHIQ/YZUzaakRddjKshp7UY7slHxb9WJ29bmMR6vZQLBZT65xlaGp/i6EUxhW6hnJM3kZ+B49
76rzQnjowEXtxGMT7rLb5u3tqr4XYfVRr0hF0KugnZyOWSHW6XDnZ8K9h/8g1xfvcnL90dj60W6E
ue1kN2HqRySQMALsREOux8oMflNxT8Cx1f4I8Cam4Ek4xsnt7zxJ0Xlsav8juubCphm40/sEfDDD
A/iLKA7BEOV9v5yhq6zX/SGTAuVBEkIBBgZCdij7HYLi0dXFxmteuwgjFh1dAis6KhKqH2pTC/Te
t8ReF3QM+JIKUvdnzG5nsrXwLgh8eulUQpzQrOwXSb6aYE3BC+wuqC2l4mq7MprrSr51oxgHhbKv
DZ8ketJJWLrLGf6t02phTtwe/6Ok8tNW1oeWqN5OWTE45ABU1q4VPubl/1Sy9bSoulz4Ayo1Teq6
GsBe4TxgpHIooLNTQZUYtNYhkmMY98r7MpKObbdLT6QCoHRYjYuKLrsX7yEWffhaoyXz4cZeImyy
NZDNyJFkEWg5kI6BzEmg2654PZaSmn7z2A0R35SKj71rZCCEvcVwjplIBRCT63LvI/mHR2LCsE+i
dNAojVPyjWDlcARXq1mQienQvhXnnpjKTiMMUNDMzwEM24exKAS0RX4xM2+lVlXFqbGReYOWMW65
PlP2JMYm72JbrVQC+GXocCKcaoVJ4HEM0Z/mfdiy/eNOoLHOfsFknDsoRVqnDThvzarcv/DSF8PU
k2oFi4JEgBt7Y/nerY+e21chiqSntUnapG6MWaTFsZr8k7TjBTifcAMyLek+UXkd7+YoUjFyb4OD
ZW5+a7gkk7GYLlWoqz8CpdaSqqt0ePORTpfwpe47IjrFAsfr4mBoxiFi2Fe1Wd7s7yE81GW1emKE
wh4tud5RF2xn5AsbXMWN5z3Wp1V0/tS3c3cXwICMkSZpbKWJT5TrDMMHqfWu779ZZKq9ioZfzL+l
RbJh++z0H08ZnZXv0LAogRsUB3nZkwAHLDOoc9vt29U21Ewj3ui9W8vDynD3O5bYRdXrkNG7OO2Q
sABDsciDdM8+bSuEKB8rGm39i8BtpK25KziSvLedna7kTcmlL+NCX8EXSdDPoBdqje2tMz9rhQbY
qFww/whluEKWmHyG7q3IxEzbveWx7KJrFpIxDSjIXBkwb334vCP/8HLuDl+/ox3+Sq5PubZXaq9i
iOwjz1L/WQvmREDKRZywvL5kN3zmWRhgKSjguAe3LnODLRQHq4+eCvZbh6agOwwkx9RE3UL5WXuQ
EjusOPaWKFdoyTVjpMD6cBzS/0BgfKOJuRk1AlBXqrDLPU8rCPxjjB7ZYIsSEaVNjVfhdjEPvCd2
8pDJYH1vqXSDIcJpl9izyUZrOGgD9SRINweN4AeIqt9lHT2jIThEUFt1epf4N51Y2EnBaqu6v6KU
rl63nlFAt2S0SigUoX+oYIYHkz5vxQHzYhUJZ4AAenZptcOfOdOgz2fTwcuxJ2gr5pNsqq9iLoBd
MkwYQKcyEGK/RPzpGa5XZLyFI++7vYMPK0NhAS7SRhIW9nMdxmejdedwsmUb0GWU/2IYNtxF7ryf
6FLVGsWCVLACGko79f5CBYjFI+/bKA1L9cPRhtiM8JeDVYYBxkDpwTf7YPVzbjRutaOWs8W4OU7a
X0EshsAtSjBoijuwAGvy2wNKaa6zOibM4vbdxmaA03LFEsYJEJg8k2o3hLA9rZg0SF1yFAIL16Za
biGLJ5xQDXFO2wsNvauoxe5A2qPZ4iZTM6nIOKULv+xz62oo5vcrgggvMF8lE7tp53Jq5/AXTnzX
xfFHl6pppvtvmGwMDzN8n2dCE+pBnMNlvc7LcfecCoUMTQHWn34hSCK1u4gxGoswLkRvhnvz3yf2
iuzm6Dmr5fqplrrJr3RgZgk7ONpk8skrO2RADYdx2OJv+D0k6Rk6TcNMh9mB/iCpkq+y7qB6sHDR
hjd/kdNYDoXZtcasPBttbLusRccMvPBcLdsxSq0bdBB2R6Luox0fe3EuRYXCIVY2XtY4t1e6O1gL
Vlkz7VHH9+bLZn4u8tDqrSEqF2TVxiEVdwlP/rWRpgqMDUXNcle5TtC2ImzLWoSDrHUNSYyHYzCk
5YDYwUFZfLhirSdy7KdOeLa+kmKBxjX8TK/LgsfBI4iFMNnmkiEA/fJ9UzQQNC6Iach7Qi3gq5Rn
Wu8xKzOZGKcg8Lg1l1F6aZjwtos64sHuFoEVQIhDj8K7W9QEjb9H67OFpkTU5lvofrxJH/nSneAL
uZtsuyRDm/9p8XxRlrO25ec9Z/NOK5V7MB7wUHj9bltIaQ+V6m24mSwMgR/1xkN6AOLbt3EHvQfV
CsHRfMcY47D/FJGQHf/cjnCqRJhqpfgp85XCFkQRo2RrDmuAv82cMItYWR9voFP7T6qsFacUsJ4g
1kkfD+Y/xh3Z2WCUgVkMjjPY3VGLpxZM92TAKSXaIYDhl8yAALvijpBefJWE1C47ylXI6MZ+l9Yo
uxS0SEhqu1PUOAxaD3jKQ/4ckGINaimho79JhN48233t0GR8rPh9Wp+7LMO/N5db9RQHURcjMTjk
9ZTaamKPMTzsS3YI4+rx/D5h5D+KQ4ELL2U0lK3whfho9+KJdpsyTUtGdC7bnyed53t93JcrqfZ3
D2529PDk/8bkZD2vRDFgQdwhJyeTyDKWiEbVtPGD90Vqf6SQclgdbltiw5FS8n2DJyOXYBw37Atp
LPzCIv5/aBUs5+P40AnEb0j4G8ef+tbl5hVVb1uITypXwv1O5mF/LnvCLqVuW0LUdc8gAzw7lInJ
+iI0sKqnvssvb1t9HmIYpbUkgujyWI/nDTWXNkNvv3GfxoRW0VfZb7QS9RdaNWoqAjsHC+YHZ5Po
SS499EiB9AL4lYsjiDD0411T93zi0POOgUhKzqqWCeuU4dHlIVaxwxC8O2Ys86a0WH4fkX5/r+HM
l+Xn8a1topWoQHzpJUFBK0kXw27oO3adVhU4U05zUG+GxPVSjqKgizb8Fyi1KjAVkIEalCZVCFJe
acpo+W4mNHi7yRAM3UuBOH6E/x72WCYhzebQE3Uw81BrB7+E+R7A0d3DgZB+tVxMHzOy78M2qRgw
FDjHWRd9BJucHiqiG9/RoUvpoV+G4DBd2qqJy0udJTOp/QOXKJsOPoK7p/NzJTeLyy0d5U50wgvN
0nQmHMqU4KYdyqQmY/H7HFMo/FWm/TP/04NQHqbVueePipd4WeZk+Z6QJ0iHiev9FwQpj/ineWq6
xztNRkVnvNVbBvK96s+8+y4aFYvsl5HcVsfEiEM6j9kG+gOKk1z7V9iJnASvj8j+k6oMwhAZAaQq
Ty8GgLTAxPa2V99fgDjZPoHcBtm12V8gVSV0HbyfhGvJQIl2QDrHjYbMvbkDZde9cbAoKt77fQMr
dAE8XEr1JkVpzuG8UQ+rnx1jR+7coyUiN7Q7efwKszJezbPcGAmqbWYDf73OpSgyXs7iA3jPbKCF
LYBkgoZRXXR1+0GLhk5zTWrAuzN+B6mX1n90pmp3Fv4WDgZF1W2l6pOOOz4TEoz0LqXu7We5rQni
YdPP/gsHuMHDLJLXTNe/ht3NTcyTUhBs9lRSJ63xE7X0uevIBkuvT5GtnvT3cKrRc3Nh0SciZkID
nSSZsL59bUChdwDA0j4IlEIJghKrb7l7OR+ksqfo0OI8rvnFYiONL0bzGPSyUMG0L1q4diXq6KKI
JdX96/GRra+KCflaqXCEr6DAdWpK1DfMJAiY8hRDLWYWtOAR3ePud1YhHpCiOdFGoFVWbpcD6u5e
lLixC5DUKQ0OYBY7pqCcYKQ1kmuigeQ1dwnh1RPG5lq//me9EPizcxOJyNmzojVO+7lfwZDUqCl6
FpyCurcbOSH2iZNe5vX5VD409uJeTJmra6I2cYW6OrLdoSQRevggcNDZUybB5a5ne112mbIHv8nE
oKabFOiA4dLLDX+1QWPMjMJNpwrg6HE7sESRWnpzyq+fSTFwoWPDIx1fcM8/X0DnqWysfiCWwm1V
JbQ73xZHPs+eScdyT7hkS5NbdtZQTXa7/vNz4r6sdZ6067MPdr8uEWEnzK6poipwrWlEvDiCBCEn
8OJjKin6KLfPmrajKoEmw69yhSGU/HxOo01rqxXXnLOsD+O0KvISX162UVxQ5oQSEx2hv3TxBffz
fZswcB+D7pXbv9+OVwg2xv4Kg+Q03MAYLe7l9Iom0b2dWnWqHbq+0w3GSqbhxS8mocDNjU7xO8mR
qcj/tzdmBDkMxp1B+TgtiLAf7v9ytHlVrXTZn/ekgDzy0QOhIjH+gU8yzvHvmQxOVWpEm4vHPWC6
nFcWinqqmpB8/Na25qTR9BP1hTLSpQHJJ/NF4nViqrN8qrHsSjhANQ9dk5cqTfsBVccV6sAHmsaW
4nTzZKc8pAQI7klU6EAlo4u4KROxCJaUY+/LtkuFu6r/NdQYVdpU+tvQxGJZu4hRRLYsK8XnMQor
ClIMqJXmYWV/NiFaOPBuumWx3LZ5nRiDc8RrqQAvQ33OOnS6QOCibloY3x00zr/GD7Qx5jJJp215
qVyHRR9cBKkj9OqZmMNaGSXIt9pS9BzjEb36oqMfyQmrlNXIpSf2t5+ghUzAbmR1Hbf9W+Yiel8K
ZrhLdog65wflmhN5EU2AJQta5QxaRmNf0okTfAB3l54wCgC7iiR2HUNhHV4i611EChLqnQElE6XI
/UL+J4wl6VYq2wqvVpurzgFE+2O1c7Sabfm3sQxKOILJ8mztNyu7FmG7/SxWlZzxooo1ZMWdl0wc
BSU7vzAldEFh/CScJ4i5VGnbHqWVxkGFSAxhle9gT10lkS0xnCmBWd6ioFLgbtIF459Q4O4vjfIY
fpq3NxyPP+muIEGSX649+mruX9sWcoY8aTrR1aax5a2rD8UV3nW1R2kk582fBjZ6ZuBUij8WYH6m
bAa7OCLtNNZZG/iPlkDmOn9YMXEQieWfyr1czBMJ+re9JQ2vKcAx1Y+5pcjuv1IWFtg0vu/Jgt27
deH+2aHLwDT1tlFEMWx+K3H/CdqUMstqxc7vLBK0CFOl6Of3wYdfoyTzE8TutRq7mvE18fU2964G
BfMqoPNn5lztcZLcSc/J+hStwXb24q6a9qEZXd6eKDvI/aBI28/gxzKDZxpU7w+uQWFGM2dNEmjH
9UBCt966BfH2IQrJcsFV5wSgTmc+cYr+nVbtkfr9GBD3TaPV1o2tU+dATWSP+Ij3kLjP2lpioKfk
RJtfNf2IztEz5xaluhJbBS6VbPJX7FhTDxBN+6UKKPlnqmu4mm+4JrTVGDrmEiGLlCP3wKkiM26a
RtOLCFOd9u3Xz+qSV1+grw4g21VasYHkK+w8U8lRQPWmRvCHsmh9dphDoVXud8e5wfn2qgCWaLG1
6L4VrufWdWE52uioZIc7CbmrAAT1gegX9Vk4/B3FPREt8nkhWxsznskNKA0sVVVpco5pV4Q3NzJ0
RmICAmc/x+Ip/aiEnjHiJxSXOmnuL02EC25/9ufZBhIYDWXRQhElDEHjfOecnSCsugoHtr0xaL0a
99ZXquawZtHx4zbo6oiJ+Xp9Qu5kavLAsmi3uxEQYXo+slLugG0SgFbIc8bZbKp5GwUtdOVe7kpd
kpKNk3MNudz09ZLSavEb6iP+XDAZ/f3F63rnhtdcfRiSfoQnduE3HWRbjJSPneyskua+F47gLdZY
Sjw9hWIzLRUp8HLI37mBXryzc3SwCsDiMonMGBb5zMlKO86WGfJbqBMNqTlzJ35tS6xzAnjyF3n0
+hPMIacrrzuCK7h8HMf2NBtgIr+i0kzRVcxS+RVfnZt4Om9McACYG+XuPk4KayMcAfO9ZE6OkeB9
FvsbplK6rBjTPLhYtjNICLlv0swWoifg+qibAsPwKJmTs1dskEclVoDDjdHsrTnIB0NTRBQ8g/KO
qr5nGspjMAMGUS5sHMIu2F2hExseM3itP5iVy/jBE9faHOndejNdJ9VQbYqu1HJ5B2jf6+WnYcd+
WlZ/uluekYkX6x9g844mGfU5frBhECLOn8xxUEIJgozu93noM9d3JzHeO2fL3/1VWjvqh2LqWXm3
BPdVMEQKaVHI3muLw2cOKtCX3rTsQsXBBPoCTCARbylKbdAHuXQIDG5kAz3FWCMr5V1L/jaHx0yo
REzQCA5rr1f/kRTHFOfJsHeLkhTaEWiwkvmirQ4fcdqruEaRnqFJJDVLEJZz4ZgLVB274wUYtUcL
6x2WXWQ9nsO2Tf+XTdJY+nvgg7POG575ONXcNALTv9z18P/vXw7UnfWNdjj8qwVooWeNYzKXpZDV
BEMO7iheoRz1MMiwljssbS03NkC5RHLVT9D86IRDzcYQldOhT0JGqDKcs87bIsM+46mPsVjjzYxv
Ven+qHq4Y5jXh/cDCe6mV40hiazuKWFt1epc40xAUZ0SQHyDB04QkDB3sy9wMXClCJ3xJrZfOZ+M
lHtEj7SjZ+MsqV6YtQNpTzDUTCPxST6oo6JcWyg5sGKOCmhuuYsAAAfrWYZRi6T5hFqJKIYTsGJW
wDH95QNWGkR+8GQB2LNxtkuT5IPCTSkNiqlSbz04urRiTRXzNdvIEFekbva8bHzITKxoHcSyyj4A
KTxciVs7K3xS5bTRUruFK4CeBNsCUIxD0UrIvvyRHQCPFLTFthI/9yr+yj1X2/QIhZEwRkjqAesC
EKnEJxOY1yT93mvmp9IeBdJw3B10TMWOXVeDNw1FuBmoLgzTYN2JlMD41YgEcSCSCMc3FQgFWcnK
QZ1mDkV/L40iowVqXmp7KKz13ixhs72dxEDNNyRo7wH87miC5hEqjMGnrpo1lb7Vu72TJj7goRIa
AZjfkDQP2yp8na5l5ho35nD8psUW/lGMK86DmglR+S7AxRJH8z68WoBOnBXyHgufDXDzK9pKE2jn
8dWACPT3AzdzAzPg2C8q3mXmk05yLljoXBWYsha08irH4xRbZ8n0MY5WcoWSLIoAoDrt4IhX/z7l
SdhQCDDKcPGZMq7jIP2Zuxc5ezYAMv9jDaVtWHRLx2+RjaMYoTF4BYPM15KJ3o6uRBLVVTtJuGoM
wJBrtwVQa2tEtL4qBi95tk2hjkasN+M+wVQqTR7b/5NwoHKTY6ub7JFw3BPsqd2zNqo+RQoPcGRt
TesTsprk8oU7kfE46V6lauGRx6FDskvP8Ar3h55kJZhAwGJ/HYfsuKjHijrV9lSRRolS2xPUt4cr
M1QP8H0KNwNR9q9CsLDlaS/1EmbQcDUSRyv5TOFWpGz3c7jrcmgZx+vZIPNOYCTvno5z1fld6Q6P
ZvE+NJWwCG4LqBs08z1AgSH/LKxCnmMUlbvSJ67oSscvTPHTPr/hku4dVo2S7zaY7YS7Wts7sEZQ
a6ZXW/i6/17FUqPKtOAp7K1NJVFPvE2l3PWCJweaHYIre5Gzvo6c87B7ZtMICXSFRbThxyUqR/VZ
Ltccfm9M/Qg8RqoSGicmD2krX1ZBQXsgc9PDX4rP1Axr80rXOUj0ctQ1B/yvpjMrl+UcpOSgTOWU
LBCjNLh+4dYtx2B56B0ehhXJlq3Q/ekzm/6CW6/fgKGsZRgnjS/cD1xxUoxYIJcvO1yzVb8P9Cjc
NqrH/AlhrVi+4ilSbtkwg+JRZQB+rzzzpp7/UP9/XuU8KTekGSc/NhIqZYmisqAiLPkj1M+q330h
FuPC+RhC/dxM9csxwvJscnLBpWCdkMVi8O+sxWDYBgV39wyM3BTjrhnFz0sAy77xGtxhLxBgK7X3
DtNit8mJSENhux3CvApryhf03ypDErxsgvW/5lhfZPBekKIMkeOm3aZlwEAz30EQagdCtqkt16F/
CmsnMlf5bbbLeaZFqK7oUMWqz6tK64vsrnDLGXEFAcJ3adkVWjHuhKa69xkHMetu1hXlI+aiJLij
tJ2oC2PJcMOeUjwGkaHenAXm1InbnI6Nn9wSMjemqKySUSX7dF1YgFDpGMrukq+aNWDWzvIvgTnq
ebgdu+k00PIJVecECjeHcsy+xfYoIlcEfO8VwhDPabjmSzzqBEcDUWzNgWtO2SIyQNVtkkes3+6I
Se0F1JVJichfCHFBsAYnmd1QjxKHfjLbyXXG2suHYB52dcfRnorGOjy07bin2IJFXOwZaRIn2JHY
9kz8MkUdNV2/5TJuHYJNUlBV1TaZeWx4p1Rtud0HIbk3ejqSlpE6ler7u1kzIBzpTTF03HtXBztt
AB3U7LWw2urv5GX2ryFaucn3UtK3+KsMm4xrQaU4K5ZzcYky7QCzoM01w3bbsbxk3MiDfe0+dtfH
kUt/oOIiimAZ4xWWwVZEdwzeRAsQNkvtnA/46Ys35kMjujNPDxHc3FchuVp8KByeuj1Uk+RkZIKO
/d+j1LQG+gQdmCpgXHDxUaQyc7LnQkzzQv+UGrSHjfyBkCZY1WMjHRu0XLC3xZWUrxTXCd9uLr41
VAQSYIKuEtl2BxSxjE5S/EuwK3X779F7w6xgzfoFH/H7wVr47sPs80p0jSB/WASPJYNP8lZy7fZ2
o+RwQdXijcviU0orm8V1F16Fk2G5FKBTOtxdelPIzy3ZmTYZnkQ5a6eu9aMDi3vsMdHOalJcb0LA
StthWq9suc9o4eXu1T/j6OIm9m8U2PvBJ2XfbPnDLzkdnYJ/kfVEZvBq66xXqV+dcH54sxUFVbzK
Nyir11Kk1Qw1HY7OS8MyBudKdJ0Zt/PkWU4euJrRQn9MPAXX5Cd+28tQe45cZIwb+iGC7cDbhdBQ
JpMToixHwm9tUscMMdKwjnklH0lySyAnpyZRfOlAtUofAvlv8dgjORHKVse6+BMiMBxtyoysIaNl
tMllw3wMG8rTX64ZHqHgrIdIENShIhaMsl+G2U637JQOJHRyiHlPcwueSBj6DhrGo9rah9q3Fx/w
1Zn0EvuH8tOBPbCfXzBKUaeJ/andzWdNgoW7ZuXGaNPb9Rm6QONNrNWCUKqhmSCISMV1kPEl6AZ9
E+sY/yNHpMu8Se088t7Io2K8AIBXIEUt1feBoMzBrEn8CO8kl4dS5/Ldxa+PYFEI0c1euevohxjY
WsosGo3b06LfBOiWzEn53dVraJpkUqNHWOUiXAPP9T3WH9y2abNoL3XLlzQLQkq2qJ8wrA43VG1R
R+BNCYM2BCTL7L3qv4xqPLHhEhliWeERB53+Fb09CaN4SCxMmb0v0zEHhFaco95P+WkRlJxn6W6f
IDXW4YdwpUCh+52j8kO+YmaHtjvgTcd56jk0zDppYmgCF+OjEkynEQKUf+7oIZl7wkBgqmfCYiaq
feNFvdD9OM1uztrnzKi68u4YEtx6aWOxMleWF1TxRVNMBnULmTV+Jf3r9QP3AEEhbRyosZQjteTc
XMRyRgrToMLhrVjX9JltX2oJtbqE5MD/uNX5O9Jo65V2g6fSjlKrFZf8AqBbHneA6Brwx29l21Ei
u8wCyeHx8kM4fHWyJLP7dOJlCjeZ3dbs7pr/hjk1FRvV0J9xpoo7Zkq088vSidCeag18pR8spBo1
jimXPJi75AhFYxYBWjDHgbNvJfYimR9Klqlje5Lv2UXRDtsj0fE2wcE/BvaWLTc5uIUqk/ufityv
XMIlWkPedrmoaiCFxKpUN297X83RFlW/RBome3ptc8gJ0VuvCl9v0t2LqP4LQYzm5/ZOEMwHVSO+
iyuNSLqOD+4/5YTqzaOx8qCUZWUYHuouIdycqJE/pIQ5MvyVrXlv5cdNWQ8yJUtS3SwOmS3+LW6P
dq3OHO8fp/Sd18HQNMXikco8Ev2vgvm3500kIZN3dkUsj1rCWL8+2XeN/ZAGw6E/5OjgZgWvS6Wi
TfAPU68XaCy4kCQENqqthbirVVe5nFInjfGfYVNMFjF5djYYnbHjTw9G/lxmnkANXmPeACrX0E8X
lbeHuLkk0rtWjojQx0Ze1rMhfaR36/dG8DsypR6MkTBpSDU1FzNkerE4RFzx4WdBxnrem784yjwK
9mKM36n/7UE1G0GdvN9bV7ZqvD1r/PSWcggWeOBJHtIBb1BsWDa2PXlUlXg7Dxl7qcgS40E3Zz5e
6jj5drpTMwinPTCw8Nt/664dxvG9OlmXcSL+GUdTECQ5dA5KkXpH41i6+0Z1XUdfB+ql1pSEkob+
uOXdI8dlOxYAIbxQycGN8AVEYGQhBHbNeeGlEYmEJrSCPUmBG7R2hRmMlVqieYziqVlNmeKiQoLZ
Q4+3kc87FxW+BkB6jhn8F1tMG0fBcHbvFhceo4Yi4KTx/y9BYiPmNyeNp5yi5VX1AhKwpXccHLDL
7976c2WIQ2Vq6jgdfKc3UgpCtYhbrEPORp0ryHQ8cOrHVX8he2IYIQCTQv1vYDkUMs2qb69JdH9x
zI1YuYlRaHfLCjt1DT9isuou5rBHx+47xcjVGlmsOsXBQ5vjCT0G5SxPj1oRhhfQLwnYHzFXPKLC
qKYOlpkodOqL7TIP6p6e/r4wiPJuUVp6VwnFyoGNM9LTQ4eOfJh//Q9hGPZd4HvQAuEChG/J4SiI
xhDyhkfT4C9W1ZrOzoxvCGX2IhGxcg3YVeavTu5DFUuiQj9NhuQZb0S5oZaDukPKRmtpWorV8CAJ
FJxe7azJyUGm6aJJ1RL2aNsvDHZulIIsH77DrghkQERVB9pTIVnuJ5eNTRMcAu9xDlm2pzmBhtrQ
gE86XH1+xNoL076jK+ZOejC8gYasbl6oYwv75Ejm3E2EQqhmlg0AOZiLvZ2sqpfjlvfevr+v1Dt8
NE/XVnSzdhXsW7nCQmJ11ExGvj+bxyPtbUxf2FjkXiu1ih7PNeofIdoe9o7NYLvx+ZzqqYRXXPmm
e2OPySHpfrum4K9PuRLZhn8h9o+89+QLci2x4pOxeauc5W5VqjWYy01sau2DYwyqaBsYlKxsZpqm
iY88V+QNXSq/oPxEWgLh2V31UZKCo3yLmwk6rtejIpQVZ/W5WCo9hneESiok771rxvZiaPHXinv1
fGYumg7trIIyiGjlb6NQto4A9prm5LCTxCw8eC+ZKS0QtIXoS3uUob6KPKVTnMGJd+iU/jz2ldoH
kQD9cMbHhRj+cbxxWntOoAFcXE0jZJJVGTIUgyyj7hVcuy13QjupOMXwWRDZBpn61q+D/A6g3m2N
v0Bo3AO2vWNP1cIW/r8TI1t/ds6xAOtv445Ktqmbk7qcmpEST+Swllbbp+czOVAOc71G40flcSNx
zE9wy+yhCoSzQrICLDANMOKwEgCl2adIK3OjjSs5OpYuiMadgxkCrFVJQZ6iXfrUI9KuVaip2ZSS
SilaKl94rnC2rYUPiYcPdoZFGryfLJMGFvBglxAWdS6q5NZzTKcLd3J5tqMIKDIUNk341BNvDaKP
2e7gCxGEWNc68K+PPixfH9VvtCNbxAG+lnZCTo6VQE0MhrLWgztk6XSjkgvT8tJI4PIfwwgB7pQw
vPngu7jBoCMwS6dTXhYlDm1nKEz4GryCtpMm3FiXAVAR9C4KTuHGg6Fr5QWcz+LIm340EDqSOVMd
ICsONo+AGlnwAQKyg9en+dgZPmCV73EqfHxE4/G4yVzQluhcqV+i9C6tlolh5/aslI+Eej8uQEkN
7ZiQcPYgJLiD2+hpmcgoaLeyMjEid1/QnMGurwSSfElLLCgAfhHu6J0SnjuERklSZ6NC3x00K/lb
+lytzsaabPI+7Blhj7mhYf3UqorGwbyxuQXxJpfNtW8Uvz3i29WRuWZIclJr6iY6bSmlIQkY+ySp
4OP6S707EdNW/cOTH2LSO2hILzcT1i1F4cGM6ziaEtSLJwq2h8Etit5zTMIhbPp7LVb/TJh6ntMV
7r4ETO2rFNz66GSjfr6jfWr2ytyjTaiSl/m+b7vwXsmMnnnPJAt8XEM3BERizM8BhFHPj+6Y8An+
Eu7xv9AbEbQEl7GrA5NYXvvmafQakdZXVW+bitfKXMnC9qt6JPPcHi0wdWVnpLJRmsP5E+2TKobs
Q1rTrEnd/VuKuu7rJaCw4TcUakZ/Ga4a3PpQQ5ysa/yeDiYRol7XUX6Jxhmsx68YD65fdQmff6zm
Xu+0GWe1uy0i+a8pUHOU4mVWF3oHbfOt0/8pCdaQNqZtDwnGe8nJU0TQEWgHTS9TdNWkqpmuB0r8
cKLsoCqToud9/g9aS4ls+uMdOWFf112FxecWzQDHyKjXByva3dB2VaZPFVw1B2uasJWmYvDNI0Tf
i8qV8/NTQ+AuBfEnb3D6z+3cvaNQtURrl6PPKA54y3eHijXkMHpwX8k58LnW4kS/SIzMUk6LSsWW
VTUNoNbFAUHf0Glm8d9LJKG5dxerxoqVZp0VSvjkBEAorFy5cQOjdNSlCNzqQ/t6f87e6sGgQr5h
JPby6m8MVGFDWnVBx5Ha85bLuvwxDHA0RsfnARSFR9A7CazMMrYjcf6p5QnDTE+21IGJgjvYVLQe
Ko5flMB9XOSDHgO9Vh3VCniUwUxc47JaVAfcpbEuEHYtosOnFb6WcJ7yEYieQCZphJ29xvLI/Bj7
BVNhrcfmuR8ugaNuwOgR4OYka14qDosvIe9NW+gCOFlDQGpruVI17i+9tXTI17tO5vJAUgKlNN7B
pU2C8l3GS71btnEFpDJ4wYdT3Y7a8t/owGBlkA0gLn+a1wT4qdslL8hFEQ412plFkIbyxlf7yaW6
do7gQs1i+UppGuYd6FdOy4z5r9A39w/4cAs+CqWNXqxvSFcedBd0OPHDw7Gw3mIz1FAz9q0hkEcn
L9PDGEc29AZK2QP1GxUvyHro9tLFsYMM96f7Qvd5ottMr+ZX5a4z8ABUeWVAAKubbqHRkCHip6EB
um/VuMYQoKgUW1GFqmgtNXHnA5E/A3SiY8wgSkL+wFcR+g9EPx3nR/lrIWxAQbM+b+A2LeVwpcfD
llhgu18L7ER48qK0SOWmKJzJEh4sQFS7N50Be2fUhFudmbuj/yYW0fl6XTp3+b7kQSC/sJ82Wqa6
myT0fTNALbzkHqlb1UPCc0tmOhYZdKdrJo2lW0OqpQIxvVrutcl91KR5quRaXJZA2s9U9x5QILwK
uWS0b750EENzlSMZFGg7b0h9K4t0Tr6LN0XMldUdg4Pfyj5pXbqQrN2qq5ef2vYw+MKOOEISs4DV
dC5r3LEjb83cyw2QQScPqIRSCmhYuxsMclWnDUAS1fZFdmPbgHIxJEQs22rRfw0TqcmqMyy0dIEM
N3pLCpqYIB3B+14Jw6sOXla9E4gMYKm+qIOGMG9Rwh7iAn0IDT4/rchPZhwprsVRmcCZ1//P0OWh
1OD5RJYoH4m+1lbURt4nZQdp+epwuCMke7/VcLisaReq4VMVdGchpb7YxcyMcqmI4iTUgu/ezuo1
EbMqJAN9Hvzyf6yXQS7e2ay6ikywweGOAFskx/o0Nan+rh5rWXf03CObw2jRpysL0Si1mmicGCgH
DU+7AAlV3dEu6tR+JUzK4+nn5a+Opd6hQJWWnr61vDrI1mrTj/NZ97tG08GyLjB9olv0FnV34pB+
T0GikwwjbMeLVcytus6oPFXV6Ifur6BrhPiDjxJUVhgKpBLmMJpXuDNcL3hHsTWhJeae8HUQaPcL
Wbr+GdXseKBsZ0vXJam/Y59EKJu4tZrpRR9PPniKMM7341zUqy+ey+D1qBVrLqUeXXB3n4QrSAex
lGnnjDomo1EAW+eeD6nkjrrkmaIpJNDW59rq+UqPp+qnMk2a4wko20kMWhCv1WA7QtpRnaFD+7dl
EJL7CTyhRxDrxoImfAxjIHrvliB3HYF1FnEBreR0lhruaDwWpAlc6etelDg9FLl8Xg32MyQ68Xdm
XJzbutxWEOdE0jeSBOhH0K5dRums3Z+8J7+oh+CuV8HPeDci9eiTxTZWYALp+G8v3bLlCEOta4qI
WRnapf7ja7ekIy2VEpIyz1Wzzm6rwdJ2foXhNIqoajbDW1xsLjv/7iPIpYw/AZzDoNdtJhxpPGn0
IAzIwAYN48f7jBEWX0s7H2/P7CoDPcK/qUzlXmTNbv7czUofE4BjWsSXm/Mh8Y3XhrzGbQEL1Mw2
FPAu3E3BSzAR8ajJB1DiJE3oFReYgDSvm20mmIlU6aXcsmxPLNcOjXc5czNXlsC5qToDZzCcIRBs
t/rMcdT/qUlUUQ+EneZ9Pf0Qunl0ECDeFqJ3TOhBHVeOk+rQfRHdzx5en/fFcatct6K9Ufr0my9W
2VjH/HoLdkntqfYqNwZ6TRJ/oWxpDgl/0m4fTHuUT4xHAYg3i/lXjt9MOmRgMuD+DMzei0FvjBlI
wXCRrW7rWyPXKYTAlSzWGbZdn1F3+CUJfkR8SgV/Er8Im24pCLasPSlaS7oi93805y8ntuJXPJJl
0tCCzWQ/pPqOELySBtvllRrZGzNCKxSNqO4hwxQ7w5pOkCwwe78BsVqkp9GNxoXYUtZnLmzq+K2q
R8p7zl/4vRsDlxBVRzcMLaaDGu9C9l4hhsNGhmA+eVr0JV44EjadpfSofryfj7Rkiw6mjxDnAsdL
z6qP7EP5ufe8QaqX5UVrnJHcZN8VH+H75eTInmH+Zf0BYU9e+4KtNFg4oR1WhX9GfBa3PTVgdseU
2aLuwCCcJ9KJEAGd2JagmGOMqLf61ncFdWmfQifj8QH5W3pDoARSQ1FAaPD9uWGiwthptAEtI3iK
s7gGU47/KYJZmBWJQB9e7oPG/wWWTqMoVjoaMtURXfUTivn7bBE6VKv5CkmcJMUKOCaBvxiR0Gx8
YNJj+iIQz/eJiF+1VKOSI+h60doNQc9xvzS93PZDLR22KqbMk7m1dS26LyF9O5rdUiLNoArX2yM7
yhWjGWzsxkfwNPG7wHqL9CuqLaeG5toCkOPZRyr/iVFNUgr+TmP+b6UNqIoPwjQTA32+CqK8/FX9
qgh4lHtFYZ3HAV1a2yHKCn9x9fC3yJxIQonlz1c8A/FSZ0hdflWtnaIpXYsakINOpxTkkoDKy17T
ixYJPn6yrluDQdCcKN/UQi/XSTpu1IWVz0XmXeRSPyW/1Z81o7E5HLJMdOUDaH821eStE4+EPiUs
yxxlbym+osNOcbqT+eOokPEFj8EanOVF66OhBgPapsyIjRMKan5l6psTm8kF7Si/+JFvtbfKb3yg
c4cfSkqbAIm5pnPF5yUJvwHv8jJqcBU4wWirkLKfs1rvbQi59rllkK1tUgeYhyG4CjhaCQMHHnW9
9PhoST+jS+RvwErZN1CdPoTZPMWzkJXjs7kaj9xhXybGGfS9RRzMUmQn5BFuFmZD0yfzYKEa8wAu
pRstuXFE9UAGrkOeoXNEmSrLoe2FG3zzg+TxKVnBkFYYnPsEhuO88EvimjWGbz10eEUlznTgpmWH
Hc8atdoOcwSo1TcZ4Y3rVxeIU3LuTiZF4W6+42LSmsWVEKe6IDYP0QEYjVa6KBG9gsIVd0iXmWih
W+PR5aWXKut8PFcBne4gikp+djnSY3acXYhrayH2Wy0q9TQWYPZq1c+lhNG6Bj0koudIBKhtzRAt
O5elCMkc0Y3VWHSbmIxPN1yI0FG51mhA/L5XIu5p2Pk2cRtOD3JyVEMCzcfGDIlZxdNGsWzDFzOz
3E5ulr7JKHvd+s5Lsduz+diCp10/l70dGXhrVpbOmbT5EkHbIJt9aBBUjgcZTRaV0Lq4h19fRJwk
QhTW1hu6i+fF2YfSsZntZKvTa8kDwoVEbeXl9ImjReSvZlpq+uuz/VPGWuVCU8I9YzWovg/hCe6t
oWkVwjeE/mosVplKS7jeLnbq+ywSbdjgB+5O/OSpi0MKtyPYO2+S59mLh23+bv+vt6BLnPUEg7ac
m3DIs+EPt7oHTksx+MdxX3pGwMKBtV25KDtZR1ZmngCrSiF3PUUyaWM+LU0HEq7JiBvhU2KVDvs2
0YOseQgFYHZ/PGYErssifFg6eM7d6p95BmNlanE9TdF/nMI9TgaB6FwCkrSqSeF8Edeoe9pNe5Ka
j8+pQq4YcsOjH1Xbcvlw5VjNEICAg5Zu6U2DPq9bFUhJKhPmNZfIcW5Jnt/BYFIFSRPhNNub6QHy
IEdBJ9Gg9frtVkkO0+eFLcR5i2Ws/0RERKSU5KdXvdwRYmQicOlRhMmYr+Z6C3h9v90ZbSj92DcR
JJj07xFOx8dGUpnZmWDMKSE5oR7cbzW/PnLuvWNrfpB/LRqYPWaTbpb3rYKP3D2ylJy8I/tpNnCJ
cYlMnDxrhOT/45YarRZW1wjq9B2SxlQn1jlRyx0PjcsqOfJvgcjFzB6UsmSTmrXUVxr734V8Aev1
O5fvymusruFFCnaiXkuIk1/MYdqkH2DYPXnUGy32QL/vlQHYpgDTbI11xynsASvbj7N64yi+32ZD
/Iu8KsUGmSCSi0uar/Iwhnz6spns8R6rMfh7O8hCuv6px8tj+Rqnobq1cDkdJKOJZV0NpTt0ppAf
W8Y5hm1vgoIig9eWUnixkg/YloZQ06sVDjv+YWg2c26h1wQkWr8RXB2uglEh6/EcF5KnuzeMWd7E
KLxKgvT4631uirKBLG00iLDIRVKNjn2vkzH72sGcH+XDWz8FgLQxFHezo6x7bA9ozeKBQUxy7j0Z
cPdiVPI7XcDBG2OYA1URlfz1U4RuFMh3ggkbe2DpL4AIEaBYoGF2Ul5Y7q0E0F4nxZafc6scERSo
bwSqvqja6wdSOTgfLUxTvVL0ZCgKHmv5Uo4iQvnZlvfRdK8WEIH8PqmwL7y9lQNDdhFmh/vJGrCQ
n0miVd24biCJyRguA5N7iiIzW1gfkuzVDXoZoivpvcNBzkSDFX+MX+f/avGoy6tab8lGx2sXkjNp
ErNYqZTry6zoDBCg5cgECaFDqZHRjc26dRIJejSyhtYDAP2nUbrzTrTTKnqcChPz05gyWjiyYRLf
aT3SXscCzxU1YfthfYjEmhcfQF2JyH2qqOd0kQ62SjYAQlRnu+7OWq2EhXiJXW2Y2n4yDxW27EQ6
YGMFrAEV/IQvSCygk8GOFshTgPK1OmhJbqzjI4XNF5YeA9iv7MKjNUylz0NhVLYN+kd70tgbDNbx
NSl8w7qC+uxHBSA7dDPm4V5WNvkWkGGIBXbFRS6NG5PTeldfZKiWBvrQ82qKJ8sP0qXkiqAsStqK
cQ9GEi8+MynaEgE2kYe03mmxFf+MBPUELtPoSkqyQ6KOjTKW4jsZ8RhUZY6oxjeRtyCzUxh55TNX
I0RTwbsFytyo7yq1CXqweKxNWpkC96n0svGa7MZuaQUCKrUNa6hGvnMu6G/c9l7TfBYfO2DmD61r
Kam9CEdoPKK2KdLrrmVFoFWJse5wgw+eBE7X8rH6gT5i8GjwDgCQMcQp8+OVq8zCuHFc8ypqnV0K
MpurBvfwRLJe5Bitt+sMipVJomdgBN2gOPg3Nn8tlkMZ0zQWdBokd4MVRnS9PT76dZI2rshnD1+z
fwVSrQeshVu9cRSlCCursZPzX4DwuNQJKgQDjGOx7IxT5YCVeFPzspSw1K/KOrku8Rj7DnZaVV+9
cMrwYvMGkbG80DzFPIwX1b2gq5iW2EUTbVIbEN2W52BBi/v+vB9D3mGPYwhJgeoBoKutk6ALaXtG
O/HIqBIcKZfsydDI1R4BIl6UnVniQGXBiV3AfF+CSYCfKeWEYvUImyXwyO2mIfJDnkHbXNebIX7q
kw67bE+OlS244fy79625CgSN/UEMC18zEvduco0bdZdbYpnJ8fpXsAwXC3OWHpD6iP6afaJTdEVn
9yjUyzugDQ1z4YI9DGlOOe0WWncMe2RdbKJOFTo0ioYl0FhuCuhMBtoP5sd28M/KOIyMiIn+B/yr
3XHGs8Z8vmI9TOyiwDOktWvi3e2XXMn19fpr4UjJLXkgRxKuSovYjr2WEoaBBWVoGgiYZVW508u9
FRGa6GLqi/tJQUMEDkd9DiNLIiQLxWzntWTOmGYZXib24VU29Pxl1cv+FSJrWjt/pzavHwZSqrBR
PgiFxaXXrSZvopMcwG3dGAQnoKdqLNLgASQ0pfqza+B1hACx/y1h+BzqsaBxfvHaGSANXGrERtgp
1/ImYcesd03CpcxVART7fA3+ninDed21hIgxAq24fJJmM+D3X74P/cTb+Fph46Vn8ONAAuuqUITA
fUGKQb4Wg9CbT03YMO8MoZQOkWoIAoCgTlJ8q/HVFOnMk+1Ro6SjyPs94mSUyUcThoQhOpawMdVs
bRlTG22HVptNflPT8H+wfzep1M1K8G6dj2bxoUn3jqXpAiVAWNQ6ercNB/16pBwxpgOSZFQZnB5P
+SSoKKMxDkCj/xYi0rrUfehKMaK5Ejwn9kqFKIO1Kza9dc+w9G02aHDTjuIJEZYpBe13J4IzaPjL
FyS1fBCCxGwFA8SIHj/jjWAdNIerkKx7fmC0JPgOffAjSohfqQDz4Ie4Sa/Ng2QT7Slvee7IwNS4
eqFtpHGcXDI8mhWJSVg0qWXqlR0gFhFI8ONmUcqLf12sXCnTJ+54WInUXuCDxfNmIPjdXf4n8MLo
+K+QxXDTmjLUS0ybxPPvf4ZTqPLTf5VcM9MqFOC6PVtzRLOIk3EPvpQW3rTcx8E7d1Zmf72TtmX9
CNkKoEY/gYWqYUJucuxwFFAyVh+7M2JVdYzCp7xvA04Omyi/6Hc5e75hNUb4ofW85tqmtfzvVB+9
65BqFe1BDZjTU8WBAYQhaDmAJ0djXUoM4pWM8Ef8zjS3d3URvtkjUTLPs/ea32whiTBWb3twlxnz
N8zBrc16w4n34kZgIFjuJn9ON34NHt06zFjWKk2Jsiel1UwNXaBSLkKTL84+W2S6Jv7cUBRl/vRM
bv/EmwJUOSzDlYJdR7vZdZZCeZtr0QGXLGA0zrMCdu75Z0fwNeMrrvx8Z9SbmcxpnNSpiIem5Btm
mqM1eppX2jbprdRwYGz9GcX4kZUCKIZ5S9fMwcCja5EIjyeJ4+a+6fq6v+M+zf7FRLOJNF9pZHHW
h0z3LnDm6wFNKBCGOdqh/GqGVAx1opPC/rq11A55x1+dpcxmCzNdpMCksU2gTdI1oRIkhPhbhoIl
PemaOtVKNHrOs9Edo5X+qlKOXK7dowdhlfFhfRL1TCI7bckcC0MulLx+YNIXpM57GtSUYRkI7Sou
Kq+50ik/NXkzda3y0iTcQm49CfTzxfYVOKwBuuvaQGY0GEyQCjtiPVAcCptm2WwBucCW3iojXRZ/
IVda+dvu/bqpsogwtuVF8aTpx5YqdNAMPTd8N2FXD4v4x3UupwoicOrcXn61ErLS/TFssljVNYnw
8qIn6/D9pJqhf7PlaUospMje3kCQq0QZIDiXSDSiYyF99lQ0CrHZDaG2Qj8T9fJOGJgE6y9f9yA/
aClgX7mQkHhbdv7d49Azv3c8mOJ7RFj3wyTaCLtXome93rmZc9tDVwYcTNDW92GgGH6A+GcFSxTI
NyFRd8Yoa3CgMvd+/i7xLT2ZkUgsWP/hY5uWe3uVzwYanzAASVLjOThyr69XWFWTImg7C50EjE5Q
hx8htcw/zCozWnebDCUW3MYuSdmsOWcXg3SGsH+fgsBdIUsfD0I6uunx4sdKVqXaTc6ZC7z9gUq6
kuM7tDvl2VqLJxWvUF78upDsaHz7ZBqnKsnrzVpzvH0hi0lmuIvFSGRFrG8ZUZgLwekX6Ee0LyWK
GeuqDmLtjSQvLbYbYDswS1xXW4rAbWjpKgcIJvJAPRvbqa0nNfOARZ0Ux25jTYRpmYQN51eAeJRH
s7UU++rqtC+j4MDYbyRCL2bnhYQDEzG15kNta6WOIGqh8zAO/ais1IeR1sIrVYAn48nLSScEc4jv
X2NWkq9k2EhaAtnFqzKRe1JLtjD9qYYxgwSnTwArx8Z26PnC6grmLx1yOL95TMrI6xfAcwkSQIGu
aBXCWTtuC6LanbVouJT2H7+vDyTYfU+MdSTPraC0/UqSLJPXvE2rgaVPoTDTO4JiGUvnqkcqSHyj
DDb4+pssfhes9+zsOfTny/xw7WnNGXVe5FujaIhcCcDBZpOAd07+1njoxbQTyFWFTMwwqmCq0Hys
TBVdSrrCPdfkAe2aD/unfOyuLWdhgDHfIyBSin+HkTrW/d319jeeI7PbzbuMgrp4pc2q4yaG9Q/+
Hv0EG8HVc3NeqFM/7V2v+2Ch6cZkUGOfmGISI0Q8hotuBh9eDPm8oZW6HfhIgHEy0IOZZ/VKRVIG
9XCFiEs41l+0PqwwVIWXH2Q/fdz2M4QG2AKwMx6eDERarxUb9wJgxM9+MfA/sO6AV2k6GiZw+chz
CJPSti2iBsXpofHrf+OFwqHylUgU6uCnbcIMqkbx0vALuRtaZJmqLF50JtdXeRX+oTZzftKkd1/D
KRHbgSKV39StaOEFGsCDycIYzxZ2fNAoOwdpSa6BHtH4FcWQbJkBR+/i48DBpZtk7ETfccIwcoBN
pFajnF/PYp3JX9YFnQNDtw1rNCieMO23UjYgyDmpfNdM8fFcuH18Et0Lhn1YGHRkeALV6Y+VwhWT
AMCyJ1eVsAHvPS3Ay/LDTZMc9u6Yo4gB7QcpaOGE2owktavf4GN7KmaxKjqaaW+A5MCYEwttOXB1
TeGpaEw9Uz3TaEgtd1qBZmi878c3aluWnmivwUYQxg5AFgu2fq/psFh3Uby10cNaY49JylDQjli6
Xdaudd3j/MafiDAh5HlRPM+D8BYn3U1FqY8fqxqteS6D2pHozntHWaBpygHYvdArTxslUc/1umRr
ZBiL8YByjC3ptIgXniPoK1blgJ5GydgNN41IiTt6HDtduIBk60XC+UDoA/wmzR+dbfLPeZ4sDr0v
OvzIyGhI+erpjJ+fDmjpM1BiQvBRWDbV90sK+EB1a1qF+FU+kz/yj+/0hvJUWCRYVmc7VuOIfOF0
2HLxt0Sq/QUAvBtB3QsLKmmkxYAu5UyqcchLIoZmk7Znt9mVDlPk4pY9MgD4lNhiPkBhljYjFqw2
CfzAgCAt0E3HWzPNjmfLj6lOb32IcXKH9ovwftd0KeeEfyXS3EnL8h3Spy9SDjOHwirfpOl8RiRE
7xoLgG6Ktw5cpnXyKB4YMTnkzK/u28xb1d7tDFS87K4HFT5P2v82RQDVVJxKHbKeDvpJVN8M/3Z1
Leuuh4ZMzmugHTZb/8xWO41FX+YbQ+a0M5JDQuPDUbJpOBSKd9PMKomRloCTnqCYvjZMK3bSI8BT
WwDgNHIri73F8OAlINiI/Qj/Q2R/FlJDZl1QnEjRQJgzp2DH55KduRXPOe+DLUr8yDk1KvdMEBbk
ON8ebYkOpd/gXq/h09radHWkUHs4LQoUWi14uuhJoKk9o2+KGW9yu/JE9QdDnMnmkhTBUik10w4V
ZUoRLtYvZOTEPZ7LnkbI/MEz3/R8vCpc0LSCifsnvHM7oeymLJV5agIJCQjn9WDli+4sfuDDIqEg
8KqrNF3qHJt1aWk+sdHgPgBzTdkaY8s2UcNFd2nwsL5RjHlS0nM+a49oS7vG0WyyetNw4LAk9n4X
FLTfdtASTTNTUUAOTDTM6J+Q6snEcFOeZwSByzDKUpxksHEYakP7f2LrVwbUIiqiuQHNtyW6wSTx
PlGGj+LKcvzDBzgEJiEY8irRvJjaQW6odtOI3vqB8F3wy/+jS7lRAlmWG4XwSLx8plbu2FugFmFq
aBRNkeRJd0pW4GrKTB+nUO4PkdSMevD80YLldg2GUXu1dPi3SgJeXZ+GncJ6cWVA0UN0Ifdc1stp
S4zsfxrgc1iz3+J2tX40mZNBKkx6SxMX9Qdnf6TCqboxQyP/J2rNla5PZTM3VfnBphfA5qH4ld6u
monhEtwm88Uls+K1RkFoTOIy/xVVMyL5Zn4VGn0io8nT6I8/HBnhGjsUPqOJMQ4kgNxLNnyqC3iC
mZcxJYF91v9XHpuHCc0MY4khPKmgTvZs7sEJMs1UVcB18mxsU58nYJoDK2gl1dvbCKreXjSOPMEK
BsSEvUNIB8buBPKcqCufh7HDo5e/4nudAk1QTf68C8hM92Kyt+f5EJY1YpP6Ah1NOigYWgNjBsXX
g1PO9yogF0awZoYBkqBY7mv3kOJ1RLQ+FmN4PgmkZMgLb8uricCy+J5mCW2TtabA8oiMGoriW648
ygDleFy82Y/1RADio0++Jwungx2Rg66C8D9AS1VLK9ZOi9yAgv+VRfZ2CXPN1tZGqqaGlnemx56x
JRQ3TOOLqCgEQJdExUQSZWBYdeHRonTD5cm9PFMU4q4V1Dacs4Uz/6zw9NLe2lnuCRTdPRXPGR6G
j0z6pKgcv4WQpPxUbQeSE2c9Y76zTTMOQKfK4Bj3B1hLX6PQfiuYzitor1HvsPc4tW9BsHzAXVf6
ox32fwCrLMBrKieV2iRm88C4tBkSsEjKC9Lij8PJFAaxCI4wIdKjiqjqp7LKzeJEUOHubURPuXJO
yRR68NlJ8me9wShmnDHIYlGbltw4lLIuN8+hLq/6pgZeZoV3s4YUEses2HXBfbBmnPWcqURiJCg6
ZDsf5fjHm0aFN5vExM67bY7fYffrQYmwgNAy+CtRf3wTfLL4HNX3QBdhCxTXc5xhfOlwQDcQ6btK
j0wIrDCEST+BwgpjroAOlL8kk8tnCgIylN+8kBq4znlZx+bajSvKU8OUh2LliU24/NrNjgSjUy6C
iNlADyvyGEds71GV8KLFKGufTmzQjbl0yCwXwC2xU357iPF/gyuCj5SOIIB22JX/XCjbCDXDT1eY
gtlxZniw+B8CTd1zFFRCLxQckW9QhBzRC2EyugXaFiWE0AGra5hQBpiVMVJVxOOoDVjVefwqv85a
DGP1s9ZbUIfD9vVOfy7FpCO33/hE2vHTsjbCG0hzKxIJBMflpCuSnLRBwQ4xHnJ+nCUyp9UXhZ2c
+sT8pHOCSYnaYNOZi6Kfb6NjuRcDSPhkae5B8ttIyL2ssQhRHx+W4NdgLLmvsPJnQdOGrV+7WGnl
o0XrsaNqoWn69qoxGLIk/VObHZRZsB8HafIYA1nCA9qjvfZfoPv3xqCNwhRSEiuxF9sLK/4qfeeL
CE/lUtntpS4wV7Fqk3qzgo9l4tqMTLXUDYHAYm0PUhjv6nEDPVd0Ow8eSJM7OBNrYsf72AunyvKT
TfXV5Wk+4DYZNOLgN8byCrVOyZT2/4zQlJFLH3YeD+jJVT0kPyn9URikd9jVcB1EUVq9XmP3zz9v
414z9/KQ/9mx7Pp/0BzP1fFo4BvfmECH5l5ub1Iu9I0QPTlVhobnglPto1XBLmvC91vA4D58x/6T
w5/JC+xOHW3FCNgEx0/35IFBZPjNsprqzZbZeOUNVqq7ds7BQ1YDveojGLKrksdzE0TdEU76i5sW
4JbXomjC7j+/+yCDjyr72C2HrTlmMnW0JI/edzF36R5W+nT7GvmbSMHg7POQO3a2RLvpETRy4jKr
LQBKD++RBAJlc85GTjhaTV5BRiyjbHRGH6zAmrbypD2Ci+m9TZyUmPaM/6BTKXBaBoeQlgaSoEqJ
hAdKyxBckSOWiekgrdRs/5Fb0eZ8HnyXxLuVGdBnRGlV3QY3BSDwsmpmVaNQUt/vyaffSBbU5g0y
J7EMo8xXG34D7bxd2pucCzIIPTCVBa6K0kQhThAzycTRBmiJr1rXWRiTdnMFZz/k/edg9lj7cRa+
Y4iUm2LKQvYERUnURovgU5IFq4lru25lx9LDUNmPPsYtoIIRYQ3mMtwvt4+vNO1ID8oxavWyjZuV
WN46tfpmYsbSCNeDw2yQHpc+qUqW/ryfWhU+EygIBCXihFv8rsO2ZTFhYagFDCTTpk2sDID/vjGc
eh5J5ZP2SyIAoHfgPc6R1oSDab4Pa9fAsXOSpCixuVSQ+EUj43kQnOZLsF8GZPx9NNtnstC3MG7p
zIE6lBN4QARztXljxRyeauATNIcsC/iQ3VQCBqbTXVFU7b8qngq04DKJs6RIsgFVyG/VrngNc/I+
tT42XA0v/YTwDqbRulb9I/PYDrdKsRc3WFsFDXmAiK+yAvB/Hq1i2A94prArWHq/EJ4i7T4Kbzan
agxWlZX/ZTnEGfscY3sAXe+VDn72DJOb5h1PDniyI0Rv6TXY+TYdeFsNCiWqtL2F2GJT+2pCjsig
SH8npTuya8Oju3l/mOji2PIImKr7vOKPoEOKWcw4uf04yVY3XpRWXeShpAdywtP5Bip8cIl5bXw6
1oNPVc2mRhep6G+usCcGwFhljM9KMrdKOXbHwNxB0r92bZ0NgCY6mBnHDxT91dMtTILU05IyBrn/
wpQS/eSCp3lQg6jJKdVzWjBQNPDBwlwwGLnoDXfldUzS3/v75Ez5d1LYiGP211EsrCxnB2E9ay4y
2HuSnoUCMixF+kJSyRBD9ckGnIibawyvr5sm8vIY1sRkARIzH8JeTuiA9WBWfsg5XQmiwukWkCio
SyTzetAqQ2m5g0tXBYv+osvI/nlCobh3+bx/Z015CqMld/MdF3ahp6LMR3LKkvNusLtcBJf/BCLz
CDA2I39WXVhRHyKED56cu01+68QiK6RDtksDh/fWziGu5PO4tCG2CnUzCzuMuLNpbmcjEMSb9ZMZ
XbBtVRV4xS6XSBfIkmcX6d+NmoFMXHb0Kyn4M3bSAaa4X5PK0Jd5Ug7qUpQvnSZNLk2Y0h8MDllw
o26UERCqnEH0PpsbLO2GAQ8XQvu+//vP3JJSUVlS+qehLaw8Lg3hFoMQ7oqaZPudHYhJibrf3QC8
FnKM+VnKOVlOGUuSmR3uskzw2eNLaYKGmNlWqGLp0ieN+xFtjpYgGryoT8fsdAh2dON618S2gLz0
D6vkmHPgMqIqQqg1qkRqFTYierfOIcBgWCasPhoBVxqsPMa+0nmhvm0s1l72BueFCPwxac6KXLUb
MmfsCXgazSgh6RFQWnsn6bNHcNOjWt8xYvUq4qj9Pj6Urvc1I16+lvcL7LST+sb5mCsitrUCZ5Jg
TF4a2H73bygxsRZK/4kjozDj0+anH0erW6VfN3/IKdtrxYwV4wu/o/N3Sx1erecvSvNO3nrPEj8F
g3Iy5l1qhBnIAiAWtIoTE6nmG4dWONL5yDx9r7MSSK4KOGsi8e8qdh7PNFHgxAvRcMbPky9Kq21R
jFONW3yXyaPkPxb6qCmp5w0JwGNZKY46M2/ORD8TBgZyx35PkFv+XwTmnsrJauR0kTPU2zMfAmf8
GOyfQRiJLtZoLwkJbBsIZ0q9BP1S6sb0qSrvT7EXzBat4/kHYsjAcI4qz2AjJwVpcOkLbsvErp4u
f1wtzI+7wkvcnj7QDBk+MYXVmBdBKx7x8YlDwjeyMTxGUc47P/WkWvkBQeLVMQkSj5D05Ego6iY4
QTG0tmN43DWqpYAUPA7l0xYLvqovjU4fBYJ+dM1epQx8dLqbxvqB/9hc7GVpS94jR8+hqFhgofCv
k+Q7VlPE/TO8ili01wRp4AppflXM3IW4uxyU7rFYQ6Y3AzUMRFf8hmChSIZP8afvKGqcxuhLI2kz
OsmdOEXLdnBIvbZ904ZOlQyrwYvTpQdChIYPsEQw5soIIFTQmCKyQNNFddmrTCipDXWwWpfOYgni
kDLc1OIDUaLIxo0jyx4a/AdcVhBGwhrFshBq0pXKgvK9svblRHL7Q9WwRYHk3kMMc9PNvVKJdorg
1P6nR4wgCHk5OjqvOFN0DtPNOPw6JKRCqFQCR+Re0NEvxGedQ+araxEBMToc5ctri4zUyyNWAVY5
FGjQgJ492hYfQ2+tmqjEz9PY+FYHN29It7tusuUkdyBfQfbMhe3vpvcrpKR3eTKDirD/RThDCwnp
jdLcMrfj4sI06VLbN7eUXshoRcfcdqS14VZjTb2nA6Fcm/1Xb1xaDixpze006bvojdmCMWR5MQ4s
3YSp3uAVIESpyr6LdzoeA7Qhw7oyMVWL0ft8LqELYfYJWxDwmTLcNdYRR6l9KAR0SiVmf3E2B6Sx
zAfFf07FTLo0bxP1ftsk7UP4DbU5OCzPByuaeS3yeKJMSFfeQwygJePorGQUI/2x3J6SPMtOATPN
NDr+p/jPLwpbNH9Cb1G4+cSmz1tWcI/SR7e1RDcCsos8gqPtzotR1vIhtf6X+cPA8pAo0MOonWP+
BRkF3A5MXQz9JpnsT1/XiZd3KnOTMi7BMsJRx67EMxYoXk+FcY+jMxHwGeOTARc3ENyTxBan4shk
Gn2Io8UfY+F5Hc6oSlHziOsSAA3mFGBaJIKqtWsw1FRiZT2hrY4JIh0QlimQSLj7akB//XkyMwMt
/P5HdwnaYxnvUVMqmZfTqmuLH8grZCVC54/8osOUu9hBdWMT59yvj2w+oGpPv1JXQB1baglfOnP3
TFAb88/zVNoLj8iOygeTPN2leVCBY4obBgtavA3nnul3UroaFIDQpWDE/Jsa4YUojXeyOuWnMXMn
nWLFcNkwS6UaqSHxD3PQVNrkvtedhdAWZ1n6ryRTA4opSdD/3x9PKPVWluY4YBlu6mjaRf3GkAT2
tUxtGxySBtcSsPRj+83R5KYeDufnWhsrIFG+54BtrnzYxyYFIVma/sHROFnPPkad/LBdVaTAM67U
sGNrTW4fsvA8D4eRfhMwRF4PkOMdkrg4t+21BCNktAaD3oslmAJsXWdjZoE+kt2y/jkRSmMIUQM4
cgYqVdtbgJDmKqCsnDvrvcz3pCGM1X3jKJH/E8thkwB2PNaDaTM0oX1ASq5LuQJ7WmFhw+CgjgsE
6biMxIvgBsONARP5dkh91sPLZC1xqn/9SdyIffV1D6Q5MqnAaaho4Cnv50IqLPPLMW7Yx8mFzJC3
RfeEqe0fkbAfwmgIpvMGG/PLhUSGTxROrm3HZ0RG8PluVfNZbZFXPPBBlLPV+SvnoclQz2NDOSSs
pHcjsvCimAu8fMHtQg2Sry6N4LNX7n7L/6Hnli/W6EkPuZ4PBr06IJwG9/pM2gdCWZcx7PeEX4mJ
G9adkcZSz/QyCyOvDtHcHlsvtzZDfswT38rU9jClP7n7+he5MT3xSS9niXVy/nzwdkFoMvPAMXFT
hYExio4KunRTi2mqFJNUQMO5RJLU7yw52w/Jc5hhQbhJMFwjXQOEUTiB+SzrPm5hLK+h/B7IAefi
DVqnNiB1FnpUOXKn2x96GYF9iq3dfKh9vkSKjjlgic9TC2ndrEK86GocdEKLq2/LVZrTBcIp1YuL
JXGzJWPUtlT4rhewb4EEnkpKLgH+LOlm6XV1x70Iks3cpPPS1Sal7d28Has6j0W4UT/ErwAejdu1
M9RdciF4ZdJEa+cY/TlODeF8Xt/bLx0wNzvE9QwfXSxDuIrMnwIHLNbunup2kZCUh8Wc5uHJQwQq
jjNbus/korR0vOJt8cAtLjvsJ2OsohWYoD5UXpsFpu8ar7pU/XxEsDxTKAtasMfsclyvqBJK5Zir
YAytUKEW3qBp/Qge5PJHcOANMz/VvUiq/yAqUc4kXChn+PVwMAxNPsa3//mGcC6LYAq/NyTpmCWA
nOf5ukbaZccDVIzXD7EUnJycRIabI/272ETcRaXRluCunFZVv4Loa8+bxgLwIQnvh8yl9+fbumYw
M4snRkoml4u/L8NCslFo0W5CIv0wE7WcEQjUX/I9u1PGPlJxcMcidX9JZA9SV7XSYXIbHgFG3KOp
QrKV9o3UvI9baPS5PHcsVv+X52sighpDBn2VWaStoSbZRX1P8S4qfVM0r5vrdS6uADK/XUOtFxIU
kMePcS7lH8EHFdAIFlJGqLOVKUW6YLopcR0NIHul3TERc9sFD6wia0cehq1tQH007wQbEfwPMV9d
38DGsBekon75oKeR3GjXhdHHJZKJSiWntP3Ic34NRe795UFzX/0z6VYA4HsrLeF/hJq3qoymJrBT
D0ETkzN874av7aUohc+OWFdTXKg6egoAoq/YPl8bMeqVMeIBW/knav4ehpPePexHMzzdAfk2CnAA
zfvug7nxaJ3NL1YMktT1svBnF1acir9Nm7BILWB/e++aY7haemW+zCIRuIQdSZz/cgnwn9fYqmwO
jzoi5CMdk+byatxWYlqVDE0nFuABy9WGj2rHGlWsTwlSCPup7WgwvgrBADbCQeZpW4kSqdThYz1e
6M3SWUJDl/jnnKfknrg8LEbBdG0CbEcR0XNZUKbCl5cJJkMUWGUFVz+s8VfbKB4fvjoHnaNfct1R
oPO1BwOUtaZ0JwiUzOXc2jxhWI/3ctry5SUoC2Dd/rApK0f2w67WnvenC4D7nbD5Kg0jRqdyxVK2
nDXQVfRPozTLvtnCgRaiLYde8jdh28K9KvyZA+F73ok6LzICkxcQ0QSQPbe2nzhkz+quQWyWDySW
mtWPLEXd7T4H0ZEcmrY4FTyQCMYeOgovXJNU2hPOJ/d/XxPcDOXdFgXN4avj7L50Zbao2EjOx8wo
22nm/nQF164fALekrCkMhWiKekFhPw/9S3uMHYh/yBphdkEVQXK9KHiXU2Dsq7vqrdV60uTAGTFA
cwqfuWn9BNUjV5SLjKmnnrT0ZxfNXqxYnaBaQYUtLMZp6XnFzDovtSz8nyDtdKPfef+/xtwMvAZX
E1cWH89/S9zq0jHCDPqqwNkK761AMEmirC/SCg+xhXYmUIugr/kWHKyEwX0Mp9wtrKd+ZzxU3FS8
TfeP1LtN4MBIYPKpw1Hc+mRGlfE5Z1awWMqQ1+7HThCocnP8jizbZqazqOV51VeG47zwdskZrdgf
A+wacy5JACQlZLvxG65zvTk/NMWfX6nldV9cv6fohFgkUvJVRMompHqwGxm8YAP0bx0UreUvSmBq
ggzM3bRF9zFl9gWsc2mcc8iADydaME64KD1yq/GOxSttVv8x6a2LCcJ5ElMeZalDMkIt/F51gSNb
dnxwpFizEKT455eGNAbDYPUbHUHCJQInyfAyF5Iy+bckazVKw9qjyfN/1bTIBa8c6LlVlDuFntG6
STH4vZB4X7G2/uCPnJRzuGEENtqt9W0aXgdM3lXOmlpAYO/9nP7KJmCvI4eBJL2in0EGYdwm8W+0
ervoBjZJeE+aL+GVtHl0iqocyp4ZM6SjRS57FutY4bQ1/9iaMxXuJcrQmlzngQSDDpdq+rCsfKRa
gs2PSuFYzWo7QCmaIJsN0LvB+Y26VoOuN65KIwmyVh4fGtbEN64Chn90ED8ET5RrEOf4o+YY5L0y
4kdBrfkh3oLDRtq1ZmyR/v6PVCqCRytMbz+Sn+f/1wfGVmcMQ2C/kT/JJzbbF3SMvgx0mBSMWP+R
rRgtXSZF5gdgv5MMcvGkP5V+1WHcoOBuXzulpAJFmKXN2gzM9roZKBxBTzOeDhfy81gJJ9FfsKpt
njM/3qRiShFQjrqFdGFIpFI3Eqn7tQ7NZ9xD9fX2t9wZEuI8opQ2f9xw7SoDQechXnbYPIGbGfRP
LRDK3JZkhH9hMukjJPuvL+403LnkwE8F8RRPQRMOwIF1RxvY1w9SkZfcmhJPChU5Wr5g3mGnnxiw
GCn94HdQxw5w3ukWqPLosRjp0W2R4qP7XYJ7ZdpvpLUfDjGTV+hYHkcYdpsq0ULEKI9czhUOfL5X
ujFKVRaB/psZn1pighf4Tdf90k0eRtCU4Rp7uztvwVyWetpRxMg2mttJlJVNCywdVn73Rdubztor
6dH5dnKwMs39oBAB6CnyYopPh/LetF2Tc7iaORHsBJ7whB3xqVXur40sJ4Q47UVbB4lHoBM1Ratn
U5CDA6HU5kLz2nYidXx6I65FTODqC9SvOWUo3CKVu9Jrrsv+khLOR/3p8eXPAs5CiCsDbp0VKhSF
Rc4Ct4YKowwQJg0Sm4ZbShkQRbsUroEIayJdK/qt5HqPWQRZBxH34cQBaJi2Tbs/elAP/OR3Vig9
8bz9/T7upw1NnTwJaDmMLXdh6xaAGROh/7PRWDPRUdKMKNWJAuE6m9M4gbObmG6JwNE3QOrrnjNl
A1/PEnG71gaOWUgcJ5Gqd3dhV4KHFWtsj+tvcIhJknlV53VrK1Zv6v6ZcuhXonWFEpWs8mQ8dyAE
cQMo/FHCeovCoqCuBKPf4xk9kf3+WpadVJkDJpdZMiByPvVBndiu9lwn3TPrjrhoH54xMXPd7Njb
/s7CjFHv+Rwj5CclRtpDdEsncoTFHYsjfHSgAWwUj989gsocBEOZxCXxFrUhZxWhdvHuw+lnIHeJ
hxu08V+WUtc5cc3VfKUXQG/ejX9DlSFv94HG9FivJBWwnK6bxM9Sj8d02sN0iqQ4HrMUo8LQnBgk
YC76BAisAUu0WJ3bSIs6JdqrY9Bc3BpcS7zvq3chHMobNMk2FtbgVMDuPR81h8XPHBNFO/oNC5Pz
vOawlR9Px0nC9nnJwsUK4FC8pW8eEK+e/E48kOSK3DuFooy2zWG2aV+DEIqYdT/wZQpG1cl84S1o
7mLiMTBRS42Fvbils1RJXrbpTnlzfr+8/ElkVlf4n0KmMSsRjF907seZ0Ia6RtovG6gur/RASNMY
p3gCSQ0jHMHFrnX8osRDzOKDNBaQZ5s7nGVTyzZAUGarq6zECUBOEu+0Ukp0jhQJ4SarKW0GlyAj
Wtc9geCDNGDea0xIN1CoOTEwQSZAMKvwqCbXGsvFR4bMnPhrEl7sKbKKoreAnYMWjeIwIk4Oyq/2
yEevxgpRGCReeRMMCdrPwkYevVUrFmbCIok5r5+NaU6tkirAY8Ni6VJW9XzF4yCt+ZNAgI8Z3wK0
5BdpVOEuSfTzHVY2mvhIJ1cm3WzmQ+G/jIVYT/6uVs9axQbuC2NxuUg3PSE0RNxchvcg2T0Wp18t
bK9ySumPR69Ch6sWIep7O9IgId6S/MxYqLgWeYyfWC54wR8HEop9lbBnd/JoLZDGOqlS/41tS0ZJ
tqUnT0M8/cm3Lqh5tYOM9NP0mzBiALrsGTMHpsDtvVGWhYYGmAbbkoL49PkTtO6MBrRY7Kt5PKgC
tb9Y4jVYxdfsMf9AWFw5YW/29eJal8dkmZObGKaib/eU+XzAN5BOSam8WQUQftKt705YIdy9g3Ud
xawYalAC5psJFbOlIBQm/T7Wa7fiIbX4/WH7NgTrHicIPXoHz1WqoS0UX1H0XbCU5GX/E14l2XAI
bQnkC55RKiFVW1tQN5daZVscL3TZenMrRrXacEzzpy8FLBhsnKOQ379+2cKsJgmKfxucS+ST0c+s
VlxojLUXJ/tZRNfXQizkXvkaSd5DWPo6f32ZxbLbb4MQXm8rULfC/Fwy0/WCFWivC74JMfBhcsng
6lrJRmtD8RyVDtEQ27Oj1neoNFderOiKEYQJxBm19/KlB43/UHG+4qfkHA3kqZwWctr5WEqGPfjo
3VL5U2W/+dV/N2yoQKTnyDTka8mJ1qYoVhp50tNfD3qc/zbe07ZzyuG4ibe1YTYetDOERtk81DaR
b19qgXjooJiOrNwtV/gfaDdhZgxn2A6YgXMwzKOj+ham5KcFSU6A1TS3Pqknc9zzELQWt+soTZvN
kKb6MKKWntX7x3mJtcCSX9/kYZfk89klLfMw4uOeB6AozU1OOV97ndNI+h6Rsn2atDwLyiedIjYo
EsEeG18zr8w8V0Gk18NJoig/jqCWE/m3VD8rtLG+ob3Y998lyXR5q/5Wv2M8bXF/bfRehlyP1wpe
f22xSNXIKx0mAHcQmTbcdAKAG42G91xcNTDw3/jvprOvuPgQ8bdDCTtaOlVIcxyeH3o9YyZRHvP5
/s+G5GUALGc8AyeGJl3THgfSuZfFdT/tS2jJKr1US3ycqRUfDZQap/1a2cNhLPcCrZ7ExTdtPPMb
X9kEKj+FQNwwST49fTJi6yPgySfpY3MYMPHofXtdDNZdHOUX4qLuqteotNFzpPw13PLaG9Fm+mqt
Xum0//OoWRvi9U6FlAzmNmXQWJRPoHhYQ59L1XrnSFdPX9ohydHf9b26QPpBb9vIukZwmdNgUNQ3
uHk4w3ELDikDwQj4r0lK3jwWDnfrCXM+WndP4THritrc5oD9ELQuUn0fg07b89FwpDGpcO9t5grt
+55Wht5Qj3XCOBPYaNAF2CmXNen4kNkcjtm/QFnfK0VwBa8LX1cljsjzRHdhWCkA/JRRjMk5Z+Us
FAVKBQ7RaTwfvFc+4ZlAfKQ2kstDfzBj1+gkuZUs0Q9KeREWD2lokePJsKVoWiwMlwGWTcGrwWKN
jIImto+OZNEnzdKQmShfOeV1Ra1CeF8XqyJfrmxupczPaDyuEvPGlGamIgcBMTM/pax2s5QLcdnh
JO6W/Gj8q1BD/IjYWshv4VEncYREt9RTChIPpcT1Lzoh7oVdQg69tHVojOridx/9XeD7xnPj4MZ4
6cNVj+srlwA/JY5Q22Ulh1IE6MHUsdjvDkS2Z4Wy+SjdkDkPSU4tvuExzF34swiTfIVuu4dtU7Er
MxxNkUbgJ0bP5apfVu0SOapqyyVxrLzlT2KvZC+LWpkR95L/X7o7gY+nq/uBVWwU7EMyWat9FJEo
M2lFr2Mo8+yB5g6rH89Q1zxsg0kmIO7mVjzzmwtCxTM2iRUZPdhDC/yksPew7EU5SaKS9U4a5EEW
wodSmC2vVSuCUcLFjW+Co+WliE5yoqVJEGj1bgxefUgnlyjHv3E4u47iqO80Fav5XLBE81DhyFv/
xJIyAJWOS9QRpErvSAtGId3ik4p2z6ocXu9auXg/GKE8ySowImOM7Lfhe+EtxiCWbv6oVqpZ0Cmh
R638u9WlIsKotuuWl6uyMsJBCVqSCSWLkcTQAS+fljJo1Xfggbi3HjWmN3wxDwgoRjd87FIxKCGE
G1C5266md7fyk+ZlRRiq8PvMgbGbbNlrePWv6ciKDBOmhkQqNYUJ/zC7nsL81FUIAVhSnD+DJIPA
pFgTwHvzrvh7Qpq9fRMTP9hnID331QgcE74z5NPOx3JuHqPDanaoSfS5a2JKiKvHTw4SyKzqdYou
myTx2sM34YwABkxltEFldcVaDXzaI2f50ocB9RroZgxdn2pGC/6czMWcJ5msuLKdr+pMPO3JuSw6
3zN44/Xexi7TE668eQf5C5AMdShN2BLtC9bDP7pFMzf+ldtUbhLLtqPrECObOk7nOF3Xc9/TPWD4
cdSvtqOJt8aFk2Rp5yxjig+IwsykyE/kEFlEgax3p2M3JOdiv1Y2LJSei4RBUSqItsa51bOEX+VT
pqRdHII03+6Mi8YCHRd+cxTW07wi+J96mXE0rlAY3a8Il4RsS9xoB45HS7HdfeVgr/3ajrpqrJq1
mYCZYtWaxlGdhSMguIebG8GvDmYhCGiDdrVAzTosFx3GNKMcsd4nAWdOzQIAvHpkf/gxYdpnXPtX
wtELVupYC2V6WQYBBSroRW75+/Al6YMKfNdXKgm1u3dAVQyE91U3rYlKyrIhD9Kpx00mcn8eKKl4
hOGZr807TxMCmHeeHFrVa4D0NRdNkZbQmQPCW/l+xisIu90oSHyBF6SmiYPjPi1L1jPn7MAraAsS
QL+kXzkD9ljM84qXB5cKTBlFs8d2ifJbZei0u1NGgQn9SpsJ+wfM1a9BLQAs1HNqqlTWFErmDsUy
DC7UNAeDu0mDWG8Bq337A69JT2bikiIK3E/m/m5tN4oemwOOALVb3ccNzxfDhDdcw3B7J0CxN8WU
BetcYnsE93+othpchh6bSotCUwVYbsIRRmJ6ArkZ+e1klAiNjV2QOrbgf1qaJviRxvMnvYg8OmJ5
TGNCH/JUQBe/VhtZa57SW2G65vovI4e0dgjDeQc8ueLKv0C6MtgC2geyyiy7b8JI4ZIAnFdKxy+G
RQWsClk9hm56kdBTd8iIumQL8j1RrJ8rZ3fGrwN/YubVmSM5YgjOQup1tP9Q7LVkb8fFUz8LG3rf
jJzdEq5QIvB0sPgaFzkLo6NlpZ2Cksr/PrELvUZZApGaF0sndHqi6KQ1zVk0HcnWokpekj4hX3gz
Zz+UxkurbyJyuEN19tFkf8gILSgXnulpJeeyjisVagvIMWGNSssjfZaRVxJQ+SINroCvJb5aliDQ
dyZjKhpJkeKXX06LecjZNyB9UhkTw7wh1DZHkUSs/hPdDS/UapVA+t0k89RQ+fHFbLd2z92D07Fj
8tQbSYZv0oIacV4N1dGvS0aAM6xTfXYnBqOeS4IjgcuKh581iJpLE5Ro69AM+Vekih2+LCOOPeGq
Ak3RqqUj+7W4lrzwmOXslXez0gZ1PaFuYjmCxSWxhnbCgzDTNwoSNS3MbmXndvXcoRwO0PCkG6iZ
omK62UyrPZvLKlgREgVD8bdA/nFcZYfSpMXub0PakFPDEkrTBSd0F0lXSpQG+c6Kc0PUvXKdy60l
eop3L9CYcWJHTzYJlMREg39Yutk4iMsv5BI1psYbsIK5J/sncRB9LGme/AgsiKDMcKHGh1GzItgH
DlYN713kw5zOCE7LLwrHgTP6xlOp/DPTf0PD0mSErAAY3YPGOGHN7DyTUHa0cHM6jpUz6sq0W7FS
v8hK9cBa48PxEUtvaE7jk/m4aljLXxIEeQRTYn5jCwoNnHvDyvBquEo+mjmjsrtXOKfdN3r1T2a1
yutxUDtYZSROSOKtzCkA8ZMCcUBtZeW5s8PwWBF5Z/HwCMtRGJGLbr6Nf86pyMSgNhzsB6KU2hjq
o7rnPy3t/gvuvAD0WnSpdimdDhPK/2nI2hMCFh97Hp5nMYYrfXcsyl1UjRCtS3nuridU3iOMV2ff
eUcphoFXR/34jY8RqL/XSud1m8w4L0eCWlii1zlIa0VypSWg28CsmJsaChqukKWUxDZyf3KWTaQi
AW59anlctTEoRJNA18WuNt6fEMHevkcNJHZVZxdoIYl9/SHmKTwPEX6skfUlRQM6CWgCpA0TWOyP
ERHhKUhOnVjUzj6GG2ypv6SPgzU6/b5nzod+4uiKdM2yzjDoxK1cOgLpG+hoP0iAejEdR8fkpHxs
tOssD1CoNR87/38hGRew02+qA8WxyV8Uj9wx4ezbzIVBUtuSWiwE6RR9XW6sX+NFrcY7X8ACN+Bt
yyFQj3OCBvY2OThtfQzlnxcSIkAVm0zz/UNLNAT1rdNlXFnwREadpHWjVSj3rFbfjvlCW5rlpq64
HXKPKg9hGD1VD9fnzVccAvDZYpzeE/PTqeT2VDcbMOcuRSvyMjwo1c/PZk7sB1Tez1kt5lF7XmOt
jUyGP8R6mfqor+IgBRXuwUbAr6BMJuqIGvRJsiDjAZEY/zpzIFd/0XAHozpwmkaIu7qMGZeW3s9w
DAvYNP1RM5kkdYnBt45xj49JGbMN5reGfI7CJHfY1Emvmv4VJn4ctEW7+Ev9Yh8EakemniCAcs6z
NizsNrRzvkDLMvHy8GAUVx+kRtJgUGZbS9Spx9ST26rirjg/kYc7xy9mpFxjsR2fjHmlq863IrCJ
nZNC45PtM46esca4hLqvAbIo2xVY07NG3ruryxhYg9l+6Jt05NGRAvRm6Tfwu8DOhieJ9tMBCjat
0Vbhc+PS3RQqTQ/o+AuLmpJjYfoeoScvK3oqwRYTEBVQVaZCyDf3msBYMQwCIUnmQAFsJv/to5Vi
nzseB433u9iv1neFk5K2WPFgI8fKAGs7KVlTizhWt2cGaOlrxZHL4Xd/9wNpzA0pTo9rGbUmWJK+
DahhJgc7jBEQLEbZh3Rntv74rf1/mySiMJgpFjPXBHls/xi/nh4SkZtfKsu5/cm0fDJAYE9B6EVo
enEKJKEedNqVubFcG2HGkjfbTLu9TQqJeIonWbesFYmBHWtFGanh59jvQrkvVBHLjCi9uecjsGHz
W4kAdUTsCrP6wFFKJorxeYKit31sLPcuNorCSCWU0lsh2Wn3AlUBFIVUnn3xm+CAV5aE9BoOsZTb
zBn56tWja8J0a+E6QXUZPrIAUNP3V9E+9uM1rrxwQDZKTrrTe4XvngdKJ1dM3pQtU3KSDeiKks8R
DPCSzIcnirJR6B9f/USmSv9SUeUZJFZMIt5tksLZPd9+Md1dAsyB5aFNfrTT6vsI3ZvkYxEmwjHW
+SOX0bHFZv/fuxWeWroJ6yk1JuV8QNbLjCH2rZYuE0Iy6iGpjOItwKaz31ZzAEMt4+NiGWaPh1AB
9XeoEi8UQbhYrSfZ+7Z40zZaqDAUINPW1yPjsuQ7frtw7A7cnEJmut9x8qrmBfKY3yq4LSOJocR0
TYktrC2d2LpzZA2P7KQfQpaMbdrN+h+tl5BDk7jkOAcOS0zdqBWS+eGDF1S1/9nTCufFyqM4RBtc
64tl8M1CbTLeTX4CUeBBJBIc0SIc2z37UJ00EI72pNZtiPVFg9ajziRzryZhm9380vEz2BX15+Ys
op4n9xn95qrYL9MZKOjYHEpf2yGdeBuxxdj+EAkeUpU5wE4bpdTA4AdPNaSR1y1VSoO8TfE9JuAu
weAn3Q4ni9RbdqKX7jmqTJNIIQKWLb+f++9gXpTwxXE7+GXMvUdXOqpkPybKkOasNiA07rNgcGjx
Q/BW9mB4vcDCM7HuQnD4TBLVyk1nm2BxLLwBFG0i86L0m+JuHoIxqc4t0O8RzWOi8ppn5iluxEWQ
S3YHMjY12/I4QMu0YRQV/HVFTBmfIJWEozxK1cBpqZ0aJ3yWj30rTMf2MOD6AlR91VQcwQYZCaHa
tvyxWZ5xLBJiwlKXRyO9enuZ3Q3S5r8JEqONJf1Yhlioq8Dgt9QdLMi8pyVJDSbdgMxSNpZIRl3U
MQCQjqgZ9EuX6XUMUYTQkKBpvGlPfD4ASUNHtWSTBEmbVdHWtjLyhnRb8DfBU0Y9SFDPE/D96zCm
KrFte+kgj4vKyO2+lcJNWnTxRKNHCVYt8q9DBADtFW0LEFk16zKSniV4a0DFDlJ2ed6feR5u9XdI
/VybuNNnlq8w50JtveA0H4luTSaNC4hv8TQGvMil/LNZG8il2mj67sdgQexakbLoVUA0dCD8gXEH
oONvmTDW2DEja8sRy2Evor2TpD8As4y49ulvg8O7nOAU5zhHRfzXqTelnt9uguhCxMIiqISyvf1u
ZvoKZlGZi1PMqwhw1IxhllBVf4wD3x5/Elc+7J3305QnURWRztU0RNs/6OFGymfzI4fy+Pfrjteq
qWTQGuOXJI8DMzQBL36HV17QjlYgWRV1PFe19wcUYkmH1AoFidnz1fc3c13sUzXF6Tdml0b6Fzo1
GAL/0MKjI7dS4dacwWfq6OQ+GKtx+h1ILgPKrzMCd9RJM8uuNc8pcuGvGNvSGyYbcfT/NQGpIMp0
wu8GAWXE+Cz/fd/Mpf9oaDZQVI81Fe2o+yOkw1aydz4vlwa9hwgdsvHSJGgIP7bhj/l7mrRFglG+
od/1kRjWxcda5E16JEGzjir+Oo2Q0wwmegewi5jVHFh4tQRpnctXFD7ubtUbImYst2B7YT/9iHIv
DkbhCLtWjiazd/KWRfq6DC7k/m7rGjkJRWKMA5K0XPngek8BiUldWtPPoyoXXmBTdR00H1QfyofK
WW1UybhwYnRdsu73AAv5j5skgfFNAOljgFgtVS7GWptecRRB/al018p8YDwGRE30aDzkCMMbcoec
do5XjgBi4xm7C7Df4I+eBcb1W5GyydRwmZ259BaLMs4BKSCFrvKPz1JAiz42tCGGGvd5h97rNlJw
gMZpAYxty1Lc6H0MWHpR7OB98gWyEE5X+0fq+PNDIlvqlH0TKXqKIDf0OdxxNNi+lVx6kcMNsbSG
2J2DPT3Gd1cSmDRyy3BV30MC49qqqtUlh0hMIwHe6qWvvQ3SUNIplkps51D0Y32yPr+qr8zAkw82
7K9e4rAD1lEY3ooxbe1GAohE54uF88qKOE9jIDC5Zpn4zNb0SBcYnO0fJtcr2o53QThMEx0j88ji
bA2f3czEsPoDVz2MWZ1klGaooSTNWrQLjM39mHa+fywtkfcBv2WOS2CWDNKzCYFjP7Q/++wy+0GX
ld5sCka7fCcQwqbWIhJFPKNbH9eisG9/48rT5ONLQi2UD3g12rhXUCUkCgjY6E3/n86uNqelm7RS
Xggb+Xe6bb9NMldnOk+1VEltJkq3QSohY2r2hH/ddHlQlEWnsUXCda4j0sR3+pYEennpGlkI9C//
+lucftMXYlRmsKAKFRvKfnkm9p8LF9zi2bmi5J3AbE8oWJ30o5pK3hBG8dRkMefNRNgoLtqN6LCD
gLh1M20K6BtCQwrYn1Xn0pHVuFeaIxE/IPk0lGjmpK9dGax0EYfqQU8Tk8A+ujdeRcVZ9pHSoNF8
DbPcsvHLl8mfdhDXAcV6FpxfYxfinxGLwobw3GIomu/w71WYAgdKWRY4esZPMZw5aDyTXLxPeL95
g+nOJNAT8bAobgLi3Qzqj4wxLx753IKB8Y5uBL5E7SpfSqeYhwqrEhV2t3N06Qlr6mNzrOZVxC/a
zsbiJ2NSlG7XpypjEbHPo69NUiMdeT+0tXcYBhuUg2sc1p5C6TRToCSO046mvKHsZcxmMr7md9nL
hfuwcdQvr2E+LVPu+gN6P7+eANQ1IP/VlL82vViL2/wPvJWmWpHmHtQ9ZFc6c9ikOyDIBdTHYRW+
Q+CDCszeCzLCwupBs5H76FwbzJrl8QB2CEHhUK9/+sLikJGROg1Ld+cbrYyMN1vPCYgmZmpGYfyC
Gd+NH7hpi1MuvDIEc/2xhueN5L3DpePR5B2VOKcPp1UJ2JtL71lNinzMlT3ldcSrngA8kwplueny
ExKUbHmfsZldtRM7u6Gs7+ylLgeUc4ES1JurmiTi7kyTxeiChN7DhSpQ2yTScSxR4pwSapMXMSry
02uIX5tUJFQwxoP+cDXI/UFlB5MkAM9mpqoMJO/nJkT8YnKLCWSrKdQvn+B+pa2C5eDoDltbHwPW
aDNISlOKddqPzRhGOUlbgfY6u/C4geZGbY5dss4eGvXXPbDkLaLCpeuiNfh0lSEn5eWOUOtr9SRv
1EPHgxWrLyH5HSUbrSRScnpgdanrkCSS6gmw0zoujk1lmJ9LUh/pVCBL7hXZnUhkKC65NhbOAbAx
pdQsK4JqbBT5tTahCc3BcimVvuL8XtG3C8fujNg1MIDjohO/roz3FdRPXJr6dsR8UZ49MwflCgsG
6d0VlZCTSr2WxkWj3aetLOTzJ7HTckn7jqLcyk0I97OPsIRiO2blflqu3nTN7tDbU+/8p3cRoAPs
ywClg9nI/q9GA/xaLoElpoCwY7wRrkESdXrVxD4aQr2N0S90uZvipfUwDmEnTtT1ATA0y64eQb0h
ToKznpaQdx7iYr/4ms1fSZdvgOXWtlp68hCJKl1CLt7t1UlsDQ48ZMh9AMCkiyRw0WJzzB2Oi3BF
Mri3L/raA42imCkCEUluf6yOfAudeth3x1t5kTFJQyRN1IDPYrFFQlQCdCO0bqbveSddxPO+Iw5R
D3u+AyxDzM5kIxzjNVnkgH5ByAObS9kNMcjHRe4BjLLZLaawRRpDKUfRm6A9IlNQxZPVkPhH1IV8
eFbMmcGXxTj59Xpgm8HtXszf6Y9fj8JTtGO+VCs7LVOlE68Kux92eXavoefPm6ALrTPdY5bxIt3j
sCBKecDC2yjk6jXibAchloU5kPolJRHIqpDMMGHGIdHhDbjkXwH2YLOfDpZWlQ+xvniOy6PKif8k
47g/cRGh3bupC+wJ6DrXUhy5loIPZNB/O0SJMRffIZD5EqgaNqbQm25pmsGZmyxP5eVoY2Rgzn6J
C9NATB4UPrQ/0iMx1fAFtIVQI4mep9o7CU9kln5CIl543bgqIWBrzijqDOqo8agjJdxBMbWEcpfP
6wW5n7yIbfc7nvUyE46X9SbVwvK85qUx3TtteZiLlqSQnVdd0vV551nHnAKRzzP93tIkjraNwtsx
UiHSjyvwUpBTyZq9nE+si2k6d+9uPNpyW5qKWXbWxaqi/sAmnsk53JHs1f5lU79fJ5Wo7nQKkuJv
2qnAvEJ71QpbAPXZRmwA7RJnyIcohGDEE/NNMgvAlMs482qnwmAf1WTrhZgrFrD9QpulZ7zQW4VM
9xmK50Q5SVridJE9MV5pueVSIOIxc06waoI29T9OY50xyKFbCyWXb+JW281BK0U7xj2Ue7pQrvbZ
ptAdXFAOpkDg/Y0M3uEHZE9uFEkOBvgh+pmVTtkJWdnbfcVhOhCnSWAQesITrjDRNSD7E+rZZc3R
YWmcJpE7g8L4QpPbtqLXWMDQU6xPMiYfEm1Jxbe0AlN0rE2iAhaRuVWySjxvK1PZ/SH5mb3hd94t
8DJ2XrhrzsnRtS9Iv4hdRJ9Fw33RrtnnZyZ3wfum8F6rInrrQEOwfp+VRzG3jSuosyJl+C49JCF3
/Yny0dK7z1Yoqn/HgFY/jHSwDamA2ugymf+rL9rnFws7jnFCrJt6byN8+OGbP521DGOYLwpEIK0V
+xka4Bukp5YD412fSEMxlZEWt6JKuDzs3i6RuON9c13WTbJ8xmHRCPelc7PQwHiJSd/KRQWFehaj
uE2k4ZBsZXvzFPCjlLmaA/NiruZ1Vn+DXKGJFGPEwyukPD0rBxBS86SYVB5BqKlDVwnR317c1627
AZYX6Su0X+HKkme9v0CjWTs6VDd13pNv4/aNSAD2InynW/rccCeYVm3k70ZZzwq2tbVXtzKBtgT5
gMLMPH8NSJbkOae/j94TIeUIZ3a1EsM45nceXoAzT1ocdGD7gcacLd7X/Rmn4iqj+pRfk7htzVcU
PjPtWa03m7YRUZF5+3HlWbc7SErQ6H4oxFD/07FPzG7nf033Bp2pGttvc6ozb2a1Cob7gB6nW1iK
e0TIGeo/SmZaJ3yRnepjwOgmNUaIAzFTJgsWLeMONTgOroFk486rjc8Kg3NhwP/MuYmw0JpOPCg9
zXEDPr5PY65CuVh2X8IDBlQyH/5jEG3Tp7MFaKDgHs+G67IxkVOG7umH5ACHdUeUErF682y3u8Sz
w9l5Qp7iGB/VVLDLB//bN/WU4NwBV5UtbF23MZWeop3X0Xhl9HxZ3hjF3saQ71ZpGV7HRLFBhafE
XG3cNiW2AQF7+11Mm899I7zEaMPJUqQiwEm2n1oKz+qrEqi0RI+7LFyA28sSVOV7tG6e2oqMJgPW
JfQmVXnJqsvYJ0/86mXfAe/DMxGrP845m+JVObId+mhKpIlmFj4/C2Rbd+gFc6JXJLLaSyibj/zD
74Mm7l4ECT7eol15CeB9llP5umGn46wz1KQw+0XjMb8p4aElWC041QeqX3fqk9M6XU1tW2EZaHj1
f3LkONoO6k975Oqt3xdDLRWUhLTgBSrTpuGOdMSmWf3fSzBGJyTE6ODCm6GsVbnySj9uGzW8k+sP
KPNGKJdnscAgWRPLUZAdMJjJo/kXcNEtaizuRq8bekZi2WyLtKu24KIKbsaWi0QALaNYqOz0qG2M
bYIpU1+0MMTZzHLhUWv49WWhUSCuDhIsM7Q7aiVjIFnyW+6YFDxFFxrKilSDAbaT2t4DE1H4TpX6
mCb/CHFVDnVVZoF7BdfeyIfNVIFC7umHUb8G3vOgae7RN1a5BwrZJw2SzBJOTkomvhSw+siHWHwT
XNSqjOSAHjyTflDFEfAgh5T4iuv9CQJ0qvfEu0r+a+Zq+fbO+CuwDc7rKT1DyTqn56IKwrnYB7oV
8W/raXRkYBAAmRm4qMJ9yvfKNj7g0R+QPDUbKXJTEvAE7fdbY1lK5cf41JWQh+4mJ/3yyxcFMxOG
sAyGWrHcJJUaEleNIyOfcmLAfgl/QC6Z6igg/i0WRNZz1ti0SXXDZXI21oKxZdfxMqrYlwVO7jhb
TXuAOYDeY6N2nqaQ9CD3ImWp9sqIw0feyEbgdQiOyWXbZvOa65f02Sso69DaDsV7MlSsABF8iMu1
VGYwOtxnsXAgAUCfpTMSM/5tetbZRZcoEnEuBrL0e35ba3F8dUO6ASkXLKNZNoha12ji8OKpK9Kn
OClxpX7/wScGggBXPj2UTXFPJKkeorRYvcfKY+YVCAbuJeLJEnR46UeXaS/YbB2TAG4ZrZhYvKjD
tBke37CpjrbFPJKGHePrEUcLTKczuOD6mPfAJupNV6/V07deBJlnbIrul9WRmsDavwzLhGt/6YTk
DqFzVb+LUHaDxAt8s2j8rYovkRjOI1fBD+CiJTIMbMz5z6tZYi/dYqEqoMYTOQd3Q4Ke6Q+TWbo+
Wycc6AdXCP4Xu5EI30Lk53JwqdrVm0g5eqlzpdIVRysCFyPtihyXltWRaoj0i+XjdiKfvNWZz6x8
8PEENG8t83hhzYmpKUY3VemrF0pKVHeMpvGX52s9RPSFyoP07rGR/4wwofoOKF1XnlZPKMQUKc06
uRucNdYaZE4LmCpwwcWPcZQ0XmUHW0kj3nP9Ew72aAhzvuy9VNzyORtHt8fd2cF7La2VrNC4QG48
Xc1zSjJEQm0FZP8IrikrU8vAhReZghqBb3RdcqF7uxK5wHx3Xt100yctAiVkOG55pQaehXL2wPLY
xeIRr7P/wCX2m3lfBJ9DjqqzBZLC1p5W7RnuMS1hBjW0Zn2TVJUpmO1dMto+WX6yXpanx/vwfjy1
QeOLN1k2xFryOs7aQbpA+AgWcgkc5B5X3mx0s8+qIkGwfcE4Oe+bkmGVzNz0dRdLYDTPH2VdzE3D
SKVQ04Zb6PruR2gfmOOKzFua9jx3buSKDndVrw9fo3TqsCdafqdq3ZopXaLd8+4k7KIiphTNTiDE
lzQkCGbRXO0l3+0kDRMzsiNCFMydSsSS5xEDvh8lpejRPkdeLkez0DeUg6P7KBAIOUlbwxkSP+yE
cjlzl+QPxHwwo2s6M+cMgeBEsLgstOiO3+G+icTeu7betRIdCdJ7q1dFd4gEQjnYuM+obmJfZWOL
dFPsKoIHddUhVf+nMnIBKgTDBwpfsIM8YOe4AShS+0qYKTJYimRR14dNQQKoYRFuRmJiy6lrXlSb
qK11apn5cbSinveNKWKdV+NJ5lUTK7+Fjdmges0bMYlyJqvB8BsVFsuuYudYf2YLE871bCjaiMkR
W68liVIEe+EM/dqGJRZmficfdMRGgpEwgS+EwpugsPeawvv3HHR92po2Wxj62oe3NOukasSLCdmK
4s5OlHWu2AEsadCIuWcivjt1ZUzXYLZkQs9PrtfnPLFdEXxJAD+1Mu0MWi+F+cPYYfkWeY5DIsqq
aqV4cvjVcVLV3zHRAkcvNePSFnmnwZp8czTscxrHgWLrwOWpX9TMF/n2Cns6lwbhpBx60FAJuZnq
iGpB5Ni336hteBqjq7vkozaYaKAcBPOUewpa6jccTmM9KpiZSXW62h1s32I+MqOOnKI5i0C63Bw2
1xp0FitIBThGkvKuW42bUi1JzXzxgPAJXYWXRG2gioalU1gonPyVYIosBQi80v2Pg4CWxocnFJw1
8oxdRs+vroPyzAnT6pQwZIJ3yZeVZZqGVdainfkM+w/1FBWQYU4KAA23KbevdEZvvrevZHfAt52n
Bsv2MYBTzitTAvdVDv3OLIw0S8ejycqvScoYaE5OuSoOL4EpIiDa8xs8n1ucCoqLteXvvUf7DjBk
/+37l9q4JIeeWfMTvD/iXXtA291HMk/3zed3vd/OfxX7bIcAKwzDK1Teru9E/+MG1Fig+0XkddkK
XVb+fMmgmAr2PfakhXMm0a29p0fsnh9KNdJYy7PmLaVZyTBSfXxrKyvAVmjt78H4dEjq2ce3M3jC
7oa53FY+YynWkSyrgN1PKHaho9XaopYWAe560owLibsYBLASDrknrUBz5T/TU/6psR+Ni7T/X9u/
OhFWgpyCoPM2UOrh6YfbJjaWwk6a8WUes3vUJ5xJxSBjMy7+s9ttSWHo2jpsB7Uv684CRjXZ0cV8
lmubTWXERSzb5ORI4iLk8Wd+M4bdxOC8LIT0yu58wJOTKaSmcedXCtSY/GCNU/8tgNH7UY+ZTK/z
L92K+jm0Xp9PFtRG7owQ3p0TAvED1YKkydQAKqAlEgeyiublBg+Iqo9cr5nLpKBn33gThKfF+O+e
L4L6zcIamWjIiVSevKFlDUvY6nwnyJhtYyjeTnqTWYxczdh7hZj80RBSMOD10N50McKX0lGSDma7
ulvpdr8sPw797fKHT1u8ETfi7Rke/FN1mFOxLXHt9xBZ7e1Cj9gZxxAYncqdvG9O8pVX5OT9z3Zk
ATkhcbLYg0rdI5JFJPNE71nyyE13g++G2PPgiMhQ+bgWyPf9OFUglCHUIK5AyeUSpSivPcTnc3y2
5jDSHfvm5nuPg4hIrd1anTRhUaTE0Bm+r+EvewzgeSj+UXxOGuIiM6bjCo5BOxtO1YNdPwXCnBQn
6XIyoGRlFoOT8mI028cDHD7ANsSW/HkylpR90XHG89IOC1mrKTC/oHMxIhfxLr5Y4HV0EbplIflU
3nNuMJwmx+xMtgBglGd55lVnODjGcG/1FH73Dn4CkpMTifJS5x6YKJx5n6OW8I9E2mmY2neq+Xgz
NPhWlyGXeXrQsXU1ocPa7DD7oQoi7dSqj/enp5NZTC9esGjKQ4r93vWQ/13O0O4uk4y/FNskupVE
BuLN6esQ9PHGNj82XqCI71uhXAF/5ljw6MBPwWMSEdtIzWt6rOySpylqMybsIhfHC7MWkMuzaVtk
iMkJ7t5Z6dKEUA7exvhHr0+f+v/kyeYn/Osgsggp7A+aRkhyHxVP2+rrZ8Bd5UGIMaj9WTb0Feyq
TEiyp+pTifUx3MUdK7IIkySnFEWuNbjQBHX1LQSC0Tky7ExLMb7Qy3iHKnVvIqr8zfBuAW1rVSUn
5cDmzjGVnOMFzr3QkD5H9W9ItqdrB1gCr0bDLQUePpW7IrvU8GqyIgeRcjpqlJERVK9jkKLVH6Zp
ExN5FoagNHihxMepa1SurLNz/gdQfmQHcrPt6dPFZ2Ahx3WyNVHmi2o0rmwTBZXspjVMTw3TdGsV
vJ2xKACwMwJ0BtNJ2Z/jIdBQ2E7Gx62cj6L0iHwN3FAVQ7M86kwD2ZZ+6EwCDOlrjSb5HsQIdme0
rFomOIije8tFUn9vkBU7ssCirYAoXOfzDqB/ZQraRv2tJ8kLoJEEiJ0WziGHGqquPnxLVshINKpU
EZDEZS/BQcSxj/OZrzJDpsLokhhmgEWmhBDCbCthOmJwySQIZ3LqSu/sN1M3CCGSYD0BH3KYyu/Q
H0mjzCDKwq6ZG7ykgrfcJ0Mxs5Uw3mZ9rmjqtg5maJHzWiNXr7EQkynQqIMZsb+/svjwV1+WxTHT
ElXP4/DI9f94+EHwDhSOTcQjxdmeb3CeC66mYIxSJ2ps4eOBexQW0iHEA2M1NClhStaH5GDmTXI4
K+WgukVajf43Wj5Os0w1K0hdq9Uy88Jq3MzV2Jf9b2MCPh4OQqMhAsti2bHuN7mtmLoN7uUcK+yX
ybrwZpieR4P6uAASyD5iOrbaBFoE42eeefYZgO0rBuGAX7XQdFJVyuY5bmkRe+TpdZGGskYMX83R
ShKeqAouuiF2tloiD6RiSUilgEkHQFmpxqnsftaYsd1ZBN1Na+B6p8wMTj0/184RXQEus7qXbutS
89/BHYLohbl1BZUAOnnEPBvVO/WPJI7Tn0PPulR8EObhrK9Jt+jjExXoEb5cQOE9HhRF7EG0h4xi
ZvMhRkfjrLrBgcw+1I539RCMTVK+vyTtsoU4qo8ziGqvySIo7U4otMr5065O9v1pksfAbEGHAcaH
s4LZymfoagOirbxofBktLsutFxNyBiMTqrSjYm1H98n4xSRezER8vHBYPm5cjwKQk/CWvdA7toWV
dKdTyWE+4kNLfIqEsHz9gGQecDlyMrqcz78aGmMUoSdholqypwI29+FKX/Mxd+2hTKpeWJcSeP1f
jG+BOH6Z4vx9a7cgnCBJA2RIgHgJtsv2i/lTIbGTpFRkPV9Amq5PlXD3WJNqLDsgJMD31OV25NOg
IO40PjLim4vsml5IO1x2dqPDiQ2PiWntLJyRCbLHBxW8fIBwDDt8LUmwuK5gNdxPmMbaSNOKlxKz
8l6pC3Pco5YvKZgi8q0Kjay8/J6BBuZ/sy1+RYO3q1/M5fCY2GozW0PF2KHXZ9ywHGmpS4rO+iFh
IfSeVya1f33CaMXGnEsDpKRDgWOWruL4zpNqMIElms0qTckSiybzcHTZk6ssEecxkAUob1J7iP5e
GUixlm53WCiKKV1SsGvI0KdO00bjFd3RgfHYO9PVSCtCem+MaS28W5RmIXGDyB8OUlx2FAM/aUzp
t9BayUx9ouXReS4ngj+gBjJ8XgGEuNndqgd+5CoE9olCuQzvoKQhGI61QUd6rsazBVTSXN7e0I7I
SAsbyh1Jc2Ds1Wrz+Mfm4v4IbL7JbDOcf9lHCAttkp3C0rFmceO3HVFwogDcx3FdYdbyjvhEexWf
wFfcJbjLT7jUUG5PBAw1BxY1OPf5UQ0d4ODjX5w09hIacsvGbVo8r6sHYFg8pEwVz48mYQDyTZ2K
rKrcUD+JGvNWVAN+fMQ5RuXLcNd+JS7/T3Ptg8+pgIaSZa2AEx2qW7FvDj6UdM/bksuCGK2JCxEZ
DYCuAmdr0OS1kTKcl2VItixO0/QapBuECbgP1XT2Wd/+NGD4idAmjBusn3mVlbFx/TvXdrSmv8Jg
vz67KNivcyCQeZmLYsYZsdAAMv+INayKphVuunCI1yJ7gXg9WxAJzayvP8X9bMkAoaPcxgAqv7ou
M7CMk7ukV/GCmUtCOMhNa05XQtHmWn+fXCrsEbV0rxY5Cac6KY093JlaZUm0Avp+BAnlLxeEyy3Z
wwVF7X/vjPBG22nFOUuNRwa2np2LiIJe/Dj/K+HHoZyuwdTYNVHS5heuqmLnur9Ivjg4dEd2A07j
foS6qLxIAEHNkhCJT7JDpgZuLCixRekz0Ow/SQrMfFg6w0HySis4CKR5EEgA9JFcVzi376Yu6/7H
uBQphLfQMFVLJ6ZV9qL/1tYk3PMCi6rzsBynu2g+Q53gOmuuroUn375Jn7P5blMlwbEpbgMryycW
L8Z+zM+CeQYoSM5bx8W3hvX6/K7bUcC7xI47upzVu3FLjJGR1WhShQNQuHUslXOmGZODVoEoCJ8p
k3E+Rr0borxdRZIzM9DuOToSQzUynh5nV+HBmqF2rQJl9N6awYOxd7D7t+/t1EgHiEbiy5d+0eIm
L91/zwe5WXsp1G2mr7ET8YFIXrSQu8uK5kvnJnDJV8v1HoAf/l/sVVKkxLDlZvrD6PX/W9kX6yro
xy+DXFFLOHJYt3+6FFnKoXlUd/uCGJvA60mwi58pTfMd5DcVzDnd3acPx4B15vBDPIgvHtWmIZ9g
02rG1+iJwsNNnR5n8X/8XpdGDqPcucqZYCFU78vmDCu38af2jgJPAVkXfHFrXS8UwEotqCvnJsTr
dAyIO2zuwDI6lsqWfePEwkU3FZwp5E9oEmLB/WE7APzGTPR83pOWnNxZBi4npdCewG7IEBaoShFm
FAqtyan5tSatLdyU02UvK+BG4DittN/l9ViqftZVHFbRm4n/ueoE4Cg1+goAIfbwARouN70WT40n
deyKDlbLisAf6EoV2uNGKZXbuT665eoVXJdfhs7w4ok1Y4QHha4Kgi7YeObY1cium14ZFhq8awpA
GdUw18xOZUHOhWcbum/Ry4AQeceUh7UJueHaFh8sw2i6d2cXHCNH9i3SFb77CId5yI4bd5jE2Mol
5oB1xjrdDkTfhrZ1P7miY3gLohtETqX0Irvhxw55wtBoOpX2/BKHSs91mY3rKwO/Uw/aG660tELq
89/StJg0RiZGhJ+6q3O0iUJJgUJ8y5TSRupDKSDeZtUqJiIyWjEybaLOYHZAgyx457mpgX6CTr3F
0KvLd2LH2RBz2U50OgJHepIqKzmMEGS6X4Ps1I3vbugxUfgyoWnVh3Oe/HNY1BhSK5KzQAo4d/Va
pLLmlaTup7TPLw/QpPwN854JqY1Q4QA/Vl+hgVnZ5TNK6IElHCDF7EKQvHayXYbIodyht5n57VbG
Uhk45C/4+f4zP4k4eLNNlF3rVMCDWb7Zh3kkkzFOtAWazLlrxC5OiLYE4qS1XEXZ5LfRQvK9zG7l
NLOUIqVKvUDTwzKCsGOd7RuV3Vr5diI4eWJPCnG4yIeCeHNJ4fX6EvX69WAWCY8RucEs5IQMQUbJ
zIcfEEA8GzqozDBIHdWV+Cxe54tRRf9sFYXFIlBue3eygaIJ+CAWyvF6FT7IFbX6rBGNza+NeEhZ
3fp8gsQ2gh9SwbKN27yWaDOfFN1ckyWax6UhtjAj61ie9pSJyS06LrjJ2/KHNOyrRPYLARd2/Cha
YyoWxE0Z/pJ2d9eYNrRj4HkI8hX163h7I5H2M6VRjhFllnK4BE7kfw22xSOhM/paY/8JRYHSVFso
4P2oPcGRe+LyrZQY12r+QIarSaM8Hm8UCqkQ3EUtBBdnGyR4zZKDMK06guo0nCcVF5vMkPVbkzBn
QnK4p/Y5jJm3gz9avStM4M/PzjrOIWbmSbG8DFL/VQUl2fKfIOB1NcbhVIuYVjzMGQIQadZ7Gft3
3ygk8trDjLl0XdeRB8ZI3edyoT9C9QJCE7dVEUdafOiPo+JZkQn1bB5O9CTMyvlzO21vQborPcRB
1x5GIee3xXgix1BZMe3212oXqFrsmo4Q0WjTqP0x8isg+cXe0ljFmsRoxko3IYzDygynoB6XjGb2
RKfDrgOm0nCQMIwn9BPhGFlkZaT/4CkMdBxhrrhQ9OGFgOqrs31DHNfyrNHi5pFeXl0TMnSLcGjp
d1cUQpM/JQtdvMg4uxveciqeYf3WcWiyJhcD5fEhlCyUN1ZJL8vU/x7wNsR7frQ2/jtzLG0zPBXV
qqzUeMa6SSHuN27kJqKDFYb6qXr5bPJtaWwIaB9tGzPk1aGG04B3SpTDyjwQqtAomAfBSkG4f5oa
1RK3b79Jozsn8xXO/1+OxQr4C+79FjLOpG16/Df+SA+9SGLAlKnRA346CbxU4XrLhvz4lTA+wygG
+B5pumXhFgdw2h47xADl6ntt4X4Gjn+wO0wLuovNXuIL9erZiW5A4xBr48pFpp/GNu18uvDU1vEw
R3InJsAc6waGxkN0261Fo/ySsr195aF0byCz89eBw33yXP374GVptl5kjQYIhUamEV6YT/DXCzc4
CKZ2eXWNxliQBY2BQq/wPAHN0hm35N3HUAdt0dIXw1Nr5QPQdjDws+0ShJBxmVH2ITU23JC5DB2O
Ncs/ViDn4tvTgfznrxXN0TsOeUG923I/MA672QGhk68w1WAkQ8gC+7GA/s7s9SHSAb7Qb5Ss4j3F
XFgcuf3+WAutTH4t4y1AW/p6CzJSuwlBAbdPYi8/Uf/T+yrHuyvyT+fMsmpBpykLSNImfyR0C/Qk
I8UCT9U+J+il44nDasx7AXgBqozwBqDm05fe8eI1+cfo0Im+DROt/lWT+IinR40Aq3nIVyg/Msb5
A6oniiI5yaRLNILjwcI9rccVXN96M3aHGTVMSGhUtjg3T5jjaYa0ZJ/l3/IU2ggD6lTQTTxOoi/X
+dtWao8IYHfYMPjp0aSd9PBSpWPAPfzKvppWam1QfztdJEwD6JG7i6NXNda0QUG9t4aDz2ymGIMH
hOEgaH69F9+5mihUty7clCbW6iQcLgeD1rH4N4K/+x0YC8Afz37bWqKb5CXTy5YqJNcNlw1rkNGN
v8NwC0wqq/jQH3WpAqkpn23k+XjUCU5/xr+hAiwUam7Bi/TqbQD2YL8KbVHg88l5KXBGrSIC0RIb
EHqg0LjHGa7eoQsbj03FWujnKOexjdWp1MeWkDWNFoU+2fcSiJdjG0m/Sh6Jkkp5TubV+bGrlcYb
jw3GY3DW9/yLNCnHNDVZIxbTeS8NVlqaJ771sFyrdC1YgRBdFqFnxcyEJ1NrbsZlWXPvt14YBqCt
+UlMxqSR02eKYmmA6XFaEdV/bhoxhGTxFCpip6CAB2+CPJrxrHsXaNeFFfFQiYxEiCvQ8t1MKl7y
bENGex+P1AY+RBKdJUORu7ph07yFphwfR63inM1FJo8xOrhFoikb3ZhQwyNdqkMsxOZ/7DuU4iQ5
hX5I6pHFmCAExJRplxmXiGEozdV2yJqNBYingy3wQo2Dr4aOS/a4FTw/hnExK33qfzO9jVY6GRKP
sci526lwg5K4J1HMr+6wBhHho5W/O7vAoTvYqMrObgqJbKQSZq6Z0b5UBQxmsGpUf7ZaP+BEmP+o
oyriOoV+QfvlF1nDquqPzkERIyiQjk3TW4EsTDq3vY3N6pcwbIssvZcwHd2f45m/NS4VH81el/BI
qbV6Ii+S6kqrJ7INBYutfAMLHDCjBKI6EmtQkjwvFGhQXLglBdLi6jLD6oPffgRJt7ix46fjgPbQ
z4P2mUDsyOEm728cZHXFJ+mpxPRGfnJr2XD1OSLPLsMkKz/Qs+51twKwRQ9hO6I1RoVRA9dyMiPt
yvIHOVcIxT2roIQ+rTWYedwW/BkIFPYxyI9qSQUkMOxr8tzAYqIh/sk23lv5LVYJzXZshFwgwOhl
rKLrDNMEDYN695pWW4qOTR8QfmBMTrO3nKFIRu8CXSiS81+L8/kz67dn5226NaIDe8W+NA2rJZxy
keCegeVTi9viwvmMC9DKy2ZRiFAVRdTbCikcgZ7ujwEViFtfwk7MGKZJAViXb422y0yQXj1ZB62Y
BAKs/0nHmXDFt41p3Qi3GIjp/PPY1Ji2QQWtJjXCZbaV2M8NOFhO7wzXsViMTh0ixsjDeos1VvVl
3Y6HjL7Key/rv376FiDZGyFComFpvRLJSANsST/qvygpT4K/95S+5A3vpDOy22S5t4lHjhS/ZtWe
bnimcz/Y9v5a8e/gG3FLNiUPtmDYLFLgOYG/rqH4SsgWApZPACZX4x8mzg36DXMWdl5bAJWhdK+I
c0EKpLCyVmnQp7YDKO27N7RCtkJnKt241zQqc/roZ+hT0vye/ARNO0kxmBjVfg2zXHz4aw0kszxn
c3PV8j8ByGF7n+Kc7vTXidAh4GMz6PuqP1vGD+y/xrYS+0RE9LWVzb02In2syPfzPSqS3lJIrYcg
XDlzPoum+nYuMStgkTRaTEqZ53fGotdHtqZGpbXYZeF52dwj6hJC1M196G0r1Yb0GNEpi1dl9XqQ
ClxhXEkze5mH5p/LhVRXxNurZlUlwDK6mqlK1FjJCYBb30a4y2/ff46rtX7Ddmhf1DC9rNQAZGdE
yJ0M7amXK9rEohsXGX2Tk89AlEqdS+tzukX+c+onBBChMAX3PycyZKeAM15vyCWjvor7h19+ajeG
pmt0xv5uz/yFrqPstzq53DU+T4FICK/scRk01L9v2D3gsUF7G20kK1fYhspEafPFhXmIztT/MMXq
2Xhw3hFZEyKzO9XX1xDcR5h/XxlFN7G4/hJr+V9DJZuZQcl49szl/mdgQ3eAAEKT/eOZ8xJEF1NF
ob/OpE1uHDuHLCPGSUvGQEfROIZaIE8LyTinNYFjugC3z6QtWcz0GJO+A/Dgug9Wo79wSJwRMExS
AGLkPzoqdpCOenVLcJjQ3Cdzi3NTbxDIRfxF0q1RPvljM4sr7hQOLMFhg9wDWnNnw9GQDlJc2lsC
KWHP6r0cGt1ou6i5P02c74D5sr8rwNTKqxWa6NRZqAglr168TGfKP4A5osUHkkObItWT3s8MHV7M
gh9M1W/q5Wz4WHdhaJ+3Cf4fGH3QoDVVigi8I0SHCO0Z/u8f4iTKb7hvz92LNuHnjxDxguMdq/fQ
2Tviq4pk5HJfGiL09kTGrUAMERyexq6fGX+oDQEqG5UhXhworQVg1fNgJTgLo3BQA0sSue4TVfBb
qH0oZj97Lej4d8QYp26K4uB7lk1O1fYmWUbRYy7aCx5BbK6QfHkbKTo89Q18pj5CRR1DhCjJaeOZ
yOiCKtKYZDMh5FD1LRu/+tOs6D6e8FZkKRwYhcLIysAr/v3tb6Wcblpcpnd7o8waFpiuRDqDL/r6
+fMjiBKY2S7LN2GHoXcKoeb/BGM6b4VvMfbwfHZMWz7En8tnDGycQ22uan9GF9fa4o3zOsclTuQ8
zbHujTpmKhfYS14+x3OGZL5qVerGc+3O41Mv1XTOLRu/0Laid/DCsJNuH/Pn/zBLOmnpyvZqSmcu
J9T9iDyyg70UNlrvwzuIS2FN8NTpuOfdVNhAMXCXSBa3R/4zQTXUwpnbOT7irlbppAEaezN22oim
8ilS4K7JdBbF8lD1s2OrGlOirXodYbsmnXpbxTeJJuSn4lHeeXX8FntXx9TSRP3HC0BHsruhwRIV
UqjNC+CmZSlirUS4oaFnz0ooYlmBp7l885yr2jsZXfncMxf4HBK7lCnK+LyCM9UXqeHv61pl86lr
BlfhrUuovpzdzAs7jHVEkb3AXWfxdJ86YorfOedJ2iPnAAhRz2hEE1qeo9zCaslHcT9mIJN3KrlG
RGbCpiSBPxaJz7U7PIb34y5dgr3xVeNkqJbfHgaeOwSk8q/p5v/Q5kUkPf9RFTWy+UhD/z3QLMnZ
bvFf/zE7Hue5zMPeQq83Gvf4m+7j2y8VTqrVV0qyN1wivVmEYEPzsV2bWazZFUPQCkQ9Oag1uUGq
sX+F0h/u2Q+PqAkVuiqGnucWyzMMLVG6yCMJra3MIc4zLbPzPeI6Co0KimkK050hsPwuy7PytvQD
WcjiZj9VWqKmCNJXaYAhVlmKdAWmIyHxgzip3kD2XG1cOCS5rpPFOl7lZ4Un1q1s7MG48rujqV+k
70rO4Iq4n1/w5x9syfXUNkFwp2B+O/JsQksdprwTLXoSBAQFneMldyeXhBv1whKbCGLnEOXRmEvu
vA/jye6LxsgUTCjLIhAIq4pbsNRFIz+N9O3UZJXsuZl/Rm4Za9I/4EovXW1Y4XkHJMskVncDGHqw
k5nIOtbRWUAu6zmtkP0TCMXnvmfwleKQ/o7ZhsoyPhkyScHZTgisgz5YbV3ewUb+wmg96BFx3qHv
tRGUN/cc0jxvnUP0VGQ97xc1BK7s+aQ1LgggzpdjbGpJZkkwv9mijeBPiGaHBlOY
`pragma protect end_protected
