// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
tvPFZ4ymtUKESqMNhSlqJPAmAb6Tp0gOHMRdHzTbAzRfq6lZrlAJ/kE8+H71JU1r
e4I2B1o9fuboJMqDE53/VyABlGyM0usdKw7hxPeex9VzWbw/jtv+xyV5BJhl6D2j
vhvBO0iX7Z3hVMflh2ZACguNg9Ab3S5ZwNAFLR84F9g=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7376 )
`pragma protect data_block
9bjWRNvevafKhE+GzmlvMinRR2qWs47bammXzCVRc/zPuxSUZS/Vg9+aC7hAXS7f
3vDCqZ/KxWa2UE74cb8Fr80fo/Ie/TbQt3EpNzzIBe+77odyGzCDpD+qAf6R876b
kP+ZQ2vVGeH/0RMt3tpsFvxD6q3KOJ1dsx58OB12FIuew1nmrSKwJIAlkpUZ/yA9
a4R2bi+lrpBOc4RKUp41Pq60Wk4PLX3ZY38feErvggNtGlpOZvEpDD3fWvjLBhi0
/vTQFyLHHMnZePKJlqqzWUzsrAVbA8qF0hzsYRwHdIKRMI+TiCMJ+hlbPsbDBOcs
VToqf76CKvWkk/f3eMg4fXKkmaFSu8WVTjI4Ri3dhNwhrd4V9QPwUkMT+suGM91u
Ok8shClMHiN7DAzWPambZ81j6lyTBRSrH/Z/P/GDIAKfm41NIZuESe8UYYfwEmhY
3XddPXFGlZQMgkOhIBaj8qmcMynPgQv6NFn1SrQLknz6S9fnJq2eACam7lUTzgEh
Z81pX+4Jjk/ha560/3bxPjwCNyqpcH770/ip7pTriXOjJ1yzRaQbEEv4C07uF6Lx
x84wcoFkshEhvDoxKXqDUwubRbxFoCWBHHnp2LOOauSQGM2txMVMbgU21YUbWQwz
UCwvdooohpEbIhPekFzRD/QHw6wBpCCEDmkjq+EUvJuSCgV5cemFKtozxCHHmKR6
jXrHleUvab7sYdPqjRDolQ6REfdGT27DYIDJT08xR6V5TOwKjSJssdq7Qc5FAPNA
7a0Mb6fMYwHOvtwYfgzlEKg4+UDJPB7MqzWrqpzDz4GSmawdHtWGzjGoRsTXT5lS
tn2XgB1o8DDDvDUd8l3b3PM40jXbcuHfORxMIBNkcO83TLsHmBNEgUmz7oTj3ast
JNrUwpy5CUN6dlgVkJF8NoP6S/2ZFJesrxWeP5HBHP9yvpoPElOC0JxEz6/UPUjJ
6AmmljYN8h7K+sqcbaGDBMRlAzZqgHwaPiASmH2HQwVh7Tknk+CgFNhprvwf6uyn
bSFzwoOGiULJKBGncdSrq7RA8dLUnz8azGjzNQ/zYfdT7B23tiWT8BfcCoKMsX4Q
MhTD7NJfqj+2hFy6d/t62W/0L1NupJVBRfs+JJnCz5Ds1vEdvYkRKNsnQh6EB5qI
cTsi5FDuLLhpD4m/mVh1DybvDyXJ9wvMvxL3bNtV/1FhaUqJgI46sNw/YBcucoE3
ywOWeZcra1rdnYgoicWsnKN5AQCq63aNaxqDzffv994Aar/7eJD7Q6IdnCmySFRX
Dz1xYHlkBHgKpoBoqeozwYv5m+UxpNEeZdykVXaWb3Y+grd/qScdr/Mi6+uIww7+
WiUkBxqbOaCFPr+pKlN+UpkbuLQ8TQy4cov3IkCpgrXg7hoBIp6HUeWOqR5RpEBB
y2ZHSAhAIBdNBoc6D/cj96ZEUB4021ufaaDa1q1WzC/U0IEy8BIrCaGIPskXWkU7
xgdAWLT7l5F8HW+BNZa7VtX5ySjMkwEqVJZzOo3Ns8Bs3nyCTkOKr3AuRBxM4w0l
EOLJCr3+hCRbdqOsvVitMoqQu1FdCcjFqNu7gjVW0XwLdxv6cSlXMOV5vsGdsUS6
6y/ncgAbhChaxMT8qlSVzfEOSwtMr4E+nVa2UkFRiQvtxlyUKkUOPT/H54dIAGn0
r2y5LoE8lLaxeKKCTUCXFeLYfmlRKBljxU4Dm00EmPMJWFAf5l47giDhCJ9haVEy
7h2HB37G1dedxsgQVt+ud4wV5d36PcSOWuyTfNfF+0FQ44sEPn02B9BgI7LsqtaQ
hiUDqSTdYpy14LPZLSt2S5re9sAlcsqWsA5sMw3xODJicl5GOYtkJsGPrCx5m1vh
q9qbOxtB8tKiR5DBGDFfmlMGLR/Q14WM++Mf2mOumXfE2rTzRcM9wschPeE1RbZR
FfYEkjFfTgW+teAXb7bZJAtKw5VaNopvmn0f18GFA1N1OO8h1Pl3AD0PCQS21cRv
TvFnxFSiBNRDbpHinEMUVO+QrgnQMu91WVGBanGYV3HTw964UUaV72qdj/Ke9cGo
N8K8AJp3fMgypX+1s0gsKhuXl54JuXBZv2A16k4SAowYKtYnF8OrRlBi/Pxghy1C
fhexujOpCm9SYDGwbfhzKpyhN710Ds7EWXgyCC8iv5gAZOV3FM1FBApE+5Fq/xhh
42KNNiZQjy8A7zKccRONcqyQi0+fiqntadBO2sgzx76f1OzfCBXD82y8//L4fJlG
cCQEsAc/YL9xds/twCzx9c/TVvrxv6olUOCBMu6JChVRLDgCNnaW4c1v26ukvCPC
q3T5qvuNJiG/3T5G0ZMqRBQyg5C93/CJcE9iEmQVW+AgXdbLksHSyVnlzzySP06V
ZARJrn1TU5VMHVliMfg/buF6/GHNpCB6mxOCQWgJqfnQklCglZ9XQOuw1Q3dCUYe
OoUd+HFu4e3Q6wdR6K/2JvCpKKb/4BQcvMn1GTlGwV3JGy82ieJVlLz4OOyZfO/2
J6AdtHwS3CDZMnWNjnaNVWPIcjYWCYYRU+FFtTZVWyaYUB/zA4DsBY27tDrzf6A3
2fttFZUXiMlnjSwUpYn0fr1KZFBQ8XWJKXE+rQjCNexz8G3XXGz1AdyIxqtafpoe
fztROWj65FrLqtPYZt1ztOscETAMMSwQ1My+1z1Pd6tZ89m65leWUsClW5xBllho
0n4NHtKGk2tKr7OEb7MgHHs80U50dB1Gsw4EMlZWEB/Vx4bfpK55gAmSFO/ENBGi
fcbyRCrHd89PQaIau5SVv0vH/enexlJZ8p5iaseX9ukF/HwRU6Y+rLT2K/NnBKOe
a5X9AEsArFVHqhwdqDa3V8HVrUuh+crnP4NuFqfURbFLb+Aapi4C0nu3yJKSq5po
s+gRPYFAAF1ABGFIgo6nTwzn+u/MTt0deGXqi1dmW+Cl+RhfXS3AssHxhCOzP52U
xbjOocVaxYcwVdoxxrakKFbsKI7oiJJhVK+B3Zk8mQFDXgluARb4PAad+GSqj2sk
4QI7JNPFLD/7W4gzk7kIHk0hXfgAny0lyOFqmbQclxpC+CbP1QVX5twLiUa8ivZR
nunkzAPjlyPm7wZd1cXv6pUPZc/J5ENmBTESfF0MwvpMxpDg3PfJ+reRTN97eFxW
TnCkTVszplXfb4nkS/1eH0YQDathqxvLxxg6MnQtdo3c5tOzK80sFDll3KC/+CvR
seFIjKnueAeZnBU9EZW/zAN6Hhi+oXeTuBeQho2no8d2qVJ3kGv/V5fT14t9/gvs
VEe5dXGo5FXuq/5Vu8uGbv+R1QykgQRFUYZ1UOQoMyc/6DRmfGfLxNOfSyI+2P2U
YAPIIgmtVxsBM0LuGiVfBukA9Y0y+MdGpmjhktT7kI3OPUwWrW/w5c05+jKNxn1R
aQVreZLQTRvP4u5cbQsgVHGAwYisjz4diqMg+ZNLHunU+kdWuMEqS3BVSLH3MP3W
2ps/y44y7tDh+EMPizjlWS8oVtprtCzN6NfSe0PZWK/EaMEKV0GL4DOiykMr19T5
1p86NWAYoqXWJp4ifdKHwIUHfKtjQbBW5zVBHzub7W0YRAdv103F6TioeU3R6rqy
sKWyotGVVGSHaZj+Hl01MewvH+71CJqfdzAXmtRxVUSBSxVCHD9ZWjV5Twkqrue9
4yyetAAClEGka8owx3/V8ZcDvcsfSdI0m6orury5xu4x52dtkvNh2/9/njay9hj9
zKW+6XBAbFdj6gbqC/Rczf8JUKBXTmI7Ha33UDWsQ8X4STwqlbprx0jSAcW2d91W
LOcdBDImoTNZYw5bkUq4o4hKvfLwnhEl05oqOX26IVTKaLVyh65hnai+qIyDWH1d
Gu6Ir3A6pwQ+hAywdW6TT981koBnHOKGrjQHUSpl15AgdocP6YkJZqst47Hbqr/r
LnNoZKmvfOhmhENoyl4/9oeShQ+IP6VibzhxBjutqpizGQUcJw+EP/TtJzamg4IF
2mwek5qbbt21CIPfaGOTpyzwitpFOV/qko3KCKoAEzIx3fyDZB4nw3gFNWaiWdk9
fmF+J/c+/yAPZiHeTjVkN4sqwLkZ4Smn3satDw5kdbwV2S/Y9hVpgfhdM3Msln/K
YAEuHmhmVEO8IXWKh0TgW/56ux8Php1Lz2IbxJVvIvSMcpXFYXWXpe3HHjdeIS/H
dqqTRv8BHxBXwkg2gzQ46mbR+oseCvy18ST3fM3DFbbFUi6cM1cEytD7bcCtMAQS
izObHZgleSL1yVaaGs39AFNFKYbwXuTZoZ2y/UzUI+f90wXUJBbG+lRqbrj1yRmX
8C1lg9CK5qkqgohWYgKjOJgSDS435J114P1kgBDarL2QLFmaSEU7A+rv5dau+eVB
qjR8YOIj7CaLuZJfv5jMNlRCiw9rfGBnnXdMXBWgj6tjIxRY450tQJ9hsfPna9C1
6p39j6X3m/EhHEjaDi5NHhqtjPrvlWxNLRYB4q1Iq2y8baRhaJayW5LtHmbTpZZN
b4smr7eceCPA19qFj0++GEQe5WO99vtkxKnO6eHbqT8+QEdnZCkjcUMQyLeF2B0o
YabvPcC39pa2Z/nNK+wGpjYfz2EQABRezaLREBBSNOqx3I7DNNTlKM8+Ew1uP33e
j/EGTtlSGbYa8UPQr6j5e41D88SaBrCHaTlG9Oool/665hHInjHbVyQs9ldcQdDN
A9RoSEyepeK2F3iMfvxNE8q8qG7KpFA/dcdUtvOmo4NcM/EevnyiBO3zPU6eMSkv
PiCJxauGgxEjMCaO4ZKhhFMEAzoG1N8ecJ9EUssuZzRyCf/ViQVI1PbKAx7BpIEI
7lA+lxiTYuQCcr7aK0cmannJx/i+TqSqkFGiKpIiNxTglbV2y1PwJEFKlGm19J4j
IoK4XAfKa71MT8t2W17EOv8tReysapGkCX5Efxlk7qJn9D8Eg+PD4z7sX5eCwA3B
z69LtJsK1olaAv2SK72oL7KEWE70X/F1f+/JNR3RhvZApRMCKs6WFEq2jLfTT92Y
vcZtgFKjtlsc+81Mc1wwpXZW/9OPUI2Epwsz9EXKMQBloWL1GnxDjolzFN71wxsy
HFzmWWFe2l4wXTeo/zoN9cXgd+oDBuzpPSy+jEZr42e9q73eJY/qi7N5HSwxpDKe
osOp63cqLUQvzZiWjExsRI4BI8HXIlEMTBjckEwG8BoNDx9V44T//fIZI++sbxJW
X6t83SVCVbtsj5B6U43qQoCocpY6LGgve8/T+INTIy5b8mRSxzbC/3stW1V6/aCX
xLk2AaHokgN97+4ZTitEIZFnwCOdjFaEkE+cfvEjPRzxY6wYW839QpKl4Gfhvh4t
awM9weFawKbuWVA2H6mBn/8XdRD/nvKnZzenWorMK/A+tOX00xnUAa8IkHvXJU5P
t1QmpEllsdyx0aWs4zfU7GKlaUxWp1FLmikkCWwbjdQzr5nVl4Iua0P5CcYDXZzf
Xt7EAEUfcqGeek9LFExq0Qx9wWr/4FZ0NMXtrYOvamhcPQomDBiGzkiy7ljA8QBH
T37TN/Gwwp2ut2XHmbXJXXE8sy8bGt5F3h4cJypeXr97tCtUBNhdQD9Xy4xZzXbi
+bd6MQ7h+bMa+E63h3c8CmkUVI6lB+XoR9OkNqVr6ZhBJEcShz84r+C4Zgpieg/k
qajuOfOiRqr8cT2bWFaw3YBzJ+hFSzt+pUkL+P3Bx2wV48WnfY4pjuNonW2fv5QT
yw52JxNeV13/hh8R61NvzDQO6EAMVIy7ruX9Bn9TFjughTU+oDMPpOvC8xDRN/G7
8G8aZmLctfJjm/zID5Y/dLMGVUjcdNeiFdQESmFErdD1npwdAR8PphuazEvCjFko
y3yMrVv52UdSyAKEywkf0tSOoarrtGrjPSH2Erp6q6i12DPvWoSAjrQweCMILidM
4dIY4j66uK48dEjeKIdojoI8nDhuOOaBwkEw9sXk6WRS1OuPSlLQjBJt2eWA3FM5
Y394BgMZntnJCSeYuOI6WQuDH6enWD0zjFLAn/fR2bJMIRsE3VrXGxK4Z9/2U8ar
enjBEvcMGGYzOwO0hLLOFZ2F09HIa6pFaqkFVks2z2t2opuV6AZtCE/fzlorI4nR
K0ev6jMt8rfQPqdmGe36C8Oe1lfSwZhlUu4pYXGHhjiwGpPY2Bg6sWqVUnQVyU9p
fIDNkTTfe8a0DmVC+07sVcW6gP9G1fNEy9ZREfQVcmtT3N5nOTCG1MzXseoxjlsX
ECmsOv5nq2AoIfVN2nUrPg7xrAfZ2sc3KMLTPQgpYDd0qaUzsFlFhLbEEYecgna3
Y7ytU9XTekEPMRP7lfGscZIFr7JLdOr3UW10vYxtkBMQ3PV2T5nEJNO0EQX/RjaO
agKPz0KF74eK/UsBbHipayHDhxw6AUhXBi/IGED6eEso5zmCr+6FtOWKiwhnlLpu
80NydF7UFliG6ygNcVX42/Hf2KDq2FkEDCo2vDPbK2Ijp0vBf30TyG1p/OxUQ0QR
m/CTDRE4WoKpH4p+cqF712MPGM9W9VUQ7uOAYH9+43kGgQbcM6+M5h6RlwUXB+XN
Bz1UHooYxHKTuKo7SMpzBB+lywsJtP0J/ZyBfek08lBXd7hYfZcmzYtsdrlwE3Zr
L7M1Gvsl3UIroqhiWHMZJ2bwqtZW0Oi5sx5xiwIri4UBVb4ZkDX18/F2GxD7lwsU
zeJvqJa528ukxJQMyVVttBtSRqAsyjDdykHLa5aU0I0kDVPujnIX2/O78UwxQmvP
gSGr67jfQ4sr7ugGLZp5gHlMGmiP64Fyp9UxP5Z3jRDnfHFFRCIfeyHyMT2F130l
w4PW8HJiRCG+rk8B5m/7q0PSe2y5LrD0oWtK5mdsLgu4imKmxRrr7HT+I3pb5T9c
cy1HN/AZJ8+jmf3jul1EmnYfKzWDSa+KxwC4v6tPynT0Y6cA7Z1MOjRcF2Vxc3cK
eLM3sS7s7M2hNpOCfc2bRGVyOu4DereYEkEB3T4+SYWWGLewUZmHoWt3eS3Z4Fwt
YujcgzdoQjvrpZEKfXnpdRYMGoIr09WTRUODnUxTmXze/NKFmB0ZmHY0RV3JGf5A
Gokzdr6jFOLca/5q6DBOA7UmOzRRUzdpleNtwTrUMCOsz5beZ6X/1qlXP19n7WJn
haWkrckBIVTXs183EfN6JAOLXdhqK0XgZ+xSj4B/bHOhH39lNB7qbffQGGLYliae
V4pQYKZ9JPbCE2YsCbuJm7nPcIrxNWmb70kVyKQujWQiveEWye/EcurXcQ1geQSq
jlHlYVBW+AHNEkcPhkk2tSBLxW0AOQUqCHKmNyKmtADKeilI05FOdTo9cNWQ/rV5
faX/eIZ3lca4ak6c0KUem1YdzGrqeUnPSzvVNH6o9+HaRW75KSQQ9192F0gxiVZ4
OfS8RXSDoJAl/o+ewqhx+o/45CAtd2ybNFkpLG4vCw2KQKdROz9Gi0nFolK3U1Gt
3QTkPbA+6/gTLFcauFw4u+EeosJfYmRTYYBGGz3xL4A8CEC+uJDGEJLJlVMLAMwP
1R+TkbMqt29JslrcOdOIC8pgbaAxkX33j8U6sQl3R3Xz94NTca2zTl1jfqxAO1hd
tkVB0ZCsPrOrSB2g+iD9yQm9np+Dy17cqABS9BMRC8NZDVubXoTGq20UI5cTbV/z
Jajqoxd+0LuEwaH6/AkXOlnax0SStyxLC92tyISAUSqnOaQF7vcC1T8V09UWUBv9
2Pyo6WjTbE/iFylJp6Sj5u4jKZ43H6V3PzXy4Ow9PUZq7W7T243SwZ94vWBQ8G3t
gnUWJfEwXNuED6K5PLffQKjuarR50rzJeoLWhl0T+ENxeB+OXBNtnFXI06VVoJ0G
KKftc+RtzaTrSPCFDqk5ZG93T1Y5Ch3U8oTRUDU/1K839MagUVRta9gCAff2HykN
7CKFpiHY463mOXygiZw+Lk6JszEhhXP3+zvn4dQthK86W/KBttdRbO4sNBn/RCYw
LPc5WHP87B1uxmuPY1vA9gu6ABSUNCChEFiQueFJdM/ScatKbc3Mptp6bL9+lvfj
97OGmQTh9SwvfalHgHGnZj7IWZW36qsyQmyg+5PflaVEmzT2Z8ffahQOFjFg0Oyk
QzWaFNbPvHxRsXCdeqJAo3zSHUr/EcTSza4oxy+DCrOVF76m2bdS+hPy/vNgBxFm
gL3S2WHF61PKfTpf2ok2DANdFM1I3UDdTe033yCFSGT1MvpkqdxSt027sTd4jNGO
+QHc9+7aQ6b8wS2wdwSMG89a0jEj0JiuftQHmvyH71/WQ8mW0snViMN/Byxrexax
Gk57MpTmU+P0mVyANWK2XdXLI4PLXVELvVdGXX4NmEqYZAp8HHCZrxlMO/SvCZPW
XiDcJFOXkqBKHB9BpPf7LmygTlMvh8GRZraPnGs3tk9/bFG8BDuOkG27mK6o26QL
oNNZp+G+Cp/xnuRI87DHXuC5a20dVUYVT0xqoYnn+KRdkyHiPqO2hgb+mjTvCv0B
2w+/2dJuPMtiSJnxL9OyybHk7pO6D72vkkyr+nizoDUZJJTAsoBm4MXOoOp4EZln
+IT6y0gwGcsA/fyJt3NhKXSDnB2t91bUJgoQ1/anl7caxJ0cNDXKjsMGHB+LgPTY
hXRKBiwEJFu0vUURD6fGZgss4m4jEtT301zFrsaKqJw4exilCnaGzgwqsSgOR7Xf
CyRR5gZxJBTIJFfvzQ+qRr5rHYy6GnoTPn58i17IsIifq2GNi/cmFraz0E++azeN
Gftaecav7FLwZLL8kVIRUBqyox0nCbDGF9AKtIoiWNx4g/jEXTFwFWBpqZJMpDaY
CyHeuceakZOxPbrljJaX2lYu06gdZaoSHXs1tju5jZPGy2UynsAy64sdQ+TwDDSh
Wgd2rEp7cVbNlsztApxvslpqU/tyd2D9dUGKWCif87E7gI69ImqGikCv1iteMjLz
TEEZ02WUIhi3gxA8XMI1eKQ8lV+IFoSdfXXJ3ykfVqj5vlsgAlsJjgIBhf00pvmA
oLDzZqwaXQAardePVVFjTvheDQfsd3sV9H8YqTRzzjWavfDj2nCNKo/zo7/el7vU
l6rrxJL5UcDA/0KB1GZOOnkt966d6Vg8PnneHfJf1chWQ8B5IUEcMawNwr++lt/W
5ZOvHoFYe2I6uwqmzKYvAbonZTSY23ozeyDBX5dIQMX46a3eRtTMfTWkRJBFGdV2
qAOXJKyt7HbY6SCnZjcDNil35mrSW6AC4H3wxeFGmY0uMyl7xiITC6jQCkNN0JF2
nyHtRSkwo6AQjCJBeRcfMZ3QrVe8VS6icZQTbJVimb1NIxLJ8BA0beddcV0CsPKk
WXYAu8Tl6UIrT222TqahKg64/gOm9sGMr5mc05jfkcWBGHboiQ4poAW3BmoM1T7r
8Tkr2N6AHsqNSwslwq5v3MCkfCodZ5YMp8QUemZ6yRKXJfqmmh6XFWht7D4GKYy2
xhkDsRQT04p5HMwJ/xBlpkDouQ8x1N7YbVAd67fPNmUUyv33q2LLmpN3zU6MFxnV
IdQcO0WjoFEpLudNdpMQn5679M8RLyH8nXHv8wJor7C42Nf4bsJsQqlhMoJBn6Vz
ZdoF/CXffQ77STjxyD+ZiEz46InwYVplBUTscakTru8JzPXI3b0LVcTI8SA7m2Ch
Q+a7qSDtfD8D4uvzRI8csFVOBHoIvktZ2UFfAiaBvgPoJ6gsxhtXDE9k2YnBYvV0
O+T7+zKTxvtQpGTGmypfESnDF/71dKBntbzvZeZqdfxnorRScGc8xlbVUK9rHh/R
VcMhoFixAKFRRvVU3SZJzIktqMD8Gl7NEaTBEJmH6uRPng5Db7mM8NRk3dmBQPx3
qhXU8QKAzWD1EiPzd/GjfpoaRftyTu15I04GAkj5Ejg=

`pragma protect end_protected
