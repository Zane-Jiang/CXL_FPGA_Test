// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oCqfaylKqpVNJokGdU3AS1O0vqSR1t+g7T6u1m8lA6b4jQPVOmCvECxXNRWF
VzCrcYDaEd6m49TgTOxWRiHDnrQsDzFOd+8l+r1avSGu8Rl+l8xPtsXAdojY
w52X1eRgesDm+2ZGuhcRgueQrkH5pT+fhD2j7zqayXqptkCK+zpoIAHHoC51
4o8RbteMCM7FQp8fTu1HoYoUyLao2ZadmRKykI1cHeu7y9HEJsV6Mc2NpJ0J
gvfOTXR6yOrXREYX6CoGWnCYt3+L9jtVsjlHlbeAoe5rghv3NkhOtxmk+C6y
kwK7YQqupOf1eijSaX2EvPdGMotHiIQyWmo8zBgUMg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aAPxMBtuoWYL4iJgRyaDeopYK9ZtHZS1da7rMyrHNkVfJ5DTLs+VupJ/Q3+Z
rAL4ZDaNhgQgp56RrZ1GtdxCVUMWu7xVgi8Mz2Vrh0beUPYkzQLqQJXYWPUa
BHW+BeuZ/cUZ95xq69RuKFO8m6qJ3O2w6QphzugBrklb1jM+ICskYn0JeAzK
c6be7Lom8hNeAjoIthyyIHRNTGPjYavNlz0HWrhsrIVQAjgdIYTWAj3vkk6v
69Gc1M1orrmHByh9+dqfOLrczmfvgyKD35V79wCBfA021ukZnYIVT7TDLZMo
TccuajEec4D3TUHKnEQ2Mlz9kcaSD3w/BL/E7UXt6A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fitw67ObKBF3CDdftW+o/HMen24rg3yrg+Zi2wxM2rtkNq8mScCRN+aLD4tF
Srl0s6TMiLqdKZ4jYhBvdPaU63b45cLKbDOnYBWCI2or6zdZOGP1Z+j7fGRH
He/rpmMcMJo4puk8nwB0DkOFoEOHAtPP3s92feIeWnomIgkEGhr5a/KpbsJM
7O18TQZdNsQNs0DaBC7dYXfhOxOEb5B1iINGGPt5K/ZxEq9xcJXFR/BXnL/a
JuvuY0Z6BbekhOXylDyd+OQ25bAo72GgmjCT7XlfY5Rn7aKSwT/k02U3lapW
ToTD44x4a8q4bWsGKYa5UJwF/jexSdBBwxA2qjwOCg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XMLvqK3D6hj04QKaUpEOuVUESGgK6XW5kC8dDZCdg3EgisUZGU7r+DE/StZ1
Rv950irlARdA6lY+EREuF5oEV9r6ZV4PTPnqvz6YNFS4qVws6C66W1Av5F+W
cNvWRbfb4YvjsnjPAW7JqvJGklD2sJ8g/EVccqUO9Yqn7asr9/4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sdLOswpI2AgCqcCIHaNTkKZAO1pf969XSlBQcQd9ZtBRQnQv78QeU3q/ug3Z
AS3OzJQtsOMon2HexuQwXb9V2l5vH1vODlIU48ll8QV28gSMN9GToBoBWJq0
WQ0y7ga+3KbjwBoThPE/rpA2T9hQUFlMGjNZq5kDag8gzrbZ8yjspEjklRoa
coAYkuvD1JsJOpHK91/FAzYKpZR1mjWd9agjTwYndWc2q8o81JP9CQqzwcTW
wt9pIWvr7C3G2HNPYtM0xGqO19mp0It68oZv477/C30P6wSAvGuowGcws8Ks
92s/GDn9rLZn/fUTLDFAkjs6RfLgS849zV+h4BCJY89UJ0kmPI24LJditR7m
ojBlkpq6QYF9WYpJChFt+DYSXi2pxPHLC0qMdVwq4V6BS8KXKFDC49iKzS/C
d/p7i/eIBj+1zcbTzKqpvPUrFUjcNqg/fsC63LxbbncZfcF8ND7LWXBSrZTE
e1FhFUQOV3wmY5Ad8uZNsuXTDeKh31L0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O+BBQ5E2x3RytWgMM6KoK5w8C3MZ5X11dxgww8ElDzlNCUErPSW5OC4O19yb
t/fbvxOcpns4CLihkldWuqMSbfvZs6UF3/m/xry2Ta+UE/hVcH1BwgKzs/oz
9mqgJTKUj7lNWKSjTumeuIGwnejpq16vwdlSrrj/Saq1XC6VP9g=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
udOrB95FoR4Vqiadfjn9sMGV7CpRRlPX9UrDhRCaJvvIHqHIXDJzr6vzRNMq
0TgTr/S9Ts3GOy5n9stpjM7X4ahi3jEkkOa4Jg1LAIdnQodEb3SJ7glIVFOC
ASr5GPk66KsR4dWZKkPXkquP4ai7/oNYPKZcAd9VsB2UISjncV0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 36656)
`pragma protect data_block
togHTfqJR2hABT2t2me40239KYmjejWOA7St9dDjS+qMJr3qtY+HcBYgmAN4
w0lHFLHDV0XHdIJbxI32jiU3dx/2ZPpT2AiJO+L2brzxxh9/Cu+sT3Rrk3Dh
t/aeFGX/PA8dekC6PzDGNSSNmK6xxs2dWeN2ztBxwDuiNOY9LoDLN00nOZZs
teYbxh5tVhi/Ku8QB+RKVBWbullrUf4VgwnYzz/B65jN2X3upXLLjxzefNgN
5CjpRYmoSnFLfwaLwA5PPvAkFrgZu/m5mmB9OJHClsf1b49hXH1MzsraOR9P
C0gKw0nFvR1+gKRAwbi8oJYninnWUqfa9kJtKbMnsS56KEi7/wa6e4dbStax
piuQG7qiHjI6hnicxYEPODzVRfs/0h3ymJDdJq4b2b4sOmkpIOSixN7N4gGv
j2t9NocdfgO0qkU1DyPETdycF3sbfSS6+lm2Yqxc40lcwnIW9/Jg7oc9hFuP
ZDYxOk944bVjq7r0A94UnFfk683AkzCA8JaQ8lfQDmqCMFctDWc0DJ+pzcAa
5m4mnyzxVyiKKopLGHzknJjTrRAsGwlhqXRHvZL8tsmM4gwHwH6FHlOkAqu7
JqYte2EI7RhXW7M33sxkC6o/5Nu7trbhGJTi9+gE00CB/HMi7uVAlu5j9EjY
xGnwcmkxQeT2dSIW1x3tZcH3n2F4+rfph00PeGiZiTUnKzFCuP4wFgH33+q/
3Nq7JWgiz5I/N4yaZyWigKL0/glA3sOjQQCiVFNNqBFSe+mF7FrxoZn1BPnV
geO9kKvIyHRIz5lEy1gjDv54s9YOn8i7nkZQWfOfVLpkZIVucMykKf9mI3Y8
Fed4v17Vi+ADFmCPAwgygKJGVQDHzwgvcD3rnHG0bN5wLiAqlhjZJ97MN8Q2
aIu4pSTGDM8d5MqvmlAlNVXijfxjLJEQwYD1Y6v3IHxn9HtcR+43Uf9tiOlu
q6uxvK9j7miq+XcOKSr7HsBOCISN0cHU/0QoHoWOm6OgVUulmBUmWCIkRGDY
BrQ8h3xcHYRsEjzpguRFuJa5zN42G2ILCBX5p7KG+Zfuj3xCqNSwBs6IdeSw
tNgeDAnbGZsy+QYwTQ3DigW6hKIKBFmMgWQICXsGGnSUD1+XM1T3W5nt1568
nXHhGonD1s3rnS9cHJWVqdVW10Q/srtPvx0j3U3gKYvOAQOvrJwl81NT4umc
4uLTIJpYnYcXYXVmEvtz/F6dLcfxYGTBTJcfMsj3I+txotSzyS49RYSIuryy
n+UPTrMJJOMXw5dkc4j9DXuHu64L12j9Eo8RGrehB9+c7YDDwIRsDdY5c/LZ
FkygsxnkMnaH//thkopMhTZloYjW91AdyEsR3NSmak2viPlHKQqjMtknREU5
ujVpFeoD+y7X50EnoHpzXJEuFNFNwgY9FmUz4O/vCJ+kTyRuEN1g9gZ2e34/
OdmyWTO77VlmHJxc/X6iMTPi/zEE77aJUhvG+0yKd/BLq+V/6KHaosFuKczF
NZPA330yGbAqqwnqIxhh4MDQ3gehTAJQkkj5ULpKL5PgiUJ6KlKE89F2a3iP
jztfFVzKkn4zgu9ghQSh8Gc6Y0FH3VAhYqEGSb7HTRVlp/0h3pgy78D5NBKC
1gi5kE1BbYzqtfqVZXb86mMQ2VgBZznni1zzZ9IsgsIWtUcibbvx+jWMC3GG
yFCr+FXNy6yBSh4ATzzLHUrmsKsFmXfNe1s098V0l/qW6l/ZuhGBHg6/FbfB
nHxNnB/mavnpfkX5YQl9DusUZkNaIOjeb7gdFhXySc7O+OErB4zxXe3r8yY7
jqAttb5dI0HhxOZq3OX0iFc5f1sFOL30uw5RMLeBF0ulIavOytwd2toyZAlu
nhcWR/8LQyck5JK7rRYwGikhBKC+g9hMvf5oMBWVI6l0FzudMxzPPTIWkVMD
drNAt6QFKRy/YgdCAzRfSNHWb3MHIWYdCTquvWFlGJdBdWI3YtTcgAvqZiTl
/1UolPG78v7L9du8QcaapmdV75IPnajmDVaEqDR5MxpwjIxZfJ0Q0az2YEo/
zo2BtoFUZopE/LZhcn8yM0zkPsYpXNLSia2chG/j+ZOZElOegCd7pbqJHITG
h3Ds2r+UCzlXPLt3UkFEfQ7cQgicgQinPHVIFr5R9hsdML+PleO/dIUSk4cx
M89kOaOxcD15PSDNdRnUSzuc8CZRMQ3tKqoe4lW7T5kxXyZcpPoK5+yhWk2p
Y7uNuPIYAA6XFqXYVy5raFWe5SGAIQBmmFTyFDLg7geMvLcMwmd6GyjcPAvv
1wzPbeFqHj2vHTAsVJtl8WOim6jx2eS3pBH2spt57OUnyyvSYPjlsn4ee8VS
27XuoFsX18V2c9JWANwiHxzaXkK6h16Wlu1DXppxdLPIhjPPUtmxiviK2LtN
tnrm1Ru1n95+FH+aqikKFFUAi1nRDWafsd95ABHEu++KHqK0IkXo/JEK59WF
cgv0NoxLzRPa+mprCzUYZ8UK1sc28D85VtlidcCzGhO2gcU+2CbxbtAwCJVN
7JRLUJR0HHvuEZgKBzAQqfXOkBfnPoN4R7TDucLxTdGj/7SxelrOWJJUjWwB
gqrIfuWgRhf8fi1BYSFEypFXQgu+vKvxJQX6/PVM6VrKOYnDN/3CMhSpn6e+
65JCC236CvtmOYlE2Nz3XIuBYKurMeydy2QFvAcDstyW9vEW2aox35QQdEdj
/kPr6/Jt9F6/1bwfUCykiiNUJvQuyw896fMm3wkQIDDxHYnYV+6JB2JGgEQk
zf2etoiCFBFEa1c1kKPC3adzlipm6xdskhg5kMz3M+T+K7NHrA0Xwn04bZiZ
mZPxeniU8rAM4BApqGE0QFEPXjRuVnwyozdV3sn5oWAlQqVMZsetMz3nmGH1
dbIeGRSuX36c3Gxy4EA/ryinb5V4PrknNZ9LsgMYf5XwHT+KaeP3qBNbL6g1
rzsvyCuI8iNIGRBeNtt9n+C6EmBTr004ZntWMvrRg0ZceSoa5PW4OxXM0q11
GUAmm+1lS0GCi1ab7WYbyrnj6UwuMn0bv/nhZtPK2et69I5/HJ/c9sHn/mtD
7qLRc/8WU/3sQkybTwJSRBxfBfTGLWhCcofnmOv8fyoJAx5AzPq5tIAS9WRY
d5cXrFwg2UbpRKvipxSAOl1o5yctAdXBI82a9nVHXC371KTOD9bscRVxjLp8
FZdCM+h2jilBtcwA/h2fFRp47mLbxlXZh+EoS2SN1/p0njdtKrR9QTCZXmEj
LedBdhYm0WsoBt5Ac/ZcGgYiz/9aIjRGw/SItQnBsneXs5U2cPvCy3Jp6fjb
MgtyUSjlreXDapvvdEoMv8sWU3FPfi2sTHTlepV6oit1HQCUCacvOdA39Tpq
9Laatf7Bw2Iu0N9xoqLTUZ61/T9Us2Hk1kFswlP2rO7ABqbHyCcoC1NCZVes
pX4Pek4xSzvTCEpm5Ac1FlX21whaKNsxGGwzo3qQeNhJyBtq5+0zFOgmMgz2
CEpDBmFFgb0C86AIcVGG/ucyuWcSINvRO7FCXK7qFCdtwPbdOLsIekOPqRNl
XV7Y/IYQgCT9gbvf40laza/yQDMgfcDpsuy2IIgLf4H/OS4HpiTXxy+0fIxq
iI903rgGLQSh13y3aIwFU8UOAshSUuYXHqU7lFf5oBIJ6Z7Jo6/m9NoxW5js
xkksarOFqz8UlSvkuc7Apqm/nbsFb5bjYxFJw7z2LrDajw+kgV0DufqRvfF6
teLSG8oD5LIimpQqJmQ1CTG3HoUK/q1F+pTzpSha0zdKqrjOx0ss5qURYE0p
ko2WnKt+Kp2u9gv86twxoKSDrfHhDi0ghgN1wfh3AM1D3sMmxNBw6Oq9pzBq
Mk0xPIAoy+KsgZxRXl04B+p/TAI0wm0o39BJK0UI8lTO/NT5KaJ9wNr5La4F
/JGnYo9LupgxH/jAU8bp9zWuuOq51Vb8dhxXPa2zJ78wkreyo3lPpc19h4iu
yuqhm6CY7cUwD8f8iKkQxBOD9ZkuEd6itGzKbw/Fmx6t2PyZHV7ElGEfDaVi
eeN3o8NxaRenvqIaotKdeSK7oCFohebrvHDd+ZWwmzE4uFUcUORAHj5MDxNj
7nLTejEl+qLi7uWAkE3sBOSmw5+PjVGvG77ok2imH/gckWtNv7k18LnREuUi
RpHvNlE9wuX/fwLnuqXYB5rGZtgjj0tj3t3pnewNMdDbctjmKf4N6rVXiga/
QcQW06jBc/7a8IDlLPey0rrUcM7AE3dvt//uSuX9h41doqepnDELall5HnYW
mFI27Y6a09kA1EwZ4Ax/TxcmbqQ6VlqfUeJKT3pg0aHz0muBxWvnM/jex0b9
ZKkj+DBUMhK5GJA/MVv8CXGM7leAuVBx0/guMV3ZhenHm3urBjvaNAvt61fK
JsRmliwFHFdojS3A7RZwrVcyxJW7LrBGMmLjFGTXpWJmvirP19Xf7C60NYsB
ym9AzrrkiT4fSd57RCOET3iQFZQGuOaGu3WrXMHiycr1ObG+Lgwr4x2ZpDV+
3XmeAIFvOniCDbypV0U4ffMj4/pe8oZedpKiyDKICfnChOoECNMMhqbf9990
dq44fiPRlvNhuBTy/2rQyiJxWOCuE70Yc2WpzTYC1mFDm8aq2HDk+Nl89+uH
uAdoAEMMXB5DUQ9P29fpr1VWxW7hQSZyFaIolMoodYO+o1TJkVFdyrtvsIB3
pG9hd9gdaoHBwMpv/H5albuzMLr70622QtQAnPs3qGsh7imAvjluJuV/i2Fw
fEj3VHORtCU6VMuZVjnkZWr10S23MFWOPSaAwQgh0IahOd2P3hEjCT0/mfMO
JLLpyKTPD90PLqD6ssrPDv9LuZWxp+zOOB6kWn82HzVd5sylyRb/+ZqurkwU
jReaeQXn3dainhta2c6wVQWrODAiTSd/wqastZEowGT0EXq33zAHvVvqsvgT
Tpjio9Ku3sMS8DBydBl8wrFh5lVbeWjSCkMzSVejlqUTyGJIUNPmL+ZSLken
tvrWDDSh25is3ETWCS+hxtIKFTjO8YvpE8SbgWQrtLyTLr3qeEKXqisG+gJV
vbcWG/9g19lbnDkfUv6YihRSG/ptnTF029kzlcF57Dz9rBemK4T6APdKybi9
dfF1Ih/M9zs9eeN1i8DCx4DbGx3Q17KCGy89PZuiS8PBCEijzgnzG/37lqZw
mXDUY4VPpqbL2KqywBGeXsTuVdlgd7sqW4Q3vyBeV/RefotTOLcVCLWt7OEG
Bxg3bAlr73wzpvzO0YmOO0c+d4Ym2iHI8NGPDKNPtG13kOQxfh8E05ZXN/eG
PGoGrM3j4muYcNa35ZFb+Nyn+mwMCRWbwLcnTl95Pcv9ptuw7St4xxsB3uZx
/Abe8PzBzaHm4BsBFJxYyz+DmXPkOyhy1dEj3lKCOaF41u9G14Xq6jv5DBI0
K7Zo7nkcK/M1TsLHz+jD2N64fD1qB1qRew1MsTwPWYfdeDmirbPQX0fMpqqB
plo/LznPe1SXZWZ9Dj4QzY/eNgGZeWjZ8FOxWYlvqNzXrXoWyb0tUeMGybNQ
E8IlzisErg3Oih/3v4DLJU9wsBTgx2epKJ9VQED4u9uYAte0WRHX7rAJ6Vs1
+AnZ6kyfhkquFGjkMG1/daYRMbilUNa2QWX1eT95t/v5Sspze+YOcbhbPYbQ
/ko8a8VUtfDnNqS8FFCOMuZhFdzRgUFVmsKjxuigSK4CGcpJhGUufxJspC2I
inkiEAIgWdpMBkercInKv+95/haO5DyC49P+1J/NjIF2byQlZvzqsUow25jK
xgalKm6mHXx4k9deQntMl5mZco6XoHyn4pzJ2lP6t3T0vX9w48qstI4LqE8V
O9mpy5FYSyJYxAIZE2fkxq3ObkWHbKXr2yTvhsU0FdcAnF7fLbbk/ZGK1qf2
Q0JrN3zJwA6YsjNEOw82dAuCSWq87p3ZdiuZplrFyontDe/9fVz/VGgP2oje
4c+dpqIzJ0S2RpLq5Abix4L8YD8wvdETXWx5tBgcC3CvwyVtN/oUSnjp0amn
tKKpy7ZkSdcqoOW7fsGtfYoOeYZHgLE2DVVcFyvwmNsMYVZlhV/UbanfwntK
wzH+Ot5DdFQRnaX4BInaJGhjaM5REDxDjGIJMHZkUAC06WEzauwmtKD6EHvX
7AqD6/xEwzBe/DuE3+1eHjgHCUl84fj6EuPZ6OXW9LcVoMLzXF+ux1dUywVV
IFAj3k/t4rQoSlwKF8wYjdCuEbWfVfocXodFcetIKeWbTMq00MWkh4I20lM/
ecrRxeWyO3gYwtj9H0ZWUredCVKg45y4NEaOeRqdRg0hD39SX712Thn0mMcV
YhBqsHDsBap2+N+3bD7w2x1wZworNCWjAhgqbN5VA60V/bQHpkocM6Tth0WK
qz0IhAmGrunEwUDf7p8fAYoKTknMsAy1o84SZzQ7uIKa1Y7n0WS/CO2swo6D
85lbcjlVw+TmcCcmVL9/Rs9zp3KSpN9/bfN6FvYSorKjWETaHVC4MOiQeRfS
6SDu6MstwncUBYcqwEt+TKGhd7NgUQhEbTr2QwoYVbxeh8zEP4kR7LGs8gfw
PdnCpa+6lxPNod93ysggEDWKd9LwYopQQ+7t17BVzmapoF784B6369xKg9vJ
qEAHtCJLZYRLtRsHqnwsL35+7OysLrsWQr3TrZMvuSOdwGqm9wnxFPjSIGcO
VMqjOr/+fDfYw/Qf9P97gVYUdqY4i2XLtSb5PhbuDlHoIeViZ89/XyCcT5sp
hT+0u5HD2uagTtVY3GymmxY76AhVMvIKoiJS4iXHtcsso0g4V5sxd/vAsd/l
2Y4n12Zt0Z/op2utPsbHgGnYPFu94QDSaTgpUiuq3/k0vDcBTGVEpGXu5Xt4
Y8gy1T6c4/Uub/O/PM2m0eOFo7Tbkqe7R6vJVoFZcKoEJ6lZfAiPmll5kBOH
NMX1Ibk3H7yagoaMN/IqAF4WrhVGumnvg2lbZcoiBE55oxhZnioU55NUjQls
MX7AKzkqo9kBnnt0+U+l2LPw3uJ6vbUACzKE0TvkYV9FhSLPT7FV6awGf09n
4FG1/7aUVKX7PiezrAU6gWND8UjJ2yLmKxt34xa2iKHMaGJllOmnNbP14AO6
ObTC0X+3uGyYOoH9ZI5dN/YOVm3LYXF/GCMXqA1k0GCaW9QbHJcAcEmyBmY+
x3yXhaixjEa9dga83g8J+Tz7liPNTEMxW/UeHVUbXj5FbPqIHnQbl5r/E5Yz
f+OrPHcCpIgzjnf+NPImLF5j1EKYZ+e2UQV5Uf+hVb5gYcFfcc+y+T3MC9P9
Xo9C6+Ji68mqBJPjEAd/hHRH03Ol9iR3lvK2Mz9lGdynY4psCW4MKnqxxsYM
V+j3+Y4bvbdr06Lmi752hf/fpeti+DA8kxynq7gqCNjd/8SYWIt4lqxjJ0gJ
nWRwyMbH9bSqgvwpAJhHmo4Wn/9BP540eelt6x8v9wQZLuBddHnT42sDQbP3
64/95YJRHOmkE+4PM2M4lELcwWe847fv0Sk4yPaHrUZZhuKiEnCkm2dhM9jX
677Ye9SyJyZCjjKm4gCyH4jXCED3zPHup0kF2q4ZgAAqK9tYnxTynsgEiROQ
wpjR6hxgd5pu08Dpd35MWBxZi9JFubC80fRAbcC6DM0Kd2xV66GimkG47CtL
jC8Q5sBlODZuqMOQmYIX4yVEKfM4S1OQY+gaOgklgfe1QkB13Mt4tlw4IdJ4
eaeckbbQC5D/A7DBgoqR53CPCjkMC7kNjjAzSg8pLvcQwCkZIdre88SRK+2V
VJK6EIa4GgnrdtTSdO6rGKOQXryEJeVFNhANIbqBk6ZRfpum1b/ec/iPaH6N
mEEXh/fVlo5L6FLZaeh//EYj6V60fDdm5cEi8WjYhcB/fQRrbmPEp/pWEPwe
0xfw4lX78cvOAPf1CsVJ2Fl/1GrHDVXfT5RqHonCb4ST1oV6NTg4DAt1QFM5
9yONjVqNvz/iJdDLlH4mw3qDRClxYiZ0VFu6+uKJKN9L+FKdGXlk8Ijox0ff
PyOvxxJUbggmzbeKNo7ZLcoYNhgukxeybW/1cWFUU9La46u83GABoOB8Kpkr
hsRkqPD7jufIUu8tp8v+Vx5IzqEgcKrotJpAoETAaXnVsmBVhwZt+7jGBa1U
3BOCWslRMIdK6WFkXEUYcRwa98a3oZc6nwShOMIMk1SJAwwaYtBdYYb+Ire7
hAz7uj85K3lylCITTD2FHI9sY0S5Abih1TUJBCy6Bag4Az7ssCyDzQkNWik3
s6a/BClVGAxQ8wpNKbR53B4puy5MChCzbUmGyk+/R5lpXMnj+FOr15t0BjOw
/GynRQLkpgD5EWNcCH5GY/jHNekXwlPEPupNJhdbYcURd4QhOfVQ9mcJrggq
O3xXsXh5tJI4P2rM46lZWopyhIeTuEEySMDBVIZc/qiSWoTOOIzghk+rCabk
Sn8u9ZKkfvWbI6xzPDZEjsX96t51+zxH9XOd9wxMw3MXcBrx9kqYAwGpdqOs
gqlvY8yycdPpC03bnBGJbRgMgYrj65SKaxbL4DMZB8zxdYkIpp8KMOInotku
mlBY/CanEqyUBiiXaHQPAEqZ8UQYAATK4/fOY/IETKJuKW4E0IliPOWXs6yR
10W7snNUEMBzbVxnlY7Ui63ZEOynT7ItsDYUdIrQypOzo/yshgF1EP/0hkip
nvBf/sOJbuzERWnCkbYh7fTErt2mOp8gUqOtJIOvi/sG1IqcIaRPxuhgE1mM
s55wGUrTqWBBR/RuNc52waJ71yNDrzfcZxWlduOWZACWy4B+xn5nXSUTTQQO
LjDnl0ILt8GREuurkuZ4oVN/lSZhT0YfOoY0ivU0Fdi294+2e5GSPKTQI+ew
P4jNiCwRRe85DBEk+gZKZioA5cFzg5t1PKPFagL7eEJuXbY1k7BBQnakjSN/
PVK3XOnHyStnLjltYGoGB115W8fY6sAPnuQTrYhHzHzSEV6K6cBf1sOzDOqa
sblXH8XM2eOiMGRhVfDYCFC88hp1bC8raK9yPwNF71SZb4bTpDI41CJ7ihNk
pPIicFifBhNiNEGwwg9ICDhik8l27Z3KkW9RhStaBmaN3k3DY9ROdJG2BlSw
1n/AWHz//FwPLhEM41re1oKKuGLTCQ9jELWyCKRxsWROoHJRYelRBM+OYir1
7onF060MmK45In3fjHfeuvlM3U345dKProBvHv6xHHNgMla+tOndc9ikTLex
sSdIKQ2Sxx+K8oItVJ56HCn3SjdapYhocDo58HsTmWNKIoK2eRzt3rHHDEuu
DYkm5JXmx+SpxxGWni2A79jhQf/cUl3esr9Cl/HTvzpgBpK2lKQZ29q/l73Z
gYCBWiJHUKbRGEn7Jp1P2Ywe4O/qP7p9zy1BoTW0uhbrDpqfvTb1nZFoiq/5
hoNduy4HdpZGWa1EiUt8bQrUXEPJ+IupipFgsCtqXGIL/IWRqMAe4Mp3XtTH
Q1SCJ+wwmkna7rHXXd3O1TSyzEo8C6N6SoH55KHzp09smvPJAriGp8e5Nog4
q6JkGFeSyuuox0JCL09gEifd3T1JcY4lrkPof2tkL1n2C4yQdsCxhTsWdZ7C
IMP76KeTV59g1NhaQbsYFMxpModbdfZ8Ini59+Y1gQOeWFcAyc1B4Dq1NaBN
iMFexS66JF3cuwrUTr/KII90CzfvYvYI7RVnWaoAh7kzBdOu92npRlyxvSSK
sSygaMJuM8WSyyO0Pdi87uTDkEBoDD4bd8tw+z2PoQU9U2rlxFpcsTfWEkcS
7j1vEDV5tU4Sg6iPsGiuzEDdCv3abi2weA11cvrm2XJXHrZ11udMQhNyN0jQ
Y7zrD6oJ5QZMdG7PyOLXRf4Nw7DVE26KHrLHNMazBun9K9U0txIo2s/q7OAU
D0t0LINCwgaKg6jjOC+bv6WQKivSCXLt+P/kgLQAGDl8fb1ei0vwdlojwZKo
Uac+IxzAQ18Ljqz0BJ/csQOLd1SrhAiZ82HTj0nGKS0gLoI1M36z6ZWY7lcL
pZ7hXeFfm+R1KWlr1CrGsQhaTg7ZDHn9xRAHWtssNAc/1VMgboahH6efmWsB
uezzTfn0b2UL0o54+k7mjwtgoyH+Nof/+yIA6nZlwrx9Ion6VmRjRqMfSj5x
YsBEElRxhVM4siOsrK6BLVYFBhoFrodRI5SpJQuih1NnXNYUEqN4Mk31v8Il
2wzNm3xIi30uFN7se4wCLWNQigJv+u9iY1mJy4tjRVxP7jaUlbaANT3Lo5zc
Rwt3kOXay0o23ZmjTJadvlV8d3JpqJzDibfNli41hFnAWS0+qTRopTiqSstk
L+l8NrX6LgkVkVkg6VojsuFG06T/bvOt/lrgynLmwfCSaPkqZ3aXZtU1wDcU
lA4JxvtsMGuB24lx4f7V6DkzyKs7SdgRUCaNTdG08ldMJmq3nnUgvwmHts5b
GiZ5FqKO14/YCx65gg5L4+e0bH8HN1F8soi/Kem9INETJLBGeDkxlSu6/Dfj
CgnPsP+42HVJvZBsQysJfL3yRKuqtP4rudqiXWjsoFqaIv64T1rrQQRrTD3i
1CRJygerWXN+u3pemUQUbSyXIlOy9Kq52QUwYlths2LknUZkBXxPO4QHric6
BdD2ptuysVc8CIC3HCkbxbLYUXNGbLinlaKw8BiwOJmEz8Tyz9YtIR22gnHd
qpwG+tVPZGqlgvJDzBXc1DGkHDekG+IpsjwY1Gh+Knedu+xAYvTVSUnbsRMZ
7qHf5bSBBMVogCBRRjROSkHMGpMf2fdBYPIu3aqjDqD0T4zsRxmBmkpw5OlA
rSNG1kj7Xsi+hwpEY6q6QZhfZCge6KTcmdDUtuuxlowDOpjgP2+s20veCT74
GGZct6YuhBc0RYhNw0vUTL07lo/DX0U+2AlyJRNAQCqdQyZs9voiHxa+uWtB
A7xlZq96cDt806YgwkZzj78MYE3IWkmwFWROEoEPNfXBVyYSsa2RnMmVbmyV
siCoxXdjqP5352f0+OMM4IgB50zZW64TQkS3Kk1FMR3Hj2OP3YteaWzS4G8c
TnmOqV8uZ7fYw21ILfleG2Kk/dkFWBcgofxtRtXnw3/vfqyAR8j1Nx4vmcCi
OlrHymeD5EjVwZ54pXpAypZ7G3Miy4OGn0oetdkvIStkQD7k73XB6NtrP75P
vuDxryUxgCGXhBgBj9VL6HSQRrjOdMNYhmIzMduXgfNTJDSi+jqTYV3JKBUo
PThmm0wY37bJa2AJqSG04VYkBP5JEXOR/HDOuxAqJ2z5COQfiFaYYoQm1ydL
6c0PIx94FQ6habWQRXmq1dWxhEn6wRe30+lfLLVkoC9XgIoW+ESk/4VyjTeP
t75uuXSw2aovB6ZJZQFan5bX6jJQO7PZGf3840uCTLzyufi6HXger3YuhLJ2
fg4GOXfL3W3fLgjZUA2+6XiZ4vfYwPNkTJNXxyEYkJXZXJVJ2YDkEO74o/7K
QeRjF9t94w3uMP/LeKzEFliq4frvvSVqg8DvXxdzlAt4EdDL+7IU5oOj3S2r
fYBP1Q54rDofO73E7QUkMxQlb3brb/ofllHGmFiscRm2fgBLFQlNJA4bJTib
Opnr1DJdutSVuxhgj2fejvChakh1meHrFywhodFdMr2JjU6WjFpfLvv0fcLb
lx/s/84mLD/Rr7dvfJAQjFGyVOBrzl2jtO859VQlQUsIsXpmCrcOFy1A5sS3
HpflfPOHBNxtiTuzh4x/9qRaJKXM3twi9OBmSrOiYNOj6QntEQnatzdcc4/k
Uc/wf9C91i7+gHRtlevjSF8R0cr3eCQJd94saOHqbVPGmedpodapYuuL4htx
zNB/3ZbrCjbZSkubXOgHjcrlqR2HtjKbG/+3mYpIgbMn0tRDoKdExaXlUgvz
COKF4iS8qAOBLusGNWThNGKCxulKT3crEPyjDyLqi3UdBTrqKGwlGKo/S/s+
QrpTDvyAlVINPXySXsjq0/6bQsZHRXjftmtkMvPZQ78mJ5kDe2npBwnWboRx
gzu3YvAfazASuRjLHf4u2MJWSezz+XIsJCrzQaos0nRIE1FxyNqPEbRGX+M0
1DSew6Vo1+5kJsCOCo9h+N7PzY7Lzcl740mdU11LxvY5ZZImlbTX78grDXe5
OfW/1LWJ2bos87fnR7IbKjus62k/EPlwmQtNvEe5IiAcZvd7jA/VC+fBQtpb
sjN5ipRliDrpfUiKXKGLUHswr1kw2iRO/waCNhgbO+/65V1xt3NvtxWQhzJV
UQpcTer/yo1Z2mZGruV01LuOTIWaHN/Mg+FBkGyduU2T7rpbD0LRGgdvGG7W
jTh53RkZDINjbcaUnq9B3z8sHEtclkshbPOyX+qd50CjYhhUHabGtCcySr8I
Sbg47+/Ubwy/DbCgREKVG6PucW2zgMxQyX9+rTwIH22fvi9vH8YUyNYwJzO9
T1aG7wX+yB+kTHB7qFhOwBFchVdFkVVZshFEn5oGGJjg8GeMM4bdhVt11Ran
syQ70bmsla6fJkcPq9+3hHiuK5dsZR+w7bHdgutDnlr9UMiHfehtE7zDrolt
zrNfPISdu11SfqU/56S3oldfcK3zpebxM6L9BLDJwi8Pv6UUF6DNMvN19NQB
QFJZAZx+URP+C2aPBvodWDJp9smJNY0CaC6Om+cRtFZVc9sEYgNThcBS9lUm
cjptv5ZiiVN/kcMk8k5L/ofaeSha65TlogVxs3mln8Cq+5oVpQEOZiNGApBC
9lwvvVL1ESsv/zp4ES9/xEFlfMN62iX/tlM/iATv7YIX81ECZyJR4Wz2fiVa
74S5lQJpizSrz/RK/Z3Rrz+Vb1pZO0Y4KYAFNV8aGt5OZLh4ZiXOCWZkSQ0i
eQYC20tvyc2A/pvj9/QKhwCqhNLQB1vgkCdCOXZAp07/BzyEzD1+wur4KFj8
0wxCrLo1iEW74Tw70YeQCaY5FY3qm+2WPvOZT1GMmuQtOdhZG4j9cF8gv2G7
g39yoiRTFi1Fha6UOV2qLFszn8CvuNnUz3u3nbOkxFJCyiVeAu7ke+kj0Ues
8XNPn4F1Ol1W5RaQv7bTe+PhOeNRlEmPZa0U2pmavnMCi87AfSFqPOiJsIDb
U92pT7K9wo4w0xUE305v7TJekllcX3GkpsUB/5somT96boZr74pEYXx71H1X
cmryEOpd7vGbjl9OUt4QnKiYvmLfAgo973PA5FZsvFG/Md9QhTV6/C+PmQlR
r/Z34T/8Q2WYft99tzw47SiNtKZGoLPX+cs1c1cmNNiMTvkL757HRMgTY8my
+qlQuC6vAlKAgcs0CCQldIkZCeapK0CNCOC/QafTTesFI183MlweSJNADBOm
rjJbJ8oKwMbJqfa02qPS5z7Ha6YmKdbv4927V4UhED57oI5OcovX50xABBkk
VNC5OjKph8aRM/GY0NWcRBoMoebpP5rM3jUgcrTe5+4kfRKij+NfvLIXdLEQ
wmyvjwqTKO1eLjUVQQ3cGKhQmRmdlquoRXEPY60T20KotSOb2AGpWPVdroKg
JiXxTgusjqKxmZFuCwksqeyBLx6dj46l6bZUHV4gYJL/S9hJft2SvwGxFQ2z
2xrWXThLMKuYJcxaRemkdqYv77teneD1uCsa+1BSCGZTlu+LkwMamXFDFTUW
lBFzJqzGIxm1Rh13csfsSbuL7lelqDgcZDGGVtucu0wFycF8Gy/HyucfLJbj
zxruZR8yOZUMqwIbDp2LJhXm/14uNX6jb7eoqNs0/Rw5ZM6wXl6YKtfDnBDN
djaeKcDwC1SEiRBRjxbG3Ybmn+7jxzphDbwYm3gFsVwNAhDMvZxMOy7i7KW0
fnQNxFBePftQAsWYlSgeZexwqM0GRXVzKmnUhMX6zOo/4C9Vd5oZxzEFHAMu
uChtwE47vC6vsPXyMI7mhlMfvhgQaFuCmL8tWbDoH2pcWnTwlB0fuWoMfUJB
kNxtdDaaXG3fRq6sE55pfQHp+Hb4f9Rpf8ZCDoiNeL+AoYRkB1UyTzxvOE74
/4q8KIIQ3ecV3bGjsgxZE5PAECEGrZe5mbx7oc3VpTNU4aiAhERIHDJNS2RE
Mo+uyvGG6DbKPeO6PCL7CSfHUS4SNWSfX4UDoBPFCaaP0FhQysiviwVK1KpF
S3e/MA3eEMbJOBRmyHNcA6d86/fB7ZhMtJtY+1RvfIy+o86HN5W8s5YreZ8u
ICvn+UwMs6alamwnMNzdi0/B1aTwif/K7+ry6QEgNMz/wECRNaokBaGyHHpC
2fSNqdO0UwWMLkeqfo/lDD4G0UbWgIS8l83622NGm1kc2EHIzDnH/FtA/AW9
DWPGtKW3PFYNKZX7QSX8hioitQL8wXgkgErxJIDb2OJSHvpZRWXwPNv+vsx2
y7YKZtveXW5EvGjaT0A8W2jdhatpsFNsxwEThc44QyRFQSbRGUXsuI7+b6mZ
EvAMuhN9Ng2EXbDOGQj8acDf8NXBHj+xGUONmVTff9CARJ/crLUPHQxeVvN1
sHJedwqPSp9mI/ClkHRjubJedT+HCZlhh6z8JwJfDNvwSHbum02BO93PdePq
cFdpdO/3sH1KKpUuZdPaDDoj1O8VCXT6Xl/zjtgSYBzfslnoRx9MfnH6QVY1
714urHlOLBg2xSyq2Cq1842UPTrEoav0y1+nT+u7XedDmAmWfiJNQhuVy9e3
k8GoxxZswdS6UcIHm57rdyaDpqgl7vLLUaQPEBVvLLF6dPBifrXJPmbsAW3P
Rqqcr9zbmTGb7D2bAkUlorC3UJAG3Wo8/vdMmOwtd01KL3BiXEKZN+w0SyHJ
HQpkb0bTd3x511zKhLUpJq93g0OXn5/cTqrDJwsax4hz4WKovQmXSIBM5ClI
L3w1kM2SBVyrshGmf8mHDfcIbJIkqvUfby8Ru1riQCYqX7V6thHW/SHKKieW
n0yA+p0ByKDReOkfqNIqrocMPNWAvyGZtBSUhyUBv+pWWc6RcnHIcVQLZ6T6
dlYpp/5/Tbv1OZikCIt/vSl0rjwIWX5Z3hcC0Is22UT5MJCqEzianpWPsSo+
NYq9BB18crIM8+sk+StXI9zR8ygowS1TnmxLMVA7DVVHvvO0eNNOpveEhuIE
1MhynC3VJiHtUB6B75tHgm4swpUMC3H3D/Sz+G4RaKWqFULMm873wvjFdhoh
Oo77V+ZpuRMnFFMu5VX37+YHYlgcTTk83gc9+JXYUbPjKFCdr1TTd60n1FYw
EabIfQCnPpxBdWw97vGIvl5pug4vsPykRslX3QcVV2IPYYBZtLtZwosx96Dl
q92M6wssI1hBy5enMslzGJf4OEE34OaHS3bKX0eQTrp9QcT/IWxMxGZd0cKx
04xQEjgroqRGXbtv4dokwMwa7wSpaciCiIVxkBpDBmeg4rcMttIlUnVb16u5
A7XMR8MhH1LSSZWLi3LmxeVZ43hkBXCOe5TMFywgpppJLHyszE/I6nFkTd+V
7qxuLIrhqLxVjVH1Jw3I3Pj2+BGCacP44nHOedNiAMna0O6A+38JoYy06GIz
1hCU5ZXYl4fbEj5/bDZeaxxN8R3vyyy6d+6u+quJ/NuPgsAKUZKeNyH5Qa6E
pwrIIhKT+ZeNAsnPfFcih+ITgcDvn53PkC099z9RNSiT1LlBm2O4hpoJqMvw
f30lsUuALQuSZAzq/WVAAUahFQZ8Vz55sQymzpu+HNz/OKL1FhMV20I/RvMf
TQVVuPrS2DP4iBGmYWWdZ/0LZRCHHS8BxI/GJFFkiwkc6yS7I1OTgNZI4+c3
7kZ3nVJ5NCEDpwD26Le/r3BvvuIKTXz35fiV9NSp7TMekF1zMtuJFsjW2sJN
Mpx0Ezm+iEKyKj2sq2BifbDbiMpv37ZJMJvk4Pg1fk949DrNmjLvp2SJejjM
LaOq9QuP1pwGXqU0nb8eQyZS+D+7L6n29VGVf/kwP+XNvb8gHqccGaPFRIIV
INM8uLCxM51SbZwWO6VKaoPav4DV4BWrAf+04QtmwFXj55HzIqMW1CkWPHBX
96VdRK3LiNwlAb6wGvZ0x6gxW9hf5C7Ly8SeoqksHQyoDxVgLU77mqw1c+xf
H1MJN4iq41zyTpxEy6x7gGzuSbV/BGIAPUCcNKt8fpUDnai+97YqS6Ih3/ak
sioLm5kvGTUkmpOMNkd/Xtj6jC2iw+yNhkaoifEvYnCGZcxLEswKhBoyTxtw
hCLzTLPssoeztKDtlp3020czoGF/8PC1Wt1G7YdB9XePWbpRfcaE7htf9VIl
1P0E7tF/723G9WZF8pRteps39ya5o/WsqYefIypk6J1RDremDhijblr3uje1
0C6HPPn/JemSLWIhIbPGoWmXSBp1OpzZswzufSaBYA5/IsESCr6CDwtIYZrQ
L3PFXUpPIXW7a7wGmvM0tJysLhUmf9Gpdx9Aq9w+6C4LQP35bbam4KC/X0vZ
RKQ7QNUuu/NyV6iyLJWgUK9qTlFVD25wVVIcUUTm2E7BxBW8STlfRpotMel0
DNPBFwfNdoyAk6KuLnQL5c12/Yke36jrTBCKi+vsI6D6v1cjq7cl1V+d3F5S
hTUt/wEZ0cR66meqxQ7qLpEfvXx6E66fZB3JWG80gdDVt2xM5qqdmQ9/Jgu0
Nj92jVoLhU31opt+3UeGIHcosMi+QHMeBn4tZWQm+/Ep5PgEmHmaqAQHHQxT
rC8iYmbiUmHPNCjpewi/e+h5nOG49gS064WMBaLrKRK2lFTnPbgadsmeeTSs
IA4fWINnCt3J4JZJdKplCSJOQX8W6VcwvvzwEnAIAyMG6SQ8tprgdWfGSz9K
R+RjqsTn8n+XGjgqVKpvgzvqGR1dRpTU3er0pUncgsHqcBAiS7zC0dDj8dC7
Xf+Q36cZTxrkDQTT2znGrTN+lXKrAkQKU/DOUwPBHqsodjA+stum/NAtkmxU
cX0P4oajaXR+EdYfaLJAbni4g4OFuG1LxoSxBt5RCLYyHOo1h1FpBwT23gSh
mLoakX3lVDvpMXGEjmrLyBHiwToqm4SRrlBs5WjYK9veIhcvLVZcJ65X6nS1
t5XOe0+X+iiPaPobFwpmRpzHhx8NpySdjDztIcF66tFDHmy9htcIVphi5gZb
2dT23CEdqXm9tNjdr+5Iqq4Oy0P+f9tNMG2SQiU5ddqExXxkRxiAc8cTCBCx
b3u0LwgpZTDsqjbU0ETsjXZ4f6sSabRDBoYyQqMMSIzGG+zNjrtrHYPW/6Pf
Ha+Qac+AaHXtMzgBlc6cMFrLXvN7GrziNNxGbmUjFE8QqV6TofUunQ4tsy62
Q1AETAcf0LJztmJ+IfpxqwuWtBsc/eMHxmWkwvMuZ++E2b5BJTLuOZS9itm1
jxve7eiPgd5sdb471I985Eo+SgpmaiK1t6WjkokNuaOkP4TqHDp17/HYsAgU
32SIWAbsjyvusjdiKqDWTPq3j8vDZAJC3o2Npg9UouXWYGS9gJgaCTRtzmQ9
Rgh7/M20LDTrG9j4SaO+GI0HYHphuRjy6sIOTfhnj2WiJfTDEnwA5DuJHrtW
JrMqusKL5+cn8ywSc1gbp+H9jPrzFxKnTMQfYga0gDgvqgHNYcldzAwSmqqQ
DP+dFQ1jTr0ycrBuySXn6fJYWaBd0kkA1u4Q0yPiXZAl+W4+Ny1AluRTTjrF
Zny1uGsRvRrY8E8d7igS5ePdx1M83K/8ZIeyLJoBQxYQVFTNoVti3TdUoxgT
bINU6Ipdzti4EPFwZh5lV43AqlLRsGLZ1QDOLTK7lCCjySnB79WOtJkMMU+w
c/R1nALM7hzcbK2SyxSa2uuyo2gQoIMyKUq47kQ0tjeGJH938lRSIFBGrSjt
EoArkQYF+IWNi8e+vSHgHTmlMz7ULnuf2s1hafVQadwjUhgJU4BI4IIYoeoc
5TAUErmEryfhps2xQ582WwdkUefZiY13Ch+3uBxaKOLLKiOkxEweLef3IGbw
xpYUeuahBAnjbfxJOerg7maS07Lz/MtN8BoZ/kD7aRU/hBmxZg/MNUcjjM7G
bm8u6xzfn9CR0En9Z+aFdCf2XCWAIeLuGvNp7M/nxQa/NHxLPHSuvsu149gV
kW/7iteEmPL63d00iGwbENh+j4KBZDa98CSXnoedkT2RbsX365uPKcq/oznx
rL1enoRBn0lazvgh39tkDG9aq6BPo/AgOvTUaAiUi75alwMAViP2O64f4c06
zHFObkXnzhX35PEl/4pTB7Jr+Z6xwdiNwroyowxjRzNg6rA5N+g0m7KoeoBH
22B1XVCvgmhTG4SlL825m21iJDLMmJmJY20MkPn6kQ2KGTbq+D3o/VWrjy94
xUbXpXXbhyUqZcslKGK6W38oj7KLxBSIQCuOBvu8DyCbreYOJ4kYXLlHyQBK
72KGzv5LODz7H7x07b14e+Ltv3rHV5T6RLrNCqN3BQW67koLqQNPIXhXlAmg
tuACzocGTHNcnofG6kAqIoPe7cmj1JbkoHTmO0fY/5B8zHq812n+cBBSK8t4
CXXCcwNLyz2/5NYKAlzw8aGXCW2ysfu4UFgJgP/zch+Ad4niIxq4kBWxmdkM
ANNxvOIMGySv88FHq6FO/ArdAGnc31jx0SkTEDq12eL7fl/91Z3YHldDVFvB
GsRclbB3zv8gfwcC0qRSe/o5c7pLZMHyHIJ/AcVSDiGspUXVTb5F8MrO9Fvs
6IFf7pHmhSEFeJ6HCFajjBMZwturI9QoOclQ03q0OQLPCQrVj/rHjp0CHzSr
9Sv1YdejE72Z6zu2PG3xHlAopOBXM8yX/39dUx4gng2cI4LiNGKsQR5+uA3t
AwBaJ5mas45A5bVQdspVWb9O25jngLsgfiZzyVMa16p8rCkmS5uZSD2nXcNY
hkukTaZhyyxDWsyn8hu0v2WMA2nHapX5k+erFLa33umeAejKSed73/kqkRlA
socEUCTpbzkA6InluZGRWsFBKq0qoovFmser+nCF8sorvR42g5flNhfO0W6d
1aWkXrkxRclhYw4Fydo5fKYkz8Rm40j/bzsLwtAZw93NwqqO3gtxsE2hj0kG
8xc/Gas1TlOB9jLVL/JxKlC9Hmo1IibgpRw7PY+wyeqv9VLcGafO0zASH2MX
8f6+PBhiuLY/QP7mAcruDVQLX+cxKYvSikyWOBltoluJwbHpnN9rh5h7rw0D
lat0P4jRQYpPj2JsYvTNGwMUHkLAlm+1jZrR+bnPYx0+ZEjyXuN9XXncAzm/
btL18I68o+ttb45JTzx0gqLCJVhiMSZyOyx+Xu7ArUcfG5LkSgwvszKzdtla
61lHQBexSNJoVqPZRRmMGy26iOjADyijJHL1/DV2ZnAQ4nl2za55IKZDD2ZP
TcSaM8xTvmJ6Q6x2ZZ5D21jnv2rhdufMCRU2zQwps+WO9J3+AmPgRoocphwT
tSJzIzUaX7sF8RQ80ocugP54WPZHQ8KwbaS0ivC7Ti0W66CNf81O0gIYx/GN
fPfszATTnryRfNjZyzuCtq86X49E2W/zCyleQ11YBWIbvFUb657dzqxCbPMf
CqOrgewxOh1oq4iPDKHzOjXZFT4IncpisaDJhLLbLgmjlgf07VVpymYEnJY1
y75NOuIbi9pvvaQ/y+WdzSdt6WkIBYyhCSE9y4A1PSPHpkYv1J3Vz637UXT+
HhgQjKs0vb70dd9KukSh3TBGPHAbMytdZHRtPLH7pMwAJOt1kMJRQBSrTcCj
BhF0fJGg+gt5X73qQaucrroRyEpaO4BihyN41goOlq8dq8NdbwT21Y0+RE4+
bxKKBuJ8mSP55bKtyGHt1ns5quEemQPrcSGjN43HKoVmMaluCxSKXzsf9o3N
ONQ7s2jE4qiFZzlthdsT8kURF9jnivSjZvIxHtRAbdmegNxRqbGiis8pUmcv
ndVNT5ZJXlK8e6He+Ww8AwnAG442Sct4AH1J/LQLwfzIFyM+u7+FQcTCMMMy
+/Ip3gO0W/usq7EjlnKTkZ2WdsrkWjPty0h6xu86x6V3BN2Sn1V7m+UGBa7A
JdyuGMPzYta62MQgVbT+2ly5uHRfYac5RZFc0UhwSI+Vqxl0k3/SZhtLfijz
Zxn1TX1ea8xOHMR4hrZ3CPHkXLOF+b2anW4gIkzTngPp6U4CAhtb2GUa7cIo
dYmOj80sEEBqR2fnVHeGIyVidY0LogF8n9Cs8kJFMlxKV6qgVR6MbdY8IAUo
rI4weg/4As8fldlwAZDKxVc/y03j8BvBKkf2SxM3INGdCowUz/Ozfhc28aii
LGdglrjOnmz48XQo1R1NT5ZqpUIv3sJbrWKj8DjtQEXzznMcgl3XlOW/P0Tr
YZwJn52VPQpU+LbKisBmVQzmQb0vTgYY77sWI3LbsKG0Wj6EZVA5QjZHo8Jk
30hXfRB7cyz743MWs93d5qjN2Lk8pepIdTATYx8kB/efSv01Lpcmv8Ns7L49
YYAMUKskwqpAqOL82T5SKz51wGC49v9b6Pmo1pPxQ84fdxcgTEEF3z8bMcPL
ksXwk7naoF7v88ZOiE7EjqWs40PunzAB4PlMJeikqwG8xZQHEr2K1kxzNjgE
oyBnjGjWSc0IivKbahUKtuiJXbogoe0aJSNad/5+fCdkU6yKeeuGp452s5uQ
ax92WQv2CYKGLR5uQIqnSioJun5cMA5Rgcp5dEj8AShbFEmrtvWmbZ+l2nsh
nXdcyvau87mU2VA8VcFfTd3cm3cDv8OjCx3sB1K+qPjy37erde/lG9ClDsUq
fixw1XtIeZGP1TC1cwHSndhs5vinNcX4nC4kw/Ooco7NR0/f2Qwf9TefgsUD
rba88dU1uiHqfKn/YioRC2ggypm/Ko9Ks4rrapNlx10TBBTmrtBeJ/SqXbsA
gu81pp/DISI2FHY3+4fKBEp9kzsHb5phrqNWDXsaJGgxZcctfRiRWxzpr6T+
HLh/pB5HxD6fMYl2+Rl4SLJ+UE2ce2DiFBhG3HVhg7cdrx4dNFW58HIiiPaz
K/Zw3CK09ftj6sN81ZLG37faqTwCdOvRi4pn5qzY75DrZpxmxtEFTyzS8FoQ
eYlqjJqRE8TxIGgIX5OKRGID5CoT07RrY65wKYt+oW7ZTrmsz6NyYUr3fWT1
+Ej60Qbhi8nwT14fClu2CjxSOZ8BF1OOAfX4e6qdaCJCyOMLB7ULDf+FRbed
H4LOIcOKbRYozvZOzMNS2Lzr0XZZNmApSpCcnXkrcl3PmXz6TagtxoPXulXf
/StEDlm68cuf2OjTdcOPcBIlCLoWVuZDJmar+omjc69bx7svsWyQ3Uty6auT
klU79jx1YJJYruQh47Hxp0AZKfpoQthKgC4obR2dLrNp+o7C8YsCtdxBl1Zy
PQxiCqyYg2bleat1zjS7drZzqDd+5Dfk+r2q3neAvaxmbTGMzeaSvKDYvvBp
C/qITou+lopMbNij9ichuuJIx9+7jZpQ7OTyD3uAp2nvLzDdUN59Ut/oz4dW
6Okwx0UhBBiTXzYgZK+fptumSIhiIpem1USZcAeNkJ1crtpypX8GBerCCbC0
02frx6reABpqUCV7weaKgyICk7CweVwSuEVnsoO9Oyoy7IOG/REvUsEqC4wn
xHHFjDPZN5Mubep1AKkWAZZ/OyBSWV/wSz3TPYlObgBnof9rygX1hleHTge0
iywtRB1j0Bd1uBzhh8MxjedCeap/xuryYfT3MwOiDj5Etmk1TetrJgTAw9VR
gGE6VbA6cpzf4a5bFduI3Moye5EHZ1xwnGkWi97jvvY3ETATf+VUUZCj7/1X
VF/YlQMRwGm2LgJvj9Jm2KMatvzkP49o8OuxbCK/QlrChRug1a3N6D4/yN8J
sfaEgPmoDPoZCxYg2XM+5CYwwK/EC9XW5woDwW9DAzol6ZSBp7qASz26PaTO
5Sv7mJJ1WN22LqMRwWkPfQi0MFfphTxN6jVhdQI2vBZtDeiAqOKjl9Sr6v6a
tAqaGzme2s5UHdWZvcjfiQAb99pCLZgZbWbojHIBc14BJ5vljIlOwhOlt5Cs
qpcbgrV+Y2LbOr0QcKxc2O4kzkucVhkUjEuUGSlh0q37EgyN7/1SjLg9M6Wx
MjfPN0ISIMo4NYRF4tFsCq8ctsC0JgE/i5z7l/hJtgX7Oz8hAUHPJErGYQWy
92OTO9JZf041YfMWuuMMzMDHBSpByI0ETtrde1RYGri/yi8GKh4G6/ATi7ic
znDeQbfJlGCs+17Z7uHW+2pbb8IVIFxh5HB+pH2WyhR5v+4bBTQp+IBWE51b
Uw0unQyOwKiDo0p2YpepXJrQgd/Upk5rIEyz9C2v613tOLlNqQedITXhaijU
x9UxrZhIw9qFZmhrZOe6HbHj1w92Z1qCTJcE8dHMI17EncMxrlcvmlf5yAy7
aW8pEU7crjfCWPg2xoCcqItlz5NeFpv7jYZJ9VstP3VwZqcBcH1L7m7BxoUf
m0XDlJGqGZiE1lqI3vWXjwAu+EAjyfRNT76HsxGwdCWN/ABBUgV/oW/XMdLk
jSnMWDIPwOfgzUVYbJyvz1lRldqNVNwylnEk8ByTuvaLB3+sIb/ddzgYXub+
7aIc8PtdUgdhZlnLi7Qzgv/pES5HdS9Am9/t++KctSuCvDuec4EU5Gf+rzv1
D/7LzQfAeLEUgyNsXQiSFRhzwHN/fqvwGWJT1lqcHNizq2qPO6S736m2JVSE
7azg6y+O9sh4Gh6ZXXisocC0akGCnKbhOwOSceP9FwNYnHZRbOT0QpviVhqX
TauhPTkyd0EyrNDEen4GfaiNf5bjoJcIW63JTCaLfI0o7KJCjSVUmcq+KhWi
s2mzzk5P7eYiSIwdtleGbwhqrr3rs7kuJKyIzheBRwKFjWQfDQBDt+H68RaW
gbyY8EAa1HJXjCQPCkuw7i4gA3P440eNJXUgVqvrCxiUkXOK4cJqDP6KifTJ
dtwpVa+vlkUrwIS+9Y/aIWSLYZ+zvaq+xeNHISKZIMij6Vwc3KoCxBT5S33E
Xpk2oNOG+O80dAuUlV2xpfW7KbQ7h0Fn84krkO76tmFUO1kA7FiN6a+zJcrQ
Eri+smvOQfnq23dIPYmWASWBguzUN3pEFhlv8BCPrrv7/LjuoRz6TppulFfA
+Nz/O7iq8V1X2Lz3qR+aqXC/BtIjQ21PQ/Z2pgkmOJSqDjM8o81NzoHdR1Wh
SwzfmNTujW4iuAajlmJI4Em6nG2ypEJv1s6ni5ELhGVVzk46yQF51qbmqn0v
guShXDCA8IMcTjOp7tVuxz5yoKLqAGUIj3bo9sveE/6sU9WUbZxvBxzH5e2F
0I5SRbgLHN1CHiRC4+9GAKgiKEd7iEo5IAkVy9OZ3Gslig+7wT6NovIOwXph
7xi5MsjybGNYgxwohEqAnJvqOAh+fUVxGPumhd9AMv4IK5IB4U1qVRzVICL5
jg3dvXmUTUILwa88MGg7obWkw/y3vyM50NO6zSNgJG0F+fhiyphvhRdA7BZs
r8ZoH4rDCPlf+WIDEh6OtBar21qadvFuxOaqZjXHAavo9KTkdrhdHPVNRZbi
NvlzAFFkz8m7oMLwJ5KPWvx2KpV7Smrvk/0uMOvHytJQKD8c6yXhaNw9AbGw
uZQ2QB5RuQbkQo6TXn/GLUqIi19FqUXEqMElVEAlzKg8IGnXGLk5ININHJyZ
wuD5lbO/Tr8IipxOHABmSuAk3j1hB10r39fgTQzf1FNF9ANCjY7haLl6qPDy
ls15u+zy62Yo60l0bSMklUjeLwzI02KcJMc53u3b60nTm0Tsby09HKMbALsd
xL/eMV78M9G4GKC6TRCf1N80lL2Zlx4flZj0tY/XGuU1h7TfBanp3Efqb98e
AX2bwD0dUoyp5FRmVPEDoXpxbMX9iyG6i9e9HQ9W6Rq6eiAzuj+iGZMYB7is
2ySeCe1Zk15ZD1INirE8GD02DoMJsL1/p8wcAeBJVdaO1Xtco2yb3e1uyNU3
Dh4CCC4+VheXMj99ZzOim150pbKyGfBwv0NzmtNXhslmBJSKkeGO61a5dI5r
+gpm93GM0I5iweVaCld8PaBuY+yInyAWUCqwZINL3Fn+A023PBH0qj7O/cu5
y1h5fHP8N+fXUJhWImZUPUxzRczK26jUbW94jqJ/taUG/XXtImGBgK6y6pVP
CF2tXQRVBldzDEiTjRlsRocMUOj4sAxi5pq6a1kdduTvJpzu7M8oSzMfv7wz
AxnNMi1pgRfEJ2jGcseP/AoV9mm97CR+wBzRbHFOtOWt2cARzsBcvzydS/Un
V3eCJCfrJYVuTxWQEeNVgn8YceGxlTqEV4Z19qbj2Cgl4HG1AuK/iJ6Lb7Mi
PFd5T6X6lDqWDYVLkw0WTVD9f5Aeb4RAgqGBlP1Hcju9ww5Rp2SpNfL3N1Cc
+6ipCTbP8MqvP5hBtkQv+AeYlYe2sfx+/mPt9umo+5p8VYExlccTuwbQLQtB
B5YiOBC0k+HU+NuSSLrOc6E26jhcwLLxeKG7mM4mVgAbFBgCXcUubk2TR6Kn
1LYQTe5JZIwksd5xyA9ujHjx7KvMN7N6XOD0eybield7463/Vo6exmCAck1z
IeFtEwjmuLOKrp8x26wShGL/TC5Yc3aHsa46KeBlDi5R8ibk6H1xdkjRjS55
cpj3UxbT401Zjf6DlTJigv70PI763/DcrIZQTD7zPq5UYp7bNyPu+AxrFWxn
q2PDZtYjVvqCd+TokUCbGeN25UZtC/0RZDaHhCMlA+QEM7a2Mo34dwbgEBxq
N1SAFltn+JW1ZpxzHAR8pGLAYv2vXCGSGcrPfZrVds2LLGrtVIm7Xw0QCQc7
6ACZOE7ZSpfq+xtHn0DFLLD3W/MuN1oDIMkW0svK+p8KUCVTEHKwbpFqDm2+
D2XyUKDomiPwZrKgmlz34nZtHAe1kibLMpJbOk5iXZCsCY8zsRaUQWcw38aJ
1Yd0Dr0HJFVDWueoLbhDucO15JsbR2QFHFwYnV423FiwbeIyvhw/J2oRGU6K
k+TGUoXqSErC6eWEoJyPip2XE2JDbgWPJYwXA3Hxh4pXB/HRnpJQ+QWx8bhq
cQo2iTo2VIcHUy2sWDq+YOlq7GMJ5+XPdjr9GsdnsCUIegC2E0IAviKikroc
NIH9DqGnnwK7NiryEawm8Bm3ccPLyvWjxAwixA51L75iNi0bY6Ai9j1Ysdtc
zmLnZEOBMPvY+MjVIbtK/deES/U3LGNQnTOSYOe+9YOcYuTvHt3DFXF334JR
khTW9Z0A8m2yuiovoCZ47GOiJXj+hWarX30QvRWO9uclOj70D+nz3D8lp2N2
S5sRmC+F8pmKUPLeA4tOhLP4Vls1ReN9QdwcJhipTeDqL8fXQo+5K5c1CZzo
meRu8QG42F6wiQD+mDjcFhGUQxODNRDZAFkiCu99PV/jxz5owW4/r346M/sk
5DcN+dhXb/hCEdhyTbmC6+Z0JSYHUw2t6HetIeTw8QKc+SM16SuYhnJYhBvB
l0GiNVVWqyd8eep1pBG98YSaTPdEE8MMnTKlobuzUgF+NBYn+eQG+erLRiq7
p/cZvGIi8gg7Dc6ZiYe3FeG2kLT9I0YOxNPBpgwp/23Q2oronb6sF3x/OEdy
m66nldCMgxEtKYw0YSturdLCzhl5t8/3sxcyf1qFJ/4vU4Ub4+Men2oJei7U
0XzwQnN4d7aPIHRqDbDzLZ0iMIOh8E3lKlOj728pHWBIigrWgaMuu1IJgaz+
Zw51BfV2Cw9JR0V/pI8LK8BaqcMQt+dRSUaP1zfSBVOAU5BPiqBrr8hHxaIu
VDo1mgNgL+LtMcgcXiEw5B0cslMnbxgbNn9O96GCRx1B7lqUicTxnZYjyiYW
AhgI7IUP9JJa+2hbgAEaDIDCHDUBbd8zIVqA262iBQ6XTgGE9vuQO55jsUl1
clqhvxOanSaumXNYmu237j9w9q1DVr4owwfSi3qjEjlSls6/KivWMTug9EiY
floMZJElxQCTuHTmKOjaxD8kQUGUtna+kBOCQAeA7hOn1n+R3TeknXlyB0JK
UMR0CDPKF80m5tC5X2TOsKZrZhE4K1Mj6WeGTLinbk6gFioeSr4crQAwq9LS
3MwaTUlAumo3cjHdJrbQocoyzJGjOtJvYCX5w3C6OFGm+TMhp2bzlUKfpf30
bCrDzpV3U5cT88r+FZkUM3EhXyupelojZ/5lT0a+KafdMYW2WtSa8n6VuEJe
o4Df5FjCaAs8jR2foXdu2l/RkxBwtzxig4IpjexQO51WS3sH3cmY/eZgjGPL
Wvjl2gzN9k0GN4yEZRGg5ejuJziYKiUU0Jk61vx0+rX5Cag64g3+beFABo0n
3/c3BjcRHMGYK4AII/o39S/EjfBS4mMdnPlj55g4Hk1X+adVAaQaEGl6lmuN
iZqTuk94IciIHCa7ZEL9Sz2Y89kSKg65e8pYTMXPZRsQYXBe8olOaJk99rWl
wQLaCfwBU4tSROgtYdWl0D+rEHzZmxE96PtEj6PVMxwCgRA5wfEGNNkxprG6
amnXYwEyE81GTsYNsXuGXg38Jr/4Qy1EJu8arRciEI35wn8b0NEfS3Xtke2P
WiZEH4Eceh1gLibnc2LEbeqwcsQHDb1t9q8WWqRrsnMOaml2zxlDhIIGCPs1
Ond9SpDlRdVUjASqg90/BwuqUTrUyyWB+hhdFU4oKAx90mn0J2O4+jm+Gutq
T6mPjFOQfDbQ247JHqhV8aP0v6JehS91I66GDxU2kwghxgeKBlkxyEAucE4P
HZ53ADgmBrOm7q+CpQ6GbgGrhaI8chgNSdCTUrs7bdeZfBlSGh3SHjUN0hqI
5Cqh8vIYkUW+eY3HsW29A3HPGSz76TK0GfFawjptqFMmDVnyFd1ErqgqThtt
0z5rkrRStOcPTQxReOtv1jiLlKe4bNe+TMCGtUKvVrHgvEaDLalhXCitG+EX
d1zVm0w/wglPQCRRQMMYN0VMQqLlqUcB4xYhB+36JjUxBi9O+fAcnh6alDoN
1GmIE4FOs4hf679k6qB8Vs76AFAEFfQYwhvzb0k2m6DEk+6oMYx7khOdi+HM
Lr2isoo+MAfUrBw5/IBIUoF8RSj9Fn17hd9Bs/iepNHFeww4po0o+XRgAdMy
WFzLbuK2+/2LTT7D3Uoz50p+SorL86z/yD7+BFGmWiqdlZ3TwnzFGYFpX80J
oPi0UVJTtSS6gpluz2JRk/XMYJLOhx+5m7+/KJR2Twnw3DYFl+c/cTheWztR
VPNeWop0KelWN/qvaLqiD4fyVHPDXwWZrVTPSAVp+6pGp213YxmfDz1cO3yo
O/Nf6JNBums7rK9dw2StBTm2le+XvDmqKv2Rd5D4/fWJ4bFpHHzdlxuXILM/
aok4c0NrPtlE+kSg5/l4B9pVd1+pzbz3AXNpcR2XMP9EYEcQLotKJP4UNZop
8Q510OdMpPsSL7tmMzMgHcrP+BoJpyvHR3UKKDuflj3LokGR8TIgDGtnmmAY
zOHbhysolCvg0HET/UbHB46ka7tFPWQhtdAxwq590gHhSeQ0kMgpAojrW1kk
x9t8CCgaG086xZgdYy0zNxOMnqPmsXzz3pGWwYkQhuAFoytfZW9NbFAtXc2A
F59YKUWe/F2IDfXXdcSOYAuN4UH3IFBu/KKs71qNOBW8pgRV0l8tYsNxhyjz
M2te/GFZkQ+zxkZOSI2Vh8yqq7biTa175Pl8kJEGnLockVQ1qPvVaXdYjbhD
PFS6haJpekImpbrVesOxUUaq23EVhAZAEURQXzgTOfvd5j7fka9bqQde322P
nqiRkY+AIAvoKxSMhBetosTxOt65mH4dvUVJZow7RjpBFy2jUchTNnUKSmb/
4Hbxf0IXT8usQrO7MRwKRRnpLqDKebwEnkQuS1gFcFhT01zg4/E8taAFTfdI
KXkYYVRSVa9oeNPJfewbqA+V2QepGNa2it1l87yAvwwuHhU8RVDX16c7t7cB
scw14dFjoSDlJ9kjDOnCwdMdq2sOoiOy3MEqcbJA4SPV+7wbJ30U9fYL6ZFO
q6s6FCLqtzi3/NrIIW71B5pM1yuH0v3bW6FNe4QZA+cp1VsRNqY3jOpHcnDd
arMKY6N81z07NGRX2DZqIc2uKxntVKYoUtFRqZzcj/J0VtUGuMiCA238gNeG
u8WsC0nTMBGut5trAwlH/CWFDIuSGbauQi3rHNpkEFJLmQF55vrRl5bRDXdj
0foiNI/OgUG5+/RX+sAwXNzbwmZZpc/+SNcbM+S/EAPDA91lZSQcunhHqVT0
KBBCxJuG/tBA1XdkJv6WL8aIdKfyXAO0HiJCCdtw+h9aQjykyXI8vqEWYh+i
E8bKUn9ZKU0pnrmcH/gjXy6yAuw0NFqVrSOJhsGNOhvn7E51aJFgEzjA5+5N
YgbOP4SInPIEFE9Ns/79MbO69pDv9A1rjYEBuGUulO7KaSf7/SiBmC4QaZz7
iyC7dQ9FyrIm50GrkwHYgzZSgqNSFj8+tX9jDu+ug87moCWKrrTAOwiZZuKw
cwxTmC+16Jxp78lI0f9W4MRsmxMU3H684QgW9YK4se9kRJgRf8AvlVYIX9LO
ZhINfigxB7TCLpM3j5idvDCDyYP/BQEeaoQAJy0k5yEMyFyuM8vU1AAfxB+f
YFo/NIkewGO0vyQyW2FKrg4cEVftAIQVvXq99lIH6vvcutuebSIS18bTdMwo
nZVLTC/rSfLJGi7xpnkGGvUlZCEQmaG9ASZLsk8lkl57hfw1bgp3BicKR7Uu
UOazUUxS93sO0FJf2NU+2JRJdSQFcqJ8DEYIFmNy3DTuYYQHBQs2MfycJIj7
58PJKf0PaX6Mae+bgsBxM0id54UzOM0pHmukhFbA5pRK77bLWP2jwMWzpV77
9e3INPAkf4bpYs3GEYl4zvT1vKAu01zK5YbNfE5bWtjhQd1vGtkLf0IZ/k6h
kMR/kkOmj8vy0E9sgMnaPQZRtn/43GH8o6kR0FgOAGRER/pFaWkQMW2tkOqU
biV/yUkyz7jfGUWJfNF+kRBxSXVvghzWQN0P5eqGepKsD5ClbrDdlzRG2sK1
f0IyZeVlsqdEJO0JRBaifkT9hDKZ78UmbTWXgrIfuPSnFrGMvsmdEcL6QyI/
lUuGYjdEL+3qVYx9TA03qNQsRFICb56MKKuY3+hY4+/LlSQd7pT23ixTtzut
iieq9h7yZ5k5WimF9waIsznbzkVvG2zP85bB6xUiX22JQiRPBwrZht4vCo5k
8TIgmWekTkCXuxFmvxNQxhAnlQJ3Lg7mShlnh9GEyndfQ4EtRAaQ2z3uNAeL
vwJUf3aX+StdQ+HyNZEtqjEFMc6cIqAaiAhk0C8RWEKebE9blHViRLaYzDbx
CsNxKGj774kkNWFXNK6QgeF2mJ7CRN6UAP4hu0nrlCQeoe8sFvhE3oMsA40E
ZXZvKV9DIQfTzu95m8i9R2iuI48PtfoX08nyeiYQxxNeLYmZ/WpBXqSCLBdf
paafB5RR1FLbmSYPLJCQdA+jDgSFiVNS76SFvD4yfOCVhljajdboLo27n3nY
xM87Ueuiv2n8q3VFlzpaF3RugZ+AzI5ophJLWRBJ/P5grCTHS3vfGAwadTyC
B1gMT9RYBeep7oBrHj8Hof0yw+t2c/sljfmkbecnBKmmnPufibD/1q8b4NZQ
ansGYL/+F53gslbtzHQGrTWqrFkr930au1oKnKJcPEyP6VRMtCg9CS4b3/9p
xB1yWLINWW+adht/70V8R+LVSqGpI4rrc9wmFXMPTKXQEG3lrbCmOwP8lcdo
7AwMeM0faJ/gYMZP6DAIYbpaeVNAta5rL/+gWCt7t1J46GSCf0EcSSoaox0p
ObAjsn7BBDbT91vRkOpdMKSgju2Q8+wF0QxxmULe3vn6zzS9egY+la30ZcCH
4gUIUeFsiuICsAOwjJ8pZ7q5uCXSzfNQFIdHMPnPuSi2ykM74GZaMjbaF9MK
UM9sWKkxvLQnAhPZ7T2fe+o6/1MaywGwX8OI8ZmmEzt/T1DXYcAW/dI2fN9p
XsmXqBxIERh5/C48nHtzYqDl5r1FsRIsbOmsSAkKPJDylXTJoKb5ipTuy9KK
9khCpijLEcyV/4Np9jXnRdcxk1jvDvtMpnykoKs/uMswR7WRz3C+VwSvn1kY
N8kYDTatQvzAPffYYl6UzHvCGrKITWI9DoWZcNQvmOrOH94CCA5XzQ8cfLEF
zdl4exao+WXXYwh+VctFvXFV9N/z9EmEIvxgjTZGAxtSYIMLWaRFnFgp962I
yoPjhhhWwBEw64SjLSqGZWQlZwbDU/nGBSDYgbEXnj76ERwA5F8cpMC3gdgw
5KQkyu7DboHysAaBRlvQiAJKZyV9gi0ZIPYzHca5cB8kK6Bu3eoNFATVo8TU
R8ERP4EBZ5OjMuhhLix2/lQCXsN0XUol9GCmrHoACZ/KqzJpSAGH0m8hITZB
FINXnA2Vd3l9ffULnlzZQ4EPMGmc994n77NKoBOm7TyIDwnz8LisRq93C323
bxq/Kvf9/C/Og/KhLDsonCpGgrDqgwX6kQO8+tu2ouwCAQ00qoV5eClpU3og
RhwSCOk/Rhp26T9gCWf/BkOWeyfaiTao5tAkYodvz8S64oSVbcAdDqY6r3pj
u2rXBGtOh8SIbFtpJTL1dypmBJnE+PSMN+zOFlByyTfgLDpx32BsgW+Y0+xW
D9QT553x7jaNdZ5JehkQe8s4+KWtoI35aXUeFp6r1OxRs7qywrC7xP95mOBc
8UozFCEbrxhuYZGMa/CscQy1TDRiWf6QjvhqvUF4Fk6X/bttr0gZ4d8ggkyd
Gz6Xvdfof4feL+a/KWN4Ib2hvj2m4LXu7UmmfQBXyMw6ZtXInN19pKMZsMZp
vky/wmcQTC4Xav/vJZBtQGTbgmxj87mv7VZeCoo5/CrTpEVqIHomssndG1wd
rvjuHwTvOqcZWBV1oZD21otFPBpysLzAtzEjhElNtsFa3mSViZpnIjACw8CA
hY+WdwGmQpagNc1slIfSthbu5J37R/NunyLf9CJyrD1U+D8YdERm6279WYeX
kHbkAjM4acxbO3L5Rq5+xNPXZfSmgbPAodM1WY3cCc/nK8/TDNfhHZk9/04X
mSOUynJzrYAWfezf3JRkY+gYkyCc4Py8Ndchg2UEz13kdrAI8kmW2jOFDonh
yQuUjOKzNoR95x/xRe1qhhQsuBMYgaNWZVp3WpaAD+m5nTu13rCp7HX0Hih9
q9LCYz7+85JT1x58HUZMjS9PnUl9G2RM5Oow1zxHyPTOXbC+ZpC3JFVGcr0L
w/tCB7rh9n6lViKptxAy048qfZR0eDR96lSGa9gjpIqGPyPIhMeQ0KONSLlQ
bk4a2ePui4iornPo+fTtyrnYeM9RJAzr2xy8PTgHRt2pVP17F4oB4m1kGMFJ
R+zF4TJR/wYlnsLLNJ+zkAnSDpcxvmWO/3I2IgW7qazT2qCURf0mQjQt70xB
nt5eGR3eyvH8flLMnMLnDfPdn7nrxCLOL4OXb1cu8AsLDM3f7FtP/UqzirAf
hcslWNi0PNHwGwsLIrJOx1DHujbt/E4RKUBiaFH3T4fi+G6JpudpFamHO/CB
aKe1pjp7Ufh/JER83H5ed7PiSgzOV1XCyUSptNBxzBgyTQNcVxJ0F/Qa6Lt6
EOPI48eXSMQT4xQlT1VuoXNqPclSxwRa8G9Nsykb+90LnBXCwpZ4fpVD7GP2
kl+wDDVxcYkY+x1wgKDx3k+OOrC+ivO63BEK7GwQGgiZ8jmsaab+79whnYtu
5vgtJP8YtpBKso20wAIFLW/vMjnUUsL4YuFZKvY7E6bBHBxko/WpzeBYvJeD
WfxDwPd2hUxWYOwrFB1AvIPOnlBXPrl7iHssrmS2V2wh6WfJkRoi9GSrq6dC
0qv+DiDO0Yz5puG8zj4r46EGLn0i+XbY1zGGc9ncY8Q4ihig+Kr/1cuv4ZsG
aC/jh2Sh28nOn4xUToZGjzGrbOrU+5Er/StzlSFm0mcvq6hZXT/vF1NAZomA
ukv95mx8IUqlodNWjVLH7rC1z7rXOS2MxtCi0FB6WmGaaokEJgRrZKBt7zIk
eP2vG1hFPuZcRO02IBvYdgCg6AO9FGrHzmghiQLcT3ecPjTu1RcZwAwnl8O1
2P3IqPtAZvQcsQwgDh4KGgcOhoL05n8VuiTsrQ0l5KicJYTXK+47U0dapBLf
lnpA46a3D3E/VUwHOOQr3PBTp0Qq0WFHp9TWI/fqisJwDXF29z73SJoC5OZO
5SfCTxBnxNlCBSdqMW4R8ZWSy3wmggaXterYIraL2gYnYTbWQCSisTCPP7gp
I5yPFekVQWviepLGFl5Dx91OfDVCEFouhisDuxZYr4ysLeF53Bv3QdBEKNpo
+x1uJHY05KVj27m5pqe7ODscaAJEvq+20vDZS08QMoFKqQg+8f9+Y9co35ZJ
GqL0Sevtaz+gvpQ1WgZSBnojbHqdc4xE3U7fAe6CH6nbIjJ0WgfWYUEJgRoM
zlZsDVO6M5y/m5Wv1swChkXqZNIJKwBwidC0Eg5pXHL2mB1Z20zlq7VK0OLc
UeDjp+9iG7ADNhvzmEpjNPzfLjnjn9cgnPwUZHMZv5HtwEa5a6f2R2lSubx+
Rh3IWqR/V88bJqnYXo+EaaHmNqH2OV8yQVhXL6mbxX90FC1PUut/q6B9ad9M
1yeOsaRDdqdiOVGKw62SpYbyfHI7jsWshJDNOrye3Zy/kURRPznZdrbpjoJn
s8RqtuSCKMBr356fwm5BRYPaCsHt2hvqQuT1OHg7IRzCFU6xDwWU0YrKlGip
UNlXrysDEDdMEt1isNry8MLskPqGUvWJ6QLq2EZChz8OkRkl8HMqCDT0nE9a
Jz198oGENXJ1+bbASu2aZVX3h61U3mWqZ6y/9BmXmAtGE3I49rI1lyF1SHbQ
mm86RKGXHLHw8KLlYuy4dHYM0fIrOcNtfuDwFhktNqKYlZChiG986Fhu8Xfy
5Uz274qS09lUdb6bFD+2egf9xp2yXQpf/9WMUHDjGkXDlFHnbDvbuvyM4Wpp
laKddXDuXQDuFflbGAbH3QhQ5QEfRhCYbrIL3Hj6xq7kUpaUJMe6XBMmTaDl
KAcQR457PZHK5swnEKadeaHKX4HlAokx05dZ6hS7elrDhyTjqAJBaFZakwPR
FPVX9H586EWGuFjjqDlo2KxxLY28wxk0igSqLH8aHZFBgsmLgnCFLLx7PxE8
yZbuwS39PpwmaSwcFhf4c5KbPAqZq3B5GDu8CHh+8KV5RgJTVGMyJ6HDODV/
LzdC0TuPgErbC2sx+ZVGOwzdKn8Sn+4uaOD6+LVhc9E5d4B64XIbHsDSRk8j
ZDQNv4HsKP0dK1qdELVV6KB1Q7LEkkOZP2+tUVkMufJQS/baWzjNy9fqLOGC
O4A/NADf7iFGRdu9yhM/0OS+dJIGLrBEtk4XRRYY579OyNm7fq4VA4fMt2cR
vaEOa6cK7Yt/9Sjy4SbQShJMzScI6soDjRdZRyheMmrQ8GSjUkkcDQYW0i/N
1At3uBmDHoavWHn++ExMVAou6NysdGTRxvrD1SAL8MpjkhUs+uUPg+MyBMK3
GQw//SYiYLgKs2/lRM0hY+Dhwgqsz1fEygm+OgT53tyAw+IL28nyErFfyjBk
3FEE+DNvggMYL1ye1PRFqjAac/+je5V27o8L1za0+VKtDp46GvDLF/SrQ53f
9Q2E4HXvK+GlrTlVX0vmfFpg/ikWgk1VYoqlaPokdowqFsdljNtsdsTFD85O
tAyfPf2Q/6ZX50g7O6KuR/DSdTkaDgNfaeKJHSnH4NEiSStifMZrSnrLtJzA
3iVpXCUMf53/GmSnoWNK/TG3dPX5BGdytnNXzHyd6yCzLW/hCDM0BFY6x5v5
pQuEDYm3UIe0E3b44DM0kjQpJpSSSC+7Uy0oSI84xpBuMPtXlq/j8WnXcFOY
RpuHRqUNQQfSstwMfwzLpTFfjNCh+v1AX/8sAzVK6KrzLFSnscfViV4IiDQw
jzuJIZj8l4y45LN5/f57LdQxBOe8SZRs8DkVvhsGB81VQmgNPezPbGXdK61A
fdaGYbs8DfZuEkskfEUcphEA4mi4hDySSL2/toeG5Ll8ncGfKvkr9ndj27xX
r6YWkP7idPc5DE8Cj/xbjDJqYPjJjspsn7OpfI1YXe+CjKBXPW1J0czqgEQ/
jI982Eqiv2IkKjc9qEUv0MeNkLpEHe3JazEPO/birKIVMi3caUojkMhI9gNZ
X2MpGNIOq42GV5T4K2SO1zpUpaLTXBRbJ/9mi+cHK2kDpAT7FwPTnNYoCyIZ
SEdfy264++lLY+SAmd8zl8ZcIt3wgwRD0yOvfNEOCMvadVLoHnkJSuxARz8E
8bBQluyDp0GAohkbYaW9G8weMqn0Up6rFB2tI5MaSH+XlQ/x5Rk7VvM2mwG/
46GMvGwWSKrxQYBydlAHwVB2E4aB6Vh/Vs5bjDVaSODvLT4Vu15Quj05xOZd
oyuLWw07SbGPTPliyGeUodNXmQA7V24kark+GHhprGL34VFDmtpKjDm0Q3Kt
SmhwDoYe1kP9zi0T1hOILGrhmwaQ/3dTt96uyqsLUx6Ls7lI6lNBboJ7cMMu
KdLXAFuxROCUcgVDVzChvOvBcF+0PcVdfn7U+WZqjhryWfFmhYd2oUJMzv8f
Q4R5kW6zvmMacBROvquSICisGO7LpC3vTSdb4YAcTJVzB1zfbu+9xrXBNqy2
v6I24kjLRK1LQQpV8Ws+omCLBvdng8ypwztZkVa361uUyms9jejGxjmG1Oqy
rhQ4CugACJ31PW0wgatS53WHczrdVd1JZHq/DUEXJNa0WT+AGG4QvfjLWn21
4zVx8as34mSQ3nOFYp0INBYn6Pm3jr9nKlSy5wFqByZC3z0KFrJU4Eiz1Dzq
j9+U3OyWmlPHfO8EnJxUTjayg75Uh+MQsG5758zriRPZuRqxz+SVRp7txSgG
U8e32H97bhoCnE9T7PHjKgMNgCKAq9z0uj1PlkUlgTmn79Oj6fb7a4j/xIPw
Pq7ynbio2qlIPJlx9YnfLGwcy75+vA403dBsVxBfzFnUPEKnOwlYnmbGStLE
uBljyYu/lrXgQgVQOuPKNcPpm024go1mJeKXLG/XaEicwEgmZD8vhD0fOoG4
0f+oG1vyrYfLgMqlWba1AMCuDkacEq1b7NBXMf3LfFxEbszaAlkMO+J49xbc
cEU2qFcVf6vz+O0pWzjR9Kd101bhT6xNDArScFK/B/3gdnUEGMFEl4ym8tms
LGkHq5ZK4CPdIOEBblcnV6RLoqVWQHA+XDsDVyivFTRrlrNwNys6AXpTXYqN
N9OOj+nABaIwjkuFvn5J9fIsSThcxIjbaG7oahJklFKomci1LTrKmR/LQoHf
LJl8YAopRicfH69sJo6o72Ek/m/wF7/ICN2P0FV3U7l0EWZnL0HOu9lXsLwn
JOMcH4ckzixH/ksJvF9o+MLR8NypoQdI+E3q848bs/T047CIz5bKFHXqYf6X
67PpbzsmtkRBPspqwWZiZybsj2b5R24Uzm8oecELYOjIl35duIVWkMtjZjIz
+tq7tqn31f0ek2rMsLIDp9O+jfVoyRqCX6o9Z3bob/5doNaPHRs9UGr1s93A
hQU5G8ijSZYjdMqwLH7bG+MHWesBRHXqC/XQdRWak4OF/GE1q6nc8wLeIIFJ
4Md0wlrIbte9wcOT367qDTCCZ9UChp3xYTEnWvcz0Z9a/XM3WJGmpiYNaUP5
iaMVEJIjGSR/h6ceGBLuZ/O0pLEkZ5euqd3VBMRkNYeUexZrsRye5vsWtPXd
Pu3L3W+yanWr5pUjQEIg4bT2ZXfc8maJVT/oGcJIzrI1KxGXXxhGM+uRvIZW
p1RzdPMDyqviVkPMMxuoIlqrX/hvmGLUiYsMhLgXG8vCsxMXNTvKQ01Svtlx
u9jCxqK+GNqdPxhtM5JSIVHI0CmO1CeRoit8gB0PgGp+gVDMUlZS/lno1eKG
l0vHNzrJUVzkDtq8P3ZEOqy7YXqNJaYjSTL0zhbjui7zb8FuGfodjw88BLXT
2E1PwK0SBPYL1P/3Intdlf+37OTUK8u0pbAHkWicY8/W9BtA/8IEZQqs0NQm
rdMREtVkHZFB94x7OHkqFXYcK2Cm3S60SYnRjx2BKFWPExgDPTQdN1h6w8nb
czlNHecNMPjrUZHlNBpryjy1fyS2nXv9Q/UyI2CS+nwuZa6ofDHeKwdHjGPP
tydyyOMIRjbxK6bf1ZyD1qe86eROXIf7h7T5j3V6gA2KUsHvXSQGNipT3sQt
4xFH7TeECSL43V4xloTWfLHh6zkQhcZTGqFemVkEJ4Q43lqvNoQ5kkdpN2cQ
kddFch33YDByW3BXHRokZQO8621ylXPewvG+8xeAYKFy9xpViUdrquoTmVrU
YE9w4V8CDeNzBu07Jue2Xe7JJkCO9bYrd7gutKlnr//8F7pdgv4pqq5nyANx
/QENZOChP+xGlVR4WF/wecWBDCfqgYk2l4TuKxi5jIhcReGUHXBhguLDXhts
qc+W4uupuMy+PteY1OiDUDHt7ykL3D5nba9E/CjWcju8Wob96EkM18h/Nvx7
Izm0m/aI67IiI64X2zJho5YmvfH4W/liAgGcYBO7y0bug8G+zc4vDRaFUwqy
xkJaTeN6nmYgnQ9wcQJAeVdrIA7rEYVt+K/3lYK1pCDBKMhwQlMIhLLbOwNr
okbB3lpsLpXYRWSU+bZRbMApCb2R9+Ng9S8qfa81H19jV+GdMKpKrSfpdAfE
JSuiuJx/0ZNESPSgMLJxrWXEN4cFHiR5EPUFGLaG+p3gSFrVwE/T9ddr7v2w
wktZpL7tcWC+SzGHK6OPii4NAnnlw1dY5qyfigX8n9qTmFsiEx22HAgWHsnc
1zGljfQMyUV5nHa//lqtfq1PgSHtupojAeiTr4TkPSANhAmtMwTdqBeKyHIp
EO0JAYwv7w8dMmjW3qbxYd+n5X4rxtkBKJVEJ7LOo7Zcy7og3nucnbpO+0Ss
TxO8YV2IBKP7bVxjvyZw4atKrbd6/TzGz9qAb0YuTm97VI3BvKtOn/JuUS1d
t2hov+YIKBqTsuj7+EhyyT05HYvaTUvEUwmt93od8TP5WkY3/suVF7hktVLF
Tqk139ehsFcwl+QHmQoiwqRGIwwW8BVPepR5So770IhAOZrn+q2sEM6CY3Dk
IomPPZzmot2BqRPbSe7e1uq72dwpIJqYtLN1oaEEeqBhG8MTCiM01OSADF0y
kh9QbVADo4Fi4hi3Pwd4Wmb5E6SJI6X1Hh4f8YfQEEc7QcZM5mrVz0u9z+UV
QYrW2rL0OGwl+On/4DKpKTWsUsWKNM0B9b4Zpq0lcKvHttqyjkAyRnjmPNRm
EMIU5jhYA77jmtxxx6HQR9MSljUU+TgLlcnB1YiQLjzA3EXnGGbQZMZcPDsV
IwaNDSJIocmoLO06v9lb7Q5QjUM2SaEjzkAvXf2ZVPwomEtuzbN7ZbTFY6Ry
GZL2Bs6IlkNHIFiiF4PfJIXgsQn26+EKSMDYfh4JMJ6u6rtgVg0wb19EIPlv
LPpkyDRcpN9PvPfaJvojyXTosGXxxdjK9UD35ukjtX74Q3KFOKhCAgR45jiQ
NiGCx6/ZR1A45EXUBg5HJh9oWNWDxmLsdA9DmjgA/mZTHuupsmSlNDXahkLH
spTxt5uy3po2O/pz/8w518GnvhKSazSsPIVj+VVZJfny8RFnfr2fmtwTG2tK
zqeQC8gz9mGn8m3yIMH6IaOVWLTOMqR2Sj50A5Rh1DGjzOIL67oE2UaPjUtT
QnpyrA/VorZkS5TCqT9uhW/kzPjXz6SFJeFSNtMBDbMQOOdyNRkjwScK2C7A
58Yi9JfIdya+a8WF6Hp1dzQnhCRVJykcbHrJX2ziP9TgR016NVSfMvjSKBnF
hAZC+4Bi3NbDKe34nZWjOXidc628XXGLsUyUwew+qY+AmKxTSgAxkNxzRJKC
8M2g+mwUb2izpve4bZ914z+bQ2Rw7hzU4lE6xxSrcfYyrLXXNVFYmeKs2dA5
Wx7EZJPWh7PZWv7HhH9lhFE+TB2/oFf6ICAQgrND5wkQJElqHCj3+fStegcR
vljdcdTwLy/kFZwkRKwDQxAGaqmPCXNnIbNKGkZqbqB7UQZZYnCn5mMqPRcH
/kG0ByUPiqI9nMDfRAObTHnisEItqxiDwEu0w3WWrWNafO0CdNpNxYlayHYw
ZvWVmZDRXApf+fPquIiWD1gQizkkKNVd0UBs3H+sjMCcJlpAQwspHGElT4vx
rkpyRhC59ZtMv7Yk+0ImkvJbHxnTaCgYLudiS/cxbTympfEA+nAiP5zJcuya
6rxgtYCF5XOnMjIzPkPCtrLj9StyS6u/w2lNV/vNNqyNf8XsiT/q4kjdGdnq
sKxH98eSX0mTpqO4EGqp1XiDJApPW70bYdK3qZzA4PPZCRi8gaYa/cqrfutb
SrIG7KJN748GhRcPHSNczJ/enms6LmQEuAVMVntH+r04kDaoT1spCnAKqFxh
eMe9S/L8ma5q/u9RLMoal3ubVQJExRdRTyO8VYp+npjtdbgcfSrcggIRvRmg
BGqPvemJsfumQdWotUplFBnIcx+Lx5Xc9aI8ozT7hw0T502V2WUudQOyX2C1
B659VBDeBkyYOP74jQjFHlSKM38xpHa5OGa5OxeCA5ucJ+rnle5CgpNPz1EE
qJ1mUHk72gRk9lCTFIXGIQIgsYlRZspU0JXiFXpXTjl3J9lZ2M4z+cv11Gp/
4Tpgrwne9WHlViO2rjrEkGl21qO48KC7NVfJC0p6QaphKIusicwQ22QLTguv
nQDI8AVouN2FymiYD6CGP055APvY07ezxKOZ205zVne/bjGQ8Ifd5vqNaMRy
6EQcIfQVC10XoPSjcdjHEa9dMxfqs31XwpNYv8yTjZwMbnzcIuiapVupVsCP
IF0yT+QGaQ4JuWcC8EcyXKAnPAXyx0gkFf23/UQHiXC1swrw8mKuFpJLXFlC
wr5D93YsTYG2xUb8SMpjicWbowMvDDh+bdAtqrTpnO9uhuGZXMuMEWBm97JG
+pJLWNr2AY0thUeS9gXkkq1gIIxIFnKQrSryMlLRZXnCEtL4RcdwHs1NdEA3
MtfaDSE0zd6WY6VXmCk35CdjZZ0C+EA9ShLSZb8gRB385V4ATxMnDFzsOBue
8LBhj9pbhHSx8xaSaOqP83jsfIummGTu8fh18TNKNKq7b3iEjYMaXdc7oivw
xcx55zTuB1kTPVXKlpggANUAdeW6fzMr17RJ6h71ahFHRQM/ysRupsh8kGts
GFYZlcPHsixh+yoa0OLtPahfb+G1FTtCDdJg/QTv0vBqFYruT99Ey2bmVeQ7
C6kJYYAHJtj+zpolJdZA4Lr6x/XfSlsFKuDaIB4YXpILJk/yDc4Wd8t7/Isu
aYGj6nbpWbqq2U0S2wWQkYenRn7IBQRbHc7vc5RXHGlj9uRSuEKTZjnklLeo
/AxHEOZHpATd0eWMd47LdJu9e47bJyRMnKuALoV1Wud9/CIW4j4SnWBVqVGk
TGa/Kc1pow0zRxjgEJ4qcGSLH/BZ/9wxlh4ul/5RgMQW5hxbqDwoVjqWiZNI
C9vGqPjhERkFQrf5w1IuL0afU7ucqRyNvZS7hBZEmruHEmqZs0A6RV+i3V0m
cXNSABuTz3+I5KO1yroocnBBF+6oUqVhAR0WuHGPsBpl8UL+Kth0fVgNNLjj
4GwBaUiTIJ2pVGu97MfS6hgSrFDgleD924bK6wPLysiVH7hDACHoM3aAqGB0
n3Zietz43ceTo9/V4vVxwCW6GgGwOH2ninKYlA3aDocSayY5F7wYNExoow4v
gRUTGi2yZVsHSCp6Zh3axyDm4YHO0Erl6gpdZ9lmUdHTRb/t+93QXbh09ndD
m9vPu/XKWuGojwoT0Wu2cLacd8qI6emZer42f0kkKh4buUVbv4ASN0oNXIqi
1Inj6+EBkyEK6QD65Bba+qZxoTRs35nYol/RZWQ8qwERFxus1mHiu+u0oJ3f
u0MHnsZqvBLBXOA/y9ik6cKrXd00QGAzeRwoF+x4MEafsKL75S44YFoOZ98Z
IBWUr5M0hJLlU3OYtQNpZyuzwgwwyT870qZs84jlMOq3bTFy37Ck/nWzwlu7
Sjaq/1KjbzCvHjHRjaW2+V0ZNiVoUB4QpIHBdmiK8IR6d4o8Bp/shKGMIUmm
GSKBq8Jau8s0TgGXMPnqPiV1efuHOm6tjAs1pK9FX6LwYnUBlcdBasOqFrHn
o6wnE5Es1tGAxK7UowwvjLu3/h4ifHoAEZBqSCvv/D2rl9Hz+Q/QciHhRF2S
OaKtxlzcMoWahQ1+ALVebHmvOLLY7bp/Xc5sNarE4VN8VfEV+np5LrUWsCfQ
jA3IAxrVrC9UENkJ7PMOgbhIIyzc+14yI2B+rHIuiz62Avm37E26NNC5BUnO
QQ6LhHgUUEaBtWrKy8/kqwOmkpuZFokD1u8/3F5W4decfC+bVmmiG9SIwl7h
PkzcpodynQayBFFFJtydhaddeyS5Z++ua6q24qkRdaPhxItHJEoga9nTmq9e
JMf7Xj7b8HLqGTRgRySVgvzrYHcjKUtgxsU34JDNlXTrx4RbHxoUEPDgk75e
gIsMSOkGGdFznygl5/QEDDFfem7UufL9OXnYA5rn2JECdXpLv3ceRycqItMO
OPOduGaHrAp99avl7WwEemQCl/gBhjuP95HAHZbbQNIkmy2Y8eFjtu/V0GXl
OBVUYWZer1wtIAmu08oY6JjPMau6GlbjxW9phfnn1wimftelE7+pL3Nys8ws
2SDwqzDop7WNI0t0bXpknRQM51GVKLIoR58oN96l4dysV6j5dhgjb4EippBJ
q+7qfTqM+J2+tv7E8Qn9w41ZGG9aKOjyNQTMOPqCrKeRgh8k21H8Fo1fc8/O
n/3y/kdbpPgxxiJwNdhKghbzkv5KguZSgB+P0RHdp2UKID2icCmkAUWF7fIP
3ZogD8woxPtnO2LD8BGOI0Joj+5R1EQpdGGh0bm2EFXC5AJ2wRIREB2z26gN
sg808BptReuTC+vfs+6qo7Z9xEvO1wTAHSHp++CH2Jp8PMLPxVr7cmc02aVO
l6eEmGYbDivEGj7PW53jBITdf4Ec0PQr0YAtIi9t0YFyxD4+s1dQ5UXLIIvw
KDPmcKRfQnb7JKyL4PWHOp8Q19QgTTY0BoIwdxqZYWVfImYlCa00iSvlMb1V
E+OTKxOdJvBVVAK60vjxBiuPbAWTdTDgjOmaCdIR595LYCf746eBWwrvOJbB
AfuU2mF5LeBauraYyG0/JWDso1bRaqfb5S47dcyI03/4WVLOMX9NYqn8Rz4+
cF6n/BeiUYIGXBQTUqI/R2VRI1qlsivng6o18Hzld2IOeQ85cOD3SjGOsgm2
v8QYOeIs31jhoqtsQmWdHxsvRE4euMf7B8s4fmitj4HigfEa/456uQHU5mXH
WaQY4EI5k/lUk+2raCtcrWBQYaoAXnhCo2jO5bESMPyzMCbf9HSYG+gfKJ3J
rWC7T69GSA8ZPimN68JKXjLU5HrQ8+DhzqNq9q/h5l4WpApmWZhgosAzKiDd
s6lzCeYqDBbUs88o9w5UzwyPysV0DnntRXX6W4oxTLrIM5nvP8ux9q1SaZD+
tq34IXghQr7p0GWxZrfCDT0B/NXaAMXlIgW9AXAwhavhzg6PsW/lfSOdcmrf
hXAjDoHRvwplBoY/hFUYeqbHlarJkoUBtR9U7ZdWkI/3cKTpYPl4+TEPsrmC
dkFRmBWTdFxgAXpchi7PKEfrpEv3+EnCW/YYfd/akP86W+lFhBDd9yi2cr7R
spvnxLAZXtqHQ4zaFA07F1e2qj4mXcYjGxrzZSErfOAJ/I3K8c9uH40o5UT4
rzT2w4DobIi63BHcI/nll/FtZJQlotJPiWBZr5P9mSXYjAsHbmEH18LiBY+X
Hcvs6vz/fzpXcpPpAzENU7Ccc5vzmCkkkN+3ZKvb7FyU/9uHwIhUZt7JK9W0
nT+0LOt3f+ZFoyLTQp5xLtHa9/yZ1xnEHeHAWMSCHnpGklT8Rfo79thz/a1N
0jrCKwlAG0zevVxJ1v9wXmaM+jDRqxj/vJO0jMV0EFjxeomURE9gE9gdZtaY
9EI+nRLkv4t1MOrV4GM9A3IzsTZjF/nbmwdieLb/e6BIsmXRffpy58dJW0Bf
3MVr9v3LmNihyI4mckE1BW4fH42AHUhBCMFJZXLZM8SNzv0yX487Wf67IydO
mMNwP6r0O6IuXSWX5dDo8DEK2t9Hin7rIkM4+8JCs6G2y4RNkONzuTFR8kUQ
/nCg7zNG2WRjdwv2EkraQ7BEreOAbiE15gHoNDchJXcxmsgryVsC2T5YjZ2S
Eb/UECWN9CWwg2RQpCFk+o8NM9C6+VMRBbApqC1/HJhMk1fuIYo1j/Lnsz/z
zwLQ3tNUgON9Kcf5jxg6BqN2sj8gm3rqDOaKsCVyIMQyQ1xtrUotYL1igfbd
+XxViFdxcy+PsrCFVJJikBIydecTDu6SKpDtnf2ezbkvXM2zynBMSJhLynxo
AZX+4NOWHW6rCXeInyoiAXo71mC7GtEUvCAUACWbp0MGAcsgNPZ4SC6hj3A4
e1EyN5buWraRYuSVmIWtg/0o0NpMNez7kVtY7qfBy/Hx4db6ipfZS3hDeONk
Tdezxql2CXgY8tu9AmomeYm+l86oomeokLhE3Mm2FFMNfQKozKrOKGtFB4eH
lNEjSYCSnZrOGcfUJG6uYp4rGKow76SIYcATn+YoDVVqPIHzL7tIKElO7W/z
250d+H/ePZ8crzAw3lK0D8VKDGKmkuoKL9o5VFTtChmSJRsIn90jgIpDtZaF
SDFyW4lOQ15HLRmtCXTtMKOqJGQFUbRpDtBjgtDERt6n3ZlW9/mfUdD7ha7t
YqZ+84ZTozLdX/UkeibU1sYRcY9mL9IcNOPxS9grQEOzuElHlj0wb3euPK2+
sLHIGScku4Wq4gY6uSvgxOjbW9d682ammwJmH6m1OdHcltcRNviD6ZyeAOhJ
61EHPqNzqF7jSE1LPrY9e1CVT0kFowKM72mI7aMyLLnN6XChXQ6cB9v1/I+a
heCDn6R4ghh3KaphAx5HQYM0/P9IsToedaEgUZ/WtBEzfn65SqhLXxKuFdF0
+FQjBLOQHHTAYq8LKrVcBAPbTOj2Wgjn4zp+F3/M27w9vZP2xoNiEI1fQEFo
KMpGmR2ldNAtzA8HG3CKemtVorp0r3TDg/14oQC71Dds7wQIuwWcQB72Yqsm
VBbCQz5HcMQ6znkob/n3bChjN5SkqTqcpz4epR5H9zF605nD5mewtlI8//ot
zNkgwcaQZhbXbLJE8txeJMNPKBj+iwj+POBKYrWX3XNONfboqrDvXD68rI65
NLM3PNweUkLR0IbYLxrlIcXSuUMEjxhzdL2JXbUVV0v7/yAInMD0EHR4d74G
lZ0K1I+W1e5k0/oiesrr+yeSc0qNe7mBOG2qCvxxYdXQVqgqdWJwh5HALQa2
dF4tLjh0SKdVe4AcvzkyvQBygt5M5ddN5mMnmUrUj9QUob9yCQHdyFFnA81q
UGCawN+Ix5MSRVokzaVjWNGOGAA+iEukQNkQtFeZHbgSFg8egznmH32G1AtC
/rSErlAZDxIf+UqN8jPY+awgDPccgx4uZoZzfzhYm3yqdG4AtFtrwVX6DWrG
jqsd2dW2G81f9PmwT9Kew4woUa9/MgvK6WDeWACvDJUe4xtHhiAPAneTJziz
DNGF2Hi88wDwIvvkS6d81ej6AnQhyt5MQMFQtQfCr9XD5lEhBZ0p61lpPzAf
VpHw0gze107MLE2NDKvndxndQVEUhJSPemqd0ws87e8ScheElMmklfSfGwBm
l2BJrOHp3lAIKwKY2zzwaCWgVzjpShB3Z1fQgYAV1ppG9/9ej2PBu+KEGCx8
+Ju2e453vNH/PYzClsZQCmEyBtTCR+uQUu8hENAcxMqCN5hKsLWWYriCMmLd
6SPWzJHnbhuqDY8+eoh8XE2i+1RtK/hkayXExf5SkiFSMyk/4zLoKcL1O9fP
ZggytPO+B1WY+R2UsFcYrTJVix1B35ssREkt+YmEUSSfS2AgvEgLR2nxN6Fe
6pIpEkN79h+2gCMT1/q52RBZjCdawYE8XDnmsABYpL4neHBG2LNuqXjJYszl
I1fUxRieksvuzdU65mBYT2FZJTFfhgHxE5/Xm3E+LWe26URydZYwAen9rx9m
DV5JxHVKh9btsDyg4gtto5cNyb+FdmnUbk203LhjdlY02+4WP/chvVphgsEm
vtVFBd23mfJTR+nzwjt/xBCWFY0wmuAehsbT+CIHwDBjQ4CXzRLrNy+ZPkS+
4g5qgWZgspzkKHrZMoIjhRoBfW+1XPe3h2if3KcjTOnoDqnEks2D2RAMrQQY
SsCg6cUGmtL2P+HJ1VtzmXs0I/Uu1AcL5BDrB2TFq3mIGw1g9DYITpRnhM7Q
3lbV8JWXLfFcPk+8vJz08k3fNROvBcIsL3y3igGYudRviFWfsEh06wtt4yd7
BV1xahXPcOeB3P99bgkhdxGg29maqVFNL0boHvP7WtAZX8RPlkCIR8GciDCB
NPO4pvhUa4d23g3gM1yVNmVTuBM806iLvhABsnheSne+QV45TYZKgO27LK9J
X2x0q5R/TKW+oYTDlKYP6Sj4PpLlbxB9l1Jv686bQqlBlV9Z1D1wesRj17Ni
2IXW4Wi4lEDA2aac8gGxVA5CgRzXvAEtxEYY/cpNvui2192/9MIGcY3TBYOV
Zv4qGJK+USHxtfNoFisBmCXyd6CANNVcOfqLgipcS1QzLshzi+jyYWwlv3xx
M0HnER8VX1aVDV6vmYyOvY7Vqyu0fnxyqAqvejUyEhcnmNc0h5fj77DDev3n
qWBYbCyGbCdbhsDww8mfkYAJFDWSHYQTSG9z0gIx9gftCIY+1G0LxjwQ5SoL
WP6enslpLJa+RMJUQs0H/0HCEMmhipZIpjhDxQSAIz+MbpsEbbF2qutS7+2+
Of4OsZ7547J6ZtITHp78COQ6T8JzyhA0jQZP1AkW9QLQ6KFnWWGpJPJZii6t
1jaiWyDO6zTj62eGMxL0uNirTN6OvebrW/F8jPCbqJLh55bz5/5Slfr6L/PT
tDP+VrTgH0Sb/efOaozy3r8VffogoCJ0CkPQ1KPZ7Q9fzquFZYwtehywhD3B
WZR1zT0pwEGppFxC0eoUyjMaND2z8c5eW4+hee4NpbWOwu8IXLHmzRWFIh5d
BMwRX/MV8hIObGNOffdoCqTFs77vPIs9Zl4P0t44zR2YplMae6wPhY4fy853
jzEHec1QKG8e4Aa8E+rRPiT5MI0dPABYj9beLrV27j9yl9qRQgKGU0qJ6mRe
zSkJEXPiUSpgQXIAK1+RETCgi7jzijXUPY77n4wGdw2PMgpnL0HpCtK4npRm
WW3aWa8VlnQa9aLSfc9OkAL5Wz35yeUPnyQ7hPXOVZ9Pq8V4sOLQFk9bDnXD
AspwE+1a23YY4fD6V5Kss6v4c8Ew/MjWK8mqjOXF4/jR7t/F1dKyCAMsb1ox
GHgWYAcGlVbV4/I44IMLrXeKpLj6iWzsqHAr70yE8vxWmE2z909gHdxcyCBm
yIJmFiz3hZsJMCxTS7nHWxAVlTkKx5Ok8OV1sccMy5ATWRbo64mK2a9x8y6q
ngxgB64Zl9pmvRo+HW6FliCnP3fo+gAdhcaxIGN6dRyTmCRD+ex8IQj+Zjti
qM5qEPMznfkZKxlIf9Et/zzl0elagLP48fy62CH6FUn0kHgWyrUYRzrKcRrF
J8VYEDP5nroiP0xx5jOeIP5M3iEiK+jbl0/3UlAf9oxCshQXcOkKS2Go1A0l
Tv6rviFrYQGo5QnYaJiPrgXV7Qp+fCZweQglNA2Dqlk8t6HB6ZME2aiMsUTy
5gNI6jH0LWRIdHB7yryw9ZtWIkbPbqeEe7DVSKlMTxQ2mgdserACeDK7Kf8W
R9eZo16Gk4tgrSarcjkr37Fu0jaaQPPaHaMsza7HOOuw1RhzpiXxd1Jr2B8k
XzNeEtCLub/BoquAsOghq75Tp8gn4/qlyDL6QeUullAQRXmbNtwg51v9HN9k
N6aiLQd6eubVRk/x575D6wrYGo1y+W2BzJNbKcQtIEz6QdjqWdKxNmCfiLI2
3Bgdwy7hn/aqDlFXwMPGZ+QWuVJdSeoEtX+qYW8k93l+w5NfquN1AznudyQa
rtpEyGpCvw8DkB2vSf158HSQrruGdc3V8x0+GVZkMaMO/5O6zBFR+gFxuXMA
Svo2roYaA1SnMsXELUIkLD49fPAbUC1+i28Ze3vt9ZDlcCH7SUi1sWremOSd
9RCmWNrPJTG2UZ1BtvK2C638aL2kIxleksW8ON/vY7vF5T2pPCynh+PifHOT
KTfoECH37ZkRHJy4gL8ltAMq8rbCsKCVQSXjt+QpGdtYmkKUxQzzz5rL5LOJ
U33iv/e4L7OycVev+jMoRLZc/30TZ27EHWvUlLdPzkS5Al4fgKAK7Qpc4EsH
0gWUzcQgVqU5BDiU+AjVPyD2rQIsHOIIoU1uCOIYGhb/+PkIrkoXYEaGnmrT
Sov6n1eYTxUOKYdtqlk0Fwbu2YTuNz5E94FS5GZn0DXn0okAzbiFGJf1T0q/
LZCXfCxmZwdEltV/oLmHg0ZnVL7TFnaNehs4rv3z5mQcmJRB9LysczgzaG/T
hI1EFJ8ZwP5v/rX39YMpSRS1FnL5kW3iYA1guR4HSxdbHVapKA+YU3/1MDUu
uo7yCbMSDCOgIzGzKtdJJQeu7nvNcTz7i9dOS4zlOMUFG2sNOlIiajPiQ/EU
32jqPfd1puFcNdcOhQWy0aBWy8r14rQbKtDNHVmaoeCIPTXrr1ASClWQpVeX
92fx+iDKDsNT76R/75NAg2XzQXLPyQdcVNPrcCwHhlPQcCzAogCIjXiykVry
tdMjDhtFroIfacXMECmrWmkF0UECiUVw0vFK2i9x9W6VfOtIIIA47q8CSDEY
AqRHu8sGrpalqeVW5uuM0yFhYPPFFJrCXeIBsO3cGarOQNwDIVar0zV5fehU
sho7ZsMIJkgu6aupPmqEQcnJxdO5HW/RkaaW8EodtwxSp/uaWoqWOZjnYNL4
VvTq0KtKpQ8Ef/ebbljRkAegnu9jA+DCUxlY4zPqPmm/AzpAqBef6HR2mK4c
VKq1xMcix/5AUaLL8aOhXEsRhz1i6t56MI8iVqG3YZymEa5S0xT+9nnrTxgH
wLU/rsjp1vhwYiP3ESeHjX0Ur85/FCCF2rGU8k7gyAYeqTQKbXWNeroJvqfW
gvr1s5kHX4VgzHzoe8BgVfundKGVP1JmJpJH8jUYTPxBFzgT0cVuIQddbnD1
aGdU0SWG2mh612/qN5zzuMgGcOAaJ9k+La++sh1ma+rvQfSMZ6J0Ow3o1m8+
AK93LGHqqFqS7xZ7Kdo6Qyz6nXandhoHOBSIqFHShS0Jl0FZzwPjMYC/Im+f
4latikGuQ3iZpvRzD8kUraYm/SE2W5W9lPBVyi4Pez/nadhA2/J6k4+DApoz
ITUoWHRbiUvIrwr/nSsy1aobtqADlzmtSKGgALJV7fs7yEqLl2NwHBqmvVdN
MeCmJxwG1gmT5pqzksTu/yp56zjCKztWZqqHZ/+rEQjoDjWiy5I29i7ajrdi
REBEYGN8DvUtkVEfHuBfdTB15SXEcpWZpL/9mUxm55xK+Odi6R9l5BU2Pv7g
d8G2gcQV+vrx3wIwpoLXSnEATuu4qH0gmgFg4roKDTNC6cc0h4izSuoNAZgY
vsIBd7JJWS5j8LGeMruP4FO086b+noR1gpgbyVmGt1lOit8orVC49tKjZuIC
37IBx4peVkjXQOvzP7qrH0UHD6DK8o7YiFU9xODH/YfFSW7u0Uc/tav9rrhr
hd00ilBeYZYz/wic+XvyC4/+LWpi6c1dknGEBrKhDn2LBsZy2fc7xcGBNmB3
QIHjg6VAmWd3i9K4x6mthe3QgaaL2Rwm4rqiivSFltzl3733V4LyGhiAZRo0
w4mZzr9nUKm3WjoJOwo+QfJ6pMBisLqEIXQZ8gs74GFIfz9NACj5WYqCFYYp
L+7si9Xuo9TuH9ThlqnlopUanzS6d8Xg8xRISPYSLk3uLkhWVJf4dIsAuU4Y
gutmkWLe0lgqmKgtl3jzfOkmxwxp6P8uQXoo2Tv3Hxrk+d+VznoEjf5b+kHC
dLe57XbfZkei+e+8cUU/GS+502MbVb0Yd+ay8FTgnXgbX/gTXrPbOPdV1ftX
HhOl8hRTHMwb6aZkOJ0dx5RqlohWpgvaI1khYRkdgkXedGY6SQBdxg0bGpU1
N6FiB9jyCR90431cE/ZZsn3NtN6auHy/Lz1xZqwzeletLoHbAWzDEibNSBW3
2mJUlsPachya2lB5b4AG6Z7Kb4LXaoCMmVi484twR0kIhbIreB80eB05jZOb
W+9UCnygdMBqdzLEk9qMExkIAm/4/JNDcSp1j4h1mq2PtauWHnJ5/CLpy8y0
GiRolaDJ8p0+PJy7/nEfR3MjoBfyZBpcezU1lkzIUmib0GHA06iT9YNRSyVS
XutecQcGcuTFcRaZ8NaMm/AfATHtbE+VG3xXpabmf91BNZ3mvyov1QiDhThm
ThCF8S9MnXy347KgfYty0fxUiUyJtG0t09vlbo0SHTSXLBKiwsmcDSGr23eW
n0QgswFMXqEeyCHWf27h+NU4jeMybnm2llww0Pazg92H4CBzsCLcT8nVOHRN
zUIoRIYACiNS1LAzXZKLiwJchIeWYUStKL31eEL9FJhHw7v9tnwrHOppaDl7
RFub4DAbE5ptx+TI61Na4tzdD1yXNRNajyd4b5IHupqFO/H4af6gegQ/SM75
uW8k3qfK4ALb2Vqj9S/yP7ofKltekPxvisFSWh1/cpj4Wwu/VxUFeKjCc6+t
51LGgEgN81AJ3ZLPFu2MeRouodX6Wjr2+SRkad7w5C8Kq0y7iVL4drTY5OGX
9XlCnBToQRQa5AniosAoP8sFegHPYRVaGTicCEB37pyh8zIQBSVjuKW4hRdO
2KeE9DGzkOs61f8AS+LEG0rO6lE8fX6ABDOwbZF4agGg38Mot+/kK30cjPJh
tO60zah7XkpZnY9IbBsENKUv4luvhtgA3rx1x5HFNk8DOxLUiwoJp02i44CB
EkM1rUt5F4UeUE0eOlAFc9tPo3in/TzYhUA=

`pragma protect end_protected
