// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
EI3J+oR3Mgy1RlrY4GV0GsihyrlJ5a84DCSoUD/m5iPTX3gFXDWd3LtQCYG81n14
DCx1xJphHkB3RfSYzgWq1Yqr6qlZ9QB6ZVTs1VZdT7GpbiCreCS82x+MOEaAdvn9
X8SX4T/YOgPEX+dCD+bYrvnRQNgIdUPXIjLB+jp32lQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1408 )
`pragma protect data_block
PHMIqO8f3AvSVeWBaHmOzb18ynR2akid/TCgbN6X6BpuiV7ae+EKeApArSixbugD
8Ph86t5VH4ZVYGPMzxOyQPQIvDieob2ZF83BV4Pz1jkVx8n8jNyRaZ17uqfnuzyq
qcJBlCha/hHycKLn4h63AjsDfugaFL5YL8xe5r3HiVln8LedLFZU2TPYG7oKbkcN
KqODmxEGsiH779VF2zVLpSvFOU6GzTr1E7Rl/M0pE31dY1AQrF7HTopQTZAYnn4H
TG1rEZvmsfkbnwA29fCzqyB6vBgvPGz7fUPE4tOGXlkTuEA8v4r3jWDK/H0PVHMP
/O7ZBsIkPd4hEKF13OjQIqMIOPxaL988SeLhKhGw7yP+uj3EkWzKB9EHiP7UL59O
Ax7k9IvSGgDPl0zT/hlX2n/lliWZRhLigueU3ZvFfYpAVjieJKMs0uebNbKzCcMz
N0PGPtRGZ9KXvpBv7hTRGmBtVDbWVyPnegv3h7PxRZGKNtCZnJN0I0nnVRTy7/+9
EsU/WFBZdMU6zNuqCs8KK9Si1Mab+pOOe2Y5TQKDPB9pzn/D1hmavL8rqU3OYRhd
QgVl9kGVKBakz+3IW1xuDnYfJhJGgCXkyUEHpK+QnpGkMVqxncn/DqIE92OzxYuJ
MCjdB6zBq4AjmVpV5QWW+KKdygCUxBmgMxIMijCM4GZDQisv69Vait9WcfjHn/Fa
yxOOFo223nUYeaRIC9cGVgs7i3C9qC2DrRiuO2AYPM0EMPbA/c9TBf2nCg5IdlZq
4HLdxRIQ8WYAeI3pHlw/o7iwVGEMc3EUti5P8SjbdQkR6MGTj9aIWZVMU91suDhB
vMqs+hlZBRxccVxFzZ0Qu8GhwEixVibXsvrlXSX461Qa7/qpvvFyMwPjPSzoC6RX
BYhB0wOrYUl8UpQH3etdn7b820KN/kRV751IGURuLjLL+dl5S8wDyRtX0LoSigzt
6r3EMhVZGjAkAGz/dmOqKpIXFcLea0fxjxLHoTqeWT82uib8JOHfEtLVbD45daI5
ocJS4wVVtkrFDq3yHvr+7t0dayeGL5s/gs4j9edF8kR3A2+RDiW/qlvYmKHTIXE5
ZUYkMuK62r4k5zLCKTYUgDKj0zRn5iLmGgaOX+ZNxowDROcgCNJWeXp4VocroEvo
IRQHc0o9fe+Laa5PBay7s/VUi8gcM0i4r23WB49vlefrVnk/P3JCZtJUAPPlYFV4
/iHQkRTirM1Ki4wsokB7GiteEb3BvIgaqhhRkZrKHzky3oMGVkH7qww3U2JdPBIL
q6xYBSElw8MbKJ9HCB/4a+aeLPdM7DicYrrpwJjFuxjkYlCu9y8vT7citztDF7Nl
xguF3N9GrrNcTcac2Bvgg7AdSox/RPFxhHvN/c70mAelDGWYGNsO37wNKZuqisTV
UP+yd78P9ojiwLk1iIYCLDirEmxrRHtuKel52pDeWzDf8Ww3QY3y1flsCJiVC+Gl
D40LC8ahcz5YFyPJVP6RGHe0LB+yJVfnnoscHsRTy/99MMSmRFe8N+UC1rzQrwQg
RJd57Y2CtHIWndQv3JDF5bQw6EYa6GEYOkN2GGBrb5Q2BPwxAuepx/su+fvaw0Cn
d5UIkcqijatXWolTSVdrP/Th/e7jWSsJG/AmMHEOsGlzcsnm80IVIDppLH8Vpt+n
zdtf5RmT6w1K2WWlikAT7ukbTaW9m3L1MOTCckMwXB8uK9MRrFNTT9JgKclhq4hA
Cisc6py1vGJHnNHmQEMzOrGHIfgXbbOn50WKYdfGssRMLG9GSj5g9F1Nj/TI66wj
u3B/wqwLPBFrBaKBkoCAXkV33qXkKU1dpuVtvOpSp1lZk56EJkpQSfjMzqWJ4BEa
4YwKOXHvTiTxxZih7PVNwA==

`pragma protect end_protected
