// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
NxeQ4cEP4wW6nHQvc6k3KXrjNpWccUiSmGi7Pak2va1g8I2eDewcE0ST7MEVzcBsrGHnbU6W6hBj
y86LVwuKaP+k6czIfctFLPj9EBg0dptAMTxPJxMypKVaIFtkOFjPObQLLMigtUIL1HBp9m2pPEAY
EvChQvFOQEL1AWSVbthKAIQRBxmHRyTA7A9gkbCT9usnL1O+9FdUA/z0UJUP1zA8LOKIUUz2KMmG
Som9bBNt6MoVL3i0JUZUAFb3LJ603+gt+nZakpkXBjQgU8wjxszuRCp4hFUt4NX/q6ekbc/P+YwW
OmjnTLH1d2LuGSca+xbhFT5idhcTcfxJbrWpYQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7376)
xe+XXBXC+bVXpPdE3t6/o3ZSII3vMRb+WFy1zA8kukN9Lkn4XnvmzQ5DufyEDBvjqlTy/qTb206U
yhYdnaXxZNRLS9j1DUi0RjDoR8jAr+CpeOCX8xk/iWO3o6t/tTIWAL2mgPAIy/I0g/TqzQ3TKW/t
yEq8yQLxLL8HHQMRY8APLtDgB9kTngUylC3wGnQR9rb/T2LQT3vmOtg+sAkP7/6inL7HeFSdQqfB
vQIelY4Blo+VJf3dx/p5M5fji116TCi4FrlkVToL1NeDN4mQdLGaP1f2PgYfwHOunDDA0chT0QJx
2CgzR/88PQF7Di822FyOB0AKk1O+amxjDq4WIb9ajWqwj7i4sTlLPoHuC3LCq6A+aMgFRegKCbhY
uwkuReQA7g0nAZ6whvIJWhtBT7yijitqtLVXrP9XeS1qjhseLKLvxgpl8pSzLoMBYxLpCohGytmh
v+aBKK3lsG4qHSzjqaPCkUckXdKtvNH83Y+CKkrs02bvEtuBJbsym5Dgandf6EbD54U+iSxGGfQm
wmlTFkcTqTQvYL1hwB+HV+Qa9NG6yxReoyL+5NEQGMap2yJ9kYF0WsYiGTKSGd3sNrcn5OZl5VIT
CbMF0Jy8ogQn9qo/MzD1xvXMGwp73ScAiZmSaXqx3ZqqCOkneoypKLWGRo58eaCji4rUbNVSv526
NuCdmTG3cG+Phnc4J63Je25Wxoiqrb5HdIJKvNjQZbgPbTjYNs7ic2a0JFWv3CzII1tl6UTNCxpo
FUne6gJ7QRFaRZcuNfk21+RaHx/e/esi526ll0q3RH/CH7UXA9pf+NRkuZWQ7lo2CTeV5DabtPRw
RaCDNI2m4YwScRYOAgvXkCxlAw21SZFKCa/kTtz11F2gTOJs7xhc1r9q1npIhLt1Zvo5cD2jALZ+
/NfvtJlSj6fTQI3gAJAsMTVX0riJCA5sx+Hxmhr5exwgjnPIGhM3qKt1gLegTP6jpDHhMEx/AWK+
wXTt7FqDXnp6fhuPMQ6TXHj54NDKqyo/EAlbTu+fj6RupTqzS2F9CPBafxvRZ+KMwj9HYhis3r6C
Q/0ZRCcmJA1k8bRL4gAcy2pCdV2BVyWISt5+p8uat6gsnLGA0nv64tmw2drBoRdXcmwiv5YhN+LX
qx7xONf8agFnPjB4RN64t0gtqLMN3J2j9OQVJCG4P6v4mCk1IS9ttKoMDu9yORcO8P6/8mVbr2Sx
ZDDQV9J16fibUiA2A7Crm5yJqgPrqdr8feGb0YVHRW+rOIdRJx8PwfAF6ze9lGQ9umXh8ZIhY5zn
5ZZQpslC7TuuVMqGjVkZiPlpSsrJQle7dG3XWkE+sYeFwEw0LUH2rLxNrSM00ZTjfz15XFuLRAh5
JoOwUEv/GDFkQz0qQW8zzUCxrSo55/U1yE1SQ4y6lJkPmZJaOfEd8/JQ17R1JDEQIb1nlrVqJTrX
cE3GojnZCFLz96pSf98dBkSjtYoPQxeqiPz+sy3vTRcVMt556XRx+2hP+rAMxmL0L60pF3aEIKgy
IXn+kudSpHbuePtAhUo0JBAHaxO12MXqLprxBnK8I98nrZDJ2Qn9QeHpE32LUl4Jc/D5ROC/+Teh
JTr7X+HyOGmlnIJ0ohlW4wPuqTU5eFbTqTy8Sot8NbU/VkwD5t2u10sBfdYNc7b2FrOo5FW3IK7N
2rGUaURPENIxTXbHqdQa5VXH0jabpKj3xILcXAzMHV6PzkbzZH/NaNNs5VpQmX5TYzN3h0yIlkM5
GXqqCVhSW6UnQiXT3jGnGdymQgvQONEKNzBbAmWXHh707cR26NXpdqqYUj7/zC71E8UcHEeXGtTA
/nv7GGqpfMBGPd7QXMMxW5AogmBkGcPnfuaB3l80P8vfGXIwFZDN2cteWAVGEvH8aDUHWS9J79vY
Zz2PezUdgqSxA7AV04wQALuOydMN+0fDEFOKVuBLJEHe5vLH3eZnPqKZ/eGIMxE4UpBFWaqk0Wro
DI6/YCv+56q2Z6xxYMoI7Q1/6v5LNXNdwYaWtYDMmdJSian+/2GbYHs3zVBbn3a9LRAOcd5QttA6
EvQ2GGvuASiz2FtGpvEKGHecBXgas3ZWvKPMO6njZiysCfbtud5hf02YaJ83zq1UP936Pi0KWMNo
HvOoXA1NSnPNlA8JHGUbL4jiicIqMnw67hyDLegfCpP2gcztfbmhSG2H5KCZalTKLk0F//RXI5nn
hjeJccazAhwoTuI1PP7L4MYHrSqOUX9yvy079mnPDhM4r4OCE7LbuJKcyMM+NyTdv8ALQIb0wnFp
4O/XtAk/CDwQjHUIrWw7T+bXaWVKzm88YDIQUp3MhMM//Xsj9vthTxdkQwPBelQTffNCp7vw6c/d
zBY7UcZD3mcN0ePF4k4fakOJAr0D4xK4T7yq2Ib0BHn4i9j5/Y5kUOqEoXLcHrZV9WWOhr9VBMdK
qk1/30LZ1svydnHqpuhcKE2yUZS7/kmUM5QdfKFwacHxlKz143WMNsWPRQAykC83MW4eiMgCPK7q
ml3pDkHeetY+Sj1/xjKvdSHiWXV4W1iDoApruNNhQXJbNtlFiya4mTKmneHc33ON8UkOJUzo8v66
IamxvmH/i+cxZ5NvK+XRuCARgB6dA5zBCC82IByNhw09lkDjl6j3YEdZjGuJXosz5kU7GoyQHgW+
cLuOthtKPBbKaLGbG5n8p+ldUBtaYsxrIsnOWTUDdIAkPdbF8jfmeVx6Ka9DD51l9zis8RYyX9rf
3Obppa+DDZxOkE/fYY5sxNECdYiK1yBcKbCGv0nbKkmLIKRyruFz9hRqSr68pCCCCYTjLgyzH3bW
vqm2Iu5SrO8IQKQZSub4MwHaX4C6fmLo0ESgaPuarSOFAMpIXH07guYxLMUJhL1LAT9JV1o71srA
GCdZ2CsyFlT6Dt6ev6YbTV1tbj/eWDrxkjaHsm/C35ACKdvE+36RnAxfvD4tcZpFdBGB5svjS74r
8FsJl8hfgG0mrtroSNWXaOC6wwFveZEMqKQIhbWK3UZuBCzEOVzqiuC6z9n28187iZG4jcaATjYR
uzqvu8HFbm6KPxe801PN0yKfQYT9738PhhwuiwX0/wwFemLiR0C6FmdRl6taLEkXugIuQcpyDIX4
J4wTJb9y7mg6NtEDs7Te/8/9HewjhMK5j8uJ2JTaxnrVNCQjJMMy5jNPoKwcQ01nXMBPDIkzws3r
Zue98XXkpCH7NkTGYd2mSQf5p7DCLE9hrZ8SSGj/ny86jVnLHc6X2u7efyAxvm2NACgUtYvcQ6Mo
j5uqYQJ+mVkVNpUcuPcD3zGKu4JL6sfS3q5kab8MEhrr2/qbZ2F0R7Cyu1LncVv1GV0stKWRBNmo
bQhd/7vnWGd/SHQf+tmS4r28Lms3uUDIA17xDTJeX2QsqRBDEvGKJeY1VhsGyA9BnFL89nXvGHk5
nD9bVbfbwLrlMqB9QOxNPPISSq5xC1cv3Pa3q9AfgA25AdF748j/+GqTkz7vmt7hwfH+FQysrbSk
xxWeOT6VejcoW/6J4YaokP9P2hAnptDBRCDN5FMfPek+w17Px06YLjdeRNSP2DmLBFzRMNwcqAIJ
6PkgWAA2Zd5LVEDcxLGdBKzrh+5O9Bgpjk1J2og8aIElvo9oQ3NGXDbNJ+gHal+XmJ12Oabig0IR
BxySwM7+OwGU/GNHYJtYziCdPzsVnJuMrnozA8aAIR/sHFLZMeHWqnJhZXSKUiYc50Bm4Is2BZ/t
R/ka3iL0OBtz71nIhoAwvTE6GCNdVHIlwfEHFR1lmej6XbuLDa2rCP/ki5PoNT0tZtBA+OpnDPyI
ocg5WE12DAqhc2B8gZO5CTqkIHKqNYRDmMItzbKOQFbHJIZjNMiXCGziPJpviagFb2yQx4mantIA
qAupbbtUteIwlbEtPEODXRerfK93fg3jSRJy433hjXMh8sSEqYXkSQ5w4a/ITC8RLMzDEg+qJLqV
haDofMnBbb2axp+di60pATIMl/YyYkNjThgGEhX8sufrZ55o+ORuDkVvswxPLwHDmvJ8EYGJEjJl
oke5hAnzLwzpKv7IqOd/k2/XLkb2KzhGKxJ9uyxgDL2Jh2dSSckhW5MRwW00LWb2EWmt8toBnYxz
Qmt8GxULw1cj5ohMDEZBjRiylKrOSY2DOZGmYXm5htRiYeKxhafdB0q6MfQmD0k+Vbkx+SPslFWB
vCDI0QHy1fhhCj3o6mxamombWoZeJqsEHtpKOpYH9KIQ/vJPwFX05rBa1ec3jIUgx2EWOxm0g0Fh
hz0q7QB/WWO96XVNN26WuecDttnk0JIpDPXrEiyK9NsWQYYBoIHblb83bRUxhcT7Y9y3q1t0VPkN
2e8T7CC7AZG5lLuEc0cZgDtFGGkcqYckmsFoOoOs4es6LqnN4iXNHBEuNxm56czxnTRS6BUthS9w
84IMZhxKoM4BwFxzxO/Bm6uN8PWysPTakDwFtq3woL5GHTY/t/I46XRKFcLXmDfKOMLqrWt8TGu1
zjaI2eiSCBca5dF7gusiwOXtQmTL3RPwLnokXOlQKxr2SAQ653xs/TVDETy974mE4R7CLP22dzI/
n20egn71KzXciVcgfIZEeZSAt0LiHLll2XFNoBj+7FTmkBIbnbeqRgaYnCrdudGQIf98BrEKjXUS
s7owpgFL1QysV0O0zSyU0vdsXdUiE6wFwm33ZlB+TgC7U/R/Wb9JZzzlonIvxJaJRaEWco4Z398x
Rou/afZFgfewcpR39ITy8LlT6UkJDjjOD5CAAowM55btG0i/2jI7fYwRVtKh4GibpEa8KLTgNFBt
4hxKuXjaaMfPqZqm6/5O/4lAOOVr8hBw6zkencRPKuxuSftC0om7qWn9unUtQEhjzEHrNUyZMVxa
L60yE73OiMRbnZKZse1HmAVY6w9+eVD20ybBAxgG7kiO1PXnlqf9Ln/jMgwnyvVSopq5PUXwoO0z
80E/oPB7O96Rhqj+9fOzbJD8J3gKfVpYfVsqZCgGNgIe9cxLWdMAjG3r5lWEJiAwE51A+DxtHM/J
iGObdchz+WgPxJS/HShu92wiI89HulJn/Q1zJmftEUoXp3lU/pWl0ut7pJUdg1n765nTH608euRr
t4OnqMpmfhFo4pu2KwbAY+d+S3kJwIn2MUM6Lv4EvBSRWjDrgztYvAZBlt2N9iiOnG661OjhGa+o
RNgwAaE6fjrrzGVj4NZJEftUaPV/QRj0DmXemm/UrimVqVVBds0nu3qwQz9GeGeuF1decf6vItg/
4YF6h5t79W5sWCcMtPPjOuqGGlOx7zFvvbM/gcWqdL7eAx4Wl4MAOGlIF3DIsTofY0UjohWAXj12
a32Z7opBSfNYPKRstgSj02McMJLUKHHY93Ca9v3t6GO5rzj757S7ulA0aZ5R3UZpk2gVDxwWdvFF
jTuOB69aQNexpgzMkQ1VBJ6h2uRgWsoS+z0M08svZXaLMn3RXVwuxDCffv1OgBywKLc7dqlo2TME
5Hclw2SsRzO+6hHGGmEhx8QactWUkwZpXMTlvCIK2evgIC/O8RIM4QvBz9bmI2O76+gyfyLQTE5J
Rtl6CDzsCFWdp0moV54dU6xJlswJDP4bOXuEhA+oLjLLgN+xRPZqc84S/epczyn71AMa6TKuZ2Oe
qyS4a3ktyKEFVhHFVPfSieN/sntfDWJgNY1IYFOqB7Ra7dqm8Ys9jU56poMNzOg056E6LVndlQPW
TJy4R3qxN2mic9F4IqR+a6YAP5ma/+cpv0ExrFpZGHw5KP/E8ktTvpxfZ5/fdUjpk9eO8y81oNqO
FxjQ49PyOsC2LPVnKZasvXhBu4xwlAfHkLChipX95cLO40zk7FDrAbfi6YSB+atxMyWu0LIkFrVH
ioTOGbnu0cZ4u/6sO8bPzFyZ4cbiQXJ1w0emZyG38RuIOVdtxM5o2mvBt5bV8SU+dNe5fJfq4RPS
CIA7Qi+W3HIhrGFOakgngJw1qqdgRJmFZ0qDhPlRCXRfHD31SQyKVRunw6oAohe6Mhj/NzRBoo/W
edOYYJFGWoQxpyZyjqP3SO8Mmg15hklg6RpmAH3UD6Ensy5a6RazPhgEASb30vTLVrsv8fo3SBml
NiM6W7cE/mh9636V3ixAbRzm0m7752wJ6tYw4hc1XRL+7tLfzyybbUsz1eCyRIbioXgtF4mgmq/y
dQsmA1hrUqdknmvTja6D369YEPv/YFT8v/ElCa007GDCDwSw+DIDu8jE6M7Pg5Bga6rrpm0Un4aR
1j+wT+vLRFyG3JR25UNV0BE4PTgJ7XO6o2QjD+nqlauVSjHiZSfkfz2kTBQhRbYRHQO45DgzEI7I
Yef9T+P82JC8CCfVZ5UzZH+Ls1FvMeTmE7VmPGBCwVmj5aAzf3L8h+yu2I+CpS2xZSBLghKFLKY2
jsugG+wnVFPaTbVx6iL/68yWY1QHWOh4sQAeIxchmdg6hhj0S3FsAjwJ18nZkNqyCtC2aIrZRHEH
k0EauN2QD3t89s5DT1LHXTgA82Rxhj0jb+5p/rwUNkP/cWQp/lmiYvoxytb54Dc4LGzmiyl//fM1
ZIcNM8Jf1E4WTroaqh+Ewz/rwKS1UHMkujmzaIb803YhbpM3PB0ifpbpMLocoqMrFNI+aFU8k6Do
YrxRM4WYkzlxfnQTQrAj5bokjYL1oYT6NkflqO6lLB18aEXQZr6ka8e6cCRijbjawCMQNQP5dhl3
xUeaVxEhdcsNd4OOL8HBMLW+2yhLDlOg6EWfa3j1qjbxF6wTedqEOiMIfJ3z9dkyJg1Ly3weE5f8
XwyBjL2pPGSOOPVk+Guud7RBPROJ67/LNFVRmDg8st2KlqNmutZ32fZ6co1B9Gu9BAQifmUqFHRo
CdvF4dCyJMbLBdEO5eOfO5B2yJbojacWKjxODPtoHNc4WnHS0/UFUK+xeb+6ZlNj70FmrnSfBdhb
1YZAHS7yLoOOGIjD3ke1TkuIjbGl1Lm0OGq8rdwj8jxTmjzx8pzu4btDDd0nuy52/mq4aNpBhefN
lfeqHZY/6g69N3G127actuzW8iAagVkP5Xskb8mg7tEhUOrbjSTcSeuICSxnfZrZjgqxscNfjNm3
Q7twAq9XBfHcFnYIc+D2gzrtL9LV5wTEA1iJgYx9hI7trKN5X/tCBYfdN7vbgm5kiSyXbGtY+DRr
/V1ZXFaazBm0ckoUs2Qrq18Ly8yOcZCE0s9rjH6vC4HuwPtBWVybcR1MNFgA9d1TdPwvVsr4rdf0
tzixSjPKkJ/W1P+Em8qtEueODLUEv1KtamB0IwJG9AdRsx7gk7rgoRLcYh+wcK4imOorSysogDhy
0CmUoEf1hUopUzu75EqGIUw+QnHJYOr2lSu2lBiTpdgcCn1rJSa/HFTQy3dSzqMf5zc7TojzMh8Y
sYfLzEM4W5s+homr2thDXnaBR3spyvSeV4jKhBlYoFYzEX+wvcaPVwV/0laMWr38AkpczgIr2nUh
JfpiVGg4CN0tod9mz+tonY6nUV1B5GSsFSCmK/r+f6GOiKcmxt98mTVPuHWPZye63q9AiaeR2zoL
uwW6wtZrWK03iA+6TwKywMT02XeRYHcPLYm0JV8R4wftci0ipVcG/oQEY8wH1s2MYEq3HfcFtIzo
mmj5IzIaZsPGhm8li+TNV2xhoBJxRNn64078ffLPvsr5/tuC83VTvEcW50FLyymUQBf18jW472I+
diu7ZQGDWUc8Ox/G4ZSbRh3c6YCJd5X0vN8U5GaQM5kMZGA+56uVjJZX7fi+RTCL8VtRehRH6V2K
rrsdSxD27kOPKlFdka0aaGpI5TOdurWKLegxerryHU69jf2cWSVsZgwPC8sBQEnN93IzZbgGDXN+
bqDK6S3yvDym7GBLbIN/Nl31sKggWo9DclgQQBmxbcJaFI/gp2Mr0t1mclkwzdAKE4bjlq9BwvmN
W1NXyMNU8Av3PGF4/H2L4pKtlZq3sHfwp/xz1fzHsnmDdfmQqZBR8kCWRoBn8XtN7z46JSZU5A3g
2q0Cndw1uA1iWhbGYD1SodTWyU+KRKMxo1LvMuMTlqEegOlrq0PjOKN6Gb1EFrzwYjD6xsHWRcZ8
wAJ/mQ3UucbDHOyq8cURBUGqHTXh4Z/s1h7ntF4nx8m/04PkgHyndD3CTvrhseYSp3mFsVvcPIMh
LxXXZsatYuCQssvoUr2mB0KhSljuGZDjQnPHu6Ven99zPsbZBohxrB3pHWIIL0gq4MdG51dYHyDB
p6Z/Qc32tFUvw3KMtglXrWo6Gz1COKUNXBEy6msKye4FLbnzIz2SDYmrhzPVjEWKgqZaGKOOv8pO
TWtVTXtz8/3RO2dxmkKZqFppVS+GlZx5YYBBmCWHu/q814TMEJAEMIzr5mNcdMGuIZFyg7WTyu6z
3tQSt5PiG8aA5bmsdHMvG+UJ+AdAXzDz5e/avLK5YHkiuxd5ZqKXK8yk+ijUOst9lL6uAFMMNCzq
x9FkXZVQDejWsPAeE1Pnse1k6Fyx2HtFYDNwBU2B45RS4ZpmP1mA8OTcr5clUvgcwK1t5qLDAyIr
dOA44NZhcF/cSbxNBfreWq6tPx5qMceo43jfLNyX0eO/Q3N+9qMJ5vtSzrJVgERcTR2VVfU4hi6O
9uGoW1ezoc7GH8fZPV+O/0wPSquWg7WB54M9BJKpSREQnVUBWb1qgWggsJCpCWTBIG1KGAkbjj/I
vIouIk0vSBNtMM46WiS+Rh1C9kUX1YXQyU8NIISShXtQLw4DVkgWIYYkxdsjmFd7g7zVl2abyuVP
hcXgobfeKRYB/holeig3BrUx/b3Gm0m2Qwe2t+nL7vSCt1qOWD8THDcyPLIN3foNeB2fu3ltbVf2
J9+NlxgI7VyAk36NLkwvY0CQOgytmWkUe2ZsZDTHaZ3ioMwJng4iiDTOs9z0KNCkCzDGpawfB695
jaDevLuek820xvzvxKjvpg5d44wdIJBCvactUJjbcFrT3i+0i/l+txO+0A4rj5U7rIOYjL3SYkGt
1+5Q6uoc78CP+LaSRJ15x/h3IIouVOw2WLXU4T9vmKySbM4NymxHHJjnK9orhrED0x8gjj6oo2OU
SgRjgk10zRQQbMRYlKjuc/orX6BhjAH3W9pBQ58l9KWUgWq5iZkDLeZkWAlarbG9Ob7y2530mk2F
pyVz7HHOO9jfO6yCKWIMwImZNLHCNCN26dSlnjBwoubJwhul2Pmtjy/Bt9c8Roia8+aVJnfUa0HC
wlTzRKyfNAuyz0edYbspv6eJxLAE7lTUPWP2V/kddBZuZZR+0xWvWjfjdRwNwMlETKmDiS0why3Z
bENq9J67xT4FhSKl0w7WPcz2ROQDdIVir+bPgY+P0kMReQ9kZgqWTEBIv9Wp1kjRXbdJ1voIMmgS
v2wtYzb1typ4o2Z0ujiu+8wKau4ZP3PWf20Gz8XM8Ycf6vEB1U3+3fKryeRPKQCtgBGyWjYPIMkh
wCbLgmmUAkXAHxE+JiK3JvAlwgrMKcLVcVyMDkgBgzHgofkIyNJW2voW2molDDrV2vPv0FNEzb1z
j4ihDt60tI2j2AOD9geMt8liwqEYrMJB1M6D76rIg6JI+Pso53jyCOtThrOd1DFyEodqjI1cIme+
22EUO2C92wIVPirLk1SPjn/f/0/eS/aUKiOXzi9Sr4JEqIBU80Xd7loEuvhWQn7SAaoCBJdBi4Lk
9MgsEyYrywmT0uqR/unpRe0o0Bv+xgNlgoWWBS4KT8jOWhOGhUpw7h+rw9bZBQIoWDL+iazVbY/P
lCr7tiEFZ0UIJN/VdbPdoBjPze+HauUkH2Uw53jqCJtYgH+JIIdk8Rk7gkIi0Z2Fbmuus+lwfnLM
gOlrNC0uAyahV7BZDItx0Xp9zqWhKn4=
`pragma protect end_protected
