// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0GCi3gIuAFA44cEwG/6K+jAEOcP5JseqYHOiU1fwjlFp565UxWyCU6j1JDhx
uyE9CiV/TmOrSCgYLldGPu2Mwh394X0eB8C2TpK3Y+YU9Hxy+EWDBzspHR4h
b+16GLOKyyRtsfHnfvae++GMFt/e82AMYYITxhop54eWkTdVhu3xdQm0Dboh
4QxBnmzNXxo9eBSzfeur56m02qWmdJpxz9Fp3K/VA2s7GwTmGdRSjIThYBA7
cVwxYGjwexrgw5q4Fby7BsAB3N/U4fjxofKt3o0mCgxusMThu4TqTPOKKlS4
B6j58zTM5kgwiNNAUQH+BNHFca9wVeY3rzCZ+8r1DA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ERvSqR2yPxyEFcp0S8SIqCiSu2tr9ARxx7bhXmc340yipeGVtAJUSJEW0O99
ipVV64SuJZ/CCrQJHHoLh7JZFOeADROWtxD9kAZtgxOuS0kZb30G/I4xfpSW
L49ntWQ3+y9n17I/i1mwlq9DN71/qlBV4AZDT2wFsN0pfwQtf6r4GlZdkz0U
8gDtBqIY8ncvAWJ5AjxsnpPNu942SajXNbkLBhBTtKoLuLEKX57mYU9I5ebT
V6gOPF144pVP3uB+OMHeEHc7O39lsI5HohlWq5FKz1USADMFO/Q37ylH4Pdc
mvDDWGRB8orJnNoCR0rl/nAbYC+9EuaWxqVuI8Vy7Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iZsZAO/LCgsrGoFJtIm7+zblsGovSSMYyuM+4ScoTtB6lcSZncgrCzZjtPR/
EC8mLUZMLIGIJq9uuqPliGnZ1gynovusoJFu9tiz6eB1MUXQWE29xSPREnUC
P5gKvU56oD1ivhFxYO29FzbklCIMesQghoJh661udaukGJt6xUoil7IyoU8t
YPua9dULd2W2JzLVbFxF7sc2CmHFrnMtpvhUQlsNqWBMKfyNrws2AbVEGMaH
X4Pn/2/pTYF/ud3mdL1f8Jv4QVrIHV0Kixh1H6Rnqv8c11snehBe8dr6AHDy
uTIL4qYE14p5kCI++tJwOnvLwA5NIr172tiawma+XQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gyhdF00KM03hQEBnBA/3mYUmxU6hb04JwFnPf4BGnGsxnAOJcKIVQOMt9fS3
/8zMgk4vJlSYSR8Fhf1lIfpC9ZUQkIyIgCeSc3ohMcxwuxW2BMF8sQr6uSfl
N/6sMNudaduIW9Hu8HLBkkeJBX1NlkAZigkUIfaJc5HMDDHaZQw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MY9t/w79KVFRpvPdZMmVAklBri0A+pH3DFy+wKgMDqIJlHq10aZrAK15HscX
OaRMl73dK6kkGGTHbUJXPnYiFQIEjC3o1pntBVhj3Glg1PgLmdZMVSAJdeFW
qa5OkZ+8/neC/yTXer0VVC/yqzGfAhXQ+T0i7lJaKbsft5o8F3acjSwflkJr
AnUQpWNPEexGpFx0EXPjkmHAxlUIvi/eEvoTyEH2YXrHpMNod0e8xSE0v659
pGTG4Zwtgl7uza+8Y92gg46d9zpchWPa4hntyg4IuVuphZ6qOIyCGbVV663Q
LPbStnrvvUrP1BSwxkLvIJrfPwQ4z9uFEtcvb4dl0xsEkIjKkwrMKetU9vae
ukHuG4irQA9YXpkrjOf2YqnE11IFXjmAxAJZ6gg/Nv2dokRNJNPAMYpO77FA
2rKF0ahcChy8ex1Tqxc/7RT2HvFqLhntTm5F2zz4W24nfeZdP/tBLCeeOKQz
pk3NpaEFzQWSpJEKOEI5AvPDPZLGu4yX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lqCmiSDqlwW16zuKQiknuQDxOhgXBXpPXXAGnFJNmSvHtBCqTLupkWJDMKzv
adpdDWXs9bFOBQ4v8NUP1uvz5PbJ3Z6Kso9jHzuCAoROjNXRCC+La2+G1AoV
AxsdTrLGW2cV7mRQ7B0vFYyE9+eegTmoxHl2xzRcTK2GTGqZYyg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gfYcfOOL3HaL045owMujkFqPuqmuKp+qgrRi/kMSfCu3wxm5AhUn9LYiK0ri
6UrzimpYewCORqDNPouUMECHJrrFsSD43ou2nBmMvj3GgHzxqchNheHy0CHa
bjrUlRTWWdZBrKeKCVys6dK7UL5JsPsyDYn+3ssFIcjgHt7MH8Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1008)
`pragma protect data_block
hFttLJDV4meLCmscHy+qwJ1su45CZ8w3/4JzCLB4W3iD60CmAP0l4p2MdmxZ
w59WLrDkcj3xuJuoxRec5dZErbbPzVE48qHIrGQpGKNYarz3JXAXF8kf6bec
FBoi0IjZDVhcuQpWLRccm0wHbPFSqp1DpK/k6zdYiv2Am9dczjLClFscxF9l
faHmoz3LNyf33NXdRm2TyVF73q3Oe97f5IhLEvtnZORS+G8HJiVkBpS20XMv
TOEn7+8yOHEIJncRtMcpxOx0rI0A7S5mjfpWUDH2bCAkh44kS+YTJo7LdUwv
Ants/de6OdDoQhuenFgR6VHqqJLmV9k2gtjHhtxnv1Gro7pLQ/aorueqoGx0
q2ZweZnC0a07ztEPDmsIwEbjQKBPdyYEJS6CkrDW4F41HzAN9WHnO2TuEgER
uBLDhiYl7ZnOu9pKV0HW3qwHSXlwIN1TXAgL0SyS64nehW8n+y3PoYKrmUTB
THnR+sLIMiXleR+sVxUB7d990fsV7EEF2Sdo5H8+erzAKrsDZpA7FSGe3+bq
viQ93QG7rnMtYSmzViDiOqPV4C2M5MQfcM0rlxt1icoia9u7al1oYraxko90
ssg9twodW051AcXmaMJgRCVt3Lk2gVcbIBp7SlR3/guRJ+nINC7Zu3Z8wgGt
3K0oNg5cBQ2FPcx8SNj0e4gaL5gDITz3JozoMqglpvrstF/Ojab1rohaX9Ib
Z378lUtWGHfBOqX0k30KtofdBd14JbHgPvOjvS6GN3v05bcnlqXrDAkhL3xt
zkAUViK+G2ne3GSK7BaW1CejDestIjntgnYbP6+m2Mj54UNN02uBTCOgY+wl
lU5hsh7ILjrLuQRObiUYmg6tNYatbFZSaDBo9GaHwwzpFpnISOBX8yW6S6Bl
FySzc3rspiSpJJ1cxGHw+8LY38IQ8MtTFtUqZXRtqh3J4D84qpfhU2g3qkXs
klDyLHmOLm+BbV+X61iicpOGzzoFRqHHvxnCyBDvsW2C5601j2DI1ieuUZkV
RgQ2jEkknrRuElIbTwo5gR+veAnnGEsBf3gNIbM+IEB4vPvbtPWaic2BGs99
ffQTgc6zbVInW514b8Rs9a896gqC6Gh0Mi6xnMsTLyvIhXsHPoPy4PrUfObK
O/8CSV5lxXp7zkEXQ4kDLHuH0MQJDd58tmIDcLjM8warBDYeG2R3J3mgmcSt
bxG4WQr9rQmSyfvimXsydxfJfQQk+Bgo8fzL1dRXbeGzNFXblxkmNB0Ohy2Y
dZdU7VSCyIgYznlVhdxiGXJXoQ5bWJHx/4J8sEaxop6i6ZSCBrX2E4HJDLbs
ChRqinlVHs1eW+C/glUnBRzI

`pragma protect end_protected
