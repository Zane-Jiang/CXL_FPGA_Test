// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
T+CysHyCOnazubOfbf+dTbmeZOsvKM9G3+TJ6uuTblHs1ab53I0XS3I8vrFGN68F
cFBZcLHhHXEx/1iRjmsgNo3Crf9UVsUGIVbcMD7GULnX+o2vtvqemTuTR9vicETX
7mVxCdnOZP/SV898MADNAJ3czbFb73pVXHIbvPCHvZs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 14832 )
`pragma protect data_block
8Hrts+2ujaajJhCgofQwxd7/rsKc1rMBfdPYf1QWcszhZK4r++n0fsEEelMvlnaN
5G2O6XoesufhVDgdqFZ8XmoZCxTUTC3f3DyV5IyyQaVOpvKT8JmZjojWojMYL1vI
aPfHx4Vbsmw0t0BpfDMv983EaOUMWtMdCxodeCROKU485ucKsAsKi/fnqoAfa10y
CjtD4/qzF3/q980JvLZ4syka8L32vLnLf65Erm1i9xybgBbVSmUj9ntk4E1ZZeyv
xS1UEuWNg+0Zng7G8YyorayeYcTr/b66desRkUO5xB4zO4AZICXVx+4hhCeMv/O9
TCGIPOr7Vj+Kvd0yjoNaA4ealnMsAZcK9uD8YaPw/LN3dFwEAmPRkxcyJTx1Wue7
p8/G+zsahidH5PnaYcZBhReejtW1m9osuUZIwr7iD9GfpGJOCuXiO08T4JcoNtrN
+ifQ4vqANdQ2iGHZHB+JF6eZvzib+VZr1+6jdRAvQCIfKYU6n2iRj2Syll2Pvffi
p2OkhmWpl9XQWtTP5/UDfDqg/41QAw231gQoEznOVLPyOb5RclEGAwl//h1Lfnn2
dRorFsoHcAc/ef9tYCMgWzRbItdGYEzwbYdyw5L7ZhD1mOXZJs1xuFquaef/S6Op
KqO7dB/5CKM4tMQggnjOn4ssD062/kQaRK3+eheCB2rTPO2vvExheTABjjLAwSOH
z/fT31FitIJt+LXND1NzGT1MK7wpEeUTwr28ZLXaBKDKbj1jTS9z+zK1OKaOM5XU
3Kqh4Q16/pdRsHZsrQdWA1lC1kTZpt3rxDkZuDyjTnEP8EgehjovQAe4mcBTGKoD
yF4X0TXcLoO2zkQvuRH7ocerEzCkad2ZDbNkmXs5yJxaGF3sYw98ZbyxmMJTZUxc
oDymknB+hrYx+DBHMZ/e3WNgSHiCaAGQe2AAoxG2TcHS0Ab3v2u7qyxlc23AUvyB
DOtakbZxmM+7+rWBqI8V6KzJSkfbsySfRmf6LK6of9AfRnPBCkdwDhSOM8Bq79Gp
RqZbZqwHbKP2JqqxD6r4qdKkYrQU1sT6VrK4wd2hZ852gH2WUxlfxiHx472z/2yb
DjcPAKva90K6L4r3rD7kHN6nUhpfEFED5yCNrocEfK6gAo6c2bixHrye/ug6kpsP
wO8rSIeeWzOZDu5B6MxutxQrgUTWugNIz8tkXuk+E/v3pZdqK6l5yKz8JLLkwpE6
Ovsl4sOhoHzZpUontdh/+XHOEnRXobg87XY9CVKdzAerQmvW7nYj7dlli5gUkt6p
Amslnl4lkI0F1Gxgas+Budvnf7serOKiS0MPKt+lapYign0YzeZThS6L5LAnp/8u
9fywVDMTxDePleqxCux8aO+jnFcfxksnCuBKI+v3Pdw76UaXGVZXRuiNIh5HfMx9
U0Oqci1y3xXSdco1pkjEysu+jdNNKLly3tnU+eB15kIQiF4LoDj7S/EURQ1YwC23
z9S5Cab00z3trWLilQQXCJyywETTwrYF+a8Wb4V+e5f1nLArx3c0BSuqazAXBO4a
UOaHLrG3l9bZ65rFokralQwg9hfZTR8/MUszD3VQACnady8MEYIL296CPjfWNdsD
EWkJSHS1DBU7ilPq/a3VTguPGaMAheyAn1EbxzcKRQFoUb2lcWfvtmLIU2FT0Z+D
7cI3rJ0Xu4U/7mTDnTBTjNRgmKQxRVj5BKcfO7WWoLy01xAKcBkO+tu/8QZ+0aKy
0XHwTmn2NJNVCJtpC0x1D2DVDvL/02SdMxFhmHbuoIcQ+h1zfKsDtRqBzp8byE4B
2EN/RRpYiWmQGqLkSkkRLc/gx+Z/2Fu9JIdiDyz8CMgq/R/Bx2qK4gjuyUaqn18N
LzH1zZyvUaV96gLjnlHUdHXdy2UZcpKVR+X/Okw7wJG87CHOro3gud0GExhaZY97
xbjGveml0Aq2+1YICS0AQyPtec8UnvQxD4z1dfCqoTaoCPP6d2HrnuAqw18hCEYh
PY12nulkK7QSTCGaBJt1/zvRZ1TmSu7kcigtY1/VVgCjLxMgkJOpxe37dKxlrdxg
uh67HLmh1sTniRrNf6X5I7mhZ+GIYHAkHjuBWJztySTGF2+VnLUxsg/bqv24YbnD
mhqIEhPzfyV5v4F5VrmFUkQOk4kLOM6vIgcVWdB6efr0f0Ooz/RRWyKe8BWV7FF1
NCNocsCq1/06atwugMdcQ8LYwB0o4YtCe3VfNvjHRdBU/03TT0luN2IoTP385jcN
JYXnXfgUI9nQKD6MUiL0te5Dfgr8al50aMLIYIrhJUow1Rv5E6+gT5rhMnOloIAc
I1qiRKfNvq/m8t1BRS7U7M9gtjSsdRibb5cCMWh7FWpTpl25yZDKEhWpYZNWM973
ZB3FsKpJ2g5F4l0InMU8WCr2+CQ0CIbC5WWDg0/JAAe24SU0ysTe+sJnEU3ZJALg
mh9XetRrotvmlX/tMaEuUHD81wg2ez2FdQrxlGp+VgSz/+qUgmxyvHyrqyr5I/3r
gQS62Gx/YOFTAgTlV9t0ta0hJuQJN7R+IkxxGO5Cj49KrbgAgmY6XExO7WyoscYQ
F6cRMo/lwAO30zpeZWZQoLvfrOFGhznXE0NcOuZeXV0wPTuWD4O01IiKhlhx/x0X
hCjdcmrQW2DXWvoYjSpX4ClGc6vVwKAjSUr4SnHIjQ+K/uRxri34TrGUOCbCMuM4
LbcFrt0y+ajfvsbU1SAOrS3VLBT5dmLveZ89qDq7DAe8Kf7ZRRjjYWbkH96fxn5E
DzoA+CqAU0x4Dy7PKBApWyOrvf8n1+LxDeACylhUcxGxYQ9Tz41NyYe56KrINL+H
Iuee0kb7iS37Ev68eCX/YZxogbO6hsfuDA0JXH14GBLIUZhLDkxX9p1Qfmt/lA4f
1czq2SsgcCK2cfbpEqRwwNCaw7l8coGMaaMS4W1zb0plh9SsoZ4f/7nmEVF/YvCq
SDZZ9+Zgudswe8eOCjjsNHsYisq9kj24GD+ughVLw2SRuUlPnZIHYDPaXwxUz2Vb
vZSHmQftBnUyMpV/uhR/dFkvbhuUgqaN8pctkqMp2NbAOlhT55Kw7Jme4Za5A7ZT
9lQoXiHqHaUyLs02vf9FZrPS5eRcPFym+dZE2Y5tHCSeYCpxWFbB6pQnqoNhJ7gK
8V/+QdcCFpK+fTifMUeJlLFagjuxhFWVaSeSCdfCuGe3yKTekFRFUpb7yrukyJwD
LLvlNXKUClyQmkasfSgW7a/BmxJFO2oXh1S/5tlomOrsdD0WXTrc4iGSrshhZShZ
hF+Arov79NYzcf26xEg0Dse6rK5tIJuQW7R0HmRH2Kt1z9c1b82XSrwMYdpXkVTy
BivtdbklkQyXdbd0gUsLBn7sHl9uC41N2W6a1KW6AFqtJdydCjU8C0F1eOZr34EO
HSagnxqq+cwmdiFJVgDw1Qm38rqsOjVb2nrcaQiO+vPC/gmY2//j3rFIX5WsC/mJ
0SZ8P+oeigCf8Q+RJnj6vGsNyvBez/OpmMH/ilgkGVUN2tPUGRWOI2DYTusQQIMe
qGoqCc8xK1yomLozVX0G9OP8XJr84mruL3CCSTJxl3jKKn+X+Rd9RUrm6nDUJ9mX
hr8jRDMQ8tQ1hDlZHVsvn9sxIUBLriXbbQOz/yglZK8oXTEqiG1nrY2zXCcuL3ma
kWMm7ARFcjyldGv+N9/kvNiKZwbxE75hr2H9ICys0G/O4dapgYlIvN01KBmX4rbx
3Nx/6aC3ciYXsMKlqeLsSNFh5115Gkm1JiRezoL8vvLbTi/9kRTatfPsS3ADm6Fd
DXvEzhnH5dYRB3oeBz+B7Tmy3isv8ZwJgz9UeNDzecO12hYTta+uDAcYALXj1dWG
rsyeUf9J+8Tv7afpLUkW7ID0EyQI13XXDQQQ8ZmVa5BzQP8Ag9BO5JVQ2w40LSXH
3DO2ZKH4e/0/rKyJDNOytSq9/VwZ9IACfKgPKzi1Jg5O7kt9mjqpxtbROzNyi0vr
OLSliGALLsnW/YoExoyIJeuTiZe+HvR6B0wvfzw4WntmJi184yVupTWEDX41I6IH
pgYzz4vtD2M7jtXE+ooootCrSoVCkl8AXeozWCm3UvriEo4s2ARvh1/X+naSyjTv
u9GrmUiZ2tzQMwpjqcEm0RNh6OqrS3l2frZ1J09CfzQcIVN8bBur8KVNGOs6EkoG
Wi5bLE5P/XHVjbOUv9ce6LnsKk0KeUBn4STFkXhGVy/tvxAS7QwH0ht7TPKi0LnM
aZrafcEgPiQFcahwa8ZYUbIS+pOWnmEKedmx6TDZgZeq/+Da3dISetWyLQXS1WU2
GlIU8baYLoobfIBl6z6OVpALLNHYt0wBqGvPQcBlLqQX8MYHZvnF30ck75RKaHqn
YGXGiZH7pjo+J/6N4WPbQL+A668vXBrJIrFI78QadFEMGK+vfiaYEo3RnbEra2MX
bEfFVQBXdt3Xtu+b7byX86iRDalZljkAZgfq1xcQKgZTUhqqsoGwsXlq6YAzdNGQ
hvKlUaI/XGjKvtB7594Evhx0u5oJWMA2AH0/WcUHRnhkI026FQJ+Rj7yPD0VZlNT
Pmnepd6aIFzfttF4XoEAquLDwVKf8IsbDhKBYduWl+6SKldmFMbW8P4cuQ9DEetP
KOn3p53SOhBdDJv9EcBS+2N2aBrXCvFWhbHnWNkvClffSUsmYlcCsUJr94Fre1i2
MqKSESY5w3H06s2jajHDvvV4BdR3ySWDERoNExy5i772qfs+rcuslp+qLqcuBOaL
LnranKtoyRbZovnJqlOiLufaBaSSUZ+x47vBfv5TLLZC4rrTKXJfpk8VzukJKhFu
a1E1jtcTK5d1LA7wG+PiLC9VOMW+US20/+Y9DuHX7h5FAvy17ykgS/hIqbdKRbRz
VcbgSt6RhBWitPOuAFHKpspZwbb3+GFXspfesy5G0pi3AlNX6djTQrc6RzncvHtF
rlE5FRdG5D6eMY6IKo2A2x+MIeS/6uPYe0zcwd9F8xXBeKQvMes9sjNtZJ9BMNlV
eazaUcJEjQ71CEe/gcQ8FLCU4eztBsHhOQ3PbA4vw7tY9J/HMMH5E+X5fZPlWLQ3
3WbcstBwx1Kr73U0wN+DB9tyAtVQrIkVy4wEvjL/IGU1TdGcbwpA0t3+f1JDEZBk
NPUybkLmMi8ON8N8j1AQ1DNoWp9fHLnaq7K1qqJnFB69f7xUtu3mbb6jRdhPbTFM
ZSAm29LOUVnqaUJdReXMTso7SyuSrWhmY62RhXDMq0wtT94xpHG2sv/s4uO0VeYz
w0NmcesYshIHycUHyCY1s9klXXHB/HiIH+dT9bDI43RkM8XxoKRsd08V1iiinS2a
EgQyOSOR4INl6OpnCH9xRLsqMBGxJWnd4DwxpQi6svOtaguSyEG9jmDU2XZzIjPL
IcZdNLRU6CPUM2meV94oltmAFusZgF4Gj26PLIvkVHjTVQxI76DauH2IWnDTpE1p
TFoP1V5QBaVR92x41Z42KwgzIuTL0cQq9XL2VE+GcOCZ3bBqP2BcHfdniA0KuhCa
2NzbrBlgGyFAKUqYxC0qTgraYqZxQSsqgJLmUVaBawU2OwLwe0ngksNMOU8E858O
rht8uQEi4syLUXxShNee7AJXWQz2bHr9IuQ6NGww0X3tHejFm73cXhckdMss3AsH
Zl6liOU0wbN0hk/ZZUvUj7XrbFCeLG/Vn5rU8GL82pe3VCTUe0Rfrqz36VuEKGC6
Azi0tDG2upbCLsaAVqh3WFbSGgFEvirDm8+sLAAa25xw1y3TgndizanUcQ8AGQ77
PONbbQtiFvFwuJRly6e9MwdcfVYsVZrbfegJiaP/El9JSobJKkzFTxOhBp26Tpzt
91keuCqywux9TXcqX6st6oIZoNOQ0thYVC+Vdrweg1+q2iPFpqNpp1PP/mOKI6BA
JsWLfDpbv6heqVkLgBlSWOTesnb7sYzB0s6wHDBfqU+DZ1HeAQF42dtgBuJKNr5T
Uz9UsJ53cr9rpZL38CfMGO7ozLhN3lsXrCR/cOM5sh/Bvj8/lOLWjQ/NK2ZelS7z
OA3amwYAqz1iIrrfXFWiHAMb90Eg5E1LgRaauL9mANcXMxQxZfaPov2YPW0jd/ZI
6XfFaV+V5t/eU/rRkLqq8Da12+hPdDxYAZObdEtnToU02HIMX21bsm5G+nMdIDWH
EMlKldZVh8eLBG+cE+uNIzhYKwC8dYrcg7gQgeLCr3aLGM+EXzYM/ussvwVX9Yj1
5fA5B7wjQOZNMX/AoMFYPGSXvpaa97UOCaX0SrbUYpDzvl24GKoTe0vq/n3oxsZr
f10TMYEiBM5g0YrqwrwYAJOtnQYWxNoOZC6YM5MMMTrvQbDnnzHpqmZduzY9z0CF
rAOkfxsk1BAG3lDa3/fpPeehYOYXBkNDmVuamcVJpLRzt4YLuLrQvUKO30aHm0cg
0qp2tiU+w2CLhn3u8sxq65Zl/P3SKiEpsnMoLEFZrSNGRsjC7NBVREas903Zv3HD
zch3UiGIK72EIXIk1Qc17htRYagX+jbVBuNvrN5+g/EpdQPXrQ+PikFksSy6+aev
87Ar9EVf333tyk+5oW1Uhpta3nhlxZMKl01i56jHK0xeYgn3DOSVBrLHpemsbJDU
nxfQpPZY3Q/HF77V2gvl8+VtX7iaWOBuAyhd89SDiB0ZfItwMWilgyQvj232hHgO
VZ1YZPAOt1Uh7oL+Ztosd5Dsk2+ZeeLXK62sKHK3Uq2Iyo3jFeg+niV+sOE426mc
Kpn+iYnoVPgSBTQkR1yzZYA9bxRUptHiQL+OIdjmYkH62jXxZ45fBYMrQyyifVh0
C9bnadcYIuV8HBxjRfGl4S8SInLMQzGmNB+wBaJI5cpb8dBkiKGUa6gFy3g0FTbU
y1sR5PZxo+9UNNWv3D/eSTwG5tTIV1qGEJh4sf/d4EmVtdZ9OiE0R04EPzO6mDiQ
Enx7Dp9rM3jQif4lmuAAKo2n5GLsoZplnuv67/Hoj3e8bUY9bu8z1cr7iP7dbzgT
rxU/2jmmIvUJtAtJzM+GO6UmiLVxqydB4P42EswdKxV2xe8cB8cCPEw3CwfGHzbx
igOVrVNmD7xDUSqnN71w9gglaHhccsnY8YD4hs9ebee+cxf9uFeibLkeccJvZhp/
+k7mDpl4mAqI8bqap6Xq3PdSBb62sMAEmt/BIA9YE40JnKU4wyaShCuA8qq4qHJN
aZ/aqavcl5rf4zk9p3HubarjietBQVNDOR9AI4nNxAMJAQMCUK8QTq8p9pbxRpvK
VIFY1/EHc8wj/ZlJbe4O4mdViGJAKVS/2Op1j5CnkwrOkJyrgXkQ1nrOW0pUceEF
zQ6ApyjNUeGioaerhIv9cZW/6esHLD/IwoEUOCa9Gf6Ug++dyFqEA+xq5yCZBWoU
UJKikb8mOp+wD4VQkiIR6ccbfG7iErSZ6GusCcm+JSpmIeHyGygcGNsmwnluaEyN
N1oZgR42M0JtFWegZtGJZfRbpylV+lBhngRPhjYV3lrgmZ9fP/U/Q7AE2+d8Azy9
s+za6hFf4R+6fIvsMc6cAQPngFY6wBqW2wlbRPW+Pyf6XehIogBXlMHkuWREW27Y
4jDs51DacLv4kto4qKEbzsZcf7Hjx4h9goJ5K1ylicYcAIpIBmsbs8wS88wHSfz3
eg9vtHU+nsPopTrm4OyYlJfU6GYUogm/1RQptg6Wg065QmdDeu2s8a1e79wDi77q
p7VHgbevjG8JtAJM1XXDIj4+R+S+SD2ZfSIBSV3RjUL7XOtZzGyQDcCoaFk1M/Gb
uggTa5Jd+TkrnfbED72QAYtkxMRnol4eqpeyxMS/yn88SF2WwRcvT8Ug/q9R3SfC
qxboJpSwiQ4MOP0So3/TZnTq4IQVUPANVkHVR7R4Vep9x9GgVdqKnFdeGgHWJICX
x+L1SfE4pvuauzy3p7DHeA0nYO5cia8+OYHzcO+2Va0VnshDw/yInqW0IxAyw0JR
T0L4VRgSKgOvzdYGPBOSRSGdKqn4FuCSMfjkzfyYk7GgHvs7OoJ5DOk83eQmXxPL
F+ixiUwraGmqC92PWPxfNhIGpZcghxSwOntsECfkGWmuoW+iDiwFIg+2f2Eu82q6
GWgYspg10t9fmV7MuLD5aAgU11lMl3XQF6MeHtrTZQLXspMNRLDDL74ekFDhDlZ3
7XMgRagZ20F2gxARJ12lnHZlMlxtVjYPFouKKj+Az7aFbGT7YCiJ3emHNzywRD9W
r+m3kf9SmF7IUk+5BHN+VylzRhE23K/iYpioYkeqZAtFz5fQM9TsTE0b/p8C7UKG
cuPl1jHlhoP23NI16YUkkndaBbXTbPsSRCggmfUSK6PTP3H/PuhsQiKUx/0ZOK3S
Q98nv0baPAW+GuK44EMNz/Qias6q2rjEeNgNhZtVfoy/JPHxVi4rnEA5hEX2XbR5
epvnmy+QtsJLhktkUUeQom+fWfnxvJcaboNYiADImOwu/v/WZXV1dqCW/sK7hgEe
wsbQsj33YCYlgiVjC9jLy3BPE//PBgm6pOesWjHlSc344v9mRvXJ/+a3S9GTGeNv
HP1A2GJdhf9vzBUqcfVBlS1P16V2Wg8bNjM+M4xwLd7PC9meMOkQ23lIwpHqIVRu
jCYiSqNNi0euZdt9Eco6yFneAy3IMcqfL5AvJltFamJI6yGCzKasbt9TLThBrB4V
Eq3/CSjNpHy5WGdzdVYIW3pddQ59WahunlregwMs/IFThhPzwpewTKl4e/qpfNJ1
iNY2qLJLHm2/u5tWsblyqdXZ7zoja2yf8JvoTrCI/+Z98uAZgonmLCus3YIaT3FY
dSFnqtMBYhWY9y8wJsHxRwWWiupKcCSUlEEbqVsn76WEXpcfiZVcpLN420KN5X38
9ck8DtNOCDY4vnyD9ixBSblqe/gCcO56aKM1t7NqOyuZy19V1s2t/2Yn8GSttipW
T1mjvRdF+rDTCyf4H/vOfTaUQ5uPhKFVd7Ndxb4S+O/low1KDKNaGUFVxK8M2od5
KBsrEr4mx3jnO2ZRDwnSSlPrMozOayZWXF9KyxEqEIzdGKSkEtD+vOnfEXJswdO6
kOleYxai6WEOQbqE0avvxe8UQD2yhnKQ9/rY2Smbwf72aoJsYfhZnpg42g10wf5e
GFMxnNsHNtqH3+x3FKMqTyJVJUjACeCHkdWJsfoulSE0BHYhntqyS+90Mhkknorl
aZJIDgfBF7fkmG8YUshYrWgBpv4AOZCrCzv7fgTln+S1qGRyHJUDHwHbcS94/Y/3
RnPxyW8fRVBB5qTmZ/HLT6w+yLjOA1O92lAIEOFsFHVPnKArthYWX7k4VsC1sr+X
9GA1+AwBXSZs5Ce4peKG4B+1/THCea9kR65FvMJNAzDqniZ8IvpYQ+UEQUd0WZHQ
7VcIRYCqDaMOdzXWBtCC6H79wh8RhPJYwp2J2otftxEHrC3VbJN/INlxPttA2f/m
msQwa0kMvNfOQKkCf6YhxuwGoFap0z2eDQmVsjKlCAglUEF1kqjuOstCikhfm+9p
vxh2L/03fhJq9cVmOCQWoXi5jKCmbamqLh+Dh8MDS4gIFRCqrmrEWyUDVMszGLUq
OQA9AuKASrBvQORDlgs8Hwg+IsmPnfMAfu1XpvdpOau1DcZh7Ss/YvHlUCjTHPLS
bKFgCupxRjZuHScHKJH3sKZ7oIv30jNNFl0gf8OvPd9wTqyy/0PJP6/N4t3P/xXf
7YmV3BjIrCVJ5Pk1qCXSeQxuqLZehf/nJbi3fjKkjtpHXcdIYpmoSlAf1Gn1hpXa
c5K9CJMc5W68A9195NBI1+yEvPdpjbuTfmiqFj6gGjbBc3l/Uj8f6ewVbEEbJkh/
WebnVkHTojadehN0QSpaj4cRa0YW4aaWiOyd2mFThGZ071Owbp2ytSkTn8BoYoVr
gSBnTEdYNh48V1+vlLsebEn4OEHx91Ju7JAedlgvStTtTje8w7LkvOouXMq5ad7Z
Zft0zHAqrH1ukkUMzo4mlIb+Uy4g/+SKtTOOGisEGTeymkKtb7OfQWo2iPd8cFca
Mor+WrTZsOEa+rjCqJpzBwZJzrjPNoIwGKuMsiVWqc1hf7yYSz6EJoA05T62vusI
sfP17/JNIf7nTDAlcJwnQmEELmlCN2nYVIzyTQJLIJqDMWMP3D2/gjPmcROpTU4w
m1fn+HTfxKhlkPUaTCd129aMOeuvGyg23Cn5L5TglRsXy/4SQx5B34fB7TE8dLHa
FuwoyYSgxf05qbIH5QhKqmT/rAuvhXX1h+BVOUPUmwwZ2aS2sJGuJhEXaXY/uYjB
5WV8yzSzigdEBzFLjpfJVxJP0AW/wNjjMMhE9YydtoAKOeE4ni1SD6Yjt0WwBNBw
rWNDuOI8cFjGXEXRqSs1iMsucegVlGe7GFZ3pn6sotdCFPvvyg/u6/YKHXBXvlm7
0sHVWeeECRXG5OaJxC6x2tszQ8gxFBD+XLVGVOdBAJl42vohM+sySDszptl98v/5
zEmTArUkdMw/SxNfgmDm/35lmkPy8KN47aMk4dSAkUZgWF/VKlRgXoXY3MVhwmGn
ep2JdWpexqck0GHea/gu2i3LRX4w5E3eEzWjkk7XE+0ASXuQt4FuihOREjjhxERH
fLzZKdCACbGdxEAMrKJT0q8UgsiIJHP5sCr9H4gAyXYqAAK9xIJhZ8EA+6lStlWb
aTSOjXMp5Aql2n/MbpDVYWi+yF+NuAaZ3IUKZUXRitParIhxbuZ9CuoDPaavCo2t
MM1wHduCj5cPfVTUmNyIAh2Wfl6/oIDpDBfysl4+J4z3pGdb6uVxup1Ktecb+N7s
1lAngnRdQRoGRHamIlLdwonE8PPcWS3SEtFCVIhi2MB4FXWJ8pnSphhhBxMGyZr2
lUe3bSB+le0s5aH5oDw6RO1xN49oMNdZkqjzJNutJv+D02bkAasAgYDzAuvlzzE5
LfuB8dgNYHO/bZujTEZiEdaT8t0sTicDfIwr36SR4sMJzKP15mOlV7AbUtLJzvHM
UqV//BZdq+mBNvNTED+lrCvpfMDBsTE5hp8i+dRbUmaDMd42FcoJaB1ezgpHoSh6
Z5Ou8BWThL2eaDR5zzxaSZQ8HwGaoBFiWLL6mNFN0BBxWJubbkf4jDuUD8jmj4US
jtxsQ17cLCw7w/SqIkpLC+odeYTxxRFxzhipPqVSjOeUC01Zx8G3P8dK3HT/PKjA
dTxieSwNznYBvnyBa5js7DxkRBdWNkaqnwvuufOUZY/DONX7IAbYeSUclZCDIfGE
H/pxmNdzyV9ajXlSK9oEtvWaIxhThRjvbDTuq/rbITlmRsz+lIVcAewK6qsBjqS9
OA1yMqtpN5euBjREv903/bucJUAR8Cbwql8Nx5OknNFcLwSIFw3lj3n0Ma8WtZWl
sGkRNDlZan9IPyP6s7KEV6H4Z9Z/XCIEzwAXIaJDA5t1PytsZZj2Yyl2X+9ePKBu
FuidtxYoYCcebRRRTrWvuzNpLkDq9f5yq8Jmd9zaObb4si3/1VNnEZI2HufzpePi
5rS1DHACR2mX0DJRXbzVWpCKYkVLwJ5HurMmQq1jlEu7qTozDUSvp7/E1qMqN/jD
fvQDjdP8Acx/ofRtSiMsDcmV/TDDmqLluUsQAPAf09yGkoTVUqF6NE6Q7xAvW6Zd
afu69zL60UJLFTPyRTx3uhL00Ov631YPu4pBQbvql4E0bYcoG4ghs2J8CvgCO1Sz
x7n+G+bM/HiOxpZVYvMaWG4jyVJTDCxNCgnqAzq8OpJpcZk5xBrVaH5Cgw8q9Hc2
tL6WqYgVBIXHORUmsyEuQ8AYPV7LQ91TKAfiabmtjcin8wC/MvrYcI0xQoJdRx4z
IbagfKZA2VBomw8J3+0bPRxvh+frdM4pPEDjQ+cWXippVxH+EZ9s9FeIjAME0lbK
+4PmBsKwZRgjP/q25GsdlIZ9O25QKV2AEYrSVmBolo5rKDJRYzihlzPdkKEV34wV
B2+26sqSFw8usrAgZsAeZRodQOy/1XD/V1NE+2DulgvQFUEav8Qn+z3HW6EKi465
ceeLYHnqZazgdgewgvYdAvg/YZDR4acQaNJh3pWmLu9wB/RJ3StwD40zgK/0nCSX
gYrib4TBdAYeAIDYO545Pb/4MthVdieVu6KKVXgWfp2FPZK0EIwWqeJoRmA72lQQ
4EVmqpvKLOMdnEPftkIJ5vXcEUB3VKxq3UggdqY5VqkVazjRIm/K662jNK+T2Ww7
Z8hP/DeOeZACKX3ljeq99r350T0XjB1dDhPtxZhAhxmlu9k2NFNFDXuycwJ21GXQ
fa3XyETXzDEnFdlXRAzmv1ie9YmZdk78m94RE+WwsES/rZ0JXcJECZPdtpeeKSRU
d5iXpxgzoEgN88DXeP8mZIa7Fv3vs8n/LPg4zZKsIbfZL4/0IHPbQQ+TpeKiHYsF
rrNqCAvZKyeassGkX5d/kyl8R+m4xiqE46Xmy+xdcyqaw7lyHTvyyozCDSGe5kNJ
yn/wVPnsZtKVe1U+otR/fcmjZi3zH1Y2t/hkKXewzDCrw8BhB5/aTA9mZNlUQV51
2Dg0CrsOFoM0o6WtxUaxD2gCeVnWyLdihctxcJAO08OA63OHd5ompNRV85amJehZ
/1KYMP19qk7KN4acqot64Yx5AzvDwohc4UIGA6PJoUtSkxGQeqryYrO+P7NaIL24
HVwFgpU5S5IN9y0gUaRfHDba3bY045c9QpvBJjV0Q2I3txhepDN4ueqUG7w5cQDx
RONa6iWbq6OY7CcQJvjcU8Wl5GF2NSffLb0HShkgN3seLTSBaRrdz1zDL0sR19ny
HqyCFES+geykIzwRLFa5gG8kGThq+B/iZMb/Jm5sD7HySdoJq0/xshs7ciaTFeTR
o+aHZk+/ehiyFamJ0v5xCWKSaTny5hchWp8Fol3meoVVKWJ06f8OpHexeBmLHIo2
3XnqQUZ9RIAgW7tNeIdTfbZcZnLnLZGHLC0LrIqM6yr6DOwNboR17XYOZX1lRaXS
rCqWiMcissh9LJUBmWrDZ4e1I8/ZyS3QkLsRga7T90T0Qs8GixTiKOayYG6yqsVf
Uhn3GEmm7e62LW8eLBFuOfqs5PvCSLyl2131atplDQ8pu59ClQ8pmc2xGDMCw7/Z
rPFr9fFEJ3aFdV5amIFCxriBm6enEOBOZUAhvXjZN8esNDbSRX8r/M5pQ4U/AiGm
k0z4XUL9pI0vi20KMfC6QwNdJYWJoePrSSpATkoAJ9rsCyWg9DySaOGHJmNiqzF+
zD8yZiN06OttFuzw9CSyIcdnGyRDpceQ0wBI1ArBDEd0wugLXaC1oHFPOkxuGzOM
yvlRkMivGno4sHwC3rMGVn1CcSZwQ5YhMQlu6cI7voPhlY7xVJBkw2e6mo9HWpLV
f8x001yEPMcj2ar0lVrfwEf8UnmvUW4IMahDeN+vVXvEl8/B12PPBENuvKV+DX0R
EoxV5Ab5Si1fwgmnJeGJR6PYhttM6d/eCXhA+xSr34g5v8zWxGGml9SmEiPx+tuL
I2thfWSnCpugx8PcG+nlvfslub9EKEsLimTm7D71PkT0oZ9RsGd9x11qRlCWFkDQ
MzUHyq+Kv+hbLnGnA+mPIUDGzQZChzqQQbEyBWGjfWafN8nVQq+rq6U8nZ+1oqI6
XP2TM2X25/luyy/sM2SFzYFcJYBqpB80Q1euaXQLPdUIC5yCb/YNuW55vPu+OB82
cYvl2kHJgjTYi4ZR0iSDSmEMKwTO3SBwMusGheSGPmWpBboxI191rIBbT8iwnoDy
1B2V0+taP5sESOS08Hs5e9d0UZMxd+ncC9A2WZ2Tj33QfIZyx9VtGV//oAfy4X5/
S897x9fvCZ2Vkfxn1bZ7BEtWQwyA27EtOcvd2/YhYc58cKnt8RzMpmJOK0fSc0fL
f3yeNGAXaO2rjum5NcQt+KyV8n/b/PSQjx9G6LhEUQEidfSdTmsbWAQ6+1CiV67E
Vp3i75t2GkPrHx+fKE+rwEIz2A+yoKYjGXeMgFDCo9xhXbTLjARpTCRg8UkRLi4M
CNspi6iNfbL0LfeAdtepqDl8LgqGwgA1J6ROsNaPRh2FpyM+CDiN3ze/juA9CiMX
3RB41dka0oM9rB9LPPqJbeYnfGimm9mfRfCXLScojV/8vMOTWOxmpPvq1XTeiP49
VYghXtq/9ZRBEdw43CsyR34yHaPZ2NXdbwt742W+eYtHtgGkDW9hlBlstZ+TdJwe
E71oy+Amk9/FoQeRhz7ZgJlEYq14+dntJbvcxOdCe3kW/8Pe8eRDUNQ/y17XHgeE
HSegmwN6BS12Hy2JlQ+6+ArE4Xp/RBvsLOGM6riuJE3whC4OK5fLcVwfCCMKpHb1
tOq5JIdhN4mSg/6tZbTQa14lkvFBjcxX9G8JKMvglD0VqbaPGUlUALY1gJfbdpJ9
HonDtv/jbtTmr7PD1ToB/oZOtO6f+g5rGbDVvMHO1gudEoBKnWsz59dqPTvTrDhQ
zHoqSgEV7AJPx1Gs6n6DdPGo0J74wgLqfwJCg+1EolD/4svOsRIyPUKbKaMUFA/i
ueBQxDd/cX5eXv2OzSIFi7clhwZmZ/mWls1oO2bwwpKM3PUrANGaZpHR+eNZp73A
UWXnAK0EJ8JUCBuXNvvaQoCio/PTzo1e3/e/KlCNgGHBqHkZq5imMHTUWYhJ0QAH
kHQp82YZUpkMf4i1XmMP59m+oaLeaPNQHk0/xhz48Jea0gRvjRPWG3n58mwSe/Sc
jUyOa+94lDIGMq6szGo+yhjMTyANk+/LFu+4YH7izMW8EQWGnlmYFsqMC0Cot8dO
tyfiVM4kvTESPH1oqpK19hLPkToUMG+P/h/bhHmt8cF/UqnPV8GGWHF7Nhf0EPz4
LkUwrt/JvAyDDgTLPtnJa8lYvu3T1rq+0EFraUc0/2pdrE8d32gT1Xvwd2tV+wkr
yAsTIeYTe9f8F7JUh48l6OLJ51/c9Iw2jEvRXiL/FGnJz+tNzK5jDze15WWnDlYl
UmmxJjGEISz97ZWz0wf20nQ6MCPdjrXCCah6Cpa32qR+tafT94RpKWMXsJcrvUmu
buwlr53FFaCV9+SMnuRzY4vSA/24M2SdbPuMkwiEBK46M74WYOrEAhPZFsfo22Ja
iDwPcitaMQqEoXZR033dxfouk1zLywPhbieBuDtRNdBuYdHzEsbUruKfeK9aowva
NHX24rjEpvgxZcMwG3NAP24wOWxv+/Y19loX6HMnwsPJ3gJHKwIFkcoUSEErz03T
mjLgoJH/04VVzBi1voHchmYIvKBWkYKZn5TngPv1SShNi7I9VdksywFbCKritCm1
MWWcLbbJybD8pQ4mmCe+f/9xQR5qqOGpXQONruJpEMN6SyoWY35UuJbLJTZf3UdU
DJe290Z3aZdT7tx17VHJhTL4fBq9piX8nwyaP2JiaFG8414Trs0sdrt/OGQY/lC4
ontqcS9nL0hHY5atdKRttXo+juD9VcDnylzzF0hJQxo7pdkN/xBGILXLGD2d7Mqc
NerOLYQSOSQDR36j3uQJKL6dRj+WdKsGkKNVrHXUID6/fEJjfFlV/M2ksl3u0NsH
9jPSrTnpWY+jaWLFTrFCk1YdxP9n3LZdoNB3YGHVGXE5htuQ1WG3Q1Y3+RVB4FZW
5j/z/IZPEtZHXkT3MDz6XMaYrtzLnZ0/gefUHyufJCDux/EC00JKpUTNgoW7R3sz
fZJRhC+7P80pBcEGUKZ4JPJPiKfgyIp+PIf1VzigqulEhCfM+hOXzZjCGb9kWcf1
cD1rkZ7lbAIWXqNikhNBqNIyuN9ZkJTIADfm5NgsDvscjWPqchGjfHeBEfZhcuhY
V/6ePhmT8PYVH+cy1YKgIqNhphfCnU3UNrEsFeibKsrfrm/dVmcjqo3ajy8ufgDd
RRbYg9NwGD9SH2Iw+vXtudIl+1E4ZGQodviUEhXt445EnR6KIyn/lq9DuWIu92BV
k7oWDsQa6vSNxTLKAsHF8MtExGSlfBGsC93tntCDKo4zj8nxTYppCebxxGCl9t54
DGPj+IDoTDbrFNERuFK0ui0m+lW+RuxMPvFnTDCvycedj2Ka8sSnnFaai1eIwEC3
tMx+PAZYsH6BcirBQHgaTc/wmfUNTVNNBwnmfkpMHLcZdABMy0JhC/mP2cJEH+lC
ROvV1ncbt5IJvvIjKVLxQVfdyYHAlD26tX2uOVaTPqydpVsj0Eo8UeRzUAJpsaso
f1ODIfOd2DqvfsUXPPcEFCKmaH6D5ve+SnBuSqNbHmP+ttpqKicimZvUdqjaRDnV
PaPbfHA/cB/C0L+XfEWB/KQ9e+DeaGWdYD/KXDjokoUhJsMKUAA2nlCvhwM0B5Bg
1ZIbKyAiJqfnpL25y6Z43lLi5xNwkNfq9otR6dkEOcqG4cgqeeFbD+7zFqOEBNon
Ci4JdAHfZwZRtSSKvx01N77oZnqaCsfDdz7Wg523BWwdXX48FXls+Y+QzyQmrTTp
3IItb17bi5MYtg4gddza94d9Yu10JaF6LWMLCsmSK4XGUFRc6ow90rah/Bm0fttm
q+Po31lM1lrZVwV/pmtU7qFlUmktcjZj9ZV6QpzfVWb6ARXTdKvrO1QPp20wG0tf
cAq4t2MQhpoG0PNirT7MnBs9GCW1j3Ora7sbfZURHho+t5Cp7Tj0rd/GDkZ7gnJu
tsh+JXy1MygkO64HONNT2RIr6hPP7IhWhpQoRM7InFktxjuWAppJ44ckg4UJog6B
4Hnls2YZznc9XW8KSZWkUaY4dEJHjfcJBwYXxpoWap5ZNZ+q9F7OKKady6tfmKcO
7jj0eefWpsIqH2cQSmleu+haxoJbxnpDhoiwwhtKUjSxhqwvTBEpXBq/GDfeuXy0
fOFsVuzy0vHxjdi6eJUVQQ24DG4+Vwk6vSu9CPlcyHXOC4jvu/HUKPVITess2G8E
I05wnaZuMOwrSCPvlgFv6EKgQtIe9hLPZVfNHbKve610Lv8a4K59+Hi1R9xDY8rf
ZT+Shpgg3i5gnKUgYa6n3thqE0LD8ZlpDos0MDvOr54Mc7Pmmi6jj2BwbRq/tctV
FJJ8EZQ8O5SJ8x3d6pIMMnZr5ibfJG+5s6TnqdBINv2LrFbtGhQEndc7lWry0pUy
hvZ20Xv+VOA98RstHjaWN4V1mV7DgVyjBVrdDyLDpBUW+tHKcXmQ0qKQUX+GaEa7
YSOflwTSn07h/uwQw7bmJvaX+65psJemu+x1VL+oKm59YbDS3caYT9MzFBTGe9w9
jY/b1Xdy5tgV1cI8mI3q5/hkd4gLHCK7+iH2iYt9FsXjjxrXkYiFWPJvyxYOT2aW
7KWT03Bbn8JtG2u02C6JDREB3zVmGmnxu4YcIOsvNWRZCuUvoJ/bGeCnSZTEW+i7
01Hu6TnelaiZxkKQkBOIb90Z1rdCNhlbi1K92idrAEyHzAeE+y7oiCIlRGEV40mH
64V5VTqTzjBysa24yYGNH6Tw/GM7+aw3slt0GEgkDAM0IFx0LNPIHAg3AgYT+F/l
I3SfPqcvHhgiTGA5LFrPV/NPZevQwlzzSmop0eyehR0CzLNvRsCI7pIyfZOBMqRg
DrpoM5A64Nq2lE0rZ+k77I3EaQbT3NAVffMlKaw0pRA1xh3yX6GntkHNh3WAOj2K
2J8oLl28zTls3D0OlH+Vyz/m2+SJMfbKgRNtD6LZTfCP8qn6+3LZzgTbJMh+UwmT
L+wHNTTzYfOAGs0ImVDXzNpRpw8VG0PQ5QiS/PYzgKtlvKmNpNqquG2yCVCOYCCY
/QsrLfzYMgYn9dBNY+z5+zL/Ci0NZMc+zRdORHcuvGA6f7F1oOmd60JucbNnjSXk
N+pMsLMH+ZvzoPnbRAkF6rrraIyYI7HgNs0euIZUARow7EXd5yW8HCRhtmqFATnO
r1KN8g2bbfW33X0a90VXYH+nlaFxNNxr7QqbJHr+s9PHnwtriuI252dIuG5cVvxj
T/JNs6yITRONAj4pYhn+xITo+XR8/teHenpcWkrvx4SGOwZU6YoUwG/gnL5IrO0X
2t+Hs6pDIRd6QFE5n2enM7AiebfrnLoYPNUVr+9hOeGiL2rZ+vp/HnJmf9z0+scH
PIP/DiLykNgLEwCBk+C3PDpSYfGriouH1F7LtXEU+VEiADubf56KNqYUAB8BfIt8
+wM5L+J7ubtmnxfzvmq/gKnNPkbHhhdNTYy+2jRyZr1bEFXF/8BId/5aNI4RuPwr
xKtLefwSPqkqX95OcLD3GV2pIUiuKjzR/3tErvkynT4vnD4UA6Ush738ByZKA3TB
rilSQQscW7ndGJXz8DY0dt5Zny81AiUD+21bB1vKy0bed6rekVDUD3zK+eKPisco
FU6H0KGd3FtzhpzuXwANhHv21UozYiNFuOY7bQRYt8ma33MPIEObilha4oHEgRVN
n6MQkGP5PiPltkmpQmpq7kB6o25qFntEPa1v5G1dqgtgqZIWdLdeeXHk+d3YtFS2
0uO/K5vOA5SANIh6cn+jm1LFhi+awu5jPgvhvrdxcacjSiQ82XU0xMuLr1cfKYKO
jApGEqQNplg1qXUUTfXBHPufMvlw4PcKdCsCVYoHOoDVdoY2TTQ7N0qyDwIunkM6
iYoVmmgYjtntoxP0/TR4I7sird3lFXs5QBZWcAN/mdI6LhhueMAskDtZ7aMti2Vv
jtJJNoBJX3nYX5TCo1by0/m1TDYCrMI6lsv1SiikmYbuayQeJacii5Fb34AWX8yF
1jv/tXs/AWjkbJruX+KtnssZDpsTpRbix0ivqvR570m6n6/i4atS6Xz7jdGWjmH4
b5jct5ss6kVtV90hsYGZaaIRHY+sR3bva9M2b8IfSYjOc8c4KS1BvTzKToG7CNfV
Ogql9jHOBhR5KiMD6FBTOiN9SMFViga7/45aI7NafqEGyPweJ4NDCAzmvehRebPy
K9L44IGQhXBbkSPIJLey5YXIZrGUE+wKA5hgwyKcedlkqi3otlmmn/oWdeDC88zF
BJECHPLKbrruwBf94Mw8HhPDd92//DbbNPUdt5XAOnCxAKxwXom8dUC/M97n2Tof
Xw++YsRKgOcSfS74N6dQxvzyFcvw8md6Sli98yr0zT8EFR1t8pirC6yFIkIjdNaI
E0y1aLFpNDqQIZ+9D23U+Fl5GvfoJHNNAxPEfldAQLsAxHtK4Dozzr/m7D7h14np
bxgEPxN7K28dH20e2GaFZxa3S4uAavyCFf6yjj/K5UQUDFOZ5iWGfLeLX2hd/Jr3
ChaWfXKYRl3z5vNNoaam5IfZlpLLL3aP9x0dzryao+2FRLppkS/qaWYUflR4dav5
75vWYIJ3AynfGW1I1kyCwkSYOVWgM2LJvVz6ngBIwhpOhd2s7dSuvayyptWLRNqd
+FH+Z8OYeB393/saMyyyeb1n+/GmKgUcUdDdjfUl+Dj6g1cNnCPSraP0w1qXWMjf
Go00XDY5DuESJlw7Vj+AbRjBYWDrw2SMTB97u2nlhgwNEB/wYf/RhgxdY9IK+3qn
tFrmdk7Xp1SCNPUU2gKaxXwfCiUj61b0Lp2p7rio+dL0vQPnQmquGxyEeLgyDMEv
AH4GWDriiQFMqe5tQAIrGqz0TYWrc88M5FfBF3tGSXMPw3poLKCUck48Ujr/6z/V
V9n11MLBXt8fdvJns67b1p9AiNkqqWtFK2FCbLIt+KpWzqq7WCQ11MJC93BFd/aq
9ikQWxNmYKditIB9/J6Xjd1iEXYsPrTHgZ+tkQNWvLcA2sw0DB5t2xz9df6cJqJZ
faT19NU/OdkgbJPJ5W+kMpwHOvov8REOqqXU3G88qE3UOaGEFi0FWEkm0VR/7wo+
fn2G2y12t5xgqUdu3H8qlpjD5jyMd5ZChRFwVq36tRBDUs2F9ZzgHnHqbPVoMeXY

`pragma protect end_protected
