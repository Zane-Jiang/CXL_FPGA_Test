// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
n3jYODM3uIZeB+tbmzWfZoBxtMvcpvBK8pBaY5xBNwXzBf7zWuQ0jfnL935O39JN+XuXxisRHgSB
vQ4VtqsflgaXAzSe5xONLDRJfmSvZb7UDNHvM6POX7zGKDOg33bkzp/+XmS8iKvJ7mz4j3rLSuJD
XRWQmTwS9GWdApzQ8hcsjSP7dV5isFlC5f1hcLsQvFlnBorN77itjHZoOUSUMpML2RbTD0sft6jx
8UGYVTVVIc6XSrYaIjlUcSrzIyu9EarA41J8riJeZSMHKiLVb/PX/Z8cvaCWohoQsZ1xEM5p9p3H
IVwgl8CtsrNw//dJSd8soDxtW50JoNCry0RNRw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 26496)
vJYSPmwWODexY4xV/ZeVzIXNyPgS14pU8DKkkKRmpyOrQmLnNChQLicPj8zF8Q4D1SOax8lZ1m5Z
/zF+uIfpOTBR0HPqVcC9QsNqa7TohBeKnyiCkV4zDheuX1jIUReMCIRlIELeGhKS+5WhBuYZkSIC
atmBIgulPP6cZ37jndOhENKZEpf3xByMZr549q7dbQXIy4jhMr0jR7jUYCD2QUS4ckpjukpbQXpt
MWxhA6Wd3+ofymmnQqH63eEpnUWgmbZYlMm8RILkV5rJwI6dxAEOY9Jm7+VgEke+3Xp83TS9kp+j
l2A9U0UnS+LIYYv5Djj0N5gkY5q3P+dz+Z6fJgAN0efm9egcbR92gMRnX+mm595Za7kPMrh5Z8s4
Nk0NptsDMYcDZ0xH9W9VoWTstfQwwcsSGZVQu1awB2g/B8+ap6t1TVkEjYjUa/Jan73384BRmFDC
tAsnukII41pCyodbY7NazUfSii4Lx/LpwDljxoJ7vgfB9qkdhLtVhv0/X1JP0OPsd3Fz4QaqZxS1
D5TZuFKiJo/+gjMIPQ0PWvlFhJBMFxw6Z0lpXd8Kj8EHzgAo17HHBNx50WCHjuw1ZquIyg+6jl99
J7AMRIVxAyiyYEWhZFGCmBgdo9QiY2M4l6DFAUkkcW5qPrWQoduTSfKTR7cnXPv1R6P1ccVbG5wo
HOdN2cSbQfWabiPy21pCnlS3BlDJw7DDslq1GScf8Iduvz9ZlyHVySgc5zwC4xCZYFdnnUz5WWyc
G1b8O4PSb4iHyq/N5vph1WU1JvGkB5D/nDaHuD3GEuTMsMudjOGCOegzDZ86Mb4Mr0++8BLTahF4
N2rpovqxkDpNumc17ACf6vLRD+8x/fBxHdx9OtxB8EY7SdoqtEqolS+yMZcKAbuEb8TgtqlQ5SQf
nXNUPvTw9EJFfHLl9lB3E9f72JjYG+/N+4bxWB/ejtbvRDHZ4mDHkGj/ne+U1h0TOwzu5GBKohYG
MVLMh/jCdQ5eLTnQYQefWfiWgHq4jgvp3RrkMRbgWdDp81+v4Ek+CxKGlVNTgaia6vqlAjfzLU7U
mfIM5Ly5OfCA6RqeEyDmO+RBxcAxIGSieBIRzJlriychP6+JAUtFxDxlC54vZIFjqUHx2bOQC2ML
J9gb41ET/JaFOSfM80tPO4uWBdaZJWDLQdug7ahiN2Q+GCvKKZEEIe4YF6aVKIZ77Jz67hJwCrSA
wqAgaukEnwoZDb/hZYVe5olRvkS+a/Hvum+KbcKnh0tPdeUpr5U3aS31qu/hDy5vx3B+g/DcWbYI
fBC5wETIpR3PBTAjBIFJ6r3fPWaaXkvOIPzEXjLKKBYctK6AYjlBHSnheJKyS7kvj0XL/knexK99
AjviP/H2fHeMGXIwZI6EcZk1pO53GToUMPlhZeVkPrzHtqbqaqpzYvz6eop2r5KfDRVfF7NUFw+O
+TIop4MiSTWNVT4CV7hCowkvIcdnS+yPgDsXf4ZQbXf9aFJRV6yBqVDhc5qJYuko7hwToMXB+TQ6
zzxoE2Jxwq+Y9bkymS1AJVh6onqds6W/FSFL2ioIGpoGxME5T4z3arPTnR4jfjZwA00m2dy+OovG
VL1QWdJG270M66sidAQfikSmpNImPmwjvSRgxSPZ8cRogKYe3Jq9P1eYz7EaXRExtAEjAFlA1cF8
r/aK5Ah7cdxWN+9gSZ+wlO8Ig9JsPGDVkIQ0yxKg3gRHhfEL6Xg4FEu3G+fKIKKn66PiDM7Z3H69
dWP4pAO64Cc3Jslu+7rQ+DsAe3sBP4pCV1/rwrbeG+O9lH+rp/NdSMoe29Ug+FWoSbhYtMUH/CNI
wWh9nDz4iaF8fGvZPhi1qcIuIXbQrvTK+xli9QY6DAvVLoXBXV1BnNbcgpi/CzNNTl4gqrllU/QN
bV4k48t/wl2/8vpHdA2O56TnKDNwUUPZJ5NC5Dyy8FMBPcnzOww/SWURYX/LDkqD8398GePU5Yhc
4mXj/571i4PoK1jwl7tBvjry3HjR2+Y3jt0aRixpRMGSKG9KieuDaKMCSDViICVCu/waoD1/F12l
UkRXf2ofSe5UHhy3EVCO+vZs7J7ow/4P9OhLzjOQOiKoOH6FHExGp1i1U1OKWPxp+fd643/FxJCy
a+nnVjH8ElcOdLo05hJnN7D2vaheNL6tp3hdV/RrB/C//TWTy0tfF0UHJ1AhPkqeB1gLAK1FIozD
H2J74+nZzdAvKrokfwkX0yyBNK2GI1uv9wx13GfZeZVZVcAAJrSTJPxcNmsdZTnEsqR3hfpRBT9O
QKsl5rqQYnwkS1jr50vv20vblqyfgdEOJ+lQyqwqt6jSUk0qHIe3+cO7kMf4/c0Ne6KtznSbQyNo
9MjzxmJc6ZZx3sZwEwVd5lh/CVGml6J/Kc/rv72fWwlDo7DXqMhw/+bYMmXs6sT7qwL3k0QFLD5K
EKZlJzrFEmfJ7TpGrzEXJmO/Oo3ljCpW9Zp77dZH8h4jGROd/8qGIHs798Y09MXk9hsxE0XSy5gS
6Yg58dv2nmQ7i5Ivi3yt9kneoO3+J0RWbPUY8jrEJI52cMx9kqyta6Zipa151UrtXiVlo/5CVsuJ
RCsO2jd8gKFaBCi8o3CdieHqaPfq+18ppVwCFjTf7pvklSadzhHrPRA7bG4qgGdXU3Ra3q0LTzdT
j9N/F2ukw+wcu0Y+4oOsI1geuU/UL6u0uT2A7ZOXQATiwcE+b/o/ZQvTa7uPd2s2XuvroP3ilSlA
tGpBVSzKPtCTJ53HK1RK8UjIPutvEbn0hEnoKcWcxzCm0owmTPmwkxE5Q/fwLqNI6vPGVRFV0pyk
lmpDFJ8ph8NJ/bxjPGj3YeMtqaBnA68nC5I1TEssTpjq/fYO8fIDrCCm5WOgqsupokG9Ww7Yi+Fh
1h6Sb1Z3T+hKMl88dCn/tDv4VT9hqNs2lqnWfbSf1q+zcMj7Fefh12FfBNFxZoajwMAj/MS5yVog
RvFjauIYmF7Y3gLnyppw0pBu5A5pKiWGwvWmLK4BdH51QS1Lm//iXv5dzReOZ49nmhvZvc4aAkFJ
c5N5ePCSS7nw6+lZVd4OfepMPKlQ+BDDXC7HO2cjG1u6gYqyVg6VZ+ILCwJeiPyMtJUbs0D4FimV
/YQJyI66I7dWv5i8R5bAAktl4rjI5RZSLKVOJ6G08E0wuENfDcuyJHij4dOhjWjUajHcGe6T2/NZ
swuo87e+ff4ELP/lEdfHyTXwxjMUaE51WmpqXKUlHu3QJmvM86BslYLAgt36gSqpddPFeSZ2iUrQ
3vaZD/4rb20i/hsu8EaXBdYXUmgAUhGWN+J7RXH725NdEtL05p2EjDKuBtefQdBJ1BMxr1O80Enn
/0pXjalfw0Twzugu3yHaiaZKSVpKDkyuBUe7H88phohOb5j6/O0niDt9dHgusXLDNpmfNWGxb8h1
gTXup0zawoge3mHR/zERStRvroAWbM4rmBzQmewgBRALukMyvN8giOyAqvAQ+OGq07szgbjNWYkk
ZUrNzIfTus7Wh1JmIjvg1duQ+q1CZPJrmkg6OIy6orx52xvSJtB/3i7Bx+2BH8gVaY1p0q1Ibxap
XYWNp4uB99Od+FjvaH0Fv7gIf2DbxkP24xHRWWF2cSxcrMzh6RZCW86QMVlT6X9BhjdGnPyGXMH7
sAi+xJ26tNaNOv2caT0NdALqCMNcIQprKkFkzIj1fgPswpelOXojYePMTQiWw3Wf0Z5nNtrO50BY
3+9rAtGCt9neKIozIsN7DDFt6uwnU8Bkrf18jVVqbZCFQ0McCSJeD01zRZrC3o44waBwI6jjuhpF
3iAg7+lzZhU3lt4QHgj0AodUDmQYWBDxxpxdiqFiY5IxRToHzI9vVXvPLRjWV9ngpgPhipSLAge0
jQqd/yITuPsCYKVFxL6G071jZwZqrMCKKDmwZkf6PPItqQ6nSEcbuqsXQMHKKzZcbnkq/IUfU9fN
bwxtz7FKtf8azXV7W9SPrARlGnSSY2+H8VH1IVWlIYS7QB8aQ96bd67oECuf7aEav/BOqkHz9gqD
edx8JlrqIZoDleCLkJUuG7uHhghD4O5c8swjVlCzyEewR2T3fZ503ugy7k2OQxsRkqI0OBikeKjU
o9CH2yHjspJrjET0XDWZ0P+hKj4mI4tgXD7hd8SLDgoY9weg/k9Rkkcoz6ozlKpSjq8EmXDQ30/s
jTqT+rCWmmGBLbyMC23x+iZgYxgaiWpORMEtUqNLM+jRSP2NenZfT+W6Yd8w89++9S8Q1lOrBzQm
I5cfOWLFQULr4C9tsQ9RLx+7KB4IezOzhzPSTXUTZBoMtfoSiH0bfdntqkQrQUFlAWf8GTVA2JOy
K2MZTPDHLv3V7Zr82OaRkuoswg30v2gwLg80y2jvddHlBtaPuPnfKNNHs0+Z6iTHBqFumrq9Ibs+
IuqQEtnjMkBXl3IOgpYPU0Rz+77Ua8+kg1Q5OvV8VBSS19UY2ewAZLK/T5YCHY3NJ9ItlY2h/TKs
FnvrK9zcHoYBO/Se8kSTjNt+OdHVW0xmma/+DNqE06IDpc7xFnlc9Z3Y581tQ19jJXZVhRufru/9
MTehPi4rS5XZ4tWzai1JxsxLiaHqDu3wfUdGly3U8Bih4CZNbTlKnfsJcdzv+cmgfBi9gVoJDbuL
GsdyRqnYTvhih7dx1BUAi21jz3zPdFqgyrsv/X752l7U534KkupWpz+IuV78j2cCmKwWUfpK2V+R
sAR8YFsPN3MiD6k+zISmVCu86G00irl1V0IHq/kIZdVNeSvLkn2ZLgPP8YzOy7AlFcJBgWxOE335
itM0I6/lyvD2GubEDrnDjnLKsowxcVlbqMmjjkB0QIo1rS+hcC3bmE3Cl3pUmUFkqY9WidjtRa9X
Kw++RjXU/B5uR1g8hfPEQgtnu8y1YUmumLG9iNDxIOzVWHIvpDxpjhAuxBPn245T9/vSXHdPSTyD
g1JDT5Yaf75GiwIwYWkfG9gWovc4gpfnDTahQLQKM9gKr914HoMVa6ut4xbV5hu7nMnVAVIrDGTB
AXKlgOkah9ChQJ1g83xh2UzgXEaAvoEMcE/B5RVdYC/IVkVFlM68NBIEG0qM+HDPRK0/5tExVhVz
eVVxH4kvAENeP9NtdJcck7uSPu6ntpNlhBMQAZeWcyfsuwUkfocow+GTkA1qxuA0WIhT98jf2YbQ
yqN+DNrlYyuNdlh45NK+v++YIyOu21tQYSNM9B/gzIp7k93dC/aq2YIHSDpEWsZuUmdHEXTPnNAd
dmaF3I1iATneokWSp1HjIgN6NN9cvqZPw0cwIKb8dEo45J1mcrLVuXpLlqBxSCQVEh0XdXhOsFM0
rOB3RpDhq0w5ce0un8U3iET4m5XpwWXnEsW+9r/pygViEBd9oYwdoEjMg4UjRdH+OHdlLSPBWy7S
YcF3u67OyenpeX5bisHsN4gX2cJ+M/9sMtvLskP6ASY8fTCwEYv12EZg00LWN0yjddjd1Y/hlgg+
+ceJj383GvJLxUcx0YLf+qoyRHVKtzirIqgz35ULL814JEYw2VD69wPHAhuEzY4Q0FL5Qgb/19Pt
17BUHpVX02/GsrHzrgW68MwAHl1en8lsV5OJJxPTL6YoE5vpEWvFNx+LU7IyrWHiQ07ccpOQODFb
+HdYSeG6oEnQ2NBiJXbe8R9T5KJQ59BwgUZIVyyPDeVLnCZwlW0ByM9a0KC1zBa/p0NefCw3FrC+
13g8xP6U5Mt/yR54FyKg9+yac6UNBUCpJoIUrknresLPV3w1+V23s/vnTMjpZcr/Qfh4TR7BKi91
6j2j+V3ut77uhFH1ezRwvP46NQYZ0gteO7D2HVzTZ2eXKnBcmN3ZPCeC++PgCtQelcjMLUgfBbtY
iGrTgT7fTd3NZMY+Q63t+YlLtlzNzPh9S4YOhhD+wq6nFarumq6FNwnVgNn4CuXuLbZXgyPogFUJ
ykdH/ib9EVjG9QhJtd84DqPGIuOvidVDmrD0TapHSWj/cMXOyy94yoPhZzY5ZiG3AtaQrkTOF4Dd
Luz8LfBP4csR+b4LDCczci8bSn8+eUEqifnHkmdJnJYYmDJk8kjOL9OZkZbDQCGUegH1LnAWyqi9
kIHL21vf09OmrR1L/mYTVOa7NdGVJw1J+hFC0uFNl5vSYmGHkibpbgRTx/WLyf4cZAzoPidbcy20
GZgD9S9wQwOfyqzFWEDx6gy29OZ8F52wA7EDZXT0+WmnxeLvpDDCI9ADj9H58vP0kxxifBsf20tj
ex/oyz6cbe/2yBpbRSViUT9b5FvXzeG/9hEL4ch8QOILUvlJHCX3yr8SkvOxQTvLfqHif6MUEhD6
HHypmk7XmBAoskXHITZ+zRD3rFmpYgR10tovzJcjLZAZadZpEeu9CxcBjqTN6iZvvimuU2rrKjuC
TgCcjVaVyEYlOf67baWidCym3ye3+xlLPsn2w0dApW0cxQRCMhMv4l/zByseAvO1Z368ZQBQnSRn
WfYxmP4WMpXRPgHpDXPg9gpiOyci3Q1xeB0otTG+Md+eEmyunM9axcAvgw2g08p16EziBrxVhc8r
qTvp7fYDEor0D8VEzWMcTswPM9qNFLp4mKzYh0KiH+mOT7XkUkEwx1xuL79rGX/A5Tm2Hg3jEvrj
EVlFL2nW9gR4LG9ZHXNl+Jh0BdJgpgwuTeQPyN6QifkHSzLpvPNDjma7/LpI0hrNfjEqMILUl7Id
2TpQQiBkwANxvCJY7DkZFcPG37USdO6m9Oecxtp/P7W7yUvOAZvx8ieyHkv3HWhxy2RDVE+YCOAG
qbKshW3WPpi0zUiIVH6ejgzSmdc4eYvmA5GV35/+1q2uin/Zy/kKGaPHxSlwAyhMh6V08Jpf1Ezy
1bEY5bHfINMV22tU7GeTsYn0UxCKJFg/OK+jZgPF0aTGv+EyU6WeCrU9ngVyXzrYppFvbPGKPtD8
TaU+Xc2uba8zwZDsYoTgkj89GVlnudV/60zheWv5pmFC78zt0v9Az6LOWRyc+ghjj2NYIReu4ztN
r1/v9ThZlCV7G5iCFUc/zZrN4AvKDDNyIlpD+irYvigMRmor5F1Zx7u32bVwaz5BHbcm6qYzQtsk
um4pMu3nao/Dk08mqfw090H2RDdlZww80Sy/RxygdXf7y8XMiyy8iafAg1MT1kZlTCpvLf2smADC
FMJH9hymzLvVAK/enJYLirYT+kakvapwi0cu995/Ac9tG2Y0YcryBPIWgLuVWb2xPiTkRpU12bjQ
jq5PQyr4DZnj+O4Ws5prULTcoIiAAjLX4z4yb0iG2Di109hLs41Np1X/Ua4tZfN0L50sp+vImu6S
bAj+HyCryxtlvpoCds2kvtQuc7dKFadDJqWC+k3Yv2ObzIzv3SAxRug8GBY/vtxxSeUem8ePTNdC
ty2PrDmzaO8Hl24ycb+8ozE8JjMXSLTVdWR3qzoPuTWhuvI9sgLjN9d20Jfx28Om2E900BlwPJX/
v7I39zOpYM3INYgDmKZUwFbGHLDxKNt30wWug9VFgIelqs/ammzp3HQWzAwwd95YJkM6cKgGsjWM
92Dqu2v3lTyOnXf7RiPEg6aVHwYYscPCUYxUxcnZG8wv9y2Gt9acPvv0q6DO+/56Dyx1qnjO1bIM
IquYrMOgmjwWQU4A7ZxBbZV0RNy7vgElOpi4ViWqAgnJ0phhcjkdZ2Nw4Bmh593YpJDiq3+duqRW
3e6HLWHCZsYgkEoJZ10haWvrA2onlqiDqV+r5pn7r6lEXann3LEEB/kELHE6atgfyFFTNCjJY2d0
UeeMWtDczoXnP7C5x4MehlUkDR90ftd0C3btGaCo21SIV3SnFExLHqebYJW/f0A/LSwYmke+jbOX
LOgawhJ8iiArjPGtZLqJvs4QFDC4i7clKTvfCv9pdhw9yfAMigAwwfQ60CusclnnnHWnBp5qC9MF
eAyxWLL1jL9rq2Ynh3IOEp0QNwW4fK6UWTPcPKO4KgyI7nM5LzsAo6MZoGZkndAjjFrN/CnJkL0e
RF1LfoDwa0GNrCGcZ1198r4vvb7338gZ+CjeJXKW/wLMEAGPCc6Wt65CJvCBmI6fueLlO6dm+pD2
a3kJWT9B0fwUkeRbo/X22sEsQAwVy+6kqV03GLshJbpOxrAbNL0Un4QxICr+cG5yE88BxSj0pasM
POJ6nBzplXfVKcMG3uln1DvGffsJzNlww2+M9ebo3cG1U/eWS59N/QC+usj3VN6NkFZJmu5Vnkez
NZeAPOCkgdZTtFk/+d8UcJ9tHxQGU3wAKldAJug03wL4PqacJ04N+q9emuu74+L2pyZrOIetp0mC
pNOgAz529B6oMvIu55qORFjptGt28shb9HkP8KTkwI7f0UuwrEC9IIEXlrRnviLrCuITCDj7Sloa
71KYwwf3vG7jvnVVUbZDgZ63fLpqM7X2Zz8lBp+zSv6k+BLtrkaEoCyDlHmPct1wq7/vmcyLYI1c
xjAmjvtElLm2hIjfsVvmvv0oPqwfhC1qwLEVMGaCdikEUBhdz9PR9lJaVKD/9PrQmSIYraofrOBs
wkvpczzj7VAZ10I24eQ6lCcDW7BA+EaPyN39OqJJTLC9PrU9f3XJpFu3+g+I2ePVnBSS9J6nOC2z
O2oUcferm7wCTq37qHOGjpq6BqufrD6+hhOJy6cLntKsK7w3/+Kmm1HoDgYdvA9XLRso4x9nIDzv
xBmnr1N+dZ5V9xjXAtLJAHntXwQUlSqJ7RaJjItWNEtUavVsaf/JWL2YmkKiR2atsq4ElnE9a04d
vkRrllPUNLW/ZX+fFwSafFMC33Pi1SxSSsYwp5D9zTYVmw5LKAFmBdIdF2A7RF83JDwR9DrH2KWE
nNOFDP/c15+pXyCJsUHHY7fqbFCdznp1ndcsOZvBtx2ysNfKB93JSmuDLfm9BfGnSZS7jwEEy6Rx
h2AFFuJSsnQB/fCb4vjCNq9WHkRSXZj5Rfhp44/mlx1tDuSzW9opQuG7HFpV/M3HV912i8Ier2J6
BqjrfUc2bMngC5jf5uqjSirnSmBmeMK52RPLSOeP7Ew8JUxjPgf2lF9woJt4o+AYQ2oEzmfNG7PS
gG9vy3RdnRKONJqa8Iwb4fo40FxL8yI1miLmY23YB7BfHbTu5xX6snk6XTXPFZ8fQLHWfyXQ2+yQ
jf+pEaLo9G3Jft7bhGBHPXFT9+Ab7hR8+6KvrvJ4vlhJguyBYIzSOGGPMZL0pTWqQLg2hzIsQFDg
Dxx/EFNiMJDS2zui3UNrnzvvkY/Rq6EQRkR/dtezSEn/aCy+c4eLhXvTWkiaDML4preqMPAErLSu
UGqweiMQLpuUkBpK60T/LHw6VpONsl9yUbFHTOcBiSsMx7Q5WCoJks3Pw0mN1OYy1oAkadVyCVaY
lFZSiFUGtzJy0YFz1blvh27VxBc9VB5ClaJjobr7HBGQFfjETctK5439z1+arD5iTP99/QwI7fsb
SoqWWrOKqES2M8Lw9g9+eFhmYPZE4e+MyoP6LUJCMHkJbKrC3kKlou3XzCIQhozg6NHigRYXBJV6
3cVQ1IKJLOh9nphZMovla9L6rngyrrNhwrdZJOMOXE68vWNb4VYKm54G5nleDaECnSaVVf+JO4E8
Zyiz+NerkdaXMlcjq8a5qD1h8lyOvs78UnR71zI9HKNAlJhvHO55L4AqG4UTQ8cQ1QwTrPzc/ll+
4L13id6/0gcv1SS7gjWJTrr9u0BYegq7pKqDFFiaSr49oxTK3PDjsSND5yxlvjN7j3bYcf84yVe3
T5AuO0VedXfGoINIkNyNLqy/F1RA27VBqWk+w9/lDo57G8VAAZjbeSGBgO+bWLHRkzZ20mQQySQv
YIH+lubPHCGswKRdueTSMzfyjZ11O3XKEpM9vDFHqH450EJB6q6zhZgGCtQPriKno1QE+ejjfroc
OZiKUY8M7v6DN70YcFxkf6nglczYbp9+DtrUhw31NscX1FC3D76MpqPHf8C8SMuwXRo7EDVw0B+/
C1ICAD88J0yJTuxGSs37Ojbd0AmmX5DlWYwv/DSEyDSyprunhz4QE6Qw6eau5Ie3wN08v9hPYP/2
9Y3dWAegbs1QULELn9k04LGBR7M9CMMRBr4/ZpfWH0dYzxQxuq/INknPdtYPXff81i4ejsbDkV6U
oJ15sz4UCvlQupWtfKbfsSCJKiC4qn9JF1c3k1gpbwtoeOMXfUPDQHQzlyySxoWxvU/EX7PFYQEW
CP8cjmyKoVwyAn+InQ/OpClMa2v9gLZMlgog+RwcoUTDglgLTIVzq2wIraLr2E13P6e0i8r0eC9M
8w8Xqv22jnrLtTBkAv6ROTS3WQ6fcP8X2hJQHFS5AyYFG4IhL1QAF9DDMSwqrQq3oAvkzbDId5KU
A9UHRUPdm1BzSE0xKw94ng3HG47D7hxNT0bDZscKgH2RAFg9qyPo4FcNJALY8pKfb9JVIaDD2G3F
eiTLAQFeXp0xv0Oz5KTFZapHCpOY+PyOgQVXC4EX4MAMbV292bAH6CcXqgdKCuceJb2kEfdeiR2t
AXhLUxZkxjr3zKEN3fz60oCcbSDqqkHmPB8B+XcP6Bwa82tlZJiKU8Td8PEN2jVhWzANuiI6vxH/
J42dv0t/TdB8JqWs1Eo8Lna0SwIFiUOeuBX0uq0YmSSm1eBmaK/BCY4plWa3v9bJo8MS+LCrv/rZ
z6Yzlhbf8xfAlYcCvjpPvx2Ji6seef0wm08iOPYq8MEEAGZ75wqYxjoPmnlZSoe0D0bg5f7X9771
19GmLz4qMBxettkI/GujKN5B+6pBQ+ppaUQ99++9uF+su7ypnPXPpZ70zDR8+IiBiVEeI7CRoxmW
xy34MtBqZUvyyNQqreolIHjUZQO68sfLqr8d/ce468w8hsj9h4PAha1MtyK7x/xHl66O//0Gomy0
smIqieAkmZjpK3KCpxYSR7RxCUZS9+cOsYGJMuoGohdCxEncapKJEZ/gKQMlzzecjGCQxOdkfx9w
4OUryT0e48Ja1GREN6gJaYTZ+xsuNaVbB1AOv5CjY5sBWa1oadKfU4hcZk5q26JGR0Cp2BRKqPa/
hvvNRg0fSB8rjpeFz5QGKVFnZfOiQibNRdx79ie8hIr1UNUIiL5bMxafdG1f5TEO1sBcQS2x4/gS
LpW04kL2zKlDNncUuD0mvi/csO+B+fbB3PyengrnWw3YNQoMlOE35mRCBUKCN3IsXluzYYqz/NQw
MqB+qdi54Nb7vFWoylXk94FnAN8FAcdrtLTyygfdaZRq/MopG/0dJy2I7fQfR+BMMDsZ9eKiNFHq
7jG7+2gpdK89Wb0Z3CSxDaqX6Wz7IxlUj5gnKORJQwkQbFGQMKBdU3X5Sxb03JWVIXH8DQG82w1s
VlsE94hyeSUirMGfsalGb4QcWso+8mcD32Od35w7NVpYk6A7L6bAoiW8SsLZ1WGBIlTdJgStHn1h
eyMgwU+DPJKr8eIOkv3zG5mETkmklvZrPVg1WQ2HWurTPUVnAPhdh0zaO+L5x9xSPhqyKfQYwev7
ptTY9kj6AiEvIJ8b+ZVI/arLErtALhoyrqqzq9/z6P9Gdn+vjqBewLO/ZC6wB/fuAlTLTBr07Z0k
po8d+guFsTa6BQ1Q5Yqsf1DN83N7XNrzXeX2WemVp/XVo2VP0BhV67RQX2Z69FHF8gdC7rl6Uqnl
Cirf+ygGDupuV4ehT0fLW1vUpcH3eEpAke8SgRrn0hW3mOU9qxLTeakeWETthvN9qnYhll9uv2wb
ptoO4rT/sA/UjJOW9lM3tXCwPoK13vhmHoOiaX816iwKlHiOwiGZZdzYVva/cE7HfGNATzr8AZyC
wzPOtW7ubkmYgQLjRtYgQyRq7P8P4QoWV3GiJ1O/kJvbGwlJEXyObbjYpv0tSKVac2+L381STznL
cdyMflg3WnjKiou8T0Xy4Bv44a5XckKJtoK2OHFH5fkzyo8tx+JQhpT9s+to22LBmqk4IQz33FOK
iLuTZRlnCfSx5Ob2LoMrQAxiwa1d0/m/V3vVVvQKwmRam0yBC7PMqAIVKFjovYjwv6ulWj95OQP0
PBUURgQwDopF4b/v0hkUaaki6Uvk+DjB94mvc0sEp3L+y09bA2nzL9OhLOMtCm2Ykpx5uirB2w8v
S2jbOniAqvfJn6QqrO5rAOVUQ6dAT42nx4ETakljxvcsiHWS/aduajgGzXVLQ6CC6IFTN6AKTgDs
tkbm8eSwjtxO3IKqhcXlH1/6rgiGjuRk/klZKhd7hgh4VV2wL/0tjyKcRohQiuL40VcdSVPq1W+1
G28F/o7bb5aix+BOEIGu9oAwIibTEpsKrgp8hUcCtIXiHTESjoKy/BVXyMtxN9qYHVEX+odkR7m8
4afBTIIM8nZTOXu7Iia4VYL+dn8cZa0JWexKqmf1W1vOh6Dvsii1XmRxF/rO+CMDlzrVp8Vwj/y0
nuUx6bFivGeRcNz/HOoIg0d5UO+MRxL0PyRaFl0iOxebqbnnmvYWDSFgg35ChCnnufbrh5g0mnAf
km5F6P0PKnygTNPMoZSi0IeMnmTQWhdtePpxzf5vNmaRTcNf2LmnUO7GNhzo/sFBwQM27I0DtMnw
uQuXOU74x9ONPagIpRSPeDQXKyKeN5TyZpf9OfKQU6YhBbTNGLEBt+LxteMMPUNmJzh4PtgJcKoQ
eaLY6dexXc8fPSQssAGDlZ2vxraN6RTNDTiNrAUY4EHtlLeYlplbBqniC06tl4uzgk0pdvCHINRO
OfInd89XkPvH995OUl8QsKUzZv56IN6GXihd0fM38HxkWoi/zOHztPAY3jghf46eAy8Ta4S0QCtC
CQRZmWpOv3Pt7ruA/eQkkkda2l7F639cLZepNFlXvwkT5uNjZRMUJKFTaklwzhu0My7QrMDziyr4
PIH4Rn9po+vUeSCJBlZg7jgI26VJ0qtZ7YXApjPGSKginldILTKflQ0sbSA38cdb2roSfF9wO/8n
ylsHsiy08kwhVcHiSVrxUO0XsG+x8W55deqkOMsgBn5RxGe3vwU4jjq5t1mEbMNjlI5VMvVe8FC4
WDIFDdeboEWCzCafk7Liuf8nNa/HfBrRsoywKoHw7PMrrt3UPjjkNLUozDND9xr3MPITjGv6gd3j
1pWzrMuwwSCzZdQDwLfpRsETk3ZLxg6mfUMlEDYgQE5OCFxueanlaHWEt9OKskg2CsqnOuw7O5g9
2kFUEd0SNljbViILSN9bjNHBHsHz9KafJmnS2XoO24zRKlq/Vs3aWg7JMY9GYtaifpaHqE+LpqZd
PN7aESnyjFbGKNPCp97z+mqWAJpeYJ9IhhzgL307KkYBLYvFwaPksEY/WbF0cBpLGkt2zdl7zWoP
mo2uDmuDBVg2kCQ0xsiIrOJGyx+JOVmPethWbzANk1KpZcW05plTDo54GqYSYokh+2VHq6k2G2cD
F7IY6R6ZPUP8W+xFymtn7fNik7yhOZLbwH9GlMEN4DVNDJOKRHjmU60UF4hd+oSdOvRdE0iHkBh8
CyPROf5OX+4G1/lgpJwry4Kwrssdy6fmrtjE/U4WDM8lY4tlpti+u7Egu/9NB17mDAnxls9KOmdR
XjZAk5H1+HLfioHb2h1eQNyMaIb77MeyC2Tf5zG8zxjv9Fqdhxk2uRlD/Liyu+DIPJregizFTdQa
lO518L9N0Il2/Tk5QVMKkN306kZB4EkuN+In8f6a5TpU8nBUClq8RHCGhypvTDtgKrbigTyT/fdo
eVfUlMsYyHWmWkghM3NT2eoRB5JOkDu06HjWh/yigi75+NS/xH/c5oB1aRQx2Ad095v0mfmdWRmI
luWG1jwkZ5XrLwSLgpBREQ8hVyTyAKgKL1gs3i/v5OATM/khMlezqb6+mXBv0+bpTABtrlO7+oUa
QBWLqM5alflywHsOm5E0KV/3pFiBDj0zxOYTe9BlwE3iQEqGmSsim2MTBh819TT/wLHfj8BTXngg
ifYffmfR3h1MeFE3Qibk3p2EhcZMaLz3LfZA9Ooy7R0LDVqhMYBfiopFg24eWsijO7YGOrfocTCk
wDOt0kRfoaLbdC5w3ohsFjIiImE67oxzuXBnXuhKBzzck2Kje79NylISBovY27EuVJfzBfo3APwr
hisOQ9t7f280F2Fba5SnOtahniyBr+0b1GZnbwkkpjUiGHgEpzJN9WV8AbmaDAlkInBjDRE6m5Ql
g2mdpXEMvvxNHaRIF3oYsX9CFvQbQTcnp9DleQfNHDoqIaAmdoSgomEuLCTEer6wchogDkS3dX5W
Y3JovfvnQIVJD4thStD+EtNkTWhbAYgKJeMphS6zNQKf6h0pLUhB/Vr/chjNsXAnMG+4+Hx1sEae
F4ftcO7iUQTxEV6tPUbqC/Vz8NDaxZz+3q7o54MgbL5gfOMEUxHio3h4U45wc2HlVLV9cKLKO9mB
SEP4v45rrbqkZvOMJYtf6k1ue1VwNywq4F2WSoxvDoK3GwobSvflzVJOMnECK8J4aZZbBEjgkT8S
eq+jVBf3vIXxT1eVi2GpA1d5oWHFqEhq1mdbqIki7ddUSRG8LxMcGFQWrCoJcAoASbv7BZf0sOBf
bd0GF7ot1QtNxxRcWUt19dpx6L9iv2Q0srIesxc4NAa7n4b1zaP1EiybHQHrkaiCUCfZxbKFiQDo
f7VkpQwVozO9yTEbJDrJl6vbWHEpZHqwqFicFrKvKykdMHnNMOzDAfmpuAF6oB5eFiIfkVZUxKrw
wGTyqizx0YubaAbC+aXXeoqzqIN5LAVB3nxOk+pLiG1U+SzchUdll3PT3bhwYUo6EaIh0ffacGES
9jl/JLKED828GgSj7OhMVmvXAlJBKqrfP4daNmUuenRCbOysCaBo2RGrU6iRSZ4nmgzrb7S/sZll
uOtgHBMoOSuhG57n3JDb/8Q/bN/PAeSz+b2iJpi4GM2ciqtTSNwbboPnWo93B8KJoEWwsnWEF9Jl
J8Cy+iXBZYgiosSVHZU/6fDuItCSUgR/G0dnP1NDjcOCxDvFxgD/Dm0sFad8ptxkShL1bAZ6bsyA
JJLBxCPGRpjmDKE8sTnZ6tRSsYzUW7L6hE3S/GrdzmgC8WaIOOJWWT7GmFSgyzQw6EL2iGBCj3VT
c3UxR4Ro9Gzjs/5z5ozZG86SP2Av5iD0yXnBkV9xa90r44IwtyhK72iID9lIVIvLt9ECK0LGBdBh
9Vo39EKrZfqDw3CYgG1QpVkpNzteIPwlU8HOt8nUE1N0YDxH56QJCDVol/3cPb4aLRiUA0PN7wIZ
UrZYZDTk2Qs58maM6YQ5siHmrRQQ28lTnlSsHslJo9zJX1xIkE3ul3bjbp53B9gTxJcxcx4R6zm6
tCgruwM8nBfkdAe4izAzkU31GYJ/CCDiEAfrv9/nG/eVE9jKh3oB87vVLYG5U2tQt5vEcLxwPQoe
3RujDlXH4QOBAh5t9MNOwUxtPPLFQgcXKrZHqZowNmgA5z88XwrNwv603bxBrGqIovxkKE4fEMsH
cmhJSt8OpI6f+yO/rGrrLAu2B+ySrA6+YQ+YRChoBOAjoskYaiuz3SbvDzP52ixuwDJAPDE81l0N
F3bnvgDWz6CiJmZAA5qKWFHHwi0o2CJ9p08p4iGCkwPX7/YBLg6eXXmvg48iRdsxSn0F0Yt9myD9
R7uuG5meRFCngu0hHM0bFGNBIzcpqcM5BTK2PdokcwYTV7wRTI6JCYd4LlqwcW7mQjr61is1MlrT
oxyJqSku9KfZgfpvo2hI9+Y+qV4JaBWl5l7PIfMtMgK3xvPi5czCGc2U914DnVTgVkUd1njKf+ge
uLPQbL+y1TpiB/fN29+VSPK35Y+AtaYVr+Sb+CelPM84ZVnVrhKbeJkzfs48DPdr2406RBlB9f9N
djD8Q+C7PhDmdrAbnp8Pr/9Nhuom3grHR7ElT0nFhGgyN7l3mX9zwIC7gdgVDBrt0a/Bxr14L4bo
n69cjjTGKanvLJiLkaWvioJ/v5Rewq5nI7XrKZQXK2/K7/RiX/DJHXm1CX6Aqoh/SxKh8mkfx/9C
gKyeh42G41jwRIxTnQmEwb2SMw7H49eZHT5w78S2pIQ76+ngsTmJZLhkfg8J3byDsKBYfznvNMHe
QchPLUrPwh9w3k4pOsWUYqk5qjC8cjJI5KyaYhaCe/JqGOFUbTKKlXKKnKjfQ5A6CpccZCaY74XJ
wSq1kUR+nscjgkKiOXwiFYit8UFuFKBBQ2SohcqJpcUraitHI0Cjb56uQiRVM95ZnnUYIogz+t2Z
wFjpngINkAWRGuMvUp0cd2KUiZgTP6EgHNOilBDuyLCP5kLvXwxVC/G2vfChYGJ17fQE0JC97ASv
PAsrWHdFs6HvhHeB6LoBERQ7HteuPld4TGeNduKfa8uhe3jCQ2AHeP4TR25tbWaIumP6QcxCsN+E
hL7sHx6cYGeqjQcmAX1gc+Q7NEzxDlPdh6tqnqFjijdLcnRBRApPlJW7aaVVTxWJzSS/7lTDwNq3
KBRY/ADUbMHJtQpcJ1DFVXbog04qA3R5Ph/VP9VDMT2v83iwmcQGlEhyJR2hj8vNOZIrrzv+LDra
J8OVjBMZGn2GglpEG33Fme4KqhGoFW7/XRkvA6Nfs2NLQmnwn2c7DaM3NppzT3U4cdz5hPhbqhbz
Db/4+370Z4IaCrnAfwuMLAerY/XAw4coczmkVGqwaB1lORxYqAU9wcnrlhfo9Px2Jz9RjekaEJrs
GIZCxRAjQwif4Z6Wv8+Egil5Njt5nSWy9vOu2oRYI2+IZ/Gz2kaZ/3EUtMpemtK/o9L+pMC08u3w
E9si3HfQ85vUizesCkPe0LXfMT0sQouoRGeim1RaZ6AQKcvKciCJUbXZt124fWhFfkpM0YFhyegU
Z1V/fU2lMA853ROz517frOpw8L/jixm8ASThFsSiG7T0/kGO1/qr8DgTexRegWU5vknehtjywf7u
BRPq9TmV5aS8awRQZHFk/oveoDO0WwCeOBLLJYC/ITDKBO7FujQQiFLVt+x6l+xtaKi+f8x6ftG/
I6aLQ/vSCkdfJaAtBhZv8U0KM3d49PHB1WytA1zbdremUNOuNBPYGrb78sVNLQavUcAbH9o+TPek
RbO7ZTCPThb/izWbmhE/e3Dj004azT3u/QltWIlvbMG/o6PFrStU3SwVWRwLATW8UcJgDTKJbwt+
7GhHr+NxidlaqsEZKh2KbPf/NZAbIz/i4gXWMoM2VqhYumrV+m7fHny64v8aSphkMIfgEcCtuXIg
uSWLYmllZH8xv3WJRk0/vGQmd4d6gDCcgHYq0ikIZ/BVG2Ecyc45vkrc/+4j8ar0nSJ8mM847FC2
ZRZGLfTfzBpkTtmUNhSYl2GMWPIhuksbr2eXgPbxN3t0HT49ys2Ql6shPP3RYaqKb/ZQ0w8o8FdM
moc5/HQmneGGadetvhwtk6UmINgcM9paSskwtDhIk9yQGcyoFQnnP/MnJkhc5Hv4dEq8+qsttd2Q
qeAlOdVH3n3qWziIJ2ENN1NlYCdWhg734z8yNZY19J6fHisjoi/+NzxXcdk17xojEHx8S0lju+C6
nwiW8rCPoyruLMyU74xXS6ikF0sU1tDL5BARtDWzrkQ9CWZRXA0iALJWXKfDGTSmzU1IvJbdAOA9
DN0p9x+i+wFWpaFhqX28zfFXbI23jy/0O/ZUJFOaj3GU2IvWwDRf4NRWCIZ70WowimMLucS+4Mvh
1ZDLS5CXb26XR7V/RD8RfQpXxHsGHoey9c5P1gdE47ANOQSjN8l0TztzRLdn9uyb10o50SHM6Sfh
KLJOMHNQgBamSq+F0rYpOONwllp/ZbHLHc95PvgLcfBJYM27XXd0anXb45uIMlvFk2VdGFt/VJn5
2MqqGJ7KaJwKUEyWnJnjIV1S0Kht6NOvG/w5ywrUX80VLjiP2i2wyOJkqcqlMrLLkEHzKuc5vhJV
agnshPANQUT/125ZcAy22/fSIwaWvw1j83ZA4yfKkgARkRt+qfnRHU+Fjo/Ocv+VmHqrqspsOGDu
o2FG480L/6o874tYrlAqVHpfpUs9aCCKlCzzB4xQ5R5lpXnqVA00p9H0ic/nsUuK+t/TfgX8iKIL
xzbN0aQ+0yW0PcLXoFndIfpCBUuIkWajhNuyrREQLom+4Sevca6KUYKJ0HSWULUvkYVx2LuLKHBP
9FZek1N2+3QL+fEW5UPp+i026t2DyS8bFy5oCtWIgVWPVKgov/ShVQNJOArjVDnaD3IALuNX9qsX
zTxike3knqNZzABCB/iZDLtAV9Fb/9zGsHHkQZDcnJE/txRzOfchlxJUJYcUTD7b4hfgzRpgL9nP
XGoTxhBUPk92jpvm8/fPokjedqEY111Qn8DXTqkkKPxw3piQxWWrV9/YDZcK/qAucN2JRJt0Wn8i
sDEqqVXVkF5R2Ij83kerDt1V1Pg7zM3MHOiQYwtfMoP7eJ/+VkCmLhOnlxC7lWHr0MmN40A9jiuM
VQMNo1ql/Yvtskmwy/A+QDmRYWS7P2JeLoYDK244Rw9OYlCXRFLUubs6uA5RmcIjT14uyf4CDh6F
/3/eGyzFMy9Ux6tEgKAvqCLoFmQEY97BF/qZUEPXYihf82g8TUXcKRmHhC04F3MzHsM5WU8Rr51W
wtXuA1qqo2iJUpL2baHlaC29LshrpBTQU5oGN97mOAlQxbg28FXXlYsukzwlR4tn2LtJSV5ek884
jnKCdPM1iv1emwUriL2Hn8K0kPScO2UfTBOxDJZ8PHC0Kc0n8ZkJysMKE8kbVvevjjE22iSePA3P
jMUVcNCqPynhzxdO8h47Z/kbXiSiW5NbtFirU1qZzNwhmnFh/NvgJGpDs4czW7SwawkN304hw56I
0s8coZH8id0YeCLnSBVAVVF7IaiaLh5IHQc6KiuNJX7aSWGX34zXdcNVh5zowkvcCNr48fhTSeqg
/PuB8rIxiCdm3KKq/NDt7JKTQvD1sSyefwU9fZJCgjNmsnau1Z9aeHQp2SvM6aXz87WSGhQ8duGU
Qm2hnu2PWORIfYSLWiShBRKtkTwja7CXvin3rXFnz3NFjInGv2QZOymyubhd0L6GuepOZZuFiztT
Vr7HkXBaYNT4LNbur1TYdp+nx0hYHRpo/+cqhyb6O65cHdbYJtHamDL52hzRtjrZCxqG2uGcDwRb
ktLN7B1k24y9Z9sJ52fViB11opxTArXzsg9jhphTpGWlMNJEPGRp30qW+M+OgERIv2S6FC+XhP0o
+bhEnACf/ZkSNTae50MrtraXQ5I9fuGCOznp49EUrTh85Z8RjA+Ncinqwo1JghnqrVcItuc5ZxxF
oDu8715N0ZZT+KMCoMiFAwbsIL1SfO8zyZ4op2iuibLNwuytS1h7Ko8/DNfiwCPauW021YTDXuzz
me6XBe8+HvNzxRdGupqU+RfaHHuFjJi3k2cI3Eb8haT6OjXpRx5XZBqVyWrwpmRABjXB5q5nfWgk
xbkfSCHIhp1f1el4d76bRjvTdo1mjfP+UDTEz4OZTtbtKebUArblYQ6d9ycAlW5ivsMjMJ3i5zIg
IY0pMokdIgvf6Sm+LnEpRY+LdM0gg9EmgUqmDa+gjXX/WB0eRRgF2OMHZuzrMhvMbwax4s4wV1mA
g2E/GK0g8v3+RRDys62pfstztPvQz20S6vDaK/9tKneRKDagMwvUQXMW+F03PnaKQXhBfUBF2j3r
9Q45FMuzBVRSPkXAQiIDgjpVEjgxmOfbWcT2VQD5ERAy1F5cc611VhnYz4654rIZqr5UaruvXgRc
hTeWdzUKHWmM9rPuZBU3tm82DiIJk4T05NRghix2YNwVOxOQW3QFLDDr7gI8isGBQ0Fr0a9lRKjJ
qOKajeHiQ0db1eR24lM6+HR/rN9EjfDsefQzoaPGFbeErPm7jEmZIT9RIXc/VVBLwKCVxlr36mkI
0a0k0JwBPVyOKr8KGSk90gBj74n0/Eu5bm0e/gl3qR+ZmaHb3P2h6kHdiXI7/1Ty5A+W/q/jfDuN
Xdy0XCT/zFiuehkfSGxH3kLW2FzdyWaHnrb/WfeDrprQtjnHJhrHcBAGHt5B0nVqkK0VRM8dwPDU
tY9KMbpixoOcnk5vRCoBi3hh8IT+I0wqkTTfW4rj9t4Htlai3t5heJqnofogVJpr+R6pBh8YI4s9
sVHgc0YdwvpLYPkO4JoPetaMH7ZcFkMieDmg+kqPcKoY6u6P0kn6ogtokW9WGJor6SS5q7aHDlaR
EH0rrlNQMCY7F+QF1eNnZs4Hb1uLPqgv2q5hT9hfn7r5IsH9nvTYLoDQtBeiyKYBwd8hkoiXVwkJ
P8ifaMRviWSNF0ogAOc7l/R81mi1TfPtHNjQIgDDWUF7GeVx9NI0AyqktQ1Vx2lfok3vz9QOblbB
zPY8HnC6/3yTwJLUVmoRGgHQyJVchDRjRT8y0V/mlXakH1GoM80OB7QjJjnxcy6j7jkwFhLt5TtK
AJPovZFnHHXnZzAURz76I1igcwNMMcEg6OWuHwRhssIRkcGSS/af9NY6+7EE+9NPAVCYTEq2Xg/L
msXV5IVJOoJ1w8iM8BYI7hLOgpmsJqYDsB9xNJAlQOnmXeHjJ2RYDJPT6450pntVicz2iesWWmc2
tDuafKNzhIdnivQMDTzxiPA4NYPahYOvjyOomcvFnSG1B+HWGZPvRVCdp7diuT5hd0fiMofBgszM
NPk58wiGw7OndydpLl1HKLpn1d4F0d/u4HCP2GJJQMdLlSLJaL7uxUkuHSn7UbjsSQm0EuK8iF45
rfmpIBhPZjkUsqUHkjMKu9eB4Q41r9vJ5y4z1B876JbRIqb9gagt4OL35R2druSjypyBnx3Kb51u
I4Bf9LwvEo3DjBX1qBcrEG2h5qhqVE+WOthQmQg7CgYZoxG2r8vtPVEHB2P6kq5pyUF4GfXBoGmO
rWIWXLEu9wAvbniNPVnS5xyEdG+uyOQc7t9zNk6H+zF9YxnNYsmmYx+9/RbmRvw0DILbYSlvcZp/
B5a9eUJ5UwHw9WGWPkrEfnZRoxZpcvUtgWg9O/3ZIzaM9fkElPcYMXJL/Cs2GGVQtmsCGZXtZ/cB
bgIRlYhb2GiVMj1M/RZ6tjSZE3pZQnHr52ngJTavLa3o1BC6paE+iYbvBDRSb11w+vgterQXH0Op
qlHNkXq/JL+FdA7eqJRs7mgNgNGmUsN93bue1/LNUbb4+7aeoXm3xK/XXuzYpFKw+VtJEydJzVca
ab2RRM3JwiYHlELsjgD8ph5lmnQXmpp8G7/9Fe6v+008xc+q3CkiUUC/ONoXDVSpYq5SLMd9lcJx
fWfFcLk00ZvIg7KrmjuXTsXlWYcyEriMYJ0purrhjEmz6ZPkW9j1NeGrB9+ooiO79cmjgkW+5LWC
m2OnjXFq3lRJCvZ7XstgCEwvmH56zSx/EmytFleTHTUq60OeHN8T8Yf1ZGmOdeFheoCx1A35RJMW
b78WQqVasIHO/FCiWcewF+qGz1E6GFQVb0cYnfxD8EqKMswCbs8S1I94d4aI/OEHohSvX16mP/nI
fF01oHOvYNATv8Dq9TtI+h4cl9wftMfIq2Am5xZyiFwc/fvHChdJ6NKptQKsmgS+gdxpicz6jWEV
gU+iXjFJRFCAdtz36iXzPO29C/fONScDvoTIGUXHZ6s8xS5HtkF2TuqQkOOzPDKA45SK7arSMHFZ
CdUkPc0jS4w5GpFpWm0YO3+9NccYBoSeGu2y92TQtVJh1Hih+uN0t89QosjZyz4aJCg0hKUflO/k
vOn4BZ3T6h/GWyMpZ/gTmgMYdmaBIQoi9uWboIMYa12/JNKAloBWsSR1GxuzWnTgCHFYvIrvhWHL
FxZJtiegMCxHCGUHchVFsiUpxVZOqDZI3M7gsa/ImBsyus8Y81DdtLKjOk9bjgDazgCmN45po1mb
nIdiWFswnWEm/TMMyS1iGDi0eFu/q5aCw3uz2F6cpXKZvvalgIrleY8sXyDTwI5ZBK/kdEof4mKM
QvH/iBgrw9snqkBq3H3yhqIJYMiGOitgEZ6Z6p29O0kx/ezgjrCq6tTmQXlLHC6eN6RpGRY/4JQo
risD7GJOOSHUp7oZujD55OiN9eSAZ4zPCzkE36T0nODQgzyjqIExbpoGITiKre4zON2tD/dcQYVH
udZQS69EYmBltYuzAcURSGBe0cByLdty5zHNhc1IMb4rsw8a/xk6Aclfq7pQQ6lmjdOfxEtFdCPU
3Pplda2dZkPfzBclgrFQOyuT3jbaH9RAHXKgSaKLvEBCzqXjaXopCX/DAqeQmPKnS5kwki50w780
fEzBYJZCsEE191ZzTHYBtp95MXr/xih93Pc/GQtOemTtcmCcssdYRRMAPZYB3RmsrNatzAurB3Uv
hJMXasOAL2CUD2sCoshYDjonxdgishDD0YcJg++GucijQJ461n0mvG4BUU/fLNSxYQ9obzgnOk8s
5M1PKLC/yLdk3sJ2do63uRd8YBxo7lIOgYSi3CwaXdOFGQ3cZ/nUeBLaxTXq16Cbc0tMKi5f25wC
HN2aw9K84mhLm3aFogM/fpIUAFjgkJNKH815hMAYlHfd7StoMHRd/v/OLdalbjl03hXexUOTBMr2
ms6F3CwrkhjnLKqMapkn2Kv3BEoRZKKz9nOHGkUdTXeiS0I2b2K2G/9LYrvf6tIfZ+BPAp4heKO/
RTG0lcktsXzv/Naa2TKtupuhKspyQGuuzOF3JmGwHS+bgZqNrE9/HuQu3J06AEBF97cc4mtqEPSc
ZDwOkSl+CvvVD6qvNyNOs3/uQWyIzLFb48m1NqvQ/b/saw2juAMbDkfQif7x6bd3v9y4BA/oaWWi
iP2hWCgtamFTKjxEP8nviKJaB7lHzNCjNxs6tVAUZzfADfFe/MKIgI2EOglFmINgOxdUcmZXQExG
IEOsoUnoCHxb41y8AJuFarNOJiBTZ7GLpNZS+g4341W5bf647cyk+Wdp+TaAFllewpPX3cTjLpBr
4GSxPCJos0UXkpTx10kii51NyWrtW9kXIYaivEPp7HvKMQJ6+q8J6cHWBVReOHf/sRmj0Yv1W2u8
MYMedF1sx85qrN98hbvAHKu7TH6DYhHcL7HH0ISlwWSpS+9aid3Pjg9QkyrX98xeJpDg4HH6FlHM
7ZKkaUGw7iFIUmgoWd9qLsChv4zyF7kQeEyjkW81lZLvfmP0hrmiHwJY5C5fVBXFpcQWwtkz3/JK
000tiWD+8RJqYRYKHneeK8s/vQpvCTYpsWgAD5tHzKlAPMdYvRGasB2sGUnkg9q1U2awGAzrLksf
T0wk0H82GQLHTienlQdndpX0Dumw2KVgqZWSXyTNmbYdozk6v4GJVaN4umtIHiW/KZrptMDDxUO4
6ud30svietgJM96dCRG2+A/+V8Zlj3/pG1HI5tIV/yseyvKHJFFgGo/exEn9eXNdEyKIgHsZcPvU
PwteZzHWc65A93eFVSHfTLsTRMxT8PbkZWOMcizaCzoGv5YMvpGWaBsFMhI82TRAkxal9eMJ5Zvi
N7WRWjLi5OWN4jLLTQ7x2HK905aEMLiESZmidw8NOHrN4C0aRfmMab7XlfERNGZRnAFXR7BnBE+r
+RLbvC/esSB0Nmd0zGgBP/jp/o4GXD3QgKZfEBd+t7k0MhyvUxJ8lgeITsbrksotMSi2K2lsfIiN
LfzR1+Yzjh+S9mJ59Yz28opyPp7Vm/GSB1dUIKS9nVFxiZL5jk6c7B/fEB3AZSmElO4uensc9F5E
3CZKisoGgb/zjYPuXSSacWqdcf5XtwIESuVUwP9HsbXp7v1DThfpiENpdr6bhcP7vnGSZSYJks91
XJ3k09/d8UU22qVj3rwGycP3j50YXxNIyg6daEgef7Y/oA0hoAKrd+a2KDJ6ZviMIqpAdkJdsuGy
+Hjl8f+0uVtzWH9j73iqe2S5M485ZabYpEUvEUjm0up0u1SXjDvV+RfQA32E2d3eP7yQI97w2eY/
B7h7BWv0oH8XaJGe9ePfLHVdvCa1H8I8iCxnpd8US0tepDaAVEH6Hvxgb+n++oEHezfSX/45u+Yy
cH5QwMIlyydy22qOtI5dadHYFjqLRmsPW+N8lhM8kAU/GG4+oN0Wlhq+3l/ziOMVInWmbRK49Hxo
FJEQerwSFgbswDOGukWMq7eFvG2yJt/j25Sreaj6Ej9ENBpfvI1w7hy4YuujSqAFHpNK9Rm+s2TU
d6DLkynETVrDzrAATAaX2MBuSBFuKT15y/4ndIkIJga4tlvHJuuGul91HMr8b07PM3eQJXKCMJ/h
pW4YxLRUHotqAJVmGJpjQOoy2vN7dv9xaYz9VukPfC5T4zFIN5VGDqDefwKeqcPhRYqfSom96dtR
2SRjfuBaWHoxU8CVi6ejML5J2u5V0A1yyAha4vQH63w3bF+DrqN0jvdp/AyCmZ42bTJvmGPtyJtt
5o22onFZ03ALs2F78p8ueH9vVd6KptoKXEgPtXXGfrbUsXp5CVq6iDPzhSidoEUq9mruSYglOgOO
w2FFyrlTkCpdAaF17sGJmA7jO/uk7WSnxQr0gOpu+BFEJN80Dm72fFm+bpR8EQvIJiUNSYXvP8T9
0RfrCZ9C/C1JksA3VkukwS4RkA1IMKw4stHG+Mw5UqZA9zXvVGjs6jCyXF2k4baJD5/8VJ6cjOUB
BK6W+hM1939QkByym9O1SZ14BSxWuqJK4+KeRWyMiBja4rTwPeH5Rm6lScjKo70Pmg9vvEVzzrZN
aV6ryFhqAl8oJxVz6a0BS4aRSaB903UmIYpi8PftW1FW32NKvQXh6y7OJDA4YatT/Z66FOYQb9Sw
N5Ns+yUrEb+X2zkooNb0OLVLnJKNpSIm57qqPRPj4aExyKjqvuA582BsTgQgZv5zRM6j8GgRTmbo
VzzEjG6QC3CJsmAHIb+VzqV1kEBkxlycJIn1/l5BbXZDUCm7Aqb0muY4aE4VNKHbGi3vieE+inbp
6lirhRO5V9xHGkHlwT3av8g4aWWmoNmMEz0N/6XQvBLeBegVCxaKU6Hcapm2CNCRwX8HRKM4SUVT
7bQfb1I+gSWK5hOzatKjGucq+Znt+rhL1RZqikF64glz5vKFTnu+2EkT+lyldU2sF/lbaSnMTsEc
F0mwa3bK1Y9c+szH3hYEkYYxq4dETcqBvIze3MQ9iD+1dknAxyt7HTQcRTj6ZFphX7gBpQdrXklB
oovmNE2IgJjIhIHY6Wxp+01Z2VeXRV2Afi2un08hGXP/AwfmL2QvEp+UhUwC2DTuSHazYZTZo3OR
m3TA5L4x4na+oSKmWg5tg7pAwh1lzTXRLAXYl8rh4rJLKGKp6HTjBAOrSaYG2Dbf75+yX8m9jk1I
R9+waIX5YO7NcoVMcx8B0jBtLn/nkKJ0k++EeLqbxfijylpIydqSZcBQP1KcuwjT8FgdApPUemsd
Qa8434f4koIh6bO3R06q1cBRBqTpBEHdvetToiLQR+uaew4NrODQRatxScoKrDoMVOxEsUQ3O/aU
nCRCW/FhOmF4n60x+5ShtFIkVNMKviyp47kHs6Ad5/1ghwTPEe2l8wY1X5L4AiI1pUT5A14foNdn
y3Nvds7O8O3hPuhPLpbhen8xkJd6LqcntrSD6zADw5MhQcK+ylfkYJJR8BlwRI9G+lf655VE6ZYp
slA6c2960YoxyePmiiMqC23XHTA9bA707s3MJzSoDUIF2cqzA0fr18j9EQr5m79MvMZ9FAQtf/FN
HdrqMXB56xeSyh0SXd8qCN5eg3WdA15MX5R/S5orVT/8ydQjb8xgJSFf+ZbD0GCNQ+q83M0R0H10
uMFWmrfMHQZV5OaNUAqa8nJMZC2VCK8jLdbGwRVPQ2ZEiyLSFPt1/h3kUqxYxXNXdBqsXuCMeWAn
8bp8BbYOoiQEwfDA+3oup0YvfL5APuLZUuq4aAim5Exbg1xJSllF5ToKJ4IHuOViVeBpIJfNSWZe
1G7EUTbY9nrCRk9ev02hoGzJa/vsXVRDj7VtTopj+6k0Hd2cVCnJd1uRJaCcE2yduP177uZSQJV1
WdEJEL8MnOs53hnDRnQD0v4e5vg1mv1DKFQ8b2nnkLyrQJGWrClvcNwdZUsJy1rEDysL7uev2wde
slLIEZdcl3O7L8rGH/ozHPoUbqIJ1fygsqmzXS1pfsJgmV0y+itYMLC7WsGXVBVHL9eDlX+lm45a
801F8qfqLzzvZjq3/vnhSwADCpYgYGq2Tf2cOdYw+88gVKX0Cmtlh+ZRupIIAIbcLDQOychlruI5
hV3EkJ5435UOXcBn5Vro/pJ5Rw8PBUswkgZkWMXBajGbY3BGqI2QpKMVR9CK4Agm58r4EqBcRamv
V59d8nRUcsmaZ50frtTfFxwdBGdv5nwLTnhWsKBDJWr70+7vD5KOODD0V1wMDS0p5E7r9J6Ab/TR
rD+ouAE3qmkHIZ9gcsqM6OTEhrfPvFgKDPAiYBb5XEeyqwvUPev3Y0llu+f7GHkfnHEu/Gb1SDFY
pXVNHX3IVdIbz4F01kM088iHfhWMQOmYqRhHqtI6UMD5ZxOB+cVTgIJxIVABU06nfZHwRDbgPbN9
zjjgPsQwAbIqC9Pq5OIzNhR5BlKmA45malUwa1DO+9H3rVnY8KExCOylbKhuiK1g6kOHjyCQllv8
GpPlLHQbJJvVC2DPeBrRQ0ceDK3XnzqfA3iQao34hQDoy8T8KI1T6EIMlOrE23i2t9aNLsjbBQMg
jTNrQpB3yvbAKWECXf4wjSMwX4L3NM0wonNk2abxlPJ2GJIDOREj372uAYdPNoT8Sd9h/Zj5iulu
N1alZ+LOnbv/upL0HHpFeD82HALkZaQpJeFd8UFZoqjL2fDMcPJ9iAGkwc+gUXiTZiGooQ1NaP/l
bqeygoIBR1FeXK8dW1KTOZbiMGRXFQd89OdWB8jyL6PxauMIy37iOSELX0TEil6+2JjKLI2iDOxJ
3TsPBOmQsBopI+RSjBwksjp2v26aMgn7+XSQ1uOKWpex0lygclVe4nMpXCBqcTaJrfpgzgN6M8m4
MjZltRP4TZdbXrsS1HZWj20hWQIxt55oCFWBH/rFBMzlFP5Kjw7yVWRkUEJfJj3MdNZeLbfyigkc
9nBDiDB03USyhq4tm+jginh3r6Uul7cUk5CxBQl6FLFG5HP/4BhMzWsjB1gs6iGbLhJU1N8+2EgP
cpfX0mzC8tAyCJtq2Ly2405NUngtqZqKDniM/jNNpQQ6JG8aUq9gH5xNDB3z6DtdCEnKSs5D+VsN
9ZQ13S9bKQKpIukd2fsDS4dwfaAMQaGOcExn7cE5VuimN4FC2fQ0cZsG6PubRWaHTu+SCV/zXHov
sl4YKRGzXHagM5T5RUt3oC8uAXt00LiNVjB4j2810f1gl1c9I+rSPhyBB16oADFMWVKwRKht85Mp
AiSC8djM8g3+GZxDI4mu+DPFTQ/+tJojaC/gRe9cMH6YIWW7h1abCQZar4PFGGc3EDlTzpbcgzvC
DEwJawQVnC8QYdvSdvO3YJLQbbeWrb/UShLUdMQj6hdvoc22IczAmX+iOb3Kj+aUJzZcu3j2MDq0
inP+A1zEoIQoUQ46QztSEqmfAwiC4EbspEy2TsABSNb0L9+GJf1JFMlb37FWuYIUavTdjbjL9IE2
4mR2kRA70ogfnhJDmqI8EEtSDDz9nHVXXdTclyD7NhaaWOGQ5FnBNBcOXy9+DIVzgdg672aevYNs
1B18fN0fU5/3xI7O5BP+dQoQAOfKCTKSZiD5bh7EFpoQIDh+7quIDzwSNn6JMqYEmz3oCWM9DZq/
ZIliaPQhXp0Uami2LMITLamraDprq6MhGj7mJ/wmNgv5ewYK5tZR10SR1TBWc302VEDApmW8RVFU
B5SicZUQ7XhjvV+28P5ojiw9nBOC9g1afhye1itIM37iB/nUu6wJEsFE+kno3NL9LsNIiMBGHp7t
0KORBWRxbEvScH5oOEYdkNdaiPSwi2uer2mOuNwjLuUCKHEqS+doQWqkADVAKFwpOVEjyzfwVU24
MZMQxr5B7d1QYwyI8HAAfq/T9r1bq5+bdh+rxoeeGfLL60wIInItzl41LJ8ZtuBrTz4oN95FcN98
z/unsJAApG+pnR/jWTXyABTYBmL39FxFr0rl3FW7/xtwCT08UNoC7Al7Egqysx/+3x9r6KVMqmw1
drj+o5sY4EBAGnZzTXvHCA7Y/zdZ1cy/yXAdSTaOB9F3XFyDZ+3tS5yND50YC/+1q42IIFQrLE0f
lu36BXjpDZy7z3Nzi9FDbP22ju4MvPXZNuvOzD08YNNbDT/NBjOhiEoS5IXQMZC9K3/nUbL2W1IZ
6KRPOqgHUwo97SKiniWtUKdctZp87FY6sLbZOBqYAEYc9Ahxo914kDuJMVRnMBR8rcmikrRnnMiH
ZLaNpFikeBuIHVWhnZLVl4uHxzNjUED5oohllwixVRuQEP1sL13UV1d7Pq2p2k2gW9+FTyZoV2gp
xNlvLrz+Yiy5OtYo12Pqj2rC9pBGkGSzUhVfnaz3/Bzbv5j8zeEY8II2ekoRzhK6vHJV6j29/8xz
JPVW0N4rVsuCO56nYf3TMFBCqwwYK9uudATi+Qx11Vh6WBPptQLWwOl1oblbgVskj9OtCrdD/NxP
CePLUu2xt5FkU4FJKHddT7kCaxOKAh5Gg4pLOCS/i8vwBsAEFfrymtsypS0tuJ30zPJVw6IFMsvx
jP52O0n0Z9mMJhUcZLzPu4E4EiXQnxZM8gEQfvG8ljN5hgby57Ce+0kGgllXRFu1s0oU8KByZCAw
ZKXkh6yhuvJi1u8Aa6ODEfl5qqFkYawg9GQFMilS7jbijg0sG8skilOtn8bDm0wC7qGiRPaNZpwo
97/sVKVhiCENWUjpyOXnADznEjs1n2gAWapOWXW6JSo7qC+4402NjXbwCBmHUUgewRRgog/s/Rvc
tLDLlkuD7Ai2QNPHnqC9/GkcMKha5WgHqcQOCzNianUBK7bZusep0NDL+2G2KF1XJizHJvCO1Yq+
od2NyjYgHfMAHQcKUS4IUv3AJrT4Ge2uCGYJXiVJGIfu5vhcbwt7Z/bK3x4JO6DWs+P/p1L1LgEn
azRVRwd20gniS6cEr97OsQpetbycf+oNg6K6YBoZot0j9w3WW39JaAf46qK9G8nE1manBGHHkCff
gLtidIIuxSfhGRdmnrR6qZSkWeqzO9JTSTYelddwHNHhrl25Y2WEQ3661U6CaP6oLgYb4GfRmuLg
RQH4ISbi6T9fnH8faDk3bKdUmq99yJeFT3LNFvug9jtu5QLvtHfbMVcc2js7cFoefwbkV0QZrKfW
ahDLr/4NO2KphPypPYIGbo9McYYhLZEVMNe1H1UqtV6Uvwgv3s6Ndp9RT4JdPYjvIwOaHv9ElMAP
TCjdAFg5/PH1TmAfcMXB7erzAwMpB1ucCeslZHSdgAfxDDvH6dHmN1krgVOtyqEFNU9aB4dagpF0
xQUrNzq2/y6Y7fUysdy62JlP8B/JBj6OD2pOJqY42+g6LNOAtUanuNqWIJIPZWkHNGS0EEaMu6u5
ZWI6kNN0nH8dXkixqXkZL90AkAax8pOpPUpHCBTBbZwSrFz7Pl95VrIUPSkL6SAVU4DQkm3d1Jvv
nrxyfnERAiiWLqjpyZMMLmE2f2lXRBe0Yc8kj5kBCevmX9Ugj101Vo3PHqcu2N4iUs2tgVsNk4O/
PGZKpC2GWb9oW1jGe32P+OiBRUUbiaO6WmgJaCCBAnsZ3drENSEuTzF3dUys+7oxD/ZA4Em45EXY
yMVmVAuHycS3ZzqQMbqmcixzg98jJx6KB+MpnrXh0ccyI8DXMMYRZjDorvtJw1AXPK6Vw1gbqlpG
xP4QElenq548ZomWGAF7cEuiDmhLd/CY6j2Soe7Qmd+do4ZL0HkuY4ceCYa8A/R6xOLHiLf+wavv
8tTGAeJF3xNbCAvYpzP8afnCKPGc2UQ3O1+1B/nC6Jaq1j2t1egFIwjMeS43M/Eynjm57pXuqz90
rWubvqgWREy+lN/jhTP5vOQwolvssOPvV1jRrXytM/s+svJhDFPOFC12ZHmZMjuFpbU+YTqphiUq
k+Rs0qXIqHwh7ckPjET38mf0r339pfbWDyNqAlUOhQAZZpKPb6HdGug14eeiuI6KJWppv5qIjkzr
xkbPg6/EMokfzLwHrSqhmX3EkoUKNO7avzpiG2ip6dE3CNnbFAB0ulYjONOk5elErFvTYqo7Gl/3
DfXw83VPXd1d1PTkqs8Fqk9xe5WrZnu/9oWBJkgVuKUpGOCrERNLkdJfrG611XNe3AKyuwBPpq61
C314A+zk4OoKnpF4RE1/f7njGFuo7qxvkTez8bKxVEq78HUb0VTNPheLd5852YIw1ln94dqaz8Mo
apiGIFaFSIRNqUD+dxXk0rRZWLXnXDVlo/wFZ2tRs895Ef3g/FB5BA3O9otQ9gLc/YML5Q8ZBFzb
oSzOR6DBB0TDP+4lTIH9etEvaDpj9ofEduXfPyJACxEBBpkHUV8ATDJ1EOfjHflsMdMXkpz2Zf8+
O5WnaPaHW/bdoLC+2RKLBAwVgurQrMmsCxHx1DQti+8HhD8YCIR5Djte8sasJPMOr20YG6SYwRdX
byAQqU4Za30Twgh54irxHUGp/YYEtf243zzU8ygg3jTdc4KeOSXrAbpmzHW6L37N58iZL3SVBWNt
arQLiOdEZeI6TltpvnOroONY8hnKFT3LWWaGsy0PGVWofzzpwDI4/KJ9QLhXMrYzbjRq/92z3VCL
iegHS1u59Wag0xlkWuLhP3BsURneHEaek29O8OCu4OeTrN/XftNPPYXCN0QJIH9rToRe7uxdyIZw
dc6gFalCdNIXpcab3XFYzak6k6O8IU9BQMnpPuO+HMk8/U6q7SctOYe4bnUkQLkPEIF2s64mxoqP
gfqBs3esZSF6bAVxqBXA5/3Atq1bCijFJSR60I50d2CM24VekUOCTxOSrB29kM6IhVnfG34r8YmQ
af26ZKo0q89mmi7/UQT+tIEnTW4kq46cnmXM3UsZuOnzEMNTPuRcu/ns4UQDE3ucpkAxmnaeaasU
F4BqJaMQZRe0ZuUezK2oxcucHwc1MFSvhBPMw2KzFRr9NCqbWd+pI2LTKqN/E3oXNlOTcAcGowcW
Fh9hZBiVBJcp3QaqXcg8n18Eaenj2pv9c8hqVzR9t9cxXoAYz22udjHCS7UNCT+SbkulCdgPI4Er
ExjFrUuAapgIyhEoCqAHH2TrKdbMN4ec7wWpzrY8LkTW6UB0uJ1exRJKdj4VIXr3yEyjgQGaHz9G
m4nS0Sb+ATbWfQulYW2/OLe3e6+kg7zFUfbaimx7j4Xk8TLOdNNwJLEpe1yITjQrOWfEjKPKslQt
lcQK98Iqyzxlp0123Cfov/+H1XoB9QHTEe5lx4zU7nOfmuWMKkRa386oh1CB5YItw1MSY4jHGI5N
ZFCFhcLLgU9/LDR1leTa1RN+FtiRnzkZr36HMCKoR8gfnZwtGEle3VBdoKXRPaZIW+ebOg1wm+L4
jix30akYG4xnPSYShU3Mwln8s9Pj/KaYiHl8PAr7iomxkP0tpHcnYugDm+OmGJ7/PBz5pg0WP9Or
/v83XMtwZAFEHIG9n6wwMmWAqacxBLGVWX3mAzKEX+zMOhBnfC52bo0O+SxWNGYwNUkA1GCRLtIw
reA07C2QDh7Cn/oLlFoKPjdlkAwhrAuBG+1kZPCNL/N/PVCcFcHjSy4I1aP8H1VTzUuTL+yYPbQH
P0z0I96AcE4R8jhPXbIW/e4a9ye9vTXLHR8vG76H1D7rzj+y690JVb/OnADJE7eOztC+c+wn81it
flgwAKJc2Z0T+iOH9VQCRcwpVMOFC2oT/zHejwW3CQZc7jdIBd9PX6tzKSTSAoePmk4JNoycJeye
b31FBRKFhB76cdlbA6fgJvXXY73FpRDDQD2MV+FOL6I6ZJMPqReE599R8wTV2OcAKDDZp5a7CbBK
iEVF0/58kKMM/E2mcpnqQWZUolb7OBCPC+/lBaE0nMJoTFpLiJ/QaHiewxxfwDCM05p30ya5EkO9
brmyOHZxyKlSCH593wXBaK5HFo1rUn27X9kHqp4AO8gTwLjPBqxdLvRhLJRJt90TIX6Jh9WCweO2
Y9iqTB1+WZHfSvfERrH0IT0QNejjYN0kvCsLaeziVx+5WLQwtep0vczBTytGvmmzGJRiEW69H7da
SvPJXKSZZPdefIDa58uw8UGSQZHR+sCWhFjw9u+NrDmcLMhEUHir7CN5ple7WqVu7FsVS+kc4uT/
XCuDCZzAsNDm5WAj2AKBQMOqbFo/0nj82K+munYi5pFLH6iDXRBqrnZPLdcAIHh95pbFA9F7nP5t
ti5B6jrWd3OPN3Ol5ogP4jThINyihWPOxk+taWRD4oC1TWFsKJSkp6mzx0LyR6ZunNqNcrZrlKK+
6wr7QmNlO3YaC9dYLOUgZYs6ciZGIN4kGVOsyEWcXikIpwbfjfFB1tWeWO1ItTYT7mRT3sEosIM2
FCSZxfV//duLDBCh0vMDmfRAbtAP4tT/kpfpL3Plltmtf/ZwE8RSCSQiscqaDgzjCuuCV2rn0XbE
BfUo+0C7smqLpoGeXGwdQQFXcjHs0xXeaVbXxDUJngcCOue4JQo9HOmwZMIqfCYxhjdUmZuCCcLi
EY+Iw4CTa1U11J6SmjstQvO3tPVcfbhJfXkD0Wzz+9bRcPvshWhWqJy10mcCc3kgz1pNjaAkukFr
ckC2zu4f3ics29al95qzWwA8sTTTos5CzON3p9j2HpegULcnoMi7iK4AipqSkiMNn+ajePg9BkGq
5w+kV9kHSDD0DC9sxM0V2sn4UcS65B7EHTXg4nWNuXjxGldBEBP8dOPtUkWXq99ObGvgbECSZZnh
PcqlYXpCPebb8gkhxZjED9ERV6AeaRStyR7rhc+Mg0nRvzRE5drW20qPDm97qbZegT2U487u6pUp
VTXekezIxivj1bGM6F5e9ZYL5TRh0It1q/sC34u9mQqM0xv4xYD2jgJvhZrcJKEN0YSMWvxDiYCq
FAD7ysHXxCCncHNce7bS95Fnn0l+GwmvcqG/+4P5ntF4n1pXa0ozhqKxae07STis56RcXzEztLWf
RTd4bvAFW2yasIrM3uZLUrT9JEaFP1cuJRuYe3+EZRejTotOKmDLYgzWvRrG/ex39Ipp1KgZ/7ui
sN7VeY47ZLK2fAbtUsSL/IZ5FJF/ytL9ApVKTDcfRDrG5ngviV2qV1hlbi5b1mk1bhJJQ861qPd9
/X6sht/zlveBYJTcKZw78L3g4RdSYS52xLREpQtXy8QfOpmYAV3pqIfmterkN/qZrOWI+mumd8fi
l+BTyINKX1ah29/y6/7K3UbP7tMp5kG9tFVFBDsTf0iReqlVwri3AOF6bh434yrn6kW7UWDp8Wpi
dVHzjTmzUnl9q1sr4PYWeMjkD7livUBMlFf+/xtn7zAyUEWt5JSyLr+XSfXBnpKpXp5dDccUA7OI
2/26gBB76UriUE2I54ILOIDHB6zKFMKMrRRV/IYfX8zF4aBz0ektr1ofW5G6fmEYfWi0se5JO0hK
j2Q8STUK/NmdiJvoad12T5gc7gdxn6VzCgIzFkUhvFJW/A03MT0AQHNB6EYHug8AsbMMglridmOs
peXPi7Nm4M4YvzvVtJun2mSPg5t701cVxj8+1CDuDhl3+wIExpGxUR539Klx/Hi42VpfHYCK6uBC
NTZpqqWh0x7WNz58lG+LZ34bwiYpdJMFIAp9xjXxkxlX81tGfd0P3O9C7+y2fykrq6iEsWx7FbEV
yp0gPOtE+E5ZHayMLafjcRIsrJ2bBKcWL8cQ6V849FVNcA+jcsZjsTHKuWBth/eX/TvMzmfJYlyc
SYfa0j7d5wnH8fwD3Dq423VVafd0dgaSXd29jgNbwXUxg+qEBlV5ki1P9E0eDI8pGGngZ/e/EOQv
TgIEB6uFokT0mHHF6wZonMaAfPQFbXGa9c/UDCgFBPM2GJHSjwXYWwux9XXum+luES4jyAWO6XVb
vAFg0LqpbkxPwwmTEkfCwx4FV2O2SRZd0CqZ6L3MQBzZ727JxCLAB/9aXHHiRIBeyiPV9H9kAxg7
7XeqOTGP05olZ0ih+o9d70QDU3xVW4wMOJM0CN4zyr4jd7SNQnRsyAaEZcprQrrzhll9HUBoDhA1
bk3GOqBRaQGOKNcJihAhFQWAgxzGxA+pWd6Dtgnd9/rLTT3pcPkmKQDGVdlELzuh9ZGbV6AQt7JS
A+oOEDM3orzd25j3a/i1mSSTjt+3uPMPGQvUs5frzGjpwyy8lj6f752NFBf9vAu+QUOAX0SxXGkW
QXDccd+sJ6Uj+r2S4vfBb94tGyZGAWZ6AkWnG79R9l4U+ov6jpt9TvboRLQH0GSdPo2c7fUNy6A0
4V5iBvVr2Y4oHKFoaI9Felfw6zIvHoXzqUyh/VlfMerXsMQkHeh415bP+2Y158nEMOYB2DRx57Jj
K/DJPf5p/pkQnpYY/qglH7Jtr2WcVQKJSCJMC6EKIoGqtom1aLHpwSMwytVDruYArzVscVkOeCDZ
oANZUWA7ECcs5pE2VsfA/iHsJS+zFf8HBRon/3t8nWStphsqp2UGX8xS0/eNtTGJO1Twrj9c1kfq
6kvuZXaLsJyJPFYJDbxs5mlMayXCIYdHe2FNSu8wB8A1LpUlDmg9R5Ng82bvElJP1ldrHgcaIyot
bGh7f2czBH8IsUdll0qSsw8efgaMOHrQHCMgkls56HA2mjafKTly/Nj1vv2WC8hKbRcBYCzK1PVz
TeTGyVUq4hfGoSdJ89CUz6F6c5gAzGPs3Wiavr+vXOH4FKFz3EWn//a8xkS0WedAib8slp7ze2AY
Po2uzRl8Rwpaynim2lHghEXOB9PBGfmgpdKYpm3l7ZiYggMKFyQEksz0ak+zBCNvb8vzBgf+wiWd
iBeqphuUXrT0xDnRcOm0HcrSkfCW0TesLOTs9oj8Jz2vxFioIlt9l7aYjEYbFBJD4Q/V88gTI0fu
BMyp69uV9zCLL6Wj+ot2JtGqgugawkWvkLVccP7mnUUYRyeNHekPGs6zADV6jLfvKjgd+eH2nxIU
zkW+Y3Vd07Qu0djZf1RvgUCRLU78SJ3x/6+7L8zi1JshF1gY4I9EZx9CSvV7WvIJdI1KXwyD5drR
ax8784+0zq4tShHOCcaCznHKXSDQKuDQYEMNjJdMylLeduaK05nuEe6+Nu9Uyv1KyQUHKGpLZtpn
6OfyU3oWMK71vK51utWFRYnflNWmhL1FSM0lpZdZiDBd+vU4kZPmSv6a1B1qH/+laF1sxz6a28Yt
eoZFg4ovpcBf63K3XG6V5sZ9sVL3eMXt2Ck93tNRQAnxlk2EK3GITPFUSYo0TOVuqK/xVmMFt5qv
b/BMf/QoNQRkfF1zduwpvujetalHozDN7AIercKMvR+P2UlxyH8SQ1A/LVAt1cSP
`pragma protect end_protected
