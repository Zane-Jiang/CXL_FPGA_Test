// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J98lTjxwjvosc6cTmj0Ckw8demCXq7foBdlhOgMfj0nkYylEFJj00uZ8D9RR
dDgZfcG/SFDVkUdsUbM+XpXbZrT8ksKaIZgTddM+hGapPJmYuLEYJLHzyv5x
R4dWqt4yIeNYQDy77v9+zr6diVkjBW5HDW4W4HlHSRs6gbs4fPvBmGcg7AUt
GZELjtORBP8H3y3YN/TRPZar6h4nzj40WJJb0zBn3RwSD8ul32we7St6WXry
4rMlw+A32guziuathPUCCBciUnMM4nJYE+EbIEop1XSNlI3YPtofBAJgYjhU
GACdElyODqlZ0o6cu3pOTXH6Rqf1EPTcDD7WW9DQsQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E6uh2AFPibILN57lna2eCd1uT+5a+b05HMj28YD9NYGVeQ+osvl0xyxQT7UH
v2B+WQ3r2J4Qw1PgWlaq630MfTVQKP9kQ7a8IMmHQRMsVhQcSyovDG50XPXm
olsaRj1HY1BDiAH+fLFWTaKm8ZCHEu8uZGCR2Zsvic8B7omTbpf0mVl2lxzy
EFN5CQP2uKr/5nQQyQ6bz8od5o1P4m6rMVSoHQ32Se7k7sjcUR1WhSvcAxDL
78JMr3W0KXSf7g3WT03fmazQhcEHt6grr5fZ5TlRprfLf3zyfWWcr3IOrNlQ
P69/YSERmYGhu15U0PZZZ/3NoW8XbbYUoctzlq7ZsA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NDZFDwbFNubSNGgfP71yjMzc0ovx2JzuZI+783j8+55phCNHJ4QTouEW4nR7
ATeKckHlauWzWnvvm528Zu7rAQ8R/CyIzNXm9s/fvXtyLqdLPxElahkUP1AM
OyztLx5jcz2vvhB96U7KqkAmn9cd6RlwSMLpn0UY3z6fTyXVjReOh2DO6PC8
fZnD+2GEwJcqC/tzICSBEGMcHkMLwUKiTL+RF8ApHQuD6XsMJP1M4iviP8Zy
JCyYy3TMMKWsJmx/00QE6yDz2rhGxKQ8jdpYqfegsFdVb/+LnHbzlaZLkLjL
tGnz30sEhXK9Ut3K7by/uCfOlLYaIPjnNKRKHJFF4Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oQKdPkpyN8aEt8ZIaZ54Vm3xE/ktCEEQSCKHK2zptA3b4pK1rH1rP/BgW382
cRabCnaqlnSORD+vXtdJmkx36qQ8D8CHejBGwuQc7MbnjMv9HzzHh66HrNgH
1dOPq3AQJx+XswYxvEOZkc+m6fTftwfUh1Yf3aGaxYTFRySq5Hw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
fRTFv/+wWZRswh7ZNgYodKcKAqfXs1Ze9uMpaKM8DewlqwzHLBqfko3fiElE
KVP0fLOr4wtRDlrbsJDZBwN9yF0+PUTOM5u2qr7WpWcJK+yCIRgNN2EmVbJ4
1Rtg21Ob1XogUWnIwf+ZyClZvQAT/V9xIXC938KZAGJCfXeSCSzTEfOYPwgC
UKdlDUJpP28gxZltdzbUxksX3vg1FzwunK5bWOratJZ1cpUu+qfeYSLDIUNU
KGyHkQvmUpLXgMx4q2ktx80tcrcwxwh9+eVuklTMncG8asLBF3s058hESCRp
YaqHtdQ9Ew1iXhHLNBOfRh+Bi9FFoQ7MtuDFLS0nonQdrUe0tkJwhf17vcyG
Ual5McLnpXmnRzV6osOHjLBfdMVgE55nOuPQ8qZ7a9hA+U8oxjkYU1j0uT+x
Z1dd8erjs8o/ZeHQuOF5Jc0nAi6vGJNDG7b5/dXCK0Y2BCg3fGXjPtgHf64I
A+SCx+soMh49knxxBx5noWSiTP06lZmn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q0oF2STO9a9n2AISgDeQeWORgOfUPyrlq6Tya8io5eB6JC2gw2KMiwruG2oB
flN86bmIVXKC+xbvSNO2q0g7dD+NS+k2wT6b0Sgz4JwjGgu+O/DxizzUf1Dy
OqHMo/tqHrqwhDX1U5pEZOZlCEQO1/G9+SUcRQOTweHzI0VYCAY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qupb1XZksTRIljiffPqB2zz+rDVTGgOxhvHhCKvyOacr7XdlN5pIS9XrPzsG
HZTZFh80hB46xKDE4UJiKIsIzI+lo+qJYpWBOYKAuKnbcSZ5+IsjmkCrVtg4
p3ZFzhCvyprUL4zP0iVCKJsJYS1G0AsqENArEMUwD2HYP9wFXTk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16064)
`pragma protect data_block
ZF4ZMIqQ49mcFCkCHSbFUYNkdxn/rD1M5b/mZCdJ1PFJGzsWStrlk5KD8Z/q
LLbhrjDrXDkWQjOgWbYxgXFiDRUflmobLOVAm1y0uSqgUpNgbIbc+wWgMJfx
cXxLZ+FkFapNcbfmyaXBzFjy8vEW+ZEvm2dYdhVhCzE7idVwRnBSJNLwCwDW
r8iGQSP9T8SNXLEEGVG/B23CCvxINKODjHRe50d/I8ZKjfaj5u6UcIe+8gsW
FsZT2bATMJ20eNx6DjEE+FPxXBe6T5amaunTNz4Ubk5Vfb3P35wEyNMRehgD
kaha5T50o/Rl0lao0kaZhM50jJP0Ggxm2kGOdk7BjiwrbO2IcQNSfzJJ3AsW
0UsdptlnknOJjx4I3Poko9WAX2OBg+GEij/OBOrj0c5zVDGH6FFy/vcKVdZv
SJ/TIWj4JAGd+bUfN/oZiE+1/9XMAMTmajFQ1vUJYrpb01UxOBY8q8OuKKBu
OFOe8nPnq8c5nHSFc/MQ9wGIDkQV3IF/EcMWsZwKp46j50k8DKXGRILHTWWv
i4FwljSzQl/8/YB8GspUBmPVgsmeYa8QThY6j5m+sOmiaBERGASvmJu/6avU
Di0Xo3VSfMoHcGf2sJ5MJKwdyJJbdxq2uEpRjlPxm71wd70bpgSYVrHmdmCw
skjSeWup8OCfaZaB51KyEDLQsuocJJQB8fDHTDKGqJMa0+00NW7D4Y0SmUEl
wV6eU+GG/RhuqucGrSbIZxtcIV+P0tz8NtOOZuHP/zNOmmUJ/3Q3np8WW74Q
PeCBirIZCcJUGZCnUO2U1xV046IOrcKC2Kv76BraQw/EceNbER8fIk4yA8i1
EBoqmCmUnrNpaW8aKP1z4A7+VSEJbtL0KPtzd9a5IO9R4za9KXSWml2tmL/s
YhZGalUS47gU2H5yIRoP96NCm1lCYHI054kqDOM9iDe3MwJBDUSvC0e3BqJy
+/1saB2FUSKX2bZCCls7VMlt+nWiigdIdz/cuXk14FGp4+2oZaI8h7l0U/VR
ubMHzQjMhRqEWHqujZgmbkIVuZeWCU/CLsNeKuCEbC5+IE4tUjWaGhXj3Bj9
QwgqMif+jQbxADe90r3oQSu/hGuB5AJsi7OBqz/HcTa/MqqirRLw3lFvQ7T8
oICZCBskZ2iKZHT4Cgf3bGwYSZvU+mdt1HChniM1jJZCuG0Ytj5bqqt4W8s4
0PQ+Mskd7XNrtYJIPVHa4496MuMnfgnOeJTUIK8Be5iOJnBn0F1wR3hBMHHr
5XKC+H9j3SoyEO6m3HUnPt0nWuJFoCmP08ZUbbuK5TVGn9Ja2KxtrT1VIzxb
3cBHXZdpkrgXrmAFKLq9aSsJU8ZKZNRufuwRs5dIYuG7hlwtL6ELqAOEtxt6
6D/Ew0csnF5CEB2BMEkSMRL5kTTil6Oys22lw3HkoMDlBudQNgSAgWmPkJAa
0jZuRUjfpF0xKhiBbROZSacBXMV1au9q3bYp5QokRsH7ZP3luHo5FSeY4CTC
JjhUq9wGDKdvf0U6IglFDZGkoZOwsukHC028SFps4AeL+rR2uPbfDXBiJz2m
Ezc9AWNmqOeA5QzDSQHrR/4hm41ue6SlJUPtC7SDA8gGKx6bJoXIihDgyxVN
luzlAFgDlC2BXtdPmODn8dJ8Ce/rdphIftKgkG8bR29BtDWeqvEjcY9JLOhw
NSGyWCxBUDJjw7NVY4L00omFUXbJNA2762VlP2gA34+pR0gzI8wg9FU5unke
7PU0quIvGj/fSqlvGaJ/zCBI4iepZpE/lU2HKsaZxH4KvKWfpV3UaiOW8z4l
4xfxfR+VH7KhDG759BS0ZovGqAZmJdvLwY+ATAG42psVTKM0NnnNBCd5OkUj
3sfdYDsbaFuCeLj8M/yktlwQns0Yt+qiH8UqaqbhUdbz3+eJ6s4MAgheuiK4
Un3TNZerffWi8HQwAUxplUsHLG8pH5g5Lm/0TgLowGJosH+s+yjWqdWLy76C
jVJxouuDKS1/Lc5vTF17WVODkzWc1tbMBktiEDPHlAvxN1dltulQ0quEl3M5
qBGpV5Sjff2AH3Y2RE903yLwJRkZ0etwOlAxB0HyI++CHUJ7jMLyiyPx0UjL
ix4ce/8L16alNMV0AI2/an8dXMbhIcKvWghzCZX4CXgiKr2R2J5JCfEm3Rkz
9ng8vicq88leYJBAL/RaJ/0bIlCu1615gBwqxEp7O5IuZfYmu4KHpceRp/TC
YP3OMkjNBfEMO4GjAunxDFdV52Utm9Z4S+1MHoxOamf2dqUURYWFbMXtarsc
zDNVfylvuK6oVsYqUCHTyy9hI6y78DQGFvKcpH8Nb4uITebMnxki6H4j1G0J
yZ5LrprIJmB8kw6P5+aQwAIr/HOEmqcx9deznO5fLeNLilEOnKe1BeT5U4yW
TX5400Hm7yG1QmNmZdxOqIp4F7ev3GhtULC57gl1+H0iZwDthb8eB1RvTXrV
UmSYLZZUVrrc6Smm2sxlqV1JrwcE78pVI6aHZVfyNR2KRY4USfHK8YBRuBVD
+KK65BqUtSTENKNwvr42f20mPlgiea19X6X7w7ce48+Ob6xihgWSB+jBO5EV
tA4xlAsBoZ/j64xIi6UskvIo7XokRjXe8ukH1L7dt8HZDLzviGSDcVBiseum
JQ/Ko6uaQM6bvyrE/7wo2UgSJ/zvs33lWE47V0kBnA8iuc5lPiHumvAfCAUI
auEoqq/LIEIa+B8pTHXADLA3OEarx/M3phdO5wAqbzvYGX/GE1aKXm3oww6d
X7Xq0Gr0eUMsl73JX2S4dIaIrCLsZds/4jfo4ez5yl19YwxBqKqGzem/nLgP
RJ9MFQQnfSXJ2Yi2dWigdTD3zN3xCfW4AQUy3OFhAp+LFAYGGFX/sknfynqx
/9Wzulb7N5fgqlV0H1ixJVvwo690olEiEWMMuZpY+93aOt2yeweJv7qvWv0Z
6xIzP1C3EJmRRc6gb5Qf+hb5EXlRDOg92u5KYenVqBOOs5Btg83piaQxnG8v
j7RwXC8REPqqnDMHZLUFcFCFqOyBAChKQZQ3SHpsPJu/wrpq8B0nfN049klN
Ol4HpeGN3fjclpQwLVRVvPsR/fZE7f2TtFRU3CrvNmvYgP3ZiGJFYrAmKgQT
ZBZdbfcShiLL7fegsIVht8DEyxl69Qqe/qedUwBzXJ0E+OkfozAUPCqpEYOc
FPviSn2aOXS4LWsI3/bHG9NjLATOvMvI1Q/kA0aDCsRzhn9SZEYVe21PSxy8
zAKeQdc+R9cQwoGELqa+WPn8EdALUFbPPx+LcyTwH25Hh/KDz47JYColIyqN
zVGl/BWOFrkSRoZpcOyhSHZH4J5w6tkw3Ar9fGpDFGTNwY3eWCG53Ubo3XiH
YDqE8WVswoKDJyiT+pfptjL4hZfBw9HMTWs0NQwsAJSNdbCMhWRNT2pSD8cm
53KatGGkZUdU8myh2hze8tWO3RwZ8c/KT4kET2hoJ+wLe88JCDlbmwCzxf78
aLxJWuVDqSuHI8UnNY6/5Bt5EyO31bDTq296dOkmCJ4cpYv2aWeo6K7GsPmQ
/6YxnDrN0YraZsUtwMyyZh5cGyg0aQgWhDDH9pX04bs36nd74igNU/Dsl83N
1F6kHKz+suMZOcOY6N3syydXZvUQZYXAuBmMZRngAfLiDBXNiMHe4RpN8MFr
9l0OfRZLheC/sEEJYeuURKTQPw+y8Txr5M6957XvNNtbugmeFJnc4Ly9/HAa
le6fCf3WE9lPCLazUVxnkk/6OIjpPFpv38IUl8M3jkFS8LnMw6l5eDuenvYo
LrBYcGoacNAMOSi+461ljfBq8ODLnY9GWUNct4FHWN1JXgalTFj/Ej9b0aam
mwUY+TMCGpB3JFq6+7WbQtF0XDk6pLsOlLfLvg9qMEhEUJ5gaz8wNNt7aVWT
Dh8GGYPI1WLF5FreXCHNPjegGGEVq0JwCZUUd/fylrVrPDod5LDWiCvRUsyQ
+Qzy3mQeAD7nB5JoAKXWyUgJQArZcBRiA8B6ll3Hi2XUKIDJZsR1b74prk9K
6bH+hWLDLbfiVrJRbQmmTzBx/P+E0Uafg3VFqlXxg58XtgjTOAZgRZ/UbxgQ
BDVxf8+UUqp+h856EN1fdO1sebOFxeU7PfGG62W6i89vootModY9PokLL9I9
QsHInXyRYd2T/9TOyp+c7/5R8/sF0fqLUT0MWQhhqm9A6uqHQnXSKeJWVYK/
bqLqNJZ5V0EPv2MnoxWWsaFyFGxMWrC0yTUbJPQiuG0fym3Q7f/7oBG0MWyG
m5fMGUrCsN1o5XJwXNpqiWG4omib+7nNwVAErRyiL4JJjiNy92KmvkVcVKtN
uZN4PfIcaOxXgL2TZ5hs2anSej4z84DgQEpvj63vWqNl7M/9DoVFthnKUXNW
0Wo7WzY1MgZ38MTZWKtJwrGVNRGxp+/RZFRUlZ2ZTxmziz0tmxKMdctxXurV
uXQuXkw7VfesX1Yu+q4F8/S6r+Vhdpy65c0lTc7W1wTJx8aMyMTZaFoemRb6
uyzHcnfLYsdIctBzjeZ9UdPnbDkl1mqHUHdZUfo6Ua1ThGDniPtGmXn1+Vmy
oYxe5uzAJ9zAr36Yh4yuqiUTaEYJznwtdP7EDUDgfSUaOgLCFJAtEh5ceKiA
2cHgAtZKejxyTiLJPBFl5kzBJdXOk8mc9rC3cFR3zeM/5t40IqFxqbx2KP/t
fGl/JS08FkcdMc9glr6K7iRt7D8fFluWK6fE3TmtxVcS8rRCBTKiE1ZT0hL7
RHpw96c9SVGd3c92HXW4Rr1C/0nwLbuM2rifdklAsFbnuB/gZU04Al6fvw9l
r9eEyDt6ke30FN+wb1fvxxxPB4eyfCx7/ffZLq1kyiCIZo3Ih0Ed2q+PshJf
kOy13O5DzYBQIN8Cdqa3JkGBFcyI02KsGt1W9r8Qbll7cfQaaMlh9yzPKFqT
DbAuVdqiSzOKolMAhyM18y98UFEGdqlzGJUwIJQDSwKQezrfmUIsOTz8zHng
4pgBZ0iASmQ4527zeloEi6MESGodVqkH/6XbxbV5b1SUrCQUhgHggQAQfBh5
EnJUzxIZkGXzeB0Yc/m++wtTVLEus93eNcKloBS8Ca7t4kpRGz7niBzbU1QB
k1MDUFR2LAUb0PmfZPK8db0pBdLdS0Sdjxksb/VNB/HrC/go2RYO6JvGBI5p
Du/dEXvvsA+ZjJx97/1NOWPAm0e6ba26TUa6dY5OAHLivro61OZPRiz/Igs6
XlKtsdevaAnXHApdPEgSJcA1gUiLjA3b6mYHhL3P6IGOblXWsc09sGo5Yucp
p0gzIxlY1pIp71pkK2v3FxEvyqTfFL+NhTKP/xFp8F+PZJLcymgj5Yh07+4p
cDFwOy49fSdrFRLYa/VO6XhJPmkcJc01FgTk0QDUKR0KDHRs0atf0tN0wvA+
/o+MV4bQrJPh1hYGCAUqIheEkMLCwMm2Kgs4HtnUuzY/n6V6CYCBzIm01H/R
Z0JC55QUcTItJ1yXFHrR8w5A0wr88Mn0pi3F4L+4NXUfKVC+xqPqt4/fbQug
falN3SnLTzXgirrC632A0wli6KueD8ZOzmVN8msNDF7t+BTbyeYgc0iVF/sQ
PaXLL2oI46W70y2Om9uqaGaeuICvxAwu0QBmTJU2Epb5jPXTOoOadYnlS+85
jsTYqiSzbhXTsiP6HF6rwlJPfdIArOajF6boBir+IsGnPvFid72USCbvOVwY
eZJJQHaZ0jVcEewl9ObORmNDIZ6dM3yw7QiLu8Q6ZZZYDvNTEOYFegSrqhnV
ntVDRYjrLNp7tKarDFQ/IcOhQrNZ7t0B0/tTi6KcoLmr7i04a/nP7WwOtaFm
NCvVT+tSGMk8mTjG/p+j5fpVT/j/ovWddY++/oHaFcnNNm5HBWxRyS9quQMj
Rn2Ble4rhcccZgCaScFak7SDr5y9nJA3r/Z8rOH5VvgvmWMKtMxG9mPgC6Lm
EzBFoE1TZR6eIY/EBIaiaA5akxCPnebexoJ9xd4xLU3gNIuUgkYNzBK/shpu
848axAyGtCcDat4lhTNf8H/DyBtceS3vFGtNbFFp9JQDlrkE0sKyhWn5svST
SrBuUY2EBioDTtByLC3HEKrMham+3R3IM4vUVWjZK7cjtdxHE+Xd2FoRlICk
gmCWga/0G2hhQmKr6+8oHkQugyUnrtpxSuS3s6iXWvnTJ/EGHbSTH1XAG/vW
s7W5ZtALxpybNdYLbsAOE30tLOp2VVRRDqkuRJaj0UGkmhWhyScKj9z+uZKY
oeYRaytH5R5fzvY01ycjfQacmKJf1e/MBAzLyPhd/FMvYtQMnBw0Mr+g7I/G
EoLCNjj2/hI4XFemyf6CJ6HkPNSEbnooRz98weOV1KVhvL/qb9kX8XGejJkw
F20mJLFKBj43vVwbuZ3d+j7Hlc256M7ZWQR+LYy/ZtLvlmNQMwaJYwQeCycT
onheknFS6FjxjEliHlGPrEMAtSECPj/kblUTUO2//74y2LQLGnU9qhR9Vzzq
TmeYkRChS+aQf42aV50ZvBwpEdB2PDls/zhRR1s6oTTkHPAV/7iqUoErvWsa
1HUTr5UmshiKqDWzQBg/3hYPSvewF49LYqv6ey+9TI1EzIDZGaJ7b/7qtjlJ
HfNWHpmTEPzdSOW/g7+yYHzVYX0sAlRzQcbbKV+2kWWR+5E/4ti7R19nfZE6
1IXO4roAdwNia0r3AwlRlLXJz792QZ1sULdrcruYEkQhhTXnvDjdjdgynWw2
lg+W7LZ3qfn4SWxyMg5OPm6/1nj41bGaQjfZFU5mR1oVIS4LKWlnBFIaoc7J
CG1F+7bbw/Qx9oWXelYREMK3PwHFzsI9V922vzFKvubwKbA+y0Z8rDqq5hoU
5RLwPBBJbTD+VDAteBiZme7ewMpPoQYCpWxfN+w4H+3rzV/SdyfoIePCRN0K
rniJURz4C8i7S+vF5vvhlPpn/4ajeRoln4Gz8PRZ/3cgH7N2uMVgrNL7hMVU
i+HrPxel/Lo6E3S5D1vlT2WP63WIMUahX6A1Pho1Qx8u/omwRwBJQlULAm9m
wT8B8xraJwfypmOWZmbtX6G/RbcykdMntNs3HAiYHITAcQ7f9ufTcM11RPTP
Zr9dhlhRU5lfCtm7NKe3MNMF/Rs2A9ipN3LwPX2oL9bg8CtJJAuqlMdzkWaP
M1Temlzxth1Sd2MMPAV9xCv+lpoJK+WCtCnkytdOsjgHadKHUjXhWN21YAl3
njju1WwGrNImvG3GbzyYlauxwWFnbVr7fWP1SM9jygIHVqPREpIeT6Sfbur7
J0a7SfsPuW+grlAK7eYzAdUph5zYNHXesBoeLixbIcfU4Gq78RlF3yyT6a9I
oe41PahggalKBKDitta8LEbexXKhaYN6tR6IFi4f95KWX5tAwfang7rot/GL
CAhO72F5eT5dQQJ7dfeSSS9MdCIJxP2oT4eYv90Ld5O68ZS/hcruEMFMR55i
8cMtJTRi+0WjRzS3kCYYJfzUMsCmr8LNDPQSiP8pmOnRkCqDrcE5/H1ZvOzG
s4RCJVV5cnT9UhKLA5ErhmCLLCOUUXd4gZEdmWRQbabvnICBsjLpNhhqaxVX
/sWXcoLC17hGVAQLYVSz6KWwYCP0prIZqEJ8JOxNYUcgxeat6L/wpNZ2DpdR
y/fgsNc+Gj9x7SKm2glKssEqs51UHefUGjA0wWn1Jcd5KlAqDsaJGStNnR+t
EwM/R2awBKgy5Oa6mhcMadawE7Mmb/3B8NoTXHieH00RNtKNeu+74ZbDnsU8
HN2bntvd1Nk7TWYgx9hT5GxpG0aE2RCsSMSP+GSkc7Wb4crm5jqx0LZqIYan
/neYZpe2JANpqjpDvk/jeIbLX0SqR5G/hcqs0qlx27Srkk2GsLn8rKknWrZj
wn6RvbZjiYcGsxSPpLo1l2fHxVyJKOOehbpM99UnBnMcIFuHcr9dU7iCNr16
n0ZzP/RGMs/xlO94PeY8CGSlmctH/cwS4fvUOSpiT8+isvYsTJcUG6/dzw2O
/C3qED5p6d9O3OBFrKoSd1Zs/n31nAHJbAcs1UtY5/v2UAIz3pryyl3Q8E49
+3BoedJtFKjz8EqRpUr22YsrUKQAMTt0bMSp7oxR47KdgLIo6Sz0zbe6R+oI
Stcxr0T+l6Z+y5CwyMEpEZan2ET2JFNMRs/pjnAFWYDueg6LhIuvlGl8VnpK
IEVANN3H+EVJmz3G81NhP7V+V2tGzTDpgdxwl8oyA7oo/a6YOp9QVpUeRqMG
sB8v+hSJLORALL+98RS890k715lbyRtd6cq96YJn2h7YNgkccQQbk3FUo90r
ip29h7dfz/39xNl/Cg7cdN8s+aIEtq4ovuesyRlgFbRlRfJ9tB9BmZ874w2D
Y8ENxDvT8/gXUmKlYA1FCquiixcM3MUbO4S2wn7x+dbhb/Ouopw+qFd56R06
UqE0m3HetD4rSDDt1GqlJgFaSBhOcpTLKgfXmGPdWlEKxHy8Q17OHQxNSe0x
YNA7zwJ5N7Ylp6cu5TooCUH4bRiK0FSFuHDDjMboaI1aqOL9EBBLWYXGTK05
zfMSqsQOdcVj+jMBDzHcdwacPCEXFvqtnEB3PEtU33qwt4X7oHDDrWWXXw1A
ZKBl9JrllEbfDrKABPGSRKI0HP6UpDHa0TBUD/6zF8NEN8wGvXQdzRDZeolo
pvmPFYGuoaJkrRNNmmkzlobownIuNyHrttqdJV2sN4Fz7cFz0p8mDzLSgcy/
6kbCyWYeg3cSU6mQVLX+m5Woa4byker5fN62X12kzKulMhzWKRi/8ImB960R
hhozEdrouUlR2GZ7lx+VKWJLQFsK70xeLBz8PzUD1nyZE2bPBsD1u6CgRzjF
qmvGcQ0Jq1jr16MEfY8kqsuVvInjif7oPYy9MCPb8/ajKNnEzjFaI2HLwQQv
qWZFhTbDjl1GYSpVkgRQqjYxwFb+AXYlADTwOpNdZOUzPkPMbgvDxQWAHXpS
jxbgM8fKGfgU/5HN00Hli+JLkJIcnkBkTpC398cjbC3vHCT57HE6sL2Uh/l4
ZI8uOTIeeby3ebUqd6Y0R+3K9reMrPOhL3zFiKb2fYD6Yg2gpu6Y1C3wUBKa
KJ7O5QT5DcjSuHtL5xxauFXY0ZHiaALkBkSDBSYel2Vn55lHG/P7JfktXdYZ
nadG159YH2qo/MDN114K2Evz+N5CBuBzz9uAIaiLCj+F4MG5ItlZ2w8EY5Dc
RfSge6PdnxKIEUXLbUSDaJ3vVUxYCtS01ofXwVrWVim+cTlYKWKBYgrP78u4
YDi6cD6RaohqCoYWtbcBUCc/LADQJAjHdUkmEx1+M3BqAAvGuRsRQFsROxRD
5bpXpuC8vVGyE2xqVt2oY8Ph4cP64swJyUxWFh7DwC9OIlmfMSWiZpLpIe9J
QnJfn/EXbvInnwWA6RLcUb42Wv1zA50WOSTlVkkJGLBJHON9R2ytJ83kbhva
UE3t4xvmqnrwAXnaR3dUzZHPFkHAIqpMBXyJXUk8eoCvBIAViUf5bASIzmcN
1A8110epS5FpfOVy896qd0vGMK7FNwYICi2Xgg/8NLOypIugtt2PaOrBbWqB
iQ7AzkL4XEtdadww8/JTGPvbgenLcECirgZ180QTxFrwkeHdQEAG5RXU+Es4
VhgawM5C9YDw4ST5KaZQfQTjaPjJTO6TJ9NA9KgAftZ0NRaMk3omrE+L2zr9
Kf58xQI1OyeONz86gCjW/pDWuliney5g0fYL6pkPx8KwDr/pxv/8aLSZhYVF
CPIbgxcSl16cdiomVuyqZ/0nLoYEJh7p4lwfJWfskSBVvGh37JhaY9A9skle
ghXLVGypCqzs/Of60iKzbM9S0IEgSYGt/8GkxhNPpVcT6Lv3jnCRKmGm7S5d
l5a23rPs5HDa71I4CPSOjMWjY8+YqrWWHVw0fWW57yitsbaVP5TkbwoTYRPq
5wXhJBM/dQ1+M8b/mC+nH6+Hcn+XWWCqbKu21cDHJm54Toe7VLtrse/UB3uO
scB/HFa107OblBujzJMIYzAUPoBWweMhqdajLp4kPgmNhfK8ZhE20VK0c/JE
1BOw3xHR3t4I2/e2He3r9hEVn48xgpAdrTVNFi3EWODHwWy4dj0B1wMQ+vQh
eKJgDuwL1Cm4DX7O4AcBeEW4h2kcJQK9Zs10feCuSFWHzOP0cUeV6WZj1kcs
uRbWpJqAEhojgbjGA2Q1M+FaeMxo45DBmuaLf4vrI03MVtJvDgXJg7enM/GL
HQN9kZ20d+QelydK+yDbXGUjKnsrCHQwbUT0U9XmfHCXy607xftKu0GJBrG3
oL4tr2f/HQimkIl3MAvIW80ZIYngYItN7xAMDduHhzaD93rF+xzaCgwsyfTh
nE2gfk4SPMTPrJwoD6jeKsdmTeO64KPjaGm6lz3Y/DvC0ZwPcDRuCeo/Ickc
xcfQmNjCUzd/UmtGQ9Rr+H3U5O/yB8XDIBL0azgABANGwDAcORyOeHuaBxZj
qdQPf+qkfApvs6b0cxXdDgX2qOQIvq2yeDrN8tisiSCIL+CUc2dP1RzDNJZL
oaQr1TF/O3BIMB4oVPiR18UD+xDj6OeldJRmIkr71xHT9WBQL/ChrdC1o+po
rUL7SFyphT6uXy9w237d2DGxrsZh10aAbog0JLmrWoTBCS0TgIBKK/nTugg/
ETqu34uGqX3ig3Wyfr5qouFi0u+QQvh1MTbPfDY1RvSMj0yDhibAq3aDIWiN
lAW1kP8ijP/t7mpc/yAOkizjQhC+DGgEHKv/2xWpHZ1op/wVuxufSblxFtJC
gGdBzFSdNJFZx2Y6olEg3/cjchAnTjt2Rd06/IdxkpRBcwN0P9fqRbmhO7aB
WNFlpnB4/ZX7YK6PgCQXT6w4lYdwiweLlhoTFJnDeQM3fLCPlBzhq3fCYIV3
LfQGwQnMCRTQHStNql0DWd8mKxuIJHqP8JuMP8XJdtbw9f2E0zS+ubMTHRyA
E3ilmhp9HnBwEtGwV3rVBPMf+9sOP1QeagOIPHMijhz0wq8rA4l+4DeFppjh
Kcc6L+3oZz4De9fB4xEHZOm4WxPCfwdinOuOwJiRl0dpTCAHWOsCFveSHL3f
aoOUv7SR9RC6db0WFTlkUGbqDjfuxthY43OeYDyvJec2hMZdD21NfQCBu0so
SMjrxP2v9WX+Yi4d3fwD5BQpzd560C8yJaa8uQO2nrp1tP55Vvxx5nAaNJmx
t8OZ96x0JP3YiaXxZdkyJALAxR5pp8eLA5ZWjtKffroupMITA/v4uDxVhwNR
S2VDehAzfQGTJWxYOFqqRjj9cjugcScDJqGZOYL10EFLCDR5ga3IbYNi6if4
1EfoJv4y47/htDhtCQq+pzfDpj+skjXGZMzTqmNRvw0Sn/tCrILex4tQ3MOo
otj0x4c7h9c6y4SABfcG+FpnpX4zv5pzhVtnuOekiGQo/9Mh5L6+c17QkTJf
8WnbWIgczl88E/iTsrzorfJVmnFu1KxUJK08C2hNGvUMD0pyS8Ixq68ocajp
SQPqPnNGHe+YeZtG0mZ6tr0uQjWXHZ+sFXWoBOJrPVjGs5pqpigvav5ojv24
Ct4P5OJT85xT0zhdftc88YfzYXVOtkT4VmBW3Dd6Wiq3Y/Utidli12tGA6Gh
U6qTXM4GOwxUWIHvkPXGRMsFnSwsf+CmrtiriyUEigrPW1WK0+27tiE+apy2
YV6EMTfDkSfxIXh2F7qzW19ipRfS2yK6qZ643KAH16lVKWDxsy40CS1NARw3
v2pettJetRvIC1YIRt/5x0OG0LBBGPkY0nreXy7LE94Yr8Vl+0Wm0NJNt+qQ
0vOSUQIXyRY7vekXRTVJcU5lMw3iifI9IiwUnJWPAk0nY2Uw+XrZZngG76yj
1xSlNC02g7XlGqkFN/EnCNiwsYczjHPF3xrEG7tCuyqR/BrmZXxIlCeQ83/Q
hiUllEEMGKnXORrI30bl1EaJUBzfcSYgXXMPRQ3ueIP7VNge5AhtpxTen+Id
h/cjf4alO5mDIoJW6e6g0sDLEGnGD8wFt9+9ERkWCm6vIGmocPBHK6ns27XN
AyWoE7bGL9L2t4jaY1xTBjH0Uh9GJI2XT3EidEPooQXb2IKJrT6qjxSyn0US
+fL7gbwK56c+z4wgct9eSMJsUuj/f3MVIb+rmnbjDDJZ4tN4veeTp1rcIkRk
wZqT+RjzMXgeuIyDFAR7pcXc1KDz3mtiFFTFe/uKE7QCai/IUY6pDycNtOmc
HPKbC6nWhVDDwqsgzvHHR+cFZWUSrFZS/IqJqveAYaJQZvn028+rf4EEKkKb
ZXUF1cH8fJ/vCjGjhk9NYbIyuPnGUypin0CcI6fE69IyC5AXtb4Lq2l3IY3z
vnlmEHTOqhV0ewskqdg9+L8CjFbMMa9g6+b0U1cEQ9NSmeBdrEA6s9bNgZKJ
Ocl/JVEPQz+35qO6Bdp3aUPr9aFa8n2NggMewhbS3EcYgC67bqg2iUzi2mYF
BrxQfBH5Dmj5vep3pgiSlF7EAqSdojstcLev6/lWU3BBimyrq+l3AknStIDS
jaOedu+9pWMTnKFjhOR7h2oR7a1IqMzsZcGVgFCpXIGzUJn4Xaag4hpeguKM
swJdcIwsvVq2xKjjZs1k/I+wQzs8EXPxo+roEjzwx/yRLysPLiDuYu1sWtZ/
JWQuLrX7Ay5SREWoe5zQCC/3EFHWGIvbJxv4w4A46ySGGnSxrMc+qF9j71mJ
J6CTHDXjGZ82wvsQ7QsNkSOPAzRqwW2Zq02a2waTBbM/SZiIULpgeY8jxKEW
2EVH/unFFh/5ycI5yN+EQYLKPSkmvHsIAczvq1iKcGxGxl4orgsnE0Gg17E1
K/MI6uerKeSzDoDWuoDCT5BXckLNJoyUOT3pUUBh6ygEt2DUQ8LsR1zvNUY0
fp9sq8m6VjF7VrLvkO9tWfgxP4jDRlF9ss5vB0BC5LWhLp1jCCV06aUYs90J
tOaCR2g2ZvbdVvjZk7abzLjBdJXoalRTHtzDcpS3mEtjAjK7MSs+7ufALq7e
gGWnTXlWlPuTPkGQoVhlPvL4hF5/nP9HTeu60cZjCM2/JkkY8994PI4UEp1v
8GPBozkJq2u31p6gQJK7sxVGW36AoqrMJqzQBSSY/HZMSAsyuu2GyPJH3vwK
/gOG1XjdMvnVa9uUe1NJW6GHKzMVYHY0Qk6l13gth2m3psaWJuVZC8kV1+JG
ahRtTYZFvCh0ICS7NPvIJse8hV5k8WR3vDJ6JH2Jkmi/73gaN9gSc0ixAk1A
sm1U4T8GWRiwJYijFkzNY7EbNTJUbR0dYxIHDInY/uALz6cJRAL0HVkK8tBJ
MxuXAdolCP39ZD1qbmvSYYya1lGyQDKIeFKdDjReokOlZ+mvzdwbVMOEXq5L
Iat8ENDAEbVATM9qiCOLO4EiADKwp4WHfJDarIEdLLk0hPuqO8G12UsrvMqT
N0u7Jm/MXOJRaPFFOQVyETLrwZWivnk27r5yE9kbiBLfEyV8G5uicj0VQVhn
tSXb8s2q+RtUrSxpA8dyOSpOvf3ljp+x6tdfx02U7MHreAOIIuFRr9ZoCBLj
mRcfl5RO29FU4t2B2bG8Mb+Ct3u6kRxXULax+Uz/4ftp8z4ufQOMT1qeHkKg
TuDnLnhK+Lh454fafDScbexBVUwr+k/Q6XEAle8+bkrXg6GUAMmBYQ3e2d9g
FNSgQTpQJrWkI66emVLWmx9X3VfTnR6AI5j4t0479HBNM5AxOmngDPIRXbZS
yB6YnvuRTgHapksSxt76PgCwMVYjSceJu7yz9S1+SwKnRi7BV9psoq0zmXEI
rwqyjTK5lI8/oMIPPaamChGn6OpKTFPJLsXQ80PdG+hwAYZMrs9uIofrLeW1
Ee9sRpMPNib+ZWQP7QSWzm+uW/7B1VpLME7oQ2vWsQfaEklc+ePk0aWGLdNr
pXNHEAenej+l9NuaA65o4UqIferl2YY+ks8rx6bw/kumYIG/FQHpvvNVFTbU
x81XO6LpP44dcqhZUn7fn1N379/ZQgGCb4bFwlmRZ05XZ7pPtS0y+hPVGptW
ibts7jS17TmXiBzq5AzDUWemez1HKcGxlhsyIO7lmfmXKX8mkBVxQ67zCgR7
iIcoytrv1MTAswGC1YQRInSlGS6mmbdQ7M3dnX4jTIOHI4qT1EzoBI1ev9sg
qSlQoTj0ItsZogrkoTfHpqWhZVE4muqujcte+nmjgGo9pYt2CiCuH5011yXf
vmfzPxqcArGc264G6zb+xua43giOtiZnkDlYKK1y5W7pyKICIpmy2oR5r/FQ
WOit1teGeNJ18EQLvmxpgjzzIXPpCX/lf0mKn4lbrxRLOhFmIRE441llwGJn
k9QrqENI/zPOswi64TQNnObSxhAMz6p/7L6uxRcvbD3ytMoaIqcoC/7mZz9+
4fOEcRnTNdHbYqc/IfXF/oc/R0vTFUGFkvE+5O9m8a6VeDwyt2nXj5BW5S6C
P5T4cc7Yz3MDwB9goetdNQJ9asHY/46E4L5O6KEKCa5ptm0GGrXSWXXmOceH
uFzJISltQJPqa2YwXPq+tB1yeejx3WsCITNUaoKkWa0EYkmIut87d9yGKL3M
wa4wRHaXOduk53YwqbMcoECxytFVUgeOvB1yZQ/q6dcupAPEhfsJUoLlE2uG
PJEwiCbIwuNEYQyPzqr28iSQzWdnysEABuNpwAN2BlVWT91NXouTK3TTwhMI
BLV0fFr9J22u9jbyqVTuOyFFrC4NlX3ou6b6ZAxEhb3y/EIXBPplgnD1Gqr6
Ql2Cd4cQ4h73Qw5yjZNHT8sCesdHqy+1tWOzeBjXaCLSb3vaQoTdlzREGTv/
zaNhlrBODST4CBUsspCxDebbGtEZPIKnc29dCYYH1u4GMIJE9iN+tOvmRThV
fXwYUlMpuLan6JXoM6XoywDjPM2fJ0mIBl5O/Ds7dCvNED18oRwx13y1V+Tx
QgRiITeWCfyqQKOLn8+WLZttgOKdegMa6wih7CaYFyx4ArxNWMQI44MTI3oz
qTH0F+fehFxxjVFv2oyXb+JA/mNGEnhOja/qoMKHQQf5Wyugoo9iFytBFbmw
9bkfpKoTekAzDk9fpwBUnUyZAqqXHPFkcxCOGfIJCP9PQJAWf1W0mbQgK/Uo
4vPCRrYLLYRwk3kR6XkumdcG65oBI4wU5v95m9bToiJE7+uUhDwXcUaORZCd
DHNxqvZ0k/nguK8ZZeHIWwc7MBGuzAJJ7PZF1hxbu/k89lTpJS0uYdbiVTgS
4ZcpyRLTErTF2oUjuuJK1VjPSq29Dbwr/bmQwg+5keHoc9aEjDaC31rclRK3
1/VnO/nsXgmNxwHPM3/OzVova0fk7WJHMRl/oP7pVbe3A+u/ryPqZnBOiMkV
ItnvHSYQf5nE2ixnCuUUF++Ubk9fLOna+vindPGNfVIMlXMkJAIuDySryaUx
dJF2O16G2cwkXGSGaqxKi28cnpBOF9UCXsYiJtxdCJMZcl0JM1lEPOr8BJc0
KykfpJQW3MVHcj4o+EEc8m3iEdJQtFqiTMlx25SjvQ2H6m5F+DkkQYcmVP3R
ApEYhDFUu36hyUrJfhBKvZRZxxGgCHqxEWOrQXT+3Ws0BCrjeIc1de+1nWgB
30lekNYIQ69AoDYm62c47drjwWAMJZw5Qmf9IMpLZyOaJwAdhOQd6bnD1bTi
lZR9jNsduMuAjtNq8Iy09icCrn7FYAo65pHMPZ9Nv+iQ/H69KiejVyzQQV6K
pEFa8Vfr0UvdeFwLPL8oUY52ubLxA44wJW9I4SJKP8DeQGUhFyV+YLH1HgnH
pvJXn+7XJi3z7UI5wUAkd9ocdcCDoqTaetKRCadnJBDrhccGlAUhxjSmRuNM
grrJLZUBNiywjqJP5+i2XaVA1plYwh/B7M6/Xik680U7n2w49du3sAzQk+zc
Eljn+yKciLJUpVTy6NTIvy9H2Eiov2ACEC0+aYKO8gy+myvNmS2Xa5YctMzE
oJLFoqkPepkbmj/LcHmKXSY5vRMSubXS/x7TEBNp59taHhKAUPmq3SEjsE1l
ynXc3oabyTbSSPblnAbAWZFbwPkybY6+hI11vbHuO1p/kjXglhqmM7ixAdiG
ZQl8n7D7MVhCTI9yUox11IUrZdIZQNFl8kae7+BLcy53FBYv94T+P2NHp0uu
UdJdQXsJRV7iYosULejJ9LSjz5vzmH5AgjRb71aqsTpKPDlmqo8RLTexV0j2
3bDmBDN7Pbk/I7rtumVnNEXDmrAC9qb8vPkCt8V8gyvXXx9k6ybSq09/09w3
OniuqTagetFbI+uf6a6j49uX1mLN+4SN7eCYyyVIspJe+4fZ5nKi3lJ1P3yY
Tgx7FV7xZmXlohhvmedRz3ve/kzRtmfruZHR1cMGg/MLFCwFfIWuKnhXruVt
aUt8UC3R2Rx2HgADqLcVdZEc3KHoKKlo4aYRncidSrS4evJKdWyX1WVSG6iZ
K5qSjKNr00/q+puet7BUxhg5drUoECnx3BTUtJwMgnZuUNlbpXFzzA1pSjEp
Li2V00bBWWfQyKuUDSAXIMc+dOBF5kw7r9JWuo+wXatsnZPUTgr4ghRdEc9E
xdMOjTDDJIxvzh2h6K2nya8kTebIL8B2+cZA9M2dLi+3vU3q88N/r9EUApip
gzqruD1N3w4n479S0BvBYvIrHEuPNwtYH2sQAEB/jK53x7dmQo3D/n6XLJXr
yZB/3L1Z2N7zC9txpR+UDIeIW91zAJM1EN9usYYyn/3uNMpz8x6UiQY0PO6O
5aL/2mPcbrhDLXxgUHmrBv21xuChZp9F2ShhQSrEMOzJlUTR29wT/Ivq73xC
Kgb4VJqrHabRnef3gfOWsv3JRyiwLHaxGWFmun+dPyC1UteeQeeGy9yGzbGa
zpTLZRefR7GQ51SgYUkdVy4YmdPDLy+CRD10T/BSpR260LiKp7XQ682LFHW/
2iDVXvswRJkm8WpcX/y83lhF1xcFLLWnUhjQ+HiGre49E2vU/FACjTke4jyW
A8mqltMpQV1fzPflNHCNpSc1dLsYulvD1JSqOuFftzSgufr0kgNm9vF4RIYD
95KnE7Y6okEZ30CJZ507rvauySYXb31ogN40HCVl8HtTpH3rECmZ3+V8H2rl
FqI6b0i31xY+OBve3qA6cF8Q5s9ivTVIHkiZV85yw1AdpmUny2ajlKTOXtqH
370rizS0E2m3dLKOSMxN7YNgC6zyFykMhAd0ea9qDeS2qIRHlOOAoWqrOa1Y
LKQ0mhw6Bir+fkNfo4h2SuD93Dh3jDSaxBrmHmWcWaCwxESVqrs2CGHeCiFU
Rt8aHIQd4w9vT+AMUJd1d7N2F58pRPyhN1hJf/c2u692pp2g6ZbkhobVEuaV
mZhLfrBhCtgztt+24P/RHG9ogoI+e2ukmNTy+r8BkfNRagN+aTPCxRjqPt4k
bIYT7aT0MCpqS8DGMyFn/EzhVaM4g60HIcAFrpAV8kUKVmTOiP/Bk2xEwnNC
lcGExOV3WzOnsQ9xbkzOif14czEm6hAjKYIqS/JSweedOIliGa3EGtLmuIdS
QtfwJcAT2aIYGjcnDRW4BvYiGWw91BvRcseNZVaAUo5DBhPYvaX9oK8UIVpU
Ga0LuEHGLFxmkRyk2tUYgLVZ6I6a/LZDR9NPumsuSmsX1A4ic9u4oR+yh2uY
rpB063maR0ds5Ey4FxYDXCPE1UXzX1sK6oKmR4mJdLzWV+BpJaR3fY1pjh16
1dNzVWoWQFGsEGCKXkajZQShiHhHFJhZ3ep1Kt04b/r0Lvi6l0hgGADoDPef
zmq68Z9qOUatSNW48VteRvK+tJ5gsVmJ+Z1Sj9+9vIb2zopwSXyhKfH/uyMk
/PlUmEUPJOiaE3QFowb9v3CHCt7YaEY/wsLr2o4s0iJKSYQe3HHAhPln6uUD
Sltc+Gru8oH15dCoHe1wv28JehMrEovcUUs/J8Vnej04KPGykmNHMpOF+PRt
rg0t7El4NIMK3mZ/OYzt6s0v9v0R2dzUPAVSKYo46w9ivEeVp5XjMcaZyV4z
X3BRxPp+EoClQs0UKL0gtA5tgI6m2OU1MFLkwVUbs7ajQq7pdamDQOTfVlgd
4PXsNuaKAT8viAY9GHIVh/qVEXL2P9EPvN2rZn55qj4+ME15k8EtMHLKZtM5
NoM5YQ9PFPhi83uv7NBycFkOSnZtIvELwkPnQxCTGrP/FaJosk2GkdaxG6/f
aZT8hijtHvDFBhLuboLvesr8pWEdxnLfrcA//WwZb8VLUDqXI/v+/zZ/BBSh
oKn3Ev6BJcuZydJeQSDFZu4VoOedhYm8kWhTttsw9m1imCaqa1LayggyueQd
uVQGvaTG2ROf/ylF7zTw5ST4gOedBw47eq8hYPBmkrx5R8S/z615CKRru4L5
057qkRSS0YP2mGIPGo5441ovrerOLDfBgW1V0/1SEZIjI07NqrgjbOUzUO77
eIw0CPoGmNn08+Kp2/uGeDdICRLX8ry+KaAQdtZzuXQ9vMCpcQBeRQNvNK03
jYcussZj9cJ+/4LAkF3TV6u33qp7AT7H9FcNdvqJsmGBuAGJL6B4EDKB9N//
CZ9ip3HxcVRGB93zqoYFpPSpNUU2e+kSR0N8UPZEBp1tFJp3YP1VYdO5wEHf
CKuwnbUJykYDQrsqCwmIlOpW2/KcF4MZlB7wR97J5ZsilBtive00IGm4wO1h
pJuaqI5lw0M1gSRSbRoGkE1MeRWL11J8o5T9L4UqGAP2fOSawfEs0+pV/ImV
X8u0jPH9dkbBBSnhQKURsOjlmrhU4of0kl4KDHd9kRc7athrxVEyusJP9gWP
MJG4WZy5O1WnIPMB7habCK8HIbMAJAWzd+2jJm7A2z75Q878idc1BPHELZVf
Nd7ld6jpQ1zW1ubfB3ksC7MKARm3ACJ77FHu7U/rD0/pp++59L9LFkUaNPqY
0aBAHwaHkUzZEZ1b8SFqXwz+UZ0r1Mhz189gqNghPAZDApnptjqQh6MCLuuy
KLUzummMEK0cW6CcoVvK4Bjz1yskjO5b5DgVwRcUJdk1233emxapsaFJ8UqJ
pkdPhZNJIT+EsUjikyX4PLtvCTKmp6llz7ikjiZnScteiSz0ZxbMD1QKnyv2
CKCFyFGEBLAHznQjzqkAarhe5CnYmEZDT4kpjDs3RO0KqtpkvuuB53g4UoCk
p1qL3JaYy83X4G1xmvYX5h8OB/V4tqLinFRimfdcj9qINgpXwGQJNRzAHw8h
n75FBUqqjAApxCnIswvgv7aPhNOfz7V4k4vtD+rewt4WjvyXWA49RT/IFjSS
PVN4GqvjAFsocQjmOEJydqSDqKWiNinMs6VRWt8rikCRAtPBdOVr9S/jokb7
vhoupD0xSrKayv6V+XUkMobZk5ZjglnwOcNfqaYzd8aa1WxGZHklnRPUVrqC
iSlpIKvO3oTuyYc1MgjCH55h8GlKxj9IXrup00CjzGyKeVHf8+NoqURBgwpb
DkZPP+bfUTZgQF/ezEvNpeiE6q6TRn0P0Q0rkh+rgD2+uXEEE1vfM7oeKOKn
w9svArMKPobf9XK9Ly3eb/acf+gmTYoH5nU6cT9FW7A+1RZEGbIiywmbyDUV
ySbQYBqSMVQpNplQKcsCFVtWduEjq8rwF3btWAvob5dxbhFPvPpjjc0dwztT
/7zAOWksOjqNmrMrGF96Xkpl8vrEwnTYCsoTn92S9xzaFFtJY6ORb3GFo63u
cYpWGOArpiG4x3FHPaw80eeJ5Z3LHBNcuM8ZPb/WVk/cn3fxBde3exlpIYvZ
rrn56LIqlYP5k+78/B7AXI5xntz5ObOuyviHm5/6IDS7kiJJL4ar3UY/ph9J
hexylSIupIwg1ZgVIylzx/JH6FlyWwqQBtJ3SVoeebWdrq615X/9FQnGSZ86
bONN1a8X6KvkrtKRNhcOiM5A2yjGExyQJfGTkOatmCTgkQ4TiCIJU0bNfiOn
rkwZzo3llPuGulHdNsMgGinAMJdEGipqvTNPF6vjm9WpUF3rhl3toKDpYTuV
Om+sF23NlC7pF4BVuGIXn2zSPbyf5Z7trtSq728xA6L6v7N/krGkXRPORSBM
GMuerjKf0jrQNIQOG4dX5Yfh80eEAIV7nObR76fnJQyRvfMGOqm/ESbmdZa9
fEEtpQc60sgkWkFI5ujoPJ3lGfyU567v79zGEzIZcFUPe5pUG7vnlYlZdilg
SZ9kvfJJomLkv9ofR0wrWGKQDCUVCOuqtS/ZHekE35xqEvUN4k49h38EWvuN
RTH7EXZdJKuTUtG2FrgI/PF8sQora3RJ5koPEprXEaJ3e89KqNdL9h+G6LmU
Ya/F9nx7eMoxEtdvbyXh1i6G/kxHAAVRzmWc3V81vnHfcgKKWmXSGo5nevPJ
NXo2XBvuysHx9+5CbhT3ZoGSRAv008+Ei86ZRQHD7Nt9MA2HpsqSakYsCHLo
c5aqzX1tLh/5eMy6ng1BLMGVXSnHkzZhHGF4RDjEjUf/ZMngS879oaJtFC86
doiiTO6znahkhB7D/7qPEaodvSpSpZU0IGcs0X6eucX3y9FAqB0kYASPtLTI
1dfllL34JRjgKh8PSZXtrDwjMv63ZhjRrDaU44B00eYW4neCfTK8kvrBFO+l
RzkfN78kxjyKMJTvsiSsSq+noGXCNS3HsFvR9YLMDIfEJr1dwEJE3Yp/SpFS
Q2co4z0VNCGpt65QQIGtUmeAF57wyZD+eTcOrmzeUaUN1gJek5+IGn3pnPYg
ZCXHAUUvx7+5a32IvIYX2jF/jHw0iI0/yhv5nm3qk41OdaSi1Kpa7LnNSdzM
rQS2MWNBjD24DN3T8Q9Dr2MdgPCRrvLVQ7D3MOBYW0ILtkVAurAezkHu3xom
Hx8WTq3kDZiWcRcPo8uNT2eLW5MmxCJyyRZhIrmZXaM4NZDk1s5JuBjqW7fQ
nbi121WtKX/yqa3Z8+T9mb4FlmE8BSvqys2yqI7Wg3WbeTxH/7LEm8PGmG+q
lii6n/lEuVFS98OERyuTvrFCdyxr4DAMUfM0wSIXtyCN+kmrOHWk/osgk3qg
/fhJMJkX6LCmBT/ZZzlwqbsWrPauQYCvgmbvREwvRjbznYtzq+89lhydwz+i
AT4ZSjyZ+SZwFl6xPhTtr7Xg70ZipsJb0tL5OsQllicgEd9KeKeqw6kt9pQD
cY0I4JW1RBTCB42AOF55IhGNAThNsiVUNx0cjODAJtqX02Ron+ODTie+Mb9O
Y5hLLWgk5g6UxeruJcwfyUvYLGcEQExkc3j23rcCz2360MXfaZ8Ruwh911Xg
pGszjzS+Rzu/97d8HyyS0TxHlw0wQoZm0N0KDmTVQmoPKwFoH2RPSfzBuGDh
6o949kqyPlRZpYc4LCxjNPZogVnOjG8IxnPhG2kzD3YDXbtoMUR3t/qqn0o9
i6VYESMXBrwqYRvSFlOylAdCiEg8sU5bsd57GVPrpf4OAUHPvEl2skgXvyXt
Ap3dKScjGqnsmTvOkvbY0J127DgOb9x1Fqd96ogy/V+CwwMa9LiCiENXauM=

`pragma protect end_protected
