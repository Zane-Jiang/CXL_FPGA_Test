// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HSnX3G8+k9Bz1/YemTeSs4pnWqBmSpWixQMkIp+7L6KBtoKqywzsSt6wdYVU
f3IyVGOm/C/Zh6vfi3iaiCQ8RJOAK+a08QDShVjUgn4PZVzoviKUT357Q0Ak
x92cFWkAu4QNbuXVN+3u4MCiZ/KLGFmaXBSK2ymg15EOx6Iw4voLfpHfqtBn
vr5KLRxz7aVCPwbdLb2J+gKUk88Px+LBZ+hfcr+G9HXfqYKoqCDY1DmoC+3Q
3flNY/yrSjlukxrxEWGvt0Cr8Ous69ituEzA8NGTncjQy/WOU83HDR8diRh2
hib51LaAnFORpuEgZzTOk4KfgEJ6auCplGE02bKG7g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LnpmVuc7U38wJuA4OJjbsDuRcqobi+mwSJaiEVLUxIG6jErvmxkrmZdw/nOF
F6FRIORBrw07oSKwwhql+ZsNLkzEv7p5ClD77zz60gPDPeoUVgHhhFok1grB
dZFAB5QCOcH3ZWSwSGNLH8Di9T+nEU5qxe93PgV3JiGbZ2ab+6AU2z9yNf67
Q544MZ/4i0vlypYkouPdO2OZ+H656G98jdrraaJaAHIfN+kxrOGHfkGfM1t6
13kh2VMH7+4Xm772BO1iNB0ZtjlNjuDpyc/yw++T21oneRY0/Du+wp1Ar8/d
5CKuSRqpBzEnA0VaW/wg2VEZkfiTo4ONfGdV32nyjg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Dp8xWvMoHNEYjdmwuj4n9F65PhSfToB8gxNt2dRtQVbr1YopaVcQ7A1IGP4q
iuaTJd3rFvxT6Mj5S+TXUNYsKy5uHJxZM+UGxO3pGPcnM2rE+29EPY2hVQZj
m+vHO8deQcJCLzePvWMkOgxWgRMaK1ZmaJUfpQ4KaG1X3IAaOZdUG7sKNPC7
myUmGbJSvPW8bDnjb+Wh4x03PG3rPDACXY+0SDYFJs32UmZa/22cTtUBfK4u
HcRpGcjsiwg23/VVArFQO/n3AHpTBfRvtv8IQgrwScpWMoSJFWEP3k1F9bmi
pe711JtsbuDnWm1NSiPsWN1aQGxs0uGUyT/b9UKLYA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CeTVJXOuKWvrI+2nKreL9zHlwh0Hs4HPShzmkuFVxmiwoiIiKXuqyh9Z6bvp
VCpRwOhExJsLWYtCo4WucE12B6Nk6sgIdqBYKNAE6ljew0pA2hy3G2/2kRsT
dhJbeZv5zesjv65XlAD5EYDd4x/V7Yh0W6lat1E8IuZOZI98Lss=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
esHATzpi15YGq/zsAkx/xxzc49iu4BoAdYZkOV9GR8408toBonrulioWhW8B
cVd3TZN1pAtMh5iNHGsn8Z6iOuDEcKzmvl/FCGjIDkHjX8LXJW2oTzXJn672
RdwYTZ+0LJQV4x8wyMzC9BIXZt25ZF2ukhBnE5yjPjiMRMk9iTObSIeY9J7y
FsoNWj+k7rfx/sUfm5Qxxb3NnBBTLNKWQ0hTDJeuk+NP3dl9r0k6G3sD7zfN
ADTUj09zlkIF4+Dlg6HzGs7sJwjHAW7VjWQWtS/rdG0gk/lJhjQoAxcc0eHb
4UWTKrsOOJwBWpuHMTXlJpWMIj/x03c7fk8ubCosWyxLGtb0Rqac9lvDNf07
/J6toIEVUt7+EHEQ5Cn3CCC2f6jEQjmkKVvvA/3/2bcDcXCASWjie+okwLgH
HVbzvJ7hdCbxYJ3ckEGyXV9nDkwguIzCuCggBj9bg0Ph4OjCM+oM+PsUMzbr
CyO/NZ0HqRpvJJ98NAlIa7w/Z5XT391V


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KPFatsI3DG6+Ar5fRFz1+q13BggExVeqQ2DBTrnms9KdP/4I45T9ehW4RAvn
Ev+5c31IRXxaHKTmzEkl/vPPjm52VXaxqxH1IA9vfxtGroEkWOOMR8hcx+5H
XyybhsRKVCEnpyj/8WHBEqxsEdV/dAZKRVziWv7vhP9rEIpksPY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n9kBTJWSjZvNO2MHnOaPfHJWLTL/lwleF2G+b8oI7vPphUecv4Eu/5fMyxtB
Vmq9gmDohOEOlfwC4A/sfUKwtOTSwy3vlpYEGdsbQV0E296dFjUOu0sePNQ2
gWTda1bmMZ/aEM/3UdtbMvC2vOvvqOGdJJvdLXc3QKJi2nqdVjg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 57312)
`pragma protect data_block
a2MPaipF/YF1NSUe7tnmFwmvmXNaMNhDVGv6a1p3HKidoLkVps+WxbOv5swB
oico104BEkm+wtaiHnKGi67LNtQuE0muAI3eaQ+LRrj90oOY5QVtRmmKegfr
vd9Xz85lCiVDqEEvT7SNx7zNvuSMD1QhcqCklipBdydtx03IXr5FG+A9M3rU
LHZndpYNvoymJA2TK2Xyx2zgp2LrRBTYmTBXCSJZfyqOUFHEmCbD3wpydTtB
drYnFHzUiINXjm5RfNFw4L0lp1OYmMljXEgoOSk7nFUiW3dC7I7OtcxchQ/+
Lqzy/uHACOcmiWO3RUOHTbwHFSCs/PUqadjJPXaFeuU64YosUPKcuDzGoLDf
pvRaNw7nI+W3cOAid9I1e6K2g4vae6nH++VDhqy0bpVSistmLqewAj7zJIn9
iYBNMlwHosPeQiTkWFiW8jori9JMBVqrfcieG6GDaCVk0uFCWtmLLBfL8/9h
q+EP0iN5+oXNZ0wwMx1bKLhwgshrIyisJME/SsKC2DA9Orj0M2IxZOVJUp30
SQDboxRuIkgplE0VWt9qRwqqtpej530pKZkQcxtITW/6nuS3kT6yAMDGyKXY
e08VvhW06T5hotIRx9b+Zgvc+4p0rb1Mk9p/KToj6vzH+TelYAArZWx//dlg
WFim25LK6r+uXkZevai5c0Cv+q9PTzNQaBPVSDQkRp6HksYUEWqM0h9nNBG/
FDFqf2sUUVwO3aewGNfFix+HJ3Fui3HA8jkl2oyjNpGxnjnq1RBq7xLCpIvK
UC2nd1LyKd5SckrZhI/fBMkbdDZTNl4FWDYJLsSN7K+42PAlhKANcSX+++q2
jVVOHp3z48/guYrn1S57XwnaA3UzXm0N5PjNvbZjd6ZuQjH8+uAqYodp8r6t
dapddK2x64+608loJ/vVvSvBa0EjlaqyiRdB1vhM5IcLWrGf6KvEBkG1BuS2
p6DER0qq96iSk8ZJGy8UO2YOsnv62TsONZfIrmXQUWpwEj+ymTTcRy8qenPI
vWHLw82gKMu/cyOXY0iFfOxSsqa8nWhiOWj2vsnO+o2tg7ujkF56B8Fqttuu
8GsLEMjSsJ46zA/xnjx/KxHAmvCQumRfam2nfJi8Ez9Olq0VfMNxxeaMTmwg
qs5wR7hA7U5+7nueD6l+RvHRDM3jq87FSLpmQ2eR6uoDcsn+cuSSsEha2eKh
eYOvBvgy7EDHCnO3VU9elQ4CUJidCBFNORD5H2T7Ys1CRrHT54JwSdrpYsq7
JeGmUVrqH3WgCz5G+eGX1qW6TYdrmqBdRuyi5mdjP+gTQHTGm1rLJotALofh
OhZn/ArkhNEEBXgK14I8rtsFch8LliUcs6XG2sdNcKyaSt49k1QwVtLHsqPd
7otSf3+DXqFBKA/ab6dncuvJs6bGM6iHx0XPXwxpX6vErHzcxZJ8P9GIf1JC
NktRJDGDFunRNNdXOQTzkFcEga0EmsOvXTvTt13EtQ+GuhZNqSBlHHFQhxml
azRPaSimjHOX7c9j/QRaaJQtfzSU9y+M7T1VhVS0bFFC4O4zYXuk+vmDWK1x
/6QGEYu76LsGD4t1XJCB8temKqNBOHoEHqydgGR1vnL32iToAZinryz6AbCX
aFJPF8lxfwwwz1wKn8TCDcBgMLRUg8IuesiTwGZv5tEh57uhKARpNKfee6R4
ZD5vth7CDJM5wmdopaz7GHNZ8Xv/X470juQYzK6l2DgUK6jN3LipIEms02Ij
aQSA/fkc58hFS3adtbIX7YsaJVIbSFqcgb/Wr5U21XytKFvdgFHrgDA87JAO
rhALFukrvzxy1a3ePeMN3WKPIfGR/ppHT/HpXHtdLWD6Ne9ba+xq/KsU1kgn
Jt1SBU++Wgy0pXlbFtzqGUmNr9O13d/H3fSwtBj9Lisg3EFqqsCT4GNUAn4E
Y5VHWbAW/qY96jXULrgoB0kAOD58v2mbPYWXksVVeUMj+HL5pHW/xIxuwBPE
DwMZj2gxcHnXvDEFckZjjIBKP7+l/mwBcn8H7GKXOMuel1IIld2+hMuvxMsV
FfTDqtI4gAPFhBKpb2cro4Top3CF9fO8mXjroYiQMSQ0vQm6RctylT42TNTg
xeewoauBe5U7ZurzL5TWV6MOfwOwkvRA8MmF37abYQtguys0kF3Z2Qt1OLF9
K4yoHTqyENPpKvzjF+tmPzoEumT7iwt6CNI7YEhOd6cwOe3XliNU1KVo/MnD
rUxLR4+jjarRT9cUGrrAX9z1rRmhpU4YHLtEQn3nYmwM8TQkrXdfNlciBMRY
1HvWZnb9CYXfd2SnWwHSTepg1WVXqEdjQ/dURA7hXX8nk+VPzNQEN2bZwb4b
OKDOCSxvGNVxXSkFBUYmBhhsGIHnCQGoi+T8JktBKfSFxpmlrzSNL6CpgRSU
1w4USTXQ1pHW+u9yracLnIqVS6boWHOzrN+PFsjHVFJfJYZG8l29v5NKFuOK
L1KFkeHtbEqgyD+SmwiWX1phZ8CB1hrEFwhMOWFMfoIa/+R5ygwHt3uFfD7C
RpOHJ35GvL8996kTtcURic4KaIrYmBZp75aKeRL0SIWyKB2yDmABKBkNwkQN
t/osWe+GpQVtty7R7pSFq50FLBb2JhIrBOJCZku2OwcE/VwZxb3zVzhM+C5v
u+Kf7udg3c95MwFkjlqRfUuJ1wUwrxpGqpfkaFNMfisLYpS+aCkylHDQze4Z
dsVwNTSk+iSvKX8NkohD/Me32cIrgW9rzQuA6ZiyukMVi05muLGPEzsOpBFL
Ww4VmBuVtbLGYQryFHswmeJs2dWekz5OYl9NrhqGjxB1ZgXh8OEK66Dk5ZCv
ZUtqLsEUZx7AU46FEKwPlPGyect+Peongz5+yqvFPprkFT+NfoD5ZOh/beGj
ULU6XFrG+vk+qoVSlkfYGPbJyl1ZGzq0NhUIW6z9sx5m2CIrhBU0wY50eby5
IYA9ypFY/XPwyj8R7q88se4+FZgG86pr2oXUGm5uYRITyV863XLsG1JY4sOT
RKTHcDAexbCcs1rm7lGNHoI0c5wDWA5jLczW5XPl1LzEhQHd82YshwuVq3jt
LS5msiUyarMncDSxuK7cmif3nGnQV6RbEbAFZcuLDNu5TUJHfnmfRGHXAB1n
sCREHBn731eNpLR7R3LO4hWQUnRVGD8wfhfaKbp5l6CN+YsbtlqJ/CowKmUi
kH0G+FDeM29GV8c0Gu9sb40lWNva1M4omNbe1NViHFNGOyyQ/IuoxmUF8S0Z
Do7jPSNMbhv+0d5XXo22ODlmspUjpggDES2Z6lXlI5wP2qgQ7FG28PZlej02
NYTY6DrYD2dAZhkzH9WLntR7jfiz+218nre/zqZyiwDLaPQd9o0W7C9TZHJr
i8dHX7ZAywg3QuUzrfLnj+BHqirhXPdGh1F8+iGcVJkDPR62AIuZWqqZl2Bw
J1XeUAC42ybibL8lP6hHjVsWHmp4/q1CgdMFnlrqAPdebQ688pPUQDHpR07q
jTV1PUyvdDBbLvINUW6b8uEv9mE9pOO/X+VgTPkeZ+F3bu3HtSIBk11APpRA
8u4+viKy9jiyivXu+j4AaO4y24aDTwSobqlbhlggIffucNzwhbJfOHb36+Fy
IBIawfiniGTwHSZCt1MgJIcb9Q9y7pqEvqBQwD8keCf9aV+jt0Sid/wW7+Hj
8dDMeACF3EM73SVn9O5321iUaqQVCkcbU73niIl4KXHvhhZaGxa9N6yj0cxg
ZLVg+tfalhpirkJjuiWQ5R38fEpSeHPY/qAU3dQpTgHIknx15Gkl9Oez5Mbv
JOz1mHodrk4zSU/9QYdTz0X1n2qVj0vQHxQNjNCtLMJpwI5hPKuHIDnD+SUL
VZX3TGHJLFoiUZPo+dAPKLnYIjrfARxd1E0DjcgE1qbDMylegBMeSyy5QA2b
Q/vnOvVC2tyemcS8I5oy9aGASrqtstvL600ZAAR4IIH5sFyUYTes5yj61Bhr
+ynF6d1W0/bkqiL3eB0jJX58zPCLrblTQUPSIILnVhqKR31cvM5J6Wy20/Dg
po98duFBmWuwmcQXwAQFUmlYPPQ/Ubq/dswUucOJHdqyRVUdrrhbjMQfbcmA
fHlgOheUlK1cROCTgqqDgExsiIr7iK8QDByJzjYYfyxVFolIO4MnZdaNVZom
+qCilGKJn8lgpXQ738zysHbVPq5LyT5cC2cmI3NSUsebun20MgGzRcn1D3JE
hAZVm8ii+4SomdzN35CRDSyqzxEWwustkdjyQHLjMD2yGCF555ENn+pYzr7D
s0GNAByzOCk0BXYGQxFNzVLp9NVVNI7d9aud7myXJBWPDoloJiJ+to0ht7iB
R47ZwY9iqSmfTqBwcNTa2cNZ+IbjYXBhd4gfBrNSVVuC0B07i9Up+rOUpANr
tS2OuMtjZQnqepWbY18oQWAwLQGBlHorp9p3RMJozlQm9ecKvqCWAcLUEg6O
ycE4zaJpgeijHFLMITGgSdVLrAHgtkIlK0bn6vYKdtBJ7zr0Myy4jO+6WAt1
FJsU/JNnmF6pOSu/VQ0gPtKoOhvc95NXqENa4c3SHahTkEZ6uR5jMoJw47xA
UveeL+Ec79+zF7HS0LXRp4cAb/9W/S69CpQJtT77pewRfpmj31IxgKEx/XTU
13sVe2rBrvyIC6xbwReVnmYjhwQxF00BqAhHMWiSOwGaXo3a1PUdLRkK4Khg
fQBkocLpjzCEkhjHaFkeRpUMY3bGACjJvvpqNiylplNccym008Sl02hCCZlO
L1FsIDa9RLpZQd/qjQjT0/DlD3HTRtgL/0yygdfy1H+UK/qEm78jzcJp5wvO
YAKRVd9/cLw+bfOVwnBbalvAebvZ7ciMg9iRCI+rX2coq54BeGon+rViz7cU
ujpomEIEkiQzUCea3KhZ4/celzrbqtCCv/Fo8WXrgCzUCu+Gib59kfZntA1H
a8zPAsINlNcTyRSvCffYuxUZEYCa5OdPxn8xz1/iGUXWAAyJ/KgKEK1kBaxt
WBJX+X5pa9+fxOThG7tXXTt0JqXXi3pOBZz/Ucvfu4ym8KFUzzgs3dtJxSkB
t5UrS14V1ZQguPacpdx55m6Nllh+0JNJtNd2IT3tIWD87lsCyH6HFifcwj2o
wWRoZuzhxWSck+JttjSWFhVpXndU1VmjDamiRcUXWk/aulxGY69846PgDHF/
03prVH2tHNk3oiassv/edVgF3YehOW85w87qEeDhuwxhKxuFY6pwB75/VL50
Os6bIFUTUTYUwT/mFlfad1U5TrvL5o8nIOZ2yU7CnuNpdrH/mgbM5mGuHSEo
QQbaoNER5xwoZ5zgAD5VVjgiulO2njO9BVUnN8JX1Z9iQEJjgMZSS/1R5Mbc
3g7rUIIKu5Mz/n6v88Ey08BWsLz9emkhejG6QBdNPBekffkNH06+1kJJmeYw
gj48oECJZvWt3MRUZWnUISqAUu5qVl/v1RswRc2apeg6aYt4LP8AEYsEy98/
gQYFVUwTI8YLYGJNeh4n8rQBQTloKaYcD1d6opqxNLZ6vSQsK1kLpqs7znjF
nDU1JuxpGoPmRxdyi1dlpF3h1fVt4r3NtB/uQfKI5dGMbdXxPR09AT404iAG
QoPQ5ETsrGX70vdAbYxjsYbafBQ0Ne0ARjIB7qEA+B3fHcS+n+u52/5jSq6o
RkUu4/yP5gGYGVmR6Zbnp+M8xuRUV8UFNN427x0FBdy9mBXOR7bVB/HJ4CoP
ahsnM2i3cd8oBl3RLjyM9K9NJ8Um4MB1IxK/B+P9v3bWvpDIBX0smQmxux1p
e89DkHiNay1Xnk7setJLGIRBhmFm+oM/2976b1swLMiVSPnYzbTuI73SX4u+
0hHMd+DhQiAx4U2fMZxJ11TvaCHlPi+w79PRtq7N/9xuk1qUkzejGc2u6yBV
iwvtMft1ukS97GOwd/nNiesLsYtVR/v/s3qCj4OAZ/oTClEHdfh+zpNZZJ6m
sGfq5fERcZT73NqD1FkEEXE/tYdjFG0IVF+Fp6PRxcnqFRTAmiSuX/jklFFj
ekA5BsGxwC85B1sy19LSxMgmEIbCYOz+VJL8g9BZqEjJPn7c0Y1NPmMV8o/T
qfaUHoRwLOFQ1xAtOCb53wFiZLUpkm+xwpDuT4a16CUHV406qspuMebMEoad
5xRgISNDQuvSocTGDNS0i+4346cl8Pv9wkcERzzLQVundazBshe/OqkKv/xl
+ZrLV5QXdjOqkhV1d7a9wizJgB4NX0SrSEuBv86+b9GegXFh2zP1ifFiIaeB
GMZ+3oN4bl0UhzlXGrTxvaMSYmHE+cxvfiN5iarFetc9NYDBp5rEiEYsLuZe
BHxQAuwnexkqQDtNEm/UoHMj8A/+GJndQxFvuiR80xqq1kWsRFWEUgfWGoEc
lcOGk0Z1WgfmA83os/+3D20fM540fccI1QRxiuHADsPjIZ1O3iv4kTVH1oi3
CpNdbZGLW6w6nHmui1py1JhEgEYHJ9kMdIhqe9P9yuQdvu0ktin1iiBdK5sA
/g3LORYo4Hkra1eUS5XmV345FJqJMXo7QT74lrdWoABbGrkbbCw2Sm3ulj1O
lN4eonBsGqlJ8Honf+262SH7VCrCwOJQmZXjb15lVQP8yNu+qq8ZgzfP7id4
AqwF4joJnjB2O4AtvzAN0W5+aAmR48UVBOORUpzKF5NvxlxNkWTzYewrjIpH
fu44OauijqX4D9Z/9dfUaqh7JqT5/Bzr74hWm6T/4nskH7UG0td8I8bsIycE
1d84gUsnYoTk9uaN8tr2VfG6KU+G0ip6ksapKVjDxwS60zUQgjjaMVo/GP1F
Z4ivBFpe8oAs0prZyaVDB0SoEVbr6jCUXRP+d0Krr0nzY+xqyGLXpr9Qxje0
bGGl09DymyRehw4nO2bWRgo9M+v7XWtSaMf1DfqZmlDrEUQPaSYH/W1dKGXL
FEweTkS4vi90t7611sRFXiVB0HpYzR3zJLAUKerSxg22sLz9IaPn92gF50/R
L4jyHmRuAGRG9G1emPjeGjtcnDPX0trdAf/p6ljwEWrVGaE3uqmt3Gc2xFR0
qpyKHCAQHP5lRykY3W+u9s0cRplHNgvZzEgDBzVOihTFIL5JWnV0e6Upif7u
Ms/mnq03fnhkwgceE+UggCdC8OeiXRp8q3CYengPRgpZTrTs8X2PABBmoe7x
0RGGy/ZD0FiBVd9vCpVzRoz4ktHdAe3hV9WpfT88I7A9Dth4mRdJkWzqv82a
YFLRNbqngmeoo9b0j6KzrxzvuGGT01IC6Pm+5pazo/tsJ1rNuMSDcmROuf2g
0/r65vuWFWyhCpptSgHRW8WFwfBxVp2/deU/7/kWoYmHBfsFaTiHDaDSeIa+
9aB0AjsLW85yg1emHx+Rn+TT4zie1gTPxHkaRQg38XTtFAjTPy62bME6fFFF
AojueQo6PNXfvSovywSoVa93HRS0fTrY5Uhj07QOvTwWsqdeDQnUaeVntnff
03nimeBIn+PWhvZ5DeRF+E4oAs+6+pEij6CvSNaSd+7Smi+Vy6LtNEyS+TEr
PUMbdEiO0Y/zIyb/7AtPZalJIwjTjdtUR8O3beO+HGmlFteWbdlqn822ZIyI
mJBqVJfNcGpCDXoU3IxFs0adinD6NHPUVLxVmJvfiiGY6Bo9kXv/3yb+QrS7
UI/UhLvzxw27rfGRboxd5C2uz/Hl8uv7h5IC/CHRLbCqc/i7VmBkvJF36Qt0
ctYnEXUrQUGa4xnty0FRCMFfevCwzRK/wGrBbHUXPfGs3XHx4N1FFzCBV6CA
I2LqrbpNSgqCSYKSpKhZkt9XMadiATe6DRWXh27gIdGXCBZwbMBd1D2pk2cj
cFPLvIchFqIi+7GLjjEYG99NJMnJpEf+JFpM3ugpeHYIiLPdE/dS6Dqhc/Vr
nNtB4/c21DY8qkrjTRDYeskjcnHw7a7eAMnD6bN+7QrqVcD1JVd62oB7o1ly
ACWz8uiy6ne+g0L91cO6Xzzv7mVAqDV0qo6KQJ4J8PgrEp5hx6VWKfmyYEy7
23RGiiCpIzYFbk6r23e614cgfv9mYLZZgCDh8U1vWJ6P90w91y6pJsh2zna+
ab658Xy4VfOGJJicdU8NLZhMbl73hOcFIvaDce0FWNvwbadrl+Beqf742zCk
V0OVh9QycgLif0KusKTTDI6SJhwuK1RPqNy/TWGTKyZM6rbvomEEWjQ+bpBE
1JunEE6LVX35CyLLAduo9plHwl9YdofWIIDomNW7VN5UXtAoyegMXEiHammZ
D4cFA5Dzq8iKczGP4sB9mF+uWZQHdX7Aqv+yhZ0AWeEb8ITIrpJ+8Prh9G6a
1dD9JU2PXGlGtg8dKNKvnEeNo6bS5rlm85NEsfVpNkFZI3dWJP/CGUgV63tj
RcLKe2BigVNZuw2pOTeqk0SRpHa9v/rH71Nem3S+UzluDlpa4RxHRiCCyi4e
FZAxb8eBy6Z5UhYpRUWpTnPm9yFXrOcpkX0y1/Guenx+KCZRFRE/HFyP1gAQ
qY+n9t6PantbGGt7VLGz9DCVJejFdrmLrbKN2AiJiKAf+4YRHNGbTfoxKQ9t
GENeBX+wB4NlA8PFKlGqzVZpaleG3f88+XhyrPkXaj/8Pc+20KkIxrviJQan
JP2vZKeX9K0Pct2dhSU2MaYJRCBKjxgsiFP18uv7T4TM5VC/3PC2gZ6nyQVE
/y1hEYyOxS9zn6/lHjK5X81jbTChx/yzTr3RFii+1h4cQPmTc6QuMdKvfwZM
7J3dA1l4AS+Ik3KuHrAv21qg03CCXAW1T734gUYbPtSehwAI25uW5DYAdb2H
UligGO8IcmOybVlf4agy9+y6eolIEY2OjtcTqRk3TlskLPegoU/xOxzmQf98
rcNgSkp7OM2IPOmw1yepI6spxtTAMm3LbxJObVxFi976dVf/IzBpSSdHCbmc
xTN97OUitAkGPpcRRMcEQT4vRsxXtLk7AmxBGOyxqiuuCsNHCw+u6MAIwsdK
eS0/4g99xZNYVXgFkqAFdsUqjxqSRvs6EhakOti+USmMmnG7dswoGETR70kh
0H94ED8Kopc1MwYh5SWs8JPy0iTvBQlIuDQGzkUP95o2LXp/UhZeeHdoSi+n
2YhuDXDBVyZ1dnccLfIAcDeLZ6QQmTbZN25FRs/hujUWbdYf6/B9iDsPq5hX
+BWjabYjd6hJT8nng8xQahX3gjsLth49GYq6n/BuUt9SlKr24lbir/bl8asF
p8/Fm2d3JoUniDukfhb2v8n5CBpP0GZqB/F2brbGMcAURiGuAvKzo7KulGkH
QVTosf8fjJ0sp/dGIhRKpFRIhobbaxydEpJ0P6M0LdMh73NQK0XE8E0z6yJI
mJR87FGBX1r7Ek87248Vg4HRX3WVe+hVKhh6AbKZsRhISlhHfWYSAF7gIfnW
Nb3umXndzkeRCjHdzYVB6BdGZbBktwoNwEaLJlIFzK0R7EMmv+ppRJl2LG5h
rd4SMzPYhNo6VVa/ByrwBNdbKRzazNinpPiZ43/v8O+htLRHHRYCI+F0X3AX
mU2w2b53z0Sh6Gy0McVKuDX3d7jQKQBtJVgjtZ43UOmkJdS1KYmCCmyPxMlm
EdL01cd2iqEaBC1moH5GtW21yXBdIfGNcZ//avKQRKjztBo3JLUJsP5Etmpl
ruBsbKHFl2yW9lqwT8cSh022E12v80usjbVpABtEYwAeXSx5+KX5TG84XwjC
oFtNPdXd79g685QCHAylDcYMF9o/u6tJvNzb9SK6Ic8auU3PupcOIFEtFFkt
C4YMxpYKQGYqpG6rC3dkmUyS++tNN0khUdDgMwGqdoSiN63Hg4g4AYNAT/mi
jvf7HZ/0Rdp27cHvEol5lSw0jxct1z2bZCii9SRl9OXgiWSOj/XYaTtME9vq
8b1D6/PN4Pw1X3LrOlvZAKDtXijzVeNLVO5ZdmPfs3PrM3I2OTxddacXJRba
g7qb6IHaOJcYuxyHhoWSK/WFx7oAz9cAKVUA2rgS5UFKw3KAAckiLJTZQboJ
8Ph4kst9IV67WJoHTaADqRPZ6Jrl/gTNatHOnA4prWBZPXy+QJkPQF2qIrdc
RhmfI6ItH5Nelo2he6P50aLGXObCHDnRSeLZ4/WLsl0rCRWEpfsR5tCq73oT
if7305E1f0fgweMYsiUvXWyr62AbKaPBU8fJrtnWrAiT8a2O5YUm/D4K0bMH
+crwsjUmSfYa4qvBz/MCFR4smczz4qec89GQFHGzwx9W3QkfZwr7GUFHndPy
vD+9tJQ+8w0zd2HzgMnXxFo5n4a4MOpxdqDwdxzpY+2TfeRwo7cbAjugNuFz
gxspv+fwvUFWJwjgywZT/iqPS2mfQGmcSQJ2u60AeMylYfu12Wn+/ga+LhNG
nFHbEXS/a8H1k7YfulBJM1gVfZqCRuDFJIK9p1f2lwTRZHs8a52OPuMfm3WJ
SXL6LQKF6XlFKpZUGknMuPyGuCiw/Le9zexrN4v9ohSObme5Dgnr4K/quXBj
GFHIFpE+Xpvdo+qcHNCkq/vncTNIuTgvCWoVYEIF2spSPlD7G/AhhQeePqxy
HFcc8Ahh1Nqvlfqtfr+CODQ9jTRYa5sac5H2mnDQjuNILCLrkyRqEr78UNBb
WpNNvkgRxDMMH10RAjA0FJNfOQHRgJZ8Lq4wJ/a9mWdhBTqkAQDcL8OsFM0R
YDfXTAZIwwhyAAazS0KG2CjDHGsbC1IoqVjhlEPzv4OnWoFZ/J2VevYJcNBT
5AMZTe0Ud3O1YAfxsliL2M8ncnrxE0mbUHbplCwHaEj2mvpmPMdXsYzb38nc
HUhDPH5Z0O86LksI7YZrGEg+kWQZDIcLSTHitU1LLP0QUQP6zOlSepry4ZXG
DRwnbTwKwQg+rplReiEDSsrkHEwYrBCKwmBsxILNlDGsbqmxeSE67DebJs2Y
UTrC7kjaBfg+kUjX6qmIH/VayOLJLnfjUBnbcPmX+uw20nGSGlsc4dR+zhkx
0t9vkB3SmD7YuAqvm73pvaOg73zmPsRVHlfkPCkNkLR94J+hsEvRs5TFesE/
4ffAQFLcQhjViXSFkJFLEJxp1NGck5LWsY7n14zLoOh8iJSD+yxtLNfZrmhh
bGQ3QQ1BEqkkIHvrv3c6sLBjGOll5HMm1hKOHLpdDaYYNusE9W1EvQfmEBvM
jcTplN99qlfDMMcRhQ/fXee7DTmTLgIG5CqfX0gcl94m6Yk7hAt6d9KHo9d3
4IPOtOK4xHJ1osG0Iw9NvWFDBpsdZaMTB8aCKikRBCVU9UdXRFtFK4jp/wON
K18fJq8e9Q7eXGvsVVLNIqGWTaA9r8CDYiG2dJn6Kr9RwM9UgwKEXU8Etu0E
icfYplfqQf7MOQQAPp29m9w+eJh2NfejhXwYJKr6n6plcLG22FfxFJiKragD
bn/D42R4EeolCWzxBDjdiYBEg5UVzqcE+H5h9k/wA33I2nNDtZzTMz0tI4UL
ayEIXr4t0xZ/R1E5EuqUKQCWap11pv5QbFLcT0qnYXCCoO46ISVdidjLjXVB
mCc1dXeHxnlwirYHoghZ/+Wix0pTrQwb48xImKA7A/i6bkuW/cuTIt0X3udv
OpNhNRHMZghExJcRVunX+Uqp0FRjDxaQaGVu5gg4OQ6UIA+3QB3ehGZMGWmC
EKhFg6bU8Acucmo0NjnPiamlGGrfbIBCY25hxR1dEFRwbemFAX2PDivo0y+L
aDsW/na5Wf4aw/dnwL6z1kRoQnYUEqcXDhZlIJb3Hw6fveJqYZffGRHI7RUF
wucsJ/JlWn2jwBCk6Hhv5emm2hi1+WvefLuXZb2STZrb/QV3y4qBM9Rpbb3c
WyU/bzA0q2VS8Vdno3KtY4+HCAWLPQxRweGBWsttf44X0qw97Jst0Ctw9WJH
au7XbuV5PNG8Ful6x9DaEDh6J5DYkWQPyuCt8hHQzMI25XmMJ4uJryzQtbZe
c8XoAdrCAT5NB1jglWVoR/ENq0zqybr6EHURFeDWKkHt/8+g3K09SdrshPLJ
Ct5YHvzA/r4W6erS7EXGxsFMmt1FeCLyB/k/VvvH5WflpXsClbiNic5RbJQ9
H5mCEXho+2qurjtC9yrFhI8qY4izymDSCSCh40KOHoTvqKo0bpSquG+ppJ/j
SWBOqGgqv78GgZiBEHYgJfqymW1+kIVF9qi5Af4SF0wKRX6B/2rN4ps0dQyp
A4H5W9Pwa+HssvijVajMbW2JT4VGZMheKQDuYzJjV9lS4m9AQ51nf2qgYWOQ
TL5++4+OnmkOZfe4jHFlhCev9PZeHOQzHD18oYrJ4XmowQWqhkAYnDHG+5eM
/2VJfCg6ZDIGMXi2MAGnQWoObEzhShm5k2Eo/+ksmrmY0qi4GCIH5sHNs5L1
obIz2YeUCH+T8c71ZvAbvg4zLNYU5SZ3QW6uRyFWR8KeuIDyDIcwJ/0i0a7e
hqSuA1vVyE1nA/PKsjgt6js8ftLp7j50S8PTPSs3E0h+uEWEI8Nzo8BlSXJ4
p7556327IkwW1sFafTtZYwzk81KsHl2e3U/dBJiffXwT4fnDuLyViwYfIGy6
HxxQBOJaJ/AbH1kcKMnOs24FDu4IDGCoJ7vlWERt0ZB3aTuvvP8yFtlqYPOf
ZOp3UYlAvscuyizs5CS9XRO6HDlDp2nOMsjRetcn9DDS6hZFsFu4kCDAMtiE
tezYNGDit8rcrfqgeePdlF90TmwB8uZA43aTnJDNscdTtHp8gEm2GBgCEvrH
x82Je4CeVUFib8pBWR731VujUOB3ig22NJK6PtwK0kJ/4+q1LS/eg3fbYBSD
n9Woqxx2A4bYXYBSFhmvHQCPIYqHbBM7CGXB0EMBPE3ElVqaXRb7orB89S5f
A+P/SUnUfWTJ5b1oOIWMGWrxTYtpGo2BP8k7O1RuEQY37dT3BkIe+F2838f0
BogB2m7LEMAMCPu1sdTt+LNJJa3XL5sXTSjnjLr8PpnSjPU0FcDsxHq4pHLy
heceOcANC+ge8+k7x4vSMadlcDBLojlklrS9AL0gf1VnvjbLEm0ELLkJ/8xk
z3eMXnGWpN8eezhTpzoWct8996qC5BQkIZ2KPEMGHhDttiDVJLyZHlMVDkMX
A/CFKWJELBa+2oRoAxjyyj+RJch5g+bWO7QX2NPi34BRJBM3YmA8PsWCGIpm
WcWMtQ1USs14MjCxys1mcnZXrcoriyuZym+wx4/gGM38Yk0LOKdEWSN4/IbG
rAPITK2C8DL909qbWUBzJoHQljvaDh+meO+QUwfFBLu0cjAcCPDJ1luLGZfy
hihwRE3pLqXdjx4ic7q+1pgj3XKrC3dQ/8zyssey5aU2yPfNaO7wukGTF7ud
iJS31jurMV7ot6S0gSTe1OyAxtmETzx7j1P3r3vetCei9lxQbHvKhzAOc9AB
kbNJA1GFPVzzsLodzZlvEFZnxl5YnJfjFAYbDh99TrMZFRnV/LNXGsa0tCVC
2i9QgxlEg/vVyAx/D3uC55pH7YeXXKLNIflCfI5Ju095GMkP20giX3cGA2yD
i8CFeRlVDQOtegW7qjT8A1iqIF97H5JPrLg6mJz6+CtdAepLQVpPsb5+/W7R
X7Q4qVYM+MANtZLP/SMe8CUMNqqmAe2u7+Ur2CCg5xUULKwDyJvSm54139xT
N1ERziapSztBQ3C2eUcipUKcNqqX571gOz3pYXfw2S3jTwRWnOFRr24HhZ45
ZeTVMETcnS8lUg90oIk6zaCUK+ikOSzjvHjPekNhDWtQY7RmGxx1wKNA8PFm
3ZEl82uKHh0qZjf/TEq9aGOTpCj89jHPAJ2knIcWiwkuH6j+tVOS5drYRXjg
mQ54rKOlji1uIVBQfndctLqR18nA6loItU/cbrSPKrsmWP/8Qh5dd7k3OXVh
KjCGDlt3Rfd2ZX5oUphjVJ8glkqjiznKjU+qt7DVC37tODzrh3J0uRrX8WAy
qJjDmkIDQrLmnezlDD0EYrxf3xAYfHd1ODs2QlLQDDOCtYOqlPze5hcAhzXr
AYiTVX9JBcA8nZv+Hl8gPoa9BDLbQ+JXAA48L8idbnfG6F8PyJLtBZeCihlx
6P3eDcqBjnefXwaCRaDz7gWeFmzuqPFh3yLbfSI2gZ974uDmnRrYiiZ2SwGE
jbn86F1TsAULsyRA2nIPkR4VDmTfGG0C8JGBJaqP/Kxh1D/wjNxS+mI0Pt37
RG1tHyY+ggblaNZN8ILGkMMrWjqq488pD20JwqrhsKZyxcJ+QA5phSrdYiyS
xpMJTgprPriPweaF36QRQ/+HdvN06NzEztEVHJf8MoiM7C3j5K/6xSUpl4ix
7Hl5UyWUx/uwFcbRjpMu5LTSWQL5rtDtz6q+lIxS4HqKNFgliBSiy43OWQmT
hGTAa+aM5MRlYiNcAb4KemeOs/GNW4otRbEPqQt3v/hFaI/XwCsbaHSTWLQR
Bdk4rkg8oty+k6fTZyG+GikHyjhFQmIVZYuV4iETC6a6PCdS4BntGGB/Hi22
JAhs6IemqhTq5O1SF3ixRcDIPuxzpnIJlZZxai7iu2lP764pGZzkHKt5IkFS
nDRY9PGZZccfF/trDUxSP94/IN/us7xD4gLZ0FtY3iaGmu6OMB20xGwLuLKV
CcJqUoO8oBlTV7kIpqgHQ1zDN9X3Gg9Wn4T8t4mZM3iEqFelIjNzCXm/zz+o
yFo9fVEEUgzO4rc6ItTouOJYWDs2Q6aP50MnrWt29J+h2452tt67WVoaH+N1
lGWuGd/ZltZzh/yIQssajoEQxkbABnLFPEekJYqQkH3UUd5ZcBMRUvMyarDw
gEWQy1R4Gyj0pHMSbFO8bsHwBCvTUgwRxZZbYBfSv3yNXdV3BQ6OwolOFXMP
av1+g/VU7rEdwG3COebj1lVcjYoIT9D4sGc2XtPRbQacNk+aKkZTcHywhKm5
RFnat7ZILDeqr1qiQ8EBXgURJVulaUstUBLR93E5aPzqneOKTlqX+Nzht1qi
ThXXBbUnLz9WijetgXkVgjqyjfXpCdb+m8ovVeZfxxrCwO+as5lN9g54sTCZ
GysGw1kAH2GPnbGaeuR7DwvHcn/Xgt+y6n1SpikAhLY/ubX3/HjmAfihL42o
QEwcD6Pnn7fCZQyaVcXPaU4niAbS5PvAp5iUuYrQWiOPzr+q6auOxRO6HoNC
ElKMm0GhZRp5Z3dHzTZ5EzdSZ8l1fG5IMOVFDAR+v1NIjG9T9gjClEaJfyHo
AbY5EN56Lz/tm8o0CMp/YLuXNplpuEJG7cwqfr7P1MWkoB+rSZ0TJswJ9798
7R6KG9tD9NS1tl4uetc7dUPSa6Xbs9cN+EgpRa0FeFizU5hPm1RhZ7bhCS+f
6o1X0Nq2j0+ADq+cma74J0xuj4AsAFB0eBFk5guiMnCKc3t686kPCFl6v0ez
QMRpV5ZV5jlSGnM2ua71YBP5vBDH8F+kGFxLaTzqDRyxBc3QenJddtiOzeUz
JgXtOT6SMgC+0b0TJpWTnnJ7oIg+vqOkAwIC8dmhAq7SHKgXn8e7w9lmct9m
t7QKEO1UzwwLw+UjuuYZG73iuA4qKncX+tdmyZ+ufGPHY9In3pNKQhLame55
ItwNhpal4ZH7CMZj1trgDr18xnPUqrinqqeVsQK0hBcJLsVUIzDXtFtSyR4w
4U+BpkavsdKn+NZ3ZewTRtnspU6b5igMsCe/xwW5X45vwuMSBFf1J8qRM/V2
wAnNKIcJ945AkJOc1noEMV54dWoaWeCTdsdIjsed3U9KauRSDr8KT37B6Yin
y2EvuSAFWrjVxlfFzQ7cQWcuUv6GcURerZm4b0jyB4PKxg5aYchPPaz1E7U4
1+/cHIC8vbU8qPosmiEj5DsqQJrn9piMA7R6j/Ofk4SItvP8tytUNNW/Xp6r
kC3ErB2GYJYRApxXC63iFQhKCoJWdPLB11wPVwxpnp+JAkke5IRTcnyxexdX
pnrZqdxC8aadoIY8Wh/1JJGSYa5h4ZIsjdhJN2uLrBn+Zpik0Ix9SpAT6e9b
CPZozzmkb60aL2gby9uVoan4wBGQumswNm54Jzpup/ZRo/6+G1WyRRzC2Huv
YP/aUuNxa1OLO9JUwVXz4kUZywMZhh/jA49Xt6pfwba+EUGnD6YVQc2TlYAH
Mgu7M4b7YUU/na8DYHDlHAmBWZzRXYQF7dHt0EKSRW1gl2q+wnPvsAPjsf7H
3JGb4iiIo6UcBohVhhRSTqpcLeIycZYBJy2mtRBWt79vW0986Sfe3mh6mBZE
gARD4TgUOl0TcOI8PKnj2oix+GDwGVdyi98O71MZOPzXqlbRwlrbAm5FKqM3
8ogxrMKR0rcoY4ZBTiVnFRDcJY2nXoc1SFnZzyI9LxkSM8hiKK/AkE4lfR87
lbPnQhLYqC3WbykHU9OgmKEUvKdciEtsskDFg75te1iquWuR3kKql/NHULXc
D38twEqRE1KBhMvfW3GBYRc+OCJ2EwWufRYI6KpzvCsqpwmV/DbefwmQJXNJ
xLn/QJubgZbsR/7b3eK78GcELz6EZHb9Id/KOmcHBK3FYjzcfEzaXYaG2YU+
W4FoxlkGHDNca1QA1t8ZCZwojG5S9NEvMXc/skknB1I4tYu8fi8QpMI9hmai
dV5CTdakoYoN8dbZoNTtVO9TCaQf6bucjJOLLM0P4ypdauLgZp+u4/Om9so0
pQLpHUbAo6vHVI9kK/2BnvMbdQg7gB4BKgVbBNABK/X2ZF2g66jRFC/GtfP2
A7baL2R054ampw7snzj3F8PIxVYCWjIL9MERC24ga6N2zvfTBruJLSvr6SC+
zQ0XdfK2TdOhm8FleQHEe4b2Qlobda/tNlLPozjEPfLnFk7HN/LGQdvlbWYA
ybSRRvwEPsVdGK7vj3z+oxDgWTT8LfINIT79CaryO9d5Blh/WmFsZxNNReMT
RKkkWRr31zO4vuHQuc6pi3/0VdHu8uVHNZQDl5ESCRR4HOS067+Si7aDWCtM
ZPOP02VsUOMKS388YOkT2lIuhsVz8lDE9mmyn6M1LKUB+OpaqoH2TKGvoqf4
ysjgBudQnN+iEXYNLM12+U1NKAMjg53zQUCEHhTj1JyyErJEhIKt/khW8MNT
s5UbFFG33f6YXPoX/0dPVy5bXXPko26N41pRZ3C/zbKxZD6YGIYuo3BSRgLe
9ytu3bngIERhjxuxHnGSKzb8xKrRUeMmvj3G2O7yRz8IiBNGerE9bMgkE0fr
EPAZ9qz+TkTqjx7UqekPD75iSNr9mDosQMlrezimghWgc8fWecoHjiY7Ie2T
E4uAE+2B/5LIJ9Ahl46EZeD2SnkVpFxk3Ys+afyxGU25LoAaEX74bW9XR9fO
nd3EKiig9UdH/y2zbTd+ljxC0HT6XEaXIJDR0D3hU3y0UD5FqqTGORi0TFfE
6ylQzqX6BYbgBBpO6zHpueOhum9GHnQ4AFCp69H9WMcWCBJw0xwCy4w+chp/
5FT7Nvp/2P44ZVN6SdnB1CPy70bt5+Sjrzx4uo0d4pynvVbdxtHBRQwYChN6
//Jia4bvsJHgj9SUPblgHqgj/XK+69YiXMJSudXr3/CYtslWT6OZe/vBuVtI
PDhhoJCP7Shm/bmrqYxU3ptiCIlWwj4FHEFEZKgjlauU4vdSA/9Bab6fItfa
LPkLZ0sAjFF7zBeUDV7LYcd/7TeDSu0hJenCPHpjfVXBwWg568qxx3zA9G+8
RjUWMnhFdqZX+iRZrdTKFiiT5L7M8C21ZyNZkPNnw9seqiPN1m6WBI5pCVdx
UY7rULwruhEFp+owG6Wc14aZfuxYVHMpt9/tPOAvL9m/AVJQQd3g0PVtYX8y
PZ6Sa+AsymoCxIiKNbjLpHXDC8r4wEHKuEdImpIpVjKn3f0Nj1dqhCP7lHJn
pdxci3W7jO17rqCuy7XgP+3QuGU8+rRSJFGGmYeYKTSSKH7vUHF7LSMYQ5gu
AJux34x+SGUGyYCC6Z+xiEQp9w2dv/olYzfb9YM8T1CxjOAI6XzedBaHHA0Z
YglaAYoeYs8M6M70t31CyBIEgvE+uuNmCSSYfeqC3fGt7MgBIr6JxoCO6T7p
FCDZq9b79VNg0i7SD4y78bmrc4dYSe7ph5roT/g3J4gpkKB/hStZ7M+xPstt
jpC77+oWII6v4yyt5AsbUKCaYqv1CKH+H8pFPQ+lFGxd153hTHCJiwmSPIq5
e9KSE70dMjt53+AuXrDr6uWo/5a1liTD7BxNTbnsxMAp5//r2wJuOs4O4Z+G
MYvGeuZn7GXE+pTDYX6zvTPvdP+Eed1TrDXRFHLQy6ecpbtxb1VWb6+uYErc
ruh1xD0B7w9+BR5xLqgTPa0iEh0ASAzFKg1KRyUahHjoSryoNBwSyJdg9fuT
vCTOtonSRBxHSHJeezPnUTbL1z0K42RBIiXf2P61Mqo8NFfAWLJdNRCCtVoe
W/2XgqnsFeUHcvyu9hPU/80gmah940y584D4RlGKvtQyRGPnyxkwtC6PHStO
IsCPvgdIp90UWBt00uI3JFbGX2AVs7N7Xx5dlfPlzkkdosl95suFwCi/8LlG
+y08fJHVz9xhvcRYwbrihYZZJm03k66gEq3BJcYQtmWAbPYaLy9clvA+WES2
VnUvx98o0LvqEQbj8K4KESO+3Vex35T+v4X53KTYHHTTGlXuyPiYaBE1vbIZ
s3RfutETAUk76BRJ3x1EPa5qAkTkneZYUDjrvt1pGrMoGKGnNUPtRk+OEKaP
1A87/ajkrOo5uys1lLiHT64lO87kjX43s2T9yin7BT50dUQ9xvwpVAyv4Yjl
MoJGWUjnWwmWkpDEiewKZkKK8AN7RhGPwsqzF+fgmKlPrHqrO6V991opXtQ+
e2z+nwC/cstdq9JVXNuEr0Oew3FvgIcjsx1LR4JY3mGNT/CM6vzVx9YmxVtW
TvW7lVYTpGFr2AuythhhCkY4+bMbVjEppx1wym8H7hcVSk77+mgku2wpu0uh
wFbM//uy+ce3uMPHPolmG30V3FpDJbuVU4I44KJzYlfLsXMC77CRrPJ+AXqT
JnxIMrmZ+dSELDhsxCfgUL+v/eW4tSzqeRbXzKYVVDLJQDbNsysKLlGjfiZh
R/j+w/6Bp1/e8JkgkFFu0gfWe/8wY0/p0zfuDl9beRzyg3XroMa6aTfajWrB
dYBIMdQwk79dh4p39oi4Pf4cBjtERjNz0IAvYDnG1Q4r2APBMS9SQAgGj1Pk
IMMNqRas7xkzwwEWhP+A9LwSlBGrorDDOWgqXFX6OG1PmR1EsG/LaCUI2kUR
bUkr/uLf/lmL6rxx19B50sFEB+p92oq+YdKhOQtQe7GlV+kyrPzWvJf12+wO
Y4viiVC5KcM99mGqQbdAiniPicolQ8Y2n6eSm+vz2GakSrhhRRlpPHdmUA4v
obChlDyRzeM2ErwHK6A5QiAelQy85z5VtseXdmZu06vInFEqwn43/t98GkXU
ejdfGtyBTCiyUZ4rZDXXbUB/KB/Ai8NVyOZbTGik0/uSC2xYeilyVmWPmLAD
DTZUBNJoUm19vI8dswmRd87ptNG20qQUDhVe3OUmuTBIGGN0gRkHGDcFkcPY
NyDJfdhKMuLsXFmiZHCIBv91DCp0wJahu4Inqor0qxk+m/TtfzulghyA7k3l
hs1dpRylELpDIJQRujNIvAkyi2Awv0p1zpgR3ybynU6dHQ3myFrY8J5v7dJb
mjKVdeMpBXqjELbqfqqjBZezviJrYSPMS1v2xv7qXL2EKuVqcoDpb1VQO7wY
fqeJ44TuhfBjiXd48bWLvUKsWoz7CS6npJM0FO4qsLeZp8CRijceyphFixJl
fHdO+9DQ5XXQ86/3ASZDXjPKku3R134WqkIIJAzzLIV3Q/aGSDH5TCYrId5B
OyAfGWPT0mRajHMdZ39oWDzIpYfaXpxVr+Pc/2jrb5ZB5iL2p7yNBu3ZvDlO
Q0EMB6S1zbeC9ByQHRFV2MrSIKyR36KO4knnUSaiaSPxJl7STuTDz00FSh2e
29UkL1CEKi2gQl+uqz3L7gdNTQ3ptRJRMt8Q9DHeK5fQvccjFOJAN1zSCttB
a0INs96rOShHSsPS6Qr6wBcxj7kZSHuKg3LWZtHKQtT7MPI7/VYC6atCa0sq
BjYiIHFGHNVYvEsdiUfthtp+3hdmOy1KtL3UVln54Nx4Hc/662GrFF4VCjqx
BtJbnCXiZi6ENcmdfQjME0oo88TNqzQ/SBZLm3bHkAgTRHKFnWjbUteOyuZM
M7TRiBXZun5ZZGyM1q6k2Xn4iY9nGBJymR6gs5xWXmQ7QKFr/Y6MTQk7C2U8
BTbsTX6OGQzO1CMpfXEg/Url4SwQBLnvwEOWr2mlxLVE84KnfWj6W+eKYhj6
71WP2kr/ZDU7puqWiys2f7UOltvfoHkqqa+3T1NDbe6IalvhCuWzjoIlsQBw
+KSkj6jaj09cxOEmrreK7Ypc1y15JbgQIOjoSxdGpT/+kRhMzWFuOydtMuDK
8//NqQnIkzQ48KX5wd5RSdpPrKrdhYzO3ujfviv7C5dxN3tH94LhD7d1Mozm
dD9Am3w2oWdZ5YAIQASmeTv4yxRoeE19Aofu/Tg4eWYBBnAmsHzUS/+Ocy1l
ucqmLsMH3dDjrkYJuxsKoijgpVkFXSLPJKewmVLb4tc/IOqL39RCfrg6VCv8
tiAQ69qxC4/BFOE/Zz2tyD5cxh3QfhfmGHajTjFqcMvljMWv+yt7+mgJQvko
zVIwKxbfVSyQbZXoJVu3jCGmFQBZgtn2IbRd5QT83Ww30R7YCsMIW5YDu4y3
+ThXTKtR+MN6iQRUFqwh2aHxa8rhPQdfGC3TaITdpaweLmIwdMejWQs3J1m3
9ZaTaOTQAsB62Ct74Gs/0I99xGiID43mbvAbu4GgE3k7SGfBrlKc2QVdgJ2P
s1ZcWaNHQzD8frhuG/JKvGaJsawtXgSEfKfx0NrDsbJJm4wdygtvWd82fDjN
TShFyXotApCLEr5ZMy/7niugy/4EnMvO0+1gAjUvVB4IvN8gBS3MAkMf2Pbk
/GcJwJwYaxX5tI2Uslb8mqfcUPnc/OJNuoM+zYLU+liV86RebX0XTC/mtx0q
FuTqeUR2UvC4auXbRWqMHye6zGK8E0+cFljZ1N5XGuDZ4lfg4E2Un2LYOJxs
38jm1XQuVMtUHRKgXkOh+FUYBewo69vSILvi8ppnqublS8Nu5cE8Xf1dEi2I
IQePBcXxJ145Zb02KsVmrQremDSq0GUC9kzPRYeXcjXpFzZWMYRmPVfwQUN3
60PzB7zTeR2Qa5vX0YO0NGbejaDedq0wuWfKkeR/2ZCnC1gh7ozbngoD5OQH
coEzwXHC2Pla5cwycDEL4V+WkgMV2kl6dIOueiTjaFlgBwF9nGXX+DAREt5o
RxIqZ06655zjSBA7Ci3brt7oJUtiqivIlRLfz8Gu9vehAkJbpDYrGbwIZf2F
dGoh1YLtsOX5IwV6MzQGxXGR9WCTsRtYbQtTHSZdQJ7YAQb57TTmXQozSfH2
y4genabVBtnyq7fc6kq2tFkqKHJcHS1FkCyhMQQxzhVTs7HRTEqwkJv+wwUv
gO9O3KITaGO1cnFrT9Qio7moUT2wQWQCe/yjbl9X8vxr/n0DnXJjnDNFZn15
8MLAhLTXqs84VndME3mYf87RsiisLqPubWOfXoOWsF+BOorsUh5eA6j47vMY
fQdwIXqSOTG+21l1BEzqdM0ts3UXCVZt9jz4tGadEyWGUo+IdrLsltImO94s
7iTb6Kl7XGVD184Zaq0SKadph1OK1Zh6Ors2pal+Ia1BfSyr0WLeeTg93up7
iz8MzQOnw4p0rj0hN9TgvDCB0grfO57MscLEjKiMgCRt4zZGiuEE8j/InZg8
XUuzr+P4QWDjKOXVblR0WJ0jhGDemg+mzEKhRGacgbLlagsl011cdnaYfVpm
urV7cjFQQbqBB/QWoLGELma+zJerAmeChnGOD+nB9mehJYib7X+tmFa85f2M
NDmYsAY5IS9iuGtVp73QVejnREiK/GF94J5toA70aYywgW4+PLuuq1ijKAvQ
pt0ojDHv8lAr7i7u7Y2e9MTdBJXzFLAJE/VAgB4l98CSq1sE30/+aTaq919W
laaBLSMffsILrUUKueuWY6PZmPLmAozoqR3YsJEkcwoiDxa8xssrczj2FNNz
POue7n+byKMUG6BoS5ar++D7hxx1AvPArWeHiPQun+SdbPvisSVifrCDoK0t
e942QjcHA5Bp0f71gqDiJ14HAsaq3wbjuOTaaVmAjvm1Wnc6MuKbGlDrwlJA
hTfvtOcih418tT/q/JnEioFcfMurQD+QQOalNMMupd7XEPSyr117cAzYsKHz
F1rbuRjX4JpTsIcCxYFa3jBgRkd/oHC1GJzExd5M6bTHqI3kG7lFYx0tuDRe
Eg7pMVI/Y2oLDPbrmeSE5BfOLI8zb/SPfOzqVUYanmZBbFJjiFzM0nICA5BB
HUUsPVtgq1wGPcy8KW77Uo2fvhqkMbBxg2t2DyNbj8Ohrqq9uq4xfbQCnPqC
pPwga+dPnf/iin0d6wJWm8AUWj4J/QHkDFq3OU0TP64AtyaOwW/4xVNsuwOi
KLUvHXk+ZKqXb1oRQR4WpV3n7nuY59fJdv77/fp/8x5i4gR7ioSZKUyyvwUK
lOapo1aW0uwY+682fiYYdG0Q1jDBE4JuiptUZ67RGbFySYfOGg6Yz5EfsRuy
lYQCZuvnMQksBSFoPCW8bNLFQ1kfHsGV3Sf2rZ7+EklSG4Lg7IoF4EeheQHP
EMMOAP6jYI6uS96xkxS1I+OqesQhEj6IqPXLLJM0VotJLYT+2fmQTfoXRbd/
80As8ZmLAuOGAP3I+PumxpmfOF6/l2NjCJ/NnEGD37DlUpjLlwdyF0aFdODw
n5He3iKuWxmJgc1BviJbJlL3CMVp7JQ7/eBNNaEWd5ALPjXdyslIZTP2pKNK
xAFqU70mCVI5YpCC1TVshKZg2H7zTQ8mxQTJBRJVLOhUhZYPPxik1O8wX2Yk
XqbVAzMOeCKfz9yQRrt84Ak0kURQAGCU7FMeuLms3loN4XFBS2ozAm+Q93+p
v2yGNRbr4WdEl7aen2chQfo4XhCT3wuDPFzsZmQE0ru99NJAMvn3WVnanXES
j9HowILoPNgNItW3Gtf+ETt3aCAEjMgsa6xxqdIC6j+b4i3R2zOr6MCqUBRp
N6OLvWT6mOCSWpoBU2wgsmRj5MpZLml+OIEAI0F2NvjLnxnWHzVCQu6+OpnO
nhwJ1kNtZ7Mi7LTl7agHmqDLkNXBZzyIXtoXCF/0sgXafcxDuBexnTEYC7/l
Z6IAiD0eX6EPwigh3i2JEETQzuzSCmio9ku9IGerZ6IhqiQdHyYRs9B8D8bo
5gMDjlbTaEueaePho0wnWwX/AMv4+Vp5ZjyHQ/XvFY7ii8Vn5u3jIaikbVWF
D58B+KTUanpA1/DQFGpIuqr2Qz1UqbZohhYNE7uzDSgXV0hqp9kcB1RSJluu
q3e6CAdFlCLIvGnJ49qCENV4jbyJ86plWAcCFmLGDYiOa3IbS9zWPZrK6VBJ
iBzG0PxI6wk+DB2r4AIAzfOu/fzSebLe2N3P/JGjmPy7zEwCV6erN1N9mqeb
KnmXGAVI3grCSvGeKzzMfEouy/iQM+1AyXrdvUvkwq2nqC0tQi/goCmOs3V4
oX5C+EpXjKVGjpSPCH8htW9fBKvdPzWLjjQ57tgbzqhk+k4yWbo4trH5Fr9e
vDTmgQHrJUkaXVGLdlv/K4Y9b2zzeByEHnxwixMjErM6D7VHyQOnRlYMWUlj
8cD3iWZ0MpfOCtDpEPX+6h79kAE8bHCEkaKbDz9QHhgZSbUVpfiGEABflpFO
JQbSaJxMOOgxR5yO+Sd2kGAEiyNZ/xc+6XJi7b33Kb5aCUJnKL46vmU2RXhH
ky4s9oE49nLwxCA1PvkEKjp+U991zuQiFjDGj3jZuAasQp2WTLFKg35Aywtm
qMebqv7u0lupQiogCkjS+8oy3OVmOiF6ZjtmgGxuHpKSY4JvSWqIPxsF6VDT
I4mUIWvaQiADhCa+DQzwnDFmmlVtIGLEbUb6j2IYtzymUiFCe0bjS+5AnEVV
bNWYvz4Lu4tPXJ2ZSpL8MRDQxf6KCv+Xbm7W0LdRO4lE7ENX//U3tOvmsz3S
ZWPg4tbXr8PsRv/CDl2+X9Mj/auW8XhCClkOhL1QlnX9fjqL42enh93Xjr6o
WFeTb1H5r9bFZwTMKxKLOCgzOEHIIfm1/ygnxE0BmWu4PJZIlfuTQMkfxi5v
nWKLatAwLWe0Snh8I1jw0emyI89Iouog7A8aqH4+HEZkbcVlqH9H3D21JzIH
Uyfbtdr5kcEV6rhSao8CUdLfsF9QHNg8pAuLwoYVldeies1MHhD0UFV2rH0j
/V5eCo12+rbzggqzEwV7jg+IPsI3ozUHAX4hBpWkIkFIK72sANn2L6fJNwK1
mhr9/SeAff/R42tcp4oNvLeYJNnemZckzgiRv1XbuyFbcFyItXZggrUUH3PH
K2f+KhMbDksygf/5XC5YiU3yX36woXPjF2KClIL/EUj0yWNOZOsh7R/Vgv+0
Yas58ERlPLiRMZ2nKO2+lvZNX7fJc1d8GPNTRZOYU4kwaegh0ypvP5BmDpKz
BrHxRsUZ6LO0Lremn+lhwXnclm9xS9RaBZh1H8ij2I4EfaHVWZuNufDMF35h
PI3ZgXijbeVL8s94Luf7vh5+zQFq86lFHs57IKCwgWMcgX4eDIVZDe0f+Arz
KhTvaGdSWHdT/xIov4DuQCLToIs9McvGg6soNvbtIpD3EkRw3iQNULU+3wrA
Lce26Aolz3U2JwcogRuWCYZXQMX2G4XvE+A1OHdZ8Yzw8WUiGK0Mw2gHkOPg
DGADesgtMlRi+TCrNbaEhkbIYWFVvnv5aqMjKVM2DOy0kEJCecZjj1dOGjiL
Ow6x9He2++IbELWzHTaEmTl5uw0VleWJmGEnirC8A/KrW7ChT05RO9y833WX
Ig4NhJsQ5xTFGhERuqrO9PO35oyBg5ITwnWlWbHFzJJAfw3k8aXIM+T7G28q
M+oCCNowH6yhMf2GokVrLBofECXrlDoxjcUpF1aRBnp9f+FzeQIvpuQxXkgd
vyQe6JPvq6xa2xdyzDJG4jqJXS0SLbYdR7cDKpS/9xAZPYw1yZxxXhtKXwcs
ltD01zZijmkie1azYFh5ClyetTr2Rh3y4IwZAkyG6mLQKM6gH/8I212MXy+7
IfqwUe7ph38IMJbLHeZzUBtVp/k9lOE4gvTAY4aGLn+RVURsD/eXOEGQ6gdu
3tjLaTX+/a1xN48wPz99UgaBN9VQJyIPYCoAHYqzOvA1vx2YdOhGNb9RSHMy
2wWCT8C1WNYAOB0dRpYFFCngRO5RHTv3AaXLBYb+GYBsb7kv2sh63wgnzayr
mZ5PIHbcQyOwMupSSwUQcMaDZhbubtChuCDTQWhIZpLPzpnTjCYpUuxlPejD
gBHwk5VZ4lIDAM9rW2PKViyKiCedLxLKkttuyu9D7qfgmZKecCxZAcm+2chu
i5L/v80LLo8jxn5bZ9vmYqWBzyf8xknJVN5oqWr077Dt1V+r3Q6URTa2YldD
FsUtOv7sejzC6UzGn9PWY6zxcY6kvmJUj9cteesF2IinxY56Klo44fqZc9s5
09o8OJXINOCkzzTx1/2LSatSy6ppjJ+jwRuQm2zRYRrFQp954LBLrePkYyXH
5aHr8ddDcVOsH9KkdghhK+7xYvpXYp1lfz3N/mCDmpZdOLmNYCqzaStHF0wR
8KLNhQyDDyV9w1FwuGmpoNe61z/zokEfEqsH29oEbKByO/Riutn5aLvfzAGm
lPaZDrR6kSba1UypOUw8fQOpLbw9nY++XU/kvCBE0I4RPrt4X23OXyBzQOVV
ka4t1lfSi3qOA3DTw3+po1PAhBuCpRSpHOXGbuhM12x+mJvAGcfEr6twEe46
VTaogcsL6FD9KWBpUiY8WJ+OY0H1ZlF7DUVc7CgUE/easeLIQeTrRnax33Go
1tN4naTcUZ6uax6FLjWbfov9z8LuOQDeoG283Rcw7UxRIoq3HAyTZdAWjwpU
hpbjDnhmrsViqbUFyMngvZ7jRcHoaX2bVt3r1nYfB+u0ZoIxSo6IR1WyMjJS
16oePmVTmx3XCyKyYWK7lmCX6qSbPPIwqpsWPX1n7x6ukEKeL6+svWKNj1qO
dcOCL+kVCzPUDEzVFISN1SZbp1iY9DZ7Gf+LL58Dl+JmNFtm6hhA7nSUgyZx
V+gkWBobyFJyl26B1h6dtDI7UazawxxrnDd4LTNKw8XSaX0FUEVIf7fbxfKy
XO3J/QXLykp0NmMuK1Un2jbT6lCZT8T98L+Hz9JrT8XX+5Wbbuvc3NIoMJvF
4ni1u6lt6vc13PHpRmwvgFzreckepwZ+ueNzcHUtQZOv6YmKdYmMwGcVhIMj
rvmP/6s45ei0Jhq74EkO8f7x8K1QhyiANToa9zSU25DytAUuLAso4hNkoZw1
MSgP3Qsk4KrfjfjW4o/67tpmAWlxoK1rnscLPly54DcDLjBcKabqNwSAZ+hr
6WRAgNZWvHgRcrsmUKPSeQoAD/m+x4oRibpZxdXzaZBAdioSq3q1Zt9evYad
t3EJb36stpNKlcMUmMbnxVKH45MyM0H1curiz/by3Q5YQRR1KLF8RsXYyjDb
aZmaufdQJmIlz+Vhj4vyQBCdry4bi/KouAGoDPintRP9Fvrsxf5IZDNl3Nyg
2uzlD2FCu00b2+opRCaBgiaTXvTnS0SwXLiPrhP/nc3qufav840cqVKLnG5z
vA9aqUcom52NN3SqicWraQ+KPOftK37DmttZX1mYycMMliW0XvVoU7HicQ1j
jwF4qoscWbNFaXEuSJdaCFeTR+f5Ay8pqepJNttkEC3VJq56I+tjVfTTRWCP
7Qvild1diEy09ou1LR9t39hUr2KnmYEuy2AsMlOsiHDB/hLfawCUJvGL87Pk
lElwvt6uClVQGiRGugxu/RNj0LWWv5gL7xqi+eqRUchAgNIpm5H10f77vF8y
IdQLQCHiS+feheYaxg4IOUTr62xv5msheriCtStP/8loeI3GJBmZGus+bBun
b2wGbZ916/DeyTxYKg2l8BcwObDxS9LajowIWaOMm+Ndou6JeWV27Y6DbRiw
sKn53rZYSfcfsUlIjtgLKaiekenfcDbr0D7RSSsCfsSZja4aekuDVJfn9uIj
mfSZ8Tcwunr4EStnJ3gkhhzTdvwn9hYzPN0OBBXdG6OpY1TaXgAmeXltTxnj
drnS9iFFsSfl5Fpph1qYwCswoYl0MqBTYBEWa2heH+xgHc6hMBklrd13bIy4
HpaFG1q78ahwcFtoj69qMVFluUtDWorbH7YTYkAvtOaEDTyLT4l8iDjjOjEz
PqI9XTnd2jB29oAujMgV5N99CyGyX6rITLoMWfUbrDuVop9vTddM2aS4seZM
38TXwePuHREZlzRAGOxOoQIIYmvgO7x543jZjWLi1cLo227fkPTEOqEr8/5Y
nXAH7b76eJ9PJ5uqXyr394lf9uPNzfouVgx1ZKRWxywaDCg4TTd6SN+uxaPl
H93xK7UFUmVLbxtKwa+q4p9aIUyuFvSyS2JKfL6nnSaBWTAbNjWC3QCOJUXy
TCZzQUVJZPX94h+LOmYDKVsOOAgJ8Sm4kATqBAqreSMMOmNGE1Bxsycp9Z5s
Sk4v19vI4yZnXQOkRqmoiNjaNK1jfgP6YtIAoIfITaLgplntqwaSV+o9ECDM
7RNH1BFMVKBKnd0J77r71ZFItxNsY4zGJBwh6xmZvxKihvWJXaY9g5B4fpWj
EYyOtYnmXzNddrD+YHnGa4mFIgUUBOky/AAQ8W12u3xlBAUALfMe+L4t+JQj
XQW7GjgjXZENzKzg/cnOa14Nulb04ezhOQKQSlAC4UQlFUspLnpnl8mQ7JLT
SXPfenWfseAyfDkZwkJTZQ7ksY7Ow/10lJ+HN0I3cu1mvi8yd8T+708fV6CL
fxboT9c6uDf/l7HnUxYVsu0rubWhRBlKhLb2+kLqYMU4c4xyqcvf39gXuWNC
AWEFkkWGXrko2duCDB1O/zrnBD2bmCslmvw97fNqmYCIU73gniSoLKoew6Me
JUbKD8ENOAwQws2I5VMrq/RCsNlAj4yAEJAYSmAXyybB8UTuGMyrIUR63zyf
/bnZvN+SEVyAZm9rPJk+z1RMnHz2Y0nXEnu+9PcI9gOM+X/2zTAVgpMyK2N7
YcZqgBmKozonQc/LeFItLbIMaYEOngrYuPkpd6FGTgnD691DC3GgoqUsgjAM
sPEU7TNjFi3PZo/6/IJbPu9raGLExzAbOAyqYcCozpBLEmTYnJyTm66mMwqk
Uxz9I2GrTqEKmHyeFaMpF6oPWxOkyccJ25277ejZRkP9TuGHJGhNBdtsiauI
jI25BW8AlvUbom7uZPTByIpOf1rJxgYUAC/9dhisjk5ay2EPQU/96MeGTRe7
sU/InxikTno4HxOTNojLvRWgZY/QM6a5z4DTk+DRNwIUziFMoe+ipSnIoBoA
df7aH87VtbEL2s9pwdofQjIenhF9LO1UV1AwQuwlRCzS1WcqsBpXQWz8Ls/N
MNDQbQgCRyArktVmpaoxV94YLQIMvPcLpxk1/yuKnuvv+B0UAliRE93NXBCI
NYb1YRMTNEe08UsSeOL84gCMThNUnb1WoIGebPQxRL1mCYt/mcauQ/4XFxas
tj6/zWheBkZbglPV0mmW6Iouq5a0NyVBGX5Ku9yEJFEiQ+cwyFbvIqrw7Dek
hAdeEUeOO4YnpnFHgxTfVw2aAVQfS4xWSeDODyKX2gfmrKfKgpx90knSjPIY
uuidJJ5wtQyyYuWLkZFRULoRHaCeexd0dwC1MD3qcHGziNig4yoqZf+4Vkxl
vw6Jdo0yCoTmM7F1Huqix4BT40jtGUD+ksD1LnpBdOhDCX87PQhlG6BMRB+r
Pqx4x417k2OW2SOrokEZxWo26l2d72biCwXSIUFYN9Cw53FcnD9u8RJg4lhX
B4LkqrUfuXfkK3VQKEKB9HAsw4pnN9AQ7hWvxp/rU4AVdNfvg+sdj88FBsOJ
bGvtl5i3SBZ7nCb2OMvw76l2N+5JOmpqZKLsEjECh2ILcJLh9ZlouDCjDeKP
ylkvuLrgSaqsVnJTJXetJSI5/WHbClsoFtkW1zRJbtILLv2YtdFa3IJEBzcf
Hnpw50hCe4czt8AQRO7oFPZcj2J7XD5fE7cUFlqDrv+RwHfbHIrsh7l4bj4V
dmONA13JE6yK1r251Mnebc+4V70sytwS8DNkh7FF4qR7bB7AOGgFmvMbs/oq
LDTotvoH5Y2WmgU6vtmbPcw7kjdRqIyvIdW9jkmUnqmOxI79Z/yG0EOw5vSA
0kSrGksjNiGCVNTW57rkosXAgFMeidi8GuJ0Uxt2+A/ilW7ufOh2DDt7WDHe
HriHRrT6H3744pbvZpEeyWafvbCG/rLc2ARlaTi6ddPPLLQdHWbLfMBq3ctd
XAkS/nYIMlGGTjvwYvUmNKmNEkFORUsYR+f+pCc3alklMJ/BCaoxEFkErjTH
yAMbexlh1rDgWAR6v5l5A/rfXaR+NGLM3sVBpZc4Av01jmgfNPYTS0G8bK5I
mTQldpgvDSIPu4gAdGuJlcYH3qkfRXPZgqnSZeBKxRavnCU2r0sbYAALkv2B
nmsoYkQNwtN6agYopgHNvnmtoSqUH9I1ApKgf1Pxyb8vH+ccKusy6xdyZFqQ
4CqtA1pCWJbpeCk8EdfxPukqIzyKKF1FrlPVN43iGZsOoedNjOAkV2w6nf79
0PwHs+A2vEOtSlSuUWKQ2C8f6SMjCFIObj1jVdC42HZypmALviX4vlznqbFe
7LDTzofo5mZgcjm+vKB973eWUi9/c2l2UghlZVCEP9jddPmoh+bn6LwW6xSI
GdGEY+YPNpT4w0/p9hcg5rpPoPNdJ104VX+gKFJuC4aSJ2DYsKnNOSfX4Ikz
khVSLG2DjlVWn0+t9LE0bO1F1xfrkOMfIfTwHz1Ifwq9TwmIuLYnpUhq5V/d
PrKZsUUWvocPbUaf450dDTEEii2og7G5IJIq8IBJwYg1j8BDi0LuMBSiZ+sE
NxoBu9p1auxepGqMKzhlUVERWMZKrHi1BvV4a3JxnmqOm44AF/PNOuqZKGTM
WcS5AgUdYcxi8bzjKMcyGmsTiTMp5SXnSwLIvhlqaDqflOUTMiV591ujlO4Y
sYdHE5yHnz4rKV/x3TaPnfiP0qJEeYzftaJ1GC+Ey9lzoWShNwdwCnfvc4vU
V3BT2d3eUMWqAKFVKaPhAw3tDxSJKBUCD4uZBiZvuM4vUCHQMhDasSzxGHkn
AFVni/Y7BtLT8e5hOHhvJEXzrlY0yHjo3ci/CuDNKXO59NQ/4vJeNNloXdkF
sEkeUZgk02TjURJh8hT8oJk0d+9vvigCueIETilrESYXqYnGVcFcU0+BlWBT
1pl++dvWVCVud98mCru05zWiyUxwfEaDj9Jvv+tf1MY6oxbeNTuGMRAT1TB/
TGyN2xgnaHH4nNi4Mx3+nx9LG2qBQxj638rCEjGpeU5UPQF1R0dKoHhd8tKp
aM8UorX+pCdTvZ4N2/wGf/07Eyg9iAHSHd2YVbmEGGvE2yagITY312y/+OeW
jqWutxGKaNOXG2iOGKyfWPRZ4JP8BafZ7x6NdHiCytEArzvmU7Ge02yLkqY4
jZ5W9FUe4afhNeG8sUeL69IOXb1Z7c/0+NznmvjAW1OjVJ5RcVSkFlUcYJ5H
jXoODA6aeM9wZOC/QiLuMBfXP//db3ZvSPu2Nb+iHQL0ysG+Zu6rIVcfQkvS
d4LtivBZy44MgE6w+v1RIAgph57vKnSfPoW9zezk3OgiIKHL+gtmkLtyHMOr
hHJ4S4xT4LgFlbdxqvqCoUXDcoLRncGpqrlrP1/TxLeTEybl6ImDtCeTbZju
O98M6F6YjQJsPdx97i0YRVFIIQO9ZhMj3UOwuZpsRcVAdsr/C2zV9ZLKrVyu
sKZxjwlAfPet9cX3Wj9LNWAcYhwedAIHwO/Hi+xYSevMrsr2JxN+vI65wi6h
fBiF+KigG6OJCbI3VMwRzYxV1kfHVntFyafSoaVLL6mqsyEgKlzcr6a6FtHc
ecO2TWFmWUf/hI2/17wN7xnY9/1WJsz/dDldqOZGW4+otfto0ctLJV3rVP+M
WLj47LgCaMnMQjcleZgzJj8KocgTpLnEEuuEM67olXAQGb77T9DUQLd5UI4N
iyWlp7Zg2aLsszWjcrk2Cve+XEXJdoL61/SSF34yrlZKuIMmQBcGp/X1TZOx
iBBzTvwxjuPG6QH6CHmjLYLMUFJZ2RK5y7RogWw31fa0IaXsr9YGQTsNw4Y2
Bshy5exePvHaZ0WGMGdxIubvtxIM0o1zai5C4/kWtS9NA/snGHzI/7/CjPIp
k4o5MilgogKqA4NGiGfl0k0TNGaxnijawxcuwjO1Xr+2+9XUYNrNT5uFARaJ
7V+Z5JoyY4J5JyVYB3EPEmErc1YPoXUYkU/ZHWsiU75uku+b4u7IMR2QCDdv
yPsADKs8hG10WfLKDsatipvmVZWMvfW35ce5Z++5kIPjEsrgX/xnmpTAaEsK
nSnz+Nxy/QcPoH2ZeMLAsJkvvZeuLm7471nEoITZ9DO50eArqPi8zGiZ2Ctc
eoNaknT+ZK/tx235qKM3A2UcKs0hlZG32TWk8V7AOU9rGayi3TShkNehQtAG
LneFK/2Y0O4E8W931flgC1L3o7KS6wgjRQST7JA75hB2jYewiAuXL3wdI3lM
9NWZDQKdFGO4QF5InNO7VlNyqA2v2DBa4aOCfbbYHiFxiyBatBD1xSaLzQey
F3ODTF3EKyBCPLBaMg7nMicxtJ55lxhovxN7irgidCBvh8Ic50aNnaRJ2LaE
W8z7GGq7k6fTlaTGS+eCGmxoc1XdhwlDWN9luX5oEOyOz7DTaJdpOaVooV/o
EUDzzAORym1QUgUfj8zGJNoZtFtp6N4lFWA8g5fAlH7Lh081hIcxorJm7i8d
DSkRKtyDc2lJToBLahgw10/jKDHqUNQNioEJlxMkhtHtaJIR8uH6lNa32xkh
WFOeWIuKrklMGjVVlwOiIEe5rsoAXA4Gkw+Jhl+n+i2AZ3rXxSExCUbHGpHt
zvPOKmNNBVd+EElgK/XYSbBfIbCbf76D1MFaBGEG0Bd0uMrEZ4i1L7tNJKQQ
ZBmfdk2beiEjkWD0/Bkpm580ZRuK116RMRuaXFIwn7YkrnyRl/zfVRhMIOUV
JPbtriooIlJhZ0qD4MHbdFzqV7/cuycqMCp1uwFffKxIDTS7YfQMveQtnjsa
aA+HDFJ8oZkTy2aiSFPSL/vV5F/YKe40TGyZqs2YjlNBMgKe/J/qhDRhR+wh
BTnosob4APgixyjsw+UbV1ji94eBWFNwEdZqKHlDiTm/wHyZTkp8tOnv8kfn
RjRTbfYzsxjNFQv9ZNR+aVa6BDhAnfJhDUD1WbRQrkY3mmDUgGzfgKvs2156
ZC1OI5+vjAKTKLazFAAGHwSghXzXz1u+bk/M8JYvN8jhtbdp6XmLC6AaGKog
soxbmaFvY/jaCCyOiMVPcIT0WpDfmVLz+OsWCKC5oqYOae73KAEiMkB1m4G6
Mb4sFH+Y8pqXZfJE0DLCukhCV4xmQBGyGIqR4HdZQSCu/M2gmWRPgSVuKpWa
36bYez4qT3K8yrUmtvmnppguHMQ7vuRvJ8nKVNBatyL4w5zIio0Pjwz1C4zj
gBX6kSMW7V9lkODi4+gGP2FinEj3Mobq/9+kx8CItKYtA0WmPkRIcZGpxPCO
MxnjV/Oss/ajLXz+xHJEdYxN1FYkCHkyfl3VFu4qCTIZTHv7T83hxu8/Q/pl
B6CbfPdV5yYwwPGXLPA1Qx/6Wyy3GhkN8OPGMKZ8noV0qWGPDTMNA3Pzy9S4
ixxGG1FYi8T6L51YLnJf1pkWDe8WTT8jMQIp9aUkWPlUSFc27l/espqU8jpZ
ODdnpM7nyDMBE34XrMgncvFj6GwzzNMpELJHFy2oFan1+yQBXJj/FdLGvQcQ
5/umciL4ianIYqNkcUa7a2K7L1/ITkx1IF8TII/xph02+z6pVCUeGj0p+jZH
DBu66D8tiJlqCngya3Uu1z2Mz8Q+eTsSHQVeanL/4jKnBV1hlNNR3qF8Zj2z
6NJGo+yO7ziVH3O32DcHgaTi2vOXJgWID798iHQ8QQSdzxw95Jt8GQvJGN8G
uSgMxdz3PpMoUd2+Do9f8/dsWvC6ulyEDBpRA1ZMfrTdXUcUu54N3dcQ0wni
bFCfqU6q9Ldc0rucsbLVQ86g0o/4+TzgRu9wiebCarjTsME+DjwzAXocAr0l
lzxRSY6axVlJAEAzAXnSJPOqUz0EBxCqJ1vwPh3p5lOAeeQleKW7nbYEkf9l
dOCU+tPdz1cPHiOcw5C2E1D6qzGdJeJpxo70n6lg7ByfOrA15CavCi4W4lpL
IxA3j5QZ+CVHjuh21qom+HtcCpgE30hZAAtIEhgrTs47iTeJEwjoVamU8IZp
c/ui0z+KvIxutKQU+nRhwOm0vho80TVu3U57fF1Labb0AfkdA67J1gb1AWgP
CNhrGYpMd1pV7oKkCUODPkqA2yUz8bxsKrkLLiyIfJbCP0IHgg6Ymy9FkXOG
OYVtk/77D0Wk9ZfbcotKh9HEweENLk1B3OBqb6nwanv49fn9vC9Je6RIR3sn
HaR+26hTTUb4K8zwRyh1dTvKkh/L3UQVMWxMLl10RJpSYbTwhejhHNKwwip/
ah+KlvHKgPqjnlVnAYrZ7YkkPjrHlBlTY0Y6RjzHUXDJKH4zp5mcWz6EzV5Z
TA8ZLV67OYTVZ/8DhrBKJnBs9Phfe4ChGu43rJ4KHFMK0XSy3M8S7d3R799L
fa7KTz6a8dKSRwGdbfSB+7DPVlBMtSliAAR6tpNMAdxPM5AZF4G0xVihnMQf
7MTKh2W4wSKmsonkAs9IKhQWX48X6yYvPD5VPBnAXZB///jMDpw0GIS4e5N2
olREzTcqLZrQLVKqt7TqtDjGB/ifKhEEs+oedXK9a55IC5VuPBRP0mvmkRIW
ijIRgybHPaMH43rzSbWkVFrYuG9crvZ3sI18um/APTUR6raE/Y6Drxc1Dt2h
13WW8WEIgmh5VKxysfYkX/9bMXuXI3k65bvqn9+4jbpzuwTQfoTDa0hHqvQp
1zCn3n8vjdvPpmbOgkaEZWVOGWuUCOJ62nFVQnoRDAfXg15J17mDPJhUYO3n
cgnIKTF+QeONNkZrmBWj5jkUaGS+81DMY0FE2lWAN5NZl3yBRoJNWmse3HQz
dLQvpQArc7n42us8MIjBJqDaji88bDcEj6FbMn/jCJeXfBArPQxqXkZ6Hc1B
QsB8fV0djlHpFPgIndESS3I4dOmXcATLl6wguTNtISeLRGDQnqjNih3iu9Hy
LybTHllHUvpWyqgMg8aqGvqTfb7U7t8uRv6cOx1JZWs0+65vJmxOEsun0gIG
MXYVqnl5+pqO5M52GB2n22ydc0dLNgRSZEGiU/NMCKTqVePYFBfVKd0163F2
acXWGLriFTi1lWrvJfLExpolTA52eeFNOMb9gtWUBlgwWcTgwjZU39GtTnxe
3SCsupumDpSv38tR54LflNhVJphuc+nGmPMmxYvLBJt7lzWVXk1fgwXjuLkV
dJEEkMDCKyG67H87aBkOd+yFROcZfxvFITFXDX6vBuFWrcE6P4EY7Pt0dNzs
HpsLw3PC5nx755jWd+XGNc54Ta4cORbOt9RfxYOQ0JeHoHH06V2yjqkomXAq
/t+a6FAur+WZhP/F+rcvqM4u08zj4cxLGb7UiV6RXNZ+O3jK7xipbEcCHuO3
MGkTp/U0BCLbe6lcDKox0fN4JOfrhrcI1JyMWoVG2dRZfbUVpM2Nz62w6xuh
lBYxEAd3Hk6YQksOmGQ6tFPiw+PS1/Q4o+x99H1dCL2geBFqLHGdLFm+MTQD
ye54eVJgsOXdf108Bz1JiBIBtJf+2pIbRm/V9tDBQvO1wU8dGDhV2d8rL7Vw
MdChkDz7Aca2wpxhqjpmCBoz9FagjoNDGacuIRSkGmtIGV9eO0g/Ii1lXXqh
b0Pra4jJGs6Lo089qEqYun0uSxXmr+5bAD+ELu9EknwElTsj6J7oF7d4lEza
bCEF7J2b7ofqY4ut+IUfNF/qMQbrO3nkYAtwoEbCriQJzYdnq+bRv0P9/GDl
yVhCXGk8hf7bpeSU7404vDJ99y6FJLLE8+6PYL1qY3taFhoRiYUrNgZkkFoW
Wqrn/IH7Bzb9olWgdFE/tEo9/sDrOy52TFyAibVOOz17BSwyF0dG6o2m8T7i
juLe9X2u8pAVOPhdyPxhODDxl5q6+Vi7OrBCWuJ87pBIdR9XZ5LjjRVY9YKH
T88PjPN4GYZFIzW5j12RxarXiGpFBxn580o8/fQ5Ya9+xnKlQ0iqCf+Xoak0
PRUW/cAF/QSydA2sUyQK5U5K9wc7Knb63HKdc2THxcVhBZ9TSponP+TpjO/N
fWIrub28PW8pfxf5W5E5TG9hKOATnJNXWeAZothoT9HQUcyMTfMaxePW3T9S
HUzd44j9njpP1v+fSLLSP6ZfTOedtVk9ke0p5o0iDU0753XvZypiGW/fzkAf
i5Gg9u7Xtp4ZvC7WYwTwdnwbW5WEx7XDCk0TB/gAQJOCWhw+oOOB5YaCHpPJ
R2NHZ37FUMix8i5vM4bgh7XChOnvlhu+7capU3Nhzdbx3I37UQuoActg/z3o
DHe93dhWBR15sd6/7bHa2xGGMD2gx75CaZ62vfVttPgZlwLvg9vXjBzNzRdp
H6qe3yN+4zznmNb36rXJrW3KldJX6aHhsz2T/bDmT4Dh4tVFnoOymVI0GLcl
7lpHFqFJ92aJpfbZKJ+3OEpML7l7Q0KMwTb9UHasJn7IWfpeNJ1x0IxHFgSz
3K1dLIjchLlRZJeNm+E5TtUijjgqa9r8sUFFg8dUv1+zZa1ie0clNPiqIdW4
yVdHgQjJv6JQC1FA+I0FS+Q6yogqxCRqv4iXySDsNE4dk3N+dnYqZApxGJL4
OdG82nnT8g4C7PszZgM1RiTrzlSuL4SN9ezkineA33eJwyX7fg3p3t0JHTnY
ApSbUHHshz4VSHJBh6xQ0k0zwj2IkKeehNiW9ir03sA4pwmdnrWNu6eQNfu4
JVIrv2bkzlLeWdGu051FrtU6zx5q0MDuhfOgYFuewBWcqULYNgTmNIKUAKm5
BsTEgSvIchslXCXevMgZOzLE5gfp8T93hFyIx6XehwV1994eJ5QrEMIUvfiH
a1Wk1Rfin25Jk9SoeYsXHDu5Go0xJkHjKCTIHLfr88n0YOWTkqAUS22Q6XOa
N6JFGwDhcyS3DCMOMvpVb0DnVX4gpepAbRbsK9jvdue4jcXbGFyQQE2eb8wl
GFd5LmNghC5Jc1cLNlL5Q+TBmYkwwgP9Ur4Id96vmMLiC3uWJT8eoz/Mp7j/
4SQOXwIHU3BSWSb+pG5t+aAgM6yAH3cfdAZKDoReeW76+Iqunnpiok3EUeH0
pUnjp5L3DGvOsU0iX8JiY/lvXvutBCTn7YU+Wl8DS3wl9wUoUXmxJsD/GVlE
++eatGu6YMh2DYAtMrwDkfazsoJb2ApBMvUHeJlxXfHZgjKhN77ZlSfBVKjU
oBX0MpZL1Is257d08+LMvbD3v43hBGUbJbLWb3OtHwATBijewA7QyyqCA165
pWVQ0czOP9htdGt5zPp6Tjd+smlphzQHODavLo61WaCneLiX9lpA0hJOFoIt
IM9LFi2t4XF4sEZttVZkqSnrqvqZAtSdVX/AR5lLehITmeKgfc49uN2ui+tD
c3mkGI46H01PAVkqpINUBCF74DlhSHzXvuXskXUDIg4VR/YFiUyWeACgrvBq
1T293NwRRx3lX0N969AzPQQ0BjnwF/HQrbBwet+gOL05abea8yTLh9OSUpe3
nbFccSZIv4np1fnd0FW0f5sVqDTTZm0BTM8pTtEX6Yk0es7kh3zMojwF6faX
aZKQBl7FRWTD3AiOp2DAnz9oO6gA7KJaIu932ZrsbSBQnPOg4FTwMFY8d86e
5ig7HSigxGPDKjXRjzD9KqY9eQ+uolze3XtQscypbfvm2a+4Ch9o05PnMfoZ
CZ9IG9u1ObefoE4voFQahv0JCRzzDwjo5fGei3Tnfe1whksEbQ8q0T+Q2ETk
kRLbJiPpAMSqWYKIDdgkzQOnP+FkpuKLy6anm468lbvpv7HEcpq514GFENkf
ygoJEEtckWBXN6nMC3FiJvM7Ax1iPTygtgroNgxio5mqaXMnmj0RvZTNMCBP
Q3WHvxXc2dTBK1j4fi/Tx9obatWOePsJNMvxYlXalpnpdWNqLyyoT8hEgDlS
flfvow3Gm/KScoPME1EzJ5vO2wpo+VAX0ipvvLs4sq9LloFCouIXeguWx7H5
4xmbgef5swI4FxAGairG+HGUSzvMGt9TVZCBvHKUuhurKgaJ5JR5z3x1HUU8
QQyTXsQowWT1O1AGzgYZVNFNNoHd3vFEOPpnskbxIxmYRqe7+FmuUoPdGv/y
1G87cI91eY+Yw0pczzS/8IKpe218+b+Jl6qpmDtZv4a4fdC5b5QwqaFQwYgs
QgYKSt2otKicX0IOzwG3r2aXwIGTbrIO5k7ueOrMtH3qEO93lHgW8W4gFjE/
E7iBSyhqvyUuJcwGUluwXmkk0r7a7zLMinaKSKVcfaJOXCrX6mvp4L1CMxnp
1QAYdUGY+YkWai226IhjVPqdBwgdDH0GBgW9nIfaenrSiKNAsm0levJUSg28
vF1W+rxmWbeMF7Jm7D2O+FaqHhHnMbrBdrqcJI/1n1ut4Z2hwAZmApzJIkMP
TVhTVcoERLieWGFbglf1Ax/+ptVX/0rLMYeUDj1nxVAqNrIrLnhaRXbJPjHW
UR6ly287t09BZa8L4OcasOHjFc11uteV5OBVP0V1SFoUNo5cnCo4egUu0I0u
kIBI/oVurl8iRRJkfTKaD7cONWr9hzmQVoVj+7N050aJFQWjoI0U/iOrLHW7
6KGTmF19A2b8M8UHTH/td/Wgeq84lpEMHwSXMhS8ZLPbu0EFQtRWr/njXq2y
OiSHJQ0rBJMTCNRCZ5n9RzvNL7IqlvHlj3vTuSHcP50qMnw/pA3oBYyhpKjL
d64/1TUhyOOFEVAS8nJFTdiPaTiSa3RYaRfQo5bjUM+/ijZA9OSWaLh9Wd5b
ISceKWWkgS8aRpRRGjJKTxt7lrTwGWVW3qY6O2FXry80UmlQKH1N4Ocr6aaa
0/mx3wAfGfr9YZeFL30/gP/2Qa0zCelnIYcAr3h23PvMvNgV5+69lJLlPafQ
YqQ55lOAPWG00TKPbqy5H94mPtlHMuvfvjkzi4qbkJfsQ9HUAyAVqU+eTf0q
a/QJmpLe5RW0lvS8s4ThEXGBy+P6buAejCYfo50gOwDgMtIxIY0rCIezvdBi
j2GEfp4xwMuDhDeRAszybujPOWG6q+5VEVyveEoisIO3f7aa8GvnHoBUH8dK
A7KMEDqDMMLF3hObIgR0j8q3K35W8nTkkJ2dhjWKbjDnJfyNJQ+YnT+Y0osN
AiGTaod3ZxSLvuldjNjqrR/Y8O2UR4tBibQ7fsGjwqP9o9x/er/ax2XBQgJk
UZyVXbvwhpCtHhDS2eFDCAGHQcX4tkExlCIyrnoa1TJPLM2vi2KeahnBPaqD
4QNy2gr1tbNYJUNfyVX+tovW3rAPwSpOR2Fr2WBRY8NR2AzcGWafwLN3Up8g
InNRrHlOILHGQKUXLZ1E3eaG1B34VJJO3EjXKEWkZpA5wC0U40HxUpzFSR+t
qE/foxMIXIB1c+zBlPpDhVQXt49zibht1bXp25VJTDmT85x11Bxrqq10zhdQ
j91rETE3xBULIDKv7Nz/7LWwrgGCGrwuFSjQMtUCVjAHNLEwMYTMO0Zj9Llh
CJF09Kx0kO3xNocMnKsomF4Dq0Ixre+SdYui1t7pl6i1WTazxbzzrlOtcbHu
qRv870u3/mGpdhQHnM+Jtj7I2FH4UGsjWqkErd5Zzu6dLjxadsC/c2q81Sgb
HBy5OTqlUd4hapGykPvUcGd86BxxuITLWk8mX6+QIHSRVUduJFslhjl/mmtE
1xOo3962FcP7elha6xuG1K4f/60y3LHKVUXG6MQ1MGKUYZgYf/VorNbzqTIr
uXAmzsUzkFftFWVD7A512CGRY4wuE2RlNHCu1nH1pnUdgrbaVaTxb0J7Wqaq
/ZCxpaN4hjhP6yvw/MNbJnn1rzkDLjD6uHxneRoqpkq7x6suw9OD4YRmqbp1
a4weHvRhWUo7VcXN+tewQxRlTQgRSArEvZbgy5czC59sE/a0J7PA8VLrR+Zt
a+xnagzcmePVZjdEmKgRBS0kAmo6PwIjO11LSmfc2kYepD3JrcJE9Mx6ApbU
5o4puYHNXq84pKzhUmg0ttRtcCSPPcZ1ry3Z5EWnr7rasj9ZyaXcPflNifgO
NTl+tYRH1uNodGzmF2P/EixbYOjMxo0RhtyI4Fv9lgTT+kGwrIzXUPPFYLHP
7fFlkY/D2MwtMImwlVHPGfbPFHKXmsNKApe0jjlPUTkEQn9eam2voilSOmUB
14tFkpTVypGyrSF74BUDCzBTo4io6m5gDqpFxphB1KyCYVGWR4cXXNq+/ACb
KNmwKXgYUZCn/e3tkgq8P98MUUjRSlRpwfcMpCpi8T0AG5M2D1+GqjUdwDle
7iEdmOi1xT+e+DENaVfdnhSZSNymYi00iJnioB/6+1eVCFAYZtgHNACD60Mt
GLGFRYfoFyOKY2R5bLCvGv5nzVZ6exD6Cizu86ECm/FXpghKcC81/0lkwRic
tkm2s0HUkmXohOMNJTnUtTZdb/VqgkYlH+ywjMhq4XHqtUAgs2mmrCkSadac
qeaVg34rfToA9o+HwgNjgCZ8uUlpStv6IFLo/vTukHbkaadlD6ZmphBtCFnR
y7WWYkJHbt1sOy+VM/28otqV9Q3dGrbE1hyeqGilima9YRGRw9/I9CGAa/Io
810RFqyUIPcNQjXBhoegXGqyv1ZNjy+KUBIxjUCqo7IDtf0xXMlMpaSzuSAs
6C/1Tq4Krw+tbwefipyRsDdQvgK9th93xPXn3YbNKBET2VVBRTCiLPFoKTTw
5HqIe+0JAGBejEfihx45tV8ew2xcXngJYRac0CrPADlq5f/bCdSglaljWOHc
YwSsV6B4lBjSIQIBg8/V935+RWC2Idba4CnM3uu0k3rEIgdUnClMs/AyYm3+
amUR0Tj4rBMsrIKnRjxFoY2wvE/vIuzIR4GsfqLDtPv5jJHvZRiB5H/866ZQ
ilqefPUmqr9XkEAu7XLfERZfBbGeM+ThOLcLfAn4qpdgRt9cDJeE2k43T07H
WduPZ20tSpWhurZ0Xl+Mx+olnqEpdVp++sadTNCIFBGHftQrVK2+jgq8Snjz
ITaIcrfaDzUyPMuto98sDcurd9oOxVM52Pf832B415Ontf1lxof5QbiDDUWV
VNo4OXLja0kkCgxRzA8V2sR2sX2L0mv7OpEjsitPs4CBOsYCqSrHkr4La/j5
VnYOtn/my9SNHRrfTXEALa2FusVewCF/SiZUnhj0sZI/hIAQQ9DLJ970eS4h
c4x1jMGDtbh29S8+/gD0vtYpY+Iy/rLXsIZaQAaFNSbW1mzsmJ3WyVdvtZfw
wUWUiR+4C/xAWB71vtjt8AV9bHbdiUa4qG2P23zZgs3P38FfsIfqRR6bfOSC
IiuMV6L4MTQZqb9O5cOVAhJ/en1GGOlgG2V0gJnPzmUbUXq4J+3c30QQJTQW
hVw6+o95aph2ZUa2ewogJegTKkvgRjfkF9djPhLe1QH1mEJF50ZnYr1Zs0J9
ntM1GtQlMCEwFKQ6ewzdajv8seI0KiO+yQHW++kZSkIB8bozpwQdcGAauDno
0k0/YMEqRcIi6JpW50FhmJMbeoj/P1/8BL/Wkj5MYuP8lkjypBxQQIbl+O/s
Wy40ZGC2dj5yaUKAAqipM86JciPdQ4JSei/l/tQ5agRHGX88/m7YBajgazR0
1JKV+np+RIM+8wxVDfTZIosqrl1qLbwsNRg2XcKmahPnyHzliJxjMMfGJAYX
vVcmB1EV4l9yKgqHEYyktLlzGN68DzEwyQPVynVt5z6It5Un7JmabFSP5bZU
YiQxJf3kCv2i2gRYdf8nFCmrPPjpZFlDnpa1XAtaiMuuEflEhOWXb4i/iize
12b3b9gw26P0y1aU1FYB/8PgGi6dbh8luPgfXxA3cwBGGC56CaBewntModPr
udnSBd03IIeh3/fqxR4ZhWgahDZhrSDtQQDARmCV9cSCvTTsGE+cuC2og92R
Gs9om8tfEEJfvY0gJhppy0xie2izdRW4yldziluUWgJf8aadquJe8f+s4RKE
rwBp0yxNIqifpkZpF5/K7FjppP0Z8RNjZL4hga17LMJdjPvtzunaKeQroJSs
xM568urrvwsjJMccTFZnKjjG7jqaKvYbDdXPdCP3dfzgqCxKAuG8xRfXDMJb
+aKBKZEI9aWhJdqCnqR/yfyrFA2OE5bH5EyEiasswbQXyBqQED//WBymZG+K
/Sj8Yi6Hldlh/yyzwy1rMg7d8FMBDZaiL/0DBOsIbSYL/ZSL37b92awl81lP
s3YBFHAt6nT9v8MJyT2ILQ3sl58z8dZBwfJswTZLiU7RNciOY6QHSX0mum8B
VlU59uRZkDORugeEBeQp1kv0sOr8g9mCH23Oiru5i/wGxI8RdkEPqA6Wi7tw
8DQxqGjYtNTe+pcb1tDtiwIfcv8vcUbQeMt3u5KV9BhRK1MqC5xs58kyUa8S
Y/sLXIGU7mG2tmKqHNFZ+E/F5svPbi95L2L+DtS2lpec9z1QOvIclmsBMooD
LPsBnc/KCBqaEVHUNchT9RlERLEF676jZ6szkMfJULFoCa0ZFuskCWLwFuxZ
65phZYvCLiGnFh94OQq3WNmb0LbFUzwRXNSuKjqD3mF9WZ5lJEuBPZIFjXf8
7zOfbjcbTC9yfuhj50d6lT6Q1ZBo1YYxbHyct4Ib9jzZQbTrWKCxZtF+s15K
xK8T9pJYYAcSyRf16UbaObbxwXHIQRakfJ6yFsmPEydCmkQP5TmiCik4bY8n
62AjqibOqCdTfhGdKz0xjLk3ebVbRuLmyAwO639Pi+512TfrVMVf3Y7rFynI
wB3PLt6etDE6roV84PsdIz6VBnsJcVCqdcFZnJb+QnIjMrrm/lF9eNoY0VGP
i/oyBT4r4I6cOaUCdFAZ0KqN2Ko8NAuKLxufbidR0ab+DDmAj30a1JOsUDaQ
bG87w6GocKxg99X6Cit9bB5v0U5vlwnTc55dkSlQHiFtARIrML0V/i0bwDQh
WWB5TNX6KrkBJ9dO9dp+v8NQ3e5wdNQCzV/X12aUhUiiIAThHPzK75Lk1xV1
hgI38N/h7zvDZW2ufO9wbZssn2ffgvKn5I2hXXcEdex0t1LCsSfh1D6Od+qp
yq8frSuxST36ythGR7Gf0H0D1JrWdlys4f92jYMiWI04vLZ/odlsFlXMZvHt
dtuAvdCNdEOCO8svk/tgPhRjD9JtJnkSafmpl1jk2nlQOaUqzrxjIm1GWo9G
isGi+Wul/MBVFib4jezR10V+2PHcTDHDc2vvo/Fu5wWHxR0Utg9amgcMRrls
+TvEyf84L3CxkPsW9i0dcAKJHeEuAjeNM3BUB4OwJMG8KiiGkoeEbf4J59EH
pIm8fuCvDjR7CgWNpORIZM5m7vbcTyWGaOKVfGz1TjI5HUwV9Guh6GrvXUvn
Y5Fa6vHBu6/EMF99m7Ns+BeU1D63LLEqdS09VNwUMIopNWfHjYmVJkA8bFy5
XzC0eQNaYYie4WmMp8OMCRwrJ89lm7UdtIC6IGT00BoO+ewMM3hHWC+cEnNS
9oSTMNzXu56GbreSoSK61ydIsDi9ZXib0EJSOiBWh7tPFKhYBSXxNOV4/bBd
iPEc5sCP/0aFYEREi/d00kqK6eNZTkrtvtAyNBM7qor3ggkhym1qBYp6yBm8
UEGV3HGGJbsz35QyhqGCZn5ze32GqIw4c+IN9GdfW3y19N1ZV8A8eBOGoBWV
sCC1R4KuaqpczMEu+CHppV/g0L5Zcz+qs2a5mlq4KCw5t1HndjlGQGyhgxoI
ht6JW6n+g4Pu34QExO0zbuNvlqDnUEN9Yp96OIUVPBibkD5r9pOht2RDa8E5
a8B7tcECcDr7//jijzfjIgGpO7nxnz5ZJMZBJ7+wt0H3ysdSPXfRe5bkzfDF
9zIzQ/ZlGGgwl1CWTrX8E/bJX8yvD06t55SeoictNxy8ac4nGjoJzBSp8mcz
k522oQBpAExh2RIagkeLvf2IbVzxVqedr4w0xz3gxO9WPWBHfizZV8A23+yM
smTdAP+CO99FpheqgU/v6UO4NBHxblnVeuTDQ4aw3SUj2Z1MG8hEisxDTHBY
ven+H21K4KnwnC6zhviDc7Xa96Z0Ry0kRvGdCfxf/0dGLkCrNlLHaRrcx7Ox
is2DS08LxE7hZjns14FocOxVVWYml5sN2+QE7ezhcBUqEE/TycqJ8ZwQzeBB
ugZ5fc+1NsP/w6hXELetz7cD9EgeOvh/xJi1E3VEFwtL8iipFN+Lx+lMaa16
pV+Bhvzszf0Zm0BZfyA3kzWkpQsUHgQTwPY4eluXc+g0ipQxgQMum7/xvaYK
pW32gAxPM8ARa9XPobI5KPzCJ0cLQDbXCBcmjnBplnGYS5ahLzJFMF+G7XAq
CeMUXPy+zXcLupGSkHBJcs5fHo/clnNp4iNSpaA1jlQl9wMNTb+qqYwTKj+c
lJ37sOsNh2LZl/PHoRLsZP9M8TfVr0TQe6HtEDrZWseWU3zQyckJRef1oeWX
5J33nTAOPjx6an3WQY8kExSWE0JOPHgUrAVnfwm6SVTkGqvk5KojLGLB54ds
6Tq82or/P9vgvwVuY4Qpe5ujDq26kjhS0flsdFNf19Rl54mYrI0IpnMI+eiP
4Hm2p+eT7Z6/iyInk4VG4nz4Ia7HbmxbG22YwK8Jx+Au7AumjYX3xpzThZj7
OnJ4mBJ1SDn8JQblweanuzRUztR379R7fxslZFI4w9iWdEdbl51WGWLCg3iZ
fGeMOeDuRM/xdDwyDDvuKgUAF+Xi/mkXd3R6WkNBJ9z5ikZR4E9r5WzNejYg
4yTcbjb3sKd6Gzm1lfaq48cG8q2w04KaaBgT6HAScsqTAnJNH5OkTQogNGK/
zknvP9DHQhXvwJtXJaJQ06lE3Ka//42OZVjWN+O0QX+k/xqVkWFfxl3XeK03
NSHQHUOEYlLwu+NgERAqnOsUlvOZAeit78kQfIfVgStVLQ78aXux/RSFeZqQ
mx7aOBN3H5HwOjm6xglmooeVoe6QNJw3OH3J2A4nIQS+cuBYfEdGmaVgIA7o
qsTF1r69WW7gPH+64ny6LJhbgjcjGJ6Rk++ddacAgARmzUWv+AG8cAVtivr+
pgUxdAP7rndYyoLhjz6ApOwNevWBpTC/U7G8WVmGzDGmdeM+I4C4jj3C0gln
k7XC6xiqIrsencgIKd3MFWKvn/H7jZhdyH8G8++eXxV7tL2MoS3ygdQrlrLK
vhh4mluTSGeDsazzJDBdjj2OhTcBQnw4a0xNgoc7mPe7WtYxBiYAIdZzza8b
DAp5z4V/9eAoxK08erSxq8a01BCYMI8LF0tfOS1ZRIzoQ9UY6kFGJG5/AM7N
UJ2lV0TpS/Me3fIoHOk3JM+q8U0UxXL0iP2i2PepnvfYFiWOARRTL7lTVScO
XhW9MZLXRTXcVNx67Om3gfRBGlw5jqLyPxdJ23xTU4XljXKKInRpD7CuEJBc
TC5ahVSan/rCW9yIGYUorfc4et5RTR6C5Xt6b0EbLAZ4k08AmiYlA3ezbpak
O9Oz+ifk0dZgaFOyEFQL3naPy+mhjXbNdK4tasm9aOqK+UHLrnj8Tix64IZy
ie+DYQVsggYrHaxSQ4hxRkz1QNY0ENwf70kPniohfqV80lQ30ixvVmzb94cQ
pOBtUct+L1MO1HST/1wySXV6qS32gSyW+XEk4BytJiysQqAAv7TpRinRONNE
PX0q080qYM/nMSCEBIam+XJ2LMr2mCWRiNeWQ0/OGToGzw4Ch40GEuKhHErB
AAN9RcvSIg8zHC5OWoutUsqzYiUORGKbOxDwnMsnFEv5oWeXkPWs9RrCXZB1
VoENsc88LkI8rgJM/vkD/j3+givihp/KQ4Pc2Ucpavr6xE4UavGlp7KaZvAW
lQqHcXFGCGcPljPIiEDqddgvtyRcshWAYzxVQphCaqWtqB4Z+w83CKvRwzi2
cPnfo8vfkvVD+KujZ+F06wFEmPbrzPZ2zHHYV91uZaZajtDxFc9R/gTh7F8g
0vLfJ5ANOrhp+ryUBTH2pUSqKW/2oeGXoS1gn+dMAw+W8GEB3blaUaOdIhRh
bl1m11YcoqyNccnWi0JP6Rh+Z54zte92zOswQr4NEuNUtSZt25DFtpzGaIvG
+fyYVB04yKYdO1Sso4I2vCGBHw6N50Ke5uEX0FbWlLxJZZTCt1JXfjPrs2Zu
0IpGSM6+QF9tpRwzEbGwpsfYuF2JNWSbeLzWvW6zbqjAAZVY2B3HQ7/6I6qR
QBQAFCuLU2ktE8f7ZuRN2qbNehP5knkrXoF4Bah1fNDA77/yrN6e1HoMCGW+
lVsQZcUDseo4k4UAce+2J8X13pf3Fo3B5mKeZZPED9ROJhRRYO62JToxkjzO
0XTNYmEoIsJlBAxJjF3giQFvll0d3Q3viQUuv58YCRBFvcZdjDqSzxdM6eI5
r39yOWrH3T9gklaf8QAWRDRHfeI61bzwuJXQoj2Hm94LdP1cbt4AT3/GPwyJ
vzDUQ0K4FC9L5roGhT+yS2G9CK0S9QlEG5wEmrbvcrtb8vnvbKwEwBNCNAlH
l2YHH7d6Rg0jejQuI/heCcsiWt7d624jRnp+jfWtXVslgkSaK91qOwQ2NiTp
ktDWA1DpKBa6M0myXCa2BoTZCHFGayNdM7EMs9IQN9ixWOmO3oKH2yRVgQZY
7GBKrcVgFB1Vu6hCsk+O0B645OcDUYzH0SJ2UpZbN3DqBXgXkB/mxT9vkmdQ
TSnpXnRGzL6vk1YTjWIE0bPnESVF3hQQUdwxSkj8MnopCFz9IiG55EOZQxLB
C0vqY0ijQQDpxOVy3uLGQrRbmvwMQouZeNhWUZvK7aIrxY8JmQkUdwBFVGZG
ND4QhWG/2x6C+AVcD2xUZyQhjWL7kOLsF0WQZMwNNqiSr85cK4XVHI3ysyY0
BBYjTTq6pcfNrXn3kufpZ+3iTH9FCXhXCHOMvx5XNsztiZBttIRvHtoOtqEu
zLHip3DFwQjDMtz3KuEChwZqjFbDhQylqbLpfm7gDyzUG5xpWcyHBtrFgB3h
r3mmdHHwyjMZXdS2FImz1YdUxJqmcUJYEW5cv2d4iy+hmb6p3YpP3saYpa3K
TqG9Kc6IZQ+or6WigigTCww9FrU8S8DQLEwxT/b8l/uliEuNX4sD9WxWmSjw
PT7ca4v5IhhHZ8TUrK8Rv1S4UHtCK5PBKj8dq2VRXZuKb/i06FLI6KD533dc
8DPYdBIiT1he5qpJ1ZmIC3hIRJaWeuVJGeU4O9+gylMlO11MlzG/AuNC8akz
whOapve+2vGrC8IIoSB/d8IT/slanQjV43vVo0huJRJn5lBMtBeZZj5Np+Pp
b814m3Kf2vJz+zED20pFRuuqEqbhkpDrGs6+FhQTLNuD2q1QZeDLI6Nt11v8
YOXJdAFE/lObI+xbZUfbouDZqrhvSXzIE/WbeaYrGk60NqdSLoo0cVpQ5jSA
MC8eWMI8yRPAO2GgF2pyKIojfNd8FxnKcWtgGGBxymgcviq2ljjk2HM78fYH
blZbgSWCun+IK05bJCnHien3VszQBgIyRkSMhlQan1FRQ7KLihTm3V1uHIMm
pKYCZ2jvco5Z9qFxmQW33phHl1CacjRQujyVzKY02E9nMkY6gU30uLsUcFk0
KZjDlAbaRtpvT6kz5KFwC4Dw+kgyFPyIVZ0zQGMxb6ugFYlDWMZC69CHDaYc
A/p4D6YKWWGK05UWxn3gdUugRLG2ucz22Hsi7eS93GjM7fTxtZ8axs3/SqZ8
F3VwwlF6PbxD4YMbiEz1aiys/hUfaN6aLfKrZS75KfmrJSy+uAf6UPY4mOrQ
wc6OUBGqqXglM6AJklAMjFRSSksRMIfuJlf5vSEwVvyvg+YEZL0VrL5raKna
+K6JgAhX0dH4opi9aFD7Lx/6DO/Ub1rXXp651dERHFwmUjxnwaWIf980jO7u
T+Jzij8SpPH5AyM5ArErSBF+QExkFQekdrRtOFXopOujxS/3X7xRdAXIpU65
Ihr+Sr3IxC5T/Hz83+cedVkPrPpRFNjbOVgWslGCsRgkLG84doeD0xFkcHxx
U7wwrC8LMUAHlKI8V/1V36booUS8e1taXrSAYjZ64NrDwPTORD18XwGkuoxE
Ifvbn7WZovwpSVBdgT2eHKYr6a1E8qv9PcZVkFu7kgnfO2JMZK89WplIMc4A
rUgK4SgddszpKpcn6OOu0cmOPWAHt+z714UfeQAr+rj35WAdJOeF4MJlC7xg
WgLLuI7tTx1/55Ux3BxI4OliZw4YCCKBTnfs/FLyyXJ7FLire3Rpfq4WZ/CU
AhbIBGky5f1KuKta8mgTs6lJ8kvDh/K2eDLj7MZPHHnYN8/uFXYVHEtdaRCZ
61jrvWWkCPWyGM3LdNa3U4GgdVkQWy0XVfj9uvV3YpMpC4QOF+PBSw+NQOuJ
SSbIqK1MMAUjQ1K48o7WheX+cN1MfKWWuAatl16Nja9FDUk7jOHHFByq6cE6
6j3f5E/JoUFg2vZYIDJhZZtb5yARPUMOI5LgPU8cobqckNFB9i31Mc/xv9gl
cNZ/gAPqNsMJT08zD0ippJkNhbqqxdC6J0NMFH6KNwKytBVjMM7bkGukcpYY
1Q7u6FzH8ciy8q0+UZWneag6DG3+HExnM5CZdoysCy/nEUIG6/PYXAXD1jwU
2B0l35zvIBeWbV9sNiSyXoktaqfNiqVVp6lHCaTirUjREmxdHTkXnfsmSnhj
D+na9kHhnfuJWTZi0pY2gbxeKThrDTaZdOGWgMtqOj+tj8R5TLjcKay98Myt
aayBC6/Z+CGSFgHVaaokKZbXLXwrPAVfapGv2grD1ID4fV+5Fk1IF00/bZqR
/Wcu0L1v+oE2QJurBYDruh4Ejv33SzIGhUe4N6Lgb4kyxm9mgvQdieBsFbiR
niA7v+vEf2hb25D4QiWv9fThUYIOc66R5YpAI63Uq3uH5qiQ7vba5MYlz43j
ggloGvzGdGfbR6APUS3wJshnfw26TcDvqu46AiYvb20sJf2zPp/Xa0NUOt59
3d4ab7Rfx9IDFGga4RuqrLni2VRO398aKjUe/Rzobnf1jh3p7ilqxcGJMOvp
COFCfqx+LQdFfKAUeIyVlKVXLfvgP94KbTd19CZ2bwdvslYyQ/bKT/5KeuL4
FDvV9jzEgLvj/s9ux6tPUkJ9s5QNSvaWUg2zloEIZ2Jg6o7OHeZAEGgNlBU/
YYdvwIUot71FtaLefZNnQFR/C6ANs4xWgRMmiaVG6Bui6Bv89JT/iC0dqsdc
50roDvP2ac4JvdQBV/WRWPmvpBLjxsiOQn3x4+gkT2m1zb6OjQw1LJhtwry3
dyhS6HjDCRlYTG1/gLipv2hnfwS2LAdIwAvp7LT+N2is2r5g/gT13CPAO7LJ
b3FCgr+QD+IbqES20OZt3IKFFcG7axlHxdhbig0FSu5V+bXYkn57eyoEHqEn
FdRtd+1B3aACsUtdWOaTS1fqWshSAl/qSbpFCoDAWCYjfHptjFAox4AUWf5F
qHErS0CKU1xXkj7nQ/xjzJbtoHObMj/ApuSq2tGNhFVNOUWQBIvNigBVut9c
INhTKKLw3vM74E7fQ1kFDpIzusE4lLYZtz4hOSXLIFlIdMG64PeMsJOwFCOJ
ef0XvqyOYldLuCvrs+OTBS5Vfk9jECNsFCMHiOKVs0C4Kuel8vH/Fdt/AokD
EcCBT2kEzxdX1NEKcjLEb0KGKoKbjQO28DRO/Wb4RjdhmQapm0JJrWwz47Hl
84BH3pPqduXBHj+z0HmAFi9za8Z+YmmYvHQ0Khw9O/TP3+vEd6W6qhvDCOVr
t+TRvGB7BV3+wxk63961+TPAv/ENf7zp0tdLhnId22Chd9p3OW16NuoKxoiY
IhH1xZvCP7DcWgWt6zlKEeRPf4EHRI87e604b/0PvLTFkQEhG/x9E2wSi5Et
8tEkr7tBe/+5PcMQkw7kCE11thAJ60/SN8LxaQW95N067QTDDkH5JnJN+LC/
Rn/2JXro453xP8VSAL5gfPgVKyO+46o2CPcKIBMN8ZvdfdZPIONrLtgsotx5
CHmnGYa7WDS5CnUCtfipyW9hjKs52dcsPuJFj5H0duPo9O/WzGtmV2Ho/GLI
m44rb9dLnh+qx8BBbTmdHXdo/tNAf/8YUAAy6W8vZ20tp9jW8UInLiwuy+QU
RuzGPBVvPuH9DBOVObrYsYTAmJHArCXqoIeKC/GHt7YZ1cHh9T10s3sY2PpH
VSiz0Apb6jH/pgb1ae9dp6IHc6HVQWi2aVoCnRTGiDYozO4fNhBV3Zp+KTt3
16JfgznqgOo8TrXRHesL0EKEeiJRhdlWlhmHYfwixbkdcAUZs8nVvzl/mUAX
CztUD55PXkchaC2J9bju9GNttgP8tPKytfEsyJ8hO6Q6pMTsMgjUSvIczopz
CjGJ4V1IV6jm92OP0EuE6BWQCWe9RuEaZ0C50ibjak2hpBFQrpjNR+CA85TQ
PQmHEE4JtX+ssx3tMyRO13bdIMKxznrB6CTL5Ia09itrjNNN0rjQ73kt0WIC
s9NtHKPT+MtHihpq9a8yYhDwrGmkLfTmotjtjxB41A4f19MT49k61jcJ8UD2
WKtTXIS347l5NiqHrYhBodZM5MsxRYOmbpRLsQe/airvWsAWPnPf/aDDlsrL
9/snKMTj4EfpbkfqPQO/OrKzzkE3wJFSg/MnwewxeQlMXKbKwVpVTP9K/A6b
hdU7DDm1hiwn/xz4dFWIWAqHhokQS5MRH+vTrmiGOBzZY0iB3AzRZGTHjthi
83NJc78GjzWORf1iivjG5/6z00B79tWJQOcz2CLdGCNF4reKyVW0wzYBBzQU
FVDWSpoiTzk5xSowQljDGAauYu6eC+MNoiDgHtCjWVOqImtFCN39L3J6/0nS
xn5qJWhUd4g77y+bEIB0cD6fjljMT2vOoZTl0Cj1fFkwHRo8RjlOeqphBywL
LJZEixHHTMYY79xdlh2qyFW5euSCQjJimJhDSZuU5s97u059qrXVzEQlphWk
yix6OOMufq+akJFdzSCxMlxUCxXx24q1r6RGsTKk5kqRmPMPqDY4gnp7rc+W
yEMOPrdKPVZHk79TpQnS7En0Tp+HVpfSVo1WcVyDd7HUqpoc1TZ4aVMZ5LDC
lXuxn3vGmOLBit0plDpjbWj4dW56dWDYIrhYUVCe1aO0ezSQNdi6vE7vKsrq
bjvDCkANippb5nFRfJb4A/qjxjObdSM3PsOpInYvH3a+5i2TmDbrMCFSTdH6
KhQ+zDgMuIiWMmbinjvGZZnE1Di73XIYm/HLMmFoUcrdPE8bn31QU5TW2KG4
Z2vqS7s4ipKtYcYguey9ebzV1l8beWunspUIBtVZkHCsu+7yNeAXolnD7djT
961cVIWZTsg83bB+/SgsI7hSaeHwagv1tRuYlYFduWkUmzBFjjocQA0XWda2
m06txERXMeP21MjjVJqFVVLCQPY1975N2bjrg49z9toyMwDMFeYUk+YcLwbw
GDTt1LPXw3J72aXvG/d0+aB9czF2IlNR5bPkVT0YJRuC+331k0wMzNDutt9L
Vjv8rp23JGIXZQ5+6qHt5rZBe7JPBClC9zWSF74WFRvkAzKzWCy1Qyf/nFCM
Q7rSBVeNNizLEStcozdEect3UpshIDYMwgJQaPSbI32DBo01beo2bCR6M1JO
JqRRVeHbu/3uIzETDYxvCCM/bS3lIV+tY/s7pOuc01D5FXpsWch7czz4rM4Y
jzXmicOB8Wth/GDGcw9PXxVqrJBp74fJsWoXsuZWM+pEKffDBmXaAzjA3fEL
36w5Yo5t8MmTbBkkWQXEj8RQuezXTFpwBMbkh+uHZzXK2TzDvOOF01T9Y6rz
Mr2it080TxmH9crSaBBTLN1wdNTZGe9DrDDyXcu/KF+uFjVaG/rjSf3yWE6m
G2+Tz/KaKn+wS1CxAWet84JKD2q2UiFWHrNWrQ+b0eGGjIetJr73hwxwZKY9
7ziZffT5tG0d7NutkfVzDXLU3YJrqQd6t2/5yy3E2jd/wei9GSq0Kj+4dElV
iY5H5B33biu2sLlaYZuyydLG3R1IOlM0gTrahN3nXBEemtbXflRVZk+DahlW
pCbYpBLxb3D48t2JLa1UPnq77BBp7P+Qj23hNCHtYBnflZD3ZPBHGcKp7HdM
m+lL5LgpRSgDySRyPbuVUyu3Bc4cr9gGj7HmUgLSNOE/tsU3K1CYpc5lFVvM
CY469Y1RcVj14qQUcAGm21XPnZSnn3d032E0WwjUniMiij9z2+Fkb2Gape2d
xQkys0etRSrxlQ6lDltovfHQvUGBHUxmDxgFGa9pNM65ZZfjK4km3Ntcghrk
vo298TVVSHkOamnfMiUQA3v17RZH/LEZ8ELmihFeFygVzjy7C+aYlra6TRMy
n64Z3zkUBykNRwXWeUPHKFEoMayDmY9zTtfkB7WyyA3NDEVhFDX2mVe4V1kY
dT8kkLzeQ+5V33q33eZYz6F1EhqHgXYhkK549s8lcKb/RBMAOqzAcr/fLf6R
CNr65+PL1WmxrqKjTEqdzjxv6CfLsSac0oLjsWQm71kr5DYzVXn2Wts0LZeH
Dhv+H0WsLWr5pizR8r74BTi2WI6tGg2htgIJQ/e7hbvwB+8GI5OF+faklGR7
Ii5xBZri2HiOx6xDGNmQRyIaYuQBm4yvPe6n6tzjSHq3ZSzrWnUJrWhfU/zl
U+Qi+7jBc7T3jYf7stT+fi6YnFMrQWyCn4dHUfEg/5seANl1F7AJ4DCkuVBg
sBLgUhVAEh2kFE1t4ShpozvREYiRINZXpYDb5/ekYHl4LIso6u9/eTy5yHZo
nXUJPK3glxudXRlJUEhcxsbPM+znUXrvX5qlvybB0mUN+onoXZ8WYsFK6hR1
Mk298QXnwdP8O8J368Vz0LoFtlpbr3qSqoscQL3MC5kIgcsTVfRfJvw2wgmX
UGpJPxA4JcGuZHnESZxnTvNiYhqRTCzJMR+fimKZ9LtoJpRCimmPnHV1mkJc
GVtrZwOw3Z72//IdgMdhTWJk3AJwLhAxMC5p6h2N2Ic9LWDbayt8XudJFyJq
xOQerDozRly4AvCbFwVGQCYsTFnr5isuzwt48XlyOzYIZcVeSi8uWPL/R166
C0qeq9M6wch5IIR2akhErOQmSP3cE805h2rlnvPuOxerzHqcQAGoCL00sFy9
GSBaDbTSV4W9C65O5Rj3Esf46shCvb3lDSIPpJQJ5uSstXYIYTGVlL40R55O
TgACdW9CxjA2nP4LtHdq2i378TZQGp1KkNffMtz4vIRupQVzdmbW3FU1e0r5
w+gzdGUoM+udD44rUOp3PxQx+J3tgHfuS/sUZrtSOZSI5NAQmIo+VMyk/T0g
BQmOSdgccJfv7uc6XFUMEei+8sPPPsP30XUrYcl/YoMAVy7wYHvJCEWtpWpx
DfoLTwCdu8gObzyxa8vPJhhOUMqI7AKFkt8XmYfxI6UxJkhkKWngiZpnRkec
aOIs+atOSuvt9kMX9AGIuDpkckEMuPEbhmPOaezgNU6UmCn6fb34qHy4TkOt
OdQsztS4QWgHR+NcVEkJJ5rWY8zlKEXveXx1XSnMyrRgU8cUz42JYz0zsCBH
m4MLZkf5EBMC3p1VuOv0QqQFfTr4x9DLDOF19UxcTq6bGrX9VQm8pY9Z6cF4
1time3yywovnkVyB7y+xnGoKQaBcgFKw8LXhmRxwA+4L0RE2Sd0luuTBb7LD
rV/4xyLC4EPlKJu3T7RzJayPcPDPzUQ4cFzWKDulTVXmlczeLjyWKiuSRCdh
PAuErOKAUm0pFW/b2+Oafs9Stl+HKh3oWJitKbNwyDV3X64Q9rLpGp6OIyVM
Hd0k7GWGABS51ZQgTfzSfrSYHhVSiaVr1xIRHidCMTWwnJZLrVJOR26L2oZv
xscq0NCjEuDyAiMKnwIxk5Ul66EtUPlKFWny8p8o/d9HwRDNPuVe28EPJJFp
pDfpv72DRJ7+Si3bHBPaIlV7mylT6FZSfZdYYkQ0hZH52J9Yr1yOQn7b1sVR
aoTQwGpeEn1wsiCkojbQKmPcScDnjCSB0gK9/ycE1Oj0kGKfMt3LC+dZkEnF
EyMAsrvYv9khW0UFCKQn+Piw4VTJx3iATGqy0K0vHa7uAcjTTfmyASesKbjc
vOMWeR2uUc+r0KGKcrKm+9tFQZRr1eA5yiI7srtMT3KdDbUzonleLybw/Cl2
A837ImCs2EF96kd+kHxwQMyqFJ7lYPSAONVc91C1zDT1F8hSKkMjgYXc6R2w
N1ix61jbdGiku5IVLSnHBmssZr1oH0OXQlluz3eH2xigRCPRiBxmTzWQ3lUC
XYzuWYb21QCbAZP+WfidukQDsxsxex/KjFeWA9TCkjKP6aYxfSq/czJHfz2F
eUi2uolIOUCv2q2n+68TtZtojusjA/k0o1/BbvbunJmsEjEusCyYBNHghho+
XnVxDZjyudsxFS6IamuO1Z6USnUTklirZJR2v12oJKhpU+ytYe968nXft93g
8MCHisr66LoZrIjGUJpCfRW9Y2Acap8EeFgooatko837KBO8WINv/SJTAmDO
TKcaqbsXmXVqXm3FIJoqZO068Dtt1uKk3ipsGOC9vWRlrb6BGkaSFPnP/63F
NJv36bbTJm//QCJQF3GtSQJN9CASzuONY6kJpqmzs59VChIQDiChv8fHoNlD
fGn/qJ18Bg8C64BiQKdWlJkfu4ZwKOMTvuvU7RoMmiSN6nIfotvAHCr24MfL
y9qI5sIuFdHvG67OJU2sl0co2FglnQGPfZeV+Q4+iQJw4cibklf+bQq/a4ym
yyYnVx3Wz0vxrtZu8/iQbQdVJptsS5uEPM+1uQzXgJXnnFFMt3uVek1OtBlY
nmRCgh+QnaMjvLkS2Ig8TOMzECIhZa5WMOYzpb3nOOH6/EJWzkzFBsFGrj0G
6fNX3tY1mjXpldKB8bo8h5C6xw2iHrOhmIvN2YJcwElUnBJPJfiRyeVS2tW2
XNAZqvOd/KhngEVx/Z4+yzDVpm6TIqTq3mmqZnLT2UJusQnmVvui3gBC5Oxj
vLIkruRtS0MFiIqbrzwyDYEg1hJt3MyuIAfu8iUoYDtL59QRDAKZXH82kXy7
gobIdeUYURJgXROjkgV+h9rpjwhYkGkHsixYZUySDJql91r1VMtIaK5MQI4O
LqiqxM2Oo5pdSlrCW9KEp8sEGJW3Mq63cNN7kcoFF2+hO/3nfF2p1io4reqF
vBvyTFditFK9N8LiTfXMYa1C/FTmgB3pkLsdTooFNDzyF24UMfgPWFYHVjNk
K47Sv13FV//+CqPr8rshJmBl5TDKjCPSofgpHbCL7ltMRYTP2YKOl9cH4+EG
EHcg8VL7U0L+nXG9KMUdrgpGfTInwWsmIx8DWX+e89zXSdbtmnYPvSMQFxsr
ZOAGjwTzvJkZjMfQq0yJRLIaRuCbH+rdfCAmvEIeopxCO6bDo3A9qivrxF4F
tfJkXMwdHzLVPbVX4XV0wj1l+TITnSg/pr6xSZM/MZKZY0bHdGxks0invNwI
htN5uhupPXGocvvV3kE8bQsyV4kxpt7S0vZp/hCBMqhtacW5CMPWP20bwdDk
tJax9bOc4FUw8zeHs/aYyp9XEb/U0Nkd6GWN95n2BPoZQksluTW4JoZ2naoT
lPw43QP6dFZj5rQReYjFEtvSuSm7/ovqr8aVz2gL5lQgnsSMgq10e/mzbnfD
oF39I8Z3K843BgRFRXdKNSonVDuM2kIlmpC13uX4YdP+P+RLYn55aspA2VBu
TFfKRgjHCwPfv7/WJsC/9kO7yohzGmFfAg6YfGuSmpb0GM6nZQXCM0MvlJvq
oz78140HmNtaMuiARUX7MZogrvyRYJbeQeDr4p6sfyhKzpobfAuqbaOiHmP1
/dt7O0mKDeKDFJ1NnU7ta/Y35NcTr5u+aYxEsk4GcmrVMszlTZZHZVFkh+1n
vD2y26i8k3ZOjJExFJaEvSleJJr9uvO8kvv95qbrydx4hASL5Aye9GXsLhcm
fLTrSb6qIXD2H9LJ+aPFHWwif6wIWAEOxOgyoHZUw+VRbSJg0n1bydImI+bo
/RoLKieKiSVo9Mush013zKataa9tC3kVR2njL5KiWDF99UQda+iseWy/H5bv
MRP1RzobBHjcjaoNzXeS+LMM0vS9yjPebkW+Qxb8U7NbQHYX1xEDWVkMy8M6
G/VPgXoqgsryMr2B+uuHxZpFp4bD0hFJTA+lrdGKZ79t5OEG7iT+X0Kslpsc
FaFi78RagSr3u5iB2rZDTLVVat3+oapSZwpFAKjVzn1urKHXJaSMueVh0b+L
bdNfS0U1eJl+pnKC491D3MOGKLsLoT0YQcsi3983jii2DeYu27thaIVDbjAY
0vIfVoATaqbYwDHH20Pxhyukug+Kg2GCTHtgn1mGZZdB2L0iZPczBdYnjvtx
oENHt/5ongBjREejRGjU30XsghhHOHdijhPCxoLTIiyncoBHH9Gilu8+COsc
Dah10vZ/Rq/0opba1JJexmGmutgdG6SWPV6dquCnPjsXV2w3/TCWLb+3D5ne
Cubq6yYwmqvg9a8vE+nAcyN2j6Dg+uOP+OZo9K0n0XZQ2Jc5ah0uenRc1knq
a8NMrXA/KSzV34Is3vMB6CVIQeYvo9H4AGUlAn2Sw1iNSNMdpjDNpMpv1RZH
ruMwdBBgJK5JoZS70KL5g7KvlwAQFXnifuoMD9p2/MoZHhvWy/IzpJBMKOP8
giUlsopuaQC6Rm6OMYNSWRk9RO/PGAE/eNTCba9h2uKBChaLjWI/rqAMEyJm
jHt+fBbjBgiuCSo+G13DRXmBdl2FpYVzpz9XHHlRdnUt/rg++nmDMjSsGzeR
rWuPVKV5gts7JMW2or9jgcbwJHZt7vZtn37kDzFoRyMiENPbUbHszdcbxfzc
LdIT24gcI+uuqkehwq+w2e+oneau++vF9tAy0x2o/gSisPc9C5ezcI1XzSvL
sbI0nzPj4vA9QoE9TAykMQpo18dIY39KuHoZHAin8za9yievvhYGYjaBWr4+
jHF/J5haEQfYiHqPSG23b14DmSyG/72CJQJEDLC6ADEuHvSbe8AeHII9YAN0
PbyI6SacW6OH28z1P59FBPCi3vdhqtsw1P66ppmXzaNBqJjot99H2cGdxCIN
RVKDy4XRJhznoZuhtuQefxF1ul0YBk+IdW1ZP6vqRwIzhAOtBGTGAvekr1F4
qCK0KOsrH0YU2oFjBlmYJICyHTbJ8syNEw6jP4xOFTOpI24pLz4fCjp1VSgV
pWi3BwVN+m6qSZxvkCf1jTKiWHPrwD5aCzmsbAk2QMuNmEhqk0mhzgwL/YpP
ILTKUYOVWtM5yBp3R76/6ILLqekDn7sC08de/uQJQKFkA0lLl7MWeJ26RXAq
1wyncruA9SDLK13+R0h0zq20onEV64Wv17KWeaAXybsI/dmMcpULCLz5KVG7
AgbHhOJkT/OTekN2+jhDNGp93WWjaQ4dQIdfPslvYjgQn0NR1OHrIbj3cUZ1
wpd/FQknH90yLX9xKjh3z95KNpKKf279kBNWeNasY444ylb1296/d/QllnrY
e1Zhs0GFsiaI4EniyNfiVcVUcF8qEC7Y7vcyCUWFUw0N9k8Xx0SOmZDLnttM
duurXvKF0HEybkbbndT426Se3R46b24ypJuWwnpv/cwqIDy95mkiP8jd/LXw
IpNkpLnYL/fGKFu7SudD2n47s7IDwOxr9Wc+L+pKW6VXZZH2LkpNsPqYSTOi
t8DY43Oc0GfHoQOswnCwPqWYZZhwszl5yRCfJwcKXDZQxT2TvntVs12rovDd
PdNzASZDFqN2kYQqUiOZHYLf5NquSu9m2tqA+kj8OKuN+9BftF+exnXavzzg
oTD2UjwTTGcx8EK+0nc3GooKtyc0q2Wugw5oyNkm5vk9QUeMncGQKLFT6RP7
t+VsvLgHgfFb2GYAJy1lBIjYpoZmOwbg375XqE8RsThqItzVzaeG9V7cYEXS
AXuzqopNCvo+1+0XDd+N+GkuzSakvouHD7rDHzckPU7I+rcZ/OmWdfWCasmg
ZB96JEr42EHOtDT0dAxQJhlD8D//M6B+8i+KYAXSlnws8CVSCwVrt+iUIv+i
28ZsU2m2JeTdQCSILcyH4dt4W+jIuDSZjLHfO0mEHAtQPzsNNDX0Z9jzqgiR
YjuRrFfeIkHlDeIhTtEpn9dH4kX0l1CGS3VoZEUYO0p4znAKZ69KY2tMzKNl
2t7Mh+4FfNEFjwfB/k0BEVS7oZwEptWvzEEYvseCxB2ub2282GkaXVAQt3b5
EMx7jkzi61CJ4arOCFXcugTikWnabZktHEJFwtBKQuwUSqU8/FqoFLofa2PR
mVs0+s7e1orjM1e++0KNKJyDRpIhKlXaT/4tensD3cieeO2ySOsvN8VqVm9L
XPhoLxWW9syWFEcfe2yLBS87fQNwlvEa6TSlO7ZS1onYGf6K2M7A+Zegpa/o
fX28Mq7ulUuAp/p86bIwKsojBwzKYcOfjOD/lkzVJlx+pupG8702UOz1ti4H
0TJ/DGEMMrkb8AI/JVITzsoCP2o+q/PD6UVNN0w4pM0yDyUe0Qv9YCp4TMp+
ew1lOZbWiD41VtkJVZ8+7pwGpwtYFaRUejawen9cE3GcRHow1QjyIqQfsMh4
auvrITq8ntiWtHKd/OLtAVkTWnSkymFx4LVU+7FOvffIhQC4dCxndmGfZSol
UlchKI1RK4/e+Va7JiMXEU8DvhwBDCX2Yep5HHTMDFU3CGQFqHhvgHYVr0VF
4KUhJ2MpqvM+7XfMa1YR0PW3Z/ZY8GMszEF1nSt0GoS1h1yLYL4YF95APTiH
aXgfuz2YEPkYcLFOgvG6WI0Yca/c9MJgsS08iDXFffNsakajS+9BFoKKatnQ
cOxxAtUy5Wn8Wdq2XC0GNfQK8f3cIex73BGYpkBUpdNfqtNLp4xfFw3vEZJS
EJDcSppQ6XAqlWT0VxpeNv/WqSWAzebj/mihxZTfB9bXmIFTTPUXoeFL1cjr
aoOWAXe5k2wichvcv7Xg6YeT2L0oAYXlZLNP62LvOurHO7C5i+VWDdsZLt0d
bAeZPdrXxk4gOf1SZECIPwM3feqT9C7qYo/jmw+nSE0gx1m2F09JkjtPgJDv
KpV06krVNzjZMqc+PS36Z/0lZ/YYtju1JIGRZHDgfoRHmTTQiSgrphvg29b2
7yM8hpMKqG0sjz6syZfgaXKL1bQpyzwBX88X8dRlhbczQVSatl5nhvhIu8PU
bAOmNdkJE3py1T86cQn9zIrjJ4FSpbkKh+tL+aZg3NCqUJN+G7twKvpErMXL
PtgsvK4qv8f7A3Wtlq2gpLJinnOLGxQN93hvSQqp5AlMfhE3xfNJjWyOl7fS
lQFQKn8vtqtkVEeAG+oJWmZtaez6lJCSsdKISyJER9lm3i3SnJdtD14Vt9LK
/yt000m2lRjyQpNINC+kedlRQ2IzkBpEUETgXrmd1VjKhyA1FMvv/WgtfLtg
0BmQnvlGXGsHqq+7QTqn7PPD53ZwznnRUxmRpfVUdarCDzwXGSbaa16bBsNE
4aRrFPtMG70Rt5TBh/E+T7sNh65HnTT23yKwugrVQRNbgss5oYNahGArQEcl
HelZliIlC98IXnIPOPK3r5oKEsQ/khtxpuIKJ51dP03lFy2asl6tZ48elHGO
1Pm5VoM95GJxoaHdXEF9aCKF3tvv3qlYnPsid1gEMJqXXU7hwL5J5sPUkx05
r9cOiukxXaNPMUT2K1qOKq/XaDiD6BPusfj7MnuE5DZE1PkapadHw3uVy6UK
W26/VbhdBOY3csgFUnD+2vbHTvkMqMsAGTvSV+zqs5ZOKe3RnJ9GwvCwaPxt
KUPGoYSLXsIM5Uh83FbNJRh6dxAHh5fSkKKzvi8VRciMv/h700Iz/4TTm/Io
0S+Tx2y5FEryKJa8P5lknWVqzgSfOLcksTcVr1H9wXo9H5FqCiLAijuB/JVi
7sLWJyeFKWdpO7DKDA2PTaI2k70yaPGXgm39wlQrHLqYZNDLMM/B4JDGf9RK
Pab8/iGAIEZb6wGqFrbEksWpVvZT6/VXG19KbYM9F+9+DuzGheH3icAoxCAK
TQXrVbdfkKuZmc60X7hxPxDuIsGzb8pzrAaMo+foQyVCc+X6oGvLQepfS/DC
Sa8kaWHJ+vhf4a5nRpMG+q36CIM0gB5StI2crRSgjAqNrMfmVHcHE/OZAJbU
NgwQbIgBuoii5KDRX7BRqfHfjh5wQ5JpBQK+1pBxfHcFzm5BPA/RmhfCYcsU
HNWaeYaCqkovxE224TMaHctuPxlhVKZcesF+PvrKCvIcDzgBkao6eqsYBblk
uBjY3cj/Mfi9eZXP9i+fWebWE4ou0Uc+s21w8Esn/CqFJRIoGJBDSsWvE3JI
qzi+UmB8fcFtrgMkPk5X/tFsn8AzGB9OPnx1fEJPzQmafc9oUYsbPgmWFt1S
kndQshJLvaNPn5Cq5Y1+sECJwMy1GFJifyTd2waDH15Ysu3UisPaq6hvuwQL
QTYjMoYV/yTyyEcf3gK/63Lt7QY+arXzAlMTnLJZqZLR8V2pcdOpvq84LEoA
agLdnUK+Ve369cVaNyNfY0IB1VdlfJAnu/eZd+C8pT0dVq+Vw4AEuTIUGV1Z
KjnaDNXpkZub9GSNZB5ql5zazeU0r9q3R3NwFurAx1wTLO2rJLLgcFzcuHeo
r3cjI/YmbfvBacYcwsb/4IA8XBeZlYDTZubIrJEAxX7lIQ9FXLrLJii4CXjZ
NJDwktT+3En4SlZEuiwhZmrwJuZtXMsQKvAgZ7/3SlZealz8upaCXFl/yZxU
vom+OlRqzYiRWp+jNTt8vnpyQH/51PNpyjQhdc9ggGaUCY9kq76ck1KCZrIm
4G46wgNBj5UMUDH1mdK0oGjLH1YkYimxPPJV8cF9I0ItZsivBcIsEBfLzUCt
UrDe6xkqB/2UtC299Qr4tQrmWI7IinouYtKL5peRVRAADja3M2k6kZPBsXYU
A8yYp6uC4L38WrkrD6ZKKSQIVrkM6O5CYqhOF509mV9rCZYiUhlmnfxmuYXi
rUki1ar6AxngzpvSTMks98sPIDVRUZseHsIz8f4c0+WxUDuPFJh+k92SsVMD
k3gVyrAmsfx0P09zGWpsFFoJ6aQuIL2qqLQwSRynvDLQbKsxM7YbqXxB3VF/
lvwcYkdG1K2y8DPWBsurkU/t5BAMGGLQE/WA55QpdoXycNDUIhcty9YRVKK5
qidA8SQFZkTjPWz52czO0bnhFeOhB54rXtGK9f7XNDlJ8wWLb31hVU4eHuxH
MXK4GIWoh17EgC/hyXuid5Z4cJ8XHbKKGz2gzkICcvVNGuX6q8hATJWwDLKt
c10PBPEMxM0sgTpwF+AKyVHZjkQy4hkogfyd/VgIDDr4hPo2CBoc6Ve9HdIG
ln3nRTPDcIDtcN7lcDaTsNc/XwaYkTj1RSbjEsz0mrmcDgph7/1QYmB3+T++
0EGY7oTjIsLwRNqKhkiT5IhwxJzmv/IoTEqMGl7QzZK0zBUIWsu905yC55ro
GKC9Jk8qZuIf4ScL1BCE7KobLiA6HVX7o8cUUE9OSt+LDvKXoNZR6x9aFCMK
frVNc1SXVreVvC47ghD5DAbwULp4Cl654rQ4nniGAzDGifkMw0zq1lK6dqoM
MKaMNXhNFe0hQkybFofuElCXjMK3bH4tR6MHTD4mjCUX5rvjHH7fJJXJOy2O
W2mAFZCDicUzdA/bkydFoZALIVx75dT+VDwcoofX4mRSCHMlNiRE5RrY1yNx
wzH2pKXQpYB8hMfICzCNIAwMEQItXqjVfzK1JmoloRmzVL/4j8FkGoLig07X
caOOO4bnOpQIf6dnydwRuQPtDU2c6IeJ+lIPSZFTpWuFTmvnHpXuL1uMputq
+GqIv0WgVMDHHGDku5cN3v7bQrAULRs5rrPG5Bi0L0PrugRDKe3G9a3uM+pw
0I60+5I0wdUzWSdI79sYtJ0ivGwvybOJyHgWadtXMJVDT2y+CkasSPrre15i
xkSowD0dsrfu0I1GbQFUdDzIcgveV+k5baRDzDthmlJPd9o1X/+cS892ccEX
kjHev61vGO2uFWrSM3k9fMBpVIwg9l0f8oZWIg11OXc9U0OIrjRQDM1FRrFM
DeIHaM/GGTaXtmQQYMm+ThHPSx3syQ2/QgznQeGE8QfuAdHYZYKxyd3UpBqq
/mwgsZn//1ETNJoBMcYthmsG0oOfpxO1CKlSQLpomKb5XQN41pwAsOp9rJsE
WdJa59xS5hdXoMaBFQFADWl2VxmdaLX132Nxg81k8xpJP+qrKBBEgZA8Z5Gs
UeBak1hna2Rm7gztjEMKQn40Msrf+yYeloaZ7clz8B2Y3ZJgwDrWYMeRFF/i
v+Fzq78b6aBU/B6Jy0II3qz+hFZoV1iDajusdowMv44G76/tavZ4f446Trbe
G+MZIJbqz/pBLBuwOURY63NhpQ6JHUZT+npjiQGGLZ+7N97oHFFAS38ovWFy
Fz2SWUGKnpezLZuaEKQA2nlKdP1O/pqU9oHm1uGxVIb74EH8FmB1IB4NII5R
vJe6R+M1OlrFWW92apcVW06PIsb2W58kd3nUnmVRAKCZ6f7DubScHuW7Y9gC
M6CVSC4jFB8g60VbUkIIJShlfDtdcunbhLmCY/3T9I9H5hijtN7gqcV/aDrb
rjGmpg0k6M76buEv6ULAYWw2ON5hPKDvKzcecWMIJzOq3MJqHkwubN6XzZac
17gYSf90P+FJLmbcvGvuWgqZqWZXsAf5GqBcq4Z4E/2BWG3fHKMnW+sMV7SB
1f4Y95/UZcCTDf5P5KJPX6KyvazDBmTLlmWsQzLL/1sXRfaMW+l63rH4PAXR
qy0kQEy8WrCUaaWJAzyt6hEqhS/ZfBxL2lsBeIblI8xbnXND913f+cXFEwyQ
q9vB0ycemDQ8rDmlss56BI/zaIC9MK9P295B+CmGr7K06cxLi2ivmcxmkK4P
dMfbP2Zw92FbUg1mqf3CLrtbTTZhOhaU/jm7Uazlrp+6XrJp4d2RJ5J//qGc
wIgHQJb20oorMZf/pFw5stLfjTvx7NJ0loWpBwyXSoDRI0O0I9GYWS5Yrd8Z
UAzjdW5GOh/03RoSXsDnkVVcFitc9CGLpPMwKkEqDPzsUp6Pk4luJMbxBSLX
N36wKZvuD97evY9CxCb6nKrLOyQwrHw3+iOkYinW535gETlx3MrKYFLSuexa
lGPcd0rHzoKt5X9bwMDpG5qy8DpOmRDoy441Ln+6bkc+NU+qiZ3pQ1jeuloM
kZw9Rpvooc9F8LSmplA1hMH4MMR7X9xKZBQ0KPG0K3LpIoCe4m9nOm6/F3lM
PvOcWplzvZbcXI/d8wUm4Qgqs560e7R3azXNORwexpf0uQjz/vsLntU3+LUr
4ADb6o9zP8fbqWSkG8KocDBVp/u8bfqZIKiLhUPN0sfwhezgr2pKv7HElSpv
NE0xe3OBYMahCkHSxM0BMF8NwC5v9vzce5FPhMHpdFMpmIh1g7TF1KFXtb4f
x+1mf46YDJC4QstZiDrSEwP5tD3qL7EqKiEvOjNuXJ8/Wo51w7dN93FUJfuj
vUkGD2efyasNnQfmflLogRSDzYfDwO7spputy+bOhPLSg0l32KfI0+rBQAnC
zuuysMKknNxKO8cP0rIELqL8K+ZwI+t0x8qBwZFMIG7jnG+pYVO4w0gwgD+5
sanPix4zWP+hsGM3y8UfQDFIF1AhszD7Ob5swwYadlLOTHx0USxOyp2vzpIF
9T5Fvyrz7/a5Q9XA08WmaUY6NVq9aMDNIMhBpVGsOINaSCpp/+xiaEmppBmf
ruMsBbpjWSPghXToGVFynHGsiMkXgstJYmIhffzgvm0K5f7kJxuMvDTXdXvH
OZ5cgMGUjs8O4swysnHqmdEpThauoDy80HX3qVu3P0YlxfBQ9jWFAFYo1uC2
uOSpHmwq3j0iyJ4Xs8gotlElvD8umeXaG7X/ZyRKx6JS1R+emj/wzsaarn94
SAfN9m8E+pXb2lGMHFUn+o2mBJK2kX2n76VqByx6Ww1FoW2hM3j3xGjPZc0N
d7cQ3ztT+RNB/7YDoHcCzlrtX/tJaMlxOUunL2xeLUOMez9ZeaqGDbUCLaNx
LRUtvMcKRHLk+FTGQl1AuNrWXDoytcZaUuAUljv2HR+QsYcHBnFfAC9TYO5V
hiJ7/nype+INpR5sACZI6qF6Eu7RTDDx7ULIOXxaQdJ9XIn5jPthdJq7mBEZ
f2rOnvCT4LvXoH0KzXGh9IJ9mJmEK1pHPriFdBG9FMQG28zA1bp2cY51nUQ5
EHoLpazyj6ORFgTZCuXc60L36+GUt9svX2EPQPwO8BAiFzLRK7YlLt4UlET2
znD+ShjHN1uMcz4rTY/iHRUVs0VSiIVoMDAsjrJnQYqzLBIk7IyK2u0wJWkg
kMw4uHdCAY2Ck3nfUy1K6kAA/FiVXWVurTaBhf8lTIOJLX8E0GNdgdoTBp78
pP5bnIf45/SiuONuVWA2YxZov83jKNLT1us6WgW221l4OjTWV5w+o7jfLXb/
sVdwrJChW2Suv1YanpEj2mtGL2wkLMqr3FMj6ACFRzDMA21+9OGc7T4krQMf
C3sHVUIvQI4rCchNZ/lhAb0aE4DzCTDAZwiZ0uOEWNTNTrFj0mAZzPIv1Ccc
gY6T7Nk5ci5v1UotVsOLYcQeV99bBHNikxW2CXHBSF9QCs1iqvm09RadGieU
QxtUn97tyRlck3iRX+Dm+5rTzN55MC9Jr761LuVv1zRgmCuz7J13PhtXtfJc
vCTNQvLDNTzibg/MfY2KQuHkTgQN4+HM93myjIWdOFIkKe1yyIb2kdYGGLkn
N5PpUMY/Jn31FAOsIf9yo3ScSpoOO17Hmlz55dtxRuR42Tglvt5Mq6DA9ZUc
wNxt6BWHMpPqG5n2XZ3iTTzTF7F9JjRlfHcwZ0T5x/Q4tF1RFXNcc/i7IgOB
vWya3h+W7RSCH6mYEM1qCmdiGZoz+H3Wz7VNCi4JbMzbRDFbPPas40PvMQwY
yOvNnPchlwQ4guM6MYnJHMMkrFVbarXBOM/v/nLjEv/IpI72dWdmdlxXm1hh
S3xJeNJt6ZBqothNI2pXy2eXiItFZDDnXguRetYIHD8R6E5LzlzCpXCxHcBn
GUKhEV5TF2ER1uszmh6RRqBEeAc4K5devEtUN36ZO+ZBKCLzCREVA/tdOcx2
k/sQyLsxl48LZRpzuqTaeWd0uk2CeqjzmaDiMnErX/RycOp8L4WZTt6BjIMQ
U4DcI7CiqQAao99VciZo6zm9xWYqUSQ8zqQ0/7VqdJZ+CaeqZEKOOHt1mQHN
+D4hj64R/vv/5WGLCUtOMKXC16CLoap68g+co4magjbRivN3DuoAFMCqvlSI
S3G61Sbvk4GAmRnEVRyaht5R1KO9L/7L7ElTagMrh9zIa52+xi5k/QFux14q
QCeWff+UaMzgXGvTv3NB7aTic6qHqUFBZN4MbyDpE2Fu0P5b/qTcX67jQda8
8LF/mwpeP6R9GLfGz8qchGbV5s/m1xgQFSnUq5sQ9Jx6vgpuuJsacGQX5fy3
12yYRKTn+Yzb/ziv3zPiYlUTZec22aEHoy3PPSLN2ofqG0ZF3uMTvat/IHAv
OLi7Ly+qMdvaQAindQrFPBr8s0x9IJBW4Q72dhGjAJq19zHnGMpw4+8SyKXp
zeQJ5LsFWQH/NmG9CFIIXsGnCZ46oxXmJkK5rVrF1F/WCLxitKM6LTRy2FdJ
OGRCluFfGH70z0fQ54gaGDoWPxLbFdg7CoyGEZ0ArS1NahWUgfelyBgIxPtQ
Wh/3Op9djz58V6F2UNxnYCDVAxLGr55zIFUG+l3/ZwQzvhtvVsEhKN9psH7B
1Ghciuu60fekFzcCmObNw0i3YqFYoKAWKHixm5VaxhHfxSfyz8NBHRmIGTHK
pD7/YrG9sh266EPGZmBZozjiMWnQEQ46jR5daIx8YfcVTmlXtkeJDXexuT2Y
ive+EM+3bCvl5QwKB5EBLDzEoHIogEX/FY5vp0lxDqD+hMa43rSFv94fQGpM
biaFmj4pwOE1NWA0jXnzeiB1Qv06IItUDPyjjxJDc0775zz5sahRMzTNCoCU
Xqu65/jGl9biibxXr7hWPWwOJwsYnnDMGfMbtmLfEXLOyIOwTrFZ1U3hmxIO
CfpQWht4H7Nobm6BpaJJ2snbuwF5VoMzSX748BNYBW2HfO5pPVkpOM8Cn7qM
zsvajZMCPM7bsy6gBzdktnvbnO9AbVTjab2iIYMiqfmRyPmfPC9b6HJnPBtF
G9jIY8hyFTqJ2JlWhxEecMTM3ADxsIsHF9PJSYq1lme+fqJSlX9IIvi9KoE3
CyHwLwyWCVFqz0IQ15a1clDTFMU04M2pkDGsXTOLSmE5T9GLJ026OegVlcee
RK7hj6tWNmcs2ztwBfzpSguCo3aqsuyiHm+6M9/jeh55yZhTqd6UGpmdrHFd
SXV3IgYq+orbk+XHmOAO88MRK1SgGYRyrvH2A12l3TmElfqLkk9BS0vI5Vx9
jGarDSClduQIut2BXnjQsVoY/Q404hekugZ+Gcewx+umi/LNf81Jrgi1MvwI
Z8H53bIi9Y16jikowrshT3wwd+uxMvEXyroNfCIQxiIlGIoZNGxWF56BQ8jH
Y5M7tDv2y/A5pX7nR2QhImKBGbOdZkiU9Vx53CIyU8ubktJMkJVhoKe+R3Rs
tJcC/+qlclwKwbWUzaQ2qmvxhVizxnFiK1vGpCdSOxssSfzAl5e/Wqr3C+LY
sgxez4t2oaxXDMOF+ZWAItuSJzo09bJdPPuOkzpV99386amicvrFVkd97YUE
BAgXD7UcM+D+OUhWNwXqMOLFI+7r6V+cf98fCYdSTRJONbK9FqB4Je36eYf0
r92FwgL4YQXMvgsJNzM8D8FTplgEebRF1G7DZqbzjAHeSqAgig3oyvkjQoJI
w/ETTM7NoNn4vMiYfC7h0vuvsuiO7ILHanCouhboNmJhQfCnBl5tu8nxGXij
kBVSqocNAqE+zLswZiBPPlECOOddoW4hjeqJw3OLr4MndVymbPYqq/aWnEnG
OeWKXR7VFWI/YIHJwsvlbE/1QduivNMYCExTzMkmJckaTgTFkgttrojCKs35
7yVxppPa7tGjHIdF20EnvIcBsa4Cix9gskYQ8zZU7kDp221IC+dZHf6BnzEI
pVrkNiHMAbUmhsiVTmF1DsYAoKiZAw2a1b0Fk7QOblMWwq1/OTjiL+SgyNXm
LBbfJnZ/7VGVCQi+IOg3VHOsAYaQb2KYyEjjYw9WR1UbKi/MUBx38wDALvh/
svuHQS5C78OFOdXHGBMl8tu7trg1kL6jHSOFCUvLWomltmB1TjWsWrOTmJrR
ZLYFDVjsd4fIh9fyqtwq5Vd7Bf6YzS6exSm8dQ6bkfMbrx3b5RWEiQw6T4aS
COnhQzCTYgFismtP1pNGDmlZkG2p58v8XWYVVIwj3OeaCme55NUOYXTRVgFE
ojHYMpJ60kjx1h2cvGWnHeOZMSlbUmuBAAoQ5b9f5HL51eue3tgs5+vo0NRj
ZuLkxnc3JpUsKG9sTg1RetsLkgyRov5GCbSDk/xykoM4CZCimtu9CscW81B1
S7mM04VFYUmqBL8WsytFzwYX9IPhJHlqGQyh/wgY2eYDXNiayvXdfCJxslTo
AChe1G4n682jhUF2FOSokr3HXBsqfaXYc8H6G+G+4OpCA3eijH9o/LBiVqYr
vMrij6yoGbOwSR0sx7ChlKa80NfCy9OnIkC2wxdiemyx/6bqseCFgOZFE6vM
hQn3AMUJKbPKtmjJC1l2kkBuIT20L3O9pXU32tFSvWRJlScviNmt5X07rGwp
D2Ub3tTumybaUDcnIoADrV5zDyhTFEB5FFEp37qD5Z6TWaXeFsWCjYQKfzrZ
v7VTdseWjgJAKgBxHVFj6WWmUj+lfWm6wJXjTFGjxJO21MZKSSj9DzCMo+DK
KMjXQUSiNN3eQNtxyXriAQibQ2Vbxqgq4WvjwYJpox1gRfTwA+IJJasarlrO
/mbasP1fmaND2kcK0dDU/6691ueKf1aMNAjhWp2+OeklWnKCo5aVwXHOEX8d
Bn9DlJMZM7XJnZjHzlfYoIXx1vyMj9GuS3STkU8zoRc1Xsv407JcAPKS6V9G
Z/SO91wnp0ACcsj9nRfdxVp2QF1cSbkwcy6r5MJ2K8ZAfvNWRwJHZn6ocY1o
DzPyJG6pM8WApGRukzl2NeVFxG/n5pqv7e9WtjKJURr77Ztr3rKdnzoFXqQy
VjkO1dN01DCQzX4H7OcdXoj6LORqjXzmfMfp67cOUta42pah38baGLUEmOkb
OWrWCBwrezqX9N922mrP0gxnzbcd9FgvAdFtHPK+7FDJMe6ps0OAm24OBKRQ
zlHbnFFRbTVZJm4dR4icshADhH+3UsjDHEUuMSE8X9xecGkfUPQRAEkeyL0J
Hn/wKXHzTlyPt6R4nkf7uPkEudETTimSwEe5wflVlaYai0nGhIBKxIH5klud
BJvvi1bxMahJF2v6lXNFmrJd4p1G7gp4toOAeVRmX70cKtUTFk92RX7XgC/E
9wcKpB06YRTa78LAm7TnkLOV+dpEeGL7I8bdyaBOY9EaZnMy5TQaoXQcDyXv
qtiSRd49kZ6ajnGPF26RjfkfCtdWbGrEXXc5ynS2DSBQH4UT7AzOwvQ1mbAz
uskVemS4AvlqiKQdNsZpoyHzhiQw/BFLqnk5tDRCd2Bi/Wk/C2QWSpadcWaC
cu9ftEvoOaNJtrTLrICF7U1knMVpTGXnG+5JQi49qsWuqmgbfktl2rL7dvGz
iteFBUVg6co8AjadkHgUxv7CtFmkob+0XvwVj1vEQov5ufmB/nZAnCoywen2
mOUSgQdfbuE8Z5lLOrxDhg1NOO9Nnlv1sUMTC/UDd9kyNEOZZj+ca/co4bvd
+2vQvxn+YGb3J0zskVdyKhWz0CyvnGkS/NHfB0mX2zZs+HlDsZ+mpGq2EoGp
F8Q+EoP3zKyKz+e/cGy/T5ujjRSNtbuo2HJRg/GENEEgYQol2hC4ROEjCGxf
5HgzRFFJ3X9RzdZcB5YO0q6uLN+flpgWnAYydFViqFITmX2XeZSc5FYHmK7N
l7I7U5VfJAfgKiaY+7DTEkK5G3HnFq/TMbjyG6eH1v2pHrgs5QztUjVHukch
4elgivfJ6cDcEVITyCQQ4IEMAv3JhrZDWODJXb/RySFoKejZ1QJEcuu/sK80
JQEpK5IFU1qU1KFt0rEcZtpfSIWchcj5HffaSSbBR0p4C1uXU5+HyRMnAnOC
1gYQkAe+XRLQJU2uAoveilrEPZt+qxshcVn6DiUQUH356LmvqU0+2HHbcMwM
EMVZ1SwEdRBlOellCFNP1NWyWHon3Tqspo5GnybSiZXptMU/LiONfUztoMWU
5rx3Ezxxr4jtRhA9vAnwuNoHZG5wgD1bUpeqJkXR2prUOm8o1DGGQhFuCU+z
yJeeoOARXrWzP/rgpAYEJSYWdCxlU/oRFZq3ydKakUPB1ZsVceAfJTjyVJK9
pa45CXm982h/cjaEvlR9Blopi0iazdhGtMdNa3CYo1UpuUgXPVdE39tZLUKx
8GtKEPr79pzvxZegLgtgzH/wSpTXwmNzBz+mstX0A2Ca2vMQRMDmXD08bXzI
IAN4mtcokx8nJEHT+7OLCpaIXoDkEVchMGK1PxAJCRHtcsBgABOBImn0lmg0
U7Cu49ySC82HOvdEHZjR+A/soX9DVOi9Bh5qltk+5s9c+07PO+xslMe/vZPU
Urk7DZVLl67wqLXShXP1RhvsAN9kK9TU/PMajn2XL9eaUz22YZbNs6YVTy+Y
E2cDlvAbJq3MSOGsK9ZaybD59qvD4ImZBt8DAR5ow2uW5jCwV19Y49+tb14D
NGGix4eOp1PBPzIv35MkibsY6i7V0VBUkp/uszYxg4gloNGgpazmyZlHYVa3
pNY7QcH3qEOz/W0R7rarOxRdSaXLVOQEVUf2uOKMxCkoxweXuuw+YdX8z6zQ
F9zb+GMGrbHqKH4fJVS+INWFXW04TRJHYGe35mTfXRACbKRPUL/0s7L+a241
JJkBxowGVE0jfP3pNg0S6ypj7wdwhFBTK8iUCgBrUXfKru8y7WJZUBynCCAt
XQpofKzsEUZyloQwJMGmDjtGJQBW4bgptLtOUqil8HbqhvKbuV/pdQFExePk
Ww0dj8blqvOjFSxroFw6TDj0YBkm/2J2Z361tymlbsup9Xtyqnq6E952YfCz
jmoRmu9fiiTRVBZH8njtkkNFbj79rdBkippbByyu0JQDOEq1cPmh0HnZxtG+
rGdJEyQeN5szsD8zy4XcSiOsgqozgWdyA0DYBZAFYihgb9abhFM0j6vjDUgK
8uxrQEVaXQovR5nkS8fGIvQ+rBQNtEHOmsG6EkzGztsKp1SwctzBT8i6nOzf
Rl56tC9UeyYgjmoz81WONEWwy3E1IP+3YAwnQjHqT0Kx3oy7pk+0x/kMoggF
cJoEUPJbKAjjlvA17V9J05fTIJhWdK8JqnF230AwvAaO+19txP1d0OG3S884
2yNQNSFX/aA8JzRGeYMC7ls1t9L5kO7gVRYrKVoo4Flqo8cJNt7qrs/EYaIQ
uO5Qj5wlCwAtKl8hh5Vbv9GDdxjTAHWg7QU5RKmKQlp0BsV/3i8rL6gFNfzO
jtGfM0POLw6SuHFHtOPE3aip+MEfbYde5TjCBLUvLoJjscsq326qebdKuYbL
R2UulMyAvNKVwMRQqV0glvX3CMOipFiRahEVjDJK+lBzY2zkWXspsDKAkhmv
oessMfob7B1tPZxVgqq2BiMgWNPZ/AbZe5S7gLOL1MQwaCd69tqdE2ys1PP6
bU+veNIBc2Be62mu7m7Mc8k41umFk/In0n9m66wgxL0zBpY70+cw2cCImDe6
jnOVNsVU4a/k3d/h77wIVY3+TiE6djHDSNjblV9kRUzLm790Dx+ratu9IpqG
DsDgLyPTwemoW+Vd42ywyf2o1XzLQ+DIV6n9+Tt6fWzKfZZwDgb89JF5vs3U
ZUIKVYBxigU5X+nlTx5tago9Zcuto/611JqFJ2/VgEskmK7mrLIVhc6AH5DU
URHcJrhRhaYXwZrxGxGLjyhwX9sYSh2mX57tQO+oP5CLZKmz5w8a8EoGs7MR
hnUeeJoF0JlJDB4usXAZjqgZByquU+uLV/aRX8xOmn/4Xy0KEFN3wXIvz6pO
y6gOYzYSgRMk3TxBozDUIe2qOjgfpB3q43pRiGaYj7GZjIUt7Vq0zDzuJEwg
20+6wyQAs4cBqoKU58ZduAwW9nr0ODLsHZjtnc3PKuRQuREmpGGhZkvs5rBO
kPjT0360o/0sX9gfWO5TMSckGDMN3nfmJK4W73PVWs6jm1ThaUwykqBfz4lY
H2xrGAYK3+fOuH5enYTNbay+adTdePSREw6lO480s13W8CwPUYSB04GHLHjv
1Og7YLIr+UeF6OmgvGdDT5T/qrdn8vVgoxwYhHb4k1KcHjXHkst5V1Mmib1X
xRej6d4K1NneyW2nBH2iNkn3z5mMmHQG3bS8PEspmpgaqx28Wgvk2XAkFYwu
difKovJnyVIlKz6pJnKyXyDtMyzkLJ/yOiuB48lqiU1LkI52xTgcYBvW8jxf
zAXDU3L5QYAH/mkIrN9y3iDu41dF6PFAGZfvhO/IFRV2BlQQbAp0+LftTe42
bqRDrYdPhyAr4PsvL+nXyQHY8n82LyCs0U71MA5+M7XEtw2iFx6eeufv6WkP
hqIGqH9sB62GjsjyBUMiKtpo2d3zGvscFv71IZDsysukzgNy4vhEirIlEyoW
taTmK8BnxiI5w4GYw1aFPrgWXdNjIl8NnNjNS2rqLaMghyoiPVspRKGA7iGq
wL15MNpFJziFbjLJOkU6BjP+3vChoKyV4na8sSg3EeY56f6CAUPrOOW/8kQ1
+o6hvxWH3qt7HyGg31zp0oDUPueQFbrwtUSkHcbp2gDdRJA2+hZL2654GGu4
3r2C9u99teAAmG1HlSbvLxcYDO/95WJSjqzfGifLyjSYy8XHW917gHGn6Z/S
6FJh8DsdIj2k/wGt9ew+WYBT3LLlGkTFIUIJw8gGtbpc3rdPPykW83pZiVxQ
YK6xTHIO9w8BX4NjIXHaPP7gNIIcrcrM5zD3z02KWgeVdOI4UL/rw7EXRG+B
Pz3sjBP0i4cm77qUKF1oHzLLVmxT6jRZbbFgThvFhEs4V8iIqKON6PIHikFl
6Vb465okZ3teFKOf0Pa3xpaGkp3iPTk7jEyNVQ9ZxzUwDvm0M/Fxk+EQpfcq
L2KiX4pX0vG7RjE1gQfu0/5Vfa6jvVX1qMpMzIuEQxiwv182C5N0cn23x1vx
JmYH/Fq/uuT6VH5kJqdHSROpZITKAbgMu8LGtPvrYBDzlpLd+t8Um9WjKk+u
wsBm2sdiuDVddN/oPDADXdDbEppoXJq9yHpU0Ar8pjFLqT/VHDZoAD0kPuQe
psq1OhGcMMHClA7yXJ1OZO8nwnxjRQcZorgUSEasjOKdgCgJo7QPO8ej8mQ+
KcXOSEM2zXuISayZ2BNiroQ6scZuzXYaK2eDqXmwtYtVmqjscmbtv3z5frfw
NNDp/V/OtyVohFG1ZF9wRh7Ldn7wF80iAp+EUD5H+PXvHHS23yp7qrfugvJ2
n1YrmNt8uZTEvFxyPOjZUobRjbjGr7nXHIEDVt8ieEaJciULl2lxpX/kOMCA
UhUXLSIOvCL8Q82nnxfjsv4gcwooXKJojstXRAnG94zXO5/nUR4IkpZ1ao6P
mn12YOPDy6UodpuT47bDOR5jc0Ant9aUw1/nR+KRLYai+XQhd7+erPqS+oKj
X6Z7LmkO3CbTmBSHtuP96FQqx90O/BMUBaqRBsSw+5qATxOsY5SZOc6F8PxE
WktzQAfVCGhgssKQhViiqesIJSkRVsbW7QGi1hXBpsgktqvMjsUvQfnng4LE
AAPeulfn6b+kRukEkvgGT8TZFNlC8UnatAyKal0kmTzideqMCTwT1gArzgMJ
OEGXmjHcDJFDQEYg+t7gaHPW9CkgO1If46fCxmf+kF4LFNvGDmrtK0nuSC69
EuE96a0aqwRxHF/jXYBHRYoP++wm9SMPes1jE43Nx751fxDnjhvvgoibdJLu
fdupRHiTuaNoplUotZRXxLLPYiDWSxjlZQgZo90wfvnoLsEezb5bukW1HgOI
5HAPoZZKa0BlX7oVdG7jFMWVhOFyzkX/lI08WjGd3gCM0VCm7nTwh+rs4DTo
s3U13sHZYzhcF/Jcm9+LpQ7BBorWFAd0lJlhOGxF6jo+186rI6hDdeUSLzhe
Qo60PH2Sxx+HhVDbBpZSAVaqBIxAzs0Mxkf5yp+dSMYt5iH0dVU8JYZ7QWGp
ar4Kc1CgD05gBjzFevFuIk+1HaMTjE1vg/dHIJQdSr+TawQxv9Z0XDHi9+7Q
GwOKjU8+vhGfBbi0SIUeEfTOW1Uk2G6qtzA2SfHn5okuiC+NqcKzPEfjGZPw
lyiEscbGjV7I0pJcilGIZhW8z0nMmMQVnyrmTu+6BlZLALMYFnGFVl4j5q6j
dVZ7OJwfWj8+b5/C3Bj/Q7VkXIOqiT/nj+coORGO8ASMdWIwilfVxuiqvaex
xRLlWKfL1VMTjZF9DqJH8pyU/jmOAtj0al6sGIl2fcCWK7dAbYxGgbThAD/r
hD60hUM6BsXa9ydTPOJuHl1yQCYbCG2rnf+WGkPPmZ3niixa4C67OtRwxQUO
pwraVDBkc2dX5f/sgNm5SbDAoJwHCMTXuITceAryM+PY5U6hWh/sr1asUH+i
Nj8nNNBKc/bu3N//CgnVdNdqIrV4IA4ge4AH2FKO6ZaFVb6jb1k3YVtpdpfS
unY22FkKW7s3Yc6WeYQ37qYAoDXFvBqeMjFu11gIrxmJTPU1saxbvZQSZkkI
iKL9QxiBwKwzbii4/iZpUuwc2VxT4XVkqzCJhmX6d9SJ7OrphXoh8XOJhqQJ
gUUvPRL7OsiypkrIk2gbccIBv+FeW/ou5oteomPIyLG7QXPB4Vq9EFHq+xmH
E14x8fh5qMG75DltZWdFQepEr7IBVEBUekTCpiM0pDKd/rRzOy+sySNarFnu
Z1rloai68ZQw7btk+2HZpl5mpXzTJ+0wRUQPCQ1mPZ8OxDZW0+XE/jrpVyra
b1EMJ5FZ/Q5x1zAa/S1DuHOpVvQEo2KAkmcd/EmCc3agDavVjt1pnB4B5Q0s
NQIdldS5xx/1FPFw01ZhZ75k749Ds2kC+HhfmPUxdlsHXb1WB6GZ01CnMNyM
Z1n0f30NFLh/copEILSknqybvAAthXJ2/9NhJiLYNXPkDyKHCUw4TD98cEkc
HQkrWKEyAId8VWrRSSbT3in2Ln0xjaCmgeHtVG3Su56eKQ7pIGtkoulCFw7G
bY6LTYw8apXx2q4FtTym124EFAjK9UIMkPz5p35jqjCzgK64dHybO6XvsWDq
No/fREe2BAS+6R3Chonerlgx4r1wQthg1sahNAGqo8jI7V6TyKbe7TAXNiX5
jX7NPHisMhUajXC+Wnrca69frb9e06yoi4BJEL/Oxs0ghzCKsdbJZagaCcx6
f1ZcdlzwrmzEFQKVdEvUn2InK44GBhb8NzXE7o86MC8NThxaH4D3rBNfrYLN
YYT6RkPVMLhF3V4qIimQpLVa1pPIt3i4SYrZPI7Gemm9wTIIT2R7SLeKtlE6
ztXt7/ZlqBg61An5vqfm6ntF2y6XV7Zggj4Qbu2R2bv7CBIXKyLvlGJsR5tQ
rky8o1zuTjqC5mnOset8XC64FFB3A+OgDvfAPSz7EEwoouHxobyMS8xNsyWO
v0LVP7zpd1WIlDm1+yEZxfYKpKJXnPVEVtWx+YAgaLJihSVkFNxJFsWBkS2p
zvI+mHtwH/s0RC+bmvp6/wBaoDlgr4Dqo45r+W/i+3HzMXKGW6zkc5Y2ZPFb
dA3EZNGTwdLTV2O13kcduG/iXlKbDlXy0P28uOhtubbaJoHX1kADZ6O+x92F
kzE9Smf5qCSgRifbdI+3Vpdq+prZxD/VxTKRvJrk+wuA6mkVv+W2jT/Ciupd
6A6UGx/jJQG0N9c8G8Bqy4QswNjRWzRT+TDDLTUrBWIOu9OA8ZoiXIEuwMOh
4KOxEOUDJTF8FsgKWVZQZlzJHDtg/xYY6y1BPWFNhIGEkke2Ky8B9Nv8Q4qK
z17E+OVzjZgCdX+i7ywjXIvy6I9ew1NNCt+r/aUMSKyVjwhJ1v6qbF/nogg8
05u2sP3tsBoBFIU/IaWRVaV9sUbeC3iiF0rfCllisKhBJEJEfXwW4XSCdnxp
ASanVYaQ9BNf3L6AV7Hu3vTtGM+z0FYi7PZtwzNsg8vl0TpOvf1EKZrews0Z
JI0oywL7VmA3fb0bxOAT9xXDcuwXboEQ6UcVur4XagrZe92FSPUHVbwXfrVw
9z4Ck32aAs9cw+dCOlbSLmCJ5tFwdk7dcDEyNQioEDw8ZRmVF1CYRLvQT8pK
mnpZHJxJeyBtln2m+Inezf/buhm75oYTHQUQRJ8xRGpThxGayxKf1KmySfcB
Ez8kPlICIDC1vHUZ3jL9YQ53HJWNKJeWKNikLVjJbZ6cPP9M7uj5AKaj9Wph
lPc39jElgH7dGiH8IvCCBNonLe3Mi2UTosN0LkduN7fXX+kZ03CHZsXTiAQG
0uc6KdFif2Ej4fr+Dfc8Dz2KV+x/zE/Y2SzQJ6OE2Smjb7fKmFv6W7k5cCM3
aU71wQYsEwIBgeltNoBRmzCffgdr1I0ksWtYYlLvE6EIWdUg6ItCCZCkeuiR
WOy/Pqbc92A+MSJ+4sTEjT8G+ilkE+ieIDXV61NQVV9LnDQxkMemO8wo6jc1
zVU4TKos2WQrVuOBfYkHyzOZX8U9MKWvmCRWEtnpoxTq3jeyKrznTZeaIF4Y
aj+xBqk16v08GB29/ocNY23/wxvek5x2w6Rprjeej/EHdjuyEuLqT9qp3rgW
UuUFUJLtTtvEEtAnHVrft1kTlQqo3HnTyWj61ENZSnOOFFggy7ePQVKLfgs3
3xcqdUuRBpaHPYcwUEF9X1Iv8g9nruvLwAdtiRpWHgvB6hkQZCdGDDSwr1lZ
S4JbOyF70t8AlJnIcyd/NCJd9VyX3tnT24Mh7GJyyMpEftE9vgQhQQG0VC6t
CirmqimJ5+1h1sqJIAJ1Vq3uM30N9pyjPDyswB8/gl2LmrUZv5jWJScjbyFX
Rykv3rFixs1Hpd+gtC5p1OAyW5moWoh2ewD4/Fdbf7seV0l/gh1fePw17OII
ymldLdrdVbAAz2ZotPYyrgULMUo/oj/I4RgtxHAGtS4b+CaxWd1d7axzuDGe
q7FKTIDS0on2q+JdTvwzwRZ9XM3fETAujK6E9ha4+mX4F+CV4977HOnoGFQv
VMyLgtGFc5XJkqpA02O5w5BBaJ91UtQSMqodBmStAbSHLtafxa8HR9j4GOVH
OhPq0myN1KGuByu/l/Wc4jfNaCU7mMwXRE/LKZ5Nx+y/r8RGotIaS4fDVrWC
HaGhXquR5lxSGgFiyDush/8jK5MhVKDT1/UFtaAPPy+CErNe/+XzT+O9ykb8
52NseaY0Ztz/ap8P4sT3qy5BgC7xqCHDCOKdtmcF9phmONX28YEHcqNgZ3Pl
10d+0lR8jbV363YflvZdUR4kYqtrAmNv1XtU91MvKwbezQbxt46UVIqPCFu0
PgMAB4iv/mXY3hO6EKpQfjlCySXaDzcowVO5lqOFjiIH9M53txPctZNPFBeh
7tG6rQCIVn6y34S0l0aSlLiBJ2D8E4zjoYbhWXz1EOAFxj6ubJXmNvseK8Vt
c4iiN1I5T2zMeP+7rfdrTj93QXWkv9x9I7C2FWavLbfJK21Ct3pXPMv54veZ
1z0k9b9yTP7jIJRyluGdWJkwhKqTLxc2MbwxoE06RNEor/DjBrmyBy5SjuLa
/TrYpIEXT3N6O57qgmzGtt1mN5InTdKZqQzjHtGU5llfgEx5IML7ssQYXr7k
SlTT+PYYm0OB9bbjImVLyGjOTQc7GOHHZZi/BxwWPQmWxEJKuoZ/ERjL866m
xQwE5P8E0QgmNon+1AnWJnhBh/9Z0vRNtdA7DrKszCsBXsHIbTAL7sRYJCkG
A2uBCxdWXKgpnqKtMeGGjdpz43fawS6ZFTvNuPZlFx38fjPm6Q1FIhbE+LvH
7D8VTkHmqRN1NaLpNPFuDPaKSQvq71t1ZJtM/5uuPmLsD99p6QeVAOtwJBJj
IswzN0D26qQvjqfV6Hajd15UARgGS5kT+9IwXd7H5/lUETbVfweHU8SZSU1B
Wv/vOsGlstGDYbF+UWVH1rNIkg/DAsO+KR/h

`pragma protect end_protected
