// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
panQp/ec2LjI703Uq37dOvJS1hdr7uEmhbwCjSCaBLp7CsgwW4g1tC1K6qAb
81NNM9wMMpKG/5Gm2kn19xlOywM/SaH1YBpNTCt+X6JIho3fIYgJiH8awGiB
4RYNzjukRHjtdglyR9j7XKSucx9oN/lJOHDbMJdGlGXKbrphdBgm/zeUElx2
OMCF1baeJeGbe5iPG8ECrEoNf2luQu7QKB5H7CaggnEPOnSRjpnroI5C/NSM
c1km8Xi5traiffXPtgwgg+iJeIFmB8SkTqy7XCsaVO0BIDEhnA7EvQmCQKHU
2BTRoXeIvbWz+Cdbij9G5EDpZ8MtWDiw2wg7KCjP9w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hLjHzLK0SZq9oB0qq2zKaBgDRpzsLBvbT2KAAPsZ20hbp14w5vlZ+gbKca/C
+yJwNVqf0itJ3+eVmWsQ58aK6mXb4gmnEcvlB9VJ3aPz58JL1Fg7pUT5+EEy
vPBwCPdL6X95kiSWIaVs9017Nbrt5o2NK/Xsz4kZKtZ00ByP6waqVMV8XVUO
uaW43ih8vYInRTwerJH7FUY3Px/F6jLswL4sUfAKN7T20E3ykpH6P2BTmDkK
pHm+dcp4nBHHOKWawaGYocbd+eWjmeBhWWIrlV5yqNE8/qa5UOWQDIZhtdD7
nVVGyUjxaH1d7BgYr8Om8vtDu3xjLcIOquQVuggCfA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ggV0boLbH9LAzLUCM5naBCHjPjrwCrm9PkrJPPVNrfgbhq6ixPwt+4Z/bhq7
rh3cmiC43JsHJHvYG61CT/+YjxF5oFp1klPuy7m1NNyKcX7ngirvhkOEX3+9
vmrHymvtDIVC1+0zGQ7fe6EtLTU/MPg+H7nVnQAwujB1irTLD9yvQzD5eSTG
HuTPmIHRpuWFzICI7qsVl067KgedKOb1ypDL6yaQZfD0dzpmFVgdAbwVdZ9v
OXhTgRbTXfmtkltHH79YZd8Ec/5OfgyVW1YDGvp1EA7MINayCEgfKvBiriN1
N8bZod7UwRJ8YA5mHMvolv4rHSGe/GAE4pRsL0GAfQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q7pq+xvBtS4wIwRIYWEBRTu30zNu+Q2BwTNu2PqM81GE+TFMyig+MJ2Bhg6L
klN52K0rWNIGDRBXgFXpJiijBvQwGqYmlgK259yI6SzktlkoFwonPPaPs3QN
0P5nDl6XvvOmXc6CB2PQ1UH2RWnRAXPGPMoVfQnWRYsIQgqxMqY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Ie8++On4Tn44kfuUBxa/85YIAB7o0VUQ+K7X6IDG7/S5ald6t4Xe0DVCqWiT
FW2cCqPLwSHmppJsY+t/9SX4gbaKtLEUau6EzaUWJb9YKW2GPb895AgPsifT
Ngh4l/dVF2dyV1kBG2Cme8jl3UJFkgCgbUbWx8DGrs2Gf1gvSfjc7vkNwMTH
lBlPOnwnospTKj1/cj3ZXhNAnJJZz6d1odyWgzGgOp7kyxuIF/71mvcsg4Z0
mCcsHy6W68dpbDPLiCaMyxVEUVThLZMMyZnVX9WIYx7Jm5AHNKppbsftZcnS
SAdxAI7d4PSePz97Ku86tusUhoT0UOc3VMP6ZxzrFLejc5R1AWfoaIaiSo0+
S1HWXkxDYhDit3z8X1mCI0Vj0jHZPK+MKEkh33JnpiTX9EzMF/7eHncGeL2z
2QwgwIWYXJMkecQqtOCQoqlu61jme51dgglc2S8DFbmiR1eSDWyRsDla4gwj
bdqvrD1auneWz22nibOYSaWy7DosySax


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qjT0j6kQwiGXbekloXR0woOufozOSi51rC6sFqgzczEPNsK6lEQ3XBNY0wMc
c2u1zV/RFvhGNcSVhOZuDdRvWkq+5FZZs6EhuZj/YhoeBU9O9HkAe+mdnFS7
DgaDajD/B68glLzh+uKdvh6v6wUUe6KGKNJRD2Wmz2mzbK0N1ZA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SZC4WXv4htV/dPOMDiG1TzyPgyz/aUWC9Jdy0ZPn9D+pz7bzObDth7Qe+8g6
0k+L0WYw1dzZpaM+l4X2Q7sAFu5TGY0CHVSG/r8aoPB/YZq/Eq2IjLBylA6Y
8oWEAfo4UzvkGtDy/vfI1+Du8lDiyzGgsuHvIzWmQphoWSvpnXA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 257840)
`pragma protect data_block
g4pHShgmz/i2auL619bfO8dpBxChQi2rULE5EXURBNYZlYXGVY3PzU4YoUY4
GLaYA+Jxc59kfDF94nmJcP7GlfnJZR+BhUAbHceJPLCuj4m7xjAVgaR5765x
JD4mfl7tEf1Lp8YAIfC58DTa+dxd6TjIe8FYtS4qI+MX+zxddiv2APAdmEjY
rPHBsZvdQ+6V2r1TN/gZmH8ag7XOk6rd+4yMzmMDAO0R0vF5RAPp/SOmLvr/
PU1J2DXPQpBSmfQoWWBdfVzuWIYzkk/bFtO8LN5XcPRgM8MNj/fTZuBi0qp+
phSx8K9aTx+q3fwaVlVT/NOuwFSQlaNKjz7+Cvcw/efGdkiaLeW1/kyaAaLr
BtIULa4oua9y0OX0U5YntqtUo0e7vcUGrKn1AfFDynNSmRuOz4ZILascAr2i
wtq5dtvHJ4xuFE9bmPv3yWp0t2osWhQ1NNu/c3u+5PP4Gm2D3jwHBsiAqx0L
01EPkVu+nx4a59FWZaYBFEX05HWGtWIb71fjXQIB29XbL4i+nJR1lo6NUe0z
wq3dHyMymxDJ5ysyDvLQ2XbRUL2q9HECWa3vk4oO5pXgHxoBSOwyYQW7LQ1S
/U876SCwBZl410lMNX64tXj2Wz1aiQ4f68pX8EDd285v24ZUJeyBzy6fk9Fl
60Atvvx14MD3LTOPnysiVOyySGjY04iby2azkB3DjIAvnhKB/Olbx7PnNIae
05c7qsdQdn/25HAoJrZ1PSSdDPUUbEtYNIXOSH6yfwJWnt1oJza270Tuk7O0
l/O0F6/+bi4X8MRkjo7VKZFDsG+cCufYZ6A7FhFIWkry3nuYg2AfWCev40vw
AlbnpMOMLGpXclK3dZErB5LU6IpLoIWd5zGvXBRhdoV9whl4fds6tm2wPDP0
m5vDm+O3bmsx/WU0SNe+0817cKRXqzM4ZY6kVJUF+Fzb0HVRGWb7LihWx4dZ
sSMQVdKnmibmHtL97HTVnWjMHWOrW5NRugrviqADnBi6XElL+8ZRUotKh3/L
xowSgk2pg9CunAsjm6Y4EjfXj9jF3I6aqU1ygMTMlDXHKT9Z7OymogzHsppl
1dANeQwu7yOQgO1Ub1qijxAJdeNT1bwo0Pbab4Av8cnHD7V0B/9yszj24nIs
QdRrUNw7hTTX/in+x0awdBWB8o3d30dWScPqG0xtpl2X2RZN7iXCSA5AiUBJ
1ykLEQS1bufVidenQ10LUBjpeusn64ye1XuPSgK1HJ809/cHDy8ynXL6lEBw
dv0cwLNTG/pfLRyNwBWm5EOkFJHW9JjprbiD/L58ZcJUp9tvuz0jXsvWPp2M
Y+if4GhnpAvqE7R26Ns26uDJwYlpdgZKB4e6ZLM1jNJ/22ZLNj55chEB/6ss
OplAg5Z/b63zvON2yW6efouXzIfYdgHUW21bdMVAKCcJSVMg+pRB3woS895X
EsYsVortFj1nY91gZYV6oLK3asHHmVCj8gu8niWG8o0e4/eEbLKO9S+hnu23
KM86vzNPByIQHFmElotI6LGPCMvkE7lnS6k83XM/lzkIW4dmdSD5VoHk+yPb
r8GDMNHddmetU8+qhr3X7sDtFjrjplfNePHVNpVFgcSY0At1tmTzy1Zj5wkx
jN6E9T39Yh7JCVUGATXI4EZ/Tae9HaVhGdPcpqIfShBhRVYqgvSKn+TKVWq+
V1Z/kdoHkA5UnTJhqIM93F5k9OTUIi7S6PQyv33Qh/OInKRX0ab8r4DHdQDk
wImDhzzgQeKIyuZHKf0BcyToZJtiB79iE6F7V9tSSlQCKV8L+dGYGWfVHgNe
6rGjrnwdofGtBRokie6uGpS0qZfObsstXjWz/0PmAzyI9mXMrpRzujUpdy1G
fo8JNRXX2/HgDZO3nWc3/IDAFTUTfw0FpOlrXMB2rsStLBWg53C+28GNEmdx
BNmBPemGRbntYadochn+6LAboqi2UBomsZ2lwKAddDYkyVKvUQrpNGxrVZxT
69RPheE+3O9LSmRgETpWbZOQrx1l8J4duQJEBhmvS8iK7wFWty1jl/Pk7GD/
fopmcTqI/ITUkx4Rophybg6F+6jmXBWwCicVnfhqOdS9cUFVv/wv+fYq5+6C
QFsAH+8Vd/8wAj7aMyQ7DxgO/QqOIPEMxQqtlOaGzyh4f4FE9PwwkXWHrQZD
RSMvU94usc2MGkVcIHPL3rqvcQ0Fhae3KtxAH9yXl50Ml7j8aAugOWm5d2Vn
km61N8XqrJ5DWAIHkKgxD+I8k/TywSdbWG2iLWPL2Q/1t5A55NhAXgpY7EiS
fSaujcNSToaGDhsM488btDIMzV29RPaX1E7jKAJBGd4HKRRqDkMThfvMXAj5
zSZ0bE5/JI9w1M9TeUjqHT60JHZVqALKlOiVlgSzqE7waQw/hQIwLGGxYe8N
86xekg13Y0SgKGG/PdsAv/iZhTzXxg2HWF1mRlSHaPE66AZRwptTIFBrhZHs
NFZOchCCoNfQpVwt5nQMFpepng9ffdWk928ijOyQoGR+mZLycPIl/5sRrNcJ
XTAH8lld4ERpI3ksrI2pTHPTllU+eekt2p9xTz+Wjw3DXj00GwiANotVCdqo
YZVM79nYvpuRsxhFzt6N1KdiMUoelOxF62zMhrCb1xBQwViogbmyTYMLVnzE
+JrWwLpyjSRY4OnFR2KaTq8aKtDGMOs0eKrXyi9HD0m/bylMIB3Zb1A7NM5L
RN58GWzLhdJFFdNCrGmCQBFmZEY6IDrbhiPbVGBubnMLjnQUWFfrx/xKms7Z
Fz4iaylKtPUjWw0TUenVKXd0yOMv3lUWGfBx+EjO2SbV5Vpujrdq1wim43ht
cPYjbpzMAmYXKgKurCNdAlu72pgRG5GuFYgCkmwLcDelsRiKaNUDiRabM7SN
LWRyqXbF8oCcDYMc7PD08s7AgqR+NyuEaGBrZcIM5XF5wlVfsDT10sWq71LF
2xXJfZbX2ZdLlGirucbzSLfSgjH9M5pSsNHPmweHAM5Xax92JwdfZesBJasi
iq4WCsbWCmwFx6pRSRR2mvjcE2EsUqOlDRLVdtwMR+yRmMW8TknAMvKhylII
As2lyCgDOrz16Bjr+cXoVOI4haMweOo2tvIRZ2cICXKKAaTW0wetbLcGCvNn
ZCn1G1qQKufJmhzs99yv/Va05EDcYK4a2WZOf32X8IMoqsqd3x2FKsP39BRS
cK4gDNl4gQp3KeZVjvlhg7w225UMQlPpTmM/N686xq62U38dxhcjMlQ690sq
rg7elc/lKXMnH3Dq3vawGo1yhiKlXXmL/rSbEF/gAx3GnVZYxeYOLhTbJuC5
V9ZUE6y9TF0rty/jCLgjsC9QfrKoI6PH7ZcZdTREmqg6T8o0Kq6bTbdMYas+
7fFqgd1vP4EjTkFRnMrIJI/zl8baneLlLW3K+GvaDKiAid3/y6PAqrI1/4mC
a7poJEDE9eSJesfm1VSk47kfEaXBwoui7UCs6N3ZJdk9y5cE3f3MbFifVSxu
KbQq6OfCnyIkICrXHCmzp/5q7iJseYXyUCkD93xb7dJFdG0QrY87lmrNDDDc
djpWQOQJp6ElBamYIyuR/WcJ0FjuW1ZvIMGTIX8zhz6htlysoa15Qv+8GJ60
+UAHlwezGCwh86QjBLemTPv38b2TKH6TrV2mBb6vf/Z7QA6krS1u0y1nqazz
ALJxZidUxgiObVT5aSOoeryvMkK8uaMtd+9B4jq+H56Dl3C7Mu3Rz4OFptS4
Sij/uog3v9QQ9b8Bj8FhGZZjQud2momA4Kjr7OYI8RFtje89xqEu4z1GJEXV
UgDH1JXe2ON7rYKOZtG/lTny2EEIZCdwjdQfrvNJHdCfg9op7Zps5YpeJBwU
TE/RCl3FMF//akr/yXgG1sw+D/9fOs9WjmDp0zwKH0XN6XWFvQhKXNBtyHaJ
fIZm8tAg/KTplkumnlr8ZXr4bMm5Qpk9ncGIQ3Bgng05m0omaQJEroLJ++hM
cJweG6a5JZt1MyxZNS9KwXVu4zaWmJ4jQQhZTm+WEI++96cfYoeEW/V6n0lz
L1X9xEoXXN07guWGWZazKhFwRjND6cCdY039/b9gX2F188ZgI26bnuvVSSEs
A9nZkcVlu15l5lZLB6r33QNjCjb9W5xXRv6dmzrFi6YUd4ImKiAQM6JGn1qv
oPYRoXrL3ZhfZnOoRmTry6ZUyrzA/7lEbjbR080KtXLz6EKcM8nDsTA1mcBq
46VzWsOXtxTcCEVyj1+4OqcBS1mSXgiFvglT/4HgIvKoyAlgZYIs2qUmPKxz
GVRrdN9z5hglqqh34Fr2CNSdUR5axKiiJ2g1wOIa0bEozs3thnNIr4BYscc4
7XPByh7mLIOAHLyy+C8jBM25U551SLPewCKTUiYxFZMSDkUyUK+McLqU9UXD
lzXtso/JhDXvji3OIy74lCnBJ5xlygjQSM+KZjk4YbQ1OmlUBucFo89brkr9
SnPGDiT4hPSQFU7kxmoZFIFKiDT1+dOUJsopM08hCu1cnc6yYSGD5dObAlVu
GodV9oN0EF+QM4i5adEbe+0u9wICt36IwJ2moDUSnTYdoh9QXyMvRzyRO9Vw
VvwUOhgr+WHxsBKxSlQhTIt1gnZaBRpJ5kCZ8nwrNPVbwtEAz9qpA+Enp6R0
tuDVhMVFkwvfQWohapDtPTG7ndpSDn6kZ4q4pzhWymn8UDdVlEe+nOQH5gaV
CIlVvVvmDlZXo+QYgCiCnhxhO/0Rt4o34tccLUHbQCZkY5MQ3sCrvVpOPVlY
FbVIhnvlTHgFY2xxfi1K8Ahqs+e0xiVBO9nti5NAI4tG5V/JXuloHbsZyfd+
kRuTM7V1MiGuVeoVW/nREm8Ens/Y724aMdziPHAggVJWrkgNC2RLj6FOsEGs
rw4ECOOozjvUFNFRf6YoBdOsu45E0+oa8gBxFT913ae2Uzfhl44exmu+cc0M
0kMZb0KT7THVFK3FbOq3rrq/0Dk3G0scwOt1zMWOUW+bxSfPQWPRlt+ydpZF
nhsX7m7tZnBChLwDJiTaoDHp0jxSwvruQVtLULz8waArgB63KQmU1/BeYiOL
IO/94gRH2K3rShyWN8w0TEU8XYLmbIGNV+yAfRnzCU/yfskHfU5Umi5jv3V5
m9ESx1gKnfcovW5LIX2ROlGBN/wkGstkBX/Yz94+CDCLpBlJfyhNiIUuYsbe
+SlIkSvrv7kCIYK3OBgaY+hze+cZQ27sT1wmMMCBnJvop/ZUEBIpQDtNfj3E
dWfq6d2gbkMpNCtB7fnKf7HbWACDi2J9mfuNrELPyAxMM4UI2E0XLE340WS1
Ifq/5jzhhl0eZu8O0oEop6pUTqa3oFi5OZWBHt65rJoE0fFZwHTzqrq7z76f
xxGy0krOvNLYQvrAaDsL/uaH6byNI40Cdsvez2imqcsH9Qp2LMUqgXOCy1dS
ULyRCLh/diHSyt+5byAJyLbQCnM0OuV0n7Ga/Ru4bdFPLzacMzq3adtMwypO
lPEB+CkGffjJPxC/7dVQDwd1LQXk28A6yDtSSQJ1gE9LbpMW0wW8fH3NQbMQ
3d+xRBy51qPB+Eo9jNEoWwMqR+B/yYNsv68U85U9GXEPqo8/p+W+wOh/W1Dd
nLpBZJuTyzSQU3XEgWldMdYCvhaV6ED9jbSdnF5BRw7WyIU5QYrJK5r4ed/4
OinwiHggSzmF0FrDzJaHqn9aVgnIUq2dLG+CTCrlyLWbulhdALIMui103oPC
iGAA8/rbpMdAhfxAyTOEN6sEr3v134G+wUjWNPt1GeXHJrdHxJcf1aC0C9vU
kjmHRlyDQ7gMqPA7VVfxpcAb8nbSHbavWUjHWAPgdiKkzPqQM6iFRgN0CDqd
HxY11E9urdsd3caMEEI4lMIm0apDK/VmBgqg48kD0D5TKGx0q9CoRB886gBF
ZCmquQos5t9iu26Jea83upSqiTpfNXJwFcVIsXfRDJUJS83ag24gUR+SbyMG
n/s/qs1EPsekD25p5tFSl8k/WqgCjmE+B6yUVYMGUL4prMNFX4/7uvidLSfF
KhjyxEyA1+YFtupJ3tuJ0E98EhfziF2DEEqXGQ+9whU+MDT58gyprL9yvKvY
K+sQVbv3bbGrJcq8BXc4bmkUEx97RJW5/Zl+k/pgQz6UbzXtj+F29bCpZCYg
eHKj5rOjQatKVO+ft7mSvDy86bnDa4yBsYGtRXsW+nMdFESFsitqo2vI5IRI
xJOcibr+wV+EI6ph1hsMzSW5fsXoZsv4FTTiSpTcrHgLbfillCnaaZDCZEW2
TzjMJ549kEctRzhpo6BWvVlT+ylY4NIbVoBQBmwLH5P/YHSNTOj7Di/9lBzr
VyzA2rba0TzxbUA9zZgevTdefYLMu1+W3csgN5ZEI2DTWxffy4NN3ZGIy1TT
XblwKLBsMexOptLzOKhEwFP1y5akezAu8ApGUjibtwOsfvMABYvT4dFjhNaU
EJEcyePCjjXxlstV8FBTrjTIPjKCilUOpDGoDFVqyFkmVfjmAl9pOl54c7i4
YEvLsSMaJaX52ZfGDtPPhmvehti7u5kMDDtoyvDVs9p/ZRDYgtU5OJv2Mhuo
eNWfLDnY5PG4iXXKO3AU6OhJAo21liTWRwrOUm/KjDMZPqUV4bThg7iMt2+Y
JebtJ9UV0QpBCGkM1VOxVO/GIgklZqUxiwL/TT7Sfq1qv30WgqmumSFKGExQ
noennF/bIex9qxmzTatPLuxEydXJdhK8yXVI1cqXvU7lPEif2o7/GmQ9eXy0
InoK9RI8Z3UHlUej0vFErIybOpNVeZU5NXKHilkiw9+2+IAKoAREqHHuzFij
DgOVOHGAPAAI956B41x5xDdSs9VoFr9dzwHoWqwn7mESfARq0GhQVm1o56/4
fXw2/HtkxbNLL3Zh/K1YUXJ5Cg84e+qwbDnUAwoTmBK3lnrrXzMi3ZldEaZA
FxznA5Z6KAENOMJ5qioOc2KX1Lhl5dYJ+3g0lkAE79Nvtux/GlOQQ+T86BQ6
SxJWCwgMHhahTC/+CKZF1Gz1Ouk5U88unPKZCWIaQC+Kq3l4M5o0BSCmPK1K
f2zoo3+T5eQ4uHpBSj8d/qqr8R1m9hd85Y4W54uNPS639O5bTUBy5jk7EXDL
FPmHIsV6RG0USG9Kg2RHc/MMaLtpXvvyiOxEgCIlqvaN7GdMjqYVIOuzcdri
5/jLVIRyCbLJ56rSLcAC78tB2ao0mtexpodwFSfKbjcJkmYXZIkSgk+tFFjX
2q5em0HSn0EcJ0CoN4JYjX4d42lCdXhth0fQ0vIxy+GlJdwEYF0XLZRbqG7M
3s05uRuid1M20uH19BFCHggwz4vTqz6MmnIwzycGDAFjgk3GxP4j68/fgm6R
8mZv2NQfEtf2MqClumb3U1gmsQmNQYf9mqO0A4YttSDnj/SallIsn7qF2pke
ODI9OLtkmWgjcvGlq5fYugdCFaNlMtKAbHKAza1iZUCjI4ks3SvZf0oHIqj3
kaCt4ujyy2UxUX54X5hr073fe6bY8WXofCGebtd553km4vGVlL6oJA8XAcA5
sSlEPvXGNjRQIyDDZ0cpy556IjJ8/LZxlvhQDDQRhXmLPT9EBkIvb5bwjjxk
i5jDvzIzRqLEFubg0xfzdDdZCrrAhOLcaF+AquYVT5Ub0zzToExFnmYdGyA0
RI8HYIr3FhinGr60X/24l2jxju9DFk9gH3+IctKasTGdRFi1NLH+yJ0sRIBN
rdSZRqaBexec4XDQkkP+BBqABacBMW87SG8s8t9PYTxUx8nuPrfMuFRq4VZK
xTuRKIxgYh/Eobo5uNJlLUTDdKgTeAH4QIPMnEDF/MsU/1/1ySq8yKsYvEZc
+7AszAQWb6/gsS40w5awCwUbXOObGqs7jpSCpWLZK0XFwo5zMoJH047vOZEp
ehmSqpwP5Gfrw7Wkef/P4Xe8KelvjCxdh4D9sSIJHWQRa8qy0wOugl0DJdv9
IMtDl2Yb8W1H1Xkcz1w+PphDB931FHEiNiLdMmCOhyLNO3iAWai3OfELXGta
zZZLsupDpyF2kTbuwJdDp2wzUtaVPxnPL1JraTOxA9OPkfo1qc9t32JSGr4C
s2LX7wN3gsd6DuhrlNnt1ncRflzZYexKbuUTJ+QG6pYco93AxWQ3Vk70bU3c
PcRqVWKN2aoNNAgg2Vqn+WRL8mcnaRHGMzu2WVpIK4E7Tw2WuIN/U/lVi/u1
vzNzzFVK7iJpfjo1mOItrKboHdUHTfVX5599Q7Uh9cF0PXcxUdaZh3lm3cY9
Ail8ny/RYCbesvPTOHBuFUBWdx5g9dZ9XONWjLtNXl8PKhocToKx8JX1MMEY
SOy9uj5dL/3ewmlimtdoQXyX9vfmvzF9P/mPwkLnrF3h+ExjbGCTcZ74vjnY
reREiqP4XLkt5y7uOSg0AET02DTphES0lri4onq5Chw73figIw8OVTjiXjKq
vn3iL6fcjpvtaaicIVzoEI0uK/ge66v2j0i5AAm4A/vZgkFOuOWIY7meGS44
mdCMQcjpgH9udptFL7b7+JRJpFPUQJ7gbza8Y8zst+O4vteKCSYF8+i8WHIg
mc1Fgg82MyXZFlyt8jA/WUp3zXqRBW4owgdGnuygHfyzhKYQPcse8BLqJP1M
AMAi3XMtN+zhvfQjDHu5s/T02U0jUKXwtv+CDrhLctuAQWM8nuHw2LoEtqr4
hRynHuPEcqD+5fGYoWoJgX4zp48aJYE5Y7pIukbmgJoX5tfJpQDWVFzKP6W3
40DziNGqLEKFRxoV2S51qku3rQORpVLUx033NstAu9pm05mq2jaU+hi+pSQG
+j+4GXwkVBF8TSEnfyY4ZWfjJx9bs9/xhtuFnnqCZbl+hCRhL/RaGUGlZOFD
/Ie2+Rt5zfiNeuDi76l8zxhjaSUL6dY8aWwbNY9nt+WpVuMPt3GjnhF2DXaY
AMwhKzOptUL/nk7FwEg6m8Q3fGjQn6W/oTYuaPHBzOxTXBv1iYZOj1GlK4ma
T3v3s7lGDhEfX84tI6v3C7yVekJk5vxsiz9Tab1F4rT0udv16JjXy1w3nPST
F+GdGNfawJw1tTIjnjBT4NWfVBoWf2BQmksGhonfItqtmrVOlxI6f87/3XZX
ZHqlUKaKyFrm+Y/uuvHjQxm7EqZ5fZLySuFnMXuPLQ1RNwXuzLr3Gi+vYJmC
MvRa9mECtEVyNscWpdzB/0efCUpGC1ABsVyN+wiuOnNXUkzWzKKaQxMs3Bpo
jKBEten1vFyZSZ0to4jZAxyuhZOWdZaZ70zasBb2HwaeEVpBC4auaeWy91YS
GWRZNpezfOWvdJgxXvvTKuxmMDxEUElMJOzep6N7Ki/OdQwvzdZeRcJXChcb
wH0haazAg0ZhqH82i+DcjtU7zgV5Z2mgyIpwQiG+3bpqEUZzWQa3y91W456l
lmD8zoBIamCCbOiyAcS2UXL9B/83kyZAy3/4VwSiCrO1fEDBWezXLoHAkfzr
zNVPT9uRoHryHtbyPaGaxaaGDALuCJj2VhRAH5O3k94BuFrNmu4EoRZEhJEf
Fln4DrytIwpNBurjYu4dbYoIzUA6mQZrsVwfRtvbRcYNGi0Wl5BgHH/PyOW0
lflk7M1s9nS9POtp8WZzn1TtIE/1o64za/0tNQJID97m1MfSSi0L04+edaq5
XT/CDlw5kZzc2zOldLQBdT2N0+4b5BfwaRKBp2T0cim8XiGyrkgvaFZSh35P
QPz44AbxB5k1lI0+Q9/S9emVuinaOsVApS92DDPoAbVVtegCBL07C9+NlRX1
NOVdlHLF56WorRc0/aXQhASww6mF3WHw1bQREKTR73LIiCEYGZIPB2MYpQmb
C5pdskOjQ9PPjPuYu+mRI02nLBGK+xKKAOADBkEwykApeFe44Nw1Jcge4Sld
D6wk1014aJ/ZeC5W8MZH3S4fs0vLUsuL/1ipqeGBHrbgz7nQpttwRbeXJs7z
GEGfxL8OIKY0QacCi6tMBSoGukPPJI77mvL8Bkp7aLdX7iLPeSjpPEWa78UP
pD5o+ZhOvZGRreRL0YXQw5F335hHc8uEOz5SrwVijebCWRV948ym8wsQ8z4+
TIPdAPJ5XS5Ww1VSixFCeKPIYysiDzwlsTauKu+3AqWqlXzAgVVD/ZbSiLpc
SCtHdZxcOEMmTlPfjjkNCNpaN5CgHTyMCV/TNVXH5VOboyJsmB3qA4zN85g6
d0O4qdba1O5YSy48/ix9cjd76C3VbIrt8TaGjKFoCNZPwlVOrtx0OBKpGR+K
c7R1tNx8ZDfFzrBCEKyVi9oqCGmEe7tPPdwjL37c8qu8UrCNWa2+fNA9k0Sq
8XRnvtks3tRaREVsfBcfwDUUh9ZLi4jpKJBVw2hES6xea5QTg3Rh67mDhiqL
uUKxG6HayfpfAwp4TdoNfUgIRKvK7yZEex7D8zetaJbB8Zs1WRJsEpyV8CgD
P2rq5YP5iaerIbCM+CIwmUp/1PYBlolj2x1VrVzIJzN6qD8kh6/0QksE+k3f
fFD2A8dO5NUB6c4pQisYtAUj1uHS+1gP+TLwctiraylkcXwAFRCRmCLXbbul
HBejpiFAPj2GJZ6uZYh2ei+JGwWGPAxRBiVQAvAOy+9omYlfpIOoknbE4wnO
TQHtF7oLpD1LKsvjl2ZlQN+Mt39wmkBQvZdbxFcEv32v8YLmNAflz+3vAb0N
vmjvmT4pNVuZ1XWI8ki1GMVjVQn9daAki8muxa6G6IYzXcVXiYByDYyeXdHX
hyR6oqzCeyibhU0RBqWPi53RJGoo+weBH1mJJRCIgrth4v2TeX+AgjjdZurq
rLFOYItXt77LNo/6266CpowpzEaGKZ8zJRglpgp5C698iTpSz92yAGYkLL61
OjN1HkkhDHt1sgJUdS/7lRVMOvykLejOSwinHxoGW0a0ZW9EjpQboGv0Vdm2
UVCKsZe0V/qvzuUs8soFyRvLZmzsG0vdCZj55H0g1ClXGArV2o4bPxs5f5b8
bWBZ6b36Ezr1LoNYtuatLJbFsSGXJSaJhThmGJmjKc15O5G5JIieqUAlmT1a
z47YZRBBA8yHiMOnWh+TPUrzwv7ekcIPbV4npzeV+NJAqa2a4xtY9pAVaEfY
/PTHXUT8CQo3PyanonW7tRjeHf+QhQlTnljWZZLK0DcPMLVe9+BfsahMjfCW
uO8TOXLWnHgds0/hn/CKJXkBXYNfZbx2EnyMtDB/wFj8RzAv86BiCawJ2j3I
/0vfK+cosWzrPZHVhXmQppyiOmHFrgyd55TZssg91k3ETpL+gRU4e/uQE2Bp
DGd1eaCw21WfIMNlsprMqchSPGxmYFrVzJcp7M7RxAqfc5udtzyJ4sDbCiFT
z35euZVm2GKOOxsAGF3pXVYTZw0+9yw9wh09m9zMxq+/3DXx80k67jWpDA9I
RZa9K8oQNxR/pp7/ofVlSBk7RULjCyRuzmBpJ/KR6drkNgp9/1kv67xn9kUQ
TtKs+nGwZeLHtlJvIx8a8+YKaq7pA0B0YyrKGrxIcacOT9UGUvXVH3Q61UXd
EqVWIRs1kZrdTJol0LjCOstoWWf/zoMGiM1TQAZGOaMAJNxPojxYzT1w4XhQ
eGD3eaWBtDkBkvJZy+H2YQzHAAAQdtPxXK70qSuxqXs0duyDrslkZmNaCgNI
sB1lUZi7ESfjr2VCgNzOymcQ24/AGJ6s+wp2uqWqy7TdJivn5F9HJ5zvTqql
eFoXiKgOTE0bQc+hRaNIHl64w5/a+HnpOVbIjp9kPJofqeOlf0j5X6d3hfqz
FcnyR8nPt/fyH71qddT9wb5mkSv0aWA7teEsaDq+8Z4BiJ/JAfhCSa/Sz9+b
14PpYEPgdfCGFu/9A9Kq1JihJIlQub+1gwNXPyHnlR8OClaD3ecDg68rdBd9
LGFbiRgxScuXDcOR6eZDRGhDnJLudbYIHpnpFYn5hcE64aT/3Zjq4yFy4hNY
r3CFtW9nUOBKwEfeVUexqVarn13hB1WX1yLopGAa88KgttVq37Fx7UIh9pn6
SknfNA9ERiOPnqwDg8sz6Txq09Z8WV7ZSNjpDPoD/6BUNJbnX4Thr3VokrLp
HvvGBY/p388cvvhxxDKHLIXeqMmwOka832bs5YOWUhWgc0X8eGZ4yCvWa25Z
yBKkGXJ9tXg4CJKJR8kdzePQlF0zEkHf1597AVzB2/LqNf+GJXu7qysHnfIR
U4kTvkrWUqq6VriIrfeDyaMYiQFwrBxV8jGXunHt2gsvyd6VP4oo4OSvD99F
Gd/S95PZ0uzp0CQphi/WRuA32KpJYayYxtuJqfUMnNUOmSUOqYIt7MtuoF2t
aXCiDSgyJVsjN8ikApHtHNAZ5iyrmteb/4PsNcUuJMki5YgmRzkAuZVytu9R
KQRwSMPku76a52Tn8Wmadn3f+RHbwnChEZVBk3BVSeMDxN3V4EXvhtTXwPLO
W+sFyiIvqwmCp1So9mRh/KTL+J40KmXRYglk7zbvbRN/fzM+2b401B/KhWeq
WpVqR2iY18OV6WGPx6kHJRexFriV212nvcV2mqAbU5kmnNYf9pfTAbg6wHb1
qrAZR2FsekEvSN2vSu1qUFrZ4QaUdEXlqrDuh+3RuoKTZPggRhyI/ujA9336
ZTTy1qHLSGmiL3IoUinrFit7KaQpvf/Izz4SWyPz1FrKJYfuZHSnnueHdcC+
oME+UlSJQU8Bk4EvPF8EJDuRoYVMoRPLjv3BzS8dSlIyOSR4dfDRN/yu7wjI
CTwnL545o6/AZEaZ8qscFcjX/OcmG2g9G88BKkHYiVhMZyuKO4xALQZcgENo
Sqa9P7WNpQJf2qXHA85Fbztb/Oc0DAgRXam4chV8UkgJCt51MdMJSH2ZmDZg
QPAy137gBNzudDeC/9Gs5kfioQW7AxdAwXyUX9QyzNtB4XuP4iejFsj0N1at
jKv4u8gQAvmzutcFgnCtYtS0/WAu5DTaTH3vMs3CaBLP1/C59bS5RRhROgbz
eWM64o9IxWaI6LzH478pqhaCChKNY5TqzEQ3Rx2jiBqzarlMrAAfyGcU5jlb
2s6KrRWhLZAkp0RWXR1mK+VjO1YJ735fCLr0Hmds1eg4TKMMXTZY55AwU2Bk
XdAgd4HtFOSw5mk9302Tfzu1vZpLJk9Qb4yaThSRky0RKhwQwJemSCKbSLoi
abTAd9Z6IskxZHCLjfdivRgnffkIMyUGTH5hYt/dBk8WX3OS8sdn+k0TPHru
e1B2gRrIzyr1ngDyaODm9dLmb/gJWiloAMmjOGjDEyieDT4zn98uZKSB4f+g
LN5UDAnbB4HvAMyjWXGBi8uFGjZI3XQdZ/dpZxtWtaVe6h/+Fp+NAaFb0G1X
3b6xeavpM5Z9IYCJoIJBOcKCY0ZEIaQqZlUTmIIFGvI1Re0BRLWMRO5RdtWj
rNWfNhHZaEGEuoiGA+DNcpNAC7DjD6UnxkL2g355toSuwghgrzxQ9LlVT95L
sQ8WmyHLwYQKIds9qK3l/RO5f9Usi3rZi6ZJPaS4vpZL0Hlr+xnblqPxyQDY
PKkugDY1iwI8NGEQO9QlLWOv5k3yUIxp/nA8Veq++vKOFqX3+TF2nKvXa3Qu
HTp6GBMBC5USLPgZzlANHZqIGzY6n2sT11AnmMQAHKWzbSdKB7jyNYhaMZKl
Oy9h7LHeq4/q4rIOX/dS9rC3AIOVkI7MfJMRgqm5BlEgRb95a6ihF4yJSMvG
+rlGEQYpjM4FsSX0WGI94jPBuywAg76RMDXGK9kqUo6Vic6OMH+AoJ/lhX3k
B759XKkBHH7SjPFjxpkyYSUBpUcJWDVFW2lhyG+1cy13avUKiZbUSOYfy1Dm
7bB0EkPvNCiSpu7mUj0FbRAPk3pzsuAWAFsQGaTXhCRFBrP87yASfNjRT5ds
839/BVo+RRe+PQOzhUlKEYUozFP7/jySaVZ7z6YDds020PrlsQIWqHEA+VSP
LTOaQRgqCtZTeDm1MwWyQzYWBG9v1Jqu2vuTf1U5/Ez8f2CmdMVFDggcsbU6
48JyqGRn+OfiW/6PlLUdzytc8dvgsCoMhWU0H8guamc8ZHSqUV0aRmaXuEFo
8clDZJiRN3QiP+V8CYSCpf3LwSQvxxS25SWEcsAcU5zd/l35+RX/IP/TJgyG
r0F94MJ7VSe9fH7yrh03+xxX/Y6KMr1Tv7gTW9QCHxqbFpBcuaKdr6TjqWmk
raonrMbQvMy+8/loQUpRnpP3bUcLskZpZivXaEeucY7gbEwuUfVjSBaneqJy
dD8UrYa+ybOuL4/4UCM+GV9gt21drMsDKVgTxVIq87wgYm0IvBUl+Vv5Y1Wq
J4tmshJae4xRcX5ZFlJmlB1exxZoBuLxyMhvRFtikA3BKRxJaoqYJuDh+Xib
Nkpth29Tvy5rh5rDEhd/7+B307iyCrErD0x/nhIr9hg5jC85I5XE9qIS2D09
MQfQo44Pa+dEWlUrPqxVKKuQmJ/NnpOkevg6DNhuEP1+JE9jWzGwG0Cqh14U
SxSo7edqlDUlNmnwdN8wzHi1HtTpZnOuYI00RTs4ueEZmSG73/BtZVz0u0yp
aD5nxaJllKrMnb1DDcPLiTUY59fpfurdsMuZNlPakLtGLV2YanFLTAgrd+N9
GDXLU7M+3VuxErb7YvR/gzvyg2t0WMbsYYq7ClXqAXIlPCJqHZ0Q/WdCKIl1
Ety3IeDLym7Uo4cmbEq5R5F1ddEMN51x03s4Bh7AtZzQPeD6T5Roort4dXnH
hweJ724d3RnHnsDvtArK7IAUAJrN5C6CGioYS+x3NtVIlx6AwY2DK5W/259p
jxcYJzcSqqv3zYwupEY2o9NNvKgl1nwsmrTMIWjZ/ESI31cspxXmT+oaZq0G
9PMnk7fc24vmcKHAyDaFjVCubr2J4nGFQSQq9ZHdr+aw04a0kRphCTqJK875
We/5f+R7u7DCwvB1QmJbHEuEn35UL/LepY1nTP9/vzBaEyHrZ3aq4vO10Wqx
sA/5MMidGhkg/6vMrg0aTHVc2x4oirYGhGpQ/3Iire4p/RXjkO6W10H64nVa
Nyzo0wqOMnytBpj+ch6Fcx+PpUGChXXVsbcZE4D9q4kHf0K4qnMuWyYxYRXg
84f/bCogAmeUeRuPrytLGptpRHntbUGfHr8pjjn2iVxTFnbEJp5+2pYS57rM
VYmdxChD9LOVQx6KnMz2GcLR1EK+hmzDQIDaLFDDALtzHbUHE8gMlOkX/SKb
+ByJFOpmogFOeUe+X2Q4lYflf1Iy+UXITBPbn7GEl2988pzcafDScbL6mWnR
qf6AM8FATGdOBPKfH6O1UAab6g+C+beECueXrtW3dGVUpzxgVOUgKyS/4qr5
l4Tsqic01VduIN1rGKBFDtp+fCEmx6kYlk9RhC7NiYYR73DpN63gGldJZEXe
GH20vo5d15QDI00eKGZORvbTP2PHQEyl44O2vHckpiZbcfnggQb0RL4kY0v0
HKYsVBP4GaGsMmpquRJgVCrFvH3QzBIwaimzldfCFBbc0V771BIi9s0aCIGf
AQ8fvdnnX8IRmIBzBW2DNKT1VR18vYEb9Wujeu6kMNpgbbvKhnLqc4CMpp2O
KpUwcrnSaRNlpJvZ4ShHxl2X8fVMX+30qqo6Zx2DFbJzSSDyOyGRErPvGIUG
G7FVP/kK/cibNHt2zxfo1fpVuXx3aY8UAntBdzNiEJYWBlJkN9l2Ot41Jw3o
Orbl2k110WcHR9h/TB06ds3/vFKG+gGw1OCWhYC8N1mloCdSGk8w1sPSzzLk
ZuPt7W0FQ5+94P8kpbq/jRvdLiPWWWPSfVmsljCidve+/B1mjvDhnwoBB40K
OJ6ottMav9iZndsZzG2OQM+aEB/vI1QKapLWLHET/sjW27p9+muyDYFMIqQC
YHCFfT2dzo6EkUXbP9+/RlsDOljBP6c+6Fm2W1JwvmYBL0AjjYK6FY9WptDy
2mSwOFJKKp/6SOt/u8WnIShZxThQ5fotXVfnuXZ1r5EtNZR4GgBX+N9k6XJ1
8XcRl9cUbHsrNw6haDWbnnacMLpnzOK2TSRmAk9tARPeFZvvrWSf9tWODdxP
AU9vH34C2QWoCpZLH5+GiP5yFEKf/mFFKIusz2ZWyAu294GcWCWjy4A9K5Du
HpJbtQA6m3FOustIWk3KQm1z6zdRWPk187TlhCOGaVmBLmN8DyZRMoO7Kc8I
NiGx+YCx+dPwMoNX6YwBQRpANlTqZK3BNyd/t4jE2LwRfKs9iNefJxAM7Jkk
BaTRrl4U8bEr4N0n1xIy9do9nukxq+csKQdgXENxYWwCeu48etTJixqJQpxW
UJE3O+alxcYM9JQYLYAK8pjUjJ+EdR4ifT+9N6atOLRqy8mKm8aZl4mNSil4
qe/PytjWPOiZ3qP19iFem9bsAIOL2gwtbSaeuFt4H3fendUBizk7v9yHb+8J
XoVq9/JY2dfzR9sd1ZCrm6gGDf7rRpSvWdRKnLU0n8EhwCtvw3fVM7ZWNxvy
hsT4ijSMc54Tp8zyEMuZZm00sETmflfMLpx0yWle342iL/lnoVlTHByVxxbs
V32ioiavf/l5qqJE9m742vP/zaUXJyWFPfvPS3RaSxzkwfFbPH8ERsakc/ME
oibEq+YEkEiTDTbog0nZRN6rHim8/j1QDILuSWEuNfeqt9CNeR2QjKbvrAtR
lFr8fl7Bi2eX/Hwc0KXbY//WHTH3sE/57McnZqWk6UqrgvarzoVAfIC2d9zO
SjEolKDwxmtT7MTYK7vlVWG/tZtgob1tf/Pqfbe0hQdEY3dzMj3Pp0xKVkll
QmSfQAT7KL4Ae6p4eiKJCKOEPi6jU1wNFwNxK/zL+SAd+o/UnNLwPgzNdoRn
NcKEFekxTrqn7fBbad4glBdUb+EBe0nesHCTc8fAx4zrR/kmesOfjUle6p+d
VuV0zPX2hCd7HhRq7MGNtfk7Vc6ZkRrs66e0citoukgfw7qYTWCgZR8myz7p
QIbDBH1CwnlKqxQTNGj3lnk/AB+Px5Y52aJfCcZD4eoQQdv78R9digvgCNUG
H/71UWR+YUq9F+gRnC1736WpOcsrEdL3V2KMRfk0UZJZLzzmRgkjwsnVHX3W
d5X7Iu092DGzrOIpDVVwMbb5OSm+Z0G12hXmMdGWe67vAQcZ8SUFY/zOfV0f
qYnXSLYvEf+CA3i4AFEHruwVt+oo6PuPemfWGYJjBHaaD2sl+nbNc3Rf2qqZ
sA7SAidXTnw17BkJgkI+/vRTaiaQlbfSW3oqPIhrcDkXKIfmGDcpaBZ9rVZG
eED/u1IoSS449bs/F1Sv9CzJjkZh8jMnRH/KOcZOfMABJM9h1P2XMEF1YNIf
kJP12DfxiPDLQJi1VnCyde9MySisBy01KEOzEwsRsMpPuunj7BbLzBsqBYDj
0karkDZlCc2FKl1HHmPIyyzzZ98X/eDzq/gKjU3NlPY+mMfPvIlTWDNFYYYI
LQpJRxGQQz4zzYjSbBFAPi2VMevmvYEaqJoFsYnD7ggQ+NI/+F2QCgZ6/U3q
mQmivcOQEoLVh23D4fQpTUS0VqBNyUQ7RMg12b3yozLBOh4tYU9npAOAr1XG
Z0ASLIsUx0EvBt6LHhqJsSGpkMCasXmvGSG8Nf6Ro3IgqfZY3Og/rAid5z05
TICY+xlaqo6hWXIQvV/cXuSjKhZFbjF+JaIdZlbE+1fGkl+r9OAItonlp02A
fm7Y0qfWNO7K1xaZyPeP26LoDqsm6iUBsvvL7vl84NSNXKC2IAsntsHbVxTT
e0VSemd6t8p7Iu9zZVCUzIGohLc4bwX5sdfm82IRIKvtt3JTFFIskmszn818
YZ+qcTQaAIUhsYMw4CTTei9B/QXI2dUKkbVAAsGTal0TRXGVB35PyeJxaHX4
/ObNWKCuBaYela8bnk9hC6CRT46lAMn2gLJ2dAb4UpwWM6UOybSogRYwOmmV
p/QeWsDbawRFccJnicBhahHIC58qsi/p1bqCEKx/6SauJSj5qSnngumIxzGd
xuIoNJ6wBrtGYeJ4uei9lnZQ7MxJziWeu4m9KWDoOEC6o5/8iY0dA674Zsed
RX4ShZ+bxk6nJbtU0LJTUMt0k51A8ygnJvljQJdZrR2EvTVARZfe5LYngmpG
etn+Nn1rKvFq3whRe84C0xbOdsKcm2UvykoXgq5GfnVtmQJubbHQItGix+zM
2Vffom0l19/pGnzo0dm5hFka9GgPd5y21fNFCrl34z5oLkM0SFGVP2vcT29J
ZAbhmN37HtBJXKbXVrMcE5qSNsCHFf4Yy05EKMnpJTJz4nVY+dx5BQknMiyR
WRtMDtCWDTLTIOFEWwmrTL1rrwlv7MbumagkIrQQKhoIJbjwkeBME70nMits
ofaIW1WrYfDE94AAiEcR/+69s2lCC2SOPUUWXLQckLBIaKb2tNtkMsd4JsFs
AunXmFJvfI3BTAqhqLnWddOwn+jJGP/ddtqswqRYZ/xKQ8eUCokfUi3mhkbA
5fzj4xltavREfZlOguMeqC0VSHLE+QgN5UsdmCMiH1wT+uVH2xb9GHgeqIHr
dlL3EPhOqcbiDiwQyVS1LRC10EFe6L+hv+f0qRh7dLgINpJJmXrOI6+a3uzv
6mWfXHi4DciQujWbPyZzVI2+x1aSI0D1HfMQdAlMRWN0sEuPtIBNJ+kq6FWW
jG0S2tmy0NGDBrscL3ozPs680uSi/lyxNF0NybN1px2Jcf9hjMqtFvqnOtfm
w5golJ7ZyPKm9oRUxVATcMEEM57tIvVj0T89cbG1HBLRp597jL+qMn6JJqy1
1U+SNfCv4Fhkn1s4qVF1oXRpjDEn61zSokmRBWYKmKPZSixvb4OahwRHV/5b
2ETboUVaQwbxVBTugr36zpr4SvufL24LETvTurOWPhYLlantbGIJOFlg0oUq
92dmyHHilDg1aFx6Le9tXcLsf4jlH3UoIf0RNHoh1oRuyBSOjnSEOvb86Ng2
f6+LRb21+Bc7yCnBWdh3h2w2UJRKtR778xPv9FyAkzyH0zSXQkKuD9P6OoCH
c5sk/0iAVrQ8s2TkxhRvB7+5/an1m7nbypk1QMiat4cocj6bisJ7DXqFFMO2
qpnDFmqhHwZrN4mgfwBZCeqc14LK7HMyq+WdBqjrBCD2mNRXtwGTasGluZuD
U5zwIdIlAsXmlRBGo2Ca7xG6FgAEoa/mHSa2YzAxbBqeHrdh9k7Bv3b5CsFr
ttK8UlNEOFSMZQp4DkXDMYKxXt9XF2h9hRcoOH3w55hJ/QI5V4ROJ4kWOU4/
JPgMhYj8Bc98Q+QTl9CzgZHUOAQ3zTeQu8dqaNbFy6lnEt6iyIRtKlFCgF6Z
ONj3oRhhkJwGC0gWhcMHI3rYStGBKWROu6ttD8PkVM7dDYXYKdauDqemhl2T
KZJ9Tq9+XMJEpZQY+VuvW22ixIQ4P2Sdpj2sb/kXO1rkJYR3tYKyzd2qHlx+
Lph9Lajs1PC5aLqgCnY7WCjudRIwamt35roCq0GQNokQ2rNJ+0UysYuu042y
4QopVLAYzVwJMW2IaeKxzk7TL9M6iMZLAG0b+2+SRzn57+htsEYwTOQPylsA
wUpPOLnUcRCvSLJhC6+1xyVb9F4/N/b7U6TgQVFQUVxRFNNIQ5jPtLAO8GDb
q++Akk7N3qXLHHvtJLjXM0JwrjepBzmaHcfijLKMDQJkZIYWx1T59qaKeYtX
BdTp7ssIQ+H5Z9z/DG2y17iCZtoAa9mIozGwI3EmBJ2GCQtbDzhK/LHQzum2
QpnyswNvdp8gLmA6lZQEF3XryXx93wFcCAKflFaac79LVCqp+1F3MXYyYQ3x
b/KAfpBrD1XmObPmVffzZOh+H7x1jt8mIYUi8jE4fCBhly/saR6jZ9RJPnTU
RLg1cdYq+sRe32mwDIZAJcg5o8ROCEl8qAL0GR84KGsfA3991OmE/o6hRbdC
98tYVBjy+j3eXRJ2QZt3VBpRXeA6rRTs7HNvhRd5ASIAloD4BZwIERqHWSVO
ie697JRlLwqsmoWabCRUl15RIlWSyQPa8/iy7+vRmakEHqVCUEl0MRUgwbAP
+kfsAorJI49bpok+m78eeSgrzen6DyO4fLgRm+TcKn1kZbU7oWG+AC3p3GKJ
JdoJT71ISy2sysBkozyT9hSjUKjd969xJ8tzZeISZaOXLvkX5rWxJX3TTr3B
wdVH15y55bREV/1oAPgZjw4oEsZh0kE/lViWKpUEzdAb6Jri3XfDq1Qyfw1z
yaufQYom61lSSsoqasTsqRTPfiZwv+2O1C7wzAN5NRCq6mmzsnRzVKtFSAgm
m9KxktRKZ7d9Rfrrd26isuhgLWUK+Q/PgLGyUsTijFlg9ga4LhBCtLhTInrP
tnYEk3wTLKpsd7NP+8TbX81cUrBdBYBUjilgORReSQji4FPMcrcq8eSTyeag
VpK5tFwLXo1D+bhQ99PphlPDfDykm4cJI4n5ttkC4lAiccxkZ4pFA9fupgXG
q5FdcIib0asB0JVPphZUfJV7g6Au/Qqd5osx+LnrMFo8zu+u/09DJljacr/p
9Zk8qw1/4O1e2asXx4SALlLAOg8rdUqdVBQTCbxctMw4kEtauiFAr7FMWhaJ
lc6MLu1vJbLV61RHmebbuY82DTbJ2Fv7Qk4HJnXX5rSQcsKRHazSfFrL1djb
ymL2DjkyDMvdBuZUKlT8wGO5hvoiCXg+aO81wWFEk5eoLdCuSeFY8zH+/6NU
F/xSeJ6jib9X6kveJxKVYiurjbBLSjB55Z4oxTtLmsJ4rqGTresM1pPJxcLe
8scADHohWPGA9oG/I6KpBDjMFNcfpSCDIrOVyWRnvxsSUZbL/LRPo2Z6VRN5
RRoE0fkQvRPh82sJT2DYnLx7R5kKIA7ALSV601hjr3gvmihfdHXEyyqPwQ/K
A+ydIxIJFCkYA1LRYyJM+ssX+1xJwSqYU8R+u+yu3z+S1WaNkcB6e1j5Mir0
aRn76KiBeuojYS2JUiP36hRltaELhuxshjZ1OhUHVRvxsgR6oYnsHbWAMxlC
qlQKcACxbWVPfGrVeA3Wt/2ohKqNCgUfu7SgowPK+pb43GviZqMYI88RTwK8
vR8NeQiA4yEKyL9MZ6TCx9loM/ThfGIwoJNeTOuLUyQJuPUNGmyraSiPoQIA
4FwL8XvdPRxMMGSY7NFD5Cpk9TkrjOBQsy5oz1fWhLIt8s+96QzQ2JgdB5l6
jDOXP+0eenVzEy+2ewy90OQ+Kb8vODNzYz0dhqJLQb3A1DA0P6S1XBD4aui+
dOyI9q1KU2QvyYocmCFAnpZLFoOrCi/+Zx5uhLb2thcmrh4EyIrfqbq1Xl1Y
MgdXFl5e4LdOhiYNGmfJSL23C4f+xMTt/tJVAbbfzlg4M2f2qjhWGebOC5UC
8E+JqD7rec7sqWG9xkhjgpdUh1bQBw3rgTKJtVZElTw5Zst1lFaP6TAPlqw0
FiDgUFd7Nb+FWOI9Yw38/MTBtBCCQfPNZC5uK1sCUyC2vGfbHNpGLEDvEk3n
o57iDJA2g4nTfmcVv0kqJIT0+XvISVNvkSQV2xoQeAzCR1WbhxBGoPMx9hUz
IvrfiN/qq2N9bt80qTtNFkJK+U+XakCvbAzP1ZNZfAGChtR9rMf84Lkj7hrD
Wpp4e9dA68AJuiagBfDp1alYYRCUxULgsY7uuqtl8TtjYCyKVTCEaHqKxnaa
cdlLAKd8ZdBQx/k7ZLGwbYytdEhI9v5dSy8KRSy1RcblbrCZnOZVINqAd5xa
8DfQRQp98dQYx9DNCg8rXP3Iof0x1fayxj+orFbx+55DVDoB/BLFGnuO7blP
WSNTb8racT64rEZzr8ufIyJaxmGGx6xtgywmecExGbS6bH5fkM6L0Pmcws0a
rfhuNSbUmsxdBos3sLo5bhwJJDBZwetxL9OjNBJQcTin17Z6Sggi/9W/HJRA
Z2qRto1slGtpwQbSwYON7LKT6OsRLUTAIyhngQmHNsW2J5Ny5L7YIz0gL3q7
AAPnTtO//EnbViYJFJb2cE5gW9+/UqJnwlyPAeLB6ndK+/Ou+GF9oLTUNa2l
Gl2xZZ/Iqluf1xD39QhTbi1ZatbJ3QATAhYXHeWCg4V6cz7ky4xFVntPX8Nh
g2aveSl5IO6jbFGoToybpLGYmJIaAbuyFNXrN9j79EFddWepnVkn15gwzSTQ
l+7B3xVMS9GWPrkR5TbPN3J8JhSx+qaHGDwUk7y7Ar5HcJx9xtziTjFpQArQ
vH43lVhb5f5ZJBQEaAGw2vdNIrYEQ9Pg6muaIcIEDD1cB2IWouh/RoMf+ssy
qQD9ucI4K8z5qp0vM9A0uHqn5hpBKJ4ttQ0SZBCKO2Hu3qawmDsWKWt4n+8P
6WpAOE6qiwjO1/I6ThSs0A3O7auXvacSaWgF7hfXFs41FFJ45kgeY7PJtfZp
iDK1ssPbH9JHqwXJ5vVUoX6CCPfxEKXJ1D+Y23ZtLOUHkA9I0VH5bb9rz0fS
pdhv4/vGMc7cqmopweS05cgKR54Q4DtTWuOXOP/i7ilpJrbzl2TKgRwzwnge
xz47IfDc+KQReOCiTmcCdYMKoQYQj5YCfQIVtfmbLAZ5O2LCbElskq5gZ/zT
s5PP5lGW1lueiiabY5Cihm4/GpDnhZe2D+FECSzwoL+sywODczAvIMTJ3qMZ
jTBj4vZDTUcqJ00DjNqwdGtwhrXy8cVq1OZ1KHEQVrE6jpwKOHCM7HWyGDQr
JsB6636eAaONXOgqsQmHxz6wXF6MKg3dIlQO05s+4H3Ofn9UB4fESxbAzLey
nMIPGIXG1MaFD+qxkCuMExXjHgAkIaupmA1ytj9NnJF1RNafupX1ysBGxATr
AZH2TZor1R+V+eUdQUz9r6JclQ0ESHBMGbTA7Ar983itgVB8BN50ydV/5xkZ
RPkGXBxjo4sqdYd/FU//QQYB2TFl2Tb+mOmhOOVR9vtlhVbf7rOhfQrYdO6g
x1NtZ01BbZ27DvOQQzLKvArIh4se4zkthGOf1+lw+z3vTYSdMBowpW3zeORH
HLDx2+0L9287wELOOXDqv+gt7PHgGJvamrGMB/uFazWj8R96D0+6oO7LohsY
UBVFiHbjqG5/P/h6uMoobFLDtftN/tv2cURugReH8uwnCf7jmIdh3oC9+xsh
g4nu/F2UqkKRH0tgZ644AHuf8xYpNAPywdZvoH81GZUJSlcmqbUpb0K3B+8j
Uf38Mb4Cc/qqNFONi3ya3nMRf2uQ89ZsyvijD04PcKJBWW9YRFKEPaOk1Gge
b/Mrzft/gZbt3FsRVcCnLJP14UFgISd1l+5g0oR63oUEheqtHvBDlDkFpqiU
r9xYTBdoD7b1ob9aMEERYGvSthFqyYq869pJS45GcX1UrOniV1CV/IasI7yL
8Q8ik0taG4SDDjNRNvcdEeoQECZwNkIzPLFeEWYQjl1cTO3DvO2BvigURRqQ
mCM10EwyP9s+1kq9T5tFJSwmPHBIkE1vfGsckgK5GZmFzUuzUKmdJ9eI1gNn
mjgYS2TL91bTJPkys8s/7gqv0Iea1wnaWWxN3+LtkwEB3d5GjEfrhkNk34iI
P2AKBg1uB1zEqEaodeNfQv6oH7eCVKARed+DYt80LXqp3Zq/t4An2Edbc3zo
LfP0rHdsLW+zDvv4rURulj6blXz+yFGj0ibHjYqjLUcUn9ODe+021EA/hiC9
wsTd2YimfMmTfIWpX3xGdJsPCAG1vQhrXJLmeqas1DGzhPXkM5jGSeiMqfYy
S4GkL7bfRHU2Kvp2soACj6YYRTSi/izJEdgJ7BwO+XT3Yis8xlcKGTzy3w6c
egbgf+tlDehUdg/xp47WMJQpflsRilipfr0ejMO+rF5fX4zDTw7gXVpBuxu0
MnSNEfdAD0iBXvfv9qKq0H/TmCeRMIc16Wvg+D+z4kBUUdauqfH08lVS+g0L
SrKgmWZYU+eAa1DZUjPDf2jLd3Xf5N1TyV4FtHVpTnSGtQLHcWKUz1PXfUrP
zEC0KsYfObqFAuJ+mkB3v0b/aLjVFZgR1jXzvuDoyfQS9YkUdm6CIiHwMz6q
2ZpjDh2eDoeMiBa4tdTGn5iY1FmIr9aOKrmFPxFH7cNxsuS52hsF/5SfutC4
Ounftrvbu29/IZ9qcusoMX/bHBX1mullVds4EBdnmP0NWDLzP8FPekTpU/Pj
rHBZzvt7YnGDk4fraoiAs7h02dbP1MIiC0IzZ//oCJ3QtoWg6gSM3ur3R1JX
zfDtITRsubVr+Mv4rnieaTYJCYgulKT9QxoXmo+CP8JyaV/OhMzbaiDJdpTD
acSTfCh/Oq2n1Gevt2aa0n/cO8Xx/sMc9AsDuOQ/REsa33wOfnwk1686XAjB
1erXqJcb4gYUo0FVUcKcY6CIr0A2RIGodr3OMcaJdwa3k6OqIt7ILZ9bOheu
XMNvJItkZzZ57RUg/Z5OgoISJvioukfhJKC3UrYocUEaI1039rQJp+UwVcWk
fsmfRFRgntYCTs/L8JgTGAtAlKp9w0gbZ/a/xmmZVN4r9DUbAURZFDzhweaw
uJH7UA0YL36AlYNivmSNVFYllhaZqCOcj95m6Ljv7p++z5CIBhpKQNrCnBUP
GBWCp8MMuY1rZxD/Yozo1MMezvkvHd1pBmq7y+AYFQ5Q3J/sgzgXtKYR4aBm
zO5u58nB52b+XPZ8tSf1rkbDomwV9+kS04F6Wjh1MEga4xUR4tf8VZ+kVLYM
cCDN7to9yqQ/3zCn74KtFuC7ZD30hbcJo6AbU+aHfqDP42vwClXVmusBKCt9
AIEuQtdziSt+S5jkpNsgNNUcyycCF+FVC9Eojox/dtU6XXnHjrSgyCMh5x8m
DuiUB9lO0DLDIXYPeJ1XlHUMiVFXkI7GHaabSF9/IIrC5i7uswKsPnix7AQ7
FqxKbjRQqkY1VvidPoMC8J/QwgIirwSBoI2B89dPH76hb3VVQI65TGRjfDyI
Vzzemr+tHvqDV2PRmneINhqPD9SiGe4CNMKtf5MMoVb808EQ7Jrh+KjobpYS
HE8y2b3JuYxLyDDZvY/hnBDdHffIsPZXtJiDrzbqS75cVeW5Wuuej2edH40H
aZa17isEevQkDT6nl7DLKfpXJzYpTMoFbjTVZ7L34gZSaiO1LNzzLdkabdXr
T7DhO6QWp3Odx1mQi3Aq9lAfZx8ihteoQ1k3z6VBOM38V2cx5rnx6ooGWM+D
+9xr/jqETg4mvmrGQ9Cr2r8YgPwmIRM4c79Tx9oloKvD9A/sMd2gQ2QQXQut
sm56DmvIMFqL2Foy3Sc9BTdfFCDFX1gDvXRQ4HSASgGzxCOlmUlYDps+OJPg
Vks4BSQHfV47rrWG423hNYXJZrzCFNnl+R/ex1jBnU8jHRZAy31MmPQgmYgp
vkHfdvw6t5hra55DbbQyLJ8gxHj3synaYsTNHDHXtsbX0EkIBcwLEFuhqBF9
L1x0SyqnFjESZqmgpWCUbCf8YZhrm24P0JV0C66vAhNmfrAuoZGgl45jj1AI
b4jJYGnN/J9V/2FNb5LxDTxx6HPFj9vyArqEesDwVbOILCP6juK7Nr7Bsilk
Zj6gNXro7iH0RHfeBdoCB6uXrgVFqf5AQBIzAeHi7m1eVk23XVVSgUNsOsim
yexc6KYPxk/Tm3zqHGC6oIzQChJiSG+8dgAwky8FE7u8OsjL3KJCpJ4k2uI0
TMvGEKHROY9X5m0eixjUfTpmd4VsLSbvWbgeAGYz/BKTQIy+kLdvY+/Cey6m
L8ZqgCZKRV3T0cPr6NlKA7D+Ew2ylwqIa96LDr5Yvtq2m1eV42r1AiUrRSgm
vPqNKs/zQ0R9mbZtBz0riT0UgG+MElhf0VPB6X5jscLF8O2Knurr51EGebd0
IyWWV4lDF/WubuVZkT/O/D7geg7QY2CUYq41FfSaEqZCZzLMAkhA9PtWAYZT
0G/MyFnZUI3PXq/vxR0yt+e/x4tvwIFSVdlJohDImq1DwD5YDOxHfW6vVz7i
GnpWbR7lkCSVnitxxUARt9m2scXfQe5za+keLIHIkmoNqGq6QYpgGnIYxAMr
8tIsqmNkjg8IgORIEIU7/f3rMnpXTgq/Pe7xddk0pzcRTBocJBZKbX54i8yC
yhogNB+40m//V0aG15dr0O1mWWNXdsF5LyKGuuVdlEA4D/12hj88K9rYmC1T
iIC6vh1ubyUS2E0ZDm9tiU77xFkzeQcoI/7+5vYlmrTHYZqmW6rNLVfsnSq7
r/1byaYKRX1FukfE7IbrM6VQvKA9FqDjmB3Z83LV9yGJJXWBmwLkGQ9qd50D
jMMgeCO3r/U75caGXamzwwuC+0hoqZ9EWRqtMBo6fsjDQsMbSTU/Oa9ZYkfz
docgxTt3X+vrpzjRsv8FhZ3M3ODlXbAzb5QdLEvWcWbySYQLN8XCK99Egt6z
3P/cGHGBBaYV8eV9J0FOlJaza8hI7Y5khaMwdCLBmjFr0XHkSJRST3sibQe/
uKXdDuEsezn/bAJDiazWH+LPVI6DNAoMmswDRaO2PAtAw628rDnLcX68U0Vq
6ah2hfcNN7RLqhdLcZlXAJqnrDpjr+oYDUaYsQBqR5VsELUJ4sMu60DC6rT0
lz2UM7u+MxiQAPmDJERCB5llS6QfJzcUDEzFZQdGL5JvvQ/D9aBVK0Xu3iOx
omOrQ0Rwr1tJIF8A+kiCxvKB2NoDWU1oYjMAXjMVWj/7Xm3Gqgo9IddzhzXg
Uv+q/LtCj45XcsCoQhbQIvMphyABBMfVY9T/cVq2/gHI8QqBtUvL2WvzydlU
c7VTMSjbCbYUveDZX1oVj4ls4NMfy11rkpbjnCIRIcjAHnqk4TYEbiVWmT89
iOZlQ2sayQfGLZVf+Ab4SDXVLJhR9AJvjq8XNB/EjP+mzgB+ITQwCdjgYWBe
60qK7DsRv237JLzDwUsyCgabLG4CFYpu9OCUpzixjVhG06TS5g88tdgLuOX5
iKifOwG3qhIGIuN3lgPVXU22KwSzKUXz9moRkRfgZxu8UsI8LZ7S4qjgL4DT
jseSTcTbHYvKG/VG5/YCwo7rZ30Is36vCyWHeIBFeKezyEQoxkeCBkuzTFe3
ma8xlzj+Xw0fl95vVmBZJE6xirsRJhqmTIi1J4bZQFFV83gnS+7mUo602b51
O09vYVsOh8UGRKPwEWRWfcu4IE2dyV67hVsx+Z0jze45nPFJo6ybGlwBVdQw
uZGGLAoJjg5X38lhmONPR1V17ffUzIwWmHCFjMSG9teJ/SNCTOv1cC5pLDs6
iIdhLVHEFb5PTXirHK0o4G2Y3fDKRW+ouAyOB/inBJc+GvD0XjfVxJJCwlYM
1RXBz5Kcn4BHn+r5q7YeZHYGbjAW6FJeT9ZqBk5/h9+/ba9swIS/uGPyEuYw
TsFx94ax6Is2QGuv52nzQu/vl02G+vRD4hEYJ8i+ya/BDVnohk4EyU/ifWU5
U0+oZtFoCI78b3zQF1xSOCtyEjXbXqKvl6lauF2iaUZs3TZZkB25eVXz7kZ0
tGUoYj+mEJuclwEV088BhM9vOdCMKMAj6D+lTzVT7aoBd60ZoK5lGZhNj48h
VpiXnntiVA1P9lqTe8qikjk+wy7y0uc+xXdMHTprvmEcbrUkG2LVQvQVONsn
BSigZOdj49qh7ZpKls5QICK50Xp5ECUyMjRkEe6CLnG7nJkpJ7GPDT8xSirH
LFGVzJgw/kGUKs1HW6Xxnv5SMOtJHi7TdpcTOyxQkd6X2m31EdUMZ23b5aBG
3xWKEEYIKVcWHd4+fqYrI7IptEGdhgG/xsgj8EN+Y3ZlHIXK8uXQEOjrnhUL
3Rd19bDBWrhE312stWPh616nojTOGkGfcO6ap6CxEe1DOhwZGYHNWI3a2UUt
PAeDIzk1Bzl4G7rBuXwS0DQb/mbuG8s2JfSEX2hRhq1NOrLQKUYJD8yg6Nfr
HwRIUBWlCJIxdxmPL6XusNgm13B4MKpdWOYG573/PRb1XvSCwZWYAvDQ+q9e
CvT/qTlbNic+YALMTnfUNj9GoxCyqIy/KcKp1VNRhZQW33RJ4vBsWAqECmhj
VWyL6lZ+oFFOFH958cGKBQcw0NI9kNgZfpQlOqBLJ05gf/+vEgFzUnjuknLQ
77p7vlw0WTBV2qiE4UaDqxNt8JdaNjBzmZj0pxu8CRgUw4jFkzq4F4q5PxD7
Ew4MpG4fenEhVs3SjFRjKeEDKYNzdyWyTPtRcyYk/Y/no9AlD50Mopa+cavX
q3fxzTH+cus4R1PfFkePcAfuVky72uW1vVQDSXl/j2lWJ9QS5WOQgnoFZ5bF
eGa7nW4pTEI7uh/f5S1KBoAvU+hyVNXjFGsvc1ParcWfiKV+maXmRvX+KQYb
mMxeNKga5vCQVmQmbKB+hfNuT2/OBcSQBb4abfnuL3+W8KkfjSWYa+PVB2c5
2bohqy9jLxjFaN/oOLVXAe12RUXebU5YdSamgPtsWz1JVwUr5RVERPdEFbab
AB9oEZoVzdk3/A6CjBnKDFJvFkiK6LRAhRCOMuOD0DKyLmTvqE5GvUaRKDq4
veYeDj4db79u99GUtCm1K1KXGXHtCd/OXKGwRsfhuJaOOeexf6F4oFIT4HJ/
4bUlwNcAYm2LU/0zZiZuZnicvyLYza58Xnx5yC5jOfQqE82VrYE+6RO6pJEp
msV1GbXWwuwxNXoUM/CQi0qQ0zXKyyblFExdTSE0qC9oX8ikws1WLcjBe4Tg
2Y2bE/pFHGgRxVgw4N3f2FrJCjFhFqXtk2eTOsgW5u7kAat+G0NQGX6rruja
aLiQHvvLhjwWJicIXXDTMQ6mghaQFt7qfbvH3AlmzKUAwC6dIEZAhuInkerd
+23qo8elWuu6klv2nKjvjOExDrrBEJFdiQ3Rs9An8Boi2yDttx2sQKvB3nFQ
TOenn8DMS/aGgrYwY+Xv3mg4W95gHXCxXjZaySKwJG0x0WOAGj6jon4VKlSl
sqrTu2B4FtkV1gX2cXmHyeNfNFDoxfwEoCLvYJVTSGy5Q6xn+ENEa0abRsMn
E7NznsaFAObqBLJ/rIhOfyiDYQYP0y9NOfbq6q4tuUtrvQ/CZTx6zeKk359w
/ITi20V3m0Ec2m6zwZIIkkrnzWe9EtyStnM6Rabu43LvZcerCnJ29xtVO/Qn
TUkVuNiSZ5ZEQ2aqTEjDqXSk/hz0rZfTYmNogOuBirXwUeqDn//aGWY/w7IJ
a/B1VgnglKTQET98Uy7wlcvo7N8r8MLQqOn4nF/ro5E68OkYskufob3Ahmtm
A8cvCEPG1Rvo84K6wHqA9FzGgswHDDc4JO3r0WA4c1Za9M8794z4amfsb05q
So9hAGtMeGf4Smp8K/UMF9pO3yz1R2ogD/5shc4bizf2adXTzKE0Pw3C2ufx
iYRN/XPZv/svAC+PeX8DvtNyGY1GyxM8CUq6PVvJi05ZtXrgFafbA+7SO4UC
aVVBtZ8NfM42yC5NQxc/i9oL625mhqPyh+2Zu4hiFcUvkA9TQa9slVDpHNMT
7BCCOAS8nn4WTO8wHNR4DDekp4JsBg1k21ybnD66Q8ag6KrnVGsanI2KSvNB
0f9AVRF7YENsLjcuTG0V/v6e/oWXSbAuj7jUwvP9nBeIu1t5QLtqErr2hII6
f/eF+/ecfNM6jy1ewu8PUeTTKzbqMiBgy45trbqADLxcmMIiV2/d9zC7mqGY
VtS36nDogXPMVWpeJUMEADLBjr5SBc3cc2PTbxtgXEuolnB8xoamuROy4bMJ
Zbe7yX+Z5ljhjPbIBnVjt+7B5lf7EAsdfVjOVaJMLyG2GXXYnlrITTBsfRSp
VkmKrf4BvgjaRFPQLJSPWeceNCvLiMEOuxRCR9aCxzVRg19k8kbRSQqgN6zw
QjGIbYakH+8qSe3SL5bX3YngfXg69gFL5+H/l6xMmGyKqGTyTPYVINDI95q+
pXPWmjCLzM5ssnFuyPcoK8Njh067nsQXNMzP+hzzp79ZI9vOf1vLB0qcHRFe
ZqY90crT1P/1h6cp8i9YTTpLdAneJ6DHOiZEu3GMmvXccC+JwvSzEiVetkZ7
8Ois2z4VRMseja8fwpp/fDQWbj0GCse8XVC9XhdVzDX6qAK4lbDQEFDl6Yp0
MLb2uk58fM8Di6PPvXzMmtg+nisrp4rwtG3znCowRIJxvGiUd81t60vt48UO
WzvK7enQY6H6Jvc/dm/MjtHnKo7Odxosf0E9A8E7uzPfQX3dk8nOX/tS0n8k
W8VVF6ejTX4RPm5yBeBnXPpJk49XGkdL5SYyYVmwO5nwQaW2oPDPm3s5U3Zy
h/gjK5Rj/bS/tgtfjkekDvXqCt/UzMXyVUcdIBexdx8Q6p+fhDfdXXyhCIAZ
Vy1t9XzYvETufeDeet7qMFQF75ej000nJfN6szNsFFnitmlX8RF2P7QNrYKX
hSOyT0hisSAGqeE9Q7jkE5dfCLth6kQa1lJfaOYrtgIKXzNbGlx3hALPU+9m
9UKBJIwajbbUxJFO5eYErt3cd6X/1+l2lcH36TKIPHOVjxZkgRcK4p92S2oK
iMmrvkgUVC0VIJmxlSHAESgNAyka8X63DsbeTp89a8cW+VRlaKDWb0nMPmB5
09kELJyLm4eIXLLZXq2MyPCJAmwix18Kkx2yBD4mbxwk3A+/IfRzOXVdj0g3
K8p1/I5xkJ4FEuUeiTJEoz3AvkaZUbKWA2FHcyeZip2TIv22gtjsZ5i0mLtM
0P6gJwQHWONcDyOKc+D6vGje6U8v+c8ITqbMiyC/fdh6ggBg2EIjjAnpMypk
1yLLcslhK6MaJlTLDS/SMBeaVGTfuDXiu2wOgkqIQXGClmzQX28pSxwdk3HE
pD3688Wom/dRpc00zZKmBZ2tW0uMqth1ElIr9lXmCShixfkuVvpK8+UHNT+i
z3z3+OhvMZKCZSfNevH30Jd8V/JDCaLkmDnMrp8XDABIJ4zuo/U63riyhHfc
MbDI79EZvas/R1KfmJX12oaYWtrmqJv/TudQqWozH0HYumuQyyEQbdKnYEB6
CR+OQUpIfvLsGIEDyz7rK9+PShw4leFuYJGgBYKhIGsqQlwWqsSM80n6Dee0
hfC/vibzZaZqOgoRA1IjLKjbbBaP0HCVDnFBRqk+WluGpmhslerPS0WzfsOy
C0dDoYc2YpFtwCqoije7qlnh+4L+nryWn/9XdINpxd9/w+x3sXqg+7LoMDSX
/ytltr8h0cVVPNSMiTUfxB0OlNRGgkJQq16nsgLGDOs/JCTwFNnNfWpcQaG0
wuqpBqcbNy1XSld3ZNECGgfcTFTX6Ndnty2Kie99PphKlKbOkxUQ3TelkgY+
/taF7a7ZOWOZXkdHSQ5BYywm98vMBaLpqxiLcHWzfZVcbFh7wXHsjg3bqXQV
OGo4AFu6psOeBwXlF6gr2VBeWXOcVwYskmx0S/n7WUxqV4gmenPYgwexVvbv
RukRJ+/OKIkSPrFZ9Z8m0nlxfQ0GcfNWYMiAwvCPJW46cQr8zv+6GTsx+A/P
GafvVf6FUGI2LebGXQ1zhW7zZqvVmI96TvaOSZWxJfeUT2LPPz7xcZ1DVZZw
2nAuAsyDXWvTvUNsiFhRKUv8eICzWDzFRm88nhCE8uIwHFtZ0udYnRy8XCEw
K2wHAjVNzTDnFu/Rtbjg9NE85+B8qnUFlTrbfGE24UTnn0kQ40KQpeb8O2+v
1kxwLTMCLOaVrAbQRT+Ie2ORTKBL2TqFv9fHP1MWWWTf+9yZYDohNigy1LiP
DLntjHBRnXvc6WpRxxd6+NoCUYBHrCiSUzaREQiFmX60h4RQUHIzX70edAjz
IwpK2IKLe7tJBXKXkN6YjncxETChyiuc9ZFMthLjJ+x3WzpW1b3X9CPYy/pt
KYbJg5gmAZcJ0i4pX9TEXFRRYkV7bOaDcAKIRodAR/ZintKemjQ2Wo6YLLzK
S89Eby7PsqCrctJVfl/hmQAozOehCGKozMkvGbfICnbn6iGNlIXLoyMno9G+
2PxGRXNJJE2GXdjWsgb+/SL3lYeBfaiVX0tAzFnjZd1TZ8ZeRN0ZXmBcc6W5
n//m3YbIZAcZe3/xtubA1B/jZZndh3hFcWugm5Bk/LbUkleL1JOMkCrlLkco
c7tRwGRVouHMU+tU/FYuHsNUv8dyZxSLYVXvn2oq72OzLsoBZ18he7oJ8xSs
QwYZNGLRRacIVUQlODMZ/rN+EqRhuWzBG5J2kwXa9X50k/1+q0NtRINgSEca
bWGFBcneomUioOIMNs8LFppZR3ctt9+iYHrW6Ek1FRPJk7iRx7GCkR/tBtoS
HMOMOt6dfBHmnerFoGqC+IhOQh7GBP8mk78+SnOja4WgF1VtMKN2JO2Dj+9q
5FRRopT5fvLzXCoowktvoEsTL60mmDWX4Kow9uMGnt2TjHVMlbQEjnhN/eQR
cnMlzhGww5NhJzcJreIw6On3m3LNpEaiyCogtgJ4nPC1CykWMXXxBvrJhkui
eFvI3U2kGu0WWte9veXU0gU8zEuIwdghYUwPoJVBnU67mjJmhKKN/T+xbuFw
s48ssOYocvnG6b3aXvsu0iUWwdYh/atTPVN7/WAbOtxiVEXcyfvtsvfdufly
YNzgFpLFFvnhvbO7RJIsaLd7QxgeMgmPENpDgdT3Bp6dYNNXF0YAUnA4txuv
G89zvymLEYfaX5ZXK0xuJW53tg0HMxra+L3D8xwxK4bqZscUVfU9sqvUAKBr
Fa4CrnNMNhXxSN/+oDGnDT0O4St5rrGTyMgwyLQn0DXJv88ydVYV7lHLIkjY
pSIZCLy4TO3DFNjjEpZCEjHgvGjazXOhDtlCB/YuUip1XOvq9whuFJAlGms7
kYHXSROl6mODRFfDEj7eqffWAiPbzgyqKYpFTFbQjUoBHNmOgnnEOOo3LeXM
eJAM8Sxw2xtckFdwKhYW5UJbsSq4O35v6d+MxJ3Bu9evZE4gpxfPMaatdTul
WV+2YKdi8WzMTeYu8o1dcEFAFHiZSazo4vqkKPkLwRrgE9T2mz4v/EkWC46G
283XbGeyutS7nB+dgnVd9uGFTI9UoEJDxge2haW7Ou8ClfJIZV0F/3be/d1R
8BZA9D1860vXKP+zlVTIhVfAnViyfjQgchne1t8NqccnGCzFR5z26MCSw71/
sr/g+L+whIkrYbD2jmEwueg2aHieZNeFxL/er63Si7ul14cYtbGlURcd1ctw
sdASf0EkHXPrArsPrvUnBb76ckxvjX3pzoxRpJ+SPFnju5A2EIuFPnS9CoVT
AaBOqiSDdI0kGq3sMVvDhEZE8ooILwV0h7oW8HcWS73KGlB2YgHWqwmaJaiD
thFC3GHtW/+ogutzjPO/lVf/6SIGRqQ6t0+Us/Yt4zXZtdHEbhmP7PJa6JrV
x1scXuphci9mK0FdYLhozCcEPLK4jLBPttv/Pe9Q8JNSE2MnsCB298K7lzMy
HUN0LOXQ8r2oPoQnVy9tZnJPWAhsmm0zTDrMFb/eRGH9wa0ac0r3fVLT7k3B
1MFp+mQNGnTYH4hftB4iF4R8TwQCFRiDClQEPoXd3lU1+6SZ66E+uxuJnGg2
WoQDLhvaHcPnH3c2MEM5+KUbIjVjNbtcTmPWynJyc4e2hvnOqelK0QTLUOtl
++aRyiYLPlwP8xvo40hi5pYVR8f8xmHqbGHizUVXf710sYp4tCtX8fjhKbHE
kbuNk5sYVWDmifrICcJ3Zbxxj5e5Gkd73NGsek8i34S4BsIte0bt7wLdlW73
4ujFLJ7/0dAu9jfG8stZcPBkGNbBiVybyLY+2ArytwWFzfoMiFgvjOFejugk
uwfYSxrML5I0ZglnGKRLCyUT1lAPXxEWL+qHI8siAkO7RlEjthKmzzhC6Ut9
QbbGhjOIoGS11/EJe6rXTLk/gQJS/Tz+dwt9xCxeeK7so59R55WsO2LpO3Zy
3gM8U7tgZ0pAIGxRqLdPuCQTQER4lMDgjjZ37mlogTnIiOLz3aOnwjNtDv5z
mtuWyKH7W7+sxY/9l8Sq70PSK1lRUHW4BL1ldPIwCvOheoaT3LC/J4XKqgy+
earvokjbpbXIk818+lygXKHud/VQa/5E+Fj8PHlyj/QijIiC0SCSPN1eF+GL
RJGjlOSd8A9iSkmN8gcukq3pym4m47MfvxmF6HILwyo1po9JbG+W9GztbKzV
yxS+3xy4xTucwHCCdY+uXuHUmzuI6QVHNGQMlFoUeORZraT0wSnLI7cEsWjM
Hgwye+yl4mWMsRlE9zyFbEedHjssXZG0z7K+TXKn7fzQXs8Ug4zgU/lmQICj
txcKgCc5wAqXCcZaXXCL7Uivmrv+RAB+CB0T12mcNyMRUm3fH6uy+HTkK+H7
yQ3Brd2eSEgXyZ5/Kux9E4qWJ90em93Gs81E5BuB0S5ICOVw4VzjOGePq/qn
h+0MUJs0dI5u9DJXsFcVJz01SBmMx8XZiS/OArK8cdCJILp1GUxMo18j8ydx
x5eHxYFa4mmxLONB8ZVmn5YJ1JYPs1yzWumfsz3m4ByP6hHtMOtlsH82GvwJ
mze1urZfjjyGC/YycTlodBK2rg0k5TcdH4MxIZf21F6rmO6VmjW3SlStauXa
Fob0rUEAjBHXaYZ3WUWrBJrOROOjF+qp0JMEYXtj4VomgCLYqzLvaJbYk55z
/8NTm/gwQsKAGcKuUTY8YuW5IlzxZ8kjXCtWKEXJ/qEXysf77yGALV1qkyic
rH6K4wTbEwS2Fe600Sf+a2bpkK3xA3hJyTATFUADOFmtwvHmkbFfcVf/a78P
tYuAcOuUr7GSTNyOItXAD1erKnQjqAwooic6AoMOq7qekMDqqWqyv/txzsGY
/cx8DWe2mLn0yMlj8EfhAV5KCd8CYAcNk2bPI74rLblWfJpNFEFTSWnvQeGX
e1SZNOQhdr2NJUSzQkpsW1ff4L+FXnO8n6aVgOg1i66hLrBO33/2B55ncTXa
+rzWJNj6mD5g9Z5xLB/I4B+uE11cgTgO6zsKRsug5MTppkOaJlBglpAg2PTI
AXrExerwohaOgF0dWDSvL2ll2UUsd9eIUJt7ShDaWyJro79bwi/4aE1QG643
LjlMBq1LjSKfOBtL69HyN45nJxTZdKqbatfvZ6y1F54FyBrIH6pUNfdSu1Su
uaeM6ATyIF2O4pDQxkBw6I5V3FTBrkHuK5Jh41yqKjsfzPWLYM81dj5hsCXq
9TivE+mExaCGBaq7ry5vRCe3KxDLTZUIJfxubS0IGM3cLUVNipU7MspThE94
VgO8AxB8APQ31L7MYY6/CPsFCEjGZe0sWjkzHi+gc0ynuuxwc+Z8QM94wrri
OkZ1/CfnBbwkYNSiQwMfm5aEjnrnEYo+HcD2E3rGXW+DC0e3M1C/GU9F1kjj
AYU5WhCGhDyHc/scdP64t4xTjrgkH/Hfpn1ZDX+7PjNNhjxWDSBG5NsSOkV/
f6Vv4IIKUUVeqgjnEkLJI18P3MrRlGV9FNYUBjmXWdcTZx2oQ68F1E3cw48t
EIb79qO7RwpSnvKN0ZZ72tyzsYgQrFb1ylZcq8vbRo78PxyHQDeNxHMfaOsK
Cl59kiM+NxCd81U3QZdsgkAZPZZiOKxDxl06EQUyTE72eDGECoWjkLY2eJpg
8QpI8Y1EdfSQleSoCgUQ9TQ/HrOb0fJ1BYHpeA6gyqpcRF511nSVtSQIZnd+
fSTa34WOcpEeqOOChvLH+pov9DJ3fL0jDwRQALdMYGPmGHPLQdOkTYFFwQzJ
3/KbdBzKPIRSikBrUNA+iAezRMemJs5gdxj7hd7FC7bMbNb7nO/4R3uqOGzL
+qWIUL8jL6oSQZ46XICDfVZY5jr2cKNxEbu2A30J8PVw7SCfO03uofmDF7Q6
K6nD9RdQthg2bhF9qqN85YIRWz1/bQskMj9v8cBRPtFpiDNPYBHJ9oe6gtKO
z3ZxotUdwibWs22IosgPdyVXs2kVzG8edBgagmpu+tE4AHYZ2oYbrtdVuek9
MkP22e+Gy4hO88Tnbj8ANA+nO5COhUquuMdfT2685i2dFtg5I3JXhGPNRk/N
GoCVqTPVbrgQHJtM19dbxPTC++kbR7M3BHENwPa7VNCPHtKHJ5IN/aZto+dC
0C8Y7WcIH1B2ac9isTtYr0ytVa3ZR/IvfmuTwaBt2EEUVYPP/Bc+dzHJn1op
M3CQ6V70rGeAwyqUvJrijQR6NSIYEjN79nsdjkzW55ppEupt0HZfTrrkVI5V
rd4GJZPmxBfVsg6VYl5WGVf/iMJVYdSTPkUjldInrQw12/FOSH1d6NlXPsS3
u5u/+thAohIKszG14tJZFnkjQRX4qH1C+5Uda/uq4ckg4IIPQK2PX0xToDf5
rrcP62jP15ywWvHM8cT3SvaIW5+gDKXEOxb2Kl9i7tqvv1dFlnMXiT8blPuU
s0a90x7Ve+Np8fZqC3E7ldFJr9tep3qRV1UZTCAh4998LEPTs7NuFmPv5IXr
ONsR1OWuEOS/2SHljhprNaahBN7ehKIK0OnRWm+PyfPkdbwv9kJ9M2fzf4no
FopxlrO1WrRvj3HJalcX7D5lo0LoIQiNkEhx3ukSGeyMCe+zWNOgbbaK1syK
VBXNCGSdbRiJCRPCxMS29hvc7pq/Y2+k264pcDm+hRNgPM7uhWN+Slw1rPzA
Xn5V9K6JfLJxGqJo5ECrGntMVUzX5KUDeegUj39jQaA4G7lHxap6LfHU8IHI
aBOtC5Xq2KI7ISKHvnCfmW1+n2oo/DbKHt8Et+paLDi1boZbGOMSlcF9VOrB
1pJBb31juN44xLa93PWYi1dl7550nCtiR193/CsD2CdnwUIDwZAtQdb3ixpE
cYM5dwN64J05NPtWVTq7ewexgQpnX1GuvCpMIsWD/tSfEyggv8tclTq4GgLo
omWssdZHHoyetkh75N8UFZNLJ4qGqcHSqzioctPXXTc8RkHmG/WY0m0o2uEO
aRcsRPF4nxmwcm0YVzM1FBVy4Ky+hh8NxGVvg1vnWxv55R66qw0h5F15gTpo
u5n09R6aAiRdAjv/S480qqMkkF0GcCRSNemcM7jaf/6TC/jUVVP/lV3mU8gY
hdOoOiH3ih0zHKGA3h6dFVUQe1DxvcyIlAkRN2pdcYvSmtIzZacDxRksZQ6r
+8x96sHuxTNFjx0vroQJsIVe6tUBT+pgK3vyXX9jqYFvwuiCSAkMqi6xv9u1
fqtYO2phZhA1mo0sEacqGvP8vYE20TODeS0WuD1XB1Bvr+HEYEszYCwoRFk1
4j38S3YhpY5+jAruzjrdfqd4KXG/5moP/FKcCYTgTSxJUYJWix9jFxlW0czo
+/DayyZCYchZPaczBEYwCJdtXq6H6LRgC5Fw+qTmD9fVMQIP7e2ZSYX6oQ/w
f4cYRtOI+0xjyXJJDPIITF1w8peoxEd0CPl/EsYJv/QYtZXoBKr5ntzS6ecn
GuMQxy2mbXeO7OH38BeoIKXHtwmHmgY2TFgsgTpidTOpcJqWJU6YzCA9dQlM
h5RRmp0hDp/s/H7X9Zo+ThIgpbOqjd8pQmokkMawwXrKnyv060ATxj3aXOGt
/timmKmGeQZJfwF/2XGvIJQlELsYhhwRfuZnhDCr2mvuFGMR9oChdd8/ivUp
Wxb8M8VnOcm9K4DN9379vXm7o6hJS2bEMo/20rf3uiqta29FhpJkt/83+mK2
2uRQm1eS+7CNlD2Igtgl7wXbl8nN4OgUj0ya4GQW7IYu+jZlUUbuW2BsO6TW
3b0i0rwhFr3RrthXEXwoK9rMzGj4J+8j39VHOVI/SjO17sNoFPnVl4ZanImi
ZYfV9ci/pmgQi89Hir2BHmnQmxqm5rp2Zf+tHVnp9NYFcNu/cOKAe901dc5O
H/LfooS1A1kSZ07TdgQQ3KjP7jX4svu6TCIjdJNiMO7pJeo5/+9anHjTGORf
Sv8xcDyerCC4VnBPLgjrsy7NuhRIYj8VfXOBYMFmiSQP8EAanvBKDQF6zaZT
TsSjY4D5kRSPrC8P1afh7so1fctNy6ggpdc2gmzSuUqt2FmQBr6ysVnGsLaH
KcWnGQS73EKPtvdlxkXiMIRdOsuUhBpp269ms4Thr1NC7XZhZVrPvcG1v04g
AUasOjTk1pjRB7Wann8DnZKfYuNjfMKM+SZg+S7NoA3bKwj7/aa0ueOPuzU+
t6K6AtvqLwQ1xM5DZ3NrOa4eoqM1ZaMtewdSlVEiQtQbpjBVELn0hLFEQFnx
1UR4p5a3uNTDnJxg2LHWa2pqSYZPIianMK0R+RowTTCquHtkjp2CXwH7FF2H
V6IBciuYzgzZ+yCkt6p4HkTmzCcIag+gNEBq+GcQE64ImoDY58m8k8GYZvne
zcAdyHj3rW8U5iWqTjvjID0N4XaiPY3OSrwUCJMSWhWQkxoBZxwBarbetBeM
4BFGFc2SpTPPblinL+TEGdastCd2XtIbYCjdA2DmQdVkc/zg4GCDq4/TW5u/
nQXOaKyjYxfQk2h0m9Fo9TIfUbhq1C0XkL+5XMEMY/ldGWser7l8qtbqCyFq
UbfcnPz6Sz+iem42bASDgiBvTIeD0wEx8siiAomfY+TJH0+ArNQ/Lb83mAHk
J9BP2d8I5y5LC2JZ2To59kSdAkHdhRqBXFcj226X73R2MYbg9gfFhb7G30QY
HIVE+GKidkn4BxUVAdo57EmtZDSvkEBRMIiwgMZPLhOJnR5YQs+t8bBlOywa
ozlzyoTApcJ4Fhu5orsYYa1oHMGwbT00NGua/MhXRfrU+Y2I8iJo5hi/zyjJ
f/dYhVzLwT6rkmpswk2qRjnmII0+TkB2EirRNMSRwZT7L/jY8sex4cCFkY8n
OIF2Oa/cmm46OdVrc0MaXJyhDbAZjiqdw7BNrJXviJRNx8HqKm0d8QsiphAt
VjMmU86NVfUtYxxmmnOl2rbbwZwjuea2CKGzPzkgR9LRL+E4cqMWnLsyj1Jh
z7zWbvLdMuEOe7bYM0xjv5DxHF4kN/jBJ1SpT2n2LGmOdkHs0NCmp0P+XTGu
1GM63MsUsIdgZV8DcCoh/ehLlXOTm+q4hlnFOCs1fknZngL9qPXpTKOtozYQ
j5/sTVUgMIqllli0eonbZSdNLevGC4i4wVTWn/oXG2CGSOeI8GrePLvz/X4P
nZLVUF/Jnm0JfURfQ1srr7ZFTk6lAcbAxWEpbK5bEkbH6kq92Fb/7ncSxBMd
QVAfKYprUcLaev/XVLZKV+OiZ1V50l61M6XzjKrTUiBJ3CjOX+c2fSWOAMxM
ZqVvlKrqhNG2og/zRRV51RPljyb26KU9QK6Zg6tJFhy60JeFZ0vJI7yU1R0m
eQQXqvg9L7PrC4LCMFFHzvwTUqXFSJ8jhK9oFZuCiJb2bARyQn5eu92oe5L6
sEZxtuE6zEf3Dsx3Ippy2gjer5IYhTGYEVggg2e7d9fRMtYGtrDYUOnQmeEZ
d9d481Kh2ZRBK7Ac91bOm1KPkbVWfaaSQdP7xDSfr+NNqvmPhaldG8HYbNML
xR1Vgl3cKMs0Dsb+Juo2PnohKaJ5K4r9uSuc/9F8I+1t09x6BXrshzxxqsMw
ccTpJajOiSxjPbFA3bi9ovTfMCpQw1CLeI77H5+TrZpM0KvwYLFKvPiathSt
OGvJrFn/Ixp0Nuu+ccDQx0grQ1fJfkkiAGnTwvqGkxtW/k/csV3M681CSZpl
bWii2Qjus1D/jVjUzsJTVSBCjpZNLdCfWoHNNwYUMyGXfw1KLltO0DkizYTI
a7Hj0Q1CJHPQCj/gIdruAmpb6FWLl9mZXXYOBbFHPFi4VwRofXaTvojAr5EZ
E34LKMcwkfksi0Q3gHaWILQnxjFFh2kvnxS9psbpcOJeORDavgfNFv/BrBYN
4eLWdmyFrVzgCzBIH/OD0hXMncurNwGeFzS8kGX8eJYV5xYXOQ8LVHu7byRF
1nuWhROX96QXpfP5QAYuDIGOlvqWSvuryAWsz46nQnghAO8ABPuJvgJEgPDA
5ItME0bUFNMaKlW/CqE4sJNsLcYxtGPVzRs7Gvvs488Cwz4z3HYlFdEpNC3j
wl1OylgQR4fHC2ynMg7+RM7Po2Iwx2vbwJCBTjz7qTFIX4Oxyz44UbGtD3o+
srHR7ElCQPUzN+PHX5BU//HsThS6jjhth5Z10yKtOgdMdWSvIkzWrH8lHjG6
jmIQuYEt5HKBQNZAu22Rb11LN46rfyHPLezK2f6In0eI1GKEDg/qmFGy+qFf
ei8l4Eb414w9p4Y5BeoRTf/7+EMdyjX5GQZa2kNvBmovWvrG+85yR5aLthCY
AQwiOpf75RFw3EVZ4jl+KSG1l7X8YME93bbX9dZin6kBVK/hXDpOg0S8v55B
DEaxrF6dp4Ks4RF1/iyt/yo1SUdjCQeU3bvfdVZtnMhg9aLO6UENYaWVb+6+
8lthiu9a8QKf+mHqaaln7L8fmhps7RGcYcghSNCMPOfmUaEERHArtYVDG7c2
i6beCEErzUprKqnONKPWNaqsRKp7s5ck8Ibb3pZqOJNHROqNXWYRZ4BGHYvr
dEs559SSat6lWva1zYk4oxrrJhxUNw4sKzCYwzACjq+2rLrRhTRGyvcBhROk
5+cj6xmk8Mig9S6np7U3rhpA8+B28/jlbvAWfHdg21vAVNzitjyr/OQVRzFG
R5B9xtNjhYRIS3p4yR0nZO46aJZ8WP7Vd1oZjdB8hbSwrHPncm1CtRhhesWP
wA85WimhIttggcWvU0kEvwcJNZPURGONiu/qSWP4WuX97MlTSv8uUEYjXmHP
ktNry8EnCIQmmaLfcnI2SKLFDVkYe00uYEmAXI5HCZKr9zYH83sBUKK0sIdQ
3nYix8KLo9phR2DBfZ2LWq1m+xV5bysloJlHOcDLv99g0+7bQP/tfZ1PjAaH
PG8rush2ylsR/zS9hfnMd1MJnFOBtkVC4Woz1Eaif2/LDbPkRZGaWoeRBzgx
hjilrqKV9b7DBGTrV+qN8m9b3hV5jhJK5SF8+49/dptRT1KaQ18c0V7BrpP9
+JqtVj0TNQoNHknmOb37aVSe1uTVM+7U7tLYHiDYX3IC/B8JKGUqBILQS+PB
HOmCKeM8qMslTmJAXrMcJL8O55QeLoRf2iVcqK9iC0eFRwEMFX2zmNAJr+Vl
z95hEuU/n28OcxRxdl0LfJ5qg5rTrPImCL8grMil8f8bX/LkzVPITKQHlvPa
GjjuZfX34tNAlQR4pvXERjLqcuV4WIflLZxNIPpkkq4tD2wZJtqzhtER6u7N
4jy/NYLTnTts1zUvuJTD0R+I/KcLkZz1aBJYJlDZLhxzBovv/txHo4nbZQPc
EbsqeAn3E6wkiLK/hZ1dx5L8f1Iw2pYzT3pZsT9HIb73wGCzTyfYAnsnDH7Q
Gi3zL9RZ2P9+4n6mfhnb8lV41/LaXCoqRAbVP8sNl4goZxSK7GDa7yWvwcX7
pdXXLFR9+hM9sWIta+u4PcXm2Ypbu8VOTIuCCsHUyJixk/gPfQ30DMi4Dler
eTNbvkcOwQJfgsxFh24QwW8Ui1Pr80IOeXBib52Q0YaQ8DCtQW34DGVIMEQq
Zw070lWBQcJ9Sr84Viv3CTJG1Tgb7Zmz1blIlYX+Yl7oBrDkr/W8LxBPnWzX
wYBfggYyHcD7S3HGc0LQQArsoTO0kb6bz2ui+8Aw/bRIRcaf12ZkqxNZAIqI
syh8hkSxIHj8Y1LrK2dv3sdh48gCz58XR4pyzxPfeyNfENpQ7lyismOozMyQ
W3EZ9rhPhC0L8vzRWv2aFaotG9SUfJvc0GQJPi1RjJW7xzGEKctoAiK5/s6U
8jUwyDU9ZdWyLQZKpxOCMeF8vhmVDvZbdjUwNqFysycII114tQRdcBA/lXtp
/qQENa+PqRPUk0tDhC6mZOfTNd4e7uX+X7dE4kv5I8QucKmqe2QWEIuAKTd0
ZXxFr7HIoEr6qt2QzvMvfwiZ2fgs1iOcc+daDDiABEXQZfUJ5SQLJMuW7a7i
/MU4btj0IHdetcGcL9xei5qdx8mwofFV4dxeRDEkiKpdWwZnSSTYZkOYz30I
xweZ10tQmR9KVdE1GxFHWMBBWHXmvizKvahpS98nrJ30BFfpP9J/i0hF9CLR
RlCr012PWb77kH/QQRq1SzUuKPOVd+WicEk0AdHVVmNXLeXLPoP/bH/Zif16
RbD++ksONK6douwUBLFXy5TTXc8GwFss6G3RA7Eqic3EKsuOVPqtsauG5BBP
pbYfxeHOQ/fQ5EVmonlwUKipPEJklVQdslSrkcwpgOb7fEHvqV0zmAU2k7/O
SU7c2ItKQ8kMgH8cbAbC7YApwU7wrVahZLx6jtELgAHDlvCDLJU1h62gCguQ
85Q8a3/Zvz09JcW+2X2q7xz/Us4+oVgkyaU1FQtUvIusjtFTatmWHXDrAC0u
u7hX1elZQY0CxC2Ei5crp7TyFNgsRBw4tux4gHgvEdkTghIHThZOALjM81rC
+FiO0jvvYkIgifXTUsulnhkYB/L76GS/+LhTfQr4lmBHsk2CcehRm1UCvLmt
Nzl1HZmDu+r5VzBuTo7vdQh02uUhnnakbaPteoSGNmXtOap3O0KeLL5pbTzK
nRn5LTsLnNRnKfQeQtkRiFNJF51fm0HmfsecR/7SgTG3WGW4KlaDszOKHnEh
Ip1VtbVx63rpgg+D/uk6xBPawk2L53Z3xwl8xYnMDt87gaf0IWD5MxUJCsji
PfN4P/LbPPoNRfuy3Iv6yUPqUdYIe6DgT9yU5Uc6ECq2n+FRb4xEwwy//una
0M9lJ5cA4kYnDRnwDIfZXWGDLw+xfT9MYrFaJFATMBymiuhe1mW5KCOPMt81
chjFa+WPCLBA4tvSb/9rgBGTrIVLHBnL0+J0ObEMHi4h3KrwB3C27Jsq+vim
Yo/R7nInehugYRMRUQYeGCXCXPk0yH7HME8QEmp14rEFlUdZOM7yvBK8sddu
fwo7Hx81oVyxT4NkyH0Vi7oytZHrvBCXLqyQRYXvNFsHEAXw+SsmIIKrYJoi
6LuUOEba2ESalNYsIJJy4eA1P4+msZJRO+3I0h9yx9EyXIvRk4g1HlMzCeYv
dr1xc4LvZXtSRXJ9X1DSHUHoxfL7i6UwS04YK50hki2nGPPTQa948zDeS+zi
EnGvM6N2uhIoxVdNExfDX2VYEgE97bICHSbFUWuhk/1BuWr5Vxx1kbrTUYx8
iMB1TCRCx7IkAXZo0G4YYmDFBY6xw0x+g6Phy7VNswbtyhurGSo9guflxmTK
Ify1Fe3Rknhrha2kCSUV6jDyT0hOglhOe7fVqTuPPvwMvQ8Z5hc0QOHMwFP4
TmkVrKYtKXU5UmPSSrQMD03WE1o07fZ+iCsBESbnHjVyz8U61OuDIdXKC8ik
dC6Q29SdoUiXtyseMSridLqPO4hXvJMlLeINBhb+Z8QmlV77JLQWkVeXSh2s
g5S/t1WXz4KfI5zbT2adi8UXIYYlSj8oov8zPpov39hwflGuZ8o+7ex4RPH1
OHHadLCuh/NpUXsYePakGiKvo+19kJrAY7syguYhPOj1F47NfxH9cOPxUGlZ
b6PdFu0QXpwiQqPv38kDObNAXHegEKJdid+WuFmXxMOEb+MGh8oHV11rY7QV
aydEvYCcgl2/EPEy43u1n3AwrN0nXtsTLspg6m3pRm7nzJizssXvwEXKtIHk
pCe3GDGEt/bo6sf8j6JbowzhUlRWl3srOT6/0hQT077JKg7wSUKJd/hEFt3j
5IeLgxew8lPQP4hkL8q7dk4FayADsRQ42kgq6Yvd/fuqu014BDZAZN/w/X5I
lbd2ZwI7T8ptsymW3zWT0qtDZKDf8mDIuGuc675NpcaXD7rb98AEDyGP5bx1
7lfEqWg2GuTv7dfiD+kmo3hy7YFqXNa69NuG60yhS3RQFtrz5b6NtunbJTuI
uwOxm0VfbAM0TUbV+I5vXYRu7Orkj4kX5i/VssJ9IZHfrFvhr/1hOBpAY/Wd
Uvdbw0hiEo+oRsE8vYvg5G7ua6jixeTpvaugT/5D+Ffr+FH7ylEJCWhY2vf1
QmVByryqPJ/mnwje8jXqp4ls+vgFvvMUBsP6t2bAEaXCVpoDdfGiySZKug3y
ml847l1pvDTxUeHB5gyPMO3cc9HZaAkEW2EIY8zwgVpzTGP4Dd/t3e8jMsrR
0nqxklOpy76e5B865AyWzJQHKWcTlA1T7fy7M64pWdyV082PnKsZO+EfO8hg
NYzZRVY9e7t9vWdceZyrSaZsZjNjCkVIKE+82j8oBlCRhZma7AikecnUeiIV
KPvbDsCOIPE3v2Jg5xFMZlW08OOVuQD/Ye5jEdVzHoEKygeWHgXvMfJLeH3X
0+FwQHvgLM27tEgM6l6T/PtOfLBoYb7lZ2ppzGhLF99vXt1N4+HH65qBezHZ
cLKUM3fFLfnbwdZLr0jkXX+FNx8H2Oufe2UGIMygQ9xSrjlxOp/G7EE7zuyf
voXaeBMlfpF3ej4mgRsCPqALYXQqClIbtz1ipFTzY34awUwrcynYVG3O6l+p
UB9YEgKhxf41C8BM4SlbaujDi9JripXuGEVSbJXLklAbhLEMj5uuCq5Q3gBZ
1uc21GH3j6K6FIR3VF8SYDVYyBcY4qkjpl70zs/JEKNi72i8vQmD3jIOPERV
tLmsvrcUQ/mtZSQEIRasAz355OytgGQbfhKsw7tCLcr55Zo1ZRKnzN69H/qp
Z/oRBSTAhE15TK8JAxyj0qypptkpYDKbLFdx8ZwJ9kg2TCTRIoI8/Fo8rZU3
yEix8ijjcNW+/UrLdoFDyCmzQopKSvOjFG0B+Mz+AGS6YobRtn0k5iXddzat
M2gT7qDyiW+qtetZMS5arILjmJX0rFW0KPrClHVr7tiqwgQ+vEy9TopVwuXi
x/G09Ga0F4Q1dOD7iZIcve9VryfieSjuIYQT2wu6/KSNxp4JZpWPBDCr7sIn
zAR1O/MGEk3bcgr25eI/xpvs/KJfZyu/Ma4PJ+eoS6nh7RlZ6ERe7fZ4r+/B
f/rHF7rQ2TXDNtJO6+10yE+KDxKGXSHtOC8loj8o75FtOeA68+Dza7zMHiYO
ldpAPuMusXdD0rnY8H1I53pdFQ3inNd7QUNnTxesAi8P/y72ID7yN9QoYYUL
fpL0nV7IHSxy5Oh+mnxSKahXBKxMI0P1bH2CJQPUeiITLMlEC9UmJBDXxiGA
fQR01jL0kA7OfAjbD9cYSo+lid1on4s3NBk17DhXp806pyrisvYIiZaGU0F0
BfTRfBycAIGsSOrT3gzHuQvOl1WFdXEIK52v7k1HXmX+BtRtHy6LUgZehPCJ
6AIYc6dLwid1E2wlQpIuh/8/6VUdKR6XiVPLkrj0X9+STcX4qNYrOBwb2Ju3
o9xFfZmWHcNgY4T4zxUANfq0yR+31Z/ArTERG1uGKK9N/DOz7kq9yc1HAGf3
gbNq8guzZxY+hcA880HzSvv/N/Dowl2iCf1bG4rgxVn2uTeTehN4vlB+5CWT
KOEpBkJv7+OSKdu2fOL7JxJ18paKSyemsmVDYQce4jzJCZ7DLMzZtWFxPicG
UljP+4pb6+/U5FCCxVr4+st0LY9qGR1trAld0sW//L2+SFkRrhSf4ucxlvae
LOs20GNQ3+oflbIuzHh9asbGpFfqenEsPb7x2gvddRKAilpb5a9LQUsaQq/m
S/Dk0MJdCsw3KX8WYBADFK2oeJ4V8a+HAizKCQbaqwO79R90ICRdB4SqWRtQ
780QxzYeHZfrXnyAa+3Bpu/0LTUvWBLklIBdnYP6VgQwZanxCHAJec9v17JQ
nSzAG0LJ+yGKbv0AwUd6ikWB32PrA+iBmq8XDpNkx2Qy2fAzlRCo6pZwXz59
t/LzPKg/ddGhwiBykIP87VpZYN2sjyFm5TOwt9jxTNHv7CnkBLbHzSEOTHwN
QuugvcOyHRO+RErMfHqqWf9So96wiHRNbV0jpIj9U9m5ZVzhyy5m2dVe2Tk5
EaM1+q/Gt3f4mv2ORI21NnzC41H/DQUmmibP0TtFlsTia7G41/qPH0OtbOT0
QYT9EXdmCGRDbUQ25hLcR1XK9a/ePwUKxqABXRi2mKbmdIYIzjSm52wBvp8f
0kLwK84ZsR4YP7gk234dB90f6BHO/n+9wYgqC+ye5LHnFnSz+E7DOImliIfq
QRZjKSDmhXLQjg27iHSqYYa9nHntMv77P7ygni4MFE0g3ffJFLLfKw6s6r6f
ZDCaCi5iQTCVpem+Hdo4lW12CQtGFy6dIBz0myCgJ07czDBWWEXOM5vnOZFO
bSvN75eYTbRpO7Bgl3tXOzzLuzF2hjgvNfPbB81YmycE5BMOIiZGJwDevBoB
cG0KGP+cFwdrLzxwJh25NrLxAYpoRzeL6PqvCCJxmCzeiUeDQG/hRKDrnFbW
PKZ3VTtTbNijbIdzfgB1fNj+3b3KBgKxLEO3faZ1huFE1C4PecaHKkWttzqV
uR858OsHBsXPJiA/0mmDNF2/y2FUa4KcR6QKascDEWwQ254VePJC2xPYHqqP
CWMFx70gyI4LLRzsPL1zdqt2QUq1GEVQPGdTSDIdclMFo9eql0kMvYzHuUlT
Z08bI3hKar+xTxVE78IAbvYnUp+EOWDqrNmKrKlV8+UDLXfvmYpNMV1DqrWA
jbV0F9sAeAOKU/+gt8uv4PHP/wNtPuOPgVaAVRrDYSwiiumfOP3mbd8DmY42
B2qBzR1BIXgqs1ADVTwkSpl5mdpEz0X1R5OOJMmA1ozkmUNmbODSTLz2JAaK
i6mXQ62xRaZIgYBD4GWV6CLxLX4f1CgjN60FD8iNgYbCVyWUyWy97ripaW6d
mGPV1JXGDilB8a68KVb/OJaPtKVV/Djhjj+/pUPMBBzpqdbg9adhnDkN4vzu
lBS6c7draLGH2lTniPIgusjEngZD54kQVFrTEti6d+hu/IkGLX5kqq2ycGsz
mk4q1gy9MRcpBagCR1fudsprxA1hhpIF2Io26PZN+euVQGMsaycTWCaDXG+Y
yK1l/44nFcW3jxdxX2vMJgY19kQgQ8DPi/SKrdmX+HsJ7IbNgeg0cv/lbr72
MCvWQyLUwQqdWl421JlJndDyvgVL+SnruMfTFA/vgRFyJJBVztFnXHj/z4pD
L7tTAMy6THht7ZJ3L5X2roIM6UZZqDrWoan2G7MpZWCuLUzooqxd6B0HvAB9
48sfdpywcCJkgpy4mJaEnTZJIUM/1jT0rPr41Rnacz39g8ViAqpmK/KgvTAK
NJLtRr7/uTwM5y1wvApKQC5+jJBBDqzKqjI7fCO3OPWNbrgi19jKNhF2YGiL
tvMd1QXGsGVbf9SxMB9fDIoDalk6Jxk1D4JPUUMf8WS0ezWelPpBhPE5a4XF
LXRjpcS0x7rnkokn1xOmeAan4yKBezGAb6hr46CCqDejnvnjebnvMRNDNM1O
ASOdF5ouxU/i954GDKe+b9Vv8+YwwghNbjc7v2AXfxF/GVA1+PCofsc0P1/E
0rzhv9MNMI/+So9THaN7yutGbeRj47ZJYXjJbCSsLadJ6YiOBU1dIwNn43Zl
iJ6URgxZma5dabr7nvmTAe9m/af9mSQqdBLdzJsS/7YbxZZQDYXTYiJn+xvP
P6ApalpDRLQ85gcGE2s3uhS9fZxAL5PeFwE9xAey8QoBn9Rqh8qyjx1D4yVx
4a88hwyqV5Ze1mkQHTUUdNEeMlQZwZr9Uuaod6dvJOnuRIKft6Op3D+pV6Gw
LVMej9x6Coua5OVBqH4L9ZDbtskz3vUfofCnLiR6TBLDsdgAJdhfMIpSGeep
TTRaV3VlSyIBwLM3IxwUwIFtZ7VOzcWrj1bYXJX60veQXxY4C2wrH7hV2DcX
BAqneG+p/svkj7hidCflfjOIweXNTwgxjOwm9JiE1k0PxG2KgzZ4V6FZQcGT
XNYXUJts11DrWXaNatJYSFu+cKwiiz6rRrjVgpGBKzDvntOgjFgDINwPEXDW
aNgRWowGd/IlaYo5Sn73eH13xNdH2XIFQcrXtrtz7uLsvk+7xPtv4zFmVH4y
TWnjeUP44+45+jPBAor1FOhppklSW7LdiW3s95nVGhT7vL9rLDizEKzq3v5H
c7qKBHNlmoQyUIawurRDEiSi1vxNkFnatm+XtiAHHibtJMhbNu4R8o0Jc2UD
BIfqFPo3azhGBKpxYfia+sRg561lJ3qnAVll/I1vYEVfHLrnfiv+CcZZhHS0
p+p3GDee3dOuAjBNzpqSaJpmGLaVQXkWKGZBuRrshpVVbtNqy5Ra5rYsdgPz
5ZwNlOwcLHRIRT+IsquILB0vUbpXtCGGwpyOthYrnNGZQz1L60KgUUlj1FdN
Lts5jyk0no0IpF4ciO62KIb+mlZHaLP/bs2tVKl9XDi9FCRBKA0uRjuHSYpc
yGKmvrW7AJLQCrYclolSJGeEdxh0bkXCDKI6YUhfGssFq/sG7JTl/QRW1Lw5
P516bq5Rd5jocdqBwQVQSZSQTQZf44Fh+8kWk2uPC0As7Ryj/tJFBVuUehix
ahyKDrSLfC10p9YligcRuEvCrQRVm9FPvJr5XM7Li6qf1R37ArNI79SF1w+f
euDgaYxt8WIsCiDWW9kwx1mGVjizefpHM+tmf10zkUVPpf900ROjLgpGFKI2
DvQVMfMfWiCwqM1X8kGbMKwwQcJb/9P3KIeXIk2FsPDkFWhCHqe06hDwCUrW
2pZI2vBLivnzOEiYB0NBiuqgW2GKvh/vQOL0edTQBtgBmU8DKuGZBr4K984N
Kpog+tr8Q/Cnkll9zVJfryOw136pz01qW+57K/v/6l/nTEJHeL16i24tJ/Rl
4YAyF+3Dzc5o735JEQFuFrLq4m/xQNP9g1iCpkcftyNIoirOucevZ2+YBSJO
wQEHqQlOQjgB4HHvPWv4gAugzZj6y5REiyp0c1FG1mo9SCa1LzepPrHMTyas
VdmKENR4RWlbWHIYDoriXdj/xHf0psfbGaXwmKEi6L6eQ3f2ZwEtcBm/YcbV
0SZniWrmy64xZMeH2pjyBYQyzFkf//hijxhVSIN10fYIX5QAnSRE2awvZyaP
3AyQ7D/AOgWUHSnloH9Y+zQXvBO8CEGKTSikA96dJy2b/jyRQe80sL+mi8iN
/DiyjThX0qjr80OwlvPn+cX4gNPi7fV/19HIcCixPeTe1RCVk6D/7Tw0JxOZ
O7Wx4/IM86srB5AFKzADcx30I07f9mNsgpuVEhYSW1Mg3NkZfqnWk2CfXZNU
ycJhkxGUGSrXeMGn3NMNDA98/OJCUkONsog+IE2Vgk1v1u2mxlny6JmW2q2r
pZWz5ekZm0WlEchtF7jMNwwHd7qIIAj852YjRO+RtDULP1aUz7cctO7R4FVm
JmYhFjbfaB7u1YSUJ2k2bdZngVZbS6KjVJNCcdE2DEWbzKCcsbat0VTlIjD/
Wg5Co2aZX1GZ5Jg/LUJ87lpiPttseMiP8vshQE/pONUJIzO+sDiLRLOJHk5f
SQ0L8Ga/FjOZH9utuqJ1T/Z/psPSyHh+9cYazKTmELHKXNjDgdTvTuxehmSd
0+4Y1YmqM7h2zS/GtMvUj+WNPnIF4kYZHxUnIU/c6P92ytGf8yU5EcZgrOI2
+ZXXge62d4dcKNXbmQBM1vOaJxh3ntLrQqF0QvBc20FkTqD8ez5Bl6HSnATf
+cL6Va2sV/o0kGRd0DZ+LTWq5RWm7c+A9deG5xwljU3A86K+hVKMKPFSc/7f
YHTY1T8AhSm09t6GBsb3bkaTOLF+d/cwgcHMlCr0f/O72rvJQpfOiErrrnh1
JtROa6JaMYIDjMJiYR+49aOR2YnsD41LI7zs7JjgtGROCHuMhoHVlE06dWsY
obfQUkdiaCLH1m0E3a7o5zkvsCEeBFty5uf1V2A6wzskLaY72DScKZ+Mkd5l
kTtHjECU3FrSqJ/EjqOy/D41ERXtWmzsKBG5rMcBMkLS4g0lx8ntNQ+YNcUs
IO572rHQ923jrQ4k8OHU1WlOeZRdELdwktAbmjQgzqqr+G+pqhdWoUa6dxMK
8X4Z2oKnc4DeFcuf19SwoUGzEOWbZFkwpTV39cow1dayhYqaDakJncNOT9FR
o45mLrjREmNeYL3PYSKMfuZmLQnvnfBEcTun4IZsuwqwS8bUepgXTqRA0VgH
oHGBg1LdOvyXCnIMX/LuEnjR0h47t98z7VJgnUw4m4wolvH/3uCK4aohHBBc
IMYFpzwf9CLDNXh1ZNC5PW69hcPleVTTwUs3lssrcWM/7UKAJI9Hz04fQZUb
8nZoRXCLYGzftjATmw7cRV2Uy8qGgWv38RMfldpYRCxZBuxPXijPtEWG9POB
xZBkaHp2pZpQclYf7FHzUnpu+kbuOsF+9uvyg/Ku9YBDAZHc3A+SiJnbWnuh
25SPXegu3qG8nunHVO0zivbNZglvsK7GVsHqHh5yOvSxATss8UvkAmDH+se+
/2Q77Wux6yRonT+pqMZww1vS1rSieBhbCIioDPR9BwQfPlWsHr3D2rVsWu5Y
ZSAXttbTvE8+nBr1cjMvTm6YfwniWUJv1FAkJB7PBBichNRO4V3uENhMvpJk
QonJGwClBQwALmmba1zhEM9A/iGJXh1+DZ8j1WzDyHpFX0gQgGIWZpniNijW
VVstocX+9p3zV+agp//eKUG/E3HTpcaihgiVEwo7bKlqgHkqt/sadLzOgzWS
1jy2jWHbZ9lDXM5WOyb+7KrABiTfsLEmHqk1rdzEUcWEUuf4kRnHEyP6UqEL
1vfhCQ7RJAQNSWGdM9gZpBAurcfl4tMOY4QZMgLONQVUBH34g3y+i++KF7Fp
BSvWORJSF2uD3rzJmhKzntZknfqiJPybPAvmfbvIqHJcQX8h2bvXRe/CjcR2
yYnqS/bHmHWk1hAXZ1w3aJQhBHIQ4SGsA0ceLD2vCT0X+mM6rlGCg2PTLNom
Ge64DfVV7i+eOpM45wHpNqYlNpyzGr2MOvfNe30Gv6EaPXxxddaAqtUdxvzL
hbs4qibLPnFEHPS7irAuUfEkAeFDP2fsYZjQ7IT4ridJCTZb1U1tFGj7gy22
XOYbI3gZG7x0XYYU9hMerybAzeCd4HQiTtngJ+sJS4do/KuieY32uDSJoC9w
SpJnhVjsftwLdgDWPjI/uRKd19qPw+aviNSO2QGAM9uRIKdYe2n3lw+MQ2+p
asw9B/K2elurYd/e+juTRz4AflPFcGN2fj0P2oEk5dnlUCWFZFiF+rpqsk4a
+fgodOVmFkKSu1SJfpg3rULAYunjU7pxzSH5meC6Ca6UCXzQwPy2/FQk1NpF
EKewLdub98yX1Va6xqLFVlrCHx9aKu61tyoADW2+XVUVgbPyB6tYyB6WWfv4
s5i5S2kaKen/lQNdlrKMDiTl0nPYxe0gXwgaXwxgoInScgr+rXRU5n3BW3xv
rf2eROIeyiihEe2MuLp/uqbZfWIcdokLbiCvrNOdlIibXHKYiGSd6npGV+FK
jIHhMaZnC1EvD94ouRgfYS/2bVOm13gUYx0z530NsJigpB549h/q9n0kHW+v
mHherH3CvU+xJsDFPtadyF39JoGBPolIsGTT814I75c8OYZyz1GKX6Mi58pd
vRqV9apPXn5GSzj4rjjeKyw/j20wjuw3EeE+3nd1s6k3g18fc0916o3gnNlk
y9Nex1A0QlVP+3V9ByrRxBuMpt87aqsqwx8O//tf2Cp8tts4ZXkTu/lyPaRP
iIX2nxDCGKwYFfFZcJxnENY5WnIKI0PC+f2J0kfWsPTCGI2gyLIUyoYMe+cc
ov7OUDqRulZ6Og6fgAQEccmlZk9MW9kdPZCxuglPoDuOY/NISToyns8u75Ny
LgdrB7u4DnHJBfM8G2ZjmPv1XwKhrxOCWXmJAxAHyB6klAatBQiBNsVaijoe
q5vPSgQIiPyrC4uMFUEg3m0pcHRb2isgQW3YI60/TIMHFpYPltqYivVXLTuu
N5IKV3QtSmbCTpRJ0CU5MtnhjyuLg7FoYsaxyfEIW3RzfD2cWbKXtEZG1S1u
1pvnbEQjgTULwmxzltMvyGoE7ZPx2lOw7UdmLRb82M7WQSsHnnrwttMVOBfn
cMNT2c4pLFh0EEh8IRoTkVUZdFBpx7C97bDKaqEGd2plwm22aKbQQ/4e+a9f
mRbxexG3WqGSc9SLQKzw98dOEM+PTYLrzxx36rv/Ta+s9fDoZzDVXAirOTMR
afCUfcFLtnmi6Xql4ntKhWuUC8ABxa5CW3rYATBhaFbNkEzg1DBOkkGUOQbh
mYVNnmjdyw1HMcpREYdWdy6Ci9uDhG9tOqXiuIKAhNOmHnYQrp3d5IfkcDuN
iJoFOHZrppuytkDBzLKsL7h75+GUBeIry7j8AXDWhErKQXJcQfDo8Eta4qnW
EhjGHRkumZjGlcIz+8kEwuikvjyHfp2K+TQAnAsyCwHCg0+6j6sftNNPcXCj
+U8aYLZeF5jh4u2tc2PEJCdotungQBsHXGwveQlUka2YR94UCBLIHbx3gQXG
nZYhKNH63uxpzkWUW1vYdMc92CIo3JGUIMRVHLkXz9miYypbZuCACGMBL6yS
zaF4b+p/eMBcOXV1dxIyp/Mn614AkPUPSLCPjtfs8NbLVYsMd5vXFfvPf2+Z
J8YSGrb8E3UMmNIunOJ3p+F4x3Yitz0cFjTmz4rWZZKjt8R0d0I3/1/UvT2X
viHJzJr/KGeuvuGaiFzHUZRdaEeh4Ixrxn8bOkFuW+rpAhscgmxffDrEKweK
x+7ILwtlYPeafCVsHdkmYsAeyh34d9qOYSwxv4vdurjOMprp7GjSui/WnchP
8bDXcGZVU8iXDmGctOzujby/BUVXKeGNQc81UZnFNGWpIldOgumqr424UiJ+
z43vA9p1mtZ22bOairU8ipMbXi3oww8HSIlMbTmnXM1aAK+LxLON1mbQ2ycY
IajK/dUflLcqOHA94jtHVBcl2k0/Nki6Qo5tuaf4e9LWEGBaHZ4gchi10oOG
2zccA7XBCEPhdEKJ7hQDLwnK5XVC6kQ0Q/GA7PXgQmaw+1eFnUFKF3VL3euO
qVULOJGvJatn2MjLLtdI8mkA7rdJGlKm3awxQxGK7bvScm64VJRw6UGo0dBm
wx/HUV/JyqaYdFDuyfrA0ATNRcAf4kjHT6RFN+czikznrRVdWZuNNV+46RBC
3wECxGr+HrI4uzy2xOR9uwwGXRu/2dl9oF4UNcfMYe5wfa1tVyi34rcdFk0Z
1JArYvnAiCmk5DtVH8Tax+Xjcg4txAPW4hT8+dMkqQYlYM0obQgTtCidLCs2
tBKSHdqG8RfXYrdJBXP2aJWVd/Y6+kiBL++CsM9WrlxJ9UvE2Pl3VsfnDxRL
iHi3uhWY2gPqRvdTwgvPoln1p6o91yQp8dpoMQY34BnIudGqKo0i67K76pqA
X2Lr9yVxbAi/gr6YU3Ua3OKWjvzb/g03Om8DEsz3Nbm+39qBTeLXGA749Qfn
Ptx0mrayilNJVUDP3NJkkAPK2EjLTppQbrKcbC1HTjMelN5byt3KLTFRdbml
q6ar9mGAlFqo+kuMQQGweC6x8khNcZdtaBOzJKJ6ikJSsnv5Po5udO/MNZwF
EGKHdmVjz/46LkMHxMuT7rVBfVY0cOKdn3Hp3qXwPoUIo/WdoxoXUdSIoJ1n
J+7mYyVKlw63zLWROnrdD6ok/sI+ezYQnYM9qxN19+GTuPNkzhPc7lzLLyhk
hIUjDPXgRV+j7lwSP+2HHbwZWTcaXXl7102eEdDjqBJYETHfyDzg/pJ4mFaq
QOA05c6K4q1sfQCmnkmvYZyOsrRChkIMcVyQrBkX+TZ8FPxWrjPczLjwVVIw
Fo7Cd079byXFLSdyTl3L546CP90mz2iDFfdn+7+auEIwzKAaT3MZreS829sA
X5qfSlh4U1bUl6JkP/I6+j4p3RnLfp/suEKkgAlsyMf5Mjbd4ePZ4gEYU4IY
UUGTkuzqCqPvAkAGy/5KBf9elMNLKJt/cqm7++y9gGXEf03lan/Q58B1TmTZ
CmlGGm0azBs/PDLLgbjaLl5KAXs4PXRvHV0FIMJwCfjYA98IpsLTGzDzuz7a
xFtLv6NHKxV0lNzevNDgKVDRgPQX222uXVk7aim2UOLwLAoy3GDyaMtDUARB
Xn6M6E06HnW9lWHUDJL3BFE/54oK2perHNSDDgcm+KwsQ4U9LpCvWkI0Lxc7
nqWfP0+bR/aWFqWTDdz7xflgZ71adhOidF5b0sMMDM/VZrA7UDEJwEJpq4m+
XhxAMkGMLK/FlbKZhYy9nI3KdnRw3k+mbltTqhfcXKBRrESPoIfieW+Es9a/
c3pFmPX4hzSf/vhKJ+tY/DTw5h73DQeA16ASqI+tXuQ5Z0YsuAs8db3xDLtt
XWCQHHNYLiqD4cDe78v2CU7OI/hATNudm7KTb02gmvPpemXpSKi47jSywRSq
/U8Sv6WO2tjhSQaWu9DkucFpTJ1VA805DV0tkkiXifSfJvfgTPCWtbLDCJcn
VCeR0gdqox7KtoQ15Iz75UAuAHDFnhE5eYID182QUw3di8Ekm2x4XFnu+Qg8
CAAcETRuYP3eu0OVopTVWFYveDkUP1hXhVdzW4Ht20Tjx1Mvjnb/3I1QEvCC
yIYkuX1GGWd0ro5pvD7J93wekPehHfLmEzRFdFBBcb0VsMC+q1Z6W+/NqJWr
PiCB5hCMJ4TEZK3NRW4JosHTNTgXInbWP8Z9MVOkbu0+Gt5gXxzAApTgbrcP
udlQXLIFugRTX/GNWDhP1srpIJM/fA4xw04pv6izDgX24bbmR7vPFUf0mILZ
iI8bUhxM9FMy4Pk7ZghSGDo2900XFaMato/dTV5LNQNcbXF81c8SWF0fAl0v
e7PwuVickcAS9mit1rNOuUaJ37Uyf6E9Mb4i6SWK+GdbSdSp40GJV8CmRdzy
p92cHW20SV+UMKgEzOkaaV7KfFByoN20NImD8Jkiz/CaJAQ7l7+A/GEtfoSU
e2j5Vnt6ji55eInExBImxOutMDGrMCIgvqodjcOr8D9CWwebY3jmx+ZtRMOR
zut2As8kGpmKMqIYaGjeRUR5xzYCcjreOsAjGc4PVv60ZQCoAeaCcIr12q+y
ngVJqyMhL9UhPDjvaJoOGqODlK2RcnZ8WhaTXWMDIdGjG+DADYxVogeqhHMO
BC8sGwn/1F5fhMZFFv9fwFllZP6Q6T+me3x4pCwISt4xKzKWiI7+UnQxgzB0
hOJuM6d7Z49tCH7tC73rQqI4DDP2M4BvjfSG2lIS6F50WoKSivY36fhGYKnX
/84ZzqHug50+oFlTBo4rehiIvNKTW3Hz26Pry7WZA+rt9yPKP501fonU9FxB
yHXEspEpfgjUriMsQV3Dq08dWPT355BBNO5ZWd/X1fsnVNsoi2Agk/Jfyxpp
Bl6skTxOOAaLCoevh8VPgTnQulSK0llsDqbstIjLECinMUNXRY6k4QH7VoNe
BiAyAtt9Ix/CprFXgHiDLO8AOnIWWtjVVwFs7lxY0RW7cV5Ahsdt9soBdmy0
6pSRoRnA7c0lFXrgW1EDBKqPI+OjmI40c2fkxrn+9zdNkJXTx1V24MJyf6Pc
UlBUj+G9bwCqmrQZOCPyucGM/4S08yRwbHUr9jdk0gP4ioeuKwCEg86Y3Ywh
WswYA0DR1mMjBDoBVEy3kO4Sq5Xy6Qkxvm46QX0Tm9yuGYYG0B1FzeLZQMne
/W2o5u4PTUXQOd27uTPMPQj6H7wpVg89hMCUiNN+Z+RcjZnog083yQ5FR51S
zlPUqK1MUKPQEiKPqAM1QasiyNig5/CQgDgSTMNlbxgF5h12EgAxE8pk63PB
0jdT9tCo4TyNMTr/B9OlasE5AkNzItGbUwZjtoX1tlGm6NXxinhhHjo4Xmzp
5QwHIydWk34CwMtuOK0KlEeWb2ZP0qRTKssjDvOH3Ql5ESCBMqXR6cMaxA2R
cClfpY2l+PAEx3tv5NPn8ky5nxZwsR9HJP1ZZedlqJ9P7SiDbkfeM4ZvoX8c
a70KgYrr8koKav1Oxut7P+CwE5cOvKPxCNtu8fbrsMewn10rAfxvv9mAgHHH
RyIBvOA0A7RhZgS8FQt5K0tt2IeamOOoOPmDvRStmmR7HEbkCRUrsJX8BhQp
e4VcMiCuBxwYlWzqSd0xMrPcB7w/Nheiv8HvXc1aXzAowOOrGoRInjNDh4EU
95GM1t37n7syHzplcpE2ka/HlGBelLstdjh1rorg+sPXIMNapUNWxCoryxmj
rcWIU3VzLbvMYqUxDdXCtAUl+nnC1tWV6RWMnSmIyfkardxZEEretcL0qfi8
UVJbuiAMmfAJe/OXYTAoEK2oaP3OEa3jUKqG0p8vRORlTN5OQXea2btFTbA8
DjGdt4+3HUgIqzrvrarsTFeMYKxgdCwZxzMkTUNCFic9pHZACFhaHkhd3x7W
SIVIuRh/KU6zwp3AiVpe1Y4HjWD1dT+LwsTEqgOaq5BNaSGN3Nr35raPko+O
OOXwjBlZnKKWwGwf0pUy/3VIjRjVbmPq/+bXk4vzOVKLHOPpvk5E07NBCJNt
Wz7NdpjycQkOq7kj3YhUt0uTnPWxedBLE+EEaXhi8J/XiV0BYzDWryrg4FXA
yfPBpDgp+jFpMod+9W2FVxs13HQg3obleZltwIM7gxFa9AUxm2cru2tTi1XY
VqLEIUJVjL9Rtq7ObhUgAd0gobUw6erxGbTRIbWiRlUdGwEuvscBpuGlLE0L
wpmyTFNYpoPi2CvUJRmPAWMGLr7KDNqcTAVhoCj4bzIDMvdJdt4Gia123UiK
4C91owWaFF0sPAQ8Iu/T9Bjk9pcJLe1TLsL2wslh1XwxoXbIbaLommAbkOjk
QRqw9t2GYt4akiPkawn4hxGzQk/G19vNFhwGDRCHPjFCnwj57BKVdw4tL5DW
Gf5PbKYPv0eYa1R0C1iFzTvRNZ3j1hg9V+fUyJti96SZaqKp3UhgqEQnNK70
NmeaRModfAAMPjjXiHcL2NAK3HosKPnZW/YiMKq3A+8NUmQJ8AnYn2kewO9m
WCFD5v3QD3I9QY0iB8U2xefFjZVdfSOKp+OAfmj3m4nsyZG7HDrFdmjnC4II
UwiBi8YgN8AiIX0xCDKQwtYtJKv1XP0h0qBRnM0bGXvDc1D4dgVbvwbRiFhy
o+rsojJ+pacBj31x8oMMFjgdued9e+/v4te7jQsUP0+1Cftbg0Cu6MSEZU/z
6ExHGGXpM1L22z+91JpA+xlMOkvyoY8qGiTXdYPNF03+cpq54BsQqesB1vgn
V1HiCmMcng38JkXdksHjDvBNzqYiDMN+XdyQAP5m8lV0ZZ9iExirp1JiIX6u
qR+N3owYyS0TjcoFqut/3ek3VdeuNhVrzdqyqe0MvKXVka90ichIc9DHGdVn
jYsbLyyLq59QyA6K7c9Jde72EiWEkXE1kvyIKaThJNu5sPwd0fyBWpKxqyFI
MEssVBs0ivKcan2T7c9tz7Cee/xkz2VF4hkCpgX8lZVkX8cZNUIao3AuHkH4
vFlXyOAAs00sHbyJYfnkKs4YoUO0u1W763rKpZ7wet2SJuax5H94BPoi69BC
nKBkABeD9WBxrzaM6L2IS5jZMn6++CsFlCKhi36bRGl5PZGgeuhPC81n0TJt
lm60OdPELRVSCvtuNZYPmAneF6OMe2a1yF5pf4hBT6RLqynK7qHPspvv2iIb
yY1kWAoUPTVes/hiEHn98XflzeKYITU4y6Hii68vbIz1ISQiWt+XeM1CbJmJ
TKZved11FAQenWpkSxm1O3fjGv6gcN8EmWCntatvcTwtrSkbBiA3KWD1+4UY
pckkjm+1hhIuHoV9oRkOcBGHj1hmbFw/iCY71a6XLIYj0ua/ltQq0G85y8pS
aOEOa+Vhremw0Q0VXwumNufu/5RWjvdw9KkXTvbsmWdyHP994Xqf2lF6Ya/z
i4huOCAq0kWbSZtOiq6oygUuXwca3FtCaaXQW3iOLVeNtdGHCyqPmke8N0yN
dPfCgVwfwt1Iz9LTHA4/DqvB3K/3mj8kpOqAu7UETDrRkh5AFPAh9cjk8ws3
DDp/F7ZLMslBI2Ct9gTnqGImtAqg1Xl2REhWtBHNL0vZyy6QmqJ58Oe2HeZV
3fshGU+0u/o8KkbzEBFHFRg9CHUsWohlfeROopCoSAXKIjitopkjiHrwjHZo
sn2dGcxnKcTbC1743tuKg7f5qMKN32Mj5fknpaxUUyeBaqlfU+yIoYcJKml6
onuPJhKNKwHggAFyj3zNf55VQ1stjZ4oIOey75LO+iV9OfuCoysIozoXwdqN
JzTgx4dWTA/faKIAh0Jf7mptthj1w2fXKm0wPCepxJ8Bmu0VVhLle5cQkavU
Dt84y1WuQUFvLplbtr8S+Pj7jmkmWWu8VeHcWn279GYui8fYrtJb1X4bEEUr
KqafENdLwARhEJ2jjYjSuh16h7vhfnAsW3wWx4+KCdY2rX8wv625u0F1kMnv
UhrV9PXvcV0QTKM0G1EhvXANwZZpKV9Ch3KrP47t0nUWwK9hailowzr5jVjj
BcLXByUTABeFyqt+oh0YndfWyZ34lCrSdFdeOv8AVKrWR9ftq2GftiMa8LtT
8LGivZv0FPjz0U3aHoY63pavlCLMWnYACOX/GdU1HyQKGEslzSYBfscLfrcy
sMmJFas+TlA8KBHI3gP7JmO4Xz2+cp3qzmu8CmJRGDYNGRipUl9Z/tnvOOxt
+xouPAOPhMNYZmx6jrHSIqnOBE1+IESJ+WuRDU9Inw03CimvYHs213TDbRcd
pXcGRI8gQG5WTyv38dO0//3yhitieOzwZgM3gwW+X5EWs5OH6wlCAblYliV1
AJXcayYfIbQ5mxFY3J9mzg/FOJgy9FOFshPsnq1IfkFhMT8XpPQ4OzMKfBlw
yXh/mZFAwZSvbg8602X2FNwmRFHQO1FdH1ja+gasT3wE13hPQGEyBRQ7Jm27
p4TBb6XMNJh/gBcvsPNavKrCk4v1tjknO2s6QvGK8Zi1fqq2geoyV0v/xa4B
+wG6e0/QdwDuCpJFEwtT56F7+Q6e87W432QdNOqoaZnKlGAvig+pAOyx8qyI
ltic87LedSdeqeXyEq2IwneEI6HtsiUE3DtaG0QgUlHcLb6lKKXmwQqGAJIE
vNe3FY64TLxEkYNVIFx2fKnJjkfYTaO3TVm85nD0F5f2sdoRqFEdvMS0IjYv
bCctYrB0VUHuYzc6MTX412JantOT/O8ZKHucmp/XYLHaySzeBDP4CNNHHaeT
WuqwgsDWz7pyJQbU4nhD0i2MH4BHuI7gigB5sY9Kj4beQZ6rzoux2p9tYlFW
9aTyoGvjt0xabOH8SfgJaUpiZBcokLJtUV7a/kps6vX709H+G/HGZU8VS87k
ceAy7HFKijpMKli9OvTzYYFiTAeg9JtdVdo8zfDO7oSnqFDtcn+WMbdCdHpR
Li3lCocIgydlAkx69HpcILE7WfVS4j45GKdoXSEKPd8hbHACZc7Kn4SvP0J4
ZnfRBUMmC9CzfVb73wi5C394oqWWjnaCxVlBftQiWLSObn/unxJOmNvPHft3
x4yp5j9yWz9oHQGNxI/7pGzbLEH5+wmIiEDG0mbgK35Mi1mcPC4W/PgWgNVM
8RVJYRM9OR+nXHZAJH4jNhlWpBV8Uy2nluNgcPkHZPkZMcZoU/GnM0CbaRsW
TVK0TEClQHW7VduCp6XoJwiQZaCFs3abNxrFactAKjN/tFXormtn7X8uiJFd
EhzY5lkjRMbVKi6QuHdyy5mHSLUSlK+hOqXor1USb8r1jzcGwFSMuGizNasz
t+/wjEfvQKwsV3rwBdJNhWpC9ysJimgQ03Io6fkyf2I4ux0g4iTY4mbJZXec
Zk0W6H7qBLJjXqy4KxXWp/4RDzOG9T5O5F900H7j2MTVz1pvMUO9MS4WOtMR
Sb0aAWCc/e6TgIFVQQGmOPu2QbzRa33vvBhG4KI9qSB1gNmyka1Bc2XCf4pO
d5+6VFg00n2e/zIVLifhUBOIIE34S2xaD049y+yhP7DXlUWIuuD/8Oww533/
wyysprI4GEpJjyWgWRHMQ8zjVrRjhQXH6x300GfAnEnJf0TWSxZl9eFdodpo
xkUY5isHE8NcLhDD/8kOT+xPdUQuMp0vhhiAPNb+NjqlOCAUMYYzWf++Jx+x
DqFITB46EB+m9OUAA688ccclKyjb0MCEC8lUlwmtBEUFXPXg1/fWag6QEQZz
7Rcu8fbsMxfIf96XQmp/zbstrlkcjKmbWCcX6cfSkhGrozGUFpSmevVBVJMA
wotMVwSusl7AMlZzLcHKxtSFCT5RxusnX3LkObIA9e6Duq7LLNjo9nFJp0Sa
XcbLT/RQRtFUeIed27w2J5l0u5fawKucKzJJxIA67xy9bgiunYeOEwP9/v0n
MXUHSB3YTRwyXx9Y9R04WdEoygChbLtXluZvU1w/Gaip2wFB5MV0vrkgnXOc
ts5GkNHCJBd+iq9b2x4dXclgF1miNic8BhRMTSqIYk8lZgLwEVhTUiH5g7xZ
DjM/OB4ARdOuEXDLvbBMY75AOBaH37c5imy7W4H1Lq76KcRgvyEBlIWMx0S5
sSxj2AMphyve2FFWsaDSy3CL3KQWedW4RNaxXXZXGznYx1cHiTLJ2MvXqobu
r1j8BmZA/5hRHk/gz74UUgP3fB111pmFEfMAXsPuxHuJSp6v47sOzBlhOfSt
7+MoPsQrcQ+j45DYf+lB8EA9Z6Dls7jIznd5BvlwJEbHbZt8iriUqWfERMww
+WbC34HhLzgwaKtqDsmBbY70wmOHZC2EMf3ukBbIwFLTkH79h4zV6FmnU7x/
ntL23MEuc8ZwPoZela13uYJf6onRTD7aufuq7jn4fUTwH487i+7NjiQfM8r5
KYZcDcfd1uacT20Hjysq0W6EvZieLI3lpNsg2suRHP+jN7UDHF8mBEGDiHbS
KF4nyYeTaT75SIeW/tRYV41wm/i1meytdQm+VRRNu/4KrozZ6J2Q60Oe+doe
2363O7QIhWwjILYw2ncgaEso1hCMIGsWyMDHxoF4Lu9/W+Bt1diHv9ZO3PPD
+XD5Uso1PDdIJY9RUuhRisT7tjw1DRaNWXlQOA8dC95+43YiWOrw1rqEOoaY
TrzHpg+oCy8GO9Z12mTekdHAM0RI2buCklohXG4hJV0vpN486BQeA+OdxabG
WDoTRhK7OSsBBKPx6LawVfv50Cq5gw5DGh9FwGVeFUk9Ztlg9MHAzTo7iSnw
oQDKz1EEXuF/cdaw7xaV+FU+nkQ/GLEYxc2uTff50L92ghLnvuYuIHJjnZzL
jcj9LIoXADeQ/Gxght6P23OI/+nR4S3i+dgZ1vRbaFwTxTn0R6qPAuRx5oIA
cIe4bJwMv5d8lrYYwyOe3x4qreIlKjX7PZRrYHangglaiTyI+24uyJFrjnuo
6x7oW5yvQT88Vv4MzKlbV+YDbeG2s0NecIoL6gZm0Sf+yZw6n4+ygL1H0q56
t9eH9QKhnjcYuIEbtNSpwh5WPFwbFCbJqHWti+77s4UExdUBwQogfqu//aes
X/HegRUR5fl3HeEbbGh+XbyT2gvtXFGRlnNNxGSUZ0e+6aAOciMJ9pEtxRkH
6lcJxnDVUzXW1M3end+7Zp/wX1fja6eCtXHXbpWBlti3k5R/cTcW/C7/aQWT
S8VrJo96E94M36InPTK+EXvu4Cu8pmfOylfZbz4bEmru1AqXqqI1ry8TpoFq
3hcSDA9bAKh4k/QZ6xTN/ecds0bJfGoIL5sn0+1vNRCLBOGepYcqsjijsnb5
ElaX0nZZCuPQxLddp/L+bfsnD4wr8pK+GVRFj2Vcr2V52BV3etqgEUZab2/u
aMyubHgMixXfAUhbYe5DO1nwPetS3F3d6qNB7RSC3c04vzACDS2xIaC3s7vu
MpjR1Y3smndOR42JtghfYocVdXXItdBE3g5aILMfL2xeNq7Rn319ky0+ga76
/aT23GpvRXOE5j0h2WdJGbfaoaXAZU7RPnPsyMePQuArZOAsodWweK6REext
GoRXIaLpQEK/X+51oNZjruQj50wUOr60knmml6eLaS28g4Ft7TBQQ+3K65B/
YQvNnR1qLUM0lE+sx/8jm4oZs1c+hNnbxaWyHyfi4+3TR/17vs6cY0OE9lyV
Kd64BeLBglwMebYShbIzAgPOdDYz0IVoz7P4GrZ4jN1bCXlwprCp71rIxcKv
+DuVU2QA72OU78qPBTZdutxHqRGEVppSA50mR+Y466TSAmS3IRx/uO8w3nHM
Gi3gWLR/7bsTXJv4Sco7HwTNg94unRGQLHq8jRHZ1wZeK0u3zbOvr29N2qYS
b0GmXdmwDAQVN+NQmAJokX6Wkqs8cwERAje9n/jzPQFnXVjimyslEN0i9Jkz
tfn0KyL+4uXhO/guvPidD449cP9+JvA7q+zPvu/nZspSGCX2rjuaIemQnD+k
FlsSzsv5ZG3JfH3xAgz6r1Wfg7o4YvYFvIQRz2P/t3oT31Hq4ZFwjVTNd1EZ
ExhJq4mgpHijXJgVA1eS8KWLZsP8OfsQf7UTfM1G0/FchGaZDupd9h8DAR9n
f48YXVt5N6CnJ4Wnz9JZUe6Jjcbwh6SN2/zbABXslnah9Pj3B8OM0Mb4nJyZ
xZLg+WpxOZt1k9QTymreuKVfGRXYZy1iXOgkt26Ey2uJ9RXL30MgqR8yp3Jb
q85BYsNTFh+vrta6wUO3Kt/5M0qo8C2MLyPKiHloYsJGhdbL5T4mmnwRJnMG
cP4KYcdWfHTipSC/AjB0PmLK94arkXho0/8S7zAUkV/I8a4aOA4pns8Y9Pl+
T0NH57+Nx3cgCTXCWvoRLsALq8/R0GbqRd2JrzJVXFTPb/XkFMrR3fvvoDjG
1Ulrzukh31vfiuc+gItTlCP6A48H5XpJlqL+QnJ6uAG+Cw46nu8AUPmqfYzg
ZPg6o6z3BMbNywmWlF/ZldxriUX09/jxTNc0QZXtYOTz4DoZWOy0j+kg29CD
eWG0K5lpO/AhOWIjwDvZ0d2ZFcX6OP3eU0qfZY7lzaYM/pLEMfbgH8sU8l/V
1aMoqjMPmCHMU70FsnmDr4P4mhHMHFXX+5mlX9HdHwHqJFTsj91z7xynRW0M
PE80/lj1jj5C3QQZfsYLfGCQ1jQhtiDdp2cHeS9VJ2c9LnviQay0uwZ1U/3e
RfIMtpPdzGQm4qrfPsPEtyB1NSn7vRycVWoRxRgw2Az3n9y3ixk2sE2SbT8q
8cFy6/olNm/MLyuJ+mwSM8hR+9pwKFkEm871OIzQF+j85+JTuDryizuGeweY
fOmjBkJ+Ngb3siXrAtRFwySfKJ3WVOE8WMhzSJ16r+f5Ge9KdHNcMUQ39Nhi
xKXE3FyNWXbBgmf1iW82zoHoDJ0AlQVENDXx5uNVd5Kq9etguFWFfeBJ2MuV
U78hV/nQjTJJUu917uvQHKII7KBGlUbNPjm+f/XLw07+n9SVgCKIz6m0WoTK
GYdEco0Xxu8cij5PiuJZMbBbfCP00J8J8RZg1HQGzcXFHcS6HMRW7VUa7DbF
YotCpuJkz9Y3wy0E2AK/11i3m8EPC9pnV/aRqh9iNtzeKOSwk5SgojT47lsK
GnCRiwesam/YYqmtgl3/l1GwhVcDZUgPkaSMf/xto3WMFgQODInwlruSYmOP
94uhRwkn44p3R6HSn2w6FrgTbwwXlzXm483aZFKr5XfYNJFm6u3GFhl4BJBh
yj4PmBfYxarNzTyehNin5Wt/od8h1ESGIlfTg3QtE/iARzgxdxpSzZFjH0XV
jJ8aLD6koHds5kDuFFSgD1JOGfPJBrFuKE8enz6JvfDXoy5bh0bwL75bNvbs
Pci3xuXWsd+HG7q0QG/Bqoq926uhJHGzOe/U/3iIIE7bGxwPc/M4tCvzyUpD
cKuobeBqFBgWAgy5sQa1NiaLw2z4/xfQVNNnFnbyVPKRIacDAsNjKSO8YrD+
RxSvRDoddEBU4IsFzex6yiIaPKXo06d0qgPqOVXMZ7SOvhKDVkKoKIAPL5VZ
efAmlWUeylDa80/lV4bf8xmAooPMTNjzGitF6WIYdWYAuGNtN18+YsXo9QyX
QGDRJcGvuN+QqzxHj4XvDtIBkPIWGpA/uha+t1BzuSxKsu01CBStoDjffjBg
XQE7crFpuFkrspEixCXRPuIiRkIxUBXS3yTpsljlIZKan1jTv5QBddEuLvt3
ACrhOc/qFkoK+xQYjPaMKekRuZ9v5ey7Z5J3x4H6NpDvkeoWeYBqiCmyoGJB
OGgrwgbJPeZVVs6LgTZ2KYU5wIb4UfSwHE2hhZ7mCe/RfewYhyqpWvv6CCVd
gXizB5utLEoeVDUL2IZaYtudZO/eaGRo1/uwE0Th/kVOetVN1CzATYKX8OsW
ShATAjRhZktLfRpoRQorPmzIUOKEAdQSR8NE6jSxQElHqLuw54hpNvz2O+50
jLfzKkM7WfiJE+OkG+OlQ3JA5CT236gDly4WBj3YyIIvp5pRO2MalIfDeA8w
FeZOWutDSKiPfw/P2BilU+PkV6sb+Osdb76/Lp+s/TmBrCxLl8LfOVFDntk1
HJ/oRzJZ2b+RZlMqvxUVN3nF15+Sx9fUcKbYjA0NrdQ1GDtxaBSZ7q71hrvb
ZdEdE2nzT7Vxe8Fnj0/DBwE72ndv8fJIjiyNasMFR6n2fdRSWGcI6cc6psVW
I6QCkCb0l9jAXxMc76fKNj4or41woc27AWPgkwqIaSoNLHH7Rano9VY0U4h1
3zI0g1fjVI8PGjeBGoMEuUX1ahj0uuN1i86T6Bs8ELVkfKW74CR2yoPG9Oi6
DfHY0FCpN7ljgolVen3ACpwb//PPSS0fi457DgliDUv0P4E0QjQAbTMaRrWs
tkFoEB/D/HpQXh/O3oyyonLbgXo+wWGztzPbkgcW8iTymuj5jbyDdZk5zNJl
bvBndacx60HHbtu/acdB5C8xae/mO6DanaEnVhcVfwVKAi2AXE1tGqPqNOkn
nZK39Do882gTYsKK2om8VsJHJBvi+tIK3yEWqO6/VVAmjdKz/XmJWx1lYas2
XURURIA4SJ4wgq0C44d3LNOlQYJgFuH98FtvjC1oTbBJ4/7ZuizwvK2rx5QI
vQEeg/Zg0iwetwxylrRRlbMJYwXjt3EEr0vGKMugg4QQbWyGZrjYU5nN8TnE
ZtMepmH2TfNQXHPJmxO0nfhn1I5PHFBN0Jm7ODxetn9LupX4Hbzqkf6wYgo8
HjsyloojEKElOWdTGa9CG+d9k7usELLR7G0oY4H/6WyzX7NXClmBesRu1nxs
v2cBXPDkgARnGBksIY/+yOD+yo87uPljfqKJAWkvsP6qUGE4rz910PsE8gay
1GarB8GE4wEKphYnJ4DpqbKuU3VEbn1GNXBmuE2/E2acKRil896Yn4Z3Rzue
h8VL2a8uE0GvUJR/vXavYKNWiOeJxiEAmK/ZtsBfqT5wYw8pITtUxzzC4q3D
9s+Lqb/3FiagrZPH9eT73B+b9PY3e58zuJUHjdHaow5snLsQBnh3rtQ0XGep
QWiBJ4q2dXJ/+PwfnmmyQE2csQ04KEpsHJd9PBR+zksrWlWgcMAXhwNtgfum
lgpqADzmFXuAA+/K6IjhWuy2hlDaRpASnKJXUKGx9YQWWGlGlxzZRPBs0m1k
uqaErwKoyOpCYP4+09lnT8OYh1IFiXeycQgQuruVdg1Z4M38FGe1kJegoZqR
T9Afk2mHv64lyBp3LPA041YX4rv/wL7trACNHdKF2wU8+RsA0w6pHXWeY5tl
6LYiTbTi1/KJe7L+izqy7hI86eSV7es7VoMh++iBAfskvohFdvgq1L5dTTpZ
jvs20AlKosxmM1jqUEi9hfTASVXHU9V9raEUH6IdxpYKE+zfnL+rzYOG9bpm
g3RrWjsmsW/Z4Z1WZ/o+smKqrkiOQ1kZYLRvLRw8e7pQdekSgTlVfGYuLnIa
AfcinjvQwqpkBWhLeGvSNP+np8O9xLH/U3BVK/bB7DuCzCRdMU0GQWFbKtlr
avVagUkgge1D1HRnfBuGaGYTqks2KaeZtrcXmIcaFdHMx/wdXzkXMcN+M+Xo
sr6Bx4aNamIjeDAB4WU6L0gkG3Uk2E4T4E9dJlqE7TiL504GeeLD8Dm+R2dd
05bfUJeAnO69Y1sMC2oV6O0WWKKZU06ni5USmIaaRaNW+PMyQjqoF5KvF2h9
S4J1sdvfqjIzi0FswlWrNu9KpaHgDyjee6DudEzkDuzyKSUmsBfa0H/hoM0P
8/Umn1eCcTUAHp3/ZxiZsg1/uvP5slNhXO1OXSVOh5/OWHQNQWlEiVZxoIrv
JIKr5bkZ16jXKh+sOOCWOTERfFpAjU9+PxNgBJUaLlTc8FEASMl3CmQ9uBz5
MxWvG9cR5e4Zj2ASC1QyuE6HBOZcj7fUemh1DB0UxcV4oeXhTVB7gmbYB2Kg
EpAWOz4HBrA6rd9A4EnINsYBtOUFrUij29ZzHt6rvsruD84w8QZLTvILELSg
JIsyo/aLURgjpKDtXZzvJdQ5e0PwlEN+5A8wKRL0byNq66jZdkzJo7/oVo+/
4PMqVPs9hWZ99WkZRGKZsCplv423kl1fJCS0joQiFCzlCaoIAhfEq7cPb2G0
tquy8IpbrKOtz43TGKvY5N6iKvYA2dwd7MjRT3UX8Dx4nL/EiF39LINfUExf
jThszZjMdk47nvAeKe9LYfW3Z/J1/BJ/rNk6j7csbA+doyEDLCSci9HumtkQ
SZuzb5LmY0BO+quGS2XqKuR+tvlA1UWctinOHRPN7rR8GPa2cUrE6v9bfj6t
mr3AuhQeUTHHsCq1/LsqtGvQIH12RUrc5EbmkyaAyHzm/m2pgOI2h4IGAlfb
uo+GqjWRXanxZdAcv5RzW9dKY+RdIchVAB/b69ZOFhEszQsVw0dSQmZf9XhI
IgC2t3WmuK+aW/hY1k+6pEsmlhyDJU2riRml2IDxcwBLBAs8w7mUlVlcK2jo
Z3CH4Ji0gxVEw1dnWLXjRhsSUo7bLfQxvDB3fTkoKCW05hTfREPv9B9PDUeB
+DZQdU4KXI24wlFdH2MZTParDqOHs9ER6jxXWXsbwiLevPKfuJKvnhCjglH+
ypm7mK09Ed9DdlPALlL/xq2eOpvOai73ymFf4Sti1Lx0QoHzqTnShG99Sb+d
k/BXgXU9GVywBTM7iHN3ejDBkayfA46EShbgChnQZqk6l43IaJQBSCJXrDSa
9Sm4SupV1FrITwGsU+Uyn1nGlLyX0Wraaz7d4M7J6ErxAX8ibla0ZaJ71A8X
FtP2zDhk0F8SwajpP4qOL+P6orDSdXkoPB3F5hMAQZlGUwzRZqCMHCN5NgJG
2qnUw2CGhUcstjaMryyC/Q59JmRiraJ7lygg7aJSsqMl/7CuAEtFm0fqKaU5
+qmWwONuEnDqJLjtOGPXtjZ7TyGHxj35Fs1wNTNnDwwL2phexvJOLq9RdB4j
4vvOqWA63YMBa4Nn4UjgQ8MQaNMbj/GwM+Vnpbs04Z+qoMV2ttN4T83dhWDl
GDidAxLRCeyp0XkpD/3UUcF+cPlaQsV0l2nnTpnLijuDn3enAaAntRE+BzUd
+V7TmCZezZQCtt1KUxJZlBiZuxAA+AXZdUU//BU1q4Ph7gsaDkRUV+5JkOhB
3MVFgcRXxXC9ZFS2StKiZ7TGsdg7ejJOqVPs1HG0Sp5YGzCBPAlQmthPJjAu
03iw+l/p1KXaHvM7ApHjBEIY4k3K7l6mRlSyVzQlxbslEVWMGuoPu5i8LRTT
P0jsl7Hq3Lo8j5wH5HZnD08jvzsHD03pKI2s+r1zHfiK4tNXj3olYbDp0hkM
X9HkMW/n81r32kjV3oPLY5/REoiIOfk4Whn2PIPqORdYj6qTC0sXM3LOdqYm
fbQXRHTbl3ISLoojksI2wjSTES4Va/awqiIbdk+O4OqfG+defMlhA7J5VUKz
WdI86jHjYkemUbKh7bFBzz1nnu6dBJ34y48/G+WX9VPLO7/t+DLN6D46zpCs
mjktXTLAzYHPltMluxXK3lN0GvxQngE2b/V9pBzENlmbAK1SB+QYPi0qQETu
GpOCzjgaks83DVAI9P4C6kcl+6TrNOaP0YjyUk9FzvJ/1L2loJn4NJ4FL1yr
SZtCSZ533VF5r+eBlKfNklzRzgqHlbo57Qz8zxpN0LorYGEN2SmvumOS6BgO
o7k7a6v1NcL0RyIbTEOoPDQyaNOLeR8/rJ3GY1JR9/6+rD8ON8QIGN0rIXP/
J2N2h2cS0tFBr55kIeFbV60QK5dxDM+lZJiRtc2cOKSbTuTawipTZO8T5TNN
QNhq1UMyHHXKmWrIWeB53AZpjPUzi5YZmwKR0RYFVIdiBMRl+94qy2th7sSe
00jKE4yLoKI3Bg8YPr+NjaIA1RA+IDcEjdKtgp6bn+/OR/dXLxq+IxIwyv6t
0L2bmu2mzCzIY0BX89aFoVQhxI598nXa/EkBGdQsmBNWRmKUlLeIhML0gnwQ
iDiSfRorG0i1UnmsUIPdEF2T7j1tnPC5TrBCo1yz5hBcY+8jLDINd0iukwU/
W47Op8l5dbYzTiMS0hk0CIWbtoEbs9h9R4LE+b95lQamZKI64NQZxA6CvdWy
yqP5qKrEIrUONTA9vqqrQyPr7nitnvHW2TJYmf36a62RqmVkaxD0gtE6cbLv
GsK/Q/9hQ61uEoozJstriAp0l7g/h7bRqNu6P5xzjehaXnkGbnkp5SeTbmu2
Pv5jrXMgoPubcm1g1eN/EKxIwjW75JgRUvPc0W1/jtEJEbB70MfDJ549BIl8
YnzPj+mozp9Wy4VUl/XQOpRn0290qq1pijdBKGgsOI+ZxuUYAalbriA0Sbse
admXyO1w+IPY78bb8kMRiMWG93Bh+I/+QgELMkkNcuAMqVITxb9DkC72YiXR
JLPpnX4W/cUsQC5FctGgLiiSYN7PcPToY3AFHdTn96ZYk0eH3xfI/tHzRhk4
gmHwg6/tSp9J4YvS3cDgsTlTfdBQOEwpI0wffKJFAx2vCyE0fgJUhoN9QVUL
CcyevxE4PgPB+wbHzTwJKq7bBeppdP/WyND0RxgpW/kfGdRMfbIJkMXxG3zf
if+bLFvtpIV7LXK7JpoaF7lMpfTfeeNKylpw8M4pwWvJpEHPbJrMTKaC+VDI
ZvHhCnmu2+PEqdjRaNXrmyaAhmx8MPjAx2gkr1xHY87Xq+Wntbj+D9+JBPU6
GgnbZqmN9pzM7Ii3enXVGpPgkOqeGWmf+zbwz3Uq9SSt58qBAFeyWY/QY1dq
naGuQr5T1Qwgh07xMOosSOIY8hDr8NMNWxZlRwhkMF5Lt03MrPqeADJYkhcX
7jtP/iHJMmTO0US8YcoF5WPDxzVOmZwcXHypRIL+M5XKn+WTd79ZqWATapRX
sGckyPFhaQM8FUXaDXBy1PQaoh2sdXdzo+YV7IArlK/W/LAITcBmM6Uq+ot5
A4yWHQ3boXMGHqF5UCLDWvxmYMJ9HzJqRkWLICI8Pn6MVuyGfbGwmq03h97D
iMYjUol8QhBHfofiQwHIEH97jYrvTWk8yXV3fShgQQpQsg5T3qySk1G6LMWJ
BRzkNuXXUJDn4QHBbSWVKF91/km8nMjb1uNjCMmEhYrRGz8ktCfni7vENRwG
4WQx1dOZaRjNdoPKe8E43ljY+KB39EyqL2WfSux6SEe4EJXItyg6wWz0lZPl
B4Q41T7m1df5phE8aEsbVAtAK4baHrhmMauVsuiFvOdh5W9iaHob1+eW2nh6
1ScfqKEOUSnGivylHJ7PR086/9mQWfbnkCSY2sYKl53X62JKF56qkmWuwqtV
Ks1ogyI9lsLi7v7mK4/UWjj2lQnWezfzK0q9yHb+z9VXCTkYLRhikkEUBKuD
9q5snLliRFehldKEvknAzifFF2V+qxHzHeKOY7GRgDZXqXEV8cKVn142BNfz
bPgpAUERy+oxi/vnG2CBn2hVS1zhvrHTF9nubFWv4Q2r0+Cnr+Hqvlybx9mA
+3CN2EeXcoO5O3vJ4l1NO2PKkPJ+JzZxgVg6MgOJPy6YO6C9oHwWh9c+QX19
acQSqIQtu9R24UTSPPENLsD+9Fi7TtYkU1/URlP0RMmhXYFdcwuUBU0dBo1A
Z+cJb342CskujCjNjPsOtp44bj7Xn+eYwmrHErsGxcMosdh/JaM/uKi1lbPg
s0Ef1lRlK8cEVdjcYs/0bPs+V+LxVWBTQQzHahz0ftfCGVU5unawUEjU2C+d
0JX1lRMDNehWDRAVkw+3aOdzVcqBIbK3csdZPRVTJ/ifnnBVSOj4t2WQflyD
aUqKsRmoKapP2xXC5Jod75BVpbKQv8s6mnjCUEmhxwYMDDW5rHZ+UP/zjHWu
Ud86vBev4nXXgY5VGqZh0y8U5k36f9wqv1l/WMK9GOCKssvh6oYPHSzYuwO0
JKPacARIkzj7DdvepTLPD8GHiLuZifAZUSc586G5kx995e2dVV7CcCz/rdhr
5SyJl5P5V5ia3xNc0+Nau6bLi9XaiB+Y3cg/m11lHP+fKj55971tOYxT0YYC
qsCOCwiAR4nsPoo4SdGARqqDB1Efj3Ng1bu2MaYFR9Uvfuv3XYjeAiYUtWB+
JIYA9Zx5Y6gnU91PTQHJxizKYkxrarPPoUd8Iu9WwOISUazfdo/3SA22whpD
rRGLGI179er4tIXyzkMsenXt9OHzSrj/87REhHpSGK7UofmUNrn77HATBrXV
ggdC1kKbiI51tQ2jQJpNYc3u6GDf/3CsKWJkkYMUWke8QafUjUzf2yACoVNx
kgKtJD4/wxDZV2rG24NiiTMfjwrlWb3Zdq7GtMEWW1zSCehd0XDXPtwvyWRm
hT4qx2kl9WNVbrLkeh8FHO7mJ1CriR12t3/PWHf+IJkilVFR3jBAZ5wOcT+c
CGSTqstowjzq+oCoC6Ww0iry/z6ctkqVRMNYdpbXs8PpwnHZmneEjqHO78bS
C+Flj8r/MO00c1nrAhI349ON1f/5hGfHddpa1hM5I3rjMBx0XWuwi07iYaYk
1/saSm9zc6pvnpGoIwc/B39xEzV47uYVG9XYcDO6zgegmcqxzEnYt6EtenLy
0wIPsSytf/LvYvzmN2ukA8R+BchbLUrYqI/Sob7B0gm6JDXpD2LuRgoG3FKL
y/KQcBi6xRJZDEMTZQ8Q33P0+WDSbpztACIuOmvR5tzOXLVH2b238hDSXoMs
npIOLhTqlSuNnzS3+brsmGd35uO3lpawlylNL4rTGxhywIdb13X03e/zUHOJ
/feAJOvnpbmeiN+9+Pr5Ua5LI0ggFsrxBsJd0evpVU3C2onru7y0LsPCuxJS
iiM5bMZUtz2uGADc/bWq/B6cmbkc8f9VhsJydlaiftLPzBqhBvIBrG8mjXA1
urEzW/2awU8lqEJSH1HniSf7E8E2Gg7i3ca0JEiM8pt3hElgPcvK+m2cMbj4
QLtCOIxZep30nCZESkurMaS5yZXJL4BWmZf3keLCeRbUaZr8LT4tK0gTz23/
CkjCptQ3Vv5C2jgS4OPDBrEVdrGTW9UXiQwu1UFLwuwB97bHBhwtPSTvOG4W
wvTGnjucFpqKBwAkKv3XINJzEWZQuT1J9Rk5eIWYNXAE/yRgY5SF4fxcsitx
ONKW+J35eDB4SCTi9dcAA3xbaWCzTLUfu6ZDSFftaHZwaAWsOw6qhvtGSJZ8
sNA5RMYKfmLMnckZzZ1iqY0/n0ZkdLmFyjfVEnXKJwqk1ThkdPgq5piDNwmF
FwSOX8NNJlENEDulNR43WKziYqW2vSQWRw7GyZvbC5R1YhGBcI7mHOIDay8w
CH7UVgpAtv8V6uEPboFQWCfl1Y2LZAzoezX3NTJOFXASPlflq7ENER9RI+4H
YFQ4UL1A4Hgg4nF3u+P2P2gp/idzAyHEUJfQeWk3IQnGo+V3pvXloVP5xMdb
QPsp2cGh1GqVrONxeoRHeX6oRpiEGtEvKE7ZgaZsbo68zfd0XGpz27fficA2
WM4b+/DSDRjDPVNl9aJtYOAY1Mmi17z95jhd+Ta4uexPlcuZXE4uxQN/qa5m
0EVFtOThKcHdlKZ0q0JO47NWlYEuCRwh1Shh6SgiQWqb0/QSWaIXPEhwpH03
CSCK4N2mAvYgrhW4O6ZnsmozxOR7y3+bksX4BNQUQwe60BkILL5j6Pgex5hT
mSPEbs+kP8RlFRUhYmO7IEdypXRLvk03d0PmbSRfLDs39/C24P1pAmHuZJp4
3LBXmivaiJuoHijz+06Qyc45VhKCq7TPxoSwQ32G7G69QSiwe7RoV5knA3Em
B3n5aTHtfRbORpGNDyuUQfcPB89qrbSACgOh5eCL3FW84JyqSmCi2YuPyumG
VUpaPnadbHYY0KPo4rVRZAMenfsn5QGaIO5Bn/23SIflPFxHTl85VP5dxJX1
brJLSPKmaDcChQKL3iZTmkXv7MwQW4wvuxSbQxPrwQlR/asqz69ljUktkz3d
Nszg46AaWSCxndXAQCUh+rq6gRnhGDfPBSq+/74u9q6rzPVY4jNMegqXWXon
3KqPRjIW+tv3UZlPIid4u5UD4NcUedtNa5ZxyY35qcM4KFNq3uOSnAtDFJBW
rrgVq3RdyrsmGIPZ9x3v8Ern7i1Vgzz7pqdN2pkhWYJeTMDFvFJPDzS87leB
guM25WSiCL8PHOQmgF6uVZlcDV0/yPInktkrNa/jmr93Iuo0DMY8lWC7HmBa
w8cN8QNFejYs5FP6jeUq+4Kv+EmgpMXJm1V5SQKlB830zLwxL9VrBr5ea3lY
Zch1paOYLJ8tHyv5sT7qgdiRYYNDf1kK38LyUiIlxdnfGuzYwDYEPK+4UT15
R6pATVnBzlsgx2J6k4Zd21e+Dz3AsHqzZGzWBakEyZvaAdUiE5oCi+h4/kQi
zxMpOp0yazs8dfC9aN1vQZm4MOAKIHDUDcsE49anp25xnNag5XPcVZgRP6nf
zzjHiaeP4EvgZk1cqnFOeq1nJFORetcftakjaB6yQZlEXzvI/dytWb+dZpPz
IH9J45RqhekKg4TpposSU4YIUScfu80s0WW0e7gPJz0x57mlxmP9+zMhxC1K
jSj/1RCecO+NjlsSIpaYaChBAxh0EHk/ww1slTnHmngVVegUe1ST4cLh/icM
ZiOqvY0Ran5ez3d2Lgr38mlxJ1hinmQLX9KNodZpAE2bjRVq9pVbp7L5cIvf
hnX2RtmHF1J3yy2mhyt2Q7p0QInqNAxVmrJfKa7DFATUCETdWDstR9SdrZ5X
fV4OKlQL1dVO39CJ81S01T7KFIivIgcD7ZFHiuEozZUuX3rrZZaK9tAHl+cl
3w7sWD+hAf6J4WbXM9Xl4IRdmPs13IU6QgrIrYr7AO2uS4f2MjgiW/Lf8mCD
7xAn8N+6zj+iwT99uYWOuGP1e9sJ0THsQHyZ8KB7jzxv5T9GFhp91YoLZn/x
y7x4cgeALLvb6880yqUOFs03zYTnkfsCwcEWsKYIlJIgyv6wdc/kMKCWAJfh
Bsic++v8hfRuqaxE81lN5mUjdrTurD43XevEqqVTUmhwzq8aVoLbM7YGZoZf
UP6U/yRYoge2C5rvIvCzpGXjGenHDFu9sGrhuIJuul19srxs+gHlotuyeI8r
EbE4HbI1Zo3FlqmLWjJZ1br87WbS+mV2somUrE5JTfX3N8jOSEZ/f53DoFk0
ea2IEPV1MiwvFvmOytjxdjIzdSoW6jeIGPWU7NgV/D4hTGka1WE1tT+QsGTt
oOSdtGz3KOGRSTLQgMxvbtIBQGKVfnYcH65PtWd9eVynQ2vDMV6lFdQzvf87
h1Nbycp/57Oye8ilNmLdWufSpGZ1t1tMZrXQXzWl87486jWvyflY4BHU8fU7
pX+S9keoiOJn4Zm4mX2R9ho6w0wIAtCbnZHjee5ARjXRhQAhqdo+c+Ci/GAE
I9V9O8O1GhjlEUVXE0hnaCMDqvMgpLCKs3lhYYp2I73esDZGlxsBMbL0jxVK
Jb8uafWtb7cpo75uzD9hbFip4IQ2I0UBCtcc4EXgRiyjLazHZ+sYWJewN+O6
PpGN0lhJ5jlPkNfXuUqhVuNtxMknxU7AtTIvy2zYbuJSymps9Wyy1NAEl05Y
vqX6mYfvhWXLtpGHr2/pKFNUVC53vlWbfOKD0rOA3NUdH4n2ychTCiH+SES7
u/cogOA3+WMEhWmGdEVvzgN0J+SJDU8+27IAD0zjDF+yqkb/wlK4fQFPETQ6
RrHlZrQdXEDFAk10p6rvuJFDN6xFfRL3ZRPgILRHyX8GNzKZDsJ/fUN3U2IY
90cqECkRWIWC1nthp+mj6gy71fSVGxSzM7Ds+SAneu/Ac5oj+kLCi9vbupjc
dVjI0JPLaFx93fm37Dh2/qKVseZoZIjBSJ/niTtUzL4MB/dxUDFfO6ZMfXi7
6d13CSlWI2ZLk8nEYpQxNzr1L0xc78z1IYRydDXqsWlLWnYpMbhGUtd/Z6Gp
/kAsfPwIZC4JaIC6eA5WWRbtOu3a/d7R57ogNrZrzskvzXaWEYFr+GnaM9YJ
sgXTpuE5yhBPQOSTjuw3QA9sWRN1lzH6SZ3frjmBPFILRaiY4lVbZtMG3i8Z
BEs8VZBs8uxqc0gVRYjsLZlOGigoV0hJZzuIYmbtclo0mHnFCwtMYxmdgOXi
IBxSkIDY9dSPK4N+oPXJY+Lto7Z3NBTomfVoDm/HhPY9qL0PDHHs+CENBx6p
5aqwggOX/PwPVr/o6msWtCQG5d3EeCAY40rcHGJj15OLRgjlZYPp43DvXc29
hVPf9zu6bUpnaqLOt9WeC9xGoB/quUB2bBABCQzYu0x2P0/2jb0Y30Oqbt27
t8OH1B104SNkRjlYFgM5O9QsEiv0u2A0cUNhwHU6tawdszCOh6J4DTXPeadP
8mCI4trmGFZSh8GEtFP6CXDTbC239zgMsdisrX+GEwac7XI9gSMGoVRk5nVi
wOIrHLL87hMEV/IyU/KhUeNhzIWXNNFInuGpMx04n5D2fDWGzR8UICkT/bn2
nm6cZRdNT7nAevQNNUtjnnY6NLXz0NehUwZfPx9TzI9c3WrxsXBSasn3zBwR
liM19CFDN1Z+uDAFnchewMi3le4K0pNuoBFdtR+3J+uUG49LhnCorUcAulqP
2cD7PdU2zq7D6CTaZGNqyuKLFwupg2LZAec0NN9l1rttQl0rOMg3gEFwn59e
4BzIK88VfSTht2W3+8Nfn7Vq43gjPdBAKXLcpMtqd/8DvGS4x2B3YlBRTabm
RtI/D/mUmy6Ja8DitsncVzq6WctwG2+Nr0bYhxJyF/Jb+PTUyV7i5cDq/di4
IhIAa0e3suS5b5HAcJuguO76NJ7u5IqUH6Z6T5+mvg0ELj+3Gald5XEtLHRR
F8x7rCRe6Clb4mC9AL09FowYPFXpxLftKh2rECxOMtSpqeO00TIGC5jr8xwL
3q2f9TfNhE6fbFdAdqfhmPRKgZFDsz5QC7I8v3OnDMDbqYMflAEez9Od/TwV
niLeeNoRpBncO+n3dUqHm7wsEuMrDS/cyut0EmKuHGQb3BbziGhyCNmaxod7
xzGl8gJOPATp4TzGtZ0dEKHJeRlfOqtKSZugbMbiouUGv7KMot0aB9nfP1Ku
HUzDu1J+yhCJl6jtGWhE93F5YZXgIVNYL6efrfZQZsHvDXhUUeZxq/5EtMtt
0PbBdOzbfPaWhRdZgnaNcOip4X+WO2tw2oPgMeXxsPco6R0pd6agywtAyMWb
9Ktd/qktgKb+q59YDVxodJz1pVLNLUTy7/HYBFn+9w8Wc5UgDx96p3C8pWq5
rfwEBlaF0d5j22K6mA8eL70Xvhgid9DI917rPa/jV5SheEpzr93MDDC7rZba
/f5d5lCYVOVOSbONrDjSFwQ82cpFc+jnl+CRZga9bCZCFWkGkrU3/H2HvnYX
x2I+pu3w77E2HEEC4uNOsyCI+WvH12krK01hH03GnTnsdhHdiZWwmoX4aKVr
9k0bXKEyk8wDR3Lft/cBwDUm5mcgnkYVWvmr+pceVNtDglTXrHDVJB0No8KV
AjNKcKX/HQ/G+XOxW/ZGsQlVSZvcE3YosQiV2FrcLnvzE/uE2/OzFr9/7ph2
JAn7/h/vFYMX4hgoIWGecjMigJJAnmhDKyxtZd/nJt+gI67OLW6wA9slMWl4
z9P42c3i4uKJx0sPk3OeMUwnXHJQN9DuHUky7yB8FBzI8stj78H2ujj7QPCf
9x6EMVJ6kYsbguWOG63sNZbgbk14dKZ3KBtVD2LWQFqDivoK2RPIeh6/hXFZ
NNFJA0wc8eludQ8MycufwWYoLVYeHXbJReKRQ/xcfiDEwbNp31jvigb7DF1O
YpYmRD5jG/G+re+X4aJGiPG/Uku74mUCktwhbjNHGJ46lrSS4MJqfDtmRH6N
FNJJd0eWcBJHwRGVhg7ZlpG0hFxreHT88YbRDGlikDmKrWFy6Ndxilia5ABb
/3u0knrccHapq/3uHNehLVrkXZQgfeFBwP1poeGg8RN686PEO1+SEyZ31cKC
V77BjSnrcVULWljaEqnQ7OhU51H/ROMY6ozs3DJoQPoNUnuBAdT17ZpkvOkw
wZhyqwqSx4sfBh+7kj1YsGI3asx7yGOjC52dvkxrgJQYCLainkX7KAxakJ6S
0fjWkdTT2EuWAbG70eMOWnfSHJgSHVk9BjySCgYkxYtYG2f7VmCKgSkms8cs
RRwK06XSRv185+8HOyXR0IzUJBcsO5AkGbzPrPGU355D1gvU/WEtEa+IkSFB
ll3lV9CHXFVGsQ1AswEU8Ef4FDL/0D8PRGCMAJInvwB1huHbUjlD66h61Zds
tILZ4Fyv+/jwXYGQRr7Vjo8mLnMBq4HmJZqVrRFttJuuvi9v5WyKGIXld9e8
2+Wp4urBdoBL6XIayVXPSk+z7Uk3QCV/LVtLSwIr9l5uMnqjplFGsxmaHFu7
zpeAKaaDGGi7ac8Gvb/+9QOe7xIq6peV8kIHAofVZUIfptA/yZjxsv+qVbGu
7wSc4sDl57jWiLxAeCxrORVdcb5or6kFgozVWG6Juf51IKroP9E5hLO0nSil
edXT8ursKXn5TDjueKcblB31lkdTow0XC7huVynFjpbPWtk5XQYdT5H5CfdH
klILMTaaH/UcfsolGzkFya5mB6rabdYNV3d6ykbmSgAqvE3a/ThgHpUibES5
FMJGjP6sZ8D2g8+EyWJIjbWvKlI9U69iFxJKcGlJ2thTy2s/zoFFCopbmunU
0gfDz9a86Pil72NjMPDZpNGkt/9kdoKLWqW3rwHQmRpEMpJA1B4Kg/SqIIuD
D2GYqPraZ4hBdOuWzUrii3nB/MovD4R62O2w7aK+Fb5YZELaC07xE0KVa/T4
QIg0DDrWedgCMtzsK2AB2PZ7miwhc7RxKtrP0miv9aq6DuwuJm1LJ1c8GS8O
CgKzWJD0Xc+bUBcY7T0/GMfB6m3zRMXUSWUM9s9hsVbEnEVLPsYs3jLiomyf
HoHmmQ3lMJpTKKvfpG4jvV1T+YfQr4sQSI1+E2yJ/ZKLp1trWFPDDj+qwlfr
qJz/lmfOZYk0gOaURDSUaSzWk23PZ1NahG6Ac3tONNPNQbdPoV73q8gbCfuR
NFUx49lSbCPFqjVaLRLoaI9hIftDYqNGpMwvy8syjcgTCLF+pckVaOS+Ju7Q
uqwaecl8iAbaSQKIe0vopFeuzjp88VJFBvxyINADovgfdBPYmS9za7i07dlB
GQkJROacFlvXnebZC8HqT69k0fKlfvl8Hxpp++jICoslWVLKNiU4031TUfY4
tj+yuDUSCWnHtui6Yq8KeV2h1pMmTY+lwLD7O07F/SDROySQ/99xisVjD1Jw
5bg+NE3rdn1xyYjKhDuKqpRacVc0KGp8HtuxfrrBSOjO83L+GD9OqwcXcl1B
Z6mH5lWYQVkz4ENw/vSO45YgV+f1MgZHEMpeZO9IC4ulx6vfcPwOlhgRvUzK
WX62fN0Nxx31PVlXGPeer/Mnn/kUZzJTSMXyA9krCxow4EzBWJbStT7hPGmg
o6eMvf6sYjj2I9RzhTeHr9NMIGLlOXHyagXw4qsGQCQo+8I6P/x4kstd4H3k
a9BoNuOLTzNkB6hT+Call+GxHhJfFQ9bWiAAFHES5Q47xCQIexM8Ucz1+zll
9Yz//GarGOVv9N21cqQbb1Ze2YpgQK+eqbG62HqB7sMYjmymKjzhvK/rIPU7
0P8m1+npuyMHmaw8Jl6/omSRhdSqHHveqL0LQaTILTgM0RAHmDmJjW5JGsCl
4GxjB6Aus9IE5joUNYEz078Ko5aeTIRFPMNgkch928E7srw0TS7dtWXKN4Kb
P4v74w8+c/PPYlIg57hB9hn/U2oehfjYjeenIoBirgpxcAFqp2hID+IddYHE
KTwioWhw+czs/AuJf6wWrr+ikB/QyolO0B5HTMkiXZ4jCeK0BvJzff8K6bm1
Z/VtzwovfK2V9R7EyhENXQoVkUFDhzpzPio1zyBdVXYhidyP7iG7I8dqVxuO
HWPXXJp0wZAOG/RW23neGNwRuqC4m2UySE3tzVDL6wl+i9db5B8//dQIxeJZ
05tBTzRmda4Y0CrqPp0MqUOANnJphPMXUzryMkGNOkoPQpjiuYZYmG3GeydK
YzcE7e3uf/oq5Yx3UY1CAuYd9OjrmRsbDLwKkzPQyp5AvLPSsLcczlHFzHoQ
5XW/L/aZW8N979v90cJFsJGIqWwQ8shxxUQj8j9u56n2BXhxTuVC9nM0haPA
WsWnWIiJMCEWvBcpcOdu8MVitYbnKWvqTX7/3OzKykG614IR9BRuuNi1pZpM
/JAP0DJe8wVPjEDudrKB5YsSx9YaTcyutI8MHxPxfbxfiws20Wv6LE4bPdAF
5E1r+fPa2aSoCFEOJGMlLDmfV/mWMYB8OuStHNYOhTXzDswJdrAyNI3oxKC8
fqhfXVHtAEwDAlgBCwNnhagu8UJsVe8g42PzSzf9T97aXzMsesMYBATDPgUy
Eiy6yZ188fpgpCUc5/0FBP3T6Im6Uc8iTexvTtieM19TlI/tS+oVE1yp5ukh
uPfgpnQnKcAvdJA1Qeom5FbyCpp58go2dOPRnDU94Dv0iOSeVHOd6aU1KSrH
RKRmZWVlIAHQ9FReTuHCGmsKE39oIDL36WSXveVJ59Zb5WgsUXU83ArJW+yt
vUvy6+CKmUvvBk0nzhaL7+rQt9EmxIwLlnSyXV35vkoLYOSp9KJTCfXSrrxe
TsucSdp61BepwwTERgKKFZo4Za6HZkucKFJdUrxEp+NcXXW1nC3rmKPLq7BO
OBJQxd3tjcFvOU7i1PJaDk+oenXPKy1usZtksgjeBK2Ua/GNWyJilbz8xU+Y
1pLlYKWRAY2z4dt7tsvuxcyg4g2ltY0uYcqTuKZieaWTYQEJozLafueGLaSN
GpeL+yWddyWFyfjkcTrsfxBuxnqRFVBXMiixQFDQrmontSqlBdzz1pYTXu1Y
ZF7AEU4nU37iU6AQI9XfRAmjWF4+hUAFlLIi1u2bIZfCWhN6/OCvdf1LIuea
lMtec14QJy7niaVJ65JJF6icGpx6W0KWu6b2zzPVxgUm9lJcAAzEazuAH+Yf
Dpe7bf+sMy42o0p+BSYBovk1+d1bMzZfATCbFrKOb5sq11xCdjE+bX31hrJi
tx/MJZA0WFHZcJJXw84aypuclrg27CqcKOZ/h/7ju59j6eur24xbu42rh1ER
DRawRGvigV4uSbtG9/F6uVSlqsv3i1UJe8MJv/jEj6uwa4cX896mSI+pYMkl
arm5le6HWbBZHYyp9uLmLUS7ytY6AxXTQz+fzSJ5XqJ5vIUH2IWy1oO3GbJg
NF/TsLq8kzrtMeuVJX9ffQ/lYGH9nxy0CEQGjETPhiOAQpIvR3gL7EX7JYJK
WLo7LtrMlqE+iVWRlYosXRBatweD1HhxCajiBAbmKjriY7lh6KNBBGPmIvvt
D7BDsvoQof9fGlCk/3Z39lezvaGRPdFALAeBir4fsEMcKGrKfKBelwX8RtrM
nYelZWzq4oS6p6EcnPqHV/MXBzvsqRaKkw0tIMUjZGjfSsLrfapmZWv9GlxZ
w7mRLOuzKjFWZo2gtHL14yNaIHrKlOwRkA3VYh0kBUcyEgtpb0e+Wx8Xwtok
irg5M9NUMdk7cOXO+Pmmq6Lev6BoSr4fC4rEKr5/Y+XpOXUTm9PYhNWdkZX+
j17G3RfKfZVf+thliz/RhXmvs44VTUUL0CcBxskqbZOiDHEil+VzkVvtLtcR
3fTh5Zxa0zDSptaCmtv1GFqGpuJNEWb94WGZ39S9jGmCGyH+Sb1S91t/nIK6
84IWh1Q8TXuu6NzQOau6UlbLYX/2HeCrdGEHYKlhcMFHSceuNkR6XGsShINV
/y7U7scIRBtzOh9MQDmA+g3GK0oIyvS4/wcZebv9qUjwfHy1vFq5mnqe8XPG
7ulPgzQ1U1rjN9fFFdVQqs0qYJcVtBKxGDcCOl0Y0roaGtnd/fIBVKM8cH1U
5FXqQiPs1bL5aadaYSiHFYDzst6su18ljN4ka154bbiPzFn9eYEGFNo2SCHc
UhLJzdWN1Zt8PkS+PP6TVEOc6RmlfsiQGHyj/9+nsxXk5qk7N9x/gOzDH36D
9S5pMZLgK/HiTbduR3/Y1Lp4eghUPbVr1aXTWpCuQfIAPNw2h7/e4vjbSt0j
C84/IlBBSDN/wm8U4M49H2y/0/mePvBBl/Nb8vMEdfJVfPEdn0X5cY0ddmXK
1xb440gZBVHJK3t1AbSlWW1B2bUz15kVnniYRBUi6q0Ff5MqOmHkoLqs37AI
iNMRHSjYTnTcHtQRDSD3xnqvroxX3zak4rbGwD9EtVUtiPLhrql16S9ybu2t
pb/8fCTckeqhd/B1kcf1/G4cB8FWvPCrU4QkduUgFBDuEO2OX0MR3W+Dl1Wb
wArptyKUOigZ0JvC7XxoT68t9UubbmLBcuKhmuUdBxfDP/tv3Nxa+zpjLhkS
URRXaCac5Bb6V1ZDuYJECPNx95BofHAkonx5c7ZGQArxyUFyrWyhzkzIBEyz
yqEY83EfF1vb/jSoUeo2as7uTd32edKTYU+LnZLAYiPdB3O3NrdN6aNomY4G
15szuPZRUGiJgpcy8qFnmU9kWvIgvyZyirpvnaLLX5VZX8kfeKUSMQ9/ICNc
5xEFOOKZ8fyaJ077USh+UGwR7G4QFW72jNPZ4xe1XsAp2g1VKzAuwWU5NDKJ
5D2VHlH2Hi9IwtHvgdXDlbB5Nf3qM7d1/kzGbvM5Tg34nVWDDl+byTkLV6bN
1UIPazwSCt/ljR+4POP1Glo1gjk1R6T0R6neoOecrHt1twHy3QedN/4HolK9
xdNDpzE698uHjBR9/fEiwQ6JFB+Nb8FdUgjHeJhbpMqMx2iz9dgybGjjrddg
Rd0CzS21T5g90+o/Tuo3OSFCpgCrJTw4/eo+sqv03kmwL9HHLRHD4pYNufrT
6bJGqrPKhjZR1+F6pbp6uCDpzDsENQaR9bKBtzRBlYlD3EBg6QzEZHbctTSm
BiWVZqXyhDOOsZQxRQI1FSWhVxz8r95E6zxWGxijSQVndaZgY/YhJZr+3SFq
5jA7/t4yzpD7M7fA7HoQIZyIZgc8o49kuKej8UhnIDpteyl26sZMTcwk9mxd
VNyaloBhcVur3E/KvqZiX8docCoekfraSRgb5+cUa2Or/idXN7YK1uF0NEg2
Kh1QEZ17cGsDBKOCpgHMFTMHfWNYv8LLBDx6h0Rar0PZ8DlX9onoFiRsCrTa
kHsGPF8u0PSC6WaHXdJ/DiTLKkup/jECYjlFDlVF11KpeHFedz86JE2wYfzc
ZqmwkeSt6m+KPwJzrLiTM3punxxIXSrdx7J0maRrmOkcNnYnw/kaud5ApmN7
7QI48xSgVgcLmWRmEB3sbsT7PNIR3bUh7xLjWbVWeRltqCWNNzqgNn1osQ5Y
EZCykrAZD43CCbWbuTuIx8ylPmUg8Qg4xsc1Dohc+hCffufTBYp6WCU632a7
m9btfCe/Z+RE68xEKdQC4AZFOw7rUJIbwpTT4cyAv58pu9bmQOPsl5R/82/a
7k/wyjJS0w6JRECkEMzMOEzGECIGirc8PfJS9SFDCSGqSIAZsTx9wDTpB0K5
IvCJNNHQszJcadCxwVgVvutQiaStpwnM+k5DNt4CpxAvHDFAaIairOzORdHl
0R2VFDMr2EUokYxXsz+9JWjJc6MM+0xd0u5tKw785U1ZOFncqFv6P9O3Zp8Q
RWlp8sUiFh2Gv6VBXF5GTSA50/BQw2XcmsTl9R73icU1lI0HExZcCEXPWL2Z
QheqaaxbOR4skP0ZIlvJ3/03nWr/HVtfoxIATQkbif01OlerrvBbmp0XEqsJ
5qSYEr2GqJinB3HAQ4C50KILsN9D8bg9csuG1gq/uAp2KfZJ/Yylkn9W/KmU
8l1xQLch9QCEMpwq4tC5ev0/Ae7YLBP+0rdrwpN3gWWi/23zP4ZVRsKQ1+Rv
pkQ9khSw4RMLoi7g/x5imhBs+NMUTGSW3abYpP18O7vrKnGu3WILMFlK/0t3
d5wtnJcpgZgykLQm2AlOBOhPs5sGPijvJvYdgzc6ZZHv0utSqOSPBTLy3d5F
waNF2+oNF1S3ScPUeIZOBWSjhbSgkcsPWAA0M73vWOIJN+8MgGOv1+rM+iqA
cZ88HnEK1yLfHZYrdN96PfL8eAJ96sSmNDhfP91vm7DGNjmdZs0hyMjn15c4
dbNZyVE+EEBJDN7wTCJe7nzOqGGzURZ4ixxwPEtEAPpPVQsE8jPsFtelzZ60
lRfqpHWI152msZqDscnXRZK0r1UOxwm2zqq52Q9x5/O3YYUxU3p9cY1dgCNB
YfNan7/fpr6kvNBqLai7gIMiDQSR4mR5SQhxRdNzmhr67b7EN1rGC64jefb+
pr+fW3LtIe7y6FVELNXLY/pZbCR5P+YQl13pXPm5Cc3yof2bPA1bwz6KEe5X
7yyLwMWdMOf9U3pHaShVu/6zphZZJ0dSmc7YBjgwVS17vuoi9Fqk3KVtvzk7
Iw2vGXgPpe0VXZqoOaq+B1s0MxjYdXpCjhDWnpoFdPS4jJE8wBYlMCZqWZ0K
esGnu27YTSGb3bjAAVwjfNBQT87He7epe5FnJ7IdPezINiiYZGh7Abw1ZguA
3D8x9nb4DcsK6YVWXJOdmA4NfaCIShNN9SFp7c6xj4xbqT00SK4nbevm+1gt
U5RWgRMq2XX/9UtxYM3sJaW5g/Xyy5FVY17YFyI6rT2K7k/4RRRBjg+fx6JE
B1qQ1Mg6Hro0ISL17L14zaSWZHl9YZ6vVfZtdGg+vnfzqmnUeDPBjaWjHAiY
J4hn9c3mQR2+eL+1M363r9v1xkJYzVB/kQiIaptF6QZfcD1/Oz0eCOcRD/5H
EaYb0wUm8bkxu3WPdkVHzuf8UQIsYeP6o6bDe/2Y366iKhzEmeYSmSfqVvhY
Dd2mlwwRQJjBxNjnhcLEF8KAUYxZ7R+c3kZdeJy1vIhG4Y3PU+ybvcHG0dl6
ClM4bQUgEgv3tDD6NCdtvdwDKYC25Hs1o33t8AFgeIABGEcaZx3QqcfKqbvo
q4NNNYJmrQthPmCAUQAnf/fmJT8URnOjnHQ7k+EMwvPV6pZSmpPYZzn9N2Jc
F/NVVkZhweWxUdyAoLcNhDvMlpQ2wXEfnHQyiEqYF4nf4fGhOl1vGq4EhiJi
3f6Anhv3b2jbEYvJucCWwAKgOpouyJ2YNTPDnVU5K6zYU2pXiT+/zyoiEBv7
H/ekNE/leI95Lk4xtiwlvYR1m21iEvYJwlUBlMnlxMFOoa+iXlR9noS/vQZi
AFWo1NTHxtMnKChH21JLtMaLafVfOjpFAce/8sDzDYpDmxWARLwx1zll/U6I
ZDO4PpCcof8O8uW3nKKi05ye3jl+CwRWsGlcBJh/56oLnanHve+rixijp+iT
OdvfzukLBGappOPAfhHWCVryLTJLuLFfEQ+SIwgILlmwMQjy6SewodKZHBQm
/QYMjGa0WAl7mqBKNHu+Slmupne+ELTwgIZG+MP/eri43yEOwwBPB++zRGj/
/lbjggk/+G9tPcrkezxlmBVbyqQwjhj6HJQpU2RBwKBnUDzFR2rkJlZMI6JS
xxoTFIv5P+dyJvgdSHNeYkndVeut0NSJZ1YfqG1RNC2XldTaPU+JKdQWRXkp
XvA0ZjudNUztU79iGSky80AtnN+HtS1h6FgDLn3D8KKjfnGIVPtYCG4jrpFF
+YUyye1S7ZXGW2cotgFoTRUImJB0HrlBo32xmJApRmW1GavRULgKrwKz5weY
dq8umNSgjkjZMhwY38aS/bkXfT4BomPl7xbiYwb6n5EHBznFaXThJCSVGVoH
xWuK8Ut8W+bCVIWz5YTbA3T6UZUxZb+6gJk+pK1SXXrLhIgFjqYPTLgMOQLK
2TMYhJg5vkWHlbQhJ7MeOhJ/VZIJaGaRNDtLb5lQlw/8GD5pz66RrO/EjqK1
ubnkQEcJ3ndGJYuRU6FB4gJr0FmRoPrgtgdr++rsWPZkaZZiUUAgDfdgZird
IQ9qhrpagg3+k/JWjW8EdgShutEZgxpwoy7/oaeC54A7nlIHo6D4ohVHItJE
dHNgB7/V6DESUFxC/paN5GKpW1b6PG2116ir65qV/Qw5lAbXLx42pB+ys+I2
LWC8YaMx2uvKNA1hGn6d0njE/a3NS6zPZabjALoM0gR9+pvl31xBrzu51eFi
fzAlTr9t0nb2laI2XoZYnIkw72OymEAjGspt9PmUxcIF21+G2ME0tfFhRQDC
C1b/rHDnmIb4joj4VwfSH5OjMidosLPt2lJx9nFJQl1611KfmH1LW+MyPEsP
wR8rtL3T6rohTKiL4+xI7Toq1bHtlwg8a9HIw7ZHJThugR2MrJ+oy/1nRSMT
NUAUXJzip0q7LJHmKbN1wiitHIZmjb/y2HgZKMSvkMdN/2ZukyOHw2K0OCyd
oonrZqFAJDmqXy3SZ/5Wg4LwM7SvPf4akTKau6rihiiBduncW5iMvYML0BYs
mL1lM/9Vz3tcMoze4khKfKwy2TfCSm+6a3KELrVoNuJ0W3IQUhFnMimHuCgP
j10Ozlgh6f+YHzNlJWQANmlBateH0CZ1LJER1o1SgSxs/ngc/wBKyBYH8Omc
T/l8Yx0oUVEofc057PtYzlYsdNuNU5mzIod3T23XOXROu6TbLATyx/fS8azW
iP3GNY4zA9totZbbNpXp9jzqejThE0gQvJZHv0S1FadUnTR+uyHusX9CJZQ+
foyRBpXqCR7ZPM7M7m3j/kdeDVFQu/iTjdErDnzn7F6P1ttzg9b3rasXtk54
Rc/LzaeVqK1wRajqxUy7aGn3Rrq3ImImypMR3lI6PLIexy20lQr82Cw7f3Sz
LkrnY7brXhdQEEc0nHnDlMzTjBquWbispuhnMafBSX9mQb14SsVecLW8AcAu
3vIJawCnrkycBoh5S0JDFNafkwwUupyAtriEsTj5SllzuFZyJy5YQ7PUNNaB
6Vk61AgliUV6HcLqzESLgUMCBLpTbh+C8z4BhgkTUmqUhS0wCd98sJwoLuff
mn6aOkHcE9YRgyIxweTFX0GVoU1WMyT6R9HLn8LDhT0UeYtdbt/le5u174ys
yzLiJ01rMOWOw0cHyA404seKJ8kxwyVV6S1l9OxHxJ7f3DrTn+xpnf2wk+JB
8j5M5BMAuzqxQngOlQJBpsncxL70o7my/D4sR/6IBt6Z1qRnmY3cplnj8UUM
s0G6/E9/E6mKe6WQxmeyYq2a/7XbXqitmGIm0OIgZHUedeKg8vGhch+dUA6D
tKVROXBWGvHWWcZtXokBjxyT12wMwpJTk6qNqr50nHhhev+kKuqfWN7Rn3TA
xReyX7KtEjoYugba9k0xKr8P8bp2Q7dylbeJ2w6ad1w/chcM221CBIU1e5Or
e/IQIB+DOXa2/SUXE7aW2OMiHFXTE0J6iIk+VBlkwfgd3J8nTbwDDTnbONcp
IfXoAEIGL6J44txdifxAt6x82yoGq1uwzUUDIuqyn337aPsHlhISPX0McQ2f
5LHttfMk1myYUDt3Uk4Xz1WRpLomek5uttNhUz2X7rA8jKwfLMPM++17mbne
P9J1XTxuIbAwG1XEYeIYP2p03Fgp0jGczjwek2vL66G/iBmiYQ7pMs/QvKRZ
ECa5D5Qj1+D77D7dbKOh9VnkNy3urw22RhwlKJnfVdnSJNRaTumTDU1v0xam
jzPfedNljh+b+mXanukJavHsSarf+2jmEOCjyI2HcI8bLkHTUl2lUdrjoLAC
+/HotgAXOop8zmYai6r2isFMwsYS0iFWZ38sJ3oSTumIlS8GZAehQnFDW1Ts
n/j4DnC8v15DkSm7T16ZqjjfmVxxXThT4AQj2V0JxTnKvDynxt2HcQbKiDlw
IsW65oEPwZSY/UEQTYf/1BQJHHpp5oBntYIs0F38l2iLyj9KxXPmjV4/ei3n
3+bYZPhiRikL6ScDjbbogALF3RAzzkX7/ZLQo+5gdsQuLg7CorC/6QA75T7M
do2puH3uk9tQW3TkKyvC6mZ68HdPJkpfqWezSTcokAyPiCC1hcLcBwcQJJ0w
xHl2cC1MmqqsfDvvZESScV7JRHkYYqZD2lnevHQgwQhJ55txq04kg2ss08hP
FKQdEVYGhSqEUGIRmQvPFTtuRMZZ7gNxHkQSSmu9OZdbGv8+SzwcSGSRX7Hv
BXrytwj8w1XMbnjZx7izWr1JoR4I54lQo26YntI/AhgICbmbudEpp90EpVUt
LczuLEBw38SlYHM4WQMddLrut+vTbJWJbLfZWIicpba7lHK7TXYypiAS7Fme
NDu9KAt8oD4jZe7XU0kTQRvnBbe2RIVVc4cQ3bJ6SPSllhWQLW9SjtgiJ2Vc
ETxcn4rnnNPwevAbDvglSOFQzgv21o8WeZg8kFp74KdF46T7e6IhRIaNTNsU
gz1mBX+hJ00FRbsDEMVjdjPJXvqllfr4iJ1m7dw1P0UZ8aZ9Ys5sQPOBLsfU
nE+PgwwxLXeUowxT3tdbUDeSylJYdjKv7/OfZz2w+sRITDURgFAXAROIjavi
wzIZu+eio4A/r7JjvyXSI0IP9RUNUj/eO5pAV+V1z8KHOuD7ZUYT26ECn4gO
cSWwb6DVNfDrX2ZI7Gjp2GLsaHX7q4P/X30jAru5DZXYW/9vKPLICl0mkzNi
gGcD16onqF7I+Z6Ov5A8CZ7hwQeQsG43tyqaDjZs6lOU9b0txpDXvj++N7+/
OZjzswPIwBCb9ED/TwJhQ2cday8df6Yc/CZCf+SLR7T3ClE4w4QAYuRzzBMt
yi5kGdbkJ1pO7+OtjWv4lDfTyH7ems5r1xc6AeH3IFe2B6V43UDJ6mc92kbB
1MMVCn9mCRXjSftRpapA+oXwb30sfglJ4FCVbwu+9IcxDIquFzCieFM3AHs4
xJKwhL+ZP4hNPMvHeEDaWcmPyQpDGemcD7ZmORuIo09ZgamU76Z8K4yH35IM
tCebTP/mgZDLF4GxKQeoztzP+F9d5XQuLfsP9y2yw89yKfU/SCr8yy+Yowaf
w7u8Cq8wdgGNVivjD+0JhshYDlIdOoxVDAYYTfdX3Y2JJ7Vzmw0OKVqzkhfa
/6fu+mqbdyAn7SXVdTSlsTL1nlkW4+iNh3iqZou+NziUcyqlJSmXmoZZRF4b
lOKd4lMweDFdRrAzpU2THV8LJh24ZxwlSZU8G4RtK/7fPi/lbc7pqhLzeY8G
8DabHwQkR02V7XRDvlvI5KNDcr05GdEMjlfWQKzPAN9z/oeHqoMB+dX17AIc
nfya88CnRbrNebkThQDs0CM3OzW1ypzjW3QnGskhOFStimJWmVHDs1lzihuj
jlPsf78y4DfZVrAX1jIyLDzQW494bVsbhMumeRFAOyirkFE4vZTC94JetwHV
KOTuvuswrdhfrcBAiTvzR14g6+b3zEqG8KqtqGGirZWjeseGZkWC615OKCFB
9wnoDR88Dr0NCC2EZkhUHq3UcYvlwF0pLsByKKl2kr+xTNqD009/F/8P9Db1
Hs4t8DL+Co/wyRlPr4R2ecQ/5LyLJArWKLNpAl/NunlKgTyG3KgP/7uVy5BP
tDQQGH0tI7BRbvEQBXQRpDf2jCBd7dXNrw0kI9pLiSKrm86szoMSiDf6qm+s
jn7OYXZNc5VQfG4OzLNdKdmoJc+MHsxwSAEWy5GE/6RiqurDVWtJySAys7Oa
sv9JMEFxDnUvjpP+fGJiBvj71cuV6C41uHBdPBs1dCSHay1rOXewOHum6GG2
jNkixaxt3hiOesn1Y3ziqm9LR8g5HSFd68PNRTSQ5PmtWiS8qCpybfJkihEY
6YH3nSzBvUFhWvwSCR2Xlmzi6+WkM2pd2EeTSaAjFJuJ88enQhP/KpLAn3nS
fgKhipTAuLJs13onUGpSAqKpVJ8wZwNmUJonO8AFNG5Cvk77zoPfjKXK3T6W
13tJ2Rt7AYIpgeBfH2WSLIikOknFRIyR2mkOFrx3+jO7yxBV/2TF/Da160yT
BfDSu8EcEz18+gLJD3DDkMPv5hvaMbazM1XjSpZNTlJAbnXikMRiGiYE4eLD
sTJ9QYuSzFRtI3/AvXB0yqkqX+2ZyTMCCrHXBi5PZKVG4kiet8yaOSgGYqT8
GJP8f0o+zUEJ/D5oKtyt/h39PSP56TTWKbw79BWqUyg+uH6z72muWa7b1for
4j0Ash9Mj/Q0m7IMTEerfjC2mAo78nK78ZUF/pmQgcuwligmNwlwmLhMCO/q
hd2OMNHlgOzNPPsqVwdhNBho9lK4KPU1nwSdSn3wPM0EashhyYDicZJ9Js3v
p+H0Zj3/A0+b1Dhx6RXowCDBUg1UhxrZmEzal4OS96pUtHVyliyyfKyoHyYm
GlbC6VvbisxWJJSM9gA3W6amg3KX9njQ7+BdUXUNe3sVrEhzPImVsA+wwAoN
rWG6PhYv97cZQrr1mS2IovaUIt5X5eRsGMndwkVR4ZHvqgOYFW18gUcinVxr
fGVwPY669Yi7WY6EGrxKJw4BG/N0Xu7wNci3b+ZM6hN/QfaFMaRnBkF76dZK
JX3vB6vDXlL8uQhmlWtTPACEJTRNhe4o0PpoN0DkNECFdr//d7I33MUJ4u+c
ANlZUBgb5sCRexhwTr+HfMxyPo4pxulZsunVBmN0OE59oEhSJv7XU6DbRYpK
J1gKuwPvyT5kJltt4CdtfkQXyEeLM5GxRfNfVGe4uqOHBNa4wu9kXftATpTE
4p7qG/OmDDbMheP3rFKZCmYw8MJoiMAoKaHo3zDnJgUJ5JK0D6FJzrqv7jpD
wIYS+HIHXFDmhtBT8ZHLaY0jX4stWSyBTc6HQ/w0o/YheReCQ4NmRHIB8SPO
CYG7fAHbtqk0NMQhBYNYAQoyma2wpaSaq7DRJXL690bCjtzACD8jZhh7PQMt
y2mwu5OMYjxUXfaO2Q8s1lChjejWA8vb5XFYZnY5NPWmdco3dy6LJ56PDWhp
BlmlqCbqt3uff9CkbekvQyQgrepiAUvL1kYFFc2fhUaidjrO8rWGCBaQ5Liw
ZB5vVtdotyVEB62I5/ucRrShvzVmeTrmKahgnCXEgDqYRBBxW3FFLBnby8f2
0K4nIaPPMOuBZDqH3FEwr9vk7kHkM4RZCd3OsapJepyOeap/JKfBtxoxqe52
5hPLgAr/k4/jO4A7+JUsxVy19EDDC0d+y04E/gyrIdFhfrg0nfWCxcpv0p2W
veXkZmKkzipZvAi5T7k3UoJ29Y1bbr13CyfAhuNjA6HASpMevDskkZMNXpCR
+4UPF8XV19ED3nxXqteGSFX3MUhF319ngg0whJidA6/JiLOWDL0U86ilbC31
Y/M4rONXfxTv2qwK7p0lrOIgeWUUrI9s0LLryJTbKdE/fDe+nQjfwXfVrz2H
DR8xtdDF81HqNXqS9xogTYNrMmAdqiveIEK5PsU5DCQ+4jtJvB3x09QyYTiY
Lo+uGSDFFmT2NBcdF8akW083+VuFmbssbxsTsdp1nnpnyRVoZGGSpWtGgZU8
jfDtUxvr2+I+i5qoiLQ/pxAx/fxvbEsJ5Vc0m+em1J2HwPH8+COWLmP74Ecb
X8gjO7PqPGO2J9WzlJmROiDJr9DePVF7XDuJFVwmXdZ+UqRBO1D6BBILlcwW
ckLSNitLYwg+1CUh3br+cr15dXFcxCzPAdtCH8+xG2ZjlnJDQ3obetS1aB2a
V+gjK43PCy+dWY+yMUxq051B5H+rJe1X2X3dgBwvvL8Wt3RdkJalge1mkZP0
nNyc0RwuTO9hIHoCOYhOg9Ye+W9XBcyUHldcTqEUTeEGtqjL2BwmLeZEOOXM
cSjbE46KE3XFzQHrOBajt8x9aBZgcXb88qDEoDNLbcZvfwbhxl12ax5iMfWX
cTjF9vmUYtatvReC5Zekbw5DYKinE672rmJzx9ejXYb3XDFSzRE4G8Y35gNO
6vp7GFoTFrDndSEknbVu9YfWxbbJMz8awnv5/oo2DBwTvZdiZLsr1SGaGsBz
KXMpTFE4brC/EmfsOZQlxU/erDbV006qYEq+41wM4oaU3aLbqh6LAFgPegXA
oCGQ9WwwrPg440h73d1nKBd09IJUk+kTzzS1H50B5H4OPRgm6CJ9QwHxbMXe
hhp6CteNjDGAnD3ReD9ZKhs5rAeOE10uMwGUkLqo13ruTiWG6VoegKwSyRbb
kNcumgA5Qmv7OoVZ/YlMERnYhpIshA4G4G0S9G2HJyThA1RG3FNzsyh7DuBp
OHXXPR0BUZ7ZPB+pUAvC3RmHQAJR/L/0GQsN8PWzWF2HoM1DBvucvm79WOV4
AUky2GROWowO/fZYTGHRwOxA2pC40yHNE7OS0AWzxp1E3EtV4nRT4iDUxzkg
ShmaZXNKiv7dQnBjgQ3As6Dc1zJoTtfSLkxWxnnl7H33pCu6DFuj0eNZyvMJ
nQR0sqr3ayZwJXsOUeGTxKTMXEKaxRmQleHJ2YodDMRJrBicv5PuJs7b5deX
ytZtFRVfTQnIuTCMLPW8Mk1lOHMtM8gm5Bujgp5KsLTVxHtrVZfSHLslsEDj
TQ432BMGXrbCJGdIAgki8MZ5o5eCI5IPbYjtAhRh6Ry6pg+BVYtszneEWpuy
jHOwGS8UTB/UHjW7FiUnJfEsY6DRYxu4DZ5bIYykHmhH8ZeQTCEmssM8LRHC
w3qmwCRaORNdVnPIT86GYISOIsW8FFkW3juzID/DstZJAm5sh1y9oYCso5Bm
IsRLGsrYCsPISsuciT87ZHXXTsMx+k7oSJbUOliwfA82UcuGuWnzGsGWLulZ
hvIg5ZlJVu329UDd4BJrc8+8xPOhPfE5xlINZrgI4LMnhjqbsR9GI7TkcKeG
uuEfUhMQ0lTXu5MYDOEr/iGoppk3bzTmM/ove04COdAq4cTu3/BTuvTTM9jO
0sxG+s5D8NftxIBmhQybTYKj9iSTkkmlf9e8Ne3Pmb4UTP/OpflDjccsEHKA
OJSl7aqtyJzh5HpODbADYjwXBQ1kkL+cmJ9xbdHQ/OR6JXQ5HyCKbB0ozsIq
DDM3FbIWMts4if/C1T57W58+s9OUJ0Phu1NlzLhfvWo0dQP3dwHxiA5HX5qn
1GQIczHnuSw4FHe5bMwE7u6p62TRz+VjcqF5R28obnUbOecNmrMSNq9Dm3iN
c/L4ymri9EM1cO8B1er8MXBd+N59V49vcwXFlzwbDOMm7GnpAmaqampZk8iN
VGwS81AxIA4LaiUp+ZjqXAmJAYH0CtwU6UPjU+KN3cmlfaRM7jttx2jx5C+h
Aez9KOWV/0RCAU30erVM28VmUSegmwP08xqxKTfFKplBJ2kKiHay0ZWxqrlB
xOSIomadQfcyudwEPDEv/jSRgfiG9qf5SXsI2ZkvD3g+/neX3aEqQ+izIxyU
TsaTdWtyRsjKKwwuT6rNxo7G+nb3s4GAF68Y0UQuwB9gPa1OVRyCkVHpulEd
chHISj+9H7J5NKShBThFULzEqC5u5oBVKHy8mW6wYD8dx1bVEu2QGJqyUlTq
lediAV/Vi2Mvi6kiJSQfggj7cYDfV6bcpm9m5l8g7+ph/5UbGGR10GHZ8PP1
/PSaeCUTDJwqA6cbVv1+pJaptpkfV3B8P42AorfN1wXuyfP0VUxNyczi1A3r
may1usUVOCQqfAqtY38s4UiaI6Di5JRbW0MGyjSz4WlWhHzVhg/+5bzg5yaD
obHUrdE+13DlQqgxLLHOQZZ2XUY+mnXoYc1/kRRhnar09lClAaBBx1n6+zAv
gR89MW3GdZ6seONNaVvYPQhzrYF1EYjQy8LsmkdjTAsXj5CwUwPWQi8T2jnj
JzjdRFkBnjITfPe0uKwLR2YsqEqhDSWUIc49rPYfIGPIvIhfpIOwKJhnp2M8
heu9U0qQQ8s0SIk1e/NOYdgx999oz06V27CwcZJW+43koDPDxozGFaHd5flf
NE49aX2pFAzNh0xWYgMV2+5Q2d5Fj2cNrFphvHzaSl/Cn0R4K6FoA/mxfJZe
Fjv3FpJGHO2rtdrufx5cAX6Vp4XO1d6FXtdsiRQMX2vo0EPFZ13pyM7ZC8Bu
k4ybZ4ga/ghLsc26hAkJWRaZdTY4kZf6O/yNxW68kULnv9lV/3Flzan3A7GA
MrY053/XOhG3Pp67UWqJa/v9TOtX6gx1tApObl0S/0gS0xBfw+4S8U3htEhI
dgvAnLB1INqi2PmURJiOvqvxHjK1TYRBwzsKaI9wxWN+U4IAzYVbAqdcZZDT
kUauTvt44bTALpkEhL/0XYHjPhJzKkBwHssDsNP0m2wokNgUdwZOEoLHZOwr
yp8MdowPHiL5XW/KiqG4cSksiAoBEp7hO8RTsKfdbK5k7Cn7NsFLh7lLL5Hp
0/gAYz+6JOa/FcoVTy6hfSaYTr5KOj+/5BuaHe9HnlNdZiVMF4YY7eCAvHD6
udnznZ6ohzZwQFpMnZLkMLYXyAllVrHb9O0+PpWErgvsID6IIHQ0nTwrRJnC
LutJGcxx8K8NlJgoY55m2gdiKfnUS2PT1ViRnVzlooccRptg6tI66Kyyyoyu
WbYGWdyR/2E44I2isKJ2gmyjLTO/HrjTC5g+pVLsR62CTnXg96tW+/Sq7brr
L5WLCkwIKjkCqK7oNvfNgPkyQg3REpygFjMtrC0xj7Lyfiy8vkpy6okwUIyP
ZobYvjXO7Zxm6iTwgJev11Iq66YZimWhpULj/PqQu+Q1fmi1Wz14mfnSyLmO
nAqE6IlD4L29B0BqRe/cde6He6qF70Eczw6VFnlkzDqur4vJssUEPtJiaoQZ
8S+kZFJI/gWiJ+9Qse9vS09SmWx1nwGpvSNIvGocpYew3pIIIfg8u9wxJ8wr
OIWy3T/qsFCT439nkW5vzVYRW+mEuw7XY07njc9r95AjXj65Ha1LbVeWkGMn
K2g8CDRIomx5lCTbLs99FhU7oqFU+ex0b0xSgZeEUG/Eu15RpNxw0HrntkCu
1x+y+MM+lGofuFKiW1XCseyORDRjCZIn1bOFUe/R5T4pG+fywFd5x0NmCJL0
Pps1cBF2Sd3Mz7hgHMUIRhpqVQhoqjuVI4G7EtsxqmpmH1ZfFT8w73ClMZru
RulaFsDHUFfUwfPX1L88Kn0mD7BzPRdRme1MBlMIxuFqxFu1JDeC5QpkdQyD
yOEDXmGvNbQ3LvBrQmJkDgL0SjcrY3oNPhCVupxqA1bNTHaxcKLEtMAa1ysw
9r7GkUP5Qhc6oglFlgPWlj9Xa6PLafUQkg55VVslVpWSNr5hQEDB7dJnWnpH
RgR87FdAVAGQHpHFK5V0/14VdYVamlwabOhlZEAjG0f3Av6guUhZQXNn/nNT
pxmXSaRDyoUhGYW6/MAttgG1J3XMWNwiqagEJewYwny81oWy9ZugZy1pZQpo
eWaaDDjHettk6bCP/YkET1OSy3gKtrqtePpeWZUBO0jeLxCaJqpy6ry8OGu+
Vnt0Sx1PShty2tg1sZfYJyTLmDw8gQLnOlYEmK/1D8XIv2QF/3l4evpqmuFE
P7KgKQq/mBhM1Addx+a0fFF/a3weF7Xge5SuT44S+ys7u4jCMgknwkrf41bA
UiEPrrRFU8SuxBOxvRibk4Vai97IToUmURzr/MrWW42qNzeG2xMd4YQT+Y82
Shu25icze01qHoAuCp5uf8PLsCOB5DxC2JibE07PgyW6dwizfDLGPkVkDgIL
Fu/JNbVPFGdD3dVgO0gqc6QOhj2FqJFRvEby0CyVeHgPJxxibCxOOFQqTLQF
Y271eRIYyImbfEODObzqfWA1MubjvOPcC32mep2eJuVpRidfwI2guDHKXX7r
sluApzcQMChVa6G7U0Uo4pdC/4HMWe1Ab0t1jyFTWPjLYif9NahqALu96XHR
evkz2+jEZcGPTqQGz/aZ8tXq4QSp85aVp8kOkbjcZlJgakplnJHbUKXqa4//
QvJY+ykCB7bDyizAgzs/2dVgbB/QRkhLxB1LSaJu9RjJSQwfsCka4ie6otu5
K2cZrAeV9aUNDN/85nN08Bt5Q2OEKcvC2zegDYK/IjGkCBqaYCDMDp8JKiwX
HRrcCnZnUodR3xJ3ddj6vBJ3UGPDCedxHNtMXZdYWF6E1IHU1cLvIw7shLdi
U5tAJo9PV/TrjirX3T4DC1moPexB5LsRsVFIoFlKPTjG3+hMQmUOIvJZPoIO
DhL8kyZRbxOTefswYp6gqAd3CenutPShfnS9xs4DrHdr807BdayeAzO8p2Sw
jUerjJSr+QuW7T7RpmtacIyjpoKWw01YFv2RySjFLC8BkQd8W+Mqc+iDfXLH
xHy92/dcqgchm1jTCTbAUN4ewmp4xeekPYkBM2QiJskaI5GV7O7ct2PxjMY3
YqCl0FXu8NNx3NRlbfANMGHc6irF5dEPy6UmnJ3++fnvsM29sWD78Ls19QUf
2s5CnKhoNIGqVj4WPUhASbLhiER32N94jlDXX+VaG0uzcFFIvKbm/X0SvwET
vV8+JvXAIFzcpahJIVmDUzMc2wIyn0gLE7UrMi0p4GykmH8Oso1NV8G+B6Fr
hggUzrwJhVpRIN6o3DWQILVgkq5qjp2Gy+i2gQ07qqjGS0dgS9NMRS7CbyOO
F3wzctS8KhfZ2JqGzug4rLd94SQGH7eLr9awWRUfbN4m8UN4/N6AGMA/Zi3i
3eJIslvjE9ERZ2uQSq0kM9iOqN0JOfn/0bRrBWXsH3mOYtzr0L0nMdtkbjMv
RBQzJOCSmRIW+RuCRC/duuRsDUJ8NtdrAa5J7YwwEzuqgzYiTXgwzFtTXLsW
AKwCL2iPEtWF1si5JbSxnB4oeIJFxQbT0QYwprLSAbQlRw6YiubhEuTY8r+T
kJPtbEups7CcsvkKLTZi04r3F8efH0ZfYWezFYKoAwzrGJIgkzWquO/8moJ7
yO7WQishDuRF6KDT6pWOky49rm4r0iaHlFezILg2ytUcpuUch0UG2pujJMP+
tczuYkF5+mVYOASeWCSDpUs9vWNoOBZ0UurGX7jtqwGeDo5ht7SdBctegLja
f3UYrcDzIpBbFjkmmgmBhS931Kxe9fLo60z8OLiQZXfu8rh/jSwIFdY07DJF
xwZIEmRmJQPicEiN3Y/HEUq80tHsb1rT54EhKN/4oW4pAKQscqNxMDsxf0oC
JTPvuTS2lt3uYchKNZbbFuuE0prj5wcqi2sxjznkCMnbzQxnBKk2odwK+89s
2rLWxzG7bcg9fT4W0z6AVEvefnM0vkXXIJQIvAe7lKiTYh3/Xwfaj68KyTpy
9Q28rwumaGw7lVyqQRqyJ/coWUD2A7IHbiUntaxozP5lMYNiLY4ScbjlYr9i
AWijAzUKoqM0dxsI1i4UwtksAZ/51MH5zWyDKIF4NmqvolqZYzaqHP2k975y
pJeOoO0ZxTjdXkQYdUnJkemgqu6ZD4ry5FfHx+GgatDKRrJYHyIvrSup1m0v
lgDYUmZcDt5Q+dwXTnHR6Cv194VFl66e45vq0hqFZJAQzq+M0h1SHWsuVL9E
beIRohcjFR22ByG/k1dA78ztXXXh07S5W2loKxm4KZXRD4NCtQy1AFN/yXOD
0nQPxRSXpbszhe32TLldWxHspnFotpbnPe0ZQvH8ddjcDIcXMmKx0BuV8ISU
vNaSjC4G4VlP062MPhZaZBwphPFL6bA/7H8hDd1XuJPjYHlEqUx7VdHoZH+i
eOJ7nt7BYTfCYX9WKdBMylNb/M1ogiib9rMsXkhZSuns951MH+S3hFXZiMyX
+nmVjLp0mBZO7Wj9W3FSSMJnSCMWiLIjeHd2vVwhdBX8+MzfDge+3GMl2MLp
ixiG6v7WzKxN0ILBeUKHo2CCvA82lNx84IaEaEiQztPkt+jxxpKMrKk+CrCU
CHC60krxlfmhzOtjc4k6DkJgHJXEtW23fNbk5gOYiR4lwhAvlK/hsjB+8aru
gh90o0UKHXx5oA6zTi4INVuRKYhzGegUFUT7o2RCQyZsSx8QYalcfV40tQMG
VOFilB0OUVpRTembtdrqMbiUDnR0aAznKNQhmuxzsbNsw8Ol6D2RRpAdMktZ
u3UFgkjfR9Tu4o0MBDkFXF/dyFZbO/5uNNyBslgbxJzP/S5NL0+Fc6rNLSgN
AeYeFopVT5KcbFetwVvVUnboLjwirVHwlMYdJm4EHX4RrFdMZmNa18y7zzJS
vul9i3l0bVeeM/MPHVOLo9oxLZ7WAosHWmf/En+oCfNA87uQNn0vJMJEVNS1
4qLOtn8LYAzrV845WLnnJRdq+8LYhtPMaqss9V2dtsdpM8h7E8pfM4qOyAWJ
3/29x4B/B0MeQufK+CKb66giCc3fnt65s+lhFuRYwcgFcuxooPYR9tkLgwJw
HfWIzz7o721lxwvmPmuF8mGy3HY8NaxOZwlEilvpaJROWs3WZNpUuTKZbFU1
z81MePscaW7sDYOD/Oql1Ha1l2NxeClentaoBaEhpk9j2UWOsXP5KMyCmzuH
iWKBop7p5p7KEDe/mWkWdGUxyZQn2RaYeatbYpdOEw4f4IdHGK8rsnms0VvQ
Xv6ozi8WDwKrbuG8Rjl/YDPE6U9A9m4KclGtz377xz+1HcxrC4f79DddC8q5
rNi4VAkmMX6xjNiFBZ8SU7k2AU9TS0IRCGCaYciqQ+08YA5YsedGrohPJQua
uglvhEhYo++bMsLLR2VunONs8nA47JvGsc2IoX+uUN82Wijq3ww5iWVQTagW
iR0budkfW6InNcQnqAo5iJHln1kQrxazBQYGNXHn+rOhbPdZb7nucKat5FY5
oDlUyGOwYoBS43ChWG3M5Qhkqg0NObaH+Fd8W6FyTtZOYu96pix2rtIXcqFf
oJejFt9l28EiWRVWEb/6gAaJBeLGZWuzvy4D7F+MzdHTEs6zsyNz3yar/66y
Jsq3rvtQPKSInFJy4m1nbM4BwPoKf62ecF0487I/KwP1AUuWHK4w5rBoRJO4
2u/kqWwt13nGldItos0rU/wRx60h7KniidJKzUbh56wlt4WC1PnYo0UelhkS
ZDoqdxteo9UHFaOEK3O1k11XoqXRMf2pGTBGnAv3bLLg0fNB0U3IBlzyVM85
kw3EcwaehYolq0EOygvjZlfr3HgHdfvS+17Eqy7GeZqjmWnT21Xic7rdukrT
w6d9Rz1WT+AfzLjwCLoY/HqbAV5aGDlbB0zPEnCCvDr3mpfU5j4dtz6UAepN
R8lgrMl2StdYXqEmyti3CEnw0qwUSaQkWoJmuV2E6bmcBmB6L9jP6X/Ppwrb
aKDs1Pur7becqB6Jpg4+U3uM00nbKp9T2qp9dZPpIZVZwDVw7iZrX13KWuJx
P1WNl2hFMUJhDOsmLVdDM3THfQRXYwK9Asa9wPacBlYS1YiAIhciz35XcM24
wHDUfxm3hsQfCdc3T06SvzqADvUMPxROrJlw44Q6HSi9xE0SMHzOgKC6xkU9
oMveCBowa2K0rFbqpHubCyYWP58LJDEDbpKMrjgj2FTStFGjj1e6d9vR6X9L
1DTqg9XjyXp3q0VclmcaH45INW1Db6gBiROyt0I9FKFHqXrbtJhEAe8IqDOk
UQ6BiXh+3CFbg92Q7QTVoo/hyloEupVfgyZA0yfWkDL/9mQ/yIxdAsRDAEqU
dSCYBpAaFaDlpdIXM3UE/E9j0PHimjMqUqd7LlB1aA+uA8sU9QwcYT6a8eNN
ojumtqwGWRe5IlWHmktOpFeZHGIXQsCWer4fXui6UoYWEdWFNitAUiC2WQQO
/9GKyMAbkDeQy7fpOxDoD7T2LWxsCQ/D6ZyuAY7FviF1bGsAaSmubMdzqdbD
Rxi54cez1J6YzIz3DWSF16+ehsyOEqe0g6OC1swhb9TAFhboAEw3rkzSseLI
9ScM3Mkok3qf+vf9lRzuqjmvOsQalDjYnzJCAjqtA44+fn9JbckrjEgfwPqw
IkpdsUtyTJgvOnD5Lm8Zo/mrdjXLvTflJv8hho+VEYg9ynk9IJ8vyKOKtY7x
AIbncmdVQs5245hQe3bbEVd1j/wy/s7A81P3zozuovTjmxBTP+z7j9csEluJ
dQEKszSOVHjrAia6CvuzgnmVZbDWxBV5z6/pSgDQfZ53mcWeqwe8AWoNyxth
hFYE22IvvQLEwGd4GZ29eXV6zxiFVwSRCclvuaOM+Ra9K3qq13mMaY10IFKz
N9X1Z4BQWDnDYmryaTWRTA+3JGh+ymAV0LBJ+oO5FHrhq8enHr2ChzY/fzl7
iMKnncips3aS6sk56ydntSQ0VQkwhX8bTMdzr+dGNRFegV+qx+1oriG7qdSL
IjdR1EM1FqsJ9dqPfOv6eaXZAe4oOKnh725px9yp2ffrby1tD2z6TIqatfBT
ba3bkrzp4HHrrjs8pP08jEYDRqfwPJpSrW+V7Qb1Y8Uhkwz3lExywR/H0XTD
VKGoQuUj3MH+AoK5zh6FG1WI/xz+BQgNBEuvHlZGiS7kakXqrsFhMdEs/wWO
tbGc8WnIhdAinahY/htpHaO7j+EBZCFZiRjfeohxxTItxb9V0KBjkNFYLzF6
BwDT62M1t3TAUyENAxcaJC+L/VmAWjb7kIJBcKA0ofW0EOWBPvvk2PINsW1n
lH5xcBj7XMWMfukqhaD/o0e9AiwDETUd/N7xzuDSzHG2uOLeUFInHTPKYHCL
V/40E64wA7U9yR8O8TdVDt3FEx/uoKVQjGZjCMTXXHR2A/FfTFNgUDOsWNM3
QsM7suJeKnWjnzsSxOMF8v/dguwTBhi2ZnMHxho6mrU585kNiuWjDxxuj60d
/bRPUWAfKSkSv+POAa2ksu8TUOJ32yRc5EWaaHbAKXpZM3Amt1mWf/VhjuO5
6v+ZnOarq6mR8XDlqJ46dcwAMg+qvew94zJSOewoUzDR1hOm243G7eqdfs+z
aObNoQH4cwXjDcRJqqP+tnjT5DsmOd2f9zMKrbthDc2WNpkwgp29RGy6/sH3
M4SSUoRYou8TXhH0Kd7A8jtQzuiTV3hzLCQZ0k1rg4o2jxYU3CJ7BcsRWnmN
GivIarW445sUEgKyv4EeIU62jOnDnpZPsOzhlHYs+cIzoNYKPoYAz9oV45+A
15HfAcQ2W64gamcRn8GukVkfCvJI8FRYOJW3q3tPZvRdWMHUXI4+vGrh9fkX
0h/S7nM2tDh32707qIZsDmxn3+7nboHT187iVFvKJ5MjSTzUKMp2LzWpxTmo
vo63cpVhdfnLIREznSmwy1hvtOPY7G0GF5EY4vK4jP+F2dT8pqGdbcDSWRXR
JvNFrPF7H/nbG4CUrM8zsJYUxMJj09GKcIiyMBXbXXIobYjXfGYumesR2eZs
ZU1hCYcv7+KMHR7xUhDsgde3y/1dIQswdWFnJGTnbKBFLbMroVQCHZ6aM9Jt
Y1zRZ0y6uzlpdmVZeNCFl0azCIpxcjzBdzphM090oF4kL8uSsiGGzkq8GpgA
hos9ALkI1W15Fc2JnNJleq34dLGi6feE4BEa3cyF6fqoybASOqQT3RAVhO8n
azfXcZG5zW4cU5B64vKb80I1/rpcDpmjqd+qj3Xm7jJXRkjvro1aVe6rOO5h
OOey/7K4tFd1duVAfK3kog60EZQyYjS9o7qiHygDkObImrRGW2+O+3B+uhP8
aHz4IFVWRbxRh1nLNedAVXeqYAE1gKzIQIQDCecJIvVUzoPb/2aUht9R0coi
DRynj1p3K63O32e/JsxGzmI7BTK0kDYWWO0H4RUAutGVp1Remo4Gtwc10I+t
aDj6tbXcc3+UOBTcWSxre2yqLI0GicjIHWkmdxHGWZTuVMTwrz10e0fPn7rW
IrHbKsd8Z37CmH6WGFbtrgvYpyLtADsO789e0COeU6tsBvO1moMzOILNDGqp
347tnIP+2Q9eS9AL5SlpG8InJ3F4Qw0mmZkLgB692mwEY7PbRHSUAlcmbCtG
miIaWx196BleoOxnmlEteSbST+N8/4PbGg/5JJqwvWQIaobpKXIv7/j2ON5I
DjneoAbMAuxULu9+RlAwQczH7j4xWSk98b33g2qN1bOBHC4taFHdndJuPg+7
OMZFHa5cOWz34uU7dEmUVPWyIZbTe9z4IQ+LbbbLFUASOp187CTqP3ncr62o
uxfFd6xvRwR7yECEbyj3cvAso9idn1yz8u1gyttUbOnrYGe5BUGKZNShe5xn
Sx1oLRL+gLaFcNqEWYFkKuzm32hNRfotSg8HRV4p9s/ZFQKx4MSS2cPGzFqE
aM5wdoXjpN0yGpEftp+hqR9GiSjmIoUgARUes4SoXSs+47NnKOAzz0c8EDNI
CoyNpV0dFi4d1tEPbbeUn+MCQC7LOr3Ll9UQ2Yl9Cl4dDInTyQPLDOx+lCgU
GycIOQcAWiirytZuRa9eq3pEJ2Is49vcCLE8fiq2qH6v0bNS7GXxK3fpQMWn
HJxVml38UCItkq/8jdWKF53EMHvlPAfcQLWuY0jMPmtMxv2j45NemGESmQLo
lBHczfEMOEfJ1/TTn4u4GCZzYd96nxGFFatnP2VqalakvLiQLqvN4IZcBMOc
NklWwNAQc5RlwYyrRlEDrzzLNVr1Z9jqci3mC6UA1BG8b9VEJfRY4VL5UyMh
qc1tucA83QXLj5xeo+4gzsK6LpLF0mKDCa13ev3KT5eDgFg7WD58wCzhFEYw
IM3Xr6QB0yE3FzScwYsltBMqx4siqMd/CAn3dtsB614GeJWh9ZNeUDC2/cEL
uVb7MJuoe69Ymu2I2UkvjAksWoQmchJg67PRu0jOmWn1FofZiBNgPmSWd87T
NcrT7fBZbtbfmgA9a0on8NYY9gHtCYZxIW2XnJuCyn9S23hOmm1w5EvT5ma9
EgXjExYCS+PZm985+4MTUDFQYZvOrLcetD0/JfN1F8QVvwDKljx53DWCLvQE
kXlMqSo3q82Hga39bRBt4vxDfl8rZlK+lRZ4506Zi+iQnz1HU29N/H1bmZgq
+mLkp23cuyfUYziX9tK3Xq8BO0YegUh9fGXapxiz0dj7/SKoN/CPKlEk/PqA
IDi7Fmj56+0+K7f2v2YLElt55Y6yn+DBpEFYLsJYvYf54tam5OvVtXHfXqWl
vnvY/H5Xq+pxeE9BreQ5lUG+IHxfd/s2ErUoVtEe3yFnGoy2RGhxvccZzFS8
qzIz9H6aAhBvfF4LtbM2xg/CnxB09NvZrA14+W1ENc3VMIA+t5XmqUNiQtMd
wZgZKmF2s5y7cnJ1WX1kuSu9mYK3bcIMs521x1TuWYcRDup25roCnC/MgdcN
VS3kQ84nQhDX8g2hnHRAPousM3vy6GKEUrvOTBSCqTBJUiyWdChYMQO7K96L
MAarGW3FOor/yqSXwT9so34C2dCnM33RnPnmHhKys+NXbPmGkVF45AH8Ye1w
jE84ZSs9C4E+spN+6ZobTqDW6ub72NanHFqI9oy2zJCLwI0oltZvpbHUBQIn
d3bjQTUMR7ScIvk73cFA4ZDnH+GlbmJMoujJ5rpKozzVlRSlsh80lyL72AZc
X7qI08oYaNGtJz9VGrCtAEipkZDuWYvEN1pDNfToWwJQA+aE5cMPveDzSKHX
WH9RHUjgpyQzt2Qdql/fZMX2ktfMPWaZ/t6Za3Wc2IWXPuDv+vdrkgmmsV1E
6L+BDNXIIP98rmxzClmhbgvwEW70kJnjoR3ce7N4/vtio8EBjR1BZJsoyqKx
DEJ/2YM/bXqCU2b502B6D7Iu7stin3+EvUrvMmE/PU+Mp9ZpNfBGjFvr7oGq
puLyLH/mDaMMqFZib0O39NdIsOWnSHkWLB5P5BYi/OCbnzSJJN2AkabxyRG9
ai9J7lf2ED2KXD7nxm0O/lXb9Xs5RZGrBQoRaH3nJpEZiNMkftl8ZrcyBUcn
jWaID7tKPrsFOZoGlT+ZiERwm4k3/z3ZbhIxrTIWvX/PFcQnNKODFZD1rRhJ
Ku3uI81YhY1i0zZ3hR6T7Ln4lWYiG3ZOzNYueW6LoWt/woHCxiVXukUsHcOX
fzKoqnM21FqavQDPkjqFmvKjfMewMfp2qTx3bkGIJdACHDtRKNBBuhVU6j/5
bygS/pumparPQsUY3csS50IshXTkEhhU6CAChFMlRuunOFQGqoYt5SAaVRjB
Li+lOZPTBs014/wCkpAy2qGHnBd/qH2QjRHcZZywQySNBDO76nvHfCjQsLDQ
0koA6G9wIP3JQ2LPXSEGiNQOh+2a/Q4ekpt6rQpjn1eYZeCU43TQroZNXrS+
BjUBdPmyMKOXahgpvXh5u85ObitNliQlyQH2oGnammgYxvYZEb/D5L1TGCKu
vrtrvZv38TUjWsHsCK+WdBK4GYWFn3AWQsamox+zqnoMstZiffAX3egFDyfd
v9fv6KByizQ75LBfHFAHLquOdcIQJOytUiEb89eBdie/4LfzqBZBOvktpiB4
wdxanyd/OTYI+15ykyfFM35Dx7Vm5QKmYnWV2dIRTx3afwMCDnB9zrU+U3A0
cBso1oUrTifKjExY+E6FFtLaLzknOCNLZJ37kKqiSZAh0KqDtj+mbkWIQcmU
rUge7M7SMAQQOJTH4AwfQuGHUHP6nH/2gZz8B9hK9XX0eMAXYHw6Elyf9kAr
1aFgn3GneIuWz+W9W+PSbbri2mB5eZOwG9zktkQoG1mONkDjXK8t9Xido5V5
OwCpTadBe+5EgWX1fzget24W4X39cNwf8+xivgltJOdxpTbA5xrqKD5W1DkG
SUvwqhW1oKP2GywRKBGCIAb9q2QtHgM5DuEawHY7n3eds1lpkC10av2lRZBA
8V/p6yGdkY1WIloij8P4UVPw1SovcjxzF6MyaqlKH0qWauu35h5P+bh9+U9Z
PT82YlxtNe3SIK02t9j5+o4rQCWpZSyVB8eGB9lkk+spR6tExBNzaXr78nXZ
+2hGGTuGdwnmQ0SphxiBFJu9Oum9H6YNYXskScc9r7fu6HjWAh1B2yrCVw86
Hq9DnYFzKmM1Gzh71S5ztY6VnmumRdNbxKJ0EQ7t1WlAg09vY/8NCBBUGEic
Jiz9K+jfLsMLlpF/h/VzB++ez4uo1wLWPCqdAJ/2DQVyGzYdO0stO14ZXuR5
MDO2Ev1th+7Evs3RhKXswwOp1cJcD6hDotp95B1r05BDVnlF9XySvmmLADOr
tOAjR5uRgHdoeS56h6L1ttnDPk13t3rBRi9EaMIcJ9iDLdRQ5QezLrIk8rb6
i/AuLgHO4b8rJ0Z7zU2OWSAxKoXJlRwPKKUZWPD4KZ3blcRYmfsMqEvhXrJk
CEQAWgTep2VDtzq1lX6jwn6oXfROEvf4O20NzlQIR+/v75K1XdVtD0o63S6c
X53qQlptfoimtgkpkPF8bdKBF1p79pIic8E7FeKCLj66kcxljs6a8UUv1lCK
tIS2NVukfORUiSjz4zNJMudck6lZkrlFMSkkbK78esKyh1sjKbluZWtXpvRM
sY0Bkkiy42dtvNJrM3I+kWLzijhU8/ZsKBFpxQap6/SdnlITL52dRWUE2HUd
zCXz97xR8O6JKfICG7+V8ShzzGi+cTeHkUzauREBXshCxBqmLyE6HIFPaPE5
q0IZDFfvxgwFeJcVfFlWx92XiwmzMTsy0RNxPYz1nmVbu/QiG25IW5MsL+kK
+XDEC6WBfiPevt1omU4WCJTRRGeNhNI5hdiAY87uycryw383oc20WVezT2LR
vYEReg8hyxIh6unVQArwk03j33pstuleH053DEzEKKqzv6jHGZHRBgB8R36h
wc+FZF4GxPPdmdqLbSxAW0/WYFI391Xui8OgOQTtAVH9n842Ljm5g6VF60eU
8XNmmNzB7gTE3IahDOZYz/xCdJU4xjY4lwaqJsZW4i+GreSv5iQr2bZ/HLuX
PiMG/B4KWPEYdf0+PEQeg1ucFq0ZZ/o099lNO3+I06jLtqWYW9rZOVp2UaRQ
AC+xedWT+bwD7LbUpSCtISzTaPmfUtjjts4lsc6ts0EJH11pP/k+i4WENpdR
8siSC4Qs44yruosogR/iexqma4btnhcXb4d20sKjiSq5/cU86zspuaWgGOey
lrENU3zGfYCsM2g2W8FuAgI0qZGymButA7Ew3hffvro3xBXiQW+sPhNMtOSj
HjYpiLQ4tnRFi41fKxJmazFMjRqwiui8BJ1xuWn7zNAjsPHkY7npYj2y3KOY
Nz3g/YZIE1UPw6WrPxvnxE9tNoxaUZgkyhnYdyBJF4Uokq1HUPYJJedmG+xb
0SZEYP6B/v1rQA8dN/E5WYQQV+DMzp73rg5qHoyY9qUyUaFPBUPXiQ01Rc1I
gw4CF3jcPdPotvpLG7kP8AT1QeDVJakI/tNUA8BO9hZVlCdBWeLGMCVsfdPK
1NOK455raTDnbB84tisQnG+BoPgeYM8oe7HsshRKCJ71d1F6XvVDdraiIStV
iLLFNehGhaBXdfQ39PCDtV6GFsWyq3brWcYbrJTwU4OQNsVU0pOKCcIkmyjD
Atpj/dYd1kKVMO11g8ty+YMRY2XZCX3sXrG+t4Uu5gjXGhYU2Rh2BCJCFpMV
x/6HquIRYBkniHkEvLl8DSbZmLVU2YRw6CjXQSoA5VkFYTjUztyyHR/tyvcV
rX7we3D+dlC6DAigQmSB1f02z9MIVZhz2w/m/x11Zq90xfEg9BoblLGtp1JH
y8fAgTbcBO9bmgSLRT6jjypzEaIQqouDqqvaM89ddC5I7vPqoGg7Hwq+axZs
99A7OGfkvJjyvPwKMDhFcMlC0NqFTRk8DW0SloPQas/5qgl224arR24u9252
VNI0xO261ZXkHc6eXLqC++cra9Xug09ET2BTEfLSW7pNyZDSzd5Wwy0z8EMq
NKM1q52uxVbi1N29ch97U3kBPo4ZVhkS87cBtcLF/qjBaCj4jEWEOwYbQmrg
MzG9/txsFpLPOGVqqmI+s1YRHtRhC3cuByB7hLe31zV9ANeF0bACOMS/Su8e
y1pUaILE/+hRcvLRR1d7AYuJxque0cNHKpn1ydLz0cDRwdmO1YFjSLHrb+89
JuIalp7PtCpeHCAlYLFsDQR1jw2KFxhG//n9t+9MRPNL/Drm+i+h3+GL4USr
Dlivql3Shia1W7JtvfLMNzwYz/eep5FjtETf2pyAjoENnHzXG1l2jcqtO4Yk
MC/Px59qVNosnPnBt65Zevqjg/Wp/Ynr6AVhQYHc1jqjkfRH9QfoOAzHZe0h
wJ1806V4rCszBuxDwGN0NSczebLx0sqrq621JTYWC323qJYiJBh0pmxq4R0I
wOesdDxn8PeWr+JlhocecI/hkoFcz/kcbRIVYC3LHamSPQ/dFmfuBbOGhB/K
rItCub5BSy6AvC7qjH80DVrek91RkAIxVdD6rzy1yCcrF7+78PXgADPQ8VNu
3C8xJkynyD1G1uz3nSr3ZgTQNSvyYy85dap1Ac1ctK5G4rzN4ubZ8zQgwupL
8vCGhipT0jhY3qSPgWXw0MEfN1bl9mdrj6hLPuESXe+xSWYRgxILwZ/mo88M
sZqRjDsgTopz5qIscC7Xh5CYPtEgPBHf1EepdLrpbLv8jrGxYyNxeA8/tXeR
nkJ/BUhivaSy6H0j9fO8sFhvcuDgMjwp9p+ytT2U8GhaE3fLxvZ3a5lsDSFz
zv0tATHMSKMoDKu/Si+j23WZJzTSp+83XY7HPO/C/sx4YP7I59tKHCnfSmTB
+zGm+qlvwewjV/+APJ2H/umOJ8mtSmU3JEANwuOOYrd8ekzBQuo3NA/JxicH
6bMSmhbgSMr67NGjQoccPBsdov18x+bk5y0vuN57vrrlDdbFE3iE32WzrgZ4
aIFY9QbM3dRNGzeS0f7uYpY6ooZZksjWtA4K0hXIkRv3kAzZZU4qnWk6thw6
A4VFWMxYSNGNWqjWIdRzj9od5oX/7RVFUDJRwFjNHbmo8+QYxpfAcKqbCS/+
lVCUtaVMLP5uNVQv2uiSawqn54zShzKcHKAeN4It92SkklsTjg/af7r6+HQg
wlhaRQzxxyDg2VwP5ywI42bufGGcHHrQaW5fgBdkjg6spuNHaKXXAJyXRP/z
xW/k0D/tBQ5rUfdqotxU1KvlcmmXwef4iKHlHu3O+mJwUVnTmCWalVYzzn/d
A7ld9TK6Q5Flue0+EYkqgSrKC/LgQ2HtfzCshnp06shg4W2jiQk8UIkxBziP
luAGseMV7P7w8kFiy8PFDPym+wG5w8O6hLkieySw9iQu4bS2bVPNNmbPx/iW
wmNoSShZ1cbwoST6SOWNk/HQhD46KbYm5HZ7np2PlGpDCKkxEru43jxkbm/3
GojigNCmLh2vKCRgRRzcJCa7hXUPCggeG2x86uymxK07MFqkdwn6f3goGwKF
snhguM0WcDW2BStsBzDkPg8/MtVZy8QmIGXrdD0PsP67tXF/4pSzZktLc2MI
YA3lRTyM8MpzGLQ22UPIE0XXAcHtY0CDPO83+lOpelcKJUOrA56ClH16xvFx
mdat1Y5duIYJi/e5GV5olwa29lCU4NZ7dTGNJl1U/dUv2C6bSfk8Sg8t1wjK
dG8ET3Cqu+NrDjBahOrbNeEX1b2STrEXn9A7J5wqTztUslUL09FpXfd54Y6e
KcySsbEdzI45/3oKREi+VsRUZKagOT1UBT2Ev5T8OinaLLzUWO+STG+dEYpm
Hq3vYoM70s1eJLVUeQYwt/aB1xo9rbrkaMEx2sJSk8RjE7OPN95aAmimSOOH
Kcj/UOvFeYqFLJzPuHBYMY+xtJz2XIScg+zEcJjUrtVhcLiwX0dcVNUhfgSF
i4Tr7p73scDZGYLAiCztwv1F2Cr6ebXl5N4gcHeu4nQZOB985gWroLrPyIXm
+jDfBb7o4Z//hjOhwMazy8jl/F02TsOBRhRDHQ2on1nAI651OOeyh3MXFmBi
tYAXYiQSRgiCRcfLxHPlxsHI1qdV8ILpb8IWQGvbFAGy4euXV4JOOGqkXrrD
yKTlQb6MWw15vIJV/Ci3jt8iVFf1OZxEbAQ/YPJ1KwqXgadFiisN/uyEFwtd
6cIyUA0zIssCv35G/7b6LRNyv4vIa6i8T4E9ToNmWeQL6CDGl1QzlbmKlX0M
z0LuNfHFfiyAlvn6Rv7fUN8Kxq/WX55N0LZDeyExtlFMHFWwkmZR+TzhJU7a
pyknWGTeAV9rkJPs/SLQoySYcIlxMOgL6LdoiuPH7xIs+ym+FTSNzDjqbJRF
xVlp1mawf6E33CBfgD1S2h8iUVHINGPHoZsZWmUycGhvUN1WA+e0qmq87f/2
ZSqahGF1uzUq3JnI7EzNO2Gce7yaJ+g1LuzYWfKInJn5Krr30pmyFD99/1rD
YFGIfIvtQmvBN6othCoSdq0N6T4C3KDD2MR/nTcVSRYRCh5Zh5hEbJO88HlO
NPJYQWgjcC7YqDm9wbXFWOxKm5MOwslAMZnVFElObrOtAeflDt0PM2QqXvds
Sk+8idaW+9lVcNjhogFVtbWIJQd9BcVVCcBkr3ZbCv9rKKQCgYCkVO2OOy++
AjspP02PsiWabNsqABeixhbtj1g3JFk3gsSw+mDXtG6mDsnK4uh1Nl9D2IkA
NC/u3ROSN4pgJR784zZb1A2uedqtJDieaWPi4Qqtkec3kK6v9QzOhzbEjJ3N
mqUgoaJYQKYrE/+AZCWgk4ebt2oJQ+HG+yEQE7eRKxRRxkO/QVub1UNCpRzB
kUvMNm7W7ZRhqZ8XMyTVouvW3QAGMV49QZcjUbKbiKQE0uUf4pN5hJNu4Qgb
mQrKNNk6qvVmtpK2YBvahEMTZo/2Rrbe+TBPIGNlq8Qv3aDl8Fm198dL7inc
4CiQ5Q0DHTm01JjwHw7dD0ASwGm9/tmLUdHIhrhHoc6ddHArp8quo7ksIlCK
vc/EMRHJi1BN7yp7QTXO+jG4+vbSChBgwOtlGhYbTGcoSF2/WXSC3EmRE08C
UBAuIzN1cdXj+U6D8DqQ5LzK+ltmqc5wIstIyxXK/Kdc+fW2TrWOzn2b11Cg
5X0Kpwz/XSFrZmSUNwAFz+rpC7fkVv2puFfaiezpxKBIWzKn1MYh5Ap2Mzil
i+PkNBn04vSGVJRLF84fP2TbgYJJdRTyM5x7QwIoE/5rrq/MmocyHPUZpSUH
UbhTGXpk7RSu5NLP3BYN0ou5X42NwOP1a6IABwUuheIftkECYq8x3iXzAdf5
6UICFZDGCBVy6qy04F8RruAlFuQb7WNk46MKnOSM6UxOS/l98JcEMuANsGjv
LtrPPbUql6oDACqQMwiakrtf317cZn2q2SjJKYPBk/Lf0qJbTTjfyJgAs0x4
/9bq8eoE/A1reZkK3ymd8E9o+FfxK5Ah+veAwdVCjZtos5iKgS+z2sNTk4Oa
aNC9iIQpbZswT9nFnQACDRDjN3pZHmFjSPPBGdO/EelIRMVWrI5WMM04mjSN
MGdk/EcgOG0CTJ/SvfFaSL73oCE7+Si6lexQRGAMnThaPDkzgVQ4Ee155P8+
kvY5Hkb7BP64R7lAoHJuYkgKXUDDLoqmOeHw0JxD2uaRDDowHhKuRNG4Iiks
k5CROGpLvE8r935eC98xMQtiTwlcxZfCcdW5Mghg0N92qN2rbCkvnjMm2zZ0
gUFXh1sdM5tbNRvsiR/VxyinjlwIltNTS9o6nGD120e7SSxtAFRhdei45G8Y
/D5XMCJ3PMVm86X7C1I+WsLDZ/8ZrIUKzLLOvoYbRQ/sgE6AVEZNlnBr5i75
aXXDS2r1z5utfj79EJETuTEzo6CT0qqc4M843V5yTNql5aK2GEN7bcn6unK2
OPu34rxwa25EkkK87Wmj/fsvcf61GZoHvXrxBkOZeXvl0RhWq6NPVjChO1cs
mKRRztMzXa//rjVFvzcR/Gto0V3AUYeaG3lOaKd5MBnX/KIDTK3jU92XJ7yo
2kVD7Czcom7/HGQj13ZQ8mSBDVkQoUuBlHB3N2PNw1HC7VNwq0EUJKLG3PXy
lvGlQRGVpE5axBVbAF1tm/9MwDRgsPCML++LU87ouYWCOqAPfDsGOy04f6Sv
knRUAxghBwTaJdk5XBaUoYGhS9tm8NCNnGqcwT2s0njR+QYGFP3N4Nj3PnAf
8CB9KunO2ZUyePwq+3xaaMELddYx78R0/Co5A/pqJpoLtf5T2Q6lG7aZOF2o
Y96wDFeLPKNBIXgfShCbFYhSbk2hjZ5LXPt4OyAwHdWblOMHavkHbm/he6tY
RJbwgZV6yKAov6NEOxN/uNnMzCUZXdRyN+5rIPu8BGmGGb9CrKqkcfeZY5NB
jx5dk/foPjSZBZCn+HwNc22j+lj7xwCIJ+gknKEAlkz2r6krCoMEHJDdL+ir
D0fe0No36vqglmHknCwtuJ4ev0kw/xgBahyS/Z//TEyljoM8AN4kqi98vvgG
/gXeyW2nQiuqEdoNQalnYSMfcP4dnOSU+1+6xUfMcGT95PQdo40fjoHP2pmM
1SFF1nRQbQ7zF2BOCwMAlSYdQ/kCQcYttRvLFkklch1wCcah9qzHuowIFy4o
gGyq23WKXlf1CEKvPBoVcuSckXWOT8IPvD5RA2cu4ZjgJ+LQV4m9ytWPKX7a
jKcJjLuw4su/ue49tPaOcuGVQF6QCmTOTXaWuoxJG5QCJz/Hy98nz3pFQhtq
SkJYcPY95N7+8cnHpVCK6JDm85K1uj4zLRshW2pnVJItDOzAu+mNyy00DL0z
GHGZ020hub7ZvkK69EfCw1UKD0KuMWx28AT14xzcBiwe2MURjOdQYf0nADXg
eeAS4MtxUyG2ESQLQuaLRVeQ9Zwvz5Hidpcxku7kQWFmrDKHpylFmQ2+ZqFW
IckscOzBldSEwhICtM8CisbOaVc/bIEmUozrPcHh5IejV3Zj15m1guEd2VOx
aP9A26LEicv19qUjxnD0jks/7pHORB9YbhQ6dfa4oOHf/JR6joOLMLeOtCl/
Mma6e5Uc46FjhGMTACbCyKtHz95rIgDuxaoS/ID0JVHDtaY756BPPr2/YLUA
Q7k6uC+2Y+ay44E4FqcseWvi1imQc9hSVhkmqL7qQWgCohLMVV7MdhQEQ+Jq
3bdmslNmbNnYQQM1hgXTRusCRZAZqr1SD5ftMSzgH0Dga8slNtiZ5G4of54l
RAVyARAGDh7rlbZqEY8zZmwT5h09TzsmypXd6UHlPIttkufS2wf+1bwPuwVe
KVIemSeVm/nw44nK8I5bhaEkal0pcNpxOyNl9DUV8Ek4o/1ksFZjgtr0I8Gf
CgD3gXF0tVGMmz7xb4Pj4qdx7KE1MJrytlMT4ra60qs88RSzpuk2Pth3x4Zk
AUh4ZD0bjILNcvm1PLMr2O2XDJHpsPi6/q0NeCxAfPUnsFW3QVTL/9AftCN+
3xZ0uHLns/WFpCVx9Ban4UioDyZ0xbU9bLm6YY+4rRYcgoAf4wnUmj1OL6dJ
AIl1nAMXRfiJDKCCxNTX1Fa3aELvj1U+1GZXwC8ThUgh6eMLSWznwDDD5Czg
ZupRkEYJoJkRR2jHCx+ZalvLUrSqXyoEVIMKqYDksT0QJX2u+vXog49knLt/
0i7S0KHWjEz3hpSWcZEpoxIVWMlYMfLJVwE/mvhBZgMmOVMTcoyDvneWgQpD
E6yzT9LP3YLecTK2I13U3PuaSFj4VoDdv7bQxuznMc04qywb8NnE6m151zUO
StyMkxKwHthQk32RwccNiRMPcDMdUVRBCO6bK1tgo5FENPqqVKATHQxt3JI0
+vevwICJt8qPdjJ5w3gGTV0m53u0mgmkkyJpAZU9n5fgXj0fUOJ1+NWHsZ3u
EfYN14DP6OrZyx54FfWZE3cPvQb8w2HZnUNxvX+fT/uSV21fpkbm24dfAFmB
CPqcL/Qj/TnZaW5oPfRjApio/eB8RTnwXk1kLQQwCdT1dhjmsOk4KAO1n7Y8
3g4Mf0hQnm/EFqBPdRgcDNetAZPsETV5O4JVclM9Iqh+8nug3fveS/F7k1lB
HmSLlfyzK6EQ071DKTnvgKcPs8yNaFInFJM+fqg52zY8Xbg61q4J6pKK9SjU
EpeZot41ojkbHCtF/Mf8gdQe3qWcZ8cC3R2BAIGyeRkWxWGECpBKi94sV5B0
PmfLslS8YXHGbPBSVlX8tWcLh8Mum49ik5YegSSDHo/MGy0OkBICOLft0iuc
oIMMfZoRugsKDmZV1q1cMTOs4//UrjGV3FFwWCnB/8+A7LNbZdOrmyTwhvpN
JQtt/fQ5ljHHlff1neYTwcS9Z3yjx7YjYJjIdfyJalknSRD8UBllBUmA/2nm
ePDWfuBquoGP8R0s/B7OcGXa3rrtZGWgAgpg6wS1VnenjZMntQRMAWv/Z3B2
csYf0ubctqpKWw8uKNb4YFvjgemkHF1BKxUArs6UKoc2XpUVn0eJ1gMklsjl
kHbeAITlLjsTlrMqQMfHtIRx/zRat2WIk7Ja56/z2rO5Fvc+mm5mAeQPkLg2
JysFeOPv58F9rTfezCYS/Gb/fbWwJDw3XCM4bu/ylN2VwNnSe3S6k2dh9B5P
bWxu+MJ0F0MaecokrcxlVA+ou8YiKSQaPqHZWvrgyJLzELf+W1KATR8ilrDn
l75zX3Xpq44txvrxstIRZj4qdwyxSR3rncDFZh6loZwEADFg4DdIwmguNe36
Lh47feyR3AArMs1vRcZNX4MUNRjeUzfy8uvnPx1Mgwq1+bw3NwYlQ88PpTVT
bdD1SuiAq5UjkYt5T7HFdvfMHL0qPm+BVMtMopJBI5ROv6D9X1WyibuKpgZo
+Yyj1ffvgZF3AohkhedJoiJfkq5LNRpHgmd5VvEqS69iSjjg6AsXdCBZMFQE
brmwFk9kjdDcqO7/3eErpmIXqLFfqRr1MLW4hopqBjasO7JifT1X788bpzxD
rBQNcc0n+WyYvru8+0UsLwS2E4dNoBXyrQ9B6qiGITTxl5/ObbRTWYrynW6H
RQoYNdta/Nchh3IJuh3A9J+/HoI0zHLJ6MMB7vtla+d/oTK/YUrt4x2n563B
GoLcbOy52J3fDCGnZ0+v5km+w9LRR47p/+KzA5FZyWmsWNd+GaoMv+4+G/me
Id2EcVYn9PdXIxNdauvMaIomU4JEypxWx7vGDMzyGKfVfhkgukHGpvUrtdpD
8MwhsneJ+OcxtXJkqEoBr29wrdLTqlU8B14toUvECqxd2Gw+eFZrory7pBkl
1hS5MTftYMsdEO6nqs6HJ0cdQzeHx9houJhY8ZHpPIFQOb/fYOlhEkMjqWP+
yyqCKXOm6SlO3QHGVdPdTH9gf84YkqXL4ybVbs/X4vmQqElRSaD/PBOZUpS6
pbtVsCz0nAGT/ir+6CXofen1CPpigRw/TvktcvwIIUlwxvU3g75a719gA+Th
xaSiANhjTJ1C2h3GUcvvXZFTKcb/0NMvF/GOh1tzW9sk7qn9lZnAz6QOI8IC
qAjmS35yCHq3MfFQRVfgJ+DPpjT88K2CJTpLelrTQpTTt/HhzApPF+akz0OY
wgXsci7ZvFooUs+nF33Eogop7qkYXAUn6QePrwvoL0s9lohC1pooLQzB4iXN
JcXX7y0+fEpHkDdwLIiyvl9KmoDSswO9kMJ6vAC5Ii+rQRwzs9vGhf2kScjV
tTVupLnuiCmhgpPmZljFduGYLEQJ5lspZ8PfD6utcyWKON4oQa3+SZvSFKS6
gC9eWzAqA8g8ctW7nIjyTSN2KDJZKI3YO8at3lvwTDYh88lNnqHZP45buGNb
rNVbE+pN9NanmOhVRwPCzfPO76jXssbUAbWErvc1cX1sr8xOXrDVuRNfFHNq
wetY66Ib6TNBx6CxLWURIrlbjVa7Yn2kKvQOMMIt2jvTDmKMlvC0RH/kQ030
RKQguc1v/tQ00dY6377NNRV+sAj5lKOzruK01FWD41LleVv3Owf1675uE6Yg
oSnaNHJVfOUw7A9XYQKrAskk1dk5OR4pBWO/hGITqk0CBtKedkJ39Y08BGWc
M5cwJWBLC7vLJq8uqP33xS6Z1CKTR4AAGg5x0rhpo3q53fOUgsG9RpxKbUmI
Nbfxh2gC0UDVU7TXI6pvQfuZ8JZ4ddC05ScMsAOfRMPvOLfpYyNFlZ0AGhhP
thrL9yNAR0dSlbeYcarnhkdI5jVCux/JF+QaSAoUgqmVumJT9UUvAZzKMIrO
GbzAQFrUyuFWiG/qvnLwFeZ+rAPRVZVd6+5L5fliseW5mZnOxyBXpJZHI4BG
YF0oW+98MJIXqFRNgKpGgueBg+3AiFcb0cRAbUmh/LgWbA5rVZvRMw8nWWxp
CkbxaBn/IYs1OokkpwnW8B8hM/CQZ9vUm9g1OY2VsXoNt2uoHbBmKgPPfI+c
1TE2Z0ryp6yVaA4y/UQNA3fjvi/mNgRQ6s2YKUdkPLkrhvuEzJNKuQ1LghVQ
EPgJNxkd5hLbqElQ6+CIrThGEPZPPkFJ2AyCmklR1Yyhx+la42YWS5Pa7ABh
+CQRR5QVUZBhEFhuY8DmJFVm1rhZUHBqRna2d48UXq6dzFSAbocLkGYFTcl9
IErz1IBh0glZ+BiXc2fpzBMdZsw12kzFhlr4xZNORXtPHxm6Qa2nhF+fp2Hc
u8VcHCBVFkXC+jov42+a/8Cd7ucjGsRa4ANpHrkyxMms648wrRi3H0hz0Jk6
5+KobkIUwLKjOiJ9m5X88ms7UF2ssBiqK6yTaPTY/bVcwkw86RxruRAsFaNL
D5zG8DK5H9UbLqw/O8OI888iwezjNFFoO9yJoPgj28oP1S4phqvrWIOt5jHP
GXMHYcnV/Y3ZgE24HDxY8BDCa/adbODejU7098g/D/SesSSYHiDfX94nnedh
DcXhYBS+aNYwh1EBWJjUHnLk3Lg2eVqd3TYTZVN0b9eLnt1FaBmvXjbPLDAo
eJYkfpHvWj8d5uGWpjhggBYiwQMLaW+VEVIgyymhxOsJeyHvHSXhTVWQI40T
tstp6K7+n2APT5gWv+Zov3L7rcrsyB53apHv+ssG+w81sKRkN8wTFJvi538V
utQoqlw0DNcrb2Evs6KYK7W+rv27nZi7S+dMVsVIkNxbVqhAkpes3Mq2CsJy
kbtCYDAlRavZ4NlERndJK5RH5stvJP/bBz/ctmJtnb8Db5W8tPgZVM1IRLWg
MRnI/H2oq0mVK68K5Xk/aHSIhPY8g0lyL07PhXBV6sWwUszjtbXpsJoEi5ES
OoS/3kTtfaiZjXswZ4bX4Qn34DD01WPxLOqGfJKIAxp4JkKo2Fcd5YFfyxUB
kWjDshrsBYVp79whIeexFoOGCsYC1WAyQFDYdbhJnLKRotSa6/Y9qR77OGxm
QkGe4Ghb/sw/q5ePMTPkGcNw7N5WysVivYXh5huEZQEF7tZyBABXzTtJBn4G
DloWYU9jyz6ZsrSh/pifMWsKZ87iNCnrHPkzPgDhanOD3N6itvwPHrDgtmMA
jzAJz25Smo4YIaIZTl269e+31FdtiWAh2A5EgmcxaSqkYbfBkoHOn8PFI0/a
AesxxkL/+hx7gtGXGZlLwyTFD/G0Qergy10DM/hNtMEYogxzdcAlIm6R08zz
Fsf3ZOJ5ZpAYgSsecFPX6mIEMDs6CANdXpi0iQN3CwljIdW3/bpWZuoVIuuk
PNVjcvKEJ4Uon1HkBJerVIGF4MQFJ8maKKzZVC58HU3Ykm5qq4F3Qiy7Dxml
29QE9DhcbeLOmpzjP35p/j50oMmX/9yN3GuSjLaaeF5k7BT04zIvlOjdV5oB
pvds2jUrabsqaS++DP53Ad2Fbc8pH0UemUD5Yj4xf/ISjvBaKu5j283sxtjW
v7E0O2is1NNkLM9B0OAQ5cCEgs9L91l3t2R7PohFSM1+o/BRVXz0uEwnLvy5
e1bEBF+vyawVoZvtGAjclB9XaQzJMVstR1as1uSHpp0j1XTBQfwvCdViqgf1
sbYM8MinKmvXHRvrFlHFjxmSDc4w6rkDj1+7qRqpsSZ3i/jZxOnvIkjOrH/e
CdVNTPVeeDIUlcnCfp1bV4+U+udp5JwGbQCSFea4o8JHP7OUOXV5kOVP+uu7
7qsYq5njV4OEdUtvCjCHl8gXqmXWp7j//PJLsXjcCMyrZ6TyWAKP6duhJz++
RRO5M7pRLr7JGXBHSEGFSPAJTFvfZzmgiTGuYzSWox9omIIX+Ob51VLD2DUk
UJZcgANvRNtlZ2ritM1KNJRVSLRlk7gumzc9hN0AADeltdBeMKYqydMI6RBq
OetvqQu7gYtCF0qwookhj9myHTtzLrwStOCT81EsLdIIaeUvwGqs60MvS2kP
Op4V6l0z57Dhp4yf/KJqFqlNuHk0e1hoktxrqfXi1aVi25RWt6qDNhwJSCHC
xvI412zYpFZdXpSccB62KGdH7jmM673l1Sd4/eaKjJc69FsDs+hmxRXrDGjr
uSczncm41oD1vPWfSEQefOD+AN6ijfQyv0vD2ChWb3C3zXql04dMb1WaZUPw
fuSXq+Z6hJJ4bVmYOitDiIm5b1G7/abN42ag3tb577lZXavJEdcKkR51JXRK
l87jhlW8QuEyQb7K3TQGOuyv9yZ/CGW1KZyjsdzvgfkacCDrA9OzyKpfudAB
/o1TiDSu3MAssc6swGQdmSUusqBx5tLc56BDfBeilQlFGY8shyQwGSc4KAY/
0sgntCyLK5sOm6hcreW+D+dqSQRKDtZvHKj8VYhO4NSPHx5zFGhLgtVSub6X
Nq8GUOOzS5zEQXPlKNy4lCZsHwLUXkIsqTdFRN2DyS5b7m63H5j3HP5LNwwa
ixLZ0caBTkz6TksNEZVqwV7odUBRV2k6fv+09XBiRV14SDI/Sg8HnNfZ2xZ+
xrHw4y5EFaTa2YBzs12QoHLJaagAg9WFgiEn+Xnx7fXIWzIqNaPFfeOHqlhk
BbtlIaY2b+hmzRNdS7sSSrV7/E3jI9DwqXCJA5cPfbukGLU4wW718eASi7an
PIXG9tc9HWU4HmZT+IulKtiJVcBmNegvtIJORu0Is0vWjSyDeWLTUMLTi5go
OSrrt9gC1+O1yO/wtVVBqg/bS3bbo1EG6fPOECzsSU4LGd9P+5pU65VoDyM4
tq24nJwdCy2/zBSmuSOyvf80tgeStLWsC/BuhY0vG5ZPKG1DMg2CCtkhv1YA
ob1uy7IQCjGNdOeCaSEj5gtW9c2VKgt+bHu2hmuBkcwXwMwTu7qzUYiJw80Z
Ev1O+akSOeMPQzucFT56NupUJXfSrrE9Uk8+9p/12DJp//VHi9tM4RCIJYno
EuVFhZPTXPziIXv4BAEX1dMHDdx2g8G2vU31RWeTBu/6BSJA74e6B92kTKQT
00wJHADgBwFXxpeFqXpBiPcMqKBX8yDgPZy3yNZiJrVQFVoVBIs7eRVfksMm
ZijdXK15HvH+RNJyYUZ+PHWa5loMhzNN59a3bRF7vAxw979tdDgu6YWCd1mU
hbCS1wgoM1a+Al5U6toYVgb2SVHsbar6yTon3HMatO48TaXssD7flS73J7Fa
zNZXhczE2SAIzbsVqhAFUBHUTIhGSJBRpWWyrJmDgTo8eARbxsERf8Y2tuXd
hsGlu1rYeNkv5CBGtkp1fHv9cpxFfrEWYlE+uKcwq27KnyK/0cgJNodsCuLi
YDu7pwf46MZfv2kz319cCS5mHlq/8ZJ/NrMJDUaQG20y4odoYXG3LoXi2fwc
0nR8QNFbUyJ93wIVTv375Exet71cEDdSQha4nHKKAl3E1q1+ynHty2pz6wq2
tAcwW5YMC+Y+ojnNljodVTMiFImWUJrg4ZeG++7WZDwooT2NjDOgUNu6LGjA
VlRGbRCzlAN7RyRG4ZsULlJUcRte9qTo6YRejT48nuHDgfdcAWJECsvgMfct
U3hyDjrqv6CWs0cP7Ymr4b3C3IZ90JtJpPZ3fYcdRJpTVz4+BXBzBO7rzv90
4Z1FaWlnfUN8DSFV1GbqfYurKubgiYxr6uj6RW8sLN2pgC6Dlsa6Gnnon3Wa
MPH1vfQCFGo8DzFdlSjGarjVlcGJCmZqsCFrWB4QDxEW9tAtEv+nwOXQPop4
+vegKMY76hwcPZtpmUA/LBGzyzhUSYUlD87kzzDB9Q+FEuAuAH2/g1wdhm7q
wKP0rElPWvKhOzR8ReWk3+G4ZvzOcbPuQbjFP5Xut7cgBDy9J8eAYzopVG8g
6mfLuNbSmlE1IGz4P/Na8kIGwO6rlC36YQyCQ4IIBAU1GjFKeXv0raaR4LSL
EpYmnWv2PeluA5JYvttQMspuSWKQld8JS1mQeegyY1Z5L6Qp1h2n3i5UYbx3
6ZvGFVyoSUJq/NhR/S2ggf8j8kl5eonfoVhhhhbijUPPY9drYAuOHlApJFJ1
PgNmBwIxZ4Ew/rGVv45dDdxd5Tigy7xSCj/cYhPCDzRjQA4ZVbVu8K8iW76A
PN4qddOm6NmNMz92fcF/gFzDVqkckXEnKb2w1kCqFt3b0zyV+pgviWX8OJxt
YgZytShxNvfkVSoeK2uV0MI9tG5D0E9OmZobwN7EWaiyiTJsm6p0YOeUSBIm
Gm84uIW118w4mQ6OfqBi2LoEW5lR9kuRGg3vBJciQhdSEYyFz3BAE01hi77A
XqUbuqygIUgqZreoHrlG4dz7PgZ0tYyc83CfhXpssX7XM3PuY+b2SdNKwF1E
ix8ebY19zuZbw9RVxBAJQmKv1SPEctfxN76JIAZ34RhYaWIUmNG3TfnTeKeB
7l3moPwACSpWJJmbINq/N40iXaikuErQ+iljAoaiNmj1ef0VkhqZKfZILGHj
28ZyOW/Gwtx8FbSvD5uTEojNfGAwaiEIa4Q4Jj6Kg90RGpUoHV4nNVA14YTo
ZdOs++B+hIqQJKKBS4kpCQnbz7kMCkge+31PWq//sZBIiojmzacsoS7bSfSq
v4DYojoGU8do3rihnfdlISBOKOXCh8+5rhsq0xZHITmFgF4qHLqGse0UEuL1
qvUjZfnKbMMp1ZAL/rYaTJnz2YofpjM3hVlQmKc3Wup+Nv0NhQSEbNAfaBId
Rf3wHtBlqoJoXat/NYYWkZWtzHUJI35BkWCxYJbh4Tv086YJO3xshqDiM/wu
+ODga2a5cndKD7clt87JpUGf5H2zt7fLQHQGnX2Uu2r0MfhJCqTDA6FCZvj9
xV+bCs93JB38AuKudICCpI+xAzrzQgXFMnYBvQfBlsgD6ZjDGIOxxSa25BD+
eRxBhxiaNvSI7xVkcKb4eYWHaWQMpcuWyLKqbpdg4IAjdKPaVjnSZ/E5JJNd
clqNMIWaxUrqvGs2hCJUpHSeeHZBcDGW3HYedb5+9Zmx0lLjJ+Sb2vP6u2DJ
gnpxUuLxNPLQj1LOaYnWrrYzEZpAZ0APTo1Bsn9fKjaMgc6KkbpzM5pVTm6q
/9jQpaUXDHklrGk6M3zPE5uff2adqGQCRxBym+Geemko5IvUCWVkb8jwBbAL
6ONd4scfs9ps1oZbaTBFZz2YVeR4pXqniMv7l4kmh97JDyjfOmh4t2BFrvKu
KsxOEZ3wsLwSC6F8U800L1pnGsupuuYCoPC5n530Sf6NfprSz9dQiVxNrnqn
dnPD8cQ6yjXcDmGTHLS9Ps2SeynxVJ3KtEJ7i1RJQdzySxmuvm75iNvkXTKz
82Khkq5dy8ee5CXLHV550Q+VUo36Ea7nDT++Izlu4cBCKZT68kCze1p5JVGy
TczL+2MFjpz82u3giBDtmlneg1p+rSAfNmepPzNDkqGo/7Y+P7BR5OYY+6TP
rK7OsOlu+bOh5uKga043qd/4Bpp8M3CoK7U/oG+SVuuMMKTjkSRnyXQW8UGK
N1xrCcQoSb6tI8EAeVys3GQy1Nhvlpy2Acaf2egylNMWNtR+xzIo9c52RmxD
KyWg8LMXntep+mNLsLeDszxQol4/gdNUBBbA9Y3m3PpZGIcwXJ3mddSci2Jy
b1xx0mH0Pq1g4ftxAlG0xrJFn13SO27gF3X43YiiGMjcDOOdTsvIhpRA9bnS
7GpbXXX/SkbLefa110uZ8UXT0ClqvkP+koOosWCjN7iN+hEfT3Y4iY/qPI6+
7LKUTtURkpOr6ztm/3jxIVf/ZRGaBWMmsp9xC/C/dUMDX5//kqlPTRZ6c0yt
WolcADKc4xgz1rnHv2HN2Nt/7KA92cHVkoEQMzVj3YywMtpAdaUgG9QkRHY1
mB6zH0dD7GeRTMZo9sJXR32GhoMCb9GrI7DNbBnOtAMhAoOqDBatnWFQOuRn
9CMDEhh7sWMQ16s1Wz10Z7VGRvMT5mDyOxh6zvZ3K7Xt4y/n0y2iPd1gZQUa
I9CynOSpGGm7ZVeA/2D8q2FHKNHqTB/tkLETDpmtGzKyMoJJn1ybET2vzZt8
HvLTz+YrZo9iIunvlytGHX+yaV6vcu4Nd7y9pgsIKWi2HPXuQe2W56TRQtOb
vaeHwfjNX2zfhFoabQdJ7ThD7swa72wTGfVwSL2MgTLRMcEZWp4jT4uDLWxL
MDIxlPaVeqQcrlpOUi6K3w84PYMJahlCTt4YTrRv+gJ4mYdf37KTCOhkkrkj
xXaE49W4/aX/41sQn8/q+9sQ70vrdyZyg8b/7uebnxxz9LFnZGSRnUTbj8TQ
8c29WNV08BlzsVvoxJkyNLf6/kQg5oMP2PZvJoHdurtv7uFhU+iPO1GLMejV
BhpS6naQN1fjX0t/bjQT8sCLk2d7aCDAcWtvJOqCRT7GH5iKw5MLBGQK8L8l
EnmYzENgDF551o63Us6taSCMM8PA4xwXbmGHXn9rqEt5ny/sQAesiWmiOt5O
Q8EShhbUEP9At+BG2sWNKGYXvsYK/qicaUTemKoaziFkU86jIXgkL94W1uK4
fcYNzcljky5PvNlOM1HIVA+rF+DWHSuR5QTHZb6GQOYxgySOtRKTVlFB75i8
+S3gbxPTMEN1xSJtHeo93swEW7Oh6tG1X6aUeLZU1MOof9bNcX5FUrLDFYe3
C2nzJxsh6Nxx/xhC+Bi6AAm6EtvWCc4KNVdDNVBEQ6Mh463CyPNLYhC5l6Vx
r/qydBICV5tViyO4n3rIzMnIDxwgIZVDYxiETj3s58VVRdstQ7tozsHQjqM+
AXHHGUtcv53VvtYvPei1awJ8o9LBWWF6YENRoXguwmU59quCPyNCxDS4RXhi
73e6/V/aTtP7uEdzJwtKFvH8V6klvSyeWBf4xeQWuGD5u3q280ujS1yTJxEe
5AKKAOe3sXUO2ufBF8vLKNDGNQ/NPwL3Bu7BoludLm53CBoD5OKjOBeLghsq
KOsTuqPBe+HzvGqytfbdm4ZVnsSPJCb7449KfL6umpIU1mpAt2TC9meFT0KC
S0FalB9SC42Oa220SUNnS6guKJZjh/YxuaCA+OmeFXuFubRpoe5L/2KwvOgu
9813UOWt3B0zyPMSXZsBi51cxZG2GfdClMrooKfFXccBo6wxpIAXkgtdsupl
QYD2Y5rWzKdBfcwzyJ1iCMEVfTc614+qdhe3h7oQX2OUoV/72bQFC1jvDyEl
FwC//EnoV12kR7HThXFijprU8Mr/1Ym49o7V1YNRudvlb6xU1b1sfyRibPuX
SIQEJEzX4PDHGsehlmjHt6EJfroyUaF8kOljKE6OzdCFeEobebJrVLcSZr2E
osYeBjLLxK/ASb9csdSCl52IR3z4SI9RbodhnMdtsQDZ5Nr0JDmgjCQc/2c4
zV6lMJSMm/ri4lYzwYmDyY8l3S9g9O+MMhHp/ItDNFCOnHLDPSYJo8V7ByYd
TGvMmfB9IKRx2V3JLNP1aG8N9XpSroMFmH/iqM/AL3QgT5ElStX9uK4WcbQr
gSSnCcwlhztOxKVgRppU4NHLLVVPxgBf6/Rg5rnXcEahNjL6iSWX/5vfer8x
aZpPAQUbBZx9aPLSv+oRbR3BeQShCve/zoNqz0A+oxjmr9ps7yEj7/jx6JTW
bc8Bpw0ThHYn9pg8vlfi9FfB6wUSM+PBwNP+bUL+UljAYG1xLDG9jCjX3hM4
mJHSkH0pV/jZuSyvKujYcASrBmgXehm1r/dcA8/3gPK6SJUf7Ds9OV/YhPmD
jAUuvQ02MpdPV4YQSOBKKdVFwLvY+UjjqU9eLXHAYtHEVoXaXIlkXJ+b7Dop
8ORYJD+mkaqTRLdvfkgW6IZy7eg7TNuonMh9shgS0Bm120sg3KVxK4uLM1Dv
g022lF+j69UNxj/JQ6k0F5jQpEks8OxaIu9cyBFbqwG+4ql8w8ckRgq7fEyq
gaYm7EdF+aJQFGN3RF5p0pEE5j7zhZ01rqM3H0EJmhecz8WHNypW0xmCidhV
5HDvHriuGfap8pQ/W3QbOzFh7mGeIzAHqZeh+1QJziB3ViV7aTIKPlPvIv9V
WRrC3ADgiL2eyVGMMsQPTE0aGOwsdkdlVfodMXd1usrTnJHeWl7KOIu9iFUe
xFisOEkpcRvx9HTQpf5kpzTdYzwlf8+UE9fH/KVoXNrq81ZKF85hdZ39F1s8
Z2CHvcl8/yenYlx+Y0qNMnGmhgXn3IBwGHx9hb6ogtybkkBJd8IFsZn8ZcRr
EMFROeHNL180ou5Q4aheC26rw2l9CiN+0ab/sd+0mZJpRfR2g2dxdQ+WIZtC
5MUBT9BKENNWaDtpW1W5kaV9mGeD2DNEZfScfa+acAGdxUBAxcDLO7q2QZp5
ZvW+wQYeWwjP1o4X/0WK95Zv5RsKqGIiylxKamPXEDHGKE2jBrz0wZhsOkMH
3W9N/K5FKv/ik+B/zqe8932hhjTbu3Y7z+BeSW+fxclxsff5NEusgMB6+x9m
ww98OJTXrgxvkZHnd4o5bvmMfxCoFHShT8/5l3DtVE3AVEtSyFj9H3ikQJXN
jzYwyWff06A36aeAQoitFM6RS3j8V3RtfXw/9PsWy6+rv5LjvWs8lmFu3ruq
6d0SFnwPCVHdDumepaGxbW+jccKAIp6BAyXVWQfjfgTlkHCV+P9wbyQZL/2R
Ojs+u4Jgh+cJ35xa/1vQo/owPvi42nQkPP4IkLFuxbNiQXmsfgyAIsU4h7js
tryz7kvQu6NfdWwhYUjFx6cOTCWuvQO4kJIM3XerLr/HN6KFJjAsn5tjH46q
l8AFUR2oYOvod71ZDk+YgJYkfYERNundqConAXGSoNy1G+t51sehx3X6zl7V
1FK+fDg4f8FJP36b2gzbAGI8+vBNhpsqekds93h/nd4x6EpKpcHPSGRHJnId
UToQr/O6AX4JPNRKSKl8dsjdxLR6wJWcblc+8JFTvlsQhhJimHuEuNF6CgOJ
LI8U2iTkSm+76vp0ia9tZqbtPTzZvBYJyIAOkrH7kFgKX1G2/uxX29a7duz6
LgI5tS/WQjzPUC6Nzxt2hEMe71lmDCcYUQ/0jB+6BSIVXw5PaHQluGgFXKbS
PpUqMrhptPuxRVfTPMzEwWkW2UtCiTKm1kROMzzVbySQV4YQTJgynYgXEB31
nQsWoVbBlypQ0XCBGX3vSindE7ToJ3BiX3wT5l2IhjffsLXq/nILzd7wcvSc
zPvf4wuoiQ7Uf/3rNiAvX4IpPCaJaLgoshS28EbshAFAr1xC3PrC9sQU8q0e
MeDq93vgeVRC0GxJBm2877Vh5YAT5x83XalhmmjYOzDDaTgwMhalkgU4EOQC
oxFdjqII+c0OcMRkesCZHrKCa5H2cihuK4PThFXFBD4zKekdw57oINvStbfu
tmAOCot7uGTu0aWcNp4TvEueUWuKnYLkzlk0UKecps+iIqt3zOONsJXV4qKk
fDAZqE1n10G4JbYCSqLhI5UlSCIekrUfqQimyie17XjENLieZYOzflN+ySnp
sSU0asU7r4FMki33M5YuwMeznmUI0BX78IhTAtEMEdFCIid4RciYWaZP0Jv/
L/xP5OtGD/ceKDvHW+BaM3cdvrMtJ88KvPhX6v2HDD9B1aeomiPWqpI9M2Xc
3RL26Mw7Kl2st89C+qu1WYGeXNiLdpH7yo0RY8dKn5W/Ns/abKYzoGTSSDJA
nGbdeMZa53D5RyoWH6YnYdg3D4QLjbgh9WzczioCJcT7RGvEA3uuMbIPx+DZ
Nw9TeVwupyJ0ZP/c3N+y5SnAflVNckRyvjV4NWxty9uSU9tS4PhpEYX3+wZm
aKBHC7Ly5LswQmmQEAAUYtucVMS7WzGaSzH6ZEyduG4FhfcdqpzMED59MEGg
zpfGBjXsa36DF1wNtoX8iboICwjFlyF/S24G0fOb/BLmIHndQpA5nFoieDwA
kvPPf6Zpb6UmyUKgIg7yYdg9fBTrjLyXulIxz/FCswXzLjGoMi/DIVrYt3dz
BK9gaxsOgYZHxJxvAyAZsw9We5SGbSbU1AbZuXn9v9p6wn/PefN9fZcGdPM8
Y3LO6nhVazrxsMQMwh2sZhVrQ9x6rwlnKNcHjgH0D0hJHSyjbH3/K2edJYNj
Phx+fmiJ2+snT0aid+6d3KXWOaLcQjMaxdcS2Gp2AECWuMGkuGzV3oN7Zlin
5w/BAEdNz/HJNf8Sf2xxZrW1tEq69BKSlPhwFac5EMf/gYyGAkczQfnaVimQ
/Yl4/1zlM/WrGJcis4Iq8zpLaWVSZ1OHBvFJrl3IQc2aVzgJrdHwsyH6eBuN
TpgatDqNr2mES3Nc4S4Y3CNF0ktCFWpHl4w6adQiz1UJISPlAFHjcW6YzxNk
XJvNRowML1PJlvb0f0iGFyo1Nk8wY/wXdqwck47Txo9+UZI/QhsEGaL5ngW7
SvTkKACbgqF/egsT9B/66fuwtmydJaKRPqwOiXclseYimeqvIe04vjHLrLWm
WhnhU6Pf2GbVPi3RvNsELvS5lHw95ZvBpnga+8dMTpKMr6TQJl7TO1PDLL2B
+NcIJAKjs2X5KEAhXX+DLdxUaQxQdRhBaVxuD8ibVxqgej+D0txXoh1QPOmf
Bl2MdIUpUofyW/GfNV38M8d8BHTvafBrn1hTcKYom9oGEhGsrIiOZpOWsR6x
A8uUE1v+TQV+XCsS4+452sx9FqWUxGKU++ZBwAZxHNWBCW1bJESmOn7xtzYx
lbaY4SLxhezjQgKRSXCa/XMN44gK/nk3NvGXQstY9yjqGYA2dR4yLdIqF/9P
X/Vs4WNGwiiZlM563HbDKQuf/+WzKfrDsd1f9YWYtlD/MekIDBmAoOrwIFvN
35UkFWsDAzb32FCbIamlsPYua3ExmJvkQ7mt4jyhOeUR1zEQDz8B/5OpF6b8
aYTyOIF4WImvl2C2eWFDG2/A3AywIegKefykP4z7obB33TSB8ucoWzdu9kaZ
qea0qa9X071ptdorGYk2zul8zb6a2OIW9NUUgjVud7FqYj7n1JZuAn/cVS9v
6MACKRNC9dIR41YtJ0MK1zq3Dw2xaaZ5xg6q4NP9I0hrQDtFMNfEDqo5XHrT
MvpLeJc69xnYirwQ9pak1zxCt5/4sDCF8VGiDtAdrZa/fAhZnRjVJ54M/geK
LgdKfDF0B5d0TGcqHENPrljZMSUJ9GexqfOy0KTjNRP97XwpjW4drfggE3B4
AvHSm/TOwh72zJZOYc/wV5inM3iSw9rEte1AkDi/D3gqwyWWPh+ftASHlr2J
O4RtkUgBxm2/e5pbncnJvtXff8ZtnnjYKNmqwwseDWOkafuTr2cW0WzS/iWB
EO2rN9er74Wq5wyv+Y2L/Zy6v3QoSUPPs/HsxBrCZveT+ZRVqAD6J7S7WUsA
cKsxk+QaCuiJHloDybhyEvR8ckdyy+lQ44E/H2FcDj24hdov3xxdbdpUNQBg
rczTY6kowF+V10/2GFcRPR7oXBdoP1OEKy5jKEnhYgWtHU9ctp1hF56ff6zX
jE3Y2HfRqCXtwajvm16fXNJCNBhAodFw0SedjYXgRB5xC1yRJZTVpOqdhFgt
S4pZGRRU7uo76K8Z8Vl6LdFmF1zAbDnh5zM99Qr98FxAOqJga3TQoIwHNi7Z
X6KM4qkVxywS3Uai4DUXKP7O9Vwja4w1BnxQHYKfz0dVq6Fzr4KzxpGQYGz2
8qklWxeT0MXhfGRNe1E/WI/UoeaxR/tHar4v3r1XqbT4xEP5/bdkTqDcVmTD
gQX9c44k2n9T/9o33IJY6ol1/Jdc39WLos9xcykSLY0dhk+0jCnb9oNnJwY5
5a0FupEDAwzDc7azGbA3cfXEtvXlBnYJj92Q9Yzrh71F4+YzUg1yfeREqXzS
TILBRlZMf/FzcJ5tcF034n8pMfRHecuZl6ue2zqMSGM3mQp/e0IvMPgqmVzE
jD1GaJZ/UAt5UpkoJgJ0+74CUsaTdlhSWNfgBjbvdakv6Bgf/TFAafpEtWIE
7LTdIMpk62LYBoiGPb+GlQQJdeR0c5TOjAPi4UKHF56h1rA8ZlLuAFPK6lVC
stlkkCXQIM54LXOHlD+DdKvdJ9tsuF9vPEzMyKVXBnMIc52eRc8eT+ndX4Rm
hB7qyAAG7EgXVj7E/k3mtoKstbL5jGmE2E+uxqvmkwFRM9cWuASNyjZBiujM
sZm5uEPn3kAYioq4/ApBc3fUCbvpsY+O+aziHAKdfZlrZXWSfuB91myQWiSD
s9WUGWGeTJ94cTm/Rs91Jnq8QyHV1tu0J39u32OPP0V3IU3dTUGiK50QQjfT
XdN8Wz+AgFGGlcEMUxudgEvgSpWpIyN5zDH5funt5NJZAFoo5WEJGnsMlYaq
ug76Mvy6A62K2Qszm5513cLbVEC1Nq8QLi5skGq9yZJ/n9GEggFSkXAusegK
75bT3JF5fkgnlB9ZpRCMGLlp8Ogq3t+cef9qlKUjdKAqeXTx/d57h9PxX45c
m2K3TrL+eRvyWk9s0zsr6frO8rr0Ixn+mAKIEaMYKlDY1sQKUi3IAGTrEvSu
Fn1b+DIs62x5GHjLev9z3odb0fB9FZ4/fLbBcEDf5NySdOc8MRuIwBsDDIWs
FjSiqgX7Egz0E9hNzKtOnS5zwP10AkLlmlDL2ZPbZAWpp7wM7ZG0tty5A8J4
+3FSWEAY6qRLpD3SB87DrfYJx5q3FtetgO3b8lj6cjWBXt8u41nkhivfYtRk
cbkvbicYRfNjopiA7qK6RgU5KYNOfUU2Vu9nbqxC3MWiWsh9xtTUYYTu2DFd
7/xxaTPg6+mGIqt1+SYPVQvCRZnurMQE0XC/+70gHkYg1GUrUKrfqStBKPtv
vsNE6oSl2k1PzpJWuOtJPE30qytlHLYiNdz20433iH6Hum/AIDLqVngacgxA
vs/JPsAFO0vZwpB4KyEAbxlbNHKb7WDkzjFFgxrcjDWrxPhTKI+z5noAsqq9
I/BiDrrbFjy9HNMgvln1bEYujVIKl2NCIeVrgRRoOVxiC/NxIwzTonJ2XpEq
UYI/QXyLN6e+FNUxkEL4m+UGsB4ApaKC7pZ4w+0LcbWr17zCwgu9IyvL892f
N5TmzkUASpoNOlJPvb4Wg/yav8I8gXqAjvmvwYj+Y4y92gukPjaZz7nr1hFQ
fsFY1+PfREr5PCnqeP7IAInTenuevKBpDs8b1nQ3TYK/Yxcfd8oT+wk3e8Z6
y1pNtosFRF5A3rn6+U9d/01FquhUZlw5TFSXPFc3/5ld7veeYw2HFE6siM08
8hSa3PUODgU4ekVcN74wtGu88stjg/K3OJPqCivUrkCKUMKSLQHJLGeSIvO7
6AxYPUE4ZSzHflnBN9NWt1kXGK1XfpSnQ6J6PmJb387L/YnKnoUQ3sGcJomc
I8Yd/KsIllIgZR+L/+5YM4U1gCXhTXz9CCbonFsFgo1Q0yhdo0In79G9koxt
6So13xhyaV92pNkrGaEx5ncnLIxDcU0Ot16PAwrreO1NybjZW9dY3JxhtIlc
6gMhg4pZuMSGumfs5i4zBT6kSY93vW3DqDceCtqyAbcf4aQFuYw+PBch0t8j
9SML3Yq77ed07Hoanql5PPzTnrKqRE1tOxbdYtY3D0ipU2AZHyQxlFfr5rJr
qVbNePyimephUm/S/iCwhCL+hfHA8gYNNZXQ2C2wt8SHUz54x2U97wy3/yOH
KE/mgjooUT2+/LwnE3OkhG07ktaDxY5vVwMzvidUffaHZmpaG9nqTgbecGO2
iQNYC2szkCcG/W5b7jm6BvOgTesXJXq83tJC6eaQR4Tdo4wx1YLhHTuq+ajx
1bis6Z9yoadhe5wH2/C4bUfkPIDL3A0Z32QqkyallTsonEkOXN/S4Lue8De4
blkSrSMepXG7BypMARtMXeftqXfoEZ9b34BY09DMekTznQL9/wcP8q5gFMLG
YqVQuA0DuV4Z7v46NS9rgJn5I9cb2/R8Xj6avcnObBxk1loB7LkrBvtDN1Xl
Ii1FgNzWPSHNSf3e5jv6pBrdRyOiQu7K95O01tbp86lFnNAdZm8/Mmn06aMU
ECQvJUWX2Ps8larr/6vQ04UDNrMKIEsfe6JfEsvHuSjFI6zaC1MOxKQNrCIz
GnnD9RTH0bZEg5A3R64+CqFGfFOJ1Vbyq/GP3ztbnlXYkc8X5BBybxHRlmHr
GDXvEQh15LG5sDKzV4wRi56isJrJOjU0kBgLupvronKRG64uS6tQ9FsmWIYg
TrhGVIhB0bpJbOUkIik3iLjRg+WXE43J7mBNQNawIj07e+f+3KS3IXmh5E5+
FputNhP9dn3MI4Mj/aoMzl/kfhRIJdGF6C7+CpcawWEXToo6XI0dqUmnMEZ4
+invHWQym77RCaMLeCQsTXlN9XFL27Rw3y5pC6n/zBL3jacbs4xa7aajKoMO
6JYulopwYcGvxXJJyHxAcyPf90mY2WgHLfAYKH9bcXxKwWtYI0Q6a+AppU5S
UZmrxpdBJv+3fCQWR2lXgH+leItaD+cCv0oAihP5mpMI3ppInMkEFJNn8Mdd
kmlFeLzY7QBnsBZ/qcvtO9PizDdNrXRpXk8D5VxpIMHVeirs+NDRwddx7A7U
Ga6tvCX4NR0e33OLSAA+ueyjxkmE2mtymRtPnigwwTATs9DxGo+6ePwqXCgm
dBA/WiNwQBsYvpuNsB1kvJz0Cuz1S0aqOdbGTaHsNYnoX95eZJUE80shPd8J
bjyxDpzqr8Kugwl/2jYF1sZPdLDEWvhJziDrMvk0id4wk3uwmphVFvGtUHts
o0I1UGDogGdydCFl6wgp9SJpHs78IrehctdsutxwQbroddmeueNUlKmJ+heK
05WdkNw/kbS154Jt3u7KNjQ/l6158HcakhfBaBTap/81q8f3t1O+L5CcPmmB
GEQRWDy9mlBkG8ibUXeofo0TYDAsu81eG4LpuhN4VFjdz0gls/ROEl1KIqzN
N8PskAf9cIEa/5IlobhSFZbjHAVrVxFLxsMg8FEoljKPEhNothLo7GjYfdI6
IcuL5HA5+UGlCNKiV4w3dQM9icYdZKaa6K428e45WeHp0n57UoT1nODuqOCt
RpEnhrROoNID2M7zOQ9WVh59MnT8eXaFQqueDQ2YVSE6v9Ct5EZdRXBUi76P
VTFp68wWCjjll5yxQWTaZSP6wc2HppX7N7b/rYiesu0iQKGP5HWuJXph7wFv
OB2TnwO64PblRYgTaqsBJ2wfQlx34l0Sm66O2eThRWDsv8NEohtgchGq/2os
axUn4VCZP+Sd1Y/0V5tRkV3y0DPUKGldkDbF/rtd7S2Nng0f2awvKVCtvk6V
fBvAwHyehP+HWC8TOfMcAUUklB6jB+xpvrfgUGrNSK9ojC87BDspybxeFG80
sgGT6rjFD6zn2/9+qWx+1botH0H6FuRO1U6S5dTUENwN4in3iMqGorXIhOF6
BZ8eKrYiOv11t8TkHYJ0kUCv++EzIYDgGmYc8gjW2/a2HZv3glYhPx2V754U
9TvFngTyAB0OMxgPdMD12wN9Xa3us8gylLb7gATzHf/W0P2gcw6RQDLjCI9b
cpxNesVq1qHrD+4hBJ7utMTycFAP2rf5vcaZBmdqQoPeFOhqhoxpj0tGQhVm
c8P5j1W6ZkyX+7eqPZpcIX+H5IC5QMj8uT1gLu/UKwthmd4CdgERfq6KTDAi
/c/5v/AFyYRM63MkjyW5tLtP3We872DqcDYn+GomhRZzdSoSKwGuZJwxVSUN
BU2VZbcFir/7XNwvR/BPXQiqqjp9WKV8nRt3Xyw7znUprAnEbjEKQHvl7N7L
TGK3BIntPerM59ktPM9lMqMeXibzmT7+DEpuw6UHYoSVGfMCkdsAxwkuXqbS
Iyfyu5Y28ZVaSuEvFlgD2bj8kCnQpx3AEgm0GkZeQ6qKzGlI/QVGA0cHky2u
yX4KXFp/85Cr1ZKfOr5iBdJwnLUsI7jwtldS3f1R5pmAqlMr5++XlfIfc4z2
OA1DUgnQhb9p68fym/wxva4dAUysZ5QXFEdsUCZlU09rg2Ka1fNnAy2BPZLs
WS0xRkMtERZ2TXkw7WKFVkIZR8uJ65xb23O5p5owQK9Blo3nL+rCPryH7RXz
3+FatEq37Cwwf7BxadqEcoWxq+PKV1vFTjlkjLhnqIWjFdXgs7WWpZKS9xYc
XTy5w+m+HNWqsJZEJSBvmeYczEbR7mIhKqdhXhY+M0tFjGkg64wN5LyPLenj
Y/0c1CGYzhIgInKxSY1o/yz2PJqYqhEPOda8FUjFkGqt3tIEXL0B7dv8/Qli
UjJ97Cmd2fDsY/0MaGelK3XM/MMtuXtXTT9ErfahdkrvMTOcjBi0WIJSbMMA
1PIlBh6dR9E1ktUPcl58l0NlyW7anjrfev9HXlc5+i8IvPj0z6BZcxUWkIRf
nY4KoSJ0QQMdhqipV4WtA+mHHybBNcseOgEQRgJYYmLzvsJBmNkqsvNCVNtY
1uP4mppHwMuxwww6rdSa6/rhQlzsbtQ2iLlURzEMNoTSNnIsOmN5SxsDIm1m
7LEA9VxJnFKflcDUxdjuEAFtRWORgElvi5nEHXxWdgs5RZxq08BOxfQ3lGAM
hmxFcb5qRLSofudm5zYhs1gHDXZ7vPLIb+Idbm+onzRDuLT1rxFVYV6mSHU4
GeQzMwcJ+KlzKxxj4jJQPs6AxaQw8h8vVBEz8rlgU90UtpysEjODCUBXDdg9
9QVXuzJzJtCWWKrwI936RUZpzR7BfkhM/4n9wpckunhz2p1K+2LXi2i0TfHn
nnay2BMUXTlBU5HBUs6ChjL1A8ftc1vzVbJpB3RcaBXnXokFIEQiedD9wuOH
JgmsKRkCoIJ/CPXLX+JatrvtYhXNeiTqv64JiXtfEyT98LpqCkXX7/rXFqn1
5ajAMpU5B/9pWSFSJ+NVPxCnV5cgJzBbpgd98WSRZhh00CGLRq9v6lDSzxZ9
Aqdey5/GRZcRnmliUzCu5VD8IsSYIchDsM4N28LxOJqbfgwpnpgbyCMdA3h+
NLmOhXhmBV0uCL/aJUn9afucAJeaHyigCTIWb04Yz+KjhGYygRD4OEeSei9c
yE3HdKcTMv6O0wfXVL1mrcYJlxWplYdh4WUYcXI2gofwWmY2LvGbqvxvso2s
mT7gXlmCLdD63knicsdX1sVNkvGrLhicA/7o0wLL7+fkkHlLBL3YzvePuVg5
BMME4oQY5FfSdPiz17IYnSm2HlpIZLN81wQxsLyd5mpbih+xAY3Llu1cKCfF
yQ1uUhq8s8XecncoYOoeA8IEXXqUpPItjnAp+gJzVALqW43qHGpxkYclsM4P
uE7lZMULN8SQiGO28Tedp7Av4nTHGEckdueHhXpAodVz+nvcVPHUdEqyCJ33
K6OQBNd1uq0UpQZpUUAR3b8zE3lnnelj2llKKrxGcFIfES+eZV/scEHOG7zv
dog3unoWBiByol6g+Ti6VbP7P/Um2cpe9wCqqZKM/RX4ybZG3B5ohvozIuqi
D2wd3PXzZEqF/oKfMYGxGXo3NyGkjbsnoa9VSkztx7K68C+Yop0qCAsicY3V
2juKUsghM4qRmSIjOiK5X31NZ0ivN94Hqi6x69WUDYDQm2OLs/nhpDJNSLz1
RKZgA0gJDhtuvbravuejlVWE4kA3DIhAHw8fJ4QDHYiD7NkSigEUaH64Cq1I
MJVQnHU6NctWa79kcAoycEBgym9rOpryjA2uT8tMSbm3nlO4rPfgFa/aFfR0
26JkdhI2Dc/1msHQ6IywtT/rytztSN3yU7ZGAwG46I1LeU7sMiDdLWxXm7CN
68Z7oW2WqACLqHGMMK3ntFwIzAKtYWc8sumQu8vCj3b/jWYXgl5O5vzrxCY6
yp7KkG/n0UIZuAXNQ46A23s/K/WgZ5JEzw9ivXocJzh3ePU6KImNfAR0Pjdp
jaTHDwOeDxR1j4qRYrzWumn93qfCtL8Bski2nA9n2RXHsG4uOtBbjOkHuKby
JaSb0TtZpb6IluB6izR5kDWu7J4hP0tugqt50dYZ9Ig+keVe5PKRU/+GAzdl
rWZeXhTZc4ObSrbKImFwauFcJiJ5W05Enfl4gvwT4V85S7KuGqWS+MdnNgJG
H6whgsvsThzS2e2csp57BNSbjPx6LTu/qyct57+FGIZePV3M2WUgc5FRJ2mq
49n2njSrG4fhfmpI/ng5W6btr06SGSGankfilpxhOlfNgUEqFZ2KVu7YyIQ/
Hi9Ezz+WZf/zKlYN3wQsfui+P74vpOZy6Omw4yadjfaW1NyiclEtQ4D9dIOA
O5zy2ei26ozyT1aGYiQVgn+5+3PW88rCi9diYTYyyOIOIpQVeikVkXkuc8u1
c6Cx/8rpSJqWYB7UAVmFdScC/suXVYz5Wq4tGqr+UczoZYtiVotPUr9ndIfn
OzGmrIhZ3QAZpoLDekGBAOpe6KbXHVQ6SxfEfjQt7AsCNEo5OdMykZXfsKsK
BxlFEzL/iiPPbJ2MuZyStnuj+S+xb+BgQeRf5RFqnDfmH0CUZq/wk9VYC5Xg
hVjEOt6RUrCU3dSYnVcz5+tVoR0GLGcbpXP/TU53MTTKrf1q2MG6hT64trqN
ipKuoMPDGq8uQvXrdbRudvrDpQVssv79XuYQ1e9ATv/hUAWQwU8SaLFnKixj
Hpdx7uyvMds87UIPDjtCL/0JCy3+mK4Pj3HkBTY9blcH+VUy3FcUZTsmEiwT
Tw5IhML9yN3oeyuNCZ6GGfzQSq8l3bMxbSdzcB3CG/zknDwTIWo0gFQkcb2A
cvrGx4cuhvfALvnnQiSFIfCP/ICKuPZPzCW8qXuC0XoNZg/GAU3eYMYChQpx
WW3BHZCIH/fRRhPTKuxpg6McG78yd2Ok/ePVfxqI/o0tN63BbtIf8XsdCStp
R28bhHIFuvpGU46T5dpP99FtNVyPHiI1hl1HAKHGQun+22Qy+WsJKFf7kpvs
x8zLytCG6JrbwdsveDP21IydmoUz3NAAJzfV/w7HtndqhrOmENcaXdoxx6Xb
XZLAIuFen2u2Ou5Po+XgdB0Y/1VlH2H/GbF33zfotrbigw/WmJcduMPXyFqC
lcPXXbItxm05+pfdfzijHNUrKEJDsqg3sANRV96I9QpFy4cSYGPqb4ZihJ5W
GQSKodIgQ9AxZuEREqJoF502PxJpQdGvVOOKIr284xwWn0Bzv89IQtO8BMjT
c2QYtGIxuaVLWVJyr3jq1jzjDARzvQxA3eXBfcs9RU/52s2XFjNXxdxo+A71
v/sOtHQQalcD5cxbdOBDi+toU0SjYYj1AhIlzRlnyHBa7UsuL1f166zauoV/
Rg6uCz3cjVg+4NOXKFAHHWIHTAUYpE2alMQ8p1j4g4sqHpl9SlRuzbF5iQBH
rdV1vxHZIsn52W7ZNpgXrJ2I/PgjT/4rMT9i3TBis/PPCuyvc/2v8PPA0M8o
429bA5khnNnql/yk8istR57YK7PO9DwXZ7KXSws94hr1JLysz/FpDui/Y9tr
weNJFoMU1uMVKwCqg7qem3hVxvn4+cW8yyVY62Ez9j8DmRbfxosNP08SWAhA
JQP0pHjRNOT/bqqftuz85KZShS8WKohuMWMOFIuTXdLgLCWJ+c463XFdjnjd
u6aki5k2nNOL87pqMpyxDM9xYINapyK19uRPAeI1mgf4Gt7r+LL6UzGiDAAl
ENaRXFLesWew5b7GwH7oC3uqdy+NAAaktVbm9svBMe91zy384Z7wzCdxNLLp
IVKlvwt4mvhl8rlTxJXoKFqiWihKvZCS0b/hkXRyu/ZGXsazcbv62d528/YC
Xnn6Mbns7S17VRS/wUWPrOfQkn54to/YMnie9YbUO8LN46hzhE1sOgtJACGp
T+6mqwxpLH9ZWdhMCyWiXNg4skJo2mug00Yftpy+mAkUSvNWnL/FJ1gCPtuW
btbH5cGQRGZB4Y69Nrs+7mq4N++e4SKg758FpKpL7ezURRP/Ehvw/sn4P0av
miYxb7K8UKKl5wzvNUt2x+w9FJ8KNRo6hwDUrD6xDQaKEveq49RdmmAyGiwf
48ZIIi10MohUzP5eFE8iVpnFNTdNNfA8fO+ZzqbQsbuNsou+1yQAoJ0Y18Pa
vHWZ855547PbQbubvJ1w2MquBCvst+Hqkm7Mb+gB6FPv4R8mKcQpxbVN48Oh
yaqcqY4Pvc3KDzP+UVUtYU6Oi/L7ETxNtTlGNKNIxPCIqKpFsxdzsY6shUY0
beIU8RaQTabvquQg5V/SXGIRX0ehq3A/LIGNwG7Rrwr396+ZLaFsWkfFfJ1b
1U5dXkItte/tmgH4c9Fg8T4wifcPngDsG6+W0c8pJZqcFcXM9OK3qSmsB8Qf
I7ydAugIYFlrT7LjoCRGZlzTQn7Pu1m1o30d49cqs8LJKl4b8EWFknPQA97G
iSYGoU3r/zRx0LwiHwzDD7bLmAVJ52z4aCOPNCL9pZOQS46No4KKr5MG+168
pPdiGWqmDAfo4tdcaeAh+fZ8QW/aSegrblkocXNNNm0dsqWAKp6cV06YMVN9
cT+uHPJUiFofGZ+OPj6/a/KsrrYb8WIc4XHB2HUSbhs1t7y7Qd54R6Xpme/P
AP8wYxuQoi0vXHLMu8+fIGlURv3gFSZEKsDfKRIMJuia0q/Xc7o+No7TRrnL
Bx1Ar/tUAfJLup/tbvrpWCZGoyndLFicy8tXbrPAfhgVJGsYACopJlP85o5B
RUCr4OXvT91/bJbSXkbKffpQ9pwxsiYZlmNgDcoZVBNc7/ZbqZqXlXyZmtQn
bRtZebalZG/h5P4yuCLcMl6ntrYWL3Sxgl96PQswoqvhg9thGdV2w//TBZmx
WuEocm7ybTeTsZpOmpOF+4jR81w9GFjVK4IbiLg0fdD8TYFMn4hrcnmvMIht
/W48I8lYkxaR87fmY5eK4vHS0dIl9qED2J5xOUMUbd/6PJLK6dbMl5fDGuji
gSjH5y6SSI8MCM0Oae1VKISrvCnTkV7L5nTaKFULxbEKCKHZUduzfXoHPz/r
fWL5soWDLoKWSJwod+bmO3h0eCouAxbrx0yU93FwqS5zJoHHAzKlnBV8YNm0
VmjfBlAIreFw10FoFcrBFU+U1+qTzltEYFN7ZSoC15CEUrecQiYTD+vjjq2e
2EKGeJJxBJfJEQIJioRdMs7tbjjdtbI68HLXpqQW/P9TSJZ09vN24U6fE5rQ
e/tdDi7pPa66loTGpe8FFSkEs4SHduvG3qKq0O16VZ9Upkps/XI63YRtFqXe
O/jz8Ik7L5l0Csu/tUirROoPBj5m0c9t0poyi4zWZ0R7/nF48HWJHbyYlV7e
H9+tNyw9NnEM1zj/sL066LLDkAGPbALeJXRI6Bfvf0Z66gSK1V7S3r7iM/kY
6Tk/0GFrQLNRSXKLgeQymAXnZdkp5KSjsIc8a1/7qVlaC+8gwVRAJoM3aBdt
fBH0C1aQjL3DoIAXaDXgyB2OqYUF03QjtkFN0aMWxdOXVHts/Xm3HvvAJoQy
vkmR+V3uMjVzDLuDS++FFGu8lUgy8arDDekJmApMX4s8aCXRA3/GTf92NSUH
xTdE8n7XwH0qBu5tjEaj2pvAgTNTVwWXMgIbNNC0xPSpm5uMq8b5ziS8FLVR
qeRjwmmePfnpHAztwAVc30dtNjVgFE7z7SGFwz3Ht9w6GcR5g8VH8ADa45mx
qyTCg6LYKbybYpwHUaBUQKbfTZ0IvIZgwun4JvvLT/M161VPUa482DP34TxA
BtILDOHRpptV0BG8z1ht0ngnXndql40aCwBhUugESuhz5A4qmxa9XmxF74k0
HdaleRCoKPVLdqVATIayj4MDamrm/mf4vf/0BDSLYPNQDZ/Pvoz6s6gNAWGH
+UKSM7I/lfdObbbknjbQKbHNF4FmORlMX3I6XjHeqH00XWnTeQgUWdr4nOOx
2dz0oSTZy0Mp8XDP/NHy2HIppF57TZk2uiQDfcekFJEJaOHtzddcgVjxTd42
SA81ohNh6pZTfdgxGJF4oVs/Jaz6g22NtHKGT8f+58JGhhetLQU0ejEWvzyd
s1AcXMUOTBHVL0d/TsWVTfoA5ONHvgqs1Og64yc8pcGU5F63K7I6wgRhbXq4
tb5oEIzbgBhEcKoEOfOmfpVQDtImULum2WTG43SwRwannWDyqwASacHqsH5F
T6FLc159iu9vCD+fk4P+7/gJdatpR4okNeU8AygN7ud4l+G7+wSOiphbXLM7
YEPAMpnn3Q+rQ2l3OkJX7KGw0IXKaahQ4ELkVfD48ml6wbbQUwtEiQEKvQzj
aCb/2/cMnDjSyKEvuPXej2W/LTQpZHrW+iqiPmXxG7cw9iYTpaw3683lnDbA
/jz4WyoKZUu3pKLxsuAyyE0elsAAIrlXOVgo2LkdcQOYBPOqAdc70rDTh7g0
gVrSFgWnwz/45X/CCma0vniPh/f699DfZjlYBt8YH2QeRp9WjgEunrLsjX21
eXPMYDMnHkzUL4v1JfujeiKqtk1tIK6vKzERHHhta7ZNrX0/60QbxIitSzFm
wzsTatUjnz4JFA6U1OxZol08G1tsyKYM8FDqxn+5vJW8gOQ/13UJh7qZNx3C
0TSFg0fEqnzFb/2+lwOjYwxIxu2L14DqmwJJD2YZuOT6WYtUbBBsrKZbPWI+
zAz+5JDBXNbAqcK9BpJbq2fi1GRrGsa/f+Dssn++Yks4kQl1LmaTfKfs7BPH
XjO+uMru23Xv6SmuoivCbKXV8rlH1QmGXNse6OPXrSBIrIkV2rz9rBUYjUs4
HhZUoYcy941xdUtkj1xDJnwram0u1A5DxuD87BSW0JgBpp6S20oML1hwgyhh
6wV5PcGzYI4B6CezT2fXp9YK1TwekRz57jnzoUcJJkJcC8Dy390uDPlkPIoI
AqMS6vx/kVP3VifOkLjQ4lhRp3WJZHA+6Vc8+yTBhJH+nC4kKJvjS4pCmRM3
hOlFD6i19H8zfa6vJIFB66rntdTBo2Cu/OPXpzKvsAPX74l3N47hz1KqgIKw
UXYDo8VfmG1mNc8285mv8w5wsFZyzHF9SP6lm/5BTXQVXZrtlQl/1+sEwSj/
PE44yOKknhuvQ2sjMpntjKSgYjm7S9p/vDWjmO/vAU4+l8uLO8vg0cXuM8Gs
Rf573wvKOTRYevFnIkBDKahX78DeAOxCyQwxfWdp/JqbfbGDj3om0MrYIvAn
CxzNLLZl7IhuZtZ4c6ZzQJ2K4ceVwvCNGkkK2B4vnWzUbAFILT6xuKAgzBT5
A2Zr3F87cWdUIAf4ghkZm8gvKIq1Ov8JhITyEsO1v2vitS89LTx8tskMiHTx
Lw1FXmHolY4+HXfxtXETy4RjaaPxNOnmzh4a2VDx0055pOn6qp1n5ZGC3yWh
xlDvBFwbFF84RibfLjK/a+u5Z5cCh/K1WYtz6/aYiA6zCzFVZqdrDkzACOgv
ImHH+Bi4oMTsHfpJmMmD8StwSPq/G8aQSs8CmOGUn3DAZI6Q3Zwhk6L+W7cz
9PHT/JpiZr4p1JFQtFrHcFcF4TGwRWswst2CFFcnG39atR/xsYmggism5C6a
U5NGD/qG90W1IWFN0n2Kz0zxNZ7aY0U+zxW/isxNWGwKqhTPs0p7QPNysq9Y
ht7RwzHLI5f4Pvg9tab0SR1pvzxliXEOBb9VENFe6+JzsXn4usf7TJT8FEAH
CS89+TjS9Qnj+dfWH/ZFMxMGV7Qe/DZLmDxmZvynYf5QxPFXvlzxVyyT8mV5
j6ipxBMg73xcCOdN58ffa5PNaKMAE2Iyod6aAqnWHPwjR/w3ImouOO5/bVhF
NA2FxeyUHwQalrhT+a1z6fzagfgk19pMzw2THKdWJh1gGVoES7Ru2NtRZbfW
ezTPEpivh4jeP4BCUE/fHZJgo3V3hTJF/R/8F0pn6jyz/iT+gH7CNT97xYKp
hh2+z4sHnmsxNNYWmPJck8ejzUVKg+q4QZQLisBR+7Mkw9f2Qv1l2zd479+j
9miJZ2NKj40SLFdSOcAD2ZYAivJexV6iHULoyya/zed4b/mi/zPcX7IrjumN
h94A1w5bPBaRTCvbUryBvyL/qLomRNufmTgssIkfyFwsj4pEZu+TzqTh6Pt1
Y2jFy0T/XyO1l+m6XjrY+wI9yR/YPQiSPMckMoeMUB+sY9DET9dKBewliRKR
EcjQCKYtAext3ZADvrjjDJNwkvzIBLvONX9CQxfpbH7c8Ehfk3mL5LJyrK7C
P6D2+AkDpGPeB01SOT7/4HVsoz8PY1GQX6gvevL6sMqPbk+dIMFeAHzV+tpC
XhY+9rcGfIyrZuJpFAhcKFgbZjUuTxuw2/eu4fTA3ltygkrV3zBpnEV6voIX
uWVTAov/jD7ooDuyOOUJwgkiAmEBkfRygEgT/KQivyudO1y08oVb3Wdd/NpS
zT8nINpJ3oQywbp9FQM9r6liJc8lRpuv/K0zT59pcXpq4MEU5EQa0THuF5f2
L17cE23dsPmw0KaRoPWPTe/VToSv9HMpQJBl7rZ43ieqUe2FtPvuhwNvYv9A
Ehone2z1obhniI3VhJaLH5feXqi1/7hanyZfKw3yHCx9SH226KvL0FPAGO1t
wN436fUQ8yX0qE/bxwvrcefTA1rBN4XXgQPOdKzGNohtSVdpugpNi3eYasyY
Zc7UPA91FHd6hMx14hwgbzJvBExtz34eMGpEgrQB0ieYkEQNsxfiZ62ssQ50
AZBUYNHDbk3XTUGznsADIPZ6ptZD0N9aTCHgKn6pGHoB7C/hv3wQT8CSo+R/
QorgcZad/136Xm/g7jkzexyAQYrVP8Ghr4sNseE5q+iFricJ/hCaVy3i6K42
w5Gkir1QjBJFCIw5Y09mE+JVJe+t0l0dYJE+z6lXGPmUcJ590dB1GshR4Vkb
3vti3lwognTG39eLxGYGV5zlELAWMc2VFi90AVHpmXANMdPTPX47YipdJN92
T25OezLu8OZln1weg0Lcmz2BQ2qmTOCiid2BswG69a0bCS2zLc8jPgkCEP8t
zliO+izXwqVrow91lcx12TWccP3Jkao0fiWFzf7XANFBX5G/A6F3zqC/IgU7
IGBFXH9qHdh93Oaz2IiquyINZ48K5r9ttO4hZp0nD14CCqK+t6Fpo5wbUmL0
MYj1nwjBtk7HFpjr+C8JmZgaJHAcrJdJgHY10T1VtgqYCpfau34CAbOQOCdH
DRBznqo6PlIgzHsd5QFRRUTPxkw8QFUidRZ9FWxeko8Aqq8PGnzW53kVtfsC
eSECgVAUrMFrgQwWOKzVJR7ndbIgGit1zm1ZUjh7UBs4NfJStIUgJB88xHv/
7VFONd7tXlU4zvqhkbEvh4h2mP9EHxU8oaSjvaWp82DHIEdXIESa9EmQsY/L
QLp7uf8sMXpiqCBXahbjan6tYtocLLdpiUktKysXVAMdr6y+WzysKZ6ZW3bh
T1K9yCxL5V0puXW9iaRX9AlySJMtXkG0zu9YcyIzxbn5giuuP6zQjQx/8+jg
mPFhgjOwzu3OdH7lAThLtZMWGqumE+j4baCKue8bq4XySwGjlgcutOPjsZiO
6SiPKqqSVz1Egu4pINSE2ZCIzne3mgyU7A0LhxLRGkzFTAlqLetzfi7vMusQ
H3MkIrY0vFhaA7tWFL+CZl2Mlv5775Awmd9YyYGel1w0ybhBl9nLP8i4033W
gJQQL4jmZb4Ar1QNsGL+vSXe6SPZoArtpNjMWEoyMNLOnrVFiLa3zzpBM0ZB
g2Ihamo9mGbNpwGxkieOnAfeayvPhZEhEoiJRFk3TsDl75l7bVoomgILKhzI
XnSvASVOUKl0IwFN+wTZCu1P3YIqoi76k6EyHCE8fUMP7Y8Ef09PQnvkyr3a
tr8XTh0OLsgIc3AJqFiTHwTdQZ1W86rL3OU47uBL1g7W32mvFIGdztrx2dTA
QFq7dT8xI3P7DZD01Baew7LNAcb4GJDCOpYm8Sv+vUgSxte3ZYLe1GevtYs2
wJeUAbYGOIpoPTrsm1660Iy00jBrrZ1A1+9aKoqt3gsWaIbel8CJyKgPiuK0
JnB2oKGtbSz8bE2KaNxVE/1eduyxHmnIisXyCMA/LE1+O+9QjI4eO0ToinRu
T9iOn3cWCh+4UNlunmY9RHBIuU33mxsuvs3yXouj/OVtJxJjhmBbyffVgzZW
2aLjsq+0xGqgzSPRIJUsTV7CAO7kFuYVf/1uZvYzqUQYeJqgcqLy6MX9rsD6
xFo7QT22xi9fDGzC5qk5H6aNpRI9Sd25SggivHN2A92/OSpi72+ykmVY3m2Y
cemdTSohczP9hVEZYf0dwRNgkhijgYiil4kbRWvouF1M5AIWRlvJHEH0JLnZ
qp+HzUe3E3nM++Lm6uqOzXv+nH876AGu1JQ9cJKkhhkb0EY/GNgXPlElcwjV
+eX3B8IOqDhJJ3eF2oUmxDucHdJWMH+XvKFFK071fIMy+0cAv4FtTGzJf6/X
1dD1JjoRFE1fc633bQsaEhJsGgkvIOA3W2QWF6Csm7QoYszD2lz2G2dLiOOn
ijYj+OgmiqhP8RF72VdhIZdDG3jQ9a017AWHxwTrYfy0n6EiLVevrjUIyw1T
d44AijMMSkWUcag5jrXsqhM/PNNihHCulqn9tEXdfD01F/72aGshi9K3yGKC
LQPIgJlAmCHsgPHS9Ju6SwxtaefTIIFQ0IRgM4v+hacZL7b3UDgjLrQO6iPH
t+b1NNiwlZSo43y6W5lnxRtSxszxX59jqIHg/cXj0S/Y8GX0TILd/5R7PNKm
dVOfMJa94NL9JoNgtiXsGsSGobQcbcAdGYWdeUF7HVcV7s+5H0hJhreBhaFq
vZjW+N96fCkRZos7eAi+AJQTvP0IYCgyp6kKW+UrezZZjtHdD5omqOJRnYC6
M94ftOm/ExpRKgoQNgnZ0WaonQHfOmrriJ3Yxdxlfctlo1UfXnXn/ptId8z/
K9rcL3aWr3PCIlQLReaqqabGJmbHcHuurj7lncp54FzzZyh+7AdJ4Tkmet85
jN0EcuOLngmT5O4Bj/BdDDkO5Z5pTm7DbPD+/gtgN71zVV8Cdr3QKBc7Qzgi
P4zzAVSetRFsitSoV3HGYR1BMRXbQcr+ZURWX47jicrH6cQ9fzfP5v0c1v/t
5vs4vqubXSHGUbUWyZ47KL0NOexPXV3XyaSUnvBHK0ovwCz9CPKM+7pL1Xqo
gTUN3xgR2qOxFiQT6jqgl0BWy1+PM3yApMXN5ywT4zRmA54hb8m5T0WBu9DO
KKs+2DDSucJ/Gz0Z6J6aSYODwF9Dugauly/N4cNjMjPkuxwFfDxwD67dtkBK
P8cLHiDyk3wyr0II9Lo2owjtT3Nhi+E1A34qxclFD48UKrTwmhvvRNil4KJe
jL60DqC60ZnKu5EKB1AnfEBmVSDmb+KFr9qD/m+U8DeiO3BCN0llmvH1Ie5E
dngQc2+lqOEoY48KmJM57ecnKdiylutRLAyyEP+c8orTq4ty2LmiZlQub2zv
xnulb20AAn2wU8fwEI/bsAYyY8Kzy0X7AN8aCl5co4qE7gldIQv3XwCXpJWU
G1VxCP0AyUOFuKxISOb7v8+nt34mnhRUPQqb1A47aE4Hy64WH/U7yLhPHZYa
EkhXi78Rr5DQdU2jpE2dNePLCgjQni/H43ZNdnvGQvdQNWAuG/hLN7KSR2Rt
G/4BpgMU+G9bYwyVnGz0j4xGsTZBUZA7/FqoCFQxd2KeKDVd46viCSVDr/oE
Q8YsjPngmUyDNbBD2YPHcM1/GLt1r+nQv3mw9RChLdbLu5NeDD02NkcHDGQ9
PENjMUuA4nm+TvTe/hOeSwba7GCSQ8nKanxf2YgYkY4CfV5xAO/1NPXwNNRz
TdMPaYi0ed/AJnPbI7vPNtZRKqtT1VE3NsZ/FJNUyPeG2ZzKL2oNCLna+LPc
o4RaKfBUh10zbzZqJpEpRPjGufLjiggQo8WEgEOA7vQ/KTe22kgcAk0xBZJ/
eNJ+eL7g1ts+WkX+mLjZpqumwZbTylF04y13SVa8dv878XU8wV3qIzzXJihA
TcZA4ikq+oN6eF9Ye19LjEbCq3NgatnxRMR8lkvRHHkAsjdqSjCrA1zkLRXz
Amw557Vf4C9F55Swg2r6U7gymyGiRg+mCYeDiW+0tlHgHG2xUxEzNRnlGgSg
IEHfGuQfPCl7vk05stbThEIM9JS7BUbKrB8KlCqBZbbrX09bbAfh92RHdf1d
xPXOwBz8/2h8iYeGTKlSTskMtwLZK4+k8u6Qgm4BaZ5uJkSVvEDuBlfg7x0L
ktbHGh/m02Xg0E7clX253e79bFoQ930HZp61Osi1Voa1i1lfdq5jejDz2sRs
HrbhPosmazzv8ZnhtVsXWgSESDvG4p3Bn/bh6r6NKvSyTLhY36TQ3tMtOijQ
vAchHbj0GE/ij4sYR/eRWq0NiOA+ETlifCgwzS0H0UiR+Nw52kfBp+dLLDHd
AN858/jmeR/Qbh8gYKPuJUPys9ue2EvismW28dbCNerYEZ0UV5EA4SWIlrC2
j8TqDDZhahGTqsBxyfyj3/k6Y3cJ22RDIbamZBKfICiWBEcuhNCoDG7FM8CJ
4rgBM/6dr0au9aouyzTfk5SFu3Au+Dg+dfNsPTc+ta+VXvMsLmfQ1teC4Zxv
rpFqAjObtJTeH3RLHXZNuEqlipSWRB9dTaVlH3hKJ2KVCg0rKrlhXamRKlIH
lfCFVu/xT0NoPrRAdVqJXAxxu8mqG1f6kaf1k2xRQMmGf0rwqNiAdZq/etje
5gvOxb1cdoLOuxHkp2tfRrK1z6uf7lnVmJ9IplGtNMof8mFK+iVoZHkoYQZh
vdVDqZtiU8NHUU7Dcu946izloJ2MoayF5EfVoqBMPgXAk3bn7VQhHOVv9znJ
mqYOHht/o98tnxM32VlqTUTkkPCRi3GVopxJIeOhBH4JprfOvs3k2xDbhTAM
8pr8yFeo8NblGbayvZRHcWlZjZq9QOdct9BN6Fu9+ITHg8dMFSFp8Yw76CgV
TDeKLvF45ALS4AeEPr1taOg05VwYJFgfGqFJNkQlzaymVjvJtBXGAoVb5uHw
zxFmkhjdKc7Nb6bCEHa1eu210IWZQmTPwlXJMQ7rliJza0KJ+jj7snuVA7Bh
7oqXAyNKm1BwA884LWxsEuRITwTgL1LVl7PQ7ktV1IWBa6HGXHtj6I8YxzdP
ocCmbB7WOHJhCt09GBvqHqBmb66ZImiKuyRRj02FnOdTU+A9069Z/EsovdQV
73Z+bdCmzJQdA+RhjagvTdudt0ZHypRUjBow0IGRl2fU2S/OQvPWYBAIYAC1
HnyunhUyw2K6/uiIgwIUpy3nTUnwctVK5TOG5zROxMmzBbpcdbCqxIOJgdpo
QWTOsZ/iE5yKkyLkea7sIYWHqt9WeeE0oWp9w9aXPDYy48WzOzMraZJflyPy
VL9ZaeGCLojZdj0vWx9EC4S6z6hC8ou4NgyGReKd97mrvHL/FRbL+KP9ltwf
daQxlDU+VJoWSaPsSAT7AT1/IG4yYzqT4RPNnVY3iMgc3lgbyyNb7N1grNsl
SVKKKOGrI4byIIoAYyyohl3sg6mm82wf4uylksU7Hc5gpqZG9FHX2UuKStxj
qN22X1KzAqRbolWIYMMbv9jZYvGHWrBPU1qcpO1oCoAPiWezKJX8COKNiErd
29B6dwk+xCkq+Ohi20uK9hr8XsrudUAP9xwyqbEPQAy8aNwKj9JsfKCt1Vy6
XMGH0M0RpGm2+mdwOtlwny0nnrEGSwuo3jyH2ajsutGt8x3Dm91GXImnF+0J
+kRu0ewbIc8QXyqvvA7ou0xD7LOxC73Vig7R3fZv1mWGaYZvhCuh1C3E8ROs
ouyKMAu4X8rIDjZ+OXqmu4TY2inbTu9pArA8KxLE473dtyaMIaAh5ntRKsg6
TRqG3qsPLyUTSBZSEbb6NVB5EGyLrXpMnLae5/GtsDVVMvHgRfHMyx1xQoUq
Z3oOg3kRrmmPL+MNdKp4R9jIlUF/qE+rvjPzLEk0mNM5vzCxLOTeL1Wy7ODH
v8bNhpmohsr4Yucq/LWTpqhf7HjIHvRht6mtHF5XKdVB9ptR0YlpPXoeqUoQ
/IRkNJbKf0DJeX6Fu1VWNISXzd1N9ogS3wLiXJ33H6MAbALqC4g8vU7bWF+s
+f5t1sp95BMILsBox2d8AOpeSUATOC16R9iuVNRpUPXisu3LpmWb54is+Oz9
xgRmLB0t6j/OqXzzllwE/Kb1R8+j7XuIciiddxQuXaKneX8cBKTIV/Os3Fee
+MDcDaRNzb4E+MLppCGdMBvanOUB63P5TXluLViQgkqwAVDtDcleOKYrOuPG
8/wr8xgqJdg7MmeQDczNqeSs2z+TubsRhHRsqbzHGtsp7iewNOms6UwJXjeV
7o21kxWGSLe2WqcrZn18XfYsn9Ub3Pcj9ALWOFMpTI4eA79g23Qmi+V+aPqJ
CYqB7t0ospkxdmCQPbhZWYnzukrCjiRgoa2ExoXTtmXLvCWMBw6UqLBlfGGF
EP2XqbnHFPSLx1yYheH6sPkCuTCTR8jwGWQ5lsExsn6PUGOva0DaH/kFUsSI
R6b+cmFCMYARvn5L+mdvy03WBD4B6ng82lj6Ya+xxc+bJB921khKDkSmKrIz
tcR7CSUX1BSjL+YyDoUVqXOnfKIAiHzJtErSrjisi1/3eBI5gXlJxw+rramF
yt9scyVcu8jcucYJv6/P4V4lCx4hOQ1JVqT3Ss/TBzMqkRV3yuaC0YvN8pI5
CncoKTj6Q2wiQF2MrhDu2noKe4QciP5g1Qt75+3RzIq+ZACFt+90F3wKEbKb
BjV6gVb7+0RKk613ghy5UYv7nGAhJOwSMhmz1jdHkl3gVqayuorzrlOu/s5M
1A71B9Vp09CX5suzMS7BAf04jArQkMbMFJj3BdHnkTgd0Kw1Pb9d4bzZgx0G
aF91UTCyCeVaYloTEcKzFMmRQwn0s+FJYJnv5SSL2LyH3ZwIPAuMz+gHOZR9
s8KImLQ1zylzCU5dDOZRGlt4xQTxAi5EIz1XC/TSD7l+9XZpkCJva48CumZr
tL2M7+iUqCOBvdrt41bZPsr/5HscXS0JOA1Z9AVqWnrjIvdGh0n8XPjtnK5S
jn082bDhCrwvCR13r3lGFyTEraP6lwBNbxS+2LdsWh7RD7ENsbChB4JQfByB
y02cszNgzjmluYvkJ8DcFzhqCnbbZZ6FEqz/Ya165uYcFKZSP/DuCc77w2dQ
hEZbnlLtg/K60njIPL1x/yI9FSHtHKIKQpzxwGX59Ovf7bAfcaVB7X0ysMTz
a/HtyLJkhaurqRCK6+KbZzNGjwaU/lJUoXkbBaw9j+r5hG4eWtzG6D+c8Rv7
fObupW31XfKIou0NipFTZXtQS3I2J3gtEBVCwRw6utIGz+s5H927dFSBEwmj
rEycm8ZSHZXoEEFNWcYPI7JSiHy8lJpJAvu8gCmc1E7c6kQH/n2/CMQHebiY
ighEme9sxE3CIp38al9A9IF5XpkPQdCLvgGyCF1X23mIdxrhQmdtIK9sg4wI
Wxmt44Sp7/ybu/S9PWlYXC4DwpJSkqCs38pDsRdK3X0DBlJAlCWkr4B9zI2W
qT+LsrYg8CcARvR2DCHFRv/XnP4u26hTRkLsvGeBhsafx/IFd1g0NostdpFa
0AamidrZj4GSTZnHmof8K9kmScfDLeKWV7P/oXqwtJVMy5INomoZhOO6pQH3
zS2/cIIQHIGp7Nxv5Q8Y9gwzkoBvlL6v01L2BLMZmD0VXKjIJKI8AoTBeq1m
nj4hzA8OU+1tocjQmT6HcgNfAKzW8igwaOqzLrXWP8zVs4vpnPmoPRC7Dsge
Xvy+AWh1wB+ufq1vkzZQi+MPKV5BKAxUe5in8zAuQce9Fr/ueanreOuEoe+M
b2pvuQdt5vrOEggXB8h5hoZwveDzpS/n0A+hllT3YBWVBqWU/qdkqdCIpyeV
pFOMCyDUwnmXa1c/4zS/83WDf5s/uGAVutlYFFuzqd7h93285qsdmutzNqSf
YBTqOhEGhEIvMk2m4fPemr8Ql4fsugOrSsQCx4p8YD+OzC1d//lnne5eNUXG
39WsEH9fWVqkGbImlMf4m3fZVn8qG1vgFoKDWpZB+cGLMhzvsWBPslwD0BLJ
JCynnU59mBe81jVjhIAcpthjkkJX/NMwTkzzOyXri5oP0aSFQGpHLittTBJS
43SCC0lGy5okAxOvb/ROfoOdFnW+e+RqhmHk7RszyNAnGoI2UzMLbfi6DDsv
sp6MF4MwfCKuKg+dCzzrdFKXB7IzKzf4x7IxVflz/2yuDx1jKuG2e+OAzILw
rqwU2sRR9z8/v9KJMRJ5INilaFF3hO7whMPzpbgXlQbf5CpWEUAuOyd8xtoG
mCKJbBA6BolU5JMCYC0LIQd9NU+unIN1MEr/stF8wmxFkxBGX5QC28q1F8vS
Nasc+IhS9quNJY3CVyfsjxxrzV+ZqnSsQD12ISj6W4fAGWlxHTJw2FiWUWdV
dYorXAkrXkoald7XGIW4/EVszo1PtG5wYxAN0NZmRncMY68jaIYqANz60zzl
1Akt6K7elZnTvl15harYRisfh2PUKD1PByQop3p2OMpsl/UjjiDX9KVUxQ09
1SBWumSlli2Kx7PI7J2ZRsdUXAfwNJFvjc/Qwt0iAxsVZZsiCuk1W9kNVbkj
GUmaBFKgfeu2T8QZIXncljXHmljuBFi3q1EY+eoLr5Z6XH4SQ+4v87auIYcw
/YlmLhl+BLmV+/7IANBgNiY2SkvxSgrV5Q3rukS4CAszFYz5MvjCWpeEvjqq
0thIImcP5A7PQIAteuvhgUXqLhQD4tVizGTliDGBHMFLQkXZEDDF/kITjK50
OXK+YhoV+k8j0w0NaFG1tFyJVQAqpYRE2x1dQQi76UavA6h43EONUDI8MQLH
m11EW7B8LnHum0TBBlcLFxMkkxTvX+hJ71hZZX8tBtrJPsj/XDtPWaTzVBq4
DxEl/dQDxqyoT3s6vs8R0KGsQSpzWLm0IbxlzDnTXBeN9I6nVtcBqJ1+s+Rt
uPG4asZoHGiciHVJRxL0LBBnTylSFXKUc2KYPSRjcSKCPciq+z7nrI2biBzc
T6kCfd+3tC3I5dIRfuIuxsNdhUwOhBSTVdXnG81QlgAy5QGUoG0FTuqSMrju
eM92ruRZ/nDk32fSEOFhmyyYuuj6ExK7p9ey6AX7ABp4inD7TCi23ScdAkO4
7CyVBBmeYj4IO+SsI/mSxFsR3ACLe/JsDFavW/Hwhnc3xc5A05BWKxLW2WnW
UhlGqZn38YXitu1bwn/wHelycuisaXhzgYYNydncf2Dlxc+tqnUjSpGSIGJV
puI8avL8+BWeQds0gpW1G719k3QdXEHXVMQS48YArO74aZCAfXhL61goEBrR
JtXHFf910u3OFteoBALSmdR8eG1cf9Nirl3JsDlArPqHY+Te1vUIK93lW0Ma
srFKL6OwBJxqlxU8ETN3dxvusMtBk4l2Xnpw77gC5NlMnaFIT6VXcFfKDeOf
3fJZ6cbnaV6pdEtnDOXzSyoccagc6yHl/7qrv69BZBD4ofSfPD3Vhx5M8AB3
4Dpa07/OBEqyP7h+9u/dOui3wUhCDkdVuNelyRHB5c/IPeoogdGmVJ5JF5sh
zJnnUoBiAtAoYYlHXmaY43sMtKicS6nLhhpjM23HAA0qJEO7CHY7RIhfpyNi
vPhjlug83I2OKI3/nxa/uTgGlvAoXnOjjXrNNHW6lIPTxERxlwdPPANYKd4Z
uJ1YJDwDr7SoQUhAOt/yQTwRadLYdSCSQnYwCKhYAO5Z9M1xgvOnzDOiDu/B
JwE9SXoqgntg9qNJiGNkmiXVyDlEZA/MbRj7lM2GqaLYpBIlm/wTO7TjWv0H
fD7OzimPIhd7mkOjWw+nN6cRHMcS86XLawQkvbajewtz24sl6MQhRbmveaKo
c50fclYbfATydwqPuXk8aytcMCXDoRNt6kPQHDwQElHvlAOrJ/JRbMZOtCbL
73+iNlL1fqnc2xcB5UfCtVz9WWhEO+htG/tZ6G6aP3VeAC80Vp3efA8xKgVZ
GO+JJ4T4w+zExBHV02WIe4zkDzTG7/pDh9WWvfxKzNKGlL5+YadLkF+WH5ty
+DaRQNofWTF8PaJjynbQwFYHxSuafHGi5OCfFyaXLE92mup8a5Aa78kK8v8s
L8yU+3uoo02pWw/msCF5+ci66EWlrtvBunWJ5iTmObnPtbqlkqPk+UPz3hKd
HuX8khJByivQ0rYiEJNYpV/d/Bs7VPhhcBknNAqTLuJC0O36ZLYyCB9PleV/
tVONuw21WcHfT6+CHFR9oM/RIOrjUexOM2e94PIJXmR9kah2k/PTA/SNlcFu
UhZSKdrIRRP77uIJFg01XsHkBQNNZt+n6k0lUqcPVNdy7MdCQ7JN4SMvWH79
CudAeNvcUb1vQx14FtQMGra6F9f2PcLZhlmQDyz1orCIRIWnuB17KYkpxKCA
ywrtErdlEgdyUm15m14jK7Y8ddrDXygbqDlIa8GmIW5/e/NdZUY9vu3JWnya
VzLJosirUvD6FTsJCoxR9eVRYqeIvD+8vDjlX+3lmJXOosEDrZD/I+pazf0R
wobwj9Ad1/N/9FUblpj8RBI/pOazjE0BFtJ9jHgnqDQumtMeQ6iblprMYLrU
0vyyGuucEP9wtrLHnz6fFfPRDdE+4EEkkzbyD1Hj5R3u3cqsPiB98qhRpbBZ
qKeEWjMidho/lLzUZWdY0pCA/kmHbZBB2TuNSe34qNdWVsgnMY3y6jX226SK
zducoNDl5Ps2UtB5zMT0SQwI/uiPvFxZuxnpiei/jL3OGYo6LvHrI5aMaLmf
yCHKNTkjer+jXig0rgUuF36MLjUkKJHxcI5dMx80NrDaUE0QqiGpvLH4sFWu
4/12vJPHtDePLMDNu+AJFkiVl7tQsy9uCjiL8w2DEJjWgr4UA+OLe8okihUJ
MBiIJW4zzidosyXEeMqWs0tPfBbysykBSyX+CsLBcs8lGF653l2YXhwvY7N/
KwEFmk23fWaiOusiQAaSJrbG+9H5m5H/3hi+S6V/fvTtgdg9IfLpVi6UxClK
s5Oj8s25iW1DkOA1WaxZvIP1Q3ztGUcjbLmkFfW2Vx83lzBfYN2kvEcfv6uJ
rTdZH1a5101gIT9fnnFVD6pEAoyQsw8QCacOgcxyFrNI/OWJm3nj0sAsBCmf
YloK/lNUMnfbX6JVgjiiUNuZArE3iuS2n/HGv1dHLNQcusne2FjVYRRE2lKR
q2dBRir0VB6MZGqBdEZZfQcYjo5XdJMCSe1VUMlH6O2QCL2uXiRjWeb17SiA
w9WBwWPrrVQC7QWUqhHxaIrTMu6mFCOWxuhFz4uXoMt/qpKO2TTcEZHpuAlV
9NaAWis0nehJVsBOAfwy3ZMQNWs2h+G0KF7V+7Q93smb+ltwc4EOJgT+m7T8
xmkcQvYN/A2gz4qw3qfHdG0iG7d4gWnKH/xnJVqVPzl1YU23cW9Ar78YgCZ3
vb3UizCaN2TFznMNcam/MrB4RJNX0PkC/EnPEpfzHvb4CD0oJJa5UWI5aznF
aJlDu8U4ZPjw5D0HCwQr30Hvs9OUIpqYnoxIw5zWEK5MvMgs4jsJRHTPBEVq
2kubBOA9L2G6TiKVZAwIzDSz5t7DQVhenE9caOTEcGCV2u6mc4CNbj5FgEtb
iayCQcPyY748R5qMqDMky8fpLdk6Zh2ApBHfEIJ85vuZGha9oHNLUB+1XtQ8
gJe22o1j0ho/EiELJAC1MFnC6ddnRNtfoBI6zLwYFFOe/dPhX2gHiv6Az3vO
Nl0aq5Yqss2ocup0VML4P8WG7ceUKeXp8atgk/kad+92n4b2kkQwxsEfNkpT
KNUGniEDyjfZzh0SPFAWnB2W1hQzGyNrmq2keJ1iqxNoKRP5sEijL9FdPSjd
YoBY/wz704SEBLMde2X2YrNKI3lCDpsv+q/zknQFcL0qm6b9e4PpnfxEVqTz
owlub3jGoMrU/8yQE88u0mMBY1KKZUPe63eUPpyqPRHd/tzbJ3+EqFGBIhNQ
R+u2M37K+ZPqhQLlKbS1UMeuCikBPQRpNUDF1z41NvajjJbWqZ8i/0Re5RDX
XfO5/PxLP3tzTSW9JF8zfQD7A0Ng10DmQtZrq4JywYfKy0tqNjUEVt247tDz
mVGCV4m7uqyCjr7SxDFgYPV1CtsXdssSq2N3H0GRXa/MBrUGy3fgFVNEEBJN
eapSq7/0OkF+hI61JLe29iTvkd01NGKCroCliaDn9U/VoqKQ6okZqSnYHgzs
1Ma6euYHtEhIHS7VydH2120lcKCcURT9WyjzTkDNLbFVmgc5/SlfK6qgU1OS
abnGoaTcFgj0lbVloDvYzGAAapedQqrWkUXWwqV4plmJhjR8ghdJqVW2MJOT
ZpKnhA8wIX9+SOLnPZljz8pIm9GjPKaSyyKpW8FfiwPowWA7BLA2k+XN7vsD
GL3AgLYVxH8pycDiZiHWejlh3tSK0ApbcOLbhQoWB2IHUu3Y3RzqhvqRMP2y
bNmiZePG8mrrpcpl+bVvRdbCSB6UcvzgtozY6tkvr/NV2aJKmaEN4b7dz/g/
1WXMjhkZpTBxvm4W4qtxaBs61pCRqaH9YtulYBj3WF9Pe81F25/7F1MAbuho
M+e11SbXoxy5HVHXSG40hcsuUvI3mAqgW0mYLtff54NZgO1dC9xyumRN6h+N
kXdotT5rnLyzfScZczJbMYBWF6nK/Xec1kJFEcoY3sfaBR3paGBsNwPfMMfj
kZfTjvWJRtmNmEc6JJ+4ZqZ3e7leT44rvoEmzKCjOTdx9uzzZjVmReAocZiY
pmBHQhOqyGbe4k3iAfsdIuIarAzmUgcFGgheaPPberMV3M/JA+XKubc+AwX/
GAgPRD1h8GXAW1Tg/3nzR8JSYjhEnW9RtN/8EZcLADPklRIcWzKmus4ymNqa
PzN+9Uoh5BlDLqReN5vjYwZuh4ZcTXNI85JSRB00OPsmccRqudth69U2ESXZ
RjPSK+5kZ+xKfQJ6xQjn5HyqRN6xXra2g6Urv0M5XChu8L3Ix+k3W2TiKtfz
Q17B87Nle9rX9hKjBJNj0EpHVrJMeM7FVd9Gb0cdIjOZsn5jT3Ne5Jygbvtx
l1Ytlv3pqQcSoBvCX4dF9+CQZs6l2xrPQeF8PRB7JafNPg8uXeynu/ojU6X6
WtKKZ+RmFmr9oDRizwbi0MUcQPML0hXRZFc99/+MdgLoJAKr0BFduf4d5MWE
dFHjd+mA78P57jg9oilcBbefRjAjvwI6uBK3Wk/b38AUpGse1SqVLm8gKMmv
RXsCTqIlCnYpXF57CynTXoyHF1zMv2qwxNzB9P0dYmAB5hvd8SGp+Hlkeweo
nAZNrhB9+DAO482qC9tVfiJDuZDJDYiC38GLzC9LYW12x3EaqbTKvg+slSJo
iKF9qpKXqFqIzPeytWwAx/sX6mSbdmM2AuAD0vTAt37Q5O/hvp4PGSAh+vFM
MMApPKZFf0Fh+q+4PZcW/TUsiuCGbc4zIAIiR9WypKxcPmvpEyk3xgyKaXOR
KzsP6sr9z+fRj9qaDyU97i8ilyG+/yaQ8EOK9rlxWvsAe+7HqfktRIS4oAxW
z/PrYvvPhL/B3NMOP+coo+kZgp7qjbE9nhv3K1ngy7I/9RF6vTdgFZFY0PYW
DgNl6pvFcB1HNTKjHRQ2VXXZoJ5KP1xWvSMn5P4qFIHbgKjvA10Aq0eRNJBs
up13exmkPbVJoiDYdYS+6eOSByG2PJrZKtExw2tm3oB7APHWV4IL2h2q+KM7
gJkF3t1AzMv95MWkh0IAp2on7VyoFkEoaIgPG14hx9iuyuJAF7bHexxPcvEp
pwW52UMH0XrkZ0t6J5I2HU3R3ujZIq9FiNmHNIstr9aLVc9EFHBT8Dkvto7T
a+05ohlj6I5hghBXaZTcpdqIUpknbN7kbAafoFvYovG6Wd+RU1IfyZG2ozun
8LRNKvr1NVL+s4kOyZo588Yz9GBlDifBZHq+aHsR8/zZMic8MtrfG76uJMi3
VWl/HYeBtI59aXQB3q9HlDdjpm+/qBE2xRqR/hCb+zaCrQ8DirYXn+bCewzd
1AjYaouWIr6Kkhqj14bmHLA/lCpagRjvwy1D7aw/VOPZg6weiYxPNL0+AsQ8
5PLfbXNuDVJciP3IPUGmRyInU6lrOCjabwk3wWsy/eInP531P5KZuYBmC7tz
lUvsUHnH+b4H1muI8LQ9UyFYPZk7vP+7YJw42Ilvwic9ebad6XTdQ4r45Fud
uRkjQck/eZqHm+cDZ2FNocXlggarVQYFFUEvnRbbmayAyg3YyphS4YU79IKb
r8eSaE18pNtXld3FQS6X3n1SjjLS6r5CGlAcRBcp4YJa/fzPbHA34ylPlJ2Y
8+vWWNuXdSDgbR3ZqAKyF9mQMyqCb9UpMhjQuGGnMNiSxoN1a3CFmaepRysP
8vsow66+b+w4io0RQUKMoaS9ikA/cO9UK7eus7guRjR/nFFuZ+0ozcdPgaCk
vlhsJhcWKjtyYonUvAoSRMYeFZvTXBdOpP9xLb0vhbQbQFdElGjTIpCaQ93J
LAMM8ReQuJsD6FDSic4+KVJOv6XnQ30N+zsLNz7e/j9H8IWK2WUllcgFmDw3
02oqOYnfIQ4BvGrDFtuMHxiiPYPxGUujY40S2TksuIm3Fi+yS6AntaWo47gn
eUVJ3v7YLel/3T+rti4aChOL3m4HnX56EB1M6F+h9yRIiRMnJA98dUTXMJ1C
WRF/wLaITCku71A5yU4oCcZCikL9oPIwLRQcuy+DYNz/1E3bW75y6K05Z+1E
UdOlP2j6ZvahPGkIwf8zw+ZQ5fVSJHw0AuXvjUMjtKDaiopYF/Aw554qpVg6
mALXvesQ9WFeRMxRkVjj1BoHcVtUPf1nThOMYzTsZlDcHyLH5OKbQvUYunJh
MRDRIT4FSFav2iUd3Il6TaA2kQ/3QxCG4h7+HlTtdaiVaiTvGx7mjJ9bwnk4
me8lZG1fnD3pz/17TFEY3LSRskHALPw4nO56HV9OVOSeeFa3DWZq+wKJ+rGJ
KGJOCbWvzxBFagOHQoPBsdYPga8f1hoxSUfsmFBvPFFEviirw16mJzhDeNtt
BzsdKwgTh+/qm92DLIUn4gC6JhZeWACksKYcgBLM5bsEftt8KYn/BinYkTei
jn8ru259aRuyJ/Zzh9yCFHacL6q11+ww+TxLZzS5DdsnJVEa2AxNCtEIB/d8
G20kN+chfOU+zQ41aCzX3wI92Quow/ku0//Kmg+cIvmf9Xp5i7AAPSGQ3mbH
I1vIL0se1HDH4PKp4XXCPhH6f6CbvQGALvUyVYHYLLX07xwRa3BuG2VUdIux
rTMdFMo6Btpj5qTwzMjWoRRjgwamz63nS9+ZWCMIo66JGo+Dd48lBfOqPCpp
H+lNULkF5QQybshZokwxGb6GZ1ztrbuAvQQn4gBWMMVqdbNQkHCWEmiC4K2x
leGHfdw19KqrH1kAqziMqxs9phP7NsUK82DbPHphIvzdZyk9XZgve8HR++sG
FacqQsBFrTt9WJoOfOFXxdh+VJVDZyMbeszfehFfmoE2wiXaXEAJgUR/j8m2
krE0z/SXr5+QLCckxccYooc9eyqM6kEaMPumnhO6kI9y2sD88tGqlqRbEjHi
+4LHZCJORuc/ZEKqHW9TE/eYe/WfYVX7tbecjBUwtwJd5EQecjDEf8cim4P/
/JtsJXuAhfCtTOPUgUPSPZLDcjvUvocFAkq/UQ3MLdNGQAv2EaCbg/HScl1t
OU82cejxDaUlaqFsLiCagc3OA8HiDO/JLwWVx28Y4HWHnXlSzC/VmK3Gz+6J
MgqXw1ZpxR3tlV7m368SNobOVbvnQmJb44kToDCHU3XS+fbpXy6CWg/P7VM5
VbB++QRcgLq8/+1On7v3E3GQOGvY4RMo/onBcTa/VBkbgKqrEb0YYz/m+MCR
JjHf0jQsS5kqoRxzwETZHyiQJEzzFQN8Z78rsatWlbKgWraUoC33USXQvaoU
T0cJvAPaR3qntPJE+BVsoHh5iOZzbeqnbUJCvPxRduAICCZ+qssXfC7jQmhl
+Ij3wcD3vSMc++oY6/nZ6gyOYrqJd/WA61eJn23w3dRoHizfaCceP3QtgZox
LHFyGglVocwl6kCaC+YxZu99viaFrlnNVT3fINtSTqI6WebQuAF4MYzs2Ald
EM0v9tCiXxP+93vTh+JhovwyGYcsw14AaLcw28BZ9656j2W8MzZzoWja+fUm
iC1vLee9hD0Lt+HSOXRuQoiUJj5RqKzQQDo0VuUT++OijVGWmts88D2KVlO3
7lmb4lDCWy+LNprp2W1qeTCqQZIxEiCd4jogIDMLbFrV9FhogKFhk3Nap8PX
EoTdTcEWI4puO4u8x3VXjzsc031Szd+GBd5UUtpMm0TR/wCCQlL29unr0MZF
R/wZ08151tHQakH6xZs7Yr0gvIU/Rpe3bzGVNBVcHX7kCITsS/SIWjdRYcEv
TuWvuJphIHR5oN8u+CkG5KK9dWUbr7WzmS+YyT60O3JcX4YWiYnEKCCKCDYt
XCOCUE1sVQnOhXbm0f0NLCeGcVsClNhZ3W2ZYEUIA6O9LlYVel71Gc2yKrra
LEZoZ8PpgINpKLioj/KCs21eGWRttA4qPLqAY4rt325+SH9sPGLbYM2fM5QB
9yqMMYTiKw5re64vaU3O/anm65fZcFij8RpqVlRRa/PyzLFQ9R3PaKV7U8jf
ECYLKCKqjYV5mu8iDTnr6g4v+O7Y6FbX19G/HmS0VVvo2cBfqNVMbrXl8XP2
B0J+Lyw/0YEiVX0bofAr+Qylmw/jc76V7ZsLTAKOz2N1Z0KpTz3ZuXDPMNwq
CXXWKMjEEivASNtRicFZBpOqLqp+xh161EtFE5vV+Mo/pxxQ6ilOdSMUvae1
Insjzth9SsBtVrfkbAhrPVt+us9YIRf0esz13Ya3vNc/rm/NR4ZWUV8xQkfP
BnX2Z8+9BOMlDxkTiZY1HCk8Nwa6ambO1OO+YnOMuuGqZ9B1XX9vMrIGg8kB
snA4FcJgm803+MeywYidqrePYMoHml8fMbhoIC2vdEz0Sislw3pM4ofMvWMt
84K2v9iDYd7Fh7McumHk1gypRKTmECIt3O/VswdDENZfjGUiV6LhydBPuBb0
mKX47vCwQooCz0tOT5j6CCa9ENz8u2d52qlHKNBDREAKiDW9yBlujJy5qA3Q
gI+7fSaC8EGfbjMCxwvJEUOB711DRQJEWTbjQk0YjEbP2q17eS1OcvE4ASFY
jvW84M4wUwjGHS/xcCK+WuZwbkfTOgU5t6dGNHfa6qGamlW7tbiM9At76yj7
I3d9p6kvMoTJUl1toRs/ULJNWtX+Fje+ChCzWNaynsjIK/LJhN30YBT4jvDB
u0e/1LUTl2JU9o/LCIfITqWmEABa/GRNiPPiK/zJyfbuHhgUFmfux+Fn5umi
2/tbGX3wChggcLJhsUOlfgo54WKdLNyo62bjKVFa/A2fIa1urAdl9yCQrJmg
G9biC9+WRpOHiyg1U0XNecl2AdiFtytDGUpWfxKXQHuKhbPm3UHgGMrMinwU
ttpq/qWO4rn8SnsrTaT8IIdwH70zcLe+mpbQipQIwpCXdo3qxkEK95g28jDI
tOmYVA3bB07/O7j2Gx93h/Uui75tmHtNYfUubM7DX3jPbzuFU6lf2YYb/0Gn
3B8jSfhdljJVmyHaDGgdfy29+D59WRMtoww/euybZySPcB5mNuGXTpo9+w3U
kfoOKesjTAn1Gl6k/duN07+N+1nQVDnCsCjiT8Rz7N2c5fw60aUS4cxB76e9
+gnLzALtAU9dDw8gCzBuTX3pGi9BRIAvkfItNk4CbPJBQWxYahRAXBNKckVu
tAZkBeqTiRre7ojrPBumHD5gpu3ESReDiS6PidN7geahJmOOjFZy+UIlgeez
6zwEzayQ1cbnw3LHt4HHghKaueXI5WMTMKXqlXB26p6eXGVDS08XeumnTYO8
yRssU3e39IflXj7FVszocMvDEyg8C0JSr7ltHEyBplyFrDZx1Rt/X1rsfObM
3terWV25OZReCDnhYXr/Zyey/EHfJmVzzOclQwXGSJquyHGVC2p9r0ZSzwXV
LYXfN3q46zOvztQzEf80d+c7R37daI+fo2Av6duQkh45Evb9aOIs36CCWXYE
yWB7kHsoZJXlC3M9MTPkgyy9CSnSv+GAxhT5ZXGYvK3zD1LjSE0hWpIsCJyv
VaP70w0duz/DOZhRk5XamUYOfxJSoyTPb52Tiggh+/HSX2BFxlMIs7+C+RPa
fry21UXtR8KA/enyO89+7skwWJey1PZOYsDP62YMubIcSDIRMW/0l1+yiC3X
z6tsv369t7CJCl95qa7bhPW5O90Qq08AzKRcreRDtaLZ6GRx7VOSnYv7YjBn
WZw1s0MeZDT4yk+bK7S8hfexTcOjs8y9R7ArrRT1isqNUz6DAcfmYleYABXE
sTeQ6gHt3xdBZ2sb+vPo1UGOOw1YSxhTiMoABgxd04UFGPp3Rll5UHYrUK/z
QC/HmOeLLZ3eEfDT7yfKNLabA9TdRt6mwPTPIEe4qtEE33zfQS1AlPpR6cIT
jB+H5twROsZFoqwYEggR0qUdiWpUo4pa9V8Ly309gYD2oDnzWHtmnzMikK7h
wzFBX2jE/jJThbeaq+AYgrSJzX54xJiyMp3aveDce07ZGdulesIaTW4nx30L
X3ODVe88H3MNv8dn7XQWmAyuLaNIcBOW6nNA5Ik6DZE/i1GW/ItV9c6goMr0
158FtdsHyWbsSDtIFUmMNJjR9MOJRZTCz1I5c4HgHV2cFCyiemxqqpFoscaR
2Kv3wu6qTmlsG1FL0ojTsfAMyLRvBLrds5jqp9+Zy1q5dQtJlUU/8i0OUQic
a9C4YXzo9bJOe1Biu75PUCLBHaEpjcz/gEBNuShlqUBxe8sqlDSu26wTkN66
e4lWC405Wz/J4lak6E2bhzPAkefcScFFrt0QRSPeHGtdATfraf0z0V6gB9WI
4DHkV6Lg3SLfIXY/qMY5Pa6rwJsGxrK+zW9+CeqqhCLTcOg46X2rxic19nGa
75GON/62nUjOmEcCf9jba7CB4Gifhl7ozNPy+TSJptIWYCkOrzOuRSadndjP
ceGY2CssfppucUGO2mTEAPmzWSWLdYFhFgcO4u89ezodAOy0Dbmq0Av72COX
bgdNWZ56KIHP/1NA4ikD+o4WlP6iqb6jHaWmp81Lc3CvhBvz8rfw+p3G5rRj
N13ns6Jh/mNocOXjQP6+B5/JPtxEzE3K57XxL5K2js8gnH5iA0P+DJAXuQ8Q
c0gM9U3iIRxmXe+f1auPaPEA2lkKi+qBprv+SJTde9kePlXa+T3mhGKrHGDo
PPxSJ+Qiq2pytz/hQUIhqBLLmMmf0zgdF/JgM9iAcf6XN18rdAebBpuKVdb9
BGtuPcEktUVyQ4Yxl35Q2slC8nQfbWbxGJpO3Lt5VL8hCstQ3JY3NQNNVh53
VvqCM4MoHsS99hqMtt5TMpxSOifhH1zWYDtrGh+3pkMXMFOo5LaxR4J6TnCg
/SIGoJt/IwO634aPpufPDJ4L07I6YmCpYNd8NDOmxh9bx8Ojfr3hkgY3JyKI
Zw9VSgHQVEq/y2IF2IJiUllB4wIFBqNA4Q/GxQAFNFRQ8SYvR1xAofFwTE4/
fb8C28f+JrFh6NgzPAOQU+Q1ycEbUUZc7VUlkiigkeFH519+mUccBd7O0iBY
58iwXaTEjwgwo7P5kYJwW5RO+PfLZEKSqCGYErtsa0CWMhu1GU6zJ7u9YR1s
yqAVsRPpWrEoTdjvP8pVXC0hTTVgTLAJ2tzxI1KluofzozioiLnGtRt3m5oV
SLtDCjNGYH6P1b2IcDl4aPXmuHNaafdNeM0rlHGczQAaIMCbg9YdZfkr5ip1
XfwAIUfbXHQ7Xks70gBigyEECZCgPxic/sUn2vCy2j8JIMjxED1A8Grx/EHA
iL9+zJGuaRxYF4glMLvbZXnK3zIG066Li+C24IiyTe7zo17yjF2i2gls8tWL
OFFG/jmgOqxa6Bran7SiNsakai8nFFQ7es5qMAcI7Q4KRY8Gu5fb+aSgzYXn
c5TYnfLSehdrrZHHFDSWuRFp0CPv/xgS/lZbavMnQsxYtNfwjKLaglFTe+9x
1HZpVLH5mWdU49CPM75FaJOrMeycGBb+FoxvJ8a0CoTekG0eiKiXSG/NxRO9
8MZRur+SFrDIiX8LfWKOBA2dxkEsWMECMNelUFFwVWfLbMWxze7tdsDwpvER
8DH0eZAXPEwyiavYpT571t44ccTTd3J8j0RWiJr4jR3qHt9lfcOfFiglMr8i
uz2Ph+GWS7+jzDOa2GTul71xZUWwWoLeWCUllVG1m4afj/tMphzzTdn9JQeH
xS3wpBaozl9nLjnKZkBy2nfZ6dl2GleF8gcZDlNDrhvNZGRZUmNcU4cJGKpm
/XU/ko8hpmGUV88K9Xj9GMY9JR+cGuIHRg//mcUVaCeaZIO/wGaxALCv7+kL
mg7DC0OJgDgY7DMslCUhayvXCcbMH3auPkIjqvN3tcuFuHEsiMOrgkdWi1w/
DjgfTJioptDCjOj0NqMUsTxKQqpNkqkiAqzQ9DCKmKfzdRDRihy3YigVzASe
/jR60ML4aoi4BW6O7XyPlIGZGHm1hmWQzN3tkSm6UxXeZACVGsjudtm+fV7s
SsF3vHC54hj+WtktUZdA3k/o79oKBf6lm8kUdwQXCnRWtFZmluApMqL4K+9I
WvgQ6YIXRX5peXaRkUubH0eDhp9sFoVEwwDj66PHANNzZFPYoJOHuY+4XOBI
TGkUb4bVxpB5qkRoJLQgdpXbtcDiohB6tXcxukEwUdxVDchOsj9DzVcEk6F0
KRpraL3dwKKlF9+qtqexd/6p5DWaEL+qqxx6uYuQk8wE58H1QUUAb3r141Kn
gxZZOBlKxgxINciWBESgTNBPnvJDc7+8mbTW3y0k868X8QWVoTfxd/MoT+Zf
7l1FL6BZa3ftXtwFjzdACYCqSV0WB0yEAqFz3E+UFtZHoc7O69IsM3UU6uhK
kkRgCU/QKsRZEf6yA8bddfxqty6duy2XqG0Q28S6u2dorQn/s2pKObQ4OhFh
eJA2+wbIjXPuA3fZ/cc0PO5uVkQrwKa92yTRArE1dXSCLyhJnRIP/Euwgju3
GANgNI8twLFpuwplpWRLJ3Y57AEu213vknuMXga8lfOyekZtUzvWDTX4WXci
yezuC2b+sD6dTSTFW2JVkGXvF7FXGSTf/SSjLbQGWRDAo2h/O5BxmQScHaoW
ENpdcI8SY2WAyelFTQmcZ9qp2DUDsJ6nV3dtrbpwmTZ1/YiBJTe5wX4GF4jZ
CcAix0w0Q3KDEYkbu0A0v+qeYkBFjZA2uXs4bIYv69fhks8Se/+ja2EU7IuO
oISLS3G/SEVl4IlIvHM9+PXmCghyax0tCoqpAi8dL4j1GHzY6uqC1BeUaZgY
GJjLOUqu4+OXJcbVQfDYrT9JO6cAXlaic5Kgcnb6oyRR99qEwAaw2MbcclxG
R8dmyJ1OjYaoIp1mpHYInaOjzbr9Ly4aDGamZkH0cTcpd6LdrVZQd7t1C/Ov
9ADei7c8qOQn28gfZ4ETSe53Vo34HP1opj/aHIztTF1VVUAbwTSKfW51LJxi
hRtvKGreIZ+FNfpJNn33KrwER5dUv62SvKqQa+MSP7RFoDwbGi9DjR+8R/1E
Daklnf0j5e2D5gfqgznd+fGFOwj3+Bq4KPBKUBZT3+y90ExSP3dt/zFbNITg
pHy5nqAw5ojTzW47rlTTZg9CD2j1C0BFkpWAd64XjDY9SMbf3JN8c5YLlD9z
6jSxN3sro+0ULQomFb0Leljdn5Wl0RDAHqFYZ/uH9Nf7NWH/V/dtwpj7KzXW
6gmkRhqqxSQlZVzk8ZOgRDyqtUmMMTV91PvyhJ3ZwgXO1pt74aqhYPJIlh4B
6N8ngIPBRUpSn5Mq0F5SjX6kxBD92FhNV52hkAEXEhFbzNxgVFstDJSEusLb
a1BD682+v43yzstd1NCox3wnivX1tZmZmFcwfUl9FYg8JEr+qoG/ByiO0rKz
ve0k/HFCI0FcrFhccm+b0lrPOQNZ8InPDGtzUyR6So4VHG1uy+ZGM5qepEz1
PSpZDlX+WHpYMls31ETi6Usj1JEe5BXRqKyAyvWdam+e9qGh3E8wygQWVgYI
uEZPvycF1kRovlxPaNCR7FsTYtmlxIab8esQslaEeHomnJnoV8YwxGYwKhsY
YkLkRUdPLh0YGmGIstZB+3wj2P+WzkwA6Fr065kcw1pogKpSxbQToWk9XSxb
HdKZT1Dsh3ZzHwI5RXkbILF8dfBK4jnQd6JszM64w4J9ICJx2OD4Kk9/YrdU
J1TQqOq1KuIl/PaqF7PJYm6CGJ2b7J74sJ0umlBcfwLXnmgXy6GOY/wXMN0a
FCSUOWmlhxHtxgywXKjLaoAxy/APtgyeRUWp543WR8l9ZQTNBEnATaDKiFM2
HAD0BIvdHkfc6TJzd0pkB+1RSeKv0G16tD3xL82zX/rCTg+W7xcjw1du7fgn
E9QDTWTxe1iMyj7bMTjMBciluNYmbBvXJ9UY/gZPASBWmth7GSiC5d7g7DBI
WHLhzQJAcbR5U/61JqBfmEMF9tLmOSJM0QBPI5NwJYEJhdKPRF6cXq9HyrNZ
gfWX3GMifs6ms3j7MvexwsXDD6pIbRYHpzWw+fztnHUwJanOWkjPrQIn6qb6
V22OXFvE28nEgR/C6PwKz4wl92QykhesC4AEejeFUlNtGD6xhHapqRoCF3EV
lTcWxV0gBYh3RC2oKVeY/NEl6rhEbgNex8USr0jFIcqKtnf0MH2gkk9Pi2xG
rEraE2ESIdPjHacWJPhHqE36XnghHKfLnoBh69hG3OHxKCYV1Q/P3U5vywTq
sbdqOfTkyrhA0a8njaTozqDWAwyKBrTDN385Y93ykCGqN1ck8WZ1gSB9yLIS
+Fi2OLcPt2e5V9pXpH7mja06yK3Kupn9PfHEv1P06/XEeDbpvRL82FbpGDwR
WZgRSsVtWcbC7wtJ/w0DdHnIaq7IBDtAoJ5kNfTgQIdQd/XZHdcHLXN5+m97
TLBnAm6UVnpshBbrenx3/ereLyC2vfs/KEd5di2kSslA9zdq7BfSqYdvrqq3
r1lXVXgQHd3gn+73N4SbDei8YlTMHIpvHLvH20+lD80Vy02s/IPmXcQWTm+S
ksrQYIjHxyGOLAF3Ebi/H4U/RjLk2ePfc8O/V0luZsli33Nk/1Q7q2lDNdHS
MN1OfTljZKFDftiqfVd4n4lX+RbweX+dYtxOIjFbHiolUDJfC8Fi3mfOyOlH
jB4R4KddunAmwNUtQynat9GsQ9xF/hXwzMKQPbiPQfxVokWm19NCSEFzr2tM
vNWi7hrBtYcgRf2Jc224g3fRVl9mxLnnEeOuHvC+1j0kPWAzC8GEP2ZQRTvi
aUA+al6UrKZqhvdsk3QqQbawpp6wSb0CwBsVvwQ1RRiSvrsMZfyIj5z/iLLI
9mVf8eEkby3DrWvgis8c3OZ+OzhSoXMdcImQRpQhv8Q8QddhMI0DDBqBYct0
oaVA9xERswblidnmaFoBZXhe6VN4+dTcAYaBhLV2Kh4kTtziyr46WSNhJ+dJ
9qVhK72GNruhddhJabSmJ8g15XveJdQeNNXjR6eQu0QMlh5bGzEyUowAGRD/
cDtLzEPcNzFajyw/T6wXVP5p3EDBQK+MonXde9RjMb7o/7a3sHPzLafZMJ+A
mUkqt9nrkYhn2SuUDbuYb1bIFCAe0y0ioyrMPHrXCWMu35kcvq7d3dC3dyNv
cKSZIrttixQAOoXxyLf25fKCzwDNTKFGU7Vi/MG7uoPmpncrw+HQkraAQSPk
pA0jZOEHCoqFcCdLLw9kKKhj7YDrJ44r49c7F54fgEkbML8vTL8U2vKYNaBQ
ovnzjyZ3UhLNNGThEd9cb6xMUp+sA3FjXkHDIqyGx3ZAk/DiOwPcdcUp4B0A
M2oEwlrJqcG0NHfbsSqWONgehvNeOSlVqRn3s8fEwcrCJruNlpL5jI1YaxU5
IzIVdfAwfnXiGBanrMhgrVBi8NA2VNDb6631e0Pde4ho5aa5VabcfuK/M27B
aqaJc2gGKn49iUo4E6Kxz6tzrIsYMmCmRmwjY00jYSbZTuBzFoQqO7aHgPxH
P3Az4w8FmvjDd79uv65JwruOInDMh+JAkRB12QzMc5S/aS0s3TUv07N7xHqz
CEBW4mFLoiDkuXbP0EdC6EiRMN8LciGHE3d4ZTqR4MRWlabF6RkMXrYHSxol
rLldbiMjzWaPv1AUk/C5VbJzioNZml5mQ1558jzm2AvHg2yl3wfkx5PPJGHe
3nDZKlGPg1zoZrLWXOpxMsMOLh9Q+m9vv3Kv4IVtyGmeAM7Kl4LwijcngFsg
rvWhrTHzFp1x47J6+a+BI61HxiQyvus7gSRvQkDRoaD8vkg2/ka+LiOlS6Xy
0RjmLY0nwj4C09oYOMKwvjTl/4cNVhXnWBae6UtrPr3A+B18cRfWj8/loexA
+VnnWxh3atf+xxzSSqh/hue5EqCFFqyT4Chfc3juTKRWwEFcg7DaYWBe8vgj
pZSMCjP7HQ2gxNPvCUPR9nXPLd5QxSRJ3BnsC9jNogJwOAlwG8zgREbpzzIW
LAtNvE52B6eFAk2wlItH9zxXObLC0D6e/CMZ2qkVQrlkbA2Pegn/dEwtsF1S
+oY2GLRm81C3UDD4l9GWt/7u7sYy6FAHbP9lRf+Is7OiFovpFvD4/SULkvuF
ppuMtOnN8VbnguLo2Hgb7AT4KSlAoexqQcGD2piBaoqWBusLbHMdDKoBcAhY
cobWGQ5BNFANl5MeR6Y3LWskgYDy/1OMl0nWeGdMx4l/A1j+V9pa8x77t99/
sge2LThZqHbGLYnGbEj/w1k0h/zOiGwsEG5niHn4y8tHgyoEMBxqxyubO3Ed
Ufm2ChYX3z2jKT1KIORvDm9EXiMJsujOqj/TYB7SsNdZSEhLFTeY15+8dAcS
k8QOwR2E2MO6WfcJSVmZvXGk3UMSPjx+MGL6QbOm4k7myg7v1EHhhAwE9ebc
XbZf/hix5sijngiy8pMA2SVuSMm6HqdpxyBN+0Z0C2AoKVnX3L1ZOT8pAV6M
Qa/KEAwqjCMblPLYITMZrAUr6RccCeix4URB7wDNcE6veRvyzvCs6zlGYKmu
RFjE0Ti5+8XV29SE1oAb2NPq62jA9OjkzyQg1hPx9gkhNkrR5hqAfel/ge3I
JBb/WKq1zlCqkuyE8dSxGWFQ1R/PeX0GKIZSQx5lSeUouMMNmYnfBADWtx8a
t0eQdo16GIHdCOwrZNqU7MwF4sHRViYdQSFaN90S/SzGdNUrhCBcZOyt/nWG
rHJKhHEr2uIOihvDzvq2xl25DOrPilhQ+b04FoQ3e98xXggKzKVOjQWbn2En
vI5Uf9OUmTPRc8lRQXuMTC6snHC2C2JBe0UsKpkdqVU7ZoY6x74BnEixqT6D
vXQm9KOIPydNlGAmBDbqfwjzBaZtNUIIMWfIscLms7QvS73QwS9mUD/kwYP5
GSg8S3PIr+sDNJYO3c2PppOVWYLpcW52/QyEGDHCbWrE5vKLrcz2Wp4ULt1i
AlzIQPLfD3o3Hjs+Hrqqy9a1gnNuyA8A66T7bDGKWqGT9Y83tw0ykj2SdoUa
ZtsPH7+AyY2lHj0getMH3J9LFcduCB+tXbOcvlA3RmkcmGzKAhRgAV0+si1a
B+/b8OlKlvVXKePZj3C2E38aNCPUvOnzsU0WM43J/DLxSYM9lTJPhuVfe1aG
pQU2vNWfk2rS0vNH7xnIi/1/c1fCMd/PkSwMpVUrqNThnMnb7wlIh+JgxW5g
hi2LODKcgYACvuc6CvILI+dni1mIRxxAz1VhUSaiuopk0LMy1Ty1SGU32mlm
d/jlCtjuWs+3IlA8ulQwIr3eoXpEMgHeaMSQ8DMZfa8fJdtCEvLP7cs7KW2X
g2NHuk16eQk8nkbUbM+oHM52bbLfHx+DOGKhwvfVzERB24KZ29ekC9KbN5jv
u7UvABnZP9eoeKQrrxYtbv7oMhWimdDJy8h87TGSI7sIQWoMV4zID1bhZjTw
9QCcs2rIxT0TwXvKIS6DJGBpBfd9c3yvrQtEspAjSDe7j0/JDIiQT2okc6hm
ujiUmH5NwObjISOQHrp9M1bn909GD0N415xIxDaDJ8SBEYN76YOe5hfYZ183
pGYX0P56/AiblBTqzs055FanEp2KlCwR/ByzyFNSIWSZbIoHSWhftcyD20XY
6t8WUnupz5lJvuHRPC/2RCFu2a4rCSPZSofagppgNBkBrvrn9auupZQoXduG
HTxASmiPXkKFxp6l2V4mYxeyT66+wkRQUQHOmzw3y5D2xT8SCjwGBX78sUFr
GqnBOYIlgsgOv720H/YccxQquDa8Z9xsEGoPN7NIlGqK0ko96E4tjHXLm+bu
pepuzq/Q9KkC310u8IWXbab69KxNRhJoiDsG/8JK+Vil6udSUjErN+4vB8U9
DwbEh64p/8bXR3nc8xgSrOmN+cHQ9nfzIlGJQ//xmNGVvUYvd2pNeuLnzKGt
x24Iyi795GQQxlPd8QWeQMCyUokpZNb/ug1Y5OppP0omZlHFZJto+zBqrcoJ
9vF7F7tl1h0iAhJGw9wejH0AACnv2bgQnjxs2M1ZS8I35yuaIeuKgcTFwHnB
B3bWbpZ+BlblhP2e4MWA4CCh+vbyljdQkyZUH20aYJMTzLw0UHRJQrQ7W49n
GsvDfp5HkKXV1RWbzb66zk8/L4Or0I00oYcTyxaWqTjYlPZZb0S6vdlG/bFm
Z7qaTpdJaiXX3OncINyf996L3qNqe9/78w6laduHh7+Zf14C0hBDc043RxUj
2NohpIX4rbqpxpRfi0n6OHNTST8ChAhFJpg13AxPvpHP571USdIWF6priOEN
+t+Le16jnwjMQtQhwMZfpj6i1lm0+LArMCg7JMaGmh3jH6GNV3k0UZEanr7y
SZqHtNnpjIleIimKG6I21CQGunQ6rU0xdovT0ThzZqk79hv6qCNHB44Lxt7n
E0Op7aPLAcONL1+XmUK2icBmCXbCg4pKUGvbjVLwZk0yHRzIDhg4NB2KkV7j
CxU9aISnEktQyKcqY4OG9yBRKJWZJx62Lcyyl5VQ1rhPBQBD1GmVvjVd8C8d
L032AijqFQ+8qy5XdCCMJE85KmhxZRopt3cX+HJruIIjWWzIjEL6fBnfENqp
0vzG9SArJuYqgYcgtGjhkUz953T4ED9y4uhMgchh0bzFRuMNeY9HwUqVzWYh
1TRZ7iYyFJyg6LI4sEs2/bfmB7OhPRrOy1yIvydXgBNhE1uUIULpDWyR8Ii+
uEm4nsdQWDpTLaX7PS/7cTPjJGJmSteokI89ufd7kZXI1vAi/5q6LiJLIe7D
qHitpN2I5xy1475l0eCxBDPYGmFkDNABMahmL804I4S6exhfI8mMn8m0giX8
gfoTwkcMS275wScjF9Dl7crgmYdwnQwYLIRHnD7Cvl4vBb/+/yOURg/xI8V1
BRNNvNVUEkDlu05JdQtaH4oBIn9foCM8JJBbn+K/b49hunZY+B4c+QPNfRQL
C7yOBUNtxr5DvJdhimsXUZlWAiwDnpwJHN0hCvKKm0hvdl5cUFhFkiHDb0JY
S5UwpJsUDbmoOtuqN99uIBtvOwy62/pFsapR/HSN6yH6IyjtK/h4lD24Rtdl
n/qPBMIv6pM5XPvpLAiYqq3QjEhJ6EUKdWo5+OmcXYHiuBMW7e441beOLS3c
/e4nM7xXOaJohY9OeG86N7dblgLm6YwOLSyL15qJiwV+SZABdiQA/FW46Wy3
kW1hvPptaVitZ+9YeerbV71uSuJ0s27ATPu+YdmEsbUVLaaquVg5fKPnQ3s1
s+lNC9F1zV9+e9eewj2S204kUWTcVrtO2T50b16aBchY5x4FtL7Q3MJ+LLb2
4/kUx6ldykKqbnIzMGhewLugZWoE1voEFc+Y7/mqcAg+jAsqJnchoRaKKHeE
nuoSykBOTIzBQjyAWikP6bRAA+Fb2ds+xJxTieQQrsAmbaFyelICqbAsaxTw
HN40l9mmPYBy+UmfnsHQj8tAu9rn2MBwc17XP3hIkXLaJ9vk4IyViKYgqgpU
OIk58T9H0alwkZUpjcT1eE7p4tCQqGBse1HJSWXczhlkzDIf5Is+NY0b83fD
Q3h8XBmISZgp+Lya6FRRPH3gDywTEHC7wCnEPA802EnSnScJWg69I+xZ5pPp
3EO5W1n1vE0faoR0yguz7u8IMLvhlYR0H04LVd6Ye+A/xPKM0A3iuW08IYFp
88JJ3CUgWDznQqTaXqU07QZfqOi1G6CGSN465n9+PnUWkQNa9I9N34WizRtf
TE/U1tdCvgb3O0fexWnN4LRvtvvsZweVuk+sBYo+stcVPxCxUu5m36tSc+dT
J912NDzB5ab7V9paopOtBIQAHWhHgvLI3m62ENXjg+DJEP1NH2WGi0x7fjo1
oMBi39RMgqJqGZZCvTOf7MWOVI2VIL1LKPil4VZziwkmzaoUtlGviLPe95UV
NTlfS8Ch+uRe/mrrz63gHpBIMVZf9o9G1Ni6Y7hbUKYUWBrNS1JstxplI+bV
VyX5se6fOBQYv1+zCQXwbivo1H8QVkJ72+g6HDcl2ZlqPAkH742jjQD3zPqk
h/nyeTQdLsDmuuXj9GkObXihx8J8529AqdH6u982aVg1mp9l1IBrSeUJJrd/
lKJqmK+/fQckezPXTuU0XJ98w1ESeSHWriQJF09u07MRMX5w9qJ+DhKLo75C
u1bCjgNoyVM3qdGFHz1ZPAU6hKhOF8J3Qa4BzHcueneu0zY2fzzNZ5+vnuc8
vCiMqbQxPiqV8nemti3d/0/qtmNiOIqeaIEKqV7UYDv90GqYKWPMMXlDy1nt
VybT1mEREDtR4xj8g9wzgKo62JokNJGTsnpRdWs2yQ3fXhBaFnyWQFbc3jjL
zKPphpc1pM/FEubEYlCRL3oqJH2a0C70z+sxr6E0BIqf64AMNhSNrDA5SbJi
Ob9+qUe1NX3HlBjlcrdw2vXSX9IdFzeZ17aRrBReSV9TDbnUM0vwebFetKEx
1+29Rui6xNCL2UUh7tksixUQVONM1QQ/+cHrFngmHS3IoACE40IyWh+08xtN
PMafA2Ltzd4zZRlznLG83Z5C4+0HdAfItNy0jmb/gGDeuvKLyK+g3vK5FxN4
EXv/qPir1josKtDQ+emUXr/j56CtIpC1ckKJYNfg6VWCE2INQ8floWHfCf2J
nsv5Q2fY9AqRIP395gP9pl6dptv2hhRT2gi9XuOQwZdq1R9szORMdW+mFqG3
CFr8Sg8WPCevyayYFojt+aDE9hr3wzRYunfejOM3Sr+Y/+Wt/NdpSAXxOERA
FfTIDdXcHCZfZl7TjW1coG3xX6S/XzTuGBe5ikgQb6Z9OjZMiMdtNch5wULT
QHpgaWzfxaRUX7C4lGq0sZwUaB/3qasOdX+8DId1rkd2rl7SOuA7OARj6jX7
6hRc0c4pAf+oUob7vtYBXyGE+OIojp6aEz1fWlRNx9U726fzW4r3NikttNEy
Y+YJrunMY3eq0b6ej5Jjkhwn5hNWTyILpkBUi0/9MS0j003e0XwrbqY92oy9
8I2BVfuLLCuLR5fzwqkO+WjulfQRH19wXSNZ1JwC3vvxvAPIAoE23MRpiRvp
sx0fkldFQx9YQj+Reh7umlexGxPlEftw68LcbFXtgcDewtV1V//rYjuGOj2x
O2BqWlJ+/l4zbegLTcioBmRU0+vY5gosRMOXQOCW/WvbzyLRHx/6farhjqxb
bnHOHXcPYghnurUKRTLajQPln80BxwQLqSG8oq5CW3/GqFyX+mj3mC4QtU5A
oKd/72aIrIYDDDITmNbqUM11PjBvnYUy8VAbcjfYjTkij7kBPuNHfGK4u84X
bM60oxPn8U6JUYcZvzz5SJaMrw22Nr3l9DG3BJ+h1bkw2l75Wad8XRYBiUEW
N2zgIOqAQfMgdL/4rj0yyIgWSZZYi3TJt9LC3EoLp9yypuDZdl7V5+MOni2k
Q/euOO9RtSieQXLm5UskHnUsBeKGfDqa6RNVoGGDka1HG8gfN+gq3QMy0884
dcF6hJ/ddNUC27TMlKlaIbjqVUDzcy3NxGbgH1Rji742TTuvoJykHoUNoIeB
7FnvrNeJ+aOPiukfWBqxQIkoycXDiU6GfHyXizICfmttnHInPvpQ/jxOo7Fk
hxPs/Fj+Ea9Q2tOYbpPPT1fCjkJszfgZdkAF1Oht1UFoOGevThLpGprSWjlo
egCKW2LS/jydk7che7vky2vAntJroYK1CP+1deY7+/qzlUB0yrrWtXtAuJTo
imDYgVn7AF6gVPbLa6c159WbQDOkpErCNTYjFMJonxoN2Io0gML7Yd9QDNDh
nSxWPNjAi2NMS1FAustCBHdvWokop/Oo1Sqc6Uj0pFgfmEwlDbOZyqJGtjHZ
SovPFo7a7pJ8inBGbcay8EOV5dohsTXFC7SypremfVJp5mjYqkXrg0jzq5D3
iHFuTXY8loHLpFFX4RkhWoR47jqRz3QocwGW8t8+MXBEPDKH3zBZvxTYeAkJ
XV1pmGfpFGikjFqOtVtBDoS2xVRAxbLLGmaNLoOMK31qxXG7GOA6EGEHEOx2
ZPLC4uI6Ua7ry5GlFMZvvkOMpi+AZGJ6Qhlpq0vhi95zCKWr8q2tNi4Z5GjQ
HIa03NUjOtC9QmrUsS2IH3iiJNhH2ftUwMFBHhtPod1URLHu1aJo7paCRo0a
SRSjFK4PbkPtjHFpfQCCrPpm1tXetOhMuOi65/zbuEddDB7GNJ5A7BAsM8mB
sIbX4pbtBJcgBj32loOd07T4bIWWr0rRN8j9CrpUEWXZ9w7MM046YxpPRvmL
qhnxWtwdWWlObmxpGH+dpvO3JXKwJnQjtrQvj/xqOINTcPevT2Uco9D3gt51
jSaHYFYEVwnluN2/PY3VZi2rPLIK2hkyB4vfy4+XImwChQyNkB7AXsn1GDxc
q0spoga19rIq0YoFJl3EEXLTTRVK0RnsoequwgQcY0TwOlv4YKetMOPUyMsJ
cjbwKxH8J5p7hkZa0BAn+e/vYSgVybO9Cl+5SsJOM5KipTlavnQnJb7hVAD7
GbRWMUAls1NJLpb/JfoK/P64BK23wOjqc8AHdJ6HnoR0MmRm7Lfy9mZOCA5U
gTHpz5zzw0A5O3Eu5ZbMWFl+3hc6tuUdt3sIbli6ToqVu4J0htR1CUYfp4uR
NUwsOZ+tEDlgEZa+mNpj1BUm/3MhCw40Y8kSYWhadCD7wbh2TH0K1cj+fk0I
qPynQ5rV/m7nce+IuPDwkRe7jj4v0rocO54dsyzMXejFKa/vUPP45ZK5+qqE
bIfZYrofvNGyvie+4/Hp4VHcHUaeSdXDTF1TVgCjNdk9Lugm/W61xSxCebaZ
+mRhh+v+MnpucJOQ3Fer8zhzS2u+/vlKapzw2FQdw26VxQo7X+Uts1mppTFo
mo3OTlLh3IMI30yJeFDvlx6WuOORtQp/NfUNm/znQvVaHKlB/nRGikR7gqFr
Y1KC5uwF4ZfqYo/HhGMSrZ2NVk3L4jyuNlX6XFljKMqodgoLSzhpYzY7TAU6
Yj2U+iYAJSL1Dz2NvaoQLqhRpwjFn+/NC7ewn0+QGE4Eft9brG8V4rLl5Rd7
PYPyPimt5mNKiqCrhNy8jaF+RzXVC8ediKfgyW9rJh3/WBolXm3kI1OEtVs2
k6hQ7rKUdMg9UieMLuAvgxVzsmKP21raUbbBLprte9frxuWG+JvqX6yG74Ok
dCJd4hn3jyLNFu9Z7BwToH2cEVZ5wzH8faB73WgtdzM7urV40kXlXQtp48Wv
mdAvXl96Kq+bMiD0t4YpLo7f9xpqOYRoewlP5LM5CUdiRq+lFZ507S82mLWn
7Bi/my/2eyM071u78gNNsrsWIHCCCL/vSmCwoWebUfUNi1gkUNqXW6jCAfLy
lN+gE7xbiDU8dEEbJ9N7QPYO8lXWvW/OG4tyqj0mOTNUohZ7rGBiGROKj73R
GrUGW11uFArNokFpHB7qussTFC7BbGeCy8auXwwry6uvsbT0X4J5LWBVgjL/
u4RiWGjbIPNQnH+cvlj95aXr2/Y2sEWN//qZmBJi6XJJh2hn0Gc6CCh6C7K5
4YaMXdA3XxGxNENcixg9snS39DfsXUm6wUnLFmaaR/ov43GowZaZaMeJLD89
Jj9PBD4ZFw6MvTpbHW5oB+ngiUtx6MqSOyqLZWMrMsuO9rZQNDACaoZ5bCMq
z3SO/igp4TUhy83RI9y02+qG2G31e7S1HbBuHX6YrA4P07337lZCjm7Nnac0
CUTBZKS607Tsm/vPJb1rg/TV++GQaMzfKGwsJ5JJRHUhJl7MCrt6IEpsT2eI
EioPL9OaoLvXRysb6sXKVU/POh0WXOIukOMcR2D4cmS0qZh7BI7EY+KaxxhV
pFvILsNXuvCbPQ60FHe23ylEiyLnHW1QlTdb7RywktWO0Kp8cKKHvkK6Piju
T/LvF3qcGGgUJcVwoQBPvOEqHyadvsWuIOpcrRo7m4Zm9QMs+uLN63mUDVYk
QRYfhrBretCBZEFzGgVu4soc/fT/o9G4JrtEVir9Xh+WubAe2xUEKH73SKhD
Nvdcco0o7RJTkUGwtPsQKgdFAArHltWqeRngy6M++hwd6CIGNAoOOoNCjVZP
IMSl6sLcBlIoubLjLZpCXGeIBcD2gznlydCLWMw2F4tWQ6SUz4fFl40JMP9Q
uh0FndaSKm7vuWSUUpxXNq9F3pBmkmwo1r7tnMSI8ZBsAZ5vOzHDZCu4qBy2
OzVJIvqO3a/RHWiZVIbsbnzzarvoB7m6CFYObN2/IxoAV6xLMjWxyP/KdK8t
L07Wl1Ta+6n6AmVGf0+tfDVAEfiAbMZnzoLeik7QaVJdoegzCupg9GTRkrSt
q3yzqNsW8WvfacmUWVASTuZ+0ih2hdolOUaxDld1POEnjn1DoMIuR4zkyuRk
pbsO1/FIxRg0sLU00bOJoyrDEJwSNMmpssNWx8O/vR4rMXCmyS7A1q3pR4yR
lbTsZWs19xQHeU9Mx860n5eytlpU8XvQ0wS5LNt99U10tRO7qCN2mDDFCAYm
A4m4GYWaBMBtupqyhH9oG9+uVegVbYs7E8opqI6Z8UfcrGQ3VfjA+oJydrFu
CnlyvLX16lqFhc6GakzTJ7u2OU1AvCch5BPeurN87YRjG7VSaIqfJNqOvhGD
8d5Q6FyzVCKRv5RQEGqFJHHKIG2xOXz4M5h7k/+lkJU3PJSpCN/9Y1FPI/tE
kNXjmE8Iy4+2IvYbdS0T1G3SJX/x+flx9PNocMK9webhhKSEdESP6Ts6MjjQ
5jlHqYP+g10+vVu0vJjJ8RjTUVJC4D10yxQKUFjdFctzwGjCZyXfXhTO6k64
Ihrj+MJCMgqzhxR42wfQJfwsHBsDwD30qtaK3d4eW6zVwwSCgMIqwgk4/pdK
IrDQDPRNOtvWY8nY92DHnx+x9uaYCnO3grSprsK7TtW+S3geoRqEtiTkZ7CN
VucyEJXfcwwkiqoPhmTUmwtj4qaaxIfMyOKFbpgZSMyaDKn/bzX2ojv99RnI
E5UukahwG03SsEMcS2VNEhlS4liYf2WNBqJ9lp/ztqX3JVNsDiMdGK2ds9UY
CnBaCybyzXMv7gYW3oBLJeY8OFMiUaXlZheeE5sMtKNUcHZ2T8MqpwbatYjC
DNXgUsKJLokl0ScldzOarkq07GXtHnX6+ZvX3Ohvfp2A1vsp7IhQZ1qUqx5/
lRwoQmG+GaGT1JqBX6mp43JUfGq937GXQtw5DgzX5LqAaC75rhFad4mS7N/W
L9yU+UcxpYihiEdOAGcid1sDQ/xdFoVZRsHTueO0/6Jy2ftFA/FdiR3p8Y28
CZkelm7In7OSPVevN8YsqSNshIpLGq2t7vs38ZrT0MLcJpCE9Ntnh+BfB4T3
TyQXRmktaWTvmhg/AEqrP1R7X7gXCDUBImrisDmnoTcqZEFUtcHuJDa6r0k7
7rkysklG5mls8PUdXPScaNlIbLh0hLjTpLdNEE/wYSNryk2O+gr5N6NkYZDP
ACgTXTHcLDTX46ELL84loFRvpubk/XEHqJHbbVsn0AJudyIuPGrgjSMEGfDU
QWMjVKhaX9cnV34/Q+aJE8zTM4j6IlWl2nmoEOxUNhlDv7tMFh68Zche5zRo
fcUf4yOO7jKaJuTnytrbzyi9Um+I32UkH/cnnVKtz2ElJfFptE++Mze++2Jg
J4WhKS2P4P+/Qp09i7YsZSCFMQ6RVAptKONrDJUqtvUkXtoL61uO3w4GIH6K
IKpI49eTok9i8rPBaHhZdrmlbKvh5uNYacnQv7yTbkxE0BVexVs2sPYmoIQs
Si6fYUpGM+HagBzpky3WZbVaQLutQ69SrIwKXYYRflqKfetY/srP9Dt8SmL1
AzB3/5r6JTakBJc3KCisLevZMk2r9Ogcan3QF0hTKm0QGOlrnEfo+ijV4KmD
h6lrkhRpFrsrgoUKwpMx4qJjcvCfmzWzXlUv4YcUXHhW3MmBfPI6ePxYja1P
CYEkX01qAhSqbf1UU/4djop8bKxCRjWQnFh1ELYcuEyEGcw2oEF+Pfek2vvP
NZWyczsU1qnLMJRpFvbA7U7t+CjkLW+AcLRCYPO+7wGEiEDbP//jYMI0Jg0L
DbcC1oDgTb7IcvDJNCIJ6jEPj00awveYI1H2CfN1o5L8AJi683esDMfqF8K1
VLxNZ4g/3CmuOFnTKBNSpoflVlimJy+MZxW3geoegO2OumLgC6i2XHb1dXgN
Nepa8U9TxKtepNj2nBxZknXMSKxwWv16CyeNLUulgcT/MhuJr+9QlmWAz0mK
O06szxrylD+p0KP7hbxAlTAEkZUMiLf6zIhQJ/E94Jd8Ls+nQLZd0spgkDbr
zhONJkF1wC7YsA5M6wujcvgXG9bx658rTuiVw8tt20qrdrWJdt4y6iQD28Gj
CIetSVqY73vBt/X6D3NoSAYglXresxPhfxF/EfabYTFfAg9QFguL/VFeAWZT
Tqu7rH9d5k9j2CdLElm+r+ZwpHqmb4QxwPnlNr2LlmbLHH4PWuIJKMAUqyoi
JntJfpC8Ku6xsNS22wgdtDnHBsjSgUIN8Tr2CJFkY0tlpk07Jcas+TGisSTq
NrZTQRaLbVBlOoDXF7bkjfEfdPebyRgUJznHo1TjmNajhDthgjY4JHj7EFYl
MrCIy61mE7ypTLl6QyOiJeEP7NtFE/vxD2TlLkhIpNnwV+jysT1vBI2wZCt2
4JD0oxAqd7c++Q7Ixablz6idXCaunNIoG8H/XB9Gt8SoVucV7O8qO87lyhvd
zuweBjTBlYqHjZk5ZhP5dB10V2YmGocBoY+pBrZYtaJwJ7mWps3KCnKURk7x
QK70hgF0SCDshNvqltTQIpYGuj8zBUkq8t45hR1KFfd8V3CziBPEyNKKnTgz
3UBXd82uh+/lj56ZkuMzOQ9uR9zYeXF0Xh7NOvCwugTnUiJMqckA/aBKC5OE
eLhAoSqd9g9rtVvk+V6ukm7z6eUA5zZx2npLHwg8SSAcJjfGJx0ncNK8Zr++
EIi86QzwA+JgmluITm7yyaHZpQtwxKeOm8U0O3crIX3jTmrr1ELFU+odhNtJ
N+xBOuM5oSzrbeOLwVKPGeiiIYQ8J6Og1QHUSIZ4OdCdI/PLJyaJstM11Hq/
yyHvmzbQ/r9wgjk1TOOFf8NRdvSxmNZipTsSxSAZ7nr7ME67cEFSuVaBIjl6
C5IPUpbxdGic4K/TfDm3E8fwmyrhxkW0EaUqw3HBt9yQyh+yenlkDnyGfade
j63iWlO2RiWerHFzSd8jyuPnrNjCTH1673TSaLNHLrhnHMVp3pZjuB83RaRD
V/etRPy/TdMgLETLizrm85VhHBNTcJzKULlwGXq1/dWrmtXuXk76QDcAMM6u
E8gl70R5P9GuLxsFBpGoYVuOnaL9A7Mq4iHni2GWmZ3ZReMCRfPT96l3DNWc
rqQqRaFhatIfZXT3dh9VnpXiDVjTui/8j05nlhl40YMVj0EDMeaEPXB+tSlp
teyl3tOB2wlIRedPkmbepzRUIwFs2oz9eizd6DGQi9FAaENOMq4AoSRmO6IK
0Ww1xMzDwiHtUMhjpldCOJMPj/877Pp7ox24gqd3VJvgmizDwLxGVV9bS5QE
sXcpD+do9y30Gf6Fdg/xKmbTd3umQDmbO+aqmSXyH7+jGHEDJQfi9e2F/uGY
XcxSoF4YnzfmvFaxEgF6jmM122MuHNWbFZTSdKdGrjADsT5Is7SI8CbaexxM
r73RT0gmsHHUdydEMYhwC0XiM2T000iZk4+w6OP5WZVT8wFB+ZKLaBA5SRwW
uqS/eildO8kxmvGeKnyNWOzFofqgFRJ/Ws87x4CXWxH+M4e4WwrJ/9a+cVXU
ymiR33VmalacXVLR5ZIjLmzvS9YsD9OXRh4jQJYgkp22Rqy9JtbxtbXUfZR+
oKNHXu/FOz6UMj93u7tdqRMgiIcC4VPJP1iA/pO+uZfxPbuz51aMIxFi+XmX
UsK0xy9mo1c/DNDVTTwFzPXY8aj2tFfsu563yeyXdW9xdl3HHSCCzp5zxgwK
ZodoZQ2WeeL459Xc48mactKg/Ez/VTtcLIA336e+/ZOreYCx+XkwhqBWCT+t
mwsen3RZQWjvIs1hyKixyytai6rOj14GLPK1maIzeL2JXauDZZQBJK9S1ke4
9ZjgNG9NjmxCLVmO8Kct4ESfWwluOqyU441sOcZ7wv/GqO1wWVK4vGnqGQ8o
Ea6uuTn7Igpyp7UMeunzNTsbb88dzP7mkw+ti6VGxqjMuSWL6rJhB8GOirsr
howPk27X0oJ7TgITtz++F4yaM3ZzHYeLg6KQH7O8TZHcksKF80gpzUDTAiPQ
qPHwX/brB/uTHADWTVJQKadG7xB8b/bJs/jyLBxorD6ocW2U7zy+MrSSg8OQ
oB7a+avwAZOgikLWzW2GGcZS2Rmm+MyTwxFVN/pi9YCWNwUTsK03C1FOQw1c
GBTEURZMAmDXVOalSyjC6TgtRWwLafQ5k5SGBTDkkKEVVdISOrmQxYQ77sam
eKhuwJjnD1LlYFOzmOskT425BX2u+YibHap4Ug5vFl445zCLMg+ww2yUTyyX
axBMkpSQQx0H7+F80KAPTpFzU99DY2ujLGVt+dCjvURgk6k2fthPLhVi5jgY
smI53GiueuX8Ikm85FynBM0skKldSkl17mYXCnkdpQSvGwa+0fMq13F3GUNw
9BZwEfIPvxKaZfAfjrimXmaQFEEMMM7iwRqm5AkEOAIqHXNf6/5Z0XBRYHLU
eJWvZgR4wkjWT13mPFUr9ScCGUbRGHlJsooa4aH0ySyxwwLuO8pHNhARCPhh
VH6iYkfcEb7mODrL2qOe2RFh+0qE9B6wtaZgYlhugv9vi24lSHoQWKHYAlYQ
bBgvN2Y2qRFB4hQB0UKrF/O1Xgpv0G3EU/b+4I0c0zJDyzLCO7lsiwN2xmep
N68ZGNneKqS5XEFT+48BkYAI0h+sx3NxPZRkisGGpZlPGkilhlkElcsKf6fc
ZqTNRNjNSZL2dn75OM/XYIDJjLfTtED8Mi7tGyyNHSQnpl1iIMRGnBT8hSkL
n9RYzJAqGznCi/KK4Li+itpV9q0aPk4zQ13KPLy0cZlHFuyHaVnfzLlKjVuk
zw1UHcxoqYDbsMGYWmVJy7PFMN6qH65CxccjTPWaP9cTgg1IKPum613m9EKY
Ez5FyEwvCHzSLwjnb5BMWe9X0G3ntagc4LiAIdCvvFCUngtJqmoeKcQY6U06
0wlLW8JCS9exp3JzLq9dfTgqJiFyJgeUnKNBUdw22wjyWzph3DDbXqCciKgB
6Ag0cOVQNa/WGO0R9wjiJayncr4GVxdW88xVyyIKfuEfX2gCXh2S7pPBNdY8
PCokkpe5j2sy/hDWHVFPc5td9G8ZPX1SImIuN6OBlPaJ4i7FajVjvwWd7r+s
mykQ9+woQWwg1Cm7QinOWE70mTVGbH4QNzBJVTByh7nlqBAyE83+ciOwVnec
Yb3E0pTPgr4dIABzSkyhUpXq4McqtuvPSMUEc9RUkEMUttliNQn26GQBzTnz
R1rMfwhF8GLSmURDfqOZaMCqpb9lzVgV3zvVfZ5ewqbJGg4y4QDNhEU6iL4R
PWF8vSEuyimK9EYR2tj/G6ozlpEJNTwd9FWrpxTrbno7XWlJQJRfetFwawBQ
jfyX9mV/7SpMu3eqEqx2sCZXsG2Rmca+mvr6VQuQqf54OskEojC/P04mhN3k
2PgyAhXiFKyK2O2k5tVVqGd8C269j0g2Hli5TaSw3g7ZJWCOb46AHMdd9EXL
ekg3FgCCWZqdy2mHNWS0ESWhAC7//mc0ayXCRqkI1C7e1TdNEB93MCW+TVez
XKOG3fQPoZiIYOZ/GdK3x0R+CiUKi0IzB11Taw+OwcAOH83ghNyzcEKEm2ED
BEBBCIIGJ1F3O4xoNBDvfzoNn73RgQPzlZkHSDaY7dQuXMoBGekhsO+xLbwJ
3X+2zeapxc5mkaLOSsBgEZJRBXp0ecYgsN+EmhW2c+AT8M3y/Ria/D2FDjBh
Q7MkDWrNij/6LEZxRD73FyuXgkOtrEyXQFBkvdCE14ykjTu0w6KbPtFC9AYL
kpDoswi0LFjxttBb2326a6VWZVHAShmLuU0f/hW3eo8WjWX/bG5NxDW7nde1
62GknubgVKf7cTZW8DvFeKqB8IUuoNYd0b/6eytSO7/6eO2/mtZA+DU1fD+t
iasg0NUiYnLXMlPfbz8KOXiFfsze3cq0bSzwPDvvIs3HFmAceIx4I43qh54f
wtkHOxTQb/PEoqQzaJoa+t4ssQJNhdAhZxRzvamlANLjjaYy15yWTQkVn1aV
XiXo/t4Qx1wY8jruWDcBQKglBG8ROBx7zIKAxy5LQ7yNctSjiBZlnrrMH67O
SZW2Q42McIdSY0rzH3/4uKgo+4iSYaLf7duRL0NUgZXNVIiYubtuhNdXA9a3
p/bzJsdv4H+IoQ0fhqZuozhIR0l07lIMG2Z/IwRkS7jnuQtRHaVRjqwVprsK
JJsX+B492YQD8DasQLDZipflknIbsa9/vbFQw+vbtpewHpIJL25j4R/4LpoC
OV1GoyxbUiT8sd406KkL44lXnr+Vvf18i9IcSuKe9QKRMp+SfWWneb1SZjaL
VZXp4Prw+hlKYloDrSOrXAnrOJEACyk23jUgxi2FIaFMsAuH3uGdx/5XLxZU
5atMvLXOrkOj2FnXnxXyLD/moN7yvgqQdmBxASXsAhey6nL+VQvRxvkxMEhw
x65HiDbT9HYQRedr4N267wmyg4j6h1za6xfbYQfGU+enIVwxY6DeWsdnKWuK
nkLKcgsMIh/J2+bQKcTb9Y9lIm5ddP5EnBRJWXv84Vs5yvdakvMX9UA/9W8M
tRoX2OksvM7pjdh4YE/RebqrQC0c0hCxHNNzrk4fRAP8YO81Uzzp3D9yym54
SdDUoSAsBjKP2a0NSihZ60mL22VMvlm/hgrC7Cs73lP15+9uSMtBcfybVbO2
PVc/jewNg3qiQpnCpgar9CgS39iBo/NtBP5YUL8WOHe4jBUzGHmjG8UzKVJW
l5eFFx4SnwIsUpe0fa0uOc92qNkL6asesPuZzohNd5wiAPv/lO6ZLUyRoNYc
R0EIUhrSnTk2iGGOlDpCpN2zylGWVUN5HJ5qXRYUEMvICTwfgpA61oSNC311
aHLMqgskXJdidxUdsgMBfQCbVqMqXlNEZdFtckD4twvX3lWW73St5W2QQ2QG
T19g7FhMgX++8EOkICRrp7fvEGzFaiV+QuO9Ia0rJzWK+MPI1eN4MggEsQ46
Av+YCrVmuJNWXlZMoI9MhNMkwh8ZWwkQaq/vrVg53HXErXTdmp5kx4H1pBxT
nyPinKdH3NyTkAvVDlW9w+i2j86UqcaJFwaJFgguKm9l/ujqpyP5MwHouoFA
OJYo1JtY7VUnYre/BHbl0904GGTASJgFcU0q2Vy86mCtZItv1BbaTUl1ipTl
MXDS3yb3vWuuHMvTyjkZGeK5cIYIRjypKRyKr0t8NPWa7Ym6KzrM4UkW4KsS
+QXaOBczLMI7wDYOeXx01WuJxIObIsE8+9YrV7mezPfIJ/gfLWD0ycHwwKdH
hd2OT0uei+cr/jKe4Sgrvrk2EylqtBI7iS0P7BxjTUd75Xrdue78kHpabHQF
q5LsMH6zqj/pR/GezORxBzjds4Sog0yXT3v8wRwjZZCGOIJKYhRuGE+B3D6I
V7I+aN3BBHTE8q4GYot+yrwsV718+Jw5kPKI4caME0inkldc9nTbCtXC7YDZ
TWDelb4hBBuVORH2G39yDxsxZWX0Dx9RNkn+3jbdYLeh8ugNS24h1hh7VyEQ
lOykH0s/hwGJERjnkSzYj134hpiA41Kh3luZNFBn05IWvGU4f0QbBXthx4nS
CihgR0fbJySdxjelG6rddXIa0MJ8HfxpxEXd8eQvYnHQohiu4fWIs/2KxoU+
NN1P2M63Kjiw2CrjIVywIsdaCKPe8VP1z/Bka8onS9lsrc/RUYu1wjR+m99U
ww13xlABTe5x97MaHKyrRRDkPdg0D1fA3HaEfTNMLtzP531yJBtJufDA4EH6
RLafL6Nr/WRrz6YjbfaTABYapP8cysUgiOKPZILu+Kk4obVK+BXsXI4SxSAx
ombEsrtbNvs+A3A3eaSbJDglI/fwq/3Cjw45bZJaAP0sFJg3BFLYTkIyr3UG
6spfgt0SNwv7Nn6fdfe/GG96E/MApia0YuTWhKL3RYn8Dig3GG+xxZe1YkXv
PLk2ZNj36u4K52l6UmzLqzdiH2Na3GxBb2zB87cT6T7IR6Qn4QXanlXrSr82
2Ktc/qkP8MsEjMaJrEyRV8V0zHj7L12Nr5UVvORWDHFSCwZqaEWpOYvetu+x
XeHYulGZZTqB+E5C1GVQ1PITdvoYcaYPQ7keku/Axc0gHf3/sfOZQI2kfm5b
Ifq70dqDcho+/Ka4aSeCph6bxgsKU68cbTmljzmeLO79uj2ptkVCaXkBj4z4
ltCG1L8vSGD6v9otSRS1UApy/L3b6DUQHHqCrOjSkRAMQdXpZEUiqlsN7gQ4
4THcwLT+zIoOPKFlUv6amUNQZPyS9dR2TWijuzw6UM7klBYo3I6Du3RjO2kU
13bu4xrwM50BmSX3xHS5w1/6j1hLX2dGNWLNy6OO++kLh7pQVDeFuEwhSsqJ
kYP23VuyjL+m7soyRKeeDlKjFHlMVjDdIZTeV67VXaTY+HGn4ppKpMqOTCMI
pSq9+kOWCRC5EvdUsmixb1ja/rkdZpD0tiuVWB0uBOg/ZkGyQ+S1naYK4WTB
usGcjf9EaJFpSZBJLDP53ARA4TIWt71kstWNQtPEqygHdVU3EOCRIMyuvKaH
sM3YTZZQII+VejvPN5YkbTvWD4vXWEACxT9BiElXncCYNkkctez9Ikv6OBdP
A+fytoJMuhIj9tYeXAZCpCxnqAJR7T2rMeaVh3hVAMacqBlqeOdtiVvUMqHg
Cl2BQJD7+vlYBkXfIswwE1iq4cHpejtQYAUixH6z0SCEbo68G7iMkrNnHSyx
gCxwu9V2IrqmdhH3BA8SyYJSn/MzCZ7WOr2tYWoXAjQzwNvM2YX8tD8UM8zK
nWsdCrWFC2BgQgA9pKRJNgmCTMIrhgX8uM4PcIBVm+Nrd9BbcBOuD86GKrG3
Fp1fpRxbH03wO8c+YhRdu5xlHNFBn2xbtz+BDdn0zoqLl6JBpl01vmEPXxyy
lDqvuGzRnS52y2UT4N4lQyqKel9ZG0kg6atffCCcNK28+9N7XdIc/9CZ9HY9
uZ9GpffDyZ8aqr60yqy6nF/k0kBMZyIgQBsS4dH17rIPZ5uC967ooqjke359
cL0Pms0o6t3P6qh0PBhI831Ms1cvxF3VkttnAxY44cdqOi4ro838eysdVrLj
xOMa0MfihoeiRFPfRcwf6snHqlutife7F8qhW3b2O4RQpf1WwpvXhmml7RBo
aLHefjnf4Fjj011+xhaIOIHzQinYIe5N1IJvKVt4a4Q4Ekj0sO+LHRMZGrIS
Og8nMF5lWUb1wXbEQUkdF6Fm9npBSrm8HUj1z5M8xQC71hu3RPDSN/X2JDSP
kqGTIj/wlLt0ZPU3FAP9VXYRfSX6y+9zVEZB5oJzY6fMHZfPe0KBF/xUWq2P
C6H4A2ON4jwxhu+h2+9C6rEw7+2RQ0aMoR0e0oSHYmI42u3X5KCqgKkL1LCM
JmcMbjZ1Dq5rgImKYZps4ogaaHpq+vDM5uhK36r8/EmMPLlcovErAcB6nbUL
OxejEQs/9WZjZSCZezsbEGlHfkVOQprgGlnVdrExmRJSIZvq630igy5jcmJg
ecKjE/zDz7bl1vQad99mdWOyTyDzovF9IWmwhPds47mOQ8DSDkYByf8Uo/ZF
aILTuUxPL+B2gt+96Z8YKkdVTJONYJoCmTlv8KK+xhfx71BqZ9mgDmJwX2cz
gYfStJn3EhrENHjhnSL61uJ2MKKYHo/V5nydJ4mWwZfP7546d4ETrsEf59F4
fAULK/c7QmgnovF8+A5lMlbddmTdW5OTMdxXUDmMbJFgQkF7PL2EbHJUv6/l
rozV37+CLLCO8v8G5p4S309ab8iwiKn6msIsaSSQcEWJEXMTmLnzFiqrfA1t
1k559U+Vi/aQ8RlGIFgEi+FYc7b7ChdsiI6Hku8FCitfitSCYADTv/5IYzGn
33TW+aMgCtyeO3T483wCHQJ71t/O4SgZnbvKwISac7MsSOvXrGSYodPLbwcj
jEqhkQwfsK8Zf7sthh+ab/D49xtx2sOnOvX4kZ336IRUDOQ+LLaiC6Yr6KKl
25XYSKztMyHo8GHwFzuU4aDShAIQ/TPlyhVTBOLjIkxxrGK6qXy+BZl2xOwy
kjLnmtXamkG/hjSwqosYy4aNfupknPKQgPulukFhXMgbfg9eWf2p5I8UPCPQ
b9wFspmg+fvlRUn7Yrq+FGnYF1LbYUSK6Xcz8fP3vy74kyz8xaTE9lyikRT3
h+7fV2Mb24rtkGj4rVYJHf2PVVY2Quh3YeKb8Iz6zWxMdiaw47a+2ZPwSZPS
5K+rHB9OEOJva7hx+mBQynTn7B31OB8/HLQQwlIiy6RmMxNwW1MZ53a/vwIm
TIxS8MWcJaH7Z5/1rVQ20GTD6KHk7FoY79jMchwxqvBLY/gapFBbbMq96MjL
VLn+TK6Lpx0jPeQeIum5TH6gGcebe/Tk6DZQVLEwu0CWvx0y8n0FOrl8vCac
RSBdpSyBSB6fV7R79z2vKd1zxMk54jrLEy+K6Py5e7ERsHzhTyDXQwxA96pn
KeZkxecSkwme2GMQjxVQyU3vfQMMhGookNtaXBWYONIWrULmqI8Plt8Z+0GD
QZGCVnV3Gab9WNucrMNxQpEqtjZmFG5j88IINvgDOzsk8c1Wv+pttTc0x8yS
abzLTMOTBJbd72MHbitbPDpOFbhN+DSNRyEm6/Xl4QkLGIceDJMoGGU4T23s
ZISlxQLvJLWWGw+Gj3d7ThWOO4HmPeqnCtdEWHAB+XmKv7M9wbhKqJSnEsUy
5JRisKUsMEQg7sd2XbokKgamVzfSvRnNqdFcTwknVBSa3I6omltRoMVestUV
sr/iVrnZs30oxzXkmte/dXiy2zO+mwYhIz0Y6cUho2fKYzuc1VTWb4LbVDIQ
avxly9l08YmvJMTf3O0u+FN0apRVTJX4WfPbD6DMAuzmY1ZdkBAIbLi+TAV1
L3WX3v4rGFJCX6epZSavhH7zuoGJpdUn7Gf9pKYYURF2sGjN+tIIfIKlOHmj
GUNMf2ylNcPgVYfIDlBvmxAhvhW0+/gJLotpTwhibIFCLApWtAPpuvLestjj
7i49KX0+J8Snfbs9pef8jpk3eHWQSOU1jfLopxj4DlYl1qnW4AWF3TMwC2+F
JfKunDJEXbLjuIk5F1HgrrfHsqCQTQWEP/o60+F+NEW3dPj5dHXxNC5guw3U
F0aPz7iqTR3jHsAsiTeYS7Vjef72dTC06e/Q007ld7ywRnrwpVAc/1di2/Wv
rVxfrw5JWxXmF0YUBt7w1c4X0QsRY7MaY6hOfj3RreX0i3fefIYjY+MI+VmJ
Wy7QAz/AYTcXptEJOscMRDl76r3yee3ijpqA0CxQxDutlDtKzrjktkPb+MvJ
k0YVt/Y+1JyynDgfC8nyKCxS0dX1MvHkAPE/qWaHca7dB0uKgp3rr1JSqTEh
OtSt/F4gC2mFknE+zwiGMoyH0hpK8N5e5y1+w7K0T+0leq7zzEgCBNwMq2Pw
GJr8Q5EIHtki4AmJ4fYWm1VKOR8lxp2Na/vwpPKB+/noEMexTbQzPFjJ4RpE
vhSMQzHqLJL2ktOtrKNaW7gmXlLqeKOHznIO8uSvuCVL2FTvyaR6PUW85p4J
Al1iefkXNGJnWjAMNBLbRWXirSXd6FWRYCYNYxqdxFh0IftyLc9h+njIeXWx
GTT7q44JVRKx6EShOwf+4c9lEwNUKa3Q8IZao6m4lqN4LhpgRQoEEl0Nyism
vYAg74BPNslNoSh1FcZq2nteW6JNQuB8cXUDAep+QXxPtNAh6RQDrM1EK+Yk
plMbZTHXJBYlT4Ew+6YHcAv3KmadnoyJ01mn6JT4onvirHskjVEZ/1XirkH5
2hq55zmSd5dwakMPTAJV5p9OMioCQ83PUijuZ1mJ036Z9QPhOoVjJLouH34i
PR+GI2Hj/kDXkcxo9c99o3aOh+HOjICEQHyKf3nPOA/je4y7EPN73XFsJB3K
c3ocCSwgcfWZ/pF8xkzAL1aCPfAcpDRkXDkDFaZ0b4TyQyfgsVlPZjvnIXFE
hSWtFlJb2030s4DZ5q72nsRpYE9vH8kQsiwhw5hj2glvFzhA6VnD2HCgDSEN
08/pVgvClesysUM5fQrLHk0w/yJrRyFvKhz9p8IlWySiBmUiAkoHGFfL4846
1KCgehzXX4Gfu3/XFJQnxK4UCOqd2AuRV5FEMQ4fHwx5HDlAZ+FAA3OMRn/6
umq8+H6ojCYy5JYPMxCndrVSy9fwQH+FW/FY39hTSBEq4nskITTrrmFXkP3l
LuZsx7W04j0UZlujUGkzXeHC3szydjWrgIrNOcoHVaPH6oEoIVbTm7AJSuHS
VLt/yV+xwWk7RcKaozHgaRXmtEJ7ZVBkBAO2ECQDNOYkwgrzVNpyz/NX2N2w
sYA/HF4aEEP/slZNwWtYPWoWJqzmpz1g1WAr/8vMi2aGAlVmdU9rAIHXjlDm
Tg0buUddDKZ5H6Jl8sxPgtOKORK5qRWU3PYFgUaFmuRdoIBRkyys9TeOH4kq
zd4mYD6vquskd+QDXlExIo5jVXl/Zd1hFx/u9soE9eg9yCIpR72fjcBeSldb
F6miOXB0MfC+wF+tSSa/kdaDnqvZUFnfIR1RHMdHPeF6/By89/Qu3ZJrxOi/
gFwelyFVt32MiZyEDmVBJRJnnAW9UR4OrkZ45Bznvv0E+1pE1V4lM8npkGyT
FjJqUPz5XW1Rl8Yb171snTt646/reKkwl93PzxpsCmeHgSXdArvOq6QcBX1u
beQGQAgNFTVJ5eAIpUMvw8KD709WuqDTI363V8CrlFoBFBF6qHCUE/mrEhiC
CCCjzX1H2UCWZOIbRo2b4J4D7kAaMBvxj3w86bpTQs3fljQ9XrzjRmJEoCD2
h0QXx4ObTs6O2fxdPO96SLRtOiyZEAGoLwi1Pi2ppbgr5BfmTk14YYlgobES
TajeDaDKyLuF9J0gUwGQvG5wx69snUynoAlfSED8QOrcc1CI3xwHm+mjp8LJ
JuzwFU6qKNgpniz+sX6ln1rc2nbjfAcOXQ1kZsWRpbitlHbY1sf6CDb9KCac
LYfRxKC3HHSU+a6u38Y1xeopwji5aOP0JvRIsRr0KGqTcO78Vqwdlx6WjvFL
xn4tog/lrglBZlHxxZ1kSnOLBVcMgZJjpibcNVukTXQ0z2WNVgivQ63MBoSH
fVD2N1yn0n05TdWR1WvoxSikwBPeWUdfkujvjjr8U/9RDix3wBzUcBaZ3w1R
SpieegzZqZGP6PxmENIQNX2vOVvFwkepQvXpIDPtfXEXW0udfZsYCvyo3Wvu
c8oa58vRc/smwzNhycKd1AGMiNjPph37vqnHzLjdZsBVf9w1RVnMYHv92lS5
QmLTjMfvhs9n2GxTU0Z3DBPnlT1TXgGgZuRBXIyOJwqGRC8b+YsgCyTQ+VEy
2w0MiarSxScny/SSoc5is3lmHTUbIQbuR40hkWJXN0PFlBnkHKhmLXirHGsf
az5TME6xTdPNOfzkorbCvN58Vw9w3dF3qpYA/hiNPPCEBXTmS0Cpv7DDx1if
NXAzytcnEplOmPpf/fS/8QQT3aqZmiy8JMBpZ4RSkBoFOIrWnTaH0w57Xg64
qgAndHmNZJtgC2p/K0D+2hetKVhnkRhWDUg/SG9Unh1xENoN0hsBRyznMBHA
nobjPiUYiKSslX3LdxwxCd/WEd/OWMaqf1PNqRrMtuR/EHUuFdo4U2VOvb9C
Fy6OZjgDYM01w8OKYY88sn/+/+LTINqH1i2FbjzObf2Iwp0nnhJJyk/ZxRnd
puOgvRqwu7+yHD8QWjxUWaUx+ndLTJ3xTyCRp2nUbCYpreWGqE0hWR8HHGEU
nNx3TDQCMFyLsauBfTUiTY4Yx1nnsvqObgT5VrD53a5sCFY0RNfFCKVh0w5j
AWtJWjwZggFXPQaTryVg73KFA1IMKpRpWhOiyozoXSZ9o/BAqjRiGHGqXI/j
nCslVSpfnTu+TZWRTcKXCCohawzvaWbezwrE1pvyJiNDjc71igrAfoyed4mg
ZclsA+wcFqDJ1jMz1w27+5ES9Er69DK5qOCwbmN6VMayo7KZhEL5da7dcXUr
994P5AnN/quXrxQXNLuXvr+sPQ3FcJg36lhqNZpu4lSNCFZMZ29XjWGMIN/m
tsl0UvOJCQtMbQyjHU4SOEoZdf41JTXxvnD6hiDOjfptGVU871vMmxgVO3id
r1Y0MMe4roGh+i/pRV+reJH5NfCr2XH+cRWelT+grK34yCfK1DtJF0aMfBR4
olq/8iAk3jb6GARoOXGIezNQpiuwhe2/yOm96vqe0zfRt8/nyFsKtpB2XnAt
La5+yc2s0u3JruZ2mZRCvIzMMxuG6nZmsSbcMik0CNbJwiuGTpHmN8K2Kgyj
/qSiBZrzKwO/NPCrEu1TZYZgV1I58/XCOjTpUIWPYeXz/G+eUp9SzCxw+Qq/
xaSZ82X6DVMmuFd01otq2zr9urrvWb1ZbQXR1KpBmF6npzUFteOJ+xBA3Hxi
ic3JXaAh3yKlagQYw6WFy6MVi+2IaGtKV/xoyKpUrMQA+CK0xCr/n19/4oIH
J72SIrsCz8f4C28iEi5uaW6gDuBCViTr/cSukXE91GkssMsQZWpAb+UhN267
I0Du8rCOBR+UMOzqK8fl6vNbSCborGolqTP5HMpIukdvqlQ7d6HCEcjJbsFY
tfBI0NiEoEryPqFgKUgszYETk6riQCPoacVAfua5PRxaUsaI2azmI2Ho3aHl
sQFI1mxQxLTyNVLXMv6PEtG/QKQgoTitR4XYddGA0gyzXpHCrwEDLK0nny3k
xctrU2aDxsoUtpdzMuPnWdkpZMmRiTq5H5NXx9fXiakRnbKqC8JvbBytxVO7
ilGa0d7nWpnBb25Ne38AINRvGu5/9F2w0jbu2R5F52BiDZks6QIRfQeJ92FI
Aw5Xn1afGqBF4XYbLzAobXoZUsXU6mM2M7yLNt/7jmYjiOrHJorn/NFxpo71
ctEE+2E24ouOE7lL8EShjTuiOgFKCHnBrOxJTrMnll+Dr1OkAu1GDu4nzyNG
/1wQgpvVhfzkFh8/H4Ro7A04pr8ryb5vkVUyCn0p3ttdsCCyXqx5bFQUnOfP
5x6Du1aD8KLCONQxp8qg7CAh2qJCYiomH2AA7y+kJRY7c6hVN01b9+30YZhz
r1hoXgUBoAYhpLoFwEaFRHFtD3aW39odWsCFPoNDfPfHlxNxY+95SacnJy8v
yGXCjqx080/ZpWl2/j1xtMe/N9vOVl+SsiODSpDflqAHpHhqVBxfuDCRJXx7
HcrNbx6KiuK+wWosfL317eiN1/hdFl3p91a3kgMQOOFDQZBKF7vU60rqnen4
VFZ+j/JOfBlB5ZylvZwvfKVOmrWdT7Zh7jD50kbo7IETrz4hqMXIX6zsDJEu
u2Uezb5Q+4cu5Na8AeUqTW1NeGw+T8JYnGUYmANxdd+NURfotYUdJ29/E9Bh
zif6Nusl7YwtSVTnnfR94nq4Tng3b/NGv/XCeIPYKhg0/E90pUgEiIMpmI/2
Bk1Mg23cINUy9aAQK1pL0xm/isl8+TfMw/4XwCW/ggRxDNgBfi9MR2TqkZoY
sVzKaySof1PwzooEjsMVcAnXB2zs3rlPzfIUM5+nVxtlvWivTY9KK9tW1PTe
gZzblh6ScLL2smoBQIhdzo980ovCN78MxzCUx2RaknviaFhSa1TwTP9nSVKT
thFynFYiIPUn7Yxp3jFUO+3XtJWy9OvooDCKjgUSgcZLUStm2wel/oectLKY
+o0U1S7mDqGWcIkEETOT7SD7PUifW9S6n5VpY12QpG4lTwvpYz+zQ9erDV2h
ZgEB3rXZPmWKrQOMfar/WtaU5D6UxG41m/s2PgyGUY/RQOffcr6ZdiI/PBxD
4czfop6Zf2a+Xw67JIsLoRFok9UMxLH1Xm2JFVNpk3tGI7jSVGCcB64bvy5P
uNYBD/Ap1+/kzdDwWhzVfPciajYuXfV9rzYXPESkFS9QoajEbef0nEI99R4l
NKHUs5+PDe0bkmXVyc7l+MTI75/noXBgW/plJj7uf56xBvkieOQEHMrgYOy9
vg4Mvi8aGFlqqble7bTcVy6rW+4N9hjtALzPHzIln95LJjHPstZddYHV68Bn
mL5Zodhq3+zaA4Tmb8FVcJ+R1BYT/5fVEYYD5ZCBTyTYD54NwVG+8BWmdssD
yDaXkqJO69vNmEq8F3sx2rExwF9q4V/Lx7vl8ZMzvHHr5RWDnGGUCaoD+cFK
YIWJ5doWw2AgNwLNZzhiZm11z/Vzv7P8Fd2yrhI0i1HCLk+dqMnhbUjjQBHP
+9ZLJY0FSxTMwqz6nL9P0rrNSJRmNrmYdqq4q2v/1z28T3OFlDP0DzE7o8Yh
NPznGFXCM2yyfebZ0/dHVYp+k3f3tzmauyJTLUGw2fWrebth7D0NffFLWiWE
6MaVxjzcdySdVEsDSQJTjfv3Dk4J2P1JWnaC8/C80bI8RtPmd3UiCj46BO6O
M/2mqY0FBWjqWOClb67b/Caqjx7Dvly3YpbOysbMDH9rHR0cJWohQp0Dq4o2
N0hGuQP00rX/8KOKafIW7Gr4hhiWgoD2AABlOtTzzGzXQ9ODUj9k9hh+dNFy
cmQ/tN8VE4+hUaCE+PkwCN/vt6KnEH42+B7xrYsBbv3sXY0+7t0kkEPUtjPn
Gh6t3eoKoO9HlPV9duA5zoQlDGH6nJIBjCCo4QskDuh7J5v74TzOeLs2sY6D
P78RtD1xqrpONh3Awe67ZON91nLunABwdSVSj7U+cYikJCT+HrQwx2ZP2sh3
aSymbkz25zMFnKnSQ3TgePjB45DPXS55v4nvlXdbdAtk85IXftaN7/YwH3J8
u9izEtg36U53HMGK+0YHxhiq5M8HhhkjAnTqJb7fhwGsyf7IVK5AOA3O9TI4
n4ljHLCbLDgQY9OmobxY/p1Mwg6VCxjdheAYKMrR3/UvjMztRFJJ+byydPCv
Dt8GHkyT9ZL08VnOLlo3F1aWCoTkn0a5MCwToUP8eIHPnytcj2AM3EcU22CL
3Zkk9KAEPpFDZS36U4Dsz2l1rReRurfs+0DVnH+R4YpqmC8ZjVBZBmkPXbhz
Ty11j2CPq53zr8yUa9Ozfq8gJ/mdlIx4tIMDUISNBnCsZepTHNUM0AUCMzcn
AzZAxgtX/Gb9vS8vsdhq8J2g1NsY98+g8B6DLrTV1+AACd/nXYham5rI/zN/
xcsK38QE/sHT5OVuIeeJx8IWWguXMfRwj0NvHGt3Gz9AvtJmNq29JW8nX0EL
BZkp+HUH4CzP0Pc2OD0poEKQ5wFvIyLyAnLuamWztGzqmIzpNL2nC/0SlIri
kVcCMukFza6t9JTzDYrK6NqStY4bK5/SLexFbkVp7KZ2iyNQhTWbIKlNQyTw
jC3yqryjcUajGaHNXiJ1Res+qJ37adukZbMd6AA/00XWRoAK55VFNmzxD1gG
6XVb7VRikDF0tqomLZHuMM8w1RfF/CoEvidG8/ryIIHZIeAf1vYoOEy9N0xL
BN0OBYzAN4d1o0/K6IXXPWjP91296/Wu1VRMdzEUYi8ZUQ8Nvi9PJmUNjkyq
ohZz8ldyvKCDutpNLRuL9osM1npmDWfnvHE6U8oRZjbwccqZvD1GpmfeZcmm
d5FduqGi2vsMMzaEOXoPkefMWs3d/cvoNX2zwZkVm3kuU0rj0l52Sc+shLPt
lIx6ALrTjmqfVOd1Eupyqcj/k6i2omQITvn4EKe5JSTCqygID4gqGgj/Hsp9
P2bxjsjBCWrQtmQQY2BExwu0Q8rcaK5QFaXNNG7DyvAuUMwLbKkNMC8uBCpA
m3b0aa8U1h9WjnNjR37WWGLP7m9v8J3khdGViicMx4+gEWnJVgCMqSKd90m7
lW2N6bh4QAVrdJaN3fKNtKuCb6W7ErEbxFdheAV901mDwgOzPka6od5tw/kg
+TmMjXOT2n+yqy/LY6Ow87S5HU9Gx4CnAkdvqrecAsTHv/2X6c32+WwOfyfm
LAZb+os6N7DdEK01yjTxECt/OCDVtC9l7LPCBtYEh073/kXV6rIaPvrm0amB
At7K8sKMS5iIPIRO/Eu+ipD4d/LkOxmjQ41C3/omGYLXQf2PEWOBQU2h+rPV
KyXy2hvZzj7gZLyQZAkJ89BthE3msVHpFSYxz6kY/IM/P2gPSuT78HXmhl2u
Cx5JhruFJa82205D7LFGT8Dt65QG85BadqCvq4a1AL6FGbetdvft5SvmMyXG
Jvo9zYoj+CVFdBA5Zhmhd1FyPGt6OhCurQH6WHTQWsDGQNv6TIwjKQhXeoSx
X/if9kihMSTaRV9bz5QB+29lCbI/9aloFCGoIunurQFJ7HWZE/ucE1tGdOkb
g802omAiO86jSwMzNgGVDSQmOpygP3iZV4HAIJXRKEvIvlIPZyQGfN2Tt5G8
i4whHsMad/smxxVgDqm3y1y1AI2H9fdBreisZVHUSORytHHTyQw00R31ZVwc
uhhxKSdybTniikUwPDrqeii+9JKH4ZP0jzLErG7yhs4ePGdnV+FZe1jGuP0l
QdaQxUMiOFsLoqVsJrcBCDGPtX/K7arlrfYiVbKpWhgRaWQDh02+6lPWzTSr
Qe5dKllrZqc33y08ptfJcUODpHCEYpif9+k9lMd2h9MwxXVOHIwq9lQ7ME/x
URoBmVVo1lrM6sJ6pQUnJRu4beLX0hfaa61eAe7N1P1/iyMJ9ttJNtie1p+n
Si6++WbzFdfEBb7hitP2AqUCZ0EJl4BkpR0MpOFwno7lyY525WypP8phpA0b
iW2cyBzx0OXeR4fXNOfauLpW5rlaysSu2IaeljznpjOz9LW633kHlkORIa6u
Hf/KJ3BelHqad8qQLPRSjvTt/pEWdxAwO7CL3FiNQS/7Bar+YWxZ+ZDY7s2K
n76AdKJHUvDhWy7ETkbSCrM1XVOKC7RhZkXwncmT9sQl3bfCp+AZsJpqdKB5
12E9u1IwOC2t90NkbHyFA28Q/LpxJt4qYDCmdhqPOJjkRU8giz5H7poTiMmf
s+6GrQt2ueyCEogz3pCLOl5q2mqiUkylJIdFa62PF5HK4HjyIf3pusrmx9m+
YMl96mAXZ6yclpJUdjTV+HnRH47KitXR3Mb66hhfVhKIIRB6Sp5DmY7la+U1
gkj/PyRDwnlnHF3FunAobC1sCduSRC/xO8evYi4gg2KKwumBNfK1z5dYbLVm
MGVVHHuBvjk+4MnrbtmpxGvJ8bWPAjP6WMkwLLem+MqHaZ24czKo76PQEmbP
8LNXtK2laWeI3OX8POcyKTGa19y5iGxiA4BISB55DA6iHewZw/5w8DA3bPif
P1iQTpUKYeyU/BK2i91joM3Ie7E8GKJOpTjkPt4kr3HfDAETB/uX/gmS3/om
Cf1+BUvRbAI7Mvlj3v6KqDEERTaJIeLqR87DVKkyc+ds8MbpeL3tdMM+iFHt
DMkjYESJx+oEfPhOPhxJgYmxI41PS8mYdSy06jxEY6yhKGap2mAKRIqmCp4D
vmWKwc1k2zae+TLlUZ4pgA01ufNoVMp6sEqQ2c3XlFuO6+sJb2U1+7WbPLxt
O3GgK8dgLUAkBAaJzJQYfNUqnm5MPN2Pq8JyqIMFGNtVqL7rnVm1MFP7PXNc
Aj4TsRqqfxIFfZARkWzvxesjTB3uHRI7zwDbgXw3Ug8RlARpd0x+gOt92LX4
DOBm3SxlCTpSXZK8gW0inY7Ozz5hOWTx0s7CQ16t05frgDO2VtwnbCCwf9Bu
7i09xQ1QRVEMhWM8oJc/l/f+vu/pf0DIBdzFLv3s5MT29c+YIs8Mxr/mHLC+
sbhdbjM1F9LIkODuEnMypPdLyktxI6dJc73ggwzOG3deo51xR7/lgfyySdxo
1zRJ3sPo6u7efYlQfweUSBNtt/AIigu8a18MuI0gxrUmfu+jQKsYVjpVtT0P
zvxjs3wp9tY3mlQt38xtIZeIa1KixISUz0UknzIJbnGafbs2SwN0SRFQ7Yeu
ILqVyfSl2QGOXZbOM2DtwnJQ6qc0h3mn4U3wKMTCq3dpEYFV8oTKkymTc06h
RWdcDZOp2w/XvEqdWeNQUSKryE6dVf98CvoEPPx6wIQPAckHXFSCvn9Hy6YO
tBrCcUWi/O84WIaXUNNVkQiCFsc3ciIIB4+UHVFanUuQ6826jjSXi8hmVoun
pWy/pJYnCtByKolI8m2Y0WwgY2iqvQflXbQfoXm5vV6yjKLF4pOl9NfKDvSs
dh2KOabEzPA/Re1s7y9oZdDXssNGV2+E1xiPwiDYoLd8vrVgrnT4CF4nrAPl
RrkHBdWSjQcpJ4rVL50eGoIOeBQamIbDo+2HiHKrXQOFtLmjrWYNQnzVRnd6
QtOIbN+dyu3m8E1TNMNAWkw0PAOw2zsyqBQUSvFRFnXuI4mMGKjJtraDH2Yi
RT0IV3dt7hxvsgSCPmvwRBDK2wsQWEOu3wD21iNbrlnOYYUodxXr+OqzqQ+4
vUDgLoFExkipxTHIkAOaDX8pP9UVZesn3Uw1NQlSjhcZtvn0+gzv4l9bIm1a
2uJ+FjtiM5DU2ngDM00rVgthsH64N8eoxpedL3JL/JKVBP5Aqu43MhAR7v6F
w43mFor1kYxEyUPV2zE7SvVZuYhGnT+pGJqW7m1248giRO9LFeiFrZ0i09Di
/ElZdYXIyh7UZ3jNpmvxMSwYs8tH44ti4Fz8OVNA4PYPFvk+vqnMzcbmCHG1
BWJpHGI3/kw+nmWTWfgal3fe0a1srcQyN0mMbYUX6uKgSBFy7p8MYZiAJSI1
Tx8SVK+EQLBWOFgg3bHw04qkd5vFR3FaKrbAta+eyWEOr1rpf6URzPJqx6C1
6x9sAr2kfSdiCC6XT+zAf8VDx7a6md0G5souBI3A9LX3zu2lExntcWQbEOmq
doI4oA4GYw5iBghS52Dk3hs1NRkmHgHDY0o2jlzAMtDKskvbNrB+Q9XC5NqZ
ckizUjUn/tMI4R/u/W4M/UMvsZNdW7CXYrWIE00qR3UE7zyIrptAwmHrNMJJ
P1EWj+lTw+O8Ulm+jGdKUMqiMlawpp/dwlSfxpo47qjbGEC+ojT/huXV0cTa
BoeG43+OPTfrzqhuKknsWsIAXNZ5wCj2aim2xr1JkJvDJsexhZ+bj6fqqfcZ
Z7dG9AQ5ZYzLPThRB4q/RPatfKa4R390MDfNJhUX76RS0aT3HYdvlx0PRo1y
XpWJ7jkrWBc0oCIrGCvoPJ+wgUIhP5tc16wIxUHg7jUeAPacP3bVlsQ7DAgn
8zp2GwJ9Qrztbc+4vvw/d0YdHik0gQEcDrNkDhZbG20KFzhyX1k3+iPgu+Yh
wqzy7iO4Mjaqe+fXI9tGC69ri3BFHIITJsZoui4LRCWrqPCZNeaFEgHMDJbt
4boHV+Ol1RrDnskpGxd0Im1GqCqzdnwLpbxDFfcsXV2KmvKDXOdqcSsc/05p
3ysB6niPKkGgcKGyooFMTNO4GtzF5SimNVS8kX2WaPxIcrH+DH4XV5jTClCw
kF8Vc6W7bLD64YX2qqipNbRVoHNFWTX7jMpC4TZHfe5YQYz/L95CoTugz88H
gqg8MFoTaU+b1DyXZAbqUMuEdOaY+MuaS9RVqg0DpjPjE+rZQPa0vQN2jXkV
IceHubcFcmRo8Hb5F7r5iLm0ihzbH7DYq9bdqIVA9Q+RdFKKq1WXoaLQCkMV
x9KowSf+uBUO2JtLK1fTX+CXoRbCZEkCEaNk3RnYW5z1yL+MoUOTTzM+S2JC
X7laFptGo/5vbDWA2kktGhNrdqsOH3NSbr/+02kAB9Xih4wNEIelLDKxnIeF
6Z6gV3hYBbdzndl08Hky3DqorYMKy3FbU/0PnyMFIL3NRRgYxRQR8Z2gn7GN
DlK6o0bHTc3tsjbBWtTP3pDz1l5VpOAyS2ap6iX5MHEjPkyu7prw45O8rGyK
YvTNtrB5kg8mpRYQgordZSntRf+u1KmF7hEjyT+PX0cSAfCBHtDrvSY9cab2
ilsc1aUmx096Xm7NvOZ46aTaj+eaoq90/Hqatq/EKY9ABEBBHFIzhRKv5T+B
3bvGxcuug6vVzDN1JdS4zp6lJrPqZWw6ol409KJPb30DtbmtGdLWSWaJ6DCB
29WnIDlob+RlaQAYOZZerzETVemKZ9jA1a4rZXSND7gbn0bH1WTFgYff75Ig
+FF7En+js9WWKcPNW9DZrxDDoYAUafGmUvYKlnng57ry2VbBe06MsirE7dTt
DVrkxH+v0teXr/kcW+Tqec6e2VvvcJNnerKA+knqhIp/VSQjfcTsRdhKT5xf
fNQJfLAFNnWl6zNk0dJ5015kzvfEqLmDepOq2y1vTlEZ/XqhGs8PpYcRj3J7
FZ8PvW3h9A8TgwsPxHbk8TcqvRSm2I+NVJNN0y6/TN98Gk/GgeF1ir4HNwPT
PHUgmaQ4N0CUilxs+kRxiCwIaM9+zg5urdFlzC2JUGEVDVpbYOkVJXZ00QNG
KpUb/NaJB20jdt237AnFmjNJzvhxLZKDkOQOXa6q6K96arJgKWewsJnODqbV
EuY8TRQg5cHditUMzXsuO1/U9oLI8do0RHi3DREXN0L8i/9EmARg3n0j3cv2
HJDttqbsrqvXkJnCQhGSkqpmgW9y1Upz4fCEjjnFI39dxxlMcdhWM9ck5JfA
3DNOQ/+OXVDl8OjXqnjHF+nGf2zhi6JMKqpSjmAgal2bJqylPpAV9wZdxKAi
wm/76XCbSJ2T0qODYDYofkbM30/gSLxUm2RB+wTktgkGMgHjCgv/hHuYMzTL
6opy89Vw54dZH4wwxX0iI7gfVyfRynDhBi5gl95MjaPFsyDrKm6GQEAP/Ake
x4XHDPPOU3Q6fgM+vrRJkSv0mHAl00VXqLM3jb1wvn7g3NWwp3+oa6f74tMB
9AK9moE90YGv4KAVKOh6g4ESbPLEVAeQsHG84Dkxg4T3RQHHfANa4fJ9GdvK
Ccrw/e1XjXCwbTrQaah5p/0DSWr+bxXddtSvxypqcIyWYamUQcU0gOViBhpi
PYY8/HbKVE930RI7HTwxBMI7UCT6IN1AsLAxWQvTrU96aB3uKj/RgSO5BXR2
naIstS9uetMJJ42cIndoHzHnXX6Rkp6Cw1Dh5Ussum+GKYPtCIohErR2I0ux
p1meDyWlNy0tpX0royFGDWSX7zZL3Bvl1LXgE6HTVcIN3oED6X1TjE1No4UM
yfP9P545K+2jp6nH1+Dv8qg2MMRY2r9A2DtpBDUn8/dAt6MBfXG5tsgCi9vk
YhYbZjP/osFCDzMNX+mw3ovGoqELV9l0A7Ml63ZasJeETvA4AbgoFHXKnRfA
PMSWYKwO7Hyab1xa/GuEceUJvsBuFLeunB9AZbrZ4CvW1R4rTmSwqhyfrSxc
3tauSb8GQcagpgSEH2QC9SmuRD6v7e1pGeBuOguzwjT9dkLiOlCbP6xWcyYl
G4Ds33N5mWn/0CeoUPFxpoLX28bgQPqLAJniNP8/boZX64s++FXNMsBRZVte
3uNa7xGad6+tTo6Cb5fpmnOW0fJaaVBsILFSSDuRAVziYPpfoD6O78iR1Vvl
ipY1crN0HFKDdPn5oOqslUKMe56KPzUQZL7eQXDE4pbIT/vlyc+LJ4xOONXC
ssPIHd7e5Ie7VIN8fdAmyzyT4tyah++P1k77vX3D8BC8k8w33IYMQm0pHUZj
IG4C7z/i6GL16+2WOhPpN1YBzw+sAFunD7QOoAMEMzFZ9NbHJFehJ6W1WR+R
S0eeZ0qRScM4nkJVqM4PMc/ihiM3CgFCkPhndhXL4bS30VDybpdr27Bz44A4
ZH2KRZjq3OI2OpjI+pwERiRZMAjQT/nV2tNUlvXbowMJ3YZsZfLmDNyByqkD
4NaMa6RPL7OLubkViPQgacy4zcNlz8JTqCUysFz2JI6/yLgM8BCGiA9dEMj2
odyfbECk3BnQWneEcO8KebMCjLnTJLFYigSq30F3B32pZpFqCSwKu/t42Ash
2iNX/cY8Vv5L50nSQSebOqbaPKLWQyZYeSNVzJBzJN6np3LkWiwkvqklnrVT
BbgbOWDv+6+YhHZUz5UyGEXZHXzQa45o05DS68VktcHAE7LYf4VLrQKqPpwp
50sG71eHCQABsIgqjhcW3hF206QpMEejPYu6vCzOBl9OobwOTVW8J5Ndav+V
gngUIVmr+ZrhNfK8+UoCLBG0sRIxlwKk9CcyZKwRfuwTLaFna8cy+FrHQa46
XvkqvjtcYgrTcqIb6TAb21jifzKSRWdQJIEM7sPdNO7ADMQoc9bgLgXl/lkQ
BvKuyIH7qX4VEWisyRDXAAaPemQT6bbcbzjlrr3HP/4ZEqPQmwg3Hf3HJ3Xn
7I0T9g0zM7RkAtphdQCrPvyUkeEMYNjcPjZp5uZTq8ddKlpoJCXgJ7ol3M9t
FWYcH5BXJCkzNiLQESeFof+SuvYoHhVd54ZQfBu7oMZh7BhKa5Bw3tGgQFQG
JoqYnuMlbPQjadiN+RxCoqW9GechMpKfWPyNBlT0RsTBcTJ8N8twb57o2J06
5PS69om2cOzuMHAPHx4CwEFD31G8zmrXYft2S0wd8RQVaL4HSPPtJAhdKp5A
DQv2ERWQylSiN+wj/dXxmTKyYIXOLRiwNtu3lyOrdJaShlynYP51ux2suI+q
0l9RIvNkdzeW5x6WbfNCCA0/hkH6Ri3Cvf6oZMSo70osNZ57gh4uG9O4P4qS
6UOctjcjsu8wcKv94tFKUkRDFcnPuf3C93GDKTl39hI0ySJ5iYvlARbyJIu5
U+K6lJK+Gyb31mfKOZYLbLE9cosmeot1A7uTJlVWnH7dIhX1gr+J5cR2Y0P6
X943vMwFSMeqYVOF6cUp2jrkIkQ7QkIXnlTVR5tpYADJsedjTv9RcZAWVVIw
4/CpAHnNhahEEdPBCxW6l80wBO7y6SyOHjLtTb1Qbasi/6PIMnyDOxBTLM1f
JyDGXmqFpI0Qv8uZvmzGPsqvI6dztjwaTEZMcmcQ/TXmbp5d46HgTC9Nhjvt
ND+KOsEzrLNk2DAWwFtiYEaMSlzrzZSZ9MCC3k9E1XDllDmcKV+6MsK/cO9V
coe+bg0Y2t53+dVLHBF6fWfVbkDUAeErKr7mditsjVmVxihIb06YbXoR1pB9
fncr2Tx2qIGKvpBs1AIK6q1HZXOHFlEmBbDE/0INqwpaTRtNMrDcoTyGciFU
omay/PxCsg7HdFKnvAp0Wi9hCXWS6vHPEbKDa6VE5SdV4sPqiGlMPgya7tIR
Ga0kVSEveawjcisjndggaWWKnltKkg23mPXHB9C5ivq4ySZwfMywZH+kUcgb
LtBLNm5DtpjmKIoLzeLxceddVvUYCASywwlJCr/MYEPoN8EuHcTUNeRcFXT3
oIXop2xZ0mHASHwzP+WHT1Ecg/2+EzS/aLtrHeuPBhi+QBVnsYnjfzPJ2Kqm
gnF8o0U8d/8+DOEDufEphtl1lexMOyqlZ1UD7fJlzOuAiz29RKg26zKWfwwU
YdldW61CbGiWjsZixMdCENwLp305wLbXX/hI4D/0no8XTt+0D6BzZhjnHr8I
McmoIUjuLc6ECHVJC1l8ygYU+4db7UfHNHQCx4qMdgngq9vjDor7/lSrcudm
GLvvIQzfSHccfe9gfo5QbyE8W7HCoGZXPL9JsSjMJIRfRYeRYSUDRhRLlqcw
pqdkqlDvyR7s0DLXThKi+Bof29Fi1htEL0MUfbwc6cYVhClQ+6e8MayqSf+j
aa7SQoAY/ETxpHQfwPZ54itgCNX4BY/MUSi5LGjz+NhlR0gz3Thtm8BK/VEx
nvZ0Vlt21C0fbw5TDhitWrEJI0u4vGawmPoW9hPYmwRUluGDLID74UYpzm0w
wZ5U+PEF6NGeDbXkAD5rQ2SiUthP4KAmqC4XnrHAU3D4CrOLoxA+Pk+Es/lT
P7mGtwJeyUbJvlgHs7JtOfpMN3s1Q5NbJb2Y7nLoM6FqE9/xJSM8DVcWFLVn
9w52gZPbf7dpN9nVzHwtWm1l5Dkv982nizEDZM5oYR53LPxM90ay4SL0c2hw
ZBWaqppj6gFp7l0hDCCSwsiQjxokW8J02/VbGqSia0q8Xh2D5pGAG6g+HMXw
oujtxMtKPcmDDFI+UVBN/sp3lJH14eS6EluCKJ+lsg4IZZ2Yhg/T6zbjIPNS
722Jliw93ZvRH4HkK93zfvJTNZNaMkcTwVVAeBxMVZhpOwKe8gutprtQG+k2
YJ3wWgWFzqvTrnv4h+LwUUp5fgOKPiJ10c0xdSRLC6BDaQ/2C0RVV2wg6JqT
TRIi1cqtMB0UFiyI+YH7Zbxq8F6t4XTirNZ3R/jBweglqEqVMepuc/bGhFGs
c7fZnc6TzVeMhOw1eD3Nl188LwY3MkXZLUYFbMPjmRlMCJVNfAsO3XTKz3o/
rPPwtarPkJGnkq5iDkZn6VhEibTEAKRwf6F99/HwNXruLgOp7yUYDOuKE14+
bd0szBM/RMPukvQZxtA3nyb2cXcl6AKjQ8bSc5H3gEK7EMrKtfSpAldEHeIO
aQvagEbmqu1fMxzyBprMBYKfje+3tMUdR59DSrbpldXru9+eUAHn/qhYRK61
qSOtoIMLxa+ZPiafoZb7SCWdxT8HXwNLp+itpiHGnzVIyfw6sMvN/cesEXm4
lHtwEpnvkPnb/GzxKHKPgL7l3GwyEyukRSNdMmSc+qX0IhSQWyG6HvPxxIEJ
6aIJbzMjV00mwWZe/IVUI4fhilAfR/Qh5+jnkv56ylqExhVgO9ty+Srvdcms
6WFc7zYEP3UzqQ/CdoAPHLE1YMXdAwWyhfxgcbfpeKQUOHoCfWBtSdbvwkz4
wrjaLJMwkrdMdYNQZ7NSy4Ote7YoIJfCmuiLt8jYlHeEMiYmKS9MtUbXdqy6
CmOk6F9HKGNfj+/pCd15N9hmvE3Y5QWPIgRhwVkBJKGl1B8pYDFwcTuucB5F
vcctJQrmK47IrhLFgG1Ja4NpXkBhNDXbN9QifuWSDPQwh/+4EP7UiaBUniqT
EmuSyf3dwh8a3Vrr+YAhazmj+DwQi7GqhiG1pdAnTkK6M+RbQSkOVP47KfiG
3CDue56UmbjmNQ+Ut30lrFQDoaOZIbMTdR3iSQ009GKyhpbeBnoB6hpYDTX7
sPmhaf403sji9Xx3Eh6ZPnoh8FbkhvQFLgCNRzfVlcI37OuPjg8aiHKPblo1
m62QVwXw091la2gfmfHqn9k2Gk3Ac/PSMqd0tayFTM5jP5CT/RXd8thaD41i
z+goqyQlGi+BMp35IoO/8LW3HGQy6+57OCcEtiWSjATxGLnphoVI7ad/L6Hr
8XSPLlqLZn5G2Ge8zWJ4FaXiAx06yLx8HtfzNbvpCdcBo7ZOyaXHpBF1xX0D
DiH/wtaVIDhremqbbeJIelNU9xU7+NrzbnF6hAe1Fd/Xe2CrYa7OyuJ3g+dU
lMjZKCAv/N/GOQT8rMv1JKNnLcNNvLXK9Nt6LRf3Q9zsxMAXYo/IV4VdhqGf
M7X8XkwGc5RScSX6tHDWjuCmk0bFk8aAuTTAUaWb/qkip4m6+/s8UykXsdBx
4hqm9wwyaNQ+3oZrnMGg2uksjM4opyTna+KJXAX+S5mdHZqr0MmSOiIi70Qk
nSGwtuoCtcoW53Y3smALzUBmjszB1tq8OBE4S1iJEQCZTOXmpwIx/bsVw8f3
UhWhfdIrBke3H1S5+1zoxs9NC+PRqa9Mjyed9oKm0CzQV/1sf1yHg8YFHwDF
rGpW/3CZuNRKeKS+MvyvmmKlOAPBE1pt0zb5VJ1RrfbI/t+1EYsajzK7dUte
PMDbCfDTG8gVW3TVHEZgB/3fqopjrcyR1eqkkAqH/t5KK1mNzxDcmDXyUUSV
Sbtff8M9gWGWjumZtRGybrqtgtidc3jaCvu8smoZUfmQuXynGfmx+z/4o/r9
XtWnoLZqicJU/hZk4SBVnA6+W7Z8nwIxKpekkOC7NFR6ah/kf3s/VVLsvC4p
f+PqRZOxoImlrMiqrZyvpQaEakYJry1zxaN58ITsM4nf/Gma4IR01XcUWzD7
L0p+QVFYQPqsz6cttlpkoyGf4W58Vx0fYyav1gBPOF/SJnSuf9TAjpOr9r1I
r2Mg+dsB2AMunr/xaNv+mrPguQnczGfAtk0hQe434NG6MC35F4YXykm8X5n2
DjdqXnZrBeSjvJtXfy8I0zgKlY/tq0tDf1PjwgaUAaj8Kme+UkzlcsxlUPe3
0PXQoW8tj06tAa7QA+BPHyMGdd+vuiNkt4QOVy8eCFeHpzyaNQcleJ2VcSYc
qZBTsaZZADf6s4DoCHxN7gRax86up2EAd8c3VwFRXx/wpeHXX7jjP8ZvgzbL
ynDY8z1TIsl2dYA3l4FqNaqbBXfKJnV/soCFfaXt27i8n/lmhaegK/+ZaEj4
8DjP7QLe1VG6nB5sZxb1GyEq+ZsCYpkO/4a7Ktqt95aEN3oEmRAinUwNH4Fy
Aw1zbWWWxQ+FCLsz+l8MbD5/vAw/9hWBd8NUNE6TBsPwqDJ9Uz89ubyGFx8e
685Z+ZEnCRSm8uaMn9tEurwI5ecZj//c7qWHEx/W9PUxkHQjaVAP+W4MJWLl
0mttr8gBLjFx+NKDnRMlylVo588X41yrEapQC5nTLpvLAbIgnPC0D3xeiaVm
kXY/lbhjD0DwkEvvGGkWUgXCTbnLzRBUJg2hkR/JVm4Ci7D6Jew1I7ZhNvZ7
oTrW4bqqVtTXSC8JYgCWFiTX3luiBuoapELNi1tGdPCTCAxfa8RAxuIwwtL2
g0x1bblFLj6q8r76Ou6q8c4qb93EPhbHqKce7vKvlr3KSX7P0uYb6Y9c4WFj
EuY7/kS8QQByRhX+lKPszo/ummcymWNE4JJhkQS0/o5hCz08Mr/FtbM+VC4t
WLGsi0WVUHkFSNwxaAK6R+YJnX/S5yS0FW5S8qlOEIMW3uBM+I+6jsag5d1L
ZtIe+9v2JEjnJ/hZ1f5u2R7Ws3vcCBdd+Ivr/3xfbzSbovWonsPkcort+QeQ
P9DKTI4JZSdJrq5c/gFRKF7IcbIaTu68J72TTAn6nPWDSI85qfocTgdDCTzL
K/FMVdLIimZW0tUqrZfk5cjHQJQoVMQYNqPZFPD8h6/BARRdAlsa7tZ6e4fb
y7H83y1eTNHHCXDSX3sE0t7FvgieYMdv4oyxyYSa0BHWpl/L43lzz/4aGoEC
3Frqo4f8y2umW2l23Ilf4P5sKWHJIveUNBMzS421KR+TqTyzPvrbD/pwHFHV
REing/gHr7MmikKDe4XUO5hjiSiO4kqeHCH4C5a6xXXhxYBkmkMUvEXWjCxK
IuVu7dVjd5unx3gx+xKg+BjlYl/iLT6kC+30Gag45ja3If7gF6Q4Kfv0llJV
8V7hFwadGEp4IgwGZHTn8YRzI3aevuo1BaQZ/PR7KIxUnSkV4mxDUkl0+SlH
d3d8Rbqj7pyFGw9Ha0kux+1t8sTqwrIGuHAt+dZB7WgvLdLZD+Cow/lwIVxq
Zan8hyCcyqVz0Hbi8F77eXp7E2kVVvzww683+5SkLVvlioybOEJJpATn47Iu
GBIojBa8qsDkSOWOIaD/FGYe8HTWwz+2YTpFqENI4Mffz11quNxiomtlnLY8
jGjR0PPlakf5pNlqUVAVSu2qGD6k6GIYvGKlBE55FEncXPUYZmecY5Yhm0Ps
ib0KQPxhjtCNaThSUt4PfE6trPNstimyWfolAo+g2GGtt/Ofsev0MRQXtmlM
R1n3Hj/WWAlWu7TZimEhmZEPT8LFpErVv6KSu5FE7wqwMyYfEeJPPsrTlcGo
uRHa7WIRNsyCEWpXHlJfycGDmKkFqsbdBbP6PQ0NeLJ3Q1urWnfGan8A5Fhj
dD0jq8pV5ud9QZA9SnHesnhMvxOIHf0KBKCOyLBGwCeDCSdPUosKR8w5MSii
WdWcXAkD3SFEJgFNIquF+I14AO6pHMRngBAOe8DSh4/IrYVsm6eNdUW4GSON
of4pkETOZSrCB9JNulh1w5nEYoC9UCLjS/CkG4ARloZvwXXpLdoZD03an4hh
VYKXqmgjB3e2ymuxL8/4UXS3psdcf482FE5Yu1GbHPeDHUM9Hed9obC3y9mB
DGZjDV9RkIryXBpgAq/6tYYqYCiS7IreVQrIW5O6BBwRfR82UsoIueMAqBSI
9browRlmdCEEFbbCf3UnlRJ7mP2quaf/Cf0UCLjHUz/kqRnY7JDvAUm9fHuH
Hhd83PmhlcarCkPSYuPwLHObiU7iPh7OF40tah2SR9VAk4/SHrdB42o3aEtH
gFpDOOh0KUCcShAxuJKyo63uInZeqZJ6jE3B5mafZ0ISGd/cx/5BCfaZhLKL
ciU4Bemd/7vQtp8XYRbcKRsfsu2P8/si7EptMS09L13UIcGApn5u4guwYsRC
1gXejVY0irtW9B3x2fobmJMSDjNk05sDIsanFzRAlMZx0DLQGnvvsApM2nb2
31l61nmCOxcFAy+ow5fkV9T3mDzhEt3u12WbutPwAacBapY6KrJ7fEcXLfKh
5POfu3bei9pX6MQiPe3HV2U8Y1q5r3Hy4jnfhY9hDVm72L/jN+XcWj9DZStm
3H6m5JFMhHqS70ig8bR6+U+N3VYjf/UwhKy4KAWKMH1WpQo+CYDwFcayN8S8
YD/7+qcOkcqSn/g7I+U56nva76Rj79pVAUzc/hJjLQV26lNh63mHZeZ1TVIL
r4fLjDagD7wlhImnY/pfZw6uReMt62L7hTGwdy17hvu6E80CJ8wbF9j6vmlP
arRJzx7swwuHXMVm175xwhoS2YLYzUtMyP3uptNA6LYpULM5q55BJEgTB75k
6m5FORvpj6Q93i0RntUq2AmtairzlhyhS8BEhQkyFYNVKvHQXPvk/Ea0eTKt
V2fxTHbak+krS9ZYNI9Tw4ozKeOv2uZgm7XuKb4JGAnbVZsDJd0v366Kh858
k1CO98p8HWZylWZxlxlXzOBBvRG7z4xg1CJNPxNb46CUcGU/H83YRW7Ki1Kr
W29aKsVQsW5gnYRgcdcXGdd3BWtDpfnrP5uZ5aGRZNXB0H+rDTBgp/mJHb34
IT8OmD3ylP39gGMd8y4yPFNalTP4xMWx7FvW0PQqT+OVU2CeCfHEFAZoqjkl
X01UDQuyclh8POWdq4BDLtPNFx1FCqf49Go8QIDLcp+txlXcNvF7bVh7Kvay
yGv71BvWSpiWx4TP8ReWlw+bW+cifsYAZaJxHKLCBFMQOeTFTxNsxQ77dMhl
hbIGqXLLm96pxcIHjDXNbaBIOOe5bcxBD9zEJShlDBe+hHVyWtbZMuHdggx/
GzKgdqKWIK9qkk+LvPFZbTI7B6TGT1IcVcewZ3DOAnZVTgKa+2tojH3rW0C3
LBNhweNkNvDdR4W2uVuvavWu1E2hJm3e4GyNrnBmvWuL2l1OSPxNX4FkfBkl
uDs4Bi4ts850GQ5F3FxycZQ/5WLw2JghxjyDAkxlUBuVQQ2ybtt9UdkOrtBo
v40JLDLQq1VM2KdHc/lXSkdlITmtMAwTeS8Gyic7DAMikSSopghJmh/IKdVk
HBOYV8R+hWxEWBsEpn1WwNooZyS70wpTN5LGbEIJ8eFhBkUrGMfLC8hkO7nT
KJSDLDAKXflQ6m75FOlK4N54/Q/mhrcPs1m9ro65vBctN0BfMydEtt7XB+jY
IgcM3vhiNmU4riog9gGw0s5F0a/HhRWlYbOrklWXbQ1j5GVrUiDjGTRL+DGd
N+Pg062kj2GFpp1CzGXk5vto7c2bwfzdeimWfceq/sv90lBBapxLEy8HAPG1
RX/lA5zRhk8iiPE2L4u8ZCSBXwtHWz5Ftq+x/QjxlVVz59aL67HBCr5AW1xo
TZJI2Jsn+Gq/sVIvKTx5hnhT9C+sXdZxIbCPtsbOyCktc1zDvEZ3jCHEM4Ti
DlICPHwRRkuysIlDkMQuxNhz0XhPp5ynRGcdE6RXWlhNH+XDWu1ZzjtRTGVY
BONbbDvy7i6yBfZl9YjdUN/gs5Ype+R0YagPdw6pbN99zQ2qU6efCb3UfgvD
COaK3aQZUnlYty6w+/FfhIBb070DPIMjeBuZGDXh0BOCccJc7NX8bWhz3UAm
lfvCoO3ylcRyUpjXfj7Ib9BclAD6lz6nbUQvQ3qdxdZ5oX6n+EKi97F7Z+x9
s8rXZWvriz4e+f2WC45lDh6P2uswVy491z/5uqpJx5pFcd/2MGpZtLKez6E9
UPAjmadyAdViF+iewZwPj6JkThOiSvCtnceXPf2nhc57YaYARNKDCb0ue4eQ
xM8rzrPFv3R9CIEOHrctaXcfrWbXaPLWV7/kUlVPgQYlGSsEgCYAQ0xEZg15
hLdvRfyyxs11NyNj9K1mkQk7BDXeNxEoovzyb2gAvHEc2Ipzx9G8lKINzKn8
826oNRqGsYr3BUrnZkDFoGwFTLMAmOGQVhJOlasDABQyj4Y1I2Zb/9tMcqdG
XTv62csylMfENLJSjDeXqUVdmBbNRP5Fv0cQjOE3eNEM/5N6UtBnKeBLq3/W
AiiKR8ga4hGLBX9Ltp9dC+7nzUCftHVeB3O6xpFectCoFS1BVUeJL94ZRgxf
v2jXi5Bia5pgm4rAsgog/FRS17UnYMY7Dl/1dZR/XctksOY+50sccwZ28LjE
qbR0bBa4jpbLjhQBqLHPx0YikV4KA+j6I10UDZz3FRUdgIIYX748Ty+OkZJT
0PNE0mCPBlBp/aCIr+d8xg4+ceKE7bXMJbWQwet+bqpIctdxKrtIH9n8ZrSW
9Br1okHlqAP2hPhxdJj41fRyKCLLKMCZDqT7+itIIQ4WJvbw2bcR3pLdhvm6
pxkRQsccyqK9q1M01/NoRRIbTkViVnQ0t95bk0xzcLzX+K626GvN9woLLwaJ
/qhutvklacFNSXlHEy1eQyi+YP1KuSApJix/PrprltkATJ5yMmDrjqKY+uxc
/mFL8tuAYyI+DjQEfKswADLzEDzs0+2HB25R6PmdRktHmdO2JS9/2PZUMaB0
QYhG/aQYzOL22aIZSbA0f0NUWrasrJNGTaSqP0vSKLi8+i5HEKtk9J63YFT4
uXLE9pN1tkQrRFTQW0QR/yceeDuC9jegl2qmtErVDDrH08ECMqJSm2Esm4Gu
BCkXN1yw4r1gUDs4ySW3pF8bLhwz3XFvhH1cV2XxDNHUFS6O0et1s9Vst0mt
RemYM2nCIsuYazffP8ka2QFOjyycqVtj3L4TrEbeRkQsSWaEArAuSKpQNkSQ
zP49Conr1rt1XVT3otN2Lg72Tqa59NeqjMvIiqExU4Q8DuEts1FF63/ZL8Og
7YuwYDMugdXZIgLYZB/Ji0+l4GiNM0cecIHB36OLwbVhX9YUwB+uWj7x+sjb
8Jla3U1ZF3vyXclsjvFz/Zntm/zMx78A4Pel7mcS/V/f0Y7smka4tKf+W72d
diPmyEOVJ4y8RE/h0Yy68WEC8pIxpcNSWBiZBvmIR5HMveEOzBYkY61qqQYB
AJ8bbSbclUGc/0Yh/sLzxBdQ4wyS84EIsuR9f7E65ABGgP0Xecvqyij8C9T0
kj9Abp1uoWL6mXrAWABRsvQHK+Xya5a3rv5ADsoCtCLYzVERYB+BsY5xPQe3
Brv03u+9nhBc/6HpGTR6n0i5p+fJ0Gv/1EgtG1m/ZM3GMga6r2tdrCNNnoyx
gxL5CZ4ib+Sr9PcfrHsocI8b4s+cC7c/1ViCGl6igzsFJXVWjgvFzlzzQU9u
ea2czERqq9oGmBnx7b2GLSpswK8IBQ4k1MLh79VJFZ7kuXYAsm9t+LyfiPIl
oqT7VoCiBdfkYqi6DMCqnHT0nBKVJKfXqiMfgE+Ll0f2Aqy2SQMs1/a1/uNh
PrUvgZ5l1rr4QNkznLnzopWH9r7AtjgbFccEeiZDbS9aPzcpM1ueRi4I1FpB
QDaXCC27NfqKPZsjCWEmwTY3AhAXxHs0mz4R+UV1mUSANW+SETXuZSohq7Zx
DyrG589ERNwblLBx5bFImuady6VSGq1o1SnzSEqhOkSzg+0+NPBroPkMfshB
/xfHzmMbaWGEokHgVPk3qXRhgg0nXlteLqewEoz2jXsnAxWc9cDvEsI/jqX1
lPbUtGLH7ojn08kHn/0JMs+RbwPZRv6FmygO4Msv0vPQUlrHbtRIyrZhXfXG
HiWXabXtmMCZncoVAVIc45OxRuTL0iZibD4pJcQUpKYFE7FckVlOpcd6zKFV
S72Wp/6K/6y/NmXQ8lACt6SgfD1HvZQ61YahKzaK+R3V9a4y/fAGjyJC2d71
fz2H1XTssxUZ6z4n2GycA9fZQeIi0cjUGgrGUXZa38j9FB85brbHz+U/IVW4
1RB6kVWg39kNdRydK77qTKudRYUvAuGGTVHYgRAcW0UQT2LEeTuAXpStnQJ7
wxBaGro9EjeMzeZkm+Dz42LTHtQPkhemqNdFRooQEuuQIpKR3EqS6shcGHKd
Sr3KiltQJqVULDQqoxKWVQecjd4RHT7A4dK609qrTGHRt/qkzObx3E9DVgq4
Fk6TKaBgz8HaNXXaoUSl8ijb4hY1cVVBzkaeFusmV1+ALl1z2UW7tzC/GCtx
3OZPUvwAudTXeStD12abslP6agugfec7n9HePuO4AMt32Zp9ItZa26s0NgMi
z0bmIcbIn7DAsQSViS9JRv8j6enu5w8CCRrXwuHTG+/MjAYNmaIpwYxuNjoK
ZIBq8xp3ZPzHzTSajGoAavN9gh9TLJ/cdRhasl5lAPGKEcOyQktsDLfVvsl5
dgVOgXaX36Htdn2I8G4yL6xVVmYIvzKmXoKvLCtrk9jeZONWsae0NANFe3BH
G7ubbf9PaNqFFvTtqjLKtW1SroMdS7/+Kj1fUQKcXEzrNVENPmS5KuEEGMWe
P04sSAtcLJR2pHRY0I578HIP2YeYKIESVXBI1RQhIqWy1XGZli1+PNtU3Tyx
Wb8lvxQ4YxZ5FtOQBKRNj3sNX6AtH6K0g3XA8NeIq/EdV9HgKXGkgkAZBlPj
Qo1DH7RIUh1mbv1xwD17B7NdDMk21m4M4S5wU1BSEH1+6UnjHTGEnOJIfjBM
6gn0yMye2U2HRDXx8ka1AQ1o3DNameIfRXmihcJEdWHndN/QOX5A3qXqTGXo
yLYDIJBFDArQVv0NCAJzgr2t+aY1Msw4h03JG1WBisc2NF+FTfRNMoz4dhoY
CuOfk3Xbb8Qs4zjj8/Ym/FcvrLqxxy6gQfvN0VLtr345WF+LW8PexHKaPYjj
YNczGXemy2U1fhNrigpfXOqhpaOg9qapntQEBOsOp4ZNde3bs227dHk1U2Ri
jDBM4Nv2uILgtQo6m84IvTRpR7auk7gn2fEDewYvMIixy5c6u8igzU6NUg0r
aDZzKw8UziMN5AhZPqlxqhJb92ybSV2HSM9SufEozsQcHrpPKY55x+UtJiOk
J30KqTEK//jGPHNsqGZnh1jwyLpqY2E5IGRusjAm7eHIVOAfwcFyXExZXp39
fnrA9YiEKh3C2ZY/rNefnOCcAIuRdztqzRcqRrRwcnj11xcTVdi5GeSJP6VP
6ftQ5SETc3S5B5gP87xvIDIk4tCm5/eDpjElNRq5u5lU5jd0GfuyrgEXGZpy
XG2XM7BRQfYJOWKMLytCIcj6/wlrxlHHsus6TjPpr7C2GpNE3dxW5RaAvLOG
U2hqdT7NBW92sQmE/PImj4wPzx2Kxjh3jGQr/Ju46yX7pp2GwPJYetSN1Gk5
hsrX/6mH0S7IVX6D3OK7nlSONkxpbDhe+BsKWBESJTjVeMWXyNG/X8ImXUda
rvHYWJtwoCjV4d3GXlSeCt1aHLzuv0xChll3LBPcl6fg2DcN9z9HBBTyJrZx
R2Gcona99tg3NpYsd4G1EQ+b/hIJPUaF1oQBGSLXpsTKP3CZDO55aSXz6XIM
eQ0ymUDuESGVHOWNNQ0o1FQnmX7SgE3vaGRV6iuXT3CXWKiQeAHXjIrIYTJJ
zkgddYHqA1HbKzlOtNx/qpjsvm09DjvcagbUxVNfkts8UV8gdHf2JzpWpkkm
yw0K9tjUK7ucLlxLIjYQc+XG4dwPcAb1Li19EIbTqGlN/Y7ShdGTBpRaST3/
t85lVI3/gQZ9W1xB04+iBX19EfmhE597HIT93b2l0KNiJTXU7OyEYJMGDdCP
3GWEb8VUDdWRLb8U/BoAvvRcIi7sH4b/TNDlLZ15Yol4Ry+WLe6JxeirkgCv
98EKFB2szYu5kaV2r1thN0SrdqQcOCkJv5XCVaed/nvjqMpSLz3A7Z3vH5hE
KYgZaI/TQ4Rr7HZH5JnzrBpG8gUnMzppi/c/jugRaaKnoxEUI6U/sbC5ZePN
yWX1xOrYPZKQ2BBzYWMg2XriLqrNMHirrPx0Q4IpGUqihn8xgjBAm2F7llaN
VMSyTdwqgnu+OCFi/6f7+T/xMH/KipZeSwghujbk6dPrAyHzpCFdDVvSgAUh
jqzBsSg2Cip8PwJnObLuW+xYBFpQ5biW4c8tk+7+rlbvcrUYodYx/kwIVAPQ
i/ks6Zgxi8ezya+MBFpjEz47++b+b3akVynOvED1hEaGejfZhCvLhI/WR3Q3
dYFj0qLMI0ruQ/gFF/VvDAIhM07nXW2ZmPVJvsapvFPkLpS2vATFDoBHE0kL
oERpABmbwLau/dFRydMtLOa7c78p8IspW4DGoBq47yb3oFJJexk/VKP+/g+o
kUDbz34csaFXZ+My8plULNnW50wZhpQ2n8qku72LkD09vg/QKKj7kI0Nrfiu
+mLMbRdysdDQpIoKJA853N+f2nj6AJ7gpSBwfVgul18VMAMAabD/BEBykOk9
umJnQ3uoNU2OcIzKCVr7VqlDtmi67GEh9n1P5iJDSeC/1+LegBtYQXMm3e+e
ChFcljiMzHqxmgBLOPPi+b5LlrOdrGn2BiwUlMqftKS3zlrDwCp38WzPjBUN
ucFVxZ7RSFTGzfzKpCF23X4v68La3OnMw3cgVRy8OJZL5GUA9/as6pPDJUZT
VsALxqhEiEoF14joCWEJrVN84KxUuq/1T2hKdRqXGFQQ1a56HRW15kRsrk9h
ZnzmbRtJZV5zZop8kKoOadnwkwr91bU01+GancrcdVBuDjpgYO2+50zg6akZ
6ZA5OCd2//olYg5Xka0Tzh+QOMvcgkWXKg0X6shrgGnc4DkoL7BpqulunoZg
8zpdG+PwfjGynBZ/UhCgljD5v149CfSsycWrEFOkTqJWzC9uDkvXn4W21DmM
SEkCLFHHnOrSNCPpjpSxoDmyNTq7MmAI78EHhpgRJPjM9Y23afeTh5nY5OCg
2CRP4c6zffALW8iep6pL7PCJwzxRRhK7WryeOeRtkSBHs3WM3+9a21MDEQtQ
e240Kw9+2A3Yb5ApqPzETHhDqy2nL33c1qzqaPZ/fvuurx7rkXVFsuUZVbpB
qdy7N6zjzbCqaEgsmaKixoIFpqhF0BO8fsmU7OAW4yIl9pAwtvmzEWhtloVb
+IqimSr8QxK896zs/ZK4Edt6qORCQ22K7cI23bAsgUktFDQhXkiudaqy4ZpJ
FembGi+8l7yklEN0CkUFGd4FmhjvI/dUrdzXb1vTA4QvQfmeB1kuEcYSVj3F
1ASA24SqTKB7Pmv8amgF4BHjtRLWtgL4UFh45Wb6hA+yzUmny9n6o3F9aA+O
YHPKTxfW957NGG2MeG2Xkxw037QGzoDXHAnb89TqKgbnUWTUTKf9BhacPH9A
QWhZGdIwUSFs1ik6pIIM1yOrdaramVumAja6b/e30UpHh5CGxMtUSGnchsc1
TpcoRqYM75mkOi++AjA/V4fy+lX07xA/2dVkhol6+tbwOg7ldFMDcGveBu/+
M5yYhJ6BkaStIXsKevN9jTsMRmZJY4832x6xCOCaOJ/tktZ3Sd6UPmNJfSyJ
ICRitwCfuUEYAYq9V9UPjjHU7LBmK2SXzCWwCGNgC2dUUpmU2N7kVCIStxFA
JdpgSGtindJDcIkGI1lobY+R/LFbQ39XuuNr5k1wZ7oKo8tU48Jq3HLWXuCo
RVjml2qEwVkDObjUzdaHduF1SsL8WwGlrmrEVF05PYLkBMVk9fmS2k5LRoyA
stGhXybbN4ZPV2qbO5Y+PvNygmFRYrbrOkH/JwLnOFjiuJ7FHqX+EqNTU2dz
PIg+ZUioL5cjXag7DEr4IVcIkT5UJsT/Wdy5mXegNrfAFvok35wHGqbh7PEA
kG/u2HrEp4R+7hb6DLWT3HzmP+rt5sfa0p4pNIOosLj0sdtnTVCEeOT14hic
xkH7vvIfiRsx8iAtnmQkQKqqJ8rPw3LGPGuj8VisgSwMsV0AkiLGG/J89hAX
TrWS5KkFqVCMJCZTYetkqtsw/RBfIDh1BNsaksMC5st7N1zxxzE9k2DVFVLW
zsjFuxg05LjM8gXr+jhV72P6Z/VRdH9Ke9xjXCXpinCtnzG2v7gBjMwwIWfZ
P3OiLOsfLpX61ABAUtD/vHRAOhOPQ89ehDhEyk+NUMtkb31BPhxj/Vjc2Il8
teXpYyK4fn9D0lpX4JvFIIbaHP8lHqnMZggsLFhs+rbhirYuuOyhwaHPhkMZ
QzbO1u50aOvb094ivoRHLxPCm9iIlncr58Y6hDHyXSgQL53dXLyu7NLJd96q
3NoFzg8VckZdJn1ZVg3cz05dmeDL5VqLcFXmJA5BBi9WxhbC5ZnVkuHKXGiF
kHgRbYHPsoCIC6NTbjgea6OWJf/xj4GMP6yMbL/IIc452LXQC1swb4n9Yq6d
mAHInAZDCWRlUvEWvnLJ3jtd2MSjiwb5zZsNhaFkqAhppcHwnTBUWhPmsQCy
KkvhAot1QkUs1Gnl6IP06fem7BIseUXAMF83Mq03zEndPNbRwBPXoX/ty5F4
Kt0Xab2wIZsh4KcSXnigvtp4VDwtT2F5gm6BYa1tCMVJJ4rE5VVa4hIqyq5n
fsGJvv/ILOiNwG1y4imZoY2Dm54tjr84+3NanKlfiarflUkIy44MqfBbExt5
iS81MUu+Z9oSkBf5/iXqewv+M064yjT2kYS0h0qXFYpT80oeuLAxYQFwiOhB
9pbd7bGkEsOYokfrPWlJY10FcPVaSlmu3Ueto33C3+haAIZ1J83J5vhrovTh
MIIuKLSInwYy5LK4cQMiqVCs1k5ZlNQMHDRwXtcUrJUHObQ97bxW9D5nRXaQ
TdONmqB7qpoAtN0SSs9V6lc72NSh5BpNrB9nIK3wvSVi6EwMokAzB+Ikb2iH
YWL/gbeHHtqu+fTbcIsTPMDj+HgoxRUrHZMCbOEG/zSo5JFSWBajslb9xNg3
M8cKthGZu+zLBPy4yBZlZdvQwij3AqWOd/AUDS/6wvTuLanDSoSDOPh8rE36
yc04DxlMVe1aiVrbSyA1T0WT35ExRSykixaZaYx8OABskwuOtbTvTGu0CpLW
pXJ2sLr24M4hzGKrHgB9y+el0nK61oTLa2n5UXH7MSPAZfqKYbmmeGZbFCPE
6eW2kT8wgv7RHXPPzbsrDC2ahrwKGkxTQYLyf+bdC2EGZeftC5VJsTPZ9IpU
Ai9tzotXJeqTgGyoHRhqzzMFHoDDs+sNuZ4yflV4e77B3AAXlMU0gywg/cui
dit/6iD25gm/pGrcgtr5si9i1Y1whLUd59/xFEaRVH6kTjpcS0eU511fjEyt
ptA9SZJV79XLNL4UghnyshpzVRI4eUwOL0HGqY9EMlYRKhBr6FAqLuNs5zH/
v2Dp0SzPSBoPYrst3X6pt9ednmTrTZ4S/mvWCTplKmnGct1Ksm4vKd5d1ZmQ
lsMsClaceM1LJwHAHxtIti680lmOneD5ylkLU+qOH8GoidOZozB3mztxtIoW
9+p0z2rf8CXdtEu44dbfYdgtt9cQ+m647tPVYFppcJHxukzCIi1p/YnShCqZ
HT98weRCcyVPfIf6PBoBGEuwrw0Xwq6UKYCkuDA3zjGyKvm0a2wyf9o765hM
jODLQjTeVVcGkiZmyxLBokJRhk2WejaHEJAd8Zq2KC2+FbWVJ3/0A0aqylWy
dD1OgbMebbbmdV+5NtEJimZYxGlky2IpAE/g2J4/02nN1jUqRRKxPBhZOaSu
9DtAUpa9JiTCFRs5lUdWCq4Kik8bU0xDv3GaaL1ZPvfFoaFUvb94eFdP0Egr
8q6UnYfR54kUriaAHRqpgx/JPEFhDgoc9gCg7c7FrY2LhNJ0vnG64Lpuodo3
PE3D6HcI2sjXUB5t1n+zjkdm8tx9WS1kZvnbLIVZqVgyzUnWEDa5GXPmlXPJ
elY3vWI6SJ01/UoVf4Dlrf2Ir8FNYBXWkZmDkpn0bKoawoUwAJCVCR14hGrd
Dj6MBmqOPZoWI8yDdvegq9aPW3wHzq+T89XM3Vfcn5dBFtJIl01sqM4gAqjf
EP5WmHAX8YeNHrJ4m7jxO0WoCYID+PJsSpeqEZ0bk3wbBsB+UQwxgAux4iEa
VXzCxTBsyYnGRvSFlVz11SjihbbWrxkRoROFrDVI7nLMNJTj14yfTaWcfhCs
j3yQKOhNqQ2Fve8KWnPEbQ0i0h6q3D1FQeOGd7idkdN7OYCBnTJtTn42zzj1
PniR1NE9blm5UH9XiIhv6ghkHo2ZuxA9/gwqEbdH1H0EhyU3UNvHq6FfeBZn
1hB+bbDMkN73/P3aa5/cPSiWu0bRKIVVefyNoP73a55c8dIr1C4be509Zo7B
xEKUmltiZBbRp2SFGjExyT6Jx8S9VwNXyAKeJeF8FFJO6RSsSuKGMWojvJ4c
C1qTsc4Gq97AIPhDhn8tSB3AGFM/a1q0w5EKT5p/NMsmTdVCzNm2+b7xHy7a
qXAfMj+TdsKomf5qopaQI7MXqxiIv+rfh473q8INvULAvx5iRWBlO0XX++WL
RXitnXAOgf8EctME4ZXBDmwl95GqXi+2UiImJw62ZelkA8MqpChUI0OjlhAQ
p49gOwSIwhxXeIYV3/PlXkXMk+BAk6Av9ZdtyoUeyzEo7oDVstcd1BNuB8Sh
NlKZII6rm58cTbJmlLDEN8jh8ZlnBWrzjdhDHru7EHbz3OgkeOEt6lYZySku
lMRQlij9smM4GM8PGAyclUQPmUERn3fcC0zqQHDSN+6zjw6RaY7y/jB/5M5A
98hMot/Jf088HxLPrKU2u7vm+LVrZV0gq8tkbIWz2rhuRZKErOwEQTCLP6ZB
aV+W+jJcnEDP27OGUTQ3IOE/9GvGViZvoyq+lv3zkqI//ocZp64z/yGlZYmf
OCe0ZGup1rfNkiu/ZPs56RlumM4GFyOzNEHJM21lO7hmzT3SfRA3xwIIIaaL
Q5su9b8HzMCp/R8Tgg/f7pwRZocgGklvvxPQiPbFT6tmf+3uplAb8Jn2bVYV
Z7WA4eHJg74BY5VPbiPnyE/V2OnM3I6XDDYT3GXoMl4aTbyn6mMR5nKQ1bI+
YI9dOq0/bzBGm3yqWhxq/ICKe3t+b3LpGNuSkNedr4HfPjsH/08WvQ2fA+Kx
xWzVZzoWZYjtiidLlN87vdoGyJsaBCnP5sV/mCihV25XLTd5/ci7qUfnPvHd
u4j2Fi4HZkZyKNFXRXLeBFj2C5pehaDCBMhHH55AjHkJznU7OfLA5o3OG4zu
s+zoty+2sND0i3JyTe6OeoWKUHEegLdTYOrMaOSonPY2YnxcIbxWweJbtUHj
LK4UIY68vEXyZCwN+2t8QafztsClKISHzb8TFFrS80mGgIgZyNenTMh/TtRP
mNAf38nGnV8afIfaI410Xj8KY+iFQMeUHDaNhXOWwQ5K2T5SI3Rrdfo/N9ki
j6bJi+diLie5zdr9nVAHSRGYeuqPWftHv6NHBCn+thB0TL1RfDsw2PiZzwaz
e/Hm9AU9+64svGMa7t3kEJ6yZFBV6Vm8up0HmdJYIS4osLIDeV/F5B1A7y9M
l/GNvCoXZuHqGinHA+u5PY8G+iQ6rzGKgQU4RZGUvlC4SuK8Sv4s3PWz8khp
Djp5QsFw4NEi95Oqpv5rr0gMRXBrQ3KOtXBssexgFkJPV/YKklFY5ikkmBZn
dovlqRSVbsJZ1B3b0FqbD+NXWZ0itmuvsed1Hwh8jykL2eB5cL0BLOLnSmqj
vmDVVcenhaNvBJlGWi6lusrE4OM3ZPRfJDH/cG23rqe+/A3EPmy/M4LPom3R
OMf+IKKke8sJSJjmG4CAMOG4rdQj0ddcWqfn4BngLvU8b92vER0yeneeX/nd
6tZonyctT7g3O2x7zHnZJ6fJFo5uO0Voa95driaBPODwT4bWMoMe8fHm5h7c
Ob5BBWkGUQkAQbGE7Li7Y8zIYR0zKr+Y7xIFs3SlT0E/9a1LZc+NvLnrZv8F
Wg5VRg1SUIRgz6NA+PFMYoCyBOaauMVbZu461+noRFB+xZAHGGuXgE6FGKw5
QVVS04P8bqafw631jqJrg5WELKA41NvFt4ab8e42xq9ba3UfU9iSkpLaZEJn
MgrOH7jUWW91gLEDyEgeYGtvmZE49Jo2ucfT0xge9F/XAp8kv99YtSKq49d7
U/RYY9Qw+PPT/W99c6OWLyI08LWGC/LFWZP+clBCorFa5s/Pte/hsw/B4nNH
xmAifVD4Mflb+WYEIZEXjW3unww5eVxAB8HO28edSlm0r+9GQjw9kXr9TxqO
UXbELKZr7DlVKwKcn8vW7dnxoeDXXhEwRtO0AynAI+KNVtCtoqeNCbOGfxES
+DgnNVAy0eKF0b7WBXGOUqaGQt8rgPrNxQh+0kcGwBTIIW0khqgbGaSr23Rl
EdmxBm70fLUrjmTdE/QYeIjDRznH1wOMs8IXCcBLVvV56EvugZGDSUjfMqAw
qGb50idsOX2eh551nA3MoGeTF0PPEZ6Ps3N+T0MCFz6jFFdiMBa0G0DVlqhM
0KRtmbDmakkZk53hwEG4RSbvEVt0DhgtzG8U/XS+hML2tajHCOsvAazkd7qC
TC9lF1A22xIs0rlXKJbAdokzMU7aU079FF4/2H0IfKjXW2F/pVzfwTBMVBgc
J1580kLl+h7TtGnexlngXPKuXS/vaBjKAtEWZPVBRMhZ83aRxjjOhtezW5SH
gasLM57wsnm/gEboB30ZkL6MXeHudeMKchPhNajlljXVwrfOm/MnucZrgAcG
2zU1Lw6mW6EMErWGJ13HCKfWKLf5Gd6y7zWxnOlj3YYhxoYkh7oVVGbyAJUG
r8EGwINuL5tj2zUoV8GIYvWCB9pLm3JrNPH/hQT+PFEaof0A5uk9fbchTNcu
/dYZDk+aJA8NbQDKrANGi30esY/6iA3A3hxq69r3ZnkySuIJ4OdzT7k2pRv8
niI0i+ytU3HnbOjlIbUdafuD6CG6THizgASy6IrRHzKrhAYaMu2qMaHzyB+/
X5qjZFu7x54tV5VtRv555jVPSPWydlBfmktAjfcUgWfurYZfgmGuL/vtTl+j
UZQRg5XFbfEUKBxQcDoUEhu76G1IPtKUaRNdVVT2jr8I7rUy2bbcYTm5h4WM
1HlDxWqpi9E1e7CuCaZBMT46Mc1vCSqVXfMN/+sltjk9PPl4agcrBECaqHpO
NGqTG/70vNQsf5l3vCEIEQp43QjU7sg/E3vSRHJSwgJfaCM4BXkGgJKcHsQl
CNerd9+5WcycMbq+bQMHH/vX2QFuLizVJ2zJXDEnrywpTT2xyH7JaG+wu2HR
6MkkQ+Y0ILihaN5IIoGZvRoLIgZm/2bLOYzz07s5NDNNwyeNhg43QR7oVd7/
t0n7A3Ukd2ldvQXeBosl0KQdoUTBNqDTe7vlKasYDhEurtKvJ8M68l67Lg8s
flKYlmaXgObuO9eKWMFdWoBW8GIYi2pc3ZhFljORwNrht3gLlGBJ8fkgfMhh
GFO0U4/giC0WVAucDjFyJah5a/6sw6KH/PHyQuuWTPOdRs2/Myjx6cx4zZJv
vErRAR10XrjVmjHZzQp0mRG240/PKgBmzhquDCXtDG+7wzKnU9/YTtTuEtDm
yF+o0zp3rTm/CS1iOOnHP5ByqbhkOIezFDVcYQbWev1496ptpwSnnYNOC75L
0Zg2TCw2CK2YgimopijChWZqMJbIMSmaUmzY0gbC0/qofVihxchlkqftcHhp
aiZ4oXfH26ir7dMNI99glkamXvT/4f0X21Y0CWH3HG3jPTBcGEsDPO25pkaz
1RnvSDbHVGWQz9F9sc6KLgSTvcH3+7KdsbsJCdZl5XsMbg61afQSGLcqhCIi
QsvH3qvU9cVSParyjF4p50uSk0MUZLU5arA8OXE5yBH+t+e2SBjnl8ZdmdZP
XvQnWt8Z4o/4l2tDQvEoEzPEw6MzsFArPtvEX4wuMHAwepsnkW05XC5ea9cB
QKryiQnwnVSTOypEu1g1QtdTKnKdf/yMG5o/aSqm7s0A7aHatUPXWx51md6+
NP97NYWMPRvrliq+l/fUdgA6oLsunn7ODD5R7b7wYxdH4WKY0dx2JQmp+FcE
bkjVd6yO7XkKnDtA2k4ZgAAJCRKmMRBI0X79v1ACagX1X0rCEWW8fc0xyOZY
9+LHQQ7Mc7nvxnBgZ9T31lGl2Dc7n+S0EovNjIwcT3r8u66ppC9XoggdhHj3
kvu2WWCs20pHVMt6oiMhoYJyJYWXXiG+ynbwFgBAxz8yZOWJhaDI3mORl88H
5ZZm55PR4XqkkytIpak7gPYIuhZu8jGM6fHbfjt5V1ArgxwmziUSsrc9ZAXF
retkeTaPd/IKlDxX5bXyFs7ARnw6MLfkyAE6ZMjHBW6CuO98FF2Atpa6Q/2f
X7RfRRHtVlt9CddxWkKJsCnQaCo9CeL4zvizAtr2NgbVcPywn7Fbt5o9wedZ
KONpv/vof8BO2d/q4JusH7se/qO30akhpG94V6gnTeRNnvcNRd56/hTfkByx
2JiWlKnRfq2GYsDvPLuegtN85McAK5FVqb94yNEjiexoriI8AzuuNvQuSily
vLiTLusYSO5yiCtD6FfUxEL8iACJuMX9xYaOkEoqL0SML0l69M7jjp650Ijv
+evhyGKKp3m2DBQ4qxNV/28p2jCMiB083f9SvMNFiNC7IbvHtNZFBNLJ7Jyi
ztUFEPtWXVZX5KhObNBnuBUJ6byHDZgUaWujuKTg+Q0ZUFKADP8x5Hx/eIQk
6Pf2iLDLExIycvJHsW8Fy51PPTaliejeVSGqJ2eARLg6j8Q16TpzM2Ts4pEX
YshYVHCxxcf76mezl8h/BhnoddpVQ8fgzwsAPQRI0shclnN/gaefT5n5YEt4
cLzfz6BQNcpKW0LcDm+S/ZkcWxv2bgezoQzHivyz2FqBO8cA38GBl+MFkLPR
dUNtV3/+lm6RWdo7nrfF6+zOYeoJre7l0tYZtkRE3g6Z4Vu1IQccq+7toWF7
HgslCdxKNjo0esmAiYS/JoicvoLhAH4VyzjLNcxiuWHK7yCev91pLSFt0wr4
i6wpJ9rHu3AgHzsEec4cFv+GxDouCDN8dhdOfA2UkEw1CvQtuh+fRwVVHQoU
2SO9e2IZZJoOKjgF9akyGXoJ9k1aWz4tPbiqDxS9AOl6ebdAY2UtWYX/1RH3
AeIgzvNPHbKH8sYQBo2V8u+UbbsBB1oWNddoTLRwIbeh+iSsnON7fLrO5FPP
lOleWjGCsGYfo37rxXh7r2cod2dZ1+93bmIibaBsoaxy8HkuKM/HhU5rnXjU
VJdiRuwOzLPx6r2aMmZQcb8h0yPdQOgyXX63Gw47OnyXRcKN16KP3GfjXKoO
L4KDgx2CuiJt4yU9+jlhNEaj4/UtUF7giO79aXgbqBKNy5iLRf+CgyLtviGZ
ri1+oOOa8g8Q/ZEoibkZGsx1P4F0HVC/EG4f4zfgheHKqjT/rPDbg/x3R5RD
omomZqhd1N3ZxEerLBpR5uoeDD4hArOu78QFd0Jbn6cckT2lCC2Ij9NG7Nv1
e1d99PIS1yCHqNLyzIhR0yRP+9lo5MsF+MbwZNk2uCTtQy+xrgHHN1PBmFP1
zgYyp9FrpLHQKg5kSTXxU9j4dgfFcP/JG3sWAdFlqWBaZqHJL+C3tXYc8bR0
ihYPMw5J6YBkOIbud+gCAZktALCX8xgjNT60AlSNgZE6w2mBsjYSdfGayi+f
vjmvh38JdVXI9iNBpL2qugHBZTu6C/Lw/vC+Cg5f8B5qqZ6N1zDjpY5vNaV8
MAYVjwiYfu6ArLrRMPk9IJCbV58BQT63orHslenNZBwZiTq5wXIxu5ykykpl
0QNZbmD8E38sFUFEf9NL6+82S+5H9z+88EQyiOVmCPmdAXp/D+1mOqnuLEr2
efGF37yJyegK9FaJGyF6637Mrpq6P3jftsY3dodQURkFf1USnOTg61ZjM+Zs
6HdU+xUTJMjlWAidHK+yLoOPu3l98kbkhufvINWKZmc1PzTWLsrZZFWdTNSC
TIeO6MGqNdETDOpJKGxmS9j3kL0/XMsuB3iPdwgV3QGXCtp1zqmwmXIRLlNl
fRQtMRpjL0VRxN5y2U8aaNFcqNUezIxIQjHBad64pEmFHsLAWmWVEi8+Skow
B6GlIXCKK8+j4MLCSMrD0HnnBrSl4NKZAOwwcuDaTQ5o6Po/XPtt88vao0q+
B6E9fmhDZ8PpVNZ0bqCP2uSTM7bTeA9RhrESHBMttpU+KuhJewPbtzRY/pf3
jlkmjxxwXGl5+vosyxj5M3JC/vHB1+4xyQ6IQkP3Rquicj4MYJ/A9wat5rZu
+40u03Rx+Hyq5yeRjlRk+hM0Vi6xJMQiNuLozM0vk5TsoafOYgAfc+y5fjBh
jTeDQHjIgoDu8WfXgu0mS2etSUZysFVpRvqI9n7wKbkHgNvWA69dbpzOsfkN
ORFmazp5mfHn08on+yZMG4TOpcXOXLuu0084fMMKaC3Oj5045sxkO44W0f8V
yc+X16qQ38KR4Hy7et+o2j+npnHv5HJvzb8tqrhJ1XinQ5ZvQLA1dKc2jpK0
Arw+ZXawGRLP3GDkxN1gDRn9i0N0U0zDpm4iIWZy7UftAgv7Z97tR6S3RdWk
WPzYdlbSxeawtCtwpaQqyn3kfb5wnXfBtPzUfURqc2HVqgg7Y4rCkFN+RJVY
zjmfSIhwXfSM8BNwkE/4iyNzhreTmhpZd+WGyBDZrwrQ4vmZ58Uqa0DDCNqZ
Cx4vuQY/UHu/gYHzNInKcppdPGtT+CLGpMuWkJCtwe2O+euMwdZBX0Obno/w
gWApewpK6OlKGS3GL6Ae1VtLXtdUDc4ZQ6M9YLwnuUHBh1QkT3sWMtlhMCuG
Z/dDfiVR6j9btYueA5kpidOJhDda7Fr24fuXeb7UBgJLB4njjuHRGo6sNCSX
jS9oIqRmTmwu8EiCsAz5laKWJIiAzzZ0yW4K0Fk+kf83y0N6pigpb15YgMxA
s4o1BtqiTM1hc6nWTnL5BHB0ZH8Sf03w5UxsOIjJLGpDj9IT/ax7xNf7EtR0
txAdIEyqFv6QXsIYmOyGJdK02M6zTgxMfeIVbKooqVJ/0Kw7LhVzi5nL944L
ZukTOQi1y9+89TSyBIE6imS7Ua8ln+ddVZ6AVRRjRJNPnMC//LofOorA0wZw
rGnmG1BuxgdpHpnSP5oRsuxKHvbhONBEe8eEU1rP18DB5eA7hO4QJkC8Dg34
gSC+WMrwnj5lBxwHqo2ojq/ox15utepgdO9T26HMujbKhXp56tBhkffF2h+2
QR0g6Axpc46f9pxbbXQRN+XTc2Gi4k2lcbPLL8mmWzs/41cGKqWvyq9yTSTy
wyzpxLlOCRwDi1GWwcEA387fAP0x+c4Lj1Rv74xvlJBJaC6SIWQ7EQ69OL15
8bpSTS41EEZc0xcRGcUTGiGHq0n1vX4OqI+G+ukZhXLhZiTMfErrxWQeU7Vw
913MVAsWu7rGJtO9X9BpD111b+ks5tSXc3s9YlAeBRiFLc7+CcSsyUxOd9AK
fFtmDLf6rpk0DSMGSFz1DED/edvX8EA4bm8qucj5L74Otyc1P4LX7AfN9QMo
viiNL5N+aI+f9OW0fg0Q2JU8Ufl8xQdHWjoEG8YTEQyxJNpUS8aO3wv0X2GO
MhiDE4N+tK3BDgU8eG+9zbBR9JVoCcEl3Y70AVPZisvY2luvww4gnosHu6qt
qCjs4psj5VmTvyI5zDQr60akU62ygISQntQ28EwuFAFWb82lw7DE77zepMsL
6Yn3fDzJG8PB5i0FiJaeNOBqlT/UAeicZphaf9TQJgTLxFQYvCFUdAc+p/nH
3Hpq+1TBwgdVzbHHIVhByO6JTxzmOjJGsa3Se4zf1LN/V7Yc2yy4Nh6Ig00I
qoAr8rxLEV3Ge7ZFjblEbHVWswkePpKrcKVBrvgCZZkE0lAaEQ/NvLnGIKaI
EQ3MFMks9JEKaAb6MfHvl8kiwgv6JHVYA3Ni+ZGz4MEoG2iu1v4X1B0s71mm
4txgWpwRR5qybfzMqPA3aYZVQBUqYOhFPAINujpTj8xUT0wcR5bypE5fk21H
/rqsMIycXUUfGO3Pr/SBCVmVL542E3KdDzMaxpovsVelmgFAj1vwu1xpz/mc
SpfAXyP1njo1znMcNCYnI9gvbkE9LWxEQq/udrErSHVGsIHQ4yl1z6affmFY
srHxRhNX4bUr+/0S2UMUlS1C2BYOjpokEOF4jfQPCrm1lEnX7m1nDgTurS2m
GD+PxVYa12bZYrh7wuPA2JbC8wR1nH+Q3ISZHE8GpgnlONKsWzcwjGa3Faeh
hpwlh+ZvHAv5W3Jwlwymh7hR4YxxA+N//Sp6+8K6TA63Hy03k8bYY0sIPFJ9
o7BBfzwaBkKGjMG1taimHXloLZJhhkvnJafbXcW4kxb0nqkBH5+Pg2gHMvKS
/xP5PoXuA+FP1+j3OQn6cShmqVWLHC5qMgbSJL/hZVoUPZuDe+6R+LkhlS40
Qd5gEsF59nWC8tmn7pHcsT/84tm2saRh8rlEH3v6aWawSF1olxZhwrGUAS3m
au9059mhwv6kV7LvO8dktTF7ZDOEYTNOndat1ySV9aNLZnVx1u0VFbgRArAQ
wO6+a4Kdn9T3HTCUkyKMfw4GeO//yePyQIukTd2WlPpekej6LBCtEilN+yLF
2G57AWvf5BbSQ89xXElq743Af55KPKseAMszXzsruCCsxIal9u1kBao2TMe1
dnvYpV4a8+Bbuq1m66zH2Ub/hpE3mgoR99EDvB502NMTBvAjL0s30/cAXJXC
JSuNY9R38Jn8dgoJlldaNRpnBEK5FaLeG65lMyctWfeEQTll8RpQRr8tlFPc
aWxcH6QKE1r2fx8CcoHLqkWN9USOO8Ag0A7FlzU//FIj41m2ErjkLmXKyeJX
Mc3I2iS/Mmcj0j61p7PxBjVMtxFaR1Se8Goz/JKfiWNIffvzfkkgzjBPjjL5
yBS8iOunj0fKasYtZMikbaLxpX0RO+OgjT+19kPOhsMUmHtej/slIrVKqZ8I
hYo8JwvTXk7hPJ8iYFP9ce9grf7wMoxjHEP1FiVkWymMrk+RqsNWWLu16Cye
6puHhCat0poXoG8Pr2E11JioGcBM0QNL1PZ2RIstBNQLKxP+pLfyjSlzQeW5
LZDxFchDMbq8yA86gs8fOfKh9Dyv2eAs45Rcw5TGlWVmSShl1cgr8hCtFQOs
pV8JKzGhRE/HvLGyW1btmRmpQodzU83LgLkLOblVrEApsulF726VaihnWhOD
SWT/iPVYDbk7wYx0IZaYBF4z8XJZ90Dkp0eN3ny3DSZNYAQlyNa+cxRs3J1k
M6O7zaIj3+lT/Y0L5nzavis3Aj+JjuVSGfuiQnC3gif4ZT8qCGZ7pjVuJ4Tw
4hlB8lkT/BPUKsw470Gj1+JBZ07PPJkqYGyPPWyUQqDep/MtnA2iVhZPNvjh
Ieock1ZR+pJaSL6OY5vgEBEzzNAyFnomzXB/v2n7AaXVGRQlq3Poxxo5eJ7o
U+RHu4r/teuz7Vf7ZR+0TnOQwR4bV8IHvA5ncw1NYdJp4IgcvIhZPm3PFn6A
y4xjRrxClaGLR6+lPeUu7dvlSRuTsT1Bz3r3TOWwhqCUEQVUBWFWmgQ34tbQ
ySN4/6Wc7+f8hFqj0puQRm1PnzkvOVSSpYzVORAs5zIG1WCp9UPNiVvKGAzO
kxgjFU9Vh62CBVpUp7IgyP52FmgS25nGnhPFiaQes4Y5osDA/k2fShzLAgur
pOo9R0/pf71GCr+qL+HhJEVw3gD+hg/vETjcn1cPxd9WX2oph0tcDi+JtaRI
uwqetRtJWogvD/LJacghWzJGi6PwNA0drnGyRzu8a7tVUwjlL+CRe7W1SBBK
W+7LLI+YxAjKB+3W9o1YGIlS6ZRNwE6J1lRk0Y2mz01Fac54/P/hJbuifzaz
rFtFQgFIKsFLz2Nam9/3SzVkjTT3N3Cej4wejer9lesPMMSYMU8Fhck6BkQx
DGBKeDtCq1WCVjH986lCupgBnNzbdo3/KC0B627RJ+7IucLpbuvQN2IheZTj
YXLbbYpkdvpqBQRKbfe6b7QZ5vHwI/Qo01v0G3avh4YumRdgVqd469F+LBvN
LzWICjozWKtWG1gKedNSHkp19JVbon6RE9JLFE1xyO5tbblqMXOy7gElDXaV
zzBReFvGa/c+nHBPZD0S+H7xo6lJNGwtohlMDNZUmY3xUsClZPyvCQOn5+lZ
MTAYxP8S//6GMGmGJNCNWEMUJphgzqYL3A081BJlzfqMag1nIOhMxSPDJAiC
WptAn3k1SP4dKbgWm2oHyDHCHUhfLl9kwhCu4CcEEeGlYsvZL/ngEvgmflfF
DP+hBDmudrveLxrCWLwvxXdrc3jiySlsX9k6bH+wXyS7AGGNMC/u2FANrzYS
H9FYzgGz+yPuLlB2zV8lbR+jRZ/mFdJhTKwTsbReHxXzxYLchoF/ypqJrpLu
pgeSC+arC15kaL4HIGB6F/nQC1lg3YokNZJjNVAxSw6QTY2YDXgITnT2Mler
+N9Xhgt3uI5mkgQXiJBdacb7A5H2XpfYAx+BgedTvnQ1O7vykK+499ZSABfL
P/whX1rhCdsJuueQnPDnBiRfX2Uwi9qXrM3Ru3UNGBx8ZIGg+i5eqtR9xPO4
nfzbsTPwoY9kYpO165eF3cDIXlNWLBdFOD/J2d5mDN1Y8PDow6EJS6LXq/Lc
uUnf37sHNJK1mITDm3kX2RtO02IaPfnhWCoZi7bYmCc3uZ8151REJTkKOcbM
RYSp00aR3CURjhBRTU2kG2hDQWccSiFgI3CDiCwhUea/2IH7FY8aOs1k4Ucn
JHy829iAlr39I2wPp6vBLMKicoHq3LDkyArkPS44YtPvMeKfj7cibvopgDq1
noVdTKLM2+i+GpmCmMSTx8cJIRJorYIBBGupF1lOGQhS+1+ivEQ+yXMl49Tv
hQW4OYIsT5GjSKBczSs2+otnv8cPjI4LjWMD/nhidlvkTb5E1aof923mMlSH
c1paE9f/xqUQHZJfpsotwmKquyUGEdfsDbDs1F2tYUE81Fdne7mkhyFzF1A+
LXmNW9mhPpN33cXnl1wxEUW2MOkTmGWTrHt8uzdScsZ3AuFCf/Bi5hdW/JI2
+q5wE6keJLbSeFqBCXXQW8lp7nRVBqH7NNQ+Dz90FRd4DHeuxhb0hP2IzqKM
UBbCXeY1Zv0vc/UCD6rHN8TRp7anAfEew6hLLXSmjYkizl5XcGcM3rMCLFKC
G0gWo0FZ/tBoC5zeOmvFnThl9OC83zJqPNf0s56IYlWCDzXVmwc7uWbDOOUk
kqtk6i2tkj75FPVnD6RbXtBXfF3HSiDvLF+ATqyRXo1EqAIeREQr/2MzfW5B
R8jeaWDV/EtaeS3jxK7gTzFdjlfKwEXLZDJKMS20wTA3jZf07FNoTtJmrrqW
HcWtbPc2EdOx40jckFpsTRXOkscqWHb9mncpiTYUgWo7u56W9cHZ8xacWyF8
dUOmXN4HvDVmNUhCpfE+MYmNQZsaMDRL36VHe+IL7299VkRd7xf2lrk67MNY
x5DmLUk7og7dv1UY8l1OS4xomRv2ljNY2hiRsQP8C7HAAUXsx9mI/bZY8ZU6
Q6kUhfhZTDxk7eSvGs2f3U24+6QDSPdUYuEu3TELCfUQ5FGdXsoIuu0jnx6u
Df/JhwvpCaotfsMcHQwpoxnrqw/zhxlNjEDWRP1EXWcuA2sbAdO7a8HDQRxr
VGnQznEPR7hzAIVCp4dva664YrXdWc2JTrpcJBS0+YD2S0Ro3WEPSm1YNKsF
eWUjFKRWo2fqRpPAV5elp3k7GYYRHrm/9+UsyruOYkJhY7vm0XVoh3wyB0Uw
qVszL3i6Cj8Mkc9MT1ZPwrXxVHiIHrjspRbwDeDiK13IuvrKBTCrvXJIxwzR
YWNnDMHQ7hMSeUpHfsGuaqmo0UDfkGRewxhTwwdXjckh0CXwnrSF9nRSSTyH
zjC1T+6oB5TccGluHcGCFApzZyXA3JA6PFMKRh6U32QpeHobnqjeSvRaN6PN
u4LqsHPsXvmISzdUBico/H14GrJrVyomad2WokAIK+j2woRwtUCM7tatupRQ
x/B7D7ECwJznVclE6m5XS7san9vuQ80+HZaSEPCHSBUnhtnguwqQiyQJwrkN
gcNLnvEf2qH4Y8Ym3pfPGv5+vyiZuqqySDaKfVCLei4HF1EEIDigp9cUZKvs
JhqNHzNCX8LKy8dAppm9AIzSG1py5kCWheqZ38xTfdgYL6EAykWW1q72W69b
NWiEL7I0+Y4kxfRT1IRs3WBn1MFxQ9He/ibBI0L1xGD7JxCQyB+3pMFHv8pu
zdEqzgb4B5XNaXjQxa6I2/WK+PTtrqRlJZ3WecbqFBI5clEGrglj1iaaaZBq
pc8yR4L1ySiQJkA8PLljrzRyaRE+wUwQzAh7ehVrP32+yVKpm4dDz+yg0My/
KcfALhZbh4rGf3uX1qIN9GPgJj4PCuKyzJBGkA4S4CHTTBKhlUWnUzsz3p1u
8AMESdePe1Oa6vnv7vkrzKz4bSamz1Hf1Wgu41Rjbqnx7gPvW2oL1+WPJdJ7
20NEx3Bh0AxIJSA1rCxTyGO+lCgaeFofKRDLWqzt1yzOtqeDU7pYr5G5Yj67
qhmnW7wRDPA6KhI6GXXIW9wng9fHPGBQCicVUxPQ/SbMj+i3K6ouHB+foP2E
Bm1Ez7R0oqLIoSL5DKyKj+w2fHG+p2r1mWmWlsJ6dJzSiD/F5GJSIsvnEmeM
932OMg3LhQoffBxiDXoT8e99BKJVhyjJ5sGPjMHCilqk+DcaozEjAgFVpS5l
I65HWqwiIP8CFhq1az3wyAc3mgpMtvpa62Xtw0CC25t1nRnuagadeLgsMEDZ
rJtOorr5VoZ+x5dET71gxl+Obg/o6lLZA+mFZsbdht+QY45tbPFhi2qQ97Ub
Rd+IaNxi+7b9Hm1pCkRJq05roEraFtgqD79eUlsYyjZI5I/QxUbZMfrB7sXB
VZN4VKRMn8M9xMbWVwGdtIBFjpx2zAU6nLYkiZCtI0oa7HujR9uk7zcqn0N5
9Tw7zSU93fTiVIIBZ+jWxPhmDyDQu3UGHFqE1H88h2Wh35zpqpRkmbY4/Lsf
eNIZLZ9+W4lhVgZr+Qj2qPewVK+VFH1OSTJ/7hwS+N2PW5rF+ihjTd5NG39w
Q02WsXq+np9GTkvWNKZagXvgKo7gxnBmzoNodaAsQocVr86QZ3+YKaomC+23
nvAdveMF9gDb6+q8GOsrPBscsyX18LAS9lSsODnoCZLnVFGEHGB7ZRXQ5LhM
1IPTobcgC2Hc5IuR+vHeBV9VXSWLUWgfXn2ysD40Ej+tvgqPPMe0VHO81OhK
EqDRR5IJGXvwCtfq4HD6baChrksuqqoCQqfQ2E10BmxItKQuJfc8lpFhB/S8
sRUI607TOYWUpTBnU3keSvUlHEpCMVGrdf3IajdlH4Vc5BYdpCkj8LFkMlEQ
DZeAVTlhyMnvPXycJnaAynLlgvFkCd95k7BD3iPA0sSEVQfg/kwOYeyh0Z2+
dOyQPgCcDnciZeeu8TRCj5HQvITo7bYhn1B9zSwXBEH9sUClyHEyBFQ8CUBg
C1fVIKgIqs/3TRmCLpgACJHv92QBadZNvO6L5g7ZIv+SQCg75uj3n/Sx0WLg
uwq3q4xKPhx7JImbNnq9KE3OYGLMXpnHZ8dAakjCqGuf4PXsfSIQCNx+abaX
pALzjYROkt+fHlG6Qd7A/lUaAT5jydPLv0bzw4kySy9q0+I5u4yxdeHb9JoN
XWe6skrvrkmpuVu6PJYREiDUZMudn5kBjkC6uxyjKsJZIWAFIJzGHcAQSQ5X
yKGNVzFODK5Ih5qFECdHccjDaHCeeUeBAivtV6tY7SSq1WYfpu9zfdA4Mx9z
TJwQ/B9xl4w6xStFMdSkS0Jhie3AR59aEK1g4YLztZ8+yf9SfAXpnoxuR9hB
RwXSw/BtM4DFtzkXDkSGOzqmf44GA7khID270HMVPkdnUZcnLi+bJ/yrzsPo
BMTf2afk07luLvhlXexttt7dRUMeKM2EeJGSnkFAQYQvjbDIJkBXLEP35YHl
oqfDJ2f607EA4MGlySTpQB9nZ+A9+w1xD+t0LGBrRiGP1MY3QKYOIWC7JM4S
ymhDhiWPDwHMD+mYHE6ahSXFbxMLa3Z11btwtkgerfVSj2RLtVoJeq7wEywl
tHzqa6Co/q63CRef7heCYsOmeZ8vhtmITHo6CddS/hpJEZ3kBkSfXH8zIItY
MBWmodiCMaqoIsABb+EpmYugrplpmlI8OUQjh1vHYQ327kATom4y5Rp1R+1X
xrGWlr4j/ZAw5835Myg6JsGgEGp/FqTqt3BSFVHbYl4Sw2iZ51AH5Y6KPsg3
ncW503h5iklj/E/VyBjY/TYu6bXSUXNXpU6q8ZJpB98APNKkt8BhG/wwHhcJ
49YTJNyR4a8gOoziz1Zz6HuOqZtoGzPuf2kaageq2p1DgcPcQIFcQ6wJkEPt
yn3HFp6wdlM3sHSx8J6J/fIkrJZEjXW5TC9ygYaibZ3OlPXVfhcQLdXNmCga
poGjet7sc6ZBfAmgYuzHG7SoCumIbczQlhNn0FVGfFw95GIwkZUk9NmgQ327
mJ15v1lprEGkm22RYgIWnD6cIPLazmPdz/6BmuKwuylJbXW8aYx8V7USearf
0IBw0N0CBMmNcjmdDBDHckQ/K8vn7ZBjIw372lPLlvabEPZLp3hUoPvRtaaa
B9kMlJpMgq62bjc+FVoZ6IRVn6gmAOtL1F13DuqrQnIQWmUvhDuMvnJsdwmL
9RAMLq6fG2CoB8DWn4jvL80f+GZ3ufWVKOVuanpc5HlsauMTr+6on4OOWZVn
tD6lYjnft2163sMTWcpv64TIxff7sBvNcXKxz2jaWf6J3G1L4Zdqv7BMX5cf
qqzxpjEkQIlKZLSpV6hEEC9Ylm/jCQMj8ICPGAAKzapjP0kcR577ppGQZ7ln
j+I63PnPPny2JnIztd6VWeZIZdYeQhOXeu/WecKS4AopFqVLw5KNUNH7b0iH
hhSEdbZbeBVw32xOI2N+ysGdygXw9trNqQ0jN0Loghx3iF3VZTquxGVzkcmI
DLcBr95MIHeYabPu3rGBesh/1ih3fe6pYSjHW2DRrkRIcem3pVjgLLMjrRac
oHuBk3mCp8n6pCSYEoj6f7SspH8h7JYsnC5tFj+RPnvlTiVA5yJral7Jq1e8
G54JPxviplk8q/jrgrI1Vue6Id00TJL5Zz9MBSZjvSg70niIHv5IJnmr02bL
Tco9B5LIEtXy1z4QN+zJGwmPMYA8CpaFmJeHLij1b+l+OS5RdeyqbYnbU5X2
UjjOm40f46FsVgejnegIXdTHozX8IFxrHN+20423rTjOwpd/Tq5ZQRl/AXfY
C8jeMaSjUmUNlZO8f9qBI3Ii7/xlSe4LKhPqRSbAPE8G29INgH5JEjWKP8K7
dOp4ajbNmtUURivaQnXjLbPWHd8Z3Bxn6MjuWgFSLA9CEi7ggsvSN09IRWJx
y4Gob+CuM7RWQRpDqZ3+VXe/Er//3V5bFNowPO24Bt4W/X1FxLThhSb5+pAt
fH9W033xjrrpOX+hgEXqjc3ehHflrNLgfTw2HyoiHMAA0Bj/prGrojFn/YRR
+SwzWRxp2yv0Z0XmLxdYJRm3HY0JflB4439OtTF6L1jjXJvM0umnwOE3/5kb
jiNemVteNw5Y4zKdS3RkunxdsdgYthT85nAkZyGRP2Bp3AvrOzv9KsMHaIMV
sjGGMkpPh21Uh3mKmfOy0WMSvStDpxvWQ6++NLofUoSo8SyLpwxbM00VZp3k
Zsg37mLPfrEEL+bR7TzE3TlJrkHLohQsv1zSml6Mj1eUpsbpCvYbG2DJT3G8
+Owts985fuMEzPvmDNp0calNHRU7+V0mvu5/q003qkTo/2c0ECojhNowBwXF
yAG9PlKjS0YNNX6sc9Y2QpliUeQoO81nXL8b14mY5c8cB1lenDywtg75WCwo
LqIJpSKVhgYhY/fTURk9OiOohUOHtT0e9JhK0jCIFaare9yb9SdkRw7Yz3dh
c/pQZrH7pqM7B8woDTa4vlmgIvLLb6ejMM7aV/+iRVVSbKy02+7BxBebnF7w
pMde+A07tVHWZ183bNGHE/XrCNMy4GkxOHgN2Gy+rZs0hRAG+3V4pYireLqG
dfLz2RXCB0e0G/FFH5ZzE77+8slxDsXDaiuBNHRqwBb0BKyNZSQhEmjN9TGr
WLHcrTe8CaQ0KSIW3wUwO1es3b+tQJeRVkReuKC7P1B36bvNuBIdcFEWCm3k
PK5pQ7bq66VzMCkXi+CgzCplYtQI0EIqIk0zwrWrU8hTpigarrwyljwiSkeu
6+Ori42+DVlnUXj5rfzmSGQGna8055rBffHUPpWvKLgp7XAGx//ReeNSX34P
mPhkQ0LcTzG8Emo6fRSNTOydOyT3mFfUZzhRlNkCZbNXAFcvKTs0+06cSuSn
EtxTgjj5gvhzvr91tG+mUQMwBi2GD0/f5FN1ELJgXEzCKxK7nT4wPegRMl2Y
ZvKyC9Ynd0FBrqxAQ+QRH/yR1UZlFU2roKHG0KLU8RJ0k2bSMwpPF10fCqUn
DovfLeSET4AGsw6G/jipYvN/ARKPzPfwsaa84WfV6VLwFLvzclP/cCdepaES
6lBUtOJvIPsHyN37oCk9N5NXOxntKsL0I3Np8EFhrQS/ONlvadaWmQ1zPAhF
qzHf2OgmbEJLFCwpklOuQ9JePuRXIulsEfS5dci5Kh7tRugN/kqIeXX6YsuI
NiXOduHQ2AVn+E//nu/J9KyeNKLD20RuFSvqt8ava2hrPuk2lVv2gtA0uHcO
1+5Oe6dRjC0aJpFvIid0ZO/Jy5zplYy5ek9H2yT9sRR1/a8Tvo6z+ycZJp4i
XKrongdQqEKe3gkMcbXKxRhYDQbIZqKaafPqvoaGaP1Anx9aN6ms+ng/B8VO
jbnl1MnO54k1jUrsAJ6axOsqQjjFe1TlwfxOw2xzCcH3pnUDSZtIurACzZtR
kj8HAEQvBthA6uzMkHhiDB7o4npNO/vgKR9CgAZqakOl2cx/jpEf/7QfkEFh
qS0KDOhaexkA/xCuNpothtsyZI6GnztpLq7TsEgl9ALTchjX3fiDEo5+PP3+
UDO7uFIToPEg4sj6rvVAESDtyggvdcX7NzfBRhl3ckZYhxHZvg8IlTgHhPoo
sxnaZmhrwRRO7JZcf2xYTU4Q4t5X+b3uMHMZLA/+tx3UjzbuhW1GKIujDRJG
rPQxTULW4fsLMUpfrDbTGrp5x2r5x6kYw8ZgcPcD2eLu8+EdnGObsUZ1RMg3
nuH7sjStPxdsJpK/93xflGy35SGEk+QSlKlRyjL74bmQb9/aoebBWm00X7nk
TfRHXhbMW3DLD8hWnzTGlm90O47ls0/y11uZ16pOuYwNCuRb6nI2NdojpRz8
UVRoY1CgSn2CMMEZg94glwOf9KmuztVw5gfOAwSS156bePeeMzyvaipCRnXO
NuRG83pzNR6bpR5fcuRAx/dy8slqw6KUtKvidjQ8QQqSoEQss+XH8xLUrlZX
sfVPDLAHqFhOCXxAKtiMIMlR13ptDv2z8mhpO8FGRQoTGo0H7PWO0pqkFBih
oy/D892McvL65ChVZEc9os/WoYrZrlmUufWA6RBV3+AsQpCmcHEdozZWqA0E
dHLiRAtslRgv+7WkGKf/k8SSntQ1TQVdbAqMpAcezQr/dc50QqiBAyHzYacg
46a8MKFSsSBVqmJcR+OlZxk3QYQ2knomzIWoJi/NQzO8kWgVcEqBiz70SFef
meVf3ABxg+fEEpHuf1+eFQDnyd/bsSQrHyDLW0p8dlrqoyCl0p++oQKV7PkA
s1S8HZ3wcyE26Mzf23XMbgWz01KubXjzd+axbQUlFPCu+8ddiuKByU6CItGj
JKvuockoRxOd+az/eoSA0NaLY2Ow7klwU04gY/7mcaRAtBVe1IuQ4aCD8132
gouM2ksrDIoSZ5Sw1+TdIaZDPAlkT9iPp9c2UK+l0uQ3nMvQIqbvZ8paYZIO
6iUT5RE3MZDsKSiM5HwQ1GzU7yd66JdKfK4b0VDTrsbQQbSmn+7BbRkSz5s0
lK4qjrczxiK854z3DHI/dGeQE2w3VXt41LElgqMSNnuhGQ1x/LMC2jWjl8bv
Z0HSAEd3BmfOaBx4id4VXHeey7HNpv/gyeDiFwOu7EDYMTMgJ8hT6C7l3LKY
QSfQ332emQCgbtb+HxJv5H17AIj/+fMrmW3OfdETapYAfw9iMTshH4BfYURA
x/n6aFaq+NDu/P78fAnvB6cxNd9H027iIgEM9r3Et24yZPeYn/nNoHtMWxvb
jAXD/4rN/RbuOg189jpIlMYDjf/btH4XpOgKPHQgQHCCh7nhGJBnYXyWahU1
oUTYrT+CSswBeUZzEGUlEslk8uuF4dTI3DsLLADlCOa88bb5e/Jg8fSaXFZk
w4aUGk/sRFKfapmpp6wiJJuZOXZgU0dp4SAewAmQ8KpZtL0QyXjqFDXQR6Jo
zOyMXKzPL6inLMPTixfv4C+nVgXg1ELwjlpzwI2aNokmJnx5ynEyl0i3W+hN
Syi6pkOFmPcVxTod9Et3IOK11Kp3u/ZDY04Vey7hwfNSppMDCxQAwfNUOvy+
/ImbVchfznSqK39jiF6gRNtfJT730LcF9pxqmfza/lS3pSKeH3joE6lXA0EL
fKh/xi6uLajNzcvA0Ou7O9SdysS5WYXAmD5OJU3QUs/SSccMaeXuXi4QQD5u
I4kFSSMD69rKI8iWZXx8H2+RAVSgiqU+5lVKX0Bk5njtww3BJWCwzwaAs3C1
fLecd2WSzQ3K6Moa18qJ3cKZdmuhlFc3cx9aV6uqVPN25cR+xTl+5HlC5+uK
j52Dt5Jd9Kh3xwi/U1kTjc2Hryq8bBW4fkvLTrNtDp0vhTGUHRzMCwfIvW/8
6v9lzSpcaoV134EGlmwBnb+AZD9jffGDxK/0CrNvYJjvMbWKsD2LNHutCP/c
+NggzjUfn3Oi9P+MGAnRHEo9MPhMEVnLBtx4L868yiyPAHHYXZB+tudUPw9Q
5ol/fYeGr1jJphht2daVW4wzUVQ9SWS6fIYVPSYoN74wyuMgJmsjFDaGKPmF
yvUjudUfu+Ae/rh7V/RmkFXorGyUvyjJB+KVc9roixmojiILIQXntpXnh57a
0J9pQ1MBrM0nRGnhFyWmgZWWI/Q7HIVDbYNA9wErNbh6e8+7/V9gRdQRqM4R
bDf1S8uCgLrxbtztaN6yE0v87UEVDbHWbDqpy5SoXXhctqwhV+UrjwXy4R/y
IOpATByXrIRmeQRgmDB16UjBJ+1Tr7WMqEDO6d7Nz+bZuufJdAgycL5yJ7l1
bLDtVynyq1xk/GiFwh0HmJn+TDRsm352MlDKNZb1/ju+5PkIWqO3pd3OFCkB
I4UKZYhJOr5etMFBi/3oGg1QCOFxK90QopgMgSApsvEOOvrI5YPGL5Bwuhft
0BRBnJ+4nP6MdqKiqZWb5Sej1uweT5ddQcRsO2pS15IhbcxbaX7tK/sDERD+
Khh4HElsjA6hgY8C2h7lqVZQaL0AZloOJOKCZLaEqJzWkIX3d/xdgqcTeHFL
xhrIV1QoJGMi0SkK80Jz1jy3hH2scevyJUkHcOcwFkX53uFsbyZ/xUlEP9uO
h7HnuhPgRdz1xUILEERiJHnjYEk5FpB3BtZqnR1qb3iwZ+3MLDMSBaY+Ja++
AJ4AeU+KTYkGsplffenqPcRkzKGSPuMa0pM0y1KxgouWJ250ENA+xclYw8W3
zhMQziToYPuFyx0kKgDE4fC8RA3qngWwA02wfONcgxDQh2KUbg6okK2axMFM
WCsXtTxWh4pNACD7unx6ENa85INY1tOzY9/gbQ6NEy79rSBkUv/UTBcjsLs6
vfWABZXaGaD4/SguCNDlgBfCIkEUIo5ILwZdLCp3FLoa+uc3zz8b0F7dP9kt
dUIZXB3/lSym+dqtsV05Bi8C7KXxtc5ik83wdKWahoLSl+SNWs2RV3BMqdlZ
J4GzxonYa73K1auy9gtbngIV8DDRuEYsyP+k0+fJ3f1iYrPY8CWdVU3k8Vef
ESTbVmV6AheUqPbl4fPV1VpOj5w4bhr4NPbbfjDncwnYuoVRSFm3TosIm3xh
2torY9Chv1SsAq9S/eUsvSQ/B1Sx0zlH0+EOjBIVCPfO4GQWWIbdFtS+wc4g
o4PU0U0a9bO09+sqApxe5kiCTR9BvVrV43LXifUeUZGmpu4idY+Eq8QT+8al
1S2iqvQmoiAUyPuw7xbBVx6O45R6hIuUzZFZUzZ8/nfiSOr87guYl0Xyx37w
1taSNrgxm6iKnyKJL6I7xrrpRzX1GTq8sN+X7Vk+s7v5zxiY4YtiqWeh3V3y
qE+2vDW12fPdYAZjLMzqheiBew3uV456d1kB7s1XIJ/JMlEBurvHn/bMBy8e
piBV7/I+bUJu1Ug/vEadCmfBZgD830KAWRxiXu14ibgI01VXY8oW9zdQps7o
Lx1ldFvXBYwg4brbnErqgorE6fFaumt2rxHjIL0sSr188NXNomQd2mE6dgn6
UW7UMKfQ8m2W+TreO4fWqUduia/j9kAFgeI5aMPF5QgOSRGn2/OKG8RIAA8b
Th/1wG4QZZigJcTkuBRIZHskyNbS44S47sEKHhhRcCcCA1nLPcm8hg5y5EWv
sDNYraH4Uj5R465b6MSMZk5bnvXA3D7Mwwgxesn+AdLUasHUxjkZYmvXywtB
vLyiLDC8hn6c/TpS3v9y8FH/Ousk0JNceRC6cnfKlAu975tNndd2tMDg/Vxa
X8L5npzjFB+vQNuifsXl6O/SJTtag+35/RghmBUExSbd7Gy9/EqeOXCU9cU3
Hi9EHNUyJG48rITKA6TVK2G0q4rd5LoxwiKCpvXWRDwtZM47IL5/54548PkR
1/KrrwJOipqdbHLX0H22SV3yH6U/tuO8RiZmUZ0EJIkGe36OEKnQVn/QXBsD
dHFaxUqsFbaxYhzQG6SDlxEPA/xCoFzKzD3IJMGXcdPiijBP7gXBU5d8+cCJ
WL6AdOfDxBR+KTK5ZFrpfqp1JQdjxXtgQXp+TbfEJiJRpX0OAgXhVwgJh+Fo
zTH0KmCXfr7yM1PdF/Y/OGOYv7lHuiX8dIVS6LUh1iGy0ad2ikqzAvXLZoPm
/qjFUGx9jKnLD1kruO4U1dxovncxo5Y3LM4s0xBO+PG+C3q8G7wvjs8P/MeD
52Nf4nwv6EVtZg3oOff9aPuDkg/WmADD5cjXR4WjLTNChhCSfVuA7/K1oU0F
c4XfgAeulkFm/xMKESq/GbI1ySZfcgeGh8U2v/O3nNsviIUwumvk15ifXud5
/cMCTOuFWZaj6wnSuIDc4lbuiojro/XCG8BN9Pa2Oh22dBItCu2uDNs53lSS
WGNOy/Aztw2Fwt/x6yxDwYyA7nXhGsVNb3hgwxRJjy0HcAbgKotsrBqBia4Q
NztM55WjnlGiJi8EZPP2QI6iZWMlhpbffk/6qb5OClZGpXBo+SqV6o6AZa6y
5NBMZF9GAsCTDOo6XCKgEON1qNTJLQDyGZBf06At8Bb+/bKswhWz88RTpk+u
O8Kxs08r2IFcsevr2MlobC6Rmk/yx70P+eB4j372MCCzMPYfmBgZ/c1t2PM+
6Q6E27EdI5WVyyvxUMF72O/VKb8DqjmXQ5UrTpmDEwZApBosiA86+E7oZKuj
o+GRAsJ4N2GqSk6PTEEe58dJLovmWEpfhyGeqhCtjrjKx/olgudyZPCt6d+7
HHrkLiPSJdXekshds5cBf3FT4j+IaSGKW3+pN2uNvfawqfBU/sXxGihvFyT1
d9bmFfEeI4i8t/6yB+2w3XARoRzgaDnQKBtd3qQQc/1rTeUKG856Eans31ay
v1o8OQazLy6ZXiiIQAI3y21yGqsJsi038DsPw03fkOnR0uvvWG+B4fuTU+eD
n+xSlgUHx62YMQqlD9YymbUB5tPn06816pQp/wjSFtrjh05Weg6/8BXi05gc
wFDNpl0/p0tcJvv7PXpeOY63p0P5s8RAZZYvPvp+w1r9m9Ia16BCyGuQlVGF
JBdGM/hDQXwr0kAlIaALLEq8dGrVXhDLKt6R1cTJNBre7c0L01o5PDYq8t09
7GdY/T2Bkwiy/m15oAvBHsNanOr2GqK/+z9Kw64LaHMpfauYAGPIODplqtsc
Avcw31sziay7Jrlow1f+TSYF0ySczDVdE4n9Hajftsi8IT6punJeyd2j6pDM
Y6TfmySDtyjXqweyQD85p1XV1jFGVaIsOGwQuv43GbluIPLu/6fQ8/Hp/Z1X
uxNRHx3j9LlIvdJocy0NDs6AI6IhI8QKuyo/3harO1FSGTFrZZnEn9e+kMhR
a1w/g1AYQTqRnI3f1pb5wbfaCKLJQD57WyvmE4Cai9P9fq87VKRa1y7VSq6N
mFlGeJeDc8L8GWKC7Bes62QBbT5YtRni3bmjrZ0AgBjkcZ/aI85M358erJGz
Ovq2FLKMeVDmexlV8NvH7kKAI+xUGx+CVCiCKvn+14YSSiR54qvtBnFaFvZ2
3ZPT0nR1xXR/wKTjyVcAWU5sr1bi5rhFl8aQnfZvVAIz6bUw5HGojKJMGb+n
UsB2xcRaERaMxpAn+V1f+XTUomdA6Y55eA0r7L7S5T1vRrbDKY8DzjQ3XSWA
cjwcmI5Emx78rE56cuBIDto14IOi3JkJG+tFJ1b+hqDlkiCYO733Z5l1EWnT
c3Tec/jCMPd7gw+E+oCBXVUu2Tc+V4qFNuktehZsQ0cub0d5Mf4edKuaiANY
mQ6xTVj0yUzq4+q6XC+UmYTsdKOO8qhC5n9LbTvmUP1QsjLlpup7r8zTxO8E
JbA2VyV2b3yBSeZIHYr50/ZQPtYZsSSSfpuUAWrUi2yCT7e3dFKEn1pXwlxL
ZZsqcJZIjevNvMF6NwkLMqEt9EJ7c5ITFm7iC/iXy/tSwfBkn7D0GsKj0I8t
jFgEA6cwENA5TVQThGACDOytxvMDBmPg19K52WdRPuIcfPCJaUYtyDihePTn
Mntv6sTAjL//HyRWEL3dDJrlkJ9LBz2acxZeqDAzY6wvS3b99zn+JnMGfFaz
BOVfDTcmZY3WcJ2bmRVxoSio7CCrO8S7uG/1ie5PCH4Ee/vEkEuWlBwCgVzt
IOZbYKG21nDg/uyonk8kiN11toe/0AcL3pjm7zSWlk6/OkPOS8o+FIgOqUID
O455BW6tjFm2iA2XhN8jfGkr8IrxrKGG57ou61WD/SYq8obVMGX11zBFUtWL
Hpl+4HE4Uz4fMQTj2drvSk+C+voiTwvWnHDk7RBVKa2/+g9WrkKeuaMrME/s
lfQ+u2hWnHx+zkwbS8uGhuk6ZayAlUZUoVywQw+D86jw0kv+JSh4QBukw9IF
06hD3YWP9Jnj556RjKbbWqbstAXMzR3GKFcKZ82wu8UXByWWUitUvZh66oQc
4WjHtBswLY594IEuf135NsMl5LxEWq5/kUAS7JJOxxdD4Q651jtL/IafKLFa
JS5zucIcdpZ3DJyKWvIRm9co/lHRfAI8S2Nh1HchgBMCRMMFGHCbR8pAZ97n
cW4QaUN6dlqSFtB7cq6p5EQU1/CsmS0Ya5m2fH58YFRYh0OBtXCQLQzssl4H
VBXL2OFR5YUk10gu5gImKmTcFrurbJudw2D0HigTTThUzcpa+KsDnuxTQbHw
ROJQTGwkSsDQAEYlL9V4pdfJ70o3MSecfC+usTJ4NRMUgYPDjax/0vjKdFO7
qTaWLWyFJR272fhFSE73AAYCZOG8FKLk4DRpjTlMmAxd960rNOHcvMqkFvW3
U8PTay/MQLEPjnNMC6wNUcZIf3bmO+WhGg38DE2RnZnlPgzaxRXHupnQIPQT
Whc5n2l4Kh3TmmozG4dHnQJLOYWBFdYrZweRuS8/X2/Mnv8dArMfUijIxiok
ZLLslSVrdxzj1BsOQxeF+reijDxKWA7o7pO05XL9PlLz6vqwXBGRHtb++ss1
z3zeuruXPxlua3o0BpPAQbtdHnsWAJZbGAiNs4RULgw+JJkC5IqJHW2r2hKY
9jwl7IQ57LgFfsPKkGYMNgWXFG3XwSkv+eOuTBa9m2PZRlzBLK/N5I4EtN5g
ExTRMYj4OpWc9gQ8COJQ2ivkWYFhL7rfE3RURazAuqXrx7ivlGIKeZomKbEG
sx727L02pKAR+R+ga1bxt85mi1BAzNqJ7CHleWL6GitsaYyR6CSFAs+7HRLL
0bYaytMniebD+c7x0CkfeFqJu6uiER3KmNCxjWyyWF8ELSMa1Knl8scS3Hk1
YLm5qYPpjkGaICDuaqF46S0WMl6a0JCxHG8FaDWWDCOke181cjFN+AlGjwAm
O3oUL6oCF+OAMq91mRbaPELitPQayt7seXeLyxE0K5u/PxOWJAqDz1yKbRgg
9M50xfOLwO/5RtLIWRZLYLMTK8KVMcPBqnkEQ1BFTpyRfYeYIRKYv3NQ86uq
vCKUHtGG9HzercN4Bs9MM/WyM0fAdWowqZthnDXN75Q3ROLFlr5IMJZQXPc5
Bht3FaZuIW8Cii0iXCeNVNoRV5iCukz4l6yPI07GymRml+J1lVa5nypzjDCs
Btr38bpsLYNHNs6xzvdcIm1j6WjYpG+/PB8vWQY2BqPTiyaTCLIk/TK3tXF0
K7MZvhu3Jc+EAhBzsJp9qUvTe/JbDU8Y4Q/XrUorYAmXZqeBrVU8ih0DYxQv
N2+KSzZcbckYXlRCjks4oR4GF1QAO1mgp4BcM7NdVo+m3MWTQkv7iOfhKCJ4
pkzNO9Iqsd4zbzWRzuX3UTt2vDxZiIPHEuxVrwNCx92ndBjP2CKMv21A/M/Z
KqBytF7+BDm9XyCaDcc+6M27OLUTuayzXQPv+uC4hVv2UDPaA9bniwLyXqzy
Hkn+Dvu3A77UsliM7Sc7StKrRJe9KGkjpKa182F25SPQQaFDE+q81u0u03kS
GqKjXCZP7WQmjny+GC7/znVZLIe+Y3sUdzjbQnzF5c7G9o1gfWGkd1p6zrrw
XNp19AbolflMDXMK6c5uZtCYJfNw03rBSHA7fMpGLgq/fxuH7w68DGfdrISg
pvLX7BMxAWwR/OfQBr3raR0FbkqfeQ99lw0Zut/LcCRWBMKVJeRCeuxfxWoS
gPxm3+hE2aBk/qXBLfTY/sADFa5Gmbghb15jS31pF2yqoMccje8ND7M+Et9V
cQv5xqbeGxCEBQT2+/A/BBN627nmteeDPIG2mWuYRFJTZ/WIp/R0O7YGVfFt
d6XMdLKxlE6r97BqDqgdI0ZO1CTX1pRwEPyh2WkyMpeMsz8bI9ztQlpTTztl
08RJDqHk+mVE0TdhNVA7AW4KgeSbIzF5KMkWNie0U21PkVNWFff9idD9EXPR
a6lUpxMp4ht/5ou2UyCLNEd3cGXeHEj/BK+6kXvYbCtPCv0sqxVOQZwrp9XQ
7CikSWguJIJZxXQqVwfA+j/IaIX8716w2l/o60qvQXTaQGslk7XGj9HtS4jb
G9ty3Jekdb9cly2HcNCC8YEccYJCqXsPXXNtzvxsGP8OM150gEnlSPlRUJrl
Q86RD85mNm9P+ZAH2o33PA2JbnYrKbMRA2QR0ty+PfIqZ/EiwrF2IZqLAJNl
wZKZPYa6ijXbbnmM7dBAOIZ01/RgSVDBF00rDsgJjIBPxPaEhHqNXfIz8JwU
BI9enfgmu0e5+lLdeXaipewGSPOH5smhdrA2H/WiOwP6/iixpQTxSmZC/qsl
hw5FjVeUHe4LmiJbQ+3ELn/ZEcQLcoyYubMATGkrr/0dJghJaHZH1GgOzbrc
bZDMvFp+GDh5F3PrEGFNs1nPXxeJFWqCibJGB25/p4b65z2+fkfr9RoIlXOw
V/M+otn/ID89I3qElETtNj4sYa5zenT6mpr1iFivsmXgbRbgCjDubnTfmN3D
1iZYvUnfgP1CxbTtXzvD4JO4AMmBVZF4WxjNk+CJRPobC0lGg+TjsRvGrY6r
SRQYIQ0gahmv8GgLI2ehRLiIaOJnZKC4UIgN04A05weH738HjbHXk/h9Z2rx
4caVkIsYN5OfZRelvibQMXYs2mC5nKK2TGsI9kb6UchKVGZGgD34SqsXKmtN
cmRfjno7Sujdd9mPmW3k/5D5kKQGHNxRM5HRIjpd86ZLffW54yTXPxNNWQ6y
Vu85QaVHGZ2B/Vm0ur9PRQvUah2445tv2sYsBkG3n1WWV+NfjyqM6vleE1Yx
r71UHmv8d3AM4y59CHuPb7Gaz4csPyn1XPUVH0J6Ws+TxMyN/COIOtNZYn9o
ww0Xi9IREgko2jo/nR5vk6MAkkRhEAvGwBU3yK2JteuAY/XnH3TDOPBj1wA7
O6ui/+MmhiL8Kfr6NvQIougsNnoNRdiyM7V1eMNi8CZMPsuhWtY14WaictM4
S2V5JjBYjw2EiXsYQTYHdVJOgFWpH4tLtZPA7XAS7KsE3Q0cGDgYopiQ3LZ9
RHGnC5Y0rHvULpUu093NN1KsTDWLutDNNaTsnmF5jz5tYCrI7TeYNMZbJ26i
RNDGhV3CoVYbGL7Pe+QLAH4blN7DavkFzd9qkozj21sYh4r6XGfGHcn3bZz+
15Yxa5bomzp6FH3LYc+GGoVlCAFWWnuz/DLGPMAAIcAR9X4MsF5HGL8q6f1x
1qLagyrOCXCT3IePBCCfdqvTzywXaN7M/GPW4xontU0vgHO4NDv9Gb25/xpL
E3MHU3bmtRmwjRcqLTWPuYsH753urf7Xm2X5DzXx/Zip9+nvVf1gAUbcRqj+
qih513ljG6J6jyYbzAd/7uM0dEYe6wwvRVwY3GkmmbErLF+NgMhs2lVW+0xo
lpGzy3ux1qSNjEwOH9iTs48SH2s8KPEJvtJNbWEp6BFGTHiyTp3C7Z9Tu1Nq
kWc58CYGa7DtAFO3qc//stuQ47ze4eO2IKdTcELcB7pDgAy4a7YMFyGb3/vB
gdE1Mr8SOvDaokPM+Oc7GnFtmG9mBS5iJNxba8JRCjEjbNwQ3wL+ACxHdxbr
sHF36lZvTygouPdndNj10RCSFbCEBiQ9fSGefshXrNjEsDtsdR4fOj2Y0ohi
lKcrCyKc79JARPnbPdwT71TttTVPO7FtFTrRbtUu2Qdhd2I0a5brZU2jquEO
+ZxnLB2diu7PmJpWIwL1zwPoZ0OGRrGdpVYsSJuRUp2ktvyff1tPWRpM60sl
J+Ik6yH1ec2i3fDifXass8dX8Flvrxj1jMwbo6XSf6sXFqpd/kxKuLNXX9tE
jnogFxLM5d4I5eYq/aERlk7CwNo1vqTJ3ERZkQCidb3E9SibuK4sYK5pNiwS
jNsc3XComy08yRhGtXK7srDmyXpS4QsN52pF6f5LBGRDDF34qUP7gnondfaX
nRX0nEAMYmH9wbRezcaKe5K7SEAjxMDZXcrWTjSB+i/nKiuoGOEcg8SesD7z
S0bfU5mm0nuwge+/C/tkCgllsc+8JTFzM3CF+LC7l5EBVS4bsPCbopnW2MAx
dynK+RZ2vzm0IyVcooAeOBU5i13NobmErqOg8y4UiN+uEsAMzCL1rspJ3J8W
Cm/nqZNE6ClScIMNQ2FxJ1BKfrDeHE9mXAZC9Oe2qRXO4leuUaUWKwYGroV6
AjEBmLtxJLeIBy3YwEH47aZX0E8rRPYmInJ7xG4lvYiuNEA0vAQ5P4yXMvl6
5aoVbd9a5fjrXj241NF2sBpOuenXfOhlo/SjEfxX2Ncf46c9t+yWKIXDRxuA
EWBS6/L+X/m3d9qb8u7GMCLG+IZhBsCxk+xIrDFoYQqKVTMtZ4vXhWDbHDef
Fdw+zDarXSb037bopi/bem206bL6mFh1FOhz+dte9VOHlZs6KMk3ew+2xI7J
JKeJ0IpKsRfLPV4iMZmY+K5lN/J3DCTuUsbMREGVSU0O7k/V3BgDmbLwm4D0
IsSKghqlvZckr6RS8edKQIOfv+IHf56OPyEzaB2gp0OowDxCTPO8q9RTXr2f
ZbIBNfChG0GDR7ckfQc34PVVTEWlFvkgGhnVLcrUYUp5zZXc9ENYe4WaTAQm
Uu+WFqr7gSb6qQ2NNe6X62h+6pPrq7+O8A0Ccw8gUro9ZO3JN7wi5jjdVcR/
GAMjS8AzIxksgoelAKVX9WcW3DjPXZuAu+joNSUkXNBtjBug4FY6KofquJrX
ku2DOAshUqutXpvKSa5YUmCDR/WsHjt+yozbfzg4xw9CK3TOUemreRBcMlmV
ZqXQq0HkrABz1jT6Rsu3JO5pNIFqCjH2Oc9qyK2TV4xuB5Ht0f+k/9f3kdWp
DUiqJqgPWGiGVzhyCKnEg1vAW4YfD8qDZFdkrfy507g3YJTdTEqMvAo7PuGA
8AisK8g0983LpKjAVBrQB71DfghXfCYucfvEPFDwQmwU45Tc3GAU5dHo4UVv
2Ou/MhRMbfrrGS2w7cFRCMGW8gfhw3+XuCSPJ3H9r0CdihM+kEWaOdKX7yvt
ouS4bJCOg4T0RMMnOTdM3vO3h0A8uF6zYM76dG6iaZfxwDuANCWhC1zrADM8
5gJ7IERhHP9/r0LRSWtE3aYOoQsp45sPyQBXs/vWPQmUk3d25jnnZb5EJGRe
1RJl+alewVdJSH6bYpkxfyQbay5bc35xfP2uWfLNVzkmPHU2LMasNdkZNuQS
pOilGAInAyvN7W3Qty93AYp5ybxlOwS2cn0gfkI0WsPVenLsC4QEunvVkwGP
/frp82/RT1EPagDen5ybluGmwwYuvoYzPhKB9QwNkoqJQxwkhfDg03bYSjn+
0r3c6ckqnsWzwsGffRFJd9h5Fo7eUj8blaz0z9C3FGhyE103DxA9QZeX1p5F
60aIbrdStdBUJxedaWcJqOsy4beh0WbyvrTIZseDobidWGi1hWY+PPL4cWXz
ApfHWLkdsMkYSBtCA1GNEcWeC2IN/1IhsvdyaWGAGJUoiqw5LoLd7Xovg8jl
K8x9GtFcHVjG5/bAV61Y+fxfeoVJRcEBjdD7Z7H4yzaVnXk+y+1CB/8e5gA+
mWnGrCiiL+aTUK3H+wDNMM/xBYhsrSefFTzbqDD4BltkkBAW9b2XQ2PmchIv
pSomahmu5P2Pc3i+xib6rb6lxOFdQKyTTPH58QySL2gtNJ9A57S9RYZ6PnpU
bwCY/rAEf/nucWTuvI/TX5EsWXOKeKC2dz9pxxSLWsBCHEuULZkiXsijimO4
swqvIV8vn4GVGbUbZxKNFA/ss21fDUHlruCSRBPdT4ac1PTnC1crVzvvasfs
VhSlEYCDzU0LiRzsBgnKavF1SA98COI4zWo8vZuLBOTmF/gd+aJVBJE2GgSk
A1zZy7wdFyMMBiyKKbuomIB+9mVfg64qOrMdRk2yEJKNGxT8uM2q7v+tR/hn
6hJu8LuHYPcr7lntMwcNZ4bgHEyb8GItNS3MvN6waQPppBaBzrnFWfL33+5w
AUXQaL5YESyMfQRmuST+B7FRG4awdojAGPi32j44pj/72FkA9HX1QPXdhhPs
4i960OPeJyjg8lTQcFXlolGDxfjwQvm5/YkzS8zIPCaL/vzU6J7uxhVYZk3f
JDsndVLj5lW2u9xAdjKoRILmj5QQIp5MuHJgY0rp/4TK+FxQBBaFIadojO4T
TUyGtwJnBQsdnauq4IiTRMH0mLHXkqJ5XSQCFQaawIHVc6Bb97LLjtUqfJNW
37fsbVl1FwvOeQT8Wv7AfK0D1G9pvxxLyEnUCanZWncmnPfTLCjbIH7LBDVr
ru8BdGFydNVAb+C2mCqqqDopgwkaEUhJ2bWvC1t05vVOzzmoqN8LXZqgwioA
RShUWf/6SKznS41+3eu2Q+b5K4YGUHPktZkon0YKeI2xxJvlUFSNuMGvH2xs
1HNqdJtbYkqkK4S08M3OTi1dTqozZjZRG/3tnVUc3V3SPFPBVJhuelh2X/Q/
iDEq2/66h1aScMB83HA/Mb5rwJQ73vY+tkV7S0AIA/MQUWqrvi5Au1eyUdsv
aDPgIYqoLSKWKY8uU0LqgROKtRXdu/FNS0MkvjPuRUn3bTuA4P65jP5OLbwc
5/RKmF71iIRy5DApo3BWp3YxZQjxsRrngBv5eXe6Pj4g3aQTIxvS+gYzYAlp
WYEqtToNzVEA/ZK4IR95Aab3JL685mTQmO7BvSVjRBEvgMPLTSGHpo81FvlK
YsobGSy6b9H0pIA7YMuX9X2Bne7zJdYRfWf0GV4IpikFem6EJ+PL8JfGnhx0
egqXs+PEB3PUpjjOjPJi6E7Wm346UHUK45dWwWrgV8md4KsGdM3Yebd9szbt
aA6vzIT0fSZwkvpdHoYRiW0Btmjxdw91XuMQRw4shzwPfJyniWIZkgSpkLuM
X0PfpV3kLYj1+ivaYv3qSwhX3La+/s7z++vWwfV6qBa7AJfaWlRqDZ++7FIp
/v9eA7+bdRzFpT4U+Mt9BkcZgqRA1PH9vJYjUNRi32Hia6r3+HtpyVX+jIVP
B+dtEVMdPXNJUAcD0XK9aM7v0pXhhJnHVBXx5S2wN4q5ScRFOmHyOAUwKJDW
34GzJk3XVItBMPrvOryU+MOX8AulKyRMCwJCvxDBpuC7FGyLEH/RC4ByTEnb
TZIhNXMqTcR6RVc3w2r1ORBMKVkokYFJqAlyEghgG/o3J0mU6HeFw2xZlke/
2cOK3ZadbUXhIYV+i3UxiOpf5cXDRD+Ow7sVBwBzUv4ew6mJigyAM+b1TNqo
XqD0fSg2cQ7wkq2NLCdQ0mnpIv0+1PHDaPr9mmTKfHvKnTbMWpL/I37MsF+l
cY7nVMjS3FA/nQLRrrN6/ooWcq8jXPTZrv/4TySRB2aYu8nY/v8sm1KMv9ia
xDeW4xD/YCnZlrzPIFfc9uRIfgQ/Li4t5+MgLrE4oP7+iDaHdhe7UatNzHIO
lfwSt9m3d8kjvFdIVKRsk9TPNZk5lzoJVlIAb8t0M0obcofu3264Ab2wqP/6
i1jKzy5+/agBIYmz+3Ofr6Wg8QLsUCO9sVKHNqxLSoSeMuJVxQ5oh3SybMf1
pTqAe2Sn96TfiU/O03BlMUXcM7FUr28IgqLUJRreKrhs+G+FlMNZ/5i6TLk9
Y9pu/LF0oE8IhIIp1QY4TqfaNnIzuVWTgCFBq+YDRzeMHWXocxXklCVTA8HT
N9qYpomPMpgLHLpu52xS3JDd6OA+19AfhPzUzKWTPkovxekesunlvgA6Jxp6
/HgoYmCKvmjJpGoAIl/YznbIXMy5DS/yar5+7e/d9ISEgAS+pi+0SvCSohtQ
s9tib1pemuhdve64NRmsTBHFjsOYu80oRUSXeOzNl3b5iiw/t1QWyHqHsI7U
3UNicDjl6x8nY+QZb6pI5g8P0+uo2RsPULKmP8foRVTBrK98uSwvc94/y9As
t8eHge1Lu75yXu3ldcpQ2BuluhcJboo6wFLpjw6q7FSq6/XPdjPJzQeJamH+
z8IZ0OYAcltTS+/xyi3r0aKIDXw9GGI/fUwrYlhtSVBLjgakp6QIpf7NfJRj
RK00fS7ZeH9Cip8HbPUrHkQsC/QaNXKhBdSxjclYkWde+uyraZmyhRSP/rT4
hEfwBGuObv8hK8u57Uwwbu66fWAI0i/ncclfhaJU/gCoO0mNhmOo3kE+j3eY
HDyL4pYig3mZE0y26pP50TtvlIPmVqy3DOMmMEqpFl49i1zL6VIwx4W3Ebqk
JjMLjNIfkSqQmbJtDhbJTj0C58oYbhT0IwRDLUuYzhjtcrzvTudVkY8bqLpV
fETMPSq79FylR+xycwEeuFQUV7DK3tiEBBDLRgVJ4MsSbn8bZoepjwf967mL
BQZtaZ/WJ2zihljmXizMp0nC9w455ST+fO/USGS7ofD5P8YZorJRRJARGkRu
5rhXSOu6qP9ivsKORG/jLQg6MBOxCyPBKPN/iw1FzTdgUXBl38p2R9T7Jwqe
Vg1QITsvsefaIlzt9EtVHwf6PmGw4xR/jBdmV8UvVGBiAR5Zk13gHphvLmeu
1hLaNrtp60ACQSc3P29r1larNa3R/aoDvnqDQ08o+H9OJacmjMQHIdo6hb5P
V2kkVcEx9/cNOThulljMUROyme/39iYRnqL+tDmsO3juDjxd6hp/o8bffzeI
Yyrou8MIOIkhi+kEfsK8miebEMhkKVPWajcAM6irb/6Z5pJ+sZUFbXsbqWAA
AuYvo6rx3Jacooxq6W8wIO/l3jz1hGayqjg0ipwCb8upIRvSZx8yU4H47qfa
q/FpDGCYFfMOhHq6RDbKRUXpCEl8cFgtdcZaN1TjwmJ+fbO74W1FxrsZLt7G
upwk/+2PgzLajJ10SbYLWPhsjQP3trDW0G7P2nNq8FIMi5a3Z0ZJc8/TLJxC
5FN2jePlHXZrCI3WNpjC0x5TPYyqFVpqyoxHE/pATviEr0+j1tTzkXTm1Tvq
H8mTQPVYNGbPw6BJNWbfVq6uM2hSXvwnj4PJHaSHYaj357nBIlX4OLqJaBTN
HR7dhFyPJrU5bQIKoY4CK5Px/h6bJr0enGgLQ7VJzLNvZ2yVum79Xxbr1FPw
eg6zUNhmwtr/iSGTV78ijofUBRk5hjBX5XLTdF4TcrdlJg3JtBknBQQPduEP
G49AKNU40dVC/19EcffG37jhJZItcrcf7bAB+0vBmo6AqkE7Ws8GwJJ92Koz
m+G7lNRfAdTFbzKZZag2Lnn6kPqXtM6q2BmuzaxYr9dEXEMm9Wve7vCdPn7t
ju3FsLvKIR06NHZx3kwCc3UZO1v34z1FPH9/0tnM/jcRNparK+0yoGVJkMVr
nbGkfmSUxLj8j8xN7+MhFC2zD8lliApfH84qbruZCYKSjKlrEBZYeofKC6pp
0ltSkemsYS7p9YFRwQnbWktIfZL3HLBhuN4CSloQ1u9jKyp5y4g1Tn4nghXx
Y4wpGvxSmrYmgvePmfPqJpT+luLtDCulFuPMf3OnubRL2yGmGqnJhnkaY7IW
s72SDsCL9HD8TI2/fmd9vLjrjT0thW0gRl/aYcX9HwJBXgewK7dbs00qgpyb
KQcqyixnsMd2vVdSbypFWfqH0cVWwe0p6zNKqh1Hxi0xqk18f6LIl4S1Nb7i
IajAiZcfunrh31XSvFYGoyrotKlbe6DGecHRevUf25xTXpW13MV97Ym0VJMg
pdvMdy+nCPzfZmYtrWC9IOS7iHIWM7KMoNS47qWap5XfS5Mn9cuMMXPIRz8d
5/v1l8+6fmlDXiNimGCRg0OCmltnxsiRIb2eqs3t4eFBOxlaLGiKAQS8y7Nl
YUrmDR/cIxiy/tF4S6Z0iJkZZ3EB/66CwxMfLjbTKHn1Cwbh2SCoypcSyhE4
k6ID8AD+duYexzIfHyAWOHGKlkRRlNnbPbiUB456e8vDS9juICKq26bsXgRF
0ijTAPElXn8u6/B7ByMQ9UnXInoQCUadFTnsCfLjdy8kLZ+/ryIEpK7m+ZBY
moCJCqtAwGU8vOFjKMRxlPBnv5jVSU0tSL+bsB8+cvdPb2SoBPZx9i42FGGb
n19i+5xSAVUyvM2Z7vRQcZ1e0u2h9qqe1qfo1itAH3iNhWwMkCRP6jdbxyAW
Qk0GvFkCG8S1VL/uUonPwAzuNFSPZH9dqgvKcn5Uep5ArTIBAqp4FAZqcU7q
GcKlljIp/cDAKcIWp+hRu7f3yyELjAyiEDGl0TPR7qqD/YJiZPGbMZbqtNu1
WR3Ixr8IffN3aEr+J/zLmxHAoRg10qVCnQI/t4R7FcictzEF9rkqxq9mWl3Y
9Vc2ZhkPwCnXsr1XUnkuTWFFicZo6wzuOTLWIgx3WKihCnUBBW1318b0fj3P
kO1245d+NIfAPFeZeEA3nh6yAnpKhHTi5lEYvA0xZU1bggl8OW85teaQbBlX
EUVVSrBHEtyux2Y1rLcas+jgkJzFVGBSxaRJyj/hClA8kyNIbdJ2bvmXFUS5
KljrapcjCoLjC8kHry2p44uYtdsuyaeqUuKuopCR+5xJ0D9iVAYN7ddcm0SP
Btl+c1sb4enEUnpewTW8SkmUXVeNRmEGNnMsXyp89iKDP1ymsMZVQJQYqGlK
Bx1vz+pxj9/L2a91bCOCI9lTRMtuKHn9Rl93T7JK5G3wUqV7rH+Xen9ESI9x
usM/XNFjUAR3fk2K7Dq6Czf6QGoFDJni+roJWwlJlDI+KtaVdso3pgMecuhC
6BCk3+gjTj4SO5qU/AZ8q8ugKjplUTVwRMyPLASwT2tVsvOnkL45qqVZldzU
Py9PWx4p7/ymbDy9qhyeIQ1F19pnLnTrUQwNdaKFpa6lMlH3fnOhtnoIWEXl
lDTfD/0V7O1La0ffaW17xA4T0nVf26SxNJRpFo87iALruWL78KfwdkWnBIOL
ztWmZlkxo4ygzDrphBIHOwaP1QNt+ckHpntwiSI7RMt7j6m8auZrRj2Vmfth
XX3yduoO43BzpBV/O7oxl06/ag20FKoC60PIx5nzW+nz5EW5LQjQdy3gjRcI
ulRAOuKXR0drXcPvtU4eCWT3362TgGl7zZ+5WYShPO4PjwRkFlPdC3KrMvoi
fVZJhnnTQCeTKFKkEfm+URYXGLPfiC+vAykPNrpz+w4C+A9bpo3g1tE0ORnm
f56H1IrkTxYBqu9024/oKScTJZGWVGGKRvs5m10hFDyUoCZqm3dcxBpCDNIO
c6i0H7chZ4GIOpY7VF3t+LzBubCyK2zp35CaHhaU5LYXwzVIwWO4pQ9FCQJH
5p78Oqa0lVD/+GIvRxD4wXF8wxIA82FXExk3GB7FGtUxNAzXi9BPBYnSLldi
agoHfq4F9O/RffFXboFL8eDxw2nUowYqKsP3wr30EB7caXUDurE9DA0/Is+S
tYJoN+SSZvSLtidRu1mAPrLk9U3+cXs68FxsQVNwHPui0+nxYoBqC3ltxRwo
0v/Dnkpym4952it+cw1RKMl43VsXMLqqFiwnDb3kou2e3axGoixU9ZnswlTO
ho+jSinS/BDopiwVr0K3EqFJWHkVsm98VF6EEt0bY2K5RJ6m/ShFXh061byM
/0NVkTOdt3tvpzCPof1hJn/qLNBQgoUcOTeIqQxtrE9KFtCGbt7MUniNuMlF
8sHZfkY/mzzhq2/Gew+86UVo9HIa+/pyrQHUdGFWlodvUXqlF7iDPbQr0lHO
Wz9xgl6OSDNJEz8QAxqEEzq6U8obf64dVmFy3m/fB6YNTmGezmwPPZPGAvK7
dPxqzcko/huQoT07SOE7Zhi1f6DSGmgkmPipw+wgns+U8TbsLEUShmTTbCww
jdcP/0f7r3YATlPttzzEHCIn0PBdBsX4XmtJQBhvdmjZ0s+p8o61iejO8NWR
lAtHmfFGeFa8/4GQ7Jc3flwojxFfBilh2tMNEpyxBwkjV8c7zfeMi/7eE+DN
3pAr68w9d9/kBdWfKLw0gVs7+ptgSSrWZmf+czy2OsIpOhsAchztm7JFxMce
dPx9/SXLxTokElTJvK/J24VkaFlApHh3XyqHvtwFgrWjgVMpzyBKhyR6UoVq
LcqVhIwHG5Jc2HkmdJA9CgKIaUlL/XaXDx24v6GZioNpPw87raRlYtG337Db
xwM2r/yh25BiSZaHLga2JDubABgwp63q150S89dB7AANzA7za8giYxAPJI5n
jPamqemZRTLNbyZOFmXnd9kwqYXahCirBqoGlLDWP4N+nozsbegTftVOSzmf
eBA+TD3Lj2EK58J/mJgSUStNR6DDvf4atEjL76veuyFDH3yCHG8f8wle7HFI
HsnrScjmNt/aDN4KD5/axgTAWmIH8ckKeV+/+pWtwGrhkT+BHjgoPsRXZBh4
G3TT1Vn37VhOc2pZQugShXGL/7/ODP2XpoVBevi6KfpNYpH0oT7q1w4ZW3Fr
2orr/Z6nWcPU1XObS2I3Pgy1tX8eujs9+jb5Sdlq6uSqk2FABbC2y1mrj/y+
dQ60q/4MS8lagEHjyVb9i7emNdU8ybyBQDRsFxfZahNYM+37i45l4GTfCI0c
E0E2U/qq2CUFp01x65cARUdKnszgtQrMtdgzFAZLBIqTJxz/Z80Qgqswx2d/
wfntagj4HPWkUVj2cB+LSfn02aYj463dM0zO8tdFlutBY8s7tozJ2WGQtP62
0ZI1SSt3wrFX6Gu7dpY1pd1lQh5qe5T4dhdijXLaRaoJgljcUjTW3itfnwzO
LELsY0pFKrPEA621Kx2HX+MBYgGeIjNfpJMrTGWjTkuCrFFqwjggBow2fFq8
vCNB2DIjtVdqYoANAR5bbmWfb0lR1JEjyLpYk8q8zzXOUiQgUVY89sWY3b5W
LeOULeXI6DeEU/yMLortX1/SnG9GQxQ7E5lShEuRk/zJogDBMmQGR8eWzFcl
FzbGJS3S240/EhDWyrQwGPDQuOAJSKieg+WKfAR1uLci44QjHEMBkKraKh21
6BSnpAEFvl7JBXoP7YOGMIp+RL6nyS7R/OHEJMQLramX4G4s5nKpFigCksA9
MWHSWhU2QwZJ20jZVrPVEfxvJjiV7y9jPXUDVWYel4Iuh6hauiUMGItEzzC3
i9hPhRKsk4RCN07bFMZi0Ho+TNMtQlwbJ5oZ81BQW2eV8nnDdcIrqMjdYW41
rxnTc+yErdvnJdNd1JZZypyecB5Qu0OK8pROkRqYBbW07y4OEMzRYnZPUmYB
yGLsow0QQGhT19qFp4OR9soAh73YoEEbEiQTNHq54HkgzE1UdGlVK6pOUnTS
ZUYA1gO77VNamEL8QelFsEm99Lm3vq7y7HVEuV0hdQslAVX0p6Hb2Eg2/iON
wWWfEhvGI5lyWAcaLNOhzColgUgey3Z33h/bzGZB8PV8VeoZKNksxBVb21MU
ncBlM3OnUg91bwet21e14ksXyFem0hQkpYZ28oJjz5r2LLOIMgXipHCItZzj
9Tban+T3tCdC/NnOVeNNYIdYOPS5d67/8l7L58O3iQ1X9crL95DmnHhHdMRZ
CXKqvuk7ApzhVBPMhWLIO2lqQKPkxKFj6jjHyjIPDVVr0eKlpRqD1WCXOXV3
GP1sBonlWVsdB7h61E9eLly+4RxiwGqIbi+OQOFLlLYGG+vbOZoldapuHKhm
+WKPPc/23HCBiIEENr7j9WzP6TzPQQKYNpFyeaEp0D9Ubbm8vKL4DOCB3iyl
iinub77loy8yCgKOws7EtXEte2w8y78JSXidhHw//2aKqSoE0kprsA/+T9y7
1FoqanNhOLjipzIYo/QvDzkYl244JBdrvXevmpKpSsmslQHZyEaoOO9aCYXi
aipMJiCZ+jjLADD/OcndLdgPOxy8v1Oiq9oSiKCz6q67Iebnq6QRAWJ/rHDB
WaufAOZEPFmxYB9Jn9EV/oGOlrY9Fxis57b5yT9AIkUj7wWvjGt+D2yCEMkC
6Wgc7qEWexRKFlJd/se3jnjhUzSrIiHZQEujsD3CMVHkjP0tGoH2MM7gPMp2
2n57Cf0o30bqu+Eb7nsUDPsMvytpCjjtxXeVKGzkIg0T4EtYCefzZ6IkWTBm
xH+v6oi7TR0efm5+DZxwZI2gqQKwK97m8xvj6c4hNCZ+5v/cQvD/siO9G/gI
99EomKtVrqyIA9T3L2lEABu3n5e03gzkZ6s7i+78Qqj+J/J0TjfDG1c7iWSE
OfuKW5FL5pq+8KhtGAvDfOlARuGy/fHsUi/h54ZnXj3C/VdnXP0PcojXZQC5
ehbUdLZc4JvDIULExd5J+c8Xe/BfzDjHcg9f8EmI9x+f97QKy1fzl0pEmVxR
YeO/1A+Y9rwGCTrL/nOAV4GQxfvs2eY6Q58xJeIYXcAVw2vsyCEEVMlZM5st
Bu8UfPkOgaeC55FqWpQw3pGVkcCZI1lZfnG+otBu5mNyItaB5Y+nkGD1U3zK
6vaA+DSXpUcfAuMRTI69IZ+IOMKNKxlK59IZCBB2bWJgcsWE5qQCrKeGqhAH
KEpVJ//sSitGjCFeVKXGit8DPccW9rjuhSi2y1gCRErflIXrVG9I2xsrX4XU
s358A02CDHKxCMt6votrKXap5tlZzIp17bnADR5LuqszEyHvEztz29m21zNo
egB4LuTCQjAHYRoFasKcAwbE2Pf+/p7Un/KWMM/oeYgqKWrjv7mXM/1P4I71
YQxFoNe1EJxzdU/vSzN8EY80suqBrHOJR2MZTef0Xr5p7sRF4fax1B2bw+7u
sKpDKUfTz0bDlyBTQd49YRf3w9idnRTVWw3rCV0F7nDAccuKj+gdsoqJTwre
0ZrkSy0ao9/SP1heeB1l4u0fZCMxsQ5QroT2eMUYyIr7vc0vG1BKXjcDM9hj
G2mMnJ4MKeNcCBUdO6IpfeHBYTlGpPN+ozEKOro6ZtXAACxOUx9C+dhAFi5V
22rEQlCfQMt0ZhsvUJW+oVAOeOhAQ5+SKz95ABodiV5JXhtXiWscyx5Tm2y5
Y4Xft6SUMcouyvTab58ZC5GFiq5gNLgx2fP/45XKjJUvx7zyI13i0FDN/3/0
V70N/ITDf60/tzwCMiT3zM/qMLBaYlCVXZdBsGraAU9TqtZIEkXZgX/VW9sl
598O14B3WSuPZUQjUex0STV3itLrNN/FVKTm0Zz9q9ZRYdQBCemrgSyh8zkN
QJcdAdmgF7sBlnf6TmBGVELUiLj+Y6z/P7b8tWnflcstds0a7FKttSjmiCTP
6JCslKCczblvPwL5ezGVOO9XpmAa+tK+9kcagd1S4Ui1i8yNd5ajaPbOT6Oe
rN2QpojXRDckablY/dURikjYfUjZX0IH8gvkFER/RF/D4jq5BCshMjiIzKD8
EPATSd0tG5uiduJSXD18LbcLjvvaExmdxRm4fNWXYW1B15r10+Gp6UVvZdPX
+huaJs5v9eS+bqt0wuayE59f2MazDqrovePY7qm2fsVB51xI4TMkD2XRUbMu
k9vyzGhtAWIUV50dI4zKw7VBR9v39J9wAKXKNhiTbBu3w+RzgWhNokgPsBMe
O+3XbWDnzr8kN1AyY5HSoaqQab9h6/D7jtls0L1SXrO2btQ2RsaBfNTlItyo
sE2VeW0hkpy9/Nky4Nsb4xes8fdqhKkE0TPatzGPgYqeA3v0rHJgRv2WfAEY
aCKH4DG5y85TcqaMaIvEskwAzeHXkytljHg5Xz7LBbLQy/k1HxQrTuQRxxqW
ojUNQd8XY8zLQBdfoRBc4/Uon8gkRplhuMdTYAjzgzqXFuQxdokan9HmuMN8
SrfM2U2GfnKvqiM7GI+QwW6JVb7Xhw7kQLz/lz25JS/7Gc00r8PLQ5Sl9VtA
DmWEcVcmGG25f565HP+sbc+b0u1vhWeNuWPSgDYzBW0IKMY1pyLeNdTNny+S
sKFNXsZMjWipyOs/1bmFYOovrxrgiCAxqKReC2EBXMp0YbQGY9Z4IwlvMVbG
mjfDw1oNjgHaUYJayUDG030WzZZXW/Q54vH4Uge2MD5h73MM1PVc1y2Ba641
AbsPSMT39mmyyZpvRT8FqdSMexD29JW09dMDHq6pzFYNeX4CLhuIR/ePHJqX
0RjY2UBhIpmfdO19hUiT8K1z4Jg/+j4b40UfAdj7DAOiGECaYXSf54ip4IaL
LWmg0mbSh1aaRIiRo4N0An+kRURxPHbM39L2wgr67I2KtDg7eKPtL3EQF+3F
a2aeCXUfr2z5DJUXkta8SpcEdRPrwBWXSEhtFVrd5+9a2UGfZCfGDietF/55
GUtgb7ebhw/e+u9UZXxB7I56xo07DPWFzp7t6L65+RvEn/QbtTXg0B5IdVAy
iLJ/oH90GmiKojnBfmc4JUTW0SYphLVyF9qoVyeTmlwF6Pm5K8YrPvskuOk9
2fSkiFVtdU8WctnvgbCRvNmphcDvFjKkLF+3c3DYmyNexz0LdOBy79oDiHh8
RSil6+2X/hFa6VCaHv5nXCrrOu/58dzUE7f5q/XqzLuiNdVOJO3TYG92+sDN
Eq2UihKDuiL3AychglTlno5VCeZ2bho+IwXZ1MB7mZpnarlklcn4hc5hy8eh
EvGLlViEIguLVblK4+L3K/yHi7vppgli1qgrnMcBwj2g0/Gnq+/OBnQKCyJL
f1anuzu3rEUzRB+IO48witzyc3b5i6bMGazf4wi7UHtRjjrbPyxcTHzj3VYe
rWVd+Ao+mOMJscxeFN+I0DZaDt+lzHtEKzEtjfP44sfnV57UhpdMWaIR3gXx
o3SnxwkqPms7a73KjuzcRsmsIfGjc/Qc+AvrLP72JrQg1IJettnwxEUDTTBU
eX1xK77DHB9CieoJX23+d/8EpwPkeinRSsHf2P5W3br78DWDN/JdL2q723jD
goFLWy1BHQjV5qDZyEc+WODU3HQiYjPl7cJtZWoIp2ju+vKNmE6Bz49BJxf1
b9vaSPliTYE9ulmioxYkD2R/foE+cz2dwWSYQ5wDUJw++h9TlKKOqsKhqsET
skZMgSBuECs2U3z/8bE3jiedzo39YetQX+lkPBy2CMLjposslxBHzARU9pQ/
THjIPaP2egftfxhfYnFvhUzXPKckoICq96EKq1jU9Fi7J4wrDiYLGUnDrXe9
+E17XG3+XyJPnVCB/heifYc7JWt0G7sMfJraKhaEyCp31KgDR53+tWbnu1fD
U+mGAHYOqxYJGFMS2QKQE9EYlm53eqkrDtt74dN8NCZKLVr1OsHXFbPnsAin
X3H/1ZN5lhQbU8BZnNSkGHh88Eocu4nA2ZP3qFGGn/uMFGdUvOsqck8fve84
rzqEvpDXkPuii/sxnZtn0ssj0uPN6K07SpGy3Q0JEEzsRAabO6Xd9nFHK+8o
c7xNxVu3Vgi8CBDst0pUn4nZGg+I1FZ+upZFMxS6/MdPPPC1tKP1I18P3Sj9
+xupywSTDDRd+Khn+lq32IyvD13IlOxzYRZHOcnwWWDBctqSc7WImYdykGAL
ar8ERDBwFvboJt1fbmaJz1hu+FiZ3w/dgiJ2ICCMvjJfCu2trhdpLSZmdws9
VDLqqcYB5TWe/BiWp48nD6oNAnxxoJzFLVAmRmNvs7IkrpPgtbKGdTc08Vb5
oaXZU92YLsutXKEfce7C7T8hxF5aOPR+icaJOOCh9YbRsGk8k66u2FPUeTPN
J38kpQub1ncwk+7rzKG/ECZoNTdzOYr5C4ixlbF9F4xJe2CIZjTE7U7ow42x
Z/I85UftrJESoEccQk3LC2qVmcL4qKbgC/E5/OFWW+azThmyKLMYwUYKc0aV
cWiMsAVHJCCidA7qM9ohDEqWHUB9L5S/LDDCiWHG6J70Sfze2G53zULcqeIX
0ONgxa++ippx1yUHzGSb4SkEDyXe91B2oT/bAy65+fUsvPzY2FMHd3GzG6ZX
D34tXfps+WHSw2XFNhNNGeVbjvWwPr+okdvtBCdF3ua1OnP2MD5hqsNYVNw4
/fNJ83rTrdN1QdL3AjR3aQ3z32U8Y44sFmUfDD9urEPdpmDMh5hS+z3qaqbo
1qnSYoW9GMUZhzD8cA1DO4XQgVxSwKiUqOPftAEEYUHsTtMJm4OuwBrs9uxd
vQaDYSTdYz3uPjeQdasmPXeyIQCTYtSJ1ShjQNh1Cu4aN0UsHvPEDO8DJD3U
BVDUp2L17AZ8uphhiqHLzw7swT8Avnehoe1ITbyULhY/P6ihVsT/FeqpcA0x
Iy/xFlnkHRD8YqYJPAnLC1j1iKn+TdiZ+MWxZmj3QmIIscwzdfpZE2x+xTc0
/nqMg97+mHpUQR5e44HUDlRg/R2K9lmab2HB9k1d+aKyghCUJEKD1ICzFd6c
OH9QNNguPAtMtWVJ5efKPnKLk6XGctVn3bCQvJEp9dIPaC0fEPo25BDwutKi
wzG7pSQcgFD9LBCbqdxdiM/ocw2oR44qvHYPt1O0jQ4rPLPe2UFtCHVcJctM
eKKVkeGhkK2AXtAOGOqT2lyswqiAYNAF6in8mEIG7hZ/rHeu+MaaAEaeOa1u
6J5vyldkUzGA4OxRMok8gHNVdwlsO3G/CdqzDw+p0YVp/rCYNLkdl1J5dk0V
/C3ZNweD62qARNCjXCMDRU+6zGXWJkHFMV/S5MAL///EbiUGoNbgNX31I/+e
er7A5ABtJP0EuBDTUNkDlNj8FwjrGvfqg3sXl/NDM/uK0eLA/eta1N9oAemH
fNjaNn2vxxV9aR+9Vcq0XfJ9KA+rF+sJZUImbO21QPFas/18lbFcHGCm1cw9
ITuEi+C4FN2YBDgZYGEUNEWRCxvxksaWp48EgB7ypGDIVL+3OOHOFawQvRNO
9CyDdh34Vz546olscJH4gL9Se5ufgzlBClJFKBj3p12d0BNnh3g6rLRJsOM5
dcoUKfmteb/tSC6IfuSZVcgdfrOLAShv+8VMHKSqEmobOL59g74KABqdhciS
5I/6lBMJsL+xmWDTDXLlmxBH461uR+HMFRcU3wptWjBbrpGrGRmyDwZjVrTF
M6XJZFOV4c+oQZ7SqGRVSwbssEkkKsBuP0aO8XpP/6lp4PwdpcTwKiRtWcpj
6zxNpWxRhkAXi0rAXxZ3qyi+2QfPS8T6CxSZ1aCQVa0wbdPrTlJmj7IM3FcM
2DeQ90B3sMMteu4s+1mVM2ovaQfaaTxpLsszQjZRyVDFOi0RxST/XtUrsoQJ
QnnkZB4CqKjpHxEYzaD1wdSY9d5s+czN7eeantrnpGBDxMjltMb8aw+MZSMi
P2505/CGiM7bzLaZNHfxtFxW5/wHPo3xd38RMCUsXqoMtTBmOH50d97+Qxc5
iQHVDVPaooj6TgKaj2mf7LqVt5oozc1LRMPTdAO5Nj88t7z1B5HR0w4JlLSS
6KAQIRA/jeNkS1a1ceIW1yDlrHuPLeAi/3okcdC0vzmRie4rYbNXf3YsgbpJ
Wm8MtL5c2pZQS8RYNK3hZXvT8vtmGL8alsgqD4qsOhpvOQJFhOPnoPihzdMn
JqExR+4fBocMbsaDXZRQQn0Ms6+6uSwS1ZaweCuDw+WhSp9zEnQnV4ahivOq
M9xXUf5gfqnJrFePEIUKoiKCo/qVvxmKoaAPyagSvIFRAuyqXYAIae1nUM/v
9rqZByIJRaQizXaWMWu94kvOklVMEZW6HjmnaGCWg//q1tf/FRXUe0keNZzD
wVfM0XNvPjQuY0ZpLRQU2iVMN10Re4wYVM+q9a4Bqtzqea4u4aV53knYJY0i
VqI02uQNapjv9IizQYWCNVzaUqK/S2aNsH+Iv7d/U/e4tub1c2mubBPfnNNF
yi0qqdV8+DEI+M3OCqhn62SLsUgIwP6CK1eBWg/SKvA4lk6O1h0cNgSndVGm
rRVpyBnTMTRnyD3MNU0xfmpIiPXEiFslDngQ4KDUo+vjn6XTMfnYw9eQ1RMW
4i5N9JX4seZZryjJu/tUBMyfk5o9xYwDZdakFDS264T0TBSRzsbs/frwGiwz
3Xg+yTSmEtrqJbOC3IKT9ughqFzIh7Ewoq42/44fuUGvj5oFet6AHFUw+hFe
JklpUDjpqFHGSuVYVQoNL1xXPV/+0uq4xHuTcMwwH9bqb7odjq9guOLqPfE9
va2InSNOfiXUdMPkNcKqANQBctlJkJtKfHeKcOKBvJD1luL5ngkkV2AoM9fn
vHV5tUE99jZE+qFg0I4u+m265PMdxtE/LChGytmJ2Ne0wuWp4v4Ij4wa+N1q
RXaTCAoFNz/IcCaCgFltQQXJjs1uLtNg8G0gLwR0rJWeeikU98VAh6UyykVD
eQMOlzHuRMpuLjFDCFRcfF4Q2DH8WAkaYTV2K4fJKxwEUhEBt30ozUdL/hHW
IYcabOluuTOlTOlHlappyh9LzddFquZ+anbDtkfN8RCv9YVgDlTSKXJ5kbm3
A5MXeOZRj4obg9fyLKMR4IA6ZUK+U0umwtlKpfUzOrk6AZ/r+IYqneuGycRM
TkI4gUjRDnk9IRW5xjFUnKM0hhRGhPC0aMqlEUwo8oyTtSxvmITBlR63JGz+
colbwPXIvpHA9IIZCPF15IdXx9/wac3/t6wUyoflDUw4TEFVt0arfq1pvVCI
ssNwJasBi3CGSHDB2pdL1cuHeBSgjxSS0XHMDb8wRh5ssvyDDWsl6WNfn2Xs
F88773gzYAVZPy+yDvMBZxOz29sLqtBzuMO8AgPrxXdqVn0tB0vr2qi1ea5L
KAZtAkI0eRIZPAgfkFKRvP/ouxN47dLWbZqnOiWaM8E+dRDUITGczLpR2OI9
KI6XQIdHSf1t+cOtLnPtu4e4T8IIKE0HJE4Ylgf5PyNCSA9KadXwOz9SdQCw
ZEFxOULhJnIxfyW34kn+97TMqKQEdU/DKIzDrapw3W2gQtCypHxeM/Q3bkQF
PqDaDv4qn9a/tWjZRAgjxUI9sc4AeQaf9XO61DMMDZmvRNcQVRjVWtR5/PHt
h1qoLRWG9mJOdBAfwWhvll3Ru9sJ5DdeRu4BK9Fh6iw/HMixoyIDjmS7mxI9
cH+y9vW2OfaXFUSNJzqCYJXWvJ0bsggiI/+koLPOJnV0C4ho1FHRY9XKmTWR
kTXvN7SvIUBiPL8HmWlUJVuGwz5nT4dZO0Z3UQ1ZPpFa1jI850KlUSVwZiFz
0+Kl+Uyxq75ltRf2azxl+H9ky0Wf6jpQrf5s9YspBbbbvheXiHi7PJTSCQc0
w1DbUsu33Y2e1e9H7FCpjyhKcVXql15rG/MhiW5rCbDNDMl2WC96GxvH7aKv
OGO2otH3nZ8ppkpMaVy6a2m9TyTYDc2Hr7KqWBx4z2ysk2Z4G++arTRxv6EN
+GbIFskmVkTBDkiQj21RRgb2/b9xRJIETZSI7IFukvwoHPhPV7p4PR9iQ2vn
oR/bJkP15iLaSpxsoQRlY90ZSHz3Fs/2gzdrLswS8dZSlpBOT0m84QDa+EJ3
wWQxtxmMDX/sakLSid8XaZ+BrJesOa/Iy44VtE6zmr1PDGM1qqpxoxlFP0yK
PVVJ98I9p9Sgeqj7LMay5Jd+1d7rfk59Ch27jyRJl7PMLCSlbkdvoIGbMqQs
Q58pGBJZPuuTn33CHBp2OiPm3LZe86UVjsuTluVVRMEmExpoa2cyHBTq0RrF
7scIRyrIYrHY3TbJh+2Onqp7YST+CmeCdHRJlDy59/Xfa5Mpe/poiCDjc1JV
5G6FqS2YGS7GC/sbYAX9ug4+s13a1AwnQSY4aQc0tvNSA2ACuEUIWYQ3mG2F
L/hV1QONB2mm8D1LovkLZzC7iP5I9KaruZRxPJKDxew9/fqRkhQGOC5BezgN
2IhFKgJnPDKnSlbgMJWPgSbTcVOnaOyhQwsc/OvDK7vWwzx42b4nVhJpBdes
fLOu0K/53Px7Wti7uSkxjRDQJ2rgBKlQVtOPm2mgWSp/+NNJezgd1zVDAkX6
0A/IHXT69PpIVt7/hQsWCmXGnAyW1v8EcA4TMrkkmkQZCAOzh+buaB9QFA3k
EpBuEsEC2Aflyk7MSN94+rWOA8u+GHM1KXCnxg+ySRFWAy3QZDJ2g0l9RoDS
Pea7NesfKfKCcl3h1NPKyzwYKZU2RHefRLQfas1Lba0OMp0C4WJ1MOOpSM1B
gm3lceo/2R/sTUdPZ+YC+X8msJy8KlY3vkRmjH+D6DbvysJ+xH6YABRzB8kR
OflLZRbSTaOJOphx1BdtrqgSrRtEOrEDNb/OhMVJKykZFo/syhJLc7yk6H+y
XcCFWBeZ8/96Tm8toak+60QFM/qxjjAaAYt3Ya9Jtq4rGpZusfX1il3sPitG
5DBVmVx48YkFFJtOn8wsDq/k85vMBMcgsDcZmhcpPBBLIVf8I3n9PtfYeSAA
fbSsYrf4r2xY39HwFFF5R6ntmqBERCipljvVre7mBPpsFTeACvYAI8L5v62H
ZLeB3l+1ne8eTb3Z0xg4CI53U1R/gRKx9KFeHUGX1PzB7Mkv28Hq7YlklW0w
w6CzUOEd8gLWJZyw5LacsCJCaEvFzaoh6v+FZxbkwrFOyVIo3D6H1T3d37KG
11rPtxkpKhRDqSXXNgN4BRm2iA+mWEhIp1HYD/3Y8847o5ESndovsvkUR+nN
4T+nabvfwhVzKEhh31IDzaCR3B2Z1+Kchg82ePsnF2r+5CDT+SomHQs05Ab7
nGDFPg2xqgzbwjCH7+K/ZwX4BSs+7Ycq+5eKr0H/JvmD6lKQLyg9d8/37aSm
8gshvwG9lPI5b97BIF0JwAaXEJMiQ0pXATS5fwrp0fUmV0wX/oxRa4/lEn8H
PFAVm+81sFnurb6wRe9gBXZ5rxxpH86ovcuOtqbPWEseW2GnRM2ZWShR1Vxc
uh9xZtowLOZPK20NqdD0nPhM9kT7BXgQjqkbPrOcsgo46Fswokxoz1EVobks
DEj3/a/hmLRcviWGJll1TfRicCGYroR7FZ7sdWNdLaQdk3Qfh9NsCFOuZm20
rYAwSRy3MO2yV3PZMnIu3s6r9AkJsbxfG1Mq5GZK5xjqlW4IJVRLkdvVTXIJ
xRvgvVpDNIYH91VOedmL6fPjHWxeLZzuzmTXIUfzfG7pk4vJ8/CoA9POaRBw
382uMBS2kO+psP/OFPf7DLyHJA+Fb9pkfpOKC/Cf969UUu1jWJWzvN2kEgLF
YNrgdev14XPSDYdwMRGFimOK99V5RnnrvrUKgSSvAvXpXo9O+vWNdLyaodPX
P7SG2Cf59mP17+hNlmfRs5IrtwlhwCYx9HA8ICFDnCDQ7ifrWKPi75vqbIVP
4x9dUBmFhYGzOLE8OVIuqhVwVM/cVBxtB9KDhXxFwALMupf6dVcghbAaVF0O
4zQ8kwI1WqkfFpHJ1pKB08HfAibto7X6pFRKdnCbvv23Y9jA3VbmHTaqwSUt
GR6pHTn/Nz9XE5DApYLXF7ON29U3+4fEp3CQUBOHwdaPa/5zedYLpbvnSo+3
v12SGCYkFwVDbT9/sFIJULxz2VKaLhb03PnSbah0+MQQ1gMrvmFUDpoYlVR8
SuJYvdQYuZUPMzCKf8Cg+H2UDFtl8WRi7mx9p6qQvClLvoL7vcv/ArpsVSCg
07OP3m4T9FzZUMEuUoN73k2+kd8J6Uhj5kGRULg/O0eCOxUhdAhHrBXt63pm
Hjy7IUWJSAoIe7S6ZrZoR//e/Zw4ZUIS6kqhac+PEQHmlox6FZdh5GzvdDJM
J2XaMpUy24OkFKQ0VtfvPJfbWzsoOJwcaPr0vaFKvXaIs/xMDnblO4SIbLAU
jkqWrBKtltyZQ7Fp+mr5HHn5hle+u6X0AM0SOqoxMRq1vTIGwlMLLjNXGH+r
ef7vMQV47mPRBeJ+RQ5G2re5mNLMsySwsivAcUy5zTapEBNDpnZ6BGfSMf9Q
HHltF3ZVS59+uSm2Zht18NPIXEg6fw1g1ZRrhuQIK/A+5YL/UZE1MEjwqLef
Rm/4TUdCDVL5C8xcya2hUnVnfsytv+9JpqlYQYTn1jUiVCBsxaTstvDFgiB1
J820JfNnBYvkarN44uJs1zanprUvilcUMYB202ld996JM710/1w37MtcYJkF
rkbgtfi+p4EBFZNP7i/Rm3qgKIOGNk6KYRKai8mvWxF8E6z+WXYrOr9KbYFE
oYkzMgKJURjmu4cW6Y7HFWkqureYHzVsVDWXOUf2c2YysJ8zRW/WmowCJqdp
9g+hdkUZLc334gKk76YipIA8hDH5xZmDkyJMvgNKgkATeLqLKJJbTv8LocTS
ShatPXfTR4Dcf/DO6bmMJJwhDtFYc1SOWR5IwmgNEtyO3siRz80t4FN/lvQV
ZRzpSL5OfYzRS9WtxTX2gm6skCmVI5Oh1n7n57BWNPOONITskyuaYRz3neI6
yAN5Se0MPnfa+yCayj3sgSOgzLgxOaz9i9QeOHKLfKHuZrxPov6glyOEklg0
XqT456UedXISI2fT+/jGejj+TMSUfM3lDiK+rH8tA7lNW7ekeEywS+KNXCCP
YyvIO60hfebFNuWt287EpAuiFyQsr7/9CKaxBREijpB9+zv19iRKSrs6eGwq
B8tQGIuCVu93IF/ndgnWm1sq6RyxERt8s/cQibXyY1mmg3PtIA9tum4br9CT
jl0udbo0FikRGBNnNhDXDQt6L/8JOizzo2NFEQ8oLqMVv9OMnADzGiJTIRQz
bf1pcWHnTZnacirztDiW1HbxITTJE//L71eVFnz2KgVBeA/6mtUuHNHHibUI
TPsyOanMfSFG1r62CrK7bGIgtz/hgEqyD31Er5UKFok2pZoKi0g9o2huHBl9
T95NH/r2uDfOgB8vOc9Ow0mUqtpsiEqNC7FCKIknZ/fDamQdBYOjyKP20VeV
68zQEZo65QTncwz4kYruS324OzHjhk2VxaJTXRJLnnf5bwkNCcZpagf7SVoM
NE4ygJIUu8vFgZYgjeeVXNCSITLZWphQMUmX2v53RTSMoQSHpCleGRz1y66I
vZqJA3ZIVroMM8uUGUDTWuefQ6g/Qd5RacgFacAQnqwNxJ8YEmFXy2HOT1E2
OMGmpwwCK6MOKr3pU3oNiMu4fX7nXVysUuH4Qpps3Q7eM5IPlEEXYTzlxJMh
SnyscW+Y8j1HqS4lhUhz8RWVHsiH1+JFyVH6BNXfHvrR3zKO5//UAjsFY2zp
qG53a1Aj4ekfhTqqj5Cycom3IcfRNMWCvepiVXuA/IIoL61nmED2Vt96M84/
qMjI+kUbSDo8my14q4Q4IJ9tCh2uHamlbl9tMPTRTT1iYhIofylDN45Mv69F
HTEhZTXDAFO4+zyTFd2GVaUVolU4e7R+3f000DfNJeh5eCMs1r7mCgiLgIZE
pG5Ij+Oh2AwGMv+/rNzs13iIeFls51s3Q72e53sJOsx8rlCTSmgM/iSAvC57
Qxtg3wC3GE/KjQNsELAt5siOVBxxkQZSJYMSET38+k7B8E+FggXmP9zhLMw0
8AV90uf7TZ97GYASjzAO1qDbWZ2Yw/4GeNO8SfLB4X6fqNGbNc4066xPUT1U
HcwateDJSl0LjOddgezbMccOShL5x9iDxo7nBnvPxELo7PeU6oY4HlMOqQ1e
+1eWGl8EaS02TpwgDbr4l53K6U2ZBM6u4eiXPEW2TOKMq/H+0nsov8Cp/U/i
kx3iFF9u0pQHC0jKULLJFAtXcQIPL/gWXy9hD1g7C180pQ83dqkx+XW1YNvr
z9MxBJpQucbLpJTDAer+5N6BppPPBM/8Sk53yzkTk3M5ZyrIkZVdKA3FnkPH
HKkiC7s7kaI5G1ckyH+fH7UQeRdlU/2NoZKBc/C1fRmJ22nkCcPVcwx6Bw6L
yYvz9ekU8e36FtShtOupsanO/77acFWu5qS3pD9eEGKR7mjU+7EuCWPbyUDp
FNstSRzcCAQ5msEGNANYxBriNAsqRLeOv6RFc6XiTdgYHJU2Gz8QzdABvCGc
MtwaNe5ugeiGrQh18jtGGe3stDimTfVBS/J6SAWRazchyi6YI8ENgSg1ful1
S3XtiqPISg+S6daujQMb2Jhd0BIVYsXa8TVH+kn/pdcavKqP6erIur1e+VmQ
6vNtSjfw0ADi4KX2dCQoMVXcixVqYG9apyptsgtoVv7gfr3LiKJZQ6WdFHBG
sA4Y9nNCDnB4gaVHKqVtjH/96zFAO7EZeCyFqtmwciHTkKX0S0gMemT2B07l
Mam5BSdB9fjFz71G+u1w0g1optnFcUobXS9RrWty81Ejqc9VUEcUmm2UeF0l
NI1QKCmo44u35Nnc6ZXmV2yvNaNUAPAr5a+GTKHbG21h09Yn5+D23omjFPYs
QlAzf0/oIjmTWESFTBCjoH6OJM1RxA0/Ayt1S3tCTXyKNH7uNCadTJyHeteR
QTP0sRgIw0ocVENyJxvKaflPJ+fFfO7nSoBO+1NRRM52CbtnwgjZW/lznN4g
RPn0syyz7YDu+ZK7XzJ25m6y1ECL9nK0zk18EHl1QR9T1AAmhEocG+8nIHL6
D/bruS18wDBaHzREMe6bt8Y8TmK9wDDl98jHFinYt/RH61ROB26Su+iZSCT+
2sOD905WdnLS/MPSGaTyKbsmcS5ewi62WiN7xYSa4H0cF0TWZRE+o820lJRJ
rb2VwpjkmxUtwoPeXuGTKGpqCzrfP7Ib//JkkZL3dmz9+VS1G5xrSNc/3D3y
E7fp9xTU+W+OYgUYDACPaHpZ95v9CBoYIM2OnnEMdrGoyT7EWu9qwBGSyldY
Ru7FryYacnneed1rklhLlSfAXG80axs8PdJn/ANtDybBmj6Z3KZKAdJ8tiso
OY0D3TKnE6XX/yI8+p7d9mgONF94ckWTACSPDyg+FtpNPUsnIfwSfD2tTYS5
cayLU8pn6tVAgIuNN6Gw0TuoyWKIXWNAAuGqMdDzo8uHGHQpqeep7zEUw/6x
+jWH4x6QOrGcxgT04usYpwMZETYedpOpUGaAcmCetPWDH4A8VuJgkBOLcXHR
ULBHOru8HhLXgWAdOCxMa8rmecTMvpCYQ5gKhv8IsepyjmTZtYL5rdwEwV6w
0+3xEwyed7j/GTeP2Rh56cpXd1YGZow7W2DuLoeDccm8AgxVVMNioH0zfAGP
U2VkDDP4sCluPqrLphKPBEtArGxm8fq+v+iy2vLgedQetD+4wUucMiMmDkn6
9b4euL9KwGdcSIdFVZYnltV84/k6QRbHEC3pTD7QHwMDSpa73VY02f9bjCFU
2zNnZC96R3vqG1htwmQ/MisdaeZ/3hqbFXmt6gTTuqK8LRvQZWgsKH0q4cQw
rON8B/tBl7l2pOqyLB8EP0EUO0FQyCMODNJc5Y9dGANuCGMLcI27+TUoEiDu
txjmt57x7viCz3U4jRCyiLnI2Qn4Wltf/XMFZNR8xSvDlrhqa+lB7DGw9aa7
m4Yg4v1uN2ZR/x/7gvAxZ30upFpeBQ83AhgRg5pDhHBf+Yv0HnzDOhhtE9l0
KX6qK9HjvKHD1Rq+vCYjzTwDyIRUCmcYUwVykWwCHihqsz3xaNsi0/rSFZaA
J1NFzadZDAPQL6W7x3vkP4uXVT1516ZHBzYvdDUIHccfl0p5XbM0QgWA5UTR
Nn/5zuRd8aSxF1+fC4b3tqZFab4pAozwIwHwCC64gTLGhioVMbyJpX1AhR5w
O3QbVoEL6ikxXlhvVXyUKnaI9UNw7dq8SnuoQX4pKmDYekSDjn0bH3XqgSAV
xbSgijoD0d5gySLpVqA4Dm+hNcIepEwXZQHJ1HLJlEfTa3fjwoNCx9WCUQ/t
ZCwmuKenZ/flNnwOtOxy9YgWJW7/Ft2yCIubDgAWGd/JV9apjpwibWlHkSDC
aRl5mvrM4eTjPOfYKYHzP8emz5regSfGMlknHlHCk6PDBmZdDZaUsGmn3EaK
y4J2IG3xdkL6+BlhSvSqIfKypgEliwoxWeoffMffkCVk/R1mgEjNq1FEOOLk
QtJuMnp7QHc0NRDuDFxssmZvbfTc/VEccxOgZ2BhRN7Dd5PFyjzVDZQuvOlf
1wpmr/4qyv00eI8cm9TJKLBOHbzOHh8hPpwhuwOgyjypmGSdwassUeDhpgaL
mG7Ay7oQA8+BmNAzjaKr/aPoql0OlhxRnklyrxdE3jlhmypgQJ9JZbd5pB2R
3n6tN7t2j4rQh0SedqA29wOVbIBZao2fpDyaon0nRWVf3vcWeGhBQSbGPLYO
8pjpIOnU45riGuQUi92BGRBYhd/9fByBgob/e0pAJ0IeiGNQfD1xxjUqg8M6
Y+HkBXVI+c/Vd0D+vifMNhHBrBPWTYVYker+l87DydaKSVvH9yMxmbxQDosa
5B1ASdsfVQ7zJ9B5v/oxiNeN7owHob0PjIlWFbmL2oG33549bIAeT48SZYg8
gGJovz59wyLumOBzwg8XDMkNas+7w+RhBAJjh1VECajeSecciF+3EdtQYYfC
q7hftA52XbbjjsUoqdtZ4LG7jRrQmt4WEWRI49beh2FEJuoR7bvCfqi7aZpX
t9ftaMKUpe5CNMnsZnCfltcbJ2XCIcv2+uM/gi13F5YdWwnGp5kB1bKCgDNw
G9VQiKnp7sOttxWiCtt5TIruQcCV/M33bdAyuChXPGi+fgm5+tkia2wxoz8q
s1yRiefYIVWbt6fEgjGukKL3oyzCDYETyHaFo7xYHdHLu/rPO6qRaxKmlUDz
lEH46f+S6qEUTKnDhci3gCGQcbbr9jR4tfpcy9hK95qYQ9wH4UVCjckrfMoV
ZsAseN4y3Y7Vbtf6o3091iv4CxrXQ002EEbiJrRLukaNBQ/Ei01wCL0KQ4c9
3GntfnslOkATYlOoA123OhlrvSFcTeZn4mxDQb8DxLj8kQ9BRJXKhnpY6309
7KUcGmrwwUYpedn5jFdB/oFknrodokYC1ctqgBAu3sqnhZZQDhYXYWpKtEce
yJZRNzdnHYMoMW45X5vL8KksYF4W7k48AXXydYcdrBtEGs0TcOzOusMOxfHg
XkJYekFqsAFbsLBbZ/4gyVqiqe89ataolG15s1Xobh4JfsxeQ2o/gYrR2TVG
3H6eah81gaZTVQczgblzcbFP7azJ5BDUMigwlJQnmGEF5vSLSCrULeEWVgTi
uqvSjmQHo59t9Nmzs0gnPvc1Gle9DrWqbw/3pJBjOgPdAoDwYEWQ0afytTo1
u4S0Fs5FC/Sja6oZHdA86/JGt1z48nx8/7GrS9huu4zM5NLklZUTiNzsLkOk
C+4TvQgAGprwM3LXXWos8QtKHUu2A5+PHzjztfg7xCx14ubofXURt78r/Dso
mQMoCDCoqVvk0Z+PMTEysfjkbxM+u6eeuR5h/mGMK1WjyVtURNqHLPq8kSNz
i8h5kiHUe2TSSuVPBndvqVOTTgNPDSVFAOvpc05ysQWay1rUPdkOWQ/O2dlu
PRCoIZLj5Wf3S0iMEaPy6GLi3UaBKhuNB51CxIR64mNes9ogipEfRtIu0awY
6KCA5iph8M6LZ/g9eUELnRG7KIVjo6X6aDNKrkmKgIqhgNTykjkH8GU5RDtO
3ejE+fAJkvFh3TigSSx1MgFLoFtdhtliTB0rVDWLbk0IwX14ztMDsualaZuN
FVs0u92Ekz/Odc6ZwtGwFq8S/LwpI+8raHv3jHQ040mks4kujaECNY1lgC9G
eCCMnBrw4lSHnpYyirDeTi3JsOGwU+6N2x7nLeP7vFNJxBQDzzdv/rho/0kq
CL2m737YJSpJHF1O5TalGWy5vchruuPSn/FitaIhmmtaiFr+tIySwU8FXGLc
NuWWidhJzmR/oOkVQmk2FAE2R2xymOZXoSk7iY2kG074EeAYiwr9fQbI4CwM
cnlR76HYY4jBJy54wy6o7mNiidwUFnvve39ebGndAIL3L7E5uykp8KxmbrnD
y8PC4P729M4wKdNluHK2efrBv4rGgHopVtBIYYTdKD7IxckN9sBhRVq2QKLR
cw3UkTgWIWTkxobilo0FWLHFxqD3PPl8v8AZ11bGWS1OdB9RAWRtbblFnlKb
qb/2LMp6ND+nPp3yKlt9DPDktg+Bi+6Sn44TVHF1yfvsiCUN9abxpoJEgf9u
ya1P+3RJ5YQVGtwhnS7c578oUmOlhEWOvvk3R39mQwEhf+v6Z7maQ7FGYnCq
D3BIeHqCCL91e/t/ua6WdsbBBxf5DOhqt1oN0tPhBI/ZW256QIIPwUVUmf4K
cfi9brxxwBRuHAiYZ5kcxriL17BPKGX91D0mvFyu/aPbWGse/GbWqaH26rHi
KHI13a9dqSjh5DEQq8soasLnzYLpxE58+3DZEFFGdXkMv7bvYHge3JpDgUev
Hts9Wm3xGH5JfbggHn0FOcCcg3XhwNHjWpFs/k9sLjKNDm4n7rZqohCNWdOG
++YxmJeJ0+DkoVf/FwIfLk7I0p33PKlC3+qRWYvaerJmBOLKO3ybfwjHyyYo
+OEn9CPjDf3foTv8x+y83Q1hxkUCg/AzQbV6JulNDrEBnma4qnkqRNdvj6CQ
uTZZmZZR8SWjBoTMzqgfdlpHMUk9pi+vy5XaFNkyUQ8wwwA2bvOBkk078u+1
6V9I4SqV+WQH7s0IkKau/OnVUFW79YGHrfxhrx6ABwrK8qqYs+PnEknug+iK
e913x5hDLMBUGMqAFQoaPWaxZodXXA+CuY+UTBBxFEqcuZHgMPypPf9CnOP9
FE68/2hBCvezii56u290CWZ+yRE0Qv911zJSpqGyzDv4Vo8yEZQAJiK4/o80
uiTqXRRNccitbnT0whGqSjdxMn+qXnEbya276f9efHttFo4Emh0fVp86j2Xw
PLD+DYAZFEchNtyyVvok8r5I5NEqE4zmnBx5m3oJRcV//J6xjT1th/PZ/i7L
ZvUS4QbericVTVXjjOtQPaQdoW9buFTxs9V1XYzSFX9SEprrH2VnG8EefdZ+
r5Z92yT6XDft6WVeTIvbujRUOrHA8I1UV+TTksMDHtCGYurpCADp6cTJ7gqu
Ra1kRJU5gbeCaKlNS6NOT6KyRBwAHjhQ5glizPlkslaDBWrKOO5gKTrNqLBR
FqKRF0FLISSeAocucpIKfChakMwPXBRxYnZitVhj5BF3frnPVkeLAZOYanAh
egJK4eRh3aDJvQV8JHzIyJXkO9UUiOQRvIUd9Bb/oFn9ZSV4GnG2HlFEBje8
3x33qnBI8k9sjeUOnHQPu76AbiEk0BwEywt68kjgba1u661JItSQuOJzNYeX
HH+JtjyGc3s5h1wT5sG/zICZz3UQnKC5MKvpwiizcKBaruwOacOoKZ2MNziM
ukkw6RpSHX+YoYKfGw4BS2oeHXn2P9wvZjevVoLoIBP/9lHwsyFtvMySG1EM
1O4Erly22y2aGUCzNXmNVUdFe1YuAMozDucY+k6yD4a2Nq+x9+/syslZDsgi
04AT3m+vFyZkcU+olXXD4PVlyVqM9egaOD1EfBeM6XRZFnX6f4UEldHbxtay
fZaf/fYOwDswFE+4j5hLvDvNH49XFeUxlN+Acqnf759XbPfbO7k4iLtJu0pq
FK40ZecU/LTqKIllBcs3dEJ8FUkrvLfcaSbb/7giCDd2oaDto/29gAO8n/ki
0S71KELi2HAgay9Q4LzhLKlaAHdZWctJ5x/eQKS6KuzXym7qYN8wlxH0wy1k
UXrzM6XwD0otcmku7hQloxkNJxVb7GCSev+g/RNXtHbjzzMVreuAMzfZ67rE
hu6414yXQSJI4XF3gRuodqom5e2W96qjsu27adosWmGAiTnHE1rf0haUyJXB
HPIWPqeXF9YT5m2K8OBF4jsYzbl2XAmQAijCm/Zucx3gGnm95AIXHSC6HfE3
5GVNI5TGpZlIhL8bBEyG8V9hJ40lQJGdbI9sMFJQWtmBpK/UCqMh0tJpzFJK
ALj9/XSoiUNRqb9747AeBal7F3rwRHsxT9zTml8O7VvZJQsW0iHw94ElTejI
kI1VCpUeHxwjfcBhtqYuLv391a1siMb2U8Xld8yYjhi1+QObXKysCAeXGSw9
9AQMfuH3Aj8xPHXdyX60g0EmcD2iL6yGLNAipLH/LojAK2lOfvLNolLEUl4L
p+UlFNlqrGSGHus+7QfksVut/jdRhe/0qLvvOW7zuj66kxAu2Yp0BTzhqe4P
hHQg1AmzanR2Ex1prTDVG6wtAgx2NhJJ5M7IsLQG7lgmjjDTq2SpPIANQv1S
RV+xcaWTCYidZmd0ZzgdvjmQgg7dNJG96O/9Sl9rzramuLAgjjXf2utuGvJ7
qkayN9CPgCBopDWBfVCALC8lpBrKC0tSpbEYCSLFd/LVvJDl9a01oubDGcu6
fdmEiJWnnFM/wUb3FOW37DFHs+reRV08WqKpV6kLawDgqM3wxF7Kwl4Nzmiw
SxNc15QQTMNabZX2I60vRzpZUw+Hoi2Vgby37j7z2eJdRK/l0tBXS8r55m9s
deXeY9r8yW5gZ5bWg5yAYBAx9HlpgTXRYi5NJXcAAPrzLLNblb+Imx3y5VRV
wVE+jkhfRdkVpoAyaMxSqg2Xfr4rbrJ/XZ+KanopGvDLgP5O2BhaU+mDgxI9
EK3e2fl06SK/qh+tw+M54ed6qnHM9YeHODfQgwyX4pIxXVv7Vxz3JrWdaeM3
DcoYqyMduCCfNdpaSPfRDYOmG4cThF9nn2VonRdKsYc5WIXdJlE1gjXniirL
FyfFbOEe/NJE1eyA1Br56ydwlwDjQe/3NL0YZonxPgQqctzgkto2Z88E3T3W
ovRqkfgQbT1zWTB1iF+GtGsGt35vZZkZcAfEeCvJMutefLu57wydFhS/Y3LN
x/gQ45/2k86QEqrTm681NQjt35tCzgsV03hHaIZK3zX684+Yd5KAjZcMed9J
h0sBRcaoMgq/aIKBN9+WPJey14MZcci8oAibv9TaVZFDTa5L8Fpl6gusnbK+
0SYznopzLJW0rMnTxvzk6Sd7giNYDeNjLBjkSJxUo7j9j19hFz5sH2wmD4OJ
ylInCS4jR/EpnZD9iEH1J0TPGINJADkrkByYyZIcOjieUSJTV+A63tQAOUz/
6OaE0mqvWXKkigkYesyVMQqJO2CTqNQfW91+swtve0hW5yx2yaDQ/h9GTwP3
gQ7nrLQoGThODIFWFoJzOs5oKNjJDW5jZuSUnAa1eWb7xGnWYhA5fwUUWf7N
e9aB8vKraI7o6HjKD5IT00OYzLSANt1U3vAizsPBMbu7tQ+EE8Z5rwYzz1UB
D5aQ0iS5WJOh1e3sswTfiiStNXh16biB4bhgkREMMtS4IFD79u0BrxBAabf+
yLqgAK2UVq9DB0q/7Moh5ElGu+3MIJeMhAe4SUki1gGM7bL+/FHnBAVJ8rlr
2xQvJ91aalFBnc18+DIfQaDDi0TaIrE+TbNiZiqvDHxnFaazbHB8QSbemLDO
tE7yTdyusrcDu2o5sg7E6aoq4E0Ve6mmt/CN4EV71iOVVAO1i50C0lA7oC3u
9FH1aK06zpL/n1o/ggSaHsTf2029DPo93PTpyCA0tdUwD8ferNguiSzXYSBR
hJZXa+qlT8hB70+k3GXbvj+5RnVF+Jp+biUNMjadG0VLYQ9F0O+9agG4NFFI
E/ObTlFQSzlh7E/ZsJ6B2Vccw1CXAz5DONuM8+3Icd7mhV03H7YNk1k6GVsP
nVWaZBFLluuwvAoodzdLcZApupLR28YuT5xuyHgg2PDSyCX/gpsldbFcY3d8
owUVX56JTlBOqxQhi97Lt9T6cPhxqQolPbfELNJ+IMzK4bfJCfTcO7rQ8sJW
TKzUQWg3tzO/8PaElx+YVfDFTtWLCe5XlvDDlbnrA6qMKD9bcRpXOoqKnSSU
m9747SZ77vXVynUomUYpLjYIdOLtshF8gULfjnVbzsyJ26Zd5bWaYsSR3u01
dfLSPQxZolil5P4eljcih2qouvmFKm+BYXTRVXiUeblUAOHvslvwBSRP15Bs
GqVWRcjA0pgM3/774vMaKS7R15sSgw7aTJj/g26HO3KUE0Cb526qe5rqPjyJ
BCG1j+z5V6yaXHynMSTxHHS4FptcKD5dUN1QvZ97kAJCHzAmKfqdJp5fqYMD
Lr9mFgrJ+jOzkodFR+uqMDmowsvL5XyKwJIe9sMTcDQuCs8pn1tRks2R9zQg
oNHJ/5NSoDiKUzucfAbysgcpeMOlVMvh9vjMLlFOkHLZtJVYT7JDQn1eSHNL
zAsPO+vwfO1JYPJ4tBOom25TB6A2ZzCEDlt4lIHszdvFajEmVe6acEQJ7USh
SGMEPyo79KMyIS7tKWnuuxtft2WNOBIuLHGJp/VhL1SOyO1MfZn/NAKIF0Mb
wKYh5quN5p0S1GyaDxvLQniHevvYG/1PhvUWy2VOawAA9ZCtDLrH1qqJHzyl
qpMmtdnXR+PAPtQCO7qDGHIZ3CAordCr8NbUFrmzmGo+9FZ3JKKiAu5Tbozn
rjgFDgr2gOMG3GU9TCaj/4hhyfOgpRIr/cULc/1nISCP/x1iN7qbWaV5fjZF
MxxY3dcq8fAxG+XgM/fcNTlx0Rduluy2D4Xnjw4n35rsfYrg3sqHoZWRHwkK
tRvl7soNDsGx6a7s8QXgc0Hz3RrktPvQOi4uMZckmp6nUtrgjLmyCkVOJHOb
ZgULD4QDWHUY/q8SBNaMT5raX9l0TwByh3lYV8C77cZitPzmvFQ+tUHMhNop
CwiytAU9STOn1yy3t1sw67IcJ4piewOxLqFVUjCnsG01UQVGhvClAGq3ZyiC
4a8pMVudt/DoZ9ggCjLbt1NIQ6sKH8Gek4zYQAUUG2K/wRJ9nIOoAi7HM7r1
Cr67IZslI88wxGmLzJ9r+SQk9EATpIVoyppKKC3lZ4dXcelGn21Qc1032uDj
dOpKG5nDT+gJQdhnDAbS7n7xvxfSRnp7GMfNUHKG+qIR347ywwV7GOIdEvl9
N7f5U5oZ238My7eZPntKUAnW7P/dgf0W3KRfkhBu/3U0w7UbBeZtM+hw7GTt
SwWYjUPuDHVW1KBk4P3xOwJsZjQpfBX2aii7IIqB20dn2CjP8/pX2vzCLbgK
4lI5KW+7CMXMj28rb+9Slp0jYzMPnfq9SadoEYno4OQsrG9/HcDMo3T6wDsw
aXXUa4M7Pe8zr5LWqIPyHwufE2svJpwsg3qrwGCVlzx/N7mM+1crdaQE1Q4T
3RQSfdUievafL1H34u1wpV1vzqsLjkcck58s7fcnVezid3lPgpLQ/wwbLXKl
FDI6rfds+IaP/MpP9Ol25t4xnWsGBH6jxsaFx9TxFQoc3QXLjlYh8ckSnOsC
YQhYQN+nCpG5nT/jQdPhZqg5fx73EdbUAAb7MGET5p9u3qPZkEEyr+3Q/7fY
23/wodFlAne7UL6uByW8OLZVG3QR6fmejd5p2bFZ0uHnVK3dPGTue9eLhspr
cBljeitmAhxV3s2Q8QVTPannFLMCWW6MGENLxiNO3uQHuMe2ShIgaQTPZmBv
KbeoUzXsESzLUokzYMRAzcSJcm57BrC0HqZJzhyNY3rnT+BIbnigcq3dFnaQ
B92U3sBE54zH8ihK/ATCaFXfUL1GYNKoqWX2mV4c8ZwmzZL6guOHl1k9eLcF
i5/4J+tW8l9Cq5ZQq0wyZn8oAORx3zqlFKgcnuw0MKHR7MDUJUe5m6/iHWV6
pfPFrE9LojdYoBm/+N0MEsuUAZEIHd+zqcwoh/LR0X8vTebbY0Lgx1Ttz6ow
UgkR8wwX64EBCyD+PhW+abQhTbCigM1JK+kWFpSbmwIYnghvrwTghJfzhcjs
F1ZABI5/79ryfpoiKYHQrIW+ZpFLvO2561xdfbMGtuc9+05ftuz+xSTunnkQ
Zf0VBVlkX9TJpOYrjVX9Ziii5nx/C7gp+Z/0IGQ9OkJDcMKpvdyP0IPo5QLA
X1xo7GwNYVojiGTv4w7wj/UEZ6VypVbA9tfK15OhCqpnNsphsw8tQ+L5VtNm
/xZnZBKKXTyzVvqpJKlyqSbrnmMxwB+vfmuXExufBc3f+c/p2UiASdm15bMd
cfcxBx0obOzWlzzjh6/4IGhU41YSXrU9tH5rULs6UUf921LcB/WcySS1LySz
WxszQV0g8kYIVa/QOXKE7ZMM1acLQpjCYRfpSnUT3jrEbolLnwDO3+8eJfVp
hmDgTJBE6AzzEL4toVDBCvS0PM6ahzLbAFHLdRpGAm0c/SDCfn2yudUEz6/H
nuOygYzrzkOwo5up69z7nWE5ULpV8VmNuG0Otmw4bV/ZLGAPz6+qe14GfHb4
+SLDyDn9j3HJw32oRynaLCNP5oiBW3gINvjUcqGMuGeC2SkMeLO7MJqUCJfi
noa2X1NaWupCDLHl3Q5nlLMPu6TahGCCJGaYXyZ65Fpu7sHDDkT81DICMXnK
GN2CmM1Qv2tPFHzkYE7h7rNfXOxZen6V+ikNBp2ho1mPFz31yaIb8NO9NoqT
k3sSe76UHJxzVRfB1/dQPUcBjcPSCXjQf+ZlMd3b2gzDX9Tp9QbFmZqVw64X
AHZ3WfGxkXYK0yYVWGACWnTRTSO2TIqivCEZiPUlgl7+34Y8Q5VFjZhdJpz+
kJ/e3NjOTzzm4ZfzxkmXJzh/U2KsEKJFJbyQRVvL4jGonKmFBT9CTrCCFexZ
G8c8QaymHfwDqzvFTWEAz3Z0V9tjVIN70ss8Hpps4urXqx5+W0o0kryKJmW+
WovZtnAVuY0qrjyMjUQjfAUURvpig9Ok/ijzVoROlxB4DEiyF9uKIokFGkFQ
dqDubCY0mYWx9iy7ey3E21mO3jeLj7xe22QpNIhYe8SSOYLBH6ZfSbA72P1P
no7fFmsQHXtQ36Ph/po9LCRmB+rsd6lf1YimwQMoYp2CMPlMeC7fr1XscDdW
639wPyFy3bZTxEpPCqepENZa22rGM+aRYoG/PaIdqErngVftjcCTC16rtOCW
aogzlQkB1+pY1bhflSZw937eWxgiC8jtlNvaHwyS6S1Q/+7a3ho3GPpoWwSw
yY5md1vjG8QTOfW21HEdeJM/i6gtMeR8kKWz0SZnZWhJDgW8CBR63PXuLb9z
pUkbWJkLtS6GKjFGBe2e20edB+8ugMSVta+gU1kpES4iFAuI+ms5iKdSylyo
iQdU/AQIAI32FfXEgx18iIBrfEG5UIB+wxtNwtpLN0YABQmRYcORsiH5reV5
omYmG07OY46ZbBc4Hk/xIHuPL++fh02bc1XaLsugtzj/E3/W/6Ww9iBwWOud
C0rlc4+3EipLA7s4b2a48yeWV1htcn2ufqTVe3iqM0NMME3Voq8VDOwG07jT
hDZmcj4R/dw8yaq/bNL119fzE6xMt27g5Ahor4cbuBy40fPoIriD5e4mDJKl
r2fA3AoDdvXi+Gdm6DMaBkFlBqugGHpxyirW6BeBI9a09AZQeihH9nLj+4w9
XbsGbbEMwzHl8f7QmHxHzXSFX1QshCQSHJgGGEK+D4pNa233hL5G6bAv8F7b
0ne6ahzeJbUxXLSbBRZdlPQOwWs7lZgmMgecQJKaojBG6PKPoDpjT6jYICqL
JJtkjXXPJQdbDrEeQLV8hmJt+2mmnnK4Xk09idAApSMLmRjfgaK2Mg/1JDlb
vI3Bsp5lggWQko3xN85rHUP+2Tzyanee48yA43ZSCyqBYfyXSHcrHvumtrmp
rCqep5JHZyuN+XSYldEC5QcJrExLMnDgOeHE71t4VhIFWuGp3Ij/gDPRwJ1M
sEZXIJcQkgDBxcXeJS7kaHYSLWF/vbvhtpkSFxOb0ezgh9tZyNVbpd/AamrI
uzaTIO/ay4po6bgW5aa0UnwutF90x+EqaVkmzmdTl7I6NHB6NrWvTE+GNaE0
WXrd1hn7rbkyspXTM+tWAVyxtXJ3B6tRdMRg5qplYLx/hlQgQFWpm6zTsnk5
OVSs2mNYoD5JXEfT9vY+BmCoPaBzxzJcDlpXZwPVM62AxZCflWVdNZWdgxxx
7msY08HoORlPRaaEnsBHgUEgh9yPJm8NcZYT05SFAbQTidMvlw7ypqVlYetR
7Tphvy/Ve6yff9Zq8BI3nqtUlE80IPIQh9bcZPE1HvhYU5/I2ZaprHdnpFqB
at4EImU0tZoqlbDWwQS0RxNqXBud2FQ7JMe1iFRKPbIN3vKjps+AZ7v+lE+B
DYsKwyrwKnJR0DO75GPY0vGJOVZkx0GwPEGXhQNfJtLULFSXfwHfkvoJI5UG
gekbVkuQ4H8eTtk0BkYJPw+bah/4ZM55bqQe0NliN6zPOCW4Jydvkj2IbIAg
zSO0hedIust2ZigtWIyGClThj5KeF+L24JXdhQVNRPwP2SUngt7kytT06PQd
uh707YRc6n3J7/DQWC0ys9omCJw9QVxCSijmEO3wNgp0q5T1E0vRNyZAbKAc
YN7fjnp4vBfc+qdncShanzkLMiCRBJy+wpmDnDJWtFczSYxEg2nHm1VXLzpR
HiGNODt3hGV+R4scCS8IDcBKr07jY6SIzfq6Ao8GHI+5qlZFxSXCgKf191pt
EmGBvPpRcc37owpmUghrbXorD9smFCxO67felQqEnTMVSPAqxASKKOhvgvyu
B/MndFRndbus8AxrpdIBJcK4/Dlc1F8+vqWao91gHBLgXt7Spz3xqZIBli+I
i2FBPQGSwHXVjXis4VTfNeJHZBxCI8AwkcykakvWWNVkRwYsl9ov1Q8kGsqi
qs4GKNPHlqNgb2nYVbb850M6jtdVP0l2Hr1NPUPZT8KhqLLltysYOE7U0PP2
y1I6tM9eoeT/3/2/uJhSgN5t5PiFkwKyJXBlWNjjoCD/n5QeCjrPGKwYDoQ4
RKbYKSqE6Jg2Of6sI0bM6f+BBUiGUERX03Y06n/L0INM+GcU5xZRvP9X7hdP
1TUihSgdlWgHRhCQZ637RsEbl+QwNyLBdzHk4PutwPnSHqnlKHqzlu2emz/K
rjgtuHuZxwHRTgHceHAXuYjO6pmQhABs5CO3gLnrZGgsM48a9h3OhfhyDoaP
Ns8FxN82jMlxqPhheXE69Kk7YtnP+RYYZ8vpSyTUPJDu1PNesSZn3MZwizVw
7MIn2jHLbjklv4CTi7Yl51y6nRO/a5eLbdH9YsirOXpeAV49xZv/i2J9bH93
K6kV984Jg0zgwDOHvWh1OFw8csNf9LyNtBZrkLXrB96K/O/cJ8HWNJ2Ks/ng
hrTG7ZysHh0LIoWuKY9UFe/OhHP2Qzo5KI1QTm/L7oryNN2egfD56Qvq6ck0
w44O6Aab63GoNE1UbfaEiD/YZOkL8TuQiGL/3oJ9keBmmmSQzNgjYeAS8xSg
4LdVHucJGNSO5xham+Bv+7s7buPjbagrES8to9sDT4FVHbUwD27j8LCM3Piq
CiZLoeelDJ0xJL5pfTgEDrDf718V7sr777v9HKrNx6llIezRGFENezLyHQIf
gFF/TaWuNn2u12Zuvk0sTHy9bW6aodjUzEL2zcbi2t3DIsNs1UXf9P5s9Yyj
2kzeKSUuW5bSKLznqKVwci6BIExycXqxXuRxzK7mclTqkNuXtHAiw0pF1UxW
nlnEt3LBn2Mt6WtzNPYVw3BSeLrp3ZJZoqoZk8QxSlATNwcH+7mkUfcinzs5
+b17ytRhUM3epFbgjUaXg3q59kg2+8HRy348wie4+QPW1jHs09OJ35Bm+EfU
We3Odw0nhn2hEnViWvxq+P5f2ixef7JyCmroFWYyQ5Dbug1AtsM+mjsU2jl5
Bb+Cu53tIpmL5eKh8OHRqVLYEOpBRUsVONdYeI2cRvZGDwu95+d5bSJ+0282
a8rNthPOe5KiuMxji1mnAmlz4NPQmK/X6r4NH7018J+r6cE1PJA4sdsmySX5
GV0gUCQMphgAJ5RANAbyS19DXXaaXlCFCKaBtx2l8zwZpcjAdaHQOXbUbU97
kWBtKW/CsNDzXHxuXuf1Q+uCZSWG8+PYgNq6mT0T2ybyOupaNF0ii1A1Dle2
fkRPwflGTOb88xYWDShfHYqhmWS6uQj+zmnrdy2DkWL8qXZhZjdCP5oJF2c5
p2M1s9KC0bENod8XJJ20NYqGhetFLg5wT68DGwe62SgT7fcDfqoTNIUjuTuG
GEfktoAmlCiXMtIy2W/zu0kebFTElDZoR0sThkOlTtOmjbkCZM4rKFcnyIwx
HxGM+CG0DKUo4jSBrwqxnjfGUNFcfpJrBCkmYk/1sOkRzUnEwbuuSg06LN8N
KZYtVFVxWgqZbXrC5fzw1F1IoU6QX9m+Ekj2L3mbl8XEuYZ06NOl491PoXv4
D1cGAuASZhMn3avmNvvNiILNZ64eFfH4yVdGONv0B6sczK77qdZeJsuQc0pi
RsJUMvU+WK0om4kIhXoJZ6AIHylr3CEbxrTJ7TsmqU9s4sJrhvJ/Yjb5OtUI
wiuS8Se+rxd0uiBOPxZFIoYjCtUSDnMZAFwZWkbMlOb9Ylovsy5sILZZBKRQ
Hssr7KnLoJUjqDLGQ8sX6q3DGOgE1fU0GBmG2XnzqoomlQ9TXeIXkF4+E9hM
VVkswFicMtSOnJD4gxYCiMIGtntGu89HtpwWyTPag2KFerSO5qwwvCYNPZt+
rFCawj1LOVencQG51g2aRoAXXVDgyTKEZ+d96dJIolHxXIUYhVbaId8B1I68
6NuOdECUDjarkpRJhzoqU9JH5VJbg8LxWSNnYHMLo73wSfSPqt0bdEwHo3W4
4x6cLPyk6fvv/fIS4WZc0UBb6XmiU+dCkAQrD/LjvWQ8E8L15SAmRt5Bijs7
sYHGMaabDj1gzEnGvaMvAqhl/WJpOWPPuUw58ysQCfd7jGx0RAtCVHMCbo64
tDWdzx6jLH7aXc77gDSzn7hNxjq2MrR6T1QL7OO5qoWDSLdtyi894wILa8mF
uhhMErQy0Ux3wyP6G33x0EuiFtMGYa99fQzTl3KZooCsVAyCuVRrzH/WLUZf
Lj3sqykAg3fcDzHIHV9B2y6VurUYff65uAx/1hSKBcZGr0/z+uvrX3TivN0r
1qGqr8E0Hvzc0tSVgXqHb3vzqenAFtTnjWGDrarh0DXR6nvSTA3BptVxLRj/
++lboAgLrfpe0aLmUaTSf7PjDCNGzsmse6PFT0Zs2oTIuSu9LdZVAtiwL6MS
GCv5R89fFkAcFrtoGDFQVyHvFMSbfiAoNGMUCoh+M3jvpv1g0NndFlTeGF4J
Ns/k/pWk/us+wezO0aeH6qgw3qTT7Hp1hEYHOMhtUpD+ufaLS88wDmL2JGsT
fMJ4//+CpUa/naItEuJlsrh7wXh2IBFKCCoIpcFbSCmss7/8bxmPPs3n1q9y
G55UF0QJLSs8Wq5W9SzZ0jcA0+pu5S++GZ2XMemgDLyNNSEXtY/tThmsIWug
JsdjRTEVSVjjJY3Zk5X4rIAvkUes4Bwr5REAwt3OD3G2aSzXOe4Qk3gVJrgS
Hrc3xqsGULxZD/pUnJzTykCnRt1XIuavA7S8gRdlvv2pNGn/oCQQAq5koN2P
scrGYt61apRZhPEYZQFfNxC5m3HR4Yc2D6edIG2mAycCXFhK9G11jPLOo8I6
9wCv8psmurbkgLQoISzZX8b5GdALkQt1o7pCcaIAIKp3XUzD92qf6DSS5jB1
dfU/Z1xynxlOiTMhjUGswVf/qbqL7fRNxCsEQDqVV0LYXlQLXGO4vpBjApoa
SLAP6hiYmOt/FWB9BzNk4eHNEPJZsCSu3ZPXNeD4gjRn5UmXdVWtB+GahNxv
vpoFYvLn/pARbCWVGti7KEWUgOX4yuH9DwTxGkoEeN5WTcG+H5GGeRokR0Bc
73QyIEC4rwzyUDSQZVkIJ8O0WfsLjQFK29in85pG98xLjScJL8ZyVCHKvJ/y
MGMDBPXsQGfK6PPJFiBwuiXvR0kNaRVqUc2TFDP+2YCYBqckpYSD27OZUuaf
oPTtUtRtlJTxv4fSU96C7fFOpQVcsa9vgg62BpVi7WaCMq1IazziZLqEzIo4
+XiLBlww4ybFAntAqtpSB/oXazPBJdEtb5vfADYBoWr8sQRLxFttq6mM/Hk4
BI1Zk3+GmdS3eO1jUhSIhHOBelRimQoeaU9th4LJbnqxjnATtnyhTjr4YJIG
Hbf+d5kxXLpBLc4sU6yap4cFWFRe2hqBicxgkTkJabYdjvkWkbBxJ5AzlOMt
Z2XP70Q+ztiJleqcdfhiSP2l9cXAGFwpmP9W1Lj3qfr7haecD/ZThx5PVtS5
sr5nxKpXBw8A4y0YvjTNKgY/yMO2g6Rr/CzoMLrGvv0tW8+/z27HWeplf0GF
zjs8A/VbGpKeJOyaTa4lXWP4y64GhyO0UUGGrFWMQBFRkvFACN6eHQxANlyt
AW3dBRmhL+uoVZBu29w1nVQO+jYBRMBHKjh5ZL5TATUL/hytRk0ogjAKbHwY
yoZzNT1DX1Y6ZJueIru7+rzyZWzpy1tUNG0jeGWQi9gmbxkWN5DBqSnkCKyJ
NevWnE5AYTq9toQEnKCBFHHrRh9W/amGglV2SJEroJq+BOUB2mKpe2peHsRN
W3ovTLcXyileWsyBSu1rQoPMtYJr7EJlyUlcLYUyUPMZ9PDR29Zh+d3IcN5Q
I7zZhqTQUU05tUsqO4S9j+c52OjxKoHY2kA0Vfk6MtWiMXJ2wV71KucJyGI9
RyMJUA6S2+if0uXtSaB0c14smhi2RzxVFaXVE7/k3sImNGWVDmC9zWxOTsF3
iRjmSwYuyxUFz08jQNfOuqeD5YbNpaLRQXc6pJKVJkw6xik4TXiPf6l6cRfJ
V1+02YN2kibQxwkYAU7EN0JNlhioSRivZWfEqSMqiP/YBnjAWwTmQy2zS22l
ohTfIjgBpy2MgD4Vf7n4IeQlg2VVDpoItPD4zZ6iBI8l23H0Kbv07yd8oOws
tLAac9AYqwgSsscmrlN4Rx0A0EZpLNKIQZGBNriv4pXPVTetBtYl92qcMPIA
FQ0XLUdonQvil9jbzeJTkSwrQMfZcvL47ty6j9uRR36MyeOH152OxF1hxaBs
PCfDGswDtIkmABvq/RH/7K1k29bvBMRXpNCmHL1CrJcJ9FOXXyi/xkf/I3mQ
4rJ3urVbz34hWZOMb4xTfZFShSuNR3SwmECGCEYNJfSppJcikjgKQoEbNCec
Us4N7IO6Jjb7pB/XY/vTTdpZyah1kuMZvWLHKUNfFnhGahZo+/KuGdoNAxmo
2EhAWtCjHnhMtY+vzcyUcmOAKaHmKIDClbByM8QY+izFBSFmrBTp5F57Ac5s
0OmKhG80UfCPdGpWo6yTICQWP1/kHPdYDhFeMiY1HIYomiySYuOKdfIC0Zlx
SRPMVbziLGt1cDHgDHmee9uXm+uKVVaDgODqulm4EAY1yHw3duWrE80EQ7vA
rU7nXaOpmn9Tm1/NX50sbAiCbyVweHyYNAeItp3ykkRXr9y+RAAuHwYeb44z
wFsD0EO4wgEr1HyIcwClI3Ac23VFk1SOoMrraAhSZwPmgZdjAHa/Yv7EWsZ8
/QtsUxfCrmuGmryN7QehKh/U5mYk+wN5zFAUaIMhTi8rLPrJBoIVfYnlaPe8
i8mqdMf9Y0LwNqXVM2bYBBO2Ti5j6yWc3f6kfYScBAN2Q0PWOXXRtkaBHIfp
Q/pUvZQdVKrf05TIP8ExLby3rbbsSNpaHHIbmOUrXUN+hMSVsuV7d1XJnx2W
07ABNqsw9Qzio6xM9LHgUMsM8o6bGN08fjLc/S8JyizohbWATh5VJYaVR2yY
7mke83NCDrElHwIEJXVnDpoCdU4FPLKwZZQmU3Q/kEPNcKmVPz3YkaRJxexe
hWNZcog2ckNZ6aRK9gLBdyo1+v2Uui7UpgjYtCQuzzzdWCCuHcElm599vlZg
Gi9NQWjm/nYlxy2k8z7dE27cwu/ug/5/cpkslKgwIIFa3S5taxLth9M2wfgu
DKfbmD78vroHjfqPHWLs5sqzM5gjEysMAhsYggv8J2O4LWkDZ02bmdwbhRtM
qNB/TnJ6QoZtlWI2AGUhRmWBDr8U3/qUkP/S+fkjHg++ktCNKkvZSKBSjHD6
LOMg2FX4P+1UrMICU5KwR813DQKJqsjIwK/Kzz5nV86xup1QhF2aSzLKL2qf
ktsoofj4yn95p9chf5AU7XxjSwuPLokF/x8QHK9gMMYIynTN8m5hPD/Th83o
tMlfdrTRZWQFIbC/+try4SZ9jOA/w5BVneIqPARtHpDwUZk5WhPGoj7Wd/VW
I7Iok34f/oQKQmdDPffRvlgiOfltbDkJMX+Fses3xbQOt4I0ZsKGY4sTUIlv
MsVsL1UxS8ePbr+VkF3YoAbuSf3jZQ/EyKpGLEZ3eG9h48FXY2DUlfkZfcD4
FDHK3Ime8b2u0mSXwNFMdLGKaPGH8QLbW8cOHgsOOca6fJSSLYB3QWNpboww
j8giYNf5Dquh1RAPyYTo/u74zmM9dp+H4ak+s7Pzs2tRamYYznjlicvQ4hNZ
VZjlsgNIXF3FJygURR9MYjsehN64OYaRXFjdR8SLdwIm82A14y2Wme0CE9oV
Veef5MPDkszFLNdUYwyRL3vTVeA/rWsgIebMNdPrDxRKjU7DlGaO5l3iyTh8
Rpr34Vf4hFRlAv8hzU7ZDtFZ4Ntl1q7qc2Q9hL860m/JWvIGjlUpg299yukF
z40er6z1VjSYcwD63jlpTyLIDkovLgzp8XNXii28Y+nvlVSbBUzsUjhnzd79
vMjBY5JFIRl/Pc0oZPVBXBNnCGTly/Lp6zIy4QMFMMJCkvM+3lg5aCK04gCl
G/hvrn1snf1a+OFmXvs28SJOptV2+ZN7EQme3hR3juVFmFG1QczPsuz9TOQb
VfW3bKNiruqd9N7EsXoiepEgfdAJhh+iUKM8IyVEYSuWXb6jItN/sU0oT2CX
8+uUFGt5NfFHsF26G8OH6Lf4vVtRjWMhTHKueITnyimaWDGmLUA6pJjwpw0n
EcSba4dc5A+OOwNupd+DRjbOLN4ftgwt/UJ0kQ2Vx0+MnPHrv+EDHwya1Mh7
nTxnDfAhsenhXdHBCz6VJZywo5HgVyQXqYPH3aPHZEOHTTiqlib7aDMDhEZt
x7qjnVnkrg29Zf47O1GsamVzoIEfBpm90PcDk3YQMfCs/yRPefdu6VeUOuhV
ZQrnqmHfMQaM3zhprkgdeIX+BhW629xk4FVcZU21Ka6keBcKSLQ7DFOw1ih4
x/pqKgVWjwtif8QsCHbfDPHKQPwbcT5vOXo8edbLCPo2sqs3hdwGikaJZ9c8
leYW9JYy1pFE2k5rnkjcBAFK3iNezrdA1ktm3/355aENUMcGUhNk1aupkVrb
5VUuisPZ+Ka26BsKymmXaypnTllciopsSItSDZ6xanqsJGbWKBfArmzew2t1
Fii8GvLALBN2gv5JpuoxBna/B2v5efmCPf8lfmble7HLh4OP78pxm4ktJ5VJ
n0iB9nDWQ//p+gblbBi6XnPxYouTrBfdj3wqGktNmRQnr2y4NKmfnUzqF+V/
fkPMvryBtLVAjvUVWZsVk45Y9D5uA9GyCGACsFfIe0Vhxv3NM0X+pbDI9d1W
RJzuSm4jmfkeR5p+f3vtJe5l9R3zmKsC64ZxUGamuuZ86avfl9eN6OuXpIDA
xQlweWRbbmkZiXJDDjesAy4aORRaDD1a/Crz82SjW40hReI25Ms3a2y+dE5R
TfPivB60//8RQboI00zv1MwpiBtWpSjXnF+PjBDavN7p0GZbQBJHCLavVNY1
P0Wo/FSgpIyRcQaXcX67QC+nQMAfYFm9GQ20EbPdXWucVjx31kcyHVOziZ9H
zdmDxdn2wbiP9NAS4Ktsao3p8S4ZWyf6B9SZtgkFTUA1+2vrcuSQmko1DqMc
YuvV4C7mtQcCA/z73J5GnPLdFGsI9P5Drl1wbwPBJsY5bYgOqu1xu+jAX/fO
T568X2To0X9uO+I5FEzwts8OkXWERN7TreCkgPgPkPTLm5kFGnXofGzYRuaX
GYYU2ZDoNNABdyacoyhXho5zYmu6a14ILn+shBGhWKMjoq1H++f9U4hXtfSj
7hAV2pGzpTnMvwzSKPHo0/HA17jnnbS8Yxcf0qhv4rNb0gE88AFVTaq0RtIO
w4ZvHSB8lz3nCyyPv5i2Co/3F5Mr66jHkum8Vm8PMuIY1V6zY5DB/XDhPXtW
TA09Etxh/S+rauc9K9Y7YNU3f38YOi5xCmImSjaTHUlcgIRCKq1A6Tcqbrof
JR2RWN3bqFJFGuQjeSHxT/xAkPHmZ9wcTq2pIdbdzliYgNOW/VHZIqhxooWW
yuTkmCfy54L6L5dl5hBj0pe3XvQKMgspZEz7EHjhGn7xT1JINKjZqIeg261F
GKUyhMVJ5mvSmgd9aD0UwfnJcAboaSJCAVXEcXNihIGxzfgcmegYzyaThI4n
HlJkoy2iror/NqDTYsI+plzpy4y0IRxqE0tQLvAwuvFRwI7JdFbgxfInlr8l
j1Zj3Pt3BWFrmdWpYFtnWa5Z1adNKFgC0045sZACin3fF/f4u0N9tjl/diSS
VgBzklqzMjI5x66XqY6LWZ9J8Xso04H6Uf+gtmNLYsHMYFePT77pKEABf5cH
byMjgidHminD7Gabw7jQ4AyzIXyv9wh3AH3PMdPvxmWVL0JQWL/uTuBw3q9j
92NtGJJ0ptx3hPDOFz/tH3K/Z+wu3oR/lSb8OTnlKjj2HChzAZqmCyKt7oBq
RVBB2uwYX9YjIZEp3coGkuzZB/Xx0e82BdmNjC+SHDsqf9ZsCl6ASsWh0akm
S6+KczufmfN80QM4DVxMBkidAcs/A6Ft+rCqCVgZhVbOIbTSrYvURbMGvfv2
hdq68jh3X3CCOSj2C0vMW85av4DUS05xWF9mzx1yFGBlP77sBWbAIHuhtgA3
mtb8LS6qYNP5Y11LAyzrks6TrkknU3CYCYVidFZ7I0DqJ3VXTJ2fQWFM7FVn
CmuvwNyQRbPCb1rH7benlVga9NYFNWJEAVTVNWow2Ngl0RRgUOEgoUzh/D50
Wl3R3GdmhOzXgIb+XMmxq9Di3Q+qUDdyd+gkxhQJs44zpDoRC+dm2JXulA3F
dWzoQQbDBYgz66th3OunPIqWOLeiOI3BzSGdlZn/mO4vVyHgDibfnUlzuwUZ
68v1dp555m9MCSwF7QP3TOq18TNoAk9vuHed9UfU5/7SzLVUrDFRT8UTDOZ9
kEAhxEMg8whlNeoE+Pp8kBeHbKn1rD2xjUwUOxvvDysQr7cPlZ4L7rrT6zCI
+2Am7xwIdevzYr8Eck01j+WTfFvuxwYJUrLOVIZYuyaMO/yUl2TVUMd0emQd
FJxM18qURFbNjWVXZzzANdAbSzc/ev/1jx2JyvYqv5ptdTJJ0sPnYC/SBpyQ
SupSoPrU6muLsVczARuRcHJb0CQj7N6Y1XpSjNJYJJinu4F7C7XRaJnb4lS6
Yf13KmrdpMDCiX66gMviTcor0aGpS9JSjkm9IIY1X8shFPIar7YpQ9NLOdpk
VFt0Qkh7K3ZM4WmIhPLL5ZsGgie0FnhjYfjAOTNmdN22fqh7Y5JqYigalR5M
gKRj0JWeVOmB7FW/tMC9JhebrHcIHMrwJcyunT4DbnwRbeNVNooXDtagJK1Z
B2TuBUwGURMxWdl12SUt2+9Izrk6kX130fORseGT+PyxEG6ZVFY+B1A+sPnu
uG7ccUo/SWDY56BXv+CPlh77CygejfM1XIy5lPAB/F9cxaxyhIuMU00MqfpV
3rKF59oDNMWAeR7bORCz7B9Flkxa04ZbCZMrvlg0aMlrVEd+XFMTnEo6tRkN
U/e+cUpsgH47H63IDpABKiuJQhF2d0iRdRFRqGvNzQVksPAtoTJzgt9w2l1H
6/RmjuF1XSqyEnjTEZlGhkoTEbNFXOnKP9Cx/XD5ykYiVEQpz3YdrkQgbshQ
rlY9jFGDEUNnx8vJHctscDu827FAd/IQJT946L+v3biZOUFt6Cm+6emHsyXJ
6lMbSPN8bQ4/fXb+a4M9LoBGdow3td9YZLHxdy2sK4iwqGfRi0v8HrWMxtU6
9MiUwysTXrDVfj+IAF76YSr7PK/V68cLUSe0peV8KOK5avUw7uOG5V2dBs8m
kzkg4plv/eVHI0BlL2sAz/1FwGhKHEpjJ/e20BMrH+MtwOa/Bkm4Z2jF4vly
X4QFAowrzlO41ZLb3v76qHG4LP2PEbw1BeMsYP9W1nbz3YWdXmi/Hm7jdc+j
FeBG+A55OQGaq24SLObwEtN9GVp2vKAAQpn8yCVmurK0xIAln42sXMy5DOd8
fJB8o6urkAkPpSSt/D6ulnz1vgYo5wGZ6uP0y+DqYQWhczob26TJNjcIwjez
6lhkUGxjxljU1hBl51aO46tHc6ZtNjvABSfUzglY9JpCiVqkcm56oleiWWY6
d9aqqA/UHzQT5im6u1CG2hxpSFntQj16TsgR9NUlchWMY7RsvnaER4mJtIdx
yuPVUvHCuh4CDbyw4qlfv1H7wOcaxzffXaJTkRZTSlxDLllFH3xo3Uvl2Me1
lbhuX2oNXOyrZzqrAP/IrhDaK0Rm9JD5vW5Wd9cTkeoACUEM8cS9qsf6pFvp
dCy4HN5UIh0bVjdXTTqNUldMJvIO08SAsGgxsl6N4l+OlYJMrE1vLF4qo2JX
ECiznPSGHHnHkdeElAC+lotBN2hGomKe/KVFmn733PteBV5oQVmFjg/QK0pH
dni6Vw8mxwqbu0OM0YQv319D2aqHleY3s5tzzx9FhHsyyEtf3KpZLcI/eAZ+
EVDxIPP32jrzMB3ScbpI42e936PK6OhS7rNkMgm+ShqQ24IF5TSMjWg8ymuG
kYsVVKx2yNFhnGhPwtWWVx79JcICBHajJbIf1zQ6GFuVKw5BVOh8BTJ6Fy3g
le7jcx+5SJofdKbzd6xUCO+2AjRATwQBWxM983yQuoGQURMRB1w3milSQy/r
WAh6glnjBvW0VVFtdormwbAWX2W4IEE1KGJFCwSsTRlNe6Mnb8ReCd8si7JO
aiXx3NV+VvW6LWXl4XjwORivlm+wKIwua+p4X4+vUJKc1m8ibOc8i5Kox343
sYXkopiNVZkMsXtaBI1u+6q0vRWsXgrDfNN6jZHdsNSEZ8aS1g4LujlJX6QR
PFlEmCBoomXvCHmsslTauACY1i8oEoIVqbguNuI3EfSDW9b8wXq3dH+YwnCh
65RG2OnAOv2s3gMhW4761b5Uw27q9ByuOWNGTd+3BfT/YCPYdGxopFvvuadO
LLw5qcPFgMV5QD6D2nPvC2Lmngr2LlPF0EeRBXeoWRLYrWi0nLQ2Y118f8CI
jz3U2cKERfYwtEwSFfO4SWyz6D8pcw3WXQFbnTPiLKt2cXsOToQg1DyC7sve
0gH5AlP/bxiNT/IG5NpcUf05A130folz3Iav7sPY56ILGh0DT9aOtVEFQtg1
FKLGn0msAfw/T2idP6hh7fNeTBrz0RHnji8kSjl6NNh02XdvJJE8T1Xs0ove
HUd8T6D+STuVNLkCplVtOAXBsFQGKQyt9+FoMapm8/J5zCVTfg94eKxjxUFR
fpH/Jr0UEFoTDwtBzThvxQg/1gvwDW/pMNm4Y6uDOJzLyMNn8faP/OY9W9mb
Vhy6EG6n46j2ccSG3BpzyBV6p0kTEh7rIg3P4UlRk0IUexn22+YrK5cwb9XN
UJpGeuDduV+yL7zGdNIwNp8NBriru1AhDHt6qX5M1+8rq9XcFAk95r3a5O32
BSwxs0yuGYBwTXHwB1tfEtnZ6K6SZvGJkOodJqIb0y2Scf+HKfU3FkCEMcLC
SNfeKhYT4CBIVGV+saz9JylwclbGnkkXDnqKb2Fg8oZ3gwxWjJutebTdK/D7
mBGXrj/i60H4Any2CLHBYCqoeVDMbDWqj8HfXZ8Drh2iJsxWb+p7lAxDnaJA
xBPhbr4p1XVmQzoUqyKG/HFo6rL9ZUoJNkRHWKGNziIKkmpBMxINfc3bUGCJ
aa/bJ8UHHyub2Z7uvs1gNzddHDrzwNAWoeZta9q+VskMvxKDsdnQ/aDWr1dt
zE3VIkLxxKTqR36hUITLLk1N8WJkLhUQvLRw2qa60LvMTjit17trkMOV9Ovr
DNcpd6JYXG2D4ajBElx3Ph47mTgboG/uNJyE6g6QhhaGrrH5zA2Tx7T8T9dE
56AjKCA6H02gbGp1EN+tLbcdyq7d4rL0Q4ssdtAeeqpSDQ3I/VDH+5nlqJ1V
jUO33476Odgy/FC8IQj3sv23W/kli9NqXDK2vgHWqiUJhv6/+Syj1o6w05D5
2pZD5CFgqrzx7+VzStEmo0xy4YrxLRtRBeoiHB7u77A6lcLfjQP/jZDSh+Y/
1Xy+Ivg7kGeWChPHkdEF2l/n1SS/e7kbhmo5HTnvZFARN040f4i49tAZIOW8
5NXEL2SmaBx4b4KfoOzYSr+YUm2MGIAs2wsoUBPXg8X5nZJQOzpCDfJ4Y/qt
wf8YlBL2BDr+011k3iktKyl1f/tF1PvgJXl6soPNAZAHH21VnB0lpooK4CWa
aJ4JBOtAAyZI8QRU60mkXYQBKQimVWJpuhT9p+Wlm9BSdNRbJqbnu0IjTy4r
3sN+sB28srzNZKI6nlp94uDKhMpvrKvYbqrLgRynlHBONXpTWte001X2qZyJ
3veVY+PuV1xKjV/557DpJxoa/rozSdv+GxQmXGQcMAfRJBF22HUXOXzJa4YX
tpVTCD7dWilXz76jwunonfuY8MD1bbJC8UVAbg2IhOpmG7jI6X6d8qNnh0Ek
FjnmwtkMqs79cmcDaetjyLMRSMjj4EuOvrevSQvWX/z5AY4Ph3r2ptQvYCkA
GfOtzC0fWCd2LNBDKWyFwuamOiDhieJ6KQ505A0VHGKMjAcnejqjbv60QNRs
7ORnHNwwPIidK1ndZycKQv8u+I+hBt9yuhP7pMKT7QQqaJP4kUHCvqMsy27q
ItWHQ+7GPJqEzQslHmL2YAfzNlgYqJCrEUkIE4o8rJScD2kymZiw7ygFQpc0
pHQPaowvT0TjIjKeQ8vtjmc7yXVS4rS3bwwKBbi6Q3qt/YFS0c++qAXGm8Wn
tZuDEezVSppFVQ/EzkZGqgWA6rWcIF60pkn5Ipt+Wj3TlP+G5hhGhoM0mDfk
5oKDWG2yTUXOABTADWFe1iU7cSLxom4YIzz/7pReNlhAhTeTbQa1D06ixqsU
BPQQ/iWJ+oWGYHFucK9/cxa8PobRPLitULJcOMmV35xXkHC7k5og5mKe/DdW
0wxBN8b1JsI8I5N0FMXwpai6gnmYgTAYBHY5kU5YD2IoSW6hUYuzuUz09qTP
HHNx5H13cT8122sKz8+/VJ+n7/e+DQnJrrx3hitHtLskZwecUoZgXxhe65Hi
Y4AKo2pGV3+Ww1eyCj7gyp/uO4iChddrnDhwQtFdvQFgycUKnxuf/c6VXKbe
szx9CogMhK8t0Zwcq1H/eOq7QlF3hmcuBWQoX9WQdPaMDOG70L7Bd0tXdXb1
yobWyHreJHxCTkR4ViUgo134PLCzE3rTOp8CiY3slto9FUZTtN+OdS/bokw3
WkgzPRRwt2QQ16diclFzb9mT/O58/XlcbOJutyXMIu632OxKNZqEvLX0W1jk
NnXKIfIB7K0YYnfUvI8HhXFFykiCD9ScDYSHvJHkn9ldS/YYRyNsYEvzizCt
avwGeEJlVty8yVI3AJawpEuec/yupe7V4p2u0kheemURQOND/NbW+GDIMvVz
wyRqfxHclRg0Pz22Cp2zLeINhMbbvv3PdfP23xWHco5XlhHExkhAZvHyU+dP
tA7eVBprA6oEODkAr25H/Ngk9KquzNfcWZYdUFgcTH6PFB/cFjg7oeIeo/qe
DYNB+7YUTmBVL4kW3hoq1wGKCronMLpmam7Kc5pMTuUTo/n87FykT+wzqxM1
5/FGwhYSAxmPK/SF3u9jIQroK6MtRTa76DAxMC2w03275MbW2EP/oZwEg1mO
Be2Rk9Wnzlc2UEeDef5yMW4vz4+fYeFcVNIH3wzUnZYG+cMOKbrxnx1MYYgq
rYWOlXksLzg+s+5bC16HDPPA1iPZBcHwbDetwgBEchI4Tpp+xjT4W8PntNOq
Goebjnk5cV/59q+ujAT7DdyfPKLPtLQU3tjr/CjRcZSV9ZVimazzJFReUnFk
d7htMe/dajZqWs91pOonO80tFRgWkwA6SfvN+zGpAn4/bE41lAkfD85MQIBT
NszJ22tTLGYzc5UC+cNh7ydDW71PNQYaQls8067sSz93Ije76hND7fLVVcOo
KT3atTqpDRUobeH0sjCKq0YyRUSZN5jrztfoa9Xmqccj9eh2OEZOQzji2Lh8
cz3/jbJffsM3xbIxwkwbfrEJngKZJtExAmpsHg94+gopcTHkdUObb1YBhbPU
uXrZoFnunyaEdMpkStj4spjwxU5M9Md2UAH8HCtYlhk5hP33SgK4cOxaaa9g
mUqLc5fqar02KwmS150dXJo5pQvhikaIERDQrRjSfoObFusUKoeh3VVIzFuM
4Y1XNFGik3hgRSVo1ghXEVALJLUcqMKXT3FPVrKZij2dgFU7x6zCgbRR0e5r
e20CKreOsCat2z4rGw4lYr6dxeGl1V+sK9CqlZKXqySpl7hztjwJNGqhuF6J
DOK1jveYyF5R02XX8GfRIKeu8qLHNZR5l9QAXvDoncfdpxsCcHPByQ7K58jU
vjohcxR2PVyLVC5Fbg0XptNQkw8Tq7FN86qoukGAlMvEByDu/Bp/E0nXH6TC
sDxGqeybrNksvGb5wN9o9Lmcr77HWwT6c6eyI2T9Y5LseUpGKXj5xf6iKtyF
c3X0dKGt9XjjLqB3GP4e03P9rwO9wsfeUxzpWLRPz1rrMI2X573LL13hIDEA
rJbt+WsV+rTGOEZ+fe3Uwyfa2s4DyVvBko2TWAnVEc4DQHCVDUfvI2zO4KIg
Ycj4zG0wG5qYiuIHBLw2/YcCtxTZL3lukb6Vsy9CPicV9uMNHOejLTFyKM5I
3SL39bV5oGwLVNx/Uq9EntjVoGcRrL+8HcAUh0YuNP/M18US7U+CcbqCc9xL
fOBbXd/zs6i3Us3+m8WudqreFihegzi4aGs8CpqV+53GQAFCuqF2VYOC5Vm1
7x6H9JQqyan4y7v202Vhod2tt0Ef7NIAnNnweTYBIN2U1uAZLF/Rwmh92CKW
+Ugjg35u5m8BpaFDtOk0JJ4jMOfTswbWU9eQlI/2/xqrTxYdUFPQbfeslatg
5SGpIg68Ay+aJeUhHZmHU0gi4sptXYrYbKfjHaDl3JeMb9gd8mjXil3y3OXj
9zIMXfItQBVWFHW+Xcgc7J+wOZ2wslINGqP7KSEbzpjP1MaHc8YEhnJevlBA
7urrO0wgNAIPOSIVOGu5cNmRygW7vZcycA8XPn4KG8OVxNtjqbRHzx4NGHQr
DWWuOmtWo3zxz1Dw2q9PpHpeP06M8RImtwv9aRiRyIr1NOCCcpnty9LGiFeZ
KvPe4vNipHOigVLi4eQbJMUmL26reiG2BMU1Lq4n4bbfdubvWeAdr4GTS0DF
LNjulkQCS2IOdeqbLPMdWJFRARy1QCV/Xf1Q+k6MS60uHjLk3j4Y7WDxDtmx
YXYczDKWC8rBXzDL+KlzCNfHYXvONu04vdi2pqOvX37uVbQVlFbhAJqsEDdS
Cx6OpF5TDK927xr9vH0aqavmvX/6p7cwWhOewPtxDCUC3uOQmMh0ghVMBniQ
LhIJ2c2qjlnGRiK1EQPSJNzMO7cX58b1nsh2K7/+whMZ6kiMwCrt3I4RJMAK
W5OqVW3UTcsvnjMElq/q+GlIDvJhFIE4uYrTXwwHBpWEGaKdirzYJkr14yl8
zWGVrkbJHZZ5IvPrzTpkNnrHHMxMafoxVtaRmQoPYFURvIKc4c9lJobGpkH6
CIqbIGYMcyw1nq5FOFZz6CGKgdybif9/7h/WNUmLV/Fr4oRDQEnmhALxmjFO
euwXfbUt8rjT5HclKWfMTAI9bier0w1Zf1/h2aaOCW8uR5iysIAriis5PbDJ
bgGonySvEnuu+p8WMC6gpIXPvdX35L8vonqOCNADtCN7rJMOi8Yil1htPFrx
1tpK1Klg0UF+9Fer48QUMHbPcT2Pq6NvVrmrZ5udwQiqw61xqhUK7TJ0aEGi
XgwEaHYpR8ernI+l1I4cT4LYd8iT/LWXWRBaxeW+tFvpIquqDLoYSk8m7ixb
SjiogxsHABwoTTVL3fhU8oSIcC2OM+J97YSG7Hje70VJFJpcXtnsoQNJuo2m
t7/biRtHI+vudPKCrzALCWSC+n+W/IXHXOSPnp8mwpTMcW4n2I+gOOprg1J5
8py0zR6yw+8wD5PGYwm+1dJsjNkEXKUMvor8Lu+dY6Mxjo6flC+3LNjZ2yOX
QVNBh3qt+qWTXR71/JJKnBkkxoCWukJjRBztAhINGTw+ZkTbDjbi+lYJ8qXT
XQ1eJnQuXZyOou+TA7yc2Uw6j+MUizuMeRJ2s/7v1o1mwnStcmoySibmMNgs
sNK6LZzUqeEVrdc2MR8RXpU0dJsTY+/FOkSvulGloovZBNxRvIQ/Uf4NYDFI
ihjQjIWVPMhI2syCbo19lxqvvbMqcyVfqwxBX+L8dw4rT/P9C9FIWuR42Qso
gN3LK27QXM6ioUE/HIiXwaILVBrz6xqIVF4ifFioTFC949qq7Z36wzWoQR7/
CmU7BLnIHmoUTJEcaCbs0nK08Spi0z2pMn3um4s7ZgPHEigdPl2RdrZ4PWwt
0TBRPyLwG1a4xVLDj/OxvwfYS8vcurEJIgi//iTEQNEaxAvbMziOJj9LxmAo
cqb8ywSrbmhh2MxDuD29FeBzSVFJjYt8MbBD87mZ02gbIsCEnXdCcpqujmiX
9uMA3pLp7GwFQnirtArMq44Fzh0wtzY+vgLxwkV3YqcmtoQ97Sg+wLAw80+5
8qoKMkIQpDB3bSadiD0/KhnNBWMkn80lPgaa3+KnosiiLanrqWnbbC4/eWRF
96YmDnHzB2pRr36hqr/pNMSXvuX6Se3lKYelp9b7eFKC3pYt6LnNVM9w5xWQ
/E6HdbPdRTeQAncqdXAiTHlujVfGJ+vGnd1fouAcQv0zeXGyC+vA5uB6McJr
ll7LR6LzKxNu0BuG+pfk9vGF3XONvfB9r+9AduWJJO8WeFuJ03eglfVMgfZ/
r3CI/KvGpdvV21fHavRjmptCEILiG7OY0uyVbNTu5LqfLAUgcuZz+N0OxZXQ
OD5rA2VCFjOlPaQQktxE53C16LCJXapQ5STyQmcG8qzKoU3EB2XRpB6w2Avn
+gw/vup8JQbpI2JBw/dE1JrgEozv5NwJhnKKxaTQf/ahVJAFXHTo/nwOlxdY
YBKqZaO10+WkiW4PqasnWkmEhxQ9o3csRHxWFaV/Ne+0wuZmVvbnjGhBADeT
LiAVPc0BNhyS1gL0mGcTVNCcACre9MzkXlijh/9UmZAr17lS8kNXZQJlSwbb
t3HwHhk3i8U+IZTYhv5Ii/5Ij9PGxW0g/4O6Pbqpy0L3r6fjjc3U19bcEe9b
eGbaSjqXI81FQps7H83UX4hhl2PcvHik0hZTRFYUq6G+1JtkhNLIsWHnssq6
ZpAd0uSus/ndYYDj6wxVZfjrsl0rVln+vlMQPIb5EDAveXouGUlbaGe12OZg
1mTtkmkhL7t7/k2hxI4/iF9rKdM9FnfkwlcM1EGDFwsfs37jzDblOkvXviyf
WnjSycAR3Ogw8cRYytOgy8mDHF1WIT2jKEoDsO2rraJuFHmOuqt3qQ1nPq13
JCz+PjXgSv+SB3bQxdgBEfxspBUAqB5T4U4+xcLePSNFDv6TgfcOgG8bY2eh
BhWotvtE5n/obJbK5I4b7zkjPZyIvVSBvrjY7nyORgoHsikEuh25fb6QBTKH
kq7ogh5mvfW3X5EoroR2KvaMKdfYouwfDcYORcnjajiS2sDjic1tAZlUfCt9
vFLjwHo4I8vgbsaFNoFP0HoOluuJJhOUF/2Xr1zy2xFwz28Q3pVYDAJSQF1g
sLWo3ZefsjBcrkzytofATX0o/OitONB6emi5ZEHaSUrN7Q3Bl11uKyb8SKr+
g7pOMobD21lbfzNKVpL6yEzs5ji+lx/vnOIjsYR17w+QV+0awWzVvZEJZj5P
wlQ/cTJFgiHIeemprt8hzy/r490l9lZAUwIBvzcsYDDef/v9/4fGFKGVmB45
srjrqOgqC6Q/PngzFZ8BtkhOhBs65AcmmeQ5fWKiYlx6EUrp3E1r+jCFBViX
5y2vZ27YRnH3xdcAVZlFWV4wsrYJ+2ZQebZHu2zH9n3C0zDBheM77fOZ371N
qDR0AFv52tWPP9f+KcjL/sucePTy+2S6bJNiV4yF+zxf0PWpP4ifL32Zv5F8
ilwtDu+G5AfcJrk8EfYesFNNcyHtT6ggZFS98s6e8N0d05sV39lvDsGGIJAx
pxy4ERVuqWn5Xvdkv/7ID/EIflJjOR1Y5rjVQ8On3pTE13RsgxJ6ApBTG/Un
2EqN8I2f7j4eLBdsh/+FY5YtHWtJUzmAkhGlVgxQfyEhcRIMCQHKBXY7hvnn
WYrU+PMIl6qlwldwGjlBJq2jOq5/Jc7zE+iY/5YC4AQdutcyVzIWxdZ2UY0a
H2m1f4+E3CROju3STWtcfYPanVs9Jpmx+z+4gJTXC8LRN8pkDDWQasqjROWF
WS1KQF+qmJ9/o5OmS5JvbZsEmfqWpy4Wedj6DxcNwoKaf6QNWDigMztzVVla
wEnakM7sT8bZnl4NIc2isZHj7talJlL1dUpkPDrzZPxq3M4LOeYn2Ned06LT
rWNjYHsFErKs7DXAnzxOLq0hQvFy0US8x+c/g8aTxb6cCwsmQMxoHey2TAJK
rlcq0+4pUDQ1zQCAJhSaEK20B0IH3Wx16crzh0+qJbA8alAvie61o5JnROE3
NfKYcoFFfXCq7XtoS1rdIvyrg1s8O1IBCY6R1R3mEbuDcc4VdI5Iok1UW+4m
+s0aIytblbkuJz8CY0kUjOkasDiXxE/h6c1BZiV8hjFv39o/IFN9yG+Di0Y7
AHi/P54S2EwfLl5N4HH5NOz58VirhC3ocFcb66IMMDRSyuOWpl4Gm9TXcfd5
gSXV9twWLUzGorQoc6rJA3ysXeBGYgR2AQCn2BiiTjM28BU1ecO4pYMoTCvR
pm7EEAh4pkBjLPtTeJkauMn0/7rGET75ps8bhEcb9MNhIw7xrraSReRZ+6CF
Koj2dkPRWp1T5iGMDQm11TGkufKEt9likItGP/i7FJxrRNtyWtSakQNo9Db+
P2ek5NjjRu1tzLjLjk+GCjW/Y9fZ1p3RkdsQF/yZCA0R8U35F+GIWOa0Xn1E
6NJ09d/+UQmFMUmmdACVlq0NSmVgLriQauf4Iih2k5re2KkEnqHGs/zd+ZC1
YdS17UBaRekSddG4OJMeQAj/eIMAo5+XZw2K9h5aF+Aufb6stlwWymKdire2
wp4sEl61S2svkIBPOhF/25/afroqTjwmSfq/tdT3Z2Rj6d0hes2vqJvoCE2U
HGy4eQPJzoSndcgUd6rqEsxHj1ejjUqkvLoOKlVLBnJhUhbgZ4OTVuOr83Mp
AyvSQLYdttICIb8LeyUu+HfJrKVCZ4CU5LXdqNq+1PSUSrx7AWfDLssJYQbF
Mh72vMlsSl/qrmem0GA0EB4kMW+mYeMCIxP+gJaGWHs7Xb02KPROQktNUv7z
W3fJL/EsDJmUrUi59tpnsARFy6Kzi7NuQV9ofSuZHfkCfmdWKKTGVCjdhqMh
by1jW+vbX8jroroTn/bjeOAjjgR+JY5UWjju7qJ99q4Y/avnlWjteXzBlWNt
mxrNNPiNRA6efsSfsY4XAzRMd/b1n8aPQCSvzn5jJLR4JdJuKztRhNQtHA9T
8rXr+iKtgy3J6pAUdi3kD77n78QmWZ2IWD6ArHYjlmNLjbx50NdZcBq9NegT
/lFnCm2egy0q3eASgnfY9qhJHTf54KpTug2YyJo93+Gk9o+kgvg79zUrEpEs
/GKL6JWdDId4dQL6gWevivwuLkVP/f/Z+KpqqAYMR8PePff6qBn0rWDDwUsP
uUfaJGPwZV09hSi/+xWsyw0CpqkfMQzlVG1zAahlEX3/mO6YzK47d3P1uzWz
ZYQofB292YLu8wKRLUsBmOKEX0McSJK1PxrLXDKyq4NP871dLXnXknrTveDo
qK7P0F5ukl+SaUs0IpD8Z0LQzUhs9qMFzE2ivjEgtRg0q3JCG+46pBJzUgSB
H1/HyAxQiQVZYttbb1UDkbhO7rA8QrqQSyjvXZUIMkOdr88EZLkgbN+161Rs
1LMxHKvQS9cOkjSIuxNDd/TCo1ARoGA/H3Wjqt3+R7pfdYm6eeivOri9VFZS
TyiwAO2ra9RdbdoBpoJo9WhKPX3sEWOQsatOMOxTZhsNBh4C+M1gX/0hXMJ+
LHXz1NPE/fW3FDTtmuYA+uJkq9ukSdShX+Voq7ySu4q0gMeNrmlY5u8vjvQl
tK8FHrtwo2zYTuhyIk/quSyk3XzhC7UqGCpNO51buXFq1/RNZ7OLuxysnApf
GvA/NBsGHsqJnwFuC0IBM+J9ZVvaKPlTqsegRcIaSpUGHFontyNz45hmrXyE
al7Pml15DstYAjzGny9MdMQuqJ4/YTDm0gxD3SeFuoRmmXF9Ms0eZZDyasQk
SQi48fr5Ho7bgoYjepnMkpsUaZI6fnMf50cWgay7s4eiOhmOa1SfxxC7u2pl
vs1KjJYzWypBK58JqYekSHScnJHzSjxD4AvP7kdr0cgg6fM4kENfkBi5bP5E
FcCrpR2jKnuev9Q1QHQ77qr8RjEdxWHGXi93N8wJjH8fCr5l4XK2TnE8hi3d
asKz9Esxb6Xn+a+zuSRDLuXFHVD25OcqIdrm+7MzgalMUHrQiotFK7vVB7aD
t5y4CBclMKYqAqqMeB8zwCevxIMhesUKwwlawugMhJVMhEN9cIhsVyugxISq
i0f00bJ/dSBAKyB7IpmQK4fUljJ1FOcHYEqe6qQLL6ejd3fX7Ei0BzxZIrC7
zGwapJsAPK9F/09FcsSIWTfCFfNQW7otYar/4zsrQAiNYq+Mt9HwDTmitfDM
EbIhBi2jxunYyfuQNbbQc5Z8RCvwSh8jASnsQCmQ3ae7U4Pns6FuoRmGW+tu
jJDhg/LpWdBGZN/Y4+vCfGWn2gB3k684fXNW8GO2jsFtUp/urY3R+ILwO//Z
FsCZprOPAA/CnZ1nKrmsDMknifwtTZCfZO25/qBlCKICaW0lmgrSW/By/V3M
ZdUdRQMsK4AW6YAzu4cOb8H6qYeF4SYPviwtW08KNP2NCVpkdSHZMDyZYWWl
6gsW/T89H52GKvjhjidmThzuV0iubZuaGoyTBehgv5AOXZh/dRdOkBn25F6A
LYkd96578o9BecuhOZlS6TJtB+dJh0fdPV+UTvRbXVqxz+yOxuatCH6Gkq9T
y5FcQl5XbntohBHD4eTLxwIY/TeLmENBuWkemaggXqUsO0iLiWA+abhSDxg1
WZP67mBlXVkCmooqfF0ubji6KhrIEU9dOYxKRyVYFX5SGwQgTi31JK3rZihN
M0aZ7Ledgl3kSNNZEKKd6fdwPsNYHk+chptmqztGUyHwHh+WFqoxlozoodc1
sApG5esN6kO49azhuSB8AGM2yj4Dp6DmvAZRcdCpywfXaDvXC3kRUog6VSsq
6TBWvmhjndRPL++9ZgUbpFlBExRwHeAZ4wfdKRKCIkGc2/Ox7JdkBR07sqza
VYu58ZY+ZGhBc4aNlR9iN7AI2xDK0r5xflgGKsdiGnnPm2OwRaeMcf58+zFf
ArZMZ0vOH2zcChzFzjgWKjG9/sHSWwtgNZoWQeAeL78jbCxKp/DfZ54fJj1i
GSjVZGsKoDovbz06yhWDnHWD3QcBF7CL1PjwUKeYrOikNRkNCUjYn8j4NWBU
CEFoNCvkQpUwYw1mb5MOCT3f0q3kkw9egLV51ddQYnwYgW2qJ8CVTz9s42q1
KG3MlG/kpB4X3w0IFyCalWMm7bxoG1vcL9e6yQhal42kBImtuw1+XiH5cMDN
4gtRK5Ms4imcUVr5NvSupVgqGwGFkpbHINkngDkGtybL6Q/2U3uxUWI3pTeC
TWXRhs9wKAUX2YzQ3Ed8oaPsfTg1yc82GhdHkUngLbQMUDRkLRAtGs9NCp7z
mXLBPU+2BrlBYawkQjRS0CHm300OsgB6rAinLo9GR0siHDk0v+nQ1cm1l8L5
FFr7cVcAoiaWLmM07po0jz3dYIrvxDZzZME/XYNr8Qd83+oQYc9O6gNNrIKD
9ywznfL7HcVB9mA75duvSZuW7Bkat+LJcJ94knX3WYDqV9fl/Il6qLCfNUbq
CtnDZ+quVdO5ZquHKtOpYzhAs/4Sg59SPr2HUrmAvxWjHIB+Y6GLh8u9z7da
twi3U+EvgB1V58Jg05vB4+bLo3SljgZgPO562jCHCOL5OF8c6ruvynk3OwDt
brX6zJXGEBgizLBZwFgc/e1yy1i6oclWQGvVld6n5WQZP1lqm0WxuekZerew
7BFfPTPNZWfLWz51AWeG63ewY+sUQgxIxlfbULf75mpZ4vAAeMw2U1wCtXHw
/Xxra36UfhjivmkwlH7D7gn+nLzG+jqxOQ0T+bPzDXMXFmuC308cIVlHTInI
x8PUg1fXrQ6Exx3G5waTqNxsqar7kGXcrbqH8OSpMQbVi1mmZNVOseJzhZlx
/X4VkMMLtnsjYbeLEEIXR4VgUGJjIJcxvaIN71ZFkVbhQmEtWANRb1LmITDf
y91JCANSd2QH7a5+ysMZrbaHfjJC2URMCVgrq/YxSJopCOlKXs09Qh/Vbbnu
Y2/SIMbdxP4DJcO1lRzWH4zXHOtnATaWvpjZNlUzyHibTv61kAP/frOFibtD
2KcC0fxZGowJ3aP23nJ7IJKw+lqH2qUidJydo2YLr7qNU98W84RPTAB1iQBG
a7P7i/eMdsayHosm33GrYTEgp3wAmwuUcIVXpLeGIQcH7gmVw0BKDv6yHz6/
I8HOwBIRc+PKcgRWTC+iwZBQxslcvOqc9s6vE8xiu7JmWXthqKWrS280W/ZK
jAO21QL+DDVXTqS2maiFZHJQ7U0fVcjruYB3SjXjS820O5Ow5y+KKhaSc6B5
AVJ8PRjd0aKL2jw7g1WoUhdH3V+o7LjVc8AoTWJtiBI7rcjSlTxkkkC3dhFb
2FZvZt/LnCOfuoKIsI40dRXLsxMvBMqQ5GYL1BunVuZdbdNoAn97FU7eHv3k
Js8NhF+gJ8RJnnSKUhvtdo+vXmobkMWgjB+iJC4sbf3rqxMpNfGb4Zcz/fe6
CclKPlMNArjgb3uTd7ScNbqjtruM+zY783QjlBcA+XqtPsWRoDTdQ2ofPNHP
oCsRNy0VOg3hSuGRvXVU1x5+6F8wmxdTpWON0zuWn/CNrTTBc2QFhd+pSalC
0tQsGbqmRiB7UrIWosaoGSCF1ZrOYSuFWdwhA6CEfbQyXa6hBjbUFfR2Ffq9
DE/2IughHHH61C2AScyTKqepZnKZqjMFIKXEPRMZ6kVjfM9HMaXUb7lz7U4q
XllQpfB3EABix124imCgRvXEAFodSoEWw4YVPZzgmrqEVpOWnuxqFfFEaMI+
X+AZsjqMeR9tqN3JAK9uaqYRcacK6QVLn6XqT0aFvuoYDk7wZRIpecrWTf2a
KlYBcSwJTvOkTQSiKYS1V2yYVT+xC94IS+HlBMtRwOW/+mh1gHqDm9kufBVB
VZtYrgIjY6ejmSoyjXvikklrUIc6QU/C5zrmC7qzqxJX7MCJWboKwOoI+uhT
0LJXE9uLcR2F7vvbNtwnWkmM6E2duDbbCGa0jnccvW1Q7QSYKRBTsRetgEO2
UrLdLp67H6sBiHX2jaRBUt0MnwBmVSsS5lrjU9wUJifKEjERGh3l+HM8Ezg4
X8310kxcwBoIMmHzONZBcbg+P2PCovp+aCfn8OXIAyocQlv7Qr9l9hUYlqVz
qT4fUYfd7+Qo+pG2KZUPRwwdWmrk/JXcanrji7o/kRpPHLpJOmotH9eAixEO
uGGlgd4dGCAABF/jco+QPmTI2S2ZQZcoIe+EOnUGAiIJVZhWIkOEM3is8EZY
buAtygoU87AYVPQGs0juHind7YBN2jV6zYCr7pfIgirfWeq2sKGxBTB66jO1
3P22aP0SBAtQSv8k1Cu+lIKoFy7g15CjITHtTMPxF5+6CruHkQi9aleXGu9K
ge8UDYvamzLBtuaJbuFsRTMg0f/Y4YzfdkDMmbTpEyeZbtp+2x8YHAuXQz67
8ZlbiyfiziAD+Ndd6iyg1ZgG8guUcej16imAw2GjRujhNewPnatwTLdvAuF8
FtnJ2Rr/eMmg5jE5dTLNHZGkU3Khei0zBNXMArDNr2DkyzUgkqwRvqjc+mcp
tdcCb/gFRkAX5nlawhYiBwgpKaVTimoMQd/6YMes0YuVF+U4/IZ0uyq9C9Aj
MMcSoqJPrFD/w40qyb+KoSM5rUBe/yKV//ZZOD7Ribtk4srztNdND1tARful
IwaZBeCqf92towMJFYsc6JFH7yCeTJRWF1DXmXhOczP7S9E54WBzyBJONWqe
Gcs/SXmzsZ91jE1ahTHWzIDEROl+t9NgBdEDjd1w7ggdurUPmQGGmzAmQoJl
kgFoiqYjt53+DuLXmvQRbD/ujSfxIMVJS3vSkvEN82ELmwLFBcvuWTLzqH3a
M2rRXJKMpHkxvCqj+09zOeWloCPkPUYt36YoCSr6Qf8HcwHOWE9TqUYKSUBv
M2ZpGbzwF/YWy9koFmhfHB67D+3FbquHY6VXPJf5lXjwy7kyj7paVfpQfPsS
6xKdpcRwuR6ErEY2cm4i/ETzG19p3hk8l/BqHhajGFTQW914kgrLobfysMIL
okAoNa2mklEY+pOOucM/3EyDjm3ezMyfgbuOUK2VJDAlGa6CWOlkQh34CmzO
BigW5VjhI8Xv3uhTBxROp/zTVQX/GgK6tD8PGPFsw35sUlcBjNaDRNF1xRbZ
B9Mmm9zakY6lMLBBiOPXnGfLZVgYa0IXBehIcg1ceKm6JIORkJqJibkb3JcO
6gkGh7fz74431VwAgYAXtx7+MDTw3xGrqAZIFBQXK/EZntwmKUATgybg0U2s
t7hohiXBpgsY/OC9MoJjJdoZxS1J/2XCNeUIVBCoDByHXexK8jgFnVz8Eaa6
yiHgzYCMOIgscm1zumYFEGW7uYTU5aYM5baZgSaPVjF28ZGr01arrDzfX59g
BvkcMKpnvT570gfFa2wC7u9nsSj0vznSzvfGXc1RLrIidKabY6KP7nwh4+fp
bZJpkeNxiE2Cq4VGEHA9cIxJKTAgDzAv6L9pFvUadKo78r4qkwF5ZYq9OCBk
62HEO3N/WHXjj3syduM822r+vMEf8PLa+RmwsF9OrpjsIJSU8pZdze06ko2w
PrUOWjDrvjE5aLimQXMsHJE50APUczRWdY8nuZqBt/Ppt6AeixrrsywOAaJR
Y8cyA0XmzIjOf3iQAaDqOSTuChDUWw/xvZOOynjTy9JFUd5mOquPFYteEH9N
8whZj7Zt/YXepFjHxKJGsxawYxwfRJcWWQ/f49Y7GS5l8MnQqUx5CTmEeIDp
PYdgeGgHMpr3cFPk8x+V00Y9/A+iXw+TFhRpxTFfc93KZBJ9nDqDRhHwoAeN
3ukMAG+BAOLY9xFI82aEW2S+BMZyTS+Yk3PS2lGE/rlmjX3CzcdQIF7JAyHG
1l2OVhsJCTvCltGPs4Q++qdPNa05pTLU+XNmqJMuECwsDrlL5eCZmUKZAzz9
3iWpsLpOxgDN8mX5UW5eU1i8OKZBzzH+YWufU4cnZHSV6dyaSvCmgpQYg2rm
PA4OlOhIYL9aIDMxLBqZMxERUqGRVw0mHtZGFMXJ+dzZEdNE5h/9Wu7aF/uX
QKgxh5kNhtKTRBumPh2NGDo5tlwVpqInwSDRbgvx348Lgp1eJRHYIZgcEnd+
Vq1eVYtfmDLRNvYIfm96qchYpjj6giO7Dh2BTDvbGiPbAlHnLjK8F23HweNO
C8n5HaGXjU2swIiQ4LTsJnsvji+kcI2Q1iFxQIyC+ZSBn2PVLJwhI9wSV46F
7IegYtLnaihXLESBmsXWs3zBAujCBpxWZlRvPyf/hRrt4GDLDeb4Wlxr64yr
Xo9cN99+ggjV63eZEWXaJhBH+PPfBdm5qm0PDh4Y6S9DYQ5lxmGicQBDflqG
uL9lW13rWoG47SNX++ye27TNmJ9F7nVhQqYl87OCbSuTCAFQwS4pD+grTkLk
rlEZKqDtFjw8KWh1yrdx+mNuA2OiPQQVdyv6wuZJa0/nGSlFQlZ9EKUf5+Ov
TESs1bdGZ9Y91KxsKfbCPGd/YvAFZIxVQ1gK4iIL48PmSQJPhUTbEVsOzfE9
NTe5Mu0UywVIzlu3Rcahew50oHVGsCigMjUuK1UL26UvcWTx1vPod2VjIKPs
Niv5p5VsH/Ff3Uk5ua0P4OHorTdL9ldI6s0L8iwMD+pljq7VvY+SGeQwTP7u
iszygyagsWolZXJ2TocP41MOwXyhspr2N0C4Y2nvkDnP0QyXg1fE5JMi8nGO
u6kZbQiescZkVBF9m3IH2XJvJlJtPlANV5ClfVwT93R8nYFgkPwNqNF9WeZQ
z0dc2HoE/W0fJvbKBdieQLE+nKIZssYqikaZ4wzdHFIzc6frfyD1ELdeUbpH
9rE/4qjLRy88ew7iXgw3bA+mxLw+woy1JrBu8BSVy379z5h/IqDsAo9ZOCtO
2z1pfC5kXslgXFlp4EN/rUHzM0m3TytZNrpUjVEUDTmQh7tLUSAV6dMdH3cA
hULgbID2t1zctbo4fCerreyfGi3uN5aEEjwHUJ9OfRIOxvyeOrL8e6WLd7RN
DfC+4c05ftLHVvJw2g+sPzNOI2MwawpwD2s81bxtdvKbBtD5CzNVBOIvSyEW
q8WBcGFTKK1p8rPxNWmiCuA5z52i9VX3coY3UgKhx+1FRItQp+1ZszkkDn2W
CkzFTdNPlNtl7OtZYB+oE1SUcCaS/goLQ/tEZ+8mESBscaFZq0+8JHMgf8ri
ZzFBYQ9otWCM2AFe+7GlsRrWvto/qX6H9uSWo+NZXwH3VLQqHtuq1ssG6Iiv
DL8hSFhwujcxS9A+EdfCMQkdY85CqcbseooRVG7GvU9JGzD5GV9vBuUaOCPp
aTR+OFlESW1Q/kKLrHMh/KBa9SM3fWPWjobCj2iEf8s89DMpHNH0XclgOSYA
T9Ql4ODOHiRZN2XxzfW7DIKkGukxjWABd0/+Sp1+rqTeyvme/w0UTQY53v7E
5sENUWolo2wf0cxaHjE+hY+9Gl3rDG5loSeVfPQNMybtyHF4+Af3QpEWdcdZ
3OWuI+6pbDSRFqTMnTON75WcF2gLz+9YMUaYD7kf/76E9c9FsDcJN4uVTaO8
lwQGaDM6dX2ktQJNi9yWj6gkMJuwcmwAnaA2/5zF4Xr0PEtp3VikCaO79wit
3sbSGrbsqkeNL5a7haRS6fQ1a4CSBUXGPx9f1HZWBEdFpC4t0xpg9M4pgSWp
yDrDxPNpVya72A2zE1CqXtE6CDyimt89QAV+ru7IJUnbzIvgLpgdmqEJdTy+
879c5+BXnE3x7G9MROaUo1E0Af3F7jAUEFi6W0/aQtsBbzWDQAaxkYb7F7Rd
A6UZFbLIM0zUYsCuJjHIwylfQdpTzSoA58E+yOpD/P8uTka7UBsTDAEi5JFt
VIVtDZrU4fE0YQqgDmnB9dxAJzxcorhnP8FW0OwbQIj58B+Z2eKUDOwcIwLq
HQsa6ZrIIKTHCKm7dShJ1B4NVmGJfOVGfa9IFplP2Y69ez6+VGyC8oLnzbXd
A95P90skewbBZJ1y0gtsO36dZILCHBLOcFPTUmD9LS1o81UYcBcEhnUn7wmE
zB7AkNT4kkqZCJLixKMevgftdjEMKhCMvzHcRBEtjfVZu71F6aNsYv4L8YK/
ZUcCnaiV2+ml4FXiYeIi91Vk+i6Z+Ah4kcs+E/AZ9CYs7Y71D6TqSBS02aOp
7mcWY8+TTXLkPDQPojPyLhS4KS3tK/pxvxvG2s8y4PzmRaiKl1CmPKHAR1Gc
9BUb2t/HEsX+RRVCi0eH0do9nKEsFSKzyAJ448XICrPRHQWt0NujIfjKFGCY
WaB9N2ThiMQa85V6WLCSDy3AwiJkd++5OejyWU73l8wuSHiBA2vu7W1aBHGs
w25erdiop8Usb2sAo/2mTmBFgEiNIl4ZAVR4PnuQG6I81Gxy5CRkNah7iBTg
3Z8jFe69gi03OM45B+GgQvbfmzLqUDawMGeTQrGLvuDK6uosm2X7M9czXLXK
jCDXHBTboyl0fr//Z9pyh/Tmnyy7zQimlxnj/DzUTGLwXKg6LLKAuj9HCUke
oPN0y3YAT8ASoAR+/gJ21iyEdz655pU1NurricvaX8kb6aEUgEEgR1Nv0Y8s
ze9p8v7fv6tWUsOWsMxE5omimnkYAoMzw2TQ6BeV3xZ8PWv7goEPRVlJI4a8
Og8zv4PNv9lQgfpK0NJLU7eF0GvTmhjF4B80MEGLFWIy252lSSxx1VgH9uD/
0JIs697x2VMmt5747rIPMSofelnltgzzWMCbpvvelIvb9AKgc+Obwj09oQEw
o40boT9Emj35lCTFom/JHY63tAEWG7z7vBqODgRoG5dKsihVU/33vdckOPW9
sak7Qcp6W2WHVCMfAsIwy+HKPRH49nSgRiOeotuBGTRzWCh7G02Y+Ui9Au2S
4dtT2btRZLIIo63LMbRlOhPIhPXlUTolUB4xB1fj7yIuEgpOBVpNFrCbhfb6
zyb8PK5wgOLtSz85PGks+cWzvfXpPIbRa+vkCjKPLMKPuZackzViC3Z43XsB
dEyN77wsmzJ1ocjQa6r1wL5NBruwuYLoT3orzRAe2OxLrryaSNH6m6Dh29NY
1OPOLrCtJtSD3uj0MeQbp1bKH1/ZtA5B82BYWgr3gljP6V9i6BH2x00OYuLN
xnDZ/HRRX01FDjlrLmS6C7tAifJiNGxiN8i4D25F5oe9ea5c3Tic0mtXBaeY
cq/avy1hxLSTOdYR1EzpYBAq5DE9xAk6+iJ2dkRIEK1pxas65bGT+5z3TNSZ
HsIClK7oYkOqNGgtZqVBlpC4cweTDBpiTAbSg9TZIFr5cu+cDnHfTIE6wzP1
vaiBx1ls436HUT1zm6t/qqhdQjPxKrd8NOdrg4va08hjgdP/yH4LzCxU3OWP
0Z8kUEuoe8LoCVuizcbbDhHZMR321jgMN06vxbByjHsqafdW4QteJ3pIO+FH
lLS4zOiXigy9glRvZ2YeZa3OvSb57FZcum7ZWe4kf2ADmIFj7mTPkfUotRY1
kTaSQHADWvDR1kxCn9lLhCp3JsLordZrmEX4z8yJLQmk5cnF8mtXYtQTTgXo
HC441e4cGz3q3ZZRxSoFjS9kh3XqqZ6FHftMrmdzjABrlQxOR4XKCfTwE182
FDup5HUDBjFwJ2eNY4IQVVolbRNlJm31pWtaMOW0vQA/coRfNKdcD+LnSNEh
a/dor+1XOFW+8hNvPxw5mkFwqaBMe9YXShgOZYjBvF3LCaTtRntjET729kKm
+urDDbE7sg5wz3Gdom2TZBj3mmdB+rrUnGnk1mI8uzQSkNmNYgJFoHQWobCF
b5VI9qbfCk64tNmMj67Xo3lpeao8vYcFHobGy1tz64FBQTg8Ch/C+d9UK1df
rvQxQ/tii4B7McYPGlLPpDawbr8SRKMjlvrPnIeNQSJn8hOqrJN1IcXKmXzw
g18JyWU0ZtX0vLi6F3pPI9k4Esbf5b1BSz4w8Z0Ve+/sYCEJEPtv90LQ079B
38II5WZYhcHJY+2+SFcYr8l1muHBme5ZsH8gdjDv8ZRntgAWIL7DWaWcK66f
xfDD+z68HEh6krzoKYSvohsyWEWLf69UjIRcDwCsfIY7/IjEz76GcaIv5XMc
TZJBCjKbe0ui/GdXmGg2ta3UCitgztDbwlw5p5uLgSdPSfIKjXkqrM+0Mu13
Bv3GdF8mDOOr3zF/EnSW4qwmLvTYkcHqtkcVZXmWm5PdpK2Yt6mzoVzSC/M3
CALdW/Gu4bejdIOQ7iri5wbg6DSr0It1zNfe6N2iatVvHQBgQ7nIlLQk1Q0Q
dt4A66xgL3X84ZDYpMo97e/JOucduDcRcMF/cpH1nwBlaPuu1+oDbhZ6T/HE
cn4ZeUld+yz6omEG/dye+cqlPk2yMkh/N0NPsnIvJhmnRfBOlQ6Tg6QwFE1e
Bevu0+gh8x63kRhj0LlJzLxNbqMOyESlH8zxCdGkFXCo89LuNvZVt9lZOrSu
lmbAHItQ99ROxzrmCoafgDg4kFXX+QfwyXEXWfdBwWByOf/Yr0IZvtAL8R+c
4UXfAn5uaGE2gZDCMxZhApBhJ3ffZEqsGhuD4Vci45WSC7T9BCD4Rcdwwfpf
eNXyvAmsWuODjkkzegc3zpoG4nsu4LeFKU7HI1TzQ5Lo41WAAnYIpQnHNhNn
Bllx/9Bm73xoLNJrlmYlldPhemw4nx3aJWdo7/HuFNckLsDrBP/03eJPVhJb
5bEi4nV9khRCgK2nhSNDeyfgZ4TvKA4shrieRDlRiUWnmvVAO0kZioXDVDU0
ulY3Jctgf1rA6Y01bDicxKvHoTcrQj8lwxS398qmqRLqhX9WU4yTrqbVZyzg
uMxWxSyu3FBogY5WUYRGyg1e4/Lx0ML+9JTEorrYpNXellgusPALsXgneLyZ
Afbvdgl0XzPLNinYyA6469hM4AJ4bCPFNZH8X6J7+7ZrBySxFgvuDGm8vXQs
R0KdIQxkHoHcvPJwLASB7nYB+3zkSenm9tXhpxwc17WaHQUdFHwSLE0wisU1
td5g8KipB+maogF3ix0k6h8fCsfDdQp4FMrEuNkM6+mXO85qMzA32EQlBbFd
jHksgJC9CEq9Ysr4e8d64biNhAmp2+ZQKUlabUJfKygjBeSnLunBN8ofoglf
v3BA3DgBWeaiog1dxoBAyr/FLFBh3uRHppn9e85Z2FIHPZXYqQeiFa9eRjGt
oCtSApxRg9kgc2ie9FMerxGMEwDE8i4Zd+EnUqVw0bSYT7y1TjUfRR1HyVUM
hDXGswmcmYjOj9zAugNGm4y9VOg5GgnUFzg+0NpxilaCreEQwTkOgA7+FeHu
ZmYKnQHQm8IxNXdnd4aNaSBBwpKfKvcjGzajvxQhQPhqfEzKlcJv2YeL8ZLy
xF1x/4U5yOyJZR4oZ2G3sXmo2mAY/ZFOyk7Da1jyKftwe+x/ZTpRIxv4PsUZ
LMx9jRlXza03uiAJ9OAqMCgkA8tftgvpyriL3jZQy3O48NU9gHhTnSe2W1rj
2zjXZLDVQHJB5kLmv3wieAhkuMws+ELK/eFxaWXelPZniOfBQLEIt67CIqkI
UId+5VS21ezCFn/HdZImC0QwQ6eTp9qQaLRR7LSd0FZ1QUG8iNNN5D1e9sV0
o7Q4VnIHrutXpdBPOTAhMQsV/7+tjMRxKW4lg49ZhPxznA5h+nzx+30D5Am7
ySaA9u/qGBqOPxPK800gIL0MerLpMKaLCRQyQeOqr4TDOhAnG+4bIdTJFv1v
JFIJYezFGE6pJpw3vNYrhmjlbKI0Zkrfc7iM+DKwfgpYSYzj4UOrOkm97zWG
q/GHpVvFcrlrR9tQxthAgHAv/K6kDRcWpoqeonXqvHVZ84D4f+nCF5+rR32l
9y5tNzsGfprteaGz4XDiYmAx15D3VHLpPKKNP8xhwJ0b8Brz6i7+b5M0ok2V
zKgr4riUr1oP7KhuDe1JF80lMTr8BCPiPFr6UCr/Gxwozq5Kj+X97JoKPDh/
4oqHfD9tIOnUM0Mqw2TdjolYcmtaiOdxvL+ixT8cYCIJQtP6+/yF2jvVF8s5
+cBEncpJo470+ykoJvdl2RD8PIzmdJt36uN3SWyEYF0y3aDv0pccna+o900V
H8LZn9lvkIr6oEeZcw/5CDVE3Z763bMVdFB5QqTL4EGCop9em26yhhNmHb3+
C/lhJAIrM12Ki83Eqxki8cUepaRVk6CS8TPZC+RxlE7hp89fEzYuW1zfag7c
d7VLeO3AklPiE1kMyWjHlRn9Q2lGTTYfmAwJxH+tBIcCO4G2XHHFb75UN2KP
puImxo2E4XomzdC+aD6p7o/ztO0u/RBv/WuRR0xSPgbZ0TmHReKSqQkAWHEB
tMh1XD37uTwc6rujn/blO43v9PAYO6uTCLGFCrRzPO2eEQUZBa04SWZpSAzz
qKLzCqGaU9SD6rZaA7IhFhvSO5Fys0B1+w04ed2C8xH6ZqBUKOwVnccl9xZC
a3OiwGTo46YJhJODb0kVsGQuMfoNVwKqRrMQMv1J9jOPIRAJxbfDg9ggAjzg
brItgmNn8O1lybrYUbWVvEbI8nJnimo+zHQ64Q+PpXwd6DpmrQCgCzDnt78F
4mZ3yciOgd5Pp56yOGKtwI4jBY6IDLzfVuz2RawzYnVHgk2SvX9wyFKGTOwp
lS4QWZ5UJFdq8lc16T8m8KxZmIZz/Ye8VEkXRfvVa6TY8opoyCBcPO0tc8vi
OoZQSHZVTdErm3LVNnW/0saW4zquB40q6hnJlwNKf9V3co+b5dDpGOgWNsbI
yjoNtFqbM8YlefnL589sf4Jx6HlrE0av6HRDM4A9sF9vfJDSniNrJy0CrAon
/N8v+h4p/Ujw3Xf0mZyNbAb8LhEmctcr9syqRFcXxxfpzewzrLkaiQC03tv3
ofoj3UtWfWVgZxsrxWuSE3h4oYmIyPkc9UzKay/IHDBV1kShnONeuZcNW0oc
kznnXUCs/BG8vPw6UH31gLcfMY5y1Ce7eTUOyYeYpgOPdBRM/lsHDz2XzQlD
8LGkWw2IdF5gbx1BP1qi5BQZn3W2kVHL27zgoKzJBpAQEQCqjwJtrTGyOsUb
ipvymQQwQIxTYjWCuHnmbddViEyqzKX0+6NnMxh9Fc9NI+TfPjPaXIp52E4L
Hgyh0ZFBLXwnsLGHrM+iFxBtLma+0vNZTpciNjsEPDRPYAGgrtR/1oiMZnK2
ThokEX8O6hl5a+p9BvK+UjmJHezSyxNxkFgq9Qvnrs+ZvGYvwJS85lAZtnDc
ACYmY9pVr2KTJaF6h79H0MnUmB2bzBdYuWI57EBDEmsP2Jg1KuBtBR7JbGk9
wkDxLufgu24U6ncBKl28KpUASG0iFBqBfG2QPJhDAuH4V95w+ZxWAAmFvbV/
uYbjFcwCWcoj8HHBJ7KWI83kD+YYyo6IL4Hs2lJFG/ruHCIGUDssP8oNCkYX
5E29HKjE5OFoFIgV1yBmwQfO52Dmo6Ddz3J+CdtTrSXVdOfgDPSKPNJ8JDdY
cfzBqcY3beqyhJhpSXRAjhZe3Xq73bA8Zu7yIuCpeJwv/sqyU9n1mG6A+eff
FzbkJN9N5FNpolf/VodfYt9UwNf9jhtwpTCxyq7GB0jjhN1vMy157vIK7hlC
NJAF867eihXLEISyAUmNPP2l+T3DlOYAgjPYs1LGZe4xDYy7SEfTVGYhMTWQ
D7CKRgM81dkO1PUlzV4nA+yZ77QjONAojKv69UIOEy6hfDamFrzdHyHm2tE8
icLI47yWL6yGr3P/9N21GwYpOkurIN7RLnqwTdswRVySxlV7Un2y4mLLibTI
gzi5gWcgKTrJcFxmZn+l4u3ts2T4gOS75JvPn+HmPm8eaS5+PqbiMP4ssesi
8yXug+F3+h7dcrKcTF79KjfHIIZGRixYwBN66y7MEkte3OHhhjw1gzU+pG72
GFf9GVwy6JQGkTxH30MZ45DHn8Xq+k495m1hPaqNe8nO9QerxbxeSKJKhgrQ
zROkco31Wzli2x2rLOrWjHQyoDjMS2PjGDg10o9v9iNa91gp0tR/Kmf2V9Gx
z+MoqFoJ4TOtHiZB4ZiHNthDzvwPlzuPkljg0dZp2VfRRPdYRv27j/fes+oF
rtpea9KqzJP292FApa1Mks5EVZ6LHWataX7COCmTpknFJMeBFjDaVifST95f
BWEwDd5PODMAPlQEo9CFgcfGeNFz6u24pQ2WYlyDjXJDNDzbkjxZkDGgtE9q
4A7hDJcgi5AXWri/JUusaVlfNaS0RHaMi+2h4lyb6xvd+2NbZLtpyPWK/ArC
g7X6UC6YGvQFOm0jqk6Z2EiMr28Y3mKqX7GEvUeWiFQ4ME2kz8iqGxAqeAxl
8GqioU6S2NzEc/EAJfm+3n431k8hA4JbarUuk1DkXzzQWnMYNPih78jll5xU
AaD/f0lTGG41Q4K9xwOEOhbMVVS70IvWyP1e59Kolgj9SvZciYZQiJlIdyUo
BqY3Lvz06yEJDOG+ZXDmxQcmhL6t6kgACkPWkjXt8zGW1WKuWmvpOzh74FD1
17lPTrX4lnga406qmSZbPJYA6kx54i/0XaX2+OstSIIkv6XPH5pTW5uOvoUO
4oECse0Jb8nIWdhXeuGZtRtv4zqsL8yKnahf8mFNYhFzRcQ1R+HtXObx37iF
tU2b6GNWdj4DdcOCCWBjrEAl2di+XQpBpms+sAMtnjKhLTzp068avkz6RZQB
LbyxMIj1c6r641UC3Op3NjXvZm3eOlCVug+SSwtknI2IPSZLfaX9feFVOmhN
1L7W/7751MDHj4QZIHxEwmf9HzSvbC4rILP+lnNXEXa/BfCRiA2m2O5kJD2e
oRO8IxnRTSIb0LvbyaijWlM/845geKrW94e6kAx4Q2cIJiHT1Sru8JwZS/ei
GdB5k7tlw6OJtOjQl9hjmGv61jfY9NEa/ot23Qh5G9H3WR05HWXRUo9xdIts
0NxplfdGO6c3qGd4MMNyDXAycvQhdfZee3TVkx91A057Zv42xmrXny1lF8TA
pJvQEKcBkkrttORUUiynfeqMax0szZQwy+v4L8dH5DGX+Y6NtRr/WVBvkgnH
7/N76kqwuok2wewUA5R5MHl4H2xqsOqpUmH3Auqu5+t1wM2U1A/Uu6SidvrF
MLOQ1+erpbSMeN2Aewcs7uvxUu6sav5K7OQmDh+pjGoyg86qXmuuNmRyBnsw
CsWFlUI1seXVYwrP2Rxm19RDVXEwYB9A7f9e/UAoBSmLwW07jgjaofJzSdwJ
17VPmZM+te2zhyaHibAZF71qc0lL3Teku756rhwakF5+L/DHLjaNtmmuS7mn
PZYflm56qOk/UktN18taZN65GVQVAl18146wiHOql4pnGVSnMtFtPwpSy+ir
KL7WlOe3kbFR+uvccBZevfrPrCYy5K/0LqffM7kPDrcXLJMx+UYbn8w9AZ9M
GN+cCHBR/xPqPwQO6Jw+6JavSU51owxj7bVJN5Ir9r7Iy2WS9caUbpaVfOri
QPZ+QcqPpRs+83nxN2jUG1I3rdsAyY+sqMhkV0FWI+gstiVY+mWaGp7P1LP8
TWGN+70SSI4vcjB//UeeWpag8YH9k5yGb2eq0zYiQsgG+fNhb76Q3HpVrNPE
7+luSGAUaTkiN51CPlbtkbmhgcMIM5r08hAVYVoH7QTwk1+uRj+9zK6R3ba4
Gna/HbRpHH/jAy66uDfF98fEACmgwASpqxC94jbtL7m0NQa5Af+NYJ5ptcKf
z8pEIq4p8i+xnCjvY741yEx20lvMEvkrWtqKvRQ0RvAk9T09f6hfsmCccuzd
NGsjl6bzxT2HRXOGedm/YWo3rfAwgShAGEDngDh0OJ7FsOtAX5Ogfh4p2jqo
WxwfSVZJUVawkfrLbfu/yotI8ILVr9sUv9NzYfOa6zjEaN/fmFTAh7y2Cb9h
9BUcjwUNy1fRKClLO9ONOOpS8LB462D7G++HGElO1ZWutrLTbSdNIsUcTgjb
3spead2ereyXwITyPOyUdn/mFEtnANZc7wxgcW/Li81IOwPtWvb2Lwp+tTcD
hzZUfm0FtF84bDX8pdv2reyBhCy3zmRIGF59LAHgy76KDNMa/LcBWF/q3Ibt
a/Fna88RrzhQ42VJjGg3bn0Gnzd/bx0+nUSG8aQVq54o3jGTOm4Cv9cV8FcO
gbFxKLr8ALSjVoC6V29JVA6a+5fwXvomifCAnLm9ZBB89aBo46zit8J04PtJ
79rXlzr9bFvdoEcxBXX2Ug8iw0wX8KD6yXuTbN8kK1S2OO6BSNMSq+qlU/de
44ZzKbnGqolwwzdWCv5uZEn/9eB5gk7ykiuVkudk3EHytLknRGpvst7iyUVW
LBJMkVJWACIvt1P2kVTr+BLxqFU5FAJ8wpOSqvsoE+B+4Y5fln20PtBhuz66
9n8FihKx0GZ6OZspbjZTMCPO3PFsBRLTl1S8k9iGQHwP9Q4wu20vYBeF4qyZ
FoOlreHnUnFYchIIJjX99EtuuyFNmGZP9DpYL3cwix4/a1kwB4xM9V99Bos1
6ZYnpNiG1MiTrpxws+kgDKZ9nMbUHEAGKzTEB5N4Os37GXq95ZE2DiiaiyKf
VMXMbE3r21ZOJIThBot4AsG7jMzLzTjMLusJ0paZvSPmJHtvx0Qru+hAeL4i
VKNHR9srf2RUmH8+XSvyP/ebuIuExokPrye1nIMgRIZZBq4bw0KeL43MzvJ7
P8t2yE6mS66NIS15Ih955Fw7xQleDleby90xEgokfZCkNySec5pSwt4uKtgO
SiPM6bSmq9UlxOA0v1eqRErLurFaIaDL5OZdmNnjrvYOpCYjIe9MWfKaEDTT
z2T9UacxzQzVznNYyogG/Vu+z/TmTeJS2cOSV+DcHkilR9MLT9fi3P14vyQF
Biw0VqoURBI/+p3zz+057kzT0IAknZKzqgCNZJnTKunZMEvq5Xh4sJWPF737
hFekD89PYiDx+GwyrZ8OYo9STc9VYokAsmIJV9QX2C3OulnO8Tf+0FuohlNi
En8QIXy14Yo6oa49pkqROxvq1f0bgjrgs1/W7YlbwIlluVd7CmP+pf9/USQo
G9kQmczWQ328ENcH5kwB/F44CWZzYLFPJbzzadkGRFG7qI53dWCi8YnlRDvK
8D35RFwGmg8w87OUq+ZbWSmcsVJ8ygeTU1UCKXimsn9AwpMztMF+oLq//uwQ
/kbtaH1VM2cKg5hHODmH/EShIc9nsm0BtA2Wf7mDKuyjOdiOkQxMGXBnGolc
O4NadM4GMrKvBwo5MxI9wo8xd0wrgNLzCA15EAQmV0m3PdN6st/WnfICDlT4
ajWtHfGsRj1CqKLeY6rq5NQi/TCcYpJjLPNY7QbEa7YBpJ38tM4vntl8iDGT
4wHxyiG0BLYiwqWtwpWKul9pwHBvC3gtmmRuiGX4mYpyWbeuPtDhqJB0xhpH
MQC9s4y9BUuRvvo3NdRC+tKeTP/Skwh1SGPHnKEpajjmTz/y4kf0w8Qbouzy
xmkEst3l9/ATWRqFm7iX4ay9J7Wu6PAMZObdGoJWIRob/yh7LQv/37bhsBRT
d7tcVMHSEaSe4+E2k6agTqwlZLVZycuTdZd2zd5spqKvERx49CAhfA+Yxz5y
qjex2Mzn7OaV/FYfvhIoBtoq9niKrAiVMlTvMfcL4Iwmq7MlmxoWP9VJvPjz
2nlERPCLjvosbjB/n4FS4TmSvdQ/tJy0C2XJB7zJLy4FwI/mnG0eDQlzK1an
9pG0yza7CvNkPWWjlDIEuE6bCmi/kpHcjb3wrZCz1oveIYlR7vdR5S/XDsJ0
PurXzeMOjJjyua0ip4AxX4s+tAMY8pekr/lJLgNpocy/2noSb4uvuLOg55I9
8aD/psp5tQmgTWCTOP8glNT8sbuxP0xLAWFYl5ZQGZ3BXxUQLUNRuAaRm84h
TyWV3OlhaCm8DlmLG0bkA83PfxFHZtd4FbO56LGYQK6dDTZm2BaRmwtiKn0T
TBdV9L+sweBzzq2K//5svO4Pu0fuyEPrkcfWRPljcCGiX/mQ4lVa8IlkjrnK
kOTJeCm7oDk1YKV7tlcWco6r10/gNzes3KvByXEQ1kBM5zF/1Zt+7X08FEsj
XxGToiRlWhegtzQUBIJVWr7oOQn8wY2KH2ZsMuJym7tmE2pOCzLZ5A/VpCBQ
MzsT0l0NhNQCglRdJlvX9jYcCaIvYo253NB7N6zKnueSi00F8Ahs2dhjXswJ
8s1MUV8pN9Nsmm/irKrtTB0gddS+p2JDpq8PAYhihjopWBhgMqC+vNMeZCer
uWtmk/y65Xw9T5ZBYofYc+jJ2LoUvCs+SfasX40YK6jCggbXDYufVPQLaE3D
tuD0ufEMOsf9o4b6LpC1wN0/X/pxVTkkwq0j/DIvX/eHESiOTFdDlI7oI4tI
GrGZGDYffjpjZRiN3LAqGMMCOExDzqH8gW5kWVelQELg/OVE/4qC7pTZN+kz
ADAm8qdtKl4VILSAlS3gzkrONx7k7axo2KXi1Qmbmemru43wM7J7kOuiFxh5
TDccQsyR0NTLaZdfPzCbIroPg+Ur3oyez+oOSzsOB2RtBXhPA5LZ25nFvvOr
tuQN6S3Hd2Px4avtz3hFQqVFU7NdCnW0/PB819EAgRM6cNhqaBKcJMMwrVw6
F90GhVTyRbbzNPp2ommXXdi2pLybbSDGEEdfKGFGzfiWmvDNk5KWdTa/ojPl
B1yQGYzmFwnKM7Nb+jaF9n4i7ZBmEWMInvOtuqP5ZPLDvsoWp34/cMAyzz1A
z/0TxXgsJoB6rbeMOK0DEP+YPnKMKp1BJ4upHqi9ctObX0dAzHxDrAd19jVi
uk9pX7QdVz3A4bNsQQsYTnpNrqhB7mCD8D5a02L4fwkB6mNhdciBXHrlZxeQ
RVlQAPv4BeDztIaibJoIoW/l0ODN2a/9jIx9kithEENBYSnWhqpG6QIZ6m98
eRxMbFX0Hf4p9J+fG9xQF3njfyi2C8XMiF31/bDYKB+W7mIZcZOIQpKCZh1m
0ZoPoDvsUrWdkETMnKlHlnOAp065EUgzeDVX6F+VUMH9tldxJE6K5b/1n2S6
w/fQiOrxFQ1wNSolJixHRoVyrS0VoUMlg/FtnasF3NYzAt9l/gEGoH6Icq2T
zLsgEZ0h8XO7+cAsji7ImfFaBd/LKQdnp/ogJcscWGSMF/1dTs3OjdTc+Anq
moFis2bZK/dRGcioPeUBRlvzRpHnjOH5YXlmH++ZOB8wkd9wCIFhc9P9dpv0
Xdekb6F8mgtlQs0cvPfrI2MWnhP3ySPntcY8nEWccJtQIJsUo34C+R0LpKII
sHAAieRI4v5b6EmBMh1c6jLG80FPJ1skKhbJSHUcPbwQ9JtcdlSfT7c7n+Uv
YLDTQslhpjo3br8S9DxtMKHlZH38VGBc+WxFdbgywl7JoOaTnk8UcvrzSKHm
3bdukz8rA8d834HN6eyXQX6EJ338CuCn1I+ZLM2/3jbCU+zqk/q2Uk2FRseq
DYPdNb/vL39mU/raJJ3ETIy45DuSY6Cz98Yv2JVr7RToL52Riqe+pMRE0swB
zm3+uLSznB/jJN0FrAYvT+x0tRNauDmAPDu32SgklmpREm8s+WlahH9bhVWS
brRrtPIU2eBTCRmgl96P1MX5HyAQ3BTSKC4XtbX2wYDHfbJNE8zR04sDgIMX
JFNZ1OSqx0kFnSw7oTrEwrps30hU00apzIQinci2SXJcsocCUABNxKZb1mQr
h8C5xuJEPngpViF8FAVOe0kCRMrKcVnH6cpXrbHxRdWOiwpvdpDFE+2j31wW
8wERtpzslENsoKD99LgyJxOQ9y7usv/yyK5rBJyLnEGQIjDgk/Dbd0QlTqTU
DwXL5zF4L7kn24h4WCZclrLnq+Ldy/1rinLXwVs6rS5hSnPm0z/nL6LnT3An
wTEW/EVZUsR7wbFJtl6zPks//T4KQMnszvEgQj2BgyOatf+hcTUR8BRR9yKV
ZENsfnQgKWKiM1ldF3i8ky+tnT2OM2Va4dz3lBZvJ2uFKAiZ5DRCgOQjEk3i
Iibb5hUcvmTmBlrV9bKKy3/T5mFxfr/xiv1n/TdUCNSREeb0V+HHW+wcluGF
CUqsOWFTq1+qxEnHmGPoNhCyNVILtovhgEz24o2WkOXmkdVWmCpioT7KXrAI
ZS1CHJc6QLjaVod1PQksXgPRkEBC3WZCdwhW9SYmadcFY5DD0eoqRfshIyME
97rtW6w1Ay83Uh7LH+RCPD9xmypXNG9jlcxZoHo628y0lO4mHfAed0ygw8IM
lbDu51D+ZeH7f2ZVtfj97pOHOUnwICFYMPLY89As6XvXXdDb9tQ9ivROyUm+
8aBgyfb9B29TLGt+tcBS1MWdWtxnRMVv4741Q/5kzZujkw6//PFXKLCQr9yG
0LkcR+c/G1+8+yv4bCa9G/XTvKdjRiOykGkOA2e9FjuS+7w8Wjug/ML5DDui
Pv58Oa7iZYWTbXh+m1NpFnLBLaRX9hj0T5m1XPnmByRS5MEWCJwuReZMXpIY
79GGB6UiP+Tv7D4F8ngIsvNwB6uD7km6xofEah8k5a2UzvS+3hwJqp4gx8D+
e2XsyKxoFKc3RVVTxVH8ZsKSeDzJJRRkICawJKHvYktrphrotm2aPQEUH3Xs
MKUTy9rLPnCma07IJyMEksZqWeNZPvp1kqxpWD0ac0jC8fr9xioFPWN1jpvi
0LzwP/KMZ4ALbhH6WbZVJ7oTp8LRfMuC6rChIHbJEluXo1izFBOmPGrrO1Lr
GysYBK2/IZGiZjxrpxvqDz+9z3pDIEwm4WzPg+tyBNMfj8CCVpavoBYv1TkZ
cbwVSZu0+uQRQevK8xvG84OXlYQdw7jsA2tPBwrobcbQDXrUr8dEBjcFGXOa
ZXuMvo5VF8icCZVItBUxMGEIXLEBVKaOG4tNJ3AjYAm6sSXq9h5e7Mf/kPXV
D+AAiRchCAb6F3W83HfbDVnmxI5WOZbFJR3uNqcnDepQvLqdidM+rokubg+g
N6gGZXmzWWbYzARrFoocl91MC80HigwmozlSVObCAaeHYgwcDE12JF5bOayY
9oHloSmWNNwOQ3wB6yd6h/22LtmFEB1YDpxezNXwqUVkvF9SY1rSFZ8ZShNd
H2uf4JPGoSj7UU3Lxzr8HrMfqi/KViRk3o9NlEGkw0khl3Wl9GeGybId4wvG
DndMnpY8Bok0XCfzject6kJVCWQWtFGggJEMP3pP4Atshc/U7R0wnGBpFNBW
0s/wZx8QftRfnf+6UVSGnHcRUTVWFaQBmWxYnddcWutigs7+fEWZ90j6VZN3
yDGq/zvHr/OjhWis4+rSDUG4Vqk+fqincD2PJiv3NQttBE4QEltcN4y0Bnrp
DAb+QFK6nYOY8+Br6pFc9Ira85B5EfXwBwuY6gZHKNcAyZVI65HQdvHtgCTW
G+z5nSDH6FuqaHSsfvi1VcxDpcVx6A7nb/35djVsd0Etghbh6mqqoKUgApJ6
bt+2ve8IB9Hw5hwjC8lR1QuhBSVmM8xsNbK8zwKAjzIMoc7xYUAurruBuRrW
4aHYj/wiR3uw8Y/3T7PldScfbgCqovVwV564aBpQohaG0SHr1kCmZ/vr8F/J
xUHa0vXQhfozHYQh0GAtk6f2mJrs4e1hBOR+RC6kulh6zVL3ZO2T7TzAMlBB
OV1pEksYtO1fH/tc4HNjeS39jMHKKazLiX734AlNgNjSCTZQAp2T0302cTWV
sYfQsGWx+O+/ZDrUjvxV6aNicgAzO6RAtZXW9Ydc8GP0Jo48Rkn6UMvF43vP
pPqI/GTdOPhj9gkgeJDPi2nTJarX6BlmospW17YPltAiqdtJ/077WwwEM4n5
y67RK4rlx6b0I40kmPtpVk41cq6SgNs/zm+TeyVx2vC5+m5WhkYgSokx4IMB
1a8XXnkk9WtUpjcLX2ImNXgllpacN9v2Jn4CmL6WdaUDOgB+F8HrDvBmHXug
E8/9tol+jH90pSDZNmjB0On0bY1fF5qStONkvx5HuOANa5kDQZeKQfv9Tdg0
xDt9iyQp4kCNKAN6pR2PJjPkAhJn2xXO9/1OehPQyx5VsiB1nSSsouI62osb
c7XBNvXKU5VvThg/H6icxIuuc6gSkDy0uj4Jho3Ip9wuxX2A14xz3c4JmvrX
u3vISibNbfmCcT30FoQa87kQDwER9p+v9hpHC/wdx9+nmeIqNjpSFih70Ii2
Kdoda79c260nbhXNlwuapdesR/dZ1R8zizo2O9ch7Gz9T9PZLqofnYkvFUnn
QbjuJN1gy5+gZOnfpQehqN3/L0yCOU6Y3L04Lh+aeAeNknRdvwDAahfsX8Um
P/AtWzJhrxEAkmn88uO8OV7wHfZgdcPL9akNCKMSt4xIGj0oGqOmpgL/gp7L
hP0WZo9qaGE1fl/tgeSD56aEhLpowwrHlKehIvghm5eThmFI8uZ19T7e+uZ5
IoZ6uGBlGd7etw8zbY3uKXpTcz/yP6PC5nzQm9EKETy7ge0QG4bisOg3RwTS
d+5RsL9IWGy+f6YYekwzBjC/hKLtXIuelDR91R0h5dGcm5ElqyrGExfDlJWC
7L90yTqFIH/xtj/tFc46deRG6HgUikluxfTUKDAObjrhoUyqKYo8Ohc1n4nH
skecmcDAFcFCH2VXCjDbaxZfHkXjatKvSEmqi2q2t9WPFAfbLKov73JFsAai
JgHn33drBIY8fL97mPTSZZrtAEb1sKWfU3VACb9kZrF71xTlwP+71I47mEK2
Hk4CgQmDwM45WMlsr80n7lyT+4xpZd7DUxlJ5nvfdcLSt4CFvnvRIVv1jEmZ
bRN9vH6TukqQLz4qLtedp4Qvtc+Asb7bHphu9WKyWlS3VBWf/rOIRtdP+y/L
03XLleqNnAXtG1LKcOHz6FTOlC3KFhWf4SsMwQL01cdpt1pA5jZokCwzBiXM
wka3boCyId9+/OP9IrAQovYlrR5GBSCJlnJbq3XSy3fFiaY7vmWk8vRoy19g
VCcEwv7mCMBmBt15doFg2ml7TaTfs4I2YM7s0ZsZFuC3pSzqFMMfo3ZGRuyR
kvidkH2pvHSReZZY4vkMTh7J0PJMQrDKbLAszI6paOoiMsa7icMIjBKrCKOf
ChWRCEsgSSH2p92H/RrujyDFJvm+ALbapsM7Y5eQtiBHsjvUcLHlw+asghM9
KFTKUPOCbOEJc08z/zA7d3RsJRFz6lVBs7ik6KWjJ06n1mRmB3BTRQ6NBioh
nUJlz28wGn6xLEGqHM1WSr3skP28baOuF+PqxkJ5HJzbe6h2ALRJO4XAnVL7
IFhCytijwbnzIEKxK+Qx2llIWok40c27dRHuhkoxqKSJFfO1wfdXtTVeOZPb
swehPSmtAufJBjY2sMNGrjCffQykH9gHxERAHf7QiwW16732AEolD8xEa4d0
WZRJ2mzo6S2oCe8/SzUWm7LjbCqHoOhBYgr3VJArBHUdm5vg2kPNBPUHPDTn
Dffn6sw55oFyXceWfRhMFLqz+TM6Mj8aB7gEf7b6nDbLI9FlohkICbAnRj/D
1l/JlKpYE6SOG5ITkeehWiphA5Fm0mgdzMkd49H3vi8+JVvkyJw4cQCdhiEx
Z69RUCq/otV97FiBBgr436sYwkVJcwKxhjhUUhXWVet71fol184n9hA6EjxZ
DwVuD8ASFLrFohgsHq2483hVir0WfyscFCzO3kyu+c1SNJ971cWM3QUcQqfI
iEq/BHypHTxgNjOlAAjuPJrZjn41cBqx+1+EVvP7Ris6AyRN62EQdeY513CF
dnfB96e5lU4Gm0HSwmH1DFluL2yR7RWLr8ZrARXdTYKZEdxJF6sztqauFPOL
r7/xth1+EHKryzApnTaLHwI0hJkCYiJkfCUFKcRZkYnIcji3jJL2uU5mNFCp
/7RNISqOGdtjTDz1faMzPsfru1Cf5YM8+FlWeY6dWAvs+ZBL8uX1xCM6ctJG
bCnkkLKJCgW9ob8thZHcR63feOSp4BqA7ZeZoT7NNX+FmpjP1ziztH8KG/X+
kF9vtuBnqESaHjmjiaa44prxyPhDbSmOazjaRAelooRJGSZf99qmgD0FdWZ0
En8PDW69mMHjHj+Mpb20Vm7uOsJC3TBAXKgfdnr007Wk92AmMwoYvGYZovgr
bO8pvcu6+kq2fFkwStZYxdEMb2djv0bMtft70Zm3yBEx3okQV6hOfvtEtQ3b
kk0CFtSM8MyP3KfKLuZ8tmoo36v4rnHz9OU7rXE4zSyE2VOlXwE6/7juSwd2
uzzF2hrdS7SxnzmpDFsXosCQx6vVOXxht6gdyPGkjY6ISjXMa6lXsYx1AChH
wuzrX1fZRwSNexVFrFsGYk/3hffts033rLv0OhpKcGuevnr7pCgwumGaifBX
AnjQJV86AYESh/RN3XnxCkO1+ZGkEguJSMIEgqaCQT6iYiCI8Hj8xSdyAzdO
RkfP0Dz+kBEkOiwCbO3+w7sYTkit0dFi8wR4+i4f+OCCgqE3xjTIvuRIkfg/
jHsH4PEceqBWXljzbvuQLXveoz+XVDTI3GHJE5cUTHCh7QyY+1f/1D3i6M7j
jsxM4LYkfKxWc8TL916urEtC0G2hk+lLlWqGILO84uA/b6oVn2+4iBScndnw
Fx9B3/DVRCH+mI+W7NwMC8qYES6RSSXPhSOrsp3x0jH8hiLXATGFfFuc86P1
hteVYKsC+vVtbJBdhTGI2lsBtQuLXixzpNFLvmRJz2adomupzQ90KsAgdtWg
6FwFqic4P+5uCRKmlQkFDSyQr05D+4QYaSJo55+dquOmzCfM9VW8o8s+iZKe
Xai6gBTBDoLi58P8KxUrKhxTtSX8ZOEGpMVEURwJWQyBdrOvpJHFTiVubM1T
wFO4D2S1ntHzq+KA82V0rc75KkQDKjd8SnDfETc5tx+4SW/EZ70a3SoHFca0
5SqmEM2EHTXmzQOzNtWgSO7k7fBuZeDRy0Cwfijj2JeTZ0IwKxq3c6/fxQQc
C/nsNBT+mADxkc0K7RD4TXavU14UriRnBORWb6Ieql0l7QPV6D/JY3cd3iC8
7G7qXxptUusSmmvCmU7MlM+RKRRB65/Bk7HLbMmsfq9xm5hICaHoOa6OkhDS
9lq+b9rhHjO4MowAEks/gNFjcUfF/bDyY4S2FGeS17wY3q0d1x1kFEW+Nmn3
QdDLeeAQzzIheqRafnQsmfzPDTbbxN1hh9Om3ym1uZkq3YTkWpf1GAFVroMs
PZnPtKq/dI3s7PjxG1pZdvu8609lymBKWO7EzgYZVs9mi/Td+l+ITA4WJOk5
546dAexjDaVcWbqsA35tHgmNaJQMtW5aB6UBJNtnbbbThcw8MqoLoyRubo5N
83YoQY+7DzUVKipm6uU/mYhIAtiXaDonyqVELE+S48EO8VzKTZWPAX1ElsfC
Wj/Gr/CGdlx/jKICmhdBnZbRYTds/Z1pch0KsU1oQSeT/XYCV4dJrJnudehK
Zp3Ds584osHq7gxMV6X5rqtkqkOU5NoD0/ydrfqmxERPD/r8U5Qe6iJDB654
zgXMTeQ9e+s8+u9HwOJT+WbssFd99GwYMA7fVssnaOm3AuQPFMaHVR7y9kZN
V2lz7L6KVvHsctw2De7EMySQlOf/EDkKnVXDy+YTq3HdBAcJG6AEnh+lDRU5
y4FdHOsq816Z5OAle7uOwFtltOVPO+kz5KvPJhFUCTSVLirSanzQNJkcuuVe
IyrqQte8Aw3kGt1+lcQO4RDx9zh97P6JjXdrw+TYcL0QsD82/SQVJuZKndM0
NNPOZ/MYrCuG7oq8tOi5KA1cDv0MXXaurBae3ZFc2ZF5UqZjb0bz03z/pcLF
geFl1pRSDei6/L20kHt6NuaaBUDFPuBVIQfBLbCCBvzvV47FYybNIdbrgjU1
zdcAkTQkInc/h+NkVAzwVvxRxBwFi+5Ny7rDxBzE68JRTtLaiiIeHyZ7ES/M
xJAz4DzzoBb6JO+UbIGHncHIPZFvBiXZhVsNl3uUFqtZs3d+1/D8wLAPRHCQ
yMa5U7gChTM8mayEAVdc5GbYPHjgEof/1ns261oLcDg3dA/qYc0A0YZmvtnY
X8SQ80MP5hr3F5enhNglS9mpQoXuze6c1fBnnHwyt/OQ2d9rMNGdbbC4EiEL
F7HdTv4j8JFdADNNH30fomN2xfxadM6e2ZEE25qoc2NebZS+KayKTBh0Tsyt
YC3C/FfgHtinR8RtrgR3UTkvGkpZb0Jy9R4NZsQF379ZsbURlJUFL/XBw99T
mV2wgEKD2mTwq7poiZ9vIhDez7FYcZwRP/tezsNGWfu26ghlYy6VYxWYv/m3
sshANcBqj4XazUz9OKpmeeMzqhvFg14M151r7BfXMDiMhecEqas3MZj7Bk96
gdSL4x0FKXT+R/cBXmhaez2b6XwwYVRIGZoxdG60mpwQLI1ozR1BhL224Daa
6bnIOB2kfedJpVpuWlYgNUU+UgpRNk1h99OR+MoUypUrXgm7r6lKgQDUTjYF
08crkCDUR8RsvmL7Izhu2Y1FisGnscsUMfrEw3qUfqtzjn2mhAvn0/Ku3PDM
ivNvC02eBBNKJhhzA0zufErgx1rlKJ9hBKorvMYwcamEcGO7DNX+7xmrn1Cx
ZSZHQVENdpLOjtJbfYMna/d5L0RhW12aH/lV8f3i5MMdApetO80QnXGd9vNf
lMbH/OzS/khZ4DTWY6tb+0nR9AwOZBTTHb1i349vxSxhi0YUefJuYZNkNU0b
xE9+w/Qv4W3iRWsKideqBjiggaRh9EBsrDGMau8LNBDpj/vXECUXdfV9jnMn
6gBnMDS/tuwvJxG3zc/e6kGLnlXBmBCMlY+LArLGMW5yCbSkP6SVaodm0B5z
UKP/F3vsVYDN2QAn8rtYMY0RClXL1eL5J8W9Y9DTNFhjtMMtCRw2eFyeb3DT
/dIK83XnB/2ciOoopv2lYSS5mFM9pcdwIkFHoorvwj4wB4WBl7uRLMiZm/lE
BhNZz7fFSQ+OUCfyzD7s5tGkuDiqmrF+nDMWRx5CUywEucMlg4GgoLbomP+E
PMGvfkmgSlap7DB9BdnOfhBwKyMggxXYhnVua5xHNqgYn1tBjSDR8ZVk/S6R
GDzTAZ9Hs3Zn5Qku+bZFmb0jr/7Lacjc1jce4yURppsb09huiK1zg4avJlOE
oGsDCu1ii2vechfLLfYS1QL2+3WvCg2NlNa3Zwe2KGEQhW4L0ZzERaez+hcN
iNvQd8XGcSTGXCLtpxrFTVKxAredIpBf57pNLPbe0cw6gICZbq5ZY13uSiXT
FffalELNx3EnwGt7D4JixYU1Wphj/PJgsoGWDlTAAk9E6sEiOhW1DovZ74Zv
Xum6aRl6nz5Fu1sgz1oco+xh3f0R47aYQopSKAedrlGs7bX0rMHh69DQAkmq
XACq9ja0bGwgctpaNl2C8RCMeOUfXdFr3yZNLO7a1wZNsU2U0qK1/F3ZjzPN
xeqKSiUJPid6Mh1C3DcCkx/DPEaM0tbXCpV1XhhcLVG+KvvTwARcNtlL+ttb
6EjcywDpPxd2/kOPvHK+PwaDidoZ8OESDlKctTggJpLl4KGDUMovxpOiUzj/
xUj1h/J96EvVBu299aNmj9T/OWk+uizKbzeV98UX1664QrSXrkRWsOiIn3N5
wZdTPT84IaVftcpCmCzZQMQokKTYK8xFeLUxUalrLOrH6ktoZ5NfGr1J2IMf
kPxm6cTOl4Ra+1jknaoh/i/ohPGiLdzj+Chd4h7NCi1eoiZtBlmyWV+6lhKv
KDwwDgo89kWCy8v+HVmtod69lteujlbwBk7iqqugOmSD3YaZ03L5/Z34zNdT
khhiWTlvuamjzOqvQYVRcUQqH0ZvM5G6d6OhEIs8yyUu3LO+D26m/N5VOehm
AopcR73hR+KVcQRnpODpVQwcerpJeYgzSPXnufPccbTOe67QvFcrx2v/bOMy
QeTETBPsb3EaH+/aQ3303rvcnwdEC4O7hSpiIpW1fVwCtMDTSaGxSKXC0lC7
dlmYLMHWzBdMidnud0l5iZxAb5gpXvbGixVdd+BUCJn53Gkh8Q+WzYzsS1mi
GsNGaz7XTGk+GYNnABn87sIgtiXgoMnoKqPnZ2q6MmswNb3jcKv3p9G+ilTG
p9sCtLvKWCF7gQo0HX6OIVdo1HzPuGB3m2xL69kTO2kUQdeP4FLAUCrDyIyE
TtQDz8hYShyGdDKc4vg6icZmeCEWAejbbQc2Tu94pKIa4iuD7YTAXVP4zngB
SxcFsUFsRGcDssAWs2Ij4fornxnTHPPf7y1q9lKkgzkaHgD8RSdVpnoYMUWw
lZWs3dDQthKVODo0n5G+MEY15KwhIm66zzCsseYZQajAwSa9IfevaR3NsAF9
DcAH0LIUpFQbXlkJs7fVIuuHr6GDuYEhkEXtEs/gVHfIJH3y2/QZlu+kf121
VW7T+vDVteXPgCCoJsfm503Z1Nfmqj498yixlYHcQHaAov+05YZ5CsgBuayS
Ue/+LYsZ/8crSdsfOVVPEHJv6mESs1ocMHMaQWZMh46vTmzedpkDd3TAhp3W
/KJ0DV6P5saDrV7JStQxuXvsA9kvsx9B/61SGr5izJKRHR8j/G+wRR8JbqUa
JNTBIV58JuJJIgcZIbRZ6sEwlPAP1G536w9v9Tm0gTddXqxPf52IhHXU0ezz
KlCD+eM+2rFZT/1zdsyGA6Rb07zTJ7yNpBRIa534+c54fyvJtQ9wH3oMAEMz
+4hGJdFLiTneiMhCm5pnl2jF4uwGQI52t13rT8xcVWbqJF5cYWHlSCYQFNBC
AAbm0bBBrM0lH5+EkyFADb+zEvVRvbfBeVs0WKbDliW+pialbxrC2pHE9Jsv
bV8NO+xSTiFlbmI7yU8vH/68lqbhTc8Espqf1rMtQYdF7jK/dbPT0HLNPUFK
0CX8+uwPthmQr9LSqh9Ck81+5LTzvnoXPf51LlLBkovFJM9JSYxcazBctUkR
sfzLBP5SLBJjRZVnrPrAg82Z2fZNtuEfydbGlp4vJORtc/7ztxM0r2gG1T1b
iwIPBbGv4KOoc0pgVD6Cn3cnrdXu/T6uaIqvF7hruMbDd/Vr2uuc9H8m34qC
gd9ZGMYK7Weaod4i9YMGQqfpBFlOr68o+sIqmgEYBfNFCeAv3xs+FEVoRYY+
D/fZd/k/3w4cuEhRU00RyOsIRxbFnDVG5IGArJ5mIAOb7ZZteBDCkfE45XO7
sW0Iy6B9RAFO66vQmlkPiT3vDCsv7V+xiCVWsqGOgIxPDqH3VKsA98XiZxvU
EK1vnTL0t+lg58GGnATXpKhUIOnr/O0DoXNPfErQ6qFQ88XRmChah50fOz8t
O0qVhiApEmyx0/WRK2cnGTA7QewQvzBZeP+3lov5Gx4I5ww5N/5PFs/lO0hA
jpICooiChG9wZsP4S3dsnCETYOnyiQDAaOMJOcKkaD0VS39tkuXGGoBmoPuQ
QV7xvYjTDrvoYU9FK9m6qLr1jlIM1MuiATtJ24zuMkNvVo9eVVm5EBUYZmpW
kI9QkbWV78UDIlTF9vR4mSfvPcs55g6VKssfU/tM7LNGpf0N5ZaeJhrcu4Dr
EVEtZJSd8byhmdJGb1S72tFNvIUUSzD2BtDDw1qRzke8A3aUgfzP53vkS3AU
bwqvFCTaNcfiyFQxYKI9HE7DO2dbrpNTSZjQyhaEcueTVusLAawJNAuOHi3/
UVqKa9xVg949IR4b/FdI0xcivuNVuYmbWS1VyKPzE0KmmUCm9yncefS91CLX
QjRKgHsrX8DWzdDWREdCA+XKidQigsel8ekXLNeMWg//DWzxJ1xjFs28ELPo
8f7YCJ2yKD6IHiOTFjRZ4N6VMt0kpNhxp6sQlMVuK8o3HTK8tZ9A9e1Ru1ga
IEAFZWZaE20GeRUbNuJMAjRl3mLJ4b0WmNqLVdE1TMveUL5iDb+xSdjfKt9z
JXiRcvMgL4ClTH4YPxUMK1BhRBzGNO7KZMqiF+hIRzVyLWKZYcKTlK2qhT9m
do4T4aOSbzka8/ACE2qGs6wVFeuR9hyEhm6QPkRrwi4Tz4xhIaGB9/tUq7nt
32zD9y+LBK/wAP2qUafsjAUm3dpffIVlR0wDRbl6CGTCJxRRlvBhEn2AQ8Gh
gd44XSDxI1/QEMjLB2nsr4djXi+INBLinmcryouAygMiCp6S7MBhYyBkNvMq
1V5CuaABaPsqs3Yg6OUL51Buy4wKgCpMReqtzxmgTngAvjaAaCkSn7kWKULy
LZNugwf45/VUk0sR8EI/ienm4tPIA88mmLOwE7DH1u1Y7LweeR9Yw5mpou6Q
q4Z76/Z9/STIm5kvgErXe8Dz+fR71Qn+JZ/Nnw0roUT+rfSaKwe6fDWl2mag
x2v+H8hfn7hsS+iOAcF+jibNfpxYocmjLPRGPBxuqJ/lMEpGB5n+xouiE3h4
LPQC8jkB3d1AVKcuVCBXlOYJfJh5sPw2+iXsao3T5tiIJSCb8Vc28ru2ZG4y
QAlpyAANe1u5yH7eXuS+YZArO/hUfMS/LR0N6ulzlh4LRZ1/DtJmOjxkUIPF
HljrFNs+RtBbqDaN1v/K6SG2gTP8I6XLsZHRGzUEIPScPxAg/1Xl6qnvX+OO
vBggPL6GPewuIv/3xUYrSpCvuGaq66JvGiwkWca1xOVKiawZC02L/O0jhWt5
SBCuP7qNUEikaKNP5Jr5hOQs9NbFdyXqIcJhunPazGp8D1Z2s01vByEKH+rU
3sFAfssOZGnZ1Owu3aidkmCWbtQ01CBx5ezVGFXX01kXzwYApIAki6iqWPJb
roQ02DPNebLMpLV7apfqyJrMHWpnRMvTuhHGp0p9RIC4zSm6YmD66VfGXkvF
SzlwemfBWo/ZP/3rUdummfrX/V9B5L/PHMdX1MCk+Hhpc4J7sk638wMqqsSd
7WTAt81ycAjdFYRzMTemTfHTzX4okvz9jspCdz7B2fOr7Qy9HjWIIlMKObS5
+IBkWPw3HY+R0bZbrvq7fkrcW2qKOwixhfaOxyw7RBsmXLYtXVtnGZ0kz10k
4IclLXGlM6i7Ekqukr4zNZcUtQc7nwfHSXloKNGk2LGl9u+Jha1WGo47Iv5x
p7sY1Cx6gjNkcRQy3OsErrS/1ITTEjQw5ArTsVTzkV654yID0CZMDFZpvRf4
j8O8t5+T+X5nb/aymvcYItMLa/7mH29FQJh8v8kju/idfaWMns/kRnIvSIOX
3eIZdIxuQYptLlIt1kHzlPZ7psmOsnRCXiD4MzIww4/NoI0F/eo3b4TnGgUW
xy7SvNnON7CPKDoE1p92SYOd7WNbT8J+SQZehWUbD29gs5WtVjLPtMBoxGBo
9qzorTzmROtgNUyAcuODkTpsedKaWGlxd1j1AIBBzR2lvKoKIlG4YymhhluG
lbnb1UcR18TN4AK++smbo5PVTjhHW47a2oUcAOTlMU0no7LSotQafZC6a4qf
2VpMRkfjDQogJL3wGvvfAQFYVY71B/BO80d9aDCZOcV5xDGw2VuvdxrQ26fB
skIXR33nxZ6CK6K8aNM33IhPK20ik/+LqgPUJ+8lUwhuj1K4oWHN3qVgyr7g
yPjJTJKMCjY5yEUfgAjRg5TGbLePU1CSLShtUVZL3RkYec4EP/EXMnDR0Udh
psZXUDOZtuqTjCvQGAGP4uxHgYHXnJinQybpLUFdbqf8hm5HLwxS18aEsst1
XOB0M3kuxBeswkigH7GJoBGSNNer26YqSgA5wQeJIQaqSNwTdVxZGp4b/TDJ
rLMH7I7jchCMaEjIbAEUfJb/3R8nNl4L6A9uvDgtP5I/zSCFpbwQ6vIN20ic
sIIWMcZqzammw9UfTT85cNY//M6k9bKLeZvZZA30VD7ImeVTtKrKaZQGv7a9
V5/zRJuT+MEDYHOMlcl2VXH/gWPyfGG6tDHSA+jrx6AflmHR/g3lxu9Lv+Vw
KxcJCv3MDvqU4Y5EDWeSJILc7js7Xggl6GJZ3W97lTLWnPW0/C4hNiD8cBYT
vsWEXoiS2BWbjJz7UY0liJytoN5ci16hPTOIx3UGngFpvf3+QwKdx7bztEbw
/wK7yak9DhkXrtxBw0G3CMCJbNB3MsVyQO96nx0j82S1kymUO0zYpaoWkB1+
AMmr1+l4rge/G7UWLIebFCyEgGObnhG86sxNKXzJqha/8URZa3pY9JaDN5MG
34dChMFgUFi7WvuGc/Ofz7qXT2ZbRXg7bfMeUai3rzg6wNGnAjBry9o87b2W
TYwnlfm0VFX/uwXpv3Q6rTMupdi6lOf51QKYQHJxHaC9n85jn9nt8YSwxokv
nRUz18RTD0U2yTilP/MFWMvIGSI/0BNrkENjt1n9p8bd+F9OH3LQHhGl6TB9
AxAVs0V4rRXQ5tQDlXeKI7rfwOlx3aEGXUpWy7dn1VeSAnzT9VwdhZ2PCkYW
z1MHb0+bvs32ewUXi+MsRmaNGgXAeBlNPrAemWtuAQVxmPfERJ/SeVskecZS
b85B660DtkXBdtKFLlL1pHYI4lytsxzyZPoSNWJ65JM69i2LrIz9AAvbRfde
F6XW1epC+NYU+P61NvGS3Ds01VQJxBsG2fNdkJjXiIhH9wPnXzrTcg3jXJNA
tkGtohFtq3ba5yEBFwDel/ueX/mp2WEHrX4BGtBPhFXYv+1EEYQibGhCmXwP
+OKPEWuwtq56aYeVuT0v4eYAzBqQiTdNLHMO+qXARBHReAztmSL/iI6VEAPY
w5GL/iq+ZBNuS/VgCe99/6D9Rlhxbu4DutqdS2CU7ZsCFIbC126UvqRxexXX
gW3h6VERgBp/uAV2SXy8neio5kZECSliOlXAwe1J6VEs64Dtanp/1PPGY5J6
V1xzEefb9Lkf94QyY6FKDWY7qCHhev/ng+jYFjA2e0frssBdvSRg+VZUUE4I
5okMzYycn/9tfqBSspv+jw/OxCYqm76kOWHRIizTK36vxF8cpqmW6A8WvpuX
XL+oWbQMyIZFhks8KAS+oRCsep88i4085NQoQjPdq0ME65+OOaQQMyIHWuLf
3aQt6pczpU2DYPEuKB4Nh1uzQDu7ef61kcPE7c9YiK8VDMuF5mKI23Ao7Wo3
B6AbloKMHkItKNkk6+VF8Xo4M6ASBb4mf6EcAcFve1JAgExxrarnglKACbkf
gYnpO+PIqgdEqn5WNuhDyaZudXBCuiWm2J+wwIwcjregWmGaJhBV534ydryV
OK6uelB4s56+uyKIDXkuPXpPq62h6BA0oj/ZxI0JTY+KnFw5EBdUPDNHkAOk
T4B5tutWmC5jSCZ29/2tLzipO5F2twSye2B19KqP49fwIggK9pliRXPfoy++
FPDIuv3Llcnt71HnywyITs7jQDwZVXTAZZdOFyiqDOtLVZnHK2Z0v3V/kfZ7
+PLi3hDIDwoO4pPYOa8Lt0JQrrQwfFPWLUyhNFjyGvaKKvNxrL/CyGgJx4UH
75rvoI8M8B2tLZ18u8SrDJvbTAU6Iu5BwRdLPc43Rb9MpDwLW8kCjZBB0T/U
4IbzoRU+XJtLne/SxTK9GYNkU49K76GF8+0SHszHQSH+PiLonvF7rNJCBS3O
vItzP47GeHL3jNJdZi3OxLepiSkAXSJ0n7D92KFmv+9da8aOx9OSEecJXU+m
XCD8xrBjs/3O+EA+CmmflQb+0Sk9qmu9O1h8HP8pb1lo/t8yTG9BQBSzT23Y
nLUzWxovQ7/itR7N+p8q11yuPBiEttSEWbXZGqxLxm4uKP4aTWWasA1OApX7
G81UIWGtezsDj64oUxjPtlwS6JXgw62suQDcEztmmdwCBT6Ri3Rztng3k2mF
52sWpCaE+gfwbUVH3FYD83zLjpA+HoV8BANAUCxUZ8JF112ECLMcQjj5VeU2
bu8PLwE6z6u0G3xmTyTRQ9H/jux7CzNNg072TLPu+IegGKEsyuNYnkXa/aP9
/3NZex2iVWAc9ARBARvaQ1xwvGefs5g5KPNQuYGgVsrBn6JI2Qt4rA8CJPYu
kfBe3x5txaLwo40PTEvTcC+jHU9M1Uyvg8WJlm3a2pjXmrJ1DF6RrPMg/842
G4N964q5bkH+WLCayTamOHlpG5/8fbhUG34gqA7guDowfI1SWO5Myd5NmnlX
fivSSjRglvzRzd5bPcfGPeqxJ0jxzzmcIedtimYyfIUsWogGO/uR6ELXImBX
5TsBbMd5GuokgBMDsexQSLnZ7XemdNPKF9kefgdRd65fnRwZaDn5HAdzVYCR
95F1HNvQfcqjTEQlHRm3sq2UCcAo2qgpq6vZeJQ/bZpt5np3oZ6wKU0NFplK
7whr2Gljz87L+aozcWMrzGuNgvuE/XU1RBSxgvrojR23oAc84xFxYN00PSN6
UX6S/i2WRIdFtu+rV5vos29T7rBkxvxyVtk90DmCHlvHjm0FvwRfw/2BE58V
/VlAQcpSb1a9vO8C4OWPNKSr8x1H3TX4srMagJgQUs4U+7AKh1H95aLNlPq4
V244Q6Cn4Elw/vrGYbJavjUNrj1UbKSXkt/rGgn+an+zV76lHjNt2phC3UXV
N+PVtjzwucfldH/oiHDK0to/QLZ3lemZmgq9tv60vwGTzmQ187xtUGPAUL8l
QdxDBtu4XzPJ5BABFl7R0LFFPW/CVpzRsp6x7JiBe9ZWyubbhbYoQTMH2jtD
baqN+ooqsxwOQyqXz1GMVigrybPv0FdHQoYChAlSSCgFqLrYZmIIgms6T//v
RbuojRxvbOsbGucderd12MiT7A2NV8YP/MMfosgsOa7QnAmaYyppssY0vVtc
ePTYmeXjE9WozGOsfz887MqKcRWik9GUrkahsH8M+XxYELiHIIT+AOep/Ql5
Lwyilykwe95y33gClQCrUYfpOg3uTYiubWRjUlSb6RMpKjZIyxPQCAGg+EkA
09U3AUI6+AuPknAxGCZ3wZKSFxHiow4l/yEJ8cKyZGbduLVQBE/5YrhWDDxC
9vypPJmLjFnPTxJMEEx57BFrfdZ9W2rw9xRQwzOnGA1WMt0hHpB4IVc/Utgr
G8zHPr7AnNere1BcTJO4SSGszcIfV81OzeHrWUWqYzgfhAQ27+9if+EQzLiJ
1rYT97iV42YdHd0gCrUtJzMv2wWAtHW4G+gPbjp1ducSfKFGoI2m/28AtSTh
JjrnRJbNiCjFcE3wxMGnHeIjG5F59RRe6InokA3zZK4cTQYFdBP1ONXDltvv
LndYhrJ3Qnj3dHLo/A2kNsF5bRRBfFLopgztAdHLtR9X+VK54YOrvNVlgzg0
2IClpyafOVWoadvEV0TvoOSLxnpUWQitxgx8XEE/oZo4i9dGf8adVNSWvWYF
qYFXVdOhAUdeHm9r5iwLfgFaZBk6NGAMYmX4/htDNBYlSJ3ZbgLq4Y9V57KJ
uzb2zW0KISrcBZ6OPd5luqnWIqklsrbZhNK37EKVFpZvWvpAbSnRNcrb7q1t
tYNh5O3sN4Ds4h2JnV497tma0BrE6QZtgn+r7BKNhwXQaQQbRhEIEGtwDmWB
V2Mfw9TjB6rPLdIHHIZMmLDZ+9jl20CkrMndFnUlXtXysqDBDTdTW5TJ+5L+
HB36NKw2zoEV4cFnXjEfxU/yjN+YrxqJTtiqCnojD70aPQwiwCfLbodX24zC
7WEQscX/9dIcFGMCkR7uVgX5dzrhNarvTvhlL9lAI50qu4UM575U6V1VSytq
ZxwTZ4F2a0c+rvwJ/jLnPdQW2cCG8S//gxvTK4teJNG+m/xsf6KF6qwa1/qd
wceiP1ygMKg0Zyx34ZDdk4phjOPLfBUZT84Qv8eWuPZbT4rkzGckq7vDy2sX
aKhOCeYTmMZ3pccMwC+oFNuFfsiODk1qK8c7KYpM5p8vkJK+aObtljLkW+Z7
Vq/h1LEan5PpranKC/RfRwF0X3RDuQUbIyXx39T/GpL9A8quYKgVi0pOOzHJ
WbaSHlMWWRmoTA0cB5inpVM/2UcsDIMcO9ia07wLmWI2dqjqN9hnpyAHMqbx
17yh6YAkI35YV2lEllJMGX7nasw50xAFYhfKnoaiaup9wGCqZohgffT+/ggU
S86aCsiJ6SyppRIxUPCvDqScCGqPgFUPJ9b/xYKqiLb0FJCOFinro/aUnlPB
odU/nSj8GncM1/EBBuLty3cCSAfD4jQRrByVyN//rciQnTmNsBNOXkS7yI/K
Qb1D+Xp5CQk+9siLt8o6ikoJ0fW9a6G031f8WKsSdUNSAu2MF2JefxaOjzPL
2S26MlVTbn8OuYutGvXcX2wpnQx6tymmimTYNSfYi9Ob6XYBBKAEd4v3GU8Z
Oyw1UCqjG6wltr4EYkbkWqLWD2WFTRuRfiW29WnJsJiPE4viJGv2rEeXJWvV
zjC9ny5gjtlBsF1UMHkdQlTrIIC4Red1rdAH/qm1n1jOt/J1tfOmnSQYXWWC
skYphOGxgPjSwgoNjQOnYox15GNhOK1Fqb9q/qOjdxaLl050z34v99Nk9cfV
Ru7BSsaa3ljZ9U6V30aOx43ohCCFWI8L3lHxQ5KeXxTBCS2fHvvymeDC8nj8
8jVSpit/but5we7On+cKXgoth92zdyVChHdTQGSRpkkHKHOmpODWxM2xPeIc
5n0ItIcqrYyJOJl3yjzmab/g/nl+4VoY+3a1hdMC4L6tZILBNvpO8EwPdQ0z
Sq8q8kgG4nW5P8szw6SEf2o3Og/TEiX51A+7e1jNufEYQHgfD4+EXv0vVe8W
fABN19SL3VcX9CQwrfDoFQimbPlpTqy6gwvdxb2HnB4dRFafbgVk9iBKh55V
qwSD9A8u8ifaNecHPoUoUf8UmXtJVxwwK7TyK+jG9qZDh7jIKfanHy+aOM8C
+l1v1t4wfaazhv8d6TpcjYMclhCGZQ7hZpyR+i4MCSL3T7M8lrhop0qfyRCg
KYPapdvv2r39rP3HefHbj5/wSHR+DVKKj5ici8x+qC9pwkOcTiYb+HjHZYwm
QWq/NWy9kg7EG+FJ3sImHmTeQJDBbDPg+m7aUR+0Jz0kJ14jNZTSzwhX4ZCY
hrjoGhAp+Akp/o9adAjv7IxVEoeKAOB5g51q/GMqgPd/Jd9eTOj7kw7ffuah
D+kqK6mqS584LFEoY9ch09Z9OYN7LwPj68sM6t1klC0+Ky0nzqOAc+aRTCZV
bY0xCPsikWCMvB2czO0/jY7elBPRAeohN82oG+zgENNTA1ravuSQ3QfHjqhW
e5mxGRVuYkHOsOkszcY2Y7bBwUvm2Z4bYj2Kvtu95h22Ow6BE5ID7p4/towD
GiGpUxdYpa+fKrSqNF8FeZHv7TvBCdQ/m9xN0r4Aw8aZiU0WVQwkaP/RyNNN
adGpxeC47/fL2YY3WhnPHagsjHVkJepnSesF/YC212qXVMeDaUlstU1jomQn
RuKFQ01VzvwWvgK8AeTpFml1If39eLbfK9VH+mmPzuHWEiRRYcb9uuGQU11q
3HDV2K8FcaOdPPz4bJUNnLI4NJAwL5aRku8FXeonRvJ01L8Y/P0F1f4C0Qar
bL7qzISuqkl7h31XUZl9iKaJjEsrT/54T38j9959+6Gc0xREOB1o/eEVq/3P
bcnaLBm1+PWqxAs0koAFREjVoCVIoPuR5ih+12yKXszy1ZYicmURPpoiWc0f
+LJaj0TC9GOCP7ClIB8qLLNvShgi9xdzfTb4Ts5R5oKj/Wwxt/Fu/FIDbAYO
PrLpI2P4IbztKE99PFwC804HfyywzBY7bT89hbiWP+ebRNfIbx8+WEnAwEUN
bEB+ftMfT7Lw1doJa366698RDa/MKbRE6Gax4phySIkPPGBBCuv7zv2ecUIM
Ba2u69E6zuI2QnengzHobd3y9RpaORA1w17bk/Ci6hmhI9Y+4Y2Xy8zCAmIG
9jRRHKH1e0fiJDLHXByZFO9JS/0sXP5roikW4BrX+W/ih6swfowP6XU2phKn
pOT41H6iXKm6qJvddhbdBGMcfu7rYMIVwIwem72BupXPHF/BSuKLNNNTq8ZW
9TQowESou4XKsP6/ES1hGQ8VXh870wdFJL5kkIC4W556RB8dTXUTyn6bhxOG
EyN7wlBMj1FEcyb800sPvR1eLMcjJ+l3dxBD2LUjRremefGJaiv+9NICJU7z
ksE+xs+X5osFqARjMg3FYacpHNQ/5RI5Wj71pWfOhq0Oy/PoS/c21BR36clA
QuNX1UofME8hORZyaoeABNk0zCet8BwGw7PhI+N1mFO+7HEBerAdoJ9eoHOq
oum5BTNEXhyTZsK0R9DD3I4+tL29dOaUQI1YyEI9EIU1QxhpnfVbFsPcxT/U
0xLn99Ga8d+F3ZAGHJEwwXuzkg0BWJhhZwJtwAmMgimZ8Qui+pDu/l0Dnbxu
7XxcePqaHprLigaKFj0BVl49YiqQPgQbY9XBIOYOurdtAe5Fo2fQt2NdBbGX
bATddrP52hdubapKpavt+mF3kT5xnRticmTyTtKlEs5vzumq4wzW4TtNs9ne
7lji/6oGj5JxT98J8rlx2mcZhDmZzZ7d7nW6Y0xVIo6VP7cnHT/XLk7kmK6E
4V5oFbxJTLoWtbQKzwaA4ZwskxJ1wLsH0hIZM3+bdcVXApyrM5lMHl/6hWgb
8VVV+OMHfO0NvMS9p8FFSG80y/f9QcC7Bj08b3obJ+x6VdAGV1tKk4YmWS39
Tf5uBj25xaQQqhaqpO3HvUd+eL33Hf1JjcT/M/vy9RmcDloq99h0iRdc7eeT
esp1n40DCeGdf2b0usXolhiuyVo3CXxH+wwgavkttc/Jb3b45S2C3Lb3o/Y5
SsfvEE+y/s70pKOtBNsDSzp/az8VfXHRpLMRI+PK9rhdFpYvWNX+GpG2NZyj
k3b7+3L2+1sr045CZBsgoYtDVIpvigjJX/+uxXNduzUGWX9qaAsNMuZlPE0k
57w6HThu3Vw4S1SPbmFyJ11WeEXgMM1QAeOIC2ewJGzn0UhyLTwgHMlvmwd2
+by425Lw2nVny2EvH/EU5dGoMdkmj/RQf5kTw3RBEiblDbDKaztbP7hHUOUJ
Uhgo+vbN8MP30GcBwbO+melbosyr0SDAoSVlKEZKGwhsKc9Xvq3uB5QWMwz7
VZaAcq72Ie+Po5yaCv0jlTM0xPkghHcPmQCbDSBeYhBSiHJbt+Kq0XUNCiA5
vBYREiOxqYKoxugjeYTL8OJv7tfIs8VQkMkBNq/yGzh/tAG4vdRUFZsr35O1
u5avpNPFKA3JBq4XoUMEpt52wSmvhqDxwbk2qqO+n4qGI2ulS+cVkOV27Oyr
TbKW+EN5LbSEwLd5CAOdDnlezrs7BuyjW0G0LXuDZfeZfxDZia1xnru/Y0Mw
fjyu6ZChQjvoQYaJWSRMAIb1gS4wTN4/SRwivGex/k4WeItWGmTrIfDxdXHB
70mLKpXpwlgSOIN2OPPA6OtSDrFdaNBl6wbR1AgkoreH2BzZW14yA0yBdg+j
PClkRCPL4JQJgf5PMZyg2LgKRWeGH5xyyu7y5OxFktsLpRI/WtZLo6uc45YA
tAEsxzRXdWIi0MM7GOwQh7wmz4/PfvFuIzVc5mVG9bTJ/AAsuq8txs8zfSSg
J/bX+5eiINbtx7bCA11UoIu+47h7Tn5R/hGAb510E/oZO0m2/b6yZ1DpbDFC
iX7cS/5K3Bnho6RoxYf+SSuy/0GJA4kxMA2wOLjMrOL4uMtaYQoTIdzCfEPl
vQQo9+hOSwvIGR22AKacQ5vjY8qqngFL9Kw7M2jzTcKkiMiF1dAOczEzlJWK
UoN+ZWXGfLfX+K3ygFNonufoUVXQBMYAwlApKhD8duOuFe7dEXZEWfqKBgvD
i+/wGn7thmmQQk44JBy7J2ogk+IjkIQiTlaRyLZBr8H2IWZ3I9WPkZGjDOmA
WqwkgUQUq2aepU2shRg/6ObfXeCj4YKuHnEQxUVstKdoC4Ppvl2265hxA0Wn
bG9AabxKro0tsimSawKW//ca2xgDlRxTPo9tNvv7f0ACoWh3uuCeAnC2DVB9
IthJleVta1azuhum5o9SypywArOTLWzMbie3iDPHXx0SPRTGhVorwnj8KHdn
pESOf4yE4ojA6SABPqmuzBvo7E7O+UDIBpuuYDH5nMQxjg48uhqPTG6R3hYg
JYPQUO9q+2bOebetCS9pp909mFENI+7vHMVpPu4+WxnBjSJn0uLNNInozwpP
CRjRRYmTsJ38cGkRQJI+jHNFjphVAXYc1oumpVHPs0O9rhwFRS4NW5yrT+P3
qzx0I162JxH5lQOT7oR9RodHX/SrfSBWQ6phtYlSjvHdiLUy4c2dw+CaqI6g
3nVNY41AYbWaSzb8B+a81XzoefAfW1u9U2g2Vc+AZRTSrk4o+QgBY6iJCx1o
RxJSM+NQ++/bSKvsWdPJhO8u2ETpP/UefpRufjM13DFwn/Kcdqx7ZNgc/mG2
ySN2hnARfVo/BLQyEskY04sZRBAOcnndcs6Z2lba7mnrdz8UKTGDFf6go8QQ
JAYQ/tAAzRQ+gZItLr6ET3Ts0im7oMJjLxPLtOlQUDs3alguie2TXORKPkxo
nTCpvB9Uc2FS/EdhuT1008M4r6Pua5V1j4ihUsgIIxQyKZNPgm9I6yCIonUC
pjbIAhqjQtjxcdOuNN9gs3BpTrOx/r6458AbK6xDgKrCOzJzvKh1+G1eWIy2
uQh4MYQDXMuA0U/ueqGQR39kMMpQtmVn2UOnDNb6rQ6shWF6nsYRdR8mVKVS
6ykw68Ag/ohzJaretoO4fiuZiqgtT7H3SEFlNsCe4X/hn3XA0FC7CbJvmHf8
xlbkVnL7ncEvI0iYkJe3rIqgYISqmT0d8q+CBP+Bl3RudwxNz3BAS48eFiQ8
OFubSe2aFSAquQ9hfx/KGFwMWk7uR1ziR/spQ5tTsBed+IsW+A9V/5iS2eWp
wGw+dyelIstggv7MQAJ4KLZUY/+sBAEXN1s6uOLbLvIC11Y8sj5oaDLyZsW8
Zt+4hKkANHExH6ZatYfpStFYiDiWijzCJIP6rb+8uZVgbHbYOq8lnM2J2Fp9
4QHv7F1utsZ8j5zLK3Br8LAYm6xWQQQjZv/gAco6KfgKSLejdydsR/BfiofP
i6abTxVIyf0oemqeWiR68k7Z1jd3Bn1o4mhkn10WgbM2DFABmOiSvEjqEThU
gtyquP6mkn7MJZQewBoILiro/7GE4C7xxy5+2HGqTjSC9+pFOkAvYoh0yNIY
TwQDbI8jj0pF7vCxFWb8nEiPqO6+GvaNFoMOBcan3qQA07tr70iUhe0VUw6P
RXA/5qq0/x0qb9rirh2C3Xm0Q18t7YkWd7CPe2Dv4u3ygpMvBWGfGqRSV1e7
j6kP6+b7/2o1fMofPF+2ULKwFrdRZkofXkn7213Oo4EEfL9CeqL12SJ78SkH
errHuXqBq/r/kLenK03B6a1dFfbUiMIxApX3BqEBZW5TiEcGeVznPZZMPEIv
qLA1+rf2Vu++qr+6SzOyVp+fZZP1vvy07XYLiKxvCQEUQ8Cd4aPhyBFSDPHY
dx01xXuRVkwofZkD+aZMaTNqLZYGAbU5M3sbgm/jZZS4iRi+nkaRc5/scuqE
yZ7LwdpE+lPogR0CN75PVXT4G1UfxmzTnjRNlOv+6DK+W+Z/JGAxmozdemKn
CAjOh+7qGvOE9k8kP4dIBwvhp8fHUFvmkVm0ajfU7zYtb1SKg1WqV/zmgBfM
pppbZJ/rBQuabnOl9GPDIc6cTKacgpdx0jj1PaEATAld6sKHie2J202asms2
o1IfgA1WuAShZb/IGS/DBJv3+6DgKhy/S4XL79NcyccASDRRFG+u+DLQDj82
kQ1taTdG4nItpWEaAjK9WrMZHe09zkUpTVHz1Voda29Q6s4fzNNJptT8E8Li
h8BC6M7o4aWLCbdmqob0BEhdAb79eCekgbSNVEvObT0RiX8BcmGP0XMqE+gn
h4XzEqWUfK650PoWDvWMLj9s88K39JR0w+UDPktlGVA/d0Rm8CU+c74gmXos
yAx8X3nYk1x3may2gRSOgEr1Z201yFSTr2x0ajpv6uJCNid9LFZiPg66xahN
0gb5nykAcBERDHj9sdx8kbVh8F6V65j5Va0YdwrBKy2BijgbkCN50oVMA2s9
7WGU8ZAJqo+dj3WqnlyF7CX+ghMCluEFfv1kYPZv2t5V2s9o587XLvwFM1SN
p1Z4PJqQHbFLsAowL9+vtES4wnk4hBDuGbwP0AL8v/F8KDeeeluGtTpjn03O
5iPQDaRPTa77EetIopEMGGEdHQ6UDXkjMoiYu1OOD27M8I6x8GB8eUlfJo0A
RfrQTnM7F1dtzQk/t7CnoTLIsH8fb4GNLi3aI2O7bor77GXbChkL9ji0ySwg
XoJmRcqSz+TzZz3gOHPb9gXmgcSI0gjsp+s0rv/QJUvpR4W8sdBZj/HQuUsi
nq8Ick8x/eb3fuocwvRXCZ4WoQvKIsNdhOgA6lTOP5Ncnocvw1JAUN8zX4ML
socgc1SArKNmkIzN73V7jYZ0ejPqm35qj7xINsYk+oTOyFecpTQfjAUIoX4L
3fs4QpnCu52qPivFC+Ty363WcceQBnsgqf6NLddX4C8su3xjsBrS5D8vLdip
c+rxWG3VUejvUnXgkOPpZNesijq0V9kjWHoYOhD8zB6aTdeOBLC9MkR16mWB
QkephC9QO4a9rr+pjQg1TXS1K9BafYjlHcTCcRFc+ClsU65dMQQ91ifu3mf7
5r/7zEEW4bLqT/wgPjfdMRQ5tf0SsjGCyfSEa0snT2SJUGKT9Xw3WeA1Jpky
O4MQ4vjWzds4Eos7+8VJTf31oh/17ayL/HNbvmNxvO9vaEWud4YN0+L/9TqC
oibWLuyVRdYsa/ZA/nqeorP4YIwqOhmuuZVsxQbBHfUNVxQjbPo8M/ZgdhEc
MTr4KKTepy4rAxYHFm9P2nb1GvXPMKi3fU5904drQ5uroTVOow46DJah0iPW
Qd1XJqLCGRlUITq3Q+XkpKgJfRTsKghWGc7PLPrRqXrA0ThBe/1AqFAEF96G
pbWoNmpSliEfnNaJGn7cXdDDvab3J7N/SS8HUBLYja2W5JD+OGY1vRS2dhHN
KC3foZNEB7sTbNYG95i5shi6RaMkxxDOpfnPYJXQpq5Zk6KqAyJ1OAwS81DK
Z1jCd/KUAdVfGFsi1gyxqOvnCURt0LYdOC+qOqryoPkPyHgIc+rgdDtSC5UV
f/nvbWb8l4uGN5Qw0RyMB+LTBQWq0+ocYetGe9OpgCgBSqZpjWvdf1IWDQ5t
I7bhdx3Lc8msNtLgubfqyPcaGVZDA/yqiALPQjcI55y5pcTMR6+3xtG9d+UO
fR5W7dw17OdxIkJZL+fezfTQFDZqrx2hc9N7jnvkYZAEbvvxDgIn4o22j34H
BRsjOTdhNBOLFCCLfv9Ql2sjkvlj6l3dgoJ19ZkXXh8KCkW3QzoxC+Dh+1V8
s8gSHRc0OYSre9dvGsjHOhVhtmb9UEcHknCv9FctVwBn1kLEwqY5/h1MeNDk
AzJlrCDnQjQO7ybKvf1gHUbeqNNki3qS+BdZDjlqWcL30mwi3XuZwVMENJ2D
zOb55SEpia4fMxR3Etk4LoLPhQ0iTQV51xjbvF8jJq9GNlnElWeeiEoPYpvD
Xhr7qXMPCXnhsuZgCgJsQCe0gYSkGZrA25qDQCx3l2tMM0qbzVVzHfO+2Vdw
AjGRPfBh+i6rMNHrVTHAHz757F3zN08BMnvWMz5icO4iTWOKamZ/viGM8BM8
lMgcTP1DT5DTdRUgyk08pQj596aI46pwFxRwJ5llM+WyN1FcIZfNgcGlMNtZ
USHbzG9dFS+aNepFGJSurZ9PRWuct+I1P3UFZMrtKmB9vK7BaN/aihIcV8m4
RbDJKFZyp6d3becdxV5DGioIPmO9Yvo1Zdlfbztx4LqgFiNuxSvgU4BovTZU
g44WL/LUW4Xkty5lww1P09wQpJDquUCiRqxSFBXS4sobwB7k7/erMI5yaswa
TdkZYpnTCkuy0K/4WJEKNCAyEXqfZWxNr4FOfTBfUKrdnIp+3qAECh8ewfET
EluuXmPFg1X5H6T0vUp4RRa95Oo5Lb4LHdOOwBX2mjmw5RotaB2kVexZ/cpo
p4pMEo3+LFepymr2/kL9k5HwzmsnvGQ3gSQJShjRDxlFbzjrHyLHit5Fd5HX
9mmNjy7/Qm7JC5HRYxK4SFT+0cS812T+BAPgjGU4G89VsIPMD9BvDQ+CZtiQ
2Hq5mCHU+tiYdiU31gQoAQWYzhibyIMDyewJQZeEcd3Pcrha1cb18L/sTs3k
/KsPOFNPFTm5zWoVxbmJ+pLLn+H3zyiTRUvTNuctq4vg3lXGS1wjsntMl4tW
wY9X7hwdL6Np5VRmoHgdEo3bA+RJ+w4Ya13cS8COIVyxe+RckIk1yNu2jSMt
vNLe3QDvDoPj8lw8SN6tUR2Fj909ixVlpezhCfdqMUBmphvrI6jNydTRLfiY
bU86QGYZTnzcahKopo8uLrIe4Xxltjk3Kdm4eu9NudhDdPh2j9ffyTdEusfU
t7TBVhbmJooTE3r8ERO2nxd1FvtvvqL4baAFw/IscfhNtnK/Ontd4vPTXdEd
ZjKnsarf+tbrm+DyjrUK16bmFwIoa202A10+jTbxLZq/INlRi6QJGeKVtJfP
XR5GVkKcrNsTaIQs68nQhuq2gGVAVT2b/sgJfMQN8lS0gAFwMDzF970JgoTB
NXfzsXkGfvX5Amx9i8zbClAWovW7vIYzq3Nv+5DmydTGKxM0nnbOxJ0Y/Wx7
c42H0Cu0dYdJOxR4fkk1KUV+MX0Ed5GczVIyBAXF9ecZxV3lofqzU6CGkKvM
plptKgkuhPTK2fKimNitlzReoTcLutUop5uNfWHCaH8BVaR2Z+AwnthAtcfl
onN2FZ1WEq6DpLjegJie+XmoDFL4VdwXTB1Wkm8xjS3cfUjFg9Jc1vQwUJDC
Sa785avOIar7zhPk/xsJBJKTrBUTN57QIpuPF8gDFNQ9tZ79zo+Ex/2sDvPh
Ddd70y6UoizJ7L6B3Rhrl9sfvn5J8P6d+7oSbOy0mRY42CaYDxGIxVzMNefY
IWQ9R/xqmeB23+b6xHSp4KTs/++AkZQUSuvSjGrPSteozYE4K8tsQ5UqJYXT
8swFBNdSmfXvvLJH6QjO8McFTZKOC6k7GZT8IO1R/qRm3TTl69tA7qvPbMgd
Z8yhEd3SYoxejNG+ldnJQ/t77zdAdPcHMbajBNHotrDpRd1ri6vMq2+Es3EO
f9Qhh/a68LSHETBCHFltxpwCIaJ+lIsLwY0Xkvw1lu0dR4MXywZkJi6um2up
p2nxPqPpzhrHtychW1IQZwA6Oijfk7hlGqwbpyLFx98uO0/RBXozSS9a6336
yskS/YLGYve0jxDK0fYl7IjUzeeNGzJgniijZIA9DMsgOuYrwiZGh4nHQJA8
9mhrR9aignOeBjOLSWPNaC2TWGyigw5vPDCdW3X3Pq7nIgM+PhwgDrxggFLo
5zo+ZDZO6f3XktpWO2pjsjyI/DSfrNvy+J6UCijoYOGDAIDla/o0czZqIsa/
Ig+8El8nIsEN/glvPoWkl304rIbPT5ApKJdUQ3UQO1fbmFO+uHdvDiEqOd0e
WKb2BKM/2n43dSNp3JPSYnYDL/LJFxLDKqpJhmOIATLswvCCZVIBr80WVVF6
m7OpaRAS4JtijxJUSv1hCch/9errEh0q1IptgGRBQ12+2NqU8s+jA3ewV7Cs
bW75rvFf5iifYN6Yi27q0JAp4PND7W1StwjaAlgu0yM2JKf2zQnjywSN9cyb
AWB4vT00AH2POW+GfWfzDiAq5Xvf4W4VVlwISOUxVpsX1sLTVqp2ADrrCPv9
NfFTzvzVq8lkbRTW71kTYCl5rhe/zA5EfTxtJHCsr8/7e4T35A2Zi39v/vcc
UbhHCtW5sC6E/TWqj4a5o1TvN+F5AXEVUkY1RN0RmZyeexCtcdUv8yX2asyU
Cod4AQCOGngWeWlwp6oqWMTpeNNRo+NhGGeAlabjyTLK2gIObcdKE2ywkGpd
xU26mWzoQoemVDiGKR/V6VwTQoJKIR6EBvBdU/3iqQKawEVhifMEj8QC/hXk
oA1YtFmP0LAK4/X5quvGxHI+gc2mqSS5JGiNXzzmIRvpnnM2A9V0F1AI1j+p
lEe8Bc2QCVlAPitUQQn7mBuZU1/jKKnlMAhO1k+9ZLAD5mOERSMQZ1b1azub
IbBc7bKddIzAI9IHo9zPvvITUBzIzJ9wK8OyG1qiDSd8+wYHvZ2D0slzb4PS
g92t4XtOu7z02cdmXKZjwHxJ46GMvLzZjYT10ewUPy4UReMO0wE898zQbm2n
vSokAOA7qiTxI9dPmLkEZepfYK5XMgnTtnYL79pm+Pd3afN1zdSnVU1bbElc
JMguKAD6IP1puunMYJcoaejnQCHb2HFeSHT3d9c3mhdrV/2qGfnzXrI49c3s
oXcXOQWu4+usKHOvfatluhw/oLB6Rot8gcLFi1ynVBUIvHyHIxbtvDizKf/d
Aebc0pSr7UeSKoEOIirjNo0MLBA7yoOrvzWxtGlW3tzXkF4EL30Gs+UeQcpw
5CbUYRjYRWliKTiL89nUe92HwX32xwmtBCmnEQfhrH/tiuIUC2Ewse/m7HJk
1ZQKKKJY1uIx+CwTuwiY47//be2ivcOnTQhsuZduadwSRiOa6ORMQrzclXU9
BcB2tKnykut7qCXMDq2Tlr164YnCehoQc4Ws2wtKqUCZ6elsw2xKr0m85MxS
IhQwKpUgUBAeeah3J03LJGP2ghUiLInWGrn0LAKp3sB1oHxrld03HdT4iI4+
CZKW2oNVngVgx73NmPy0oiffmbXVEq7AUxXMyshapaSa+ugavqmGWQZmFBBd
pvN3cCC2Oiv0Qynx2q0hSuR/Uqpcek5KY1tERtIokx48VtYGB4TAHRZ9bfRg
BS8wisI4fwWWGj5uNPkF34aQamRmP1cpw830lbgrZIi03X/gqO7arMH5JKGI
iZmHkTJ3PlcR8tgzfq7Aj5twdKYBvAlaNLVUYVPC0v505wTFhYYLqSBPxQ6L
1EmNx0TCCKCi9y4RqRd1MM9m0EpMTGPbOv4Byt70rr6LfyImo1zqG/mA0zJC
+lRTcHX/U3SZunLMk1j67QBsxF3beGx8m7h8bTN36ieGQ4bPDau8TX2De0AF
QBeIgVUrzK2OemQ1fMI6IYOPGjvz6iev1GP6JBTH0wVvoOh/QpJwIcFVXWJq
IApgrTwiBgOlrrrlXDlgbhH/McjNcN1BvNX6d/NqwlYRKSiUidwbfLgI8lAG
fF+oYZ4Zwbn+leX1ottLQOg23OUgZ1WT/LErL6vv2vsGwe4p/GwSPIKJ811t
KTdlev5EensHr6kCsRFVBiWQwBFRF4WZ5gxSoVoa1CN9yjEwOk4kaJ8iB9NN
hdvhCgHJoINnWGc3WMiJU+036AVLtmv1LfceRnY45uTWzgc+4afvSU2ivugT
BFI8UxcgLzjXmR5YZMfQaDarXILmnHrNJ3/bsF/ySdr0N4m+LIIt3BgGhpwq
Bf9TZu2w7L1RpauLa6SwnlbeT+HROFBV6OgLYpcMqfPozWnH67bNBd/KKmtR
FpOjnojAon+qN/SADKJ4Klhqz817utRcT3j1etBSBfqSuyrePZD92r+NMsYh
c+eiCN2L1dvobg3iyJXEbdHdCJu/BjaoCQNPyLV7m0h6qfhMax3d9iAzn/LI
cUeGa3vymqjPvGE3Ul2oYwZ22z5ili7+Ne2mNvSsRZdaOmEmSOYUtUDdk8l8
QjBHD9KPdc/cmcc4wt6NdHGzSAvpjlJ/VFqDqwyHnQ40WlTkbl0GVT4TCnaj
7669AY33+8uJEQHklNAPC9ZlsjBzLT+Gwh53UUwhWL0QE/Z4e2QjIFskhODg
zFXqzVUq7nfHf+i4W49Uzbx9l9VDnVAYDD6XSRKDnrD7hhTzqlXj3PJCR+lG
lmWVWKuwjK3XvoX8ORi66Cr3KwzcA/kk4apd3FrGGUEYsB11XK5gfqDq3KVa
tI0+NaoyFToZIcbzjCzPkrNwcywz25HNLMDtruXZjAt6svCNAxl4t8AN5omu
cfymTEO0Ey94aAJlkeUKnmBXiA1q+MC9LweenHYTJluAnAPnhWIdYbat6o+N
sQRqjC5Ow1W1mqB8X1m5SPyxSN5GqKF8Rlog+Cli/eVOUPWwSJWv4wSX0tW0
Kw7Jo3tavWcqs+G66u2M3nZnenjhmLv68lbfI7ERtL3c8SvpMtdkEy9uhzsi
tbu6orOP5+RlJtWGfoDbzWAmioxBWT4FQ5HVFFEwDE0y5xNVrEkAZUmQI1Xs
As24bShxjAqkAtqKXQnaVqhNCxdaCW9DAGZN9rQz/RUqxhqSUtpO3eKy4ONG
t/d4svLRo66+crr11P8e9CfIy27Bamj1u6hWYeh7bKSJPBI6aF0vS55OzVgz
+ao2sD9tprz6g/+0D+3WQaFv0A0FY2JeW3VXaLCIX2A7eZWPnhE83OVbQ1u8
813LH0K/EINk0H6I82XQuxC0hcT0JDz5ewM/SLhMYaQARy8vh+vXu8sIFWeL
REnx4F1qrxXH2YWGwIYl6qhTH5uQUgR5WOfr+6FxjBekoN6rXJ6P3XKJpsfg
qJB2ep+XHSsLNPZiWeENYlbMLu2nGiP9h8vjdQHNWUbZGCJJEGwbVx7+Ruzr
jySkgIeiS2nFZLtj7wHAdn4iAYvtb8cvJPcgMKSaBGXu9/rZTFAEEfwMxA5c
rEAvDCB/GkOUsbFF5/mk2LqpVcxaMfWu1vimjMOkc4Ls7XrjTH/cR9UIuCk1
zWsG2hTQ2RmGJmGaQlohWm+A53HKyUNEFfA7uxtcxEjvkW9CFcUa3gNuD/uH
VIHwtmfsdd0BFDffV+cT0TgraWlCVWB//VANeJ/NRpXBA/ZC4mNutl0prywA
BG3eKK21S9ih2N4VX6di/crlTerileFf9gJ0dMonIeBwBi3Pgd3Thyr/4UlC
g3rdi2O425djJureRpISV/vN4ssvp0UCxwjfmdoeCgEvNoqDU8kWKi891q3F
2zPPam3zAMvgZSO811or4CvpOBWY+5ErxGXl+dZxbB4VS0oemtQ90xhyBob1
1gYQjywHPINTxnzBu10o0Y3IYvhXhSaQFQjgOQDcu2MGc2aS+SsGKtFfEdtL
5oFHzqObhmkfHQvmpQaOgMapizF3RvYMUmvInJozK/NcvXIEs1OUo3owmiN/
zugugl2RqzYvpKtW0DjPVtbrpO/OjeXCZXGehxRkDI/BMu8cFMkeGrtbdst9
0x9j8wuszjSjmgQ/CXl+4gywHagTj1LVK52Le5VZPLTAYTe7GXsSeSg6WqWg
HdQhGSN2QkswtdhPQJoR3X5Ok+nO1VlkRt/hvU3jdPqx50f2JSWZhrPF+QSA
qQNXntX04qdFNLrWz3TqzlYFFYk220QHnc6RsKmbbMnFpnTZpFbFj9scYxbY
eawNyHvsLvzqMo9yfenDBGI+ymYwRJb0BRIj8L9m66Wu8fb2CgqXDrN38y9o
P2S1wLAnE/5bvQ3hHFej4DYhu6Hn7PuHQaaZPKmDF1NTmJ+ABkSx2tnnLxjI
/frMOKZGY3g9F2i219AIp8Cp8yb5c95sWUIwIi666+1u/JmkoQPimG4OeZCp
0SSTsci4N8LTLKAvAdRCx5pBaocOyHfFl75CfvoTUZ3tGRVUMGwNp2vEsrbb
JdN/0cVhZg1Ive8eJF3MMVy4saUpZ5svstDjmVUK72Rw9aoYhBe7S5JXbl2h
crsu+NNXGTJCAZ8bfgKI0wbh+ufdt5A6Od2974K7+vHSV4JZIEmhXBDZOLgn
3/FyyS1A8ViXhJhmt9quNwhSLvcFMVeMNRWbf0nsUpxJUAMRszbftf4BoxM5
LnXy8tuPGtAULrfXiMA0GBBa0hsaygIpOrySytcu7MGqIYz7t12JrfuRXm7M
GJnJjyaXLkDFrNTnlpH4TAWqftoezuh5O9UB8yo1cysbfBpmt8be2wuCC4Se
HeJuPTLWWrfS+3e91LSPWMlPXVFCOPx6HHJOPNHKIywO1TL0Y4w7UooBH94p
9YbkSmSeUsJanXx2Qe0q+/I9QtIFUhpL7GUrbAldmGdS6a9lvWDsxTlQ7ngb
NUgw2LisK0GlEn/8vn0Y0LYfayXXXe5ZY2Q+7mYZ1Ihy72PBSV9Z2MQYyUtY
aq/FpnBDAz2CNQk7NYQJehbimKcr2EzJjzpcN7bHVG9YY3c+BZwB5OrrsbQb
hr36soyNUSfVuZaR44G8JjtXlaafGNPGtRfIVA00emo3fIIxdpcMlgCcvM9Q
/n4bm9ywiSjQLZsmuEK/Od4bPaKRm0+rvFDURNB0glKgyJxzFvYI8r57+0u0
7X5m49xIsbiiEUC/z3w5qeXREsL0cARQrv22I/rCRb5ko18ftMsX/cltx1Q0
A7qLSHrT2u8nfnTNd/D4QudHxxmsqMXPCiA+qdQnb+NOMMAnh1bKUo++bo1x
vEKfHkpHf6B/Pmr1J3RnzsAwP4zsRsq40IIqMDU6XURlbmZ2tBHH6EWprZHZ
3REAXwaqJN9FjTE9E8292a98kLkGn6TNoy87DluKx5bvs8TAZlQLY6u/l2nZ
QFEzalujpHr+1lRAGzmxlIovIzfbWfYoX+gp2kkQjy55MgVXrX2b7rpru9Sq
sg/XnpmlFBwv5df6Nx+6zU8XxXloijzD7we7GRX/EoigDrW7hqztyy9FE3xP
+TPaSVwuDSOqGtc8xBPOy2vcLpMgIV2KEEPPeWsCkY+yGZCQQLxa+/OBgfim
0B9YmmIDvLcTMYPsT6Tb/B80k7bxVMeRGijB58B5PWHXR1N1voaSRTMUuNjZ
r8YGuNXSN8oiKmqJ8F8i5O9RXJWewbraR3/J3kZOMhRNNFSPF/U5Ur5Z7yF5
CbUTJqP+zRLmDaqR9jNsxyvLRsO4D9Fz7x6dTCZxacwJ7ZpOoWwXUUJpLaB5
Y4ZtQTfEGh59YDuGV6tZqNt157HoLScuJERMlevvpqd6qOPP6WxnZQQ/ZouG
rDl2zGDvDMTZHxwfEZx6PAQVs9rarMQbNhjFRlNmWbIdib172txbvWEZU84h
sHEx5aJxjy3UvJegJlZeCJSedxWkqE+jyBEZxx1FSEugEyfxJg4nTrNsiW9A
W6O6G80RPIbQynAF9ptlY8eimZ9FrexwfUHID7d499vo5h89CiVx8io9e6P+
hL0zf5v8M5fRvzu7K0gZqePBghvXU20XvhcDIiazPSzq60PAZS+DUFdv3E4k
JJdephpoUx9OwPH6p4buDtFUFWzZv9bluQMMLVmz8Av8pGn0wOLxMZJeYKHc
IzroYfGmHwygqbPdn3GL3kzge9j+XThqGm9ZlCm7FCnemI2NPJIjF2h/8ADN
0FeWURjNc3v7lMB70/NnebwwAPnOij3sdbCYeleVjO6g0C7ffT4ZZG5tAhFI
VtcMMB90oGAFn7poUJhZ1RHqBqc+o4qYqhCLoX6b5K5gYUA5g+uPwpwwEz56
b06g7shU9V0QEqAYfN5pgdgOzN1rrdTl59v3N/SSB3khpCZuyv/rR7rcCJhU
hTZPrsCqnF6QAlgFysgEG7VqOFalhApkO5Q3r42T3lBhzMNxX8JILXSBVh8y
UMq8mo7srNxrDkTL/nOj0sAcTJQCql45pwODvguwak/nDIkTCDF52i+7K+8j
s1c5yKZLfVOEG8IC2XQyiNL9hzNn3XgGVlsgxS/wn82IYJovRA382C1qQTWx
7VzfXO6ynyB4cLvBpgrY6Zu6avomE8MCfa7CLUzkzXAK+Gr+S20O/Cq8IljG
yhQwOn3nTEz3z+GPW5VMksy7Q+lCvk1xBHH6FAiSrUBUEqkbTALArXrOFHrI
+3Qb3H/Eryu389WZbGu/81iKXyzxtziVK5o0fZg9OiDHt4S8EggewQVZtkPj
m87LgwpZN+fpUMdz4TvAZzvKb6AXC68+calHpvzF0xzYLLkEXQo64Nlq5IXQ
46GEfwVNNj/cQdE5+UTv7hXOwiUmMkETbuRmyQpIEoWm2E1fb5AIKXvu9kXi
Gi+vnyVB01PgULdVBpaJS8ok2yjseXgt3Bun/Re/J63bSFD85uIWepDR44nP
uhJ+nmF0sIfkV0YYjcB/aU6HjTePrS0WHKBnUcPtb/paKaB5sXkg9j6PvGhi
uczklWu/y6vwzs+UYldFIi5tBUZud5G+Y55ejMGWqMbCkH5Q79WuULfpKN84
dz2hRiQNz9cfsmgixTYtrNBx/EH1V1XMrevQwHzR0PRqkuFbPhT+wm6m3l7J
Xsp+VaQsoYMbbhX4BAX+qfAVivVtznzK/mk+97JfwIJtdP55ZGcA2fIrHPWn
3fvttRUasXNhwDTuOIIF58IbexjEB/rDpDXSbEXfxerzlXsNnrpEqmywDwWS
hsYTWH3t6IDMhnb/ag6n8bPOmVUAQ4bOjyZd20QG+3YJaujyf62qdSyC7P/L
vaKOjGY8s7Ex9uU5RQhOrAzIx0FwIpjN3Zbe/1dKozbVVJYCyACZ4TwR4AkR
xmNRcwQ5Njcumhi3gbXdJj3Vr6QqyImQmNLI3TfHugPfQArQmSZQ8m954iI1
LquY2+1+A8c6Zt/sXmveDacwKH48H5ybmxPEPtTjXmkhBwpSTTjjtsYuMzNm
/XffJIDXm8zerTu/C4mMLKtryGsYm2FwKlEJNuq63ZHvoJBbAF5nEX3CY9J6
hOX14XT32T8rl2kcUq0N8WXlMauBc+x85ExXeMsHpPSLz6qUtSpQqgwKxHvO
LdGZLJht4VqONMgrIVNp66ZIpwr/iG3g4vjTb4Rs7A4bkblB/ZcxHJXNciR/
rfF9Vy7NsjWL+pj//dy7sTQpfNHwC31NbnZh4qaG7VuBqYcIjPir2TiqoWa8
1SwddFtFo/GisZAHX5VwaEWFc7EvhH67AgVCNMFy3L58hQb4kzAfmNREpyjR
xuKCkl341DkEVbbrPprYd3v56k37qZut4eOb2CzU/OTDtFig4UEjHHTcvXxU
MXlK3L3ttEDkE5Wh+9mQOiVFXKfLM9e2W7lW3kt8RyI/+tSTaNowuXeEf/f8
ijLrQVlawHURswhn8w47xZSdrh1HlbKa4I4rY+xacwgCbk7zP6ut8qQzrjsL
faT5sQESgok/oI07NDv3/yL4QHgIGt5H/jxqn1ettIkaasHDXI5Xj1HeSV2g
U/X3FD9B+YCWwFYO1ZIZ75XcceiBl1sUUv7hyWMeY8bTZJjS8BDxhO4iY0XV
B4k+1mU+/EBvw44XuVMyerQZNxY7vXfq6ccQnxTJjd7Ww5j7kPxQb3uApkhs
izc6vhqWwlGq7/ptXBbGFRF79zN5FlcFwEgPazoHqwU68r/vBFs+LhhAFCdP
uLoegqLq7PJhJbr2QY5JZ/PXBK+swwOdiBZV1WPcvtgnldhQKv9bhgWfaq3u
QU5D1oYV0hZ+xwOaZg2LdxXVDfmP/ppgFGaJtCYt3J38F4qOqhAl6/X5M5uh
0JTW1bYU2TzaBjrUH1Fr0/DFDpNk+ndI/uJIoXzt1DlooMYdgyj6kPoiWW5p
qgSO+VbMaSABpOGv3N8Lq+CYu3uqRvOxRiARm7gsQsKWtEDmi29VsBhxdRsc
5yd6BDeE0x0kab9BNp59VT0l8yPZvbu9kvzjlgiIsrTNW3vR0hGKEuaFC35P
YjMjljP+dyJwjP0a4FdPf0GVrWOX7TQ7/0+qKO9E0P1DTMLqNIxR1C8kr2mE
i8xT69u87JFeyrg3t8QLgsbFVsNPuOgYnbDKboI6T8dJOSlCXg74mM9bCXw8
RdKuTFoyEwjgoyjNUpsH2HjG1ks//5UYjkt4subvyJoURLBpubQTh7mfvSR5
twbezH1xaYi0UUtWuGuVZKLPNpEBt/1G7JYvz1WoSmuIZxT5grKwpAV2OWdJ
yKAiReDPAJPRzsSaLcRDLsCci3wvcBT52QlYCgihO0SQ0coXBaUUFooHEQrF
qkJxBj8ohGRpSzxsf4RWoY8aIR9R7SHs3TB8stdNzVdEMYk=

`pragma protect end_protected
