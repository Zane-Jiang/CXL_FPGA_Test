// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
rOnRLNW6wLCyNWJmkRQKdun3qJByVjzcTr1YFGdGHnf5wEAk5BKj8+yR3ATx6xon
UACXaX375OOCsT1oV2wXVg6YIkUHiqB9fJK+SgxKThDV42kZF1MZfHqCAcR6BJwh
eSKAEttuULZnGCoq+a9VzRyviI43GIFV2bz5L4+CKLY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 29360 )
`pragma protect data_block
xv9xQuK7fWbdNueHuT8RwsDFu1nkeqWm8HmljZOY4fGos5tBc7wQ97EJrZONprZ3
6Te0t6nbuFSRhE0rPfGYDR6+EtfNn5s+MTSnlX1PC9Ur0FTkWS9nzR2jBd87SLhH
K13AMLwjahtXJS5BOkCTOHagcEzkg+dARwKBnxqsrYrj2bF9GyBTVm4T7UZ95bv/
a507xX9WlKNyWKK4SPjp0gdaSRTetgimu3L0xK7JEygC2xdPjzuBuacKAZrQoVrl
Ax4wBy0ELyKTqTMOx7k1YE1Sc7Y2neVLOS66DiAdOE24zA5aV6QRMSEF748QQ6i9
Y0ahYPmz8GhuAx+5PFqaf3rX+ajSn4ZKAbq5Lt5qjQHhHOn+7hP/r/3IT2SaoX0h
cQZh/vpo+zF43O0vbqV8VWJJXDIQyE4EzciXB5hoSPvDsiAWSIEOuIJgxHARNrbK
tSfKcoa1Ux3P2rGpSRNKMXwLdWyMdXoyBXMyaBE9SVvVEg6E5SrK1tgP5TGNDK9L
KpYOS7e5abr88mBEu7tXjkMQGrsjBEm3gKbaa4Gk6Fi9V3QJkZyXXU0NjQBh8JQj
9f8VwHAP7apRMD2eRjyUI5VG3QSHzZ6DGvYhI5W8QH8+1CthhjpgQt6scJHUgp0I
xlnOGXcAmQ5Y0MO//BLJZ5d/H1ZMfaOQUdvrvuanqx52byo6Cv9zPuX9rDaYANDd
Sykk9Z3nX5qsNM/8SUxzEyIfLB4Js5Qr4Vf+uGnf7d5as8lda64zlotvMLo16Ksh
CHIVhRCEACZWxEMrFbMzO6QTyLbsLqIZF3sGn7IFDKk4+NM1MdTiw7y00ycgOMnp
jvJRFSYLN5B2Ya1AUprGa6cwO3DrR0opuggWlr4iVzdkkHJLTQLAvNlbCfm0yq1k
f3fQrlJa1ctDqceVtyNpqQ1wUEmSc8cDQO+HEv2hx2yzuAhzSApyQqKTSvzqSZXg
Wku/T0BxmxK3PUdSp+qg9gMiyXc3GRvzzptlamyhuILqv6LEBD83MS0g2+kjU2l+
9YXU5+bVC/Apn26pt7FI+HeEldOiUFqhbmLv36PxLU6DTsfRw04tC/rC5Qs6SMCp
eBtB6gKZukT0pL3qnjPG7D5SMBwQ0gTM8DAuDwEknYXQqyzfLyTXjRCJd1m2fAD+
Wnt//1IIydk1bNgoTRWeZZmvbCLdEDWdPXXdMoAkqfsbnVBKTGS4/odmJAHG91pm
ZmisDw9wjRYlrcypNr8nImfkBCQcAMWckoe6d4WLf3FzrEOr+yy5jewxLHKQBUAP
OimCMbqHDGwm9k0Lg1qGW8sD5G6CdtI403XwlT95/980fZk3i1SU8YWks5paowjp
B+KbCZluvCGQERt3/AZgA9eG63DkDDyMpG+M3RENVjZXn3/uO3VbFaPx+AMLvNSQ
b6TYnUxSfkfefk3lNO4iBzjVnC8uCYtNXgTrkjw8ROwBt3GrcJUwZXaZidibryju
bVeJWJKdpLUov3iqpZagvb2qLNQ2bIXAEZ7LHCAHCTd3zFnbZ+WyrbEZxLBVbDJI
HR9M7gAxh0BAo97n8V5hFhFyK0epKCx6OZbNKVjTs8vh9ma5cxPeYZn4K+9eGjhn
p39a6Fax9HOAeLDnOmFKkkykXVWICbYRPx7k/HFlDY4A/zDM3J7HIC1QJgDzkE7g
Q8GImKt6M1eJJdv3oNM3xS94l214ax1wQnMekxiUSP8A4chu6NdqN7WE1BOR7PNW
fVa9u1G4qoaehdCNjZMLpQB2ADFUeg83qbm+s4WVwWUZKlYUbq5rAbrnMrb/VZM9
D7uTLUp8BxTWGPzFf5O2bdKSUFZ3WCrRLFaRSxirVuVrbezJb536qVNjcKWB5ZEG
n+pLMgL6Q7aWuVH+SC1BMlpW/raGUH87RxQbdlvv029zHlFkmYCP6fiNeKml+cf5
WCryzS2E2EV/aFkLg/1lt/++WWB3yqOvwKKAbnJ1aWk4ES4zP/Qm4tK/IbBK1GVN
YlVTBkT82x5HWE4Ft4NfaJ2nLACBTkF8zhdMYsaXmdi1+ad5yLb8kHbOTmmfrPUf
f/SJQeZ1t05p2U9ds8wJoETDlWUKYbMMxxeRIErLgzcuuRi5yZNpeFmZyxK6xrJY
bQkbIX8KRkny0Bf9IUyTnNpaBeat3ZJOjtmUrAwiH+2gzgCYigW3FE58ZDZ3r7uM
zSuOrkr9yfB2AFNjOcBMDka96Wue9Vq/eAgTLwM+zmQkbdBtyToCTf9IbBshIpIG
q3cMhur2dp6KVrFZKq8dBGWLkIjnNqkcuprGKB9gQlHQhhKkUM9ekSkaIZVH6u69
W9qeSB3rr3GTTJ3xp4sSzPFBtLYWUE3BMaNQqzfBMkJb+3bbn1kJ58dNMQKo5JF7
4nwP/kSB4TC7EvbZ8Rs0n2lkuW3vqW8fdO56ECScadliyvo1RRvKwSuJ6yNSNLzp
waM0MElP/R/gVqb6G6PqhcWTeVXrI3agAJFCAngSBuBAVXnuop87qjJzLU7qPB2T
CefZ7M5TjOL0dHX5PqfPKVtpBblS23Z366rZlXkHiZPE61laZV9gRDW+DqZr3vVq
XGAlXRAekINNCUIxQFACdjuuckn6im7uMfZIOyDByzhPiqZA/pSlIYywLuqrr/3j
e+YQlsWsUK4Zgs283oToGXCsz9C9oRs/dGGgVgVs+ij/j5EeQAK+mNGBA6A2f07S
V+1/IicZuSHRw0HCT6VTyAv/BhKRfbo+s0KUXGtjOeu4w1WfY5kNN0G65S5thJGR
/wilQfNqPeWRFAKZ5X84A9cwtwhFZiLCbTuMMCG34+qHmvoFp5hP9YbMnh69H+Br
3nnjvkPkxvqXf1Tqb11vVTTqg2Cu2d3En+4V39dM8k5BmTPjuVzPHF5sVK95z8Z2
mjFdIRR0Ddpz/itfAP3RN2tdhdHNLUj7s80D49Lek6m0L+yBP5/+PIc26C2TWbmP
OBOIpKH16+oAfngNMMqKOkYFgu6abcqDQ30quytRb3zNBnj6jtY+US2OC8HxnKxn
d0yGldPjwiQNIy31pejzMQ9SrDZu5wsSGoCCXNYN5djs5fFDd5Mv/jukfEBcNCwB
qsgIocXPwkKGRt8LNdN7ONUBXD5L+T2vHVk98vA0H3ZyDUnRWueHCabjk8cj7kfX
ZMkJgkSkGshDji/ItT+Xggs4NX7wBBRBEMa9OJZCtyR+4wJYuaMKCxTo2Xx01Xcy
JAlzL79wiJVMm5fj9JuNV5J+seS1woFHkL5AAOCuBY66/grHCue2HS+DKzgjQeky
Nt6DUSSTXSws7ntbS8XRzJ9CPVp+lUKkYdryFdJs6xRCI435aMnz1I5uG2n7DLzm
Gx0U6mBpVSf9ymV08f2dKgXmCnbLRSpjgOicI+ojG6Szhe/hQsixfH/Nk4KfDbuf
mBqrI6qM7SSDd5p/fkv7E/9G4SixIs1NBfYEv+pSih/EG8Hj348nv/oaOSf/HxgO
PmfphB69f3z+wOCt/tSSGqooZbwCdP1YXkvI6XcfJ6GUkWASMiinXm4veEis2at8
Ct2FQfXCVIKxr4/HQaBpmOcAdnK9P6DvPGUbdGaaP1yjsyTTmeJGFw+SbuuBT22e
cPzo5LAO86oM+Q/7GDwaHVUme41fPFpD3f/c6zIbsZXk+xa6RI3VLFVA/fvyjFSO
dpCQQiW6lety752O5b0xkuvnI6Srb8N6mzSQkTL5AYwNgXBIJ+Sq6za/grqOi0ei
hM8IdoW8oUc2BKEll5O3msSDuFIWuvM+8JX4XOXtAGEgPJ9F5NZ9o5W44XVM6MTJ
kYJ2Xx5SfoAN4CPu93OI4gKAttsI5pZlGQK5ZDDvlbDbiRv6HZ3bQfbISAqN3ZKp
U5pQG/IXNF22moLv8Cla0K0aQWEhoy+Vf9P29MJdt5XW89UNlCUkq78K4hgIKGnN
zcq/m1/pjFaZvr5fnBRWukRU4xL4qKseAhEZIblFYBodYX0pOORgfeBOFOVmnwXs
bD0S4b8CYVzM9NTjbig6brgmW2rnUYnOcx2g7O0VG44glOcOctnci3ncyLiBCq66
ApJmlaVsMksvAFSJp6w0aP91RhNR9ipfnUn1f1jg4t8FFmNR/a7IqnoZUFcefqYj
vlmRfiFKWuDnkCwLd6nx7JcsXNrCA3itSRHPLYf3T2Kx+8U76DG9x/mnPAtWOYM5
kgHuZtGt26PV65gQPzJDxTjgiOT3DJY1IbBn0X3mRQQnwEr2PXJieSuTcKZ4ae7L
7EFzTNGU5cWFxV6DgUBgNPWeIpRfd57bqjCzrFON3rU4mZvfFDsVI6FcVBG4j6I7
di2ETTNs8pkIQ8MTkzW5U+LQEGy9OnD5mxlpvK/Uq9ZpqFhO5jcmV7od1l1cX2wU
KC7/uSnpGHrDXgewrkFzlA+UoybezT80pFwFWbvRsNPVmI9tS68fTid+hDqQRa2X
uVNR1gfM2c1rAteXSdZPOPxZjQcj7hYc0gHMltqSn2jlGW+0YYY1ZWbre5EQB9RN
zvmjDNiF5xQB/OUfxEYicN932W3e0FwjWKigrKxhcLBkHdxYZLB0jt7b68Pyx7TG
z4snszgrHzg/oluWJYdogFhiz6tByMYyF2dhH45Sduy4konpq8FbTjd0fPyUC6vv
ocmppT7LTTuV78zMm+MRLRmSbnlM95YCJVgZWK5+ullUotBS+PyabDvF58cc++yJ
lZKHl7TTLrztXIlz5WjQvBb1QXWzS/qDJfBlF2kiHMN1BvITZuDoFH1imYyE0jKP
2z5Y9xNWEsqfotSz7Kk7kIbP0EYo8JNaWLSNvAvg+7oujARto/Pnok8Q5btwJWSt
+xHk6IL773HB1yX1s1eZFMJk5xwHC3RIOxu+U2XgE9caa7lkbzsqkq5zlGMU0elv
fURArQ9qUgfz26RqL7Dv5T24N1h+lj6KZVqJNxjHh6nOeCham2ShivpXcpFQMp7h
NLQrN/Pz7iDIVCswRTFDRZ+hIvC+RL8axxOsXmU6cv8KJuJSNRssHT/jbVLNZCSA
FiF3yi6z59ObY362K4OdT9gkqoZd1XFr8srwZp/CIA12lCnM5xdIYhtaeBJagVeL
EmroBfWipFe7yOfoUZVmpNpL/PIWmIEq+iObiNmL25d+ocRfV0QepsQ3D6dm+wLk
6ZVVD72Nd1LN+dHl+Ooge5ItC2l/Y+z6bzx5BH8uZyONgjJt73/06cws5dVnAs9W
YEXvqlAUWh+tBOd+VF8TKzChw2eBJ84TOduZ2rX9IS+IjB7ZSi0SSspCJJQa7W10
awTguAJQZrKCOl35bK4pINJGxNQDn07LpG95dhG2MbupDmkaPndqAd11UHkDmmfn
Pd9QprW6Bbe/V1OZ+zvJvqQ21O68aaybQ+LTlaHFEagk5Rtj+z1MQt7QGzpRX2Eu
NL/VeeHgJOG7ewMkbUbQGoWNTNHGVFP6UmpYHIkAI/AYZJKr0n/W9eoo02UIsVqs
k5kaYrmR0ImRx3infzEIhjX0AnESHAlL+UhF0+pUO4Iu3bhNOuCFjQNsrmMI2Ti5
06pKuh+vQ5+dBQ92QhE0O1UpYyzrynSG5cHxhGHLFnR8xtaefxeL+abTTx4M7TvF
K7Fd8T9aaGriwgv4QYyV5Z6s3OmNaTCmW8kEZo9LGFPuY7nYQ2EVU7JqHHlfe5cw
r6jLVB3rEArBq4TkWJvAsJ4Hj5fmYLiGNCnHnxZTiQKGAmcX4p6lRhmranZnqI12
eIihDdWm2KWMG+9WRXulbwL3ECKTcsGsEjXGdc4/KY3sqVN8hGIOMWW4SfeCtOEL
BCjDO/FDXIr5P7k8DT27aiESkZt5ququn2uE0raTbAE54ouaI/fRv9IOu6s+mjsK
fmzH1ihCzu7Q1BBWYo7jhSoHKLK7XWkhxr92rWoPNjElCw90OAfzbAnQSkuzaq80
6Db3SIoSx5sNFSkzYZbxESz1/cgTB5TScXveBWfCyJ1vilz8Ni3eRWeFabWXtPYn
7D58Si/VXBn0b2jTX9dZIJeo4LAPOlkgE8xagcpatDX7GgpkNpT7hkeWDAtG6Iym
aSo14m0avo9cQjal1UArqToN3YImFwTXlw0RD4SY0CeWzPLhIknGIidZRH7jOse5
NMpCl7ApAF4MrwkmZ545MhRWGUNmWqT0hgaygA5Jgf5vAJXAk4a0vDLsbRTYRCca
graAUwb3+Leo8FbXkGyqXQQIHpf3TvEQkJ9++i684laQvwOrWFcHjiNs2ivtuqBK
YFM+XjkyyY/uoPx+ZHHKjVFWWBHBfAGz8t+ySjPx0ADZxSgslCehUzwtZ/iNTzD7
u6/doP6/hwCdv3F2r9snXvSE+EuD7918I+51Ft3o/pf27z77kalPh76n4AEQeKzg
BwQOAj18Urk4bKzM8CPwNcbUan+GuL8Dk+nxH3JDibI1N19TLK6yLlAWVO4gyY/o
I7gD8KLo0EJC0iw4w2IcFeGcBq5wWyUZkSPE3PMjD8KqMnfKmC0udSsAGFmo1W8U
yG0g8w97r3ThR5zCUnxO59uf8bYS4H7RtEfWELgDiu5pBLOTpGTKp58fQPMN8IjH
7IAEw/9IgxjfYTg3RHXfGDdidCvaf4ioKpHa3m4MmPQK1X6mapeBHLjpoq7jObyC
eHMVdj89V9Uutycu7LpRONlFrE166ZdiPI8QeeLCFCZJzP+61cEVcuUnwkZBEHOj
mA5RcKgTMfc9bcJI27MJjRK40ENCAUIBCwEt64iOvCCxpbQvTG8ZIhmyAZjL3BOb
cvpcvrx/Hznz1avWVk0jzwikIbON54y97GY/CLtEVD/IBarsjGXICR8CvY7XCIzF
guwpoX9PIB+a93nTrDDBiQDp2Ay7YSCeYtCPn/eT6R2W8gaN8fwnXXWMhkyYrnWo
tQTML7h/EKUtd958pGEo06vdZwcXOb2Ya3FMD8bFcjopqb06N2DIYirkxfmUfavS
QQGyB+/HQ1cZ3qOhQxqfirSJc+jE/IK7hT9dUq4Xxvk8idYTvosHEg6Xhke8z9xa
b/J0MgkqhBvbw27l8l8+xCwefErPvBBjL/gEKd0kinl0PedLAtp2DThH9G2JmXTM
1X9TBm3ZIyhU2nRMt5bFDnUzK/MLYO/TuaB6xOrG9I+37BaKgYGN6P4TYcwSrnT4
e4MCj9IMd/o01XiC3Sjg3iYFYKpMXwVFA5s909LREe6v7N6gndNNecv4bJdvgS/w
NffBeu8+G+2tVvkIVryiEgFG3SClnOpJCsumVbAMJ0cbLJRS3RoC7Y1pbdBJBgDd
lUzqo8rIX7/5GZ7LV0uZHbC3ywjPAPna+2wpz+6uYLJ5+OulimwrtxzXTDvlxTZx
xCU2oMkcpEpSsbrM6LE2VWnOpB0NKtfgMTXMlQorwVwguxgOmNc2AMMixn+JEjW2
GzVdNCLQJWehrzJi8tY4pCjaaHlnSdoM5XyA52ZVrjiTjmu1xoZwOUg55MEtVk+Q
g1SBxjOi3Um5xXarhpJcnOjaimRwkUCFkeCzDx3HgsmqSKhfRb5yOulj4bGQIQ1S
fahUjf0LzxZ8DB/rN2DAMQHIDuwvhb93PZ2WvpbJByQFQwXLBXW0LEL2nNaL2aV/
j0IS3dDwav1/MYIuRFipplpeO51opzx0Agl33R4HVmyKybDXltIJxDckKQAmLBXf
T7p604lpgumanLQS5GWk8XHFK0BHdyQ4jphgSQXJNjLvNG53X2AAyzWC0E14S/zM
jWRQqysFTMywtszdFZJPsgGygRBj2Gb4I6tf/i5Uw6Vv+mMxtEEzmRUS/bbyq3+u
ry4bmxShVhrcb2rmPn/nWdWAfZCtH5FIF4GR91msy6p85ziok/eFDyvek3gDT1te
m1O96Mgt/+SpLbQBZ0XvcP//9DUr6TuyY2ff4TNJjPqGdYZEJjsZ+xobkZIogWEv
jQrcbK93OKxBNhPvY24OHtAe1BiealMpbR9xa18aVBctR4fWuW6FrwTbtRDeMFl5
UdC8/a7jtvoy284K3rdQ5vT6hFdga0LQfcq0hULGbqsuOG+r19E3gdu1m87QaDa+
Kjb+Fe0MlUPuMo85BM27G8/K2p1NATXa0Lnu1isGF63TWJHOQYN/vsN30tFIYAyC
4T5/wg/Mt8+T2SNdWYDgtb07jrDBv8S/kxFaggPZ2cGZ8ccWDNIjjSDg3ykgFH9/
RYzTS44RyhcwY0iBpePdtwzH/0hpwahYqnwOWFrowztcVwgzGv0M61FrvYiW5Ud0
gCiDznjw1OZgBoTORAe+ew4is4wJQ6QvXFmOUv+NY0CNWDpSGJzhkHjjTAmbzfVr
Yg+ogzoCvgUmIgroyoxNdsbzWQKbI0lAfdJLTUsYQfn1SJh42I0RYRobMKMf+/Ob
82WYFnDYjZ7EpkD0qnq+dAiheGLcwpyuIRpUV/7cPx0Sspt5zS2vC7QiaXgRr/C8
/rx5Q75LZl5jjSGEnHkOhUB8FxO+7iYWoqbtg0y2DGOXy5SSEhGmZ/WnuwjjUuSK
KcOmomgiiR+/gqPNQtiUnmp58fxSB5z2N8oDMKs9/SdUNtCbnsH38fnKQkJg9b45
BQ9J9ICdO7sit5pVmD2uXfvrTTdsFpClzXW8yQmTPUHE6O7rN0tl5/er47CDNPTN
GXzU/2yt1ogp81gbVzjFMHq9OkAUsd0fm5TzZxdGab6cPLVgrVSULEVy2hI3syJc
BMI6GSqQll0dmRqEnjMYl5pFA534VTSgir0Nl4Vm5m/G1xMKzMxCeuNrKhh+ztVm
G8LbR/mvVTZUoe5hS5SELVV5jxEcLKe/tbz7sFFqtR67XKyygAipJy9VIDEYZ+8U
tcOn37ZXU7hKm1iOrT3G2+FzZGXdnhtwmLE46ogPhYWnoUkqoX6lYo+EiqQviZJX
IZmUfOyIqt+Vok6KRO9ufD5UQ5ZnC7LjMjPd4OXY1bijyNhcHg2kh+EqQ/gN6Cb/
dBkJ6Wu6aDY97LTwcPGsxNzs3IT5PBQrCJZPxvAOwNP/xBifwi10Fvkl/L3lKu5L
s2Xxv4L+8v+/IBZAn4UJe75USIf0AX1i2Zf/llLaepxWEL+wDuXOl15SybNIueGZ
qyJa+9pQlf/nMYWBzAqvgsL62JRqGG5VkACkjxBb20smhPgz/3EnZZ8D3XIHBdce
84GFNS65yOdhNjiwRKEbnFuGQQ+o423Tcfeu7VituLR72/N5vQrnOV8QmR8wtInx
YxeclT7nKrrMce3ryrBx0dOasp5O2HK5ZjbQyKehsfqLQajV6+uc89DKG+fnZsVa
kxK6fiWrg9J497qDaWl1JCMgrTYvVwcYk5IElBYzQHCoHvNPWNTeHw2xPkkunJk0
s1nz+Yv6exxiinYtTeMDBpgmQYml6kjLJFCGR6gdMJdz7V1+Dd5MsMU0u9TLRP/E
jSHrBv31Lwj0MeGTMSnOV1oFg/CDYh8B0ItRjMDJlk00ijBnCM9oqld7DDnnkZ9N
NdAM832eXWnkQCcMuOnx0ICSy3kK6SA8/nYPyVpO2odJrSbTsGv685cca7beT6Xk
hMCTC2BHFgZJI9Ey5JdE9DINIxsMocwuVIsnIDQJ/DO6hmqLU99uvkZvATT3SazC
qxcWNOjQ4uxEh6PWnYnbhLBOwjKY9h3c97hWkN3ScQKjqUFxu8rFnwCOGKCnt4GJ
DS+CWayrekGLBelx9QpzQhA81G3Bm1axRY0x9LUgfIJQpOe14TotR/bBiHvOr9SF
E1oJuxYXRRJvjhODFq3IbYqYMyIy9UMltnQEnfb/1GyzwiuiMRIqvaZhqe4AwcNr
IP1gLQ7pg6ex1sq5M781aHSm/FElZo8hG+dWmM/RVfxesVvGDw/u/FK+yy8LUuri
IDFLws6EEytGpgSZUMhNIF2rlfB2YK3fbiRCOzoSvEFcJ+kxq3Ok6jjNBbB+6C3S
4vsM2Xhyti+p/yMTHMtJjOorkNYkIqwAJZquJTbOnJYqow9wiha+bploDkCxzNR6
s0e4lNvwHRODJkC6JPy6PM+IYvsqfq7V8mVYqwwIP/4aK7hvtftx+CYTy7ESDjGe
saPd9urPMVqSBRaDqSHZuegVchJRBpsP022nz+H5a6k7DmkGeaghPDO+SQsRs8kP
QQvvJ3aKdl3B4jwihqgSukwCIyzJFdslDI/0eBIGmlMF7pDThQxEYPrHkJQXUw7i
4jqhsDB6c9gHY3nZsjJGqBkTqmLXRuihWRsqK+v7MRo02HLlaZ//VMgv8MPE+0Bm
ud73zNXRigGQi4r+cXyXHNcbosP0UcQO4hyiq8I3/3ln4+cb9c3GK4z+SYjoxCYe
1M1hpzyQhntWfeLtgF7U++lXHV/A08qMiWusIyX5AvOh+a61YtbXXib6Zb4hG/c9
hB7OMP0SVG9Swm6b/2HWaeev+nKmXmrCL/ggmCzhVcMeAAFJawLJQPt0BaA94vV1
oWQEBIwPEf5O/bnIkvAg/Efv0IoNY+vHzowakpvfFDNU3msopKKwsYBiDYilgvuA
wkH4rIrtgpCwckCYIKwXK+bAvUbfv5PyIp3k95rv6CKYoHcwmJ90WaZihHgUjF0/
xplw4LZ1WJK0N0p7hhyNr0JoQHUZLsv9sCSdvZdZ1zYGCinp9HUw+X8/hn/8HVMc
60KMWgrKoLnW7o/2QJUsyk6uVLK6keU7LemqBekE1QtUgg4nBaOCiHeD/RoZYh+a
s9PQRPu00ewyCl0G09X9qct7jn2/6OKIFgGSf9gLbV1Xdu73N624Bjy/y0chDVOd
oKbtYHYb56FFPxOMHxvclTfywuvH5OTwBmZCMDQ3kzjvgBXfkQ2sRYJNZZh65Osn
k6rnrOYjme7IgqSmr8Sp2NsYvzFB+uetD3M3RPz04/MNGOqmXSj9nMRXoe4zBYDw
6vsN45RFMruay6ag81+3BZJ6m7VBbekRXwRg1BzoWF2DfLdDeD30ZFTmnPZxGWUf
mfBaWWUkv8Oo1pmQ6YyHA+bVpJt9A3uX+yOOwlJ5nMCUjXaGjnhjp3yAz1cg3Lo0
3Cd8GWkXY6naMUbzQWsPY5Fw/ntzHI79CNXfvnt6OGoHfD57vFOp/GxtDru1EZ+3
tPejCtPn8Vrw8N+fNNswACxelBvQDLOzkqJBVRyBXBi3nhYZeqtFUiywFXK0VwP+
TU2kX+d6MQ5V4KMYeyGk1FOA21jn7EDrqNBUXUurisb1+pXThRs+QO/fgWcGO3VH
53uDBjV5r5HGYSvroJyDjo0Lh4zyMsu733BWy1vIqYs7KQMdSovHi7217Ry6wN5Q
SK6uhydv3tE5RUXtE23aBJvQNNW1m1c71hMgY4I0zdCTi7qEzWb8osykFoPunipM
xMA0YSE+KISPsszFGmog4i2l5T3KoKTmF50xXTiLj6xY0xpJzRD2gLUwhXkH82xN
JKq5Fo1jgxV3JjHGaQnxwbdVTRav4GrnaCAAh57Xfqys2vmFIV0r8009u6MhzhXk
5tgshgxz42FnUi+ZCSjQuvDO3pP3jVtAudNE94VFgYV0gkS9COOMzaWo1nUF5VRT
zEtPdBGXZiYgRSzqTngPqRDX/aRRKuXTPaOWXBgodZYYjsRZhyqwY5EIEh4UEYy8
oIMTOrqpnaI7Ji/DWBcz0TWQqPO1MTqJO1jRl+Q65bgjh6/ao2767njdDBtB+/RU
KIVQSlIPjO+cK8jTC+kXPWfTanEENUC389Fg7Hy4zePqaOXE3gOHw3dEdgSDTUX6
Q7Ty+xLsW9P1V6mzmiMdKWDbSIB8Hsa2cVUMgUbd8wPals63SQ28IrpfXB1K8VoH
KOHLwOSbC8DhEIKaM4DUghrFS331iTxw3lIoNEvntZImosBJJx1VVugZKUGc0Jjg
uyDfPF8ke8uQ/8kUdo/oLPM5vjEkMy+eoR00rqB2zvaGyycfqf97G33Tr9NA8mNf
FmqGUt2iUQPxboo87hxoyrfRZ5g2/7foi0ifciPnacdg6Y5eiOxAIWEpwXLenf0G
uo4qEpSu+DfuwvcWIRDShZwrrnUQB5yGxrVAFmrDpM3Fhc8+ogwRrSf9cpepuZab
HX1JT6/lZ/u1RChQYZ47Aq/dM6QoF6D7DB1SY/15ajKkA3BnrA1kT5a/lyTyDID+
z0wSyfyF1gljBT5R9770Mf93o1GkSeCmSxGr71qPZFUdK0IkgCxbkabL+DWXIT5d
OtRbIV5Ga+kBrzBMExUNCQvlbbPmKI/CguYeTUE0PM2eTMKfvYBgKmwoYNJF+Lky
EQ9HmHIRjznFwwFTMhNxSLEMXyj0cIY3p9I1SiLBERkh9DgOsvi0wvK1AbEA5NRE
FYxoyeNcOMksKPqEoHfNfZnDQEOnnO9NxZtPW0WtAM2aUiXGHGVpO0rNQ54hFE1x
qinvzQp9dTMq8Ht/tJZ/3ZwBYCkmz5e2BrwmY85QRnnjjW85tuYnhG/xIcdlGzia
nf4EGJsJ0rN0nlTLCJP4uGo0Uhvsyvr1GGsyCJlWbfUjEz06Sjac3G9eCYVJe6GD
ouvRVpJPp/V5Iztlbha/gBXqeLOcfi4S7oa6FCWM8l+thvFiqMDO6NOH8tUb6yi+
7gXVZtyuxTDbVfyQnpq5NepwGk44Ez0kXElN+z5mOz7u2sDID1rKp5443NNt5XmJ
MLFhZ7LgJRsTUQYGPnFYJ+VVTBK7EAuloO5DSfcUVNc6fSnZW0NGrdR1n2Nyt8jF
FC1ZCYW/6UvpOUwZd+VEcNrZMrNtitcwfKSkvWPUpXJPVEBPnU+1B2jgUegh7Aa1
qjmS6LblSI2OsggFRZk7hxrneEolpbeh/LIxwmnlu9XpNiiorpj4zHkg5/pVars6
yiLyvucSyZK9ey7x258Ko4eXkmh/K/wp4u6Pw8YuKDXxlIwuL/0/cibBWp8JFV8u
sP9WXqCdRBJGA2UL/5JfsMrYuCvrFbwPUs34OtYuGWYRCEQKsS+aPOG1rXEYtNUC
o0OgFtbYm8ckqvtY86kU4TP0dWYQZNoRbO4tG9+0yWDOlbsxNj4t+Xjxp+6lpSIw
AfCwnEX/6PlCgSnJs8IjA2KmPtn+EX6vbvO158Gxjy5eS2ZAzooAZ/e/Et3BdagJ
8BJ2nDjMw6AI9DhUY0tEV/NCrIr36bqlC6IHkDFb6wBbz7EhaRWULQ0nIr1yb1nO
kBAlmOnEw6XZJEcKk7C+RPQAie1vVoLEI9gDTjtxFRJpn7tzcTIwHu95RCrDNTWi
qnGgEzUcFuHWoxJoiOnwfMavcyD6qcGMTjE5sVyDVd+t723U34LnjrXuhEZXkoNW
UEbZYS2iQDn5qfKOvuu8KNuofX7bkgTqeMoyDklIAeatBXBgEV9WNJuS7yRJvxwv
a281US3vwBsQ3Dk9X81JCqHxnGZjjCacWdjTeBmvoFvYyCTyfFf87L+f/mxEaxr9
R23ef4/KyMfZ6wDDAtlJooBT8F0fpHb56wf9wzEOFQMaoFpUtXIXDZj3oIBLn8Ir
KS1rvhZyifcD8zD6Yj3rNdLmYlCVxhJmEJAJOZG9vbWUi8QyVa3A9ztzqCP3okV3
zNDbEmPeu3IwLui5RsOSrQX9gRHhMRQW14PXdMZ3r6qZgSw6QxS9ic45I2uSfjV+
hH+UePvK8snJagVUuTS1fe1na2NKh4/3aUPV75sa4gJJqeqE/Tgh/FERgPo3vKVH
7yHKdE5aKvstmg1pkgqyz6UzTWkLHStkrpeOJECWIN+fJ3HGNS8uNKK/ypjSYl6f
5N+zkOXrWawh0VXTTDbo/NYT34nAUy45ApBwsEoWhWFnM+FHaeOIJi6nQiaqYP/G
dEkgLUp9+mcKQpXWORrELHKKK3d6Jblf12kmNe7Bj9mLz1aVkDIVfhfLhDqgmnRN
79m4Rc7X2GXNV6T4mjbZIRaeMEvhZ6L7jkY/c4WL8EkHGplB0RbJUnqCzMdWyBj5
Almf2LclDPox4uS5buW5bZKLlp6DRtlRl6QQPM25yzqaOyhuRpcOuO64IayiNRF+
hlAZWokQiK+m6EbgjcOwYdSL95552FsvNjLxkMDB0VHQn9Gd+uoPTZxbW6nBSmnL
EpuULLQbz7lXGplvf3l9ljQfO0XjD5TLXZc8TKnil1a9RSvBb72wd7RNvz1cCW3T
LexZdDd2IkfZxYK4fZh1bbMWvD7JWCzW91APCCd+0MjEhUtrtitu4fy7UOUq0D0M
tau3oHV760R/Ng7FXPcTz35SAGL09aZp+57bfR8tWUGhFXtyIV1UScL5KAAdnmg1
GFO2w8SrToBz+FQZehnl3L2UzcAcYGL8yOazTIsW9dJpoHYduefWtZ7YfOIFpr84
QEQ/lHq+5Nfok0pQ+9SVLP5Zr6VNQQlEKXibIVZEvxrClE+VQ9nqCkGiP7MaRMD/
0kH/odkjJW6VUVhxdOFq2zDZN99Yqo5f1A2rHDow10n0nJ5QEdmeGQELT7td2dZZ
11bJJktdicIBsdrakCljeR5C69SpWfl8aI+F7EGel6zF4K/ZRoWauumB+N4jMYvc
xaV0VNHNu3a88JtTP9otoPYVb7lOy6O21OJ8MmcZbkToykaAxBmJ27Yg2/fzDMQT
Z+ipjF34qd0SO5xXO3iIwoHwWufr1PVSlsx7FiTs4QRe097E/b4tIL1jLiNn6rXT
ZvSDdwfN2AmpLDwnggLzRLB2/nZXEu5eif5siJOYQeH9BLnAcIszBfGMJiFlDDDA
KKwAyObcmcZ6JCAlMYpYtLsQRjEvA49/U9plnyTMnRkDWpJyKCyAcp3yZhU5yqV0
xhabhqIvsMjBNPo/0RlJhlX64+p6xImyai+sQkDG2L/1SzhvLfHP6Fdz8r9iCvX1
85J4g58Z8cLnsCHOxuEgn702D687XVYgh8oi+MV+lM/J5xdA4tBaIoHEOPvltzIj
dMMuUFhhwfFivnlPy2VEACfZ5iUAMj5nruxOdZbAHA8fhFkU2jt5ZBCPkdlX3Fko
gqGW3ygOtayVKAlWfGrz/OlC+K3Qme9daBLg/yNy/GKE6hPLe0MZDjxmEyQo3lrA
ROOypummcEVgLMLHMwB9K++1laLZtqGsqx91SGPaO/KhNk2JgGErfuKQtBD4F8K+
54DTY0utVaBu4f+6vWeuIfZSHsQa8vh7iTpmnXYLdaJ0ycpAI4XnkvEifNanEcMw
mHbsnRGdqe5DhYd+oEwthXhTzU4ulxzxalN2tTOGdgkyGMWL0dlXCtVGHcgDhw/l
UNQonEtBYlkogO+ubfKSa94lIsWeu3QLi5I/aihgtXKAKorETm06IhZr2zriCpgx
8VJBVvO8546TZ6A88xIa1rVsm0UBHq263NKrgitS6HTmsM1b66pHpp3yZOYXYqj5
Y1WSJy0crCtiUe3eozj0ymUwxKEMBqM0ywaZXbNGTuF0njQ8b/w1hKQgJLTO85NA
vIpG72oCHwcFnMaxZYhNg8EPhOwH1UD9scyRRf+tEZTOO1bds058seGlAfrKQFji
obbCal2orh7clRAog+vCfSpDdwmbsfjt31Wwn8PbZwfRWC4wOzhXrdUtJhi2j5us
F4emJHz3dhGljQI/PcS+a2J/loNJ1ze2cF5v8eJcb+HrSAP2e6MjRRQ/FxKy8fLr
2/LC0PLVqW612nAEzIt3d6b29h1dQuz7PqSfGPwDWqnQHMfwneWIzKyalO5uF/NC
26Z28FWjWJ2BGM7Od++oZIfuTQLETyhYHkEF9PsZ3WbummmyE/16q7RBrASVkRAY
WD7WwI2JI6NQ1JZDg1WwXHbBdbRBO2OVMkooZmcOnfkZdD1xAuTigjUkdPjJOqjT
/MAi/J/XGlM6VjwtDE4uZh5Mag4N8vQpPr5VXwAfSpygt9f3uImP/pQcaX2eSeC2
KtHdDveQLAMjZHLZK2qMrOUlWNJRiYxtuyFuBy4E2XmliknLVBLAMCc4Mq0TMzGB
9q5MdZml546tUHG08ivYtRlcW5L2V65Z5zxMv4IHDlNsX0eD0NDENCIpIzaQ2BJt
MI2KuUWiyuslieyOISVqJ0Ff2g6SNuAMpBGrIPkYwVgR4l3Cy6pB0kEeV8sew9te
l/7JMTCJTqq6MoVvxtkwdkjLouc+FWevsK4y49li2vgmvt2WJFKSWHYKCBUquB4q
c7RuKAu21F0iBTHDJGdARYqx5lLuQQ28ccqYTyKC3osqQqmdO55BsnMqDc7tH+DQ
c/qy9L7Dtq2gBOuXLQ6QNgaog1IrnahMVX2dTzgbJCE6cPmj5+2ZOgwpfLAGkf+H
bvz0uJXopZODG+mmwL+JsBiLhWJNEJBC1CG73SKm1ZzI0s3K6UEWjWeBby4RiVbG
TcDsK5XD/kaJ1yiLzhboZygEnvYpYZMnQzXOq0BHBU02Jvn2d1aUC+1VEbuh/4B2
/LcohhHwEwZmDDJxuwZaB0gqtpEI/Ofa9byLMHw3CwuDN/oWKNlKPmb8ZqMxd+vy
MU7frka/ggl6Oml9PzQ1oBrKGGDng7XoUoUH808cf2Lmm4oHEJuZe700TGiDgjhE
K53uLy7WVCjCj46hQt9dRvV/xh1oHIv8tKG2hyZFgHe6ppvLEX+9iZKvMSaID5DI
LXpj9+MUEf9vIOz1sONTnpgVQXEGMSjgLywPTKpeGiMT7qP0YqDcK+/koNe4VBbn
Vr7syvvE2ndScmPCGlGgPg05vCATzE3XJI6t1zBz4D/F4V7D3hAcpt8HfvtMnohs
hDCQbhkGuA4IU7ZUSJts3bJtRsebKQtn04WWsCYjYv9neWfok6TpXke1fSAuuUYe
T5sKf9jMqgO3LYxJkIjbu/LFE4pSfFbTQpGE50Q3E3n/VuK9d9c1hOPYQQ+/4gOD
K/IYPPGFyZa/S/fm+ebmcoyK4mEr+IBYOpl26z3NYYyT0ZEyhciOOSW0Bp7SdRqh
4iF58hE7T6DGYOuK4gqzN0IV9WSHXEaXW52JWSgYYoTDv4lAEPpwW8cT4xPxC+Uc
jDKkugXSm7KWVbT1dZquDIX5mox93OSxigZq0unNlh0lx9oWeqpNtls2LDbh3iJ0
lzh04pDcgRNQshZDVXo1GYN5VpFffboNj4/QU8K2zhJCiQl5G98T1UzOOwU+Y+Xg
ZnwL4pFvVN2bdrvht5opI88rC2O/CVTukd+BJfnKfv7pHwi4UZGfhFuHeLbpd/05
K88vWgDuEi4XWa4cwJHC69yvY2+dYMI598Q2pEhLCcv4sfbtmlKs5NBf4QlhFE6H
Q/QyfCQLPlpTsMeDvN0ED5MeQm44KK4dxA82I6akdvCgGHJH6jYetuUi/k/DMDAq
i8DB6DNTwYlA1/Ub5AtFU50dkZgG3NMpoaZxol2n3ZjtNRUc0yxUdZUEXFMzWAEs
o0en+ieYwf3lzAETUMwv3GcFJiIAd93REACPOgHa6301I2HHgcAdZhHbOcSY1Nlc
Su/2TLWQ4m4Jc4RF9DErQ7JenvxtSsm2aKlJEE8c72nKJES2r8/RTMfdkoTEz/9h
oHWLHoWL2eDc8hHdXYiasC0TQdK+dB5cAK9KnDQc/Ieh+4+aUA/9R1h5txVVDXn4
AxqmmCNqXFCCXwcAjJGt2IM/jR92cLizUgZlv6pl68c8jV5yZzfZcthc0K1EPdP9
0ILSvFMCulO7EA5RCcglG/ZQsVOesDXkDNgw3KdrLDlGG/7nIBY6xgMYQ6OndDtP
LPgjoCr0kns4OvyK08qWd7u7uD2vY1J4qt/w2K5whmbl26bfKwxFEIkK1OanPKEs
SzVuqJkGjcETcTjPcnPegBDMqXHIqDm0lMEqTE1lspleF49myj8CSYJ9+fIHcJzo
NeKT3NRpyMzpi37NQCINHIekTD97h2RC45mNTMyWrnf3dUDeAisnjl0jF9HbDDzK
EERAaneFNU+5gMWiFOpTb+PuBvnIN9wTMzfzXbOUUqRTh22ycAZSscPhXGwD+h6l
65s8TDiLn/N7TCqIuJhW9eDc39KT0CqixA5CsYrWE3AAZP3teOs9+fgU2Uj7CEfv
snZdnWk2ZaKq9N82KLF16ZuxcuFob4NZY/CBjhY3N1zl9Jj6vtF/+yP5tyOz00U5
7W3ju3a1xARJUDPyKqTmsa779LamsJOILsOWqH1V/y+gXyioylCyWcYNb3WOhBdm
zFk7P2GTdoIs3mZ6ilTcfLmgxqu9sT/mtlrJWSy+YvL2mHCExOubZ7aKrZ2orxkH
b5KhQ988Zjk0fMV5usgOyK03gNWBbX1bDqRPsVX1YR8YfqCk9NdrQbp7cmAi2r52
jAU0pp7tcs3E7qXAMr5mJtv1oHkcvRaYceW5/Drh1vHrjeEp+VnLzgpx8AWwC6IQ
c/h3OWXeizGOQuippx09jYEReXIybMXOeDL1hJAHwC2o2Kq5Jx28/r5P/9AFjnZd
wNbVpqSKiPLwsraWb2Oixmeqv9jyTs/pw76xeUko8KGUihxzzbLSktgBaBZ5dowz
9XZrIgi5YpVmdQft0vLX42v/N8Mgqi9Znc8CpP9hlYOG2QZ3tIC7zLhsghKrsKqX
/jhIXL3Cua7YRYF/G8XI83NTBEAjXcthZ12g9fbD0MMFvwQgiLLex+8MLM+1XKF0
3s6maNBY/hWadPuIG2JlKyj7kUOtgeHt841OjILxOkchSt9Ru0ygeGvyUqbfCq15
mne9aCVaPo8FVE5ofU+2cbiVM26oE2rUSP3kOieD8rG5j+94SXm9BttJzmEDVbP3
XZER516Ivw5QFH5MmQsLf0KRS/aOJhZUNjK9xZ8n+lxYfeThwKmuzjDbpbcERh6+
j9Pk83INpEe8gWwTazD5fTmnrKeXFxWEzZzox9LKLi/2jCcdwfkQevlnVUdOFw16
YKgW+UYgmmzDHKz9qgzJkMdGhhmijXvJE2mL29eUjTEDCnD2uAqT7ZokC6fK73Gb
dTRVPJpY6YhKI0e47XkTFeNNk6/ID1d3n2OoFQd/8bRSLNNGOYGp9uUi5w93B9mJ
WBkhNn3z92faKW36ZXn6YYaWjXCyXgq25tEvywj337bdQ++dGQ9K7ZRy1xgHRZD9
yhQyIGsBUPaowsnl7bn3v5Lg9rQembZ7J9wbrEFB77oPHr7jgM4107w374/aDGtj
5Qiq1SPMH0TeJKZQ+6Teouex43/gqY4rk2ap83QWuUzK56kyycH6GK0YXWo+S5hJ
jQ+dXGwnaT+Hx9FuSFRsa+mW+ms2SOqSJvPULCpqfpnK/9SJb6BdP0di6zujHJUu
1g3F7Hjv83ESk7EYkp6XNEFP+BEb4+Hr9ZMzsJXeKNk+7+YhKBVdDF3uwV4kwagY
I99PggYZLUg7GN+IMn+OkclukbNb3KD597m7d71W6d1Z6ZleN56x3o35aHAwUV+v
KqgbypEp4CGk3FEe+xYJ8MnQpdaaPxmFSZ5OJ5+nHakKjNRDs/DMSqcLre3BsZ7f
NPV6fBHh9r/ep9vqq84VxMY3J3mkJrbTDywFqheTdrX4x9dPkAE7qeP5Nqkx3JTR
kXkm0MWfDwBXzfiFX2jWz8/dbVpUp0f+VSZDp2+rCKLEqht4SKcYfs+iukVi/lza
0qSd7Iwr3Tb1C986p+3t97MCz34SXGSBphHDvj5n64tzgMfvs2B1EgHPTkmFx9CQ
DIw0CFJO5KWhpYhpZj2coHnVP+m2RmcbgC1vaXDj8RgcF2RTJTw88nuILUKl4PjQ
qk+i4dZ8pWjuX+rt0Oqz60rhVZ2x6DddoyS9YwFGR8nm74tRZ4OABE1M0g1DzBI4
ozglpwaEeu55TdWUxRriNxebq2VtE9STj2vgfimJRcJne2GgZkXPXl9iT00A7oX6
2CIsedKFAP/tKrM35M3DfLR4cui3Y3SC0USMx4qf0KE2RRoDmbFAZXP1fWDiHE40
ooPpQRKaB+9WOwUXwth5XnxRfSzyYSHuXtxzFdStOIvgwQ0YdVWFU71nfSpbP8Kp
6rEuXvkARDB3Zd386WuWxrTVDV4TQ5Ip/D2MDZp0mpfIGVMGlC5p9bCBctC/VNqY
bAOAU/wSg8Zzk5tzxA0WXD0+cbFoTm9FleBsFqNHm+rByFQPirtK67mVLBurweLb
D96wAbpom7ckPRpXkKJZt+Jfn+C2M33hGkzfX+oAF99Rbu2ra11PASSbGsv/ZM+a
mHL/H1OIxWbovmM8EMT/Fnw19BKgXxTRGFPmwTTDEfLJhLwqQLCcA6Y88BQ4iRX4
4Q2Y8qBdShPep1LysbpEnYI1/80Gyz/39oJ6n0FGM3oqILS6Ie+dYL2AgSyzSTld
awT/0tcjFYLfQPPW3neCVCELfZ80YdZDkgZ+YMHjRmu7hGXmQdagnPTtU7VmH/gX
tFfM3Az8mdrVxc/R8AxD9uWLONybcK0CFzjYkMY7GnILoVBWMnqDPVb/q1HqQBZh
cKKcj0uWCBNbqUqdCoE7OMCkdWiRrK6kGrqvycILKIrE+tEzEGNYOfpt7mTPuxxB
Ko2LIi6hL37feTjOn3+iW/lMvyOZi2OW7lSq/PuEHJKu1KSneyyzCDzkoaT2dGcp
04vRWmZZ0aDT0EmKmsKi9V01zSNCgExnm2CR6rGRwjvvfm2CujVkrF3x1fZr6yKJ
OqgZHCEBTo4PAP31n1AX5/vgyZ4jVawX2GI5R80zal9fi/YpiMFGDri+OQXjVvCP
3BUY/uoC6ovhnW5ytqP/jJ+IpFIKezEy1W5As3gyV94nzgeIMqW4wh1B4Y9A4RPW
RhoSEF6jt1uRjGumFU6W1ibZ4ejb7Lrij4EH3q9/QzIPWUfurl5UF44q/XLPPn0K
dxjV8jpy04shks9V6gAtZmefUT3N52qGFTB0zkIs/Sq5S4+1gwxg87kNd0UnbayA
6bkSTaNB6X5NnPmMjfWcF0rm+TIMbVU3I1xJeFUPWW/aS/r/9tIwKvxBxEgpuGQ/
ySF3yAwBXlKtQII0/OB4HlCaLN44Ki/ho+tAkyfjju1fFYjbpyHecUHiMgrqaM0F
+SrBg6e8AaLPsLUaH/QFtrQsdlIYhqDJ0xeFZbYaXBH49Nwa3IYMT5F7fGcG85c9
U/cFwqcjPX2ToRvQ6lVXHB/ZDj2uFI63f/c0r5AzgXPVdU6kSwFz7ZNvbtdnYJA1
UfHRLKbFwm9JuRY22JCNHwyUulFX2cp688Rw6hkDhEnzYICBHTLCpdp8FBP0nigu
duqpcU/a93N2g+KkdhdHTtWvxBkyOThGdsTYoF3n7rPNLIothUTg+POV12EnSn13
2RScZLW1DremN23gvVSjiwMXxE/QnyUusCJ5cpZDMlJefEKJ6zXpP1FpL4exad1o
isjO0B6YG7D1FPnALJV0sbvQzPGzNS7v6hsa9Ty0sow7Ne49R+Sv1vWcKRZ9d9eg
dPlcEdsVacNrXA/WhFmBEnjdPKZGXmzoWumfsCH/ketee4yPjitRVmeytbaqNlUe
ifQ47WnCkmS8dSckVDBQXVeSMJkOFZms5nK/kV1EfBLMfBucUC7BOydJXUTEsRYs
kJNDUQjrDUp8KeUum6thypixJ5rdCeRVHI5uBXkquQ3cTPW2LVAb2TvHPUkiIKdR
b8NXngjJfX0T4uCsVFXaHdv8HoySUI7CJz3vtEJ8P99YbQniF43rwXR6o0pwxiZF
UyTJFD7olK62KVKCQn/vrB/V8KSyC86PG+K9oXz4TC4yMMV20bm9Z8H+8XzThmPb
LO9rOCL0jzOXWshs11fjVl5x4YemJMi2nBWt6TfRZ1q+Yd1U51iy+LwvrPNd+3w9
GDVhfY3U8lYX3N2TVP906qodx4FBRQ3w9frPyWhURf6kAl+v1r4hG+8wyZFqHTL6
xQ6R63mJikYsK5jHbXHq24/Y4xhNxTWstzeDKypKz1SjfnhGdCLKLNpAJv9uQTj7
7e+qvSUCgatNbYwvmHjkRstFqKgOwGXV5xI6DlArWXrpX46meRWKoybBSBgxal2N
3yMN1vM4ZDkJ+QrfqGmYQSKzogzK5WZ1GHkDh4hJuPQMzukJrD5J7qztGty6wUzu
MuMqkwYjdchfcS3Jbw0q25hlRHFa4xLvnpKwzQ5HkUGLmEMoAhIYQBm6OHZXppQu
2IDEPM9EfrYLij9oMP2medQiP/sRc35O5WZd6fOsO6n8koWa0wTTpC43CQWpMss7
mWmIfcI0eE48hJ+EDe214qKpTvvXL71wofuNISwm2Z/Nzrv7vKqqRD6Fbjx5iD7h
g3hbl+dzMiuFVMYgvujJyT7Qagc53kjhPoBd/iHh0QUCBqZEsKIUKZ+zmnbCY6E7
BkKDOraSMLIREc9OExqAH4hT7yguP6xP8jPLAGXHWEuaSfk+Z+iamOxPsJnY4bd/
CajZvDlc+1qYoQj/KTp2T1wv0TksXGM14R7wAYarmKhfyQ5E7jlvMP3YOntokj3H
EkAB1C5mutxIPZmf3PJc7rt0P1HLHHy+IYHqvmTF56bS4SLH3ScnmuniNRhLJYTf
SKpozwiFbEOUtg+s+yyIzIiwTBEw3NBII64TCZfa9CE2mStCfxU0ZR7eAtCpPTUo
kg7pqJPkcdAx2UCdR2hF/Zxva5YZo/wBpCuOHV1hrB+OQ6yg94KXFYVyKe3fz6ml
/ERCveQqzy65Y+W6ZE7KeYMIIzuZndWYIDivQaXbEl6zU1yHrq+n3tamMCJvMgTV
kx5RLDqwRp0e2Z6YTu2XmMcgtQjrTjX/Og6qYnt7bPPvQkjvAQ+GaB1bjyBxLgwd
6j+bxqea5L6b7Kk8PiKLtxswqRcCs5CHRBU1axtDVPQ4kT0YIAAIh/U/f6ec1bDw
VilkMLuFDWtEpKs+IepMmpHmmoNOaGBxSdMHnxTMMatX3kJt12xQbOVPQjavni/j
K6FdHJ5XRKwqnxbNV4sq4P39ro89LJIYwp0VKjOE4x0bYT8bdzh6ub6oOLrB9ZIW
raZrTXoFuMlBZOckujV1+ZLeiSW+V2wXsl9eMsa0HoZkOqnJyTBAcTyH9/Naoc+I
0v6DWzCghVAe1lwVqh2MuFmJO4t8I5yGSN7QbtjqwIuLPeJatyClwtl5eT0Dgyt3
E+AE2U6SGdZq2L+VFqQtoly6zGuC/tpFD38JwSWkTaY5f46BhzNYrOesebxsdsVF
gd85uo+jTRJ+bZ//XSjPCbHLiX96T9v86J60DzY58OjdryvZmKauaWABRoQelEZM
i3454RBQv3gkrujjkb3tumZjChkomlLmwJz/AmtcHcSyIMJpdD+T/D4GgkWrzUhm
dun7pZtuR5pkucNMRqJ7637t4Ss2AekN7iq1jwKd0hKHhRyH3SgK7iDsf9GVoyX1
/h3y5UgUC+8DfLVgyQ2Xe8PLax98lExdW74AFh/nJmdajnb4OxDihDLvGcKwO+4x
0XEoaZ33kPseS5Z8gHj8atHRfzMO7JuT07AwW+zWYFmk84DDXn79CSTdbw1r0tWD
31f8zLrq6Xsvxvtgtnl8sS4rmwsNbsq92nv0Kr1cs6NE/5dqchCsGlFmiYUiRvDl
ztE2rKI86BbcATVtYdW8ZjkRkhB0ifXLgCoFx6/O0V9CFPkmtUxGBq4oQQqK75Ha
4MLyHDfcf9oJE86xQzNdgRR3l8tqetAxlhOYoF7eDScPwJzcnHwAzoQ4FQbCR+LJ
Oyg31xv1HfM/YuieOojzie3LCXUJKI+9RybYrOZhVsqPvT3hfIBqFNE/Ruirg46l
l2qAyuLqkh4aLmE8/+unml7nS03lONrK633lrLk+tqjdm3FJXI5finAPvDOODM4Z
6BZz5/9UePX/a7tvZOsmSiKrME7gVKWrLnax7yvA1rWUnRYHg1WEouuYrNrWqZRN
rBbRqly86nEUoC4R3MuqbS029F5yY7FTBEoHqvD4AL8mGjsC+TNvS6tIXJXDCo3J
ZP4kUqao+6h1V8oNBgLhfXw+Qq9XLZueR+m5+mroo2vSV0wVQ9CWAsEv+Fv7Q3+J
udCagrPYAubP+cOkx7gTwziW8HohbQR2nzYSpN86h0Igoj7opAxjZyfWXa1bFN4/
C5toJcxjhMRaRnban13ri4aeUjyAAzrxN0yROYL5NI9Em4L5WFsvJf4jNdJk0lnA
AJxBs3MtEPEUK0W7N8mbaca+e96AOf/cgXvR6Xt5gED2bB6NoWb3gibPVNjSZJ6Y
i8sE3Vf/RuDZm3laZrQI/sKt6ZqjsHidkkD2sUcT0tVLaJAg742/7NQupuf1lrx7
HedsQQpWuv2vney1XBvHAR4Dr/VQBu9tuJ+hcYGdOLtm3SWzAHOHWTyba4LgZ0LD
X5+hqNxSsnsGgm/BlRgEbtzN+25i4lokiTcDQdw1FChUMznZHk271UG57+juRmH6
6vcSRIU2/k/tNnwE8/XlFzTjBYoyuzaYqBFScF+QU55B3Xvj6vXYKZrbllSv+A0S
9JGCOsyAHb1IViCZDsShM1G2i8/stp7wxOLyrhE3sxEsujZoCzYGjiRjYWEKTpu2
0/mZU2FY/H2E7sV9Mm8iIy9hQmLnnx52n6zcRg8QArPhpvzDuWcdMJCHknDD0EEe
mchhNjqrWXkvDFuiozgUAX1PBOtY+WP/xzAnEjbdit2evZaDwNkt1YoId12TWpbm
IWZ71TCiVvUmNtT2IkYpjAE21/8qi7a3J2TglBLKp8G7UH4RfQXJTIetokft7dGd
/lpH1SHhbt+N08bYHGqnqLrerj1T9hViffpkRKZYuMJqBNvy7+TOVOV6o9pfAFEE
jafzbEH5T/jA77QHII8aX34r3BZr0fNr6HZZLll1Gg7UKIZbn32m0Wp8HqNBNram
oZgvRN4LxnNETDax1QI3fPs313qlZ6VTuarhPO4KspIjwaGrTm11BPwG7NxvlZvd
cVcgI7MMtfqzDnvK9eYeNBZQiP2vlba+5lXAh7dHhVD1xu7R+2iJtWaWEJoEKcSL
gPXA+1ZED9JY2iP2whYEfTDl9uUwhgsyGUeD2WWmId/aLkRhES1naIK/ADVH/o3I
dNXoIOELef3wTckzxSb5MmWubJ0o9JxVsnKTiEARXOuFh/oNjFgCVuBjsgjsW3lR
J2Nk7kXfGqpbjVr1/2u0mo5Pvj0BvWGvkhbr3LGMXx3oGmkB5IWRb5mJWVCevEb7
h4ARCT6orsxjNEjK1p856fzXRg8+WmVjoItCDcG5RM3n5s1uzK5WvUpaJOvjL0ju
lLHj+B8lln+/jPJTqsKdf/r7kqo/nJ3acJWiR5QqmbdKDxIZADaeW8dLRL5J/lhj
QJHougVcJpWYwzR7447LcTYeUkly8bhZ1U8FYmuM0jOVGqX9UWvnKO7iUSk54gM+
rd15YGcjdv/IoI8M24XZv7acZIB7D42TlnJ/m3Ddc4EyJ7J5VuZaj2N5XTNm9pcz
qR/5ectj57mBbHwUkwRPKlbsKqRkzwmPPj7VYb1iAi8NGaLz8+tUP/UQZa06y2xA
setAMrmOvitTlY/GfNiSwxmVVO14pXXUEf4Q33VKihLCYuHGgVE3XaEEgvhMGFy6
B1kmb/7U6+tSaMw8tQb6+ajZvBv5oOQHatwKOC/jLYf2ee1jir1x9azyk0lnYl25
8midpmi53JoxBzawiMo1qUZWzQP77jjGkJp3pZD4e7e6kpbwhW8GfZ05e94pOE/G
EQnNBjIiejW9SHl5/qMGikE9LGBgEc3N9sThXXfGF/ah/GEkp4vaBlmtMZXhm3Kb
W5DqYeBr7e4kUtgHjGH1xUUPzUwpGWOh8JDGFaC2R1Ez27cjPN/2bn5PmWSAXdrJ
Ak/ZIOdAtCjFaH6F7obe6f6z5jmfOuc7h1ep6VEV2ZkT7FOHhe7zYKuj5TWAcqaR
YNwWeEPd2XNLzTGOtURx+NnwAh9CgMOfC+fcTty8yX2muSG8rzw/LXjoQ0F+Ei0f
pL91wEux3hgOz7q3IGdXjqgl93hNWJUldRJan4G18oF57rKgZpcFV4pP3+VZadpc
06St4qBL5FsTOJuL3GZxonnamaF3JxFgaILTnSjce1ml5SayZdQ0c+oPf9pRDDI2
+8CYyuH4GhpEv520q1pgp7ClQIDo6467tHEzYvuuW3rrSvbm6aZHolBsM4owXThx
vWXx22S9heuUzLfY65OjFa0h3sdFp5XztcpexmpI//lJ6s3LYcicJj1lXjouS0jx
D5UTNyNlDwd0+iX+LGhlWAMg1IxC3gDgjNCJ267/AT0fCL6cIuQKC5gOshTm8Wr+
A305BfSc3ldHkzKBjDPGSLHeWm4GuMZJvr07ELr313M3djMkJloeq/CQ7CwwjPZ6
tnh1aoBmw6dvYHl3Fl4qBuV3KQIU2Ew67NMew8YOM8QHR31Bl5Y8/KtvFquMDV+W
RaTWv0QD+sP1FgVD3BsteCzOsF164wYkuDIKAKx738g8Zzy5SMQlB28FN4bF7zXH
/H9ZhfJu4vaYCcLo0K9RI3crrBnn4cKaRClXefjXKCWexdy2C2zpbOfTjOr/bYj6
JyKR9jcAny12fb1+A9OehWC59pF/GNI3Oj7mNP9/uxoUdKn+G88mfZSFsQLBUJtX
Y6P5ZQO5WZnB2OKfBq8AoC+uw4U47hQ9tkARrNi++oi9VWgv/D6Q5PtFobTx2+yP
hZYR9ewnbtFXZkqenc7MSMdcK2L0LBS803tuFKknaU5xyQ7hoMKHEGELV7dAIrU1
HhWJV99TyJAyPautidfC2m9E+3CBjAKlEjfPHfBc5MpCVBxBAfUV+dXqDjIaKvSm
8t6+iIeZiyLP8/9/k+LEbkbvbJefDvEmGHb4vFuM8Vx/gipvQetK0wvGdG35mVVZ
SoXK69ABBY9dglM/0FbfzR5woZEE4HaDsAB12+3yP4Nxj2QmC0WYk0MpQJqw1lQ0
qu9/OWuf7z2z1OCEAjMIceUTgP33bvvYxBiAa04Uu+kaFsa+q3YoX06u9hvcIiDi
tYjaRNfEJPQqCZQNHBKzr6vObnN+0br3ccvrnOUvIB0IpjIWnkVIWYgFFhxVAc/h
2fncgfyh119nPKxeShZCDKlHsENn8IIEUYrHXdoGt9P8169419ssY9b6+bwgnGBb
afs4V+r//OLc6riclX0yZGUIK0ZnyAsQeSgv38JX35KojsRw/jYlrKZVXAA5VxJA
Cs1VFWCR9Hob+VTds3OzvIcsvAzcQmejCJWmt4AMu2WxliukzTiV35uW+jI/PoRP
3Nl5i754Jv5XPZIBGR8C/TqfgBMYH3OYq/f4ApRmWg/RytEH4Kjv+gzjpOy2Qn0E
Ql64MrTlsmdIDTpeurNi0BHT7DCE/j/NIm4rDWjtNkKpupwgiX3ohjy9I0SdocRn
m3FoSVJDxCNvGxtQlomnQE6NyrTEFqPAVZuhofq2/Xt0mUvtz+C0cYb+gBt0TbqG
04LyqyK7b865LPD2qecY4LeZJy9IsDHVYnhIZm2UY0up2sKk/HeDbULhtDqFVKmA
xDb1qMieFV+jaBRWg364A5SvyyrzXrG/ujCtXJ85mQ1NdIwk9J15+192vbPg9cYJ
cDuqUjBi4P5OR4dsGGK4ymA+km+oqvJSyBN+JKH4jZzL2hMxih1fXWpHRydVu1Y0
MNho+iIZd1v4fyvZ3RZUvZHsnhqeDaJvyMiA0EcrFwgmIhk0XqLCfPLFj076jsgC
92bBIFsM2QIt7qc7M8MPM3DLi8GRiv4t1+OzyKp1ptxa+BdEPLab6u5aQZ/50p4m
7bIWMVkFnyd74ENwXMI38lAVOJdbf/O+euQIJBH3NAfQHichWlbVzdb5SzdRnJB5
q+sidjyINkviRDh7c/aEwqXGe1MqQNeu+ems8XK7IbleNwJQVUEVShHbzz1m4sAv
ShDy6Wu5E9epXdbsJSqLvGAKr4CcZU6rFoBidor91oYYENwmwB5qqH1TDnprvxzR
ymxQ+7xnZkmT0pJH2S0O0iB9rqWy3gpVhDl0HsBaAP4xFmKanwchWhtFYqsFkvI9
Bz79Y0HgGYaBcHwecnPxfVGoLBLgOGuPl7sOirGLHxCvgJOeDYwerElggRtFebo0
PAj5mIzuSMN1AL+mjkTi2+cW3vsHprts2HzpyGOGusyFzDlIiZZqz5yX0UtvDW2E
Ib2ythIW45i//q78hDvZ9BKCFPQxY78rImxtE74P06iWRYrbc542YOXuqRLGL2yN
zGm7LoGM1Xvx2CTobOyvwTRyPeNaBcfPOlZaKSS3XSmiscMjTcacb3DA2kbYUXKE
NVcIHKB+8XMskag26DjKBLQyAk+J+xhZBJfmoVVd7Cxn6xM8rEQS5PUS5DaMFHzJ
CUyngHnD1lDaq1MS6/3OjfMn6j9OsPyVq/f+XO7xraqNQaTsqHX/bWeiwF8LP8+a
4OxurlZtZ3kOCmkziNrTJTZyUEopn6e721Ql7DVnvjelOPAUvQYfDMjfcFkHr4lu
FeY+4a5ZOZTFTDxaph8aLWt6aUdAYMhy3ohLCb6uF1pjfvlx1ynLqu2LlSStU7TR
8RAmMsNRX91kNurtiHeePjJf+0nja+tTQFnwDok3SyOuyBWZluRpHKtRLIR1ZDrH
M1BlHbAKqa8bqN3c1Mpz0o8pRECZfUbn3FH7IMCTvKvjFeMdfjwNu2z9sfyeFgPG
FZBgNg0Ed3Ys2nhmvG+5Yynb0VTo1YsmXNdhm+uA0HD3n87usAoeRqMinngFZ6HY
Zr7+D6TdngCgPR3ksOPHZ27mKfyf5OsdiBBSIc7cn2U1k/c/0qDn9GRET/wuPUT8
48RA/Enla97JUlupViGfxykFmmdUJkY84xvL3sqom7TfgflKXwh3BDuaWuh8U6WV
WRFP8svClcQ2/IFjqjQDVEnYRtG6NfpPuVHPGDZ7K1CDxC58dWAotS9g0XYW4Rdb
i210WGaxX8cjPMYmbwsXKHUJHDurvEJcc5XA+WY93IpJHRxqfiL7XalovkWGG/4E
dVfokmalhIiigSrbAsfItYhgJCoedbUykMNW+4zBG3qvNxGuw7gLSEXG7DE3EDHK
aT4DBOyFCrE74boWzu164ZFLocr+xVtDpcAtLt9QXmURhWpCsGr0F1rLYjbnbAe5
apb42Ewzqm3M9e2arFPuDH9P1H3TQX+jaEv+oSVUFWzRHHtGlzYT4NylYq4FtasH
uPFEZRDWqYR1BSB0oP8H40OjKh5IpSyu7yEnVCUbhMP5Q960afgFIYg6QH52Izhw
AP8iGCy35e6JjwrWPPQwrAzIVfM4xa6pN/DuFmBZZ0ZY5lc/qw9+QGQWhH8AyAFr
1XktyKlBTOheGqrAM51dOgcUxoqhCqMC6es2pSJB2aogJQt70BCGaFY8OIoPNXxl
ZqXHws+tUrDvd/IKEspsgjhAwyCZXGiFcB+pAWmFe0foeJEG5qWtd1M5y0c8aNKa
BMNmRsCpU1nAd/Tn27sG0CUUxPVU26l+FBobWJVUBCaWdeEd5GR6f3Njnm5S1QM0
owHJbJAYvtRK0p4tt0JEtb97C6Toxr1nEyzpDc7BYbElXezyMimxsYGQ/4yMB8oj
RDFb7ua0vsIS5QT24z9X5SaBZSwBfSFqbN7knLrvQwm237Th1BGzFS9FSym7LkBy
DaETCCYb3Y4LmFmjlZlik12YbWTAXDJp3EeIHlNWhS7TLvzSnl+iaf0MUQs9JMz1
YYhRqPej12q8yROwi0qxxIS27aOysR3aQc8f03PiKAYBEgnf9U4xCKoZ6S8UDog7
BMilkHtCWMhmkbOCS1GeEdSE81WFHngJp1eRScDkxWOvAKTRclKcwFT0fSYs2E9Z
yOAKvv1kl6jaK23AfBBnotEK7jQR8JMWYs8t7AQ413pnlcMiUPKjn19Y5ds36+kh
nq3TU+loEIIQ+VrLpj2aY0tdbWC5AtMSbbM1BsvH/irG8g3aHaAt1x6At4gFmjy5
WEN/LOKmv+TSqixYjJMFJNQkfBhlgc6E9S5qs8/X5gOv/ukAlBOb2lHD1x6kEwV7
I5LMWsaPt2V40JYKvu8hQ/vEvJUkhwxBrF/s51F06RZJo/GJL0iAbQ9/dvd27H8Q
io6PPtZDUsvVCgqJO0lhSta+AVMwRC9s21m1keP29DJWgbjsFZvIvFcG07VJeP3L
IGrC0zdLYCXU9pgI5u1dKjg7rfyfHkofDAJdqjLKhqg0QTfR7QA+UAqo03NTFXAJ
peExRCfS+AyeyFg2dazT7ZCoPzbTGx8y7dGWjtf73YmzEozozJhvLl06+H3DlEOe
7ncXjaXfuLp1/8nO3QCozRBNTmAtGPxzTF5wErNTLxSIoCskHMKPgO6FDjviFmML
BcTrtPSg11M5wYqvo1Yf+iZMYXhmD9xqWN8KbjPBDJVKQpmhITs6DRWWi/5IEeva
BYv3aXFQEsOjfmC029EH9id6Yy/TgpuuRK+9ah6f0vGsSEvK9IEiBEaTs+UJz7zd
rW6ZF/VTMtB7TX7Ka2CWXSVsdCWQopf6/Fe3b4eIbO5kmgty7nawAscbsoQhg90G
Rd+err2PsYrWZj1NiNE4i4uQpY2yr78cJRCg57TeIiO+RWNP4Db5ez3wHovmFVdU
CQzEzFAFc6Uwfj14ONN2I13/jyG/MCWsiWYy+f8YHffOtFd6Z3ljtXqBKWDJS+LB
nNsELynwjPuHROdg8KRrEnwk1Sxr8Wu/PTBIpreqnLdIAUADgCH8FNyLfYMeQdVA
fD8mey9R/FOPXClnZoZ32vyELQOspskfWoJrwAL/yIu+aQLk6CYO6Wp1JiY8SrXZ
Y60On5KB/0eUxde6TB8G1j24AjjHLVTuz+NlG0bNdRcZq2dC+tOrK6Zlj3D9Q9r4
8QHOQznWU/En+kzM+uC4xQK3UNfkHQSvpYXa77XZQPOQF7PH6dF/Q1UpsUa+hhhG
hhiSmxVFbDJdZajdthPHxEznp0H6wiazUmH+QMAhGHRD317lnsgZqm9uihCzgf7x
tbpCZDQbt1/UoMAsD5WXdK4jNoTjlG7uFUsS4MZYlgFxz0xG2aExPuhfZWCrneR0
MJCfazUypLeYE/YBnhN4WMEhcGHlxWQJhg+ENiIaaXRxqQdULlstVfq3r7SpvGDE
G3IVfOw8QrgpqMpQluXxsIKXoaMB3UqhP0hjnJI+XkHJ3hp69gnZFPNjDJf9+fi1
1LiCylUNznpS1Ms6OxyHDQKMcqQZG3iTANJHhSqiRpBgZXFVT7F7N2Cvs/nwTOFM
SF6CtYeUqJp4dDa86Ga7/wIRs5s9gRL/qXfUZ5lLbGJt+vN383heb36sdMmcjUCo
zV9iV/uwY1TZYh26xveVKoJQ+e+drJLgQ1tY8RIdTpPaDVAKgXF0bdTmshCiQBjb
U1XFSddkMVTwbFSWeMMM+GoHs4rT2BLuB+lPE888sf4TkAlbLdo1YNVYvwlK4I5R
HgfykrRzZJErRwiclvKblqJnwdoG2MPaAbKyWpSBs3irXuSVRxg8ayT1/IfYLB6O
FaNVZYx4Glytbs/7QvMy60OiFTXf85n/nZguuhw9lg627KKgTrP1qJmcg54jFIMd
NAW1qiqI16jCzpGC0+kRe3u00ICc5e2hFPJoSEJWclYXOn+12dbccWlyfK1Ks8of
BIh1cO+gMwVahjXzNZP834F/2X3JOywefXFKtylsHUysPS1P0NnurBEXVmeLQxtY
qfJc4jbFW/IHRWA3BFHXegMvLZqoi8YMZ2O8rfYUxJncO9TLfkOurGrjGuoWpqCd
ruzKlcubkTTvEzIizjlm2j9VPPfamffJPz8TKKFNWl5QOuPI452ApO6yCkqBP7Hq
G4i4z5I0UG7gq6B4EFeDoS1Z2j8QIDADZKRd7y5p5Olj017Nw2kgi3KzbCwctyqE
I1aB7sFS1KZ9HsthOLWG0nLP+ej+Iz8XxTEpbkOlFM+PP4Gg8YrK0knCjvLxCwre
yGS//ktRrivqhLlvcG2DEtkCG7XGewRyiZGBlx0gEnj3K794UOaHb363f0aWASfx
E7dibkxAes/BYJT3/WEtnpyO7rX+k73UmDsJ/Xp+cnuPp+rpNyGybSOTg8q2SZ2+
rMvnhfsSxzA7D1ueLq13yLgzKttZ6JyXWAco2Yky7oN3ZjqlhN/vWYMh/tI1sN9r
3GwHsRwWozm9KibO+ey9gOQykoTaH/QWujmGl4rmgjLZKhzMbM7TNu6v9MsO3qLA
+yEGRjEW1uV6e3/0Sq/CxhbUzhnjwEiNa0vxrdYZzxPdSXzx34MuoqvAbDE9hcR7
cJIVkAqALaLgxdVXAKC2pMJVI/FYKvBQc2xk58KVJyP2QF1idUIz3Nb7d5ecdAhn
TB8m9BYbQwUZMxUo1NDHZVMkIjmf4nxii1Xay/rToRPNs95XSyaRSgz3+ELSVXQ5
8Oatw5IFX6feZ2chncVHb+vsCRK1HesqYSbhHkKOdy3IPE7KtF5IFRPEzHEBs1E+
NT8ZJlMPO3Ob9amS49O4qw8o9FKQLKR0f5aneCk3k+d1g/nZfmDrFNgAZNYtCHr9
3NkZ/Vp8iNU1Es66CV2W80DN22FUS5xe2ODB6gAWrAry7pwQPgIedj9oX9PcZQzs
yGaGJizx4NUastrjy66Ha4vwFHusiHuW10DbHERzwrIPk59sY2D392/f4LrrXpVC
fyafFp0UHz8YqbsX/RC3ek6N1y2pUrEsrE/+GsXgjKuSpezTXQQjvq8/O3ZwYChu
z4MIodhIytuj+TyChGmIZmD56EGH8UVXoGmdm3Km5JZV0DHzjnfeiGkD+jWhTdBg
YdPtrVpUnjm/P2Ydp0CiblXJZF3iFiZe0Hp1dW4rQIJdAsi4jIQz5NpCEkT/E73k
/6H/40PUMzFBjRKQ6bJnMFwnpei0KZ4yOzDMFdCZHQXhztu45J26CtdN8IqzLk0z
s+j77u0YVmEmEOhUFOoZeas3lo4wZStYB82Dr5M+Qs6Vmvfl9CV+2dkwTC7OM0el
bYBoJELeHG200Q/UFCRLVEzX5Bxc+oqsOt6BIxnfORActz2ABc3Z6/bmz2P/ER1R
CTIuZOUTjCvSxWLtPFXrMorMTwABMSjxbX0umLDeUKqjOat6H2vDHm/DIGiLcigY
OR0SiR99EPZQpB2LFJ/C2Q5JfaiP6Rz/QtZLHFX8HRcGIp49xZfhut+D79TISUu0
wb/JKGGF7aob2B/KpGgInaKP5SXo3s9HPHZNh4YsHOj/H69PMpp/iSlwmx2cSdZU
CKJL/w8kMrwqckNOBYH71iO0jb3MSSXnc67MIR2JWHKFLeEHsL2UWxxzqgzmIBAn
1Cg59N3HnIWMpEot1ulco9UVtndqH/DgGnKTZ/U0dJJ0THhE5NV2RTXaJ1msEPpL
Dj4EDGYrdoxoFuRRJWTECvGgmt4nb1gBbzEc/mX/JMENFhAuIdMlbuSh7nTQbpsv
j5vHbK1Pd+umZceCZ47G5/EXnjYOE8vQrOywmr3v7HN3s36P2yhjq+paAxy5S0HC
tqxRwuHz7+77LtDOCO+fwW/sbIEndkn1pCi7fPXmUxDrZL8FSBY0WXoTjBoyd0ek
9MGjtr7tNkor+THQpELCp1AMeJbbR4ClZqhxAf56j5oLu2dvDxTnPBRj0XvT84Ty
oK763j7i0rjqmTN5JR+M3HYxxK3wShWTn6v+tKTYWZQOJJD/JKD94a2l+BW1xqsY
2G7pSaMnqgy9cTkbkUMSwaZgGQSIDZEW0+aN19nj9MpnpQ2WpnwYud1xxrjGd6yj
TEOeaXT9irTaEPmqnnvQXytwqWhOM6mcAboqUr6PELLUnUdC0SByipeWj48kHxbv
bjuGPKeX8pAAqouLm/78wWVw7kpBZvOWd4ZGlqnhb+bv0mqzD6yZFMEvQTmmpfaY
3V1XM8vVdMjkgbrmH252HxtpCDp5dvuvJnJHU7ZNGMFiiSbr06XKTRsC9tmJ7WYT
VhZPsbO0/VqVii4TUgVgDGjfnyu+hx7aXd70oHXUTP49Km+61Xgt5En004xDC1tn
+iurwqr9N/mYq8lfy37qENS695lmdLoHose2c3+4T70GlOfVIbtkLjuLQAKzAjbt
HKAuGBW5ou2LvETr0O6+s33U4/q95NMrzf6X4F6KTkEbpz8P2oyuKuX8/8TfDpy+
A7A50dUXRZDA6iaNwbhu7bLYypjweNwqNM77CpqmEiW3WPG7E4/T/8QI2ZvY2avd
WMcPZcqQ9l5/xsc+LRqOp5E46s1qKXMV7wje3+eRpu71GR3dJpp/29N0bKWMOk7q
xr7NVAP813VhpaLCxA1BFtedhan1zmGh8KAdWLWDfrcjXRyBIkWK0XGH3y3oHwEc
qIV/Laiz1kdy0LSCCAvaqCCuCwoGNAWz13NYRaD7YRmVVl52j9ZQjpARq9RAI3ju
8DDAOtCq1onII/bmtv6gQFBdYZaXf0/VA8pbCoLffmvC1+z8ScE8ivzWvMQQOFkD
kRyKqDwI1fjPe/Kwsm3DBJQbaHWAtEuUyvITmWKlerzpqsLH2bQYcBOncTozBU1C
fU5vDzdB2Qy2rqKOBdwqQC52X/TaG3fwyFwmB6fxinLI5Vtb9nJ+hkePAJvTGdXs
M7tYzI9ONmb1dWdI6FAx3OrT/5RnTLPx4LfQJdZJSyJJF/U2B3rPiuFOYTpvx2o7
Pp++msqyAPL7fC9r8ylJiST3oufVf3oSNTS8iXSnlo2/emnNFe2rIbr94sXm89dS
+PdVPPtH6G+BUKh0hof8zx7UEmuw4bhEuT3SFB6MfWmQcLTckKKz/YjgoJVjkSYO
YByRme0CWwyJV0rZfpEoJCD6IiDOCKOBF3+kX2cPSe6+aTElSEO6KIJ8qW2jc3wr
SH7ScN5H4TeKN7VolPMjZv2Swxv/Sz/47GDp63KPv2ijLpqAAMYrI7nrTJgCqKaQ
Dc+xsvkKSGeZXj0HXiFSTO6O2ZDydg/huHNUb3PLs2XJUAClvw4wzRrxQa17HV+x
04vx6shJ+1XzaOY0qFsspIwpLU5pRu6ObQtitF6BwhXutbdicKp9C9l7RzsDzrkk
oF2cRrxOfck3kIPhABc/FwH4M6dlP3uDqm1sCbVZniztRwIjIpSP/bfPuJIMfD6d
SriydcNWY43f5P/vkZ+hVh+DJIIwRL0xlp1rX2FlXRBjN9+R3q3WtmA7lLE0k+pt
dqbuGNDbYNZ5Zu9kXVYme/1iRBHsEVE+7v0C7449lQUxUUNw5c+bFQwKQC55ae/T
KGKvjtZKeb7QgC+5LsW38tSO6jMe3qriHsRN+T4CjCtmg3EN2DuxFUzR6trdRxMI
lOTszc5cmeknhK0DUPrW3UlHGY5nI6AQEthymjQpL/w/rFlemK0cwSMhI3GKIbuN
0U6ghBUJ1Gf9GrZTeOZKja4VdNXOF4RNVJQ288a3cx8/B5NaEhdCBiBdrW+dnEe4
3sKdIv0la422/QrQ/aYYll5XV5uzRVRrVa9F7RPy0K2c3CtuadY/UyVcssqq012o
ioC2MokvYKqojvW34UJ+XHIz5Z3hqy+LymjfWWky+MPrApqS47hmk4Br+v3znD0+
ltfE703GDvhplJVrpGBMvwkD5k6kjIrGgqGG9atmmkj1j1fwuKVt6q/a+Ro1LbHH
ASKAjFZb7ap4rW3iqw6DpW0qW1Mz8cCVS7RbTC8iwmqsKb1aWQ3tFW+bXRw/Hsr6
2loQk420QSPFA8aNNaNi0wye6RxB/XpLIhKThylobInbqO0iygRtMAA4HTVQvvq2
9iBrt6i1hYxd8a6rSE+raDJfT34FvVcBYZBQdaOvWLMauKOpThGa0TTxBtxPut5s
PZlKN+XbZ8J14C4+xWS59pq9CWSVwi4asOrjoAs8BpwazmClf+EbrrYeVB99oaJf
q/i5rxggy4iuLeBNXTlFhyy/MdT4ZLyz6uVIBVpAKYzpEEdN7/42/yvxDNZiEjaA
7mVX4yRr2K6q0bXwsS0r4+dU4NfAdAE6AIAq8asWQufrEz0Royrw8dsIecj0/tmw
a8y+uJKHBV42LbPk4N9UvwWMAUDfb8++ax4vt9U8Oho5xYzRLykqm73Mdo1yQr0I
cBufhydpLjd3ErbH8+mXiId37iB4htnDnLUiIiS5eCjgmOyetPj3gegV2ceiJtkX
4JrrMmtST2eY8ALyQMFU/ogpoFxf/sHqFdhCLQfKmFO6Z+MWaEAVY/cS/AWjM45r
5wIxZj6ci1SI7lTwDxe9jm5XGZ7AwKw0uLxNH7J85DTgv411AJwetG3QPyxKfu2X
tkAL/TwU+zzeLA9qq3GPvsrlTmKZfFOb3Tm7si9/UgTBo/x1oGyd3uzcw0BB/AUf
Em0En92TrvYOyAeVhd5WUD7soaDv5lqGgJcmthBhHevjnHKUDNKk9wRuN0da8qTJ
T/Ump+bizSby3uruors+OuRBsbeMka76mpcKODbDMvqCd7p2N/2oQi8WzylNTF0n
5fNh2WPo2G617vOivvrddZ3vpw8wB8LWLV0Um+bF+deSR5rTdN31K3s2kfzPvABF
jr4ktGwcRTRzImEuDp9EaQ0M+od9LhvYsVHJ4YoUwxRli9JfZDQbBbDeQCNDifa4
CRYaxY7H6tBcxu91PukDX1RyvNvcnMJLPLVBEcMhCkRKHI+Z9Y0Hb60HbkTk+50v
rCH8mAa4m1yHlhOr5kCgBxoKP0q4lb83knSQxYYBLo4/qimsC3CH2cSUk+UbY+mr
B8y7sCoptUxTKcNPuBsemrF0cBjJ3bPt2f2vHbJqoiHWX7yDBQIdzqNKWbKm157A
0KpTGIZwZ1AyuNkFcP4ZjAqGdd3tA/xx53OAiykyBOMYyF/kZgTmuGb7X0jd0jop
/NWGjlo0qeOFwfpv2t/71o2zD9LWiifBLR5rcEYMr6AVxQFL1k5s9+PbdFD4jqE/
la1pxFUXJgeMVs1zpkc0xqYamtvbXNyO4VG1d9SFUUyFrC2MT6PXIltTaAb5oi0T
KbtSOHCqmvfXwAJnwM6Ue0PkM5oJYR5MvY+7Q0/obiZNG01SboVmz4HOzGMqDNkB
9MwqUJR/B+j/nzM7xvA9WBYniiHVjgmdhHp29YNxG3POAA2W1wj7pLK4+mTkGhCJ
UTmRcId8e+DRVq2YzVoVBv+l37ZJL9jFBidyMWzW6H3Z70pXIpA7bNKe9PsW407g
j9fjED7gBHcHix2zmwbbN2o9PloKg7Dcxr+Eh0nsJipHItdm7dK24jYuc2LWJMM7
TbqX/mLEMzsiwTN52beUkWLvbqa8s24RKkcf7aYZOC1HcM04Ded5TBa4iVD86pSz
JVXoxz205We5EZH5h7mXPm1YeKQh/bFn1PDDlswo6DNofpvTxAUR9yjQDTSGwE67
uo4V1xWfcToQUbxQ8pjLiUDTewwEslpk4teeT4d3YsOhGknkbCZK7iC5F2bWoL9q
CBsybScZaE8ZKvvcIFhE3cBV/ylNLdyStmjHOWpt3Dt2vOwi4PeprtKkRqJUPZc4
8UM5k63PXwp7P950qvDs+9vYwwv4CF43KbdyUvq2AttbyxhB8LnlQY/M3A2I9lQq
oWPN8nIsNcTpWS5jrmmyuHkBF6FEJB78vwxkcH7CJsi9bFzeb7XEhgckb3dyOUc2
lp/keF9bXFVT7XRyCpzro5mFHGquiRowd5Bpime0GEuDoN82T+RmkquAwIixW0QI
ygTQHpHTOEtihaZniVGZ/D5Huo+VY7lmB5ZCj/dACdLqm2KHGoVlB/Se6wc1Brw6
6S46n5cVKe1wzdOaUqFGJwdtbt642HNoGVnYoG/3H/PdI5jmen96nXPWl3M7MMZO
PapsnYyTEYU1+6bx0gJm1Zngy59wFoh1tO6R/GQkCE+0OhTbBEUOG1xBohFpljL1
NIkibxb+D4fGMHB0t3VkIDy983s77RP+hJxf2ZbabGzfk29NSYGM0VEQ5wDqQXdK
EZrnN/BRyz7NTgUqhSYTduReveRHseqRwTpckd2Fd/6B3m7XChTieg+GuKc2v83U
KgSi62hNdmZd8hPLx4HOzvhGcLp2TaT7+Mue1GKjXlhPvMW742ygg4/CVeytl7o2
hkXK1mAgIW1EE4kbDIZ7t5CKZf6pl2MLwLRmVZLl6AiY+FFnvycaqUqP9o9DaaQA
cLYKdMCa/Wz4zT4x39kyQbz4r1k/bHbZi833UbTZ7UkvoJJ5mRpvztXngW/SKg7J
tiRhQKV5mX0FVv3gn9H3KMPy2XCE9CIYPFZ1WCzyVbumZvspz+7VH8kyXgeq7jUJ
PDXZzXyVnp9QxL5/lNIug9Ycz+gdwuBAfIC5SQzYf7U2qtWO8oHhGmnTRfKXMEcW
jIHSY/6dQE+S70JXoQvxV7NxQLHAO7EeXxp9kwYQEB2O//cpsVYG96B0fUXCED1G
BxOGPLsacHQFn//jND8+6SLL+D6IKJq9/JAil5PurvnOhS8HHaFZHhWg7nzfR7Gl
/xNdfk9UlJdO0rPNfkWzM6B1KqUWJ0eH2sqWfowN0y0WjearF/0TbrG76P/SJZsN
euiGHWTB6FY7nGTjYCKXDKCBv+GjK95fuZ64HjbehRSul8BmU4o9HGpjTQMZkoEi
zgRgxSYlAZEqYQlq0TqEOSmkW5M79d6xrxHAskk+a2QVIKmwJlAzrFtoXGwq4Gab
tBH4BF9LYI9GIgB/VE0BsyTPM53pdn3o8RhIAM4kHz3B4Co91ipepNdwcswtFuiT
rbjfH7WbnHU1pjVa7DcKrR7l2S7lJzb9SZEqekyn0BlmVqwm6/T0z+GaYJNLPbEH
v66Hgt+jkA6M53TEzWYsz8rYBkkcN4OXaxQzDGFcm5cVtt9q8BtcBfT7pgVsFbmN
4CT0mpE6ebtl2NInVLo6zSssXkQeH+eKr9mRlA5J7qOBWZnkjFpSv9yDiAd2YbrK
woAubGr7X4gfndjd4iKVxhsCot3wtL8AaBskcVpYm/vsF8dvG/fTVFRk26ixtXp2
6bowC/Jw0oRXfHJ7dSSl43nW7u7lt/T6abSrwbjWcwhTNNlJEdl9zknU66XWmfRc
OfGQQZUqy+JOpA2L3xKMWsyMzQ5g9/p2Y+nF0sUM2zabfX8P2wkaaEj+MEeAH1wc
FFdny8xEw03uwE9gOkb5RBPMzfnk/w4Y2/MMWRY50NhRhkYdvSpmCK3s63kUgoMw
dtarE9KEqfleC+fuG3u/hiT0CI0p5/glmmmpWUKocEwlQDtH58keokqwpIZaYsVi
9uVMeM4omXHwZ7ptrwNQFrUB3i7LOC3GKEBIzM6C9JFtSYOujrvfFRo9QgfoA68+
ZODn51pwXM/VSRPfijKLI7Gskvx3hxClCFXZ22ZePpaYyNolKqffRvjcgfElhFi8
63iWIFo3MvaWaGPhMmY/rkB2ZSixvkme1shybKlycJKKuobKCRCvtIqyTInsGI0x
HUPhhEdr2P5rP2E/971uCkEUYTXYqFrWYugdhmlluZPYcBGKhZZhY4U6BpTZUmRj
0HtaQbrcAshMjrRRreoXvumpPtyXNeLSpNjArwzKn1g=

`pragma protect end_protected
