// avmm_interconnect.v

// Generated using ACDS version 22.4 94

`timescale 1 ps / 1 ps
module avmm_interconnect (
		input  wire        afu_slave_m0_waitrequest,                     //                   afu_slave_m0.waitrequest
		input  wire [31:0] afu_slave_m0_readdata,                        //                               .readdata
		input  wire        afu_slave_m0_readdatavalid,                   //                               .readdatavalid
		output wire [0:0]  afu_slave_m0_burstcount,                      //                               .burstcount
		output wire [31:0] afu_slave_m0_writedata,                       //                               .writedata
		output wire [23:0] afu_slave_m0_address,                         //                               .address
		output wire        afu_slave_m0_write,                           //                               .write
		output wire        afu_slave_m0_read,                            //                               .read
		output wire [3:0]  afu_slave_m0_byteenable,                      //                               .byteenable
		output wire        afu_slave_m0_debugaccess,                     //                               .debugaccess
		input  wire        bbs_slave_m0_waitrequest,                     //                   bbs_slave_m0.waitrequest
		input  wire [63:0] bbs_slave_m0_readdata,                        //                               .readdata
		input  wire        bbs_slave_m0_readdatavalid,                   //                               .readdatavalid
		output wire [0:0]  bbs_slave_m0_burstcount,                      //                               .burstcount
		output wire [63:0] bbs_slave_m0_writedata,                       //                               .writedata
		output wire [23:0] bbs_slave_m0_address,                         //                               .address
		output wire        bbs_slave_m0_write,                           //                               .write
		output wire        bbs_slave_m0_read,                            //                               .read
		output wire [7:0]  bbs_slave_m0_byteenable,                      //                               .byteenable
		output wire        bbs_slave_m0_debugaccess,                     //                               .debugaccess
		input  wire        cmb2avst_slave_m0_waitrequest,                //              cmb2avst_slave_m0.waitrequest
		input  wire [31:0] cmb2avst_slave_m0_readdata,                   //                               .readdata
		input  wire        cmb2avst_slave_m0_readdatavalid,              //                               .readdatavalid
		output wire [0:0]  cmb2avst_slave_m0_burstcount,                 //                               .burstcount
		output wire [31:0] cmb2avst_slave_m0_writedata,                  //                               .writedata
		output wire [23:0] cmb2avst_slave_m0_address,                    //                               .address
		output wire        cmb2avst_slave_m0_write,                      //                               .write
		output wire        cmb2avst_slave_m0_read,                       //                               .read
		output wire [3:0]  cmb2avst_slave_m0_byteenable,                 //                               .byteenable
		output wire        cmb2avst_slave_m0_debugaccess,                //                               .debugaccess
		input  wire        cxl_compliance_slave_m0_waitrequest,          //        cxl_compliance_slave_m0.waitrequest
		input  wire [63:0] cxl_compliance_slave_m0_readdata,             //                               .readdata
		input  wire        cxl_compliance_slave_m0_readdatavalid,        //                               .readdatavalid
		output wire [0:0]  cxl_compliance_slave_m0_burstcount,           //                               .burstcount
		output wire [63:0] cxl_compliance_slave_m0_writedata,            //                               .writedata
		output wire [23:0] cxl_compliance_slave_m0_address,              //                               .address
		output wire        cxl_compliance_slave_m0_write,                //                               .write
		output wire        cxl_compliance_slave_m0_read,                 //                               .read
		output wire [7:0]  cxl_compliance_slave_m0_byteenable,           //                               .byteenable
		output wire        cxl_compliance_slave_m0_debugaccess,          //                               .debugaccess
		input  wire        cxl_io_csb2wire_csr_m0_waitrequest,           //         cxl_io_csb2wire_csr_m0.waitrequest
		input  wire [31:0] cxl_io_csb2wire_csr_m0_readdata,              //                               .readdata
		input  wire        cxl_io_csb2wire_csr_m0_readdatavalid,         //                               .readdatavalid
		output wire [0:0]  cxl_io_csb2wire_csr_m0_burstcount,            //                               .burstcount
		output wire [31:0] cxl_io_csb2wire_csr_m0_writedata,             //                               .writedata
		output wire [23:0] cxl_io_csb2wire_csr_m0_address,               //                               .address
		output wire        cxl_io_csb2wire_csr_m0_write,                 //                               .write
		output wire        cxl_io_csb2wire_csr_m0_read,                  //                               .read
		output wire [3:0]  cxl_io_csb2wire_csr_m0_byteenable,            //                               .byteenable
		output wire        cxl_io_csb2wire_csr_m0_debugaccess,           //                               .debugaccess
		input  wire        cxl_io_clk_clk,                               //                     cxl_io_clk.clk
		input  wire        cxl_io_rst_reset_n,                           //                     cxl_io_rst.reset_n
		output wire        cxl_io_master_s0_waitrequest,                 //               cxl_io_master_s0.waitrequest
		output wire [63:0] cxl_io_master_s0_readdata,                    //                               .readdata
		output wire        cxl_io_master_s0_readdatavalid,               //                               .readdatavalid
		input  wire [0:0]  cxl_io_master_s0_burstcount,                  //                               .burstcount
		input  wire [63:0] cxl_io_master_s0_writedata,                   //                               .writedata
		input  wire [31:0] cxl_io_master_s0_address,                     //                               .address
		input  wire        cxl_io_master_s0_write,                       //                               .write
		input  wire        cxl_io_master_s0_read,                        //                               .read
		input  wire [7:0]  cxl_io_master_s0_byteenable,                  //                               .byteenable
		input  wire        cxl_io_master_s0_debugaccess,                 //                               .debugaccess
		input  wire        cxl_io_slave_m0_waitrequest,                  //                cxl_io_slave_m0.waitrequest
		input  wire [31:0] cxl_io_slave_m0_readdata,                     //                               .readdata
		input  wire        cxl_io_slave_m0_readdatavalid,                //                               .readdatavalid
		output wire [0:0]  cxl_io_slave_m0_burstcount,                   //                               .burstcount
		output wire [31:0] cxl_io_slave_m0_writedata,                    //                               .writedata
		output wire [23:0] cxl_io_slave_m0_address,                      //                               .address
		output wire        cxl_io_slave_m0_write,                        //                               .write
		output wire        cxl_io_slave_m0_read,                         //                               .read
		output wire [3:0]  cxl_io_slave_m0_byteenable,                   //                               .byteenable
		output wire        cxl_io_slave_m0_debugaccess,                  //                               .debugaccess
		output wire        debug_master_s0_waitrequest,                  //                debug_master_s0.waitrequest
		output wire [31:0] debug_master_s0_readdata,                     //                               .readdata
		output wire        debug_master_s0_readdatavalid,                //                               .readdatavalid
		input  wire [0:0]  debug_master_s0_burstcount,                   //                               .burstcount
		input  wire [31:0] debug_master_s0_writedata,                    //                               .writedata
		input  wire [31:0] debug_master_s0_address,                      //                               .address
		input  wire        debug_master_s0_write,                        //                               .write
		input  wire        debug_master_s0_read,                         //                               .read
		input  wire [3:0]  debug_master_s0_byteenable,                   //                               .byteenable
		input  wire        debug_master_s0_debugaccess,                  //                               .debugaccess
		input  wire        side_clock_hip_clk,                           //                 side_clock_hip.clk
		input  wire        side_reset_hip_reset_n,                       //                 side_reset_hip.reset_n
		input  wire        hip_reconfig_slave_m0_waitrequest,            //          hip_reconfig_slave_m0.waitrequest
		input  wire [7:0]  hip_reconfig_slave_m0_readdata,               //                               .readdata
		input  wire        hip_reconfig_slave_m0_readdatavalid,          //                               .readdatavalid
		output wire [0:0]  hip_reconfig_slave_m0_burstcount,             //                               .burstcount
		output wire [7:0]  hip_reconfig_slave_m0_writedata,              //                               .writedata
		output wire [23:0] hip_reconfig_slave_m0_address,                //                               .address
		output wire        hip_reconfig_slave_m0_write,                  //                               .write
		output wire        hip_reconfig_slave_m0_read,                   //                               .read
		output wire [0:0]  hip_reconfig_slave_m0_byteenable,             //                               .byteenable
		output wire        hip_reconfig_slave_m0_debugaccess,            //                               .debugaccess
		input  wire        int_conn_clk_clk,                             //                   int_conn_clk.clk
		input  wire        int_conn_rst_reset_n,                         //                   int_conn_rst.reset_n
		input  wire        usr_avmm_hip_reconfig_slave_m0_waitrequest,   // usr_avmm_hip_reconfig_slave_m0.waitrequest
		input  wire [7:0]  usr_avmm_hip_reconfig_slave_m0_readdata,      //                               .readdata
		input  wire        usr_avmm_hip_reconfig_slave_m0_readdatavalid, //                               .readdatavalid
		output wire [0:0]  usr_avmm_hip_reconfig_slave_m0_burstcount,    //                               .burstcount
		output wire [7:0]  usr_avmm_hip_reconfig_slave_m0_writedata,     //                               .writedata
		output wire [23:0] usr_avmm_hip_reconfig_slave_m0_address,       //                               .address
		output wire        usr_avmm_hip_reconfig_slave_m0_write,         //                               .write
		output wire        usr_avmm_hip_reconfig_slave_m0_read,          //                               .read
		output wire [0:0]  usr_avmm_hip_reconfig_slave_m0_byteenable,    //                               .byteenable
		output wire        usr_avmm_hip_reconfig_slave_m0_debugaccess    //                               .debugaccess
	);

	wire         cxl_io_interconnect_clock_in_out_clk_clk;                       // cxl_io_interconnect_clock_in:out_clk -> [cxl_io_interconnect_reset_in:clk, cxl_io_master:s0_clk, cxl_io_slave:m0_clk]
	wire         hip_reconfig_clock_in_out_clk_clk;                              // hip_reconfig_clock_in:out_clk -> [hip_reconfig_reset_in:clk, hip_reconfig_slave:m0_clk]
	wire         interconnect_clock_in_out_clk_clk;                              // interconnect_clock_in:out_clk -> [afu_slave:clk, bbs_slave:clk, cmb2avst_slave:clk, cxl_compliance_slave:clk, cxl_io_csb2wire_csr:clk, cxl_io_master:m0_clk, cxl_io_slave:s0_clk, debug_master:clk, hip_reconfig_slave:s0_clk, interconnect_reset_in:clk, mm_interconnect_0:interconnect_clock_in_out_clk_clk, usr_avmm_hip_reconfig_slave:clk]
	wire         cxl_io_interconnect_reset_in_out_reset_reset;                   // cxl_io_interconnect_reset_in:out_reset_n -> [cxl_io_master:s0_reset, cxl_io_slave:m0_reset]
	wire         hip_reconfig_reset_in_out_reset_reset;                          // hip_reconfig_reset_in:out_reset_n -> hip_reconfig_slave:m0_reset
	wire         interconnect_reset_in_out_reset_reset;                          // interconnect_reset_in:out_reset_n -> [afu_slave:reset, bbs_slave:reset, cmb2avst_slave:reset, cxl_compliance_slave:reset, cxl_io_csb2wire_csr:reset, cxl_io_master:m0_reset, cxl_io_slave:s0_reset, debug_master:reset, hip_reconfig_slave:s0_reset, mm_interconnect_0:afu_slave_s0_agent_rsp_fifo_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:cxl_io_master_m0_reset_reset_bridge_in_reset_reset, usr_avmm_hip_reconfig_slave:reset]
	wire         cxl_io_master_m0_waitrequest;                                   // mm_interconnect_0:cxl_io_master_m0_waitrequest -> cxl_io_master:m0_waitrequest
	wire  [63:0] cxl_io_master_m0_readdata;                                      // mm_interconnect_0:cxl_io_master_m0_readdata -> cxl_io_master:m0_readdata
	wire         cxl_io_master_m0_debugaccess;                                   // cxl_io_master:m0_debugaccess -> mm_interconnect_0:cxl_io_master_m0_debugaccess
	wire  [31:0] cxl_io_master_m0_address;                                       // cxl_io_master:m0_address -> mm_interconnect_0:cxl_io_master_m0_address
	wire         cxl_io_master_m0_read;                                          // cxl_io_master:m0_read -> mm_interconnect_0:cxl_io_master_m0_read
	wire   [7:0] cxl_io_master_m0_byteenable;                                    // cxl_io_master:m0_byteenable -> mm_interconnect_0:cxl_io_master_m0_byteenable
	wire         cxl_io_master_m0_readdatavalid;                                 // mm_interconnect_0:cxl_io_master_m0_readdatavalid -> cxl_io_master:m0_readdatavalid
	wire  [63:0] cxl_io_master_m0_writedata;                                     // cxl_io_master:m0_writedata -> mm_interconnect_0:cxl_io_master_m0_writedata
	wire         cxl_io_master_m0_write;                                         // cxl_io_master:m0_write -> mm_interconnect_0:cxl_io_master_m0_write
	wire   [0:0] cxl_io_master_m0_burstcount;                                    // cxl_io_master:m0_burstcount -> mm_interconnect_0:cxl_io_master_m0_burstcount
	wire         debug_master_m0_waitrequest;                                    // mm_interconnect_0:debug_master_m0_waitrequest -> debug_master:m0_waitrequest
	wire  [31:0] debug_master_m0_readdata;                                       // mm_interconnect_0:debug_master_m0_readdata -> debug_master:m0_readdata
	wire         debug_master_m0_debugaccess;                                    // debug_master:m0_debugaccess -> mm_interconnect_0:debug_master_m0_debugaccess
	wire  [31:0] debug_master_m0_address;                                        // debug_master:m0_address -> mm_interconnect_0:debug_master_m0_address
	wire         debug_master_m0_read;                                           // debug_master:m0_read -> mm_interconnect_0:debug_master_m0_read
	wire   [3:0] debug_master_m0_byteenable;                                     // debug_master:m0_byteenable -> mm_interconnect_0:debug_master_m0_byteenable
	wire         debug_master_m0_readdatavalid;                                  // mm_interconnect_0:debug_master_m0_readdatavalid -> debug_master:m0_readdatavalid
	wire  [31:0] debug_master_m0_writedata;                                      // debug_master:m0_writedata -> mm_interconnect_0:debug_master_m0_writedata
	wire         debug_master_m0_write;                                          // debug_master:m0_write -> mm_interconnect_0:debug_master_m0_write
	wire   [0:0] debug_master_m0_burstcount;                                     // debug_master:m0_burstcount -> mm_interconnect_0:debug_master_m0_burstcount
	wire  [31:0] mm_interconnect_0_afu_slave_s0_readdata;                        // afu_slave:s0_readdata -> mm_interconnect_0:afu_slave_s0_readdata
	wire         mm_interconnect_0_afu_slave_s0_waitrequest;                     // afu_slave:s0_waitrequest -> mm_interconnect_0:afu_slave_s0_waitrequest
	wire         mm_interconnect_0_afu_slave_s0_debugaccess;                     // mm_interconnect_0:afu_slave_s0_debugaccess -> afu_slave:s0_debugaccess
	wire  [23:0] mm_interconnect_0_afu_slave_s0_address;                         // mm_interconnect_0:afu_slave_s0_address -> afu_slave:s0_address
	wire         mm_interconnect_0_afu_slave_s0_read;                            // mm_interconnect_0:afu_slave_s0_read -> afu_slave:s0_read
	wire   [3:0] mm_interconnect_0_afu_slave_s0_byteenable;                      // mm_interconnect_0:afu_slave_s0_byteenable -> afu_slave:s0_byteenable
	wire         mm_interconnect_0_afu_slave_s0_readdatavalid;                   // afu_slave:s0_readdatavalid -> mm_interconnect_0:afu_slave_s0_readdatavalid
	wire         mm_interconnect_0_afu_slave_s0_write;                           // mm_interconnect_0:afu_slave_s0_write -> afu_slave:s0_write
	wire  [31:0] mm_interconnect_0_afu_slave_s0_writedata;                       // mm_interconnect_0:afu_slave_s0_writedata -> afu_slave:s0_writedata
	wire   [0:0] mm_interconnect_0_afu_slave_s0_burstcount;                      // mm_interconnect_0:afu_slave_s0_burstcount -> afu_slave:s0_burstcount
	wire  [63:0] mm_interconnect_0_bbs_slave_s0_readdata;                        // bbs_slave:s0_readdata -> mm_interconnect_0:bbs_slave_s0_readdata
	wire         mm_interconnect_0_bbs_slave_s0_waitrequest;                     // bbs_slave:s0_waitrequest -> mm_interconnect_0:bbs_slave_s0_waitrequest
	wire         mm_interconnect_0_bbs_slave_s0_debugaccess;                     // mm_interconnect_0:bbs_slave_s0_debugaccess -> bbs_slave:s0_debugaccess
	wire  [23:0] mm_interconnect_0_bbs_slave_s0_address;                         // mm_interconnect_0:bbs_slave_s0_address -> bbs_slave:s0_address
	wire         mm_interconnect_0_bbs_slave_s0_read;                            // mm_interconnect_0:bbs_slave_s0_read -> bbs_slave:s0_read
	wire   [7:0] mm_interconnect_0_bbs_slave_s0_byteenable;                      // mm_interconnect_0:bbs_slave_s0_byteenable -> bbs_slave:s0_byteenable
	wire         mm_interconnect_0_bbs_slave_s0_readdatavalid;                   // bbs_slave:s0_readdatavalid -> mm_interconnect_0:bbs_slave_s0_readdatavalid
	wire         mm_interconnect_0_bbs_slave_s0_write;                           // mm_interconnect_0:bbs_slave_s0_write -> bbs_slave:s0_write
	wire  [63:0] mm_interconnect_0_bbs_slave_s0_writedata;                       // mm_interconnect_0:bbs_slave_s0_writedata -> bbs_slave:s0_writedata
	wire   [0:0] mm_interconnect_0_bbs_slave_s0_burstcount;                      // mm_interconnect_0:bbs_slave_s0_burstcount -> bbs_slave:s0_burstcount
	wire  [31:0] mm_interconnect_0_cmb2avst_slave_s0_readdata;                   // cmb2avst_slave:s0_readdata -> mm_interconnect_0:cmb2avst_slave_s0_readdata
	wire         mm_interconnect_0_cmb2avst_slave_s0_waitrequest;                // cmb2avst_slave:s0_waitrequest -> mm_interconnect_0:cmb2avst_slave_s0_waitrequest
	wire         mm_interconnect_0_cmb2avst_slave_s0_debugaccess;                // mm_interconnect_0:cmb2avst_slave_s0_debugaccess -> cmb2avst_slave:s0_debugaccess
	wire  [23:0] mm_interconnect_0_cmb2avst_slave_s0_address;                    // mm_interconnect_0:cmb2avst_slave_s0_address -> cmb2avst_slave:s0_address
	wire         mm_interconnect_0_cmb2avst_slave_s0_read;                       // mm_interconnect_0:cmb2avst_slave_s0_read -> cmb2avst_slave:s0_read
	wire   [3:0] mm_interconnect_0_cmb2avst_slave_s0_byteenable;                 // mm_interconnect_0:cmb2avst_slave_s0_byteenable -> cmb2avst_slave:s0_byteenable
	wire         mm_interconnect_0_cmb2avst_slave_s0_readdatavalid;              // cmb2avst_slave:s0_readdatavalid -> mm_interconnect_0:cmb2avst_slave_s0_readdatavalid
	wire         mm_interconnect_0_cmb2avst_slave_s0_write;                      // mm_interconnect_0:cmb2avst_slave_s0_write -> cmb2avst_slave:s0_write
	wire  [31:0] mm_interconnect_0_cmb2avst_slave_s0_writedata;                  // mm_interconnect_0:cmb2avst_slave_s0_writedata -> cmb2avst_slave:s0_writedata
	wire   [0:0] mm_interconnect_0_cmb2avst_slave_s0_burstcount;                 // mm_interconnect_0:cmb2avst_slave_s0_burstcount -> cmb2avst_slave:s0_burstcount
	wire  [63:0] mm_interconnect_0_cxl_compliance_slave_s0_readdata;             // cxl_compliance_slave:s0_readdata -> mm_interconnect_0:cxl_compliance_slave_s0_readdata
	wire         mm_interconnect_0_cxl_compliance_slave_s0_waitrequest;          // cxl_compliance_slave:s0_waitrequest -> mm_interconnect_0:cxl_compliance_slave_s0_waitrequest
	wire         mm_interconnect_0_cxl_compliance_slave_s0_debugaccess;          // mm_interconnect_0:cxl_compliance_slave_s0_debugaccess -> cxl_compliance_slave:s0_debugaccess
	wire  [23:0] mm_interconnect_0_cxl_compliance_slave_s0_address;              // mm_interconnect_0:cxl_compliance_slave_s0_address -> cxl_compliance_slave:s0_address
	wire         mm_interconnect_0_cxl_compliance_slave_s0_read;                 // mm_interconnect_0:cxl_compliance_slave_s0_read -> cxl_compliance_slave:s0_read
	wire   [7:0] mm_interconnect_0_cxl_compliance_slave_s0_byteenable;           // mm_interconnect_0:cxl_compliance_slave_s0_byteenable -> cxl_compliance_slave:s0_byteenable
	wire         mm_interconnect_0_cxl_compliance_slave_s0_readdatavalid;        // cxl_compliance_slave:s0_readdatavalid -> mm_interconnect_0:cxl_compliance_slave_s0_readdatavalid
	wire         mm_interconnect_0_cxl_compliance_slave_s0_write;                // mm_interconnect_0:cxl_compliance_slave_s0_write -> cxl_compliance_slave:s0_write
	wire  [63:0] mm_interconnect_0_cxl_compliance_slave_s0_writedata;            // mm_interconnect_0:cxl_compliance_slave_s0_writedata -> cxl_compliance_slave:s0_writedata
	wire   [0:0] mm_interconnect_0_cxl_compliance_slave_s0_burstcount;           // mm_interconnect_0:cxl_compliance_slave_s0_burstcount -> cxl_compliance_slave:s0_burstcount
	wire  [31:0] mm_interconnect_0_cxl_io_csb2wire_csr_s0_readdata;              // cxl_io_csb2wire_csr:s0_readdata -> mm_interconnect_0:cxl_io_csb2wire_csr_s0_readdata
	wire         mm_interconnect_0_cxl_io_csb2wire_csr_s0_waitrequest;           // cxl_io_csb2wire_csr:s0_waitrequest -> mm_interconnect_0:cxl_io_csb2wire_csr_s0_waitrequest
	wire         mm_interconnect_0_cxl_io_csb2wire_csr_s0_debugaccess;           // mm_interconnect_0:cxl_io_csb2wire_csr_s0_debugaccess -> cxl_io_csb2wire_csr:s0_debugaccess
	wire  [23:0] mm_interconnect_0_cxl_io_csb2wire_csr_s0_address;               // mm_interconnect_0:cxl_io_csb2wire_csr_s0_address -> cxl_io_csb2wire_csr:s0_address
	wire         mm_interconnect_0_cxl_io_csb2wire_csr_s0_read;                  // mm_interconnect_0:cxl_io_csb2wire_csr_s0_read -> cxl_io_csb2wire_csr:s0_read
	wire   [3:0] mm_interconnect_0_cxl_io_csb2wire_csr_s0_byteenable;            // mm_interconnect_0:cxl_io_csb2wire_csr_s0_byteenable -> cxl_io_csb2wire_csr:s0_byteenable
	wire         mm_interconnect_0_cxl_io_csb2wire_csr_s0_readdatavalid;         // cxl_io_csb2wire_csr:s0_readdatavalid -> mm_interconnect_0:cxl_io_csb2wire_csr_s0_readdatavalid
	wire         mm_interconnect_0_cxl_io_csb2wire_csr_s0_write;                 // mm_interconnect_0:cxl_io_csb2wire_csr_s0_write -> cxl_io_csb2wire_csr:s0_write
	wire  [31:0] mm_interconnect_0_cxl_io_csb2wire_csr_s0_writedata;             // mm_interconnect_0:cxl_io_csb2wire_csr_s0_writedata -> cxl_io_csb2wire_csr:s0_writedata
	wire   [0:0] mm_interconnect_0_cxl_io_csb2wire_csr_s0_burstcount;            // mm_interconnect_0:cxl_io_csb2wire_csr_s0_burstcount -> cxl_io_csb2wire_csr:s0_burstcount
	wire  [31:0] mm_interconnect_0_cxl_io_slave_s0_readdata;                     // cxl_io_slave:s0_readdata -> mm_interconnect_0:cxl_io_slave_s0_readdata
	wire         mm_interconnect_0_cxl_io_slave_s0_waitrequest;                  // cxl_io_slave:s0_waitrequest -> mm_interconnect_0:cxl_io_slave_s0_waitrequest
	wire         mm_interconnect_0_cxl_io_slave_s0_debugaccess;                  // mm_interconnect_0:cxl_io_slave_s0_debugaccess -> cxl_io_slave:s0_debugaccess
	wire  [23:0] mm_interconnect_0_cxl_io_slave_s0_address;                      // mm_interconnect_0:cxl_io_slave_s0_address -> cxl_io_slave:s0_address
	wire         mm_interconnect_0_cxl_io_slave_s0_read;                         // mm_interconnect_0:cxl_io_slave_s0_read -> cxl_io_slave:s0_read
	wire   [3:0] mm_interconnect_0_cxl_io_slave_s0_byteenable;                   // mm_interconnect_0:cxl_io_slave_s0_byteenable -> cxl_io_slave:s0_byteenable
	wire         mm_interconnect_0_cxl_io_slave_s0_readdatavalid;                // cxl_io_slave:s0_readdatavalid -> mm_interconnect_0:cxl_io_slave_s0_readdatavalid
	wire         mm_interconnect_0_cxl_io_slave_s0_write;                        // mm_interconnect_0:cxl_io_slave_s0_write -> cxl_io_slave:s0_write
	wire  [31:0] mm_interconnect_0_cxl_io_slave_s0_writedata;                    // mm_interconnect_0:cxl_io_slave_s0_writedata -> cxl_io_slave:s0_writedata
	wire   [0:0] mm_interconnect_0_cxl_io_slave_s0_burstcount;                   // mm_interconnect_0:cxl_io_slave_s0_burstcount -> cxl_io_slave:s0_burstcount
	wire   [7:0] mm_interconnect_0_hip_reconfig_slave_s0_readdata;               // hip_reconfig_slave:s0_readdata -> mm_interconnect_0:hip_reconfig_slave_s0_readdata
	wire         mm_interconnect_0_hip_reconfig_slave_s0_waitrequest;            // hip_reconfig_slave:s0_waitrequest -> mm_interconnect_0:hip_reconfig_slave_s0_waitrequest
	wire         mm_interconnect_0_hip_reconfig_slave_s0_debugaccess;            // mm_interconnect_0:hip_reconfig_slave_s0_debugaccess -> hip_reconfig_slave:s0_debugaccess
	wire  [23:0] mm_interconnect_0_hip_reconfig_slave_s0_address;                // mm_interconnect_0:hip_reconfig_slave_s0_address -> hip_reconfig_slave:s0_address
	wire         mm_interconnect_0_hip_reconfig_slave_s0_read;                   // mm_interconnect_0:hip_reconfig_slave_s0_read -> hip_reconfig_slave:s0_read
	wire   [0:0] mm_interconnect_0_hip_reconfig_slave_s0_byteenable;             // mm_interconnect_0:hip_reconfig_slave_s0_byteenable -> hip_reconfig_slave:s0_byteenable
	wire         mm_interconnect_0_hip_reconfig_slave_s0_readdatavalid;          // hip_reconfig_slave:s0_readdatavalid -> mm_interconnect_0:hip_reconfig_slave_s0_readdatavalid
	wire         mm_interconnect_0_hip_reconfig_slave_s0_write;                  // mm_interconnect_0:hip_reconfig_slave_s0_write -> hip_reconfig_slave:s0_write
	wire   [7:0] mm_interconnect_0_hip_reconfig_slave_s0_writedata;              // mm_interconnect_0:hip_reconfig_slave_s0_writedata -> hip_reconfig_slave:s0_writedata
	wire   [0:0] mm_interconnect_0_hip_reconfig_slave_s0_burstcount;             // mm_interconnect_0:hip_reconfig_slave_s0_burstcount -> hip_reconfig_slave:s0_burstcount
	wire   [7:0] mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_readdata;      // usr_avmm_hip_reconfig_slave:s0_readdata -> mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_readdata
	wire         mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_waitrequest;   // usr_avmm_hip_reconfig_slave:s0_waitrequest -> mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_waitrequest
	wire         mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_debugaccess;   // mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_debugaccess -> usr_avmm_hip_reconfig_slave:s0_debugaccess
	wire  [23:0] mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_address;       // mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_address -> usr_avmm_hip_reconfig_slave:s0_address
	wire         mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_read;          // mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_read -> usr_avmm_hip_reconfig_slave:s0_read
	wire   [0:0] mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_byteenable;    // mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_byteenable -> usr_avmm_hip_reconfig_slave:s0_byteenable
	wire         mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_readdatavalid; // usr_avmm_hip_reconfig_slave:s0_readdatavalid -> mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_readdatavalid
	wire         mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_write;         // mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_write -> usr_avmm_hip_reconfig_slave:s0_write
	wire   [7:0] mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_writedata;     // mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_writedata -> usr_avmm_hip_reconfig_slave:s0_writedata
	wire   [0:0] mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_burstcount;    // mm_interconnect_0:usr_avmm_hip_reconfig_slave_s0_burstcount -> usr_avmm_hip_reconfig_slave:s0_burstcount

	afu_slave afu_slave (
		.clk              (interconnect_clock_in_out_clk_clk),            //   input,   width = 1,   clk.clk
		.reset            (~interconnect_reset_in_out_reset_reset),       //   input,   width = 1, reset.reset
		.s0_waitrequest   (mm_interconnect_0_afu_slave_s0_waitrequest),   //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_afu_slave_s0_readdata),      //  output,  width = 32,      .readdata
		.s0_readdatavalid (mm_interconnect_0_afu_slave_s0_readdatavalid), //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_afu_slave_s0_burstcount),    //   input,   width = 1,      .burstcount
		.s0_writedata     (mm_interconnect_0_afu_slave_s0_writedata),     //   input,  width = 32,      .writedata
		.s0_address       (mm_interconnect_0_afu_slave_s0_address),       //   input,  width = 24,      .address
		.s0_write         (mm_interconnect_0_afu_slave_s0_write),         //   input,   width = 1,      .write
		.s0_read          (mm_interconnect_0_afu_slave_s0_read),          //   input,   width = 1,      .read
		.s0_byteenable    (mm_interconnect_0_afu_slave_s0_byteenable),    //   input,   width = 4,      .byteenable
		.s0_debugaccess   (mm_interconnect_0_afu_slave_s0_debugaccess),   //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (afu_slave_m0_waitrequest),                     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (afu_slave_m0_readdata),                        //   input,  width = 32,      .readdata
		.m0_readdatavalid (afu_slave_m0_readdatavalid),                   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (afu_slave_m0_burstcount),                      //  output,   width = 1,      .burstcount
		.m0_writedata     (afu_slave_m0_writedata),                       //  output,  width = 32,      .writedata
		.m0_address       (afu_slave_m0_address),                         //  output,  width = 24,      .address
		.m0_write         (afu_slave_m0_write),                           //  output,   width = 1,      .write
		.m0_read          (afu_slave_m0_read),                            //  output,   width = 1,      .read
		.m0_byteenable    (afu_slave_m0_byteenable),                      //  output,   width = 4,      .byteenable
		.m0_debugaccess   (afu_slave_m0_debugaccess)                      //  output,   width = 1,      .debugaccess
	);

	bbs_slave bbs_slave (
		.clk              (interconnect_clock_in_out_clk_clk),            //   input,   width = 1,   clk.clk
		.reset            (~interconnect_reset_in_out_reset_reset),       //   input,   width = 1, reset.reset
		.s0_waitrequest   (mm_interconnect_0_bbs_slave_s0_waitrequest),   //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_bbs_slave_s0_readdata),      //  output,  width = 64,      .readdata
		.s0_readdatavalid (mm_interconnect_0_bbs_slave_s0_readdatavalid), //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_bbs_slave_s0_burstcount),    //   input,   width = 1,      .burstcount
		.s0_writedata     (mm_interconnect_0_bbs_slave_s0_writedata),     //   input,  width = 64,      .writedata
		.s0_address       (mm_interconnect_0_bbs_slave_s0_address),       //   input,  width = 24,      .address
		.s0_write         (mm_interconnect_0_bbs_slave_s0_write),         //   input,   width = 1,      .write
		.s0_read          (mm_interconnect_0_bbs_slave_s0_read),          //   input,   width = 1,      .read
		.s0_byteenable    (mm_interconnect_0_bbs_slave_s0_byteenable),    //   input,   width = 8,      .byteenable
		.s0_debugaccess   (mm_interconnect_0_bbs_slave_s0_debugaccess),   //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (bbs_slave_m0_waitrequest),                     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (bbs_slave_m0_readdata),                        //   input,  width = 64,      .readdata
		.m0_readdatavalid (bbs_slave_m0_readdatavalid),                   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (bbs_slave_m0_burstcount),                      //  output,   width = 1,      .burstcount
		.m0_writedata     (bbs_slave_m0_writedata),                       //  output,  width = 64,      .writedata
		.m0_address       (bbs_slave_m0_address),                         //  output,  width = 24,      .address
		.m0_write         (bbs_slave_m0_write),                           //  output,   width = 1,      .write
		.m0_read          (bbs_slave_m0_read),                            //  output,   width = 1,      .read
		.m0_byteenable    (bbs_slave_m0_byteenable),                      //  output,   width = 8,      .byteenable
		.m0_debugaccess   (bbs_slave_m0_debugaccess)                      //  output,   width = 1,      .debugaccess
	);

	cmb2avst_slave cmb2avst_slave (
		.clk              (interconnect_clock_in_out_clk_clk),                 //   input,   width = 1,   clk.clk
		.reset            (~interconnect_reset_in_out_reset_reset),            //   input,   width = 1, reset.reset
		.s0_waitrequest   (mm_interconnect_0_cmb2avst_slave_s0_waitrequest),   //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_cmb2avst_slave_s0_readdata),      //  output,  width = 32,      .readdata
		.s0_readdatavalid (mm_interconnect_0_cmb2avst_slave_s0_readdatavalid), //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_cmb2avst_slave_s0_burstcount),    //   input,   width = 1,      .burstcount
		.s0_writedata     (mm_interconnect_0_cmb2avst_slave_s0_writedata),     //   input,  width = 32,      .writedata
		.s0_address       (mm_interconnect_0_cmb2avst_slave_s0_address),       //   input,  width = 24,      .address
		.s0_write         (mm_interconnect_0_cmb2avst_slave_s0_write),         //   input,   width = 1,      .write
		.s0_read          (mm_interconnect_0_cmb2avst_slave_s0_read),          //   input,   width = 1,      .read
		.s0_byteenable    (mm_interconnect_0_cmb2avst_slave_s0_byteenable),    //   input,   width = 4,      .byteenable
		.s0_debugaccess   (mm_interconnect_0_cmb2avst_slave_s0_debugaccess),   //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (cmb2avst_slave_m0_waitrequest),                     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (cmb2avst_slave_m0_readdata),                        //   input,  width = 32,      .readdata
		.m0_readdatavalid (cmb2avst_slave_m0_readdatavalid),                   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (cmb2avst_slave_m0_burstcount),                      //  output,   width = 1,      .burstcount
		.m0_writedata     (cmb2avst_slave_m0_writedata),                       //  output,  width = 32,      .writedata
		.m0_address       (cmb2avst_slave_m0_address),                         //  output,  width = 24,      .address
		.m0_write         (cmb2avst_slave_m0_write),                           //  output,   width = 1,      .write
		.m0_read          (cmb2avst_slave_m0_read),                            //  output,   width = 1,      .read
		.m0_byteenable    (cmb2avst_slave_m0_byteenable),                      //  output,   width = 4,      .byteenable
		.m0_debugaccess   (cmb2avst_slave_m0_debugaccess)                      //  output,   width = 1,      .debugaccess
	);

	cxl_compliance_slave cxl_compliance_slave (
		.clk              (interconnect_clock_in_out_clk_clk),                       //   input,   width = 1,   clk.clk
		.reset            (~interconnect_reset_in_out_reset_reset),                  //   input,   width = 1, reset.reset
		.s0_waitrequest   (mm_interconnect_0_cxl_compliance_slave_s0_waitrequest),   //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_cxl_compliance_slave_s0_readdata),      //  output,  width = 64,      .readdata
		.s0_readdatavalid (mm_interconnect_0_cxl_compliance_slave_s0_readdatavalid), //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_cxl_compliance_slave_s0_burstcount),    //   input,   width = 1,      .burstcount
		.s0_writedata     (mm_interconnect_0_cxl_compliance_slave_s0_writedata),     //   input,  width = 64,      .writedata
		.s0_address       (mm_interconnect_0_cxl_compliance_slave_s0_address),       //   input,  width = 24,      .address
		.s0_write         (mm_interconnect_0_cxl_compliance_slave_s0_write),         //   input,   width = 1,      .write
		.s0_read          (mm_interconnect_0_cxl_compliance_slave_s0_read),          //   input,   width = 1,      .read
		.s0_byteenable    (mm_interconnect_0_cxl_compliance_slave_s0_byteenable),    //   input,   width = 8,      .byteenable
		.s0_debugaccess   (mm_interconnect_0_cxl_compliance_slave_s0_debugaccess),   //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (cxl_compliance_slave_m0_waitrequest),                     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (cxl_compliance_slave_m0_readdata),                        //   input,  width = 64,      .readdata
		.m0_readdatavalid (cxl_compliance_slave_m0_readdatavalid),                   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (cxl_compliance_slave_m0_burstcount),                      //  output,   width = 1,      .burstcount
		.m0_writedata     (cxl_compliance_slave_m0_writedata),                       //  output,  width = 64,      .writedata
		.m0_address       (cxl_compliance_slave_m0_address),                         //  output,  width = 24,      .address
		.m0_write         (cxl_compliance_slave_m0_write),                           //  output,   width = 1,      .write
		.m0_read          (cxl_compliance_slave_m0_read),                            //  output,   width = 1,      .read
		.m0_byteenable    (cxl_compliance_slave_m0_byteenable),                      //  output,   width = 8,      .byteenable
		.m0_debugaccess   (cxl_compliance_slave_m0_debugaccess)                      //  output,   width = 1,      .debugaccess
	);

	cxl_io_csb2wire_csr cxl_io_csb2wire_csr (
		.clk              (interconnect_clock_in_out_clk_clk),                      //   input,   width = 1,   clk.clk
		.reset            (~interconnect_reset_in_out_reset_reset),                 //   input,   width = 1, reset.reset
		.s0_waitrequest   (mm_interconnect_0_cxl_io_csb2wire_csr_s0_waitrequest),   //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_cxl_io_csb2wire_csr_s0_readdata),      //  output,  width = 32,      .readdata
		.s0_readdatavalid (mm_interconnect_0_cxl_io_csb2wire_csr_s0_readdatavalid), //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_cxl_io_csb2wire_csr_s0_burstcount),    //   input,   width = 1,      .burstcount
		.s0_writedata     (mm_interconnect_0_cxl_io_csb2wire_csr_s0_writedata),     //   input,  width = 32,      .writedata
		.s0_address       (mm_interconnect_0_cxl_io_csb2wire_csr_s0_address),       //   input,  width = 24,      .address
		.s0_write         (mm_interconnect_0_cxl_io_csb2wire_csr_s0_write),         //   input,   width = 1,      .write
		.s0_read          (mm_interconnect_0_cxl_io_csb2wire_csr_s0_read),          //   input,   width = 1,      .read
		.s0_byteenable    (mm_interconnect_0_cxl_io_csb2wire_csr_s0_byteenable),    //   input,   width = 4,      .byteenable
		.s0_debugaccess   (mm_interconnect_0_cxl_io_csb2wire_csr_s0_debugaccess),   //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (cxl_io_csb2wire_csr_m0_waitrequest),                     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (cxl_io_csb2wire_csr_m0_readdata),                        //   input,  width = 32,      .readdata
		.m0_readdatavalid (cxl_io_csb2wire_csr_m0_readdatavalid),                   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (cxl_io_csb2wire_csr_m0_burstcount),                      //  output,   width = 1,      .burstcount
		.m0_writedata     (cxl_io_csb2wire_csr_m0_writedata),                       //  output,  width = 32,      .writedata
		.m0_address       (cxl_io_csb2wire_csr_m0_address),                         //  output,  width = 24,      .address
		.m0_write         (cxl_io_csb2wire_csr_m0_write),                           //  output,   width = 1,      .write
		.m0_read          (cxl_io_csb2wire_csr_m0_read),                            //  output,   width = 1,      .read
		.m0_byteenable    (cxl_io_csb2wire_csr_m0_byteenable),                      //  output,   width = 4,      .byteenable
		.m0_debugaccess   (cxl_io_csb2wire_csr_m0_debugaccess)                      //  output,   width = 1,      .debugaccess
	);

	cxl_io_interconnect_clock cxl_io_interconnect_clock_in (
		.in_clk  (cxl_io_clk_clk),                           //   input,  width = 1,  in_clk.clk
		.out_clk (cxl_io_interconnect_clock_in_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	cxl_io_interconnect_reset cxl_io_interconnect_reset_in (
		.clk         (cxl_io_interconnect_clock_in_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (cxl_io_rst_reset_n),                           //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (cxl_io_interconnect_reset_in_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	cxl_io_master cxl_io_master (
		.m0_clk           (interconnect_clock_in_out_clk_clk),             //   input,   width = 1,   m0_clk.clk
		.m0_reset         (~interconnect_reset_in_out_reset_reset),        //   input,   width = 1, m0_reset.reset
		.s0_clk           (cxl_io_interconnect_clock_in_out_clk_clk),      //   input,   width = 1,   s0_clk.clk
		.s0_reset         (~cxl_io_interconnect_reset_in_out_reset_reset), //   input,   width = 1, s0_reset.reset
		.s0_waitrequest   (cxl_io_master_s0_waitrequest),                  //  output,   width = 1,       s0.waitrequest
		.s0_readdata      (cxl_io_master_s0_readdata),                     //  output,  width = 64,         .readdata
		.s0_readdatavalid (cxl_io_master_s0_readdatavalid),                //  output,   width = 1,         .readdatavalid
		.s0_burstcount    (cxl_io_master_s0_burstcount),                   //   input,   width = 1,         .burstcount
		.s0_writedata     (cxl_io_master_s0_writedata),                    //   input,  width = 64,         .writedata
		.s0_address       (cxl_io_master_s0_address),                      //   input,  width = 32,         .address
		.s0_write         (cxl_io_master_s0_write),                        //   input,   width = 1,         .write
		.s0_read          (cxl_io_master_s0_read),                         //   input,   width = 1,         .read
		.s0_byteenable    (cxl_io_master_s0_byteenable),                   //   input,   width = 8,         .byteenable
		.s0_debugaccess   (cxl_io_master_s0_debugaccess),                  //   input,   width = 1,         .debugaccess
		.m0_waitrequest   (cxl_io_master_m0_waitrequest),                  //   input,   width = 1,       m0.waitrequest
		.m0_readdata      (cxl_io_master_m0_readdata),                     //   input,  width = 64,         .readdata
		.m0_readdatavalid (cxl_io_master_m0_readdatavalid),                //   input,   width = 1,         .readdatavalid
		.m0_burstcount    (cxl_io_master_m0_burstcount),                   //  output,   width = 1,         .burstcount
		.m0_writedata     (cxl_io_master_m0_writedata),                    //  output,  width = 64,         .writedata
		.m0_address       (cxl_io_master_m0_address),                      //  output,  width = 32,         .address
		.m0_write         (cxl_io_master_m0_write),                        //  output,   width = 1,         .write
		.m0_read          (cxl_io_master_m0_read),                         //  output,   width = 1,         .read
		.m0_byteenable    (cxl_io_master_m0_byteenable),                   //  output,   width = 8,         .byteenable
		.m0_debugaccess   (cxl_io_master_m0_debugaccess)                   //  output,   width = 1,         .debugaccess
	);

	cxl_io_slave cxl_io_slave (
		.m0_clk           (cxl_io_interconnect_clock_in_out_clk_clk),        //   input,   width = 1,   m0_clk.clk
		.m0_reset         (~cxl_io_interconnect_reset_in_out_reset_reset),   //   input,   width = 1, m0_reset.reset
		.s0_clk           (interconnect_clock_in_out_clk_clk),               //   input,   width = 1,   s0_clk.clk
		.s0_reset         (~interconnect_reset_in_out_reset_reset),          //   input,   width = 1, s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_cxl_io_slave_s0_waitrequest),   //  output,   width = 1,       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_cxl_io_slave_s0_readdata),      //  output,  width = 32,         .readdata
		.s0_readdatavalid (mm_interconnect_0_cxl_io_slave_s0_readdatavalid), //  output,   width = 1,         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_cxl_io_slave_s0_burstcount),    //   input,   width = 1,         .burstcount
		.s0_writedata     (mm_interconnect_0_cxl_io_slave_s0_writedata),     //   input,  width = 32,         .writedata
		.s0_address       (mm_interconnect_0_cxl_io_slave_s0_address),       //   input,  width = 24,         .address
		.s0_write         (mm_interconnect_0_cxl_io_slave_s0_write),         //   input,   width = 1,         .write
		.s0_read          (mm_interconnect_0_cxl_io_slave_s0_read),          //   input,   width = 1,         .read
		.s0_byteenable    (mm_interconnect_0_cxl_io_slave_s0_byteenable),    //   input,   width = 4,         .byteenable
		.s0_debugaccess   (mm_interconnect_0_cxl_io_slave_s0_debugaccess),   //   input,   width = 1,         .debugaccess
		.m0_waitrequest   (cxl_io_slave_m0_waitrequest),                     //   input,   width = 1,       m0.waitrequest
		.m0_readdata      (cxl_io_slave_m0_readdata),                        //   input,  width = 32,         .readdata
		.m0_readdatavalid (cxl_io_slave_m0_readdatavalid),                   //   input,   width = 1,         .readdatavalid
		.m0_burstcount    (cxl_io_slave_m0_burstcount),                      //  output,   width = 1,         .burstcount
		.m0_writedata     (cxl_io_slave_m0_writedata),                       //  output,  width = 32,         .writedata
		.m0_address       (cxl_io_slave_m0_address),                         //  output,  width = 24,         .address
		.m0_write         (cxl_io_slave_m0_write),                           //  output,   width = 1,         .write
		.m0_read          (cxl_io_slave_m0_read),                            //  output,   width = 1,         .read
		.m0_byteenable    (cxl_io_slave_m0_byteenable),                      //  output,   width = 4,         .byteenable
		.m0_debugaccess   (cxl_io_slave_m0_debugaccess)                      //  output,   width = 1,         .debugaccess
	);

	debug_master debug_master (
		.clk              (interconnect_clock_in_out_clk_clk),      //   input,   width = 1,   clk.clk
		.reset            (~interconnect_reset_in_out_reset_reset), //   input,   width = 1, reset.reset
		.s0_waitrequest   (debug_master_s0_waitrequest),            //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (debug_master_s0_readdata),               //  output,  width = 32,      .readdata
		.s0_readdatavalid (debug_master_s0_readdatavalid),          //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (debug_master_s0_burstcount),             //   input,   width = 1,      .burstcount
		.s0_writedata     (debug_master_s0_writedata),              //   input,  width = 32,      .writedata
		.s0_address       (debug_master_s0_address),                //   input,  width = 32,      .address
		.s0_write         (debug_master_s0_write),                  //   input,   width = 1,      .write
		.s0_read          (debug_master_s0_read),                   //   input,   width = 1,      .read
		.s0_byteenable    (debug_master_s0_byteenable),             //   input,   width = 4,      .byteenable
		.s0_debugaccess   (debug_master_s0_debugaccess),            //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (debug_master_m0_waitrequest),            //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (debug_master_m0_readdata),               //   input,  width = 32,      .readdata
		.m0_readdatavalid (debug_master_m0_readdatavalid),          //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (debug_master_m0_burstcount),             //  output,   width = 1,      .burstcount
		.m0_writedata     (debug_master_m0_writedata),              //  output,  width = 32,      .writedata
		.m0_address       (debug_master_m0_address),                //  output,  width = 32,      .address
		.m0_write         (debug_master_m0_write),                  //  output,   width = 1,      .write
		.m0_read          (debug_master_m0_read),                   //  output,   width = 1,      .read
		.m0_byteenable    (debug_master_m0_byteenable),             //  output,   width = 4,      .byteenable
		.m0_debugaccess   (debug_master_m0_debugaccess)             //  output,   width = 1,      .debugaccess
	);

	hip_reconfig_clock_in hip_reconfig_clock_in (
		.in_clk  (side_clock_hip_clk),                //   input,  width = 1,  in_clk.clk
		.out_clk (hip_reconfig_clock_in_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	hip_reconfig_reset_in hip_reconfig_reset_in (
		.clk         (hip_reconfig_clock_in_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (side_reset_hip_reset_n),                //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (hip_reconfig_reset_in_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	hip_reconfig_slave hip_reconfig_slave (
		.m0_clk           (hip_reconfig_clock_in_out_clk_clk),                     //   input,   width = 1,   m0_clk.clk
		.m0_reset         (~hip_reconfig_reset_in_out_reset_reset),                //   input,   width = 1, m0_reset.reset
		.s0_clk           (interconnect_clock_in_out_clk_clk),                     //   input,   width = 1,   s0_clk.clk
		.s0_reset         (~interconnect_reset_in_out_reset_reset),                //   input,   width = 1, s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_hip_reconfig_slave_s0_waitrequest),   //  output,   width = 1,       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_hip_reconfig_slave_s0_readdata),      //  output,   width = 8,         .readdata
		.s0_readdatavalid (mm_interconnect_0_hip_reconfig_slave_s0_readdatavalid), //  output,   width = 1,         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_hip_reconfig_slave_s0_burstcount),    //   input,   width = 1,         .burstcount
		.s0_writedata     (mm_interconnect_0_hip_reconfig_slave_s0_writedata),     //   input,   width = 8,         .writedata
		.s0_address       (mm_interconnect_0_hip_reconfig_slave_s0_address),       //   input,  width = 24,         .address
		.s0_write         (mm_interconnect_0_hip_reconfig_slave_s0_write),         //   input,   width = 1,         .write
		.s0_read          (mm_interconnect_0_hip_reconfig_slave_s0_read),          //   input,   width = 1,         .read
		.s0_byteenable    (mm_interconnect_0_hip_reconfig_slave_s0_byteenable),    //   input,   width = 1,         .byteenable
		.s0_debugaccess   (mm_interconnect_0_hip_reconfig_slave_s0_debugaccess),   //   input,   width = 1,         .debugaccess
		.m0_waitrequest   (hip_reconfig_slave_m0_waitrequest),                     //   input,   width = 1,       m0.waitrequest
		.m0_readdata      (hip_reconfig_slave_m0_readdata),                        //   input,   width = 8,         .readdata
		.m0_readdatavalid (hip_reconfig_slave_m0_readdatavalid),                   //   input,   width = 1,         .readdatavalid
		.m0_burstcount    (hip_reconfig_slave_m0_burstcount),                      //  output,   width = 1,         .burstcount
		.m0_writedata     (hip_reconfig_slave_m0_writedata),                       //  output,   width = 8,         .writedata
		.m0_address       (hip_reconfig_slave_m0_address),                         //  output,  width = 24,         .address
		.m0_write         (hip_reconfig_slave_m0_write),                           //  output,   width = 1,         .write
		.m0_read          (hip_reconfig_slave_m0_read),                            //  output,   width = 1,         .read
		.m0_byteenable    (hip_reconfig_slave_m0_byteenable),                      //  output,   width = 1,         .byteenable
		.m0_debugaccess   (hip_reconfig_slave_m0_debugaccess)                      //  output,   width = 1,         .debugaccess
	);

	avmm_interconnect_clock_in interconnect_clock_in (
		.in_clk  (int_conn_clk_clk),                  //   input,  width = 1,  in_clk.clk
		.out_clk (interconnect_clock_in_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	avmm_interconnect_reset_in interconnect_reset_in (
		.clk         (interconnect_clock_in_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (int_conn_rst_reset_n),                  //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (interconnect_reset_in_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	usr_avmm_hip_reconfig_slave usr_avmm_hip_reconfig_slave (
		.clk              (interconnect_clock_in_out_clk_clk),                              //   input,   width = 1,   clk.clk
		.reset            (~interconnect_reset_in_out_reset_reset),                         //   input,   width = 1, reset.reset
		.s0_waitrequest   (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_waitrequest),   //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_readdata),      //  output,   width = 8,      .readdata
		.s0_readdatavalid (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_readdatavalid), //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_burstcount),    //   input,   width = 1,      .burstcount
		.s0_writedata     (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_writedata),     //   input,   width = 8,      .writedata
		.s0_address       (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_address),       //   input,  width = 24,      .address
		.s0_write         (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_write),         //   input,   width = 1,      .write
		.s0_read          (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_read),          //   input,   width = 1,      .read
		.s0_byteenable    (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_byteenable),    //   input,   width = 1,      .byteenable
		.s0_debugaccess   (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_debugaccess),   //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (usr_avmm_hip_reconfig_slave_m0_waitrequest),                     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (usr_avmm_hip_reconfig_slave_m0_readdata),                        //   input,   width = 8,      .readdata
		.m0_readdatavalid (usr_avmm_hip_reconfig_slave_m0_readdatavalid),                   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (usr_avmm_hip_reconfig_slave_m0_burstcount),                      //  output,   width = 1,      .burstcount
		.m0_writedata     (usr_avmm_hip_reconfig_slave_m0_writedata),                       //  output,   width = 8,      .writedata
		.m0_address       (usr_avmm_hip_reconfig_slave_m0_address),                         //  output,  width = 24,      .address
		.m0_write         (usr_avmm_hip_reconfig_slave_m0_write),                           //  output,   width = 1,      .write
		.m0_read          (usr_avmm_hip_reconfig_slave_m0_read),                            //  output,   width = 1,      .read
		.m0_byteenable    (usr_avmm_hip_reconfig_slave_m0_byteenable),                      //  output,   width = 1,      .byteenable
		.m0_debugaccess   (usr_avmm_hip_reconfig_slave_m0_debugaccess)                      //  output,   width = 1,      .debugaccess
	);

	avmm_interconnect_altera_mm_interconnect_1920_x6i2ati mm_interconnect_0 (
		.cxl_io_master_m0_address                                          (cxl_io_master_m0_address),                                       //   input,  width = 32,                                            cxl_io_master_m0.address
		.cxl_io_master_m0_waitrequest                                      (cxl_io_master_m0_waitrequest),                                   //  output,   width = 1,                                                            .waitrequest
		.cxl_io_master_m0_burstcount                                       (cxl_io_master_m0_burstcount),                                    //   input,   width = 1,                                                            .burstcount
		.cxl_io_master_m0_byteenable                                       (cxl_io_master_m0_byteenable),                                    //   input,   width = 8,                                                            .byteenable
		.cxl_io_master_m0_read                                             (cxl_io_master_m0_read),                                          //   input,   width = 1,                                                            .read
		.cxl_io_master_m0_readdata                                         (cxl_io_master_m0_readdata),                                      //  output,  width = 64,                                                            .readdata
		.cxl_io_master_m0_readdatavalid                                    (cxl_io_master_m0_readdatavalid),                                 //  output,   width = 1,                                                            .readdatavalid
		.cxl_io_master_m0_write                                            (cxl_io_master_m0_write),                                         //   input,   width = 1,                                                            .write
		.cxl_io_master_m0_writedata                                        (cxl_io_master_m0_writedata),                                     //   input,  width = 64,                                                            .writedata
		.cxl_io_master_m0_debugaccess                                      (cxl_io_master_m0_debugaccess),                                   //   input,   width = 1,                                                            .debugaccess
		.debug_master_m0_address                                           (debug_master_m0_address),                                        //   input,  width = 32,                                             debug_master_m0.address
		.debug_master_m0_waitrequest                                       (debug_master_m0_waitrequest),                                    //  output,   width = 1,                                                            .waitrequest
		.debug_master_m0_burstcount                                        (debug_master_m0_burstcount),                                     //   input,   width = 1,                                                            .burstcount
		.debug_master_m0_byteenable                                        (debug_master_m0_byteenable),                                     //   input,   width = 4,                                                            .byteenable
		.debug_master_m0_read                                              (debug_master_m0_read),                                           //   input,   width = 1,                                                            .read
		.debug_master_m0_readdata                                          (debug_master_m0_readdata),                                       //  output,  width = 32,                                                            .readdata
		.debug_master_m0_readdatavalid                                     (debug_master_m0_readdatavalid),                                  //  output,   width = 1,                                                            .readdatavalid
		.debug_master_m0_write                                             (debug_master_m0_write),                                          //   input,   width = 1,                                                            .write
		.debug_master_m0_writedata                                         (debug_master_m0_writedata),                                      //   input,  width = 32,                                                            .writedata
		.debug_master_m0_debugaccess                                       (debug_master_m0_debugaccess),                                    //   input,   width = 1,                                                            .debugaccess
		.afu_slave_s0_address                                              (mm_interconnect_0_afu_slave_s0_address),                         //  output,  width = 24,                                                afu_slave_s0.address
		.afu_slave_s0_write                                                (mm_interconnect_0_afu_slave_s0_write),                           //  output,   width = 1,                                                            .write
		.afu_slave_s0_read                                                 (mm_interconnect_0_afu_slave_s0_read),                            //  output,   width = 1,                                                            .read
		.afu_slave_s0_readdata                                             (mm_interconnect_0_afu_slave_s0_readdata),                        //   input,  width = 32,                                                            .readdata
		.afu_slave_s0_writedata                                            (mm_interconnect_0_afu_slave_s0_writedata),                       //  output,  width = 32,                                                            .writedata
		.afu_slave_s0_burstcount                                           (mm_interconnect_0_afu_slave_s0_burstcount),                      //  output,   width = 1,                                                            .burstcount
		.afu_slave_s0_byteenable                                           (mm_interconnect_0_afu_slave_s0_byteenable),                      //  output,   width = 4,                                                            .byteenable
		.afu_slave_s0_readdatavalid                                        (mm_interconnect_0_afu_slave_s0_readdatavalid),                   //   input,   width = 1,                                                            .readdatavalid
		.afu_slave_s0_waitrequest                                          (mm_interconnect_0_afu_slave_s0_waitrequest),                     //   input,   width = 1,                                                            .waitrequest
		.afu_slave_s0_debugaccess                                          (mm_interconnect_0_afu_slave_s0_debugaccess),                     //  output,   width = 1,                                                            .debugaccess
		.bbs_slave_s0_address                                              (mm_interconnect_0_bbs_slave_s0_address),                         //  output,  width = 24,                                                bbs_slave_s0.address
		.bbs_slave_s0_write                                                (mm_interconnect_0_bbs_slave_s0_write),                           //  output,   width = 1,                                                            .write
		.bbs_slave_s0_read                                                 (mm_interconnect_0_bbs_slave_s0_read),                            //  output,   width = 1,                                                            .read
		.bbs_slave_s0_readdata                                             (mm_interconnect_0_bbs_slave_s0_readdata),                        //   input,  width = 64,                                                            .readdata
		.bbs_slave_s0_writedata                                            (mm_interconnect_0_bbs_slave_s0_writedata),                       //  output,  width = 64,                                                            .writedata
		.bbs_slave_s0_burstcount                                           (mm_interconnect_0_bbs_slave_s0_burstcount),                      //  output,   width = 1,                                                            .burstcount
		.bbs_slave_s0_byteenable                                           (mm_interconnect_0_bbs_slave_s0_byteenable),                      //  output,   width = 8,                                                            .byteenable
		.bbs_slave_s0_readdatavalid                                        (mm_interconnect_0_bbs_slave_s0_readdatavalid),                   //   input,   width = 1,                                                            .readdatavalid
		.bbs_slave_s0_waitrequest                                          (mm_interconnect_0_bbs_slave_s0_waitrequest),                     //   input,   width = 1,                                                            .waitrequest
		.bbs_slave_s0_debugaccess                                          (mm_interconnect_0_bbs_slave_s0_debugaccess),                     //  output,   width = 1,                                                            .debugaccess
		.cmb2avst_slave_s0_address                                         (mm_interconnect_0_cmb2avst_slave_s0_address),                    //  output,  width = 24,                                           cmb2avst_slave_s0.address
		.cmb2avst_slave_s0_write                                           (mm_interconnect_0_cmb2avst_slave_s0_write),                      //  output,   width = 1,                                                            .write
		.cmb2avst_slave_s0_read                                            (mm_interconnect_0_cmb2avst_slave_s0_read),                       //  output,   width = 1,                                                            .read
		.cmb2avst_slave_s0_readdata                                        (mm_interconnect_0_cmb2avst_slave_s0_readdata),                   //   input,  width = 32,                                                            .readdata
		.cmb2avst_slave_s0_writedata                                       (mm_interconnect_0_cmb2avst_slave_s0_writedata),                  //  output,  width = 32,                                                            .writedata
		.cmb2avst_slave_s0_burstcount                                      (mm_interconnect_0_cmb2avst_slave_s0_burstcount),                 //  output,   width = 1,                                                            .burstcount
		.cmb2avst_slave_s0_byteenable                                      (mm_interconnect_0_cmb2avst_slave_s0_byteenable),                 //  output,   width = 4,                                                            .byteenable
		.cmb2avst_slave_s0_readdatavalid                                   (mm_interconnect_0_cmb2avst_slave_s0_readdatavalid),              //   input,   width = 1,                                                            .readdatavalid
		.cmb2avst_slave_s0_waitrequest                                     (mm_interconnect_0_cmb2avst_slave_s0_waitrequest),                //   input,   width = 1,                                                            .waitrequest
		.cmb2avst_slave_s0_debugaccess                                     (mm_interconnect_0_cmb2avst_slave_s0_debugaccess),                //  output,   width = 1,                                                            .debugaccess
		.cxl_compliance_slave_s0_address                                   (mm_interconnect_0_cxl_compliance_slave_s0_address),              //  output,  width = 24,                                     cxl_compliance_slave_s0.address
		.cxl_compliance_slave_s0_write                                     (mm_interconnect_0_cxl_compliance_slave_s0_write),                //  output,   width = 1,                                                            .write
		.cxl_compliance_slave_s0_read                                      (mm_interconnect_0_cxl_compliance_slave_s0_read),                 //  output,   width = 1,                                                            .read
		.cxl_compliance_slave_s0_readdata                                  (mm_interconnect_0_cxl_compliance_slave_s0_readdata),             //   input,  width = 64,                                                            .readdata
		.cxl_compliance_slave_s0_writedata                                 (mm_interconnect_0_cxl_compliance_slave_s0_writedata),            //  output,  width = 64,                                                            .writedata
		.cxl_compliance_slave_s0_burstcount                                (mm_interconnect_0_cxl_compliance_slave_s0_burstcount),           //  output,   width = 1,                                                            .burstcount
		.cxl_compliance_slave_s0_byteenable                                (mm_interconnect_0_cxl_compliance_slave_s0_byteenable),           //  output,   width = 8,                                                            .byteenable
		.cxl_compliance_slave_s0_readdatavalid                             (mm_interconnect_0_cxl_compliance_slave_s0_readdatavalid),        //   input,   width = 1,                                                            .readdatavalid
		.cxl_compliance_slave_s0_waitrequest                               (mm_interconnect_0_cxl_compliance_slave_s0_waitrequest),          //   input,   width = 1,                                                            .waitrequest
		.cxl_compliance_slave_s0_debugaccess                               (mm_interconnect_0_cxl_compliance_slave_s0_debugaccess),          //  output,   width = 1,                                                            .debugaccess
		.cxl_io_csb2wire_csr_s0_address                                    (mm_interconnect_0_cxl_io_csb2wire_csr_s0_address),               //  output,  width = 24,                                      cxl_io_csb2wire_csr_s0.address
		.cxl_io_csb2wire_csr_s0_write                                      (mm_interconnect_0_cxl_io_csb2wire_csr_s0_write),                 //  output,   width = 1,                                                            .write
		.cxl_io_csb2wire_csr_s0_read                                       (mm_interconnect_0_cxl_io_csb2wire_csr_s0_read),                  //  output,   width = 1,                                                            .read
		.cxl_io_csb2wire_csr_s0_readdata                                   (mm_interconnect_0_cxl_io_csb2wire_csr_s0_readdata),              //   input,  width = 32,                                                            .readdata
		.cxl_io_csb2wire_csr_s0_writedata                                  (mm_interconnect_0_cxl_io_csb2wire_csr_s0_writedata),             //  output,  width = 32,                                                            .writedata
		.cxl_io_csb2wire_csr_s0_burstcount                                 (mm_interconnect_0_cxl_io_csb2wire_csr_s0_burstcount),            //  output,   width = 1,                                                            .burstcount
		.cxl_io_csb2wire_csr_s0_byteenable                                 (mm_interconnect_0_cxl_io_csb2wire_csr_s0_byteenable),            //  output,   width = 4,                                                            .byteenable
		.cxl_io_csb2wire_csr_s0_readdatavalid                              (mm_interconnect_0_cxl_io_csb2wire_csr_s0_readdatavalid),         //   input,   width = 1,                                                            .readdatavalid
		.cxl_io_csb2wire_csr_s0_waitrequest                                (mm_interconnect_0_cxl_io_csb2wire_csr_s0_waitrequest),           //   input,   width = 1,                                                            .waitrequest
		.cxl_io_csb2wire_csr_s0_debugaccess                                (mm_interconnect_0_cxl_io_csb2wire_csr_s0_debugaccess),           //  output,   width = 1,                                                            .debugaccess
		.cxl_io_slave_s0_address                                           (mm_interconnect_0_cxl_io_slave_s0_address),                      //  output,  width = 24,                                             cxl_io_slave_s0.address
		.cxl_io_slave_s0_write                                             (mm_interconnect_0_cxl_io_slave_s0_write),                        //  output,   width = 1,                                                            .write
		.cxl_io_slave_s0_read                                              (mm_interconnect_0_cxl_io_slave_s0_read),                         //  output,   width = 1,                                                            .read
		.cxl_io_slave_s0_readdata                                          (mm_interconnect_0_cxl_io_slave_s0_readdata),                     //   input,  width = 32,                                                            .readdata
		.cxl_io_slave_s0_writedata                                         (mm_interconnect_0_cxl_io_slave_s0_writedata),                    //  output,  width = 32,                                                            .writedata
		.cxl_io_slave_s0_burstcount                                        (mm_interconnect_0_cxl_io_slave_s0_burstcount),                   //  output,   width = 1,                                                            .burstcount
		.cxl_io_slave_s0_byteenable                                        (mm_interconnect_0_cxl_io_slave_s0_byteenable),                   //  output,   width = 4,                                                            .byteenable
		.cxl_io_slave_s0_readdatavalid                                     (mm_interconnect_0_cxl_io_slave_s0_readdatavalid),                //   input,   width = 1,                                                            .readdatavalid
		.cxl_io_slave_s0_waitrequest                                       (mm_interconnect_0_cxl_io_slave_s0_waitrequest),                  //   input,   width = 1,                                                            .waitrequest
		.cxl_io_slave_s0_debugaccess                                       (mm_interconnect_0_cxl_io_slave_s0_debugaccess),                  //  output,   width = 1,                                                            .debugaccess
		.hip_reconfig_slave_s0_address                                     (mm_interconnect_0_hip_reconfig_slave_s0_address),                //  output,  width = 24,                                       hip_reconfig_slave_s0.address
		.hip_reconfig_slave_s0_write                                       (mm_interconnect_0_hip_reconfig_slave_s0_write),                  //  output,   width = 1,                                                            .write
		.hip_reconfig_slave_s0_read                                        (mm_interconnect_0_hip_reconfig_slave_s0_read),                   //  output,   width = 1,                                                            .read
		.hip_reconfig_slave_s0_readdata                                    (mm_interconnect_0_hip_reconfig_slave_s0_readdata),               //   input,   width = 8,                                                            .readdata
		.hip_reconfig_slave_s0_writedata                                   (mm_interconnect_0_hip_reconfig_slave_s0_writedata),              //  output,   width = 8,                                                            .writedata
		.hip_reconfig_slave_s0_burstcount                                  (mm_interconnect_0_hip_reconfig_slave_s0_burstcount),             //  output,   width = 1,                                                            .burstcount
		.hip_reconfig_slave_s0_byteenable                                  (mm_interconnect_0_hip_reconfig_slave_s0_byteenable),             //  output,   width = 1,                                                            .byteenable
		.hip_reconfig_slave_s0_readdatavalid                               (mm_interconnect_0_hip_reconfig_slave_s0_readdatavalid),          //   input,   width = 1,                                                            .readdatavalid
		.hip_reconfig_slave_s0_waitrequest                                 (mm_interconnect_0_hip_reconfig_slave_s0_waitrequest),            //   input,   width = 1,                                                            .waitrequest
		.hip_reconfig_slave_s0_debugaccess                                 (mm_interconnect_0_hip_reconfig_slave_s0_debugaccess),            //  output,   width = 1,                                                            .debugaccess
		.usr_avmm_hip_reconfig_slave_s0_address                            (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_address),       //  output,  width = 24,                              usr_avmm_hip_reconfig_slave_s0.address
		.usr_avmm_hip_reconfig_slave_s0_write                              (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_write),         //  output,   width = 1,                                                            .write
		.usr_avmm_hip_reconfig_slave_s0_read                               (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_read),          //  output,   width = 1,                                                            .read
		.usr_avmm_hip_reconfig_slave_s0_readdata                           (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_readdata),      //   input,   width = 8,                                                            .readdata
		.usr_avmm_hip_reconfig_slave_s0_writedata                          (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_writedata),     //  output,   width = 8,                                                            .writedata
		.usr_avmm_hip_reconfig_slave_s0_burstcount                         (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_burstcount),    //  output,   width = 1,                                                            .burstcount
		.usr_avmm_hip_reconfig_slave_s0_byteenable                         (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_byteenable),    //  output,   width = 1,                                                            .byteenable
		.usr_avmm_hip_reconfig_slave_s0_readdatavalid                      (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_readdatavalid), //   input,   width = 1,                                                            .readdatavalid
		.usr_avmm_hip_reconfig_slave_s0_waitrequest                        (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_waitrequest),   //   input,   width = 1,                                                            .waitrequest
		.usr_avmm_hip_reconfig_slave_s0_debugaccess                        (mm_interconnect_0_usr_avmm_hip_reconfig_slave_s0_debugaccess),   //  output,   width = 1,                                                            .debugaccess
		.cxl_io_master_m0_reset_reset_bridge_in_reset_reset                (~interconnect_reset_in_out_reset_reset),                         //   input,   width = 1,                cxl_io_master_m0_reset_reset_bridge_in_reset.reset
		.afu_slave_s0_agent_rsp_fifo_clk_reset_reset_bridge_in_reset_reset (~interconnect_reset_in_out_reset_reset),                         //   input,   width = 1, afu_slave_s0_agent_rsp_fifo_clk_reset_reset_bridge_in_reset.reset
		.interconnect_clock_in_out_clk_clk                                 (interconnect_clock_in_out_clk_clk)                               //   input,   width = 1,                               interconnect_clock_in_out_clk.clk
	);

endmodule
