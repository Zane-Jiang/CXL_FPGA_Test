// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E4KnbZwe/6lSZ/ISRKvVD31nBUumqsriYvlq6ZEbMVmQq5/s5b3DdgOQwiDO
2rhJQoeYJDz5Ttp75chkeIhvDw4xoO0KRTrDS8jVlUR+EHZnfHh88BsFsn2y
mRHg4ck2tPz5P36apC1ZehfzEvWWPYdNGRG9mRZj+fxoybgsW4/s/UDq0u8s
umr41SZltvf5tTCXZZAY8IXeOmeVwYMUD9gfVPR+7TTgjLp7veAVFLCcW66+
btdS3EYP3vJNB36ru7MZo9iuqyDeVT53H4QeFFbTe/63VuVY0qSfVjXWfknh
ggV2XYsuoQvA+78yWd3x1IWpMvCrq59r91cef14riw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JtvMM1gj1WDpdH3VuQDmuoJ2x+HXXDa/vl1Wx7//Ag4b5VFghdSGah+GPRDB
nw3jZsqhFyAY13wac/16/LwL3/kDzU/RBg/gMcrL+m9K3KPhNdGCR5M2P7g5
TDKIKs+BqJvd3eqROTa04I1QbQA4RpSShmaTysB4koBTIUCAgDb4x+BVC6Ld
Vj7cVuqBp5BSsjg+lC5njTCbzIVvi6ejlb4KC2R8EAi3O/z/aLJPUewEVBFM
CKGCr6RBkMi4Uo9q6ujtPjbECzqoHYXLUipL+oEkq907TW+/Ttz9I2oWwAEo
jszRO3hvU6LMCFt1cB4TMohv2u5InZRDr7WkUiKGGw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Vkeg0AqbjK52AizoHHiFzY02lv7zfDdpl9esHVx4T7SxAiPC6K9MDuUwga34
D7rGKSU3rl0nL32bL5pd050vLh16n2wjjLwZQffQqRBZYQ8//g35grd0WP6J
kQXLsROsH0EFnp/5gT0IUzElvU8DG9sCqnOUFBaArj+lw6+T0FZmnTQITDOQ
u0Av551dbaEVDs3FJKtEXfuG74ZDKbm/NQ7Q/LKqPLBFmFgvaJddqvqwT8f+
f73QisiibMOTgS/58W6pEVsZ7BrXVnw4mY7tgg0uj9cHDbQTHMUh66/04axX
f25D0Hu2CIvIUgBSUfLZQFOa0Xn2CKSKeq/CJJWFVw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WEeZDTG/K+TLYpQly40ZNbS76dHfWvzriJ3dkuv5vLNcP5J+LwzqAOn+XJPW
E+FuWsWZV4wFisQDchxQX77nPwK/UwWLhZ4W5G/U1NR6p1pT+BJdMi06D4v3
pM01PG7fgg1G7M5ZnP/VyGteyw6bYhFP3JQUgplnaj+mnf/DvFw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
d1pX9T6rW0JyQfuM7LvzIwQ/fhZdsoJoAqqWmCmjetZQN1NV8BPDL60fmDNJ
S5SPK6Vd2VT93YRlflTzSBSNmZch/fVAymhlRV6fbelrTMgbWotrCbGBrGSz
SqfEOWi/phtxmJDu+9ylOYyRMuubstd5PcpYkme4Q+dAStBPr3YHouc5Zp2k
k/kZG3m6NGsQ1aF++O0/ntVjvPk2DRyrrUZCNV6ZEGKOacbdQ2D/D9UYrdYc
XL1gOq8bH3IFgrMF1KgfX3BgBeR000/Sby5fq8UGFmRGNnOSGaHMeq0cIRgn
7g9sslTgC4s41APqxGzIpEF9LF6TUVBf9dY6kC18sYfllvUQZqyBbJxDiHA1
/AaGLw5VPU+LTIRZHJaYTlgZlWjHUauIsnurlaUpP4a6CmwT/puF0ShPXYye
fNGGAu+Z6xiZLMZkhOAJYWIvipMtjuNzUeGRfKWf5h5AjJB8w6FBb4Wjtl/M
xxFiw5J1P2LX4q39ZaoMlvova/G2tRI+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Vzh+DN/3M0kiUXRMGIKOfpMqqNA8SnHnSRNI7iPdRg0G4KvooFSiL/KohKbf
fAwVnwqyDAVnO4coHqr8ty+Mj79OGtu5WUjVfT7yfKe3RleZN1/0M7y4ZYb8
PNFgAbdD71vxwltJ6ADIHgsoeuCqEcMlguXRT24RMgjpL8Loy0o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aoRiqicwXFt1HK/0+nFQGfZ0r9U0hAHh1PrvM/+uOtt2IjS3xDW7uZQhiNDI
UJxFI8zK2TqSXgxJBdbaqKPB3ffR3IsDXqRq88BzjZzK/SpXjvjSFoIfvcic
9Zpf3eaqV8gWV6m0wDOY1OF7pV6ADSksK8HPCyIydlG/euWPoKk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6176)
`pragma protect data_block
O7LHkAJ1XwjlHyv6GyL0Yh3g9v7nX2jvwKkUSB3+QWsEtky25bJRxM8FAQIV
ItTHy9qPEViD9hfZAQ6C2aKX3WqPhrO/eNgTMelJG2YNxbITewYy+4EYkb02
ctAdibgiYn932c1C3+OfLBd1N8BqoispMZGjn2l05gpKA3Wuopzg8wbgwIt7
5xmdyGj5rbLc4fqpzVuZzvKNWh3kOcV6Az+4vSzqc+egHZAYaifEUE/pP7SW
DI3+NlkA8pOoc5A3K+HuU9qy9naFeQgb0j7DfDKD1jDsIIN9NF3xUH76DZO7
/5/YJDP7PjqujdjvQO+AZGHpovzCDyFPMJJqrOvEuk5lcW09ZNNb5erEBDSH
IfWbVNaeZQeTCLx+hBa0aQO5WjOY9vC9+8jQxxBIBqh9lf8WgM5ZkWhkT3UQ
YtFqjYT8/W/RYSF+zeXlOI26VCHDydhNkwTPhXdd60hgVG2chcftHFUr9vR4
Ys19pa540s0qK7RSEUHU5c/lSEZRGHXGj29hbQ5IYkXxkWkdq1MRWsYd7FoL
OsoSV9vGCF8YkNJ5T2RYSnY7+2xt0PFsClSnpJNt6/KW6b8tqfzHDtjcIrVX
0FWteckNTO+v8J8y5sAKPyn70+hhi7fhpdKNyM2VYAljiKVo6BuEnKSPnMkR
KjMzoCQkF+H6Z6mjGSHNOP2ANZo03TorXp9wyxdTYdKF77FOs6WvbvDBxkF0
fX9Gu8SV/+4KsyaNuGiy21wyVS3OH4Sbsb1rOl2aIcYeP3oop/kFa6VUgVVB
DPvsp53gTTrQjUaa/WaTLSQe/6nQvvQRm05rgihI2cAhLLcTT33KxBtgaCoO
Qpt60aEchsloV9Txzzdp/+lRAy7X50yIhHKjeV0997yCY1cAYGKUth3W4U6K
psnzapmsKbgOQTIjTQ1Za3sRt/0xLpRBYdNxnlXKrnTHdPwFUQ8f0XphyShh
WgGWckOrULyLWCM0XUAH4jiKCiMA6E/F7T8cbCM0pw4VGuobfte/xICw1/bP
gf2K4v9ZLKYv7rgbJ/pbjKgfyJQLFJAu79iaLxGuLYJ+og0qeqZWwuPqb731
9LbjYsimh97wa2D+SzlPtEtULvW+53vhYN3XVH3rE2+YdGsCdx2WyH3O9v7j
imWRC9nZkfJ3I00hGDUrjphmpo4nrCw26h+RDBh+My6MnTLiXzgdz1lBjKTV
lqtXU+Ca3CWIips489aUrIZlFDcCPWEeTTJOZLMFzlR8O+bfFGFeR0lHEc2a
6PzZKMChKBycrqbXQVEO990vRykqiwS/Bb2dpYPZ6Dm2mFiCp+0ZzqAJNJcv
Pmz7XXOIHAopJy97nh/hQ9sjGLhKsA5jJS/WwNKjypEo60xWSbRuljNPj08J
+OVZlJWzU/ulg/TZPQs5Z5rkOSIjY1ukoY9WkM/Rcen5OSFssCFDszFMSPVm
IZQtNKvTCFD5NZbb47P3kXF/3EnoTc64qkPpIbSmKLb/na973no/HYmyZmcf
ZnCv0YtuiOAYw1Oaw2/Wzd8J2Tjf7zS1AE2WoLehUO9Nk1G2XG/BP6kcX5HJ
Rjwl53Qj86q0osCFrdidnAVobtcsWBsp1Q0JkDqs7ei17uWP6B4pM05gmALA
oDBaMkDreRPXcUbYVFZrcoVGH/N0TdmW9ECX44rbmzqFF841glis9ueuEMeV
TYol34tBwEekmfmBrccogASlW+akhwlc/Qf2+odq4KXHHMoGiXTelnZSu/h8
MMFSo9cPYm6nI53wDGDdUMqDhb2ilF6ea6/8krkVW+z1nIQ9NqMzHT+Eic9g
cJ/1cN+aLK4bWVc7HWiQWL9GmDLmdX/jW04k+WFp1Be6yoXtwCzkSE+xdI37
guVlxEcu79ltlL0uMMZNHCNsGvIyQab5S/mEpieCAEguTIvgyki6RQ3jCtyi
KH3PjLfl78aTgQBAolMFYol1CB29omYYCZZxdzX00scTwRmR7ZZUxTqDuSY6
P2KKXk6TirzaM8HBrM/96HxYobRPWCmFZDnquz14jE3Hu70ti+ubpwp+dnVF
x5YF9Jm6RYKyNhCxo++VkOE+eglMhCNrr3ExB5WstIYIW7DZGrrG2BqmGzih
sIkXaCW/5vt8gxxkk7Cfml1zCLq/kRVn2Dlqh/QruPbLWS7jjFRgXTdTEAMr
UdZ4wYTlaoSKK6YV1R/m8EukvA6U3LGHpKsUwjG3GmnUuu+EjGQJb7ierjkG
DYIx+MfztgZvLBWfosSSsF4jIkrg82XEsXhwb0bv+GzcWAm1JhxI3mkvmwev
2aYx1maVedbuBF+RVDulyGBVbBDeAOONlpdHYr+PZ+dZXkZdC8iwulGaAAxb
5tao479bSX0ZE6dkzlQ7J9FkkLx87bJe/7qgIBpnXZaorkIy+IDJdeCUJoMo
yZpbLgVcx08IlY8+C8Wycz6U2JXbde2g/rt0+/70LK1X5wqHwUOA2TD4A+/h
Wuqy6zXTQ9wCnowszJT2RVj6eMYgLiqbMV0RX1xLxL+V6efUbWptRkeOqxNw
vt55MS5kFzf6LuF+M89ncms9guUvr/MuGSQfqyvXUyKIgv6nUCpoUAnLyndn
09Q5mC726KliFVXleQUhDst6xQLOQdBELDy+yBCF6cOsbYrn0xIlSCaRs2yI
eDGFbUAB6DjdVO/RpBaa0VjABUy7Gu17VUdz6343fPcTeTU2CK15aL+V7oDi
f1gAVLujSzsO32e7tF7kMJ4IMUrw0X6zCerdeqcGEhEm00eIdP6TNpRxD6bq
NTgcb0Dx/itR5f8o1TB6YEq9OVLozwEULxtzGVdNI8l10Jd1lQY7AsDX3AkP
Vp+V2ltHGdGwUg0PdVL+vJNYL7qJEON1E3JWIC48xqxCz8dfc+w83CO1mTIN
hSpboOROVsMrfAs5ZxhM9mQvlImIdCrBlOSONuH9L4J5VbsTOSmjhgODxjFx
4QF7eGybO9LtXKhzOIrOWpc0gL6bLQBxs1NjVEoJbWcBzf+PdFaHF8F55Id1
Av4g3C9C7AOJMDWYq+fdTuUo45uTP7aOISpxAgGPGKSZ9/0GUjdrgj9zARct
5CSK2CHmmb/g9Ht+O1e1vyMoYVfO4ZC8huzTkP9nrhbIdbwnUAtA1gunYuzI
xmiHqyDEjPFKHJ7F56nNBAsauq/bODjZkvCo8PSLnvNUAqcr0PwDjqkRUof2
86dGL96/JMS6BJ/OoS6JAP5OYpy7I96ztc6tdQHkWBrVe+xFCD86KILmwXBn
qmGkOnNsu8ahPmo1bUtT9CJU5K3eI3+OmNU9s/6cJXrPT4diqKkx6ly87tHw
xCF7U/w2c6aD+aIiP36hk1icG2lK3NIzYXt4BtD6wGHodm/xuCWekB05jRMs
n6cw2wk5eXj7pfkGwfG+SZtmBIeiKUCEGzrXIQi7NsgKpe+L/vlFeDF/nbfI
NDWr+m7RxRt3mD8hhm/Mg/gmR1vVTO+JXUQoA0VaXrAqPzFooOPLDPyLNpCt
PIsKpOeF45JlElzF4s+bi4cYynsZNGRwJlFlUlTL2r1BmcZ/Xg5eOBWC+r3o
qDbBR1WR5LqzsO0UvnAlYUrA6JmcVAbSPcKkA3U/TmHKG7OXuRD46c1DhqMT
1L8Cci1lbxRY5u2WpP4NENHHlLxP54nDU8ZaBRhRO7SGHX1du2i9O2qayo2Z
oZDeucZZty7kFMZwOqT5E8pxZ3LwNECohJbG2hIJT1i0bW/6jZPxvrSQgfRL
ANEXABC1wxGnFbnAFIOa97yZVxQSUs+3Jwp/8TTLz3d0ymK0Ozr7McuTP2qj
gwI6fcd+ZG1MJCUqYEwnTY6nfmhHCMWWCR/4s3AXgupnLAs7ywq/3VATdSaS
bf2igfUTdYEa0Q/LReJWS+qmtbPURp86eMGK7CMz6huG9UQ3bSF8fxxYmA4C
neiiw6sLbfHMV1iyDA9r7ycOfExYnbRR/UYm5NxaToIFP7wlPBbSnnt8J6Ni
VB98Sq0SE+QtJQWQgimEJWTTHcSV6wRABOIk+8+uicZd3IX0j7zs2ViN57X+
kA24X03JSfGi4FpbqoglOKzlQerJBgI3G6mZLnV3CyIK0gd0fsMotDs2FaUN
RWCzt2QP20gJ01Updj+YLkjoawah3+zGpOG6sFX9N9W+0t7qoUKX/g/NjIGJ
ET49jHak44uTVXZX1kWZJdlAVrRA+Hi+r1CriQ5WR4Bwl8sCohEAd1v/pCAJ
rRZ0iTG9YPJ7hpd3onBQLu66gOeQitxhZ+sjb2LSR2oe3m9ioOIvPu5bMIId
jG0MRsl/0m+BK5YLjt/7mdzrDW3aezqlu3ZMlXul2PtqFQS09X10utLTMCav
KVm/74oi735Zx2KpFe24gRt1irWsGRHqyEHKhdgDRVPXFznM1E4aWmobNUYk
3QMaSARe9PqCFSWwDbrIqXCw6fw+WxCWIV/No/5Y74XZti2Bqy2lRPkGKmFu
ZCm94Ngxr4A7O68WZPS/D7kozUIcZMsw1DtUXe3GYg/lqDHK1UbmJg6r/Pba
j1URPdg0Df36WaWpZnzs4gPpO/cnbcOPUZsOiTSAnp9cXmanHYT9uqhAK+8r
2/RVT6Z+T45cbn7Nptxr2OiRGq7/bXqdlUGT/cJPas9otI4CPOmGt17/vLQa
FxBaFB4U8a4XpK9W642gxMhs98cT8LQQ7YJJyT142KMmXg9ees9RZjDKA9Ma
SThgOiz2jMDfZqWSAVq16hI/+FsV41lsGCXc/SR6xQf/5TgymdJJKrc+oDO4
mscIxMHzgwWYflrbdMsqaiSuaRYRKQK2KmSu1FOB7ud627L22+t7VNKI/0Y+
G2AeHzDLqhl7up7SuYPCLiQYU3x8DR3vdJiGm9fYa6NJe+kn8olMjRXcNWZa
+kcHyqNjA3Rjm6ztXfK4ONbHjcwYZn+a8YLvcGtH9oT9FOFTeN1eKLqP7AJf
pMOywVORE2udXsfodbfh+XHP+M90xudDssQb4jV3OGq0cwf8t/uE7u5/N2jt
3rcg8zuEIqpTYLi26xlyzrVIlL2+3sMbGIiDPYgFBbOIRWrChw7RiNX3yntB
AXqVnvcEzEzmUg1DrSPUKA6R86uAKeQapxKO983tnM4kBm3E4x+UwfquSOX0
vLMaG7EqUKC4KSBN6QwEZo81ALRQ9XW+tFfPTnh4S0M3JnBR2JIKLcbGT9Ce
s8n6M4WJq61sMCTrpul8rRH/SfDtDbW/YWRvQkKD95k8jmWrVQtBq2AuMxfp
sOKDyWJBrxdk8hYjMTSjz0iionPlAVKAWE6bAGm/+1FKXnBdrnD7fNsV8vam
wmX1doWZdJr1htGHCiwglsksZRC2IdFwBJusjAcVZ6EVluG68XjiGv4a4FfQ
Fty1xkKL4UNg1Tb4Zk4lKmubno/AskpSeDiJC2Hz+S2Lizxm5zQiwlUKD4sJ
8FfT8MRP/BSJ1lWndo/djtpt+zkSR/aMGlJtN0Y778d2BwffMgIi19eSNgKs
MYpegMm67kphn9lcxCdKwQRc55aqu+imn8N75euEN9VpoytngvrSCk6utE+h
utRMv3pUJCHmh0TZDJQoKrSgVQykJk551fKszTmm6SR+3/HLwqvucEYfv+iP
7w7kPlgKBVi6pjikIjDRiCaNRYGdpCkdpkVKmxF23FPGBSx8nV8GLAzLszF0
17/fIGt77oyifa2WBwaY7ignJhopxrv+lxQZV126yHY0IR9ny8zJF2HIxb10
KWUfUt7RGvFvgi/fAtLTmJKRMQih8JKRQk9IvLiifD9IDeBtQUXskyiHheu4
9e2GO8R/zbF/IlxuNDwJNmPX41NzOiZqADa7MNVF42cUTTqxo8nwBwaizM3a
H3By69jAuEPBgJeGLlWA/zwDEhBLLUCfk5c0uoCTJYjuDGotOefNOx/CBkgN
1UfnKlKFyvWRgCgjDZXAUoYH2cxd8PFR+YB7xs1z8lLg5Xk2FG/HO4j1AQ9p
BtTkwfJ35oVSEQIJJx1Hvlvpp1vrJt2uGv8jvBAGiFbBqF9lJtSLZKKmqauc
tUwbR98PfHrN/MtW8oVRK3jqaY/baFqXGWIFwF3y/QqhutmoWSTEyjXnVmBZ
hVmyK/DTm4NiysUdsviZA2tGehN0qzxgciOzt9Mvl1VK2m9ufIMcKYnmIRpD
eeRKOz6dPrQVD/UNAP1CIKqAuplaoqtbeNaawirXrERn4PNrF1vVTeSW+bnt
ZQI1a58wpIE3n9FWlUgkwfvOCYy0KA9pqb905LSYmuDGQSUdDwy9NV5uM92d
EUBOumOKO+TkhpDxjD7LAOHcqLHlq3kaLDZl2zJfsdloW01eXTPUN4Q/DSHi
QeIgF3pJ2L2CIG3lxSP6b3COuYmb4Hh2621b0KBqsxSAE4sKM9NRjQltJYZZ
FXynb715YJiaTkKcVI9eVU3hqO0EwkahP4RBJyJItAC/MFjvU4x1D7HbflQ2
RBX9jeYsrEM6D8uM+rTHK4eT+MxwKlBNPMAHyU0E+XmXvBFIeGif9ayz+Q1F
h17S96lVlZnkjVSd/XmMWWhh4i6rW9JDqxeedHLL8nKKToUSf6rUBmf/j5Kz
XuNIEtpHgSiAwbWRFQEj2nyrxyvC5SjuwwTj3BkNnLZjjOUoowR1qb776H4x
Pc0lGwHo+W2vJHhtPIGaOII72ttgnccqv/YohuWDO75wkNNIsnJQYWADKSB/
MgAxRl7AX6SynGNHNoLxRDnS3yd42scFJAcwyIj8eVCmrBEXsSWK9jq4egqd
Nx4/dkKxBae7iqEot21fEaUCTJySB4szuHjJYrPb//icwOc8TDnIRZCk9eMo
cigwEzG8d2urppE+wQUy47tfEfOUGeK43i+GuV5jGndL2m9Tf+ktG/Jy6/NN
ZDB0DNoF761kdr9aXrEfCQZAUMmeoF542z0LT99NKspl403iZ5S2ycN5b73E
adXTGiZkdhXf/T8s7cucZH6ON2djDf6TxKIQoexpe5pmPOGLfP4xCjcagErF
5X4ljRJiSHFV0OqWJc+b9c1cdhmwmo6UdhoiRfCqrazXtTFrhvs6P8ybO3o7
dlSf2MzFdKIAULIavvyhRSPYUm8IOkLe5aqvjDjypVnIoZVDcyaINxzpGJbl
+4PJcJmcON6qKtfhnOtJf6pr4UfbeyTEn9qEuZCUsJnPk1h5b3mTYYDOJzMy
WywLt0LJ82CrKqHlezT6pqbcLKSL6fDgnHGOQSHNfx4UZfcM64al+uQJF15G
+iO8DTPc4B/gs09rgijcUJE2XPHxU8N371HZMr+BHhwIg7wLf6yESOsk66ss
8BsiKyNXg07J+buH7mNKMYi01UdPBDIlstFGHPSC0EetVw56ayOaqcAMG57t
LbKbG940oxSYeqYqAcoDVUuLoRqT8Puaz4SifDTzSkf6vNy6CTn5t/p44D71
2y+PO1n3CpJCkJCAQRZd0N+AnXXHDeyf3U+drj3ouy8b5jisEnVZ+LzQwyQA
rDg9IXkCBHN5UoSoYuo8YVfQNWasIkx7LcURlK77Qg6V0qzpXyH4l24SCENn
Wg/PWY7P/1Q6srDJMu/llYyG99fm741AbNY6V/2ltCyY80eaTGIzC7RSTJZz
jyZjjLy4+KFGY81n6DVz7TUMH26OU5hM/ahuaT37uhV/M+Cp3DcbPgb0wXk5
m5cdHRRD9wj3IkpOh5q+OB9Pb9wexIUuYqbISWve/M84qTmJ1ZEVwuGbfWDf
QhEM8HmeGOEcWok3Ym2NC2gCPzBZskY7fsmoX/fIlrlAv0lmR3o0Wkvb+Df8
Vna9VVVmAs+972AbHZNwY4R5KHjKNAhxQEC40KKkGESHVJEQXA6iLxskDkuu
z5WETynYYzONLlGpG7Byu8l9HjWGMebTUToTC9BlorQr1WoeldB2l8CJfr1G
J1ed6Iybi+WAW/dGGcTGVTDhb3iTVcH/i5zd8IAHe9Uq3KDbUw4+kx5IcfrR
W7UhZjo8EjDcP7lnFCrFXUMqtbgmWrmr7bsvSBPsy876jH5iSlLeP6aOMDT7
nlhWC9H3TYoX5RwDFHyhy6T5N3EiO/3Pw7kMx1Jg5yHkDXfwACE4XCjA8R7D
iFgn7WzVnSltw0yPh4gwWjwBGLY598DsBBfY0zlPX+rhBluwayOR9AODCVBo
AM1p9JWdcNa6vWZVcAOVEnbRkJdU2bfZ2AIWvGoklrKcl9E8f5GYnc4GyfGn
brcA7ZE3yri5CRCDgq7318SZcYdgySgHuo4r/HHV5/vuO5uTdnX3hGUmjrx1
gdbVjXBXUmPeNnc=

`pragma protect end_protected
