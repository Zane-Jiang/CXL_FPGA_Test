// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Yxs8iesxSTaPGz3qm7IBWEjIbm19ugzGMVba2MfVW3jEj5+ch6M7jTbQ0i2JlmPy
uMjjetuHXf22LnHVKnRLwCp7Tq6PRQ+w0HYHhAQMW36bVMUG7nqsgqvrxa97xh3G
1bGnro6nArM2AVGKwWLfkN7OTz6Zb6f2g8TNMfngaXs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1376 )
`pragma protect data_block
/rf4WRLMSPkVt3TPdHBL4TsP9uH84V41Xs/dWhF8NiF1MGh4PXXKLQtp1eEJCij/
Yk1Iz0ZrM/V231qQydVsM/ElnWzRoAFkPTLQf+5xnKjpXPFqENKDuhu1qPsyR/k2
FUeCeYAkcY9UcIVxx9mBJZIAgKhyzcczveM/UyBBZ0aJb6EEKk68KmkQgtwHON3X
lexqJenBy+3nF+5HcILZNvOc5oRjPkkC57Puen41jXtO6rxtX11i/aT5Tg5hpJJc
Ux6AW6Pfup1zaW4VoAOLQhBX50Z5Ek3ce3/XGGaIDaCfpIEv25UV6s7PzavdBHCo
6uAu+fiaekgdqVvX9HktPSUZmDarVTnMCk7LGuZ38Yopp3amKnOfMa6Ue+/l6tmq
fV4GTcVaDbzeTvB4qRF/HG6gJ/djeBXyvfXejNstEB34QLLRJQd0EFMHnBswd+kD
pY4fmhlB8AiPYf1wNbOgQyfxGRsibVlUHqT3JxlT4yeswwdK372DNc7yPre6cB2C
MBv2SHZJm5lzBW9XmR3g6LOu3nTP5hForD/L3w/YsLeOc/1EfUA2bYETtz1+Y9Vu
DSiHoixBsxAcMyxRQERfjvOhav7X00SNdp/FeGkzqCGxyKczMztK3ZJbMMsmRWux
arZrCiK6pdCg8MzK02Z33ZSVpxc4vbKqEK3FKMYsFJJQAQPTYkGlXYj+9yzLu8nH
/YcXysaZ4MiIqQQV/b8Knt5dDY1fmO2AAeQyYuXVTlBJ9asvcLncW3CTEZU+2R1Y
VvrAB2EZ1psb05XFnw0lOd8xm0HBTg0A7GHesJNuLl/ojV2JlXZUhRZRefunIl9l
2QBAWZnua255aMtpp+WNMHl3sCF4duTtW5YCTT8aGlIG1hNVfH1UbIb7n/0rr9/m
uoSyTI13Rht0LZGT3oj42O6noRqHsEs5xWmBGLL+qpSRPdETTuhIQJoahMqlWPea
1aO672n7xjxxoVPWlN8paAbmUWOai6S3EDPp6gQYW0uJQXPqdc9oEP8rn2DfP823
sI3KNI7vAxt0XgJ148PQldfGOOLVQ4zS5ismJDOsgc3LORDUbipM7hnoOqRqdoPS
MgIy1KRSwQzlbYF8Wy2GQcmTR/AzQSU4LAfoWnnnbYMt50lCRqEiJZ4era9iZNSF
yeNJV4x5ubBP1EkYuWie87TShesreo5gHE+7PJe/iIRLsJnN2HJjZYtEW/SAEiqH
+ZMew24NAEjiJg8wVKs3CYT/LuZAZAyHNA4OLq/tKZp2YDFCZQiPRCaIgP+Rwu9/
Ig5vjiZo0CU94PkXZKBSDJkP6lbNdWVc6vwLgZAM1oVZFnKp3UyVd4RrzB+FTQRm
M74b9RTolQuJlepr3HUGdbMSR1g9VWcUcb6KJb0PYUrm8vCEh5wGsQ06GnVBWOq3
lq4VqKcz5qtr1pD8JD2wilyvObX1qffmUm3rjoF0wUzSnBW3xaZlD3eKSQJTwTT7
fLj0wnjjWrvCzAB6FsRqwpnXbN6PRr5rVLDNWCRYNVzypdI7lMs8A+av6LxHwGH3
71LQMtQ49ANsWv3T9qXSwn6CVvcOH5goSt30HKEGBfVASw9n2PlU5EVdenUkTnvN
3wI5i/zEr4Q/HdYxmJn24qK1VHxLOEm6uuJRtz7s9+ypueDPPTvKSDwa/2hp8I9c
PyMHqEUwCAxdyOhVHlkFww7ykMWS+rgB95U3vXsa+vMo2e6blPNwbT8AIVujRFY+
cXyyGYXCX6pjI9dMgpbgn8exRuYBSAcUg8TQ21iRXlRecnSv6k9BKDCHE9krtKoW
jd5YsfygKKhWEkpZ8LeUXVZjAx1dvpPX1JAlwG4T1Q0=

`pragma protect end_protected
