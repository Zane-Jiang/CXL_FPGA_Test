// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cMmyt+AkDOfIS5H6my7n6ZOmGYar+FgfJ7z4VqESzn78oorlOruaeXmxqWem
/yD7zucuxr/Txy6bvC0SJibo2gynMICeumll5BWlXUj10Mue6Q2S55GQNZTp
uUUuNhIb1H2TFvXiHlWmDWYvqVOSN7XoUkU3GMZ1ESEY/Z1MCAxoWqzN82Dx
MkDqrm5mXDuIzYHHV2AKQ0m7k+UaGoFVNR8SccuCgNdJXkEFQx18kKQjxCOp
UQ5q/wC+HHBSbvUWOYXawxVo0sUKKv80oFJq/92wHLqObM3n89pD1hefRwW1
ltSFIK5XtiGC3ESc3yvJitkJ6z4wZrKQOPqYe+NOAw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fOOzdjQR9s+NxS+GU6YZQLx6YBlJ2pjkj0XymxtIlqOy4Zizk/ZVoPPNm9Ca
lSW7rNwfL3d0TzapIDBGjRqX7mCM2DD4ciyWeTvarr7w/zrS1DVryKZpZ3ml
dFrgT2mKH96Mgv9eLII3kA9Nzyr4wYUL6ePoo3WObR7+Rhyr6OnRKdU/baOk
h1lIpQMci4cufMivof+5RR6lPmrVUJBIszrFOsoMkO08UwpmSGJt+WBugU56
wr3q0M0D5ZTep+fe1O9P9tSTHAVNNBbbN888f3P4GzC+l86ulww50LU7gruI
5j6/cvE7wm/ccZdJ1Zm5vUX+/OlvE0ZXxVxRNROKAw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gU7NiyPhqpqoomf8UHSz85FE5OQo0j7EAGHPrIWsVGSc0ygfDdulg6yiD1Is
4aI3MIqbwGntMlErCMCC3RbgPqx+/vdq4Wibqk66UhdLebOcZA9Szm1cItjE
qhWaIZ+hGNnHUmUCwQnOlY1Nmx1Wz3YhZxNsIXYEodzPz5zM6BGCFuGlrmxF
spMaHBR53CHYl9oQAnERDEDXe4AYgkwyS95+brtEXlqBpFhK/V0jofylSxko
1ea2kXg3z+fFhxmq+9U3Yfulm82RtlOzh6YgPJf/U8jHEMG4eJetaklXdbJs
wqbWP7LiauUrpfv8p8JqDJDJoQgNH4Z26Ni3N8fyEA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AVFvt6gLjgkPkqEOk8dDv9nP6bdCP0KcvgeVve/1e9Kq3CIMsAJR5LG8lLXo
qH/5PfOpNITUgxefxje4dUPdrnYl0/pyaURzBiPbbcT21t+tGQIb2DCm0Tq+
HFZjlFA6MY9PIA90fTGIh7/utgmVoVk2EHSMhZPBV1Ir8XNOAOI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ezMHE3fraeI33kEM/NA9MFLebLKjPFh2s5Yz087e4z2nQ07QRF3F/UyW90W7
K7HNTW1G3tqcbnXoPkLxqXT2cCIrv6hKDXkzXA8sJfznzpPdru/kcGWdS8tb
tNFkeV+kMtTs5mK9821HlPQ2QshN0kIGuyGe+N6qT7V9SsMFwDjLj1YVRYyq
ikguyaRXx4UIKNNuGSP7ORRjJlXCkWU+twYp6fs+Yt2Y1Kjps0CXt50afsaN
SNGf3QwHyP9qPE9JhKYD7WpbhqPVDEBPJtsZ6oLp3Lrn6jawROo1ND8JRSV/
b3uSKMNsXyRmlA28R+sUsrzH9TUqqbUt50RXgBVoS/k90gPFclrpQkRPOiu8
kl/SQLO3BfZOC+8EXKogmPzP2/rJECJ+VYMBA8H+whP2mrYYSfIE+mB0LphZ
zv2F30SkN+4l5aca8qe5qIy8Gw7OZcNC2fiE+ezwju/CrNHy8dsprbBTgAZ4
gtpywke/6z1xcWdBzOAZhnqpUmFC+xR1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fdLH1mT68KjGttpMLDY7tLLJoWqYkGfQiCz/WFLrEx0RFpyrRQvQlHlZRcJQ
UxrZLGzIeNpd1YWfkVYRD+1+WfDtxQNe9HU7l4Co8cQi7TYmc3FiHv71N8sT
2DfDpQeTodFWMfqGQX2/ISmIhncq6Ps810DQg0Dwg4J2IQYCrWk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qx4ayLFY+4jxe4jLMt2/+cLLbAl1owPLspv4KFvHyFOcfexok+J3+veFvQIb
+oKXhokVgv384FdlfqJR0va7AaedhHaxcDg3ZSx5/gQOOLBZovZ1wInFq8B0
2MYm9U63e9zi7BAkG/rDMjkWCJWxjeibIdDAmwd3doO6r/NgSKc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6688)
`pragma protect data_block
ndAPAMMZwFPkUiP7vTThKxphXF4sYoeFfLY7Izfl1xagoDaiFjkAjsnsrxO5
zYbpsJItPwDKCXOYnm/QB/R9SKOpbDHNXTJ2pAMH2wNG/mW70iDrP+GDpUBu
0N5e7wDSkXp0pcHNy2dMWlgLcGa1W3NfAbndaK4YJumsNRWXTUjLztV0SQuO
i/zikyVsqTx3u0i8sjfeOioW9DZD/oZfkopHu3yroNV6PPJJrpLDzPZs2jnJ
YRgcznG+Hlh/1N7UwIwXnPwHg4BjGSQmJt7rp89FVmEvlRuR6EPz9M//aakw
mCme9Ex7iOg6sHwOfSxK0XnGw3Q/y4yZ80BxP2UpVdSAKx8soZiwW26WN/Um
Zuz+JYbNrWQTcC1zWQiWEILICj97SMihJcySYYMcupnkPTHU6AP3m2hF0qwd
yd5I2EKkBPqVjzSR+0WVZ/8Nwg0Gk7GBSCkLPLZnaj7IDq22kiicylO4ZeQ8
ANuJ1pWMo324vpYRvwmvWqC1Fgme9YA1vQu3qAhIp1g6AldRmHANTtu3P1Mb
Dkv+IatK8yU3nqRfAVHFdOEArcHJE16fhz+GuNEyNaV76sNMzTa5I3U7oEef
d3y6EnPQgasovdmT/FEoQ0k/GlDcVo8DtcnlqcoqQp6cYI0XgAlh195YneyH
6ibXX6+Wet3etXxm+MNa8baycPOOAB9WLQc6976EuwjF1hbZWktix6FY7u63
i0uPCdNlIypmZXZSFaoQAWdbfDdADBbbtsS7pjhVCHG/YZyreN0loqah1Q40
Zgil7c41Gf7xdmmwe2uB74oV79vyK9/xe7rOtxKL+u3znVQpkAOTIYVF20pl
9e2czR9A8u8mA3QEZgf6bXf8RTLRtmeHfomLgXSN8BcA0JShXFKE6tG8W97o
cRCvgGEfWf8IqmdIwqBFYucWDqrIrvGWBs+Cc6CrlHKeC/NG/i+OorGfbk8D
kjDkl++VC9wE7eFuL9lGkZzoFz4x5BcOkllbnKKs/Ez4LZ31VUtNlas4j22/
uLl72FqYWpSvjP7I0M7XbNjeB2AV31b05803GrEqWC+Lhzg3uh82lp7DuiwK
A830yyNa206L/yrS/1SI+S46u2jpoMQ0++OZGMLpCdEDesnAHmagKCz0/aWu
aDgPH/hqAU6HABbj5FpEhG0pR3/GEFiKalIH4ivIKAvusQCjru30B765Hef/
ilPRh6oipuzYjAj78ioWiP9bDdNzdc/GYGa+fS86NUFkU4dOLtdAMBZwDP1I
NOGF6xk7TkcJ4gBPpfP3cU2iYNCeV2hCog1rVTS3l5IRQOV6tKcl1VqpWPmX
Mdr5fFlB4jWot9RffFGgqSHiZNjZkuaNP2nF3/BkYpoisnjA0bAPyWxt6Nar
/L7UDcAV46v9N4phOm6JQmiKyfGv/lpeAe+7JG1OGQIq4BJYPmdOeomP7Wn0
4RUwgLi0rDirxPk1lG4HV44WJdDcHb7UCjNmOvceLtB+rmtzesxxvBme4ohs
E2ysfgd3pzkRhjfsB9JQef7InEglISt/aGARfNc5u4qdgJAccgtaCI5bk+6f
MrBudAct4pQ3+m8GFhjF+R6Z99Pe5ZdzFFzXHD1RnQoSXiCPbmDDVQIyb5vX
6wQC0wx7XaGWqrHgDVLHhHtm21eA8cTgmmaLapzsqu8rUrEmLlzGChaLdqoO
WBW5SQOzLOVrRgBIUl5/H5C3rfEZ1n3/TCqUOcUGmz+MP9UVj1qjZut1RQvv
1rkEVLFI3cpZFmpzci9Ja8Qe43X+3UN6UUyWp038GChO5tMQ7oUz0qHG92r1
nLq6RrzX7prg66Yt8fgFudI32vuLIgvj300I3HqTe6ol8aoPxUgTCb+lua4F
8OJAsrq2F5Pce0h/V4MxjcZLCBvIy8FvA6rghuKJemFqFiRPfmbCLJpLMUo2
FhPEKxRBESvu4jtW/vfuolIciJnuC4fxMGb6/Ff18K3ryW9VFaCXV5/kiN+s
yhRANx+1Syer6dokxgkoo1lPM/R6ASQmgfzmi88HuryXfhoeC1Iw9z/V5bUV
7Q1PZoy+bvcn6uQylGiJFnMfmNFFCm9OQhwgMcYTaBkgv3ZfIQhoa58BSNEF
a2R8amzdRCeJofMW2qkANudbp/poGRe3xrIfpQB0cbXA2S480KClHhPLOYAP
DqgybCPSAj+KT2EjocuxNePxwO+EaFxlyqIv9MmV78bv19dNCUv3MuE0xtYx
Jw4jCHpwXpjnU7o+2OpQovjixayte/IP1jCUKbKYV6I3uETXkG/TINE7fUV1
RMng30Nr3QdZebBh22H+yPxpl1AiWzF3FcBE+58jQFAB24ct8idH9nzCavwd
k0Dv/iQSawJkHrm3+7nkngzvnhO3Mqsm4Cx+xBFovu0666oClvhS7ercMt7U
BrJqWkRQ7mqvL2etIylNOt1fUayRB4NOqg94lEBEAXOTjeBJscvSPSxSH5uz
+TlkVjhKCdsbp5GjilB2pTuztNdaFbSZhbVsPMhOnLdhY2MBxyn6vxK9e1JX
CW2Q4X7yxb85oQsSXt7gtF+0koFbcm3H3CnuIQ/YIgHLOCIynA8HbNbAwowj
uvHthE5NsIqseVnTVMJvLlZHztwmFxvmVycu4kqxu35+htZouMybj6UZE2jp
SW2ys17SXMMCWAmELd2V5Kv6qehGQ7b0xsk0tCBBmEsdecVzPYUOB5GsyXQi
pcOgrrZ+3c7tjNvAkcLvLb/ytqCvgs9hk0037/yLQPUV70s7/jrCuBTrVj+v
BELZv9ufR8Wx1iQVN5kjviUE/djCVZ6E+OXqonQm7pGJI2Q0s2mZsR0rWWz9
XjGJGSZVwMaYW6MS/c7SAZhUd4VyNWkRKhfJOkDUagi6K6rWczl0/bOODg0l
eljlMABF3YCu6609qHS/4t3lChNtvzBmQrf8xME9TZ+Ms2VQniWkENVRhKaZ
U3HPPsnCG2CYOxLxOsx/lHh7hnxF5WuIK1b9Ov4Z5EDYkD2woxQw40Da4Qfg
Lw98iPGe6PTHtaO86aZTK6EQg0L3FINSDa/Nle9MRwIAjLZdxZRm+B5Q5KEU
3YYCSiKMJVniy1ejrBuz5hGITV+BcfEehKy8VYRYyCX9VASk0faz9VQee18n
GDgl66vO4aqrxVVio6DcCqtydP9TLouTNOri0SUh4tQRm4vahv+56KOQBYb1
DEsgKm3cOzVSOYazv07jWoqo+kGvAJ8Xcw5qPwrrCxKWatUZ/r+9eircdc5F
IJPharLrw+LJCU9WkS+fxjg7j/bEtRkH4nzVaPchlK3SVrnrDqWRY08HogW5
SLRtLAcR6r+182ilcpBEbgzjxaLep5TXSWdxtRQKE0wvNMVhGhdQyZ91FA8J
sl702/CR8nesPJkyBIzhVzaILb4Wbf0bIY9buGeJThcsmEQUBiuBFaBbmrEX
ONe1N3lVzWlcVFZyrJi4FXU0sQ/HixydmF1YKahmp09I/1nWxkYR0+9/g6/R
GjlZNn6G8bV69egLTcFrrdOPNUvbtdNO8lM1638NKW9KPe0lcrEhoDk8gA2f
8I68mV6fa4RgWPnaCnyQ9DYtuXbyILjUD2yvA/prmRv3GqRgX3WYs+GoG1j5
wi6m0khmma84j6T6kN330qJjMSl+xDM7KBtT0IoCy9+3rhoCODdLbDvv2m74
QAJY2+pUb6hYjPVpSHy9HTwId6zH0MeoZc3V9t520vzdRjJX06t/rusMqadW
Vf6+IRdDdaZrmXHdegyeAC4kaLcncQBqRoA7VoVyw7L57iiayKR0AnYE72j+
MNWokZrreRaVuZvMxgP4zqcywiaG1h3DSos4noZNA80K9HM5kHF90QwjPxzJ
fAmHK6JYD8J14HsYWZORpKQLGQwqTtM5Wz9jenNzfIe721JAB73/DORw6VsT
tHMzcnjZASbaR4NfiHLPGtsjxiREcj3JNFmJ/U7L33AG1EItllssXC+7yxWC
l/pyTbSXVGWUSuhDFveJI76l7Sbbe8gT92GOEAQG3Ft1ArPqKj6B/hauY9aY
BvzYMx2vzvJVu5CI90XUOti5T+41sEc/pCL7Zp1uSVpAcnECAwp5yMnSRYgq
QL+qmswaidh6ZzuO4HQcbpF/XWt8+Vtn316g2aAWiEmY5wPPR20cAqZrPqqB
oCiyYAhi+3Uo0GubfH8BJCptvUYtGpIE+FUHJyBsTavCzmm9cE/zoxMGEbqL
Yj/zuKYMXhij5J0yZAN8S7rKa9FDvh7Rha/5H+xqPhvfp+OHsqKHIg0gJ+0y
nxIey79dvbTUxb4eKc7adXdTUxwkXvxFyBtkxZZvzB/SN74glFGTMjN6xE9n
KAADYRerg58ObYprWORU8RNjN0UlJX6Uj6qgVYuVK3wy1Xfs1d7I3ULdP/s/
kK9XzLYBGVmbOJvvmgDnGsko5j9Ef7wY2kpgTpsFDua861yt+2yLXA5gxCgU
JxpH5ckPEZwbhpbBMuFqMvM9Sk5nK88v2KfIsaPDjKWSs9gqHg5T061xs5J9
DM3GFOzWRN4qV1+Se7mcT52mQGDa5YqV8sterv07zTd7Cl8NIXM0YO7Iu7pv
S+1D++yUk3E0yUx6ceFMHidzB7N9iQuoJNJShvn35DQp0uYMHkCNw++tqAOq
lawzV5tKPAYH5cc/bucBq3U4cgOVpYvqRgOrW8VeaQzWThU8/k23GpmCNPwX
N0tGaJOX1jZ5MIRtWTe9YxsbiLXlZnqp9M2sUeZvPG66zK4r3taCL+s07oCn
MfRr9FwQwu00l+TD60oyVZ1/G04F1DSOCcYYTKdI1gu6USYXEFX62SJyNLNd
y2+c25li9qZ5LSkrshf1Asbk0vCqxW09SJ8APb9/xSkc+dV5YcEghP6L9htb
viVE0pdOqIoEpSw4MXyzX2ZjKKZbw9AQdX1VTruFlP5XJTYHADRLin0pxb5X
nxMNhfAId143lkjCyaZUqa2+ZPPEHPZSBK0TI4tNOlJkOi2c5SY5Meum2y2b
jgCUVQlWyWmOYEbIP9YVtmHhxHn2oFToVmLvlXYjfYwzmclFjQLiSKege+aR
05h6Pp+b6edCKBko85lwLz9NSK9b+zXIYTOBufkaGj6od0au1Mt41h8rOPnw
6x6ErIZECbkB/NDcjzOCG9iIWgb+wdbqbfJfT9TR/+MJOobtL558acV5MvMy
huEi2Vr2HkAxDm5/WSlui5BdKl+u08cmL8u3BDe7S0jpnDkoe9isGrNjhE5r
ak1N1/l+k0qvvTBvBFbYSeGMDqSZrbmWTNNpM2/jUBLiXt15LRyg6ehj/GrH
Hl/v69uXli8blOywAKpWiGHnoXLe03HQt2GqrIJXuSBTKg/byfVQfgRCsTOZ
ykIuWYy/VCXhFpwF0D7lABmw/jTWGqCcTYHbDZn2kBP2jImejZG/WZ+QalS2
F/+vbR6Ks4WQuEJc3seukD0cCucqwTOZ6q5hhyjTiOZTEJps8S/6p8XZMFRZ
hSaX8K+vqgRzLfasQSGLnBNOreYRiNyMWE2lKzUPTf6CvALvE1WCXLwWpfk7
bszhqZl+i+PO9oD0iC4s2OWycjuI4UumRhbfcz76crmxJV27bJZ8o+MIX5RO
2ejRZNyj760i6CzZn6i9bvE0GTxtV9XrKOURMCRVEEvkh3d4fS1DQme0xDZj
618+P3sgoc3B9lTcw5lHUN2q0ZqBpqSu5lzuxkd8svSGuWqxCT9qlLZLVV27
CaSxa+j1KgWA1lElVgcZimcYJGZLwPsMO54MCvSCE3vBuAHfnTV50+VqKBdG
BGj82Y44oKOgs7OrVbbkVENvMippVmjhJyjJgfHYGPzVRzxTHq23YFY2M9/b
2Oq5Uil0jSR04GpBnAKjsYKHYXiWa1M+B9bTWmJYahPUqpj0l0jp9A591ueN
QnF/ZNQvTDiGw6PuJe9pdEAZkgO8r5nwYon1TCOtg8zroBZjQ+S9/XkHMKP2
GdlwiehWoPph0BPNBzyESMtnO+c3ecg6SIKG1QeOK0UrjB5iSfnVc/TYAF0V
+gojt8cNbbBWlCbboAC1HftKag/bRLIxHZBsK+2h62MJqYEqaNTK5jCuIkTt
Y+n0kw+xxwn7NWzl8l1rRuaMrQGku8p7dKYclfKKu1PQZ8WO4qOHG19wRYv6
7Du01U1i6pVMs+ne0gp3MfVChfC6ZOIdgROyfujmqikZ2Gv38WOWhPINmyFJ
rGonN7vq1LzPN2UxreWzzyLB7w/1jMbc+EV8A7tXEGcS3lysjpj9h5Bd/AK/
cOQdjwKye7WLaV9zBvHln00sK4bvziajmPoAPWjmh9DjCYcUhzR6WTv9GN+o
jr9kSBftNx/HidYBobqS1LrEZaN8q4XVoABDvTuv3HaPXraJLe4LU3CT1OPg
9Tzi182IXQ+STci0sDlloX+diEcO6hU2Dht7kxqGL4973Lo1jdErx/IrOhBx
m1Jopdu+zeIs6HEt7h8+aBNj6rD8+9keTNh0Shs/vVyMxqhH0UBJ3BvcfVX3
QCBJgZE37rEwnaA6RXtq9nY2q6jzIlhIOiFQugBTwIyiPcZwrML5tJThE2se
ZpLGsdSqK6O463xXrcbxq4rJfsklILHsr5CpzkT2t+tiBLs2NbZHf06wikfQ
QQkOBPeZzkTxPr44T66NhazKxj6/gKKzePl43mbR/LZngRmxAoG4sfD3fqy0
hCAS9MAsRCdQxIANp6BcvP6VBv04LE9/CgZR7l6f3rPydB938e1sQVMLrkxc
ryjYCi/ozimJdNxjynkyKeR3/MfbHyPfI6RP8joQARgmZqk7sGdoE3cHj83E
BBrUJFb8KDwnSlefmpojxSrlGxG+/0BfHJpybPBfvgmtm9WZYCF1guoc3h5K
WoqTp+16D4vSTecZYCRPEK/EQbK5lMP7qHlvOLMNYTv+u9lVmoHccashkezc
Oeaq5Ms0+zMy8pqalTh+7I4pxHd7VXkb+slX6V7aosO6VzgZbjy9vs1QDyWw
RD6v5hhASg9rc7a2OLvYHPDYWNEHfkgyTz5qHZiyInwidJCwpgEoYxZZ5qh6
KUJuerDJ5O24CdsSsA4ReXAPek/NzzaXpgRahYcDhPVypNcqzhYdncAb9EKe
WZJ0OAKwusYsHXDxAHF7jR+WM0TO2XMtABZwk1OCe3wvcKcG5t/lKnNfuBYZ
Z31f2/3kwf6p11HNqcpBGaqkWG17TG7AL/QrJMPZqeLTFuulih1QfyvO4b9N
va32jtDNX+MeXd0Q0RUTrK6XRQw5LOUVxCNXSiD9t0M/GliilXtc+eiltlFQ
i7JWohMq/Nqa3xUEK7mjzfUVnm15iwlpUhzmcegsT33nDssOCjl365RUFApN
idsfqBVhwy5wWL3DTMgrSWb3VZL1NN97TUWVdJ0Kv+uU9Rp82u8RGm6sed93
gdR/Czd/oOFhhGIRyntYHQEEnYrfUyXfK2OgKvQng/So+z1qxzjM/L29rqAk
kmNTIDJF6bR0urkTz2T5J19szxfx3lSavFzl+ZORlTcUF0BUurOpVmXrzFI5
vk/ThDzrJYeansUrc3eesGYqNFTdqR//5Y82Y8pWQX4drZOPsJIcN69JGRol
xMoxB9PStjCm/yjAWaT7IBCl6G/t9lxTRvPt88ePxEZKi9avE7TKZwQY6A3g
vzuM30aIcH9YaXSu5hpFMcI7x/S0QhiA+etNEw8OA9GxFiiNH9QhERJy7Daf
/miOT4pod4AAtiu0dIn8s3hfaROWY0XOBCV/y1A1WkvJCNn02HPtKf6+WiDn
Uav1LmIrkokLw/h9Ly+qKjf9A4V4gfS0+AkeMJaDr5fOEkdsgSmAvxTg76hj
/FArPJda1PUqWKHpG0KGUAOwUi3hm+dU14/HDYuwR8fuIAoyTWlEsHP9tEPF
P8a+nEOPyihs+ghVSf1RvViB4t8Zh+/c0LICqAsGkuN5bPYBXliZzsgVQ/EF
B9L4SScPxH6Vmrz2ETBJK5drK7xHDzrn0qTyM6mPij+ppICEQvz5j6zcXmPS
v0SjxktRAx9TxskGVe7t1LaqCmiOIvwpgcvOHM0z10f+kHgEMG7XsRapQlTA
r5/czQzvmvsh/OHqAH7Ar3lhyQRgTUanUC7v9v1c5WvsH6TcAAr7/0+xqkOO
Ck924rnhpJLFt650M3pBBM3AD1TTPsOLJ85zNfOB67UVKsQB2aNyPzr3tVsL
HsVotIlLio79pmLvYZ8AeFUcKb6VUP/8a815PXE+/hgg0cxXsrWxj9S8z4Dc
Em2gq3nKm8n2J3eQgsr1itkNdXOFHs5Ekqq/4PLzhw5RDWagToQ1a7871aZi
0aUKEK4moYUPClzhbtjMC2C4i2N3q++J+I8bYSqmKGG99ajLvJrztYlOhIWL
jRHtJ3zYmMvElcgnPULYE5VjONrZZTPwHN8qmj/LQXI4hCK2ap67rub6T7I6
rX2yT2ciSOETNIuUrqGoGe5QoWqEAjetrb1gIXazf9NtcpDpt6wy9ri3o/bK
zqvsujR/YayUu2yAXhY4axBaK1NZYQBbF7YMAdMzpnhrDKi/fntci415SKOZ
V3uGRYpeLZ4CbkF4VKvxGNqzy6YjbwLEs7Tdp6BSzr/p4MP5z19D5JJDf6H/
amjWLSLnR3UPanXjzNIlsWOEKUYdHgTUnNRwzxovSmEG/MiUWnEwmh/NVW3h
+2gcAOi8BTUkmnPlXrB5LXGa3lPmQfTRRR/qBu6p7M/EiKhyx+MY72zTjJu6
C0YYt19Xupeobj/C4YHa+V8+MBqDyRQU3oZV3Q8eD5mwBziqdI0mhsvEzs5R
WTwDswp/4AGT6yrklxgLFT6s6aqB2Nk/L0qiu6r6OB5KJhrtSJUo75246Lkp
AvDMFHTHxy3hjnFCszhiwyJETAx4WwxXS5yJGCmGDF+UwJYwi4MTdcx2OaQY
ERZthkjLDNyRXIduSyUbs0Iiv5PurkVc2MzjBA==

`pragma protect end_protected
