// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ao/KQ6+Q7NxfSuChp/uhI6L79p5gbBa6r6fVQhmMx18b14d7DAIcUqX0Ns2o
PBchYXzwACAmT3krcALK5kV3ucVfgFhy42rGFzYIRab7hM+NvAmWSWOYlD05
0S4oMVlL0Yn2NhOVHbGruIFFbHsEJDCzarO0DuAh8fSzN6xNPB14dHFzqOm/
7dOdYzKrHCCagk9ESzdYU7kKVT1E73JIOC+ygQ38lr1qP4rcdRy2OEaXHcMp
zZfSEN8TRv10fo6ksaAxP48SjTRKE3NE+gE/kCc5yqjszLO4p5aVJD7fKE0+
ZTcgpcbMtfGQHzsmV8LH7muZ/rgDNqbULjsRPRroKA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AbHlCcTlHkKxQqUe2ZI/JLyul7IDn2bwnQ0JEGzcOsDgeIZ42HEIKIB17cG2
47loL4ffSHItZlgPvl3O3THsnGkJlAvQ9ulWYFgs0Sf7M6OFTdEuPs5/7jVl
Q2EaUxGNAoZstZwcvNmiu19KMLhPB/5a+kQ0xnjWFI0VKLit00+W5NBm5kEx
tfid2dmC1ZBuJgaKXX+5U+X6ilNUzXWbZXA6d+AjcJyqYmBT3TQw5R1qqQUF
zVyUydYfFoRYLzdQ8wvGXpz3ir5JCWxXXoE6YB1sVpclxb5mdBQoDxjo+2bt
qRUBjLlvU92P8prMmx1XOKkd9kgv+ISveYPjQzyqSg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CaGkmS1ibuUk5Gfdq1CS/Mqy9ExBMKlEpORdWAWxWSEdNYXJGKbPL+Bo1uQx
kAoKhtyCc1+OhNyGvRmJdPotcXUCAiROb5hj/WNS3358asE7wT07c/RZO41P
kzemICuFPLpZ9Io/j4qQWo8WYH82hiuLsr4huuLQaSawbtC6adkmh18aT0im
V43FZqsCmhPA1xqZSAOAZsYlSLSkhArFKEqWCb78mdDC/MxK2YIFBBM8Mezr
1spnP7rVJ2Sv9K/a9K3+BEagGtoSVtWRn5R8Iv7CEDrEg3MJNEokJJQIqrwx
VJ0mSZkpm9Q7+dF7ONTDiumnE4fH162OTaLzerY2zw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pbZD5qybHHZHyxaSYseO4iqJY8RBCu1zrhG8ZZrv7WvsvGTBCJWAf0zU0Udy
ucMIB66ZOmsj5De87VkeQbEzYMQ7Z4pPgtw7ueVwSuV1RVY5di53MmZ2SaEQ
E6IyCuS4kc99r+zwOVnIv7qxUmKYuXvcK1h5z325aHaCGAIai6w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Wm/mYvL7zPNn3UNsc7wug1jjzpZbpHk361Jq+iyKyacx0VIQyk3fSGeZ9xT+
9vd3SqYbXprkxNM5lgDzyngiUoGHjkP8Uu32pdXvYzX2026KtEWhohgwgu7k
9j5xzi6vbm3SoIuJmMsY8dlWeUWGgzCXOwyr9JiwNMFzlAwCLTUt+uuyNjyI
Nn+6accMreaGLGoBHfmYQEc0wx29eqgFs/PZo+JEt9PU2N07wJCXmhHrp9qn
lVL/D5xsm41wBBzFJ1/uF8HofIUVADl87Wty7k8iTqEvzolQCgUoLIXWheMi
LmeC1FQYenmEs01ykU6Wcv2PcQDKO7IJTNDpiSOex9JpdeENEQygQXDj2xqG
O1ttn2tyglAOd7i6iyVanVwuXU/qQ6Zkogyd0Uz0jaHoOtpf0lmVlkBTWFdr
gvzXfROxcwQccKUxS96UpKlQk16L58F1ZzaICHynini95USiBIqJEBELdjKu
WDDJHyi5Ckdr0fZPQzOLR9jirLp2Ihs8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UmNpp73Azp6upkI38SxQssK8Jp3aOMSnO9M4egPX3BHbPJ5LvDTNIv4ZPVtT
wLNQo0hPjgee0wOjVdvbLIsbgrQFHxyHR0yHng1PqTNcOdUhVW1L392Y4YSE
FzjLd8T3D2r5MnUIcOLteiZRDVSl40/0w/u+J/q0AZBx2goV42w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PnRNuh/v18hM6I+RWIvDBlFkdR2crmy9pmbXe+YEO4zPsndCARAoiNo7N22f
22XhPh+YK6WMpN6Wl7/PyXyGQSOP1+AYH/dBdImDc/D3TmpidcmtqpoIDwoM
GX9fpB34Ub9ZyqVN7imkCUZO8alg2+WnDzCFwCHMaYz77E5mldE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15600)
`pragma protect data_block
F/Xdy9b/tfaVFg+Ia23pXBZmsmp9uD7DaX+79gMlxlFbsLkWqrSc88kYq6eb
ZwaeXyicLuVeC22nWePRTdLxHDOdJKWmD8XOiW5vezhw4TbhAviIHH+wRcB7
EMnUEoaepDPOQZF+o0ATCYHH8f0HxxYv1RvKehdevnsDEdZU+0uZqk2Tken9
CIj+fLh+ZbBcbEOPTFglDcXSd/8R6UBTvC440eBsjATYsrD6b/UaN3xUk+TH
J9zaXNv6+rCmS5IiMFPY0U0rUa1YVBs3kmHgnI1m4QBB1srJi6EVpAMlw5YF
Ct6twDqi3zJSI5Z8AOtDlvlqotwrlH8hqtPLNbjzcC/2D00opOUYdRUEiYDK
J3AK3StpGYv8jFFGhWvPhUllWFo+Ij5Svg1/58SHVUAVkytS/9ZUEgjKzEUU
vRlGbH0Ofbd+CbLCmeJNYXWeilzVpSwWB1UgnOXIcO7++Rt78Ru6UAZi1c/e
KMIVV82Vv6y6LwrAPXvL2SIEnf8DBYh6ZiWvbuAJQaK1rcnHIQfI0OITUXl0
ZfJI4Y55ctiTqgnXF9dHNeshdOwhMKaGB/bUdW5fauVuKW/dN/h95dZDmvzx
LqJRA2lFKVPJIHgwnMNJbsOW0/aiLmalOOlzmWwayHpY8Xa5az8r4FeVDMyR
y37xegSReQcEkjY95/8TqxuWvaPCBzIdssvAhrn34dyYPfXixrl42MlHaXrM
gsvVeADf6XCERW4Le+R07w8QH65Z+/mV5y5NIyAjkwGstQZEcpoLzEhz3IaC
cnvC7y5QZPWeL7YPVKEtr6734J7zsSzk46Oyx6Yx6DUQOR+dnOoI2Yoe4bL+
sD1Fs+d7lfiiR5n/MdOPw9eFF6xAteOYTdaN6a2nGwgdIcPaohc4toOpjTpc
/Dj8b2oz1D1EtjZED+gejLkRo1TWpcf8QKlmaIfjP//629OoHvUTW8tuXaE8
p6bSHC8ZEvOXjs8zZUxox+lCf9ARnOxgGvScwoCPy9ExpjO4g5d9vVTzLHhI
qPuZy6Og76OuRM+cnWn8F+/O/02ljwbp/5QWLAjEXAkGiTrLDNQM3uCIsuhm
nVYIqQ3ZgcRm9mRoBWh8ThWCHyP9ufN+ko/aw4Vzp7+nGhiz+sd9/fEyop95
YBas3UgIM6YzexCbUjPiUoO6nfGSRTELmNTp14lRFXyyqIZ90hrWDQPNVicf
TRpMcASZLQzM6IFs0Qj3riU2wlK0JA3fYfmowpKqHmw1CFRji3eW4KbkL5Pg
aq/txRgBhLZpXGqxC3DIRWpu9uPq2W1aTSV8VoqU9E8u7FnzTxNX5GNIq7EJ
KQvnOb4cFKhtXBSo2rAyht30vmAt3hy0y4WNzMNrWe+58NtgJvrQO7rVYFn1
CrV4ZnEmGMW1S4AHgf/FzRtl1gzSVDrqkMQHiXvwzjYP5LxR875kDKo5/pkS
Stt1IaxW0TzoZ3y+d0EBSdlTgeEKsCnPgyYMn6CcsVBG8APrSq7LBZHGmeHo
3PvnRhFmOM8mBvpslhbiXTEzH+HEEX1+KamNLkLlfr4M2u8EoV/b3sSv1PID
oEx5qqK77hTZQFomzczud1CXRZRm74luZaPDmhNEPl6oH921chcR9pL8GZ9m
3E70sV7cztDQFdntvKCOY8AsnyduB93sO3l46sRUwO2s6b4pkJQxPgZ8fZnd
pgg8o52idXusq7Pc/s+WCh9cyTQJ1A36jUa7ImRjZ+u0tAU2V6PZ/DiI7Ct0
jZyJuTkm6sQ82b2GmvK0xoxIv1lAAQsOlJ1wbEI1LotqbM0AV/McfmR6BAOy
nVfJGvTrZqGC5mE4um/gnUcZ9hbJtsy9NEWhS9akr6pNQd0WC93HfP+qaoso
aZZvElc4xMULktUOyaUfPz4NiUMJEYJfG8BGSBMg6ezO1W8ZM9qtTJtL9E7X
QwNAzKbKKjkFCLFji0oKYdStlFxdpg8hSmwQaFFkKR2MUx5TVAyNy4ACOep1
iveoJnM3K5lPDuTm4vMjT8BNmFguzXRhc7uZWzgJ8Zql0ECAAgDFm546XBjT
F5Ru0MIW4b8rb1WW9gqbQbeIyXOovAPBrK7Qle37wY2CvTWq4OR+TZHjCFNf
YdxhrKliNCaFb55u7z5MMgDDJTP7zu1/+Bkaoj4RnH4dSECJBhKOr2PT7LDK
k776NG3CdPtgqh8PNN+To3MZcLb+fpQC+QfJRnmF66vnfjBJGv9THDd4g1Ki
MIzAMhsy35nYUwqVeHufJnnDVzlfEz/Sop4PBEkUko4YZ0l1ExQB3s5qoV2Z
HKCau5RtNdzMbpyP3Y+clnlbp0QGEmh18BnFhmmUW8UIcVw+1513/z9YImhE
JVZcAAZCjLRY3cieVvHSr8nox/aBr5dAApdwYusZkE4pbgF62SY85SlkPinm
NMMQ5kfmzFA5AlbPvGLZfVRqEoYRR0wwd0VhinsPuUN9R33lJoChALLvMDBX
O33aZ3R7nhD9xTDAviq5RiYSaMYixtunXaW2iYKj4QLqtikL0S6OajhIoGW4
O4Mh7g0w8K39syP8f9xx4HwE9mSSRNS393WqyCpssLEKiicJ0Fv62Uc3CEAT
0Eqmabzeiadm8/aBnquAStMc7VAYYQXvHJmb2paXMi/TuyEVhOWH1coSR/9L
U6KWREkTX8YhEo4xLAxBHZqkTM7sG3uhqEchi1W/NhSoEtrHFEHakXtx+ekz
UOIo/fubZYSk54NZqGkES5Ix5V4Wtz4+LGQrQ33yCTwEE9VHvwNgBnbcN0kO
nXt4blyLBaKGjCaEIRMx48MlVCxOJUMkhwR6IZ7jdIVBlmOSvpKRXr1AIZxr
HxOYjvc0+GoMnfLpKIcMtVCyL2lskzwgk6u1naG4+Mu0RwExp8olUeZGZKfq
Clnlwh/RYKCC1GjsT+6IoFMTtAGHlA0dVJZRaxZ2I4+LrLR4NOE1zkOXb63o
W2zO4O4xKem4rlbeyllU6pqUaufYAcMvoKLiCKtLq1JxZrtppZki5FdyX0Vt
F5USECC8D0+ThVKzv2hdoDvLh5gLsjw1JhNwDXNIifI12X6P0B82Cjsnrh/I
/d3kiMVVxgqVrxJ1zlOQy3K7VrJMxjA3h3V84U5PItuNiLSGO0Xi2UInKP0k
D6S3diNz3bmXm/grsXJX9DmjDrrcNh0TKfxTdphzajT9NgXXpbRc0KPTFfdk
zCpdDRlZ2hBhtJRDvmbRIL2FuuTbs1rF92tvRSOAJfRcz8T3z65/zgohb5GX
OxSy56LsirUv0muKlpi8ll6R5YJ3F+ot7xtJQoBGeiInrkg/TwTRCVnTgUvu
tIdiDAtyCI/gdzyevdhCYuP2ZAgujsfADML+ZG/bgk/dFO1CWb1mIscXOhiD
wNTMGbMAi3rEAQBoavZszqHFlq5a6zNMOenz6iP7saRqxmTTGB2uYXRSBiLo
fYV9joWqzG0B8MHbzF8wbyOnm9BHooQc8fzGiZj01EF8HRW0GlOSLXN3617T
JCjsJ3gIOjwAi7a9nYNWKPYrg+D5HOIKI/sR/hwKJk9H7KN6PYjCKoImqUjD
EUMTqikdzpkTjct544PPRQ5js/Zo0fsTo1UVjISpNnKOKOZXkLLOU4OxNLqT
tmxVEOI+vXo544oz0yAnXXvbwRL3zGpDbcwp92W4Xbnu6nVVQoxGeLUmxGTA
rgoD1QFSG2+Q5aJ7PvMkWZsg58C4Na6HgV6P7I6W6mXUZABfPWvTsKwF3yyC
Wrvhbt/Av3drkO1awjEOJqrRZr3fPWcd/OIZGxGIXhi+Fj0O48iKeGF3hzel
0ZYHOovJQNW9M1XDwZmN/vqOPSpYkkWCGi71bWoPyFz4Kf8MQHAsvJCAVYmb
fcDPIWa/5scjgJNhegv28bqJ72/7pOStUCVS1Ski2Eng/O/C8BrBJguT+/oZ
9x4vesB3g88mD4M2OMapTz/oRrLi3NkJejmvdMQv5uFnETkQulP7ihHqy6Qt
hZOnSuDrsbQ+P6p3Yc39P4g+Czs0vEM1elb4Z6McO0dNMjOYyIlfxjpc06nl
f6oPFvGYSDyaJoN81rPSSopNbeQ6tS1qVhiEtHdcFCIHRaa4+OiFKmaXYn4/
+GauGyN2VIyFZe6IrzmRm4VQ1LRVtY68+mRYyxDwKCiRwRwxEb7ESAM8DfIe
eCIeMcn+g2KsVYXANTOAUJGU1z3qioHTR80rFJVdYKtQZPML5+5xWqJMlylW
/rsq+FkViI3sPEJm8qHhrQdZmUT6GCqAhLW/FS95IdVDMI/WD29n18RnN/SD
8j1gsyQcFVLwC3uf/JRv+RdalKB5C3UpY3JrXiBcsxgqBMCD7i6pPtTO6Qfb
eM+y5LMGYsDxWxWX42FCtzFyMqAqPDQc3u5lUOXu6SxmClDtuCXfIn8jgZi3
9exjnQ+Br6f5no7uYUFBYBiaEZQI59+5iS5ZvS73rmofxvQ3tOFhFAOgOhZ0
mBFiLhFT3rgZRTih2Kk3FJLbPgnag1VYVuPcwRHZ16DLWtF+Tpk+cvSfM3+L
dGr7HBkhzXthoKUFcZwO0DgzaY3Ir/d+kppqLFqL3eO9aPy5Sozfm2PcBw1l
8ek65X/C/v8GM+ZRqbQd4gXCcNtmYj8P1aexOnciHBJe1+YEP/UJqidKFHEQ
cdUGusMI9ZrxUzpFc/SsbTTo8IgNXvTg/B7JdtVglqX+gkVO94bDnEQQ9wjZ
tyQVgQqKZASzA1Y5e7qppjqwB+ijL0ib2CD1YGaVnl/lxL7ATNqAuXjbaQi6
4YN7c6X0eXsvyHu8p/qAuIhps3jl7lCsy3eWl/OA2IOMZzHg/PeTEDh1UKR7
pI/1znm9i0vh/KdnFsfazXXDUK2wbLksJLMHcXSPOEGrLLI44a/qlACt0KMS
vjYjCqE5CjAr6znPQfwezgQXt6eMyhxP2Wt+/7qAPNjdGIErSCMKPGKW9TBc
Qx/BC1bquI0gEsi8MmolSB+ElB6ul1NoHF8E2r8r3PFBsFfpV4m3xksTfIJ+
Y/W512wbA4RkZ8SFguummPfwTESKSiKiKMfZ8X+M6ksJ3Pbg8uanFirJ/ENW
gqt/kJFMj9sJTAi1i9hdibDHEDQ0SQ2MojQ1FclS8j0TXugC1A3A3YDO54Kb
KSEvdY3cWVP6t5J9u9Y+c3IXhpjeL1LYAgIm8Nr7JJb3n4FYpvsZmgmb2LAU
vB96vDkDbfhglziEHWVjIB/wrO6TCikqLd71Q7gs9mkmGRztN7LX8pq8PUXd
BQj1DzEBcqQkt0MtJbZDF/cKxLl8xPOw9iyUOZCvkTrbCHmzqS2mOh1JVtbR
ofrsUIkO5s2DHERtAh5d5d2CtAAgK5kQndUFtm3sNNo8Wh5khYS521Vx1Lnt
1C2ddQY/ZwnbK5ye9R2UzcR/JaptdzwttTYTWQW8ho2+MPfAOQqFeBjgcHdT
GHe9kfxm/bx0yDoYgVEery/sYuM2EhHFCQaUENa2LQZ+uor9zBFuDTGh1d9X
dT7Evz2LXKPA6m6vGIdZoPXhk22+2zdz4K9vRlIBJwEEpBcrNazinTFD7Z3m
uRRt2MHilx3I0Vs/J8eldNigr9G1BRUkZfUu4CxPm7lMfdQ4275F2sn6Xtuo
3VPAbnerRlKU9kQEenAI0uCP/Q7sjls2Qe/LXAjp8w2s6jAb4XpFT6FCMtSh
YIfMNN79JpKa5HlnjSMmIM7o6kviX8Rnfn58u8oVAxBUsGhgb3qhJYT7O3Td
jRFY+gT4aIIu9/1IM/798VWq15+kBjuhGah1FlNAl5Ib+tzsur/4YFUmSUSL
Yo48cFEZ7Urjnjv7ktfwaeIPsKWsQ5CZTCNtlt7+RS1kbdZHwXLNiAa70ngd
P14o9Besd8U0hHXxeEc40hai5aKKmI473NUT1//hYpvXQUdTkBs6WZH8Z4LA
KbO/Jx3fMAIKAbGgLjHc65z00u6m3EM9WRgi59/KnhytQi8sYQZfVuap2Sm6
miU8B9oXT9jv49OswTbpHG041pKeVKBJ4BzpkGS+vFDJxw1UuX5RsKno05mr
Xdvod2eZAii2yEY6Vu02MuqyqRwGHIx8rG6LOEj0dZYHZOj7HZhUNAmb5v0H
tgz+0upqD+wgrOmF16Yy4M8ZcKJKO7WA0K7a5tqDdVTMz0SQ6PjK/SiY1xzu
IvuPr+VMiUSPY0UnM2heWcBBjdHWXVXHFnERJN3uG2LggWyok2ksNPcRxkdC
X0GwqGjYbr+BX7B+ap0UHhr8BHD2a/DpszZ7EWQU7Wbsl5/eBUq/0r0IDe2C
LebORRA/Qgvfej+DC4z0qtHxK36Gkl4hIPiZArWYwAxnfoxXAxhLg9Hcr1LW
B67KWyoUPJI2Tb6JW+t4tIDiLyntcLcgr010xIccZuzsFXEHhT38Jvpi1mJS
A9cikZl4dRFhW3HNEEEZkhAipKl0EqWbxE2mjOPoR+nk6tMoTEwlNu3/JimW
yMuyPze8TCfYwlQpO5XlXoQ4yS3px8pqbAe5cAri/TB038TDbL7LoglzFQel
746hco5gXxqU/dM0BBjNd55aRzioIlIGMD1P2jrWDwXO1vWYz7kyu1Dsb2a5
oiGmd7l5oF4mnKHKEBfl97QZJRsHkns8uJQgtOZ9GXoc88WNOIqrr1DHp0re
ol2MjRNYWuxYFqrSZd+Ggii4+rQSHmrDSt+u6/RikQT+BmrrXpTmHVMbDMwk
+w+kIL26yiEdIhc+tOOgoQClEZrntF3uIml4ushPBGXSUVpus4r4JjjcJTEO
2HGvlshnmVrfl5/a6SpQWp3VQOSZzcHQ/RcS4rqUiRKzHvCP6Uae7MmCrUGD
RNSQuuHdpE6om/HZSROhQ1GIpqkTOj7HfBRiLNTTd+jC23vVwNx4DuW/n3NS
hy/b0bK7FMtsRVCn/uGr3ZLGHyHHF9EzAC+l46YGCT7dfc5Rn97ijhBnDmrw
qw3XPXdzm3XRtSWG69JHafDRf7hAhmASAyRMJLHIZm+jroWAEsLQSVcc7vJT
kThmZcIFXSK5g26vB4Kbgk0HznohnNzisdV9Quh/YipZDugOSYpu2GHgaP1O
5QwbtpWk7KxJiKQTU+eDk4rGBv2TniocNW3w/z5iaPjornI029q35wwpp2YV
fiPf6c5y7jkM4LE2rUccLLRiuOA8H+5043M8Nji+y8co4gZe7JS+v5Cc+5jA
oC2Mk+FR0IfZrc3ynO2YmV+Bo7nTPZrkHbcLuy1qB3aT6Tdk4jiqnoBGMAJU
9sniaX/rtb7l39Eu+zqXvquguuyppW+HhSZn2t7don8DnqrHjL87ODbqjwv0
Tv5V7BEFWOhFgIwHJPl+R2DhQRIqw1jLOsLkGxZ/bgupKHe6/7YZzFb66cTs
tpJgeFdVtSQyRCGeQISlyzpodZz1t06+72IcDhcfbpWlFHebSMg/F+PuWHUR
klxAs2/tyWJDxUeMo8CMlGlB7mzyuW4wQLTaP5VA5Lh+hD1j2QcdjXcMADCV
GN52Iln0zSVT/Egoxx79gqakm0kIfZ123orMYzt9Ns+dkHkj/5UiqHR5Wlom
aBFXfeCqlDbA5rEMriOjeRvkKA5CKivx0RaosJmSW+CrLVwLoUVR6wXFYkx7
WRZf/eohkF6m2tvSRhV8Ou0GV3J9tCWIHXg1zvVaTk0vO7HwfMYa0C+Kvwl9
WNnmXjzuo9AB3r+nFc//VHfXAFQao1vZcRR4n6MN4+mhQFyuPNLQ7J7CsO7F
lJCXJAsVjGIQ7xturSyZo8ixcCvPYg5FnkbOjZsYAf3kuY0vimN7LyV9UPnh
WwW1uiUd4r+k0OsQ+Rwy5xdbhQ2UvwxWycC8bjX2eDgbrmpveSBBK6y0Jmyr
Bpi+jd9XN7xnLd7y4bs7n82hjGh8C6xr4SgM88nOXNyLnIhSWIfKPpWqY6ac
CapHw1sbdeTiNmp9LkNDgB7JG8dBfrUIhBSBCWMnRsqyRmYrt3ym+zR+k5K0
meBe53brLKm18VDe9E/MrJMoWiaDXiyo9PNE0hs4QQHXu27z/28wtvhasfs2
2FZJvMzgaUI7sSPid4kXLJdtxZN7bOtXbcB7Uoc8H8QoWuTOnD25QpxJMsEf
rQ+BYm8LP6lbRtit30hrrtwY5Ght7QNFzsa3h8ce+jtmjjyk+SbDhXynN6JM
nKlpbvLIxQXo2GpoJZk1TjzttI4YU+8h5dfR9uosAphZzuiV/9FXpkNJuD2A
JqYrYc3cyVsto/lDQ0m1SoXZLryoxtsJkCwvIoskWJuMZad7vMoS4suyq3Xg
oatClgni4p0G9vg8BWF01JU/Px1qpde1BOE/+mxpr2wLlTNKrF3k9sTEmn7c
pGHHPannS/yv3f8XEfc51OEkeW39OG6pouV8eU30is4MDitRjz/vEtoNdcrN
c+u+Ou7v3up3XpKLKbawMRip1iA8JFDaQm6uCxBYGq2Yhhxezzi7P79MfMuy
0dXKawwOlaEUDS9xxB3vavAcXFOExCoOf2Nv1o10JAKWWfePlLrcjmsCgmHY
kjZMlPwcpr/tcH1EFsk9OgHNLeCdLVKXhVlxQOHZ0xhqig79a8J5EysndAaR
+YuiQiEXTRl8EdA0J1aRQrwxOcdXG7SyfaamLK4duJNJG6VdzEM8UCx0Mkoe
NrLIr8Ry1vxLACKRJhTF1xpD4dN1wYytrqgohtqPRLxDPrSd6srCnqGhMVmL
FrF3aG9iM+/2mWCu1Wa7dHUuJdZflGyXUqDzrXAvh7p/nII8S9+y0NBTo+Um
2o1XAHATdtTIp6F0RJeFu5sJsJIFOw1TS+BJX8rveMZ9wN+8I8PyS3IJlOWf
EGKqz2Ilq+RtXTdee6EVoHDl4+eB6Wnpy0Dun7CQAogWiO2HKsShpw8m5gcc
JKLKYdYMPHx3UZh5nW4cO+0pTLqE2ulM1DViEwsn8NGZgBl2nSTDxzc/Htgf
0HeMEtPbRIDK5Ou8p6gqmX+aAHC+5HOdp0AJEkoFnsjMuD2LALx7eISOhpqF
ZhiqxNygXw6gDLpled4SmHG76oo5X8MC6/ZPN+qlWFUh8Cm/hGEstXHeTXkD
di5z0ti9mGbpqTAichUEbenf8yz2Yo02VQT2bOA3OGVf2tk3MckZ+DTphIV3
wQEdSJWgaUj8npklbijJYxqt1wb8vBtMcQhzvToTRdWfgMqkNAiahI7UYbhp
J88ERBHKWyGY8COQt913B1yIzOyWd96yjLUidVvQv/cIUMVz6H2FlDzUFYUA
YoNN3Os2s+lKDuc5CwyZN1vuV2jsbfuzcRd64RwkGmgtLdl/PPrn9/z1ZsIV
X7+7QQBKeKGs0PIJAwsljpDA6opoB/S4x81jKfkKsbDkYPGha60q5lKsO04A
T12h2wBjmxnLXpga/Gs1W7ZMUYvZ6anTlq7tWldyIK3HZL1jpYmiBzklK9BM
pOQmnPtv5RfE0CQL5g+2ai7cTGZ0xTGS9Y3FqWMOaBMX9tcuDN20xQy6Sr7o
rJ+a9/RBbuIZ0w2ZgCpD5oaCBjcvXscCqG9+EsHBPEMbcwOcnQbqGQ3ZO2/h
26IY0u6lZZYlw20lIBigxcp6uy1R7KQ8iYhNAg9h9GUrahS8JcqjxvF2uq7Y
niFFtk5OWaFP3l8Dn6u5WNt49Zhs9mzU8iuTH2cVrW0udgoI2qOe0ZPld3xL
6k341QoLLHveLAbYbyhcMat4xvV0IF3R+vfXQxRFahzuhEiuaipZ7N3yj4Fi
wNxPiN/bjpyFSrUK87s18D345cF8ZIrE1MG5u1h/ImMxykNQJlJvuCV3O6qd
n7LEx8pd7kR3THt0IfYQ1bkmgZiFnUCUl8hg+gOEq3+9JXcAItVLrWCKwki0
jMG1DQAvG85/houbqrg/sEnjGHi1DaV/kSlrmvmSpYNMCp1wdCBcmhmRV+7N
wtWuUyKTvZ4TpLQehD/vguGc0HpUhh3z0q0d/hiWQ049aHuJPMZ3N5NELiPH
UGWd/+Iu9Q/9pSyGvSBNbqtHMBpeaGfvIysLJaNJ1Czn3klEjffFJ9avdVkz
MVSmqkKUxC/VxJqMgHJn+MliDkc1pRsWTYgRSVr8+X58fkINqhGeSJHBGmAn
Ja1NVePu84URXi15Bjbcvlo1OSEGKZsXdKxImxCAF5msLv8qf7RBWfMjwhDt
nTUhAxom5fenkgetow+t9WXVrW3lRSgIMLNZZqLW9GDTNiGxhPz+r7XdZi7C
+KF10kK2qrBSa6fiq2b7HtjpwlImUnA7puX4DHrPz2iJ385EE8cyu/3kQAoI
cnANnLOAP/scqsct8Ht4GMwFg7ebaisi4dCDxc6rIejouAkuOjq6GNJieHoQ
WEMT8/wz3lahga4EWPBixEkU4XyqhsnPwIW8hS0cpPEE0FNOvxiRBMuUR8bW
ZKtsT3Rke+2Loosi2n9JqxFXSuNW/mIANi+8TbBsXAfpu5zrKOPqFon8hyFn
Hj8GSPv9Sl48DF/djTBZynX5nYPyswYvfkKGs2cW3OCjw41i3I6FBVxSYwPt
00t4VKJ38s69QXK/WyOFXAa3z3IT6kthM1CBbkXHqZqOzJMTbxz1bEZTD7vB
6p+6wj5b79UcH6o6/LPoQIW0EDTfR+PGx5nt9eM+7BWtqLrR7p+So7aO4KLv
52QfFGFuFjmrR80ZfVUOhF0tx1PrTGCQ9zXRYOR1FZdxFrTjv7VYOpUy6g9i
/ATOl5ePFx7o/0IMfoPxKtUEpIMyYVrZEZY5O1S57nTZ/t+XQ9/vIbEuK/wa
8i1oMipc6JjFfNyA9OJ2HvfnXfwgVave0GtRIrpAw0Uc68qcrErcnBPtdLmG
T87y9zYDp1sbXwvQqVqxhEx3jk/V+EeTgcnJu+dySj7TSA8KamgQn9odVnCp
Em4OC65uSrbPI0v/KzxAAOjahbPZ30putbJLNq/yLNAJiPChvb0BRWxBWuo7
LtAyHgIOMcRefKkKyOwcm63wbRRpaXOMJlF3M2unFoNO8KQmduLlnSRSCYuz
3pPTrbq3Z1dBVTf7DxLhkNot1NKuP4UmFOqjTWXUSC0vXw1gkbVwlA8PhK14
fyivzlZ1VoRm5B3eL+QAW4ztrlVzMu9u50+n1vAdhMqyC8pqK4f+BgideiRh
UqwRbfn4wEhj8Rl2cUxqEABvJzxtwHyCtxeHHFZaXvtuUYqfkpV1ZdKpMjEg
7Y+oB506984H1PNChXFxzf/0Cz3M12l3fa3OcmKCYux5Xk3mMMJ+TP0AkIN+
0xvfgydvbW+tCktSnJvygmXMr/Hl5w1YhwblJnyu/YTXv76jn94YlsitQ1rm
kIHfJ2OfSXhpmtWSh2oJnHwZdpn+WyatLR1TxSgSF5qaWheSBHDXBEaXMc9B
p2uDAD0WoWwK5PPCVFgJy7nfgeLIJfx3BTOCH/nqkjasb1dK9ijQFMcz9mpy
IRsijMEG1V3gI8iVRyKzl3R37DoDGUQHAMyp4lLcej70pBcrtNAJs3VfTt9U
mLOsRESS/lrMZj8zWGsztdMeQyznCM7IBpxf96da3FTPsQSJhTE3xFBqVzdC
2WVvb3ngDAPwSzKdF5OAMMW0Ym62/yj/ro5RtGmaczYTl1y4HAl/BaXLhjoc
JIz1wcu23X8sslK9rioODcp5WOSaL9R9O4kbWGzg4g8o8OYuj5y0ubp0y4u+
8Vi7MY/F9ipoa9lxR9sd+wMD+rjO0fPuUpN0AQvf0LdsACxH7u3fZg/N/Sv8
F0/95/dnb+A1ue0Lz3qokP9DuismPt0g1AXIbkqOHxnMh7MjXibrl05OPe8/
kMxnQb+5/0dYDEoK9wOW7xoe6MX1fHVJIej10c+TURujUHPo2iziovoq/3A+
XIuAr7lfhkjGiVH+qqnfs+MUAZviiDabJPmf/rFDwTSoJBjKS+TrqWCjTkYD
pzPVeq9ol/7sk/CoNUJTE5msFtdikKLfl+0GxmKzaoEfmzTA5prGYsyWovwx
ad+DiznrgQuZb1P9MpDZJZlEv/nnlnoB6OvqDw5bbA7tAhfQ7z9qCH/Ksa2r
ZDK7d0yZUIRs1PfLWXBNq/Ax7V3bivHOOGavPnEWn1YIuf268ObOjgiuPhea
2fj4QWHacDj9xke8i3bKZyz4Obap8LeY3n/SBp8LJhzMsfV3JGh4PHQBBed1
fUOppZJ0r3k5SGgfukYfY5GVXqEf/Kw/XW6rN0QOoKFQZeJlnwGxdU97aevA
o4ekSDGtmy5J5alABXXY+QsU8Jh1A0CgtuJ8G2oNOt2nHRxTT82HLFH7eqmc
CxQAafTCnE7mSm6vR5mYXsXVB3JGpQN1VGOtgFm77djyR1Y9lCZZ01eNFpfd
FZckg9j2tFPjUacM/z4gU8PBNqSlZued5Tm2710JX6oGqnyal8C7vLFrc5pq
3TIjlUoIqDC8dgZZ7wZD2xp0O1uncZ4ZWrBFzlEB9F5cZ9hE9nsBD+kiTsae
lP1H49taDGIRnrF1VfIPoYKkXPQJepBR98rnHKCIDfvgJzzidWOreSOGGLpY
7NT5jma1bqNvpcvM4pG6LaA9YwTAQOdqFoa8wLDR0PRQn9Ll1TwDRyXFZlpv
BrOTRFdBngEgjgvZkAHE3yrU1M8dyoEX1jMn3Ppd+cjtfocbyfl4oxAGw3g3
l6AaJhe4LmhruMhKyBYh+ihFOmawQl0fOpCuo7lSNTs2fcfw7F+77fKS6i6w
EShytZ7NItqOW8KeHtt7bHzFi/gNt7cKK4ookFY0NiTS+2yxudkNozNnQ2TL
nFMra4qSg4L/yUeVJ+Y1X8ZfpO/SLyJt7E9VN4uqtX1k64YDJzU09Xffe0g8
P7PGyMtz+9rIhj3PqXvlw6aTsuMSeWpFoYsAxzQ60w16WTaG1hx24wU8HGsZ
SB8TA9hKOqQjIP0GK412lKd7V+l4dzQdaTQx0XKkk1GjjuCdhsWniSsvXvYl
FL9jDTnIFDgbd+NTSaLRFuoKY4bgzsUS+bMNtDVHKrsYUmXYS8Tap0VlMJhJ
x7Te+ybY3uTQ+F7qFxne5VXF+NxGJ2N0eR/GftT3CCkh3mGR0ABtsXQ1sxoD
ZFlc5b3dwUYHLiTUWirfxw5L0SJGFQxGLFZla4RwkK+uTKeiM6pQdVtpmMxm
yOjjmKxOicysda2lyLLyA3sK8cLJfzCUkzaOYvUncEqcZGo5IzFxkinzqR/j
5K/Sop8ysuCTL667/+aXAT+KjgDC4oA8K4P4t+whM4v20CjunvMj09IB9MvD
KFSIBj6Lfo6Y/zRJuADEGtjZ3PpGlACNQwvsrk3qa/QyTLdz6xrFQmFtrEeY
jMqAUXBtwWW7yTslv9VmXpwKb5jqYUP6MjcNBkbasex1nTiGYokxgzpIN2eC
7/UOo91qlghyB+JZNQzPiOFUyj9LMNubTKuhqCLHJH/L6JOnILyVQx7D5Q35
RFPS2LKftjP5ptyomgPhEPkL9239aix86AbCArdYwdLwTEylWyS723EdiY7+
53f9buiwlsa6m+LSUgl5x1SvoyMNeCFcUeWTwYeykaX9Y1CCLAw9mN8ZsyY4
gJucUU6dAjNiFgMzzWqmfY1GTMjXFvuUo4or1jt2Aqak66QPvNJ6AWkOjkn5
husTkshRcFB2FXgqu9rQawx19Pf436et1bEymZh3yrrkaJXg+sfPqM/nyled
MM+MAnzBdS9fYH/5Ry7dg3DqLnPfF9PwxVv3/syOVqcMFLIHJptUnQ6LPd3/
h5bE42FU7BFWhGcUqsz4aWHwMgtyvfRVnNpibRODiv21QBFF2CzZ259lcioa
rnXuXpbYTft6bC/KWaEqADaYCoJUhdFgrYIcwrf5ZlqSvVyWfLSR1naTa/Bz
N21WAKsBs0Y35x98eviRMquHO/GTSSZlHdwewluekaCd9h6jn5yo8xRSp7Jn
95BvOIOvUR0DytJcN1/qBp2qEyu6ntKjbUfIN5QWgvxQfpUNVBAAwxngdFZP
i0qwlm9QifQXV7BduL7Oo7wjP3ZN2tG5C3UOWk2BYWU/zbWKXHR852H2w0t2
qJ75GmlfQ8aAXNMDcI+0kCJ45oSB2euEaC2Y/SUB9vm2B5DIDjuW63M3wthq
Xh77dRNQzibrPqaiq9SLSEbtq01zA4af51wNJgPgrd49F8g6Cn0z7NUWYVwj
rV3mF3ZAaZBJycFuzK/55ftrWvi3Q6wV/AYVrRcynfMdG/baWXQ7j9cwmvKX
1NT5kmNKDDJiUpUHDWkfMQphdh3CLQRBcBBS48BbI6H1SRjWhiEfmDMYIGdv
5RZTZqt8xsVb8WpKOs7cIonceH/Qe8NrcUaXEAafFNkRnnEJ8bJdXLvNYJXs
kaGzyrno9d0GM9VBdlq8x5JqHPvf/AdYV2LQX6MWLrTLeUnPgS/4yvn61TfY
gsuVjO+XYbn+yDwXw9FXF4XlFbgf53w84Q1SGbnNKeigX/5I/a1H3lknvke6
wun2O6FkwS/1+oQSOydnkFYqcJmnOjTYShYELlhvZaAQmReKiPUZ0JiUf3O+
KqEuhhYfi0RC9V2Uur2+mI235teA9Sc+FkQ+1f4wss6l99vv8xwjz8T7dD16
G1OStZDSfbMO4JfvqUgRGGsCEuEgv4sCwk9KQkCL86NnYXF5Nm/+htn43+W6
+z3NG8koEJDGu+eZCYKwj+Mmaat1AWYfvUBNvbrnuIS3zb6zLMDiqlXQu4m0
BjPOd6yTRG3aoZ69aaf0WDOg/qHN98Ozy/IfoK3D+7zUwVRBLqQGsCPqbv1a
E59XgeaNGrxErpMdyosGLzp7GcL3ShpRFJ5KZ2jOQYy92MZDDOrluNrBYuNl
oqJ57IC2+BIrkX+73mGvselXRY3SXOpWG2BZ300Nl5K79K69ovrxhJ+ebvJ7
xYiw0nWWMzqA5kxC7pEXhDuvIwabEKmbLmMJLOEnz6x6dZHKh5TAJEHYyHzZ
Q9B3WWWopbv2pWkP/slgOAiMCzwjlrNtzScX8pkGkmKEA+t3Ge5ipLnrMXNP
A+VvZ+rd80CrjAJJP6IP04xEdmGdQ2aMKwj4BPlBDGSPfTcKZzEV5Q+mPpo2
IDlsxtkxJBrJUtMIOP2kAOUxI1nVv+3C+Y9LbdEPsf8WqHb0SkV5mf2RpJbt
8s17FBc42VBEDwzYs9i7Km8AtrzGjgqZe/qo9tNEhFWJ+4BR26kXcQU8syq9
BcejXH+yGLLggC6KdiCr1Vc3/7ggzCG+/fj2TaSlxmCcRJTQJWlnFfUchJda
8ltbtdqRjglfLa04MbGPF1WW2CdephMHQwORcwkYFeWUjdYdLK7Qw8NYE5WS
92dYKaXaC5AwYM4KxPPn41K6Bc3+BgKfXPXXSFOoZG9j5CYERUidx0NASX7b
8mdT0gOoyEgtmzwITJD2z5SVpsTn+G+c19vk8PK9hFgL31oOrhVolRn8pzY3
G3X8+qChGMQNBIXPUXE/AX7Moy4mIWW0ioFmVMMoklYhpgis8zTBfwWJmrFa
XyJX2HXS5DZY/wOdnpqwALZ0WSnkkTVF/3ogqgodX96hc7hv1N9Wsd63Xyak
ds1/rE4H/nRY55lvhv4DsMwHz4hkiM1Xgc+kwjAJcgsj40vVB3RS6lViGMPl
kzKTwI1li9g1R6K7LvkknRxLZaQLxlZkJpBPTOgrP32dSMKAxzMONbJUS5oX
Z/koBpcsMCEZczQ5E7Tm+FJoxF4kSg7BdXzA0XleVfaZKsOxYKAC/h8uTTrD
he+d1WHafoTaulaJi103Aq7FS65alaLM54HrAIoL6jino5nWmy35NjpeGQQK
0TWOJniyGJdlxU8qkSecnY/6UAAsN5WA3w1YS9F/mKsuWoz1CzT/rnpeyUGk
AKt5V+eTqRawh5L+L4sXWshzBp2DLsni+3krR0Ogse9rieNolrQe/H1Cf40p
JfBp2lqgHc4vEMD4czx5RC2Mo9YGJiiZolT+gUjgN1MZNo6JLXLtTe0+R+kK
Z4nTReNaBi6WlFZdF0NcPxXlugt/RIZDz3yraXFcWeUZgKrJj5XvPPF8HFZ4
Wq5sl1uhPlijYe0jN3dG4kRyMfnNqAZn/+Ct4FLGzYKrUUkZGnK1QuHMQS7/
0Q0C1P6BtzkzL3DqHwQiiWpCNOpI6CRH8grtFjVi/DYdXLquUpiW8Lru5fn9
I76364mDiAY1MTfYyUzA4mLIvPlqm6GBJFh8Jrw0rEw6HORfJFKjEi5kGK5w
gkUfk3gV+pIfMEpKPVe7/SdL1kfF2heA0B3EHiXuDzI/a5ehy85VLkWkXRYu
ibFg+cp2StW445H73uuIkzxJR6F/+i/Ui2zHJBQ7HE+fMazZGIZHlYLRAfCY
1zh2LxUhNEQppeJdhxutfNciFg3M1q/xsNbeDulkagBhM8J03KvPjP3+4F3N
b4eP0aEKw6/wuyrEsC7ugwgPv64EdnTDKez4h3qu9TC0/cWMZMP+w/e6w5p1
kfzqwdCXXUnQ6xzcHnhx7JDOrRzsWmmpAX26Zd7NRhri21zMJqlaGj/np83T
4XTN6oYJ9Y6Iw9Jz+dBznvKl88QOWjQw/PMvXIxCLHc+WdpGg4/B5baS+aPQ
412+4dntITPvmfJ7MrX64MchTjVB8h3Ynw8AJRLmkXetrIZjeIlUbPnfPBI7
DSDYmDsKRnH0vbH37ujfL7os+eWb82+Y7AHvGgxFhuhjpTIVunRoxYZaRSWJ
GceXgeq62IaRixEC5zdP0Cc+VWREudQqAKrIdVFPLL4IyEVnDwFNqmMsCRlA
PXLno6XFl2vqbE9K6fW9qROw+v9qtKZ3hWGHJJ22rl0OgsW4kIXktYHXBFZM
7heeDgnzVUOlSa9d5cYbGq9Y+QtPFfbOaP7BtqmZpWjNmonfeTgY2I9TC8Zr
GUZMDi1RO3zqBFFEIEkvgL5XLPmCPQgrp3CtFpNfq2kIIlvw2ISqo1K4guNF
AvA2z1VHkpHh8KERy6152txuKOd+/UVRfLtXRmOybUNU8AtLNL6rWgEA8SeM
u031VMSKodgISSGg17O1QFUwyD2GwmdL/IR6RSaU/kGn1S2jrjxEkZS4GWiS
zypEoqux/yf4oLak0B97yJeywhsAnu9l77nYrWGcSdjbaOlZ8AJ0eAhFkan/
849uC/y1tlDAR7nN88fh3qQpXaejf3ZXAxMkZH1m4niFdX06ieWc8TuQexi+
4TCRzMiX0SBUEW8qGXl5NHV3N/A1g434cqa3BZDrmsOtbSjQ5S4t0Ar+8/5Q
uo/A2Uay9A43l+oHAiQLqMEp6Q+ROraQjSUS1RNrLzYRytJ7FM/4bkaX1lJP
nmatZcCF03XLF5HIgFASxOLHWiA59VSjpvAe55AmSTVD2S1pRWMXYEaWMKZ5
bGZDZugc71RoNI1av7H7RnC5RAlmJzXor7l3ZW5po07j64QQ5HvqOH0JNLdS
4coiSFkv7NpM8EDu9B9xf8PYj6fyg5o2A+WvXf7rG2Pv/xjpLwuaIYXE5TRj
xJg6yBN1xdhSXbIlZAmXOQk/Y+fZqh5mLwrU6n1RXb8oWwclVND8R7MxTMRl
7f9w0LUVwJtaDnWf7y0o59tx1uE/MA/Z81v1EscK14doirYTqHVkl/YEdW/4
QojZtTKpC+3RitPQDA//zp7EXbzAE3CBzg1g9LHr7fdtfzhiTs0cC8dxddbQ
iuGWeXktVA21aOTN20jynTycisLvLC5xt50yVfEcngu/7Q6+SiAxLlZH1ndY
Bqlrn8VuYsFEYyqS1hzJS7Oidzr+dYntZb+N/zIV+Z5RW+pq5+5Sg1HYKFGR
zjfzRt97WKBWVyu2lXc3rlkWsQZLdmSlMyIRYFa3FhsCCT3k7VB8HMelobBx
2eCb7MkSqbK1b6CKKUQeTxGMR5tXwo2cQs19gg9brvW32jkK+XtDsvdVQhLI
1NV1WMCUcHzWfMOn3vUY2mrzK+CBRonLZ2yChWieTGJIblmvhz/LyFbWsCEV
PeKCyOzTnV/j7Uo7s1LS2SL3X1kx02MYnawpTZqyLYQc32Avf8bx27YeB1b/
UMZhWqscVH+h4XeYcW2MCMAJmBI6o9KNNJTTsV1AClqsy1zhk3cJ9qxAJLw/
g8qnsDwy8Ld3wl1tOEHM1f9lgJrahnq1IVeVg0HBiSiRpP6ezEMceBfb/dx0
w4iZFI/6HXR3hOmS35+bDvxFNclfGwwP20vc9ke0AChFoa9ajFW9AuTDhgxK
BJI7CFHesR/9abg2gYNCuMx0yunLaDEVqgkXBLfNf0LsSyzKWsCWJYjqKRPE
spO70GNgC8TSki8UqK4/0MTJyxCEeVMgmc2GxCOSSF4TzDotLmSggVWGaH3p
xC6qZt0SBFJpU3A5J7FG+b86C8TzIt45McWHUk67Y1sfhAZHdzwWjxBscUfH
PCsjSRiNDCrcAQytO+DAiHmS4/NwVFV/0QTd6i8zSCmc2vErJpjBVSh3UV9W
3OBvrh1+gLbG8Ytvb6PIxwuIKyYPiHNTVNJUTDWtwq+saOu1E5enngv+Xy9S
l2M6/mFRk+XBKCHtYejC6JAJFOjjJuejct4Wijq5pNLYIt8i/o6eDEOZf7Z1
WE0uFb1v40WRtpybSLNdw527BZ3CMvWnEl2RCympbxI0YC+KxGhS2r62oX+G
a85Lss95cjMkr4uILfvkfEKl29ypXAZWdpNER6yoSvDwq0EwvQv0WCzMg1Jb
dEf/WBEumaBrL6Y8Hopy0WhiALuAq+CdlicmkAcVTtpzQhsfZ7vxH9OTvrIs
z5g5EBY6lY+cuQR+/Bd2anh1ltRYUye5b3f4vpBcipJQGJ9RcRtSvoFFlr9U
yDuVhp8DMFCMolpdOuwR+H9lQTH6WbYNLJIaHnHF2tGH8PuF3VhkQUbODHaq
Q70hBqyOrT2eZRwewwGkXwYIlC02jJR2aTU2rcRxFJHeUIim79usSRT2s38A
5PR9wACiXmG5Zj+jTb2eMKmhdIq8SNIeVM3c3B4MFmA32WVO7gVDy597dyAk
rTta9lC3ro6spAU8XIgcuijKOrm81Gp+qLgXM2qJSQCFnM7dWZq2WRDrIv5x
KRHXiFy4JCA+xTGzjX7DtVn1rpNsA7lBtmSO0CvhQGymOzBrktd7NuDSMkA3
W8ogmBQdbBuKMXuWlMS/3evxVRH1SPogb34fcd5OThSlYhdo9Ixka07Y/Y5x
p+xHYqtXNE0ll2HHRpNrkFaUi0wrIrdEa1S7IiQUxV1l5LW0skw6neb41YGT
9cTYmkC7OcUxFzvu0roqIpyqZxOyyzYH36bRPhFUF0oY4rhnyAvCvQ10gGiD
1ERSvOiIDO6vAbvPWF09kTZnhMnfCyMbOaZpcVqw4PShv2YiIeg3u/tSgNSN
K5ubf/5R6LyRGL49/4NsANehqPDoztLE/f+zGe2IFdNsHtneGMTrP7P8ozhE
ZfqDrza6Kjiyca1jBrixwauZWVxDRKDzJ5cfoOv3+Rz0Ko5DsaTTCuJCucdl
yfKqzGn9vXjbY69EPyvsZlymlasbfBvnuch/YnCcrpiNkj9XEvz86xFcuNR8
JLQ6ZNFtRkBYh8N24OyyhS18+5vOBJN+1eK4M9+AY72cD3l0u4U06X382D+X
SqlGFoUEai9fnya/YiX85+6OVxqHwqrXqkRZZz9gNfKsVEP+F8KAoWML9EXI
K8UGZQnVCiTfMyLpazhPbCpSHm28muP+GNZvo2lxM554WS/T+gHpRYPY9VZ6
rId8Fi2H2Sfm2hYVNK8+TePyim7I7DKUnECGMvG/lkyRGTMG2co9xz6JNRhJ
D1e3kc1tyufkHsPLDfynGbX1i9/CS06PDNYwU4OU6ENo5fLFBxQehnDK4kAf
FHdiNXl5q8WjdudqaDN96v6XURtOs7nEvEfwQuEUm809797kNcGdktzNnJ/6
GjjDoYZaERkah2cbZKPSVZ7RNkPiuY7e6ex3wy3RBdIoJW3ZsvP0fqxxIzux
+MttOSPqTZcObumeW/ngly/wioO4tGJLJ+T/aDsebJG+069013MpZ/8H/jfU
NgE1ChyHYcmRrMk0t4XgB6VK/OArgVSlv3u0ADol5ZXgWuwcfZbB8yw9k3qz
7k2OFsx1BZisgtY/RNiOht1hsXS3i98BSWXHaaJqU5+lWu/sIJNhpuetPUDo
s+WRAV6AO2FqSShy/ZBat4QvfY9A+M0EhNsu0t+nG08Ix5ZSjK35XK3Jdyrm
dkr0I2bD3T91oZqU2NfUkXDjJxU3Bspp/wAIItwFDxicvNtWCQiCQlqwFjec
20WitkR7qvHMIG3Jhl0SxeLPY75lVuBiW5iL6nfysES+MRyKD/UfteVx4Zbo
lZjWlaKB4mHrDQRIkgJ8+APdg6+ftBkn1VDLAdIMykDHPD6FvZn1T1VvNf/K
vgr995qROUBgzp5vbYo3LMhZ0b34FLB5mnXOtdIAu3iaVeiD/aZvjhBR9jd8
xNr5q1IZKfpZYevS3DVAWYbYqeXtpYnRTViS+lmf2qxo3REi1xTSg9Z9qbzG
lBG8XOMsgaUOD5dx1Cw0Grj+XaYvMHFk2QxxSh4mlBetVRMT4a6Nsu/rqStR
M54txcc3lXxmXWeFwB5pzaKwKDf6NwoEavRXHzMkO8ZPCBI8hRmZ0teOiUv1
5kmqFshMpg9+4t4MWUWsIUkGg99EvbxuOioEFWk/iAiB9iGR4067PUPdVklU
Lj5uDQyEzcmX6Fq+5lMthX8bAMcNRUX7j0WyehzAIY46yrMxMNFTF75MIPCQ
+FF3VzpT9FmctKlG4f2MxUhbFJXkcwRdJTPfZSPBh9Viv/Sea+KrxaAFhN0M
V0oRZ3BXhn6M+K9H5aKe7O+MisQBwFpiU5qWia0L1HXNNZgWGoMnXDrA5HNc
WpYYQ6hNeUdG3TIAx5XwbTxMDaR8mlY14n4z5ZGbLJb/SZtZpXt9Ia/IzHLT
JxojAIrav1XCVkhKipbu9HB4jeQatSkdYCBLYp0C

`pragma protect end_protected
