// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iS/h2B7vueXO6TXgM5CU9ULlBxbYWQ9N1Cl7OakzF2W3LQ9BzIrRNvFSicla
uI+RFdJGl6rnc7492vX/i6hVGLp9LUDGBkwbwx0Ak9ByXorwaxWdEOlDX/bt
3R1XPiglkX4etr8dQx4wp7nX9C0VTfe39t+TxFEyNpSiPOONMu0QE6fQZgzC
mL6DBjAQZbTPUXFBQ+va2SSTmGZwXlVh/b9GoorBCufLn8X2kKrMqYlI2emN
2fRzdBwY+CJyCb6kKruGzaJE/C9QWpnPREPGN0M3ERY5ceL6mlFz1VQl++y3
DQj4ODReDb4uVb/Ope5gyvvl//KJ6GTp+f7WY6YkBQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VdbF+kmvYwvNS/z9Xml5iwWGsMCAdXbFt7aOAfyYrbhTn9rrd9uClHcZShpK
8+NuthFn9QXExGJZzEE7nia3OXqaPePMkDinTtyVwAocYQxURHcM/zX8u8kV
VuO7NajU6sZ6JIH7u9+kdjAZ/T+eZWCsvJP5ay4JGn/G0sSlJWp7mCCo5vRo
Asm/Cwhoq4zBS7VLV8auy/lfljNFBU3XRazftsG24BPh26vj9p1dZdv2IYBB
fnIyWnAlgaPhr3hd2CjeLMPkEV68Pfw7hKPF5H+FAxQlXofKoCiAr99P0XHD
NB1DBbm4yUP2KLvizGWIt7sARXC657sFRito4JRqoQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iCZ9HnSHdI+yEMZZ2r606F/MojEGr5jCxJ3er0guwVXlFKRWN7ZYGqdiZ41+
kLK/1tseiz+A2XEzy+FVOxXHSwyj2iIOWxPRgTNTJHMWoimloECq4755wAue
k/GoaxhtMrAUi4nLlEUNro1DotGtl5gJ+odOpyNaavzf909GB5lUZjqvqSCa
sSh7fOIiGHHRLhoKDGgI7a+Fc6cm53akmLycxH8V4aAqlYYGd8/rRN+06th8
IQcAfH8IQ+V5cxwWFlanmuYh2UPSYIqwWz6GqzPq5tKzkWkt4ksDAjSQ61Cf
eUdZVzJW8ERdpGGuBc+Yqk8YoMSL/XHuYZOXO5WCYA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MYmxODL0d20fuHtZgVUXge83PlR00mRrwBL6WMGnd3F2jCGK0Iz6s/6QYbiO
tQI/dJMNmsymZTVMZwJD0LXRUEddG7sAFSHseUShMKWIxy5ActhpwJweP+o1
1I6EZl/0lGbIyPYuhvNLSI55kIBJG6ElIx1vCe2V5d17cf5v340=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cN6BHOe/IDNZxitsbqNo0ROwt7vnMwUaSqLqf1f59fbNGZIBb08k2hmgct/a
D2KmlbIolaPWjQOQf0lj/lH4Jvlt/qO7QGFK5eY3oVvqH0tF+K8pa8zDQCbJ
UUaAQfr6z4QkGek7CsYIlS0W2g2oo4ck3eiBOSOmPBads53aTaNTXKM5F1Sb
CycB1ECTHEkNlTxY76ro68bk7Ee7ckpHAnmJxhwasYCa/zcOHmmR9x1NzOBk
E98HSmuxGW0ASTeNTJVvIZdcATacFyHVVRXTRN/hvdzhBe/OxxKPxlt+yrSL
f/fF+8zYPTdwwXGw08x3U/gHG3GxTXYAJ/tcMyQfjYCUSZ/Vq8L2iEEXfkaA
5mAw8uifaY4Jxri+TAQmU0MkYBXMAQnsSWnpgwE1fPapVcFzaHbcT3LDDnfF
UulpyRivbfMjANdI/Cm92K2tKmDp+HDpuc85zveV3gHvyeHp51b2yabVSL8x
uFHRAeTnd5OmP64trqnaRL0BhuvEVQdq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PZnhzfOgcq1Yhxh2pANH2IbzTJviNi1sOlvaNfnkVPnc75sj0Y1YrpbZwtnk
L2PpK8XACe8U8FQqZxfF8f7/4fikygO50vpeOc2MC58MRHEI/UG/3cz/q2z9
6hAYgEu7yi3gLNq6tDD6eSNY8OFo6VAyJVf4sNMlcttDKNX3vPk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g59bE21KgA8ocNwdK5urU3MBECoc4kWIDYOW5M4kehU+9dPrsKx7iZBEIf2Q
7ItJMg11LbaDJ2qrWIyBMdr4yXDxyo96K/rlvZyLR9gFWpNLuAHsghdoTt3t
11l9XMoDE3rB5uQp2UbXg5Dp3UISx6CKbqgl+89RkowkmK9dL/8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12512)
`pragma protect data_block
IDUCV6n9Uu1RTCf1CZ4ubeWOTKJz/tUV1z22GSMmJseDFvjLitlJmhKz/2nY
zRg0EOYXMK6EFuIxDiBD13Vc+ai2o8pb1/Rs+KPFkExxWLkvFns5sLP0n99q
91GunLIL39mXiLHkXmSSyhlKO1wpmzdqBab9BccEHNthcbY9nom2LCiitvIs
n77NxkpGcW1OtyqPDyUmAtahttlCqfKjmKkbkK67ZTd03V+LWgrXEXSQmoOq
hX6eP2K37BcnViVrwYxMEVbGA9uHD2caBdwm6LH4kFHDoEnaS2jn9V475BU+
38eeIxFC7eXd9WfVr/DL3ecp34vFXQL3IkU9dxONV+YCwYjA3SaGFukJuG97
WwWTIvYsE/8OOwWQoDz457Wh6wLux+vkKJdLUwv8JpTIYw+ltQ17T7gqxlZ+
LJMc05CczprZ17ZKRYjQfINJFdcnv3Zs48ZWbdcEVx12K/U/5Dv4XWAo+TgB
hx6TuYlbf8Ft76+lPBwVUzFK9u1uAkwLt27hYR5U/SKcU2VPeuzNRTT4XRwU
37tDgucFtpxGkILx6ePb7M5BMrVeCAQhA/Ha4Lg10FU1S0wKYeFTFmVPdZlt
6Ec1E4MuehtO7tfWr7XI3Jdbye03d5pMLuo0nlDSkLrIw3GySwEtWdr3unyH
f5Fd4ly/KjMclZstDN6M0aR2lTYYZdlZFgbTrkp2iwnoKJX3sHpVMnjVof9g
+Zi/l3DWqddxbjgvCM8qqmtqIYukoWjPjNMjMLtGuyTEvkk9+mb4azz5nIGh
F4oWbBcx2hUdF4T8GfJ+MyqO3bKViyA/rv4H0PRJNoQjOVg28pddgZn/Rm+v
cCYJxr120O7QoD1WVRLQNlmElY23nrFFa+fH8b3mXqX0PGfeTqb2fBtrpm4+
1BF+q1XQgheOy/FRl1nwNAh4LDtdSwQbcrf3dbK/HR4qAQvN51inR+tgfjt7
SjsCQ3YPWDQEV8StTCd5qIbS6PrKoecNUJ1SD9LztSAQY2jCKPag4UwK0lFX
Mev2k1HSyS6txt8RIWTG5Jf1VvppoNcD5ROMj9j2APkZcxgP1PR8ieT0W0Xj
5pGnzg8U9xTfIGHCKJF9sXK/FQJESvxUwLrc73OOZvKo/fVS7g/4GRr5+qpx
WVKpXSPGPC3vdsEOuntCBErb5JMplp3IlnFJE/AIeMNtmZGOm15OE8+LXYda
/vX3zMu5SP+Hblt4tgm9V1poxwGX18bPDfah97Kg5ezv71Lcki2eFQ4QljIB
gkzmgOblyInD/YsMikibDdjNUEjO43o0XcN4M3Y9F0XEJOV1++t85PrrgILh
m22ObyeaKkiEYAsswSPeHDUNwROS4wYVoi61kxI91WvLyMVXNoFwelJnJSdT
nE0ZcXzdqa2Uuky3aLR2ZCmmMDAt6D28ZgLQ1EQIbk8MwpNIjGQ+q+dyludz
SE8fEn4sopaXtFdiC7gmS4TUADF1Dwut8RL8EKbs0LPsBlhx6NCkGDGRkdRd
noTkqpCA525vS/8X9PjLfBjSDwJRQHFZ28ZYX1OgaYEoF8Yi+FQUvqX8eHlX
NXKM86JXqjCg4A/k5Hana+ZEe5ZVj5kLOhSA92NVbZtLexPLDeqPG3+CxPaD
12eKFPNoyUHB8EjT9+70Vz2YSkCxBByb/O1QLZ4bUs5SxheUZcXZ61aCEn3h
ZfoP57Yeu1fWItiu1SxHCve7VyWjsN065v6mUMf1PmRpasK9cfHo795UvvTJ
ORWZ+2JRs1Wi1mGhvLY0VyIEn19RJNJ3VItN1eGLN4ktIaJj3vpJC0VnJgT2
J9xqCV99LFwSdqNLz+hnsG2tUZEzvt+xnsZbFZpGUMdYgu5NwdhEX7/Rd3OX
eKS6gHikchSgjauMSg+VJYhuayqzIYdlf4cxl3xRZHBhgLo7FrQ36+tXkTuK
eDiYNhbuSF4nvIj1X3H38UYH/j8BMesjfcmEZoLWviZ0wX6X9ajN7Q6IqvUY
/YZQla0LG4WZQ0uHx7LQrO3oM8hNR87nI/l+0PBA3KU0Qd67gOMlo9Eu/kiD
hftHp4uA8PYEDYHNw9xuBlyWhEAxs3YKXXgoi3Z0Jq8MK9+tXIcm35tOQcKu
+KQIPXEu0qqL6HZDIxpd4f7w8lKTNkOmdhWo8EWgiAvFuqLHOaMiIrNPQWck
lpejP23h9sbJfxMqKtk0ArWmBgHFWS6urWuL/1XBykTg2VzsJUvYCJIFTAeR
VXsMrJjY2kCiIX1adPdUW2/SH9QqSVuD7tHPe8aT5qaVaph73DoTCJ2wJjfA
aMAEv4GJZrMtDXpB9DuA9TPCkVRD5khr3FJ0DafmxIF4qpsWtlLCTMUDSbbX
r5Xvokn2XqRykr+eMOOv1U2EWwEt84c032w74JefdojVeNsTfUErxupzW6c9
UwzYIfNfPkfoKHlzT/yP6YoJYfPuKG0bi6qUBBBehm3k/wH+Ua6AHCMQ2TBX
/UGdbRvxhEXWYUhbEnSWpm/2ajX3Nx4d6qKZEu5xwOKRtWwMHdcgxi9uW/GR
lsnVL2sAZUtrh6nkGB0wOApT30Ok/tiCIDlgDYBgX7j2M5yi8WcEiaJ8xWE0
ASbq+xF1jz/sN6y+/N5LvI+iATDIzTo5zPrsUsKshEFVrto3YqgSjP6rK+HR
rupzl8FhKwN8IsVftsMbzrfuhCgIsvNaNsAgxnNU1BFQysCwylygQLqsR7A3
kcrXMUkvwIMtrXy1atplB073UxBOjgwzW2iSn1xuCm6/AdIhB3EiGuOwTaIX
nRVjv03veUrO/A38hb6rhr4pWshjr9Zl8U51xJLK0MmHedxqJscCo6uRZPdn
XzTx3Szp/AeJEINE9usi/a1p3nI6Wxl3HV0A2jqWPGrtQrPeu2JtLsr24JV2
ztdW8N+hSwUIVTOGwr68suKsse5q0OIjmkSJdfZZvuN8LkVpGn20xgyne6cb
t8AjExYJvBgfB/XZCvdeuWIXPIw2m9RBqhbXjQ6t51/cfyfgoCd1BiUCeqnj
37D+3hZYsno+EZZkBUR/ZftRvpngLXy3PXqne2bkWoNTzFTCe/5j4YKlvaTo
g8XXQZNxUjPQ1Bvu2IYXlyeI4SqBD6/Jk+M0+KqUbu7d4c9bKtVnvnSVGQE8
wd9Q8wIkNiajeeb2FmJUKl3DeaqbHnda0eAUqawi9693k+INPKckhzHq1UwQ
kFG0LY+MdvtuQp2ZeBKcWKSHd5w7XGHrc7LsjkIm2yvDC5nKracCP3ZglHzF
vqM94cXd8/89ytHyQf6FO2re7O0QhEp6h3mYTMMDO+tXSJILpadIkdRrn1yX
2CeGbvpAUxnx9kNBOkpu2Lk87BG1g145q+n/wZZGr+0p3DnvkG8KgqNCFrSS
aYJi196ht8Gy7Nib8AXkkdeKGwmzonaceSZvKbTwhF6UX7axox4G7pCL5GAd
/kebiA7XokJJzcR3f9xb4SrlKEpIGaq6rU+CUcFWQ3F6adeD6wVFVhv+sZVL
fHlsigKFKfQ/GjqOKyMkkgmFK9IhrHl2af3aAkNPD8/35RdP7f7065NLajea
3IJeIhCA8w8JsZPnAtXqLldiIJ6korgahlGk4057RsKnGQpTPvqf+Op4xxNv
6VMeVhffGpjXxloZpijxeKhnPt6/DeDnj9dI2M6qRa31B+8SaVHndM7H6SdI
RnPmIy5+hlDSSiEdAHEb2+P0m3Uku60MjvjMIdusMCBQhsaVZFgFR7SexMyg
FrbOLVbNjky2H+TDLseKHAw1YSdDe0mYkXtTmMUHshfFcVfPl5YKkpGHqbOb
cgFEo9aDC03gpjMPYZU19i1TSMEVfZyILJx+qVy1Qm7H+sc+Z0FxisMWc4Pk
V5uVkz2JTckgLQj/6nGfb1MqD3uGcwsCqlvZZyqBjUTTTU6t8Eq7alGFykeZ
Mn5bJtzWj5/7Ez42PbifYflcroF03Lhp36Mh8j2TmU73Y5NDLjP5GkGqOVKV
okHGn2/YYObd6ucvmACVjuANNJ6MY3grKREvafy0egTEqyu2NlpT5D9vKDkG
FN9ZZzunfo7VPi8+6OZtBnhVG9VuIP4oy53vrvgsmF78pDuRBxGrWD/M9Q1j
k/ZkLV/w2ZgqjQODBcHtoKY4Ar0PudvxbLEFzKdgLHm+OE7/J+KzNnTOQ0CQ
QTwRpnIw7H8NgRPjDGybiiYjN6kXpFRO/O1/2xWoFNzUn4/KsHSMvTp+SoBg
Rc7f1gi6SSPKOn+pvjZ1V2KrGIlAt5IQMDZheCyV/lAMx/58OUk5sPMaupld
j44rBwKpMFOrcMrQWVkba0IdehrxswILM3a/JqV6OhetdI3LSNkUptKyvfb+
o3bKzUdm+rPbQY08XIxt39mtNez9bbij02vQby7B1epdVVY/O4A7+lp4TisR
FSZf0sNj0mrgasItp1+YD/VBEYeoluWtZuQSNrNaHNqIpPWnPFwaCpAqCG1E
NQZN+4GpWPrZkU3jF+gbKiBOQbVp3zFbnXT64Ze4z5s6PceB5C26vrmzLIH0
DIkm5SPdxmpnvQfRta24I2ASOOu/reE6a7pUogIV+MZeEO/+RfbfRYThTA9i
l8TQBwrqXOJ6xBEfDiYlMKTgmPIE/Aph6/9/gins/3DuBnVwaFgSwUULb4h6
jU5UyvxoGfgiGAGY9doJyiel4gqY05doq07CtneXdNUp4fzEsC+q4LXnCaCY
Ra+Goo42ABhJxBi7sp9dMEv75GNLigLi5ImaMWivh3qvpFvfuyIoeoi+oNvX
5DTxBO1++FmBvi9EnKzpK6J/SYMzAYHxPnDlGmmK4sN8Fr7WxlJKUDPceYFw
NHTrXGG80Aqk2XzSgbzeS6ITWTUUmZLhirt1NxyEtIzc8vjs64k89fko4n8U
SbpzSvu4GgwpjLV6D7lGVLYby/b/YbaXuMK2hp+fzXD0Zjq3Av8bi+V2+A4K
+LQgWySs0bTzuuY9YhNBxSj2WLW9VcThbsy1F50o6mg8yqwcOYStyJgVyNQf
ja87QG0iU1hm5jFXWqwnNihUZkXpSk99LmuipFpg6vBJo+GR7cit5029A5T3
SHITXtKYTwvTWTWdtMN42YwMAv9So6saz2b2mNXCldyO6Efgy9zw1g5Nkk0w
ud41DeYtYse8ZNf9IV2FyxkPwukREsWuwi2xXt7gTcnKV5YFtA6AcJdRDAxe
fTo90LbWWak0FRoM5t5HYS5lx9gQnB0ydKN6hTI9BDKAyshkFEQTQP+kE8sj
ZQPgxfV5evDjSaIzexQPQWY+toGP0PmYzKbhenMuqnOi+Xd7VDGAch12SU6q
weVRc/C922ll59IHwL4/ktjsSB+FcytbS/fg6Nf2Mneq/lv7DUzYNNHYSKpz
pN6EsfkpVdB0rderWehb0cyISHLvkloNNP1M5aM0P5u4N6DfAOA/XdcXFwYn
BNmx4tZb+poK90bhFqPC3WFeXx946VjMDgB1mpwqQgzTaedRFWkcT7VMVBVc
iC8IaC7P52YNk8eUXiktPcZRwGP/D0wN+ypeNCbA9NXciR/o64Bz+XC2OXka
iykvDPm2jtCeWETZdZaLvUsJr3wxzeSG/8HOqwypm8uaaPP6DmQNl5vkFwRX
DDCmn7A8LTWtyA3Bq3yVoNhTOpov/Psgr+zSr709uvPReKd0uYdYrFxPBDO+
kzUIfh/xnQT7+iLjpAulObMM0dHe5FCQbX6FD/KsV07uv2yEpoxss/FNAS/z
qZmxlHMMHa7SaKRotn4Vrr63ryWzc32+WwXTujPxydObolvNj/XzyOfIcgH1
ZWWX7ptUsVKoKdOMgtXXDt4RBJDufWcFGrSH47aQiwQ8EoL5x3G0oAfzsk8A
TrLrvbXujkumR4VSykE/VQDiCcIIrmBDxKjLtcXW86xh7ZbF4MyUMs9uty+H
qUz4KtxgRS4qfbcD6LeOKxaInoXeRZO42HQ4b1VhJ1L8HdK+Y7pJ59NfOgvI
FI6wJdYvTzFfkutOlYAyMahVvvOlx/lEgXk16dZNiQBc8uCToSokHXimdoGr
H5xoL3iCRKm79gf0nmINkU5X4yuk1IoPqdTJdqUN8HD9/3O69UC9YwKeREex
ILZnFRPDzOM4cC5GRSPo4ji+hKN4q/Ce+bxEs7r4ocaB1E/A3I+wjQ/e1B0o
cEAiv23XS/6sO1QUyq+8ArH+GUeq7xtsdwMHpvuOGwI1dsMKMKrcjgiZXmAL
+voSmTeC8dUr7VslPI1MUS5ZOvUWHxITIjJUlIkojw7W1aWbW5dwG4fgXspO
8kIsdy8e8zVcgGunnypn+VAyZyXacfgQDnG6NAiroSSAXeRm6pZp7sl+JKN7
UEEADeGDoe0vmFAHrSHC69CqY2TsX3HAPbQtyD3JUR5zuClWn43ybJ7e3qFW
OJZ0fHRCleRA1CY/lQJ2ew4rj8iOibJASKH8toHf5uUW2UkdhPNQ5x+ahzSR
ZVjY72jSUC6JoPOkQq6aUnDjKxTyD2pjxvmeiLQ+I1RI25ZtmQIGbT6cGDFh
yBKEjzaBI1HPdB5ZVdz37/IYT6hwpYAgoMdqt66IXhp2aFQb5Z6b2EyztCQg
Xk1fj15wdr9jayynyBQC6inqtwDemQYJY/KGkukSFa6S9d5OrAluugVn+lQh
qo9trUTgHtCFjA/OMcwFHYwxTqs6sWSQBsL+CzFtld5+hrPKjGrmXXNceA6t
CtSjoebR3RZmXHBw99FaI4ILf2hlrkMWz85oGvYU3AeqX1wbUSbm6rdzOLtu
6Eirk80hIRTD86Q0oS0HvD3zjrk6y2wSD6mpsjRW1EdIY1xzy26VwgOKgsVi
kuKsZCaA/VApPiMBxm1vSm6KSFuwGqhjcq66zMBsbSZzmN8RDFXUdeEtv8KK
OW9nc4geh27MiEUNjqhRcfrGi8643obE1Ny4Dt2W6ALmtHWhg3Vrnk6Do7Ye
Ftkjcq+SdnmrpZ1PcyNTRiJpr7ZBu4/CIQt7MlwthkCIKOeo6IcimfE2kOvH
a/OK1RylZ0a7k+VMq0q6cbwDsQgv1FX1ByiIST/AQZQEcuimE3w5WsCEKuBe
PrqvrEbdVA/M23QlOInos4BhOJKCfTJ+9cOTeJkyZ54v3kRN5LlB6GwVK0oP
Z+tBRKZZOIhS9/qGZA14zA3FvKGOKdaRCSPilRvb/sFJu8nZfRk200SDQ+Cz
mZM/HX7rkzQ8DqrJ8At0VksjC1CcGkO3vdIbOZwZjKveYUBonRPx/x8x/yhl
Ka3oKekcMNvg3n+FENuyb6Eq6Sjdjzr4NqFvHbOvkZghNVJiouv8zthEEAdI
jCTRQKkBJcuv/QLOF26oNHvurdsI+b7jugzZs9ehnl5c11IrvkIFs4FkmEz+
0cJ8c63ZwtL2FhcVq+fsFUspj3N28Ry1h7zG2AAW/uzRka+5J4rTAyGF/5wC
6a0VKuz+vDBap/lb9Q3cxBV8QO+9UNMELKfypOsOz/9Fp28Ov6AS30a6QYUS
TyblkeC2o8RUrOIDzoFG+1NGEUQ71TeAOasE1nbyaRpDhUBdZMJFuAD4tWqB
L9+c+ttRv4twM8ezsJFh9ZTgEEnGALl3NksdiVvKOHAWz3Nx0RzLBqfhGUyW
NtPEZ0PzdOF8KsQ2eocwcAv6kXxZ5r5bfSgvqbRMg3hhyWrXNVmBt/LFWYpE
5+lqTw1Qzw0q+ggLenRH0d3u3Iipk0uX7aK2aPadogjWS2/nO26phZdPVlEB
Zg6r5e1Nqt+f6kzSfRcHZeLkBF9DoQSSn6nvA5QCoRzwsMXTPuxBj01XKUaw
lbzquRJqdVJG6xvDhBhJwpWLvDqkL6rarZu3zHiLsGhM0IB9WRvTeIWMifpb
X3MayxAzVdJkaa6i79HFMqtgoL+0WzSerHZIAqlKTQNRTwOBQLfNwNdh/pG1
K1bH+TcBxQ4h4P/40nvGWxkDUQep3ELAOg4kCU0eX2Ej8E6yNrEuboGwLW3W
v7spM5aMWIrwc7b1c6sYMA0XiiXfRCKDiCuOxpQ4WP4A7IwPEmj9XgR7HF7S
lga2U64pV8WdHRZ6CyLLd+u0pnwsXSquGGSJq7tuS4XYhuqLTBEpC96SXjQp
37IG+C7pwc5WOXGAD08HkAPYnY5buKEnCDNOG1t1uqGfQMkqCbRihNCC5aem
Fk0zeaJQlzQ6WKLTsZLD0TUVXdE9BuoorV37T+3xR5bEN3VCzl43zl+ccDBy
xAJtirn8proKoxOBOVVNpju2pFiYLkTkadLYksIxE6R9hDQ1XD9vYmXVMopv
DlQePiv7wZxN3EwGl8cAPazgiDL1896DxRQ4Xl7dHe7WZqZqH+MmPBzMdvXe
CRCFxZgY+vy/awdoTrk4n3Irolq226wwHbs+zAGD/V1mLbvKDnAWaUpJXdJZ
cBeE3PL26Uvl6hCjcx0BIexhg7w19GmcP57fiwby/ZNsyx6EWsDa0OM4JLz5
R0u9vnbaiyy1gS3YrVwmR2El6mXFqJ+Kk+tOi4f17RN9wZebqvDEH1HCY98S
bLPpGpD/6UoVWdcw6b3ggfFphvQ9WAgUjwmQH9GcUl+NskRtoMM8I6Iy7yff
MAdEIdjThrp94Fn6H55t2GSYRwfvAOLVP7EZaEltuS7q3t6gCocsdBPpLdef
NLjxHy3txXprRc7usruj3FczwdkKxA0tEe45T++2CRRpihuiZyMYImo26xCl
G2erAQD+CZqnKiY2M5BzMygVlcw0BJA+TIHNmDPlIVX5Cz2MzhphoIzHZmEN
ow52V7GHdfG8BPomcMTYMVzcSk/C8mQULlnUlM8HYK+Lsr1naDoYHDecXLvx
fJT9R1XxEF9Feqj2TiCUP5NCwCUOD7ivm2pQbtRvPrS40YQlfTdcEuwyp1CF
Vum8VOTAHWvalii2JGCED668PF6Z8DKXEUpuSUcNoMsTiGn9iJL7XH10D4JA
9Y0YWVlPSTp6ThkcWsic1QSIYn/wIuy8VyLIQ3tCxTD9QHBv5mHKr02+Ir+M
H4Pe62DDPK2IS/04Sc/9VB5UFhdZQrHKpFLUpppqh2IMPie1uBXmdkQfyGMc
pIjHIxVHiDXlJZyspdxQtVTTKM/7US+5PPUYRwPBYzhjySITtZyrH4pMV/bt
KQhyIs62uD7Gq3gpTUTz4iN0RFwpqevsgEqOXM5CjCM9mmbUZ5US7iCBsQUP
hLoKFBsh624h5eMhz1fCLXp9Npro+n+eSZikfbdd3fNR1qNqoZ6FY473LEwt
Cstm9qMcFGpLL+ma1Yu3adZQJM9Z3d6+pXlVyRuQGwFjpSg9/Ygbwk/D6jWl
T2cpcpAOZiusYk+fkJJIVdLD17iVBuYtltomBuXnTS9VZTxTWbN2mvnl74vU
0ZupKMBinxKP8dCqteKR1LsPCiCWoFCXAllBpEDucGuqJnDwr6qjaahN27OQ
tBhwePnw13mLUh/wCVtW1PGGlgWPQ+7PSMJR1uLbDLy8xEqFl8DN4RdYdaPg
B7qUJbLIAx0wu0HES8hxiOdosk8iawAdO6cZ8xx2wP2KzsTg3+8efY3d11Je
ku8O0N+rO1kN/sQdRdnR9EzVOwUSLagqi7FBNN2OHFxQW4wBhkrNy9++hgdk
Bk1YXpXzMsyq1dmbktLtsy7f5EOMXbmDaNrIPg0yNphvxsoAaD3AWgK9sp6b
UlCIR/Ynx3/7f14Oi/AASN90cjChxvVy6SwWsSEzJjZApNsMVuTvkBDY8m68
6ljGf/30gCpsGXh60NCA700wQCTy1I/VWoD/1t+l1a8NC8EnvH+2ABeN/OV6
iFltyYMeqwdgZBnm1cwXzBiLDRqO7L7Y7E6gSu2EuVz8wbFL6g8QDMKhtp/j
OAtJRWyS/PgMGzVkKE9HxAS/9qSLDn9CNVgPuPtHQJN1pG4rOjNWIFIUiT7T
RhaxXgOTTp6zbd/VICVHNTPE7RccdTgK5H2JxFxLSpoHNKVTg1oQ3bGlnjIn
3Y4HrpTZuFKkQQBETzSRyD6drlXGNkEVKzMA+RY1jfWTCv+q009vTNbsKpsr
8w3hN8/BjSXZ0idqlvekR0Am2McGiguXOEpkYqx/EJEVVHq76cJbHVakOuZI
2+43/+YWdH8/Rvxjmlot+joc9SH11GX47zgMoZCw2aaVzRyK16v15MVL6xW5
V27er3BU1I9tOX2u0zdQccqXa/e4nHa6tkrv02UzZZ7crTFDSG6VdSLAHirn
259dB0wVZZUU8PvmTY4glUaQRPlQb9g2xFpZoQGzI28RJEM6Yiz9nYn+DNh/
qWJ4//tX72tzoT2vYOphiGxxOCjECjFu7n5l3sQal5Q4uKPR9YO4/FeisGiv
R7IJWsVLMMmracj6yZDPclit5zvaSQFdAjC1oZCGRsp+jYtixcao0KVFT3Ie
Tf3VzmKLXfL2YsU0zLYzxgUGbhrOllsBcfQenjqHf/oa0QyvX8520oYFm0oJ
UUKSgq6daUwrAghrMmgV1blhwbKPXwoOkle0mEqm42JkkyHZnGIVM8EL6AOx
fg1EKiyvt8007045hykNzSv3TV1xkv8svAbPNj8eh/DfEtURb0q9GqLWEPSJ
3PZBKtknXl7wOuy5wBgzToa//vL4St8zWpSLeccqoDk1g8qoG6v04zvXvE/f
3dxPDcvFuAWW5RCGDqmYgvhKnfx3FyhtvvZz9jGKjooBzf/ho6OTReA2kEgC
WSd9uFxCiknSyXAqHVM+dyDneYlZEX0F9d0TSartIQzo3zzIBkCgQw4AB8go
3aqUa8eCGFpbHUnhIEtQ1PioccvFLALSVtiVisTyawCCmMaMELHl0kwruf0a
VLNniml7FjI8b8ZLQxY2CdO7udDH1wo2MVLMdZGam1T+yS6CKEpUeDjbulp2
cy9O1MxtFTnlLRQhXeVZBAavxJVpI02Pw2Cs7afZX1RQY0t3D9W/DP90c0xD
gVH1C3yDlPomuxlYqtgw/MkuGhqC5d67f2hApBqSKjB3H3659J7t4CzJ9GZd
SaqK97BEJDZGkvAzJGCremBIUwpcgveSPRtaAnJiMSdMVYGRZ1DY/2TKosMT
1OxVZJ2ySl2B56LQoolPST4n3xTlRFKwYUrMzpTcY38ozeRHMb/pxJOg/g4j
xF1/lfNaLgWUanPt5xRLsnP7K4jxiJlnTSVnZS24mBBiRvDD85KZYqnOG2Rm
CY0CbRzJh3JY4/3JlNIUkQ1XVwI5hMLOcH1d8vpZM7VeeJR02TuUv9wXapkB
pHSLh3MQF+0Va1Os+yM/v2oaRHAEYzCeH+bR1GzwdJzB70F3Em7ytxtuxIEc
MKZ1gOuMSDFIaeQ8mJGP1Dt9RJF9mEbh1RSSM77oIYY/vGnoh+vsJC4E94hN
0WqXB4/o/hbd9PvSYTsrEV3AqsIxKnXbyMKRToEhaG2U1X0Ew8uDE839CugT
8lHiEdzb/gV5ZWC6VJuxEMbfj/yFL1W7LR70mUSraCxthM2jTlP07lz4BmSn
SJxJVOeTNDDAiJxGHckBIYDHdCSbFI0ssg2f/KNxV1nKQAURSaeIcDbSZ8CP
MpWZk89OEJYzrR0QZQKavhOiXDq9CV33icSayTKDvA/FSzqb8EYOL4W1Y19+
jwf88ySTgvDXf1SH/T3GQjDEXXWYedvqxiH5vTXcjz5QYOOpyaKWjFB/Xe3N
jAL3YUyfKDeK4+CwQsEc6ISBSmEOA9tUEcnk8e+omCnrBjU3NaoBqcP0y8+5
r0C852PfHQ0/DtiuKkBkDokO6youfxZQAXd9o4huqvSg07GcE1Pz1fE4TOkC
raDq1SaTprP3GTZf/qateQ7/oqfuEZAoz0DkMDF2PrO38v4xH5e+RiHuoBm2
1tUZdxqRjR8F3fkF2+AdQ9Zmk/yLHLaBBP4YPh1bl7YJKY0p/vwR+JrscnVP
babAqe1yKSvWoEQo721ocBtN/UH+uL3Ru33vndjwS3arnxu64zmpd9oaAfzg
pUF0qbZzDF85zpWD+9X97Bj8cyoTAL7jkR31mqaMRGxkAa7Y9Fv24+T7lL+1
+QCBc0QpIN3nAisd9pF6NPUBlmF71Nk2ZrsKUUcSCFCVZDgzdqVNc74HHm9a
6l1byDX9OHZ9h0JB6udgl4HE0srXik5pKRf4f0LMNsiPrLkbw35PeIqXV6TZ
YTPEXMxoyjbob6bSxDvi88rLdMjv/FGF++XGlcDTAkj5GGtZrMj7cHTxWqMq
91+XKgLD8YTbLEQzqTaKTG6WjRe+AEG41YSCZhp5q1rOrJiCL6Z+lOg/ywqn
agJOx6mgAFx2wyY5++WbmYEB6GlZlzYrX/R4jW+CCuGPvqWPdrd1RET9Rc60
+qqYnoL8lnHNQQVT8MapwurQ8M9ScYqXJl5cJyqSEBJ060UKlSDsGRezsDGT
7UJcgDftjt/dQrl8vdyRhvqeu+R1ImKmGhe/+hsRiWTFVVq9sw295GsGXGZe
n8paGuP7REIujXQQcluAKErf0Zx7SztwPChcBZ4uOUz0z4j9fGkikfYVSWsN
MxAUID4RSdvVtl7+vWJbS3bx8iG9edFa1ZLX9a0nMuAv9fGAW3FdKE/66MLs
9XSOBO2ysf43KeW/zKKVLV04uznKQgqFMqBen2uWMmc7lt9wo1spKIcjQ6WS
c/yabO8bcR2QuUK7k8hKywcnfZEc3LSvqxuyBEpotqnP5ze/bqaHYt1gq8za
i4MQwXZLOLLZL09DMrcW/Usp/UtxCK/We4pCu5Zxq1SObOK8K53KUl/z/KO8
fWgDb/LBWMnwJOoAY+QZf46oUR0MSp3ZY2ZcLGixyb2/Aj4EcKZwc1Ecvneb
ZpPvkBvfHNBl7xXTu4j7XD4/BPuPcDZrZOR4V//vpM5/FWIJlI/JxO85lgVr
DT+Jtt6Oaz1Qp+IDVg6mNZbh8MzsRiTGz31EZ+0bzf2uB0jZZfcc6z7DETIA
fINA/u3se409GZMFKZaj9jLmwRuT9sFZe6nTt7sMK2on5G7Jv8yx5CdFYw0n
UKBSboGQ/liLeUJkdVsCBJ78Br8j+mcdFbKUKBjY3ksR/nGnNCAvh+BakOBU
b5z0YDilTOHWSZd/sWA1BJ95LZxaXe97AgvzNNz5jvV9fB/KPLyqp70GMnDP
ZVCypLjCrmefZJd+zkOpIIbrGSYuiqbMCp8kkFMfWd+hcQ2euu2rN+ZM4DNU
dv04rmIOFsB9OoBxjQ101YUUabvMVQV4TJ7Z9tKH7FqTt9zkMdi+KAmwCgsE
wfl1gyLfsptFxUcBb33dL9sK2ZIgqpD/ECtr+SjrH2NI956ksb3IFd3hBGvC
DJsxUxgQNF6pMqeDG2lNBH3mqkh+iQwn3EJDjaf1F8dlqg8Z39A8OQrvqj83
mRuCCj7Kn/oD7lv6zd0dyoxEUHR1qkBQAbGF0hY3543lzkASxzNTzySJyp7u
Or8CsoMi8R2N1kFPaE78Q+3JJzQYl8VJVCQmpCF0JdNd6pQGNuFUe6YKlcm7
TtUFkz9R9PPmWtoux9dFHJdYqcz8JzAE0sJ2R7l6r5NIuN5PKVNpfUKXw/79
LZdnIRxD4YMmzdUvCkWAcZE/PA+pJNnL12TpMorAYksO25jLJqyHr8/8uo+M
xa3tJQa1QDk7uqifGLVvhL49bqhudsVX/3cR7Agszn9F1qaLqkoWPh4EeBac
9TA+5C9Jb0iKzuxmQjEtyxw1HUoskRmw3PbicGkj5sOtFE8XNZuL7pRwMcQR
rZergb593zpmBkDuyCOEQI+KsfT0iIRUxHavC1wmkdaF+Btakbn9cTGx0QXi
MJ0xYwmDBkDCGXFV2xktaNqA5NMzMcg6ivgoFQAIp014Dod/89IIN463Faum
rTaa2vr5IjhQ+CztbcR6NrrQI6gS0UxdBqI+AijOZro+QoeEfC3knhmtrE5J
1b+9CnxDQcEpcROsIJraJo5Mfv9NedpfLl9TRhMtL/4aiF4rnlls24O9P8/i
68E4fRotQVErGUT9jzxNlH8de3ubIiTJVX5kDUB2c0hyStt2Lq4VFJfUP5p0
yjLzpJ/QEFHSldHJWRXf4D/PUtgoV0PXQAK0lRWpQ4ROsTcQyeiGprB1T3/F
zfi519Z6Lm1+2Y/LopunDzsjkc8b3kTYHVmUgQ1Toj3THtmh7kIit1m2r6c2
mk4ejg7EFqWo9r4/2JyO8wGVrymYjd36Gz4C5gzT7FeK/vfO+CvCjJ3vRmSS
Osyg+hxkPWHsuvZ/+U/IoeFRtmeMw1qRt8FlFPVbxLsExk+TZVV2l55X5BjO
tzvd+yf2THcgFt7AI34lCaLDZZuk8apCq5kpu11o+WcP7TXQwkmYFobbY4/Z
njQs+Y2UKKoKlta9bNyAOH5XMwZ4E8BKxTIve8bvsxZyBMRdV4c+vlgNEQRC
B6fFgg2zKs2D+1DY5OH/zpIhbsio8DChyXliJDt8rcXqObwMV+jdcJruZPj4
WYNv33CpOgDAUa2tiu5xTQx50XWEWtjXbHi22UjJK9MyPU1hHaq5LA9O5PoI
bqhes2RB+qele71m47cEv+RcOCJBds+wp3RiitGVqXC5TgGJecYrzS0P6iTi
mno/MaZzP5XKLnflC3XN38hFgWzVWupX/lMPZ1PMeJHk3Xa4f6+WcpkqnkQW
/8H5K/WV6U2Wg5bLNcWfT1revjOYtw1QVPA5/Go88awHmM75c6waCYjBM84J
kLHT1+jfUnuW5H6ivlWadzNm19IXUO07RzYfD+V0MZUsd5XD5hDh0eWWHkVu
7E1fFdUdng6eTCwg0sgAuO/dfVeM3DVdMkhhaa9DOllEkYQt4K9Cy47ZXbGJ
sxZ5APO1FYJ1tUVDw3gSlnNvVJKw8U6DjiM2/zg8ntPmMhDi4ATZN/5Xkijm
bo0fAOGPZ8MKCFE/fGMTG3Z4Qfg8vpAeTpA3wgLy7IW7IewGbM9LRaA5WLg7
meHqevJsREjTcR4ldRI8vgtii/afzrO0qLYxN5NeaPyeCEI4X/0aQYMrADsf
yV+7CV7qgF24yYhUCePPiXWuLpdTk+Teb0XnNWDBiqKNg/v76X/WpEFyF8X5
2TzLTxDNmj8qJO3cPzOe2ln8KrwOJNlNz0wJUgbNAX/5uNlyZe3iZDrgtWwe
yHJT01mcrIN7JBO59YD+6m9FsfKnIU9ORqfhOgNxaKk12+cCqOqlfqnaG+vS
Ql7BG7U3OirfE+4KIbMDtsfdpbxNL/Z517IszmcXt1z00T/lKD4wpcZdLwP0
/v5cUfSO84ShWu9lHJ8i0hmcU4KF7+65eQkaaOU3NsoFZSazvnWVCXNdH/K0
fFaKYOt5Po0wwJ2xeDkO0AWX36hSgbJndFn3klu+kF2x+5E/TYYnnNm0p0Sa
fvFvirqtrPFoU7Ha1TIaozdCr0EmyO/z+vNlszewjgzB3nsQ6z5ARhnuX+wy
1mEwzm2USaRDiTumW41V8kouH7g5PkoTTvA6uLq/WjXxMdEY8M5uhWW7crSp
kiVf4BJrbagOcp+NocJwQo8h3ST6QPpfPcNluQbEIkW69+tt8eUbh9Ly8n/r
ICTrSkbD3RzvaP1ofahhVv5pTqcX+PvbKPycDJ9aD6rD3a13FEhRLHt+TChX
4RLhTeJSYW+daAMFxELIh/Ti2h0gz2hb1OaSw1QTFtCxgywcJqDXEFKpkas4
8nB8DfiJKu8nWoAJSMSrKtznV/TSTP4lU3ZfXASrP0lLzyWZ5DC9hHDihv98
LM5NlXwyLd//HYhZupyugyRAMSntr5DvO3Wnum4q81x0PEZyNhWu0j03f1VE
0KJgKLJhgGdj/Q7Zis2HOq49MH8vds3zvXvvtODFpsX2Bs0bgjZnwRBlD34B
1jm+K1ckZBqb+huKmY+rTDTPDUKOBGoCtumWM65pk89wiQSCMBD00RIBr1xy
PJBapIjm5hlfKZaXBlqB2ELlkW9z+67tzbuCNwWVZM9/HxV7QfWotaughAqg
EUDUat11YR/DIAbYo1F/mGX1EO1LdlsyOFnGDP9HhSPMvgAo4YbLkGMmeGQc
5UwTXX4PhlZtRuBh/W4l6EgLxwAFxLOiHCFJGLPokbNkQyRhOcnc9s47KT9M
QfyZrbBZnD0kKQe/HYZXf59+unqxaqw/7SYevVDHgp5aIhbzyJ5TUgY2eFyR
hDBAJVEbO23YgMLx6N+OomvK5gZuQuI/jq8rXcgO7GdS0XyFGVsxBVBgKU2k
1whJJLplfY+41nY4oYcKzn/LrZ9zH2m/tLC0Qb8EXCYuWtCaBC3MB8T5g9vb
6EwCIUosqcVnhG4GKPHPvRlat4OGIOFhrtTuglCdsDQth6bjOCNWqVd8VvK4
EADu+EFve8/6Z0JpiWkKPbboDe0H/n04/F6uI0jfcJ+YHVD+GTXfdLTD46iu
6xT4+Dp0i9c/vDC/uIT0IrvHpcfFL0765l7V1L96f5qwQDaaKgI/RHhmBRqM
3/XExsXQ4fvDnnYbfN516XMjPQSqQYO/55rcPEVXeo8oVQeTxwj24RpGWAbA
kvdFcK8lcpSbCTZ4oCrv/Nv52gqg16unNwZusfRzJamHHQ60GFy3S2VuuSW0
9s3/ru1/RxxMnoNvFIdxTnZVdCBwHZ/fA49u5eaVFEkSs6qHteCDEnHoi2Bw
lu7dJDd0NvWtmVNnbSzV9Na3rWTkP08Ym9Q+xzCDCZCRkbnZxmJMyJkXuRXP
hOorQ0gwIBzEcXaYCMeUWFITuxorLM87hSqF2aJIy0G0+c7aqj/9vozzYCWK
KO1q696PSTf1OiMF60WxFNFMUCJSKV8VIiKVscIgmA4wYz3J8CGuQG2BCNd5
4hI=

`pragma protect end_protected
