// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OAfSdWQVLh0oOsVeNPXHA2SKheoipyAWray9CCbRLnss7MvRGBl/ffFXSv7A
ZSw4+AkTik6OmnalSioeFYIIXOhWm4RwRA6b2Nk0NAZVw8KOdbRODXFKQLlN
VAx0u1pptclnIrud80+4Q3h19ysqheZ8o0O8jtE8ISKem0dfZymBFtOhqg+v
AfGkAZ2yeh2gsFtx/wCI5n0+i25tjJtv4NG0JXRpZ5BtA470MiaK4eIwcO1F
KMhBmpvhtXbk4s8d85OEAMQaEps+5qtAVSsbIp4grLuQ8fNxsEXiYrxki9NG
pfzbfvdg7sxmVsAKp64KST2MitWR1nPg9St0cFinVw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IZvMSCa7BWSLfVJmlhgx6c33SrPi64/6wEVuN86Hn0DqI375p6aNqdJOE9Uv
rB9wjUar6W/kKTgvTep6s3vAf13QJUu+fDP0bnrLSHqg8F8vKQbMMfWjksAL
MlCZQc2ayYE9RkRTd/U/GFWtHqwvSye08QfUVaUbOiGr8lJ1Cs4gMEAxua7Y
LWtmUBhTkTYXHz51rmuhFk8DI+VyhNsUZGVdDrIxo0o7Bx5QPpAQkLBbbcfR
g3JdysgwmJd31ctMZvvSQ4rUJ4fafCY3pb1MAQ8eVMhAZsI6aARElRhYr1cY
qI9E+8nX7VK3UZ0wwewN1TdeMDx3j8xHFnWfATX5eQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ekfhCTYd4m3I6GQFi8untcgAksRWCrwPwPgy2WfFuxX5OmfXM7GycSVRIMLJ
6hYUR5h6dD33i11VLoy76Ha67xzSb19FZatexQGxfpTGxAiDjoHQUf0el997
xqeWf4FCLBRKIv0XPsWuyVTQYBcSTw7zEXfaaOjhm+NVXLGqzl6rFFU17ftF
k/ab/BDudsm7zcEovjpWlJ3u+xGqKolaWbPdM2dow6Eq3fmsjhqo6+Cf+Hus
qihO083PtX2QokfzKW9EYMLG3oXOcmgk6VZKUxruWUeLQpOmeONfTjm1Ql5c
f78gmwWgZmylA86Keao+JuFA/O3RIU/uz3T6nnOXXQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GreQdzENvcN/InodB/LVRFZStCuyUXICfZjL+AY42YMv5/k2HL6uKiDzalBy
TeHWRXZhmsfj1Syo3DyVAkAjkFyNvnzZe4uxL1+nkKXrIKN/M33/sfFiAdy0
n857FPePcqOKu3ryVaNlQ6v6C5m8I/YGxlMN3WBkvD8o0vgw7Nw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nKSbc3Uy700xaK7m80deJDegrAQ8SmwosJgkI/i0M2cZALW2YTWsYsmim0vh
pF7zxRbfjFytxoIbMyYwb849obtZM63nhrlH9HabNkCNtr5IDpWgXQgCeM+P
hoLVdFqbF2qkx+7BUC27k9qzF9LRuXsWffPJxKD5IIxVxK4PsCPLhHINQe72
WMFcvamV4Ch1zEOS4NIB+U5w+7IA4w9hlqzgV7ge3HKW30+xI5zX1956OC9U
s+oedGd3c0TIJcnC+oXAQA26hzLQOFmvQBIANncRO27OS98K4FYcYhCTmkA0
OJeaZrhCLJ9VpSjxhyGF50HJlfLDqeCyc3C0ig2Zwyccv7nAtJsbRm1iG1Z6
7zhIbyN5BAFt0xMTjxr9JgTD4tKRvoXJKN+HpJL5ouzNs22jFtTvWkgbdD4m
veI8Yc8yzMptS5gtHbnhj25rXVnFayqeXP7jHDu7Mvj8fIetBH4ByLH723d1
cIe2szLTkopwPy2Q3JIJvpd63cpMxYbp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DCeFel4oaIV1Sjx/woYTBK74PqECqmPosiRRtbUZK5BP5mStLuxDXY2jMjwb
5CoW625SCW/pleWVx/Ogq7yQ17jnllj+xS4cU2U18k8WcidBxp1TxRPquvTj
IC6celO3TDkpacz1kfLsnTttnQrUZ6DyHQ8uA7mjvtKEFRBXPBc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NxsFT930MBDDd7Ra63HAVcfDud9P2Makfg4XnkYt1ZyxNj09Zjcs24DyF4aG
DfTxi2rnUuTUAgbNCSOJbOUSQWShXdOOw77PKTVsE+TgbJFtA8x3JycstIKd
j5vO290oFB8M+4UxWnW8wZ7xPFr+btwf2WFgSTCBI+Hbrk5F1Jg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15760)
`pragma protect data_block
7LW7PyjUn2URiGPNJ0xWrjyd4nI4C/qXI+kiv3NLqWrpZ7UTbYDa6XFbUnpY
E8uXG1nyaeaPIAN50soDScI6qh1vRg2TEsL6IbtT/XFWX2IWIEhCjp+yL3p4
hYqrPzeOg6eqHa4O/Q1ZI1qC5mfNihw2NipeixCyS9WGuUz+uVRQkFQ+SnIA
l2tcKgg+CuQVU1NYsf/tUHyATNROelqHfp7v2sDQalitaKckJ4ELIPWUuNG4
9iA7afFrfQd7ZDP6/NUzSDB6YfLtbDNRaNQiv+/dRv7S8yrQI/75Tl5P261Z
HWzzA5g0j+zeJ7LUM+e05ok/aqmiSv8LhYSRS0FH4UcXWrlPc2OnqOAYWo64
U7IAA4KSxdWTlgd/WZmdDbbh+0OVJ+bGFMkjo+fi4oJX6+AbJMOalSKX1vPp
6ivjR/Ebr1DdFmoGVttOvMzDIGZKSL46fMS1fSmgmCmrYxqDCMo7hd2dkyym
yVSBbNmj3p9vXzEz6NGsp2KlNC8RoOSr/XZLGQziVfkZuy8x6C/m+KPeQ2VC
tujg/1M/S6LR7W8EWzXGta/Luy5Z8x5mGA01dVm9OK75tUlP/1Py7jAKfbLZ
KSMUkB9es8vQ+GcHV95dBGPNPCKHbPoUz6hTWXMeeNbKTsFEAq5MdGLkdUD3
GTEKc5JuA+Kj1XC5vrnB6U8erHcoQFR6rRZY9UVVWNf0H7KRwyM+IutdHRQH
5U86PyiGicvEBKOp7EQpQbE+brTvatcKVwMt+EGpJxys90orvhaEw8AN5nwU
kUs5TqFDeofXC0w7qDmDmgU7yJuVT3khDqlvPt/2l9HveiH/Ef+x79b9sEEm
k4WcAdFAA/SifAuTEbQ9moqm+sT5PLHPvdxB7VQTTC1fyTeD2PrLKL5cCOWT
evzVE2v1LRdSkleVIju7qAA9rHjnCdPHsyuZdGXvvU1Q0EKQc9OUHbCWGnlD
5XizlImcyY+/LDxdSL4axKyNDKz6h7BA4/HUT/aRA5bIumG/K8AT3gcBnBYh
Cdq6qrqMixSKiNj6JNCbfa0pQhaOQkLEmDWFSVMH7zEiSHByhX59C93K52hI
AepwDMh0i2f4nGpQ6KQ3pMNWNkTMDfiDNFhadYTb4kqxrZvfYG8B6By0jzZt
Y8mhA6UL70yZXetS9NuPIMSFZrI6G1ggWpwhCIgKMW++g62ZuSGHtpYikm8j
LJPUvwOPOJ/2WVr/7Dft75ZpE2r8BDO9NoY+3Mt4dZvyZ86H9DPVJPfsqF0Q
LH10BNQEKdiYt/BR0ahDAZnkRRxZfI07rAra+9tfgk4N0dgYU8j2C6N/DfRR
wfminyKrnZoYWjznZBPM+jG77nwuYzGbqE7DinTTrY0dmcF3UMw4sWRz/SRI
qjWZ6h+v3GnZfpayfh8bnkzlLi2C7wX5FqDEvhGymdkl7q/QKmJl2dl5HMON
nMK8SPF4S3fnizigpvblTMwpq16yqm2zbWpMwivH87R1NkPdUjMpfiWPG5Oo
4K/Ni+ZBg5WgrxHCFpQAHrYCnMuxssvpwlgHS9+KP3/hAZ1XoCIAKMkFXzIx
X5l1SM+AnhosdLmEZ6awqBCDIlUe/5FV+wDtKNGP4Vkd7FosKgE/VRRlMpaj
d0KDI69MrYoxIVj1z8lyb4XPMMS1G4jfJ/fSBRn1vzHxIjvJj72e0niPpYYF
6Rm7zRTE9lNj4IBsZ8y+Dm1i0dqiqY9dznfBAbOnsmPoeQ+1Ofw64kQUoi99
Pr5B/lVHRY458DrSq5IhSG5ZjyRoKV+ekIWutqxM7cFurs4qER7uDBfJl2O3
9CQoORKl6nxbbKY31nY+2uiqMJouqQn/PZ+ges0kwa0OnAtNFkRNwT/Kvtji
LDVD+g1WidnMMJh9YY0A+/iXYQb6JudeQjzDefb6idIyw3mIRq1n6Yh1MRwG
KGjPG9stCCr9beK9+VVvn9kHKlFwo7lbW8vp0mBh5N0/hPgSAhmAR6/S7Z0t
Ds/hEk0CPsuFqyAGdM+spFFoKnNb303/ENrK6G0SskCiqC8pMjek8O4q6gOF
GfP2wERrPm2GK1vZ5c6Nk2y8jUcntkQ5tDn4a7p5ry/9Yp6ETwCtrokdo6mj
jcq7lLUDa1FmrjmEVD6uVlxaccNKOp1sdIfm6xY5uKUMEq1+Bvy6ktYKLMog
uw6KlPrfKCoQOyMWf3NuWdFS98eLhSJvA7UKAl2AN3Bp/ncSTsuZNQj6JXiX
N8xBMPy2+FE2DAVlAjcPQV4B1zD1APUFxUXaEsXHgaFEvGjHKr8qiVe5Bs62
cCtrV/mAsVvpwxmglueu2TRZLpD+7mLTUdMpBScLbHw2AgZszpQ73Nr3SWY2
oPMBQWGBM6RFVlgL7YvdZUfZd8uFLCLVKTO0iavUvUrEhYGcq9S0+KMJbT7G
3eHotIerAaxSkyrPcwM6kiJUPa72XCp4JV9detfY3MA8MWv+wiuGyP6hIGR8
Ze9PuAyY7HxBEkOwNsgRuycrFRDQKgJezIHW564cvpYL3peHYRTTxu/lftfB
BUTMODirGny+iI6ZLzc2UrUMpbTvYj0acUFWDR9CLjClm+nQROwFaHifjm2S
NDz84GCxiRLHgVAXLvy8TBUI3no2XHSe83Me8ZuJz6H+tLBMgfrtu6iMUUUN
CS+WJqhjmGJYMgJTLDl08aqjsud3IuiuzCfvaSokwqL3IWmfO76j7YghBSdD
by3c623F1tprziA2lTzSUkVuxgvHRbFD//gITwld5Jl0kzmXsWQskwJAdmAt
Sg1OX/lSYfnmPQfcZcojJVEKZnFX9stolD4pESnaa7z4i9VXzQwIZlTWj2Jd
WZtnykGqwXd7VnL7Fa03m/gI+NLZy2qBnqqzcvlJ4bRhnbd5zJJ8sy80FuwJ
KIgGrdXAp4xEORGKhpPZeP/SSuh7+HeF1BqKKm0ewcwe4lAwlVZhgz12uRD1
cZNZQ9qWglu/h/4fsGQr8cyQ+9vSpUaI0S8u/gwtTRBAM6S9RtWMAc5LvrYL
iAnV8DiFSwEpw1CTHQfeTvThcSqpuroF/XBuayFSzAyzqlEjpxA0EGz1QdKh
pECoDXx5jBVXQs6XBfkR7MaPy2ij9rdg9PT8hIDr3vmlcmN3JbB5xrB+nc+m
DNrdtBqOE05wZSTP5U2MVyuyYvjz2YJExEMhaCIfHWCoTyZcvDsDJXIJP6wN
3ebI/owMWr91vD8HOZGPMonfCURhg4DpMaSV2aewG/Hf1jDD0bule/7Yyrti
d5wqSk5COhe/PPa3u0RTHjbXKtv2K2jAfk2GpZuakfyL6b5TzZ9ASHrsfoAJ
RbksPLNxTiPfnK+zi6J7u3xDoLLBM2Xrf3rExbm9kImWC51KfAQvXx3XHnPE
YpD6ikSGsMSMYFeYAfhRH74dVSOkDPAgkW0psSx14WQRBCrSRcimMEyt0HHL
0jA9n7ERC1YOdU/iRw22nlBx95CSz2IpcYrnsfAlmUnyGJgMTGNRweGS0W+f
PLd6ia3AQToOniDtKCx8SHOFlkXiuok4iNVC+6K0mI+spAfS+yHx1/Hzi3pP
ZIWScNKycfOcs1KWlHlJgdkY/XUQrS1yTFGUeBjrg49meEO/gDB5aP77GhHf
jH3YWEem7qIdELol34mvePd1XFm9Gru1c317fT8YU/cPn0HyhUaXF6g0gSzf
HJCa/GjJxoeRixkia9BWx5nhTDuoGjb5eJww8NVkCG+edpPue6bvTaf1PdvJ
QjuJRa+xplKnIBAPlmAm7XDXS177coecz7riMP6mye5X1FYcRw/3OGIvnKK8
rBlETJLmjaUVl0DIe4MvpbeB+dNXfI9qujs8GZLtd9EMmDG3PlEHqpsj1Kl3
0EbgkOKegs1DFlZoBoOaF09Y/mz2yVS3rsG6A9uLX4GrawZQo+KtFVrEm3qQ
+y4AnE2g8FDPMx2J4rf/U1rS8bURJS96+IW4t9Zfd9wQqDqVierAbjrW4vvX
+e9u30CuRK1Ss0hTZH7uZqgRttPqydINfSYL/0gVN1TOhVQMrkLekwTS9RKb
2mzHdsSfpjL0n3z3MN2rolUO2HvByXMyZCJgLsp7yion5Pbd9JRJRQKdT/HB
EvroGfcuYQdUW7uMARzJonQcwd8Lh6ihvLbXf7P95KtfEgytlBB/msWIJUC2
x6khcFI2n2eIbO+pxJ0wKq8VsXQwvf2VFiPVQ82hyo+LeXpmT43fTtKyGTOI
7vOnCka2jDrSSOoIdBwyiqV6qE/oAcH4b331SVA0vStfj3mdVoPG7k48neP9
nmfUyncWqKxK+HvoCXFDbXE4prbcQuuAtHXnFr+n9T1MS5cL+KWCFJUDrbN3
+9YIbmqQR9gGU/ZxmT1nnwCFIye7OIfurWR8qC2HUphXpCHia+Jl5Tlredhg
vFhDg326kx56zq/Jcw7K7OxMuZ5unhOaJJ1ImdHDSrJqgKkQHA+tknEb77c9
fi9V4FpWltMtBsg2Y4S11FARDEPQFpVbt4rgvZzZnQmtsTAhpI28xMySLiXv
oncTlCIvr1Izb+rpuKGY/K30seDiNdHu3aADGR98bCVLSrgjOM3Z0N+DG0xd
L8X7rcMcET8mrR7L/1Q3VJ7sJemvW0ciiLxy7B5m0oTslP9KDOEgRkGCLhW5
zk0dNw1tjABk4RtpNKvjtF7TvBAX2r0QFVAQ+1LNZ0p63beXtsghD1kBDgzn
4jMFOdssV8N3QxtUmKblwSQdZB2KeJRM1XGSL9fd2ILFoWFr+xOwlPCR6ecY
bEo/LhG6mmSHHLEngNKa553uJYUob0wjmqaI4niIPA5f4T8j7GCa+fRpb9u4
ptsrkNN2BLDiaE5/dcWbH19Wp57VR2xnW8MwjIIcohz3gzn/JNOsrX85hkGg
nPc5EbKoVkJzYZwQoZY4K6NuIX9bQjMZYv141ep27WaR2MLpozGK7sYp40pV
NIWy2i3t/JGeRSyWtz1dRlW59L5nk64ruSEsNZIhNpBfD3/PO6WP3c3O87/b
a693BU7TSNWJhUlvOWA/1zykv1YJ1nAyiIKY0EwK611LFa8k4DTKsj9NH+TJ
X1J7gBibE7BSxvqLSIjv/1MvsFnNYNbS9tfRuNK/hMHiZnhG4iRwktizMZ9N
EDq5SwS3vAaOnABzJza022NDS7WjvMEkmo0Pgx9KK6SZLkbC0O3yYB8httDv
3024mliW0pfBw69KFoBp1Zn8IPEIFEzUlAIyFvuCu2c7XAQYV7VgePfgVSm0
YZ0gKzNTeUSxHL+N4YGbRp0bVyV6uVnRsCAH4m5i7uOlyJYo1G3VeWRF56VL
gvhbP3oIdikQFUQVzRDOeykYFxmKrSbREZfH0Yco/H8a8TUf9x+BRSBKUPih
eLyPt9YUg1me9ymJIbJJve4WQDjNQ1bcwd0+iT/uU+sRuN1WlRHw6XfhggVY
p+atMDkfs3blZSX82M/6lux/mXhkVOjfjhHDKqR2bWDehN/kaxhcDeK95lvm
PIHWwLRWqbe4UrQ+JG1TbUPrH4mfjNQU8B5v75UUiTXZcbR8TqBf3dajCA7U
nuOIuREb8YA/eDre5ljYkrNObs2Fia83pHVJMebZhWoPhOpfu1j7AEuMx/Lq
qAqiNaaH5/L0ouf9EwR48ohM9hn7FbHFdQVSomLN51JVlJ/DsLqDQiujifjy
pzPVK6TEZNwBhNcydUj3GGoD4aebGFS9bmW+t6oYbmVDV1o95qF5S1BNwv9p
QHN0P/1aMvQhO1pY/HT5vD7qLAw+qT+stidebyg7dgQxL3kLPuennFNWP4Kw
2WETUdvvcaPXWsRifF/Fw6F53SowvvfCgSlqX2ZyhThSuxtSnbIsJzUtf9mN
aKvPygWxlMw499n8IQhc+u/ZJIZno63LiyBCA8NJybuNIWAhZHnonR2+5EFC
u4RpRWbNjsiS7KUXsp5Gvd1jzQugTtQYK23CT1ola2gsAZqLmPIQbgTiYDWU
fpmpw59Xp0QDPSehW3eggxGXV8tsFvOSkj1dHpYOxyCUx0KNLFJL6ALaCqv9
iYqiyaw2rSDv3cE4zyrnBLHPE/ZoLWbZk5csEZF18LRESBCigqPqOh6XS1w/
Ax8NPowIHVjwSW023ijXNxwfz6HMVApWaIxI+bqk5wxKb+0/QczFlbIZANl1
nLw8COsCxxpT2dOMbo3OnYEZLQ3Q+Z92lM5s0U3OLGdZsDvA0VC5Gu/gLkjj
1y+9kSofaYpF4tsj2aqFxJCjce6+3SHTpUZN0dmNVamIfucd3DTTN7P+FXEH
e8v2chCDuCGrB4Bf0CoxeZX1IBIVpRVyFVNoyAN+I9j67u1ztVj7WncoZGWh
GVEn9nJz3NHdeC4S+SaZk+g8cgH1rAYHp9Vi4eHXR9KaB1S5xrc4uK/rVyGn
W2vTLW49TQayOqbI5wRtVzsOy9lnlqShlcS//63RtQBzkCpSh8Etb3NihFc9
ZoB02in4wEd2g2S6BRH0/fvh6qCF1R+QkgUaMfxkbtymeH8VWnhsBqP7mcqa
CaI5LOKLKW4X42/ZOymjb1NgFDhOZQmNCqhqiCvUbmaSrb939umixKoH/A1E
aPwJo5yc5Dq5Y3lSAywAff9pPoEYKxU1TqiA7wx7M8IdycF1mkk154jXUlEX
8Po/0lv3wCJXGkkvxh+/qjVUJUMTWg5Ag7Jh6ndjbDJ4d38Sv+wqQZ59lV2n
TFkbD/KBfh+DQznTVCEEiJQ8pZtkdn/DoSI3Fc3KMpiHkrFB7UXLtIYQjY/+
pKQ96BYDJIqGIwZ8OAKC5ZCwnU7EyyIovdx+VN+0eMlBtYexiS6AbBq2zDTJ
fPGl/P4dq+Ncud8M81ABV16k8hxKGojkDf8Fud2h+ai5x9cCcv4XwS8zDEHo
I7hNUMjiLbA+TJd5iyE/mFR8eshYXlvcSxyw/HXrJqS/zMxGwvFRFSDL8SqG
sSuLJ7XK/jncEYpY6g2cnPKXsUsSVS1dogbMYWNOzfITMMTa4g9pvgb/iYZh
Xm8tdWsTC8I7BS/zGDFAXm2ytUs6/+HQoJHR0bQDv4yT5nag8oRBPydn9qAr
7+4KMxLJMOorrWRQUwatEO/Pe2AG5CXIkmG6I31/hGc7DGKS/lt1HG96i13G
f3h3eB4KEMB6vJedIMwEOJ8cIDuY2lugv4fwDNjV/GRn3fhgjcJ8rLxu1Q7p
eqUo3J1NjBEjYz7T/2QSA9V+22bs1FF4Zw40M36gX312uBODEslPuon9dJjR
bHuFzjwNi9viysx+OdjRv+ZPBsIzOHRrJu3V8mlGmQ1AbzbceEWEscII1qC4
C7Nli9sexHeAtD8wOtQvbTrGLKBwDa174WNADlS/cr3uVr47fOMl185yxTfM
+W4D0QRvHtuKoeGktbxMNYd5b4aebur7refDmc573KDEiYA5K/HnAb/YxeP/
13LRAGRddr8lHqn6CI6pV5/L4IIFjUHC6sU+iCsfKxnAaPd2Crnu3vKxAxjD
zBFDB7NDJWI+V+STRhRyjzLjnUp9QkpJda91HHXnUwMAkdUoK9/Om/1ng1dH
9QsqUIwET7Z5+9lYDdo4YaIueA8KmdDwKL8qQawwEFKyZZ9bqlzh08bC5N7A
qScroNXiMYR9D1DcUJ+v+8Lq2GZdkUERBpx570ZFFRTOK3w0UQgTG1ga76i0
LbZSlrMmIqbVeyswsz9PA4tlRNHYvyCEc3qUooGTZ5TNrBQjBQ1ENM20Uz+h
2A46/sFPVZzHh647nglhXvJT7Lwc+uCWvTyFhDksOApUjAa7E3i+yNFCqBkl
715jT65lWldCV8i5E+27OfWprMmJrO2LDzp4WXzHjbRZG+gmtvKeJ7vcMxjb
tqbaANfBdLkB4mz7Z9F1V8beM1Vj5+Ak47PzUG2E7Faf/vAFbHTFGhIkmvL5
q6Hk65UEzYgUjjSzbLcU7FeG2tS5nelMsHEw1y22CHFGwl59uDh9eV/y5Ujx
JIb3pop4x9JcFifhMBMlu4zvbuF4AOPqi/qR23f0rae+1FiOto6n8yNths05
R+FsN7IyWBgC7eE9OtnChiitcXEd4hsuciVddZN3qAQ3F+UAHMDby7N0HeiI
1ejd0PodMaNoQ5xCOncVNmExzZpp1o0xvciGBi/Q+VDSMQQ3fot2Q61rXbul
P+IN1CZ6iv1uuv7d4YRFycegeKwsTqaEuEAJZ/jENgOQAYg88/ti0ystVTIO
hfBZT1vRfkSh9TsJp4J+05bE+B/PTXN6zuzfxrRuV6yPJzcQZCAach8XlzB9
z4x8HLkcUJ8xI+zhQYGnYuQdtIzaVsILqqrscCETI4if74yIPmZ7GE+0NfXQ
oofqDKSHXqYexY+aHw8DDcMCzkqP8DYDS4ZilRg/AV8pphh9e0V+TaH34/49
fwrIJ6WMO2bFkPUQ0NansJtuHJGJ0/cuvUw8Wh+FxNveV24SCdOfqVyquwK+
wAetKWmxlSyZ1XSSXGaYqV0Udv3yLHTneUFE8Z3LzHhKg4dUAJh3RyENwDOE
n+2UhNQbdfb1xnLcK/soGd1hzoh2U2mTZ9hxtj2czN5mqIrT/lcXxOeb0XA4
OXr99pY2NCNRoZUOk1xAU7Eh+BT6m4sqw1zpa//F5VK3mwym5DENcsB0509T
DzOL55OBciAPQk2ucR166BMaZIW0KQguPzA6jNjO7EK5jUMx5Wqu6E4zwJhB
2KIpCGxAbw4X53EmFeKwV6Z6M7wkLL2XHTaz2C+ZOX+nzFooiMB+X8C4rGhW
iKcFkYKDJQDvd1tJ9mZ+Rm6FvvlT02M76tyfivbZ1GN0bhi2hKgPlt3ryi6J
k2crl0kfRVAf7noeYeTKljWw5RGv2ZlEOdqB8DYVYdetk4Qx46EbEuT7FjOh
oivGJsL049Sr38RRicLnJL+qH7fA5mOWtZC+hDysLtFN1BEtim+FOXkOqk/k
WmU4E2NpczmWVQUR/ywVF/JechffsUp3in/UnRuQqeC4kL9inrCesg55yQWW
rZ22anZi7BeXcbE67+4WSHks9qgecUFNQuEpkOcr2xo+3YoH/VZo1uUbIh0f
CSRyrACUsJ5a/lG5o+5vxIpy1xbsh3yMCu4ukwk03ACWROyOkgb4fTrcdQq+
8s39E9cRAisDw350zikXiqPKCZj6RWco7GXt418mVgEGEFMNgoc6CY4r41vr
ko3iEM9M2vWwlUaBZZzYKbooNirOJtTLT+KUTzPWafyNnyxYXKL/vkr1YMZB
oOxrJ9DCLaRu39WcTmjG6ErYVb9h9DOtmuyuhoFLXq5KeXh4+/hKw/OX95ZL
SnFcbF9BTe3EB2lVKzwoiEC+b478CKdIBFnh9VBzrAAjoHELnRGiyjhRY09+
JTt2NRGSEYV0EAWMePQYup2/XDWFRwVj95S1TJg8FWNQGtzz1MMXtzo9LuKn
j3/XN5dqa6TaIT475Zkmxo24cWDJ8x901s1S56RD0y/Jb7TRx5fg3a0DinrW
XsqPuY5h5H6qZqDe0bD6skHD/5fo6SaZjdLWVm17SMG+ki+QYZsEJd8LAqsq
an/Q4enJ1Ga5SHbqocY5E1Cn+2vW5ep24p7y/9ztouLq8RlT4iPUXUV1wQyb
zXXLwVwOCBLMjz5DINgC2gKsQlVTspKmjNY7xOWm/MxAI04DudumSF0+PuqP
774ektxT0vP+9fUm2nkDDJmJuSM4N9wEFHS72yVsUIewClCXlqCLDijHyqQy
QaP2pGCxv434oBi39vP2qVul4pbGcBQ1Ps4d7BdD86A5oS5bFsdup3Akddrk
J4kAGEnxFPURuzP85yl3pGxYG5BxXZbxcz1WXL+QEtNoch8e3/2v2hVY/Mas
Ew2h3y4EZBIG96E39Vu5DsSe1hvRsM3B7nWIDvcHsIrBTJcwz/zCyxGhro+F
TvHWP30irIHwfN299BedtPA4ZdauBB4QxCKAuakP0W5REzvodhOEUfaF8/jM
TkbhmH2lA0Y3jtfffVn0Um+yAWxu/WcZW34kHHsBjGe+BY6r1IRtOcm8ArRR
c5FI15dAIe/PkOEs6sEaGYKEXrEjWatf1fGgKinXzCNq27mDudia6wD4dWTi
PgPSwYupAu+q4PADnV+2OM52jelMlHdiLUpkh0bbILrcEMDLeDTHpG3aTnlx
KdSOlNjID0R0D22rACNMwwN+sqs62lIpDHdAe6fEAeiPYL9oyvTrY4rrDEO3
5v/wsiQEGV+8dhpIRXtdxeO4d1YFI18lhsTatvufkgse0qYcNeiYP+dYDtC0
27xcg06XVLo0tVk687EleOlHHxNTWLQbeo5Dv2QdvhIkqOOS3Vt9teS3a51s
WekHlSHDLhapGLCUsE1FJej0nQSEewhSA/+dbu92htRV/DWME00atSW/DfTG
8MCZfpLmQj8fUbW7hFGZKvIsY+5bkcQgdr2xIOPcKPZuPSmVJUCJpmVrFx+1
uAnbjkX8KXzUOYk7T/a/D/Tea/jDbaeipFNQPbWoy86seZWOYj+LtQ9Eo+41
kiBUFwKpZcLqmcYoTLg7c44O06H/MHBuoMUiWIwWnDoXNa+V7G2hYyVXH5as
HmJ0eRAAahByzsPfVFTpjEhjAh0xbUyvFeX4JO8gzrcqsJiVNqWJJ6z/9YZP
vbYsJAemwZLOR894ISEpV7HMizZDFJvmJTnbatt2aFIN4VQlsGfFBbow+Yh1
5wm0CFqu4iX/ZFifzAVk5kv0L/GDFJRV7OeGx6IzhQLbFhcN7pFpYQvoHz4U
PCJf267DY5ybxBudrgclv4bVxUW122evf8YeBFUkhpaRDQKOPhZzZMTjCVKG
P4zWtotSj0zvnp3Rhr6QfQwDcl24sYbFwSm+NaJlpoO4B4h0i/PVmu8ssuy0
n9VdHqcKEp+f1SPFeHj1shJAqM2w9spymi62BAz+5ib+eNy6KGZLe+qwhUlD
j7xEPXV0INL9QgtGccZnSBlcvUpnvuJFuU87nc4DZKz0lCQW9I76kqZOVRz6
vfk2IgegetP3GM9FFKMx2oYMhMp+pIyfR7nyPTgi0PBkDo8SGSMTaDLKo+Ib
x+hGcen1Kp4oQgZmNtz5hvkhfsjech8TL+7PKkS5tHJ1jVD362DWLZrMBWHb
MadMW35gpy8ovX5RJOI/Af73pe5ruZNyChS4lSmI12LPydEgh+5zoaaMXa8r
RNyn72z7KbUmKPa4RKjGtwgs6Z3qaMxHsDdyj3eIwTF7xRQo6kCCUlKaqQpx
QTp4TaK8GSa73xdarmGev1aTlti+HulQz4md9kQxDLR//ew7RwUaN/qI7T05
7sQx2zFxzSGLvAd4niI2Y8Nohn9I7kS8Uo/A8eHhAArC+eOFFObltjxZIDbA
W1Tt+MReE62ivd0ooorwul6G4BCEv8BQtuSkAWIy5yYROYjNmnMXUMlk94zj
vwGHF2t7/Eo/dALk7fCClGqapvdbZt4OPkLX95CWKowhpJxYWAmh1CAhO3d4
oyIMuvDN2H0+WkPfmezNvcSYVYmF75E1ewfVfHGnSJv6fD9am2ZsNBCU3t6c
6ZC15iCkKyvCE6dB9a0lCNnPA0tmJstCo/F1Q2WDG3KuYjklw/Hp4Pf916My
gP3PoisFVa7kmDmLVZM8Sj49iPQOokGjgZvOpOjw26XrQUNMxfO1EddN+1oS
IyNLhLmtsyTRxAfiIQkqvmb/KgLWHvKERjgPDaXQH7cgXBHHtEDUMP/2BLAd
B4E8AL4AAxhi2J9ytzotM1d5tpt6TUABvLo+s9wX4ijJxGDmgoYni9OuWOrn
FoiaOEoxdEwzxmDPAudmhIvpKMrLJD4MTsn2gUII/I1qVDhBMpp5hoVhYOHJ
lleXt4XmEnNZDdI1s5rAL4qIZ3rtSy+J5Sch38qr1dzaY1cu9wG3S1/rwePt
BRxs5cpDrkzymRVCZ3HyuKIxgBmxHitgWcXEtWp+z0Q8G83q1qjGThtwXVQU
lApxF72Rdml6pKnYCuQzgOwnteaiuABuU1XO21gDgJ/5szCi9h9rO04Y1lCA
zE301k8bXkxmqsQhl+ahDLv9V42/LSUVwQ9YUT1MJt8mPex9yMRdIurn8uoB
ACibz0SSkxFPDsH8FWPpq9kFKGJ+vZW/+NZ4D0YdlpjTrSJv7L5TkGRbchwp
rW+kD9SBAFW3PjZwRG/4XUBijqZ3xZFb5OlKqPda3jsRRuNzvKjayCEB3rEE
Hn91fwYAPBjuCIWtBwJCr3YqxTIp2XH3+umhuO6Xc9bHxmko3UCu9lIhmScW
Zkb0xgSO2UjUbNwlsLqEXOzrhzU3qElZuIJFPlRnB41BjVdwuulQjkotJCQ1
AjapD6FKqvw8fo8BgoLSAmsrrpjAlbaic1Sa/Ov6YIVZ/X+yAYqsldxri834
rA7a6KO2RlJ9Gz6wI97SYQ4+N1+b3eUSm3kA99YWy3VSZoge1RDZgUdMoglM
2Lrao6BmczCMM0qbBG0ztgWJ8QctmDoXCfWmg9ieQKgg/0grXCRq3paXC/jF
9COhWg+fscO1V09cX9HYcOyyHpdQvNioI7DhnNB/nh0oC3rPASnzoEqirIWu
8vFx1u9JHgwSiBzhZE0/CRmAPAp/yRYQKlwSRyE1sMdum38MP7QHGpX/L7YE
I7ZMxezQiGqWiKKV45yjtyy888aZxf/N16LGSyvkejjUSQ4Pm1E9uGF2zQf3
r1Bnapjw/rJetI9/xz9cGJuqmjbMIbVYEXoKM5eElQTgqXMluoAyYRBbdw4u
+d5idWuSjNT2Uxx09QB7ElHjJHtaQNg05X5gg33FVh37ZiVG13zWp7EBk3/e
D6OwCdPebXyhQM4zyKdwgl/b+7EbxCsNgk4MKHigOSaVMVVOO7mVDr33Ysf8
wI2azXtsrJXu+TG0zIm17LcmOMZ/HVPqj1S8xvO2aKasgqtSF5Xebeftx6cx
qOCNMuIAhzFOlEY7uydGQOf5+JFviyC3q5wWiJpF1r2wFIiUX3DjlMjti7qW
VRvhPM7iPkJ33LKEI6D/d9Fw+D3XUaxiVBIxu0/iikUPsk5E01jczAHvrJpY
kHU1rlgOxPZgkYyApdHpW8eC8fT46JeC7dD2oUcAryVh90h30ucHtd+MDEDt
IBUam0kMtRS8PHwAOryB52RmFwnPCQxx0KkxDQRqmlmxd5wvdHRiaoHKoVgV
Y3fZ5f6Vrh+ynKqSN6Z4xhin9pgLPm86x+gDNKRwrCzX5pNw4tZvQOil5hN1
jvXufHd928xqAd2HAG89PHVcvvxzo7XxRKElYgC/nj6OXU/xywE9ajwIecXp
d2PwplwMlSNydanyg/5S9TLxNdxSfP/wu+uUZ5zyiRHtiDvPQ51Dt/MLl6FR
FLwdKcp5QMwOQNXJjR2D3WmODq2TyuUIrnbORsFoddFtLsWKyBL5h3GnI9xH
gNrfQ3pLugOWCKb94p30j739DGV6iI3fQ4hfn9Ds8N/aHGYUws77uwIEJb6A
xoLbUQUBHTEdQpTOSgQkRQcLRd+Ruvwdk9U3OEIYFDcrcE/FSCg5H15zS/6S
YUUFTC9hWLLiKzeVGwzGR0ExiK1I0T7EByeFeMGlLo+k/ZA0qA9+KGIMWXpu
/kkKWl6NN5Ytr0IjPDE5y+EkHkeRIYD1Wz1ZaSKFk3SwbpS36qc8LfWXCymU
wOUhoVqUmJjoqZUReP5vSDd0/nV8zV5j2SVCleZvAkKB47sD2ybhrO2wuYgg
fsCELba5H4U7V1xCzTbY/1w7wBubeRTQHNBeBZcC45A1Ok2lVGqVXkB2WiNh
Zdk0w6oEjrhKWZRy3Ozwyw2O01SXFoQpE0wCYsIY5I+/ng/QFjVZ7As7wqKn
cVHqQfwwku6znB4zZ8UoJN6cWTifqBW8oofpAaMMLw/E07MhjsV/MUeBcmmO
C9w97uKlbUCn50fVR8cWFzzeJBMPcPZVJ+QilUwZfNvIPV9DZNmAOAgg7VWB
cTDFN+KI8mmvd3wSyb0KQQXbw5YSC7QcBRYCbGBStpCp6eOrGGhqV1PiBnAI
gZEbTL9wjb5r6qJfms030O/JalXyYs9KvlKgH5QUIvkzk9F8AhFJjOq0vseX
t9KeKfuxE8jg36cE97YXzKER0HhHYdMR5Rtqdjet6Vmuo57mUGMG5e16sJLu
htt4MT4DedeEwm/lUx9KEZBb8OEnTG4agVcWaoyfCP3cDt1i+ncxvtZtDBWB
DyG822MsjwN9+dF9d9qm3191vnvPiO6DTOwJer99SZ9MORez5a2FZOk7vXeC
b/cF8FegSi+w0IgMd6D8GRJ1UUD15iS+JfIISAuGnmxUmEWV4yOeV4UJXkv4
2qt/c7gzf7Lst+6rbH0c3OCVxKdQU2Gx91TB5VYwGY9lCGgLSrvV/yM8id6j
8034vb4UE7hd48ysUo4pKiV4g2+g51SHuHKl/nnN9g6po3Fk28n52yORFdvP
9T/76+m9XkihjE9wiU6mz8+LRHo6MTilaA2h0YRsLdMAtle3o7FpYRvMzJL5
rOH8/tQRYDysk+PLaXmEBO1hiAwdj2fhUq5QiB4XPlw84RpfPgi+1ReRWUma
QFYrU+hUbjHYJ/9decFJso9zz+K5RB85QHYRYKLHxzT6kl+scLup8wUI7OQn
PA1bmxqifuK/yRo3dgwBf900RRKg9QCd4EQSFAfCPGzUw/yNeAyTvjK+iyBH
TfT5LVAWvRZz6zSInVQ1sMmqTfN+xf4WXYJCTVlVGN1GCEY+03z6KcXAVdvH
Rf0cK48rJ+VG0w1oUf/ZmRO25qKqtdBYldGNEfRjbBcro/+y7xjLuAXwLkMB
EXK3f7D0xFINRnS8j4j87nhhbCrgmgz58TQMH/FXDsfl4lvOicxIPxgGjxeE
kmB2G691ZP7FlSsBMxWA9mm9L/QPasWNU1ABNsDa6TB8xpSFMGyKTUJmpeHJ
iiu6gKJ/xfb2qdnCF1byMFHu6WCzq1tDT52P0EN0OdqoKHDgmp9r1Q/hA/C3
R4/qk37157n6R8FJzy6l2bFBC6HUMT4ZFBKeiNkPrjLpipitzB5mjL8vHWd4
YVRGYOrANDQ5XePoYINAhdq35dXxw9vB8toV427lx5pb70DUOR1zN1EBiARQ
xBGGLw78YSqhoPbl+ewZCFdQRH7VJQjwXZ7DLBvyhMnbphFTX62BSYiPAXlz
KlDYYfuDBzXLEjavEqIdYQfvXAZKmFaagwLCDj6dPjgBeT8O679NvlV7+DRF
8vemnC6vJ9amth8roL+zzzL2DrNo2/NRLML7wLVRMP2lERhovGxPxmJDkd7T
dVwkmKkWQoNEZOFdm3YW77A+bh7LvP9DKfYpF23uaa5ocw+6U45YqCzSB8pO
CApH5KDYMoY2KfxI6BcGQxPPeVTsFPg6NQ2My7jjjFxKLGwkdpFbEzrs2xah
nWso5zw3tGDcxLI5zEfMwEDIrocWlXxt21/MjO5bWiUE2b6MWB8ZXUQ+hQjI
CksYR5tbObO839tZuS9TRaoQ8WuS48XUGEDQjhUNYXcsO3F8NQEWcY3TvyYM
RiSy5m1eGp4t+obvTFaDA2ySn34f5QXWDufR5maWY3y4R1njedOnl5oIsXJ4
ZZGd6qCbeY4Nw/yGutWoYNwaV5hEoVTbsNtaaJeBB1p6CEbNb+i1LdCv4iV9
qI4JUySrc4gqC8ExAxC7OmvRJbL+34mKe8794NGJsvCqJ+tnyXe9E30Fx2+0
IrEsuKstKml86FeCMnhCp0ZmYd2z5AI2oD9bVITHynRx6UquoqFIXKF/9yAz
OuY8VhiIQT+BS8aUg3TxiZDZtnijii/cnQ80WARhzzlsk4kg+ssNdAxr+NVr
4VivZI/Z43/WJSLAVT4u1LYM+qC6ZdqS4Aau81jbnrqUns0Qlg/pGj5IOy24
FNGPs3ygpcBiZEvEFAqIGIrXzBfIlMJY5aHC4LsoP1CHHD38eHImNzCTn4tx
NTZRYyXyCUzMbWahev47Qgf32SiVPEPmfZ7CqGpGWpgAXnH2Kw4clllNtZn3
0gn1U0yDVaMPbnVbCfR7iu/Au6akQPSh5qXAHghtMANi1Z3IbTdtNxRwfoCM
yG2CpEISeVbRylhqE24jmnjgs9zvB4iwI6lFbyMwe67h2Fa9cdJFyM9OQ9Qi
1YH8RglVwO07fKhGe+d1R3K8+Jgj/Bsc60mthWwh6eILTSFc+CgTeMzXneHR
WSjeFibyt3b9yGRFCqe1mRf2yXNaK/2k4Py85RowllByn/rXRgOtt+s12ZJ/
Qy71CfCqTBGwew0p6A2L0cZZVKo7lWO+fEksG+1IeJTVda9J2n/eZ3VEgSgz
hx9oLcZII0HI09kzFMt01rNCbLfYEnjgFHof49Ct/hzj+VmQKanS2bFhF1zg
5FmD4fgw09Xk2wont/w6Y3ftrnoRpyJJlj0X3QAEiBUic+IXpMiZNfmoY4IS
q3Fd4hchgi2o9YG3Ab2xC8fvBw0zPIaJU8P/e3qzipGkBuV22WddF3Zuf4Bv
9Sk5DHYwrOvPHfBIszpE+59S9su8MOPQZqgrL+q/hM2L0PLpuW+kD3snm+Se
CaSGLOMbYxjKy2Zn1V//pU//K5zaMWsfeLMBiRlUGKkySgZ/hwW6sW65/FNx
3jquTQece2qEtroMNdDW94PaZU70MdpIhpBc2MlM7/9rEuU36jj9dzJbyt6k
vKB0d4jsxIGfxAmYbaYBgvx+3eI8Z+feNQNZQ5PTxpd8nLlSHn6thKGGUyA4
3H0rIeON+nac3t2jovIhQJWnTJEJ0BXJ+N7jsMcgvxRKbf6Qbk+2eVU7SME2
SRpsZSy3g5NX/1tmDT//gHJkSqyaDaiOMkcQkcC5zGiwwN5d6S6pKqkW7qtC
D2dgv8BaIa2XpS3jAVKdoSWAsviXp77FdVEiZMMdPfiEtYIDgZeUqbxhIoa3
7daNkJbAUcZnwhfa8aYIIoKiHATSby20e470yCthzuIenuPDu1ak4znviWTw
c7mTfj6i+NDrO1zSXIGKUabd1FEypjHkVarT89gYX5yHW5E9l3ZDqRhK8Yl6
pwOt+9E6jOkPXhoot5vqFhI7aH5kNwFlO3lKugwGXVbc7fZ2Rr0Pg4shcS9K
6U+JmOV3l2vvhSbhMGIRK2jWAsWfETsDvQB9yFtFJJjed5NDSIcHpob6gLuN
qVwGahB6Og1xDCVpMs10WOba29znG1JOS3Oce2RM0hrZ5nMTXdVdjzf0BnuL
RP/6jfXNlznQ3F2ItEm70uawDE+4+b00SSTL+SpCAEBYI7KAsoBoGtw4y8Ef
Y6UM+W3VwXiNli5zp9jIFgUqlTX49y3w7bXlXi1vkRXDe5T3GuRsxs8FO2qW
uwMq4V5H1PF/M/ldUK/vMHuwbBEokSbG0cz/UquvSkIYEeHtHDnopLhRmgBM
qI0d4Io7z/MC+NwVx0K1oT01GHuO8l5RL0xqSLGt5ptkGqu2C6oKTpY1o8hj
sYxl8rkGQf0mgOcsGJfz6yaPsO5cMYkxUbD6tujjCUc5axDIs7/T2kTY5lrT
nAH2dJmhzFGRi8Pc3eOEeIA87f80eQYB4Pfu3wbKtwhWFfvzBsz14mOwCsDK
bdi7XdKeNLS+gg65K5LRh+OnL8OYl0qNGze5RIwrVun4ZFOqlc21gv6RqD1A
CMtGxH9J7k5L7/210YEQLqV7HRp8KpNDE+yudo5dCQsT7VVJhL1iQ2nQ7UNz
Lti4UQ0Z7XqWVjPTavRn2w9vzYFVrsd5G5VvXkQfObDNyEmkYowI8zEudNI/
zi4Z3TEKjPfPM7dqpLsUNyqe7IR9rf+l8tjG9ciyi6LF74VeIy5gA6tatN+R
WGSGUE5fBBF9H2h9nV6/urhr1rpvXecXC2zG+uBUCzBh53fztmBk6ar2FdwC
ffbvni1Dh/QVJhA3tRgh6SjT48A8J6Y7h0RikbKjYqxLKudEyEYqnd2Mk265
ezI+AYQnYN8Fuiclv7xDREco9UDE0OusqtNf3vREU4SZwiwlG1AQKIRl0tHn
zIskmNL7Ms2E0W4XkimtZK+10j1uebw9v6yregim0mBI9QACYfuTg+uPKPh5
8DmVy6hP7BVekDH1jve9uZO8cPASZeMidrN6JxdoBp+secIQppO2hRb93hNu
RhZi0I7ygHG7n2i6NRC58c6EE5kQGh1qBXpeEAmAem9HqmUtmIjO2ebNBw8b
NGLrSTozNIr7MxrAZFvESNQInY2OzCIeSkCxvY2wOye8S3DXmSPpHhvxn/pK
KvQMbPgKcWaGG98NVlh31COIUoknyzr36X3lGcYamfE7zK5du1Tw+E/48y5v
x770jTIdqmrCJC2K3l6eAxu7m/GFDAGF+kTtusA6Agpo16p+JRelFVbN1+vY
50VZ383NzV47eVsZycDVunsZbqWZba7CjQ7hYVqkYnS5ZFyMyQJenxUo1FcX
e0NHgmDvbeFv6NFgFxthxcESS+qhsQUuPe+Z6PVin2FkpFZKDnVEOVy9V78R
N6iNeIfHzTHDX2v3schr6uJ543/3p2nQ0/cNmOT4v3lIZ5Fb9r0bhBj88tCb
kr8V/HoO/INM2GJZU15qkoDlwWmhacS/Ci5Zc4j141UAq+E+J7T7bpHFV/am
/9z1nG8hin0PFKO0mJHeKxsBBVHrwjxD6/UjutDvLuoyGQSbSuYWqk05/pBr
43GadOSqqUnaWT/YYNOCuOEvN564uD2rqhH+ZaOP+Q7QLIctriPe70fAMh0u
xT1ScuyYF0vGOX+BrnU5RgojMqrPF1h3KlpqT2Miok4lZr2E8OwDg/PQv3je
5j58wz/3td5xpvdU+wQ9kBMFrm5SFm8idVduQCLsJDmBClc6MD7n8CMCuYNE
01iDpEXyMerOril/7TP/DuBLJy4o4IfjpgPFzZeYoq1/pzKY0iGELR/W3nBe
WOqTzlqqWBaFr5bsLNW9fKUmpaSV48jV9PomtEnwf4P5xNWkTOqjhtxvW57Z
Sc1MOUaz37BtylJSN8QaMfUzTilsKJC5N9TfmP5JjllsuJW2FoDPv2DWSOJB
hFTD3d+vFkNyqbwD6zyWP+clceJb2vFmhADGUApY0+CRvb+4o4SDNghVT8Wt
Uy/9mE7eqry4J0NTWu8q3IAywYR1an2dlVAixGy5vVaiRkbS64X57fc5ejbX
/EGeI8jF3r0NwG3Q0szejNlqlpWBb9e+smMp3iPvT60f9j3kWZNSSSLm7ofX
YPzCt61GURPvDH6aICAD0+rXTn/MlaMVEh2qcoTuNPOBfcdDgqakPyNEqqdy
Yp6odSTzpuMY26kn25JYPnWvxf0OWj16DM5+NqL4taJJoZBsd5tceQzAERwY
xzwR1J5TRB+0IdY7UqiBmxVPPEim+4o9nj+be4Wsg/0wU7gsOXaHjL8LcIhi
cctN0gk8nHg78oMi8EcS7b3meC9C9B4BM8OAYqqdW1Dtj/BjuKD7luP+/vl1
u8wAFBY9D/xQInRb9Gt2iP64A4ik2gPY4qOb3IaFZ/YJ/Nk9MAdbxzsCJm32
UtDxipao8nGyhJeXSvTyj8L6I0y3r71qHf2WZcAg4dOG/9lpDw8aHy0PL5JM
gtZdOMYx9KigD10EBNr8XZAeisr+A+79WRK7C/D7p1VK7Rxcwf6Dirdqqi40
I4QlA0jd2Q2edw9JqRFrB9MOXXOOpyJsC+ju1Bv0PzpkQm/uZQ2WEjjPkLZN
wE9uk1RVUGU7QxCFH2bo2vfMoFopFb3EJ8jQsF6+768I5HguyTwUGo2dLTJW
F8LU4zVIOwm8cD1vdkNiPsNFqg0GfOQA5PMp/p6H45hFyHfhXfIr4qCuOkvH
YI67r109itCQl1wCEiBsNKIeUjjbZRkpk71aHbLAcLNjQm9GWTjAKZI+peGU
2Wwr0Fh/339AqkHJDLCdy+dBFcdXWrrx+kW2mG9LPNQUQYn5xunnpNryKTxB
dL1akkKRexfwl+EzhYzE6Qj9FDur2KR8zYBchWHdy8MMPs8oBqUcZngigpFz
mJbmDJctvHr18eZc2NQ2MeXD5N7otoWdkh6n7gDWCARW2Lwe8XN+VHYVGM5f
3WGeIL9AFJ58S3hgIAjy3h7tgkGGN4a0UODdHfn54ZwIHJErfFP5IzFUr+UF
bUGtvoZME4HTB271LeywEbL7BrnvQzAvjRJuM+/PkA9oTqf/axE0zXLitoVC
eGxSWK8Uw5I6RTsKvq6SE58KLi90/RIXAEsFpFAouzZnLLwQv6t1lI8qzLZ8
ECV5rnKpC6fT+c89ZwgUXWPzVTrOlQk8F2dqPOdVIhrDsHp/A0aLycxcbwrk
mGJqQQ4YzIW+1wragBaJXWHaxwVxhCU4RVUR8swRwTpfIvNO/wKAcZEqkkpZ
/DP15UcVIYv17pnQoO+RhiNOtN1XXa+oTaKaXC61VqRm5zwgWviqbAGqgVWa
OhdsD3pLL8pcQ3r/+DCaovV1gp1k8HDnDA7G95FF/wmnfXtgUknmVxgdaKzY
9QXF464qG8iPbEOmwMP9O39w2p/B28ElxjF61abLU7/D4TjPKyl6kdRiIwRZ
7bj3ipA7pQFVbX/PPthWqc3tJlzP2UqySfBSSVV3zozIUN1ZDKCxInCadqhw
0ygrAGyAkoWEoeRb5+exlGiEhj9nUuxQ+VFn4xjF6tL0X6SBSLlaO4lbHysz
Dcw+AK97BexI+O2mTj+7h69DTpZbLosxuMZ5Sr5epUNNBWiB91my4d258F74
YaluvkZTcWr5x1W+E8NW9M5z9vy9G2bsmFwEwCCbWIKmvalPERL5+k7pRYlr
MrlD56ApGliHgC6F+qGaqCxjh0WMc3ZqahttX6M7iJyQg8rfDRILDU7tDxnT
sZ/yQF28tdcHoQjUTv/UsjGU8ligKVuTFwT+CHDytywXQwFeNmR0ZfmJTpfu
vfcSO9IAVyHYBgzFuBbKA/AiJqF25sKhJ/Zq+2AqhtrjAtm4MXqJx9N4hdaq
d8EnvrkZYpQi8cwjoOrGi6bUS58UvsfVFKAlW2ppfbDAdYr+cdPxVGlZopQX
4Wz+zcqOZaMnaJep9r7hcLUapCOChXPzyzXnkJSDRfweqBGHByl9afqr0aXW
+r30dNH1O+g3yS5dUd/cz2PUu9SDC+3Q5gRlYiOPEQ4j6Ylk8hKz3EdwtkgR
X4DjmXxhQQiv8Q==

`pragma protect end_protected
