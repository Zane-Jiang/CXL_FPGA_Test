`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
VIh9v08U2DoWiK42hQVP/6zCllBiBsBfWu3M3IBIdAH2A24CvpHSnE3kR1hIsgNt
s72ASLCWGGehCgejcAsykzu9RmNEwPKdz9HUhxjQ7rk9U8LSF236VLHVtLCfWxR0
l6gzB1I0UZo2snBLyOxOWGwJ00B5d5BbLWmWM7oBKmY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
cXqC7ExQ4kVQtjGrM51j1gxmJL1ah/Xerz8wOrXO/+hKuhrN828DRHlWkq67ce9v
FHTsRerspYb5V/bqUtIjoe0xgB1U13+VpqkRaAtM7f9w21Dnxyk6sHTUlJ5YAcWm
CimGZopjhJZ9Rbv8aXae/SWcHhQyRNetXbskWZWREpYobom81boj7MEu0bOnP4t3
oUuqWWHZtao0jMLVMMU97cR7jff9HquUxlmSA7QdZMUUQCz/tgWZ4kFr+L0l31Dp
h5hIJFDyp3kx+9qF0C08VbZ4ZChCbC9r/r/moiHsHFiDPOWGFKB3XbMD8wYd6lpD
zfialYozS5yHr0/hxOpQCfNI0Pt9FM00kAZVg6g5nKHItsK+NNA6AvzFxYvTqke4
dxwrNu3+sld08hm2ZhtDkOhjm1Oog7T10fz4OVtql0XOaU2hm1nWFz2Pz32/S3DZ
XbWYCCmOpJ2Ff6W2hYNJW4K6sgBEGLeqL2kcVS4phojpohjJ4IMT3M+c7IZNQoI8
6vS+pXYrVG0eKMdL0ekBat9/M/66qhZtg4CJicBQ5rxedduiLGhdN5/VE6jCmSda
r+URAVBPX6Gs1LlKYd67n3cNMujqpsBDbQdhecKK5/A/rulYgGTvTV3vSu1wJEJJ
2ihU4eWIR4olZnCez/dYJUoK0MWYcMUJAgBafBWycJ5g4d1YuH+jZiShT6PtKoLp
fMnnyB7n1tifsinkgyE7nK3BKn5y3Ko+HCr7RDAe4kY2T70tcAG0LG0uzleamWpk
2jyaJDD5mF+Y/nRe2OJ87tL4+dLhSZ8JGzQRiIbureg//C5XvY+LhtV199VCOpn8
t0n6qoWmbDi9rjUN4FAu6f9ceT2dmTVKXiJjjgKz6wI4srNwugd9pr5JSiDR09xf
w4EVo2gqee7lq5kPSZnL7Skbb1eMAbKUYALBV4CsDg497tw/hA0t/vQs6M/3nING
u73zg+Pu+Rxsa6XrEcS+VS1JK8um7ypUl+rIIX5ghKIJzpKTivivAOMohASY5EBD
duy+CfXuN+N41w5ZPAa7Hy93QmhaT0Ie789VYaY7ZFkGNGE+6zWwsasy9pgHvGZ8
xnP9GPnbJaG+JPo8XDot3+Bkp9MAd2ZtP3W1snR6bQz6Ci4LnSndkGRdPLpwypZK
HUunOhnWWafp3IHhnr2XEFrPa/XyN5NkdXkKsonMpvt9yU8Z+ZzY08jrZMYx9QzN
/g557ZvmeMYcXSbdRyW0L4rU+7O53sAhMUw7PmezRD/wDxz6FOLFqz1wwefZCnNW
5x5Ymn06DyZGBVS0PPO3nrRABqqQoUXMUzPJZY1tPJlI1nIbXLDTKOVOtfDvHQ9Q
sH0MZeH7h7FPFO94OKvlX9b6iEFe/sIY/zEfnHBrXWuWv8+rtubrkwzWucqg5ns0
p6KOgi3GH8Hbt0lYDBrWammcS4oLo5nq6xRTMFkj8/AW48yHlJgEB5LOc6rHxPwW
Qytiu2Np8b7Ps+9JnA8LKAPzilauukPzbCSBaR+deQqqLa8TXUq8tXM2QggTBOme
XNUhiola24FhQwdtPBiYe9HEXSfxeIZYtobT+VhVlPvGk+K5lBhefZ4gHMzKOqCU
RHTpWzl+wmaBpzukU0jjHOovRnUuH74tM+3dZGwspnoylrrNET1nndg7qoRf+MfL
veuSTe15Ca/t8O3fCAAO5V2om8QIItraUNDIdOZd62Af6P1gEBhaFwJzCbjEiXGD
/rq5CvF8Tr1YBWdcxY40+59f0td5WvUmyhisOxe9+3sDNHqs7tktVwCGHIHJBHsH
F7pDDKWxrj9iz3M8MwWbeHHZJakp4nZhAAbSGLLdZlZ+LSjKyhtcBTUpvPwHzSUn
XDO8xtIF3wZd/nQDHDhVWjoCaT0iAop82bOpTEtLtPoQtKdSH5qWu666X/fGHWZb
wPXBY+cPXoVfs1k10p/n6chMQvlj4W2zeX3/LwOQ3cUkPkIrB03kSNY264bywdrp
LBsAwwN2Ez4a43WWY1BYpFDqQRdwUswO5fVvC05JpXmYRjPS7q4Q6EgAhSHyozoN
LQL0yUpIZUhWkwjPQDvSvgy45RQjC8+jaUbj5IEiS90jXJKOfQNaax+ezJ3KY0tg
6wfPtFYDww5XCItauXhgcgAVx29FTYQCkrhFzz3JolpJ9wxfyqBSZgqCCvzD9231
RvOcsQ7fLqt0yi+WDwL0BLT5i6illSwnAWTG28SSrf6fyGGuafDcUR+FM2ahRU2O
1xtrNfVW4rGWNQ9E5+Xb5VLXykoOG9zSnx0CzjXOCAkj/bkpUo1uFuq5DY0Gu83q
d80ELN0HZZIlilOeJZoVe5ETK0uL/eKwKjlvOnmTm5mj/cWRPPmLB+rRt4atCro8
Vr6lSYmOkiA8Yxfs2M7iir6e34qQUyRvQw48fMLllmEFyB6WN6fFlX3I3J/LeA+3
JdFvMEeYo2z8dN2P/QXvCR2PouS2v68/xwmAAou9h64Rhlr28iKr3arCqwtyaL9s
StwzwwjMlnUgAKNUIgKeQ99hoNmgwzr0VpPsX7WWGS4kKrgJjbZNZ9FfZhFCXYCR
0wz+CTbzLWMC8yg1OSx8djrJHDY3nC89R01Cnm2hsUd5mwvofjAm1Mle9XDe0TFE
yvE1A1fjzQ9cmsBDrDZhzDC0A9AIWPLUEZIrNmwcol9P65bywJxyPy4ZKBvnSFfs
KI9U+5URUkCeuDFktP+BzcGa7kjb644Xacc8Dod9DCOmHEZSLsKnM2wPgyw/UrPx
a20n4HJgIEOTjSkJu+sqkL2p46g5ziGjVKkeNRD68UslBlGUz5HQ9W0H0is50xWa
982WHM0Qp956dpHsDq6naXOkz9SRotQqPbYbd9MmZLG+ytiSzBkbX1OmIUEyKZs7
oh1Nyn17TzlRtOcIQtI/SJIEO3CHQgPcG5BfRAAbM/DYsg0Gmj8V5J7noTwX8UmC
u8qYEzAnqx3mQTUCUJrwF3jRo0qmm1t+2mhp84+yny8WrYCOCFYBY5ml+5WkQpUa
mNXio28m72T2ej60HvOk/p2oZSNxH2ySOgZh/xL1gTEp/JPWps2ebrSQAZ2ogZ0X
gqVYEcspbqsHihmaCdHIrD5N9PzNppQ1n+8fKRaDpv/hY432ka/GvtW7CQC9cLbM
ho3wgaNA6QXbkSSC6Ej+xCKMKQTkUNn1TtqXelSWVmgGT/hECv8qCZisHz+7bNe1
Q8i3w1IFNvMsnnJySgAwP97ZgvqQiMMhW/Gk+QuFuYzwJ+nLNo5Kj4AAWA4AFAVz
bzWUj09WtJqWOvw1F+SRa1vN10PE4mcixGAJoWM1GpGrcVCAf1NAxchdRjxS+jbW
ubjyEJdwtp3zXZkIEkW4iKz3fRKwi2zH4DdHU9fcl0Th4HGA8E43aCszmvp3jwZv
Mx83EnR1SvK2yQ9ExtbZ4j0DPWfCR8Ekx/8Fa/n3ywA3i4Spjk2/rekVRG6dE3dA
rRt7OuV7T7xP6Y9PZMCVisw7trOblH5Sft/9phHIGM5PNV31MN+ZXtIA0Jln2926
Jp+P8Cn7pDYC9F5/epHSWZz7MpkqLVEwXx7x/mOSPS8BrJC+Kd8RZtEIZDuq4am+
r9UTFVpJAC2mskqYisYjuw0Sf9ophdXNpIvImbSMWuy2YJ57qp1qbA+nI4++fxz+
ljtnnZOx2cvLsyfY6f9OfOqBBK+vAyufStcNFQN37smY6qvlKU4/M277153PGBDA
PTd20gzgrcAY2qtlQo9y+wnfB/R+x6j/XBfbCiXaYpO9EiEfY3lj4V8a8FextcBM
KjXpTVdDL1m+gjQqlRV+4k1W+mYGMybXzji6sd/NYIAXPcsbmpnUa/+VI9gjqUn0
ZZj0yEa4D/2niVQiFojvKkqCGjbAexGL/1Iiuqqw+NnQNGoW/OD8YL6ANlVs4vtF
c1Yubf6yMtVlTgjbi27Y77B2enpp3JWrGSKpZdRRkPGxeqjS3uDuEBozUDTXelAA
vGjVgaiB0Wq/5TSSjFL535pjZsbdj72rnDZtWFntGeg/EGBMEqq+K+uQNRRcj9te
Tx0S18LHjUz0uORzs/uboGjUCAgYZZl4AKI7/MUeAd2sxcieehTK3i47wru1+NGi
qnclhGyWtPbu3NosAAt0eFGDvatlF0l0TLDJ8qEuS5QjrenKlpwdvO0k46KzpCC4
ti7qk6ZVF5KTypIkEr/fWcDTDZON1gRZInPrIOnnwdOWpuGf+s5cvK72qyH7JWF4
zywsQFo7CgwJ/9K7xb7Kzs1p1UHNUEIJbJ9IkXavFSJKd7B0pnaKhMpVMoxJwR7l
v+BWWRBU3T/rfy0fTe0wm9OAlb08+t3JYqP9EdCvcvQJ9kDy03awALrbp61UgrIS
vDmANs7j+Vfiz85HYy3jHcUo9YSPcj1/i9pKGaqrUlQr1NAo9UxKpSoBhkDRdixN
n8m71/5Y/m2qWmf+jLJmMrjN0g6llkHEcfMjYkrzmo/MRkKInCbN6fpSOfcrOMsa
K/SYrwiupYAmNm896eQ8aS7nL2X0oV3He9ZLY8XcGawfQh1F7+oWKiptdmoWha/s
zLDsGr/uXng8OCHbeR0D++R/5rsexWLkkj1G84zMGR52w9CRZSEelf8fHLGCwBh2
G0zTlg2epuGkgAAyGcyCfDABQKZrJuz8l1JsVs/ktaTE+64m4VqYE7fX93Iuw5ul
J/5IBWWkDSrmzzREwJpK0VrTTNJaRLRMUdTjxZZujG8oxsJARoHCrWfz5/jN1ezv
I6qYyuIMi/aaDdtQNqJVxjse13ZboM+rSf3qh8TyHm+s5yEqVfG/chC45VSAesBH
uVuHSB6HzSn2efgy9QIPWB+1B3iGDmM+UIN6yAHVx6bQgazzwCI/Hc0C+Mn3XeEc
WBG4kSmkNRjP/kfEzjByA+rYXa0G+I+2x1TUIlVAuBXbs7mKF8lBQiixHx54pDQP
eaEgAmlf04FVji1v4lbrix6IhxDxrIWz6OB/pBUxGZ1Wov+NL4KNAZKGqBJ5h9Bw
/z1ynImoSKS61fMMxJnh5i3ez1h/J8CimkCGtCxKjwCJYZToc3jSDXIFB6KjGVzE
fMXqLqMA4vfzF8F+RLKrGlT6VeCdoIC92UmJFI6kh9BhNfwkCe2K+gczEgnXQsun
M+M8MKQxzKiLAR8YhfbpjAdhG63OthFj5dOi8rb15jAykPmGPhZTZgYSwScnOwbk
n+7OhzOl/c45XeRrwqYYpPDU3+5ctlfaFd2tNI9/HavqJTzi4bUxIax8EC4hp64F
VqovR+aNfHGcSC1LgjaOBp5pJT5GU/yDnkwMSfC9Hp8tSA+QoBzdjd+7F1ztLetd
XtKscFFAowy7BTeP9lu/Ii9d5ogG/uOY6/GMhH0geX5CSyqdthaUFt1wdyfofroP
gIQkdSUL+xiADJ5ZUGSGwOYCrhfr69KNDHxQMsfmlZyoRyUd2fB9ocy9qoARKTt/
+34oedHcVDmB9X/6h+UlSAS23cRtUtnmiKLWtzwti3J2foGlZKHU91yVex2w9Oq0
RNzO0FSTxH/kKWXVI40FLyDGxCfidyh3oKoHf4y2H9K4KmhB/AKX1rwHZUdvwZ1G
BhlSQ/++OxQB+WP6Tf7uN4fHa0VNyx0dfHuVg08B9ScBzHAd+WIEXUf0+Zp1aO51
Uek7zedz8eFRr+qM15sBrO3uveOCyD1cmuMnNQcedhgcBX5ZFhkovLefqQScPj+5
kigsUu84edkTjknNfk/zzCzum6BB+G/UFWild8Cd9zC0Gc/1WNGAZsmar/UJLsKc
LUP4GOE/U9rD/6h1aFyCZj+cFddJU98CkBzTW4kW7VlZyI0RsncaTglo1xh86aC6
UG/YgqSrMFqJxo3Hhnn/lAl7bzWDfHu9m7go29pp2oeFyKJCuKTP8GqUrxj1K5Af
8kNW6nBU2TLdlVnGCBSdune/mW7bNzg4IrMcd5VWX61E9j4jHDqc7/fMmBUnlOPy
mKb+lgkL9kl2+4S9VZkYboXuB2oRYDtaCiZBWokRZ1mo4fYpQtkjBsdZfZ9t9dYU
b9fEY4m+gbRDakCG3sNN/8V7EasByQW2fzqYg4+zk9wvBEwCr4vktxUz411YwIr2
P16M5JQ+gGxQceD9we7HHEN0U0ejJTzDVCftXLyTq475i07ezD8g1uqdnR9GgpAP
8Ac68rDJqoQfCNeI3Ln9SZ/sca1JCcxE6UBof0dAeeGQvtd3AK76nfH1SsuNv4c4
rHIlVU0Sdxwq2rvEpexUw2dx1EiXDwz+rXjV6uu79+8cUtMOpl003oiSF0qLqA12
FqM2IPOut9Ww/bzd0+OQnJMHNxgkoOEf/kp2BHLnsj1rNoIKM7yGulqbdAntpJ4R
5YMuiF4YKEtY4vxaTo/wqE7h5JjrlKyn3TPg5BQRW+Nj7IkGLTvu80k1ZiM5Vp1o
XKawtO7YNoXky/4SoUe2Q56W4ZC7nYD1lx32NBZ7iWAIAlfFCKH081WiTb3wFPRy
d81+DE47j/0QuLIYwCNaVV/pDV7OrxN7nyzoaWjzxO8HISuVFBgq9GSfZ4kxKhC3
KRiEPVT/ELAnwaLGJdMk/vhgJVTNXz7h/sQ3GpMeU10DLkjma1ffT7Gpo1+RTKl2
Vqp7PhM9Tj6clqR39tL9QIaQ/WAHUdkoTQhze/CiFhSPLB/gZD+cjDb/Q+7TQvLu
jHUFY3Uxz/rU4qe+AJyGjp+iEpDMbJJkUNBIJz9ROHvTgz47oPP2atRjorLTg3Tu
AOWi+++mJTCFPtIcGRdsd7EEuBSJ9l1OCiak2BXZynCpx8Hk7w+uzE2wzunbcbEC
fniQq9OcV3qOE1snOnlnI/wvXoTYCdTGKTsw1qeX6fHCYJyNfvZfxBU1IjPcONqo
G5zhkG8DIRFPsoo2PanxVdENmUs//hJa7sBxxBBBAetJU/SRngbfySjttKPWx+08
Tqar8NzaR/cd+YHXn5uhZvpGTW5RidBeJwmtSLhXK03pVhUwWPJL/Aqx8fzeUnK/
beRYvi5sua1efuGCDailwjKUDO2hTzS/ctTZpov3kXHImNS6o3KfqDE90hinelqI
4+cvJQZ7uF+T/Ygb6gzZT337HbEBGnithVVQk+qyk9MPVsCQYNuEeScqVWwljZLf
8XeoukSS1Id1BlcjPT026XNfaFhVX/aO8IGuAFtcZNE+pU5lufkJorYe0Ul/SXnx
9kLFODn66IIQxr5zbw9niQmaykRSES3/wnCZZtCW3Z4wXfHC7FEvyKF5+RSHmWtt
oycOxrokAqpsi+aKJxBzCJCO0vYznR4nJINeVc/s5oXW7IKurJXjREll5OsirffP
8YrTi4LOR7ppB56usB/tirqr01ZVrjd4ywE7/w394PTC65TakiJbWaf6KZMpAbcx
OG9JuLDgYgfN7CMn3k9lstMrPTFR+6zwqdYV+YvhabrgnaGBWxcgfIDVwbgJgAVR
19BRpQsNQLSLh4CGmqflqzrncEHf9j2x36e6I6fbbJ9x+EO89Bs+CTUWAd27TXx4
YpcnDopPYzGV2zxSTwEnOug+MvkXG+3PDW8788ilthG8spkVNiBecsO7YLD73ewZ
gV9oXMsnyvc3ioMcVIBuRX7UKB4IaqaENX8QRKZhcpfmikGlz/wOC0IMkP3Fw95x
knExqQLSeCQq+AqZM4nNIA75Nqkae4W9VdseJRBpZ0z3MCUC5EgOeCZgYln4RK8h
FT9ehIyfgXhAsy5rRvFKPCmLtutBpfqvY/ddaLitMAreiwWmHDUw/lt0RBn0V5Cq
QqOL1gxwE+fWP/GDn/LXtCxKTL9LzX/2F9Ouhp9zV4UA+KGuo9eVF5yvmUP/3yrY
9N8Ip0VqpOyoQXThrfwdgICsMDAYtUw/UJG0IDfvaIgj58iYzydsLvSwYL96dpxB
8PsciICdS4Tn3s+FCFO5rYvCQqLqcMgY0Mv3JotJFC4VfU0pJMq2SBgd1cGLzQHt
JCVN8D4UARvPH5QhHYA+z5YIMfaZgCcX7FPPVvLSJmG1nzXuHcrnRiKiW/CWxxZz
Av0nny6maRSPqDCBEWWsr3MFnR9V3m7M0GYTJRx5H4xNfyHQm7mGKmFPwJmiXSUZ
+FQqLrVAAd+l0iqIa/0oTuCgXmCtK0x4mYw2bqveZagEnUvcCbvE3VSbXH5Bulm0
cGB7uKWB5SRvcrJ4RBlZyUUiIgCjMfBwBWrJaECTs8N9EhNelFkfRQObPvHfBJJg
6SRxDaaFMxwvA2RP4nwNmje28r56Mm30e1ChV1sWRcyq5A5LEFny1tbrdOaShozH
+As56WfrMJProtzgWTP6yeZWRQBAHU8Y5Kxdy5ygeasTn1cf5lt+gOqflVmtPpyF
7Uhequ93C+sN2QH9h/cvf3pYEw74BdCih6sZQgpesCmVFd3w/+zLaNdGjOKwEg1Y
nfPxe2QyV1Vg0a73Mf4aGaXHeG9KGSqYxqOTLc9HLhn5Q8Rj/qi7dtcZEozx8JMy
zIEz+nANESq9pofle6/cRG2rH37wWHMChdz52u/GLd6fmoIWc0kNH1ZkbM1utunI
GrUstG8jS6U8L+SlUKv64DBTmQgcESQE9EeUF8fX4E8txzKie4+gQZGXCt4j5MT7
4dXVLKhp/G3zGPCY7qFdy2lPz5dVTd35DJyAt1d3pvQeZMuRI8QxYeD+YcyRW8vA
bC5VCJmXoCOhwd95wMiItjdXxdHleeS/8IzOCPlkR1YMcpjHHI145pcbkE0FEWMw
6U1aQ4UJd8cuI0JtHVhRkmixioWqm+L4xGLQzVX9dS8jdIh2aogOqqmJoE8ZLfdP
HupLWWQneuA5sZ8eM6s5so33bA5p9Xnf0g/6NIJ4KFQad63C7em+F+5LjzaprYvc
w+cM51IEvG4mZtmvS9it7LBNUAZpL1F4H4fBvAgtXBE/Y9xq+nrAen5IJF0JifBa
dCHFSk3DlZeOIEBQk31NizqSh+0Z5a9QuldDllWWRXvbaaKqvZQlePzTBuchK47I
FxMkNZQpL88TLNBhMt6aFPXVv9Iks2KToL+QB4wzrwAdlkZeKXz9FkteJxq06dTD
/VONlkDpAU0gsn8CE0RiH1nP4d6KSdRAN5poTSGssYeCIYP0i8oOwfm/L9GO6C7G
05xxDLwkT6V5CeMIKlGLeTeWnFXGoRgamE+HcEEcdBC4r9uL3XlnuqcxXI839Ues
zlIuYihwX4h5KOYITJAUUbZk53+TqavY9xJz+4AIf3Vb+FtTQRoOdW+687+i/BX1
wviaJjSexIV/8S/43bAUVBS8LI0MFT31SoOohKAxTOuZR5SN6ksrPb3eQtukmcZ2
BYNRIAGrSpweLopymQVIoUAVbxHtpta+rD7lEc9tGh1HPLIfyb/RAVnrqvTiimj7
yp61s+VgSOwTxtsIpK3yyVhuD3fMc2asYPj2DjDymnW6HXAY7SPeoK4jxW73PWFJ
/MERjGdjBAGtFrm3flO11JGx6nSqbfd0iNgt2xCRLmkBx3NpoJzpNjiDd1jByfTW
B0EbsaHVZkLSyZuV0YVh8NndxqRAr/fT9MWmIbTNd2ofpfG3y1thr/7+vtenFfMu
nr8hoPByQjdH5vBG6QFD0tr1LcMubzWR6kFhXn45KbZN837o9vf8YwIVslsORKE6
tbIhYrtQJhuRAIlevCD/kj7Xcuz1aVvEcES+XnVLejvE1NzavOUGdilX0pfUgfxi
4UbcXI2x+B5ISYd0d8Bo9eOkVlUzOS3ORTTE5ZNJPQjx4l1d+ncB3kt+65grbgMw
VGoIc1SmdhAdwomh4eOErZrv/jyjZhhWYEfNVP8HpJDHcSqIsKk1y8hcrp13pbsY
iOYqwRtrcMrzyHQBmyQ4yXyiO4ZQc0PquWj8hC96U0AUhDgj0UYJMWVFY4k7Cq+U
yVh1CUlzrhFLxI9Y2jkShQXtfPcS3hzliaCLRjL8UbbYJApx9C2z+LsK6ls24sv7
wjN8SqfvL9PtPS/JN1etd06pu6TlSm0WyDLcYO+5w+vvaGc5M/Cs1mqXvts3YpcV
ry41Wyafrwc+QSv4aU+J6C+rcKycYvyXmzKG0Q30hsU+zAjk42gEa99abdhfrxxc
NAOymITOeBEq9OpgWFe0zCikuzfEzM5JeOwHJx9v9KO9GWyXhnK4riY3ovkTsxIz
lc7z0Nc+NA5+9O9WVBT1W2/P16IGxGwOawJRu1iJDIL1gRkI9mhid/zAXQPmwH6M
2KGH/yh+WYME218cRb+xFYvcdNFHPK0uC77zIrgFLtA8A/VqD5PpXn6cyp4DnfT5
X8N2+57lDI+Lfyfai9PNeYDFgwFcLU/HxewvVzPqXcFeQuWFQfA8PhM9RrIVeTyf
05CxZw+ofMLaFZKg5UHcfwX1OcPkOgTLI7BY/lYpXYwDNY0hFFdGXUYC/o+yWpnx
YitkmEb1BCFEjVUsAKClc/etwPXhbJ7uN0DHM3A9daHuBQB3HnDF2xybRshO1Wfs
YqwnefTb2mj+WGSppEkgog3maUCsmIyTzW8Bw0mcTybyK4ll91u8OXtt7oownZ1v
6FDOF3CCrD4bo9mpTrUQ13CLNnIPxKw2qnL6FsPI3Dr8mAzB8qEMZKZ3PS69QVy2
jo0l/fGHkvTs4E4zQ5JwSHpSSX+hwD1MCHJf8nN8NWVp8oI773MADwob7gT3UcP5
lLbhnWyjjsiEhAAcrotflRO6mPyfiEFm1BdkPC9z+Ip676duDRy2+kFaY/W25DW4
a4oakkdBhvtvE/gVVFTXZ2vy0FTfQ30c2kOKjRXdIsTooO8Qp6ITr3cPnp/eekRS
43Jeu72SRR8Vbx5U/5WNNRTNIV1SXSn1ZkKW7Hl8bLXgW4ojttp2hx95qDeHikGb
hU2tz4zYJi1NgQU9XFP1AV4DtdfJkZ/285Mv+uxB2PRAsJ4G/tvLFop+vSb754o9
Ce1UeZkU26VOV7mUV9oeigvq7LOpL27XJqDOJ45uOZnG0KLfLi7e1F9FjHnkDOLs
YnnyyElaPqSEGNTUE0SQgwbrlvSHuAZgfV+L+f2BATDNt1h5Ky+s0p+1yoWirUhU
yrsDvPjP7BUWiOnG4zILVDzTS9KWTopa9w5GtH41gMSTjgh1pq9E/3dIz71mxqRH
csuVagSqgptXG7VBOZzW0T7Iubbi4c2dEVohVTvcUyT2aWpkED7AYFlFY52VDys6
D6TYan3ZYUZL+W5i4/wRb0RvI0oNdf9x80PlodsQXYJRLkXcC8RwnttiPPc7oI8s
A7jXaykFixhj72bwEERwRn+hYw+GINBE81OZnwEJ+T9JajmMoqDOeGNsAbMFKcVS
mgjJLnkv8zuShbt60u+khKMzfq/nH8lhGqmCfewWTIY5npXjQLfjkgkVsRb3FZox
7f51iHANT9iNg+95PA6Ip6wpDBeM3/tTVKbu/gmkiL2oukJv6hh7WDWAIrIqzq8Z
5cI6YB9tKGJmhl7BJznc9jBjH78wL76WrTstb7HTdnk=
`pragma protect end_protected
