// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
DmjpLKf3Y4Z95XWWG/YawYchn6NOia7zwpYzAQvpDKM5yVHDYw+Gtml+U1hhd1sz
u2Ipx5/2ojEfPF8qeDry3Q7JsFEELx8FdEMtTSIPfSftVL2zgsGXdRykLaKzBOR3
6MipbwZrt/eayV2tOOrihBy/7wEzxv1p0VVVGPBku7I=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 30944 )
`pragma protect data_block
ohtGnU/Sye5Y2PGAcfglxH6NZX6HOPFmeXV3ew9BMBX8Vyto/cQwe719wNnOilj6
1tEoHmchTjV1DQL6DlIDwbP/iRsBQF2qJ++sb/SYkY5IvBDp3QHmu6Am1l9uURtt
pDlHllwGDewRhCBfrHJY6Uk946YM9ZkydhcvJWmZhEzsVNvE53tG6Nacy71gRN+F
JZfdmxU3sl6lme9pGdcBUedvZ809qq0z5FtzT50wtHTZXwBaNVWriTzN4yK10X5Q
eOonuXPMmunA/d4KOP0kIwpzA/kdgCY2CYTl1VkEXe8iFcUN1v7F9pFy/IOgPhw4
aEgzF3X8OmlZaZIFm4x2qL5OBLhrI//8k7dRjPPurgDlMfn/K+pUctSOZqTYE0xP
mmVXsKNEQUw3KUgPdgBtuOvY8Ugv87tHY5W9EXaNy2nqE+dcCRytSu/YMkTtQmed
Ye6V6tSQGgPZL//dQy19ufZwS+gHpVzCbBp1zoFJIjVzR3r1cB7AzLQKuHvjw64T
SRWsPk21rqb6/3FYW4W8N2h3rpiu5al8FkzToi1/aBuVmQn2HBZvzjyBSYpiQU6M
TYz0dW5RJcisE7V0YTKA4yQ19lklSrIg0ZhSiyVjE9lW/iOiLsDEkzqfOwapXIiV
33vaEjjQgnvuUD9X1JmOswM33Beov9uPoT/nhmErGEL9Or3Hcs+QTX4wMGX8Xgom
NfnjLimbpeuu34+jzhnizMo21lmNZ9gYy42rW6bCiho7SkEM9E0rmIINOkDPyddV
SyB0zc2Qm93NEesZAfjgvt4X11+dPVMBJt9eT7bhppV9Mo32eTUcsenyqO6yhy3P
/zFh7txeriZfDyYI09e+5Xk+PxRB4cM+XkGDsN6LKoWpSEaL4UdP3bPyDVpueL4L
+oAfSfWWnZXvgDDG7+vN/ufmH6qwLzjD4F3LynzbWt2QuJVZeRXuAkydvO55oJIp
kzDpjhYXhBfFSOwlnd+hROqftgQlH30mBNGrjeDqMHhZs/q6+hUkreu3qb18WCCB
RXQK5IQvq4VGyvexxJHY8fArVIk2DXLdqYS1WyG4iazrokWyTxeHwBPRamV+QpLq
hIwupTJKDLswXoslEqHCFmSDSHDy+wQ4hr0l0n8OfkExgmy7oBomprdobPc53sKK
S5thOqu3qzYgRgBEjX0VXvvEpiGFXJijNFJZJO/2SRgeQggvkrFcvTh/X6z/6tUS
CIk28lDrgYHoLO2vli3Ni0PFFyYjQmzsqDeI1jS20danDuMiVAJVeBObP7fvwvie
TJppTFF7mVrPyw0nUDSyNAT9UjQNTeWOIzYLYCtmiIbwTb/wRnkIdI4Sv6RE/AKJ
36tU9gBIR9wIZA8i1VrZJXnzVFGlSPeQ75CwPiiYxHax0DNxIfjQk2YkjT9Z77g5
riMW7dDZ5zkOp0LJbFAa9pap896yRKs3igXwANwngIKsBHe24H9GOcoZrloXUp/5
/2gTAp/sediTPuhWkUiHHEi6zT4hExVb5COBCxazh4lAN/kCtZ9vS29MKwUwtuzG
n+OSCRx7I/LICWVjwcCbuQQyfwrp3t7LtLY94LMllMFDRCDimAR5W0Cl391mmdqU
5zx6bwMD6XVSFAuVBhIIUjlD2O2xZg5RjXmi2ezfW/eowFXKgpM46qiZ0hsGg1tu
lsm+I6G6RmIpitJY6fzBiU3904XgUdFNvMzrM6af42tYjm5YoaqTzcZoFdpbjs5i
Cv7rkzmuKN4AswOFTrc9To/Y0N33Lyte6EvTvNbNY7Q8Q3qnYdDfD85JmJVjG1xz
8Ouvn21q8ZubuY6mHolIAo5xsUenb16/gKh4JFVlJ/YZMD24rmzJfWeohOysD9TC
KyEGLgrlYpaIK0K0ymMMFT6s/imojF1CCh5zicXpcOvPSJpSz7VfjZljDeTGgQk7
b1oTsS1tR2ElDbYJjvaWl32BBzTuBtZxzlKM6INe9KCH3noyuYlNG1YgOa4jufUS
qmGDUAS0I0oMhMBsnh/AKhqe95hyu8RF4DMD3URNvvID6dUB5iWDE3JNjknXO4x0
rm1P8gTBnAB59pK1W+7xt/YRixM4/YS/tR+BFHJmILlYzJzcQXP6zK+6x6mZCm6G
E4iu4PPc1rwmq60nRuVydK//TTPgeP8iH0/H5RvXeQZ+8SANvzESSD1J3I+Z/EBU
coMQf0M9YJpWNcPKHiwrct1HMVY+XHmk8hOAg3UfuHDBaPsxxvge0j301Com7KV5
iYL7owKxNcGR0PmF/OKMMqPuVmbMaszuIh8waJh3P/jPHyvPAjVHtd8kRlGq/qKO
qgdUXTYme35bIpHm9+VdHAuVXTbsErccMDvFuc63oIN5bMCr8YjZycDxrc5T4lBE
olwNG66x2psQVWHkONXX90h5qyWaytuD9GAvHSz+QQPJV75cgdBrPvQatP5apHJe
RFXyAjwCWRLSULJ/cSeb3SPV3ZRaYL31OpVHV6XHEC6GooOD0x0nppQhhqXp9huo
3dFyj2lx11JmLHp1RhbJZF0yezaISHWdvyWMdLZcCZcFPkScXcGua6YwfYGJIWiv
ATwR7btDHBSf1keRQloOnKnlcg1EeTtYLF8h20FGfb27Ckk8tngz82XLcPnqM7mn
iYZmphiPXnyI3pQr4IB4urlzpxyBvMYf37IKN/KbVd6nzzjGfU6ZoiNrnSk4opjs
8/yXF676LqjMnuy5oo1zy/EaF3aFGN+m46Q4wUyaPiBZIbgTjRpBCs5Eq+6guuk3
KBiJwJDd5gggqSTgF4EM/QDCIozGja7LRUFq0sWxCPbnOQSqD6jl7j6ngXlTJTuc
HNKdaFcf7/NJPpuOaaVZ4Ejbviy5a4J0aV5ZFw3kNKuBxaHJC145GqwXOEZHWJ/b
bguIGoB6D1IZmHOdUMc5RrECFlEimOngWQDf7i7ZO0L5oIrI9787IuLpoHlkU6C6
UuMXZa7IBHw26x66eoybnpe1RAMGCzdOHdAe4Ap5v8I8qddx3FaiAiTPRTwDRhgK
YVShwn3hGlL6O+PmfcH3le3mOwrU/bWZZoaB1T8ouB9tFItNloAitb0L6CQkJNYf
dB1p26KWKEHOx492xPWNsfBYck0iB2DBrKvc1njimBY0ZntqgHXIKOxPPHTWPkFK
ZYFkL/T2TuhwJ8Jg6dKT2w8LnG8digJcbKK9nKckRbY/y8PyacsjW5FCtrH4HViS
u412tl2MAyJ0PQgUodyqtT3xAPDOsASe5IMinrdpPcsBi1F8I1Oi60QtONuI+l1I
jVGWrts3rJbpypuAg8d3gcPnhSN4gnJv4FdeVM98IPUE39LZeQALoHbH9qDsPs7p
gclUKsue5Inj3yQA8G4tzudMsxVQdxeCgzn7tfxO3BQfe/iMQJEsqJh0DiNsMs6j
fUc8k/FE0nyS5k13SnpFwosfTP1a7Pfoa9twZabvTOGHZQqAom5HGgzwU6f5+ysA
DlIkD2cUlHwpVb0ujc8/vXdBdB3c/5rAQ6vPun0C5NAiuN3uFaO+CRDgXc1Tsil7
6q9kRy8SkZGZR9sSfqfAb0Qlt8FAtGYSk1jfJ0gKWv0NgVXZQ6/mfHFLd5bWBXJd
GtW/CDcx2k8MVta9bj0sK2V1pgwiLtYjNhf28v9/ZJ8SeREyUCVc+1E5ZB0SXRNG
T3KTuZFSHyp1BMWd4oQA/9D+S4dktOzzKsYXTN1w+8lrrp7st4Ff5jcxuuRpo5jX
w/6vhqGCsIJ1XPjVLanx0KV/PIb+FS4zXiX0Q1jpxhf2/6rbJcVBH2zRNTes02Pb
35d+6CDJrlvpy5OurrMgJ/jRsIr8utj2erfdP+CyuLw5y1s/ibBAL4rIca82HQks
HSdXADIg3ZJZx5or9/LEKoiJfgdXqpfqLATT9G7zn7Cte0WmXO7/fCA3jUHVsCmA
zyedXSl+ft+oep+AQsp4BU7O0na/xyIYMNdtgkkAfLp25wWWE641Et9/UrCnsOZt
ukvoYKXFxYtXG+YOInP+NyA+HHQS7yn4Loe0ORQGmkjXubNw04LD+N8ZuEoDhd8o
L7S9hFSQcMMUK+t0o+LU8N+ke5OZ7VI2HnuHvLsmgjRrgFwVHzTobVWIaXRyxHnM
gpYU7w/TrcKY0UzNbfXtZIHdy2I4ZJIDm+rou8O+cSH0Q3F5OEPRRksXXeo/DGme
EeI/BA0AUeSWA4hVl7MU+awX1FXPtXtR89hSYbdq1loh9V8E9mVgmq3KuUBEoqCH
VyKToHuJB1tOj8A1acVkmoMDaInkdKJQE7sjedpql7ml/retDa3GzDKVw84d1+kF
1HHDKpSitd+vDwKNL7G70YvehQcd65+yXpCMSHT+e1rIw7vGvBE7OAQqJg2WwZtL
cop+L7c7IP2WnRl/hwE2N3Kiu/6/V0oxsmLYlIu4A2jc69VkR5/MUIgsyp3jm1Gc
uhsPfGNJaT53ICzYvauWlHbX/P8SNfRFypV2tPcKDsdZLHmsVo00+RRhyrDCMmyz
PZkTI243s6JXxRdVWlzliVx9lPog9sH3mV37jqxoWZCdXpESzPW/duuNQbdUvq0l
YVmluJ7fyvCM2wOxL1R+er34jHmRg31jjd4I00AjqDtsuQKNItRsVi+xHamZPwy2
/mZma3xUKpQ7XzuUq5jJnFOrXBiMtxXm5tyIkUQtlGKpk2XZlwe6TgzU1gGFkobA
DmQk6dEbCDkwxVq6uJ5lkll1deSMYivCdnLwLQl3AJ4SlHOxZjMPC3H0zEq6uiB6
Cfj9D2+MZiFLjvnTB+6slfNNHe34jO+kdRPBT5IKjUB1rYyE82X10v5rEyRZf1Dj
zBNhAOZgN4+IGEJTCeG6hXEwRaGrCCYJbUIlGG5OwgB0R9IowbbkGq0B5osbS5dY
ucLEMzeu5Z9amKrSVMPdvI32CtFAl8bxkRmvAMRprq+N+0KbuRtyHsw6u7gz8b/h
Y0H85T+FAle/NvSdrVpndhUHGunSgrM/sl9k+n3oYvqcIYh7go+GjLps2cQ/GC8Q
8PmhaaDMIsWwzNyqR/JKXi5Fxf4eICdCZWH6IjRk6R7zduFfer2Q6z67jBQxjs6k
vVTUCaAcKvP6SGvYG+3FKz0tFGCd+ApDBV1gaqKkxOJ7jFmcmc23iZo5nVugBqvp
P+HiWEVGyFwldInT/sDViIqfHd9FACaXGIYEzbPkF4DUMAsSVcLnqoXrbGJzPIO5
bJGKD/9h2CNCmhEMSYNjKWu83xc/iiYyLr85u8RC0+Krv+qgi9UYWJvlmiX1L8dm
I0+3GuvvngxyIrzzwnXGYCEuB/pRfWp19a6NaoDLojfgq070Gk2iDKChZn/awRUZ
EHDzv7kPYBSRmMb/c2a4naPnojA2atGXmI47axDQa+tZkszsTgNZQdEb/DQZcNCG
Eq2tN4JYv2U6c/1PdLdLfozgpl1Ujld+r0b6XHWNEB7X7HiYo7O+k7zlej0a9aYu
qziRcdOTKP3EDTZDHl55sM0a2NEq9H8ENws2ptk39wjdXjM4D7DtnybYIrF7+y8f
zW4eAek6kKCj9Qc17ouQ9cNUl6e9yAnSWzFSKaVvbML/3B/zJo6uuz1ULVjYzNi0
GfbXxgAExByYqOZJ7MNMV1Fb+umjxLm8AXhjaPIe6pvaM5lhIBivsO9xgxjJ2WnX
sw48wnR/zNpEd22VJoORC/WehFDdNfq0ppRPG7kPQnxV22H23Dx9XC1CtXd9KxSW
qI6STacdrlRoeyftkGsWgqW7zD0rSS4yTfRpP1LxUe4bIq+/igZ56CtFC0gAGhdI
KT8jZp7X0Mhxc+SHXVn8Q1GLPvUvArxG9Y85S9USLKffeN78qb02zYxCuJDko3HX
BYvyhCUG8LAQSk5t4j5IZnqrxCxza0onxruMwOxda3D8AaKSk/3R7CopMx/9DZo2
SaXmQ/hrfUC5FztFeFAjnmowkT+lg6Nyck4CU1U4vIZDEogFyoZq/qqnPknGQjzq
WICh3aVGDnetNl+Zel8iU/K5RHU+rr0p75X3hU81t266IjYCfULGKe8z6uFws5F3
G+Um2nnYvGZjP/BNhfnxavj9nbyeAUmJVxP72XS79BzjxdCa8R11d+dDqJuFXNc0
EpZAQdUHahZI3idPALAR5AL2ExW26yIsAKTVwuWjflbNEnHqPCzj73dWWRP/v1Uk
zVu0cwTh+ROK4wVN/loVagLSCz1SKLjqDUYhLRpa7Q2nFr6U3TQLCJmSYvm9VBs+
QRL4JxfGktNgMmqUqKI6/T8d6tDlt+gZlwdvw8yDOR9+bv5RVczuFPQKYMhQalY1
12seR2/zfvSugTSo/dNL5jB3oKAi9QuKNfkJdlYyjxxYRJykJzTbHmlBH1Dy53s+
n+FB+5P74HYOv1khoL2NzZGHABEoSAWkhBxGMyaEUaDnE7/lIi7UF7/nyRqZfLrw
Oda3rWvz/B4cOOwsyKjub3YlqHzG4wce61Zgb1IUbo5XetM4zIAmJ0IuzzZ3YwxO
ieVuUZxOjLuJm9vgPboExrik9LQFEgZv94l2TqzegdKA4BIghhlx3cNnVlqXJGgj
LVcHVOoEA1fRFijslr8KQyG+qfQqp+X6bDD1uPFvHTS22DJIQxZUY0M7ZzULtQJu
+hn/pSkbTgoCXXOEhfkSKpSRuY8ii24KN1C64aDIbDw0cs7Mltjc4jPBlPH9xYPv
VywedrISyvPZgqQ98JdUsImZCjZ4QHafbhqJqMaOOSAeWTVN7lawAeWGor0I92nd
kmdOd9Hn5HSVQNvgrW60zFko4LVG1OHwN93zP9ZszXlyjooWAf7X+EeaMbaCBhYY
2UVU5ffMTW37nGBx/1abv9rdY2bUorpM73BK7JSRCgWRmDORkT8CBN6lllsLN3rl
Q/exK38/WjR0v5NOaAeyXpzeE0lxR9L7GDYyURoz69Q9sQRSa4D+WYvhAlVfJ86A
IVHvSkgYzW3nG3M1mUUDqq1vC9XDdgLenbMgjlLscmevDuxN5jPEVoHfOW74gI3x
vVYAs/Jd9wzphOX9V6ZxNxMKWEV+6dlqciOvHifLCelEGa2ZdFWL1ZCBKkSnScJ1
tV3ZHnkvoi7tkMCXh0kyy5VvYOix+UvcOZ+M9J5dqsB8tofZBhxcav1DKUNmXrG9
bDyIhRGCdaxDjLBnyqGz1HvpUJMWOIH97ztiyD2k0/qEbqmlSPohAeKwjOxIkKKG
3Vwoj4oAX+2weUAq1NrmLQHH5PrLtkftXv3WamY/9Z+tUZwS40J0zXIlousWuNgR
cz3K2KF7KGkrNsjoqfPPKxcaHmA6a7q35UozJaBXWNv1nDBf/ENTFN4n/jmZatds
EzzuBbPXFXB72A+lRcJCWaejUr+nW+g7KAPn3aO8MLy4oCrQo/9sNzwwM53DTEuf
//JWvamoaZXVy5zzvBlqQsK2E7NUUL+rjpe0O135SpeF311rkOvyOPCU7jpJDzbG
yDLF8gT77JB8ZGNgcv5ri7CCTa+8Pz/SarYz7kEY75QT8f2v49ZeK7i6JP9xtZJc
PjbwSUC7pI5Yzg4OMc2C9sxHNtE/WM+UiXxupWddicr2/S4cG28QSAhY1K5D5Sh4
NFWy8PGvKKvwP5L973kaaf7Zk9xNUpTW05ZJTUygmKJiQZq3s1omDEgVDUYYI3ej
Cms+CelMO2s9mrDijg2YGjYTYAp0XgkLTBr7jGK2PuaWx1yVTYV4+1IE9Sh7ePHK
eVMZnEM3tEFWjJ5JWCBjGWZ5tL/UlggnaYIIpYS6nkRQgGs3U66oLVXquDj5GnWU
5Bjkas7JJSgMaarvV227Xgd9LmGSH8y9Oke7Vo90gvGjOPezYzCV2rWECPKu+7d3
6l8nhvfJL+9WkCrL49BjOaQJdjwXmO4/EfoSs6wjovV+kg4CU/Z7z0EkxLEMyhjh
DmXqinVlG1PVZrVpEdXSIPln9K8mA5rjV0SEq5/mGPVhosxuMj8xfx6kl+GvZGxn
eah1Y/vfcoi7+hrKZMqMkEBxoGxWvGsXGL1cixQ9EIXbsRcQv97DCbLfxbEvINk4
fzmKtpdFxaxxS9nFt/6V6d1AwPfWZKOUTE91Xn30Uiibbi87s8N3EfGfZgBnfp/E
11xuTq/wwADLMSGnDdakfbfEtuk6j4Ju8mnoNkWGXH22M7dqJ/Hs81Z8sWRnfEw0
PokgXcv9nN9LZQW3/X6KWzzsFY955IeXJgohAkZDVe5tF+BG1XrCRH4lkHUVy/5/
qdvzWPd6otofvmWv74Ldzy7hkNa7x7mJmNX4TN/q0aj4dQ4ZNpto5j/O28fOd1vH
uX0KHhTkGB0kjgPsFA3m4WT9skCr926GnqBVXbJ/UQkDaGRXif1O9OWByFbPe7SP
dbTCk59Mh+37g0zFs3bs/u4SirXYxw9Jl4JvrsAHHHc25LL3OiTL4vj4CR4sTnx7
sY6HWPQ+rJWyefPwm38sA3Ox8F3v4z6KHtntfglx5owbSPogh55l50dSZmJlreiX
Qiwxy0obfDo0R9bfF4KTiciCgRJuBe9fpMwBSkQHvIgNRk5okRUvrIpLmMjy0cZx
DJtCwDzthbEnB49NgV1M5q5n33Z7E/1Irx0P0t4nEjOxfuAiuPHoxCEG+ALkoIO1
7cpqLfA7Cmz3iIxSeAQdyUkjW/kde0SklDYQTgOVvEDZpcHFQVv/hOj4Fx/HsZ4G
6JLe1quOT/DqD0EciZsBCxLT42qsLsLSTdSUsVVXw4D7V5bvNLUGD85Rv8ZgwdN/
s/W/28zUCMrZDQIRji4rWCJCkdnb0QhxryKYdmGcWqvwY7pSSAYwdhM7tve3zGAs
45OPYMDTviYcSSOD9W8GFtKjwLDlduHTGKabhX/Q4ntWdM/ohK1hZ3nkgjA3PUwb
kyUmJiqxC3E1K26l9JOxYyI9zjatd4/q1cQmWue0PLyfhEPCaCICNMR2Bgla5wKC
VlaiDN14xMroelS3QGJ61jhvNsIZZf+6zraR4dJzgsncb8FsJBqg210cnWrQsfmR
MqBY0sMOXmoDYi0uJqKrUe/nSm3du02F1FPWk2ySDLlCpYgKkBWs4d4T0M9hNYTE
uYUHOCZLdvBoT8zcbd5u9Ja0ZkQjj61BagrcQOhetsknKneYndrv70T85iTRkMvi
wXIEJpR9NPKWjBrw6Smu406ZA6AG5pDLSJrCX3vou9S9W+5k6EVrY4pBXqXv7KTS
nHfqNCyuRRTWUy+V3vSY96OzU6bwMaWJhOvAVHsbgs1k3lkjc+WWB8t306XEWbHl
pkrxdaS90yn0MtqvId5URb2sO4IXKGE+0pirAed1NHzeW3O6Hfm9ijc6upXx9fXb
VWCQjbOtktKJkSjSDdE9d4tv+kbB+2Br2tOwUfQjIeuVfF7b79UiWZO257P9blE2
MHPsMIIpoY8WyRPnGHyiXqiHGzcuDUYC7+Rs2GCKGeyjDDdaB7P9oYv4DvyS7dBe
SLI3FVMh58qneyb+cjUot15A0MesAvQebr7z8zoAzQncKvfYhYNZ23LprU7Dlxfp
BwS4GyKRlT3AXLd6Jj2QrIBV2/eLYAu8bfCAs/LJPS0BaQqqrNmpv80RzrmvqEQe
ikVk8NKPNrXrPE8RFJDsc4spvEnBryi9aFZ5EdBuHgYrZKcqleoly7tvt4bL8/tM
7Rg8DiayNzskqy0apjcCkBcdlPxOxJTIRmYfIlku3l12iTwAEem4iiaEPqX35yIr
gyagih20uqlG2CCnVHb1vgOL+zZ5Nt2OGZRf+uW+LvngnpMoSgoOu04Mkc/OMIWN
K2K0+M8WrEz9hSSpvEer808eR72ILcMrrAnlAU4PTaY97k7iIqcPgjRUpvPApaZK
f9vR/F75s4U1sxGLeP25jrPqqx4Jwt53Y3lvbFblCIChIDx2POjB4Kv9cpHhs34S
t2od6bt9LZ/LyZe6m0nPV6ZQjo9O65HbsOaa6xY4efsbU19tt72x87rkdZbgVPMF
mb88ZoEZTJUHGHlQIdb2cZvlZc2yJxRyNe06XqwMJZ1YvK7p2WGEaUMob/c/aGCa
h7iu8Bi8FxsXgS55puAKEPn9IhgoCEtPsmsM0TbfzgDru2cLfgvjqfe2/jBsYcdV
aNm2TLeZyIZIaRgbSk/KEiJhznLZxbncEPGIjukRObCnPGqazi9wNhGcqdbIDp5x
n4Ive6Gfuidvsm2qr4M+tLtPktHFDc7W+VcnP8+F7GksNX/UOXRUHY9a9ZUehYK7
rC+jH+ce/TOBoJcAEvF/NHEb/N2Z90fJfMC7WTqy01jJjs3im6xju/5o297/cIdu
nq+4J60jaY3UW7chEq7zjJz//X6dIQ6kBZSAh+Oh7gcYOjmtq8JCdl7ugC8HY1hf
b76hITAEvI1NRH+KE7dy5UkHZ2SsjQLjykwgD3WwjbxfYIBlj00bBHoJf+MRo7ht
xVSa0C9TBqh7DR8oa8N80Y6nPOD1g2HBUdouY5MLwTD0jNIMFIrAZHNyvxx9Srt6
sBC5+YLkIgCzmvlgZcSIK6OjRq9tXpzjTlIxJI2ejj50zqOLqmGnri8214jAYBDP
Pq42p2DI2rjBOmWUixMigPtYLMOuQBZbQyjellD304NXic2nSxPCBgsQwXs/rRPk
FGnoyN6bINuyHSiIHakuCKri4+Fo6smMu8Rd5Go9CYyeVfGegjtZoGLCPqYnMogS
h5n+xLD3ESMTTdJulYXVLvV9zAxVRttZ6qzz0qzukAswfD+BFoVIlIHktMWqjIH7
MJOfFs+Ji/sW7qqBN5Ml5zbhqetBrZyE6EJ+yp10QyZWapIt8Ew7zyEI5kCgtmHg
yBWCjf3YerYoh2qyqpLgkGDxjHaTDNXt3INtIyhnBP1KLpDePGmAeGUnPhEtI7ke
JG5USkVenCffzmihPEqGR/J+ujq+y+odXUkL7M3GCJBUcv8NnElihn6ctXzra5jA
FwT1yEQHTPDSM+iaLXqkCYr8ynGQ5YAfH4QtxXQW51Lfou0PFwQZyyxYfoTSLGB/
lZ80zix05NzuWsXTSoIugoZwdUV0ybrAZbX/o6byxvJrPLkmAmc4BAPt0GpW37ma
bssZXybxVtR7AErIsaoYNWv6tJ2XY8FitomvhjXUaoxLkvljzoinm1aGcxf665Bp
CSwGe4J1l5H3h9OCuX4Qw9kE6oMSn7rJHMDbd7C1Jw3zUxQSX2lbXAPEQCJUXegi
ltCOfbV+rQx/Y2v2lRJv0u7v5/i6Wo6OvFv7e3/osQPCTAckRCWKQYeHcJkpT5E1
o3DGsQetOWTwMVHfrDm8k7O1HvefsJT16+1b1L7eHcQqBFMwwlwoPP/ofR3Hng7A
Kp/7p5vLORsuzTzZb4vPrpL+EmcGylQCxQO2/LVFeOGWJGLVOXGoq7sbYpll22jc
MkJ+/l8AbvhLBkxHcIQAP8vGQMbJnZ5yNibK+K39gGU8tIyURdWT25EUGqgWbQVn
oq9p2LzFp0WHfsO8q0LtDI+rEADe1kWGraCcC0DVnlA7swXdtcgfBvdStB62NRQ+
tCU4FUkfZ6FF21wpa3e7Jc69oQS6r/NERgNHl2otf+2OQBSgg6daSE5ANhZ4YjIi
nkeJPDy977Hu+KBu6au0Bpagbwyq/giCs7P0Zib9Vk0STx8j11TM/zyMbf5g6XuT
TJ1lt0kOebYtIz5+oVjFR+Hv9+HQX8QaOFZMga25DvNooWr2NpNaEVahZvDxigQC
4qmIMubloC+E+h4+MqxBvQbDVgeUiWB7Zh7dT+1iVnFEbjNlHJnZEJJ+v6PyvVuk
QECBaDb+Ban8m45sba5MbaFrn62QzANTtcVCpAV/7bBxwydmqVY63+uWj3hvmwLA
9vBGov4P9QmhoYAdg476F/FUhY4cYm0aOShRbXHGTXwGWG+UlbQltio9UrTJ3VC4
82O2ANSDQtnM0mEM3Xy1/75l00hqpkeHX/p+GUv+AQxabmWO3I6aKBHp/2U9xnaD
c6QOLuUr/W4mqSiLpUW8/tbF45uujxkiEm+CSjGn9CIRuGU5hjBRe9d6DRt5s12x
E+VMjYPfsGWo2EtzHPTh/0FbC5/MCynRdF6YsSdo7VyHNJfNYkBx0lpphw8EqXHL
OLNf1yOPcG/Zy1CFp8+IwT5NHRPKigf6w+SLjWmFiqWSayhImjLNoIlhImVahOdk
DJnKRD1HdvNp+kKhMF4bS7gdYf/buzzKt+W9burFIA7amSSlxPIpYOICXJnpNAOB
WN8/9Fwfy/YJ7+B1cmzGfad/zbIFmuTsIt5Pafy7wkXlQ4nYPFv+Q/7HRP7CJQus
K2xM9ii6Ber+UANUQPuG4/hmdrts6n0GPZz3ijtYMXafq+qVgvHpEePfRvX8UwNk
cDBsPVhZQv9K67lGLCang6E4twUbKaxsQfUX2PM0VWNN/cQN9UbFhDh75RvzNCNg
Cl/Ip6Gn6TiQoeIDNqu2003TFusSPOONYFPwgY+iw5owRDAijJkx3INfOysSeE+7
IhkUKFToAyAocaCTzwAt1BpVuz+KvQHH4C7OVGx1nSRXHdLz0Y2YmT0PgQFe5aSg
vQ3q9Xx3eOFvyYTjhfb6y0mOIR3oa2P2T8w14WQZWP7MO8Ot3HcrKziM7XjmY0xE
L6d6W6crQgRH/6RLWr+kf82WfaaTYk1k9+7oKquql/NsAw0RqcN62T7KEH1h1NV3
+JAO9GNlJVSK9z/BbwEyg9Eer0h7rhwqiVSjedUhOu7iHfg9d309xZ0GmBlrE66Z
bN/l35gx8LKt5zl8LqfORybpNnFST/EDBr4oMGDYX2yKdnVj0yyz6O+dty1wu90e
FlpM6JRqbFjlDJ5laGux86WI9jQadPjp4vVHPS2LO+TS6K/9RNXYBVU9GhmlbIaE
JU9SvnCxnllO43o/myi7NlEc5RD88OXpgErWWQJ+usvrMzqYQsbMVyL0epTM6WfS
iiMxtfZ4uNFyeahfPMvyw/D+lV8I7xjnPWaTBaT4FkvLpUEhLg8t+/SNZOJfOlgQ
7niuwbWZJicvYezyjOB0iToPqMg5vFq6EjFCeMhIA/2o4tAS6yJLuIwuTO2xZc8C
311Gf2bw0Zb8IjDbj4dIed9vq1wh8zESCG+EguQtlIRmy2yi26Al1Ju+HndaIRsF
0DdbZR9ooaCCxyNVAGpahBfJ/gmXHHGBTGv3NcmgCLkLCMEyaiKQ0l0XDGB0/CB8
GsVMZA0xfYyuDCCn43q1fcPORCz2nes8K3mnWGfgwTEM/Ybtjh2Q14f7ExNDjdZs
bZv4VudWFVIg8btgfQfC+QxZmWHVxWUiKWkDTVBrbpR/FZWVRKfQqzbBjA/B/uIB
zMIIFU6IPfkUYfMetKHJrQ0Y2ZH7QLYtq93uI6Iq99STrQ+1+erCbUQldIGYRzmR
nUnDpcSwhCG3Pe2sTqfXe/lv3SYeXjiCCFsxxmNDC6/qD8rlBCCiqSVEoATUziRO
sMd3mub1AEh+E4ot6qap47J+r9wyXMOCz0QpOdLBcJ44y6e5eAGFlZuwKYEXZn+r
2QVznXROqWOzw8XnzOG1/BCog9fbJmYQE8GO72Ze6bFebcZLT3kvaI9NRYtr9LZs
z4IDsOAcsksw7sUpqrHVbu+uMg6q7hxlquEmUehePFB7WquT+Bn10wi5RODOch7m
MqkbSnKyAHdbESYs7tnu6lXlS5GgyAAYH22th4OBDdBBt7XxwmahECqBZ7G2ICDL
QCY/KQzr1jOA+UJ3STaoOh8dXNK0d2zckojen/2vo1uaJIa/gu7k3i2TxGBYk4I8
s8EhOU9q6d0sB8rLbPeEFub9slkHWJFLq+9jtB2nX9yLb+bsT+Im0xYfFT8ccd7p
+S2R7SrRhAEmYUfTZh57wUs5F2v782bZK/N5qu2j1OoC/tl5GhuXXFCPET1DeZZY
W67DaQEnabge2M68Ws5VqOFmozHWFBof1k+5DU99VHydQTcPzsXoguzBCL1jkXQF
F+/1+Gz/9lDaSMP8FGxQFg/XgDtG4XkNRfJ3bJ79XtBoBBHnHK6k1lMHDJMhtJtB
n0zrOHR+XlbNKqE97dixB94c07r/WlTQX7IetxtU/MWx71v8bfr9IiONYkWSQLev
wukruqqCuHaX4Oo2iDu8aDKrs/rg9sDleUu6hLWFQ9B4yoSK3VmyZimOjqBsNbzT
iu9yyrcl9K/6kFoT96TmfKZG8ek/gl1Jq6cluwi3s58xTWtdUkuz9/gCSF9MZT0S
G2e2qp1sQdzcJFoDrlr81mEKj0kbToSByaob7y+birGU6QUIUGtaZvc78CLqloK2
yV29msrwCRClqSiWIgE3JveOiq8BukHIKgH9BoIqnQ3Zf1H4giGvAVr0899jJDs5
fburRTGGujhQ0rI7Xv6ognFTqEXS+It/DuYAv0OTa3AUvr+Y3wSapK9nhhJagtC6
5E8c/PtpBrgW5Sj14SpVORwOGBGTTgoxJUnl2hM7wcttbKbZ7Ld7lmjTdoP7G/Mg
6ItS1Djmcjiqe27exE0zjqXxSXTGngxgWi5Df2aOMsreQYMPI6CcH+kXPHaS9VOm
WCRCW6bGXvSCXVU5yA6//zvs86Mtr0J52I4M1SHW0LTx6qzJAfZFob5cqreL5bwX
Rutum6Li8QOXQ89D+MVcazyPs6LpJqSe6cwwK/H1RXlvVM0gZf8I6F20mAiwcm+f
e/yGXtyBiP7Yh0lKWcUmmDxaZwOdGkAsMwmI4qVldHOLdTE71rB3N4ZFDfHoJ1/z
yBfnD4saYhggR6fsn33DcuYcrhpdFkfNZCYfCThxFCBxb3c0mk6zNCYRlklOROy7
shGhdDQ51NtMbqqmICKZwVuZXraU50caw2nKISNxJxvlmON1qxo1wDuI2MlpTAZ9
Pb2hQQPHugP8eKmUUJWLLZtm2WDRbb2OAr15qNrQQ5F0uin0CWPDL08Kn2m89GZK
Qh+u1xTFI5zc/X+5YDcTKhWqschb5YfRifuFQpOk3qP8fPwGuD0l1NS9kMiHaM8S
T7dcLEEA3qldtgk2fSZunoB2TT3dXrnv8bx3fXhsi/N7GBRQkC8ZC0tOLQV3N9Iq
OJQhJqZ/F+uDUeU1LIU8fpLoPv0dARytPVJwOb6gpiYeYcFdL96gJ0os/d+DToNb
P4oRIrUUTiC9TvLArI+d8SItfofWfjTGLL/2GqtgMCp+DiXXe9xnuUsm9uRF4YD7
YoD4WK3qlhmBIk5zrvBTkSCrTR/FN4VWPs+eal0sausFyjrEbWfkiUcfwFMCG9jP
dXJR9d7zTiHyu7FeMIGzqTUYcL9hYj6EkxpRoxetxPv0+qC+ZE2Gh7NlE/XCpzNp
A+MGkPorZ3AHHD+Ddq54Q1pGPvDGe6PkIvK3X+ZBYOhkvFg7Ohov8v76OKzaRbwd
aGesUu1oRGNYb+hQ7dqtalZiz83zLNxlA/w7Q68dd7Or88y0DrWbuZE1D7xbg33x
fp24sBFnYANYtL5HSqe/MDRlrmUh6D3GVfhTnL0WxVu7MfcIt5aT6O7Ks+MSrMyi
ifUcFNTty8rn+vubLv7e5wni1B9g2HIQDQ+jA1TEyIzrA/IDP7Nr5lCclXZh5Yo+
nHCfs4r4n50IZ2FRoKif82SEWQwKC4Ji/WcDnbanRE/778c2NR8fLsN5CILU/ae1
UIsFZ/X+QKYW58uQVGd+H1MM0iRfyq1s2Be5+nKkCmqdLnGeZf0n6dTStBC1Ftks
83wdN1dmmf2Pqn/7RqtJLCBHT2zoeJp2rKrvxb/CTKuNn4JAB2v7w8X1hYFhMrqg
W3UjEdFZp10BbXi2wwdvRUd2UlVj3R0hFB+7Hpj5VecyHMsCJDrrjQIhxBJ6P/yG
Hid5oO4Vd8U2baw3BLfvsTtThRamA3s05AokAaaDfLy2wB/ixFO25XsD1DmGDVCg
SNiDMNqB17HHpQkdnXZhPT4HGIElGj9PA47fPjoNX5zbZnzHBmn9pUlC/yzqbbkq
+jvKC3kc1c5BvolDEjdLT4pYQeSjGI8ITN1bFsjJfoDOKqrYDob55niQKgsAPU6r
OpGzwh5z/C6lhFugLKOcqvAmyGxJQLDxSFyVF47UPUSQoB5L3VnFDLMvfdQRNLYs
JC3DkxYoRKfyUiiQjA9gUa8raBZQrqsFcBg6jVXUREA5KCxR2SKDqxs8wZF9C7HM
eMfxspOlyHwxw48ZwbjX1HX7/oZ1/xgFq5Xlbz+OuWfIuqYtXkqd9pLmcTlNt5qd
xBDet7DKSHzIXVHNIujHK45LajSHhyz1kn0CUsN9RR54sz+4YqOB5aD/PC5JgCuI
U0MMsrjjl3SvM/J5ONpC1jurwYcHGlaTiBb7DuJM+Mm6bOqZT6HR2Gnzq4rx08UE
lX6+MMQH6P5t7zJCIGZpBQuDvgdPqvssYWb8SFjvgxqyxqUZ2M+GEAmJbu5vOO1z
dx080rAhbm9VX2GU3dIq3V+pFBuZtvSZHr0SFl7MQzRhOsdV4lI0avW+6KcdskbM
5UlOMjDCBuyONCBJsN/waU2qMSUtBMaK3HrlBES4nX2yFfdT8Zhe9x+pXbAVqNIM
VK8v/GzxzTNuAe1J55PovWAAWjH65wKXf3RSeSiCK/cpZbn5KT3XBlQ7WJC1k99r
xkiuttsbPyT8/U612NfBqLdTQqEopoqfKj9yvw6+CpA5WoPunVuo4tCsJlWxByXj
ymkvA+mYagEeNn9Ah3394D8Vn7cxrr1L9B+/bFleY/cr8RI5i0hVBLI3UVQkZ1qF
LSde9FgfH28SkhnPcFRfgx/Z21xom3cES9tNl/UJ7S0B48BGAaEEuqANal3PafnQ
3vEd+Fyjl9AjXfDENJ+GSDzLnNifteYSd9GhWRTs8rRKln2yeTyB8YnN7vG9NymL
/wqHlHYbubvCj9/zOKmnizqdW2CJffWveAZ/Ev9HaLejefREi+BJGn7fo3TtNioD
LHwbsfACK8qF4il2ThxLb22rL8rTBew4zytt3mdMZ92IWsBy3mhO10e5ZSzzvj0A
VM4QxmGolf2CIb7VrZJ/Wh762N3Va7nxUmWxWdUUPyKsbGtsd8wl/L3+Gl7pX0KE
9uUKSBPnFzr0i65QudVdDxQLkWE1tglJRJjBKup5gkMmQkLznkPFxzPoFcCJ0R3u
Bu8X8tyK6T0P2v3vLnTWyfIDc8CkFe3Vss3YxnzAwP4cBnzsf7JiwwkqyLmsvIc/
9Jmx7RJmOslGIOyxAfRCputppReO0+wduqgMYktKr+d3wFOoSDh11lcnnD2fMM73
tzZ9Frs4pE0vEZSqyDdXPzJ2nLzvWuFbKau1SIs0GhFjyYDF35lBM6ytthlff2i1
e2oUdn04DZoIsAv3b0qBFyF3NZbqlJd1Fx5don3pr1DDswEt44LEzsXEu0y5UlPL
55ahL2xGs5xT9QTL+TRYasr4qRmn1ErwsEC1spMWU93LsHIwF2Cx7SG0aknTfFvY
CD0+P2K3BeDwOO5a6L1imbJ5fJ6GP/7tkXGxSSHQwASLwBXKMyPS5aID9ng9LTzK
7eNjCQ2uxgtESz45ELyYN73SfV4/E+/0nyD/OyIR0n7lcahqRypP/XbJZ2tMVljx
I7kpln7upX9dPiCHteEaMEk/aAAF9ho+ktZ4DfPVyXd9gGC0IVZw96OvOrTIZ0ED
eF/j7ldF+T+vwWTN3MEInCkDIPdPUsJKDVO4QqmYDz9G6xpWolyrrxMZqgv/V6BE
tFt0qdLkL8slYd5IlEEVTZouzx2U/mx2nPMFeTIf/e1xiyH4iRdFAFuLG33t4aWa
DofxiiQsNH/06mXDv6yti0K5ZI1U+1ApQrW9/nra48aahXyKUN0WqtmU8N16yDuZ
fEDEztwSG05vtxYxlJOaucmJD53y7NoG6nLBPKsgWvca/X+fi8UtMV8WQJ7W5Fgv
QdglOO20cyxPA/6JUdL9xTBp4rzsaLtQuIp/vhlnwbyesd+rtjspeQGUQaMEQeeU
qD78PxrztgFtGg9jTFCAsaNDo/pcf6YxojBa1IgHrmwHDw6V3cWBe9baiOmHCDhW
4lgpZas8wExh1q27RUshWzfu5ehMbqXno6BhxNymqPH6u6h55K8sjf+PcAtU0voo
K5B414UDzZXfQO6OyBM9eMQoXOCanzYtSMtn4wYXOTMPGGXg0rROVBjkOGK+6O5Z
KDioJ+LVmqEL0UjUs0oyQQT4Ht9fLxN3UzatqCM3PQ+DxFdCaytqAQ6dxqgX0PUk
oNbHTGKE/W6HR13r/4Q+U1GXuxkO4zNwz8kJbkAQAwyQTQB4FiN4DU1Lst9R/qyA
KwlB/0ejxqrTGG9Qx5KPY932aO5obyhhWl8hemtOI03cHafIDIFo8h/2+TZO2COb
ubDBbqp+25GpXw7Zr4GAUnMYptXNn5O5pT2yJiSUJnbis/41vJV1HzNDgXmA+N/Q
/OjWBLnH64NQui9XrCBPOkgQsb+tYazehxmLz/oLD0IwI/zA0my+mnCGWQI2TxF5
Vq/Y8ssMNYkQB6b0Euxcy5OkzQUzldsfEHUfAi8J+wFKmdM4ODS9a6SrIlC1KG9P
fyjS4/aOkUuDLrZaaRt4F405voVaG4Ufs88dYGKjUqGDISywfaJc1kYvh06Npzaq
luWyqjto/SxaDk1R9HnoG1/t5s7ey1gDxV9ZZ/ImONEOsdNyHH0N6yBSe3RAP/6O
dx60bDICKwYFwSGnaa9iGDmOYAlUKTZet2nCAYK8iwvRNNM5IkTr2lX8V+w9unTx
/ClwiIRWRJPWTgjAZNdil98qMXCO+ekevvWGBngpK0kTdhNsTWeAEjzpRHp0e7Rs
aCcFAji5AvWiDF6T6BvnW9yKlRK9xBwHnGn7uZvS0Wmd6PEUE3GgoARuaGfZxvE1
gWL57hidpJbK8V6g901dax1s+MStf2wf2ily47SWiy9mXnBV1s19mMSJmo3H+xtj
AtqTnyaWcRVoiUjMYq6qb83KtTpQW4WLJ4q3567hVn2drGzL7bijJzCsUhywT9OY
MmSmsgW9rqBzjribvIBLQ/5l6tnBtM+yYIQ9NPn5CXsZlrVaKhQzxJaUXC5wZ7HJ
nyPLTVD0km11+vmY/sIhtmJ3yXe3dHBAmvys0K+A3UkHLKbCFqfcbKnS+AuHezRm
tdVJsUk08G8Ql6APk1jHi58KJfEQ2W3/5bxuWh9nC+qiHq6JLG0aWHDpNJucBziJ
4hk/adDguY2ykpJ1MlcFztCcF0/65JmI45eBbkNsblIfvg1yzvnwMwsDGJyKwoyW
eWTfCnzmOS1Fxjj7v61HwqusXLa6Q7GjOnzLwMGGZxrWmzUz0TfjsoBrlPFMasNR
mADVe/SE8AD4lH6+TjK2uMAvAxP2fvYSZF1ieqMq3xcaU0V0SL6QFML7UqBWZW98
dlfac6VWohqhF/VELdZKEareHH+DVu4GSQmHxwmQg3K1GExxlkMLdkUQGFCup5Sw
QFJ+VJbOD+0FBBvosYgsYM8IGFDT3VBxqSPMTKHdYZnscJX7qfrb8CC4t7IFwgmW
ui3R85o+E4f2vSLj/VeAeD5vFFB2NnsYHN4R9fwmsVUw6835QYH3kGO6P6867xdc
d81IA6/+gKMBiyuyQThlr1KmWu9+8ii1WRLG61+QFhU5mNrvRzhLnN0p5rYjf4Br
v3CvGg7STZ3erEgcoRQQPcMTQOkBoBKe9SZhW5lW/9CUNjxiur2+KbpU2ncbWAw2
0d4BTG+xusDreydZPCbVKnZdPVqXpd55ONpd5+uWIucOcI/2URcogD05IHqr2V0d
R4fS3L03DRyKHSCs99exRjVzV3jO/qlyWyy+7VTDutme+urrFpDE5frvrIRXkACE
4aIN1VQ3D5K4MOKBuwDgVWlRcb7uezWyjUaG6qIw1H8sXwJbW2AHrOuK2n3t1X6H
vfHe2e6KnehL6qCMaiesXVnm3gg0y3mFIkUOopN/iOt4edKu7/McYLRWpLYSMtDa
i62Eu6NbVgzCkSjf8oEZ/jPsYIDb2iFVZCsiUXIKK0n5dtMDT1d/6nWInA5SQ7fz
QMYhY18O6dixtAErdqPAzWwZNp0dQs6rKwgxKBi5N24V6xBgjYCmb8VQxzpMwaeK
vhHP5Rx+qGJabW20PdT2ZwAdoMBa1onBzIXNRusN9rjagHTborvdIvMvXWKm8K+Z
b0UrbhDX1a9REMDtGalZzZ9UKQY0OrMXSWe1nUMSfn5GCRTeHdiMd9dBB8b7dzr6
ccs/STZPt4wCa43n4hxTtCTgm0joRn4fSCh+zkrrYQP9//i3v2Kld7eCfSdun8b1
8VQlmX9IcBoHQl9sTk3bAX4s5342mHFBumHUlVYb16DguVjFxEa5strV9ESbSjYe
q3VzFrimETpQItaIzB/ubnjJ3j6Cjnplb8F8FF1Coa2aIXxtn2PSceeKKX9iruIR
xjmfKWf2pX0WKvi0YBR5hb0CgeMvAQ40ycGce6KBz19Ps34sXSMrEPEIfsiHtUde
9Cqe6UBhT+Dg2kEdMBnXSjsGxmpAS/jL+uI48LiED3QlHBNDiDxJWETmAsyjcPxz
Mfp8t/dFTt/GUPkdJqiSLucsFNpNX5A7AgYZRWpkB1C4igdvtj4Vhjb3FQTR0id7
8R8XYTMvQCCyNo9lxKQXGUo5ae/aSpEPEfdrLv5fSSOmhHlMi9DicIEco/ttPTrH
yx2vpz4MP9Z7FoVDlJxGuYIpnsPQPbIY7Cnb+9RHWQyW7JeYOstM3L0EKDWnw8z8
9kBBNUSfHRGQ2DjHZsAcLYGHEbGmzvL8FtrjIUnVSnwV6TQqaqoTNfnF7Q3cTte4
P0D41Nfo2vCEj9jiKuduV0+nbL2Ju6YZYEtidfoBlyxttoVMaecwZht8aWrqzQii
nI2rC7aLM7ev8axLZajN7N7Zn8RV6rtArZ5u64npervJtu07vQxR9MsCTDFV8XGA
3QnKMWnsn2d9ec+Lr6vC5ydkZyltWtGfYNVHH8jDjEgAmHGTTwV4cHdPlP9Z+myR
z89+W7/sWZ1blUN8akwVZZDeY4sjZNnq1sF2p3/F+hJO0nhaGIRGsbIZCLHG69sM
vG3aYH+hgaWTdIUOnUqYY6jGwASHyhYtAkOPeL0UJIqGgFUxrFXolJ9vBmIpkqld
zKnEtrLlFwwqs+ilKdAxH5FrxSAkUiGAL6DQpFwmW5SeLnAdUcLzRPrzQZvAwBqx
Gl+xD1Qajyr1TTUOZYaPXa23au3JsWDiVnsnF/YSRILabrfgdDwegxMKFvnw0eFD
uliO9WrFllZaAT9Rb0fqzcu3PPRILyu3PrhaSOj8hilZaNX4hrv/5Q7UdAUXNTw8
ckcvh/IgKxAHBdffLYzgjA3ouU4qFdNCavAk9KLF2aHe/ATkAVM538FNPJMqM+v5
3+fQKGQ/A+9rDAbOHgnvzyCL/JXr5RsYzKRzJ61loW8QVI0a+NdaUdWDvIIdgMu3
rQR2uRlcjdpCfEnfHTS5VDjQ6tgf9b1hB1t16a7RIup5L7/v+4X/MVzNA1mEs9TY
BSAoLlTIJ+RwOCUQW1ZTYymwA1RjgyaOy3ARe/CAHG9Cf2YDb66CQXPa7ofuvT6K
WcMnsRKJAKAD2SildHMwGjassl8bsxc1bnyTnQ/WVHjL9QsfGqrIBX5cs7QAy6RN
pMXddMseB6AyuDTC8evf9w618TBPR8Z8qredhxwP8L9sR1dGgD3zccBPdBhl0YHs
pMIKFDzy6og9Wu5yW9/y4Vor6+sOQiaWE8x0utq6lBmu2oT7PI7hU+OWbmMhRuJP
aGt9R1sa1NUFqQ9+LJDqOfZnKqnAskPbQmoSK7I3KIG0Zhyy6K3X1Ie6xBkvucWg
/hkqpq6f+ugsXgA52pfTsGaRy10zyU8fB6s6B+u+uUSgJN30rSRIRlTnaPmjPJnx
GSas9J5wjSLApofRLSDn0l83AoKiPH7fU8ImuaYVuOmAcDr/gq5zhcOh92o0jbN9
ZqC20rP9r/K2a/T3FoW84tKc298QoiCk0aRstLKGfRtT0Mag9GNQ8vMYHqQOb9eT
7mTEsstk9KY5m10ybsAIvIh/t6Ds1Jclrctjzwzc3NhFogKGKRm+4SBI+BHi468Q
Ftz/JRC3fgTp6gCAreXdmXkMEnxr6cg2dG20v2wufOzeZwAdfkQPhO5MX11lHjdy
y8oOGycHkiOynHlblytT3NaLUjILP8qanyaqrAsDbtA7fgB8YXI6p7cn++BH9LCO
DpxQ/XDkunHjMbJUjFbgHcN5wGFKgfNqdTOAZyjHgxHrTxk1lSR/RVcSeBMrHoRd
e3GnbMRjN8UPAS3wok8rtJfF/mFsLpz5/JU+/X7uWzbNvKlv2dNgcGpzABfT1gzj
EH63jtAe43k3uvxFy/kFnGY80F48l9ruw/HGq0vaLtpdcyTgzXOLpuae5oZU1buo
GzTClzdcSmGK5gDoTnKPWceclxFwgAMW+ToYf4qw5LrE0fXnujPvVHeQ1sTqg78B
iOGeB9nQntc4iXC8xdH/oWTVLGudQIfiTY0UNAhQLDofHXShBTNiqJLZ9O25Avpc
W5bb/6/jqKkcYkTKmbHqdc3s9ggf8xt60Krbsvkfev7fmH23hRbk5mH+qZ93Ozfr
/JT7GYFmD+LkJuW+VXL7p8xDoTUG5x0N57rjXNVm3lcd+SeQyeYMOIb77/MJiH4L
fyxcj5iYGX/OCTP56IxNtSRZhDrdo2DDc82iSBQNT+ue6TIv9fVsiApw/qusHXPb
Wlb5QeRbFRa8u/17B3QSuwoQVpA6IxTHexmMyULZ5gEH4BT4q3g2XD+wIy1RWQzR
PM2kmOdt5cLAVp6jF/5H6eY0qclMEvZspYHlqadWaIOKdnVkc4Mbn9eAW3iPnW6C
gu+hXds5MxVpBO8tXh4WWovNsvByAlJnodBqn3QfTUGluvApqhyIytW+Bb4HRq1P
FuoCTpEj+gg3sb8bDa1In4swBroDeELvoVuLxxwr+02VijjFy6iVhf+sqEO0szgw
Zbmg1BQ6Yv98M+WziPg6nEnUDqXTLhysNF2to/LM19o6fX2ECDTg52xG42Atuue+
ChsgWxbJrzFzy0Nj1esMGBGmtk6OvcgaAbL8h3gixZf9o7LROYIxZ/wlJBigpAdv
ByzF1QiBerlDxZt4F3xXeho6ikObTCW3/3Htntq3Hen9TIEIj3l/1PpsrsppRE9I
bJ5Mc80OgX/ZWnTBLmGPlGbrnBnyR0l5CcCLIllUp9LGPJ1gCB5H+yvX8vLxIb9b
lI1+IU7Ya/yjuWdb0oI3+naJb2JLxun37+9xRg3poReZakCiQKbx7IN4cCKQl/Jc
o+8y//FfS57tR9rmb2zjoiBk+yJ/C6xAQfA+WlSw8TBAOYZdxjZmbK+kP92YokYv
5+eWvJdcD4SmLTDvRyR5Ws2eVIdba43QqRB+eWf+Pst04V/iVWTPfOSkvroJjQhq
i6d/jffhlOdOPyLSPbsUznuEcraurQixS6FeKbKapXTHBSWNjau5bDsoMx/BsYiF
CpB7jrhfJk+5HxW8OdKAvL7pcEeavVZnUWryekrdUEfh8zbajoVCTZkJkGdjuOkd
ao4FstW0UKSue8QHvSRG9YSGtBnHKxkMdGGbUBTdqFhgmQUYoG1g3hDxWwOd2Oik
PtPjY4S5sfPN8HwzrBYE28qkIWBBxmBV7bG1n3ND62ptbxKODhG9nLPXI7HmjB6U
8Vo20qYg3Hi+2TPHUD/MH22wyDWzQO0/s3OQh78UVAorUKDoTgHnYpvwYWhV86MV
1AS0EGNTydjwvQa6IR9CdhemaN6Lud1B0zPMPHx8uIIS5aIpLkqj6JOautPvtMJZ
eG7wtd3ycLmBPA1KAdxnlPXrXxjm1pQnDkhOX6VFBCsYww90ruWb2okCsQXm/4Ru
xgEceJmfY+dtfQKRL6bTYf5y84OqsOv77dYIdfjFCElAuIGGAdchu/z0yo61buys
wT4QskZQShL9Dln1Vgn4YA+XVK33q8b/EM74sl3DSvXkN2XLrrPmiiozGpKw7/CI
Jz8NTmhYVWjDzIY3/YcFp+0fmneetwFrnUWyLHlw25AzsENAoiCam4XX9YbfkRIa
Kz0GkGDVifLiljNS+QAwnTM+BxEzVEwBpKKTc6JAY4trYzrx4XjW/D2+b6+raq5h
53k8s0FIXf21LS8kKPG4GmXFDEM7aCSgFY8UoU0EMNfMs4TLmsUshOsS9D9KgTdI
GhaIFhso6WyMRKj6R3pRLzZF0Heot5uqI5tI+AAn4fXuUdzHrLhsYUk8Bs2JvA7/
SdJUXxZeXTWUfIx1tu6NseFACV1Kk+NBYezAHy1HbyMAjaPMD+yk8Mk3GfQX1Fp6
8eWom/YI75yMr5LZcyBvrABDuXd7oZna+QwABuLYLuAWZzy6pu46v+K+ES2Xud8H
A8oLjKMcGGwajn0GAF5c8HJqSdjoq5iGHjEt+VKVbxyCnCPzAj9m7O+22muhyiAS
4/HXsYHrUrU7CyxRDILjglXLXeAZlbNmFEv6I1tVomMuFZrHDlo6wFJ0b0udYqIV
zFXJZ2gDG18Zbq2w7Fc6LV+5sypi7JuBrixQKEXRsMbldbb+Wu59Vw0IFu2pkMtc
rZynuviR2C8ovJpG0oX0S9niCmpj7ITW1RX9SAGpXGh62GuAJYjlIA1uAR/hwBVk
LC85BQSMEzyoicGQIkAKYUFIrAJXJXc2jqdirL6UbCMIaQf3/kfxSVOtNdAmHWhz
TDhbULUvTdj27yKzzkLf5uhxKIXe4/CLOyClPxV722sY2KWvyGD5TJ+1K4G4uBF1
lWzZL1598DL9+fvhN1AZVLhFmDRwwXW1AyBrLB8oLDa87s9OejFagx6N6VnIFCrL
F9tI+FG0dLuC+L6OXaW4iiZwyCyPemcQwSESI97GQU9zuk56q42C7YIPGmdqhqdF
1FzIHMbn4eVujJI9na9qfmuhNZ0Uu0VlJEiMRattL4S3DkxDmas05Jk3q/ImQA3G
s8RioMBk+rDrEa/0BUgWOWP0f4085K5qLbYPyWLC1pI6jI1Yxwh9u+uYDxEAeRMT
mgdFuOnkWEPKO0jKw1oMcJoGDD9tXiL/r0KPswQjzeHrngCJc1mNQvPeN9jaQckV
fGlhh9rv2l0zaB8qI8Cz+nkcjaaMhXhADqN4vFZGKG9PEQf9mmGFqXhp+vvACPc3
MTyTA4WVKMI9srfDu+5sgvqm//MoJ2sXo/ymLfdAqaMgCknnsOyPCHhD74yN1PKH
584+JttsKpqH4m9drTpjWJYQt9w+iibNrwhNJiXqgnmSUnYm3de6eFT6QpUNwdhx
Mo9lVFliX6LVi8TrmGWwiPaWfbB5uKbxWqjTKrKkvbmR5hofiYTZEESUMgH7ISFF
kkvTQfyDXZ8IdI/QbaosS0DGasiUVYfywpG1B7sbPlXdQTA/IvSbATHnuR4AFPpS
JXhYyOgoFMq+jLRiLydz1m65U5HmtfEJRrpn94qdUja6aL7qgzV5vdsWsIgu2AF+
Zlqtzd7vNJ7WEUWtkx7WBb7zDKyqVL/u94LHvV0tE0ettsJK39F17dK17AZ2cAeg
e5j5lvFErrFHwPFDYpVgKt7c12DbnynElSAWMJIzleQeVTWqu3ChXtzuk2r5/Ff9
dWJwvl+/gcFyHDbw88GkWfYxUAKmqpc6K9onfElEjnYTk0ghuKAfMSoca50nFGLd
vAIQFp6Pbyqu8kloLUylVY/37JF2pZXUNnoJQRFjPKSOPZMOgcYzHiRT6UJy/GaS
ukHFXQx2F/103yPSAyV0ymHCvOna1O3D2g/+DDYgOrihSFrjjw5tHoV8PhWy/cU4
65clggTRWnyE4AoF4yVI4iv/wHJL6pQSfFuZp+XvCzTTu1Dre7bGSGhMjC7dmdyp
rXMxNZApqeDCIcaJP1khpTi1OIFOUf36sTOpwjS8OGkg5VLy2rIIc9dKEVKUWlIJ
bkTVKm11o02IpgU7J4sSb/trGBlqElFF6a+AZdVwi5MiJMpSi3YBcYrqYNxJWCRK
VBAVNtZ0vZ3bd1LC9OJXSkNhsaFrpVJx5uZ1kjvUiOPJss7rS8gFItRzMjXwwBD2
y3W24jDqnXUZgdgO1x5ZNIGUYG/3+U3nvgvpYdC8YoEYv5oTwZVykyDMT0IFnvuL
GOLM1zbYVojEz6Dx+SCHI3zoVSj7W+3z/CZiHxi7l/hbiWOcJKb37CH4+XaopP2w
GF2AgJbQahAOZlP7uqZAk9ciay2xZ7cRLBcvrzV+sjwyqQKGvXAlcNFZ3rDmvpXf
xr2z5Ym7gFrt3+2jRh1i45YXLiuItKvgCoqebiOcChbiEQGMxL94k8n7H7adk7m9
aI3HQP+V1xUebL2XO8ixN6rj4jegyQ3jAoeTcJL+cmrYWlEh7pCxZfsmaCYt/TXo
j69HiPpGcIuO9wdwt0WgLLhToOhDhaz6q74s5EJdoP8GABk21RvXGCtYx9CI9d/y
rASVymn52ryvCVcmaZhzXxA9Y4SB6eGwWTk7fmPr1jjq7liFvWy/0qAAWFcEGSWi
aws4TzmCiGIvuwxyrQeTKBndfgS0lLT5rp6G5Z59BiacJ1EMVfspXl+9dAJwNHSH
wsug/vMTIlN8o/N278EIOPxugOIdVrAo1SJ4BQtVFNeCOkPZuUqvUq7DSNEc06n8
Dba3UZPGBhQ3MXe687DYF9jp9iNuPQy495kfjWD4vVEX+wjZNQX4ptY24BYygUX6
GxAD87vTzmZNeNDdJSLE3DwhDknzKrxkVj9/DZAT0Ab8lVA/yRv8lt/Ofd9sOsTn
nTxJj5In3s0rH17+ZMkgC2uflieN9vkAG69FnYinWiOZFW//u/5hHpxXQnwLdvXK
18k2WAu9cf64tp3W3dSCgVl/SXuxrgWIhOVXDZ7061gCVOaMaq2MEEVurkDBK7GY
ArNm+jdQc+pP1FBTFktngGgSo1xptyZU1QiBo49kwIi0+tcq4pqYQNidZ9My0CBy
DQPBPojZll4nS/7AUfkD65pgasVVxaN5dRyBU5EgKiBiKpPwHged8GrrzNr3BdmT
9ql8Q+3GZ7dyVlBFhdT2/wKg/iV2QJj1K3HyQf05213+VxypAodgp8PoxONbKF8P
0FHjJ7j4FEw457VwCC+I2To1gFRqQhzcqIEpDDVD4UO/6MMUtkThnVxuOajLBX2k
etPkMU6ZeJ5yBlmDsNI5e09YDUSgaF/GhCTBdmo9QBlkbgVaqIRh1DUU7XluKo1e
1WJD3BWB8i27q5KX2sMmsTw6aPeRAoSUhBfzU/D1tHOqAALjb/s8sLE1mZ6TKROW
ZniTSo78UVn2KDeHQv5Pf3bsWNzw0KIb8tDDIgtwys797+9KtpPrWDtQIup4e28t
deSpSjircjySIxTw1SQFkzECUIfG/7k/HsaE+6u2H17nbBPYtfbiYvZiphrARMh5
kJ8V5oi2pkeLsoyGumrr21qi4oPU0WnindJZ6/OTm0+Vx8NDqs8QiQBc4w/R2pG9
pf/8CwEw4wLw7yBE09TJIV2r3ubx5HWXYMoghpabMl+ZqNOtRxmjPNfQbq99HF1V
nKHZHcNoJIiN4Rom0ldL2cEfOQHyLNyIBfBC66WhD0/LnasWPh8VnrWFU3zaRbaF
vHUnyXKYif9c7fTa6zfANIdVTMYJp4BQOGNIS+9yL3BVYHArXdOy+SdrIxUlZC2l
6C4u1BHAZlxQHc47IfWSV+vMXogwzvFGS9tyhGfLYgW6DG3UDyFkJKpLOYBzNpjM
Yt5R8vG5dYmKg67WVe2vMsGlKAHqatZAKMHApO15I8o51gho2KUmLB6q21nRsAZM
poh9QhfE+bKoZfnOqsnnQpsTFnfFQ4xUfVF2Bej5BNoxCJkIo0LuGz0Q9KOamqUJ
kfn6Az6+GjeWTnp5VeVFltpH4bu7AxIPKtmnj1tRJCk/BH4meoXQzCwBF0A9Mkac
Bf9+FDlbWYovJKoqT+oURa2kff7nMfpqe0mWg/LzXWijuNDASMqSXlW/9aoDJGm7
uZ8XaFYRjoeHues7US0StVOz4BvZzQN2p6BY46XiullFf6RYtlXygpxJm3j68XO1
6xKw+iXjlTRsawEagBQFlFpR4SGlDaGQ2SFnCf5DEh6HnMd/fM4o6JlmkTkScbGA
H3nHXEIv73uzA5tIInzGoswWsjnQMaP4EwFw1Xc/hsYHDHhzirDZf4o9oZhoN4pt
WW7WUGi0cJboW9FGeKmojgkj1ZZkNVXUVF3twzZ8PmXHFboZtKA+MNnCk3s5fBzT
i/EDWkFkdH1ciithh/Zq0vRp6EYHepBdmTDbKXwexhxeQwmZxASBsaAM/5iRaBa9
5E4ADgal/QVOOapjrPx9Y2auWY5gbEI3DpMuX23kynXv78YxWFIUZzybZ5syj6ho
N/uORTZY6j2st3+Wt9e+BzpyIkr4utKdGgBQILDw/RCjtAYXJmD1kxIajMAhlasv
bAGIpydLKwi44wfkgOJkDMBv+Nidx2xcLm233lrGOOnJ7IlbHrgeW+ujS26cEUoU
Rh4ptS83ipyoRCiqEujjIGmqi+bnwwentxaBqt0YrsJ9TB5NpLBC13gPhjNW6X7A
rM7VNWDvsQhwWGImgoGhb15gHTgCj9P9s/pzUuYGeEvp3XZtnsgExuOXTF5H2jl7
Z1/JV0h0ZhY+Tc4LZ0LLa1lSMOBdJ4mcqfBpissQz5FUYw9fy5A5Vbah5AscNHjN
90egUAqTj9DJU69bdAtHMhtTLMA84jQppSy18l51SA4MmYaBuFTw57qk2ckdcLdz
TugMybM1ElGKuROpDbBMZSEVVZAX8GWGoe08DvXEBKVbn3NR2QtHpgcPnU3hunDO
/9fOyFjf7cMydNMtyRA16hXGFBLAzbvW9IoSXlcH0vRjBsRymnYvr/RFibyQ7/Qt
fOJnM2HXsPluG5FV1XNjT8UMRJ9NvGeiX12xoxIuHGn8IrvRbuX3QRoImX2Y5hbc
It1HDijJQjJOnAU0SrDjnZDUAad6t57xzqrRtWUHHkiIPhy5sWSCtxwBqt2RkDnB
/PZ2A41B+qvmw/xlFxAVDQx5GlzgoaoaG/hYp+xcFsGMUR5SV02NY8makMDdu3Fk
areEwx6sppRt/6wZQaoU+m7P2+9XZud9mlR6j6rTtkjD3y1878OqYOf640tRRyO1
nPXpQF+8+Hxwi4fuFxDlOFk7k8C2t3mIs7pq4EP5D0MuD607rVqbixaqlzZOTdiQ
/MJjVSIqT7VQxgvuOHp+v3MKNHVZ1dAlhWxKBkVG1alfe+ztHKoLz4iU5yDJgFvc
ezR0+Snw+xFsx/3JuOSSKEXlJ2YRtiokdQEtzb1HRElGQMB9M/WhwNLRVe8LYvQ7
Lh5qiVhPTyl0201lQwFllITfQvgM0Gd+z+FQPS/0s2VLA8X38UUX2PHW8WwI0C29
gHid82aLjWXbfdZwu8J4DA2fXaU5eqWw9UOxtsKrOdfZxuG2F0r6uOSZVrCMPWWW
tzETqqSTLHWtBHgtf88MCrpxv5Mp9/EwwB/ayjHUzyAtrld4tbwNzHaalbC9lAqX
XTjtaj7tdFPLm+51NUQc3uY0GbOUg+JotwDZsDYZK7Cb/DdN+vkBnjVX0Q87rbo2
63ObZeEafln1jboXzNYPxMDUZph4dNsnz/CzyQJJm6/8VYsecV3mrQbfD2dm99IW
8w56c1KWPQOpg++L8tLU51q/0OAiCSQlBGEDFnQH534NOA4ig2/ujRBxZCR0Z7BQ
SPfLcbz4akYUDnSfe5Z5aKCf2R3ZSTqomphI8c/rXNFui1ukz0bhefMCff7nrG16
nGMcPkoCxJFD08/nhlD6rv1dOvStPuCDdVZf9F0b/fi/zEkxW6zlelepyd5J7R2b
zMTEZhinVaihf7iwlkGLa2Oq4zUyEAHLJmoBgrSdhUhqGiuERkn/1adCIG7W6H02
k3VovcZ9OkpzSgGDdPyrTdJBES01qYkVTQ0COm/2s3d+dO4PdZiEQG31L/O6Ky6Q
WxzgSONfErUwZ7vdlzaR/Yi6O0Y3eCGXkOJtUCb9cdiexjv7OR7oEMvkeT1Wm5gK
DML8SEne+DrmIbzAHGW9HMeHPYbJm5K/t3hwVY7n4dgP1aXmNxtsnbXyaKsWZyWJ
Kk+OOSQ7/DJD7aNNXS4ehbw1k2AybihtZ9PBYWMBiQCOcAQ7iKq+3kIDVhpQ72KA
ojtjVD4w5z3t4ZwAVpGLLzuUZfKsmQ43AZkF6tpfU2qUzp/WKZ8ztTbnET/duz2Z
WNpBfXTcgfgYhrPAvYuxyqQfJaA+6NWayqpxCZW1cF/DPIZNZeU1cnFElz5LM8+c
JB39HDXFVeduucx2XtNKBJz4ADGcx9MhR5F1mxWFf9+yUxlzGeZnwlTEIwkz4UEC
8CYd7uICh9TARFOEwsoEB0W6E+bL2r5i7eMXL3MDekpNOuuhtaijTXr3cg8HNkgm
D9QbkOHC9BkSOV3s7eGmv89eTAHEeNNHDc75zFmrhUkKh6xov4x+1GPXCSItqi5T
bVL3XGHsngWiyAnJX3+oNVp0pFY8SyC4ioSkW9cVNahotmVF3V++x8MapCV0OOfj
65YGVfJ5uQiTkrTcsLVZ6fEE1PhsryzkH5FKSi3KSIYLQJg8o45cMYvzJmyCfj1V
jrDVLZgqzZsJNpoMolOXlMqXGeap8WzXafLMY0KEmEsbVgoIkeBDirqODc24KdEy
IfdBnRoHI0AlZ/t3nqDaWUx6n91zxxowQZQiGdWWx1f5r5hN3A+PqNWzorjSiUCu
Th7GI+i8zauhEJz+2WeGA2V31cR8nRkYVZuxU35HuIINXPevRBSK+ByC61DyybNa
Q90MR6BhxFVr3UESWjSsXuogj4UTWs8FoxkDePQNSNLRASrauq5yKx9z8lO3sTAt
1cgfEJ+9o473nswmuT+P4zppXR315+znT1g5706o2fc+p8KezcOfbjrOt6nBY1OP
vgHOgLOTme3oImIP1W5PliBYcyQ8TdDCJshRxl/hnQUfhCng3S/gXRhoMZELwD5O
UEsG2Y9ZI0jaA8QBFMrTKGkcfA4XmNHlNwFr360Wg9kMJy5QmTFDU2kIzKW9Db8c
AuniX3ao8F4/uwteiDS4v5lOkddlVuuNVs837zguVUkzlfuFCC7Iuon/xVyuu8PM
7eN0WysspDCC2XguzrfO2YZgDQSXyyJTvpy+HZILxHHDD2pwOEKR55SfYJOUt4Ht
r3XP4WfwV85PvtXoCWzhyRGAoHyamQ17MhZqVrjciAuub/s/BX5Lx9yAhkmIy/A9
ydgO/L+7ox2rSKV2WBtGNx17pufpn9EG1Kr7h0atwHiRb/FbpK+dR1WCmGVo7HZQ
cwpqYy8+CQh6e1KlXBm9rsV+teJDrJo2VqNeINcaFbaxpXo9cjiMT58Seyr54rb9
iqNpHZ8mIo+9NaHjA5t8PmBcYpQNthlebjh0xfBjXAWk6s/Jp0+nC/onDL1E6orj
tz1ecXYL4RRR83QlY5KyXN5wyTibuWJbQ+0olU0w3bMdvnc5vZN9/mYDfZyhiDXk
AY+bFA4bl66MPMMx8H5FdhDe15Ns9Zqq96bWBp6snW4SDJyEpswRWC55ZxucxIwO
QUBINcwfLN3iN1XI3xo2gtm+q1JBDCjLoaR7zmeRpHqEGvodQ+jV+F98r1+JxKXp
vxTOO91pq3fX/7j/VdAruBiIUpfTUQ4cPgddlcs/POBM6MPldkVWceLcU0E8hZlL
MHGv6VR/Y0wNlenplx/CIIDYOzU59W0SStiby4nW0jAD3qBbB8DxOTturyfbl3Nd
N/yLheIpUGPFMXBpSv5ambBotnncTdNcfaDLCj7tDlssetDIaiw89QEGSk4ZhatT
+kSIFKUNvJLP3ENNmULk9+bQXiKwhKIMJiaMRanOfroFTaWwKCBTq0sK+bi2NA+d
CVmY3pgA7Xbz+E/nLWzKFy+BD7Z8cmnfaXVzaTFCkqL7upG3h8ewEgtmxRblhj7T
slnQqaTckp7LlZHnBFrDCtBR51KKxyvqtoX+E5yVuXTkh2LVEtk6KwbvpFmzssrk
bsDprkczjZXCNzP4Qvel+VEcqJmKdwK8XQh9NfvLQNNLeTW+f+VOFk3bR5mtcMSJ
LOTIjHylTz6UDmM8rjPna1oFwjp6hCKFG6TUMKIP4O4c7MXusIvaoZkbLIaqsu3u
umlLG/1jJJQU41sQWtd5J0T60nJQtC9HMr7ZzBLAwySjrc90aWc4VBmJIYG7zoNj
ksLxitRPPs4+GvVDJc1qC+IqyBwOQNDDNS6s9jSMQDMjxSGCV0CrrpJvAIBbemC0
EhUN2OKlwScdxXmBtzkH9sHaMUNFNLdEyUKi2W8g8GodyuCGF/sCsHs7ZfMEH32n
ujWxkT3TOeXnkxuJ7mOr5RVYxHu5TtQQqBUwVdIUTmaxMTcip5YxrGv2noZ+7Lix
vAHJZ2jXgrIwRHgZLbWidmGPigkVj5ZQVhuzqZ3zkNQ7D/WL/ja8x8nU/x8WBZXo
7gymkXnYRUyjHAV8XMD5OxMalhv4Uo7zRaCFjDNokqpoBcvcn2Ya4dzOHDuNhZVn
vuuOsf9N0mR6u3munB3rRT6KFQe9gknb0X4kWiECALd7V14d5zdIUYJ3A/uhiqY/
GereBvelMWnr43T0jLFpXwKcnh93oS+3ZQa5l6udBuaDtAX0cqys5gHnhbOLPqoR
nCsFYIeY5r7AEjtzQMyWW1kHWxamjbDbPvivFqtcPzPq0KPWRL1LrRblBZI6xdHi
QSU59Wo4dbLHoSbrR6o0r5ah2QEZR4Rh0fmEUCmboVTpaPSTjxlF+QkmYRCw81AK
Dpz1Z0gJadStRZ6Qz2fKRd/5zGUEqKAHY4wUofyLKKi2h/JgX0dQ9NfwWoEt1qK/
IdHHtPHX5+HTp1phT5E7coQjVo2oeVigPhEIKoW96g7PSCFZZTVGkKv5BRpDtMoA
MIwDPYcP1QqMCDQVeGYH8+GbY7WqSnZrXB0i3bfVJ7SIyOJFgGfWBPETsxsNPWrL
tdlj+wSwSVm3aF8VeMCTIz93Xm5IhN9yx6VAZV3HmBd6OfslVT8++9rl6pA5nFQK
dGECB3bLDrFdHB09EF6bdgymX6Fd/M1wJ0wHuIYx4ihcaPq+LOfjLV0qO7EBDeSw
rb6KPvL6Tm3UUv5M8xPGuaMaG98GHfA3Q2WFhva4/NSkU6Dt0+5bSfja0M9Ylt3H
ltMgVryM6jzIjji3chkelhAr/nCVfZQpEYT8Y8ICa2nRqQvkORAQnOp50EopgrrD
1IWDk9DQ9kFSiewBJIo9S2hpySjDTHH04mB+Re8js8EW5pmazQEqFEtiUpfRDveW
YLbqTIhvY4JLY2JC33RjxJW5SDIVLMuWGFL3O81w8T83R+iPr1QUqoIVWhl9NzDZ
8H+evqgkt/azTgofZi7TSgmP8a2dpE3GYf4rkr7jksIP3KjKg06KK6Gig1/D7brb
haO3AT35fT32DmZvcDVOJAnXdax9BIVReLGXOQy3EGdlF3D08kPPihUlMd5CCP1H
IAb3Phf4DZfxYy17MsraOqE8NSzggoU+0Nv1TgO/q1TYB/OfPgOH0OZhy/OFI63G
iI+x6rhEsMhtB7lcat/8GHwMR/UU30jOgYLBSNcx8QAxWTvhc7yehu1tUst2RLyX
hqiCxpACR13rIZj4u8ujNzo4cHXYYXT7yOPag7uTzfEjQRQvjxTUB4nal7lTLo6d
YMnMS5Dtb6jr6EcJuAcJnNZwdRFajDBBKXqzYRdiSyZupUbUctuharIx+b96aOah
3sGkfqFbRVBAw7WRyNa0dON1cnvdyO7HwfDQCtDipk2qqnKJMwMK+GE3EorJw8Mt
R4gHWnxqxpt5nQGrAyi/j+pPc2ay6ZybNqiCLzWCh3SjMJkakJhOE+cVLBDplikx
RjM4W8xetcc824RRLWjKj3nqG9j5j771i3eHr16mV16NZnMM74X55aKICht7y4ki
Da5k2WuV2S2k7eTEEkUIZXc4qXc6d4v5w9fHjOL0vCrVIJaX/Zv1B5NQe5r1Pmjk
lzj1SChEXlyqrXLwTADMWJBEiqZq2ZfrIY6fK/Qie0JXPdTFv9w6Rcc4xImWBpFK
liME74RFmtWpkcgkE/MKxvp3El25XAX9B7xr4s7CxilBwG/Pa9NYJFrP40gVVFCa
zbrJK7Dd8sGuOfrj3l0g+Tjjh4CcmHp5A8D9UH97EGnSCtRIAJ8pmOIwFg+q1bhr
hPR9P4jfGHlVpDeWSAUs6mbzWW5sgUrIg+kkr70+t/km5UrjzKm+n9hGGmSxnaov
gJx1hy0NVLGqMLjbYIQaGcZUdkoMzlRSeDXTo/ENfSAC06kx7l+qil9HCidcPnhb
dPaQZjhO5SMYnzTln1tYjmjGw4ObcbBqfBMUozX0MKoDF2/0JcBkLVQokQdI5Taz
qc0g44xMC/XccPTKuRvRFScsqhx8AZwvr604C3A78BH7t4HLD2sMUXF1jzB0SijF
Vay9LEdlktsFpLxaCN9fI9VZOEbyEVlYvzhGDCep9s/Ott5IPPdpGVeF9Zxu1SAs
l8KsbZyONWeNlIqxPY//jZ8cJXqDQrHWGo+r2sl56u22ff8SobjBMjXoCtdO7vz6
78Iw1hBVYn4qmTcckwBSLyd8CPoLMA8iO99wGENF5/vdUxJXnAe+Em/5mvYq5J5d
rob+pefs24uC5loN+j6y1FTDAQRafqeeSP/xjOwseEHzWBwoZV8ntpwbSRvHy3UC
axuSdCIByL9P9BBCy00iPt2SWMpB3SodRoPw0T5llFiOQ3DSGMbECjosVCqV/CAn
S/UyCk27DHZvlLrh7f3Exc4dKxc8ZwuKLtIF0qws+csTBK3ZbbrRbZsyzLEVq9e9
7OznpjVP4SRMmnPFHtjRBSJHV5UCyUDuKdRmh0aDZ7Lvwj2HGcH26lAb1ChZbIwU
EA59C4Yj3MgI5b9cMW3FWnxL4pq9ClghLxq+meLXFd6hg3OaudeSI29hlhx2rG5d
s56+M1Q90jmy4xm/6WpALASkoZgXt//tUYdKBb2RkTpI985qP1eHqT4r55008eUd
bpTkWy2QkOKU7n95DpTw7TAewG/KQfFiyEr6F53PqXL8B79UbkgaHOtb3XZfDXop
Ussv63WzPIbL8HLQGYHuUvQnE4eH6eowxTh9nBBAmilDjlzdtgJvw+uEC3nCif/U
qDmIrdcISxB7ad46JlZ8QFBANvpuixHJHbTBpWads0omrHl3K+PK1RyUUj9mQsfR
lDPbVn3hn+7aiQ36hfT8sbEPKSUHzRgUC/3+eN7u3CUQAIDCwAcOtLUSdpfpQixC
XlubklMLuieR3o04i8zxgjojv23K3vdSiYi6oDlRkGQ9f2x2JNltjs0Rbvwhx5vV
oGfQi5yejikE5mvBREaBV2uc3KEYMnko1JjD5g/8ULZWdqSlDdp2jPFCsGw51CKK
qox+sFDSONFp3zDnHU8qMvbkU3J8SByDVwBCfhAUo+IkauZhUxoYxCXNZPfUoHXz
r0AtcPe/BfpsYmuDV5ifnITDRWPbvINGG9/dg8rI6c9RcITlKlVMu9tV+h4CrieH
PM3nPYbd0P6uQKLAc0zp6ra/aP9OI0+mDAJwlF6bAwt5Z9hcys5//fr5mMZhnYx/
X51/V/B82AfykujP7mPdckdLxx9p7iXjNuZUezz+/P4RkdVHWshg1by50cvQXUK+
fRWMQFDFePUImGDT1Wsp7RUbYEA5HidXv3oMzdQ4C5eGTUcFHBt+t2VntRpLfSGk
GL+o3DYOyUkq388v13+1zUrUx0Q5F4bPC2f6d2TOjpM5gIFDACKNnXwHRZvmyAEd
CuPb+TuLkrIq7b7L69KYtEEvS5XkFHGd1keDHAny0jk+aYmosfHKQ5ulG9wHcjV6
AED/0NAt5w6QQ9I7eqyr4T1NNzkt7s8n9ro4WAkaJQftKKujkPYwSPT+BGJozvcw
Bnrnqta6/m8P1UhdYxHI7RdG0Yirf3lS65NTTdj2SSo9JfdiTJ/2jlWqX1EbUY+4
oXPZXzMi5Hu/94iYzMWgXF4ywmw6YFLx8gM4I00dMp8j/xJSiFJ+e4ri+wTv5Ufh
HE0F/UMFUQrQRdwNtazjsEyA0FFSmE1e6wGmMXDGzjgnDqmKWTcSP00XRZrIkhbd
fngKYdnpX/94Jt/8zBkUxLqoewnFeOo3XD6K4xNShrltw5iQKHS+QnWqKU5+vHtW
YjezKh50l8qyz00ipoCa4Tm5xIfC/vcLaEkertWO3/70zK5RBpNud7gZE4shbGXh
77PwZmHQzswYEeb5eS2qjx+vSXtqa2USqVFkeGZeFznVgE1sDOFr7qrZyNQFU4I1
lOr0rwof41MeG7KAKfhtN9DDbjootuqMt/Ek1i6eTN0UiTawL4F0DbKQAeG56/t7
wUhPvVpHeEOMihnOBZmRfnSbWZZezK6+4PK5RKLKelpH8xvomzWueD7ht93QLsv/
LH9GafsaQD3N6o5eXkNXwqbA0Qf1Qm1hXxLbcocLNbbDjSXF3f2O+cnUU3WUR1m9
kluCsw+oyO+SVA2CJb8iki1akzRar01hrrA7UcugmrBG0n0MIHGOV686jJe71rmM
P7fbJqiGZfETsnBfa51UV3Xtw4VW64+w6krSU8JqVIAMc/himkAQLGvzGvZV3/6E
0YHUg6mXoMA5Xe/Nuu6yQupXsbh+282e0jhY9nbFPi3XxsG7sw7dfXYmYmlFxyW7
Gnp/o+mFyA+GwSvkuGCG+TS50a2Rtyx6gUYcAmC1ak9+YqeXt81h4p738ESdN4i3
4m6sCSD5JbR5X3BHaXLUfQernJcCOjrNSJeX1OG4FIJkuIuMJ3AqjmXvAwLS5ixT
X7cj0D88/Kh1WK/LhKUctmbk3s64gsgZ6Bdk5uW1UlNpZHazx3XOuBP51bvkFXvE
Lqf7P118EBw7vxy7K/wHIrdyzXV2ZRn/2SnRLfQ0epKIyeFjoLeHDM/E/t7XX94r
aYeU8flts6JpYJbC6+BtisjNEv5gUF+1HWGsXi8SW31lnl3nTG7J0GJjdmdPyGge
rvNR6Y11SEgwlam+ZGzTWIsCqj9jlfiNT2nHzV5zq8s5veVYt9iVwflPVFq0Grez
W4aa6E15kJCOZxXQ6NwoyTUizu8ivrd8SjoIrjyGSaG7IKoBtxj4gnfR9laQUidI
jYfNksJu22qMhicJpo8KjhSfrhkoQoAwZx+exVO1hLIp0daMbDvnDQNVr/hDENqm
W3JDa0gVLONvsPS2WoNc9mIsXcJ61rFKW+BwSgJ0EZlHPzGMAnUd50m4VIf/erl9
Kgde1b9VZq9qzW+TQtYeaQRWTf9O/uEWD+qNQtpJexq2KKJ79Pw/yQfKgrxmxpX0
/ZOjA9nq7+kdbCi0TFZQJsx1EeOhyexH30yHDWI1FRVUH+FKvFP9aWAvqQqfqH5q
27zcFpg1OsdqH4+1zFnsCiY2LRU/SGa2A8z36N9MacZ8tfjhuLWW38KgchdcifBJ
+7pNB+3nR4kyoiHgxYOdF61IXVZsBnrTPr9jJF/FSIyJeMTEgg20XHENv8rs3XTm
odw3g5njIvyBBEFAe3devwn0HrHgbQ4NHRhgnhFUvGVdU/C7jEsDb+W8YH03i/fk
34lYf2LolKScP3YX3QEjte4xhyGcc2ow8MNMN6ddLto5YHDHkbtqr+9jr3Q+uexI
nbzjPQr6KHJnYj9Uu0Dl9+YSfOwAl6mqD7kNge8cFmykURqiPB368FQB8OSit195
JnVo/Dbv1IGlqU91PtdWJ7HPeovQF1Ej4hYatwGH41KL/73DjhVMJyKLpNAvlIa/
bK98S46XDj/7NgmFPOXcMzvFjKDj1OqW1joZEGLKpQe6lqyPyUmsVOA0E1WrZRce
/AUkhi7lXOue+dojAu9S6Rbjxzn8ueXEyrq7HP/Qh96Na4AA1GkOr1fHImmQhCXF
8StTKeGcZNTtm1CqdQkK2OEN9yBVvwtWFzjWn1K/PH4DBE/w+j3EDD5adm3TAukW
+w9f3RbRgc05Tduxilk987kLQsVn1+UkSSMsDST6v9MokJ3COL2M+6MeEiKNG5oY
5VgykG/bIOULXYzWaIu9PhIZxr6/iM7JqAH+uPfyRnGCIsuusB3RZSiJmfnVCGve
pLcauKRZ1WCA+vMn/PlcrnnKw03dLu9YwnaGSXxDWcuKCKlreAKQFOBeiC58oX25
vGjZ+SnGvTh2clodh9adT6/iFG8V0VOkPaeuqPMLsI5OOgPWPJ/otvCqgIsnUHjT
OsQiD82FJpfwPskRskSnSwbDb6xSUfGaeSQ/3s6r/x9OuOyLZymV/cO4IY9nmvON
3wvidA08biFqNyCnrxXyUKqJZ0p+rmr2YFtdNoK+JD8a2c3vOXNwJLsvkxMdM12h
3XatUUhF0gATDgaHC4GUv5ihZ3nxRGUez+oJXJ0NyyR2agzbTHQNg9ILg8wkOJDM
VaVvTdrP3jTNP/zD/dyabgLUVaVjN50dGFwjPfdB6p9s3GHgvs+lX4nScNVS9DmY
4mABgkV1WfUEcJxW9HVtfT9lSfMLlJ+6YB5vM1HBQQGUJWfXaKDYhpEdBY+YNRdR
jBr286Qi0DnSVEiyk4h/YdfmRAHWNablsG1wC3b3Y1zXb0erJUg3T2p8yGws966C
dFeWU13ywwANF+syT1eg8CrdUD/+yw2KAOEMZYWm6ds5nvAMQhPmDdFnRLqtSure
5vkA/Vea/bVvhEfnqeAzkmvi7NHxhA99qFB1bQ2fly9fpHPc7jJUpO6D0P+N0rGV
GLjxAoYJYIThAtqq0VlNR73qnR/LZVWBcTCYjuY/YJqhzkmuItCqDmkn+sSFFwEz
n86nZo7VfnkiQ8NBS79u2fj5UbCoDVyl6KolyfgoeKcUzYeWQ5qDZbcc/k9bcAPj
q6nXrd0FkQ1v0U4fNgSKjSRUKEPJs5Vllu1eXPgcpwP2af59hZJW2hQlEyiNs/ug
MN19Ec7SRjh1Pxn/ILyFQr5X2MbV1RK5rYm+sGcBkCpdzf+QzO624MVJG7TbgbLf
CSRwROAM+0mK/PbLPESicbZ+TLzkRjU9QY+O03nM8CYgA6/ODcLpuzVk1P4P7ZzZ
iU61Oyr3C0c2EQvaBKbkUXGIK00O5iJWw6u5/rdEhZz/nJXq9HvbGPcLQV66et3H
xkOlGPLgTv54Cd5XmC8dPWvTqx7Qjn4n+p5DxpLQMkCAji57QxZPX1YW7464KPGG
huwycurn1zPjO8oMA8xfBLs+YQ/AZZYdwzt7hr5oRGv6zcK7dKwYIAn2NPCcQp/I
Du1wUrK3qfzMT+O7e7KddTk+tY/p2iG0k/AsSpCIk96B43nUfayonpazkhPe7e/U
sfbdpCRnkALIaNz0QcgHi9pVi4xxlnEld1iK44MmPulp39zgFRqLlTrAsAJCOL/k
ShyifvL4n0QIGSy3CPM1ghCuf0lP2pyOuq4jBJ2pp49yhPDb+0kaMAP3aLWH5s4Q
Sbsd27/VlPOyRbNCaA38yBx+yqzLHTYReFNKVLf2Zkgcs2VeuyYF0lqErh32rjqj
c0YqmewTSuaAVZkEgg1gXbfLVxwappb3Yx5eF+H4YMNyLZ89S3yc6DWZjAvUj1Jo
0oqcWDkiNSM+0A3QMgmJxoi2zHB89UbkMRvAOYx0VmaGSCZ/Yg5AzqyekNFsNHYX
uJVfUZs/MXKNrPwS1MRRW6Kbfw4YhvCrq5x3F1GObEcUH3SjCo2FcslMEUvSdFvm
qFSAxNjWe4CmffC0u7FcZij2CyErXpSFpeQRh1j5S5ovYfZniiAgns2D2wL0t+I4
Zzfjnlu+RGzBBscpNrv6WIh1OjSODa60mYevOheedpkdw7l2nIzyRWtMCfM5DmL9
pF+PkHSZTpQfXP3U7Jl6Q2oRrJjaitcZJau1Sg6tk51cmqzmLzzpPHEs8vsGWy6a
Y1HlyFvBw7xDX+HD5WwjRCD/o5rHPp6Kwm713+/m361mmerfHpMtWtqtfH3yI/0F
NWJ4MBnWxwgVM0jlKGyYc2kg3GowwE9Iopea5iicH3duGmIlecv5KkRu8NZ78XJ2
nXrhfAXDHfkZPjzv5eDZrj4/wAjNX7bO7r2PxKFv2b64jG8jqHqMA4R/JUuhZnBL
j2TmeKgGsaexD1zUyTYCyY07iQbSgl5fG2ms1Yiapdp4dsHmIVMLtDr4A2YDfRVO
QHKMNu/Z14SWjEpei6PMpBbyhLnU2fvfpuT6xPyDbSDum7oEm9ngO60dRbzJ7thp
vpo0ig3vsg+fpKqPKHRrHhIMptzdQ2/wktDZMhsg0xqp8dtUXxBUitzZ5iqcXnnC
bxKIvPMGGVCJMPPzjp8rnAMo5ofJVrDjeqInv2LzNn17ut6Evoyks1kR2tKY6keY
hF4xpuo8cKE2licQZVU86fxpiXsuAQ94DZKQwH5Pux2WnKufSb//DkxHkafqfWyz
iJRqGMg57MOLTAi4J4G1jXjdiDnFQMH4b0Mak6U3kZcjvgSuVC10R92ZATidnVZA
tlE44ocXWspSoag2fINz0zlq8eyQdSFJjlP4kC66sjG4n5YJPrCpxrUsyq6P1HEU
lHTgk3dnSaE3FMZImMFDnUwrDm+xL+JQG6det80RI1PCuuOTW3Z/7yafhFrRDf9J
c7Iz/psZam5xHBSiZM/RQEuZRszi1GRMdnFG0730+VDFwYbFzsEK7wOP6mzu5SLL
weEaGNJ7fkmMxx2QLtBTgKMvM29ZoAAqKmPRfGnjZYSL/+powkzlvdWZBtvAAYBo
UVpF57Ezz8qLF1z5IeO34023AqYUKj0A6ifJntTr+v0vTvokoZdRIFvNLfz9vVVa
/TvW/hryCvz+Q3HuZNQ8ooC9L0XyelZ0KIoyRGn7K16r7XHuqhUlnWiNXlJZC/nY
nIeQ+LqpDk2dEZr+bsyemDHkCOaE9GmHCHBD13bOhk895idSJJgVGf2xvH+PAveM
e5bDSpRrS34yOSeorOo7cLwFeaIQ4G20dQMkCT5nUlokzVInnvo1z6qfjD/CMLnU
xba3/lRJyhum1lkiGo4b4khakg+9kry6hRGft4kRuEQ9ENfqw9VHVdl2r0sgIsEt
gIsvBeakY1mqssU789m+JQzS2dhEYJqnEU+egDJfF1pfmPwMKdG7LoqkQt/4JoFH
zkR5p4wlPyDHMW0F+2isRDzMhFyYaCZsUcfsOO0PECeGKV+8gUnIkfD3Rv+CXoL3
/x401xO/BmjXrMDmP1FgrGjmJMsnIXgqmr16rTn5jhN4VNIDm1BaEipU98bax/tn
WHu/t3zpg9t4C3jx7yeXkaJgL6MzWu82yC6dQJe1vb6aCJJ02hEvWPxS0ux0Ex2O
jgvX8rYm+R6LFopE4aSti/jveV9SricLQ+NbZtxihO1KqCbjjKSGH8Qeo3AcLX2t
KYR183PZ4+ZyhKLi8kcrlDCvulpy53Cq8FECu8K3E3U=

`pragma protect end_protected
