// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oSsPuVRvGqW7k/hn6sKy8XP/P+zsDVodVBK/HUzmdQInJIZILqpS8pqLIcJ0
THnOTEfbDpcZgeZhiqcaAn4/ML4X5fO17fOG+Qmsxu8FiUhnoYrOt5P8W88q
Xef5D6pvOl1+er07jFGWCcTsKv9VWDgg+OHBdC10NtymOUp3QJGkLj4pVhD8
Y88pWfbsqfqHlOgMhJR5jqJ++JBY499yibaADNJmfyx9ozn9Pgdp4YNXN8iK
N4idCEI3GrxAun9CPndh82YgFLcGsNDIDlMAiiWbZA9BPwxY1wa8xVkBXWyP
13Nf7VZFdgd3ygVDduaFD1GCKeCp6J/9MVtcsWA3JQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AZCiouEUI+zFp6EUlRQdjLVRq9XDHOH3wwIWljnEaRXDacZSnU4wu0hjYnmD
tx8RfnseyeXUIBL8gv6apKb6OlMbGg2x7gbPfNuvszHzpcypB1zNE5E2ll50
ZXGFKLAnyBpICQmi2q2Y/G4r1Cp3f1jsefgMNUZ5cUr5jUQ6CXiHmTd2y9YZ
9RAsPxUEuKsa5PwhU+FHMnvQ0zFvFX47d3+YhMr0mAwZPg5pvw/cWTKAaUX3
0SqZjKc0V5Vd6V8xZu4TgK+uY3XW5TrAxhEPO14jBCDuu9dKHQTxIt051n7X
lUlsr1rRn5SIKw/RrN1JaFFA3EODIuqcszrpR0b/bQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QKEOf/1Jw7xig8cCvKii8ZfJbiKhCqL1i5/g1bfVDmAE9QTOOJ4JezIoLsXM
LuzPcdkmmgdSzCjuFehmI821qFD5eL07Ej4qUMr4tA0XeRv96mCRcGKWeUVW
2vYs3ITuTq/7UTsYOrN5G6/yVyUosvv/SWF/2uLqQE5o6q1pwkiFlcU8WZpb
fNCkkanJtknzgMQK1mQz51YeDzRgfxXnGGwyFwHrHkGcW39cGzZcTmtt7b9l
NRDLJ2oiz78U9XIHIs/7bpSQFpuWZwFTtRIpfL2sLv+BNe9uhNYNHNiIwAgM
GEb5bwtxMy4FZIUIjw20UbBcTamG+Zcwfs/a8ve0vQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DnkOuaHm+aNs0gxj+1tvtLkcPy4OD2sy8NH2fOCu7x7DRt9TVUfdGhfoc/eX
m/2XF1Ob9/t+5nElKqTsRqYYwwqqrR6dhpqTsvEZ9tHkvF6t7scuDkqjdQkM
tS+g4FLpYxsrx+zOeS+dOU94okmh3qW3/3NZ1hXZ9cpxuJ2FJgU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mhrpvdtBo9JujHnGF6zRRW/iQW2smTG2zd4YLmRA67wUqkgjkzulA382eB1J
SN2EdRsaGxSdXh7wKmOZe6t1Ep16IoiSIEanCKN51/Lzmp8CRRNW1zun9zHc
Ye+7wjRcpQVjOuCYJGnrzglxOqhZ0H/IrnY11Tubv80tUiAbHHqPWjSH+LzL
WZbi4xM41uiKvBglDMfoIR0dz9LcMgVm22uthITWfJVvhHw4n5qeqFwgCgJs
MIpLzA5sYM4z7hbVCoZSxMZoszdsg9hI5tsYz8jjh1LoPEolGE1zh+roQbhu
K0/JOQWhhAvD3m8/gLVwU5RV9YXkgrm0RQumXo1d01vk+kI1jCAIKsPa1rwa
V9YDtTvF94OTmoACiNQ5ihtuqwW0+2Ys5UuvaFiHSNGEF+L1MaqbRXSfcaKF
7bN7xyzAq0hTHQKcR00A65WtrocA9WYSIZR/XIJLKQK8cooox7uRYsTwE/Be
62Vs2A65mwuG4dTzWtN8A1XT7vTMwXEu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G9f9q/XXnWet6mviW09H/bxDUGHcl0FYA/YddN7hjLGTE374uJLMvnzT7IIj
MpZDBLeu0IM+raYgUbxmB1eyrLyT2mO7qUjVhB6ocbQD9CBjR+8EB4P5GMvP
rHsLGAS5MQ2c07liCAApE4X5qyFt6OTyjVjPx5niHUw4leXDNV8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hwimnlOO+SazjuxMV58zoFg0HBRo/5S/9tU1vEPOG1wxVfl7RDlh8gYRUIIH
aWOt1eHLbHwdWPc+mHxpXDq4iO7fDNVFkFvgBqAPJnWq3T/N2rLSPiOcpZ2t
lyg2g5TinluuAiLw1z6Fw5pqIgWWmgMNE4UIwBVU3ZwG+pR6rJM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1360)
`pragma protect data_block
xdC4mB/SEqwN/qGVkEPB2jUaG/0abw+kPPFwhtS62Jia8B8ONVUYsAyIfSDM
obnKhwnoaRj3Y00kPmjSm3jPWe5JOUonajj8rgNfgDnNTWuyRTTotzFHIL7t
nqub02m5pGnkZ5ymxkvfz5ME8mBwQYSSqbPLm7/OJhH3oJ8mb6jzt+SLnnP8
PY+7/YjgM9+FNHOCzVNrdUyXO7Z8RMOiKiJA/o6zIQewyOskyJhZawtGUtGJ
SCXFamE0YTyAMLYqAKrlI9R5EhG1240jpvZcyGUAbYcmOkR5813YBP+FXvRp
TSwpk2ax2yjmRdc9Ag6NNUjDktSgCSkcZpzFJrByWdA0dZn2N+Ok4sXGHJe6
L9W48PfMJi3PaQU75xl9MgDS8N3laH2kt77JCXJgiqXS3yRhi27rtXoxRyzm
+qLd39QFY14Zk4ixccIY3Vqwc5hOSFBQ3NWF48ErHpDQephV7KKEzJIBQr6l
iyAkh7DWdUJ5KU/NHdaEqBgIxWwQgY5/K+s9MIPtnGSCi/KWXWcSrfGaoM0t
9EvzquN6xZIrBG4pMjQOVkHaSGVDIXxSoyrDuDGi87sq5pLFvBYwFHqS3CVH
3Xjq85X3RX0rm1wQFfo1YAg75Qodso9My000qJfFdV0zMICfqu5Pk2jJtHGr
vQkPH9oU6QlekVFmw/XGHieXukhL5vabXeJmHDKOp5RWFaErshRLlQW/ENjn
GlvJpdJ+47fiYJ7WXqMiYJI8dOiYj5YYwDNpLppeJbSdsqWIRr3Z7AurAN2K
1xxsj/7k9Ot2dR6eazKqODBMPu4lgH3vGhCZH/qlUohnsWDH3arkl9owG3H7
B8CMR4I34z8dl0DZAvd2FkWBh+0oDMS3Y8q4fZvBqccFdxmvtnGejbu3ZAGr
d/gjh45V6r8Isix3KkZRem7VBtsczsJC+hrX0LZ0DWJiNAHp+9Ry5oTYF+yj
0Im74EFXeEHS/T9kdox21bGZbpYBMRjcYSCeK4ubEamz85bgVihEIonihjHI
HMwrJ+TOWYR2yNFu2H3N2lVx6E68NCpptXpiZ7eRsYyVgRsEbj3yKoED2NZf
gcMdUB1oM/O2tyndOyaEawo1arWXHDbNWAz/i5HGw0W1PdFs1tx+sP7AYZUd
MT0W4wDliUg8PJKVi1jKx8E9SS9ts6UNP3HTFfErgyjji/VHJ/td7rOh7bGT
dvXesFWyyqdgrgSIIrYO17q6qM7FXhFXxnbogsO2a9PAdPmHtCUs475hi8/+
z1gOOwUAn+92iUpOekmxUV6JpNhRyNuwzouR4Lmme/wfRcwuo2gohP4rM6aC
ixJp+vzRXw/vejiU0qy6r5fMAyhV9rEuIJuaudg2cjYW9b+Hbvs0kT/gwykT
cQH6i3vG+PdtQ0yW9gOsppTbk//5vWTr11uP+4NtxS024PXcRNaJXY9YsDGZ
4tfV63tr5jH7tox2I0Cr8tjl6KDcOYu86bCin2/MFEZlkYbZ9bLq2n+avvBd
Umwu66pB3zAps6qBwzK1LVMfbBH9RVmLT0X8JRXuM4K2d/38O+46nC+sn2ss
imn6Yy9YJbvWMbgf0P4iBAGThUClFatHwRpJ/fqvQTJpD5eJXufh8meumMo2
c4TqaJ8LN/T0yOhXliswoks5lpc/oy8rOvzT+T1AWJ/06xL7kxj9m0jU/gB4
iTkK5OxmJCzT8gTtejWXxFBSN4zk/ddfXrItMtnPQ0glxeK5TBZEfjOea0vm
0uG+zr4pIx6m0oQsfKqar+dzEvd2fXbsLoWcR36+gKrQyNpuc5x0Pi3GeXKM
HcopkYhvP36NBA==

`pragma protect end_protected
