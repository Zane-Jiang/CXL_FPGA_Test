// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bh7yTih8SbRBznoJql4H1rUkUivaAPRh6WBaW6fle1x8BdGPE0sPRa3VmIFf
9ObHVsbdYv7f8araEJ/+ekbmJZHFxA9b74Vxv5N117KGNjkutP4CmLPb48IY
zVKjOta2Sja+nlNPZa2/nxJ+RYLZs9Jq8Q4LgV9Cl4sj1dGW0/ViM174VQbD
Ti7Ui8GOAcQdpVaKTh/7MFsmrRYe1CIB6KIiMBzhDlMmhNK0N0YheKIhGRzd
d/AK4+xgpXTPKwNzOeloonczu5Z6wh4sfUE6+hJaXPcucJjyIwaohWtTTp5g
Y0O/kQKditrDXD+Jykaeq38LXHaU6DKhl+nEYrHfwA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YoyInsv3mjyvwDNk8yQH3BFvY4evEf7Wna0QYImBEUM+r1RmVIFNCqJyqQZc
hHhurreXyH6Ff5om5+OO8/whGdhg7gIMWXhGNKaDXhgb48HCKMxhG3Fld9XN
6elOmz/bxEgghidPdy1j5tTjC65zUWctrn37V/Tyb3KckNhmNXzVvcsorJJY
YT86k15q9VByePrW1D57zBUQ/i1DBHe2xvX+Yr/4RIckdpQBq13AY2QhUg9C
JO1IJHovb8uCZlEmvCYKaTl8DAM4sdk0ZdTwxollgoSTlm4P8aFBVoslHukN
GKpDQt2TBj7qBWuNJzrVjM4SF45C9pFMpTncGbR+Qw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ce7DaR76zBcB0tzEajnwarXjxfKga/I28S0CkjMzT77mK/ij7t3+hV0MiZyc
vn+GEtqm+Zy8F0q4pDH36qz2balTOEs6LPMo7/RuLZGHyJZUinJl9jq92Y+u
nplgMGz8Zwh7fpYIB3oV/r371xOMi/BzZs/x6VCEtFWsUCztbMNxa/Xmw6jD
WZeNCR/MsvETk45yg+BE9fI4q5QXtJckS0lpyRuuHIA/3sQLpIMrKeV16e6W
bdsVA89HjF/ATwuVzskb3kbSPx3fkw0ejtXADOG5n4Pf93dh8MUYHBPBf+cE
dVTzp6Cgu0C58lWnged1NEc374wcAOZCpgijPSuwXw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JytgS7BjmwQQMlk6jFbunnSBKTdc/HX1/pDpJYvXzLcKK31kKLMpN+jFkoUW
SJ2RzNvDeg94oXtJb34Ovy0CZaiCkEgtaiUvQTXpL8irQAi05DnWEKROozVl
OMF5XDchOtPSEKFr91qtpFVcCfo/Rq9wijDvZP0xdRWsGiNaEgg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jyo0Tr+qq0kBshTwr4RFuO9jRHL+4z65YAXTCamnt9EX3jYUBg/WnfGLn30a
Zn0YScQQRMlJLGOYQnSnmWrNjDVGPGOq/LFuhDTXtLRY9w9soRWa6hjJ/fEP
kb6GTnQIo5p2GJX+TI3MQ3ZhqbkxEzpTCH4jCiDa4Mjqp86Q1BRmVN3D2lbe
G8zb/7NjXLMARczu35bvkUnb0B3AKes5bgg4XymmWuWnsOAZAt/P8P35tfpV
G/WdXl5R387yZhbbOUQsv+jMx4XMQ0c1fmC2Y9TZivVZ2c6++RvhhhQEzxDT
/mGDPskNy11x2JzFwJw/PEZXZrKl2x7u/6K5FU2aK0P8xK6v8vWYj/E3aS8w
P6OtCDNBJFWG8bw4v5ZMJGWSsthn29gzYTcCBHc1O0/Q7po8vdcPNgJbOxGa
4zo0P13RnfY0SkzLxFarkN0En4mUamfoC1t8KR/hjjHpgY4GLr9iF4mR8tcz
lIK08sHeiiWQpqESezENPkIRVghN5oN7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bBOxRyIHL216ODMTNkBY0s3nJyioEN1O8SEnOIHLey5V+xKSmp00pC1+deNN
8b3GFWkXYG//oFWkgF09mXq8EYiqhHG7Qop8tOhpfckowGHKvE06/YK0lith
3Y8bwhyZe03D2uGWwtsY7rSykVqT5DSByNdcv/8dMeJ9dfbvZeg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e/zZIpiJfpVxXnuxcxM5MpS9j6lv5YjONIWG1t0iIrAznLCM+hM2agCWX0MT
XPqPLiWl0Y3k1TovbYrMB0ydAZROYozPjjGbApQ4IAjEPSwydHwSheRJ4bWg
SS9jyz1SWWLt4yJv7CWG77ou/oVF6BbEX2xopSLSZ+647YXIjPc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14160)
`pragma protect data_block
MS4DOLT/SicIe8zdcizOqOQuooljPSWqmuPa4DGDDRGFMc7yfiSlRyC8hYeY
QtPI2chdZzypyHEjtMzHpxVHKc5ovWWOiTucZ3dui+fwH8W08qntRvNpCX85
kjl2yEEssCMjaxhGmRuRkYjdQ+Six35T7Wm5O00EjBOMJhVpdG20cjsNAGF1
1sdzpSjaxaY0lWLwK6cvYeGHiMjOTiu73srfsY5FHvtz8QoqabzQxGmQDxr9
Mv4ATOkzkjPQ2POH/TmUXL2CUzxB9pSowqCJjcW0bB629ZPxAksldX/Z+t3h
ipBqBHYvFqJkuEDpNvbei3hfGFWTBKMyXImrKGFjXITiGsIidTgfdu+r0+01
tAnpHg3kXw/pzKLcfIlVlsEmYwNSrzGM23onM8HR0GZ0J1FUMuIuMfJGb52Z
N4hZuR6GRKvDooaby14yA9+zpB8KobsWZzbmPyNAy0aOVqGSo057YwA4O0d3
t+Z0gym3cO8/OPPlTU8Chy5fa1hX9KwJQNMZbIoY4OIWaU+DEjBM4q/7Q320
5GTNLe7QhYXhmeFpZ4OaCeTjfSOwG1aiZlvVnzlB/nwHvslcdzgENTZghVt0
yUV6EAvOVetsHTKiy/XVKOMMojMmio6Ljd+enn0x6H8rFvgkg+g+Q9r1W3nB
2rFP43E5DfiStvOYkdRmv8HjyVt3fAYwGyb50aIxS1CwFa08UTWpqFnk8sbO
mNWtOicluQbKrYy+c0+eUMuhS+eRgAwt92uegPW9XGiKDiHKrqxCss0D9GaF
q54PK/8Sh6mFH+dYPCOavLiAly9pr/5VNJXHzYzllEZ0f8XdxwN39V5Fdn8R
nAY51CPYkPFFTfSNiGfx31C83OmdQgGlusgBaA94S3idHcivOuGHzbankU7l
suOjYMqZZ3aLwPTVMcAL5ZzlC6muDbuwKjH3/kjytaaOmqg4I6SbuNlWrX2d
ILxnsljyv8ofn7BN9hi/UkykMej8z/JWHnujMJyHQgbWGakNYtutIhIu/coR
NZR7MIt//L6Rfmtsvp2RtGK7DBPyYsUnmi5nuh3vtn1c1/L4sv6qc3uq/YGS
Louqtph322I8TpbmoiQOiifSzl92LaP98X6PNS5ojDncFjurTPi88qkKAKJg
MWgrrP12mG3+3ubdsUOz3wDAss+1AAWEBjCzg+AYsP69PoY2wQTHtdnPla4a
x5KJ0pYpVsKQ80umKJQcPMoQPx2ndW+hr/wz6WOIyp0Tr5F4M4S+HtKuKMWq
3b/CaMrY2vXigCdINmqVjLElQIrFAIEm3R24GdoXR0VymCCv7Xf66gbvUdH1
riq129ol82+mHP+dBsz5Hn7K02YH9Zxby6TXdsL00XDGvjAWD9BjVhAsJfot
cZgZilriMUlOKx1qArPKLXLHDYWyGa5ZzM+zz6hlUkyJ/CcLOkmJCAllpa+T
W5MUksjk2ZxXiPzgJEx3H+e86w5N8zvB9CZoQ5G2L2xMMFfHEU0dLROY0L0a
Ns/IidhI/k7fjpMt9hAruHttej4ITU6nCFIrowCJ/6CfXp+0veRmsUvAVIIS
jRvNEM8Nz0K4hKj9rzmt+wa23Txf1CLo7lDEaRPRS6TYYMS07ymaQOyoB7+X
FRsqqWG5obKjwIT9HGMvpB8b0BruTVy4TNlk9+4Zp58lX8wE7YcQFPWf4kYx
RyItND+MTl4M93j+O6YsUPrPGFOWmMHj4Zv08HNXcTmGBtHoPPZpDDJoj49+
lj7UNaXsKmG4afrFlAeIuySgcJkrb3GawaXyqpOx37JzwtxHxx8Kw0ntO+fH
zgiTbXpeNQQ0b594GZdTItXUAPCqjzG2JiN8t84W6aWpLaLe/RHetFQeKxZX
gkV53ZTRKAdujAGW42jQhk/ahmmuXY0rfT9Tpx3ddBMDLZqCfJjz7S9nVNKW
oMFHvni/wH9ph5v/zrgtWjTU7Qc6w1aQ6DIbZXBj43yvtvBJBrwWgezLhwGF
cuG89pGUv3Tm+ZnmARO7gOXTfjul5FMFYXl77sEW5cF0krPivlVrgan4XnWW
9PQsj0Xlm0/D2jX3K+TDmwvnAnafBzgnjIZDcfk9fU2BI2ZzxT0mNZxB2F+8
RH0UZ1wl+wugGGd7m9/4bj0a7tBaLNHbkS8YcwI42NPeVjLT7BAqLuGYfms7
AM0WWw7wPL8D6NUWE64f7ZHNE49jSG5cgNQKyfu+EDGqKAAJ5OOU/cT05DKy
oStuWtstGoKxpZnxy49S0R/fYP4k5fHcksyjYnoPKUJP3zBIELLnQnUuZxoR
O/lQD1Q/lB46YJVURn0CEKbyNVgtMVNG+4hkL8fNLPNzaZoBK95B/7VwVcel
o3G3LHpyy/yUGZyM5qp1LiW3hOHWmpx1VX//Xi7bJ4WtH1TIVDQWMhS70Q9z
H1+4467Fo5voBIdpOcJf0vN7kQHh2dMMfqxg7/Q1f++HmLvzEeqvzMuf98EI
UGxSFmIFHfu31fCvzXcoQyjzVw+zeLJEWqWKxS5gQ8ljdgayeXLey/0EGp8c
8oIbgW5Wd1Mlsjs8YIWaOPX6BierSGICbF0+JHfiPs2lS9FVXTvlt4iPuTY5
t3ki34W/o6AUmV5gz2ZGdajRMaxhaLavxCTVhdDktGLY6ub7rD1T2wvhxPQy
OMlILoNDvURCuihS3hPziG7qBiixMFDsTYRjlTca9z+sdlMdlfFR2tq5wdHZ
5MOUOItiS3D3GzI9C39RcCiLYSvhvYNpW19rDxqsLkCA7/ABBC9cNHzpFfpv
3lzLUEDSbYl9s7quhPYJ5pGRw+XcTNzigCAqskVDrVYnuEpYDmoZH780+Cng
NTkmds1I1VgOB5LVKSxoZzJTVWSV1YsiTjosEJB4+n7v/ZicrP08XZ+H4AgG
FfnbhrCzw6PL2QOsyau8wM6GFfkvmhpgkjiPuFqwF6ArJakePGy1ByzcqeGN
Z5tFUZSgbIFUscbr52JPmjBpMlXXgxDmlfLuu+PBRtxYAYjjJINAmv91B+P3
/tZJlIsk/X0Huzk2tj1z5+42qxMOhzz+lYT3GmBh1u2ce6OcPTs2w5wnT742
m7Dzi8eTWmFynDp1E25a+/GRvkrK+55wSOIumYffMSSi2Vv13CxbFn1Pgyp0
Tvhg3SgnI0/2CEr97TvPIK4JuQxfrjlpxw20iljGrsytGBJTXe7a1kTLcLU9
1ZtuQpNHYtnR9l2pzHxPs3W2f7//DIOCUgUk/5LhtrPYCnqthZfJthz3fu85
qmDM/GeMA75KGUnslhYfWeD9iDhq217WWWmk2GUltav/seN85a8/7e4MEJek
ALQkty1pqEO2uQxm35LnbRQ1ZiSICsLscQYab5JokKEej5LFjLwuLxO9Hmo/
HkB/7cjchNR7UBduH6c+sLAOzswtE8I55QahdAga4Ye5q9ju+cftNu44o7yp
rRLb6YH5c2CZyJjGbU57PpEEsOLDfJLFnbaDxbFNaIBR2wJL7Kq5YJyaUtel
/1p7ve3/MOjQ1YTO8lsNc4tjV584U8AZ0xVhz4fmXcRHYN1ZcJK2I2GTJXVg
OgQeVYal+9PHi+skltIxN7LvtSk2m+s7itlVydj4XUu2uNIGhNQqpj/9KqZg
1+VaURVyYIOC4nqWov3H3pyqhxMroydPn/v+/qKoPgJ/7Au1DwptAdYDBtT6
MsqUbchRlXBnWbTcIUD7ofk1uMr19WDnh4Cna+8U8OzzVOZs/Ulb+Fo7sb0b
qjMbgrR2UapU7hXwXaDxWIEAmBXrL30h+fN6xG6vfbBom+bfefGceZX7prL4
UwX77A1BQUlgFMIHSzHV1FXURjSIavbsuZ5Oz3wvdiBrgwFGv8tjTFXMlZLs
HeyET8UUA694oKbXFpRAptiv2oI0GLyXC3vhGQYuI0N9/9aajpCC3yScJsq+
tVKf+q3Ft9l5/mhW3iBLcLyVAZcZibW/VX4vFai8CDcfdk0eiTXXJ6e+nObj
L7NfvF8Uo6pv8eobxSoOLqZkxbCLcSHzNt8TNluHQLWV5ngk8rXaGwnFcplk
NhlBFYdDHz7f+xDxPspMc5ebsa+4/r+2dlxpDqtGnskyPlQh0vb/gaX8COC8
4/62TDpSQa1JVZTwCwpZOGMx7H1T2vs57IW9NZ0EOyKPL1lJimTSI4loNnYj
eVYnYJjjbDJx9WHZ9gZUKjFLTxicgUzVntuzgKl2M5rqKte0sKc3SNRSM89p
btm+LqLpJu1ltO7X/NB5V6Lpqg7q0Xzp5IxplngV1iqOq7e2OFy4/blsD7Do
/yOR5Mv9IMjqM6KFUUWTFLzmWxSuy1D/xERX/4YEzpQLBbViWhXfqa9CDVuh
3ZuKaVSf2CcuyaBldTpEIxSj+obgpw6OIOAY1iGIiZhTY3ojrBnT63G0f0sX
Y0M6h9tnOCb/oyayFHIfPjnv63WiR8anY9rw0jnkV+2QCjXsCGYKUkwfj98h
CDV5OgkiauqRbschrIUDR1w5HWRs9gcwURRmvZrRSrxW6f9Q0VEmuoNvcpZy
pJZavXzpRrhERukBqMKcBsYRWp4jUlXTTcLHLWi+MoWqh7J+wSJwM6f7MZzH
iTaiWb5ptJrABAWYjvXRU2rr+AdFAndY6LQoZhAdJOYHEZvYw8Cm2h9L6Y/Z
6awmKJDaJrn7MaxyT/cZMN8CaZ/oepXB1BDqvr/eSSec+5z3Cc5tkG/5DCvC
D4QHqtUR59LZNgTAy6LzMNa59dPlpy4r+gP/k9jGf2jMM1ANYFk2VobMvpxB
U80B45+VgoNvCyPSJxIKB6f0CfdSkpIPtCUmASiLN6FuPH0fNrEAOD4lHWqf
uPWMIBTEuv6LRspmobUKYM9GaPKrEJ9vc5pOIZyhaxALAANpcipHlX5zbObF
o56IvKQd70PxIUwxa5igQBBOuwugRhauNdnkx0l5KlTi3106KFM3Fq28UZOo
G8qkChB5frV8YnZGiNE1JjYyNBdgniSLtBcpjEQPSH48eQzYUM+9bwzdGZ5h
JBFJpON8lpFsSuBYNV0mkZHHcnmmF935ZtNKAKzlD/LJlPFhLVMs9VSXAGaj
RLTLJtJu447xX/bk1QVauk2q8fHcr1P9AUkMnOnWnxGxrEyHt4LfGs+RbJwX
SeTe10Q6AO8B/tgT5eO3rBgx54EUEi702uYV10sjkndXkxfNaV2xeewYxb31
WRGtQRonx02XfLj0cN9/dzd4ROu2tIGrxr2/V7A8etMwDx4nzoek+eWmFeOs
I9ENAA5RN1uCYBBeqezArYcoe+luguGAr3SbfszTZA9zD/mzV/1MiBSuyMlc
VMW7w7KuVL64zoALDlHfa1v45XBBBLbIsMBQvUYBsxtTnptNh8E3+N00MTHW
0RGACDevEzhpt87nw3Cn0XaP22gOPXt9093Me2jxloCHdYw0klfjRlWMYQVQ
KUoh2uvITZ8shOEqfqRiQAZLEKXfoML5DeKIjIuxunteX4Wv/RW/fB3dK/gG
rRerBTjJdtj23VslXqVH14g1JOLrB9zW6GrC9BTdyvFfg8QaJSfoH9Ufgp+B
nkE1P5uEkUaNTQXgHPty8QYZ5vk/4kwAmzCYIm4DFdjlcyArgx3PTRC/MFmU
96Nq22z6lyql4US8oG2eq109C9EEOYTLyTc+b2u9GGJDIFDi7rE7Q72UIIHj
TWV6EflDiJcdI1sTIeKBt8K0vkGTL0T2lzWTgF0YTfEH+kh9ccv+sk9VQ611
7z5UInyBlDPlPoBTBc8/3YUiXnbsBQHgNGU/TM8esrTzrky84Ox2rRO2WBpf
tj3Sz/tb0Vob+NOacaYj5KTdH85YQhIeVJ8WQmtyR5da5p3hyxjzLmqr0HC7
lXBp8/AZwbblj3pWJTitbHm1KsWKFgEjU5G5wptxkSV8sKotWtLKSOQQPuJJ
f0gtRsxiRkd+zbGqjudyS1I0WA/NFlbBYkxrRCQcNdui0a3c/j/PWGXpjRiP
Y3WTXzRAwgh7vwojZGFOv6ZfoIZuMYfQYrzqPTfoVMQkRPpoGdZ+VREgB1XG
lJSL8dmKEyUUbVAeMfSHWw0/b/7gD8E4igDbC1ZIbQC4itwQuzVk8fWnRWyl
cvohobMf8wV9SKQIgKrHSJIxkS+55b0EoN5T9sSUiH/1K8fo3ZMRKkvyCA8e
QG2McUrJZLaCawamyJWW4n6JKD6r7Jgdtt672kMzeHwArZ2yMIV65NQjfiiZ
tA1djQkDGsYPlaGt97iLJiCHisu8O7zZula/7YqUUVrEFQpLvGvHL84exRyD
rRH7jz12DkvF5syfkld2LHcCko0880+WEkORbfnwYr1hk+5iQoUs2+n/hdzM
wdBZITlXOgC+WiF1IdcXKKfQokhGP4IGMX+1GjFTcgFL12YNDzRmHr8Ydh3E
hkjJjf9oNymGidS+di0+0q3cjDJaC1jdTzL6BVq8R3+z417WUncEo04wdISX
Y0y23ocw30HCrRzGJrexolJzhxWdPgjhVt5PqT7CYeUDXmcWaQVmOuNuiNYv
yA+wbUQtc/noga+p+Noj51VKbzawrB7odcmrBA0Bk4BczTu4WG/ZP5wU5S+i
c79gyxIF2PypOk+rr0uwPOJ0AX3Fwm8A41aTZ+cBz9duaztckeVvS7+8RvBP
8VOhsh8cN1JyGFiDA/bwhpU7lGnX/NW1DNkBJzUvzm58LfYOXL00hCHEKMaY
ocTBwS8aA/CZjsad4NaXHaqOtK0aq67UjRK4jvQF09eDwf6Z8iBh/QUGie8q
RZc9a1k53idXIsMtQJmo5v/Hbc3tJiaUrtkog9fMNQJHzXIxEd4DMruxhlNW
6AUzofe8BQ+WViA/TxhlUQUsQd5NSPXB1AEbJ9xWxdMWfodic33nXJL24udg
k2WfPWairW/kSdsMAw5X7KVKPoIsDZxA9EsPouZpuZf5IMgfhcxPUZWMi1dm
aLM8E1hFm9AViPhdIMVYatxp86CbelKJoDrq8Ozxhz0YnFQxssx8ey1jsWzz
O09gROJcqsl5IzF/9d/qHSpt99Hxk+/ClhsJ107t0Z8cApmybhuA1fBIaKuz
ibm9jB5rmuH+EDXgdL20acPXDa4NtCbvJtoWG/ef58Beef0z0ShlH+iRhL0S
RGO5VMJV3jQZI5WPiRu0k/vP9QkSCmNHOjWaoj3YPqD04YySz0Aap8p6iEBj
u8LDwSs+BWRRJVCdUzFINJOCk7IRmMsxl7ACcsYaN96RJOD1UetAGKzaem8D
Rqpo2HZtwC+TnFKHZ2OHk8HQhZO46jm+l7lKju3b1MKXUbBfktgYdYqkJ54q
36kkY9gYBNf/WEsmw9uo7WB1Yh9/9oy0O65cLOYjP1FQ4RDZ+DkxMz2+V8hV
S5nqBM1HC8RlBExnOTnXDoy0f+LLGqE/0M5EDjDYv4vq2scLLChja6KsQ/8G
X3JdNTusbqGd9pAvToAn8HA03MfSxroERSnBW3/BRvLHX1G6p824xixponDU
K4yNClk5cAy/4AnyN4Hc4/4Ur1R0gK65olYnfbbB3N2wsMUgtcdRgU/nXAEl
dBayMKXenrJv97ypt1QARieLzS52z0OP8J4S3zimaO1eJSYyWFzHrBCuIHjq
qnR6RgWxXnVY9CNt0jRxGqrz+F7NEX4ERyOSnOMfz9oSOyKSHXLlYKYIFOlV
74bmfpX69tsgq13a73pXxkUMXGEdQPspPWpStGw5M3I4yfeE5A0LKQskAbNa
jBGZ51V1DhI10HBdgY0aITFjb+iJstjL2n2Y7zLMTYV8nFzWBKFyFC6Hm8FZ
/QU0zFK8aEwOFC5gKIJke/5QP0j4i6jqrJTE6jQNaM/XoItHuIF/ky2INgXy
q45FpAVMjZsovrHEW5t9DzRsSWmQvVfABJdxx7j+oAb+O5NkfZcZsQ+3IAuP
cTu6cQTof3n/dj93mjRG1kvZZr/Pxd+q1eVvoZWxxbVQGHVLKzBu4vgjng6F
keiiTsg4gMizGRuURdhetQOrMK8SGwjUnpRSKXG+VREMR5aObVI9nbRiUR90
V7TfcY7oIVkZ5fMxtHPMU91v+QHTjuMxaMNcjA8AxgTHeOXwGUr+OlArmGwh
j401ZEs1LUfUO37OVe2B3NdMHZHMpyuHPxdtP2AKMo2fsZJ0HaB2qlhxuRIi
+6YjG1ESanyiawiHpyTR/0tc9AzC5lpjHqERNXWbPGtbk0Dhw2/9Is5tQDx0
nDxRCeb5lPytYeccAJpf9VpkZl3kyKrWUqAQmHNELUHC2L2OZMIDNv5c6kc0
qVkWl/gKJ8NFPXP6fAKtzFQcX6KdbA/zKNbZo9idMuvmeFG91SFhKu87vP21
1qvWWhYoJ+anA+KjdO+LuqzEsYo26K0/jzTXbOfHtAbRb6l0Ffwrn++FkwSH
/Cebk1ktBzUL6UwilnpmyjMGoqXnStk2AarKba6CP/UlMMOn339pC/3L4iNw
o/cYYmL0XapGRy2OS/C8DDcD9u8kWu4ZIJIE+QezwaMAT8oVF6nWjrotNok7
82+xxVPdSTE9yW8+d2xzPLVsraGhq/7f0rbO13K2nXDjCqvPN9w+ZVWz3ysF
xTBAs+8CEnyXeOCfJUDp8yUuyCxg8u662+svtoSaDrxXNCOaATMqmw124xiu
6WP3Icggy2wa1hG9PHhjAgh8N9GEdpHLi4B+govJQTZxA0EZwReY9fUC75hc
k3Hblj4mkaQkLu0XKRvVdmVTmmWKTrS6HQwjIYJXFezkMQp+/AwZcNf6/8d0
LPh5ecLYDKnLyQnBf69q0+33oCV5rqqnWjemCgobhk5KC780Q1bF50QpRTt6
767AiqMouwTFc6p+0dGUR7t6VMRDHFI7eLmxiz0+E3V2Gen6d/EBD8BZuTbw
jOTbgurUKd+dHQuk+MP2ufy4UQvNDC43Dd0Q/Nm3qaJUVbiWpQ8HkOCWavhC
Ke3xOMXn2EO8wrCdi3vohFcbkQY2D1/GXU7kTURy+jjcTUJH9Zblj/nTUNzC
S/MRJSxqOHknlRPH91EJ229BeuzDBoFAlkOQ9pK5LQHtXMNst+vSu+ranLNc
Ulo6JxwDKaxj7xzLAshQA1kMv0eGQFU7ozgEvd8cpi7HNVkeZxADJUKyvHVG
S0QdVlFnw3ai++3myC3YcGf6dnSt/V8iloLJK0GGRIOxTJFHRWrTQSkEygJF
5h3hKMMgmKPefDhODjuRJbjP2wCY3i/eTJmpcb1DQW8VZCBUzPghWX/dCuQM
tkNXb4kiR3IUte4f/TTJiOl5ZDK6L7YTwrGxtC82MWSl/Clvehgp+4fNz+G3
LfmcYrk+jw85MrZO0nRasCDY2KB8al8HUqjnhgL40UW+Kfh2VShclrYr7gbu
Ew29AYr/Q2i4gzzPFxsjOarhFTscLEnXNXP4LesGXJFdEWj2OusOpk3UoM2D
h0/fWGy2dnk4cfU/sGO//INbUhDRwVHK/P6jiVOeMhsmmFBoJ9tFvJalTQSA
nloKMfu4d36J67TmwDB5pCHDG7mcWbl3gX9S14ZYqkKFohlbtMbwR0Rq9DAy
kKJnBa4g4gqfSjyk5U8aaWITWJYA2Z3X14RUZ1rzeX3T5FfKsp5y6eAUNiTQ
BCxfoSTHq5xR7KZu4xeEl9PWh1aGFWCagG75BPCUzPJevHED8TX4VACMTTNU
R/VSumSI9Pu8zgOQB52anD+LrvknlcVEfzTBmyk0tlOkZ50K12TJmQnuZKGg
zyotgPRnKUYT/Nw0uBb7971dNVPyRGJCuYbG0H4bjqfmKNGu0AEdwbvIUWj9
rkpglHJtsl0rhDaLpuVC91Dv6U7yfHDmh6LxLktDuodnzmrDqhZgfdXCrMQ2
xzz2OtnC7f8VnLeZN6FnV+OGm32DMW6n2q2FGv33akz6f1uf/J/FH9eVB3jD
9/+bpHFKv/9mC/1PqrU6tODVbrZK7Jd6Jm9jcLcGi+u58A4exQcHjK1Bnua1
ljqzOT7B5k6IXVlHKgH992bHGU93YVwwImdakTlyNgFnzPGTREELPfRyZDzO
Nu1fWSLmUHKzo5tzBYeffUHKOrrQARLdolnGqI/Qzr0++Mu3nDfFsyXz2YfZ
iWbm/TZaHLV+k+hr7U2VSzKwncyEpXbgRMA09J8I/On3lNNZPI+JtPgjiHSj
URugW837jjKgwyFUixEi4kU/XS4ip7O/d/wJaD/Td9O7Dmk1kMHD+FQsgKwJ
UmwXgM3HDzQGzLil+79PMh+1H5JxxuJWcbT7B5oEXeGf8RWqPdYvIiBDOglr
OubN65eRt32eYSOK7DeZ/VXAONxRAIQpCyWfGP7APrw1qrsR0jPj/f1arv5N
53Kp968gQoWFVObi3/0mX4/+rSZ4ynEoJgDc2ulud4hucTsux+cixhUlIrGY
4FRFcste/mNk7hWCBE3EGt9pfKVlNnk759wbi2+RliJf2OTMIPdgCP4JoIM3
R0bJhiLJPSot/RNjMrvMkIqEebVQfus+kj+6xkvD63Lg7ULzhwdbR/XydaOW
pMbOuS4vdMJMJf5EGuobm5MBf5lTpbkToIsEA4ZPimEabhFG0WX867BjIVx6
9nlWsAZ77HnfAhDqLpLKFTeiYTPTmdLjxg60OqTs3mdPlZoPPTNUACkfKDat
SEMFqmHyQjJ/oOtvAA0ZCQMGdDkTwr5wAnUWvpNqt/aTxSVHFNnz4xvqiZHQ
EGROiHEq/GvbKGlea2wnCiDoPf1YX645dnCA+Hkx9dEAxbtbmBNdvzuGnGO1
pPWytkKzuwlkSw52cjhZeOw/mEYumJHMsKte/yi3u92Sj6SQo4F3cOdEQga9
frpB3QNqZkTUhd4KQZgEambt0G2L+goB1luwBMQutCxG93nC4PFy6nOmibkj
WncN0oxe99WsHo3RRMmiAPk2L5aOb3J75WxzsUh6GqL32zVXX69R3r8h90xa
6CWvwHhdiP78F9WlMhStK6hJbLkJyDQKQ82ULmyL5RQReS/a7r3vf53KaUmC
SrtFVnrMkdHB7lmaZP21s5wp5NQotaZ/VdJmgudVd9+lMjJyfS1BiNj2zLS0
wU9ZyvB49mKgfPzs8E9H2zLezLsb+mJInjuNwHRqKBIVZTaGkwPaBeNye/fG
ks7jpgN0EitPYgyg27aY/8tk/BlmsOmW1ov3NJOyfLER1/cCGTZPthj3lnjw
gQmp/+kgPso0+0C8biWAxGLnwJUZREo8XVNvSsxFH8efiSbSFHv9jiTSmeR4
I9vLEbNsM04l4X91cEQZ17hGkBSaNsdtEz7lC3NcS/vnPskyggpKqD6hKDL9
Minm3WFBkny4Fmye6pPOpljHMFQXrLpLljTejz4fT5vf9VEizagayi/dotj0
BBXhh0cb4uMOjgDQuTTFsIyV+mnNb5Ay4VcmcEJTRZiN4+2SASydKAvxpUIT
VpAgcCJp2/lTEpFp9u/cB9OWbx/BReCRrleL+XK8+bpyt4vijgCnRcUMGyGC
3onk0Y727jpJlQyXILYpK2+ooVeiIytVesgHBj2+eg+z5UzcfAY8XoRtvLPu
Rt2nVVNkB7M/uZQUoM1f3vvRKjH+n4O8e2/CNRmgrgfz9ybLwcNmxJzsu1PY
un6xurkmW/jvifnmUxguKDYYc1egWRHSAsb2Ljl4tW9tVfj5dLHL8A/pHZ2s
H3mMZxT3eGkotvXp313MlvCyKmG2WEdAvoJRW3qIgnI+V2wqLeXkgLrbG2E5
kp6cJfE/wPBV4G0gLgXB60COIm45wKmdMdTo1rZZKlpCIUOzRD4Q/HJYMQiW
fVY+4LGSRus9/TSftxIFzhp7mpiGpjMjBPBQ3qJqfb5JaAu/sMypNVJpZGYt
Eazn+jsfKTPIyzsy1HM3C3E/KWYYnJ+R/BkJolKLPTkO40H30C23JOyuAouL
XSq/Kf9JC0A/0zyAJ3dJdnCGDj6K2mm4QbxfaZsNSbAvTSzr202HbnrE5Ri9
7XwtFjpHQOJraPu3UgrAXARL0UWYD0sNrhOIFvGpwa1ismjGvx3slNnCvyLe
eEOYTO/ktURL9tZcFqgymT0j0Ue/HpD74zOYwhbL0Q5zVBASEjHPfI84is/O
I5UIF3vLQogFe6c9flWRZ4EHWQq+G9LfJyzOFYeMRbD4hWwi0dig9AMk4Ly7
kdWxMTo0ELyGSN2JBBUJzIyaHAr3DAzSjQ6rwPowIUSQAzLH1bkLWp01fuHB
twFd7xQOzGpDnbffnEB//7/5sfbgZnP2kvWP/lGRPTg8kXmXET1fGNvXM/J6
HY1SDVN/7v/dqdWIjZ0cExPaijGphrtMX2SVJTR0x53LOb6LsATj7qMWjHvs
z4G0LsfryooQJWsnouSBcouNOK/qurMZR2eg/6jHWcCCLFG104rhXYK5TT01
8dwjRE8hCQJsXyiXPE6HEyYJuuypSs2oQlZbT7qpH492HA0iF++R1TuVaXJ8
ycHIO40Hpp3mwPGHPBpj+o8vmfnJ4GEle4HHm4aPtLb3kAoh2qnqc6sn6+gw
JnDQRShaS4vpk0/uRxLHFz6Ax8wpniK8ak+8O4oRubFP1AqRsrA0k48BnR5d
d7Uc2fR4xb/SX7kIM2o3n8RgVA5aPuFcG8Y1dqnoTmYe5p9J+FAll+Mb/DJE
SElRnHUKcaa0+711HEU4dgVe7/e7pDMusVvDE+KR4D3aKaHN9z4KAkckQ5zL
nTMufmA/ik+FNHeecgoquLQ6xrBCNLdcziyR2qSG/nbM1Cl044eFd5PnwY7u
J5brzWvevQHhYqIfKEJ61TWeuqDqhumMPlIJLBgWIKfqVwXpctLNHq1QHq3s
Bl0xnrpOxB/GNt1S3L0pJl+og5MfFSS/TFLe77r7WXa43NT/q6xwOU89JvqM
gb9IlKSRtch7szUi1eaNcBLNlOhnivoIELRonq6aGTCEjDrQYdhmBodJRtmt
2FSOLuSd1Gp3BWQ4XV8xc4c+qvf1DjqVqzfjwt6XRmGs5F58nTmhhS1Ftpur
ceR/H0grx1yZFtARJJKFstRUL9QBMkBq09EyY9rq8UKDHSHRz8pvCVBEdUx0
odzpLtrtzgawfL3dMUion2ADea9l0HnpGPBA1ESouDIHs5s5ekBQZwTMEc1m
IGhUPSCNhvkHt0EJvpaMrsx1Df7O2tsABbMINadyQ+OyLfJhSLZ6L2p2ZF6V
6id85oqe4JfIHrhftAMni6/WsWfxr8Ld8bF+GxUCqi7SyhQCdlGy7aS4FO/q
ouIXDQlNzfSOnroiTOBAlM6+KUc0GhhHySZGBjpmAewjI4znZ3yNujfD7aiU
OSjtlv3H9F2bSIx53fT6lv4mjqDp2PWnMvy8JVaIMdQh9XIGZjwMDmr94sKF
0qrrDmo8yVVla+x9lYP2FUgxoRPPb1ZwEeaD0eVTNtw6PJSlb562IYrP7uIS
Xov54Tl+7/utm93m5P5V+WNhz8W2GASdFuuhJ4QTYG7SBkwD/v56pq4wZCO5
9Rc6yIbVY6tzx+SOL0jvvPQDWFsSpOUybXLHIy680fb7Rf0ZRWgyaP9bm3eF
7+c63LhIMdSU/5IAcgYgRUCwVRLLEmaXBvmAIj+PuD9NBXWc9d30yJwnKX4m
DV4pZed5N2+VIHG2qYhB3SiXUqtz/6nF32/QZFFJrFmepfAcik/Q7k7L5Omv
KVsJTl5vsac7UnjFD3N0ddqz179DFY02BmDv061QQ1OvsZOvkKreXOpQEejB
ss5QIEmJScaDMVutOeWbyGdoW2SwwLISTM2nNl67QNOAFUZzDsLWj6SKTCk8
tltQNaKnczjWdzOIpVTOuj894Ljh6IS5URdwYdu9nqnqrtL9XbDr+iFedPU6
bqBLfPJi31uTRJu86MHpwK0Oh8qmkK8yqn9YHx45Z/Msrk/8MifN9pKcyMxE
SozutDjxeoGx1OSdTXdoaiK0LRHdvk1eaMrNZeh57w1Ge7/KCwWhfrcx6+1g
32TvDH22i2F+uZNIs7EmDX5/bktS914N+usb2pp6i9Jaitzgh6eD7lC/a26M
3H3rrpATqhd9LDP905dfTM7Py/nu4JhtN3dREVi8Co1+5a6bax1ynBVysgOM
ErRQxXNy+LpZkfuDDyYpZ1VHp6PwSe9FR8zGtC5A/vqVKO15nLBukueyxEQt
wEJNAGp8G1S2sQiThsM6lZm149XVujW6jdV9d/lATOT00gukFRkK9H3CqvgH
jyXhCBjfqlYWjxgfKhVDmKiBI+86u+S7bI1YvXur5lIcGcyjCHmfLx2KZFJt
D+0XKNdqjvf+FBCnl4PUVrc9COQWiu7rYhK4aFDEFjZymU47Q77cRVT4ajLa
2BKtm59CFoKrUfvhjJlpEKVqwAI9ZMrLmMrsP2mpQWrkd1pxsHQXchdDu+w8
WWvPxMib1m+2ANvZuAOjTSetryJYICPsoc5GT5Y0mH+K1toCb0JL1KzYv+AC
A/aQRd8fVZImAHme+4OCTS+Ca/+ToRv55Uz7gwr2LLMI27PFanoRG9sA+ehT
hkf3RuGbGTpIz3aMEjjwZv5MVNrerTLzNnYKQ/mplznmy8cLP0caGzyKWqCq
zscl+gcT9YLobDI5op5/oNb49lIX4z4fZ4w6OTXAK1RauEn5QolRWZZxpDhC
sfNCNTRegBhrPHP/jtC9DOwTE9PZY51XMKceX6WrM1DKFo08nJbIza4/pTzi
0s8KzkOegmn9VatgdluIpZMLXgl2d4JWdkF6FPm4t9BeUdbyra94UvVzF9GV
uGNb5dFFgoacHXhajPorSKEK4bwImwGOxUzdW4BRUGZs5iGsbGZAHVNWtLXO
TvkBZ0v+IBcmuNC7iTa5brwlN3bqDG6AuUUxZyBfMD8upgIy/sqosLNes2ge
fSgtv6wZthdDprJQ0WfV6Rgh35Ldl9Uk+530kAxdRSP1FgaWsiAoaMQCzUcg
xA0/pRKU0dF1SzGEQPuiusH68/DYptRFlOF6mIP59ur7M3W6yY3xHBupv5gq
w8Xqx6aMMxiGF2VbKahNgX+gV1Dm7BY56TFjiBtGGuVi5XHTTxt0XCFAsLmP
zXMfEtK/hm6FH5XsFU8r77EPDeUywdZT1bwy9Im0OdjpsjWnsCyNOCMBbK5l
wfAR2Bu8nWKeqPECkjmGTJsPD1pDqxMEBdY1GtckRQ6l+c2emF1Z8C8Bq24h
N4t1QHLYH5rHc9xsiAnMQvmAHoSViYp2tA7W/X87BAgO+Y9KEFss8lZs4X/E
h68y4O+JbsUR7FGSUNrUZLu5nbfSFp/ofHuSoXVA76xriKeQCMRNi4CGDMw3
DB7NCx1UJ0yOyCjSJYL/Gk57FHikRM8rqftup12TJUOQ+KLoEEBZFmziZSy3
LUJbfYCl98Ex3AJTxCZjsxueeMrDV03fOMhzlR3TfFN8IGEIN8KRjNKSXBkZ
Ri5h3EfFwx0/0dnjAJG4K6/OqCHm7n/dsPTUPU7AaVpHf95uFbnJCz2yjGFT
Quy9od5fxY2+JTPfKijlZgLEgr8gOSMD/72OUsWpGHMPm8NpPNuekmXkuTMy
pAHujDXyE1swl9y31HGbyJQSQUNLSWytBCrWeqkKYTLi5tZhsYQ/CYmEAKyx
Q1ZbCV5wVF+EjEz3KR8fhTyeHI2/eUg6vpX96OksJxQ9lAFOYaCnVqX8Hn6R
2IYe6BNlzMEuLOLRl1xyVmIqLXConau3Ebh1zJuRpMi0/NA9m6AeqOKaSuST
/Ijy3+0Byquk7v12uN0QbReAowpO8sFE7oiYu18JpmmfhJxyWiGvG0rGIfhs
cRRaodc1PijQsEQ4eXuQ+gZ4ImWQjmEj2ijNftrkyXGZWP3dR1XhmKTvYH8y
AJ5/im1HKYrRLT7M4dttLgdniNpYyjfnvqvcEfad0hnIpj0Q04sF1bGaDewv
iCIobQf9YODat2HaXxFA8RkqLfYjXYq3JRVOqW85yz2tOgDSZuXKgf2ILJYE
NKH6qCMzv3rD4UvyLY0dFRt656JZO2Nf3QIp8SnU0bcyG0c/l5kYXd20zEK+
Usi/8pUaLUy0ECiNma5XdANbwmOcmTBpkNbvULqOPKztq0Wn+c9vLZnqwDS6
65G6kOIDWCIp8/kUMUusROPVQ/MRzz1CkiUPdLc1OXTRUrvcTXUxOEE5w3Pn
ixxl8A0HXypwFFbpE8SHDGdTe7Gwa9+kS/E2nBvMnXyc0K9d9qPjEz1IxCzH
JOlWbv9USOMgJA72tzeodDIJ7Gf7WBFmVccahxsQRAtRsvKLKaE/Io01ARl9
C0NEv1Ii/W1MKHHpHVMevrULpXcw3JCloBe49prsXqsJMbOWZUo6kZ1s2sLG
YHPVdTOMY0bqRkbkB4gHlN1oDkLpOYGSF2UKDnYIJpc0PWp6uiH1GhH3ZOSu
EplU3W/lQWVIbq9NgF9vsM0uemwaSGqnkCMISVQ5HjSryh6wSAB0XyMwYfnj
TsgwNvqUMBsd+hDwivErAXVHKixUp6P3mGjDZ5JqQVizX1ugp0ybXH3RYmuw
IXXfOUHOZOvjlRutw/MKxaIre43djYLH5mBQ4i7tvAnBdL8rFIZjFvxYDpq6
670Xa/ykrQM3yJENcY3CYbjJvJR3DnGJqZP7JVQttqeFDmsG0ZQw7XP4cYs4
Z7mjOH15hZ1SQpW4ZI99zXTouERK7ckojOaRKgWOVA/poni4jt1FPdK3C+0X
LqIevEcMxFWB/Mq/G3XjVellUXVqzOUKiBDyqAt6bAMGahw3jbfF6yY/+8N5
dcy8uM0CsVbd+72J6x8tGBa8rj2JiNwTYSdKXsPyLcnNKVoHWnZMNw+8jbiT
yw4cSeg6fsGIaJPQD7A4ae90WdHPJPSNS9CcPZOPORS0C161GIt5cEhaYfiq
+lKgKWCA9OOKWGWLeZ5mmOKJN04qkAiZpI9annRAJRB/TgLJ4iEOPHpIZFBV
OxrnyZrYXPnIW9tffdimH2TUj0M2thQqp89AvpLfqk0Vm/PC3oodAD2BfjX2
yiwth4t5+N0onUXpwN1A8tHaLEbJWtUIYrsa3zuzg/BYP77VvZHyQZ7rqUak
x6WUuuJxZhVYZ9VPnBGJmVit7nGKi+iRHLOQtCzgieffbRUUdObBFeTomZwA
0rYW2nqDL7vTmLcFL79cyJWA/oxLvNwpgY232YD4/O9I1NHHSqPBv9GEmHjz
gvDLHZmuV0U4wnO/Gr1W2EdzdzWXQKrdz3Z+bsVjHkAOHAbDO3EZGlN/MCSD
S+H8pfmbDHvjnvTsLq9gfBe8zu2F8nxidkVEZQtFpaYsfAIJj1TB5BGCbtkP
Rvsi6QderzqWFGc/6WexiSK2OM9XDvqZu6gtDYy8aqaNw5KQubAbxj8YY3U1
IpR5vfjP/fRfqsDAz51/4j+JUHiaT4NOvsr1VfGQPObv9mtIgo6KntqmzZqo
r20U+AEwP8ur6y46/kPIMJ15FBQBJhgeNw46g4M6SljLcu+YA84b2GzvAkWQ
++dOS8NR1S69u6CwN+Se/60hCQbXFRcdwrCME+D4xaoMvUc46rPLhItGa8NY
4JGqXm/3/aDR23jrXrWg7bAIWE9Fmc7tL4Tj/hAbABpfn8ao7ibLfdnogPk/
PkoeSdu3Y4mEaMQqcFuA8Dz4O62i5+JOlNFjgAOTTJ6vZfs94mguKtlQq0iC
eBb+dcZCboK+6SiGEKH7MQhuolrPAQbfXTfl9FzhJIfHQXNxJUsud5vOFtOS
wprpcwGFjEdoFMloZk72yUO5qrs8hiQDZ+EfcyBpElr+x8ro3PVPBrO0Wxft
12h1nG5GtpBMZoLvy2HrvuvIQDMiDd/jT5UKh3QXV8BzjfYoEfWC0JX7wG7T
WFbKHVPp3mYFk2vrjKC1jzHC2YI06QV6aBvrNXNpcdml+4sKrRLFzJKHRvB8
kHmHbrZy7iQQtvWhsJDJWeix5zbg551Zht54uvJFliWIExpRfICn3eRLP8u9
YE6TjVxx648Vzn0pzMWyJbsgNFi3Pceo03G7EnBtXqMBYhu9BvKSBwcmlIL3
idpc4nxZ5Mz80CNjvVscnrErKotcHy855xb4FYRmmDr+HCKaZIm7T92LT1Na
xrLFd3HarvRMwGPsO3cBe9rrUzr9ycB0/VTZpJf0VL8sZwVj+RdaltZh+3On
zLS1iDpM6qoa6obJFAl0Kx1kXZGxJTPS7z31VspEh1+zMRRcGY1RlaTAvxVO
iKjYRDukGSFr3KrJUVLB5ZW/DP1mwhG+RKQ9sVvyCLZ0ijzuWKPHHHQzdVNs
pA7R1mQewNsWToZy/VzkpA/FsFmUbdl2pzAaKqSRmtDF+jbXWxrrog63GZZ9
bpNafACj4cX6L4pZwAkGarPWq5WHasT+OCHXXpgR4GclFiNUTEqMsuknpVJi
mbP46bIxrRRD8HNrjn5a1tOBAZeC5myLL+vW+h2YErjuppsEBnniwt1rCucB
+fQefNNa+GQPYeJ0fDPtBj9vsU+Wa6F/ZWCyLIiQqZH0WeJvAgyh59S8Rfoc
S+6CVb1Fex2+QWR5zgZlO5oCfwKpMhWPEzjbPnndpqTZFujnMGdY8aw8N4pi
qQQjKdM/R+1vq7kbE7DltlEreU4KBoamcsajvMNVPgMkH1v0ohMRJqreHgAs
rgtjXX2+62IGR79MUI0pZ4t6gc4OGVRdQ/T3Jekd+8RdzitCDXvEEh6fJPrX
4sjDqQpy+Tu1ms34tylTw1Epfbkk141UlZPLKfzHxl/sDjGWOijkORHz2q70
UpqfjCBdr7vV7vxp4ozK70ASXb6WRQrX1Q/p2hshiI3p7lTewDkXMTyWRrXY
6Y8kR+hvgzcVpjKwp/m88ePwSZ8OfNIXQzCmZRereP7CPyM/VJmVJ6+yrAQd
VqUzOUPi8BubBaMSvb0oyI6z+gALGTJCDOx9h62ihipDWj4B5fYTGwmK93h5
Y0xQUM4sRDznFeQLVBTSDPpvAfPlJaqfLrNg1b1G71gksEaOx2h7IdihKqcQ
2OOBdx1si10sTbnzlLvVhSdpyr7m+zQQJxD8gdNk

`pragma protect end_protected
