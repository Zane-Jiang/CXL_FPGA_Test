// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LAB/y7MGWe1Eq/JbpK5mkWbQqz1jc5i27jRxEiYKmTRH5EsQsXtTxxL2X21s
pjTHC4roiXbCI4elTCsdT13kH6/4Oz8NlXynCEIzr8OBdzJWH7rI9umJtHKP
QRC/JwO+ONLLTPfjGfsFnTI9qh8mOFqIr8UcBXbkueiK1ijpsYneBQjkWnCw
sk4hyBDZY7M1ajJHKJHDX4dZKN7o14GXAYPJasx42vze8klG8c2XI+KsLipe
6z3tXTworIqqj0Z48YLb63+r5IDv6LdsmB9PSP2zIZulUWM48IV0zuoELrKg
IAg1oGRJN5JHayxtuoh9H7PbvUtGw26/LjDMhDqung==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BwTJvzLeG4T+bCUD5qS7U+obenzzVs7KOfgNPWK/TAUTHWDrKTQuajIQ3oXZ
adY79yb1z4eB19ganB749R7bfg7GRXgCdpTh8tn15ZSCbCqVGz1VTj64z4hF
vUx8iRCx856sGr12HFVFeYpp9AlCRb3tE7lTPkM+5fBli/S3Lj9EDcweUG9w
a10dPZZ/Ylbayy3r7f7vOn+U2HnwNJJmrGM8pwv3Pp7KGPZIz8QwMBLTVvYs
BxAmfrd1vWPUnWBg2FD9mHPkQdixidsQr6E6Bz45q9q1v0fDVTzN/vApvRLc
Vu6PrjYjC7Hf8NNKjBFuDVSbjlCDUb1CXqsnm+6Lbg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nn2NJVHO4t2aRMPCCP3lRL4LATe7H/MzWfmf6GleHLDTq2/xXyCyUedKHrbG
fr+7qSxqdV3KGlEv/93jx2VI/3PD2FRGyn5vOn2gmIFBlX3Fcf/J/YQWdVD4
9cp3uQPeFXubmoXycLZOk5Qg0pQ57gQS0aHhvaxiLSRCK+5ibhvyWT53IGAR
KPguDa2ulPaH3gcOTzEMjepcQ++gi11Wn7Zek7po8L3wfr9fxkkr3p7IW4al
/PPMTVvDSZlRW4CI0ehUxgAcU8YP1/YhnN2gU6YGOayRQ7PaD6kpB/MkqaF+
655iQ2SNdsK2xlr2a0eu8sC225S4g6k+fXgorwqKEQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EkyP7we/14tX6Jh9b3s4//sjWLP7izucAfIXT521Akm5j2p+wsf1CkHagrI4
9qhkjA3ixap2TLBrPRHsIEgnwU5VL4nQmZOeKCrXt0mZieHVt5lrI0dwbHIA
SQo2+C+6dMc3/xqMdiVtKB/i3rbl2JYTQhAZGtMnf5V8fVd1Q8A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JL5BuxaoXGQjHbJ4pv53bo1BrynuSshw+7yk4jONHcDSmU/+DYxx4+zcrQWA
ciuGIAbqZuNS2uj7/03o/5pNAyHH1Fjgm9eQFEYIUK9B0xJHCRHc02Gw41PX
Qj3tDnaVoFv097gReCyoQH6uGS6QiAXvDfItEXrqKbRLRScFBsg7pRBMjEIC
zc+Ymj7ZrbkgGHGP2Y7SC7m1upvkVsM32psGbhw8gYselR8XeUzg0raQwJcA
AMKlwDoUay61qLH8+3jVVqh+9F//wRSjsljsn5Fx+39I2gHm0msvFgkUxw5r
p806ubRUJD1HdX+tIRhAKzg9zyUKpCwyE9jTsOfKRCHad/9fkwvCR7hcgcLL
mmV8MgnLGCxOUzmA3k0BeOS1wLeJu1JAlQP7sWT/4vpSlMuiISyK2VT/dcyd
p6FG/k9j7N+3jGNnIHONzUgd6qkxAzAZ1wUBu5dYCmDSwufIFrDVtsTrU+ax
KSrji5b4vAdf67EKLeG2FHwvfNqQg/pq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YpgFGuKxNU6esB06CG9VHSwyxN0jH0/RVwTaKGRYQI8W/QjiF0+9zcifsjTz
y6/bzW4DkwBUY1bNeZKyBRb2Mzc31E8vAtyDV8dtkz2ZmYdPAYtoHBAjKwzl
NtFkXq0o+BbSb6ixft5ajIvv8vxen86ywlYxU/tnkMGejXOmeJs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SOmhUB9JN7PtWzLjEx1QVaFN5FjOdWJJwl0IQrVM0bKU3t90N3C3qFq8MbIl
cRImNxj63sZMawwOlQl9Xp0/llL8B+AEai3k3JA7RKBBqEaIIMvuA4ndhI64
A//tPTqGsGdxZ3NWxf1yIQqs3zgky0/MJ7YNxgksGFjoHOcjSlI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14240)
`pragma protect data_block
SMnltiXxK9AoDHR84dF+cW0/LQ+kO7Q5dR1EX2km96meXCKrk6Dgs75unuKj
HL6AASsXsZZ/dd/Pzb6IFaRUaAUuhJNcLP+LMrPUKAbZV3bGd/W33JUI1qK2
6P/RFy+xCAwEe4AIc/8sG9kkf3H2ILaTJ1GTSTBS+5nR1p2hxrBPkrsAwnYT
cf3cHHQ2hJMKKdJ5PTutP8P4H9nxF2dqQZhjsGqAgmMUAAkDWbiKLciOEmCd
IsX5ofrut2HCl3lPQUwrF8KjGCTPTaEQ3QvmoERShmxXBH8K/L7WOKwJkqyU
/tu8SgiE9gggCyx5qmeCa80h1nXWBs85eqwmddC6xtIs7ArAW8wTsxpJFpT4
fdccfJYGFlKdzlSMxLawe3cQdHSC3iZiIx81Lo2ydbj5Hq6iLzPBk/YmCaBI
a7Vi6psnhrH9WHiqztxQKbg/ufMDbVUBuNJOaebncw9XlQad3ZAfdJVVSdJM
QiP36YaeKNNTVUcEn/UMquSR/TPkR/SaiGh8iICKd3lbG2q+k+lXnWjKRGK9
7y5gLl3mF69br+ERfz6IS2zRquWIZjoMIdmMYfJkK1esmKHSdUiSchgN6jYO
XnTOBzdqid+PFV3Gd9UQ4ajVa+zjhWtY8BpXtt6j5fkPoYMVtHHB8h2gQkhT
vFtuclC4Az/CvEMPwwTRjAATPwBsFLHeLO8VTd/Z8pRrUZJL8GmR30nOF+PL
YAT8xQHBQHZXUoOx54CxSG7G2bM8Z+btZouXOj3Vsl1mgXZhu4Cj/vRZ0g/R
it/oSXsvxyzOPDvkWBSE9eiZLlLLz3qUSeJ0gujbkqiKET06EkbNq6DTGyEC
Lh6SFllP3xrL7AhFVM13gxe2Xr6u7JwT783inJlzatlWTl8MQ7wLJSMSs0on
DFKMDWtE9W3NVSTvJNtCCXanPSMIjA5e/PHL/3G3wF5nN4y7kkFQ4IXzF10d
7LKPGrEbOHBL+QH78AxcPPxK2B6FWgqs/2uQsy25tU4e1vjVbRThn6fPyxZf
LtlJ4soicONXoNP99VVDseG6CeYvvuBITHAk+rvuNO5qOiE5sOOKQIN9rOEs
c3bPwsDu0iUwi/ohr2h81r6m2lh2T15G0QO0TtXNw9A1G1zfKieIUKRyPHLY
Z+zZheuLQXs/zdeVvEQlmr1FDQh1pcBcCNQiACQ1LmRJIuNvzPkNalCxqqqh
sRIqFgtfySF6BygrjA+3lV7tqnJU27iYoqFfo0CN5IJTY0kNmwEuova9Gt8l
QX9hTYm2DoIHnsR9TAoo22W2fl5JzIRQQlt7yc4QOh8GT8hvLMv1kepdw9y1
mnoEqaMTJpPSnq7BZoVJYDBRKOSZ5moRFaeE7H6gWvtzTmfLtIm6ZhDtNcqu
AcR6Iouu9CWt/PG6LdwzfwxN2pqepZBq99ABXPyrm3tS+MTfRhwat+dQOYRx
g4KTwSEiCVqSC8RbSGRWtTtzhlNN2K/8e2d2F6DtkQcWSUZoC8ntS0TxD5jQ
37V06lOJp58WcF3S+V/hV+zZ80S8FF4YYfQOwHUY4xj6TQP4GtE2JBzm2RAJ
kN/tumvxqtSymeRkmA6ZtuV3p0KsShzJER1PKm5foPW/mrBwnP0JzsQFQyjR
qK36Vg0/ygnLDwr96O+WfC4rQqgPXS0U5iYt4RkrxiHFN30mHQgrV3w2Vh/9
SuAwwgvrzbW5wjo5t3K7PBUHSi5rKmyY21yG+iDI2HB9ZAaYlGXjmq5boQMW
2xI2WnHZVGiNB3AHVG679e+Wg5Vyw3DEjjNjLAYLgHzAQCplCE600T+G5lVs
ejMLKENYnYoX2J6BOqROIbEI7mB3oxDhI/4QFMOTJdjiH0/k1nErV73JLAAh
s9Prc+E83PfKh4fbJ1P9FwGJzt5JvKZEIXLwWucTYalIR0DcjxeDHDamJRaK
5DN+T726oUnEF32AgdR+JpaDp1fLkkS0Rz8pDuB5KbT5CJsC23ig58mRC3fK
WL11X9QUqk3Ika/ixVAOY3O+pW4tbpR/g0YV/ET0DmdFKMLePogOi48IaqcV
IAN9VVQxM1B/LiQuvQfr+ewEN3ik/DI0zl9j3zmlxVPVYB/uVfMorf181MNo
I2XDw/PkavYYO6K+PeL1pmybAjPdNAcGJhLAULWRQ+iMnCnzwxKdc4QwhZC7
QGLHP//i4+B6lMYwa8QHL+a7aLkGFHME66k9rIZRHrupOTLfsT3t6Mp4bfru
mBxxewdE9ee1wApwughZefOcNGkHEAzAJeeIm6fP6Sv5Rss7H0qfGN2ARVHN
IThIG/hAS9+MSLrutB8xAR97GnxCUxIiXiQ3I16yWDhBeuJXqBUs61DLcZN9
Ak6zh5AQa/M+gI/+y0KyfCYKWAsLnfEaMg9zjZmtGcuuWvabeXIYrIYnoVEx
53owiwFX63mNUmnwwCPPVpx5/ugqzaww/DDRcePauaR+7RGLQIxSMvj5hQax
iydw/tbSBMu64Q49TOA7vs1WhcnbvbsRotPOy61Hb1uPGE14XauOAJmw3EYx
QLdkRmiHNXHAcACNmLZLZgFTe8Hf0OUSbATBeTpHtOwYNX5aYNKM7RoqaI5f
mH+KLkZQW+0Jlgt5gTn7YTrqh0lhQbgzxPEF+ai4ALrdT29hI8JD9MIZG6hM
876CpDENYYoNEvcSOw+TlRDVRmWWWBKa6OmytptUB+8SyG6Y/HaqOl4Sie5m
IwIVKEsolli4DjEkJHpmZojOJ3Bo20kGuX6vjYkt7UQZN3PMoHff6WH7vnW+
+UVABBFg7jz6/IHEC/A+qa82s7LNKIA7GG+e8XsgbuukmcXaTwnG5I80/b30
eAqcvu6oXSU5lDew13r02hS3s2pnCJQxslvm88++GyHiumdFHD2KcFCS4kpo
qYOt+ShwTlff+PRp4RuKSKkpIcjhEFQqN8gI9auUVakUB3d0hmgDCGxHxMcB
OsKvuFLMAly8mE3irwBSRb/mHuom1CvHZqRIXnfev6A1FRIw+tMX9C+gZe1J
31zwhed78P9MvrJNMunwOcSsnAsE/VxY5keKN+YbW1dpkoyv8dmkVDjW/mr8
wN+/JbeDxR4lWLq7yyYtGK5hGxeuglVU8QVf8WSYA2riTS1U637Q/HlN/seV
gG36Ecz05jPVD0kc1gknu2lfkV72XPIfAX7T3+8im6+ckpLNNrzT6AkuSK1X
YOd7obRFxMvGQIfTcWpRSIE/Gmw22ztWbv/edhpVPQQEfHoA51Df8zw11IM9
NZO68cInTwM9PPki8lfPyfCfyZ+HA9nOzLQ+32kBcgo7KkmcG/+CW5fMh4NW
uGKjWRz3npTxUKx8N0Ic0lb5XI6E/ong73Gs8m1v+B6bvzmSjvtN0jPi8yIM
e3QBXM3ukLmUfIBSVaKcFHGmrPPANIyJA3slBHxoQw4uMUGKUCYScK/4kZjA
AZ3tYfkB0Tfk+YAztp2iUrfsdvP9bwijoNytTWz9Nz0XoUe97AiEfltH1pqE
uzOLmhtEkEFAdnVWVMWku1TYHsu/HLx39TM7k6E49mUW6UZw9pE+OElFUqvZ
5qkLgGvGgovHtu/5+/SubTxUXBlos1ov5JSpz/Gljy11N8Pg2Nf8CEuFDpZ+
FuWXnnBPI0cJAeLukIYQRb8GfX/8hpUCJb3+YDgA6m0aX8sGNWml6Grm09ef
OkILN1ljwnuIvl60XPnqql/rpEq2pB7rPG7WDYuie6FYvGLPEgJiXOO42HBv
d0hLqLg7n0BVsiY9DNa/JzywadhKpuoD15m53PgWANzr0/+k8W9Ve3PO5FWa
Q2IOLsyqCWPB35PAbiTuXNGidJ3vhwAzJWxQeDGw79321CfvD89fvZzXqLoZ
vqwLH/CO2Zf6vZVESQtJY8uydddfcojSi7HqpC5gOkvDxDbV+xZvqgCpc/be
BQgSjkYAKHYybQoCYllWNSTyDSMz5EntI4eD46EVbw1wqpozTIVXgfO1jRzi
iB/GMKItkx7sHuXojvtJT6EUMWbsRKpt5UlPLmsGUgi+KqXF3sMOGyWiOtnP
HtpAIIwDghb6cp+zg76P9O7Kgaf01xmt/2n3EpyoTQH6tdI/fIYJOFIJ0wUS
T4F9pTnDKIfbcbO5Pe4FUqQFmTPzyGmJs4M8w+k0bABMIlrzN6UwVuzOeXbC
V1zyQSQYbckRqOwGpIzqZtKcFtRAbN7TL8oNc1m91aZkf0oWQ0cEpzgjDOz9
VC8uYseRjKrb5EPPkdtcoShnRltnIda4Fah1Siyd5JEroh8DqT25hTWkdtGR
88myviQA850K+dCxVe+mdN/5O3I3Sy6IvZiizHhA9gCL8fUewipamjw8xH5V
jrI7M6xpNUaf0xPYJfcV9K6mm+1y9imt0BnBhKlCe6U8YLMNSgFpodNDXLm6
jtPJMTJaOT8lNmcFW8WH5xtVnk2JJ/H2LT60zWLMoSrMm7EKlhO/nfphUx++
4i4vIdlHR6r56HYtPHiXodBbfEPDYUR3J+BgjM1GIa5gLNJ1nMGkbY8vlwUi
nZ56O1jnwK1mX/nfXcJviCPzndHuMimR0nkHdivoCzc/E0x3c96t8Ar83MJB
VbckQ///Hrh+U+EVvIA5hzk8rqDSaM6/tCUdOBaGw6AzoPgtlCpWRniiBjH0
JUK3BKMa2buGjFjBNWagZWxNgqTlYUaFYqgdqT7RyF781ApgZIRRjRh3Iguo
CbIpXRogHL3VgKhAxCUef5njZLzTBBIQvcjZ23eB3EXTnWLOlkA7Pc8aEJR3
nNHu/+DxIgQhQLKojhe8hXSo4WlCfUOQl+mCktnWDRrDnDFV3L8R8J9oVV1B
QxE6EmJ9ZRaPH20yPPY/JuLph80NT0IyprO/qOq5+gD/J9sGmMldFfW2LFRI
rnPW5MybEODAQb9rX8ja7rh20mdekXu3rCWquz54Al6z5Z3+eaJGg4y5qNqM
2cNRJob7fr8ZbCLgbq9WrnbTD2m6MJOd0z94Rww5F7tsKfFvpSS8Or5eOK2q
it+McClLm2mo1yvxfmereW8o/0pIOIrMS51JTfcqAN8yQH3OzoiojPeylfoU
xOkQmTjSF+mB65DXUyPUFe1oCoPw2oCRdhiDCBwe7vrmy+46c5/8wbq47lLY
Cm0aUz2BI8x3JnZOj0fO9Tod57XTiyGffiAUmNOTlRZn5KP95QOcYWllTrnA
mCGqubz9F+FcfgLdlQKzPJgrhlBvvC6nPioPtg7IQdxsyWUbQadbm1cMv4Lx
Bnv7AfOscRuychU8uryOiJuWGTT7LhEiH1GzSrrBWXxVc891cdSoxGihhbz0
fEDwvdvTsUpStiOrHkq8lYCJiRyrjza5NV3ewC8iNQqPxgWGocUUGPF5M9dy
V3EkMUhyAtnx4stGWrCmtz6KQ9d3vgPE68FENi+kYdhjz1XzsTFzvJDq7AHA
llzD/2+dGpRDpkvIKlyXozXCqw57GnkOUEOjqboFFAyh1jIfYiHwaAtA83tb
rrloiF3KGjCMG6yhlj4a67YSATzLfSDj3vP1MGHCYumiveQKt2NjDlhl1lXg
Kzd9sEkCPEsIgb/K2nko7qtyH5NRUjECHC2JqY7isSngq0w1CbQLGBanT15W
i9N3bMi4KLEV3LmB9VGvW2ojO2bpI7+6sNLS8EUDsLnk4wKT3xOGcpZyBJRR
ddqq3nLCAfzZmeEQ2da+3w70x3lRLk9O4PI4gQbz2FDETITW8jmUuAwjWdKN
NLhyEQM5sLhVEoIADdSJey2g5UOV/H2RDLbub9We8b4f/oaqD+AS/TpSjh6+
k+U3alXq+VYqXPwXvLbjKhhcCPeNLs+Z1PQ8jvZtt5kCGRMSYm9SXh4lWqfz
3k5byMQ92+Ijc9PGuSIcV++8Za26OkvmfLrZDPeZa6j3XtYWL4ynNOHgvJvz
SYEk2lgQyHwoPz5XAxot6c/oxtehcBNaQ5FLKiFaVquNKNx3ZeBNIdNGEhBV
MW4Ke5nrSn+uRObOsZ+417FZoPPNC9e0dl8ofeaaz4pdnPvqwiYRpQfJKUVq
UYX9TjQ4sdOtac3bmVeWW2AvwsZixT1N97pqDnky0TKxKjmKRzOorZi9mbSA
Gc/l3uba85yRRg0EiIJRdlACFdMMN3tM8m20QaC24ojScsDNPHOtWTERta+G
QvQOhHg2mk5n/kXRpSSLt6IZVDK8Byq/eOBo0r+5LzYUxFRPtyHCw4Qw6heO
3UeMlRRKNDFqtTZ0xgUmrt0JO9mZJj+mXKup8sQT1HWIHAqC4eFpU9fAiHgi
rP53xPUP//u89naXX11YaCBKHecQUfI4Pt0NJf2aUHhL6jiqIR8NfGhl8cqq
cCYpzv37waLZt0WNogj0BoUfmWbaPVtVL0kljG/svKN66mUqwNwpDlMiJx+1
9ZAq7UvpeGS2TrdcF6TIwZcRedDJKRuoTUOYdG961jNJuVe4b1/8fwvoWSP8
ih3NVwV/gTYkxLoNpNYhGIQFNtRr4ynjhm3GkMYOeKJrPufKnNb3iS4zSO7G
BBGoWC+ED+Y5s3iynfqD8KqSsmkjvo54Z0TsViAoYzXKBgFTT4eygqSIjQpu
sfYPTMQ8gi72Bo/gNm4yZ7iGfpxcFjncxIqZVOHc2ivhXFQXao/NPOhg7t7o
FbllEvAwrS++uNcW3yAuIW0IwuIJjdkAsy7gn2Ya9jg6u++g+dQFfDetf9Lj
VlOX8LH6zQgnAr1xxEFgfi46XS/FRI5Scc8uYl+OGEHoU87//Kkp/Yl5U7lm
qpVDEbjBmo/BZpB5q6Sl9K/sFyvP5KcHoCp5/SAfaIoa8+JZrtuuEwHsgdr0
MBHLk/KCVknI4YagZ5PPDe5myH8LOs7gjEJzICicrfx5V0pQS9UFoWGgHVHD
uDiD3ZuyJXih6FV3mASuaMeYh4L3gywZFOwZ9Y2ZGVIsMXq5MeupPZpI0/U7
ilfwn+aZB7QZ+48GrsgsgDdxvv01fha3OgsJLJblFmLUt7wnoN8UZW5vXKV4
JoXcnMIGkMpaxPjbagVrravPc1SFJArxTSEuDUNxS2QV9NqlUVKdy49g9lhh
fJ+hR1ppJdeIMroRWRTWjKYgZjxfUjNNVlP57vX5yCm5RnJgOEfg8ynApWwy
XXEinV+JbldWNHAYd+rtQZLcYZVg8Cfl6xIAbeWxf7RhoHVL1GjQky+QCFYj
ltINZhXhsyWJuNb0d9kpAuVezwYunMPpP20RzdRatbkwi6wO41n0OzaDxazH
Xv7AqoEUdvqF8LG9MXIeOn20Vemm9iiJowzinA55ydk4EJTBs4CWY0jcB+Hg
ZvysT6+0JTEJgwiKZ/SMSv12qebBFN1QCpsk0I0p+/gGfw88dR1i4uUnTs5m
yyXMuW1xKggqXabFhAy3su/PeUdPesx8WP9FCAqvvLyaC3o+OeGC6RqLBiat
SIHS9qvjIbf+NKfGcF5gz24o2ZdtLDRw6FYqqoTNHQZQ3/iu0SYt26u4LIhN
QZjSdwWELtcvgjJKGjC20noTVN8j+AKIO9do/eCWJ12kOka8km2B/50QH/Fs
Hc5rev2VIJqjxWh/n1wb/j7M2fgslv6025fHUYGYrgldbsPUYe/lFJ4Ve+QE
/CkeB9ZzKeXBbVooHTE74g2RKAMh2i3QdTnHB7Q4BgcSG0WgSa+vwWt5cOcM
5Ge9DId2TydMBih7DUhcU7DLO1go9WXsrhCDmioeAqlUo+zXhNWYoIc3LCtL
PkCX35WS1T4La8ERI7ubtrInOxZSjI9viz1dKR3P0m6Yyw5NLOC5TQ1L+trk
oPtjW44/SfSPf1MSbeR9YSQcb0A8YXryiAYZTc0NeydzamNIhAD4DI7smQYt
9+xdpFtYGKWVCQqZ22muWSCGlzUJD6X9hRIAmQFBI7XFbw8aoWTNTFxAoZcR
xXPgFPerFUt0EY/mNJLoxTIeCO+V4FpHviPi0ZQbF/eA1btAE2xM2r666k9l
1SC3aPVxdABrb2hVLHG9K132SYDERxeq+D3EEQBeDfY/aGK00SR6ZsA7XP8Q
NiXaTOj7qcq/Z0ubIdmm5uU4dhUEJ6GGeONVV+fen0OAExpSlcD1P3c01IH1
nRZO+tO+uPNfLN4CNF459vcIp8nLkU1ukkc1/tUrB1huLQUbP6gBRRrSkitp
UcyZWLu41Bn4twuliodh/NVpDDDnrR/vmVH9thWsy9TtHqFepCGjteYzF0iN
Ag/OZqWlMPbLCoi0vybVhWkqN2VL2h039nXFddRCoqCX7U6ccQ+IpAi1pRxc
JAAP6xgwQZAjp5/OFqyrkYPylcVNl5SNmzPOJnJXoPK96fgSp4cU+nRuxKMF
KPAiOn7X+wMzjNqoFpHs/B35zEBp60LYEaz4xsYaPt1NR9tH0TZOkU1GVJz/
7UB5g5eEy92hfwwmACxRUXW5W8OupMAf3lBf9FW3cLW0qqiILrfy1D2Q/Abp
9pKSm7HnI7kbo6LVu+xWoODqpR5hI49tZEMky1lRdcMpZWW2DnAHoC4Ro1ni
pEbxcEfxDUZ568hMiA/MhhXjYZX4mCuL646imDuw923393PcVXNAE/Vsqfrv
d0NUOQYN7ApcU1bTe2EYI9xJgzRTlmKpxgg15R/zBPoHoGXpOQbrjEFUp+BH
Kk4eA+dekopuR+IGNEY8+g2cEKWE+C92zvbORWnVMAIOvUSzchQ9EzhqnwMs
q7omc62fKyB5wSAaorg9NVciyCcyoAVmmRyczD6CBMCFxIzo9uAiEC3lUVMB
XLeMMk0tO/MkbrSzTh+4RyZDdSkLpv4046YSt2as5U9lKPusFd0/1PuQm5K2
9I4aphjXVwGkn52uLgAbSxmWDM8Jg+E2qa44nx31FLrYNFmtiTQ1quYcOUNl
7BvkYZnB8PnkDtJetwEDvQPsOJRnfO0ypa3IFvekm5kolt5cv4pIEzIuLKzc
x9OFwi3vhSefVpLc6eD7L19ACXgj4isN8nMaMuT2qkSJP1p7yjs4MhIiSj7p
Z2mCnZaRNR0Lyp/A68qSwA9v6Eevv/UWl5dCX/mo2FCh/hw+yDhNNh+/yeuQ
9OSkgE6/eS6DtqNdgBPg2wUfKbqNXZqv56ki3s6zUunLlJfyQYEOqyntT86O
Cl/VGWOso9TMfxHPzB0l8kO58Xrrd3tuXLrvntskF8dL/tsQUjLtUGKaV1+0
MJHrxkpxRfKC2x9EVjFzipCTkgfUPfQKf9cDR+ntqkDQcwk6JKYGCL3I0IA/
YQzhkcK2OL7sEsWyprJpX+VpZhnV5up1Eng5psmYe26svbFmBnhYqUVpGnp9
jfwohGJsrSDq0LFfVfh5AD9e5TSFZRYgxBVaWmYQMUtgfNz5jXh7e8HIFLzJ
5qgf7JZ0r/bQG1osVsTZUZS9g0A6YSlFqVi3aU7sKFwSwmSX4iPt7kgyW5Ns
fWyvxkUeto2uFLM+XFGrDlNmutnG6eIrmqab4W/KlZ1Q8vAJtRQaDau3bc4h
VQ6Ykf/fbPp2X0R+LHhTuHpec6F2k/XXRF1f4PWe+dvD6X+EuBpufvqGk82+
ohPn92131OPCRzKKv5dFF8Rs4yVQD07ScHeLyN3lRpB3P4dEV+uUBHVd0m66
VlqDx2cEjjbXhTsgjCkZZsdtsN8MA9zZCxmyP2V6vVzz4TZmM+vs4+mMugZk
v8gVsOiMkgtI7F5sLXHZsOAvtJNZJ0eh+3Jg5iHH+4xhd5/LwEyCnJTrl32g
Gn7rIZfJ2qndb8kMwiJKKF/wpoEjJ07gjRZKPujjV5mMclnXiARW2a1FhCCc
w9KCg1oJjR6BQjy6rQLSXG1d/r16ZIfg5sPViMAd85p02y1zrfrKsY8fME0E
WHtln4MkLwNumBas3cBjjkM8BcCnU4Ujt/X7kduV0jxlKDKimZ788TrpNmZV
te2WTpZoMOEK6F/SSeMZOJTuJRloKKxr5nGmOdUwFLbaIopTuqnnS0pobeIW
Z7QF5gN4evDusoaCKh4PRqnRt1hWn4swd6AqwBAcRNJfAXocDVVNUxpPYgWP
0tNfesTVSvjVquv7O4ITY9giZAJIgIC8TAcVY8N+YIZsNGD/f5zEHB88IjVs
IdboJrbDbP1EylHbGgD9oK5oyAyw/lj0wVlxT9FGIKvcqskkZqMhH1aQqUKm
nJ/mrD9ZFdyaRvKRomWMCpjvq/uRHmGgwoMXfeyua4PK00nXuKJaBx/gGdUq
ePsGfITUR6+h9pyeKdGec0/YiG7pJxkOibb4vpaqlz8pVwCJ577G8kh13kDO
9ULxgDxgBBqmaQRMi3LOUCj/yTlstiaY1woyCfUcR+izGwcSKijOP+ehl0bn
v5uw2YuLXbzOcBEaEt8a4FxYzdVNXGbXdrZ9iS8EsotQxDuU1zaGmxnPJG8p
4/b7iAlP9urVETS8YEHzzhDfbS4oK9gRqaz6gO5GWB3GVZNsxYnAbgcpgcyg
Pcv9cSBdCubPpDIs6cchRMxz5CHo8l3CMayBf8gQytBdZOjtiy5MfSrCKM0V
9yefxliFj+PHH7WXsst10LK40VAylvXxzidvK6uR7XreQTKzjHuSyi8yAwON
bZtEvZsDRxLis+cfVy/CQPtiRxQkc+9IFoGx452XhFKHGFt/UQTzJ6sLINaO
e02txhdIqyB4dQfPNtADegeYOwk9KIWZFwaDubZpXzl5f9HqczD9SyGaAsYW
OusvAwmonkUjowyThlk7XGLP8zkjcz7nee77CaBLSmJws/+wij63w35fAQNN
h6rkee7cFcuf7dKykVUGct95SM+LwvpTIoTJ7m6GsrAimO79u0rFQ4z1xs4A
Ny8lieg7+292hV72w6Q45fq3DBcjTLJMw5kk4T1DdJywNuWtSWsjf7mKhDas
HYXPC9yL9GXRPJDFAiDG6S8OUV75xBiuuIg2uIxQndS8SezEx7SsbtXjUb1t
19WBixOw6T9vdMHzhr6q+DKzWlob8blifDGXgAhOvTNGXqM9l1f1V2xxaEmx
BrxxT74dLaQLGlhB2sEEeH3GnDcGd4N/bA/uHmxRFBmROaWKc3KYnABIwMWt
nC9Fj4U5iww/VMrHuw4F+Ke0Q+iz71bBYNeiBkuKC518DFjAxc346mEjJfNZ
4co2HX85T/wtpVvtnaVd+htwzQzFboB0QAbeudwm+XoLeWh2PdY8UB8P195b
elhKskmqgmGVzKP6ytc0VpIozS7fYy3Xvq4YGVjY1xfxVkLbnQONll9K94fe
eXCU/f+goPenZMS3ANAvNjKxw5FqFIxXHIVHzXyWvdF5hGOY5bxzuuowVeys
tL6gLUWSjse2z3LADh1mxNxbGilN4eFNZTMsrhdRMIcVhDg50/zohY36hdZu
IlqlUPhfKit6Mf8Va8LJq+tOqTNHRnuSW0ovWz9grtWZhF3Df7q58Hfh90aa
xrabQHj3+tO8RZocR3+EgnuacgR42ZsARyiTGAx+a8ZOfvbJvvbTFa095kJG
mWmJVYS8W4W7aWMXj8i/5i2DS4jdLV2dkhg2MlncPfPkIuCihrneqqELmBu2
Zo4e5wWkKrXtU5IVkIt3p1dEHlwxA2re7OLiIhjUXRPFTSu8tBHWIeM9ahNZ
Tlbx1jqCcP4sWAUInWaXbEXWBAkKMOWArDrTEgeYmyycuAw8mqkPPiWQypq9
Gm6kreuTjU/JHco5tQUWxkZz9EOj+pfqUvROH1dPzjF+hL7JTO18X2LJ2nFQ
zzOUb6dLcCT3ADgqBHf+ySeCzc069fyNVaBMLy2TWEHB6gwIYZiszgTjPQFp
I7xUJLyltQifcJH7y/TgTITGlWVCrA1PZQiUTBuaPFKchwOWO4gbUcyjacus
3DZhNI+VYf1tXInCbJncYUySnWd2u4JBsUkhLGHasRBzo//FB9yKNZ5aeSXk
VBa27JtWt59XOrS+kIVfzKnYtSXHQ080rwX29RaNYTzVscIJOcvKyFNBMhVd
DY2W7w+sC8NSXkCmx7arHA+4JjNhxHuMZJVFAHiQ4Dbe60tk8mpOfcjvv5zB
LnF6p16Cu8BsXzYVjAKonESGcGWH3nTM67tYzEWE7M16hUFIrndJ5bA57Nrq
FHl1acWddnhmxsm3fEhNyymAkwMHuidxAVuY8x8SdSnseda7bPYZ/1CreWnU
p71hURHjoThu7c9wVVflT1j8EWMzvWhXz8tA5qnyPGZEFfxc8OzniGJnzRHw
2UoVbkLYrTRu4d/tROqjJIfsPgghw+pNoXPYSzqtZNMAmMwlkOVzc5BoRq5n
l495AIGtL8Kb4WQYHfPSXU8ositw5Bd4VL5g9A5u4dc9Sxg54ioBnihKTc8O
YJ06Eot9nDAeBfbhXUmkOH8oNSDniM6FEsBTA4ROYAw0G9LVWFOqtyonDf35
KTdjN5FYLeKmru+JMqkIEUvLLr0HBwrA1DTztY5DMoJse3SEndjQjDBsgygR
3sGZp8ZbUHEUClqQgriZ7br5ZLehRzVOR/y4ANaeDIPEexPFOmKJ1g8tzFKM
6jFomfWX7MwVIKWZeNJpEagpld8ZqkrEjSWLAguuJB4BnEH3NnBbUCFCYjom
Caw9z5EXBeH+ygMs+fy2+mPa9M3j2+s8UfolTK0pYB9OrPsUvMzO7Kz0Ggcv
uIE77yn0DCQpniRYQvyu6rJaoNfr879n0WHVCQ1fezngWEOpX9Cchb68S7yA
DXZfV8R3X1y2dKbWQBYR8k8Sxjmkd8zbl1nLrznim85cWqCUiLrBxFrtu0vz
iNANQCMTt5dwY3X6T+UMgqfUzuep9NWJCqu3nLt/A8wb54RItt7xFVfCD9B9
YmdvLGgm9MQXNlcVXzSiCko/yKc0MtLtstvfAbvR7eIPMlwQtPSzcaNq6aml
hQUhPHr4JDZfMJV1PnYDcqgmi0U12SEudu+BhsutBJzDtHFe769FbMY/5xgo
/ed68tlmx6bLbmdO6yiMl6qJzuGLDkPvxGNTfHBJ32Al9V1x2r4IC+6c6mjw
a1/byvVDpok6oU90MmVOi9/Qz576HwdAYRWvpL9gduDa9eL6uqwiNeN4vPBM
nnUnI3SusbDjoX3G8AAZfzkjHaPsivuVnj0Qt9cuhZPrpnMw+uGZQQgA05+Q
c8ZRyRkFSQqK8dpz8Zhx4NOvp4lA2Cebirrue/n56xOz/py1FuZks/P/1dAO
zAk7XMZGolTB12FgoH5vXqQU/w0NLv8CTT5OI57/TJgbTlhlhPyb/VtT8jaF
IxEfonBwADVMBwjQWpvfmUmrynDkjihq9cZGxfrFBLk7l/YTssOe9bICHTFO
ci+DRYwVPS/9wKHO3vGb7ngD8RfTw0bkFaqMuTqvLEcnPr4oaPwFAG7GklAy
DeM3S90JeQlN4hwgIyIBddLcuOcCkaRWK5nF/v7BVZ5IQgQeAc3ZB3+F3PuG
ombQaf3+fCw7Y4t4MzQCVDvQC6oUpzPTHXnRsrIP51LTmDAzh1xdKi5gsnF8
OwTSGL6GY1iZz4bRYaUR8OI+2/TYie5jVKKJkR33sL+FlrwUnb9BJwlASOQX
b2OvItyQpTVRoLkB2YRCF3DZ/OIa9bxBIDXgCJ1FuUo6lZ0PLhUrS/dAHFpk
oreuysNSCWSLBijyHG7jkk+Tsfhe5l0cgGTQeO1uGmj6PQGeN0XZ7xUVFco0
QBKVkKvehEVYVts3YJB7IQCYKHdrNnq3Aj1+a/1S2lPOeIRNqgRr/YWRkURa
hcaqjua/pLizl3xmm98/FZmAOVPVOFI403s8DHDzFHfGxrdqKxHnkFVZ1JLJ
8eJhV4CGAnrFg/bRtL+J4kLXBo0ZTWkStRg2mLne+/+bTVeUCGb+LXN8bPOT
OzWckJkqkoLtP/5nZJFzQ2xNxV1jdpm+Bm/0Cz2QGSk5Yykc5Zd6lVzpXYHm
2P/PYUTALwfNpqpPq6JrH9cMqZMq2YPUfiwm3fBckWqQ13TGXhV7Pgq2Hr2R
/nvyzWxt3D/4qFGaSfcxzPzOMdwuA2f99wr1b87TuGxZd5M2TmtsDqtEoUIQ
PqeRzjLjaLc1jPTG4xPMiKfw2VJEuhmq9N8W8sEPKnN0etkjX/UUioEmokvd
EdpnWRutGTfVLsz6hf8iGFMTSKGGX26B9sIvWRDwVfGZPTR5B9sDdwfusfME
IvDXY4Y8wk5HQwqTqBx4KhTqmZF9kJB5ZX8FvWfaKwPe3jxPNcXrlHvcJJM4
HHh3gc9kNaWMZlW5uSSpR3WnXszQApeES0HJPfCqpRcbcD8BwiM6v9CPEfGL
372R/H+t6HSOlYA2A2gQCr7vQfvzSE/hlBEhRI9E9N+We5QdqsrQtE1c8k2d
0tj07WSAfnLRuo5WN/EjqRUJZe+kdNehTx4njLqqrzTkm2ooXDSZ/RwRvNfd
ef7iSHuFHh+E0TVehUKhRTIunx5AtrPHC+d63/kfNNtn4Yf2C7W6tvqapSCu
K9GJsjyZTaLJV2UnMHWflTlEnlE9ZazlbjjGhrLahs9E7dEnRhASmdF4AQ7N
hsYXXj56aRLqlm/GJbxNfVf58J3LlbAFD7K0TaVpu7inRsd6g3nsUKwCdWgJ
VXd55sXvAfSeQ0jG/3skj/ih5B0xaIUr7Zbfg0H7dHFzONKxFWugX/S/yxlP
0iyJRyzJiVyCpfGeiwvT5wqIoTk9gzpkoUDRnutDBwU1X7ZotECkfKAZ6FOS
6+QZ9GTkpbgv3BSX3xPqagm2WRQJhhDSbhAXqaG1k9sjoH3L+gFz2bG/8vJD
EXN6oFE8vCUmZs6NS1LvHWJOMCSVCyQ8Y9+TTWIlhSq+ufNvC+cz6HijvfLe
lXVkIQnmcmZXqf6SNZR+DDisV7bhj87qe7FJTfwiC2vZC2R99KlfudH2pi+h
JxAWRKN9NFaJiAga/LhcsbhSkOPSUmV5cFeHleitgVz70gtgZM6otszBYPuh
jwSQYAbwlWWLzLveDTDFU/1cRg6yuQS87hzaCgredh/YgRftHIE8m15LMr5u
2l6KqjCtDTM21a0e71cnTp8J2EA83vbvGoQ5R5dviZEZQZxSMPnsSfks9+yB
iNV1/AIYlYBFZ9Cth1XUnnCJ0qSTXiI4BgSyDPtRLR+cMxvSuHnCDsy7o6Qj
Z3cmS8ttytrV9RYCtyqMy11Y2uLVvzocSOMbuT8Dggtg2dxfGw2pwo3y/wkY
ANSCL+6Olz/ikfxKbbID4pA3czPSnL0YCZtPbSbignbGQQpugt0y4Cdwojkm
48YiwEh1VWhw3SIk/2/L91KjJ5m6/uS9R7igoJIjkIcwhaVKX/b3Fl9ES75B
4tZl+5sPY496uo+6IYLUUWy7cXFD7pSxzw8QQsRIlXM682hrH9b4GxmTCZUn
MblB2IlJwmHNyca9B8epdcJFa0tVljkCULj3DOsuIKmSG4B2cFYavlSzBDzt
8YkDRkvZon0JO2Veu85G2FBu/mzrRr8cqQL9OtUPJBl8jo+sIMNlZT3Tfudj
1zbtMq++Oz0uTe8zZm8xayjlYB+QyvNZRTs7IlrsF3C2nWZpPhXSCTuI5kDT
BbEdsvBZcjYjvDXP+iTf2AdPr0JBL7s+wSyl78+pxpO71yQ4ZLFahRDa4wYo
Tj7HlU+/lQ+txOj7bWLT9E4aVgJYRbLgnhSlgAXJwHHNH1zX8o3Re69qiAJB
Ei8/IsvdhKKD20q3K1lwDVL9Iit1yPq9w3k2axHTNbM3CSApUU/Kl/VlULgA
JfyRlzdlqb7iR1aTuCHR5oFGuXjHlSDvwg3ORLyiV2EpKrdVvbh6gm8TtXyU
O53+Czbl+wYhJlQrwXF6B0pLjL7i4zFSRQOu9Z6GuOc5N/k7n2n+UUEbeS/l
+k3FYHokdW2nLNox2G0U+MEG9ek7bEfdLOubtiUDjbVFoC36Gyp9gq0eEOs2
uxZ544l/rxVFDq7LXrcN0+JwMxXI+RBoOJm39KpJMxu147DkuwBK9Q/wJ/Y/
zgMVmBzfVurqtnUU1XzMmSgRQvyNs1hJ34FrBYaFiRKV1W5oVhkHvQPQkt/m
p87lubJNI1WhRpWgigwZ6uZJiY2fHRM57ngs7nyVtkpKvmPvL4OfzQ2Aroui
uKycowukGpZJ5pNWEAXX2odti6OCxeh3njaWi9H4C6mWepOMNLXIfursQmOB
wRUz7asILic8Eq/A6zB/M1bxsOp6bR+xt3fmoJHf+osBmhiTUuCdMNBpW1VC
tLB5MgbiGNYiTDK/ER75NEt85tUzERHlsFgiSnErQ+RE7CCx8oKRS7TtVIKM
K4I9ux5wueO40kS7W94UbSltIsUURmGUvQ7GnlRUwPtXdqEmarDA5shz37OR
Ll4VSTsrj3E51Am5F5wR+Op4Iqdga4QvB2rA0V9vibpN7ZfHqY6EABYW2yMC
841Lp04BNOn9WrcFINwMb9fUZnUYhrGPYFUB0aqjuPuoDwtMt9OQaXS09rhJ
8JoTB4zVy529S+XG4YPnhO1117iqAWuDxI5GkK+hRri+gI0mBORgS6bKzbpp
D/HJ7kuinE8iI2RWxCX9x3BWYAGxNEy2JIR5WwQEZ6B+vagSwAnRDF45Iebb
lPkmwCHH61FwAEPiV0dPjFSMn9RgKKllmzqg9Gr71mJfanYS6WznS3IgFmvQ
B1PwfP4q0B7chA/quvE8LdF+p+RtqY2ozeVIKNuWKijMfn669KxV3l1/n7j7
m6FPuWIUdIS0gdnjK1s0jE99c0eoMB93sSlQeXWX9z9BNZag4V7Hx0z5ePil
/2qGTlN/kResowO54DSsQoujHT5QXr7H4OypkGiZShQ7hpRR97iV7PpY1E9E
x0L1Oo1bUoptvWK4Kx7rhm5OAVt4yMrmJE8KYJcyf4zKnUtg0UsUtnXmJHAQ
5D3pjM6LPVqmmAA2f6IcBjhR+vueJoNcL0TAxFu+gHeQDjAM6GvS5H4O+MDr
eecMpaml52aj6gilg8GFwVhbVo7pbg0IHusmdslWLwTieLDlewV7ks5baz/1
4MUj52kfmqydsmxViUPbFPMRrAN22TOv7E10aYCV1SgSICPCxz2Z7rr5SAdU
HFaz32H5Nvqz53U09VpxZmDLe2crBCpv30YseH9SNl8VwXrnyDLx4/HkBWg2
ovY7ozYIaA3DaUXoosYjOATjaRwwsLv2t5Rqvx+ZaXDpnpHb1TfT/Rt9TVMo
d+PT3JsLHXTDDV+UnBx1aqyIQBAfYDgjzr9RCXdh5FBn9pw+xDhV4JTrb/t/
Aeay0wm7BYGUjiQNJgzZHzNn9j1MZhwNUtbSYVY/Qn+Aq9MmM3Rol3Xs1Ipm
obNbZYEi6QHZ/hLpqORSbqII0rxNrU5s6qwS7mJtoOdo+8hM2ea0xB0bXlZD
/RPwCDxq3WlNesxD2yNmL1B6VANFaMj/kiB5lACjHnjRlARhoKE1xsBOP8um
lIULyGFnyhL/LGnRP+T8cpiMkrU9hQmzIMVYvXyxYLH0weurXdEyn+MrMQ1R
JovhnzoKabBFFmj4R6z0U8hol+J8k9oeUtzB4UNImw6FXarwP8xwxRFtMyt4
n4UG2svFjQghfjgQ2aysYYrl4+0+UDuTMS6XkOgHTaYUcz5u1xaWTR9tGAqa
dsZ2O+9zDOXymIQXU1YcqsFnxWxVovZqlVU7tpkndChLCQOf0GG5EvLiTnX0
NrPO+LQJbCfJlGozs6+6oFCaXC7H4HldQib1/pPCMJVjnjk60kAJR61EqUen
pLMvYwIGeq3M1L8ohJweGA1cPzSj4K59JlzIjm/1a/wK5oaBrbK3P2BEHaRR
qhmMaAJWH4WY96p4fCZJaMT7iGgU5iBg2YjpIEKrPc979HMojve+YAZoRHUC
mU3x6BFDoAOp1BpPAzsXLepiNgWYjdEYwTI5hpCDzy5aIf3rD7YFXvCE/n2k
I8uZcQPerk7cLFThijsH5E+VCHXXysc5rPQE83Sm2niBj9LfZeAZbCBYnejt
lfJvaG8beD5DVC41dPFTmpSed/Elw3Jx/ajsKMiBs4AzVkqI/CaVayCJdFLQ
Gua4fXifEGIRsR1474Kc/Mz+Ovty3V/qvUvKgLwwIXpzNmvgRekYr7NMwia3
FFSSEu/ZdYBLis0dr5AydNs9VncwQTcb8fYQw5yPtUHTwKuFWN8XCK5Biaxm
mNeuXFwvQ10TUIP8tkx88CXcpE9bFookTB7VcIR2q8SyNQM55dgu6gPjqRea
W9Y5JveZSrJzcQu71JAMd9+KoadkwSj7dTHrF2Da36XQtMfRm2jzfZCGJIbr
qFzbkUnTsB6GASNP5duy7IhW0+MMBkTjZJudKN5/RxYzpYjzifAqIoC/YZYB
CVWqZsdetNq24OXy8zmItVV1mjpW8aMuEUIha231X9XmrNfR3ba3eBb+L8k2
hjw/UbX9A1dFHCEXaUBTJPujLHRcQCgHrBLVi2gSSm9hnvrUN+epR5p55wTj
tt1po/e4caajWAH3Xp3DxPAlSSMiaJz0c0F7hx0SlVJV5Lv41SUoln0x+aR4
vbzlnzXlcFDQMAYkQKG+83tJDjz8VUEnKC1tY8PmxUrVO4SN8hQVtPSI8BvO
3Zro8jmU6hnNHVDyOncED/WhE77dqXKitzkaYxOnp9OVTkmlFXIiDBZRQLUX
0n/fV+zmGAHgDveTmjE6xLtgm76aotngRBa+mvrrvrQD+751RIX4MCEzgyT9
Hh5ZSdU0/kGpx6locUZHU7CDKO13Wsa7nwNS28/++zBzXz05uR2kX0kF7cd1
1LAxc8JFl6+rcFPPTYRm3ukdRZ2iBxjAMm8kGXj/wzMRMeACP8faWk3y+Etp
IG5YVnUTaYm3aXd870C1UjJ1T5TaECZ9X9uejawYou5z4/B8EQEcBugvG4uH
GhQJ7LB9Hj5jy9tOwsKBA1cSmd72KZoLHnckx9Jn/hw8e6fMfrY8r1lPyE5b
MA54wM56QJqhjVBdB5ZSP5X67JgNx8gd6NDT0Nuf4lFgfjGkGY2OOvUQc+Sr
kJwQgh21n0xSw+8v21pPu1ZdJhui2cisyMLhxhV/ztvAuL0l/PgzrHHzaxcy
7+tzdiDQjJRxhY/pj47Uiz4xN/XbPYWXaL8prmJ2t4M6kk2gVs/+KpG3Pe/F
MZ8KJ8fB24kZ7UvOR043KKmNiJY=

`pragma protect end_protected
