// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
T8QeKFvoQmzp9KCK3nrEntTAyvQByln46vfrNZcRAvyimys3/543s7wkTsvK24Vk
BRGctsefJQ+ll1yIPFi0d5en/eYHFIPip9ohGY7ydJKqp8Tf7NGJV+yhD2Z2ysJg
lrx3wAVaiOdD+QX4J+tMMomSGMLnzE+h3aGW0vQeCBmTnIzuT2hAyQ==
//pragma protect end_key_block
//pragma protect digest_block
8L1UkojYeKzISXoqzCOjv5z9tmo=
//pragma protect end_digest_block
//pragma protect data_block
gmPgBalnyhVklG/A31remZYGAxiqtNr3Y0F7xYl4mPa/2TEeJlq1NapaBwuXGEju
eLLZ+YJc5KKM3Q+KJhfK+6/c0TfPfrMOL63sl3cW2JA9kTkeWwb1Sd7Z0eYtWHX1
4yUam/GLeBjmyeE/MBgwvjyAiNJCMs9ekNeKLAsJm77Qe7pmvBaiyCnu25/n54VK
sD6Ej2UXdO4RyQ3q4U/WJyuuSx1YzlpxRR/W4euOljaIoBRG8nqKY9sS0jRcCuu4
D+PxWNOCXqHJOzrd/3/ZqxBsSfTgE3h1RMdbl02X2RdJMumtb/xvLPii8XjfZs+l
SQqGHUCgZNgAV0mg4TC0nFREJeE7TE92VhFJhljE8L2kh9lMlqclsQXwVvrOuuvN
t/v/BE0bhArdRp+6TmN6wjWRVPOJXkpkGv9lteXb1d/HmHpcbtJDhTRCCwm3hVwd
Akxr0ZZx8LNG6O6a1zmpwvRKogLQwnJhTkvjjQvWeauAnDvsXRPR0elZa66VNPiL
6aGQKY90/cN/oVLrAESKjUK5WurWdzaxnV8AqNAJB7x8buWPYXXJClkSXw8rO7n4
PuiLDYc5P+4JeUspCBVklQk7Tg6kC2floFHufDzh/2tlNneyRBauOhFrakxvIJ5S
iWuY6iidJnA8h2rVTilzn6ZHhSo3n6FbmqLG2iOddNKFaGyJSP/ud2D0psmxZ+Po
WiFy6PXAEDIO7scJAB0Kx7i0xGZcpwZv5NbGxIryKH9hiwiHYYZp1kiR7BWef6KQ
ULC3Memgf8GK3NlIwA1Fpy/6l5fbaV7ksgkiXzbtI75W8ZgtKz2jUm3yepz0xtk0
iHSqSFXaEJU9jO6DfhU7JQeu/ca8XGbUOLvKIYFEoP15VDLWTFZk0niikGKtsFI4
iAs9mU8OvGLruMKrTj/duiBx8m/1gRgY15Vu1UTKajJPt8F7ILIlJDPpiuBQV1x9
ks7MRXp9SkU7/F3d0BXE6/knsKSJ0JDXwxgumGlSQjH4/CwYhAFFeJQlsLB9Amoa
adbWdcl/Si9KHFRRIRk5mSXU0l7nCBZeqeSf0fuNW3f94vr2FxTbhXJ76EuY5dt3
VhwegQfPUaQxDhabonSsIxqsNI9kk0Q08J12mFrmic30o8dsICriJrz5g6cOhY5V
SblifjfF5455oz1IOBDSlIk13pRZnZywjMs8lAtsVA4GbGgbZmwr2g7HovOe6pab
TvUKioBsMhTjyZmeDi3Ig5nJ5cOPBaCW1x7l2/cbZCgEkcdjjnjgz8Ii5MY74b9J
DP/T7QV2P+VwtnhWRMcgrgK+Y1lds/G6xHk08FGri/kVaCmZP4H0lIlZAIlFbiSt
DgFOqkfP9GVZxsud8Rct0HD/G88gPtSqYVVlfbxaQM+FRLImglkAOM+WhfiPpK6P
IlWwxCckPd2sVT/HwLfUP/i6EiKe/SIJF8RAazugRuNaV1e5+O91v8QQ1mY9GOqM
+1F+abAfxmdvCyKD4LxXf8Uq/+b1jTBMa5rN/EbApqdhf8fnT3+puvQ+J8jTM5Ka
vvRMtL30VRe8tx1VaFl9Gu0LR7lnWbqf/wy3mHMMlPIdNiRN9SCclllfvyXqCGcQ
nm0RQPEfzjELZW0IAiX1JJdLBDNBa5YvLY/R63xfnldrI8bi0aKE2TR8bQRH9YrX
Eu8cPzpghnxMvRZ5x5pqwYGJ7Kvt6uuziu06mgfRC0OIaZ4zkVxz/DmoJTgXCrCq
BS3DrojIpST520AnrGRAUMwirZnWgcrEB9Y6OMuOn3HIKlOpif3npGebU+kxqfkc
AjiM3gTmEBrdGZVYLtgwyRyLpDOTy6ST2HPBuNupUbwdgjrZZ9gofs1FwMNM/TmV
HvgQ4iHU4mj1hHKBIHcnH3toEZfFKLA+wbokbe38Xi2NsE+lnaiY3Zz9FGBnIYuG
aO+unIypTxLHzW6jXOUtUzn2lhI+ueBiBJRx3pF/ujZYwk+3wCpdZxJKSQFAmkYe
Ni/iiIFkVcLCqOgqkQmcKQVGuYxUH0rRHmBFBMlfKNXDx9C6JTRxDZAZr99S2vlC
MvMfPu0mWPzcE+KE3el4IYIhHwA4eXkm8RfTJ9roKcQzPWvky8FkhUpJ/tyM/01f
CTG0gJ570g8ocllF7pET1APOUqZ4QCypy3yiakYyJnoEI5pQxHGyATdv5OEZAHpY
lB19zOwfNw/l6/HmioaV22GixWY5UiTG7cw6ICYx5yn6S5gdT/gMiaKqyzulXkqz
ACo4JBjQLLwdALwWzrCmW7YUm+vYQqH0JaSaigePl5EWa/JHylw5PFB7yU0HtUAa
OwkoKssRBQaoQRWLBlonxhQnhkMYahM5oAlO0HDh4W+sTCaL7XH7e+2Mg0Q/QHae
ZYLJaImt6/J9sir0B2Y37gBcTdicCi/GDxfh7Vry/YmQtQP7aBXiKY0nzhU68aAc
6Hhsd7+LLTVsY5nquPKUy5EhXAUwMt9EzDk/suzTEd3tizfwrIHdR9Us6IrR8oae
8tNOpOTEgTkeL/6iAf/dWFh3uDEnYzN3G5XtdBjWWep/KtVz7Zl5B498aXyUn3O/
naxpS9cXTt+cHsVJDsySZY3P/OwNqfKbNNXcUQos0oFyJ6Tcbpwj6HzII/S7qUxe
ONPPrpjjsejtp/ElDqLg1iITayDEvWRsqYFLLOSlLeMENHVdAB2wIhMpcSd2dygp
OI9FdSUjzwqHKcCbiRFJpp6JTPwS8Mn8xzQugmD5JI4NkLUu4UovyRlj1sVI8f1Z
dZawgen7XBevFs6HM0LZbrSISW26yuPCImEalxGK73cnNGnMSPtzVOnzV6xfuxHQ
KrIfaWdMLx8MY97qmTzwwAzHgJyQNlczgkGRmvu6oor//6D1mfC/DM+wQuB9d6kF
Vr0FwTGWNQj/leghNRRkK31fVC2V1T+CYqeHtVG2vIO4bKIX4JfiHbkufVrdBy/A
tnIx60HeAyqzclZUK/lr+h62Yi1NxOXhDdZ5gd1EfY0tgqCh5q/1KQiaf3RQBLzD
4lAdXYn2hZrCH7wmARloUXeSIfYJ4zb34XH/abynZ3djHPvGv2aryCnd6g5h4PH+
MEhU46dnEcaONqeagDCBh+frRLpJwmEo8qWFwjPI0ZRZzn+3xPCgjLKJf4bYm+sj
McJFDx0DXvICVPIFrC9MXSC4Ya9Epo6J2lR6I4oyZVIp45n3AdOsuhgxpynoi5Sw
ki1Lpv21/e616+EcD8323BdXYsPNjVzNyIgoKTAdylzRKq3PzziyN8QpJjFcO++h
hUO1UqyaQB3PE4NOKADiAI5dQHPNulOJrYzK1e+VBGQUrkX6aLiPjdltQ4BjXlfO
eA4EZp87A2V2E7Z2icnpTqJOuLrXX8H2ew441ethz2zx2zNR4MiuWG9jNBiPJfwr
+ZN4Qt3tazq/svQCYZfyWIB69khqh+oTve8r4+wf1I5rXhutYpfVjTmY95QsbDOi
m5TrX05FcjNbMB0UcFLJeVO7iZNDLIcuBKyxM8InlVDc6YerpMnStjkD5sIOr3oQ
5BIOY8nuwqc/7nXmtfBNG1KOhYl/OxDGiLZJZ85+go/UF6Zo5A6ZvavTB65WnNfR
5mo2UF7krasrb3pNNoa38Lka8aeFfFQMt9scS4cEt+x+0Cpr4gaXS6nXFPRYiGy4
bgW24dPpp9cGxKH0xRBggEUyhY8hHwvnEz4ouoscyzGPKV7CnMAhs9pqibHffib7
ZHywwcUWdWbCFWGVfIIKmMMFu3twhm6gmSYGjNg7kxCeO6qQARy6GF+kU1ouhQLy
hfafyPTXn1tdXg9DJ3GKKqNTpvWAAiWYFHHfIFbGOcfad5L69m93J3yONaz3Rpd4
2IWUW0K+V5OhWWw9cdsHz83DkC8pm+kLucEuz1batTgh+s6LFJcZkHIvODpBHV6b
h3rJpiOoJBHXBfZCnUaAS3l3CG5fYtaGtw3w1HUB9/3ApJCdWAYdvNV/prMsvQDh
mjglpgER7JuNYYjnfR+lr1oyItmbTQ6BmwjIwmH58lQwwvKqXbZ7y1PzLnjL0rDO
IkUd1OGJjbraJXvg3vJXUw3v2DhGio02+Dlud2fQD85yGXCFmrXj5/1Ud93/QMpZ
9vwNKRB5li2jnbW9vjqVkT+PthWuzODCNSGI9m1UN0V9I0YYJ5F474QtNMXOGaD+
RL2BFSrmaQaIM7v2ZKN77JybAq6AzN6Mr9cSrl2w+UcANzoRBBR5ZwYOupJsWFLa
AT2awwDqkq4kac/RHlG9QM5Juzox2F1vVLk5iFz6YKVRlxNihuhyjU6Mg2ituO59
N1twGuN4jL56gAJ4kaxa9zq9lls41hb6/CMXy5b5HJlXCrIkHp189cNBlfMb3oSh
GQ7xvULGjgAaVaYJDeCkatPxBpbX4axISOsnnbSiCo11G3yLEZGhlRQP+JKw6Mu6
gJG7BW5dJVc5IBxP4QDs3KoiMRBaoacLljrTNqvN48dNjlc6ta2gg4l0qE0n0a25
aDmA3AivB6ilRw/GXI69vM+tv9ojb+ws+PaN8IpvY7C2cAO+G5TiFsOBpk+6UKXS
LcD/b+Mxv/ryCrRV2R4OKVOapYaM8LBtZPJSzHd7Ypkyk5tXpTOC0MuV09RU55wq
csdmdtu1s6U4HASUd2ibv2cc+JQ6FPrPPDlnjdEo/ppPuLv6cns8fF+ZiR9jA1VX
1+rr0wowCTta9H1mjDsPV8NlzxYBxRVMEDbkaL3w7yIXq56kqseHEscjWvUsq0M3
G5JpDGLXPR6VABhpABVqCC4Eftmn4IixoNS/bbhSzAAziiN/gr8gCjvCvBcpFb5J
Dp9I9eUgXBx11mvFHhVoL6rOQ5Z4lfICtvndwc7H+EzSHPloj8k1YjYEru6cjUr8
JeHpNTpMIuNxeHB19eXw6KEHZgsIbtIo9bCpNQKi4l3CvvX1EG1ndXhD5csjUUea
t7qggNEw0MsqFGbwWhhhPTKLiUKaURus+aYRXhki2TSVhChI74l+iWenFpG9C2fv
bmnUFML6J6kKHOI35J8A8F/Wwi66k2XKWMjYoMmgsP++Vt8jsrvXuPLs19JeUC1l
2dkwIR9CGNne2CXx6H0ktvRzCYUYmOmZ5hBgM759hsg/OZ5arfShAckdwVgV94yo
LRXRyZ1Ay3t/qCuoVnoyhWq8fzuf4L1wzw8LNm2bv1x5+mBHTROVTn8QhtWcq8zK
kvKqmrhdLw6iC0pw0m6fJk/W0pE5AUvRpGyBzg/j1Rd2OmWxa1jvVXkD0sQkMAVw
0JOQD8Eui/ZDa9EjJN3DopLJ7w5T60OAyaNZ9oie9dD3cEj1s1Q0T02BiGTrkRAC
SMS0m6cJKVdSxY7FIqmz97J/H/V1HsbL21DltL29a+C7DYo1X/mYwM9ucRqun5Ip
6UxPoYLg5B2eZpN+Gllnmm+Ge2q9nv4dCy8bWYO1O04YmijTGIbw4vuaDojkg0wo
vXGn4zjfcS9TLFxfB3NS+O/zLX15YDVBJcJLKJEzXeq++NKoSmHz4d5LIjT272Si
qU+yjefSXHT/nUwmtF/G4NjGCLpRQ6Ab7l6t3dUPF0nYpP9mewQrZ9eFwDnctbmY
z/z80f4VOty3+zdWYQmLKiKArY9fM4/TPk+jJnJwlC1/pvuCph6RUj9uLQ1OVi4F
8mFm+RT/YqcV5CK+41orxrkQZTeZv3E3WSN+GEc8HUrSkK4lJGNar66nt03prnaI
FLd90V/+GsJW3R6NPiylIwG1ByUWX9S15OkjCLjw2WGlYOxENxf9g5tWcmddIyRA
nJMI7BoAGflz6bSLktjcZNbFxOpFPtCRoSpKDMPFw6kt4DgRTULI20vAdBUsyLo/
U0oNXU1zsB3wwQ/gEX0xE+hxZKfE7Zm6/NDDxEdGUrFj1NsPSKoRzGLoF/761J7F
KqAgElUcVRUMGc/wY//qfORTayX9iBVBsS5cuDJnNpwMSQlCQfJUIqrqqqp9PEs2
FbP8Sr22czjuGStfEXKS2MC8UJhX/Vm9g+v+wl3YclsJ3KaJSUlDdCtCEgK+K/iY
6YhEoGstHhJ04ptKx/m95w7TceLW0jIVsa0HlHJSvhZxxBwhhycNVfCGPdrqC5A7
1xfJX3G1UG+sdPsTvmNU4copEZ8FMz/y544aeGos4DTWhuQNKQuX6k/w1+l7troQ
gBgO4kF+S/1oGJZcWHKBC3D/fAbxRnAkshi7vwB8AZ+/xUnJ3nAkam/CCIXkHVam
SbQRsyoWMqPaXcHaP0Q/JAcZ+RaY4cfN0IB1wa3MOAmZXbT0zgoLiwzCRvfrBn3O
FFgvIX5wCvbsucK01g1RPiezhnNrIGpc9pvJUuAPu6mdy8pnMfKLT0Q4vRwboOlH
97ZoMKx5Jfl10r96lWdRWrJ24nZcwUrf+Ge/+vtRVlKJMVANu+yCeMlLo2/ULDFR
0mdjeOVkSBo2FR/VN8Orc6GM/GrhX6/SDTQS8sMPoHtL9bsMI/S3qGWeki1NvuL2
tArKraBDW1mjxHdHrnx4IoE5M9x3HIkM9YCAvajdpaDhQYJRuMeRFJfaNub5GCSs
nZh1VEBAG/IrgEOnqdm7uh+wGb/PGDdVo5h4Ff6X44J3phvAFfzIYrjIdWPKQWAF
XIrefo1AhawU/1sMCqIXGWLdnBnNUcjWq0kXqqnKs1IjWUrtBHqh5j7La/fhc9FA
VZtyZdSmnujyEG0NIE5fAVxrrP0XxG+a0SQjcQLbR3p1hDF+qNI4DCFhLPUEzE3t
sXv0ut035dFodQB0vKPpyqGUusNuC+6waX4DyhtAQviKt74Tat4Ynl0+IFXJJ1lC
1E14D4xXcpzPiUWvFR9tCo3oUgFxkb8ackaCazfs53tdV0Ceqzaa2P06AthQ+nrq
U2vBOvTpaXExy3nw6aoBVGNHrcBFt7sSbuTWcDrLYhfg+MWrIB+6ltNxS6q0WIR9
zMzeusJOUHXCTylXKwhOm9tZuNnQlY/hDt2CMoAudCyl5wWFYu0uwpKWXkJ01LXJ
HbBDKPolFBjyetSnMm9U/MsvJNvXT9YOKls/WAgAKv1rhUizWgeLo8n6sCUkBCNK
W9T2HGZ4ikKmkwV4ROd6PyKLGgYPcYxC1N+DXsekM1mey7dGNwbNS4V85/We1NUn
zfw26/hbs66ywQVg/C6vcgu56boj1VV+ctGFVuBkkZIt5CWW5jmV4oOSMYBEsLwR
iImiXX8Ym07gCEjomPJ9kcxbCzsqIr0flUPsHSiefRqNF2zLSWtkkTVqaNt+mQGr
gSdSxpVtJf3NEgwBmcJbSafVsS4oqs932hbNEk6FkvT7sXGjmD0otZBhMe72OcwC
nkR4tMgTSY9rcitVLbmMlRd1vHcsCrHjIzV0GaV/98iS6qA704nO1jMEtM0nvKOS
8VUkztOOIQTw5kHylsq5d1Bd+LOqY5/xWWWpKELrrGVjPHD/9Az50O9tpoYWIbPj
xSvt0GIccDzD5wbBgj/a34Cb9fuZXdEYzrDsg2zbD2bNnk+gSjtmYfBqHRQfad39
wxL/KR/mIKHqJ4OQjAIFdfUwmFXJzB2zKPSTmXodqn4cbCMmSz+tdAabzjMChR5g
SJ7TN0MX900VGQM0oRaxXf8pjscGCgY4suMl1zyKm+nUfI7YxfEIqwULgk+9Dd9q
8qzJSBdXb88LKAtYVtAnLIDPJim3L2igVBzaRK0Xp0MhD+8ssT817ct8ht24R0y8
N3uJh5CSevu/B95wF+E1ciX654rO5opT4SKU736pAJwqLyW0+tD7sLNVmFXAgRz6
LnRRALZzpEEtpCkJ95XIZ41J6PThgBXj3qo7WHyEvrSJbQsnjOLpIYqzdXxjYjPj
4y1pfJn6tuSfQu2T1GSS15rv0ELExWNDS+4dJA/oRnRYM8xtz/t0i6M9morZnWAz
SX5fdvjW6+DGGgRnTqyVj6gbaP/yqtta0Dn6UrH3clNaAqUqN/ykitEmqJhmQ2OS
ogMC4665JtKukgiiiV07FBg7bgdCaUd1qsci4W8NK5u90C8Zn3IZgQ63s+uybHOX
iQ/LECU4SMAMBE3H52mKi2oaFORTjMkhG+b1GatF7aVGg3hcn2nCK4UZt/fIYJHC
dRKFkQHDdJ8PDfg2kSiA9AuzwmyYBSWcVplvCSv6OXkkfu7IO89ungn0ew8faCeF
z02AfFEGC9CyiB/ogyXC46q1mRcWMIaTsdNyNg+MhFrp4fwemx/CXmpGSS23bmqZ
TcrMUMKrFYk7acJhRDQvv21KV+TVZf07dcGjBITlJbz2CxY5FaKTFj7wW+ETf1Bm
Bwh4pfgNfMGqmeGqG7cqBZVsL+vSO6h9LG+Gbp/NnZGEaV/nYKad0Hub+YP45hNr
/kKwi32CYnCKfbWsvTlW5gZ7Tk5egDj1Hw/0bRf+lkfKNiJbBiOvBTGmyEfI3yvX
i8d4CFH8NM1/eAbCbHKIn7qP6KO9kgod/lpYQwIrjDioBweVC9MasW70qIiwfSce
bHIZXFb9URbNB7Ne0d2EZAtDCxDbyO1k1CJfZmEYNto5MnGQa8ezD2LJl68CowSi
zeNYm0CB8N0XpowdHpi9MSyOPauK/kqueXNSlg+AZeD70AAoPnzMLNX137dOvrsJ
vjSSJPJyUj2laNOHew0k0etwapUVKOC+oVhAjMgG0zYuxfJVwaRRSJRFo9be9ruP
Ffa32vptkPJ0+S+O/ScswboYa98oeVw5FLTAKkoehhxwejSOeNMAA3PjJZJkMyf+
o+uBfuM0dbkXCla9lv3FaoPkKes6ZFPDo//LDRdFsW7gaaD0IK0uOWVC9YqEv9tJ
ePvE4TUmWe+dYeWmqKTaouCqbYAsOdWQBCcGUaOUr81P6bW+BNw1ViTcpIWlZaxn
AexQSjmxFzE9dCWH9ARYx2EtVNmJ5nj8pLe5EskAQJwUvrNp+yQvLCaRPDlMqhEJ
PDX5h3NEVSyuxCMWE60uhmE9P80Wv3NarOMCcZX/DlF9f/Qc3cNoyaHA4cK1TljA
oiHBBsk3pYKXLrdMx9mftI+rCfh+g+xCk+dYZkzuQmzIR0h4pEijsL5xeEUzqDuY
pJj7tWvINio03Gs4g3u/aE4I4nA0fNKQlQWquglF+s8a4vv+S0gGK66TVBL3b/Uk
L3KBAyY2xvt/MRWFNkwZ9B7B7JUzsjlAnx8ilZDZrhJ1VdRQfp43+i97E2oIHvEm
cSrUEQzctlKursaptRnKbyECKxkXqet/FquL+U5nVroZXhiDA0HITrm44OV7yEhN
6/Bscgcp0aE9Q5MJOEFWiPBoHfvq4fB+i0qZ8YXoLavvWY33FKOFZpGo1ukXMGPz
CPwTEaTz0gB3tE7zazdOZAObXNJ2MNqvj4lM1MSqAFJOm4yVPQ7n892MoW3txTdl
SOQazppLZpMZnnZxYJxiQe01553JlroXXAy5JmXsJqv3x0i5xmzcaecX8yMfDE6C
5mNuhhy3jdHkfSQNXABKbZNloBLRNJvxxWF5aD/88vkaoLHHe2GR/gvNsRY7rNLL
kHa9uqaF6A4FrJYvip9Bk0r+0BEbV8ZIn3anEfcY0Cg1MTeOiqIj1BQwlOlUFO8n
XOP/q1EdRF7CRX5xhMJMXYK/VEmGcI55xl8nBjhmvMW3DYzP7ytoiFP6ZFOsa6lA
oD6JApKYorygCNpLVlRbIIiui9WxVN3qb0hWtD7VX6xKICqrikhAl9ZV7+zwTDXZ
Cq1BY9z5HsHxxooz1gcCDz8uR1Ix/bL8OAGRXmjFi/DLQWNM86TDSJEbZzpBrz0u
9QVNe4T6B1MGUp5SArAsDdpPezp+ID8KZuW80Kph34YTltKLUnvrs579TdtPnCma
UYbMd/IdCMlIc9841k1rzmXwzWFfFsBg4lzoIF1zKtXKuyQ1EbXx3dRmjQEhVbm7
oaXKRXPVeJiPXb81F5oK7cWbV0aSSNfxhONqUVQxLEY9MnY74r/RaY4w/o5RspLT
f2laFcTy55EjQ97Wc5fXigy5c3I8OieAnfd+C8aV1YQJ6etAEpGz+s2R3xMaVQWJ
SV5VKQ9/nIW8hUCkgBoRL0glUUhCdfIFhuK+jV2YdVuNOB6DLgs8qZQC0oI5/nQw
j65PRg1dEw133j6asSCBZVnt3R3qNmjA1Tsg4Cl5ADRF7unPZazJPhtFUAZzaMhg
veHPla0QFjYW4MxEVOpY8aWtIffwuBUZrbW4AwTeR1/QW2QpLPOBSq3DoyFKqnlz
iYOr36aRataYyqaZCJrbxGNmmcZEtQ+qtkRclx4tGvNMmKNdkXOjLmfO+Zf+xBVl
/WPkGn/ueBuoOigbyijIk3bscBgmrLOpwkpueG7IzoFmzyW7rxMYLhKChEpu0L5N
YMUYPPVDJaKWkX1YFVPTzhJ+VzvAIi5/pwsISjSRIs9DPCTx3Vvt6tnQOvSsI70o
fBrbrBtv/bNwqyEtwNu17rBt0n2WIOynJ69WDWbR7CKS0NL+9D19cv5sE9dZgvCu
fQwiRimTa67kGOqEy8TTJ1ZtpmFwjDKJbYz1avoRBXz7HOFaR1Y82bVVJht/CTb7
xB3CM7E8YzEm6md4HVrbahpOcdLRFzUIKeVRSuhVgJZAMAbf6z193JTGJg7GgRD+
thtLDt113JSE9yAbJ7DXCuwKh7eNhJpft6uaQanvf/pPUmnr8lCH2iQINS2rNZJb
fjRtdt+LwftkTLJK+mjplz+If3cFSqNePAASezA2ed+R/kGkS63fMzQ6ymNZWmaK
Je3taLIP2tHWinyQKDF1wcwUEdLWdVGaJtP1PE8KMyj8rvvwAw2Q96dqKtOji9Gb
i+ebgCsHF8lwm2Q+94Jwxjl7pfpDAvWpbNulNIINq293IDSDdXE2pI57Yt2Obg6F
H/UGJW4Q2N99UFqWE/cMlZ1YqQNy8aO2WbzhtyP9jpdCVE5u8n+6Vl+eHqX+fb3Z
nLdrWGuPagjxvX//vN1kWUUf1r3bKb7aCoIAwNI4QTrs7g2Vefh9X/08XFvwGA8S
A6heoVhuLpCehnP0KHdUw3H4R5w1hWrt30d9pUB5gn4mzQj5TiHb0HBNC+y/t3vD
/f3ie2KSDROzGpEcVOT6FetOmROvdmVUQzaQeksHTqkuRpgwXt0e9iEh363ffsX2
NwYlE9IVKljFaoMlqSh3Efkqx0PwTCW/7NIUKkMnBYgmi7r5oEVeiZsfiu4SR4Kv
8PKX4hMt4ZE9ScI2/Gp/1UNDHRcmXKfFFkzpsYq4MmCEJ0UUCR11t/haFs0TsegT
2ww6gcMDsYVTC/Ohtf6WKFXh8JDXzFxgN7/ZU/XEgy2FAxH0M9Ba13yIM5HDNyAC
LywR+f299TvG9Y9acNzVURsj1s0DaBv28XvH+ShxTvxrpNVnoAJJv5PeoYpWjTvh
HADqFkNzBJma4F9g6kLus9dzOuvioKZjHfgiEsNypmVk0MpelodKnC8pmv9j62jE
Awppq1/lYE0ICoKi1E76p9uo9K02nK+poMWGmFeekbrAf12Dc81L56BJTH383cFm
i3KuVqWln4bOco1dEM9Yp4LG1Key9KwMMD5NsthSnMyQx3CD9KsxHAaXua6ZBVi7
3JwV1iKcxLl0xdZFZEVv6c1phj20k7wzmHh9G5qA5N4hkDHsWN/sqzSJ3QQjlOyB
d5UAs/7BbQw0hmig3J3vVVkQoUrRS5yxZR9fuTVps0J7KiMVM1rT299ZxxRI74nZ
NvooH8CSmSgpgbmmKkMvnW3nsfLpts43zHvIJsCaCIG1QVOeQuFz4tESGyHRL7iX
pVVG+Lv/BKkSmxHAPil/NMgFTEV4gW//PWL+4kvhbCO7tOqvihDoUgQiXpGvm1Hq
xdwcozcW2j0rQG7dhfboFFhIabLTtz6jNSDqnhuTrqJztk0/kmBWbgGFEZlLqJ7n
AGM/l6LEL0oY2A/hZ1s7XO2iF2KGhYaTAl9bkWnRMaEbnl3FqBMroS3ycoookbgX
lbg0w5gOlmoxAn5G96WSfvbMZhgH8UxzTqEdHiyeLib8FnZ/doPLPbU1gCEM5jTH
zMFQ3Md7Ry8KtWFctpkMlqd3brFYTxfnHjLIF8RLA9UCeL1Mu6TW2cFpeqfNt66m
KeMfgmGRT38CnuuU1gD7vhFnuBXpkUgIUlpytftFI2jX+QJVZJkJqeceEhPKaw1G
ab8jsfPNK8czs84IqLmaNn92zaDwUKdfuEAyHsKPaefhOYiyoqXBAMDiFi1eDAlN
u/IKQ3r+AcH4om1fX4Uqq73EbV5Kn4yQZy+Rf0yVkegsrJPvejbT+MnF1ZWqxlT9
51kdElO463iC5cn1N7goo5h5B/2+eMO+6col3O32RVsWSi55CWYeMTJB2csQtxYM
BAwH2qsPr2z4JowyCYWVTpIvkfM7KZxSVj4nlvYTgb3eE3dFjh0hrDvLSG0Sfv8C
QTu4t2kpqlGgI8EMXrjtCPX7+pBL+LFa7b539uCi8fKwMSyWUIyXGF5Pkb7vbdxH
6P8RLH9pHVRp/xkJYqDEoYuuQnh/g1EFOvCA4sWnQBh1SgOgYGukOD6tFEeTZbNR
JRRxsh1/ueSMsBKmEbMozT4KciuASVFD16sIFRZFOMKiDuY4aEjCjI6ENpiKNbcn
DFJ8byeh6tGDxQmbdhQsMcUk/Az8Un+fXHLkd2nl71FnL68EnGA596eeKklCTmHX
N7UC1BW6cypvhEqMw82Z2YOZMB5fkOdz2JFteBabocN49EbSKKfQgPYFkV0DR3U+
3ldfU3YyCiK5pnMYYsCwg11YIjas6Ml6cZR3j5GPuWNANjrad4uDs0Lrb1kttvXb
AtND9+W3pXZjIxSu1MSgwiO6DN8BJDiwZw9gl84EySP4rH+nsZOakBC+yX2LmNlU
8bUIX8kGNSic9mTOO+CpjcsqPzjLCupoBejlR6hwn8W1njOhzD+Np8zoeRXAMorm
jrCm9sPHqQtUEBM6TM6FEoRDdMc0HsT1+XCuQ5VPHPXgTgRlEb7Fl2xZpG/P/xZ3
Fzsvvup7XYzJHI9RZOqFl87Qv66XwCbZxVpgg9PGwP5lMj5Veo8eOrFS7KoeBzEZ
Evr8/ub6TW+zeglKpuwaCzT1OObN9ksxFV0k0alaX+qK+g7AhdhYA42u6vmrriZN
ScuCeTxRAyW5/yf+lnSMZQTv1NwaP27ztp1asNkT/qtogQmudNW0fEPqHwUgf6uh
LhTMaAR2JHoPPejsGsJLkkuAQ/vA1/iGbIFy4GFjnsDIvckgElE3IvrP6DtIM4bI
nR7JTRPzubAiPGSMNp55/E5PuUwl2sl72OVLyadyr48MN7pyBc69KD9nx/u/YnuW
UHrleB/f9rcKo66J2roGQbIDpnsktRKmOPcvVUtjAlJgbxoZS0tarjMlAzfBbtuX
g+lTl+lKOKLT3yxhCpcoENtVFwmnzQXWekPM2dUdQYujbNptS91WLI6mv4H+dcz8
YvJe1HPFM8e8nO1cQSwJu3SB8bi1kOgVjVRmfwjTJPUR0z8vmoEEcL4il0ntZlK0
pX04hhIyhgo5RpYMDrElbtzkXTo7cqBLsdAPgu7J7vOcyvAoJBc7XJe5x9TtfVlK
nMChqUuSpXy8PmJE6o2f0VRNR1t1tf4Z1G7iagNQULrbJjVYCd+Fw/WbQmWVhxxb
AwCaE4bBG8ggXqHI2noD37zQSiYaz+zhrSkvsHgvGypERb3hXtlWlwIM5dgIpiZ0
Mv9DpQ/SuxLN2yvzHVujlSvWPP03cCQOtcJFalWLFIbZR0/i6F14h//3ki4KKhIZ
Yjx1knzsSg4ZxNImozxTfvnu+I0NSuPHjquHzJktRnPJl7ck1Q4Cf4gvWX07nviw
U8XD3gCsG1/se29WT8xPviGPGQxgY4IL2eIitSg0dsGDSpV3fuJ51vcw+s7r5nJQ
KYCTDU9MiOn0H9ilcS0kXAobTKfSTRFyaUVYQqvn2Kd0ari1+/SEWQ1k40IxxOUv
Nyr4ykUerat50cMbmg+vwibPQ9EdF8xmdoYG6N/kAqe/C9ulR8nVlk9WDPEv9V37
G76KG0xG5hvTZ4nf1QcaO2wzYEn2r46137ScVPflMg1mH1RdYmMn+z6LGyAq1BEb
VvM6t10iTov0oTGsz6lpkwOf6LWKyUoKlduFeSMyd8YDzrflMtGZB+8Y1dgELJQo
EpzhqrE0vF37FBPEzwyJU9bu01jJVLNDLFSeEv6Hck+/ulNaI9N5wpeDyHaQ2rrQ
A7MmsK5m1f83SyFPnrunIOGg29ekifCu+O6XvNxns+2YhjU2YOsoXGkCcodvx6mC
IFiNVY/7zK5il7n0iVrN7afTqP2SUnZPe1hluzFP5fC/hn0bm5FHD+QbImzqw00H
9q21z03oNOM9fvv3fziEBfNiOg4cjhq8QPKi6iF4eAVVYnrcvNXWZzOs/eWJIRXS
6leM/nx7dEqFTPtQGE9XThJ3w1MMFCfzFJbhaHEHxkn4iCvLNN6r6GLMMdLPDwWw
haW19qfROXU3H8qn45i74XAIBvJZn7tYHG9u4CLi/N3kgwSt0fRM1HzOr857JQrv
3c/74+tpkJGMRn50q8PkQp3KxrNI0lHZkQvDE75/+5rVqoD335MEuFWmMPNl8KiM
ojci/p4l4O2QElVo4qoJ45oflGw5OVpc03NVhj5T/r/H2giF3q5ZQavVUb7kUSot
KPAT0OsbW9VvYE+MRa0KGvKiOSSGQQoVjnUNO1NpoaE0HGW9PHqtv7X16ZBa1hp9
frIrvpLYU6zfGMgl1GoUl18qg5hFtxqAc6ByWuqgW7ycrAHW19BkLC3kzBu4kd3C
y+JFKecJ38mPy11vXwwyUwSPfJtjbLLfo6u4+H+w7ZI9kj3oB6M2VMrY2cgBnZ2z
Z1qz3/FVXmlm1sMGTy6MONNuolJg11HN2b6y8VnUxQ1bf02/htLAUn8sGNff8rxZ
qd9HA4O90fje5pzEM8JryAqQ4JJsZZRrkh0edAzc4Oh2/H+KjS1oS8VlTdgYbUsk
igNa3g95UuUI83cbKi97QHxHfIZMFewRMt5uQjmPPY2cgDAIInmUckLJ2h090DnU
W7A10PwXg/jPNgwuodw3J8kLSSspq1dySlX83KHu+IUpnW4NRVXpJ/BLHp6f3m3N
TyTn/nBSkX6Y8q9BL3Ex1Wo85Mm6i9QWubB1UUQZoChmiHaNIpLjQ4tH+U/HcK8A
zuoTceR7syZ5wBRGXa293hRcwUXqM5tiXglnbmJCoz85ENHKBAUgju4auH0fsJvj
2Ty5ksP/TGUo9DYEKlHkkoc3t61NJ30Qg78Pbr18IHJPtgcb7yXMjgJXH2A4RRbp
UOL+WRRqoR6GEOoePvmSEe2jCyXurMmPFnYBYDSh2J8EBfIiBKIrxKkmswTpLLJh
Oe1UurXzFImDvj3Jd05M2rlTdl8v8AsndAfSWbnqxNF+xQuzW+Gozx1545YQe5SK
iYSAy7SYWU2sU0YSOY91WcCCi7bbFKKFSeVes2pr8GcAvRMh6/Y/jkw1fKEpYf84
qLYmI8p8kW5gSLo5bc6N/LFm9MkZFeP9c/EMuHkN0Y8Vo87Ezv4K1GwxmAEfiRWd
tn/cW3Tf3ZnrPV1nkltLUFpiG33B13YbuJo5o+Ab1ASzXy5AYEJYEGs/JWOdbw6P
YyI/60RCJeDXKzF8yQevaAz+DHBi83+dI4r9vKPnXUW0CoyyrnQOEiLRTnSEudgw
DGJ+4SZuBm5TAiWshdnKU//izbi8bckPtBpSz2DBorgBFkWMk302USHOiL2vZHp0
ZlkViaOdRxf+UaSCHbvUj1enZ1O1suxEW7+58XltCdXabobCuizNq1ZPYI3DPjGc
17LwM5/by6aEdB7qnahRLR9ZlVBCqGIGk0NkkhWweo3kTDQniaii0OiEOUb3Yv4b
yAMUBBpVKwMljsOW3PkQ4cR8iClEh3d7uOZOlVQKPp0NjUPQwBPacoa5fI/1NKzP
Tg0BwW5EhgVx7kND05ZEx95GNOw6avYB04HbofW3R7FUciw4QW+N6RodVphNliwL
RxVqGFarfj+6bXrM2CplwH47VWlmcYuz6E7rQufKroQQUoIK0EefD/Iif+/FFHmp
kuv0wSgPe44y9cUwyD062aZuwVv5L0VS6TS3uixDV9fYTLio2khdKX2Ir+cbc8rQ
v3kTDjhcFy9hgODn5Ncyy2uSTmLqfNjw8dcV1Vyo39+xuzGM3QK6RNIDhPtHF6Xt
RIt+K9GA6lkqEmM9Nzp4cXKEdmzqqlStvqOqNRqcw5fTp0KNyalZsYECf+sIJ3ds
0GNeyfTRbAdz7ivGo1mxjDYjGMO8P/UI7r0HtYpxgI+BCEuf1ySlP+H8c4yQ6Aa7
r+NCCCFzh0DFdwe0biHSo9bFG8zct8PnstADtMKjtiZqaDAY+fi4FDiyNfgiqmbW
ju1nnrAA3r2HNnib5d2kyTnVP9MQtxzAlxkNjfgG2NoPeq1OJHvQKtubRXFYmy0B
utklNfLfIZpT7OOOBLDnXTyrN1/Lg0iegIHWFnfpeOc2TA07MgcPva8MJOxP1byB
Po4GO84vX5/RBrFr5hPabQmk5ZO6w+NO/cumFVlg4NxEPcjV6Te+Y7XlaNAgRzjL
UnR7e8eYXeVn5tQawulf7hsm99wivHoPy+ABDn19HyjLXIDeuGZUaGRPWZMc3BOf
tE71UNgi3JkFO2xm1sosFDiwYMH/4gyk0r/yjE2ZDWGTKymfqZP7wqKccdtd7B+2
OweAIe0i+SCgIwEe/aYwx7DKcnnr0VKIldeBpmaZPav5EWaIFy9StNue4dnMfapv
giqmljgPu2vM+lPYW/YGX8jJdi50OJft1qlSstUlUwGBnxAJVZKgZesa8QBKhwEc
Jm2Anoced5gInjrBYdBq+05ZdwJj3pYLZ2pWSUoCeXoRjNaMg9Gm3DBcbkiZ+V1F
1pdAitGd79zQ8wyL8J4sl3DS7615ICb46CA01gA4H0Fbu03f96EanAMs3r5x9zt6
qI6/yvX4nww6/lGMP6NTcXCgGXXXELfEeQI/4xvGSjUwNZSNj0D1/iQeumMTObLf
8UNwbx+Ev1ypVn7ps4T6DxCSpPscRHQLmZsuA0vvSaPoPDuhDvShyjjXR23TZj9R
GfsGB0ZF6EYVXluYAH6E36/lqZUehXt0uemfV01reJvZxZ6mTIDsf9mv21bz59Ne
QpTRlUqIL42H4MyKtYAXzQMK6MmwAjaA6QcL3ugpXlwI7Y0T07NAT2QFlTylr3BN
LcfKA2jkirUEfw9MYOgaSatnGF+Bx47IuHNoR9M1jEKBQCDd7wUYPBEQxKIhMAVn
JMHlqN+vWlOk4znMExbr/SC8jW5PUOuvw8jV2goy4y63k16EnG3T34uyK9X0Rnrz
PEbtxpu8RdI27UobuwQCe0mpZy/63TyzJU/N7RV+5cn71NquDq3d6wVWZdkswqjK
wSdSZEnCLS7g39BKCi1XGPIhWVOrbgbI/39B1UaZ0AXFLaxYUCH1F4891ZFFqcLi
fJdMuBokcZkJ/iKZq4rXr/aAIzrzn///AZxIum5XV02SnjkFu+10BKl+V0ktaM+G
ahVb8dclqxuDaxyv6ZH2ow/3YkK1CCcLnmh7/HxUVAMPL2uhc2o6xOLWLabOPFIF
XJ0exM/G5gqil3JKTKVKjkVVVkH75NkAlSy8Qbyj7wQj7MbjuF1C2FxbkyaHnIOZ
5bS3gpdgK6bJ0eGvl6RyE/+1bFc12wrQv60iH4bM0C+ayKbdffHXGIP+8XyMMSQW
kTaAhqQ+MiWheG0Oclqykv0vQ7892DkJyxgy2jfxRdqEfUB9Yns+bWMo819mRMkc
DAOPGAWj9ELH7yq8W7yKc65fRDxxZBvZWu/bzFNvGE4YrIGjHWPJGNhCl13Lpke5
q1Wy+yYYBtguArC2QJQ/vpUz4ACKwBfblSDqwmUYT7U5jj3RSHgFaZay+jOea5mx
tpicFGofZmppnuSV0J9dHaDIDK18Lpx6xviHBmt69EYmJcGM+pNMdBmVSWymJrZF
vW3qS6UxZeU2F0WuJv1bJVSOKAUIvBt0sS3xpHd9k5jQIPo57hAlX2K0Ocj6eoDt
YegfE7pO9/36PwgYjW4TdsSj8RsD5SzrwTsD5CBhEUWLDvNu6scb7ja8WiEglUi8
8LK3g5yOYRUAmP4HjVAmGxtyH0mtBXJTFBSTzqBNkFgIVc3lcB7DuMY67nE/EvJF
ElSmbGxxacnR/YYI9c22s7mg4lRnPlIhVw7N+F01GBhAuUC6cRU+T8wYXozdYOY8
EWDuuTFz5/6Va/Ug0TMAB8/Qq+0lTujdBvmeYd4KgG/lT84bNHWKi+p5xaC/Rsrm
uJjddsW91pTg8xTwcmr3LGkPQRb7b1Gh6PEqYyDlT5Rw2eRRCnGvcMK6i20leHeV
gZTs8WZ1pw7fSWnrli4rWW017Kn/H18//qyOvrpn58dhJbH0vq4+9cCMoU9TeAYJ
fjg/PxO11ZMSbR7+R1lBiJzhq7da7LZl0/DabNuUPCrth8RIYak86bRFaLHyKkbA
XOV5QCTDsUU28upCDAGWTV2IZbG/88IOg0/U/ZF19qz6dfVmQbwYmrIq+P9A+yNu
B9DPIRivjBSfuFM877uzr3xvyEuIU4g2Fii3QL9oO2mk9ayZw3duz4PcobWKYWeo
7taWNMe4zghXnXFuCDU8gV1zK8ttrDv8I9UYldOHp6Fxt6I+wtXLrkQNc6ZHfw1y
YCLGI/J1kjXKfKbMJfENqBVexXLkiTNjw+lf1Frwcw8R1sPFJPQpZ/r0nF2hJJtD
TREYabgO+S0bi4fBiKS8vVODuoXrOmv7bvhhsDBVggqCRBW6IlndojvyyUR/0KfW
txbQAL/s39nm38yw+JNj5+3A0FZdpdSUMsGAv2Fyxov93ex2WC67nxr8cvNhbysU
AU5w50k7TKyatzovenLku5lm9X65xk7gI/zIRA1+bP4f/JrV16wBDDuwnNDrGMUY
JKM7t/IudcmYYsTs5CmU2JUnSIOWYVE5Jxwv6M7fN02Y0PJTeVsqBDLkOrMKzX5f
etToqqABYd+fqJdfkOP4mKYi308wLn7spfibUBlloSMu8uZA6LdUslZXiy2R071P
NngUSDqGscFZLkxz9wDUIA+RxJHPQMZzh3HJgy6UqYCfcPTrDcoF6GFcm9HN4AXz
woH/V7yluJPEC1zOObguFncfhCW0pefvnpcmD5AMiW+6TEGbbDL0nEtMSGapcp66
hEnOz5JMCdqQfdFDAjdmMKuNLKFjNN/zxN62QUk2qeGhDtz+vaqvf2qVSW94xfCU
D9NR5GX7TOCLMG5sOVDVSKZRoWcv6DD0LlAcJ0FON/eq4G/sI4nsRvL4xS5j5GHF
zGFLF7zn+o6SCQsO2p0VegnRhpSz/PbGzlaVrtCoRSfhusIuBZsn3PBGyS9ioHBO
polQ4PS+GaWRVrMRFY4IzFpdyqUwDvhlaeQCL8J8FHt+KpXodpJGPjkDbZleb2e4
G0Gfzp8L6UymQ7U/eHlKj01gv2T0SFEoDqXHhMPRAYQIvpM+mm9Y8Lt4ypuXY5cO
sfHZWQ+k75pnHsK9tgVwm9wC8fBnrVgOX8hrrqqqtltNJQCA6OYtRYmZyiNxMfGv
gSfSvTtHcz/xCmqQlW69svBzbUOlX0IGRunZ+o27kaxooUgSDWT6P4TnBURNDcb9
oc4eJDFtt0ucnhPTCkvsoJI/nY5yV+Xz239QjLndvBVQe7cOQus8EpQKydWjbjZs
uuRBe1/NZbApybDt6hImGRkUaf5Na8WkKRIDNZAgih1zCeHT3Yav0NYYdnI9fW9R
vjSMfuA6lAI7XUz4JMvL5qw+UCFFvU1TffRQUckDxghENdUAwiHCcnu0DKeK8f4e
oH2WXnMQWtUYICZZgXj09vcegeFsI5oYkddUyuBNAduIgDdpgXLaOKvdWW4PoAX/
Tdnx6Bwe46FagUS9ZpYEO/v75b9suw8YoFUikv3wT+q0rAZDP2blA7rsO5z13HGi
jH79cJtvrEwX3vdI0VxbgtsTNr2etw7PKzziCGHqsp9YzN126paLhuCaqOnWlAKs
+XoAMO4TklG0yNuMXfC6HEYFtp6usScTCCboUiGpIkLuviegRQpxCvdmB5nW1Og/
tTbJic5P8NCHOdMW9pS/xsl/qXORVFf/pCLIi8+xpEntBOqhmBpG47/MC8kjeXz6
q2Yf2PDvIPkDXdhEKyhcFoWY2ZzCHatDRk07YOz5pD3rdlO/47Mz9o5qvg0Uay34
6dYoPTHM14kPmJCyCNtVm136uta0a+ZoI+Qfxm7sLoYdidH83QjJHlVdk0M0MvXn
/1mM0lMp9XtIwY3DC5GkWcXlbEJmC5mx2jBsr3BWyzZcF5nJ1RwyOnGopMHA90Kr
c9YLjbA7Fm06hhsAG8WUgnoTb11fVvYlREVyMeDpQ3h6sKt0FhCk9TOXbsvraLHk
VGEmMnn86G5FsWg1GfBxxW9bAD3orXZmZCxBm+lyRC3+QhtT72gw9UdOAr0D5rO2
mvk8ogTVWBhT+qr6nlfDoBIvpgDdcnxzq99O3NTBQqHWxi8vwx7O1oeE4w7hg/cV
nXmXPQXNsc6gaQvlyBPXBpqZv+qcq+XHorQHscQ73VJtrP7qy+oiJd/1mBYZdbv6
GP3ev3Wmrr8jH6qEuUCM0CHKcAEAXA3yTYr5XalhNPmiwMcpm5sGjNi33hggybj2
2TErDPaUWBaM8ifABIyuXHdPIsoLLT+L15pDlf7/lWjWUSxE4xsyA5Ml2Fll+JnC
t/pcsKXP/Btgy1jZszZcNq5lssPzCBPk0qKbTL8QSOnoFMuvyU9YY79iQQuYWULr
FqFFC6Jx40mbHBoRckKp6cAWAE+sCcHvZYTAZVuydkm9aOaYu251EeLx2enUuBuC
nL8lKIvb+JvB+n6YiXGomUlqIVWJASD5fyK5NNuWy2qw1I7SquVYlXUxq7zRWMtm
XcfQuF/ouYv5Wdg8t4b0Ea5SNypCxOiIu25oa96OWywi8zLJPpL7nEMFWT7PWN4j
Olg1NI1nuNMegQkPSr5OEGlFascvuKnIaTfn2tj0rTXeSQ+Af+OTqxurrliYxI9b
7ogpCwy+CWqU3R9NAQ+hwVUgLV4XshFkSc3Pfqt93VZYLMikl4nTEZddlW/z+Aoq
dxB8H6CsMvYhGj63apBp21RSQfZH79PGz1R6STTfm/ynDUAcx3FfnMuTHTmVkbaD
3SU9Lnm9ql4bixVgpyzQrAfvKu7kPOh1jW8JyB5vcKKY6AsE0ZU/lmat58owzZkK
k9QLfvof0FOx9hgTIyUFfsOkAz2yaT6tdVf4SgqXxLCgqtaiyNn/jpeFGEDAHmdO
taQ9a58PKSL5vjX4ndtq6gOQGGuyfD4JbawRrgKJ/G5pEuL6TdO5mUMfjGXVgaAq
UIchod2uky6miIaiiosxDCSALs+cDGpTmLeJqd0CBMddgx2CZnJDVceCwbxOCiAq
lwiPzoGUht3DUkVo67Azi5Vz2P8HKCBbKIOHu7V36fhAxSOATIl8F0yX6daRpUyb
z9nz4YLkoSODFQTeoin43V6seg8W2XI/njg4bsu2GgOwi0l0efVNG+YBkncvp8JB
sKwPHXRZGqbVV9gU5pNShXB5W2RPwgKDTK6yU7yEpO84/lkQLDMkGLlHZtGBwsvV
qUBT4bp1LekoUOSrQDFGfMR8MZLiW6C83Ls1Hgq4mYNRWFbu27l/WNTnQFrjxqPH
is/Tswiub5VQfnAVI9TdFyFK9Tgd0X0IKxNHKdiUWwop17+1RzyvqmQ3QHBuGrD0
i7EmxwXASrizFHi9AOv5oAqAcA4Trv4KrNOKDeKOUOraVyVBDqtefJEjNctOsSnA
OAuJ9Up6gY//ROqT3etvMziVZO+RRZceqy28GhVOPfXLr8Amzy7o18kt4K+x6wcX
M5c16ypRuYRVtLXquZtgC5hDMMofmHDZTpr2XJyo74P3u5JBUtxfcNIfBQEfhoPd
uhJuMH8cgmI2kLP5Rac6Vo8BejhSaKhrzSV9ffTq5KlC1Rt8jSLXy/rhjf8ptMVZ
MVFGRJ0c9jwZiQ7EPmbDRNUSIfG3MLSztgozy4dVxQ/Aena7dUwMshySSWBa+FAA
7Ucqktx6kpC+d+5acKW4i1GK7FQbGcXc+uGhmt9gXLMsiVz5MzllGpbBxFR/hOYW
7kd0IuvGjfEysFkmSzf3SCeFddLLJ9eFQhHWAzpSa4kwe667suvs6hJ+5jzfi/BR
dI9FzTBuQC6v9aAnQQd0Boi7BkFXTRpOGu0zahAUmaXFh193v5SL1jLwvQhWmOfR
9Mi9rEt6Qhk0dWUNa/sHpysnxHatBXl1GYTDXZWlfWS/W+po/tYTAYpJGStOOorX
XYRcIZP6zAePdrrKmeKUE6dczZQS+yB8Bq/vtZ/Dtps24NWKok+DtFYg2V6mQxIm
BWwK79uR0RWqOSAy6sVJUOQTQLcKNzHe2888pRAvE+hM/cdRO4WKBgiH5EzW4A90
SSFxV3/slMYSqks+Qf6uoIR5ksN1Pwl9o9VSGnWNGanSaS5RxJaKHFIhecpGlL2l
XmgCzuLcLFagd1+hesgmYRwqvRLuQST82T2wT/W+tXkNHtxWdWz0EuMUU2RSbqwv
pJk1+FJXl3rpMY5FFbTt3Yb8wA1AdkR+kiKRj8KyHqTCrGGKFwkOg49DaZvNKDac
QS047w1xt+6v2RCtQWHgO6i3B/Rzck8GaPMZWtr+tV/ehNANCTo+z10bVMCsG4oJ
aKv1hSGByb/cnwAHMcOc04LAZOJCE6pXu1aJAno/MiWHyRR9cJAtn8vSss7kp/l0
AV4ngOtIifd/KKa2DCwne29MlbeykgX1lfAJkDBsYEoVCCGxb9+SdFpl2Tmi8Gn+
M84aNR0yshJkjWmrCHGFYpsaxGdJr34pPWwErOEXIfbq04l9z6IgqI6oUl21lm90
b1ZIRZKdXZQzVQtJep2qDsUI4m8bjtzBpF+czeWjZ9KEopXILgXSyhFJ2NbwSzLr
uJzaoik5w/ufpT8gO4yChOeb6n7HhvWfsSyuwBQoKWcWDirK7tMhALWu7lip9+vW
aauQeW/SiJTdmyT6eQh4+9e9+Rn2YEQ0GMlASqktoicmH2ITXzrh4FLkGO16AgJL
IvZWTapsAgTFKOJk/0oQjxwajdZNQvDwY5ExrFDVg0mgYfAy8rGTFnaliX48905y
K18ostVzZPunj/IRs/4a1t34ilR5YImyaTVLgdTOG879Mx7EoMwl3ToQu0MXaLdR
j8O2lQ9gUZlHt+VzWtcVg/K8Edm83MWaM6FnQFdvp+KiDjuZmvA7X4LHiHKnVRLR
/7pj7AioywxD5MouJoedrLG+LPr0Gw8NIIcfzarV9tyI15zT4k/b4E/Mwegj05MT
09C/5KPow/i8ZFq4RGkzOeNGX1RjeNNpAwRUawnflbJOuFi6yu3FeJupDtX2QST1
WwZsjdjtSE9V5rjXVYRhqzpeK87vPJ/OuuyJxz6p5LePhzZtYft+kkQVay6l3E7u
3ySKBwjB9QMMXH+Sq+iNtGqSza1zWDsgdjl8TxZsi1bivsO9QvQBh7Rb8vdoBCI2
602NmJ4/qOXhZb+yHF0MEJMlQZYQCbQhwzDWrguDe0QvDhNXVPaWgpq20zE6gi+L
hewlhJS3yJKbqKvTxbWJ+kfkiCpoHvg1tRdrnx/ri+YGANqDLlqSMKXTUiyFysjM
hAGXl/Gk/B76TC3fCTeby4rX6zazK74IlGrDIDwxBxNTlIxUUIjDZAb4rkoAl7V3
orHD6deqJgjDgxBmFnlqn4HDTi7ws/6NYDUB7Hy7XiE3JP7rS1kNwFp0n+pnR5x/
oCmHMsk2nhO+UyyvR2iu9smEXSfCPLnSfMVNhgB2yzEuoyYEzF1iSkJ0jOGtndwq
BLhyic0CTCWKn48+RDVinSB8niEksv1nWXubIlTHMl4s7CbNRE+UF1pqBIp7no2O
pFDo3QcyeAXrZ/mF7pFC5J+RADqCdRpArOvm8IPOW8MO47jq1hD1vGoZUMTL+shd
ZzMDFQDgK9WFPNU6hcOrC5KupkunWkzK58JDmPHYzI7hszQi2Xm6Nqlpa5twC+Lv
v/EX8TfyqRCakK43RWTS9VM2c4ygbRoF5dpR01s8NV4YrxxBWKS/KPkLiPFPCgQ+
6fr6DNJ8Hnr56Ccky2b6C3W9Ze56/6NPT7A0ruxCscwky3eDNDOjVrg8wsg8oSgO
mCPwwRVqvvmCL9ryWMccAk8zbh5pBtqXL1SyTqr1LtygM2Jt3aaK2FSC9RIkm9cd
3ofnh+qf735TgBeCqvkLyveRfAUhMN1v9IaZIjfTD4CCnstH2lvtsKEFVRe0JbOv
GSk7AWHKcfVguOtpzHFBzIKc96zsXYGOAiae+DDM+nVme4CzHxYI9W8nnbe9Pu7P
Lt9RjfwgM1m3wtWJybVAoS44ecnPOC7TItvDvuUFpU8PeRd7pxtPoRC92bS7uZVG
4g1piEmQifri79+vzf4W2oImOIeNzFim5iO7aHZBfO5UMIMwHtJ2Ae9lyBDfQwfm
L6ZLaBcLl4gs3XJ9hJB+YylTW890oJohxROPnJS9n0Z5eYogS21MVibkXdhgamt/
5hrGUprC0hwmpsp7wtiUemnomPHtK9y7iJPqbj157kn+NMYQ92+s+FNx8ixrlDim
brw0IVJWsiWzX8qy3GkahTkrTHRMxP1YSAH/uqPmROspgJcrQQaCDYKdRUt/tajd
HPlmadaQUyCq/Iz9OhJWmaFgclQnyV6HdHCdlEb2rr1byzms0wKExK4jGhiGLpXf
Ha84Ge54MtQxfshLR3hIRmHQmu7IuaO6Z6S40HCSZbMV8FXbJyE8UZkmKV28HUk9
ze+Bvu5adepBXvns3Sm3rPk+e+mvPlYIOSroLFvqEX1fUH6HLIj7Jryk9+0AUqaE
/LAlw4azb1nEQWlQi4Z7KUNmmFIE/7uPwnuSLMyJAZ0uyf1q/fV9moH1+cYC3YYL
MfPSsA45OC+fvX1tFKpFINL/a+QOOw2BYWiMGktIvMF4FGClDmuxkyVgZseN2DZk
HqBZIj2IjdIeW9TSLXZl5wCD9kwV5YYh0lder1JFmR5lhQmVz/xfiaQpJ6msAb26
IRHM4qMNKYYhtJISQ7cc3FYmcEzUAHZKkqjQNcHWVZyID5tjI8NAAZaDBUEHA1wZ
NVMW0KSyYfcUiHkIGqwBDetg+YQcQUmL6Lm36bJOslrGezw1G8L5Hdd8HPlHC+rk
UiL+cVKIR8SCrmaRNK3fznPJEPMqyxCJTMw+EXzIYHmcYtMym70BTNAYUB7dK36h
ypNwT6tKVDxD29yiRDHzW9WNLAHu9Syhs5D3mIACVR2+fa5yOEcdTpovmmDLzh1r
f026NCZDBy9gM6ikCfmvhbVpTdCrqjPkmROXjuOHlIzCWWxX21/ZONvXDSU+Eiut
5JDBcWNp3YFd6cDmjrudLReN9XDYF1H384Av67be7Tp3JuVCx9R70upxVEgvqOV+
wI/kGWkKfa16wZENEzDqSn8Y9KwkyzPEkj6swzJ5QlwJoEYQBYkvR2xD+MSsGinP
joiTzNwMsS3xLJA3vyBYs2nbsDLDQzmoRics8fCEdNUG6dTP0pvWH+BvCgBI9e3I
j47Jse+Gzemhmg3JnI8RyGu/2LibPpqOyrZApE3KlS7Ka/+6+o3t3yW5cYxOVLeJ
AlHfdhuhWBzsxOn3O9x3yvTzuj7uehGxPW7ncb72CHZB9FN5f6Pg8ZR2SEiFpfsj
c6hrT998KUhEaq+OnyYca42tbJSxYI3ewwNHoQm/qiLn5ow5Yp1tCnBP8dvLPyS3
FgOr8PsD3klQ1kbivfmZ2JZ6SWxqvOCdkymZxylNDYU+IgUwU+dMMVadXaCop5LC
huK4M7FvmP4NOqMqy9e9Qfs+Gxn33jFLQK9j4mRhe4tVe4FFSv6x4nCLsCvHwuyp
12ZTHaKAvHLmFoUIsVuZRaNoWaZ14Q1RQArMuDqMwLWIQc+EvPRtpsCje4hM2Elq
3rxEc4f8+nc3askn2YMNb7LfgDai7bPdfNJwz9xPZyUsanDCPqP3NEW1K1WVc32G
jtecpa0oiM8E3ub2FxJc46rKdZXNy+eoVp75h49kYZQdH5O4BULgFPrWN/WtDIjG
WgLIYby1Zrxop/Sr7ni0/38Xa0iITbMIg6gV/QZGT3tUR23tWMdatORZ3K6q4tz1
JOAzJsDr6xAbYaa/bqiNsgE24lypTBjt2/jlFMWuncRWTSl0WCLaMBxjjHhgz2VQ
2OlRuHxCcIPlaBBVwrOT8TdG9kRcuCe/287/sbxjGsLMLsoBIew+jVa2eu25qQ2/
vTtMFmM2LkhB8USWtVnLwHJVuF4m6D1FheNTmmLIwgHXiE435K6GCQesfKUiQRf7
SCk2jAOCxP6q7WkU+4QpAYNY0jwDri4LJZh5IezOdmJbtR9jklI885uS6OykW9FQ
gmxuX680IiKYmucVMhHJy1dhJS0daY00JBjw5F267qeYkGBDwt02UQ6IabadGI4K
Ojkp/VpwdA+0t4p+oW+VCN5WYS0noDdC6XHu+x1DsUlA6g7tQJ9p1BFTV49EZ1yi
xiBHknGATr9pL8Y2gCw6QB0gwI3y+9omQMIZPdB1C9KUA0DAtgWYaSlaFDaT/oxz
JeN8z1rrUtz0QvDhGjXPHD7OfmXUDW/YNERajkoxD7eEQb79WkyllxIjAjMlhtbT
2LZtX+GPrbfk1r/lJY/AP6WsFQ5lLMbGt0gqpv1cFBZ7aL317uWER9Lb5qSMf/Vq
CqVNNyPeyORoURn5tHyfEXwXH53iwB1mDEBo2RtCso4FEPS8axZbXwF9aNEq4C4J
l5RmCACiRboBLAyb9ko5fSnV/ccd4gNyQZV4nzMtVNDTWsjyv6zMTz4hM6j1yeeT
43LjER7GCIEbzCEBQPdb9/lxZUQEHNmZiOHVlx2hG1WRhjo/zZ1vuuwti/oR57wR
Fb7Y16TA9JGngiDJYepPkc7rmnJlLgtkLfAcLRX5A+YNKZ2KlEpgPD2+I4lmKq9P
WSsPFyAe1wX6990yjxriEBlFFi7RAjuatNXzhtf2beLJXMSBTn2EAbjCsllqWJav
apFcRvKhwsalHZbzaqwXQkZ9418+90ySiK3x0Xm2WZwHDuQoKBcR1DmiYzZEIyD0
t0sGU33WIXx8KtfRIJ5s8PVVVn/1yBEK3D577Sr0xuiHxocsTiWFjOgYxruZKLzD
aEm5cWIKiSbXufhSsANCz4NJWdPorvTLbgDJGX3Or0ChqlSqJATVm4afTs8jaLE8
+h52/BBzqFWjlWx7DF00FIC3z+8xHflJhUoB3AC0hAk9k37cTAkiupQJKdGsSFYQ
HanHMJ2Yr9XzOW1hhEr4LDBIKm7u4WXF0SUBYmP/KScZRA8+UhG7k/tG+dNsMB74
Z26+J3ljnTbIdU9crTJ7tC09biorLPEdXAtnbHaQU4UzWJkEzTaD+npsbptdBKRC
a4e+ICvke8qAygAZNA5F8aAFsgQp2Ch/1Io4AkxzxfeRZbuAvJkQelY1t3K6bpFE
XKgVxCIIuuVy+qPL26AtwsTTdVn/g2aa2umZppjwaxYOujI1vg7P8asPYpFwq6Ff
CXvKi24GiA0BnKbV4D8yi7SPUR7nxvXXROOROzVIM6ZPg4uRfdhuPeIpBZpUT3s6
dwajlCWsa/6mMY1U7S5SR+jf0iagyQcnYPGg6Av1kHt7Z+EJ+4c2u2iqqH41OFmX
3EExb/pcvg7+OpMIA13FlKfCLt9exbJC36w3MTdUg5yF9BZyJM5dFn0BzSXUd/jN
PFfSnLxhFtglIOf/QhYrdbguJJ/9TfA1lWxZhG0/Tf+rLIsSOB88TNL2qV2MXJYz
g6TihIe6be1fUKBqAUlg8r/BjLqQRloXkmk71w4M4rWpTFnpvTof4w4NP60ybU6S
ccQXfqh7o4pnVJFAuSovD88Tx+91T1X+hJ1n909Owt1PG+9N1feYK24SPwZ5rW8m
rtwYPPLfreOPC+w8CwTh6XE0JtvMTipfh68VlxnlP8uiwAKoGNhAde1O0d0dl6LH
TokcyE2PF5dZ2kaYBNThTreoNFY2r1jVN2OVqJr3MAdjQBwOuSQoT214sPLhdGaP
5v6+7Okq49gWh01yQYZY8b3GKKOufIJYJwMPB07npEc/mYMGOITb1Y2StnH5JAq+
WcYPXI29ZD7Vw48EUNgptBabPK6SaCp94lcPKVCP/sZYRAKTPoJcQCS7unyhjYY5
HBJ+DPnyKpgvBaIlz2e3PxHMzjX8mqOFks2AQF/3lfemTG0kBOe3cR1CjHLebf44
HCq6wZMUnhKj3f6XtOooqf6MCxjgPqVSIswpxY2rOcUx6yFpKoYHaOkTV/2KbePN
VOgNm2gwoDwnDzOwAbodhsQ2mRZ1h1d1+SHB9mwbVM7lLDfqgP7sq3ATcPxgiCmD
E1SLz9hdDF4mm92sGoHOqJwyMhczwsKAI2JWGTmYVqvPNYkznLiTH1c8YeV8b4B9
T4pbTb1tF/7XJVKF8ygGyxBOolLC8oriIFt6IbrnqmgeD1bdM8440ipr/v4tuEyd
Qy2QrynD/TKA5l8AwlTKqB0vRErecwOS7VjjY7Wiob1exfbTDLO5f78OxjFkYmpU
GP9EDM3rxLkB6QvGstjuZ6bpxqD4Emk1DmtNUiDFxN2mviJP/3akhU2/84r0r5Qz
JXC5Fa+Rq1iG0pfgbTwCSLpxYj6B1rqA2MNjQhJTRJdp7cPud0UxrBcw8B9Neolh
DC77QeHXSUCqXNj8Xft5QlUny+KrSPj5lWvcT9Dw4oe8IYrhUyVKYsbXT47JFy5c
Oz/jb2i7aArbtOMJ62rgpnAsBnxa570siUybL+EQgWOddUa2uiijBtHncI/cAw+S
llZIzXG17aCaRTb1dOASiJXOnpjI3VsUA8HCGK788o/ZkDbnaHzo5rzjeCnU7fMr
4FLtQ2aMnM0Uy9JeYklAj4OipjCrxxcP8ipwJubZ5p9dQuyU8c2KQC7fFs6k1Vhu
TabgqsI2rlHHPDYc3oFW9gIQkUjTxGRO2IoPVIRfGfQtW1yh4XFD9eZ6m4ZAxye+
dmXV5XCKn//2V1waCnNrZ9V4Ge/u5Nd22I7if5U6kEb8ZChkd4gas35ijsY30mO7
EdRqriVaVwVI4+U7TGqyUjpVo7i58m1+HoBuFX46m6eFE6q33cUQ7ggbVSJ/MQMP
P8ZrlTpoiYjBvBON/x2CHFf8l2FZXrTwV7FWItXQCf0XldwNz7xu6o0lMWFMAh6X
LRqIUEl3d6zEmmT6vntogGVLMQUzDyakUxHdaKkDb6aLpGItynxHezNMXYR/XqDk
swndEm8xWyMyvYewUwIjDAZf1spoQZZ7wWWfnPlVUynSKkT6yeDTW8s6uSaeNoEs
UCClBHXQoMVF2EajqlZrYYFkgEcN7V/46Ohs3//xgLDx35H+HEj52EiK0nGiu4hL
gY907XV6jW8PF412kP1VSvV5M0MhXgszoPPgzRqIzP2XLXYRznhaJ31ty8aG7e2u
jUg8+JTNBQ6PTSyZYIEdnthcZL1Pqc0cWQiowZ5NqomstymAVM6di14AAwauORtW
+6VCXoNDQmTkpjfHMHfBzeN2h+J5D6UqrZP9KtJyOhY8gbNpiUJRH2mCpkfexP1A
kIzKyFN/jWMrX8mJUuUThmJSsZN4/zZp5EtaqhAz+l19NohYTcSQoUxoQMg5xfk3
o16rtIOxrGDz3A9u0IWy7NCs9csl//fcarGmxk0cJgpiDcOnqittPcMGHGfkYUh+
+a0gx0a8mCO2rD4KVlOiKOsSeZ9GCOci5ie/bC863YxiCdNVeZx5TzeKdgBz33TA
oXhaqlOxxmFTZMsUgTSh6D3XuNKHRe3eRAg0F0+1HnJdD+sXBz08/7ELHnL6+9j+
rSgPgI8pQGJEvPLopsy93JhmQv84zrwquUdlruM9i3SfhbFGTBgCfi6Nqqgl/wxC
TOnOCO5PDCeE/mDWRDaiYq97S3bIleTyc/aMi5smQkfvdPFtsqXVG5oCA5qxKnEA
PFSmbHBne+ezC1rVlEtfPNNNyCnzcvWIC7lcMRi6MVur/yTKrxwtqWDCTx0H9dKB
LbJ9zEvdeBkuUo3hODpH+t71G8eSOblutk3eJ0ISERXTJEf3mdWs1oe890oRN8GE
sLp81bdXHfNcg9I4NcOsg1UyRpxoOhmXXURB7Ko6ynu3rkAdUMVQcpxkem1UUlB7
X9cURP5xdFEOmz8h3U4zreI716yVJUHPJ99hXqpWGZLoEjgoQMe+GocF26J408f0
bIE57FCis1/WpNBHCndzWZ7IOgqiUl7/Sq34303LnCzocssLdymTdzVnooMCssER
YyL6dHo3YWaNyfayHK+8QOhqUXvr6mbdArCs05sf0BjBkco+JIJIBv8uoYAQkIMV
uZq97VrVTI6gTsJB3GvD0cJtPKNOw5JSLVXY0GrdWmpb692fboCc/4abc6gpK0HY
EzoIKJWOaW+FbJ9/XWpvwjJIy4T5bkVdrvDBbynXpyW+O/jN00M9BTPHz1iOQ/ii
uB/zLUkkc4409g5jBrcAjWuN9ANgFS4FxOncMtMjt9zzscXx2joCFlNgzDMf2uq9
qPoxs+lhnT1cA8XX7CZkdpjVIyBKtAu7Ok9WEvAIfThU04np+EWA0v0jUCAxW/zJ
F13eQle7NRd9xWAjKXNB94UdB38n0CroS1sW9QXTM+vVNDb6CUb/SwWSxFGVvf/l
ZZdtNt6oPGUy7+MY3O50+ZIjgEnddwYfWGEAzJiojddKaECyUzKpio0f7XVFA629
fzhzn4Z2EMeDO3AwrFYl46Y8doVu8eIjzQ+3u5ZTajiGrlqeZ/NrOsCa/yyiJe9B
on2W2+LeWwu7DcHn0mC4ZMbkdaAOItLGWiVMwYwR0Zjz63/QVKYBN2eq6JLYDdkL
KgenoJNJXQ2Be6E9yjAFdKm/60I0KW8JwKOPg0XsLDcFUdqtQAGCnU1FkCxnzy3w
/HAJHihGf0CkrOJMnABuStjADVSjadwPoJNgQ3b9cUPy83mDa4TWCcab/Xz1CYXd
45Z9oEpRTM/7voL6KYPYAT+9sW+4jaune4C02tz9NURteurleFalrIIocTn3S/Ag
ikIrYVl10aPTEG5iGU/3gkVejdzj/rGaONRaQ8yQP7HDwQSHR9Z9uoQPc2vVjoY+
jvfsDtjZNVYRBcPIZ2YKgDaI2uiX3cx/dVdNv7n+O3yaCrIzEdj00jQJAf3PMEig
x8e8slasWjuDbFouSWfhDbqIPnqV23YxA0ov5MdkBFiijVvAYBThgX9R3uStyEMK
3/hs5oLwqxFRbRGVTzeQUUnzXoqqD8zIK8H2fa3zOosD/+lpqkVf9e/YnddnAzSQ
sRY+AGHojf9byko1aRMctiakVQDfv0EgJsLGbm/g3cWCZWcZrQcJKzH5685P4OBf
Y8GItNEyAsovEfFST9xwNKK+w7bB0DjDYrjBIePNB9O94tQMyw881KdXn7kpjzK0
F3FEktnvrpLQ33502SR9jOm9KnbGnlJfRZ7kterzFncBqsyAt6zZDKMdYvGDx+YT
nLWELMxxmbwxGddmgHyCKuUtyIPDGhPrkAe7h7U3YTu1EClzSH7gN368Y3tbvfV0
irE4mXENFpWew6lfl6Vkz8zNdvXmEs36+aMfmoAGYr9SFCM7t5ovWOzOev5Hnu75
MncEHi9hf0kn84S+48WfZ8chMBKMOo34Im/RVfhbnPv/W6cJ8TB9SLFssW6Fybxl
aGw7ADGhGpl8Sd6DmE3BIXS0ZPE6yxVKj0tuOY2wVaFoZI84jpPnMpnGe7yPhIfN
uw8XZSGERq/wW+jhCUJXUQGIm9WfcoPOCaZ4XecVajmRk0UV6JYE7Z2KLdNybgb/
AEC5GwRcaW7I2rfEWqSJFc8qhF+Kqr3ot2lwDBa4TYauavYW1FiM5ghmvA086Nil
JxXySN+0TvIte5rU1q66BIKJ2gdMSRH/MPULl/s4Usn7NDIt0WqiaceWiO++3yvx
4ZJWruZAQrEVDSy0/X72n1EMxNDSHQa+MSQrF0gApdwg5Nw+xtWQ4Z6FVTVjXgTp
tIzHgH84dM2lxC7jiLjg4mtZulGKQgxy0/p2o1/nIn3FkQs6MDCHwuHrtSs9v5rR
JMPDp6oAInNie6rF2hQKTt36T6rWZR9rj0P200H3B18DIj9hXYvSFSkwvv8XmYGr
zQIj6MBD7RNyePArxmW8lHI/Z5RaKUmbKjRZnLLE9hxX5aaZ6K7kKFKUaP3zJ0BO
lExJKSP5JZXpvDLUq2G6uBruXYyL3KnHV/RxGy8fsBhNtMQgBEZ6m3oRR5JP+gmh
mr4ns7Ah+29XGjv9/DrGzOj+CQsD120ikLCdZRDfbuaRU/eib0NT3y1Ml4C1Bm2t
jpdjKXOiDIPKimsONfblA1UAIuhJWJSB8nIC3pDigA/rqtdTBJzQeev2o60KKWEQ
nZ3nzDTgEcuu46oSnR043ZW+SQWhhXGwdEPv+Drp6jfz3QLE6VNUS2M2cjXxoRdo
Tf2AyHZkAoliVKDlaiLsdl0MNwKiKBelf3YTc26P2zqCbE1934TPQyRS1430xy58
3Y1+XN4Y8kGz+TEpc9ZWjUT4JQj5JRNg9ABn/Lqfs+PMGEDnPkH0fUz9xHfC2NP7
4Llx3t3MkvFbmxbpCD9ckMxGbHXg3OGTOogJawAdRHCuQH2BtT+6n33Lu+EgQyTl
YDZiFtRDegZUn4OAYlnEX0BFWlfQ36PXwV13ShbpGmgIUPhOMzb7+2Lvku6okv3y
z+MUrFtkAG9qiEIeDvUa7rz6T9V/In58BzPjMTyup4RtEJd6vhCs+uzFaEjZEUGu
VSrCvSrU8rIQzFKiTQFjgx/0k6sJfdYkTsA060FHv3RocYzhE6crDGjUuqp6Povo
vKHw3KU2+/AvCJnIGrTFjiYTFe9CE6rdSBkKlMYkSSDh1P8poUHVjG5s9C3x3K6l
5ZHzdeK7hka6uZgYa38jJsroQVLrR0umaIVanqYTCqFbl9mJIEAcaZF35qZ2mAWr
HDL/THFSoHGgVnl50t19SUjBG0SUT+VgIlWNn2CjX4IqtVY0D9jO48Fmv6x7Imc/
fVoisgzyK1Hkb+tKFrn3rF8eSJt6L8YWiz8NOvyP6RP1cPqc1NlCM0PlA3RsTN4f
S8i6HFWwSwmtwNENU/TfpotWf2okjJBMjU/j+LUvndKjn1lA6I+++7Sf3bCA7rv1
5RxdmSnyQSDYRDHoZrgp1QnegOSCzPtxrTMwwXgFIUXcT+ukCn+7OahEcPws+WiC
mkrQXbaxkuQywABwVJlWEpWxr+ZcmDbxk/ezeEEFhnAM3HQnBytgNW2OaknHtFTZ
3eTwS7jRx0WHw26xRnWAYeeXsIY8+9MwY6WggJlcQ95eOXFe0oUpFmvVeHdb2Y85
DawXEOxMd7Sk7hkrWFVdGaE+AfDXfhPkBD64IDshP+SCxr07Rag8667QQpenDja+
Zyz5g1qjpCkcPcW7J3e9EIud/+k6B9LM+Bg4RF/TgzsVKQj70iFz3gLco4t8qqj5
0ndv+NceNZ5KFed+X6xtP36721PMVUPbFZn9DmQCCvVi1pUZWauyIsd2nPhO+Wwy
zVXOibj6nMiAKbqt+cg77R7UGcpmu96KSqQE3lj0ogF5vfe5ODlq3qZqS+1FKiWV
R1pq0ZFTTAUzYx8u7x7WydsoTETqG/I4Fx5yooIp5yAEHqudAB5BfTbiJgC6r7BI
4WP/N0quiUj+ahWxadblbaS1AAwgDQB2lozaClIy9mgICd+Yq91HhR8/cT+fVVeI
0lE83j2GZfF98o9JnQorwJ5iiBJJ7RSxp6mUBoT0r5hXhR5BrTP1JGU+cDrKSIoj
IUyExKr8DR94W9RaavROkKBJzL9JwndoU9gJqGBgkVd2HaUoK5PmxyzUi98TXikx
kPb5zGQgdKt2Rv39jEfmBn5EV6gell/gLjuhR/LRTTfOpu9Ipc2IAkYx1XlLfEyh
WCSNFd+Q/pnBQnH2+kV25wQDi1w5R5XLNEBVYn/yvufvXaZ1U0Vst3LQ9592vQfs
k+/rryHdoczrN/RWfFUvKj6RL1iza1SVcarvE5QyeojCdgFnbbgbMjftE+EfVNwL
RtT/BiCBVE2GisDaoS0xERDD4buw8qgbJa9wyeKGsTLYk6bry5zFbwNBjKvjlKIM
ZvedubRLhqIMbodONlBKjp5cJeiZ4RBWUx3oqcI5C4RAvkLUzrbloU95ZFEY5CAf
gNn9zScbNemOEFJoLX68uw4fQ0xJgtUSJpR82yhmRO4rvWqONz7sT6o2rITneJpD
897YAVJZ0laUru17sFGHOGpHjJvxTbyTThMmcTjS8kRR3spBH5i+rILD0TSFebFZ
bvBI6uUUx/hcTPzuveV9FS3artAbOu4HlXY8fyvDGIyEoRa/0E/2lPXz3UDrDuqn
bA/OQxWTnpjepazuvOf1Apo9Zx+C0PM0aYnU6WU1sXKf58sKyEMV4tLddM7dYzXq
o0C/qrYMdriiLdGCXE1dnPP+K9P5Rov/+S8ThtQHT9algGs3hsfcz8DZehRwttMY
Iog7XrYG5owF4Aoexl/s1h6RZqIU0/2RKSJaWxczMkbbTvc8PEcuzXvtHjg/YQQt
XOp6Ht7gd22uLUN3CgowgOl8S0xtB2xiB+IN+EPGaGNbmrSWA8RThn88TWFyXagW
bWBytfqCmQ66ZyjEEW/EL5AXCl6k4mxZEwG/JXu4ajJDPT4YnGpNnoNMgp/zT/Bo
VouWNQ8ySitEiH9ZliksoUAmwIvgYcFRQ1rFdp05iijxfQV3kXKZRD5ZwNznP5Qp
rNedPSP02njgHserRj/klgZy01+EgfEhx1a0Sl197JTle7UjsfIhLecERRcMx6tI
k3kr3DSouWDPF28hRdjDFOPTWhwEBfgXAc6THjuqalWEuk1ag9AWXJDAsVkzenay
4x6u1nplkuMlELdwnd7DS4KR8D96n285Cx1gMG9W9PrvyWP2zMQd5BHILhEX+W3I
WMfPz/nDfBm9tbBdkUIqwGO+z5V0Js9EzvsSKIsPjhrIzWpvxqsIrwyMASMNQF1L
FHRJJbW8mTntZzAi7+xCdhEIOCMNOUhDQnILc3wYnk76sHhHee4vTwH3WcCAyGzj
DFH8f54Ky13cLrcK+B+le1O73s4ZoiPrkWS/xNbJTwP61AnpO6bhUGvM1JL3PF9V
a23QMPcesVl45rLwJNC/n/efghLFiGToIMnhowqcgtGSdw7VFcSMZPrZCYR/AIrk
tYmn8Zue+jKMc7PrvqxK68BYwvRpd6S2skasIQmk9UTtHg6zO95ZhVlHnkAggF+8
MiU/aDvzE/s8dM09Hrx5zjtcx3Xu+Ecn62lewStAbh1a05uZr8o4lxzvRYqts1wa
GQ3oflLdaeOLm93CpUtKNKp5nPBqWTI0Aaj33uYmBJsIs6UD3I4ru96iXo9uakgm
JkvdrVga9TYhEEt3vILxIgIN193Y8JhbGtESkJUWQe7owXH7x01nMKkFxJw1Dm4R
HFBmzMk8tv7DmtIKN0DPVfzU0KcEZKYn4RfgwCiThYlVLlYqNnbTPwtNtiwr+avf
ZhQ3UV7dy8CJt2FYRHeFi5LQBoPKveaaXigoUPoM2oVTu2bjzRNjGJtfjTyFl2hc
/vFnbKRQoDv5qeYLleLkqhTyqkV8NQ1pBymIZZR7Fz16PygYk3sFZRDyLSFOaU6P
MB2V7K2pUyfxI3cko6wqMpIbWZxQ62qrgLL+dOyvm/4n5OJQIT47EQZU2aA98/Jj
02JUNVOHNPsnYEn0q554TSqH6dUAn1c5SlBel+aMYuftviw0xg+pKSsE8tOdEZxb
5qAdnwN78GqYxShsB3EVepT2jPC7yAMQ8uWJCYKnTePsxnGMS56FF/MgHd6vH54n
NrRb7PtILWDiDnHlwXwODX3NCxkOqvChQ1tb9MzxoeBZZMY7PkYc+XwYxwQEJogP
ToFXE88ujTEUBgwLwQI7tvJI7lxL7h6Fs6eSSu6237w2E0ZDvzMbPo0K42rR/fua
zub3xwKISBtf/8Gq9aOOU+hwsCRqz9w7j9PXBk1fKcx/SeWfhiufEQXBiZ8X0fPq
8T6Ulw1aDKxDGpbZ6lwHEJdYs0G/BfNPePw3Mc9A8OFZdql8yiRx+e8irCnFvkDP
h+ewwePnkJ86uTfj+pka8dh3MoaNiJbYkPfzI8Hz42XxnPjywqp/ixsDsl26BfGt
n0Ut2WCXe2+ssc9ae/vHb7Z+UV8W7AoffINuMwBUqYjNQl+6bEfb83x+EaTiW12J
z47sHxecMkKh4facnJtZyB5SDdk4YegX2I4Zjj/gQ7ah+Okg1yh5MeR3jXDwKww3
3o6b0WKFnvcKCMJuJlq5BI61Os2SNrR1+Z9CEAGsh6bVHEzM21Q5ucunnp/xGrc9
ZnKlUB8AWGcvNcy+dbzZ72Dr30WFHzKhU3haBC1OLwN7gBl20Hsg3A5Lko1qwsB8
XmT9g3zBo2uJtbmhDVSszap1QxAlaJzEImB0ij8lwXmosFQrvyAVc9aEq3H2CmAm
bHF7uI56aks5M50U97j0F8MbvkhnY2EcFbCdE/7mKLZ9c/xYHlKBv0fSyeuiyXOQ
L6i43+YKXeVislBOInALW8Hvop4jydlbobvK4OMES1zuRUaN1StPCt9wsqMQVziy
hID5saX3iY0Gf7Qn0dv5EFfYbYhCmgU05XdCbAQhF1DdFqGKhAFqun0qYer0ymSC
jjuPmcVFFcUs7Xse04gBUF/PniAToERoB6dfdM4vd52msSJukW8ZFCm5GhSMJqLV
s8FM7VuxkoGI4kYJ/qB++vvsbQsizG5OWTW+hVFUd0oxFLjLktyAg8FH7S8eKXjo
/8FvFcuBlOCgX2TV3BpU4FzvzVdT9Ndk7xr1jqT4xO6ITgAextjkBw/0mHxepil/
p73bOet0//O75pnh1lfwEwSgEZAIYZ0Lg1mJHu6SNgM7IJtP1MdQxQ2Hp1VV3oQJ
+oeBuwIf+szwCk6lCmoatz2H8zvqY2rK+NbSe2rqiICRWdtycxrK8XyH4UlkFQnN
WjEgBin28CIi72FnA6R22GOWoDqT3mkt6eQxJvp1WG19UrhdP6srhqxePuiazWSw
t7oWPBrMmW4loChtn2T3hHPFemPkvFRjoQiEWnSEkKB+T8vUHOzSoLTjpPWTrvHP
RG+vuqWsGePrF2c5kI2/WnYbffJedbxomSlY40d6yNF6x1HHQhWWuxGsdSy3heeN
E3sB8RkW67Fk3id2MWg/CR8tH0mXTUsZIyILlZRnsV3hDudcrvH6YAAutRt8ccLZ
ca0IkeuKO3t7krIHznBfytkMf0Ygec/uZ4jGOei1aQlHmZ7C7Esiz46i9IDkfu4i
m+6MdSrNxbIdr1w5mKcjgOD7zQFJXwTQXMtRTppMLV21QP+FAbS6OUrq1paiEhp8
p/2jJ5SOMprmBL+9njmi+wr3etSWXzgAYvtOaXgLvREUF6g1MH2woiTdY7OCssxG
Uogly3hKhQi6j1j/iE7fOOkqGJJpb9587WLxDA02j69qg083PxkqNkMIsH2tUEOl
FRhpMgq0BhDBJvue1GzP8tif9m8M/KphosRZj9BbiDzkshZOu8rrMHJ3jQ+hVRvS
1T6nqXO4ong88IrlFFuohdFKoDzqTfCMM+594LMHd32By6ygKxje7A1DCC1ZcLTw
LZbqVyvS+bpRSLurW8XFYhEtyAvzIsB2vuPLMMjZJvgbSxmJgyEzwwBuIcriBzch
C6fHGJKgDSjyhoIYap9bdZHU0s0WQtlHemZyc96aCbsGpVBb0/DOQ2Q69Sk1BKm7
AT0x3AMNdsx/jiRvEIzZhG/CijrgS6P35LiBWErQtat0lxuNbtIXDJcP/HwZTRuv
FAK0b7yL707demIEtnD6NggUzI3ktGKqHgqp2MzGC148kl47Riu7xSHMf5jSMfvP
uhHm5FL+Rb0mFhDjq43QeaauFT4QRJsKIrxb/Gi5p9XzifY5m5eul7kJyvgAL85I
CgvMI355MPh7C4Pv1ZWn+YHLjsYx1kv090m2IW+wo2hIK3i9V+iJI6V6dQbUY5TS
IKhyRERp3FpmDSGoaiP0bNej48z0NEToLH/eWSVHFzbJ37/vkfXBywcEjVIoTjYW
x0ptJGrHNVAAenQXTIQNTbcjcaFeXGIwYzEa/gACFIQ1YLATyH8nquCKzKMbMETq
EHCGyuynhG6WSMOcvcoW09t9kCSVHGrZEyIW+SFePL2nFC2rv9o3XbG69DSbnSKB
16GbdxjOy0mzcQVacx8i4pTNM4ZfYavFlSDfqczw2vNw2cQIUd5/cL3+7hDyPt3P
CqGtir/NBTjvX2YioZ1doOjMfsxu9cWl1p+xCzNq3X/2z4dTWEeea2smU1qoar3z
YOWLNRh6AHBDT+L4x87nMVkH67670Tx7I1w1UModUZXGFhrWYDeUqUSFZKjY62C2
+ms77FlAMGItiMAzV6moqbdBgnuTAjJxa06HYSIZJSM548Gl+iix/ydn1yD0iK8I
vl9RHqvdXm4AB9WgkgQgR3LNm66jC3xIf1hCUMfjrQM85MfQKOveCGamiGG3ggeE
yQb3SaDqmWmIdMije8Fzy2mfNAF+nbWi4jbeeY1ANbLBAtsoDK0PC/VBdwLgWK+m
GQrVqoOUwXhaq04+xdVW02OsFp5ccCj0u+RNJkIv6+/YgAgAuhpwM7IuGMwUbrId
Jh32fF1neJ2+n8JqL09kdDA3lQZDe/XQFi+ztdXCsR/FIwtaYHPZavjVwlI7itYL
N1XOvJPoGN305kundRKVqdQVVnzyX25ku8PV1vfgETYW5I7COYLDOaxLZHUL5uAw
23bgzE4tFcl1hQLp8NTwT5tLuGaOu2vgFZ6mIWZP58K8JZCkJmew/PQjP3181a3Z
mvyZsboXCEVIQvb6bEOXVVsedhemVOQN+Y6f0fYSTSKOV2ystP6LzuvPeY+nu/+g
jaXSxwWZB3w+6Y1nVp+fNQcaXsJbyw1WN2xU/uyXkIUqukAFgdyHzMd8zcnsTXEX
rjQJvYZxQiiYztf+V9VXVECBxORankb9VLBDDDFwwYPbedJbBEfMtDmIwh8DAZBu
znwk4W3Dc8heqOMy0DBZQM08b2y8AsgbT5AhAf2J9AYsjxQUYnZnUg7QM0TM6MRn
d5J0L2VB4rkDx/dG6NystcQGyvP8aUOcckLHS7K1e+TnJfSYreLrUcGePZx5csCN
JXZBPY4qFWwhp8+iTXBMeRqluSGVcpygUzr525mi9zrgU4VrDGfkKRdUigJP01rB
0uSvF34JaWF5hHE95t6QE19XaDQBqrwoS971ia2rTNwNO2FLQ5Of8OyfFjwcYPYC
7sb01sQfEMWrW0eXck3geUiYnR86qeTu8XjrVRzpbKXLBX07Ayh493Tu/lmWGQhS
I+aRLV6JB/FtEOkNemYvj8Kks1qjiA2XY/Y79JAh1oaMIqebRI68fmejz5kDgjjH
PofmMXjBZLkuaPGhvKarBJq9m93FDuvgrt+WoAjloBFOLWL4hof4QCovH7U9Jp2B
Y/xUG3jrBqv4vRG2RIuXGJdNuX7RHzgNVxalPFKCNFfjDR8hI9Bb3vVAv8u5WN9p
VVd0dfiTKHPhvSrWjdGbsjykURRiV/dkRQmod60Mhuc9e5T1IISHYLODoC+JkGsa
rE+ICsP7enKrEGaclgkCax+UndbtcCUVjhtZhvrPrALVOj4IcMlOP+4ZjdKOAZ5u
N9xFdEbvaQYLgu2iMXoDMUZTy9yuyuM8BKBXG0eEGpqEl/ju48slbmKxh9onX4kY
KaIoqzrXYIJFzKOPDa2eiD5Vgul+nF08UI0jVuBzEZnB+0FuN9L06MdqxkbzA4nc
BAKZlC3042hrn2OCoT6wDd7dIZkT1WBzWrqmDcZa51BrWHO5ysnnC543sUMDC+y8
wJVNRRiZDCdfXFZ9shk34n5ivadeB7xURVqyEPUoYiG3WYPISFgYCofQchjMcMqX
x7Anx6JVQ3w3mmoL4KiHZkPYCWqZ9TOmPiOnZUd0GjPVSCJOnfHo8JmmkJXt66wT
dZJ4g3OOIhIUuDCitaVmQk2+IjOMgdqiO+zGyV+kehK4K1XSTpvluXY0oL1sWRs+
tOALbZrmn+k2gDBme815+LnTh1ryBrGj8xN9SN8AfZlp28Xi2JFukiX0DQN1fZMs
USi4G+gKCDxCSmRgKIX1fGPXnqPZ5XU10q25ScHH6kufnKiRhPDYbgD92aeUOXJ0
q97CBne4dFA1Wn3KBb58krT7wspdbUkk0Qe6IR0v9Bo10LI1xfb3IC2P9ggoazAU
eVg/382NltkEu8puQC7b+8d6JGWgZE5TVd+72zwKm3GureN0orD5BOkLdxggda6G
hEPf/s/kudZvOGhN2Hvf/Io0JeMdb9EHzyzhlLilWSvXa/Cgb2QvCbmMhWTBZEOs
TZw0RbJPgVBTAFYAo9MxRP4LAR6kCxjDM2qxq911t7QxR4ly+Y6jx9Gtr/T02baX
/rCSJdfoYh+tUaCSy9zZiZM2Mu1KhpNmrqldO2iOAp3nCw44CliEpYBqTdp5H5dg
pIk8+qOV3RJXj5Rts54gMa7BoeVDo1K0X8y/pYsdmNJr9LsotJud8YF/Y/11wwtv
vfy+MtIK0ROi3YI1r4OfpTYSGx1F9VIQSwNxTEfJNi/viL+87kmp2M5qn+v+qHEE
MGUQRRnGTWNpSIk01g9vBBK+e74mK+4wwF7cjmVbrRXmEZio4/mUlBTAKdC1gqkr
y/KFTfZD8MpR8apg6iqWYdBxpQzXRbYu8SvqSwC7CuqjlAIfIllbZnVmuusgIwE2
nfx1HH1HCva+d7zm+9mMyOwu6DYQdWRYr/NBIW2TrMLD4uEOLVqxcnaDhUPbDN5+
s47+AP3O5mBS0QYc0AnHuM6KUt3ya8N76sBfciAcnY3qc7hTIbeuTBMUonVH+Dlh
RbfTZSaYTh6mZACjPXvvRZH89djqRzwBjA2HfbDDVZIbNn0RikbLZtpV38nKULai
px7gAusvPckyy+PhnDRXzrC42iHv9D/8YAiUPjVNdoyugsFvOAHo0qdkyOCjHYwO
7n/JmWrdXtk+zwYrYZ7qL2gheCg/Yb4WxNdGD+cTOLoQqKAbz+MDq6VAfBHveU0X
uJld6AAy3OfDLIx9oV8lesJcSl7i7w7szt3nYMWdOrN4z6fHxIdYGsuyt0tqZg0Y
ZTkgwVNyaKnwIxzwLYVINTsLiQPvCjdJuBPuRw/sRrGbNPsJyMFwLE+xHqead5N5
tMLciGt++MPt0TojKDykBrvguo9L74EQLxX8dmM39xyY/p8aWAfkHe8TWAahzudc
pt1ctcOv2AIj3ZTTmmyJLniRVoUxLxpRurW7ZD4H8xNS3puZB1GMqwjEXl3jIb+B
mxHu7Wm/WDIq1vzmSDRTxF5Pdt4v7xwgCggS7VmTr+TpVDY8rgbZ8ehJWxkdIYsv
F7gea01RmyqfdDFESpfcf5htIeBP1VSHLd487g+3yGqy9VGHBRRxA8Z18dQlOndX
TVIdTh+fNOzF//DSODoFnc60j0e5UnErR0oMvERbLThb1S7uVLksaL6XBg3SRos9
Ld8MKoFX124IRNQBwv3eDPFnaslmSk9pJScLqzgqOj7zTIZ4+fEPNWObCoXCt9dp
phRRYpswE93KerRGjpZFtbk6MQW3XPvyQjhnyFxJkrKY+olw14VU8fEApxMx7hQe
qEMpNyUdisdx+gnKN+/ziC0FWUGWuANZl9pI5iMFZQSSDcMSf2N6Jh6GyNDKZXPD
5nJmjJu9ufyo407FpMhQRzTVbSGqsOd1SUwj9C3eUCyUCTnnwixTUx3D7QGtvtgX
RurvphWokreZwEDHwwRDZo5zksxtO6ih/LcW7zHUBvNSCfM7s89tkX9T6cDTjYzo
yKTT+XDY85I5lnsupkuADuNxO5t8vJGUeHbo3HF58GkWmPZzsA8Gh4fh9jsKJv4n
N6+dP42nFPBBJ4Zz0XcRzRDhPzLtYm88Uwtp7iBa7trE6I0+l8ggVz87ukhTlZD3
fgsNjxLOodNY/oo13ByPjQ25FtCoSy/3gxFCDPAn5p6egpd0YLRnFi9Xpc3Y9pLx
dmbzP1+Wy7basREikkUkMsWH3pLDgEptiiyvWh74XOHzyhOdJ2mMg7nWtCSj+Nj7
Rv9Yd9EyYzNltits8tw74OVYX68Aw6SAmSkWqp04tC+2fnaDp5JpY5bzfcNws3kU
aSsbqQb9w2pvdzHWxtGgXnRlJThit+imFdzZ5iHtZE2VrYHFBd+kJCe1KYiT0itP
2L4qhApSQVeo/3Hqtp8Sr0003FfAKDht9V/1EttTeAR1NLcynRMKwl5GPFqg3cuS
d/oVzzqlC9DhIrr/LN3IXLbVw7ptXItiXd4YHwGa8iyR5taorgAiG+U3Q+yyO3WJ
Dh2nhNk3LXRSYnASiULRsY9DVx372czouo3GFX/5jr099pshYUZ96UkgTMVhLWIr
+pzJakaaervH748UBJjHSwmyij+9swIb7eYh/NUxDtB6HGgYfwP/sUIokR5oW2UV
pV+b6Zee1Lf7MU0I7rXO3pTlqPS6BgHRMZn5peXBOfsh/bJq3j3KW725kGTVkTJJ
cZXHlNBpf1AhYhibzqFcR4uHvcCVS1rOo+jJBJLbn07bmA/rAxOLWFEI9ZN/GdLq
bdi6NJ7eFN7psBr2cMGkR2Ux7t+qbDycFNExmqJV5JCQSZusydhuzpUELMZFTUM1
XFCcDmlJYCqbjgm+ZGsyH8q22+ZfN6v5cnvDF4Enu6a5EeVQYY7+Fs2sQO4531rj
KWx2K+JfWDGBI9DplJiiHgNXY2Rsco2aSbOh5ynwRBkiHLqTyvfFsSLf4dF+teGo
1afcCb7rORywSGq8+6caG6V58M48SfdQdPqkiBoecg90Ljowt9S6V2xVGO8BNRRE
CkCDJF403mLQEFhwnCCwM6Y8/0ohEj4QCyTubouG5D1UJ4Uy3V0Ay7klWnD/NHB/
A08TMnrO1sAcRNh7lGZHuMaUXAmMp6H73ArtAPSfHB9Mrhg8+u19Ahsa2g9eVthu
NO7Eksv/svF31Eqi0x41ouTh0e7gPEowMdeWKeQeeUBViMrGjxxlLmySzHsG2nQR
KuJ6t77yIfxOzr9sgo619AShNgT2L91rqGPi4dHg4Tsbi6tYxnlWOH3INIZ/RhOD
WyoPMzoacqdBG1+GgsXoZNOGotrPdVT6AQHg71O2zxkJxSxaGw4QfQTOBo5fwiu2
6e4L2FqY+AXN1g52FY2AGg8JGAEhcVXCWX4w076ksSJuX+1+QCECL45wiEzGcdeN
Q1U/JlrjTQa6/tpRFaHShrFO4LmoLx0/cNHCgIpa0LVj09oxv3vODJpDRu3EBohL
bQVu5D1Cel9u7x1jn0TNG6OEOhPT0BkwWCRCzRLLUTvTQ7H/ETewRletS36e795U
k0iQXpk18Tm4NVtUtOtH8ZdBSEA/3K0XHptHkyb5CcXxxb2VfxAVoPO+FhVYoHa7
LzVe2eloEEcFt5pRQE5WX1Bz6JO2q6p8RyCvkFZZvQIBAcP1+atfzAU+/Ge+0EvH
aRlkBaSQiWcLt4iC0z9iwMOdiTQAQNVieXzfZqKyvh+4f4cfePNVsQyFR838SsCr
vGeyeqLI2o/hxDmTB1AP4n9YbhuOb/OEDcm0Z1oQC8obzTYzHNdIPjOsYzh+vIC5
t/M/39ZxZrXyTlEFNtzgCa5Ccs/RpPJUtY+QwHNdva6FruLQXkP3mSTXKPiz4sao
q309GhdgW/lLu4QYcIFIgBrLbyNktcTRG6WBGez5rjxE36/IwN6IHAbuCtPAwQb9
DjFY4DuTouMl1jza2WrWnmNK9DK4HY6EfrUToRbVN6IcMIjP1fNabwm+9ozuUBPq
1ga5LR1r/NUkPyr3l6vuHMMZy8xFhptNEBrqst6nwagx31StTgipzXk2vOlTRe+T
1lg6fSAlWn1ZohF/Hn0T0a2VBt5tVMyEQIvjCLTzADMeCjpLR7TDaIxaovBSij6z
fbqRmJNd7flHf9dkuC8A56/8G1KK8hF197aemZAjV5BoG3O2HFztlLgI+t8/1noA
vs8383yAQ879DKSgn8cANcbB0bMjZcOVk9imLgRTDuQJ9Fd+6chrHhwtlQkPMbX/
R1+E3WVqP6pOa8cJzgLjSNrLCYDpsQLGF+G0OrmfaQVhk1NihiDXHrvEhcseVf4d
LhOXSuBv+lPsuQZb0Ne3ZxR7OJaerr7EheuxIGrPVxUTqCECkeqrsvkEAMOdcQQH
tO9lUQzcugj2k/4NqGgxpkDXnx08Wx3rwPFU/AWInSdnFWWYd1t19IT/9qq7U1w0
0ltQiKrztp86mNEMtQ4D/nnwlQ77MyKyX/lMH8VQ7NKAtHNBgXy7niWb9x2K4++H
PNl49xRlvvY2PzPBSA75yPUnIpHEjeYn+4tqTWYo8/noW8seL/EvBgmAVlqwn8tu
TTihnTLT8BABRxhzHCIfSLwwU6RiMQtEI2kmKVouYdFg95NGexLHJ8IBQMyxQOwr
uGWyTy9i/d0GYBTmrWcL5Nl4a1Y+arURsaW7rwtPmnHTUyVX50t1SYww3/OHQHit
Ksq4jsL6CS9DGHRfN0804ns4XVca0Kd4z8tOVrBAQa/64SG1/tr7BBHjMjK/KL6J
Isr1O1fGOfJcaan9rYPrblh1+oIBern2oUbkj4oWhXHRg6W9jNxjpa6zWVhSFvWO
oCFddh1g+tJrPtQeooXtR/QTOa5+q2Vgh3NW/VAHR1xKFwsj3VpGnHGGuomewae7
MwCsrU1BEpUy2w8CgRVdNDfkUWB0EMBIwcTdBMxvobCIMLwLTaiqoiEFIeviW3qE
GsTgeEIWUtIIC+28TAHlX2CNxc6ausuxqvpB0t2It97w2O45XrT6OCSTJqOT/vBa
8fZLosvDeIduSrfkJFEyZ2bhYfWNzFILmZbE7Kd0OWJ+mn3n8CdZoALu5hj9cVpx
sbQZBlDi5dBH6lJulO54mabqZzqHMyAFSuRmmuicjUueN+maq8e9It+fAnFyuymf
1Kc0Oxx4JdT5EplhBEo/qdM7CZAyyvit7whwynk2aNVbwRvDSCMnNUeUQ6KeZoA5
EX+okaCFChw0rRPmhq2Rp7Etjw20YgjLdeEVEGsO1dY47gWm6phGVHmOToKnhoNl
10HpW5oKvh4QPIY3eX7axlz+9cVQ2v7/V3W0LnwDtz+2nXsoRegxFBbDqiCYyLD1
273g7q0MVPjckQcApOLKljykncbyeszGd6tAZc6POaKX4adKfmIbS/WYD/ccmxnC
Rhuo27HeYRTPEa1QdsZjgZWFiev2zuDI4XVEiY06Ch6XepNgVX0JL6gazEHSH6Nm
VKulQpBUXH9XVZaOdg7RpYxAY2MCXby7FKwHnA23OkFvaKWdBM4ZwNdnplfQPi6v
hVNHWxxRwiAfl1fFMQFmDhVhxzjMe+hRQ8raWK7Iji9KcNUTtHcziWCa+sqn09f4
TKdJoWL5BNabwnMn0sXD+MY5bf5iHzCOaeQ/bHx7eT2Jrx9vxMLTmZrzFu04moPk
jW9FX2ol2saGCiXWP5HyDG89525Kt8NeyEDp2XND7nxyBBKGLVcgKMHjkKRtpbRQ
GrAkN97X5AKO7fmyqjgqL2OZnT39WlVg+vQY6ptm0tIqoEAef5oj+9R9g4G1TkIV
AdsxVxcrnE1jlYd3ROYXrVp2F/BJUUi6QgoViSlNPwtB+6um7jGlZ87UA708dyGg
n1Wwx7VrJ7GO3aDmDmIwkuFcxX6DB1asAlNF0ejggOuLpawY13lp3SC1CNy/TR26
DbE/JZYRAVfkChYIbuvnsipjF7iSdeRKxE0Zyu81UuB93AyYmw/ek99sIQQkuUzz
d/W9uHDPgrhEBjT587MqoHaBLumrcVSYmxHoIQklZ46JvUz0TETA8iET+2INKut9
BuSql2Y/jTfFqY8r78mI8Gd6gDwwnsadEwyC2bkcaOVbVh6fStC5GH+AoRJCczVW
H07SkmJf3q1Wdxv4ZpJI5uAyGHQ+TO5Uth6lpHOWgRrfAqf5Pz41Ut/o18DuZOER
z5C+XuxRRs2bMK3b6Vqh1maNkMUvwolUWOfcsXw5pXCWGUvrSmV2whb7eKs7BLKH
nY5VJ7L7MFXJeDJuD855D2nldcaGCYAazsojF12R9DHnBWAS4v/whJnjXxqB9mxh
GT8BY5WAaPLYfcw1eJ3k/eeaiY30GNrjKPNTo3sE+GURIowHuiBZ0jZ0ELSu7W1J
IkEf7K8hzdOB0BSI1O3Z3gyiz8SI45cUDZTXVKGE70bIWiNKwEvaFKz7dZz0Fa6c
JhwOC7kruTbeJp+pjeIHhBQsb84RNWwuffZWQrex7PLuTyyNy5z9n9R6aQ5pEqMG
GKhfMfbRrQVHYS9QYfa5PUA5lZNUldTETHhgXIqFnL5x5ytr/6N63T3+UpqasxSj
B56pevFn8qeBpRkyo0gGiviL+W5zo3HmaKrvZ+E74zIIo24QY4fbraNtu2BjyYs4
cKSA1WGN2qKrx0DET2HOvZZLZWvbYW7sOETPbays35mHY8iDv/9SaDPDfg3XqmaJ
V8egmEqx2TrFUEOI4wkiFQsC4OlI3/38ObOMsz7q2mo4csBi4AcSV+vypHUZyHPQ
s0QV06vq7kGK+THYf9RNffeEi9O6zFq2SJx85ObkGbOjMZQ+39h6Y97AFh+ybvla
GbjfEZFVGHYMCMY5ShBxb2Kbni3AkA352VQPCmMYwMwLVOuJVUDW9upE/AhOkgAA
dpMINsml70qlJ4MW4UjaN4jzgcoddf2ZTG9CRI2J3qODFz2jYkR21QcFrOEtqBbb
xhVJQ92a3NTNmlftEzKw5HJW0Oy4iF0Jlk3YixUf4PqrkjXVMWh3uGbenHCO9s0z
nUk3rmn1kAduuB4tSul/xb9+pdYsJyIRJV0hA7W457JlbCV8SVuoBlhIwFazskQf
odNK7TRV6xC5qwisQAlO5GnciJr2R2F8hmnGtHJ5mVdlZDoR1OFavG8dNCsQqnWf
X3D9YbHvyqtIpTKnb1oDluGdvSQBuYHOcPq9Ei/fofa4OH1cxZ2Bz5UR3qCDFhvU
4QRXyg7rqhf1BYup7A32hmodpbswf1/1+ctc7WhHh9CuHhQ4yBpEdyW4ykVoJYYS
+Al482dJA4/FmWCkkTVI4YWBK2+KX77RoQgr+Ht7yA0Atm5gfH5Z+khcYUomsBrF
TzosEbvxH0dAtetzB3qlxYKiEfE7SUo2hdasrPxuGpqVkColdy1ZTFBcRgR/wreI
tRNkSmiRGxzmwtEpftc1J1Xq4AqatvGBfH4FufJrQyzN0GQ5Hfbg1g0CaJZJSHEj
5NYlT8b4oExrDIe8d2ZUZlSLdQGeSC+hcd/3ssgRRcKJseic09z2AvlnQU5RdsJ9
nudFQfhyFR+J4lu/W7Rmws621URnO0EA/Skh4TqDQIoFAjY2Txhpxn0X40IFVWCu
EmQ7W4CwG34yrAOoVY6XG+5dglSwMYQ9CBOWCaLTVvojqZ3dSRX64R3fnuVzcOpG
D4pIbroALN1WQaLd1l7cNJYqxJiOlwn7cmTniLjEO79C6osEkTwlt2yer3hyOi4M
lG5VtyI7ALyXxqNVn/kjhIsqMI+YJPwQ/GAd9ZP3FIzunf+032J/HMhtBFXt95dL
nrvBpzlR0WrKdrDVJ/pz8heq1Nzu9hxUDn/KhSsGAKSqT5xCtiE1mBefkkk/x6kA
y5HCsAi2ffXqUJJRitgqEkibHvFwkuhhw7n0rzDBhgKh1dZ8pyIQ8v9wLlLGDnzf
aGfh+gHBDszcAlHJnJ2LzZO0FLXyBAO6mRLkBt8ISoUIwx//h12VgKQUHB0chkvJ
ZI7xpFk1rmCh811LFJLqvIQ6hzww2dWjwJgUj3JSbsoe58l3Q/4Xx/tsDwcWjnwU
R2DkykPVlEBQL9IH0QTkkG9bKze4BmdPSEXhCS5BpnuncvBCQHALzuej9/end5cA
24dCJkMa6mFEBAMA+Ochu7eQYemxZnR1ttxmgOq8oef1NFpHfLjbQyHHeraBAEJB
1lHJnbHxoBA3FXBNEz9tPizPZFKwcqoHGAY21SrZPPLIie9CdTB7ZXFyZvXviDy5
hB9VT5dblJgCSahgB+QDhGSRrSLwis3ai/SZ395z5x0letZ/vc11rOgfkYKQgKeE
tQMu4gWDkfVG8CO8y/jyEd1wmgDKB2o8bnGLYbkDfUeTAnTlj1gJ+OVZ28OrDKB8
DI1BbxuiK9t88SpI1+nOGjq1owQI04wVlcumZ0LgzQ/lb4y/FhghulB4osIqtXAV
UV+44CiouHZLVhAlTaGidYHlGwuzJRh7/UL6mXZH0p/M1ci+fVnETewKNKqjXeDa
Iggt6ARKHIMIaGHXxGcqvkqmprfNgOFBZ+5Tr0bfI+ug10eU+2ERa0KDFP/7O3Xl
f8bzjI7Hosj7jxO8p+pCIoZ7jWk8wNBWGmb6pFjvINU3EEJPMO2FPNqZ8L3suMdf
27RKAHfv7Cshc7G6E4c5xRJjxMNZBpWvB7rAKwtgXadQP+QsqApQJpbt+rxsnLmr
2J8I4J+0eTq1922hGQ3qMUwnlWgd6pIt24u2AUpU35Xu7xYvjfMFsFbBghmd1WK+
bDwu4Kp0TLpYkBQw6Ag3OfFEC4ftcOxqdiD+7z26r+ifhC6d5whYHpPqomrepS2f
tnXkFGn1QHqQdL6a6w93uE9I5NG1/uY83bPdCPpZs4c6wbHvPi/mthPxyyW9fR5/
D+GwnLeav/qB/4ZFR4Oweu16jSLJoJi3QH28nwmATtg9gfDV6wAlXfzh616S4N9z
ZKDRdz9xr6xml/93rRJIGARBqBRRHAYL2alug1CQdeaZzBRZ24lFh1OZtbM20zIw
7oKQ3Q6+DgzTSXVtIge+lfEF4O84NUNY2pkjZa5TI5Mn+Cz3hyHrdlIBubfkTpz4
ltvEdc0iEEHbPf4Zk9UDyn9HmSC7EiqhIq9r5X1Pv0TXtuwe0kIX61HIq5r08gps
ZH92Jstro4IbwIeWk94g5YTgZJMGETI+cWFKRKaGvvVZnoxEsPCRwJFIWbyN+kTA
+ofDw4dVWr3p3+fNAt+gBOArE4M8nkJTTjC0Mar+MAWCWaMVl2LXVSLKv89Zwn6a
pw0K6pLy3OcTkHSomBGkYgiOtx7Sx8nVMqw0Ygcx4ALkgREbjMhU+6l1aKir2ZjJ
J1qbDx8bl+BugN8WuAUSl+OR/fmucgYaRjwmWK6Y18BuQSBxoVu3zV6jdymxcJuR
zONV1FDxCKMcfpQEwGt7x+1Kmg5sqwd/fRMBGJV2my4Klary5k1a+9x/MmlOhCzM
hdHH4F/attf7YhmQwQnwfgbnYfb8pA+6shhvvQiD3NIttI+Ebak4NUuJ3KTPqMdS
jSknxdXfrrGiDTguJGKwWGzgp0i2OcW+T9YIEYJhqTt4fpQderN+QE3YMBkS7vRE
BtBcvPKlbRDzbDmsXOObRoXCR4JHt76qh5S3U8lmuCkGC828GxoLTKMa34G0XwPZ
r30T3cvSteQw4srO1M4x+QJEcyucO67pEZZJDnuteyuqBeaDzyOrgBaDLhvuZ1Cd
43QYbMmGbWFq0DGmhr8225NYa+6/TkeYJ5WXRh6BEWZi0Od4h4MCsoGb1VLcpcC5
Vwiy72R+oNLtdXmsswZwwYxtVzeuBbjXwTb3ouNPV6zBZiqxpXiGMhXlt1wcksrq
uqn7DBgbKOyEORI6NRZmlgMuuCnbxjiKebrDcvwnHHY+wLoJIlIIzmwc+dYBsJPV
dLrUb8nXOIsqBX2LP+cWntPvd7Bk9NLAeH6uzdhehw4l2GKvhsl/lIHoXRMD1+Rl
u1QEO60O6TeHBZgjFWgpfkEA1N1GTNcqu5m0gFAKJAcaVMHJWZ13VwOh/fWqMwo2
p7clExKQFNQo23+CaRA6Tw1pEij2yPhoqUe+Pcie2fzngTU7AwZx/dAE5Te3Em+P
EYijfmDcQhtr1GSFjN8gCnp/zR7/6b9tvHCHwgAjkg3cGu2x/e39HAY19AMkOaPB
2L/c/9EqUF0AAIDSDmXIF8pkA8NHG6couIjiEfIN8zT8ypNlWNzA3r7H8xMriVto
+QpumDMH/y/NxGjWrC4cylW9g8SkBaz8KdBjtXkU0F63hkYuYSEGqGDtsI8KQcwF
shB55/arOuzssAYURSytnv50bi7TlYymvRavehgq6sICqfmjQVT95Pfm+UVMSt+F
lOFmIUALimGhyk1aaZxnnoaoRV2Ux5V09ZZIB+To0zjMs7dglWnpskmC0omqekPq
ESoTevfBzizu0YTdyNzH3vnPAdIMjO6JC6rq7JkP8syhycDm4c2XhXF441KvbCiV
AzJ+j93QejqI8OhPpAYQtzMNk51yqMh0O5n7xGn3WWlAyPVpas2+wrEmoT6MVDoe
N5DIw2qIc1N7gyiaxW63h/2hl16ipqLT0kBC5AjkIx+0nZyUrhGg0FjSe/JboQjL
Xv37kWvXO0VwXo5HmLrEGA7qI/YdcEQEddNNSR61p+9HY6TFKxSidUHBTJNciwE/
NN346v1xpW1jX7CgWPky3l8qPx1YXzKws0p3YIQ4UC/iMBi64JKGAd0XvE4L3kqb
ai4w4yRW5sWrcxrbA+giJyXXuZGBc8NuKXNSxN8lb4OFc1eMklDNz4Q4dRPRhnKr
kg0VWJrTQ/fFMPAIdTpjE4qNP/H352vgc81xprbyaxUR32yXESChE8pNkSr2jCzt
acKNeVVbcL+sMxlFUorhLLhmsWuNTxrlvUIAZi2V5tlb7tHOc5KJxxcKc6idksNP
s3W2fbZm86bCVVq6IYDuYxIehnwDPXI+5saq8TqGmyYxwLQqcpxOPKAslsO7MBAS
Ped2Hh7URyWn9isYZLIYxMYYPFWWiaBbgz+mu1C55oT/kNCDVBK1Q69fqUFGpzW/
1VlHfHgY3O4ur0+/MeK+/RX9t6bGyTmRmL259tSo3jzasvXpbYUxyNOsvmue39kM
YHiTCOCy4dv3MIv82/7Ebbwu5qZ5YVDyol3d0Im2V2uZZl9hJcasLTl5XxpiAYMt
aKTcsTSx6/SabvJykVChgKYSCiE3en5YzNav2U5eXXMAr0QJ1/9flL7MvVTs4oOn
22OI0G8EWypJrgyA549axyuQEIRAZS0+X6DXNqznmqpYMzdrAeBu9mu+Jg/oR7fE
meLd3TbwHAAGbsO3vAka+t2X5GGzQSKLKqeEEBeX4+CIdYhBP7ULg0h6L6rBN0b0
NK7xQfx5qLMm7c3chOrL3Qytqc+3yL4IWBF6DdB76Q7k2Cg20Qh2TrTzKMZmyTSx
DNrMjtN6k70temI47ccQnPCh3KtiywXR+0nz5W7u1ejRlRVMUCWmI36BUkoRgIuc
WLe1XWJ/Dv0UFIGr00HuoQEh8iqgFrMYGrxgx9y88U8fgkpRfJNVV3Tk5q7Bka8X
9qp5Ua/txBa0S60eu1QuL621yudZHqjXCshLR9M9ZoBeSjx2iPB8BfgnHq9ZnTEH
P0T4TQLceK8ekShz/8/+hA8PW7HrOLwmVJ2zn/eFV9G8rW44dCqZ1f413lhdJ2Xh
BphXMUdZcTM3k108u6YjiCZS/zmEAJnyzkPx4uTLmg4GvKEfPQ7JvCT0DvUViuMx
2wNskV05sybwxO2Kk8uBFXn9dWWmugLBLwJ9sC3vQeu9cboVMVeDwRe7HqpZagIE
UNzaOnsImUrrpzvFbQXLAj+UTDEu8q7jbYJAzl4kWiOVb0iSi6D31Z1P32GyAjAo
QCiEBVhPqtr8BtQhkKAcVYQuVUcfqikx7f4qwzxWGS9MpUf1j5a2uegAS1TgWcPj
VcLdjRWRQ6PCzZm6WAjVHueP7sHGNzst1j/F6CbgC7X7VXKPiRvSoC691ub6pGCI
7axNx9aWX2PDrfCNMREMjS01L10jWmQlBojiVQfEJ+++kJYVgsaDhq3DP/mLUAf1
/hRceRhK+H9qGjWgiCt9jdFXFdf2QjhN/4HSVdYrVyT6AMwCU5cGrPvpb7hJkxIB
sG65DdnHwsEL9AYTy3BHKe1eMuex0SIeMjY3J6KpERtUq2F7K9whkK0+md1XkD/h
qiaflWA0SIZ7cm0CKFUMiQzTJl4/xWv8w0AQ/tu7ay1uQHazn6bm+vbedhtkDCrH
aRAKZqpCf0pkNQNltIkl+RGbdPHKTvdd+NpUrZ+lXvJbNJS83xqAMz/IjsfuZN0p
WAZvvHJs+Eg0/cZwJdHA4bVhsHeyFtWBXgym/hijYYH7llvhYhWxhK8XpRX1RwUB
qbrjbdlQA/qaOJDq0Auf/U1gg8S7Z36dDiiqmHm4ib1c3LzqPQFsS3Ikp7pjKwaI
ChfjHh9zo3mlNBeqZ2bZIZ5GyrCp7cFAU9VgOixuBs/WoQtwE813LI7LNFvOXSi4
PKHUyCGzsgys6Zp1ILKX/0LzbGGHpfGmZiNqCfMJY/Lp4WMuBcQyNmZWhI4aZ0pl
kpsONvFuvI81CWoFAH/5jIxoYAh5uHH+yx7Md2BEQ7fnVjLGAtTe1qIcM/btaLje
Uy+qPdEHbtF/W54s6ZX7ZSGx2yCIWGl3pNEgZFiceHOqo8nHGi33k5boGpdmp2Ig
OlWB3XLZ7P4DC5XlVi4FrUaCbAojvOxYEj2ODOpO1N18ue1yxDw73UXkqH+DUsbf
aa4OB3wL0M7nyLo0a2VOlZR6V6R6Nkzqne0xUC6oYJ3lJasRc6XyjfrjNk/FEl2f
Xd8DJ1xWXQErGcGcLfQmq0lePbAkLpfLUe4Y8R7QpchNgyOmhWRgv7wQ+w/cd3/c
Xt/iJDDVqe+nNITy9TFOyVs2XSpmPgMXNBp1jmmqsTRp0PgImvWi42DTOb313bqx
3QsjPAcxR80hsLcgE1vV95KdA7lBPlsVQHKLszJmycljWIKocBrReg5KM/WI9cWT
akby0mq9uxBu6A3Jg5s7roFiCCT+5hUroRQ5ZW+H3fR9oRJoQu2np/oqOU4rF4P0
pkP1cR/UKBjZxbHopdj22ocfaVKe13ovq2/hSI0aQGkHi0QmauIqxpxkwKAoHZUD
OlctLkR2PelR8ukhITYPjk7QyJNFWLqPztwUXPYfn8jun1ElZlz7YHxC3ASAxjba
nqEyEJkFBnxg76wWlspJu/S22+ywgPT/JrJwRtCbQgLUW7LHNJLXGFjGnxPQNAfk
31xTgLEpGRg1c9cErqrq8ultgtKA7g9Vh8HOCkayW6G81/dXmOZe/VZcUtA1jLiM
cu1xNQrP3jvXLaHDX1rrMjqCoCHEAGG3AaeUapMfxDEuYMJX5PJ3/pYHhQ1nsN9O
8gj1XKbR7Yt5vL7AeiYAYhlgEfYRX+NQ4ZZ+fAU6upm/ZZI/PB/LHtKNmxDiHoRN
/x2JnJECg6GJpNWfFStTkOBDo8kKQq9yQ+/Oqd2N7POnez2eRFv0VYku61wr2LLY
6QfI0igWCggdZA2kocEvpaI27hvUWP2a+yhQFp2FcyTZID/CPx7n4827XTrKVCDc
3ggmV2wTcR4ByBYDpEgKUAjJek8G/jucvMUXWCm1oH2E7UScaHgwYdYKkFRPY1ce
ac2RsvCKSfOykFHUeEAT0ZeiusP1quxvb59XC0xrpoDLhtohCGRfy+aLPGJ+y2Kb
0MvOLD62OtGSaMMxHcbN9wrwB1hRR1XIDx1fGWHZYauZWSC0ZHGkxxZg8EfXKGKl
XoOWtIYMr7m8OJ6KqupTTjaTvFz4SYDKdwQmTAlhyK2WDwyJXwtfTFcra8ipON6h
o9BBPKZwapBSos7Bf1vMihw9jpiE0xAwif/nmb5BUCy1m0Ku582GMeZvpwL93xA9
rJDb3MRNLAbdS8VnmeqzBOzQSDvIdZoO9o31d2qkfFFXlqi3dTKBVkTqQ05oJMUl
AwtZYc25paRZdcnBXerjY+Qt1L0mdGBwgWOG3PDbHZNVuQyMrKonGS1rAkIHhxBt
gnBUXH36tEuhAaIGUNxFwDTiDBBFqZ0N8wG9xhYj0pp8HOM+w0g/tYuLVVlsYDnX
vT+aWJVkaqESYbTOJarkzyOgadyXmquHZgnbWWBIP38mvpwyKAHWYU3LJ0+IoGrU
8eO0zj8JzJUymtDCV2ZYQ+6fZV5bcwX1BbtxXQNcl4JsrAt+LSVEbajexeu/LAvb
W1tiEDp/WcHPzSFEGsOfuN8FNKcx/7K4Sv0ZI6oVAXfDBp/y0ZBFEmPyq0ngPlQj
Yc08UuK/uRI9CQyMOushvX/D/0sjPH4b/mMwWYOd5SWiVt/3KrGBTdyX/GXiewWG
D2z0+JKXmqwIlszEUqz4B7u3FMvhmoOgHvAKgJeuisgp7j9p4cVMG21l4qi00Ifa
uvTgHP5qEuxIgCkkXPYMt+n70DJpX275GAJ2itKIrHV7nGhVO3g4bme/gzL29/3U
RWvu/4BrwIvROqBz+ikwU7VL5s37fYKL4hvj3NHnij+OWzPbkgpeyZ/Ia0Aj+9Iy
iNCXZBPt588cahEBsHhfUnKFMWELXtXnzggLFP9g2nHQhqtrfaIlPc8Zjz8aZVgZ
BuzdJJV7wu7uSqsdldealo8ZDjbltSj38t47b6yYqyes9cWLCjNHmPAE5V1D/MtL
nGz0D0u+rRxOZPfdilJr0P1hrb+m1nqTbaq8VrW9Gvni6ZMIQi7Up2StrSYZlHRt
psaSpG8YYQ25e+PaonJ6EzFiYLuTOX8KKoyZ7ajyjzykWX5hkS4AX9h7SwJMyocQ
5YAoKei5GEKCX1QrHJ1F4qadkHuDLuYEZaVq1YCfBVK+U60SA6z564qBPF8hYqBs
cANLS5gfgWBfUWpoWVyKZcIpkATQehdYpO5ZaTptriw2CqfdbpySR/aY4f2wAlbK
06JGuoLUX98E8K27mgohkyOLhgGvPFx4R4CFdEfrFFN/ToRwTapIyYpIZcqqDF/M
o687R/4kl3Epim9Phffg+JSazoy8zpbx0TAZBM1EB4k31Vz8+BOB9a9mq+zOLLWJ
24v8C1VEczsT9wXMUQQavZjx4Va5mTzqoKad7+EvKpvYfpxKA6W1TrnHMTZCb7xB
Ha17WMmdQpKTU41V1HdmXMnMpJa7mx45yVyBxYMDKJQb//23EhqX8hRTcIl1PWn3
xzTlMq6vOfQMdvGH0TOwsjA+9TuaNYC415X0Kmnt0wwm9rvcducgHFhaFQ1w1JJG
X+8PuY8Hh2/eiwkevHnGATpBPzq9C3IOZkGJjWixrbPafViJmJJl5srE+MYdGCB0
ldj3krAy1MTeGi0/vTQHN7X3cqwX5RJBeKZvIRqil0fnCy8QA7HqdcEk2HabWymr
gZmBpoQn0teOqV4PiUAOihrdU80IVTsYJXRrl8ARA5e6nY6qHUlF5lc+EXKh6mDO
xz6mIq6yJ/18SDMw+CwR1/qgR7KH2qsHLFyqT4s/otOqFbrBIZg7O5H5lkQkD2MP
YfLFtH6Sbh7C8tC5mJhDCYRUz7XwZGGWCLBAPu42aPV+Z7xPVszfCdG6z6rQUZDZ
pc2ZoUd7EzZRbd8NOo61bv6vtS1vT2Y+QZ33GtlDucN6sWkGNmvT3CPF7WnjxXZJ
7M6uIWlFzVwVzHiSqy1TWTBfnYc8d0VA7zeQIquxPsRo7E1f00oOmDghefXnh6QQ
5iueHuzpV38QrOMTMVJjEZpM6Txd433i2gECIhJGpCQAviTdt5IyQRspiPJvuT5S
ZgGYNi0R3Rg9IDIiRbbeap21DK3STZu5dkcGi+OtYygp7u/dceIAj/adj4/g3xjc
IoHt9FCMDtYqQlXJ6G9vhB+kxxTuu5xukFJp2ZuUZLEh7EZiQ06/FmaexRnnbvL5
R9vQVuFAzS5T2ZtcwBsd8yajjB0Fm+zXhaRon+XwIZDp+k61ZvIViBLIG32W9obW
RQA9hHTnxDglUj9deWEVCNzy09Qk1hn216XW0y56+0wdtEW6y0Uva6F9xdFhEHV6
sTHN/yV8De2sAqxTKUbrqjWkNFZexsfcmU79KDNPe79sXSqlafhd86V8ODPVWNiD
OOQVVv4T+CkHPDW4svxgJNCdIsyflEF6I3R17lO2IUK3p6ff8bvxU9N7qgWoC8IE
OJlFb3w/3b6cnNRYWAMxuWoDlNm40coKcG43T2AoOilFCxVt6wkJhXxMLvVysODq
yTaJbWEJUkjDqSx3JE2blUPHYSjiWgmSiu6rkg5BJCNNb5j0Rrd3R/RaLWmmd84G
C83GVKHfp/SF08KzUNe5liPwMikAgnyRZFKtH8fGfHj5GUbTMdp35KePAGAKMqOi
hRpuVnwEFxug9uckiPz01dpFUjF6zKv1SjB6s00Rw8diduecdWWh6YgvOImcEEo5
ybp3n72xnI8RU4dzE/5XjITu/MCuiYZH4znJOyuPybmyOhTrneAt2Z3EVC5HwnmZ
t2L/QwQ3NEyS46Rtg+cTg7Yl6QKNnFg5EMveCYUQKWEmkwa0k1GE2sPY08pz3K9k
AYfvq/+b5OgPS0HQXVwcywM6ibxZhQ2vldtl4CsxnZfCPwF2JB9V8pjqoCdYqv+M
uptBfv0sdjazsk9qW5q5yZB6za+oyyTl1OFC90Y2iVhXBqPqRpwhpsZQWm9lpZTL
SHm7RRzsj5dHbxfDzYtA/eWSFH0aDth5YPsW7wx+CSpNaa7jl6nj2uWOHUyNjCw+
vyPgwUYYpCXPAtPSkHRSH1kIbw7i6kaNfU38jMlUhaHhoqOcK/DgUcl0TFU0dP5F
1gff1idO+G2Nk6ccbXt/IN52cgdXiO4M9liwnPTXqutRmbE2UTRPdMwoPIKEEokN
BOgtxZ/lS+mcxCO8TIkaX+JZ6/QUDBiuO3Vww96N1eJmFQyocaZ+fznXmIPjsvyM
VgO4uj+2nCVleMoNJxgP87C6wpeg7vaBi7Yjg5st6sIUmiBPU6Yb0wcS/rRv2W4T
/yH33CoZITnbACfxPXVRrFa0rYQV1bH7kg2tfHiXDPzBdNs7fdk1eHU3I2tCApXv
tHiU/bGgJL3x9A4Iy4LH6O4sVbSeuUiS5fh+UYpucqRZ5xXUND8I1PKrJjxVj+ZF
O8v/OK89F7olX4Ouql/Qgxpmg8ntLIkUE5esgcIs642XRJdn//tIAUaeUIwuysjh
x/fWVQaUQ8i8/IsdJpHucCDiyljoz0M5c+Hld9C0+zLFESPEvYH6DitfYZL1U1pC
fsj+ytCYV3YOQAMkIEogwC4ReW68IBv8gR9dYIjes9pkOKiY+Cpn6R94Cw3gVB++
k3UytikpYK2f/4r/XSyzPdb8MkOrRKYnSHgKTxtbts3TixpRPQ3vU8+fazV1leoQ
XnrlEAkSFwLf4ocNJ3vnCl/CDgWTx7Vwba03aNYF9tFqFETvvPEkMuyD1VP/qA1G
8QpIiYrMzM2d8X+KbO3BoEJ3mxh2xNpq8qQ6QQr5qGuRvP3O6MGwOymmT/lNwEIS
fPZ3s8GrEx6D+CEJ62b5zeV9fI79rD7Cn61EPz48886dkFWg5GIIhJ4tolb/ZDiO
WlHPwBVG0NGZ3t2S277+IcCHo27u0D5qVA7s+UiDLhgnrnLSKbg9muWQdWFP0l9a
W4EN7Ih3XWznqRWRHvKQP17H/kzD+UHn6wrjnyL0L1jqXCmDSw3XGSouPtJesh4h
en5bPdCzasXxtEMTteBBwkRG11GacUmT/pLwVNnSbcX5VedkfHlJQlDW9SHghsOc
XT/OqEFJM7I9Aau2IjJvhOVmArV21C2QpnNw1ulXi8YNLP3VgVM75RBADJ9eb9jn
lcC1lUWqPbovB9CFWC19/ks1BgwJdcB4dd/J7mILv8Grwtg+B4dxeqFi4wRWCz0x
5GPF++SQLy8l35D3asw768/c1gZrRTLnvqkYz9aac7VcABsdA7sm62F7mZZh28vx
TxxWxDAkc5ZyTttPb7+iTcnoOBvre5ShpFGHykHvhi0b11h6fh04LapCubYTUnUV
1HOmgMPc1pTObsiGgKCgJfd0OoGHsRNd3WrqtvZtg1Og1tAkXeC9ZNIJ855BWJnZ
U2TAUn02r40oupko4AT3s61VXa3KbtBVS8Q+ucOqmc2ess28N5wRVaCxx5hckBi3
J4EdYSsX+AwIFFY0Jl23EQx1S+msDt1hnWAV7Ki1LfQeGySKvxCaGWd9cUQMLuH0
oYSciT1OEyVwxDUCDhyqxV0yzs2Bpl/bgiAGuuO1aiO+L9gmnF362Nm3WVKITm0w
qMhJMByI9CymvMR0gLS8/IoiTeYUD3jlJSKP9JXUzzmucL5H/fDRmzy3aaNgfrC5
D5HBHolMjD2yqfaupD3neewf6pKJ3r6w7BXzfvztYrSZaLHxtC/ENIFiyfdrVSzr
DHcVEc1kOFftaJYHMWXI8ZS2IL6x0lpb+Vi2nphWszwxu/OKvYWCvOZPqMOZ92xQ
8UEIF9ujWAKTF1Vv1hdm6+N+jjO+qxte/bso7vpySgh6kaeASdiijpE6RnjXpdhJ
kxvYWQwICLS1wjRT2xNJDzFvCc6XvpV8KNcprmdk232QBzqr0bUgf6sJN1374KQW
cLTg8MjsTcLtDcxdngijtIH91Kbby8cg1+XwRdXOMEdSH019rZvSOakGNcnXH6QN
6eFves4S2/mAZc/g0oJYJw0xRloaMmtD4G0JTAzgHleoDjBSC3EW8yY6PqFC3gR5
QWCwVbTI+zdNunOKO/C0vKHaISW2PW8kTLtaRoY7ieBqaOrWNUC92kQrpuTQ1/KE
+cspkhE9YUkCeJ/1r9sj+aoj17rGZV4NM8sszAsOWodrrIH5KVQP9YWEdZYpGRiq
5ONC+BZANBeWuLpjIgYS/+3RZZH2SvLAbZo649XAm4Y0e7yKrzz8oNFpIoMALsg6
+CZDI0gNTnC9KS+LAUetCCmjUsch8g2fy8iibwJFeqUpXZCqt/Hnljf2BMlPC8sT
X7UFHl7TEFqjY0UrWVZEj9Au5lpc04NlfgGljbEBDwT0raZUTEuctqyRz0/03Gq1
LHQBvEIw8qAC+6SErbkSzx4VRHZwmgbsNfHc3j4XfotNeYjDsZpJayA63b63cNVy
DP52rZYJEyR9uE3Ihe5suJWan2xQlB4bYJ7CtHC5UaScXkQACPQh9JZoXCie3ywG
3GquLIRTC8XkC/Z7s6wvUP0BIswoOQUVbaFyhzPNfuasTF8QkzIcB5f9NlVA4Cbi
Kh0bXK8cZW7bW+VsAinb7WZecv5t2ycpdWEa7VWIpeoCd7tzYvOyuC6LWVsqe/UD
Vq8b/4vlyDfEco+cpUUF6+SkjmPu4Hi6dFT4YjgmOzOB1eWjJ1JOsAQYMm7Owffx
UJ0ISFbJ2ZQ9NMAIpnHtIDPwiVtnHkKNlnZH1IAC32+8aZjfZTqQclo8vKlSJyhb
AjAJ/jd+N3SywwZaNF+ARESpqSqjRMhfxgNskbR5dxBbCrAyV5DsZwlVsk5c7FKf
lImFJrJLUjIsJyMUxLW4CFaeQAtNLu2W9TKImhF0CcL7d/Vzf4CETqL/clFDrumw
mIYPChR7IaFZvZafLgERvVz9o7q2A0PtPwESt8SW7l5SYiWoyccxioSTv90cVn6C
tQnUO6/17ynMDFgy9YRZjfGv0v8Elj2HQmTdOx4PHkGn5q2vBtiiTa9HmXZN8HCz
C3iqr1X7ncjNVb6xhdcCgkn84+yb/m1XNwACO8CxrN2xU77SDcJVviG6htH934HJ
ebBhsGEWzRhOJwfxV4dpeKY4Bv2MCXyiP/1D+/77H6Cl24eaorB+mIOYlA16SdAb
mJCk0dLCwR28IkEMbI9WSPiYt5KrVFKZwm9NMImDns/LifcZnzv/c3M7eoReaJjq
BKZgq8rsJlR2vs81EDQNv8gcSluS3PoE9oevwCc+SQGIfzYpHeFyUvXEOf8Fhr/V
8ff28ASyiMGmyJaLQKuQHT5Mmo3AjqUdPsqAkoQDDJtnJ03TpjnMrpOxSv3mz3de
I2aOTCAWkfCqDCInfEGVd7Nxbi6qNlcuDyqVtDKmGHdcQG+r0FHEcMj6KTFbOZ8b
zgHhH0SThixVM3FmGtiLdw+8tCWtnpQ3+ckamcFQBNXlKDILRF3fkk52boBKfL48
/tgVSfck1sD+Sam1/HEoB6mf8fHXKEn7tOKbTo2WsQbxjyFTOOQ3mOaNSZSeRFS+
46LgF2s0E+e1yPZsQzGtzZN0hH8s2Dl2NYIMqWI8c6fgdlEXFoeU0xh4Wowe/vgk
o6/0ET3PuEpTZKyGBCWXTtgkYWwPHEwi5nr83OZCnJaQdmuriqDknxtiv4Jkw7Hn
7+emv6dnL1rF7nE/4tD+F3H6HVMkTv4wEeqMvZEeufuB6u3GAXBzKnfQBBXVcB4p
3EyRAAyz+rf0GSGwp5lWL90gE/ggB3YmgK3qhybB5cbjWzY9fiMvcSg2ik8hFrgR
P/0JPbFCNMMG8sdPhF1cO3x1YBVbbT7EaIJ4yNmMDsV5H5cRj12+lmI2awBV5FsI
o4P+WVHLJS16GQYa3DzpHhCiFG5bPI+FheFYBOBCYU3S/FFJDoRELUDMAB2Ra5zu
vK6IhKmo7MD891oPfxG1sfuywV2dCEf+Xrh8IK4zVBZ/YB53TjzQ4o+eC1m5/wTL
TUyzGW80EUaptoKzD72MIQcWOLRHOIQQFOAGBq9W3iFUDnaJOcwGxYePnekupJOl
PzFm9nBmPNgYAsjY3/g8wYQPph5k27jdEXwap9PDZKVglBLd1qWaVgIMMfXn1MSE
/hBzHaqc+8cPJvY7AiRl8Jl8kNVbv3vQSFEcDBqeh+EnzFSTcxUwaRtZ/hOyUaHX
bSEcHY26BmP57tGgMDeMo93USrWrfGuQxX5pSgAflp3oSoISwC2qS00AEw0hr22g
04Mw3AesX+YfeWjgXFokULVQKwbQ1Uhyxq0lkpSks+OiwWfYDNcIqc1nJChO4o/+
Alp/lgR7NDrqP0mKeyhLmcxLrspJNH3Z9E6TL2lUGV8+PfqVHKDhLMzb6dhNYoyw
mYYxUOULnudDfFgG86BrNcgOi8MJZK5ficCZx/pffNRqWw/kBNvlH+Z+GrdnN/zV
9KTGXDwg7Qxx3Yk8wKw9Ri5CElBIPsz624UQjsrMG/CpqT/2+Zleec0dy+552Iuv
bJe6KhA0hOodQcPxPMk+VHTptNhZ2POADAZ44GA8HUzv4cfwxWDcXm1lxO2Qwz54
p0a4810Qq0GLHYDgkzlB4A+v0u4VwMUQ3B2PD6jsGjXC4DYJ6FwGzbeSyuqyd3vq
gSpOsAuDER7uTa4fb0f3j5O9udrbWzh4lySRxqdUmgKiJ8Gx3WRiuXyKjOgUuD7n
gtxLxNxmYqFPoo33wxetKIHArwtfT5+Ba9TViLxnwp5dHPcg0f+Pi2hyNhTvUGAH
HVf6IFEPlnwdZL5LRPJp10NLTdKNsIgjUjCXMh/iXd5VMH/45EBWCLa6ikQHQm0l
AfslJYCcj5qW8OGckecHRKIF6EwC4Ud3UpVd/LGG9TKB5vMtt4Q72JFweV7/n4zA
KQZ8RMi2b9IDuzLgwYrbvstHQZOwMCTvXY29A7gx+6qXtSop7H+JBrltdyi2WTxs
QBNDi0bfjDV6Bv76IRyMSoirQChAbvlodnvndIJFjag2xRHYDm/NOU4/wehsiUw6
Vbe+TiiXRjFiNSNVmXBiRisF/+lyXyvWbzmvKbaZDX8wnOeU2C7Uz/wYHzqo2D1B
JTki6MuAkYQ7gOYNeG7Tswz3+j/N+lp+FZRWN9mOhtlIz9/FgQDtKokb4ItGJ4PC
cmwiPCHllF5tm+SFOgyeZzRVna1GEXayZN3DFg2NcjgCAKDZ9VoMhtZrV/zjLhBw
e1kToD7nUm79tfPsqW3PPAwwFmB8zQMlk/1PAIvSWBay7kCPyU1X2JvIhriHu39Z
OEoTr1pEw2X5WaKCioO2BK79NnYylm1fOMQgs2xxlVwPzuh8gW0bm7wXK1vHmwIO
oY0bTiV+rbK1XLnJAqJBLV1BMJ2Vc+tWHXqD+hwuJAUn2Lc7d/HItTjMarvMEqCM
a1tu9YNKPyZ7Fualpwq6d2CVi7vJr0fEPscy4KhhFI5Mm2ua6yHGJ+syFSKgoiyh
cPaQ1gmL30tbix8cAR3k6jj6NL1VP1ntIgpgCOi5rFJou3OE1zKfleYhnc9aHcEh
WPQt63YbbpMj5WS2qR4j5pDbxkYxS9rHhOPpNSXdMkqq83VuYYVY7xbP5ElTVQvJ
XNWVXvnF7PCE21dfTsXnRBSE1GXfe+mMdOtyEBW8H1uM+fMpzU9AUPigZMYInj1i
04AMmfGHLo26D2cqPEou/PX4/EQwshko7t1NGsvLgNHuHt1wLHvCIGfimyFJsdI0
/QGDWuZuKDEW3cFEkUw9NdS8kuPkHifvtVYMyMnQJK7KqTCpLzvsHPE+ZWSphXDl
9xp3AwrZ4YA9gqlcorARnICLtkaRthWSAmpUU/Oa9hn1UURlLdE0TWJUGaybUtQY
QJeyzH1EI94wQTUAiEScE0HV6iqb4wxgOJbZ7bKJpokJDLNl3KuV3+4TYHhTlBqm
7u3IdpC+JXxqXsz3J++9/z/6jcBGy+o3ssScWUX6o9+c3x/D9wXwtbuTSuYlCEKM
+0A9PkgaKIZLZNX357e2ltp3oGaReAOYjfiQEQjXXiKKNgoQS7+s658MQBHmN058
CfWabjyIeSWumlQFRMQjl3TTbnytqphbeXOS4/381jJAWZpKN8OIXbpBezqYIcDu
7GtFDGvw5GrQNF8tGnJyeNDo4xGFE8GXPfpGNVz3Csvy6QjtNpw5b4dl3X89aCTi
Vl6QXlpLCHsKkk3aIQUcxPFgM9KEgGJIqcmzOy+TWUsgDSzcCUhoHmcd3BolmpAy
nDmrGLdQfVKINips4PK/KSLPmC1OI21Weo7T7yOYmBGmh4FAScKq5aSl4l9H1jRv
GI9ZI+WK1xHZgInQ2v9j9pe3hSe2oxhJNuPQzo7e0Cd6knSnBXQ5Y0En8FLbPZV2
Wi+oMqKXo6V/mLWyzsWVNZC8BlVgisf09EJZ6v/umE1OznO3eGbILwJpwkXokV0X
zB3Xc85iTg+ITzlwsF7PPIjAcM5MFZz3z8OCjG/i1ayFMtYvweehABNyDn6HgdJl
0nyVYm3cgBg8SWwMiCQ+f3NmJ5VFvzXMdXFgSFuuGJKFDqqnefFKMRanXI9KR7h0
SQ/B1UYt2zw0mp+Oit8//BFfo9bzIZiPMg/SCy66IxRUZqO6o814Yu2Xuy9owXWY
i1kaprO4HkIR6G9u342K9XrCnw8t9ZZOSDYhbtkLhGtvkMJY24TTcQvzDtI8IsaA
98YwSGdGKRkhQ7GLzUYGQ2J5jovJ1UlNb0NhTxotKpQFt0o/7KtTux91f+2a2WS5
hQgaPnhh3JcKzKfA1D2zWFcLS5bYBolYECSQ41ouiTNtYom6V5zfgXjj8+vkF5E/
RuRFxgi3SOBN1RKewOJbPASac4ArnrGKjyLXOBylRJhLm3ZSH+SHNVJ8Fa1s+70m
SisyYbwP9H8uV8UR//Kg2LLadPHJ5f9nx/KZPun8ZD2Hla4vwny62aIj9O+g7082
+TqYHJXWL5jaOZIGpXIy5sz9fNXLFkdS7irSzlpcTq49NN1mYIA47KWXqi5Bdv5v
uCjzNU5UZXLdn3Sk4z6Ry+FOYSAfvp9yql3ixjP9Yd6zK5e/IqPr8ocrICTogSxP
TmbyM0l4rdWkjfgN/ThRI+46hLHZz02tlzn/VP/nwr1HaPtFQ995Od6KDZDS7PhS
duX67ClSW5uoUnV63KAX+i+alVJV/XeyBq7SQ9rE7CH8kU5rsvfh+lxS/DSNJHLb
50ftuWcMhAsTy7e7qrUg6QLBCzgWjhfgatid6WkqyI1ucWOR8cXFYQN82SpExN5u
NygYg7TwKmNHn0qTr3wOgbkpdCF6HzDDR1mGH92YhtIDSAzPWK8whsgKYTrpnnEK
m/8MctE1Z5oNbuR+vU7fZODrWGLaW8yYcFw3Z7N8GsFAbEMFNi9YVM/zkb51mnVD
Ger8uHTtlIfUVJgoNKqRZhLJ8RvJHt9Ik2IbGzMR/sSdA/fNDEruZhGpk9x6soW1
UWGRIpz5Sidk8tlgQ0AUeliT7cUlK0oflrNdZjMDY0+XZt2J/dPDbCpbP+dbNre4
vADirpn2AcKbgVZzAN3vgXuudGhOMugB1dmwkk88pZD/SPmE++LeMTgenO4Zmuhx
6XPfb96llGv1gXWewsIjw8mUDa9K0n5MRrSZvPEFz9RyMXkgMqKeUfTCB+7wWEas
JShRaQd7c5D6Ol9yIgrAELCecOCMXJ+zV1v41OlhFZllXAjtY2/Ccu+YNvzSD4qp
0st7rP/2DQQig03j41FQQ44P2IxQnxCbLv8EwODoq0THT9yaD4yh3xAAT4xajR+3
vPXc8EhUVE7sziPPyUPvf3LdD+tJVB1ytqE5+SPjIDoaVSX/ySw/yTGXZlXAd5+F
RgDKbluXwnKKUpe1Pe2ZO8XkHDqknM/l9nwK0YnzupqXi1LEIbW09S5MM2QWDk+J
Cl7nrqI2cKC2uJf/inrWL6JY8dJQ8oSppi+UQQY8d70OPrJutu7s9Lo7OnAAdKAX
Q6gNeu42RCJWYTdiD62V/IGss8OoHHLv/cG13GzSHywTj5I1X7qX39nZ5L8FLyAn
L2DGfFvKAu7kzny98U+bXkIQud5ybfvxM9d18U7EfezzkO02akCViqlRYnmuPymd
xnOUE3xdjW6aNcPlAGIb8zsGYNr8xgJCnhb6IzqkSb8J/e8mpm/AwscCbn6coRVh
4+XA4meg1s8a4sDoaaTzNW3Igl0kWEDjwapyfNbeg/bStLjUt2Y3wgTl8J2Bh2+W
j3ksdCrjnWRmsNxrjyWjKpUZ+emtOL5r1b1nFgf2pZ9Eq3TArpI2eVr8TcbJ3P5K
mSpJ1HkXEF+KZ23LtHix2Z6VTskMWVknGOaWNiJQ6mPJSZs4gRxelB8MHhR95tD2
7tcQQkEvHjYexKLKJbdvrHbzBYyUjVQMXZW9SugKCB6ywZvNJtp9uXfkgKr+rnyB
Gf0ADLhSuIyeXuuoYNKJaNO8RWuPA0ucOEawXlz7oYkpOFHJ+4NsYmPHTaQUrZ5d
VssRpFbTgV0RUzKtmXMYN0IUTZdQIgLligZBF9Sc+3sTxjCZ3dBcTbd7aCfXq0pK
ZThujoL6ePT6ZXAfhXtY7/+I+S+SjoJagr+ojkZBRjy8yAda97kOXN7aWsDXa+rL
ilErWixtTgk7vDaJMqMMHxSLwNRUNg0Zbc06Dv6dcvEIhj8ElEN+i6eEdJRWMPAX
1aY0XF8SnAeV5vD5SDWGNAaYtToGeyyi0oigolHtpw6ASyN2tskzYGouWO6whu9y
fS7N+NECtGbUy8eNzms5/94b66mxMRJX1fd0z6KSJggGjTqiAov2hMQy1c9jrxkp
K0JQSRCMLIRtixB7FLDIfFjpYlakD8qccz3GdLBwgE3HPrulEqbHgiHqn/kIR9sA
4ZpVerOj1dPkU1rwxPSlfqinpI4dJ4iUzfr1vuhS3sfIk7sYd7a7CDbLqqUgj8I/
pA/0TOCmuiAu1zkGKhUTunLYzFnsAzV/824dCLy1G7jbdyEGTc1oz9exe+J9Uhk6
vft1P8N+N9pDvmiFVpYgxsd6D4rsPj+cxXOb9k3UhE/o/TeOUyDwi3Q0e+fI3izC
nMiS5soohPaYQmjzCRdicmB6sBjqUdPRXuip6Qn7sU119VulUbUXeZlWwjwo90iC
9hqIhBke/Vy/SMi4q+S0tbgITE2W1+VMM/sHSZFm06QsnHqnK9YQ7ol66e9F+qHQ
zVR5P3X7CzQYQD0BKFyLqzLddnmHZvLs7tgpRUT4W3jye7Ng/g8kD1xgZPqWc/cn
vw8wJhIjW68v10MWjVZJNw1Y836GWya+OgyXrIQZR8gtQPvOUkgR5HAQAZChjg6Y
8TzqS4XEiREuBaBQCPdpr3OtylLEGItGvEv2ah41RPO+GlMhwxbpne55n7THH7uF
VmS8m8sFpnwMv1TmXTcWvXaKc9Bxq0HHhgkHyzInCcnuEbna+e+umi0fP3oyOhDm
5fFYV6DKwwYfLN/OX1S+JISos1clRoGDQBupW1qvBICTvF3XeAtCQViezQ9R23Sj
pIgK/BOSVuH7D7svOOOpEF9qtttpvWa6138aB98+Md6kqwoIYApZWFjrtYZnhU88
UcdhTQVP472IPQD//XxEM+bDZPYi6e8nlk0SCBagrRP/0A24vFD0vTkclBxZQoka
NLxC7Ny7qklTqRgyvYVEE9HAeG1wbL3v5TI8WntP72by5z62IPDgls9bnF92sPpX
WwfRf1sTUlAUptdoITwGEnWuIqxS8sDNhowwFV2tz7PVVvRsTnE06dTnS43v2kmL
Xh0odWL48Ho95EcPZqOhL6FcNsPPSHy6Pj3hbfhxlyUyAaiUCGbDT5AI7csDBZyp
EFHp3vJrGECan+zudtY6f3Xv71mIHLNNYzb0w9k3TnPqY7lQz5BschuxZmZW1bIo
SguCefC8Ncyz7pyYfVsMfRuxAYcOYYLSQ2m+aC+6nZd1kxliXjV45H7Iy5/g4Uom
OWr2mDAz58o+OAw/5nWgpSadeZlUedST77VHkQHFBEyz2AMzuK/ngIvR9SOj1wxy
DCcZ226mf5pHvTfJdzHiC9GyHICypXFw47EBEQl+iaAWGYRD/BOgJEfxTWWW7CiL
wiqLr12gCIJSHPtm78myv6CzwdgemZpsM1fDrn81bJ0bC382tn9z9M8ihXJXcbPs
4Nam342cxfkLu7bRRKwe58RkNAGdcMJmiSxQqLUh2a+eLVEzTvaPBgaKCEg7ZESG
DWvALRTzUfBqcYX9qj5m5ncCYaCuPi19XcwbN80pnL3K4YqeEvAU7q33GAqcxylc
yIFFOS6cEWFqY5SpJNy2wO9NWmTQxRKUPi7BLqfdoiEdXw4tE2ftkmBX9drGILxC
Ibmt8AQqHvJkX0mByv5FAe5smq/we0Pfkn4xFqQ+cJacnEzQr/QRij/VNV0Sq5Vg
CgG2qBO4gueYpJbCmxDxnG6FJL4tXxzErtXUElLJMM9sGNxGTLciLi/z/gmcqeo2
JX/IFVrpnLL0ut7QlvEY02unn/ZjJdLEasi/67c1y+BQ5eOCn+KN6aBz8sN71hK7
3FLf/1Opgj8LGRymou9FjNkjZje7pQzNAmxz8O0OWh48mEwDrj0qoPRVoS1GvFZi
GJ7fqbAssvljJ+FAYjsviU0l+3Q2LQYEJIoAjctPubVGyzIuf/5C2FJiNwuUc2dl
Ak/jRA58Lb8q+fDaU9WL+VXY1W3LvWxWKyWOnObeTWB7U8yEqY1dZxK7Kdub0KD9
EmqYzdUuUGmEjrVh7bjXRDPys95M6xaSWmLP0txE3SDxiSCc+jQUhEfNafmSDO5Z

//pragma protect end_data_block
//pragma protect digest_block
1XYIEwZGSFza+SUScm6Ee24AZyI=
//pragma protect end_digest_block
//pragma protect end_protected
