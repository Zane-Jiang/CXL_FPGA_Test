// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
jj0W5IfZYHbqBOgY3w1K2HuyfUB/0Dov/PqqzUqji0sOpPhi7AbiZgCuIJZNs5xhZvU2ifqOP5h/
yK+7sUo0t2pbT4Wphn9KhdCdTjLJGiCoj92XQCsBi938F6bnFtoQIO2DMCw+hz6VntQ+jI6wt6MP
nvQl1iJM0yB5q8I8IQ8LLbEqRdm5bcPAXwrunxS+mP/YlZA3LfEWttJLfLforrZS1qy1NABGqVxe
fYtMF95xp+AYIFcA4wzZvmdbpIJSVRT/578iFm5cGi4+CWpk91sxYyPcOJcv8txPXRLe/SFFSTnI
IC8QxF4/B2sjN360zBWClu2wku/ifDKPfTFPkQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11280)
Q3sVrIIo62Nb6iGIvkEXDJweMZ0apmqFQZd7YVSzbHT4e12S2qEU0/0VdWzt/vIZhIqlhztTLJbY
L5RHZra2AzI7KeN78tXWZ8G4BaNK00EkpmPGRkiyZACWD9p9wAU1/ZeYq0sQI2Wqn/u6kBDk7VR8
6hsmYE5uh/9YedzplrFQkZY8GE4/yglQwFHJrvoxDl4zp/9hSSs/7a//wuiEajhW+AlQmznHYEll
DHBT+FeA6WgIEz9ttyPN41OPazo08aTEJmLo5ovziFz4mzl4BTZKmcczBF+KiCi8Be4MIHoJh599
6wcls6jnEdrElCKxQ+cgtgO3WQBhpY8wnvczDauP4xtV2ljb6acuMzxwcEnVKZ+olS386Z1WJRZ1
wtIgyOooeIJaAls9uuXToOrF91nrz58boAHNqKetKqad5b3JZi+H5WOcL6SK1CZ0GfGl4EOutCPn
HkNdnOMAIGeC4qCOQP5JoyjPTk/k+uqxxLGuRDK8NHNPS3Go6AXvmYM/CwGXKUM/2VBTUDV/Fkja
TH7W5xex878w3wZJbNTn64Zvmo0A3i/SeUrwh1/SQdJDAmqX8rmBpMBCvoP8kf6zKkBc2QhIX+EA
SZJQ/P1Z4feBZKq0Mx37UoXLCIK60YQJyK6GnyimitIZ8qRhpa0GEPx8+RBBLV6UEG3ok1KA/0Xt
ocBBPn8YEZ2ThoWMZ5KSeEQG3dQM8Ddv5tvCc0fClR91NwQxHUnFO0YDyD1aLwLmv7YiqHHL/skJ
ngD53n4KQBgqy40qPrA1Rc5gNebWHn28VvKGg6KCJserAbdKo2MvfHF6XAfDWtORGWCUlnOyXELE
v07tCd41LHHNFtK23sjfwinX1wtL1p3MPjODG3Hh67ITv7RKJmewW8az1xN5X5MaYKoLS50IEvv+
CBT3LD3Y5g3r7iOiQigzmnZm7pBu99Qg8cvAU12QGoEW3ECQh2g2NwKz5UqgBC1v5i9ryaqIU1iw
9b2TpoBDk3r6eXHNhdfqWw+X0t9hpgnsRvHD0V09DxQphSdxHJKYT6D9EWRQ3BSqPcRD5+iX9kbJ
uinPvIQttOqjPn0dOihCE5HyGbydzf1ipkb1uDa3PIe2sptheT3fSkEf366Sc6dll8c3wIFSUCDG
K9SebvnRgxaSHVwA6Nc3+XJLMwroBY0z7yEkxWZLpnsjU/O7MTZMsgLRyCUsuBVLTmj8Egq2kJS4
UH/IFgiCzHOoto1bqbIu4Aejpfk+EQPpEBinFod1kJ0cUZMsA+H3whye2+DwU15Tc0/tvQNZPvAx
rWQreDDjadhBH2yhpuHPTvWmWyPOHLH6G9I7uYWH31a1JXSHu1nX6kU7sg51dgGMBsT8xN/xiRJQ
QkHJjS7kGeNufEnFDFXhpDxmmT0rOVn6T3lm+mxeaXWSr6sQDt6HlgIcPFO5lKfdGSmMXe4v6Cv0
6N89JmSgdUzu56BV32RQgYLIrQXhk63WtrbXmyONozjuitVgh2oGEWVKauJdrk5G/Ko90kVpw49D
UVxcK78P/a7FcJizMJP0obfOPI7U1FNwZSHI3DeQiqVddANOvLzkNkwZSOdwCUwvIsGT6SfF5efn
U2WiaGeCQoAUx1Hv+f8w0J9bNjw2CSsX5Rw+mBt0o7fpB2u1ZHow5Z1XmvbOpPWKJ0gJpxEZpoal
du7j5YZmSeiONq04mgsdvoez7rI10bQivRojGpWtzgd9/wfMOWKEGH7S5GM7BKHCOoEIiJuiL6Pu
xroj9uuV3fODxZ79HgjocWqXSSKSWHNUnkSCb1tI/3rrK46mMWKjZdE+UPuNTwPi3I/SEuovvbRE
aufWuiJX+Y9rB1Nwiqjml1vXKTdWWxp5e2A8ct5XBTftJ112rvQr5A6QR2B3QGlL0xhZxL2IBUiN
KLBiZ03wznQQ31DFvR+3Dis7EG4c2slSpamxms80erQToCmCztohAAg1UCkMyi+sjDeQt2I+cohe
XmQ+oktp+1Gpy5qD68Siy/kcZhZAAI1GCJLT9TTiive0MLLEbo/kzrLfuJhh43oW7ekKV0kePvbb
utdxy1Tr14lcQEFIUhYCEQLKUDvfxS80Vo9V/aRs8WtBvTzRiWAfHPcHUfi36o9T8u0I+0lABALD
rcaFnb/jhpqk4BYAw5d9qBtu+1DDyZo8GqoItPMLhgWPO7DJlVqz/xJOQTgqbKsZk2IgH3oD3I8N
+3s1lCr9NPQ+hrbt6AeSAvlaN/TSl8zdT2YCSBPx/NAi8wSa0hpvdcAFz8ISv9qtLjnMZkPmvqzk
76Gw13zdBmy+NthSxv4yVcMp7mHcDhklXkHU2n7tJ49Jsv3qettqgmPqygyKmg61+rrkFv93aO6u
QIofdT4lL/UXqUP9v9oW2eEeugZjb19HlmWFrGRf90fcn89cl0Vs3tekMd5hJQ474qmlcuA04iyY
Xms4afzys4RVIrK1rAm3BcPVh6xmX0AZVFPKFd33aea6oRDblcgPjm3txOtvNdSoZNBMNPERWUyI
EYzKxaIZjtjxm4juvUumf852d8PZxA/cjArQhB0yE+iQvpHpAL0r2BiWJYzprMl4u26Fsj3GFoms
8Iq2vxeO9j51tH613QJcWua8DPEH5CE7rU/sAtqcLq25xio46Hu6QEwhrOKP1drU5h/0UDnQftDx
HmmeFSvuOLB/kvG2qf96XcQ2JbKLPtaijsDHRaTEzEXyvMUThLq/QFvx27wGQThhHhHGoRij3q5X
FaaB9EB2X2TkTNmqHspHjLkVJINsEAzlyPRyJyBFjoS23HVQJtcWkXS3l2QArL8XAU4PH8Zwq1r3
R8vTTGe+gTXWEbYsMBjpbmRwzrg9595yPFhNrm5DdIAzt3DDMqKzOb58YaHUJQvTHrA6pKS+9kbq
sUd0ZkZseBDCICY93dCjyD3SzVr8XHcQEW2CJNqRCFxbTIx8jTX3yvDKQlzZauNe0WasN6XOZ5aY
32+gIG7E3a8kM1Anl5F3O6k/23ViSwtZ10xjWu0sjytfDlBzVpMnSnSBKO7blv11oDPnrW0Gijpg
Hu67iZQZ2Xg+39GEg3CWgPtbI5+LQul7z5NygZnthDfV+3d5EVopE39cQ8BEDEqMFm8czbb6eEDm
ofeqjUUltNudgM5g+oOs07tl+UBrscwLSf25yskaUhYrB7sDZTFH2xmHMBIx9OQurqVCBHxnp7ud
GighD2siYOK/YCtkddAvIO87e3DIgAOkG5qMZs2wOf1tUfvqZo/oQLizLGm2yrvOoeUfeXarXQa3
vvM8PuhPbXl6cHA6azw/5Nr3WnjSlmqJDk4x9m3f78f5ICtC+/c/bjq54TIJM09QvhgrNya0bnpp
KEMWU8M5kv1j0W+etsoRKBcAGatOu1hfib4lJVKiccBXBHBlfvfIbEceEhd5jWQuyNJCKPyOyvWj
dOsL+3dDJstY8gsHpa3sO+D/PeX1gTZKCoMr9cao36FuvdrZ+cQsDKgZ3m4uWi52ezbqIJfEjch9
wvmgrEoqhpuclI1385QkdWDEiPQaS7zvzmVvnHXeorcwi28qxrB31OgQhPaIFuMx0MTxDbalPGrs
tTchOJLDoYCTykWsfjMai945CK3zztcvoYfdvYl2cyR4sEloMsJjD+UAMHBtRzsLQH3eZ/cVqEvY
oGKZrA3wNIgGf3C4+XrsMRlCRmQIohhrUfZL1GmCw4nS6EDnF2DI7yzA/XYKLBFHoKUefTcUpQtK
6xHkuik7z+3k4Z1dY+cgbmkRftt3ZJjQXD2wuJcFuRb+KPmTo2BScfhZLvJPVnF3qxj0uhqlIL9p
bEom5MOsLynI9HmmtIzeFRrh0UhmuJJIDKhOXA27w1b5VZvlhCAYQ9JZuHAnpQHcmdggou2qdt1W
prOudRfDFd6ipqz/NL+7DW2iz6XflC6XKELgAoRCpfH5W31x3S78AqeiMusSf+wilGxN7otgc7Sn
GcFAWe7aGDxK2UO+BZZcY+myyGE8FP4PqR3Z5wNN3cQJ4eLUdhGzz1xbb8N5Oq6Vput5DmuNe8lB
T3/MK+AB5rwrPiuBA+89Pt0rd0ELfBBfOh/ErQ9ri5Zn6zdbq1H2ah3bWXq5vt2WkbrZOqWtHNGG
k8nE/2+HW16FeRHQQTc2zFM/LqeWQC3gMBLnWvXUY1RYK30TICPUBpR8OqDI6MIZJ4mwvUtQn5Ij
rLDEzB4Y3fjvAZ0gliGw39rwvpQNnnEf0KBRmrlDJ3F0aWzVS1c2WoZLuPnCKD4/smuaKPxJT0gG
FH/rw5OWz7bC9L5+eBV0j4s8Gt7HU8OoI/WqPv/Dg9HVEV9RFNmG63RhUB3LdewSZq1dSEqg8SFY
Ekk3c84cSt8VVTrlDyeuP0pPy/03cH7592vyquJKtpPhl9qfLwEKra5mBzVmtYlVm2AZsPD20rtB
I9/kTjCggs0MysY8p4mN3KH1VetKBsfR/vSPSknUq+uzZxgI4ZF/DYa175+qylQun44NBT98LCly
ftTCqBHnhohxE0j/VfAIGi+hknazIiNVA3NLMdnoK5i2HY5GHkg+ldV1f8EA8Vc/BI83H3u4INHW
yT+SigqLozpODozBKItyi21UVNo1GdGdLXPbNoSovWAquUxRSlbxwTKsYb4HATFwTZgctW7K+5i/
P3jUrFWOTho71n16NU4iu1EmA2XM/i3E4EyH7UJaA+Mypa58Sb5OmPnNHJ+YWBa/NMUhPpqUkzE3
sb5mR+3RJsbHSP4B3vlf3QiKKFduW1iMIVtf3JCD6zfe5FRTj25rDK4a1mEFvd7T5MpYhwz3cb6i
7fpaaN8dsaLIYZN3ZHHggn0vO5pWco5V/ktPsZvVrjYeos8fl49NSvi9XyZTpAgnqgqJ8Czo6GJW
Fa+3X74tRBy5u9KoxD4nQv2lJeA/PHQFJ9e4/ZgFKbDXbK48UNARhF3XWkyLkUkvlFR4YcTQ+GxZ
VIknuE+cV+0Mvu3te/ZDuDBJe+oHl7uKyOKKO4RzDJlsL6/Np09ZmxOru6CLplfy4QRt81Ktevey
TZjlG84/PWnSVXvjPdAP4sY0RjZVErYhsskValGTNOjqN9n/evFb/yU3Ksu8kssPNBCt/ezMALgv
3KLSFtwcVjt0zIc8sWwdV8TB8hK314GHN4nv4sYaPorlQz/+/ilJUj1AtIp6fE5Agb1brE8wLA2j
xoMj13YBFZ1qlhXJKZoAH4/axt5tvrmHJdqNwn4Kma4kXH6ReVCyL++JOPJeOnMxGB6Gz3i1gDXW
PmPLrX7u5jkUf8BLOjET9ITYkoYwqZwNse7NGEVRG2cOeREadz4cg5mEhPBDji/OLotUa/cTF8wN
ExihRagjyHRe1g/u9RycJTDDPcAs290OssHmBVXrI7ujZ0CemA2cEAsmEkCMoEpR5egcDXj3GL9F
qqfeRxNP7ztCZiOR2xsmMCyCGvr1jsMFWlX/sAgKXoLG7cYnzROVnCZ/Mcp+6R7Mzet+98HxshqH
8l0pojoxXyMRlpGfmZU0/1SThWP01LcrtZwwJ8d/OqLwmIJrLLWuJCC8A9ArlUdywG9fcGscBdaj
k5ZN5mb/NEz3egk7c5+HXH+iRvm1JvKX1A9G4xHf+h0hUqpZSKxhsckAY/5jBsNdx/E9W4ArZcTp
9BPM+UWV9FJNjbSmFpEbMZ30fP7QrceCyXBdZhZYTRTs380u670/e9006ucuLB4Qu+9dcENsWT8+
lHmFOotdtOJOMwBtP32l/u9xVrGgLlq0i+UmlCPDbsP7VbtGkZaF9xhaa1j/8+CoX3Ss24Oi2M9X
YDIcg9TVvYiSDdKtmxnrhj8/PJwfsqKPh4exh3Zye8+zcyoqkSsXPlq3wxHDrW6AcfJL3qfM5sGf
cr/5v3QfeY4oDBFjLDKIxldn3DpShbBzB2g0lrXlAHXwnmXsRShbHtOG/DvAHKUUgatVCGSm2ozB
iKQyatwl15I5g8qSxhy4WUIjQUer1NwDPkN1g4rGrvD4t7R15cGHBQzZWhlb6gB1AoTnxMfcmjq8
lAFNygADDQbCY0oPvRcPXbbcWDZMnnhO5MWE3cbU3SYD3pFCE3R8lnRwV1XuMZeZPxMkJTvMqhnh
rSdVk17JSvl8hjRFP0Df2W6PivLSWq1nXzTDKfH/Dxr5OiLEZZMMePtU99MOVAboBIqvM8hqjo/f
lKVqYfvfVuZAcbfNr0Lfmvzz3dDYAHHImcwlTg89g9gv8ESD8Pfw9Sj6d0X8aF2jma1ZTS8Q4y2U
E0DB9q4IGdckgdXPB1QYnX5N91W/gBP+53fkk0Jn7fpYMiLobSbVPaUyWNBjXP7IFvhO4FGEyEZU
q6AaE+NxbzFplgc/FgtuJ7AhDXk395nHiWdXhXk634LRIfxAfUmwbE/izTFxZNnSXFKblywiY1DH
1BIfByY/WzfzfKWZ1Cl1/cPtYPtRL1bU9a6oATJYo7GE7E6DSX1pIDw1MI1wAxeY0X9+E5yFbXBs
D0p8u+kUZJ274+MD4pZty9iaLtoLT39iz7ZtYK2H0p2Ao9Rr/fZeuMJNTFd5UvRk2RgG7CcodKpQ
up3YZf3MOu3ob6T3byV8Bqa3XCJatXMk6OWYadlBtgr9RGN7aIEM3iVRTzIJBzLzszax+RgUBSAm
77Tu6eYEdJAYEPIzy66ZXEcIRoZYno4qaioIXA4SfhyPb6k4urbPpsHSGzh43fQF+8GZfaposmBl
BTavRyotRLR3jTkrDZ9I9jr3Xw7FG3I45Hk7uBLiwFF6LXdBKi9NGn+LFGcMP2Bui7BSzPhhvNFc
okkmc1+E7tMr4+00N+ulK94WBm2fCTXlxdcaOtBws7C+mbvoK9x8PFi7LmgDH4o1kQUE+AQpZSJs
dBxI5HLoOBthh0dXT0AFQDM52KJwT7pv+i9oHb5ELKLAQ94za1vOUZ4hOlx6+bj4VM1hK9chsDqO
pW0vpFxpJ/ImLh5lzJJV6tCB1QkCtL8O3Gw2XP+zI6hJ4u66ijYqIVisHZHr5wV1l85SGfLWM/9c
bbNNWo6RKoEfoiBPqZtXEcWdsm11KOrmrI2joQDx8feU3xYwq4LypD2xRL3ukP43NBr3K8OWyUNv
mfkH+zyyTdkTx0sRCHm+rMk8jTluurOpA1jgjzFQZVw0xSSVXuhRMQt0sdZpjY2mZonKT0LUuqGC
SKUUIX4qsM5NTX5vAbIzMYLLhNV1EArFA14/ERLyZrtMf0GTLdfAbPjVttRZFZWKe6HOMLmg8zA1
IOituO84QLkYk9OoXghJ21mgntcyttr5jUkq5/qHfRdTUg91ZXlY1VKhuqKn0ekcDvMAsCUEW8af
r46Vq1Cjt/70GJq3Ia8kZuajSz+WlbWyDO/3Xm7x3R82HY2IYrIw9ADSwFg+xHdl1BkIZSI4XJui
tpFcrlCR34JAn0jLIOkbAfbqB0v5/rGqNDduwDDcCc33mPdbvXisXfjHIR6JdfNWzFIymIlMagVs
tSXr32avoLCCpWbkPD2UAv+/8trHj7exgaKmnVAfYbpP+QfSmRYhhIctrd0bCv5dpIFkfyk2+7dX
BOPU5yVbpIUIrFKXlQyaUQUOvI43uRoaVlpXhRwjIAmCnvvaj36b1H41xZXAuxJcS6kQAGh3oHNI
PaOWLCS4QFgPr7o7pb5I3IPcOkXC7jcBFejvaKT8dfgpusRrkjlxkDajQrei7fNG2Z3BFO9ROcvG
P3b80jwFnACw2wTbI15iKpWyhTdgaLiTpJbLvBUNcMWxVgnqwvs6qYKDqwmLNuYN+OPvfi05sx+h
pTExvszI8HuKlZGN1eH2ZlOZjvgBJ2gtUKlh6Th1nJCBzOQ8Qb/uzLlLdUiMVopNK87MdVGLc/5E
96ICYSHFwA8mATLT6hIp8UNQwuR7gl7jNVhTZKsbb0e6bOseS3XaIw+IWiXye742SIRR6IAx2D8E
IwKduLNbkaQURao/Ii4BhIqzGmu1DX2GLISZllXpRe4KLaKZEhr6o+4GmNqNZir9RkoI+1GnvTYF
ZY2gq/vEhCbRCn6haoVbGMLNb5c6edfrthyXsR1Sz1SBtz4ByxQKUXlofzKPYCoOovl1Je11YAkt
xoZLblCpF9lviQRJAY1nCPtuaRbrKm0J4M99Ye0Dy9cS/z18lFqmKyGQFIbRxdUNtODxngTimvjy
HtMVnypejWjflMFYCG+ATGazi4R8UP8SCK2pOKs4AK9xhzBc4qoTcTSAySlUXToWRQDFMIB6ekuL
vwSU4lua/av9/0xZvMKYlx3tyv2qxSPJk13egAPAmFeI3I2T77JtqmC98y/0U4E6yqgNYOU207FE
0VGUHMTZ+APFi5YHYqjuxJXsGMayQt/pDpc1mQNrBJcltC6LABrKXSYhcxdAnGICmG/l8TpsEhVV
ftAwy1GlG4D694/n1ng8tlbsS/nEU+XNo2eQIu4V6k9sNLmCjbDOzLB4Ay3OvBrTJuUUmPkWMaL8
cFIBoq5cM4hmZ841+wUfaS2E+q1ITBgWXCQJwdaK0LOXZBklH31Zd3ixHaybj+98GvjYFcqBirAI
9K7lqrnSka7KHlvNFe/CjDW8DrZ3sW5VgNJ8/oGpYxzeo/NGtLr0EAFg5CFc7G12u+r90GQq+JEk
2fNFSzBylZG54W1e6l4oEhoDvU8X9a1vZqhOL9xXBD6lAZX+ejfLg664FCBKWJsGhE7cwVhR0np8
WhrNjouUUZYslmnMupXYwK3ESCz/06Uv6V6Ymnv8ubXYIrsTrf2zdCmre9FLd1UnWdKaNdOF8AlJ
lGbBoAhFKoJ4lQxAm7Ivv3/jaf4+4GTJHQUT/wPUIkb57lBZ6bpN9t0LqaOH+DIzfZ1+Nygf268O
uQ868OSvtZleBkWjY1l0iNAGDsEGWJaHSw/W5M6Rrqhk8n4DNxzmvlMlKDmetSkv/xzC2MFbbzYA
YERxIH3MEK6E+CKoxOzwQ36KBCUvPT2pa4nWoAzi3tfzGfEVBdbvziY+Dcim08/dyI7H337w6Fs5
UV2+5eqiBzQxYBiwKjSmnP++Qxd+VMHALQReEAw3EldrsSLo4kfYl2PnFQUNCzMCoLmJaGbtNDKt
4j204Ip/HFMPmvyITApNQPUcCjQ0mEdqCahZMNAB+nP16gUPHT1vY4SEZwAkAQJ8pkcWnk2a750y
QvHEUY+ByV4TcAKD4BEoBA9nA76DqNHFRPhuZ/cjm/xvMjOSHMrayO3fGoi2w48MQuPefrDZXDpV
0WHVWwfX5iWCHvYz53Getk6EhoCQZavZRQUG6SYcuo7iQtswOqsi2Gpz9ApyWO7zwUra/NP5qsmF
3rhGFTDhRooxoI6hJ05bssS4ACWVi7Stoj+50vqC+Dth6PwX5Zvy9Wyn41IwKQzRNCCuP+MKIji3
HI4Oi8s4JzWK+mD3YFmpANPwlURO61nDecyBqhtcYt45RDw4QoJG/MCyu8ZrL1BYFj6MDvw9ODZL
LMn5mZ4BRxmxz1TWUQ/HaXXKzseWqoCuwCaibIFal+IEVKEXYnEl/Z0qdBmGpfSf426Q8lu7sMp6
wDLFN7/thPAOFjqTtoZAJnxj3C9uobf9ryWhluJokfYmwU9dcccV0/QVGcLSnaW1WvHIL56g1xAi
EOwiULcVXTEUhJo0ZwmrCaFNEsWql5EZwqeYcGGX0F/yn8xCK+Jcof/pHqTz6KB1B8Z4FdXV74vi
ok83gpAFPuYs44FpniYMYBRRTAWUpcY18AeQ5ab33vuugNRWC2JSN+3PR8q0hMUKnuNNStpDH1rB
WYUCTu4YQNx5wP5Phu/ZvASyQXXBaLWE4pzMue4eLUKKeSfyAAGwL1b5YwqdEyW4iZ99KuMccmYN
DM8cGxlcMvpbGcmuzftyjWBdslFT9GYCV4ssozeacAPn6qd2SeGMNprX7wd9TJK4JXYZyhCEjdAQ
6+8rBjD5CjZA8ywxs73CwFaOiGv2ALj9bF2buJsst56ONH7t8MsRhDsJgR0vIUWN0Fn0qgMHQl+i
rtthSL83jS/drsTwWQhIPQ5Ca4HKf1BxOzYqY97zCN/XIVy1fM9OXEDPp0xx9GGX9qz/LLUsYv5A
jbvlBp3l/jaHeiXyCR4VFZM0CfuhPyZmZmXAzXK8bjfNuOCFEjjeJLurqAIOQNbTvz1ODj4cgF1k
YlTqeuBelsTVldU1bm4wqpDz0ve6AXSQQ97ZuI2nvRkxHkwEnx+gJ6KZnu+lkj7hd34AvW9Z2zSs
Wr7uAGMCGWLJt8U13Ag8AGQS3mhFAVWV3gmajpbHihWJtzEImFzEzwGOymJGrggOflKxMpqqCXDQ
kjix6b7e9XVfiFBGRCF0d6GBN8M+OHGOuxF1fLD9y6G83BF7DHbl8rbT45IDfPY9ZZ+r704nQhan
6WX/gAFfIZP+Q+ZW7Oqh17B3602vDy4hX03upuNNGBnOvSnD6j68ZxtctACzajUN4CHHbjrgLmel
5qis9zm2N0uxJGJ/2YWENrqPSOiyZt++Z4Ol2whPo2HiWWJDncfSMZhZix8VfdVyAlETctX1M9fe
J7UB3cFSUdDWact39Tae7AAIGEhIQ+ZqvAY2oygx9+kyEAeHpBUSWsxMTxzNCHss9jhLS1Xc+g3q
TBPmxRZAMlykKeNGTz4Ts78cdWWnDX875HMaqdHiomeEipJ/LgeG55N2FstoX4NSysSw7UW3B+Sl
DvNzSvi/5aWLr9eESNs13KixrCetgo1OVT/n1g+Kl2LWHCpaBrLufjgTUFkJHNioEjSRlXrViU4+
Y3LW+odtNxouzvVddNL0m3bgwv/QOpErpqFcSVhlYbDA5l8IgeJrha0EVWzk1uYttvCVgm2A24DH
B4TLo6WwTL4+gJCbo50hwVH/0q0NT9spZKlMtYOjZ6vMbuEpQBg+bjyhFJBIp72fmpGo507Ie6F0
kxcmIMRr+5kGb6bCPv646a6fkfuok9nlHQItn/ZUx64Naqn18n7SoF37TECnYPNQQBwNT56nH0Wb
qRwgJC10cpsMyxzmPU+WR2XZvNZKHJasjVfs3p12p7Q92zhJa/yuC5VKPIVxZbA1pNUhmJoinK69
cBCZnwpuMlA92fVdVChPuFvGoUAOtStOOdZtkqEsyHnf180+AhJIfP/IHL0KGevS66Pr2Ywebvu5
M6reugSIR8satCVwfjnE9uDZRlQ4iH+i0HmcZOdfs4XZdf+IVY3tRo53n21898Q6ivxVfEVwCw3I
lYPkTzpN/MPH9vuBeihWGpj61B/ItI7OZzWur4FyU5ImwEKVEoct9I6rdTUBGx82S+BiB/FyubV2
lJhmam4jO4c/8J/rhry6V4GkT1vNF4Ooud43XAmxLnBzbQt3JMZ9OGHk+ss8LttmwQQPr9j/t9J6
su81S5vEEAs0im0JhTJ3OHTL/ukoMYZf0FJWDQaJRM+5/1Q8QucfGf3lJJsAhEXZHf8/zh7nGsv1
ALB2/VL/1RdiDiaVHmnjCknwrkODGSHRMKazqSZzFSN3oLSHr3kFCDDb1JNtz03ksIyiG8CGOK3V
m+1QyQecOpTW8ovNq4WDqei6E8rNi7JTpy3LQ2dvAxhWOI8n1yYPSIc3WTtSwJkZBCSN7dlqBWBP
KPUo1jFsdTSQByZLLe2y8mpi4mqLsaA2GS5WrQXXXqKY8tpIllRpnwZb0IFaPqnSFKYUoiteqRkW
Xdz8ixbEi6uxdwA3RHkbkPCwyBET1tBPQVKD9R9yO8kBlUW6WU4VX6IOIXL/B+UgA0J5hCSNiIih
uoHceJJs9YULVBEiMSxK+nWtgbxZ79Kdro01GVP8fX9LdT6F1TuJ4Lj3WUVMGyvnAhUCG1t0Kfb3
jCmt4w4mo66SUSAnyTZUhKTeIp8e/q6SO7Nc3UQOWfgkimeN3KysZeZgoF1/uPdpeIMgx0dND2w6
YhGbeDsHyUecF16vq/rXq/xp2js+1TdvRgPxos30tRDdSKPLp+fuW6sxAE4R+8+dvOu5aVdPZ499
rnQt3RHvdj3FbTH6yj4ha/UZjck2TbAv5pi0E7Wb4I2FGUWBbscAa4DGTX2yu3djp2Rvr1Ay9hyw
qs44qliYz65YnJd1WnAHBy6RHmY/euH4jmOGVxEVoy2ubry3eYT2EpKQN265O76cRiIQfNRPo8v1
nDtlnTqOilPNYMX4PdbUEc36TKhofgVFu4Ho60yF5B/9qGWjVFa2HJ4yBzyK85Cs9B2vNR2dFUWT
m7wEXk+Rk68W/69b3Pjhtrt8RxOonhtTHxSDGqGiYNBE40ulg++OfHMJsqk1nDKiS9J6PrVFcL6L
nif9R61639uxQkcc54Vyl+fuADRDHwCbrO+w1oTI4MNU6+Pa7DSZlw6RroTf88kNb+neRFuj1TO/
tH09ixO73NyGvPJbL/f6TKMRQuHjhCoELeXjiX2az6GFTM9ZaleevqWbOjpCGXNgodSUGjfoRvqU
vIjRzDS7k3ukHNY5ugPY2nvHbJ6BCCQx3D8fHTSPz/dOPN+qJHpe6QnJZ7u09/lPX81oZQj6i/9S
SpfuObmoFP5RtkG7zUvKxMkLy6tr9VR8EI9g474VisfsuJ3y5AWh5RhmsCKDXgkh3MUpTyZo9rr3
XtRncqUJvusKbpzpaDZrXZ0GD4Pu4SlvlFe55L2erxB7C8SJGGVLhck6de/u4PKrf7/Mzlr3nofL
51bZUnbIKoenfsmDDPp/3NJF/7Nkb8dpVrpGt21efYHe08WEVjeh7p2cB8QdM1WdLl06tZU+wRtW
9T8zi0nLaFOb0vMsJdQsn5Eq+i7LhJXM5JEhbKbbSpaovq+5c09qdKzR4R5zSOfzo3vWvwhi4J1l
qCV6tEbBGz9X844s4cZQR+v7QBukY8vqIeBs4yamKR+zYj1+U7B/BlKZ1jb5i6o2QQtCC6yk5oMg
RzVJ5d4xGo7XZdq0llLF6+JxlY6GB+zFJh5+bJY+bmhcNpAItUZ+f0lvFClC4emhHmLlQ99Pkabb
JvbTXwxbD16f+FJzw98GtRNbGCLU+Ue2LuH0xAEhzuAq4JwZrpXsXFMqSNjpVH0+StJwImsqxDL6
nPsvUA7FEm+oikZtYuXOgh4JMiwzYvgBMGtBSsHzODqum4Q6JUJillG+n6lo46L/4cJcoK9pLyeT
caLv0n2GU54Aykd53BBcf0lUjhHYzViKtZa8FgoILCPZXUgTkShuyBSqRXp3VQcDHBkpI2MkpB1K
sWdQTRwhyQDHLZ1LN4wrNIB0Gvm9AUk/t+uzm+Az4dDysFCfQBiaDKBzwCvHe2726zWndOhX8onI
pczcbJv1SoSL6AfTAV6+QaYmiIspekzXqiond5PmrruJ3laYtnXMnGNgC1Bl/eAG/tPXcJgGgwXA
knaeNFcrvrdIWl8LxrLWi2H+CiM4v4x1LHd4/wRv1JX6Qf9VQTIaoxn6Cl4TBKoGym4nE9uMNjIG
daBDsFvtRoDQ6NjFjfzbkRXbriCi7AgORszDWIzXf+yiEGxP9UVfyHmM62uEndsmUiQf+UH2Em/8
2qrYtWI7+wRQp9wLplGUHtLwp69ZGLazgTlV8FYDlbYkGkcGMWl2jgtMwZvHs3zMXiITbOEjeTer
faLWK18/pTlXDsDZlce7dxYBwG/9bv4ePl5raFtYFwB4XK7ocPWYTYZRYSy0+PD6QC1+ys+kS9rA
I09kK0gLkYWIa20fuTZBA60ZKxNb1bLEApq9+TGNEdK7BoZiIOYoX2gE7/Wu+GzncU/l/lchEaJu
I55Hu5clpxl854D+wRw1uKq04H6e+up4E87SkxqNFISDKJhfBX/4EVAENjC15yAEpGuC25w/CXV3
xkmL/Blh7b8ZZFgC83+el2W32obIMw/zE3uueweq4NVAOlgwxMcOLovlD0DvXOCePx+yLQZkT9aS
sIKhhZCuQ6pt7mgVlAAQa3hkoTEMZiPag5UtnFbdPFJNBWGqvqwuk7+4QyCJ1nrBU0sOHRpQ9An4
WHpgr3/O339Vx3WrDOMhmt55Y0CJq2xeG30uuVbh5NEU8cEs81MHRW2aKfTLNeOrDGmSwXtM4Fbt
WraFzRYStMXi9SrUHyO9x/XGwamtvKFza0LqEmwbciBaqvZQAGUGfR/u8WJhpla0CyJI9/bGXazV
w5Oi15gNNyP1oECHuDmmLwsq2HMbSXfxIsivcS0aE1V/cVOuabgsEXYZw0aVVuZS1vKZwczV7mbf
h3ddLzvttmZzygX6MiZ3JmzRRGlvFZEMWqq1MouqUOgYmhOukIA0Weazy2NTDnfMg6tqeSA9Wl15
t4zYDr3XEW8MVekykcfz7l9JvUFJ6eunzSOrjvCjbUBtytnj8vZIdupod2DrXOvealOBluW+MsNN
yqctvY5FYF/5MrTDqdPM4wYPQ4/utD86eE2/JEunpzHYnnPSt9UFlXrdY6jtzmJUP3dkLZgAhJ6k
Ebnt+7Mr45ZyOCHLcJ4CPVJF5HKoa3deLs+ujRr0r66kA/JtyfUq6CuWpaHMiv4tv0By7H2Otm9C
IJB32V/nAjC37CAuFcI42FDfQwza15SqpGJueXouynuO9GfjUCPoPFaTAmhZ2wYqEkZ/v15FQD/q
kZuCPGoA82W4r3FSOfz9h63rHSXEeRu/VK8P72wqCHygt6BvrUgU9Xji6RgVPygoXyiHXRRrzPjY
yNBeIgWA3pZdhxrDs9R0VNh/z6JxR/l3l8OGqezeWfqcZSvWcq6Z9n2cTCJWtcVaTeLy72HjkuOL
8YxT/dc2cg87E2M5tPIAuCBDxds8jpqoC1IU9YwJmTXPH9YiJQLNmoyaONQv/vDY8+YpfvYly6MZ
aOOeiQglaixKjQooOlB6wBNxVqr+U8VYgj97anVnXR40a3dKoLtWKLDUiM5OUrLLq1IYuKPbyptP
cNLxuXRVP1zC1AmQREyt1Y44aXc+S9Pbif2412f/FmYHeTnaYB8LoB0yDoMUh4OUQWWDWdWgx53i
HgSlFfPtpclk2lI11FI1xGetD55fLCBBRuLi0DPLWFdOFijbGg4X6f3nMB+4GaaAwyQOMh/lsnD+
H4aBx9Mna8pOhcXWWx1CX6lys2vHqVcY+EyG0nSJUarjCl0tSBAvDF8ypbqpXmsDmYt+
`pragma protect end_protected
