// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dykjrOsd3CCYLdSIlekquKGZmF/CyyZbuaj2dZlBC/pK0c7swMh3OfaMTBWJ
IfXBrZ8u0IPGTdFNLfbXU7SHOPUxnJ29WR7wtHjNFn1yE8OZeB0altL9drhk
Bu48bnrpQA7PG+awghNwDub+k17JGtbAvwuu9Oyj3fz1dz/xvH7WCqvSAGry
q4FUdFHRDIB/9pSvc6L3Rll2rg6F6vlvbLgAEgxoy5lNPGbfXV5Ko6bdStIG
cD10SVEZPNRO87HPF61STzG9SFC8Yc1MUfb9ww0r8qyxQ0xnRQKDoq4rjp9j
uw5Bl6SQjx0li6eSlVBzeJPF4dGdsbMyR6sxNKXGEQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hTSOA4zXwoprpAEFilW0BtPQ4Xoc+XK8pG8dOMuQNPoEiIVDySRr0SSp04nM
CwFt5TDPu/Qvho3nPM4+8fOy7KBHAAWP7qSCF7nhlE7tpRgP8RLkkRWLs4MF
ohH+7GqS5bRwjquHYydTKWiEt0yZUEVcCUf92IhTVMosBMur2JRqUjcMaOQ4
hwQf+ki7AYuUAFp8jcTQxYcA/8FLmkmxy1se+3UfFNnLYzhD9IJLnVawXjZB
aaOPYb2vLgVtQG35uueeYbCV1wtPlDUx7Kzox+YZ+w97nug22cYZwonuNSHF
S4nHflOpPl2cEnT0IWnP9Ll2apBvIQFc9iiAuxlCEg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bEcBv0Tlowy56isDCGw5hipzuP3w7HozioT9g2mN/8/HUqqCNGuEjAAhZXwJ
YKn1l5KunvbQs/Ayj5UMLV9Ig+E7jqLDt7rj7AgosgU+I4hnXJCJLIj1/2iZ
epwN2vafbgaHUYfzqg3UFuHvpNX8Xn05f2ueNxyhaAtab/A4TKezJGyaALag
g4SKDcOAUSnB03QCiHDZ6eTFRoyUmHlGXPdEw2b16vS5hGofcPxatNCc1XPb
jMglSNSncWJR3U4X9OUvaFAFF7wooiNwcqFh2LNQQnersk5hGHA2CR+la87L
hipHe1P+D/Bhd4IASamZ2IeUq1aLwyKt5mCOUNw84Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OOtrATtzXpgYWYM0puc9cAIhAvFRwka3os5fyOmPy5fcc4W0R+BiNGMh85fQ
XX9d+bDfv5wzKw3hJYgH/eJ4tu7OiSXwmN78Xqmml3ybGZHwSj9MfMWN5/3D
mgCEZDJI6MMMyWBKBoVVj3YsJR6roTf4vpE8w5pRavA7+JPk1YA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LixPeSWRz7tHX//noykwkE5ot+eCNz87D0vohR+nP+xNzJtj4fFmH5ZAwc3L
GnSZRmFPq9gDfGbNaUFpcyBwuy1vPJoUAeDz2wsI1gyQyOUYd29IrKGrsrYg
1Ah+jm2+jaKx/YFOfopRGtOY6T14YKahjSaLacT035SenpmHtQeJqLO/sYBy
AyRVI7BKmMShkTKJaj9cQnTC51oN/lc7/WPGiDJB2ki0ruOJ/UUt0qX0Ui8p
Hk9yxAGM0y36KYmiwAWmLitZAiB0gfs3E/hCu+b8iKtGm1OOK7Ub0MlQBxut
mPNg9ommZlhjTuXvZ2jeQXyt219Ixwy5WTbhrQmNXl76NEtGsFsXNTojynPq
cyp7pAP9M64S+EV7UMsYF9y1+ARwy1UaqfXImBe83xE6jp+hLMA6UtCEqWxM
KZulNdus/MKGRPcL17p6+enHaOAI2p+SKvfXQYr5u+fxxWTWBaEDBwEanfva
5s232vvfHkcm+0mP9YpAcMcXmimSoTE3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NZFMJ87spYeDHxazhCSAGRXZQCsGTwUXg99lKC5VOQGYz7QlMSVDMBw8LC5Y
lbHkrXw94JfzonWZ9UFcLpOxMTxOVFS/syNLf7Tg6JOfQr0oYCrozFKBBqU6
AqC/PTpNUDmYkbi592e5VuYqso4qs3by2ul3xBpur1YMtjKLBzw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jUaqLx75T0O3J/SRvlFKAqvGc8g9qC5YxHszCCohOh+yYlEYMhOONe3lBIML
qPyZn9O+/cYu1wmi6aAMfdEQZGgokY5zDvJb5L1BN7pOohiSjk7qahxRCH8h
UfJxITu8LdbKwHL09nmd6OGdCkMAbTM7tNoS7tmlhIynmyC7BHU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1984)
`pragma protect data_block
iTaO/amfHL9d6hMUpfoqaIA2ZySPMh49V/drm2k9bzZf2MatbhYvUaBQEd+9
iK5LEkpjXExbxCyzXCVDHDCyA5uc/nt1Wnr/A5WhLrTSTdJIUBH7gGT74kfj
e8F/4NcpqPHvIW+wlMEYOUUfDC5Gi8/0T5Xvl+gny7MtO6UHf1UnFmDa5n8l
6ryVdBpFpIK7Wc0nHGBj+WEhx2tvoDYNKZFduIrCdvWHBf1mgT4FSHCqUJ7B
ZhUVsYqeg4Oy/mkNr9fWhJZ1kamZLHNRW6IYJuXQUa1NNHiYOiTkAcIOutL+
hH2cDpIxqogk4W85Yw5nDpyO2G72zkBCYulMagfA0vP9eOguDjXlQ/qClWlD
lV5CMb2XvlSwEaMkkFo47xMjIv51fbxUG+FcmnuLOoVnxbLsiXnpAEbnJJ3t
CSzuG9nLAk18cn7GxOayIb7YOsckn28rK5ztCb3sUfnaHccJDNvBgOlSiELZ
2rP4SGFqqD9zdQKshEmg27Z2hpzpwDvvg+40c5FF0T2wlGh4yO7I73TmUps2
kiMvMriQcO3PDkmxlEDWD8AGBpISRAqqbI1MguxjQFYEUVK46B+nKU+daxh1
kY7dKkVV2sq1iz2mQY9dgvM9vOaO7JRglzEECnqYcH+KQmMjLmsaJwIKQp3L
JfnY1wRNi442w8GLJgfkLaC9xvT+f2rO2RJMNz12sf8kpBboQu4vLe7Dp3bd
sRK3909IwV8+yRBJ0qWq0pgfM8hC4Nubrrde+7hRQ399//VmiWBA7z0634Sx
LTZpvrOlQzbpXYa01BkKtN+nIK18yXsWcNPofbV9EOmYxckxH43AVmokMD6d
jVDfyqPHPY9z/KBdctDKr3WdOZQGA5FktFFhZW8hvBGguIlpym7/2YMrVEyJ
/AqgZzpP2DqMWMtGmLZqwJ3qE/ghjv+ADOLgSIT8pJLi+34n6qthgJvfNoOi
bJLItCEQgIJDjBQS4IpTNQMTOqCxV+gCiB2I06yHMN0Q5wWNcu6i2OE4JQHC
u52JnLbV2nrG9yeej4yuLZDYC7cja71e54pj142hpSgpOsr1yTNHtrIWHs7I
oJGN5wpHNjX178X19dQrfZXrscGmTkg0T+gLxw/Yzh1crDs8SDsudIPAZR9B
PPBxYMFdMvlSJbqEQmXajWUtLSv+OmBO42YjtrEsA4+ZcZoTMFHDAhL5ZY3K
d8FkKBVCCCiUUx7a4GuFi9NQAL7nrAIbU2f3JIxm4Y6Zx3ZLEqhdmPEZNEX7
yF1a+DiHmccf0AuSfhvGUjcx8k04tIEfl4j4O3xeR4sw3KXYJzJkNb2RrpNJ
AjVEq4t8HTpbo2A2DbCEl7xOOjsR5FVuGb7Xr67WAD7orHldsguHAobsjiBC
FX1FRm5hFv5Cb78AWNlEyndrNH/EzH1Ock6Uo6Cu1FrIAevrFHGf0sXoN1Na
9o/nPhRrx7cVMxWVtFwbS23NNFkbVnC65KOgjdl+MoPpJpmRxUssVGaFpG5s
4dj5h7ii6DpK4NEmIGG/ydkpjVkgShH72D4Pn9Pz/7A1fla7bo+m2aIZuFrA
djk/9qDRkDA34uKb2fc41HW9qJCDMSJrFf17fb3OFdbVhWg3iP+gCs7KABw/
Ng0BZnMIUCim9zcTNnjmpDjU73lDbLAZItlk+hyBoB5N5zT/uSlQ/JrMsIG1
s9SbjVyJjhefQCNljWtVlOar7znPHA4v3W7RDxAJWtLW/4FTFeAhjmXShlit
WXFEGSJtqO1Cyps/yeUAImZnYG9vwkMSCkkESVSK9FjWVuDKhAQLLjwOR253
geCDr1YirHBnqSD+aMfgsq/zInu9EqxM5082OMaJWKFwmXPeXLPKaXXQL1vD
nQ02v7RFiA7mpSDleU2wpLYxNkX7dmdimHMFI0D07MSGUYCV8ei8/TDXqXWM
QuaEfFXaHxDerUuex/tDw8ZMUWZ2EKfVwWA3cv5S1Yk+/Ypn/y2qvi0tD6S4
C9588/+QzAmSPyQ/BCikrIQcB/usvmpwOCoGXjhDyiCeevBrEuUl7qqOTG5W
zl5o/UjN+l6+osrLowmuy3/08GQwlY+2nI6GXkiFVj4gZghDg8CwS41boHmi
KedMiInRryVPxgL/H4PijmRclIecLxuNA0RzIQ8lcLsPKpcIzm1+MvFcA6sZ
CEQeCRr505x7kROMjOICU4202WwcvlcmyRdpF5Rsl9vCUGw4IHXYL/YC6uC+
4130maL9Ri1i76wfad6qgkL3k2lmd6A1eetx+9eVFrgTwfGClpfmhciHUUQo
P5qJ0x61J5RKz0Me3NBSVVpMDMfAKDAD+Fs+Nc14lpOoWHnQo7S6tpgwYJUb
W+AwX/pKEpGjQuSVAUi3m2v4S+3/ow4EvBhZCF0V8aCa71G26ctUBJQ4x63j
wl86pGeIeJ5Z/vQFjJq/zTfVU7/zguSCMAh7n8+NZBDrrIqxI6zu0xv0ZnWi
hf+vLnEcniq4QilgDwos0198cR+mmZ9QySC9TVW36a4DSJiISalQLuyklNfe
RAzZhjAe/6xN5Y5W3Mp8nVUzBIzieGzNkvMKA8Z4TTFWEaK/YuJzaVKPomRh
39rS07cIYC51ZXi07qQuxzX/mazbrBqHyxbBk0QSafmNOn8QlSRboy6pIR5W
mOt01g==

`pragma protect end_protected
