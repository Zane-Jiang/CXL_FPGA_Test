// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
II85kubGxyqJC5odVNMfVCgdOD5XBwJjUaKM9CfOnQiCOQ9teg5g0US5l8yc
UC/+v7W/rHOTDmDuzEdW6mgllpW5FmN3AK3PjEh6reIG2yZKrMwbJqkMaNeP
5FNhpjBxJhAxPGuSki0NTvVCXkZyNUUzpUW0+pepBFCGyacuWI7GOJxyCCYF
ddt440OGIhXyGMJZksi1xwKY7MEjIagNPtoacayOFFEwpsNIBekPORR+S6lW
NofpyaPJccyhqOVs7AikHRCmIcYkotvol/aZlT9C+D82bElSrgKSRNP0sN/D
LSd5dMtBuMyw6wNUm0bD1ZGKr1FpiOTR43SQlZflpA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pINKHIa/gZfYCGhe+WfrbZST7ABL1ZbWQrLvvJoDagjYN6Nn8y/qhA4laCPr
qLXedxzhLd6DAz5n29IY37jTty83gle+ukyCMHqmM58e32RqaHs6CTfe7oiC
PcNncJuV1hKq9Pvr8PMAoBpnCwamGgGGzEQAiNlfPdATHVxKJq7iERrhj59/
5vkXr4Lbo9YZZu58CeuOtVwVie9fS3wAp/+crWSbxmReRV5S3FVYqamxUgjb
dDxNQT9MbSrfNOLiP9kOj07H7/Y+YLJ0gbFUytkNVByOgn9MBq7ddtaFB0Ee
6NtPBEZm6uiWm1DcHcYFMItcPSjnVWmWzBC8ZxF5qA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CTjlnvv+q0TsI9xIcF7Xq88QnR99q98IVL16Z9Fc4n6Tav04DzXRXT3T1at5
G1aMSrgSOjUv6ERLkKG03KxdKbF/taD9JHAWTDWXCKySyb4ljl1URYxjE9gJ
XPaHn+J9tNtctKp99XgpdCKBPYQXe5up4z0VSrG8a9qLcZZ6688gNvvAwjo4
6F51NhMotYenvq9By0W+6hFLRYSOOx5YBYZJFpzArAL4/oAhC66BzKFKuTxt
eLtsIFVGOT2zsT3oqouvREKkDx4Yg+HMq+L/7IZ6LWHRk1g8Z2SbPl7LuHAj
WI4qT0Xx6me0yN+deW5dubWvHuaeaYNgH2U5sYO8lw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PfHqYv8oCHdkwFZXOd90/bL4Z7jRthApw5UbztuPsM2TeVIr7ddJV73393PG
36dzaIRr+I4lsdzx0nar4XWtKJzylshnoMqQnJXAuKdS6ps2zisug/mkH+3k
PefAqPbXtGWXpX9dwquyFkcL5hZobBaCUf9tJcug3ziH7raB7XI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
acP5bd5wySqeAtIOeWpNgHqMLpNd/+SFD8IChHY1Uq8sYnHSRtkjLBneWMu8
A6qfaJOz06Oo9qXwYgg599v821yvzkGEdm5o390s2d+Rgv1dDakPlx53qvFV
aTRxUy/rC+CzHM8AkWwL6YMh5JuaoTZX0XQpuvWeBftgse/UJc8tP34+o7Iz
r5+G/i5cJnykvHtG8GrG+ADdC0vXm0jnQB6cWa6aLOsIYqHZY/KPGYFHZDs7
NNHhC4b+YM+Ga5BKWH1U7zdaZP/VVvP4TfhEB8pRRTvsxnBzfJDbuk1DuXn8
D1WRDhjbHzKH16ocA8LFkZQHMkWtVXShcHzn2nMTH4A5JAcR3qxNYfBjUdNm
q+iC8s/0e4L3mcBnCzHj2tcGFSluPtlYCcoAEjY6pjcPm0B9VidzzAbCiHxP
pKCvolcA2s+9iQXHX+EFSL8CkeCCvClQ0PdXXpCtHwUXvz2p1QGXt+4VBDm1
l+ujPzP+koFzpPaoI1+DcyDzgnvx8Nhi


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FyuQZPMmAheP+OuBG5rRFditLEY8OG6fpbB97NyIyjZC+BLBtmiCCuEIKw4g
HBHoI1TL6GgOU3ehipe0VX2pDc5mWTjf8nwZKtKOyesEKTFlaU3Fvbm2Fv1y
1QRLdtXKhgnxeyoKS4JjlreLd5iamBTr5dR/Z69Kli2sjpZK9+g=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D85a35AH/DfoQnYywvi2Ko0F1y7GLLckjeWZVSNIdQilcde2mr7JgUMBJ3sl
GXCj6rAb2Pl1JBxtvnN6pxXvifkJBMW9T7vHDOcBZek9nX0NvfOf6H6zT5P6
Q/GctsSz066632jwIvP0zuPaqBgsfw6TLUzwRdXQQPud3yxU5Cs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 329984)
`pragma protect data_block
068ro+7YuU/8PsQiJuPs8ARAzR93EuyA4Vo9xwKGbVnQmY4d25bwX8ykaXWx
FahMH5PKNWICP3cMmwD4DODCGMNl8uj2QM45koxDrvweXC6BBTSLYNSg5/wG
KcmdehlkzZjc7O4c622HiyHBlNRknbdMhU746EnzrsWZM+eSTDg0ekHkYjAT
VEcmwIu3gzIEvX3QNExmtVrtv1VaW5aJztHxbVEOpUKQ1OjZHLTr8ACjZNMh
aOsw2fs/ZIl7tf4VmLelQ6SmfuQ7LYnwZB1NJKgKvAx1e7QHiTxcnPcZZlST
6lJ2QHm/kVk2gAODwWROFYSgBRXmBbQZ89/ZSYDHhGWbyZcYqZfY2TPhSamO
H3YwOOXFG2bWi+CTspCpWkexg7/rp4FZbpUpsYHZxWKaZKURl2nYokBYb0IU
LZu63jL1c3wg5qMeatwJAi9zQjrnym2vptlZuqQ4aZTqjJLkWn/3i66xmt5P
bs076EK91IwYtCFkQ4IZVoNUPNCZD0BJGzAwrtz6KcoSNairhtszyNtQkg2Z
liw2mmB3jaSJcUZOZSmjbGFNK6LfgtaUQFx7mtfdZkvJeBEPPd/uDCmtr61H
NookuENrxkhLRKRZwLUK/xiyJ5VV8il2mv4pNzXfrVfb7NV57VNLlK9Ba/Q9
uRmbScgmeSK/Rx6X+2scWtQ3Ene0SpGabjMfuHUxcSFyG0ECdnoWCpKlzcP7
L/BIKGww0KZQIBpIX87EYnXfLv1jql6frpHTlVjjob/MaZy0llvnvfOVeTO5
XzgDBRt/Xdo+XAFfxtQDy08l0Pd7BGh+MQNf7S4cCFgCMbLWKwlT3R6TWZbH
UnYr26rMeuA2npcKWlYDEZwH1hmJxiJYmiEpVWLZdB6nXDOY9XVsCArkmg1V
yarLjZY8oax0Yah7xxUwmCTyVUL9KrwHTvidlgXZZlU/iqgQeg1NuCFYpsTJ
B2qPnoNh1HkrVpzN48NZLiyLNo0y/2VVeIS8UBmNwUKUPmBaC6/Oj61b0DH7
qhBhzEBtKXaPhro9RV1sWCtMeFeyYn220bveaoi5YHsyb7ihtaj75PkB3nYu
lwmosT+iL8ppTVphM8LXsPPmk5R6nOcucw1E3UV3BNpaV0UZlKuUIPpay1y9
Ih8N0VVoXYmp6ViwFUB1mYFalMjUhPorRXcPolUrqxPMp+ljIzVFd8XTRga0
xGGXAB4B6gy2R3PiixKf7NKtr6fIyu29MzURZs2wL2GBdBW049vZmehO+rQI
yXymusy5gzx5XM+a5VenlkSBpmhbOicSOn44+f1WO2+3FooVA6WGXrAJcdna
VjGA3ZACPFpguWdvJdSVo3FM8leAEI5HDba3UrBBxdUqkyQSA2yiFATx37D+
RM5WXc7uzKRy5oXR6TFbZFv0jlqE4D2NKYpXdDx7CzQ87D5n4OlKHN3VppsP
X6fhR+loXt5ShjNWweH2VSkJqy6IpaSDh96MrFF0chWr02qo5GqRgV1IK2AS
qRs0qV3PM73iI54BI61QnXLEr2XA+MZWbH6mXWLyXZhXou8l1a5ECChcKMRZ
cvXE3gj8tgu2fYSiwKjGXv9DEU0hJWRtoe7JOm5g3Arg4X39gGyLTGxcUu5+
1vFwKmnj13ivcD3OEMNbn0+FjSeBO+c9dxKErIv2v0wkYCeppSMzLPO6WoCz
q6SpZkuG0IMlaoJfwnXlwwMPljml0lM8+WGIcZXbDzFD4ofJ7Lul8879bgpt
p6DXHqkiTCyzTi6xBx/VuDuUJhUBCrcE4OQejDjQwVZEP+Rr3e1dEkTfHeio
r8VPxRW+tI1zC1eGjaV3Y0IW2+EGR1DFtt8ZWVLoYkEx9AklEDl1iFjO/or9
L+6vQ1L0kD2/u6aJujkJ4VnaFxPQVg9IgK6y+3CebAQyN2WTOo0MlxEBUtYn
Y0ziXvUYb7yKIixHPGfN18+nBarI8PxXGvvSiDSQuF401eFnBImlwmE8yanD
TO+eXCF+mzPjxGnxTbx1nHHm5+BRmbzGJDZ+n3HIt5Lwtl0+g3ui56VTnPZa
KLvg5LGesBg9m7dF2ljJv5V2HGGvStZ2OXJk01bweLzp4d5UjhSj46dTVijI
R9T0ovEQa2O5wGI7JyEGiOEdQfAbffEuK3OYBIofIzX8ana4bjGhaTVqNJbO
j7bILtE6O66zYNiP/e7tpICC7xrb9cm4PpicNZJlhe0m27O5t5n6y+BO46Z9
Rw9mCEa3zoei3uxhmSiXcPfGxKm2r+pnNQelL2w83PCNQ1zp4tD4tJj2r5Ef
GsERUFx+3HnpBwvHsGlok1zMqGMOahOnRmEq4liAwwCCz04AFSjPnG5nFOAk
Ke8Pm9G+JZWRolbDJ01DolCDyeTddIvG3NZwKIs6QHliG99H54pAuEcEK7z5
yx0NP2apyvxksCfWZDLQguhuY3kpXqn8YdzJ7g5bDTb5Yaudma9Zvnoisl2Z
jfz2LmK/lZNB3XQTloBPsRQ/nka3pBoIuiw6fLRNBHvi4nQlTL1bzuk66l9B
UAGMmI5gK4jZMtQ7QSq+5CPO9DTAHpc5F8IhxPtDm7zBOIu8jlhWIJ+F+7+7
b4+W6ZRlTDKnmd9gPnBRSOZzVk4aexPXT+FbZ5pLhbjLvqPgS1MUNPBjvUeY
gOSKE8GmcNilL0v+Naqk0+8iFif3asodoORHvO0t5YBA0oPVvxJZlBQbgg7M
tuWIE6Hjdz0qNV6Yx/PAbJsO2ZOTQZjHTEeCarNPP2M1u3ktwQDHDlzf6Wn8
xTA/1sByJlmVgHcHDYvdMsalbpLBTcoc+5TiUAd5ukmKJUSU4mnRQLzb0yxf
08NJ3agJvApJpfrGjyLDfuZICp8TvHJkxJivEuL0deoskaMPCYzxtCFBowB4
e3iRz+gY56msNL1G4fY99hBmm1BW8g0LEGGbpRyiqqzWADv9IWvUE/KHwUKZ
wspDTRh+IPxYSFo8wjifp1MNFENFRpR1c8s+1IJfozCTm1KhOfVTwjKErsyf
hg5EuCDiXtWfhDzEVL0KBsHnuIbMJJQFRfw0tcGGyseHXwlvwLh2kUJyRDHq
r2MqPGYYxsk1A2Vfd0QLEAt3xp/Y94csEPfuQjRq5Qkd23UasaY5/2qmGBGq
Q0ePd255uCvkAw09uqQPiDGDPTV1oKLxMK3jdDDCfN2pabdMxioQiTYQZd9Z
oiOU5KR7Z87FOMtmyhsNdJKYwcb56ndctkRWTFqu+H7ykhEXKA457/ORLUIq
B9f3rA+m2xhKrnuvF1STArvgCeSi0cP4ew8/v3rXBenPq8t62+/q+wFQ7fnG
iRJIKfC56iI/OsU/Cmzacd6nXpyYYQYzZkUt5Woc0S5+sqIpGzc3DXMsuqaH
08TD87qs7TSb/qEKcs/gjxRGf49VxfX/ZX5nGWQYyJyRFgG9XFtAhwdEPJcK
aqkUNj2ibQfo8fkuhlHrgX2ovCvOqTumry1EoMG+tjjphujGbVvmIIGrMyKi
buNmqkNr6eRrgnDJZhIE5KRErM9qOdjgV+Y3vsi8+XekUqRefbF6UIQPRGWC
kTe4WDAjvTTONl3aEZ/Ou8Dr1sHzTpIZcakUnasuofnikPX6liD3MdKovPat
6sKXklLpys6/GQX2NJRSL9c9HhbKfpgic5PU1btAoof49HObKrbsWvO+1XDK
alYmL3YUbDAI8Xl8iegiJNaH9MRBDeVOK9/KYfW9wE5qkgQU/EiXLaiYJoww
vaSRaD17HXO+SGNMLyfR6+1Vw1B/orcypbJA5lz0x5373iRdDuHf56yMAjR/
4LU6X/cGuhhpfgu4lRtcEdiwQq9lseBY8zzTJvvCINjJCw1U0b4w9cV0cS/i
1fho0vnLryjXPbL6WpnCPk8U00xBcWPH1wNaco8d7UwAG1FF7pfblTDczVzH
Jk0npfCn2UmKnh3EyMVx4tfsurZKLX3o7Ts9kCTwC9N/2zIIBvqpzTk8DD9e
ozpN+jBt+ywbAKAarcCDkN2LATjsrtrJr5tETB7ciEfeHhEGvA0vEpjujC5x
IHVRorIkt9mBAC+NuS52HBl18Jjqq4otYJ+3qF0Gz3YCk59P3YN1jlmDiDog
lgRFnc/AdWti3t1so01HbyxfW7NbP0WtuMCRagGp+dW02v1UsB0tktIi8PfK
xw+Si6g51CWK5+X2flEr0MSsilWW65ROisXKyjYx9RIQqToGCG8lrrMUmeUM
BjsUJqnDArVZSNf0JnDQSp1C6ia2TVc/2mRn6uEGuak2S+B0CZ6qew3d3L90
gsxJiL91mQAup4NLkMbGPnHkKz2LAOwm1qzcpCebKODQLCkmNOR2vicii72Z
BJyMhEB+HVAXbJIYMfXXMQqEkl0OCxpf2KEFF5bbLJVQV/QDLOF8EwUThH4R
AJbE1COC+y3jYxQoi8UNhSgM2olLpj2xj3NjQzHvuRLjfA08QSU2GJak90s0
POdwpZ7cZpl/kgXu1h7IQMnH68twYP4H/rsCCCiKtNrlEeHfKW2VuGkaLXF6
FKR1MnxhdbxZSP0S1nh76B5dM4nBtnl02yPg7ckSXP6KqLTs58Agm8mcUvUV
OKOnZUbXPT3fcYZ++iXApkhYZXaDAZUCA2Myb5xFuO78Lq6vCu8PV6YAB+hw
8xNKm6HB/2bqXQXiKUwfNFPQeajbJO55jDIRo6KAhK5JNvawUgpw+qIFPq8W
bNyV7S1Gh2vEIxR9UiVejqjnzrAV9CrtOecTcagnT9WyJhoy0JpFmjfh+u3G
pvDjOGUin0TDCiUbOVRqyiq/9Krlb0l2YUPYykkALi/XC8MXq6iIjLfEKexO
38Sk5kB+nfVch+/sbCY1zGXSuJKp3iL60f1h1DkN+sqsCMTN+mmA3m4zZKjq
R/3xuhM3/SNSm4lKeKrfLs8UzOG0nst1cD3h8E1/foMWx0Zo2Pdob/PkEa/O
S0mQahiz74FZ+W84y7dY7zLem/oo/dwfqe8ECmkRKJkQywivoV0HxVmKkasm
DJF+8CaZHhrRRdhhAtjLt66m3UwVLh7YDomWGkUOvZm30S8y3CkhxVWsq25d
s/r/yF+USXJN5PEj7RVWREOp6AMQ6tG2Z27NmDlkTg/Q4nftXisiHBrfcb4Q
wBv02cgtqBJy+QoiJ3BtpZeYqFVBytKPmuJFwASCrJiHWDTy20KA2cLyBIex
W+t1/Lim1Xu5XfQ9d0gRQHL6omopajdkceMjtzhp2Eu4O5YjXfwghQtCWhT6
nT3oN3uo9y9BmMCpSo/eBUi5W9AAG75RdEIQawgztQCi9NTFFKDpzMbz3tz9
z207MaVfoYDP2ztk9GNnLCkHyYOMAf3pG4IiLthTSUjqtPa3nmQjnxCkGEjb
rY16zs+GfyLrV/T70stRzxEErEdiPGN84aUS+fuQdaEw+5RfHniirK0EjPTQ
LsoD3t7kc0X90ruzFIjB09p8YA3z6EGsp33JnHuNfyl7q+jL9PEnSiPPOAif
P9hlYmpu/r8kOXCT87113PT5+iLqM/rsdrVeQr/yQf+AcmTOYKgAENKPmqZf
jGmx232tm0wYcG7vLtOxaVtv6xAEA5SzWSENeldQ0+5f07S/Ap1ehUUld073
DCmBecMn9tZ6+ZjTn3xV6pLF1KdE4qBYFaYXQKBvWwjS40WwjR5YlUMblt+s
nxNOEf6S3Tc05Akpz/OkNBcAeJ/ZJgv/LapDcRWfJ98lkYpaZaV4newXhjEi
XZGwser+9kQ2XTnhPww6KpsjyesZgcg/pv1L8rCRExDoN95mhPohkBEA9yfi
ncHYTBWhY/VOyUFLpkokO/9U4KgQxG6pPag55UDVkg97fKll48LcaWsdECFr
gxK81RkP4FkMpGS7LuumXi19omIB0uStwFkxUp0HbJb4i3huz++2wzNFLrGB
J6uPhrN9tlKnwfxX+cdHF73Rtjbp9Poldn7BDa9ulFbJvmuEPSUlpf624sT4
omONXIz6c0qUU5jNdVOzLLmig1hXDjpPUcZlg6Oq5Qz6d+IWTpJ/EX/ThiTn
uLJ18SlGDQBkWV5FRZKDeA16H4pcaOtHJ9ANWI8DYB564QvY3Y6Fgi0R06iw
b0ywQIp3JtOqY+z5wOXJRh2vm3GgseiT2LarAY0bnh8t5zuUODoQlMSM0Bmv
oMssLQB4pVVo1/FOThkevg8h9lcsMyrYEiEhaSajT8PDQUe/723CFl+g56fl
GSqBUms0xOyE/j6w9GTdindB29ibozeeNBd96b0zMC2TELBwD/agDFSChAcr
T17dbQWFkuBxXaclMDF3uq5fBByl5dU4+8XJl90memU11IH0oOKeEnhMmTYT
YUDCPdK9Bv3NjvZhPDQYXiDxavaFKSX7TX3IbGgS3DD8oiag7BB6vaC3vP0z
Lt2VjhtQn63+9qk3BvbU0r7r4aNT2x9XZc0HjkRH4y+VKcv1xpnCs4A0Citg
W14r2diKVaitlK5C7AEcGV1GEi08/nRZCMmM5ahWErRDTEOuijXVxm6pi/eG
VD62oMftI7oTY5pFfI+a4zNteCD8f+Gho/4FUx2Ub67UXqNIE9fn5OoN9IPQ
LNT4hdeCN9OVIwQ19ajMjCd9NbMVdJ6E+tIav5eBM6IDI6vicbm7gbPQ/4Jh
eaYZqRUL5QhxcqZnhHEfk1g/ZBBTIeIBgqmq+CBS321p872TjJKABhU3s/JS
wkF613tap5BrDSYNcT3ZvoMVjzJcAnQrOML5iw31wi35HUg5Ah5TzDMgcbWe
RRaRWPhOBB6cGv+i7tqdzTSDVuz7U1AokA7YqpQOXCIrxXXh7HPWVrfdN9nq
Y1B+Bl1Ce9qpKzu6lzooEXB9WICZ5SlDqP6mUakl4KI9gYCKa0GkYQwjou7D
m5BwTXQ7C7vpuDvxxpC15NaO79QjRWecAxqgFc34flfd/f0FB9BBPzrokECH
lny4b2Re5bCICbIKqrk7oSJ2pz6iwiO+T7WBV2PK6GtNcJv8vHUh7K2+mHVO
WQ9ZswxRxVhMC03I3OPGp+CjHfAYA4e9nECWNp6dzxRCbZ1Tv12mGR8npzuQ
gMNp7tdaCs+QuOgL6xE75z5UQENBRKut+SVt5LhyH1LL31rCENutSU9hH0UN
sbdgOlN2cV7p/YvBkK9iJ8a1WtgfCmoQI4r3BuxYLbXWp/6SgxMonTy1Zt+G
vlkri9/ciDQREITIvx/P5NOG1KGBzokEqkJxaz4FRZLYWSDcKb7T/fd65DVs
5O+B3T44r7r0kqlAkSdrhuREZyIUd+9sOK9Y3RdBdtH+PbMUvbok293T/9UP
b9zsZwUQ2G0+ZZ4Qx2izrYiz1DFaUZh19IF7qmZlbiZBR1jAL7jhlEZsk+f8
FpJMkk2LZfu8Yj41kZzlPcBg4m/TCAlzh8+dSB2eASlRBmSyx/x+MeY3qSzB
pPmSMuHp+zHsPb8VDR/CjzaTNCNzc9xzqtObDO6tfMo4pcoI4Yut5f82p48C
VJdzAyETKAZQ9A+Dyr6IxPxvOob46HJSLLQ8lqHPpF5fSUhfNoq+mXDdaIxt
evHwf2THVnliYEg1i5dY8wgfR6dDYBrWU5UlpLz/zZCppYPW/BBjng7ZaXS2
Um7f/MViMqB/8D7rMuzcLD6DOravznyPC5ZD05kW3W0C63/bELhsMt/KVcpq
OcigZpohSyqloPT+UzKxYewyW2Gr+9y2KXwWcxSRgZFrv9Dsl+aJ6CmzNePW
+baY8JTIuR3g53etY2VoCzdG6gpFhTP1TeJEsrvZ1GfZBLNVW7DLYzir8e8m
wPhKdGk+wjus1yB1iKEfNy5YMWceL8+5wgDgOBvfslr/i7aXLN1H5wcdAaiq
bKRHdqecfHaD4WPCK8lAN9dtyfUtoW26zWyvDK/RQYzm413OxbH9f3o/eHdm
xFGcbfN3DlDimYAHTXIBUxdgeAen1h2fcgoBgo09Aa4mcLHUPxs1FC7ugCiU
vcuphc/kBmsEgMTbIF8wsj945w2LMxYQ8qRQHBBuMVyhGy919pc2r3KCD4Tm
gaMz+CXPYgJIVjr7sWIrmHH3Bd9hlOp3JaEkEvVO5ET4ewqNLsoWrOYsNmBM
pDV6FrVJohxAoOOUEoJJX7uN2fHHQXMDXEk3EwYTkye7o1RWRUG+96OrR6qd
Xd/bFKkNkfeQjKfKd7OEEYBSS2sMd5Ty761AbcPBB3ZObr1b/Oxr/Iq73qIJ
n2bsrordUjXgIgLcDWdv/LKys6JAJDG0d7zksqhFqCe4j/NDiiKjWHKGPPRG
6KpqUDlR3ITFnKmlrVnedpDUxDWXYVhx8qysTErS0Q40CiwLXjOYzudBVZZe
8s6d4jMjw9zkeVQafM2tkC14e5qwP0R1SPXDFrRlsHH9ME/QGyd3l0/Dflj0
rWyfbCUWka3vD8/RFwOKN/yaCgitcfGoePbnSeLrKzqx1MDx4Zn+A8HTQeG+
QgBgd9SvMnwYjpHHFJGGqSTsF4eDH3QHjLJAzFUpKD9GoKQI8/jWQc8SrsHt
Oz/ejv11DLy2Sk+GuGAR64PinkD33RFelXbSoaUvbcMP78uUBlEHeehaNRgp
G4VcFXdOrU4THMkgN9MnU4ekzyylNDEOEHXsMZsuLwOq/b9gP7QiXxuDGhE0
FW3maR9Z+qjvxKSmFKtEh2bK2IA6RSuyOUgzaxqCTPBVdOQPe2TraeNHFBGU
ik/7Xt89Mkj+wshri3PC5DhxbMVwuQDkVCcN7ORbb3DNG5XKLkccP0qZf/I3
BpB20ZLSrtPoHiTlW/K7PSzLy0CuLJy6DUfdS5jubZBue/HUPbD1JKQBWWAo
ZipyGFDJditoKUQOm3rpDxPwALWh/8GxjKuVgxluvKWu7/+9ES9CVoJAgZwj
li4cA5qH/KR8jTQq3jKEYYAAJc4r9W2+kkfu1gTXrz9gPME2qYyvSc5R+Vm2
MTY9tQPFCBTfbn8UoUKFiHAzG5jtV8AfHOLD8gpY1PiWZXuuneMTyQVawhKZ
+t+Ju4K5CP3FrXsnsZcHITzOTMpTtL5bMar28ZQ9FF8PpSTUXXwe3oOVk20V
VOXV+TfeuDZ/FqW5Pa27VAiDN/CUHFY1Og7EbCBTy0yYejt04DEWwCUTzNC4
VKWPmm2aRjctOoivIklNSkpeTkpQ3Jbe/0bKKSysGOPbL7NDR5yOvAPJzlIH
nQoqVeO2IKYnOx1P4HgEjytiiZks+fdnRe/B+/NEEeqbSqyYpfAFQR7WYS7H
O1O+pfClxpnlgX+z0pwLVteaBWLdOn0k9WQsKszr1cq06bjI5iI80SOMVg5H
UBmeS2vKNh+oFAEC0VQybDoB4oWLd3AJteR6hvxc2zBhpHKyPLt5BTmSC1kh
UOft2OVUeyKq3F7wNoxSrohJ1MtTK7kX4x6HleLD9+qPNV9GuEKbsUDGZ0B1
FatlgYDN7+fj5ctx/umzeK94kZAgM4e4euwBNblByi5NGVdNWILQ0Sydq4YC
jKGOnzv2TfXPwgBnBzWFIOxg4o7LmpCrdSUx7qU9qzATWSe+b0T00ruPVRSp
0KQrGdCSeo9oioCo5qMO+vI5EuXuSH15n/FIr0+Itq+zb4Kcezwm4ekgYLXe
OVpyKeslhTymAr5ULeZPY/4gnopGEyW5h/nSn2mnYMYBMG2ZWHSUXmkoSLSa
nrr32PCe1PejgonxcYQ6HkYuxBzyW819mButcJ8MrFXA2MyMTudVzn9xLHFq
dYxDtqY4sfqLVMG0JgaZT8RbFz9xbrAWFyLDUFLql6FjrQLCnBofpR+k7r8T
0XMn2dl71vUl2azuLV0YRQu5O9wBpr6W8b2VJr9EFcixX0GIp2VfIOABccdB
u3LOZR6cVDa+ysjjPgWp2V8gp8S8NqITvUOHDtIpiwORUBx3AHRcFXeLm6AN
pZ+ntgoZoJv8vmCnhcjB/RgeGKqG2zm5VwGBdJyts00AWhSVP50Ni8oOgL/a
HkO2yike4hPKPRUqrN/iZMqeDTzbErJ3eNbu65E08HQ3yX89ucgLTI+zEjev
ENa8AYWd5rPwIiOi3gCqFArcV9lTuJGDS6WJ+tGb1I+bfd36Su4R/B253kln
4DcsrngMtmQw+mlNC/iEZKLahbdYdedLMCP8vJzYVDmbyTdxUfrjSpkGm5RE
921JaPvP78FqmMSx5fbQ65N+puLP3CUWrjFszBeqdGAEzQrMad8v2xtvM9Ke
CvxuA9kBXS3bhF2ZeVlPo6X+L+BZ35KWbYQEHTSiP+Sg9HtLxuFQJbjtacpQ
W/i8/43JSujep9nj80pMFXCjfwvM+aAg6dqojqkVY+v8iHgEbcDHx8WSsVgJ
0f7OqbVFdW2X95v+3VYUj5jHrQx3dj2SvCGtUdP/V3cn8i7nX9g0YRoINLRL
WSPLa42qSM0YDSwOVVUZsg5WxjEUjbqK/h4E4ekYHe2GI7CnqddSVfKBsA3g
si+JO4fHFYQZRU7P00PaxL5wsKYMd7K0fpLil8Ux6CFlpj9Ecae9oLs85dT0
CLRok5Icu4vK71NtB9vySGVXVfH48zuZEm/bEfWJrSiVcrx4+zaS0NQmOj8f
1HYXQpN2Jw2/VsnsKihsXu2FFHyFntiNNDhNt0pjkwBp17nKPXVzjo0Mgj6c
bD9rLuh8T02xNyU85FhSwGojUi60Ly6HQ3T67xPGg1WpOfxhKHKyRapJiKBT
iXqhx+ibwInMSxbkJ2RW1kqdVmSg5flqEiOuBbOsiN8AnIDA4JQxcCjHzc09
M7ja25LyHKQsjaMUHHxwvllFsh7F2NFVRV9/4S7mOpubXmeJHBXTAIrCtNA9
xcdn29CQbwh3GlM+RoFn3PeU391Un4tlAY00G5ZeoB3YEMKp8Xzq5BCtRKBv
ahsAsNim7cmJExyHgm+GNbg2YfW1luDWhLRYh43ae7PWm51aodwAxfPVMSc0
etqMdGRYYtC7lnfNESrBsXbrpNhy8BOjvzdOqs2kEtcHNeiw3VoX3soqWbjj
g2U6Ns5tn4nE8QCVR5UsrRDkxjMkL2W8pDU5MNZ3gyMMtPrm10daGjFLMrfv
szRTgZY0BiMeitcwtlnODpY2Vja2gC5nQygjwjew5nFWWBqbNwpMsVqbKU+1
yaNixEAkpNw6B6ZblhgfJhXznqbUIf94RIVhBhYj0r9f+vSZdOCfq5b9urch
CbnOUnjD5ko/0QnBuzCKITKYG+VdUZl5/5rz6JQP0QspOXKTOycSzl5SWr7Q
EEKdFm0hwmQRymmeDCO7mt5on4647sqeY4yIirhNSSrRrVUXLg4mdHqTvanl
JtIMyFErurHSX0/TgrsIe2S06w1W9srkiRIulxB8mSXn7p69QYSJ5Yrz2rdB
MoSnhWV82sEDB7Mhl7JNrb/M0gi1Ha9ngf4V62D8m2mDtyHBDNcJxjVdaL7K
2+ImxO3rbeD6cQvEMt1xBPDDrgd4PdG2P85PJTxZoSMgLvsVm9bHimKTmaEi
fAvicZ+aykkY1G1PG48zFWa8yO5sSEnYo43W8icZxF126RCYDtyTz6G2itBo
JVJ1Y1oNCfL40i5NRbtqBJGR/6XBrTPryr8eQovXXtkeNY+BJU0RXbY1XPet
OMBLIHkcX+Yvfl+0PzDbDXHOeF0EKyJpQQ+H09IMUaV9unxuGtJ+vRdl/JKi
Qenj+/ZBuQd9z8nS+sHG87nRgBm0wU9w+Zsm6/OOGKif6aFVptK1zI1LP3vu
VY6k5CmmNoCt/4CRfPjfCjOTpNby72RiNJaCPmRxBWQy3AmCBUb6huD+2w0h
xiOpjqeKAxXDhXBHuOpwHRPyVLL3Fdv9N9Bzn7Xyk7NJIx/E6Borgi0aA1fQ
fPSXkclXM9IOWi5PuWdiu0KpsYJzpjTQ4k3/Ilc98d5TToHdWlP3pC5I3x7/
tY3ReXTcSvkRLje3hEwCSdnC6tWUfzM+rOrl6tIP4ROM4455BjM6xFyy2eex
K7RafMnO8IhEELyf62ez9CvkRr4fTRv+ejHxmViid3QzmutM+6jRes0hzqMA
94l43tgohZ6MamYBTG/WAmxRMQutBMX25OH/DO3TQrKmInPK3aSNDXjQQVwX
cjsJ3mLgi9AoBlqBcIoLxEsCzyfY37nAEbJcQSZdbPHK7rZYf5PtwD8KKASW
wxHAZgAhxtQjJ7e5aDaorwbfvmlj68bpZEbVpTfbYiJZCI/x+v17upoj5Kql
L6v4mSV+Xh+R0fU1AJjxHwrTW5ygltZWnHH5Kkuj/oxQFJxmV/xuj0rDmMki
+ZkOFezkiWxtocj7lVQjG00vNYmAXG8ih6o3OtxTDAdn/ITaYK+lNvqPSXvd
5YrHGJVtP+uAvh5V5o2oNUw8MK17vwGz77BKtqueFwqqhh1Xf2Hl11x/CG2H
8TMd490Xpmvz51iuNhVBe5YDMxaqAcrY0xJBYHrIT+JXx322sp1i9J4ciGk9
VfiwZu5OEkN9NcX92f8AQL5oY57aI5RzW9H3Dxwz8ZtpnAnRhbYYxM+xfEnx
/PTzgJUP+6GtHTRWc4MTUaleKHVQqNRqB4Z1tSIDdQkyDdUh5+KpI/fOnqXh
GSABGa2Bf0DX+qEwkPjYPvxupSBHl95XLAtKZyP5XQZwklgf423M1bD3hCp6
BjbcRNpB2f76J0MkwZm3LLPKadD0nW9ZoNvTT4xSTo8R/MzTU4U7sgln41Yf
NI1F3KqmD32gc5TfEfHu2afTFlzZipfLW11F1WFUC15aJAyatNFSQ7Ukre+k
ZCN7iR2M+BxpGpyLVvsORhq4isQWXGiyL8MB6m6CG55GwiZL7qpAG1gRhIAW
vU2hT5/Np5Eohq4ggIYrjtPhSJl3Qt1627BweiKr16n7aeDgHt5bfMKhWoa3
lRkt0DRyUS1jRA7IHG69VqQ+lqsZQWpNy/RDecHRM8pLAM++ak5ThyZpdfMi
9ovdhPZCJNQQxoRj32D9VKvWyIdV7e3kBFvtktASLlooIPyCmk7XwQ46BmzA
BoT32zd2REKrW/zLbmvNl1UsWEULEVefkDx4Zljc15P4lU+1k3tqwfZTWj9k
n9DsPM9suilC5CPrD2z5CxbEH4Bo9rKJQebMQhltVSAyLWM/8wdJ6OZt9Kdz
3k2iRrwEOWQSl9jujoPG/EaNENSu82697qcVXYJwPWXPlj+k/NMYt+powKhL
ivQj3TIAcnGkKCaMbmfBs7N7AmPjQlsiDC8zsBkd4bwKUXJaLnJyZnH09rCJ
FzcfJ7XX9/kXs1F3m0k315PtDoFMVZCv3vwisvvD6d8d3uwhFs9V+97ozqc8
shvHm1w60mYNDlcVe46Ja/Sd+ge2ue7hUFUNXg/EZpqhP++QpO5EFIYiBuMm
N+RU4ErICScAvHCP3CksideObblvz1UMSRfPUFovTB1VglKA7hdGcj8KjaPB
PU4PydlnoLu9VNR5GUFNUAqbbzyOU5UtleLQ3ukzzbdnrwdAZgEhG09c0sgm
TN/Dbk0WI5VUsanCIVCdR0xh4MEuU7Qow1nVitAku+1GQROxUqvl0j31UpOo
sDId8Hv3auX4Zwj6bO5O3jKcL/SoxAAoBwWJgyVAap4Qf9G3hy2+YLpAnc/x
RdInflAb+V2UDPfLyJqCqewLv+0E9Wvz0uqIV62xjwgwUbeyXFeowELn3YSZ
K/0ohZpYEpbph26GdZNs6XHUw2Dnda+DdqmNH8eiQcs5R5imIB7D2PQY19lK
jCOtGsnPhraDZBq1a4Fs5ZKTv/rdiFahfZcl9+m02PZvl3nKmK7iLMAJJQZn
OLd7mpM65d9uELFUTowcvFTqm+vm70HLv+TY8zI6MSkolDju2cXvzbGUMMoD
fqlzIyu7X/GfPPxiEqyOk0j8o6DtB424ajVEyBkMLEnOKCQ2eHtagVLX3aMa
Sti1aL0QO6RLhLM9zEWwAWQv7hT9nP3pvtU9/1Cg8K95IZvQ/SSszvQhyRPB
LnbLGqb4dUDM40eqjrYZqsJbTZyXhp9oedMP85cL2r7jUT3IfUn818CgTt+V
4r4xzSpIp24rD0m8k193Uix2x5y0eNRlOxQndb4+Mz3ViYVHVPly0T70E2Kb
CakRaoOLPNk0kIZG7W0enE1m4xGHWJkDzg4nonhziG1GFoe591gXALIk+0s6
fAB32gq3RXB2m7yPyanVdi5qE0NRkI3/WILMLpFCImSOeudLXsQ62jupgi7Y
SpiBi1C1bps+1lk/D/Ts4hdGqSQPrxJQ0k2Yd688kCB5+yK8Pzs3fi2QMil5
3aYOFPSk4fLDKD11WyTVv4q2ArFOWEeCwLYv96Lo0O5EE4dgS4WJGq+ZmRhz
Iw0J+ZZYDKzMyYDqtqB3SUqP5/VxI811IE2C8SBql25MGM5kMz1RHpWL9+EV
fZUx2+irWhWuPCLd2uh3ikUdZ4pGT1hQC/uSH7X1WJI4b7+S7nOPPx0FNDlU
iXEhQBnDulOA1QeWqc7oOuKPZoa4032hOVdJXQ7MPmB1zS9i2lA4xNhpOfau
KBNkZLMOzXvuDokrJeT31COGR6eF6EuEb8sb3t8UlKU4IupqIGqO98NDTCX7
pXdNZzzD/yPj8QdU2FhEHFIq//ogGsIb4a9eZbbzJZ99lyRAxvTZxv6TMlM/
mjJJ+1PdDFIgjAi4RfqCT64QyEsleJGWq+B5Yoa521V9zMw3F3W7YM5nzbMi
7aGkIo+2rA95EVYIiAt2To85IGIBE3syslYRLuhiOSAPtFb4RK4gJ4E7KeZf
IyhvNG/gcLhDu7Xa7NPXkoVJPaZlcFA5FjHkLpXKXG+NvXYbP+OQPKzwRqWe
rR35bZrBkpAjpNUD5uwxmIybIp77wYr110xl+5+GQ1FfgEuJ3XlqK7mXgDfM
uQ3abvaYIReOfEltQ6UtYSzq5wv9WtC9a5LNqPBBoPUE7AAUW8F/nCF3KYZU
cgw/zhfRjbEo43sNYqPOoZaztlwlgV28tgkferlcCyw7gYT2ImBaTH7hByH1
7/hqGyPCvXL9MO5MtsTGZuL/lE3YZR7hUA1c1qO8DKZO63FQngRkeZImFTzC
tzPAyIkcX1UWz7IzvgBKW/wxdGwFr3zcdfmxlPXjVDsONtYFPb3WbwDaTFHU
NgQLfXxN2siOpeafBl/Pueqpb4DYYcXNzsSIzD5gK8F6Ic1Z8DFrgoIjAdEl
J+NOD4s4Tng5zi2np5h10WXzv3pCkiukbm76BqjOopokiuLeG9GHf4RcQfhp
m9VsYFKcZAsMmRKhsXCMrw7/R5t0heUPuvftTr1ZvJZV1r4VABGT2AX2hEGK
2WOJDLLWy/qI8xpiIoGPipbs7i6JGcToaBrEemICeaYHW1TAp9LjXAP5kB0F
3tAffNvzgjKMW4CgovOPwCJGFvp0jOggkYZOIawATP1Ni2OTjDp8oeWY1ifh
Ic9xWBwvL8LDQhvNPZZdtEHxjaklbWy2+QGtjJSWPJg/dj3NwNz9ULTuxHia
lNNcjLPTk+27yVvCTPapaWuKVhPMniNIB3lG7qqVQgA8ZcgHPGNbpLy1rXhC
JhskcvwpeCDUutQvT6anOxkACHySuG4Xgwbkg2NkmCvYRmHT7INL2MuzX4L9
cKdJL6tum1oxqseB3BeqrFvkprKn7vVcsnSZ31HabkXsoUBimyMyvuUpIITy
IgDndksKiwxBvWBpWOk+75gZCHGSgyKnmAsa4GuErzduHljpoqLiHvlXTP4e
YZHeHkVEf6VOulwyQnRjbRqE9wm+4cFUtUQGhvfkXr25Uza83W/zmdXvVJ//
vuvc0Xu7I27NtJl7y1Wq5IbW9DspK8S7GXBidq0b88626dKkkFzJyjAyG6Ry
46YM3bpN4AoftL/JCT3lKc87ijBu/EgqdrQmpEBTM4iKdWfnW8+xCbTM6JQY
l459PCBfAn3qa+pb+ld2XMeAFF+1S8vSiJLcJLM/GAwY3CCL6K36dor/kDgL
9pjuVvgNSHRDPNumHLIlXaRvCtUrzOtoKEDS1fuXrYmFxZGn3XBZ53TxO6PG
Xdb7KYDSnuaAnrHAxMx2fRCGLhhDZMiiZlMLhtX9lLl1initN7dIwYlLKVOs
Dneeq7Pcfk4xyy4+g2r15cGNBvfPwQgpihgrOOa30e2Y6SCCPeXIQJ6q6JSg
Gelgsa1wIvpghunM782xtkTWh0UMjV+kN9GEN1JiSXr+TeL81/yTj2SkZ8Xs
Ix3tA8DzychOYm1kqxyWkzbkgpVPyU72qPaLFr5EqO1XS7Z8bfyjvKafP0EH
82VpfBtTTEP2gCdL05Br5Ev6QPGT/nPW5um0OAHCAD0u40xBKOylHQmCg643
PTcdRvyrg+w9GCjRxWrFUOgFnV7H01QALUPwo8e+bAjCyLkYZnFlhg5YNBw9
iybEfJZdXCJmbQXE86nsGUVkbJFDzrX2zOPZEAX7ITZ0ck3I1wVwnUv8U05e
H1NZRY1sAt2zAfj90q5RaPo4tQabAW+9xmffmEvloiAD4PNPB50R3JVkXOyl
0magsnXlRenmyuJWp2qi6zOD7GmeSAO9BGVV6T8CPv5nQVLeRR2VTe6CtM7O
d13ibxPquOzY1H3hbYXtoDtAmMvM211iS77J2Da4Mc8+bHPao9ZfXAZEGT2P
fQXAXpVLz4lDkweWe0EKjiERHXsei4y3UFxgePZ22YuFlPdlb3EPb2uJ2KWc
5dy5iP0f5nTUPr88Df6crAgYCuI0GwB6aK503LYhjk6SELqkmJnoTy2tcBqq
hiyjmglXnDyB0kgp4MfXWd6agJ/TB3H081j8DCEV51dWGsKR2iQN9AHYgvT4
NFLoG2hrgxkaunrMGt/+Re4AvKa7DKpEZDTEPHK3wRWTIbupyzzekQ4i6uHu
GiuCtmWyQ1qbNYYEs3TaE4T40y/t5+5FkI21ZJ4cieUvFLcwTw1Rja03nhRt
RbTEh9oBGIfw8u3M8xPZSnrQ16KAma8kX0BybwwsDQROKlT1aNyT8v7zebs3
197VntbPHVDs3k2Qjn7lT085Dq8eY8783oBBKtlOg9spMohz3zextIpKjTMM
kmzjb2+lE+KOGpjGa3MeLdkpPnJKHfU2RVZxBjWYOt8BVfeSB4rYWpUwepv7
gcrUNyV2nvf7RzcdzjNajOuscw6jISGTgx/uuNL4jh1uJs+fbkb592pZ2MMI
inLPM/Fwt5cCsSmBMyVXUjPZ87Zn3EvLlQqZEhRGA7ON4Zp73CeXarg7w6TF
CYAIbZXicr2Tq2HCsI9yueEbcFLzVt8U5VZ66TfJRMdwzRfJ96ymtLjWlpMH
gAnPZNHFuvWXlNU2YtM02hYmE3l9c/KjCJVOn6mKMsXka/LO2afpqcRSn9M/
uLhi++oiZUiJBMBlnGi3NsuX+maLUwHMbj9DmqgeRRnAl+uSHDGYpI4rSVuE
btMNuxCEG1/ohCLIIq9ex6iJH37C1dGONuaCmJUYjf59c0UU9L802KFOOFY6
iUDgoGqm0S8dmyMpfWCPGc72g0l+ohX75dmbQ/EcKFCAHqLpIaCDUXiH9yjG
HpPAA7uixQB7hgsTM2RYPBty8j+Wnedt7JmtNryOPj5+zGZbp3AAx+uafsZA
tSvGYAjtTP5K8bnw09YGvQeaRTjvEe5blpPGpti0t01VrpBOi+X6CZ+ucZ6h
F1kNUqPU8/zndHtl4TMHQZ7gGhqzPK2Lrd8bhyjO5DtRGW9UDxWSP7rTc+o7
Ke5eCVPh1q4gpQgqTNtfGVfkDu93lpdkTRzMdCfsJybF++82snUPT27/JD9W
EhNSpUkicIMw8mJv6hwy+kS2aYGs5rxm2WjkQzDL0s5Fyew8deEp2DkgwL4Y
WG1qnRTK4iaUF0JdNw4oFDeRoXfjbPrxPRSV9JA02SOBO5XvrEEnD911LEJ2
aEIxzwAjvoqexPUxmUor+vDEge/rXqS9r3lB5DJUdQtiU+nDEcVS/LSTk9AJ
z4GGsx9yVHVlq8Vlyd09EcGhu3MPZ/1NQ7m4vpuUK4+tuUVc5K972e15Uco5
AnKJJZYzj99rYgiUZL8rF+o9Z8b73NLSRrW0VcACS6XE7HQIjS8TzekDvdKK
pvmX4Yoqz6eXXltgMhA6RBVD4XBBPk9GzVt8sfAi0/bDoLx2OQwuGcviNBCM
07Iwg0XCbZgy6+891e32Q2/bARmNSxIj0Kk7gUvemRgGKdbIrH2QsKAGVZvk
wM8DfPUh/2SRsLBmWnXzBbazcNrj5Erz+cj51rljrvW+p+4Ugh7x748dUS7S
hQHnlDPgqSq5UywVxEHWBaLp5FARYdRW2Tsq65vT8YdOcUot3hYwccOgCZ+F
Cgh0iLqWLwEIY3N+pmb4fplTS+zBRyJVIqGjUeYfYWN4tSBRQh96VjwmwHVX
Gk+OoQE//fj/kEG19tn0dTTTmwK6M1DUivP12/ejHAxakqgxQmyer36gz1d/
EbSH2XKiiBGbSuVhHalvKtF0BFMnFoUv95SZmTwJSNnjfiM8JUMXRWwqlneg
QdALzz38tVNJxlR1GJZDb1DfskZ61qpqzJknMoQfUqryNn8Uk/zLEDsZs64T
oR501vBiB/Fc+WFQ1Do8zmcymRdGVOpnAAWd2F/I+lWBNb5mlh9EPmUf5ixk
wxgLFtb6LxqXY5bwrLtRI7MWOPGO17dapl9+8yCXk7SE8VSGxjhBivz58/Wj
fLiVfoMPhYUyOXbnJjOnyn+aNQyUvRyb+VvDr6GMxGf7+gd90eNLFGHYCCqX
PCjPq+tMfN+3apk7Z0iYxZVkOfapfxJqdu/EUPRtXSBCSv0FmDVOTm8Zly9a
0PPFHRacAXQCMYHj+Cd6QWVaSRzuCPdZaxA4KJ/+C+4WT/T3BXOiFk9CMnp6
FchpCKpHnO7tPaVXFimKXfplLT5oEennnQ+p9HBvzZpA6Z1lpA+/wifO8IQT
XriEVm5BqEp975N8TQ9++IKaLSnD2rs9OJgr33Cs5bS4pEr6yqR+0Vl6nYuE
YR6hTistwwbN4rY8sm9iFbzzFeRDZpmob7FGye1GBd6RpebzZg72tDBwIaxt
+yhuTb6evLg+CwNG8kePaeR5wWITFEF/MrZ1UQS7+p3B69yWaUy2y+yQwuc5
AWhWuri/4McBkJm9tekT8Ke5tyAbMK/LMWsJiwHoANRjcvdSvNcIJ9QDYxQK
dn2uVKAG3GAs50ddCC1IrMaX01/HMrQNhguUeWa6FTQBBJZsbO72Q/AN1Z0k
Veno+JndsLLYgy0gXuHtOBUiNPb6ZYxQgEZio8wnb8odglp6jTqvtHJzYOp4
NlsgoFww+0xvU1r+nbL2l3a8OEnTTrmU5YLEveup+g3w/l25cnPK5lEXtjBD
s0J6O0vSqV5VhoqGzUTlLSltUC5SnvlaZ0zr1Vg63J44E/Z3y7ynylFV3fhi
5NLdUXFOQbUK7XPVI71ALYTYqQf3NAqKF+Fy19SAmWrQlebLtMWlQLkTr6+V
hllssPfIao1f8KN5+PFxMmyD5qIpOLdB3yUhiiNsHGFS7XLrFyriNgl6D7Iw
FZ4tfFkoWIDoXEQIWVP82/gQDu32Ln/OPJ87E4NZRMI1PNh89RH/gANWUhLw
OyLSN3ojUMMfPqMa6C4J6XPrge6acvBuvcN9JQcjLcBAe+p0qcgC+9yCO9yu
beTfK9ikMkGsStqyTx0dR6CwRIwUqXsLr/lAEf/+UwiwhJlxm4jh3Kn/fHNM
I41jL4/6C3cYsWZJAP+30SRmSuwNLLvoc1xG0eHqfdxovHsNFDiIw97EfGmS
TTIxgwPZcPdSEuWKyQqq9gkt2h1TX3e8mz928JVEGRwS9kpEwSA0oiVbUHBc
xEqGX08Crz4FuEEm5jYXnEK4TJPN5gZp0UzKCl68arBxfRSDQJxOG+rOMcm1
24wt0fTfjg994wUTQZdo5V0UBEt5KXcz1VDVPZ8LgSR0Y9BMOxHFBU/ZeDqB
URatpC1ROMG+5sVyM9wPTksdhjdTRFL5zJLSMr+vC6BAfxcqgajI+uq2dnLI
O7fzPXrm+3VbqN8C8Di5tyaHIxLCYd5uBSKFyJB4mb0xRyuXAJimjxVv4EB9
tgvWrCuGp24VOMClrhwWJjPd6QySEn13xbhX9SK4TJlODMA7olEzI7UEbRyG
TzKhamTK0yLxfae9OLoOg+MwM7Zfb2zhAeUGdkX4RQqkH5aMzJKoBmP3GnT4
98ko+dSiER/J3xx1sZ5QrMS4wDCZYl9Vp6rBaGc/ftc+av272xdn/8HfTZjI
HxgDeetVgF9Xy3rPyFsNLjpRzjdBjqKAQzhXuBAgk8gSWDBuAsDS3VRjbbBQ
FfUoGwDW2oyK9Z+fMsykjK+LNCOdZSOhnASE53JYxW2qjHG9//gauagl+cC9
iyBaJ9CKUtl9vBamQ5rOzbjKOuVw4iWHtY7QV1MThFR4iIO0OZn0vwNn8Da5
guc06OYggvX+N26DyfwvyqcsHv2eIjn/iX4HJFb7eyuep2gBFo/y2KDsUatQ
f4p6WAXiICARqkchLnkoIrvZmoJ8VyeS/uA16hWn3D7xVHLa00YMbHBMtf8x
NilTubs8t/13hDfRbmJJAEoqLbO41dcb8IhjBzx9HG1/anGwKxoiJsAWWZCp
OLtt9dcWsB1hUOuW60UY9QyylTq7aKi+pL1i7mp6BtCEgF4vVw0dnwFXUwh5
YgtZ/IbAVCTNywszt1+G5c2HNmgIas4BPmVhzvlatpDyBWnStJxlJN8mO7tg
HG4C87MJfPN1d9wMLaVy1IL//gXSv3uQn5+gGdExg0kD5kmb80p0D6s1C9as
cLihQ/muHEPXeFRvnfpVjXTULCwXpOxofyD6NkL48rQBAkqMjHr36LTXzisV
TL1MGO4EETpee+CFeww+7a/BUakQtHwJyksbl163bTpofg/JlsaNJ1YHa/1K
YCqlFhs3JYEGA+7QdiyVFxEYzAx+8O/eJw9U5mYWw5HoKsmwQxQCDPjLRpjH
WdpI/Hvm3AD82nkDzTAbOAcQhD3Us+fm26ylR9BaG3tnz8WNgputfXeB56Q8
KBnXesJR/ncVdUoOD3thqNkG/TBAEqn7J/miRIe0JjhE8wO+CraEj/UB3YND
+oNX73fGM2Mn55wzWiY6gIvimaF4W0tU4PvVbaxlkq5k6qElML8Ysuwbb3MF
zjOdjseMQbVAn7d6ZKNRn+KA5Hqj3pdx8kAP8y8qvZcyLgMrqs2LYWnWSF5o
vpFgk06arFCvHSSBq3M8scu6ATCXX+WMiTWcYlNLctklMQqYcLNtiK/oYado
lX9d5U8QA0ct4c6bON4u9bW/qFmKJqqz0n039g6gMkKBlNmwYB0OZ8m4Rsz1
hqsg32b/NeVNVMiDDVGUj32YJXfpxlx9vwwAEw9QiGeAQF/3ijIT1uZaXugu
muP8/LtAmfx69NhQqWHuO8mX0G8YRe9FwkD85lfTf9ab8w0sxRk4StU2pAI6
MnXGAtjhDgvI+DDZo2Cl2iH1z+zsr+jos4n77vJvGgzRUzpTHPQ9cKV4LUUk
knRZ3mNMYnwFbeC8t1bm9yOccZPNFddOQMaTJddMJlUVm+wHOyHxCiUbrZxP
vi22HWWbbVvqjU2u9vS7bYT7LK3w9w5gruRGMVhvfnM7qxi+YkkFKzhZPqyx
sIKo+r6aJ15zBGma7lQdx15Ywv/wwqS6Vm6YwuOhGid7LFWksmaXmKdV7LOO
DqNvc85e5o9tolcnWWgM/wnLt9zoLccB4Kl4Vc2rwy+kQ6NHXULhrB5XhrgE
lAdkSoTErui55Qrh5hdyt70xqpvOqiQI3fA9aTlRt9GCC58FBVmZYgrSs6Dh
K0GQRUgcbuxRACvVGarMQjg3ImM9ACZqYHylVZxtmme7H0cbSikAbNDnmNXE
zz4/znFqOckbQXh72Zm8pcCNxWRV9Z8ZE4MKiX7x8eg+3/clTgn9vzQyciab
GTH2fwQ0ixBJnfcgizaZeKB1bv8B+H0mR4+njex4GAYwQb+14L1T1NkveWvx
WKlYZ36WM8SLS64G+ofBrlHI56yzOnzktFd77ClxC8sFjQYALpuXXqysRu0Y
QSY+iq1RbSOPvVZLBvALpABf663qOhehbs7DPIdRKovxMld2wBxmRi7JHLdY
J3HJgYP6ukouqFn3tZY/8P9+efZlpVn1pYdGCssjcTMAldkYtjZosYydrFrF
+1ZDouQ6z/uhKHtjByNDmwD6W+kn6XpyD+rtd9WF4c91hJCR5YgHt3i9p/3n
ejW4u0vM8K/trJ9RHoPcNLQ6dYJVPXJRfaW8EGiS5Ho+0us5u/xnYflmefR7
O38qzmpbfk/w3xZc5B6xPN7jYHZRExegisnz4bBQCNdiwQCXtUawjwpenXOe
H3dpecFNjmNwoHM1jRf3KZoag+6nBq8QPYPSKjccIrgfOgmHlVfSx6RwG3PJ
LIwQxpe2DeNvnKfrKSP1XO0bObBctnZPO+awxXfmd8g0AfUNyDDAG2GjxL9Y
CVtAvmNtTvogiraObvb9MYjFjQCn5PxvvtdSMiOgbYWOpYVbRUbkOo9NH1yN
ruOAYn8GRInDLRhtyED0h4LkAf//P9SfGqXYEN07VZDmSZjUNsFPwE8inxaM
VPIhy5RXDVO7X/6rgXSqvHROR4foNj/LAe6bnExzORKiLVQ+gZ34lttPiuiN
uN/k2eIuEG7Rx+pVVwbT+myaC2AEVyCl3gFAia/EkTc1WQDif8dwKHCopJEO
Cc2hJdilZXoBtNsy1tujAUeyc1NFIeQZY+FuaarzktF4XI0o7jRwiIMwmrPa
V2PxPjqkEcBDkXRG9ZgtrKKWB6IwyU+22jTOnzFD1n26tnzwmgK5rZdIoSGs
k52UFgvrsldKI/xnm7rMkwmjuxVk7uIkEM4DqKcLT9JfqkPsNDCxH5nXLOjG
ULl6KhXOVgYM4hv2hfbWjqmAIXA9nK58b4O1qqi1kRdPKmyftjdDxpN5qjnk
cihxDzKM7fjaJvoweZwnbh84oTUeLh1P4WS8VaLcgkIWF7X2KTHMojCOxDr9
3a53c4f5HdzVsqt3ISR1KTOvCTHpKLJsYigsFtJQ8EMB1/EHfzsnQEz/6BwZ
1bNV1ZAJ2PcrNR9hPdvuTyNad/Ec+UBrXI7ATcwQ6c6geEC+Ds5IgUAW/6iu
G+HldsENXdySAQXVPumJM2MS1ua/RWrch/PEgDpC7jnXOeUxlNIRUh9LxTrK
t0czZuF06CuDgv3oKs1rQ1RYJD/h6882ZEhtnxEgTI/yaWqJ+jm7TBJnOhRk
SJO58XSsia78pkRHY3xFMwgic5LY+Rdl29L4453RHgJmXl/s+cYNcyQXlAcI
xKFX4BnyUwzJxBwX3nq8kqFCc9X25kXcmrsvQvKqcIGrx/EBYm6048eZq6sA
nCNofeRKNEZnP1uEzn3NgrCSu4SsbkJSEAveoxVP2LOjtH1v7GH6mtIy5mh7
3SUe1Y1yBVxjiOs9QGPEOam67yfWlHVrpqpb8jb0JBQFnpEGZy+Y4nM8utRw
hzVVanNDebcZRAdxjYc/fAvupEOvEe3wmdcK9UhtzYH+SCr/Ryvgm+tkISwy
dedvNPkO9K4cl6BmC+n4l46ph3SmfYCzrlVmmPHTz8D6klh7YXG29Yidd8HV
3BtZR4CLZt+rU//gFw8qMt6duVUbZdIGqSYjZMWDJAwnRFg1xoZnxWLqUe8B
WpSKhQ3ubCSMs2eXLIoebIaHPy6EzZfoOAtcGh2v85iUxZCgYXgGpyHDnltO
QhWe44ikopLnWFp+E/qkprl39UegvboPb+rbCXtkEAUslWabRUWSFY88rJIX
XXkdMJcutgJOVfdnabOzScQol0SLgh6GXPh4NbsQ3gvCP8cmbFtBG52xSxZH
0qzzpX1autiZC+fmaQQhC0A2MZD5HlGWyY4Vsnjp/50tjXJColAgpMzHK/1B
7X+BlZLo0adK/3ojjWnAhD1CXjTgpBOsqBs+p+NVhVN5TCtORLXQJStjL5Xr
mSOA223xXBSmqxBaD3pzgi3IYLIzO3WWyct9zFombLo6gxUZ+aQWp4VUc/6W
l1oZypapi/7yiASJhoOzAVIqqViKjT2BQdGZKiTVnTzyQGEIU5MjsNGrE5xa
siUsle6MpQ+VK3eRxTKpcYKEQaYachJbPq2YYGyqyHok3B2PCUBLzhxQkvF6
qscvUiK776AcgNiol+6jbtNAw0N5HNHwmLl4YXTfaxet8Ld3WXcF3ZcPyZtt
CuOiofO+pttgmJp9mawvpBZJktWIWh3Yx1PsGQVF0lkVXKOZV1RJSaBFHjqg
sJVxRNwIMn5n0AyGi8HA17BCmtsjVdzh+As+dJtc7ytVOqaX2qZfwFnbv4xF
fc6RY+Tu1f1+F1kbvglD8RC3e3pGXFnnxv+FG5HMyiHk1MRI27P4cE7fTIDw
JFRdQJc/cb2YoW/3v8vcYa8kuxrJoHtYf//4rJkf0P1u4ClyVlGlH0S4/Rcf
Sgj1pYws5lL9tyU8NUa+wbvzS+QYRwmTaEZGYUhOH4u4LO4a5H6GOvknlUGP
ubFVHOp2ulkBoXsoFdlfAc0nVUSj+DwlURC/H1OpjKlY9uDlKmYa5JfQYcAe
i9qT+noJKgtijkCnneB87IPPZXOUiNdVdXShZiauP4AOoiEa/GZtYptaBx4w
R4CH06tCSoHDIomgCLItAkC9FXFmVjiglpJ4AblSonC1aAzxH0vDkIyAVbjD
aJD8eJmK7VZU4iPa8mkJ6bpkHoRD3V35EPMgYdHgevx0pASNEMVdUEh6UuJh
qhuEExOpRC13DtIfXJnkcPi1aM86OfgiAv6g/jmjn2LWb620zjEFGdMWJIsJ
9JRcMBfGd6Oa3YjnnzHMWBAVlNAnB38zmxwzCjMckJo6AEBKRw6jFfrnQf4r
dJTxZHcCzGZ0NBzGJoMirgNcn8WHQ++qbLGp5jZ/VzpjJBITrzpWkjPWvaoG
pLZ5aZJ+gdcd04JAT3/OtdgH2gNOSfLE8y7Hze9HtssbcDU19+t7Iw5vQCvR
UNaRR5L2Z0j1DZKNH3jYrS7Z2Vgr5JV8CWfCyGXuZ9A6vb1jT0lliF6vDgFC
WcQbYOaRoKcmwIrvEXgNcIhJWHyHH0xZufrga+deG127DItCIXD4csmY/jF9
Fuq2UsMTUHarUYKy02WtqXYjDNOCGc8VtNitW9GDXhVlrKvCQeUIJk8MzF+W
L6d0lan3DG0xWfpsqZApq14mJpz5DPNOQ16kdtYDhPDIznfrinvwK5vZaXot
6NyLyVAH88TLWRXmz890lAyMq8uT8d1VKkLWh6Rm9k61nvqTvN9dFTp/w44b
jQ8adymJiMiHj2I2YC7PNLDLWrlllE2FOF99qwGTXUbyhSBdymFZRhG+TDUQ
ZL3fpecVh8ANxpApgXVHc47PPd5tiCWzGb96VdA7ANEhWTXdj5rzvqoAdu3I
D5q4JQl8qxA/i+nrm3VpHIloUFjKAolEk9kwbzSzzGOpkwEwEHJ7UhTbkate
mhUbm4y3ObMz83rDvEtt4gOjOYcU/nwxKvh+xEscKE32lE2cmC/o0V7aLvad
m+Rm4ggV6KVOtARCoPBOIaU9e505yUNHq5DFXzTDSuTBWjn+F/G/T4pfKIKN
4As1SXtiT++I6f+AlQAYXI/n+TByLsBns/fDU3H+KDuB919CzDuYjWrHXhjQ
BasVCxVVbIu1M4JVWNhUjk1EXbWqhhmrwl6CH5qRbaFtVJa0YhgPKf+j4BPA
tGtO9Tar/lKq/XKZkJa1HDsgDPdOPcWa7gY49tppAjSvnfLZ/8/xEnUI5D8F
8Ay60+H1rEKd608en30flpo/nnHh2tX7TnEWEqqRpSEvxdg6cdPY75Rg9NdH
wZ8j6lmH+wWny7zQmzajATcr8SVafnubCXixy9wvYEdIgqDTGAdd+YK8fkUD
jNAjiOU9o1oMfDoObD49qUdGE1JoiI8IB44N5y9XI8NpxHQoTGz8sGSVPHDf
YNdtxA9o/BNkBUkg6zTGz7Pkk46kf8MYNSTO4QK9J40wFOYPoXDVVZfokxM5
qwdIPxFBrmhpy5hDY0U1uaOhz015vvxUAZMSAHv6rkWTXp57oJoGQdQAULC5
INTZFvfSMCIY0eRrYR2B7Fx9QXsR0H7N7kfSYLGd61xPFFogG3DhoJoaexFq
HT7xuUATPFAwqCLrI93GiB2fWv4qL4AAmpE+e87TFdOy4jK5quYcoH0VRrUD
UJ+h1mrCODF/mgRNcSTDtyOseEOxjbysXhviW5aj3S92aWJMlGl9ln+WRr3q
Uq9HOw94QOpRQwlwrXLQgrCNO1ZgyHrenAasL1nGOKRizS/Y5sKbhdS5AJwj
O9FFdLdj0cVtYKXZVLQl5EppMDbQ10C18mYbhydbkcjOLnTCl81Zx1sgN9BV
M+pn8Bp20YySffwzDDopRMBprCAsmVJHF1Zs1nLhBrxbaFVM6Bf1xf9niw/t
Q/CWraATeM/giLNZsBrGTVXJBPS1wo9A7Guq0hYkjCjylbQFgrbObGzf9mkz
t3h68MO7qWwOt8sSjt+ewlyiTU0d7gZgp2lyy7UiIsZyza6uB2nfjv2MylFk
U5oP05bsIF1RMx2Fx940iwG/UwQkggd4/cFRPm2Pj4Hmom7Sd6iYwIJdXxz9
NQXKKxQF2VbFd1I2r72h3h2iHC+btjyT+kI1WAluxnryPgHe6FpkeUM3mEWR
N7N1mEboxJE0f8dS0Q9AJyDXtTYBF+YH6q6x9hlLqrxhNtO4U0mVysCbT/iH
jpDSG2vQ20FRaROHB3WtCN29eZIg47PqV3dH5+3w1mApbEismyHgwbvaCUuR
mfGJt9abOG318Fi0sEeIyM4u0zT9M66peT0X/HBUKywSSReYVyN10x+rwqUb
wHkMcb7x1JW6K50rLGQfDchVOPzSHGq4czlIu5htaQfl6vAL7t9uxeCB2ic8
zBSmiIz8ryZILvUK3t3KdPSObZo4A7+cwPUAM73HZ1+VRi+xTt+CBQOa8cex
kULsZ1E7kjxW5UrHeNc8DmS/luFDMK126oY1zefdwHcGHK277gNMkuQpY4ja
Q2/N4wAVyg0fnMDE1+LfDxINVbIHmngjg9YnxObW5dU+dmlpM3ajqzx5ro82
VcZb/Qhs9DRBq0WXWVDgz+CnhrXOmNJi5h3hz2N8fw+wbBppBj2bX6Qp5dEm
5VX8oPpfcUsVEUsGnD+8jmvGXlDkVx8v3jQnh3X6BWyPMQTxa0HDuzJ+7CAx
/ZQzMjNctoyK3RDtJ031HIyW6pHEsVTlh5GOVlJT0WVbbJ+/wj9ThkRPd2w9
QfF0P3qBEYcQBKy96j27DlTmwK2GsTIZYt1M8OeVeIeQ7c/wRh1zCsFsBD8X
sdox0lpTmSY7Qzo7MsDobT1ya/S7vky3UObTQrLcjQcR7Go9jsgGFibSupM6
qkrsI3OhBr6gVXbVusje0uyrr85mkDOHCFje+juf34Qif8BDKrcFHClB/GRn
fuCDNV4of1LhuIt3DfKPNxvePmJcCsB7z9UO7PfdapVY6/9XtDHei+kgyVG6
524uT0h9InBSUuIY+NJZ+jwi/7X+5rTIm7YWilUdJREJYBVbpRK/k7aoV3u/
uWRAva4I33Q3N76G+bUzA58BxCQEx8obYQV5MsA7i+O5HLXtiAUCzXaqkRxM
UZ0ll43L9WqmyZU31VnWiJ7KDJJX5yOY1JXJGlwnRHQ9dTzSvNmHkYq6nECJ
gOkuchQsFVM2GD+Hm/kvaLq62M4+qfuA0/bRLYF0ZwyFhA6NHKg/gNl9+ZFd
2IKvK1y0cMa+w+lQRgzrJkPb15iswLWMIPDC2nlLLZpvAMntCE9XFkBnaJ9C
AIZ7eUX9kCkojmz3Eeo6cSMdmIyrn+UYjjc7c0kPnqrgDRKOlSgMTp2UCQ/F
FePEoA0RZF6wmCjOaG0UdzZgCgmfw3FdNzahIFNR2O2hej6o2TF4U4E/MrHM
7OsbFe2jFJ65bLAwbqIbJ0Onus5KyQixcVl5o983g+etFgaFTsVh2SgQtqhF
I9fRYsbmyJU3CmAIP0zhpiJ6zoLEhR/OcbzyzDEgUrnXH/HZELhe/gMFRPIi
bOWkzYIHDs9AzSKblHlV0v33cFBSTN/lM0TOiDqfYI5QGiMCjkJcDvpb72kY
3mFlIe4TQPt0ngqvgFBCPioUPZe2UO1BRkqz9X2gVQVC6KmaBXYfS/a+kbnw
/Og5y4OCEdBeZ18gyA+6lhZLQOMVTyI9rueo2B8TK7DcgrNlttf/ZiPgKRAz
k3aL0E0/ImuBNY0QRyV+k0I3I1O9NuAgc/nEebyZ35AHp2D1TrTfEtNXxdrc
WsYCUfiwVliXhr7HXzL7YNpleEurVynDuy2asSVDCtd/la4WcqUIIhGnG5Qc
sM9STI3OB9o6n7lA8yeNjCAYD8TVTsYWFwkK9mrzOcv5wilp/ZuG9B46RW5s
1xIWw/uk322EZwCpGKPH8aMHavq5XWXRMHMuaW2MyM/WRl2YEF/YT/7+hEh6
SRYq3UP9Ez9q6xFm7TLcT1lIZthTmlgapl+A4ScgxlmBQ/S3IkHUSQkyr/Db
MZl1yPlclx/TK3F8QnDZZhszNJpEJcDVBAscCZLymqJU+Figevpvj/tgrrXF
wTs6w/n2nmL5sJdKEMEupSLVdhUa4TE0u8nbM62nPzUwZv1JEJe99ObDh+CM
tFGpmzz9FRWnl2jkRvgrP0NcsBgYAXf6h4keKUS/YuIxSWVg4M+1CrhTBtqT
1yOOF+JIAPjUbt4BOUkRHkw1sQ3c/3wvkNYtiDPvc8fN8GdYtm13dV6hgp+R
rnt54m7ZzExz6mCm8E/Q6EP+hxNFrYtfHh0sqpeD/vr5JHFALDydPLk/Hqp0
GBdDsluJOG6Ivs76ccwH0YxjiJb9xf3LyYWbdZqNAYvvbTFwBO9W0D9uylgY
9dqkZMVj+sFfk1ohLYQJR8wrPs6zIl6fbcCz2G7yg6IA0FHidm6JcphgAJ1Q
LizddnKEuy1MUAshxSyg7N6Jn2/5dGUuRuCmlKxy38aOtnxQSa8BDZDo7cxK
x2dpsT1D+TfvtGA1Fe8Oyn1McagdLZwi7EBzDPRGgNfuLZ6V4F+OazKK7ory
2ghN6zgNfbEq1WTeHUa7ri5ik8w1pgJfvbIah8+ORN4Z+8DuUGgL3MNNn/66
oeH1Pe+gesNjLfHCGoBUKfHHmZg70PQkTskaML0Eum/6n4PIJtFrlXW5I8g9
oPSe8OHFj/1rWYqBEJEUCwyiXD1XWYl++0nqecW4FbygtiltAMt+7NBE8LLr
/0jbWyLv/zugAdZUEpvXltn/Gj/3724sMOGWwhpxge5Iu3njogmwFRzHIHqF
sNhxvhFMIW2vnD6HsvWIOGHzH5ylXHVVR1JlGQNHjytCj2UL36OjQU4P9E05
TZhx0BemUVmb8WXhp7i4Zkzy8Cl3I2VMCvAqbHB076ac68aY1Rt703B8QzMI
db+C7gOmB7qGVkS2rfpM9Yq1AlZ2QRS1tlqKKY3RMFzvdlbVknKxlf+At305
OqOSQwK2MsczxXpN7Zu+DFv1e1P0ZZ74sdQhyxn1RSUMmdptAz8u+SpV30J0
Gs4XE9XMXlRLdJept+bqeCCGThT13IJen5/naK69aK6tcc8Oltq/92cupWCV
LQokq/tY/TC5IUK3hSXrob6TxnXe1l6ufVz2ktv9jn3SKNWpOcO1xC6FgDC3
VNtfxhowoWsuwAKdHKAJ/BXCxvhb/B6IPeiRI/HdLcjL3Lw+hLvey1I8jsNR
Xmqw//rFv6mMsTE9cVgqes9UCI8UliErxrfoGp+pj2NHXJnw3ljpCikJDOrv
t0TE09IDd2F1+kLYQ2981XE52/NflzQOhRX9W2MClluKYBzF+VpYIhu1omfP
ZXB/5tjTfUN3a50wRYH+OpTIXDN/HBr2D3/sJu2xjLdT2M8JvGxAXcXm9gCk
b6kbxodGitQ+aP7ouQBdBZ6nC3fCVkc9I2BH8qPlChB1XII/7O9XR7qN4nMm
2G+a0f2GFnU6lfEdpTaBitTJ4uaCMd9nA2CzcslZaJ8KeE6Fzz1mTZ1hmQt6
cQDYKhYUG9Dwb43lDWaHKHby+pTrgHt1ERGKweQGTMeIUpl05zTYrghk76vN
PmVkbbhVgpgkW3/OamwJgnO0evwAWubs4EluCHuDj/zFWr8yUHoRqp6+b5wY
KHECZUkjyPpX82s1zseYcJp7CBma0uljSyhTDN19PFPAYbTxucX6d21Bgpst
nQ+cUe7a1HU5HnyJ7DPzEVKKE7FctF3M/uRpa/qnPuGtmMGf7YWWlhOcRWYI
GMA79Ofb7b4J2+jMEl/9txyO3O0OYezU9SvIGS95bIEihgswms6SkPARxttU
gYWz1FdJIVtLzKcUF2AT713c1Mo3DPfjiqNruuYq1l5srnWxdLymg02tb8oZ
XePN9pdbqNN0GPXDmCaL6NfjZ+Ybr5jy+CHyufSgFuXdkqlCORb0dE6L/BzB
BXi0hptXqxV33AFW5LCf8rtKKMs84cuKmoqqk5p12bj2Wke6YQklUbP94xrg
KjZhTB7c7KP+5lJr0gB+nVq3/48xGlhBCXLP++Q6oCY63iV/kkzqalXFTpYf
DGpa/TZ2JTMe+7TQHkDskSQbrjxqWcA2vkZZK25VJE3ec7gI4bpzM9uVxrj8
MRjzm37DV9nB5doc/N0miunzt4SguB0wYr6iAsrEC4rEGymLZsFxrWHh7+ru
zxY2Q+X4CthNaz5NGV827q1SWXF39HYe/5kkS+nrgANqHhsSkBWwE1R8ynNB
O7kUBS+grAOQoKkgSwSkvIPbEm1OFul6/08i276n81ZW53/lwtM3vfK0I6sN
84I9obIymHQ/O45p3aRQVVIQW+BIdj9TfrAgJgEhum22O9xENNDev87pm9WL
qEU2z03Yn56KL1n+a/KBEfzCnzDQ9SfNWc8EDcyO4A27XbSwYyOxt036G7z2
nAY7HAPWD81SsO0NUer30Vkgh3iftwyF0OsC0ZnmNkW1L8CRc2wUCkT/nH3/
uyhAT3j7m6Wh1j3wTQDvLkODAUuIwhssj/mqViImMIzdKTPgSukScaUuO7Kw
BQGRqoMa/FOcettCoutXZyQmZdmPiSuB5kf740g9/YToderLmm9qHBam626C
bdzG2voDTgmJlcDF6MpaPFYOZfm+ZcD77bRk8yDaWIziz0d8F7H6SYvf9Wci
+7riR4If6siptQ4I6lwX6+jR8+R10InwlaV7Ipt7E5uhFf6Jv+e9nQwwb+Lv
BX4kpsCU5xcQv/3vuJPPIa0gcXWUXaeIAlGw47E/xeNwxQyU2Hy+7lLl4DsC
CGE7Z9E3fG4fFx/fzwpZJ/ylf8cLi1bfWzRcEp0WVHRofQnNWEqd2irWCco8
eNG3oydAA5OtmjiPGuBNmM7mri8Y7CK7q2pWwWXrkmbPVSX955OgTtaat1k5
JX74sswagTJ1wanGQk0Ii1y0oX54uImzqvESvwhXMltxhM/Ueo0yRTjSTOyU
ndsyPXQPMsyN4D796c8mgSS/EZNtFyKZaaQ/LNTfeUvTrr7xHzAFE+1UK0XJ
SkUo63CLtwt75a/5NbVx8i6oxvCgtvxsHXKjzwHycwIIgaiyyV4dzLE7wd4w
KXQlAERy/TK5yqIsi3HPD4n7W4Dt3bb9HppzgYwnYsS952CLKjNB51pB6mm9
mw27BHVPMBGMlXWzgybHfrhvUsJiDrg3sVsQM16vHFKC3maSwIYctPNmrAl4
MGzchjX9KIxR1Zpvu35MCs2bYF31TyswQITCD7AvfNJaAk5PIGfGH4hE///Z
Kvmr2Hu+1ROxVyf0sezbLxHqepcYjgq3W7SrlfNTKVtmx/BZamWLlBitXGQT
PQKXCoammhevmSlfnkWy/2uEi98TNkMd5oYgzbShwcBhMgHckyIOPdBuzJuR
wHkerENeeiHYXtmuszDIqZNgOm6oKMe8NaqSm3/tnjicoNHTkXDE1xQfH9zI
cqCIKKW1UAjh3+nFFsW1RS7Y96PSJqVXJeiI/wf5ZoEj0PJjbvUg1fZe5p1k
g0pvIRy3XfnIPgPl+FTz109hTeTOTTlYm2qYSft8cg/zxLEnbvgkTSlQiQud
OMkQqY7gkN3KT2tiYZg/MS8Fc7D9WjMilc1LYBuznfy4sn2K0awTmqlgX6Eo
PdEvznkZ9IJy5r7EJNBCoLMj0ZsCjwkmCxYFAg5PvwUBQXWQumSP1UtFRq+X
H/WDFySa5MLi+bZ9HaDgWsE8gppxGg2tRfUSdBgNUoz85wVrWzjUXu+DUy9C
8iT71lT8+1Ys/utFRioihU/JasVv+XisATdTQ3EqzdgJNMESro4dnoFg1mO1
2yWdKF1TOc7GJRgpKOZGYU3g+9U0xF0goTS+Rui79T/Y3L+qUzGWCvrT+LPC
z+6SGn+qU2fDvT/+lTRoXb3zOUF4IPkJH6Ui6enw4K2uEGovThkc0vgUDQIv
yUj4KFTPQ2YYYouAD+iOMshANYj/K1l6RAE6HcLzv3D18GHorKHCzu5a59iw
TmQwtfYMYCtdaekCJncC9KQ4CldUQIoc41LQE+CdeaVIzB/40D58pH279q9l
dm94TgUCgMmisdG1c0Z1T7gt6FoyX2CRZY5AlTMqAcpEZvmJJI/JLe802Z70
xxG9MH5zN7Y2cgaXo45ILk7GFc4Ty2KMnzv6QTIG7geb30n4/weiD3eNnCNB
c5PqJ3VwDPCyq+l8RG+HDobzhlLIs2dp4kwHNW5rZL/nWC7L8WtBOOxjJKy/
56GBTyL2Sdsy5NylDDwPAhB+wLisQ6Xg+eOMYA8XksIOpTktCA5k8BGbrEsZ
7iMvJny3s205Jch1/0TltoT5TA26fwCxWqRbFjnK12bu5yyxM0cu8mMQaIbd
qzKQBbdigEtfxB2osp4ldoxlElgzLo+VnPhffmAmUF1BI2uIuGMprDXRM9OM
Lw17ER6DrRUZNX7hTEcQ/RSK9UDqptiVFphLhDo2dtNuYYOgPAWN+P/hcg4v
mXQAavhEvk7ksmHPCdRxqD29M39wipegM0PToshohSzIa7GTjV4UONag88ox
IH9DE0v2HHckwS0cRGGatO64MRTftEMdSZDLFfHPc3yrlVXz6qufL42Yvkrf
jIbvJ1Cw9MRGTSwJzUoqp3sOK3BAk7cJDtTRUkv/zaweSP61NgHZa7lKyhl5
1rRpcK8vMgc7Ig+k/qWsBgQjhQu0azcKVRDXTdPUaZhNqYSi8pB+TLl/nFP6
FIWFYb6hR6wXETzD1wWFAAGubS+muLbat6PGLywylMWDKzDneD4J7jrzlGlK
5YY9yu2WdfKadUg+Ou0dS2HWwv1ql293aId7FN94iOSn+wvdDiakn7lCiPb1
gqmV1w7o4rh4CxinpF/hDrmXtFeFwVfsTBrDiTwjATGyk3+g9jFBI0/EZY2w
LJ822lr+woZm3zbOWw1QP9OxWGIwtR8qH1Gsx3ewq9TgCq+d4Y34qJi5OLfn
YgLg2k59zuVTUyJvg2bsxhfnNe5oJDo/7yvoPxBKVd8QelqzzBVkdYeIND3C
AJ9sxu4d8HwDvfs4V5B1Fkxv9UtPUF8yKgpeYNO8snScU5rGNM3Xf4tJbJv3
pAZAsshmKNyaKgrTrw/UBDcoPzGOKVkQFIvq1uhFLBY9rATV9VGJ7MVCK4/3
zfwF/IgXje78Cv5TRQ9pd24y2TAszHbgO8IGHBTbpC29Wm1HdQsxzwpqaPHM
+/hsKdO9lfCaMnf/du++TmI99fAnFqXrfK+oTHRe8+YHjwd2Q0JZgr99RT+3
t7l5KNRrYpR+X6imIJKhZzTwcJ2LAj0vQVjZR64QTWecoGwq/X7EVd44JqTh
Ou3kMpZ6XSdbEG9Y8izVPfvgSS1JzPavOwkoVI78nZ0oUaQJLJEPGbRhc73s
OOmnyHkIyRO26pcPXAeVKpUyiGSoIA93DScdcg0vB+IkIZaSalpbUfQje6CZ
dKkAGGnwUxgVGCD2WTbyhRiOgh1fArepd4QSw+SIKl/zggMDvbARjp9DBSqp
eVqSnaxOf5zQrpYvS1ytiz2RCj39z+mACRSAH6UkFyeUsJwZoRnHEPEbWrEO
8gKMyooypL4BSH37fAjKaI7PbhD8LALo0Bk7O4N3//YoX67zSBUWsxeskQOg
urxVRNSMFhlsW/l/kByODZw48At9EfHey6SiKK9PbGqyRebAYtX3SxWJBiQC
abp3jyp9QmX+fF1CDBxdgDVKBCv5CnfbiUYBTDcxqDOJDHMv2z9Zzoom4rLC
bDhMDopu/xNxXUbwmEdIWxccMhq00+lKkD5E/2LQWPPM5DL87yeGx+S0Hooq
0f90N01rNyV762rldeFLH+2b6A+vvIhU5LQhRLGkdXFFgaSdWoUuyL5XpWZ0
Nj+IvBVK7VHlG5i1wuB6hA/wa4WkGI7yhYggvhZ2gZIFBIeZc2E90W5wP/Wc
pr92Gw6cmhA6renapQFhT7YVvWDtR8RQ60V4R4proSC9obE0kBtOpZaNhnDn
MSoH22qb87QfDdjbWcpk1MUUKBvG5g3O8K63/QYd5OBuQ7G4wFXpN5oyitlU
PRB/TtaClvNRRSW32FkHJF3uduqHcAY8puA8RAk7yPWblNWRaCYEwK9x5ayo
ioSRU0oIIl8JJ7tP98I1aX0L/3rzHWul4cC06w21U/t9Ldj8kVnNzM1YyZR6
C/vRktEwqqAxHFLEmt0YMV+OakZ3i5etQlrnCFats79RLpdeD8k+e+2CUX3b
6X65u8uONtjc38ry7b4FCwFrB6APJFeBwpmCYi1YX9OYuBc1Z0HQZND+CRXu
gV7KUys9Rc0XJBwJ1rWbRXeWsrYVKSDxMNrHKYQ8UZefC2epwFY9pFVtI11N
6ZixqwDHpvC2CKb0uMKw9azKM2/vxnskPsU1B4+MFOKpAhPuwhLN4P4sIdn8
5SZw25gFpsy4s5wv1xulDPROdO+qPO96nO2OgP3e8Rto5CGEedHLZkDpjMXA
KwHSheMquMKc3ORb4ocXIh1M+r9Wv0j8eFdub2qRb6Gkh8qDDsf2sDHyWA2m
xrdTMNmPFfCucf7TQ3UnqFmjeG3B2oG2qbjkL90QJXklWk9GUCEe8n/3XzeC
ySCkqcWKD/+1h/HZyvH3GtcEhWV5BqSX3ShfAxdK19vI2voaQvrT+TVjvB2l
ZUnRUy4NulzPMpGv2cr4EzqyZ065qRYrBvwegWm28nMAMWxG2/L0tqONV539
Gmd6rehOWx+Cy9fakS852tRXKvSafg6qGpahF6XENlSBgF+ciST3s8kBYKey
exNZSRM7onhZtgbBEZ0HfMolpNm6qOw0DFqv/5cScG0UErFTPFO2xUPAnXUb
zEQXi5tqtJtheTFnaDRfE12jxtRUm6DnxV9rljlTvINEyjTB7ZQ/F1DOQtbF
l/qb+s+uLEFV6UO7oX+mWyRIFiSK3AaIyDEpVrp5XomInzSV7yNIgFqoqLQl
I9Z6O3Y2c/nFbRxp9zctFeJG1mO8yPX9Gky5lj2L5pBHxFjSxb++NHPsXcRY
4vV2YyTzULr6qpKuKpO5C6ZPi6vIsU4XIEcfW82H/aBkbHlz7Xyfi74Luo0+
tqJJ5EuMx/F1SBRMWBwK9ngHp7TyXCqwvOSecLVEHvq3v1OumCBhi1BqnQeD
4TCmDZQgIvjNDkaagi8CeKX+6zVn5IMpe+KZjF+ZXBEWU1cyt4QnlpoCn8n4
SC2ZZKVpiKCCKjUzIDyHsVKXA8zsYhxEIzFEMmWFH67w/zxIcbEkr+ApCYWZ
jo1Ck3mOy9CHc+8QHbVhO9bNrrgQRLCIOLd9RYGkOUfUvJ6F003HzxI68+x9
9t0xaiV+4aAhgas8HmKTQO1B7YXFTbiMenoMpCWn8BtEikzrnMn9+Nyrg3Uf
AsY1Ha8XMEnXl59po/f4i27K3KLc5PndD+iRthpDYbzHHVjxnPH+MS92QxCX
MGdc1hmyg8ertRvu0S7WqTNtdqGO0LQpq6awhixzCZ8BA5Poef9/adO0kweU
GhudBCM0eV6Nyf8R6Xiu5IFNjMWXXc8BAtdbpFj0u/ThuigXF5kNyfZCsOZX
Jal3heEEReaFvZ+n7FCLZrfQT+mOn24KX0e4nGftXRsNlx4CLUG9U9GTTUjd
eNzuQeCjXzL71n2jdoLZluFWNsPlEGVjmV99OOG1RNCwSbFAvjxsczesfMk1
oCeWjenwkbWDypVz9xbuTwlbo4OS/PiYrcQbjwhdSPH8uLPG2E1KwuY3dhde
FfA8sijDgoT9Qw3zsAW41c7QOr3RRqWxmwxoW0Z+wD6mM5m/Krk0JqJoUhXR
i/cR4VmCZJ08vdwjIXblrjQ6x0dQCLWnac8WAnmoLoc8ewGW51RR+RpZZuiX
YFj4kZOZIV2WKpH5vX2jO7mdYiFEm2Ty2YzwMicJELd05aWlcO5Ue0Rjtkrb
OIjSgqHYHqKqDeYgiPtObbUOwUiifgU/v5czz55JGF1JRYLmXIpBczBZ7t+s
hAnm501PR1trRvCM5jEi05b/Ncvb429g7BXro5bnNU2SgPRA9j3zMeEsu3gX
xEvvp6oqRumvtXLYROFyIVa7DuaEeQntQ5yzz51uM9Rg9gfOWDfQC267Ynsw
lyWPcbs8vOpS4aOvdMiyx53y+7A1DQ/uv8Uy6yolJB8znhv+2jzYj3xEY6bm
/Td7ldfdOTrB2Y0ODTgd0t2Qqcj4IZxX6JynNNrJzF9pk015lbO4fvKJBgoC
hwUS5V4cipLSIVfjcLUbtb3q1uY3ZxFlp0YfLUG82Tn8NEOB5zZ2WEETVU03
3hcaz46rIxDA1YxmMcbvZ/tAVOhdJcBehBVlSy4GD9KT867mFy5sArAc0iRd
m4gVPWx9PbVB488M+wkEITAAvvHUKlRCrz+C1zZh7x/6Vw2iLBbT30EKs/nh
9DLXSqDfa3MzHqUyXL5ohFbt/U4MN1KDu97SDBp/0e8DspiXBgOfLX7bndNF
4au3HuYlXkuJlaLd0ZeI6VmijjbmawjovFx34KdEg5AK+zLyI1srYINK0tJY
NAgmI8aW4yLNS2kO583uZO2nblfCTEeMtYGbmYIkoWHp2oqUYPi7kpnT/YRp
Qv0+VLXciWqmnYLFYkNGH5ftJ0lt/1OgfwRxTUJycJopUaZD+Po10V/DWzOQ
isA1J+Kbza2vVP3pSo25IhBVPJUNUVQ0s1TVmreO+yBDWN76YZ8R0goWmh97
CRh7/blzBE3hOi6a7TeCK/f5+4wvG+WnHb022gDvvc36iFukpTVECJqglV+0
BMUoBLINsDtIOKIp9ivGhwhDyPnm7HxDK+F5E3gatxryBGaVn+JGJ/mQNRn9
FXP6PkSG9jqf1ONnxqTO0dN+Y6OPwXG0Xl3y1NmwXUO+q9M9mwK6PlL8/PKX
eq90xzkjSbjOzhrAIF7bkriLKSmo3MODhHnxTGqKxNaAbjVIAueL4kk9lazw
uoOPYn73r0wh+2+M365cLh4MvqA3Ab+5vwLLHKNMw84gfGdlQGJOzY/WMyhy
Ae7JFTrRGIHW6MdyPmlXWXirCh257+a7AXwPvBS7/GReaAzoPZWuC4SMB3x0
aEw4wyq/3O+84vmfZMvFWgjYQW05F65bdJR3PQ680cO9KrXDv+SVQYIWwJow
PpKiTgbxymOKGsawNBw/UlxFK/Tq7tKqEffMnnWr13sc1fVNhBkVyslr7bDD
Mg+roc0rDHimPQvs/evZR9VfyB5v4zgWuXnZ7saxL+BdPSQPaLq3ELQKL6Tl
MzhG9UsSJvUSunAJTM949VewwbsopP0k/vQH7INCddgayafM8ZxMb162GaCC
5haQY+PlChaHOF//Z9/xkP+WLBy8ewhpaNGSAfX1Cnx8F84uYuKDiUTNu942
jX+QQaEJz5YftbLuJ8PvhCyxHxudiZIRmEiHjoYFguRhopIoB7xResUBHC+W
BlVft9E/czWgrTADZV2Bt9gyKrd6PG2wKjy4J4nXefXT2CkB8kcvd4NWAEri
Knsmw93tBysnTnW4eISwI2aMmTJv87CvEsOOafy6MSPZZ/1m77XJgwzIjp5g
+QZpTOUK1CqLCGQrQlBh2xbZPfvEe0NIy0v7KQ/ZKCCSMVSPzF3311DQUUOk
tW4/+QR3C5Z1MaHNtS9baMmWcG3S+KHwILLEf0gQlD/C5ZX/pKHuzYw9pXAU
s1mFZi+ekJ+OxSv+TtvqVu/7i/9KEPI8Dka71hf/mAmbXlD3i3mmVWYl0/Cp
K4PjKyey2JiEEo5ygmGiwNB239ZE7OP3Vo/oGzeFzCjrEdnLvPutaFjTXcYX
BipTCavXRwGGFwlAAfT0vJ361DqOd0Pe0OgS0x7HyPTAZQKG8yfyKqpbElem
vAuzpadBCLYNcfZARgwJUki+h0QCf9yQaCsyGobo6zoGFWlJ3jVzoCh/zXVT
qZ7Mx+gw5nz3bv2S5/QTAO7KsI7DSI7B3KfaISyN4dixRNlSkgTSiSfE/5zX
aSj/HVm7U5QMsKGczL8Qo3quRGbEw+XHfhkMwvw+e8nt0SOfNHdqCjiQuFxZ
fbz5gLFARJ9me35CUl+6pZvL+fGv9ZoAZ1NJKzk/SMy7+vvXECpWJ32ewcQP
5S2o4aoCt628uCcTrq0/N1eokh617uaVNLSYqTcdm3AMqL/EK4H2RDhPQaua
iMpIH5NFf6UZCKr38HpZrFpaX9tyiw/LEfYv3JShKaQPNOHcZVcmU0FBh1Gc
0ZeH9CRVWtMyssk83eF4zxkPhHbqfFR6Db12zCFSYEtc0MbKFRxm3CG+JrgV
wFfKVmHASo6TmV3sU6wqPBW95gHtny+GS6955LX7Cmr/gshDsCMLxf33zKF7
Th1sAtHPRoz372Fh+umMcfnNUHdjElBZShNq72J3/mqXNFlDAKtNDc5KcDRb
pxjyu0RSW5YdiyXZAPUVsysROtT28fmA31QDsMBVgh+sykDoYx/qnDqwiSAe
q2F5hzznsxeX+gR6QQ4QrNBmAy4fS7wogOBjLcUxuTkl69eW/W3GVxcdHU+o
4gH4Ger8Qg6Mi3/rEQDP0JEBilIl0q/7zZS8PTXujEBxi+5CvkZxNm8RxE6J
Rw7kAc8/OyeN1Jljnjyf+M4dRUCby5i8gAYaj2N8R3+A1MPB2NLpfvJh7AHq
HQW1zWkHm7u+4B2tQEbcLAmLiNaBm6KAZFYzyNWOY0+wtLlifxe1n37NRH7M
lxOJfkC2zk402qmWORMTBxSyzbo/CeieDM2SpQ5KVIri57C+ePhPUWziV4+D
6GzMKr10ryn9vbS8Ym77TvdVVeHCTJQAUbo8sZfsGW6tGz9ov6cVqPB2/npb
4tytMKJv8MAJxs/ppFQSqjS7il10Pp1MCj1iygYurRXZgUnCVikV2Dn890AO
dyQ39gjejiVdm9kxVExTQE8u9COArb7wq9iLXlBPPJWL2axePHoxQcsyy9by
xZrspNvfzlAWv34AVSc7/tmmFJ9K2Yz2OJLRz3HlwUYb4K/p4qSk2iZmZd+A
NwYUqd2LCRoNHDwbij0DtZoBflN44u8nNYPC8rGmR8ETRcAZ+r3pi97qgSlA
eWn+rFVPXJrDmNt5TDQ1H2tE+hU+b+uaGTp09hSp43kkjCePvaiJUUxOvj3Q
XIlSGQub6YuySKMn8fr06QJktHIifp5Jkv1sRKEPj30kWmheBUsHcu6SXAQq
xS52kakCIagtkWolc4y2rxroAgQ5sJnC0JizaEP1aTVMWsp7cDoj3lD2Jat3
BZKRBHNDz98te6RS1d6lPt+w9++xtUBLQI/4+4KTvj8khyNrQB8d0rE08xCU
9JPIpb7+IvFp+6ee7MKiICfZ3Ek/1eEO3QzaRaiqjcbWOkFyB4yhD9kd+ygx
zehC1OYPNXaU7fuJyDhsyqCxp4ap4tA0pauLpB5vTGhtiuGYYEbQZDaxlvI/
zCQfTCnjQysBY+TMJcgxIBcZtG87NKNlbn1euP/XEcc3TvDBc02ySYD3a7O2
zq+b8eDIRH8mPfCJZDlbfNp6pIzdJDKhcCKxjvdiW7yDvy+WLkLlusFUuzio
jk0UN88QqT4tbruXI2tjZujAIX3jcnZABFu7CmMhlpnQczkjqb0P89kGZEbL
BESYuow8I/pWYx+BeJAYjTKMA7liLnfqVir7JmLr45WK4UWU+PVN0eH9g3n+
H3jh4j359JdBbaJISxIVgLmkjmtvdq70L4cMzqGvo4m/dwpnoYoyttYyCUE8
ewwb+2NEscGuBVMzIDWphFEKrzU4HkdVvvXs/6sO4pWhbsfhsOiljzOM063D
ZIDFgBN9S+S5mgbEsqWbGI2I8mi4aF1dW/18q149zCRkHQJ1MHk3vzQh9pfg
yLFfWOn/azvHq6hkY/Y2+IJ/4Y7Jehjz9gQHE3kkvLiWeB7uMBWb+j3buI2B
nQRDrllINL0ofDczQcSk6K6bLEWP23MnobrXyJWdKUytAhEzBEkW969rhkQs
pqpgSYzUnT+A2pg3tPAcl6CJbk2cqw+hMMCoSBEn/4VieXd75fSQNKnftEdK
qnzaWwHcr4dbmlJJ7TCtTIcJvgwHXINz9rgAZM4GXXkgzDoyGEYpcVZ1GCHL
5P8eVWbOT3TZRrfoFNyADqs7ClUcLwmCN0Ym57sIvwDg+DQ3+dW6Udpcrx/K
a71/IV3VQTV5LA9bs+Ot6TTpz6ZcgWVNufZgeUuCrURuW2mI74IYHz9QEfuW
uIy8wKaCfKkOlJ3lIr0wWw6ho1e1ARgLD7HLOv4WL2XTiGSw67rV9euyx399
S5Zd4X5UPbH2H6uEZvKniJX6/wk0ah6sgTXHB6GYWPqFkWrFAB3JgoHmrUEX
y6ZFPfK0Gc47vNHdAAPQdfXFWn1JWYsZCAJmtUH+z039CUSsPkZCZWizuecQ
l9JncQuryvGdueRyJWt8s9Uvg/JLBYzX9zK/9rAfVNJOJijGrst6W2Qy0TD6
GFQXkRXzgfA/udZdhFoXz9LXJvSw7dROcbrLjlEbsTDshqCMDCea9mqv1+Gc
R2DKN30YU2uUxnQz1ZNUFZmIhloHg4mWx1ZgJWOHu3jOx5rJtNdWoeHflhd6
KEHDm8Wt6mpsdbxO181ykA5JQG3Jsz3VfLg8gM5wORIkVLveXOFZoQVo8+iv
D6jvfBheZtmQEF4cUHwme2yjkee3ZVQetK/S9GowmED/O+fSVspWgMUviR1P
9EXfh4KOHsolOTQzpvBoVdULAELF7lTly+3/pdss2NEE4f+yvLHZ7TxuOMaZ
2q5GXxQlgqAv8I8oUsDDaEt+EcUPTVaLaxUp9sQAcGViaAAsp6b7+M7xu8SV
nfTqe9beh3+mwzGBwB4qDJpS2sw+sV7izY3FFetPsh6cazvZh8/Gd7yCz8jt
A+EElK/YfC1fSwUj8D6SPb7Rb+djHBwWERZKmm2RfMQ4dNe7za7VuU3LpNSa
9gsobfRWELWTWw+wOe9QCQAS6s7XDRH2Tc7CbkTEjax0V7asPMbPosjji8pm
GBA3n4vwAIbInyDOl+yZJbP/Mm0OkPWd27Z//TGzp0Y5gQK0YgjlRXhYeLTv
3mXuo0HJ42pF9M16ju8ZVP3xTgpxLi4gXNzKVRZ2uWAvcpk4JaREJfTdsLe1
Jlz7xfpxoOcxTXEUdU6vu9aCLZ6bot22HlvF1Oz/30vj2CGOxi/vCJizyW/t
GLJWxy50ahUElscbNU5jm6sYIvNVvZ0G7bXq/NMT+TWVcAUrc6H1Cp8e7fQC
MgtGKn6eHSXmusH1+l2jLiPJnFffRSowJnF2OgJgZOWc1YylN+z8eizFAYj1
yz5XWml8fUp1bzXqBfB22ZWr0IHzGH7p8ww2EmilzWyusm3DAVJZMqAPkcN6
A7/v/PRvfnFSuyVu0Cu7rlBRYcHtTuJReMkN1hEP5oOiaorJjpasWM1tX8B2
RHEQTOnmYTJwrfh1tJ1tGoIKmZkqUkJHyIdlxOntuV51DBNSoigFS+dGTZXU
H6yY9aZ/1zRxJRu6YoexgrfeK69NjrSeXTZMKBZ/XDlvILFyAzRZn8ucgRS/
CI0UlsrWmW3lVja/rsOIhFCe6M//iUvwuXtn7vEB06O4Oia6OSLnEZtUcolv
kcyluJfDuW4191R1dy8VG9BM56oaL620DxssrkeHgmuLa+G8D7Fbhp85SGps
RwitXqgtp1InaxUwTmutKt/Z/EKeMYCi4WezxXenJNruiWb6RDEoCyze4nxX
t+26SOK3so64JcklQpoBNvgYiH0sXH0qtcVvpvfNDIPHi4BkN0pm7AHm5ZZj
LXX2kjyr8DDlzKYLEXRp7OmV1aLy3JRTlJF7A5i93bu8xYIZV/BrdhYjl8Zo
shFNVOIBlB6RA3soZOt0RcAbhD93nLpQ+sI6GrW0aZdmNJ5gMSYhW2aK4W6D
l1Oa2kc2osixJOrLFr1hatQy6spUIGRxOXdXhJ9mTRA8Sn7H3U4VWjVoGErw
9zT+1HGD4qE4CZLfHBhhO36CvMbkQrYvEJ2fndp3xbw0DYE+dXGO/5oz6Oc1
u0AsnX6TlIoIPBxH1GkzuV2BSok84RhM2FUJ31m5AYceTWjXyGjkolATjrsc
UkABp1jzLDakzGQB/kzvRTaAboH3JSfVFJATxFVza33GI3zrbaMXwkTg+G2f
ItOQapeRffVHpD3tRZ8CyPOpesbrbJbhj4DZNghcqniyHHTua5SA5w+XMHae
6Rqu6fIxzI2Dez7+q6/RnQsPu1KdtS4B7UJyMtsRtxTSSJHmyGYCL02voe0R
3aqwSnmxa2pVLBxS0IXi3nT1lY04I9WchBaFjCyHvym4WUURzJ3jJfyFwt9V
rM8DIDoYMDJohCbUlykC6nhjhq30VLl5U7lRiKeWyF8fyGYilYYXhYVbPTA+
K2g2sJcbM9x9pmacRBp45UOaTrf592WMMhdzrW0dFhpalTPDsj2x2FpKLrd7
YoCQlNS6BSEXXXnjEmwL2RtVOwefF0eLJ9asHl0BsGMr/LvppZ9j8OSn5aJh
+vXs3NVbZ2rFCFcVFBjWBj90wK70cSeHf2txaHKJs7xObrvlXh6+Fz5dXsiz
lj/DUF4RrOwLmyqoyCP55HWaZWIdIWTrHBdoyyE1IqihkbOSZU43mRV8qHsl
jbB+o/BRt659mvka4Ca1I5tvjPh1cydM84IjeTzG6+XKbY8vZUpza50LYLPy
Je3rq4EUY+CCoLaMoKKHXdHKCDAvLv8T1EnrIul2PCRAxPjmDhrcygxhiixY
X05rZ7z3mvPdoXLfOgAQNVW+Mvz9eqK+EsdzhJj709V0+oDp6rUcbkeW8lN1
kytZARJ0ipiPC+r4dnvHCUATE37npzlVSFWh3Ag/Dqw/9150FNYkGp1Hllti
gG1usEGrhh51+AwUpGMVEDDvDPm8m1RqPUxzufwXBMriyQfOvkZnPogONvy1
d2RZV03Ex5QGRmFTudJ+10ZYoQ8QMRr32F2G5kxRHb96P0E3ihFrcKB50YAE
TAaOpmBvBoRLTr2qG9034myYyV4tGUA6KM66ZJgct9AcWYcFCwlMXGXAG4NQ
fx0vVySY3C0/fJkUFLkKNBVIQyl2ORjTfzlS9pXxmQGtkIy6CLFyBaZsiOdt
I4NeZP7LYw/NbZnl9aoUZKRvCD3FA72OhPmKF62P8TggmtyNA08XiUfp9GFH
YcSEIj2zjP7XvW6cRdX48D6+3PMYNo/sI48HkHLJgDYw/B0BJAP0qe7PxPop
3K0EWS4Ny8XxhAF/zv2G5R5KGfjBrGa3zBhpTspBKFIJtQnyLhqqPY54lS7W
mwq0P1T6r9EQN2l1Qc4gfrTPpAnD2mwwNNBtSwHVwfZVRMrbZQmP7fiBOqws
/pjUhdRbQZW90ueKBQA2/pY4dd6ULnBUEPwBSFg2odPTeiNKHdDYXPLJeOwL
Rbl7jRB/bzjiiOiGc3RrN/Yj4Gw3BkI1xAQ3FSNwUYSKjV0nfwf9CuwuSsza
OQ0KxaH1QGnTFirskmx8ltTfFVSLmDDIpq2n9pYN4A19csdWMokw/GFEjWm3
vAiDJS7IaEbsTts1BoS/B5WnfDLV6Acb9Lfa7/pi4n8uzVUAtSoCqMBm5Jaj
FWVcPOcGlljakl9JHB/CHcvUANERZ0x07U2sfiLoJ35Q6DYrA/6q97KGLe9s
58NBDqcFga6YTGdtxhGdaw61z4GqSmnxBn7t9lmg6uLyAvvftgArMOP56fmP
qs+0emVAkmqy0/NG7KAmyIoxEJpM1QgN2s+b04zrkWXio1WuPRINFubZJqay
K5LgA9RgiPzh3yS72UjyttzW4ZF2LkOxX8RzxlvfAzc6p8A78m5388olyZT5
eQOLgAgjEWQ/FyhXQnII91YRyO6GWLc8s6pWIklxaq5llXhP6cbRTAJyWcUb
y2oVl3gH1EKs3GxEPHTZiwxSnyeKnrhsXCAw/LSjkzn2ymkFUi+x2W9Jl1N9
44VpBU/Dm0LOMnuaBg27f2ibb0Fm32s7RWxakujv3ByHeUOltK5LJ/BUIpUl
6/NuEL9vE2CzFlObeB/rzD3vRU9myzzSFhz1PkrqW4ISfERxZSZ+8U1TAP0T
uUkibUdvcmmf3iDeYwMFONq2MI+3SEGzrxeYGqVRrg8i9GH54RHmJ+ZMQtYo
WR3ABIwNbSTOrFvJ6T0Y8N3GhjXIKTOqLvVmzzHKrodKyUgVmuenU2O1C4Cf
1+yo7SWJE4SyiUO+D7FjMMlZUN4fg1VFL7o0xRCn6um/HWO52fj2hg5wLKew
51FXvlEWEvd/oKM7CpvhJtoAAsK8qk6uuyyLZ7QsIqzeWVdQ6j38MM53oxAE
NYUGSGnulnBmxZn6HfJBG9hkIonfPolPq2qB37l6sqEnlMPbvBQrFjpIeL2q
zFccCyDlJyKmo7mXufEF4Q9blC9a7SwDDBaOHk3h1HFMIoXqFgAmbyj2t7Qu
y7fgOOIXHj38yptIKYWkW2cCeUSdK9851lLL8+cEJTxRdsvdR94yogbKVbjL
fpnQd8BRNdvC3dPEfaal3nq5CcMWihYkfrAeiRvxpzDdF6alyeShscbYlQTV
4acWkPvChxldGQR2OmBlq1Fmp0N3lKfemcawSNxOI8/RLvCh0GxTqJ9LDezr
89c7NBM5qi5a4U1kkRVcYtqzVc5BM6LV81p3CA5DtXbngSktvKmvYNpEEiQH
okeMSibG1P0iazZv+1pYJ2e8G9bbRn0vMYmoANifY3PxBanp8Q3Lxjj4dHJY
cQyzK+NU6lhAJez37oUE7QBUXRYh3JvcnAv2KtBLX8Xrmmd+Nsm2LfE/6YTQ
liYjuNJsgZB0tYh7ve7Qt+utzOnDW7g0oSIc+MwkwvlFLtEQ5zLRZJer4lNY
LtkKhOwP05kUjuOzZRpsjyMbRIBWp0qh8v+V4VtWt2DYQuCCVwByByxj/74T
VhaBFHuCcTHYbBuhyU56vsRTWFw7LsWFOKXIPQKSEL5rhCS/30AI4WM0Imx0
UnDqsgSpAQsQTAKNyOUG9r2fXPQ0FEjfA9c/okkoHp1o0rlOXhknp6sH60ki
ABYsj/bzAwUoDVJXyYdGfMKcWLcbvCOXIdxTQT3LMM8Zu6fBJ2hRRpUzJGRJ
3ltFao7zb3ClH02uOU8Src2bIi8RpsT5bDVNQz42b2YtE1wSRaaZ+b3AIWha
JQqv7EMJTdbhJ5h1H5I5wepAf+fQrLWyEg5HjDNHf6QZCtlV+eOKD0xbwZyS
dWf0IN/Z4jEbsNfbwcsDekoS40emk9qkpn0AGPVok7VzXRlp/nxxHnz08/MZ
ZMxC0NjM0J+NBDDoELhb9pnu1vITZmDCZZnzw9EYN2uJflzwvmAtCjSCMqCX
0iVtOaqTnONl9xTcWDrfkE37xpjHQU+A6Pg2dTtEbgkPZ6Yt6LI7Of1HMeSq
uoawxi/ZuUYWYrlvFtEPUOgh5q85qQFJE3XiYjL7SBiK1b9APvR5HjK/0HBO
obL0h45g9O2vVMBFBdDbm7m+0N/E6KbTzkQeEiTTWuhc93vLK8D88Ebj8p+I
S7wxOZp/fJs9TQonXcKzaCC9Rxj3FzKjSvSLpYKEd4rH8OgKyZqEgnv6ZEI6
dFKSZwrZ0B3M6EGExfb+5gFUO0Q+BseiIoR8E7cQN2OIm8en4Jm+0nnYRXRT
rCe21YBlXXzsr1727ZSEfXACbZyHbPka0+pgzcvQZ90pOMClA8sPaGaHL8Cn
IKIZ6ktLwvm1n5Tu6ouJ6Nx6UOCJxM4xkUwQdVe+qQiLjUYG5eSsleD1iy/L
tn3ZOsCjZD43Cwi/5e41rgI/sf9y6mcquEBJaJbxIO3CPdtvz7ie8PbwBDhY
8Txw8UdkuVYP1mA7YEW9M77Kyj5zeE59kucC57PptmlIJhPMEHvk/NbN4sTP
DdgV6sHywA+JcG/ZBocC/0ajrvuLUKOzXnKLUq+L0CTCQ8C1nTarRlo5CsFO
Nn7ijOm510xWWtHr9hEXwSs8K6K5RjbYB3UbG+LkIrzsOHY6xUKnrI+Male1
2+7wrs9tZmlOcLzedhBb/QNe+AIZ59E8URUrVN1vSIQ5GkBKuFBuhYoUm7ro
X6Y/YdYM3grH74vNSO9lUKoZwv4d5SERCek18FIFuAtsjrU9u12F5C5OhzqI
oLmiSrZcadGq/oIjY7ZJgWu8FvZci8C1+hTBXG/IdJyI0Xnndh4G3p5Pru77
Nj7hmo4iZZdknQ8feHkNCqqv/qnuh8kEkBUyVYprJi/esfvcDGUgrqOsLRXT
fh8r/yM2LkTnHge1LsK/219N3NkL9bsA5JDCfVb+JQHAbF2Jenivh5w1IquY
hXt26oX+BhHDTORWlQBCcq6eSYqwtxUVuNtyXiXu03jci4nVcesGLFnvT7Rl
cmDU/Lgth8PNHWmn7dBjcs1RhmRaIvFadPiHlmy3k/wEwTduy4vhLLrIjqQr
YmXVcLAv+usr4ToCepcOt1Pa6cxcImFBoam5KNzMIdTpy9nB+719Zi/Umuo0
+GSxJ+9VWzHQWz7xbGwJO5RcBVwhEuhnfMjPmJDSUGnbtUCU+RYhQv8ySp1T
9jrLkF4UVCWa8crZuk58I7jOHYiWgE7woRcKWtAsACdmZ2bfoIj0dfdGqJX2
X3dAfiVS7Z/qTE6bG9AsFjfmguHTZrJTN3XbbitRJ8lxgBKxtiNrobRc895/
gbQqYy419buggIBf+6MgRGnCd38dOfnmKizu/Jvaba6JZxjKsCLfHlHHuqgT
rcJFYOa/i4ez2sXjX3aad6u+Cu0kvwo4z4RlzLxiSE5ludgzUyoHuYqqpC7e
wkKCbHZnvOYmZZFv94VcYm+5V5B4H0fZrgJR9U2V0XAoS3InZzQS3fSgDVPh
xz71aYORFsvskMf5YPjKmddDZgT12oN4UkSyRN7/tl9lgAmlucwyuUfE9IQ1
9HEeMhkbA+8tlJqq1rXMJzOLB+/hqdYlZhG08RpExjooBWhy6CfLqYzUAgZL
eM249lXNJXkp4Yu7KNuYdcZwCIWD6RK1VHd1KRjb6kt7qZ53seb3he1vUr9I
7uF/HRZ7Rl3EHhN3ynjtENpbjcrlrHJagJlVq90VsCvO8kXruXcM9DcnZCAv
JI35NAnjJH/I97EGs797Om7Iv9rZrjyiU459bzyBO+V7CYd+pPBQb1B64m+s
CDTnCz1cJj7PZyfpddfTmUs/enhwV/9kGVFGNhjonNbnghcJITVwBbJwdaK8
UiwBooE4YHlNZsBzHEIQkKugJov2EsOl5Wa6zDqtAZKa7+FcbDc0M1moMqH4
opc1DszC6GjA5nBf3FZ5iM+w0xZ5KByPNak9l/i6602gaBqoKtcBxznuStjg
2NNFYmGADq9fkzwCZl6x2u9y2fG4CHCzBvcHEDR36WXdRXRCbOKNKpGfL0l7
C/ePrQuoEZC8JImVinFT+dRGcwwo9RV0DxSSPQX9zFO0viNFwixXui9toI6d
VAZnQrUeEnTyFdpu8B6WmVYaFEe2nuau1J8yNv8bFaHlykTgGK70nCR9pXDT
PMa+m2UcAfZe9Uo/jte08HOFw6Wxq+daqSOfo40Y2mqC9vefb5h8/+HS5ZNv
ycwp1Unamhb6ZYTdmZJht+wTpXNaRIpFMg/CokuLPUEg6fbc7R4/QZaBMUE9
Fn1LFI5i2ax+0R6IplxFQaMx/TvujiQlXiNQhGCkxDIQq2dEjwhqs+WcGxpc
yA0fNS+CecKcElt6saoQmkJG3noGEvoKvLLBaK9wvFNj3nbOhh7flz81JPmH
Tqh1BylrhB3IDNBx2dDEpeZlEow0ditEcOH7DyHKxoBOnYkllPbs0jSWLJOx
12wVgMouq09IRpPRqGfE8OdiN0QyxUJPdFNvVVOSzZWktiqUCrZ9CUZ+yQt6
4BKna/va0e6tFlJow+e3iA8vzVCvjRiQk50Mkm52unvk3SIXikm+kP275ugP
EVB9cU6HPjVeBFb8XILDANZCEaJ4wPqAU33w1BC8k20DCO+HAT//EvYD4Jge
zjOwbLC2x6avtivjcWvcfjtVveyt2NbkW2NyMJ0X4cAsmacdTN1jW4Gom475
WYtJjl3Wv5dXv1l0UnJSoEjjwuN7RbR3gCxyICwFDlwft7lH54UeSOrB+jVx
KkV5rIYQuQT9uWFM/b53LelEHPbDD9XmQC9XHYklTq9Tkkkgu2AjezX8yZnt
+1GGKxYFDh1DYgFgn7jk495jKkgntY3d/Y2ZwKMY/UGxOqDAD26/xDCzd6QJ
tpAoTJbncJqQcFm9SL947Ki7ooWOildi0Z3oSh77Cvyxs0iI+hdUFsgxgBxj
IMhN3ozA2zr6aqD0sqfiVso78pa9CoB8zg0VCp6Cy1xDgAgAOFsoe8dUPVtf
QfbArD5eJgzTAXVcansJxbgJWcKqqvur5MX7Vhbgia26tMtwfS3H9XAz8unW
Y1ZYOk89JzTvXJcecKMjJkROqTs/r19In8UHRfSv58Bk2qiM2fSLaHg2JJSi
eOX+svPfoVTYiLr+AY6utiY5wioaboi+RajuKIovxB97KLSwLRMca9TXQ7BR
BgneQvb9iCand+5rUo8Y3yCEiquDqmSJT213vHIedHshQsAA1zMWEUXJWpxb
zGOhkFAljXBAewnaPRgeqrCu0nuy/3VohXDPtGj0o0UL8H0BV4auNVRufXfQ
pb2bqAX0Sx03kc98NfXGRQWVd8DRCkqZAXlEID6Gvi+vB3XedcZp3fdVWcxw
35EIwkLlPoHJWQg7Q2blODtncumE30n6y9kKXtc+CmRSXc2Pv/iCVnxm/Y2h
basrar/Ural8FTX/BDzk31X0A4IXuRpvGeEipfj5HMpEeRB2FceZ4qrdPxsX
EpqgDm+Fha8ZDF2t5eN1adEKzgthOQUprj8iwLFfW0Nnux4EuVqSnbGwIlLL
NXPVONbYw+QS5JI4ygKwx9ieFW84QRkUlJ7MTJxgjWJ18QI7RivXpFjwv8SF
CZkJFknBOelonGz971Q43oMfz/l3yMqkej/DsUvEPgKSOboLW8/mIPLxnlK0
BzKKLNrfv0PuyPnX4NnZvPZ9r9/dgUQrWNuy9Hc+XYYIyRuCCeaPxxGnbyiV
NvZzG3lf6SOUi9yEnbepEvmd8pcTHT9+rX9VgN/io4oGrKbPBINhpAeKbyli
CZWXiRxGkPLXnueN6itcOkM4pSfMMF71Ig//znJjtXZChynrwlanP/N8XN2X
ZsJhkRI7+fayDyNhY/urd9z+cbzZsaUvCVLWWMVFtmPb/VhIDr4miDlBARU0
jAnlGfE9GUGPDgkXugWv37sGH971pI9iAguwDwzY2T2+z1hPgQ51oPXkwf0y
Jbto5wkcwf/3lYdSuJav/2KaKII1ImLn5wSOwA0D6UaujV1Rfrpq2RLuCqSq
YyXXXOG8b9mE0KgZwzOEp33aHmVeiX4boWIpTr4kF2y5w857X8xq8LPKGZIM
drPntcU6U66M+1qNZllud1x3EW6SuaRCB00R6k31lZcO/fiupXRqAI9i/8MS
SktnQNCVVD/3WHSkBnxt1G199sOh46WKsDtIn1XmEa3MMLxnR1hJC9mWVf6S
O8RANF2gcYQ/n1zra68EGfMvPdX8bAY73+4yEoOBaQ5Q/cmBh+kHCmLAwRO6
OjH97eGtSB/uqS/sbZxQTTnt0ZhMQjbgfnkP4voycVUxeaLRC3xBIJVkM7cm
sjhPFOIjJNHEO7HzoBkqGTyP7QLmg3JkQENKqN1qYOqMlBwptHNZjOR6XKSp
Q29QNEiBko3PpFms/PQrxI9/vEzo5ziIkKkTXI8Uu0tuaZyTNAn2RRapBL88
3Q/NoHuIwyNt1mWN46yXlOoV6e+UvMnprOpvsdCcag+HySpo0otkCwn5bpIn
nNKf4BB+/xBI6hkn1JpIVVHfeLMSqkBIk5M5pbxXN+01oQlHcLgCYU2ilFbl
5abfBrvS2v9N4vaEJKzpVSHROGMaHGM1j2z7P7N+BcQeVgowKr3LVPKbuNT7
ZKJ3M0jb/NcQZWmBuJLIGXyp20Fwf1GXY5CSiiXKSL72jk2+40jHCZUWFNIo
GVSagToNegmC+KPCIcaY4W00CB4qJIQhVGJ4IoJKlIU6vfvPPX1PnzqNDZ35
DvlaFE+L4zFk2DTPGPYk8gBXLYXFQFyaUf74ZTTtuh9MpphhGHhgf98C8HpF
FipJcs9BvRcu0rZLCDt3dMi3nZENf7jp2Elb5lqgGYGXfVKuXGa/AhPEuzw5
iiss0+2ijgifuq35FcYfZpy7aw1YTE12q9QSFuY8E3B2iTHq2HTDei7IPRY6
fXrm4ZmSFPzGTthaTYP4e/IlnoLocaLS68YfVYmPrfVTpsZlpVfK0EvdmDPV
1nJBCADXDHiKC6QfHtYlNhdM80uEKV4J5HN6/Bh9Mr7Fw3uMYdplymxqCLvA
A406ZyPbxIxIkqnQpbC3omxeGPqxqeTzKtQgDL0oft6gs/+5TtvMUwG4s7tb
BSTZpVrZ5bYnnHZu8Za6NjFT4KUyoC8luPBPMx0zUl7zylVAfDH9u0Ac/GP1
1R37QfdkfVeRwaYnjmIGBHDs4cguJl/8kB704lFX+FPuZaknnPCE/lWynXhf
MUkA5yEl40YZEu9UF6AibScVVGYG/Yup7aXaxSURpaiz03k+nV3Vgq2YD1n9
sV3Bd/w/quPIDpYygCDVT41BrHgNn0cgApRqaNav7up8yUf7sHYmDMGOtgUK
3i3kAZ5hfDW4EWktqNWIf5yLg+pDRiDKIrbJHOogfzDlcNxu9DGetWT2KHbb
vFHHAVbi0p9nrIpE8JLe9PHU8ZyLEj/IVxpcL/UMC/n2rqYE9JGRxnOuxm0S
m0AIZwN6fDxy+PDWrLUB7FdG2mWv0c4b+7fNsCHcK/gTUzeQ8A7Xk2BwIBLu
MFwb9wys+KXBJj4bcM5/Qptj0vFbH5/+8xLZsO2TqdtjVndbDIIm8d8XOVEk
BYa/cULspEGi7NtdVDWDCfxslVUJQ9wTef2Sf+IxbxNGahYG9h5pVr7TrKmA
hXeuKWKeKKULraJjuSMbO8nIZq6m4QtDgY94XOFhaFWHp9v3V3c+zNrFJR/Y
0ZGIwm+aPhMBoXtq3etPxXFHATXnMSEH3qCIW1zDyef1zXDDvBnqo+z+IrwC
9ZYaGAzGjUOc7/gUNuPuYpY/+27iesnbxiEwbYwgLgSisjXFRD4XeSv+awiF
GQb/RQMnj24tNMopL6C0Iq/wpr6XgISDS4eYTKfXqCkUO9WEg+c6NneP/y5v
SP+Bk7Osyj0d+PnVIKD9GRJasGwwwUIFOY+UV4yCWmIY9ZP8D0hnEgekLsGc
b3jat+nUzaht+ZDvc2Ie7vd9xnWFqSQzDy2XJASk8OFcCYsyJigY7RH6Q25Z
Bg8aV+0f3Cje4CsWJPC3+bKTfJ5eIflhvxUW7DyYwxDgApKk0Sb51msAK8tQ
9dJvL+1kroPKVu4u42JQIHNWLm5mcc2GaAEaZWXtWZZOpG9Pf72K/GuPwPN/
5nZ5iEhrFEq3Fjbvy2jYU1J5CGPUz6EreLHAh6xHyi5mYFysDc2Ck88aOmYh
PTvpPHk8UC0PBZoBpLxQiqOFiadYCODrfiPRL6ym/lpp+2De5lLvlXGPA1WF
uyicue6wWCZ6US3RbXlSxD7PRSkcd9wfStrILxnmeQMRaYVTUenVC7W+Fpji
LdVvZHk9BLtQjBmtJz813SonQGei9Ivc27UVP8Y40gMl21sqMCgRLfjSnYg/
9X7WUF1CtJlHSPyPuooCy81oqQ8Zffw6JqhGaZhIcMOwvmDmaMI5waYPbqkK
iiWV0J0SnNEKZcGd0NDdTqIFiS6X9k/sKC/vGvXu0KAUTd40kQt9HTTgIQEi
oMQT2+RSLqRTqiVawH7MFLSzTq18PEKtuAsx+vgSz0WjD5SMdfASRZUcxAdk
sAO+mb5AGZ3pHgnv0roQgo48OnNUmBK/hUgklKYGNGVskVNeli1fu2qTB7tV
vFpV35Re59pKHTGrLQb7JnIsz7Gs2W1osfsW3mOFCcY6imkpNtt0rOiYpuv9
eGEH98fiKmhV58NIINlXpBlIqbQkKMs4SWBdaaK6RDMnmbWOn24JxpZrracb
WkAVuYvyTf2/w3gZlN1gkxZR6ldZUmyONZoDsEfbCF+0IUlyY3AaeLNnz13X
N8EmMhKd/Pqu73jIzKV0EpJsr/IWNn/M3U+aixiq24DA4Y5yI9YoqD0Av0lg
9Yb9BzoEhd0kJ4UhgjiwbBhyQ/FdtoY1J21+yWg9otvlduzgpPpsgbDZKzEh
rJtUX8n3NElBZI3M7SzuWce84QZgr+exry5t9fJoQdLtUo7o1pHWK5TEwQ5g
cByXaG7LfdGD7E09qzbzeKpB9bj0vhQ78EehVvc3kso8xhUyOpGCzlbaLrnQ
4jhXOCWdvT7u4XPGzxcEkHc8xQSpBBB4xbJvGYuH0NiQUapy6KjEgDoc1pFG
4pMDXTc/5tJgT4ZvjhshHVY5lBK1eXGBn04KB8f8EBpK72W8g/7uwJzltw2M
eAlMQf6N6ofN7/HmMhwMcCoMSagOBTYz0w6SLy2znftkAJnGltTtLpD/IAt7
Vgrh80+hv2Q7padUyFUJAJVYUv/Bh3/vWHNv+OJEPtTuoe75Y25GGYdKnNgM
DtPfWK15R7p1xPNrzCEqp81InhfttLrHYr8ZLxPHb/qhBcF30NltqN82v2Yi
xbLlQWrR3iWPekEN624vswW3HlL4NlnCGdgMhgUEoep+aHDctH+IFEGQNu1a
FX8v6mWXtp8Qc/lZg8SQguYDiyOnawQ4P9tlVO2Tm4HH2u4W+2myPYYwL9PN
OFcYNpeb5ygdvByCMSp+ES9+5DmDePJbN0nc1+0aPlJEA10UVP5eo/TgaVV9
ls+6xzIVix1z200ohqbfXEhNHcJaRRb2fNmvXl6xSwUrnlSe4pYWmAOkTupv
e1LXZKqJbFdx3R3hiVaJ/FuiDUr2Pb5NCPsicaYEPpBlLb7FtPYs/KkTBvmQ
FWtoEvOgMOkR2MKvkF8jnt82zQ1jMkDznFTmt0fKekYgCyh/OdD0qzQpQKDI
qyEzunhW/aALX6F1glJ7a3llxBnHfNyVMu2l96jzSTZCeaHJNr3kfP8pDm+Z
c3Pw+cyo05DWkVyokofVBDcjtQ5N2FmS4CRk1RauwbCM+6eN/Br5Ii/dLJJG
56WG4F60DZUH3C/4kWlh0U5M4iMajtDSHMYDIW3bcfd4izVoJEdEf0ktlRoB
I8GgkbAHRDts89I9d6ZSbE/9XN333SoXJRPrXhNo1UED2vKVrRLv3tT7RXUS
X4gHhhamgprqpqOqchA09XO2A4EVJE92vlJmMK2rtrIQGaWX/wu1GdbIxW3q
HjCTqOcKGlzmL8SNfohfiGMhZmn5MKBp7u36kY67Z+Iu2YO4SL0bO+WplWpR
ofIE4h3KJi/y4P5sx3BotxIztV7+d2DFsaV7mGDrwJrL9u+ZaiIhQ1UUCYhx
ot0jyW4MZPgerJQAENn5OpDmjXZT1buIJWqq1v9AptgleBUj1WUeJaKUAiAM
sDSDVoAa9INNuNjviEgkQGx+qOhfGLu4fEDzKlMUVHoh25uxKu1dMFKB3Zyp
btn8l0Yk8pvazaPAU8GFnU8iNEK8mB6Yuy1knjxD9mNVvTuNqsjW7zn9Axjl
0HEiX2C3YFzYg5NfAMQwETvXPJBipEzyNjpkjX4QzIsdwRTav6Ey5cGIolD8
qyC8C3Rpl42Xgd0tD0MpcQDddLkVChU0EfqpaJwMGB1gQ8BFpO8GUqV2ZXL8
eIGaPuC3tu7Zd9DIZkUU7fmHObQ3cUXkMKwQ5c/lumXDTd4+mJTdJYySaR0L
6CwBwwRN5/oLZUOXX35Y9WcrW2SBhhOuoOexRH6LthyumV+9vldV0z1B6Kae
eS8uZrDowZZ0nGoL+Ug9fG1cZ2TACPrmtljOQCd+nNKLqmxBpvooTHKfsw8x
fGeQpgExl6sPVURl7svXSFZn9AdJzDyRMeTwbQch3cmOxcM2+y6T4sZHxmVv
BbxejPmTLdCdneVug0HrPW+UgXrBByhbVivMOJn86YqNt9OkEHD/in3xGtFF
GzwbqCy0xFxKeuvQWd5QzWsh1K3ZGVHXQc9lGRJqtM9HG2nNIlLb1pjEPFHl
/t2Iwd+Bp7rEwqCiyqVGjb9CbsOIMqIEVFU65bBRcFtpjLLsDId6rky9PYSY
59ZeDtMVygGMBBwwRh4yMO52muE38YQHcBSPgVSnt7/g8YJFw1Jau/lSzLm9
a0glNAWnfHcs5pNvTP7Fgr4ObvuPMbvPrLkRjGHa4S+s9JanyPXrSzpYsO3o
Rp6SCfSdoYNlq3QvSw6j+GpxLRyQLDlM5QxH8nXUyf6AByZMaun6a7KTVgBl
3vAVRtGWjSizvWHwked0MKZM4xjP85sK+q/US00awXv+pEGwpoUKdh1aMYVk
zWUg9yvJhMhS/aULTQTOABlHMOCZNC7YlbVajClp5oUB89ci04LGdaxQwveT
V+Ym1PnpsidF0Mgv1Zbc2usIbgjvWfcQun/auAQbdulIOwUSONzov73E0Dp4
k7/Vzsar2RJx9Cu/mLUliOSuVRsEjt7QaI9TxZzi6pDEaBUxLbVJnUZqDjx7
sC+lw3TuNVGge/Kk1xYrqQ/8txkQqi+dzXG6TfathdftfS9WsXzwpolcNEyC
z8sWKBDEK7e16xtrCc4R/IQIoiRq+3kF4OKe+19EEmn7vzBLLQ+sC5gq2T7B
KN0Kx5c08Z3r57M6fbSCByEB5padAU7jOnp/DJ87i1P/fLdwz0LhuQpVXEyO
RKNO+S++dUEO+sgdOLUyvrkbCIhRaiZwlZSK9jrxOIi6FQnrgdfK4I4D/n6R
4j4iG8jI3QpkMPo89j4XdhiaPOnU7LVKayGjgB7PrzY2RF+NhlfYSX71G9jQ
HlVaJ1NrxcaVfxfhJtkNT1Ud2kU/F2JEXTvY0EbEsHMf5k3wR2H2cjK7QJLt
Y4hZUpWKTHFeNbvH38YB6JhyYubPYSE7CGMC2QNhFibqB0bzDrNHAEPAO7Bx
5VdiZxoyRg0ODZFafEy0ZIcQ68E2qPKvtyDkg4b9VKSJxd5CFH5epl1cIML3
RKr3zhyT6i11cr3PtzUG6jNzk6UpB+hNvdjnEAhYgdtR59CcG5N80+mI9PQL
6ibH2j0wuBRbTTTW9M75P4IlYcMjbOYRlTLQytvryQ3TvFbyf4X5iGjoIRro
CPMXcqxLTviZBJDl2Ly9fDOWdvXYRqWjDXDpeO0KQ9OBvL5D1ofRMvaA7gIy
erLEchZEVIzmBCkj0NDMJyiStRi+f9a4eXcLQNk6lzjgzBPREvFjjqjq/vYf
vJSla+yirvadUTAfwk0jHgbmlCJn/n65wK3p+S2ehs/qIOgEboA75ri8M7Zl
Krby5OguR3p864Oak7MTvWmGTny1AygRmf4XXbkT3MDMhMFSc+iEvAWR5wMY
YKWqv7g/QROed1etpAKF5YP0qUmfNghDPCjSwQSGQQZLhwBhauWh1ublIa6C
SWuZDN2pSUSdehuXGGAUtX8WhvTqpItILSidIOpHASYyR/JU04SeI6dAi/ja
ScXlWHk1VY2vq9u/dXiTHkq0aCdtLS2iCEaWF1t9DId6nrkNcKM/c/cd3Y0t
w3SANBJpTkcN/IiQtEaJD+uw5Io51yMGqGqECdqX9t9w24/P6EK85XnAgImq
zuuNOBkI4yCcT6aEMIGNMW1nHMNvnE9KvFZxPHnbQX+Iwb+HN8MDJWfsWi7f
iTAkLVOpc3QJZ2GLjQpCIACF7vvlcQW0HtK7HmJvFm9bYRN8HnV78jNkDRab
0jQoQVE1gAatEZWc4xxBoq9y7mdMnEWy4qmLshlO72Uk/mPCl/AoIZ/meOah
iyW8UOCyEzDIJnmHrhWuL26SZNnoYbeHKUcJA00YgkR+Ou6KSVyY4qZdiUyz
ayvXVpLSb7BpYucfjPDEN+iI7V6G433n4TBP0eMUAXVo2fgewwrOJElITkVC
7BWNdnLQb5pHzJc1tiTUPL7V1QGxbl4rKI8bgcm/BfjNoOOhPEveiPaY2RPs
aw3IRLEmQB0H9/IU/0mOcKkKibi1YLddneMS1npIPr76VqpnfNr4zlIFGNuH
cerT/Em56MxNzrqdt9Sm59owH3L9zQndM/689deTRuR5H2P/uOxa0RtoxBw4
4Yn0ZklSQtWAaZaWhBqWUmGaDoIpcnT90J+dvtjlpVzhFXl5h1nPXpEleG18
0K/GLlXM+pmHsTbCVDo9wxEbKEWM9zNsIBSltDFvOzToAKJgtvGJNyDJ9DHj
6Qs6ORfsXDYqYt6LR5xXpqSsnSzqYo24y57SkHdzQXryhMg3tJi/zypVSJfn
pQqSY5BHHGxaVteR9YvmkMm5I1vBRRg5W0j69lKw/STkvjOSP6Ms7XDWyCfN
MTZrbyDRbD3VvAxeXJxYZGOk7106Qowwvuu5PaIxT9/anCtKSYObTgS5xtOI
1LszZ3L1efzSnRKf8cAIC5BRMnXR+ZseY+QCSPr5YlC9ZCK43e5l7FXY0xUJ
Od9xGwVagkMJVfYYAZE3mJKUc7KyL+IcRb7JMZOuvxENDkSPKyXgXk0yUTWl
2GQRDMCPT3BsVsu1J496DnYhZJ5np1SGp88iktvr4MW7QJXgOBBgB1RxB5Iy
bqb4DP22mhsmmOYFuK6ToIYojtTfKlEIwR1x1LwfibFiL85Vqu6sY4dRVH8r
bHGwTPWN0JNoCuaJaraqaZaaC/Jp7fJ/F1UvL+8eT6jx7Hb77FQb51Ng8vXZ
pzvZDexfz4YyRFNT/V3PpQuhApK5Tw0w7ZlyZstpaqnSmoV1E+5F+ibT4/eZ
5XkoboyucYDymXLAAy6w1adi9dOlG1X6L0BwL2DsndAa63mVBezAKtRsezEr
h8kWEi0RH7e3q19VdC2sdAiwNUUU/LPov9AitUIeVxV6FmRDjUNcuMPay/aR
EYKwSr1g95Ynmrx0KfqRhSgvi2fxtKE3ItsrUDkqqVubC2zq69ipxCNawd1Z
obtiwwXzPQ5aC7gBxZRCPWGG/23CTiktx7gKCOl5J1+Hmt9WgmEwBFR8XB5Q
Wd9V8TJsb6dLip6AUxohLoyhh4R1TgywW639Y+rSSwtb/iYqaY2B7/PdG46S
DZKFbNXwOJ0AlOzL9hZ4qNxRGHkTDLBPumwATJk3Z0kIaGB1do+2ts2tam8h
2KHFFXHLUgmYldIaAXku5r5GjG7L5fJgtjEat1Zcw5k2smNd7wSVmX+mdq6A
6nTp3CiTZ+SZBmSB/xpSQkj6aDKjwpfDR/kerKFKU3DvwTkhyqE6aib7FSGf
Sa+J0BhnJblWqi7t8G6UI5CIllDf6sR3YArAl5Eot8BFYitvzAy3vWyKR+8m
vW6Q6fF39W7KwKTK9SkjW/51RFrh7gePzE2SmESZpkYGCx5mufW3BAmKpcRn
kT3lwiaP/J0GsxdYbd+VsOYFaLvUhdskpIi6t0JQOnxaQ1PghN9qipSQVXcN
+ndsSv1P0MqjwX+oCXpJ8penT70fW+1o48yyss+4DJbOkWSjpd4jnTLT1Wab
GrmmgSsTHA5KZ3IQpK+y/xqhaakrVZ4O01PrMY7ZhwcU0gZb1rfjk9IMMWDI
XvzM7t4TwafPWInh2Wp8Lh5UtgU5MalQ/X0dJiRVtfzPmfCwp2u2H5b6grU4
UDCQQFWIYP5Ps1bi6XhBbju1mNL/RHHGuzNIKHDhsix/VUqgf4advUQx0wJ1
egHY6Ei0P8wvQ3NIw99ql+dfZ6g6vdx3Fn51wwqgoX0UZW2441e+VTCR78iU
k0hy7CF4ADf8tGAcWSxvPBbaufjH3+Uc5NBa1Z3gA6HVRiCeqqtK4IJKa7aF
Natyhwi1gr032EdicGgVG0z82656AXwwshRNtQMxkRiv63TjYO09pER+g8Bo
v3N8LZyDVDgXN3JnJNNpKkC3uX+gEwF2a/eGZ1COtisZgIYkFg+8Q5DXXRK1
T8fFpHfLfDTiVeirIM73soW35FDDhyjNPbpxJwMi6Gkbvyyjdp195DBJXjre
tSnqTAuB7ZNi16dscLvtrSjZAI8NOEYgFgliSFibUtfX6pRDFeGNHAJgxKWq
7swHkQZX05aZBE83UH9DCODhaibHu5DtcT2MmYvjJkYgoLjqI4B3DCkzr591
LPAoUp91/yf5qMLX97k2+hyR0K2XKWDmmFHBOWPJ+b6wxvJjRjhs1dgwcC6i
L0tfPnATnQO+sJkj78CyU8qKcf7URDcgbP86BFbwCUuQSrXaSNMLxkS+Kj5m
pLn0++xJXclyHxBC6kdbLSXCc9bitQF1BSZfIKZyUIGPaQZEBKGwKeH0dxq7
/Xf2t1vOfJ0X3ZArVn8LnFnfekq9esP1LqqumTtrYhdHpadG2JypQAcRQclp
hGTSYj2U3+OQyV7D8bKvEYIADo6kvuLiGHfPU9QuY0Ca33OMocaZ3aQh/s2M
nE2CG0qsqRjNnkjDkH3H3Z9oDiDJjchGiOatQ3Yg2rtZ41MdoCVLk3S9wZk4
4r0C0EQ0/EwdP8wNgjMFW8MmkQdJCRkQH7G1HTNYS3eX8G9BNRtthfYW6xZC
VeoV8grLI3GgAT4bJscLHgDR9+cxhTVz2ZWg7R6W+bu55m+drcJjtmaRwWkg
wR7Y3HHOteAjerDjzzwuvVg82NCsWuQbPLD0DxKkdcrLqlT1elx0kuAcyKft
Y/aFF89RUuUWu+RZ09Y4kw02LU2oDKHakGUCvZROzv/lnsLL/MvRoxkiuXyz
DSLR+7GmchECKXLr/d1395ePWT8o+o4lHXU9O751kXecYmkOJ+vJahWf45yN
ImaAiCTaMnC1ryp+/4VXLOwx1+0f8N/wtL83pCAqQ3G6ew/auAaAyB/4SMUw
ZL889AkHrRcJ7w262TJjcjEA9+Py/PGkUJAdprweU1eOL+5vg53Rkeyum4bg
16MH3YSzXz/s5Kv2yJZSuq46xkS//GjK3jVoZ1VH9MWcoGoi664719kwA811
uxCfua+IRlzz9uWehVOuzIj3lsGY1BU/zbk/cv6Q3peqSCnFjJrqe0WoMQSk
r7IQH6tPRzh57h4trS3fGvXZyzfy2lv3P0B/lsHllz4NToy7JIcu9jiMU5m8
Lex8vT/ueAXe+mV5Jn32H4uQiDIyTq6Gn3MJYNoEbHNi0VOidaC3oUW1yuAe
D+L5V96ceU9PS4FSItNOrrtC619FRUkm7o3/6QmE2GNFq91/yNdMCLDe8MC5
AhJYZwDZehq82jerKaTxhZg2dN4RW75RIhv/7YGsJj9ETGKJWyGmth+iek31
5Hv4mDtUAin8o0rQxuZpAdcPsZjce/3uBFQytTIoGCELoOJh7TpjDs1Xlu6g
HPZDZEhGU9X09rMW/U6qkiWQtwUcjm96vGb+Y5xuVmuP08g7lyHijYNUvmsI
vN9rdV1Sxzmuuf32LimaeKuoApBAzg0ug6QhVFVTsX7k+p1n39V6KEC9H0MD
QZUaZSNaCl8xwCPn97iSQmXh2kbHKvqwnpMrCZ3dfnd9x6a+ZsHd1ljtMfKO
X4No1wFfwkHTw8YTOlWTRnoS9dZC4IzuO1Pu9inYy6Fs5kte1fNlrSEWqs9X
5uSuG9TIcmk74TxWFTDlVUzZBN5WbqZfQz85NDYXHh5EHqLpBlXVoZZPJpdT
2pOUCBu/r/gUS7Voq21pNxCh6SqD8L9ysMAWI39weMGvbsdzTTH3uIdSHwPG
3gvTLU2XW/guGSSyqsSa0J1mlbgpabpv4bwGWfbk0CU8L7pahf2jTa+9fQ+8
Kz7ATFe3MdyVbGL5u/J/rq7JiVXWig6Iw2IJwMioUe/eMNYqJLrihYJvywd8
1QP4K1XRV9G7KtwqICORX1k6BId4b5ef2qvKFtvLfREc+pWLMOVqUlNrt/8D
eohywEGQhpFGZDb/qMRacXpRauxKH1U0YntJx9pnb3foNVQa0jzcBwqz7o4W
DjO3WrJ32j1ZqaFaZ8wP3iv7NLaV29cHJSqqDLwq9PXZJCxCxUY5jXGL5f/L
n8V9Mcjb2VN8Y4Fn8i3Kkp9Wmk7TZDKchf5i8ggClaKn/m6YC40TcTcw0W38
i5XcN2hSJTnVguRVZBkzqEKBs6cShfl6Lq7vDY3OKf1Wiy1iyQzRVj2YHlv+
Smmgxz0jLwjEYU9Of1zuT32k2LSahASYWNkegbF73PSc+aRMbreBrzfoCjim
KS8aY/VvJHFps/OFl291wSlrqMs8k/iTnYJU4kl+e036xqHNyg/r43SjtO7y
rgAmRJ2oybSrtzp8uarS0Q/YJQaTHgEuu09mvkuiYhdcmq5OA0TsG4vIJPBb
k4gIaVm43IoCWFQbbEN++W5YtmdjV9qPPxJfAYVTEIXnvVfpDoOyvxRZcFoK
B9IArMweDV66gkRoIWZz0xVQHHcf958ZFbhlBJu8/HxiuKnYxWfKSRLfLgur
4RCT6zjyOE+GrtK9dX9sM5hP1VJRuiEZ4KHz+bELNwjAuirXWilloOoP2dV9
JEN4asNjEXsiMHWb0dJHSXHoKMN8e4rNZ95F74e9I0U0DzI7yR/3oOfjmSK6
jKqB+MA3R/IIZDico8w+/05gfLnNpKBVN5sT0qSytBzM3+38DUBhLkvpztKO
vC9yXlUqHi3R5XsInTq0YxKgO1NFN5P44p4365Z30q2FP1rPr46DRK1z5xSD
vHMnKIvM8ThzsTHqkbrrcuQiT/MMqLXBoEinhowsl4TXcR+xQs7bHTJQHL3h
Ijszg8Al4hsmXptqtb8fmGuR1eeHQW0hLeOJ3AUtNUdpwZ0W2NpPdRfUU2Xp
DWY0iuH1iVvEGyM7W5dAVE9jy6vOhZ97kGeqRvUshCe3OPJVf+Wf6nzOR+ll
vshJ8ZzdYTxheNX0wv5I+iSyegojl/4avlufYVMmqwg59gJds+C8NLcKQxIR
JSD4Euks1Mv+pD657BTS4pXRd2xEJOIv6GtkNyE10UOfctqm95RBvZkN03tg
kfJvCazKnMenN6yzY59wvPkfcrdrXwJrBs+yDOtg6SompFB891AbGo1aUWgU
aqVw32V0X3TWnCsAFN0ofUhWHs1sOx4r0+/QqK7TCTILBUK3yMR4BzYep0al
OIyzmreuuJe+sUC23me4wVRVsIpv++bSx+kuL3ALTKT5aVk1jPyIFlIDbWGS
/nSNkXCI02w/LIjZlACclzZqm/KUYcQXX+GvmczYiDtYLNNEPU/FfenHkRlC
kIx2uufCSl2nTmt5jseNLePuTjK2FOucXAoUDKtN8CERo/y8F3lT6/7Tsq/X
Zr82OF1Q63CeJbiooDv7dP8UAG97n2ZYUGYjtjUMzdXnpTVyo2nQIH3Prfhe
DxVs/bzZtGgkGVO/0elut5+6tKnfBBfQOwh0z9aQjHj6dEoWiFlw25vyqDXd
e/awGSW6Tau88WFbmc9GHKWnV7yh7XYsdd43pPLkNsKbZ11NHAofECRWxHbC
Fr+X4OW/xhRBEfeCJZ8K8DIkY5vL1GuIAWc7fxNKCTQZUZxANEnubEcmJ8ee
s+SZHQahYC+DJiUD2wvfSO4HxltzS4QWaHL3Sfty3RsGRGARi7WrHhDuJqU4
kzn7a3W1yFYfshhkiniYtp8srx/hLC08mS6RKJZui/coQD44YNu4vixfkhpO
QOs3rEeTzXU+31FvhQyYxVer77Ml9FgZD7MjPMril23XBT9OSKSUvacVn/w3
o9hW1ayJx3eireqT2pWzLzTb6nCXBr8nU8TzThUIOvySC6CGQ9rxse3bxWZm
4e5njTPtoaz1b44HHCm6J6ffpImHGBms6943yiTECRaeYfkvSuG6IkBQQzEb
BBEooDYcRa0fVLA6uxk3RW5/nsW7Z0rprAD8sl4vVPRSFay1XgEiy6cUEPi2
Nlg1RVLrbgfdiOyft8MK/FGNWJTgG5Vmrsh8R3FVNsUVKzQI771jSHl0JJPg
hgdpxVIKpnF3cUzFTmr9GHz12hbd/QTm0sKPtguyaqXZkOV64bLuSz9YodH9
C7H55bPFRMrVJP1rujTddekHVRS6rRrR3T4dI9cUUCkBRZH4hPlVUFJt8+Rq
yCRFXkJ8phK1DVvxVr/KgPhcQt5D8KK3hOO7qHBwU38Khx4ao9I7KKZLh01E
bdze2sSWmn5Bs1FGOCXGaEmtp5qPhLbT+tZotYyfm2bNml0qjp4DSyOzgm/6
AIVBwUmw+qT6Y0Id9V1EC+zl2p1OhxydpJgTvLeg7NjFc/Td7W6nrRnTtxBg
wlmZMhi7VSjCVmZyO4IwC/JR3wCLoI9MozZFu4pED816xwG9I9QleV3gIoPr
NoCdO6I+p1yRDQmLtKFOjsbeu56PyYE4VytoiDGhWBXmh2vo1lkB0uUmWZJ+
601MGlCfr8dL/fIo968W9R4lBfToz+b6aGPMHnoMwrb+TKLF2dIMIWE8CP0Y
v764IBFUHAejgf1kfcZ1mpaZw3M7K7dSc8xoI2bCwjE6Ii87nt/nrxOFQrWY
gqRCqLKdsHgZ2wbYnDpZL7YUB+25nKzmPuxEg/wz8VX3jZsMU94oKymeAGym
7PEnqZsT1CcL716zrG3/e9TigiJVOF442sCgdN61X3MHGu8qDa/LpJRb9H8H
w5mIT4bgJBSJxpvt2lLQVvq4mIF15s6cfAMIFTloUGEDd4wZpmWzAiwjAkjq
HqO7S+yh38Th3qO68H3mj+WwT3cPQXcrWdUelR0zHINDNzRomELG3o1E/N5i
yyObXrMCzMGXVfxHkgeO1D6I+BvCO7XJRzTXo5+hreZfC7f4uL2uxCbLyClK
XE1kHXY+Lr6GcGbCsKbC1AB4f2tHy/jUhokncW7XWLku5JAD/i31Fc58pRen
CvNmEq+6w4v2LHwteY0BSBGQuwxg2Ics4sw5NGNreVLj2sAnB0FeXFrnQUHD
7JZ48M0wyGp5EXNS3KCED40ExQgAjxhQTLMjPgNVaaONLRC1XaE9FtQea4Ny
HLprsznARMQi7VkOb6BL8FYL8tGViig1VwrnYLIgyugYQdOhA4w3HF8oCeYf
FjM6PkxFBKJ+YJBBr/Z5LI6AszJtKY+8W/XoiShql+m46wiMeHAfadjdurHh
5G1FjwpqpXEoPlhbjlxJFDIb0E0PxLbjett8SfUJBGW+kx9Z8DHcoJNf96SL
sgG30cs+vQkq/Hm5AZnNC41aJfSSeGOhGRCLOrjaG0EzYmRZoAtKTw/HonGo
kKAUrT/l8K2ZqMZ+bx6fDCik4HULhS5+IHL+/5jfTN45UlW7tdMVwtX5pXlQ
FTpJ91PPWk6yP98zcdZCpBFLrMM+ibs/lOM2fr2YHeYCMD+5FdImvln5Dam1
Br7AwPyBNct4jfwe9NSrHzrlepm7DvWadW5h4QGYD5uIRoNyIQ3jx+1cdtGk
9bhb2Tuk/rHXMxoC9sP3xxkJdV3FQdfVQ7q/lGaxOITQrN2CXwUK6oUR89eZ
PGJu1becN6tTx/m7BFCofhtFUUAkxWJI8rxgGDNEHOR/2DEpc1wtLOCjqLUI
MhRjrxO6OPgigaUXklikp7lTfLxXM3gqtwSTpHSiS6SOX3SJfunYA5COzApe
1kdQHXRhv2LkJ7xFZfNDPXirdmiT2MwfYX8O0m8XkAcJIPuDzYV1W8QUrcan
B8WEQLC6d2BMRH/5N+8N87Rl3svUO94wbR1bbJw8gyZkafjOZyC1UESzGvWj
sqeha+RpJFm9MpGFI2Mvaz2lLYc/JMCYpXbXr0QOBaSIwSfDtBY79QZJtXNM
ruEtL1gC8nKmeN9gtyaz+JRgbm+xv9Cpvw6VUyYqh4lDe1re0y3ThBSEppK2
F0Ed0jc6BSogx9mvIfpmvh0YZYW0DfhUJbS5lXgpn2QP7fx+4zBVxDXt5hM9
pwg4FaaTqIvtZAJqNRS3xlXKFrr1EiS8v8oSdMMlevN3ANA8RLzpR+Q9GgG8
hGp7R/HnpATUj4ZmiZxw2ga2MUq/qWyDh3EQlqLaA1Qg+7oExgeA8VTjJtMp
Vy1yjHAgiqeKBTTqYvTKOt33fK7pgtg3oOUE/dqJYJnpJ3I8/1W50GYBrbzu
lL5HmLlL4x1M0yxRm/xc6a/SA4JhV2vSCWOoYI7D6OvZc53lOKweTJEtxj+0
nCxRZgtKK3axFstZe7rHr6Bu3o4uvfsg82kvpHcwQYN35E4mg8rmyygV/8+M
4kEDLfbttia0qqHjLC8esoa2dbaLoc70UW/1GufkIvpC53VR+Z12MAaSch30
eO6Kg6jBXIj0Rfj57OanXp9SDO5XPRKT/gIG5i+cJsUGyxq/5xf7dtt495xX
FtzPoYpIYUhwkKijsME2xnlnZxPlYfSmiiw8yEnjVeh79zGib83jXWWLLza8
le2vamvVUa9gfCkn46n0VivqBHpdXfFQDaDUy53b3SAm6+/H8aeDZ0VmLUc3
HeXR1WHZn0ufztljNTGh0SCmE+qrmVImkGQlvUmwDwDkzwCPCadviB8vBQna
hwfyHgsM9jqL+l24qkls3w6QfdzhuzH4+tH97qjjWoXTjb4S6R9z4GA6y7BJ
eaW/3G78kHpJcRFgPaGpDwAaJOqJr3u3K6D1YVfWWI9ew/EhNuvlzLUHlcw8
SHyJmdJ1T3MnazMr2fnI6sbaFRF++Y+B6sA+9XChqLASnNA6uDND/E1CMwOg
3Hw/4w9oXP63YsOXF6OQZue3/juVBCrIbJ21nBKml5T/4n9XyO1U5+OjoZiK
bfrAP1cuseiWVUPNn626ni+Nv+gRSGmScm20jDepLsLhgU+RlCwxXyzwBGy3
WNGOCZ4Ds0sbqxPpFfc+BKQXIo6GZW6mAyJVay3BnKf5XQRNLcCnw1Le+UQB
g4v/v1Y+6s6QFD9zRztqCkrGuL1NKujOYTTEur74cetmWLTnUNRlq0hFF7BT
d4eApwNpBokl/m6pAqfFgv1nSccUK6ralnhC9Bl+CwJ+LvSo1f8z40wYgGQD
0lT7OSZ3x8ZlcTTJNmvOCQfwk6maiYBr2MrqR4E4CXWEHMEWsCEsbhbJP17C
mYnyWTLDimPOB5OD3vjCBd20qkaxx82om0Hq+C5KomfeR8ufVACYfiNmmnGP
rt6jlEVaAjMLgfncHwN123og+GAaxDmET5Z6gP5MAFuJOS5nRLneM8/zdlqK
l0gp7ylDqjPK8zS+Iwfl2dAMQ+7eHZQpRPbwwX+I/8P1bHGVZAPHCaOGqtaF
WLXYzOTnVQbw/Qsny/WBS8epczLx2iL//nel4cy9ak0jzVkfkPVP8Ms7v6Yh
ynBzFAMYNu0tRGgladwxEIi1TMFS5NeZ8gDW/04nNDM6ha/5kA+17ICRAnGJ
HNwy8ckhIdaEEKahL4i3QVYQp2iCWnjHpZYkTvMqAyZnPTt1R9d2be/tvX49
rndSfv6QQNsseyroPq4aQpEPAzmrJVyoYVsoj0bXoM/Rubx7tuaSw81Pn+lo
zsI/Y1qBSjZBOvZyMEIZ2d+6jHaNAr+5J8RdqrJrAAAgrYJcw4lYPauYSIy2
L11h3hJ771Vds0AnGVQCYidW6+IICAwdFW3djeX/zcJZTvYv0cVPCE15N9aZ
QhmxrjmS9hxcNijLhTsBtebH5K4feEgL2aQAEg9ezkLV8zN1f4gmd7kj/BuH
OG7Ni4TzR+4CrQvxHdOfgRwBa7wB8YNv7wM6tGF+m76hCHArOFUKutSEGwjo
zLWLup1XOhop9QTCeGceRnKIE4JrkUOxHaQw8TnX4BLuHnHVSS0Qbzjw9lFs
L+uUqxmGy/hwL1P0lgY2KNYxvQpdnC8oidM3Yj1NIWMebKp3mwvo15Daf0z3
DH9mmx7wo0hC3VgGG2gU1BlHvHO94rNAL3I+GxF6/I2nlukzJuSkhDgpNbCk
mJL1Trdl1nAIms32EMnJUP8Wcdp5RiNHSZzPZKMotVSeRnPpebfIl32lqSKY
CZvBkkiYId9HdIPDbwaTkjooTtKdMR/Evb0uOcVW56ZkoLPrITZic77gW/N1
4Z67/ldyl1XpLjRJBsC5s/yPzcmmbW7z3IGTkn4/h0FQZCf6varqf4+mw1d6
/9F25oQyt8KjnYp+RdQJGk2OSpFlTJHojdo5yQlaUAsoRgUb84QHaciRrey+
CzwUesRT/3ja36mStNgu1xCFPUquJV0VAiCl4trPU7zJ4ghvDu9OJBFIpT28
TxE2pmYf8p14QdUUGQ/pAKGG+XUxQb6CqX5odBZbOh9nUW6ACDCxtMF8BzhH
MhNH30r4OMZzGZzTK3vHGzXqBF1rxkpVaMvSwbU69h0RQ/pdvW+g9IvEs8Pq
Yz17T9fZmqb2aeQzn4VCKBrzVMEYnbaI5HALYO5aXciZ8U6BLpfXavrgkNrs
F54rb0Y+n5O1rVYNdwd5zfqwTQMIwWdl26FJr7LcWdhqmInnBZU9ya/FdBob
dFVpBA3SJtrMALTpMKl88H56vPkcj/4A4hW7/32RkIV+JPA7s7BPhCJrG5zw
7pErt7ElwIy/50+8P/ANK9vfqTUJnvArTT5lmRy6MukPIZFTP0LBbjTm/XyF
FQSyir/kEpaP+wUPQ4lBARNRsI67HbeocDbfNaTODlleetvsdLVUFYT1ATcn
K9AmhjnhTbgeTYNrjEuPnbiokJhvPpweoDS/CsREhIBJhPa6tLkZqPh9SVxC
L3Sz3x5WIzDX6zdsvagK1qmgGwgDm7jUNMG0irPQtXgvcUPIIkRCxkLGvoM7
+K4z4iRABa894zIluwC7Pdryb4pI5bDkfb5PBxjFO4SiEJLPjeko/08s4kPt
qWmzL1AZD2FjYQKDCKAdjW/CVB2xCPL4PQx/7uqKBCGD2gmMmyo5sov+U31O
vHvtRjoToXmUeQsQDwUF88jOxyD6bMZBtepareOJ6eVAdNWbwjMtbHJOMtNE
iRLvkmHxD14acVW+/5r5EeQmB+hn2/cPXbqyPRTYBtu48FO90NS6MbUdLvke
2wcqON3skPyTFzzphYmfSooXcIIL5ld5z455cGxukXP260tQiHZ9BrHdUGi6
gCEdfljs0RfnIo2DepnAw/lkVB39Wo3P6zWTH/grLVrom3LPSm/sM8w/d2TO
Bi0B5dh0JQ4SsBtvG+IlJpQR9YjIW6R1fdSsLfnhFLCNdRX2Qw9DEgZ6mwwQ
ux+QzRjwVVZDACn38xuibkJLN89w74gxiHIAslUqCCG1KRAzXMEt8vvvo8c0
RvNx2uYIMtcyUOYsXV8OsNLVlDOKQgjGhmVb2EvkgPaYvP+OLgak5VioSw/V
QhCQAb4QlgQog3/BgWPXl0HnEyu7P0bXms+0RV6DIZJsHqocfhe7ZrlPWiX3
jTEOyU+eHgtlExNjLSctBwVZE/h9/NIBcL8epUYJtvM0ngRW5JaNlndDpGic
quMq+Q11g/g1gFA2X4YtvjxkqGlbVakfPs3wpxWeQ1s+HCs8TWSDQ6ajRp0t
yjXYlz91f3Pvty0bhbhDcX4GfKtQTFKz4aGq8+KiIvgnMO8jN2zYC97caFLe
l4V7nlXE3yBuoJLZlH1VbPNmDeSxuIwI4ZN9O9QC5s28xFXVH0qJGsyGdIeP
iql3j09YmJpsM0XQPAFMZbjM0XP1EyRD+MKqi22yqlnBUHVrQWcJ22otj1Rg
xn8O4FJg3UlYA9oJCdYoRZsY62qZcVy0pk7yBgvPHkR32swFBdlYxj5Vii3Q
POKJSvQQJvu9w4MNwIWQ9rcapHSc5kKrL4u5pixFw7CZzQYV5lJbPQUsP6Gd
ZFqGHBSJwpFULIJilsJVGTO0THW0yrUfTSyQ0eqS3NJZfoUxWmlW9UiSruC/
vyR4ytTu74BfL1/9EYQG5LKlVVjN6arPOXEtOuoEpFip5GlLHx9slEYhl8+Q
JqcgqrPrd8BUI4ucHa0eZ+Qn9qSlXQw91bzxmhUZMfP3eTJUt3qcocnHFznr
DxJwNZyXpe+G6OxMFTkb9WVAiwNWVrD7OckOPDr75HORQlvA58TsxXgmLzod
kTSTWgHUQVvfvHSDwpcOrD3JeNiebsaKZIveK+c5cz0vNadFODqYBat38RX0
ItqpIwaCUMdoEDsYd04uLpAq3BRkFgMasEb1goM1sqEHBv77OWzu9t2U033s
o4OLWtHHZR/O3rciAwghI0MGKF6wMQ82e3QjHxR9V/OpU7CJOx5xOZ7G3nS3
Z3E6MLJ3hFX67eYXxcZ9Lk4o/0LD/4go3UvIUXK8AYs6S6czeHo3EHdivdMh
GDpQX/Ae3XF5b4LxrU3CRfwJHtRywD1akeZFRGY2+fXeWeHozxKa4jNGDKRD
N+6tLTji7vLGSZu9EXNWxz0LRF1hBkkO2orDVp7gu/q5uK/P9e9LxlIKDiip
6DRvfHHwZ3u2I8xyE3co62afIIFSCeAnclYtsr1PSvMnyvOfSfI3B8XWE8IH
q/ZwFkxjYuVYqWYn49tNWvUyRBd7+sfmj1+lxMpAIot+1yLbnLftNLjT49Lp
ZoC06gcgdbtItDeE/smSx5GPB4SZGi3P1tJgAXI0XXwWe5SCE6fGeEaJek6z
/3Ciir5WrAbBxeQ9GKfQLp0jKQUkkA3CT1LVs8JTUEdmDHBH0XftsjESx8Oc
KwXDWRs//L2plN8F1WYoy1Y0klG6Qvt3RUNyN7gHjoXs1G0apL0zbWU5s/Re
lbjGvvCpTFHVRsILtKZfHxxH/fpXdswhwWmCDGPtbI3AgZ9+UbZWVMs/TPEU
6Tzeg4nzJgEmOZFpDkVBxmjatSHsYhS61/G1jslpKiovetXXjp+9L8FEisKs
Q9KnpQ8OYhh7Gvm3KqyImAo/OYbVWKS8YtgPscsR2ogfyt7gFi8QrWWkNCui
vrfea99m7AeiOiK22CpY0Z16zZsrqm9mRA31UXys5z71q7I+dUHI73h23HuK
M50lsBHmIS7lYNlGHi7c/h24+trgFGjqrLUcM93kct32z4EIrHDHj0CyXHVw
aonaCxzhiXDPQPApRQh6CvwfNC6bZA+Wl+gpSJUUqOpu3OPmqvEgSbn90fWp
n1PQ4YzJ65aXOZav8X60tWaQFY/o5X0633HJZmAelknJHpbk0iGSFWh2GZSN
jxdmDtIcggHcG9TkIwUwO0rBs+rVOg1VIJ6XcGz27NgjsAYjm2hUCsQ2Pmx2
I7/9z6399UbwRcxVPgA6cklIe0M2iTO5kScUl4CW7Jf0PpBxV7YVOxCrQ2z6
KzU3w3v4B6y816GnVGlHzbQgPP/9VSiGcVJZdhFDQ4KNoY5l17rHElORd5sx
wzVVRU+rJaADvcEO8JrO7qAFy0nlR7JKJ000e+rcEV3ntstaNnHa3mCY3R4y
S0UGOGpIjDLArcqrw4cd6o1UIC1M6/2+njRf2aPC1yzBJ/z/pTmim9MCHE29
AnbpsHVJHWvGOARtzc4FH/MMXb7b7g+qmliyNNey9jKhHvaxqI+eUCiU2+MP
gMStz++6ogR2nUAQiA/f0vQ7HKi46rLMzvkTDUB3GRaaNuVZhUp6QOmwb5l8
o2Hib2NTmDwaRNSWeWIWqH0ftlfRLiTrwFqlii00o1i6rXwpYPB3N+c4T3d0
FxHIC9IFlLaGI7029f5TiciPMCOKNG5nmVgqrMABsbHT8lmB7VDjJqq9wVsv
44nVLtkAEnTJrNRaistqkXf2uVaMLPBUs7r20z6gpAq5sM3zRAZQYuvDRVIk
yipFS8JHK7URKDdiga228xklTVKbeOdv+3HmZ8SOAKZZa2bQWz/qpj9Hna/K
iTlELIWaLvLv40L9saByJnmaO93ncjP9EYBU5ASO2c32OlOoD3E0SNuTNYBp
cgaPK6HadHhno1zihwqRNsQ/lOZYTaIubaWHDRNOk7vC4XVwn1+bZJvJU4yF
A2Bu5nbkwi2+bESuhm/AuMiFaDTW0yvZVLsq3cI4qczQwvBZ7mNki7JqRaAR
33mwPDFc2SvXlimYHb3lg37t7YsJI89nLxRkLY9BjeVMl7lKbij9BRXHdGvX
ypdlE11syESy3ZuRl7c8E9i+EnkXeaEsQ7X9LP5KZHXSBQ4I64qePtN59AMi
roZhzkgqBgl9RVrjYS1lOvE7fTQoIxAH2r7x/AZcSql9VTHnv6Tqklg4a8Te
gbNElIFyHoEwUT91NmZq+zivU+z9g03Moqva6Cri2aNbeP12kQdNH1ZrTUAy
Sdw6bfdyPH0ccs2j0hRkmgQTU2Z8jdFt5SeirJG9EvIca3fUWpEH/YGbB98M
YBNVHZ5B72RsbpB+JBh8789cP4qWI4tajxGAVDz11o7osFaMznPSLU7v/u2P
jQmF8BJ2I1XWYzPUO0GhWzp6fJlnD90oLSGmv8Sjx/WjVfz2M8Hnzvo5SkuX
5dL827a4B4rydEkdTly1JqWwv9eNakpPRg6GHBt0htf5GEYub7YAKYJhq+Sq
eY5QPNrdcvBizG9pu0CfM/n7/wre8EfbVPdt3YS1uH21+GpqdrsVWc5BCXm4
N7iP7tnUekSCLvgrjVn+QxfVELuGGU0n0I+yDNYA3Ke91lhSpuunrcUAu9HA
sNEHr7sebc4zlgsMS7gUMg74DbnWOGedtO/EyWrRBsz6MeVYoNHroYhxFLC9
lerRVFH8J5pj35ZYQpe6aZU25ayzoVG/0kJuEiBf4l+aB9vbzNBBD9zsbRRA
wBtcureRdc+MiTyfnGMOMzUgSvshKsoAbvTs8CQF3BWRG+HdZmRKycAC0AAh
kwNFIubr6CoxnvNokSV93iz4hSSU5hbrmCMbk2h+WPylPskB1IhvocBRezTR
/mnQjZ5kdnjjVoOtTULIUt0MIJ6VDXfL8L8UT37Rf5w92ueyeM6prI6D++Bd
gIiwBTNfAMWFTsQTC1cRi0fqnyTPM6hywZozVHhnpPCyRU6G4mdsZWtum6Dz
GixXIlzLm8DVAAKqdwEm77lQ/jthsXi+bzLkAI6cN7+fuzqv+9kCpdFgwb6s
/n2OAhFbDcPwzns/40vHpGMKNVlXeRnLvx6zsEGRoVy3XLxH+jXxWfprBL4V
yZ+SonVu+TkMe9sNObRnPwb+yto8fb98hTrVOD1HSERCEzFQ/bpMEXAjumGL
60rvi1/gxQQmf2aAgKkfRS/+/N/tntO87iW7P139a4Gt9ttjCuWwI1A8raGA
DsRybq410+C+Bt5Fs3yR3WH3YOlgZWfsoLvYOq7LoUB3WIUICJD91E/ZG//u
yZZwgKsE3OxZOGhvCG0DBuYMTFvUCsdDgePaojmg3krc3hfbhQPcLaKzpuk8
OaDs+uJMslgVYbDwOU9KaAXIvjMtgsXQU8aIEoGea++mNFJ7z91kWZr+oGeL
xHDvhBSxQ8WDhOZ4hMjNtiG1wZtzceRqIMCQGHNFdIPtFLjd4Mr16m+1AgjA
mZhDKOREHK/D3pw6cUGdfjo43VGEtVkYivgNLFwGLQPw/7NeG/Pv+HehK0VG
Wn16EH69hzjyD8Z5Qrd7SpJCgAI32BW8sm+k1OCo0WUiylqj+HcIxESWWVh0
/B8sTvr09kwNzjb0YMRaquipGadHx+QJL3GvuBwLvUv0lAPDmbed4oEJI9JT
5AzDH9RgfkCCrrmuRn7yFrCgEwpjP+zFqhh2pmxihrnsxbZSNN8nnm58Lo+S
ERs3ZSn282dsVDkV9fhGw4qjUPvVSEczPzc6sk8LLEjLyrZwJk5j4pGP5FXb
G+g0KQ9Y9oOTEKbHCPrBaAqzYzvMQIflEqoqOTGCVFwci1I6irAFGAOwjn3i
1t7Jxm8Or+YSP5Z6xRgnbFufOL1VL3W885ABVP2i0Wsw9be/xoDbTxYS0rhz
j2gCJsBKbFGV0Hq+nf5erJc1Hj86weJHP23C6E36ywn8hgnweikQJ/vds7zw
BH3vanA7k4s3o9xBaNGgE9b7FmxfDcyXjNPRQfdDqQSt1mlZ6WLEE6uWAIVK
yXjB544RJ9PqeVg2xV3+221YyKAt++GocoESZ2but47sCu0l6xr+jMvQMF1U
Op83huY/e5OMGyXltawpUkey9bsFJgwpa0fBDoogBfG2/dnac9cZLaXH8OY/
jNYSMgGE6S1niZ1Znq0KpuYAD9BVi/WVYzHzqe7AFs7Zs0/ui2aTcMvhspt4
RBC8S0GKqZQMqZ8gDHqHiFl+iuN8nSQE3wZudsCwN2Q885wSQLc3FUARI3Ib
rRudHGjj8r7f/Kz91cyAe7ygyNFiM+x5NN0HeL9/RRfzVKIVkvsUvWJmlXr2
pysNzB3+fD2JX/9NhaeRg38ZaKW6XOFs5tbTaJVsfH8+7oBqVwRECwHUBC/l
NNvvn1J1qlvQDxl9AWwcw95ggDlXVKjbC82iXegPbZGDtpXVW1eyu9ZevwSY
zLSMbxUgmVzyBo6dULkoWKQte5un6bEBjHhXlugA0S/BreEHekUz8eKJkv0a
itEHt94hXaCtcB+wa0FHkBbNrdLV5VcRPRlC7M14HlALShrBYn7lblxg2xu1
ZviF7S02MemDWIWiFbhSIPcqMqL7H/r8GgWlIo63cgHWzoeLPaxu2tl2sC5C
xi5ppDVoL73N2wPSslcCVSbK94xSYNIhyyZORsjKv3IRlKykgeWm9zQWpPRh
Ak59IuN4iggg+WtgAEi5euKPP4TwvnFZr5DSIdFQEZnpPFigGbIgcO7kxRXJ
itjz8k7AE2Safl/FuCfQI5sZ/MQzYDMAUlh4RYU31XXO+N7Xy0IFqkQNsGPu
HVtItM2CDYMx/+tYL9N7sJHw6BeW9mn6uU3P46fjmY2PbP+L/g5RiT90V/8B
9hBnTIlOzj5U62halQ07/duV6cL6X4tuL7CSudYy0eWVd1ai+xM3AsGe+1Ka
QEO2MIt1fPgJLpw48gR0NkgZdlO8bLO97lT5aOdyXxfmJbOg6Af4HNj0ekhR
Tanovh+zEI1EDacMy27lCjMEXFZeLkZ5OJf0WUlKjxbZvKxHMw+gmOxabmtG
lI593kW+UClVHop2Bq7aTk/KJSvojVL7sRRRmN9iLWmIosSCHyQErwyNtN/A
kbr0uzLoj4lGlcaMNfeANMQxbMeOREFFcawKPiQ7ebdLvGjSTKsPz2AFYwPR
ot3qhmeHUKLcjcevAvmJVnYaGvSYmPZrXlXd4HkTwci03/8PrYhCyFc460GU
h7AF6EJoMXxOcxJOBDlGxepRJxuxiGp4H9KCP0wER64CONNUGmDEurgxtLBn
xaLAXTkdQY3d1jNpQngKvV/as0/obB/ngBC108rELP4iyj0+XNPC6+1FZV/0
xw7bM7iEsyDZEdXfCZwuJUevyJuxRTf6UL0G1XGaHVYu5CpdRFYuhfZhXkj5
l0IbMJt+oz9glINex8N5IlFolvGSTP8uQhcuwS5UjluYdxjlUVwCAv6ti9g7
LwSx+RQ1S1BgUjef5BzuNkcshZ1BjPGw0bYP4DTfHtpUlQYjGh6SRUqoU40b
TTXZHrCvbskUYGUILfXB0vIYzDM3jNBb2Xj+WTeUueps8Olm/eqGx96rxUTA
rtMabJTnScdXOmGqaa6NwppPRtxF8d1jhie91nUOem0ZOGfZ7BX3PMGI0uWg
dadbGSWANKEUVnAvNIZPMEJWd8QXya3xW9SP/gQCp9690Ff0YcMVCe7dNHka
h6T1o+EBCZl3uMzF4+CAl5uUcfpgXAFEH3/ypnWvJxXHYgm3ZYd4wADt2nTQ
h1DShKOTEDYRxTcecVc3M5lBLzb8LnPcwMFELfHvOvf7LCd7K8INp/I6Tna8
or38aj8BRVsKZXeyjvfNC1Tz769Dcn2+8jgG9/Gjh9U0Xb6tnrDtFhDq/+sA
XXLi9HeTAbVjzTErWG8V6Z9bSnvLAyMVoHR9YXTS/jgB6m+T43QywKq+AaTh
rxEDPO7Kj2manIMhtXGGRL1oabog8moHIQqCSncfd/8wiVaft01/h/3mi7/7
qPGs3t9K/Zt97aKtP/aHz2uvYnsnvuE4ys5iPNRa5IGJmqAnj2MoFwhbpPm3
DJ1QYFmERv2KTPNEqFfwDieE/Y6yFpST3HdHbIj93XD4WjlOwGDJTR4HmoFU
FHdJpt6VedNzOt2/r7/L98FIAmD1zIputl6SgXqf9oZmMTFLdFE9GHq3XYjK
9Xi2N619am7lPNyslsM+/Styo8CSyq6oQHo5IlIVL21capcaictI0inqDo6P
ZcSdLWJsE3j6xclOAfgFIUmUj3X210iXOGbqypf2UBKyWtpT97/WX9cLjE+v
BGNRaYz0BA7Sb5QIeFC2CSxi/0m6RBZ1Z0oiPfF6DvMRNRXytD4wSZ0CTcqg
g/0wkxfkB2M5uvT1kIWKChyp4P8zdxvPrOzhTyhAsUGrNiu4IYfUiY9WvTxM
gWi8Opc3fjZGRc8OswpGmE2NeMFBus/n7ifO1jyQtDPpk5Z75Sg9cdhJqD9E
uWBIiLAfnhUxieQF+lrbfyiNQ+PfypL/Zjh3LtyUl0U9ZSEpM+7Bxn3CTcZf
14GbDRWaJI9QFqncEzyqpajE54I4Zotxx7xvc+lruVn69hSFhaW8sPrbJony
S410p4h6lYv2eeZka0o2zWPOBz2R8y2UbTd8ayAyMXUrNtmn6VU2rlHDiWpg
194jX++CKlvOoBTUWeTltFT6nrshosLndut6XrYeP1KBenCS5P+8LigFPuZZ
asHeP0v64iJfyr29p98vXJ7nJv/r2AzJdgUqw7+qCcDILiCsVsnil6xQPFzA
L+ud8yQxgs2MZjiKawdRD3gCHOwzcnqPPC8W/k907c8D4vt+JQnXuJ+90XfC
TkRU2qFBLFGXDu+uu+nIcd2E+W5Fg5UvXnx/a/cDvw4ZyXymBQsEuPAojOiD
ytXdbC1R9j+eWKkAoe/Rg+C0VwHMF4nDMXGtqvevHDR00KtGFl4PLvl0GYCY
swndoZ6o0yCsxYHImzrLb8ACggGQQWjkyMzmKyX3/i9i6Op1zXw9m2lOK2Lp
pokiDqjZJm+rZ2yEuk7/TD+ER1Pnq7jS2pi0GLUQm3GJHV2U88ZZX6l3s5Yc
97SVnE+1xJw6S8jDuId7bXZRYesin2f7s714hxwGOMWlujBjba8BtmSnF64G
kpMN8MDr6Frl0RP/FYvvcvzPm2oEhRVLq8kHJ0nNiDPCmCHwg42pMCrcnCo0
PDkMsPA6LlBi0AZl8X3uaphcYekpKkBc92B+QyyedeUuiqliA9I6YiV51qO/
2WEcqEBUzqGIjUG/HM2jGZEMvej0qWkI0nj2I3iYNq2Wp+rstIkoYuG++czm
dY5nRgQvQ1bCjoRAKtMNriY2FXJoJXyaLWTq+Xh2g3ugE/HmPI7xilFD1DOo
tJkJJzWKwFtUcs9i6vYPxtwkPIpTq1q/2jF21Qp6p3Doq5siADLyWD3qfBNf
2VRVfpz9Aq6YiaqKRQXuIvIRHtFHK+HvaYkFNW/mo8E6ZgFiqtrMGBdsM18C
10+WPmF5+QgifGbgKez7Cgs3fjppulERk7P+R/dBTfRTYckh1chroD+uZowM
KJTf+D/2yQCZYB0E5BRlADKxJoBte8c8wi8rqNN6yeJfGEpUNXdQYncD5+df
jNJcHX/nHiEeSvpQK2bii5m24sD2MkexuRE9ve++RYruCVb5B5NMSsSVYxQ/
wVUUyW2vhHWBpIH3hdxZJk0Iq4mo6zpEEXqtMSAESre/YzYuztq9kqBdWYTC
3bej5xffwPvOvXx41dAdWXGAr/wHUUXLZROUKG8PLodNrop9xXNI6/BniV1y
/X/lbt9Wvh4mBE282WFoFZOxLd3CQrj6veWP+TxKQA4RkvMYudMvxeKahzuQ
ytG0UsOi5O5sgkQa4GySMPSzF+lS2yk60OXFNGHyoEyLA6M3zmuIpfDYQDoO
PBruQV0tyJoJD2h1N9mM4c0rY9ml6En8KYYD/gVxzdwEVRj3iLLUGAOrNOke
zqfwqN5LNXEp2whIaa6bgmXYkXom4N2E7ss+ejGjI5ivaH+8eWLWT/53gNVD
gwQ3M16YEw9Cx1bEfRjsAZteEjk9/J3hN7nn15zk+Wr86DYWUF34cc/Vskz1
DGPB1+3hSdPRvF0tUBoWBJGGuVElEBH0x3wHdwJgE4EHKJZXjQeQm9GbpwIr
ycUjGt+nw8A9ciJ908SstOtAbhsztXCXjxY7Avin+RuqUNCFae+OKx58fkjC
8j1rlTuxzSKJP6Cyul8WX/0Y4VLSXZbPoF8TgKZ8R94Oh9Fo8oqAfXw17kIP
g80VTBqBbW8b5J8hH7JjFOhmi2wPZ7JIwnXfINiFX9kBZKUkX2/7fzBQLRln
o/bGUzI7vVvZLGrI4DASev4McQtB+/3pvtQ/MxuvD5l7gdbBWcWi+Wdkn4/N
bg9Mhc2G2T59BdjdMnI2EK1tSmM3V5goCSGPZBTUvCamJfrDj4yjLqT7umoX
oWeCLJ+0029Ix3QRgj+eIDNvIZq8y/gkh2TQ2P9hcrRg5kiIYxd+GHX4e2lI
qWd6VPV13euuKB/Q4nW3Q2PC9m06l5V6QsTXxApUgct77519wCgNbva55x9n
aYnc+vZo37HDkmq5a+pN9UIfzsy1JWq7e8gJBAsBDBcsKIEYoSi+InppaACV
kWWKV4aQGMAWxlPZlvKCoMJK6/Zjat+7PaE8mqkAMuD6G7SUT+VahmxStEYZ
XOmZ3nmagyzo3yDltRFSITEtZ/fAdLnq4rnxTjVx8ItHSDPe5AHHrTdHo/CJ
qY5UH6qixL73mV7c2Wrwx6y0/Qe2IsCSnnqw/k3P24k3AYW9qcCS/026IXIe
jOOF9HtjMhponTWjkaV8lFYK+auoLa9Myhny73nkEl0I9ooltt/T6MtTjQTE
WrVD5p2E6ENhy+maYUvRKR+OzkWGCyTPKqXah2UaMl80rXIsYImjSZcx2GPn
5qo8z96JmOD2dE4t2GWYhNoOb5kzTjHLyHlX4AF1pYMO/w9IsjYZW9e+iCiP
vLh0ooqZhjSTmldEl07YF4nDBoYkeS3vnuoEhLZP7d0Lsf/G2zdXsN/kGFE6
pTtG1HewumHXOke6eN/tbuFC0dZUVScpEiJIE6/151/nqyCYNoxZO/gqqPvp
+ckI0WB7rebEIFnMIlQNkkwm6OIj83uSHw3o65IMAb4dFDapsHXHBsYdRpMa
Ad3rB66WvMMNRekP3w07UAIpENHsroETHFFi7KMaY+VEAiHuEg1QgYxNCD8+
BDGkF3f5Ygs4o0AQtodSWBdkHZoQ/SfLVXf1QX2TQvd6+16rBDHO7cE7cGcU
/G4gRVXacI6fUP4W8WQmFjTYQwWTyzvp+DucNg6mTUUHbK5kTAHsap+/fBm/
SVpbQ8GqjNPdY3QsjuayIWOk9jhdIKMfp9oJE3cuPOrbJ/Y/9mOej4Bm/yqK
B3QH3Vfg6rxJlNmEsWOUqdmxWz3u4C6RKz2KEzGNILWLo7twU+Zy4b7Pujlv
3NgG6HlRnM70qI3Z0CiuhCyhhgqedCTl7pM7EqKfLTE95PDza/tn7itinCOd
esaEOkcRblIy0hQ6TUNp5HslDwn2WtrNW/K4YoFWpaw8vL3Euthjmgnme19B
N1IF4eQ6VrncuHJXV7Sa5akWVGo1nB3BNdWmhoGRmzj92hQO4OR5l2gqG56y
UAc6XPO/sLcp+18E49GcbJk8VofRo0hseGmf9K48yJEUmIDG+0EhSN18dLtz
kWFzulvrH5YpHqSTy4IqcBHtmX6hpSHxK3QK26BH5LRofTPiwMcxoa2mMxzc
ncaRbPike2P4dx/d9YfJVNiT3+Pq+QXv14c3cST7oIQScamr5JHqKkD5LX+P
9kcbcOze9klzCh5ylXRiYLE7eNpEWwOek/rAajdBBnEQIDB7beKVeEMUF915
3vc7L/3FJTD6OLNpcqtMJvg2WIA9yaUpT2eMvPHhif3CtGmb2fEHHTJIyxKl
XkE7G3yVJVx/2P875aXIopztaB36SOIgLDjfCJGP9/ykJmsvY0eHs4q50A4K
OdkSsB6kT1lKgR55ri3vnVaMHmOJDENV6/mt3OFPCW4Hg+fZbqlfHcqYZTP1
ahyZTS9mTfBxjbyyGhnVR8C3f90Euxi8mdzQRtBMF8CJejhQq74BpOVDzuL5
V9ts4LbLsCikLW5Rb/D8jlV0KUav7lDYhbdgV5HUB7kVyqJQ3rnMN26Dwvi2
JdiY6mq7CW3AmbwGR0YzwyognPai13B7uH1EMRFKdbworWZicWf6GuuH+GQP
dEx30O6SUqdOwoQDA7gTAo8gH8vNyue76+UCv/CLNU4AiTVrqGOEvRMfynA5
s7D3wssIIB3RzjAA2gM2+HLMV5Q+YC6OhGzegqVQK+OhO3Pr+yU8jbuUdbYi
h03j3lT1KYG+2mVjpHOm1WSK+Wrdoosj39h50IkfLTPUhXHfSggta2iEJPHS
GcgIa9HVcicrtUqeXT1ytR8GvbHTBULIN6BfVRY+L902sqyJePE9zIFKn0i8
/Jit4nZDSNh4R9F/4rFQmLotdekWmLvIolLXcAdsH+ESXEPwb64qwUuIVSrc
BJjMn2kcrf+OQXuQhtBgWE/uq8w1UyBOQc0VvD3ExcBkbkZWJWYr80KpiHK1
glZSd79sepwCqKxccY3wJvsVWHp2dqLmcpMpirMR2p4f/m2cQzZx4NeBQ960
iTRteB3sWzd8VBC5J2Vc9EHEfF/qohX3K0uDwCA2DpmJBfmG2s2qrY30NtQd
3DK4EXGOnnvvuT0xJUhcUytqSO9Ii3DKnLXuXqvvST198wyqK+h/v5mDH/qP
/Bn3JQmcUUsInSijTraCmUafrTI1p1m41zGg/GaC+pnWy2iYfLSfz8ySB42x
s8x+LP/C+Ags3IXvKgJVqiyFuIfz56laUkh+DOXemLbbaRrTuZV2Tm2PO1H7
6Gee5t5hKMqARPizMFzjVjNH2Rc1ePclXPy15Mowe/g+WA/yfp4WF+x3OQp3
khDns5jB+mdqFQ42eoWxWSxI9tGxqJjwHp7A6ETGE5EUgPvj8myC+E1LdecT
PIvXqLm3djPHmksxg/UMxYnKfKobGJWCyW/UIbL7Tmp21CbWZvQGsODiMBMO
gRNGpO591l69Oj5o/XHpLGcVP/Ho2WfrN6W4/sdbN6uQcQAJ288hC73D/XHx
/yEmm98AUoANWeUIYkH4Q8Y28gT0hv9d5xBJ7K2lMA//sHRuym3r/XZ5+j5L
exBFWaPL4WrUSr5pgissiFVCsR0A8u9h6iBBrTcPgoF/FLmqgcdi/+7057or
jIZWFkBMrHhRY3Nm5x1+N8zrZyPdkNHvPFO5INWyKSw6qMfCy3t4uexeSrYk
XNBn98y68Qh2kaVu1VN/a4TMZwGojSbk177tIGVeMlzjpG7SnaKpE6W/ny4N
poLpCi37waKkef5R49qt2P/zawnlfXGiHg50B7SVstp6KlbPKfmuS9BNb3te
V2l7hUrbS/ZiY0oFIyyNMExTmeR9zZrufKCd6BxGW+uIg/HDxmDeGzHI9Czb
aU97/K4irLwV1eEgzoW7s7mV2HfFYJSWHerDeouA63YhCmvGd18jVCuJWtW+
TmhKxmvdlClqZbVwffA2m0F0Z3kBcu1t1D7sElXyG7vH8jfpaCS2S1iBu0p9
MwfSuSaN87e9IOlkva7gfEal81xz3h2GUHEMHiXRIDH0vC6PCYGN9+Y+Ul4t
R+PpWZYiMlrr92IBozrqKeRafJVKxQSgH6kG43BnRZdBkh4Veu+2cA1Eo47R
msWPHnBYcx/zpO03hMkHPGwQ5ijEXcJrkuCVweJf0dSrA1I/DPRrRAmaSiKR
fjqO6mljdm6Rjbn9mi2ZFB8pdyOsN1W3bd8Glh91OtxCoo0EJclpH+2LXmEV
M1kIO8mSd4E1xKz7gQsudqhfXHZnbx2lwLt83oRd3O2egtNaGkT2WI/X0u26
DgXRoQw3OcJnVNt0CdmT7WQHmo5gJad/c5hdkDmP2/+uK+YngsJ4P09UTEzh
53BKagrDGCQ01bAx9yZBJmFe03xHpNL5QKQ6CWFot3bzytw34Mg939NEuRis
KoZ2+gQDQm4ikdEosI5557OTwYf2LuAMY65ffTvSOxaonS1yD+CBsRVe+Yhp
G2TpZGfplA+qFWRRhvWIXRyW7FoNgCp/tybFa+6EDyKbRHryMKgAjfWffrXx
d2cvhDBpC2C5zBhB1eNK/t1hUUKfGdiMH52Ul3NpzUAIdLgwKK5KMFJSv2od
yXx+C71DNHqAXkxGsemMTggdV98ZaCk8cWY8UWT1VqpXhkZM2CsIv28WA6Oh
fYtHolvkag0S2+2SJUOBdrxpazr2bQaDtnJLl1JzqsKsVmS+8se0AyeuWiqC
agS6jD3MYD5RQyqGZybxSBnMnhn02FoD+tuNE1H6/X8qfBURQH7KHYJNotbS
ctboYBzH0XfvHhHC84wmwWqNlwV+zVXgEihmrdBNIHUdjh4bV9x2fFki6gEn
dgNGwYwXifurwO6a/bt3H22DjAYxrpSfxz3SIKkxYjILqPXXNDo57slWgZsg
oZguqp+YywtfJJ+0rDVJEGLbeI6XauP8c7309G8rsZsDl1Ra+qtTmlaHQ3xo
RYT+qWgxMNQr8J7YBRDFQ7xPRnk5SloNgknEgBOy+2pzoId4ws3AXKwV+Gyj
dpfTYo2upWhoRRPU7/URdfJ9uKHsOkYLb/laPOTocGKSW2YLRkQiAUkh6l0l
nk3LBFYMhXfHxztdBZg2VQJneEH0ZfW6Kj2vcQXE8+F6znuNdJ1nvurjfcwM
g95hL7P5QfEADIUowClK+zigd2SB1rbJEBCfjt0TD93zx7D9CPJs2cCUOWZ5
dHsc8zCknTAThlMWiTpMOEv7x/ETAbDyr2Hffw2tRCbj0fbB5kqrCSKsogD9
CHQv5fToiE6VmLkWjvI5ijFwGA4icm8BZ1G09gDtxE8ZsgkBGu/5cNesU//p
V8K2iVczSgeP1LuQY9//EPGqslIZho+SGPXKh0cm/qBzsN7WxP4lN+ixBL8r
IcgyKvFl2zEDlQvX6+nyRLRHP3SLvEetQKKurDsdU+nTQmNRnccI7mx5VDc3
Nuw0ZCwc7IupIqmNlP/kdUuktKpDQFqVMf6+fZ7ClyzWyw+TQpKgQMyQWNLW
WGp05lbmU+4JsPRQJuXAAEeIngwxG9y0nk5+qWuFiwu7Ez3/YzXNfnpob62w
BYNzy+ilB4tKGfD240/A1xKYC+LUa9+Lr+OetvlOxbNPLgZx2tU8AR7Njl5T
yOlmPbpwG0ile76is0Nt5LMU9RJ8oO8DoUuQq+ijllQnZAEqNqtzpHKYKU0q
MyxIKd+2thuskx3ApULkOBdQxkfG68psK/zK9cPeknJPvHDR41JjhiNFnxS3
BkYY2QQUEa5l+cBvPS2MfGwbvUr/wLYcuXxE1NtRjTOmSrccYXyNhhagf6yh
2NL4gBYudQE1Bla0tzxogHbLkYMUkHLoGbyoZOhsxfXAqK6QtRNX1T0nDY2K
Ub3WodZQLs+XRmem8aMR7Ms5kMJPvdHb3VXj3hGnUgOL15XeCAFNuP24JOKT
ADMCxaDTuVVanOUeIGDKIdG7bs4WDrrdppbDsLIl/+tVkkcDqgYbxV5wQmid
kLuPHb38WOO/47Lokmtu7UxyxJTFvGWulOe4BSQD1pRcLWUYOwUjOlaarOhJ
rDmKE6wXUYKdrw8LAPN6hyxXAz8FuCFmnd7hxNpMByRSN4VuJxhViSNEJRr8
xg+foBXwe4SaZ/gL7YuNj9Nc1UB2i1BabXnikztw7OHn2pp5/QOloI2siA9j
9jEmVtdlpxfD34hptY5lwu3gqKSboujk4cOCXH6P6u3/Ccr5LfDUSHKNLj76
V5RTULAmYsTVQF3v6VNHjJfY7W7OVrh6hRcFIBN1ggcI1Gt8bWmkJrMxuJJN
HQJSsWOacWDEb/itWzfQLdIebts1nmwrUAkt03YG7Pyv83LUudychPoXn7n/
+r3LqTRAXJaOXXGBQ7Nj4IQTWRvDMbGJDJukQCNjPH1e5eFXJ0UfxCV+QTTH
myUpolGZLo+Ea/uszZsRSn8pSEfAG3kuQVUfKRE/VPgA1sQD+EY/yG8fwNxz
CL5VbmMPbdhoMjaoBWC1cTYgv/tZ8DYe6leWw97Zdn5dl9KFK6r0VA+igRxS
8hbsuxyuzOCH/LbvE3SeiI0hi+KrwE+jRR3TPYpVnyuQBKzayk9YFBksrNop
J32/ErhnCp9s9FbJyQvzWptiGFWbVOl4EfwdMIaUzKvD8PzNzhiFMoCjZbva
p5tjiyzM6Yw1EDYZAy+CLD6GHreCjUZpemaG6BKejovxaKFNu+ieuM2FYdwd
il6yZKYtGbc3SwR/ZNHXW1lRkl5UH7emq37TAtuKd6ptdoZD7pTO62TJNlNl
h6UrD2ZN0rGh4+kzlez4bSwAlwFXkR5E3I3fIIe1Jw/vV/QGN2Ay9MAVKHol
nCndGpz0fbveUoItI2mDnGTpfJ4OwLNi0/CbOeqUS4kFQ/zwyau7xbcqOAiJ
78rYIqEk3xtII3cpf8IsSqqHABHYZT8RL25Mrlp4lHQu8kjYNcV45CpSjQeI
NnY53PH5EFF7jE2PYjZULL8awFNaFD4kt92efjXFk8f2kODxC1ewj3N47N/Y
Ab5g9OM6hUxdYNWv515PgwY8tuENnhV+pWZ9uudWqN+aRnfDqCAOetBtMnGm
q5iWP5zwIe+vCbBI7UXOa5jb/sG4qe0t0Mmy1sC17clxwEpTot7OGsOWbT0p
ZNAd9Daj10mp2Ck9K2Dmx2/vldE6pM4SLbQxDt9JGm39DL1GUkbGm/Ne+I6t
0lsObsQTG5vhK3vgpTz+0HRrgw2h0mNyh1AjYD6Y4cMeP2QAsaPjJtU9rXdz
uqh4GtrzezeK/D+MZMwKb950ruZn4wUuLGhTIYJus0qIDEXYOR5apQ40Irpd
t1Zfha6I5xiQuOVNA8tzYeERZW5+jr3uerWCopUlnEbagcNbM/Xd+WTJBzuS
PyyVE70Ct0tNVIMqLq+303vMuUk41oHLoMtA3NEYiJXVbZCv+2CM+HUQc34C
Gfns5Vpw+oXVekQvcNvOIxG22LXJKu6Z51+WlJ4k5BEWPoHKZOI2jSNSo1Kt
HaH0jeyegpyXC2t5Dyo65EBKY4+SkkjcYCYNifZNd6kxu1FC0FW8r4NfFAYg
1R02UO8YZcU1TBnVUVQIRli+RxyZ+KkbABuN+UvDta8Nbk9T9yPweQcUoVXX
KhH74OBMmhA+l9bJB+n5ANK2umYk4MJIcSntJYv0EWw1QD3ADZbiQV45TWtT
WuAfDFTBe6ImcLAXJk7d2FOf/gJlTQB5xoOWpDyhndThC/dEdTyA7C75cgOO
YAfonpr20yfL+y1g9Hy136+lRhQChspm4HPW6qtNr1ys2mmZAFWwMndMMDQn
fq4fRj3AurhyOjh7Gk3o45iHsZ9sYVXGZtfeQUgj6JG/kWSXM4xYt79x3dPg
1F8cYkEVmDo+s9pMr5aYcLocPbw4i+jRNw05YqhDGS1btv5i883LY9DbgMPo
t/7aetdqdsSwT94RlvFv/44U75x03SHRyJI5JvIomMoM67ypOSz5sCdA85hq
9wkTlwRejsu/c3QPJ0QSEsmyb0GkXTWIlCpIZ8FMJUm2wY3M2YNP95v1WvKn
lUxfJr7jBDRi/PkE5cxwZkphDFR+2/rtKaLRBEXkX2wyLOzNGboauP9BCcr3
asxegkHQN5XytKzHdq3HL754flBMNu9Y8PGzyXfffMWTr3NmwqluL8W3gcn1
uwpp32Cj4ytf8k5QP9e/tPB2jmvCmkVuSR2EQXJQOR50G01YN4jZ8wM7M/Ik
rlsQQgeLD8g905W8ZygpZ5FQxtPhd5nSD/AY7Nu6uVKOk+QbIOguG8syRFgq
HfZc2HWemeBy8YhSaPSIQYWhTCrBTM3gGo1rXOxHPe0OvpsuuYnMr1/J+KV3
ugLShtPjPiy53D1w4s+zhgP2NlE8QiXBnDMXX0uPgyIGPV5bPvhWlAFkkLv7
kbhiGA1CK16taq4W9X0lfUudhnwiwI6qreQ0wOxjo1Ffojip8jjdrVbbbZQx
qN0Rmy2Pt6GyKCrLGqnC+4xNC2f5cLDnjxXGgUSxYL5Tm2+ZEzKzjfalDc1x
YG7MhRKGPmcRBK25mW6Ldluq2/PwCUQM2wnmBTBYDe4qCXSSRYVjnO78+NCl
pQtJaWydapddu59KVEqZedI7ogM3zoY8CIwLRQHyXscbpRTyqh1VdyIf1BIk
Ht7s1spOM4/jJLPLj6rzxKDI4XYgrvpxCQ1s1WnnfcNISfbaD5fXAF8fYNcY
5vFuwa0IXpNzOJa2bXs4ffNJueSch3Qe92LmbIRtTNOx4MLGzJJpn48XE+BZ
qzVKRcWE9ia82E1TzEu/KHmfaPRY1CjEgpuTXq49OzgPtPGFke/Do3I5fJa+
uXiRrpWz2PU5R7Owli4dWkp98LvYTprlzuSdTwh66in182L85y1HKLjcn/YH
hNe/u4jW6VvgQU26VezS3zR8aRsMXvRbOGmSw8cxi64Rctto5zZaWh8v+b1m
xcjXQZ0u9o9Pw/fqRdaF1IoNTyQGqZlLgE8CkSNYeAcHz5GiwNr9eSM8MxUt
u1NEbYJj1see1S6o14QwTYgosHJ8k53hxm+ixxWr/1NtqrlL5Ex/afO9Zgly
tZZp+AT+/XPhFUfR5re7lVL/fpfYwH1cD0Tyl8Lbs/5kmcBb4tsRd6LWfACw
YX/k2xjPfpiZlgf7vE2nRXrtm97EwsSsqaZI3EHwptUNsqj2zt9lPx7LRFwq
m15jiN6O+UP8tnyUwCseRibmRyweQmqg3IrqGfAUEzcQKvEDeusm7u+5DMTn
9txg10mNY8ku7+43ayRXsO8UtsLWo+aiMgFm5hMvd5HVoC5VNKeuZpg7cs5I
KwhBiOwiyhCyPJ8ki7jRK3gu8jPo8dA+GXP6Iuyh4YZB+qSYFm2X0pqEOcjC
ufpOndrHMRrj7HkeO02IzUbQVdNKEbLe5ZwAFzNSom09DiVAFSSy3RI7tOFf
TUijx5vo/HYsSpG5o0clTXiNMkvmbSUUviSREKucRUhcpwNOSeYmjN35IeDg
0LUZbJj4RXNkRdoLCfcZ2O4DkkYLKS6Ac+KYsrKynBT1QZ3+cVNhVdFG7u3W
oF96iUF0QXLQ8V+5IzXk1Ce+fuFha+ys1E3Sn4PM9GLNkGmjzeIoU8wbgfc4
WHXOblwKx5Rs9LTvmCDjjI1tRMr1Dnp/z0j4rj/if2u+zp+oIdD2YY3sBcov
eeM40AIHi1/zR3o2i50SGfTjwRG3WhCadg8gdLrHgkjCikU5PaxNQRxsLCpg
HvLg4GzcvXYUq0NJJyZJRo5TbYHuZasqRugSxDWR65MXWxE+eNYiF+yJhlGO
t/xt3HjQj7SVFHd8gOI3TpVOYLBYP8M5nsetU+ViGDwio5dWXuQS1KfZ5pUF
tzqdRl/0VRDGdLOn5JDKhT+JCQWwKy9kU6wOZqvXYbKzOn3Rn70tX5ctxTSA
8n42aWSgFYom7+QkXzCca5o2pc1O+WOvYMMMLIwVPytKeYirLOmAjLWt03KU
5LvjldGBeZJl3RiPHDrvOIG1YZgMeYVgRFaAaBIdqe2JuKwAmARHF8wYb1IQ
4+jnliMiXNJaTpdsaYMaZzIFX+elZS6UvAgSEzZPSdj63EhWXimLTk6xCQI5
Kc2nInnKgUCqc1SfbfYULc9xZQRLxZmr88jPgBWJ5kJLkdATjJ2LZ33+/t3v
nIje+sqGLbbDjZy2V3AKJpJ2G7N/hbBTJF5tAnSeNgc91Bs2DLS0AAIFeTS6
qq/T87fXvh+mmK9Z8Zr5f9pRzsKrsi6oGX77/bkoX/deaz6i7NA0rCe2FxtB
IYMZB1XseasSjZvUtT0ZM0+NmtKyaaLzCI4FvFlB/odk9agU6VToywUnxo2s
9FoikRfMQQItGmcSPNmBkE81sKYSjkIeJHpL9nV5rIZQLC9ongttzmAuunsN
GGQZtV9tpg9Diacb9tsStutxZeLd9TWEBPBAjiuO6wEUHijToAbtoDhkHWbk
rTG4fnuBkIlt8yX8vfB3a6E9UOky5eGf2bNMs87aGA5QWHA8zbr7hwQjz6+q
MpXxeTa8fxPxG1OmOSkLJphxWvOEI9VpJAWEqgbVLnYTCP8OhN/McmSdHORe
0qBedAaiAowZeneFOTdOiZKZ6oliaVh2PWyw2miBPC9MhO2pNUdt6cEeAmF8
ZeG7btvH9UhXD0sDaIORJyNmhCBXFJVRUyUJSPjontiVNQffJfpTU7xMCIqw
m8emN9SuxgHvCD7Nri25mt5zc+gcQdXcf50Tof7BAu3vdxxo/Zld6MqZd1RY
ARgHwtJBmXOIYLf1XLGUNW0KktfcEPxXUaeEjb5/YPtu/vRhvHGoH+DW3ARn
JTNLdqbk8H9nR1RPeCrnJ5dnuDg/NTyH8hxqHgmbacaKlvpFpJ2F50WPn5kW
WYXExc3YIrdxQNjXmoaWW84cRTC2D6aFrE0a5sYJ0lyBmgsN00xkTfuuyKlb
RLvZh/I+NcXubsHdU6zhg9fENrmZ065VTkTDoNM6/957gm9iJZzXeFOyc4cP
uvzb5Wz2upivInmnaeQgXrIvvVbL/pI1MQ46TF/6PgV+jOSIJ4NKs0RoQyhH
6xzc1krvyS636iA1dANMB3MA2cIcXbUJhDA813OZhqRabLxMI4/YRKTFXhtI
L2KjolkiIJ9Y+CeuFCer6+5b2wstdDOHMSWtFo3wyOFpk/EjluvRgkUfklHb
hcuoN74WKoZd/eUuzQeP6gQiUNp8BeV8RoC3I3joO9IJHOZRvQQDnO/2AShJ
kGJcNjvyHqihG7CfrABYPkI8ejE5CyHMDAsa7UnfK+mLUTFqdLUiqZLvj8mc
C3cFbnp9IedgGXa+zBb2j81ipMwgx7YLrUM6bImWAuiESAfJSBF37FOGf/ze
Q6adQp2EPtdnFunJnXZxs/CifznV4ppq+DowvASl/seHKy08CDWSRRq9n/GW
GH3BHOHvJrnt3XR71/OrytB49/cRwtFM6l+myBp86Jd9Obh+H/K/1WksA1jX
wCY/INezv4fRiJ1OA7KJtRucDRMnrTPJdssdd934qpikPQ5CIdyO/gKpUOCL
fC8ItOGqh1mX5ixh+PwE/9c5xxQgAIY7yp5JIFBL/33nsV1lJg8PHcwYP/W8
Bovm3z9eKBo9gRJeuZ7wp1DH2y/f6eSqzNHRM7gRKYiszTqsxbSnIT3T5dFc
INxvzxW2tjFLoqjwNm/uU5lQrlCdaQgOGOhDZHzQ0nUKc2bxBZaweFt5AoAZ
hxEwZFnV1kaVRw9lTGgb3/TPEIIPdJosN8pXs5IVO2NuYF2mzKeHAnu6Rvla
L5V2qvZLuq1SWX0VHzUMNWiDCfvE1ISFPv4GVHaxKo+Fpxh5/4IZQza2mnK0
+INXLZJI6CF54o8fayAGHfJIg0dPbwWTn6k1mnTMMYlp9zrHX71f9i5eSF4C
8CJM05LPxcn90nJCzcZ0+F13mnMIwFu0ab/YfQ0lDrFICeeVDVcLwsFAWjba
QjoRsAmX5GLukCfTA8QiBZEhher2QUdhMX/K7Ly406cyDMgccaERLhyxLj8d
5LHgSiTLwzKACUAsStqjBeHraymk8LFRDiHWcg2+btSh1vdhoqHtkDJCy+nm
MXMskk5qudzU659OJEPXPb1gVGEZfGVQxNuH4KSVr0I9ufzXQ2njpBoaV1o1
oZyO+zSbmAxU4YD0ewgsr4mXdwzFNzMiNaP84mfiD7hyrO99Wm8YLwAaNfVO
qa+xsNRQuZXfeM2oyeezsAQlWOF9kU1dk24GuSC3N2w0K+PhX1H8Anz92Bg5
e47gmINyrWZDCnfx3vHkV0BCHmyk/onVWVKXyr7dCA63hpMYWbPyJNQ8elPH
HelBjVRDfUEzbi2r/tSDaX9TLkCLnRKJot3I9kpOXn27VzTdGVpygBAbLXjP
Vk5LbPJvyW3MiUyezB28QVsUsbpqqN0otLX8uNfKdjBpwz4I4ABBOAwZ/ahu
tO8L96HO9Gplu7A6KISrnBnZXxDVagfYdViJS4Z5UMO03tuEbNF8w6AWf/NE
Uncv08AY+U7qEb4/+PPKGPzrOAO1ZBHledWFuh5xzKstKUKHqylPPwXL3Hzm
TjtMpwbzjmk2IfFm71lWtjIAjFHnJa/4IPoBxq0fuVVR386flpzw7HOrIS4d
BjUkWo9v2GrVxDW3Xi8wP3keJMrdkbAgExJy2UVoDlJe76BnFi6QPe6S5xZy
oU98We5S796UlE+ovGHTvgbNuIzWGb6jdIpbSVM8AfM/LvXfvr//xT6/nu0L
9fZ0yxpohvsC0t8OwVY5IBNA8Yo5STD2uzr8jy1qyUUM0qozgWq1giLOADl0
+RTrgVc6rOt+Rsbqw2JlGJ4K8RUiO50iGxUnSdpRJO4iE50JYjjeYMs/OiBF
uGXO2QQB68d2V8SM348D5LzBR5Y89M8UQ4Zq1GcVwmhqgwumCuyBzmneIOTh
r5F0h2VGoJyTibIkfXEdrcVMkBQOGh4tdmuh8Kn27SV/vWC1PpvyzB3Uy+qZ
q+t8dYaYy2WQKjF9Mvjngz52XL43EP+NskFyTXi4jZjmL7KcYyfhpnrtJmI/
G2IBMYqi+60OoKsA3aYISwFmAdJhd8D0SFrpykhBMUedS7SSHNx0f9k+OKyJ
08v6Kc975ktwxX1D20yyRmUhSVbZZWs9qUhq5lJE8JRf1Md3E3HD7A5HfdgJ
5UKSFl7SUOeczBKRSe792iclVaOdkwykyFSqRxtogh+DIKO9W7xQaOOgttop
tC/UJeeq/652nmmGo5vdLl4q/IS42rGCwOts6e+idzXmFYut6THwcsdIlomn
xG8LKe4EHCpQ5Aw2C+Jpj55G7NkOt0H/9y19i+5SYjvbalqg0Aym8NrKmeGG
+dRfyTqcHk2eio/pPLEpHaWWdaT4PDBXPxA2+Md2R5L7z/bxAW2Al2L9f/Ch
r/Alvm8GXCxuOmnEerMGDAQYAcOzMUVvaNWUiPmCPsj71hHeILPGvbG9tbo2
/K4la4hkEPq4S/mFNmkRZHG1Qf82dwfF5temW/pFA00N8BicZqW7LYSPASWn
Rq0L1g6p8gBI2pSCz5X7XkXoCSgDDTA3Ej0t3bAvpYeYeO+j31jXgcX5tQpe
VVtSQmsb2R3tRs0gHVrs85DsxXFWKqe2IAPzsMb2cf5hVtWmEQ2RNfn2a6d2
7CVgklxh2cc7/bbX8uFYRpM3xiK01XSukuukK4NEqePnPcOusaALxyNvGPSp
DlAvE3O8laAL7yxK8S2bzly1OIGMp1SvvBE/ybjOf8KRBu0tA0/jqgJQzvPf
sCCtaN1BDmQ9Axa/J9UKhD9B/YNICfad2GaIrgMGPnL8W43IpyM/hpQoG02D
1goZFXVER8D2ef43dfeZxiTRCkkmrPGRPBHNBpOWAtvHmjy57hTGUwAWt22K
4zZfbPSPlwMZz+b6uMiAWE6LpRIKThsTvKtduSjNnQcQpcnmet9j/hNbuQqP
gmxYKVS0AK5rH+58UbVZFObd0O7CsGcLfzWefOkL2xzzG0wowdqVeSo09Jav
Yf4+rDIw6V9nl8K1GsGxXnbV8kbobZdVqJ8d0hv7pzUw9pT8wxlc9eDOsmUA
EXExJMKZ4iiaulC7/+zfHVH5PV0wdtlmyhggtPGR14oIcqaHVd5WBdTHuB01
/+Vj4dE8bTXMxlQQgrfvXxHHPArn+Z+8/dtkpMH0AGwAKGOdlifaQOVeUSZF
MK2ayw7bOKCwKTdEh0dC7qWVh3AvuvcCEqtXsuoysRtQ9UyyfAj9djxTb8ik
XyCp3YguaxgyhqHN8Yf+yTV6U/W7/XLQsIPT2sX+9u4rEL0wKDAvodVzGvxy
mA2bUTdG/uXFpAlYy6FNbewgPXODt7xCRnHQT9LJhsUIiQkcbNu+nuUy5V4n
kFvRoSrgWFHogwSUH0gPCddD5WpekY586X+M6ZP+n//Wp6WoBX8WF9dM13Pq
YafT22XKijEbyLZ3EDkyApm2Yx7bUTdXQ37WzuvzRuRwOU5mecY0eAmbZIrs
pbPkKYGTQdNj04B+jPJTh5iDQhexGFKAlvu9k/Q2i5EOTVt77a0Ss9Xs16KT
unZG1LirzWIyvaRJ8LCriNQiTu1DrZZIWh6SZVfMBkCLMzH5SkFfSw873U58
6U9cceJ3GlCHsLlh6ctdGLLbN/vrVe2k8SO1rAusUN4SUycVZ5HB4U+s5EKz
IYqrJAbzSkqCVGtGLIxlBrhhmqf5JVMXvds8fBsTVLWqCitpDHmKwSMvgKLW
enDRXNJpaa00RF07h3KmdzRftJlWSlIs28kW4kiTDLAsjOLru7vVYEFtl7Ri
S7M0y6pZMg3AB6vdSXbdbezXMhYhKOQMQYpuozDcLz8pb8xzyChal9rpm9NL
8sGvUQxvQmmEcAFp8H95FWuqdruLRdwtfw91M6YiWFuYbvVRbckXeGm8J3Oe
9tuejOqtf4aJQiYJVb5Uxed1ib9XQEUkL+aORoUolhfqlAahTPCIpc8eiaCj
Xyar8bOdIYf8J7NkHlh3WOY+ws0VJb9hpD+kVGY5D7Qu6OgalNNQGFayHRnU
aLljVg5BwNyjI5zHloFhdpNHTIHDaaTaGq/enjNbNKm+oKQxrSr5IYYCH9lK
4HpeXoACIbbAhwLh8b0bZ2txJobf4YcszEjpGqCxGr5WPAqr5+lPh1sxagPD
gf4R+QvwcITdEPvwKGTcEoL4Mc3+w/IYtzvN/0jlAkFe13HqKcH1+2ol6I+E
nttFOPB0eXn5iycwUOr7WVoscrUtzBX8NlTr1jfKfdwIKyoKxUQ46eNgjbjN
AkcxkJ7sd4W4DcYAfiSa289W0iQITsfEK1hXG54UFYGsVkDieDFSy2rRVQcF
iZ4r5udl/eVDn8ZN30uHIRNNLrsW/PWvQx1ihkYQ0P0eVg+Lq6kCgtptHcck
myPlX3hqiIpJB3c0FVB0sJxoLMCWrT2yyybKzfynLJ4Qmy6zjA0qBDaBDqvX
WPo/5LaH5T0nKgw/zGwmtCRVetGtYfWK15z0oLm0xs8+jUKVQO9TZOEp0H2y
ZSKotcIUBsfpPBBDLDlekFskCPU4xOVOOTJ6tAM/DysQzW4JcRKTPRtFF6g/
3J+WEmi0l16JHxr+Gi4QvK9wmS33dREkg+gylFKVEqQ8LMFwI+NNp2j/EcLw
4djJcrxfQvftaRau7uetmhLZwXdYr7BFqVxmJnf+Eiw66zFkXFRAGe5J1BqL
ZJi+DY5fuwMudJ2OIbm4pZX7qXiLe1hLmn9nsFyXk7NsFgksWofMhzglKwnx
r5VQSvcz3POVJFN0EaMR/fZdnyDfv8bAyQpev0X0CdwKnU90EJ5sFSbaQrz5
mVujzSAslDIyHo8FcEZVyvlACjLJeOUgTQydVr4z6eH3tcS43NQhlMnKVMV1
cHvPrztEtDGKTm1h9aO5RL2pP0u7rBmvMBTTJyXCtbo2g2+AKQ2m2U1rd2OL
B9Aia+22Qy2fGkTtjNK4jWuFNk/ZBX2Rdn5lnrSz1CFzUehXvUNtCjoUKzWO
3ZRLW/zyjmPkdyG/Ux5O2KD3D07xhJQxSu0RCd0S9rEoTRIu9NTgmJd4cfYt
TIznmy4mVs78g/Brf2ohsu1HJLUc8rAfWUfQX/R+d4MTxltggUfuefiFC0o/
CAASP+2ffD7eC4o+O9mnwpwB8i0Wcyq1P0xVFH/vl1gh9vwMwuLXYiG/H+CA
2bGjW6rVUfVuw05EyYOIKSk3ztw1DNpfRTL9ZW4DmTFsCB4e0hL+lyuqxbAI
TbDwAPCF6uFGnaKWdWPZXPOKAlUKdXckIe31aOul3O+FucIbrlTL0ESQJxG+
YlnRRK9w/O3CJKT0iJf3gQFS6N4LY/fkAv3bOdWjn6YKDfMfTTUiM2kAcf2S
2WptiC/D/sQQ5o5f5oSqScyxLc4icdRh5MfNBSgajxkEFHYyrr0a9ay5Ti3R
EbSWs4a09KzFPMTnwoOCBmXmcBl8CAV2GHvyXrhb1ZDZTvZELERmKsE46wdq
vy45jfIsijHJFd3IQ8MDHcM6WYoM4wz8M4KgkE6speh+Sl6EF1sHxIyg0hAa
S2MFHRyvUYfKgzAG75elRD7yl+NmSdfTAB09GaFC+LPdNPa/ugKRcaLw23Nr
mxIDmu6cgmiFaWVqgcnZ8g2R0oupz0OZRL5rOX5aHbUwKgiT0RsB2bPQUIGJ
uf0KaDzMkdW8dICYm0rF3SGuwnrKpVdNduEk6N2ZLysyZEIzYaAF7tZai/KU
sKd+56NOfG8p8imkgnxWW9uNFh/jcgq1ZOwJ7j3gOKKhQvNSp56D0LG7IFbJ
2elK9NR6J7YBSE6vBqX4VvGQxX7VC14KuG2F1FdJshWgZ3OL28wHtlRxE2sz
xYyZaqmEX85cxibMs9zzODZ0TeNKLe0V3z32z9DD0EPwPwXjjwfD8cUbAPT0
jCeK1rm1uWTh7AZmL5dBTWicOJBjNMvorYMivsi4OhQC11QlcMp5wL62apwR
Meaf7M2pykM2pt1OHpXxG16sd5iLhmceEoZRApB90a9Q7HyZ+dYNJvh4WFXX
YO070Jsk4VilCgWc2p0rSBBHUjyFleb6mrxNY6mISUpN+5zh+hTh79wrFex/
qEuXkathGMElrhu5/BWryyPACIBeuoaUILKHgZQWX28eunvzER63C0eri+xj
UtCSgddelTsAD9J4kXTGheKdmNxa1V64JhTXCWbqIJyZV8tjGtmJjuwTL+oT
Jvq6DCwhFLp3djEKOAliPrZHSgkXxuURU5C7y9rifZvuNrHQctDBf9g5idD2
I59L0XzlVDWY3M3MqRLnvUXUPqpj1NTJKJT0iYTBqO5goMQHW8s2AtXZq1BV
UUT1dh2F3HmK4TVs2JrcAqMZaZiN1/4OcvpToyMX6PJaF96AimODGedsO3e1
8hYbjlb4tSa4BEWC/nL3172b/EuqEZlpyImo65f0+D/1couvSql2BrD2l0Y7
3+FzeUKjzTsvZOLua2n7MEzqo8O3a+j7Povcw0necrrHZXvBQAByn4mhRseO
YsuH2kUjyK03pK65hEGuM5VCfI2Xm+BNM68DDGEtpmvmwCMdjzo7g2yYLqEw
/fjSQUIkIA+kp67hUxggqRAxwZEwjMcxmTVpbmyo8PhSF5yvH5K5skXhPvkT
zIkEiV2ILTjgBJlXlxtkBA8fNwRzpTQXDwtHduHbntabQe2uejIlAQImZz1q
e2KTVmXxEOtioSyNWo0BCrWsGyLX+mq7xuIan7ztwXRx0xFz5B15fGKrNmUQ
yg4KrNImK4G8RpE6YcBmfJDRaSkvzUt80b8vYdr9Tiq5deFdA+MBULSrXyz/
8rnL9JqPzBy521WSw4tEHZpaY1vQbVl+IbHVDFAPjjUzPkatFrRIeKXm7Sbv
giN3M6V77GAY8qSo+HjP2N5vMSbbdjjksgXLiGYMEozGpjSWHdksRXZB/4vX
7CsatiMNWdqdJxOJZ/1Pjt7Ozt17RT8SqgPoi31V2xlji2vBJXBsGTJVqW3w
ScZvRb9Hda1KJBkXhNyTLO66nmG251JHnefuYMayAvbUOoBkQjjVHj4c/J+4
yNbDjXiqL6eXHjcF9onRqphEQ8PisM/g9C9o/IJlsPCHeCQO43En9a3w88Dp
8tqKUyzzEO6QWI5zmjI3L0BJDpbhmCybAM6aD2UCumoW3xlEVSsG4idJu485
SRFVd5OBD/pLknjbz/Fnn+F/fcxXc1UCHQn5jbwhd70paMFzD61GO/GFyWuP
SuETpemdmrC63N6yATgF1wDctgK3yhllxyfMsikcKmbTN0zDs3J7f+BJiHiN
2qvVYkY884WYLDqx3ni0mQdI4lmVRl15Jw7+HxvTbVRJ+OCWj3E47eTRWcJ+
n6GOfUeL27Wp01mziwgTW3bAuh9sa1xLwXGRrl3D0ZuiafwxEMQYf3XJUq5l
ixsXIOp2RQIlvBlU5tS57nnNNSXtz6VQFRi8fxKMuvg0CLOZbUdwUKYdSPZF
brU+KH3jcTe35nyxG0bGtFMZUVIJv2DwPU7LaGOSXo0MWF1deCFJBubKesrQ
2V484uZw9TB8rhLco1BKJf5Q/EFGYw4f6lwflM9sstTj5XCBvTHKCR22oDw3
Ue/JTGZyioSTQ8/umd1l7ZkVQtRur9lwoNYn8gsmoj5unZ0GF0URdAdp6+oz
roK1lQ1N9cD38/jpj2ds63fWFXIxvzw2MVZzE35rtSy5BN6Q2LsycVnZ9G/V
bmgTk1b5ZL10Bxaq47oaOg0fKRo5NGiF0mNUO6sAdq1Zir25xZ6sot9Uu2Db
7Y855/jsgspRTwxzECNd29dR/83P23097eGZgwcAq1vtzay8nzrp+2NZ9YBh
olw+MqZpcvmR4Xj4MzeL71KmgYOkte8adr+X0D+49p+TYXjqedwd9RTBX8Mf
R5u7TfHTnvCghkZXCsf+A46S7hlWNpMFRYRWfTU06yW+1owJkMmbbdHDhwiF
ntraIRANTy1Z0MHinEVv+zeB4R9WTCZfRaMAdzQ+T2NzmyqAzH+EA56vh0H0
vD+zq/VQ5RFbZ/4W+rSLugGhD1EpaQG57N+SKEvalZnyCB2MZwZxkP7g+7r0
/zhSNIOrpnR04V5EpJwBTJ6MPbuecLK/l+BqI6lCEYwinKIwN70AhsVdCodU
2JSZghTClOQIPO7S2fV56rvcJNcMYUo/N3eEMmDZhQRq8LskvkQXQZqj/4ly
bWK/LahetcyGLmkTnRAe8ie73389ZrL/GIghexA3NNXvs5Oby4z6CnSBMMGx
MSdoGGuB3VIsNi4u/AygGjtT//DW0bqHuKZApQFpvucCwN3Y5RaJBwxLPDJ8
SXaI9VuNMd6qcoVoALbnENES88tl82j3TOyIo89R9pmPxycfTcUEvslkjQ4h
NGEjEJIJ2A+RCsR3ehHveymu05sBiKCg5F9EpS+g3FLZljOhL2vGqVJLmp+k
gyaFtFpi6C6GiAFnmflSReGzlzySuGJayAyPB55n5oFb5FLRFO8H4V4QHMQ4
BdkloB1bYRpmM9b9dQE2nbyvioyy8iiL9TiYGg0sOeCCY/rQf1d9wV6RaKr8
+AyuB1i49zNL2pp90Up7hwddDWDLL9OuhYd/BpI0vcO04M8bEDfBCgHueFsP
5yhyx0HZP9aTuG/z0heMJH9cbecGbP+/RaixqdN+LPuo3AeMt2kBVIXK7gye
fho8F3TVYTnTTpWLjDhZeL7+g7AYTgNZJStLpgI2tgEuJZoua6iudma+DwmW
oJ8NijsyTJPpm4ab6YX5spvVTF4x7GhRSjzH7g8lCaGKm0xKVnNZuraeuxaR
/JqJMA7CXW2AfQS19ZdE3UofQLczKtqGoQ+12DRROAehBUbEt8GOcKHzXcUE
v/I5pJzOt0NdBSmH1t8hUN9dh4ZHDbGY42NbE/+QEomfo3C+O8Q0kgRcnK6v
HAnEXtyCU/vHZBNr2Yd6yrUqpy9l7Goj720wX7ZzYiD57oZG1TyyK4g9LonZ
z/yuosljUG6szNt+v6sVEM9CxTYI4O6UYmZaE9qoFhuyzvtDjOENjN1crIYj
Xp5YQ2O3K1aDsnro7kacZPTxkcNn7fB9uPb+vJGGAbDo5aNB01JH/NKFfhY6
uldT8EQAzF+R9fPLY8ebnuWlPbQa0I5OIZObjRAOgfjSmiQc29zYXfx5+9pS
OnKlFDB3OARykp1iL02OsrqnjjKZPMxNknecYvpXrC0qa0ivhhW2PHJjQr8H
QfMzL7MQ50rsETH6dQBXlut9+10y9xIzYQBujC1S3TgfA1j6i35zNIN0Epak
cP/x8rJ/YhGgy+EWO4EuTdjLwXijs4Kc75qpQKzc8Plolrs+NorcA1jj/GXg
WbLL3qH0cxLaPU0NDvKY07OVnpAO1b6G9w0O0LTYnsaoBskSSKgNKfUo85Z5
XTfcr92WTSpkMJ8aJmPY87V0u2cWb3mbuhblLl891Gd4G45nBki+oD6CAL1k
6sdZ6VY+d4UP3Bd0aZgXXEu42X+Y5/LpRzoQ9AMQR4dcAajIQaZ6mcrtw3pL
srs1KI/YDiiJ4Df3TtD9/R39USvGOPnsBlksYqCYceb0Eoy+i6K+SFCdYWPy
renAcnfdvWm2sySpexVN4RZACS8yZYoCAGecbugtUEJt4SXtH5AK1FqTt34X
8W57Gis0qd1RMz22cLJ+SOP5ycJtN74fgZbdqn7xNCgr+prL9Cxh6LFrpWJ4
QCEIx/6ApwXpnXi+FQo01Db9YyoD0bZXzzI4HVqfwFwOrUIM4Or4joIhSS+/
xIusIRHwJ63HwHHEcrsRDnO21oF135w/epRGqKecgXZ2g7zMtvcs4GUjT2oS
754yL5jQimpV8+iE/xXTVKfowIC/wHZObaD1XW1lwYcwWgu/RlG3+OW1+tYW
Xbx21HLH+LDMYSn+IRUsAF4iRB0cZpNGmN2m6vtEsrnBwj8WezDqRohlETpa
FnxD6WmPATk2LV9DdGjXUnadyNPdHHYROmLYtxvlnjgd0DlpnHQKBKFZNE2L
nb/0M7HkKMwIPQGatr4gKxy7ACSTSW2XZuS04mzfNCl533nc6EWuvSe6sGgl
B187LORseHbUQVAmg4e8dD4gCyQPL8dkvh4tBzIi3puOrFHJ92/iF4t1EQOv
aIcW69VRNSqHG7L2Y2+4ETUOlC9UugaKKyEQ+JWGv4GcoIdN/gj+/g8Plbgc
mO2r93iuCuR6U4HwkI9gxO2LGR7z+lmz4NaHfMF9NdrLKFRpCdVgdFz6SDzv
ElIUeW1AwfYjieHKBw4b6PJKRP8PrtTrnB/1ktLutyYye2LTkosOM+vwRs/j
wN8MY70OXtJNp0OE8RbZIk9Mj5JlsFh+bnqWdKHOnJdM24M/xPfzYEuaZA6y
3Iz7ZK9HBxFpIpBEaCwrS4rzwCiaispBw3yPdNljFgWhKw/6/ZjqDIFE8O1z
3Q47DuEO5eILTLs1PhFem0JlG77VBT7kM2sMlQ43z9DrvO2WqiyaM+sc+X2u
XhRM9Ex5GoO9N9KWB6yWXP8IhzH0eNLJ8VcOt9ytuLNOqD9k8X+lCMKOLZNg
6GJp8lamnz1Rl9l+/lTA62QBH8ZH+RkU/yN66bqmPLuIuOinyD/cRzF80frV
sNppFtxghLVyNl0vZFLVz/gEPGAcPMm4zhiAgdd/6CbNXzPqE+W1ncTF7VX0
IWPX+9g+pnLrlr6NngaDogA5qjylvXgoiRlmP/e6edQe6K8Jeb8SGjc8ifWz
xQGu3XvqrfolKp/6oRrnOg4C0riBxqJFptkzAoW4eQprKEX0B/l/ZqztwD4l
wb/vTQF5SxuzUa+LAFBkGm3rcJnornGrMlbtg3BT+MLh6vFfPgFNx8u9H6JH
Pgqo6NtX1HSuw1hL5UIoAZGSKAVyj7cxLHa/NCTO4DHp+i+/rms/+Rq1Y+9L
IBwEDP+Wm21W+s7hVUifHUwzZ0Zr2sSjVH/Y87KBcJnd1AF5crRsg1Ov1IYv
2Jubv8oKM1z8uj6aRUgAreJy3f08sIQ8Iqvey+AS6oz5m1UQloup9sFQ3ZNz
taxSV9dwcTz3RRsLOpq0KIikvSADtv2PTqbzCtLw8k2cCkLl6Ilnhpy0aqvC
lAwjMHE0ns3m57EHNJJ1zRJqVSdVBEBkzo30AFtzg+fBthA5UJpzN0gmqk31
hVOXOHfnNuheEWzWpBoL/cVZBm/zlZt6CgFMuJauM/liLWzx3Fbfds4jn3Rm
rqZn+mIWhZTTxlnuafUsLGCjuJZ+A+XvKmQxHwgcKjearirU5Tqvrd0Xwz2I
WE4QZEyb63TJe+zZ/aI+KsoivtLLvXiDyQ7/Y3hvJR07ldijfe4flGpPtqA4
X/gKDB8HiWk8/sf97gGfWGRoX36dTUMujMqjjRtHmP5w6pAwDjo6DzrmvrfL
0KxPQ6BoCIGQzL9XFyNQq3lY3gyxlnZ2BlWbGOYhRHmLWzzR9UbkCHLtijQg
DN9WsPtHMYpwbd478prD3ffaFMe0Qw48xmtduDSqrPQkCUue1hb7AfpBgK4a
1kHs1TanZRebPBBZbdOg9S5ZZzcMRAzq+fdtVD/vWXIRABMkwe6ka5/+03M6
XjxfnTVrnZFvwkQt2Xy3m87G8jDBEsgJPA6wz8G/pQ3uw4zwMwuW4sA1OdA4
wFrvNWeP2d7t0mGddp1vRjKP3JaXRw4lF6hqCmgPXU92c7h12b/Y4ZiRcovb
c7UlEQWyPkt+rgf1NrYjOsACBVioXUd56Utu+mJX/xuJbHmUy2Q/dP9XnDTi
VdrLy/oPNHBsT+pigErU0vdFu+HvQYGMixWr2HpISe323gnw/7l5DkARCF1g
QMcJLRcS/ERAodsE83/WTt5H+IJP64uDknOhnqLaWZsW/9htwVORw3B80ahr
gAkLPZXTEB0cym66zhdV3IB9hQ4845FsU+xSeskxd3H7OvCEm5Z/syt9xg6A
3+Scwn5IoEMOHEu5FtZfsQ8Vr79QH1ZF/8+mkcsdOhj6PCUIHP8H/HSJuIvg
GrgnjoYJCdwePxv/dVCbAQV8jKD8IiGfUdWlA1Ts4HnV7lcjrEE1CaYpEgij
xmMFlp0nskmg9IOIxKVET60denJwVrBMHClzMQ4fSyKcsGhyJw4X+hLe2/w2
aJ4sorKsc4CZzo/288hvqnUhVGi3CxbbySERemhgxaLEDYG7uZBNK3LU9Miq
jqXpo5wh/6SgCXF2xB/+3acbokmbNcAlv2Qxi5nScFHTw5TSLHllMMsIKL6R
BMd17u1wR4CWeiaweE2UWnVR5tc1Sxfafiem2gmJNuDXBIIPKo495cR/TjEk
Vcg1wbWdjSb+7vOEVC7rCytBm5gBviwybdh+mKxkyUNs3TymBfX6zxjLYmu5
Tuhr97O7mV6zpP6sciaEZP/zDn26qQZyCYps+mC6sjra6pcoYl82gAqZBKJB
FFyUl3SDVQxQuxXWy59itkGSE+wyzq1jyzUd2QXLNcyCb8+w+U6R5OwrRiIH
rHhIRjAv3ltx52n8qLpCdXV46jpUNuthIksaPuPqfmpoSuFUVILqJz8hAQHn
rI5ch2dL9VejT/d9MMlZeMbocXGIx7vH4SI3KK/gbX3LgsPsE5Xt0+RPvtj7
KToEr9DD7x5bbuHpZIxw8xKzoO3PV5UtNupnOAkoLGFZLAM6Ox7b70/slygg
JctLDfOOOY+6/R0Dk94KLD1NcVFk32ux1NLRTMiKIw8AAwaoqfk3ed6OnU2P
A1q1kOq7Z1rkyXMkD2/eTJvblTvdICP1o5+R6ymP1hx7qC915CRLtPnixUI6
+zRqXXuaX+YDGR4q7k8iILavm0S7yTjgku69anMGEP1uKx4W0/ELETvuxhmY
0jR/FgPSW9d0bpW7l+g7NmtoqPYesLYVO/PXUmicDsIG9ulSwBtAnoNx12ld
aD4gLDJ1GrNsZjBz/MDJDo59xzhpQvTxaulZXEmhsBTnovMUiyPdc+o46tLX
yZ9mlycizSw8nBFVpwhfSW12mFrdKNocyvdm9TgrHJMuZv1lYuhaKDa1Eq5U
jpGpPZ5DqhCfXKIEo3aAWO1T+3Yi0H79mvia2SgsFptYPofPnlpNY5QiMqm+
nUNJ5oiNrfQPiBKygqesLuNZznKCr1YRZi8PM7bG4lX+KFFllPcPrmTG6hfh
mf9Jf2brbk34SKQc51suidDi0BKYhnQydXdU2YDBhyfnUuo1JDu+pH9N8bYr
lNOsnc+KJhel7rRJKRoypB+dljSeRl1DAuyWanrDgam3X3oJyCkRKFSpdx64
gvobZk0lW2ehdAJojQDAk3qKqS0Np/PvPuYVW+wa2YoH9jrfjkRb/RdiTNsY
hsqPxfdfnPc20DIef/8Qb1/ZuHXN1/AMXgZE8GHl1ij7GdB/f3wxTlJ8WGCP
tG4KV63pQ5C3jl0tVeHFp9sLn20gb78mO2NKqPdp9fCDZCqK72YAqsxIS84h
Kd6R2IBw/woORKAlI3dDAPWkVXkefr8KDN/zwN0ghGGkCnGVH8+1RTGiaRUS
5h3FdRuR6HjAVIC9rBppHdrQdtjRPHstEhyB2rVSGwpRCHxp9AkvAGrTutMI
/f624ioVRbadopZA1ba6Sm8qcRFxIKd9ltBVMn7qg1r8Q3W/2j9hJv/dVY+g
F5SkmkFfPN+GUWQ4pNSucmsTY9hp0V/pv4Pf1l4mrtrBdunUwQh4ziHg31Hy
PofsTY6MXulzVUXzLpy1bWdPoSvLpx1QQNjhbAKr5LOXFgA4QGstXFr2wLhP
QbmEGg1rfVEGUzbwSJyATjk4pYJWOmftZ2dubjjULir/Wh4HcAagdiL8j/S+
3t2J2/1xlD8V7gXW6J7h6BTTz8bAvyxPe7vHKZUrE5OePb4XIgso+4hJPLwk
+05K+6LQfluI5WPoQbu22Pqpg/jKuxbP+ePx5xb6sa3b0WlX1s04KmlbVFo1
9ifFyX/H6a1lGEqMiTkjothZDg1cTCRcKc9DZjyGMbSspn8jhCgqVfcJvpRG
9Nooaaoo/VG/Y+ajsVLE61dGuMJcTeXFY3ShpmtylhE1lPke3RpTwE/vugyH
XjKbA2JfQQ9gTFexKvivvS3cYYFJFNOMW7RnrxTPS57pmtlhI5KKP1uPuMOG
4NiLASRh4+1/bqFscaLcpvbmWKelaazbx+zp2iZVfTAqPF08KpNehsI4prcz
jfjbq0Rr2bML/QY/lfpahv99sf1qZnzrs/TzxeXpPtY5i/oiNxRHwgyuyXky
9KuYB0t+oeSqGDa8RnJ53i4lqrS4aL/duFAJ8ZBAI/3UILw/F2xnxt9aO7SN
OfpG8AzPMFSIkigD+5YpH3Xp1CzCmt70KN6m56nOvaLuNQyN6iyjU1PCwr/7
08V+DoskgHWcgu2+wG631K5oRY+J4clfgup/g6fo9Ppawm7UeUTOUSqh2jSy
b0yF1OEUBIQHVfL1BfK2D/PVBILdPnLt+MES37jwHUbZ1MHhsgPBAUNbt7Jb
hxNdVwiKBGt7/bKCX44/OK3ku1edRGX4jbsSeeRMe5nyoq4q9JzwGjGWnVB9
z8tsny83qmwZibRSsg+aYw5HwRgHMTBBC++mw9z1LX+vYoQD/7KDQV+DR7t+
FHVaY1pm2N8hm+LUegcvC+6Txgmm34E/ozFXIxRIjkMPjEh/2EBmeOqSjxV4
7QLcpzPX3wIb93T5DKzcOjeTul+L4YmawWhbV0kRWLNzDuJKK9BcYR/T7Kei
DOv5FZkgPBWlJOfyueMBam1k5+YNi+z2L2LNmF2df8C769/ycesG2pPt6K53
V9AGPBUaM5XqxhPaIPm9OVM/O12OwJJQsM0JSzyhfmvuGIaY3pBzpehXseIV
7+SnW1AwTGYEPK701+glRpk3Kw+Tf7fk56mRcA/u87fpKjdStAk2wbSMNz9U
gfzkEfqTAAFb2YpAT0oHKq9PehdEud1CdIJJ7xX2SppqaOShaLfidGcm1F4B
UiiXp7+zOu8tLe+cuQ2eJc6ISFrEERSQqnv317iXsjGQ+qTqdNwD19G8S3nt
+LZ1InLadQzVJ/OnEFCTOedbwnhx7ld3RLsjlIQ7qfOOpMLCR+HfuvDDQjRS
bI3CJh//eRLsoEo5o5lCoux4y0eVCA0S/590hYikJDeFxrS+OQ738dxa5se2
ODPu6asmHOByBg7BZlNtwYrZbSWglul0L5ug6Q4VX92Mrh57s3VMM/kp6Txt
OftDNjyAg8HCVJCDRcG6BBJj6AOo6abjjZFVpq6GNqoTRykfjRxLp+1Uu2RO
dbtdIWgUS8R+kxDNdL3Z3YSqsK82ix9acFhtZLgjC248F+rklkzRPcKx2n/u
kXGpojIhRKhlAmRtS/uCOYLOcCsRcYATPRxYfQVumhh5fwyFC4UvPDEeeew1
ZcP3Tja3RTIblHC1t7HP/wFUqn0DtAOXM5LDRyZsxIWewLO0sWMb4Az82wc/
LR9xk53UgPSRwE0sM61DcWGvKcNiR8JapxhHkuzc+2/CoGJPlLfe9oJol0N5
JTctYEv3KKP0IvbUcO3jBtBFDYcHtrDkZ38+9qWTAexlSeHsJ4pj4lXTnIRj
d+fjJQzHxwz1XQ1+QcQ+2dcTe/PZveT9nt0tRxbU80ZAtoI6UAvMvo7rQIdB
UN/ORM/34h4XIE34ki+3k7GdUlICI6SHOf56hCZxbDDwdKWPwayURWEHoLyV
kvXUEy9hk4I4pkE14MVWjlDHEbBD6THJbWY1xWheEJcpCH3Viu2VtCKKBvQf
CpEpzj4V1SpM0AZ2OJ0gdNIopxG5vys/wDkA2u4ySY3zm0YjuHkVOumKmOvD
IQjxguUpWWEeWWI9ExPCqgDxkkCHHcotOkE7w6+kQ7kUIthcOe8feeek5Pg4
qtmD+yEygaZSgjkfWQjl0ePfFU5Fni6qmGAYngFjPyHswWQAy6BoD8tEosXG
ySQaLP5vxwToWlvgaxhCRcoa/aastt4X06T+1BOtAVOE1q36+fDStTW0f2tD
mFhYgHgCHHhnGlSPxU3KKaYHp/LE7SZt4lOfSpqSdwFftTWqcZdYZcpclKnB
hx1C4F8erFTp9wUeLe5pZu9VwvbdVASg1Z51eZ8DgcKK1mir8qBQYVleEU3i
iGrObcJji0aSQqJEAlSQa6pqggEYnoMl3MvDf8xlCiu2NxuLwiZt6oSg3ZQN
0s1JbMRritdBP6F9FGSahk7XVOBnTIwUD0ZLiWg4Gk/v+x4v9buQ23ol/fqt
+TNlOphKXoqtDh2BxuZp2T4CEe6e+P/gDaVxvuFfPsvsVcYksuN/Yxk6qkN2
euh4eLaSHKFpqQbbapXy4M66/Oo0PCiVQgDA5J6fb8f5qB1aYZ5KBYltYTR/
yI+l5jtIE0EEhzMfQmVRr0SnLLLcZF2xAD9LWbJ0Jg38qphFlcgruWWovyAX
O5gBRaeOAxkelW3+cT+aCu/JwofrRgXvHgPdBzgeIeVVkJSIwuh5VN644lND
qcviOIRBjJs0zf+C1cBhk+iwrfoR8mbg0Z3LIhXVYu7K/wY4fJePLFLtMZCR
u02Rbd+6WE77DfB+QKaDcQY5JcVV8cecjPMlNcRdk2+ijSh8nfjrW8eQbsVY
M58UYgWVK2dVW3Y5C9ucsHCM0rmLMXXa6sOi0Rkf8niBziN5s2RiDHN0S81f
rG3SGTrQaJhR4OiqplhmK1VIm1JtyFnZwWnLSZ8/nxbCzWOZ4wBS9D0LzdWx
cohR1EoyRYG8W7OosauuyMkpc9g1uOJbN8tTQiEhjwo1F8NY8preYzDIAqnO
vfkXRH1ePOs7QM2C/PLtlXeyg+oCmggZoZIwC9CGVDJybTmWrbooHtVLuYxr
agade6VGZXvpNEr84w4QlW3zKzMep69ZuyVz/PghJPyl0r1rtnqOJhW8LP7E
ZtFm4BzeJwvKkAA6y/d3HyrAncAmXYXrx29af7SkOXuS6yyd/o/DHm6T82ei
5W78dr7u7998oBGB2F9nJ1Bd5bgkQz2VPvFSF4OBYOJMs0yjoYBTVgtfWm1T
0iz354h89TCmvINZRicfG4pYLMQo4TGHxde81hDT2s1RHVoA2kAPyvDRJ++X
YIANRzxT7VK8X3yoC8mReL4PzbUOGriVbY+v1f9mhIroZaJ9Ns8cfiwsX+QQ
t8oeaxrJBfopDi84ruEgEAC3U5Oa2SS+1FGi12xGUk8aYNvtP5H73L3V7FoL
VW2HVWOcrZgeQivL+wmojQ3I1XYGAaHOf0GYbEJ7XnMYzQXdGD8th8ZNlV6e
N6cxcSNrLTFYoSNP1UHGASNjy6RQuSl8JnJY+DOn9P9MimhIIGd8SEWUdmFU
AYeUBrJ8QdTHTF519l0mhnpk1WZs730MJBbioAqp9+BC2wQVdwjpeRTSjtRN
Rt+ycwv8/0IVk/u3NIS8DbhE6S74SoPPPpT9DdVjTD8i4bXp/PEyi0VWPdbD
GocpzDgEDk/hmyO/mxzrjBYW5+zUOFNjiOznCTWNJlYqVN2aNmbptmwV2933
1qRXylyRsPTuVUiyo7NfxqYboo6L5Ye+rtc4esgHbay8wGOJndorgwv8lTis
wgujdpT4N+YlxNPQPVetQoL6iz5jjNQTX0SXVDjqIYAXCsOvu++MmCxHDbVe
9OH5lFHYR8S2/6mSh4KrIf+tpgUjJUT9PGPdALeUSGOdqtQ+n9xQIEisHX7a
wyA4DP+ass4434GxrYKVPUocMao/eIZd9CjFmVUFaB5/JduTa2H/dRMRbuTK
g38m5mJSzXtuPFRyCsPqU0blv1QkGJ76dTNxVVCQ4H/TQVISAFX8Voqekqgq
mdbNGq/bc4lbFlviv714dl82iVG5g8XHO70uo2C5uBL+PqBrawTqv+12CjSs
G+t/ZIt3xU2ZBh01wxTN7l//euvs4PgVvQ5JJrYEAE6soUpMRzgoR8UaqROX
8LPDEirwBXZLOh0SkKuwznHCGTi7cdp5pghjXo1uFVB6crsyfvB+7YJIcznE
zxDEBIqpf5+AzWOPMcS08rra0lSEwabBEg21kriFYn4U31WUBeM19bkT+2Q5
xHuQTcp+GF1pIv4CNLvWz+HeNgK1HKGPjhIC2wVFFZ1L/gZN5ZUbKL9KAfhP
kqOziOd1q5HQbOd5EWDAjMRu0FNVN5otrFkF1NIpjG0VaVG/YxsQbqnb2MWV
wu+YwgbqpwNkLj8y6IrGLNCbkIy8HFzd2a+YhslQDPieUd3YNqhcV1ZLaFJk
GOwaWa53kq07LcX+WxLps5G0IiLibjlKlJdEMuHEVI0zhaMETWwCh7QVOTcR
m4OesA+oXvQLSvsFkx2vVF9jav6BzLepTvb6ESIn+HlK7HUqH0jMhCpEqxO2
aHUBWzvdcwwdPSxAe1KaOLFieQJGLlvqzC2Yh9KeU4u+8i1a/9KhRj4Thtcr
PpxE7cCjqB0+v3OPfcmtfqKU5Zkn4PuCVvZa+88DKV2XiEyvXkgpGPGUBCUF
4POQSJgynRWjmoR9r7SX4IfCD6HJQbk79EuftOYwnit1iDd0DBS/QjU1gJs3
rz/UdHetAq8x9oZSSErZSHEN3GLVJvsAXOKNYlNdIrxpuLshInBg3fD98x+C
/S/zlwZw8Tzap1MV+zu5VgeuVRdpMQblvRiSzx1cErfHTRp6UYZCu/ZRcasI
wIeJsgelT4ltZbGuntOfpK56vt3/8kJqGGawZ01tmiyLiZ5763l2ngwy/OcO
DJkE/A9ZjGCXzyyathmaSS560moXKqKn9rW/0sbmQAs7oz6qs86yLNGQsvL4
X9it3bL6/y0QbPh6xcBvuz24IfO+0+rT8OUy9oTGaKr9UlD+3cPZYuN8K5UD
ul18LmdQiy8VFPf58nZFyBOQXahrdgLjQAR/vZ2YJkKS5IKT5wJ2xEHbLfc+
+mk2X2EWKMQ1i/wc1J1XX6i0MIFbokdhJZC8upXVWVZks5x+yG92cHZFVl0V
C64woITVG4dCgi13KJlmMb8b1nsyiZrwNAs0OAJRiveiduvn7nYOv6rmSqnY
lgS317NdcfaACHAJn6Po6xl3w7U5KvFyAhPOQPCG2bS8yoTiOoFMT/6pDGpC
865Oani4D0ahmVS8YcTS+oAodiqOsqzoAfrw0t5mD7QcdtKUneMeFWLFaExA
nHuFLXNRR+L67KsfmAnMg1Eif/wkleDU8x2uy2SAH25srLnkvd8J+n1WtvzS
Rd6skSF1zknDk9VcgO/t4sBDlfcW9NEfxgNG6zqMSSmAtTJPJFtuw49ZN/hY
4SehaSLSzIPwTJ1VKQ40VKPa3nF3Hc5Ja1LRXxpgeBh1cd4938s7/oTC3AWg
mCgF7vVLXIahumQeq3p43sVErw56fIUoyhMbbPmGDFbmehO6z6rEBUttmnHs
FSI6+vu1m6rvdlKdVCXTExMMOOS4TkcN7hakIyNr+LVaMhXV/7sAEtDB9a+X
cEndEQ+7L+/udsxiIQvIIGcwTQ7HC8eNbeV5FUre8e1p5p/CC2BAhnniys3R
xwWsDtNipocqOZxlqzX9Q7s6wEZiVwzIxprUjQ0kRYodvwWEsmB7QCsF9uik
IqDVbCKm8z3b1wulmzYGlD9+9vENCePQRmytZoxgfUVtQZBaf5ACzVmNVOmv
EPMgmYvvWum20fTXZjlA5lp4Gjhmq2JstLyyoRUv4/9AMfM1gE/YTAM8EyNg
+O2txKJW87LUYNxiY7RIPpx/e1cN0c8YXJnA58UweJxDK5W/s6Ssfur9scgS
SGvSTR3L4fImH8LTGi0YVymOorkk+otZ5BEvOKZTR06LXleUs3E1Rmnv7orH
+pTFnhng6zyChUrO/aejA63d5N6caGVCqAnngFu2zrxS+ELVihJVLp9ovBZE
tUG2JMzWE6wEN8t+bCTQFi0ZwPbRHjQb5SHWCR6rKHPxBLfnbK1fDSxQ/dJJ
fHciht27qiXgal5Fdjndx3M5ZPiyn/kb5oabIk9FanI8rBkNdbjXp5JvCI1H
02mdPvqveS4oi1/sqqnID1S1paHA21JXIYQKcdy4Dnt4DMgmREuWgIyVOkGh
xVJTdGb86i8UmB9249/F9F3jab/iu9mU9xEU0SraXABEYVTyKku8Sqnlrz7l
qcq/mTV4t+8fICeIV6yglx3AWpq48KykfJUWJ+j/SLvmB2gfNfK9rAofnMGj
XvjRxalnyfV/xAMs3BWTZN51hC8EdWuQFywFhNpQLmDuPW9+TtiW3rXpx2Hh
noayS/awchHujfOlw8Gn4d/RMJhhbWO0pIgObRRLdqq0+a7Hq+CJ0mt0M2si
yGYtBDa+mARSu23wPK+K0BMZwVCHhMdb+Z3SO3tKGGIDu4S2hMyRmBFTR47X
Hh7Kqt+iGr2lKAzRj4G7UuoaV2Pt67+l4WQjZutOF06WrLF5lpdW2vD0RDae
og/+ReH7VynzAS8yN263RUz7pznDFeKZLhzksziCdZxSluQ4uVk3QMzcXVXJ
nr7nbmQC8/hlQC8SVdzN1pPbFHlwkWoF+JcP7PTCicfts72OGBqlT9/ljf2j
SF4UYwmZd9u4ad/ngGeUDO+JNG74FJwYvpwd7BTCk2GxMrKtRcC5HUVbbTAF
iUkfdTwQl3gI79eCImMk4wn4S1EZepRzmvVRQW4kSOM4F5oGMrICUWXgSJXi
wDV82ua+C7rgGMAR3P4lg4U/APMibulEjFegVt+Z0RSwV6xhkI8UwnkZZIQl
1cvBoNnX7U3ENmHGsV8aDU+p5xrl/mAWn1k0pL7uOMGULuxiKOceUqeG+yPI
cfM8kWQ9OI3F2j40eXeKPL0PklENGILEYiEjbplsijVwQ2KRbiHgtHKA3Ycl
aepmzS0lrn8GXmPETA91MB0PjS6iI4RY68G0EEmMoSOGqG55fzYtRWc1UrLM
tILOrN5p7M9pLpA49eevDXA2yGJH5FLxqEpYbnJF/qzSZjdS4okrE7mBls2A
SM+bxwh5vouGLJirt9FYrgqLWyVpFUxWXLWDJkb9q2oqTQsUZR2AIXndy1sA
vAMTyQTG82WRqOTfafpH0LGqTkj7UmdasfcNcnxiUqONq2ANS/yb9CdH075j
e8CqSobmh8mX5cqxmIznGu83D1Jm1Gh5cr5bBOuh9IFNaIinLK42BkZZlhWZ
lpxeOTd7xCNZQ0mh0YhIdheuLdgJLvv+2v1bSrv49At5VrPwHw3dgFFRGi+S
d8aRkzuXJl89pUZXeHlvfpi/B9ylHirg8MMWMnVzCNd97i+KHRiUMkljVAyM
yBA8yA5B2ABgoBCasS0xCvGhMsUqR2QoS60xvQ9yhd8+wQu46zWuAljX6DMa
qWT8ap/3g3WJy5U9mEZEeKHb3cME1FUhDXikVTB8oK2aqb1oESQXA9KdtQ2b
/NmUgcM1r8CzUX4VYnCNq1KlVi5sP8as67IAQXwB/G3IUNTyNjDckjLYlOpT
qXQnqygCt3i3DCa9BwcK2fSSoOcFdSqkhNpTFwKozKaSAdIVWswHVRTwhMDK
CxsLa6SsZGSRAGIWnzkHpnyg5MZukSLze5lrJGBANv6QNXvis1+es2r7leYi
HzewoCpLGFVnIF7x+b2jz6zCid0PttSoyrFis1dU4yYu982Q+xywW5DrZWHQ
A7UPs05v6JL6E8qROXW94LxD7QfBIARJL34dVpu87S8KBRec8d57CqbbF/a5
xVgKAuySp16354l0EFgTpnsAtK9O6npP3aGFo/5aoy7O3z/bKyBCOM87ujTF
rM/4eIZaKf3TzIi/q5k5B6VpjztsGFrTl1pTWK6dQQYvhEvV6kCoeB0u/tyb
UpFLpEc6zBELZdFN77MQJ2KOi23wGPCEEt2RXQl7n5eZcqwEYIle8lOH2PYb
f4XreVGGWzv4ZaY6B6zf17tdYzFEuV3SqIK3661Bt3goNeKqfEPDWESZmtyt
ml9smuGfqkDl5ykgZW9v5w4nkyvsx7AUuXh8i8w7UEaIwPnPASk6ZhN4HwSP
xPUPYZ2ByT73vrzQQaueIltfx/3h/9ySURxtJsGrb9cmIKpokZqx4NHvQJ1K
Xy540etyKXUMWRg5UdcVzBgPgWQ/OJSDGgW7AxK6Pkg8CTS4zJD04ilRSs2Q
gZ0ljsCJKILrU6JctIZNT/U7Zw5rnkNLdxr21wArPMR4KaWTa3fJ6T6KhhAR
OBCHpjJU7gBxHNVp2JTGblWC/ib05YxPtXc+qD8PyBE+I+dKYR90IHKI2aHT
2OPA08Yt69W8hVHJdfvqKfsTOIxBo06AYy2Bz1VkzmYjQ8pOD2MGLLD60dzO
EDIp77f2qEKHBB3T/qAjvvglDvpFq1v2YtK/McCv0iRExD2QOLe5OSDk7wIn
2yAwt5eLKlYBCtSqGtTMK/m7lJAEioG+KAe4EmV9y1eQpBTroLc0S8KdMgbs
gMDHGfbxk51qfWJUszTlgzz+RIwXtAE6NZxYNtQ/yY7tMaM3gAb4GL9A0+u0
ycR1Xscfd1MESGke9RviO+HQwVDicthUSacOCm34/L1w3VHorJfR4lb7vUQZ
wfWD5JTB9rQ81v1bqZRPUe39EBXLCEqyuewflFl+P0cOYDRZmzn1myDnf8Sv
rCmFPxj7QKFy/En1FqGop0i++H83Rzlm9PJd79R6ZSR38vOTjUGIK+TLOWkU
ORB5T0ijqRW4HbAhNhk9Y7Ir64OOE2DboFssoXJ82DNkmXEeyZHP4bxe5lGj
pKB0SQX7hXfVNEJlYMdiLspRKJNcR9yMHy10dScMdKPMO/Zhe1NFToVfm8SV
LWiLeG85LNwn/XoH5RkGCLyDOi3kj7Mb9mNQf++Bx9in/TfKTwXbRS14PHgp
hOsmi1SjaigrNe6wBcBz8ejfGWzq+I7fguo24IdJeDLMRsPDEdX1HmiUMOw1
M7vqmr/LfqMhFg0nCtfvxgeFFwNAiDA3993yKQb3NlPrNcAyacEBTL5GDvcU
HEBhKVggBRBIf5sVTDdYfNCG90gnEIIuvsCMzKuYkrti17pgQxdXPLxW6m1q
mDqgtDKNoBHMGGevObDEUcx5GKhe9L56OsRxWwaeDGWzp1alSnEg1NTMwFDa
/3flCdTu0JFJ/Qq1aSVfDjIAFX2HZL3g57CiHHEWk4tsWT1ONZ/+WQHtzJzk
BuU/9xtJ3z1Koo0aVyZlpoMCmRcKGKR+TiCOQz+kE+OGwn8P94iG9Syefvt7
sxr0g4EjchzFgtCvRdkbYxnEpqFQw4lrL1ASc783uoNsSbh6kzS1VgXrJ0eE
Oa8SZJQPPyOF1MQ4vVrp7WOhPZov/vTZnOU2ubl7nGSQ2BuXlRSIgJhovs78
G2W4QMDstZWwHu69h6lr96ZGupeMqnqdlte5C3m2njcEzzq8DAeIqeJMvT7w
AHUXUoB4sQkK3NtiNuQJfr9Hgvc4kzWmAEjlYnWP0BJN/rKTBWOUYIwDchoT
BbJeoHsgsZM30tc1g1FiwP9e/y4Z1U9IITb1HhdV45B7fLj/BnaeT8eDH//8
n8RXqGLYwIp9m9nQenHuDi0wI/xeLyGMajjYJRBvZtt6e9AueF08/YAwIvMo
q3YUrGn86HyFvPjJ6vJpr4tZrJSPBUfHdWpItSN3FPuQsECMev3DBEXJZKd9
HKFdoVomTn1DCRLWr3avIRNoI9vJNAsNCfUCbQROQKqku6pTvUUYwo2KFpdQ
SxGol0JP6umhxAyaO+DQbBUUXiMe2YJdK8m+R+9UdzTNcSuwCYWQBPV+IHpj
b4fTJdOC5fbMtLx8OOShh/vNihWwwwjkfxOXwQMfXUSXfbj9jGEiu50Uawjj
iusK1H8ZF5XExKY/TWNLHTZg2sS0m96ougp31cTjqu3nAGlbeiiXF8K5LHg9
HpErQ5dIGAoulVEIQHteuZLct0oPS7K3JghbhlFUqj2sLzckigLpgWQiGIY7
IRoa1N+iMeXCgnwpHv9wcNw47EirC2fT8e93dGyFSeaVwSXcWuEgStNrDKca
hCU0ow7N2L6tGjxQb4KT0375iULw987LodpF6+CBDHht04ZgwPhCDgjj/cBl
sT2lNMWNecHQRbfy3cs5+AcKkeeQHMtWAdla+fpchskb/kupZFkCKXlI56j1
+kLglyw1pkzFvd0ceAvAasqzWHL0ebG22Jzd0EvqdfFreekLokkwPle+FkBC
BXzV7KXx4y5Y/OyTgd2UdgJkd++pTsvCbzk9SpWGvLdLztapzCJhYSRMCSeq
S/sEWg8Axtc5wIl1eojhvCPHmj/96LPd9pIDyLv2wPBH2hvM0WiClCD5TIHw
AxTmQfYHFxH6zr2WmpJuZy6M5FcDzsjfYJ2Z6YF5A6GFCFRSBXsFMg1h2/m2
qsZbI1JrHACFYzNU8ulrrT9TPdLSSqve2JcIVJi6tUfN+nfN5myxzETI5t9f
6xNZaQuRPRbK9WhFuvDxQbeeuV4mmv/a43YwAp9C3swpMHeeQg25saBMvtyi
ePynafWcebr1cw0nJswV68jljQyGCsg1LafFdbeyPXOjlMmcWAQypzAZfUR1
Kyk/iWSRLz0FA4/XzNTn8CVlWVOJImDZ1bq9GHvI6OnGCUF+7cgI4//cou2Y
5RbjbJoIpq9KYpr10S/ZqLKXPQrnjP9ara8ivYs9XMIHpP+iOc3L7etd7xkr
dlJt7vwl+9UCm5ctbnjiHgsdDcRzGGa4lc29gcN7/JvnHfLe9HLgiNFw0ZQK
QCkaG1vCgaYXzPA8kSE+PiOHdWJfxAmgByjXx21Tbk5pTX6H+7TyVfMoS3ov
WcpgF92CpqXe1lxizgIAiEXYIRwNtUn3cytyPaHQ3sahpc2VbpWdAMKZY2jA
TCyuKuGQbCNYrJTro5Tv1P52ntBywKMaJB3uHLG1oZJXURGJMQfS1UqWvTKZ
CoLbJ1pEau0mgcbs54t2Z7Hu/ahcgZXC1vEeyLNEjorYEbWLnybfgpy6jwKZ
uoJltH1fgoMYGAc9adupxbtwcOFJ5T3O0i3oa6UFW4myVkLTocMf7EzwrprP
Zj0XDub2Dq7gLZCOMIf545nAeehmfUDJuoMsL8Ln9FVgFxJqgaNwiUej+JVp
2zx7ApYEd9+VEa4koCKltEa2NTDIWJe6zm51ikyM9WfzhYRqlL6UpphM0g5T
azH6W0zVv9Y99B+jrtDQdqYdD8sZEy7diagoFjFh/243ljD1CLZnzq5sc3YO
HCcCQy1UwdWhc0U3DWQvLO1+FPy4bb3iW69Gcnz2Db+EB8OGbo4RB1AbbmfW
hJ2ptWHtJJ1u2agsOW3jwCS25DsMUI23Jcb4hjj2Sx0fEuqnLl/smb9C+jIg
1MARFwnUQZfDf4tmaJ7PbrxEV7dxdiOK0yYTUPnqh8gUqpQDm8HDdpvGB7iG
Cjtt6b7Xo39vptSA7zF+P6ssfJWyxCCi2cSmEEuYRIAuKetbBFMRmirV+Xqt
5Bu8cglhOsUD5AfLZP5rLspDHw3sRNpUA57llqmuh+az6dYk+y0h0Rho8+Us
ZIckmJSkQyQPqIYzO0LQcWOJI/NvIUCBgkd0NRoF7TJRJBHLBYijXXiZDHgO
bqbHzxIeIyG2OC8pqJbpE5Tzg7EArtBYPQ9AYY8VRwnNxnvqjhSmVRtZASif
gOO7/YG968QfTy+QUUPceOTRHc/4e+lw+aRmyoDFVXyOrY50PqE/j9ap3Zc8
8olXTARDVidGmsjKtDb97k3jF5HyKS6rtfmMPC27AW8eS3yLKa48+QsJYm4v
owpGcHbckg7yRugjVxZB2+t6zO3mmva/ae75dSMLiUyH9dwSPU5J667pE976
4nnsF9IlkJ7yEkh4WuCSnv4RFs2tHiFGCFn+B/gqCXrwrUtgna+fkY4cI+JL
xjdshQJfSYBbouPNDtwke2yv3woDW1X0Vo0a3/NrsTyfzcq4Nc7KK7j/ViJZ
ekRiFuwIpGvPUbmA7l2OXLUbEsSTFzWKBzEOoNXxzbaVE0G//kSHH7dUen/i
fs4vd3A1kl+APuMwrTZIVHqSRGIeT0tVQ/oaB88+/kXEx6qkJ3u+xL6eWV9S
uXOvKreFp1ZkWKHbrgDZVbF3b2uaxoVJaaKH0/TFPKDa7WGDkVavXacuAXNK
yizhmp42BQyuCA0WyWy9hFxIZS1qFKqp5kZywpTfx5C5AtT95bGv1Eo1hTBW
4HKb4HCNAjCJsQWhmE1gcjUxN+xWuOTK1mutjcqjG/i3FkEJYvCz/zJWrsCA
gCafd0ZMkIG3nBqeE4wrjqYeALy55q06k0y2MXc890j7Q1cUdHnD1xS6HFsV
KnZB/eC2VKhPlvHa9B/v2eO+WUKEWL2vRguNAa5LnpOiXGWI+oKN4qSuXna/
vUeKyxakkGTNRTKBZznSiN/zvno6sivFjCgMazUKWSWgAZCnN3mK3lkaM/Nk
WkaXOmNTRPqQ9s/PVb+saGXowCV5K6eybTvHO+Pd0EbaUAm5zDurjxmOt533
vQCV3h+bWgwuU+D4+sNWIP9UxQggC610bP828tifqY+7KKrt7ahJrpKUIwYv
jqakZsYEpqLkSJncN/xzAQBscObXtG9Ovwbv5BLQnrVqvX4PkPPqRlTN51Jj
uwAI9CFgy7OQ47fl2eJjhGLQ/ZcTtn/J9wBLhWMc1qbawtUCsyZhYlz1RxXR
kihoruZx0wzVfgT81bh9XctjROAdli1aMfbt5wgJnQhKu8GONrvdwbwzX7/k
CZBhtZvVqxx8Ml0HzAIIMOuy7/Gg2TRV6h/C5uqzeOj6We7mQGUjNU+QLRV4
A7twZHJFbnRgZtaieI+0M4BKGQxM9NOOYxbjyX4EjJ97tOkDvstwaIDSET2J
DpYxS+snoV7ywc6bmeCMFXmw6SHrW9UBs/ZqACK8oBSgnMaP5/dNrj9f7rSq
l6Gal8fXfQjwXqHSAO4Yeb2+tF4GGk4P3sUN5JFTnQRnhcFhM2xMlVaIlpM8
z540UGHGs9/BokxIIaepKKZ5Irk6IE3YMkxFm0BHdcFPEJ9Uu5Tdrs41d1mp
wzbKkmo0Qhjup6Z91JXnLFNlofu0iZZlm9iNfq1nNB37HV5ivw/6ud/SaWGO
61k5htFfCYxUGMoJj5jvFfcMnotdE1kL9QLo3GZm8oG2MWdK8G2VtRLEvacA
WPvKwYIMMcU/R0GK7hIQ7WukK9O15EIt8qzQtm5qztm51rOMPN4TMb5WdFk5
e2FJe5uY6rpf4ds8SzWUUBJcwaQaS1mlv6zujK3zilsGYCylctnO+3A+jXIG
sxUkE6TXvMcBj5EmhK9YzOSIOLga8VejXzwadOgNHyarzOOREtNvgMe6FcAR
E1Z/YSrrFY1BBq5RbX5TccKh16AahJcr8RiZhzyL7smMHSI2IseUW+g0VHgO
FDEbpBNlQscdMS21qAB2Ov6hkmu7UGvIw66/k0FqB2lYsHQeaa37GNfIZ1EF
UFYoMaplSmv6WX5x/CIGTZ+IutQ1WgsxH1SdTl1WSK/kPlJ+vJl51z/qEs0E
4KOaS0WgFO062jt4Se4eOiMCF6+rDTb/xGITwvG9d7WsAqvEfhdOEEdIGyLJ
qAOhPhbXjL7FWndtLvA6XYfTUZUv9xx1NaMZ/uBDOIWnehNwT+y0GXh4T6zN
TtWTK2AlOE6KchMZd/pXtzBvg8LKIjLe+eBuIJyUW0EWCNuyxUnTQ8IzPLjK
mNzZkK1NXjBifvVWjSao/eVhk3iV9EoIajDLGarpULYwGFinSiIy/qYdDs29
9Dn1LHTWWqd4e7gM5FX0egguTnBlMh5pYAfRd05XgK1b+W46/YrmmHvXfrmn
FvpC6bAppQNpOn26k8wvKeL61A4ab1jgo5xPlzXHw7DGip+yycs7iQRY0rxS
g4D7i5gpRKheTeP2YwJUscikFS/1BGUpj14GyfQ/aVmJQ1HKUHYJY9I+s6Y4
K8YFmMbHJkS1aczKdlVX7Sjj6eQCNpHh3oW09JEpTQfLlimjr0hekgRn/Ewp
dXsKdBTXKQFsQp9jk9UBXjfFwi6hqbiusxA5ZmP+KFQTlgeGNHqTRr6hyYb7
mvkdMRIoLgRdoZFy7Ju9jojvSvPMFmMwh4dqcjZ0nR5xzeIxTDKsKBtaGb44
PTGAspm2ZijnPq23O4Vx/ooBl/HNP6/bd1u1f2OQ4dSET9MZG9BTv2hYme4X
B8JF33hWm4vleInL5ul5G7e/wiVDYw6HZJCWy9x5T4PXefkjYo855jY7Kusb
7430FHtuSDeinEvuvv6TiVzJatu99D8FVRmUQ3PaNmA2D6+lAmjJ+l/NVegj
n9n2Glc6xBdjqDTmjQmXYfXQ4mTJ74DHeoCO0bOigaFBb2DZt9WO7Lc04DoY
cmaW8Rciy5vgEQMM++AFRqeoM4fmu7qY2vYVEdywWXgbOKsXWbt6co4A7yyf
b3li8iBSfaI2JOMO5t/oQ3F6Eo91EYrRXouJhg612HqDV4hKB1s8T0cvzrTH
sxdBRLVl1fSX6gaxAxQda7JQCE2IUtd9Yn1Xk5jEPQBlCmy2j5r0OCg3YdaB
OjIs/c3KpRtLZlvbwdw0Rul2VFebbR/a61nBCSgTf7mvFhNaHuJUi1Fafl97
BykI4wD8un4YOQMxKm5DVN+bJhrXFMGXZ6TNdNIBeQBgulCIwfq21M11Fg0U
e/WHo/xFGpE44Nhs+8WkYi2meai/PwN9JiLyALAx6oH3pXwqyx0/xwMwO1nO
C54PwD/6L90XzxUz1QnlzC7p+MBJs2/u8RZYShFzuwSe/v9fEWj1E2lOblBw
CglV6w32kU05e/sHos9h92ZNvV4J26smGpX1vuPp5RSGMwheZx2gbYt6vKxE
72sFP97o34JbSNKrW5S9znWpyf511CpfWhq6Tw8CL7N3WlrfOQp0cUEO2bzn
JSYwvsD6gy0SeiaAxP482nYwsjD9ewHgijSsNhl92czjgm7IdOke+7Vr2JMu
DoEq6HlqHunQORKdKmSX0L3rdWIgPtt91jwQu30w1qe0eGFgBiDJjnCoRi4Y
hd0F7ssWb1RmAVIIzIqpgHkfHX8ExojFwqL8UVoZeqU8e2bMFGABQOa3oln4
d1CLYegFu5YVUgCEn6K+NeygeqIhuH8XtLMadiIHa57+HfgX9jQqTqiBWfzI
JmdU3AanOB7QK6bqlN1zQneuiSqyQN3ebLkh9VnefiiUtkVcmNiSEUbMMo1/
Pxi9hL3u4bTVK3eNWyrMSfSEYL14YqYrZJG3E6nNQ4DOrxFo9vWs9f69I+4X
fr4zIV6bBdDTT2u8Bo2R58U4TMqyvB7QFQaMHrmUCn0kD9bfILKrWlp5PV8p
tdbqANScxkouHiTVlz+pF0/lnUEKbKC+ISNlD9VbSCvB0XwCqq8Sb0OuVNnj
nETh1NEqTu5xTtIO9L+UaGuPYXvTTPDj/udjC7f3nzfcO+DS2hjK+MRFXVP9
OGj/sNv3CbcmFJZbc1+TkDQCeG8ZwWpKeNGKJ2ht9YCO9MXLJuHOoDP+H7yQ
aE7YqukfUnVWNy/zGdD1ttm40diivp1gEE1MkJvU6FbboYpXCPk2cCHSXkBO
U4eAhupYEJm4XS56nOhMHtAf3Czlch2EqzvQTsYdyIKmPmWUQX0TTxgIKAAk
PyCpDAJorsIgoTM6U0hAf6d07YCZ7l65dreJpUohNVfjmyNTi6m43hcyWzyO
qhrhrI7gvGZpU2ABcPIY7EoAEByFHa0pvIdYrVSulPVCGYxuxGg64hhsvEf6
gn+jnsK34xNlBWcb/wrQqf0xg9F29Qm3sPpFa6ISILmVMW0xRLiLvx/fzmSH
fmPoOJfpj05z9vbbZ5MuJlTCnF1gLFBEN0iCij2jx66QThA7+swsjq5f/WLY
4pO+OPICitdIWGxJEp9z8v0+XZr/jMvgJHAIMPWTvz77vH/wckrpKD8BXJay
SArrpfjThltI1yIf2eW9f4UhAcJNh61y9uiI6qqPmw4yDAYmrR7lNWf2ffGF
0OPtW0Gp0rPSvNhqy4EHsNoREJLP6VFzPaAHqDqzk5yuU5MNotP75oQfZHVm
BLL0fyvoQ4pyXqGYXFLJCwAbN/4ELgBZf1jVX8fScT2pATjE4+mZBTCXQF5V
KhTlIMVHZ7TlplCt/+vwbMXvE11lYkVli7iF3qDDodD2bg2kKJ9PxL9NWm7F
u59MKz7DtW8K5f/hTskzx/G7oDhq/cxHDF/zVl4EVoP7G/EIx9bfSUvNmEdW
SGA/im7T1WcTxP3Jf0rOQ9E0rYOM3p1ood1vfiYS8uv/+S0LhLR4GZScilc2
uRGB9JRQxv3vIg+GWAjgo3EPR/YkKK3HRJO+Dn4I1MFalOKEDi1onsudjfDz
uz6BsQeCAN7yrPMJfTa4bZhibvZbjbLrR7WOw4i6hKyyxdRIGPxTfPPhctt8
wHNC4ZR4fYJOyPz3F5bW4a/BSePkNilZ0FRHzpPsPnoxP+rS+ww6C0CfnNOs
q97WfuompkP1XtM7SiGmXupKk//vHOPFt6kS1skiihTCVqh47yB6KdtOQ+l5
a3fAnoQI06N0joOeX3osx5bzl1WfA6oC65ND1g5Zy2DeANPxlZHMCTtMm6oX
3S/AvP3UAHJcUtn91KfeXaMvLlsyPCTz/JbIWPy1WMz+TS6OBuRCtSmSq/VH
CS+AWE8gSNqGSjKrYcgIEmKDfg3pV/GsMfnP4Oi9XTt78sEbil+aQvPdddBv
POuyfkBsi9x2AWugCjmi5oVeTGW2JxEz65CPObUrN2Y+92tGznOF3s2g6JGa
YEAxW8qB7In5OkdI2FNa0QhF+mCTBE/FVTZmh97Qx1Ep/RjarGMAL3yQ2iLb
vRfX+0VTNrOz62vcMTmHYz/2I4A1adQsjZkmd7vwOAqtv/GO/6z/iMFwFOpT
Y3rOIxRjFRYiZpr5aXDA05dp1U4w9KZ0j2Gyypuu81sU6eoCzuBsUC6DYoZN
YV91wW7DFg7N6Folw5JjmgT5YX5SIk0Loi5SQVimHJM8FvUGwV2jPe5BTPOy
jkIV/CcAxfCDhtXQ1K7ws2jAeL3hxnbYWAUQfSuh7dM987yhAilN+x/hYaFb
uusCTtwtmDsenDtiscshZ6tYjJydHKkJWrRT6N059Hm6GnZC3miWEzq7z3ko
6kHzWrT/HJrvLBEjy2Y1bPXssw6uYNuj98uCrIFBwac87Zpq77GRrhoqURIQ
26kyeSZDZIG7R8TvV6JiJJpNhCfNIpaDnXliRqMwKduSxAxXs1nKsCgZ87es
E2lFkGwCFBosaX62Pqns+1V4NMA5FbXK8tgQkUfEQzW5sZYUANNxEC/FCNdR
Yi6O7rWQyjs+DhqdHCbbdJ5j/SdYeDYUeXp2XbkIoc7LQfiRLq6N+y4ZKgmc
UpyvbALUqLBtuM12ue3VASQ7tRxHDnqdBgDULpZ9gKl6UGSID8cRkzWnvOz6
AZBfwLtJPTPiQZrMFoqsEna1+DglVO/WIU87Oh6tI/7wuc2WFqDR8QAaJLTS
65aNsr3xWLGHHnMH6wuFG3I7V6dqPmoM2VF8QC2MUO6jKzhEdoD3UYuR22qV
i9U2yU15zNuutzEsmEXrxlf0sZpBDUwGoeYKwFIv1dJL9CUOugtdn7Vbmt7f
X0wu4FXLmnu3xLlAJsID7VByYT6BdXP4yCQTMEf08NWGiFmdA1e4i3Odj1fu
ZFg55s5fsT5Gk8emTlbOGIUQqdVT1txA1iT4qXC1GQDta9LRnJN6hHg/0Fj4
9Vy9WmnF1yTPxFRczg9D3PooMrVPRYL4rxTgvVt6wSwcpups1DBfqUlazxYK
sMl4CSFDK0LJue1c+uuctmb0OYIZoyK9/dHYtRAbiTi0zssiWLYpKv9VcqkK
LFn2JOJLFF6EkYKFx1ltHahSDVKC9PGiXa9orswREB/32crfWR+vqZjbDFtQ
8WZKwiG3B2UNMtxFJnfomsB6EfiIi71nBRNmI4fj282089cJmcPCzj/ARC/5
ipFk7NuS52XU6m4igWOs8XGKXQLnUbGKv1KZvIQZbnbugAbjO1hnLCFrMU78
mmbGziYpm4cITOadntXC+OGuWlLYAMoK9YxF63qhKTei7tLM847LDqV+T8FH
XqFcLoJaBhKh8IUQ4P+1jfezBISemhfWz6UD5dxbwmt5dzkr9BahCRAmN1F9
M6UvACA+vIXIk0SNABuvqrsPWOxC4DVauVSBaiZQd1Hau+JZRprX5CmSysmy
gAyhie5Xqm+qcPWMb6BWLZGs+14Luzxz0jRg8qUCIIziQWvNbjM48JHAaVMb
NTkt5bS4saSDL7xFJBnEwrjt06ALpRUG1xuiiNONFXS2o2vl8yC/dbPqGE7b
NZaqrvB4LqjDSLMQdnc17KFVnbiYjaV/W4fWicqjfPHUCizS8VBar9vnLVr3
dR6z0Uu4yYjYEydu3DtZBL40A4c54Myr3437vApzDdwos1EbAM94uZf9QNXV
lhJXr882R+M9cBDTqXmXuD1BL/EgVt5IuMKPNbFwj5jK72styduTgt08LiZs
Xw5tk7hIeeKtaaQNJFwInk1zZKnkmpEZl/n73j7EfnAkrkTYEHcPKC4emBWY
gd9zlMsnPqC0OBnYHJl5v09PrR3yeSx9lVECLfwCn008qdM4LXHupeFtoR7O
R99PvBw2obx7Pc1vSb29twwIMRdmPrtvzIBBsstVH5sP5wvKB2XAHNF8JX+E
okOR2jMGZobIirWllCIMWiI+ad+nuT80LFJXHC5d3XjiSrkoJuFS/nfw/yeM
bBoBYJWbRH0X+zveQ9OOMH7Sl6p36i4IWejilccTX7g3nmek1p7KPnuJQ2WD
INcxIEbkTKo/R/SxHfzjDlkNK8KJd+3fNT/lGmgec/88gAKC58fci7w8Hdsb
mGWu7nJ6hPsORR1KGkoilURu5a/iJFHT93vXi1sVONFo7VlWBtr0aOC2SsIl
04YLCAo1M4C2h7RFKXPVtUC3bR+g/oT6u476515wMRG93Oe8eKYDw6eGCNy/
o2T9DPBrEfOHgFIoWLZX6CnITcNXA8w60cWyaktZ5ZIEgwKMmSH3TSv7hl13
wg/v1CgsuRjANzAa37lNWUxmrEaAbXD6gNbbz9XdCMxs01xg8/QGaFMdeTNf
WlU6CPH7KSNhXl/Nj32JBA6bHNz+BA2luMTUwLgEoZtYl313lb/ldADjzsiU
MuhLdWPpY+p2g6FJR3jIEaBLZP355HB6H5IRKvQfgwVXdILMN4K67iu3CRNo
ndNmvR3ByHzuatv5y7Ec12cLUwAPm4BEtD6kw1xYhO15LOktXedDGNtsa6ec
JIK0Y0x/2P1gIBBcOahAhZAJGFfO+VMh4fY81DzLzLozfNj7ULcRo74m6Smv
Vlzxcqu5PX+ol0MWdNgOtoRWwCx3UUh/vwnAs4NnxPwZdgJSbT/9gHZ1LUfE
svXCVGzvuegmF30qZ8MeSRCodxI2StytitUHs3Oxt+U1dd9GY3spvheB2BpF
bNQmZaKxpzKFuBHU5qa/lQdtgJfUnYYmFYMHlvM/ECYSpF6EpAqh+1w1RCIV
UbvSSqcbu0WMBYk7Q5YtrSEHwRA/zeZRWJF0NiWo7iGlLe302nhFd63ya/L6
d5gcFeESZrDUIVM4O5SEZI6itjcIqzv/jnXt5nz+EY8+EHxmt8KuI0QNmC1r
CAZSZbsQZ2S67nl8/pKZeEI2TZVMr9qrwKaJh/F/lBXDblHQdGvyqVXGhnNl
/8SB/cF5c7BnPJ8R/sfeRTbryBqo7c8aYBNe5Eu2OWiFhML+E4+17oHGv56/
wWtCQMbpA8C6UO8XFFbvc312yiEWqk9p2EuoEhozrKSQOu0ybMJV1C5cU0bA
8qBZpSrJJ32PLHEwIsWTCtlW4AsHACShhbhq0XWldDk0QAyifsM0Z9QiUm0s
Z/AQwFkmqxLHTAwNZoJNIgnQp33Xz3OnFwDVpczOKx5TZ5cPjNJdpuzZDMOx
9UsUoVGLgaHGRlI2BbCRkC/EkfF0L+GFxPZhkifn5O1YAMExu/WtZ+qheLBE
TSWFbrZypXhTxIFnKRs0N4dtbDazcuOIlSBMR9zqBrGOt5qWXk2cwBLX+2yK
BtuXwaTI1xvFyZub26ZRRAygofLFll6oaosYQTF85C6XEtGkRqYcGktDFiOQ
OjyT4Dw0yrJsIKajH3n4OTAEe5dcRkPFJKcuay0WSu/nL1e9MZgp5MOpICKF
9vQJ6cJCFxwDdl7OkKNRSKXZbDtrF265z84lu31LCsjL6UJF/N3OX7FdnrLT
zUSZNdzpM8SdlaIQ0gEqGOAIudLyzi3JEbW66pep7tcJ9GFIpwJxciniJyJn
CKATqKRiL+ruGSgPjX6KLsuiw0PJxebxztF4T5lTtxqGzOjVfKZEnfjWawqS
0NXdOzaiZG0FHCI5iajYPQH2JraasUI2OxL8USzMB1xvAIQANB+92iZe9otv
/qRrPTdNv/+rJLy1/8yXy9sI8IBaqR59y2FhsIpS82ctTWT09UkfsvuBB3cv
WDRzypN3eCdCq2e/mfvWfh7R0i730SnnMmzNMMsNLbTLKiO4tOVUNnykERyL
HKmWtsk7OHLcwMnwsLiNH13ewyE0px27WGFJLDBndHPN96/Non2GaXrvjZFP
1Xd4hEYWKOw/gbyyqfhoIjHN6Bf+PKd6Sq40xqU8t1DokkUgordsTvq8KMPy
JSjzmraPwIfxfVY5p1A9DTWmiNE8Kq/39cQGLLFCVQDuVWxaBd0ncMbjzKxc
XoqOzsU1XdhUOJPLQ/qo3Ba+lWOb3j2J2kK5pMq5OGhl7gMczxp8XwRXrJ3J
1swlvv/drzWvvGIPw1HBmDdROZnUydK1yIq8LJdDKx8KniYF9QH8Cjcg2g+p
hzNRkM6KwA8N/GzqOhGFWNe/ivq7Poh2/mH0kkYW4MjSPhrH6uPkyNEWfNKG
y5CVWxOFaD6lLRWd9ddGvYlt6oVTi07ZHZBqxUY2nhNqcB7ybq1Ve90Qqoey
/0uJWgRUQeyR4nwYJR9WMzLW2qjXZjVaJduXjvAxXCGCfJbIbThVNmyxy5aa
hvUqEll006fcd53gMmFVaeL1XO5+zMCLR6aYHrS1SexZwKV73ySz5dZ4/PRq
BIAjbw5iP8ycG5z8JzLwNXwEV06Vg8IagBLnGS0Cmz8oePpXHaZ6ZcLhzGOj
YKZA5450adakuN5xcUCrZK7edtKEwMICyEfCCxxGETJzvnvdWvZkX1cOif+x
ExDvzWdXFSvz2hygJJxk4jmE6cLqzPcyuSZfChBB2jz+ZY2kaxjQbt1LG73u
ygLGdSuIwIcccCk4ysQMjBbn+OKtGawugcHS+2pDrzRSt6FVjST4H2CBhmZb
Cykynclv0IuoQgfsz3FuBNsasNvmL8uImKh7tRbOnru2EVUEzBqiKjeKMgVI
DSLu9vbzajW61GNt8soffYCL+n7Jy5yBThdDVW7lyDeQfzKdRcff7TSZyHX3
1dULRiYNEi8zpUDWTE76hzrZXlSvGVWPU4KFqH7ePGG6cb/6O8+erwnKxvOB
5d6Yt26FNyIpvbvgqtD7No6vu33PcWdrUwT/mzYBACHl3zPnU7ZZQHYZYQ0n
H8vjIaZO4gyfTRLccKxJHcDactGe4VNv8gT8TbJ2zDU+7OYuEhYgZT6S+qBn
Vw1NOrlcrOWHj27GoFJa5XAtM7HW68X3LLCnCO/jxgIuqgdjpQHFjmhF2vCc
Dlu5tpmYQFJ1dMxs29RasLEZABooEzl4r1wNybp6QeHZkg2HLe78ZTg6bBee
zwnjDeaZNX+1168OZsBnsjo4g2XuoV0dUDDceVOrQlDJvt4LoZQ71JnG7tar
6ywwwwI4jK6cYIFWNbhH4sMjztig3z/K1XvmiOsZ8m8NwtXn2EQgH4seXqoX
nG0z2Bvd+KGDjLUraJrWtS3ssaUCoYnOdfha6rI9o1kgEuLmlNX1ms10/AWm
kv4T3Zl0D3C4olUJb6y4ozOBfdD7l/KTAsZD6OLIunGt/Hk8mNC9umso6L38
Zd/S/XDl1wtr2paqRIN9DHMbUEAdYUWGq3+pcPnm25VMlhFomQhrgOX5oEAp
WtUXs8s1MBc6ElEGWWMyvvCY9MJ8fcF2hf4PC85WBDZ6DSdp4cBVMFFVCq7H
pCiUSslHgT4bt2apRPgL2358rGugQD2oF/dKOtKpqduqagJrInKxXb5M//Mg
pXKopDQ4MIL0vdJmH1sTVU9xwfvg3JL3OuSOLImP5KrMzEHYiuS0vRbl08xy
Sm/TdtYDRoRWR8gTEv37wIPUZLOnOlGn4HckhqCHv7lP19zOp3ZiPASWxygN
WOta1tGojEbvOXyUfFoQeIKn6y5P/BrBXansLIDkXkB6SYR7j+SlVQsZpOuC
FS1LjPG647djt127u7lFNegXPdGmrBW4mxDHjXL01/JRsUT58yF2onUrWJQl
wcTzQPeHA4E6Ue50arGsy/YadWmwzQTt6SjM7L452E4+3vNKPqeH3Ce29f38
SX3noxX+WSkm3ykELp+oMbRqcUIYHQQZpdS9UJTcJYuk1YFqdD0DtZM241Qw
CrASTaJc9ZJKfDm+ZHDdEAdKDE/Zl/AsY968Ckem+5Fm5ZMC/z0g7sKdTEyv
8+wQ+xUoh5tKz7g1Qr3yPwjjdK6bu6GJh3ySiut7SQR+J52rE4yUIXp5Sb43
agbx+a2KSwvNmSisoq6gcoGL1kA8vYfRtcU1cwvVFRy+NfYr/95D5oktLc4p
pQpSjEaUrEwdge5JhJOZ9TI5pfVLxKbs2L9Gjfx/i/TSfRIz4SD9vPX/GGfT
AmMEGMTamTi4gJBPe5TXLn8HgC/zNFaa4SuPHTDU3KUpR+oqDEgWsU6yv5a5
q7d5l8/g4oSx6RRsT1t4P/mbPwZls/EgOkLGjBjtE3KFN92AzNLr4oZUB3l5
IkGr1N/RM2ZuQ04od6/Xy118C9hlH6knU6VXRnUn3omjGs4/vVZi/nzm7N5f
4sUGMvxvGrzKHv0n2g0vIVC8B351OpibX5sOG3KIYM81Z4K+q7TXHC48kteF
oj8RrK9Es44cLWYbUxx3mj9fvLchR7ujMFRvuLKo/BivTffy0i7nuL8fikDQ
xaXMeKzoag1zLvt8QccC7+a7vo99wxv/hfSMsdpvJjnHz+fasG7yDSgAq9S3
5TlTTWf1jeAPb4enN2Q4w6tcmra+SEMzGf5xK/FcF0P6/3Vd6rafd4bLvbjD
jdQBDPlTLzlYQfzbmP278/XL0qSNaxRN8PJhNpyrA71TXYjO7GYL5wH1ID7k
SoMUiDnYgYadQgPmXH2mRvBDdeOP6T17RJZ+NO5VxkcmzzrTZlmcwzbndYr7
2Hkqh4tq90k2rnUu85DHigAhdmODLqQsPiRSpaaPJjOb8+NoS6AS+Z8uyshK
UBkHmCi8mPuURYXdX90zCfCOZe8OqZX2PlU9vhPmaqYFD7WeLFVbtj7YW8+r
YSP32iWmTS76H25hQHKyEmsq4cVGJdhM8hYSxfazwJ0jyeI2CfV1ueuKrJiF
7y39bM0idpIk0fcrJcvKAwJxKTak4LarmgihotRe3epNJH6z3ZE7rHGwagyC
4Sl09/NrjylUFdPt53Jw32Ki7b1jS9tGAYvAnXg5PtHbsUtX7CJmdUajHWEE
m2O296NM5t1OXycxh0lr91Rtk4JXHpz0JLVpB1MsMILL1dCGwpQyCHEQSqTu
oGOYOCXT+98z8gQPDO/x1qNATqX4KjsTRZ5ybf5XzsHiRKCQnciBjNzvK1Wp
82O8eijmHhKP07NscKmcbEKceyKSCxaoh4sUDijl99L7ws3pkE45TYHK9Grp
eKiAJZ9VpO4muRBqYdHNUnwg5AZn6vjwEVIfevGjubQWNwBbagFAAAqr/c1m
JWmzsCQJUKXzEw8qeJv23W0ahN8mAUgNiX6IEjQboVJXLUS9FxB3KIK9apgt
9HLKpDDqRIQpOtJZtVsdFjOFaI8DPQKH4Vn1FGpjOPJMCR35NYXVI+165i6L
hSueOtOUfrRbimnwIOWYRPeFpqagG1so1pDzEuaufNjFuyVDBVE57dJMB9Vz
yGeoaN3MkU1NoiCmYZoOubCg8Vkukx3BhxKK/Bv+hDukkvZrEwIIEoKBUxXD
R5XtNPwtDLRSYkEwui56xffdDa0n38ftCEEGJG1aHxB2S9qN0uYpcWP9E5iJ
4rjSAPrpP7zapPpHvtR1Kkl7Y2+i2oVZ22l1d+r4GPmiHdDCxVDVutHTjJjv
/Rp3mSNyBmDGa8ji3rwInOIm+Y7XbCwsoeyW98nGvZpfWSWCPBITd5Je9xdO
BhWAnK1QE0Inoiyip5i77z3xauo/nuO+ssfiSqsYt0tNzwRoEHtu+jdbfiwE
Y03RiiRe4xjgo9uqzrZBJ8rRQL6sQVzbIli276Ae/5WzxuXCga0jEZP4xtCW
4TVk22B4bDcXEYwR+5EHtC1bpvCf4lIEZoa4j6anS/3Ca/On/qEN2M0bV7q4
b6Tol5ANf+7qaw/5Xryp12+uWnPuU6L0KNJeucEQKBLCjmY6MHlvG3EUwgrr
YqtzaCMzaZoNQdKgq96xwFzzq0pQPthvwO5Hw68La2OUVyrQ5pH25P2zmdkM
gaHsQrmp8IzjUOkFyWCdiCuJpyvL4Df0sjungNLJiomxAA/CRFy7KuNngSx1
VfWguf04QY0Z/cMCmf5Dc37mSoUZ1NMwoimIctGWAZaWYOhx90AxVJsjRiWu
fWRVK9aGtSXGE3AOOiosuc82lu0lCcRfSLD1utkAnvBQZCVxiBwXqOulBSFH
V2mlcjDE1V7XLf5id8yNaHyxe+RBSqVSVtHb/C/eDxppANiz3mWsuRToh3UN
eDWSWlt41VXg/kbaHa0uAQ4ea/1RnGb0eZjVZjF2ZyNYp3yvHx7nQFja0cp+
bhoC+adIrpJvUIgz78S6PggdMQxqs15pDQeKx3HuxcPk4jUGp+MLQyQmqclU
KVTxRX+dDeoVB4x5wmgF9+kGsq05JNZzgk8xrofDxv299ogIuuJGOkTarHnC
k0cz97knkIpPDuI/rWgebtsU6b8fMnHKSK+EEkvcHDARHMWuA2V5Khe0ASFP
2/8zqNRUTexvTonoeU7Y1ncdNEkryPHUrd60VGaZRON0t26IRxrlixTBcrVj
ScFLAzKh2f0UmDNhkzrOr7qGWuERD6l3UNQgoFg+ZSzg6ErqEA+JDbjESODP
p/nVJfeQ41vHxPaRwLP+appshT70SfwJF7naBjjkLNnvMFGbVd5Dc3Vk2F0p
aJlPFV5RLv4YvTD/unA+AGpYzy0NdRQd4EHv8E9ExTNSTgr2++7qhNfgaVaX
1CY8csPnF7DPsZewn1H8GBvkxxaft2fEFxxaTlPfErMPF1XOPMq/bWatvcN6
cqQ+KX4D4fKweWfHQGxZwg3gaECDxkVM35ysRSuViBAx6taLyeZR9ZPG1+GL
4Dagx4i5oaFi9nbTyKPlEDVSNcw7B+levLebef9UcpGRKEVkSz5uHG0RXx3Z
3GdwB3Sdven0lNWn+7IUASzxL8A+WpmKpMWM8sbsh9bZOZQ3gE6+pV9DZGNY
KML5rTgaop1JLB5SA2XSW98ywhhIwIhMhcNsVhiBBIOV26g6G4ACarMSZLF9
tdKIPSlRepKZyBIv2GGfI7aIAIG/ZwjX+czrROfhk8nSQzjN0hctWQuqVDZP
71PvVPaGYGIi4G+4zJHnAfCXL7ZYgDzlmUES/JHMnQ+iVpqxrQsKb9yCJYpz
Jozaw6h5Vv8JBIThJtOPVtNaJT0XSe3M/Btsu8vI4oLTaMJVDwalKau5KBMB
ZU1kiIC/ln2V/abwbLJjydq0OqklfXBg2PLYqlG+DyqBS3PW1Y8iDhfJYtzb
jz0nmd+e2Yq7Sq0CtWeQolzeq6CqQrVN6VSUsYbwsyBc2t0JNBWFIEUrk2/2
uj4pP4z33HbNwGC3QReDIQ72UjOaA5jy55XPi38sX8dP4U3b3GmSEFRBu08G
7/wStBk3QFSx1sMaMrhCpuhP+jtQCJtGTYHrWbrgSrkREInAkdTsk2uL8IzY
KAyDk2dgVkm8L3JM7EI/WsCu7L0C9zCR3OCWs0Awmi1y+grzKerjdEDZwU4k
sKzV8YKhZQ8YZNfK5ttadYIXTQsh1ixpTuTTHXBBdHjyylZ+ujCRUNiy7ISc
GQmGcX7mqZt19DOYhiQncQ/drxWwHJekubDOVxw7Q3Q1jM5HI2mso9uXXPY6
LD5Z4DTPp1P57U6rwuwwATS5V9eWCPKE/nYi/tggSbpzPb5kn6dWv4Ylhk5j
4vt7hOyJLjfNY6VDgfB1rQ8ONAsEb5nXAGCW882o5enz9LxGi6h3sCtDtTvP
z3YK8K34WQH4bkako1ggkNDFyE6vQJfh1ysI3FJZ0h64nIcUO8aZ39gTXfI7
3HjtAZLsp7Lbkm2bJ6SLjVkGNqEV7EuljeNDJ1u6+d9h5tL9PRrVKTeWlGYT
iDCywPlEx35OhC+QxduhAycV1/NFdeq+Dp8BsmZJKqeaxCkZjMp84g6VcYDd
Nn0SRehZ3XEeIxz8oLwvhq/sSxVoJtefhrjTHn1LtHK2BdBaCyUtuuQhX4i1
eHAsmYxsfu+BDuBRzu0ASYHeoyC2Y2X9GAP0IdGiSZyc+SFy3o8Q5cRXH1WX
B4d9W39NvkqBYE+hh3vSNWOAHcludHhYsS0MZoa1saqxP0ZOBY2zpN632+0C
O5Vzgd8/7dI+RYukfNvmkLMpPBbSduqdGYEScki/JS/k+4Qepd+xq0+Ik/a6
PZZ7hDPAp7dWWF0GA6op17XwtNPUaxM1/8qzU6eZWh3kRN0RO2rvgtWEssXp
USN69FzxEmVOeWuFyHKQ2lIy+aqYnafdH5vLGuGx5vw/8m5rfBgw/pBl1auI
1dtt3ti8/cdqZrc+M5OKeqVTXKYxcbF3foxoMFMILsUMDchikU/1GuGn47W+
pSF8qPSW7X4WT9oHWQ2zZHP6OCPOvUPX9G8xrlklKLt/UsKaKbkMWrU6FTtI
htR0BbYsuqOH72uC1f93zRPJAO0J8Hecqvo7G3BbNtJGLpCRgG6q33x37fqg
t8G0KOdr/jJoMSTOzMuNoMis2CBuGy6YZMFjhHp97slK0aNcJiGv0K0CL09x
o+XZEcsWP0Sjd804R0Ahz1gARqfsH/VOmfuGrIMp7E3oOJkRWziOpbW/HKC3
DXLnOAFdOm7PEH37HOjeLGwvaK3Wp1W6yVGaks+hjuYR5lkPakR3c1GO5c/G
hXtb3eqaZup6nqCFRR8kQBAzq1wvcKFrxa9QXu3AkSrbscKgv7iCUrGeYyFU
2BrfOGKK8X46np2h72psxuKosBQ9i8FT2e08Zwe5MiHB2qiw6O+YRIbO5LBP
anai4zdnjwI49zqHgH8H0g8J5iaAgUjWf+ZA518WOaF7ii567Vzfma3Zo5QD
pNyML4IJOXMlmUq8+e6TFDZqBTRrNWt+ACbVbaV8umyJZzNECGi/gItJC1Ol
MymNJVqN5H8VmPWmOh9+7jpyxMtOjqD3gDXuLlEj0IEfCaIJm1nunUwnjpJF
CuOlGNoCnzUF7TZExhljxki6CHcTrb87UhN37rhyTYdNhowenX1OdAnaf28x
wO4QbfjjqqJLYd53OWlRavCxL63R2mt+aXhOeS7ReSGfQeQKzPCnG8mW6v5N
NIvittkpjKNndjX7pkqLCIKovIrFNBCR5FJM/H1qKkNuIzsNdYdXDgH1fjSA
v2dcXHWclKtwAA+3L3pTuqRhKdZy24C5IUCdOVKp5b06sncTs+idMeojsRA5
M2cSrb07W+GxPWvtFsiPF9RtMEFNMJ5DDf4ZbK0QQhtAoTFjYSoLbQBDdnfx
QWwDZfKytWwIYzIEWqe0dTebZVEvDPll92ykSipOUrvVBv6c6NYA4DoxYtAf
Nd1YiW7oUzBTwb5WbEXsZltvYohxRS/+kFXDoEHqK3EiOi+4oujbo0SNcLU1
L+HHmfreEnBvIrv+/5Tg9e1pl0Atx3UPL0Y5hi2dtY02ReuFvsvfzgA+F1v4
FUDRDL52L024ORxFcU6FpfiD7imFQuMEYNtqnzV0BLJEwJwK3iqaRsu32yf2
E57FOzSZqVYy8OvpdjX6HmmDeREQGiDPb1Sgw/VAYEe5ucew0i9XrsOpOesg
abC7vL470DDab9yEB8RgyabdxWqmZttwTUMhivhszqjFUh90dxsCh7RqHzpj
KOgNAiPjPmGWmkjX7bhdd0F5zVcbhojzEO/5xXpT3FlY687sKnh7LtgqCBZb
V0yhEiGTJAbv07EA3Tb+PQF4+bSwmCrqCE4zQj4f0LxfJQ5Vda4QMuQZUwJA
W3ye3KgipVmzqXpeSA9jB9ILpzpMvoAMe1phSvsw8ZMWjhNjFp/vGtV+jwAH
Ns08aH0Jq0AfCZKZqxnRF/D8aOxCvHpxIpPd00ut577mJlVc/zbIINdCF3+T
6zN9tYzyzokShJ5ekDXO3ndSayd6oYHf61oqEH1r1BGJGtuRzfP9t6nooAlS
C88G2HlMoP68istd9zbKy6mTXCVz/r73+FL9DtB2VCf8eGCBAwazWbHNenMx
04tQBHn3w7RTshmB4RJHTOC44+p6uk9/r5AUccU3aq1rYKB8l14iKL+fygOY
D5vu7dtO+7qcPRP+HenhSiRNdc1i7n+fiXihKBw7nYuftHA8aD05dG+Xef0o
X+9wg/xdJg7Tj6VxLfWswKC3sSte8jbELuQsPJ0cg2XQlCoHPtszliHWtL/7
2ZRjVeZZO42tc53Lqv2Rten/+7RdTxiXUrilcD00LS8//Ja23WVWVEQzdXs0
TAsBQi7jia24Z3SfazY2fM/vAezETtj8jfQynBTFa3lvJZpeMU7U5hFtRhUR
f06tJst+u5D+wisH8kDCnfy+k07rheTbSQOzHCBalpBc8RCz67k65LNXDDhD
cioGS+6qFXKnuQBnTaXDZWJdniyu3Udcg4uc1zgHVrSlhrDa1FT1OHlbzztP
YYmL8s2DrFzde6l9w0gL2D9rL4hvgKfReNKym/6C4b5eyVtMHfM+S4j6LTl5
Hiy4pGQVX57xppL0SRaiT8eFIUwoFCGlE0pq2jznrhgTm8nf8Sfu4YioMygJ
2ZQZUuIkVeRjn0bngoydGHWechVJpx4wjiXclGNHzxZMm1dLxIdLm6CepvBO
hgts/P/cXkQ7SuU4TmGJRq6Erdb50ystmPw0jgfVx2acbc0e7ZsiF8BYbl5c
TdnFuYDQ5g3aaTlPy4sdFJUnYJp+KgHbnbtInV8PNDBPXKyGKWb3SPl2/jye
FWc7pauDzKCj4Tc8HGY3P3H/z8iCADPNfmEzRq7gRqHciZSNxEQXAvjMM8GB
EAE4C3riYKySWvBM0rkL99ROaWufcYs7slrPErGDjKEhrrjFR9vlXzTI5Dw3
67T5WWZ9VSuC3DqZzVHI5FA68BjfiCf672J07aa9Moju/pwDMbudxD6hqM9w
+OOn5+Zhgsqhm6bEasLcoNoPIYqsW+yTi6PqQP6w/tWo3SAm0pFGvjIqehr2
uKOri/qWXpFVGW5S5bWQSqm6gGlEMJnfxjhWcBJYelhmQH0siBENkM24LDI/
fQEv5iS22GZ2IeoeqioP3IPDROxH1q/P7Hhkep32TtNJ3FPa7DbDFOuv5WIz
iKE0s4gN29at3/fwDsvayfZP4UIoxM8pDb/MaOQljMP77lfy6wNFQQFnBgAq
o5PHlY4ERrTsw3ZC5y8cEoYswVjh4Kfzy0AQ1dyWmcvZSyFBraU74QbRLwmb
um9/rZ4lfSkeudDnkMNNVjWDduslakMxt8U4TH99lKEFlvQFJZAt8HYDDR6S
q6HgtM3ow1X0Z/HSViu3yDUCrZNxFQIqXQIPJ8OYYyByYKHIZz2DKAY5So5a
55okKzIOc1EXGi1WzGXhvSR/ZS8tqz8/pclD1RT+F+msqZCi39u5xiyaZKE2
7Z/PnHmssYadJR2qnBwVebqCRgvPb2vh5cj20DjUokdpmcO5GFMh3TmYsx+t
a2SsPr9UkygdHqzr00J/ng5olWxVFxrUoR+0nlJhLQZ0HShWRDoYoBidOP4a
6nmV+gkVlRXv3bhNPhPIM8PqgtutpyZ7HoVkJiQje+6edY0I+Nk+dsvuF740
TvZrzI20juartKkOmYE6B3fqxAEXAf4T4CKoFyY5yCOKnnhp/HFPeDPe3RjL
BfroMcqF13T50ozIkMcox0IFsia+IbwDxbPWIH3Icc1sWy0FgZJDhNFmHmoH
WIp0992xekEvnSQy0nwSNuRAMwow4tpczHxb7gVc5yGHmIrJqsdN3g5Y3Fy0
SwAc6pjyFktL54WS4ugI3LKDuxRci0XQACwbRmxpYhbSL6jZt7nB8uI2FApW
E++/mTCklWt7/RjNP9U3+Tt+iz1aV7i4mZ3CmmdvrulfxVzhXRlbr8Q2YgCK
xYwE+l8iLzC947ym2RtPQJsYGKq2LiXQsllbFd5zpSm/FUhrm5hnO2llfxP0
K5rk3EZ1SVRa7bVdNTGfppR4gtX945C1S7NRtolWCuMT4fzCCpgEW2hVjqA0
SudCxFClUrZAN8sjJ0N2rekvyzDqU2y9YunUghe0lm6RcYPiEr/Mz/yMNCc5
hWdwBqvZdCQ9TzR7x4JByoijUBw3b+9CIHfmVLRWnuSdLXGkxhi9CbB4fHRw
TduNel1Pi73lLUhX/+yvDArSeK5LHmvXgmOp0dqI5z950rqyenLsnOXpT1RE
aTAXJqskJH2AGkv+G+gGcO5hZWv1hQ8pmoYaYXuQDQLTci3o78Cngq0E5WAG
iygBVxjG1FNK4mdD/nbSvoECR+XpF/Cp3KzqmXV+RfFZP2wZzruTH7o8edOl
jTbrag3iwHaiH8+K867Stcy0kwlkPjVCmaDp7MS/p5AskH2NXxCm5rzibp5S
GriYJKZmgkDxFxbsQngnhQCLUVqWtmSuK0/rtg5H3iLH61VEPXKlCezm+sFa
4pTEFbCZDKuSkrehGOURujnKXqWBzt+rEUjJOr8jWEVt0A2JdaufNyYNryDA
0F4w1TlyD7OHloSbiBH8BCJfQUHXQSFV5XkC+D/YwgZHNGPiXBx4CzIG39+Q
skG+3+qQVR0BQcH9/4KxhHgptRUgc22C7Qnoyltn+39mYvKfXBYR1Cr/X1sv
l9SHHMBL3Cp/VStXxbkbeI07t8tCa6v0JbJWV11K3v5U/EULSB1yeDEz/tuo
KFGcfknZjctY5N2No++5m8QyK1GigMnQG5d71REMPhn+Ici4nqkFlgCkHRXL
fhqA7FEWev6bM+PXdA17aLA3JBJw9fTotcp6DNJ5gI9c+2XwA3LhJpChExW8
2G+dC3XH2pJn+grjt2RKrzFUhquXFIxoY0sdjozp3+dbAfkBsK5II2xxbP5o
1cVNhohASVi3UmFSldfbq3vpgkkHDklOHJtveEJuEDC68PeApftj8FkqYiKd
YtoKyM0tvFrMYm0UhvzYtn9eeNUO2GwuuR9vpyPHn//g0fcEt3eOgZTIsFkE
ZwwYQWIi/IvfzHGhYmWraDwAAuwLh73HzNLpZVci03xTqOELcUjdIZX0sFOS
41M2rHwMgXomIHfx7R/oyWg7PU97pu33Zr/G1hw5hcKXrd1s7/Zvey5yzqaj
C3OghH3lKjMewm9VnF5xOuMp9Ao253g5OUyNJlT+2LhC9F6x6V7u9wTHUu59
U4EldR0Zu96Ri8LpikZkdDFj2BF7SUdIssIp3QbLKX6hrKWT3f67e+ZPtBCL
4nkh6FeOVmtMXq4J4mghg/etnlm6L+iH2r3vE/6OBW8dKIvcLRvjL8F0WS5B
DtLNYBCfcOC9wVTgU4oCOpesQ2znVp9BIVCRvO2fgYgNJ5M84NscNcoLQOuc
ah/lBN7IUgJsKa9i1XcfLfF9sknQIb5u5+QOXV6a5eck/3eDa4XdDeliABhi
EC4IDgfanRFveuoDOUiWg2QZLoSTh//JpOKOOAMzjv+iQiHYjx++i4tl3760
hEE0gGXJbeHZOWgVc0TQFBoaOyAe8kiVCMnSxxk4z977NH63jq8NXc7Qo86y
fwAj88jSUd51ZE5ExcdZXM9aguG6UK3jHw1XxXrRzmQ6dnAsf0zHm2S+Yjc1
wMUq6Jjq3/QXL4kGg6zF0LXDqxKbQDgxEzYxLSEIa+ByqTNP4HLnY/jkL3p5
0p3fkjIpltzLs3sGUfuo+V0sPNdeoiGcllxWcgEZrto5J8WNxZX4oZ6/WA+t
tTpJBNVdHHDeHZ2iO9c/1Z3+X0hAWjeifu2I2sr3VfP89IhFxJmRQ5Sjnhkw
sER2b213l4rPHcYYl4pHVPcD76ERM23y8IRBEODNy2dXhZAG8Czs5cv3Ozh7
qu/iIhMp7d9qYkayt8dE8l08DP4VeU1ylB/06DzUqmRHptP5Zw61aBHFpyII
LzLNU3enA9n4fHLBhY/rE+wWfou8oCuf0jVqwv+c2uhAdRHtN8SX/SQWhKzc
TUt639nRD7CaSCMYnN6X2qz0wHcpFWy9MGq27tf9NrN8U0l7++l2AaZsgovw
gJ6LV7Qa1qlNdax0oc/VgC0ZKXVpwySCKlqGPUtR3E9nRJC+MNIN48zznnX7
ZpVg5WNUXwZnRlQ/A8P9b8g9uD9wQXxjIY+rT7GzlMDTksa8dg2npXj7kBOZ
9RBCTAG+PTAOu3O5shazSQbthYc7Ev1TI7aQ+x6tALjKc3TkTrlbty0uX4IU
X4NRFfbS9q6aiX0hmfzqX7X/v/8b7E7RB9Wa+LwAy5N3AYaJ8CvTebrGhqVg
Gmbq51pJwIANg/ZuTWLNdF6k6YKWlnStcwB0knTZaCNxuyEnjSBKi5J1l35o
x//+w6fVh/oXFSOauLz8L9c5tWpg+h+3BQ4Th+zoNjDjY0ShbL1RGs0hStgO
el2SIPmAaIvEd4QJ5J+5IriqOFdcQKScz9l1ZotgyxPdFrzuJq9cQG0Jd289
xFH4trN3cRCX6I/GAtc9tqzSquQn1VxWutCsQhlR6McjvaQfpXEE2kLa24hI
ch9bLE5fbhHORYWVj4BSt0hwpocn0f1RkskAQ07ycHitxCLvTXR7oyln5e0V
1vfBE4mxdpz/S86mxjRC3+4t+bXEKpNeJtQKS7BsLrQXPBEgwIBfIJZb7Ytp
SNHrogArIRcPlpB+/d9dLvUayvwwJhg/hhsXYe3dHj+VsDzDM+bnWEVt/hZQ
IRLdTMlRjqWm6nIZS2uA8ZC5iTPsEAJsaE3EFT2QmrZHDP77RvCAr/dS4R6M
dfEaN/jWOgv3xC07GIEmnePMttgeKfR8BZYKOZ4ajfwIX8iXHkNy0OG4aLWa
Fx+5ksCQ5bq6xSkq3xrhIUqzKIZiJuz/igf8uB9WhOCb/oOk4tC5p9KZJ8JH
F21yTCceO5QNBdEC+pM9bat6AXLCJAtHR7G5SEk88a5mP9qsWYF+LqUoISAQ
e1PP9Do5RftouF0JIM6cVTU6Iiu9FdcNnLltNZgyuQkulXsNGU6+S+bGHKuu
qJUdpDCxDwUNwALB5HUjoly+3hVBkToPzhQZxoWXjoqeatH8+Evazjv+G/3d
dx0UGzzuSoVK3uCr/dy8oV53TzCtDk/8Y4se6aCdUMVVSZcU6fnML8X4KC2N
yKOTqctA1KhHum83tLN/Q9gTAvDQ+5bUOSNBzVgOYNoWzHgUTvkzBvS7AeH/
TPIa8KoUFoFJXca7VrqcU8XuJsJnXrTuF0nfAUpOYUrJvLp5TJr9i5P37H6W
v3r7HHMmqMDrZ1ocKjw5uafVdAz+gaEgi1UL51t8qJNnOsw5WP4wXtScAAw6
MZUg8xlqE9d9DgijFK2ZBmBUht46ibBO0s8Q2HGt7UF8XkTx7f992xMkEVJR
3JiEbjOgQKZ4zZhhPjjBqeRLla1gBy9avN9w3Yu8wgWvFqFfit31xIWawnGF
xYtGonSDBxSy2j6O4sdv5DZwvsXIjnEx8f+8XsVWaMJT+29UvDJRFaKRSQ08
4yPYBAGssAqvhcMuG3as5ERjsMMgqeKzykD6m+fHkp38fshralmlYrNnSj5P
ezBhYF32ePn78qKy9yNaVpaJukQD/dBPLo8oFfZLBgv5PU/hwcvVSVXvEG9s
27PEWM5NAufHFZsaft6w1vbLkuJLELWKKfrv+aIIqItx7llPOimPN5QPqBxk
MFKkXMaMwY09ExzI0KxDMOn77au1dBPFY4p+MfYYtC0O3R8lPyl5UVunOHel
pJmuWrEh2YpzHllXb9vGLoEmmYG5j/dEJyutdIyFbzmtktUmM5p3/vvZMNjY
ghmxIVcHi9N6NDKYX5X6+x+uuBtgnvnG+0Y75BUyXe0eY3ZZdhiaC6IoB4BV
YzG9j2+n3aU2OFSkj0qRKt1H/QVrIMoXl6bpBs6NpCgNexd8yB9RW4zo6Cfv
Ws7I1n+mAy+I+WyWYVT1d4mm/d8IlUBemfzR0c+8Li7Qmgd+gmbA/sFk8RWu
oZrBRFJnG4G/Dn/IphHR5YV7omLnDwehL6KFoiAwnCgUnB0gxGaj3wtXM6V6
LwSFv4Xs697SSrqv9x5mxNrQBYVCCYa9fTAi5+h4WFumrnnnBZ4IrBfitSVC
meQLlusBk8m51c3eMTuqmMlMLCUu3ow9WhDH0Fccy9I58GTVENjJxajb7ijH
Wtxkfid1FKIt8ejWVJrKC4E2RVMiQoWGXOjCcht1Vf2AMAQ57KLfNJbFA1aB
OABSzJsDsdJ2sfP0xjZeGSz1hEVa56Bqhk4XVsXrxPMaYngduVG0rhynIMxN
ARMFWO2T3+4BTQ0Y3kGOionJGzXV4PYzpM6KDHUX0vpAmqW9/2if4lnA7Xh5
pJhWaB9OP8phkWPVzuJzhMN3jfu3yewK9hBguajvorwGM2YQQQYzpZUKbUUx
7H1diLWEkVZv524g5I4Fiheqlw6ApOD2J2yiBHQOMbGokrgL+DRw/vBgc5bQ
4O+qtnFWkgTstPj9QjMb21E/7Se7pO3cgmnXbg9lXP/FwXNB4gcBf56R7HTd
6Z8nIR27SmK7A445gfAlIRZ49mC6WrMITN8zhy1qqlwfjT2f6Z9ZbRMVpZAU
lRzS6VWp0Ovl3hyaoVTfMGotXj9HemoFFyW5ciTKHHwr+dHgeUAQ9+AyXLZJ
6KUq0RQLK7otVWBsRlq+CQdyFEPgSpLsZa/U7jRLtruBuJDhRzLtXxE5ydMG
xM72m1IRjUbNPiRiFUTWStndRLES7AWd9AQJac9QsQVNlkRH8ESQqce8P229
bYx7RfLWiAPseiB8fMVmnSl53/PqhFl7Tz7t91LUvr4z0aF/Bbqikj9R2NMx
3SHv+G3F+ZzRZCHq8VnKpEOYb5Jhx30Cn6h48zrmLjvmxcaWU4n1XgDU/JhR
oSK+kd+ec1WzFgLwA/RlZcpMSmDL3RjndBsVsIZT4ehnGIklItcEd+FurV73
F+xLP1PlZ73vWcFgVllDsB3Q3meA1TYgyxZqZOsburhCbfdGoRosJDIHfgv4
nlEqsDatI5PhMTEuofyeZ4US+5tNRJkaFHfP4NwwhS148duexVrIyfenFXl+
JD5AyjaL0YS8yyEFdWxFQFRpgpKUAPDTimndX6ipT/gGJh4Gl0OyIQV1Z9qz
n8whAkfyA1ZS4eHUxOc3pTtqg8eFg35UYSajFuMJDTFoMjp5KPr6OKFUuJix
cqePZ248aemVEuBpqeZ49cXHt3sqcXKmzUJeNcWOJ5altamjk6mEgBZAltZG
IEWcffY5jrwTym1nDX7P06C2YHKOXkRn/IHHnQ49Xs9ACXCwck8KgNd0ozkX
E+G5LE7TpHmhB9sfJ62cGFYXPNWkTQ4myHu4B9fQlleSJRn8J2iJlHNbOn2w
msmyypeVIpSSL8u/ltvLUfCHaFFJlkx1qXq8q2aotsw418knfl/fYE3Im7mR
qfPs5ewv42crwLsq/9T3PSvLoI9RnNjzqVsauIIACoDlG98KrdZcCtKbwl9W
LGyJX6U6w3wQGgHdWA4/wCFVSWztKTz1BXYsdDp2Ffe1vskh6UgD7FdbeQh4
Tudjdca6hPNtWeW3mi3FKOqiu4+PYWMGusoguvocQ50lndB/4Tx+0+MUCTJf
bzDkoQZpMyP1l+89KbJrDhahkcBomQqaLJTAqq6Y9Qx3pEJtMiQ5EwAGxWkd
LvGHWipLoowaOPc2O6pKO4odVBiE4Ct+KxluPMFA/GvdnesFh1cTXZFMz8iA
O8+eB2g3Ane08mySVNLRvd7U3T2TgzAjJ6T4d7dfvm7y4iQQN6GtnqRQm7Pm
Clpmty+iLzsZUi88yz0ao3eXeKtdCCthpNzUhPz1fFnz2gerVfKPGlAV9q36
+EdDdO+3RDuMayo8VTpBQHSeZ9y0QF7m8yhcdl+TAka9qnL22BcZuTzyVofd
nYtqfUfCRhLQBZTzdQkMjN4N0f1KYOsUiE+79OdqmUihZDkoi4duDSeXfDOh
zyUfDmJME7dMaS8cXViPfUJWP+rjgo8sJ8c1DRxMPY6VRx0cxwOZcPmYllPa
r/hl04cdoDR2wjqEQB7Q1gSQxPjMDYB6sGvBShfirNK6wZb3gyRL54778v/j
5x9T8PB4EJVcarYZXQNJxLk5xxy2RwU1y9o033hBPwFxQ1GHTmwM+jX9FdPT
9g0j4bui73fjNBi1RBevsAaUejE3aO/tsEgMQGvXiTI6M3ZVnUgPfy7nigDm
6uBMWigVLeCFU5U8hVhAmLW+hXn16ytQQwZRtBdx+GaJL91b3xvjpk7Y13pg
AyJR9n6yt4kyj6OqPfI8v3/qHgiqv4ixvr8PygeDDpkTHlanwl/Tgsn3NKoM
zTc9ueCeH/GvHdYA/cJB8LRcedYWBk6ZnZ/JkoyJT/bQjPWkDiRMIuqga8Yr
YvHhC7jZr90VsgB9lIHoayxirs6eH2FLbHbneDCLRMcIGK4hS0e21jbHVcj6
JA9jyMdaq7RZyyQPr1OIoOee4p+svY/s60HRaXi3/lWYQr8SBfugUnmG4Oba
1+wkOh+fOt8ZHEu7aKtmQSKTNRxLqo8Jq/yaqAYZJ0RMZtpoHUr1KwvyFKxF
yAk+zmcM8Xa9DtPG05wklXkffFwO1XbEQtykSFMXBSGulwK9a3AvbPjwmmpA
oVPw2xiCXFGAuN21g7HrNUnUTAMmwee9OuJy+qVCdLKHZZSNpbBJP1pSui4o
LKENL7iAyem6tu59l0xXtC5gXtVN8t2+ZAlZI/B424kiUMWuODXVLXUpn2y2
SJ0VMtHQJg13wvbbsKQMwfDvzJEpIeFtY2NLIPIjuzYB1YZuXx77CxJAmDnp
v+m+IkwircJOcowGm0iXmBX78YqqLmFi2oSJjFXOfY4Bb14CaaKy7smITP6X
fYP7q4LX3ZZbYWMO08oHaE6GCsz/iO9+w5b0zrg5VXr0dDCp2idiP9yBkTBO
UGk6lU3cc6/l6ygvAGvWqgZ06O7tNnDSnJ8elLffV1GAtZu82NNiVLuzOh5g
KdM7YWWernBM1K22uxTLoZ3cJjUcLQI+S+HW/7ilmYqlsV6sT7xRInTcoyj2
4/J49cWEaTcC1Xd0e0fwMaA2c+PDC5Ab+sxZB/kJwLFkroXa7S0iW9WAJi4G
+QIf3AZg0J9z8Ag7eyEq4Nwx6PUy7XAZxeReYgNTBWyyBWUj2wjF6M2smmlp
uPTWnAh4wQehS7U5rJGbzsm359RKwv2Tl9f1n9zdXq0uSa+aayU8o9KPvWwY
8W5Ul5HeonXkN3FRNAPUUTO03/mDrO9xvbZ4oMsmGs53s76MpUD6Qm18VhHv
wK7AKoHvHlCtw86BBYaeasrXrybCh8pvITcAhqFgYsF93iCQAiLs9ptbDjIN
d8jCuQyVeiHt8UzMyuRgb8XUOfAuY0fmfarPQAk9/zFij4CcySUpcIHUo+Uz
qjzjRsJiAVLsOhLQmbkPz6nNNBj/8LzlBgX7ApMi8b3RHW82v/XJi2ymxKCk
lUkBmghTzw+F3tHZ8GObGSy/UmpdOvKvIDy2TiB6aWhh7cTXqNBDhz+Nv60u
emhebI8cnkjmCqoTzNwkaE/+ScbEtg30781ZI0JsA+/owcjR/nXuBj46yoID
WOtaUSz/WP9k94Kqfh222DbgKZzHLeMBfPewvhDp51kzqJ9V2DdDxBXMxJpu
3dxWjpr6ZVLksnfSsca9eRNxjr0C4drTkZ+7YtIzGcEOsPDanONcGco+kiXO
H+UX5LZusOLb5f+xZ8BWZm4RKhPQJgYNml8nVG8yh4deW1IelfhohH5qYI/L
WCfBqax4M4jmPwaOw/+a7Ct7JNQZ74oXm2PB5H+fcC4RFL/9K1Q5P4/u++mo
fMtx+BQ2mk/G1ZVE9LbwkvpKhCPzGH+A2Mi3AKW8yRKoFd9CUizhK1+sNXDQ
LnK5o2GeWVxIxp4ZQIlV1L99bFFtdwXclOi795CXDMntwwZBpA8Def/EDvDL
h9GJ270Z/+xc4CPh7exfM4u1xMMG89Wfnv+P1MaRHv2waynmi8bN/Ow/olB5
qgQmN51pv88Uwn1F0q9KlfdgajH2bJ7oAvdWl9MPUrIR9+mu5ua/R6HEHsT0
8dk0b6AuJ7mcjkMNKOQByVxxJbqEBzM0B+AoUGQbaHQeAuq98yTMSmg/JNJ8
+xNK2UF91DnQySeZS4L4xXItYZSELC2QscVu94YLBYZsSg36q+bKh+UAFcjS
AGEm+vuQD5SHBqPRPAPGZJx3zIQAkKLp1K3O4XIxF6eMxuhJyiDRF3Hm0bXz
5qjyFCpt+xh/dFKG91Dim1HTF8Z2i8hlNilL3oHYYIY0RN7/U57zRRJNX9+t
kt1nNmPjtpL//e5afEwG3bNpilpdhw0CDPHGR30zd1njWUh/NH8PMoGpWASI
xsR+JhLm8jxjz7tVEpuLOCjn3Sm2Ps5B67ikwqQ0w0O7IZ6Mi9jChbi2BRlb
NJTXCheibRyxlErgERHyetkT1H1DJv3lc1PxMDQiEHSE1N57r2x/Vuug7ra0
wTM/pDgq+VzpjOwfBLc0PsHvWPFm+OP+7kXShC6Hdrt0i3EXp3GA7AnZqIta
yX58Hz4sfvjQy49Vy52t/FtQNVJx69p8REUR4aBorC4OO4VMHBn2m8MM24mp
pmZWu/8sUxnd9qnxXu3nngd4nexES+bAytkvviiRzOP/kKNmJvUefoRkgvRL
kEEHWNdD62turyw84AaGDmWBJP4VOf9+BZ65S7/SGuenLkWYr5u7L6GPvslX
ghoyYvxaqomAo5iKXOMUnJDytjWINnmQ58WEpRmx6PAp5Gz6t3Ndy+uCelu/
dusJouIFD58o9c/9CWwJ3oDoSTbIwJoLEAQ6N1DTH3DufDpgVPMVz8qz9oOS
gH3iawCP1682LZKn60XH9TE8W5ZgxFsRe4f45W5sOhcuYfKgSCEAxIb161D9
Qa+3gw7K+5vQsIue5gvAcf09J1CQDEhrcujHjemUYkEblLtJv4NVRIUXZl8C
Ku9ElltWNwjhFV4XBs2ef1tMk3ZpyOfurlV+iEmJ8QzrCMo+6K28VR4ty/I9
NeLZtRbz+HjAsnWLYbw2ydswmEWji0M29Bk3q6GoGFqYVGJtkrZ0eFKgeGDQ
gDAk+cEPm08OnoUbZv+3ho1vxFQn1c5lJFiFprdPcGCN3Y2/7fmhrz18ZRh7
cybhhx0O+4iStuG+uc9+YpnkvysX2csMhe74t9zBsciNL0woRrQ2HoZIIjeD
jMSPmkPFbbAEZVSxhIRjmP7k0t9mUh5S7+od2BQnOtyluNZdZPKHGS0W+jsj
680z97BwZg6f0Loo+slo88q2wSRd1779qjHGDfM7zNOZYVYzfeAioqvmDPBR
KvzzDc4AB6fptwjbPiA/EE+Fq9zgpQt5nfaIFTu6lR6/tCpaC+8yaj7ltt6n
U/MLigm8jzgctrjEZNP2zRqjSEh0CD+tfDEjthnGkSGFojCXcRACKMhqOrDZ
94dUVb/MPzMjx2Bu1sosKfj1LUcejXLmu5L6wuMEHY/iDLvbSq+5eYsNeMn8
I9ttNtdX/utHwf1p30XzPVpWntPcy0m54xPE+evAeGQwck0EaQCiiFmobXeM
A9YsduJ8VtchmnnY6Mi6871+oEj6s6jyE3jA1+GkT7Hv/rjJTUTp0Qx73Qzd
EKGteQZsXbLgIaWzartxgbsnTdGUuhlRnJFFZLZAFz/ajPCUKCMvGpDnxmH9
Qs2/i+HcgLw1vOVpzWlY8d0jYwkB+xaWORKcj5a/2J6KT/xTaklDqW046kCU
LmcVDQUadHcr/Bj246dUik2mbVQfHVDY76ok37KxunpUrGHKcm+DE/Dkd4vd
3bPMC0rgmKsG953mWIMe6j4uLqS7tpRq2LCE1znD/0rBLG2E57w4C1xFKAN4
turDLj6QKvjYCk5tjm6R1NK6TNsQygK61NcgXmNAqRIuZYvZKFwP5gL1YgU+
0KVsLKoWFgQJXr/9rBFr7Wxdhb+bJR91rn/IOmBAo8HWrbsNd80Gvsxdrep1
PpE+bdWqExF7w6XrtNcpWXq9u3+JKyFC9pna30W7kufvJ+PUGAtM63wzEjLr
1edJDbTScM2zzblNRawIU6PzrLQwE83AtKDIgxux2YJzu9YQx/j4PV7Y0Mwd
Yu+770taf+Ek1/c7EL9To56sDVnUN+eh0DeAJsO4q55SSJJl4zO+lr2+lZQl
nPnsqoN04511h9Lg/tLVIdKWYt4qgF/7+jutdZo7W5PkJ3S7NanKDXbOtExd
rpUxAtOk3Ez8AqyMAtJ/X5vUAlsy4HOslc7aDP3U2N1KKD1N+RGaHVHYFenl
XQr1D2dd/0qUM/wk3x8ZbyW6Yw5v5PTOeHEYhHKqptEbBA6X5xrZAbiBPdfe
UxDKXprmfrONVdiq5/obk+6gLmrlxqcFl41o+2TfqPKCJ5O1r4NKygL+xibf
lKhtbkmjtM3xcp0GziNzvhjtocP1hhk4TxR0DJjzUf+rwr2X2YCcp6CMacF2
HIcMPlg7lXuTSrWSpYRV4/vnLOet+0OYqqB+ok/y3+PaG55EQLVrquGP4Sti
ZDulesRfPx8Enyf9TIacqsmNWhp+zQ+d7llx48Eqa4WckJQQOvfOKkpyrKiY
avQXbqXHkWuqaaL7Ra2rpROJN8dLD1if2QWQWCAtSxHmI8aBy2BpucYnNYhB
m8fx67JuwzyjKf7F7MRxORtwbv3JvwbK9ca1prGBGBUZ/e/4iJdxjo02KHEd
6LF11zyrJ7MZXIGA9NzJpX38fylC5KE0frItSwHgppqB1UQYWnRtUHA2DCSP
aZTuLtnm2SsELcwSlIgyO5svQwk7fkeg+ClVXOZA6Q09tuE/TXji+JuEiZE4
NT9ecqYqX+zY82e8IjKdDX36M6j/kjrAtyVNL3MGR0lTdm/URsV+BWslwyOm
+EKpLN+P6C7+t07bl6cRQWpoAHa+bnlOtEabh/eOJMeh+uPprPRM11kzS1rR
0oPan/bbyTL9gkE5osf1VnEgBZuqIvRjQFv9oAg/jT36F4TVmuhcZNEKJaRA
vFohwGv0vqKq9VXuBQZ7MXcrxya4uyrrkRu0Qg/InEa+Zowj3MUPBEhdhRdU
EsQ43UP7N0ORyLgTHvthSwPWEOjme11DWXmcySSMvbymLgMYkzsrqzG36I/I
RSLAo4FIe0Gc0DOAbIMp8UOO4E5fbr2m4OvJM1aZoz1xXQ88GinQ1eI60b+2
5r3lS4rAxvn9GML0qVtt7w9Pp2cESTEBWY+ABgYKJtlydEZkYlrXOXIKDuss
9BnYVFR6+GPIPKJO59o1FKfVnOdfONXSvSHHNYaiJxPCFzLZwwKrnOvhjZx7
Tnpd+t4QpUVo63Ly7/Eddpv1PxZrdYclX7bKQvoCdbuNt3MI4RkDqqvBELHo
aZtAAI8nZWJ4gc21TuqFn7JXW0YUc8tPXekdF9xQjZLfSDK2ajCjq/OlvnJP
N506Gzxfd535GU05b7NZ6x3BHw7N+K2mGQqY2IqCLDEOl+wXAjE36wfMrsrt
0cTNJLVghD4T9/kqvfc6M3B790labVH573zC8ip69x6RR+znQCX9d5lkpmDQ
b4cwzp+jm+P4hqwTAlnxO8roRJpB0+/7PAM3bftI181NyQ2xum3kRqY/JU4K
Ij892IAcbtbDriO2rUjy7n01cwbMSV7zanVTQvNfFr4dNVSLsFDFPfQhM94W
/1Xqe30Jwd0hL7sYhE3FfN0CB4+QVG3YMLC/kZqCDg+99Q3Jrdi4qtno2/cF
56qSj971ZtdvhUV09fHH9lITRBNnoVg33gt8leR9UB3EFy7q3XlJ9R0B1PQm
XFXeFHh9IdByaIoZPUBzKJ1lBIDziM81urT4eSuuUcF9Q4iJFjK9mX3Ab1qZ
gF00ujAtnQIeF95cxOZClZ6o7QzL2/Q5TEE1gt+8+ligbl6DPTh4G3oZCVqR
N/Cfmavn1pq++dfWccQFDq7gCb2rD2Ni9qevlJpym7nGszWS2y6lemPuKTyr
ta7Yaf0UPEd5KtidFpt7qia4himOcShJXGa0NXBeFeIXg59HM6DwDG7bvds6
VDZubRK7hjbpE2BZlUfs7kKf9R1f97xdZNaRrxJ2NAuZWLcbAf7MH7NjdKL3
vO70DT16kjSU1uMAX8J+PhDzN1yHW0G6Q3ZjGA+pr9xZcS4dVzJExCkyQctT
+b3vre2j3xMDkUORNeupgH/XyKnDYV+A6lpT+h3FYB5B2vwhMZd1gYkD0V9U
4lFH4YF/ImNE5H+DDGJY+fur8dLT/n3jNUlGP+umxEzIWijecU2JD0J1k4uM
MhxycNHpl/VhjJxDQUUpCbHgIIAM9KjcqoXFnUZKr4FqhQwj+pBphcRqtTV6
OhIjcL0rdsko8bT+VbXCNnSW7o5n4nMExq+61kchlzgkqNKYp8N6e7wjBowz
jzqhvIdKfaPJRgCxizE2R2IvggH1q8G4qO7ynvOQk+oOmEAE0ETAZ9Tf0vgb
f1glk1v9gg0y3pL7gWsQgb/vUg/+9+z208tUjSawle3+8XiLVYj7BnNNSDxU
hU0u4gMe98rBeTRUS7/zHDuEOwIW2FTTPCM0QCSGa04cxeY1lTeKgDIRu2mQ
kqZTRN2UQTZvCHI71UMfQu17L/e/W4R2VsHH9WDdVyWZGkkZrJFHG3C0m6pg
T7jogUDzDi7yWOMROylXkAUF6VtxSYNFA+mFzX2f77lRHlKeROj6A1O9CUJV
FHu9lgGOxXtQEAho2IMfj31oqwpxCv5r6iDcINsjsSJL0dTWqW50p/fuGegU
E3OP+I8K/IsvTU/VF+cwe74MGN1msh7yICXvvlXi96x4VkyFjS07R/T1C7Ix
ptpUHq0VffSwr0VYKhOR0Dk2JRUGpT9SZIqwjnXUVAKKXjY180I+4BOZ/r6u
zpG0tUcqEL9gn+CQn0flc4eQgZ3xj1LIAJWLVXqgkStAEhxG1KzyXxLM/AEj
kLY+y06Zh9hRjMzedC/As3k050ZOTAmrUHKDeAi2DWw2hP5Ibt3XgH+dCJxO
KAbcIU8/i9lLVJtEMuGIj2D+hOPIJSq5OpG3PxnUbiv56pMKJIHE4QIAfrT4
4SbgJrG8Evkn8RaVmpbPah27wI0Yxb95JsS8uMusvk50PN8RC0xTs4EGZi7y
R9LhtPndu/+RzcpFZ4z4cO5uEP/zY63XDembF97YQTq265FEgvq+lgYGo53P
xR4Sg15KjrTemSJ++I9ZmCLLXRH+WWKJaAq69e3yAXQeu1o/iHBJFcCHQzsA
wmsoLLrau/3URBfYfXYPUQs5i9GpPodoWrG6vYEYogc7fF+lnmDJetVFJKIf
DCuR19QYRmTbnAlp5HFNC7SuvNSZclEcmRJd/vLaDw8qQU+c1rfaJ9IiLqG3
0MB4rvHfSlgTASU4gsZI1N33q/8jXvQ8tumVfvygHv9qdF3jJEP030MRKrpn
Zn1rGcPih9r0TbwUSHio+VW47VZlJUWVDdvVIXPybLWOHsLgWFck3ZBniIa9
xmJ7dDCWkth6BxQDjUv3LfixRlxyVwsrVV1pDl5ZgV9WI5vIbyLEsUaYJZKj
LvRoXHoURMRihOjlis5TxEkUMJnzKoSjxRDQS7rYOLiyHgJ7kaVThhZZFovS
KQHUixbjmStEo7fXKBMR1fBvPV+XsZcxrIGP4x7lmKHOfGmSGFcGugkYw+7P
WQ2slIsDcrmKVrrK9ppWxkW+WARrg9YKNI5HUmwpJKtPHBVhPyZQjLSV6iv6
HB0dsxPC517cpdKshrbCgX01C7QE3H3CN1NElkT3Z7cuUHHWa/nSJFDUMxk8
jNKQdtAeoWp0WA9LIeJmMRhcBdj+7DMuZuvKnEs0bGAZ1d2WOTky0rVtl/OZ
0VO0fkXv5i+0G8KPRORJDmX/Eiz73NRUGvhAUgHrN8tFKVodoLg153ehVRz3
K4Mt0xbKOOTzULmJLBRanTF7jRNV08b3+O3bfOues4UiZvwGEDj9Kc6DilbU
JZuS7JqM/7qFZFORhrbYh5+dVcZGLJC82A90dAnSnW293KtZf5ubMy4anNqt
eqrJyFT3NKPiBvUKT6OmUfeNc/FeAORV6lyJWu8+rQ/gaCsDMGJAjXwEAP7t
VTTQyFAFnObRGKhFUnC+ymML3i/mqXCQc5hXDxkgBjIYD+7rWjYVAHTT8f42
AXyyW45qpaHeTz/+eNj0TQwjUOMzvvelwX74C2DoEFsAzMcR7Hz6kkQImzgq
/PwQrC521Zk52Gzt2B3pRiTdRTJLQPJTKONiLbEnrchUZ8kXjZRv0IkrUXMY
Ag3fQYHBLeCOlljHJYeKr9SmQDEjSFNfz3Fo7jvu5WBxWJ2+pZl0EiqK0DKs
wDcmMbBY5HJYYERGuxf93M4jUdAX/cyLzgogaae8iegsJI3oc5s4Yxd/qE9g
YXzF5HNJUXB7tDSFNhtP+i8BXDRy+rwtl3WNs1+D3k+mHJHnnmcRXUhC81z/
P3QAof6ObmnVeSmi3NGYSdDeqLUKIKsbtqhqgkgBUQPe4LBW+CtK+cuUwKU4
FaepKaY/lP8Quz/ws3+tEJstohTST6mT9wKrFHFI6Kb1v6PENmh/k9F1EDPe
jNDlM5Yzoc/sOOCpSK86RV1vtadKYVpgggTuSh/V9hmMCBZy+0rE9ripP26c
1GlNoBQq3MXFcDYu1Wy3M//IOwpLoZzkohfQ6bnvR2OG2gTIjpDLVOpp34o0
olH9+2oOWnA4SsrPTKX1JDKyHF3C9FaMlEy2+/anMvbR8SGbXXTanMfkvc6N
5fVDTt5RalnBDXrso3X06cJdNNgf9zOCs1YUE9Gz098YsN6Epmts3eodGPD3
gcN1L2VRzxWVIM+yjwe/aPdPJMhGtbBGCs7f5XQJ+zvVCJJPLIR+Rt3/BA6V
MtbkcrM97FGZWqFERldV0E5DTZi/bfNhWpnAeT6G08YEqK7I8zDIYJYkpJx/
eUIJULY7R+w6Mlf1/i9TvMZvyxZunV1eFslT4trKtLmbEkSYSgs5mLM1zefv
VwBlehV7UCGoH0/qNMpUpCe0H6RTFjtmGs0NR2nn/X7rL65TkYr2zSCv3U7L
Ui54Rp59mWEHn6jSAIvjebJ2oCG+Dj8pPBE31C4sBYdFIPeckWku4bRBbFjZ
Ak2RcGJr6WDOYbTqheA+F4+W8GirKG55J8AckDWnrmIcbCY78yPQqrXDOFIy
RflUlh+LB9o1/8cnpDfkuVtMeuJLK0W8NEAa7MoDswwVi3hVwORiCyhunZso
Y0lHOwkckw51K+TmQSnOV02t0sHHNF8qYXceyGZpBo1mrujR2ODH1mAsJkpH
oj1bg0NnlE4gWVCgS25VN5V/MNQ8rQgn14nYPGQpMWHfDnbqzBMr5V8skN8J
dDR1JUepqPLHdTp15WtX9vrBjv8MYSnX3QwLm8ttaZ+FGPowu+Eusn+qW972
Ni7N/didPrETIcYJgYImd6Gpgj8RQ43GC2HNV3+ogFA8zfOsVkukJtlqPfrB
GYvOnYU2lDA+sXUxu8oyhItBfgzUnzceuSrW2iDpCWb/HFxCV3JQflh82/h5
kAy9wpo8gt9r1cOLsvqv5E/Bb/Oqb9ubhGLoz7/bUIdNriuw4xd20c4RhVQ2
cyH1mw4XPrbAN9L8itqbH9e4yg31Frq4xJHujQKDgDvG73ARP0NgWaF+CJZj
N7Dq9HZ33ZDWSU9MXSncDWQ4BtkYa9YYIVs7iWpYhGCA+M3CHJV91Ot4J+Dd
3tyD3DraLVTUt4tvcqa5pqpB4qxbALIRcoX82/CkOAM/LDuTHpbw38q1UUs1
+4E0ktFBekmROLOl3uG3fYmsie/0NmTaW2SYPzJAE9Raub7vEuMqdrZTkye7
1C9q3UgUa/ij//idPopKV81vVjV+Rye5EezO4cwiaAvXNyzDwGuEXQICfTX3
iYAAxUDshHThAB1+FFk/+hgroNahj35UB9b0YZo01mkWhC/5O1ml1dMFPUQa
8oJP3oFdg2GHHTn9rERnkk0DEaoK2gaivY9+P2w56MNkThfOaix0DQ0doGWc
6kmdY9DDyikO91zfbg9cK9s1DPi8IxrJHtESTVVKIYYLTmtqJZhSqffYq6+7
wSZciBIEayWVGQIaDS4AlyJ/cGkWnt5dbaLAwqciC/+fZCHUDXstFFIz97YP
9DDhwnGQcywvkWbEYx8n6ocIk2/9cowLHq0IT8Q/IwHjOwP4wvrlwWjjwAyc
CkDAhT7nE39GJegScigovGo+dRo4WJrXnOk+msjWp+J6sY18vlchiYmO4TdR
QsCYUnmzALjEf/Cc4uu1XOIwtbuy0GmWFTZ9Rh2HGfJeu0ubst5t6WnmKctA
3CFymqvjaNhq6Ie8bmxA+uBkvY+DggXYSazoMNVCeKf+xTlICU4D+Ct3jmTO
echSPx3v1waNHIbO3/i3RuM9d1lwXxieJNUoT6m72kEJXxZRQEQRGH6sR490
qay1eOLrpRs40KH6tH6QA6pVdLJlAtB42UBvEipPgJgVI3C4pAUu8dQiJtbs
cGd3a7LXFORr8+HBrtATch1AYgMkEKvTqClbbGoVoz/nZCHAl3WJyNf/j9zH
gBHbg0QHvqq+5cyLrAvGBq0BmMLGZl9S6G5jurSLA8fImo9/+t5yksLKQbgO
8NUq8YC+hGNiGGU2lxV5CBQVO0x4sVmTi+JnMGr612FmWSRUuqg/vlaU61v5
sfAkfoC48HA1W/ySIYENlQObs1tyYFRfM9yzNy7iJuyni0LJxDLkpui/Akvk
sA3lPWqFi/w0VCmWVFdWNF0kgVQSYOOjkPB0G7/e+LrwqAmDywZlfoGk0Ndm
T++/UjETQnXysdM6SRcZdRShmoI9l0/W+C4+6zUXr8FjTW/qw1b8EyLv7Gg4
xvyqXie6yKoIkufcmG+5mtYpciHLZs5FtpQnF7tAAAXAPHJhTt3+fHbDRx+T
edyHfXKE5biZfj0TtE0tJjZi+3N5dcrd+pFjNbAwT/hkBh9ogE+ktzhbzgWa
sXsOgBOx3AqpAM9g9oa3N75b4n8iDRw5PMHVEL2Q4fXwg40vsbH1WzDvWdwE
8DU4Ednhds9MN6lxpj+TNjPh8fSmSuCPinyONYr0IATodt1mHLE4/X5Gv9xh
f6UvI8bPlG2UU1MfGYncw7hCDW2IxDvUpOeY6h/zJMv3RwA4XlvRRx7jGCWC
BTe2fGb+jnVbxDcLQoZUaR6zF0iCMzlVGcQ+krDl7q57Y0ldxyNEoRLi+3DP
ozXmwYdGD4XB2vFHF3UO4j6T3/mbTHxoEQuG3WpHCPm4Y/fLTaaHlEhRFQPl
XhdpOZmGbVBGVK5pOVZ+ZAXP67YDWb9wD65C/W1M3DFncV29L8yvSDW+LOkz
3NT/EBZO1Oo0deI+mwQ48SDCB4s3UR/wvuls/hbZ5Yfh0yvRD9uouRbspQup
Bl1vOiHesWK/ySzQRzo+McF7vD0jHydj4pjZ9SgNQJAd/ITDuuhlAtrX7ujY
umWSCxjMo+rXuCDoxTdewGd6IAE3mICnkXxZTYuP3X2JnXCJd1koWhyKaJsE
2KqGJfPooFNPPVqL6wcF7NDDnNSBDxWOYm4vklNTJoTdNVw9hukuGv5Jyxyh
Z5whHgd5NUFAFBTEUKntQMBrZuTmQXiG6y/by1ayEKcItwd8W+AYUb7ApzGC
OaUd6VefoLuUkNwMb12UkNBx9HK2QasWiVQORQyS8pcKNJxWUHx7kxgid1OK
WEZ1QZB+1bd9ZlzuSlS8RTRp4sFhSDDXsEDiCRZ6diIzXbeZmYedgtVc/NUo
pvc+lx51eOiO59xr0ZWVyyxqmSSJFWQdxQjJDIsuXilhHZ079WjuhrTl/aXn
JpeZOMejfceL+TE5eynI7LEb38/gDQqZq4BJ+d8BW78uTqr1MnDcMDf+sUkb
Sv6+77z2P7UlY/b62NoMDrJSt7huTu8jVeM5m4OB1ZxbMvZZScflaiOtfGyW
VTnwqp5f4J9J303DaZJ0LAnuGq08FXIOYHWwbZblRlGASg8xLenZzrVj12cC
Q0imt7qOL9jUqIAaUFgCIpvmEIwY9bF17dt5jqDaKzDawjd4FjuOSlWsSyIT
jpRUuOgjZFJbIwDOup7021MkRiRVSxi63efc7f4VjmB9HSr6kj0KRo56eJCW
9U9AKpOGs4XyHzosyiWe07sbcjOhKwDUjEvT4jQLWDYl/PFt1lQ8qPdUEH10
3rPWfdyRZdLt5Qgd4IR4tcL+mZeuUGxOckO8mRSiw2ofk9QwzJKcPxVIqn4o
zOuhFBo955WaW2s3kF4Q9dD2QOyLZTMSZmSjKZiXyDDsqZYLKr3TQ5e4FDcu
SYlavKOCVLPQUQWYDqXGuIp7ZcSXm8Oy8X/6x3/Og4pteyq5sLl4e48IpS69
QxcMSeJyX7iAbX8mjNblVVApfHQ3afOAgS0VoxiFb76UdUryYuqeh2Z+Ukoa
C0MuF6tcbrITexBTUS55bcoS9s3nkVYWd5fzsatszqWuPHxniwvri5L+R7gS
1uTbVPNtIPv02WQbSPXGpxEhZ4JSxOR5xSZRaOwElT+8dMvZeZEn6+NrPUPr
2krhR5ogIpPZvF5cJyARsHIdIHdbaCCp4VuHJc5CqdaGEF+k5sTShacwIYJf
7dqPtJsAOkyA6CiTmUDSneMcWsQXJtha4Ldl1xSy7UUXJSQwAfjhblOswyOF
GVeUIkPv7o9Glo56+3Mt5WAsXsRt+HPkCUv/1CMaU03cZzMrlCi+8MYz1BhW
PUFJrGQfMKcaR19KVSR5ZxQ/6cXfx4rwOeRLDt0abmCRhyDZHcPhpyNeOmkD
0H7NHQyXW5X9WBLoEecFX/dW8vRIVyZmUHjRc7HtRoBiDl/cgd9xNZKQYyJx
uuoZW5L4j3Uv/kOmzAfaGwRjYoJVt/TGpGmaFD147rW+k5cBx6++S+9w24qR
OiSfwaKBu5WB9uML1xb7fQZsQbX9ReZwmS1XS+K9ETHqt3wuSIQEff97IY3D
T4KWpHTFnkwc4M1w70/qo4OFXU50AfxwE1EYtFml5XrnDQafRgqBPmdycZve
XAOuCbVpQnN03SE/cZWcDLqKLPO1DhtVsy4aSvkM6/k0yVvabo4+OF0ONo7Q
4fjqDQe/ZVvWc8kdBJAX8uMFLPMJIn8Q4uEjaLjc46UXb1vPgTsrLrwtCLIl
h69df8P85zad1jrV9L21dxPM8FAqwetIqZuJkKW5bcnjj6fs4LcnllRN94aq
V5GID5lDMGZZC9eJxSTxm9OaatQ4DHCaVnfVN0uSYKjrUMq8jHKqDb/34+1L
/jILUHqkSJCYYjXGpXzvHpvKExaKbBUZ5sLsZT7NzHDdJGYVkz2DwnNvOby+
kIr8o4d035P56qr8JFDLvEW2UowGc97/p7IFNFptPvd6MVSo53DzYrF2/JlH
GNNGJXryEUeZJoq7cCHJWXg3y+oVgXlxqUHaaQRG08+sp1nAHlLC1Ig/DX+G
irdrVRFCX72fdSEtvBXKNaPAokjxqvOGnHHxertCgyBiPtdfiMUQelFDLMUB
EtOZSHgKCXRiQARKVM+5C/knoo/yAWMD3feWPYy3h9FhVBtLzp4UadQYzo9V
ZSi1gzqv3x98Ht6rYAtdN7ysxJKYSMOExSh7XZ+hQ+T7iILK93T2wi9BaRl+
bhagUbV0IrJGUg16R3biuju0/Hha/Tx7Q8nIHd07QiuoQjDcmdDEJ2D+UCnE
Mw736EVHiJTuZsOkmF/5eZOPwQkP0GzXd5j8CSOE5fD3IKIjBkivUCrzPg+S
JnTJrSMdOY0n7+fk32z7y6Ef0+NxTD2J4Y1EsXIO3ZREmRdkja72AwItMoDI
gHKuTc6MrJ6hjt8VUE0uTPH2x1z/+E2aGWvT3mZ0bF5X2JfHw38COdgXeDVo
ySbJmcKUhVL+eU/+uXaOTg+fGAHjXGpljcuZKy99VFsMEbTVJOMETXvqPHcn
ZRSIh1d9sx8W9cjoEkDygVbiUBR/gD4KwBF4BxjYB9IB/gEz5vr1yaJ3Btzh
VGsEuFvyFbjO6uGaH+ixcTR3QZKz8zS5G2gGxd27m25uERAwbsU8fdDmEcya
pfex6HOwHaAeOl1oKpwnTakehxCuLl8jufxL7CyCtsiYUhkRcUo7lzIby8fe
xXu9OA7akiWPc52rnnU7Dj5Re1NgZMkeAi/2uQz5BLxLX+pr+6ay7UboSjLd
CCm/C03Mkx5vu07Q3OXZv7Y+XtqH3Q4ob/LZKsVlJLXh12KUVFV1qBCwGl/g
rXiI0xI8axLJrpXWz39k2Vz0pRrXzNIUIAkWs8PnQp2pdpgfOWNgxpL1G/7k
ycb3vhgRIypvIlfHE/njFcgelb0gnKf3oK66fNtOjcCboPc+9nBCskbWjgqE
+Usfk1mcA6zxLl6EaSVwexZqQ9MOEzn5QCS8vuR0zkWRsgLSk8HNmqs8yZzL
Diw7PuIIymPXSuG0kPSVIyU+TIHxJNpiy0HgEO2dg7AbDtGw6O1KymWheUXX
FwmYDxdND0gFyPH5hG0DZQamOMHP9J5GFvaQoZyQVknbLjyuBi6g92ENTzqY
SBuvuvjSFs4J6A+WasuJKMuwTmoOs3oJjJi6bmlw9sRUU0QnKlQvW5NCgR9a
op+SgW7P0nsv8S9wdSP37wusi7W1IeQOPQASvblpmxqhe9EWrb+VLwyGH+f4
oUTPPYjdlhCkaTNIsqR6UOfGdQJef3TivqQI3OSnL/8DheZpIh+5m6B275pU
Y2bXYEqws8IVjdhy1LAqQePLSm0iaQdLCEnoWt2PjtY65xo+IgNi/HueeHn7
dTXV4FDCo7as+V7NRDbNmvX6E1rYUlRNyN5vtolulJNk0SbibdtmniDmm1pr
Nqq6fglx5VgGwdNpHlSQKiElAnhlbXgPyqUVPLdiW/bED7ejTK9kZZKbhcLi
Eh2lD0pgmUIiahcUicmI81vQKhekokfUZtMZGQOzKhwi41+at09SL2ZD0RiF
6fg53XD5U3OVqisaXgEDXvchwemhui3HGALQ+xAeqKECXu7kSTjqGIhh9WXI
3LoTvCtge3acLtMUP2BFq0rWvlQ/m+rPrMx/cfL9xDYeYGccZqX3sCcvbRqi
8xLPVFSEfgQCogwvzoK54mPo7Lb2Km0kV8gBOBtqCeyyOKKqmKLfb49eRsYi
kPHnxwVIzfrFiqkpXioz4JEjaMnbVwMDwpo5H75vVtyh79vLDpBAENRcLsSv
SuMcvTeGGJWNXeGSKC9iWH467ON7bfmsMl0W1oJgjsUeAc2m5RxZGRbfoKUW
dB3bBvIybS1OF9jUsQL8tiK8uk2KRQGDENZlEIaMRl4Vv99lRuuCmfHMw23g
l0S76byFZ5s6rKSU2kos6dy5Vacqn1ZnIQo+B0XnF5DXpoSE4WR1/XCOV6E0
qcBwUnsvl2mdPLyynKHZIcVV+mLc88qfQcAHGVr1YgZUpqKmUXPzTlDuc4Ah
Qq3SMRh6hQE2ezwlLPSrdUWl+4K/agCMpW6tRNFSvb7Hv7JtKwb+IupqMHEo
Zc9TCbIhPtMHXBeuVfEFKXLjGh6UciC3iVw1Ox+sQAhkCPO9crkeaRmq4hk9
HZMkNocTZPKU8n+eNfe+A45dD7yNB6AnxS78Hohe9BEkEPUJIhH9m5TqT7Ns
jOBpHnxcMjvRmhqjnauvIMeT4VnLNex65S8r2bkBZPK6MiaaIlJN2Xd1YobE
m/NZqmq8FbEfTNAGzmiOpmyd+WLaK0FrFnPhYkSnPtSFkJDHvv6wcE1VH0Cf
YfCPlu0SjW0OOVlPf0wAkE/KZFFyQfFGcVoT5ocI6Be84ykOC1YJd9gbMwp1
k0hd+hLFgigZ87hQWq55Y+1I2Di/hliRnQzqRRjIWB+WRlHEYym2CRN+D1Pz
WLeI1vELXcqMTwIDifAECzV6e3piO9f+OBpWyGZC9XoBwpiPlDU2loRj8yTI
3+oE9qf2BR8MmPRJTZ7Y59CiiYr1aI7LjzCZid+yOK45APlbj3rI6P/qnZGf
tmyr0tOH8o8k5YRmoT4oudr7F1JHs5oWvPTTzCuyA7ulShldCKiMehvJd/TU
FZcaq0wMreiYgvP4LE8WHsJWCqtXMTVuaTAxKWUwq0xul3iz4UKKIL/8EoTo
aBHa86DIKFGwHyvGoSI/oMtqvFiXNUm3uvId01zgdtvbpoTykuQbOoUff7Zr
V6ssBZySrqR9bvLfJ0k2fOHsAow5/FRLHirOUOWPK292fB9kXDw0nhkHiLiq
SDeoEAu+PjYy8YjEoXu5v5D+tbRBbSck5KIad6jERbJj4WG3ptZo85daLsua
u8xMrxASYKNK4L0nApoUMqjmOxexJ+oPaHB0MVI2rrFQpPLgxFxGk9QtivdX
C+RhEqAy+2F10JhOBkNNtjhoxOz8DHf3baF8ofLvN2KEcIBMArCr1esAz50A
tMC+Mqt9Ba86T0qITQ2McKP92riDlyWvXhtBsWlyvDSa8/Us62a0TpVTCtj+
msIMgWCXwQ2mp+GNMn28vUP0loQVf7QlB+UVpix2pKniqXhgfpdanWkZ3YOe
dfmq/r1zOJX3uYH3yJylx5HA8YegFesPR59HCULpLYEwXfeWfHucM+1pK8at
lfl6hmowNK8jrNvdCBB1dNo0d75/MKn+7iAxmDEi490i9c1XDVHrnMyVq39M
/1Ed/aCh1+icSiLCMLD76QRG1WcOxMZ66AVPRQc7rRSbRl81ivVJusVfnzAi
TluXGRfzLpj1OMXXnaVXlyedJZolisiHnQqj89+Woo+V/tPwOyXNfeCgeIKW
mvb+qQj77JthMzez8M6RS8H2tTNE/TfYWF8tdnGkR4BOFYZ2nAjINEJCETPe
gbxm5cyENCv/TcBkNZMwk/3QG/yMdLLXPDZI+0hxrUv7n+kX8rBNSdV/UtDi
sOfYds8onLaxjAP2qNk770HrYJBtIhHJpjQTmXns+pPR9CtgPvbE6axXFMjT
G0W+SQ4Q1fBZTtPuMU4z5+UCE6Rfqgs5W+3a695cTv63qT5wBuD4gbMJfSaR
qrZdX+/cKzBT/n1AqzLAMGM1/y7FsB5DDzZhdBwtSH/76aheWdSrRiGJnWvS
t0nsjRuJYms2iqzx0VWFjziof0sq+ntVMhd/9alNxLJg1gElvNGeG5IeMG1w
3EptvXtTtFko2YoAF/gV55C8Yq2iErUp3tU/SFoEaNPLYde9j2566xbKoSa3
VZCw/Ib/sVUTMsL/ZPIiPS2UKjia9GUedRUyGTS9N0tKqS5wv/tUMyua4f1l
yQP0KOot41S57AvvBXuskGOcZVe5ifCk19fIwWzEDUU3CwXH2jHMqzzRkw/F
Sgv2FNuM2x/TunY/zOdv4e15d7JTDZjWhbe49jXoxdJCpmBV6SDiUJCQ/+OL
xAn3bvm89kohTvIgJV2um9afJbQCEbxN5yKeDXqzI6hXQUsArzCdRESIhh7+
SpgexKCTt7vzPcUQJgh/UfIxNMmkab7IqQbLcA8AhCQi0wcXAIr96obpKiGz
0wU8AJN2tsYKNPp95UCo+xL94BuyjHbXCDRCk1dB5oyNpIIu6cgZOxF+6cEW
W1HsuQX29xqyIop+h7AeYQ9M3lQhZbY8FS6syLNb75JGD+4vkLWRdwnqK5lk
zoOFyvky4PE4DWqyIpUBOu3CRNBFURv4S/ZeJTKePnF+Uw1LL7m7XCfFNv8E
24lP6Is1m9SZzVuN+9Bv3Aqb0y5Kb//jbIgyOhJY9jeEFOWrHgfy4yKdfb1D
JGktmekhVP9mWPUyXCzRgRavP2RFT9KdwgyjhLEWG/YHkmA18QUjnKOU1t8s
hgT5xEcr7fNCXrhIRyio5a1SAGpTE022h94ITQ15ybhRAbi/uqMGqge3Ywhm
5llIkSKrmOzutiJ9oAGYcc65LCxPizte7d0VDX3fKkCUaI0+VCnGywKtNnI5
0OjAkxwgGJLLk1SS29/VLY+4eKGOPX2C8QgLaUOFUrkte4GqmJSVLEo7dFg/
Aw112+2Iqkokica7NmoBUIrnkRZTDyHR3QfTcRGm60KSRD/IwJMazLuun8xy
ip1XzrPhzw1+hUWCuy1PZDyApfHLalw3YwLY+WpTfYZoEyu3+jhrqXvxMdme
0sLpMlH5F8TRGmQX4FUkEx3n708aVLqc/QZZL5BnhyHsaz5/TMx1x4igfhB+
MVpNl4HSwrbrW878gds6PL9m8iC+FgysvpQfft3bUheoJS4n1obNtpQ+xFSw
t/gNDF3AnNwFwy3EHsm6GHB0GeIKW1HgbVWYzXXdSzObw67CsUg87ZxfWXMS
v+oYDkuCtmhQC7iZGDoJMgh64xVZi75gqoNhZJGN7W5f4uypdfiQHcUGMuod
PQChy2jiQTk6czESRznYJ0IzA1IyevueVGSrq5tQEdfkLkx4ejypJCe/uKrc
ViWOuCO74yKyNmdUWmY+ZVXFfRv3ksVHSI36rEScIt3XfVY2DOZM5rhnCk7s
vBNDsh1ywSOSrXKTKb7KltzbPCADid8QfJvcaq70yTKZ1HwHUD5PdOoNscxf
HL0kCIMd/YUwJYmv/T2wr+Ooba+b1ZoPNV429Ro5zkSm9fzhOUm4fiorAw+9
0xXrfvb+MgItQZUhK19WneOUlTXb5ifDsKnkMnUV7Tbaqa9MDTfhpoppd4Fw
O3JaHtOj0eCzMC2SWWce+ayE3EUKN6RUpSn4W15lHK0F235ilErGjr6ax67C
5MY/FnZZIVEv5ijI1EZiZJuC3GQ0QlM/aMwmBMR+JQAsD/4Y0BrbYjSUEKNn
EGT9sa6/ZcY9obBG2GX2UakbqdufnL7JpGKaSP38moWYt2Avmy9HH5tRi9Zg
/XlCy8OM1ult/IMtMWG3QgZV6hgPBkru4kZBeWgBkki5zXit8sYvKdlSUnod
0fD9EIzgdPxsXY0hpcYPVfdfRuLdNSyqIsPV7tKhW+y+Qxy3Dqqxhg7cs7yw
WubjF2XK8aqwUKB93sXnexH90YuaWHuxNFyqWrfy4QB6B4s/oLcrWT/1dJcP
1/n/j1QFHdvK7JJv9Nx+onPGhub94HuZ+LTKFqWGJnCMM1gotPkiiOUXgBBE
kzfg2eLy2fnrcRgpIa6HyQftk09S/QvQNrjJalseoe+OLYy9FSenh7vqnwxh
6LKTKc0DkcXGxJogtz4uk1DY1MKzINlTqKlD42hFfh3bey3VfYWGByohc3Zk
VKV36Ou53sgB3THMqJ8hKMecfbBvdDuTcyVo2pScccXEsP64I6feoAGS0WFl
WfmMlChST9Tr1O0PJDfESYxOGnuyNAe4WK1f5MfxQky7rx+zak5k9ki56r64
On1ORifJvQQgB3Ujswv0on9ldXAYDvqs/jG/Q2333BVqCWnZINDo8LthoZnx
4xvmNrz5f+cBHdNY0GZXBLl8oD45YbdwBPl8IXpb7n/96fBwj5eruLX671jQ
/IqBZKvOCHZovoLbHzJ1FryC24AvbbaxI5vPpZMLmQFgaVHdEFzVR0SQGLvK
zvVmBSPN/P0pGfk0TWBBMXFvWY/kbUP/oR6cJ3SLJdhZbxwHvF5WvAw4n8vH
hn/gjnTwFJKJGVKf7ifk2HMJrZF4YgOfnE9WRi+K8QagIK66xRYBHoGBdwZn
YQAeBAYxyIVH5rKUvu636Nt1wGntqULTneTZXYFAloAlCrg0ZAeQCTjrS6NR
MbirQ1+A/ZmRlAxxbRL1qBrAZi/aJmDVKBodYw05mL8oG/v7GJcrGkgf5inY
UJPpxNXZrfkWvX2Up+3Nkh4iSRZKKlkrFoKwkqMd+V0ikqYQY884NnjhHQxh
FAh2C80nK2/KgQ3i1R05E12yuZ5SFEGxZ0pvJDzbCsL7rBhxEw3VwHrg+svd
G1QbEq8SvQ/+QVBsUyrVcxwbEIDTLUUTXVI02gll0FsfkjNAg5Y0BC66ep4E
8m/q3abOt7b9/fwsdSH2Ub25jWJZZulEtYRKOz9LVGa7+z9J+j5HZ6utKH3X
ymLRGCOH6z/gHTIiRToyLH/fLf5+hXUM2FgjEbqRmHqnjPmN2O7b7J62wsJd
YOGevZe7tziHok7zMKX2Hibw2YD/cgO5b0FvLrjlKVdQepiGWHUMy52Pb8/W
Httoq3dGJ3lhNL0WOwN8PN3gF8T5OkeO9+DQHn5AIR91TDQWPfc4AaLPRAwd
WPa0SwqXqs8JxMWti19dtV6hGeRpPTpChuto/fDnpsFdm42fCrwho12fdJ2N
fowrMIekZvN270adSOSIbRY7Bogz9QvAEId9nl8eMfk25YcOh0j1SKykkKJw
JXlCSWu2X0KH4N1vRATI01JKKEzIkWcnTL5y+Ioha/8ODNPTjIqgQkPlIIzq
9DUVNBKfaPus7sBua3k5cfOcEjvH6QucyRPfplpVOG4LxpgZQQZKQj6kNcaw
DxyGDRrUvFgb5Ud9O0Iucc8baWddk9jt+qquUpz5YyA0c+DBrTud6Pc+JX3u
9MXBVj7K5xaYzhDxDWk87X0R+PzMFKgZFLANwfhIS9vrwp94c2bEeoEzEOaH
9MvD2d0+TKmELqBwA1Ihz2sFZEIwvn68nNNpukWFmD61DPKnXuna0dC7P9rG
Qu16FIZFFGY5kkQ4NR5McvS8dybXRWXYvDLSu6TRymWZslEFD3ifYFTtNUqj
HXvPVlhms76xxcJ05tuG9RWzQPKwTQdaHhBQbfQo0HemRsI7dQaib8Odb8Cu
YBs8w83ZlzvtFRlOvFK49FbsxlJqoZepA2FffJAMSC79b6Vrf84LR68j1pbL
V8lczcF/uNK+3pQdUC3/LnE+FHeg/NTH+vVAz87cuG/OHBlGd1DiPOOpg4Ky
px9ESY+QbZozZWHWEKZxXyt/ZrxXtA3WgSQ9lPyIt69mtybgj5NwyOlAnnfz
lS5mIhH6/WPna6cH6UlKnmS6k4G5EpEEKcn7xeSnHD9c9AWua9n/jXfUEesl
Gzq5tcEcYdidyAW0zNB6H28ij0UA8gZVckRIXJgMR9T861WrceRx6Konr8Go
oL9zk/LrTw7BEf60fZu6eM1cX7pznBFthwX4OYEnFdBuuEN7DkJZHhJLGAf1
pX/0cKCFyUX3CV1V/V1uNrb14dR4MqoXYmP62/p6fwovBF7ULei9NoNwPjEm
sgu9+h8wYJja+xPgMvxOzEPPKFVNN6hJX8LIIqub9q5tbuUuQUlJrMKXkkAX
6n9okxxWElT5lzLzaIk9zhiVGSYD0xtZr4WSmZhRd4hn3oFS5i5P6J6NcZ+K
LOB9SA2QLSKA3Hspig7ahLoQlHpSRT+h2jYM8ay4tIQ3j35J4g9Nm4TCM8Ej
VieqaaAn+bgTFS2wtMJgG9/vW790u5Dd1ikLBlfpuKBxk9n2miaQOZExe2pM
XLAmQ1UNEXrZI+BRX12zV9KzS5tLpP2Xfx2YtTQ8DlCDe69QO1dhjx6djYDn
Te5qj/kxqOVNTYyxpV4j4AGYwApew5KFSEUd4uSK3cqF+RJOABrbiVsQHHpf
QReEt2x67SWd3Qpx2dJvfGu7rdXqfsgC5MwKaUt7eROIflVCfC2XnYKU20tG
jD9sXDmD+wLaJ7IUwsjvRr/f0IQbYpXCUVGJB5jRwW1sNmT15VLY5naTPWWM
CF8MMSPoXAxEuGjbUBo9ZusYrabnRQxshigQHO848Ynsdz4uSTki46wML6PM
9r7BOpdjdLnLN0sook8HqTivAqcuam5m0/RTrLBPbv25B5A8Cyj/09NM7h0b
meOHNFb3yy/s4uvBdm/oqQ9N/WZLx+xvCCqqdgqo5iFtdQg7saOzT6/LNFS3
firRE6IVrmdiqzDYmaSDQsiFWGmPXFyxqd7ecJ25TkcH8mvU/aM33nqdLtf+
6t/o0Ur7ViTiihN03NndJNbeUdHMXL/sDq5Y6B5XXXvwFFjBZ+Im+LfCgCLC
xdsMHjxmYKrL2AZspEJAx+o3qcByNN/1QX0nxXp7ntm62hxaDnn2l4ffTnKl
cI20H1LG9fYNR9b4Yu/fBnsE1aOeH+kVPfMu7S6aO/MSt+lZ3rdNHiAkMCna
7JzDNNv4guccL2rjoBpLtZ/u4wRt0pjeVnBYUqiKTWpzYB1B78wNzbKXAJHR
v8FYcs8um3bhHwXeD+uToEg0CeKNMjQuZHlNy4ezgK7b+8d4QYiOaa/SOSpQ
we6Q+w44s5+5KWuuMtYRaMdCuNNgdsS7x5pqs/msjz9eHVtexUjA5EG3QeUZ
81kiWIt4Nc3kBGpKUGX68PKuqj/BWDMeXHmYYytAKaMYCKAG+tbm1sIBewjI
1qWZHiFcm4HcEhdZASz/4/ISOiHloudwbCNLnXPN+jscPF+4B9aMi++bCg72
QYn0uIviZJiSMl4V7akVPvvYG1j5WUdxH6N+9Tua9K27nxCwTpqEzLZWuzcG
VRgdoh25t43nzRZUWUR5fG1gqXU/dtgxsJuzrAvNhU2/aRvtO6h9g3gEY7vX
Z8AcyPaQ26uY6/0sB3ZIH5D6nyMNNRcMP9iwqvdbDawj586OrIRGa4rR0O8F
aNMaxpYtwGNb/Hd1R9x0FE4EuxTJdwu6hWhu+RfJ6TzQpii9RAKJD9iYC/Fz
9YxsfmawYYDkQSfv4bJZJmMpMORdniUcIo+1rq4/MEoYHZWXWm/E5dXEV4UA
t+lkC3HhK5X9vZsdTHLBWOH5NABrDmdUvEix5Y1KhK1gLydGQPprJbu87rLD
WEvAax3x+0fQnTTLUZz+jooEITn9zyCQ0biWBQFz96xok3KGP32+zwFDy2tw
uJpCTArTWz524ukswjs+ZzsDjdl3Cp+Hm2Oa5lu/Wg8jyuVab54zWDG85IU9
VHrZbMuvP3DrEMs5DyTgbm56SeHbF6cl4dGIo4DIaKEtJw70/4if/J1hp0LV
k6gobQrLLLypXTPWEaADBwbvPtNpUfRpJjQvxi2TdAEmaQFP8QUrMEA1ZZjR
b0hwPawAqfxhAHrT/nH4+E5zkzZW1ipjdYkzDxtxbnsmTxVbKvXw+Y72e0gT
nzo164x3sYRXLtnZzrA2MgPoP7yB2YX4AEKwp+AtT0wtNmiMvKvjejxNkRc9
SPKpX4tbMiMiadQclncGzwTHUp0hN7FBwTiwyS1UqimL/qW+iCYjyNaetyOU
HBZaREGT3Hwo6jJOt2NKz0RuIhSFUytz4c5aOpatAnH02UG/9bKdQpwPNlV2
0QTL0juL7INrZ4ZX1TpHyiPzs4PwtMHOEoxhIfnbj+lLfQeVR1kozzQvM3dJ
cmED1H8pA1ujBijyipfK6j4nW+IVn/UYv7HhqX1K2nwik87LF+YvLGqA9c5y
3b6JR4aIBxCdI03V1Hc1pFPe4FPZWGU/VGwjO6SkLzA+TiuucjfHeMV+N9Nh
0ZYFc/gRRtr5FMPCgNuxPta98EQfUSlyr3i0upP99SRX2py9b2Hw0rv+eDZg
sTYxN5fBW4BlzzTdTF2BTNbNMsSm/OmxG5lKD1RkllMIj8aH1SxZwG0WdTSL
ZV2lg57kdST87CM3ntS2DtGaeMU1tkJFxDLj/0CRo8+3KFvZuLEwY+DnpzJ9
6m/YJZNuCKcdnCmBjOPBLd6ZaGdk9k3M2mQ4fyp78JnYc0+ZY1oTfrp7UMzq
CCT8cEDhYNP2ckxrWK8opIScSudZH3LWgBuD62xvI1wDFvQ7ilV4nhi6q43t
H/0PMeb0WEyKAwlOmvEuXg+493m8C1VmDToAjLiw5p6JfgDcrfPz2+K6uRYc
/8CfegJCHXE/4KX/q1Kf9XdeEahXXSwfdgdi7SOdiL4zWwrIMruMvS5k4wk4
hsUyM56ouoZRsB5dGFjkNiAYdQ0cVQgavq1SEwtQ0ooqFL2BBbQQt1Hx2fRf
bVzinO5Iujc7AAsnjV+4JQvz/quuMCjX2gs/4cSlnrMaMqUMblo9XwQfsFF+
zAh9JRH+IJI9STXAq5LTnu4xqJ3eL3+Qh3/PqWKXoF+Mh6un3tXJjgdHgNjY
GmUhXvYqlq8XHC4ms6Y/6DIYCqG8YVST5+TxtkWTKvktRfJX4ruihqTvV6Kd
wKY9+tpk5qUtUptmixxFRZnZ+uNFrwntlg8oHoFAqmJDgFL5sNGIbSL9OJYG
0+wPUGXKA8nFXny+KMdJwgIMY92I4YoWmJ1KcLRu/xXx5oB6r2JiLLSCaMIe
Kau/oo6z7ztcPc7L4MtyorQAKlm/HN4jWoj2AlfCLg9Hym9erivLfjXCeVwV
nSEYZn5CnPvD3hMeazZV7Ow1LaKqKu788+XVOM4S0+k4khnMd6qppOH4IHF4
0yh0UZXXjBns5OhHHT38Ot9XW1EbAMdqfTr5ka/XQz0T6ZmJbFlf2upor5rz
xJ6WhuPO+HHsOdJaHqgUvtFDZ/wcUT3suvbaLPybzjONNIyBeL6GRWoZZ7fc
Y+0zkxj23WrKFVsy7u5QqufbIGT/wAy35olYZFl3YqB4nYK5IvV6XdLJIerx
OSULLskNhDsaq7Spxlyzl//7TeRAWD8CoE1DHWR05A0jMRg/cTD7Coarss+m
0YqsXAiwXzP55pdkimTrp+AAkmtehTRt390zoue56jylHdnbs1BZ7+TiOu6x
xBTOWBnJVtBrwQ8DiGDBfVGLf1Z5sHHial+JYs+91DGehw/qqE73LnmIYWUS
Nzgi27fdYBudkFDdlWb2PnoIoq1ydoEG6QeHkOYFjNvuINieX+AjQVusMEFo
WOC3sPiheoIUebs3rgBZQE84s1EAlu5qkgSN8+enJjBgi5fKjgSzhyj4YkJV
pfUQ/BdZtUee9EmOeM+1TXAQi8inz5QqRrc/dgAKIyQfiZrS5QAh+LZJZCVt
uUc2wB/oXyMLaMFyUt30q1Dzc6e39k+lrVnvWlCIC+gDLPKio9X6QC4o0Hk7
/pp/BIXdr0jrikzGhXT88RrbvmnSHQX1/XFDvHjoxjvzrWQrUrzUXMEsnUys
UnRu589FVOigOvHcX6S9BCL8h/Bna5FYZOmPm4w/pMVaGuNNLXcd/n2hut9R
tmSx8VlOmvgbgAdybWBvrX5quyizdEZLHARwNnma/uu6+0defl0DS4+3G64c
FZTvrNvGnqpfRaFHT/bkSKC4++hENioptFgLjfYMzLWbjgmnbWVMmkNTuY7v
OmlXFf+jpPlcfCkZLphy4UIcpsGrm3AjEf4LHWFRsbPx3dvlrApl2x8Bt2m0
WOPu0pNEnOlnGteNF/Tsx3V1RZo/xBEnKxH4hGSvbupkhpBsNvDcBOlcnMrN
WTmuyh9RsgDnb4koaW7/4AoItjkSw4V5ky1pjs/5HhBkkdfHlZDm1uqKngf7
shp9rRqoREkaNIOeasxuwLq+KJDodXAYTOn9TAYJsNSmqEHM80U3fGokV6Tx
3QJ/WZgMPIo6dx1GDAVqqIqpELQeVspqDuiAK3i7JMfYlKn04cFOGP9+KlqJ
c26KVS/LzhBHMh5g1P2+gY7LR9K0MYihW43dWd75ldB6BVcux4kA8JDvYhGD
iAmuoRKXn2Bp8C4zlHTKq5VbuyM8hVxEOUBdKr1gB5EYwJHqzqu73/Rn29VR
qDzQGK3WCIGIrqNn5bL8k9L/qgJJIXCquq/tBT70efy0LBHZIu7p6QHnR+Bb
ivNK4YOB59pZqxr5rwFxZ4XFXudP0/KdeqvFuXMVeW5sPO1ZuI9k6lzqoPkR
BUMCfYAZibrrqLSQKvRCrS86/W+yCuPxv9Ys2CAz7GpbZ8GvpjulRUgqKlUD
LBnMFzGEpJEVLM5tBilmgEGlmxxMgmrooHE+Cdqdh/yjr/7W7yoXldGREwjg
KWBVbNVuJ6PDJSSFYaIK2QuxM/qMaOJB6hXNJi/0hCPBjKy+ZRX8Ww5AVjBF
71AhiY9j9Nu3bxZaJVknugvp0MDFXEv4cPAQwuH9PUMHXD4WFY931Y411IiD
k8fuW9MrW6yG+hsYlFmKRnUYpFTO0LofPTm6o2C+H2+khPgWsZdYW+0w3BiY
DDVbnRqTk8WY1SGvmWPQZuLaMUZClPRop0LHosACP3qPt/BiTJB6V4wJA51c
yy0DF+GaBitF+nnUU9U090DU5rCEfmEZrPItF1DuNcwTJUiDFpwyLP907BLo
+aOKGTogyQWGMUxk+ixQKYOvD/IOKmxDRQsS2DEj3evWs1GeiIdk/wL6Ll2a
W4+ycpe8EzoPmh2a+k2s+xmFAaVkGz9g1Z1zTVzIWutgMJ7vD6S0vKzC5onR
nboCNDcnmx9yRZJbewCn4tbt7SJ15NgHiJgDZRDLs4985XYBgKzao46kY8KH
sqHX5ZwBpFLwlLaT/mN9sI7Tp1Oiu12EcBKwKZmo28GbUYbXi+RCziOhDn6U
tRIWiXrFga/pCABYTuaBxRCVISyRpkiZ1O7HH0Y5HEDos+090h7uJRFfUhSQ
LbfjfxfH7wuEK11tE5X2bzM1UgnvJO3LJ4QycL6yHTc+q/qAMxNYs+sg5j56
vryfLO8/+K2Yaeomx5Lmke49NLbsO7QmIkIHZfebDyHR34Wue49WtrZyRuw/
RpIRDpb/+bpXyaBWHKY9T5Y5yQUsR4TMpQW16TgGYqhdZh80TMgjyy0DU8Ou
SziI1hkbmBmxiY2geayyIKM8KzMgCDCXgWNt6mkVV6/xXsLrllK3uBy/8Jr6
9H2ynoLj01dE2anm2HXGiY79nGEkIWcD0Wl5kcNWWADJUAsArWw48pRC5xSZ
GO6SnikljYitVwI22F5yRq25GVH3Bxw86Xl/HtqLzoFPqteX8NYF5fJNt01b
sFFcUhO0dsAup2qfpRpxQgkPt4a5S1SlkSqnHtZKAcZVlz5aZzE1oWHaHLAn
GYjgcrd7DgyoaVkwrWFt+MyoBUrqir9FYSidxK6ssWWx79Jk/BONm2rp6b+n
p8ql1TaC1zq3uoCx9efALpwzsN5Tn0YCId0JuQgwoyFzLbhE9FoGC1Cax1lA
dl6wJXLedZzbZ7ln0PPdD7wojK0XCI7EUwN2tGOP34D10aPnboaJyTtfJ3+n
LKvlLGKTzhS6Q4tafpAoQmuMmlztH8yEM3XxLx4rNJ6bLMIr5KTZPx5AXsAI
dmMAzsr0WfbN28uw7mGCEMSb4w86UGI8bjHEHD2SZ5xFN3VqjhB5J/zfkTNf
sxR102V89lm8oCdsD+U83nk9EuPPC+kaA2GbjWNRS6aqMziyFyYXSCBJhNri
7/Ei8ssexdxGUOol02BcNkAEiQeR8n87K33ewOHYeM2AmYrN7kuxxYxx3orE
TgmeMp7g5JnWzvOsGm4zPlN9730f9l9UI43cxHhz4p+DhrVuL7D4wIFrqHl7
q7OoCE0HJ9tWDfuN82saSCPqY899FtsTyt9krKN8+WtCDQJod8l+s4M468y2
2DvcA7yz6Uo6LvwkiUR9XYoxZ08LiTN0youNhi21wsC9EbhfT6E7gQL3csIh
90TI1SavgACCQRuUlCzFHAY/lcv6cgTrZMXixfyH36X/UrEFQlLiH6wXyZYA
aCsXTKTCaNeXf+waudk8pnEHbF83I3CkHarSCRcl/90PhUmD6/4otHNKis5i
76PoEBkzApsGQap8cOPzfZCluOaQzPUMorbVcOZMF/JUsXjw9joxkxJZtGiM
awzpw/ESWv0Mdl2F7GTog6dVoAAKsJHREekWwDHEX36clFKA2yYYtZoq6YWl
EOh4KPUdnWFFNYK7ySTCHSmlw+/R5Pvmd4hqP42Ydvw5AoTLt0ShOA6hjobn
sQnnqemGIpDhKomnF0Yqb9EvyCchbK4uF48YM8RicvrmSdZm9gVxjg83FXy6
gtiti7ZFj7Zr8JQGwusFZrDq8AylN10IhcX3AZiCa/7G6VAwHK6EZH07YAO0
8A1ccGwA289sN5jnXkyTsydCBYWSnIBjbo6ZBn/JW+S+xNCNTSXorChmJ6Lj
jOz/X1XG7fP0fpgGILFLPed1GcHVLdyGjixQKDesoCTknWHYYMfXJDX5axq3
ePshaIAcGTCxCDZvwwwjMR7WmfxllzO9fSq1AqKDgGrWThX2BBheyyxvBfDQ
4de1XHpe61FXdzpRG6aR7x8LA2dnFMp8uPKriEqsz6rMBpUJFU7KM8SqyHXC
1DD4Ao/5C5kiG9SH/j1pIwvgp+v+IWhY5SrituPBQn1b2uT/stGKRol4oXrP
Hw0aqQHl1xfswOpzAE2u7qpaNONvu6nkuWibI1m1RBaR3PNdw7bK4ZOEB7IZ
m9E2FzgfwSKqZO+qzbQvMTKrOBwmut7cKBxbPBSXcHfpgcjPtXM0RURvFbxT
5FHW+81Th0O8Nt2WXB+PAt5oY3QZb9ztrXZMhp8oFnK1j4O4B5WWWex4sB0T
V3B3jm8Ml5jHTdS1Q8QP2xMvx/M/laPHuZl214vzfPnfPF9k8bfPrzioBNPj
veUi89AdXst6yTCOuiXrpt0flkPFrRDNxJz5XxcOWzOHtvg24c/0XF7FN8c6
MmSK7A+3t/4OBe2JWqBrzw7vc0mY8ivrYvsntKk0dwlybQ15fA3yCkWSk1Jw
QuOqP7so6d8cmnUJ/w0lc20TzK/5Bgp0A6JH9Ae6uj5OXHE3WISbRStSoc/B
sJoEwIDan516lxYihKaedm0+rMzekRqvcVwb3MnNpfzSDXUMFUOfTFShaKat
yRq8pGRMQJi293rh12DESzequY/Y+XjycRqx9uEK57uAA1+SWRLBtMMULE2u
P6YYL9B1rv4jdZPL/pmhhvTbCIJUCzIMXqzz4xp5fYj82BQQpPBzYtLYAPtf
5OAzu8ycCuJ+DYyiYSn+tEurpn0wrYzBhWBq1Ad/MipVw36hVMa8pL/3cv0V
lwRLHjxnmRvIWjcMZZ2T9SlwB1yrQqQR8GceOPmEJNW55xA/gLCSz5ghZ4Mx
4nCyq9BNwpeaPsudC+QUHw35tALaxENc1Gyv+1YrAM5l3vBvV7LeCLgjy2Qu
9SyuSHEfxrCqjTb1IlD3LSRhkPQKYWiibRVh/+FbA/5li/QBkTsv2KqfN2Bo
K8kijsJaZTRcLh+2agiYKU5EH+8zijlOarP+k3xl9wXAdx1/+TeGFumdaVdL
iP25NGwzl01SyFldW6iVc29gzU1b0arv9s563E0eGX1xQTj6cJMBcDoo/ErT
dOTQesIaAJeUVRQ2jsC6HZt4VP6zH083fWwF9dKtMLJU/tDEVrtli9WAsMro
FJ5Ycw5ojQCR+oLoDbBrkPJPk3EHK+OtXjepeh8ATFRdk347a9Pa8A+V7mWo
2QzsjwC+cc+cLcFxsETeuJjyd5wnn8EqsqMsWzVUZrZaWnpVN//UlingDP/v
UDQrvWR2R03aPje4Kg5rTiFuv+fP5M7mLdBiIJfMQnbnY8OOzLJovcPlXkQs
8obaqzpVHpFgaOCAfOVkWq0WK0W+Gnsz2ZWlMOCEgwqrUyJPDS7GGsjdtUCh
vu0BzZADN9T4DudPWkPx49R66t7Nk4VzTe0Uwq2//5ytNzhIiGDuCo5G6CA+
1xhC2rOqc5M6mVUG0AyBFRUwkxJ/YVjp3YzrdB+uWk1lPP00kzkQ78O/HkDS
u2peJRs1LPXsquZqMK0a9pUf202Gi0BbxHGmtJrydyW1Ns0jM2oH/sWydPU4
7rAy2P2jG3pVMV2rbXhYNZI1RKl495BdMka7GfqnObTDbHEO3HARRNCUF4Dt
H31oiqjGQqIj0HeElJJrJE88uGdrqmBYQTXnRv2jFJIsCXNTA5aU8dLWPuXl
RQ+hY6OG81YKkAFC4+jLL2RtF93xJEJ5NLzQUwOR5Ezt8Rodej7zZPI7lbUV
1/MJQl0vyKCZj0VTfaemF5Am1u2jptQMgiMlqSS6Nrx3pwKDgegR8vLuqoFi
LiBaVAlUpdz3yNu+tOhSryDm/1Wj+JUo4Kmrh0MPQhHCJ0kQEmBqRc/HhM51
nYhSIKMbnUH4wzlxqVsc2518I6qxYeMZkKOmVTYoei6HASwAfBiHKc9fsZSl
ng4V6ngZlWJeU2DTsFK+Pc1rRD8sDhzvIzh6HE20Hn38EPnuQy5BnxIXM7WF
dvnAtwYefoYsrnicfV6QAKVz8fH4q1UyY87PoCuLSFWA/y7G+2RuIw4c/2BK
KZrDQun6+zNFtCPe6mMfGeiakF5opUp98Ga8eGUsNS7KH+KHcvvUaFmNXffN
UQD31mf2PxskjikW0IOE2bZ8Aa5fp2xzgFZqryWGPWFkbkBu3h4JiakiN0HN
+/WmxBC51FoFo/MYIDOTmuhWtcUPSuUmeXvLSkU4gAF7hJvGSSYnKHbVVmoI
yTjQQWEKDiOt3bJItg+FPciwnVzgX6yJyMbx3GGBhiaEX7C+Q1swG4Mrm9lR
TEQUIRXYS9wDydiuXstDr5ZpoFoqvNCH3j8dbXI0EA5DqElOYhb5zFWPdP62
0GA+rT9it/iW5xXqTVV1jXrv4jWivIKuGzLr1uqBL+cmviHyCWim4X7rq+j9
2rD+0r0oSNXtBFAUCwkFOMM8B4FWR3VoTwCJvD7gyePRbW6e2WpsOhDOAc3D
iUJ+xEt13zg17PEVrHctzn2aQGVON59SAHBPdm4OM3B7f9i6wJNSFzMgVuMt
WTtOneGrG/H9PGrwjTS5qHXhEuxd7htw8So4sxmszrTOlk76XM2Ig2ddL0M3
qvmbGjTL6RsSzAuxkC1hyxUVO0HnGzjTLDZDmr4Il/d+hI2bDt7ryGHKUgIi
zO4dhQI8BiH5y/DDKV/kk2wE9cxBV6YQK3kbptbGFXkVmD2U9pqqKLonedkB
VslRIfTWij0EOhB7sUnShN0WDl5JovxMTHsjy74Iy2bITjiE0tfKm7cMRmSx
aw+ApsZlJP4BQUjsW3vtoa48iTKNB14WC3Hg1YvLM3Jn/SsnjEHmuIVi6Obo
M2LUosEkPLa03enCL8khxgswqT4l3hwFW97mvNo9LxFxGpOB9NfSSJHC4sSh
hmblr3s9pEPt+qLJmz7osjSuB4LKoG1zDNkFAzCTiho8L9ZMyHmvq/B/hKwD
/2DF7wyroD0ZTtLFVjKYcsVrIUtnWJsCoWXTYTRsIn8gGpJuxw0+AHLYdBEF
YI3pt97VCqk8+1NFrCpPkrfyORIlNj5bwkQzth8m0tOBwhRoJ3tEIWhJ/ydW
HSMFjC15UFi8TwA4AujgNDr7bfq6KIUzjiGADiGrLozoZuy0lUY2H1Zm/uOs
676vP5wYZ6sNwyRhrj4/y8flXE3CnbnrPJTUh+mXRzF9AyY9l3iwm71XWukd
/7ITHjExyU3CJVTlE5K/bqvIqM/6uSYfvGoNs1HxG6lLGvGtW3X12d8l4nqL
iQV5aEr+ZbDtqdtUE/bpJuo1Xgv4jzGN5HhNFB6PdwlBNBZdAaswFRlH23bx
3WIoZcluSFrivgu3GURJGbudSe3lsHIQ23Hd/bFHqVg6WiGIUxPzz38s0NT7
wH7sd/qu5t39zP6gon0E5LcokvVOfmkF4zmpAORo2raABt+xpHBiu6/IY4Ov
XyeaXxEKXVtGgyfMgt+9Yu/tauaqD6qmy0HunsqjU4WJ3M3t4q/wUGtRccHU
dj6h1Kxi3ozniNMprk2OT2jjiXXWfHoEXz768F/lKb03c6DFsEHxUFQv/kqM
/g92I6WXpnYqDSXlfMB+kcTftn1pA4fpxIONaCQr0VFmz4x/uSPylqb+/xzV
xNwggY5jpPJlaZFpPYpU+Quhc5cLsJXfR8mdJX9RjAJn4tFWDAQKITUYSzNP
s7DAAlhroWYZua6tX43XQTcpDH8dkJUjeairi8lWjSU8WIOm4QxRyQ6pthl3
2dVZgp5P+AjpOR4kpxpXK1l68DZiWXWkYuhIUkre04sJTgNdJhNwiBm18Ws5
pkw1vGi2SzLpA6B+cgy+cvi7MUpNOelrWHIoYJ3VMjUyV27Wd+1+Ec3nP8ur
zZ6QKhq7HAeX9qRS9DSYo/k6EvgJlNX2UzaonOnXsAQHvZDECqsz6KEJ24r8
84xeETTvwDyBcjh+5hI5TgyKNs6tkTvn0hXSj1h3NDgSAcQs/DpL8MiKSZtl
JDGkxaixzEmgO8TtVwOQyb+MMyjGf6DlZ5uktN1eIfGsIH5m6kopXiN7aa28
X6kbR4gbOKafbUdPpzP68bvfSL+0xJP+z6dUB54J4sV/u1gCbJlCZAdFQFDN
UivxAJvapTWNlM62Eb3he2rJbboBflctCR83VcM5dVKkOIfZA6io2eAs22QX
hxXFWuRUu5JMX2z2mDOR+W7Ih3oTG1rGSw9tjpWU7KXs6OvDn+a9n81DD4eB
BGrnDypkqo14ALqoFJ6L/JVximtjkVvm114OGQD3RYPMRKYl5YfPTRpNnFyS
78l9nY2GD3uZaIdQgbtShiK+8LZkgZ746s4O51VJ6zy2w9poZEt2xpSf7eMP
WZDuXRX4F/YZVtjQuYam1ZVNjGCDmy/uTJxTzGtTmOWJCtH4XfJxNkv8NEbs
itPsHVmpKRrfDqieccc4QOWo9rHoYT62O1oR+CH2LrbcNQ3RUvl1vagF4hFn
b+JM/NeE+V0vUp3SOBVJfUuVW6Qa602FC8BCO9vbP9ZYGdLQfAnWVd7beJ87
ccBx1qZRT7m0P3k+IlPfqLbjsd6AB4EcJzMhD3mW6sYuss0N54tDhp8Z6w0r
IW5eZO/g3bwYt8fmsJeDLLdB5KUz0sap3KqorEybkaTWcxZX/DjminVIZx6u
J+0vA0ktgv9U4u15MaPORb9RbKFdmRaNgN3l95nQ+l/0wzBnwGOR31dc2DRD
1tcQYnYr46y0PoCovjR7NpBGoYZBdnsrzVIKuWf52qTah+x0dAMJWFWhNuCP
27uGVA+k4hzftwuhk8/aOaLJx/1OF4GKymCmSeaHn15cDLntrIwrH9F2uOMW
szdODywbQJCXEXqP2dQeRdRx+SfQQdqVJc3mverAsaIxp1rXoeWJ7Q9CNnKF
lJSfIHNin2QmkQJg6+zpVciOUsC/BHXfdg2igB7twZEUUkucqs0+/isz05Z8
OYYtyBXT1Hvl0lN713msbnAhMfHT23ohyyU+uBNiaEwLM3YQ9QjrcvSdJyaU
1QooQEY+/SaqDGpFX4AiutODeOW2ifQlebNwFGg2OehYDmT/X8qpklKIMKdk
hHY+zjr/Ru9UH+tIE+kG15d04UB+m9bIpotgp8cr8VfeGF1hoZug7QQlF2HL
rhw09F8UFHFaAIMOsOjJwHQnjgi98s/Ls/dbx6PRcIB2Oh9P0giCUGcQTxuE
QacsLbhimw0vfJj9NFUYM4ZHeUKLfGxL7th1vVeWe2q1gIppTUL+slXwB01s
4TN6Oo8NqLg8VRazaZO7iEypzrGBnexJJv8qV+0rO2cBik9bG5ldlLw4ROc4
69ybgp7C1yFNIDnUcgj0+cdGIt+O8vpuZb40VPVn/bZOTZpGVcbJicGMqG9I
XE2pTDX+r3E/SPLpXhoU89GWa74z5yxy0YW3y//19QMWn1+vB291aoG9QFLG
rHE7XAwm9SXaNHJfZ75M37GKAN+h2802OZN80vlt8LgoHm14yeo+TlUtaOwa
9fYIO/Yki6zzWir7E/kCDhsUKAPpTTOGQbRX1ftitEa1NDKHfmVccWPexbzC
wJcpTZY3irtu+a5+im/BQ3kuPfbBFmHjRphTKi34TDAGrIj108neGqc9zM1d
dd5H3jQ86USh9u/AgPFb2+2hAfIE7lT3OeTwQk6fL+KzLneVB+s0mOpNFb66
7PLPY3ypmuL7IXLyO3IG8o9JTp4+mNbWy/621U82vAinoyMgmnDuijV12fvB
HZlMTKzQvh6hTI9N0G3NC+c0NJGdOnRAVcS66U6d6c+kcLg0dksuX7y649F4
YIkK9+7MyinB7rJH0yCX/pqeB7OIAYbV9QqifSWsgHZ+is64RCShvoAceVKQ
FLXDw1ZYGz2jQWwSkxOsrDD9bzs6CtTxp8/vwXkKrmQhrV/ilABo6cu88yZC
Bw/YhwUJgyJU/dPfBTH0G8AycdRiZSgb7MTvfCHpA9PRxIpRghem6GmUPgMS
Tafsfmwa6dQSbK9Eq1GWT5uKAwprboGOtsDsSxVEhTT0X7BVjEqRdf0ZT5Io
AyEKIeZnU90p3kZOXdZCeQzPKqDq4StanlG37EE4/gYeCqK9/ByPnhihjS2+
mRKc391SBKEBcDzPxQzDeTsL4fu2z+CfQe+C45gWQCttnRVB5EYLvGdEQqHf
BLbQVFB6JKrZ8OFsCYGm1/FvXXSuDQdyLLaT3PAfa8uLXwvqenR+WTgE1M5I
rXDivyoom99cZFL0hKWkvEJqBPNfKi0w+ywYUtBgeCia7Vvl1h2Omq8E4C4t
r82XHIVvmYcnHJw71eHfTLW5uSwOP7MdEbE4FgJFpEGCBKGhh858eGIhMUj3
aM/goXV38S0oEO1lo2O0/HLF8p82Cli0I1x5sIVShGekVRWzfqQh73PE8ENe
4L/YhHXTStEixuy8eCXSEA5YXKOJKJXPlS01N9v847bAqR2QgTtOGK8Gfvwa
lgfFfzWa7bHsQsNvQbWMN/UGS0hBQG4x9AQBnpsyDCcHLUbUoZR0tSIygOrO
c6Lfl8U9/V7RQcr04MHIAdbzeUjTuUnmYDfExtPc8EYuAXAYCTZ3jmKOwKzh
PE2parknPJ3NH2hve5dYkLiyHYMw2O0ayhVGHZl0hosgvK67XkFFpg00MpE1
pdvhJqV+VNbCSrbkQYVS2ogvudLRUlnHXnrL+XoCMU7+Qa8dlx3jIehaKr0O
3wSHUs5q6DWdlDCr7MRdPNTIQRRXi1NxMmmCsuPwVcf6+c8LpWvorsYGLVYa
3HZB8NXNc+UT/eZKOkdC1P2NSneK/lfFwWX4rXdT5gOO/NFQX3TAWfAfyoUS
T7FlWCKi0T/5sFuE3+txGUACnyMQb7u5XrMnhEEmut7vkIs+SjrEG9DaXTji
CsnOItgFP13DZqHsS9OJb0yCmKE7ziDnp5fMGdWof35qi9idoA3vHj9/ra7X
jqvN1hLwfk2b8zeOrgiehZeUUlK0Vq6aiau6haOBP3toFNZCmhdxQQBHegXk
neSytfalPeJ/JdNkep1z+/9O3kVY7K/DZfYWPdAy985vFing2E4NDyNGe8XI
xvpHukGEpd9DprJ5eZyTpSOh6HzTl7U1OVzyXf2oAI5u9/k7foxyP7fi0eta
JN2cnU0Zb6vjwAmNzuITf4uLFtitaK08PcRbD6OXPvEOxDAWMH4k5G5TOz6r
rNr3wXZTzOUMO9rPWSv4aLMJb3wsfYYt/cisws8DJTfNS/hIjbt/Lh35xDX+
SIJZRK3v7CprwhOBnJ0eAC0rCcU29AvNv0VmDLh83VXcN4uWt5fIwGB7OJdb
rdwZb1cnlvgTf8w+Y7iee6igwT5ENqnZ27kSjutWH+H3ca32N4BN4s1WjEqD
L63SxHPW/r1+vMWzU8/M7ODlIO9w8lYB6bdiHTlk3/Ag44EsN1g7cv7rcGgc
WgrpHp4PpOcjASX3BIY6/ZlcNDg9MXQ+GfqJ5gEhn6eAx1+13tyKdtNOgxEQ
7o6zngzrsPExA0MrfRU68abHPLcwWSI5n+uhlxGLdDUBGxCqPyZImJAERKjO
B+57qAqhvZY/HnL+ZDkhtueJchtWzOkkkQrIW8COjRWLwCk6Dfe/bwiL7oKg
3Nlkpvj7Tr9lnr0M98QFSByb5CjdQULwZMbiNAiQl1enLdl0eAQIuYfN44nb
S028c/4mx05c7m4Onksu39/PYbGyencCw+VBj5t64I15KRjVWZr7IEzUHiRS
8QeWoXrI3C78abszXy0ntFS1ekiQD4OsufWwv/wDb+IqVOyLMCRNmhnAnbNv
QMcXPuKfTi211LppKr01Kbyr3mOJEuSLSJDz7d2wDVJG1oGlMSgFq9rF6S/c
tH+aDAyQHoiGYnxQAdaTpdnZXlZKyka6uH8bK7tAjhY7nMORJ5b4ituP84Ua
Sx3AnepmjPV+YCLw5TIV8+KLGHwKngKgNTrprPLrs8wu6bk+et5ofMYgjG1r
uixAwrU92KR2HHYCXE1b7yXx1ZOBnepRDUOC6qbRb5v7u9QzUskG0ujvQxcw
kZ3FARavYUJItv7sxwMFW4dV1mbG1I5ju8qfRqL6U4bTrqrZFoBxW+Xlhz+U
LYPhEnjw6oi0DklBRY73iMW1KnPy88YkPGcKTfjn3lH3UgEKPIycl77MKkIP
dD6T5jUyNQeoOGZ0z8oFhCObaXchC1p1sUtY4JMSX1jZrw9XfWt2L8PBHtXB
K4nVjb5S/DRrSFtml0vQF/LKByELrdHKY7thOg8kMFzzMlLEWA1g6tXYJtGy
UNwN86DE3Bu+2yBK7UJmkQRH4H+K8WBZPe8MIy0HCoeIBYn+DdXiLZaJZegp
FdAu3jfY9FieIufSC7MBwlOvtGMTH2Orzgo00SZl4CfNXU8EquQMhDxrDlJN
JU05J9zJCMMLlsJ0ZaEZox8HpNE8JkQKtrndSdQ/zR6w8lj2Fm8Nl2Nmt4wi
6JHxiRgddTRgLYFfjEdDNE4KAzz1V99P4ZJMS5HuoTqIGYkNxO1m33PRbuJ5
Dr834/kZ6hiCjfqH+BKMa48DgHQ2iVRnQMG4qX/igZMvcKHgdSTk5J1zzJ4K
kO1NBspuKf0oZc0mH6PfUOk2lMzfVx3TNlVjuNhRzaHeF9eXWOFpgD1jD/4g
axrMgb4lZftz/vSiN5t3WxlXmg0hegKPO1UUjj4FKGdv7ojVkcoqhH0tJYo6
PSCZ6J9JSIpGkNSPq3hhqp8ftOBHsBd+XaOvv1qlKWngypLZXBDQb8l0v77Y
kN14KTRdfl1aEaUPvttocedK0OGvzRg2H/r4F+RlHoBolI198kzVfG/N5tdS
1sz+dljGUYy8d1w2OhCPszY2DF7NRvJXVROghkpz9UVO5a7tyEXli4YH8nWI
rZlkI/l9dtdD/o3hKfnW00KyKlU7dormpxUD1A85VQGEXYMAym7GdDMkWUR/
dFAzCV61Zo4UxqHRaDk2hPAX6n0VwMsRQNA8ZVeM1w3Q7UGz13nPJDrM5I/7
ApIjgYFkgaJOmPwRJqoY2Rq2DSh6cD/VDZAvdf84htSq9hcS8REyR823sQas
JW3WTG9KKgKYG8OEmkOAUifn9taHdBR0Arh1TqsduS6/eBMmaMmff4o1m3eO
SGJmGYmJT2kyC0OzJT8MMTR15Fry5Gmt9mtHwUsE+GojcOLCk/G/3bgxDEuR
n7A7GhVL38lkypvX973fe1WvP5KxYAG1xlZOu7jde3Ip0tZ6ijfiHONpedi4
lORUf8ayh/a2yxJML9ejqY6JO5kPF0NwzgpmFSfAdlyqrOBYnhpjq8POV4mQ
f58mMunjqF+A9p9QLOmxO4zTMM3B02YXbXpjVSWXU0JPNfT0gvr5pYGswIAh
kko/bSncvWO+AnyaI19wmaBEk2krx4RqhAlHw4wYIcVIB0mUnNu21kpCdlrk
9ThTu9VT431DwlhMkKizVpSCp2BhhoTnvaYC1C33mBeyqTLJmCEhpIpjToIP
NjEoqHvPPwPLjIwdtigSq48HEKAESp+t8v6LwctB/+FmDAA0cFaRMPWSkkwb
l0mB3fwGkY2My53236XZWnau/tC00O0d3ZKuXkH8H/Lom825qx2+FzsnE8D/
LYuAmVLa0zc7/jyGoiVwhBfdM5qumPwuP0ULzkigj1TxEFzhdeaOBuC1zGDH
KrSImZaigBQC6oD0vNhLaG8L9KEkQVH15EyCThZ9KNVqyXmY1TmYhUG0sJgp
mePWeVC7xY7Dq0WswuqFJQNq0DYo8U1Bx29dbaJDMDS8wcyruOSg0pDYd4dD
S0l7Cxm00Xeqekv2xV7r/YoQLnVAjacs2K5OqKIinVtz6uWW1o4/kcjwmJrr
f60nTE5OjfARaA9EJVxzFAPZJxoBJ3TUUzVDgJhWElKEsr5lTyseEql7ctHj
4T5jyyJIxQH7b8zgw4nJB5GZ+lFqZd9yGg9KQjK7eCVcPau7z6yWc2hhOIik
jKPg721H+LDdVNvoGeodxwvcyphEqZYkncNJZJ1RRkYVBkS5pyCTo6KPrs+j
9lKTIDANKTBwXtZ/sAzvaGD2b9rSAlGzuVgD+hdkrgPvBzXjoI8u9gEgOYNN
NqY3eFHApJ21u4gssM3K08czJHhToKJEjJAu9YkOMiphaYLKGEPQO0fz9/pe
nm/K2ZLs4IeyKRv8QGRpduiH1Kc0TqGsKR4bI/NgnvrXbeIVATIpKiqqSWac
1Wk0/XEEu1cRMz7VpkHrbqDhuhaUxpCp+CkJ9TMtosJCZb/o5CFZiNo3aIiD
dc3RcHGJJoWh0Ni+iTGe2X8WfLGgTcWAnz/10VfKn6bQgiJynDJpQ1Ow7T5Z
4V2SLyyHLSqIN6ipTPbASJspBzbh/bQWcLqjV9LIWZh9fXz8Fq/CSsKs0tLP
RgANSA4NHybRho2qqCh2gErzkOjj1Pgw2M9wPxl4/UrkYbHkE8JUAR+55FUE
Dqnd5ZlISJeRuWRyfugvEJ1QwDLekI56zEHkW6QD2+TLknsMwtZ7xgt9gSvV
TcENoD5sLwclXqhUVWg9isAWPUBgrec6TQkPP/utTRWFe6+sEsyeuJsD99Nm
ckMtmNOQlJh6sb6B9FHZWeaRTu7QkTUJlbbn3v4U1Z8S38Ek3O4+0j3OCe7P
uNBmbav5wqqB67o/Pq4dihp3mKcSDSiq7QbRPmyXL1vg1uNvK61vE14u8kqO
r6ZmjGR6aO/OViGJ0B6C84+kg2EbEWHuYzs7uLOBRUy/JAYi/lFtr9kOJDDC
qWrGaFvdpPZwyo10o2hFA1UTvGtxX2YfH9SvqK0qzPsbAiUObmSi7dNUxbN8
6PuGoDOI59NYm1yNRo2HzN1eNZcIqnoBid4FZiasWsu/0CbvDr9kmiAKSUsq
pV7phjI/1bnU6s2htXAvmGM5hd51t7cZXAxSCc0FE9yKlBVXXons+MWqZfda
0cpvee3XFAUjC/HgP83tMoOwE4+HqIPvxQ305C9YKvg9a58Y4X3jXC4DULgC
zlUf3SD+IJYlMYy7zfsbnI7PWbLRw1IudLJU3L+p2lU/J/erIbaaooll7yiz
sBxweN+kh106u2IvtiaC0rsX8qsgiHA+AVP5x5BcD03vOpaRPL51FAqhITMl
6hQhJmRaefpx71SLRzhwF4fZ9px0ln2QZ6fxmr/zPKadM6Ikf9ooHlrruCF5
75vmyxzhhYA+PFc0kK4BxgLYmHpL2t5Z8GBdcQ7zbMeOLTqaUbKe6tEU6+DC
7JXiEoSP4owXwI/ZnIaULQZO16PXxN2LoOgder1iI5xcScWsvgrinixH3xDM
yqYwUSshbUozXNiol0qPA+TlODN8DQvcLHc8IPy79eZwiTGyAY+PXSdgWKHj
Mm+8PCiAebeJ/2+Xi4Ue37P9hdz0jTt6SZFjH3k/bzLuBK8IPDQhoQfHkq66
YeSk6KxscrilFGU6kkn+2E6bAwdS0A5skmLUYtA7j1544WJepVEtwM7oadgF
Xj/4xiwD2cpdbZEnfGc6z4zBljdsZVpUcXlxXG8hDbh2JmWvOUSmJ5BiOGWY
iRFtIxNfjCsXIIID952Pk1CSrWO/oMUaM9cyx/jiNwieSR2Y2GXATRoOkNA1
w566otXqvUsWeMFZ/0u67HwJZJyDaNuuVnhfMBVT3+9jvfC3a83JNXiKGPWi
sOWAEsPfwZgGDvkd/vzYCs/Z4L0pZqCMr4mHbRxhcVEop2L02D0YKZMhycQu
DQr59hBVrcuXY5FvU2MpnZqoAfzUohLCaUC9zugBYaBIef8dtuImCTNP9iEj
8hfW0jtNxLxVfj2J54G7cF8TY8LgEKB29oEECHhqtGDUw3YPIT2ZzEFHW0BJ
CPnYu0hBhpFHw4FvhDHU172VqwfmFMDoaVBw4FEomdpasCheerpzg5YyE/Eq
zzEn545fVizZRpkiLtSOvtCDQChjRGEmTZv3iTmM/9csh1M3LQFT5xVQFVwT
nJKMxmATqw08eaW1xZrrBtZro3s2UmDfll4DR6Hr0Xp07aech6LUngpYoRnD
n9O786IOmc7yaNw93GLCIDeCREOYZqF7FA1ilj2o+IiT5/H2NpkSIQD7KD7k
9xZ9VhvspJWCmRb8TdArDzq1SYhKPQLpPGYakE0JjbncTFp/AasMzoW8Q4uD
JzQfHTi2ocq1NbJOQdOcIEn4o7/6xmfDHO6CVOniuuccrXcgL3ntgHNouLix
oI59uYWmMD+l+XuB2Rd19ylPVQ6ysc9jgwaoI6kY7fvvx4nv2xOuc14Z79QC
p1uGr/e/p03mO7axpH9OK4MpuPFM2vXXDEzeZFZ46dAZD2Gb+rwFpe1695Tt
bVKjKRjItGMiIYLDpY/EyLWilRxAfeUfDd55qKhRCrVZJfMZOUbuEJHKKKzC
/sDaxogQGsdZMen1GjIgXBCgwoH4HdjynxGHF1ABoMoQb5EaHzn5Dj2dCooC
+2JBaNjdVUTYM8YG4Pg2ITKOmjhlKaF5cuu8b1KeuIKOXXqTU7eNT5gc2xtL
z9YZIMWTKw81/kognwwpFOJbMLTJ+fG1t3vPGJYwcXx2W24DgizbfnCGIj+f
H00wJYgltZXHJSTHKF1unSMBcuI8nJrec82IiinN/DR5MIcJOFW5zv+5PXa4
VE2vwqV6DXHIn9jIj+iCbBwmq9oUUuIEa119IyTa5tD0/6kn9fNlrk0lsOEW
fYQ8Mo9mKRB9slVpU4vmKeizN9vPHYgCZrXi3CjeohI5iwLaZkQmh1phiB+e
1lF82Gg/nI4GzCz4GrGsRiVQUAnZ/ZDeo1RZO2T92aYBWQ8uyyNZw0ClxoW7
WRnyFPTMZsRk96plXSALOcfcfRppjsb681SFBmSenSWZ1IbFnNqNpBwXHwB0
z/GxGgMhejR5njEdMyieeCCM5O+fvvTJUNF6wq1XD0dv+RLe0uhc6m/EiZp5
yugOYtMBUFs2Yge/N1d3Ikm27H8PhgHYbpnl3aO48gu8j4y/NlMB/EEY31MV
McCZz94dCL6S9jpOvzy2OGTzLZ1LSzm0bG1BQ7/GcI3o81M4HZvXj9BtfyK3
b5Xz3neZsTTuVOiFUhBKmJWWKqfia9apEjdI7vdFgJ+p2icVKiAd5lkjjj/E
gw6Qf/07A7aB4YtTMTjX1Adl0R77X4vIysjXalaw5Q6UhO90+6SIQeJHedmX
Fb7IFRmAZZBO6+J/WFuS7faEaS/XTNEQ3DJeB6MH0wsh3wd1BUs8SCz617MY
clGkxngn1eS3gNH2Z5vgIfhDVQ+vQPtgIBHLlVXRNR4MK+Q8DbFY0k8/iMkO
V4By96c3YckIWeZ9p7bKHXGUFKH8DNWiXAVD0rtokuUgqJbNHkWok7zBDNMw
FNDijrooIdLW4Lz5Q9oblpryNOWvklQj5gdZiwfOsjkVsb7mKwx4B7T3wVF9
Iap6sZwkcvO5hY54zrg4bk6dI+uSucZ1oRBknm0QqANAC3fHjjkfZwehIfYd
5LdGy1BSZzAEbRo/hgsz5mZeH6WesnjpnmEZsLOq3+/9MSE9WpWYtQic3VvF
E//4lCiFkfI8u038Q+FPn/Up8LkwjI7AHFOCyaecMm2kxafbzG2cRG7LdyRx
7VtRVzthjnqZEPNMOEQK4hE+R2yBzZwLWytVmq+th4fzm+0orBRBbSQGUUtu
WN76ocAuNoLp2YBZm8JI1E0fN3uYB9dujr1BZ824Vsxoqh68w12JKsM73rsB
+wGOPLH5F96++P1g3Uaj2mWjhY0qc8lpf2qlDkkJJS4bbZ8wUhH5A5Xb1ZEB
vO8iXFQn5OmItR2aQrwczUP49AJDaygm+Yd6ige4RuphDVzKAWlFn3wzJtM0
75pYTfrrxZEtcdmtrPJqoi98XLJszkNWzRdBToTjbiAfWnTe8yxoN/CgqhVU
yDlHLra4kPRFWFdJrcVO/vf+ee6wf1Fi9YnIuV4AkSAvMzkTAkm5EFS0MBoD
b44d/QZLGwIRc1wEoFaGbpNQubrEiasoxVtpZPuhsk2I5h35jaTGg+wJdRJd
UfxDfFw+/KNAuOuwuVJHBH8AHEg+pkPFVDiZY63yCb2rkcd9f2Nzze+QmRB0
LIhcrG6c8S+ReTkQVjwtKZEn5UzEQ63l6aqH8UYjK28Bg/D7MHTZrwHQkQ0p
mDh+Xpj6bxFxSd32kE1hNrNMMWvVoR0r9iGZl3BvmK36micZeuOKFP2jPDdS
ZF4bqHSTKmUFXw7WL3gGRpQKJNMnU/shLKqYlbyt1Ejk6NFVXizL8TpvzZxZ
JqMCtmzIbX15SZl6ODX7h7k0YXjYB77btvuBuSecHEUJ7ynW8plDuqQHW0CH
hLCZWdf2E2UaBTYgb+cZh66ii38NF0jyqTSRsolQYNJCnSRjST5FSiqIm4e0
fjl4RdtoyZeU7YS7FG8NCipYV9zxlGJXZltqiZ8PMbkrJ+Dp1D6Gg2Ly8BbL
OFNLuijT3+Bw2gM+G5sVJv3epD8VhkzzNy7WnqwJjnFX7cQw2FRm9l40+ARM
aYaxHZFhdTAybzj5+x4+DfUyZSOtkK4b58K/AE0xJ4SjnWkbBIfBpMwutBVR
2H28xfvqhjHEPVRvROYK/vk9L2TEBKbTWUg8cNwyBNaOyL/2eJ42W2bFzbWG
GhanZ5jhUFH/4aDQbApcaq045AbaA7tAvYC+Tkxb8kRMs5G3Oo5bTSOSgDGx
BfQOfz4HBi1AFrz2Xe+YsgvIwUEPvBQh2BVVGpPx5PGqCXA3gMoh9SaLKXJJ
4E0RBV+nSrnJVtnpCw13pwsZWwAUyMSFDVsaRSvgyVYcj1QflQezlJE8y81h
vTFn6BaGTa2JWSrl8Clu31u9QjdifADuf7VlpKzm9CV8p/rOcEO9wVlHhPRQ
/vhA73u2e3XWKjIkkh+5ll9zNyi83QIYYGfvSJR2LzEBgF13pLyn6+TAGI0H
qKwiR1jh0P6r38DZRxmXktBfk7CbrRz4g9SGeZLmHq6zNi9SiFMRAgPmOnN0
yv+ddFCNnSuhMywJZk8zZGnMka/H86jD605JIBBecTh2X6lCJMhBbmVCKH8L
CHXImgK7tLY31O17PFQhQ8tF6OaUxtarxttoRikc0PKLMLb6Crg59ssyK0GN
jW/Pt2g5gKSQ0/8SAaJmZcnYYy8aAfZWwran+p9sVerNaG9Xq8mq24hEXvZP
P720ENZkyKNaWWZ0imB8ytxzNryL0WXXEfABWM28uepbZSbx3OJ9wICsxE7K
xQ8fs61oZwAqMgw+O2tZ+NT+423trkyXzqpmeEat3mrnEMDrx2DTMVO4A7lz
NKTJdLHcca5IPA0KmMt0uozKnCnElaFdZ2yvDYxJVQJYAoXsKiOvW/459FO8
gwaFOm/0UKt5COQvHyJSNFbtq3INUe64vpelO4KLApP54wCeR9oKlXIQ0EYw
PUVozI7KzgYDUCpkMcvBHXxqiSz0BBl8eVqxFoHMIAQ1RuNSNDHgcNdEo/Oq
DKCPr/BoPLItm42vxvpp/EBGOlGMEoE8NOciK2U0Gi/SjDDR2QLvgCHx4lXc
iB86DUCA/tta69HdGT0AKY2c+SgQ1VkzKQD80sBQI0RpaQ7iSVr2yYJa3do2
RUmQNmTg2OoiKHuh1/ER255pPromdiueEvHO+55unP5QRZvtG66prT7lZXP4
+EuPsCeR1JNu2JJdwOsFQfhVNaVMqt7jE/a4ufpqXzzqivwLdjD3naBRJUFs
wPz59AvogcEXnD3IAMLqAvcXvlaUHpwzWkvNkTvyXRu0Q6kNPPuMYQ1GPRIZ
JfGMHv7XJH526FVEMYg30luB3+9Xergw9sTaxJmt4/nUXRq8Xmyyn/n54oCK
3Ih0rM7tqVNftm4YxWfZ90m3xziJnIrfPqioKQUabj0PSiWEvZpcV8YLtLrb
U/kWRc6gC0APfnkhvZf3QTDiKGa0p3JHm8yoGNbnedTmh1la2Qno8j77/v56
LWTkg7vv4uqOU3XruJK35IIocw5iH9iecNjnDi7nyANxGZh41kNFpYuQD7I7
dAGyzk8xjD7FAddIXNpA9k9neCqZA0595iS5d2E/PAhr1XqTAmDsBydCjz9F
f70w7XzXtazQEtuJhVnuiT8/wUfdK4/yxLU1rVIgTXxPZvYb/Ge+4YXmjTjw
bidcr8txuEakRkGIfMK/f1sK1Pjccwywsz51xhcAfuzZ37DnD0q+aCwb29vp
AgWTPGNOPagImkVVr1Ra5k65QEmvY4o9r8vZVvSqtdWzij3hdqVRciQ/7fKd
ACFqE8LnWxIJSGlxCOT/MRchkE0M1wlsXZrtKYdyTLrDdmpw0L9sT4nOgTa7
W/ftly3VNgMATxdVWbOUt2/IhRXMNPKZlA+giPVnKcMW+RNaOOB2A0zQSjMU
ZdrtdaC/nv4VHcsv0HCa84DG2rAfd2AqGQ8F+pQvBz4Ie51iSrH4dq/MLgv8
Jc4BwfBgXYF+7zlp6rwoOHnqh+FIMEP4viEJDKjfR3/LKVBbJU27NgBNLPyW
EiWmQrZqWvZCi74RjC+I4L5CMzXX7rNBy05X/HrLhi2qOQN3ZqM41Nr6GdKI
wnBwUXBSW36BqZ9S0C5+bYwZU9drDwBCGPZozd8iTRnIVgUsa8kNAYQx8xfc
O+gGgKTHt1pVjnUcchlXSw/NGVuPgAcsLS3p5ptz6ADlcc3YC5+/tH3WYXoQ
/fYYqs+uLUCIP8AZ3L8oGRk7o9TdZEPlOBOrTxmcqEYtyO5Ie/o/zUW88zk7
lUUvNwRJig62EUNwspdWQPgIYCDTQSZbv5mjLn7sOc9IGBZ+LVRItXFPK4PM
QmGmKRCz8yL9bzlCjQuG3yzWsP5hebiEn/bXpXJNuLGEssorHSQghV5C3GPO
ZxxiUDQUCIcELAE3tzjZ1J+Z7pNsCAwM0ikrY0MCx89Jz7JS4zFhPYmj7Ztf
/bFpnxNrID4O1JuGic0McpsIlKr5JAcZH9ddHVwdJRDiWVga/ZAf7kPlh/av
w7rqVn6OmDtKLu7xnYCpe/eJqvD+6sEhxChUrpUttQ3R16ig18yLPP1x981v
9ZwS84cvkrJpvinMiULOGUR4GaJ5fNHh77DeVwXbjtscKlAclqtCG5KwtlxS
hGuby5lt9BDzI03Nl7qM7sSYCLNPsMAnJ7eGs/BSlwjoJOONd7K+zco8ym/l
oYwOLcTz1CNYi4M0TFqKjoeshDnPDoYyZagdTS5yCLbJcpulSjZJUXYuBxgF
/Z61q9UEvrW5H7Be3uADPnz4LeHf6bImGcuW/vYzn00ZNEYoWhgrOzvv2szE
d0tMCn57RcYZihLgw3s4nLP6fbjK6ZZuyOT4dtETO9S4Ruas94BBCnlNofVy
17XW5BSv0ZvNfCGVwxi3TeQp/NolrxsoM9QGSzvQd9MD4bqPiN+D39Bg5q2c
FOEpu8q5UuS3sj/wTKe9lh17bJS6PSE+QUONd9ROMpEgZp9Gb/7XtPop/R0Q
d/ATcRePC2SHqllTnD/xJdfT9I0gHpIB6yYCahT5lAeqFGPtpJmt2atIWcR1
FkU5uXfZmV26e4QBMOxVqxiNAw6m+Hmq+jBEDWNpN8CCsrxDH+W+qknnepNW
vtbJA8oWzkHe6IvSrLPzT3XT+pKFKFBO05RtlYHIl0EsN/bdbul5arSaB+OW
76wfcSjWSp86jyCe6kbKYp5PH2XWvKoHE+vhYhW52ycdi1z+MCMQjoxdbbhH
Fm9cc7q5h+LlxtqGb56HQr/rY3KOIly9iSRsuATrr3Q8bFb/OE429mNYUSlN
0M1L3BIb0UoicpdsTZMzLR+AnDXIYAnQv54Xk8xEv3JxsvwIWYKlk3BjH1p2
YSo0yke0nSUl5ygEgBQoGCPp9oRhMaWUot9COhVazesR+v8JiPm2oGUPaBq0
RR6uieBOporfWuVHLiESBwD6sZE5mrzj18oOourkX4hBPPbycNL9qYbP38ax
wCnnsL99siQx+RcUGt0arqN3jl94FRf/Cr5ucaxGsFB+PHv7zygPSC1AWPnx
jIg6uGtAGU+NA0YGeL1uluVPkt3Oiv7v7Q7uj0vaWLotSnLvXsN6rWGXShhv
oIEI1o6oxPicPSOVkexPbG9rfhWT+IdDkXUZLrQBAaSAx08MizAm9nIAXpHB
TGyxRKAg5k7eM8POTalHfIwsxIrYF+IsZEjHBEAJCpnSLdEHBgz5is+kj3WI
NehqPQCq078iPoEWakxX+LC9x9BIhiX1Fg0hYCMWAZLBJiwAYRFwtMmacQO0
vAQTeXCDD6YoXqCb166F2c1ivjeGNNoe2vJcj5Bhh7r5L6jvdtdJc5pjZ1RI
ytuSEYMa8yfUvXpQH/JC7Hhx6vLaFlUhvKk/VlZZVioj25Dpycf6Lk/bnIZp
nDAbeO8CHeyNtMfeY8bof/D1sG7xXW3hpzkFyIrtTJo4k/Eya4OiZSAea3Lf
DHatMSAMztdDmHloerQAMi6CNRlPJfooIBdlc0BIwPHXKMtk5KdWATAZYrCk
0FoVzpdA7z3kp7dfrYXWUtU9V71UrS4BPCAielNqoS0bqcEWVfAFBFuZ686m
POgtm2OzIpCKo9NpGSF2eS3bfUBB6moDLKPO0yt5m/ox/tWR931ad7Rxc7sl
efaTw5wplE2e+dO9v6taqGTtjAEMLuguNjoRQlGu431u3I6o7t6RvnJcNz/D
h/oCerXVATqV1rv2i2xb8gcGdZ90V7EzzzXPR6cFL40IkfULxA7nvrckJCbD
9RhFUomZItZRUmm2/2Cta9u9dXbMOFLK+NCcwqG5V7OB5KMobY9UraoKVuNc
jJJIYhvLAUxsAVleke8+ZdySv4NLc8SL2tXatp9rzH5BfIlGPybgY2sAmerQ
4g9/ea9+FwV69jrx/+MogPY5dbJ8LTmgYh8LkaUOqCD9Znhah/8S+oFaBW0+
2NqPWSeVm2VMEUrdxiDtcjKjl1WjrFQj161eJ8DmFKDpFcIEVmprJ0/nhjB+
aoSK/rEEFyne7q0hTcM6S3LQN8+C1zCBPgK1fm5tbUzRHMyVoGDjIz09l/Ns
qz+F0S2ltp96Bd3+khuJPXOjoXaKIrx8Sw8ngFJ7e3LjHeFxk7eeenV6WLC+
n01pqboGvUpsrY+WIxshggcynZzUMxM82jRSV1Qs6s+QxYuHAn4hrXIZAXgR
FbblR2xEY55I4gtub6VLjgubyQX8nlf93fSTirmBqGfo41e0xKncBr6CPV8Y
U2s92E3xLAJSMNEghtlu9Bcf23HFPwQ8i+RsP+9/Ed4wwBfKW6zfMPSByBNx
f7gLlUQQ8WZwY/JAIZOy7H6kMy7aO/Y2FCzFeU/LcQ5SGlQSE47aoVPdzc9F
5pKmfcd9Gxpbk9rTWkzsjh5ooaU4Z0xmXtgF8Inaf+P3pLDx/89EOeh6up71
Pl+vwkkgX6t6XZO/U3ALDCz9CHQNtP4l2vuCo/sS0iWe04DXTyPcr7qpBHm2
iU/uwAdhW1fusJlSGRf+e4wYSUuDQRB79nH/AhYJoWhoN8gI2E/fbe7sSewd
5zPqkkTPGv+p3oZdcAUHa3otcIfvisCndUi8HAUS5/0RckJ/gpzJ9ANTyMXO
a11pHK8mbrRcBeDOS0VoRmVXluCDHNmYkGUt99fysyVl9ywdsdSTqW53NfRo
Rd3KXNaErZ/H9fk9peAJnE/+w5iUblvtMt/tayL/t0sw8270k/07kGs+bESU
XY/OyyaRgLJkBEZ0XeqQdvNadqwutl8X15cvwN5d8tbwk+YjGFKKWzLgK1un
C7oshFcyGlgjaa36p+y6GfOn6bHQKiRt92DKqMivHB/sWKcvUrvV7HoorKVF
XikUpxRUZJnH0W63lpTToYNAHvzH0UZId7bc/owvKU6u0rZvfLEWow4RnHGU
NUJaMbSVgSA68TTpdCcA/ABkgQOCLhSmSC+wSdZ1gI9I9NTcHNswWi4rEkZs
wtHmVvrsVpyzSwFkkZI4V4DHh0VuXxyuZrfOFRazmdlWXlEjFKCx+HxBHPN7
fZPvDRFwvrZVrSvrDD5rXF+N3A9PiADqt2wXP6+ds7Ok7ihuYa6DH/RBUw+X
RjmnOEBW7rOxDVBQS3pAqLD6nsjI2CWZdriBFUBxxHrdbDw0YJvDGEKAtmk7
D1cyLjP4Da9EZwzE5nPNWpNPDUFSQXCf32pXMdBklJRCmQ6VEq9hKYerV1wJ
0pw761ZqmlScVE0c2qvwgvWITICsqzbNXyg/aXraXJX+OyHUBVrjBtkrMb+8
p6j2t7A8WXBMIeYEUYyGjhGAm0VDWt+5tMlDGTGuzmGYbDCZNu0Tl0gD5MXl
KP8NJYSwfHERakboudKX/Vm2kGpEp/if+hPqI3xcId8Nwi/Rpg6iB5+Y+rfE
1YC8/euAmrRqI+j1P20aok3Y9SLBO9S0anmRa6ov0CHRnvTm+IaRR27t3r9B
fJia5XjHj2mkkssksfTvcLGF/iqW3vXRnaA5CdFrblq1vwACiuegLXAfqzep
I2etuEMPR/KHoGtxsoF2mGeY4S2usYI80PX/xgZzxnNlr8sjWajO8SVVJNBV
9anS5vvXkUFhMfw7eBJ1OJHEwq4x82iRDEvsOP16bYRt5/GkVodVYMjI4ID2
VbOFaCblmyNaMJlSw5CTIskCTxQWwRRb42XmqOiKWBgQlYgjjKc/Jx+EwpoZ
C/hku3cU7iurf2VluGBDqhVkR/0lr1KNTSHcfPfEhrtpZlPwLBH9yWLPnt7J
7ld1k0YJUpMqfd7EwAtpKZDY6xfCy0gYGs2hcnkQS0Ewm9eU9xEdOUCzHP8J
nZ1LLxn4G2A0veQehngIjBv4dUxJ3MYMD6sswhjavlaRKnsDinPQ/16ceg8+
nRKJIzFDt3gbckCxpht+wMhvFgbGKbbW0YoEhwRUXALqG6s3HAzLupt+JuJ2
qPz0i0mWEqLk4Xrwz+Z/fzIO32uHecNQlikTrQzOsk17gOA1JoMaiEYHtfoK
k+iK7/c6db7A8ZmJZe1z7XdB18LOnij2awRm7kguH1g17h83h4YaiKxznW9/
MEIMc2A/Ur5BHVRNeyJTLYKsnRuG5ibO5Y7Ct6opHcXkd/Ua7s7KFpOWLqhd
aJuV09xL1HDvBVy5A147fOg2+wXaHj/JaL1WC6vZsbjQ1tXCaHbFSErMkDve
kq3xMQEoGF50pnAvmZHs95tujKXP88Pv8elzTG2LAelAAaJYktVL4go6s6eE
7JdfqgcYZXDouIfEOQ8yjjvbyOUlR1RRKbClXN2Q8kGi3iPxz/UQqiwT0k5i
3DMCoMnHhAc3g0wsvUVzV/CY4DsM24shMdgo9cQsNZewr87DBQh8ARHpeaqZ
OK7T8IEV5iF+BBSPwobAGHeB4VTHH9vcUfMvOVeEFtSEJ3XWPiArmI5JJEQi
Xbby10M/aysIWQR2NQHvbjLPBem+5hi0+0t69UajP8C4jiza6GG7bToqWtkz
GAqwfX84OHXL29f4u9IA+raThjJUl20fhvCjNfDUHacuJpM1KeZdphFjRLoY
l9YyVR7D734a/Zw0nO1S/oh1bJeqpxhCE9znOkOnjUhB5tt1rZb4lFx1fG8E
jz8es25rbraRiL2nhctpRADCjVt353PsdYAp78Y7zNVeJq/AiqxHZF7htHNJ
ZYec3ZYC6jEHrPBsgKpn6w9V2ysRRFJscYSZmfZ+82GZuqmo6Z4lLIVYhj5S
3UKuWMN/B48inr1J1OCoZxbAbnWxfKFSGxcX3m2//6DNYpA02NgRlDNf2ZJV
Onf/bLKyMhmQIcvCUSYF/js+B7KqK9H2nIOqROKY2/SlkNzdXSqOMAYrF9Nq
h9Z0hk8/xcYhitqV40N2lRIbJo0vI4PqsN+kt5CZlag1GM29kGutX4Z8pa1f
DbiX8XxUO5oPDOiV+XTAXH/0cA0Xgmd9CUIZCO4go70EMZvN8nwqVYYec2gW
vYRRE6tL9038ak4ZYxljCfNyhkCJa6vIX8Fr2aEZjlIGEhF1nsdmQggcIon+
BwT+lzGPhIAGiyv0bmXf0l8E1Ag5JAlYiruUTGJ0evw2tHVSRfsNrFdRJF6B
KeKwWJUKEGDK/OfRaeCCTwApv+pJPgryy0vN1k6RPwtG5F87bUElNA/4cGYL
KpWH6ShtH9lzcSmVYZT6CD6PYbcjv//W0HATHT9opMPNskB2qK19WKbUNDY3
hoHvcjY4Up47LQm0yAyhDvHcz5Y8eOAlves7HrxFVxvivVQzjfMGvTvJDUpF
Zx08sgRJDQ5n48XHEW0/EiTvnPgmyUpg52jUfYp9NHzd9sspPPhBpcn8gDS7
/zHfFuCfr11Ss16RGhqnzExd0qXb9t/dMYHD1GcGlb0XzxdUhXjdcMDkVV46
X/d/sVvMK8ma8zqSd1HkNvg0FnB6KPFMxS64hSHF/DAwGmirA0dnJfP5zzwO
2kHGGUOichxob+l8wVwASTEMbthX2Vi/2RlIv6fnCAoM+72b04sXgZtcwbFw
PpwOTDs6kdp0/HUrRIqu1K/BRI7b5pvvp6T7hIB2zpiJqv0erkf8XjX9OBW5
hcSgqjAAuOFEJe/4BUx91exxmYtiGLK2h6VgnXVN4INElZbWWfJ1LX+qRDHl
9ouZEf6TP2Pjk4lf4kAvOVwDjeMJWcEWCQ5BeTfob5imKbO2ReZaLBEGw4Wu
mymMqaX1Fo6A55s/rxPbz5nONI2YuLa9SiOqIYI4uR+FbwIngvMKRGTGTjsY
IYVyzc3Rh/fjbXX6ohnf1N5fZyzHXbuAbSC5+bBbmCiBkJisUcL7M03eSUCQ
VIp1BWbJ80bxwnV7rKKH4BIZ7pmZfaRd+ntLiqFJTC/9tZn01qrBItvtewg9
uQaIOB7zpruXCjTWr80jfYrNrQJ/TATOdSfjWc/cNak/5oJ4pkColVew8xWn
zL9UoLcvrESv88bo5G6ewvkQUcM9H+Ib51p8OTL9pTBKRGn7+DzjHlZ/0Z7E
owsv8eAUWv7VbXtK4/m3An3FkB6eipaZGqilSPiBg8shokzNP4Kiep6DXlxe
61jQmhBqUtDKdQ4620qZ9HZauZrpFyUDKpQxv/adgwHSMlR5k94YH4oveaUU
PbI+c14/iChM5gkk5T7KNU+017WrUe+HcOnOoX40pN99k/RF2pDhllZNSpuN
KtA7vKAxM5TlajoYRlCi36BknsdKSLgpAJwtfgGNA7B8W7U6/CyhdnujAA/J
zJ+x2FPJuGlmix+FjmVM7jrQazd7iJZdgHRAAAHgSCXFOe2jQInjJ7W8i2e1
9LBrdcYr/dEKFDHE12KYd4MssHfuNV/8LVX4+Mqqi2/Vwu3GSWtK/GUeK3jS
ECCAkj6c/vI+OQ+3shPNKylTLil+Udo0i07YWaTc8U1+mHrgMANjgAwH9fYh
HL6CFBVmyixT0o9U2diYTWdjuC9krvuBJJYWZtngIrqBW0RlturO/GRR4D7N
heyHY02jptuY5PkSYzu5txVozPLx72glAapi/hVuZ2SWx8gXrzLmjH9Kg09W
zbpQWJXHQD7PKXjKtzgsWrTNrkbNeO9rghnV9TFkG2xr6nyHm33kZ55UYdNX
meDvRGFH9+hA9+kVjs0AOOt6hKHyvKC8mUitVVJ8m6MyMenuXRU00GT8ZHUc
1Ts0SJF6YDg9jcr0GEuAJnzRPzV/NGmYXbYj2EYNTkSvgpvqmj6S2WbR68xL
uP+dV5yNgZ0K333atygmBkshJSIyEtxqUkDKvYsx6DqM95BCwvML/yGm53pb
1diopu+susDqUXJG1PSmIp+YP52O4Tg/CTbVMNPdgjbWaEYcFiC7uF2qkFUy
TsxaOpDUzIH22MsDiCKhNryCxIk4Z77UjQRooUNyepQ07mepkG4MekRQb0LH
lqCsm2M13i9aSWRIbe0LNgk1qqA8sK0SOpOXjEWg1EZjli+F4ejmgyDnddgd
l4AItE0RxrIgCYKYmGoO+bJ+Xnt0m1EXGjsUk3bHl6J1EeR9zbD46Z+SKdwp
1IqgkqmrZLn5+LWWOYCmolXvA7oXq0pRxqmwIn84S4je6W9oJL4uo6WrLzZL
fwI9vXJNhlQ35AIWS2i8ca6xb3lek84DIIfxOMRCYbd9hVfgR8lNyyuGHEm3
IKkluXIJjwku5O8VsEvqeIlJseifCKRlg3S6xAeECYEzIpbHTeXSvxqWvTDG
TfeoHzpl4mdSDDm2K2McV44HBWsarIQ2OI0O8jXkS/jKi9DiwT9sd1GDAWcm
JINJwdBJc8sUaWzu5T3VZyjJ+9lAQc50P14nbhVF0ZkBs8VDZ1qqigyZPHFy
hUCTEHoav7IzQL4KM3yxaC//+V2zh1KYMl206/0IGGhfVo8DoLM2aRdEei6f
JwWY3MhUwl13ZNDuP6Q/wJAiVtt5AQ+NUkUZK1yeoR1oD6KLZxJxyFlDd30R
/sFM+8tBXDonuKII66UcFgy8+YJqkhu3hSEzDtx2HgPYlE/QmX4dg7UU3Lsc
fhaVaju7NvWbW+nMvcn/AdGi3vJ5aWTm7Ua1wrU5cOuflxs7IPoHTbXAyi77
NFDi/c9FskYKRjNKDwRGqUCVrsVC7OWuGkXQ98qox1M9fgbmjIBvhpHOeW72
W5P22evwJoT8EAjnF6ttGm8VKEryzSoCoNLyCbkMYVCAeJ6fIOjw2N/UEBRs
+1jK2w1yiAdwntM2ymj40VZ+JGwatBhqbTB2l1Yf9cGR15iR1y7LAhHPwD4A
yHs8SYoWB9JL23hJyapAVagFA3lYa9n5ujwhfgEIxiXxHfPtYiZtE0Rc1/HL
2Dah1DTYPt/lwy3gHtoUEI5l2t9JBzlxBm68W3o316AZkXBnwB02SFwBdmg4
yllhwNoOLTNpZBMZaxidmMqz19lc7RPVFJIVt3ydAF3nAzuFdOgqskwyMxvu
s/hzwppnIi4fYUWr3/0Z6fJ/svUnzUWo7tGW0mtuZN+FDAOLJvPCkgKZbO+b
2OdFv5ODBllKy/scPTvXdmmOJWAiBDAUDogMjxeNOcBgsW0k1fearS5XRRgE
IFwR9N88XgZY9LL/AYFIoE/fgK5G2ofgr5NU/5dyo+S/82jRoQcUSqKol8aF
gPZXWr7MZVeVAjiFwKABP4MjSzB8ETFLzJ8yjfgdQOV1IvxB/QeAoAwKayOq
5Bp56UZiJSpENz0YYny4oChF9UCf2C0Wx/zpp0DNiWr9Pj7YNCM6vQEn0Rzf
ii9NAA7LeWU1tFjwdGUB/SFP5DWWzf7WZugstQ/PXLZ69yfOUKvxxRuAFNzs
g20LqNSf7SBR0V3KoMSQXByJVrmVCF15V4tF10uugVh7PZpHlJbNg0vwlaLi
lMEZIYzM6UJ6GnWmzomWgL94Qf4w+4NJVEGpq4Wa+3Lzf3XOpFWhUNkm/Pzg
jd6faR+dzVoMl6xTreaCq3mDAeBla2cwW1b2Bl0b6otgE3Lf4RxpxqkG8z0E
ED8WZUaOwpyJAtLSE/9qYPOEOFLgYhjuuhSHhvNqtZmWKJ8plYG1YR3eH0LQ
bmhopMp2fy3zIR07opbIkERs7A6G1XWXS5YYc6x4+OiGELofKy0sW/9Yrb0y
mTVF3KPSp4wQWsGicjgaugkAZzt1XtFqpM+dDaL++PQZtzLAVIQ0tlIfuQlS
pdqgA9c9wJtqyE5l8+oEs2YG4S89kdL/m1rkH/GamWXPyM8uwPMYwq3YTUIV
IlyfMdxLT4vBDyzo1ZqofvuKmXs6wKCxgOxkZWBsJO4WZmN0B8n7umRMJXh4
rwzD717WGXWctI5fSiAaXjZdBeQ/6/ya7Txds3tIaevPj4u6CfWg8O5bT4oc
C5VbTZSBRjn81YofTAUD1if8Yn2jISqAlRnIY2WiypQTrLajZ7e3VIeNFlhZ
CpO5es88NKo46nk7P1pjAfaZArBZnYatUbV52Z4Ft1oeACGWeycZsHJs/37x
8Dda3Pl/yZAQQL0HPXDkTW+C+kKTCt8nccCPWYaEqqpS9ENEOXOvhqR8uas4
sazAeL45Z81pEfvgat10lZ03KYdNcQy9KWFnMwC0m6Jy0jRmxc8AcowpaxyM
1jnTuITvdWx9LR97Y2/OaBC14NCQL2dbXn/1DI39u6mWplVx7khKZlYbG2Og
/Zr9Hj56EdxcFi4rpPBAoKjVPY5WhzgOURgXB138at3whDYCbNTZd2BAGpQ4
ciG5Bi7d1hg+BcJkvx1sym8MB8rlmR6YnfZCLIUin4eoMzs+pHgSfcHo9Cpx
ExCyKlNea0iMK/k/wcSxFfCd6jmAIb0iL8iMRfgVFR7lIt2QeNNJVTOt39gR
k7Yna4R/BnL/Vom0ENvx9CQFdIGQX1sIGb+6v+54D8i9RVA+LWVXMi5/PeI8
LpUm3W0NWBVLoj+UINRcxgfBYdia9OVovxrpVAZ2dFzxwfeSzQHHRFCDTy26
kMdXIbDDkyQVgrObYhnS270FDJYst+fHM8EvRbBBnnBG62GeCr1haHeMbCGm
4a4NsLiFg2r2FLyhw6bs03aG63ZWLeOz1Ynp8X1JmzrA8ctucPE4oXsTYZzy
acoLeJETWT21PnsZarFPzHbC84P9x8Js/v7plBOfnW9h9aNJytAw8o0MXNzJ
ZxuiI0yDCx46+7eXzwW0tTaY1nNT9t51n4VXftvL8HNFQNBKtfTSrA/NRm1q
XhGCUbVTfcMRDAJxARLwdCHdnbxrGCE5jCVsEQPMO4PjCrdaMx+iEG4fCGwa
SisDfOF3zH2tAomlomWSkJDwVSheQLMfsssFTS0/yCC3Io+boLRELkq6AIwH
ma1ruOaqML3x1t7+jAdgTXDpQ13/zOZTOo5dPcNHLPm6qkJQ8+itSTESq2Bl
oujpG3nDLBW7KdcrIxHS7jxZ3pEGInXBnzP7wef1tCzNKPJgdh/uo4lA7kux
RUY/sb8TGW+OAVVctCm/zZWdqpJL55FPqasS4hmtXJPkH9K6pjYeVKSWqMNI
mkhk6Gi3rvcyyWY90NTc+lWvN0o5D88fBO5pz3qKX5J5M/s+ufxyJ0OF2jVQ
dMhMVYwMZMZCpBzEqnLUX/hbTtSSZfen8Wyxx8OjO0RywUBj4Dx24GbHeNjv
79l/31WuN6K6y42P/csbWvIJU+Pkmun00c4daZDPxs0Efyc/OxBCHQvCk7lj
DZF5/gmBdAiXbGXQ3cYVGHxzM8PD/W93B5aq/o71e7BjAs6fCHO0+iJ+FLGU
nkL0PKXw+4woE3kSp8BL5UvKUeVupxMrnEISNSucLdINmbQI+Nr24M7FHyzh
/lGIjzUBRcQMkbCXMXS+RkKGm7HGYMK5STfR/y1hpsD/H7c3gMeDl6968cHD
bPkAhUh0pWCtvBYo3+SiJG5Iot5X5NwyX/3xtWLiX+5O8sKEy3WAqcsWbN7u
qO3IeELhdssKuli7JeYOZALogq0ozLI2pJ/NBb6bZYuH0DpNsKcFEDrNLT/a
zZxSel+GuzXUqGm3lBX+KAfBgKcCcQ2Ojkq6cjOSCsYpzzKZwTXSfVfwkglJ
b1wwyHZWfTHYRBsit6DubizCQTmmBY6iuhDFubgUddsl7vjYNwgq2Pl64+H4
sH+57ptCMX9d8ZTEyNgWJt03EzSVRHyklS6dsM41O0eCRn62QBUUFEFfsjwj
YGq1fAic2UzhQHBZaqC4JMFJ4emGNAVZHKV+7zv2u/9zYY0654n4ykjqFooc
Gjha8nEYIP+Mzb79DtF36YuRoeI1n+vd/OTZdKcuHikhjr6jMre/zIjQZGKq
raCGQLbK6Nf2S7i54qh6Qp+quXHYGrjqz8E2XRUe2QqWnYLMuIhdrteW1C8n
PN44FFEdDTXu4fnjbYHG+9UnOTnyAfAWIz9u8tzzn2ie+p3uSrdPPmxzaKCB
ipcKOMArILH45YdURvRLZRD7C1xs8s/TPpyFoZuEtnK0QovGcZJ1qJhXYgQ3
RFtjiS1Vk8/HNeSAV7xS1B9d1lyDBdxlXjozEAVJXEwGNIZXKlqs2iMo4EN1
UdPiuAMi0BZFJV4+MjTEeJ4euby9XmTkHxn7Q1k7mwYksk6XUASolmQvuzkS
Cv4i2z6Iwo9mQQGmhg0ds2n2GC0lcnbLtLdGNjaojXKT/iWpZBHBJ7MbdCPC
rZYq7lxrWe+SUup1U3+pr+b9SbHHAbkqpplmtthA/PyVjk/D+M0/4d+PH/Q+
TLVVEJaIJGV/Q18bY6QBariRJYFwSbv3mnrNkC4wuvlVOHlypldxfxtVj1Mb
PnuxBKGPLbkWYjxFy3DiR3ihp/bHHKHdBum2VCE2aNtKXG8rzceeWnxiAJca
npns4hWntVaLUQAO+PDzs5ZkVAOUWBV/tiAnM0DvgDFhSRJsC9LqajR8qhZK
HA8M7PhvuIfA/1TwpLdu32Y8hZxsc8NBivzkfZQth1L2Z2zEjWTgyS4k1NfX
OKPiKEY0ZR4TXKn1fPUcjv8/W4FIL9aXxQeVP83ISvkRg1RCp08N9WlQGmKd
WH8HwFinHKZZloTKDJjXviOPKLVYKZAcrUeXoHjyDWri7oDYiVF5+KrZSZKD
03nHJjurJPhC2IAQ5lvX/HMhD/fRopxnXNzOj1YHHTxbhJ2kmYCgYIhEwz8h
Hu7UraJSEBLMbSvCMErDGJj3Y71k2q+Cw5RIhzeb42zO7hiaal9S1T3L0Pyp
q6da/tfGaFp4G/3Ak8HuB8nnO6+i/JXKxcsrr/Iz02uiyjegRgpaIvAjxkaV
tv2idGrLv5rI+C+lyiowRKeo1HRoID22Vl+Yyg1hIMGao3kZZuf/flWbC+Dq
lqEKqkv/6Z148r5hBT4TeH2ndJUJjUMgtXhfe9tJ1x5VPjMZnt4w9M2XGQtO
2+UE30pUV5AD5vohAtxmHa5CE71o9rHf+sn7S8ts9RGiKp9QS7FVCNFeaoUR
vYraNlKbDVWaGrlEe5ughOTTmaRQGOIbL9HKeelQ7Heh3n1AbT8L9tYYQPH7
z2K5r7LLz2foxydpUtuatSX79qxFTEH7wWeZM+a5g5z9tvXTLl+awlD37EtD
U+E+q9W7U29Zo8ZF9eoMmDs60mMj710OkaY7UdCw2M26czqfgZo+NCbsAFZ9
NyZ9W+JLOZGsNkkzYDXI114RJTrt7aaPFbQuaim2SQI7KYgHe1Drpoq5wi5D
i1fIpkyhBKYN8ht/gwvWBuEesLLmcBGTbkZM6Hu65Qb4ye3gzMztiulEcMCM
YGuBlFGF5+6CGdlwU9dNLAfuUAwsDna4Qm0d0qHQbhVF9ATnrOo8FrItAgbT
DTv6krHlfWIUwOts9wEf19kxzcVxIKr9VOUFFvU2CvJuFcE/iwpNTlF3mcIt
AxyIEYC90BZ9fV3TE6BCuMKNsamNGUvCEInmqhk0T4kmk78pfmTdKu45P2eD
yPc4BX7oehb2u1p4BKyOPoWY9Ht12t0i1D1YX8tvZo5EopevIGJLaBiLWO1L
xCQvPyglYv9parxqg7QWpiSp9kQfxoq38k6KuoIzOaUdaA6mKc2TYl/EXfGy
XRKqXE1oFcucMklaVgWTAHcOmejtef4c5Ch/ohsroHMgLRp0c5r9Rz5Lq9CN
zotJ8OprMJuOEkYB9A/9m0qdZ5JwIBprTxbBJ0A63Jicgq8LiVGUNt0DIvgO
ByuG1++tEBw/JoGs2mKtEqzMLvlfcDORY4jNN38fpfb0g/bQnDMptPmdB0AL
MIc6C2gsFuKq+KMOP1OE5SGzjLhFLBdruB9aeaS1Mr0Wau4bFHxuXyILjQPT
IGA4cPx6z5YfgZCr+tn/R258WssmjmtLXaF0pjiO4oLHNEd+NXLKgqDhZT74
j7rqobFCCXwVsmPNrG4U8+/IxEAQtsaSQ5wGTZEQcHGl8cir1dlJggDeOH+d
VJ9skOsbT42vllrdCfGpPytZZfkKxc3iQzi8e9xn2pJMq3vDNv8+cIKGYUpJ
U9rUe8UycNzd8Fk4TiiIYvEv0GO9Zr9kYIFMgCCTSzTeMDea8bbmbqnsMrAn
UFvpdjp0WlNYcbe9/7g6tO57aMms7/kCsiU1rQrqt8ah1uEopGuxNxM10Jfu
kDbHpZ2GkTzLT8k74TYGyMEPs9+FJnTFccFV9vEThrWwWR/4FtrxCs2YGPzI
dqwoVv0Pyh8IifNiKbD4/9gO52YclD1E3uC5rShK6V+QHPDmbQ6xjPSoBitu
8kJY7NQC69SEuzQPpvEYcKknnLYBn809Ut6OSO+HHN3I51fLZoVbkg7h3Gvm
g+0a7EFqLN0l7eIAWniv3382ad018i2tEU3+zmzx47vxuVE+V6eTXPBotBvS
ApfmrT8BtAcsAQPXpAPDv++WPtAyK4RV2hF9D5faiyOeaUofdr8TPhkFSge1
+AnNXLJZiQ3FgQVKpGnPphv3D8iuhHcmE+ackzW+EnPFdNXBtA5hM8cSJdaN
vbjP+lj+oGlZXJV3Rc2fkrtQv5PKQlMalmfbXWULHMMz5LuIY43X0p6Eqf9R
LRSdFks9ViXiy3uh57tOSEFAYSUYfuGLiRAOSaYW9Qpb/fjBlR70VnR1dKYH
KbVOCJiQuEvxJuyS9JaVrly6n8l6JvLMp6kBXSSj/v+yH9B5olSW2k1IE/Br
niv8BykJEMNydIJk7Omb6FLyTpSmJfXQcVjxNHNMH+6zFNFAU/raMbY5UV8A
hy/0HV6TC4S4SatayJwXvsOOouw98z5QTrp42BMhE0LQ8K6KKLv+aYvuFUDc
DPjessxW/lt1Dv+/hW6ovEa9kd8TL5CKPBaRVfIKam7m5/PhWiIRM0GejQjZ
+v/kxe3hwGUdwRMC20H6Ks0YqIpRwamH/PmvciMLScYrKWug9ZeoWSH3Sk0A
mmIiL8LdtQXy0r2pCCdXQz7/Dr1VCE00x/0xk1hH7bSzP/UAFXpNCNI/rrbV
YxXhZ7GDDlHPD4HofjRhTd9u1XSKNYweir3WZ8xy3RBJJNd36xsXCm00MXhG
egHFN1XadBog3WbczcXyo7kgHYWqGbBT0zyfNjn64Kg8qSSwcSjORCVI68+k
BIeJM0X2dUIWrjVkqwN8+yLj/vwbAmuZeIqoJWi6WPKmi3ty5RDsb5rflQTj
shNaG6QHlw0+XSP6ZG3OxnPOUQUYWHQXG0IbDY3sJkI3olMWrbEZetAYmrF4
JcEKvh5UhQKd/bXalW4865KaATmq7+br7lWe4IbIMS5HSzo8jOYzobmiW9nw
BrTGNr8Dvj1GXcdx65uZH5F7Vdky6xtQyAebomylpW8KpTFwvUurxsaY2zKj
tpyKBXFKmXFG/n/9/ifqphYmm0GVJNCmm3LkV0LAHJNH0S+RskVsmpU+lGYC
XOYKIe4ihnjOqP6nw0iRfhEPW8T7oeaA80+JRSCU7UEJEHIlBVXEBo06ahWC
tgtlThDHE7PV7a8zL7YeEao2o2QX8XbnxBX8wwxXANIRsZQDp8ZSxOI2fxEs
kS0zrFP7FjcaJbYMMUeF+yzwxAXWxt402v8H1MnvhTc53NqQ5k+3gkBeYc8T
ng+Go+Z1pRk5PhmbHBtUajmQHwloEdd9c76PZk0jHK2Za/mW3KYfMvJB/M+g
tQh3XSWybp/rvyKr41QEzw/btiKuhsdS2YvA6M5GkACqrLVz4YbhomBs8Wos
LNV2dcd0W8+jP+khOfBStk8F97QWS27AwgCb5YhGyXuIc1fjJfxJZMWPv8kh
IlNUJHwsGq2LzFega+HHXGnguvXwKIxCVYxyVNqy6x0GRY+tbOeqoReVLh51
8PybWf8qWca+EfKP1PllpNAWbAl1SLfLJGqqNGWOTK1kv+2b5XjGNCStFOkk
wIRg2W726up3fGDon8AXaWwKJ/ocbevMKGKLV+5FYqhvtGUZdTPfWwdnwbwO
/836o46X1GdTjgmBOrILyLZK5VlUtXvmGUrC4BzEXWpErwb6mpacKuyFmuiK
geSjTj3Stc8iCYjZDNsNdp8N6kLoUhtgu4xO+s042DSgQZ3pB9iMdgrM4D1T
trQgfeBQ9ifCHFin8Lxt/iCpXPUO7Om1uk9L6Mj6JRcR2iAmJjGzQ6AGs2AK
cMI2jviNcp9B4uvhL9c7lgS2BPuYdlWUJMHnLvsRBK3vv+N97F3Vo1ChtXVr
oGRSGxIvc2FA+MZSR0Ul1FlrK2MNhzFQoHAa4YUOhGZF7tu64IC3GfxHza14
FYqzjD1JFVC4n+hnwcTbzryZxV3chytaOYMhl0f8O1KDlOcmnbxp86xX4JIA
L+ODeFvCJwliE21x8misGQ53bji4d+pYQOBiCcCLAKlrr3/VbfxXTh4zUV87
Fd1MA8T60kYJiw3dK4V2uc3y+cvOMTzx7Ja66+Wm88mijhi7677BYBEBgxXU
2A/H6u8t/Q3ujq0I5xs8iiK1MlHSnTETco3t9z8g1Z84DCwbEzbZ5zxCWghZ
sQoUI98qkJo+f0KdriISiJLKnUmFVnshkMmmHZ+z/ObJ8tzKO6bUURj1X2GB
f8vhaWB3LUaPp+wqAXpxT9WZMPt8EeVBxwfsy51I6BPwbkeqlxh1qul5hoaO
8QWsUvM24vjBmyY2mT4e77X0Za0iSh7Mc+haTjF6K2TbGUeCDs+4H48tIKnz
P5qsIuI4rIrkhOwcOePpR+0XofCeikK+Dq4Pr20VWyaelvIa6sdWr8NHxfFT
UA6gHFBHaP+KwNI+MhyXV1Qlz/ES+5LL8zk9HZUWEZkx/kNEDkCBBP0prWaQ
nB7w+pTzJNSvU0TrqqDhNywJR+y+Ji+1+eJ6zK8ReLiLxvdpmWgLROYTiUBe
K2iCODuv3XhFDHXe0Zf5VY4RiFMptrT/dWhVQys8N9dYoWis1PWstTOX6f42
PyNFz5ZAOBDopeFHUKddfViMj/shOcm8wS2cHchZQuEGQqGvprEUR9N2WohN
l3NKNaufhe4CDVGtDTMVtY/5ZpySITHA7VrcqQiqWLhj1H4f4iZDMjYVK0MA
kxcFO2OYGixXVMlFw/7DnVfP2/aJW8l0gDc7MXm+x9ti6+ujqFNP9PzHNSF9
zq9THL84VbcKR+XQV9EbNVAuxu+ixcY8NuxyReE3uyw4Ti7e0Sb6dwtzTJci
TqcVbdRdPH+KMX5xN4ZqKzcLhnFxzywDVXkUeRG7NwxtNSfZaG9hpagzIJj6
TdLB6Lrn0V3cZzmAc5KcsL90GlcwAefHPns+ORkq23tZdJ8SzdDtB56WWzoa
a9tA7rvCIob4YtisgWdj0idXfMzXKf3ijGZpfLE+qEVX3aDgVwVCLB9HGHYz
eMxBWRPUbdPSVdHinAiseOlsuzbbGpVe+osWdytszsO4GvJTUd4qnclFuPm5
SYG5SdGQBlmBbSm5Jkra9F48BlmOGl7XiFV9L3X5+7FtNnLTCLjtFYapVS99
V6FI5hbwVmlp5NXkKRhJudpvr1NziX314CkKglO07VkkaJMSSr0bmmHCZlZ1
SPQrSvR8VXpAvVmFn/sLamjzRwz09heOOP2JYCvveZss633nqD4TsI8Esjp7
jLfQx/TIWOQsSyGpUTHR4CloSelopOk6iM6iQzie0rjcRe9AWldWQc9ayYxZ
+HEeetFk95PtCRQTw2ruScTlWZ5NP2V+DuRglZp3kWGP1mFRRcDvellXTHYQ
Oc3ngdGc/jG72FlfyuygZNaOqrxhuegRHwS9ea9SWRFDOhyA75c2XfUEX465
qM2ziAMRkcudifIU6pJjc1xIXsK11L8FFLK7KKn4f+vWkfZhkc6qUWsrNLB8
Hv3l0/2ZcRBGiSw49oToB4R4yOcjEHsxlz/7i9sjGRSzbIChmVbLoOk/kH8V
0EoGNuSDzn2l2pAql0eECAzB6hy4+AwvlQj7QKlORvvmG7tK/tvNKypS8vAQ
MjCyFsk4A2xjczfgVmLt9IUgVpqTPLpDFpRCUrxVWLpCe4Wxi2X0P9G0Tl98
okD6IMD5xkF56a62PHRiDs9x4AQlfrM3JIOaDeJQW78/0txtLbTOaDOElSoe
yJckQH1FDgsOQdrQZAZT6yxdLzJM3+lpWKjBeVmlJgK4bgM38krVFt8yrK+1
IDwTGyE+3nuZ64RPRc53eLgE5SxNv5qO7Y0k7Lm9j2PJLvZcleCbhuKgl0qk
CXHEy12lOYzNEOrsSd3NgK/KU9L5Sw4RoJE4p7xuDavw7PDTAzp3h74BtFeC
/93jXiNHwHLQeny7HI7aiyj7E3+OQRgVGNUuszjCw9cUcqOZmfmxN8N7MfGI
S4BNMou+N93NWeDPZF9yFfBtUTbqe+/aV9dIbmiG5W/a6MgVjlhbFmcRk1r6
vPHmxpxCsj/k53QVzHJi/D9iHw9m9az2cSUz3TZclrEl+ITy1KFf26b7ediw
mjLBbpbTYWalh0qo/8UM7BpnJYXGyhIWxQuvRNtQN8qk/t1I8Ozpa8K+3Aiz
3hoTMucobVr/hx0TRCK2w/E9LmuXfRXKkv9OKAIPbz6H/Dim6JWFOtp7duYJ
K/jO79FUGyCkMJ63gONvJBqj7vaHpJEvZO2pOytOKG+EI8oiCZXPgQsIkBE/
5XvS59gvGW/bZxo37D7NZ4wscSQC572AZW4Gu8o21FvRvnbux2j239qyqmWP
loRPSghwuE3Km7OCoiyUY8CEzBsr/G8QkbL3tUvQoIVuWYlzfCJ1e8pkh+nI
L6LK/YvFNDm0BIUdoMM02UbkLwstUfV+Ui/zGzul3BjuBXFbHp0eg0MUSba7
XtuDxDATIqyAA8ce8P8yebNPiiDUV+HmPp+5ke9AJQ/ixf7UX6D7ESDT7Iiq
1E5W5VRP9w7Q5EqksICu2xoS6Haiyu7lXUi9yWx/Rf0ay9qxJ2V8R91LIIPW
jLMSC4RGsb+2J+/+ga06h/Qg0FRhcvmyTUh6K0AqJ884fcpqLKLVrUJNUFya
B0p1DNEeErXKfQ3Gj/hHc4MqrWCrbvHuiiHiLF26XmYRo83iXCk47E8SxiwS
cJEfrKASmOjMboaB3crubaQi6RXZqsDCKV3kfLLn60wBcZf/tspkatXkSuOn
3VN2EfSbIx9mqg0cM7S2YSHk60HT/qA/KHpqosVu0nzCdybtmfqZd459J9aU
/2OWz6GYDydBn+WvQNWWwbL7Ce5EQXs7GtdOeriEMl0jnWQCWAxYHBOeDQ0n
UCMlDIRQTF2V5hBWw62Qrc1WSfZn7o+DABWdhmJXPFZFPb22kd4o3OQlrB3q
5Q2V64vKUV+AwSJh7NapL3ZBTZ7jtJwVkjQfMGszr0DeQM/U8KhW3FvzsUwI
5N+NZyd/GKpdJPDtCusKklAsl83BbJWpFb23S5NahWhKoGTwWBQsTmD1FJgI
n9b++4sPW8Lat099xZyFLsA6yzZxjN8JDPqQghhpCemUeWzx1ig65qxgELfW
YfMoh+Dg9yEZMXo1GpARriHjy9suaBQEo/s0IGppqdbbQELDHOm5CMXq8YbV
WErmRmnUg9slYYqrB+TklsBBWAJesd+HO4nDT8FRsTlgl70NSfjIGotmg4ze
kRQEcVo0nMaerzbvLk7FkmGiiASQc1HLNElUCVa19zebp7skD6TgW23RCU3l
uXGiA198tFLwvY4ZzZYORv8HNaruLpIKQKOLoC1oZCJ2+po0PY5J4LlcN78p
96oU8BBF3mxTWed+XXjZ3Vp6m1agYcxLA10UehFlu1aVcJueTB/0urtpUU1a
G5DtUijzKzefn5Cp0QjAXJdjz/rPIRPyhpk/Tq/yj84TVJFainmT6N8h9Kg5
TaIINkKnotsoJfHJ/4r/ix5uKuIWzEywNW+tpQOMfVdXVWn7/tihCDY2+ail
ItJMOi2vsHrv8ioAcDfE4qAoF9BnB8m6Ac+o1/ofuc/yU5TBmghsq/alIUq3
1cVzqIic7155Us8hAETfQq6MzILZs2Kvc67tSwD5gvlMARgkTOEn4axkuf3x
Jyv2HeXnj2RQbdH/MIX5i0f+QXmn+I/00U2XNQ3oAKNVh6Ss/xWuJ1z3XA0l
4f4anNpLLSlsbXLQcnw8CnkUvxNIiF7YzjfJApJBRI+JImlcbaUho3mkcUWH
PXZzFCRfYmB5t+x/R7ndmE5ISNarl+69wyJc8TJYN+Tn19MoaqXR3jWEpoiX
HmNHoGrljNmvCVllVNQoNW5eXMvESsG8JMPq5HydtoSV8opAivqGvSNYITRS
QxE5xdxzY2/YbpJJlvU4B2V801KVWhEZzuXKs34tVMX+3DNYSz0yGw1xWr9y
SQD6cBII/WPUUtdWi5FCBM6gd4BxLV6xBEkKxI0wAig+IMYW3YAbWeinAhMw
R1G/SMfuGBl8tnyXJPoBdjww4xdmd/SCpROfGZ1oQmdelYkixXv+qHnkZe80
r6nk3P49Yw+X7Eb8NuW3v1FIqIKCkr83AyKCLzModOZFiS5zBaZYOmHz+H5Z
lhrPUGOluyjZ9zDvZsANTFOg6je+rDGnPo+h6yJQWPvqxMRobdzgvq2MUFZo
JZNw8Wu/eDFchqyehUz59ELJyO7ZnEFxlnO6eSQYt18CK1VCXlK9qs/GJk7y
WjQLuDg4UGY3EpoD3ksCKcGTxAD9s6BdppTGGNbOBPtaA/JkxpkYru00acPR
Xcmj7s44OgQ2VRnm91LHVufM8Q3vlxM4hqpXWy0NTSHeQP2B0Hg67nnEBZpT
UfqHXvsfBZHi0l03Jd8+4W1XeRd/mcj6U8/rsuRkEMp6gQVcsi5fbdKJV05N
VsJcKiy6rD2vYi48/FA7dqhDzE0yFkf2AOp+XR/WjHTmo4bJsCuTmH1KLv6m
Sd8PmrRUeyER3jea4bsfDbq+6iNUg15tPq1CxY8mFR3xApSucXN48HGyafaZ
IrNnlF0paASRo1gWp5yOnwr7/wlfe6ItJDTVZ5NtemauVfrj4gqrf/4IPu5+
c1y3RmGgN73yhnwzj0Xxirf16LrBMSuudHV7zveKi8zTj/y1ExT7cdGjEbO8
qqFnvyFWwXIHKVGSHCfL9N+OQVAn6V5kN95mxfuTqGIFlZApQDMDMMFn97nR
bnjhsZefms0ig+8l7om6/UKAt6UXx0hUlw7h70O7QlFnuinXf6RaOtQzGZxe
81bLiQrS+ohT94jsymONx1++1HvtPlg7ftJXdR/+6gGpayWQeFxcEkJ4jhNq
UgK8atM49scAuwkm2SVzCnvw8IUtdx7uts5wBLgu9cwzmA8g0nkJV2IixIhJ
DHSQ14Rt8Q+9eOGd6cPzaSfEKuETEDFZCI9MgbRI1erq3UDJmEdxbvyjUclg
qVjws9YBa7dKROK2DBZLhe7U7u7S5qOIe1uFI5eTPY9i2HzGq+mXWdICNCS1
BBba6Smv7KSXN470kUlbUCBUpXS8v0Fi2ON2DK89aG53JgPhQwlERI/QwOZ/
nBKg8B+NxVsJaGXm1lNFAoUx8yUyjHMJwxweBuMcEkQoBUT+tW1FH6vFDSIO
wUyQc9FCv7PShaRh9xvPkc+QXQO33Vs7CpTFE90CzsKH/W4+L6F7KR8YGo+B
4juqML02HzCK/ihGuTNLBV8SVFnzA1vbXNC4pX1x/kwze9TDK8onxMERrNpi
qgFAwcWIzyHkdyrCOrEQTPQmsqAOmTZS6q1Tm9UcIxTA+WekDVDhdiCH+Ihu
yjg6f1UAVzq13r30diN/XgQrR4SuyKP2HBaPqUuMWRg8JBNZvZpT6IetRVOe
WQgvZAVkYW98LvAKm4Ejm94I9I1gI1kaSKgNLKkxrI4zMT9cdMwNStzIQdeo
ZMOzocpzAp4c1VSep95lUnOux+zzHUXp14XiRIYG/vRQ42phnTwBiosd9tF3
B03uzv7pGSnp06Rnb9sFRk1d0Bxr9Irzm5jYCJu3Mlx2VZKhfLW6KJsFH8Kl
QtlqPkkamyPTz8jyaOXwwEUXS5tlRzZZIVWsXVvPBHqvn5GMfOTK8i7kit9H
n7wexl8XrBWi6dRYgqwrYPpjZG62ZXPmn63/K7HQi3hKQDMZyW39QuS1jE8V
DJTCXTMVUepzJutn68jbxs9KL5n81fngQDQKYpSwfOETYY/PbjbDilan1VA1
BrgfGK9kwMwHe47gLE//f6Kx1hZlb0qdZdtspT2WkOPesG2IV2p3kG9k4f3O
0c2ZQNNyCfaMFA3AzwtAmXWwywa6L0mLroPRZo13mMI08CJRC0yMR3rB6sGO
lp8ZIoR6aQaHwB8Ex8kzpNr//3kK651tZxiDlk0/paXnsV47hvACPEqCslPI
lZgUWyFaOBmNfB+L65ivpym5P2ZCdyu7NWfLimv5SVZGwAhDEz1muX4qhTRU
Q3KxFvtTz1PLceu4Xp58Ofp+AwoxV7cysTvzi6RibLFeQm14tHx2u7KY37rK
hoANSVMoHtHWBCiGXK9LLBOLzOwScGWvGNPkNLZ1WueANIIejqzxa6FiBmp7
nFvCeXsEv/SlkgSb7ZuYKXYn6luP2pfsgXlAPS9/kdyBT8Nien51DevRJwcb
H8FWqInYihZ5Oe5a6c8+9FH6sAKrkXF69pU6tXlzpS5k5VaaBtEPXYg7Q4+d
T/LRsh3886wqTgaBDwuQm1nq2PwJ2mUi3hDKTQWvTLpl+i1f4ShvNfGDc6Mo
cn5cnUoSBNzaknzRiePjYaNTsezJ9b+7w1ohbKrZgv7WYru+b3qTCEGIqt9F
lfZzKVH4ubD+UkZq0cid50R6zZ37bLo1ce5C0T+PNxys4zb7RbB1DYBcYpXL
Po4+YQ4M7SO0TPzr59ZigVH5nU/g55EQiHsESxplARFjHHQjNncK6y+KfQMU
xDDa73DBzBUl8dAjO//Vj5kpw1sViH00tvSr+Qz4BJs6zHbHLhd8nwJ5bF8G
CCijziY75BNGRGCV9fBzuDupZlstUQ9bkTEwW7b0mmB/sSAErgOnRmAgYlqg
TszbBZc3b7xfQXbCHUs8/NICA3hpYDGAoFV4Su/hnVwa0LIbAkpWnAD5I1RZ
5XPi7uS8Ed/8/k/izkX+IzYes4s6gngjAglzcu7tK6g7xi/NVlswMmJ91TXR
2ApH3kZtjhfRJ6FEtzfRexR5kNEQxU6sRsiEZ8eP5/qVY5nu3htct1gNZI46
4p1tc4/9qzRI6JJNicOWNnh5n1YA3quaHPib8FmFGBPQyvVwSRuNm9mDEi+Q
Lkl0r1WIJ/V3NdAH4p6HccjnQAJjQMo6GwiltAqz7cRU6ZvOcrM/IxdErL6I
UVjpFLX14nY4AeTqeM/wcx5F/1pu+IjYsBTtOBW6iBcfHJwy8oZyKpxrSYdm
Y38meE/yvaOmcMF5X1A119QTTdlxqg1SXXw4ZHp03fAwWt9Tj+VMjqbjJAZU
HGiL3jBk5iqOXcFXWGXFsSMdo+bU/OiWEhgL7p/UQoZtAvzplphIqg8xv039
7Fada+BMtXMjMDuCMiizcrr4Xfsy2CFG5LS395joAh2xMbw1Y/sqLunvvIPg
9shnKxeRcFf1Jn7pGT0IRHIcb1nRdxVLbg0mtolDjgRmgP92RO5yDIE0zt04
4wBf7o0CVnMPJ5ApesnWXVH9T6Pk0eQ69jGhRD+PsrMLVA7MN8v27wAfu4UP
MStL3TL4U2174Q6fMsGK5njrDznXj372LaTOSxYiS8eKmm6NwekHYYbqYtOp
yz1ANX/Z9T2QQAjLrxyA2XjorYQy0CDHlLdPQge7f8F04/BohBVgzr6fUFOE
t9rMDFscSqO60AS/xBRpV7OU4zj4djCbXVixFL7phtpV6tVInFkHM6DOQeVq
I+6rkHdVFPgJNzWpqqlMZRFVuGp3a13T5KXf5BX3Y2AsXIwfvB1PJNrj8rQO
bg0aylnl1qkHz/BuWvH8kdbC5+ZsxQ0qKO6cA1CHvNR3WVrmT8OyjXAd2Mvu
Iyb4bGaxB36WGFcCZjNHOgV1qCszdWVJKr37S9jcptn0ZiG4LMkr3OmU9HVK
izSWucSBEu12xmfOOnzaTzclzKzHdQtGlC+IIaDrsWPS2q/ctg0A+YAMUCMy
3AIonvnm6/pkkcFWm3T+fhvYSe+/plaCMXRKy5uIw4gLmQ+g78twb1kzeyaX
56wlzwNyyEHBEU12IAl3c5oSlFwRohRUPpe6m/3pjlKtrLdz33r1sIbLhs38
9P3jnKuLbtHPkMDo0y9axB7JgK91LseUSj8AMpyJ4MojEzKYqlisnCUqyKNH
04+U8VSgVVrb8mPCxqcWtuBF1PXDeq60Hd9YkFSXsx/06r6aOM2pQX+5lyto
hhoslHVzsEOkjZNWA+dO5btE0RiUO/ApLctOjdmDpQyLGXvvF5zRy5eVo+7U
r2SJ3KA01/sw5Chk1Lf98nRNL/dn8NXKJepRhO5xZ2evNGtj6y5u/+399pwp
v1ZSg4CwoDmGfGyNBsJo7IJInzgrvdMIWv45Skg7lvYa5FO7eX6nt/n4DLrp
feDS1O/ht/MKF6i+exKx0H4pm5aABU3qsQ8VOVn/V3XTQNTJrTClBv+eDJ80
v+Kk6MmwiXdtDTC2T6g7H2vqRbbUIxyMKL38bJ+w6fYPtDRARts8Be0398u9
waZ8gLHTXNl4XhvG4hIqT2RLqemln2cU496vYontE6zvq2UvFm73XG0d9Yu4
xlzR7tnz5G0nlGHBh1uVv/s5CAu4Y32qOuTId/otV+VNOEXpjmI5CdRRgBb3
gMzMhFSNDCaymimiVyTfUD+vU45mIWv0UeNh7udnhUQBO8OamzPTQFRqOD56
GJMHQ4qwa23XhQpQ2CnTyqqGSAZvnoDfcRl7lwcV0aI6Tznc0dulfeIFnU5R
nUuiBAfS4PYt3/TZvLi2+rA/qyjqK5lu26Xi4ksg5SRgHbT5K+byXzZVG1qK
cUd7vyLuFkpOso9g9E6cCPzH6SsSwxSApg6NeFGxiuX7/TJfglC6HwtRRiH6
Re1fs+5LgaHodNGM1iikJ7s8ks+V4v8hOeRv3T+SBMpBbXvBmXqJe7NVuwHi
/kLjXeiTe/8CDbUM2SxTZulNxhR1NGlDfcXoRmEu6j7jf2d7XYQvOR+/N7eg
OFgXoyiDIfzaACzRmVQsSj7+2E/zsX9B8DjtxAHaR9lenqbGrSal+UlmO+6q
0dckaHHNqalBZ9JdDUacDHXcN4n+8pdKLwE85/3BThDb62GJCVFitt1Ri9vX
i7DiFi9JSU8A9gJYkVIWbwTMvGLWNaD+zvnR/tcCwKEZpUJa1/SOIR5NrEoQ
aHXAjvbBrfkvG8XMNr+/qyOocgBMdhye7RtqZ9/HaVyDLzidFiOsj58bSYVC
TrmRtjkwmTrUzAzuZNxjiZ5DQKHQeog2WGE4L4OwlO/2hiFaCmOaLYCAP4Cr
gNuIRMaU0OZfwjD79tgbp10UCDutzKJVhiIoSnBVfTjnkl67sVjOgNKQBRbC
yREqp0Gdp2X7OdWDdLT1Pdntgd2hNoHV4iIfXIgMI6y4Pw6wFQVkS3kwwFCl
ek70hpw88BjwIPc5/vxmHZaVZWmYZs9RbyXC3CuQx+sj6w+KPC7kQWC4WSk0
wgrcXgkdukNAwMl3i5oahaE4NLNr9B3HEf3O+sd6cP4VV+AsoOr6kGigbhTs
JV34DM5OYDsPBeakoD2qJVaDsIdCL9PeUyvQugPVLaKJCtrZXe5keWpLIhFE
pMJVHEXXSE1Fi7l3dv0BOk+uSb7MX2rBqD4aTkdtvNCR5kk5gmMGYX0CWRFg
ATn4R0+V2JVeFvNe8zJOqtlMOptg4yEdi3ZubGqgX8XG9NtjF9KzP28NLTwg
VCoGnpqk/B0TtOrFX8QUDma3x9Ge/QgMQYvOcQpvluW4n9hKH1iOH9uIgPjh
f2B6lesa+seCLo5iBjKCmriJ4wfzUS4orDDbbbxtsBd1b6WZMviTbcYWMPxb
wIyphYLjUqQpiWQ/iMNLCh7et1ROeq6INhakGvSuqe9OKbUMTbCKA5ewsScu
9RmV4DbdIi02cTHB/YFNmdBzs1Opd4u42vWj89fhn/trivXFtOEFY+UV1e9I
lcmhdm8ZFhdGwnR+lKYlk+A/mRj36E56ri7R8jcBm9RFxbH7is/EyHEqZcq1
A97d5jQFZUOp39AvplL9xQjPpb5MUfoez+zjxVtev0MwgWVlA6LAbAKFVaV3
H158CicH8hzp+gWy9UtSIDf6UCR/D4/RXPcDWMcOKiTlMjK6Zwf/t8QmmJ/v
yWiN7XF7VM9qOwZA0eDTcAs/Xpu3PD5yAaeTUr8iECDYUIsgPLozMV//e7qH
3j817gwZHn13FQFdhVc+7gTRwVdMPmFCu2uCTyKkLsCLVT3LZ5NRYRQpIPwg
HYvdflfIfOPxQfKBBL7wp1mxCGAFC9Y3ccQ5J3wiB9uAdkxg+cqfX1gqUC81
Tt1XMLTJdnl6v2TY/1hHrl3F9+OirHSx6tJQg/rpFIxtnW2UzC2klN6O89XP
xRxztDJcSOBsUMIpLn0Wcwtc0KBcZqVmRrNSyoNEdrneISIUqjqLV8A4A+wT
9C7B9H6XpQbVvJoR6GhjHvQIONkZkYBj1woclupjnUsSvn3ZupimdTpxIMbt
qxniuLncvYLkVR/tPuuKlviOY6VnbIm5sGsk5cvsPDwXbNbKTz2rzmL8uDiM
SvWEb8NWIyTB/M8FykrEIB9xD8U1GQ+7449jJw1KuY3UaVW2IVOozQ/RNXsu
JnntwjaK12a45zOJQWZUld0vgGtie1jMkgSBCEWBQNDvMgYLHDGxEU1+YOtE
NSQBsqBYMJIjLKJLCN6iQSum5Ik+0i04Mof/K0Brl6YsMwrW76+oMrDZTe66
3ljnn5sove4jaFlsFtnkDhEguVX8CWLCxMS/iey7oG2v2o7JQwBWwuB/NN+R
k6ZgbCm+LRzaYSBHyEMalRBDvuFLylVjRqBRyLUphm/RPyioTi93NwUwUUE3
c0ZObIuugFAhXj3Kr21XG/W4+VpLlWEFko+xKPzH/lQmLZU6P9EMKeFRSpGb
FuaZIy8s4Y/YbM+E17CQ5zNH5Ent/Ql0mttoKGH8rdOMpELjfECDRyuN6sOR
8yWbJekA2zgFgNxv1w7VwxFEkjnFnQ7qMZ5SolPLQzCBLnlrVbERYM+RmZ5t
y3ZI+DNUYVBkSB94EIp9ycXaCiCNpRpKGYuurgn0MJueVBHPL3rwNEgv8ou+
WoKM3pSDAjGHd5b1DRD8rQc08U3tbdbBIFwGfejLPFtIl9+7F6IYPdFaDFBE
rZ3UyNGLAE4RrolUFGHog2SBOIZ09G92oCQAxMS1VWtQrIkjngqNHZvFTqVZ
InucwGMxv5vtpmTcEZmdXGaNFAoYaFxo/wp0QXLsEcHdcZEt1XgUUbrhX+l/
LVppRwwsMTb1yBzISZIa3LQjZkQLkYUHkOupkzpdHHuhqKg+1OytIgRSt9+3
d8qyWrRpCiCNz2SbQ4fQKezH6I9WX0De7EOyN0S7f3DwSCz/daCyotCEwMAi
Vn6uYLAY9dM2oH5dQy8LKDjw6zLs3wTk14i4ulEuJ8ASPqw8CRMpTaQCCWIH
w6OWQcq98X0Zi4RaTkFRZzxvPniCtIrogBZ07iVVOO487TEwNUM6YYdOlmk/
Tg2kuMu9zccGK9XilWif1mQXiLHG5eV3jCfJkoBYu+IyvGcoOMEYhFxtwfsZ
gmcbsRh1qqtSzuX+0v5h/qaF5ZTkxZAs9+in/ipO3mzMqaGNDRBsVOfHIS6H
wZoHn+fw463F3YqazHSSK6F4vNsXJEw4KljmrsG4k5NZWi4P2ZO7CaK0Mame
EpGXz75Aee54SzkFQjNwX5twwVtcaFE/n0sfwo1eRPQYCMHqv4YVTnJKoD0x
jcjAkzZXwHbU3ycbQ2/ck7oUfimvrwmAOJwlgOoIXRwvUbCo62p2iHtqBgDZ
GcnhglO0wM+ccnCBxUM5LaBt/UOLJ/dgyz+k3uhFhNN6GzdAbMtfGt/u+rn7
IscuQAsRTTo4H3ehzd98V1GXZ6yTXQWRv9RKEx/6p7BSdj6VNa2fpRuGmqLj
VWVwif1t5I0l8IXFb1HH/HQToBW5RF+YMiS0pXBtuvaRHvjez7dZG/SCle7z
fUOVjSmB10YWLwxUeuPSKKwMkAaWs93H9S4fFfP9eVJ+m1MMrwKZOLDminWM
R9Pn0i2IO+xa7roTX4WFxIR7BB9IrfqrFEU2TusHnAZSY8inNywj3OzxMUL1
W24DTKsj9mgzecixm5c0kOjy/pJ5rqZphmPvu1rnYdc8tM723lTNFdhWuh1O
xmhyrBo1PUTa2ND9a8TKLvPfXFJ9dU4IMnxOL8njsh81qpofoc7isMpmHeI2
H0OKwr3U4XEjTY2w+6WceCBwoGkVixA1ub1NGYHOZ3zLHFdGUoYfwqFTpca9
rlbOlnytu6nnVW4OrjFJk1G73tz71LhgaVbnFJxItrcAsjE+vAbd0O9VeMCh
4isYRPcfJ9J7eumpLpSQlpeIqQMc5Rx0452gO01Pj4CLyo0pztzZHxT2TC3W
Da2fTxFcJOnzIJcnvTCbv5PHJaWRt5l/WHr4GWpMZR8vyGClIvVKzEh7iVNa
Ar5s1Em3hLyXjFluCbvp2rRj0Vxwwkeww2ysFrIHd0YU5oEE1Cc5j4jNaTNu
bq9yZE0pnygdhrS1HxX3xpi/WTbERQObdUMhieDysC5z5u5SBY75Ll53npH9
dJOYC2zE5F8h527LAQ2c+rgyzL95l/vPwONBf5T3j35Mnjf/ttKBycEIxx2m
xt3FqkcV/y918LuJ9N+mQnuRxPgtVeb1mTa8i0aA8HcfYtRP4I8Ac99a4mnf
emgV45jY7Uvdw5CnjMeD2ob2DyiEb3JHkVTWsc39A4Yq6qrB8bxRfP0W5LTe
bctVBOd4qRnM6xBYyRhLmz2FByuD0T7vcjBwLLLvpy9eCEI9I2lXPVxNmXGh
f78Y4P2744TJmI296J3tFouDLkwRcg0jPpvzPgXwUqjV7ed0Cg59+a/ZhUFA
swt/CriYdmy0V07xAcZAaTbjafsfS1RSkNFpNUecLCoyEy1hyTfJbzjn3wOX
T00hmqmYz3m5cEc/PJBmedwhbCICE6cjsrdFfrxISuep1YITCA3wkU8dj3Tg
3fM+uMH8vN10FscGN/1PL0p//a2Eqzu0OK9+Y3sw56raI9g+7zz5lgiB/lkq
2aNmvSgBfCZtMx40C4Ud0GLj7B5CdN7UYntGilX2loAUKO9HIg9ILQFDQEur
LpdIC/zo0jPvWFtrbyflhkI9lKaB0XLWRf36LkbuHJNd1+EfdeiHXcFj7YyP
Gg9ee99zCW3obhoBpyq+GulFqW8shyVGKqcy+KsF0Me/o081eIuV14m9tro6
AkShBdWA22s7z/1hKHwASGJX+9u3SXLsRxXQQv5RQk9y8Bdtc9ScTIDOXXz7
J3lcgFMle6b0wI2rpR3EAZT/D/cyDYV7hAOqhV9egEd2lqTSqftHZeZlELBc
sA8jW5JkHui6gCzQm33e5zn8vC4e0tE0ppP6SR9qXTn6HzCZ9Uh1IP5bW6hi
Y6GI4W4aG8B3ZMqpclsWHD509p9x1qnNZ58CZFIl/0cWyCRZIGquk0C5sz1c
y+d6ZHX2O+haa13nt0G2aMV4PyUOsEKtwV/sBKLqQqSaWdKTuVUTqwAWKAft
TM160352o7tB51sm1lv1cfAOicEuzG98dWM6gaEqDFelJ/2Q5E8zSQgjO5vu
ftgRviWxWkOQS13LgVn7VSqBtlUpQhLLaxcpEuulLNEOwtgo6djVQR6cA8W+
ETkxZ7rrAiiw2GganO2zrqBENn/KdjhR3TW1t0NQsCUzKgTnemayhbDuopVL
pgMSSuq+hGXugdw0PY3DCmHb72jdVCdOK9OlT+OxhdfQI+LDqwkILfpZ+sC4
f5MnU0JOvD4LSYvHasJfY4cEN03PBGnXpZGXLPr6pZwwDqgr+7Toiq6rBH/O
jqmVlx1rjuulAu8LpUn4L9GcpCSYA99AJlXM+l8qstQokAN5Ow+9xKAeQFNX
7lMH/A3dZZoOwsAHdfcICfOK1J/Ym6G4hyMAwDfRDNrEEjcAS9RL4jzLWNFh
Ho5n9v0vT4s3T0hKvUw7QsVErEYpva59WyZjzE/L4Q7BfVWAw0vRqjuuibyz
s59ipuzgFyYUGvOkC/oT3qkrTPZbsYllS3edOomG9GIlIxfv+/TFcAxMrt6Y
yErqgcd+mmfCpSIBlCcOAgRDVK2+e4K4lFMmIGeDoepnrYxe1rZYZ9fXD93T
njX4mWebkDTmKbfG44/Ykfpbh+JwqgZkmy/V9kV9ifVBbv6rixG8QkRKuuB9
OWQ6T5Gsn6alrZe3IIQhLB97YYRSJ086rjfhlhGjUTVKtgryfn3JjKRPSjlv
d88V6/3vrSfmnoOlqjNhrOzWNX+/7De5pfYsTzLfOfYcR64RNW/K0kVlJs0s
OVPcMdzAgGow6C2pQE8vvLSqY5NQKtvslB2oADA4gGDZ5yFYIZ3/kPJENLe7
QZzfSM6bghgfFubfeYO3lNZKxijZMigqae2ozfH5BbcyHt/2+XmIrK1/nyyi
D9wv9z7MpekhFgE+iFaPfES8oRsIvXt6vnHN9UTYzHhMRm2ikIb4FEZJO+n6
FOnxaP9jTm7Gh/7z4m/RXyew45djJjsSYDSbFJ+fmuw/1+EcROuUxBVigzGH
PxfC9FSGpx1oKatCuH/6gmsQK3jVZWygAqHsLCtqksBjY6BwSdx8E77DkY2n
hCn+pLPKEYQR8uFxod86gUFqnwqGYmwA1Jsb3YTz8wOCg9uXlWrMRMiglbDb
3tbMBH7yh/3SU9k1gKKQvYxztzyHYPUsuxdEMyl8Pjs7p8rrQGByEniXPWo8
B4MMkvmckaxorL1sWE6b6AR2h4prP3d0+rxiwNxlhWGlEk4m1M3taV5d9RXj
y4eCZ6dwubkkMDqnZIQ0TdnIdVDK1993wYB9OsxKFumwob3um/8gnAGfmjUf
8ZqaSpnzZLiFgI2aSC1gJhme75ZOZAOYUXfu/cpe1bR8xkU4uhKvjCwZDmQ/
PNSPyg23HJ/FQLWBHo3KpbPieSbSHzxYfEhW9Sh4TB7wq1XlNoONlScT0U4f
IzeGjmbMtrh0/pFEq8V9CPXmFRZnTkRGZDcQdlekRvSE9r8Ajnsw5Zcd7zBl
Jahl3bZmYuu2x4kURqHgx3RpCGxk+qZkZljD/25z9ay/RTdC+71q7KJRGnnX
yAqjBDGLueT8oeE7GzPfLwa2ZbR0XYSZJqGVg4BQA1NapEHdcAfLQR6J/tIv
LAaWzr+afVuywXTLhhhfZtGKZ3FDSS5yhxXmPaeuVK6+WPOzLgqUDaxgp0+Q
r92Sdf3eQOJXL2R5CW6iv6Z7TPMmf7yTWN7EpzA2Tsg7aQjPCAwXyE+7HFfK
/PeIevUvkWwEX3Cb5SpIjBvZZhAdBxCGO/rmwwVape4A8/+tZg/PFTPSC4c+
drTmN2JIVTFz7nW2BT3xusNhALfoQTQwj+6PhjCNBfU193vtaEnqvCr5sBic
UmG2UHzRYoe+l0OiTVRvWXZtxff93RaKlhDUPvBp9ufC41v+HzPBW8JUBzja
DNUkc00pfsKpuPTYNHrEzDh/29JoC3c2pq/6LWxYh5jgYQ4cISr4MUkoCGzy
r1S4rSFr4S08AN0cUmgwh9f9319fAO3q+3OPYCJBeyvexlf9aQ2opIB7jF2Q
nTGfPQOd2k7+nsWNVK0jMsGPcA11kG3FWRMVvTM3cNiErQtwfIeUMsOgLtb8
d07w2QOVOmh/cchPww8SDJ60IWCfznpJoVGlGHbym7BQF5LEP8JALKts6Kg1
EcnfRT2NeyW4kazizHUwvqsuSxzqzhASbJagDlmaNCG2t385q2Xnh4voz3by
3jwPRf9V38PQV1u9C5YzQnM9TB16OBpIJX5EIVkaiZ79Tr9S2K40bSfAuxKv
p7yl8k79zTx8kvs2FXR1+Zuq1csO7XdMHr2vCrWke6iOQvCkzELT3V6YTL17
qM1Nd2tRujMECT/glQui3Fd0KgaT/WciriFsJWJOKFh6L8yvzHWF2QeEW5XZ
nieL2BqP/n/Wn0GclqJbnrDt2O/Fx02BTW7cd130oEnvWLstr7tFrtSUOM5i
rEJSqQemuC7yKmWY/BAHk5uxgmXsW7S2Hm+4Ch2O12RDUriyVi24esaFm3eu
eZenhCKsj8A0QSARUzzqa+QTTD2teeKWzafB2SfLKHr3pA6z/nxQ65ilN0Eo
hI2MLldPcK3Udd5znJOc2dWzh2KsFtGgVvNHutoZMq8bZxOydebwbBayOZ45
BlRXHo26QLoE1bDVRikBH1lQXgNt5JfvOlfCdo3OhLxSYktSglSrqCcHIIoD
VU6rAgQFarLD6g3oCAx82OGFyKjHVkJ44KENcWHJWKlF+AuGldMYLySDvt9O
kzZtt/2HuKn0XbJJGicWYpLuZww5IDdS96XcPWEOlaO+JSDSLoK2bieV8wKI
LXWM5kMH4ESo9++r3XRr+Rr95/jm2N5+ggJXRdHH5KeVzLQAu9ggTIQ1wj7x
tou/zq28PCE3K2uc29wTK9wZYJtcJyKu2ZrdEYegdrpO0pWPWfqMuZvKjeUb
x0agAM1NTOvGByuHiYuC7J0x7cjtwggJX0H24xv8val/a1gvknztrFvAvlc+
RKV29yRDppfoSLm/PX6HY6mfr9gd43MtedBpbS5fLlLyGXLgEH0EOfj+i7+X
M6/ZupWqf9uCp3p7wLjmsYv39lsbdnmyJCoj1sOKpZ4EesOhQ1egYpLnb2Y4
DvuGyJZq+0kZCX+kQoFdve+XN28TwmZVVpiCTSueYzpC0wKtx7zJM+YauPY6
emjHn3IynGLvlbY8ZFefnD6C3xN0dpkulSrivfCotmwC2w/9LEgNDOnEhrhh
ChpGk/cjZ91n5FTkxhUSStl63Wft1YXuKvRMsDlUCBTkk4EWG/vyjsUIKWA1
1ey8jJeZJ/GVpBnRcDvFGWbz3FHU/bsdu1ARneJiLRdWuq4GZeRd5KsAQB5q
ZawBWRYoWZt5+DLPV1Tp2rMG19LxphwWh5dJhqOIZ1v5mAN6mHxyKEL34u0f
A4jF9qnOsksofZpLJ8f6Rwa7VSgEnRZZAjOJWMcUbM3nN7QmEETs/SVEoj0+
bRfALMRHcnOP15xZUjdBfljRK8wbFIM4aOdDsA8UrNg0YBGhINh16jSXIFUI
L0NsCh4DH+QqVItC2OtbZIp3ub650NsL5io8KXDjt+a/TZ1st8cxPUXb3hMu
VHXbbqxYbimK12LukkIWkSAnqzOtkkyf6AhWFpWPlilnX7d9uHiAKmAeNMU1
x0fL3zwS6BETXsjGDkR89u1jwZAyV4OBiUmubQUW+jsHbZGwSC2aP3nARzVk
tu1EUj6q1vWfAu/zMPwoTSRlJaiBbSyGUgXsptJldj5hz02zvepj6KAFCAMe
CratDmIIFhRhcG6/0bUYYzf54yBvek6rwvhH91vdFdFvMuDlUHOkXOeJeE31
EjJ9Ne/ppUqh7mKxCz9UYGZM6p3iYZF6c4Z/COEnpsmAuqJShDPlXt2lCeF/
PhTKQ0qGzvJ7xuq4X8NW7ZNR5V/J0/RUUyI6y557+Ga/dShBfVKtzYuQrYlw
a7EeN4Rr5jNZRY75seF/XbVDFKbWY4FwvN/2kXzIGnMacM3JYlM85Hp2YUsN
xW5U+kPj4SD9/yIAOipn0JXJbdm3Qkoam25mIXpTa0zd+cUzmnZ/q5ShP7qN
hRruBy+prXmENbeTnXKobsz9YXB7KYXsAqNdhRvEAdroiWqSE4BDYpahKWPJ
hBLL4GR6yqEiRvHTfAZRShOdaL3/2Ej4SgHwXJYYnlImVM8FKPN2+BQd3zjv
o2tvpHSu7OrU9A/ZJfaLDv+anh2oToTAR5NteNhy68Y0w2c0TkJFIz+Opd5i
Hxw6iThNXdLSefEnY8mQbxJkyPgs0kDI/03v9qQUgsjn7s0OosYjOWEiYLLC
mhKQTix6jbmfnwvIu2EpGaUrNZRRZBOPUIqNhyT1bjt25FKgW3ogbeeVlpqz
IyZUXoQA9UH1WfqOP0K7SfS3mEoiQ1MqcFsQaY7MNGoi0hIwtlWJ41GiJwFP
86I+3wKR0/zzuZFP1QE20ldeZIQuF3HsLr76H6GhpUw5ev+68jjtdc8EkElg
lEvxID/JQMCWoLbSzo4V4PApbbZAZuR98N8P/U+tTGQZYHXfrfXXSwj3lYRX
Qq40mOVg+zpceQ4SzUh8uOcXdCJQJN71pVRetVeYi6tuWWaFidqlIrV8lZTt
AEHfnVnlBLS9IQe2bvGk4PS+Kj9d54AaAQoGJc0T4LhxxGRHpqZWmTwmZ4E7
nrn1V4NBZGuelErPO6JVyzIWBlqxnTvX60S04byQ0TivmW+E4A1QUU9Pyf3G
XuIkevrgQl7RLve2RsS5EDTN7PaftV7fh/8BqlsLtXdfySLlmSFVKEFwMSSg
t2RqPhTDJ+puozsm2w5ml3doZ53izL+1iZa7S/wh3ugbwbUxJjM8VXQZS2Ot
Hfxw+TZZvkCLAijAi4x5il15Rqd0WxGi801swVzL1OzyK4jcjtIqhHnkKVjm
4bJZz+mMAuhvfq13PfLDZOVTPRZqDNU80pF3hjSxMwjugAlr3ozdARRdFSpB
RAWBgrszWziqw1xAkLrgezLKhm0+FWxKai35MVoxvUYBEKQdQj7is0n9geVn
qcsBmwxEWbiLlF00nvrSiZ9tJHROzRfNLuucGedOAV9rZMneZJLB+bHGQXiG
eb83ZTPzi4s6ISYpL/oExa+HvUaPSPx4tcTDbZjksV8jHK7sGa4Vg86rkWIg
Z2t3Saa7quJTmGNOJ7FuJKsiD6GOXMD+JvuYC+s/8hAJlw3tX2CKffojKVIl
oPbe65YCQ5+C4ly3kkdhHjqrZLFjbRpbz2z2Q6mKRGtPXKpIz2zYcVh7OlUx
p5nojsapR7/HHlvvb+hp9ocmSIx1bHtS7iveNwDai0y/nmKolLNGxjRTLufL
byD9T66kJ41hlvbHeLuYQl7epospivIhRkeI0V+X3OspAxSkWz0X1d4oED/m
dfeqeszu0aU77sZrPi+Tvpokwr+Xku+TrjxYfmXnTi4YyGRCtuxLEoHPkIY5
ESEMJV/vVYi865zth7/JZh6dEINLahc26TkXR1FasiyhJNcc7m3bAVPoVUDf
DZPCcJPS40m5/nHvWMRd2qlKEBMo7uKVmwTTHMkzL3WBUp+Dj43XaXIeeHQA
wxZjXmAfYjESqx4VKfSQ2yUVSMrmKKJRBhb2fMCA3GM9PzqsXgt0t2JcEtn6
nbGxZyA2XOXQ3gEHFBh7jUh8ueMwYsCBud9hpORL7MVNdZvlGposUx+6c9mF
/U++i4uGwBC6qP9yj1CkZ5kH4/H0QjjP6fwG940r+JJjLgKojOQmLURaKYbF
oJIDFFV+zSwZ5CcPiqsqcz8JU+r24fZM0pBLe8V4XpafKDo4ZHnthRUm8Xxc
TErf4E1Wi56Hl54sLHcmntUcDw+E+oHEDhJvj/tiYl5+OYf3psIFIDkvDgPP
ERIfcQ46jlzd18YHZQ49UzHCwbhWxpNNIt8u9NEg3xbhS3A+8TltyNTh9yji
v3YuSd01ciIgrAqYB5gAYFeAlzmOeP/OuEs6/YlFczGO0UnWFltIs891cjvL
hr4unFninhdiMYvg9K51kkU0ov2zxuG1QB5quYIfp8KtyeFCnv9Y2bfDqhQ6
4/1DMMYYQHUcc/zX5Ahaxgu5qsBxa740EOVBEkoWXl75ap1lEBJsD5X95QMG
x1+KfKiN+BmUcJRG8PERDSGe4PA+4OxfYCqvg8YYSfrLw3W3KwcwPcsqOLz2
82nihWl2SZ0FKnRyY9VbOe/SlhSBr1jzD+UqDcIfHuDL01EWqGOqBOE3s9ap
IF9wnnha5hVlQFRnLsMDIvvX0MUaQg2Hu9E7uZAVxdaBrlhp/pxcl2nJ0U8p
M3DPVMPwk1S4ln9X53WEGi28s70k5N74btjnxnljfM1178PyoVD0CFzLJZim
yQD1bkpXzIkucb+zkzAW/CGI82cnFU88L6zg7ZaOa77HfE01I9cNBuYMKV1d
9riib8i/wwVu5lzm2YM0h5Uq1Lt7Mk6QqfUJHZtXGaKhkpNUeIvOfHKpMiL3
H1m0ugcDHwDm45AcRbAYpJOhEIMa2HXIWlf18BLzXhwnb5oQQ5TN3rjRbFDT
xgQTNT81Wf2DOgzuMeX2WTj/RwSb2kZuNyVsWAD8QBurLPvRLtwBm+Ige9rF
qre7UuKxYIBTFansE0A1icQQBrVhp7zDrhsa2cccpUqZJCYWqPDtY3d/CG6T
ognagpOA4Cn7P8pv0yrWIj1XcN/m/iEEDLBG6s8qe6YNL+k2eHZgDCD1x98Y
nj3MPrCCTO64Krmjw8P8gs6ggOKBrzNzeYcgKBz4PDeuI/3GtlBG02BC0x63
cHDwV2SDt8Oxr7jQ8YhC36kKHBlUFGuQmRQXiBA9ZrB1Bh5svezObHjYBfO7
FWKRpRzx/wnJzNdLE59kw6cSmvnVAEBybmVubzL7H9lDzMPnnD2P3x5OcOT3
Wzn6+EW6FX8P8ZhXokxUAjL/vMIHbJUZuzymAlEHx+cQgZBBmoHxXryYGvM2
XHHfnClftH4p/jRLYbJgtcAzg50YToHAblS6JKZfCTLewxxSN8474ujcUX82
kgOH6+Y4UNUtShtlTWCEJpPcbLi2PW/LYCnkjOYpd6JfvMOvyMpywRBzJ4Om
3/upECvZehumd7p/7t+g6KvLYmRptnT6VH8Jo2itdegDwt1E6pvZAWwgLdtr
Jt3G3tZi4MHzcoWcn/AkJjYefJ2JsUpVCZheTVmbIP4s/9pm7+9jnmhJuPLs
8z2fJ37vYxoWK3Zpb4Iw0Mky9iTC4IrcGBOUcxVbFHv2KA871s9SIunplFfy
XfUXkFnxLSdAPMEr3eS7V/1dczKZJTiKJHc2kS5YHj6embh5O8MX6cwvAcw6
KFzMrUuFXK4jUZOHvAHjI0UZ4pcHSqwyDucuKlkRLqoDoNXQ2nq23mbHY0Vg
y+Xm46j8UuYsxc19F7F04VTdzZQCxZCx93Lq3MStzAkwAL3IDn1l6Jj99Mm/
H6KA7316yHQkuRkNjSY7rKfKP+JyWLg1lS03oNRqk7hI7qn4dxaN+WeOwP3W
oUwOy1Bm+yRy03P4Xt40W4JEQ7GZ0GS72wG5SRQGMBkfwqaZFxRs1/Qii8kh
C5wISm3mUAfNNLx8Hl4j7mjOH5OsvEdSsA6xikoKc1n2nU2UTHiJ/AgNK0aO
lBpQafhB7mzBzaD5Rmjja9e80kzLrRTZ3E01sfdIeUslF/5ryQQsP0VSlWAH
1X5oELjUUXNlaSWfvh13RD96eXVPNVZ9BeatZK13vgcnWE6BxOz8ZUaMDmr0
pRimoIf+rjfxAFtLNOQvGpWgwkdrt3FJkhlntaLds69IJo6wQ+zhlx14PacY
KpK+JcgNIK2D+4QA0JbMYVWIdBQmFGoFyUd1FkU5PF3npk4cexp5XDLHEijB
L5KeMEDP9zW2gOnl14Ky6He1lmkHXquYJPc/8kbbUCH3PqGWx2/4MPXk+UEn
crvE8JlVzlFy/gyNGuYQagYzK+WqWKe7pnkqv59X7kRQCShO5PEhxZ6aEeS2
r6puPTsEo39oQ8UDb40nx4WPKGn6CQExT35OCKENsuKI/pxnc9U30VL7L5xf
08qf9vJiJiZ6L1E+2RcS/xFzzE8UNB739Jgo0HxSG/Bl6aAErjClz3ZKrNRX
YcST4jyT+gLI8o6U70Lf4gSkrNdOnmM29bhbz41u5/HF/9KkckNTaS1dpbrW
S4buUB3rMuE8856sDo5LmC/x9T4Hd5vjqt/nQkJi36DhYOnmde3y0HU4vrWy
NAva6GgQ8aNJJdeeZY8Jg+MvRHOF0G0PLFoS1kpUu18d0KFEkFf1lAxRoNIs
l1bZEHsMpTNjByfBKZrTNFlU+o4E1coh1DPbGSSWGqYID+k0xNvytM4ungo6
DCPoiP04rqmdEFoXTuWo4KtSW3OtxhqzDG9rfjTBqeQgvHkgjYvtz3UPn03f
wwkPjkXr5BPh4/HC8iQQb/SVieXbfhE4tirf6BE17J8l+t9nOB7PBxiXSrq4
EjLkfCgQwzRqiDoQLH16LlvMduws/J8w1s258kuWR9YdULEbrH9jw/AsHj2D
00GrnKSdjKRJY6x5VjJJ+VzgPT0o8JZ4L1/yfZNJ7Z8x+l0K1GhvYzIlO9xd
+f77OTSnJ2epwfKTQfgSpFIDKI3vh6v0+izakpROW3UekHuZcE/feWTQIziW
1TDhLC78ahGnyV1L1YBhefn8ErU41lLTq+dFbcP1udpbWrotg6e38Y2ujRwK
C3tHUrMJC4YpvlkHFcJ2oEWcV5B1tqVkWsje+gLwkpnR+vL/y3p2vvIXUqbR
WGdGTC9FJ+dlUcK/Rm/QrtR8ajRuEWRY5bEL+QjT3ZyRiJUgZzy7Yx7xv7Fu
4yDCo7QoqrVprutqO4UxXRdPYP7kI4R6VPPB8GGkXeadhAbo9166SZFhW7Oi
IBHh4xfzRY5qwygtZ4nXfiuuAIRY7Z44cYrY1z4oK7x6WXaKmTbtPeaZeei8
Q0dqxuKW+q7jLkdZVTafQO5e4bYLPI5pjQhiUskR+n41jbSuIMqeMA1X1MSj
vI+s9bDGdzPnBIINwVCaiO7C+1Xr0owZGnZArrs897aRZMw+oBW3Oru50osB
IYYsGu+tBXA5PapPD+GsakG10DU26YvBwDpTZCbU1bZuEcWTS9pH1WH3k6b2
bwuPhcJvy/T7Lf1tt/DQEV5v5i3vznlwd8EvT4b4F/AeHygZu/3C3+f7ZTOV
J2bpl008ggg1Z6mV85iPCz/eGfGnHb8X4dcb5njuZCBvnrslAeN6T2URZveA
epjjbobx4rqES+6zvbM9I13e5g1laJhstq9k1TYqQWA3EJXthX+80fUg7x0N
oIiK69eRkowKlUhIDMxmVNq7k/ZNTtkNmnZnVWkepnupa3XDeB03wKqfa7H4
82nF+DkUndaUFYXtLUV/3W44AdXFfaj150MNqhT+pjYzc6+w/QYxk9X+egpD
J9W2cGKnEmNOYSiII97/vffI+FJ71TydmFZS5RjDBORpEccgU0WtvFWn9v+c
1pgIFDNEBz9AYMN4eHxX+tPQIgx8oCuDQHfmNaoXF5Fsq3e1AU388Me4AnSS
Nm+oWrqwqkBl84Aclw6+HFIL2vP/5NQws/fmEUaG3RcndraxPsrCn3jm7MGL
ciGvomO0GT9z04CrbsI9CmzRIUpXxZ8LIYgWY5v0lRSr2Kn5G7lTjqg5/K5B
nIHVL6UISKEAIxgvEJ9vJ1PzsOvVqHuoTKGODpDHjMqKjXrjLN1nOFPhTu9K
ZoA24whYt7RTLjvfDy/dqUpL5m9q9RhWwqwkhmVC0CeQPjkRNYro8yzqGAjT
B7qjPgh01TXTWF4xDtJXW9qNSwOzInX0th8pk37YifQAjQKuEq37J+I0iZI0
f7qXVqVIhZYZHARGMupmz1UQbbv717551MwgzfeJLwjOV/V1rYHT40KZw9T0
KPeEGY3dOrn4WNhczRy4jvbqENqvyxiGiD48oZ7wRj0t3SQ2HVJYJcvePkJu
2rq5mxWIOHDFKtGHQ8YtJCix4KXJTvM/c/wHq8lv/1HNeM8JHh4u6/KS/Rwj
d6vTPfXSxjTbA0+n2JxpIfTEy9OPQHZEFo5W9kQXWXXPrYlIZVLxRY6bw3Qn
pllt9V41QbEheqgItQCTSFzIaV9DDtFl3a2eh3Mu7XUKg5H9HfdU4iRLKMgm
sDi7hM2utJSMr2WZuKbRyALIDfvJVFv567WllfyjKSQNHCSAIwhYa0MnoMH9
/WC8BVtwv4OdXFJXfeXvfo7y74U6lpV6GKW4oTZzFOp2IFdAri7u1i2bDfyD
FjpsKFwYxuRQ2LeqoveIFBNWpEWoWbZMnEdSjMk366nnZpF1+vgCcLRtTzkz
wJ5/YtK4U9NiIQSU1Zovmu3lEMUgnup/qYu863cj3UUZP13YV9h4ZUzrYWZU
O4ksm0DSWEHznYU/5A7YIjXjyCudcJv8ZiBIV1Bn1F95jdMz9cfbfQ4zniDa
/gX/dvK2SrIHW5XtVm+Fw4USonKR9cL2Nzjv135GDd/+vsP4nkJ69qBnj9sQ
xLUipAsmgwzoNwIqaV4OKrHnHi+zXS2RyGSgYtfph1vpq9WCS+zJooDiRjmJ
TwRxOP83Pv5pgI2T3U7QggPW2JVqzKqaKrQmX7m2Q4XR7MWFTeySdwYjgoce
n1y6hW2jtILwt6Wj4OZQRpAcWRM5KjiQ/JYOPV8BiyBUHOEHbTzl7N0dMSut
XwcCKGL6/vEduenKHjdMgD0ZCzqPL8wQzaTsRE/MyGQbXmi2aGcSkeYUDjVB
/Rtf4sgDPngGUhCHE1hH6Ltx6IQNs3Dw1luRzbTo7AMB42CL6v3zsf5q0LCs
nnujirSj7CV5OjA2KrtB1Xr+cfX4muy5L7Q4KoUIQXfOR5zz3P7A0QfsysKF
LPgHJpwmjWdistzCkC5lBTHWD5/eA8NaYdFz80rvUdsVtlUfwVwltCuiayQS
baSJ4kfemLFayA/HNVbpiwwvYob6AK8+E8A+TnAeg4vZE+5Ovym8aNRUHZ1m
VcDmYfGGIMqDff54w2HgKSp/acY4WR/k2wOhelcGICUvw7A9ebyaqFbumAlr
FP7OeLQSpREST8r2ihUdG93x1DrYYPlJDhP2lxgHZAhWm7I+yUCXb3jpb7+v
cdnYFpidbG3oRruNlXfGAWPQcUEMsAIxxvWgeDSZUnFAbQWy06X/aTD8oIBy
U6NWGJQzNoqkhrXsFY/oSnwjLlD2c7NKO4aWtyEJwz1MraZmcv3yXiQgm7Ov
94k9jFqEUMLOloO1zOXJxRoBTwpw4YKQ+C8BXmB0DjuWWPPd5zfwrVK9ZGj8
PNzI5JB6UpxVcaADh1NlGU4R7P26gEree2vmWvrK1MdaeLsFpKFkFOBYsfMJ
iTFMqIR/gfmIIT+WvO63YtvSR2NOA0xG7mTZl2nCx00eeTT4Ega+vxzVSkQx
eQpaGKzlxraH3dzzIvpvN44RwG/wxN8P4PTGOI32jkwHBV8clsbeUK0FBI/8
6coo9KHDot+3D0kZxRx8Kuq4w+tqNUQSnZmhJjBNcxBum9xJo5XuRoD8AG5t
Ezcui5oQgvOw89r27vqKI4xEKhjKV7QJdTbwltd/2mfDEgnhETGLxosYHx4b
YstczUbCmbffGvZfCE9+TnrbSopeChUNkue82kxTADOizMovYDQYVzYxLMOb
/ScvD972JJJu0I4amT75npF3CLGAScn0hewSHmrODXiwj4JqtByJ39jrV9lO
nbcxglwzmoT589U/OsBTWDbQq2diu4zKPD6/PGMTO1jFHoog4irSrjRYL/cA
od9E4vWQgzKJLu5PQ2M3/xDjPgeVrga4VaKJJhtK007fjAL2lXcM/T5TyY5v
nz3HjHG7IWAIvbnkYXm2EOg1fosVpgUna/gS2aPN0U6RXcmGKwbiv97ereuV
w/vQYE8eRPSBXfEu7Hw/TWE4nohwQcYPDHqfFbWxRZgyVPwDJiRGHB9gDJpx
B/oUll1T9uqauIl4NnRyzwvdWaEvqXbQvM8kdFsoN1JEHaJZr+mF4pKROqi8
bOGVlBS3RpILVQ7LvAQUfSvjxmIpRPJ2PUnFgKq3EMs8dJYimWvXOP0amAHf
cHxajTb8w+28VBE2p1lqYcjyXdfpMXJSuh6+PftkNySjfI4mTmdPixz7c0gL
p1smvEiVYGtr/OhjEj3wKOgh/bJjwsX1PiykfXQQHlgHwrRJjlIDfMoWhm0W
tboWYx9y3ONXbMtUVtqUXlp7IkykWiUNjwSk0MhWzRrCW/zWCUKhUMiAZiPP
5X7YEDP9wByWd4AaT81mSfSyM9ssq/GIOtpWSi6809CVXM43WbDyFP3ZdwWu
kfmQAzu6NUBYV3Y1IkmpFCenKGc/eUrygADjqJIOoHWsrPBLAzjA3btamXKc
vJwNAuqOL6/aUh1yuSsSqHxhJYd+ScFywTPB/sGOhybZz5s9IL7H4NLceIB4
qYomXUNB7X7jWIkbaygnzQu9O1FC1SHAh7C8tAfu80UpMe1j0t62KZM+IA+X
H0GBwQCFE3w5qhh+AuP63BZLDaUozPxukvk2/KL9YAXOmymRQhXCTWt0F2Uh
Or2h2R1qYsGEHxpJLcb5mepDNfdUSSW90W9FQU1lQFKUvaPrFcGKBMUiO3D+
YA8DsFgt7B5M+aZ7Lhxjjutb4hjbcZy9jIX1+CEMJ3SxBZ0OK9IMr0wViMzI
qy1u8TZzKA2KMpdU9q4jXI8rKUJ9zKWfk8ALKI/y50Ov3BaIfGFlAdQ7FGh8
jA6lnhm9yT6NOYsDf/M5dDLfL5y/Gox5ttVzIUYy8mUtghvKEpfAhEANbr8V
6b5TrVayehBmVNjrIFtWe9uIyuJI+Dw3Set7xRP905IhgZsdmmleAgZdZJ9/
rCnsZXRIRPjDYrShDYUFwiAcPRYsp4HkWIMe0icSNBFWlxA8yGmQLiGGYVo4
HRGlWSt2xHYDO2bIQWp9gNDoqROl4qkFXhiUkxovdIi1oQZsiql19tGLp8XQ
r6alhBBSrf50VrXe3yikTMiVmATylXcwxJaMW+VdtMaKh2MIDfTpvvFk7kur
JESBfQ9I+aBC5dq08AYIHRjpLr2WGm2l7OCw1e2Y7xCpmOgw7OVg2y9PVOoj
RRCOLzsi5dWISrqrEuRLKyjAKthD/ERwXaAzNrU4wH6vjqybVQqqKizygdrb
v8Oc5rsBimoR1XEYFv48H+v29R7aoxE6fZfSn+rlQPdDYHwr7tOj6dhULZ5c
OHpb0JD+ejozn1+3ykteStqX3q0v5yqfc0DSl6e2c/RjSIqWUaq4IAjoSFZi
QyQT0hIvvoF1G+x839eWFAPTp62NQ6GDqY+QMDsB73EOop42Q7gS4MNsY7RY
0kNOR/op17ms8Ral3RgHllI/3J5z84VHl9uiidglt35Ii7NQTxTudjCPPGbr
O4h8yms/vLnzVw8mw/k7xMVaaiadIm7obC3I1IkFsgSuZgB6qt3iPFetscov
HvEmSCMIwzPGheHHEUu1W542r+IyJr7oDkEXZquI3Bn2TRw6JL8otX27Buse
g18jtiPqzxE/H6fNsoJaN7dz9pvu0NhfVNHmKYTMc2Px927Ctv40bJJmxWDb
Ke+hy24Ga0blmlxUP4K6T+zJ4x/ul3Kd+5rQd6bm1yqjeu599yEB0XTCHG/3
KJdBh6Ck0lkObt+Y17fTRDy/mGXJFa3xB7ajrG6bbTP3fa80PcbAAXRuRvsF
LL+PVZinGUhnH7jatfxsU65FV0uo5+8+hxFgwvHMlX7MweFLfAFd9psi5k6U
ptucUVWI+acBxW9XQukgWUncVJXx25HGVtAs504pdp00twikMEturAgtBnE5
FKofF1zL9Qn0koRv2IqRiRR+4g9EkNku8HjIwMr7tre2BVulq8cfzQORlQyh
Gd3tNXcanCgR6O7Gt/aNWwRgmsD2ECAASicdlAjXmGPFkvzlI3Syywnp4CZl
o69BFVC1szGBZSX3OYLneM9ROeYyJfDdQWnDNH4qFXRBQ9bHcmwEyi/NgLbH
mpTx6ctfvm++KDJPf030Ks81sR86uE7fvDxkS9eN+79PYs+fc8lwCefVesBS
3zOqJTnkhHyGCvIBpR02VIr0ulO3qhXb8SwhAIyNe5pIENl5t5Kt7ajaDIeo
RMNZyP9rSlvK3CEjoLy2Hf+eYrZF3bFZiPeb6YDI7hrx+PV1oJ1KsNGSt2LC
yELMZhD20FtfxtXHfSsug82zj/ZkkMVwrYANuDkigvIqBQJ8IF1/H9GI8vdG
0AQFYVWJAIQamDYoq5QmS0q75Yl6z+h4ObJs4OL/DbM9y/uuqP0/I23U6gIv
iAcoJZ/1Eu0yNBo4DRa0//B9uYJObK8ibYW7hPsV1hS2aL+mjh4SJ1tkDWLV
bNqb0iC6IVOaiWrCH+Xk5ftKqwIuHiNbIsdWM3RSJickueTeKpbn2AHW2xSq
DwseovDtkqoTfoCOZqBBL8YTp4IGtGOKfoNxaQZEZSP9EBXQ+J0yk62X1Y6r
soLDUIu8jPJ98+ylR+/RB+MkgO5AYkWbsb4iDDKDeYmu7p8L9u6ylK7Q/pSa
hdlukUzQiAkdaMjhyWSFWgluYKZ8IlroUy23l3Wpn2bzYflQ+Ta8ZuGK1i4e
/b9netORbw8K4t23Wmntz7XFzNPbjalulxZDuM4xZMePPEQ3GVbCdC6+lHMR
hfLNmxVthcZVFjI1EtecPttDtdIfsfm1/RVvWhe1zX/6HPHzsrL0BLQhDFCR
UZKMTjE6OiNpFwlCKrC0G6RCvPxaVwIKvFBhWoGp/ycV2MXaUi+sbOuOS0EE
IVm0IHU3beaFZjzhD28Uu6SkJVkz9IRnu2ez1ff5xBEkUKi8dcHTjMVf7d0F
NVWzcUTUOkNPM3OuiVRbbjDiz2fy6H42CTIlaiTyZv0mkYH3soTxYew7Ixe6
BouUcn1/aqQyqbpS0p1lUhaoAufJiJQ0YxRn/rEocpQ/sNLVHWw+q5AgO5RU
U0172LVJ8FcvYnoZVIU7Q6y5eGDrfQzH6d1WPVgYcY+cv/viKOCQn0ekpYEN
a219uqph355lhe3nVukgNlquTfwhGCTyn9p2Z2d2KlxA71PhknXtOpzBOMI0
EASMGLUgh8cEtZMkfBhNdz5mwM9B/MLnQmZGKKfGreyfJ5SKUEt7Rpf1/Gzv
hcO5faqz9iV1FTHYtfh9/u0Mpdm2nqpmqRB5T8fpVdm6tRnf1OLneO80x+Kh
cqugfeeA8pfZqtW+QEsB7E/+TMcVKJUaJjBj2C1YIYCkzJqg8ligmjDBQ/56
HkNLPghLihstIaXvhPlP7HEw4r7qTlrboLekTjghN/Y4i6CzDQMaDj1IVNmP
bSl3xRzhX8zHzK+vDRGvjhV20GQhoFZRtA0wMv0l5FJ0G2gk/E4vjoGAT799
JnV8gD1ep4FkAC9Lf7jz7uQL5VlbH6WMZ7zgc6+BTFpUEBqaukF+x6NnlwMe
QOoYad6UUm3WJtOklnhzTPLfYv64SpYMxEETWevRM0VFBOtAfYDgMJZN1nPy
vQ7PlF4xwB72R4VuBXMi2HfAKBTwLhM/eWmLDbrN89zKYzUeGtuSpWYnbHUw
Eq7UT+4Ucx6ndcPbqyiBMei/WRO7AFETF+IoOYA6GFScgUUHwWXHpOgUTjb6
Zq9RMbWgHB65WlIFzDpSti97yitmI9o78f1jsQoJO7Agda5x4xpvD1tCvuAj
8qmBuM0f7j/S+8xeVeR97pdWY3Z0QFTde7K/VEt5wyBduSC5KAHNmLyOWXrS
3eOqove5t6c5AiwiGONwa/PsTNxuHCiDo//73vyGIbLu11MUU4gmtpDIOpfw
2nKqYZlE3JYtmNobRVyrorMVOUZ0/Ymxua6rj2350o/z+tYy2YYQYf9Qz8oJ
Sf6rJHuZQKUk3wKu0aoB4ySaqPuzIHA7ckK0OrOop9+RfbMex35Q7OzxfBSN
aWy6FCcbxAn1SWcLhQN0mHK968IffLSqd/QwAZjDnI56B90mDWwhuJUVJn2x
/iirtEM8WEeBD00X8sUAlni8Azt0yeiJyaNxcJt/pTB2meU3i6slEV4FMhYY
c/tu/NHM5eatauWWrP5XEtekrfSYOV/a2TzqN+nsrltWQDPWok9GZoCD13ed
iMpgnVM/JEv1EiFzA774DawigHilD2sSCq61nAn5h6BCdNLSes0DzlQyB1K1
4UqOLTSztYm0J7zpMx7hQh28OmmRaynC0Xl8OGBjEv+/6YIydLqwPv3FgDvj
1HXI8135S79IohNRYb6giLaVWuYAG+D/DINac0wfJLfJnLBLKFqPLyWb7r3G
2CeGpyx37M3jjULDsCMSS6xwnzaX/iIqLiqg+RfcbRr+jNXW2heXSo1CMQCi
X9dqiNbek82Su9FCrEHM1CYxF7bRqXJ09kNSpEa/y6jdtcQFkNWl3CT/Zgd0
Xg1hcIUHIP5E23I/e/LPY3n+XkQiQyUWq0gk2kQWBpfCKzeKnO5d6OYcCTCT
gAJVJsbWn0gLPSuKju0cNn+Rd4CFLbbHpPjIf56znHrCDr46tfq5WDzUnVtJ
aiHh9BsJ+HQ5POcF+CGIrl18tt3JIo8NehZLQGx8uBI26JfNNi6/kFNX0CAR
Zx0F7pxOusb8QPCEJi/5IE6QEdF++aYxFm3LdPivwE4s5i04Fe0R29pkI5xZ
UTwNUkG2ISob1lSxcrS9BbDavHEgjftIUtRKeia8fGBYLI8p99VpXCRMDqmO
MZeFbGuNNBnB9FTUAB/aP/zVPBOC1fb/84tV3X2iM3o9WU3539n35FGQ5P7v
uUF6xxguvzreLEuHO96K4eni5+obzO7xJR9jFG83w0iYhDgOruwOtlmKRdud
uA0whyzkVUKkUEipCM4iTq20gdHaZpkTXnzg0x5ed58Fpt2U8ekkO1gvYxuf
WLRotfC29F/tD5f19H9qrp1FTRCICXM0rb+mqJ3CHKILzaoEh4ykfL6fuySm
kDfrILHPe0zC11qc816XfD5NVSJQ0C3G8ZlycoqtLBZKo54Iu028Lf9FG2C8
H0MFYT4JXrUtnA7+OfWcvUSeV/Ta4KbjDIRbf45fq34lgHFaJklIw6TYjZfT
E20mvhBy89BiEQBmqyNvgxxwuD9vkDXKow9+o0iBbRnnqRy9BARn6tz3HKBT
G/0ch2S51H1FmtVx9iVrhkoVoqZVx6pRWyya9yO0kLrCVxbjMykfpxjMvhOq
ZSVTuHZkyDrnwc9yrBFw5BEXtbii+P6o+SWdSvmxbMuvLubrbVfoomDcADKy
F5PZU0W6i9IxRaNwIQmDLbmEbGQE6pleyhNu7WXV6m7qhEHV7hJ1e4IPxKs5
tyVPukFZLDjkK8DA8hdQk8m/JkDmVzLePXH/hHTTFQ73vog/krAMGxg/jG/8
GrNPyX4D5LEtsKQazHhqo92ROElYiOZZaXqV15RDZU3utac6vaxZ1CKrAXCR
IyAzmnorRmQk/Zp+vObumMNbdOtOla426mAE7uoGtiNBt3ctuFq8ttnYmIvQ
QhPyaQRK/iloSC02zlkZBdO9M8FCwMzFqDHDwM5Lj26qSTvSC/NGtswbYjU8
f1hbBK/3NorVET5gocOP2wuDu+4hk5rX/QxCodSYxlolirG8RvIuSSMYlADW
hvfrwNak+FNxuzodQSyYCyg0038edr2R0DN7DfrzeCk/7QqA5aio118Difz1
BijHs3Dgd09mTLMcTZknhjZGuFNZqhF4jc8bAz9LszvCFmtMK6sKtNREigSy
kBH9GG9hIfZ6neBWRvfI/w+A4jePJdpMi/uv6NTk3bNBwEX+OLP1XpWCr4OR
p72EeyvPIyA924XkIOvfZUZsIOBOcQuIsgntkPaZ9jXpgmlCPkUf/GqiONoO
mEQM6Rw5t8EhkmmyQ9/mZFSGbWOD5F3z8AWfdn67v2aVjjoPu7u6GagSu6Xc
6HrzH9+QR1rcBen6Tkhh3AeRYh5MkLhS8pdCSDkH1ykvxSTGagq3EkjIrBzS
TwJhjz6umK8nD+c3nqX/L60mFtUUpBtxCsgsQ4RoQCFtzn1LCS+MUUouZJ1F
e3XmVm+BUykEfo0W7Jv9str5CrSXt3LVMBQutMi8/EMSVhwk4bgk6w4hrHr0
aHQMM+A+T1d0viKQYhOeAbMB+AzjMoTFOHpv/ZDNamwuJFWKWTbMxcisoKbU
Jtni1m8K4ivwzuUZTf/TzLbpx+BhaSKypDc26TV+1mzZRY0kgzTNLeaquRaw
NzUVgLew5/Zuc3mrZkcfb1cX2We1jWl+4fAEqSsBr4dnvexX5PDNVUSIbW09
1hA+Mxz7PyOtyI/kfXM1h8st05A5rFyzYscpiWlQfUzVGcMeEO3VRyi43vSh
adA2p+G7Br1mskNWHdKq/TwtjJZ0wf6dUGJGgwwLJVsYjaIK953SdZTxTnxg
/1WwC1rteEth8ErJDDobuOF8sEkAY/wm3YWt8/hz2S+SkeAq3XbfZheBg9lm
OXvR3vLcLIaEQnrdzwxXRpw4wQ0pGsvomjykF7zVmk9c9jKStgHGI+6hiNDF
Wx4ZrPMzX5u+RovNhoOm8pc02cmnGv73Dj3Y6yCtWg7HukAtH32NvPp8Fz3C
CfHqyrmJNu8GC/1Hu/imcZ1GvUc6J7+8Ht1STWp5VsRIlJq4SV08875lSjnC
mZvru35ZV3nBf/nB6jFT/qZ1gszjw/HrVnK4HcWOUKuHjJ00gdyS9ltxqXk7
UnEVE444SV2CGsXI6+abUpdXzHIpe/whPw7OPLiEt7GbOnG/Q74zz6RllqlH
vVQlLKNaohOQQ11R+TPYuqM+fNALF4eMzE1NCj4C01Wf3jy7N0TzbAfHF6Xb
NdiMehP0kmkKR5K87jJnVgxXvX2JVOON05NwUBkmxRRz+lGGj387peAVHfNo
D6PXxO/xrLp9jFHeNfaAgP9DgIruD7U8tXGWclyxqW19dlx7GKXme7qZvjkt
Nv5nxPSk6wPKi/c1TzPFhqGxC43f3+1dV/zzk6nTflqc59ANANUyi2iZ0Ccs
OT2ZDHjXxvsV2Z8GEXz0soqyFHUfhYn3+RXx/Jxl6TGg9BZFrRfemqpelEv2
eX7Yx7U/0RGND97bjcqBbRmnwqyVP/hsowU9F1ZyGRL2z1M27FBVaFTDqODs
zfEzFTxNA5dycP/5qQOK6Ge90YTHF/tMhHW4OQeKSABrGTs0qD5M4mGOtNw6
aD+F7/J5sFQ8G5KL4aC3Eto6kLMlum5hH/gDu4ZKPSpFXxSRtwaiDJ4wMP/z
SgENIeeO4x5COAcZB5MF5LY9jxq7xUU2FyUpj/rE+YdfaSrR0L+2ewz66jRK
b9zVe0bMXlMxjIXhOhrdYmMfVcnBrD/c4Vw4fxmvlBrucnn8kMUd39aYKXZj
gF44kIAr4q694TfGzt5Xbk4DQGySTXkSiercghbbxo6vbrcJm9XZazoUQ9oW
++WMzR87Bz8hBxjNHV3dFBGOaBaK5Od0JJ6srWOADbxjIXbT14TIfaQQrKD9
nAhFqJBjbhhI+zld+FgxKnMYpeUFaCCSvqFENn0rReMPT9FCoVDm3hYmSLVX
MOH+zesnwXF30BQ57ar37gcgiCsHrPyRlDhR1DKtMFPsAhSymR++u0WZVEpZ
byqtaEbAFSW11P/IiF0wtz92q4qEcVKXqS65vFDR+fgaJmFQIVxqIGO/wZMw
8t+Ft0w7nR2/dFFyaRFS+7kgxrzLvN2jbR82c8UPW+wb3qVejbCrJHTRRS+L
1t+Q2K0tk+mebbsOoX+raUZ9wMb8N7mfWFDMqNDzsFI5KLhgDMKJu2DiJQsg
MlPS4MA83SXarb0H7ZtFU/BUhy3TVGdRZWnYjY8h8hWqJD4cKUv34e53XRl0
BazylbIBxF+LrAgwnv7pwI3QxVacAcwhxv9ugI0MmdrBQGYVwk4MoHsxyHkI
ub4Xtm9we/AghId39KebAQmEVfNTEruiqCGZKOcZxUkhyc5JlqvizgIG7zX4
L6y8hKUqfkklEyXFFZ2FEGe5hBwp7j08t8V/mXE6y0bIA8+GhgHhXvb3+YNJ
y8MN1vf+AGhOzMEVW/AoNPk1jcR9PXugOHrCGPvEAyDMHnNAtFeyRtiUXNYI
HGqYvuDjKo0mYmygcW1RvknXK555d+8oIDTWfYSlKMfMuOF2u6ABHAb5ixj1
3vzzFuQpDYRqBqQ5s9cH9BH1mjwj8PJA+28G+Fkh2BE6664PZuPLeltXsxSr
lv7IcivDaqyQ7VXWMRqXySOTfwL6C3Sbwl4SECAzUfQdmYieNQbi0UGdjfOl
753EOZz4PycsQPaskI8z9zh1j6TELRUZQY2aR1ZCH8eDs0lB10CEVRxrP4Af
4/SuDfXcPwH4C/1hhi4oDLmkklt75XbZoPTGkT1m7B59CxJB42U8fBum/P82
qW83D1rgiNRsZqKG9TWYuKTWS+WSxJ71GSazcyit56Q8BnvuIk1v+MIwCgm4
B5Z9ytfzGdUIbONyUt/d8Esa81q+tbpj7oIgBMXworC41QGduGKkFmVN2zCm
/GxLn3bkikRPjx8ftq9ruFz04wtEcGQupXXwLyKL5VQPGio9MTV4l4zFF4CG
iVhUOGpp5LVdOwuRxrnRHFkHyTeqvkak5+WYNmIAVR6vHVFkDBLAC+0nM6yd
6QZGcvm6MmTQLzCF9Fz684JRqjKAk+oiSujm/rp8UXSFAvD+c7Ct0r/WNA+G
p0pm2lvJaNGU9xToqRCvpHjCm2tfjtCsFMxPWflOEhhoivBcbUmiwk9h+aN3
Rtp/LvONnsUgPrsn5HRxb/PQJUc5a7pNzbTMMDq3qembJrXLFG0V9KJRCLXc
I9xz7W5qhfw6z2vW9pPbvqe4kceNQx6aywIZj5WhHs13iUpiJU6bGnf4XaDy
ioy5XSOwVbapurAGbsOaaVflCaYXVRYi01YcKmTKGcLrnrJvQm68uGElDLbz
QGCQpwhiSo5FsvFtUfkG282QiKFM1JyF7/yxf0XNPCGTCEtqrSclg94lpGmV
OdMItG1K8zgWw2NH3E7ULtBsreA8xC0QQrlZY/DsL5B0K5pp3cbrqLttyDxV
wE792YD6HpqUr7Z4Np/x9x02crRSE0Pn7GF3um8xJ8YgtN0HAwZdzaN3YK1B
S/pHdRazRqD8JGY3Au/UniWXPTKvDe1+H3giRnY8s+JL4HWZCRfls/aiT5L+
c4ICl5g6LtmDHQD19sN8jt5VqjxgZNqlqfKfdaTRWGirZm56gMMQoZi5KCed
xLhpjxSD1f+q2s9/a+AGjMXBx+DEKMg2MxvkpS98maD1vZ/owQroXnwV6Q4o
/DswKBmv5dxfwn6J1ktYzXfSbcj5jSwzk/4Ctu4y7c9XZAmM98XQFgyf/jrT
U0eW7ohR+NSJkWDnIvoUUp8NqX3XTLB8Bnr3GzTEYdVCFpLIFYtuh4JMd7XO
8AgEKMzDlz7VgTNRkcAxQFpQHbpzG8HEvqHjC3Lt83EwG9hZHGK3o6dgOMwy
EjG/n2X+igNSg5KjOZv1ofMtgrRWhj1mclCE5OVtovmAwyhURo0dM0X0NsI2
mKyjd+ZRO3UAXEEvPaVHgmJ5blCkXLKt6tRY2D5BlO7oLrgPvcjkZsJkA/+u
YeEruSc3ZiOgWpWxh+lkOoyjGhgbh2T2iUJ4Z5u1I8KMdzru2i0cvIQWEpfE
7+eLYjA4OfH3fRvTs+s9wKCry9mQYFHWDWRWFGEpdSltvUadI4TjqWLiHiKD
d6xVLAf8Tf4fs0szDLhCTw3ddIHaAZtdNHjTiJ8YHszii+YKAfj4NnX+ND9P
WHUGFXEK89p4pu9G9Ltymy5Y53Mtb/Y34DUdCEulCZaSATlhqTlN4CF57twI
ZPosEoF+YDfvv4Ly/pVDfh4OudKAI03mtMh7T1nLfnExuvTqSc7loQpvEUBF
RZCs8HI65TNqzp0zs6Wv5Xbdd5ZUZmJNkUV5j7FxKhbK35DS56JJeVi85Zda
ALYPCQCiEQlrFQp3A3f+pQJ3Fj69AJJTB7vWY9oNVaIbui27H9psy+MqhYX7
pWj8ncBhC/tuXXjJk/UFcPe9d5FQymvtd5JSkR2i5A84nyTuJoxWBF6jtP/B
BDbEJl+aANrlI9oJxZbuqJLjng0oGwoKxuhGIZ5Ph+o4lwvNb2vwr7hQdWKT
OWc6++hZJLerjAoPgH/v4EODCacH4cO0WRYKYp/Mfx99zU9g5bAKbovQPbYI
ingQOXc+UF2Er2cGxoH3+4Vz5yOlBPQnyif0M1AtFSM2BCiqeOuf9atL/nyU
OCL9FwO3a35GvqSgz5YTSSiiF6W5YsQcb575ASqKi9idyzAkYGGRimk8PCn9
3PEatyweEZOU3sAHwurpBRS0mzSnNWdWPnNyVgiMcs0A8xikJfylUTE2gpck
s8I5O/xKsxgg4Iz3fOrFwK3400iSobZh0sK6J3vR+l6uOWdiwy4KCbq1PJI6
BYBJ/IEYYpylOKeZxcgcUbDT79s1U6BgJO2t6wRZPFz493IVmJtfFqQ8Ksi3
ksCreoMXGyEc8gQnWszC6znrqgvZmYJ4X+yQFukur59xcciMGRhGf1o7ulrZ
F1BMS6BLeti6pMbn/fxkp6ui7IlF1ZKMyg/AMcMG/Nl43dhALMDG7BtVTDnb
B1ZwAg9mYQVdqWXfPxH+CuFYOju2mEvIT6AebnbJlV/LSbnUtwkFr7uInGIU
ZW4hyQR+IeeUxkYG7fMA+2ygQDVonA85Qeyp8PoAV/pHvGSKeIqpa5FkhzFi
i+V1Q+1p+CC5XwRVLBjxHBm2/gQJ3DZXJ796pXTXj+LUbr2uX1u5ZCBgmOwF
vvaW+bJeT0tXltYvszjc9X5MMwggH1cH2d129RM4aAtMjp408S1mQLeOjROA
9kPh+32Ca8iVk4z597/9Xn35WhNJPX76OyzWunLogcxxbbBI0QHbhT4lDCZy
iHC/kG2YT6oFL2bd3p+Be8LZMz4EuXTyRZoPfcDM9+8n4yqbBJE2JTRPc8Ml
+1hJF99TSGC+U78VIVq4v8jQZyneqBepBu9UZGA14b59UNmMGnaPqzM79Dmg
wPFfNtQ+BouR4HsIBvtIxMW6z7Se75+9452wQ+1uM0h/YyyT84+MYbFkF5xB
4H4Hko1rOeBicFyjHrqHuNZ3TF2p7vJu1j5JYF+kt2QVpUdxs1uNOAybwrrh
qRLusCAhSETEnFDWa79cgXXTB+2WNVAd961QHIS/XjXkH7LT9w5OYJy2UoAw
Xf8HE6MO1FUQ6avysJ0Er+i7QaDDpvtsQ2UWzVH80SlXzatUsJa26hI04lQa
2o1XM8JPCdYOPzCtp1GTPY8SMv3tCOre9F2JGxltw8O5miCrPIYUu8l2LYE/
kBVePmaEwPG0VioMs2aLunsYoqCnfCBP3+HcFP7ml0M2A+z7euF55qTXbuPU
wfN2G2l1ICNml4biBwEARzI4s9dkV6fUhSUyseqwC9rrIpXIt6ixEZhKYaNQ
HLF7nA+/9O6aFEpBt4+cRUyDYggQhvQGZOF11rfhWzGJDp89c42X+2UXZ1ey
sJVG5KP1c1Wl1qxiYvLHehxvvHpsU6nvN4BE4w/xc0smCnrdfipr12tCi8tI
bciT1dimhXQqoIz4A3dRJ6Wf8JcFq1cXXK9CVCSr1L7GzGo6V6vQQ0gyJbT2
yT3co655PnqPOr9ljlyePtUx2bX6rwdLIGwZ/jCm9QamRIz60QlN7pg/wxf9
0QWDgsfg7EwA1wuj16H73uQlN7zz8JenklFH62halTJYotI9G5nTG4GZI/z6
/9V91ZFLM6bsXHz9vy2DL8NrZVtEyPzsmQZ605nv7rvSBO2UkY9GEfV5uyUy
x0CR/mYAzGS27MLw9OxTiW4cni8gmKipV2Csjm8aLgNb3C9kWeL72vmPlCht
Hqr6Vg59bIm1FnSBiWdkraiqgWWKgff+F8lWD5sZJKlZkcFpxGldUKsl4G2b
4L34PRFQ+GsC0hSdTWilFu8TdFHfgD5O2lLwasee9BJkKiSiEYzogwYBKpFV
AxdPUhfyKoxPUa64gk4wnNqCm2RJCu6MBUg7DpcotwJ0SMmEC7R8XdAVROyM
JPtTbxn37CUWdlegi+DqlrPa/yaueBPHjmX4qCcjFOWBdcuCak1ISYgA8NWE
f+mdmvCtYh9SjniDznLR7jNhh+C9FG8BoPdB2W4kmkRUzggvP4xC8yvN2pho
GEW23fie7MvuUYMIeHGb+3B8/RGcEHnTtxeMW41rsVOA9h3XckL2kTXXrssH
c2a0jU/lHnq2rTr0JwaXnr/pdV4j9ZkMpXp692YoR3374u9IRjFniOCIRzlB
OjxzPMzCp96XEvOj610mNiAMWEZnkdt3EHkIHNXin2eoNdYva056xlrdACul
P+M/iqnKXJpOlFSyX4q/J3alUPlwV56HWpNDTV7s7GaIw6ADDFCOvDoFL05z
2EE5+l/nQfi0ghdTqAsfHWYiVGfMoGFyWeKvNed4+AhS3c00I6sxrxKGOP0t
Yff4RFp6rwmmo8mAStRO57NH8vQ8v/bv+mqkuN2gWLMW1+ysS9ZLzV1Y8tAQ
YtkcbnvsbX/DVVM6vNkNUPDwor38mNRJRj7f0zlOVHpjJv/uxv1Ze4j5E7mW
5PTqv4J++Mqdkzp33GF6vFI+q0WCMG3ZSIYt5F1OgBmPZc3KaHKEtNEZgQCX
0BWxnhIfmAE0VqZCB518SLHdntWNDraCh4DD7nVaTSxOj7V1GQC2rbIEAWgz
aHVuQFqrhcenmjXi0QqI/xaloVzRW4Q4i0OAUrYVGcAWuXPX6DyM/LxuDxBR
5OezlYNU9yZNS72gWQ1mluPrdsp/HlKszIAWW45w1bcsGjJWAy3C2zuB7Kom
lz3FSCN+zZrVRzC2BuzLXwZAe0ZYDGD96Whk9b4SrU38oZz3vj5q7J+nYQ52
HVjy3+AMDATTxSvTH9BYMpazTLeIMaU7qsfTL++1dvLSTN5WM5hgHcqzKmRy
SjBbEw2eWmD6EvM+bj7PfmUpcHjjGJ6gMK9/VTj7G1qJsYj62u7er8o4aOVX
9/YpxijyQI07IjjoKvWmqt8fCCgismLYv98+pCPq0ETJZwN6qoa8TY5CEiGg
lU6P2VR+1mQefa0V1ZRSAKzsVKqo0MpZ9JcKMSsWX8I+M4YWbiyp3qGHxijW
/Fs3/984ZRLJnzmgJtkIsYT7n7e5DSVEbvMXe/lX9utJxC1FpG2lNSsPHexr
Y0hQHURjzL91jsqbtTL0aOVfFr0Kn/vQW2W2wVSTy6l1/NbRu6jI7n0qMsdT
g+GBL+rZLh4hzb0ZAV/il5TV0I2YW9dD4zU4GeymKVuvN/r5Wn3ZyKR3ZMVa
ag8Hbme4qbeZEURRpe66v6cYFwM21ywrrgI+ts7PrWUIteFkrwewlDAHydxB
Al8XLSaIxo/T8asFvO/Hwx3u3Fg/TddGiytSi8haxcnTnjqsRQbLkSzXv63F
pgOGaAOMCbavwHPwUZGajyRe65wdcG9XZ8+YYMPL62SYVjVK0EOaxwFzx9TT
WPOhhCkVWgxII3jSFP8JOlslow2Qyta6JLL72dmabjKIOGz7We+jbMJqxztB
6mCZNgCdT8EmrN9YFJnySaCOtnDT35OPx+84tT5Ned1wWKeY0Qp6u+tSDvD9
9UUGHT436d/AdvCZGCI4nUR5qmKh07M9eTrdMmmedkUEptM8Mn53wMAr4aPY
UFUE3cHu3cd9qZdNxZYyIMSwHnbY6LoHiLbyEwsO2bQTDQv+2V8GvZqUrRJS
CawKKZKV1cQfAiNiiDPCd7u045+lVJhywA0EKIl0SEFir4Xh+TuZpG8nJ2Yt
Si5kOM6I+M1py15f84/hG21YJSAgnkJQIEIweTZmHC6hlZwOCVkOgjMMpf6b
1kk7C0+J1rSMFZQusP+e8aGPXdiA2sS4JcaG3jxtXnxXXAcagUdtQEbnZx4L
YTh4JOIDBPbgBIZL8pcBVilF9Lwvngk7gwhGEX94pVcDqxHVEhOntQow7EXo
YTFJal1YkGqRAi9So0nzWv8/vs+9FHGUeXzdB4x7HVeOcnlFZVe79nhrIgt3
h8R3fUXwpNGcawow+I6XDEgG5a1VqU0L+DFTxPjb4hWUS5AgELrUoBv1flTH
9gDB0wwT+FiNHPyM2PcftQj0XG4VlbhTc6uUznEiX2naZWLrVxVfn4UZCAAQ
2bqDaHNqiL1hZMKWTqScvm98IG9Xp3d6NCzsfci41b1OGjEXjttf610IhweW
BTVMTyG6T0G5EVGKjbCIqKg4DMtG3J1mVJYnUTaMcInay++/49ziUx4y/E8O
wYgJqf/PxkNBYpkwUPCVYPmv2eLR0wi6ybM/afs2d648mzyxpUL3plpXEe2S
2f3flQtPp+hRpmmlAGoXrbNC7M/ybE3uXxD0hIMcNCCZSJlspjJd1nderErL
vTU4PEprrYLNBBZseAX1rWxone8QEjGpQyE9hjA4pVDTmGfEdsGoR2ZA2IS0
Y1kceSyT7GmoFZE0ieOW1RoVdU82jPXYrJAHT2RfbGV3SZp9YqCmIEyQpvT4
1cL4XKk1MAwBXEJ6Vz0cG03e6mOKTHD9SZSYvNIpyvIHNT3nFi3eM2Qvzjjm
jHxAA109CceNGlHS0LK0V/3g+fSO0GF8rTwxoGjkzxP1ie4aBUDG3YKl7WYD
mUk4e9fiBuJPn8//nvIbavcQiwFl1tG4/jSJh/499r+cH/98sRSHFm/xZfkN
/GVONzMaKG/B6JHW5+BGEFJd6rrHilbLs2/FMmCHbVB3Bg2pyYhnoEgsUu6V
+mPurvNEqxoKa56Ph53Gdto0MRCPbazZO/AU/jv+GfXOb0lMsX/7K2Nvtsk/
7hmqw3q8nEIdNtqsjpCIU1GGR4P9vZoZEvq/feeOIsQ5sw7RDCPR9n/Vn/KE
rKMVVGBAHwhKQBOazuXp9b+3jsgRoFXkGZkW6gnrCqp6iKFRDhSxVsR+5Ddp
RivbcHTqJHZNxLkUDSz83J50O5I+Ckz4FMjd8WjbAXIz1LXfAuWJ5MCMAd+L
EVNJREeMRTrBVjecWs+vbgI9BY2T54IYmuRbxPNEDkpjadyNil7E6hRW4Rqd
4ivLZeLCVpJlq6ojtis9JWdlF84jXcm8kHnNWdTn/qPNj2bI3OSSLZk6g58q
fzz8VZAg/uMGNVUcbgUriOuDM3JxUX/qQjxN9VrCMOyPM6yDaeAWUyWw4YSC
8HKYZOXw9RdjgsBWlYgj1ZL01pH+1Vq8EuHFuDB0DkjCo5WHiiWll9A5xO3z
Kn5PJgewPfofzWD80HPFZv/2VhBdG6b9FxHVMG5Pd0QYq+rT3QNC1gkbKlO9
D/lI9XilSO9IGDdKSJIXjXxxc9OIzLnvD9sQS6QKpulyiemxqbZqPWULX/Vi
DUTIJBt9J4hkBqBPnbOWtHRBufIwni1SyusGmCKRVHHFZa5HiZ66PPYEEAXt
50dFYqeCXOuJIufA4RUwViR3VqwUrGStuABhPe/YqktGqof2RUlPUkc2XI0U
fo0bIA7rlSoqZDOQVIu9L/uPEgk1FjOcS8IArunUyMeh5Fv+3ZEoFPs/zVZQ
utYNhHF/ioIaiSPIwCSGu+TX38tnArv7a79KsnR60qjPKYhJcLNM/8ttMHAy
GEhksUU3UnllCxt1MKHXG6YMfP0wz3JU67FRvtHsuIcpLKqwC1YYy13/EKmR
CepeG1duWcuaH1N10ZX+CFHajwOfLeRnJiM2sXJd+gZsK6wEPcwRf6UepgKU
PQsBCQSXTKasdr8ulAFKtOl3RjfWh1UTF3IKcELJsqCqv3MBXq4F7MC75Jcl
ojvU9h8v9bsbt0ztZ45TjbCf2u9EI83LxvqE6dRc20K/B68YqlfEd+XMwAuO
AA1kTBOVAl+TIK5+5KqqRomxU3K6Kfwo486kME32l3lAVdwLOF/W118PQ47E
ZB+yiJEwt4aWHFnAXMOU8uUzUqPmWHTD2ZEGH1CntB71JDzzv34yKN0jALgK
pnlZX4kFExuLtXawphJnTsv3ePeC4881SzK+4/KLc9dbHjK9o5fG/tjSdPwQ
o+FA0DHzoSHgq2j0LCfV5k4146UF7ZGxMVhYjJoEGpJbGnzW+fUo+Omu5/y/
4mrNp1HQBEwADNHg+7yCr1d8oLsRD7KJXOAFKMnOPtwCH2HUcsTxmIeuSUBN
XaghcFkjmtwQA7o8bnNA+LI0QHQ+0OIdGuy5Lw0iuCQCixXCrDci1Ou4GsJ3
wzxhFmKZa7NsnBEwR0bkUzlK7S0kcnkNX3met7oeBUDqnOSJNh0fkTEwGvdw
fLuRArljCSrv+gPb5rxc38+dVbpMPD7LR3yp9V+RKuKQfn/wUGU6sPeUhu9g
Q6aZZ051CSI0cern/q0Nx5L9CO/9amtSLlyhRquf5GBaOvRndtVH4UCL80lM
3SSdVai0oMLxExwb7nmZRMDKYx4h5uCybOSruV7dirOo+X57DtwFx56skLBB
ht4G0wues/hUMNcoZFMO3Uzn06w0ZvlnqwZ4y8E3dhCKgzvCvrXBagUVw5Ck
PWxft3RvzL71+EL6PFHzrOLmZNZh4ZszBo0HHVxUr1vGtKFpZA9OOeoE/ARn
n1NbsouZM4MeRMS9v7VUDy0fzZdfvx6T8TVCMdAQBipGHFSb3LWK/Y+KNerk
LfZmtKDhVP8diBoCsUsM3o9rzIXsatvTdCa2OldNSpatl/1x9Ub6BTvexmyz
SBIUSCU67hWNQ8A8wf6u1aW0qJOLFVHHwmxbZ1IGR1md4EHyU/9t+XroVVj5
H7772jR9/f10berf6GbxktoFQOyr6j/vevBKuHqHu9TeXhbP4zmiXe+2TfEQ
zDJEx1cCDb6yhmyX6aJJrVmiHA2ZFvTIKECN+CoJh7N3QXqghFEzk9G2Flkh
N/B0PeafJ0moY5r698CNQLoUk44/aVkdBG2heJ0v8ExV7K/M6v28U+/W/JwD
bSQvT/T1s23yQ75kSNC/QAeb8wkKUDHjarKW3NggQVmNL5m3qf9otFa/JZMc
/Kqmv9h5KWdZyrkc4OihVAumklgCRLFGgQVbmJrQ7lgU45kEGB+MC69Ute1u
QdqCZBzAeXMMHpGqvEIS10bkZtB/eRbcW8JPe4WPGx3oD4LhK+8e43T188rm
MUl97bIRx/RXPsykozuwXgLcEZrHpBwz0Onqc+/VBkgwKq5l9S5aQw7hEwI/
leIP4jtVvWyx1YIpZWd+1h0HOydx/odpWHrWU7jLFoX4RllQYHyZ2x05H3da
lVboACUC+Wd1ufwHmGrNcvAltZRCbLi+gzWxY3NATQmI4kWCwL+0Ejjt7JRK
8q1FuNzhZDHPs1c5agYLSVZvFZbhdk+xp5LKKW1RGj4Ul9R+f0Y8iXHTPlO4
D9K1DwURdCNPknh0IvKbDk1avqMUzUYzgsIBLVt/Wg8V5pluztesGSWLjtQ3
GJJUmuE0UZXJcDUFts1hKH1n1EfftxY93s0S+eMYkPHLnzkPAeM7v+kf48f9
jJWEe3d2TKgiuKeA5wamEcO6KxilZnmpIYaeSh1mUxHS9To/YbS4x5xK0axc
pIlg5SzA6n5detsqNpPX6VmPN5fKuicMp8a9Kf8l0VLZ59hAC4ai2qrzR8fR
CRdva3kdU80/3O1qwGSltygCiOiyPhRcwEK7DzhW1+z8jDOlRaYaeSAh5IUn
nqS7b+E4opKdu5PTAWwKxJ/bSdRHZCgSNcz26rtk6OxNdlTkTanqQrAxgDvl
y0c3Robdw39CXFnT+VdxDkIDSYPGCY2FvbCgnZ/9oVMXdYJzbHl8x3yoc0K1
JC9plU8/M2euBbRLVpeCZ3r8GYE8lKwNYfzszYBzOrCME4SgJ52jQlAWEwbE
YH0LsN/S7LE8lirOpFMkxtaFmv9IXoLy05XFX04XJdAYunPX0+RCfJPNxLA/
F5tkHIWpVHCwkEhBdCxo3eKcvX4dpHjVItEr8m/yroUJ2sBLoF+SF/+bc89E
hYUiclz7Rd7U7ayIU4Ge1335I/loh/VggUkiwelkmwAPl9lZujljp2KM8cpL
RzSNkNGopSZSiU0cJ1MRHJxWk961mpYmABUEE1HkFLrmI6+AvGsDvDu8Fjna
aVQrkKpnf9TWLVGE+/tw/h5AX885yimNMW1/i2DCyGj2IuZcVjI8h/VEnH/p
VPMg6p0lko2ptqjegr6np1/HJNkL8Ie3Wqf+QgvZx6pq1Dd4tGDx5xcgn0SL
H3/Wp8YgZsd/bbWf1xlHUoB8/yTWVRr6qeYgQingd2TH1ffunZ/a69bWywrE
2xDz+1vi+N9CGY/deU+ZQCf+SpLe1iMdRks8NYXAgeFP00Si/Cf1x+AX5G0h
0jFT2BDRpJ+XatmJhshU9CCJtbwT4cSEKA7uAwU+NHe5yRarMeRJ0u9CTElS
4wJitYudHahGZYV7gfIMOTOOM0pzi+DNTvSDFt/kUoDjFPx2RMMjlUOr9vxo
V2ibN42SNM/60onqEPFwyAggGPTqaLNtH4rfKlWk4WKEY8UZpe+nAJaCNK+g
jazSXQE6tPAK8Cr4XuEo480+NFzBBTze3cliwizOl4WJudi5c6aw6Ht+ApRe
pxR9uwdPcPoipDkJejnc7TfPi5AvtXRyu89swOOvTf6YkQDv0CS3F2WGmY1m
8771ouIne9bg60o0a87JJDhTkcdv1lSWCwVSQh0S2C73tOGLOKf7qypwHWox
51u0gJwiieCYBC8UXuqI952pKkzpgw3S8kwV/TWyIO/+CZjNLBJB1ivMU7uw
yXeoHsCH8ZnT/9Tvht70BbtJjVNOECfiolm4TdF9fpDXpt+mqEiJ7vbJWLKr
ZDOPV5qSLDTgKjkfRhdO4BaQQCgzAff8/8T62TT4qI2WPbmOgtML4zhD+wxL
yHACFwVPnej3cCCemmdobe8eQa9poUw/G7ak5E7f76x8dnViwpzs9gYIkdyM
R8YzPmG8mRteTanRyKaHdzGMuDrFUPMxsdNHuknx/rtd+0hZfM/cmFxyovkr
78xxZPSaJQz3jtIhlXeHtZiUHmWGGFnduavIYCdJ5OWjASlFaVCmBTHp10sm
ACd9KpOhuNsIOcyQTuWuoyGdcpMYcZfKqMeS77bmGDsl/epCuhVbXXXFMqmO
LN+AgWwb8Z8tB808O5DDuBpeISBIkyxLfqUStqHSXgb8qhYbCvSiMTh2J3ra
6/h4IbG2rozgDnt0kgvDbqbhXnMP4DfnO9LnkksxAWkG/n+ZvzjaA6Lj1Gwk
EsHq+I4VBB1dED9+Tt4HW4fkp4TgyhEZpHioL0OZ5GuZOTX7vFcf/pnsLuC9
aIvu1OzzSAGPLt/LQ0T5DWrWBbLkURWCV69KHHxxG3aX9X/nhKrJkpetQm4P
TpnGjw7FoLYqqzW4rMVh7kC7lsiqRwpuvbK7rUNg2T3UiU4yjFEXN46uyTKJ
1P6o1yktHxFlAB7GT/srmfLY/JNYw7KwC4LutNxk5BUIVRIXv4LIROcN19cE
b60pH2toOhdZj7cVVeWn7iyUS3cE/OWLOyvvH+iXkmmK3km5QwBWG2ttx7X5
DbbEjIsr6R6UtltxJehCT3cajMLQs8SH0Cth9jd8k17I675xYhStKfSmqFiJ
lJxkTJ1BQWTMxv+nZF6AhsiGKShDeYduc+HRoIGuo8KRimODwcQI63ogRwdw
mJ9C4NzjPr9z3zmd+Pn23ofgFfXLNcthMgz71hYVl66YvFdLroUJ3K2JPkk/
3gZyDM8v05a8fb0LZ2rbu8t4JAwgFEil5ShjuIJsbCTWFTN7ePwxRaAI16wP
+m2UHd+qaDYC3tpTUw/y5m7kotAzIav86bCtqxofxoT09x0iQ1KCPKlNDpWv
KdPosvSfSKG8p5msa7beXmmKMsgDNpu5rLTF1OWVumR+scRWffNuxp4oX/tY
+CYA0JgI7cJrVHxgvB64v9uWI5WueE3DfgOLtHB0Ytt3fJ8l4COWWrRtiK8C
syJ+6Kmlgoz6ncPvePqwLWDNtldD50Z5HMVivQxAjRlIfGd8Exsh4COYhTTD
qXyLxvPWB20kEsCLAJIt3NGXXFOXwteU8BPVyG4rIfaRV3FxHJjh4xPAVd5A
sL/8hjHKMhIYaJbyE7pOzzfGx2m3YV00/wwfVDxvqxfcXL9jyov6wT/5bSC6
L7G5Wq9EAUvJVAFigVdt781cDv/XDX6IcijGSVJANadeQ8ykw7yP9V9bV4xY
qBOAQ/oR/yfsnT1+0EMOWYDj0+mbCmYcG7PO4+XHe2TR/wPhZ8+v2ZXHzv1r
dAiB8Bfm6hc8yCLMhoWZoljhKPf+dqyX02kV0x1/pD+AzuxdQGDo30sAZpHt
FmH/Mi+xHBvGAUMSXr2q86S+TNAocVUxbUMhS6uAyD6kdaWILegzWe74zVqf
UwUNtjU/ST7HPgLHGjXEEi146q+NmB6koR86lv8IUhYZOWESRjhr+cWDNhlO
lYqg585rkMkWbdY8+Cn9oYM8GClFyGeBTD7xRZe7/HDcamwQRJwnmDrQjjDl
I/4wK/Iy9PtwGB+FVxHZjo44F+YPxSfm4yldDaHL8HzRXFDC1tLgDuKU4t//
WDYAFJ8VjvRMQqBKNFMbEttULj5sAOFrqyUQ+LViYHVKtK6sPkfiR/1j31mD
Ky2jkwhaujWA99VsYKKZn4+hlETjQTqFqU07NAivgel+WupAxVPzA0JyoSEj
QkRwmYaFzzdYg8ZEX1v1IhbORt5anBbcVMxmnVSG6OVkJctwYi5cEDtWG1k/
Ht51wGrXaxhtUKwxN4CllKU/6fBO9tTDO6LIdUu3WMr95XGPb6ohp4nXOe6d
XchiboAkXmsnQqQSE8yVAK/bxcO5n4QKZEIYKxAAz42ao100/wcK6dzUA0Ap
REvnth3GOZ/wu2pgPYN3SUGgDkg3q4uUQPIyChDPOd2emk0kUBQEMT57KaAW
ubVeM/RZ6rTTPv85dV9uNiUndTYeZtyqTULIUTRXyIdE8mkoOxRRTHKJmquD
RoQE3jknkXgMzjjP7WWtZ+QhSwo96v43QDm1iUEJEjWT0+L6n7WUgPJ4BYVl
da/6b0b5FleDPDARwJSkT14LDnEa0wINkoEYNTGRoOdhrK6l5Mll1Dcm0d5j
xorQGh/+l7YB6k9sBRQlsMM2dr4WXwSll2Lg/hOOuRNN3Kw9LCKWmNYXigxe
a07cK/JvMNYYh/kv/oXLte+B2MX7pR3oeADByIQyu6JKcVJ9282Eyc/t4WCV
4UQ+vajp5muxE+V4MTSVKhJ7hr7X3r0bWNuP2lqaEW8863WsfZwR/BQ1Qu+O
hbiaSYbo3J4xAStuxaYRPlpyBFLxVhk0vbkCTtP6vGaNxtWm7uw9gHCQiqWV
vbW8IjmUp1Gq57ubxHv2L/BLIYoX8KRq9snirG+wzCE8Gkn+AuGo1gX/Gayv
BlyEM9QXY7fxvQHSdaID0yFrzr3iEZvfegXER2Gbf/WtqWBuIFj/VzQYIWNe
j5UhQWgRkeAu6AN/yxpz69bG2jW2d2DJe0vHwdZ9aZjwOZnmZanBaPI0Z4Qt
1JUnUymlg/yg6PK4ZdICdm57Y6hC5fBRNYaO3V835efQuusIGRsPL2oQM2Oh
8LFza1NS5AWsv6RKRhreZbgIE0a6U/jMOK5ukgKoJ3wh7Erdvixbe03JYgPh
qUyug9z+0xl/UjtmZbNCRhKbrsrCe8Hd4DFIVbWXLVvV8CEB4FNw5slCABfo
BQGs9Q2Xb8FrOxvFYEF79Brvammhi7tB1Q5+Tfp1ARSn7xYb6xgA30apSzFi
tVZyMGzShk0G8KIrs1AZCb3wNg6GAOIT0rYPrySNG4efd0L2wcMmqXMmsi16
tD1TyzgXYZ/KG1ItPFrQy//P1IMVSivu+JWlAr1FrAqO+M43iaQY9HN9KB/a
9YQ8+6L+UWMEFhInfFEA0EIFzGey4wDQOBSvsKTuHVtHMHMy4qO7ra7/nsQ/
0+jnInD0mGfAJwLMaSF4J3mSoQrO/ruWlXLU/mRfzeMXPdZjFXR1SxHeRoh5
pINxNrWl0wqvo8UR0y6QWjlQDimrCAPTlWsnAJAmfVJqYu5p5DeTLnR92Uci
1cBwDMkGSRgpdRSywUfDoM3WFePJLwYIcE+lWAykVf3uuVJf1pvRc2qhKC5o
Z1baeb/AqbRWNh5IvxSZazCqELx1IofSBf9Iq4I09zjflnd3yR1O1NuZULJk
KGJ3tA8RySHQ1QiqvEQ5bxY7UZFhNlTs3IdhkWf3ZasT2u7i8uUAw3ldJ84V
laS5zxM9bdZGWyih64rERu3XaVxf18WIXbik7trFXeP0wMus/oQ/2aB85gir
c93+ciRUCxq/69TCqpS8AenGHF8cmcn1vmecDBDA33gjxbrnRZAdNsSN/3sI
wNSt64Gqh69Jd1iexMHQvyGIdfWyXIEppc3gX9q4h2pYdAk5VRYLfeGnN8a5
zruyPS8nqnVjBaVY4NxJUY48UFRC3DqWYLAGEghvu1JOd7ICsIRBNo5rC7Sn
Px6CxwFk4d0zP2b+CfogjCnZOQ08X5rK6QEy9VM7vhSU9+VQ/j3n4m+xZb7n
CyszQ7R8MVPXMF6B1A2vwId5U6scEIwzM36iMvt0Gm+ioVRFaXm+DJlElqKa
/CmHphzbbW4wVoxPIS05twOyedIIBvRwwsP4zR7nyKcnVboLOxOyLlMq8Tu6
B3m5YgQCUY+mNubTOiSMw+3/FaUJ5MhCpg4MCJD7TNtUoB1+xRofgDqdhoK+
X/zJ7m4aHzutHL5OSUHLUwphxbb/mh539u8VmWEFpIynt5mdOA0GwMbdpDJM
McrrU5udDvHdUABuCU1YpPpoPnac3ZCakz2db/x9LpWPj/LdsYppI2nVUsbD
59OBUyADS2jCt3sSem2R3YQY14jB6UiCSpuk2NF9QSmRGUw+fdkFGjgfcW/X
bRwaoYcJEh4XI6fcREajGyQ438HCuvGaR1DfoQSZpF1sAMFL1Iimd6n/K2m0
9WtcNgjGtb70WkCiErheQd/H8++NRYFsBMPu39QNfhrm/zMQHqqjp1+5Iqna
EDzqAjLRX1fKo72nLy8wFJfk6gzAvZedGheNWeb2KZ1sLKi4815Y5JYLXQLs
T3G0/IZWFWVPDYhwQtPESzyneznFy3iVgpiM2Ya5BBi1lYFnT6ZGlXm/F4uS
ONDSug0DH8/J+MXiiqhqSY9WNR6ZbusJKLqBRPunurnD2WO6KOw9rSUmGejA
+5TCOiNS6gAqpNB0TliwGxdauYQUHiHu69tjeL3CRdGmmWvgjGFTBVOk+BsG
9UMtZD2bbJboWNQQaQevRwCwyzYs/M0qFXYjSpncl/2WLfk9XfAbOZv99u9e
viyvY7EZHjCTrRxjvgNjOEoBLdCHZAn1WnMFB5T+KyIHES0MFKo0kccq8KEx
EK8nwdSg34dBnaoK5+dX5DCXsLdq0O5gWM00yxeawkRNXGTq9dTjoAhNZjc3
z0OO5udYxZcE2t7n5zjmLKwAFMW5nKnNCBJu85+Ii3nGLd5D/wY/IcKdkgjk
QYdob8/ohUhmF0rNDXEKW38ehTWiiMnBfaOJuQ4mWa7upVR9Hgj8NGMH4PgT
qwZ9eLM7pJnUOGjUfAks7za0hJffPsG+Bs/9bFc23SwCO9wjqSGgV9S+o/aC
/8x2xxdqo/Jy649dfBFwDcKsEXqfgEb71DUZYC8Ch3U/akArpTD9SVn//jPW
ujTOwH9ZzO8b8TeUkCsKQp2GPccQ+l1SEizhY85jliQCUsn9PsvbVvlTcUV7
DF5BBloDkOBYJmxpCLTFd03vUQLGp419/n0jNYjJYRhf8I5KS9t7qu8kLUDX
mHlL0wLGrirzGGVksKlPYSRr/oVtjbgrksF10AAq8gWD1aIr7l0KC+XjDLEN
7zZA1pg1m6g2RagSDKQouimU+3n5NjXi3EsR7aHoocF6rpHSvVE1MBqqUBYU
fROoS3zU4HIJKWZvCQMFh95BWAO/OS2Akk13biG9qYh+0gL/osDrb5mxkH0E
BVANyVtMY8Mf5a1lqYy7nYXgN1W802+/qX64q/FTHu8p4Xxxd21hCjLOcIbB
a+1GLs+zgTThIDpO4Mj8Dyw0IQx16fo048ifkXhu6pm3MSfMn+NgWERwMzK/
x+IX9F3ghKKqSEZ0SxG6vMb1P29v24nk/L/+BEd0blxhSXaUmatcnrnYhjcc
FmThPpTzxupWePNi+OZjZ2/loYJ0Yn3kzmglCPKMAKpwKH9rlonn50hNH+Cr
HarF8HueW7DA7ndU03aUSwO68rqbj9bTL3UEvblra9Io2Jq9IM/gFENb+MAT
QVQPE5QcMpxqd76y2dYvlNTO4G3esg8jwijqeTCCwX1eSIR8tMCQrrlHWWWt
Rkdm7tCV2l2lL5z1an7Kr728okZFfxs1EVtpZhqwbjZUZKSEw4mg0D+qrnUO
3dCwuhvc4MnanAVlEwQMnry5TZ+311fU/fRjDL2NjO1S7CNLA+4Atrkvn1vm
d6TkrcCUbcgnujyvC35+aCWzLTvlpUFMwY+Gs8nuGkB658H3/kbcV0aXHlal
KnIGVy4a2P86NieFJaV9e6jpdjwMW8C1X+r1e2rXJptY4H7VH5jZkFtrEbRK
oPu4cyiKC7dWulL7GEH1znchkW8tkvjkwPJg1+i6pWEr83jBEtmoplcHvXQA
qJ3Qf7IHJ/IybN/SBq+ELKEOmms+WLIbFY0d/OroFZunNEsQ6ighskSSMyIY
3spmm6q7bi5f5JO4LmBuYApb6EjAZ9aUtVSOoczSPuVzfHJFRU+09bebirBn
U3Gxh+EBUx0LBS6YHbepWeRjtcG3m9UFm8vQDSpWypVJM2RmjYky1Bbq455d
8DCLvChKDUMDlDjuYkWZKp/nIGCZnGAE/5kOyX9mz1BY/cf/QoDuUQ582+f6
6SDT8DygeIVS9ySmhKkNIl7KVfwg1mxO0cxyD6Bguqom9w0I8ukXSIrDfQED
dHWc64fhpgDEjvAiY8kfB7jJ21Zn6Ce7JAOJwGiZ6OqH/Dl7gNAfOF404TH+
MwzdkK6sLVWXDXUMumeghTfnpiwqJTCN5sRq2X9Perrus8bOLSIVJqtwzomj
3tUqLLdbc76QZ9JJaijTf+r/xlM9LoRolg6408Bk1tpwuzyQX+j0f1Qq/DEN
PQbmAqvA0hGZsnPP13h27Hl++D5gIagoVGDLNWYcMq+uRDa3FHT+SV63qNWt
FxJ5bP/+TVzj6v2dr1bXDrsGRr14jCOiOwKdYuU49Hhva8LoSU7WNvbSZP4v
zWtfhzzrPqTvBYMkQSN68R0tUzmkY5kDWgyRy7CKWN6nVY0+jF0Ywpf4hbab
rHPmhooYD8AHeu/KOu/ixocsb6R9Lyu76WW1L4jEird3rUVGI0of7SFsIgAi
zx/yDAu8qBrQyBhmWlLM/Vbz+50e6LAjiBZxqE+rmZuB8ibUKpGOvhnlODGK
+BsPoZQYfAO2Zu99X9S3HoisSY8x9vjfYByjEFJEv99/+IPNdtr2O6d7XUxl
+3/yt1GBRiAEPJ+sjz4+yA7JQOKBA32+V5aLwPxJN1iMpWdRleH+JPn44HlR
PshfBTbNWcdmaqdcrc1N/Nl7yG20Jj9Da3l9fbpl9G2w6kGqiuSfJWvvyXG8
gnQRe5uPHTNwAhekVwiEgnWjPl/3LrrgflPt/UTPc9s4Xcy7RYTFu8/MWyln
bjE/aP4SfvxTi11W5ndm4NWspY0NPCTAQVGi+frfA5FWuIIXFebrztJOHYWP
mWtRUrv2b/NMktdVzcuQKVcL4R8nH7SZ0Nce3egbAz/K/RzKtOBjo/87MGWa
18r2r6oQvbxAG8VGR/iBapEMKynC7gyeJuaC2v+im7kgST4rnA55g0IX76H5
BWSkWwEx0W7dQ4ScKMepghXEawq0jiF5Yf2XibnJmoEjrArXQUnfC2AIh81Y
AHcUpRTgg7tbVfpm0wkt8fhUic+finkdyWB+c/UVVKuchqsCrGUH4qmTe/xF
UCfWMjAWggD10hJKIkcaJmN4tA5PfqDp5cRcHRMsZz4tx+2zBnP+QdIuiaAK
c2L9Q/IAboB83DsAazy8CYuY770qhWGz5fpO7rJCgZ9+kdwwfd1mOdhBRLA1
KvG2X8MdXONESzWZdZrp/HEWwuCQ+UEfqYlIjST78n5j7/znDS0WcJfW9mAv
dTjiucxK+ufAOAFyZjk/mybIkbnwyStgqOjsjqowSlj4CWleQV6pS7Bhcj7k
exSeeGOLEyty04ixUgv0pTmA1wvkek8nku2O/uZWCy4aC1rhP4OiyUPRM8Dy
WG+d4VDjGa2Qfohsg4wkvflauNt/8tzGqh+F4hcj3+A/Nx9/zVx5cyl4dZbK
yrDepk9MQySwmMW5vUEmh+uqlnOLF9BMV3KyHyERqKP+mViBmWlBoRrzvchv
yPqBX0Q7XzZv2CbeCqDW7WfjMb23lbcsq1R2wbLdQIByqNTuLJtJijXG6Gv3
tJqNOhHmJlsHKa0ufB9m5yC0RU5Z51SoZfAB9WniDRfsw6f8XIfM8OqykyPa
dOWoFib5zGGGkXRJEhPtdGTGh46Qm91EQHzmODBut9nSDgBqENypiJ01chjc
OugLBbZJNetzBxLAYfGi4sQLiJPdWxNy0IZ7WUM1YakJlZdOdtD/PhcrCfB2
JNIKdBO1zLJ5XbzNFJMQXQBx+95m/Kgyci2ENrTiANDZBUuQJAD/gM9synFQ
60LwxyQJr5RWs+pi5Xxf3aHiZxM5CI3q0Gi8Hx8PXnqS/YYMVAKf4pvxE+H2
EzkjTbXJ0MKn1dsnmGhVCZRcK7WDrQTIta9IOg5x1ib5VDHDBHhFJxFQg3AV
cpukaDPRJHtA3yCDFc6nbkcLmfUqL/VxBxx4tZ0K94el5+QEnWLDxBXR6pED
RESrOXLmwD3Oy1dWelmTcAVLy0McRlT08Rq9eqPXaiOEhmE2+Rv0D7JGBt3n
QFtqzNOpY44xaedvIpiuijD3QXV+jqYGtjZgJ/wMiCHlATFbNEWuESaZ0zzA
dMf8ILmMEf8WRri00pf2NtB7IEo+UQUC282d4dY5l4XRxvXoGXe/1kYKCajY
/MDOkVJpBfF6AvS91IWuom96BjpJ1t+BIT7UJuk9ry+OKVrGYR+NXHz1xE1G
uEIbcCRDjrLWIQfVV8RekZ+TAz3E4C2fncZ4b2IYWdPHiAUM/Bj33KtXYgW0
qOunpfy/NWMJ1VZrXPwwwRJI9leZ+AwSwH9c5WHeel0MI783x0+l8awAtt9t
WvGfxRP9Zm5W0knbHqoFMk9fTn71j3RqBUdK//dMdDufhnc3i0/cdW9vr3cv
JBGI6AmhbEqfQ4Lmx85KTdJ5cQd2dgh53cQayJRz3Ccm86xu32ayBuuPzSfC
xrbpY/rUIX87fnEM+ajqrKE5/3E3GJSjwopw1hVFOd0Zn0TedhEBMRXXg3Bf
5MWYlK/CEt6OsM0yAzGt5SSEgzPcNWydLVXfKp79XtFrTMvEKAPmsb50FZu1
GxgFRYtty4pG+zF5qIfwzNtxI4TqVKBVkPnQ8Nm70xnBgaj7TL6Yu4T8yKa5
0aXyNsIjtdwWhxxxSOfrxH+dttPjLrn26r2NOOof9ZrZ50IaXFXTnV1MJ1Xp
bZu+m5FyC11x9WRemJWDn178zT2pKsdc2BdO6OKeRWkGO+AR7jdu0xww67TR
+s6p90o8teaW1jPdInRInd4WYmMTapeHPYaLzaPlzBd4kLHc8K7U80JRt3Ql
ySJS5JJH2dtpSLqYlNazF42HTPa5LTQ1SwKn0yfUC5Rb1yVpYBEXkVT51ZKj
gVxeGu0IjrtaMUfYg5jMEXJenu8rmHQzCwoly7Rz/vjLsYYqT8kUpZH8F9jl
x+yBUNssJJOKqRFRx/9Uk2u+Pw36/kWzTqGTjaUZaqSHCTmDQlewRewKak2S
x6WXIJHDUv5oNwv+gROEePZ8ykzxNpAFWsgFl2j2weDtkoKDP0ourOyY34mG
H34hH+ot7U+xTqN9Pr1imhhJ1W9aoNgTx7hJOMx4I3rtL9HfCvUwgBqsA1xA
Ixg/5bWFn9jXo1zutBQZLi/ehSkBfM5qtlTGkSt17REYSwzBLdd+a8PBN2of
1R5BKZP6qtFDPELlgMZNT/aZxsj85rxYG8lQvrkGBPjdnKdd31iS3CVw0941
0XYylxCQvNoaVPMrtBxhLbQ9pX9zy4m4Orc2IZWOuSDqRRtYpfkaE/XAG1gT
Pfs9lPFFIL8QFLbOJfFg9t9WynnaBONjIqKFSVMyC6K4itFR/IYzj/hrBaTw
KH08N5Sq6G1wWBgsOwNICI7zAr+smfWBcGd264pp+dkDDqf6mwKTCdTx5blp
/I0N40SjSdiNoCYJ14T9t3FoiET13sMtf3/50RYkMEkwaVEaaFxrFA/i37zL
IPH40GtqBtM3xB4Gs34EUw1QL7CnMR0KprcpF2jRaijEyPUmjRxr41NtKzGt
5ShXNn7PFKCRragfB4fdT+ixTAf4w3Bd3NDULRYnsilB0tIyZIM8H1AHtdyd
LUIcX2YhqbUtJ1KleUgO7P/qfvpX6MRgwrGW/1F97IuiMInPhQ1PG4GsIcxb
Ordu9mIw38RH8gmmdyYOM4AkGR+TEbvW3JsUxsP6T2SpE9dTKWUbytXDo/1i
YyTeDb5s+enFcWEMFqiEZhQwl4NWSPn2tuc9egaWYYT+3rDaCyLlEK4q7pAH
jXK2f3VD2WTP3L95Vkzb5zVEFRWXbXddXZCQq7zYkI7TEtXWj4RNpZl37e8S
Hqgj9LV9CHkMO0CfqHGRGuIWlj6HqR/z2CYjN6Z4qaNNmed5lyKE6cBmZedD
x4K79HD8ffKZflC8HmfrRR603n128IYsk0jxBin4p14ihmVxATzue+d1TLpx
aFC3r5yI/I3l1QWcoXXPvp+6C+659fRCB6c7hgLZMEAJ4JaX9fyiscF8Ps1U
ZD6JnM42q+nywsDSqe0TGrfiY30d6J/Cq3OaxZZtwYnplXgIAv/T11Fl3Piv
pQ4SPkGWluMT8yR+Q0JPdSStM5kvpIJ1IqY1ckPaRF7Pnk2ReyPfJZX1Td9+
iYyG3clh4qcQcCNk1f48cCMQ4O7clKfuZPwBDUCnpF6eas/hpx8q/rDV7gpW
zqE5Mt5k8sQLChnobRmRXrUGKj/bALREUGWX8jLPHocFkSc17RWyn9MOuufV
jUjbWnFUKQVYUhQ5MEO+0jPcL8dlolHeWDMdjI0jqvWZEZfoS+6R5uGaK77H
/9hP+CsSDmX52gtT+5PyJupmhz2SswOTitPZ9Q6kSqHebhcMzD/KDJWJvgQ8
OXVYi6uvRnYROpES8sDE9RhTNAI+BiCkc+kpJqXMYo9eDwV+KgAggQkvF7Fj
4I/rP6s5v8kKf13rHFcxUBNysJq8Oys5NSHYQfl1R7Anu4u7QHgTs6hI4icq
Ci7+/HBAg1Ryj0fWJI2GT7WLGzSQIzK0kj8JPfMzShCt42raqITw1Z2knqrg
u5WDPaJT9ZYDMk/tFEKJvIpfivsmzLV9wmujuBhW6+57RsmLQRxIWZCshD7g
jE+nUrg5KtRPI+z0q9Uale+PKzfmiuSfCZ4LpJEj5C7EA3abHZjhlXMWlr/e
ZGrwJOSWVN9+zsRqECIk7NwZd53aYvcF1MtA5AjpXCdrL6cDPvoGoO8XxgzO
0GsSdyCviMONaf8+T+R8m/pHiq/Ef93PPy0q4ucDsDm44UlMoh45UdNGJWLd
E/QG7brVsIOja553kU2LI01qQqmW/2et9J/izj/VWfgaUOTQCFeG9ZVSRMBZ
8gP2xpEoLgs9KDMiVBV9OX6lgWtCQi2AU9yZjhziME8dlErrB40U2wDixQ7I
nVQuflmiOMk0wJpOax63XiZTqbIlNwtrTPukXVsOwxBI8orz/3NQDiQ8TmWo
1SuGDM9q8tNPd6TpVaogEAXpUfKb6dQJUrzpbJGAkRs1JqkFxk6yvQum3gDg
zH5FoTdR2Y5mxO8Qh9iJw4Cm9ZAfe5a6HDYGl/ODPX/8ta1UJxOZDbkpvOxJ
Kd52+EWWlCLkGHCfLavLOK34O2jfz+yg/3NlDhrt2De+tn0a2I8Fnr4A+H4c
hEQUHdFNDdK92wpyuaxpGi/w4yRMxuMmb6m8tATP8Vemn4c4RKElUmP8X6OP
EKtGJSxEZgBlr0TCnS7a1Dl0eY5RC5AYLSw44K9uRmIM0Efpek2e3osBN57H
gGtA5zn6x9Ugdclg+udPuQGzGWpynBrI6Fudi3Gz1/TP8B+b8q8a46fgYWep
vBTdKW9mFsFdWkwWmu0D2mpjeGjzFp5a09bq9/Umha5FdqDhX1FMw2cCNCBu
KVJhnA86Y7AxYsLa7ZAwS7wTKSOPY6a3r+zpf4jgZ2Dt4/am/DxHgsQyFxgD
c/YYocMwTRnAbPL7cZ7z+nJDL0xg4L0/lC9VLvuo49PwU0AT/K7qGj3g+ZNk
6ix6Mi9qcqbBynlToOZwHXmzmHyoU5cqIk3SeQbehUusuUP01inhMtLxYkEX
S51gAb5lETY9ABq4Ls/yviagD22XwE9EpNLXjUYJACnykPdqvHyrpJDKBwGh
T2K3WAP865tuCUfhQxbzwt1JNr2S2LcpGoeTiWZ3K4v2aWDEwuNaqChATIDH
4PYncmZkI+3RKLUdDpVqZEf0LUiDmP6WgctYeTejTBQbvDvBi9l1My7PzYpv
rEAT6dB8Sf+wQM+GzRMyh4oI/KlYTNBce2o7I9new8XfQ1ptPWdkJMkzmy9e
/jKtpOWFsf2Mfrno/nOPePGMNhbPzwV6LDRozDtZ2GDpE1arx1PPJCWrXgkH
nupi/NBAg/LCe29wnO7QbzeZOoj5fTZX41z+r0/5UCXRywB49CZel43w3URi
lnwDld4ZnvR1oZHBDbT4wMHCMcT35Wz4XAxtiREc+1Ze38wsEgrKV5l7lvBG
qPRDIC8Xf4Ez72MtTJeGjWFqSz2M1iJWhOXYtXF4AsnfAiGdAdMU7Mvqt/Wk
MvDYWiV8q18LrcomwM9R+aBN3tChNfgagab23spe1xcDaauNdJPeQA6MPONI
mB26/tHi79yB0sWcDnFTLohY381dZng68/g9ITgMPcPAfCWVlHYsWQCqF9/Y
9KusA3ZZ1R+Zyl3jubuy5pqKTtvrPslJSs8CW5Rkz/R4+WFOwysuL3aQM2UE
QzC2++f3wC4cAxGaSFXBZNfEmK12JdmIOhUecX4ipR45UavpDXiWQC5voCji
sgoghLYPpeSGs545nN4Xs2vvw1FJMgrJEwec7e2z7B9pOYcVA8lghEwvUBBF
TlwMvPOzCDE1rb9bjOmYf/GZU+Bf4UgKvy1TRP5WfrcCtBqRehQdbLpN4HDF
RLWe23204F9O8jrXe5IC2NIANJ9ZIu+jdvrNbnyiGmJ9NoZ4c4clhmqt+SzX
WQquaihLNcGVgHlZgSxw7MoW33jOdqT5aIA/7hbo+SE9YWvsgI25oERs+m7d
8duLrrJiS/C2CyMThgCcXOf2KWQv0ohpv3IM8rrUUXIm0HEpJa5338/TMvPi
MtryLoKwOFKJRhrmbdThSDShvoVnm+0L0BrngA3Te4bdL+/m6V3J8yuxi+FJ
vCH1EabHA1phLL0M5SvhioTofxr1W9871hg0gvJvaE6X5wMK3yE7NZuFmzEQ
Ng8Z2EQc878ZxKxZiQTVrLSpJjg+WLhr0MEVlL2adaQJp7mdBsOdCrUvAuXX
7DBwdk/z67yHfU5OVGzDV9G4P2Zw6BVmuK4v5Dz9a6VHqPW2Vet2StBzlSiX
oUnGwXw6mF2S3jKGDN0exV7L+qjkpJg14ZBP5ydDYczcfReAz/gE7rAMDbOR
+p5h9Z2YczP+paniNUgKJTcbz7MT+xq4ZckOtFmKnkxQFKOxrsphvGjyZS6J
NwY9Notb+yc4QvAKtHaEevgoEfppcrDKEglc4AIorVE2yq70Ay5NsOgZ07bK
gcdI2NN+iOHCREQu7jIbyYSO9zJ02SuQ1bp+yaC46fSsfz7rKnb7qugVgx9W
KU8P59F8hMGMbaLDpcJr1ASXiNWMFAWalwKbgdrXwoTV+Jvlot2yLzN2D2LT
JS54S4f0x/wLAyscmTMB7IXejsdbJCoDqY2vYTxo8iDraZ0us+twe51KnEdz
OHy3UuIKc3T/XMhCwI5AnKf1FVAxPxLJ9GaHy3mVl7EjPbQgncZpPrSg/0Co
yczUj13/z+mV+ySqfdQlac3/7foeidwOQH3+JHJERAsBeDe+axzlRKNUkBy9
T2nKK5zhvvAXM74vRoQ3X2Qo0aNKsRNRMLK5kF3w7VXJbtpDNveqgvrJcZI3
B3FeMyDjGji0PJo3wfq/poVJCAuHImF5fqwR1wEe/urNpwOV8Zl/QtSZgBD+
1YncZGkfBiGU8C6pu0pWxeZau3DT3mswlHwoheIuz14Y3f2jxbVnMXDqotkJ
l2yUrYOrDFjY+2MO6dMS2vfLe2jOohu8XNIRCtfEDq2i7wQ3P0XzAnlDZO4n
C3NC8qu6KB6XQlNjFZ1YN7W02MRHuGWiRn4skWQnujrQZ4r8JcA85CSiCkju
JYjpRq6TbehfH+gwLnEacVX+sIK6hEsjIgDINRl6GbypnSeFhabv0wUP6rkf
pu7F1dGL/H8EPNYt2ZpfncjpRmW/CIAKEjumtVaXT8TrzDi7jy+TgihWdAMv
tQnXs8XzZhL45FkemJ0IM+Ib32d5EUuGLfJqDofdYhUL8YWRs9atKSgZQcxF
bQpZP7efFOnkLLCvZAI/nAdKqOiNZC1Rwsq8Exh4Z/8XDckeH/5tJM/Vbcq6
Nv8oI9iSzewBx91QOlk0MDSBgnHf++vEzc14wDLFB/9Kwb3LrJgh66YfEfF4
VplFLKLsVbxkNoTsUqsavYKasI7kG5P4WDgxpRxVYC7mGjiz7HpC4fZXB2We
3qrjs3orWFjDviZewhA1aagtwQvjR/Tq8uLcIPLHt5cy8P4q6Ef5TWpSuFD7
IMi54fpCoyMd2LCpowZEbAW2gHHNc8LUJtQ6qB7/U8CAxSBDzwHMOT4XaKqU
eGdkdqasskQpxKZEo9gRd1x3ylLStC7db/LBfxfZbmiiSmZCPKkIHIF7468l
AA1V4qU86z+PDeV4hpl60IbAAG9FeKGZ3tsgJsth4/2VRU/vky4DoxjWf6iU
+RVbTsJFVns9rZDW/stuXWcMe8hjmc1k90PvsslZoWP5cZKiZ7RIEz+CvA8b
pc8dMtWDVaGhWFGof2JSTNAsDrEIk4Qv2JEzdVGWYw4aPVicE5gv4UkVLPxr
07F40DbuOUfhuDR0DIGsqQEWX8K+sJZPE4pm0hNIQwzxCiKKWn/UA1WtoE0u
OniJaqotnstRdu/PlcsvW0Bl3pSG8YGKLaotNpXHoCCnQCPk57Bg5gkkwI93
iADaE9muTqN6iDezezEb6FJmFO4jGs0Vgz9Kzm34GUEMUEsHsBxdabL1XMYn
rkrHD/E6NQKpxDfBuAON3sLTSyRuq9n2c3XIDME3EmsYtiJ+KQbszwn3AJGr
b+bmhwVoYPS3UxxmA3lV6NR2HOhoiyRHeQz/0fDTVHtHaQAGaqf7LTrHfNA8
bMErh7Ipji+ffNXB6HdL5Fngddwp3QmYV76YPoJphAijjeLOVo9BDO9QKxbN
pozduyLjgaCaTC58SbYaH22iBZtztau7QE1LLU07nFNM8vQEFVtFY1WUoPlV
2EpcjhG7MvdC5tfSBOz3p5R/cybFUpMFMEBr+XDz2EXJLpI4KasHTdDHNTUu
qQPjpwXHXObdAhdwnzerlDT/UC4wASFFJNJR0uhBUcLBoi21H8Gwh2q5/nL+
kUcMwdnXH2UpulbAOuz7vWS5q4xeplBh1Jo6G3WYRM5OxBkj+asobmJOw4VI
SLi4ps02k9uklSmVy+1r0+PE/AKaZpOdBlcAaAad+DiJsOTT/9Mz+UmU74FD
aClMKuekWbNaBYARpk9Vj2Cej0A+J9M1AcuZDnfsjKZCAiny/mB7RE7xu/5e
St3V4hkbyS8CgJW+2LidNn1enVimdaUnhd/zAKBM2Ou9WvsEIaPyMcBMDz91
9qljfEt6FLcfnlOWquzP8lGt9dBknhSh3kS61bCo5LD6NP8xWCW8dMrUFzqX
66YU8bCfAjNxHV2Opv3yNL/9UPsirPqlrvQkM51tOHh70Z9U7FghW4soyRcT
zvASau8AjWoSmQ58IPK9u5PCnOZ1HXnMJ8FolQdqO5rD2T1ggnBk2FYijhWl
DQcwitylECF3zE+3u86e1+6wdUwgtID0Pd+2x/4JhEIFA2q/MBhUywFqOZVF
JnW5catHaUZ3E7kgZRcl9YVyOBs8Ee2XoxQG0T0X1L3qKEqNnDmNYZnyX2Rb
XxNORjdfXu1SNnIxJ/sqEsI2N/VbWkxH9xIZSSq8fTK3/X18aoTiaziGfPcV
tfJm7Gpsuion0hbenbzYKAQsykDeFAOytWI9oEhzugG+tH4qrRfk6hwYq5hf
ry8SBy3ytT6Ko51uPWmlIod9uN9N7N8jesAsGPynR1UjbXomYr8B6PM3/Lfl
jaMAN7yhEWARYkKC/QBUEwGqTvybbQ5wUfsTOOq0JhCnqhIPyrM3gS+uBQn7
5bRazyK5mVao7/cHmUEeiQnnAyfRmvx5FSgNRSJXtIRVKZ8t7wN3aMjOpatR
lMrAAkfT99384cTWjlX9V3BtRAfXA6325lB4pdSq6b3HQDv/v9zPB3zVwzUv
A4ayJ+PDs8wgvLWMi1iauqcAQBEYl3UtKPcn25ADr/e2o7GpBEuj5L2B6X13
vLeONCmcYgSH4H1fyLh5hNl1Njz1X4WDivT1PZUJsPkl+azEebtRohg+DtFJ
j7SUl9xrMYtXffUmyk0RkC0wQhJukSqAnH7wRUhXp8TxwT/0yWjvAIUuhHIR
wLtM170wOELBL5o8oKj7oMB8JG7On4Icxlb/bXXkHDurt5mAIiKBI6KvH3c5
VmsDeXP9XO7lBObJsjRXLl/XZ7xyyyznrDnG6GQ4U/Yq+pCmNOvUEsTRfj7q
uGgAxDJ6+4zWZnwm3BgFwO2IduDIaxS1XrKmjQT8vdpE8LqRsLAtuSOYrkj5
i7BsLQiUM+q/gZb1PtkZcz7RkDvz/IudXyWLyGD79QGnbKwl0+pqNsMIoKmJ
ACguOb0JOdNnX1Uozy/wYb+PrvQNcmR4gBxvxry1WjfPjsphKPAjytLTGoR0
DNAVa07m4l6h4b6RRhfw4mLx3RqEleUXt/rls9sRgeNuu7Ye7ovRZdN5A6VM
biPhsEenGSSWOJchdkpuJEhtv5MprUQIFo75HUZ1KNvKNeWMsogyVyD32HQY
NKwJXPa0xqbPRa6NzfMZU7R8fSd64vr/q1a6N4Q5tV26zi8S48ie5V6SaQOL
JcOn7yY/hCy2/zkPpyaiL8CwkeWlC0Pp4ReScxabU5VHMe5kwqOyJKSP6WNb
KOeaS/9Q7yIdKerF6J7DpX3x7uaj0Zo+JBKWIKjE2NOUt/He1TWIm5FDI2kE
gJPuupCCJv3G9zC25b/2bKLLrDnryDCcTBg1/yH02H1jSHsyq55SvLPK8p/3
Rt/HZYuF9cRD3asKASqkvT0pb+TBdxqxAJsHlfv3yaTVNuJm0FgFLdSVY09m
x6XPwlIO+Us1kPZmFh0x+dFVzVIot1PSrZuU5EwYsDFGwTZLp1e8nX1VmzsC
uMXvEnj8+cd4TrJe9l6YGTYzc3yhqucLF0g7oovjAnD3Yq5etQ5fOU1ooYVM
ZojcLXFGXtIy6rPcInQaEHGqDRjFAY++7PuPjKrhIrosajocRXO1YEW2H32+
5yDfRm2OKSmzFbQnFkDGrSYX6xSCV6COlOeUTBRRGsK9nWT4Kq2oqgC9TRE2
dVPOz0574k2s8i97SwgzIRC8rDqF4rpF3PEOFrbB8yVnLnGuObozB9dfmtgO
r7/VLlyZVUTya8WB7Bc7A9kcVdJUtQEKeQgLtIOe/MRUrGCNxccjDPIShGjw
Zhpp2pFbej2PPlGUT4VCSsiKW1ciFxTuoSw8ryDl5NNmfT2uPHIJSn7skvW4
fz7uFizaUcGXsIkYikwy64KXR6qqx8TW9aJREcM5FdHoK3jGm+4WjlHv8/53
NBo1c1Ii5qEwefzgEh4OY0l6M+q08+qO6nRKOFzoB/sbNxLNvFvlhQYT8zvi
3OoSOSBS2FND+c4FwqrbJigkboBdkWC8AsrnX/E/OGwQXdQBpO8frMMZ6pqz
gJ3upRKk9CPripJ6QGcoPBE2UYoQR4i+RrRCH4E+G82jzU53azjzuHVHWLUx
Y+on0KZrNuJK/Oc2Bmf9wVCNyU8iTknP1FPevVQdk0DSWR8YRsPvgEw8l3bE
6pynxLrP6ElL76WiYoEmrlcdqtdiv48eUnHdXCn/pZyI304fgHPIDZFQI716
52XdmzQHvrNcq6LR7KB2k4I495jZFyAmzZ2j+ftp+ae3qBtrzAFibFuaF2Vp
aviSy3Y9y1ehQOBCwj93xxFtfaRLmTSuwYrrOBv43EuebeAVn1oUCrWU55vh
wNCLKfzFL5bM3usTsm5B+CneuiQFDeGvxYkD6iEFaP07ZVSgGOxJFr7+nnhT
8yXTe1enLUltmOZRw9uo/zYs7BjFs66w6Xd7SJ9JjmZZNQFmuwwvJtW6/T5O
E+3uEHC3nhLvZaAWclagvicnPKwnyGnVOkrNpcn77LrTpU7tTWxqoz6mg2QU
7PWkfe1QFLSdkYwu5KCRVXZc+V6AEUGhehG9MRI/XymbMS877yGN8vAwH1YF
XFttZCB5s9n0sF/gOobmSg3wdciGf/+hOBxD6tmLT6utrw2g0dgy51a/qg1s
rz0a8D2mAz5cT4lBCav9pmmQn0s8XrwUuo95aoWpS3ovb4+fR0tegNwZ9A+g
a9Wm2T4u8TENErqHj2ONdySj7Mk8Gncm4o3htl/74HoAF4Pmz2T6E/aFJepy
4CL9em3hplwrP4tDOwR+M8WIxgBmJalKxQvP4yEBlhKxgAB0mnGa8tHDauCA
xQCXHcBbEoXfQKyFBwoHhdz3gEGiRWjwNFLtBwTuYl22HzPDRJoro0AhMjsK
X20wOu7bLoNWlkNPcTCzzZUawvZJlCz+TOrS4jcnGWmG4GL0AbOY4q9MdXq9
I5vTJRfSlnfalTSCLxPT2RrILk2gE+ZFDMfAkfyx0IZfHEyoBbKdUivhhZj9
4jgGkqlNyn6oyEpgffwhIlCYz9KDgRZ0uDSjBM2fZC1jtENBky6tCKm9VCwY
KhC+Qjx9EyHU4jIPYy/eSYl8ZzWIqDfzi7vOB7pBqtAMqAKQGAY7j9kUKo9D
zjgK2fucZIIINLepTMQ+oL7ecoEIdSKg7PopB3mOb00gOQll9e0VCJoW7Dae
0xSOJVT6N1arRDRp+U70nxG0iDHLQbsyYopMfmXkS/OJjodS6ufCt5RRUstg
+Tppg/2ZbgoRRDym0z1OK5nuoNKqG2ktHGFP7LVss3NpD1Ccj8EHi7mKoCBB
hCRTOgyaO3X5MW7cgGJIkWNzvElx4gpbjCoH6SGI9ONGabF4tlefQdqfj+7z
YEpcy8wUqvWaFTFTpm6FR9TnKto6r325Z9OYOIXpl3xKfZX7/rwRlF2qM3lB
2ooDaUqQip3tU6CZn0HX5RocplkrBmSjgrauo6JJrHStac2BtJIz2Gz54G4O
F35uRA013Nl8AJa1IYoBk936IRKjQarKbLwX4uvxd7NVKpwEN5HyIyB9tleE
hjThm67NM8wa0/ikw20WJ7EM51jKdyFj/ALoKnv0Q8WKzCmUuYgUlYp5WNnB
dcSs88WcenYaxFvv9lkwM2LeTXGrAWLvNL5YTDFMQ5ri7gzwlTNPvob49XTm
/2GtLpGZfpMwoImSjnDQANnvZK9zxNTZbNprylg5eAD4AzslneHulcX+SC46
GICF4LjSbmY3Q8xgac2oNaCQNC9WiDFTuzADq+y5QvwgYM1b46TYyf78UQaY
mXqwBN3ZydPayIMF27C4M0dzY/azHaMo3TRhQiLf4KtpEUh52G4o5k3bI7qb
mPNnpFZkqowHKx3KDyxWD7ozu7KvNPWQsM+StUIqhWfmCbspcMyl/0Tw3LQc
/b2r+92w8csti4RzoHJOBRPAw5viPwLtDpYwIk+k/Vr24EZoal6xMqLEddLf
mKkPfewqDQCOA4lWfp5+rJpWwY8ms4aTAZJowKW4YIrqCD4GilDFcTyoGCPO
v1rJUyZ0ZYmx0rqbWoYZxDu50RNI910FOhcIuJ2AtCOLs0JtGtPVm/JspOff
rl8fSbewtEl5YpashZRG9GYoDA1upUkv/SdVgRW8K76VyN20tmQC/ACRh7z1
fXZIlpLPJwLfmMJSinQW25EM3R0ElNq9ozFKPel0ZOLG09U6SHwZ9bRMC/VV
Tn0k4Q3lW0m3iuyrBthDvg7UWJbvl+7tYQ3WAUAc32dcpfEHjITc/ih1BgnB
Oq/x1LjepQjWLpB9aR2dSDVSpO6/yuKilifj+3hPMksyJoGprJwIIXzFyqt6
O2Vyw0VMrUVnYPc6+EPIXAaVoXmI1imtDlGb3IfiuQXPr+U+6o/ZOi/71aGJ
HrotgpvuI+4sbidKW82dZCODnC3SXCEU9qDi4JLX5zpMtuL1moDKuqx86C1S
bZiNUuvQkfaL4LtsXGoLmDSBknt1LFfeyFRMgfmZDxnUWiYjbsQJnvwmbWgX
po1lio9qR8ohx7fbO1fmmHD2DuDLBGT5VoUYH6H+YfIs/EfrbLR+r9aHi8kE
+htQEOoIL2sE196SqOYTng3B26f0FrY+NLwhqDguVwb+G318APdZPtbYLHDP
9rmLxjT+YFHS5tbfi9DGV5Ob8crI4uTQ/qGuVmBcx9Ob0KCQUEFS8n0i+NYW
Z135JUN9wsLMS3b4T/fH8+Q2cf7EL3ULJYSKddlkrpRk3f6wrdn1+WEfEWoo
sKgE3Gx8eM5fY8pGwuPTfOBu8JIFU9z7jzAWUXXOC467Yxwg1tefuJ/Z0Wpd
fRHzLBP/FOxX+IlpB65Dka0IzEwRVSdWdVp9oLa/aVF/H83nbn/rIvxXX5xZ
sIKrOq6Yjon+H8DpsTQrpE3JCj/tqC8CPfhTZhJEDevVeaODdlgqUygPmSps
WsjX6TEwgD0gsEaKpGCPPttTcPlfHMm+pt00J8KQ+BIkfzFtDpUko+jVR6vh
BeLxc7rLE27rJ245a1RZfMJAWKsgHZCJ6TUkOkvYALUZrkZJFJgNGrkOZFBT
pgEQ62PgwD1dRnjcD0TOGoBYw5Le5G+WhBjOymrIfyuojDLpotRM2+Y4LzPM
bR4i7R/V1j4rogIBsfB/KlTL5FYZRxMOBg/lMlLIzdUYeMBW2PmJ/K/tFc8O
85TP1jopgto+TcBeiFKKR7pwdzzJFqe5UYbkYIxXDLwflr5CNQ9T0yrAY9bR
DBNtUmD0z4bALe13+U12SgRLP4z4MUg7JZyp8NPvfIA3atlv4tI5KE3hgia1
lKM8OW5yST7SWCnvxK0xzNlffsFqJatgrbJ+4CkRGjykmmhwAs/UnQwxvvZ8
RsF0bL9LtRHLFO0h1nnqlE1vLoY1/NmJZ4Xm/hiro2uE0oMJMTzN6jmuczsm
/7JBvCEVd8/puXk2HncT53G4h88qDnhdKPQqQhm8nJ7UgI6CbHozD+W6cilG
9YyRgJmPHbMqToQ+Ie4ugprdS8yQK8nBLRzLPf+SYNeDQBJcYDIHt0M4PXLK
fS9NhrDROlPVfWWjYXSU/4kGWBnkDLMH2s2YpcC96r5PGoR0MDVPKk6V+lsw
zCvArhbaxs5C9gyW5zoYusQtcfMED9arhZpsQSezlR8LWaFsaVhqga4pUs4R
xDizj4d74j8I6Jld1w/H8JUKv2W+gf1coQYwEw8FkaEOPDl/7YKmpoE86rIZ
zhpZAEljGcVM515dlerhe2pVaerdqIzvkYdVl69xdlcJDoN/2Pcndy7uf0Kx
CXjLW1vF8LQbBay/GkmrMBUZnRjN/48/0VUPg1nAsv5LiMagHjrLG2flt8tU
0dEf2eT/XTuGgjrMAuR1AKfrta/D4a1hoPYOMr5dgq1RPHoAthZUAZamyepy
XDLtbPgwZCBQA+zHcDdCuWqCaS6VNqkEFrPNP2EoKPi3n5y0o6cyJMYvh2wu
FmbU4VymPGUBALS3ldQEDA6PogV+bhzOBvKh87JNHwHf2fbIR/dMUGklYpva
rXT809EhSknOTE/JY8enQNzBbnDw1+RtzazHeX5auKHpBcsS1yVN0zlGcxH8
AffyyKRhhK80B+8xEcuzuvna95+lkWzHmk/vNjisXOfLCw6ygOp67jIwXC4S
WmTu0TEnCJ/3GvpicnjJ1xE1kUqCl6X5ySleZbPmIa3folBJRMUW+0FOYztK
8kvXEAmLIEPUdWTFagbciqQLA/ogA6J+NNTktjykK64o2c13S100m/hdfN9N
/006fbcLDZwdJ7ksVPZ2zATm1RsKIEOZQe1jfLZH/6HQ7k69ac+ZdqUFt2Yj
D9EWa4D6i8HakZVbOB8YsIZwSFqA6dm0WUldP9MCnvVxv0eiTbh/ldYZeeQ8
cR1TubEMD4dJ5o4roi07NlD4e9ytCUIKR81inxPqaVwX0EuN7/emKNQwghzH
J4JS3gperpQZIH1747x6pGnAfb6iSWvEQwraqDgSps/LMBUTJtolVZEDXM3T
ZalQvyMqCZcsX3JccuptWZPJqPD7WiAVv4YJ0KV04lbEC+n/lpvFAdmLJVj+
dlfU51gaH60pH9iv72ouVrW7YTGDiY3erWRPFKdqdgAb30lZ9c4rlCZYnNdr
G6HOvBOVx2IJOPqjFL1G8yx3QOE1XKWjAfPMq3ro+gzzCTE+Jjpifq1k/A0d
F/C5qjSv5nI/1z3ssADIxzlAMRjnEK+j13ESX0io/jcPDroQ5HCi1vK6/nRF
6+AUzcn8vn/NtX1bJ4x7RDCKU3wmktHt2WBeDPE9Kbardxs49VZXUDvce7Gm
r+3u/3Aj+yccnN/cH80+SFlMImSYm4pZSblVfhazZfIEdrRrQ2mhax1aHZcB
Rli/Q7BOugGKiQk3RC+c90j+UYb1GHcx1P2uMt5OM0O+vnuES/jhIdCV2S5N
6cB0QsGOiz1Cdtx7L9woxR5gILnjR5W8vcEeXMRY0C4HhYIV/MkQ8v2Wn6lZ
9Okvi3GpDb5+UbOWA4JZhKftD4Ay+mf1TdY8h41XYVKwoybCRpKMswHjMllX
NIvwcIjBIC6DdoF8Ik2xmzzxaieS3aMdrCQ8RNMaiaO3F1eLsD87vAPsyF5D
SYkgzFZv7H3X6rzrMWiSWcNIwXs6j4jCZKdDPhmv8HPg0l6N+A8Ye8rlxcOS
hUyMYV6N4SkG8WGDYqvo/hmODtoSskLWbyxcoN1MHIyHcEhNqU/t56bJUKKq
thOK66BHAxrvBzc1lDrIA6RX+RcArXVBOMoBcJN4ygOIDhkfGwok46ZlTt7V
XR2WLZcjmNfkWR4TTpWaiW0LBIUSiloy238BxTInwHsDuTQInT/WnQHlQ7Jm
kHXGNlXP7FuPV/i8V2ew8YqLsTu/Y4IVkdyqXeLOhqxd4PpwTjDDcM/wrHZ+
aaS1g0b7SvFsxbaPr71hqJsL+ZUiLU4WmCo6Qv7v0Qip/VsVgKVur4HdoZ8b
NQGuqm08n9Y012DlLMjS3N/nfXjnQ/H+dk+NTo651d7iRE919ZBcm7UIZHmJ
XJIztGauHPSuV+upYhE7aTwNDLaHuIx1TQgPMfzjkwRohsELC0NuQf3JnKBT
f1LSD/wXaX7t/ezljFPgc2K3dD2JSRyLnVAcQmF7eD185jxK/suo/uJiaB/u
ibqPgd32xQe63Af5vmztRAwl7VAVakO32iHfgSh7B6oxdZZenC7PoqjLBafL
Z1RwpwDCJV9MJvW66eEUjQx7M41tVvXlo3H3Y0M3wKlNn/6D/pgz8ivgUTZQ
umyeu2HHwWtTG+h8ysUv9z2H1FsfW4EAn2HEHYm6oQ4wxI/RG3aGUOU0FQ3b
IZYIxpbdO0mesVKKe8TFQQY1qBvlee5A/2lA/KftjswiQV49dK7q5j2fvxm8
QUWBNdpFz4/oaxdvGxJWBbNPwpfeiUFflPRL+x3KPnYAYdESGrAO21XiSv0Y
i7SK4hXkcnUPoQkM1FvMgGOxznhlSJqjNnjIM5syyaBqW1sKk3EeySvoyWe9
XGhX7850fMGq+Nhka+dyCfpUEZN0bdrBNglMOS+K1p3twUmns/e+QqrgLJ1X
Serz7qzisdIjBRz/6sboZ/kVot3WgVlotp0RAejEle8F7O1Db9fRwznda0n5
XgA2/NKaNoaGdfOr8L7V2hwfddWE1EqP0HcjhkW9834PBR4NOZbFGsYJ6oE0
t1keszXL74PQMFIdVubwAPiDVbVffJCB5R2UQkQgYdPfoODghDlffrDD6jSk
nYnVncyU7NdZJ0tETqN8S80AN1FGUQYlig91zEcUSI2jGA7KuKx+svMZw5ED
siplzpeHN85jQ0vGKIcg6+bd2wCL45Rl1lzR6syPMUVHnkFU8G8lGgBT+Sb/
EQsLUFMAfGT3a6KWs0zN51EjZgYpyhds7o+nxk4/I2Q4Wip4r8m8IT5Pl0eH
TP6cgv822Kqhp6sw+VgxKzzKsuwOnYoYMs8vvFTZVoHeGcGOI3IJ5dYMz6FO
ydYZ8SXwTKMqrh9E1wxgwvYUFr3SzUEH3Z6Uo8l1fk0I4LDXmfZLDUfzvGDK
WE1PG+kJRQ85yt9HVL2oD3vROdNonS+qINYYCqzGXGmfu5Z+I1em9Z90AVlB
wkF0vEEM1DzaY4ByesTeuJMVYzoWU4IqwqJ64cR++R5JhJe1o3PuwmZtkaZg
7fWNEIQ03F9FHV4fmxe493hQrspnZW97lfF1Ap1DRD5K50F+Dh5gAZJI/Fn1
LAKH285DLK2jPYsbZcc/LR1AzD3MHGyco7jKokFcemB/E3shNM3L5eOYltRe
2V02gbfEy7Hez+dcaiaIZdLmNm2h1Q47UyTvLdjPnZcWZbnNGGf+yrf1wfLp
L80zNhjqznExAJDsiG+JDEOuRhIcefFzlnNypUyeCXOoMFZc+oN1tbj4Ng7d
ovM5nzb995xAeQs9oZi/tvt3lN9Ok6wynjRB1GN3+SBiLywHMi7Rl2ERDpot
aVtB7B0GN4Yb3/e6S4g16VboaEQfNN84cxbVY1BQd5o7Difxlqrt2zm4YrA7
o1m93ywPcFFgA9JHrs94kfvP+RAoV6qY9cMP+yV0wx2f2biadhQHKgch/YW0
IPkFncx/kN0lJYRT07luYYk5uLVirqoJ6VRbhbhtNe+Yi8nkyVKFsq+d7Ul6
pT16XkLFrqZ6ikdO1M4PQ9SUm7kChqPmuI7yzJWhjntEG0YrA2NyjoVYCo0N
FphZi5J3Qp4EFT2XWXh5Ef/Qy8FD5i+LnwwjddVluqfXNyzhbx16DFoI7y7J
EhbOxVKqsqaERpH5pz1iXlan76ihm571Sfc2m+rJMlIu3d1bt5+ld5oqJVyF
zzNpWtFEdQeAxi2gc5EGameXV6wKwmkzPqsVWTwGMgYwOhdBeWbCm770Ng5+
tb78KP0YYzl2bHAznZv1EuGNOdlDja2maYZWhmG2lyRy2h1eZHJzowIOJz8g
pX2gA16dT/wSzQfUxxV8oIxrsri+MaS/KyWRB/ufz18M5S27JaR3JqHp0ayP
azDYgAbufGGWQn6bEUNYt7oHtd5QQVr1E8X8zPdPpP2NxM2fhSAOVXljC8q8
XNWVTyWxHeSM34k2cYMyAd1mbtabdkXCk68w6z6SJhxqKxRbLc7TsBAcpt+n
J01D9tidMliGCAv7gCrV08VTKJgX/zbvx15sSY/iInJP9LAOaLZ3t3nmiQtq
h3CVKjHHJWh2Tyx66K355Y0VGYm5QqZwDT/aeWkq3G5tuJW9T8lDo+LDiaSV
AnXPEz+/ALFt9E9T2kIJ+SgB9MyqiKyF8azOe/rrctAcQcE4E74gpmCchl/A
hXAe83n2zXhv3h4EuCscipU2MOPaOlGU2qxTYvdHDVZaH1qE5dLSHlBT9NQx
t+jn+cE7iDGSpS+XO5eiYuM0b4wi0fJYd3uu/w9Glmqgbp/GmpoWvT7ce+Iw
xg6u4FeiA2yJ51oyodZkrh/qLnUo1JGlNxBpvpkzcM3FWoMt1KwlcvB2Vcg7
ZqtUAjoLqY+0UtrFyEvT/9DM1MkSKzL1iBo7RXAKqWnvItTu8CzpYIfkUpzh
9urmGcH0bpr2RrvomOG93i54tkapRGQNitgFsi/H43KblVEyf9b/otc5kHk4
oojvjggd2Z8zeUaHg1ZEbiIdho/uZZeHK2G7iwEoT/5MEMawSKfc3Zq7SdfQ
4qLEmfXUiw4x9msPrSppQDXoYi9isYpWZJy10VKU0Xzzo4Dnrw5nn7IU4/io
iN6ANESx7q/semx8rtB8/2AbLfmZoqzZDC4Ot0IcG+QbXCvkvp2RzDDCdpfp
vtFP0UHqO3pFe+Yk3yH60nLsTCOMYiAhf8hwdYNp4fvcAGHw21YSeYngH4MG
XL7pWEmwlNTlUysvbJ/IVvuef9w9Phl+8m1jmgWN4L+BtjiyUnacamIZobCk
8mDW5eQEq5X/amDFvlTpZpeTDul1LMvz+nODDOZ/p18UIVh0y8dPI/XDnnKk
/2MocNfbiKTW0lBlCJtuMH6JW3HAbigKLUDxlnfcaetrI5Ivx3OXEyqDXyfw
VpIW72FAaYd0HqDl98Njnza1oQYRjfUuu5tIoN7jTHEredPW338Mb20w50xg
+cw1Rqt/TAEAjgZ/qi+2dKYl4wZnXcQeVi2XcQ1/psZ8o5rzz/CSazMZ518V
EemAlyDMzW2Cv+e3xLKiG72+/ZzQokjVidmKFV4Ooj7YlD9L4gle5BTNjb6v
RGE0DAOchzNii6oUXiuWi91Wj+k0IayD/OKEmwfFzc2HjDdJ+UzPKq1er0FA
YzAAbmmPE7hREehnhl1nswJVdf+YN0jVVFpr7H6cw7ealpknA6Zh5YHKdGFI
9lwTavNyskJMxBNpMgFr4INxcth2p/KcMgTS51VelB65yTbsMeb8Ws6uLhHX
bXeAC0i5KbkJObowwFLC3m4VwZ+NR1E7mr0MorkSiNebg+4Rd/EJviAkL/Bz
f0pikgopkdJezsUVtEjbEW3aOrxeHD/HNhYUeimSivLBOsnMlhovg40h5IiV
EbjSLVUbAm3kthzWr/j15bs1FSi4kF7RHdfnIdU91L/Ksw0ZQYtFFSGhZlku
l+lo+lREbKnljjvP7Za2QJddOpzNJJHw/AhWKyWSAx2q5OjV8XpuF/AziozO
Sr0OVC6PUUfnTnfKeYeRGCYjQdRnk9E2fM+3xWph9cy/Z/gtmjROE2fSLXvk
cEfTeYB8pKZUextdRur+19RrGXnL/F9/klZtxRRFjp5EphsNTxJu4u6IzKSs
mET1BzUQZii6C3DporOd7Dhsjmten081nfta1EKHN3ibie4o9x1OXZLPAlSV
D4EuBWNw9kx3MuobAu+KruSsT9q+kS+wUYfJOWXvq3ukIP5P68m+Prcx8sag
G6mojQEdhmGBaSOr+IsEbHjF4rWF/NAC/y/CZpY71LX9DP4KiNBToAvOXmgn
m9deJyxLBk0K/PhGLqtYW25uHQNz9JvQDjJ6CPPSTGVl/CALtD+rUquG4fND
HPv3j7t62sYfzV+JKnwMDJ0VND+4ihjJLFReFwTUowSJdsJYr5Tb9plTmw5s
gdyhHIc9cvNwxkNLS+KH6Wq5hBFTaTe//OMAr46gcGRQ7R7xAv9AR1fHrmYZ
uoyjRizg3HO+k2XSi525fBwLt5R9ULpEmB5PrX0UHMoc+o/XVI96I4KhTVNP
MdqfheL+DrPmDJSSNznsuVZeV+4Rm93/1Qf8aYss/NcifDnb1hvyE+y9uNg5
qVXHfsnZ2gaDVdrLlH9jdV2/kXLs6QxMQGnddM2bMEDs0UNTSb1bxiR3dDxs
8tFFdvhaqAf+YsI0+vBBRmsww5WDvmU5LYX2nTa4utu/haStcNTXoy5tTIPs
p++6FSFargAKHg9GFIcypPluQ2j9Vr9aTjaT+4AeVR0EwEjhJBVQzj4vTZNK
k0FqEQ21VEzRxZT3KmyyHv7eWx6rv99IxDdPAsIj4pmppQkD9zHcglTu4e9V
EXfAmG1FN6O9s8vxePPJ4rpWmyVafuAo9NFLF96xgysr3TW/PAZ/IQfSRCLf
LJwRpzrT1WpEChg5+tgR0ld0C2CmfF9NspfBygqfqv5UEvPodQCqfiWCXRiV
PTMB+2SKJMKzzBEYjb1ePI43er+JQ/y1fwrUbXpY2gREOXyx3QY40IZgr1GH
jPD719yvxEj7Xg8wA0GbKPBPElFzVn8X3P55UQW+1gRBz/fcesh8mnLuOogS
6SgEkxnlDlVyOayK1SHFqvQaWyb2IM658KyNaITqRLVWvuVYOB63fqpjDx6I
rmr7AK2AYFD36k7RUPoYDLOhcIvENJ/5VdbXuEfJyh6X3JYfqBVEeTig53he
PtQwNHv5Cc67EjJfux4pzzAi1BRSl7rsYyN1gppkMnWWexP/sBj5tFNOgmT2
ipZcm0LvmnDSyZW78zbfFMQbm+AFhA0vX7WIyUWQo607SeDrtzXGrwO1Ffzq
FAjkWz7Q0kHiyqVAE0JlCZ85ltCR671UxVhXnVCDUFHk2pbBjF/Knjp5XY+k
jNRsHYJCxU0ET1BD1lPlTm6sJdw4yfnI6Bltk4FD4bX15w1saWTLCSu/Qux5
JbbnCFP31DQ97vc1t8xig+gokHwOdgrWs9c806wDx6PQZDA3aLPa7paYWWxk
NshqAJINBefUAtU4R82yUUl0XzFH93bfihEkKHmeq+vTmSw3MzfHQug+k/mk
4XCpY1pu4ZlmZo2otwWyQIjbVb6RoQzNiJR1yHx858hDsHC+CCtR4hVZH/FV
Y384k/1495lcamqNVcWAgfEq3xCuc7yUgKfbFQM31xBVhzFuS2KZKBENECBx
mNHqRrw32Z9nmsPn2UJlouYCCcO99tWxvVRtxMHHiO3nfSJdjdo8p/TyAogW
cTGU3ua8CXl24Riaxcg995AaxwFi/T0QyIdJEalNL/WIlfWTK1Wq3k/kSjsj
B1SR5BSiA0wRaCew5B2tLIDjLFJVFVbHjdyzv5VrJWua409ybePwv1weuHQu
u1QgvnsK1szzW9PKWVi6s+mHPWeCXBI7DvYKvAU10fG9vdnXMtQDhcg2o7n8
y0PXQgDTUbNABRMs4FQ3mJexPjPTx7cNcFoGHLFaw0a56H6kBbAWC/H5r3w7
iIxWowqg9SpLFg9GefI0XWPr0z9hpL2zmPYuWIj8VmfzHFdqeR79rXt6qTXD
6suD22VPrACTjV+JJ74E9lIS6j+yYQ6Svl+gUvyK4y0TffZBPG63VH3I1dJ9
9WzVfdxcK2rHukHk9FZWgqreaWWJp5Fc8/yfyLC9LQC7eos8mOjARAjopVaN
XrgOiMwJ/OrJYKmce+j6tZ5UOWj/N0HxroWCdDbG3nI2UOdNru4Hpr0DWSOi
4oOk549wZjY8P/BMTXajIPHLWab7HX9bKMUmspWIfps8NxciwZF2PV+SEKZe
+hV+JlG4/cNvPdNRpigW6SIOvKmAFwN3cZvzKJXJMODozVXkjIR3MJuOSjLr
zaUUwl7Pp7mfOmTLHY1bfbxTfEYw9m1NNPxf4GSTxZHP+pmHQkax96Zktvgs
XJDVZxs7jM6Mi+Cc0vKBSC87DCqztK2ZYcBk0TcYewjj1cXHurORCaYqRgHB
B7N74ptJV1+1A1X7dvhryrWWXcKgojH3Zbqn/wuR+hUQIS8erK9t6Bbg+OGu
1NFBpciSmZhPUiEPlRhOFB7on4jw8KlZVCBqExav8zgTBkQFhiAT7Hs4L6xw
16umbzF8w7jvvGp0pWazUMUbLWgSPINgECYLLCldesuhZVrDiXTL0wHp8ySM
4hdLimq0+9PjlYWrbsCpcXfM6Y8DWUdec47IHpBasTHHndeFcBcyNVIRtt7i
EGPF2cnoHbjPpx9oSy9+57EYlO18EtJpkiTV1INueTzi+wuZxjSEmST8b4xp
hMBghAxl/aCOroJixnVzh9aZZtY8UOyewGIAIGNGM+LbR3O5Lx6d4NlkBGRq
ZU4VgzHjGL3yvP5GIIoZezrgGaPDVVfuWOG2loHKZ94oNjPd2TLYmPLSRkmJ
dSpqyGtdyb98O0qnnaBhvVCY8T3maevYwnFBDlXIBTp4gNIkyEDPqVY7PSGW
B0BBggaqZpJ4ryNo557u2pvBwaMBEVb8UMak/5poUvBU3qk52DuONIerpPIH
bp2LbBr/0BcmfReZO7VVOmSyxICp572fwbAUHaD6AU+W4JYgS4NKwtsqUGM0
KB/6r31u6AsstnSBFzfxNFi+5xj+Wd7JQW0ntgmmtXIsmRYpLSUnfqFNt77Q
aQgbIy+13JT1G97pNgRAHbCAcj9Q2XyFgwIKaAw5mkZ0sx4eAAMMTMvPQgKS
4pGoncoYnDvZFm58mSQ+E4EJrQNqEQG9PHAtm7hzF2IlmpdRi4aa95N19Cvv
DgjgoYsYGL8Fcv+wsXMFgzyXXUA8W0QrN/FCPpfhS8N5sg5VK1Wv8PP1Th95
xakYRyHZ1nIbicPvoTjkBOBgaZrhZ060WhC8Bjv1g62iIUYQlHsoJJMO0Hs6
vqRDvS6V5jZAa7cJmhewYvHzD8r6/CfKBciy0JHyNxCvgs6W1ewOYRp76QZy
VmNhupp1MSDzYF14XiboeS1vu6GrPdCG/ERhM3s22yR9PWlglP+rhoLWm7/J
4Mtu9+gASkbITFkcCWFnTOO13Loo4Ixbx+QVZ2efWt6zjX5Xfsxle+D0CqND
wnY3IvfrE+K7Cp5EQt9m1lFv3dyHF5jOWgOX+FYhq66fA2g7RglBW1oehcpA
LsdtnW8tvG2etpJj5SigRaPQO+e64PpIeB7I4urNpQdgJNAuEWrkg0FO+KxG
8m7bPfo1QABC+6tObdXsGBoC5M1CZTIkK8ErXOAIx0XyeW9ieEO7ilgGKmO8
yiQbUfA7CjwQXo0bwDdVQxJzCrzUctWOnGPUuBLxbqHb+EkEF6/kxZ6+uWwk
IR1P4E2zvbK5ctYHjvT+raEK/B9uzj+waTzfVOVL5Y6jxapUCw6tZKNTZWt0
hDu7Ake1/X429ySJdMcm/PtlvlQYswk2r/fSsKPPzNjJ/6sKBUD93HsvHEY9
McZr/3W/WyS1KLtlRdYtZ8Y0x6aOEirdxlgjsaqvqAZoSNfo0ABg40JwidHh
ex8iBpOQZXGtcDQMcDPl78Ix5v+OntfYlG6Xfilg8Hq40tBtgIPN6di1Nz7k
LT22BXATh9Is1Y0/yCOAD19we1TU3l4PbeZRtv69pm2GcgQH4PbvhHfc8Srx
D8RD7zqAWeYUsoO2WBg4/0Qg5Q26ym8UFXa7XP5R48sGU0rDt4TApuPwjV33
6Iv9Ws/XOxoapozVb3M/COCyJfBTCfCqYBTKDVvXYBaol6bV27t52Jmavnvu
va1Rhx0bXAkIoj0Auguf02/Mzubkc2D+M9wD2szFebAfJtr8QO6CBp5v+DTc
Pg1VjswXhsBPOCVikb3PWqCbKFT2m5/yuFPOlTcAOqgQgQXhwS3zc9oi4MTs
342mv84EPJCy1GUDccH/gbGa0zSeVwRARYaVkERnNqBHo/XAWo1I44ir+Qij
y+YdF9C73fDMbX6q5p9fb/T2INYQ4hbty5PwOqWaK9ia7hm9xT8VtmH7dW6D
HPuatJk1LhQTr2PnqN1to92C2PkorOz1pMuabns8Pm1d4OcGRRV8TcMIoeG3
FNvCU/pY8T56baeXzZaxXo4yJ+bYM3P/2+6i6vWynvjyFynLIBc507aysJYJ
i9K97yMLVeoxKb0UD3qe9nFb7N9wwiBKEN+P693uHq4/UI3R3CqML/4Zv2Hz
ORjNHWaW3QSDtLaHOY/YlveA4ATKnlYEOlM3yeEm+TgxLR0PLoVBlnWWUw/h
hq6Kdf4WnL4bGBbQ2MX3vfMf0qr3ia0vAXmZaH2kQJ6zXy3djufmfFgEXNan
+G2bB4ys5KRAGPp+LEwnOvWyv8vUDCv0IUWvkoiPITK3yI0szEqP4O9YQfK8
rJ3c0SJusWRmsoVC60Uor/0D0Fy8RpsR4/YEPH9iElbW0QoBiXNuCYR+iIq/
C0g2porp2aZjkCB8+BFB4uTuMqmNecy5OsGOysHcOJjGVKVGy9Ry5semB3bW
jzSH1tB2at2qE6n0G5I8TfJBmduSjgPA0OqBNcgmJM3fjMjAxX0aPl+8LdJs
2mQNNc7EvR3MQWIVS1XGSMRGkWzndksP4aIr0L/V+s7oMPpxr45Wx0GH7LpO
BV1/3CMFdDABYWB57zbKuG1K2LkOMIpxA5ILK/6hqFXS8ZOcNf4uPj0uWc/1
Fu5ZC2BZxq39KZfmm/iElh8bkVCjM0Y8BVYmR255CoiM+Ay67cEA9gugVbNN
lYAhrwaus2iEzeDdSC9JaNP+k9zOCujecnOvPbH+IZ/bozdetmejT/hRtwPW
qWkgAz+fv09xeIN1lpMLBlhltJ1K3belqsrU3fjEHIA20fM2hNP4BT/4aprr
zlaCYieerl8X5h1LCpYjGHysfQCTeVwPdJNy8T+cpQe0wZmMngGrUlo/vm/f
tDzAY6TptNC2Eos6qEHeq7SnxM+b/zZaIKNcS4qjc6tQqSpUPtK6ObaH8Shk
TMUptFNwBUkq45Xn6r+KL/K1c2u09Wc3ZxvaWE6+C5Eo/rAXcCdAuMtFSxQs
+zwIrTBDjWUMj7rSQn8hbK8FtOj6g2SHU0fgP4VGjR7lvf+iuXMqrMtfIdgZ
emP0c53vr6hn1kmdoT3DMWuJSF8ecoiy+tTPR1r2IqlqD+GVyuCWarrJXNXt
8EzyNCNcqtCL+/rqa0mpYWwKRNp0uQER+S8Aln127CtpIrK6niEj2svXwb/j
RSpJHqngtH8o1cLsPj6YjGtAx58C7QuI1vCAJE4kshAzUEOtnyjvGF4bi3X1
vRLA138KVkXzQEU7R8YFecqXpsG1RP84EZ9E7cJJoRzV/DTBPwYuuIYMbGTe
PAihDv5Bn8uP1QraOJ3kYcnySDm/3dW8KvAROAVGtlqIU4WOAglzGN4GGTT+
qSCTInklZlwxCXtRUlqoKGlsrvABILUZT5INQOOgaP5Gtufpr+fJt12Lx+DB
E2EAqIrUQ9T50lzYDfZwfHxTHhNsGAvX5Z4Wsrn2sue9mitFgQZTwhA/ZUkk
czOoUuRoI6jUDBOfqoeSRv5k16fntFmzNRejhfa1KPWofQI3FDu92HJXIkLg
h/UQUUtHICVJ/wKuI5Ir0s9psFN3N8WKzlPTRurjfsUwZKqQydHwLWyuXGph
LLNCmr4227wnYSLvJbCAVrKkOMl3B6lHRxXdcdDsxBxR5WW81vhdgfD6ENyb
KIxQqExfoEXuKgJhJ+/y3/6nj4FJypWgNUGmHTEsGh5QhgWEDcFSj/VoiMVx
UB0GZOuF1xgdhl57K+pbZ0fm6IidadEATylmawdNL2oxRaGEkuuhQnJxqpzD
MvqUiIakmyE0QTDY6jFzR/21CZPYlRXgvROCHWSV9AD4xfSNrNUcHqA2459d
0Xb23R0ceP69rtc/XzdGlIcoERsYNv0kOxNX0zglQAT9WC97Mk0tZAkhry7/
o7qHTVBY6VMvGGDL0MPKnwbKAS86mJ+pq4ncnKdpq9c4wk99aCuqL2WUNzyL
k3nivADnWjT4fqtNe+nQfnhwoKV+I7y7qa9WMs1UMs47d1YIsOBbWFZ0OlPC
eKuIirpTsPT7YY6tA16+lrQUgMnqNCwafEG7QSHqUz4zZ6tISEUvXlydbcho
fVwYLBMPw04QXEhrHtH3MqJyddhPTnS4gu51dC9KzFVeG8Ni1yVvLCYGBI6b
SHzXxoDSRRQ9gVMq0f0va1NBMtlcMnqZAxcmlfKU56Fvr3FDU5RPStB1eXEr
Fr2OZxwyBZYyY5vvH6R0YR65DbDVY7YdMsv2eNrNecgOFpZD/BFQYcdzhktV
6RIlFO7vY4FtjwHxFdhQooRvZ9zlF4t4VY1gbouViEsAHF+b4J9K1rDjEUQ9
aRsszXju//lNfgkNPajCaT8f5RJ2Yyjoew5Anue1C8YDj5VqtGxklfR/uHKc
ITX0zgHdWXYkezVYWqecCR7gYlTV1mn0rN4IqK2faT4mE5kQT40I/ha3SVvD
FQMSLjVuT1QTJV4HeN2TT57BHylb5uQOvLvqo++m9OVJ1yTi/Kj/r+DdBbCK
Hd5euWPmQucR6J6e9II6iAMY2+r7vDqKHomJj74DT+oM4d7Cn8a1rdIR85bW
1x6r1veh8dRHHBAK+KvVyCWuHYC2Lr0eXzAV3tsWtqMcLwaWtaqoTOP+knj+
g45jn6Y5PGRfrVUrCzr5DQTgFuF43jgGZ6nVE/N1oEM/3sCCmwpgMpVR7yJ8
XK6pY9Uccq5nCBvXWg24G0BrAds7JTN37a0LUGdmOJfW85RrjrX3p+BHG5hv
WwKq/ziDMzGOrG70mym/7iF+y0Oeytsmk4z+EAxaZ+4aHLhFQVw0dDy4aP87
Lpz1LFHn0lUVeDoN4+k/QiDkCnYwADFJG/slpSZIaR8Lb7Nrn3tqVC7zAX/f
lisCQKFXwOOh8Y1vuqM+jzzELIGRFy3/+t1NxlYYKiiN/24tjbuS7XR47W01
rCFOPfQ339zR61X9/7NpW3J1Ec8H2LFZg+OwBKGwAhetPqB3LRAR/bi2wrpG
1NtVk8F1GuV7+s5V4FWkH+8V+04VyFVLaicXd9E/am1noP0Ps6bcu7y6CuBu
/CNmdXNN43swP3hzHZXXtyWBgl8YKUxAYq5Yom7/xEmZoZuoGLfULjCiftsx
3o4KDlsPfhP+xhkHFiBS3pnpHJPBoxsFfsSEqBnrRYOVm3DWS2mdKA2RM0qa
mu56P9STTfYiNHHnoaJizw0GLtVgRj+EsqnhQX0JNYyAPIgwSMEdcHKvgI31
JLXiH/TbmBjGZA3M5vE0nFgaar4rwmwi+QZJENCrGX76l/7gDrHlrsdT4aDi
auxkGdo4aivAZFWFFA3APuO+F01Rt37EovMyxP7KJAWSrsIjcc1voglYCOBg
jQ7tt6UCS1iah9nGdn5e9TFaNkgoZ8t0VTkkwoo6U2myOh3/i/0fgTYMIxbN
GawYmLQJgO6RJXkY4fxtkrw8C5SUkEmA5pJj6iDcZdvD8cvMPaeZHX4TXUjD
rUJQQM8t5FfBtBXJbvJhsxKbklLyTjTqLphpNNmWfgc5VNXg8fF8Ujh6PP4m
QNfV8J0+8F7HIA/ycZg+7MK79b10HYoVULFtGgQz10Ej4Oa+kuGtQC3WaWHB
rj35Afa62LDqLHrILwXtUQPe91QejQWPMej0jN34FtNgB4D0AD7J/uFUxix3
fFKZ+n5NcH6YPFGXH3TnsEubpMtiVo5KliaaCYG14oKyX7PXxt/djZ1Ql1HC
YROntocbpOza3vprQv+ZIw5ypV6zw73Zuje4LKX+ttTx5rHW7pNhxnRKTSfZ
M5qDFpqZV6ehSl9/FbvZSxx/pyF5jwiIawX9i2dPizPT6PmeiZ40ZVNnGu/E
y2pljjMAOMr5m5mdL83Qq3Fmel6FDs3OkDEbtbrUpcyM3LyXOF/uzBoz6a1z
u5uGfoQfrcwenTgfGUTvYKKgnfurL/2bt1k4E2H7hYd5joVKNy214XD6HOzA
P9y1gOAc0nVCsmlx9qSoWuOtRsjnGcgPqowVVHnNEYxMFajG5TgNO3bknnxi
F+2uQt+8pXD+GBXegkZSqpoSBXg7tmO/LOwxya3fLkRbYfPYgtVxtUJtrLcY
iYLLY7sS12KjF0KIEXhkYRbOMmNHJyeQRpepUbs9MZ5peXUU67B7buP4xrs0
xdmSVL9/IPIAuDccmx47eZ68UFcpfvogZEff/S4y6uNXK7tmORshrcqSOb2c
mLaMdKqFl5B6fP9I5/FbNxnaARTZFkSaHtsYPlk0cu48LG9RuPDpHlFWOcHk
ztGMpUYjarbVqImsXXILiIyuO9/17mWfMiM/pcC/oiZQE/zNBCaXA4NjY/n5
juUBUOKFKatySUH9mOwmWZVFG5fzG10ytwaVXPYA9QnA0/TN8utPR1B8isZ8
OUuaxZKE7ViOgoj1n2tZ5b8HS9/Nt8NVVTzF7bsIbNEnLYumfWqxca6CmrWr
66c9814S+k4BfZtRjvCwTquuc2iHSnZaM7FIliSsP1zi43+m6tXqvCb0mai8
ut/5GfWcH3JieP6EdsLQ5zuNTgo6YWloIzXFNQ+1HhA22fG6u5baLfAXp7n1
nvJJV6iVkfzRnzXveltzO16jG2ZniJzxDQA179oaj9b4Uv8kS8AkLVJ9N390
PlDnt/kf5C3M4UKtWqQwFn5XF2NNsvE7ypjU1peDm+9MLZFO4acBn8NO3MCA
mxk1zqfzTMttMtdw+I9aDPNRjS3g62BR9FGADidT4p5biSn0/mnzew0RXE3l
tCbraWeml8u2eZKHeX67DVMIqBR9ItIhLj7jxfvnn7FtQh1CGtZqT0TRXq5L
+5/LhFNYnOlot7SRrNgy1wIijv8GL43bl2xgUoxn3Vgq5px+6F1rKEDkgXYS
gBO6WluYlmAcPGPs8P4wAS2wEzBcDBLvi57WySPMOVwbDASMRaGhdAshmPHg
c06Ky3VXZie/A47WinsA+AKYHL/VvBqEqfYp2TA1Uv2QxTn+CFWski0FLpzL
GQsRYDj7PicWYEXq7yVUR8gv2FTuJ5qs1KXCGGBTklLo00XR/sw1SsQHslIL
3fTEp+D/gZAQ4ozo5jqfP+4wu7GKnRVVLdYjvbnrYBzWZOZ3Uh50UXON22xd
BQZCycyYf/rK97jTpXT3YGkkodrlzbMaqSn2GIUXMUVhvxKpqnS8zJRDjvsQ
gpLOTNnixOlSGXIqr34Er2FqgRzjhcFMxfZot035Ax8VSvNXElB7m3zoUkBQ
o3Li3wKv5DIQziWcZRWzmR1Tlx8R0pjA0kWH+Y838hWiZ44dirHM92PSTF7D
wC6R8GaRN3VPVNx//Vxzy6dX/lEgYuSCgEUAzMc6mZlOFF/nL1kjCB/f9aLB
A2cu5w5xqG1XvyZj5JRtjqkI0XdZQpMSjUY6S58BrZRUbxVSC5sSEqfdOv4E
azzuEX9l8t61985zFBediFFOET20DwUh4mctEyfe3Wgb0hU0Wxp3pQdG2qXW
b0qAe5A1P7o0TrlLj26Na4Esu7UAOwIall5i8jnk1euR8yaAeP/dmr82YYJj
ikCqkoLVF2PGpiNYX3oIoSI7eYObBrNMemOkz11YQHo6izeMQspob7aU2TaK
OqUf2qYti6/VDa9gJEH4/nf7P6PP9Wiuq/Ju0RRu7dD47pDBEUbhI/spP7cE
rXlIDJIaqc3qbvs50JWqIhqD+a9LcfniL8U6zTo3/XOYPwM0tnI9lQI9/1hZ
8IYQ+zkV3NDO1GrfDNg3azSBHWFGk3YZ4ZNTM25lzM/tGQuVAZTjUTp58izv
q0SuLGv5Vb+EJQWlARNR1+nfhDmuE9dXwx8bLSmvmW3na7Vi7+iP8NyMh9MP
P4ZoLq39YFYd21DkKiOgGmwYbQc45Z+f8tuAgAj5bVKsKISZQNeM5J/cej3i
JzUdPsLE6kSexxVH45zJqdYoaOCR+59cKyPWrEkehuuMAsRY8qxkwAJ+bUO8
ZPwbwIeo93DMmTzmqDU7pXymwFrOpZakx9Mw+d0QPZCUFOsREYZBkJq7t8FV
d+6LNLb2dXV0nPIvf/wkE3ZvNZtLsPb0TaYhKwrrliHJcPqUMnAKN2FfYe8K
zlB3oVXjd47PgYCwxiHOEq8ndLmg52Knf/fPYLUQabioXqh2Ikpie4NENV8s
IUWJ10OTrIVe5nQ0xRCYz3IMKHmp2JVd60Uyr2MWG5ZCAgEaq07NVa6zHARI
LgNAD5bL5yxPbWx5wlCDwViXtMLHfMY7VP9fos/isZ50WEGqtw/lM2m3Oa81
KXmfel+Vy0SDQwu7xfmr7Fa8u5OHESfRti3hJNXbhByQafmhynVHCJit3QEa
rjop2SPWb81VnEao5C1LXK2R7y4stf8Rl0aynrV4byDw9bW2LZJnzurpX9Uz
fbh2Upp43TN6EI8vB2fmdswGlOZ6UKTjRlsJDn2HN5zd4OmPw0cyboDssaY8
YgIwFqwmhM3HmaCyXTrWmH3BZU6P2JW9X2ZCYgtt0lNrDdlYLKkhYqEBnlFZ
aQDj2lCBUwjlfHVOnr6tz02O6SDcnJefI46exRxuJdl63TXrsmgawpBPeaCj
NtSg9S6jNxg+Gv9wUigQOnBfmGyh2qZARc/iW3UbkYCxta2fO9th2p4AgjTc
HaeovF5kwzHtz4OsvJUfQODEG03zWpqHChxmqBxgNXSZd4p9bCSE3ysnRAn5
CT0wOmWB79ZX969P+qoS7sX1A85FAGjO4C4Rkwg4A3bqDrVQf06Brkv7fzrD
n2U6PLHjqzJORiu3Goj9FxYMBSGyAiZ6MN42y/yOVQGtW+e9r1mXAGDuFyYC
+FExrg3Yh43bXkVA2dDtR8KPNQ5g3tKtByVFXUFyZEtePapTS8AjzXFeWi/5
h0g++rmQXvCXr0yJDiExMlaa+od0dOsBXzvLr2ob1QqiB1iKCMFT8vOgu3t5
iJ5YhXdPBVD9TgRuwm89r/mEHDGtLAmD8QmnTNKAT8kaSJgJKpEpE0TewzJ/
DoJiNyts2uhd0w1ddpKlUdlGn2b+KB9iZqwrit+MEEna1PxXbw+60E2JB0vr
0WKkRFSLiZMMgJPPEMw8NdV1uyVxjwrj0PKrMnSe1Ua5ZFxVJ5/ZP00oXkSt
gypKJLbDnupVke+4qqbykA9esHMruXF3IdokoLMJPh5KhHr0uh0pTEchz7Uv
P3e3tdHJZpUowT+z81WJpVKTi4KxoLhvhtPYsPuuJXShLpdjymmXom7Byj2C
rsRJvk4K6enJviAA4U8I2cOp6pdIvryvrd6aJWckZEA8MtSa9xnM3NyZ8Y8W
iYQK6ET2extktjB4IQrop38zuBK4eBsuUAE5WXX1TbzBYlncegqVbhIlUL9x
vHIoIl6EGqadP1DIB9qiSFwfjtjd1zGIinwFPt8b4Kcu16Ii4nbFaqfiSe3V
EcoyIkuwmIuOtX3fWzN2Gea6ka0gYYA8y3rDLtxRWfjoAkJ91ZMSuAm8Z/5x
8V18H/OqH5ojsotX8pkc43Sd9FTAKcXTP3VJQGnF/PrCSxFzZMtB68YqZHWj
WNdHxCKSrJ+Hfj41szYNak1Hc1bFfGxFlS+ZDjvairqyQJSS4NEy/Rw4M/26
c+eu8ARkceNamukPFpCjJMdQmxT954fK2PZCaCo3SUu5J2k9ovCO4HusaaDM
tlIZqAXHiNCZBo3XFzPOD1bPxgR1Ffup3EDaQEgv5lahydiCG1awH9C8WAlr
dBvZ7DITDLhJWb5vqdHlTDo2b1rJGo6oyPX3dtTZDP/L4ftSJMpawxkOBzEP
yjf6fLIpQCpF5X3Jc4hSfBjUqhIubAi1TvD9BHCtEzcFZ7odWHga1JcwySux
G9EVVR8w/emkkZY3nOzOshvF6vL4pqgrkxiDzNIaiDhxg08ta1NJ2KCIikr1
bdy7b6oz+exBERt+SwEN8RJnPXNxSIAKj4xximr//CS3KbfhbBh+vdnKfWKr
/Xisr1WY69zHdrqRwh+Po69eTJkKPb0/WlbuPtp0eBmcJt5Cf7p24C6XkYLg
Y5VYDZfkLSZQuc/tsh+iZ1ygzffqjutyPhApxf3fBJ/lAkMpNPFvkYxzJEGI
u/RpQSc07ddOAWVkJWcPvpGjgmquLV65sXratxZJuhZEa3f/xLSR0e3yLq4l
CUUxutdsuhrpz0CJIvH64BW487kLrDFknyUHnKDiKKOVqXj+d1/zvwrQJV3C
ACF6tphPNez+2JgeM+4vrBvkwEaENqojs7q+Ej+qmZZUj1PgDXjRRlGKL1dN
pk3zZyJ/qJiXJF/wEdMEs6pcnWYReVhL8hLE9uOvw71Xa80NCV3ILDyuc0LW
r8eMMYDBT/cnu9wo1iouogHUQW9iNILSiNjzTvSxm0uBP+qcGOPL0CN66gox
Kaf9f1nZYWN5isLRcVSw8Bcri7jxvtmQlWM6iK1/JbAG7YzeIbGpepfgn4CI
oY66loBdkRci8hTzyzc7bTgbSpTR/+okFQ6GHcB/w40hVIpZ6cbX/Yq9AXz5
B80tiFHM/rMZ2GiBbbxr5jODTmiZME/NWOHbVnHooqhqUNdZwNfldVr5hT6R
xNAV0Ls/r7C/F7xreTSxliTgXe8wTVI2GbTNdmuBGxfTndmV6C3vDVzdqg8g
y/XcRvH2z78uJstEFUj/THCU/ytJiOAZrvnycuEWzbnW6po820CrE5EwHWpq
dm77m0coL+UqpqntXaRbJT7H3Ak6wh8I7AOh/dSrX/Ye7knzJCe72rLBunr5
Mm0VJzyKUy0ChASdrIDyFRZk1tZHbSthVTPXpFr5TxopK5rupICYuXpx62po
QPQ0RyHtXQVI3PLImWq0Cw5cDp3209hzLk5ZsbuuZyX9YkHON5B1hsTleYla
V2NPbjDCQ8s3ogjBUSUIOpuJKkdi0cfLJaRIBMDYSAXaTyS+tzWycKWPHuay
kSybft8cd2OHqoXsB/5pKHvZY9o97V1YMtkrb7BchLBdPkbdwEOilu+qMiGg
3X4AVPsk7jb1yfy1aUFbkZWW404xnJYo9yMM1yOZYFfNRfDt17pGKLJr0SKX
SuFF+3sgQButGggnOU2V0HvDM0lgcyWFfB7Xzhe6HACQ508R+akTmfhceFSn
gXIcVP33Pu5m0azFHd3gn/z3iwgXuYdZf3XioQmwyrxmXEI+0ChgvFuerKOx
poeg6fL46LH7s6NLTB7+RhtKR0/HkIUHmKJV5KHhnk0YtnES6U7zfqvVp5qA
+qJK0m0N9eQoxZkE/PWqTtI+eYeaEzigYzKg2Dr8LiaFOouOsa4mX+Qc5xky
pCc92kgbXsgXcUkktPa9YFObX6/bu4sSlznTswJmKMbgI5kvSOZna6R/TpAT
UpWuQOgWXqIJVa/3aL9GWaLnJAZ/6MU6r9yHcezEGhiT6m9NZHgCiUOpI5nq
ijB4abTLX3+irReHyMJuWHX8iJjkxG3U5Q83wDo2I9HM4h7ayWOWlhi4mBhf
LxOCzmA54HFzdbk5W6Sm0b+HGH8wtS5Bl7iS5K+LHlgY92L5doMiHu9RLW5c
We6fRXtgZ9ACPd12OrcR8CgtCkt8/h8sqZ6Z7fq1rcbWznK2rW+o6jYsZR/J
nhwCcaXIyy6uojDgVhYZ8yjJj1cUBT/uPRkaQV3KmaM663cI2dB0XNlVRGBl
WAUJuK05IR7VCsh/SEBd2ilQzz/Y4NCU7l8X1COVLqZjS4Czgbps8fJJktxa
PL4AvH7Oct891ppp/bOKujBli1zp+LUV0OnUNNRgbWtcFElanBmUMMByfqAc
y8I05ONzttPMR+RINplrk5PhLzWGnqtixuyvxye6MDYzD5Zrh+rSkfmmBN57
jRBSugbME3FWdrSTb+D3I1LxB1FP8DFnGGTPEh28Zw3iql0HJc8ZseJlzWqn
9owdoRlYfd2CHZ4P+XpYyqMGIU1+4xMYXBUKM1idkK3G4ir+zd8GdfeOT5Pf
84jchwBFFdWCdtVRG/3FEje7URYUWlmGg7vPKaYjp5ROtSgsLIQOGYdL2qvk
lH7nV0W6REMGeJqUHfNsQAorzHunoD4oMBn/+jySJxPwCBsCyazTb1bn92qI
ErXCU5QFOTBD6fOuVXaxEoAGVUJ0V0CKZLlUfBDTEgKbASJW56fAZSZeOGAF
60P/As6g8IX+qk20VWxpX7ptf+mGq4Zm63/oZx72SnXW7g/LVureAP+nhBgJ
lsFmjhY2MMgPSCj8Gv5fD8iHb7Z7caH1TMf2gkslv94K8v6Gaw2NzOLyoOdX
FSds8OIQZ6tUQhKyzil8mXn5p/rgAwhOR7I92dSMLstW2yVcWCoK+wKyDqyW
2WsY/7WBim3090y0F1TjtWm13D/s7Desq4/x1ty4UWuwSrNQeFjNgU4IiMSI
FlQaPrK/SEus1aSVm15EpKWo4O0u9CZvObPL0Na8Ah0Rb5aQCq3dg4kM0LIM
y2GRRipsfb4aDEwNAsGeIDyrYWl4cKM5YoPC62UwDMbc8J4P0S+TfzJnJhrg
tgl2ukw3g2NnFGLb8rraXJYvHwl1tCEnUG9DmeWqXIy9aOEc7dEWnGERYqVV
3gaU78l6dcHTR6VeIDLMtC2N8Gcvk+GaQbz8A/D7FUqvukHqa9j5ER2brSFS
KoEQ4amfUeIbWTSajSRjNtjE8vSkRwBkD7UQx6bqEQILWEoJns86dwmJ9RQP
TXvJgBwkBZhXO2TBiJ6/cLgF+3Np5K48E/3FwR/t4G0GHW+aO1he5Mu6pwX9
qKcsPqDnQ/AgmX2NggmhK8CwzUT2KXe4VqxsS6lRQwrTL4FDYj+xJdcNhJ7Y
W4Qf8aUVmaV5s5P0zgt45aLK7sGOuZumM3g2J60eyn+273phJXv1BFp6KszU
ERxEA+JWTcHq03KoKfJxwKuCfDHXiuNdTz5rWHkesXgP2tCEjWQj1JiAJz1y
siW37mlpblQWwTg2HQaj7b4UPY2/yFieHutWPHdLPyWzatCT1F0A+i9yk2XQ
FZhZjWsqPRbVdtxjJAQht5CpUIhtIOsDEn+vojxsYuMnZyNDQb640XrGYWtk
V8ziC5RXD3WpGEeHWa4PgOCCDIpgQLUxyPed99Nz2faXQBiUE3BdF9AgMfGg
Vx8EXlhYtmQiX/q0k3Xgsg88E3HYBtsAO2uVUowHQ7cVtI2sYgsQ4lnaR7YO
oVCTgKWCxZHO8pc58o8JWIkzmtmqb7qWFgU5l2K83TS+IAh0w1wzx1Rd1Qws
CvbeOENyfLz1bBXLgMr8yMqZzIx72M/OtfSQq68nIoEQA0TBphAFFfB7jpM2
ey3i3594VLbflE21q7DhCcBz74WVhin0mOXoY7QjtVq6O+Q6xnlAlEOUY1tf
agSF304SGmftwcwjGs48XDHznbfNX30OvXHLNbleJqOwGhRSoY26QlZ+Wjwc
zY6lXBmWYvgirsFruWy2z7n2Lzs3xK/ox0C5KUSrsBMZM7m6Ldx2G+Bh3Q8s
RR/7BSmYZySEw/sF6wSrAfbzxuuJj0fM3Q9LJ+z/V7Rrsfi2d9mZhGAZMygt
lfr9zlS9tiDQcmfoh8k9jw5HuxNdTO4vnClv+gImrIHUoe7pkK9rgz3BaXSC
qCf1az8rXeUUnq6MBO46OFkccwrVzleiidbLUz8Jcj0SMHUSKDvMJLXdop2a
Nkzdpwsxxs0v5mzTVdp1SmW8n5hQjLskdflCQR+6VCqIANqrN43VrYa9D+Jv
ExvmMXWqjbK6e9nDGtUgur8kJBwv4DNeGjnxkvueGNylYfijyexbgL2Q4MH9
n7mTgtmArSBnxXYf7UY/MERbeFbjw+LZWdWq5YqkhVK+HVPMuPKE/OVU0Gjo
d0h1ixCcMUh7Rm+3GSPankWl8qJiEw4m+gtmmdICbtGgQQChN1rn9H091RIN
iRVpcP/dSCf3X0lFX7zUaWkFZhoUtgBsTZaFDLOfTUZ0uTFszRAeS6TdbqT5
Mk0X0n82xYY7NqsS82/1iza4JleO7X7vdrbQ5P6UHXn6TfIa1GxD36K/rxk5
uhZ9MYTK/zmPyDsYhx+8oycdJOIIlc5NdreOvmATZibxPfW1Wh83ze7kQcdu
J71BhCpFOZo33DdBXvCwJA1yStKKDJXcAeln9vHQARpQlaDcVsXMEGMc0Omz
7eiThzSlp2/S5LccbQ8rMATxInidijVxIVdj530WTANtmH4llpp0gd2rmsIj
4cvI+De3KR3XBzszbsT9qC1qKJP6nitUIg7qjLSV4YtQoO6nQKFTz0QOlBja
W6gIInTqt21C5SPqn8lkAXXoWxyWKxvvKe9u3xhZszJF3WtlwDjvC4Z6nej1
ry2ncbvP/BzdOqigrmOBvzd7vIV+1DyembV+gimlUFAW6dYb/kCSfUm4YEjL
EGq1l2pRaU2ocuAPAvWoFYu397CVuBa/Gyx69hNBk5WvCuhcYSho37Kb9C0E
fFY+xxLPS68UlGEbfcxkTDK1AK3MuziPssQn3BFoK28QOZaxHErD9p0cs2VM
JyXJgzFXUuaRohXYEwEPJ7SdIUwEkl3DGlGEiF1F/Bs/ESte4AEnrScbUr22
5NcIn5DVm0CYE6g3EcHMusuK/eeHtb5Bn2BwTJy8BnfG0a4+bO8gHhEvJv1s
50WPrVeXA5cwUQUUQVTlhFkPxc1SjOdZEffVu0ZN3sx5XyRHT6Tols3dNqiS
2j3G7aP9kNY4J5mNcnRbB3I3afqb81XDZY0CTrnPiRlhrsgqyeiW75YR3x3P
t2XB41PKqx91YbDihmRbCZq44wLQYdtSmFHqnkofOVKyFH2omiBogAnOal6v
uFleu5juH5tUCx12H1nKSEALp50wo+7mIB5vlEZ2MJl49W5AWsMAPdZhaxqC
Lh1ohSEC/DPYylXs2DCNTlILGIvhATJRW/XqrRU9QOq7y5TH0yJuxHrEHqRU
1L1SwQIAoFP4GaQ5GjVvBUHINpNQXOv6ArekP+9bESm4QQlX2qidmW+tRt2j
VbVyZPcI0Juz2u+RUX74ZOg0n7NLa50A17lr9OvA6ZPmbEcXJbLfLh0SEoaq
R7AAfNTVLFeZJJ+YC+y0OtXFjSlNVv98rUaJavWE4c2+Yri1WHvGVD6ohlkR
a/mMIUGicW+0whyKJSqMCm11zC50p/zcxc9SjhcjXsuDsBRwkbl7JrtEiZXd
cXDv3waDfGNZaCubLMuBPu8xDNHBjLuVbW6/Vn8DinmvHVqX6E9XCNGBFRJT
IEVqzuZun33E4G/cOvcCnrM2R6hdbxSn/bMGlg6Yp50wtqHpd5s/clELu87J
ZymTerLWH2csjXR6L0VljcDiECaFlEjLHOjzP6UdtxkVpJNshAU/TlyqHvDM
AjCeqOfJR13P74UfzFehMpfrDSJVeHiPbOx1bw7tKHvqwMfThw3Y1zt61uZT
eqYZQ8BUBJFvzTJbGkg+swtSB8CWBQ96OfndJBlcPOw/d16bzMLYSyPSCpm8
YLIF48XwJlPKaasHSg5ThgHG6SNba8RsQRsXRsF0xU/eeW/gpfqr/5enZir7
mQ/CF96iwckf/WMyvHQevgdvdcS5HiWjA5wPGMnHhoqE0gLB/icA/CYLWvUB
y+3R5TGGWuMPCZul8s8i3jcqIJT4XG0E3IxZVab5RVZogUHxwV1bdT1qYhob
SS9VPakrMBSJmE/50YR6x2jujTaouydinV+Y9E/3rMoVn4pwtnw8kyqU8q1m
/XCZ1eOPyOHWHXWngPFMgEOZueWerzFsTXuWEA73oNypq9El6w9kGL9qXp3M
CBD2uyAJgt9XmLnIEvB9o9+8nuWuPSkSk1jjq3C6fWpDoUKVdseZHKH8mwM7
ecePZ6ssuai6t2s9IpAPBefUhRfwuLVEY7t5pVacoXREmrOZ/MHM97K3gPDd
U/g2N2+7BcH8mAJRCgITtEA5hZyOYT81YbFNwemVTa6SVt7R/7egOB/7RGmt
XtnBy8ZD3QeNrz1Sv5pxP8Nz+4L5+qsI2mVrzOYnf9uGMkapSERDQWCfrXJw
kvrNbwHX7WUCjHgTePO9tvDldvaKizC273LxN7AaomBTHNvwcn9d2XKCO4Zt
ZMR7yW8P8CCZLhKt+KFYgU/WLf1Ihe37rZjQ8WazY5r4Tmym8kj5niv5x5BW
DvIeg6dBJY1tKSKT4vg69eD1sElvRfCEWRgPFXIcqwUgz/ZeNIl5zV3rxb2X
HIkM8KdIyU5F5nCSxWHTvsPSDEynHx107+3JRxp0FsLNuk5Q6EXNPzfjLqx0
RDvidyUSq429wwSN9hX7aJ2O/nD56ujo+SJ3OhzLvsT+vZLMm1iM+9SetMp1
WPX8+huvkh/3jMHEDGqHmw9qhEr+Ejed2Tvb2tFZOEQCdZTh2Pjt2E/iVXcs
M6ip43Qxi8/O2e4l/Y7Xn6qxGcrkOcrtx9JVcnvz3BvH3Op64/BuerXfgZ43
Qr4mLjcfMgd3QeFGv1Feuyq/AXlG58ONqwkE3gY5xoJAjp+bybzkCJioiDAM
ivuhSMWf/n3e+d5Uwh6cFRgAOC3mPG9QLPJ7KXAbcwIJ80vaM8ug3ap61o5J
FpXZcEcSEqE3Bp33z3zjWkg9k93XguxwMwZQIRGbJeKBicT9jdiF3T75CIsD
bcEfKD1FdJj4mbgynKl4Cv9M/ob5UgO/n7d6gBHWqWQoFAyl83/9FjggQ08O
ex4uOv2TiAZwBSI/ZMPI5r5051SFlvXYd8Xxcx9zNmsk4zAq7ZqWCydKmRcP
mq8KWtF13COMff1Si+s3iHqd1gjXx+wXeMKMo5R2jFCTCH7iEhdgsRukOECc
LqOtimkx1V/k/cViJPQE/j+byZA0LawCeXAGtwtda/2KngdfWsOLOeLy68/9
0gLIG2XgQV6MjN73x3cokiLWlyXJe4eLnOBoItmMvqeqr3VOgPoFiIXgQe5l
wyN34w6f4ZuDRf1dqbqXSSp6QsRUZ8hmid05sbYQT3H8PNwi0lJcIQBPnFpF
63Hoqhi3FKXv//wxUypsGXstQwKfuucCZgviQUjr+8T1/mGK7ty3GO2cYD0Z
FVdLArjCnjbG+fwcdurAl/yEVnXbaYogGm1+9RzcHi/Wn2pMnlVOAlXI/E/O
FjR+fQPr4rE8r46INad9BERoppl3hKS6MWNcHnZqaFBzaKIW/A0uTzz4hEfq
GVF87+23bb3TtzjMIl8a+1axLmD8uLOET1ggHW5512/ffcZ/ebwDU1RAh39a
F9+LjfqWlKVdicAh7nqWx4rgj6EL8es4xqqlGgGZwUSAmNPX66iws9Ex8/N7
tkjqMi0WQNXxzXt3EPFQhQc4ZCYns+8RyhB+ElxToKxWdZda4mfgPlE+7gO3
9RWsPNJQtNtHh8nlkV7Wf9bC3c3l4V8G1xkGRIm5zQwJ9dN7a5anWsvhirc+
UsVpyNBgcZNBGXzRVfu8y5oBibD0SeWrtuGAt77XE2ocR+iy/0ouj7mLZPY7
DXPj+qrXBd5nqrs0feHqoqM9DeWIA7hpZuWND3ptc+mPfnxffnvKHkI/YRii
XX2I1CqtovHWuJ/h34YWlqsi7glY8AMOF9UTrqzueNb56cRgAwQNEJ7ERjnQ
1Sv2fsMgQrM9JhTBlKXIujLL90iFdp2j9NgvLvUhbQ/sBvUi086T7YRm9xe5
A+xHqhChStg1fC1Fe/AfBIZ0WtdZmWcSiXF2HhXEF9/NQFHTGHc/FB3u9jF1
odSP6XNbhQnKzDyY+u9kq/bGGsVEqyc+vOytxiIbUeT0YeuA2jqWVtE1C06g
8OMN9przbeYBDLBMPhojmsfcfA3Yl57vkFMG7UKPnmYD4WniX9aX3beP95qn
HRMDDii7Hhqj5y0WrR1eFMM/L43LpTH/9vZt1m6eFj3or6AlBM44vfBNOZkR
nnvTs8b6l/EXIfn7wqgpndGjHzazCZdHN0zxNcQQ3X+XTjXVretAr9YIpx8V
qjy1DMDC+InyGhqbQQ87a+KAul8MFTS82iyst5m4MwMqkvKyJrzsHZNvbLeg
bjt1TVaRbLjRnC8BLC/wmf+RdUqTXm5YHLqv5p0CoR+qDUygXXSXoLqmnhJ4
eM6PSKriD8CSV+YyGYEuFfPb1ADiHbeMtWEyoXx9FsClFFffOlQ1UNyOnmyz
hyrLYrnpWp5G9rzvG5sruKUhwBI3AwnaF0+bdCSzMI2bSL8QtrZZRkEYVX7w
HHouxm8Zkkp2jumo0c1cjROXrmnGcrw2GFzuIwH6DGWaZ+UaAzr9PmxDzQUo
6ABx8wGvw++PG0em7iFkvrjwXtbGT5GD1zW3NcjDNF5IdDlzpnYQ2oJAQhni
31Qdw2zrP2OnU/x+4xp4cGceglAr9o83Jatr+0Df0IM31Z8/POoZr8DIEYhg
gj+LEsafAedZi69wXYqx1QRQ/3t8uGYwC0I+KT5OYtLiSQBWhe1Xh1bxuvos
JIIBX/ckPX+k36+hVqn0zOAimH+hhAc9aQ2+kfNzztOTMELeic1MACp/+iTI
x2tcq9cAma/JZlgfnA3RFteMvMMePmZzFNUHhbvl2Y0uE5pTGm3gawAu+TsS
LaJXBCtJf3CiKn+Wwekq+W/hiBDwb6/Vvw/yh5ExAYB7dEk6ge3kBKeawMk0
rskt5Qvh/i640ATgXMvyi3VXHpyeKjtafunGUh8gkfNlL/Zg12V0GViVWoch
pahQZiu8TPiB+sunNlY9LVDZ3WO+5reGqGlTh4TO97Zt95iDo6+WWO8ciRAU
ZXewWItTsigc+No9NxIgHTzcWC/L5abGVWTV8JtBEYc87mT+V6a9roOETInD
VirHMR0teSoaEuI/wOFGTBTMSRUT98ptTwAQYEpdHXEcw2Yjxu5/E5ngX0vz
tV8LkXEGGaSOiYkCsSfPXi3HIuPJ2KjD6e3b8VP7QAWiHF1IJBQFB88OujUz
EOfZ71VlYMR5JWwDj6aTPSBbWpE1NG5iJXRaMk6vAYkL85ZLTGgxBqTZOhYc
KGKyRzaSKLHzOtRN+4Un4iuGsdqZyp2CFZyJi4rBMFpYwHQsMk+XPwK2QGuG
W96SdPWuypV9rEtoiRL6ar1bvBNGfhq9pXH/RY+HLvzKhucWnPpPfZpivWzs
qsWP/SxT83SRipMwkuN7mZR7np0+5N3QItqEvLjYcE6yRKr/WToXERn2b94Y
3+4oHbske6KNhrI0RnoQqHhLcjEDe20nZSAjy7Pm/gFZ7s37VyRn38ejXGAX
1kGl0rE87haFkF8tvNzu1G2a/MbCb1xGcJaXsL5to1Jsa+suw7gU9GPF/KE4
USom7yRoKYlQQpiID74pZbwRahGulC8MivtnfVjeh3AP0i1ew67YIXuabiBs
ODRUjmvYfCWrJiB3XhKyVWE5FSG25IC6SQq94Z1hZDvpY2RMPqN5vFcWPBfz
ZGhKAaHBIstV7ZUmqJtg9zsHkq3a58BysyThlIeCEKLAJyvA56mWvjFWDyOf
s+F0EZ+cdLcjUqxm6xI+k+8WYRogwNC4PaKPv3ACW1Q6OY/voMwr4Wqoj9tz
mF8lELrFaqeUgdV085rp8iQiUTusu+UDn8okXoCYcakhbeU/qtVJl25X7CoA
7EB+TUb3h5obTrIMelakVhZg6/lSPknmjjANZ0EmcJYn/x1eTZbu9hYJFpXc
Jncst39+lRRaz+f+GQ38aDeQu2u57b4SxgaV2pP69YzyGaQTi2rIUcCfUUHN
AMClNfvAtJLbdvFKAWlxV1G7vEBL58A+mQXsdjHrRKSCBT5hmvT61Rfs1LWX
ZPuvEDqfPOT1JAjrwge2j3Llx7AsaNPKRY0Sj8UsS6odR+zlvu1EYru00+OF
W58wLoKt2B3XZr7vd9Uve3mX0x1oN6OVbnVa/FQrgr3oqa4N0Bar6luE86os
EW2bISFSvAotU8pJHA6qClRE3MFDYAPL7ENNRK7fllt+MeJpny5qiR7zuIi6
gWJlNoHGyvf6RI6YjUzLuBcwhZYXz64t6FHVILBQRSZl0IUn0G+qwWZtBk/U
sySQOWoaZHVIm/mypzJxt9ntRnbc/HGajWCDC7JsFQBPjKXJw0OG7kAfWylK
+J3u1+onMVH8FBdjKoKd2dzrBlB/s9UinTsjCzq0ST93rz1GW6O5/X1eqNhG
yZPqduxZVTufyEhAXOHWtiEJAw/jP0JsObR+UweW3DgIG6WCXcxLEjaXzgzq
+bDEfWih5ywFCphdVs+WLicsevgw2ux/rGY3qPjmRCTA1Gw65hHsMfaPxM98
Fjrf7p0WRRd0s4Vpg+Dm6CXcDhXZfaCbzPEUp+2M+oHxXdW8A34sz0HIJDD1
Sk38Z99vmd61ni2drsoXz1tK+CikbQP+l10PNxw0eWJWproEeU5dB228c216
+zYgZPKVPgXpHGReNHhxPR9OoIECfzIglaC3Q6QLmulIbDdMG4WYcreyod0Z
hWWriRdidyhO+dJM6krW5927ECci5iMpNu/WiiQ2eVZYdwZ3i8e2LcYh8qiv
Ome5EEbRzXbAmE6vdlCdMlnnTlcr4O57987wzBRxBKMMIb54WzTIeFDtLR+e
08epavV3CsfZtIQTcsU7pxVBeJflO36w+jfiXFdY6HoIUY2/Vvezz2+8uURA
yflpYArduQJpqU0IZVV/WB8OfKP5huj4ildeQBH+oH5ihMDBtreWy9xQQi8N
CBxyExTLJcmGFJYUqaKH8OaSiFhULL8Tyn6JXa0LqZx8SGZ4/FCjwfJnaoAL
VSg/S6OTJS4gZHz7/C156rwd6kXj+QgJSanvj+y6Asm0IseE0uHboFQqRmyG
D1PdlUl4uVUntfaid/M8ZQUcaz1J+YYLr58AY4OVDWJjWv0ocygHqE1xoIG7
6j2jxzWVciorNTJBQ4aROpzWPp5h62qJpX75V+EIUgDVUfsX6OK7KFWCOexH
YPzRnaLDRG6t4Dy5wYBsecnUL5cUBZSpjS1sAr12k4/C3CJJlZ3MBmXOP0mQ
+txxuY8jJJLjP1UMgf6ikWjvwwUmEt5sYF2/LYCp2q/5xC4H/EHuPruRRLR0
UNEUFrNYR5SM+uC2W1cQZUi5cSfWB0Jebe+cmnivrhmnlPV/PBt85Ym8+NE9
P2dv4ZkyAykq/H/jRQ/whbpGVFsqQ/PC/uQ/FFtdfFd1PADk5KX/gZcYDuF3
TX4YPs1X4DBYj933x/KlzsQ7fcSKpjGVWBsg4dfD6n0Hq83bUligdasBvTEl
1IGol5+OhsGZoXAyAhCXWhQSGkOm0ETYvkJspuXxir4TG7sDg8giZ0c3GaZP
tNdRMvSWbgOP6Ec8G3vvRNPZKw5Cxlo97x1IFHi1HoCwqYkkxIyCvqigz//e
4awfKq9C7ZC/HhLUCX97Rgltu5acq3JkoYM93/dYeju5ZqlilXj1m19KYW4+
wczDvTKPd6L/ko1aBZOpq+rbiwxOoYXGb5Rq8KrtEMYrLqTq34cp+jZBnudy
kI0xaKiqwoqd1mpRmhl3docN328D2ZxMCKxQhvGlP9SBXytij0Hbkrrsn/uv
Coonz+2TDWNY4eQp7E3Dc+74np/IWEiqY4rZuGAWPDawOWDICd7pknDvCOZf
bbM2Qg5WxMNlGMzJJn2AP0QFmNHTMuTWhmQPuZwghGAtsk19niQ5omKcW34p
WmV9ozoNHmwyKwY5gYWg9ZD58IPu/T6A3GFaoQPqG5xTIreZilTxMt5CWGp3
tOfcfaWJopUjSA7qBw4xC0j9RGMB2DRSSGpSuCH/sEYYF36CtmpkSrD37GAE
EeHRvRubLHn7+fU8HtMlbOCubhKW70YMvk4LwoeR6zH4trJUHLwc7AUUIy7K
GwayPrcgPBRmtsq1mKrKSvdS2L4v9St4M9EqnlV3juN3utcbmdJqr8fwG6f+
oTeOZLzWkeCUyLVqQ06ILXkJY4Ba6mymQRRjTd704aA02shEqGVOyv6OCmAR
t2jPhw0nGXnTkF2GvhtFUl70Dh+WDFriHfobzwcwxSVEg0NsOPlJ+8RXfCWR
cbsgCxtlhNa1yxhsMWn3oRwHcZNatJoBgXL5uSdgfQF10KjnBSq4WOBkZHtw
eKo6xPWAtexMNMeZ0cpszeohGuzEKCw2qbaFZe1OZ0yJakfq/LGs0dQxVFkF
WFy4RedGNfJv93LYpiFL4fWNGyotrSCTIOVgJ1WecUugs4o/k5F6NFT7GSMS
T94x4Ys2BRskEviebYbeTxg9ZrKeslefR+BBg+voVs/XBPf7M3m6+w+MDVp8
u6sj/NWGwISSxJvHBTC52UJcgosffWZqpNKd34awXCbmJhbxblBBIKkYj2b4
e9mT/oL4l3OaQINkO4QiojR2kkH/r7XmWnIcpf0yRz4cXKXX2UEGV95qsdZQ
SXnergHwQLAC5wgM/JqX4l42aUc2axBXmXtlx97cuiK4uAlpaSheLRIACuaY
YB+6LdZq0l2IEnM6DQ0rEB35wjx+XXa7+xoy18brET6bZCcWlfRR3rjBFrUW
J/P2/7psCJLz3FBkn26w2iQ+uMCh8BPsAH10G/Y2DNzyAsVJEIi1RkDn5rad
dDRCe4jUFrDIHKoiDtqLwNRsAXv+O0H7JAuKer7TDfSt6Y1+iTN48ld4L6oR
PfGh4Htykk3niRcnMojHnci1kJdchU8+F5bcHhCEDRARLMp5cJH/dOa8j6xd
VLG2sGAMneuIv2TVs+A215NDQ/JgkX+Pp9iG/Uu0/eIdx5Vf1UW3aFADa4qD
aaxT2/ZcrW4zKQuS8+QvM9bfCxQCGHelYjnWvthUE10wB7MRYBZP6gs0DDlW
HKpkiGAu1Ev+sjvX/QrjoObWikKT6KjqcpUVl5lJqSvk36diUBSHqfm8jrYt
YCQG1WJ1rpcfUlsFyfplvAyyL6ReM/hzLzEe5FF/jeC/pB1hGKUR7Ysm0aOU
c+6DTXyv7+/uJ+Kc273wYJmqwV9EO59gwcz4mgDMLzMSAVj3Bt3msTUz0p4Z
TK3R8xb02hCDeD++edOqCBCtkOl/4bhXVJRzo5IouWiO21gq0OnEMUBoBo7/
grvFndHXt6lN+gIAEzSbYPNikX0WyvoEa/9hKKl0SLWuLiApaXPS46UslhdK
EOEPKbvOIsvs2qbDT2lwlN2jRB1B6MNdad3G3iPNGHeHsfU3KcgeG8ONpnLH
gFCSor3pau0o5v1VX4EdcD80gjF9jopuD/BKzescuyHZs6R/RsgH5qp+8Emo
pI3ho2I2SIm7jjNDx08GHJsfHcjas1my1LQ7Ynctt//+JkatGmrdCkhuQbfX
spVLCDTmH3PWKnBZ79yRSulgOeSJ8zPGAP0vT+SxKRW3QE7JAWOJ4GZPj3Mn
qe4tKRR0rGcYSxP7GzkrWHQyv4Y2O+4QDiqPQmhqHLUhgh2mH+p2VXi3GWUm
BttAIXvzpYfSXnhtb+Ub+mFPGbUydCQe+PXOA+Vd91pKOn43eHQaSYX4iXo+
blhYTJ3/ITBObis7tevt031Ocj5hbKdW1nADb0dM9NQ0q8j5SiCpV/F4cNw1
Jla6IUgb4L/ZjQGVJxUZS9YiDH4V39GZoCInOy7td2w8UFtetE4fFMDoJz3q
FKsTGXq1pKoc+6eQ22t7Ip1P/e3yh9fsIqOvQVpY+hpOxOh8NiKMTeB4yoOc
Yi/eIuA1YwyERC9NBrI7LFNqFKNou2r0GS1/rL2j7UjU9b/kIH7U/AdPC4hc
d9/z54W9PNttgW1vlt/plBwe7HBfg+sg3rTDeXbt4g/yxGp/oFWLYxKQjojf
EYXJ7p3RJHLOwi4vNlqxF16lJqhp0FgqW/+cDgMomXw6MaruJpweqQnAwPit
keNRYVdgHee0yR+/aszwA+yq9MOOHUnNwFwB7zg+6YZ6E0hBoC5rtYyEpelA
dOCZLnclMhXt5ekhWEYrEW/w1DH7tZr49rQJe8+9jkkRCBJggjEQ8tc6pNUg
AYZq01pHeuKoeEw0P2PxtobffDAbGPmBW66LahRiXwc7jjyvwpRFO3U1k4/I
icnCRnuuopDf6Df/FsEpEDLdvfQrSvgi6ZFr++6bljca1SPiZMb8HXKe/Hpl
imw/aIapc7bsTe/OJ0v40zPWBd09wxKp6MsElvbQFBAJCt9nnmyrYG+ZkKCX
kgJxLFGCpo7BUgtund/JVEovHqHmpLOdb4xVsaVtBUmOE8O/JVHadNy2JWfv
NGt1y3K8ixNgkXiNt4TRHA/vuKXg46R4bwjOy6NSS48fE54SL+CcLfbJkjWc
BEeVINkU2XQBEFy0+1l3WsOOpKIlJWPgLKRwa4+x/KRx5JDbPFcVM39SuYwC
GhnYZXi5IEsO3p787ObuIvbGu1CZg+dzih5+p2HK0e6ahlSB4ZhlbfcyX33D
boDgp1T2E8RpCgMke2egwvV+j+H9Vf0nniT5R70ct3+pFH0vdNFRyfKznszN
8HdRYsJZ2ol7StIcIK+p6xsIDlSZer4CTz0apUkUbr3k+/AU0UstcaKwAbKb
IGmzY+2vi0FFAsST6jwBSswCq/rCTFOB33QqB9f+45YJIeEdElQhy2mGKe1T
W55OsUrsSV25ig+q5BV4Qm5RTxw3s507o0dHKqhDhha7E8LYdEnP7Uvi72za
bCuS71Oq2aX7uu8rvSWvZHO1CF2z8Z7jD4hajRJ2NNUBJrqqiIueRz7gzsI5
d3Frb6fX3uChw5sLJqs0usEPCSeY3v1G4bTRtb2g6MukzYVlcTKaDD4b4CHB
YkfpD+kFZT6lHOvOVBZXz4GYP8eeZj6YZB8Rh4IxiHO844wR6iZhZD9m4cdA
h4VOlpQevBr6GcfnKA6KqVzn6j0itMoS/HMHKPmTOr52h7XTeDp0lQtYnPOK
PO2VQnPjgNfTIWzKv4A/0Kn/IhhgxWVk8LemFLzmH6um+05kOH3KMpIU/4Oz
5jp5KA8opju04UZiO1zzgpUVRfoMTXw2XQlHmVqmQXwX8Or2K2jJHkbMQ7Oi
75GA+WRJ80ZewHzy/cPVh4DzlngV9MaYR/LSzkrCu1fsv/eC8qAz3IGX59dU
l35m+iIWjPjcBP5alVKOdO1fzcGhRkaHEUxzpMzzMHPmXoz5/bBLFKeV8wqk
OVxVND1oNB7Du7+ZAX/ffTQRpLldSFNVJSsqd/XmQ0V0EIrndXSuvD05GXbC
mGgEPaeTQWcPJJxCANuIiSf0mxXB0D2hOw5qD9FcqwuEp/Fhpj1jTbQeV4zW
KUWn7y3K6D106vHpyaU0U/TFkpH1WE0z/vf0rsP/QiPYMsgJ85q9PK5XRVHt
uLU132LtAW9Fgo9J4P5DGzSx+BRgW/qN1GhPud12UiamYPvu61j2LEp1OVKZ
onh4G+YZDjxbXuMNQEcfOAEqU30vEls9fNBTtQdrQlzPpBxwtqFEemZQyMZ+
fPFE6dT5d8yNwl27csW/lEJTrDI6YKBcHeDLV5hXuM46xYHJAH+pCQOiUW8o
rujHpfxcSvEp3gMf9FCTTAJHu6zMg3RWnQzNdKQOm8+snhJ9xzrdC+hF1ClL
9M88TZtjE2dv3gHNO+SYtqUxUTEvceelCsTbyRdG5bh+Vl0FTvXwYgAKdKQs
o2gwWD/1B5kWjXINFg78ryZY5k69kpairf0u1PLb03t6YR2E47bGdRzWT4vF
Hwv/zYlORtdj3zb5v9TRZutfN+l4StSaZ8nzT1EnrUGVXsHlmj9QL+Gujg1e
UqHpEUK3LFx5RL+4HY9mwFq5UIaJ5FM6yxdLaB4azRBfNU4xTpKPb1frCoCH
D+09rv0qeJpl46Or55ml7YVEbkpPZEvYp9cdHs/jEWnHW5AQEW39DAhKU4EK
Y8DipKPt5GsIOSGCUSxn1vjaZaEWnBmlH2DLLZj0BS+5I8c2fdt7VHEnNqnb
e23UyoL7r6TzHFyZWuFZxp+OeM/2cVI8yUKQZNYV2Hs2ax9XE0j9iD64f/pT
K7FHb9S26JjOetwtIt0n74OT8aoRIFdk/lifHgKE7BPcb0xpxxo0TlzSSNr4
cSksjUw+/C15M1iUjb7DK6HALFcxsIyhQBn+wZMThwURGlyEvqgatbuHnpLw
JdWZ9Osg4duJaZKid873Yt4aC6KAUl6rPzvsRzXmln86sgF2kebWurkHrhtI
361WoYsSNDhdmZdn0hJNMuqsjYNJH7YojFobLeHfOHURmoeFBuSqvvPfZwhY
zJkoF/ZM3ph5rHWB6ucws8NMaCLHlMJeczBmq4Tw1o9oqpv0Fyn18Ufqk5iJ
2X7s18PyuAl6Z+E4Phphc8fhY5F/WLf0//Br6lYB43Py7pFT/iXEmLt3YiBQ
knBjbh4nx9XBEHgK24b3TSWylxtievRGIBPgRGjqE+JiNwse3U8XaSK/Vvjz
ROkPVbbgppTl281QBeTJNovZp5eHRkpRA/x0ww55VCkJmSVVjEa+X0q1XqSv
HjhEtfIQ4zRu7Y4nb48hq8CF/Zmo3IwlM0q6AbKqLRaVzdyiBwq/ktCG0ZTH
M/hPWFZ7DjJJg3b8Zpo/f32QuSFJzEE3cEMEBaQiMzqTIHESQE/HQne6oQjI
cibF/CHGlzdycbuHC2SS2kya7oZTiV2R3pQ1V4BlbIHvR1aQ77XlUbkTHBo1
TltQ2bbhnrARsoThRf2HwW6h7KnJUAKHq3eG+bJrOmqiNv42OHk09HlPCZzy
IM0ODbhQvHNBrbGt+SCMrWaj3qPqQqIcZ3gJd1hqV48t8PLwGHSI5LoCt5zg
N53u3kI/bqjkZ5EWsL+3OSDQBQMzCcN/orTAhCxeIpuNBKVad47f4y3YJ0u2
x1tvNhsXWrAulbxKU8dvOxqzyjCSngln1Um2uLwYus7VrtreJhhWcQhbJasw
XZ5IobAvfH99QgYgsxF/2+AiwRp23g3EzPoGirYAc852GOJQXzjZTtWO8cwV
W18+nHF3AEfRvqkwoXtshW22H/HW1HF72yFh+K3crRZqSqA5+JmATgqOC1oF
Iq3lkReUVJXiCTbHrisl9i5d0XQqqAiXCOLqY56xagvIf5/cAbwYHlzJ4nxr
NkwQEEqBHtT77x5lXVaqcS4Hpv/LySM/IZUhxP937AwTnsogNcSS7aONcyOL
KiuoCVQ1cebmzgY/9mxU8Sf72hc950TMs2YdnkGUhomjbva6kuJEiz5y5M3a
TFBuNxmLX+9sFHdWwiFsGlpd6Xj+RcS2lXC8jnGvg8suUwlHm7tvBCNZrAXs
t8yUgAGdx8gUyOnTM3qfI05B++c+9BP+BBnpv6w4DvGVcCnWoiPkpuJ3IRUh
dmd34qShhaFWrmNC8W/irrj6CQozDhVLu6j2omz5k5lNZ8W1ZhVWdJ0f7XfF
sk2aH7iz24ClAcUUMK+E2Kf98w1RI+ZuDjh18KEP1ptFIGrgZdrALOOYTWFb
wcSGS5HDg0XoqI5hcT4Mp9j/9v8qH+ADdSqq2WeO27qYoD3vN74P09LbaY0I
Uuvq4azCp1VoVQleutOcGVW25BWbUpI/D+Bo/iC1WTx8QiodChtl+EtsP7M5
c1VC6moMcQnt9qn5tRmVf1dfjyBgWpTt8nmr3o3+aKglqjBgxeeIfLeWP1K8
3sGbLRDm73WKFOZHM4wUrTPSr9+AQCIx52fmR2Ye5anTFduA4wF+ScH89HQp
YBj4n7DPNvipTx/ayumRLXD3u01JygN03WHAeKorXqWJkC1ua48ypTJuoXn1
ZoTJF/hT0y0sEntVWkmSKsrSCz4S33LUMucczG8+qcqFNfrJeA/NTfxDF5Su
HLGyPcWhK5PlR3w3YPTUgr9ZryT4zIvugUg8fgDE4uqS/3ZjR7FuS1GYSBdh
ot+pG4FpcazLkAtwYl899dSxGcokc4Htc3L63fl3GN50Cv7+HHEPPpZCNoaO
jMQk3MQpfL0WNAiHRqlEWnxm6R98VDEjIAVFu5t+GhdhxfFoioc1sEPl12Lz
dTWj1wySh7W4Qi7hS9JM3amjtoipPmnpTabxQokFiqCbBr84IDanBQ5rwsIc
ptS23dYTB+0tjPMLqc6D2Ym4uohlVA69zg5iWPNgt2Gn5iJCSoDT0CSlBebG
9SBhqCMJyxazVxW06L25s3BRCOcS4FiIDHNtseO8D7a27NGSEGnGN74XZMgn
H0N4/wcck0LIIV7p6812VCX8piaLPQOT/+NVnPSibN+PM+6YL17WD5mMVGA0
uMscibXYHJYS4yCdIYl2HEr1QvRPbyoHwC5d+adb9iyl+ATarO59KVZIMTXw
7Ox/2mc9E1k0D9LH8hJHJ74TRvko9XNJb6he9iSBd+YwxcPXZUe8SoelmrTk
ra0jDzDzjqH+TYv3U4/CNd7mIi/ExA1+o8rbx6IZCSs3jzXf9LLyGfuWVsAY
VRoHcU10FUCWuxau2MnjYC/NSz/0KXTBaVqB+F2+cPElcKpxdgxRn06PNlJn
VPDIvC1SbcS5mF/RQgi1VpPzriTRAm7duW7h/ATlvVE+h+x9m5cTIDQF7ySE
J5U9A0JN8q6xsHK/6Fx3aKVFpbmJnZ/5buPoaM/foFmyo+q9xhSzLsjOExGA
PVEbmfu3WppBKBwRTDijie6BHfCgUUKG7lw4kXKdvqIrT2edXkojWsWkTR8V
UvBFR+NyLBDpPEFXaS9T8x1ofUwxwt2aAyn05pAJP/aTgWSc1eYO8RZ9Au58
qTIbzxSEA7Mw4rgLbW1xde8HxDZg1gCulAwRz2E2mf72v2+35lWOHc6AgVHt
V3dCRLi6V5BEw/29ZGXH6tL4U2kDgttudLtvxGcEXybFA0wG28mT8ZdePmY1
O2fkA+uXuQC2+EZjdy0oZFeg1R79YS2/AmYeuFysmBYCxn1Y0clYkrwcLW+p
GR4qR5Fju4oHl3Avmw4/AsaFFlf65aI4/xKCVzpqETR8vAw5IKnMLN9mIlMl
gP1eJ3jaDjzYjm6cvhi1Rb55owbQMOTVD9KStb1suQn6feYjClTI/CExAPUb
hqD+KgrXdCeFf/Kvv4fSjCLdhfJ+cPZDILWRl7TFEd+eb/iKQnQteQP42KQI
lIqnLCYxcDjh0BfKRZBs4tH6QeNosOv9218O0vkMHjeOLJjI4/oTusAsjisH
SWNCDLb/fci8JTx9UPplCUeOmhykwH488Mx77EihTVO902VW9m8538dLUEZo
jfHG+HtqLSHycFiwDLH89P++WPH4dvqyaxuZmDDoy5elvHBz/9MUccmLBIT6
SOjmA1lpUes6BfoHvO9RPPAki/gYrHMP5bUU34YrakGRl7M+w2LCAJJEiCP2
FQxf7OyYbwczy0OR0TM0QO0FnCCPiVbONdX08qpLbvYlyu81SYzTq+ZzSm9d
2F6lK2kSzpEWnaGMW/4mJfom1yp7oVyDOxnnXC6KYNGs2wabv0jq0QXw4lKC
1xDWn149MskBFcv5laPMtPC7xhG0Tyi4igGSsG4UgbCivOgKrTjS2xptjWlf
kIHHiv18WKjG9Jf45kAUmFYomQOvLLi2mpXOnH5Z+J+Xb3wcFcFxPpHMOTyg
XDSa2qhzfrBUs9mrRtMXgmzzyyXnMpTuKk/4taG8vuZ4SU1EebG4bCMK3as3
asLiNXTysQ8Ykj+aZNzFrJd67bEPb0wMiIw7lf1UyZMFwNIY+LSF3whUJrIE
ym/q44u9f/Q5hGlwqZVXEz80+oBJwEP2vpmdzetNLcJ1ph3Qmq5EtSKGyI2P
jTahN7Qyecoifp1tnTe2+lu+OArUqoxNcahUwvkeCquWEv2Ay4YglfiWNzwp
rkQF4YKT9LHuSaHlUQ8zRvFkFsQpcRoLZfULtbNVLuEVV2yPH4lrn3v1py40
Y2y1qK94jftHn8TJG/YkMA5+H7EBDBhn2A2sKgVX72q7LzxNIURs8QZEPuXM
PTByBuGVpbAyZaV7B8v6CH92w/SwLkDGjqum9WB9ysIaIkK+ALeptBQlEfLs
BFqMhRQjJPwgYM6DvtzY5cE5IoSqe2IWqrshaB5L59RcwHi2rYqyS/goyrzW
iDeGWJjKuLn4fhGTlIClpemxVLODywbV1h+8Ebi6ukmBKbwTIvT6roWvlBHC
qKnZwq6d2Pkfzeej4MuZDXEaq70qxOsRjrFYeuShf8S/vFaya4CSUiM1HocQ
c3vyq3Ai7rUCQYGTMfILPEzS45Imtr9HOIHdYiu19SpPwyQHVxoeK9iCR9lp
1Y+DGm9ZsWMBzlntsUiCmvvvgk7LCydd3OiJFb2pQUIu2ecHfEmPsuQdVpb/
TyNFI7BnaZRXmpenyVwo8tj/XzvLVIL6ArP9NevJLf/LTU33YMkiIHgKWrQ3
yiQx+CWLsr5cyNPhYsOV/jM2KK4zH2OzDO4ejJMhDGjCExG+Fz/+as02+pHA
xixTshzu0GWJhLeQUdT0rVfEvWlpsiZrtyKLBs5NrTma/VQtsDposnsaEZ5z
K6xjn3Z5TQmZGFq6P/s0Z0dlXuwDQ7g976/6SFxi79TtCgSJy3xY9O+Gydq0
60Lvqd9gNIHJsJ/qEGuFJ+zbYOtIxQB72ybA5g8J8PN6hvFmX9sDzMD/DX9z
s/Gqxa+EznpvkMaD6/Zc4PqAyOhmxGi4vBI3HlD33wr4FiOC3cHmcKjlSyj0
QCJszBKLx87lbMzAx9ciFCNv8HhDGzVvlFiVARo91GTse4VHbycJkjJMWlAE
XkwO8lQDWOY6Gi+uvRcCrtG4TePvWAW/yS0mJGV3wN/w83kkZcVBot88oU65
EPKTL0j7uSG5FfNxtdvQxEZBZ/8R6yXkHfl4gqXpCfyK7LlhXbzwrz0qiJQf
tEkhUKc7GYL3xi7R9vCcsLADJTvgdqDtoGtXG9cnu5Ik0RJHdGwzuvxGin9s
O+B7fF+LpBaT9aBwRQu3zK8V5BGXOoRpNCyU9MWe74P+zYd4tDrtLNVVsSX/
hmYGLYCwe1yctow8IHJeuMg0eiBFeWpZNiOfwHlAXgOH0OM/gKxf1TjHgpkO
/uSOGG/n1XDJUJHNwYC+QIGn+tcX+YILva7F+J5Cr1kFcS7beNw2Nt+gyiXm
bMkVu/mI31iYHwSog9PQ2EP2byTDhU1AN/zpLbxK1y+HPAOYBxC1FTAg27/7
USpunGfgSP9G2lLEsDQ9z86RHMBG8/WHV7GoohyQNxwHXjZGFvhyeloYW6Dn
zR17gsHpVvRLUvfYZ1ViRPhQs2zzdWWWWcoW30vvYzjWrGCXr+1Qyllch1K3
WxLEGwgUo3yMLXnIROdPKJO9ww2CJdl1w3gzx9vcN5hfuw7hDuFp24kEofGm
8Y1Jww0MZj4pwIUD6tqdaEbVU1zmKix/tSe+yRCMA8jiw50ByWzy1hJYm9wj
2RPc1FslisQ0UX/tFOvdSuZ9FUuzScZ9hI8b/7NLMxVKvMJ+qRtMkR7VCzQw
94BbJQ63zyMgN8s1OpbtWTakSe5Fzh71w05slgGnXKv6doUt7ll/Ln54ju2h
RmK5u7kMSetARlDlWBe//KOd9FelWHZU9d4fJlbquRtzoo3+wMtz3bdJz3VP
9Q5mwji588jKF5IFSLyucsl4sjNrW121zeBoJx+xHSot8B+tF+lACNS6D553
6+GM2vVaMZOuSQDHIASXOCKfUlAQdH/fwtmEEfiSHVigw9yC5ljM/8XgHrMV
WwNZVuNSKERdLqAUjMQMZ0654DqXMq9CUzx0dKakUWu89ZjxukHckQtGGcDe
32wNJSeFVTKna7duxCxJeejgQ9JVfREMnnwYE/AVudMbixRsalUco7o7tsvM
M/DJytomDoGlsYWoZ0OKouePpv9KpkZglDxELMjXy8aLmAQBRQ/Y28Y2fvjU
dVLSjQAkj6KEB/DPMz4eniCvGF7MEtyxQSCFicdrsv+0JJZcO5OHyb/565h6
IwsWWnJANTgAu3qKwRhH27jYY5y/77kyYPoiSqw9mGcGTe35zJ9Nwg2OeD7c
FO3dpsIaMAlYVtjM7J8BpSPVJQf4M+Pbn3Nv7+j1Aaakd76NXzcnw8/dFZe8
wvdAcAsWA5ufi22w92HEPCwQ0JVcbXgjNhttMTfEPhBZtMYeJm+bNJ28ICec
aIPhpO2yilYbCCzxOXDUWf0Xy+6OY4l0M67H2N9eM5QlzQjM+f+Q6I/HMWTR
mj9V+oNsks2hKvP+s6htB4Cwpbh01Ke5HhQ3SvygLbEmjghY6VWQ8BJbcLoL
wakt3a1VznCu5Cbv5ryvI95nYEJMwrOzggBT0dZbmspibJ6NBOANhx4nlbwU
RVAXuoTIJ3spXN2rRJxyJj+lT3xwFC5kfMcppyWO84kea789Xn9IODkkfLKm
3hj3b6z9KurzMx0rjpb/jJUVNPVGmjRqPdq+BR6T+yp1g1ryPK1Zh4QmRtJ3
LCQOLUSYZeXmNat8SP9NG+vfO55/hn5bP2yHdXgjhkY+JAOlkEQNiiw+kNuJ
NAejDnBXOn4PGU+L1xanCDNLqlX7lLAeODnuudWUMqE1yFGT4dxzi/haN9ck
hk7Rvi5xF1Nv4WY935VnenGcwJZr6BsMeD5zvf1tkqsHgxy4hmxezHseSg7k
i2aPSZOLFFJjOQXBmY0NkTYg8YIiJttjxemgotIO183BrW3U22uke45vAO/E
7dchgX550HRW1agWBUDMi9rvFS/YGwuGv4ypUgCp1gPCZddEuzVY5Mq6itwG
FaJ9W85/dSK8IIYacuo60GHbDy4RYYB9km3HvzVebVUUXNNOJzFffVuCDlGV
wIZ3IdFrZTSwNfWUsv/pCNHy9z5xXR33QSq6VQpR5bbU2wmQ2IXIOCJ5r+pY
QzIoaxZNpcB+Ncmk+Gvl2TvcGVP+gjYu+L2vikOzysvTSmfUrHXAXNs6CQWe
oZegTVKl1zwyb/V2YlI7OWn13Sx5WJZRYvmn/MnPudFuVkPDmtUaSbSJQK2M
azt45OHKVe/KFfku3MJa11HhiBCpFbKoDkM0O3v5/sMwOIcaq5iO5Yp8r1ev
r2OPWUgmG9191Jv9BuDNByi+1THoB8zy4qoRBsb6bu0viJ+aBnpooBhRiKl5
lPn/ef0eWkLOO3vBGvd7DDWX/j9Y8rFs13Ed9hCrlRjPiTCwpP/O+tE6RzEA
dtytqzdK2KJsjWvIZpzNdG2NEwNQYI/VutIE3JRbw8iaPmCId0EQOeg6s9jn
9HBGBq1+2Hj+0AsvrJ6WitZvEerAXeSQIWvzUBDE0elbDHYM3USCaZaLD6QC
/a1MPbKDk4Q01e6k48DTMFOq9N47oim3pbzaqC7RglpSucuY9brpOTkxwXlh
07XJTvyUzA6qfHXa8nvzwcDjS8vNSfVky+FtTeU8ZOoV7n2GJld0nHgvwKLh
tjhh6G6SBoRe4ckIjQ7yB1x5ZgqgnBXTl04s0Dwdx3WwyrCbBAVtIwVpXU5y
7uOz+ep6terR9ZaFz3kkc84Fx2G7rGg80Jy/AI0Hr22xM7CO/kjnHb537ZuP
h0q15ZKn+ZZD5nvFduvgiAogRHGa48IfEaGP61Gfb0kgHMArUHbjhvC0mDs2
dfQU9HxAvhB+91nV/BI+NBt7759XS3IwyQvXSbyLay7wMAWCPOOvXX2wF0eq
4w+AT2hUQG/aVuduXitk8+Tq1l/A+mqE/QtyxCFkz+soQEikUBZEaEZWSS0D
/LW+WvzCy8Lg3tRtHu7fuqOENdxCIip0fv/OMF88d+gMBnLBMrtuu1UmSP68
jO/ZTaR2rOs+uX/ytS6+nN9M482AX7mnkYcJgwVXfINDbm5uCOmnmZmsAo3+
jXzR9RChU1PcmfnlRu93gGZEl+weABFDDawE0rvpaPopBO/yOFI9lawSitRT
4HDZEYv0qxVz2XTw69tzGgplD0I2ZWy2MAtmg9ZrDN/jg9vNv5yq9QXnhkjg
iIJtgwSqkiMY84AEda/5X0WjfO6dsnYKpGZNO7OMYc3ZoYI2j5Nsx1sFJxiy
4ois1UYMC5C2fuf0iaqLV3l8eIDMn4P9xZ5Pc4MKKfyySJxMNUKfvekeXcQ8
fx/A0BI9/R2bmpcIhEqqKL3HoK704uzD+vrsoohfzuMoSl919F3jXzuGTOeO
MiIBr6WgJYQi6YSqnBCHHAwrphYFqwSQy33QSb50uN6hOUSKnQs8/mI0RJcJ
5WR7HrgwGOCwnsVqWUx7Cd2mavlc0kM4/jQ35DWSFvAtUtYrNWc5WKki5SLd
Tjl1a6ABiwT+9SqP+BqrQhOzJ0F1jJ3SCrOWLt+Q6uuzFXY4p8yMB1FZjpZY
9bj+OzSVgxdmbr4sXC6CVXizyFpOQ4Gicm0Z5yTAjUpXRe4VsU6gzC1lVZcX
dUF3YBqE1aElIPhoSI8hpzM1rSnks2UOWa9K5UXrlKUt6RaHLLQ+5GJcFkiI
CWgeI0Cnr/bRPmbCsxI9OrZZcZciA7FEokchTHTetxxb5Qh3aPWXEuzXVjWT
MHzM6L1v48F5TRLzZbzhgWYvpNzoc0B/01R1SD3EL1i9Bno8XtOzegtfC+Ji
vkG2RyBSME4XOxJY6qAv9z7uvxevebumdlAJCvihD99/1fSAv2PrSTedImpm
VA8Igj2ylSAdM67Zv2Vy/oGvGiuCxl58i/b86RLU5RZD73M76c6TeFx0az7E
3AcNxb0RlJ5e+EvRVK0DMkUKRxjvbdeKgxoAnSM5covP+Z8aOksaXrDGCdGp
/gkubhtQjRuU5mUT1mfK2IS2yCVWk/LPfE5YE2AJkcOVKbZB239+EtB+tABV
cYEsbF5W2oSnqIQA5O7e6d/uusuO3VhHfWrZEgMGrfpN0/E03NY7DDELjg9C
Pqi3Cyo581WPGEpgu03QUvUWHHbpiW4te/eZQvUEc4WxnGN68lRODDnrezkP
H3R4LcNp0wtMkA9xiYMWDMi+wSkCW7YcjnEefTzMRE7c36DQhHWeIwJdKyXY
XXYBZADvDc4bCiIw/3C/ziQc7sYQhGgGmei49vb7VMt/a2h9WN9ViqLzUnKu
ZWo91jPJPNUmx/Eg/rYT6cbjEgfK5+U8mztuB/+ZMRKf32ccDfNnMa7+ZSw6
pD5NSr+ij+4vk42xSxkb++KYUSi9rKvcNmYCsSMwilsBRCQlD49alhwNRtEy
/iJX6MZRRHsagJUf3tCjONGEX5RgEixaInfmHj9dDsh+LyhvDGnxUGUYi0Mb
oN29YO7oQYhNqEM/ZjB31PMLhst4acslS21rimA/8odltH3BXT1GIn7Z/w23
NyWOZ6Ir8b9uOWBBeJ8/1lOXOJBvvEeABG0uuIHh2yyLkdtKHg090CiMj0kp
J8TQnZbZr1aaYz8gQjQc1dga2aVvbION2gw6DwFOPnf7GciWrwbRk/UCZhP9
K8i8mZBNZ808zx1U2D6xIZY4//uC/Cc0PklyU+ZLz8IZLf5uuAdgW6RLoJ61
XDRa+UHvA7uHPJYhZ0F4hcM8Hso246MYMCHue8i+LIIBhnQExU17y8I8A869
hxslOodPz0NdQg7Cc33EyGHrR8xB8LsDxjl4GeN9BqZSdXcOowcKsPaF/Tg3
2I7hFf9uIWixZ5EhhzonrbY3nkIKqGcIh8NaGc2nzVRNR4Hz4M8kJdOipqqB
15YOPHZOJdf3CSN6ViGgLJAxrWqwS4IrCiHsU/0hjLH0MNnGIbHJWLMXg/dm
X90nfNDM2HHHvkuei8itdt1wn2nMCDsdqCorq3L1yTHieEp1v4fmHPClsOV8
RyVx3Crd592Yo/6PtP7VPH5eSDExLlQh+ikXpmrk7t+F0m+/NJATVAW2t2/3
h5Z0RgRAPyhD0jevGKYUyuY06oWTw0DZVpSMy1Ktsx7qNP6cAPLNfdW/BrBd
LOSm8Ml8CMMTod9QtkoTnpvNXewdXFKvckSHMmiwhgnjGqTMyp5aytqf7Fl+
RqDeNMPzYwzu/i0+09mB0qvfbZ91YgrCYlUvJbJhX9puXEdEgvTPaeSwof99
2DNRf/sRacMnSGSV+NdE5M7bSL6ZAsW127u3FMLn2nQbuhJvMaftnmNzs8BQ
WvHD2QKQ/p67Mkfkw9D3cVHXKcsGlvBq7uC9LgfnZgJ05MamLoT3JC3Pq77V
E5AA7GatmHC/i1NB6Pux1H/YzsjuVYBRuzuwCvkvt9vzmMG932xJatQcMEhK
xRlyvRFfh1KUoV9bkMLXQgpTCLFASQ+N8uYaeKRiElCOLfA+xd+XpUxA0r6s
ctGlFRYzM+bfUnlOgxXWAejDnlH+XZcChJBsvC4UFSzw8iyp8Ob9IMEmrlHx
DuEiT3ptSsLFUvV3V4HSbTJCu1peMGIqPG5o6q8+oWhitFBBkZj+ePiT0013
6cKEGzzao2ZB8P7ucoqw+iYRmEpBkPYnHC5l5TC4yeQvBZzrVhtU96UeHPKp
vRCe3fy/CkDzOBAfs347TbUspbL63VeIVOKoddZy92Aft1HTXIrk7kVUbO0A
WeIGnk88rivOW4peAH04JL2k4Ce6rB/SlXXx539xhyQap4KhzIxXxGSlI1/M
6QOTbkaIdQyF6ofQwFLLWg2EG4Vmod4RMIE5Qhw8UTXd1RplGMN+4E47q4hn
OywzOKP/jdm7pRcmKvVgDLcFx0DeT8okmaRCjy2h/OmsJ8NzJDDgVh+ISVUd
EIaYB5QwywgIUcC7R55rwfLzO1/FXriqXw82nGTSRemL+rG/KWEDXsK3FaUG
toNHQC9EOEsl90h42hJ0UBPWUf+j6n4aBc6IZOsjmJtNiTth3jYOAbAP0lGT
nDmVo1zv1VHZYOd0+ITpiU3PddIGgPtr48FnkHylxccTPg6tCrsr5IYnv6Kv
R9wxtKujstXMsdh9yS4sNjSXlIpXH1khD8Cq+6pxjM5gHt5w7Z8HUkdbJLB0
tghO+uO/n+9Yf8KtvGRPkSxyuc74HSlEvsuH5gfk0CmLAMwwM8tWFazIiUfW
DsUNQQIDCo3bVn5rxrSvXR60b+/aylYDpksnjzz8Wy//OyPIOideh3BMqttd
qDINC209J1Y/m22q5l72liZ05OVJlismvXfRG3B6oqUvOMUvU0A/9+VOdKO0
/MbNsqpw2v704+JwVKhvU2MbVGOsnbkW/V1k+Ef67d3IVRbpcLHcZmAs/6kB
cBrI/wonIzqCf03NvNHncPkT6HdWIk8yQMP0S5M/KBvVCVdqiaWmaiFpKstV
d+KNzfkpHhW4lPlEhtJvSlQ2XXv2KvM4sV44ypOPTB11ZTDqEboRpIkaHPOb
Z+Js0lUW9pFMy/dqnL7tIQrqk8rzuWl36leYyy43gBS5esH38bLWdqWxuvz9
T1Jqvy6eZg0yEtMcJn2CCEWMp5/hODGUdiUan6wBDnctHc5jQsTLp7QBRq8E
WsV1YPqvmKPSZcpf0rnMv489d/dmMOE7GIoeOLpVoad4o8v9RCB/hXQ2biGe
ThFBHJefiHcuV7cXxWz0tuyI1KvDWFWl7+gftbPczoGIaaGQw9UBV1ovvQTI
v4+8hh5qnQpYDS5YkyOKzQUwXeWfFUzjndj6tjcsspMmuRDo5BoUW0cRd4Sk
FA43K6wZR5KUxdGGTBbf6UbpUh4Ni1sNPwCpzfNc/AyeyZvaEt+oY2yXJ5wA
DgTf0/BJByOI99KuNV1SeBKlTs0RnfwxVDoznPEnXIUUBbIU0GbP52i0/Aan
Rvv57p5IIPjoHfNQcTKcRYV3aUFjzYdjk5fnyZsg/xMfoWPac8J2AaLhP0OP
mD0AvPtQnV5jeBScMRL0eKS+uBrOUXJPH2+6ZLEmFmm6chYNxLN21Zk54nJ7
K0/V8BqueYkcG/gu2k9cebb5YXNVSUSaJpXE4R1doOqx7ipYkgWISdJYBkXd
uocWkNVI7E634vRVrb1LdIoeTONvBwXYIJtu9uxl/wi3judy+a0tfb07Yegg
u4cPyFCz3NHYQHd8QsMblC+iplsBqUK9jbsIYk/uVkryTlZMi4/2dBRTB3fN
/BhQ+NAbJsDAtIiqaom8Gm9mKv04HrzpsKEHMNXonV1R03BMLcdp1rmdpGvV
PuCsxxuDPbcCF+mYrn8JX0Rdq66+zxkZmEJUX4SNMzMQoceJMB4GUo0qiU7S
RWP4Z/+HYEPriugl0Tk1ltldRBKZClVzIt7OVAAjBm5GGOdathyUeDjOjzhT
FJQOrpyRVXRdvwR6ULs5tTKQDMDU7M+HEqWr4xpHyzFdhv1MdidBbX/Sb8cq
zRJsZUuV3BYlyoAlIoqS1AalQJs9YTQUX6VM6Po1CNlwN95b9E6Y9fawmx5J
u9p26IKTraCx9jOA7z57+ZD57JoEpQn+L795iEui6Z3ZfpMRkNOPDzWTPRfy
SpiTKRTrDlq8BGde0vT2I7cZSjnKyYI8VzEJnilma+N6bi31cNZBYzdPckh6
AfaPndpPzUL1Un3TFGWsAMUZTEBjQwjwHmQxo9V6Uw/vijznXPTA//3pmpTp
u0bIuWhGNdpy7cGghmgNlnTNxQ1XP9iKIlZBFv+L0Guod7I882iX7LQPdCx8
yNGksTxTNP5QwQtmy6uytnNTqyWF7txC8bPBF3ZmmtiwspwmGpNSP06S54Ay
HgwWJ+SwMQRDblzu4CAGm3tFCXks+RkR9OisE9HmMol34DM42zYk35osF1Qq
BBJtBNTB23hSgCrNYwzTrAXX+FDfbOYyTAMFhW4wDO1qQq7w/VXgNnf9SVa3
snehj67oCAbSlPiwleV7idIGq1CvRWmQp10EGlf6lotjLBEAmx+iZy0gMtt+
1VKFdBrOnrlBZlEApE1Ld/5E7slq3gtjvwEFlW9rBax44ak4q2e6kamj52ho
bAfI2mmqrE+qVUre4kq/jYQGWfSPNVMUH8XfJFqAktgiCAnH6Hs3HYRo6VJm
mVeO5m9T0bTw3XARRKSXhh9X9dSx9d6o5NShSUp3DV5KKgufE/sFENvKieel
3iMbprrNr8JXKFtLQBCEm79zbq+RPSlgREX3nTA1y0VntJ2JSdfSBsGdgFx4
5j5mkRqxB7uB9JFCah6kXODIvVBv8DbI5RjPGxDTAL0je/EStJrMoVCR0DtC
s0+SbnmStAUy3SOYMRaiTNLB1fc9v1fHFIsCnffR69+tCcAwYFp4DovW2+qw
4J3qYsPcY1o9ivphsVrzMq/18yD9aHqSozmY8o+W91xp8qd/0bFKjRq5mKQl
ald6fYWVluNMsjI+UGWjbOwVj0NaAm6JDXU33UoKrP5OfKsTuKVMutdsdVKt
iV6g3PlHOXLuYuu2VGgiY2qtta7n1IcKYkmze9IYxR9MI3tANTzVAb5zkaL1
3kFHdU7xi8qIBQVuWh+c0Br6G5/Vmmwb3UFjhGUzPUfJVa5SZeghosTHiN0y
qxJwRsxKnJEw/4CmUS1EZjDpOtFdwFMoUBw6aLjckb7oFIcxGiuZcz3AbHhZ
/JPb0vbYv50KDHYn1qBFPKOjTj0LEw2Odq46f3c89/42oLl02+ncfsbFp9oA
bjcLta8mv9jkfCSHYiLBA2BTrmNOC3eLkpa5ytPfxP/75bNcSDIArwlIwxG5
zWT9UVDGkWe0PN6TZAgWr1T/SxR6WqRbxwnOLlv3WKdPfHb/Kq1lbkMdsT8t
H8bc6dZMGNTY/NjcdYVwJD5HQtuNXycNs1tVC3sEuSL8lmsTN96A/T05puSc
4Syx5M2ZNOkFTls7aVsUji0Z787RnBrXgSW9Nn/8WBIKoyYZZQH/AlQFFIhc
twkHAWGBQTTkksJ5k1zSiDJ5dFbYmxlBfYPUeooId8aLvBKosSJ3put70Ft0
iaZKcMJaEC9ZBGcEzqb8cUFZLwBgY8f1qU7UKgjANL3qVdeA0U4hjJsd9a+G
pjRYXtIrqxRAuQH8VTyH7tb/oT/CJIyyQEnj7jNVSGIx+f7PDXscN6ThVi59
zHnRpOFrs75y4xIvBDIOuWL9yapUxIxXzy/LVaXY8Cfge/chz0K30gnBCnzB
gMfCMD404B3CTxh4W6uE8BsWjyziLThvjo+miRXi8y5Bi9Y1iFZJunMoBtyq
XqHw+wPV0C0pIzVrNDG7SCzDwDC3iPzEdF1BIZ35jBM0G4Pdeq0U2DXvfJcE
/iE2RiQ7n3MhZ4VYDfY9aB4z1jg5LcWf0LCvbvfrtsisMbeCjbFa38FEthZm
jWUchmL8wvCsaUNAt/MHu5GOpCK328PoBF4/+tR1xGGyvZt1kJHGe7VUa7YL
XNI+ERBVHcYMHf779SZxSqI7qocqvV08oKhJ30B4BONAQLZMWzl7t4W4t6jF
y/Hp2uN+PlYOgaYFMNA3nhH+bD6MSQDK+C58tZjZo0lKSq1G2bu8+VdLJuBl
dUpV8g/+KFlZ6zMw9xdFItq9WmtqXrDFio8AJsFESFE0LFd5ZL4NWZbCqs5L
ipwczkzu1UCBa+m4zDJbBdbMFBzusqNN/h8c3Pkkks/l46Aff2vl2gXGYtk8
0e9rhvq6sUIcOVOar1ZM0UgC8ByORX0vVzb5gr9+Q9FHAhvwbNzYeEg9TCPM
mEMt4mgHu/GYeCC+QnkhC+JCSLdmvSiU2quhmgQSxEPKKa9hMjycSOdqhTRK
UX3IRpOWg1SKACLp+pT1/46zrnk3SbMoLBcosdCEsjb+5wxc0T01aNcJfzYh
iF1y33TlRl25/EqKTnitNzBxO2cpKm2QXl/VNmvuQ4eVjEYm9PuLQNJ0P0Qe
RfhFvLbISqqmjma1G2t2Wo45g8r6cArIGEoe82SapbFMvUAGGj5qgVGTUU6R
Fu4cTAdQfr4w+KvPX+NXOmK+Y4JGKCfy1fr5M1ee/CoUOx3To5azmpoEpuux
T0lBlQ/eSkBy2Ggww/m8GZwi2jiGo2v/rLjWbW0Wcp1Hn0I3gG+3g2ZNqF2n
GVBEcod9OvPhDnOOTTkMxspML2EvLFbTRfmfgHLnbcr5l4zm8Ror90XPWQsf
J6OjBVZuV6DMxN8Uh+b8NEzuIdMR7Fr5MGLrC24SV5Ay2Rklep4O+uZ8HZG2
kHuXNQlJK4GGNgMhQRfr8r3EWB0J0+McwLxokWztBgWNpf+pHVr8lnwDtUQU
wmZfkzmza3vk8jVXn0vjCWuqPMj7HV+OSTgwl/BMDMKrJC9+oCod0V94SF2y
DbC/tm3HtZfOlfcBlWpEbnXfsOg0VI+9LY+E01h6EP8h609StG/5xws06YkU
6CAirK9MLNXC+NzztMZnPs6FjZffyrYQtXugxGmrCtFNxb47wFVk/t81784t
xQ2s981vb9QraXU/16VvuoIVNpe/F8zWp/O4JJ38WDdngN3qIrWggix05boD
uDL7YOMCGRs1qC4Ay7fQ/MIE8LvIJmWHASidQNUJpu5erBZ7HXVaEwqo7XkU
sUgC5ZCfuWYpCxr6VM0/3jZYZeb4GUqf5tu5Dp0w/LLWX6513uNE6Io8aOMN
1ZWZL7wtJtcu3tll4pBw0zfVwtXm8XKBv1Zl7UaIQweXls6lBPF/uqWjxMle
kAjAnxw+nsrypq3AobwnANCEfjO3P1TUkwxXk/aevDwYaoSaP7eCeHdAA7da
tnUF0Xk7eLUg0xxcgVCxNA788fgQnLbbSucPagt8ypY+MpW5tHViHsKGJIYs
/1jDByXdpHQ9nQ2LrsE7q88OXwhWOpJJlA73Dx8quEmNRVnqR642QbbTR185
1lLfSweku0xdX0KB+aVwDDAKSji1SjJ7O9U+jJKq9MvT1NBrM7I5CFFcPsiI
AYYTMJJaWunxBc7HbS75e86sBWnV5H2N9kvl2mtYpZf7ku2Xjgpii0e5ST5F
xXcs2qsKyqKzTGWuThnPS0Y9HUWcf6ow2+McYbC15LTBvDv/xiGXDnoUAyAr
CbTwvr8QkqrJUi9xR+Ak4RRCQbyYc8iN293311wOiCPJvsAOglcL8KpBjJM4
UKOO7kVqP2dXQacpd/gnX/TjCkFRAcPBVTT3SB+Sjg8bpJSP/hBJ+nxUSqKb
NQNB1hrfeVbTJADwydhMAyiJJEUa0/ATEPofTR23Av7cW7weQsbqT4TsO4T0
VkkOjUhTgNc1mjiep1To/qwHiGr2n010hPWtvdBccm/oCEByg78XLWJVYQD8
yAMsiF7nBHi8G1xssE6K9dlOYS43H5KhlqR3iDseD2U4MABL4TAhittiymgy
ydtPVsKRAy22eIC9lHPRNMs4qwcboTCzxeBFKEuiknClefu7h5rhMRuxkdBX
4jcMg3NzHUY/iNHoG7pI4mMEwasi2zGyI23z0fd/NiRqIgzVFzzDQX+xuWc9
Gis4mtD32Sw0+RYDmDytUXJo0Ll96zCpHbWlK/PFi7Bb62uHs+hxjdS4ACoK
kdmfJ0QBCDOnrGLRS107LJpUs6cHpq+fPhLiHcK29ZwdDrOGLU18dPJdhHM2
crAIMcE1j1HV2I09tpuvQNhhSIAIwrUsEdcsJEMjEgGkJ12nErKskpQml1oM
G3tqWpl9vu4Kb/UfiN3ob+sN5lshdEsOrg4TBrgUMf7jsL7AZOVqlo+AkM1C
Oie5ZXydf4uXrGIMWvTt/QQ5kqrvrnBAnSLGfJ6BF5EhHtwoJd0AgNl4Lyut
0SA8SsluwAD05rGy1GMFV9fOMD0z0rcowZ1yQOFBtED1jYDARQZtrg4ZAgvc
KRjO4Dnq9SWR5h705yEU5yjjQpQLtX3TRtbmUxg94QENyPJJrYtTHP3v1PIw
O3/YuTaer4qI2Hg797efcHv7ickkqBRvvbv/JtAlynMsWcuumPB4zgCU3XWl
BDh8Ns8dwAP1Ml3TV7Id4D+N5nJXRYS+BCR50KhNsH9HOjf2WreifT32dkvi
3Af+SP3hiZLqssyuJj+GcroMOedsb+eR3u8L7tLHe7nY/hng/I9PrsuNr6sy
P3WngnKI/aVK7mHwb+0usbkOJYlyvkYy04IB6xjhBpzsnr4zYRY27RtdK9mO
7RW51yDh8fDwMV+BeWyHH8msQcV0Bik1r9UDfXBXIlr9RmVhUn1u+920g0tz
5d/Zfcj+KalcM1PUrLMuTbJzMsdRc2nLx58sbYDu3md4AaSBGCbnZdsw+Ukk
sA3JbgfGiRb4PFOrsmoRCp51TXrlmS7PElsQ0EsG7i5LreTL3vA+sgqkJi7k
sQ1DyzpctFKoaZjgtzI9SgEItylCizNxDtxCb33SOrPskg7Ov1uuQFXqth0G
jL5RzyMA+n/cugxbudf1P00dhk4ZugVYEpmfASJodNzNWd6GIHcd7efcR7Oo
ho0wq7j+vu7Q5tfqEoIHiQuV0G/9JS/cAVKfUXbJckK5sTT6hDBiRUSLhZBB
X4zZfB8MNtft6XEWxjTLdwVmgt7FpTWvx2UT9hoK9+akmc+1hYPLc8osUlJi
IaKj567WFo2RmbXASw4UYjPkkkXg0ipZ0NMks33Cda6WX15vD+DPBKFjtwsp
ddvC8IqBg7GoYo2GdBxdDt75LcnppSCOumaohg4qf5xQAQXhWpfL17FHewvL
EtMKldNUTSIjqrzi/p04cx2DVVTJR4G34kPAb9Z5sv3HXPX1WonjbGneq8Lk
QOkTade2mB69U8WPLSFD2EpXFhJL35U8AcmcX3Qt6VrnXZrWuq6ikubk4Sdf
Xk8NQRaDHVuV3BFnkXYgakZIgCHdWVlZApxRXg7eVE1Zlw4/tXxNigPMJRvy
V1VwGVbj/TAAxHsrk5Ky24K+tU1CqOOq07xRAftJey2By6BQPv+Xb5Jbgi8l
GniZALbOreqKC78u1fW9M0CIVYoCxOC99gUneb/n44atGLendcGJ0RrgOkl8
8RooxTOxtACs460EXqJWc/SJUW9SSYQ3ijxlFXjfflunjQRoKYKUQ0A62Czw
3E4LR4soQKpLwFMrEb3HmRCxKec4PIwkaMpYGAz96NcxLZozuU0toP62JxmV
Kze4zAzQR70rvKd5VXG91guhfnKm4rZdCwYv6FLLJWuEElKUTIRnbI/Klmqh
htaDnjD2vWKFPUlQir13rRu0r6QxJdWOEvcrb4LmBlNGb5orRVHXlcob+7Xw
X0ye76u0AHSd17GxGR0Kg7PO5LX8iDP1lcA4eixXzGPUw7WBZHl0vz+9Tvec
QRl2YJISk+OuuiOB6TrCkAKpTGl1SSuka19iJkj6pUZr3qp3gandPileaY8h
1I60r+dfQALGWLrVhLVlgl0ieRgf+GzPlGCdGmf+tJWUcQ0wZ7bhQFyeINkd
KG//IHpjwG5sMFQFYmKRMeLAVTYFGMp1flC6i3gi7Q0I9oNdrBZIAYJblRrk
HBRJuOD8OOsPGOyKuocSFb7onSRTENQMWK+QMsHBMvexGboJx7WNCKCksfjA
5WREoUTAhbnvIL0lvfK/z9GY+/vAPUr6GbIH8rtbeR1g5A5A+xiFb/3v4teT
JNl3WB4QyMeUVXWImG8xRCeiet+s5w/NiH9otBHsh8P1PupHWjDJKVNgDun2
XojIEv7e5pRcJhCNud8ubIFS2nyPuwCa5OC/FBy7sCuxJFcMzByiRyAp91Db
rlVmfQL/aw7/VrVCG0PZj0PtbkKa1Fo+YwwIk9LqfdOORbeXeuHqHeBN57TF
ysPECWLNnjRvxUGrdf6HKXI+P1SOUSx1heyR3NyjsUaZdv0ReDbVjDDx/43y
RiVXkstNY0vVYj6VNy0X3iJ17Ptb7v8Nvt/77phKFAaHYfJ3ykczx1S0jgb1
YY3h0fJqwznkJm83QK3gue4ahIhAQVW2KN1tyBQkRWPvz3+14WhMQ14vrM3w
KHCQfovbGoctKdIgAQJ+MugEa8hb0dbwn0N67hgpsi/f7CK+qiG5iIhNNzto
jR+Zz9NkZURrpfkzSwOWv9dgJLdXbHb/EN+hx1YG7EyCpUOE3z0c+PwL2PSo
3DTwdW51GgDUgfV2GK764tOFBHXUUt+9WSDKv4/xaL1JfFTo01LkbfybTnTi
p0o1Xqa1PPHkVgO3WSqyR86GBXYPl3EalvA8IuGObTisRSsNJFqmMie1Uv3o
TIZFS9oxxoNNoZqFDO8E1xyGz01ZfBkEH2llHnzxr9kJi74Cq9b/kpPUZFFQ
IILlgOcEb2mIxkGbKu5SNE8yOXWn7j03DqizaJjYEK+wilpiDlko+jhGMg6l
Sa3tfOLfsS2YfA4rusOyF+LcO4BvbuQgsLz3PDRQ0bFna541l91jj/1f9Wrp
9M3KNSPkdHNH/x0a3CiYChduibHIsD9v4skBiBygAB5qI6A8mKPCaw4ZHdz5
oOcwlbnHJZ+RZJ3Ltdko5C7SJVLV+FYkaoKc3RE7/xlj7pczWI3tPa0e6wOy
npguHc+mI13/Y6HGB3/mw2wXObZFbcD0/a63pGbz8AUhicXhiomAZt7OYOPJ
QrSZ9URlyeeXcFySVhJwX5Qzvn5mX+/iDLaQCzv/bocc6965z49etSZKz01o
PgGTxHFTURsr/jPxmFA9bT51RzcL66MppxA45HzR4rFy8OeQdpM7l2jjDYEW
q/VsBMdrbq6znyWXSmpJ7kNdsD0jaZTx/xhZ8WKss2vc1//kcf9qUM1H0is4
4naI5P4xcxqAxFgpag1J2xruuVgSbTqEV5z6cOFXquDUqtMZN1Os5WTFTbSK
dBn1My1ro2bjkcSPpqfolkuopiuJBeepm6oGr8tMVEm6NWach8NG+oXIf4G1
UEVqVX2UtBgqSu1bFM2Mt+zZ6T9TPLCeaaxoOjF3yN8Knh07tEBr+qeJBOVR
FlqgiblTrzw4xiBe5fLGBwXs36K4fjqrWC3Bj0WwJidGXg0/tpYK+tm9iHoe
sCfrZPe9Nozpkt+ybIFDiU51I1NRDS1Zok5JHPgzgFzwm5XkOtuKvx/WhcTY
T6Hrp1dpRpY22HRQyVpVtq8pfUzWcK1gzUMrfPeyL8/LBDP3c8A8Q6PQ27F8
LR8W/j2FCCKMhxz2wgxj3M6xgyHxW4B3SjG6iLKbX5W8YDPBib7plRAi5+bO
mG4ZJFmSy8X8z0tNut6h6Zmsl0yJgLzkjdWyK7qhXava/sqWQiH7R6fzt1jS
Q6aEReAUEIUxeRuF6BQd66zp2H2732tBNO9WIZFNHdHbiZ2TzoHyb8JAhYhC
CG6BJTnvHbhJGUMgmnwt51VoIuD42kK+Y0NQFdbcXgVym/KuhgELFC0lwz/y
iJ8mDfCyl3wcINQ4SY7fYiGf3CScOon+PxiE2Vdmo7nx/aDvFb+JV+SA4eyh
m2cnY5dBZIjeDxEAGEr+xRIGewHB3O9kZAxnTDbuDVipvX2ceez+2EfEoepD
hh2AEqGq1Vs700b7A6D/qKmGy9cA/aykMhpUZA0LJ/L9z4fDCtbrYnaBQVO5
o9jiq0yX9Fe1vzppIZc/tUHEEY8CN2Z932SxaGT/r5K58hv+Zxa41WA8ZpNt
qokg9Cat+I3BOjFmPc+RvVjx62+NAJ8GaZgYz3pMchpMQeYKc3i9IkxaCg5k
jf6LDxRFlZFTseproIfqUqhw3roaht/14Tz6YBU18QFExh1rSXuUv4WEvmCc
mjH18NZXlNfM+00KIAsnYXzNmlDo/9BYqq9/OJUjVS8OF33xK4s7vR4Goje8
LZPzypsPeZF31Jik0xeAdMpqUmdSSUkCwYT0Bq4dZblXWJ6RvTTUkS/3M9/r
OmDKLpxmnloL3Qs2BllgBnyn3pDcPrbG+NhEtRuE/YTQT8Lh17rT6ufUVVry
IhWjxkMvoPmnRjblVMSbImPpLNYl9IVTmxO1Y26h7Ugk0oobwtZP2DHk78jI
BW1YQaI6WiJ+qhaccnLv2nYxa4ru98zVdgBiaOZ0X6nCe1GkN0opZDa6mQjv
IVJavSOCef2DAMsHP7YR996WpGAz7q/XRwp4Ebl5sfvqGtXHTcghXFoHw7jO
uQTODNDSU7/SB7QUYAUAfQYeMw97xp7r+RwfjSx3APjBZvSP5OcQraUv9CVm
3N4pxgrsdVTtr6ZK8sK60/M5IYZG1otmCl5BQ5KCETHP4UJBnx4gPJWVrcHv
i7YkQs7/JGX2LDB+fhDt7gnpHPnRFm8Qqv3pfzoQKVdBQe2T9sRW0uZtLoKJ
Z0QaKKEw7L7HOf8HIn5rqhQuZqX08NOsdIuGEc15/X7OQAwJct0tCwGUEqQH
Uy/2gBVc5v0C3XgC7hrCzw9TVK/EzA0TQXmhhDeluMRH/hCue5QUYncCfdQT
UJ55QOsCU4rV694pZhQvFD2wVNj4Kapj8YFfIXy18/pPS1aHgT9arPCU0GBg
qmGQKht/xj5FCNJPolbnHyIv+mPf9Dwh7xAUDnb4JbF1bLZ3FYLvyvbR+ogt
FRw9EAyDAoBP8jIcXaIbKDdB0FpWqcOvn2GJWqUxckDp1/6Lihf64vCNuD0S
H4HvMJnPiF7st+0rU0KNBWAxH9oP97DrwL1oGFIhSTSOv9KwkRzBYwHvu2id
Ztkc74F1Qqa6O9ST5SvnbHZoE/km5lfPkeQRbAKhXWti6fTRhVLK9WUjbnOL
CzGKqsGG/labuOR2Q+igliUd0Pi8OULTeT88l7TkXT8svhYsS1PgqdTtsjE+
H836cUp8rU6lyMtMqOHh+NS4nq2pXrqFMxMZ6j5F4y5EHF3CxQC8S7pd0wXO
d48SGT7sOkl5rhK82pKnVTEnyqZaRMRSVjP+pP1wsGX9ww9ZnCDz7j2/A1rI
ouRvhwTWeZgPRCQAmnaKyDfDn78Jghr04sw3mUcIxXtbLQ4oKcDmprzcpFeo
C4T8fqIkaxHF1lQGqDFA79JaY2BPami1pKsckN3qOL00OeljpY3Osd8OAwLo
QOMKnnnpYdBHaCceO40CF4Q0vP7167GSPsqWfSNIOfMXoJHuxrZPnJS4fiH6
VNYKJZmIgB5bOtCTP6bMbmxgm4u+HYE/3/aJObs/vgxhd0NWtaTSKYRkarSs
1QbHM5J5tANaS+QZTl53XGQBXHR7WZZ9cfcML8bsRfBXT4/BxFSrPDLYHqtY
PmWDiuVN0CN6JXYzZvcFpPHL0Ss8NaTE54sto36e6NaWW1NVasgRpgWuTqCD
g+0YqzpPIQqwQ7NtRDgm7VYGlQLbsZA+b+YCVslFMFKV4nWUMNak98UDEXyL
0yc8Dk5XylQBkG2tSzVg23VN7PCtos4Hb74NLnfQeC1FeqIajDlpa5jm71kf
ozj1BG8BPgobgvF/YPSv4sMagE9Qbzh5i+UoDWVsNu6NncZ8vWeSFR6V6Tkm
Pb4p2fmVNjC9Se6btHJ0yGuNVVMwP6O8B9TRxHs7IRHLSN9mCISXveKQ7Zdo
RBlU65RH7k0802G0F9S+nrQLNp0n/fHL74Fo/89tlFSwY8r3KNrt8/R+4AIT
i/qkOizlrRDIsFPXzhEkMIZDjQD1KWZSwTCu3DWv8gNj/tfZCf4anVoGUWx1
WkRWNIoYudtbpVsjYj2NGplq4nJRDHOGzfTtdFj35WigHbLY51G4eHslEFvo
ONCtqOAuY/GztvY1IK+KL5cayQ07SbASyXd1AmkDWhqlDZeXNpQkn3D3zFY1
0h+iGW0iUwmW5xkq5RgizmDCRT3WDyTkw3ZJuRehZ3Oc95QNotgKxbd1ay6u
JAXsGsxl3M7puyxyZwNsfgYOuuMAPBbwgNlUipsMKPMzlQAM2i/ijmpQLOek
y8TiiDjqgmJtAgIWvB5M6nhZV+wiu9V2v1+7zs2GYkY+08YJWaMezqBGMjsd
XZC4xfXPn3+CUM3W9DcSnsLJD2jZ6XDpvqX/KTcBWUhLh4hc/72wXcMvVRo7
kne4FyVOwKefIOqq9zJH5nIsWZqhcRvpESglFxaqdiXbH8OyGMl7hJJ48GXP
97P1wn/vgxgr5GipdldnWzKbXR9CGaMDkknqrDgCwTVUMNAJ9qKSQ6YpDcB7
9FNn9RZ0xirn4kpk5HGqN2oahjVYfAAYzPi+zkKgcFR+xj8EdRUULlRVpCYD
pvdeciEubgAw5qR/NT3/wS4bxmlxRjEYxSXdG3Hzjce1CMGwsuS42mQSuMbY
ZnH4U9xXb2pt93Id7/qB0B2hZhADAlfgo2MEvVh0Tfrphl2SFd0HljNP+EDb
VYuMHeUsk0PnRq2sOJecf1NcvVrb4RZ4N0EFTLdxCvzCQiMXYnQsX2Yydo3U
yt8EFCp8JMGiVqeWFUjFwk0tm+PdPAhRzCjgCQ4cm7PpAca58WtxYJ0KV/WX
PimKVgB5FuNvObHIq/dbjE6DmnBXezwSdjHHqs3flgRb+P51ujaGWB2cysvX
Un/7177DRG4Q/sLBYFW9y1xhYGnkFDjX6ivKtJ8wLWB/6DObtAVOTvH3yYdp
UFf72AOs8MyjUqMxWWfsMLsBUfefFJHA5DywJhtoZ2Tv8MK4zlVJG44NciLZ
dBq2lJar8C+wApxGBRWkSN8mWw6AT3qYTpqBBQCvbTxoKfKbE1NvGVNSnrUT
rOnBSHdEhCFlHaUzNq3vIF6YShMNOMEQSbtVI6NaSoaS1bGodjcq8otNrvXa
eAhZcepUATf8JnWiCmB91+QBb4ATqYaBu1cixptXB/NGXfVdJzcV11e7dguT
EDHLdIsyDHmdVw0c80wm7OCSJBDTcoHPOn1KehuYnXs5Xxd9/SWFQLhc/gd4
NPldtV/tW4xxAwNUuPKGk5O3jav04PKoCpy7hlERyNiSYPONG6ESsS8/sW+8
iVsQqwutMNqMEZ9A9TSerMHs5XyAvDdEjcolSYKBJxM5Od2/3lmGm+5PCxX3
0Iapv2Y+sQaYWOS6IBEc9/smAVi5Wun2WqXf13T1ZvmMhUyRiAvtwBYbCxDE
yfZkSpC7lqEQUXMlIoWv7pQnlhAYVnrVolWnosaVBaU7E03CXiy3XpbJXCuI
uTWrdngYGPJm+EAW4XhZrguwTZJ97bWU0otQW8y5U51GAuYYytCaChAuK1wj
Afkg76ZV04/XKGocgE/yfaTnIlhrnYCxbQC6qvskS1DGA4udhHhM2Ia4fGje
zJCtoXK7zpQYwqTwD73/1k5sAmkx9VxKz73Y2xzjsbId07TfeWcr2ytvSyj8
v9K8i3iGPf+FaY/QUV8JGiNvpbX2kgDF6FXyBKgW9kWfhfvCiS/OdL7D1nlB
U1Nsp6Wd6uNJ1n/OohotYAja/tMzkKdGW+0oV+s/ryzOup+m/+/99G71At1I
P7TMFT85QQi/9bZhV28WtL8RwDDPTQy08SYWe9kyGTaEWQIm5+tTKk1A0S6r
pDXv+qaRYTVVlyTMq2cHk5mXFkexevKr4W1wN7EvR06HGjPHG7zmlwK3Zolt
sg8g0IPz+VfwAD9+08tUo2b+th7Z/OBlUI46AjaiWfEqifs9an0NGlt6ksPa
O1ugR9dSU086UX5WDIptXzc1Fm2zwUnqUOZQWG/9xom8AlP2cdlkjsKHgYwt
rVJGUKZKX3HFX54XcNkaPmo2gQ+XIjCPY7OV5avNaHsZSvUidvhuP5umby8E
186ZSYa0jvptfg3oFkDvSt6rH4ZC7POZ2MhRSKUIOOu7RSZiTgZe+ezmftlM
kMRPpKEPyvrPDC52NkZFQcwBRsjuDEmZA7j66+NHHYDnbAExSlZIWoOQNBJZ
II6RWQiO5KiLn/RSv8tIdjqDdzCaDd8IYvT56d5mQCqeFOmbJQmJKYRhaID/
xh+ziKpZABLBJ8ZxjtYNG1Y+PU09wBZcM3qx4TZxuPaY6yWCGOgu9UuazRjr
nUyaW6OfwPQweeCNv/noA8Bqt9TY/gpNEYhhWapIU5W1v3KD8KUqpqhDc+4U
KocrXgeimDFQLGirjGCoGoZQlUt04A35aemxFDq34imLl6gAyW3l1oocPr0s
uKCunqmVZRBNS8qe5LRest5GM/npmIcprQIxHE7P8GZVpnqPG7pnNWp1yS4x
7pT3vn2TO/g+pX7oJvFWpaOBZHmg8VJ0xqNH3q5TTHSIlI8z1h3Ek8KBERJH
sFmjInIOJUItVEe5pES68fmYnM1Fr+OJ1C4QPs3iF5GO/BPuCTkJleKu+vyI
AFqtOV7TCmB8rBwxtGU4bk6V0uprzb3IvwKDVg5FUcbjW/Y+na9h4e6S7czD
zQVYAtBocNKo/Qm4lpKyVPfh1nJbUVvULE1X7Z/1uNc1rFR2p1BQHON0JvYM
Y+xFN7BwRAZinFYvUN5zCyfs7m2asvAPs3wgnZrlRjktXQ5Jt5i9uEiRCJC/
1DPDNsTLbDXx6gsOz1sAeJWKdktBNEJA+iceru+UaFLKwqtT/IHJOj0tzDpf
dj0VqH3LF+yz4k2WEEDDIX1CqUqwSp7cc2XmcqPJely+ESYPvxNEa6AWRSRC
jBSsKDUk49ycmvkKHeSdTDdnzARd+/j1FjQDkV7PfN0afZEuOLANL2Eif6za
gyZIUl4ar2KpxrI128vZWwoy7UnIO8QDIG7XVx3GkL9Guo2JjpzMz1IAF6b8
BBiBVwGfRyY0YobTEMoD5/oGiENdC+0U+hT0u+YexSv7TxngsuoknhDp13jw
K6H8xkFraXqyeqJiRX1H+SPKBf3aTVjKq8uak9afwReJLIfZE6GPC9OJUSKn
j+kNjMVt19zfccPN2O1KVTFuSdWK9oHcH3rqoOeYRwB30OuHps91bJwS7e+X
0c6tB+1kflGlL8b7+SBOg6XJbyK6rIRE9Ogp5nu1B2Ft6snV9fyETgBDGBSJ
iObWo1iLcuBD04e/3pLw0M+ZahOyqIhKc88wkScVZ/to0PkT5CUnX/8pSd4y
GOEVDj5sANeVVgHgZ3TWK4UWzMq5FqSA9TmH0hERA9Ia1/KzIFmi2fRtTALA
5PogON710+EmHqS1AcbVM5uGhu2uw+SMgVQySDoSt+fAPe7PqP1Cnjt1K2o/
diCuQPdVqI6faXl8yJ+B25Un5jMP5uag0I+3l5XpuGGobJvG7iUMzZPrUoH8
vGo2rLGuJ5c3qdKLdF7gZhFQ0MVowc/3Enyl4NQ5F7IXCv27NH7YAJghdKW2
4AOJk6hpkUswNh8X15ghzCN7CrnQCJC6JXWTt/UAP+ELnnE2+w6HZQNNLZL2
HqYFFMX2u6WZYlROTO0N1nszptDdyjFVFnM2kybeTdMAvRQ6HK5wEV8pVe+o
4NUAcmSWQbeGpzONBP1zOr/T2WZXduiidv9qRPH5d0UdDln9a+laW/Yo70Hb
pZ3u0JmOZ/PbR707XzdF5o1X17MoDOk0bO2eW5AhujnXBrNb6QDBS0XwuPGh
0gs3DWF4u+dEWfAUvjurbYE9ACnQj8Q3oA76USKasH/tpLNTGVI6tEKfJLB8
fAxPQz2H2AtsTL5EvlniNtYGuogc8u74UPxzP8SL5WpT6OkkI+W3ZkbtSoCY
pej+ALDJv9TkDOxNvONSbym4wyMw+WyJng7gejdcclaNhcwjNrzcc3wOxvXY
5PchnJ9Iu32OOwGFbgACAiCrRhogKxAdHpwY1h+DaMKnh62M0wtx52uOgr4r
Spo4x01qRu3ehXKon/rFa+LzK4BOyj5h5X9WW3z7QnT87KhxUhMacvJEceGj
7pvzeqXKeJy/yw6Im89SgQGk1bmoXy9Cp6iqBQtw0AkHOF2/1eUEwavSV4IX
71mixFbJwP2YBjdCNmuRa0+MgE9XY+kGv7MXAZ4HkyhJG7o3FNQaju2aYhSa
l9WMYBnLXSEturrLd3o3Io8IPzZF0JpsE9qF1f9c2YcTile+MNUPg+rArIbH
DfQ30BPnTJiq5LbyaKJUkLABFB1fKgurTT0KhVZ75w3yWlW82yAXuszazCzd
n38oiUyNYuwDt8OUmus2RjnqfgpDTf+6R0fxDHXT+8bzK+8YBYG+MFA4YEfD
QzxlZGwXxErse2Ha+YPqmBuSL4E9wbZw9SSXkSUV2PROTFkO6p5YAgG5DtAG
nwwSSarC4eRjSGeWCNvy16j1zzMk4pz8qEABRFwjBTF8cUsHQ46nHx2JXiF8
1IRta+H70VpfGM/0QjlAxrRS4N6uZKf8m5cs5e1EqFM8t0adfwl6K5Y0uGbO
5fByafj+LB7TwrMldLWu5oUvf9OXvQWkOvUpvwT2CsUNV8cpHRv/zGfGzAsW
UWGqEJtvqeKL++3z93T6y0La5x5BXUefZnTZgB+yJVQWRWTxRpdZqPNk4Cb9
C/Lx5T1+0W9PJZI9PPr3KEIlpD0/8XtPbWE/oCVhNyfABJqXyO+u2uuAqKMC
Qi03OcDHkDY5wMt7k4Qyr1g3LRGLwUyyWtEvQOrByNus2JCO8iiFSJcPlGfb
P2ZsWm/le+yHyh8ogo6MGHVqylaa0IdXgzfBxkrKgJlnyJ27J+BA1wSZt+Pv
kBRWoF8zCdSzofpGehzGhkkvUpDvV8R+GvID1llM1irhptwNWvbHtpagDITm
wdhkkfmGpu2a9Vjjs9lYrHXxUQ5GOfiMtYn3VZNuQ37hTLKxL33DaQrL7irs
t1nJfIZ2BRGdHQqyxMLFbB3Dx5BYrffiTOl2y8D6Ckf34F555+erz1mDfkkZ
8PtLve86cMc6rmVY7Z36Ho4/3AdnhDfZLrhDaXTV81TwbQ2GZM3gGnQ8Yo7/
jKbf/P0L+b7HkPi6zDe65YpsOIWbk2IyBDpU8yHCFu+wlsW5NgjLJaYNlnQG
OJbbmdkKAdycen0Mzk3ehESj222U2APqBplr52q+akqM64Ru8kEYc8FReE6G
0pwWQgfgetDn1J2Vo3KOUvhOCI1T5CI/gZ63cUtFhE8is/daXgq1GPodYlhR
ySFqf/whOVwiYcl8dOaBL3yh/iRIoY/tcv7qh6e14wxPuAQU2P/ChRuLBdtI
PO2+OQLMb7NGfRWKzosniKF0N8e+zAkdJHieslFxpGkx8N8covi3TjPv+HG6
gHV9a9+DMh0t1GvgUSirLVFg9nC138qF6/X3wgAToeCaJcN90kyxN/N5cl8m
RNdgVqDH7metAthPHUHpTi9coXIWuv2014j+Ra8E+kIM2mfwFUcFBnwRsIhZ
eyJZFgGXRI8bZUZUTRZNfZeWYNKmohVO6DcTJvHDGE6ix/tXTLS0nQ7zQLa4
xTGgA0pnhT7szKylPFL9KvXHmmzwqrMQUoX+4dPL+R64+PzBRiYJGRbqoIqQ
Q0Ff/6AgqAvI/QrMXAorfJil85qaHLoUIaNb1tIlbBPPF0NgeunIG057rhr8
Yc66qsXyMF0sJixwQMg6hj9vvR/iVUyXE2oHv17vY6QEkfzn/bi4ahU4WDEb
rGa15OD6HRxewp290QW8ONd/XYPGbgsOIWW2LwGWpSHUJ9Kck7kM4RUMSfne
3nlf4OXjU5Ztg7B52iTNSrwXPxJYQnpqUgXHD/XvMm2+yCln8qIuE79QL4Jj
5INatPoXZV7+I9otk5BBzAU/zH0IRNf4d9KIehzCOz5vLQqhFLM1oQF/GYgP
kp25IKi9BMlu2iq5dh+e7XaZI9dbjtyvPJxKo5o0C+sJkO/RnRX9QrsH63ux
2YIv8EzNmwutkgf9TSFb1igETKg7zFBaTRh+Y+2h2zD6dlFzUj0Sd1D4v87h
95+iHFpJkRU3+fyak7mV54TW3+fHnWM53X2CoqXj/ts/A2i2wqfdfMRIXPXl
1d2UKRLhaygxf9bJp5/45s0d9i1T5Pm631bVTfLqHD01rBfAS6yDMubPYSqN
9jf80vx8jbRKq1wNCWR826IYh2EfmIJgydXXH75Z6jk2Sv6Z5sbHgW+E6eXh
gRFOWlzhInLq5fPJCZgk2CnL57+lLQatEzFldMuwvzB5FlKV24SsTReWrqqN
pcC6OenpbMAZmN/Cn57TTj7EmSCAqiKOzkkB56wXx7MvVwPtNbF4CWWmE+mu
1+on2iOfRDYU5YYjuvFTxX18838WTYKc+MuDsfnaojq2x/4ZbkCdP2Pi0nFQ
LkrU+RCfA6lQX3oECj09bisdoEbJrKkXHhUGzp4dYOxt/aS0XrhPB67vjPPX
QIjHizq/m4ajinLsm6xMoq4Jib3QvUQEFNSoiL1uMn07BgoABcfmA3Gym3OP
2vQTaGmZBBECsr9vneQBKf5eVAcH2WuToH0Trm4NwgWu83GvABMcmYppPU3P
8OI658Z5JPTtUNWQCvp7aGL+WonLgMruBlJGrO/7pCMHkczCUk+rEjABuCl8
ndY/1fP9XZ9q/AnV9uJG5mO1YxXjsOW+oXqyOjsgarNQM8TCRQJ764ZMGKcA
VPoOXcbr10g41H96pDGiVj4eJB1e0NIN4QPM+/E//HtNnt0P7kMSfsOOjOfl
ganNEnW/bOA3Uk8i08n32U9l50Py9qmtUMADiFyxGMm1DRBWQxinF/5d7n7a
SbWfNUlL4QDjvZZkzabMezyq3CzyhhVqFqCsK8JuV2ezGtII/a3FlfU0pesa
8xk6HpDSRv4A+hGA1c2NEHfs/tRFkHbOF4uwnDb4jSpB07cWSZsOwXx4jeFU
yIv7J2SgsGrY62N4Gm5rzacl0gkz3W4Yg6+ax1d4fXehXOMI8XGMJM5fsR52
KeJZJ9JF0A9xplhxUdG6s2UiP5VU/5DNsZ/4pndxXdgc8rhHT+0vwk13Ok0Z
a168OQbpvaMcClvqjZC0SsujxSFwzThi7plmBbOWq6uRtiPhXFgFznEJtDXW
Aj6M1x93uGqEZhFq/wft5OcEFQu64WSr/b0juRaUmEG2osjUmW5O3/TEQLvY
HyYnB0lDQx9GMB+c2ZQKvsGXDqN5EL3dseV8v5HlysJTFBEBjCduIu9ONMAe
+7KEdgG6LLcsZsl6wVCuMbhkWAsJjw9cwFzhBYGiirhblTXxVt0YT+G17220
GMhhBTW13j8DtJwaFE8HIFjZ087aIXMTJRppgFH1SRSDA9snBjWz9P2WmllN
mv57NlTmn2r1wzpfJ+1m5BJ6IrddebROkorPA4WbiyUNU3wHyGVJaCHC1+GF
Tf0dUHZkw3sjk83hmWmcN6SHTXdeNdLShbC3/+FesslC0GMmyXyBYogR6v1l
H6Zeprfj+OOQ/Elh7o/l/wRHEra1IUqMolugHVaR++ImcwF6fAla0WE93PIO
NTe/892RcwmC7pvDweBLfFgNto456LAxByG1kE//XOkA5zT8Ro/K6bBil77b
VHnary/uREPXmTAo6rP1RjMrfqzy05xQ0fiLOY090UJKv04x9ewVJu8n7I32
DUlfnTDMMlNxteDmWpuscbkYHJT79JT9pOwNFFq9a9Lkw+9MxZPYJU45qURF
e+8LTadulp3J3rkVHjgnVRXOnr1uGV2H/4382xb855V3R/2vsr8Q7ovQVcpU
TMb/lY8Q7Fs2quw5OjfpnZnFzaT/xvRpPip6wseGbXaM+gOyGbeVBWxppF9/
C3kk+d9Bo1MyAEZnFjymBwBxmdanDHOYe5mEU9N4VChcE8KNZQfscpX5ogaa
QcRevljEEdcbEDa7Z5KJedilOV2qJvEn9q0hcNltyny0+8X2dS7L8OFt86Yw
FPjf5zWDZrMwLNut3RWXblo4v8Z8lgzqrRc0IjqwPJtXbK58bspIIIW32mPt
LnSPH0GBjNAgI+zC6MVlfWWx52+pnmseQZSkF0YC2IyfA9GtrnI7/OVUmTkX
ZIOEWpe9yMu6+sPd+fdNP64T3p811yykhIhKV7p6pCPm+/Q40biTdaxZBd4N
IAvyZ8G8wFVAI1Bt97DC3HYXn4xnnoWP6tHJi97ZA8F2k1Xqi61frGGnG7xP
2tiPpJjc7rkPKoKZ862DTW+ySZRzKFpIkg6i6cuPHCq4UkoNunR/XwAse7pD
C/g4SphDpIQBGM+uV1LWLYDekhgqDjNql37NIRPnbQKvN27v8GTxMsZ4FcyT
+CrDwA6bNMQQIYr2N5w6ZO5faQKM/LB2EHhFor9x4So7+/ihzPDOzT9TlXie
BMTgj7EQApqimYTWsn8FEjnYwT/Ap57hfd2At403BPj4Jc0mNpuuzcp+TPE1
Tmy72menwtlEopTv8spryCXWIRKOVKI7pzsRQ7qOKRQJ8C8Cz5NyHUNaJIIh
3jHt9BdpT32KaAj4Pl6pRGcZa/Qv7TVBNzCDOONr/8St2dLvShiHHmTUBYjn
2xFDt+rvZepS1YEM/t0jzP6OBcXal5GplLxXw9RE7wSC3NqMjASLv5GO14b0
hDJSLEIA6pkuVvAgR6AXreucr7MSjd5TWniDlHHbH0yREfgD6jXuw5L4AV0I
Q8Kvq/R2bWZRHQpqkMgxHmaPyCfLCrUKrgjo41Geb9KLI8rQvtcd4G2LgqVR
cb/vbHEJhy4k/tQATkEt8FJiM5mI5QBK3DbOj/B0viZnP0Vj2me3qJ+83NFS
9gkz4Ja59a/SMaevUt16dHBiBU+WMrLq8QEC2UY0AQSl9sSekcHEiGhn9rUa
Ny8WB0l1YLRp1ZyUWxkIrfr2lKpZrvEOQ5Xc2k9+cv6WvpBgdY7sxtxDMFLA
CbsYFUXZenoQxiO00IOLx4XFXsm+Oq9CQ8PzP5Z8OseDm/GG/auPdkyeyV5F
m3HLKcvb96tNZMr1UUOuGZED8464AABk0o8u/klgTgNBYEiChV1EGAuQMkUe
UanJTLyV8g+OUxGYwx82O69P9aB8OYjci8rOLVj7vXM17OgY5umQ5wjiaqB8
QuLFipbnfHJX7YejTVkuoeXpt2eggu6+pxw38ifysidsms3nuBi4Ie9O9s7R
0uidqKfLiPMAwBY9MIC8Yaa4VelOgjcR/C+tnJlEQuxSKUmR3lc4nTQvFAfW
203tqfEUUNVjqHewWEGUkCzeXylStw3vjbYwyZUeLUPnTDvARAShMhT58rL+
o1TYF7qZrtNQayXoy8acP603Xrd+vEuv5gQh+h0rfVNQ5x/NJy1gjWto5oqx
SRWfgIVgF7BHNpSQSMyIfZGVi8nEpWYu2WI/fWuGol5NCJwxLOYlFqaZaKPD
QsLGv97LIW4fwjfBwf2Ror36rN1XFmOZx6tUKC8AjFtx5qhPDNAtezrouUVy
X4CRq3Kv3WlO/TteuwEwSBLpBgIiJyVFsgzd1cdr/K0LRvMrE/6HrTk8eaq5
KEjo258RV4JaXWdliEEdHKEKOPt/tF54yB+F5mLJtVoLqlLc1xoKMImStLgl
tuSMwo/oXbFLKYAcOHAbpp27trlp/9mLE+lCGrgQx0+PoKemYlMaX68IMEHD
fbgUMoEYjFGgSd7nENCh4PDl8a5YAsym9NojvV8tTU2Xk1rIWugFJ6gaG89T
VmsUvQhWLtH8x7cwaZjpmxZe2XZlqR4om+du6jcmN23Z0zvpwlV6ED/XLXUV
ARfusU/cAN7R5I6DZBBYyyFtrEerV5gO3AmpDHNusbo4WaJfZwmeWD79mfMt
Ee/eodi94IZQktnwsLAvRK4pcaH1SjbgloEv5Qiipo8/h6hhGWurBVdSLJCr
COTO3K/uL0vfqo63MvlZBFZoMLG9uSxvrLLgDZzW8UiPDLkKCv5/DQ1OwPaz
HFFtDiqkuUMFmOldMsTyAZOgcDz9pvWm1rQWwiPKGxxHveihqjxjQmTdCnVk
btTnKP6IUM1ZhqQ5Uaeo24Kgj4YgQbprwDpBtpbK2CNq4enIXtv6BZZCHivG
hTsowQUy4jWToIiJO48crvWd1LFBje16jOP9RkwTRMilJEEToLCMEJqQ4YNT
FGX9yxB119krKWTSk2MsTzyWSEe6Pawzd3+sJsSOsGGLA+9xncP31KFemcbC
yHmQYXmpfZPegNf7Q+EGXpp14C1V48HhDWebEtHPnK6RO5HheRXx+G/+iUJr
ikflDtiSQ1Dzn1h57yw0eb/5HzeqemRSjXNS0RVP8HfRUUPyVWuN8PAKMGyQ
qkyKX5mh/Jl+YyO9UVg+tHg6gBdqx4DCrvPuIBbT1EbPdREYfQMvCS1hdGIA
DtjDuDgzbtu43AEt0HmnvbaGhfAKUsJTj6YUw69dPf4GTlnVe2joeL4saHMK
W6nN28Nh0l9EPilE5EAJiNJk7FNXYgeFbWarq/r4+JqzJyukGId7NnTjABw0
FZHs1YgdMKDRCX+sLQ2QJbNToOmotGs3CLF2DIjNMoK6WY68uw/k9bHRWOZa
pHFNnDb/j7ausCwimQ1AJTOL06DiC8ucQy4SUsrKGl8AQij7AZN79lyyY2Tn
KwLt64JS2RC/CXgONnQYEyoZnj6wdruI84JcpW7gu3I/mxmJ29SODDkmK4bn
DUbP+9JsWPlrRy7uSE5ek3sXDTFbuSYcOIFEc+8ksH7gjMd7jlRM1wZ9cjb1
Vc7SKuvjaDUIRf6w6ZDQcsBlmbrrE87c6VoOh58x0ToiAU1Rp6YK0hc3pXYA
M1a7By9QOnHAzHWEJHLfoDB5dxES55bM5xd2SKd64QxKt7ozuMp0XaX1Bnga
sq6yi4x4GiyJlfOcxD3kKXgebW8ZcIScrwX+nPeiFNRaL4qfXTT/2w06oSYg
9bvWdIiWVTkFyF57T1JGeEwoUQuZ9j0Aj0S0Z453+wAwpSRzq2ufZe0PIKM8
YrxQzdQuJBEy+bSfs0oeg2vPLpVgSEiFwcsMt3tftiOoV79epvdOaYBiKFUF
yTTuwXclr5A0HYVWHdRuSqVrWVfHfZwKCWO/H/br+du3M0QswWAHD4PiBRfN
cApzzFrYY0hcQ1STmLYHucX2QoqJ6Rb+L0tPdA0NKzBFg/Gpdc8NTrjulng9
jjA3TV7T/FD0s+GPo+uGQJ8hmDI6Ss1wN7N4Xsdo/kpN90GMg32QNuqoPRrv
mLUwmaDR7G8pMDQ0pOZCFYZhJo03g3Fxo9dIt4kg+GKrcpH+ABVyytW+nt7X
JQB8Qwh/mSFJCyhFTbpN0d8bo2RB1+LUFWbNK09la3CzSbauvir6+npEoY6j
0AJfzBI///WZ96GM7UtlR04iyNgk89KrG6jc677BUUByjCiE9NVlLejK0DHm
vK1iiQqQ6G2b90+s7SOnlCnJmYCq/710hvchbypncU5jRlsngv3KMgCoEYZR
VKs9V7+nZBszGhv0M4cVmZOlUciB6irchWoEOUtW0WNoiHt3Wy9bvWLTyOiA
vlPEZ+3IatSPKfvex0Wby3H6Z+kQOro69g0E1mGluSm65k+61spxCaPwmaWg
9G9+c8xZYp47e0U8GTAGNCDpz7nwBc+BtwSnPWaGlwnTSgSAigL1GO+wSr6E
+WMaSrGNwQKCF0XjeD1uM+iVv6LjakUFb00CjxCmSXYizQiT8Km+yl12sx4t
CIk3g5CupP1uF1lVVJnrGry9p2ACEXRZWa5miaPtVba70lVtUuw8Qw4PSta7
kmUe9GQ+nkbxPeiLtB/nnX2+n0VrrP/DEN4URtAUZ5z3KzO5GSX4Z/Qds9ks
qxgYJnh7wwfFQvpee/I8iGdY63lk7KW4AUqhoRwu4biL1/dw7s/Mz5Ehp5PG
pGYfzvyF8PmgjAHbzQCQl6HuGZB1vetZTUXDPLJE8jcC3l8rEXJAKA/t5A2E
bus8C2MR/aDPmtDBTM3K1lm6eAYPxbo3Ws6lQe0KQVX8d7ALU2x1IMjQE5Hd
adm7AcF9s69jWy03t9mRx9XEHu0u62nht5RiOYebAJc0Wv6lByV6TTRnUFMn
ZYA6w2Rk3C3lI9rZmKROB1qlfuJ9FDjtWoAzKTeDyIYmiCwDEH2hAjqqzY/C
E2+BE5clY/qn/qm4Na7MUYJ4Negtuhor82dsZhVKtvuz688p78/y3nQh+1Ui
LRdw1HcIX/WQFR89nUeiDq9TW3Q7HmarrcQ/ZaWJecnzGgJrZWmoLp0CX4O8
1AIGWmBvYmCnAsmaSn4u/25xLZr2kzo7ABWXekrnjH2Dyrgv2zcJYa7xpjHH
K60UbmBHUSUCoIizbh/3nTk/gB/1LKZXo5pseybDY3TKdrmWx8zpmabwc8i4
5Xvjsqlo3YVlzsMrX6WXyjVQCIF7sk7msgEY6VdodcafsLvYBrSK0e+TY1be
SVQExFCg/5f0JSdPptdcq2aTF9r5uL3nDfgONmg61ehoZ+JoJJOVXxIQBacF
olUObyj3oCEhsyMEu1HOwEsmQW5Pj7EIJXUu7H3gZzNBZglAcIjLbFCAHoDD
xOQMQ7SxTXaC2ajO4rPkfLolmiUqhnahaWge0p4xeBftI/z5pgAfvvdI62zz
m1/Cmulx8vO0XimxwwJC6qgoefbhwt3NwxUYjbcKVLMmMYjWYjMpCjF+Y7AO
BocSrCI62jT5k2GvZPr2NbRB1Fd2E2IkfnF7LDcg7qrxr79LwkNBODRzJmYB
h1on/beWZ/TK0HpcLRnVjZUgxz24G+/gYlkjBce3ytVlbWyWBrZin9jA0Fr+
Gsl//LB53ZM0I/be1Znb2GMFqKqe2AfKfUcbvpfif22olVJewAvkdbKAxp4s
NfPVKwXf83BOaYhMr9OXCApy0YxHEJOIi7IMu0Pj9M1Md6ixAI6VN0Yy/BJv
2EAbTHxTql8GRGwd1nzy6ehBcCFHbkDwPAN5P2niTK9zToZmwl8dRBnbjyEH
OTck/0sTfePZLOO2C1Tlm2WvhfbCjtyrXYqkRBCNC7C58mxHpcHT9xtYTq3t
Zl2oDvsekyfDaFDjqYrgwlKS+9WirAeRLZ50bx5v7IbWtVrzTZLyxgnuq9ux
wQ654B6I8I9Sb18c+TfIQQveyGlzx+5X82kX356dJSgn9+9aveYxopXXqaFQ
zQ3HIpDUH7l5F872JAQJNvjiEnNiKK+kkbMq0XUL+VWc5iGvD7pubeXNaoHb
A56Xk6TdN2tau/Oy8t2c+pVf2zAXw3dmlyT7GFr3XeJb0aWBV6awvotqY4ox
xHCDfWmnGAHyh6QPuPcD1HKRYOMI+TBr7KdCXdGL06BZ1N8Ve4cY23xDCc9W
JLJEx2MN+VAZ+FCcTldC4CMr/H3CA098PKvryP2ivCfeM4UHUI7oDTWvPgOg
QQWk3+WJJzZCn6c6OZlXMNRSjJxHs6PFO1lNaNDiPN7t/0dwrRswj1nz/sF5
fZ1klsl2kw0f34XO/+XcCqjdktz67qop4g+iJVaqEsLMCPIETKNVqjPp1HHW
us2W1MNLhG6GpowDrNFlT1ZFS6q9QcOpZr6zzSUPpvQkcZzRXtAVF/mdI+Lm
Es8vpdJuvshfOUwc7A+b4hU084Qy9XBS6bAqtLIgA/KCoUrsquO5gWRfZsRK
B9vib5q+qykkxmJkcclLBfWwuDdREXdk/ittywgeY+1Q9qC4QEi7xiEwPK7w
k61zWwr4Q4X5ogULnzLMnjkel6lm6eTX4gcm62DI1WpmqZmKYCU71PvYvf0b
9eE9NZ1HiyecacT0hbpLxTMntFCIIejOpOex3S8iT6sMeq8944CaT7L1ZqwH
ezH/6keUq1vEfMNO4EeesTuHwWkiQXkxor8H/OTnQrAD93q0bRB+SEyFU0DO
nCEFxyun8NrcElmqDP+/i1lZbl8oKRpizdqcGC5I7MFworXOqmQwunyg/xlL
i75dEb9RbyOnsy5enOI7uWIP9KE/HtcICRqVt3Ie3R6q9tSqI4Ef8ZBAglgX
1k3QYHFy68FzySayWDK5ebmdgD6mGg4VHeSEZgXZK+sJPOLVZ6Gz9P5DX6/m
iz17FXy26O9NcxkO1rF2eeFKieWnq+/or1LFzHNn9ErN/laToPK2R8SBueee
2GS591MypAJ9hwcBe7oe7fVSoGtrkfOmyfELVEQxe7tzj5WwiVgtGWpoF9Dq
nM7hpXR6d3lVMV0QkUGufuHOEh2bFEh8ps1EdxCYLmRx+iG7iFs7s3y0cLKz
sVyMvHmiFlr5wU7M7QA612WDB3yr1cXXEc6ob1TC94Yh6NeeJJ7QUlRiDkuO
sO4pYSGUHloUQxfs1EdeoouIhEQkOZPsUfwzEh8NiDBtxjwRe1oSMN4vf9NN
/2msDSOOMbJadMKf/JEWqHAjWuHWDp5Ilpi+d1KVbqakuG++WbO0vIc7MFj/
kW8YC5U8KBYXCywadIlHNhnL/nYaaBZoepLEx0IAPWwe/w2tLTw2IgsXuWU5
GXtHWArD+89SjVhCbvnXAeG23LvWc0FSQaoescVr2FWhkqtH1SCw4BrufIJU
YtdGg09HnvgsFrQQpO3Rq2tsia5QlMgEx1FggZjlwXhBsT1kQZMYQC+DRkab
FIpv959mqJgh7QlM6MnNj4I9TueIhSLr4YZ/IdBxAu9I1fQukpkkfU0p5nGB
9ZmaydNjSpcITaI08y8GaOgoByReaW5U9RXXzjobHOLsD4tQdNaQ6DBEZDhg
rdYWW89EGzg/IFJLD+57KjphfvljBdOfYUQT1tzrVV7NJp57wVug18AH+NoJ
TsSl/ihQT+N3+1mFp64xavp9iY2HfwrY1Skf0ZdhUnZwlobi6mWxSWFwgjcf
Eh9npLtECGDKYWvIzDa6Hq8j/E9jR1ZVRRBvrFUbeMSB+3MEfAds/nEDUMzF
WnfgygSyZdokL4Q2oR9VjXoKcFOmU6WIPaIPXgE72rg+e+fzlXNzb3dmQCje
lSW4EzPtxIDrHEYkG1ZseK84/bR014VoXnrp4z+PXB/DnpbX9+K+ayG+AbFU
6U5ojXkw3CzWJp3VJuJB72UnwusvtDS/ELt3mtTczr6o/xgOlwncWsIyaBkj
IlN1U1+yOk2IS3LVX8/DcDdg5DW4q/pMVdvB0DLIKNWfcIsSKSBfSLYPOto/
FdEFd/1Sc1o0pA6KHCgakkh6oh2WZlfMUKH/OhCGRFkZwnu1jgHVFCQZ0rWm
G+09N/tdk/p7nBGkm+nqzxQDlfkFBJ/loWdbcF1snkKDSO6d19JlcjZ5JWkE
5IeaZ5vBalksymnjiLXWAQp9yG0FeIvQPgPO0k18JMnpflnfmkqTHFiDiNlF
alsMhLQzDJQjXPWWzAUMgTFuVHMd6Vi52iUKn2ApxINW1GjTmKq0PuaLclCz
ivZZOL6KgHcWBZIKVTdVSJBAZrGgIGfOefBRsmjsUKAl0hOEyw8dHyvAJPr7
K32d10+Mih2ovQO2dmRWz+ElpBJBvFRz6jH2Fm2GnCPPaqayz9hV5C0fmUG4
BqJ0bQTgZ0bwJnI6AoHigWY5Hy2oV5f3WnR258wLIWhIUxnodHLULkY78BeQ
Y2EpeUPkzJLdj6J55Wox1jKxUAmxv0x2KOlmopjqXJeaFhqSk6niBXWtvhNR
V4CXOU3aRdnwTwRwN8ezg5nQN2eyuma3c4Oydf6PIJHAFaIC+sirikMtfeyK
/ecGlO6UiMqEywAzMVpysCPxrNnTt4OQxqNvbPqCJ8X27BVGuuex/0J1mGvN
5youHPTDkpGzjCz6XSXP+vrszgWbSwFpkJyMHCW7PUwQRDMVxW0IOWWiSUaf
S3vvpclCXvm/i4ci0e0gHSuxXJYZ3BrdTcwJMB4bfbhOBoc0UEK1kKON+zyU
P2+AqKebwe7TlUFu58PXBBzgshML/GNdv+u4yFzq5xR9i6IjFi13W5RiZnBh
vKdoP9YpKCzgGkvF5ek5VrtA5XFcCmeXUUhqCJcM9q5fVKENg8jvW4h/TsLd
dADvZ5uwbeT/i84oRdUweJIffrNgl0jv+/qOUMOnff+h64s4kaS13nEqT1pP
0yV/NnALdEWTdlEh6zVnoaXDWPb529nM8IvwdtRP5yLKWiIeg/d5pRryylD1
RMNiB0cdUlpsVMoCiP9bMRHk21uroAGoT2hVU2JUHo3OGFyGfgsL3r4aiuLL
br4OH5WBIOIq8Ntzd2vohYwerktxHmMRBmR2FpEEki+8c7DiGOepVi7RExk0
OtlzkTj5/rDA6hYpRIuE5uv4pNWT1saQ9EUVjNwtM+K+VaTt46d+uhyagD3X
sdb60hg2bcpIe3zU4iozgzO0jxiKIZ1Q6KivcR1qR5+OLgmC/o6aV1WZ5+Gi
0/73vz5epyhQmFwI0BFnoTgLM7+DPv2EJjP/WoibmUFLjZwQFkfoS/4vN+RR
cl8Dc2b4OtYIEOwPmTDo1W8NDnoFQtbzJDFX1mI792/zQ5LKVXtuQp0J074u
RujrHFp79CeEyxBG1shLp6PIwo1cRZshz4NP3pn5O/IWEspL5zu4EhETLiYY
fd4Jz1zfkUdCutsGOPQCtBtAkB0R5rL7ZX/s7kdvn34HlwsGnbtKpCC8MaMS
EeSqCJ/wIXdEz2rw0pRMErbSEfHIdh1R/aRnM7qXG3Iya3Y9+kgok/JSHs0b
kqOj0EokYeIdv36vpN1rh4PHdG6wZLFiPniJE5hsu1Q4Z8bVXAvNcfZUNLRB
Stbx5sCVosESkV5nMsBaAkao3wRluCA0+SP0Kh4O75vLoND6Qh/93EaYSYoq
3Xt59hsgrEn/TzLcyETfpd2Wh++i4NfW5f6ApQnTWppOd06vvBQOuPNWgKNz
kQR+MwDVEbJStIPekNkNOPfq0z7CsE3R3eHUHRCI+Yn48r8f+VFpj4HMft4b
OO/FBLdp4gFC4Mp3fGBgiI9evCmkPiQ8aloHkQDpPCs+zwU7kKI54QbLnZb6
e8DMHhf5d3KBBrTIZPWfRvt8JPG7ewDxs/EsNLIQYRkvA8iCUQ4diRP+9rE8
siL+rWndyxEU3Q1dSr6calnDUXXnbwCLGONWnMWnQS+zjPOcHUHBgY5cS7BN
2Jn8vGflmpZPj2upRqoq2+3NIv6FHgS320iAlT4AZgXlkQhpzr9/2i6ovVoE
EpBDjVVMR92NIdHK/RHA49OoFVhD/2myaqOeS+yteJ4mKt2FY7CycBxVWAR3
lumjrEC89XW731qyMNy7YRudDCAb60t0BkV7l+IDXyzvkWpYW9++AShp9nQd
NsWVQypXkBVN0RNcjf1Uav3G7hSIFZIuJUbo5eUjuJXTG6ZlijWBswLEaLgi
pMy5Qk4HMV9GeyUZc0r+PTMlyHlje7qX1YQS3gvDBGc6jN1Ty7JWB0gi0lbM
9vTV0pYiNJ+H/Id4CaU95PQYuwMrSC1HNGuElWXmFhw6At7PwheQrIvBOEso
jDuQwNMy0AAej8oJCVdbIkt+CwRXPTnXhstwS3QivbYxyQYVmyyOgaUuCSHH
l8+VO1TkIR/KWM9a9AqykO9gkfuz+OqyECamwHLdWCk7UylSDPXJoUiQrdfh
APh8JKLYQcptcwtTWsIM8gZqa+fEqVTljA/nFQRKIylRLX8wQu32R8jK2RLI
KGPVs2RwTj3Kzu7R9i6MBokiXHHPON+pyJ2Z1aP67TgK63VqPe2oN9iqVKLW
HhSYKr/ytdxOS7qMeDK9i6lOxImq87YCUkzu67SK/HbnGcMwqNu0XBI21oIj
76BaCqusznbxA1hJi6tkJBTedKwMbZ79zymUfFFg/oAmOKsK/RZDuOyywofV
zlS4YoypYTxsjlM6e6aYb8gZasYVE3TNEqvGngWA5sWQaGfH701zW1h0sM5m
gZOY8al9j8THTktaOncCmYNFrqgyRyml6ND0uCXUQeSJTPEovgSViQpU4J5E
VDUcqXown6mnRYltM9pg2o62g3M0ea80otsTuaOR0VUXcF5ZN8qP4TKmkja9
YTTfzudmv4/1uI5Uly1JFvAse673mhQl4McFxijssd0zujx+qYqr7zx0VgvY
D5AOYt3thm40CjkzCzZ8qNqVYMLlD38o+nunyBNyfYC1hBxwn5rLBDDv3CUl
E76U1tUfUl8ATArCcsoJ7//3a3bSgEztnRB7fyBZei5vQMem5xPMCvP9Q11q
L7EiMmd4OcJJxDWkd3HOS68xEOwhETJRUofYNce1h4WeMVKGwfdOqIm2AR+f
ZWkAHra98V6RU+7VTYq1WcQEp/BuVxaUlT/x9zPO3ANoAAc0AI1iSykWGU1d
nilDmgW1Rh/40RV3zEsEuyl87r0RrOPMEgUi87uF/w2libjs38AVoJD4qIe7
pupYocUsfqY81RhnwlzM26qRR+1iqK/zEhn1jfpEztX/18mrXECFSMJGEZ6L
JKJsHEiD6VyxEFwaEJh3CP55Ol6cJBPfrsVXJ+l92PW82uooE34RW1VF4uks
Eg7VRIXkKla+45ZoO+cYndYv74reWCN5ssCNeJwQFcKsz71QHZixTfu/Z7x5
pfdn1UYG+q24lySL/FzU7RRyCmrs1d6lRDL6rnYQZ/VDJ9wWMQYLZWXWGdsH
BW9IDnUxeh7g5ph93rvlxBLaYXJLRorrhimVnnUG0cJTPd0Psg/PPUu16Yk0
k1Eb+q2Vl6hwVlhi1cIVifPRePNBFe+fKh2Bsu6tzgnHFe3xd6XjCbRa8XY3
G5PD+J+wob47PuT8UmQGlNJQXDZIKuauKrSyStzv3n5WOO07EwAf61addbdh
aBW0NP4/S+JIRDUjcMPhtA/cFyNljFJTg1RoPXXogVsTtuI0q8a8gO0GlwW3
Jjo7L57fEA9CQWK0gMQnQkQviOQ3a8A4fh3MJX45AQeTIpeofEoh0vdwC/T/
ilm+dHnrXKwCZxG3qKmmxDijzC0gUEK1q5MFV5wYj1CaLVvYoujaUmZwKipN
62LtEpuOHwIpr410OtlkUZe7LRcdsj9df3hkRh7cJZYM7U3oFG4pHvKNopLN
J2MjCxErRN1ims+ob+oHYns5a0187kG7v39KYdugQ65egQPgSSFFnByvn+V2
2LbTEXkGzAA4xkNM/TRNDj9KU1cNPS9MjY7G96rTnl/LAYZgB/uxHriJwS1H
r7s/8EB15iV0zmMAXn4h7zz7hB6tMTHRJzqIe1z3dEvTNs/Y9waXtbwBV7km
NWYuBInVoajmNfj/L9SWinOeXUocc/nkFiyd0OSJiRsvc1kbb9Pa73Nawdjz
uDV+vwZeaAI9phGILrYilO3OdwR18ZmwugZPPwIf2oAp1VvGhaUnvSoaEbIt
ZnpCUL33V+TGIWVf7h0+TzIMc7p/WCDOkP3giTewjwsv7BZKQnLpZ9vIfnNX
Oq04XiBreJXgzvgpmIzbkdDJdzxriUB1ncbKqpCvx6a5JyRM8Ts7FWLS08mM
/H6Z6e0+S6D4PNgN+Zw0DLc3J+RA6xj9Bx6TbmYhgi1KjUjiYavP8ROdrGjw
oXmdfg91AEYllwmYwssXYOdcMv7jlXtZ0SsheQAOvt2zxs7mrk5i2OhXwBPb
GLu+j+pXeEYkyg7wMt2zAlJXloSN1MMVxX1Lf4ekuojgCzn8jeYbDLb6Loh/
ZhOEPt7xQCuBzeV7AzzosGYpnVVRPOxvEds9ux+fhmwrq6RYRVTUxz+3LV4G
C3+fGfmj5T0FnoBxVoDFPcOekqUc6IcyEgBq5dNDWyNNwnO5tYv8XtuYAPRM
vOpgbAu2eL+/HV7d9hPOHJRlbM7qMbvoXNIpGPFl2Fv8geJa4o9ulmrXyPl4
KDWK2ZUR5gsKXmM4bHlWQu6gPiVc2yM0V/FibTDaU2CfhFUGKQZCm6mrNucf
JnjiI46YMMqiBDPsSDvno1fB3X+6k1YXSLCxl/b3uqgVdQyHjpnU57tqkyvS
WUKczrePj9WAke3bvtMnLVllRgC4KmDEhk+Ni5xDr4hgtfhzUReFf1eLMFH1
+APshvluARxcg2R2GElrRlTGzCa70olpHD23OEefRgZPPjeDIkxtmp/LrR5y
YnfLuoawmXVLQSkioIZSJ3gaCZ3JAE4GVig7Sg2iBtnWCHLlABi4Jtvjw8LC
5vjCd8ZoB9CcqvwMRXMzDueo0zSQFtxr50fYnobx1AWx/V3bjMEaH3nSvry8
Vd9aN8Suv438nm12ZkTMNt2/TN+cdT6gSdiIrIrMN2vdlbcV8fbWMpSB7H2H
UDSY2Xsz4otTtKFVyDgh4P0JCOebRIzbzUYCtg3fQmlXHJtmTKdQAVs/dADV
QYP9F81qCWQA4x+KtbwoxyB/8Oy1FiKHr2uqX8aFz9yLM5+BRxxJJhSXoL1e
0Wc3b0ukXAlk8xyMcnOXj2FllI4wJVhOH+UD71/kJQmEncZ8ASuH6gsXfnfI
CdAwPgKIit1wrF2mVGzgS+5cgAf7IEGd9cqHGCIJihQgXweP091NcEILUAxR
L832V/Pa6xqBprid58EGkvCjOofVpk67KvJzylI3PQ3DHjqDZIWmGtsllRcn
P6NJU12lPPXh/K1zC90xA4yCyERS5kZxlYyLHlOf6UnuFdzYmCBbNU+WJSUV
dP4K0sd75BASh5ENZwGOmKmlqh/zfsa72DJYkK/1uBYgLBmzp4FmwMS70ZM2
j1lNEb39XCTFKjzoqKCHHefIFk8P6cAEJG9OFn6yllClCX12Fp88tch2B1lV
N2/PvglLxke2D0kZACUl1Iycyla/l5nQszGayN2Ta+DH1siXsQnajldVwEoy
HpZI9mRKyGlThZgiIVa41CvlJ4zckDfG62ceCaHKL5upBC5n+2xwz8TKbDsY
fTkCehvnrCKTmGDsMxOyijeiO9LKj3jmTzEmNuuD2KKFQuo9MYq6M3C6TfDW
57EIv6q7qnlGpaedFLcGgjBMJRMBcsZhs00o8RBxn5GRqBurSEFIQ8PWNSsM
ChLauQ9i5p8kXcjAxcsDhMFBYRKTf5UEW3CtC2MKC+Z5nkHuHP1NXZzbW2HV
OOachtc1FNw0t/DphD8W82Q+Qtouhpxh5FGkZZ7zqUwUtCesgf5h71updqxq
2pNjSNSLn6KJQ2ova4vbPhrcAiPtCzF7YSTrD4lXa42ZJi//xyO8TYsTZJ4C
T0okzbX9u2bfMWFVU5+3vtb7vTg2Ay4Y7g1rZgWVLUsSOUb2anmE0O3ujZzD
VQ4LeIu0tU+OPSiDTKvFqEaTsx191XZRYplH3IpxYPK0CbcsTjfhrZyCPRIj
OiVtSjB+6CYFAtDiKEurzkUpv5Yqf2I5JdBwEAdUhPCFMc7M18JcbBrEFrmu
Ht9zdN3Rn1rvo0QEI7O236f3O1pVYk8tDgAagiUiggXnUxiAGKHJG8q4hDWl
iDJ6cCc+eEL9ox6QZek8Zjqt3KJ96WG7wLFvfq8/Hd/kOsmodgoNwMbGi9lD
VMYz6qGmBumZ6dXCvOpRzKfq2MpqoklVw435gIgM3+yQQj3wBfTP8py79d9M
AAHAD8g22/68vY27kfktcTD63tzfz9v3bE+kuh5mECcJxyxH16OdG+niPWOM
TIQuGxOstI6aD1/ELxBPEbH8B6EUqK6bSxKCT8nxXJR99hmLukHFScn+RTWt
0h8Tf8CLVsfbGkX/93lCOaPr+YY7EDDONN1ceDCzcJWhzpXbs5DVY4pKX3ln
IBiwkOR+C7+QM4nUU8447mF/G3DL2q7DzspQagc16F2d/OE1ByrkYVwI4/6q
PhuTjhS+cWyUXH0UMs3dnV+oGITHy6PUglqd0yI6byxrDMxSawyclCFGP3bD
bQA1k1HdDRVh13kbvFiYqzJkVlzp+vUNhqCnEtqkiqJDWotF6xUnbhbTRK6j
cGlZPJk9NeJJ+k9mhrbakFwmZcLcfuSFPHKi7rPsmcd7DM7EeqOca0PKv4UV
AJ8OLSPh9QMv+/yhawI5VKePnGaERdhw0SjxSBszfzIS/q5roOD7IT0Ba8Gl
V/MOk0ZWOUJoa3yDYAhvThvqZz7KXrXHbZgZ+9aWjBwdaGVMLW5oH5rtd3SH
f4NgLypFx597J5qeLWOtomXJxUWGQyOYFqiLdJ6xS0nPUXPjpyGnjv1K1+aT
VU4bpxINistR9daHH1uSrE2zoyYg3J8xiZIPjxIy+6fmyTLm7fzoF7A6SbGG
0Ltx2FEgfaBUB7qs/dU5rgfAx/54gpBlFwAbATMTTtnIFFgujvTDmQEj6cDK
8YvSsN50YCiBQO1PWp0xSau9h0JIRH+5xN4qdvg+mFPGnPUaRDSBghTc4yb4
16JWJioaC5Is2XK2iitvMPIWdeMkzkAcTOWeW8Bvk43qA7v1BNdwQa285cBJ
pjJb9hxCFKuKYvHnfm9JTWIxkGj54915Xw+XcsmyO4q8iE10BDMgNMGdEveZ
P7w0LH4d/n8N8plXt4mxCafdAFyio76KqskRxGXUwrPaFWtLslj0sH1rASKM
IkMR0oKiXFBL9DoKeYsoFQGiw7KXO37Myt9KQC+nkHmqIS+9DYStlqYmFbOV
joovYnQCIrBoIFYirxiHiXlkhpzS3V3x7OzwNRdc72Do/8ekhSMTlvyCXMtK
OR/kLvJXpCL1aP8TGLFXMvmbg82d39Ys//JgRAmy4DoQuxKtb65hc5kf77Ef
tmTmZJE+b+4aC8REu/jVGnlOi9IPOvh4AVza7fegPStm/EqXvJ11prLb+z9e
QVSSXv00AxZy8uAgU4kZPCv9zfmz2W0KSqpj6JpbXQmBx+WZljltv9UH1UjK
h8vJ5/zQYFj50XDOuWgTlXGxnN30EEvCofipaOgSoaUKjXWNrV/30/czPlfP
sWAzp0p+UutyHQt3DqrwKAQd4m3c5MgNaAojUP0SNhmad9BCy1Y2Jl+Npwet
X9x6rgfbbnL2jhFV7OwuRxQnSlmHPNOrptQLLJ+DT74Z9rUHEz5KLnALda3p
Eapt++BsDi6sGLUInWsSeFI9AUUancOdaNGm2FaQWrvVH0dPm4GzpBI0+ISt
PMEvhCGaH1EcbT3X7EKIJTD/uJ4eyThnguunQL0NrwxwtBSNHey9d2hfcCZH
vYLcc5AnIq/juX3alb/2i+KIaQHsYwqVNkDCQzXOkG7wBwMS85cF8R4jTPvp
jLg3GcWg6aFepmNw77rXWWoDIxhmqRB15nYJADVOAO2PuXCH5LdpapKwBPyI
vyF4Wmm2E3iQVCWpX4Ps4AzHe0CK/uUsvsHFF2PcU9ZwkqVXKgcqHrtaW/5k
w5Rb1UkbCAczFvxZrDnDKb+skswdDI45bkikDwkbycKu43txl4XhSoBCYyoG
rXUVnmqkm+sGHKvub8QxxcrKffePXi6bvgiS4CDRjN4gxJhvcXm3yKp+MFqw
hp95ONzbvYexPb6bf467tqcgWE0hJKMgwxKOYmoLssu8aweKP7GR1gpP67RK
+/A181T0kE2N7Ygs1hqBzDd17sdF7nMZUHZnK5F19FcbuTDf6zxPK3lgSq11
hfI1WD4y7j5OZHSL3EcLu1se+LJVlrUe/LTdadN7ehJBzNHalZhqCJmGwemG
dD5fQCovJAIW+rXjabCAuNT3FkWgud2YFzPmdYb1mEiOcJ0OTN4sk4uybhIK
M6UldsoIBQy+6GQpgxCEW+SYun44ZuLfiUaGeHg0hlogPM8Bq6lhFjTu294e
7ykrRxxd9Wi9w7g1Gs4iAtzTix/cRiWnvtZf9+p9Kpv0eB5fsCIlhhM75/Bw
c5wf98jyyCt8WySeAwUp3GkTTb7uQV7do2x/V1pxy1XQkFbZI+WLRIv45sDg
/xPxRyUQ0Wr3KOnFZYEZLlOXrFjyro55N9ZQEtYgBFa4iiMfWpANt/pQ3Dbp
pExbPQO4o7AvlhzjuFM4+xkjipyQpG0wcV5FUd9vV45eI3cq0ojccaFwBTBf
p5vZh1SrUmbppTRPCAUOjVCK5g33KsVjCCc3GueVoB1KeFHUMknHwImh5T/q
h6AypZqIJzVt4khlYfk4ZXnMrtAKg/4/Nbrj7nknMo3pCClSY1sdFxq+s3z1
id1ChBmDN9UMFaPWEd2V0oDF5ruhZd7dzZM5VJjZadEXOpk9dDCKXWvEK0KC
sguEQFsoFmjF2y/ErcURbUsmPGg2q/qth9Zs32ibr2+K+iuYi1JlRAkve3sI
vN9ZQc3vMlEgD6A3ekq1+YzPX7vDefB0suM32TbDHcAtChNEnbX4dOhqpRN9
BwYrr76so21arICRuEpu1haKx66V1BZLavm0c75Jnh1FIWjmPcCvBeG0gaLt
IHe6K1/MpfQQZHq+v856YfNTJqIizyU4HXajRBaEihn4u7vw46SDcgqMe7Wd
vbjkSJyrR7LXshfitlsw3IFIMtYggNKI0+JkVwGOobMuv+r24cqRrtiigdt9
39RJ1/UFIV3ZasAzqv18IqxAUUwXvU1SI+KTMP2zl/xuTgwgPuKgk/N+R/cH
xi72T8m95wnR64wY9mKQSfq8rthYiZbNRUooXjBlNjx3vLYp+uOelWNi6xdq
HkVTYFTLE6eEKbs9Lo+oOPh0KloCH/NK6JOoPfvt0acgVlFjsHu9UYOzYpPc
5vwR5NxBUTWsxxXf3HpTJEe6ClVTVn40kRQ9kc+fLcQ7mvJ1sZWMqmerz6NJ
VE0c2jOHZOzGam3NJOlVNxKyXCd732XcGZKPNGdHu1OrDgRW3RYZ3vNEMh8O
i7T6GfvqHF9J/eiNSfvlJuv58Hj+7YxUTZR7qxMDkfIVV5jlTz9Luvy07zMQ
/EPJkHYJwdlNR7xTlnYgvS/3OoAHUR6U/cVOMGoHXb3n8fYixCbPyegeFBuC
/PhdpONcva2z5G+puj1Wjsx3nnu6GDKGAg304AsVSW+nK70Xdvtr1UIwSTja
9Tk8A1S2IbKFXxBAD8lbrtqkYqwURkqygeXVa7YG0mlYAwfiBywxteraPQAl
dEtLfhADwMFBmXR29u+d+CgG/8Y+tMZcJKsGgdReO+ATf5GlMPXqnUycQFm6
3Th+frIUK1UxZXGZJF6kWeqkgHtTL5aYPsdBLLTSjOHFaC2ju/4ZA9kI/Sw6
e9WIpuXWQDXCxLLItrS6RibeapcjtOOfuS4XQIe9ZqA/tyjfPG7WtXIOTIYX
uzZVWM4/m58A038LLoZA8YrJH+NCjVs96SnPDms3gJjtY7wAUmsGXN8VDRjL
8RvdCjxlmwAXE5jGgt0jPdGYncnP7KbGjfymGwg5TN+2BDYXXiKXlIRrIWVp
gTKUOVoKHiLkI0pjNEEXsWT3SXznfi0+i5s/v45tDvhu1VYCe2Pzp3nNdkTm
a9Hjyj+rO63tS7UA/UuYpEuOQpI84vt2jcDQU3PhsZuvrz73vjXHNx8KjLL/
2E7rwHhk2XFHtmJHH7LspltbmTd5+CMfT6L5zeyCshXVUX3ayyq7Dz65oNnq
M6X8V5ctmffPs4XVD1J5GWitU2vS3GJVhwuovRB80wQxRGwRfqpRI5ArxvPw
rlEMIJowPSWesympmTJ7YCYLzHvIJtEJ2ES7MkcvTiMprJSl4j77yTJwDKu3
ky5+VbovoltV7DQXQNqRlK8Zgod6LaicAxGcoUqt/n+uoU8zdFs5rgrczE4T
l83pNwU1dmrMieboM9GAaMnHZg3k1uVaLgFCMXrrUo13g5lDqyh2XKvPLfwu
DadsoI5/3sunX2OniY1xbsS+hdTEbWCX9sc7+A7BDHiLn+cWUmvog9e6VY7U
vxjzQ4wHNK1+eGRjvzB8GiYevOhCZ8HYlgR4DOgREanRBdRXdsfknfIcDt2T
4lWF9u81PKP4ijS5CGtUMb9fwWwDKYg3IQZmg/WNIS02zfHAA2/PdAf9flqw
rsAL4LWCC/0yXM6VkvJhFw/8PsAZy4DPfICH/5uch6LGcAw9gCMtiX6llr5j
V09CIJQs9H8PkuFBXLB0iXl6Xw0unr4EFJJX019q7jdUmbl19wSghXgO+nPG
A+1hpblQPD9PCcUGjwYMpD361bp7QdnErYXXUP5gktXfP/2r0NuLgpFvld9c
1hRU41w0BHD+0ZYzFRZrUP34XmqkMmrn8tedBhsUsiaUBnGD1TRtYIWnxS1o
oQBS7OMsS0JPnyrWVB/oaWmsHADI2Bg+XDV8Y7ti8FIbi4YCPwyXslocXrc8
haXkb/tewMAAsvGSiAevmrLjeRNLQdbIH0Ril0pqgaaKD2hkzW2HQ0+tyLcK
FIqsjUHNMeOIZfV4k8tqIjBwjjvkxF8jep+cG9fKMguZ05pPgQ7EqzUq4S9M
n5w0YZkC9rDgxE8WJKXihigRxvD51azEc1MjKE0R94Zp5zarTjvPdsrWB5Hk
DdlymD+wraqTVt/SizCDHaYYwJ+6uAuVU6e5r/tgIZGafNqCbRo6OP960H6X
WiFiwWEGLVyghAuEJql70vTYPKxd48iJ5ob/8ZbEK+sOc01XJdp+klOmPVkF
UcilW20yIo8laHwQuJesGqol0i7v1dbU8CQWzCAgEvag8iClo9yT3HRM14Kb
BquX8p68szeIBns8zylk/PaDOeXSg1bjbcG7TltGSQ1An6YYjJeoS0JuZg4/
ozMl4hQCn/i7Al31im9TxAK9OH9H1waHC59yU+nmA10S7YOhSkda65j4n7WS
8es3pxwzyEySBMVpqCm2jeYHHgxKAuuK5ZYu1oZq3hGax7k+Xm8O97ZGR88h
pQuFORbxgjHDioN04jjUl009p1WWEFwSq9lBm+mk2v1tdRciuKcsH+cfTSJX
oMiSCTOlS9Kp7FDkcPUJNffaIJ2j9FRLhT1UcvC/GPdEBrYZ0CkNK0HRHeNq
lyDbGpYv+J5w3rsnggpAOeVMdlqefxGCvrJzejSiV422buFtcTJp99FnVxy1
nve734F/0KAfvoMoBGx6PBYWxY2W1axvzJkRajjnqy9nPDux8kzbPHn3r8sh
BNxuL0M+YgoatVTK2OsbsznkbuyF+dRNnzmRNd7FysEfdWxdoYMuIyalj+m5
uv49bcmpVPA/pph1Os0A3GntVrGhcHVUoYVcQY6buS9HPo7LW/E/KqznFGiz
UQ7OUiF3ahW0EEO0ZcqzkHEd2YheCbGMCRsjKC6bTVdqApfwoL5Z5awfCLO+
vX1ua3f+X1XvuJK6buOBHy7EHiAsZUlogtff97C523eS7AXtoJC1nxO3+A27
2VcHcnd56CJt3EzmcYO/9CPbYleM0LsWlI543at2MOpQzaLGIwWTcIdUAWQH
OmOUv38hD5WPhQgdxP1x8rhidIg8YILVVCHJOw7Eb/WhLeo8JtFfzBotPWGm
tIZnxAHuyDxteRnhbbjs5Z7msJairsb/+/64+Zn7P4mhPspazTy7EA3xCc1+
k4agErFpBZEyUScq+0tPwpqPjxzeFD+uRerX5gsURn0TzMjSpMlAff7thPem
TnM0o890Qpr0qE/C+abtuzjBBgWG01qRpQq3EUwU7vlai4CHctOVisP6h8SY
DYx5FSZWls/OwQ+03m8CVh5xJC/lS85VLg9s+BM3ljbN0aqKf6nTJ+OV+y4F
XenuTQZSX42dhoAxofhtRj9GXG5aGRRldKg1RkxgQcvAb5kyXJ4cMttH5O15
KjkEECt4cvR/kTnuP5gxkz0pN6OV0yg03twVmLG5cQCNpshfTv7FmwVHv9gT
MapfZrm/VOlFNXYD4fn3p2tQ7gvPNS0GmDrVh8x+DyXJirpbXVw75JEqp8Uj
ZBpDY6YR03HC8Yb57285Y30INPbYLWAucpqPEAnBZWQBhVoDcS7OEc0BxikW
kvCb3Ibg2Y+Dk4aekyqMhPoLRWJACsye9fvFt4F0+0ap+Yv3X10xB7slNotX
+AThkhLFmuLtoTjSCLoNBbK+mqxDQ4OW3fpvdRBfMR4xMxB3XgOlKETHyY8T
ZyH+ZKi0+b7Okly+eIIDXwsSiE3M3K0czgj4oNHLJnsTXZ04zqxgD621Ijig
YHTX7E8cczzC+DTwEyVtV7XPVDgqSieE6r70D8pu/T12ZBaG7SZNgPdh4crZ
nR7zjEZqZjU1mqYgF+3y66s/22jGME6CuP08PakJs0H0xllmfK36DOhw0qi9
UtaGQEozFmygw2gXeDaJEpA3WVHKIi6POSdKaajfUf+cjnqALLKeTfzgX5fO
1d+2+PojwmUTu2LgOxKaBP9ulNNpaKEAepZnLQeqW/11jh3T+4yR1sYUcGZB
yI9T8El/Y0lbcOoJFL2A+zaosKcFeFH0rdVWaRvpLA5cXqYajAbKz6sTSaPH
0dH8IUKO20ga0mwp2580VLcuNzSig/aFE635FGkPfAZyAVYymHLRnkFitv3w
1rruMzHADrsDeNRHJQWxYFl+EFfsVAZ79Hvo8Tw9IyZt2tO/RAZZl4/BOw3x
CG57TO77SNjOuq2P+eDCzzFGUp2Tum+DH2KhzzhunEHP3jtLHFwSkFRqsIQi
6/QU3Z9MN/UdRl61tuDN1qGK440CDXBlFEl9sJ5qp96Q9hRmRCUMTCnObduT
D3EaQkXv7rB+gL+huZAIeliaVrWAfP/ucfNY+JJ7onLgZ8IWawI5i82Co4+r
GqD061QosMYqdsIQOGi5NHt5dB4WRp/l/YDNogLxf29riH4NV/JW2ewDTaZu
slJyXc/57kR/gFWXWn8haf55EZrp38dEM7pmSqGJs4UL3++CUgJnuP29cryy
76vY00Oug6vmYmkMzahnD6avNHB3540ZWsCzveCCvaNMqqJx+18JrxYqwP6I
Pk9k9dOQhVshTvkblyijsc5Zym1A9zd7nEpwvgAfrcyZD7Hc6o84A+17UCTp
+ioip/YHBacJopYU1aQuD122SM2+rPL3FFNTG7fA1L+BkVkznzGEs4MQEp3b
hDy0WjZyy2oHDKjtLQV68nEIdgi14d/xfBdgEEtmijbSKlOUVylLgGQ8BMjo
cFm9Xt9gi8jBCJpGHlbHQpE5CutyxiHVsnsk2kIDUi1qhZkIE+RJljf7xGnz
Q5BlvnhScrDd8fF+3e23Or7O80gXXdHGs6iewFz7bfm2pTnmACg5yMYqizAG
BMxP0Fh6y1lF8t1wgPx4ubUZ4J9WFWxY40cYAxos3D7GJJENImIac75oMy1P
KQKyMbjuhYvoc7bmRfUlttbqyiQIsM9SFyTZ2Mjime2WZCXP9gPxLrpJQNDv
VyL1DW9jXrnXp0mlYqYis/uxIKpoHyZ/xNWcVFVBW2HZgvlo5l5BvuHSC3M6
3iPeUx1cQmDzn9VZxggepD1UubTVnZLtcSLZbGSR1u1Sf/g71IxtOIBgypv2
V80uMNkSgdkipkuISYI9Y2qyrvdOb7HIJJOiy5ZiLj0rbJrltnyDbmU1K98r
LI48o7LUF+2SwCeV931Od/XH1lvm8vhQfiHQn3Gf0QONA5+DEBIKM5yM8krA
KJR1qliWfaOIjv5WnSmLklN/KYe+Kl1ZvCyN2wfpQorh2zq91Wyv7p2wz6JV
LsJvToB3eeMy7N+jB/Hq4WcRt3WQXrLQCtmdoR1NoELCU/DqJA4kO/ezw5mQ
HiQOtERWjL7Dr4+47QuB7gsJsKV6lgIVm8Ln1u11jGgR+DvjO20gr9DExmYq
CxOkYZVQ8E2x1AheRC8dIYZs/oDyb8w4jRVb81KW/4FLMOyThU/TRvUu/C7O
43KFwnW7qwKG+rQ4EoMv59+GjAs0CYIiWFdF1Q66d1eKa+bJUcMRArfwLzjp
B9yW6q0hZUiT+3tqnSLvS55FuFdpuCFN0j2DR0mHxXmNzFuZG+nvRhPVpXkL
fvPAVKZIcBbamziSY/3aBTCd/9hrFmA6eNKAGRi86homL9FLSmopAkMyYdaW
MO9PZ1tFpsQuqCW8siZdI+eY6+6pgH61SJS/kPgP5mjskUhdi4SiY9OzGLA7
4C0SODhfyWReUlY9bgu5YyrhCoEal3UPukKbtrqcs+wDUC3DThJv/ErzPvls
5/w2bRQ57N9GZbBlSyqs7vOOxusjSxwYPr43ZRO7rzMkwLFzNYFn8lCbKLrW
b1x1UhZtzz1WXDyRiJdYDz6luXYKaUNKPGohBOGuPJzyxxCJTjfTTPbP3JS4
xW8MbGxcbE8vj7zXgD3laCVA1vg6uUMnS9IBosVafoYZSQY4/yAnI6VAxP2l
mxixSwrfLqUVElM4i2neWaLM+u6ZwRkpgtqXITi3Fj8gtvRYQ+3ns0m5kW4Q
VswwZmUMYv27erfWqqd3BK33Q/680tWNtFlElCK3Lggv4NwLuHhCml8wUrxj
ZczSAfajeFny+NZaGx4TnyAxSdXlP3EHKk+qprrFfSXCLh2GDJ22Ad5QryF+
jm9i0C3+9Wr8KLHBDYn6TfaDrNqhPmV5ODgI0lkX2B/AtAoolSK8DbchZ/Ts
yIwA55Dkvgo9qwPUaZNH9vndZAfbQ+0QF+4tI7J2oUpK/MaKvKaJPdNFGxHY
CNQUOxMtptEu36Ai1PLR9DGTL8GyVLOWfa0Qz53cJaXn7vUXcTT7M9k9aQe/
WLul4heMeDv4g8jdak2+qApVXwMpBDE9SVJtMsFFYc5cEybR+NR5qUtDY2mL
Mqu2m1I4cI1wi3WZHsnH59JPIDHXWSKqI+nOFuPkmZH5Ykr7AUjK/UPszii4
3++6eVRw6Gzw7APojcDE4BV5byutQpY81kwbMeIFFDScrf6o+eTJXxuDsDim
ArxZMhthb/ML9qGSLV18mDBvDRgVofoQg1+7D5QMumaFAf0Usjh3n2T/lEQj
oieg/oXstMi2x+gvVYCzTRaCxdsrtXfdYpgMzBBIzg7YvY/DLK7MXrIgA9ou
pH8fJlrO5NayzTWjjFr94wUiyl0S9R1RfS8t4mES5hBXSW90pNxP5wht0PRu
pl2+ddytOBHMXfL1dRivabiQYpuEVuiqx372g9oHeTMmc/TXCMlc7T1N1vGk
LhAQmWZfxkhz5t6fgpIZ9az6GhdOZVga570rj+lS714gRh3YI15snk25Mq2b
toOlMOVUof4maz9ceyxb6snptnPprsJp4WpmheGSfoEU7pAsf9/XgFJmzyqo
Surbjkl5bBBhGlbT2TRxL6YxITQlIo3++O9aUGwfi3Q829cTq34yeJSuvLvn
stMSz5J/MhBbT3ION/4QWc7PVRDGIx27uZll1jADF+YCh8H258YgCr1KIFKH
fhgjahI5H/BeYen0wLfVZ9x6Xb13jDhmIqkbC+bgUUGQcMMwu4LOHZ4ioLn7
JWoDm6xgQZza3anehOF+5JKyzHBQ3FzjBpIgzJVNnn1+OilZiYNqJWlhTERF
UL5Yf52GodXxNCr564mjVgeRuJXRSYGTmC6cxgLTwg+Y0vX/NKi52NI/mzSE
XD4jmulxsd3pl99B1C8onBpbrk4/ss8HAPKM2joabACklsgDyiKDB5saGhtT
EtK9RI8ra0+8LzIQVxp8NDAKQjC5eKVFz/H3Q2CKU/EdHcKQ0AArQlI/r/4X
RgM8NNhqYtnHMPb/PTglEGF+ja8m17nsxam9X/D+H4P7QRA5B1MQLqc3axSk
d8McAD0//S0UUWjl8UAqyUKR1/MIcik4e/v84Bv9mSTtQuV8S4BgureaIojO
VUw6STY/eIcJ8ADklrBwwnFzlzP55yELc42dzZRQuFhtQ6JrEc4uUfccUdNT
kDooy8sRRRPgGwgxLF/d1PeHqW+20MX983JPnxpIT054iuzePO0WJyV7rSmi
6+xMINR0iRBMrF+h1gIjcV9F5IW7y687ATRf5BAupLxbTAJqHvFGiir5bLJb
/qQaG1ORkeoJcJ+G/gFZs8i2oan60C0bJoBjgTdezfjEgsNUaSxn+oXBmDxh
Ceys6pDhmlSRoe8HXasWavfLUvO0kEU119d+7AO89oAKr4qfyhB2Ryk2hlM9
L/jpsLKQaepBGTqnmu4V1KACudXpmyKTAgVMM/+T+RGBuW/8BzvLPvC+h3ca
tNu+4nWUzdToGqspJKvceyysCGPdMjUqdxmvvAZySj1NuxGq/+Wki2h5dqyn
DU2sMiShmDjq3/JmxK5dWsj2TvEz0OVtPMxw5xaM1qyqIsPt0TwAfIXAHHIM
AqJp/5d3g+WWdCkLABKM4PUc8xrauRHqCtkjIoSaH3w2Xb4mClzbyGJ7n/SV
DRGBm8gcjnuV/jSA8QPSqUB+XbqPnnl5yaq62wL8C4GSTuuZJLAzpSs0+eZD
R2RdyjGirwPcy7Av6hNoqM60OcZDICW5w5YwzYScuuQ6Ngma9UjjQATMMGl9
WxwqdKR8sBVKuq7dJ8emifK4zYS9L966lSpR2dJv2euXdD2NAiMc/uJ1aRtu
SdaNqyU4uiZo3NrsBWaPRHZjJzrhIaj/hl0/UtWTszuXyrIdm1dh6ojSEn06
K0j405Z3bYVjYguQf0FDCrs9yuQ0+ZaRBWDkHZWz/xOw6l199cbgo6aDMQDP
Xa2eRY0ueYZaUE6vM6c6HvyGWCToztyIpepY1c8c1+csbkzVd6UrVs3dgqYE
KgfJhiODto1MfWsnyg0nm5M7jHhdMSzCILu7eCIbwNA6Wvn07SxFIzWSKO8i
PxQM6+09hRLz4lEBJyZOqONb/5rXz3alCkY7yR7cytmlgOiITlLAenzFUp5e
of0yovMmVmQnmn+I03KsDaAvVbEUtoc4eSkyeh3DjI5pol1W1ylzPTjwP2yp
F2YPFbMrB/cLm3CInDOQ+TdTQxbubHQS+tYomdwqK6wKGfjTw4Mq1DAeMLsN
gz/QMgE+ZOJR41WTpTzt7ajxDJK3nRfUZFY2k2+KHr7J7j2yGfEEwLMqtVya
sHt1VTzFbsXdq5x6R0lwhUprRifHneUS7NJ/cokHV+MVdM80evjlc4IUl0uN
dm2e5rycUwg/gP3VL5gVWUAAcVQJn4yFzrfv02yfyZa7/jv7P2w/G+SCOKui
i3Bqlxe7rPU7R4r8T+QI6Nq2mY2Bycr/A3YmbTaXUP6X7oq7w4f8I3flZE76
JNY4Mqgh9yfaFneWnRZGtAuDZpPAGtNCU7fTSjxPSwWPWBjEANrqUTeZxaBA
Wd+t+4GoTtutkBn3f/LJccYcrDTWSO+KKIcM6ScsSsj5ikea/6Hyj0b+Q/UI
G8e3F1+uN1ZOht9AnaCmz6nIBgiMtZCUV3qoel+YeUCqfZy92uoY7h5smeim
mzNIg7fo/n5VD3xhV7NIAg6GnaROIVrdShIAuk1Xn0ml3tuzBcQYaVvIkFkv
wEVKiDHsBwY+iFvQ3b+1wnB8tvqAn5qV0fgrVzpoq0MmSR8sBXm3yR8/Ip2P
mEO7T3/SxF05AKsqDI57G2lSeRCCEcf6h22MzxyVwcZ4QX6TzDbIi/jJzZey
INR8cpyzdWpFnIneJ9yddKHMSl4+BJrvuTdeB6sDGngZRcZfrLKRSeXxCVv/
9JBy51ff/sesJg9AYcG09mEASSIbgXgFrEomhv1PV8fEfOIziYuqybofdRkU
WEVXt8NfLC9ppeDiZ5XnrfFBiVI4giZLuqJXPmSugtChEDczdYRN3OurSiu9
RJ4wJ3mWl3FgNup4rSRZpYS+6Hd71soKAe310ZGWmIwB8mPoyFQP/JZu5ADs
HNEsjqwNyn2p/7pil72tZ6/fK8uyW58Zzo8ay7a36RZpLBUSDyYr+IBMmbmQ
q76ct/wZBpNXxpa6TVHN8zoLfwGEqPutzQnCDFK0mog1phqfa56Fe1dU0guc
dHKiGvEP5ycMgUvDK/zjJuRvbgr6iTwmEBhVQxWnh70sKHQRGv8r4nLnxHrm
Itp/1NizenatQlExHyfYqCIwDWJJD6kjXoeI5ftDyRpqzdUL0FF9SHML5CUN
6EE09RGjqsE25Iwg9m1MSJoiP9pD+ahXf9mI8gbtebKS/MKa7x2IEJW1cbxh
1y1V8sAR95ADPs4SFjRf/fG8IzTOcanOyXpPrN4rSuiJzmLn9maDrKhxGLpS
tLk9roifW8EUTIW79BLpNXyVxZ2tQtIPstUe4IdvKLFr57TgMKmGoMR6X/mL
EV12kQorifaw5W67NiPaHJtATsmwv3yrgg9TIwoALL7+kuUkihEa1o2rKimT
KZAFFNiHo85j2kybDHsS4and+tq3l0troFGQEk8yi+QedD1zOsp6mg5rN7Vs
wMkEKueWXPxj90V92mjDyWE251WrljDce9uRH8DmzBtJ+LnAex58zfjXT7UE
+qbeXUfsbXMSdh+z4zPd/on85QYn9qcq12DAXN0fBAPiVZICFo5GR4I/ClAL
Fq1kNZl99aFJAuARiQJXl114OEOX3piGp3oU0XWQMRD1aF2UAdJ7/iyoBAwF
dJDe/zeSHo7nGpEzlAycKRy27Ytc/2BhdNDNB/MrKVfk/25tKGCk2x88UoFb
rZ6wd4Y/DnLHqrD/pdxfE8WR1uJS38ZUIX0dQc4ceERg37Hiy4j+uGe0EdTY
Q5F0uUqo/HuC81yL4ztP0ijIYfTNNGZcbbKDDodRMO291whlxacMjcseCpqN
tyJ+HBMGJuP5/62VKdl0ty6yfmuWcIThrOajOSl78MLbFZrXPzOsS1Ov8/qO
fSZHxMjSiMGqYQ8fR1MChZiebVfb5vzV4ZhFgcQPm11VSn/zZ0fNYUNBss/0
sx9Kr0OH9tdEPy85us9r/3SG8oFyLjK/nG2rb4kNJ6axckGnVzi+yC+L6bbi
dcYj4H+KPLk80xL9rL06JuDruwLfGXoRjvS4Z8mVnvL9o/TzOL58H5MPZXZ7
FC8QCpnEy0Bo/XhjvlP4mgzIVo3Ro/t1rFSG0FqHLjWtDn6mdmNb2+jM1Vx4
Uy+Bbs5ndhu6D0CllkJ1b3mhhQSQh+ORPxgw1SKVjsp3mMCzJaJWSc6wf+Tl
NNzns0OZQkwmkM24gzv+m281+187S9s0TE16Ak1rd1FDDdCdnHCGspX2SAqH
f6MdcMJifPVPayeTAO8in0Cw0s3GPVCSu4k5tKgS9dkbkFBfMNBSXfWmW/Qz
LRkFaO6d+3mM33QMXT6Z6oM3yd9LzpRK/vzKB2gII03Z7mVmB2G6NEXH0aYb
TkV2ZM4BG35aACiDW6Q54XyNtRkBd4Ccrh8GNHC2rI1y30OpiDB9m5ATjDgd
kzmH5UzQiHXq4hRvIBTV+lZgBu8S1wGxtRPtOYE2U8k7dAnp01YpRQvibcq/
dbaDkY9aeOEzZq1ZaVUZLPm9A6ZiOv3xPyihMuIunu8j04fux/ijdLXpNDWo
EZW6pH0yg521I+alnBoRmvcMvDLGKjnotDX1E39CPXwNOhM1soQ73ychWJoK
wee6yyP4cn3aWh5xCx3KAgIszwPVM8Wz3yV6g/1eQBgdLWSqkDA0WYqR90hL
BxYXnKEZiyPdtpqYA19dP14GfukTJmDDBmVVeIZXmhwTBe06lOwLZOcm3lhz
k1azSRQffDOhqTW6DR0S0zpJG883koGl0/TzCw0ASJx9JAZ38K89fmApex7i
AA/XjitwRbTt/SmtfsqUSneaznn1IvgWDdMnmySqS0u2Fyigb1q9VB4+H2zP
QipcyY2uaSAqQug86zdADSlIGZ8ti+LdnB0gZ8nx3VPffQUOSxKBTFfy0qcO
jy41mnpW7SYpwsSLvQihzYA3iI5VREXMBRIVhcFWkZHeZSmIgC4vi3IjA6FT
3Krq9QOYHbYBWAU6HZ00DtNWpgO1I39hQ+8OcQenK+FM/yJgtKULj5Qvq8el
54BxSyPYNmrIkpuOtPIe8Hkt0YH9dL1yTqpeUM+ws8cF0r2o5X8bxt/1AErT
ZK1MIIqTb1dno+4QID/F9fduFhoW6K/2uy0T7NkAWUFsderhuTGc/OrbBvIt
wwr94JPcJZ7yx/fFu3i+WZw/O6jim6Pdxxh4y9N3w0EuZnEMNLpChLPvnzg0
fPOsV4sy7krlRFrHhCd+jStBSD1nulR2WLjIosO9LeF7u5DS6RiZ57FT3jP4
Fyt/r+7H0zLkiyWNgrRDCdldpl7VAvYkwlpY8bZ0NgP4awwZudS2EMkFhF+p
XkZuS0jLmSZZnLaNv2MDadmtMJ8LIMVf3rzTlSXkDJtSCg6gzgwKK/2EER6Q
VarQaPkkUibcDSyTNbh9ElQxOwcZ1/gr4hOEwbV2zgHcxc9TUOBu6YPUugxS
geoSHOPFE5O+u5FroCoPlc0+2Cu92NeUw80LvD9qBUUCuOpCknDnniKGqBUT
AbuxFGy33CQckShhzFuwQoy4eI12FpYabDS/5UslMUrLmMsKGwGCnH6vou18
tS3g10xSPSZk+7UgDameIT3b9LAiy9VkchBRk/VsbudbinsZSDFBaW9LZ7s4
VB8x9tOFch0pU6zKfzvQX4/AahukmIFbxaD06BxlSlAl3yiHYfvk9Qehv+gv
1itqGT7zAIOf9YLzGe4bZus89ExfAsifVM3Vv0YRc3e5rVbt9bIMC3lfEYMS
sA9r7CiL+wrOAQdMOrNyLJiki82CQxtmRO72ym3+QL7yxblaEfQI7fSRC+Ua
Qzx0Uh/o4OOuztVDrnZ+oHDfW95uMCcM2CSzPMjyYUJ/X0UKIoh06WVI6FKx
1hzHKP8ginu5cbKO/moMVV5xx3GNae8hxqmblsF4RxTDA+95C7g3LEtcwNk9
ZU8oeZwiLQ+xUD04Tfp0Iydkt/l7rt+CkAjMEfIE72K2P7T3m7QrlIEU3Z9h
dQq6mbFBk+xJC19/vKtjRzlAzUhN/b5Yj3kQONJTTz23YemfDgkH2uFNpeqQ
5DciwnP7J8Ym3fZRGGwwFfOcgVvRf/zgAS7iQmwOM6Cn4X8FiECEpUEEKHkv
sZInVUi1mR6Mc3JZbjvrs7f2N/xfyrzj3UxFUvVFBKeJHCvdW0PFkmejdKPh
zkWwADx8F36v2ecJgniJl3SQyPrDLU22VPm2WJD9O1zxhxrt36sUJhWJzr0s
XoB5GA6BvL/8vHzem5R9pvEE0cFYorBX8UlGpIYxy19nNyeFBDt5c2ehX0v9
sRg9K38moTyjLXsM3LoYN0a2TaK8RFUA98kJkwlzyQORy/g7WVBRRs3WJ/HR
WctWuk/uR6uxblFFj5AhP9PrxgwC5pR4SH8RWzlA1akELRi9eQq5ZOf1BT9l
UgyutomvOq5ckIOf57PY7vmjde4wdDr0oFc0GWCJU1gzqCBVx3Tt8YxvbWFx
vpz6UsCWDTbar0VDVTARYz9G9ck78QPwG/04ENcGdxLcaO6xPwgquGJ3moK7
dXU9+ivgPR7o6KtRbm/U8iGZX0Wp9mW9QHD8u2JO3R76G0RRJxVHPdIVz5TX
MKy8svdKYWlX3n+Z9Th/kR8PqPMD7fWXH52UjP2nNm8AgDkGzXUQyaAeQ4FP
gi4tkiR6Yn4Yp4zYehMyNiJot61AImucJR2sZ/F/XwTYRw0nIEg1C0svY95Y
Fc/c2m6xKmg+Jt+lxu8FhDrSqi+ZvjgGt2kH7WUVW7yXBD0tK6315jEMwTcp
1Ik9nMYExH6VgMeB4WFO6+7P+ekL7rt4dsClXw4xs7wLo4mV1B7pHxxjzhbF
Gkc9n18TQgNkZPDhMdgwWQrrppcj7DKfzNlLDspZ+CmxFFJE39g5JSK9kmwE
sAqjmmeLcBFFNwiiULZJrQYbSFY2Ljkmig+5pkxLteKh4J3X3HNPxToBys/j
Ko+Poyos8OTJrLPSA4A6wtoP8mUTVaTD2QUb1togPk+dfeC4a+sQIB84eAXd
Opurjrb0wBxnltJUjkELCG2SPSChB2ycA+GI02Xf9VFgcIxYdIqxxmQ/vM/Z
XJ+SNO7VcUzpvdp4Jt55p0FZOfy8QsOxahDj+F1eGKXUkU7sR1hPJZdq2VgA
Dz2eOepzybOKG/jLe89+Io2o5n4L8JKlmEyon9kqIcxvSzyKOLXVO2qKBoHY
84KRGzQa8THUJ3cIoVVbjlIx4WZGlj01aV5bFPKyomCyqUMwsD29zbAM5HVO
SWW5rMmuy+CxSErxLMqBzQD6hI+gDm9QeLnJxLJ1I9R0d3cL9G4RZQ1Nd+l+
VsKWX4TGW1n4hfhQWuNdpgSLd+DpthKRsHkr37kTgQ7pT/iHyrNRTrD0/uuE
XETzaPKsuvX39d5pk/6bFMrWhB7ncHtnsUepNaf+pQ+a7seFWcGSB4sSSdeX
ls7BvIxHi2Z6kccYeAT45oG453uZNLxj8CjkebG1pDLAx1gBZAdwi6OzwVyW
SnpYXSphDWyChJG4ei5E1ZKcjA6Lr/31EwFcOwkQNmnS2lAjdpmfQPgh0zaN
PiOQFVYwlbsU5UJqNZNUKT4M541oNGHHiJRwd8azx7Td62zDTkVxoiohFshz
a3t7Nlqa5sjvmWLkqcPMf82cph20glYs0ZinJQhvV5SXbV85h80DkHgbycVJ
hBHbMZ/AfqT8MGD6IFlsbn8lvNCb88rjXM/3lmerymyGK6k3JpTdQuGCheq3
OQK6RUAyHG6J3sOFgK8lZssqLoAGjkvlQQc67aQdPFOCs9TBAu8xnRQAqBAI
lA723tDNCbryrL1mppdRojM5MrcWiTAa75fAP13i5tahrqw3qnjNby9aYIJp
R+eksZdPtfGJM329WKetaARVoSM7wrbt6eOmzKUApC2X1ryo2+bvak5Z8wkj
eA458iHN1k4Ucrf4a/FkCoJkrqVQOOZzaU1qLwjVTX9jCRdEAqV5Qif9odfT
Lo7lS94da10lvyIb8DK5L09ibC0aeh/QhBAdgu3KRdFcwHXmO1dkwXtqOVU+
vM8EW3W3JMX43opJHONVjZGStaIPFjVoYsAYL+bbDb3nTEtP68QQchuTkZC3
DcYTaVzJuae8sLJpKtTte06FXA+1rpwOfySjoYgtB5bi+/6O5a+h4M2AXpwE
uDMoTqgvQduqFhLYXceHgeqaRSw43nrv+D+J71rvP/FAJEfJp999Rvq2kMFx
1nke6QH2Q88pnB1X6A/sbE7/H3VURsGbtVKefu35ZosF32IoF2EAENSYu2ht
Ju7C+P8mkGS4XzaHZ+MdgTVEJrrpqah6CTssuqejvXwgL1HWxzSlfy9G5qwj
/8EkQ9gQDINoICWY/NkaFLHUJULVuGaXAtw25B+I1QqG1yloY5+3e+IxGOPQ
2wEVRn+QONtk8eyHbLqFN1z1KB7oaJVp1wViOr0OOBOvQK/PXT/gY2+8qE7F
bL4t7KImeyyHlZRNTxhsSJSHPeAj3CPTIDzzM21H9d1CxKac530pFz1Lo5Ng
ynzAmyt9iabQIHZUO8NJ+CsrMd2KV5jusqibfrV1gYJMqDOW6ajYNYxv6qmB
JILOnOSBsnV/PpqJOERM61/j+WxpsWfrer9dciVnJUdTnkxVcSiNa5xxh885
A08PqJbdJxuxZzw4XOrONTfFk1vJZzjWJio5AElm3y/3H3+J1crSSA9cKbGh
RkEd0BtmKTIfQ1PFER1dnWSMA+LECIhUp77/Ifo/f652w+1XHkmN8zcLEEae
3+U9E1Ao/6WDhN9T9rpAxN5cNpSmTcBtBmsh7Ment7Ppav+XpsnwT37Z18gp
pU/XtB8ELuYERdwgXdYX++F7veH4RwUUWSqoOEL/eXRxE1yOC+XXzV0cbax9
U2KpPlf2//eLTCJT4faRMDN/0kzqA6XcpgTLhZkHuE9h5YKZrNNnMkKzthG6
QaRzVujwQpA1ynJnUq7tnvz4WX0ZturNXdzxpYUZ1TTaIWmDCPcmQ6zk5kC8
KfI5orTU+3y/uTvDPRrUAT4H9c0mtNaSMAvnZysvEUaHFrxfAXUKiOdUSeKy
sp5u+P/TjbxIghlEFHviQbZaKzoKIyGHDKG9ffFeumGraMC5z7ywtMhtCEXp
yf+VhjKY5mJhMSKuhpszq8e8g/yel1Ufq6H/on3zlnl+bizRm+SDw62hZuW8
EUYm7OUdyq5RJtpD9vGK+lI9dPS1WdsVDFOlX5OyKqecHABIDJNAj5OFZlq/
hhwXGSmu5NPS0VkJVuhx81kEOLpz+L4s1FngN0gvfk2ctmZ3QDNEoZm7KSsE
bc/GG+d475xE/cEcxqbcEHzgXsDoCdqaWcGEmo01KwmSr8BSnv7UlgdqC8Q1
DRLK+cIho32m/NersBs01KG9fDA/zny5x65sjAX0wH3gVOgJsEuF1igVKUFG
bxOZV837f/i0i6m+BQYvuY++USi84vGxKWImXWjVIskqBX/8s8WJ3zXEVEg4
YKw1iSiyuIcaTrjjulUp4pqJ5ZbeetjPCqO0CnjarqdMUGR1zFqb1yhCKoVE
SoKiz54hO/RXT1z+Do0oU+vmA+0pvEOocgBwsw0M65qRNdQsRVZ7Q7izB5+F
wvnsM+WDwgKyXJeE7l9xOhq1xGsprOtR4C8gQcSyPhK7JIdDlYL4z9ONkts6
jaJAlx14xvI+TJEeGQJwLSNIgFKu30L5oVjWrQXoy/iAnzl1BkJPG6bYrQiD
2CtdWrFg7FuJXJ+W+WtbZvl5iYU1X2hbUlB5mcM38lI7ozKJKGZ3sTqvrqxX
gcSXgZAIkXarPXUjym00xvIAn1QXGaJwLkvyYIw2SVHKR6sA2ECaw2mNO2we
tsf9md1TElE14Z+ljeSQnShXCEeyiLXXm/bMBOsfmNjMqdVo4TqK9k7RIj1d
+EHRG4IWtq2znYbHMrjESxAdDT86B0NbDaO2tYeU188fXEFzy+zz+fWC0RSz
4/YiqY5zehV0wShdSgHQKqUat2BDRMvSAxt2LRvV5gupV5tmOBHtg6xDihuI
6XIGLbFyQ8I7SaNa1lClZlef9WKDA9dZZ3LQxpUEmnNoiga6lm/S51fheDyD
IwV157pVKFg7J0L0orYJFaSJGV3NEWHfxFbrenbYjxHRMElmgTZAmvdtl11w
F/mslIP9nU5/isiriZgAEf2CtPGy3ZVCAQdoYebnr2C/potTKhLN4caZK28Q
6Wjzq5UR28RjIXmMBTyNAkeN2m7zt7f8Xlxde29ei8DjhpEkf7F2UDLrhtx1
L2YqqGhQk9O8I0w82Qyyc+N/VqJbIsao5J23y8CCgmUONX9xQuBqUS0er2Oc
sobtPprQXexOO/uYhD4PaoSo/4oxOt/BvrspAC4fTnj7UsHWegdfXI6sUgRF
o94R2urjXVMNpc0Bgg18i2g6I0sHlSG7zvHwaavydpvtPpSXd6NxiiKYqowu
satDM6tNn7CSNYTl0ebRbeEfgW/AL41IX7AChAqvT3UCRdKgHLWqB6cEHM+0
GMWE0mN6gkuBkJ7X5O3nms/ViLKBelEEmWdfnYP9KHqbg8K2QF/DH3w/Fo06
nmejApWT4GZUPUnmAuCfFFaoVw2h24GjcCoaJ7aktYxuBWypi4iymiyKCPkT
+WVElc/hlil127MzzskGUE3ofOfzduYhEW63Uw4Xifel/ehnTSlBSxv04IbC
pqKfddMNN5LeHCM8QXFN4WljtGWaXUrsB8CFlK3orPpCrXRL8IAb+v7+B7kn
fsnd6uJXDBfwk9vXwbA/HgG5PibVadKp65tkjCLS8z1cU5IMdOBrEhUc0tyb
THnk7+4d4ehZ3OfnY198K2D2bEihPhT0z2JWtbW815EfCSTKhtJXv0neUw5f
BBRVphjuYDzp23zyTbDMBzRJYx2+4orNyrERAJnMlD3/8nDVnoxAynZnKGPw
V5P4h7jRMWl78Qx3BtSEXniYkiZOYLQxNXWJ1ceKxjSc59heIqRUW0AW8n4i
ucdGRtwIShhAvjQN4PSSYJdN2CCr7jAQf+vUyZDHwdEJ9+Cu0IRx1nKW9t6q
3TcQ47xbla9jlcQrmPa6MoV90fWAvjwYb4WVoSlpnmKXN75aTugS269WSrI5
oYsFuajmRUtvApsaCrG+7jTi44FaE0eeMHLPW/Ri+9x8SnOLanB3FSfN/Gtf
6DU72CPEUNlIO04G6CHlUe4mxGZXr4Q/8rqOayGgKk/ZOUtl2HywjyhN7fUL
NTJzdCDgjDVXXIWZCbLaF7SzHizlKflRxjmN39dEWbb7QHSupi0odcdgYs9M
dufKkFXFLDaGPSNdb35u5ImolxykoOJegeVXoXqWd7YZ0ArovXvafoaUngKc
qPB+JFVF0jjP/XR9KPoL5c1QRmiBbrhmwdrsyf5cJaInLyJTg7iFYE5c57m1
7RrWppAYcQcszPyEAguVWmhONMoLsDhpPTKu3QgD2UHKX8hbt0nO6LCXUmmG
Wo58kyW+GKjGeH6ovhkUt0toqa2hMI5uepLtvVFD5ytCNziEQafQxgHGknXJ
CqHzndDsZ4FLXlTBj1qnefFV9AzQn1eSuSxARfO2FhXWdlYWfyUCnft5TK5I
8VTTJ8Ux/5vbzLj00/pGnSspWZ9ziXupyKgH1wGQn7b96ghlHQvjeBg0Jaas
1X0DMPvyP9zbZiLhQwIABQdVZycrP0muQo0RD4LdP3ypP0wsshtn8/CuM4ho
osg2gnY+5eFud1u/d5KHc77CCSq3KbI6rQuR98xvGeyBgufrXSZO9CBOg5Ip
u4X9MQZHq6DQV3px8ZShq6VI5nQk8RYUsf9vmqfxpGKP/SMlhS5DLNs02v3M
2KXdiANLZrGgR9x4HHSCBq7VvShhYQR/RaI5FJ6KDfx/jQlIl5I+bWiedx27
NiKp7wJQ4Ak8dPmTTUcrXLj9Fzlpz18QGx1kSAUYfCB7Wswv6iOhR8Fvr/4J
J0wkF0OBwl+b7RGLxoWjPxaqtDIsQxx21otJafxpkPUKgdULS4hILvudvoLY
y3orD4wuuC3iS+SHdobvfmdGYusTUoz2C0FS+2LW/1Zs00I5/ve6zzjL3E5U
GIQzSwjb7Nm7Ytcesc95A4YZhhtS7cU4pSCOJycqi8RTWqikuW1T4xMkvj6s
jRWo7ZanqQ2gGMI8ZcXuS1Lgox2hYnQcb0zfy8RIXRdnV38A38snMTZ+tyjz
iQx8bagJ8F7IeX5y9BAQi9ts4ZLev56racoDyDxoDrcEozT/46onuHzs9aqa
JsLFyYHjfufmNlQgjq6UwVkg9MXAcuJQGi7QX8oXwdq/V5fO9OWaLzwFcyTl
dndIsSo+hxAPYlG+u0fkWzx9hLpv1WNF4U6DJtZDSF/8klvsdyJAmtgZovMF
O4tDy59hjlsh/bnJUHOEIImCliW47cI0/odgNgAu/SVAfIx9meOCiVhkAZvW
6+ouaCn8HoJxZtRQHnzHcufVo+mIRDY8bTmiO2aWksSfDTrdP6YVUZJmZlDa
sJ5+TtnstNkEJFuOeDEJVjA8QSMgrR2hd9ICnYAAsrGPWRjmAWJjDuvmILGL
JGXxa68cA9MHQslBxFMn+CLqx9ZHVF1OQ6imXObnlzD/lutmxfMs0G1TM1nn
szntMUK7dKFAgUcvgyb2G65N5WWwQtJBfFIOOEG/SksUHo3L9qjzy0Fj0BWY
SpFC8f5uOTFSGzRsgCqzxlXY3JKNo1O9/nErCwci53uFjNfE1o9u8cSVV2pp
knZ3Z9YoEYbg4sFEVKhMIbNls4TxIVqrSK/m9oy1O3XLt3KBTheO0DU0njIv
Syacoc68XnsOP2DQMJ+s9DIOwN5Y6NO7SNKaQLrFkw1fdSOymUHODrqoU01r
3KX/BoP5v7psxQ/WdeAEeuQNiYW4QEWR7y81F4uQRKQiF6lwyWipDwF2//d4
KoCl2FKCt10ejyFrUn+4ms7xiKTAe0lAIMlvEpw2ifGgjPxu/qe4xBCiOu/w
acExLqbpJSwXJsdgrs5OzD3KXMpb7CdnMz6IqKUzdosoPp2LF5oErX4MBWVv
oggtbjWlhUbTu2Ch+VVcrBOme3sgGp3sPqssOeky+WI5/eSZP3Ec0X/GAw9J
8SfIFlGxJNe4o7bJ2lp7pHFdUKFPPe0xmcpL0awJBEp50yBrBb3hYnBnuTMZ
6vXh3JuC4ulITcSjrN3GuqgZMzd37D7yrMdIeF8KV6sykXk5tl3uFXeSQw/p
S8H8ixKK1UFD+7H5Ia6cSA9CfzjlUeMLbrDKXTdieuRoiUWHmptfnwp47zYh
/fZGXIU65O6LT/92DAn84487mxgCMkhzRT5znJYQ2TQ8hPh6IwUwYd3XeMoI
1hbrwKsH1BQwe6To1Ms0Zb+LebyfTvR9vLGTl7EYY1qJIx6k4xcconSkMfK3
QFi5smSwWAWxKLudiIaYoOTWb+XspnlFBnYrWzaF6u2aCNOjVckmCPaERzYv
FGt+UYhpOI7LDe2PMWkvofo7Wc1RkaY38pacNa6W7bur5icwH/ZV2Y1fat1Z
xP4QoMzS44hyqdXEMtfBHnZu4a0uhICaXxrEhRkxx8bOd2lcI0TL5fsDx3Rb
sekR6AZo8wllD6HVpvTbbMbwudEY7/s1YyeTjYMoKIqWmdd9XQBv54fUyTaB
aeb+asXWX3OVkxUrE2vSemPXBeq6v5JAN1tXksjx64fdrbC6RpNWTB9+aVKg
goelQwNv9aJdbVHcc4GsnOWeVk9NCe9iEfqzuCWEGAesU9GMxUGX9ByDYko6
IGWpsaRl6TZF/kJ1cfUNvRgGV7trhCt2Le5B7b5LjqZnpdj9n4ydGs69Vixj
ITTBZOVMpfjAwKttfRl1CFSWspu8KzwKkSTuWem4ICGre1Vs2xJrQoE/OJs3
KPJJNfwhbU2z/+da0f9+pntU8v0tNJHplZOicKPiWOehxBG2rrY+M0tzEPF4
MuASTh10fA/9JiUq3xSYrReBSaRBqJDMyeO4O6W6iAlCjMpZCkwWx0v850T7
vzNbPiNQO4s9g7xmNvvNQf770FbQ7aV6AqOy/ZGS/gPcdwyZkvEhNQZrfTOu
FMAIkmP2S2K5FhIgKX117envRDEg6Gr4jAcnWB6DHBYsRYv+6+dfu77kpqfP
NFm5kteoiGINKopaWozZBpjTgAUHsk5SOrdr38tRbR6aTcvSj02lI/gGKYOR
J0CUg6Eu87OGpNVTBErmDeKsOWwKlribxjwbxHc75Wi9EyordqXzWUEsIdRk
Yry4Lc/4dwh7S+fCqbSRGA8DkdI9xf/ccwEHMqIUppRgq4wJwI9o5aHsUB6T
tTr90lOF/zPHfp9YZmbxfr8ROeARQcjXYQ4B9KPt1/Xguieo2411+0exHbl3
BdevEOmhkSzH9e7wN/fEOIxsCWiMBA8s0nVW4B1fiBwA/sloYnc2zSg5LQFW
puF5J75GaeEJ1nnxTYjxqQW2y+JTcdewhLtceRMcGLxt5siuTJhRaH9SjQ0C
yR5DUGDDL4KdJBoKw8+ehhGfUSaoktg/t4OxeAYQtw/YbZBzppVgFTUo4p8g
3RiYjQTpKZy4mJro1RZC3XaeMQzeTOoa4Sd/4M+1vyLPpPlUhK0FaHSsXee8
tjTjlvsXrhz7zBx1L6mImypRACp5veGf0Sn4UcBuGzcT5bPQ4H9kQsfLO5uF
DOp972C9iFYYfDQh1EhBcnYIrR/fAg1skdj6got5Ezh5hUoEe4V6PInLpMw8
CR5NCTGFMW/VlLTUtABkKCqF/zpD0+F6vXMth7y8Dm6jqcbFLwRZzG0HTHPD
tfkeNotwe/PHAlWKlAU6Rgai7onSrkxCAbqRlywxQiYD1n/0dZTJ5Nt87NLw
nKL0sBznL2ocWO//XhC+drBsXo99C7I1hBHGLywRuYaslCUB88KC82oz8djq
SxCL/UqTBY4NcpavfFN9OR5uwT6swHX17KaRXe8LHdyavwx1O2QjTklPqAen
wVIjAIe1OPuJyaNaAW/qqzv5PeXwnKZe6baMBSNKToudboiBL5ZyoOhJSyKH
Rd9U4j4nupcID54cqF6S6+14X7PvyoOCuQeOMIqobQQR21sXpJ5J0KH7dBD7
Q/Kj+NpZmzp7G8pp++/DWNZUVoZG5FM9p6KL9YIUR8OEFOEhWrWvM7CVJPIz
krY3qEX7D2xtauV/CO0Psk7s2Dh7dzyieyWscc4eHtTNljl9Y8dl/j9cDNT9
ZOu0aI938NslEgmFYTm6CYET74TIQzCJzF2joEcufXhkoHYxQPMlSpX7LHNS
VdWBhbfcOcf5IjkbZJHRMDAX55udSx60rqTp1lsgT5lm3uyTzuXc3/hpOVsT
sYtQchGCmeall1yU/pykMiPCxxaqlweRvFh+Vt9yhxeKi5Dg04dej1Gf2hI0
wEN0SLGMwEgZvzwBLg/WgcVM35f5qt2Y0yXGeSwGG8fXUfPer86FE/kh7HrA
CXq4x2HgC2jEyxBNsuD4Ohnf7bc9MNo5A4NHnnD7hnlmmR2ADbohxWJtxvK+
o4UV53bJGnwu6PE6KXeJoefcFIzYq6j/XoaMLTa3DEp2YEAxmZT0XJlH4amr
aAN5P574mF08cgJbWfzVl5XD4Xa8RQJojQJ9F9ilfnaQhARzlSAL3MXVdOak
DyC3hxzC7fDsm7f+hlCHWrIXQKByRTzEtlFt9R0uG7iPKlHK0HvvyD0RToPm
lNNNH2KiNDVQE1godfsX21rxF66byNZTx95nrFbvChI2hSBrHS7YS4U/s0I3
XXH5VSmbiH+1TXGCe3R5w6+5B18qaJCdZ502kH38WC1rHCuEa4MY46r4Oibv
efBiS7MfzyISia6DbHN59Fg46VJSCMFw/Wy1eMJSwfUb9EN2rzJivRoI8m1t
6zutyAH6dHiURRabWW4Fo18Mhjm6s1yq7WaTSMLEvQxCX/v/p20gImOR4N41
NhMUxEGQmWMuRD6Vk4vFYTuN8GzxPG8sCDTXHiQMoJFjZ6C9mQrfonjcwq7z
471P29zCrXSMulibqmDVz67RsQxaL2Z+C1lb6g20FrqLYt+VnpR0ANf90nCd
nkMYW/e4fmc9jPisOQg44O+oIscTS5w2tp/bWNbZj0GdbbpcMRhB58OoZA4V
QZLb574YJy/Kew0HwavE8I8IR+DuQ2CYDScYA2J4mtIfSgG5WX7uPMKGh56o
M7Y2LeFUqhSfcsQMK/TsXdNL9c3fU2Kfe4QMw6jZ+gdidHEuiVaRkqMIkCB3
nvFyE7C85kj2XztTjusV9gaE1+7l3+ZsHRqukxX4ZyGcdrgEbhDUCu494PpJ
ves6mD+cB2JGUx2K0/nLjcJ2jvTt34Rmg+sALULgmhBTAiCQAVJZBGCnubz5
AYIyUig1Pk73ltl36JBqkoBbVSJJvJUeex2VblI07I+WYQLLehuJYijZqLaV
CE/RT9OmvsR3P2bxAPOGYNLrkpamJ4UhgIkkFz4mTodm+hyvHWjH7QZnPkvT
RFzXE/CiSbHqme8/dYY0m+vFsoabFGmUzQCJO/95gHXsIKvAl9uhHgJY7uaI
SrRpZaoDtZ0hPVj1nVde6jfFtPMa3kKXJwRczCKdF8mSdwilw5btQTHA85Y4
5FlmAASFUAjakJzvUMir8R0xhHFSbwZm+RF3kLnnA+WRENL2t9OBdYpTc7Ll
sma5NZf8/FmoNw658qLPvWqBZa6ia/g64xioODCDTYzPzOvYcWzjUm3UyhnW
UjJqVHfc7tvwmYf4oU7cFaE+YmJ4ayzesxlVf0qaZRoZcfnfIvd+6I4ZDLEQ
5o/pZ2YDMRPeJI2QQehbTEjvwdOCeUuHJsh7YHTmNtFqCYNJdifsAbgEO1xC
cGGaVnxYcr9rnqH9MMdjJBlC241om48Y2rTqhKk29M8/a9jwIkDcG96+HjCS
0kHYRPJ8dFQNEcPWjNHCm4UZbw2vmhhSs4vi60RINifFAyG2BgvqC2mRAI+8
+fxKzA5eJ/Fw/gO502XrIpSCUsFzD1y/kOXwIoLNhpe0X8IlYzfVMY4kQCv7
wKZt5z9B8XwILq2qaLst5sFxWSPAtegFApSsCgRBUTouT6bzyNKl4ZiBJ1A7
03Gn0/5cmBjlO/rosr/gNy+TJDh14QcJi8kWGbFCcxRq/V1wbGhQbpKEF3NT
Xn9YxclZF4NiaOXcI/bxIeYqp4++L3trRQbWd8/9W4wRsv6Nh0LHzrkeEO2M
N99TWWZcOoDyrmwBoMaL1yOurm0ryMHg8JCGM4i1AVACuAhwCGxKLMgCZF5g
M36p+mnHm+ubgh0LJVoUGL13rrjJLEGvMdeiYVuURl9ADfSWhEIovNTb/UHb
b8Vyts9U8Ol8i9MlOLujnHFvCCoz9nQBqK3Tb+rfIpVbW/TverxvQvHSaICT
kMIWI05bWyvJTE+1cd1rTXYF7DVL5xeZWqA5CADJG01lBKiziHgRX+WqmmYC
Eco9wId+ffWjPCvuClmGHZv1o1Q4nMDzAP63mP8fHkSHkmhusAM+v2wZlsmD
puEbtOUsftzzFPa9qi+Z3fJ4aVsk6EDJZx4/DyXF6hc0e0v6oD1Ihgwrg3uN
wAtdrMglVAFy8eI7xpOIaeSWw9pSy4Cw3/WmKoh3RCROlFcXUlRH5ffdrhqk
4FwL4CrUgNEPIRAogeB65jJU2teha64STqu0SI4HSHWny1L6B2zU2uRpmbDt
BsatSVrN+gOyMuNUzTiCFWfMpxMJ6aaYGhAmiMMqhlnnCkyR7s5Bj4hiiNMr
cVYyN8aWXezR0axWmOx+1g1r6y+Atrn6r0GNKlabl6B8qntV84BZ8f2GQ9kc
i59eQ70ca6BGROGcD6oKc9AM+bvb68YTOfpo+dEiXMPUPxd6JvyPRmi/OMpi
s/k+ERniHce5cZ5SMNVxSJTT3j5JLdYTS8p3xbvcfcDLH6f0FeG9aRU8aMqu
tnpUHKkuwQ5WAOhxiSEtx4S7CxftZfDtOAxEtEKPHMUUuUdthdGXbOn/gxd9
M3hWbmHb+MSUSvY+45+pzQTnmeELPQHhBZGFiZSqAj0Bcc4eqWrhNUZT37CE
Ck8C4cQZq6QmLCEsqGvuZcWZOrO3Bb53RIvvaVtn2IoiulIKPtsgBmIB56kG
31vb3Eo8cZQPipgRKfLXK92TkP2eqARvBaJXmtojVi5CYqx+rcI/HxZ6QmX3
7TOgqod9LcRc3PAgm8KiGJWc+uZQWkLCSiSE7kLXQvGcDir87r/xAH3nns60
9d4LMfLvOkfHLxdGql34vpp1LiFyG1LUaYRd1nf1m7PP4/u/qImerqK/VOl/
c9yZIJZaCLdMJydO5tqOYXZp/87BAPssvWIwK3q9PJddn4gPcuE5HSa5iFJp
u/C0fPwFu1P9niMKu875r7usAWdFQp4lLd710STDomxlmTWcaGxnyeW1PPGq
flUvFuGhD0eXdRhf54Kj0vo5/YrWTtY6BOO4TJTr+akYrAwojgNpgrOqkpQ6
nvtM57ZZXAEordYacO3X1sMk0CTvQ4TZe8HrLVNi89o0sefKYG+W2Gj+10P/
geIesyjMVW7O9FjRs7ewXkeS+mHNC0tsBj8Df2XDx/y6VEPDO8j7DIRV73bZ
20nGNfBTNht4gfZ19FFWwTMwDmKdi8qJkrDUBtsbug1cKJlQ9QS8rcN0wfY4
YMI3RfA5Dpbd+hyy7g1MM57CfRFaBz+ECnwbWgNsKQhQiB1g/kxKZrG/gZeL
lFUDLMsoZKSras4xMT6XDIm5bkLIXV4scSzfBBdx892Ma5yg+eP6Qm8yW3Dt
n6e49l78EF/pOcs667bhxDOIwYxER7apkNdOmFZzE/tD/nKoxL1gASBEsYfa
w+LSTbkJnQeyVjPazqSlBFDynU4SW3LSLExIx0tY8x0YLgqgbL27FwXmMzJo
9QAw2JK8HsVNlhUg3albCKl7OxcicERSr291Naj46UrM1loJWy6G3Ied68FZ
3plVP5YJoYcivBVcbLbEZXzeWJFdW1x3vcqWNwu6ZrLGHy1rSBvZILHoCfoT
qoC6esO62ytJp3LsXQZ3RJ0usRdoK7lp96SSFf/d3Rnt787PUSas9w9h1KTM
2XsR33njGKa7sScuRMTIq7uAwfNJI5iGZdoCPU3SI9ErEbyvqEaFGVxGlu2U
k7Mr7To+3e/rpWHGwcDGZDL+EL8PhtY422Leg6YeMm5joo1HdoIbgwPMhikK
LA8hOZddPeynBCuvp8PvVnLYaMz/ubydc6XnGBfFgJKJBSCVkofHJHKftzW0
rQGcRnlZUwMD38rmcKYXg97S+G8iOKbMVxC0eZjx59Aycr7+KSjPgBKu2b45
ciqeHO2WUHyl91Maagsi8qSpVijUfywSPC3kXIPsWq3fgB7GBPvEHJDrijF4
xDMQDGqK9a96HPqZmeu7NRNO7zhRwQi9g2DP/n6de779r6mRwgEAlhSYHuZX
ShYOC28vaAaPrQQE4mH6aC4itWP+FVSfZ1ht7TCRe8uVQ1ww3LvEqMoTq9+s
qKUSr91wxv+MsiJw5bT4MTwTYX/A8BN1hpofZtjOT8Qdx97LgcuPbY+sACii
Tg8cs4VmiFRJI5gTN5Ih8dfUw+wcITqXWhGuESjpJiU+d0GgqORDa47nYIDr
+VvlXLMLc9ItPANroQLy5W8dpayBkm847qV5gXTKflVk7kaH6RCk9J0bq6gE
Jw/drMviWGJb2+jfb+AAPvA0JB6GenLvomCXWUAndIgnuN7OOZwSLXQFZVLk
ztxrfC3RfWGk15lKn22IYxPxOgiV3qUK0IGZdYiZMKZxxJhmj6MsL6wte9nh
6e0xvarT+dtvyw3ysrD7VmF89nwLoFLL+1tC6GJ7ylF2leNASDApB525hhd0
1T2sY32a+DI2om6ZG+uQDN4S7iHcTV9mNvoJAuJs3nl17O8/GFuEvaJUHIxG
FtDGhVKOtwTuIxMG+JMFf9dTs5sHCRogqFUY70Wp0acqtVJmZDucbdHY8rCR
m4aolOUJGxRzGuvQenc6QnwGV2YJ5LEN/gaP2AiUhLcEy5gM+M0xW0N+nKuc
pRgYPV+93fWk20o+viVOb3ngnpqgIJgbuk5e6ZPooC9n4RymiEMqOJ6Fw03Q
GgTlwQ5p5ZwFQrxN51CpvxZPUnxTQX5BTwH+/rwRi4p0TMPclTz5oBBlsF1q
t5OAWF2vqm4kzjxcv/E+Pspbus7X5OerQt97SLZaP37/rv1rANEq4ClD+075
mBQQHLYul1DqJEx+IMQVmvJZTtXNxVPPpEomHWZUW9XcjHVra4uJ/T6Z6mzj
xZW33iriUOjDw4jP12nY5CZK1I8xZclHgTGOi6arGY1dIW1tqHosxQWMDfZc
4Em9SW/mB8mACQ9o3bGlGZhOT/sHsxfvI4nsBaBEgKdKYm3FB5YyZSYdO7wz
t4Sq4/mc63e9vS4pCD0/OZ7FD/Ol1QDW6SWgUPZ8RnNRP78e+6GIKp0AHZ8Q
dyork6rJzE6kG1MKI+1zChnLby8kLKZJAQmXXTKcWGskZQRITWTby4SNfWLj
cgx3dnrHobu130X4PQTD9U//ri9cqTMJoFiGuM5xA18X+P3qZihqLp8yQSoA
7hSCq1B3udlPq9agKFHH4uM5sNS59bo0AwiEY/FAOLtyDb+imv591wTzSoA3
Fnc/RGPyp4lwlAKFliOGy4vjE1EqNpc4S784amH7Ncsbnc9VhvceNWuq8/4c
ufEhy9bcboXvE3JTFTRTei15v5t6DV5D033L6NLG1ExG1x5iWXeoM05B7Wm/
mLsJ/q45byAnu/tDPpO0pRgu76UB8u3NLBpc6bY9PsYW2VaOiqJ6lcoDVwOX
H1BzkAOTLRUZoj8tb6p69UVLSdp3APi8/G3Y9pXxRwj80d7NeZrZAjV+RA0k
mIUSTREqJz0J+L4lgbLIGdY/PGkC39LFMhBGDKFQjrqiQFFrQGOS+WhhmmBg
vJLbDgtHwoIIjzCx/Vj0NOgA82j4bgW3/6Ly/5rTjghlMpQAwPeTwd2jtxOg
C6H59Q9MFmyR5RRyGW/TkugCfve7eycuOn+0yNzwnxZbOci8EZCbuzcT2rRo
s6GEMROO8qcGrEnmL+lDddhlvA1E+T04LekHG1fEEpmxIteNIBSE47fEjeUr
dhNoSDlsDxAmmtLievYbKFEzd3IGYFEJn12fLi1KFsnY3NunPedNTeB+kgCv
4J39AGXYGjx2utRHZJ+UNhKThrrBzBwmCleMi5iAo3Y78zLa7YP6LsF6OupY
tIJQaCIspGqRJHlAzkJVNfQoOh0cqnq4Qf9+6EloCytex0b6ufgmQI9Dhskc
VDHGvqAWkqObN/Rz9KJzt03kkcf6iKtkeAWq6rXcZ7amnqROWAr/OG2Hd0w6
G0mxcTEju6ZeYy0ahqwmYL7spBw5kAqDqsi2bWhHTIvMCeooRsf7lxQo9pl+
VP30LyTzAmwyXS1jH5FM2agzxqJzSEJ12CnnLnoGSyaNnGkwEiA9qY8JtTXe
JeJ9O9q+0iWse9QGPH3hg40iV6vSScD7wbxPWTina4N2EfR2AoTg83PltabM
jQc/TBdEIhkeFUF4A+4mbw4PrH9s9QuAdmUHy4f/Xt7XeYhbu4PwnYX2qK7g
yqFW4WJQcc35ZpgvqgXxxZD7dzcR4UpxssEjYl3c+5pIqInc/QRIEZnRjcb9
9cEPJA5MeQsVZlCkY5tm02uHxqRUDT9BunHfCBgA5LSTEmYoraWORTMAdkUe
iHE/XGf2OheL94F+T8aN8VP895XRL4Ze3u5U8+5Wi9/HfN4ibKuI3P8SBpkj
LKId+7VDKK9aS0soYgUxl1hPftsZGiYKZUEmDyvJ8c6zl3UxgxLZr9dxBN9V
La2ZdhjjZgS5D6r6o1GXTxt0YNEUOCVyfMBX9MAMB0eujkMf8ulmnl0GgR0i
PCFg5ChPjLyveaa+w3el3TFwae0TNf/2BHmb5Qm1gUcpnvwQOGBm3SPSgLbV
1h+vq88yFSZZ50vKej89xZZ4Bq92Te0ChXHgHZ4ktempxelDCEc6+Aa6Fw7L
DueH+R1OeZs/JJwcFNqcvCRObFv8qgitTytUmySMUvMt6tCEmjrcir1uoIQb
xKATodoTT2cfq1tA4MWqv1i4FakIQ8c4p/Bw9oR8N4EwyD8u4vh70cM6lSSU
qTkhHJ0cPhaJ6ouvBin2MpiGNn88jSn13XG+IFbYf4wZ5OftI/NGmbNsaZxZ
q4eZwqTeBOgJsHiMqT6dx1UapdPRCmhkltbNI6IFNfqqRqzAYGLIKCBQXTM7
pAgUVWBLJwgR2Ds+4UvcpJXYc+kB5wn3KtFKzdky9HPO2GKu1eudVTdgWZCJ
zMkdqm5+w/CUGH4KcologVsHDmJxBSHj7zzRK2QWdMcJXsQqjdTJR16QB4gF
3N1ejnXZlQ3q3YjGOkFrz5rO3zoXnpvESOXIaqOOuYKytpAWIiNQ5NLrS5jg
AcmDrTa5UysQdMzRxAeCKnRYcLc+/MCNUMzQyQnE2G0LHuq88pWG3ZBzZHJA
zHNskM+oSn2RBg1IWiYpBr5TyI6fpeRZwigl3xB7Lmi3+JyFHXJRj9Vy1IS6
IAyDFLgNtjcGMUnRDNnqCvus0/rN9m+mCcGA2mSxZ8/CS9ntxVHm8zLsCjRh
4EdLquGFyxBrz8mWBpotG0kp6SuQMOzdGN69oGOLUmbjWSVTrkTigg5YQSJ1
tXNfTSVKXGA3SsJaMfU2P+I4IW9w8xLh2gybMiW9u4lnmjR1rGUB9yrwhlKq
rjDGR91FCebPi6GSVBXPpAwQjjkL6fGWVZkU64lbNL8fJdsTUoFfn0hr5zDE
8fjxhOTVEzAUCBBCDBaNhHlENrbzDIBV/SdxJssJKO82h8zvaggP/KCwwjBQ
3FcnpGcYLSBMSKYYClpS408pCW8P5MQi054PJyaVDgq+x10HYWWB4/Gqkx9/
bVWoDhHeIF6qTfnKw4brOQKGwkF4QlNDkt9i5B15p5CGhwa5gYEmJ9Zzim4x
6wmHnr3GWrFlQNo2JAbY0W0WoeEfIdpVj3T1Jn97P8jFBtUv4DdT70OlXgug
xAiF3hSf6MkjUAV/78pnQ09Og8VctNI2wTYMYd7npVqP46o6VJi0RtT1bqjc
25jpT3oBzscRXVXVeJ8MLU3qDXIFGqgdRTdO6nDlwUWv9C1JpERyAlzVx4S2
xH0H7cN76eJNK/dTsc2Wjn2aoZUnR8+AMiGWirjQSHqa2eQI2UUpJj1naLUF
cqBWTB5Bmyf5dZUL4a3/ezLrrO86nLa54FdAjPImvaEwaV7MV6wbYmj/sNor
BIH9G0OqyvCMLlCxH3FX7Ta38ozqFqcBNQOItmq08SuNSNawHQWyOcgDV/Gm
qDHgEK6YYjTiygCZ4jp+RQyD6RmGTa6RyM7cuHEnZE6y3XWiPbbb8KFuTizM
RwMVTqOJskpIq6c5kk8Cgi+P4nJroao9e3YJpfRCfn+vVNqXM7w855AgttWf
+nbJqwwrtzQih4vogJX/HwTK4J/vTWKHfobGu96BPq07CiQNJ+altxTme0c1
79huGw0R+Sn7UZpH8I4WbTGm92qWEB1+dRFd9mDtXuR7vP8/og7UZu2ZecGN
dDjPpDvFSfy9LaGC6TdBBeQ9ztjj2F9f4GlxCeST8nV+fNSzuzTBEDeRRDkA
CDQ2tfOpbdKjZCQLKa5t4T02P8S0P2O44iBHskDwQBLnI/L9DR5OfNb5ATCq
sgaaVzuAg6yQn5Z/kG4Miqsx+ihXLx1vAvy5M3C4bMQoPzWtInggfeprgVc6
rKTHD+dTSCbe2YH/gJvbTYUKDUSVST6rH93utjZ98KVTAmw7AuSKWVErEU/4
Y+rkPsgNuPStZZxENvDup2xs2nsZgu/fxngmrrRyGH9QPLKND9wMFrEzmwYW
sS8+Egn3cGlR829jtVJKDiFmrlTxdtON33gewj3/8F4bYtlC3HjG4mZDi8Jv
F9eQlbrBXWMd0WmeFPkpEnsz9MV7OE7EhAd92BHnSbFJ2OPMlEUD5IABss9y
/VoxF4sVfyAMn+nixmtWCYhA1aMT6sYmiPlt9JWt0KUVrP3yUdsLIYyuoHTf
ByvdFf/BWqHwlBUf34xsYxtpfgya2S9I0MnH1rZ1yOcFMFZ9fhZXkuojOuPc
+aTVP2zSS7kfFNFAJoH+wSZsEdDtNXvwRCuhgpejWiGvsZHQQ1dtxC019STu
4HlzZdDxKIWElozWmm4l1Cc6Dn181uqef8Ue4kiDr+Jue6jT4ZAPU/WmPe2g
iEMirJrZOmfbSh7/Oi88Xgzn0qUWM07R72GfiDqD8z6X78dBlZt2xtSvxi5Q
u2xb3ojr3ybov32+tT9j14vEslaejvmEJfWRUfGagmewnhYW6pdlb0P9ldmJ
l8Uw6R66Np5f4Wzuecvy8s2ZAYLX0utZuW7mUtQQ9LB8lGByFR4kUOsuMAeG
hwhQyj8mfYyrlRYAH5JLbglOWBgYL0kA/CxYm31eiEidiCrXv2h861gLgxua
CFMxPhue497VRgt4HBVbU9VftjD9Kr+JJgKXHdMMYTknIl1lMUWHBipEPw+U
RS1NeTBLx/VwCiFBdvbU1mu5Zz476M9vGPSyNpSGOCYw3F1eaxvLygVicFdk
/4pKPN8mwKpKdxJfuUuhW8Jnk9Yw+sOWexM6/AYsdsk6By4bohiC/ZwFgOta
HvlBZua6GIqpoFV3UTdu/Wn2ZcOIhlPTcL0v2bXNpO2Dg89dFe4LLN2mc3q3
v9aEV0GYA7PWcLdE3KZpoRcBRqynOf+bV7OqqZSTZySh6M6QkuVDvjo/j35X
MCsstNJHsM39SGRmHvXq6IMPtfvu290xRPQ3wfM30KHaUfgkfDqBZe9WVee3
lzccdPsrqmtcQn6bBle38hg2DgR6R3/iOCWcBkW2avhwXzC8/7KF0hdseYpc
K/Q6GEcp9i5jgWeJjnwV3EZIZ7g3VZ+6dhaM7+lJrbk5efqvtJdGDItPjxYW
7O8M+ep+QCQkfOaRaAPqhI5zez/EX8wFAfRrVn3gBlYR1+SNN1VKcnMBdw5s
lWPJY6D9AzCZwOVVTmnWz6khPrWC/RkCTR6wvS5U3hKeHJvTfA2Catb5dxYO
5fIZNXC2FoypjZUARagvNjgJiZFe80cjpp60UNVL3QABhAU1GPUtwAALZGrZ
J9nX7sa0ZXun3Te7LWwppTRIJSkw0AFMgjBoQOgWNgjiSbTPc2Dx2LwuhLdZ
Yd1B7oUa9mlR/qu0hfWwH/cdZ+PN1Br6t5wIWINrcvhGLrbCcJ2oTsPf77mm
8bkAa0y+ggT0+cCOt+8+L1Yy9TukMklBLP/XXhwdJG1wbV07tYIj2JrlPQ7d
vOIc5YClnu50x2RuRlCb1xnl+xiwEggMUxqMKp0EuD1ScFrOHNDg83hrluXT
wRM5Sn+sd6WZtz5PD/lnSzyELhKN8HhVGWRekQSk1XVcqoViGhWBUEGBHhXK
FvRI2ZGm7V9HHlrj9dfLOqxJDA6EMfUleNqhuXKlpXCeVVVgB+NaEf7cJA2h
tcPEXOHk+zz4sx7Ukcpead+HBQQ+CAlDYJksxPd5uKh4ZvMII+WFEBAd/kge
85UmKZqBUiULN5W6toLjDRZR8fn/DF2/4NRyoi0NmfobgXHQDpQ1v9ouXaZS
ohxKaBGFMcKLWpf7A7bkivgGJElx9zjfZFIVurIdjF/kM5RvXtjFLdkp/CJI
ONv28MxjyEddmF351FgwDnFB2RJZJYTw2S4wj/cIHvcFM6WEEYyyCA14r9dA
ddstJwlLy3I7oAo/vsSCLASlaK0idSRoGjAjs53Ig0axbqsCWN60kNHXM4kn
WNJsBnQ6g0Ajt8sPZ0Ehg/N7zcPDZ/Pd/19cgScmqYKYD+RQzzFiDbrik9no
deXqpFDWorL1opCv/JBuyMHxh2IhgM/TtmvXb20ibA5poGlix0qaiRRFYdqZ
9ai8wq54EeNMABJFCBPXAdkdsIrzCAzwRQHSjcuYx2h023RZNMIKLZ9AhTTI
tGmg60iTl7ZABHw/ctRwiiIwcrccwf+HJ2FyUWTKfrsP2YbDa2/N2veztXED
od4TH8GwkH4dy99VhdkloP+A00tr7+OMBBpdLTUzuWQRlLQkxv8fB78VDVIu
SIDWl9ZNxB7I7h3Aj1EpgwmOMMX7q/Q1fYdh5RaD0XX/oRb/c/v8UetaEun+
PwEq++liRsqFB0vHQz8uMv5+uEqMWI1jlS/tzi2vE7yPCv/7TBMoEXCupmqr
oJNLoFv6DEy9oSq0/lhrvi9M+CMWDU24YO0+4+DWDB1nI8lHnnv8GXu3kvaA
fO9Qqji6Uvo1mIRGFsGRRd9UcPtNtKTTKccZRcICcGrIohuRaylskmoKQNdW
wsYoLOACVmwd1hYpJ5X1MsdWHazi72cVyxleuxf4WvaDl+x7tIMyZPQkP8qE
pTUJyhjsg6dSBes96O7EIqOT/nWro4tL/+Ddi4jR0izSGjo3EoQkf/1sQ+sH
MhurX54FRzcC6e1Qk675guFDvNpmEO5KqH9tHyZ1FZyEEvYfaYZYKnbT9dnh
W5yH3avYg564ehgidjMyQo961jTRtdQt5h+kK93GeX4RN3cMfz4a6YX5VE/Q
ZjWEXm5i3f06iXRjhwZ3lNwxG9aoFZVv+y4au49uygjaTzIJ3BoOBaZdTXZo
YU/sULkRr4Senp6z6ul8KNUOLfU7jaCxzZ4eIBsQ73hTaq20ikCt/cKo49Rg
SOGnL7DddeucqaqQ4q93RcKgdrrf7Ng1xnjBssna1NbtZ5vuCI8I9/ab7OwU
qnChjLLaucoeaIo9APfASWwwlgqowKJvym3mM/UX1XyvKYAZGKkatC79waqK
PWvH3KxRUNnpRwDpN9/7MRDaTXiLNAj7O6jZk6aqIVQkpCbJln2dLKNtc3N7
qzTafuBhtf7WZa1/xmbWaEzgFRXUmKIHs5p2O02cWCOpJUGy/ji+xnOXwtYT
dn3yrmi8Wy6lG0d7XjQN1L1gT8qlIj8TQtI1ASuCyraWCXiVD4CNYb/sfQ6U
wYnERizbZ1pAZIfav3RCu9rKFcP2/8RB6OVAYbFP44oCBr34L93ZGZSRv4/0
A5CB9ipmlc8QnweoMS0rOViUoFMa2CHfsmpTBBWACqz2yUttlJwl86JggUZV
B+prpUGjyxShn5tuuGGPvxVBBsWf/aFojqKDGDYKvxFTD1RULwt9/gc++oP5
1DP0A9SCdfBlK+N++qbJrBs0Nx4C76wLYu/97eSi7u0sabCH2fjKz1aRDvId
JcI9i+KOjrvsNLEt624Ah18QWz6VHaD/aSGT6H3LSDol01pgpT7xF/SDReBp
9qrf02n1W6luZt3qb6K4xHUyguol7KVxfFdzg2+ZutX62unQd8KzpnrLD6+V
xheNdHeqAmpEilvsUr8qbedjeilux9PQ9IpO0AkbMa4u0ZXtC+xzXbY2NVOV
CM0zzgOjuw0ydQzxQFsHLRETNadTLh6j5JuHj+6sEEgkFYTatt2rvbJFf0lz
iQVB1L+0mO802KCv+o/wH9FY2236SW36h2mCwP2rCvzvjkl3AnyIQ/WH93rX
oqJQDcsMLx0Ih+T6ylcXUyr9jeIh1UdJ/r6fKP9Pnbr/XHprMckyu696/QwE
Z6QDNG3UtAimjO+SbrgTyD7sXPXsCF8NDaRJsIg9MmT3Iri1tHO7YaToC8wj
kHEecAFtQnFEnHL/1fVdPUt3Aqzru9G4cNaLbS4qQTZWOQdCIQSV5R317T7J
FR4lTHdPbAOP8Oz42ZhClH6FXFGDjmJ/JUa/cTNgT0ZtypvEqApGVwAMt3fV
XtRI9JX+FqDlkCZOq6Mv0aDIxB0Npvv6GRiVs21sA4q+4dL8ZB72bmYHF0nw
Uf3oxJWY7DjV8/6NqgW/nsAtC0ILJ8UouorH+DnuLAhoWQROKVQP31RZJIrH
Rh4OLM0z3qYaF8CeODtdD4ExKFBkm5sflb50ynTYHAjwEOHjOuaXKqNKkvha
z9GJiYyufckW3OgZIXm7IoSe2GoS+k4AuYtCK3ir6iWY0ARWbNpPDyIP0NLw
Wtg/X/+7UY7+1EIb96ikS9P8Kx4wWYlvy5pKvv6FLeoT+GZ1PE1KdSfvnzZn
Vp/VOKnlAtdROXp3lCU9MD+hnL6Irtf/XH5ddy6wegbHMw1EF+uvpdf5pkBX
+pR9oqY8MefJYfCpdjgnwL18dyzFwxEEVVBzPGCsqM83UTdBQAhrXftyr9rA
Rzcr9rUZBmLfwsQHHXqR0ZGUH+zIyrbMrwKW0mHsephWvs+ufhrAFfKjPV/C
C5Wd/tAFMeWnTIdvhNtpWwyyynmI6nz5ygYXLJXCtv6Ga4VsJZKwZtT3PESI
PGxs3Xmfw/u0eU0gODXGsyWNtIO6HHA/2dmwhm9UZCllOWLmgQrn3irlMIwY
b1FrWcuIUAkWoo5i2a1ad81JMNNy+mq7KrZkaHXk48G/w3LtwJLlsbsws6l+
Vrn66IiVS+HfLvHqaaMnomuJTTK7L77ShVOulnfXbSXv12S/DsST5d16Btdd
+dSuRIdLZzghaGa2u6jbLyXw7kQ6bXbWzaAIOjyOh6zy5CK/yPk+6Zp/2FbD
V8lCcoFlvOmDzaqzvGWBW/oaX+J+gV/Seg1wylSbijD6qVmBqVpLb1/vzwwI
/52c67IWJMse0G+4Mwl/PwIC4NeQkCCA/PGc8xH9iZpJcF9163JOwIq0SJi5
bGanDzaMdU5SjOA5hfRBdx5V06ncth6Eg/jUn62xol8PQ2cVh22fqemj8C0N
SOETj3bLHE+m401fjoZkerKkd3BxF2HKBjogAZ1KTbc2Ig/Chbjeowpmq9ke
h60de+of14RBHzL5Rw+jkUxRuTR0Y+ky8dKiUogXIXwr/np4xlNtOpj7dwxP
zfs13hGeGHDZUYory6CaHGVH/HMpDbxRXor6I+M90rjEhtGE1ZizduqcMRBa
hDxYwh4Im9Ms2a7wp3KJ2tf0XqfifU7OalNcDbyWe4V2bQUIITZ565OWBH5J
PbPrzvXAZRHytk9+u6P8oF8gYTBCwwCWpFxKnbudkJWP5WYTfSC8HBY3yZb+
FAiqVQuqkOxmZx/D5nf+Cg4aHC0+xo1jQ802SpD/nEWV0+PHFYWOGzL9Af0v
Kz8DqzcnxGkujEuvrtTfi5MxxDhLDzgzbnUOYPw51HAAw/oF2OHOBq3bs0s4
kltl8ut7k+3bIGNY+LJrkwjrCSPCt6SthL4LvzorXUDAqVW5dQ0G7j+V0R6W
1BEkYHdkMH/5F2dE/NQt2v1zSXi51F/7cOVTZFd/3tZwiDpOUTMt/Kn43Vbl
VsDFJUvKKF2y95ZULcdMMRx3FpRjCba2yMhDA5CtgSgsYXk70Skfr4Dfzh3z
m8YDYewP1th4CThVFQTaJNidnzi76DI4po35AxKwUfbb97HHFKcUcKJn46IE
+WEgq13iRD9TH85U89+w+nFz8ZyuENWtfc/Rfz+bx36LMOM0ppH/XpdhhL5e
oR531HmkOOyuR14pzK9OYTjnB7c2uausRLfodYV3B6WTkTpmqzNTtkgtNjsc
UD1wqHWJ+kdeKF1aRUKzu59X6tzixuXsdOuw+a2Pg5c2I5DkjZeDDbWxV4xc
uR6qs7iOD1YilQnfLOnL0ALFvehrieiP5P6EFAu6arOmoLiZ0PIoUlvoLHIV
4OV1lcI3E794Xh+AuGW48Hzf7OFbcLiXubujlLwNw6X2Voj1Pbvjd09RFQlP
4ETQ7Nhd5p9Lci++Yy/hNTa5dNpVWcbNkLciDRk831qIViixY6ZUphLtSEqd
KcHCzSRqoiFvAWifoa+KKyVpcxUP/HPFNCVHa5cU76UA2xIo/Oxk7L6m9T/0
DTcQ4zoYCXsXeDmqUEuPn97AP02IFjAobWuJekmSFBe7+zjzPvM9ved2eo+b
TcfR4t0V4UgBdNHOWMbnmKAwZv2qyO0Y5azy4Yy+MGNfojpkyNz5YByvw1cc
JVcIJgO5bYbio+arfyZHcdAmlJwTZkjG9mHw1EgLqc8/mPtWfk5KNc8NBSva
Sn8APIpLw3QDAVN7TMt8pBnbKJd5WSGBLl6cxc2iY9PjbP5VyyvTBhcYTWDD
Ng0jE0cSEeviVuHCwVl6nTTo8CB5oAmvveBGjnS9D33o9fRuw1C5o0JaqmRm
pSQQvyTgEn6rPF5WU9oppsIc64tKKnodTARkfIMuAxMZ8CR9vfKZmkY/nsVR
YVOGzJsLBadXwOOmb2IgoicMy9HCaPlR5zGwEivjxL87BNBSO56cGHY/xQzO
gxbdmwKyunvD9WZ3w4POYy225hcV7BBGDFaKP49VWWhRi1Al24cCtckaair7
qwXnqGmbG4muKW3j1eGORdt0OVqrvfjc3Ky45IE7RjUm/akvzPn+FwK6lMpt
JABKagkcCUnMHVP+OGCOpdzgZ/QeC6pwA/g9rJ7+y3TVol8XVCikNayy6ECu
9QJttU/yIrwKyassmhfMYekOkXcoZgocgYlAz4dhsav10pX3idH49sKFw5y5
U1SQsMcavYt17jRZyw/73C9bo+/iChy78cCddMIn0nVhZrAYkqIUZddQmZu4
SzaP/n2e1BcbEiVcpsN7P3vIQ2s5XqBsBxdJhHK+DXG1nJDA4P56og/6xG5M
BYBM3lUlqJ8ygMOooNYDPzieI/zs2vbArq6MoS09rQNJgjyMNjyhQpfY/oBk
z0dK3YkcRWrbACn/rAMSTYlqI/D4mCYLDmmHNeDgcp6WCxaDMT90C2GFF5hj
Zwj7hsQYlesvkj3hAWDbAMwbfA2i6COYd+8EJZKEU+qn9DSNg9A83TX9JHAB
m7VPlz6x8pyFrFAoFcZPb6eqr3hl39z38qljC91n0dV03ANTYh1g9uHUzreT
HFCCMoNQPYwrXsOgY8Up62hqzo4BPs10hbz8WYc7EH5Cx32yDa1IaX3/C+qU
YyiCJJs8J85WIZfJ2nmmwy5czgO0NwuyPTTv7x9pQsu9xzPo8ZOLXoVxah6U
UqbSwKDV3fAZZMlmwbLAqy3NYUuAwVrg2DjAIASIYbk6AfxTCOo7Oiie/y2r
K5VH99Y7ofxiP1C1nMUzJnob7WT5cttpv8lUJ8HyniN7Yxh0gI0n+BHnKpgz
paRPJB8gbakiS+grUbZm2p76BNzr/EjSmEXPFBgrZFown+hZb8dxJx10Xoun
U6SHT88YgO5z/iDxGYMUzTMR4zfxoQTl5+0yb9T9Qr+3FLwcfRNr7JxYr1Kt
SewOuOT3HQu7a+AMPW+Py2pcIj5eYeUVJx0tdJ0bYcLFe+is9Vf0ipGrY719
v8xftKwenTHhnQpgg6ekdAFpHiMvrHWTaT2nna2Tp5IhCmwgLEFyrcnimQZb
a1w4UmI2tiT/fFUCYPF2G0U1bYV2A7OOzs1qYNtnGcXMSCRJ+XQGjYcIzm9m
3fjCHsTSwgpp9D9rcQNbRW8tnN0X2IZ5Qt37KoIo40+XVcxSNlBJMX4Aou26
LTUWx5Tne0Y8Mvhvhps2NViGTrYx+oCiIxyH4ZrimLEx1Tptmv3qK3RWzPDC
AL/BD2mGvJq82uqkW5sDTPl1VI1XnFW41n0mlWwD6H5RBaz1Ii472udvsHOm
xEfMUiwc6ykWbqyTXaHB4jpjmbflhufjPHu8fNXFWZAd67YpYqV9NQ1fI4kY
HqyCWE5aa4eDGtcj8jaC7PS8aha9Pa8XEEu6SXJcu3Qid+uqI1VuQrjGv3zA
4qiTmjd0dNfS+9o/i7czaU2/bne59Bjn5hLucvQKFz8A+yZ88X3lBPiiDB75
W3QHuzwC/xS5ZzuagMm5jiWrOJt6Q1aVkpfDgdK8aa5wFBkCPl284Z9XfV+x
LuqJ3HAUk0KCvSiNsWMw0OP5YgsA9JGleXmCgtowYg9fHg7E/60VqBPghU/B
YVfbQX/P7KVjTcOJV40Jrh/1UFpuBoVBMuXNOwCl0emlc6Z5EJ++RyZSCgKP
5Xm4+mOp1f7vr1C8GJXbvDgtwUrCSzr4nF7RbWPgzycI7VqFy6xUp8KOnOOd
07UetKOgseieIyxagUCw1s2pKn/oBT72oP48LtFBwWJb+alCpcOVHdaRshaz
XyvhfgwL03iHoaaT3lJwxqSt6Eqo8ydwEeMo7QKr3n9SkweLZ1YdjRCf3vEH
hn2CQL9Z4ZS4Fn76wTXZDp/jJQZiKVh/BCOewJB2vFYaLNFiTcUEG+vGFUCE
O6wFDe7s4EsSmJV6EvB4R3iCCIZwNi6GAwE8Y3cpdFtMcx3VeuBYdV4AnAJC
ajEwvJ1b4Lgi8as/ja1dvDxxYp/Y/aHxJbnIYEadymy/milDLMkitz277gGI
NHWyY5Gbb0xiDxpcE3QbNU0GEfj14H2c8Jd60fdo+Khh43L/HoUFGwYe77/m
72bwLhelaipSZu0oHzt4Se955tKXeMjYYB5ZvlyaFhLD8Ip52C90Oa+eiE6I
Jzb1d8DF10Be3JpT6S641ORRAs8JBUqwnvAuKH8lDnwRXwgWrwMLVbbispOu
h5w6PAtWpthwDts1g/GbWIiBAoelQDoR26DZ5WhveVl3hZvCFVNqPw4esQjp
GQzXk6RoZTkHY9Kj7FBXM5wx4gzZflAvxk12fxvr8k6wIssVCVD+PiyO9W9x
C66Y32nXXqZGld2o+LT6r3bwjuRiaOpnqQSuM1bu7hI3BBsiXf4mWbl1Et+x
efz92m3Bf9Nk5EwsHtZlUvsIibRfYU+8iDQQX/S7v4yPouCiaIKfO7gK/4FP
KIIqj0fgXIJaGe2VJ4Edve2i3Jw1TPL/HdCvkgP5e2VVgJdVkdg7yBc6r+ch
G2cr1s0e0nmyzdQVDZ1AnntViBj7TvWHUV9oNrLwqJNw+Zucl0OCSla/+/xB
o7omVVQLxMcCKYI0Tchjm7zS67FBtR7KEbqBJ01guiXzUEe5Ur+Qzw7svXkB
V4Itn5ig4n5D2utX5+NCU4ptEjrUexTFrpEEjS4LupuHi6LHEL0yNuxZzv2z
25W/ZjBZoXjbH1FWYKXkbembR1yVhrNC4Ic/lclkAiES/XPi60qJSGb39qAQ
hDO2cc3fCyK4rwvI+C/c8owFISMiZcSiXARUqX9SzMczUVXeMkDwyTvMcRo0
FpaCdoDhnGhyc+ue1M0yf3GaQs6yCmF9buaDkgwlVKdOwI2YBbzuQPSMLzgx
OtcJgLYLAyDuquwSDa7oU8TKArwIiOQtCJtSQ+/xUJTnohO6F2Q0iTBnkkGn
z+3vaDm4ZEqd5IGvl0GmosV26g+Z64pYvx73661cnALTZwQTCzqDH8IiZoFd
0VFNXRTFB9D2ZFatlqmBXiR6mxJdQaOmQUULtHVoaOY9Ir+yoaBDfXFe15I5
AdEIJdAKg3RXIi9uLy11DvFq2LRiCbBrGlMPZfcrpmo4isIMcLuNoqBJU2cB
VyaaiLPMlqngfUFLqP+6tEP2ZrjevN13tUOaVds4+j9xWuD8f8nZwp21QTHm
bGrBiyoCcRSY62BnSjX4VC0oPrO5CaENQxU84BcMXKygRnVcX4XLRRoYd84y
uynnYXVVSiVzjpZc7x7YsAtoNb6GA3o9ODRjatVOdEK+lBbHSo7cf8hixdG8
o8yVI7SQgtwF6RvsuVIPVtJmUoUx9D8gi9nT5ke89hmqvk5E3ui228Q17L41
qH7mQHt5ZDubBTCnWZzAYGrtng2/624thirZixeBvNOg2RT2udoUaydYX9GL
UBwWI+PaXkLI9zQHaemzXp3a2QplRrlb15EWx769czHQzRU2+99jfKuTJJGG
4qvyRZQ2r1MDpZ/mQQsacriGrMJF2KVlH9qKeRUBcaTc27MvG96hyW/HTTVc
C2TUjs6tt17A1cGQzeZ6SMBQ6lUj8GHDwW0N1xBRsBeMAxu7FoXI5gkiQ5ep
qM65ZBN87oQyQxMRoAiIdBcj18Q2zMmtLyy9odOD+rgr7Go+H8U13oRGCakV
GYBFCBU87oD0iNM5qlPo7ZQBvhvh3cdP73gepc3k0hOXyq5B4+FbDXcakjTx
QpIJvEsRrcSizx7Wpw6+N4aYsxUjCGf5UR4zzeao4eY9kaequKc6ExNpTIgl
AddGvjrj15hBYZcKRFtJj5tOldzLV29S2fg+iSnVMQlyLSxej7lq9yeogaM4
DqFPlUka6GznPOvJJpGU61RG/KTnwWQ221YorU+Y/tPKEkY4ubZBQ50aC1ca
HcBT2vcUBkuDzdxhcH59XWi1rFZiGG0+eHqVwUmAfLYB2EIqRcJKetjRI0If
fUBGWTRmUlRUDOMvPBfo3WpvJRL5QDB88RkOyXRO1GzuXU3I2oyaTjSK6J1m
27Jcl60w1VFnxNpF56vWSTjrRn4UkJUa3TI8JNJQyiu5cb06DvgRzsrSRMs2
opmqU5jxpYV7jztFE4s8NTyUr+df/QyKZywv6s9ko+d2iWeol0rwW/2rSHIa
+wyyrBln/hwi2wR9VX1zX7bC4Scb4vKkY2JVRbRsdGO6nvRDognk2Ykxjgl2
i4QkRWv+DHUyvxt5Qo/uqzk22Pjp8bWEjQJr0MVEvT/x8UWFv1lbC59KVOGo
n4I0drT1upLQN9zbQ8CHAhfWQdgC9ia41e6wTKm5EoQEiZceunNpR0zGKw1c
L6bzWSTCGtBYnVSImr8659GxOwY6pvm4gjShcdhOvL+CKgYpZcWHPB/FVHG6
vpzFNra1ptYZC9ApViwJBnbgoyty2wr1ePbXW0tx9xTYGbm530Ra1z8PDDiE
0TK2kL09WYvaiejweGWY2u48h5yuYJolNqJoAjM70uvn0dEe5gu2vYty1Vdz
fjATgMmeSalA/AeEW2Rho7Lg3+5TuSo0IPhAijDUETugRmnI3mRadDVUuLAO
rJXhMdGnB39wEQftFiftFT3kw78kcLz929vqmcPWyLN/PtT/O4ZzITBWyTgr
r2vbdzxY7MI5J7NguIogyqGOIFLFvluJz+dcOzuDE0ZSz1hQyA61Jd5dYxQC
16LDXWsCwJRsDDg8ckSS39c8LUsRWmQKoNdMHrqPYx/s/2QbF+J4iF3ldUVm
zRmZuIsCjnM3jpvxAOd/i6bl7CeAQ7mmyenT/G2S9O/zTGeSc8l6d3r0dYWv
Fyo7kbgEDQv3NKQpEF24uhzqVendZ29cVr7oR1bng65/ifgvB214hkTKMpWm
+onMIs57o2SteLXRNxijUlyjmvqNvt++xAo4XwqcmzI3phCwIvHNQJ1vWxgq
uwUdW+uxFw6Tdla4KvGJKsdVcWDKHNDkVdQOmF2BM8BsW+O/2hoQoUjnPrDf
tobilRIjDi0HcxbAd4K9BuUmbH1SILz1THarQvHj1Q4PNMqTi9HCI71pg/TO
f0hprqfUpe5iiN7oJ5coC7CIcGTjB8l8eaDqA9VVfx858hoTvqlZlyPDhzIh
UG3nBe0gArBY8P/a9MVhZayRgB3P4lHLc9BmESmxFIzv63IA4U9b2wCg9zqy
skAtBN9QZP/q113nD4I8+Xyt3PNPiNkGvWpeQwQXJho9V3gGP8bqvit0qTKG
k76ykCN2t5OBk1xApQ0OFSGHtB163ul/ErrOV4KmK1xWxk4ZUBUrliO9/61s
525G+LDHriaDULq4YLx6Q0HvR6yXrBjvULIDf01n//k52E/ESd2QGfe59+yM
RFBcVZ+UhGS2nAs9pocsVvStgNpQwPHQRCymaJelhECDY8ZGnfe1oEC5Q3ZO
/ly8C8fKpAoCsn9oDcHQloQZ5m88vdUSXGOh8RSX8Np0NFcE8KMFymvzJ0oN
sPx9ZrhB4VaJ/VyAXshEwEXXk6xcmF0ksUKCOpf3F0gEEZs+aKQmDxebtcER
mrnUXFwacgOTU1u0mlJvNVlMcJdyo6eA/SASrf744OP9vJlmIdbLGgaEa+Wq
/6GzmabQF5II/OeBXJJjVRZN91wPHtVkS87W7NZ87WmIKxmOkdFJZR/mAi4B
tRU+tmLGMu9C0n9f10Ns5dJoQ7ZwHneucISMotQ4Zs81IjsbuxseVYXr9iTC
gcbEWLIHSyd0+VNqYEQjkleg+KoPFz+cO82FkUq9/EFFEi1C4rXSaefOp+fd
jUvkGj/S1q6nR7/OcrN3IO+B/jrLbZ9LGbpjt2kLz3z9GUPUh75LU7qsfXAK
gcqwUmMx4xdWIrpJSY9bHLz+ha0P0CJ69u4jnprsVcWLNNXycEO1/UxyIBbv
YWtH36fs0EzjO8CQSkR+mVqxGWp7wsGuBhJJ5CZmeW0DSOV0qQmXy8IYWoDT
mS9dHV+pwipjKosoIHi9i2yNUseuDAbW2oKo4i7eBCVQQh5dn+IJFMFMIRky
aN4P5W6RVy/iw03onUqFAZMUsmX52dCnZtnsPP7hrK7QwzaVtpYDkPAbjVfm
Dy2N76M1wE2z3o5VDy0KfBAoNPj2dJoaShQc6gxwi/eRPZZiiAZiEcrdV46i
mVxpX5LUII4FCkHl+0EoLmP0h6SIg9EADXCNJok9nKo2rwSzZh8k1jCoeZnZ
goaTK4A5QLjQAiLBXYmwgESDRwEjzT+GI9v8yZyJnxab6J3nlExyJAb3O9jp
92zEZIZt/oOcbQvriFilaFHQMaqQJeFJOcoGZD0pxolNRwK5kQI4YlPAD3cf
YSVh5OdPczluWWNVM7UHLI1lbTdUY3yaP40oUM8XdF6b/ZEKGnPnIJnaneWm
GYMcxAIVTJzF55SBMCc6zrctznAq5s5UcDkLB2i7o3BFwQ2RM2JdZbTZhv5V
aAtFldtURoUIMhDtR0hVybGXQcyp2ntrkQRQZGpi6uOjfv5ygFJ/xyg8R1Hv
ZDIKjVkfk9fxWrIanVMQKb9Fs1yWRc9ksoM4/uqPZ8kz7NawbJ+rk520jkPw
zzNYrhJaczbOuHeC2wnwiNnvEtO42u2Z1XM5mVwiGhmkQY77JZNRgzU3Ugmj
ZVh+cfM8DqC5R9W3h09bUUejWA4UA5QnTbTAPOW1dzualGUkqqqCTDp/NB17
jUAlnOgJEWs+8E//FdhxKu1dN6zGnp41dGuG/O0Z82Z7628fOmGMm8ItHgUl
Loo+04rZM6sFZlClCbZPwsJYtXQ3OuMDZ/wXNqPkiJ3JUlkE1kNgg2IJpKdM
uH1AUX3FcJI+baeT2jeUid39suylMLGLifpNbOiBj3d1LN3jUyjsPRKw3j7p
0QaHHOnasyekEqa4Yo/Ke726DjmN4KGLB7jYr3XqKjkiW9/7ziIDcEzDyIyj
i/zR96gKaM6Aiv1Z3mcLzAXPD2GRfpwS7E8eiFFrMGVccH0Xvs3V2TRQXPk9
8b5M/fJwCzxcCuHshOSx/xruwf4U4E4LushZH0InAQEOxhJtJkb7Uu9NqrFY
7i2u9CK+BenOafA4YJ11N9xHhm6KP1E1ojb5+d2tn5X9R9Ike5SapUDO1vQ9
iGnGBlHXhFE4JBWhXsovdRxqc5ZR+II44jC2EWVd96BxvBpm0nztYRlc0NWw
OAXAFF93tBVF9GL7oP1IBcVZVwOZdVh9U81tZ3Hc164Qj99Vrd0NQBMHTw43
gylB7Ix099Rcf4A+F5RrQUnR7po61tRINcSI7PLn92nVsEaygF0BqLngv7Rb
nLPuJnPLo5gdRB/+uQAx+pI5SKbW9KXVVuRvMGXPx+wyFMfgH7nI5iyo7qn7
KJRzPEYHkd4Aql1BtgZVt1hkCYfEvkaKm3S11sfnrENW0Ded2nfKhPy0kCkm
3LO37ZNnAy1abMXwdcIAKt1rsUhJaZUMYkqNaLG+hjatezkJC2jq0mIfhm5H
N26gtBsz8w0choGUIWLRDf/bSY8Gg2o3Hq8UmWxDFv4jSWj7gY4cWnNxpT5F
tJEP89gBpnga44MAViB8eCcZsf6cIftckeOiSgfVPJLSDV6OiEsP7Yp+i3gV
uTXU+Wo5lkvRUDaRcGggMEk0MWZtrCLzTduATXuvZvUMPmt1kva9zA/mI0YQ
x3m2uGM9s9paJIlu+KXRVJTVMpVLcyemno4YY2LAy4qxVsn8aPSbc+jf70E8
KyBnopdRbqYnrShHFE3rhPcMDICMORlNvj3iUzwkybIZZM0JtR54LHTY7fo7
lm/ozUavonjZG5Yd88moe8YjFIE89wRD86qi3ihwmmVtFZu/2ez5KhIQDPg7
X8rIengz6FIeArTgoDfVR2hUBRrnZcT4asupx3pv79rtfm8e/CUz5Oqxeqoo
JrOR22fUQwRIa+S8yphSaDgfa2jgkcTaxoAZeR5DFtLSII71nScxi2k24el5
4rzfQB88fjvgPtozC6d+1YqmqIETPT5zLV0pooDEFsdTmfjak16NYICi5mfT
2vzxFdgAZcpheq7+pbCmocYsuPO+1FZc8BrgYbNbE+mh6E5J1e+8jkLtr6GD
DudgDkJ7CyGsgnS6v36fmrroTnNk8nI0cqo5NAS1OC3WL1Hho79AW/Y15rqz
HKpXgAORS+f15rf7OJZsegqwTbmkhcZEp/ubu7QTreWtEKyED3C1t6Zv/p5F
ZIWhCeA4BCDYYLvUXOy992AxuqPnq2Qvo5t69BFLuvwVyb49fPvarvjPBO1B
M247l/YZ+2NU7nbiFmcUrs7TCicV+uup3l3wUY1ELnJ9DndPNrbEegYoP87r
E8NEBWi+ephHfP8+EWGMleieDLqLBRrYuKxHN9lOn5PAK3HZn/GyOCl/3A2h
arvBJk3nT8gcg1TumW3hNXNX3SapRtt7k3V3i5hu4nzj3QYOTuEkB5KPSVs5
zj/IXQJZCjSYLTpado1X3b1F1jHiQAyiJRzPWftH0AfT2mTVeBakKpwT3TcA
af095mNjWLEwAL5glARjxHd6GRU+aZiKD5wAimfIAs2R6s09LGoX7zGmxXrZ
ztSSgPnCd2tm1SZmQUE1WPYZjGVgLROPVi3nxKvpa8oHbAgQMrlhrxpLIBtq
aIafVgwfXvRXplV8G1B9DZTypUg3yKv8zO9LmBpQc2BK5YIiyvbsUFw3EOcK
NXHRbAhkkHVaOOSmqd/O+4GQ+42i18936UFnrbnhldc8i9S1ozLACZAM+kHw
IZqvSVhe9wYsaMMMdy46PATuDONA3VNvmXDFfEoOy3tPeIE11BI69ZkbpOF/
gx2zXqEnZH1l4qriB3q0Wlyd32s0jUJapi5dpYU8mu56TRksbm8cx/+amNqZ
ooz37cr8fVJMaYIBWP1oDsUwpespHoOFpR8+g6CluVSYLF1K/R+BxjhKVndx
QaieW/q9FvBxozVgL2JX0iovQZo3HoTWMJtBGUQyxnY2D8RJIk8ZipfkeF+y
QKXJfszIdMhial+6vBxPNrKOQl8NYetnvCraaFu6x9kZXz+9+a+qkuqdkblA
MEz41LgKULVNS2SvOTCUpIEzT/9YG0n/xSpeKe3RCJxc76R0f/hAmCvr5Ud7
346O9YZm/1OtLvZniRX3uT3oDJ4klkryOrax4F1cC2JJ6dzBmZu28G/wfioG
Ms5c3uqnbqSTHZQkOQ+g7LlLRMC54T6NZKGUFveF3B7/pv+WOJtqwT7/8foZ
DXTtNBSUyN5ZDbEKX1Gz5X0MUxvrY2Bpa85t6u3J0yL76dhb4h1dO1mkSCSD
evLic1KFHTFT1TPSuGbnhZaSVy/jZ1k3MqcIcwLEACaD+yF4ANu6UlujRAnl
hr+wgGpVsYd3kASHl+JTmEY7DdFD9EYgUq/CEavJhr8f5fAXE/uhFtGShTfL
ujQar+GZTlyDFDo67LuCWPWCgrO9BRAr3oYmm+6B2TQHPX2jLlFD4gFgDz28
cfS1597EGVOoXqzjFRlAojmOsX1Z8bE0sDMXppgljnP2rr5pjaDarQpoARmv
0sbIv/1Sl9tMrBLhSIOpXxcJj+nl0PYwyWQ4z/zA4ZvFO9sLcdNpWHiWZ88d
2dajngpnFY/4tzn1oHtsEBzMbbIK1EoYsmjQVg6JtrNPaHMoKqksBPfdfXqZ
EwMFAMpyFnX+cTyOePd3f2+cIWhC6mejB89XQKj9i5nw0hs5m/C+27+3c4yv
s9akjTqsgTHca8EG/En4XMPkBLUo58RdtiD2OF2/p4wrUdlM6XY2kf34kq5X
cjdkbaUn7bDioSdEtaenmbfqZsrzDA09lw3LYzIRVmDKd9khWlJ8BkI6pHyI
u7/9lY/XIvxF+ERS/JuKmERw5i/FjZ6X1HrCf2rPQgdfUDakIgf7+xuc+/L1
tdRgkfslnSa9no7tVOR5VQXrwUKkcvbA4/Oiu4S4LPXdPipJ7J+UdPnq/G13
SST1Yv5kCp5P6IlYatgnjst5D8w9aBsf/rnQ3CpGITeca2zqfGzTICtgJ8hY
AmUh6iPjnW/VwvqHDKcgHW8FAACuu3wjJhceg8gJ3wYfXZEktGC8Y1iPnDth
RGJbOcgsidUyY11bohSjhLDMzuV/dlXE5PBxryJH3/2quk8ZSezS9HNooDRc
njfC/JgNz2DNW/hpXNM5WHejifFWIAts7FbewROjf+3rL6odchbq8Fo90sJu
bjcjFP+w/P9wz2rxfgGN+Z1/t8qhWUe5vgWugtzyAmcpRDr2JX66puZAQiZA
M2iorsWe2Q9tAlv38XjQXDY3odBk6D3KH3tbbTHE4AX9E5dwdMSlwNL88Pvr
XYO58Tm+/chEaE1rGgjv2wiaUrcjM2hMaYtg5vIX6Dv2PPjEepshtFr987Zi
rK9wsWMloQW32xLuqnlNEy+LvdXjhset0MLRg+b3ZyGBhQC5WtIAUPOqxsxB
1UjNplzvaky6y8YjFQ1Ewl58Wzc9X5nhAZSfQ5YSwH/Y65LfgDh4zM3CiIjy
YF6z2soG6EUCZKD2UcoEUGitQ5d+nb2EeKmOTjIsPY1lFt8+CRn+Ys+ZFt8l
aLpSg8GnbpRUsLkFfmLboezapWyBtGimuX5p2BjXmskAy1IqqhG2OUvdZ6Dn
0pUNRGNe9tg+jzOsM0xnaBaQcn5X+/ZD2CXMjepvgkPHeOJeaTQy0COAc6Bj
mXuz47J4A0RsPR/czwK/K+7J7wBVeZS2G2TBXWhvZDzTmETSCy9VnEu6BbZD
AFDu/cees7GiSkiIthkV+y4UjxMbCi2tliZmIN3NBIN7hkUyozqo7Dd1176K
m0QksEzJzHsAhlT/UWVHOUBGKh4QhgBNOOkTDa8nWXbglP2vDzMJvNsdQxb7
I2xvFJw15912bvuVEyBRVxh/l9RqGobwoiF/5PNVI561QKrZ9JSqZqv+h/q7
K90dWZ1TZJ76abzko8NUFrBmrOwFTKZg9PN+jxN8TcaPOc0QR+vMVhJ1zDLI
Dbo2cgHyPML1/GiTVi5sgF58afSFbUHecAwqi5NjIAHbtfiqu2v0z2qnX834
sQpjXlPuUQe8I/lrSyKBy5XFBHPWFN7PyhJW+x+7+CyMqE2ZQbdjTklOABN2
Tnvk6dbz5t5Oh1fFBK5vNqjR7Y6TrgT91eciqy4ZAZqpSO0izAy9EfqJevrh
EvAYVXImyYOAMLTadILxgQ4ffU5al+nYSGjhllsIM8FipCU5upCFHWOBvQsE
Hd7bDcg7JalznlBa0cN4qKzNaKA0cwYlv4KLd4adE9gdl0aGnRJLPWLvN1cN
kAXv70aCODY098Fk9z4Q5/x6GDu9epbyJUDKn6Yb9Ri98wdiqZvPDasv17rb
sDAq2VQ3VNQROyfxt/O/Gi4ma348yZzQcq19L9GqY6h0lBEqdKrXvokHkeKr
86ZTZ/GHdCdrXab4tXrUijOT1lvFhzA0C/zaQUGUheBd7v5O8CnPGCyerhID
TnFkVGCmF2daAp5SL4+wAQGaYboDmuwCWPmWh8/X0m5KaR3FCTJwyt5RWE6Q
4p1rmtrrkrLMD5gDj1/G9omJzzD/IWwu6VljrLvZsGnIKwkSV4wR3N6EnOcG
vMlX8nC3pR5pfYEcvjbDxjz80JRqjEoTkVQHeWBzuUKV3XHtPi/viLJRi2er
Siac7bHAIFZYAjj+xwFgl30jat5W2fFsY36Ri5OFxz9PxQzDBM9qoQ1wz4bk
d7f0issLTos3Uo/ok0kvUF/fIVLlqraHtwmzHU8v3kdeVLmcOoCk3xyiTdmD
t+rXkqPXPX7L7XD/6ALf71C9VldCIBA/jm95wt0AaSm7Y1mXc5ECD8rz+Ar4
uLBpAMpdXUOE5Ju31PSnWovoGU6TH3pzZ45Hcq1FTCtrdNvWSRIUOgvp52C1
F37Ax5P21FprGdH5ejElbhMhi6XvBTITD+3edpUZ2hO5sG0sIozFv7YxSqqZ
VnNMfOUPwGwuFyWuoVYFy8CBfQ2rjMcSP4Ux/68762N1U3AMnxYzA7lVT39U
O5PXPJOSai/E7VqYWbSN0GmEGlVP2HFc6vZDhDGK6qLRmexnM8yOyybtC+vj
4JNUw9GZzo6bVdnWbcwDuUJEiQ5a7iFlyRaw84jokVU9Kwm1sLi8Vtt5EXFq
mABN5XvZMJljTu4PIsgNar904zPwR32oMaJVCTvNSRd43t5yAZJaOZ/10Qao
RY4rNihIILCr3DgT0fPoDbxEqHtQASnrbp1QRkeZ5iUgkWdmxKuOqq7kzCKP
UULkbMX7E2TRmt4BjHwStG26TKZAaQ3N1lnvMOMXhJJEIL76Oo64bpbp6m+x
nGKx6i8HVxXRxzhm4m4Ctc8AdeSHRetVTTIYebfA0nz16JimeD1xU4coyAHg
x06uUkp2WJftzIj+SF0/DHKPVNCvpWBoWPdJgbvgWlPwFt+0V9XJxm9pUymm
ZKmnMuJ92k3Q9Zx4n3xo7hNRHvgV0dVycoz5UlBTTG8Au5Wmy/I7Mf3o1UsD
vmjBA+m1HLUv+cXaWTVbMB7fEaXF2kHNsX3sikyoAnZPPVlLUEpg/Qv8pAJr
9INj2nDjMhgnAoYD2Vo0kikLSbOOC223Eb24Ccw9iQTezICZux8Y+JvcclKZ
r+f7502IJPBTkVDC9s43RsPHyT4e+dEYbIQT9s52WPesXyokwK2FFys7uzX5
cDlpkBgiQRIedqre8GCHiHbljTjAfcFLTkZ8aa9twdN5GKFsviIfC168AZSr
1U+6ha2RmNyNVC6FXp3tHQqsJGYwnjqZu1mg75N45b72HKmxoWS6QKwRd7px
IwqhIqm2uQYiqpg6GKlUecCDe+SOCX/lyCR9OAteRKhKQu/3rUcMy+z36FE5
pTfyjGbXABD6/GYEMtsVKw9sZeg2pISxcCoxesxy78eYVlkkmOPmzShVfraa
gYwTBDN0+UrDQCV2MJVtMRuWuLtnn7s10Y/dScGtd2WOBMZUxAVYVAWLQvch
8rNY/OZej/ZGjGiQ9Fw+Z9p4RKxY6IGcR8ik+7nOeiPZS7G4jyeB1MCdWA3R
ET2PpnfrY/ByHRequNwpxfgH+vrbEyq10GDkZWLAME5jyL0FHcYLIy4NXGmK
B74jBeZXlUnEWKwVIiNOGTlh22s1NpV40Vk1ilzz9DRUrLOnd9wuqxgv6lt2
gNzrKMrFKRsnCxYpeDkm1dZMNvMp1ejTTioZ3O6F9N2++klpUz54LuMSCRqO
31HuZ04jkkopqG6y9VapwFNJg+61lnY06f/SQ8oHgtdj2jRPNguFnoVcqOIe
TOt7/LxymvcA2Mbwbqe3V1azTlLtiulln7kTAiq/ey7m/NVvc4gDSLn4sFGW
N0Xa7V6maqI5b/rsnSRzXdo3fc0VVlLfDuKT7Ua67uCtmuo03a7hQHBDk4f7
3kQALRm6DrAU6Q7N1YO9OGvLUpZTrPTIGrowcbaGQxXZhGTqEbb3l/TjrX3Q
6bkZ1o7RyHDwkxCrRPIYYHlF+3WZXPOEBejEopKZfjDuaAqwIwlUr4m/dNWC
2DIJr4zj5VFPAv8nseYP650zU2MeCKVq4QoO3sEXUjSGBxVNGi+9spSKxSoS
g6G7WEiiWwqBSC+2EE/kypK/HZT6HBelxaU5xFdweQKP/xDP1+1YYLAG13wi
g9PptNhR24A5+y59YlNPtFX8ebLfXa/tMiLLelcwItnJPNICoQBIl+KnwmIu
JTPzhkVoXBb40aWfIukja0tiVVehdFEA80eOyoSAzJmZkZbhN07Ch30xjJzU
fdjXEuU7IEN+APDbXLAUMPMHikktg2L1ypERwlg7tpt09FZffLSOw8nuYLK3
gJIqwotBhp8yVqD+c59zZk6+1p2dybmTpPBrreXt4se9ZHgDN9+R3i5S9+aB
lJCLm4dtunwLF0tPQFYT1plquzhXaDPnMthJkn7+T9vfK3QU7j/9hc8O8L0+
gWtUgXKEapl3xrc8FXXdCO6UMB6bFy276R9+2pLbRMNikpz2wIkHkD0iIq64
2STfNN6QVBafuMilkEV4k/USgtxO844MENIssgtJpAXx2+TnKhPYjyvGO8k3
mg7qZ7WJVPXl2bnYWJ+JWnEs865zU445T79NbWU1eiYC2QTXWB7hVDeKwtwq
umfjr5bZR62N027Tg/KPg5qoBP/LU/v1On0Ccy6NBkelcaf/s27hGNIwFhTk
FbRkHf8j0ohVu2/rrfDc2c67ts0MJ7ufCe+Nv2P2i+4F+SL5R3IqUuLIC7Du
n0E9+4YeUcYzwt7+mNHHEJb4lqTl2JmjfBkXTkGZD0OFwq08nxC+oEiemaEr
Imb+5me7yr5kwBgy2iZhrxkHCqsOzYWCfoofTL1tIK8YlgtRDMwLsuFjxtbI
S4eTTInbuZ72wFflSXc3qi9Tc8uiVbYaAdzbxoRjWVmhymr0CIMPKwXCiqFY
5iTXIiOXpR3EdZFRltrKBQRB2E2QBAYIsJNPYLqWK9hW9kew1savPK3zJ8vQ
P6olvmCLYAW/H3UXNhSQZY22H0mxqcyykUBDOIl+iePzcXHIMALVXhDeHlt3
DdaKN693hWxoXR2/MfIKQNgRmzSXYSEXrGs6Qej5PFckc9h7ECwR6xfk4fly
YHSMsIqSTS5VLMpNSrY1mHDvgXWQaJOhjz8mITWF7J0FM7NZSVkw2KA1Bgmw
3XEO12LDPMNwvtC4qW1UilxKa2a/sk50rhILL91Bg5sr1ReWXosOERYAFH9w
rjP/N5uErHhAasOSg+Z6C/Ov8g/GZlkmzx7qnyruSlO1YJEvla4ttqFNXhZ+
FgBrX1uNgiont3AurVm/JYr37BoVjTioJoUxZlNJEmbyiyePpnjW1LcjClB7
vuh6SfRhqJ52tai3xUiKoZ5iZNjFAeG9XgvT9mtXwT+4u9+WOxBZr7p/XT2Q
PILi8nKgH04Ff0l0lrjHWyr24OhkBG1uTGXuPnRhoDHG04T1e1l8nabJR4Ze
Z9MdSJ8FCd5U4LMB8EO9+mDJt6ln2YHTHMs1hkQjiVDOIWbmBqZ1zfK7eqGS
+BcRScRaT71iUBWFBuwfU3Qtt/1qiRmf6KeaS5cXyAATSwc204e5z01e87Nc
VL/tTEhKW+X08bid52SVynNuSz2Qz8lcayt4ZoBrAuL7NI9UWr12YOZCVPpI
xAPgYcJQQBGX150CxHFYMueJ/TaP06FccjSZJZfUqcBsUWqVIfCUCGEsP0vV
jP4LQNDYyZ7vlRr23K8abyDUB+F139dsDNbK3+7kV45SKi7gr43bxH2ok1Kn
pmg1W1K05PO63cfSa0d+crWYc1ErApV+nwA6jf1rsyyemy5gM19bWIq0pa4u
rsBOiv7b4bI1QI2ai6yLXyW8zJZIIB/1WrQFxGeT+8/W3qTkr5m2uTo00bvY
PXkPlLFod/6uB+RJQ4Ba5t0coGiAiT2Sx0eEJXQ87zw170oBvqXm4C9jmOvk
o9iJ7S2qJtyOPOv8J+9h/3Cc6jaUeD8RjvGiLn+bX5dp9HvJ+f6sfit+07Vp
6CnNCHQddbTiDtqddxq89Fg1MoZmldT7tORJFpInWXxwxZqx6sf8N3gJH1jE
ijtTikZeK4yJy07nzbCVQXGFxcSxkOZhfrqjyWc4g3ekSTJ6MXIgUrAX1Epx
3xBACDT+yiB/wxGbW+WF2Neo6huZSs1OhXjlegx6rjy1Q2xuZc05+8iHfzeU
mH1/9P+JY+J7gWLvhUyPruAfKJIKzPTGPNdW8UpAl9o0H0LRgkbc+4WpQI4l
YWkDSCc3mC2lS5CBOuKneYuXwesVG2lNlujLIGcMXYK/Qur2AGd9wAH/WZ55
t2qiqwIDjeBN7M3US4Tavf960l0jSchCYjYxU7Bb6ohhTZgbR2vMZNd26hEG
QGY6UmlOdnGIXZcNqbP8Qun/avMIfAKdT4i/8yKZVCj9oaBBeCIn8Cd9CETR
b+TYGOOTI/FTpUwX7x1El4FEexhVkP8VaGFvIYsAjcE69zeXy1UWta5es5v/
j83yNCGDxROiCahOET8pPyJFrKpvUv8oa8GCkn95JQWOBuNkIKSprYYc7AMX
AttjchbdGdorCDhuansv8/EU/tpgLmV1XAZ0BAdeh5sw2FCBgTINXvFV4Bet
k6u9GcpRsGfnHWRNS62x7HPkMW2ul8VHOfWAINn1qQvCLiR2zN/wo0/XGbOg
Rg2G8DWQhm2dU/67BGjonG0MhFImDvl1D4ghS/jFxdqBLDZJgLSt4Xtiy9cf
9YJtkE0mOz5k4bXQU5TG7NXgNqTLYW2tXFQNx1JHotA0nxmtVcDIikcx4MMu
wZ9oMVUGVvDMGAPER3MFPhC6brj9iJZNAFPZiupaw0maCGj3Ts30gv7B9Tog
taPpsWvChtLTxn3YPovKy22Pts9zrgM9GFK/bDlTuavIm7Ft4PKQTPC4+qZx
E1q/nM/eEtk5Zu11j8CV0PIgoVxZnu8PYhlClKqsq+q+0Cp1OSAeAeABnkF4
ZTZ/ssWj4g8CmxVkTeoqa17KZpOjElGUfjbs1TYvQwFPfa70rggW+CtoOQLQ
X4WVo66vDHXm5oFf4UnsCr9fh4vz7Ft5B6zhC3tJ4MPMSmfpnogBEdby5TVC
uOwdPjKkSGWXQkumfE1sbXxiZNM8Lm4GcmYm8xlKZw6J+CFMD/CCfd+lrXRP
Gp4lJElTJ/cMXLVMQjE4qV3Vv3m/fdzmAzuenz2wwmGw5H0uHe73D8vk3sdZ
bwYW9OiTkRgs7R+oQBQ8CekmDWLKWBD9Tdt/T9nG35+0AfcrDqHYPym7/xW1
iieuNZXZChl5p4wYuSo2Mvy9ZV3mmloyN5JTTWNTusk55jvBLzjmsc9gug4+
5icacoiLe0gis1nCaX8RHFdfKZXqPjw8iJUF+bbDK/agCONCdGU6G64M8mPV
8dE+MlOtQ3xtaCdChPtA3eFkUYrMfa47RyWZZMHZ/Y2iWJDb1GAmbMBnu/oa
BYYC9ELKQdGvMy99meEKCW3CB0mLN7x66qJIAffYIddmftO5LYa2fx75zbnA
3/vZny6NGHFH6IYlapmv6mZpPMIg02i1PiVsXXJuyktQHfoK9Cb0m/dpOjoW
5jzQdntBaGggpko8dSGofpe7UeakHzGIqVLyLvzIUGc3XsSFsRnexgpJr/TY
JAa5g0E1yzFg9OJGl+yLXz3xg0V7LH12hGuAVNbEFQtTJ7kvLdijqv/9yMbE
Eewougtlc/InyC2MZ1EjlNrDYFFDYp94dYL1lDebVW7OtOx+Y2ixmvKvefwU
fpTW+3sXogVPq2ut52HSlfIKxAOhhp1K4e9i2SVYievvaPtxrk9FFz+m8Gru
R+YdttiCpJkSJ83FdmiZje6+MEhIPDOEkYGooy9EblRuasD077vnLt4SNrvr
WxhymstNp6tm6E/d8SnNanxVPN/7BlgufwRNyVAEFwnFP5HsxfDaavUV8Fdm
lnJBqbBHhayD2eDeEaMInNNde1CDa36YOBJMZvcG8oJqyqDIWWs+OEGeA2m7
naSdzNFA7fz4LQorCena2EMlqFTemJJX8BVkyNE9vlpML3lZANHce0F+Nlkd
aOlJS605j8Rn4qsZnEGm10KeZkRw4iBYGLpB4aWexjDFaskhlnOZV1gcrulr
YL+PykgKR8KztICpQzSvYIv3KqjFCHOOb87G2NXdqixfMOA/qWaHCa3CSuxm
bcCMemfZQz5aNqt8pzJqmjBwWw5phRObRy1wsousXQMQI7y4w/WcOubCEHqa
gjLAn7qMhumAxejIQxURYMuwTSxIwHsq0+c55MMET7PkTEIKFUMZvg38LQTu
vW5rKMG0iF7NemITtxvQDy6IBxuX/3L3MXeyz1x/IMTJIdTEKjmA6c88RJng
r49BgGc/lAHK2rfJJ+2FLDu5Vtw3A4uPcvyJKBJtBbIChw/WVK/y+2ehaP7c
BvqrsA6vaLKeKGy2xHjplC9pA0erV349S9bf1vT0TxL6iLPwyyu7C+UuoDcr
HQ4K9XXWtA5mFs5MmF+mNLSalCjFVrPGoQ9jTgRet5/z9SGDlQ592UFpki+R
35UctwH3jrC5IDq+Hltz6fThhg+zG5dvjciClL8DB7wUBm/37ZcIIQtB461u
VZ2d0LDWYBZ7EKbAxXK9gm5TBIOyD3VEVKSicND1/7QGzMMeurBP4D7AhScs
bvG1vybVoqlpBNnaZCh//PL/XA1qqNAhv+rNAs1DNIkPVul/DywFOqaURs7X
VEZ9+fBWYw37A/nP0dwQbMCFYcL7yqffaF/G5eY6D+q3i4zgtMdRhup4ulsT
9JRQaehSj5Ygrb9dFyFuBQMxQrHQRDzO9J35equAYmKbKnAwYDorYHPe0kLb
IcUYTPuNa1cX37Mk54jieshXgtRBaMjEabyQicplVC+wqlk6Z+UtY44XArGg
aRV7v0KYtSmM2NYTjFUUaZW9rbQOS0b43CCMN7Nr/JUm2CombZ2gC9V8efxE
KeSNsAuJKNNA9umG49To5xgVP/Iu6xuqNeB5uXJ0lPPh4RTnO+JKD5fo7Bih
njE7Z6yGnK2TIoKRtCwVAO0re+3Mr3I1tnW68JbotbIf7XjXZ6s1dz4PEYVm
8TXxXB3DT4WWEv+DBs9eNT4isPQkZe4DvkE0bkH+hAJWgonAUPmZNfdHHRJG
LHVBVSaYrtT+h6AggNw3tieZL3lWGawFDFF0zk3BmTsc+Q3R/e0119POZKM0
qn3rKBIsnS59nZ1oAtgi25QiEYaK44zyf4OpP1PSIfDM1/C0M00OalglwyK6
Kj3J1FEWHFya1c14lJcghusL2tBducNfrYRetAEyDNq9ypeHanue9o6Bff14
vUFUeRRJtVRp2D5pvnv2ATS+fp6KzlQSs6a6Hiic7MfHWId9SxQOBsY1Cc7A
MdAE4bF8MF0yEDJislzWRWzLjtazloQC0gUxWavsRZrD3hO2/eKeY+NUMfB2
Qi/B2yJsJOx9OVdS3K+bhhe+g3tYTzqyjhJQ5RP6U69ZASM69xkJy9DVodeJ
oRkacEg49mVn8EK9zBG4ssfVm1R2pKZ5oGf7QZtbuF2Hhy+yHdkb+KxTkiyG
tGlbXMgHyLUwfSCgeP7BLHTJEiy6r2ZIUUeJYtmPWHrjJBezSMHeeD0T4IaO
MRheAMuxxavyYqlKOkpRmK16yrN9XiOmHKkP9csD4YMvUZeth5Y0NiAoJ7At
AQrOc4Kfc0VxHzoC7gXsY26LsUG3xovCagbpPRWejsbbbcGff2RN7hHLIJM9
oGKM1RG6uGEBwR+8VM4ezDCVfAEjdTgUcmZDHE7g2N/9Fi/aYguYPCb5dBkE
QqRs3CDj7EwbBU/WzUmnEpZQFX9WG/d6oPGQLLP6XEIYYhwSVwLVIeSnVLpN
CahaBKHPCEzFupwIQqupAABpExbC3/Jd1z7w0RWm95QctP985WbsesHvplUq
TTBPn8BlBvGhmjKZs223xt7/RxY3bb8HuEGXFdeorXfvUwn+AKaxXV0/2hoS
PG7Wvgdk7Y5nvcmuZECPOaOv4H5a0OUqYSF/NSlAHhPbg3gNCfnQbEvWu3G9
cNjQSLPvMfTMHOJ38TvQtWXnEioZlkrbLqE9h9iBD7eqJ+rgXNtoTRDTI3mU
ppBshWo7Hr3Wz0PQXkinJ3qOs9pb7X++LaKDp8jNifNZB3XA8cqCPo/sI6NB
6UKUyv1bu2kfY/MPbApzrcbNC1zA2BIukaneRLeiLS35rQFUWbLDKVxnZz1X
Ad0W5vXFuyK9+o618s6vS1RWwcRANc/KIr4gK9vhvYK74ZNqD06RqeCtcpKF
hlzCE5wDLoMRws46kz+9kecy0GaX7gKaiwjeMWbpOdZ/VEvK7DE7SwQmSQ+u
H799n3UqiwCZUG/RvptpSVOPkoC/SyNzi1YA0YEE6pWfLThP7UQDBEq8rMQo
1NfruZpo3guUkXbzGcbwi0T66UxDlUw6/sbG38k/oMesj7xw5G0Y+MjfvG4Z
ZIfxFdaUGxdY1kAsZgKLUpQGByQ11ERdncViAiIbVolj9LrxRK9u+0RL++l9
1RRMyQVxksvRQdqGzXVbNkth0OTYPcYPhqpkymTR9yXhwEPQDxb/zcW1S32V
7YNekyTO1brMhwol5y0IBixpbZjKpwQQiBCw2JZInftthAoNbIM7cVo8PREi
p0u+g44UFlBdSrrZm1pfMh0klAkIXCmecLxijpGHrdxiz8j52nvWAI86ugCY
bOvwFyHli/AFGB6AQdy8zEOJ4FWjDwhOFUrOJ92zSynC73Mi6PdZX2X4KtSH
38OTxKVndKcee2Uv+yrzWcftxXXUv3kRj4DGlJgQ/2jZQ0Nx4h7MuDrAy1wp
Hejy6aD1Q33DGm7CsSEWVWiC8HCQMDwQoI45poRk2jKMYt/CrOl2sdcI7B/7
m1H7l9YW2uzxHGEIp/xkHX0Pv/Ts1VqajEJImIMGEuSg6KIc60eE1S0Cowp8
MT/Bo1Yv2dGM5sFI6wDfYmCPS/+dTxB5WdXDwSXlDpwhCci/rNIGzcrYM4HA
diz1VGK4YQK0vnpDL2wko8sBWMmIQ7RfGun/LhbZtDX9uzNmiF2AwKo+ihCH
MhsoywBByB2U9+PstMM9MFqYTv753gf/roSxmLB2v0mkl/Q6R/+AReCr6qEw
8sQbK9He+emitSesm49/SIi12okC/TwSjcf/4WedwFBloXIiClRpCT3e4uIF
0z2/jOT+IC1n5+DU0c5Y11zXM0E+Wx1hhvt1zyOfKD13Gap88iJmUVT9MDiY
q17v4ODeYDOAZmcKJb9fNtwPQR173LzUeBt8X9TFIVji4H18UOfnGUADebOI
HwvKqRQXOYMPXkBBCvtCxTDwqU+wSGZRXLa8WzG4nSaBmrg+8Osrw81x8c7h
gffzt7CusB+5zY5P9Vl2cySiRee1vojCezDmjIR7Y/Gr3Hne/wwXFIxD5fzb
7EyCoHJAAcerMX8VR+1VStpz6KeKkUxqJMuj2LqW9uJvgeUnllFzU7jgAFLk
nBRiUDyUajDK6k1zsz6LV1j8aSxTQaSg2RBmovzRhx5TdeAORNrp2RY7K1Rz
zxhbBpd85esVQAyyJtidoz0hBKjrZev+DLzZoGpxyYS1We7McbyvXW9TZ/V/
EGWFB5g8VRLdiFqeXHJPXeuvZj/+iONDqFnmFVM041/NPcrHnPTOGW/LTOAP
UBIozn8YVQaPufOUEuT/1lWOoKxUl05uhNfQB47A7ITCLvLFwYwmj88G+IfC
AJ4cnFsZrMmCMvihbi+vZXDtL0UUPOimtbYiXqlXVLHxIIo8qCRZotFGjypH
/2xNFkfZxhjEg0W5iy1k2plMOS0GR+YebVWuWjV76+t9oHhoy4OQC9b6ERmE
uT23kz0GQGBIib/WjYxqhxVV9vY8rw+BrD98cQREM41KUfrz1TcVuF6punlk
TFeawMqm3YEGLITmhANidsP/2A0MgqZ06iJ0EIZps4LIklUv79ETOd4vZ/Yi
76SP/g9fFSsRZfo0Hn5UoBgPkW+Z+wkBcA2MXcUYOGyPHowxprVCNZVEV27g
CgSqSUEk7q+nohulABSnao0ptzwD9cpAeW85y2pla9tmMaHSCxIK9zIM+lCX
AsmDbW5rNDC128kKwSu50o6A2lB9DJ27I3uVseGQ5GUSYTmsOOugyz+NV21F
gnOy1LNo8twuqnwSSJK6U87f/HGQuhFGyQVjp7qt5nJ2UiWp3WSVcIKkohH0
6StGb/jlMwTLJ9vj2nbgCwHNUxZE4OWPafictszHec/sjerTNSffwOfdelj7
BMdER+3V++En7jVlYqzC5Tl6rHCNzOACV57w25wF10kPAHQhsRpfCqckaUa9
kq4w5E7bwIcb3xjyYNph1hmNmVxWn8+hxbPlrePeg/fNJ6hMyg1cqZ40MQWy
Z8owzVZ7KaHDYjHMD8blSN/qWKkUnLSg9KXU7xyV0MfTZHxI8vWJOqqWjFcj
eeC23yycp8inBaRN1OeFjgNrORoVdjTC5B7RTkRcKFc9pslewycg30C8N43r
S9kjnZYkkNS+dCPtejosk8Wpp7melosBoxykd5pjvE3Z2ql7g2bchVY0Th6A
16Et6ZerWgLSfSoQhl/yF/fYrafjBEe/cv1rE42SU1JmWC7JMOX+QNaWNKc4
Xu541VYofoSb3IyyJmQ7wIOJ9cJCaKEqgh7x8UErJdqQfLtmlQstnc9C8qNi
2agvKC/XJ8UW7unhZIgsAT4SAXgcY4zU3V7MJ5EDAd3uVYwrXMGh+4CRA66A
8GxxdVhwzFYxOgwoxUAIr0y0lxjjKU0hTdZ+t0BXqHJmfhKbolOYfaq6ts7a
Du2Ek38P0cjEAXjTnSky4aHlpw/sIcnEBewinl4ehXpUKCYTWNSGGTJkFOn3
Lnhkw3XG8RwrnME6fNKTHFB/0CX/W44DYZJOGfnmX2uMvSjoFuuZj+zR7JTd
lLNc0/yPI89THrQ4wZDnKKfmVOu1+k9X8Ac+mrClDU6H44IM5T+rnJ+fDPWO
baZq+YYHSwYf+qdeAY+mFuyR5TorYIek2W9Gm0NbKG052sLKFnWbqLru+2Gg
FqLk8uWkaL0utLLy1EwNPZGEFLpaLAnRacNTkd3gjOuE48NVwezma8ZUbsfV
bClHuJqs0evm8TorQwojJuZxX2Gam3YiBbv4HtTGeiGc1hCYHO2QeR8lsKo1
Rjzz+S+vznvIWxKeX96/dvKEXbeGxBKAXfbB9EXtC/2CwGhGEh2oV4IEznBd
9jrQ0O6+1nM5NfN3lri1Gkzxantq75lihJ4p9MlKZgBXsaZxkTqm8zyWiP0m
K8VBISoc/BLGq1+DybD0lz/bS3amhoQoJuwHSs4TMr8JjV66x14Fo2jCp60+
6rMIphMHtdqMACZERUZNFnG7vufIQ7n5RP/LQioLaemYxp3D2lDFmkfm7X8T
3sWOt7+fYI8Vt6Aoq3T9EYKHBlpSKJGp38sqt1VOIFtPvkj0aJ8Aqfm8gsnq
X2nmF6xNSFfw4N0g5sXgtowGGV+h9FTsg9vsEgfD1NRrD6FKy+2Vbn8V9x8g
OyLOYm0KmEMdjjJ+0r3sZQHIiH/yVdM74D3zrF0X7+ZY2eM463sx4ry8bXmR
uyTL1ZXf/iq7ylfN14ESDB0mJLMWzR9JE6j5cfVLbHWqvktYeWGvrYA5XIMM
BSFmjlmBFyiNbtBOH6IBOarSGeUkFdFPbDwcKmhgEBQ4GZaA7uLbrzagu2BR
Fm1Afer6UJ44hBOI9T+jvENg93qzxFVtgmIXJdmb3P7KrW+wbRaufzngGp9s
RjKYvY9B4sM/UQ9O6X0FejOqsxWN7bVQkssES/2IlXlvso5BPWb12MLu2ZT7
X5Apkq8HzoYjYBQvHx6p3RwONeyOAp3wctnybhH7vLzMRZt26dRVtE7L/2By
kRAQ3fju4TWtL/gDJaD6Q5pc7NZp1ctCOZd+jxkGUo6UruI/fz6gBP1MwJxL
x6lfULKe6gzfnpJM7pnjuwZHPMyVkNh2L4nf3Pa+psfnvaKXfbfR86bUGCIY
I+y4/O4jpzV8TZ9nsVQUitNEA0hgnTfeA4/p6s+GvnFu4Ppwri2qv9wl5yS7
4w6dEiW/Jc7uP4TNhIdhZFvrbptZXbq9r3bUJ6Bf+Z3pgh23Glx/vLGsDpm9
xvQOBP4zYOV1On76gYVV8Ly6O50Fj6RU++Yn1MoEeGeIl1DPS1ONgUEMiqOM
v7xBTGCjuBcmuo+XcIeUKDuCEjOHwKvXwC9hnQfio7jDVRBwGhlU5cvZAcEZ
/u3UPVzkRqseq01I2iUZRQSCYx5BRX85YfcmgtBM5NgVIltpxan8ii/HPFyV
FbJI4PG9zrBPX5qg6c57uwxSFP9gp6EOcuT+PLgC6JNJ2oEOesKyEzhts5ow
pBQh4ykcniIs5E9UGV0fMCDQmRcVHNVi2XYAE8AIJJiDO3opeqXGwv3U18EO
TUco0VN6drgJrsC5iK8lqJi0Z9agr/TE0jnSmr5n4GMiqJh9/C9FKc9WW/OD
TH5YmzfcAuiegdegCcxdZ+9BiMGGuBghdFMrnA/WBJCmrMmW7tTS5V6OohOW
yIwOTBqdaTBnzHePV5gvaoeYsFxc66JOMyfH+c6ZOADAmsT0COqptulLHt98
gWgCb2yDc9aq0BmsVkaMy45IkuFDYDxmORs7gizVq0IbaQS1zk1t0H8axK+u
ENzTNIltIH/4/twyPdFMgYrKvxmH7KRq1lPFCzbI+FwvCVuk/2nCJg79gYa2
T1WOHC0CEhMh12S2bOhnDMGX7+6VDn2B6EoFJfyZR65jFs8EmCrPHxEt5PIR
aY0newqgehv2TeR9YUv9IMG+LFe/tU9X2SJUE60WA4B0edoPlwq/CJs8scwD
6Lm7HjH3YXtGW1qCYilJQlZyrRpoGGwnsY9yPlnKORFN4RQ8jCenpwm0oaot
UMajErwXbRTbUlUt1UkKOrgN8I7YDzfD6TTTI722+rlP+kmbzOEUu85JBzvi
a6XZes6prmhZ/Ml1KEnseEPH65ffVLIX5NMUQFzBw3qpC+hJs53ViFhJXRaC
Sh5RwQ65EnUe1AtSFoLmos4+s6vq65ZBRlrTW7osNJ+qzGHCeKdP25WHjYxh
8kklBZd8C4EVu6DR5WV9I906NlU9Ili3TdC8WJlc5AoOjfkqn2q4DboFaCbR
78NYNrshgF4fZ97VRlDDwlts5kFFlKBgto8NQt2AS7ece2vCGv/rMIqQQ3eT
hsbdjB4DA/u1Ysps94zyTojrZum7q1JWGFcnDdRQfIzdiGyOYzttSxk/yrNs
Y1XnkViTuGRIWW71keegVb7Uz1U+wC5F3P49R37AFHZxd4c6y+N9UYRC2qUu
DMY/1zdeygL9ThaUu7gaSv0slLQibkyuBxNSbWGWGHn3O1TE34H7CQYHFOAa
5YYnPks6EIZaxpedpkVUIwUFgO7Pnt30u+0bT/99QtSQcVovEQsXBzJoUSRG
o2o0QV0hxVRKHeo4TJxXDhwhnfEiQ4sZnooI0OlWtG2a/UA9QRGsFvpYlIXN
S92JUsVCh3g3R2ccMf05SrE68OaGKeZq/pxmsb42azpXgEMWDkzmrzTSbrlp
uVfprKQzeIxwKci5PWyFs7C6IYa+dgQZC2eq2bRXh1sxE+A2w6ftLruWzhlq
Am0/OPMCXORpDclYpG5qt+jaAyub4hFiJlhJyan2nU6JSt9QdfzAgIvV+lwE
ean269WmtZEfZIgER/rlXbASyy6Sz/CFfQcSRLrOkKX8PTw5YjwpSycfVmfy
JS/SMAmycy/OWoAioHjPD+qa4+rUG235Gx+67jJRynnZAMqpNRTkWYN2Ko/W
2XyBWvEVbe0sXyGpDORfPARt70QQBAyY7WCgRD8y99Q3uWj1m9eCxyoZzRtW
0YKh3oUBTGf9uUWhov8RrL0MAwnmmH/XG46zKHU/oVWmB9eWxdbfHDq1SCgZ
YLrf1H1eDP3hRAbGwXU1YY00TZfYJeCsa9fokE669YsfQ1xMerFie3q26dlr
kVx6LfunOpTIybYuUic0/bcV06iM5zAI2h03eBS2zcWG+4aQoHOBlQumUM43
RuDGlkPnZOifTAN//T8Gyc3va/UzDec9UUsOw6Bd/msVjsLU3nAPj3HHBbm1
z++cJloOgIzSt9vHM/quwizp+NtE0rFsJ4+uJmY/vLHad+m/UCKLommOyvUZ
XNdI6HAVqdJoM6FjBWBH5WogJCmOlC7Zb/RMCy0nJS+02tI5uCW9xn8PqNb1
hITwfLPJPf3J9RbYIQ+GMukdk4HASNHrRK9+8Oa+PJQzrh9SnHVqNIu7wOn9
0HP1FUHqa2vAE+HrILeoKGhcZ+PX5oIN5pnawtK+fGBTbkXZqk2fZ/8Kg/Aq
cHQx4YdDXOz5m2JXBQ5VF+NoZcu38UFzB/M0aGN55+hIU0AAhaQKFHcwmGr1
V8Ai3oHWU3QPE/oH0kDbJzdejSwgVYRspXcFYHDGoefyp2McsfJwP4tai9dK
LhfNt9PVau00THSTPtwBUWk4qj6coM3P3+ZWYp66LsyWmefKzRr9+Z801+n5
4OSuyf5LzpxQAp9OvPA+/t9AgLPk6kUuYZMO+AJXINwN4aP1azToLhzVuQFf
mNhf1uA+ryWMXIlPRZiG0yupdjaykvRnEUdCvJlTFN3JN29eIw1gr73Ttcw0
GWY/os4NO7xMndQA2C526FXQ3tN1cCirgX1y07xDfBPL3QLEOFl8jPtKgN+N
6tjjFDgPySzokxjHb2VEAVUHsJOQlaeJ3A7nNZD7kV2GAZYhw5qwO7BPSmdS
etlZ+EZqro/abvkO8olAwBWC63n8edS41JKjsDMB+Tb/2yYg29evGJRZuLPl
SaDBjF0WPWHY8utV4qF0Ce8W5pHRhMsA/D12jvHHa7md9c1jvcY5EnBbkLuX
2is1W9DtCovCvgC9MtKnAVu2ZCFiHL/nKy0TT6WFdk9LWKw7sXrbrzTdCSdp
EaYzGXVyvfDezBAstRfOSrmaqUDAwHEkiyztnVL8a/cHa+9L1tbTPkNVKEwN
BRW2uWL79ip54R4xi6uNM/hIIHCMUThfnaCANOHSRFgSTbY756NWLJOl8Axf
ydD4PjBggqRL29GMjzZQHAJvVICjmyMye30Jkjj+KK6M1CGlBTdMdQloM13e
h/pdaSNGNBuIpdYUERj9s8/HKcLZEaD9zMIWhH4lUKTDdmuldnmwV1tNMcm6
XzuegUJkgJESw9oBgl4v4FMsu+1zcuUA/94lqvw8Sk65GuJxiSXKmbD5g2MA
rSxm0fDW6tfr7k6Gw+WX/LlFL7mKK9ltf8bfUyx1e+IsLGOZOp0jdIm0fKEu
oKT6sUPXGMeX9olUr+99pnTbyTHrxfnWIx1InN4MPz029TCuwsihHTWmAloj
RESu3X+K1hcdvuwv04iE2L4C8vBUZIy9uBrQahdgEP2vAfUXS8V+yCf8CqT6
VrX/oTxKiG8tnGRn3iiD45Jmna0qfFvjq1COhupiDymHklUMYdF/dX9+akNM
1on73ekdlDV4RwoXk9TW8nCbOoVTSYJIKiILFEQlYSYlxqWs3kmbouXgxg8q
1HzKRYP+DknqJQi2wowd3PI+feklUwWiDuoMlYgHHZ4XrF/ePzNtzFXWiU4O
wdhFD+ng3MY3HM3fOO4ST327e5yXwl0FZzX2hxXZSCdvV3sHDYQ4ma7AU9fF
0kO910jLK3SnNDjA6gD9GEdczKhqM0YGzSegjDT9p43z2FyOiki00D4tnWS9
4XQI/9RiCdRIigTyRVdKVQXSP5f4miMfdpnHTDqhjo1I6ZwKiEbiuPIxTKJI
xdn3iEwcamxxJ/GXN2d+Is3lER+yDjrPG+xenH9d9NCE9ODx3WLrMvH+Vut6
1L9rQSdAdEyIORMDHhq0SZbIZs901ENVPAmAv6bPtrqXhw/GqsDmKf4n7r/4
jb1x+zG9uiAlEr1wmlIUX7mQ67T1f8apxu/NO5g+ohSdCUNFCy71vgXaRxSS
FJmYXGk8ZF/hPN5AenXJAXykZUHBG0xYYhq7vLxlZ3DTH1dnXbFb7KTD+koR
zKKjQ0952jiCgo523ejSZ6Rs3OPuqWh3gWT0gUbzuuxQhr+x6lVbWDcTmaY1
RUFsywIian/AuQI3cyhTmxLiKwHupcsU0nmRUs/9Zr7+Ft4sgjig7IvYmCNk
dGBVlm/M0buS68Wq66UekXcVZJr8x99UveUWbO+D0ol7vi/+U8gK39yrATiI
uoMRI+V0JuRCUBFvC3IEekTUqmw15a3TeP3v6BFlhOY5ok8k40eLn/RPmoND
0wb8Vrq0PeYLwf5241BT5YOjMD8Re5DwAeYo5Q7Qrm6g8fenkFZm2VBXo/0H
N5pY36YsydxCCue6397a56CIYI+MxITnaXyaVZZKiWa/PR6CbG0rw3mYqRyc
quh5IGYCe2xaOF22Zq9s9dhucyN0wkKD/UvjtE0EV54EwQ1lyP0ECtEAQ5R9
iK+ME+WP1vvEQceY9qHqOZOtGslEmTSIAJ0kgQOz5bwH68Jnpm36JBMAgs6j
hnx3EDSVnZFO0qqcP6ZB94VtgmzC3k/ZDI91pni2/MYAxyDhRvciCthe0hpn
tnsOAVSTxTycR1Zju7zcu19rmigZdZS4L/ZHqZKijysjZUxh28+tr456BWXU
fEnOL+BbwOSvBlmhEWbwRRz5c5XiQsE/K1JdKis0r/TQPdxzt0lsOarjRerq
QkDOu0bs2gXMUegrG/VPg9YWHnbeVRCBRjvfZemFB1SSK1aJmsE4eytmmWzb
H2Yupjw/U6BqimsQhfzNOfr8xGW9OmlxqL3QrZQud1Nlly7cn6eDkiWmfJuB
t/Ptoo9DyqIweCoUNJQrTsCw54fpKWX+UVYdcJF5SyYlkr8W+wYWnmFCuhI7
1y4gpW9GRsBT8z8x+3otAifn0sz5c/A5ebTA5jk7IhfGNcYaOSrISE6vp5OX
mutvdBojljXN2J5QwcRBg3vsgr5teeRIBVkd/QIiNddMfdpngyfKgo08MwoO
ABKvCe5E2ZO/+Rk4UPGeumtddgJmiwzMDJJn5ZML8KJhNvtAGVOUlnoQgzyu
XnMpXUzz5kKmU7sM3cdtzyvCt+ENrOsedctuz1c9QqDREBB74GNoVoauxaqX
2F+8mdUK5CUWnfipqhtoLTE4BhbAoCtX/Sg1qssOy/YmsvfX/e56TOq3KNtq
hNHrgs+pyYUJdLwG3aSKOWV6bOfMOXIQSAkNeinDze4w4sVcT2A9y9U1AQb0
YDmYiVgpTD4rdu5KKwhjsQihE9x1jCyrQvuG1fbfQ7TiYV8z4cpUqDgGL3pZ
rbuGFLsX0+19cC40HPNTTKVMdLnoLdYLYrEbTJdjR8MNR2kA5APmSdIWHVZe
bjiJgN2NLq56MX0A8go+UMoRvgm3/m3hB1pXQvc66DXIUOMV++Re8vzC30sb
4FbVg8fo9QQPMb2Gh6roIsDzojonTpeG276ViyP8NhJ5NcvgKFAXD9opBrV7
FNYEaDkMZgXyNUQSrRHSNiMhWg7uncJbjbzLsl5olvRD+mf5x+HNhLq0Fvfy
9gce12DLVps37/0FKx3W9sKJA6IaR8k78Y7cvJhP1ZUn6izE4Xo6AYo2j4xV
2mTrV1taNgAWcmI1KCNp4InLCkBe9SPW8B0Ub51itbw2j91PF7x/fN78GoRh
JgwxyUU4d6QiG/D6u7VG88oRTFQIzcaV+IP/lPCaqbelkybfVgvPelR8cxGo
qY/XIE+65EC9aXQT+UfnuKTc8lqwiwhi8pEnVMM+c9tNUuohsc3e0jzO2L6P
dFR0VROymzqhj4Sigy6C0/rJch6dxaPGm4BrkopqpBznSfraUYE7+q2+74Uv
i1BbYvPRfJmrkgkvKvU0+J8kXC2MqyRzOxytqHfvn42EktLZZwXI5FCeHKgU
luo1AHe5RxjPwk5am/tqobTVtkchnymC4ex5UNbHJOiVO5f0Spr9ZV71GsH1
d/J7gzMU/c068EONxfJfllkJ49L4eACmZNDYN4bR8I1T9ChsLH7XvHtiKASs
rJWN4rhxrv9xpNuhRB4X3SL41c2OnsSMJ8JxXwx454NuE5OQaWJrKE2k071O
7grGTYPoU3XMbxMmt5QO4/wm9PbcmVcXWxeOfcoACEgX9tuVa2ujPZMYOuYD
YdCm2lOeXh0EjQFxCI+RDXkqk7x27sb9C9LrNnSKgaP/VOFjPNarXmB7W681
IFdorNYJ/xdkuNp4BqJiapDxXNCPLkIHlGJ1i0oxXBOuS+uVxmlL/cEdNL/p
Y9eYTZahbNALm6giHdztYJrcKO+wboBWgBRhTGiijnRccQUdb26ZFhtA4Gy6
cZFmhKPOgpAxpjKCIhvLswCYpUwXK2EaKW5B6JkPQ5nx0BbEUKZ307x0JQfT
BqQGo1CaMCOJFW9HZ0BHiBYo6gX0g2ZKabF4/bCvRvrb6EXZuB9LHqIl3VJK
YNcaQ8tdtk1tbNfH+38C4MGY4icx5oI5hFLJUgBbE9vo5EEQttsJf9u0nBf2
qwne1LdWAJly9ul2nBQBJ6Vcslr4GNaHQQU9+KMLY08nvoYxUf5zFHpnDJzn
iaXmhrgdHwlRoF2NB9J9AihQUV6qwilMGGadWs2WyAizXLw4NfqqtSH2juGF
TjBdlISm1GLo/y/21eWK/R4g/xQVSkDFMi6SRw2qTx6BfoIHGkWbI7S/GF0y
nPxT99Shvfb3q9k1houqmnLqFpVtxNfCwqdAAvv1HHb2RrhbZHK/3ks4385s
RAAW7wlSbae2a/2xOuazVDv2NCKmo+r6HvXGAGeHh983f6Cj6l5rHsma/s8L
MKlPVmNSlvD2dg6i0uPBUNcsLljMWeKylGOsmffUFnf+sJMcHYZB/0yxYFtm
rhN+aZclgnFIG/B28dIvho/D4KV78pnpjjJcZf+stun78sCWJIb5K1OKbDrX
r3NLoF6EZPuorcD/+b2S5ZXWWsX/mouQ67LujQJ6rxXekAAPo2MCweRF0tqy
wUfgHFu+IXFhUUB3XbghaCKzIqj0rt0bk2hxlyWRYNp5dFtXeEeTkOMJsEZw
bpjw2XsIpkpY8p2p5I+5ej98qaKivFlHizEB4d16Q2zpi/KnqO/As+p55jyH
RSWwWox9fy3r3HRw8k2mPVb7PLI8v7kN0Un4V+vDDyQJdDq5I9l8U0xheLf2
OirqSVkzMATp8qiBHVNYV4jJsEk3F6+14/ToWMpFI5L8JLUOBlyyxhoJ354R
Nug/8+LrPPIqB2a3pelCb7fStGkEjVpnKo5DksZb4j9SSm1lTJaupNL734OB
WCzE3ZV6JwX/fexCNCfDTkm+3SwjxpbfljS3DbvinyhpV1PHt8PMP5gSuxkJ
KkZpZe3uP/irj/rACenIJPSXTZC8h7xQCmVqHjDrMU+qA0p1aaKbBp7S+ViK
2preh2pIMrGrquOrF67DC9FZnFkEgcqIOdH3gKA6a4Sjq6Q2qkhiE5gEsZns
nlbFWLYu7NHTEqhNSTLVJa9ZaMztWswZhy5MAG1FIXzkci0sHfqgQZw5WUVY
gwiD2e2PbzZCs5qYKsv78rwdjp5zbplixb9geZfCFJxJhDjAa0J7yv/g6/OD
rZa8I/Cr9IzxhTh7lpJ2tVl+fi8+ns2AWC61S8JoBeogU8l728y8yeWNn1Us
vJwSEvLw3+SC8BiO0xLXE9FJpXhklTyvZ5KDcwMHP6W8Mmh/95Zjw9nowJgS
gEoIY80VaxaDqY9Jf7qkvsF928pndh/FJBIKjVJoBjqXcqyef6S++QI19xJf
rlmkjTGqw+kvlg9nCs8DMgwvxcKX5ag8o1+cQyPFCOojfZtObFgcLXBJnRRm
wvf0HiiCdvHIBEm9rKS/SkBMh/EprOSHPBUdvGtqdIXLjOulkLPFOQDciZC+
tcVasQsEvvC6VwoS4IAQy+GjN5S9/1QjHpcm1t5BoW8zej0WjBNHObPtznM+
Ac85cqYGVY/P4BpdJ16erNbW1NKuaZiB0REHDauPV/t080pFowFQ1Oi+fqAA
whDf/mpeWWg+djH4Xwp+qiaw/SvHC+cKTw8fpWtSK4+DpTkB70Iv7C8ooUrH
AFYxefNL8K7vefn6OXmYIA+x/op6g08hziOKSAo1nhZe2EGOLHPZjsvvuVZp
3O0miNkRIXd5K2NBH6cij2zUyGyBgxR2LUiTgPNCDpSk9QnanNrMEWj4rV1n
X7RpzN3OqPiza3FyiDt4eQ+KsMban4yUQ6ZItD/fr0hpC4RSAX7dws50GUTB
IJPdINXuTvaoQK2oi1DIqnLoYdyyQSI6GiB2b9LygftPZUuqUQ/xQcTfLQea
y5jKU5NmPCy7r2duLhO8S9IPmrmb+CQ21Y2n8CLu+pwzHtv3/orhhOk2b0D9
LfVUT7FS0GuGhEw/GBz9XrqvjtgVZNCCPLZuyx3nNq9czWLJaecNCknYuEn5
r/GlIH/AdZSfxAvQBnRsEhe1vkq+ZS7FYgRewU26iXII9zgvsyy0/og+NWwh
jUUBYPPUn8hg5HDUhR2D35a4CcftGibnMHzRztzK5QCYleyAwxlp8tXD50Lm
0VoexkNYSM6CKCUgHQ9VH4G5KpddTHBEltZ95aR15+wbwoZlsXaCKtsle4WD
zmeID6/Cp/uyb3HRJ0ulmcyJU+XIrqXh8lt91ihRuPVWHe/cTQemcRB2mgsO
0NddQBEfSAaXzZlQ7sGZ+c0Kjz3zgwFvXq/MJMiuhXROC8LNBx4aSs/NLR9T
1WySc376akeaDLgfMKK+FpYsD32V0oHKQ91YgiqnPriSVy7liwSue9DgB5eK
SNaXhOdHwpgZUQ2yDQtPPgUmcDVcXFSY0pRj6L8LGZDO1OzC+SIngw1Itafy
rRSwii1fLkn19kVO2s+XfuKT2zbGAamOQWumllIt6W1HV8sUHImALreFO6LF
Eq+/ueymOQgy1L3Wp9AzRCID4ZBaMYR9hCXegUtfGg+HO6BLzT9QaMs6CVLJ
2ozl5SYlTCwpF6cakp5uSY1G7SBd1sD9Jx0a7AC9mgg0oxx2IPWyydYVpCj1
6ypOnj206yIqz252NzLV3Fd/Xj5uBN389nUOSpd6+BoCi71M/R1ZoLnRDfos
JrYLCAmzK9GXbG2TPHHXkgr/dIW3XGZZe3QxQFO11zKDpOKm+EsN3q5aZgf0
wFjWZLSKuXv1NzBC660o9OfQs9Hqk0pT7r1EvjdvoME+AlMoM45rc4dSyNRm
0lTuSpBH5aGy/MAzM65Rd2sz3zDKvKKCqqR57dogbcdwFMN67fknW9gdHYc0
M5lfV8IIaJ/R7lQgONC0i7Y8jcu2jopDXV9wLfbf6G9ofUWMZjyzfKKakqVe
MR2rdCKbF61ANpcB3buQ9w1Z0WghUeWilpYHZl8YHAA+0nRYrSQcvln32aVn
mId7wbKX1uCSpXYl13QAHdetygCdNusntAbvNWdHsmyJ0bF1GVmteZjMiph0
2GyPkFeQbXv/5yvqQK/Tsthvhe3fU+zildaKbklyCAOIIDH3EC666oR/f1OS
uUhQPwBDftoufVGnMdu1OaqjfnbP6vYEbyLEJfn/4DsT03C5Ohkzewk8B5J7
/apSU50iCNwDKQDex78Yc44m0AaIYxulXbyrPrmH2ziuMffH6n3wJHU5fwa0
dAcFrLuB41+U9O3xT9UjC4b+ADJ+tX7/xMVz9tPInvJ38WXErBLs8Al1LzvT
qVvfDOWIEIuKV/gUVHAOqk+bXgiwct36lkGVS0tmuOmuKpm/ullnJO0evcd5
MNBtGwT2Inm4c8euWFVrpHXnOKQlsVkL+s7KfL+vQWB0Al8bcLQ5DBcAQMP7
btHyIL82A47s4g5fNvyvY3lqQtk5N+hgFsbiUmr4Ou0I5nvoERnzTCuJMxrq
YcAw+KrvxmdSztVNICbMa7WxGAu7ahTDFrJiHHrS2wDzY7Jxj39rlL8BoVwg
QjQuzSGdAgD5PFrqGYNfyy84cEGeJ4Kz71xCAOGXWw6cWh6ThUeIYzgQ9/cT
vd30z38MbPlHDUP/baCPJ7EzrDLoOXwi4yENPe5XlbxqSdRhzd7T0jkmvR3Q
/wA6trmNidjRvyVo8aRBygGas2I/wsRczwb3zyobymT0BNPqoS1jUm+MuAsz
IGfOHHquLYmkPQzTnJQFt0PvIff/HFmjr97y2WH3rrhLouk+Ppbz6XekK96r
ndPJxcM6q07lPUE/OaNgmsnZlfvrFIJEb0UIS2k8tPNQwgbCZbX8xkcYGqw1
JCLMN8BIAPsNj+uTKBMggemfwjW8eeETsltkqUyk+miAvu9FmxR4HMFKw6cX
POwyB6EDcBU/BpMFSOGRrDsGw78fqEgAhuOZUDQ0vjuoemzbxpu4YNFtGvrX
gJynYZjM4NWlH9xs5OzHTNXE4A5XmfU6r+g0zQrIDGyG9ncfRGzzu79wcIvo
kBNIdrh81FPK5HvR9PSIj+Wl7hM6/rB2Ut1PSFpN9NWtSYQP93VXkHe6ssds
xArMWqygc7bryP40yITlOnUF2axNBXKBxyhcCBQJxuZpmgsnM5Lp2u1pf2A0
yZ+MUo5OSOflw9loqf7r4LP1TFzG18RU5+YQhTW3v53BNk0jFbmqZVsADpU9
9hp57H8dYCdRpHFmIrPgfqouQs3l/Ob2scegkJxWWdlSiFtJXs84gU2tmdvk
GNy7Vq47sJsvC04lqHjNfpB78JkISmJdsGdcF7oue3WkhCQpcElWhpubPXXy
BMVqiqz0l3VvVEhXfsTvyh9PUKMzR0EmW7ENA4uPEpQNh4IZdvSnSOVY8qA7
btDpjlgwPilbZ18QSBswX5YzOSvEIFgdMbXxIfJeOgs2HZT1M2jM+Bim9A7z
Vc17xk5+XwbiEzRMuwKSWo6Bz2ukNt4Y+Erp86bxPAiAv47X42BSurVv1gms
19eH5ezuWxP3bXUCS4sRzx8NdkykhtnV5cwdCBINojh+HJSnRgA2n/Q8brOH
vOyi8fTZ9xmvMhAqgm8EmwxahvzxG5TriuTkLHffRK6c1+s09bgTBjuInXOq
17btMm+dHyYBOc+IkanZUuiwMObhvsL7vNrgOb8wKLTNSgFnPSiVf/Z36NBU
P7aOYt8w/c9V+aneVzT0hvt+cxXh508oaqqTWDCu392fvi7W8TGzQ0SDrdUI
CmTuHJz4XsSXuks1LRhgP3w8+G7nOT1aFDrAFv50k2f9j4NWOLQ7UhJz6KM7
i9LPgEX87lauZuOaGEzubG8ae62dFPKAexHitxiuQZg63Scog0uE5IUvyF9y
KyfE/0M/5A96QGx3FI8rgj5X20DfSYKPZfnS34JacLKnLSMEh3KphchSyiji
ijI2gJXc5GkLRZlUG8nApVzdPYlqjlZhqr8RWpPU4ESAhfGWN4ah+nz2VLXy
IQnrSugfTMeGHtKMBVqubsuqogDjuFnJnZoqn5tn8uqyx/GT50U3N48jmicu
TgKAekMNmCxrpQ7tADzXVqhTt03SsB/gTyT4/tLRn2dpueK17BKeNAoHUnj+
TyZYT1fMYKyurrr/iMVHPEoYny4J/aPy+PZBIyXDRNcYmUidxtKHbIozBK/9
37NMWrxC8eFawGaxUknN4Clljv1LOfnaxvevs41Ti3haW1zjWtxinaNBOiIZ
+CzffiKzCGh9HfnI7eJjibfReujg3X50zjJKfuHPyUxSDptKqTkykR2M2BvU
+RrisBCfQRADzdQuropeK0Slu9gOpydgWbzkJRgJrGvv3YOG4bRDhLOFFEeU
Beib9fpAZTkaai4oZZDWBrweYBV4ZnLbUsxZd+sStxnjSJjdLlI6bf+wXXam
rlVnN4YKemzpYndBg2VUFFrK/A0dTRh8VAitdiNxNhvci31v4oxHAAu14v2Q
6qaa35Y2ieDE/ialGDl8WpcbUaA6h+v7LsILKQ12ao7TQoOO/0LUrqW1Ix6p
euN4fASJcYthdjYCeZFRC8vhxCvkegV42glbmISVtTaZpyW35GVWpc+wVr+w
xpf/se4j0KVjqK5akALGGwRCsYuPfucnoVpRYRlp+yKOaTrrkhn0UbzfwlDy
eUv4yzp6nvVOHvLFuB6MEv+aQjkWrVRaQbECAjVotd/q3t1pOPzHKmbaRx6b
wrjtHVgUQIv81ci08Ddp2UWwcnOK78T52Y8vPipghcOmMgxj/bShcptSrJsE
3DxknGXoufOMqQxR66TBzrxhizCUy1T67Vyrvot34h7HMIztR8n5sZinFwIx
O3vTsDs+v9ocjIwt8kLEoaayxKkApZOUwaICHAhjOFLm+E4hukQUMO8xws+k
ouBBkWCSE90qMDOVxAJisJXGilzLpIDKYh5FrRbLJ7GevafV5dZxGl/yZZcQ
xIzbit54rc+8mWoEO2Z2+ElQPpu7uoQVgCfznnFlfewT05Tw/n3YPT8tVgH8
Ua3F5JLQ0VD13QO9SQ492Cc7zA4MLXhzz9a3Y8sRosH3L/alVRKEjyr9sYbl
++3SCu7xu423fHYSymmeKpzZeWAJP5NZFCJiKlLRGEka6pIxrgLRXrXmSypZ
Mh8PNdP84gZKFZmheqxbMRTmlW8RzHzQiVY95V6ZiH+whzUm3XVmIDAqQ11R
cR8Xpln9Ip5G0ZKyBiqq2Z0PbnCwsbsuCmm9J68HSSH3g5gVfn5mmUDVFnOU
GmUqHQ8rm2ri7C3Or5uidC3FMdU4Y9IfM+gl4KFgP4ZP+OtagDn4gBGMhlP2
GDNk8m4Kyqt8L49r15ERyAEGLfl/KHtdLIa/RiDptAe17P2+lMgd6NxjZTCx
dP71xtMXBXl4K8RUV3qewLqgfqCrdGR6R7Q4ceKZNQBzXRKwl72UpoU+91It
Ry4E9PIgvP36SWP8QMR7BIewFljsFb8eQ0eNNIPSApaPd9ysEVki3r5AOns4
2WGtLQlfPBxiIS6zQ7S0kL4Fry1wxGXISuWsO5TD11zhgDOHST0fClsgFVyh
7pdO4kwI8AORJSThN3y5GGjWcXm7xFN+jwb8PVJGYCqBEmvD3Blu0uvYwNMR
7WNceYCkXOdDQLLBkLfeQlCWrlnkgmlh1fPMbLY2S6dxQYXpZdUnQJ8xxhPs
N0G7Kk48DKRNXmhbpDkG1wMUNF7dp6oHxoVGp9qdo/QLR35ZlZybP2jtSI9k
RXYPQ7nsjjGSOX+DsMbX5wYlM9YR1G8iofAIN41F4YSbU+FFhm6+roSjl44a
f/7ggxeaX/05Ce++Ov/6quUPobPb5vhF+2bT+gzVmX1rotjQ2h+8B/GsvBms
ODutIS+lUd5NeYcfpQT4aE1YA57dAD+5UndikfBw+d/V30iiPzq97awgvJHK
//l5k+oYePVzf4HyUDnGCZWZEmzhzYEomgttJQewjyc4rHIT1MKlHW5gH4vA
VM6+V5i1mLtAtB91EKtrcNWwb3CLC/jvIuKWRRC4LyMtGrfQdUHOFB9c9FMt
FJRRy0aEzu4nOmIKfvk5keRCI05Z96FetvMw/Xuhd7g3bm3NAo4MXI2zErC7
BV9bOO03WqcEvtEkaG6kF8Y46hNays2eA+m9+FVg11D7/OXzFK6FDIIIUiEs
ttBGqCZiwWMLNDbKhuTHXp3VEp1ZeimUXnrj/H+bS6X6GxIGdCafqAdcm2o0
6pQLPQ9T3lm4hzZ623NqmA3+sgQiItDONkfMvu3j+5Iq/ICWcjk5k/r+aakF
yiGepAjNrYKu+XCY4NUMyICJgYcefzTuYBiiWRph5G+5v4c6gOtcCEwhelNM
zjUEHa7Kmd+GuX/bKO2EEeoAxFJDCE0b1NUTcrZVdK39p+H8N1kgnBkzvVL5
JJ8k6Qld5OxrjoM2qqFDVrlVbhoSzCJzW4mINrIo+T1UakUw0tg+pT8EMo4X
opgVFtCwS8wOzcR8E/wB8ucvnkD9/JqbxaEmGydf3BmlCdBKEL1WHgFhvTye
h9S4FVi2ITaCc4seDKwwv/jz09pV8FWfs3Le/9T2WDgWWrH58cFFwXisCXLt
q7cKWUMrEwjRmd2xZzPO9AcIIgDAFfqqle3a5MnYEx/8ZPAhc8KLhJItd+3y
fNwh4R5AmNHfbQ6ILwxffpGA0svV+/UgW3XZ/+01Y+0plsRdGH0oF+0njA8u
8GJB1Y7B11acLCqG1ddDnTKIp3laAxFluoDKE6O8/si6WzqUBFNQtIRKBobW
3umbCVxlR3ijO4T7zcdKs3UyouVelpB5Ugx+umLuQ5Y/tTEZy6epfIIwz/Ig
PJj2etFA8GNWyexuVqZLzv6ZOhO4JYmEn4374B6XJjhcOh6AEhzz3WHZVYpQ
jRxGDKv4AaZubwE/eagzoIzAkUUngRCBupjy+n68RsK/sSt96Y+sEQ1B4Ua6
isIjhVdTRPmaHD69SPBGL0aUNmFKFrRe0wiWPlADyYphmDgTz+K43JM316jh
JciHp5OK2h+HHBxkncyQrYOziGeY0q/DWkgMBXmIG+rMBmCQa0n5YN1G58Oa
mzyDeYRHqrnY2gDHuYMaCSjWqm0WgKvMj8padkP9VyfoVD4jprcCcjZdVUZK
X+SuG4XK/t85FFTnMvUNNOKAcEKTRqJv9xpcgHX0rJJtwe5I33JeoDbPZwI1
z89E2wWPboQMySbjSN1AEMOHpfEAL4dFSz4kaGktBYWAvLTyiNMW+DQQ4CwC
ZyvR3fDmVwTdvu5uEDGf+9oSYf1rcBMQdyNC9RtgEBJ7e28OQMyIxHF+db+h
puGgc3Xuq0hCo9u0Z+agsM7G75z19zB/76o6LCnBa5tmFFiwYI29BM9WkL81
CYKauBaQHR8KPBzUDO/9AqBvDuCkiheosu3hMVhYjOJ7DNxuN2bTDwtW65ha
LZinAgdMRfyZrIdiyWYsWaCNXltVGFULl31zKDAY7qTN3AsI+r8ZPvAort9S
vlj9nq0kDOCSlKKrZmRunk3dv2z+jcEuy4c1VfN07dRXYJhGXR4/29jRZs6P
6JWWIJnovn8dD8S5X9K6lc7yTaVx+MCmdskE0jdKk2y+WHHrlAwXnjG4ITpx
Wo7xLi8t1Dhb9Z5V81eFFjXXoGck57IYBNcAYJBkJ8MEg4V1BE81mOFnbPoi
i04GYWU0m4iwrnd2t002CyP1bFYGpKlZQ+rfJ5dCNV8ZXdKf6w+TRI2qzK5N
bZDidOKx3Zos02Ba4Lah0zF8FUbLUpNKRQp1BViH5opnOhqQ4BejOatQru+L
LrUTKcrMetak846JDRwPNzy5hMfmxkXdtrrGE5F3tNkADBrbuv7fBSmneDjP
PrR2Qu8Iucyphb0QR+GNaIaNQjCs75369sLDFd4H+vHEAMd+7T7BD7qkkTAp
UwInK3pYVSHD6fkTKF2df8TNGDZHEF3lQwi5Pu912N74m9twhmZlG62uMPWm
0Bm+fuJv2rEb8XRSfSnggcijlFiHyutkhNeT31epcgtU/eckZwlL4p5IFVdj
MhKeCxBWyM7q6BRHQKxrHDVmCJExelqKGisVBilBlT1rEMp66XV9yv7F73ek
CWCzzL8TTQb2LuvZ8yhJ5Zzff0t1BM3+knylxCAf/hZfGItkN0JBiNrloxgQ
qdEEV9VkijqN3aaII3hbKW4MbBS973VB5aIluPi/ZkkionC1EeEOO5vO6AX2
lhDbzkkAA/HTRYZ/cvsp1FLmnApSRYDfUhvbW7ktm1FmewTjXK/9Ncwc4dgJ
nuCBEg8PbskeNlkVkROu3GjhMMqaWrge4pHDTBgsig4fBsejc9HLS5S/M4Zd
0ItDEIRBoD1pUKPXdBfy5Azc5NbNndY77YiHUp5+w+PHBYpl62Yq3ErZSu4g
MSfDjHqwICMyup2TlklW1OuhlF1GdWaTYolRuEL4Q2n0Bva1Ybt4JF4UySIs
LYG1wAmBIIxyG4jl8jo+nH5WrxwXJHGAHgSIveAuQwD+dKNtglvEOJb2HqL4
vdhAyQa/ETZAQlUIfxqJYcZRxtjkLyJ0c34WqaILvfJVWcYcJWEmKmhizTBL
RAqTfJiHmdIexh+A51b+k3OSyHOLwlBtmGE+XsCaAGRLFS8qtvpYa4CCFXdo
ven+ctnUkChUMYHYxdz6P+JNK7hMYxAcCiBUNFaLRw+uyIEOlGfnTEs2QLf2
Kgn8NkAnE4dduNC3BuMYfR7uH/Ggwf4mTCtkf5pGe1mj1vsSlat2P82k7TN4
m7kerzOKNTxpCuVZz+jY5Z3sWfls5BkwnBl/wcF1umOm5xkwGVoiMZsRWoLP
xEK20e8XE7dfzwfBQgphjcfN8FJfUmORR6nnD7x4c5er/hJWeR/L1vNJICRi
8oepZEH0L+78jEyRApC3FTpNIaD8YaafoIWpgOKZNNvemkyP4EPXheFJua6k
hCTjggzb66MjAWKL/1AaKXkq9FjeU11FTZLXn6jgE2+YdaMUB+HoAYczvVR4
LaDMIbN5Z+DHnSfGfipVk21RtvZu0k0/+MO1wm1FXqd6ZOh9RrF4kt1rawCK
UrQpoh1rdguSgH7OX/4NoAar/j4ykr+cKyBMtZAuY4/t90GlS9/RUcAwD8Sx
UaCHpypltHKRsFcFvVRkrX1YTb6EoaRcJCStxcfOzb4Q//qErlHAWGlG/Z9x
m6WWC3zVvgruBUs7/4tUv5zeM/kA6He1sLZg7W4Tnm6JlkxJ6ZEu3irk1e59
p4vON1kQn+R31Ne8rAGn6nrn469cXEnpipPZUDSK95P6IyyE3K9tNhewzSb2
sc68miu0+E5924PYDr6t+sp19mSGZabsOSyWz7RBzPmM/Z3rYAn/5j6PM1U9
B3x5eyX4LCIz6xCw7/UMq8DFda+ROK/tj+hdQmLsy8VP6s0iq80dz5rT1P3Z
zK7gMrTtn30TPgplq2LRjbNXXNi/7PyT8Ga4LYbqGcJHdEOkoG+HSC4KsVot
oOIZlsFBBfyzfZTh+iayvTZ5Egy5XMYp2zhGDHpN/mOR0kByz044wiJoHrKi
m96yxdao00NFxGp3dnper39cVqDhvjFBEmZeBdVUz2K5bn4sxjliuudOYA9N
UxUuecZJPYUCdP+kMiiM/DN/qdQq0307s4afQiztdxxDjdKGXriXs3cStPo+
yN05bEiB7Ua+aKWljNsdIuBJYmZ4MkvJWXe4dL3bcJ9/0pl06OREweAvzpnc
6E9+GlfZVqzmiYbeiDz5G5j0c8z7HW508uTfGbJ4M1GvF7HOaF94TkvzRH8y
5NKBiSmLunKyI3oOtA0lQF8NVJ8pf1ZgdokU+slpOjjZl6b0AXYH/em20BaT
06Kiy/mMFisIHxIy/Y1Z2M+DtWGHrxAieZ+S51AKpjWoPRVat2F1LbV5/IDw
TZ7jV99SL4M3I0BXbUz4dIvT98BWhG16JGWz3QKz0D/GMBbp7c01bQPl64Xv
4/BXDpEcU4TL6trGE+xdj09JsEkSdtHupBTUAu30vBwR8PxaT0TonyaiZ1yv
XP6kU0I9YWj109YLTtliaTz/HXTX1cwhkx9ob759JLUV/ytGSuL5Y7QaLiy4
VEhMAPrrBoPOKbP+jeoVQPxQMVU6Mr7gyYpB1bt0A59/k6mH5Fz6dSBwX7X/
ZEjaZuvwnompbR8DtmE4L15GhqROyuhZ1EvcqJGy1e6jorLgkB3GDCzZSZAh
DmLNH1Bn32AI/kZ5UTmKrij+CEY9jweXsTITarlnUJcHDJMUZjxW7A8necHi
ZaqPIL0MXyfuLVk512XJbeTH4CNPM7GuiCXYYMsumGbQyq3rPl4wOY2nUitD
ipCL+9Vo2E0FgGahhw0iHfST/DatwQMyhvjVoimfk10CI9fhRQwLspnFFuXA
j97FoDcUdOem1S2Z/n3qFRGOAbo9dDWMe/7nLfp6Z1rRlwOfm1sqF+y1Uyjz
zOxK/+LNYJ13eIdCg4F8yO/FoaxsKBMuh6SBA4ftj+WiQj0TP4JIVo691U36
SSf5rFLMwdkXMgvjLUj0CTFlSxc9Xo/hgzwAS6cFiun+ifQsovXDt0dqCRTM
+Kw/Y9ItQd8VvuG9uqNx3t5yRWzj/YQ188tELD+oLn2b+bYcivw3O5jS02SD
3zpK7IX40Og3w14dKARPXqb3CW3NVD2rE89SWoLJDEmdSboI7IbR9RJU4Kwx
TNbWro1XZvwSEluI0t9bNAB4fVl1KUZdZGAYKPTBLuokmGFIWv+BIym68iQA
8b/7lWlVAaNXr94ZeaURjJW92QOwbQ9Rrqi6cwr1T68E6fe0CvFefuULf1dn
gnt/xX/ZhHkl2rVKTJYpfLzf9WvghnBv/BFcWfCXeVg7yhq3pVON3Yw28ruY
35rb35qO9Uq4oQwrmxUoeRVBmB4+5+lE3sTX88S6ClWcQ01KHYGm2IA/cDFt
5YHqCwlKpxChE3aM6ALJp2nhGH+9ts8m+QOPkR14SheNRwmPm89v7oH8BsPo
s0AZI2w/ylQkDw6hveJDhF9icPM4X6DvhUGPijKzuoQh5ZssGveWGKiVNUd+
ibeUhZ3rXorZBwwMVzDblvzS/MiKERhm+kQdBy0VZl51Fz8w+5KIss8goQcP
ZYP2vDlWCwbuMJsJNSVNgaqotvR/Pndyr3NUsA9Lpqh3/NQiYJ0Gm0/L8mHX
F3HOWxR90iwA49o4I0KLFS9rBTSK50vzOL71YFtldlv/rYIaSIrGhqKOixNk
tKeTKqdbULxjL0g+hAayHp04xaKxoX/kL9XNkZZQbbc6xChEZLjVnk9SWmw9
toByZSzvQCgUT0MnqpKnxDSrHFBuhQ/p/JBvlm80TZTWAxQQNF4MQLJzSIPq
iPYfCTf0U5m/Qy+FhjW7Ujsu1Ovb5sPiZ2g/JjVMXol+b8iIXZXIUzNayOCR
3sujHvhSRbDzfpvF/9EPunQZmB+COGJtfVS4stfy5JO11+D6zenFBROUztSz
pwts5g1z31BVFsla89TjbkfA/aPzp8dT4NjqXSl80fEqtLna2cy2Z78oW/pR
m+zZmYhT8SiKIuw3WK4MvopwgJXETssK14HwXzPUP56OX4z6b2yzeJOC6l1H
D9T902AwZNvkv2XyfaO1YtieccQit6iZS6OP0R+WIH8xKgkStZDy+KM8qJ7U
sgtkCs7Qqi2vijNFzv4C0xp8sez+vjtPqiMYAdGMWCkz/e/EuYPBtgSAZipL
FqOxBqjrPEypWKy6MOujzqmcSDXrBK4blqTiMCC+Uzp7PL3bYw9m+P6BPldS
XyB4hEFCEu4MzZhVU4fIGSLL7pYjiPOd62+uSHbaG72LAI9KSFWKhnGYYJZL
1JXfpgaLLnCV9Ra7RcWPhB7EkrxKJkK2SL7V+iYGBk+yaA++ZhdtgvCF21Bw
4J1SOvJ6Jy8HhiR2jQ5J9NeUYQELezdAVVTM2PXHZcEEwRkUUZduzNhVChkq
ChbjjJl4FN5f3I3olkBPHc3j1HikmgimEfmJ6JbA5nlpQoE3ae3hdiU/24gD
d4CDvlO0DNp7FfbYFR1WurD8GrR1DWxUc6pJW/pXI4xxEwIeptmtVjDqwVKp
LcXlQCBkRJa1+Q6NRPgknhOAjmC+fLUnelzlvgJahRuZMj7H5bPQUOQYPiL4
fyUuW3dkv57bLChvZhphUroVI9X0K0O9u7fbNMmt8g2FWFaBLvGpifIn2YqP
Og0+oqMWBNC2UaX9mINLiEUxtWyNVsgBjzBd+QwzcngSb3ARiYItiXcd2XUk
pfFKWkad8sr4Lu/y3F3XH0qGl+UyAVb9m+dhgUdBwXPZ2QvXjdS7sDjz0p2D
7Xz7sdVFP2NJ1O7n3uGTlg4Jd5AXSI4WusGvt7vXm6XXUykGnJcDoyxE8X9F
4MG5VVPGxlr5G1+2usPRw46TK7uK3FriY3SL53B6Y0VvvLqGtH8WR8OIYKjp
Jt/Vya5j82j0Gv7k9era/PZYv8lu7WlSKmhZzQs0a3xgWDr2EyOjkHNU3Fva
05cJklMFfUiTAEiGtnW5UcIKndTX/u0UHwLiS6hPILk8EowlSq9KKjQM/ulG
7ftEe3RnezVbwL15HQTysQEZfhPhXaO3viK/EuXqWRaxVtglxo6nzxX0O1Q7
ezghtg/GWgIf+UK3Zfe4tJOXVHhN5jODGIp+bRERWdzAjahxbI3P0tKifYso
fg0OuIBmmBD9uBJ+GDsBidPQKAGZezfWeDCDxPC2TuRYFvbRinkKPpv3RxT+
haBKXHxfSTrU0Q9fGf+e26WdV3IAiJzRVCIiiPLVmBYf93G/NW2IhUp90LDw
BBJRd3vAuVYQfIRq8Dm7Y+ExyG+T4SVzq40/46Bx9k6mwCpSR5NwmPEZPaeX
rzXaUiL8ky9CcMpxX0yJ9TT/KyWVgc2oJKjELKgTo7Ve5fv5rCt7R6cSUdUf
lh0kcn4ulGbqFKmEdk9F9ixtRyViOOfdGUGD4eAGWQZw79BV9jQiwUzGWNsH
T68DZQNvmvCKrrNgHdP9UYmeXlVHAO8m9cPkm7hetn1QKxaEXtPLpcG5ZOMt
C0Ibv6aXRRD2V3Jmq3SoXfZqBpqtei53W5f8dznqPMunhOLKMEDew2Y42Fc/
0NLXilmV3JG/7EuDkFyNqejM2XR++2AfyPCQznZJRUca+Z98ulpK4b17eoGx
HwE1FhrLxUmqm+paR6LDx4h31koRSyWTXuFBuowiklRHzJOP1Kk/FeOsG7Cl
wbhWr2fFO5+TK4c1iYRD63IrPECJyoVuXnnN+7KFN9BzrDBdE4OdUKlwHkIV
T7PiqOj/LXorGKLuLev/TCDXzPDbS1PJnjDr2XXrmDoCc/yyvKFkZPz7558A
0P98lxDOBubSu7a/+Hx8NVc7mSm75mGgjUySEL7xi/T9eXMGoqu0YjEf8f86
HA0LHgD5zNMHec60VTDLrmVTLqmEI2DK5Qg3kbRIrBCfoOdBNssrWji7Zz60
5f9810dhnWUyv2l8QVNVEFM4HweFv+8awDhyw0LDcwsDHCCJChF0RA09hV10
39rlZc7qn9S1WSIaa5qVXhIWQxjbvBNo5vrH6odXB9PiFEbKbs440DNF7UuF
rtyomSctmixBnRV99QVVkL/B6i+4DzDyl6YtDvfeSfOULPN7M5khAoO8eLm6
HHiOnW/U2xzuvmub4iLvHxVe3drdlFYV8VtQGKncSOgc5cft7n8QTvaEbOG2
1jEcOlK8FyncdBXUMZTgRmbEYc8sDNwPzJcLsJ3vUWbUqjQbleUmdnJd0fnH
NYz3KVyhiOnxzxsgZo1BnYdnh5681UF+0tbFZPeDjE8qSgs+dMgnGqwM/Gif
ARG5WTTVRtvV9Ugs2o/yudn+ibOgEMoPWs8Gi+46uG+PZZF8SFc04MD/55xZ
Q/ZhX5l1FYzgDMFYKj+s0gHgyKrm+abLPimD75XGY6jOXX6NaSN86c8bkxAI
KMHLrVcFkhJJ3Mn/QRyWMLgBwiowK09RkTUukXbEc2zakwWbp9qyknKSiCwE
bWKkvTOb1GM2YXWz/7LM/KSsgWwk/xK8JwwT26r1Ky6cwU3klg6PE9Lp1s68
1X16aRffSuxcIqg4vU9taUo+OuVZH2N+GwQmynjgDmnZGzQux9UZ2Hv++6al
ghsY8Im4t285F0795sZHJdzxkUdQOdgqoE+mIVMpfSPaB6nequOsiKuzgZ8K
YIYC9kmO/8jDzxweuq/AhEjd7BfzxFesgTaX9jVjtEGnU5WGTVAwQvLSrgl0
72rAsMp76iHctf04LFPLugpMFKn025tZ5tB8sBE43WMUlEIFgoAvC3OQxtuq
32Awmm2fGLOMXqZNlf6R9KhdQCjupCsbToi9ksKH6l4HOEKoIKU+l1TLPOip
ou0AVQFI7pnXYOGwoBJMZElcTH+jBer0IbWRc+wxwZ0KdMNss4RGqTQ3FX4/
hgJVQTP4i34vILDkEHExUNThDAK5jE/bNrZ5wt6AmFBup6nyb3/x6NUgNBZY
vyMLJxiC52bMuw5KjV28iF6w9QiW6lZVQBE9g2UobsEfnRy/J7G9hXAR+upW
U3uqhpwCghBVwJqfn64N04W4wA81b7+75RU9Cw7pp+bXu3Ra9mHUo1hCabbf
Ye7ZAkIZwtH5X+7roRbnw1ZuItMm5ubq58jfEnQkxNrBhpU26D5oou5gKP5i
1VvIgAo8GffSjlZpZR5HHC8W+aKK4VHbTUH0WyFSDgd4pO9uoKA+tzEZikCI
omYtfNVFW4PJSbLsSnDcTSVHj6Lv2elgNXov7FU6T14M6WAFuN+i1Oo39YAb
RyTiozXFF4ptQpHrfsQFLYyONqagEagXtDXCJ2FOr93PY5mjxZ1ucgbgpztv
JpwGPb88s5qeK38UFku/EI4W9xQR4HLq+edFFrtb1tfqHdInuVJLTWdzOUvQ
62T+zpmhTxOJ2NzSHQrQlicHat01eg7vAgBwyMvS6/noERMxkBSjtRZnTDuy
95tDDP8UPt3QVmbuKWfuRfNU3Fg4IpfKUmzBxC50M5fJa6+wT77z1LBSwRpL
iP9Hbdj3cUP2PHcHqk+70/UJ2J+MmCzQgrcSCB8Zb/9zxP01FO2KJNf/ynMC
3mJwbBhSCDbluuTa2KoqYZ3rr0fwDjC30XTPk779/EOHRJexSkNxDPZIQYvp
L/coHHCjmVe5jtnUVG9uCeR0vxKeUq+JvBZxrzU6mATcuILgtkbbJkRiB+3i
JNRHmybuRNa2op6XL/a0SwQpXkmAIu4Hs+IQUp7PVja8nwyiHDzvwAJB3yQv
4qD9HJY6dphfuFQX7WkSSh+8KyzbrzYa0zAVZG7o24a+cgc4nR8/X7OaVibc
mATPAs4QZDCQ0XrU+JqCE92YYGuTIdjUVXoJE3xlfEIY4KE7V4sJ0YsBWXA/
67yZqC9cJIsDiNL2l38F7UNJG3/W4SWoJwPXGZIhhIWns7HunZX9bBBWdaC2
K9jivFpfDE9AQk5EkZ9xDCX/rew2FI9VE7ZQs16HHvfj7C2LOy3SVpP1d2ys
d1MlEKdgS45Sr48rb0QaO7VZ8ck4/Dftdg4w79odtEqNY+frPN7LU1sClKi5
wTB11K5AcaKIoM4UWcNwLmwsYUaNCas4aC0OmMxnaYUUjFLZmZG9qAcZU5u+
ejh+peYevO6IyJ0Xz1fdROQ2vj7LyIolHXC1AUrUQ8tP04ZprfY6D8duaoFA
fkzQ+3PO8Q7W4RUONNZ1fQXW/RtLwyLqaj982VYYaAwgcguSxho29W3IIqtf
o3K080Mar74hC93+K7wa0iVI0TRBwfVRT/ay4qD6ukziyyYxtUXb4PZBvgdJ
TwLsAoMISh482d7MEikDB1EUlVrWqbvoWRp3PLcp5njowUH8T2zJYYKBIw3I
YyTt9XlwEh4LryQZRaY+9SomAYPeV4Grw5ZCvxJfyUWeH7IKy4rJ+CNJif5D
gL7fQmN4IC2Jea87ZXSW7Oc7xhUP+VX63jp03TElWoskAb+/9i+pJqyOi1ff
vZv97Xi3+g6WLDonGWhijD1eR4r8tNFaHfyKvqo4g1WJEdKzfhFSDrgwf8Ji
cD4mkrU0O6juvazvDQh2gElqQAXz7SwkN5uiSsKNRj08Edm9STQ/1qoEM1SP
ltKegQdFIPo367te/rF9xPc5Fbolx87mKewrLzNMf9uyxMRKY82CiuaDREBe
pfFhbrR/xd44/4BEG7olEfGKSI0s0gVSTa39IMrROq3DcRB7Aj1qGVKcFThP
FUanfsrmJSPudS4b47o6pnqh6FRYE1LAl3llEvn92nMSNeIKQSREq0824hnq
y/Hip6wHpMLGLygSi3kvypQTf5iOCdGJzKAybGtdOLuEkQsY3tmB7FiA81aX
A/7cJ6RaqXY2UCc/njxeez60T0QgopEDYn3Srw0xWj8kk0Bum/8G58YCyabZ
wnUthxPpoezC2potZJP+09tKionNAs0L8LhlfvPmP8uVfP0Z2lwwpF7YCPSD
KJV7ylCNskhCoD5HHhuyUf9uUR+ppfaOaHhx47luoO/ujsPfylGBEr2mC23+
Uwuw34kxkZSlhF4JaqMoIqfsOpZPSM9vivUbfLmtXqQjmwvaqVE2z5zFm+7r
6k8iYulWm8LAiNy9gLZJbceLEbwxYBBFdGHJUJEOCYGQSaH8gDT2r9vGQOGh
aiGlF62jxslaWwhJBdv3HWSunWcSgQfhzfJjGiseGHFDv34FM6vsqyyXb03I
XQkKbxsXQY4xRnkMg6zFhKaQkXvQk2+BA9D19X6VAba5woYNg2jsbLBk9sIP
kfF6p/wlKVnG+1PyqkhBhek3qpoij/MMGMN0uQii+3akFeqpSMXrUd2BHnct
uNJa9OeUeHWC+Xa7kjKQKcPMF8T3qQqx7OJG6/AaFb6oB2L92IQ+DFyzxmP0
ewdiln6bnJayOkOURCOb8S0GEcEV6ZJW9G4uLGZta7K7hEXhvbC53/KgjDmy
wnu+uq1+PtGrPnhXP4k3ucuSPqb+drGJ1ATqX5nZA7I4fTB5cVtRZRGseyMX
JovINi1vLKFc1zLf3pphaxEdaC7D18Hm4zdkeCZZlEZGlelMc55NJTIEw+nL
hkiwZUDRK3MzfiqPK3ixVVKDTqAuBeJ/NTfz8AdLBgSy/GgRc1WfmreEUzyu
LZoaR6UD3bps+hkDiiBWMhwO1bmNz1enKnIuiS/S7eVh+OridPZ11d6Hx/rn
Zu6Yv58J+DN8INTNz4fArrDcs1kKILPH461+JhJTUa3Gsat6XZyZ54TNNOk3
TYNpBNthU4pL3xbqocliK+gBPuSQPsrbpQMxhAy0gaSFDTqB+JdOQ42yKr8u
p+dEb6p0C058gA7AWUUn5M0ncsERP3DpgM+gMLWH0oG0h+6BphtS+nmiNBea
eazKAn9YVo3//nqfKh3QhfpMDUtBO4/Ekoy3kL21TusDDxWC9BATH1Hs+WTl
Rt40ofEBE7dhD18bnRCRhO7XB/1XOTBR7zfjBmga1UENgxn5rQlSxUWT0kRh
ayx3QDT2B26qLrxNkceuop0FtSi9rIeP3dJk9Lz2mGjZzeFlTPaRb2hnLqJ4
rZ4pibZnxhJ8249uRup12n4vVrEq5NfK7kJ95Fq9n6RImsTTz81p9E5ExPRS
II9jrvSxNvnemNQwNmwApzF151yLjnhtjOCD6W6T/AZpW97VSau7jNcWtcs1
j2UFFqmKjwv5UGPe17SghR6BXjUJDBsHcJvfJe2dulu/vAT6Kbfwoc18xJIO
LZVFC2szXFVgUL09b7P6eGVz4B8Ilp8j3UYKrnNBrEwxuDJLecNPRWQQVYft
ccev3hiHiBLYF2JVKPKnZ8hm5XNs5e2cCiegmRRzjaQLT/q/Z68WBPTn66rH
GusMvp9osEb66fWvS61mPI8Uv5nvf9rNVVKwU1DvbSARyN0NFj0V5ZXK6b5H
cxFo3NCNZO9lu5yXotXyqG0QMkNRubMvCbcKy8IycufzaTbok80Vs2yDVDsm
mnTEItrC8XuoOwtZx7OHr2ZdIJUecu0ZZ2rdO3JPaRYxepUxmYuvdz0ZV+c8
z2DRp4dkHYsyhdWdRM37FrGwVkzbAr6+7bXxztzvD1wBKT8afsgZtQb80btX
nFJL9r/dlDaI4qhFAaHNqX3qJozCoV8yF/WhSumES2RcWPkUt/UssleyVRb1
FTku3sW5JQWvRhuhr0obA14T4fCPW+tkpOFz3BY4NW/BcJGOAC91qHqT/GT4
65Y+zbydyxF+vjJE+KjaooKeS3QZS4Uty2htVc7DvGZ5d7A3ETR8wPCbji4G
UgVMArs2R6vT6YthkIEfibo1nIVdcINFiN6P9si18UPdxKpPS+yZD17D+ype
y27jISerambzKqquIMhc3avyfVqFO+wBd4X1DBiSWws29gLMVXMBhVvIpcXj
mx47QbXriOQyMQcUhNLo094tQSp3vmE7HzHh6qxCkZ8+jF5AfloNZy7oBVlq
xhMJXNhxapJSX3tkk/YGwQOROT7EjkWGDGct2c6UmTwkMcZSSx348huW3Xpy
oJKWrNC1RvN31TK1pFnm5HasmxjAlBUzHKsDJZxnk+Gp6YnsWPRyB+MhZdmG
O3jT8ln6kZtiC44umKdNsL4UQJmfMF2zpkpvLsb2A6zRJurHXNxkMGCcViFG
bOsMkRBFD0zuK7c9A9lnwpDLYQqmNtMpbxQhYYsmu1B1xHkUlEv8OiInpc+d
h6HjxgBMFljIFg+aOyJ++9pHc1xYPCMqt3CzJ0Pb1SKlbGH1qSraPi7l8nG+
VSUrNHmLLYd+HblQfSAozC85ggKp/LN+F4nZb19dNAADeblya8dIfSW8+vY1
pQ6r4CNrN2QgVZIuoh8marQIHsxp8zHn7i/N9PkeyR+4LLrNwpXSuro+TS0M
cqPm14oebGS6Jcvd2KMrGynrUvDudmR0svUUlh3QzRRGT5u/XghPAkcd/v2z
VXcUIujpSgKv7zxRWb7Hm8rO+ZyYaDik3yV6h+ayazQcirFj4PsLWOYhqeNQ
c8q5UsvD4hVXpkVvw4RYw+klMRyiDLatMWadnockYzZeayaLBzfjC6OwKZhq
/iG+9nCeDo7kWdV4FL2hh7p6hGBwhMbUDQ4WBmSFTytKUQAunASExuOl8Ngg
m1QjNlS58tQEvDVGXXN7t+vz6IkGfmUFAqzI/4s2A1wJy6Ri4DeAwhvPWSDc
RpBkaG5GDagJLAHY+HUrvGln5g3l1a3mFZFP8w2BcUs7Oy2Opo9lZAcijehA
yizF3JN6+07ojiqYUjZbkFTleq+ZqVmGsMIDWWuTMaZBnCd/ciFEI28Kq/v/
RvwJ87lDwlfGsRXwwraBQpYRmJ5IWQsygz0ftR6nBtksimnWWk0gB+Bs6y9U
+rsP38CG72iNk3534wmI6yf4iXQGkPunbFK4KskDheWWVusKV4G0G7j5pSOk
qogqbgNchAuWq9x1rpIaMD18FXMLa6j4ZM3Ih7Ddu7nkd2OfmPkpqt5d8Phx
fEFZdsNOdXe6M+KA/uT3OCSnq27Jzc64G+HbY2E1/hyga6/DV2Mfv0JO7u8o
4xdCo4SgTe+rtjsX/V867ctjJYguJEjV2pWDb0foe2XYkREcByN5wB8Xjnwk
sjkfdVN9gHqWDmfWQAe81sst3C/IXYpww1rJRu97vL4j068nC689QctS5Jc0
4sGX8oFVOYi3h9Fp5rTpctTz+MGsbwRzEp24JY1Mcr4sxdV7ismhAdyz1ZhV
uBu0XYp9ID2VYHxHm2TqJ58z2n6+ipfjlyYOQMx2DgUDfz34fYrtkWNrYEup
TUysIm9vuui5ATLBZ7YGZoMLu4W4HPYVaCJsFhWXqnpsouGXRTaIwNfFwoJK
oKMVhuMr7jSlk8mBsktfr84bYhV7NAgiu+uMfnGpV5MoB0j7dS53z3oMk7ru
VtOb/t/0bsiudix15SdvLxSxi3JM43QlR5zPqR8G/3t7fnelZY/t5LSk/vIa
D4o6Cy4vn6qptdAs70Nof8XRNcO17oWE1+B3rnOOCMCTupJ3QAJOfickMBAD
hHX6maxH+xPUZ1S5T9RYg3PDYGpKfzs1BxX5K9xi9xid4N75IPWHyfd60hnC
+JM5yUCb2TNedPCsRbvDZpRsiahRlcc34W1E/PImXxLIQSePsZ/YgAb3/PRb
e9CugBPg+WwHVck2+ARolW8IGe7SVc898K+DkyJfJLNOWF/D5uYQBErlk2lk
R62vUFNQPzgBvdWmn2C53GnPjaqjn1Ze1us3+OwMMlvbsxN/ZfUf1x+fJJSc
jCFbZCbjjwk3YJ95s1tcQ3aQddwIkW7p4t9Fr8+krGRJOIFrO+WEUqXJqE+Q
YB9TYH0ms//u1/OgA01lRajTmgWi0lVWZhjMAJabdlLixF5l+DNy8uWig+y5
PXk4TVkslMnJuU9dMaGXRMFhNF6cV/zZgOOlJpoy3Rh/0J8FSSJBMroR3h/Z
PAWdiH6JOlfTy2YNf2NMlQM/nvywS7Lh2iA4ORLrZjVQ+ON9ia6u8mzPGfGq
1Jbo/HrSmFM3XglxdYLoD1r1LUTGyc247tAVt20kJgs3KjUmS3p66nWuAVJu
nNVNaSqlhgFy+zbrwPSsnB9dyDjZsPjYKex/YlPJQv/91jtP+qiFT+2Xybd9
AfNLnvn7/dfv+FUIaEMY0HsmUUDqqKeha70vNlJPIWiJE2jItBX/et5atDu1
xPA3ezVFEYBmtd457uieLKELJznBFFYz2iXJX8C5iwwxZxRGFz1obDTQBI0Q
QlI/yjF+y1uY1v7FZk/pmqZi2HR8a7WsNv89rigeo64Xo+UhQYMKba2gvj6e
fpidizHiYB3g8qUB/bV1cbreqcGecDJJ/lgiNhxRdaViW84JFMzBw1LU9JIm
pSkwfe9D2rtN76u51JIdDCGbbRZhRqv8feNRoB+d+Dj6JninzK8Bx0lfbDvU
/0xmeg19p5LzMKzX83DgjqvEo72hpEO3CqhOiDqpFGDwAYnK4rt/3Pq/QGpU
lqCBqNVoWBrNbtd6Htrt6+v8TWfqaPJmKtkYCnp0bXR+8qDP/muGVwUoy82j
IYgP+EQ82Mga+zlAROAZdJyIUjRrxoOpK/98oOrmxS26nvuAUxmzHQdVbBVf
hyD+G10NyrhzuCLrwiTtOaW6Sliv1K7WiDYVhVhNgGw6K6dkTqrwC/vvf+bW
rcn94Y0Qz7aW77glIiX3qH4V+1eRwCXDqPGWd92saOg4dP7dknwWf7PzZc90
aPYBZ1u6w1UBNEN8jxQ7L2TGkcD9VUiDAi9nmb/nzVqARjcrDsFqJFnOLZi5
izKBv7exsDok9wrG0KBC6Mm03JphRB2WVownMaB063im1ujmS0TpNhkOr5Gj
pyj0itljP1HShq+Mcqo4o9IJUdawtBIQ6hW+3ZLPj+83gowmTOcYsCQt9c3q
UjAuY4t9mHOIlrraCBzeGI18COGiZbPap1b33h1ZSQgq0YYt6KoZ1XWgSjcB
NiWcjbaGxxI0qfpjZqfHWf4weW0Errn7JVFnTTVoxOU4xmllZbAuUz6ntId9
wyUfs4VaYTe3oEFDgmS6D5S/c9UtIFqohsoR35/E0/Ou942/KjNjs9Y0Sy23
v9e3S15bnNqOVblCHElyuI1t0g5Y4r9NTEzqh/VAUazPwkoRlJa97L/I0oDs
htP0kqzHflgObDm1ccaUJ+HLikB/lIxCkyl+apMESIVGynnVkh5prrsEusS4
uDnigTkgnTfVgQkYgv7AocvIx80PAxrRG5cgL86dyUZJOUJeh82nU8nHu5KV
LrN5en1BE+QD21651BC1S/1rDORd9M/4+ovP1QBXbOvM8VUWAwZbUAdzqWN1
fix7NbKlr7ouJ8Y/Dzk5R2DHPVf01uprXp0hu0cJt3qvuH8W0GLgzvMAY5Qj
AYo4o7yYDSk51qoAx5xsb/E6U5JUK0w3R/Xg5D4M/OV1fw2rQvGwZZnGPkjl
0SiCJAV7Dy9rubbinqafLoTcjuswRW/olTJSiMfLrU4rMMxIXMl64gn9LTcO
t110sis4kTr1pSWeox57Eo9Feeh7yKlzrgTQmIMUbhhAMoldfM5NFzR2oeap
l5wjELm+JoQNpqg7zpsH8AwE5nYUiu5VLN0NbiKPUELdrD9ObCD8StOkEN/I
U8cfWplBxdW97zBqYGU7NwR1IEr9sVWCxg06qw6WboWn6z098VhoRbT0OFcS
AjtS9TNnDTppGy5ZG+mZHqBHii3ntkXrXjGr5qCZ7Fvw0AjJbd96v0tRmrKD
E5DNVITAbLY9EOY+Q5z5ntiAqlik/YDpAv76xYWre2tPSuIQ+AFCJPzIftBi
ip9X6ocmJRR4RV8OZcRCC68UNkc2p6aqxaMFV5yO68p91v6Sy68YYgsAWNe6
Y7+ANiwytXsWrEIZlSeBlPlbHl/95YQtB8cC8i0FRHQjzLyE1kYqtEbjCx9+
BXQLiwHp6swtpaVu8rTQ3zOwGz5iWTEg+wKw60isR2lf6MUHX6zUzmcVUmIM
MdnNpNeG6nezLBxzA3nhpbRv+C4oI+EL619XFDO/P2iI7GSk360j/9XT5900
B2neNR9ovSjoBF4rQh2G4viL+gH7Q7qqCUSqxc8zZJEGtbnmaYo9nU7KtM8m
wKkzp5GuzBE5gymNQJ2AmiR42+Qy9BpN5BZw8U1EiKo01HkOdKUzMdVStlHc
LJ2uFeuxaC9Twao5m3N7LBFElMLs6tKXtyrB4ZGQ0qFYba9YyQ6ud3rMZbr3
C4QgnYI1qqKzznUGZed8zpmnmEpGcDzzYlUqg/D4R+dZRrpL4JtjO/TI/cHL
jbSqkzRejTxV30UqnDtj8YwQvZUBehCuN9osfE9y+Z00dYHyrH0SZUUw9yMB
lpXdNfdX7dLLtrBty2BVaMCSlIWpcjfn0VdwDGCAbGDgTgRNhay3eVd0WMc+
uhba35gGrNolojQfge+vLrJdJkQSV6McVePhx4atzvYRDSWr0Z/9puASdvGQ
7w2FLCldj6WN14/oKusrVnQzzQ0/OdOYfHsQku1bq4+GcPlfE2jxSjiKWaZm
TkfdTs+HuNxfw5H720qWhQNZC0isd+gkIsqbtGJB+PnOP7LShgw48vNK8/BS
Zq2GgtcinIsOqysp1APLPk8FxPCiK18SYIUjjqoIb+rMnlv+/fugxeyeX7gd
XdXW7FJ13EIa13oH+DetGIpohtmYET3Xpy09GQVWbLT/n4j4kLgZGK1fqmc+
I1UNCV/6nDy6gg7g1dK9tKnGJhgTVDMBb9AH7Z8WgZ8k6m2BNclhbgOXH7+I
EZEThfeYqKixDbSleYJh/L0Ua6SwNQ0yns7v1xSxhoOqZlrI+8NTpk41HYde
U8e1D1dFTfQXkZKPeL7AOqq2GUg4zezo4X4cfE0tIEy9R9i/sbbO8mEKZH6H
ot8YKWtvv/YB+Wp7sMf5B1XVTAvDMZE1Sypuavr/EkjeMmovrWuIP58EXIyL
yvyxNH16QRtDqLMFbbuR3mq1t/Q9pPs+5EZUaCuOXjVCiucWpUT0q8qD7a65
nwbMEgm73AyoRZRl1Qg5UwA2DP9X+OjuADbCgQ90/p0/bqdESIc8fex6NY1D
g5eN2vTP6OlG4Al3GqLn3oDrz/us4z0G+YiMCAE2rq56jjCfM8t4RS7Zxis+
M2ayuBGy2m3+j2khC3RKVOyn9+LLk0Z4oabwJti0v5GfR2cvLEJO/sArBs5H
YFcVCTlcioFwQt7h4Yr99yuSw3u/w71eHp11b7n31wGlmMxZN4SO2NNY0Okm
3a36UdJaEGiEWNEAtIxRYlkiA4QEo8ZJKeZ4qrw1vwrTD8404zL6QSAecEMh
siDXCd0WSouepWtBo1XxX+Kk6MaYz9MxUBA5YKHwSUnTT5tncX1xdfMV05Ce
nt5l4VD/y5K2vniDIsPxvW2wkOV8myssL4DNmxowl6FgxCgDzCnXtgRKeD/T
3H1HUHNb+3rgEy7NXfxDowkCwgiMi0x3GQGnOyKAEbS8Hy3AcNN1YG+Taa81
bGrPwOBSEqZItCtvojEgGEaDfYNNMCJjmpUNLLpLQKU4n3H8SxqbrIVKde2G
fjT6bklEHl71jqpJa1LJDVUv7v5WJx7MhwGKY/qEXWT0A1XaUmw1GFi/x4jZ
np8HRSGfV4fLzAmfI+1PYX1CqIS1kviHB+fXjeFwcRWPIPqeSyJlp+XNpsg3
o5LHbz8B1GK08PEeI8SZnVsc93N0FX0mWhBKw9djQBMhujIxNmgqiGzTUKWQ
A5IsUDqZ782MApBvsb8kt3vwj3NeNEThrgk/QLankGk3wo9rnovYkxrHpGzs
/ftVzDev+RUcD0URTNZAJi7B9auT3/CUZwCBPJ9ZCTEhXLsh490nfH6U8NSB
XtupMZaqVx7Boblx7vLU36Skk1sCTTtotNaXlrmVsq1w/oRRkAIRg7gVCpV6
4jprR/i/4hrJgDmgzCsEgj17DExPX7VDziO62Vt3LrV72JpXtdj/Qv4ynTwX
0mPrkxD67fnSVEf4ifRW6KPlDveoYbLsc7egzIAeqsDWCCDXEC6axBI6HXgj
a7qUsqPDvOeJsPXjbZbi7TxeHNa9QQGi75//c9U564od+PMEefkEfEx2CDrs
9V5+xg6T08ulH/+G7MnnXNsx/ewYltA2zX1vGdQe574xcdlNSDrpV3bdlNzy
yYcQjnKwqBLfaoC/tRH5skTdJSJFJhDddfuYOVcvmSC8vlGF2jjW4zOHrJM2
CGBT+a3r/mXBYev/N6ylmBrT8qRr/7vqxXp9M4fFo8OP2KM3Kb6jzuGnOGZV
xDNDNaDc0KyOtvAYkhGaC5FQFrIYvErsJtf53UeSKqCrjamXQcvIjufazagh
Kvw4a3Fn2ryclv0yoVAffFAeeY9bYjOQBx/iG9RNcjkKxEtmiD0cbeyccm+G
GDASmQVQSV6h8AERoYf8cpemBXuQg+GyzTRIZfYOeGAdEI7ERcTB0AucRmXW
BU2a6OV2YL5sNb1mTqRpnAHjvYgZJfa17zwdBF34OJP6RnQqHMS7rM6bSOjE
0TaHQ97V9K8AD6n2YbafCGqgzzDziVNwVDL7vkHXRzC4b2HG0O6JqV88UG5J
aojzdEQdZnLmvUjqwrueEuMiSF+D0V+TM1ifopo4eRz+XJ9RqU1xf9YxX4B+
Rc8Bj84R5Crkup6D/w64wXIlPOydvltddl4SIXZDiCyArNnH6Xt6qaGvg8NR
ub0tj2IJecwIqUjA47TSH7a941y5svbGJ1uTSTBksat4/ke6PBGbIQ9yqBGB
ippvTeT89GnbtMaA47GKL8/l2xAtDsRJpNgA/tMjcZCRGmgROVQgFZjpr4no
QNfYe4JDiEmuAwWPEqkbJivTAe9USpNG6GfSyWZLcrwhmR/Sjmx6cYLMnaxZ
/eC6pIJYlQcOKviTz8Sh1HxU7ZQG1k3DTu3sCXtNlhsT5CfQGfoKonZ6L8Dm
QcUqdJ5Dd62AuLgbjtDNciR9sUZDufEc3nsCpVP9WJjZyh3c7liMk9CgN7mi
eoC1ge/+GVUAAAExQu63ZqBvJU/IY2qm8t0R1gEupCczcuz+bP8N/YGzgr+k
ZSKUslehzR84H1wwMU+SF3teRc4tZHdsx35xe/bvwf17fnxJ1l2AwcN8p3/R
IY4GHKXt+wXW+RyarIJhHW0RrWmk95JcdF5XLfUNsy/BdsvzsOQIxFr9HZO0
K+pHVeP/xbJU3G9ZVD6Dc0m1em0/78t0b7oMkNih3HGmYbEvHsVLc8beRFG7
muqI+Dm6iDft4dkXKIkcyedJ9Xmv68fziDJCpn/H7L6oXZTcMrdo+vvrM4+X
c6rTL02VL/yp3zWpiOQEjiVjTzruC3lgz+b7XBU7+4kZ/ssvbZJe1PhgHEoo
jJIdNU452ix18gVSiei0hV8qB27NvmYyWu36MRqr9B/vRBaCSk6g1iw6mK7F
pMuqEVzx3+B/0dORoBtxKqAcADPb2VHj4MmnXfIFD+e06X4/xxRTce8ja498
llVeIQuO0suX0+EyVdooootBZSjvFReQqduRPilkiyodOM8DydIez1NBopgP
CIsCtyOrgmTswcMGUy5TJb8uX6arLUoJ6ZVtcI3iOPWSEvP+OKL9C/lXkFGT
KmvJWjj2GaOjHqCx8gfbtKJS5A/Dv5qLkMsBIzPnZtUsGJsbtAzZFMsc1CSB
M51M/v1L+Y7yaXHxlMZmS/YKFshycQQq0b6aWKqfUaQsuvDaGAoF3QzLoTuT
jx3WwSJTbaXltY/R5NfjhF+lrFY3/yeDr2D2TxOOTNKDM4Gstndb4QDXuNnx
VeTyqoP4jFWkKKD09mmlkHOr20wRPc8PHFwCMvlAnp5a8dCz6z2KPWdLMjHO
/FLjhzGk/Itoe7Vx8vvaAZY6KudC497aqGq9dKAfOU6lLl+s8SLUbDhsIDjg
7sjn7mgRY4DV0CwA03zFVEGtJYbxFjwDQrPgkvldeu8ZQqRAU48rL1jxAOzY
1WQqLWay6CNFcRiFnhCrD1At3BqJYwh1QttORlaIbGLINUVweZkGCZ8QwBQX
CiiQaIQO1rhwBJIgPljnB9XlM40IODjAv8iJyzSe/EPq6Wd40tQyCsBjLtye
OruPF2FqtZpNbFNjMJ/V4q6QPqh/VanApYoAFgtvCH2B1K21/YiYWJFR6ptq
CX2Bbv642OxjcRBx2VETqy1mRoJepch+LHNpr4IUr8gsK0SZVUES+6VCJglj
Y3KpsQeRyvw6b6IU26qKiogXsSawVsW65ZhgSOWV4Ql7hmHTC/WytUCUFoX6
WLyjv2gaQn+UA6vW3viYHbXdfaSjwNaEgR45AUBib3mBfEMk5NBaf5LbfTpy
KqbNotm7W1ycF7Gf1EXa0k8tA3mMguQ+nVH68qLibEk0A+qd/3lEDgkVcrNs
2dEnXuERmf+jivjpsXU7b3H3ogv3UyW9CC70+L8/Ye5lgPQvQWUagh8C1+Mr
wVz59422Dm1moRhHvmXvKMgiqm+WX2pZr1vKMOzw9/9T3K51oPYbiPSpkaMQ
8l3iFA5/4v805jn9t99bQlg5mR5epv1cFB5/6xs6FMGS/W8m9mXBZeqqJryi
K5RrOTL5w7AZvXGIY2L5lIwiCrwZnL4fdMZgi9CO6Rey7HMemvZjyAxsKj5y
re2R/UdrzpxpLwSFSskkyH0DQH6fNkdBLovvA2YE+58aMXaRFuRYAeobqhDT
xdGR1vzDv00nhCl4sLl3XnhY+Buj2WM8JfWS1QgUm4XmtaW7GEQEdGDCZfQ5
dHp6dHtttkkkvUsd4jbr1AasuODtxe0VQWbbPuOKQe3EIiJKRMoD5fmGWhEz
gTe0gb4NmujE8jqZoQ93GCVrSVHdbTDpDd0fdw+ZFwNfD/6uHd01QpvZxFaT
xecDfqVNoocfT0T/cV1ngX4R/Zz9t7Ri90PGCkfoiV++zUTkBWWH5GsURpsP
5IDuM6+6N5zujDEhZY3sT7CUQVUgdiEFrSFdO+oLEQio2ENWZYkdRix8u52g
RiMUgvXG3XoMTOM549z/Tn2npuvYPDsSv30FoKTeFJ0EVKjkr0H/iy2vTUVi
INm0zypBFIgppn8lhi1CcdRwe1SKiitfNYcpt/98ieNwwc5Y06B357Wnsl3R
SAgqXu95fYk1NjcjKKXC8HIqrePe3GKeCHQ+MPQIHbUD0lAT0N5jCmD5JCT0
qP//KrjckhqE5HxEZSxdhj3zS7/AXYiCPpPnspgjpRpxjKoKy72vLm5Tb1ua
5bDJzhaK8xLwr2In7FXu1126SlgLz7P4jkX455XawQQS5l1BTgEJ0nrXeXz+
P/DAIlp7R1En3yEzESdgdGSBKi4mkJpISLfFIy+Qc0N8QgQ/KkzNzVsM0KvV
Gi5ablZANSLxFUZiO3AVC8Xzp/IqSrleeBcGiDUEtnuwKXuBkyE/QTGU5jhL
A8JbsVXLswrcdPbl6nWvF+ed0aom7hPQxhCZZ1ZMoUflqruktvy/w+Aiowk4
fHgcKLw40eRjIln+rJB2VobO0sb9RHf5EV/02WXZn9u+lGJXhj1KdrKLBs4+
bBHrn5ffdcpfpWdHLdhvq5LCZ4KXlIotyBLidGbqd5vIOvOZS1AQEeYK2ydn
dc3Eg4zF+4jE4WME6rJBkGr1U88XjWoRhlgITkWyjeNn+5PkvaCbd7p+4QCM
xflwjgfmtPlSmH7TNR+qZ3yVW+UwfhpYe23n4E1zgAB/l5sXhx8FDEF4zKL/
/OvmfAw/n1hfXzamgJO2ZPfyG+pJJYfIcHLFBCD5XT7oztAhcg7l4ZdyQdWi
trLLSHgnbTwIBgEnxgGz7tiMvPU6hOaYzaeJdcFDDDFpgy4ZH683Orrb7vaf
yL1MX6FhcPBoraiKtVT7W1X3bfmWBkZqj2LmjbgjjR68m5w9E/r4zlCZpBif
EI6ZqMkZINa/pWO+z3ZxTuZ6SzLGaSHGp0UeASlFpVqYytc2g7nTIcGX5+ED
Jbw6AI6GFRz81rm1wGwCRk+j9IWUdnwz/XpwkRhBE4JEWQ3FbM9lx8O/ktZg
DEN8A6NQdqOw/6D9yMrgqEHUW6RJ5UzA1YQuYnkOOlhN1xN/Brw7WuGEQIkE
OuNmWSLm6ym4XPXv241jzq2KFA8FNDfsNYbF+XoCE0H9AkgDnt1x4/auQ0oc
27mhVvVOsxR0XVZNSUxzK7U4QQBRUqOytLnJ2CRLj8oe/4CWqZqkQblwQudn
/YewJeX0YRdlrZYit+w4KCkNaDKrlZBdJrm7OeQ/9Ul7tQBuvNgvDEmAJmFX
Mlkk9QPLcK35R+YETGfYmeY+/mHqEKrgFZt6BR/p648RvfzsNHpSifIYdQgr
ZipLbtSZXUhLCZT9qLZWs+st/hDB6PWls+cOlSyl0cfRo1DtrQWdickVFF6b
ai1JMVOryDqaZxivrmvLcLe6hEL/SP43bGQYK2ta9r05FOBsdNlhbwtlZgxQ
yvfw1fM1E7rlW3/oEQaLshKL2yqw19oN8eO55wGaVuOJ2W1i+YRlLHhrYMmK
yhu0WBPZgpFzNVYXSMyrnquPhmreIUw3OO9iTPPiAUIxz/gbOEipOLZrQdt5
J932cVF1c9CLbxZKD2h7ZH8mLlDv+fUnK2xzCF7Js3X+FFGbzsxkXxsPG58U
asDvmdxBarixynF74yEo3Av/T40a3Wag8SNcLW7Zny97zG5LweBcO3q5PVG+
q8sKTPZSkG7NmB+xsXSfGpThyZiWh/XG9VpR63Rqgz/GTZjm99igzXf1+4kh
NZOYDa1qHeSCajMxtnEVAAGLJwlObfXIrF8Oa/ioX0fbQN10mkqyqsPmIuKa
ljJGRnX9MaRr1dfsilTBs+MOH8m/UZms8CujxdCuaGe3jzjX6LhNIqjrQ4SM
CpD9O+3nurf/53fdHYUYyKzRoyKOpH9gEd44dqIjuLNZracK8bU2m1ZgB395
aHtkarPV8z0FNZe257Gnwwl62BE8hi/Oq4wDfYtz27sKqwTMREzt7V8M33uO
dOXdtXDgA4icAPhnnOE62QoEKKMavn0Xe4dRywisVDQPIlWxpLYECa+nidhQ
x6T0bwJaSRzwL/BdROM3caMgOe1HyGSFc2/ttGVDmcQsbTakM0J8MV0edFVp
JexckXWFDvMw3Vz9YtVIy/rYzkAtSN49DBcelxWkbWgh+I38jSZ1rGURQeMh
AC4dM86F9d7eyE4A90NtqzmYgheQTB2sRNflH5LKT6of0Ebai82bxCY34DRj
F4qsGwaZrHIwzvPyuknttdi17q7Z0jnH5GN1H3SBALYCUaXTDk+YKdR+7nj8
Dpp1K5ubleRo8JTs2BKlTf2f2VeO07UvPkTR5m/w7iPXPswNAhzHno9jIEEQ
Uf4qD4PGrrwb64R5U3BcFtKsvbKMhjeiGdLkcu6xS+mO7RGs+NHaNkvn2Box
+PA+6T89sVO9B01Y+pWCTDq1mbqk59rknVcvyxc6u1xxSKz3c1Sy7t10pZxF
nFdLxVooljWOcv36ihHGvZAXaHzPyAZfuwqfaI9N0c1cPy3GEUJKG2c8Z7gJ
xxnpUpMAOPGkcA2AdLiUeXetROLlGYmYgHk/77V1eiMEXkh1v0u/VkO0uP4i
EGBkno9Kfqz7xZzFb51nNWPfhgdmn/2qoXmgEEn9dXHxeRqjcnC5g9x5+Zz6
SJiYS0I6bk4ALFlxFjI1U7pm7HrQ+HnMi2XW6Ibzq82GYnwmcBB3hWgIuZpn
aw6r3wVmYlFF3tnjaEqAiONgfKkyu2i/84iAFuDFk/sEN72B2WLvIsGNTVEo
W7hEKSJcdVlqu8YSZx7LDMSFklmR+jQ+Q6ADhamQS7vxvEXlHYujcnPzTR7i
a31MwCzOcib9RHyVbHrJGIYtTBBf0G6SbSZrm+ZAmN5WvH5L05lwCnHdcTL7
jzWB56CeiKnKCAfy6BPtml2VgTTccnASpULtDyEd8W0qAdM4c8XQf7DCQKWs
sBCqVsYNEF/Q6NQItRtFpV24Onws1yujVw6xsz/yJ1nsjAPnbcVdS+FtUMLZ
r/6hD32ojnJnKivS6Gy20UAXOoEiuR2cvxM6kHy/1k9Q6IoiwhHMn0F3qYJa
qSAo2itOBu2XqINexSyNXHo2GMqiOEr0qBQ2yXw+/MouXZ0DiaSwRROo9bZL
qyXOfrhSdUEbuvPGxDuCPI2Xx7MGmiKbYdzDKOlq902sbX4MUDJTJKho2NzL
yb+/9LBNIytXrN884XCSR4RCmCi6H6Cfikkm1Dch+z0liiALtOVxI6ssjc4G
KxDKQvnZzF6M3ocjW9GkEuuI4kpySxfMQicmX5G1L7DAlbGk/S1yJmgKFdMn
W0sqyBiG2hk6ax/CCH6M7Bnm8ZbyaHoNCPq86e9P4UCPLxudiXdAezqO7tr+
GjAvxiZBErrawYl/MgexwXTxWvK1SFrGt/QsXO1lUnGJkiVRCvXfyZaWiUL2
o6iXI2ofr/jPCI3NRslbe06+DKrkEgWHa/xD59SyKwkeUEzo4/wsZ9R+3ENm
0hQLGkTr2HsmnyYU18NNPUWG0iqDZ84heCpwLWbu3agvJfCY/35yVFiCXt8F
0SPNRs4VO0G1uJ+CUQar9IjbhNdPqpF7S2ZwilYQN4Bf2GmQU/E9EyL/eiAd
svdROulUyaSSWXBBB3wvZjt0vSLr7IMQB3ejM8fyL4Xw1mKTHYPiI+2+7/2O
1C2qhsbIYwllphV/mQV4tHyXNVvstBt0Beg/VS+Ah/elcvHX70q/sqa/jtc=

`pragma protect end_protected
