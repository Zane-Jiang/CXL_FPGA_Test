// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oycLspEz5kHzbhA2Z8pCOS3aFZzzjqJL9+EsQRj04E5h19Hyxwgu3kTJiNbH
GvGYOJ8rXi7y4O2Y2mLLTlT199xYbgk8ZsKjUwCAibbS80E/ZESG5XEydbGX
tdiNYeJR4x1D3ZiBM5UwBN/HU65zZGtSh13KBQ7e/oZ+cAB69SKtAAbQz2a6
ntMy6xQumiSyMVBwWYZKggdBAFApFmxgkH2ug+7/DoR3yJgXY5oJj3Te0rTl
WPTeXqo3YiyGyFor2kpzq92s2TUNmHxiE1IZcOK2qNmoDy2LOjPVZBizOgrg
gEMb16oH574ZArLAtz1Nr49kWq7RTYWCF4SupUSO4A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gWCe2OTRrTDTaIHhHcrcLKj1fy5tk4uOb59aSrGsea1Wr7srX0H4WWh1N3XP
J/0SQWqOhUBEIkwhF/TU9qf39sej9PHonNGFsozhYDN0yOGku6gRVEXnddj+
3OmgRDkLcVU+MOukgUQR78ZpelrF3nHn/l3mEk+jesNs7EzaCq40KzTHHk6T
lucI2nOBu8gIA9NYtU1g7LJcPVI6NDyB0hmPumci8SuLAUa1TuJs3RVIsZEX
w25FFZCIFDWbkLdGIFnYP2O3RkNGjM5ei4ncXvOpffxkeT3z2y1t35nx6uwM
UOQ04u32HA1rg8cS5XfiRUdI0WoMMKyS8dCIu7Q7QQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KDI4ODKzqco1haX/B6HOIwSm8WeC1XHKPaweAjgW1vELdztrqCjHXsJxdxct
lw3sTZzjy3bi2LQ5Ojelj7x0MrBq7Ev/GKfe8kz1VyDgoY90DmUYzQb77i9n
X78bzagyl6gQRkSqgM3QKcvvy9C34PSetR+aShNMq/6YEkeHh6/NaPXaU3DM
rQrz17sge1MaXK5L+xRNWq87+8qMcoQUcmooH6YLV0byigzWWZ7gHthGaNgD
8RlxsH5ZdTIq5bMgDIJOhWCkg+LKfLvhwhAjWGin0qqFT2lXO5LiPtwSHvw2
hj6NbdmTbAejkrO2vzWViN9oSrIWe/CK+tIPn08CUw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PEvI+UxVcexjlX49HmxIqdBME/jVoXxb5W9P1bv0nxkRRt/YhHt2LJexE/Y7
Bnwu293EXWx2FTRHJYcK9Dds+JIhIt9GxRpX5TXMBRDo3Az4hvqLwdeWdUzH
QPf0GM4Em672QhvCv0txwvvT1p3JxskpTALMvJ/wHIFMnYSaEVQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
BrCSi7q5l/9c0Euye0aVI1T0rl5hUgZF6Dlh32PWqokx5RrYiS5ss8CxWoqW
/+A83fF8DAh+kn9dwLXwzkOXuEachcvcGpTNVhsuG+x3MUrkCXl9+y8jiUQy
fqgJAHmE87qE9OES/ewKOKkcSZXoNdu/V353G5ojy4cd1KouZa/kfGTO7G9z
SlsRS74vfOneHS0czLfWEEvLftSq0YDf2FkMJC79JPalROhILUNw+UA6wMrg
d2ru/iQhIXTUgApclw/5GhK/+2usEMSYC5a2X0ySBOVbO8HlHv/OrBUL89d8
1NLg7rdREYZ+RL/MQj/QzT+Up9+DCmju6QGFO6KWi3KYZQK3GtWaNnLuIhyl
IE8vCtFn2pC3RUg57sGeRQdOJj6+jk5rtgSpVIcXhpol/I8MQVHwScBC5Es6
b+JDJRR1X7+7xo5AO4fWH1LoJh1qgVamYeTg3U29JjrF0b53deu+a1sSvmGC
tpZRTwo33SdAEdDC5ObmaRwI0KIzNY7H


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
meUupbgvD08GBhKw4Yffn+qVTO6nZ3xs037iJyin1AhuibbjtmFsUpzTuuR7
ABxZ2j7zVjjXFjlyWXt3SzP3X2LOi6OlxM5cSe7I7TOdUS3tSy4Kr06lOWfk
Lb+k5LOCYmBziyIqeEKeFc6+hfn6dBQZVj8wdVbOSNGQ0iGvAnQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D929+vyqU+myJ8QwXRNEIeAAe7/SJNB1kMX47wt4RK7Ee/osKCgoHgvtSWdQ
vQcJRL59RZk85aXCAORFFnUEfmsPHW2wbtCKeGuscVai9MCkNc3cH9cSwRmH
xLefKKygOP7YLDPUfL2tAEKiNBeG91D6K4lB/OGjNftMrWMVWKs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15568)
`pragma protect data_block
zo5BjpcpdRplsI+9t8Gf4YqVTRUEzwTIxVOb3Q/UWOe8vsx9u7CQdG1GzKVI
/rNdUkszIjvW4vwMxT0l0btIopcUQRPkvh/nuJVXRV2YhaRaCI7X8qanPo3q
WXOuJDgvKx9+RSPdpaXjo9R8QQ31o7oKmsEUFRa/zIlipreiIcBVKoWEg6nN
lkwaEDRmrRPT4z1meReRFrQGYY/vwFLpwbVKKzD0W5KeP8ZtNxPf+2D7lei2
LtYh4c96dQJrARHbempejYkmc8UJ33lNgKS+S169Z+Zo92EJacoBbKKOcTiX
xe1gMd220CFTttKcePVX3zHETKpH92Tz65TA5qHZ4RJJRX9HdhLbzxLbW5J1
AVsvWfbOXT6moKO4TJFZwNROPnDrYLU3+SuK/Lzl26vwMC/PV7vujDKPTghm
S3OCda2c91PMUV6LySjvCGwP8eHi/6hnvp6WvYhyNy3gKk/gHfofmVesORM+
WGrhqb63zjJ2cJoRRoHEG4nkUiBfu4pvDl2QWOj3qfAsI8lsCjpqpBcFK6wC
LrNZrj+zWqy+i57EP5wvDWqt1FSocLf6vbHY8GKAnXEUvBdTtCaAN71wvl48
vRuzndndrLxLWONrzEUiskxOgLCDXBb7Eyu0M7VVrPTX2rvdj30RsqgdIZCf
S7MPEhVqJLGIKX5Uh8h63mHu8cjPl+E4Lq9PUFLCOdxSagoTIC20Yk/laVM7
Nm1evLgIaiIdMrPJm7mnFYv0TgIifWPocrzIrQ5SxQwg4dUpRDv0Y5S5Og+C
DbuJY2DzsU70dcsiw0xoYU9z/8OgsRa4OvF695Y9tqUzfeC8cejjdKDruIL5
lzumQ0wGAgGOMgWq7JZi9GHzG4RoJkW5ewRsgK40bVqO2hgBzrolzvzWI+cL
df+7G1ZuSFWPNOwqVz8zcu6P6CldOHXesX30nrD8xQJNMiuGD6ts9OH/WY9l
dspaNxVkfKg/TqTsXnaWGnCqbhSqL5bwVDcGnEwsBu9ZP5XkkKj7u5Za7zQD
wVdZvwLgASXMMM+DMxD6R6Rgzu0VxLF6iRPc4/OBDQP+VH+1UOoI0w3we4wC
OvrzWnq+NcwkjblO9vwPi8Gl1xmys+Gv9Fa6dYu0YSHywgU29ba2eokmDFzF
tVNZ3cb/SgCgbd597HJTgLosAomejOQQmGC54SlmrdQ9WgmqsH5mhHj1sRoT
Ktm5+0YAMA71To8Osj6MmFzc933eT1UhEzHoly8BFZc9qpXJN7TXHIpq2AXH
E3gFq/aZdJj8ZZHZPjrY6lnRnO4PinigT2+Xoyxod7Vl+3VgMAGs79ICaMV1
26QdMFaQFIghg5cTkp2fncxReHhifeYt/xibPwmRYdqed7ce57tmJYINro4v
6ZMNWvQlXp26ffbP0OloqPKg82IAzA0gZ1aiuCv4ICBM/wnVGRbnOKRyyU/Q
+ZPm4mtKJOq0JG145zlx5JU72hGSi68ryOcoLsOSdz+Dx+UrwdqN77ahZ5Vl
2VEBz1cFv2q8z/oSCmhe6gL002WRZI6ht8p4zYxXLeREIWX3aErtXIkuX2Wu
qK6LQaZceJHE9jPSZ9tri0Xyw7QSXhb4dv1R4IuUFV8XRE0p7SkGQCDzhsjL
5AzlS+HhrUOBOcsz6DfzlDiUqOWkG3w6/I2+kat8HeYMZCA1EoHqOLVdw/vU
6d3+Mwxvyyfp3+7EVS0sUXD8OUOF0Cf8ETflTU3bf/M067CDU5rG+hyTTrAj
9QXPg8qVnlKAaEzb7nKjhx+hsB6/SE6hlIC2nv+GPBgtKc40ojVI+EpFo26I
R09N13mapxh7X3a255aID5y7OjkF3t00+Lzp1q1Mfa5Ng2qD99tIPtBqv4Pt
pQtujiFnlVez/U/Wx6LvzibMFvbvuYSKS+W1+/U0eHiV1jiWhb0JgTmdaHfI
eh66TVZfkNCGOc36CbtJ0zMyHu1UXZxG5gix2tzEYl44IO3+8SHhO1ktm9kj
U396DTb0jgPFHQLaWJCPNYvG4wsqAYConnHmVc6CM3J/qz/UxwtpHCRlR788
A9owAA1GLEdSglDGTU3yjK72dPQHnIAiQ2yByDsxwAboiMfanGHxBI0pw+4H
VlEShRcvgJYERbt61GGN6mClHNZ7aotewivy7VlSRWKTbp6yCLSoIEvzdd7R
ZCMfCWiNKsjhiyY701U5ddQ/zc9l78udlW5Ty1NdHt8uq1QeOITQOiL7sJwX
BR0lY6yuIomiUIHkBpjNM31y9cYpRtychqogJSnQE0Gso84yY44RiPTrWNnT
ixy5ROx1uRfrrrAZJLa867WPCNRBPsHtnw1dVKt52MyH4stAIhsf4p+93TCB
Lqi5CUkVkKkobBJH+U91fuSvroGWmqS1kaIdaYTMHKVF1wWUqD3oqJQhdcIw
qB+shGqdnfjO+MPeDPlNvCaH9MuVAYn/QTWCNhF8BiPXQAVvA7ufne79/ZSB
cxaboqSm9cKUckgiFTsHZTHXuvB9SspdjjeMGF7J26/sDvjVh4Of7n91VG3m
gO90kIu3FcGnW4/MqFFIIS3Xau71ddbhWoJztgNZ4glAes6N1QHjxYtmp0B9
tRPazamHDvU/FV6j7g3K9d5RUJmq4UzFcXJayxhk+5MSCKrQXSwPZLh1tNXw
dXc75FbTRU3CDgnxsNVZIZu2XxffeJrmySloDnalMt4VA3TVlZqo7GdoIGS2
JcfJGDqPfJlo2pP0sgVROblMKdAxHJuq9x39IxFGDYkf6ozyV0Efop5g5VTo
uqZJWKROE+EVB4CoJ2NvTYkZCBMRR/T4IHnt+9Vx1/xaJzw0YxPKntcsqOfW
BPTo6QIJ+eithmOfErQgpaXw21+fsvCqKI8BRK7fMaTUeNQkorkhb5Z2usUr
hgdUDMM5Ym0MtSvC4ijGc6SitjfftPpsxFl0DvMrMmnrVqcVdcAJ0TT7cDYr
QODGf2oP3Vq5yNlhJbYBFefRo7lDfyJpORsLq+VGOWcCMT0UVgiXrsYXEvkz
7NEdK2c3uc8S15Y/FfJ9q2Ws0HIcVXlb6stpx0kRNkso0AGEqJ3Q/ypRkAYU
mkV2YbBJrAgHw5b/Q202r+pu1sTSEvP55X6nR3KLQJA3ZUsJ2gPr6CETrwu7
TvWodGSUu9sRTJnIh3IKsMuX58+aOop546DIxOnUjHJJONteLek73earlNMS
R7gQ7zbYCUmuZmQd04xNHcF1D6Fs8ixmLQr2PG3kRAbhMapBDU63hMRirjOR
iLtQWdWWMpQHYPI54hcXxiiZAZVukQ7wgGx1+ehB3yssdZS36xHwRpQrjBSF
+WlfeEIhnYj1ZIZGqfnBp2As+q0g75Feu/hyel24yGONvPEzvYRdP05bzkbz
x2VxEE5FWFrT9rFL6vOQTgHDM2ZCuqqvmJjKd36TYiuhV0q4xi6lqieIUeVz
um7FNszTK8cEAGOakyxDd9W3Ulxvh1y72tTlD6ojZ/N0I2xFVxjItTU0lLNS
a9LBfVfc/k/S7WNDFQAkXxa1dtzC3AR0dNdf0WQAjMQowMYU9QkdqfWbvsNO
aTMKUw+LRuep0Qb0MZE1GiIUYpBElPJ3bNkZEBoEg4ADscd7axPp/BIiKQEz
YK4EZxrLKcZSxe6Zg/jZS8ABYCBEFnpaxAQsERxLXmgJdkKQ1soplxifB3kE
P6jUDLyKQxyZpzZU4iGoiLEWwagzERpZ5eHXrmOniI36NnXLwbzkLIY/fSMS
lTDHSJm1p+GyjRixfYAiaoY+ez6tU4A4W56kO+Ww9wxDfTh6NxBUVxIIfw5k
rz5nY7UUxUxe8ImvfhUGahbQ5aSDUmtsZ4Cuxt0SeUJ+s7yRa/iYOXE1FrgA
gV48Yd2QiXHrgzr1agvgGk0b5XShziVq+gK18eZuna8xuOU3g5s96Oc0bj1c
ouxStZATEBrQTkHgtD27UbBQrSlr4oUeUHlfmGGRgGUwViV8uZsKV+/nagDG
6y4U3mIZmJtZY0OawW6Do3VGVF6+/hBz6SxAK5CfGGSx5WRc7sLNvUsddTWD
WjAnP2qdbeCE27u47dJ0KHqKGj2RMdqe0C6FelB4y/xnOjBhCIYDSb12O6EH
Sw8IYLW9RLLzsr9gGuy/jglSlrbEFwyYXeP7RyP1msITvMpsM2cvBRCA6Nmc
iTXpwsFbfqNZu3RLOfmTf9D92isRFa+PpnxbFj+TlIylHoXARGMHMFTNjFlH
q9mvOLF698my/xSlvFViID2qPScBYW12MtCsaYF+nPoYRKHAFxmCbuXWcNyw
wGaIMpGI0D+szGMBsFvy72IaN5olYI4lVOr1MLtWynDnxl7mGx8J5BHvh2Yu
t1tWyH7aIyaXgGVL2I734Wqs/B4muD3FRm/gGjuT02piugk/Ghr4so3ltLBD
J/epbmO3UL3QvyHxiP9w2VF14FVlpHp8AlRkIYy27mOLCSkiRDDvWFft19l4
63Bg91BrV3MvVwACd1Ebfx6lzRgk76oOP20k+3Ui7XRmH0d/tncv1ltoe7oG
cgrRZPf/QXFVstSuHFuyE/uIQkYU/c0PCgmzE4ez5quYBGcC9Vs+Dt0xXd8Q
+ReJUXzpwdXUD2jopCAZNsUNgSBASVrlzy7yK230knuqhxozw49u/gdoVZn+
bYyXUTVtDZavGUoo1YZvQwDl2wR6eBmWKffpdVLz3twKorogi6b22AibHoOQ
sZG+R3hRxml7oQ5VerNtUyNvrHtYdf3voWHD38WYoK/CIERhLFb1ozmcysOI
rNsq/kARiRRfBz7JO62RMjbf5wm0L6va/EMaARGrLxd+4ziOt22k9cq1yjby
bZ0AlM5iwHg7S7WaLb9+KmSo8ix83VPoVgaPB6b/ba3pRabnHPDa0DzhKomj
DB8JbIutxoUpY5tzsgkvtKwsHtTXjKZAjXUbIWvFaRT3n+x75bqb/iI7bf7i
1Iw7nRzPPjB8vPTGCf6MOWcs5Q3EZnIaKSQlXseCbvRGtQGcNlCIsTliDrcg
WnEVVkJ1RbdYyDoFJtEpO9aTKBDw061wEdNAxn7ky35sDXdsT4x2/IbKBKZS
vB0X4j4PWhfeEaMa6YMRUfLMkZt/nmotDhfmizDVol2fHQajgJx4sddfc3Nf
e/BIuNEcJUq52Wa5Da3BIAitKioSKP7hJ+IktEVEmXQ2MzAJDTf2YlJotZUv
y/gc+QgRNqtkcXCepqOkKsu6bbhMqtJi1fg1TC1WKQmIh/aG6GGkqhRe2t/U
2Ysaj/aOwh4zGFAr81qi/kMUZ3tCY8lDaNnuzjPAZbjr7rI1GVd2Qyc7mU6h
eKGOJ4vxBKg15H2y472bSbQCZGT3lFqC4y6Qcv5NPHJyp2p7IX7A6syGUbjP
VJsUoYCpJC1nQJIlyWKKTw2ajmVA3bU8ZWApVuymMjPyOsEyekeOwhvPlfi3
dBchb+pqnShfKkRmmlr7xJG6gBwRG3nX4LFCsn2dmpvkUq+02uqADPmXnmF9
1vnxE4PoHgkMWg3WpshNTH8VytHbcYmGwdoZmYvRSaiYPSjpCJXTh9nF4HkH
2ZU29gu1YhF6euO0zVjfmfpEJWPVjYDPbOGSTGkAMm3fHfr8UaW4PNPvedVB
ztK7Wqgm9PXk1OujivYVUCzGCKwJ6XIvZkOQ1hxOraGpoF68kphP3qXMAYiN
PCETUmd0ly9l96HoBk2CjgrabVWN+9o2sWNSOdiAggtrGGJD7Z9CHLz9y3sl
axy6NmIxg+bbh37S5Fu3gFd7gpJeF7+Rdg2HFkk9mCbSyn+LTcgxlmSIS6Y3
lvM+KML/zakZm+kv5Mv63jeHTlUoHZaeVSjyEd43YMNA7XKFn2uPKSitw9tI
dx/kXqZLa6ihuO/0SsygqILZ5gsmAHY+KFyLXQcvmCCManJFAlzod3LGjrrb
IQ9YqPoiWjs2DtLPpqzqHvBvTzCuKxhmQYPpnTUQc/2VbUVewrGFEt0cUnu2
P2bkGmhnPjux1nnSOskY+8zJ5GVWnM27jvtlkfM/PJ1OnxDFD0NCp2yi+n+x
st+4c+3gxmt0ExhIX2HoohUQjhSA4/VKI8EtdhhWiicQuC40xH86qatbURiZ
E7Xs8jvzvjIK61dCgVD9IabBk3URbiJG49xdogcN4t1+gC/lLReeHEK+acNm
r7J39eJdWZ0fJJJrZ0ITqzUoOXegZwuLBOI56DO23ARB2c2zsH+FrCv2vJ88
TUz1ruVPMU2myJZMPgVKXfVQlgwCOrIT9euJ0OGk6FTrO6lTnXKaZM3k1Gmp
6OgW6v5b/srG3873BqxwbRW5LIvraBf9BqLwRThLqJjtzhLpUh0VJakdrpMO
yW8fXzqAiM2oEFOILeEx7IM5jFCvVxas3kNdLLkSHDchdnxvGCmTleh79BWL
C85Xp0pUyOpfWIEzgxBIHebF1u3u/a/S0BQw2m/O9ajQZhGQ9/FMSWjFCgnZ
y6D6cPwcw2omRnpiBha0aSPoe74abCSK8KmFK+SnGw4FlAofXBwLycwIiU4W
eogr5Vd/3/XyfXYOv7QUm9MNo34w/sBWX9BqmB8eUa9YGVnc/Og+GmrTm7I0
Ummbf3VNB0qlWIKYG9QypZbzumqvrwsJuEvXAavMyrsagI/+F2SOYvh8NAUZ
z4cThXs2lvd12bZGmgNXxv4xFvPbfENLZSnEbpCTFTuw5jqDDSxJEOgvUT+x
V1UO3xZVxaFAACH27YlaIK5Z7QZI+LmcXLP3q85zhc/vMB6f7UNfPjwEjVp5
fwDAufcbIATvoi6JGp9D74HICntGoOuOOF9+/gTb77m+i3IJ33eEeU204+qZ
jg3qpOwPZ4fyQ2R/m4vZP7D75EAPfRR8dhOKqZtRc1bTrFNRylMTJP0kFWlx
5eY5VafKZdTMwasq5uc2WU5mGxPOtpviIsvblXnEqDwXYKWwDemJj/qC4ah+
VB/JXLQXLHnr+7xOjYW+AURSqRxvpeyQA7cyPZgWw0F6plpBh6Ne6icAXnAq
dBTVcPMKzXw41WSPNv3kdLDdZ919xNui4SxRhf4raMw42lHSpu7NPuUdvZ/H
GuW8YgfFqKegepAc2tUKhf0FFXVALE8/853wnJTSGqm0fBTs60jJx83W86Qy
JkgCvLoq+F3LdDAf3QsKpYrbhu/7S1zNFc2uETCMi9XHrlYyX42f0cNv1QQT
4Yapa3/TsJndIut/qTQPtgX++Zr8sNoRNA1c1sUR5iHSoSKq6xXQu8RHCf/a
mzn+7t9ikeJ0/Mi7ZGkcf529cxHSod8ZBFHHcQCjPlQdW85a9KnqPiwWY99H
o2tMNDumNSZUoplMh5cpiDKL2G+dueiFw27aYWKxBDb8E7gmqgZmwZrkBhEb
P8iiuFSxSRC3XutpqPUuhmGoy79CU4I4YfbfUw2PzKJyyS98dYT0OT0maxVp
E9NU0gMIHbKd8pdrSWk8JLKTPpEMq7S4b5PxePZGQKzAqs1X72B/ZmBgvqtw
qyfphCvnAwEBXO1cFydz3iIDJI5Olq8Y3U0/VPErssqZG2wS/aTv3wh9zmCe
J5xEnaUSIbL2hWifC2/XEKDlUHkmgdOBh25a3zlGCrkav3OrpR33E0sNv5m5
P3UIVBzUUlvfYpFDDF/ZQcRTnCu5rFT42MDC7yn5v8vsdymjyDl/rj5a6j7S
yjDOBnjhcwAuug5yofvuWgR2XHw30WY3b7tOcYqZmRvWnJ/Cv03Ee7Tn+6nN
8dtnnw2zJw+/gf/LIAYcZLFZ2EutxktCmosZC5ZnGGQCcDjh40H5Dtlz4FGO
aKOZuqo/7jhz0o14dXzVYIXdx1uTMPvNuI4h4LwmCOA0es0Gn9VLWJj9lQIk
HySoHLc7WAAaBbgZMC3HKbmw/uqnkkHnEwkPimApDtjJe2Sakb6wwEkanhSe
0CbA56mYR1pjX60fcRUrq7ZCMUX+H1FqTiH/h6wcVzbYQ2j4/P4/3UPwEO48
BBO4MrcgTjpdMG2ZBF9iATkBC0n+T4yA8flMjc4xEv/RjjzJ+gfIu0F/nEZ3
F3L9JsR6npt92xM7J9Xk/HChZO+Txh9RYH1kW1Oivd44tnIuv+DDYqk/sfLj
DG6LFnIYnql5jxQ6oyilbQmaYBYMLAyC/BcrUicCE6khdkTr6ZnhzWa+ykzZ
uku4QxjNQ1OBiOWgEWFFAdwMAyt7GSP3lp4UwnTYcVmpTryiSLe8B4Ua5IEx
RoHpAVkmiZbLbLyhLErT91jSKmHR+f+Ax5vJ54Rvw/hHgPJBVava6pcC/UHe
nAqdEYbTD0XtxqLsF6K/Eh5OK0g16sqPjFTzoTbK9Ocz2kZ/NYgc3TK83Bmb
3haYg/FJpJw8ck54f/V7Z5PMbjkRoQR+aACJEUHGe3Q2Gqh0HCrtUWN/wxOj
0Z0WME2hehQ/HCJjpJIdXdr+535CaadX2EXUUdhp3TYQfNSUiZayvHcVBzWM
R9RXhiSIOJ56gz26/WgjJnd4oaAGLFMKHqkZ9TAbWjrPS516QyCcWJy9YajO
04spvd8JJrWyd1F1n6Yg2KDVJXRXMeiGkuICtrqVnooaOal89PVSgRKj9jMF
6kaz8GNgOBsYuAjYfB4Oh+q5v5I81XMtUODgPfSd6mdtQ5SpwTFpxOZ5XKtt
r8fSJHR6lWkm6DU9PhlnZrIk6yG8aNzVKc2JrmX5AU9gS4BepJJKICLg9Koh
DAPORdE2p8rO7oMX+AWybOZc9itcifM4AYPr9Qe12ruOKt16P6W7S67EcVRm
Y4q/30IjRzs17H4IDcp356UnHHf9YtJnSk10e9ST2hsAdEs/pWRAPblPgR2c
w0UdaDX495JECpaQ7sV9I5NAAeovsYR8j8VF4x7wxIN0ZoJ2IT7OlaA7YInL
cCFQnnrK3k6fG3uA4yhFBuXCZBI9fh9QusORk33TN3iOtylVmQ8+vAIFyP5K
PiNgHp6gMx+FyN86hexeyXAAQSLKeQXQW4YUEit8l01VH5CRkaATnBPyROSi
LPdAC9u/j7d8iWD1u+aUChTP59Sey4Vf4XVot5AlgIOPAaJYziII94KPdLfG
0iwSN+OT4MR9v86s5V1MFBuEIOkvwdLCXVQ+iwXk7Ylsv73MOhoTfwAmfzsN
ifjWYNQb1nRZej3xV/cCJXnR/iJ5sBwNn+wx+IY3VzmM/jwm/xDHfBV/DgZU
BzglzinWVR81fqR4e4SsGDw15nyTZnchyTxWuMl0rD3QB4snCXTvFeFOjXJT
J6C0c0LSpEnkyBnCFHvoXstgk0WG2xXQS+WeoYoy8tIhNamLQiEVcZNTDa9C
dZEbdkjqqTVZJerKIM0aOeE8+MY+38RilQqvMxJS20JnBBaC69qbQB/4nPfQ
7vQ+33cVXEcHC98VjIDyFghHdSrU2k76Snv+4+8EuOH4PvFAgpOdSXcOou4I
HCWb3yiU1yb1Uc4XOCAeKsfLwMOdsi3YCsQnXR8dqVwB4i/wR8GRFdB8sEQV
RY+BNa49t7ZueqwWnrzJglvuBHtc9rYn4lyF9VjnhlvpJa62BZ0BbXbkriX+
yUgiaOQ7uxfCzXxBnAhxdoQnaStewWB8V2LNO59/ynfaW6qdWQtgikpXDDIB
Ud+j48usf/fJ3TQ4cVPesjVo5sxeja7d9WbMypFi4JLKpdlpKleCoEgqGGpv
0rfQ5fLb5B6m2QaXwlLxochDz1Rw2HiQ3zHcI7kv2lIlQ/c/cuZGlIZTDMxO
hmmwGSf7GHV/Bwb1a0RcZs+AUYcIn6DFSr+U3PhCa86CMddrBVRPwSs9F401
Rs3rz476MzVf6sBcsVjinmfzibGoRMW8dGl132jsEqXqJdMfxSaPKe8MPs/b
qB8etd7fsoc4ZdZi2iTWYKd7K3MmbGuq9FRJM1+aRQGVBlLVQvpkSEYMWHJH
b48MkmxsL1kMUnYGHd3XVzrhfrgYGMg659I3EAg7ujnTnGkBLlO2iwtIXSSS
DxqhLRb2a8dDvnreNmbt4JLuJu2LvrXV+zpwK5FvDEMzASGeY/z2VSAXzAg0
z4xV0px/yfmvSGUMGUEGtdzTMD8qwAC5dsOPKFhRp+2tQMLD0MYMoVvTrFSM
0pICJRSOmzZj8xt+bKDxq28gPmywmPWYIz1XSPWEKiEeJV+MwLVjzHLQH6HY
71hMJ0rU5pJZyBeXvXNd8c/LIX4OjJsd0eSUMeQDUgTGSKGafi6uicNjOZ1G
T2GqB2ebZ2DVT/1ce5cua5Ha5WAXlXB0sriJnRqs/PEXRMAoTxZqiswK6Ick
sWIQmHpH7PU1qvBFo+TEPNOmpALOhuN1zcKLgzJioPyVvjKpnvTmS2cXNkNB
7p23viiHzuXnI7I+/jT5PfdEqTcRjY3VhiSCywXcrnxUBHiE5w92vtKMmVSt
1xS/ur2AABZwiL1Ss6CLi5/wWLYkRxYaXp+x0KvPi1qJvYiqbXNz+h7AZZ3K
Tmci/7lSpcT66qX+FHyPSycO5xPxV+SSHpqPMpsfona4HlTrPi6Vs2em9mjz
P+ORmvKTvdYLEOahBmREOkqD7yvGjsZQiM+AO/lxZQyrYjtDkLcz9avAD+OF
YdKvz472R/7pUV87HxtqYCzIGMft2JZiCJPOvSrhqlP41CYoRfwdV2UuEQ4t
A2IDPipNajh5y5PM9VyL+5YLkPTcvvSJ7DW6Lsf/1k0N8UZwCIwtjhFqqWpE
uBVC8vjJVOzGfIA0QsaO6PByu1Jj2Pb/9bSnqQBpR6Yb7Kj1kBp6aZu+Va5X
VLPST5CeL3W/86gZ7blFLqNCGxKqgglPE4EDJyR6xWZ8J+oDJHvUrestMevW
Stg7EVawavARmAz8Y0IcwpRP8Fu8r3xLyMAyxiYem2AifWNUC/CI/dr7Oe3E
W1lkyItlI5Gzj9Iajqhpr8XCzy1mp43z9rpkXqD62t118A6UqkKTw+QQhfUl
JzuZNayYoc2Ynn0S62NnX7y5YcxVh26PfSq7BZLyD80oBMv2TWQ5yHc6ImtM
KTxX1KYFRj3NNNPnj6IMmhssFKsKjFStave+FhxCRFPKKuffZLQujocRMK16
lu/x4gxyeDMpaOeGtfSoe55QfkeICi+UNRPPTBybpYo9rMRnBN04CRVus4Oq
SE31CY4z+Ssb7vS370NSrI1UTWxGGsDIabGzpcozjkqYMSc7jZuhfB3kMe03
gxAC7FOpX9ksWeDmQdg6o744lj4YOYCaz6wMbEqdDjp+z4RSbRiyFEhwwvt7
tL3G1VPzXBZZ1/YQzGnyQvm0jZ/QPVErTqLN1z82zXuV9i9Fg+169M3jzeDM
wOdYuLJAHzLpQ2bw8ORo01YXCzObT1v/v2HsYSKQWV/9TRgQ+xqNWaVM5zWe
zgiClmqxR02h32vXQVdrXNP9gg1jSPWpg0b9iMYYhw+Rr8UwEmnw8/CA8wFu
c2pbVceDsIt0tBQhDc/pJh+7sB2+fPCnzjPYO9StffL7VgPdzhgaWT3KnZMN
suffo1CuhLPy6lkcdf8Ty4nlzI9EDlS3ZEy6Hr4H94Z8TIMR8Zkee26oiNyL
XofgtpKyYxvFzBo6Q15tNs/3o7hd5GIdABUtPS7UhR7VKeK0MzVmYpxsrwRH
Vm8Fv2Rx92l//ahywQq39o+plChk1NE1ZXSdamsuQ6LYSR+LgkLpHHBZ4Chc
fZLwPf9zB9CnTMyx5LWsDQmcsWxuNfkZJTJ2kIC8Scw//ACQBQKSwJE1BaZH
hNqz9PIaM5WsNKmwnNFbJtKjYhzko1Mw0BhlFK+Uu37LE9KqU2HOv84xKqd5
7B/CBJryTBTjC/1rhCsE7L5VTEFKKwGLbDLJhFuVbR18t0zYuXDg9EVwkjR0
HCOVaixFmw7VEyui9uNfvXt4nxdGUhZeFPlbaqcv4foyZbqGsRfDj/Kmx/fR
y5Nd4ZiZqCap856IF80pwR01na0esrrul14QjmUmbP9SMzZb6VpRfyQ5nDsG
XbjEysbQou6oiHm/CJrsgSg420OnxzFlJiC5VJ3fYu0I3Yd2nSvm2VzyvDK4
bugtM0QXT/K2aPQrwwGdoUN+k448iRX4uhjm4/a3o4KKxCs3SyiMPJHn1idF
rrvt0HCqV5QSKabLtCzEiOAxaAdTCMaVminPci/kOaOG3CewoRfCdTT8feHB
9geDYK0Nra4z8E2T8tzYiwdhMhQT0NR4r2fHHvTX1SVcZUhhstwy3OxRlQyg
7kD5fb/nR61Fa+uZLE2G7C35lTwLJg4W9wejLwzWfGv9UHYBoG9kPPIh3Zeu
18h9faGQVimEIitRKP7rA4LMavdLaRBgn/DFU0bIvRIZHNEWEDY6B716oPdS
ZdV+4Taji4legf6NO4C/TIcdEz+GgyelFb/iJAGPAeBAderRGOg2lraXj98p
IIEMuwFaVNKYpwyBFqcM3vBVnv0h9lhCQgeskjGbfMX5XXTJRkN1G4nv065m
vhxC/8jKgw4YavCt6+UOgVl+MA3Hwro6lPagPD92gB6wqoDH2KAotQ54VdfP
wlJwKkda6xfX6fU0RjUXgjSc/4zKPb2ARD6MIUwvLzpDV4qX+zDIWV8DxpIG
9NytlmZ8mDvDtf7y97lS2011XYPz2z/Hoq0N9kHhTqduCKwdiJMEUksIlRWB
EeAN8D0wjdtK2j/oGiw+PjmubhEsjtSkIWCq2s464sVRaIzhsT/Fq6/X4sv/
0fxjIuNn6VR09oKzfeQyoqeIuoqRhJUQM68hjq+kCO1UYCBOoD45uhnXK6U8
WsHjJrIYLgPSJPotny0ArkGQYtSLr7i9Ny7jqW18/KS+671LUiTx8IPn1eqp
69rTbO4lUCt6IJHaL2Zg5Vc9nGlVn3pAMkUkt3JnVBLaxi9jB7+33DizceWt
zBsQ2yzlJTrJkaNLZaz2MADD262k4msF1niWSGNy0ylPMgDM1oPaREueYGMi
zuD/5YUrLLAAOf4upS9E5ecHch6bFnjQB1ducEmszVbyDEdzJJ8Bx+/zL2/X
PS7k5GhVEBlxMZeZvMK6YCmgU1iJytn25LYPh1X2MXNWxIr3XMrDWTVR61Xw
Dc9+AKZoBuraoEArlA6VPvncl6oeDm3pgsJPNSS3iwUd4kGjWjt8bXBqu30U
giugcmclpHrlfOoHUzXkFdYD/XS/m92A/2sz7KT9xEb/z4TOk3uftmbmpbfx
5x3kt2zEQ14PYt7f6BBje7DROFVJOyRmKpuHCmI17p1Lr1u+tRCmKlUzj2d9
NdzvmJ307Ata9iHqv1HZ0PWAfWBDelNoELAuYemeZg8jce6b2dFwj00+ABv2
9qYgjiS3hffnw/fWr0w+QYtUiSgsMvWVDZ0dO2eChE6BWzTga/4Hj/bzHMoo
ywr6aO59vY1RFPFH8ppNf9CvwCSwkC3eJDacB2z1LvBT8oRUwWeCXTV1FVx3
8Hl/njfw2umUhXdwfop9EomdOow9cZPdbrQiXAMYUQi/CreG9pR+hQcdf+lI
8CcYi9yEYq+3r7LJ0HsbFa3RPFlqEr49qqIXRiu064NCLsSato1DAj8pG/lR
y5WldCpklfI4CGwTRM4PZFDrRWbdStq6iNr6Uj9366m63Kk3fhULH8Ku9RyI
QgsIltHKbjqxSyMsz4pZnwZnRkrds+ba+TTgb/eMHswif74tHDT/pQFJkyrT
Mwma3D9G7aUHb2rLv1W4SdqKavC8QAPt8Sb6afS7bmNyLdURgsBUrAq/wPy9
jfwVOARDtMor6+Ckg/7d60EsJ+4XosDqn7UaoDHIPLMDzotuXnqcW842DBon
wgSfQLUu8ZE0c33W8/LWP4AhZxVti2m22KMWFsZIUamMy6mMtxhJoxLKb9sq
OyrYK26Eae6ikh9CCKWfS0p8kBrLXHbYHjE1rJPtkutITw9Zf8YnJG3nc1SJ
s48A3tKAw5nXnRf3wz7U2Fy2t9AoMhiCdEdQ6uWP0VEM+ebDU72XPWFqZrwi
psjaBVmD3sQdyjfVXpxsWx2PX56dkzehUANKfvgndLE+JMTSQoszmYzQ0SxX
C93sUmMMN0fwjREdp09d6qPYTj3zQKc9+UPGITHI2dGerMkrY1TErgDTQPjS
SuINefSfAK2oORLKaLjxq9OBhfiAQUySK28pFCZGb1MRTIGEwHDhgLtrvpB/
IaqccVZa/LIiEZcXl0mhOWJrKfLJogpzcIufLkgpHWQ+5CvbaR/k1MuYx5kB
ktK6IXi0uFJiwbpcgu19Po/vsxsI9srW2immyxS7nYu1Rp4G4o2EUfjHUtKS
b9NvCCKfbe8zIzghVwoRuUZISL2NFFc/FF+lqBM1DHEgn8sRvcwWYq7I7r1z
IsrTMZVhPVD1u28RJF2k38SG+sBDWoZjiHX3rk5/Q3S6nMNq6odhZKFW412D
S4w+NFiv50EsiLCwY4Z0kxG79iMDzG0gq05JKaVatIHqCS7maC9rzuEtZxbT
lqUk6U9ymbALF0P76tLPspKVzXgQNm+9cnlnl+hf6uOZ+1QHhSs0JhDl02fv
txkmkBVdLlU9/bnY1scgTxybsNAFsjcd8R4JRsbh1zAFrjYv3hM/PIo9iKfK
ECQI2V7n3KvTWAKC6zEW57glCfFdKlR/9ZjAdy1iRYHTdZIGUVXZlU/U33Yr
DDFczw94NHuvuBpxvEpt7BQRlMv4VzqZROE6qV099D45hOLSY7JnksgRILX5
d7l74pdCpyedSvkCvSkJkbLrLIfocEnuc5AqB0cS6HrNz6G6Rix7uiW7pZNo
2Be12Zd0e2IDwvgv+l0Gfy5UUFg1qGXbTksQX1FDYXp/MuFD677T1l1IHwa/
uU+FZzFs5yVPx/JctrUk2RPZmHK4Wn8Qt4+5IZaY7rRpyDfNVTw4ysenVQv4
nnj37/18pHhGjddSf4O4WPwaCCVCXe+Cm4BkTODPzB4xTo5jN40PADFtAktm
y2w39isbv0QZAvSm9VbvSjYQjR6jujhJsPYJWOBzAbOfw9Ka7Ybd0mixgJnZ
HzWOtGguvlbiOUYxtOeYM1tAJnunStMsk0KRBrncjLTbD3szS1HQjxbiWExw
EglKKf6vAHGSNspordaunrbHCsUv0ifMB2xR2Gh1d7guDX19sDslVsh+vJgV
+ufP7Kc6AwzXRlEL2coF5si2oxUu6zR1Zfnw6XIGQP7eK2bHidpbmVqnZsw0
HjjmMmNNI3+A9hyOygDsFOgN0S91RQGEyhOfAH4dDEHZy2wLwMl5vj832bxA
GM93DGYqdWqO0IS68rfIkr3wRfZMFhQjSIQPhBjkE1D3li73CJlLNWoATfO8
WYxQM3jFHX//nzE1UfWeHi6p9WY4WIiO0KTGTOkNq1vlRdmRfpPOczHrki4Z
6hFcDuLRiJ07w0dycuhGatq9gDMm22Sbw+141LA+6lHz7nPJbOmmxsgugPvu
kXxa8iIkxl+IJmJal9SFnVKz14dKLSy8K8c9qXmXum5MEqxdrTMEpAL1Qf5K
wonKOsPV1F9uQxQpuu+QGcrag+kN7sQjyHsmGpJp8G9RmMqDGZn5y40N+2sN
DfWZzvGJ2SsVOTrJHpHe80EfxrZeyP8RM02GLOsDS36PpItvcC+NAYFH4HEq
WCrX139dACbARrRztd+BwaSYgO4lkVEE8FR99lgrMRjmini4OptLDG/eLOy7
EZ16Fe0wdAlkKSIFUQIRx9m8JSL5VPYEdwdcEgSn0KSygHxCCiRFWvWXgTBb
AarXfslWF8Ftkyji9fq602J/kpDhFK9ELyLxfSGStOFH0d3bYWKQAWhqofnw
xvH40vf/9O3vdtCuE4soacObRIe0Ix2NAejd+s/YQNOZgPdVH0WRKZ2hTngK
b8u1XHN5qmrhAhRKE+823ceIx6WW4tLyjEw0RACxFP2tokUeA1KD8xVHvUSK
u9BUYztdM3sBV1Sbils/q3UYcIb5IHOi04rHhSxA4WtHe0kzQdkKZrlS/NUO
mgEqLKenrTLmaFil1fGcfNQW+u0B/0Wt3E96Vhy/AvNTj9QLbOODNDRgzwnO
vxVKs8SbZq6qd3rN5nfaXjKwK0/DcJKtX4KPH0UP5cE0iz7M7wYEsuVS9Ofq
ICpbUWUqgxwT/jWIwDWmE3Sa642cvmr44NU20K0abqpLpr2RJIFHoF7fSwCl
8lgg0x+jvYu7x3YXY8n8iVb9DT3pqjnDurbAF0lhjiRHcbJvRNRidkFNDJEp
2iTXqfBrGbMuOLLk9hjgNUcP1lOsqLHkfRFG/ispiDWjh47iIjfwqU1/+Gbn
jDDRpdLkIDPOLulSBzGF2kCdlWq/dZugqNkAQs4XXSX9WjilQQHY8iziZ5/c
qHjU0OFN2C3Prwoh02wJWltxxhZexhvGo+ZqZAT8JLpCo7yil3ntV7i9kEVY
NYxno0Ni3h54JOQNkIG7Pic+vmTDyekuhnPDQTIYFhDAYJReW5BKhYV/Gd/q
eyJK0s80ys58G2QKUHLKZvz2ejo6eUh/6oNwqN187903VXNyyNhJ8cx5VvDz
hX0Wd8iV7L2yZSwTLrLmTEksip3hI7sX6oc/F3ZYbE5dNTCZ+Nlns6LRS7bd
ifwbZivyENuyYxl9ZjObTObKkxvdEsOPmhk3Ho3Yqm03pSq89GiX74FRVqvY
8kPYKKynsPed3ZggsVuez/koQP0VDkV2km/qdtHxBmCp6Pvz5JGB/6v6im8K
0H2CbFwSh2JFF7HPVqCNCgBxuzMvM7E/96e7M3XdZ2WzNUiqSKpA9EbPTHOU
2gqWpAa1n01+5OT04DC6/ranc9oNarPoqhzJ3EZOCGBe7Ni8tIB77S5yEKNY
SFQoxX1L6yjA49a0RW8r1XZHpQpRpq1E7jlytYAJZBJPJ/OpCOSH6fZc1rz2
iERPvF2WKvnFF04bn6UinKB4V/lwji7SsoKe70O+7rvoA/cOyH+eGaoKYnpI
77LM/Y8vQXU4qoxSWY2ZFIUQeh0bWrB8gjAROhrRMSjf7P//Y2aPluvW434f
tttZ2+qIpWcEh/t+RzGrBsfvsTdZ9SDgMRVEdvY3kdjn4RCdjFob/HDTkfoS
wsrMlB3KTitvHqj6vUZDm5xeUYR68yQnSY9+Jimh019f0O/fKA3T4lYvMm4O
6uTQES+NWGOjjzEoLELBzZ+wH9qvS4O/qJ1QoW+9AJzcUeqDxKp23KnYXQGq
BOPN8yBJgWl0sNdHTKf6PptMS+5RVV5hhSmbGzWfbLmTtqoJeaiWJlhaHB1c
5n7qzbeS+o5iyOo134+R+4IPIvPamckL5hojUq+PLsitOddo7E+EEeVeuN4c
3AGh3IaX0ZiFIHMrkRoifgfCTuMx917dyFqMgIQhDLsBQlrD7KDJXGe46sZ+
8Jk0S0jkwq8Zkk9WpTomlMz9F7LKHIwUx+OKq4MvnJCxEnA6E4C8nPBPFiuJ
3ADpa7xAoAPJCbKrD6lGcu+p76Hfa0k7A4jLQHnT0Gcikc/CFTJR8i0s+AhJ
oZDa2iHLOjrIJkaJTVYRTHIiNkWxqGD6ES9qd69h97V0EU4M96611HTWwVfN
0AXWdK6A0UuB1XjHQO1AG+Eqdn1bcQ4ChM40AssBJX9QgZqNKDbOAHcOcn6R
EpUxmcFzilUvlYBB8MzQjJaeoFy6sxcTjEWDNZ9tXQbKbQ0TVDAoZGu9bItH
BtM+4OjNa4Hk1e7SO1JGV6ebiPpFmL1CQ07Gl8XWs+GjetLFEFPXAN3Pd/YW
vgswMRPY1fgndoXEccciW0Gb1MrzrxhPnh6RXyLicFX6JnclKwyt8RAXjsji
xhp1y42b2LcU+qxsgsCSft4saPlGpWeGAnemQBzB7E9AABCdaV5AAldi71iP
ZACFybNwKKvK309o5+VZ36NdoDvqG5Gl/zYWqKSdvIb78vYPns/wOa1eLR8k
YaZz1KEbXcjdil9xt7TCaYiRAe5ib4HYhkpWNC2VzDmS7JMkdPZ9BD2J0ZkF
GahzpwtQ41UpiXUgUQtRxWkCVRTk+wpWAlBwWvmneijg4XcaidA+JbxbSvrH
tsWeov5wGr3rwrY49jL5+Yw+qPJEDaYW3e4gus2iviLRXWxNnyA/NGi7+4WE
8q/iFBY49SWd+sdP8ykO76d0DaTi1J6T7eNyooTn+oIjyaqe/cLZHKjvuvwm
Ne51DbBJkJ+FVvHAsNX9LGqP9GcD8KHsz5fqyf8Kc2cinzWJ+K80uGNQISlz
xw3yhNQZ+80ROmXHaFOZcNzpcWMkzbKojIlqe10QS/HG8/UVp8kpXrgHClx3
SNokYrzFP8Q1NRmhR7FTPMMJSB1VT5ui46zN8gmpKbOEh+uMsFKvFMP8TJ0o
GUpUVpm085IlXIlBs75Y5pjgic7KgWsDM0ef4pUR8k/exKJziEYpjMznSiIq
rPq8pMMPYAgu626VQMQ2iZb48SbOLZ3BN2cuXYsZHMlv6NyCmpC7XRI3n9Bn
816y0loNSFtRov3YAfdDCRLsmXsjunfA6PQrx7WD+KeZuVH7+lTxe1WVpPVX
5PSnxZo+lIrbUVwLq+CWhkGLZrTcBymUl5DgvnF25s6gshSMEWJo+Q7XV4uv
C/2g9nowuWGKky6KyJK2hgED7Xtohykj1hVOzC4ZipEwivv6bec9Gzgiiavp
fDWJuzk3j2hYwAkGcXaWFRQKYD7D9txqDNadGMBpNw9lO2A8JA3usdhweKsU
f9I0HtMJE/LOGruNHipL1QM9H9b8tG6y3NTUMGH8Rj1NpcB7QmhCfimo3WDm
WyI9h3HXluFyiHa/QJbMZwGPnTYyJiX7r6qYKAzajZpJTBr3WtUeapGqQ5nG
bzZSbTRsS9zC2yp+zO2+Yogk9EB+xoldh4ZYN+LmJTSLpOi+2FqUlQ7YsSnG
TSAc6mYhK9Q0/7rPP/wSlfhHxzSOdNHGtR/BVD7z/Bsito+QBNeFdCkJ7/tb
hkVceJmb15eJ4EtYvfHmwtXNxBvVfuaDL1v6UEsWz2p/y6GvWRdEttHNpy6i
FgTKH8Q+tsb/fqJ0JpTD/QtGKVB7uqh7v1/usBwSXls5GXb3mGIczUTPl7Ko
1Q3ZnqHypGH+/exDx+tj1bEQ0CxQcNlgSnMeTy9Y37mjwHTySSQWXenKgcPA
s+dDjsA1wVJkm4jdyAO2ENEnB/0ybj7/MuJirUGKUcppNue4v/T1ZjyF24ly
M7gzXIZeUHggyLMzrhWr3QHNqyUL+ypcMJqTtS9qtJSQx9+tQ0GzpHtGunUr
GjTVCNAPtURXBGqrMcCRFEnzUKTvW+eSMV+MtenJpUuD+aF6BvpEVuRdgP4C
ysoZ2sgQbNOXdmuQOtaRxBVaAzp62b6uMkf2QYFD25gvO5S5di/Vip97dqLZ
Yg8XsUXyhMvqNWOyfPyQ9FxGQVuU5ZNy99mi+VzXy8shH5/6H3rlfWTBhA90
HBOUxseI87V/pUCQKPsFyinxy7yDDE2EKjm29uO0WsYfLxH/jlcjR7fUJYGt
0PKKX4U35JJ/xibBxpWF08MBnSqFMFqPe5OMWjkRfSmcXIncumSEhpkTk5K8
GULSPX0UKFXCst/Nj8zSR3xzHNNSXT4NwxgABFutDb42MC87IS+2tRs4YTZS
BBPCrgFgJmlEHhc9vXLP4EZm/JCHvgLsarnW/NAuaR/BSxLvIz/At9o//8y8
rwxpR71nW0t/4CIM34Rqnf3rsRYAQJphw/qnjHdefhW8dnVeL9wezqFgEjuP
jnTXu0ro7Kr0A/iQ31g03sFjvZf+339XYQYzFfnqnPcFbq+NENy3Sey2hx4J
iKKAJv+v0hfiQyb9Bkb1/fInVYAaC+gP0+gK647m4+3SEvyPh5/M8lcIpJSY
Oxl4J5c5mDW9Ork8FTzcanAmtQKdONlslAgcAFVweU18YpmXymv/+CRFBtge
MUaksXQsQ2TyRaCdB9TL5PJ0v17Z58mPMt5HDjNofS8ub1exrOLlBccL7WWw
oQ7z+JO6TiCJO+D1l4D+tmg3Kq/jAKyxlPW1b9RnfvImrMcw1eSY4bl+UcFE
cRWjN259h/3H0ZnJfuf92YPP1uvLjVkCjRNC9usEG2TyRuDYBYR/tjwl2dZt
6JdMegken4xLjmUj4ddI0BqiMu8k+Vdg884w+Uy1RQSdFFUpSPx+OC2ZXIWx
VGCruJky6l7D3JfXwjtahffcbPSmsX/ZbPxolSPmPiyx7FqUGvcKEoc8628E
pOpsJ0OxOjF52a5ufvBFqYJNudJhgY5GBHPCmHLcEtmcv4V94oB5BBvfLlNs
LKMbqi2IOIv1zvQYIp3FZinbczH1TDtjHKBclzD9kDoyrsRDwXHavf76ZH53
jfonIyoSdVddk5QVWi8ObvovFjSoADE9BOpxzjtTA68cvzQ41ex2Ozvy4MT1
0HbSNU/PUVcG52C9KAbCwXKcAKsiGpHBOq42HAZ4vLUnIyrtVO6bbHpqElOI
HJqlzmUneve+pCOaxfsIPsLLksvkTooMjqknV5ujO1HQiXSdH8hMT4aKkrj4
OpzBRW4rLEyycD1JWAKSNRDNxMmie6b8F3F8MKYFU7lys6kfzRM9biR3bR11
aKeb2xAKpmz5Mw22UplK/orVQ0vFVW60Tq9x2VnL0NI6vmBRAVRZgaRVJyR1
+PXmiKAfzDc3JDIuhbAAJv/23WV3h0QOF+CER21V7Ma1vXHJ55Q3VB7sAGoJ
Rwh6FJxCEEWejM3tjr8iL/cwpAjlH6DHxXIcbDPZkFzA5R5LzLjxtcddDvLj
3U7WY9R1vIbUz9wMj8t/aywj5um0Vyx5PvJ6SmmlZdNkC13m1w5yJshynfPM
3mhT/lZdstoIR6VJNfEgVJX7ihbbPWTk8NNlhprEiDIw6EDelhqok8+rj8+3
WCDm31HhGqaP8qPUisij5lZUUbw+MtMLV5lYpcFQGTfMFKduTV805bagHQ==

`pragma protect end_protected
