// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
0ee1xLheXXoW3BRl4CJ6o1bhY+T2r6WdrmvuwwquH5QX4cIVvSsgDzQi/bsdEksO
x6X/fh74oIq/hRS9nXFGaYlTjpKlGis3fp4HvTBlb+UhIoQuacZUcgOnAHF1IV9i
N4/SjduWrzliBY1/vSS0/cuFmeWjCsZ2w3tcTvi2F44=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 418560 )
`pragma protect data_block
dkn+mG7J2Uufnr2kF2JgfurvBZQvTT4jv+BD23h3NZN3ecUZ8GMPPRXy4V/pJ6kQ
VUrHbgHXsNNu1pWfngjYQxHrpUNQvJQd1zQTvlaRw6acgUDMSlumLwXAJGHdGd2p
xleubqSq2NyoBUVgP+soxxNQgzQKkUEK6ewO68Qhb5AD7HCVVvCoHvKy28CBHcG3
mi2zrF1w4S4u91V4i2AL7VAGhVhS6H5s3pn4LHfnxRxxuDcnxywLEXFTP206jJE+
debypYo9IluUvXxivhCT+lXJ3UDWTjCdQqMEuq73Q+8Fwyi61jNmmzaWEyoAZBhF
0PgmbFb3ExmnOf0eYXPBbr/GDVnJHKPzpfKo2LsD+xHA6ODzUgllbX0/7HO8k9+m
qGBtD/R1+ZXoB2k6Y5LGnvB+9WoxvpCYbl5FTDiQEudsgqH+MGzziikRfUgapQ6V
6y6zyIWrc+XfSKVOxO1ku+HgW+ZZtOHPfQajuX1GV6lYD+uuHuONFnqx09/ioxqS
zLFzf70VWJvQl+/gqktq+/cnr9y/PEuvvRNUSUWnw6HLgfFUECodQ/MFaPvk3y4V
CHva7G/NDhR85YT6ReIHHGEeJhwM+iGl85BIVrDKYySuoOl3PBCS50L5gh21/IHS
GuY83Jq5jiTR6hNPwNhwDQ7Uc/j3PloXom2MKCEgnr6IQlYpsOA32HfchtkM9XBF
wbhoS7+dyyphec99cQSzRsvGBTPp5ruE5s1REj2sMiyApI4NHo4gm968lJQtyqcZ
H3lw/ZMOSFq/mHSDcg+Yed+lDHzmeh43qvAHgxlJu9QoUf1kQMFfU6XBQIjXVIw4
Ic/F3EiLkkVoUcQ7M2+RvG0b+OkWnPK3k6TDm9N7uGIit0Pf4K6QGCR6Vg+hPhwj
BP/PuKUcqtb/GvQs+A20mDENLagNzcV3bOpBbApz0P22muKCnHv49PBi8IYI9s3F
wpoxkG8J/obsteq2eaP5r2V9QZDA33A6ibLiS0bI1ThDns3/+KR+56biqz0AEZ8R
t41fl8r7Y5HXNnaoBHS+gtWF7NQ9hx/wEiHx2fQKIuHODMEsj4PA/C0BEN306x4o
pxlLMShxPJr1vPafpLZZ/+M7O8ONMyGQykNBVB1Jz+DMLjhBGK/N7pYnROEeCL4P
a0ONCbimdob8QXbHj7GG5EzTdHjLlC7TTkBcCJNAFGaoZyZRTbY6q+Hv1FCEzxu7
ZpbuWox44rwSz9+2WN8vPyy8XfibSV0dYVIOqvrzKrEbxLjDpcwS3s7IAScH/lY0
8YeuAEBKHGAp+YFfS1pT0B2WhJG01kN511eexoTu3/4NKgg/xDGllLNALkElVt2z
GTLuZrd9vjZF6nckz75WaimNFFxUI/jArcIuzHxL+BaNW9k4C69hAsFdScPN/cEz
CvnOi28mRUmMYHITDBdI5tItIFyv6NPh5RInm5A8eEjfJwQ3GvjcXCa4eWcgdfho
VIUVwqpnRRrP9wG77dRHi27twMdUtP2sYxDtA3eXVt1W9UgmeRrAHchLOgFx/piw
hPbD16uwBlXNkn5k1hj3PdjQwl/KgqQbDTMka1egJFiv8bDG/ha+WYyBIrv4AFcQ
WgAT8lbuvWmi5tI+EUUIQDYHBZ+JeYimm+geJZB1+6ge43cRFxsvBFwHdLu80NxS
w+aii0b857mMm68BgB0mk5vD7ityYAzqRED6l0ogLkpOZrmj7l3Ahmr1GwZS10h6
sSjjKLMvFADbzy/PbE374oJOexXRMOn5U4C2gIOTv8S+kCeQi3WEaIi29f0bXaHb
Qs8enWmcGfyG5UeNzRuP5nbUQvGYp20UT891KFv138lJTR2PMqRtScdLzdu6cyyR
o3Ni8IUouR39egDpttW1gA5BxOHie9wFyvITYFOx6sho5NKGRFzUEj0MxWI6beXU
C6bgNZvZ8cF39rLzOcAH1HFz2VVOqKd0Im2P58mDlTjX/t6CgbkvH/CD8ND8hKWP
3/JKev7N7xGdHJWiTSKNc5JLudNu1l0ujVXu0z3Fo45yV0BSHe4LPAVyTI0v9bdW
8SBg9SiOI7c33z5130Pbqi42N40pDNOunfEU5cqxc/U5VRGnSO9f76UdT0muWfzz
+9SQrCT5EaxLg82xJdG+Ve8IQWMb8RNCz00tmp7fxjSIB0H/lvuzCmVcpk3kDAUp
o9t0BIA6EUYgUYWdmlYdnYv6BYOZfGfaqF9Z7tsYkSONlr2cGot25InnUaliegUc
aczktmqjulBhGIhRZ/SOBU9BJ7MZhJSBuBOC6SnmksOrrbBn4UWcjUKh3cFVjL2F
/XL/VC2qykJ6gxCXHwwH6oESPaexk0FOX5zt3cl5EvH0UnjWdEoE56A6jnXqRDia
0jhRDLlEcOUO+4fVALRs74CYGE0PTzURgR2SBslnImu6DLp9it/WJsmXn4ss11Sk
2R94wX7hrl6t9itvnw0nCFgUY+x+rz3TzRIj8eJg8d//B4JvHrxEXXMR5zmAqUIM
4znxQ32DmikASD6/yjuB5z4GBRAcPDe9mpYcE9TL/vic4HTy2ROg3nWlayBvtLOV
NThn1YAN9T1afqnsUi164nCuxlIKcJSRPrmHYl3hEsy3IFzoU//taZX52i6a34KI
0I3HeF82/Sz6eQN+15o6569Ne9tr05WW9jWI1Anx9YO2fkJA9Hvs2FEYaFqHPuoZ
vjq1+zfTmIfi2FeP2d/ygbJHi3Xk19R2Rp05BzDZPD1XA3K1xinnCHL2OK7l76vD
Ss9EzQMctah8nKJqV7PKNENVRtLayKChoh2jRzmgbIgiHWBe0P7ItDC9JaTW2/Kb
Cy0ZIEGXKPD/7stRQr4dowE33yvUE+N04Zk8cmsAkPss8nwfMf3HoDyV2dw7Ah+5
BxhpMo8TsRVqMSFe/PEw2/WNnviWqWH+ACdbdJch6bTpRTvc6ZcDxr1QA7imPTTv
zvOfbxBgxRwYWWEDqsXNntxcDbxyW5ShdZ8hr9TRnghE9ySd1usF7XI2gvaIlkVJ
jPMzySVIt9Rbi3ibZCvRQkE3rybmCS1/8YaS+uIrjtKL1rMZ0sWoH1nJsdfKCUvj
6JVkW4cBLtKdyVoWnMNpPuVUSLXysmDS7YKx0o9D6dMsC2lM5vnwoBGI0Mn7BmBU
Ynj1+R4Y76BWV2LzFB4durJDZ1c7jOlEHVnIkgJEzXEMBTIUwtSICkHhB/XnNWs5
IaMxKQKJfmR05ggT+OXgMseEpv4JVwNXqklWDokriBRkeYePgxY7+LV8renoY7gu
tyv8Y88XXYhKkS5UCD9nqP7GrnSdoI7WDFHOcC/Y65WHlb6aGRTbt5wjSg0t4bb1
rKaW+yiUivmduCeHpd8FlvzYQdda4lrpdi9nlvX+CbHt42Ttu293zzSbPrc7al2K
4uyAc1EiZglpq4K2ju0reT7Dr5szP7rPUO9K9IVQUFDnwVup6nYaLMT/krNG6c9/
U6MuBXp99QKV02YQm6r8BXepGE7JiJ7EOmRRXSBB92W0VD2lxiC8iMy5xsVc8Syd
zJ/MP5fUQchjHA3xkIImgDAvKN7y8Rz+e9VhP4pL/Siwsv6vc4We5c7OGhfIWdcC
JRH6jLw3YkhJDzFLKMMnWkm55HVtkuesa4IuGhlgNuIBov4LVfjDU0+hJhV5Fhz0
SbgN5vlF1/8uAz1s7IRDlA4EviPRnLmO0IRIArCcl+kRTlQgL2lvBbLb049WapA+
1xeljMCW1il4eiQYT8zFlwIzg8DKN0DutxHNp6cYuxgte64uu7ptOezWwZHF5psg
eSNpR2hDHpxDQnDPWnyPnWQE/uUsmSRGZ+YlxGglK9jZerq504kLHoLaTcL2jlqh
mprJwc9CdGG6wtEgUuSpewwGVsM9ZpLVYOTBP0qBx0wOWXAfqlhCyIfXInVaKeIv
l78U7Fd0hBJfL5Q0WE4WtHC9CCuTW8jZJd7o3GhkQvNegu4tyan99Yhh4cqGKpOV
Gr3k5vwirbi6PRh3yGt2Y8ezI9vVOX1Hn+whLONYfEfb+NO9UnE7934vZvKYu3Ki
24qcDu/8Y/y+kICxk0vwHVF6j0XHbjb5aB1K8TMgjbk5JtDK5aYmdSiACoN2AySx
8U0MYGWZCPgL3ff5sY3WSq9+wqQisosTr6ihGjyYVxEyJe0LR7c4v9IUt+fw2T2X
7Lrjxo5J9VckKGCwTcmYH2aaSvAQ3y1UpDxEjyluax4KDoJK7QaExgRCV/vt7lYi
eSHszqBC9nDC5IqcHZPrWsEUZJTpniFmmGWtERKvOM5IYqyE1mvvCcaCXxynDljl
xL3Jn07+RnWnknNMEYgjykkqb5VmbUZ3Fsj5qEMwPc3jwIfK7YO1wVVREw8DQpAD
+pDKRbbrsZUzBfTB2YRRwp+rfqYwP59Tmuc3wfC6ku99SG/Wf6WI0kbwyvlEnQJ0
ZbO9Hkkd1wBFpl65HGaeRmzQ3GchMNqjGudbYOVkifHofjPHaXYurCE3heKryn3Z
MIlZjtAWtvPEreON8X21zDeRiMn+VA1neFdIWbmcuQeeTj1vyAY9Ut6u8VzfNPOF
6o4UkqiEvne9oX73R5B/eNPA18sve3xJux8C6NHLim2HXR1qia1zfzK9BVU0PRgY
kx2b/Ruvu5z9BYA4XRMtOtKQ8XjaUGEvy2L3V5TyPKe0PcIN5CcfpsnCuok6lv5R
HhSks3hfOQFt5+aR2zQvfSZigIHNjY+xPWDxRHDPaxs2c19sh/BcuIn/YFvWVt9Y
Gm7nkE9q1dDnRihFDD7WdSgXGUMKE8yKLW4yNAArGlsPDmfq5IGb0SeR/uvyHCzK
E9pmnI3T+GWP7ucplJ2v7gicHIi6BfsZi8XMzp6i0leuuznHd2JcN2K7m1MyWSE8
03c8dYRPjMLUkbH5IbU11XRnzSam4oWq5u7Kep0WxHas9yeCCnliIpvJWWBtcg1b
Bdto26+Qq+0VdxESlcB+2i/OeERTB0rwooZU1JjlBCDaj/lA6ceo6AvqCiG2q+7T
l2wXSHkJW1cLGgzF/o4SgjFYJvZkbu+m4QoFHxTgrTo/ubR3EeSZ84kwf0BPSn6R
gBDBhw2cqPMGA3pUy3vba1p79f4MNj4k9fUDOpxzPnk5HmdYq9qD1yIf0LiCoTFN
wHyZd71ZFS7P/pBW/AiDXiylhrxuXA7n+T3pZde3pKLRhSRjMDISfO9sgFf/jEcG
LOUHj3kVr+Din39S05fe6QmCgbRi/by5TBn5gHHiR8KSnUdPUiYP3+mub2LLICUP
eN9nKFn5w2l7rto5R3QG+NQDdlIK3DvdcZBEhQfAQbFEPHTOqo8VR0IATu8iJkjq
Y1SwPttRV6EKf+ZaPMHrrXKsXoL2m09LDZ8jyz0OMjKUEtT1wrqCaJ/f+Buhc01Z
Cep7czyBp/7/8bws3vlMVP2LGNVJ3JqHMv1lOcb6tgJKTbnB2wk1SFZuMOztJGl2
71/SYNrnSmry3XkrRvZdh5iheb0BSC9w6CQ9HNHDTiKLnDsMABm4/hMpd4yKoZ2M
yUwEHfNozBt7MJZHsOfjzdi1R/mNC174Z4TJyYEEzVYnU6VTio0NIZxbEAITTyNx
5JV5FD5hTxHR2owIism9xRZYapx57HscncVtrGzSPzqUk70Fvw9eN6eg6prKhiuj
TY2mgdzwsoztUvfcJCpdPxQb6U9dF62v3U9pMNYaWXdWE3WiXUE+uSxjiH41Oo/U
PREiHPhtrYL71P2jy/TeA5ePSIJW6x8drcu/pcRsK8MUNzdzeAnmlNLx5Dh28geC
8Zcyf+A980NZG1WdpP5imDfkcWjBayxqLiRpJ0YK+jlYPcyQKRnLIqKHg4uQjxVu
dEArAaQHqElQtAWsPLMJRe3JRfaErKOz5h6Mo1bsouvksxNZ/rtwNQzUCYDov+Kd
mkKeZf/No8sE7S3gi2IGa9NBusyx5/H/Pf2BIAVM8XaJHuloo+YQpsbEJLPhONiF
WefXULZFFBwYlT2B/NLP8NeOJPs7qeiPxNwUDiu3451FdKniRTtKImE+hSzxT/mk
9C/MvMj3OEe3yBLZwdWtlFdyS/ywRn88aZAysjYN/cgUNvD5WhrWa4sehkeSGzNz
gNQMFKLq5xpnRqUULyrNtA/Jp/svqpXR39PyYTAcC/n2o/Wti/sDArXqC/nmz+qb
byrxm/Y9JluDiufMoXYpW39ibg0yLw8rte/D0B7PuTCio6SCXUqCpYjLkBIBf4Bv
GxJA2Zgz4YlYEcdfbMVHwlseqD6EcA+wldl6UYmyGX+MDkm7ZlCGvmBjlcT39F/z
PonayOZ4Ogvvve6ExXvMV1X5+O9lEIMWwNemtOhBVxLl4nufzSZrT+nWC3JUwa/c
PahYnGrn9T1HAPEJaFM/0P0Bl7G/icy56dMuPX9PGvZfJhSIr1b9UJd1CvgeYN3A
yomy6NbSnLle1G8gtmLgH8AAwULddcNDUMJ64Qy9IwmmcXoiPNHrH7nb2ElyHWBQ
vLuNRlYXhurSvlmy0SpdGeptcNpy8mIIcBXvSzb14eSdhV/DYhGJMAga1Nm0a5Gx
cS/1uFhr7RI7PbEEhURtQwD5VSV4Q8a1fzXS2Jb5VkjlhIgO50kPkcgOCI8HcunK
rtG9tHnohDFtlupTO70aGgP72wpzPJE6runOWv/k8b1IvCf1WnTXHXsp0wR2iCOx
rS9+nohED1yVX9PmFUTOUtIfU0i+fy1A2ynGthWh76Der9/lLSrzr51WhiLc83Tg
7w9d0k0xji1ak2ZFxetW6MeHOO+k8h800th33WODYpcs4OU5tu452mWCL7qIbTLn
qxmJbbXkPogUYRR0j5aCbptcESOSdVqJ00I0iP7vH5mCoEBxZp2BrL9gjFMYF65T
MZepilxy0/WdhzcVlj8019mNQCzNQaKaIg6ywkvE1c/rYQ+6j1xZ57rfXzka8zCb
HJCUghH+mdltPP0QYcMzwF0GZv6ej6o/0w17awnSpIYNRlyAMf42x2YxYHS4LA20
c9tl5sdHA05fiqCl3bnGgH2a/SlWUJh46J/5EzwNrWAMbW5vSiDUbgiAya+44emT
jWUz7Mj1/s97s0RdkBR1MP9G8vaghqGMT5U1QZOkZm8xACFMJO2eV9iWRpzN8EIj
T40K6I4UUEwKhSoCY2n7NzesZwTiiH65m8jKi5qa22fr1XoZ9YEBF7esI1e+MwRL
3oEmXgedpwal4RKiR8PB8NoiJSADyjs/KO8vrYzBHHDdp+WVBLwzqbXm5iJiLeTy
T2jRAAeKjGoay3lQ6nJF6a6jq+HU+QRqXt7WNWsdxZSLYA2AUePnhBUo0tQBDgNK
GlF43Qk0ANOFyTlemvqLw/4iKm/PDimupdhIIzJTrWTqsOE2YnIVn0Bwa39TOEf3
mUYctcI2jg9GKk+kAJ1e9GFna+M9+/5Wq3CKnrhz9exWcmsWiUbVeKQLV4m8O+bh
pOcUlQtuJjeakvb2l09/Yu7y1PAR4AgjWaWxuAIJJVPpVmBPRrm8SCjRHKp1UUIf
mstl6cee8qu9BUis6zwcZ9lGP2G4j86UtlKw08PqX4UH5380qqNykcIYS5QZgBeq
NNsRSQXMpW7v87fDQXdwOH2qiLroxMUaBlZ4UvijGG0VNtqCZ4vBUGjVSXx0kR2y
bwWvZhZ2ITI/hT85k3J6a/neAdQg2/+xjHeImCentTcfbn0YInWN+RoNiPI84Wj0
HovOgndYfYdt3+3ULutbxA5UwcwIckz4nKqv807YBfU7dv0l/ml1crCUE4UTt1Cw
km69TnGBoUMxnBES645In/ohujJqU9bdq4MSveZXoHxG8ZJHHO9TjFtuk/mmtIcB
j7ux7PRrzU8gWfyHtBVAYpsczegbuPHqNfCHAo3bC/3ajOcesheho1aWH7JWnSUb
Y5gmWCf68/OyuXbMTYfw5Eee1kqI4ywsEyN5E8dYLXqtmkEmfxhH9rf+YN6ux0gj
1TlpyHxsrwgDb2iUcb96TUx+IvC9R/bq8Avb/7X3yHMxT5MVPjmaghje6CbxJUrP
C46ThMuOViDK6oZ+VBhY2HFcPwfEmpV+eJI56DM5d7wH8nXuRWWOG0iueAUJ4rcx
HyUha2HNW5KQpo+/62HAgH4KxFU3FTj4yDZej3ZAT7C6FiWU00QseyvdFcSchF9l
a5bCOt5BDSgODYeO1EuS7/1y/oP26PRJjqTEKz0pVXUHViKNh6XR2FdRl2Dryh9B
JSPV6c47kTycZvwK912/O04hMvhjOSnhRb+CAefxhtF2dNf8MjnPNTRzRVfJlQDo
K6W0TlnuGXOU/NgWa63zpXHUIyjZq7cfGsldOcwxPGC/ZPj+lMKlr0DZgf8w3eeK
nXO0UXXz4tTVnQ7fTISpOGeO5Ok4kh5Q7kzVCZikCZmG52YeFwv6OdFHEJrNaxpI
cEDSGJ90L7rHmKZuyi3crSWTdl4UFXpExph1sw69PSftWseQzVzn06ma6mkOdi1j
TXc3aA+kRHY81wi37Bc4oAMNUPTtxhX7DBeTlO9OvOg901uL7kwbOXMIMIyhWmoo
iZMiIUYh6SE4a3RTJhLvIcBxO90hIXwkvlr/2PDQxCD8Mt3smH3Cf5sewlZiTsOm
F0HRGgmEONsboLGRhB5sviNnJ0+MF+RX3t/NGteABpS+9mWFzD7QS0MJnEKEzn5H
VoNXsY1lFAdpDSiehOsGa4+Jl9/IF0wDtjZNdIgHMVuF3BYbp3g+VA+c3BZvW9wl
Fk+0+Mc536nY6rdHxTJmqVZE99H0hP6ogar+Nzq5b2GPQmw9hi/SSeeFX1hkSUf2
5h6br+/Sq5qvPHzAzklgSu3cw2Ah/7qIsv87hb34fEKoVaNsJQYswMQ003UBMR6O
sIqqe6dc/YICH7aBt8XLb7ErPSBA486UiUN9dtN0y1rrCXiTDjtXrUaLMKGFyORC
TO3LZ/E60z3CbUc9QuF1LEiALLYzGSApKcH52pMfKls3UYOrrw/2x/Rsz9OCuY1p
jLk21rEMGJKjJpgv1MZsgLerAB3LklENNp35637cIvsNMxe8lKSi0bwizcBZ4xJe
qcjAqYaz3MZSphL5Urla0/+QheCe9/GvQtdDacwgUQePRiU1zYp8ndCDwVAi6j6U
5gEsplZxl9fy/FXXqrVeoqGOY1EPBrugDs8s/78T/zgaYpnIUHeQne+RFt418a94
Y2402wGxFyYXJAwTaES63XfrHwBUIM21db2TvR6Wvc9hh/qqwg90NLPS/hR0R0Th
dGJ2gaz7xEnHUshWqjmAd93TOtgVzmWIIv666Qx14fNJeokccMhnWoLrJwRRQihj
z/JyRrXt03IVBojvVEaUVi36IciDO74z7JxkUAO95nBGgr2fqmp10uVEW2avP9L/
ilwb+pBEmRJgMJ/PFp42aybaCBuOEfqZOfaIDAQUvQKcU/OwLMSYplHSlTNR8BeS
835lJqqDDAk7IeQ9D9tjphNm3+DYCZHTnff+ZyrDi2CyOrivix+wUj8v5aDWUvos
TErnGSIfcvvdDnaJcjdSXX7MK3Vx2Lbe1KLX4YTjtOUaB8x0gb52YK0htnHseGHD
5LgiMU0BQkZW/ggB+J9Gc/suua8TTvWn3ZNqkYHtH2QMvdk+WENIVsX/JLTU9yn+
NPHTGtQ4DDAPpW4W2GEdexKSRuajQzuPtaSm4mSpqbTx92gdkgVTT901QRv8SD03
ccgIP8OEi44M9I6QvtkOvG2m8MOdIFMHpPFkT38G0lesIUinNcEeO/9htpiJ7ib9
MXTSPgTCKYmtnf3dFTpHMUaIuCjDJIdKCz0q+wKDeQJFqF6Tj8HozXsrlmw1pkC7
iXoiJe/ozE0V2ie/PvW2bMC9pIkmVrH4Vd4NAuilxfywJ0bOj7i6jOt9yjZB8p6l
1/KSZv8Wo7dg0mmdVeIPRSkH/OyjSi5cfJ17Tyhd/dyuOA1qFuV6Gku0lrZ9ytEv
mT6hwaMb+DUKR+6uM0OGIS7fan+2SjCPaUNVJe/deF+jNGIj8a9Gcvly5eraVHDX
5K64OS8anVZRYcraHFajHlgLxVI92webcSmn1WuN6vZXNoOIOXVN009tnMnmw514
RnC69r64bvRUS6Eq+v9KouZ+CQr6ZwIZkTW3N2szgPHiuIl55xGmYyAxc2JMLwSP
FXgOTvYtYAA9jD4zX5dtHbgbwxHfWKKzb+lmhP0vDXVazgn/r3oKFGvp5F7H4c6U
8NR6QlRrl3bBEcK5E46Ly+5tIH3LchsGMJzAp+OeNNC3Cax96lfaTQ5llPAQdFot
WeYpKfZJFHVMdbPmJ0mLUeQ1XmyxgxFXKNNhoJbZERbSVOoFoU8v3EA8u+AjquoG
Qob3UduzquJif6TH8qgrY3dkmbjBKqxId49cq+qIiZWPUgsN2y9L4FU3uPJJ1nTi
7YXuaxHQrX2wPVIz73YnkiWfcp0VkyXKcjY8QshA/B81c7TRjZ/FRZsXe+Q2N97L
o+FRbj7CXnykY/ON3zw1vrJCS+OlImNxjx/sxl2KhBvZac5ikjsZbdQLrNHVUVoC
gcsamM3Gn7xJtK/SACyAQXA8gT1tv4TiI2o91UKmrPxulUby73kI3Nm/O1rry46t
XVs9GvQ5niGSid3yhXkoEl3y8G/PLemy+ixnSY0vaRgNeq0faR1yMKlsDhV6riMo
IE+ZUVVT8Xbhx+ZlgdE7C26zpYlhRCWfBhrTxbjFAIedbNmnKHA7IVuiA3zNqvyr
CL5geMBEhr6zdpR+Mu1tXD0fUMdoht3kuAn4xXtOqNHhoHU+95gCGp8Q9klda329
FRnqaz0Rlh27QDyNMikDHHIGXqOC0qV58o4V0pG5eKV0lWQOPyBspVD4HoctEgNk
oBGqGx2XSvEF77YwFyCoPZ33hoXFQksAZQpCWQv+6r3zgiJ69huYXB4cdGADgthi
3Sc9QIKCw2KrkTk4BvxB/8VHAhgwsSR2VoX6Oc+vTl2Ml5PI3sv+VLV2vWH51/Jk
ycflQJOKBY46v+BW6w0O5pM1UNq+kKQWP8n9rmOS+Hugm/e8yFdEEzaPBxqEZP0t
qLcCyEU0i0hvCwDzXV+Pr/j57Ykd54S1xpseRHwVPsUb00Nn+SYOS/r+0IKC7spz
D3FkmjbpyznR2SXjCL7NkbHQjV/D6ljB+rrovZjJYzy+t1CJwShhixmrX1d3k37X
yfqwEKjfsOTCy/3KtZcUjrh1vc1vH+ric/dHk/AkOyCPekYTLD0MhgbflXd5ApSI
ExR16mKq5YWjmLYXWvQdpuDlh9/m38LpBB6e3nv0nIZfxg3W+Zb3coDlKAnPpvYI
SxQCxxwPsO84gNQrJx+xLBXb5nix87SS1LMb7vtE0+psSr4UVxo/l8IFHWGaS7Op
2bP0NJaJOl6V6iUDyGU6QDK7pAFAZSeA6z0iytUkaBepd0tTCIeAQNBzxjX5qLtg
jeur/WwXO76nEaBCcnHVcPw/8BhcF62xZsUIeCCDG1pTIFSPrmdC7HLteM8grRjU
1BdLsUcULcUwTeDXt8aaVu/pwY22uYiBIF7GLmG6K+kVCrbH2ksOP2c+akp0n0kq
AC/1bH/x7WyuwwLLS6uQgNImBBzLdBK1A/fIRHdXpxhg5QeIPT5tvVC1NFiCMYwm
TwdZmO1a2GqvfS37twYkwOLNneDbYv+fUf7YItDr3MVlYLXboTR6hmY6FS39QZwB
08SM1XXm+GKWz0XKUH2qMi4kDlqhC2kpdXWCys9F33EP8tgMPvMVwEIVdwl1ci5z
nih7f1gDJD+/njYg5WuWlWc1j/qK1SG4ZF8MzCELD5zeUK7ev1Bt0QsxtGcJHQ0D
KvhFHqC7QfC/YWuNsilbprSRcGL+3SnA4MVBhmfGvmTssuFgK/QYpAV+PLG+KTAI
f+E7Ub4FUy7WVgRy0dUpclKkT5Uk2BesoMrjny4BSag4RVyCHklJhY0/3cA+UFqX
GEANJM/xTSORQfhoCpRK1RMpV13i/al9eNnoccIASvTAtVm+5ZxZ8/stNKWJFUAa
+vj2db4HmSkarEBosgmqycIQOWr5p6aMUcm1EwWIZ39jOkNYzMmgGoGjNa4NocxH
kTIKRZfGZdCThxhblnKWsLDRMfkn4df9OP5ieSyhnQ6IgSjAG9+GkBS13gpf8bO4
WGXGjO1aupoYu/EuBEYDvV/l8WdsRQRu80Bgfp04BM+TIw4JyZ71FfO9EDeIBee6
/rA3qfwZMzYmOMtj0xtTfnATV4jNx5MjCpsHFj1F6M54v5psb35aPAQhq+yRfkzE
NprznojrHH5fh7PL8HrLq4qev1j5NagpPxPcKdhtd5BmPf6aEY1h7y3pIufNjqtl
4XWaQQ5Sql3H9LUfutotJohmNZoZdNQvngprwDrbBuLy8WWYG7JXyy4N7OtOzkAk
cRlMy4mFIo5R/jLwJx8oWFVTYYkvX0V8rg1PbBSGikYLw76Fvnpa0TuRpVuGd5Qf
yhlh914B25nDRFBwBmV656IP1P9VNci5CxuGu03HSY9sOCF62d2dCO00XBHuziDN
P1OBBnO5D1QkntGRPUwqALoolZP8H83DWkOrBya/CYRk5OiR5lSbrKFOWNc/lO4R
ZoVx2c2PYgAHRvRiDonVMHeg2EN4Pb3s8FK5jreVYmvUB14HBJgtpxvfL6HlA8LO
GqF4+MpXVKgO7kdzm0fB9sdjSnHdS2dHl+JRAM8dHOHS1G7rAC8h6Cy2aRzy0PJF
e3pII5eNQEx6xftkWRee0FM4haFWZQxBpbtqHdCSAiSR4kq6/fN5oRHNoxzBsIV7
Jd6vCN+Du2xOiWmxKjL0lgFSSLb5Zr7czJ/BLzOtkjpquOTAV3YM9DSNMUtFHTkf
fpnMuPrHuQGOf/epED3eF2g3Ezpae0NrybRi71BFIyPb5i42TViq0Mdg6oUJpqDP
bfNCCYq/D0aFtwf07PA6UEO37408jK74ibQveBWaWkvWnRo9GGEEAJA7KQ6yoRyF
ESywrbE3EhMqkt5IeaAaodUTBs+fG9+MlOZBBOHjw9W+SelmJ3jb5X+mIzm3wT02
I5UOz8iHK2jjO68rGqCClyyNuUgdVges0Lng4ebRUK6FulBPA3RDq7DZUxo4FJJX
FksW6lR9wc6CWs1tUBAfmIzpfmAOsWIqR2S3B9ITjBY9Nfnkv9DgPTRaT/izEDlt
SOKfYWkZELJ2G/S4KBO++/RfOMy9ZzPG7aDsTxTZq2Mw3gaNreGMc+03aC7EbCbg
XaWNibufLYYDL4zvx1TRGr2Tsx286/aBEwERmGvxd2dJ9ieGl0BfX8/4YNZflPGV
PI4g9OFYGQKosohFONDQuoEtJ+YzPJYK32LezW+onZRf+2B8rXRPVoOkSSbNfTXA
1KsIqPxgCvw7BsK766kabLCffjA5XKrdChkBByBqXdZcbZ2/4gzjgy3OJ/7fKtuw
Crc4HjjABDmccAXN/ykTBZJfY8xOBe4CSzkq4g3jcqZj353+BzPkESxyFsVgth/K
8HKVogLBZHGFu7m0+JH2PBf2b/Vl0YZYn3pI4Ry3ImT+4MlGKY+rAS7rHNtVO1Hi
7w1665uwzpBR3tYxTJfEQTpY6QOxH1r7s45htSYBhNZX+zM3XEh6IMlR1Js+svRD
jlvmvGhq+rjgnxatRRaTAVdBdCKGH0yTJ91b2EZ4H9H62VFgaxcDSyGttgXSSIWq
EzBxpVG2ybXqLOqmQms2X6o6FY45GQJXk7Mt4hQku8cN6wFPE+kwdETBgm+G+SYw
1dICIu1jOY0+icwD/J8EI6xoUgScv6Fc7jQCwicFF8qDgYmkN2AQmDyf7hZL3mbH
ksy4QaN38WCPEn3bz9FUIj36RZeAT8i0sQDU9dhB4+5UTxur9NB86RiFzaGD2nY6
iXNVYITSsuI3zEXfyN4Z6oqjv7FD3aRe4p1Dd8mTCjDPdrenQDGStAxqvPciptQS
IKVVfuhHD/yGF7j328wfXgNnKUwz+33XKF/IUaNO2iIfkXUldmqjxlWQmt77KhP2
gNktSxlI9X5D/+8nBvhJxPDBI0fz20VpvaJsFZgWLKJlgLgDl0e+utDu61zswVc0
RDOTakvyUMQ61Mn2J4+DLpAxh1D7DZVh91LFMnLVsonI3FJg95feGXYgfsZ5e8R2
X4h6c3cRrvMw2BFwvaP+WSqFKZvi5b9EdZRdPn4zoDVzqcLuJ8LtNSgrmEE1MSXz
ROe4CpYCPwa54xA9wwp35dVouwVYSDXQ17o6NI08CVon2uitwC74w9ZsuYZFhHRq
1FYdQvbq9MzKeJFg291KCpHrHUO93qvJQMQeIxZJFgFCt9zNGWnMyHw78CS7EcG+
hhb19FgyWL3zmB5PkUv2RbmaEyQYTr7zyAuixtWYWI7SQ78HjmpkjZTqzbK66d9E
wrQEU6O9aMuetxnCvJ8yr6skMD5y2MvegIsQBln/CP1SYT2mzFUCp9iY4Gbjp8sM
lE/3OxkpDZBLupLettfdYZus4YXVXh+9hJ8WiZcLHVAcW13DJ1iEcaKfFeF2zhVc
R4JTzA0XSHxLRz0iKQ2ZUtjfq7TSw4xd6uIDQ9OqBGagZkZj9oALHTTqWcCwe4b2
dmTsIdXqMZvMHKaRA2lVKxNdWka1s/pq7wF9qN9/sq2SWONAsjnGUbkyEwRBxd5o
fuZSfDsMagL4Ffk6+6W494W3gZyrF4c69GePe3K4+WZljV+hP0nKd1Kq1WZHm3gn
ernrvZvzoyf7XzBdFQ3z2YhzhJKZY6NNC4MRZ7azheJc2cVn2R48f/B9P/p9PSob
izVEV5rMv+2Tr/rSSR352O2vdyKWDWpLwqntWafxN9RT9jfj3tKrxq7o3ks1T3PK
Pj2Vi30LOyWC3MuE/IGKrNEuZwehck4lP2KCly3hesWIob2FVz1CSDvvXCSgrSpZ
QTZXYGlcKf97tWiT7/Yjk7fRyU4yy596+YtuY3BPKeFihbnSYdF73Zyf5P3klnlD
JkKHhDFEmwTVavtouOgpx5YUmfPl128MBxp5wHfJ+I0gGN9zURWEGY83yoBKgmbZ
UETjsREeJMIpUxVWj3QpiQBAmp43EBXNwg4OmhPOMAA+N8URrXx6cAeL8a7HrzOp
OjKyk2/Dlh5xj74Ma9gMGOV9QLno8/m583hRusGk3dM3twc/tvKeQzwZsm2KQGa/
hVli+jQ+dGdOtyjgZi/O4F/An1/HAegEg5oF23E4y987U4DIC2pspVc1Raiqqmo6
U/VrlEqqyz7N3ATmbXkjY3SUHD5zso3jwooGUECw691iCjU3BZBQrnNjXJONsCDQ
zYnoEo7C0C9ANxuDbNSUZzLM0p6W6Skt6IJ4pysprhSZ0/YWbRhpJ1DdIR+/VByS
vO5RC6OCm5h3s1dBYf1DMvsay/BSIgjf/kTwM1XeV0bx2zl4MqGMTWnhSFe3Af3S
NiPfOh2FQyZScuqnGC8GxzX5N8UzFp68pTUNXM6wCo1a7rDLcA1vyXdDj8Cez5vP
p4Ce1m7Iu5biKav1b5JHQygTr/E2VGCveTxqGu6vWzNHqAk5qDB6MdDd/ebW8vdY
8kyBHG47Kes/UrXUQC8JZZvlft52KPL+7wVqrb5WetYc7GZ0aStSjtWdqBInJtyd
tCt63n+nQvPHT7O2iiU32E0at+osnoYWwDV84Ihf8D+iMzxKFEFNDvGxgcSsLGo9
goY2FfxC3NlS9kJd3J2Ugesusp/hvi4KgfjqsDrx9Mvrr0Tu2HrSJ1MpVALciJ36
wUOD4Z1nLTZ+Pe3rNrlRpqW/xfo3GRNsNpxsvfv52LjIP6L7gKlIsJFmLE/vWtoW
BhwET1+EMBHOpS/yLmCGOsT2NiggFTVzG/Lyqrve5GzwvNvh3NDMI9aFdAyWiMwQ
IvWQYJ5hq+uqZNmE3xFlujtcnmo4YmEBz1WpAQ+nW71kknENsyO5xGF5BjN0JGyT
FFgt18PlWoQY01ELOHEs7h/vh7nuYi2X4vxbvVImYwy/Y6UzSUrm+6W6Y9bBfgmh
djus/ib8livenf9+IJGs0VqG9od4TJN2M4nGzLD2ts4oeXJxR6wzath968q6wTx1
FqIejiK6ut6XNLZ59qsgyb05P8m+g3n1yKhBuHKd+sQQfce9D/SbMwMoCXzTXxiT
iMTSJ0dNloINsTYoF6t9iHT3DwmR2rkDxjUnfRAHv1HQipG+OxToPMlh377oPtKG
J1pS3j3WgWt3c8e6gdf1KQRnCsE7xe2yS29b/nHUpk+yfS/n/63WSQCwX33T/Xua
tIf95LjB4ZjtsJM0c/ecPCY9nPrW8n/ums6SFT8GlGT72bh2FoxKJlCBAq29W8F/
5iXUiVD59LKl5CBZy5DKBsH3Cyf62TxctdcdWmGxXIGqYoe6FuqJW+3rp1gkfSPW
wnQ+ZGG55k6N3hhfzQi7eJUiJpYFn2aiN942U1lc7PFygZjpTU6oV+bIh037qZy4
IN1kcw/h8M2bBmjqaXgC1F+l89gakHr/38tRnBbvBRRl5sDSHCr2V+CRYfgbvm5O
TNfhx3+2BL5YvP7giLDUk2wGQueOCtqITcRJcF0SRoboFauVtx9s04l4m/5EIFqT
k7yP0l+JjK0ps6dvXqiNp4C1T/w/Fnxy/QlnG/lpjIBSoR/JesyCJy83CniV31Ho
8JadAUh08ElJLyzgl/8uTZrIdjiHKLf51fwxl0F+IGJqtUBrUHrWRYhlQFJ2DKsY
nrdVgjqBEgUV6sM61uTKUh4VecwNqAdqym36uI0dPDL9rCbrtlxy8gGST6qsh5gd
iT07IlTGTnzlrFvEFxZFMPnGDjeDG+9wgwlaO11chcnMWfY2UT+zWpj60bdRjyuF
jbogE9Opypjo5Fo8RhjRnUWC0k3IR8sW5OG8p+E7XnCzpL4VVFrVjGX5VZcWNlcQ
8ttopuxeNKEfTPvsLSNWaJkRIxf6Qum1ZFPAcVNGtrLdczuxq5/DTQQk2QX5X13/
BoXyUiYvH9qr4QKEFHqBAinvOlez0dQXsQARQokI8EX7HLgNH4ZsPe4ugmuvPJ1m
lzOqT9JPh4/h2lI2ZD3tqcMLQZ1HtTca7k5YSfEmF1pf3oeijjcLsxGT3KoFjrVl
eV/JzU02177uqTK6VksWvqm4ZR9GpzzeS7dbbxKGAbJ0hb9FogFHHqSeLRqsfyF2
Ywo89g3tRlwgLLApaMpWSWY6TC0kKYp8Vi9/Af7seY8+2oFcYpUfa8OZ9/DkQjDC
Xcl1PAAoPg54tezpyB6O3Gp//9mbhCRXs3lZvvj8SAZxVGbHaT2DfcAGOZeyKFp0
9zDP1hC6TdFld/jJUy8Fegb2WWJvNmAKwEvyRbWrDC5Dl8TRvlHXVuXpFD7ccviL
zd+IPs6qsM7LpZHTJxuUyD9ML2Ey0DFFqSWFmLf+wg/Se5MjsHUfMPF9Prhqh7bz
qpwlaBztPWi49hwjk8FIfvybM9BXxAS/c1eIaePToQreJunBTUxpxMXcYzk3oRjB
pO9wEW3h8ELknC5KXtfn5c79XDIrFcKX+WxTh5g+9yH2nKkSbZRWgLF69vqADfnz
dztdkThvRk8IovBwTfJr6R4xbOb13cN7OhMHONoRhtU/MkfWOdDACi0b6DHKAbVS
ufaOZhh3lVSzOKt+Jvmu13sJz2tEvXMqUxBCeIuNrGUPdv1Bc43W5OhctGCFWAGG
iYw+pp5y5bUs8Dm4AMcZEsbliEM1yfsaMi/tdpJ5HCTIPF5xhdtUheYMrupi1bYG
1TFeZ4H+WF+oGayWcPzr5ESeUQ7aexncQJzy/C3mI2/b+lV+q3TLD6WAVJe0J9Uv
NVxfaK5RsH/WIf8oL3ZBidLr8eOz7ba3ghtZpDJV6JoJhN5ldH3cfsIhA+ZqCqrm
5W2SQznJ5HPCknJKjMuZZb+htaWZHsvaPF/LnETE9c2vc2IG4tATKrSNiEkMaQIA
SnhOLOLVlhxwIiVMQ1pIFsuPCRYWta2Ufk/l2zQMLLwl4GAhl1ie5p0VIL0IuqGX
caOYSqZxCHs7ovWqb5WkXAXuOg/qpTWo7+GUwmgQ8Y+HYvWwyGXhUZDCMagwzegS
hWrgYkCuAJV5CRSQzwYEcHzisg0XO55GLhWQZmeDHsxjnfvwQTL+Klq1WNMbhn9m
Ab81zEfp4umTNraHnJgOPFiHp4Ussz+SvRZIg89ESFZjLcAsoriAnMdqWSxdIrJb
GZQRXhg5P6OoI1JwWWcw2QWWEwwN9haDps3MhwBxkoC3LEzjFaWX/HMi1M6IH73k
ZDaly9xPwzqFSWFpu9nX8CU8pOPAwsoKMBgrIfyJdbKnm2g414YKnyZEOvQb3nR8
7hp6s+MybkDCF70o4At3+UcsWhZ3muJ20QUhM09K49+Pgbnq5SHv78e+4EjjxxFm
zaGeI5JlTb10LF8CJj35SXqcXfpf11i3cJeAqaqFqoG55PrLiJQTCKXyq26e09yF
3kYGp/W6zfqx1/LUREpkeBuSl7v/u+wOp4R0UgNKbHzVgBxlXYAcFdHFTGlwCT1D
OJN9V+9vswd1Z99fap61/A2unty/kNhCh1X5F/aKz1pxfWrpCZ3J7lssqUQWjzCN
uLttXbhDsMDScM8q0Tx4ne0mrAtpQb7cv3SesjHOFlbUk48745onfgWEYHHvIynw
fJqCS1WRry4NtVhTYGHBbNpC9qNkadVaENHnyQYa+gKnOoGeB4gyPJd7gf+lv8jZ
8MnpMDm4BFM9DB+rKVNj/DehPPXBfJRUgnTdhAhIktGfQHt0ylzHZtMkTjCvoCEm
vl+EUXWLVrJQS/6rmUDpPmd8cSUjuQJ0pllzHDZPQdBvUXp2O6nKLhFkiVhnAvet
n17DnVG6qyKkXU97f5EUbW4tgZNEbHBitgJx4SUFDMbL6MSFODkuvrfeKmw86w1J
pvuo4utwvntOOuc8O0hAop+meR9H9S3EZFewO5aa4bxMDB0uDFzQtujds0+Cw411
xQZ9zL42ha8KF9JMIzWDzy6n94ymLFkiNi0vW1Sx6sS0uv0mJnkpujptM8vAT/Na
F4eZtLelHbEtU5loPnpdKU/9pduOKwqp0AcyHaTWpC2Sh929yNOLhEeHaHC10LfL
nuVY52Xwl9eRNhd/3U6R931iQqSSNp06zjLMO2phAjj6i0CWJOrYOUf8c8/xFBg4
agLCm7+l1yrHOsxHa5QWnZmwQ2zN8vC4p9T6vr40ES3Y4+xv8y64HSVNDavRQRTy
HoaiOln6fXTGbNP0UB+Z+b9POfRgeScROsQYp1j62J2gj2HlRW2TWUkDJrxOzGGW
6l2TtNVVWLY9tBz14XK4HYn5aY1Ao+Pidx4Hc4O+sB02weAU13tXT6/O+YNd2/uS
NJCe+2sd/uCiO/BiHXCfUZi60ULK1vxUzDCDMse1E6P1zUzrm74/oPmPcLaI6r9C
9fKadsZV/Zz8jtS3yyHnCsT/abmDVQfJsTi92GbEjbB1xmzXJxBiNNbhbycecJRL
SmQ1gEMP+i7ux+GCEl98Xx2wjjMomgm56MB8qBxOPmATDx0TxWMsjNB30A2V7q3c
8jkMwFZdxAOHejz0c0WZLk/Y+ICqFAe+9eS2tA/vM54jnPsuA7FZC7U2gincIVM9
Pj1Fso2dWu/OJ/bO0VpTnbjD/LAM/DvlMtmvH6Rw2fpP5TI4wnpyJgzO5R05En8U
7RTyq7ImPvxBW8a/0IyvANUWd3jTdDtD2sMJzAC0vXcZv+VUMeszgpy/h51b49YS
izpABP0yVyO2oq9IOEqm1D6bois5/Rwcuj+OucAnM2a7/+OcyUy3kokBcRbU1Rot
4dbbzgwvKUN+DtXkN9SmEbLS89utBxeKiVDhr4j0SnNs3N0iRPqYjs8M0qKy0Ni9
xz0Faw1IEkXRFpmBhCyLHWW/CgskX0dPtENvH+K9k3+MgCpz3Akma04Lz9oYihDy
ldjyTIcsT/hayKERSQBYmRBnWH/JMDi0cW1FnWmkewTXDnmfUi8+qoYLkPhaMlo0
KBOegrzv+cgCgpWwiHt9dwPlRg0ZhPw1iVdkqTtVd3FgTTo1tsQUzHyXHJWscPxE
x+ylHvmCBOjk5Mhb+lxHZMj/z0dFLOlRVuwFpZA7vOX3eqPvAxzBl3SlWWLkGnwK
lCkxkaklBopQeX6ISiOuLPrhksHrwrsqJBu8BQRbp9oHJN1QN1XQYrrdG/VFHgok
pGCRbNzbUwCRnSJ0HsoxZ9e4ryE/TtUhlbtSa/DMS17qJ3JQxCSYEvko7rZnQpmf
E76gSCltWlT6rcAQaL1mXEVKz4g7+GD3X1HbtDJeiqEny7lhbFH+XD6+2Z2OsmJP
BYzhNgJzO70DmfIutuNRQVuHcfHL1LDJrc4/HsPLXyrXBlBy6DORUi3xF3nAMUeJ
DS0JzF5wXuuC7m8omfEQZDAlTJiFma8kc4XB65AnjwoQbqRqneJ9F1DVHs2ylHqh
66dUNgZs2b34QW8gi16hWDW3TAr6jKMk+qddwMWdYCZOAlTgq+0Vi4o22oS/+z1t
dg3MKXF5iiEeOG/5PgU5Jo50z3gRjZ1ApqusEOp//k1T1zG7HWqtbdPH1lSjlI3m
Jnz62Ckk97Wtr65g+jX5nLQkfKHrA7bvNaM0AY98gyt4xv8TT6cA7lh2oqXu/sqK
JHtirLK8adFHVrztsELEMM0+/zJpM8zjb1UHio7jqe1250F1MeRivqYpWWdFLkzo
vQ4wH8xF6jMVrRyWMQ4d+Naq2Rv0vUTl3eAnzl+0jFo0NOZzqG6cRK89uEWl87OC
j7aq2NbQHMl+BgO/rb5m9FrFS3i0AAoZ2Q+8aqxnpl4LoyMKf1nnEWzSTyCckvrx
tyPa4Gr5HVtih75+2oQSa4AtjLuP0CxG0YApsZjFqfyR/JBoYKg2SCA5ysKzN2Jb
8wgjpbSK021Ih7nYDgezdtRqcoUyZDOF9DzEwH2pIphfDnVLFcDszeLWCmPT+F+e
ynL3ATXBeiWR19Km+pkGmwgibal+TG1GdpYaixAbR4QZtg11rRX2ooK/AdaAZenF
2utoa/1VC9phECp+OGvSi+GypeOde2Pdp5J01okfWl06TsUAK2oFdi66KyLdLGYH
d8Hcp4OXdtL6TerJMNV9molZVO5u2MGDRwvhNNUb0CcysVFcRrS3v0KN9rOhAM59
mBQyJ6G0QxV3lXAkI6zg4C4UxLIAZwjSVYHyZaLRsKN9sUWIN9O+uRS8GOD1OyUQ
rzC8yNzL7GL9Soh71etb1Xh4jULjqCMemg8k7tYweHAdzjQeMucd3hkf63TYUDPx
VEL9wBliIo3FXlI1QU15dsOqJMZxzyy1A6IOfXSxn9TKU2KyIOFDd2mHgm79+S9G
hkYFzPJVHzEIYHZzH4I2YK/ucpAE8LUG37C5/z8ojaRBGwTVzydNdHWYu3xk9I7l
ktZIqQEi8lcQmqV8C213813TQbrXEcmrHIlNKaJeETxRgJ/W5xU1kPy9clcfXAS6
ybFatTbhlSbe4fHL12cNrG9VCYXwvT8qL8Ly5Gs8jd9Pnb4/mc9oW+Wau8DI71TL
0pyjursanTdaYQlSF37vagcV6RlNLIUi6aGgThadNCQsPp2KTlXIQutt5Ke7Qwz1
as8yNV0l9hhUz/BLDyUnJDxiWvKSsg5ThQUo0vkmpC6L0WSNbmzIl0TtssRDLa7b
AdcJB+Zp1rTsyQsfG/7rz0cUEiIl/WLKRlmE7jq8gUVsqdSxk+Cg+G6YM0r53L31
G4IWW2V/gxJ0/ortjzEACuH2cGTx+wei7cDBC9YOV795/XdavBloCcSVn3g4rvf5
OFsfUksWncx9wIwxmbhCAq06JJ31rz87M6j5uqeka0yGx6+ZN6TLv4vJhg23VKxH
wdHthCVhhYntTI1Ieb1ZhoInHT1qaZTx1HwI9FSJHwIKOba2cp9sXVp3+RhICaZV
+SdgXPHgygRWJ3N5miUBM4TCTFP9Uf5lexd73MnB8JSBVquHWaMICsX8LEvyTBBx
7trn+eGupfJ0evnxU0BfHzGRPulIKjIts11lNFO/zmwcn4bpvY8Pfs0XHGzDcpaN
+xxGdWWF6IZbr3IaZYqVbVxcrsYX5tlFp2FeAbM4dQ4GSUprykH4DQf8/rJ/o6PE
yNfMDoH8wELt6RSBJGk9uJgcdUgm2i77N/cS6L3nHkLJK1Iv+m+0oq0VbkYnz4op
ej9VsiTywaQyMWyDmcdItdfjHime+sJSsBhDR4rxcXUQTJ4aEec3oyUoDxbNbXlO
Q+HyDCYV8fN4frk+5pwj1Ptf2d304XmqJx4MoA9QTRrPXkbNEcLzyjGUVmIrjX5f
AX072n/gnODI8JoDb21810NyIWVdTHFc7jgQNKNiyRHNjKsw+Z20blfld1wxcY7A
kLxcLiaNvCh9QJnIPhc+xqNoJeZPHtDM7thDTbuBQTK4kDI3RW8gCjfxydvQrmsG
FicV7R0p63jIvc9JePzALPCr4JqEHydKdIyoUgX2oWou/68n+e1G1vMB5UiFsEKw
6dlBCgPfraQhAaZqj0buu9KfUi5xHAFv4kWzcDQ64HjItX1v8JTwCW6+NS0yDAfC
6exG5qQvgKXD4RpDxQBwzQKjd1/lSyVOrxHpLsBzu6i0BzptgWMYk+UjK8GAczdi
rLGIKT4+xEoC71KrMyB21yxCHtRCDIebj+KNDlX6dUk3C+ybFz2vLES+Ama3YjOp
8VHuUei7AJ+qnWCH/nG3/EoYudEEqrqpg9Ln7LC+m77HDFXJv/I9Sd9Ui18w3X4k
pvYZfpLDuFb44H2zBkQGOoIw4ix6JvJfr4Bc1miRAUPQqKFTXuxuXrpyRLm0QMVx
eSjJon5SgD6yJ7Lq2EyTbIndco3Hd4kea8E9tdAUBMQimZJTbUCyAT7Gf7nDS/Q4
Bm6X5kTnIfdmwlybWvkBejqDOZ32aVrCg7SEg+f3R1kpiQYkWCwuQ33B9LLGjuc9
DEQ0bQagW4Lv+cKmGsoM9yYpPsq7G7nTLpAFdY/RZ1dHuJsFMpZG9LZpsH6xvmgv
CvNOjvDC7gQCEGJj/RufTiQEwSDHodoyu8aAFgCPw30PTbZjtWnSOjnBC+++dwxv
2BYDLzqNj+c4o/W4t4SzbMuoJ6RZZefFQ2Q7KL5m/muHjqi7kk40gvipfPUYE5fk
8re+eNBG1QxtxZt1coEYduTJHqqL2Pb2wgwXneVScmVr3YZmd5VluNClIvLuinuC
qS3VtAw+2zWLcmcqyOWZihY+COk/aRZOnNydPhcU0TOTE6ZQLKxgKfBdx5PI+ucf
V/sKOsRm4UdsQ+zCu+Xmlr0ekVT9iRGvwGM39MWocbX0EeYIr1YRXoOfhxDHGyeE
JRHGW30CqSdGFD/ZZpPeUUQ3vy0NBrVGIj+yq8PqWKhqj3Mc9niZTLh13VfPFwNQ
QBuuLVyVaQSyOa0QIMsePQCREvzIgzchNq4/TaFkMhr7wSdzOSQSsOvV0dSmrduQ
I91DoQEHiEDxMK1o7eM/l+5e44rg+GqxYxgEGv0PaGg6cPDvIsGjNsf0kUqo3UFv
pAHDARSxxfP8JV7vgZjyJCKlgK/ljUd+Q0m21hOvKsL7PWwOUqyRgOY7rLRg7hUG
XzYL257xR59MHkcIpWSyY14eefb9JCSrPMHwb8ZF8RB9z/GLjvp0l4GBr7UMVwf1
rrs+2bNIFJtK4mnWb6ba3Apskrc88WOqIyE3S1iKHvkZGz3T7IbVwK4Di5bXZeZ2
B1Mrv0braygK/wua/T+Bsr3aBGWJTrbGtfZuw3pFwJEzhU2FTOcYgeMd3cQgktjA
m1Fs4MiWSErXNDsLv7qnO2qLQm2ty8xOzbCNsYHIHWI8kAKoIHQonK8++X0iz8Y3
XyBLBXs4UlOHk9SBla5ho/tQY7lYWWM528jSSRMC7ob/1Sye3WM54zO+JC7VC5b+
I4zTsw+lZdKVsVSDr6VKLXFDln14od6cB0+rfyGT3gmzh1BBY145qiM6lGp5oIk5
cxlstXdhbXbf6rLgctV8RaiqFZYcaVtkZvsF1fHf7/2+ykwuBoBa+uDnBPc7C46j
c1mBF5qnMYFVg0EVo/MeVL/sARFkeJYwXH1j6rtSPCR9/lDbYIO1EWsZxLhIOUUW
ZLFgiqy/I1z/wfEC8vlrnLAmb3i56BdeunRA3NvOZJOSroPdYcTJXpjhUXb6irg1
Vo/UPbSzYc40DJAeuCR9IXa30jvDy2p0i5YbIOr0Ggqv8ScvYkcmoqj7Sa5AQprR
zrkbySt1sVuSIKt+p54al/9VP5xfJWgd5fWwAtGW/j1vl8Y/Ci4Nss/mwzEx0nf4
BqtaZ+1huQvcVcgKsUO87Yz3W4YGSI9swdLC+cclm5JFHMbqh0H3AtSJSYErPk0H
vvly4eE9f774yq4wjnvIyqYQlWFD3fiealLc7OAYSL2Tki8FgJljA1pk9tE/m3Ep
YjXzmSinDq/aPSgaf+jTJhz+l/tjO46L114WUgfxFvYnafGvJx8socNHBfXM8kTa
t5VYBw5rgZAfSb9ItPnzNRdDuMtEnC6PY3Gt5qbhMVrXs/JgTVOtc56+1Jej3ba2
kEjXVFGQRFa2nSm4V8lk0AX7mCAwJla48uyHWqItEaQMziebcFMC9vilP6UCBEEt
CmqqrHD3QoI+r0wca9JqczP8CWpV/Pr0U6btVqxBLi1H4au/dUvyTFV3nvMcfXHD
ShE2LPtE3j9Zrv0nzrryNzugUbszvVUaYEsM39rRstd4nnHKu3qAm6A1izYpbNsd
OL9dNDmpNqeNERXzWoperrvAaikCr3d+QnIDUI5ffhQbLmQOjOk22ygYLXuDxvdT
4c2CMyGunM8Is0P5SS8kQgvbpe1Gzil2wdNTnJikOW/uM3dQIv/RreRBczy+zoUl
ya+rTzxI9OcvKfVkYwrASqUFPJ4GZqI1N83XXtpgxB6GYyETAbsasZgL9O2IrQp/
tmUzLixn+tQdoRkOb44U6YkxerykBgdpAwj5mgnR/mP8crNOsxlXi6jKosdgu4MR
a5zSCx5DjJhPnglBsRWEhMRrUIkig8immlM0Fzto/WEmhd+xUQhRFjIuF/aKDiNA
cawuPGEplRISChuUBRMJxSmNQ1a9KeSakNuhM8jUh0zaz+exWhHt6WppvDwg8QpM
qC97vFb/GgXdyOVlu6ZfsMWwGNgDlgwd8ZlkOGBEg86IpVz7/KWZi0XNaPunm/wK
zMQN2Ffi2jmSUuj8jfRGOkCWASkf1XQW7Ug3Gf/tyJFlT01auynv4Yv1oZ85t+z/
LS3vV3jbivqNRj95BeTKxv+Vi67SABEq7DFKkSOIPpRFqApMd3khAPpev6ZwpEaY
eD8sog12X5mHMuqeFi+t0d+u+hcTf+1/3aacwsIGP8ECf6yPfk2mmodLRpdWajUs
5GJA1jzU4ke9FFrrKlcFm4K+JILh/SSe3OQTp+uvA1Iqr8bYTtoTzq9Dj2NxQdkT
xOXe2XlM+YBdi3YPdwBqIP0G9f9NH6XVNHtNupTNJshb0Eb2q1YNiBKARpPSAHbZ
lUV2gH7FfAerOV6zVnXmcGa9nS6bIULH6ckEeiJfS/j9NN4QDvV5L+LwCPmAhG/f
jgc0SerdSN3cQAPKVBaBLXxYit+5pzOz3/Sc/dpt6fajIa5G16ou57BzLzGJuDor
xy7a7ylcfRll+bjFH3NCZNP5hkneCUcw0G8BsjZlaKgGiLoreyVDHWjCma2oHwFD
ez1Oq9/aR05cPwdOp1FzeB02fRPHrjEFpVK7Hdtm+7WnYsPgX9Ei7CELU2JmbRZL
5Cc1SKi1wJ5Nb86TEJaNuLamvDTyuSWN/Tq+6ol0Uoz4xtY40UjfHevgErdpZf+z
5qXi1/1FRR5SvjlG7Y97nNIBdFpsIzbzp/T8FFSBv4vtNQMsJOWQqvvDGPmtbmoG
P0+xoInEqlrgYfCgPPXhtIZp5Bu+ThrPB9miJv8Uc5kBDWGkQcKL/oRyJAAD9T6g
QLrHTpdfIuz5qoXHRO4xH9M8JN42ZDHYgQpqIhzkHxwg2LjN0EAnAnCx2ZlBIaa8
xLGf2fBV4E5sOgiJz8jlGW2eqZBIW5t+zXwQLNzNTkQNDl/52N6mZ19yQl2bx4CG
BC+yv7d5mO01fjlcXW7sPVQe8YgcXzariOCNESnWBsNTK2g20fo8AA5HoSpOv0uR
6gLnuEDIiL8lTdsXco9IQo9qCa1n/hokPeFShSjcd9lB6A5JTkZ0v//ekgdXjJN5
IOSc762CCWOtP+OKN0nTrI/5P1vZAXvkbMVJS0xPlLKeL7ZK7GXv0Bjp2t4tmZaa
D8raEYR3/XPaAytUxBnXldW8rwgLlpvUUeZu1zGwp1m30a42mXuZY1HTpf/pmi8n
IvwXbThPRJRUXBfNxUEizy1hySCJqZqVmet+AB1kt0RKrvUHMrQDSFADk0nvCOkL
2Pa+T31UNnqPuwtyi3iL8j7+0KWXsu1Oec5t+6oqeML6tT7H+8VesrANKFfYYNy8
5aFeyRcfa/5dEAStmgF44F1evGlDSQv6C8L8jHqzZ2szURu/vYZ7fzR5WyWiW7jR
UOaom9GxydX6h2lvi0NG1do6hGwmnUt/OI4+4c2AmMULGhWmi6J7W+zcsnhdyuou
R2ZQshCr3/7MriRFT98DaMpALuFOOAUDHfLw/UkCkw1qQIwg0yve1upnuaOt/BaP
cGJBZ3eSO+iNCxJHEQaz0pxbAmD1iSwxtQ9Rum99om9JoYEx7+Kzxct7/ss/Y4W7
cbSLHYoXd/Zb9aQyn6cWccliF3abiQUKF2829tGleV0gg2wzkIm43J4GuIp/Rqdo
E0jBePRyzH0wS5N2fPaaX/FZ6z4BE3rCrDIF22BUx3H3kj8nrBGb1OYjVtiV0iC8
SqHLydRPIkOdIeMWkC270VzHyOpCXLfWz3NTp0Hg8nVLVAyKW95ol9PNpmERX2pF
JjTERO+Jq8FNBIU9MMpkUUess3uI0FkAfWbumcrxfrFCZFPS25OheVInYGOpTAEB
H3XPUbB510TwspYtRbp382oOCHM2u+cE3jDBLxj3eLPfTtHlra5SSu0z4gmeV1hq
9oDv5aQ+KQwXUn6XU08k6xhJy1VK7Vbs+RyuFipvYmWNnBvPQSHIktZkd83tja6e
kyG+NYvuBXjigRpzCjDnKv/iPfBDdw56Cq8GDsm61Nj+X4tqNoTekLo4OJ5qkjml
c2Hyd94/lABUhAmnhzwl/urw5NIzeB6cThw44IS47cuM5TWM0kQkj1XJHK3sVm7u
2G8QR/vWVGkX58xifZsAuV5QRE0R9WOuhusA0cpWMyuSM9FhIYLX/iZyPIB2oCim
Iz5FWPf2+PJ2K9WAIx5uOot/tFP9vj78Q3mKfVdDY6AZS1yTx+Js5iuD12tnRSSy
py/TfU0TTrcbzCoKhJjqlOOfcz7a3FsMIQoL7gGOh/g9rAOwZmZgPYfxXQ0PIPYN
kjorOu1CW66Kws/aOuLZZ5z4nyLyfxbCva2I/lvHzz3nN28c6OQNHMAmtpJZg7Jg
mCI2tuyoF8jYOqAOB84005JnJ2ixXZreGoWryHM6Z72TMNHN16+ux0SLt0XWmccL
uYY0avy4FCrmm6ujzlafB/TvFV4JzKnXQK5lLcY22PdCj1GN4wZg3ZIqe6bFexS5
Y19vAO7gXCMk1e9esib8A+UnMxoqDLehnyqOU+AokNEXSInGKvD+OwQH8fFTUt9e
UV8WlLSUOIe1QwDEMey39oKE+C6B50TQjmmOpMOZG5tTGrtSDXAY2paWF0dZQyWC
7iBuvKWF4BBrVEX9x7hj7nvDcqK/jh+9nbXcmJjuobCXvp9OXlvf45+LjQJBgfgU
2PDnecbaNAdGOFUfQdVeja3M0o0a+D1y7FnSZXnWRT3dX3noWwBpwFXrJiKkBM2w
/uyTRVukW7os1pKVuV1Wnrb61WQnDgRQ3U7SMzbwR0n0xKndujh+wRU8z9SFIzdC
R6PV6CvOvvIDprRPIjyEbocVUmp/LxZ+rK1/p46jigCZWqFNWPqz34v0G1M4AtMx
/K/Vds8tNdiNDyvot3RofP42bXx8rDEoZHn5i145xy24mTUFBsZ3OWDMSiILVnuw
ovsFq36qvskpHcWKq5Ao4i4zWPsht+rvglkQgjIDuOvWKPiGB1TpEDwW25x/++pJ
aLb3sYDoPRccZYU7Pb1O0VfCAUShhvZW99MzpXp1tFsF23Pn+IYS2fTqg49d0wVw
I1H4asYj/AoNkr+9wD/HxGj8Q/p0F+Q+HXXz8bRCXX7W/rVGGctoATzzdMSkGaCW
NtbV8AcqXBAJGzonxF3W+6hN5dn8Qda3PmYRlu8D44ig89kvaQqR2W3t1yg/el1V
tvvY4H955MrnrBehrsYLBFlyf1IUzTnoNTRvuYQcR4MXDc2Yoc35oX8roves5y+W
ggAALVltTDmDsVVDQiAj0h1LgFQ+IiVG4qWNoU40CDERsOornYbKokcWirugOfpl
jQ8kKIb74bp4T0lIzWSz1awGis3Fla++Iytjy4ifCXWTYyUPDZYDhvILVmmm172x
8ey1dJNhE8ZlTAEaQUEMtmqpdyRnzptUgku7vECwSIBjTLWcrBBg1Mvk3Ip4a2Az
5edrOdBdWyDepVb/twTI3lp2m8h8zyymQFA4BwWflv7snmwH2EqYXqBZOfHKSA1j
QHXuaoNw82huyvd6k1097woMO2OUHRRuBXQ99Li6YgoEk4YjOfcyTvrpsxMAFv7N
vWmEwqbsN4xHfoE9X9xr+vXX2seL8v4AESOrVjYdrlKmTrokMvkInNDbsvu+dTsf
7TWFQ/oEsyKTBzgo1p9QUkf1PR+Uv5pCbRpEa1oVzyUGWfAJojDUmd4KEHkIsvK1
M5Anky9cC5cUNuMMb5cmwi6jigtmGHpLmvc3R99T5twWu3sfa/IzWLoDsu8NREFf
AbwQ4M8ve9Hz7GlIATOC2333G0shbSuutkLBVfXWJd43o6gAzxNkDEMHXclF/snz
jCqnGlRuIQqVyyjoxSRpC5xmTBicOxJsfIU5cMoFNNBRBHHLWgCTrU7tICzuX2qv
p1Fi5cERz5QLJTbMY0gWFgMKaGUC6fKynjWZMMHaOw9w/g+4e7InicvFNXbZiSh+
HY/ByahFe7h9JzqVfU1QcjN3YgX4K0yC3LbV6VjbvZQGTJmOvYdc9ueIxhKRROX6
0+FSACiYz8V1yiGkyBltI2eQSZzh6h5MvgGKZDnconYi96H7F+y79Lo64uxzxoPa
kWXSVVRXK0ZrM+Mwm+7yAvW4L/v3gBXPAc4Zv78E3e/HfMw4a0jD+c6IH0D9cZb/
tNpd/vVJStH+Y0zrmTXpoz8uMefhvBcwcWgwJVDQf7fYaRQhA/LLjjlsT6oOsyXf
kCC9ZDxpt8sX0lkxy7U9pKyTP5wHWSHvVlnsH0teysNnO6x4RCl9pijRMuMwbkjV
3AFvl1KsvMLiN9g2aXFko+Ins4L2wbrRnA3aMR/5dbBiaRKIU7BgPyjkxFVn5Txn
lrH4TJc+sy8J3EFNpyjTnJEoiGfUx+nOO2kZYMoVJgl4H9IYvYoLG7565kGpwUWQ
+eQXzfGCLRvYtCeEJ0EwCoaax+wfDvTk3SuOsjERplsR3lqG4fIjc6y4plrghxnS
4xKB+YUDQXw1RCdDbkFxjRfxKElobR5G0kwstVZa1kv1WC66/CEvHJfJr4YnCHTv
f01YgoDNvytgbTzeQr1LS48/r1M/5hXTTStncSJ19apXbprKxFs6lr8BVqrnEivp
eW8rVlPnH5MaJbS135mvzDB3lcOrFeRN7GYFXT9/EOisWC04P4zeNLqoNNO/tDhM
qScxs/IKLW50Ve0K5SnRx+E109zUCVPiD+arFz9ctGh2f0cbDUC6bR6yt74Bp4Vw
allZ5mI88nIMjmregGrZUyoZ1Oa/qdinJssGyBcMEKF37HRCV8+3xRm3HHVcaN30
7sWTPyxoIcGYYH1dJHhjWpG/L4l0ChFAHfTImzSKke5nyQhmdAv1tmtcY6nMrKl8
m8Daipq8HBlk35Dj5IJykmn0+5Vs6lfjfWpDcPyd22Mzh//jdePx0xy4fcD1VSQi
BQQ01z2uFpfdAplGOZZImSpLO48lGK3bviYsmKFtqKX/zz7YTjcbl6WedsZHmNzo
ypY5hZbfPPU5cJqQj6NCd77p4/+l55hptRomd30uZt1G3a4vCWx+UIpvzTb1XKPw
R/jzINzNzP4J7v4jEEIOiblEHaYUdovH+O5tzeyex5dlgEgjYhxbsL17wVlROLq7
F/Zx3YnXETAyPMrV+PCNkjVzu8q7MbWB6EjI16Wxv3EDGO90jKRu1YAadqBtD0wM
R0dr2c5hMXKNIBABr3XrYsopM0pJf/mXyVjSggW2t7LAoCNB6I6nvWbX3PkfbSRY
TMe0YjJKTUpHN0SfRvrLZ6Ec6064ykYHlXiCcdvfFtnzEEzd3/oymQti9+e4PxDL
c42+oe6r6PO0VsYWcYFtkTPfry4T/SM1i6fBdu5+Qa/1KE5qDPdZZJbqtuui7vPw
O/eHgl2IHBjz1sVHcgW91O14eY48vY0nlwhwbUi8RZHC9LUs+PGLoU0B9vUacFsp
n6xvdM4OZp1JXbWq+ctnuSHq98pZHHKU90LJZwY1Hxil1Aj/BRUdD25Tnj6g+V1N
GmKukuhwOjUSaFXJpW/5vxzQ6/Hj8K/EBuFsMxnMhXZaxHupmJv23S4jeXdj1iZX
eU7Q5dyw3wPLYM4d/xHUtuoUyZlVnQ3vMU9w1EJFKSvItUGP8eXUvtKobAc6xlHA
HmSax/7OvjcP2INC+6GVlnKVstJsSLn5augtlSJFlHCvTNCPXCOnGfWmIhAWwTUT
q2r3iY/yB6Pvxe8MA8HV6c36qvVcAg7Oiq3DOx8OZAdbGIWP2ggK7lx462Qm4c0W
6d/03FyEO1FVngllWNFmEI/v4mNJPWYXt1A2Shlclwo3X68F6qyEOizLWDSX3bTk
dG+P1NLCi7Ne7WIACcH6mX66u34sV2aKk+qEA9NWv+DcjaONCtjupL1QiKVgOXi3
DWf1L2tpOBtKS1d9b8VFOqPxZItzuRvg7OoOnjzk1XmPfcQMxdlf5vLH3rf9R48e
h/DLtKL2iR0jByBOoWUEztpEa0IMIagyYZGOwZQOUpWb3w0EF4E2Venx8ca7cm8j
nZvpQTKJ4T7dyIQVjrxIrleAarzG2fdpRMoHP2pALIeVr/UwoQgXvZkTMC9bO0vb
Cqf2t02NvL/lxFtCZuDaw3oPxCYyCBhaoyXdRc3RnfxOwUhGGpBwc5G0q6lfB1kL
ecFm+Dzl34Mel6Hvw5fsxVzz08elHwAc7WCfcl6CAMJj+zR5UuRZwADsfZ3LeV8V
CkvANuZgCLHNCOCM0TRyzILUDuAaok4xQVbbw38rPmK8Wwgnz/w7X5kl1+aeU1Bu
uUHehPsqGFJ99WrMJFIQVZZtrx+vBlAC6SK3G4tg6nsb36UI8Lw2ENhENNFtvpRm
Ac7yyZYwgmZUrIkOtdI+I1xIrelO5qOedYhh3qPUyH74Z8xLe3hgAHv+LRc/ZdGJ
yu43KlM8C4xv2CIT2P+f92CiG7SycMsPVMsAHyc0TcFXzv7ifctUefWRD7cGtwji
WGKkVo9Hn9BwA0Dd+aKLpMDLfHXaBANP1nsg18FpAdPQ96IUNIHYTnK6/dJogSnS
BFP/B8e0iq+hVweLZK1Yb5S5++zcvUlM29yYI8bQ3mrkcTB1HxperfziMZZON/5Q
sXI69Lo2oziBw1sT5qsQRb5wXVBEXwooFR9OvLgMr2HrIGffU0VzWnMfB9CUcuF/
qbBgDkJ7VO4xbgCIGLJ34W4XyU4VXuiEu+mVFqKubbPQV1DBpAd/9+pK3cVxlISd
Kiz1qBoVaHpZ0FMcyju5cabiLTUmn1SZlEz9ER1KEsFVMgKH4C20irNnlyluGiGT
b78/eaW9BCWuqUUks5NwiwmSZCUFUhoWSg5GNT5fT0uB4cMqBaxK8+XQphNC2aRL
is/IqAqggfx5LY6dqkEiVGULRSVq7GrdyTRm9WoLSu9HR5BR09PFARydwvrsE4ra
1MYDm8vjKf60KgenbyA6OZwud/lZCew/yGMvWVlhtMeQxJ4AL99BQbhjlFHLvOQ3
+S7eJ3rl9TGYVHPq0AOY9Axp3d9LkewziKwZK5A8C5hkgapkgYbq2mGWrJSdZxYf
tPba/jqRcwzz288PWMToLQ3eRR9chtAcaP6D4zGC9uodwECKc1kh8A2yp59cPDIr
Ee70TQ1wvakLjovRlj6n4y029SxnH7RINbIsRT99iquZoH5X2g0FEdlkY1juxlUO
c2pzwFgOQTye0tebISprnk7eI8GEAkxC0RX6Q39ILaJiBFafekubAc/2Ox69RUTI
DmnjrtIzgL5h/UCT3D6/SLHaZAAzAZeMqJNRs96xQSE0jIsfnM7zTD1A06J4ji8x
+FuMj6Yrc3Vu0j3OYaMKjwFJmc+KTlAjp7Oz2CUtA/JMD1NNidiFfB5HLt3ehwqJ
sOg4q6QlZkDMCPMtrVEPu9mH5Mh8PLQ/MxUff6p3llAJSolrLEZdSr7Sjan6BwHw
bB+Hqk1VpwILSws9vRbfMsSJGYWn6FzVwi/bNHpcajuXqi5WZ+7yoz3OycTDaaOn
QDDqHknqun+v+VRRMqmM3tn4BY4bXkMJSsTszSYra1OclDk16W+Lo7r6AQ/fbXek
wZKH988od1ZFtnba0Zg26nqdCujN7oQaM7OO5Xsu/A3bdywaFKxGDpCSDPgDJWSP
1AVT9LxFXMZlwVYMjlcp48NmB8tu0ZDz+dbKK1OQ6WttFc/G6IOfMKAmoHgg8eNn
XwqvpjERkViYpTIDBFfqAp3Bg0622+tyKnIoaiFheNz+8/+RShYhdxC/7CTuQfa2
B4cZcBM9fUWjW4hZi1vfFHmHh1bbmVvMdM2Do+87KlRINuoX9tDfSoE6akNcLUUJ
nSQ109+NdYXGdAZ7wHrMwpYS3rSrxa+f6++zqqfqWvREkm9CnXVEr6ecN2f4/7TS
WXvvM4U+CpGScYaWJ13snPWllfJLqXQjEnxNkle6zwH6myhefaW2x8gYvbAH8tPK
o/6xX1TtRjoK5Va8q8k5yEyQTarBygrRKinPPZcEZSnGNTb4TBWH9posF8GvONgP
E7sgTCNqzjzlMRkXth+jEE6zD9FMlqzpskZ+Y+IqUr+0jqsClDCrWXyYWuQRkda5
2VrV0mSzXZRVDcHwQ5BIc9tIWnzsJCJ3+GA5uRza+rGPyNDjlFT6Vvirn8WuctHi
g42G3f3iyog2LQwpIa0oT3VHz9GCtgXHDIvfQTGElcJYJOj0zrxK+BBlv3WKzhiM
2jtXtHzf9kOjEvMIymNaRLDeiSD7jNPCSyaWxc7bD4B64o8nNmuvWDVoIvOSznkY
ZaeCqEWOx763RO3zbi952ohYgD2vwfV6DwASK3TZ3pQRLXtYBqn9FELVjKNUhzGz
1j8+eM5+Isb14m9hFqzPyfZGKTo+DYymeE7D+mRYGFX2n7THaUXTwDOIPcL5Yioj
cErThwr30uRqr5+aOqbX03y+PnLRmEar5uwIiUklIdaeY9GteatlEmhkqr09n5r1
ZMcGj7+6fXIv0LszhYayu2Z2kNDZOklNxTutuo+3FasmcppXN1e1M9R9dmBSaHOg
h67opgR2rtbtHYlm3XgRgC4w20ErjQw1fQfPK86VWv7m93RnXNcJvL7Dl83iW2t3
A1kWe7PSzYtLnobyJ+tLrpw+ZFsH/3LJSfepkP2kDkEDl6IoKr6GRAz55Tbf/iE9
P3MXJzcQgr4g76OP5Eh4hv1dLJlQJcaH2QHm2hZUbf+eGW6EJpSvAy+eOqMr1u4T
Canzwxm46O8s0eQZQsU3iwdb0hU+C3V5xt04sBYDp1HIcPE0eLaBe2TKLzeQpG+8
+DQdHBTq9Ged/4LdTmsbgLQruCxP6YaqtSQxyyhoLMKD0lICyI6FCqkIg0U71K83
BCAG9k89BTImI8dKnpQetMzqyA8i/Mh6lDIRrMPDK3zt4PXjnm2n964QnCWh94gg
+QHGcXaSZBx9y+5HNp736u7kt0AB2FweYf/xd95F/UFAKEH53pnuIC8A5wycV+en
ASkgEiYV7WBEJSwuQEQBHwdS9FK5GkCRhKh3QktDHgemva/RsR1yYNLC13uSPVt9
NfM1Sbn1XCrr8ZgXjcc9R4ARiNuj3+TB7VMkUkJT8SYsGnOpQ8PkM/aAHFyZFYqg
DxCvJhEQTFPIy5QCM8Q4E5TXy8T/pI9IXVkfzEetxoQ8HZxeuzXse3pHwTvsTGgf
wRJHfjMuLW4t6sV4YobNS/lZwoJ0KPoFCksT8wC8DGbBsje5KvTEwzlJ0KmW/f2f
lyOj1jGNH5BBoZIx2mr+WT7lfK3XHs1ATCjZSVXYQnmwPCFboup7zfsFq8lPfxzc
0luq4XeIHk1Tkdzb9i2QxEk5Q9RlROv9GWgzrbKNr5ImhhXRvUx4MYzOQOFf3EI/
ACQKNqyZ06HFIE8duFfGHPs/cBDkXhznfQ8LnJtZG3RyUOOMSmOGHzjlHw81EV7x
cnkhMXXmxWUQsMlMiwt/hOAfp6ic/rd7jI7hslWxpu5C5uy+YRplv/qSLkzjo9GO
63LKe8D439YeoIhwRya3TOek1NT7VL0wgJK3jD3y9bwxt3J5g2VSrFGgTQBLTxe2
DkcVofRUJKSsrJJYru87VLgNT0SLh7umNPg1qSJmZ8kfh6/GeLhIIQM/bURu1tWW
azl2w9vvxF/aYMQLiVbwoRkka7ScXVaQePqPwfoXsAms1OfT0AbcTEg0Y7R/spcD
eegPCutWPgvQmjz8ZM7QyhTij2EmQboqlFm9IocQ/6dKI1ed1VjL3OoVuLYbrY5+
1lOVXLIwz3ifj83GX0QxFbU/XjuSrqW/isEj/4n53SmeiCeIbY2Ji29UHfjzvCW3
jG4S3ztV6jZkNSNs8DcckEvGJXTr1jc6sf3O06Q/xfum0mW6nLfbP6C8LVjtRbK9
UpUqcAGQTPcijb4K0ZExvmWkAY/M3/j2zdAxpxyDQilmg98GlRxr3+pH/+aZ1sbP
ritrfLvNudBcSP+UIEawfa1KAC5psf+GL0jTp2kk31hUUX93Z0HP+E+nN8HsmFXW
raSUutiaSY0/8JV8fYfjThQ8S2bsIpnaJU1MsMk+K+pqtUdNWm2FMoEVJ8XKlf1j
NCRaoli1Mt+uNcB/2KMnnji0GB0EQLzeWqXllpV63WBCWZYPf9XYOOwJ1eqNHtwq
q/bwYFsezFwLb/jqLbfXg1t5MLpFQSgAFFj6B69Ht5tKNzcqZ7TPLfar39N1rc3j
2X1enNwHjmq0mb3EI3bhH1nj+gYUZXPjjzEfAEu45GaUnlHwgB+H581cc1Q7abcV
y6k6q0u8CE36+qgdvBSZaOt8T9Hpg/rxp9ctV85HIjpUEfLyinaDy/yL563Pk/MV
/6QmosVF8sOtNczzncL7w665fbCU6RBqDpzJuFU6VYRxD26Y3W4Hvck+tjkhLWSK
ZWgyHjX41RqVfmpORS7yjndRfDdmifUGAcUerN3+ECVVVw3g3EDu17sjwwkZHE+1
wierTHF+53i3mCMmxhOr0fNUQdNB06QPU1f8lHZ3v5MVogN0DNW47gqVmLlvHbbZ
gSQlwg1Twy+bJOszmzIlalbJCgAxPFHW/xAHKguvdWQOyj9CyGluH2oZXiJ2/D77
6PIL40Bb/otTN1Acka8uziwfIQPoEsC/qS7ZcWaUFBZMB9Uaqb+Y05nieW+zU03j
UtBmtw0pSwO9Jz7a+T3sXGwGnDEMkh2UKR4GAkwpm0Aqgvw1l8ienLIYATLvpFC1
iV9XJEhZtVtLBmNPEyBGAsel0nd9vw6xXyMc3Tkk5Dpr12XSLr0Xsg7ygV5Qsm8M
5xyImE0WPeG7LX77+ZrrZH1DNhM0p495bs/g/TxJPkkKQSnNerYPchRhSQ/4aRzK
haFmFh0fantmp+xOLdRZw3D6f6bXsTg/MX943Kjkqm8+p8EjPESWDrErGp9ZvcJ4
sSghqdcWS9MZglm6pfDK8oA98YhMBP+vOso2AC1lHrmYTc4mbpx0DZdQs09Yo91z
1zPMX0ctAvD0Qh3UVUP5XHRLXiotQdJUBcL6eNWhqSnDfUavds060g5g+zonwKAS
zHZexJ4d8hwpMhT3LP2WLU8l446h0lPN8yCBgPJaDuyGKvA1ES2IgvGa7aGpn160
3VM3qrG8ilEsu5jEHdD/bCj3mbxMzo2U5xF76xyXcn424d4qskBQxlM0XPZ0UQDH
7oyakPiqwXlROPbQgQfZotkR6IuhYbu2MROUbADgMiQimEEbgWoTubNo5070CG2J
RfO9GwGVfP5y/9mlLN6Qr+0Q78sUZGpJtQP2fWxHy5pQ9FHz6aTPr/+XMMtEZFcF
46L3B5YmZHLCnigwlv+6hLfxwU2Sj6he6lbt+Fi8S7jWUm8c+Zq9uBZ0mSZHHkB2
VKQSziJWF0jroW/D4sAaqigKLxaAw2HMy2y6tV2sO+hWASfSD0WBqdPpDzdml83v
bORPl9unx7ixHzgI7cvzAzayWWmuA9GSEfPBY+VZWCx6D53vG8u8PFowQKnKPyqI
8QaoKp26qZBUcwK6bjyOOEMu5ReRuDtJyJGQWOhHHe72nL4INf5Y4QrnaH53rBtf
tbvVXq+YIgDY2Ec8Mo4rQNnAb1OS3e9pdzYoXZfqfVyVICA6roEW0XJ97PS893x/
VMuWqVKea9lo/UGvFLjqu95+qjBbvpBKjEluzIMkpXcj4v2sE1fAWvJhy7Jgkjj7
+UwgW/99uClty4UxgYmRiYgJklhJ4kH1dKv9jXu8DTKY+8icRjWw7RRBaDxPaL1C
8dFmOUYSb2jkn15W1GO2EQe5NIZfD2usJJgyWhd1J4+Q+NmRBw983QihaR+tSqf7
Kj88gl14IQiU61Y58oriO8XSXsDUQ63zb0ca4To9xKQCfy5XRrPzpGTGL1urxAX/
YvATEpS9eIL0dfR2Uaw9x+di2AdGHqS8rtvLzC5FDj9NFDzzuuNBdM+9oMaE0Raz
em3RguqaM20IpSa8z68gJJNEQWIDFIicHHdNeuRLTul+xS5zI8f9YNtjt3wePbev
NuneOMILZXZGtc3pDMsdq5KpybT0FDtsH9LFMsUMa0lLI/xRumhzucSHMuHF4tpa
ZykSP7TxW9HnGsh3BPmsCeUgnXaNoj0L+OQg+JGxcy/8wYm05PGHk8twSUxRu1H9
6JSCFsXD4jqBltg8qWK6J6Jb3UeURecv1X138MJqf3NaxWFbRxP0bvFbSlKzMYDB
JhJAypp3zSoizuOndvkztDrepJUfDNdozLiXaYNp46KgoKq0EeROOO+BUV1sKMp7
O55hBvd6XIxLZtZnb8rPWvI0a+XZ4YkfdBOVEBn/qoQzxlzG5dZfqArvQOhHY+54
37YfT48TIw6dyyUYVex6lv9Emc1dqdqinBgjIdfARmbuNodR/NEQvlGddLPUZajM
ZSZQw3smU35Jo73afbUYN3N/yMjaJdMIOjfiFJgfl0AQMnfWCkzfYe9AHvbdStr7
i58KxD3DLh8bSPhyyD47PMGu2iiE4reWsdgmEvU62zuVcB+I3XZ9iLyLWOKBRV//
yyFAvNb/kb13OoAxmY+igrhgl5cRXqqVl3kaZLOKI3fE8HmmcaoPg8gwrcbG/w2X
PJ5IjfIYV7bnY1m4TgYh9lUhcMGHEAXFu54Z3gNT+YgmjRebB/pkXsuvE7JxUPTq
R5wIhS8eYF/W//sWSMp67MACS9iJzQCE1JX+A8pt72H+9iYxi02nbhEu1sKUPk8u
hxQYqCIMnA5zL4p5NdvPKA6919c/+syJLsY3QnnToXeA687BZ3KvYwIIlIdXR4Gl
kytdHnYWbyYNGTi1ppZZ00PddhsGmh+M0GtZBZDtVDCdlgRbvzYIuGdaH5H9XCaf
GAb1fX2ikUNKoHdm/ob/U93Um4IJ8a6Qhsnpc5+bQ9CTq+LiP/Jc4QNW89lAwokr
qu/mAXybXppsygDXEh0HCt6Ret8Gwe7U9GaZBQeFztPItwTkuskly24AOcwEqX60
AJf5XLxnaNQCRHUi5vBjcCVFXlELoZU2qQQe6lPmIzOax9OTbMXUH/Onyjbv8iOs
cPzvKFE7XGmZQf0qHF/SLWWzGUBBiUa+qXXxh8g6H5/GThuzUdW8LGmdBx6kdcFL
aGNdhuFv7m10VAXfXmL7GqCydv619isAz4z7WaDNRdEFGezBs1qmhIMgLxPHMKe5
PmpLcepaGOrQiQG080rA/rzG/Whzr8FsXgF/4zlb2wHug2LYV0XWCxbgGH+Z0Ruv
lR5uxZ+nT+O+jkoos18Y3i+1RG215D2NMgKZhpkESB6sKJeAW8cBiRE33myLk1vx
FP1cOkcBf10P3kn7OCXU9bwyty9x147BBGD0vMJgIyxLin3dI+imInlwhb7UOtAt
Tt3K96R95i58Xv1EFPUxyaM2ISLWhfZ8Z30U4CxziMJdAsNcDm+dCzCmhi50l9Qb
y8haoEJcfeHrnGKFKxg5CBdvMh0pJbLgbHMbiqSo2JZ/HwE9m3+8uSivnRD7qOnx
PJhR+SBEmibQ0r86unhi35siplFqinmngV6vIqX/ikPkuMoE+AyGSmzbk3wSvR8V
oXbaukrk9wJ9GGNkgVYedja2NmP5hHinju3h97Auu29xB/gImrPaF3ihaq3Tq/QY
3TrHF8rRzChzt/6nvLiulVxn3ysEOA5mmzxTq/zWvksA/WTSXn7Gk3K7q8ekiAj1
pjI4lRbt92yfknI85oJoVG11qr7qOFog/su6ME/TrtsLU1bUZQNneSUSk29rjnNx
49QDK3zh3XPiVfFsX0i3qeXp6c4ioXr49maw49gbBrxiQp+5fkk00KnGFYGZd0Oc
+wNqbM8hYgvtjdzH21RhyxeaTlSQVi4fdKVVHzVuO/28Pcq1J8YRQD916qYnosvt
7A2+Hbw1S9bjJ1iI1xEL0rntPYKNEHzWBqOVTtxck5g0fRQ7SsEiUPA2YBp3IyDb
43rWOQ52A5dDd0dgayduOS+RwoSJQnNO7LitCN8D/yi7YkmUelb/jYsQCWkReoTD
b0y7qE9ZTp2tedyTGe+haYLgOPHU9A66bPZReXhJoLrFV3vvmMOB2GXQ+i0it/qp
D6kNzgE0UuVA8dZE3AjW7WCcRzpVOq70y4P3Q8MS4TFQ4AyaU3G/Y48WiqFcwo3c
V7gc/r3/b7KuueqyKdCYJgsQtrBJRF0mUS2NfZwzPplIgFBI31oa3Ce3PQFlcuix
k+fotme+ZIvK3HCfShrSqSWGmeqzSkmdCmqkQdyK2X3ZYoXQ9wnCLkKxZxhyRf+Z
Swu4B1WQRGA+lOSFAQlNtUEc1jzUphn5Euqiz1XestA6nkkiuR4LCXTB4JivajFi
RlRN2nVXvdPK3LQAQ87wYlS0uHbvPIJPjtubbWCZQU/l8efFdMjRoXLcPOkTz0qk
CWFWedlaBb5JsZccPKULJ2hX4GPJ/3JbgkSIRC1IoZOwVMbAuu/0xs+Dcpum2/YL
dDEjUa6T1XeG+264K/CaVyzPf/OXpvps2UuBqTKdObUWPXGfWQ1rEFsROB7JE93C
twNrkek/D7HAweVX/sOYjw+Q2D1bjLJZbV52bS9+yhc88IUoZy7Pl+UpChMFu/Qr
XUkZ78g/UwPoPM4mqK4CgSqJZT1axx94+klLTbnJZya38SlRZGAasqsDFdg0XDJX
0PJ1JEEsr0QHlXzcv9M5d0tKnvB2ppDAHm4WlAKuJWD6Fh74H1Gx9OBXOea7P47Z
2cKu1Rr6iDjrTJ5jrrQeuElSQym26RdOeZ4rCWxMfB0rVQvstbj8jxSWZmmVnYTT
FinjF7iqIng3ew9ba6y7J/xLigMA+4TAu11tYyVay1Oi6ztmEUqhjfPAPTcZu1iP
lCEdgK2bn3TJdrjrzEX34fRBs2fU5yuSf3wg3c7vyOyVb+zFEvZ5U/KhH4Ajn+tM
s2Iax1s/UyhXM9C0/M8XG/Bpd3I65WZQyMfZwwNxfKZaTTmFst7qxvvxoy4KT53c
bbg47GLJMcw9d9HMxAxW8bMEASDb/Pkst5XJ5P5HcgJWHgjgOuvTibK1p8YAeTaV
bm63jiV0TDCPzFsJEqfy84l+GYRBc1xC0B7/b9rEvSXqvIKxiaJen9+V/VFBSHWW
UkVNKaZwhRIyLAyeuzd4P/KJtwLHrKG/62UxE5jYook2u/GcWBwKPh410y29afHS
mSOYJW6Alu8xzcdfp51Tnuc6jWAZC+L1QQYAVnIc7bXHv6IrcGo0OVzp0k3PZEPA
iOl6fQy8R4BtLXeEsEttNqCp4FShG6AUqIBuJ8r+GFfvAoCggrnUHXHl65ESusF3
a115XpJPim1Xqp83bL8MhxbSK7VlkxTqFJsnuQtuEGqA6rQMZwz6AdPk6sYc7U0d
i/58abr4JJNcSQd826mQGKKgEcO02hQpMEvv3LjsaKFRRUloYDbpxMUcfSfqMI4+
E1n9wH4upckXQu49el8WlvPUV8jer390Y+aTQjBxuOP1/iCKWFiVaYURfMEWEMyU
73s778CT1MwX70M9F5K5InutHa5obIYQoCGDUccnBuhoZsXkKsyUboUgyD0xAXlm
XIVbn/L6BTjr8QWzZ1E4rJnJzHbEOyHfGYcsEexJ7jVScaJy7vmtzENoOvWGqGRR
9RP5M/kcfbpQenCnNqMCe15Gq8TqUV4w+eFxmxCdTkaQSLKnETScjLIAEEGt5TFi
n1GQa69nPPEb0fHeauXRe99+rZJT20l7qT15MNk84CFv1KCFL7X//lEtlbf5Y7Ld
IV2g0BOpNdV8/kIlbMk8CysaEOIWmO1QJSPFxS5aA54XC6q64iRQmnkeaCZoJLLp
2j1ovaOQdGzUb4FqErQmesYQqgLK+Ea6P1QSxhpKZ1d9YooEHmj0f9Jn2l7MNlSE
UwKh+cDpLLAtOGEpSB+GNRShZySVnmkiRo5kvtAZf4RtQN478KwnDM/9WKZKt1gT
n6vrMhNIck2S8VdyeaikxTQd+MCkW2VMs4vO4bYEm7tb9q2Ce9O6D/tjon80vAbn
56a5lmjV1x32QIxaijE4KFtzN1WoQjQS1FTklF1QACGYx1fZmyiXtWvOJDk1hZmz
nFYcjz25LOf1Wk/BfhXvJKKnWbyw+qU4sEUsinOfmWsXPmAqDpWlq/F/Jzl+OIJM
mea34ZTKeUwIUajjYb3cpjyGiSlclOvM/60IK/7kS7iE4vQECg2ifZqePffxnDmM
eWctaSBmzRa/VENBBkCpuSZpyotE/QES4DIcCNt2MSWu0wcO81lwVhBqLaEGWGYT
I8Q3b/qbNbKxzHuJfITXTa0GWS2pxOoPgsvfFK03is/QsQb99lWdbXvR3ni1kEG3
Edtwf2BF0WPPdVj0t2xcjRRk9dU0pd53V+5oS1POGHNlThHRLwcl33JT3Ca9m76b
RTHf5q5HAf2Utbjr1GXVMfaYf0txr5ZD454sEy/uA7mzXrrPFsOefNZjjVxGaycg
32bg4FvIbFQtiBgeEkmkJa8F85Qr+MxYH5jOFmD+vGG2SExyBWZt+nYUqnAeH1YS
iATZIhNqLjJAyIOhvvAyASfVBHPFOjj1OcuNvyWLuO5GwsgI4ts4SYV8cmrlXh4q
n6TVxOJWjsMbAVowekIoR8iaeSCiRGfIgnYMoHVRCxTnXdnEON6Y3JvTTcB9qm0A
AV9mlr4dCdKfplHIGswwAGEP8YhK7COOditYcNRXzum+4EGJ5ts6ZBAhWKUp7CN4
blQBPxltiyHWcBCAhVzruO0Hpob5oeYWYATJ9jgoZUkfN08sP/KY4PtvHirH6EMq
pMTs15bZRot+/Q/HGjGo1oEbbBDzJ22uNPWjBfbRTn1gZ/RflPoyq+uWPr39Ga0I
qEM+LhQPo8DosGalSNHJ/m/dt5A/tdYQaE7g3Sll8aPsIZw7L7wqTF7TfhyDx+nI
LrQ6nAd/+vEW+arCUGtQRbw3J0T3gPS7RUchdlO0NpfoO64nK6gLRP+uN9sLql4q
VtQNxXNCD+u0Y9VzAmBsrqrs5daXr8V2vtUDmrUewozCOfQRohgQEuju9PE6aoL/
afupwYkVT96hqx0Jz6MRSkULKFhul4QQiKI92tiQr+zc/r16iGPLfsroKMSkKyTS
qhz/ZogMdEAqixFupzE29+YFjnQa5Q+TElMNS2Xz/L3FDof8Qe3TLdhMjgtYkJEC
I0+4ef+cAslUivdf7Nn1iaVfovleLbs63M1vNfFpUaJJBjH5Hubqt8fzUNCEKKdw
fL/8uuEjmBrPkd1u+hpcMlbahafvhYjoKoUGPhibwLRpDZp9XwpWisOchcP8260r
m4WG16K7iacFFlkCbzpYZYsw45smlnDkW8jZgsnEa5ox3tDKKjiWR6QELMhGukSX
iuvxIYy2WOK6vf6GFxcePWQk5qq867ag6HE8T5Gyu/xM45OgjuJhRKtPnVAbyPnS
hwIpw+b+2vDT22/zPF6CQ4iB4MJA91cpqpyx1CGCQUZPLPQl6FixuAI2DWsqnKCd
lFmfqU2mqx3JuusLliILOQz6VUGkoLP1OtEjBRXuugS4eSeDRy7VcYRiAolD5mdu
QEumRk4yDySI1CvKBSM9iRd56hxwG4d09OsGx+i9dVtlYRqHnVTfNJrYQHlOCGGy
9yckLs+v5GdAVoredHn4uEqpOQAFtBn6Nx//2Fn11sY558xzqE5xWZnyGlVrd4y9
fOzFFjOUYTbwEo1XE/mKpO8G5STv31+jt6uJGV5/qRo0LQ+9ClAJrKhID5nBYEPy
5FNre/ifAF3P8L2UvZ0pQCoVaZW2Rn5i74hNv0//45d2FVuC8yIi9hQ1jcw1y6g5
/lQpVzBvwxkn2teOJUXT11cQ6Gs9bWxGI5wszA9yZqCIepgR6Yp35sTzD5Vv1wg4
Er27dLdLsG2oarLpPle8oWwRzcoadPMADqT/iuDnrgS3wIOrvyBbsQaAKFind8ok
UJua0tLzHM+HO25SJiW9HFNx8oYsvVkh0gReDH49z8mFRHADYklSW3W2oStlE361
jBdSM0fHAW60nnMm9I3nHs/TjbldBoqfx5ZJt5BKQCo4rGyPa/aEKODcwQZJFWZ5
alcWY6J2rFCGQkmDaI/OkQFzFNdOkTFQ0olNM7ICqKwOo9j/ES5sfNP49T4rJLmH
XO2xGwy7bjkY0sW94eoTQryrclgPAF46ayJJX6HlN6h6ynUr9bG/My4Xr1Jo6Ukv
8SeTqqxN2LS1xcBb+0rtQZf47Y233S+HrBx/VbQhV3FdQtOJKTtzNLUgA8vt4MrB
eJ/trWX4kVYEaeUV88RYxUJn5MpRF0hnr8TeadiYu2/5DX2KI42/eZxQkPw0Kbqu
rgF4IFWNp5SxTuGUbTUVfFktpixb6K3X93rPgkbU7BFhfpQsJWBamXNVPMmUk7Iq
Q9d9/GC0QYJni37uJBHY1sIqJIJt4+13PnJgrEuQ5fRlL+fHvkkalNMo1F1cYyBl
kFrq5iBQCBTeJQAQ4Z8arm5jWie3TLfl5SoGATlXz8HHiV5eX1BFkSCO1zZOtc8x
Wc15rtORLHyrIZUfcpRMwB0XIW8u+8wtpT4gv1CrgPnTSLVRwbm9NhI4739gPcQ+
9mWbTMyx8cjsAYUd/NvENhr319YXMUsMvCNZw9+mVHTzhkM9DCjtYGWWk7rOgNPh
DQKphwshs/Kw4xo5nrJI64nnmwS6l9xE3CR8r7ANpAMDOB5/CWirAIVe7oYMkMey
7lGVEaL/F1lSgy8B86TkSpOz93WZwNQZXRk3Qqr89OqJEfTchZH8hYozZWLFlORL
1piuhZYjNS80gQNP4SlhFwpOBhLf3rblCMmWSkQkmWY8F7cjLNuWVcwwVDUJjAco
CUyNpLjJC/O/psyJRTiexAEQqWp4kGSMgk1gf7P/OMeabijGRThFQN6d+fpYFaax
+GS3SGJkqD7KY4rgQbLcFLI+4r7HpnZlfrBp8qYz9mld+MxIAGEY5PDK/5XdElAi
kOfHoDx6qk8YHIQVpsjkQO7r5n0WJmwMfU97xz8yrwQEN5MMLf5Ff1lDwWNTiBND
6zXZaP95aKtlI/kc8HDu2PvOr1r581RfqE69oeO02Tsa7oHhBvfIzpXmgOweYciK
ZmnwzNTkuA0e9Shs/KY9Mgcjqcad856CPiW1Gv1WWEovyvFhFr568m4qAbNma6fv
oPsU2nDccAOr44xiFAjo5kTZ5DEu2ZJMAc95GNTflHFwaAqBydSdydcfXGky+j4l
63EdIzRk0ZzOkoByEpQPCI9xcGAlm8Nkz/lP3zfidSwJNW873wV1/tCpZU6wEsDL
G+8V1ogpwl8LbSHjxettoeKWUGI6rDKC6Aobi23KxuXbHCk97XWtxPbRHxWVKBzy
eR+Kuts6CyVEPyQ1TX69Or4VJ0Rzgo1QoITDk3XyBVAuVd+0JvGEZ3p1V5N5JGxt
2OgzutZPu0vcd2pCQ6rjNW6oiHaG/5DTe97xjOgEoA7ww5iz8cbnMYXr8fabRQYT
gIovT7WTQwREX8ZCSXWClsEVuQSTliVP4ezBPrEN5i7pU1wYZh8VlXLGeV+Awg1C
AIT1c7HpmfzLA8FGYR1Nf1NfeG8xd1D3yOLI3/DKN7IsfqZijvjN1Ez1ncMWdB+8
RR63YGonNS9SB2ymnRnjybHXMoShZ7NFify1DmLyMJbFxFmk52vsWOwY7ztNsVE4
3L1gUrRTbLCS/5mHBrxAHDcpiKzCCmiebod0tf9Zspsc+lbUvb1d/RSF9OfXMsaE
rrH/sxo0YEfnQZsjUjphhz5TkQYAoQLT2YvQC0VcMt0gcVjs4kOReGPC6kSSPrHb
OpqTTyqetl1HZTmxin4hY48eeqKRbNOCdT9ZxpDDIU75CSJYf8S0uVsLpYA2exgV
ALCnITidUWsWxZTh5Tf77G1Ui6QfcQjCZdNBiTVUzuw7x3nHCloATqqu9BvbfZje
LEbyzC7TtIj7RMa9s8fUVjaCxe2u9KUzwhOKEjQnDyjKnJz6weQgBdMZH/3G3Lax
GCFEKlyXPdKtpT64OCemh95+7HDf9ENHwqfgkwrWyOFl8HO0K+JXAVUazwVWeOpd
z7Iy6TVZ/647sTtsyZ0ZwJBCF7reoXfYbS7u2MAlAxXf5syyU26j1TLyWjenTcTA
b/H2DnXUnzFNgbAP20ABNR0Gg04B8hLWvEiniTalrh2VJhxEX8abj0YDgkWhAeTp
TihtqG3KpGhorZIZYNHMAjEKChUOmi5ttzyF0SJnWacLVwjl9eFZFp1d1k11GEzE
U+bLO8Zy/Mzmb/8zKbbcF52Gx7xAktO/uawsry078NOn4Llml7imublnanvAvgHC
R2ys11sZfWZX2lEg+JgSsV/rR2g1NYixfIt512uNnbHUKPVmN9NSUd0q1bY/F+9I
Ba6fhkdI/l6ihjmtGl6d6UhonatLC+YOfSRsy6qks1Xxq5debA0P3TYW2duN27Fv
8xcW7kJ3WIz1IVYwETFNtaQm14eVUEtPxlpZBVP+j0uvYb4q+VuiyudcQ6VQFUsv
nT05+mMWJm7aj454QxlhR7VIllQXbCFSuKZrLeMGBdLl2plbJawFHgReg3oXT42G
9J3FObMgew68dHlQJ6hCw53IO5U1HueWO+3G9cg8XehJReMkgc2s1sUp8J1q6LJa
yt5im23lEBD7evcZq0FhPuoqR0/bKssM0wVFCQsun+j388TgWE7xJmz8zOwEsDlw
aqGrMzaIawEQCl0YkRCYZU4zVt7Ww7JQtmKJYh5qYsrMjPXY5BlhCejn8PvMsmpJ
FJTCLnvHxQPegv8PjeXOA+p8eIgXc37i/GXwR+YFTTGLwt3MoJIrhiTaefa1ZYNf
V3ZW5SShL4LBYgIHv9mCfLT0Wys2eGxruwmV0/jvBTU4CoY1gNFvLYg6ZbZqAEK5
CQFF9guDfmc6AEySwoFi+Y/Ezo2UBMLlXImOobWhwhJFzVJdDr9ZkcJpfa1GylMz
35SvmrVhOB9iC8uEHXFHh+ll0mbC2/zL9XC7WvE+UZ8x8rA4uJP+08XExXgnAAkR
wCKmTz+ulnc4MeaPnRGFxhYhcbhU1VAWGXT31JSP9g4oSu11BByWZ80doaIUv1KN
uPfpQFixYQZId8LwTNDOMEBh5P0yQYgfnCSyDw43FyRo6O5ftq0c/meTUBYx+ift
VjrLeINLRG/uzmfScDfu3L/5PXvCqp6O7AlhBzFqoLX57HDQQ71AyUWUhA5ZLKr9
4f5BDgTc6JqtlkmD3KLEtIBgraMiEFs4NeTBWDquaBamyYYKOqlwvhe56bzFrK99
/UMO5wVPcKrhjDeEo4M0OhFcvoEOqJmlg5OaXe2YVVmY8s4Ne7qzk8jDJLp3aMz2
6X+KkAnh4xD1S3j2DkNRlnK+O/VeAdMpZyADZFJwl1MfR8YT5p/vHxKI8iuI87sA
HzSMR34h6ems8YrughK6hnNjXsCipVDHS2lyLhG6B5xSfrN0A1AX/PC5h+UsrZen
FtG8u3klkBwkrGQxe5I2Nb8W7EmVRFIgyiSfRafEDn5Dsd4S8Ot2/hVFhR/eu5/1
CBtJ+Fgt7/EFqvwRCB54e8d2a0gqv/LKVUU/nWoYsb6XRPkrpq51+098u/L0LeGl
TJIBlCqq3h95nPOYi547n/zv2rOxOJnKm/b0qj26Dhpk2yDJsZmPlr3gEwWg6P6a
gRYri5wxW1b/fPDCxyl5GptT07TWJNlHmKg/96Bk+Hi0KmcSnJT/hpkgFy37BdNX
rbEscJj0dADXSztKUXC6lPih4MONQ4q9HZdBBvhr59MW2CSNj3uIhrLJLaGioO9r
ReLQ6PhD60SblI8/idcNDUx/pmnD32FZo/yxyajRBpXBCrgZA2+8yE6LZHwDPKDP
j6nS02XBgle8h3TSOj/xN6atyRtfdCTkwv9m4EXc/YYaPIrdOXpUBQKwZj5n9lrq
2QLpft5AwKY3xUuKuypy6E5cklFz3ap1m9ocZYcggW4lvWFH2mfWengu9n8q6ngo
WhpxXOl30KEEPNaKewlngTTHketNumbNSuc/N0dBGrRPqf65k6ioUruNv7sutvxJ
H2UHI8H7BzZBOAtm7KVhZuISgoR8BpIXEC7M//MG2cPrr4rNK1wzBfh7HNw8Imrb
UhZQMd8ZwNBsqXKDsTljtIBl82CqlAD86/P9upoqgR0STbyL/IfY5W+Ao8Vb0o3c
Smu49J5BEDGTNqj/0/R3dwLSBJYqD74yPM6Z+kufJ0QsGieqC7/xQ7X5v99Xjmdr
c1MAPqGpqE3Vs4tVHuwK826sIfeMTqapJKWjCHmP/gsiPsYb/Dw4Nr4JSIeDahCZ
7gcVO2BouGRzQDXMbPkKUjtf0hWkAzoq8KKkkrW9nBCi/DDYn2FiTUY2eWZ7tiOg
YuXVuX2gDkXeCabbEwvu0cUKN0kO0cFJI8sGadJNVzjSBuGTw/7YjrB0HXv1Vcwj
kJSc2pQ1Dx+2rpuq9X122jL9CwNbYCTkUSLMl4KHbMeUdnRx9+oe6lcHQk/0aalx
OpaE53rCmvH+bYf359sgN4l9wCN4uBeIQpj5y9ndsJX553oxDqporM0ThcFJQKB/
wbBqNrRBD27PtCeTcfoWQHN6LvWIYQJfOCG5ZEVK/57C5cpGW6fak9VznYJPqr8C
cu8/4Hw/Nh9D2IIigi92Yiv7WwwA17W81C3Ay8BcTylRrz2AZxVwAy6AFYcZVkND
KkK8Az5fWhGA/wmEeA/jOfzma6qkrQykjw66fY2cVJnPzlZbAHqhsQ92PykRP83Q
NX+urpiLlNZkt34C2DIkHlHYleuK4ZTr0UYo8Db66jwQYCY5smWAcz/pVKDjKN1o
jroiNbF1QSfQJ4ozDtaLpLX20KPWlCkMRaYOgZCgm7+mb6BG3vs2avM0O0KGXhVb
v6lNGVtdgcB1IcbPFWrVxGf7mQsuPQmjrGR6COJfIfN14XqbSCj06qdxM1Ffj19S
wEdsa35k0WPO9Xyoubr8UTGcdn5/PjVSQTkEUTNDZKIJoXxw1qqmDWchk/FiouyK
enYwJEGFHQbe58Uyaltfbq2EqJGbW6J2Zaf6P/+cN5190pkP7ct4WciN7CM/iXpR
9d3m5qZz89arLEDWh6+xioPaqRN2Q8DZ7Yld5lm0Zy+kortU80e9Vz+LawAr4FCk
mbggYjjD2Bc5Hb8cRynTdYrHSL4uHlshLg4XczezRCS6etlJkS3IvvwaZLeRqAT4
+17zqtW8gBBSmsAcr+8ZHvElaS5yxEzguAL7QIWXfIbnjNhuXG1eePQiG2/eoXWz
cDfex1K74AWvqs4NQrhSVgjomcyBJ2cIiqQYiDxAmMoBLHhZ0PYx0bCey66q1YKU
fDp6yTv7N/EI/wTdX7FN9XW8hYPAKm6lEhvICvtbPrDOHbTBKDWhcBGLQyIxUDVk
nvrF/QUEFM7OWHeq+zSN28KNmMD9WJWKtXQ2+/M36bT98M/KD9J9lv95YB9YjY6o
JI9P1Xx4QJe51kdyjh0b7VRDjgl+vRlidT/m5/eXUn/UKM7E8J9NkZOJbai/L9f2
2Z9f0Xv4L9LObCIlv1nUm7mEhnjv1OcV2UPgMDgg/Q6pA8t9VKJCfuNZfu98UV+C
vTKoxmxpXkuQ1epnUkVHh+1KIbf7JPySG0uwTcTMR9lBnrytTrjgRFP4PUdtL3OQ
gixuQxFRUAe5hQo35cvYuUQTdbtX6wrRnQ0Cat4qVDoNp8OpsoyyROPs/6oivJMp
oO34uR+Y5CRKnnXXBx4ueOj8+mClL5nLFJ2WoXxZCrmOqM653hpWqUt89Wtmrhq9
JzLxRGZTGW7vnMSDf+GvCJjkgzoW0B4cPnVbKMXeBkncAipdYhRLR52UwzBJrEK6
YS+EWbccQXu4Am+RodXsNYh/svAegcg6DYd9ZUjttTbvbmjfWQucyR9LoJZgWVi6
tXOmBcJxyXtK1g8yTgG4erVxHGU2k9wr1/WeZBVdT4vpKARgBQrcME5dozatNPSe
q4do6kcQ2Kih2JfI/gTMQQyHakSSBkB8fEXe38T1WGc2p9Z1KpZ4lvlbHXCo8iMf
VgT9KYSNsl/EA7Clx2NAqKbSAWJ1Y+4u32lKaldDPwRhk4tikSZXWI+VMDdrLwp9
dyEHLF+FkpCRrU8DlhiOJCAWahItBdwiBFq8tYZOPaEO0MQNJCeDZhtDaoPNdPmF
uxfruezinTtxTJO+3ldyAFBzuSF2J9VWNowy5nurFcXUjqPVFfTeNOBp+mwZatFU
F8waPVGvMmvipWQyzzJuqAH94lTJzCPFqd4BtaFewHRlfu0zpTu8uGrx9xfVZC69
RZ/kWUAnU3tm2Ph3v+cS4JlUN7amLSyXxDP6G5IIfv3fy8GV1H0Jx+j8YEC516ML
VTl2uEhcfypYfwRv90gtlhYwkBNyu6i2/u5Fecu/n3QeXmHjI+pIKRZlGbsPTD92
3pZzDXFxCDxoHkOqd6+T6X9Sttjae07SyVYg8dsjAC5PsFlmeN9mHM2qASYKRJ7l
4GaKMRfwO5JXY3rzBtCrRCKZwTW9WojQ2KB2tR+p7xFT5vI7sgACjmm3UfD5co4M
i7LbrFKKQAYZ25rHA5kwidbrwAYmdm3X4sTCDvweTX52FbLQl/0zJHgRAkojdaxe
6FaPmRmJ1MB3tGpwn31ImGpZU9cNEa9mdtPz8SUu/ycBRQfwKlO1YUXn7IQ8nvCu
7aLYH9oTJMVgjSxB0VFTprQb9BkLTFSS/GsH2GoYtcBD8OB2Cg4fsi+cc+gXje0P
xj/OPoLQ4h//onSVPMWG7ox84Hdp+O3anc7st5zmGis1lpoVyBuNWihLDeAGkykq
61W1lepKT/9CONJEc4mcD4eu7WW3yURXrsLsBdKeo/BRce/9VsIlAxgXuMYfPv0T
c2sY0/6V9kA/mqkiMtX4ENd5vpMff6j6QyT/6iHbULGYTmYrGQO02FbfcV/BzAYH
BhQLc1lpXxMMfXR6U6GGABDUNYgRaThRmTKoZxYYdluvZ7fFK6LGPPN9M/EIUeh2
P2MXBggqSFjwN4dSLD5oa2LpvULJF3Ssl/8+cniKMGvwJF/p9cJKEuOVWFpZ9th2
sxyuP9byKoVfOmTpTOeTzUKjQKF3NadpzsHHqN1YHQ5oJ1h/CzBKCiWygJ1K63YE
p9JKaNNokaEfrs6vTKYuCjb+MHCBUamJDXT+PO/537aBwIGCA6PnczEYMe6/n5oa
2OVW+r55fad35X/0kD83XmuMcK98TY3wleRDPQ0wujHS26ZHtNbNKN5MmFg3dMfr
n+XrovDtdrv/CvtDrqOZ3TnNdLIhPKkLZFzreu5AYobCKB/7+GYGHNkmxkS567+U
fN9CqQ7imIg2WJbOzTTdbBqpcN08jA+cvkiuXE7acgNnzt9QV2rH1xCPf9cEcth0
5GnavE5OUi8fsFndpY5L04YTJAlJ3oOktYh8TqHVj2wWm8Qh0AU6e2NTcw409eN1
XVnQAfgAh/b8Ucmx1F6Su7/m6J4E46IwEQyri7F+G10C1k4I7b5fngHOvfGd4gdv
NqlpFbImKNkGtTnnAYLHsFYUwxNpfowFy/JwFulcti60veiouoqV+r/oDSS1/jKb
SJ5nh8zxoCF9fqfbQFFqztNdsCbMQ0LwDiA9b8s5ypNwm234hhb7QNmQ6R2XFDEg
LSaUT8p3Rf650/UzjHSCeYsR7buVg6eN6END3tViTXbN6g/NkNWDctIXxkocRJ0u
H3/sOIM7OQex4z9QYkoz5gFdWOTo8BwIg/c6cABgwGF/AEHy2iKpVQ+Hn6i27w77
0zrsj7tc+A/vVOU1Crrk8F4Zrj6Q0YEGNSIMymGWohOIXx/nMwbJR5y6WrU5aaAw
WHrm5ENyogwSxkD+4aDQ2rP0Kv49U2CKcTVR1GlmpwChLze0k4JxN0UFyyBeYiap
2qU452GeD/JH9NxB1+kC+4KW/kBiLPAoQx75JgKby3PlZkFQ+53SzCfhuM/47unK
nM6xED7lRL8jqZCebrtROTkqzOgcLGSrQkKAZFBZQvVl0XV7su14qg/JrAWRPpUF
FCAs1de5DWeibeBQJ1KNSaEUCSh70hl//CqaIaSs1F5iQ9oyaCVeNWR/rqx0vnr0
pniG8z1lo0Yl1Um6K1Uf19PEdUuaIA92+Jf1E5IhzAuWR51bPUbUERvoJ9TZbDRt
yG63SU9bl/q0QzYauNAGJrWZNLtDZZaOI387AeimLyidVrgHqvfxMdNVP6znMJOA
Qyar1zMW32XU8uK7BxAfFaxAF7Hl6Q3VK9Oog1H/GspJxCYxAtA+uoe0beUfsx9R
D8kwSlX+Ij/YJVnXOikWiywO/pMwjsuaSEl2eJAOWsgzsnj+oXvSRQhFH5OmmxCQ
KAN9QjeeNVlGOri8t/QC7KoX8f75QBmcRKkFjnl26vSkTGd/YOZqbGHILwHe3RMj
jsUJd6kDfPEN1Lkdu5Tqrf7ygwsr3AMBSwb1OE0uwvaJcfSrhJUMlJCA1XQNGN68
7iFq2/5h+a1JbTowX1o7rL9sKi/jDBMqeKUhj5ba0n5/LHAuj1SB/9ekrWoGy9Br
0HLOrsLmETwj25R3inQPDNeF8tM19hrDlO4/frsLC73B2TXNHiEtEFqaUmVS5PHp
DwzFbjw5hSAySlsWKz6iQ279huevM6792LDtfZgzjQGuaA7AHuHHEJNRWrGvJHWl
1I64snckDx2qPbTP4rYtqkTPUd5uLD+YntKN30+DJtVmUMV5pl9BNsxv4/hzcX2B
B3QXSRnmr5eLf1QL5wWpJkgqQmUxpXeDbfKZYYS5oXBpbbNOz37e1joN2dmDs8K4
tckGF7HMdWyZ3+ROPB2uK53Tc+ne3asLb2qnqouci+dYCRkQAm0SMu2ybMROFgZR
M8qACcpWwKpr2oGT9LytcqMHBAswTy3D6mitmuwZquQ2qpIpiTQoRf0bQPPfQ6Eb
VaPukEs+B0SWZx+xddMVj0RruULx/qQhtAMk3YHyvAjeHag2ysfp+R6kuBEgg6wR
H0EQoHrSy3pdw78VFRn0XO2FtYQvC+hrwjr2xDLCbnWbCBNZUuyVuXekDRPnIOTb
5VVmAFotai/zVUAoj9vjQi6EzoEaDKH7uNWY7UzopcAgdftoi3mgw8yCQakRiYYh
/A3TWDpdDTsnZNzpyUcbmX3WFMO2icI40eOWzFXFk4CkNHox7HMWLp7SVt6hKuMm
+Q1C/UbD7EZS5lhU6it0QUqMw3O1AGtouGYjr6nMgC4JyU0CqXhWGH1Oh/rQ4rCS
HvB7ddXWK6gncjNRAB7GONlYO18C5hNxxevkAN3dc+dczvclUm15BC3EBWD4eAVG
iYNx42HsSNUgdPVI5BoI7qxrSx0Z91iMNQBdoxXBbz9uzt5b43rOI9/bIfzsqcmL
+L/2KzHsQ2ZakYJB1f6vvxvGTJdiu1UsutHyJnpvr4zkS81GJCnOBFyCX2i8d2Hd
fqwyF8hyEbfLedE63IaVqFdVC7kkxSDjyZkSx7iwvrXGhX4p3qB4blRt+eLL/TUP
W4cNPwDQUWJ/KfR8dWtbmo9KWVdcPrFZ5pQ3nCoPydNbldE3pqD4rOddWQIETj4F
KyjyhCv5cQjCYTteTDp/Ei4ZPfF2ZnDMlzexZ1HLM4GgSt9HiSLKRmjPEp4bVlF2
AGk4iKgkNKOe5vWGy2Yo5bWJ3LLrdbsXMrdCsPmLSAy9uQN8KAj0xvFiAyh5gr88
EzkwW5lsDN051l2EUciO1RbLYiftJDfngrVLH/3su83NgsgZ1PDmOx1W4gkJFVn1
UJh+dQrd8kmtfQDtvr36nmXOLG2zhEyIBurmsDeGmwCHCdrYod+1ana5DvRT3RfX
lmb1My8qpdEN1D9XcAlI1SvXUs7iroH14on1dRlfgNtoecBVIigXX8W55WhSPVeJ
oANcAxyovOGQRboPWQ22KMnqxtJdDMRxEHxAi5NhSMJW7Mqad6KmuOmWan6MYuto
MS8ljTr4X98pKzX936HavqM53DKWpDNSLLHr8LZw4R7zctay4yCtFnBK8RX/v3s6
c104Rx4YNyynRDhOLoddAd4DFjiIlGy8Dk1ISBe7gbTz/9JLvitX+VK55jdpqEIY
tBLsG92SdDjs3j1t+/24bOjurOwI7QrakJxFhVoHmOXRYUHZ5oMwhb7+U5QmWyYu
r3Zb4HhfkFv0fGaz9xqlr3i32ZMvgiUAZs5X4YdxIPS6QX2fk18JRRAsuMUS5Yvu
ZZLmnF/yGriaSIgtSnitvCqArooU0mWkKeUxwgtZpkH2jRY8sLmqgCIfrS8rNitV
+krxKE8wrgFazhC2ZPBG4667tHQXMMpNORv4CvuHOMtdWYaRtbmk/mPN7FSHIs0B
uei3lfWK44D7WaCsCLDClPOe4ugOB7JeMe2VMIlSDigfq1p5OePf/R3X/ffl8B7m
OTR1Kovs66ohv9n8dV1ufPKU6dz3S4CD7VO6E+eYBi1lnv67HJiYPz4NUKL78qxi
9HEWLSiN+gMpWtv/jK6JAiqIgohIVlBpXbXy8PbV5fqYxlzy1rLSeVjdXFaq02+p
vv1FE7ZPlaq6DqdmGfC5JtIBJ+sWCCU6ch4CjlhhgHMD8G68Y0vuHjJuAGqklWe5
zvexT/JOSHaPRtF1z9As8QGpzB386XlCgCHyhS4CM9E0Qdx+c/pzqmP0Trgzi53B
Oah4U8romD+KkxzGo+HaBlma7UbHRDHdv8ByDhHeadqRz2+d2PsebTblWlSRivkP
WUjY7m4M3/gog/up7RwoTunslqIfFWcotybWcm0Jowl85WjfEJfZqK9NdoHkhP4j
tOwT/LVLjQHF33q+7exvqW6tjoFskgGttt97Poia0MNIYwceauBWNXoN63sQm/+/
hkIyP9oE+XoXjHDSHBXwVsjuTgHjvbig1mRCLY7I1/05w/YzPtn0UO3MbKAHJkxr
Nq/wkEso/tVySuub0HLsCgBaNxTl7X7xODzaAYzVl6jJ1z/3FqDP4mP4N+G08qGn
9Bbo+bT4LOsRRfkQoq+hKdt0rJb6fbka1bddsSav7vKLAzLSUI3pssgVKUqr1EhU
ZyVxC49qKbm7FxRHMyifcZUKysU1QKXb7KBZ1fUuKaPGsCip3gIX4U+G0Jay6JXP
xNUW7oc/dy7KL3lwvVAvr9x7z4MuOdj+VCS8cAY8EFgtF0sLmYapaoFg/RrkbsZj
+OOroWVtBCjW7P+zkcjKQwGtr/4LfxV7u9+jVq44vSW+3MH8b6s4K8RW7smmlqSB
ugJCNJdARATvK/+Gth15CvQTh9DmnRpmWPzWiCL1yOd5XRm2DSGAeW/Q8vyACDUw
X8/Bw2tvjJBv2rYS1ZgZrc66NIBkDuBpdgB5lI4EjWJ9th5xKp+CP02vjBoLiniG
Vq1MLxU7hRXbvI6Vr0bZZjy1bEAx+qkOKVSrlKTdSsVY5F3Lg38bZP+S/iVpM5Qe
H6GNAY6Ib1Yo82ar1NhlzvO2uocJt/Ce122XVxw2ziosXuzx/ISjHuuTaZgsKhjo
Zl26xIfr73/jwQ0cClxfnDSuqorQ9n1Hk6Q+Cswwnkog3rLpB3C/nKqtxRV8zykz
1973z88s5unysMTvrRspcRZNZvrtod070hdGubBJFjzz7Z4trObnM8LjArWR9rPM
lqWkIY8XlLTmrxsNDE3AWg13ZdeHPOhsr8b0GwZQwrWum1IPmxQEBU/MrZ76oPrz
AspKIWwl1kag1lhTZeEf42ZHudxwNfT3ZQ4b0p69v00G/feqAxF4iwTLi+PypVwY
N2hKUbB3vxrJXdTxYc41+xN7GUmjWwvYt6fTGQl+3ykyWFWz/w6XuWJgRLhi6Ssf
rHGXEWVcJH6fUevFknpPZK1kL3F2E7bA8AGw9gc9DW4eI1AuzRHJ14Cb2Nz65EdT
6J4D+aoyYZ1V3u+Zhk1NYCj2UlPX75nIiMryaLwoH+prQh2QhAsmKOrsSPwqIsiw
nUWD+4G1XNeX1VNcBTdIMrr+D/1WV6M3Zd++HCnp0q/4+RDpjTzN/da0rshNgtWm
ehHX5XcTYfYIpUvPWKwblkeE7Lrhw37CqGoYedFOBg6M2VkA6Urnb585kAn8q8oj
jZj1lQMzmngKOps2FojQCMFKSoGLHQRXBoBSiHaX/ZANBC+oVtdn3ZQ9X26+1u96
ilx4paG1uFuRsS6vV7VZce5jaGzl6s1yJd54RicWW9v6EwUNWd4dHaOM4xjRYLwV
r6muP6+XLIWDG9EKt/liUWJa6iDMYFOg6oVgUnQNJR6duMBfBRefVEU1V28JlJzF
294oIohRe3zRdCFi9e9yCQQDD0VnvI6Nj1B7o1RQ2lNQtnxAPkwHCzPQf7wPP3qq
tD6SAkZJGM3DjWhixcpDKLbS7zkTNBBb0TBnSkcyQ+2uqOKwd0BULjUkOaicWvia
GMBRq/EQOFjOsujPwEgKv2gGqy8IFBRwGMmVf4M4P2cVdj0/ovNSLzKDoI4ZR3V7
iomUOffvxy4dE6JJNdOCdqZi/kpPPQ9K4ffA8/H+9+84DR6WvugoEWUS3DHV+inQ
06lv8gThBHijl2K85bn1/qArETbOfs5vcwTSwiYiIfmJuuEsBIwPG3GhTphJZzb+
735kr3MdJ6UeJEvs81Y5jRSJTpgGRUyajU3zXYhni0+2UBIw0f3iA2EleQUOwX8H
uu+GAoyUbWxTx6EAbIrVcdj7C8yQFmuigpYfOvYpiSPZiaLvp/VIexbHlPzr8hTZ
trqFhie5Z8yMS9W51OfwxT6EyREDQxbZ2yorR908DCG8PhR+X2TClQI1DR9cUObP
H2QntRsKwz9T+1cUrIT43RCrmguSkH9u3haY8qgpZBjDk1zu1LQS+rzkf6RmEIeH
rt0tskm2hvvnyK0xByMfgvcjroFMbsqYMaHuwpIbgrKHylc2EBbYoU8AAA9iV3D9
FQvy1lmPU19wQwAGgUxQJZTjFct+vuJJzQ04aCBTU9W7Smjx7ajOjpWwQSVjdK+K
PUhiHxLdtG0uMwXfPzjOF4hJR9Rp+KgyTxJD4SXUJbE1ZuyGzFwthQtNWhr4djP0
l6i9taz1wBO6abOBEirT3L11kyCLAbnPl5Ep1Muz3ZOdW+SwQe2UIqlWCRo2Lke1
lMRoYgqbWKMQuQrEsRCOnxGRg4tiFL16glHTQPD2Rbej+VpXLAkbJiov74IN6TmF
R3QNeLUazCbD0WERnUxHPVhAIpqpgjtIux8Vy6sKKhak3g/ABDiamjnLv8THSmab
PpMFAije0jiUsEaFn2bq7S46hrhopsupWtfTD7JeDoGMEKk3Uf148Qq9BGunuXd1
Y2fFMDVvBX0WFU4hDXwv0M9ZZjw71NslYJyOZfM5bDXFjKwjOECeiZyJk9DkmI9O
xpsGlpI8TyAxHYVYc+6sNm4FE+s1PL4zYVgTfLMrvp8BT+Cfmkjz09Q2V6V+FEOf
4EThvEacmzyFdz6whl6P7NpFbByk+rSy2rthEdhBSohQVqO8B7KI6BePH4KjDsp5
v2Qs/dJfKhIFhwtuokyTkjq+yzxLtjVwUyluNLBWGd/Rv9X4O5Fr6o6YIwqNfqSg
h2MPYipIsntugBY0pXjC5jjWX4roeHHvkqTmIycCZoT2+PX6abJTURk1PfRJXTYE
YLCFkSjepJRHZGoLBml+p45hYbDiGBVAqDqkczvKJOx+SVW8m7VS65o4+4CYTEBA
QLHz0JbQdyeTzrXV7dMeNwGJTS//ga2wsVO6Ay2pMCgTRDnrboqLum3BjzLajDyv
R2GB7cuwUgD6AkGefsLGvqFEhIb1EjXoaJJ1ovht3CPfXXMltp8Rvvc3hrQqpXES
G3j1PMMtxioYtEnXZGe70C4KYH87lz9Todom2aL3eLwmlzncuxHoKmxxA2cNyWBv
l8jynuTvnt5PqCSSlsDfvLsAEFkt2nU/0snkpYAk6LA+ujH4j30NBXiiX7TwlrW9
LhRJ2WDO3ATP4SIgmNGCmxQT9/MIxnP0Q8ciHCECs347Ec2SbNh+KEZWVoINryql
o4FUli4xnBiw/FPfSbSiW7G8+lbjn//s6ZQJKXHMjOzxY0Z+Fm7k6bE3rzy7x5qk
vMZa1nsQdqQNRSzBEyE6P9S3+KMFl8AeoDFJeUW47fxE2sHqfOQ9DTOW2gMtRdHt
40TVZi06WPxghTahWEwrm8O/Ef11Kq2+tl7lhaRtG3en2PsOGw4HQhzxzCk5KZjn
KFUFf8wI/cV3iGExVi1rxp3OJnY5crakVPHEcAjaO+21K22JvreslRm7M78276as
pFoVnepP/M4XM0YUNcIexp853SRM+c2MKQK/sCPoX7Tlwe15MLKaESascgKP0KnK
FRIySc9/2zOd2fIGjHo9o2TlbPj4N1z87LHxCd3Mpl7R0XLHGPjVEM5yvxXhP74R
f4z/zM/vdUiYN+Hs8Zg89+z6kOBwv+wVnx7BinbxZst0yKHs3j5zEM4ngeky6xCd
PMNvMP53rhwPKzC1PyLys3+7qIjTLVdG9aC45y78J1je1bogVLHFGNLDbSAj8D+k
GHhQv2LVRgvNlwycVr5uQNdhx7YBRdYo0J1XudZo6yGPip5cMpYLuCGR1yDJgpIG
ULnaJ8K3AF8b4kv24fxwOfSUt0SflfFNYWwTEy5m1HqkXlv2trpUaIP7vJtmJwua
TeWEwsPqUKrqM0+U59V9YyBWWfTWMTF4hPwggujgNyoK+twLbUUyI8H3jwqWxSc6
+q95T3zPxlKAwpbIxAhVwekGP1KmQX9qAc3IGhxEqKJ3Y9v2KjNxpM/cg1qB7mBm
AjfVg91Au4sozDGyIHH8tOpnwLVrGvsDobvMZHMK5bU/WG3uPOrSqb+Se4NhikGI
Yl+TmncxFimIw/L98otil4Qo+k6gmKybC0Iu9UdW6jFlT4LSVg382gszxskbZYvr
V6MG7OqMQmISI9RMRvVZWCvf/CbbA9IU+u6JrHHUFTIyOBGnjpB3vyRBmz6gDvKm
aSJohmdGfJdKE7f+FKIz8DE2vaIKl5ZTk7Kig44gefFabY46YkdLQelyyKjN7W2v
k/9lLC00ANaE6Mx8dayxveVBAVV6SJquxVwuu32+qmKp8PDN4G4odxZMByK3M5CA
T6lRRt/73GC46TOxdhG2idI1TUG87nc5AuBUgJoh5MwZZ9bq+fOdl3exLWxITHXY
+ZFYFuVPfFPCn2v/i2owwmZzsdqXknHaY5NNJVicoahPr/lc3uWUytQ/ISys8DjR
TWf6aOinBujY94nWD2gQHYqJaFQB4gM6DYRPQLTeWc+AH0WZUTBPabWNES6b2lrl
JueTx29aGlPyUG5LGuFSybTmCX9HLR+XAtaXs7+RAHom/Pr7YVKpKEb58aeueOan
6GzwwribaXBRoXsIs7K4I60UOmgqQ3AVxETQ63h0xN7JUwfxANTmQwrlLy4FaSmr
DKSVyhJaBDDiSmF1WLffL1BHtQ6P9DgAMgG87VNn+I2R4aBw64dTa3p7vN4f3Yb5
tt0gR/LYRPlBI4EhoTV1cKtpAuXRlVKfJKdjsl5zRchSQiHijhSR2VmPk7y2Cjni
gtauXd/C0P/gQkcGoTio7Y4ZbcZdSBcY1K/Vtbf2R5wTy4DZ3f2dLnnmbo+Ing5M
AVQkdVMWC4nWlSJ0VibZL0ltQGGm1ZniaB7WUeW0LayMqLoY05a70kCRZUL7+Vs1
SeMcJOHC6BRy9oUYDPOq/JQ2y4DwxxvuRKfIodf6B0wz0PZfZOPXoGQ2YDD+rKUs
cDZOx0J1fWwILRaCRs3w3I1XIltTh4jmyuVF2q1+MWjqtD5oHs+LJGPQvkKeAzqI
bBAGcy0fFWkg5r2MN9nm4jIf30E9qE5Y4QXhcXo6/l6yFF+SQzaR5xybbI1oCLwA
BDzYHYn7n9pAlOjSTrpF8YLVBO6ixrcUOu9UgsGus4a0+E1BBoIKJnmr9Q+Nz8Qs
QgEJR1s3TEumq8nhw5axEtscPx5j90qqJvKoZ2pKp5uwhwuRLRLpWYV7xL+aG4C/
h7FZbLlwpdPI0tgsgYc387bZmrw344RdTuyqOt634BhSdtxPvFmJiDgoJyzvLWn2
3bajhppMczprYJgJN+meQYCPf7xwETbZ6pewGisHNNUH33+xY6cB2PoXpgXs8AAg
y389Gh2Wqle5PEhGxpyVr2ZQ3BHXbgE12IMEuteoT653I5MNwSgNWSDtpESlPfTY
5ZINF3lOkj8NJafXw8iGKXxKsc1cgqGLvAWLLgzdFIZBTrB7+9cSDjf22zoBBV+H
KYHkchkqZszFs0ZhGfFJAPWVodjZPtE9rJMNGZevnpS3INwfOGuiX45gTx3NCmXC
aKiKvaFTDzo04nDIFwHExSnsGhn0WmgliBmNzXTMtp1umifG5UydzkinCz62ScJl
GEVF9ScYs4VJ/iBsNz31kfu+39fQPK6A5f7wA6DxY6ErSyvsJjyc7OXjsZRN2x/O
D/gUc0O43/BfjGFvu6uD13RKS5N9fem8qzqUrVJlkvDecFk8kX6D3UkQ9k9Ylt6H
T3GWMMl5Gj1Zrmte2+dG3qkvrcm/19l5Ngn6ONKJGh6qyR/jc0LUxhA8gxIklIOQ
WLsq6Kz+JQ4PTnu6Qa9oEpBX8Vhs4bWuIhZsVr4YXyKeknWbO7UZ80fG2YAv1OQh
+t3opO/nAbMf0aO3oby6G9fjecIbOSthSaWVx82ywb9iU00RlAceYL9PL1u04GeN
lRha6XIRyY0EppfWX+x5hGmfzQPI4Qep/pAvqvKEMDhmZnuYrDXXqoGDMa3SBj6Z
24Ckm9QsIii25P+s0W9V3Sn7pC9aCR+tSwxRvJasEEGFbhl307PunVRM6wSaGc6X
117Lo2GFZ7sTmnT1c/As5Kv+1RXPtI1/TSqaxqaKlk7wscdc/XSQ3AkZLOUZqZvf
N1fFFLY2iy0Np+WvPh3/LpdKjXwSgdYiSamsAlyLdEm1lT2XUM0ijIqxJ+G0G2if
fM1a/ojBewXXDBXBkR4IjArUKRQVoM0/VYKb77bZfK7kPVv2OnkmdTGkPkcW3C12
mf/65uJl1jOzusdoEt95XfxIswSAN+ZATq57l0fbOXjdFXri+2ESxG4kUacDtQ+n
asc+UFI69plzRMLWGnLtDke5tOSwZY6YYNDcWHPQQXqvpITXc9zc3tJIKipacarn
E4B661UJwUCdlDM4EV7FGMPPKB4O1ex4yczRMxk0ew3qxZQGDDo0vLR/64Jd57L9
aXyBd5y6WJ7zclZuLLhrZ37AlMHxVAczy6zLouTz0ilb666SnRkCrZ14Dr6BkFKS
eHQJtNCf3eAP0cJiIiO3bTvUA5QgBnM/i4tvSd1Aq4WNTad6n3cyaBLXBarE2naO
Iz2eWvit4lXIIhFeURPrUqO3vcarrsrmc3lQaQlPIqj9nJD4MXhFAyxq59O2N3kH
nz6PvQcGuWTdaTk5hwGZHAW9pE/hYCZkxV+CkBaLbzd4PILpZac6EC0zbBKcmq2a
BkVuvSDJfuCE0W2vQACQTECyomqIwU/zoitf0ABc0MULJnEuonpOwA8GKfVRwUmV
+5ej3fwlIubqSlwjZNHzAQE7gIq7AS5ztdvvBlXr+iXtjHpPT/8nO5c4qTNOYnvK
jNDZBgDI9oaRy7//836RlbQk/o7mmvv8OfySaSaU1AZdK8Y42ac5TwW6/KY4itqA
LQehqswWNnd3+7GeLa69JHCiCwlLWtj5V2mXCYyPkkNpZZmxwdhHiFoMvfYA/dYS
hd1sN4GWMf1JTP5pFiDvPvoZ7Ylzhsz4LwtoXnkhbYYpn6z2h5y2aPLerI1NwoL4
tdR+fulErfgzMj7uLZ7PzSJXMeKCrGSJTeOPNY1A/T2Lnx1Dh9v3Ip5BGtRF56OO
2MfZdNgku6eK5kAHhCsPblZ5fo3Ed0M4Q8Vh2Or5shULhhrv8LUB+MF0ETrdTmA1
mS293DSLJtnA+NXJ3GOh2IUKw5o8+2TjLOP/uz9KwSVgEeiJqWQwobG0C5Lnh8zJ
Mqoo0uTUETNwShp+DR2CPStkz+pVMI3amQCzdM24boPgNNOIzIR3XjcZc7CZyLwN
njm7HTyugy9YsRrjgopi92/0F2BaBzQpf6tqotYRAUBBH6l+dWT9Yg5FRUjWj62X
7IUIGdp6yFLSbJs4eWIbWIVFuAgUhpPVzfgWGYmGu9Isr1jytiOdgpk4r4X2LasV
9cqqN94f9cw+Fon5FVK/fAdmh1guMU6DCesP1HXKdxYvE3QsFEXDI+Bhg9KucO1+
ttGGWLqKFtYgJKhuExZ29EukFEEi3dnNpWibqnNyZv8fbXo0itV3V7edfl/Wg53a
p2PZ5UF74GcKUQnu/Chthu0ppidvI5GGO93kHUR7m0MStCvfdjWvPADHqh7lyreP
Nqo9mZ5SsrqsGEYqhVEPlcD0Xr4wytisZ3Pa/KNN5nRLUltnIky+bUQpHYet9oQM
YvyyQae1PkQiQ0FuBLluxzNBj9bcWoCDz2A5KFwBG5tqUJFro1qfUxIOH9lBDkPw
9ZIQnG3+DrHaVp0Rm9G3F148rKWD27U2JZV+dDXcGRhTbZS7GSBecNLVtfMqBgU/
wYj8/tzdhRUD/PFxo1Gi6Zw4gaoqzybOSB4Yd+I9jA/a4aYZUQnGiiieK/eIHODh
lt7rYN2bVTT3ZXRgHUa/koYDzcmhDVw2CB/uKECTe+J/fERkZyR9SltkHVODFDaG
4EyZ1MWsb+DWvcaP0cyUAwxX40XKDrKwc/LTo52Sp9DlxTf2rKZG65trb/9hEgP7
xsz6M7dOwOaLocMBH9qtbYifPIcp5s838ECaMmtV+y1LsZpydIY+AqUbf3c/qBcl
yJwB+zIZZsItYrQPp/EEU3Jb+SA//pwe82r8YnqMyBqrrXSRFzJ2lFWX3RnqBTlo
fB4qCBUzXL5b6pfScnP8AbgXHdVdWqx43pegARiqSxEPcAZvLuViL3iLC55p+KQB
d1UI57xL1rb0M1Uh8BkJzdW6edKSWZZeFDIQGv+MSXLFKQevxiVC3N4K3X9srYW2
i9xuFbGuTF+CbWkx8PN3AG/MAPzNC2qxicu8OGVnCFFOUmpYZ3cnOQEe3Z41cZL2
um0rlO8VvAK8tBCuyxM5/XHCuDRbe0ySbyXvfseuvRaTUdtNB/U92BS6xCtmO8Pk
CMz0/ZI7eu8Ux7KiTiQojdtb3OmLkljoIYwg9rGRezuZ8FQuf8s3uBGLJgBIWg7z
+1AVPP+taA/Pi3g6aMTTUL/kxKBdvdGMDAaVmmMlbIldVdLXQav/TJtrwWwyxecb
LPqUGOjBnlTkGbkaqOY6K1uGwlmPyTTLfsjWqY0y/4gehLTrXoJV9JKQexl0Gq3t
Pz1qmsN4GkCS++OujdIThr/Jgppsv6R7ecX8YAzdd+HKIiRJbAPaEbpNEvr/X7HY
opkwhEhpbvXJsxjUxhxWdUOveD+QVhQ4odLOCMk13of/bepLT3nL5UmdDbDZq5yh
7I7OIMlHW9tjwdXEYmzYitpSvoOWNv4R4OL3EwlBcFwZtDLIJzOWeHZMgSBWYkRO
ZvEic/kZZNw/mh18K17XR+hVhMYB3DSJSojOt/nTKKoQNazc/VBnP1/NWlyWgHmJ
iHfijmqSlKtsWCRr401TIpR4kkYsgxUjlD8zhPdYf7+MyU8WeV9t9WdvK6mGUY4n
w4JBs2dZsAyOwBqeA3bxzopXg0h4dOv0bvV55P2VCaH+/H3Fom+ZMdGdRwP2keyB
cqP9IBKGnhzoleH87YBOnbPIq9gFmnx87oqHGurtsZDEwxtbBxMeEPOyF8RCxxtV
a7RnPxACY9xtB2MP7Jm24GrxJhnvIWXP83B9j0W9UzTSEsLHT1/6eZkVvmxBfuTa
DAHsIyudm9+KDJecW5BYNS7WaolqvljsU1JhPv8aT67Dc1VMyZxnhBBtS+J9vZDt
pMyBNOou77eNL0NCgImJwHelRIh6T2yf1kRZSwRYOgdPmt4Ajpj5IXoLJFEuMb2B
FYqSMMevc9gmBkVy9ZDOVBQ3WT3+YM7k9AlEta4us+uu35n43ac/kvDMfsWNbeAC
kjl53p2UCJvxduaFwJFJUixofPOikzEJ5SemcHmKAxNbUGDqb3R6TIzyGM6Zb3Fh
JxXAF+ijYFWQ6zGzikeXXpkRAI8fvgEyitA/hW2Zk/YED4HB1DPSQY6lQgyviKZQ
ZcaXsZUZZqcb3BwLiZCJLzrLinGE4VVdrWXKa4BxvR3co2Bk+pd6qIvXxCxFV873
SrxLLdkZ/Swta9mF7KTKkNKMiq3GYdtUhfUvVnPyUCgj76xwOrgMofYvUrhitJ/I
+A90gg2+dk68Lv8PTxgrOVpt7ke8nHCwFd9lIiMnHNTcYm63XcP+HBYQPTembIha
ru9Hr4CmHzjf4KughcQP/NXd1e7huA0t69CUgnsZOJSByY0wl7RE8v4OF0q09rQh
+016T6D68/C3bxZKiNWLsIKkquGgN5fZoLrlfaOfevQRCcoA4JzTd79BtpA8fCNm
I/xWyuq0YQ/3aysmn3Y8LSW2e+MiiZ2G4A1s7LwRU1wHfdb5Rccyn0dxqASgaGqd
ZHhumkznDuzHy51pXWiz1G11cPP36plEmMc1atucP1btvC0cQlOjtNTx0rE6xpF9
cawv0vF8Xq9hBrYt25MoxaeokPxRzpNTb3tLRhApoUM+844dYpyZNwWJ/BpcKVeW
X4FZGV+fez+F3ccqunJ7l8kLXuKTYYu422s8+9LZ91sAWADJMcGJrZqleiRlvVVH
eetgMZqEJx5X6PlhFa7Mn7s9rEtxMRkETdpPqYRiSJdtjxHKnd+sNq6XUs5712nR
INXS+ziCv4MxcQnx9ICVXps+/md84DE6zluNvgs+KqaG2HoH3jSU+3MGmPgExoLD
JEQSa6zCaYtVvrssYCItKAZxKyaLBvNHv2Ysle0bVyPmgg/yidL57CLpvnLXoqxQ
kmzi6MWHwrpBEaOi1Whjdj77+PAbYnHMikpumCta9zOP/EJP2JJmAjeqqXaePE4Y
JqDXsdzn7nhIiHwcFgM7WP+r7MejPW128SohsBlsqZA2Wn9dzZOLjPI9eWWSERwr
aCTdRJQAE7wOv0Ep8QNkd59RaC/csAjFLkDs6zenA4qhfjeV/RmdD4xdCB2mEkSb
oZgW9/WDJOZ4LoQheKRLJsXZGtZVsXeaMzUNCti4xZfosrneZeD0+NzwLeHsEZNk
YEOm49z8QUwFSPGM3DejTh3Oc0zJzSOaB7/cLlRt47tPL6ECPHpGDISofmDACfxx
2dDfLnoH8vCy+0QGX5GHPtpmD2O3JzqCSJfQbmN0MndLzA9TdwxrQzKJWTt8iXun
nsOPLl2pzy9pzl0khTVKLoHUGuaChn5xh49gDs4JkhfJzQz67dY7owP0ba9Mzr7Y
Y2PbOI7YRlvVU3+hB3/Jve20vmEYh3Gnb1vUErlfcfPp4NfCeSVtakghGiwC4f/V
TlxVgjm4U/VwuMI/Yz8b2xY/tSE8VeXKbUAl+1oF3oSUDZx9/p7gGHaPlqm81epH
hWPMiJ2xDyzWc6VplXv7n/P3LmqVfSA/7jqddjjwy8YMw6PUr4qTvmToXwREE27V
6VYVGGYDoTu3WDX/36HRqgoZCHdnbzZWpYXIH4yz3xjClLl75uXNcoKwxXNaCB85
pbVHAxUqbUBQS3nO0lUC3zQvhTGj9IIBzJ35EOqvmok9Sg+IN5nDHjVgZGJV7kmu
fb1d4AGupUXMw+l3nrkMPfzg07ZG2Km8sLsDAljEEgRrpimYR9eW1OnpGtsjTHWq
30LOIMTcrGPns3q+N4LVXhIUfXmWKZHLD/V0+QZ1xeZWSoJV5WWgfZ0GFGGQMHEj
xj5jCzJqW+3eAk7cBB7O0rBDF4ixCSrGneFYeAg71h2uuUgODF1372Bb8hfy8lG1
xvw8mq/gHSoE4mWyPED6zi2ByYRZOTzMLjhEHW5uqfdcxIzq9Cai2vFA+VB2K0gd
6bGSB15Qb+fvZisCfw+Bly+AGZc4PmsQVuk37/U2vBuY9PEj3m7MRqPxsOPISBsh
hgtf+xp9mxhnm/tZ67c8OQTGBJGOE+i0fMAPOgGT2WG4Cqd4VBr9d4zxb6df5NFm
dt1kk0mSQqTpXh8h5X70DzssddGHss6E6X07G1J4Mx7t4fEWZGOo+psodE2qOovZ
m7HPw0EPl9thdJ2S4Q4CuWm4W6qmVIw/GWH2Xpamj547TKli/j+xt02n5c7vsejG
lHyF2SFd+6dVFhetCmrLiKDauWR6UmbQqv20I2vykntzZ+ww467TvaBK/HgvZa60
65e02Vu5ZIeg9hEDUMip8MO4O+6zN+n2Meo1rnNDocAk/H1j9ieEsefUbWI6IWlL
6ceEv35+VSWXftWR9fXlP8uIsnO2DTzSisQIY7BIs3Wmu2oJtfgZaholaBv8TuHM
leirxx+MhWVp+pA2e8u5OpEA+SlVs31bRpAR7HFRJtXy9fEQ8NBIru4u/CcheUv/
YUBiKXxqM18nITiQsRuwzzuWy0ACyuHXjjKkT8rW9Op7BW9Pt7stX8hvr7O0bcU7
lwbsARo9mW+q+88faioy56ZALsc8KNbw9Io3ICKYNhSleEPq+t4KA/1tz8bnn6w2
tP3qCsFdjUS4RUVBp18QQj1qbldJIiw8+imE9jd4ZB4kadUZtOdJt4ukAOXjlnFj
KelqZg+8U90wskXIWxJNF1KnZIgp/1vZyxNGA1DrUvtltjvsADGlfHZKShOQMaNu
h81y56AB71/a9kYNlODG5BqTvXm1zKjX8VFjWpmVITumVvG4WFvWVUMQfxahEslK
tFx3SDzgSg9at0fc2QT9w1j7s9mqlskIY6enVv4x+QXZQtA4oaFbgCYP++M3Jikn
ZxwiQo5l41nQIBCUZ4RUsOvcWs7wfd9Eyy+KtxnuCQyEzry3bzgFZ1vkghPpU0Tc
+JqDZ8HkTdPtYQIB7nY2Dl/NPnEG2ceAzR/soq118sHFHyOTyFJw+Q5aHix0+au5
7TThlKplgaWLdQ/p0ZjHX4cvtTH4rnRT/gL+But4gDhbd7hKu+BVbr3hlH1rGGmv
kuyuRZssbegNRZW3sC4kvCCFw28mFNyYkBjJXXGMDIOJgva3N4p5GueuaHxVvla0
u5uUiQcGZ4JmSzmvY5dJn0v+Y76ZxOyVEZsSaxe0TkqfD4fL79xFE70LmCHkl5Hx
BM9036qwv9u8MJcY9Zc0HhW5lwKLcADMScwYjcJZOkuMYq4sxiInCEAaLwJfXB/Z
KpWuEkNZ791zO1nCKaWlQXElf1MPEe7tAAFLbWR7UUXeWJAk3tyiqqIw+ro4Utpr
Ens4bwihCr9a/Br9BX0hM3YvwBIoyFPuLtxW5MxdhTuZ2DoNK4TKttgs22CtwtBn
iqNNGh/UI2c05N8+/U2tKLgGBdV49GtXE0cbqmj4BccqE364QhK7Wle876N4FmAP
0iQhtG0mK6HjVS9o8uBWkT2dmsakKTrERme0xq9dkGeCggvDYMiIAl5MEa0djVN3
wVnhI9wT48dw9PZIxs9Lii4TI87oSWO5oQuC/L7N69jDANOpJVaQUjrts3wKCO0W
o9H+SXDS5NRNJgsQsLe7ELZxpcRu8lZaesi0jneAsWlyEOM6WbZDbEje/MNYfRIw
Et24fu8QbIGf1L3w9wikLHcHZ0LwiY7lWKLLp5+fu3oUsXISB07M8Na315BqVkIc
gDS7I0rfPskZPehIDZweEAZrVXT+/bF0AyjSD0W6W3t4Y1xm5trhW3U8YM5SmRaW
ue5MHvb/f0fNc9ArYo2UoZ5QqaG603khEIe5W/TlLF2JtcXaIV8pTi4zY8VXieJr
GTqUKKmcLNEwYCv9jO0DVOILVElcOun03Q2RLLXkNCmQz46fCWZ8gE8gLX8WMnAQ
4r+eOTRaupuIgztsv9sVKx93ym5VUrYRq5F6ynBmvrBGttRuyisEISSBGWEzKU4D
5fw7ITBmP/GObp8IqASxxUdkPEw8TABWMzzCF8jN9R0y4y3FeorJA718LsGkv2cA
oTAP10GyA5JIEXCqhJteV4UPdpP20BL3y2n9qHzyQ6APosysDVQvSmHvYe9xj5HZ
P6IEApPy/qJ27ofP8PFOLaZK/zIWUtpa4lyfsDLzntEeF8nUP5V1GyIbkzMdZhOy
VTU9Ls0QFYB4ksjAzNyl8IXlIOFDVdym47z2F8GpVi/4Sk2hZ4nPyAcHb+FIIJHW
dIeUsyduQUMgpD58uy1SL3tyrDmqFQZNpATm39RJO0HYxl/It9w1fS+anKAAhODv
NMMAvlhDYOdHiVun7EGYeI5XS4jLGrYU4vbg7QCnEobVqr073rEgMVbbVwlo+M3v
DMVa6FJLQ6wJxZ9hjDrBUb7CnVo6rYCr+4mO+jvSfXoD4rF/6hZkAHi3WTxcOQtB
JGZoWms417gyTub9xu9aEzbYhbh2FH9J0iZF32XmNENuHtBPqCL3xf0vU52G+9Sh
mfszbIo5m0ii6QrRB/sP47o5hk9BmjY9Jjj/nNJCDM5xkTc9lcLhgj6I4ymKG5yN
gUBvjsvRa065gvxYaq1zGdmZjn+3v2tXCupm0ov5HLI2ewQJSn1BcQmczLsEdQi9
0JJ6HVMJOCgcRRuq0ldxxLdgGhz1TEQy3ZYpX5Ho8g1kFNw+GOhDVrip/HlTTOqK
piHkNA2idQeenFupsDXOj1HEOvTQGJ9giTcXGE9r3irW5pjZfHnC1cdmU3lVlGU+
BdTsffv/ZbyewELNT9WAlhpHhh1dfNAGV3AV85slqJg0h7EcddjXcmmQd/ZYXNWh
9tjFAAl2He21sQR/hP6Bm8hMBgOCwFVejoSRjSuMugitg8gXWRi6NQyE8Hpem7sf
HDhLVf3dBYMc3M1ot2YpS3jwX5N9fv5az6URV8TncNl3DqgR9+H+nausSbOPAJVi
wF+GmaOETYXScY03Pi1R4+OSCOeKcpVXx5KR13cUOcNZLhoJKwW4q3dLdHmTTbEK
/j5E+1Opue+jby+GkluwqHVWQWg83T+PovB9FYEFiQ8pMJkaid0fiiGLhdpRF8P5
PI9VL05KST/oxue/gGn4leGhBwOtDSMZNxlwXqi0T8wzS5sk6rMMzsDwHWTda9iR
dW/fzZ1QXuIpmDOi+SE3END7UX5MI0jVnDfJOTCeayev9OTGiIkBupbw4budvxn7
FpEJmR297P1sD8r1oEW5YnfhoYTVDm9K3vtwBFV5ET00fKNC8/q2XL4oqr2bfryc
h6leWy5VMBRC9fkUj5MFoa4/qmYp9vScjyd+jvAD6QAGvVZFRiQIPpMRPAZBy0rR
JVFEOtn4a3ME1b2j9MDSJO5iQcj9GtRikXhHA2nCvSE8UEzOM46GwKMktrtLmPao
cnfae4fTy3atzcg7ab19tgPawpcm3qyyexkFjcsHTOCa+4u9DLl3+Wg6tKByj56l
fBghAq9ICl7woPLfdtQuSOSgL10Y2E3Da7NIxEBBCw771jugXnOLP7UeS8Jj/WHp
MCpfgNjCkgXgE8NEzEKiBjvtwVYNi2aVNCG//jmPcwyl6hKZ5pXjpyZc2Vs98efl
/9gsHhFgbmNpeDOlPfv9lDxBe2UPDI+HlTJEcd1iXIPTG47RlgRU9W+l0AFnUrji
k67orUJXSsZAlcaQcULZLHO0I94xXxu+ljW6bZPOboUirI4GMkzNxOjhczf6EfGR
0kGHYVKDZAXBSDpLeYJTLPyZGc+7YVczg+oMRVDm3RjILnL+Qah2o9RdfKsn4s7s
42iFuvg1xZcr4X5A+1P+Cics3KgJRoPjy7c7UvKo7+3IsMqGdWC2h2Q2sqrjBOhx
LigMj29StQcjJPL6noyj6MHOjadZ7LwAtarHtcbBKA1tzdf5OYVA3WAjfsmev/vK
i9d9XCJ7Tp5h+JTzFCef+aRr6uC332f9GFZpsWUo4kiTgGt3ttiLnewKljQOFWd1
pLcNigqzjTVs+21g58KNS/0II8kekbzKQGxVtBHZmJ33TSLURO2EpBtl9+TxbKP3
QfecbQuZnIy6EbbEqxTCCzsD5gwOw4BO790Tv5Iczv53B2/fSOEWF3cgmKxTnif/
MppEfdir/0SeApqwSKR80JT+2LRgxhbAi6TechUj6bfEC1J5NMjrdjtcp26xhYBz
ZAdv5VFjfVYcJzAJjRhlwLsof6qzUa5FXmmhs/I+R48m+jTSCGkX4QbazrumB6D9
66NN2wiAwdncgCvmWdz+1hSmRsAsQsa/6bPZ7uOkLn6gIA7fFSgcIfOxqOK2N0f3
jvspkuh4kOxsFhOdQGPvW/LMGl7I/Nr+6lBdM0Oh2OzGkJq9YvibDZP6/VTRK0VE
C8+e1nHUgVuQWJLPEDsjeOXv0RpzldspJEdoh/qeEfTIfgYCMi4K4d8YDdlOuhgI
5Q1pZ9KmHyQf+j+SZs3z1tnEBTL8JDpB4D89+z/3V22Iq2c1MHum8dBPmTsCbODo
allJe/Feh1op6SxuCElmi0UGEC5fsm16EEJAP0IcLWijW+C05oNor5M+DhVgNjkY
Z6rd7uw62h6zWlQOoT1GOK68ryarbeMmVCQnYXsHnmTBe99Z0cN5E2bzYctfbwWY
JII/SAH8Ubry2tHoWZVQzr0R/u3bS3SVqrFaWp6M794/OePrGgI4Bx/F2bzeh4eC
G7JahBKLGqC+ozSDw7pRh9R0yPL6XVwD4EAiseM4Zkx/7n+Hc31ToPT7NUm+Y944
qceCqqh+mtugOq63YCTz3g5FZ5FNX/mrW0L0g9VsIL7+WlPyEXUYIOrU7VTPRrxf
8mm80T1Zaq3y6DSZbDEgeL99pUbafMHiL1dtpk5ul+otD8f2UQY3P+/wCFdago56
tOlWFl5kFTrryhATqzeKqGr38ezFhsrWqUH4t7rZgzpSLe8DIZf8syeixdI9lEoC
V5ICB2/cb0tSoV5+RpiXEwie7QDlJn/TvCKk8bZC4158xUWUfud559O2oTGRWiAF
WDm9FnLU0SBnMdX1QrPLaw3nvWJfdCBaCktWDRww1aliPvyi0+U1RS1ToJ7HIVEk
v8OTR9HnL7Zc8Z7PPO3Z4AsOSV6UlJbn1r0GtpXXQS1jU45C5KPoUeabp5VSOpoV
uDV+Qd0L6TpDajmhfeDbJZGbcbbHCAPD+qA6qxkUJUbbJyM1F7Fvz6+SMPk+WpzB
K5rJFMmv/MeP8wTwAMxI+1+IwLTMnj6sR2pOKnT9wg6hCXXBoeQbVgrN1HRRq9za
93ZFxefSVfAujsz2pY8mDEljK0O7dh89KPLCVvyMgThUpwqKNm6GQfCb81vT66kF
J08UI26G6GdxcDbzwLk+ShHmE7BGbqPycMzcZOJYghwT7wJ7bzCwnBxbMrfZ79YM
jwcOoYIH8dFguQPAcKPAMiAwXHuWpWsiUIn0ogl6o87JN1WI9Of3TaSQn6gyyBo/
qpDeALTntHX4oBB8B1I9lQefzJdZ4cpZ9MUwclYgdzXahmVjCECFipOdtLI13eva
7f4fgGaY8zj6c4dtWsP9tyA9w0+apypjKfFZYOLy2nvPtFSdgX2jSpEwlpO1/PcC
Eol+bDIfPGcvKtCJVXseQjfReGVMhKYq8/CIdxqA6UO3MEJPQ5OiXsBqclZA8hKm
83KYSJsfsVpv9K97VoST+pal6xIyfycQt+uBkwHXW9896mKqTmCEWMqw316s99yD
A5HCErZHZLy2VdsFS1PEscKIKYV8UvehPaM7AP+4lp0y+q17mEv7MvuzAxuExhi5
g/6VH/X/zkxHyfgchwRSO5Qlkxd0LCU/hiHp9xndmCsLw8n0oRXejt8yzAGYjQ6l
z+ahg6WU6QASr7BB5lxrgtdJBQK2syRKcqXPf/emkVm/3CvDRwx091hlMSQzryZ3
/TiDKdL6RjL2pciO4+qsq8vzGRBGG/JtDkY/VOsL+Yfp6ltOSfZxasAm7p0BdwIs
QuBGCHtlXa/YWGUwtSfaBfFJYTv9dQevpHPJCDsOJdHMwUIvUkglFC7s9348ictv
KfNBN+bAP5/tj0hxqXQxU/4G0dOonS5X01R8on61TMagU96fkD9+172oc8UeVpyl
bT8Q1CtIiuZnHmn7t4CohyiO4WEsXCe4UE8lMn0sjnt7+XwyPRP5w0Cj3v/pRXaD
FH8haEDQHCRYpu05bPfji40+CCKliLdA4+MPNhtGRTMg0P3xDvnGG6q34e3t1N4i
V6OQVWFBc4GGJ6zufTJl5AZ5B+0NlFGxBoEbbauMHULBmFeFehMOXjVAr2gidz3Z
pW4gngyeipdPF66x6Hp20kx76PD9PC4/qZ0qMpoSNjqUKv5Hm97YuiywyRyLL0R5
XGK7VH1H/WD7mVL21H/nrzSuNJGh6XT4nS10eDUKP9hQ6Akhdn7XemnmGfTj1zHJ
v166DWEv00EWYzT5csZ3KTTc1wLqQHkINXoVeG6XxwALp56csK1rdg2H6Z8bjDFW
DBOCZItVSh1Uuaf6vmlX6lKIws5WCn4JfE6pXt4cKKbDFMUYjV5mqUBSr8pXsiHj
K2EBxAFYnwzKbq5Svj+Z3QU6OedV+KG6KsFBV/aRKoHimDLcLNlo9TgQ62LzJliQ
JWcjkstXA7wd8gqgCHLnd9+sJof4N5YhCXXDB3tBIa/MPAmx/H8LNvbaQzhWqr09
AuZna7VtWRS7HnaMDDb/oUgIe+PsFcZssKI6PvmnE+4DVMK1MFh8t8Ets1X2Ry8t
6m96Cn/e09Xib+vE8uGokIoxSaGtyY+hdZxZyo0XfcC6W1zTdUdfpbrGOV4uq0m/
cThu+cNHBt6QaSU4jgklvwFWuPDAZFiqvlctAe2vOe6p57kkL50nDaJJtC+scXa+
hcFWhSD81nK3i8uw3q9Unrrr4cP1Bij1mMjXgOUo8x+dla8CtIrmnI9vQdW1DtiC
CccAHtPJVyEZZqMo1IOmxRYkp5+VJMNeCWHDydoAQ95ROGV2chmPXKJP3SlRXRIa
K+8hHcDWJP1A/6JzlcZJ0TiVlibcq7WP5nr2ll7eU39spgYme6ToI55Pd22AgYK8
DT0xVjmhA2Kr8uFoOhucdTkmj4Quksq0vx87mZK1LiVHloEPa3T7/Kb53hut6aDh
/EdJiU2gjxjzP75P11BzPEslSZLeZX0c0iNFqiPOZOhTV8t+SOKi437/xhXaZEAp
jDY+o7lenfERbQluKPo0M9pDCLOUZtGolJ6mobS6xDKv1/+TvvmMJxWVkX2aW0Ei
wSX6CHECCkS44qiVOuSzZ8DPj546LnMtuUB58cKqOP8bwF+ou926YvHyGLNKWZ0B
XIjZebupoff/WSkU5GsjreEkUyJVejZ0SCIIpPxJccYkwiAaehlg4garJNJu1t6h
L4nK3yHkRF8E4d8I0z/Lo8QlUkAUausKFosagFi6WrtRQILV62yxDNgJUxqHMbUs
zCt7FDv1LwU4rUqxaOTX9y3emeFOYhX011MQChF5UZMZ8WoVbLBXTOHITzkA57We
miro6npM5WGd1zt3seseOxWJYorRiotWVgE8x1kCeJhJO7vbikuPbwaviYBiBnUs
Fcop/hJUBQUDA2Zhn9LhGwxH9TSwIp15pck65bzmrQVPRH16VfSGobWYYELb7bGa
I2LgLJMujvRmp7DwMvCc980Ylzpew9uOWMUwFYZ0bANipg9HjjaWN1gJIOaq3erf
2AYEdhf9w8HXaUsDOVDJlwx861NadhSdklFHBsB8OPoAKDVRmkGV6SkShHhACVQF
szZZ20zyhfqr0OrVhlE9XgVByUtwZQ9IQI9lkO5McWgHeoPoy4fVhWJ5+CDo7GQa
2b2BJ0LD+9Rn8O7R18bCvE8wTHV8BVSuzkXMOIoA+WZ+L9oav5D2Ov/Is2vAKbJd
zb3Ok5b2SdTxCnvfh9CleLsMwMEunRvqw/sU1luH63mVWvqOM4PaGIyKyCtZ2D97
yqfdZeBVeJf+VW98MO89FmxuAx2RBjTiwX/onvKgzminSY2iDQ7P9e/wTxB1dzI/
9G5KXzrGUnx7flrj5zGvAo0Hlx0PfY7bqbEgY32s5zLY1kPTSJwVkDNIipb45lzh
i31EiLo7L3Ku/eHpc7lpRi7lTKvhR2u5CPnTwO8kUTXTcs7sdHkNxSrUJyXOIE/u
6R70AxIkaYdXIsOYyByEM53f+LuZP+LjsqVlsRZPf38LRCX+cJ0F0XK8W4Ad7hAz
aau0dqzgtv9xO15FXrfjjlqyYxHVk+BBHqNpfn5HJjyJuapeNWP9KByvjq7vfxex
svufwDkCKYGPXJx6PFZot7p7zF+QUUMgL5+N97CknmyWxNDl/gtEKhsWkaxScN4q
KCU1xyVLRJK6f1Q5EOpA+sUWw9Nn9yPdJ0FUNyV9kqC8kJmfMCpBQIzusP9e3K+o
UfXkum2xZtZfKP3RSEokxDwiV/boP1RfNv4dmG5b/XPii5jUXpWi7NLZ6TQqTlmF
8e3UOsanCHMJwzCNRDREAnyhPoMl7uzuncl7xF/JjdPU7Lwx7hvU04Hr1aqtDpjd
ZP6cDgxKU11wMmSrFU86Efg0c5xtkp1Di0ouD4CaNLCsIIWYOIlaAK0p49MdaFxo
+RhWqHhj42UwqU6g90Xjiun65vELjagpTvNd2l0qMNCdSCbHWEed5ZiTmyrl5Yqc
cavwUanI1KONdq/WfE3vGm0KNKBZwlrKjeGU6U/cCOBgkVKT/QV8E53L/XxzwU2v
qRzgzikyURwtPlI1gVzdKCVz+Acp7UhAiQgr31Gn5TQeXUz0JTAMFUEHxH7ZxDxw
bzj/fmDeVZt2EuPMWyGlWQDbFMWMjiDEPPy89rGdUZqLWrsCKkqSZ07k8zPzkij2
dBr1ZpRMGVlUxBqMPQiqbdYUbxp1b/KqPbpLtb1zruuWrGgb6WXap2bZgEfnI1WN
o89sqJ3NNn3rY1dA8UWcjW/I0iTm7hLGNhfwXw1lCTvtSXnrQ+GfAP3BwMN0gdhL
gL3Pr4u5Y/VjTEF7o5m6af4pg+PgW4vx46syOf+QaNcMdWzCxBa6BjAtRWOrK7pH
gnFNF+uHtLE3ODoHkvZI7yUXFSqvDcpdb7NH5mvbJtArHTOrez9eXx8TVTJPwBzx
V2EhyVcwyK3Mx7Ljl/1EnBlSkyOYLjFQeuZ9dSI+papxY156wKAfCnnEYwNZTtSK
sZKb1tv6ybcF2I9CNb78UBPL52KZG1BZjCT3ZKTNY6F6InMJGDpqTu1/MoTOHoPt
eXQgvl0vpS29rl1ZHxQHyCedvfysVDOlkZJX/e4iW6pwOqRXIo7lijWFhtwuOIgF
KXGPS3ucZrFuUiHA49dPthK6AgTbfeZvT5XiuhWO74ykgNpUvGcNxcKxQ2cTHo1j
iBVn8qz/y0bjIMa8hgc8tyhZJXkMoTWaGnPTN4KjdiN9UjyXIecCcUs+LiLouQ32
pjzu4+Z0mLRuDTvKEDQq5v5H39CB4itgCW8peuyZbMa4FAhOVEcCzsaK83Gl35fl
h+nhkS5DcXkxKitVsVb44efsIRs5cgSWXczYZiCWn4pZ3L/rFubWE4YKpNWygfvl
L9scq7oyI1rIfM9jznpTMFLR68WOQ8+ge9+0298xukb6zSYuyJbNQSePObJEkB4x
toStQHfy1ORu0wR67WTRlc78OLrKRxeLYd75daIT16mG5dqlirjv7CUHpQarbi84
y2S3rE3iHgbBRkfL0qAOx4g5UezmuUK+zqsk6MFqlutoCIspWK9JCADQCHoOopEz
XTtk6EzxyW7A3nxk2O3xIFj4+whGI06OxzNYk1oF9ahsnAnoyvaP5DHs7RMdhYam
ywhl5spXvg7RA1jDiDZPlXBknBpn07CV/tKAUPY5QHBoTE1SeyllpwOyg0NvMhn2
5jSdbynteznvGz1MVXI0oKbCrtNTkDkCorIETzk9hVem7/43m/LGHQZUscnKnGXx
OSn+XBV8v+LUr9rPLsJnjmjvoEidHhdw5z7ZThpNGkd2Vfa9FEpB6rpEtETNY46j
/+BONg4nXeU3ihl/ynx8sP7YV+zmixc+2T9Dvc90XiBJsHorJpEGy3m+BU11rVUf
JqBY9V4dyuoZNppAJkKM10+XOyP9w1Fx2ruwtWwb+KjJp9j/XB1hnlHNHdrr2V8h
3oImBumGPXPI0I6FeUQTPq5Ne0VAXoxzysT7eNhNLcNxF6fQvaF6CBcOvSmM605c
KrtYFMd1a9HOt8byndCS4ulRIq71GAELs0mB1GzKm/TS2HcfRSUBfLLNgHA5HsTD
OPHVFfJkfxx+NjDw0FgAI+gR0K5IdZ00ilqYXzXfPGH5cmoXTj6/UvnK5nGTndy/
fQm+srA10X9yDro795PxRX73VtYapOnMtpbDlT/qUaNoZI5NiGuW5Iu01/pfTTnH
Jmq5k3YKHf/qHI+2Jchn42b8lLhnXaB0+cs0/JqFkubYdazpqCJf5eEJ3x30cmWL
dI1gAfnZXyMM7nxncxaiOr+BVEtEZ8mB0j2EbVk61Uc8EMYlP5Gjoqe4EBVJQ/jc
7oqmWNmpQTaJpY/CWAW5QtAr2ic0SOOAkdyZi+PWWANJZLBoygriDWp8ygAaUTFO
6yzB4Vt2w0AZhaI43vNrJandk8/0q9mAh4VctAM8cCpTfFHWTkaB1PTsw9nu+DBj
F9OOaJIl7KzyfE69kwPbAUNlRzv4NuoGjkLB1lIZhHPHPOj9gy1pygUYMkIMCmmP
wMxYPMSW9Tk+HXTCZjlWYsOF4Y1sMr9ht5+oj7P7rs+fmUls6nNOFxySDe0buMOE
aP9fwpR4GJ4HPyiJB3P2+96bJDIYelU1cLxWHxCA+RUi51cvSbTSkMLgjgqAqXZV
LHe+3AU3T2iTNK7Npc8WxNxvNxEjuO2aVd4OFU+ygF/V9ZCkUkZDFMMURRJKUSlT
flepN8QswbercYleKAy6N1tQBPTJYoSy1PcweYJCbFvPGfO8ZhI/9baiMc6MTGh+
yam8LjO5pu8mbjvHDUWjtWPk8n0cPi6um8olhtdcdfJjl/ArTylsAovQ/gg2yCAC
q6JwwMDFeDXc+4LpbmzjagT8H1KlTZ569yt42jEzlxUZWgobp22RSuuswKEfqklo
jrlQq4mXfOaSi2Yxe6USJC06brKF6fAIhQ7YKBO9X+gZzmLRAMWrLAlNvYHlUqWv
26WI75qAWvkT+8Y/ioY+XgBY1ylCXpi8KCjKzPAuusMT1wrmx3IKTxmcm/JOThwO
bxXt1undYw2TGdt5p+45H97BUR8XmaPJnXCEc9rMSk0ANaD+zrl39dkCzpLFgLLg
WxGEkJktWeke0LKCy8ule69i9yV1XFZf16G5xI9BQdlWsvQjqNzl19ckTF7pdeKx
nIqYCW+B/XY37fVO2YyqPONPv7ZcOkrgPQtxnyiZ4hz0xhwvfCnHG+AATHzVQW5H
/ckFXycDK2W7yBoosvjHqyZZQI2wVDjSzhOQeEvtdA7pdyVqrIBEk/ueQOqWIA+e
9gnCsXZvWSBpkJBzneXK6agzd4pl11k4UpGBu+SgxBNy1ntJkVCb2XMOVkxztyS6
/1xxZmfiA3vk5yTcAF+TLzDhNZsSIOz/jvr2D+UoJsSO++oaKRl2Zx4m7HbTq8Uc
637nx14ivycEl3b6KMKcD7B1CAb1F+IDFKVmLzd0zELujqQCSOmUADq6JnMRqhIo
xN+3dp9XclenL2JYDROey1Ih0vUFXCdczaoJBehHLM4kCfOywR2v6+hixYishF3P
lr8z3P0nSpbegys3ekfB23C8rM3b1awqeJu/bK2Hqru1rsyqkLs6uDi/I+nHNFDP
MTZ2Y9j9XTbLqQ3+eNUzeIO8q0F5PXjcQAA1hmJkNh4LnVix+hi4WUZw76Lg+1wV
+rbYLK1W576HE6xWR2w0YeOFJK7P36CCuCykyrb2rP9lggByb+7Fz2DQWbEbFkOK
4JMgl6sGAmLfyrPWtuHkzhF7YaqhcpdM4xDN56EkMnv3j5t3ueHUQC4BIwakEkJ3
Bm/K2Bee6SNBM1MNwxCVjwVHdlsEdMPK961bIAJISZZZZ01ThIavgkAEfJUYfhde
+qhE+oNtkRID6G14p13ClSESlQlmxPf6ZezsuzyO1q0JCeFL83hZ9Y7AHLmtmpdk
FQrEg3h6PyECKv/57cdTw+0Dq6FNkX9XtbyH5RnLjDEpvQpIRMpP/zFzEShWoG46
Uj4dw4nfbQJHnKUNiZNLdCAfoB/RXn/lDtnQHot3nOZXEsbD7Xxa2jaHY1Vg8r3C
14d/QsuGjG9ULIZd1z4jpyEty3+ssaDdPYSTFWBQdR+5Ng98KrpYfGlZEkVZGggL
FWlIgkNVMN8OhwJ9P1fWTBLdVEtGwvTc8rb8AdSREqBJyf+EPeFFyxgPSuIalott
CGz+0uDk459Ma7PqlpQXZeESU2+rdPuXxj8CQ6hHiikcb3zTQIVadjJn6LkzJkyA
Vgd2f5R+7speoum0mks2a8umO9LN0JGrrHr014g6DVaI+lHsFzidj6rEZKWJVKGD
S+tKO+L75/ZGwNmPOvYlRPhNCfr1tcYU4mdnQb5lJxKyUXfz1LCyos0Ji2Jng8e7
qUD16Jt/tAyaty39538YBWP9IwbgB/eSLmJiKTIIaerPiIC+cmL/CFqTHnbxnBVZ
JAj4W4rqLMSBqR4amHfGvT43j4EV4xryiywml9hHMInc7PoELOiN4gk4BWrHKIyX
QjdUptgCpOwH98xosEWj1Y2hirkCFU9jG/i46oyRnMXoMHmaycvhIovnRnnbf3JP
TgXBwuzJcrhbnxKv1sHuzG02KDpgtkqZWncogNTn2iE8Rw6+SgbZ0cBqjpMUSqzc
mTRgu9fd5pWxjeS9b6TVjuQV1DULns6nbpaPluzkLA9JeC0CXE4MBzDNKaIvwcFn
z1G+PaKA7C2Feq4zgit2BTiHzqUfr8sQmuBsrhdB/t5yohnUn1BVWhoi1b3MA4G/
svMov5B9AaOP/0VB4xWMRITVydk/r2ca7rFPUX7WoFh1eCVvjssYufKAAFb6cy66
t2kpczLn6kECXN73gQKILYhSBuNMTSKMD9Q57bTb3AHXiWyKtK7LWV2jQ+dZSeJ5
M96MMGYKdFlvY7D+rlMFQSsjtcQSGeZ7mbwOhnpG0Brrr6NirrmOZS+UobvBQ8MJ
tBfLbyzQuhIaPnSR8Of4+LUjXKQ1y6D42pgmo+57//AkFSBCJT1lVSn37hgF1N4U
3Y9ZdmpGQ1/I+5Pnj2MrUjvA7WLc6DGNkk/bMofDdwmJ+4yl9Ofqij1ej6uMYxsz
1NpwHgFkm4wn5SfSdUdt190JYUYwTqKfmSfxrWAjeAO41h5eOKcHs/qaG04ttP43
AIzloBGjJDRAXcSLZSJWXn7QjnuUFpbNeOaw6N44MMUh5nSESVp0PrL6VC4FuVwO
ys8tW/5gmaZvM5++iF+LMWqf+LyQ9y4QjpR8Y2GPntsb0C3CRsbuTM5EFqiQejcJ
wdq7VD+5WSNbc0PCvtgJBrL+P4bgkdpgBYXlbNQm6dHZ6PIeTfixxrJKpIpfvgwh
tYJNHzXU/i3blRPSEH4T+VWzWmmrisOxVOzngB4u8k3XAyfNXERkThR8EeMc+qlo
0jm1idGw2k0CP980uDFzMXQH3cDe7ngGSeY5XFMtthujvdlInxrR6OMt8V+0/7he
FV+e2e9Pw3iWwG6AVJezoBrKvlFvCxhnAAdUm8eUizrldiF0SBDmBCyxMqUwNaT7
tUEi6YathHSwDYlTmKDpbkg0Lv1l0pJi6Jq/JAZHliBbr+8kJ5nPdBek6zE12klK
DRraVQsVMLlj4p0pwXkwu1z2W8UpyY6nkslmqGnQmSepdE1eFDL4oSjYlm4X3g41
VBR+qgYk23aQfVLkKYq0PmpKijpTpznDQHjrO8Onb6RFPub1TkAn/tVeOevNa3X1
UJ7KR4YquuCjMhMhmDL3sK5aUAM2FooRQW8Lgc052tERJs8w9RfmwLqmU8QHpvFM
EfnR7ukkTMGuun0N5iPBsXcGMK5PYYdxjTH5I8nq/MQnysFHIZ+2h9qK97DT57Li
D1cnrmll+C5VEjFxVSp8PKW98nyL6Wghv2JsjKsBMjB2NmWhzNnRnaaPO1kjnNt0
0tCE1ZMyEu8w6sk9y7RGxXUIrgQSDtBG8p0JLUjr2hXPstwaL1eSJt8NiDo636eX
n3K5FPqiN2H53KxJdT8hxjZ+HZVSWimScFxDTVodTt2zmZkG6GUi517K14rHGY6f
qHEtwJ+u0JL4nDNTc7+FKN3OzrwOBrVAeWt8kQfDaeNGv85vNmGWCVhIGeSuVelP
aNwcZgjfINxKQrDrYkfpSUx++iucyWz77jXYqKIXbTpEPKXP3V5ilUr0lMtAGT4c
8ZWAShiOcxsHc72cJdJleHJp4QVrpOzOVr6XH4dcoFlOWhxf6gUm9afnM9bSzhNr
2HWOmxeV4QGKWxtA1Wl33otoaJ4HEm0tjn/kRDWx/8ErJj9Y2Tw6eGxSMWWhbhcj
3d7553bRmfFQM7FbdCvnJbDxVYtIUqANlH027vKNQKbVRMx/EdATNhIzvbhSzVCP
JsECdridt2dpnbHEKFF135NV0L6a7klnBqIbgaJ+uiPncjlzuoPC6vzFDDrU0RvA
COAsCYIi8R6IS0sdJpJb0u3VFce4S7DFoYAl/JxMeoiV1bE0Yzd5BDDG+AkS7opg
ACwV+iPD4M1BeABTnDxTo2BA20h6hnec31Dm4hLANbrS2M/submlJzK3vyDHXiTF
TFIvyHvvBWhoo0+Otc7Ua2bapRI5u9AiVAkXMHF8104ShhcYsGX1+LXowUzzj30H
t8HBn2Xzht4bHObrzR8d8CvYorD+45+MxHv1iHE+uRQGJ2lSbxgJZR7av53RDlDT
bxo2tfve5lLf2dAJAtiDeIA75BK3t0NH9ibPO0iQtcdkr22Sy2WQ5D1p4wRF2u+j
0QpzWyt1BNav8nh1XYPWMNrMDQJE9x6Y2h1JVzh4dqhJyGJz7NNj2OpwE40/BxhU
7FEQEycoegf5I8xWjQmbCMdKS2L2ouZ4IuFqA64jp7VT+fAaNo7HM9iNgK7mX90A
HSQCqDHg/1DwKOtvtCqwekavYFz+cnbSqu9qRbSQWRKBja+5YoRoDJxlmJm+2AhF
Smx6+ArhNjFhLOngPtD9XBd7mw4aVrviRY1eKn31QLKgQR3Ws7L2sCU9rXhjJ0r/
T3utdlSfoc3bdFnfRbylxS+9oCXx0tYrKKUbfYcWa/jV3GB7rnwDX5QHkvaRO34j
9C/92PsYZPRZdIHWyU0g2L8e5GNfvGOGphQJ2mI4gjZ9lawontuNwQT/hCWTs62y
EDSgRULoZZrktYERPyMMzPakTH3esW3oyjWUlveRwtyVbUy8G0xE7862BSMk/bJf
GXvxFCGPORVP1uKijwh90vtQqYbIal8aseaMW/nJBeq+iUXYtJREkjb9HfD+jD6l
JVqvRQe79+aOO1/7gy0uQ7dyLaUf8f9KOMHAlSOWbkI4NJ1oTTt/lsWbWteahZ4O
kdYsy8yBU1U0JYjyyfPDjVib4AsqsxERNGPkcjSocIU0MeNXC9tDhj7JAtcaYJlN
g5fJLaZJrF9UiCEZB+BFwHChGbtp1QZ67fOmScZaxCuIo7h1gfZqqpxqzYqZk8Xe
SbOTH+9dy3634s6SdwPE2WHeV0SUvqotDv6FNWpwUQSrpBLV1QlML3wskle5bhOO
eOn6kWPy6Kpdl8nvoy+5kxbJuvgi0bOwEKCS4J/7bnPCCEZO3gthrgX69uu16v25
srU8/f4+XfBFGxnFh7IGFLLYLA0InjIF81C8f74DQhU4AFrcVQZMRi2kfvSa5Qau
r5/U+Jqs3480AZZ+qcJ8OgrWKIGfPwXviDRjFGCc7tFSlkI/znw2XWVw+0Ct53zA
+H/5+1+DL/TyN3rKwucH5/YiXb3QvlPvC9U7PJ+qsDaXVqIT+qFt+c2gjGuklWJE
s6KyxnRqsbEypP1DL115PmeOQIeVoEkWMIQ9yPIIad7cmzWETjxbyh2ph5xWx3jq
uUldif1toCFeTUdpzd67Uul3LqxRj7lJ5jmCqks1bUQ0nAHpsxAnZy8AiPVD/uYS
q/SsSh2G2pYmjE+6lxbU+xTYsOwXoI9/5gIyXz5s6SUH5ZZJA4xADyPuQ7OrY7tE
WCcFyEWBRoVeNGOKM1cHDbpxzKI516krZ5ieLS8iHMqITqP5AOfq5qyjG2+zj48B
rgHPPOCqKWri5sWfbFRyF4waVx0excxqOrfTOUwhN25P9ZAkOHfo0IZMF8g5ks3/
0aCo2NM8RT/hStiFK6TjlwUGf/ngwvlxtfL9oc9IALtFA+PU9nejZYeSUPQqsH/6
AM6ahovArlY9GOY4eNMU9JZbKtoq/Z9nhuqp8EOpsIT/5/JfHAHxlppmGqVcXOB2
7V1YXJKs/tIMW3ZHZmUqHnQLLtW0f4heldqfUws/ZIShswTbxbhjZtwNQkAE1Bsf
PoHhOZzRyr2OPy9wfcvFOGmQrzwfELfRl5Pc9YVhjTPrL7XeaNFBwN8VshUGvGCd
KJyA8+btiTIZsqvxz0izTFKCkyxg+FdMMCxS42rVSY7iiaAMy22JymJ/4wKPEW1j
dzQt1oiorkMVGxqjYVQ1mAe7fMnSBkf5Yq++52RYsgV3MZof5ZDA9Pes085IIwiC
xWVcb1goaESmwZEVFz39tmpxpC5p2OaEYj+wrU94BM5GspIoZwp1PeBANW2H0/qz
taiHb9z0/Dfry/ZrLEVti/K4UChGwYslgqyUpgQF6jHKE5tpUbKMO7Bi3YPTEn+O
tlwBjyLckmk2HUgFBDp5gjv/9zJOfxY/kJy8Vi5aNMYCl0Ox/cbduzrYtv8BUgVo
emK6bxex01eJn88imO/HXJqYALB4IZGfxTepMxr5LdFSEPHRaMK8ViNWNhxFMl8O
nqkRMLtyeKu3DhojjUYD/yF20dj9HPXAwAJjE1rsz5yg4I6NOum6zPCpXKmytBKn
0L7CpYp4cabEJtUFIcsyTZK6jZfGib+/iWBEZhz2CwyetpDaZkgtuaE8yt68QrYl
XI1U8r/f5TSX820/QGStYNLwaVHkPZCHlcbl2/ZnuU297Iu85W7RzO18FgGqYBg+
ltpbmdHA1nIi/6kr2tmAYrkmahLesYW5h2LdkkA9r4m5OgeX8n7wMe8yxKJZ55Wl
nxMoKRr45SRNO+kKNbGQ2pmC8eY/2mjzFpayvpFqn84vZNbJ/gTvOITT7qdyEbL6
e6R/oJe9Swguo0aQi/8ogDjtdQnlomDLRuLls6iftnt/He/eWHVCk6c0zz6yUIVO
RWUXdiAbMKkpyQC+J/uhaRJurDlOwt/nLTutIqRNYyJMTU5YSXSFFr7O8VLscXNl
8gcDBTWtvNQ+wHi+A0twMid+ePsboUIWkVzu1Vy0ZWFCYK/aty5MUuIuXiGn+f5L
Xc1KdrSMMa4+y194zpxABoIhgAlvBNgUjhttWmK0BWwgxVtotm5SXyw8irSJ9Lrl
mtcK4LK255O+5PS5J+xSk/T4xOAaUTv7yHEBJQpDaWoZir6NLaGnG0xpl8eDqcIr
Wvxnp8kiLevnx32SntuX+SvhzXMJeM9oqt4iVfrYS60TP2Rw51yyvMV0aQ7NPqKp
lXpdrtRvBqM9enzHB8hjM/x+OeoZYYRler+oSJFzdocBBp/71mYBqbSqV2nwT2p0
B9jw0X91PkTI0diUcHNEe+COB1UbPEXw9TbrxPgojbSTjMcnRj/GqdDcs2ucTt6j
sIvaQGDTTGaYPm7miXOcSe5KkJ/XWJmhAnXc2IFY3yR0cQTnDPFhrr3ohO59tomJ
pHJNIBO+/WqnHE4WePttAkeLS8B0MKvBdMNwlKFeRHIst1h5ZGPn82tBmNrsDu1B
17N9PRAOcMCGQT6RWEHNTD90PaDQsAFWDzUelK1EqiHJ20e9fC+6X6c5XcBqhe4U
sF1jxTaMdrLKp8rlVqJYoLjsBAhZB/a+Fv9DG44akI1+gA9KcE5g3lINlfHB1v8h
1G6Xbt1kX2Py+YXAmhwUQFFxapn/G+SJSIWWbNKlX0PqxwLXO0bWGzK5E0rIQCdt
ppnquTGWQFICg+jKRCBKDRD6o1i+mg9ogRg134r31moT2abAPuL7X0Mi67kc75TI
bRYJEOGZimDdOJNoJrzV5pQrQym4IxoP4DU4AH5+jDNpQi0Kh4CeKyPTESZQia5l
yMVoTd2ZDv0VP/gTRzGqqcFFDYKuv1nmUJzf+A0oDe0nbKJAu/Jyyz5uMvO1xkgE
zQtLY9gDl9CSBTNrJ+g3sEACTh/z9EY6u4bwX8ub11PJYBUmwH+vJA7VjZwygTo8
9DyPjh2yulAf16oj0utWKtU0sYRA1GwCoymTgdnBM+TzkK5woPxzRe6AaQiko73o
+UkdzN1MqYTVY94iYNJQzGiEHyRYk0S1x07r4SJBODFF7fS7RsGTuE4HW2C6tzOK
ES8DbaqyLogq+u+ZY6dFf+sUuxgQdhzIhnQi5779hXVwCaXmkPw5IZ8S686skIYX
uhqXZBRESo6LeK6NOIQxlGfNcVs7cfdji4VqeR9CrzLkNGkcKLNy/zYT287EKSGI
9ltp5nJ/C0zq0cZ05o7bSQXkU6D6caDT5ulZarXbuyj1AyNYVqlVu3H0T+j2HC0+
lNbIHqFFArH16Di7ypTkhuOdOR9XvdjnbvqXSZbtCBHTLI3RiP9ZPChV/2RHfG7n
GXYy2pvO0UoBTYwE4vpyYBhwCOb59yFg3ZxvWGXHF4SeONWxO6HxHJQcEqQHlkJh
0+IPh9GB9xKjXeRa6HF8Bu2YFTKelq37HayX998SVeiML8w0Fte6EyXE8z8+8qwd
fFatBcIUdwnnwV5QajZgaIHngBC39M7FINgSQeeEYqD2VahJy/LxQEcjuUwqF4NU
JJkKr6xUxWtwX/6hwPMKaisvV90Gg0P0VqPc2YMXKOAI5TM1KfO9VQYEcd3Imko6
Omg4let6dVK1gQYkjK8dLIL/XFJQRwXkQX5vy0y2v+TmQGLiVyU9ew953egmK/tA
0Jr2wQQqJAtB7DZ2wTsbejlVTGpnduPNR/Tu9I2IMxcWna4+miR9SIktzr1EuN0Y
vGfkyumBexxR5UHxozXip8oxI4T0XE+s1z42vzXr/Fd/llsJq4zWmcgS97uKOxED
z4hwRHv7ok91iPF7iiIQJBSXu3hcrDkwp37U/vp+fVRIVtEk5OLhu+e0v89DV4sd
GPNsxiTm6yHzAC6AFpSNyAZn2yICurrOFgTHAxQC7CBzmNCXfjGMSXjZx123tlQn
ey04hp8yxvgNLFC34H0pMnBPtL8fmeKOi48/E8prz59/Hj5qz7bl8Nai9ZsEFy1M
sJfclNpkPa5oAxEP5tXxtoUaoeodbz1AJ6V1AqtxsCPPb1ZX3O2TIX2Y9bvDF+Q1
sfIUFx4vW9n1YKwKcS1x5hE8C2VLNFfu2/lnq0g2DT1R7hXM5lMp55yd9hs+JDwd
WKuZojHQQRDJ0lFO1nV3IFmsmT3PfRpfvL/vPBkDhoUxyPGaN6xXvSQ6xWDwigBF
MAsnmWGxdFRaEyHZCJF4JEkdW9dbnLbiJXJDojra3ZmqBpzBAMjq216h05OGorD/
gAuMJHFFQQd1m69TDY5UAE/eF3djPK1Ri7MNMPZ21ZMDWM867bR+HkoibV3m+c6j
n7oC3tr0QHl2o8jWch33N5ycsu/2W9AwYBaGwuoV5UQbMD0IaBZh4tAVe0RWBpXy
doNxZKwrZawmUJO+sITmsj5vryyv6Aot8Ayn7Zl7UhsPuQHOKlHxCddhp7O3zTxv
Om3ETZHvftipgE3OI84e/RQj9W2AdgowEx1J8BbpWo1yoVEM0zI7rBE7x6h5RRsA
bdSov3Cnt59slYwDtrOznuFql+nmuq23M/NV/NoRUVMA27Xl1UIk9u8IkkAYBcDY
dRsoiSQ5vua4sU4W2f19qB+DKR/hWn3s+zTiLABCKCNgazXWeoZjFbHJOJC2H/qH
VPF15FK8DzZQ5vX7l1qjAZJCZne4O4TjQz+4ETuFyLy4ljlhW6X2ucf16nOmUOR/
k/eWQ0f8iZghOP3eVcInSPBanpDF+MOuDUO1BMyP/ikrewM0hBmYns3OZp0CJxI6
DA9up28eZcZP/x+emiY0oXXnKCI1N/ktv/z+tXVX4733U7yBmTCumRGJjwZ9FrIt
TZIBSlSvy7nqya/8cHcuSQaKVQu9lZvZErS/uMEUlk0lgQrRdpAvyJP9ddX5/hGn
EoOfjNodcBpjGf26+TODQbm7FGlquU+By8unQckQ5i4H/hovWqgCaS7ELj+1D73I
qJD9SeHKybAsXqf8u5vmcM3E3WS0n/dNeJ5DyJ7et+SBX3RydziCGMqkxkgKcozd
qCuzs/iak7/NKSa4WlHTV4d4VFD6iAltN0RxDDYlhN/1EJ5GxQh3w+mpgQAguoU9
wsidMkMJUyYFngwQop3QLOqF3J2uNAH9GqLGMdrQc3Gwx60l+KbHwSe+6jfmbjhY
PpZ1m4BFLH0Qf9ZLUm3aydoevh0kyKe72BpdeTuQvgbs7XcfI17EZ3tvzF0fn2md
ki16QCG/h/+Rwih+j7ay1zyEW3ceHE1NWq/dA659M3I5oy5W6uEM37Svfz+B3J1l
2Y+HPkGZdlCKL4Aq201rKbW0vpMLV1xIAENWC11X5/W6oMk1r4OH59KKXN5q9wzU
S8qecu4wOBetL+BHHPk3y++m8o1lAXkoi7CG5rvgKN27ZjCLae5ndEFrCRg6OjXQ
loWTbyPZTLdLOqhJeXTRpE7+iuc14tqD35MnT3IUytbJQvVMNhyp/FX56YF4i/zQ
aHaqkD3abHgJmOkvshbSUrXQfGm7TyADy0zP/lfDkSnXigh+XWH57+W0y6NV8hco
oyiz0+7auVtHBO8tEpEsWdgt+Y+I0ZaMX4cg0PfyAzpTmVtIHaHofHyCHPRecoT+
HEXL1fa1OfaqzszseJJVbZ3ouwHTTUZWQUy6fe4JG2pzn8Js7bS0YtpLjknbcB2I
Wb7IM2r8o5guk7UVz94zTrmOHoTJXqo2DXBhHYlJCox4GXVlBMK4PMzJ6JhgxfyW
L0wQuQ7keeuMqbPPAwZnCUAx0IJV7kX0lRd1d5XaoTV/rK7joF8s9mjhDwE5/6Ht
Py+n2hrHEKkv8gHKBtDXXOW8Rd2c5a0dR8rh3hJaBKnpa+wa0kyz0bFXJWTi3U7l
tMNdLbI+HnNGyAc5W1ioQxX1SIYXVMTINLoTr6TavspTIULWcRrFtCNKipRAhfEz
0cMzJkjzaTl+ruxeNRXT5nqZBaQ7M6pmXb15+yD2fYTg5M0lnFZPVx6wVUr96Vv9
d+kwCsy/qvmFU3xXTd4k8AGSmeTs+4DG4Gx7lyjEfl6mT6Fy790RV3ACTOAjAkHf
Lkh18Em1HNIrDx6OE+tM3Lwf6wwkEpFrHWfGV0r35FaYivQwTybJC7H6yTIkH/v5
0SHKH/wXtlUnmblmX6Iswx9DAm/gx02yfCXApo9pMx08TChTS9mBhkZzxYeEjCo8
lEU7B41SVVtEoewgt+LR/vKalLVQBS69bzqhW9E/DGhb+ZweUZTiTtHBJn3bmABA
WTrOs2tBwnZ3ws84wlC87e4XoPwKErsyQ3uGqaMx1kywoAdyQ4oyvw5wGPZFa4Nj
YXEp4pQ3fM1nN4a5IxnlKH/yitK1T7OH/tgGCXaIJOHXv5P4VtYsuzcLRO2kdK3V
LT4j7EFSZqTIeWTQk475JMI6OCI3RZaTSqvL9axjjS4tbwqPMR/1+aauPuOe/e7W
0Wwmvmentm5bIeBagWWB6zlWHmQ8DZgTY5pulVK1696oF37TFVNKkGhCgYgQnn6r
G+pk+oyy2hzFL/WsVnvCL8F7EAVCzZAOzrp3YOYzxdUTRZkB1EyF0MAYEoQ4THpv
KRNL97hwZlG/nJW86LQqpOxk1/IrgWDvQlq/otLBIqz7kGcayTyyHKy75TQJK0RV
CyDIe52UNz8bjLMMbbJVs/BybO3lfCu5QrGf4j/LhJE/AFVbueo8jnKMxYPCQQQT
KAvOdF3kQy6NUKrWSM4BN8B2U+BNWu5U4P4oCDno9dwU5kuyHzf5zAI0sHS4P0qH
F3QNSrKVfYbyQG0LSjCpXn4UMZ2uXSthe2xcRmpz8xaJybsgriaK8B4faeDfGYMR
aWNUQdekG8peeEoxxvGmAh0XdHdVqRF4nnwS0IxXvwn9Ig+v9WsqFJBEHynnjPpV
kyFxuHgkHEKg0H1lCb0wld6wLLPgMAwzCXZOxh2y4q14Y9EWyOaAQEIflWn4tJVL
5cz4jCWL4qEuZ2EhRlUIyFhjx80Z7uRuGyUfQ0TtjFtKjeKmwax/jQa0aHWemz+4
89hFwU3ZhUmWj4ZIRoivFpigshobYfKkD6ydvHSYkBwRCYbhcatgi/EUmaYAj+PR
BXM0f8Y+X7iUuq9bc3I+p39CoSxfjDfi5bfdRfPZxHbwcPrdnoKchanRYKZwW5Pf
KThBRbrRGIzeeWjNr3eWOxecilLIDYF+NjXeODonfWLP0kbUXQtLaoq/hvJoM0dI
KOYYHTCsnG3o4POrwW2OHMdVzeJHEgNNA3YfbgKc2gDPcpcw8+a5ZUnJntCwdWMy
ePgbvXrZ4+o6A2SiZp2HEXylYGBNweaB2sBCV/SGLhy1wCt9v86q4v5EdMsTwOBN
699/ZAm2VFbx1IyD39fhZKa7+Zxo04dpoMpQTbHX4db+ZH1YvOyMxE3Cx0EPiybj
Tg/B59qJF9rFoucNIwz3aMDTCrGLGi/cbQJAegd2QoSfpNGzt+XVJ4SzlnVVx6U0
j7gRZVwCmYF/1GqZ6l7szk0b438qQ3YJtJ2kliQ2ULwMiLj72dQcHep04hXzKx3e
bTyR3EFFGpPNDao1dSouGYwCNEuzLyPNr79fK7av0aJ38WA53s9AHf+KOupaOTZ7
uuFFAzAl2Dqfink2E5Qwz7qBYVTU+RN3/HXqvP53Xt8zsCpKwudCqEtHnPVI8NlT
i2x+kmt9uCuJjVhmveuxXA65lRXwixtIZK8PftZeclCmuqMWHJZuT2h5r2MnuDJW
W/4xQIq+YAIF6imvldju9pBbMod/AWJexuPBxIOlydYSOXGr9vothirkVtzYle0M
BkiPDXTBalrAMVIet3sla3yxNygNBkfaLPV79YlKzbwwK8ChKPDwRnAslZW5mhVD
7ugPxGHjXCPnSX9bdFNvwCAY8NP2/SGknV4AheXrfmW8aWTfX1KlGs8yvK47a0mm
J72ro6C8qFBNuqynaQ0i/0EEuJBsK3x1zo2KDUpgV5L+sBwEyUIgv7cX3CS/4GT0
0rx419wCizXJ7Aymzy1VJXpZsujXQqk/urYp/xjulmuXXIxW4j7q8MpPmqxo7rgm
G5h0OQbWHrkq4BXMSvYSZPN/pHaUvNvsDEcY1xHEB0/qo0B9SMYYnsGbbjz+83NI
c2XJY0+28Y16K0lyEkEvU1rBTMbSjuhXa08lb2vgjPcqCxDxidKRyjM5r5Nnw51b
GhmmEAUSin2FDNxoTb77ttIm76ghcqYaAY394vlkV1GP9uu9x9g9UYcy8MEEb1Um
zGjjEQmfwZyOUM0xmjnttooX2g2Nz6E3umQevzTCDArrd7Qb+3NYGKUuFQwJvq8M
9G4FgILFfU831elUCUJTjD+mRwvh+BBdua3NMky/Lbv5XBOPRXBELz7DxYO4H62K
odUIcbrZ6Go/Fktst6eRahVQslGKpZPUZPmjh4pMAa4SbLx97hNnQNQg63czICLN
Bcfz5hKcfAKcWmuo2enL1zSod5QuxJPkSFdQQePRldSR61cqW/3E+kOB3mGCJBis
/aFoCjyoGMmkHOOfojtuuOAL24LzlqASO1n0aMCs9Zo5xu8n78jP/yXnaA8+Z29g
NVV4fA7us0kMxy2VpwmLQ0wNLPrJRcU5WKrdT4gNb96oL57QifletAma6ArM3SL0
3E1hD5X8jKIQc3ZZiiKmLV0odBMnu9q21wrP9rmfJ1EYo0TVfSNJ2sYr4IHi/8Qv
VQ1Om0PrVYgNmI5tPS7QJujY8MVr7iyi8jyWcetXebK5n6QTPM7ow0+ywjR+bmvI
E15RXrdc22pCqXAZcy84nfnjLwoS0vJX3alt1F6l4OlFUrlqSOt1eC1QkgkROKq6
5VRWei77Xivi/KhXdkigOVMqOX3JuEf/QFGGO2yiWVXB2FyG9YNeaR7VzC8UrBFf
ayHrvit6ji9cDowbCAHICyJaw6lzBxj7glPKIrL7r7yTZWlihQ/CqpsCBgL7xETD
Q1cEPFDAH+WHTIbwYPM25da2SS+D88znGHgO0ip57FV4CVtyT7se6rTOdsACvLZx
x4VoI+vcc2ofhj5BTLOGTewMgHPojV+3Lpd4gZVp6mFZ4z/LBJPh5dpqER1grtvG
m/0o3FNu0nMwUh9T8ACaNTi9lyVu9c04DyuDLDM/P+My9zESlo/R0jfQhrBHViHR
qU82FT8B7UOIcA4mx+ypWQ6Bfd8FcJdCcf4KcLxy/pHNBbALxuHKbM4qnL/eKdVe
wwJi6GKCKeb6+JmGBTL1DXqnbw+LNVyojB67acuLoDXuwq6dim9OmwQwlkUb/rUn
QQcar0J7bRZZNTjO3iNC6p6FDx3NuBQULiDAz2olfwMiJPva0PedfoAckL1PhH8K
EK2UtHM0n88vUQhmTC+CUvTCu5N4Uto5cR1KIrcGkSt2bnF744zp/d0z8femBF4P
/DOHde1UJ93FrPk5K0qULc/xrP1PLIgM23CZBSuO39LMY/FY8amUZRRqw4vcgDEJ
xRnm3v+GhgrNOesUwjM/pERLQ+Llw5fsimfPe7OBpVu3BKqv9aD3jq3aLVctX4Nq
q7foanAIjrU82jAyeB+05e/KI2erZ/rdGhKmXUGul5BiSEqG19gxLvwHrqKhfcv1
Hi1iwA5xE25EYuDmEMRK8vZKGDdd4UcX/ZgD4NStzR3Sksl9GO8nAECpLA6Q37F0
XVHBV47QSnSGJ9h101DyrXFo4knZFx+OVW5XLtNwL8wPvCMTgjeARo0ryiz2mY/s
ST9OJi1X3M2CXKzc+ipLhqL/Rskg1BUTAq8cjs5FTmwhWLzof+UymLC3vKM/vLQA
h6Een1QbLlFBLyB+AsX+enc7VuhdczoN+W8FmObnPR9gqF+AultPjIXDfjgWe8Bx
dUeMnJcpNlaPEhNtT/CDPMWFa2TzV+YsfxgKjaFp6TaqLMp2ihs68MsWjEp+ot3U
0pjZlafeFuNympVUyOl+CMkC8HAxDGo/1k/T6flstqxI+M5x7coqhZ4M+cKh54Pg
dCE23plopG0s+iJriNgZnlW07epxN381+BEENoFVHLMZ0ghc4MQjsRQY3tT4bWPD
fJZvIE+jLpBS0TXIJnr3uhm/pd5/4YUmfOiuLVSTTK0TVTO28etwrv8N/I0GKfLJ
IKzQWvyCfkKW48lWpuyTfY1BB9Qm25F4qUxzVAi8Ssdm8YjQHiFb0N1bM2rqiKqp
I4MaRdWF9DklCKEEvCp5+DdC41OP3/iQeWPYBUcy0z2pAvlMo3AN067NSgUqTArq
wI1jIvzpvIuprTwkWgMf2W4FPR3S9uHCLk1eSC7RfJzdUKs6MjRYmQdBeT/KJS1n
uX1nHMsV2pF7wxPXShCTabencvRn1Dx+y+eDv0grqm9cY71DthWMqzvHqPgHTJNE
WIzVt6EQZDFqjIhai8LAYqaTg1YQOyhVRgKTZFq+gb9bVbI7bLWX4utBfoICk2dJ
bvGf6NFXeCgLNNg29v/tD+nZ8skgu46vOUJm8+R81Smr92j7jYBVpkEORFnMwszx
Ws0AvBTU6wcr/qaoqbP26aIzxggLqI0nNjUz/AWU+dDu6xrjAfzz0vpvOPi2S5Z5
EXAiX6kUTAsDrGajRyUvR9COXKMucs+XiC9pCys+3Jc5jqzpY6QxWq4O9spZOa+M
LuEUvOY9Wsa/U2uIf8nrUuwULpv+ZxNVRcrNlhI01evhNTPA/gFmb6C1is79SnIV
iDIxl6yuZawlL8UVjb6gantoiZdMLuT13uvlkOQjB9W3NqNRE2hUh/IU5bAnHiry
0b2QYXA0Qq9t4dXTjmYt0IuZt5f7kgeypwL1RR1vk4UAlP6A/QdFIUaJNXCU91Zc
JwVwVsHdfTfGWldIh/JxF4m1Y7/Nhr0Tmk00Ym8ncSxfgxzz4Jk/4qt7/NMJ5hEs
NfezbKO1vNL82/PlNWVW9mp7QZnbDC5uvgEMjdGEoq5PBbhkE+L4Vgr+hGuxqIC4
/4lZ4abFMn2/x+x/4pa00wsXRDDzczvlIWj5AbREovg/Rf9uMxLx4JIqZyXB77BK
dxMTj++0Ff1WQLnBOmYZWxCsVbYp8hM5Q/0EdjeqA4Y7ANcfRygZbh0Qan+rnuQ/
VkDqv1FLUpJr4LUPiL5ypJWyKQ0IbIccaS2V3qn8wSOqSeWFCcM3sOzITJ2HTrTv
8rvF6qWJmID+KhDFL4nePGGba3/Lz37ZKPG2E5bhPumLoTmfXBDAi3AlImWRdIBf
WT1uxhGuuJIXuEzn7GTEm+A18VQHH3q4HF9czYouEVFvvCx0BIO40/CspXKpIMP+
uZm86knYFf8LzKull7QXunIZkDgHe8rb5t5G4n0xy5N/FFNN0AubmGtbV3o/a56V
nIBUm2IXw+ZPj7JHYZrY27tQ3MBdXNzlhv5U0wMr9KjY+ugvOrkjEPCjAcd+aOD6
r5Yd2Xn1aP+3/Kk+R6qUCBm4/S/ukdxEOiky6l83DwTCIsx9szQFxWN+oj41QWtW
PjD0DZF/uok79KLiF6ve9ShOKuODm+LyPCq2HGlYfP/AiPdJb3dipfJJMoqqRbCx
CHIUcezR6bzNot2AXhSTqsEjlPnjTaXCmS+Jcz5hDPVEq3RNUoR3KWvzodhjsRAa
Y0O0TqP3ChFDFIwt0WOPDyPpBcC/IfkiC9Gu9+GuhypowJLViptH6hlrcdqQr/ar
Www+P4VyjySE6X9+0moGx7ASn5Dmre3tnZ+zqyC8kvs6sal/V5y7DOfzc+t/qjTK
6EFhYli4Sj/ZkpbiQsrdoATGIX8PGGqFQlAfhibq/TggARxBc6F/mCHr5Cx/laEg
ayb06XBKtoKTXGt+2HTI+wUYHdtR9hc/79omJhQxjH2iT76hYvO3oYdzlUjHseuc
ChfonjW+eyXDSf4X9Wmh3TRb6UVtDHkY6rnVUIkQmQnSYbg6d8T9POhMWQ4fk9YE
B+852jaoFX+2IeQFNP4VufSjy0dB+EPtsvmSx0nJifPAB6nPaKe15OnPexkWYCbT
EFYVV6CxMRrr2UpnSfaLOEF1N7dlsDWIx/mz8nhLaV+A2Iozu1aFbDgxFjHTnZ2d
TgEDIuQnXgBmXqlFYa0EU6f4alf0O56paS/xQVaqwBLmJHn7zd7XxVTez8d+c70O
2g/92djs3RvxNjWztJO+X246LHzoXSDuwhKiy5S/ylp5qaWDl5s+UcXv9TAnghCD
gRNlLSDEHpdBO1PbSwSpkuP5iBeD9Hf/qKp7biA1GT43tKUKofJH+6rLk+sZuBjG
3o3LctF2Yq40YqcQCXh3L+gzzJuKLUrqluWRXhTvmYr44A8HnP5Zn4JKHggFT9p6
ZMvHXYpCZaZ4Du2IaTUuOnO/YH97F4BMaKkpekgYhTkAgOBRtnOtQaQqavXlbRLV
2ToNRAa/MMRNcwMVxoLZtuDnLC8VkYur9QQ/kbg/dSAYtVKkmA6t/UdcNlqEcSjC
3Kl/ZPjUeHlKc3Epzw5DZXOBWmM/YM9bc0GMvHzS8XnETrb8Fo7RrOG34UxpJqpv
eSQ1fDEGUyfCCpFCpGeveWX+7L9nw3xegistC9tJoMup4fgAgG113rK10LZeEMGk
VqcHgcgAIk5hEOvtdHJoChhTgOTFh0w2h3xKtREr4vSmloW5AQsZkUfPj8S4OrO3
ophH6fa3+WdvFOhnRY0y1Pn3GhlSbDDK2u9HsZYjqT12JI4O1IfQXsqpBnzDWe8D
zOsIPVVA4Tkq/sbSvSFk6ZsXo7Cix15s+wnm1e3hk4PLgBqFrI31pvQvGSQN/vlE
IimlVMcziuSCG8binoZRbm3NEmiAajvkzD9sH5Wuct/BXEyamLewyTTKiEjqoihs
TRlQ9RBvb/U67xNFyYOdSOAVs90PKrjWsMOWLHo0WveXYFnxmf7mZiD74WAxgHWF
LS1XR5R05V5leKhPLw/Yg8VQfx4w1qKdf0yKnFWtOdGOu1Zq1i337t1j126KYpPr
K13vR8Euf/80niVKXfHscsBzZCdp7mhymk3F+LGpfx8jgy0fi6wb3dBzllrwlSRQ
ncBYxWCH4nTsM3omS/nWt6vjjOtD12B/aDcrm4K6D3vfr0Fas93bQPiElkpeSb/p
tXkjW7o9nVd52ewBBybMMt41SvFFK+9o0ElQ8mDVq/l45C9VhFhEmbn0/FD7ODg2
ZLacCk2RV/Z1en8n7tZ0Vi3vqmvB795tPeHKR77XjoLwkzFVjb4d0uwOMZ0nwc+N
pKjbgoikVSO4Dqn0AsU8Jsf5ZO1Obz3hcI58HNXqwpCCLDTxzKv772bqCaMUUtxG
0f5JHdakXWE+ZeYtgD/QHEfsLyD+G5LNxGGQfrv1DT97q40eQf/7DLfVInrMgzGy
HBfhrmUjFnFhWbYZ9+7n2QGwEQdEq37hx+FZRtpAelnEEBvnqVkSMNrVrxCc+EUb
QEKsXbTWuRO57iceoTofBolYKWYTiZ0n2knFExZPuE4aFIaEAbgfwHNeEes9XDF6
wTOmElmfLyXSG3a/ySAIbGZDGZX5400t2ocx/uVcUg3HVTWkWKJV7texf9TDr66g
UW2qC2TSKgcThVxQuCOs2dY1N5NM7uwkiAYFP3kTN2eTIribBMwT6OF5+J8S0eFl
ZZTlhq36PQ6PFmGMvlH2BQUYMio7CQr+N4irugrt4FIx3P5HOTYz3LeB/a/OTJRo
mShxnqD/iJuN9O0oIUilVDz4C5F/twEfJVKS+qIkOk2Cq8FpX6gCiuBjlYsT7P64
kzTqqpIZLrJxW3g61ah6/27PpjYCjVZsILF7ktjDWjZmes8vIsIasg7sjDUlpcRB
mzZ8JyEWdPi0mGlRbEEXJLDAMxuKflbyXiM5xrqK+pCAqL/cccGitTe4Of+94NIy
oHzd8TKz5+Wkqsq8Np4uTQq46a++Lnqd5fqLmAQkfzXu3BLZxSdE/JS8uIPlLEE1
0Gdsr8oMm+CaqNCYnrnP7IZxIYIFiZC9/ue6QLIiSDPNhUwjY16mu+4blJYYq2Hs
JS/KjRGih8fnsqaQxXp4NfBM+Q7WCmSyHcMPr4dLmaTiMU5g5Zl7CtoJ7/vSzsfd
CqM30A/eWEszZpZREtYf7DMZdwOhNVkF6/ddG7GOKpec6IfKixcVYVTPr3bCdTdq
InR/Xo+EuPwUQLS+M7mc2IFdGhqO0LI3tB9CzVr5XD9hFajMaKXPyIygZOt3PyQG
jUWcpxKfrACkNN55wXmZg+yxeiUsyiLQLhciTHMbNHokhkc3Maoex4bDzYG8+TaK
22vQ4XixH7irHVrCisVpg6ZIxWPKqINaC5PioKeAgFatJsIsP074a3960Cs8jxBI
LmYSMp4C0PcJhFoM/AhNvHXR/6N1TMaNw6Ua1oazov08RPeNVp3fKvOWrPAaY2sN
vcrzro5Xkg6BsRDadaKv4Os+D6rZPqPCAB/NdXyOQhrDUtoIGVeLb5eEQ4Y2X4ym
33BrrFZOTAKxskixv6ZHtMog9rqZnE5yTSrYlARMLooGHz6cR1jRB+ury8BfhsS+
m8oqhzWCu/PQlchaYGfpMSLX846wD5e4Jyx4DAtkeMaU6mdkOoP+WSnPi4MiRBRN
qtVyRuNEIQXg6k1EpJxTXxqATbsS/2ZM4EMrhhXfLoW8kQP64fdl91HPtCKRpNfV
iInKJApJmlTquMuKe6eKBc6nJoD6TnARgOX/wkV1jTkL8LFrox94jRq4QmTG46Dg
UWIns/Z8mUlnsHj6r37DTqSjT0FDDOGaHVwq2Sos/Fvvfvx0/Kmf0+ylCrPtbCtU
YQRxugmIlOvKBMwxP7SNOaJ2c5muyZR8VXcO+xMLpoJEwu5YadqRVXyY0Vlq12Od
azjHqO48asmpr/jAhswNoSVV4/rXH8N+S1w1GQB0nMy0PCgAWqr5w8XJcRJ1b9Fm
FqPioEldEMpA66n3yGLBo8XvoG9HggJWAu1rm6SpD7L3248FEsmw45nTAsnfU2/X
iPMGQnPbWn16OQAU2pGTQFLa7CWoCHL5tfKDTjF/Y1OUBpeJObPGARi3Cydzgy4+
HeAClteZHVAY9IdD7lh4a0fkhO1N76JqGNuD2Ldil83dvFeHsSDZA/BVdk0jD2mu
w71kVe18ZSQUNdp5E6pJIbQnD+RnnyMz56fq4SkUANNGXz4dYlr/ybFabUhUZ+Xz
q4He/rS2myG55Mh06fLwJkrL8fMNkMXu3kG6ZJpCNQ1xC0sepR5JYuj6y5N8+mJz
Q/uXfpub5dcTBuHUM4vVGCPd4zTEOwMV4wtLpfwp51P1lOb/duGtCBjE0UXXHH02
PLahCVMTPwfeV4I4v26O3QGl2NJ+omDqvJ+twOClPGQHqKwkzVxZEfVj+zyCSSAq
inKq10wdi7WwpziregA4N5BzqUxSBd8W3IbtAaIw3qnuug7Pc3HeNBBVhsAnACbt
UAmFAJ+iABG9xjWMpVoHeYUniQY82LiycwGvAhs4rVjU3JhYi6YXa+Z0QJblTWkS
+0aa+kuXP71KyPR8WqOY9z3Kxrxxgo7ZloGm1GHd0v980vBmhkR65ueVvHCAKyRP
vAYQ6mxjJgxTbZHeGT3v/dTU5x5sWbjj8l7ateQJfBrqw/W0wEXNx9ou1QnGzegv
Y6mGMtCJTGA5yRoEobRXZxJRRis3zzwnM+FMF9+7cHdyPTmUUrHp/kXJfLVX3Ho/
UPQTZM2bcf3tbhc1mkVoYYkL92f7IUUZs4cCeGJuyYZZChDqnqtWtOUbjQzP3Vml
CBAuS6CfLfKAj2ms9XHeiPD+WRMJCCRWNVplSji8Dqg8GCREiu/6+A39xaJAAFWh
UgpTg+E443bQtLRHzYlghRG0BlsHW+l5Iw3SbADENQqub459T9VPScfke2HEGW9I
ixtWU4y4DG2hlgdqizlD8GZQZFCyCaITITNhcFMNX35i7ORKZjsSStRGcAusPEy9
IsBEuPDCZP5re/JtrFHZ+QdsGFSXBakLHz0iMVd3CjvCNU+g1JN/Rv+mnxgPB0uK
iBXu1PEbEL91+vkeis5iIYaUs1OerSSAOMWktAjldZCOMw5RZBT2S1f/S/OEwr/w
UdIp9TI3n/4310NR5FNdoRHARd4U3GPJCLhzX6nrhyxkIDJrOsMxrk8+ea0DBYWG
9vkwepmI4KozPeUknLhpr+WA2sygbiNMiQPf8n8jwN9rgdAJPmMnR8PCyrkdRb5l
nhFIgEuaP3yR7QPsd1u3J5B9XWupb/LW5JOpkjkLqX78GN3buvMC/cpR00BXu0q+
EEgfwIpRe28pelhiVLscnq0ZhCvVC7KkWp1undrcJzIzeI54qQLfcnxOuqiwz9Ji
tTLAUnfBQhArW2DuONYzQivv4cprAjv0/fEH/HykzWtTg22Uv6Ktj4Sub7bu6GTb
bqqJ6v2nkwPBuLuWDq11Smr9iHvD+Ey4M4MqBQSq3sZ73Vs1IFBm/iooRUgI5KzC
BiyalHgMjEgDbZr6BDx1r9KEQLPbCZzc0Fiu8HapWfjaJVUCexvoZXX+gMqjq6xd
wMh0aVgYwnwqm7hxtie/eab5gjRKkHjNAxUprM6N5DX3+TVjJcE8ljntA9eeNkw4
m7Xzjxk3skCrdFxlIoPaiWOdRrx+WtyZ0PD6yxhhL+yLy4QE+v0tGuh97+XOmQmb
eDXhCLJnrnXD1YoX8dM4uk1xwVdlOWBErsO19oORGPMbAUY1JdwXs6WsFnVQoGTV
Fw/d+G7TChbb8wQHzDtm+GgSYkROCEW5A+AWu5cCYScbFLWui9qzU2lhQxKX42de
T8ipLh7Rs5OK39E0PgmRkq8TOpHD3ML0C5FIJ99hmDyg4pMT7olmAMyBTLdnOjdk
MwQvNrzKKSu/Wpvl1Fwq/Ndxkas9zri3DENNQcVE3cEI4GMlC7CgRA5Mzk7ytkBf
jF0bCzp5iCyboriwoknBD4XG4wUtBquXUIOqDnt9cgVWof/vxWhVpzbCiWonLc7a
br1f+LTiecGds8V0GsN6v4zNGUoJRqTvTjWmsT/tbFtj9I88GP37tjDNEURPENEq
7jYv8UHD0J9Q77trkeNUaFKPu0kYuI5Si66M7/Y/xmAVXVdd99QjQJ5ZvHzBnX1g
zvF+6YPQAn3vLITYn9cXe5SysHQ3Zrwk3E/b5s5BKG7QCmCz3kIXgvjLeH7oYRA+
5LST0Gk6YOk5g2ckKGU8GO3nz7N7KJSfeXOItuwoLed7ylMk3rbnm1cyp7LiBbwN
cx77smFWuRG+xYSjvoQfbPsURGvGqlXko804P4z/T9oVY95Cycd0VfnmzuOhn+OY
pR8ZOZk8vCvMk3oNyI/z/b6PLr4ML5YYEchUqcCSVr6HtronTZ39LlGTKNDsm8TW
+A/6ttgWITrWO063MiV3Jhxu3vcY7NyCjLWUAOlc1rFuL1jpMYqNmDHWxsrZ8fFc
xX2QKP9kL6CtIV7qj84aWaaWwr074Px1JblRmQsOgXH5Gc4q4DT2GaH5GkDPWX92
hnZbp/GGsB3yBXUAG61wJY0OvV8JdwSr+mF/vYAdhSqrDRv43b75ohamYbd2G0w6
/o+FwFBx1l8aSc/VoP4UE8PpGEVZ0rcf1KfFdAAn+EoW8I2USXTUXmpE6SrjC7+P
w9hBJbhLm5NpNT4y4L1wQv4ZJoUWJyfBqd21Cc+9tdgienoM1G5MbBRbHYpvLooL
g6ivoe3PRQOErkvLhro/BeesxSvK2qgtJNr/0g6+anHg/c/36xImKhtpkm5I/9Oj
J9e7Y8129bMAZF1QJ3Idl+dW7NtV6FSdb3OIc7UYeDhGZpPJY+hMv8s5E6ZB8ZHS
Wc9E8maTbRNHXQaauPQZCvJuRpEr7H3pH53vokP6kw/rghONqiz7uJhErsRqbPhG
/9otIKL30upfO6EjXGTCDyA1GckwdcyDWiuqSvYetQGuT/MvlJ87rj3G0d05aaTg
Mbdkn0dt4sVHHpP8naO6e5a/yfSiEhdqu0RM3qRVdvZ7NA7IvaE+GUH7qHMg+L0P
PXuJTx0ycxJ095X0gXsO3XY3F3GGFxQqGCaz6Zvj5rOCFu5s2pZK0Q2fAv64dS0F
/oa6Wj1AZKUomECeq/1B3MIlWdEuvbGSsGIwOPuogi2R/DYp4R9C8cM8JMaL3kFY
v6uirdBgy17DkteQq+Ss9eUNXc37G0+UnUx0qZGsbBArje1EjzjNMc07DL+N3v7B
jCFk4hZGKplh+IOE+481kFuue1A/F/VuU2GpAw0R1KCO42yHwwUExeIMZ+PYRFb+
83O1wumQKlLHFiLjpXlSpCPJ5NplF82Vonp68JqR5zt1WiAuVkVtHYJouh36Lz6P
AXcAdf44DdupcohY9U4wESjaqRsUVK5AIAIH81p5wEXk+yjYb6eBjikwe2uxjAzp
vkiReFjZSrch4PO8zlYael/fM128JBzWIRjQ8I6k2DBmO98TpSoyS4T4+fyUGQMg
UyHGQ7+F3G685mdnhsKpPEVpWDWl3j0GFfGRDAcMdIgelIj6NAhpldgsjMVc19Id
iTskcBWnts91AC6hYzeqWX93v6KfZHBDWsMSpMQV2PX6xJjbb30ISwvSA1570/J5
BfIiGXl6erTDrFPHz/8XsyFWC92An1ETXHTJqTS025rIxoZb6W1yVV6Tzl5ELGmf
iyWd9IGNEhIQ8D2UGWzXeEJrwpKxYwm58xSg5QDl00h7NyU/Bm8IAYgoaUt1EIy3
q1jHnYnajm2zJwsyUoKa9yEhsAz/b59AT8Y7LpM5bUcYYIaHpaykCmwNf8+Pf1zI
db8xA/ZWqWv2zIOoBzp/dzkRvKkcnb3nzi7OU/Srv+jWmBQWYw+t8UrzZyFPdmUi
4FPhfT3Q1rZUZmsFYcK/RktZvFIDjsZTeCaojp73plf71HIIGr/4W1fGHUEYFYZ5
ptHiRd9bm+b6TIqaxBVbF+XOlgkUrlQWkfDUyUvwevVyi09Ksb2YVRCy2/5nASFe
Jp+n4ut2I99HzxCX8SCUcF7R/m8N3qgU6k4LKq2NFMS97k4MgYF76xHSWxcGfIHv
K09ZxhCeUtMQq35VRKrijS/VBPFx4iY6msmY628L9qqwZMjMghqE2LvEOgk+zY2M
C0mgjGJ8GsNCFTevqQGUgxuG/1NCVXqFuvx0aUuUANWCMm1LprqaDimvaBPHpDRe
yjAfYhh/5uVEJZFZJ3zFzO9jwRxDnPLvSklBOHpEiQEObIgfxTCnwv5SrTLP38jv
tQAQzHSXBi6RJKGDCrFb6YzZfOi15npxC2BoxnoN/G4aOxTyWSq9u7sYkhNSUzDl
BxWHzeV9GDspGCGuQEHnE/VvlZUG9XNN9YYGFT0ZFX2WR266CxiMnfzIczi7cq/Q
CQ7hdioi5BkhBtzfOA1RP447bKD0xR+qRKAK7Nx+AjtXZ11eOX3j9Qjl49X2DdWY
qbXi++JYBnc7h61Z0qZNUpG9v2FuYPbNBXBMog32kvrhP6ZS2N6u5vgfPymdN28J
9MR37YE1irTf+Y2jbj4/sbBSkZy5GeKjaXq2tMB0ont7NtDgtsJTzS/pr/gS3qJC
cFTKrkvh5T927yaW4EkF6KTVEPWby15Q/nnYXYU62Kw8XhpgO+ol1nJ3VWveN1MF
zWfX6OHCocoMTeE9gibosEhSD4VGKe5Yf+Ip6LP1D5cfSNKf4Ca3wRkwFv8FDVaq
wFcdjPvvneyEnBPef5lVhgk2L1hqComVxQd65IVgEke5bME/B6UK2v3phqCSwlm4
bBUEY6VyNcNNajU/Ud0y96OhXMMNfk22og8P6Nhfn7giPrUF8muzN0kQq6uYk7Dt
rFLUeJ5YP0lrnkKPzMlpCTQnffQZ4BgXI/XR2/djoyHjdWEu/ubms9KYFQ6XZE75
xgeZlL0oVeitka1FvreepBRJqq2mln8VO1XUNwNUrB853r8DLgJjIrNTH+a25x3P
KUOTOO/s0Icrnqh7K8W1LdpkXomibqS070hsDgP1qCrH1iHeqMmU+Eprb1nnpol4
bB23/JwUTaKw4r1ghT27wFsB4tvfDkcjbkW9lAXhf3vcuB9Rx29QLSyxMu5NbkQT
6HVH1dAwoMc2HsPnn4JyMwW/AwxqsC5/fiQuV54UcB2j6uCiBTd0FQeoVviwPDL8
fN7NDK/egqArLDeSNYWDofAmmbaUUm5z4DkcVQqkwPfbCqFmikT+9fs8zbPvf8h1
R0lFX9jghZTavr5rs+IKtdjURYGSSMxg9ZHxGa7FBhv+XdDRWSRp+F+d72Q06gIf
mKioblYXHsmgvJ9O9+ZMAjPC1iZYvuvoLTVvBwPXdSldPP1xMIUY8Btnh3mri3qv
KZwthEIlOU6pyAyvJcfchwdZXFRuHfreL1iA24q4xlr0DGLuhIUPAnynnQjmpI3M
rQ6G4BJ2jBAwEpyQ+UW1/4YACfi0UEAvQWMn6ozILkOtOPa8Qz/eGLXAEl/wDXYy
VGrHc3hd2HvlBkcSy2XSLxa2EhiMUKZEuX5NObj32GmnoXlVOPPqUomj1eoehdWj
QHF57PPrY4LtAQq1bODbeYFqLfJrs8Gv78SFHaQ4+zKNGe6ZkpaAnsOEQrM/eLdN
g5bqfZbu0I6Icj1kIxfHG5F77j2G8GetehTjTlH445ED0WSv8TfZ918o/cp2RneF
q95CoGD/8oyA+suT1KWJi5V/LqQSg01xU5WHi+w3+xd3SiY4hwj0tGo89ywrzd1L
V+xe6Jxuo3M2UICMkHM9WMSO1K05zah11lpe1r9ViCxy/P81Ent3Bfb5GrnNgxUK
ZRadphjaf8ZSnwhJaSdYZCKFpABepRtUJwjkH182QCtI+SGjbJzmR8AvA3g6SQHu
6sgSxZa4WhzFi2pIQMWfLShk2XvYztiD9yLTx51nK5OyAfsXhzaTOuQA7biZvFkN
ksxfjL9Nb54V/3xALL22sP4Gd4hBq4JW9Za3anuF2qbbQSazg3pfrhCidr32RLRv
L0eQdj3C5xMNHmrh8+Ck8QvMN8O+LvoMme51FSD9F04jyB7myPZ+3WOIomTM+a69
XxgOCfMd22mCgn63LPnO3z14dZIOLy4yJbyfh4uexDGy2RdUaDNi7qssS+3EFA5Z
k7Kr2vvRobZ6hqTS9h5obdYC+o9RDyBtvXGnLtqFutWP57cjOT4NPrh5fynByJ7f
GdLVMiNRnzrlA+71jH3RkTI4B10xjX7VoFcc+MW/PmpEBYNZCEDwTbQgKNUB3+Zc
ftZSvx/9hFj47kBipSeHMNxqIV1llCvY6M1K5vK88ZEl8bI/xhQB23Qs5elHKNzp
SyE1SI79U9seHc/qsi4/TUdt3dPSVT+JMdl1+Scjt5qeLmqdSnwEz1yU7ujAYeeO
AanxqkUaRJmmv5aH2WSYkKPHtduMCYnmF2l622hsw354Ds8C5HMNOuSS/0JX6Iq8
qVBHcuSZvX7Q7M1Npm/J4jZDPyJQ81IUDQJz8xOt6MUcvNtQ1ojyLCg7F/nOJIQY
JdY4dsSs80baV9QTlQ5XYQAajbudtm5Tqtz7+5wddZYK+YIMSE+71Fngd7HaMepF
rPl/Irj5RqNODUIrnzdmHWgHIVqa9sENPBdQf7r41UyoNY29ZY0UjYDkHE2iDTLA
cSb61mAUIe3BNxVEyPYq9rXgn/Bo7gR9u7j/hcQC/n8O8B+ci1PCUpcPRxYXcvvo
qiu/HjZDHXky7VfGYTi+06zJfq0mtzcFlMi+49NJCVL2hFG1j9mvi7fQJ2sMbGhA
JmaW8xt3t7YlRwV4Tt/uyJYaIb603trW63fQE1qMFouNaVP+g1lw/Xxb36h49IZO
BtuTkNDJIYC6GBVw7Ste81ptyEvaNwPMBj5X9h/HaHTTrH1RqNmygKVHY29MxNQ/
DgWG1+S7P1JGrbKRs7SxyILUQc5cm+XNZ+uRyFY9jKtH0qtfIE2KMmJy51NnoIiX
juO5bh26fhAQ6a9monSyGuPufapK/EnJoKl7YL3cs6Nd3NH3L6mNfX6QPgp5XIiS
9Cpb9UJB5L5u9yc63VGooIKlnIi+o201aFCS4XluAlcuPDWePu3G/yEFhLc2aw5N
pWtFXW3ZGDc93URbv168RBNoZQ/NC+U2WSaWjInS2kXUWAx0EEyFBa33bxkFBcLT
bxm50k0ZkWmbDPnfhf1uji0/K2/YUmI3gsLISrdK4gTg2RDLmXis4Kg7hWMt5wFD
SwtNSaWqwUN5QtU5hwXG3AFulf04+/np8dFjtPiaEq7w3WGbPi7wzBeJVmAbuFxw
dQjKj0YyGdHHbzIhX66nMSlTrBDuTrd5WPkh/U+AqyQdd7C8XwzKT3yR63cRg7tb
/ks7NTNVJx3AnBn1G+dnOaT/f/cUKuy4WT/D9NK+3goRjmlxpyamDRf7fDCRNKaM
q98Gv1Hvy/Vb7MScer5jEvKron1N0m9cC2FQeEQz8heVj0zEcbxIMEEME4JOeUNA
Eh43sBEEW+LTRrYI6WoKyhhHNJmo4BXLxzhO8TP1Jf59tEyylSHP5ccn43IZJRqU
w+eeeH++QaESr3MARb48sKSm2dwfob1bhu6lcghww37Grxx/QGLoVsKbqoT2USLB
UzhOrSjb52KMaXkGK8u344s+O+SMaY+hM+7UtBz5U0O21JWS1CKUtgVO6xzFZL4t
jnO3K02UKfUA44LWoqVLSunoDaMzxvy0t/18X3VQ7sJYaWVrAFUM4T005yp+5qzE
bc6K+fBKa+gtiE6cHqw7GLSuNcs2GVleBQq9aWuoycfYfzMGa6WsYlgNhE9yliZQ
EZaX7YRz19UwrJQGy03vtLDcypPlGXtTdgAoJwS7ZGLX9s+x/2ZATud7OQlebwEN
p5bV7lbOfCZ7/DOroavIzepsPIhbP4u0cMMIhOoMn0cCNeQM2g+M1GnGsCUbt78F
2RU7OP2+PnEktBLBt6ekD6htZX686sjwoB2DbMp6HvUDniACC4A9WTQlDVcLDkAS
vI9/3SAoEDkykw5/VfNYdgEp1ZLO+87iXHEv8qyDc84ULrLsshfLPOWdIaI1Hck3
r410KmyLEoUC2dhJ8sDeGPXJuzaQjgzErsb4DRfkL3BT3eSOaNNlXYkRTSqJ6MPq
OLlqIETcy0soGX9e9Z01rfXHk5yFg2TzEvlNqBf4O0gbLVEECWHWb4zdDlII/ImZ
h271lYCPnRJElz5CFS5ew8i7STAaHFl1cGUh1HVZ2PT23uxjPSmRJnZvSY6IyM9g
hp3s3YpLj/M3EbM9wE9YZ98ecGCDTopWYPAJ4Hr+Kx//xORWEzBx2hRUbXS7HIwz
ZsYgmobH6JAOMBuNnpIokn1smqtIYYg+wj6Xj6w3ioxcGY70OmD0YGPQFkoYfXxd
RRh67P1WGJoP3zDj+OsIYxOQQ8iX98S7RCoMKlgHGWIMU1O8Jlrl1u9HtNi4wQ7m
ji3FUGr+w7kc9Ad1CIVQzaChW5hkpOXtmcn2jlLFwNvfd7t0sxTbz0Zp/PsbwwXm
IBriV2rKJGfx08oG0xLECTkpkA1cxFDjiqBowfZmY6CvKdNovvzFGQHJPK5TfBo8
PWPQV0p//phLt/ZKxJCVVi/dOx20upFb2TjnpxtifBG8AjCL9bVwPPU3xScijbz+
BuhOZP2LsyqZMyFJcaK5FyHz3agzuvqZsaY8clbo0SkhoALc0/Mmr38a5UkeRzN0
BQhVonVJji0UoWoOfBEpWUQlNtC2NpIYLuSxrW7qOFlo7qIjwjaawM8EarSsKq2q
U6HKrSlGDuYJaKwaWlLHQ8wWsXDaJU5mFPiKhbDO/0wpbUOxCmASQVcdRk2OxmEd
r5BeDyaU7PMTZJCbrbKrlKfbw6P53uPj9RvKWjYZ1WUIcMpxMYUncwIHNSIgOscz
Eem5i9gHPh4yt5dg6wCJ/kzxipyWietYH6OuRk8Q61OoVVJIzAwFvqq0NHUjAJmG
pxzMtNdkPvAFrnTMk9V/ijJCYlqNzaWy6lL/48uU9Ld0ce+uMt/15s9M+FTCB/nh
PpPOXQ7jjauh2YJVMeGdVHa7DbkaPZcmlHlQBNLiN9ABXqiZI4NH+iWR78TdBPgg
gZMXAqmWgdB/4juog637SFKJXx0z7ahdvdGMGnu5o2vOdT3yJ4iDx2qlZH30TeUP
DVEQGaYb4GXMpMZo/gSRepbL+fw66okQ6B43+nNShE5bVfemWIeeeQ8lRaicdC7q
7MB512Zesagf1jV2nXfzcYGqUt8CY6+SHqgVcqT8Nv251vFMFaoy6e0DImy3Ple2
Z9VOCekywk17mXge4d3hUuYRFiqHE4NfjhkQMB5eK5GUAecGV6DBVWxvqrkSvkap
uQ8Iax3OPulyR8UuTGDnEfliHIJWvp7pGXvzavhrCD2J8kt6L52P10LbwBPLqyHI
NCiwYE19kZKgJzGbzgoVmmdcGcB1LaQ3RDFCByJrOeZY3E7jJEPKcWrbYiY/BgjI
AKrVdJIzNwL6geBUh/dYsFUKvXaBLYzz1hnJuAtKEk/HfYtMwgAzyD8iQ2LxpPXv
rjtRUVxYDGaCB19gnORX2FfnbeW2ndIotp60pVrEX9hps4rB0N/YB7uonVfrQKa3
3s/lpBULzsD+zO0kto/VSetscbJxVVpS2E9OlIIQ2VzqlS5o2uVnb9DDbkQVXsB8
q/Iw3n59G6az3A4NYNErCrreW6XSDRy78UDOf5tFIluW5JduIEfDayzMprEjFXRS
Idt4ZOk9wDJ4lQqO0moCL6lwTrAcRgJex3BYPyqoPzJhI6qp1epH0/YIgAld3iNH
+uBsMdXNd97BvqKkUqph0+yQXjFYYgDdaZyUbZC4bz0LguSnss2s2SLh3P/1DGnt
Xm1Yj7r4eORi0XYrv4+Jw2rr+ThlC2E5Gcox5rh+dQc+XkwpDiU9sz91Bqnthfcp
tRmjjASrTRjBFCcsopZKJDDi0kJnRaC0LF30jWOi2cXbtKBz21u/o8HeCsT00tAG
12K3hNUd5TTHUhxFEF2KiOYhp793P8dhsJ2Fv9l5hmRjvokX+kXVXaHPPIDwMeaq
i9TnWkc479MC4H2NEVlsFHSAaE4fSmnidOASQa6V0JWQDpN6zEsVVTAHZRtG6R8l
egEbNffeilCm+Ek99LO5mzAyKSQXMLuYRFxQfjOIKvUGs2l+AspGSROIm6DMJFxr
a+qQIElo41cFtPwn85iSNI4REECLTHdq7eB424T5bSaWONhn5tmiuAjwea9hHfjC
RS87hGBYuwIsmGkXHYXfvIUPIGcinPrHelnuKP+c+7chyKl+Cp7yEL/WtNiL/O3X
xAmJExc51T8RLOzWyOoTYB9NiRhrhl9VMJ/ckd6kktpsG5QJ0lDQ5pPXe9M4dauC
LN5V8ENd36a0gjxbVU0XdLfzOeVEBDa7kjn1yzoi2iYpf/mRmJcokAniWXLhxwIX
ltZhRfLy9UwAAURgbGNTqVbRJy4Z8Kcv5InUz5J7SMhw7Auh/sAFSB4bgXPa7s1m
J/rpUs2xV6UobKRctsbaHXf2ccTccPyqlnVbjQq23Oz4OVyrk4g03PpTWUgdx4EG
Ra6dfPaE03Ga3jBeXnJO2F+9z5EH/mG14wak13tjE+HSJAOr1epwFw0vnJdSgDJd
w3U9xgJp2YklKNz/RyTgOxiXq+RGpeqhyyqN0L3+rHkhOZEi4mX1alm4ENMHrPjZ
enAThmP36IUhBLUfIZs9n/G5gff1GAAgJEF6FQ2fVsmqWph61JhQc8p/pedAd4ZU
IClbJOjtk35AOxddRVVYpt6pBlEeUTa3A9Um1EoehF3sybEzYYvlYAbAyhLcYlLg
/z6Qs9S9Avjxie/f2BUKb0bN0XfwMlJ6Evlx0F5w2I0P5rnte/7ET/3pKOyZsmBf
+ZLkSjQCnOGopdftfU1wF+J7PA8j6SQxzxQy1moAu+NkjXKPjsBhwVFkXdkit1XF
bkOOoiJR1D9puDkB1/iZiGJF0dQ5kzrKGzXl2JBo2e8ZE62EInJRYQ57NWwr/3Ve
rn1RL2zy7M4ISWLGFTD9xBf2RBQ8fmKD538xfG3cg6/nhViw76CqqmLIGKSX/7yw
8PuDf8m5lWoQmyE4mh4/g2h5rf9fu5J1BG9MlmCOxIx02fys/BKGY4UgTYdDcT1v
cpNq3PiJN1kgjdb2VTE6r8dVpgWzRS1OUNOAglOjxo8t3828HZQbuW2Fx19CuRyy
cQDbxPiCRyI5uV6CvyHeEPQu0JBxp8XBMrPs9H1UpNygTp99ckpy5JC2AcsV4OLg
1inYMFeUwFUO74yGXoPN5V9Sd+yioR6GLxRA5qXJPZpMSLAMS63F1/c05aktzEJU
9aQVJvvPNCBdyRLGUamek8EBmz5V1EeyQer/jIPcOrHTPuJ3CPo5EZ7LHKHAvek0
vcWVLpS8OGW5n9T5vqHzfHvWeEVewNw8bGhbkwAis5N/WQrYsx/lEhv/gLllt6J4
GDOOV2EPCCN/bJOvszabVKT6Y2ncH8plqjNpElLDbb4qHtB2mkxyNqidL+LZzUcr
pj8Rks0DD/XofUfc2zy/wxShcx2jYnvMLC+xN2EUOnRqpYmng05ryUFtFAwPqlwr
dUFf/CSSzRyobH1VzbMOdby9/MguNYGC6Biqml0IWPeaK5mVP/kY/NArmUsT4Ztc
BStXOMoFRPtUjzZkMMD/1Zz7/3gKblE3hBQJHQ/x5YvFBLEV2m1gOfnp3jLjR6K3
yVwPpvcnc6WSpxGWCEcZgQjDTJgYLl/zb4+NLMmLTJpOHDBhhjbuy1OGgePbtbqm
p5hKLGBolIveQeffbLre95Rjwe2gW0Pe0dNxrRZhBeM9Etf/CjyABrK/IwZAXzy+
cWrb7cBmLRQsApQzbPAYyBhc1JsgeHWGxImI2Z6pN7D5Fx9CWFYJZmxStR9Na6IN
MuyyInKqZqIfKtBFOI/sXLpNj1955AUqNeCQUuFJB46g3wKT/ENjRceI282dSY0r
GhzHzt6Iz9p+3Zn7MzxACUJhy+QY5C5KNslrPXVzQohmXo1DEY8LmtCbugUuchO1
g5/u4vaQh+VB+vToUD3toxDRM0kNOFTtb0Q1+6vziBMk96bCFxwb9QVzuN2rvWEs
7BvvdaFZlJQrxP19BA1ZZslKLqE7aeN6XZB8Gdx0mQd87Ttx/SEI5fvwLCr/SLNy
aMYVJo5Eqbv/toSjG0lqvU9lWxtX/RH12nhUA79CPGJsT9hCwn+oXPnwXnEuSFMl
1Ac9QlJ8MeikDaPr5/2f9E46fU1YnY97q+863QE8LY4JzznuIfWWglG3fd54d5vo
7AbpLaLiJ0qbOdUY4ubPEoQnBK9PNq8iVqU3vjUKgEE34AldRQatkRp3yL4JWHMa
iF8pRNEVe+asz7X4xE8votAJ33Zc7uqT4oVFfuemixhBeq+gWBGVlevVn4jzU206
ZVgmw6zPFYr904ev9ugcpD4qvPa1Ti9/pqQ9yk1JZI+g0iLWcNy9dtM7UMmedBLJ
Y7na+XT6EoHrg+2tk6w/q8zfZ8VDrCXMh1emC8jE37xfLUN/KbJYdyoC3cM2JF6b
GgCf52oyIMURUBmWM3GgZeUBIJqUgsEClEb4XW45nIl1CnN6Us4pJi1hB0ki4inK
HLwURXDgP5CfgC9eroW3zvg4zHs6U4OwzDFcOqNowRbPkwwZvVkoqNqVtw73BWlg
j6xveraM32l+H6hxk9AAfb1csZ7O4bkl9Irvzwt0uD7iOKm3uDkxdff+mMVpzngl
QcC7RNa6lDsvzuBxgVU01ztkPObETqCLcUAwAZUnnLtyDfdpTdVlU/4fwBG5c4x/
mci2DeC5wV9SksJf7vwuh+LkLTyxLviw7qtLn3VvjyX1Hwyjfw5lo8neT7a21t0K
1km9t/jiOEIkW++xFqxXPYWEjpKYbtmwUEy+SLTzSHeQvbIO0wRp/cr4wWVqf1Mt
+RDKCu1j/ec4/98s9x/vR2AzJSl4sPnupOZ0esLceRBqZQ8erev/rrE5UbAFgKNI
HJA/Jpfo3J5lqDdGbj7YsXARgYsTNV+0bWJ4eLxO29KciTMk1ypmeslkc2JPa4qq
AnLR9MXZmnPjYv+Q8xt61oYjDpWcpFdo2bJlQXBiJrcQv7T0KP2TCB6xsQCKew3B
BssiOwEn/he3EBrpwnDJYbvkKYX/ogooA7v3VlP8gLU7BVt/q/OCnp9+sho4xsiL
fAUuFitNc1hPao1vlaRN2k39xA/O2+6D20osi/DDEhHAHPyHvW6cxCJVNG6u+4rG
zxzuLlh6pL5+y4Nk4LeWqGdMA7vzH8Bodo5YC1xueNa6flHaVpc7h4AlmplW8RRi
YvFlirwjte1QtsnJaMDyLUBzuJVpoiyaufgiTyOPy2b5rqxe1lJi+k92XR0uC8Nm
wbrpjEzHhyZEqpaBoulsxXHu0he1F/GXS+qc1jNouyUvsjAaHGRWawBjbx1u0My2
0FCVDzvzUNT39cJk4Q54xBUIHj4QsH/mVT6zsq2WmG1RYwZQcqjDVzVzIHekgEUP
2OnxFBb1sOVMl8i5glB/I8ZxqkBijkEgELvFuKLvRhy/Mu/m7Ay9IGIJuwXBn1sZ
lEbZ68NaPu126D3vm02cCBy+jXm2o86KLjo16de/WIotYhfb6dMUqKyHBqa85VIM
viTbI/Sp1CDui+dbNM7hJmpKsRHrRIzi9Iv+pLdUmVEk5Od2f0zSVsyBzIPKiJE0
bfiAw0D5Kd7Yx75uxYp/SJF+J71bJ9idNm9GrZOTeRJ+fq3lZFK2mFAibejXlg6M
A53lGLgvA8XKPsb6mKrBF6Tx3PUkAbK0dhixnLSE+PkkNZsIKohyezzRnGBgvfGW
OqytwRhX6ITkUSzlHuhc6DP1VxnZkj3W26gTDwRTvAduIz0sRlkqtpnDDbhVzM4E
mq6+xqf6j6z8K9m3Xk6qmniNZ83JVB24ZmsVRNSzA09zWmeVzRAgs8+sh5l792hN
I4GaAImwmksEb5WlHQKrAhDrbYgxCWKWKAxY4oSL/rya56b8CNUBXfOrWrHrIbh/
OTFG/ubAs43UAhX1G8jyCUC2dMCycPweVzgyoqEtqrQQodyLcVwUlaixL+9u70u8
OIJmBbaEWnpnKKC+maWByzfZbuBhbmYfUP6juSm4l93SqTWs9D6JC7QUIN43Mk9H
eexmnI75/40sou+NDo0P7nhWwJlLVnpN43oFNf30uG5GxEMKKJI12MV5fzprW9yF
blJMYWpLpDL8hbmfiDdR6v0RafUsoNOBcoFgms6Cw94b5X8a3hD3f8p7rvvntb3T
ijOOlfF90fua6iCzImb5gIeQCnTu8HypmU5WIEmlGXx0XxY0JSYqcnA+7VHkD9Lc
RIm0gNtyo5iGcy7Ed0o5CjBuDyOWGt3eidgmznNdqh+PMjjGH4YzqBWTmaTBjWa7
60iRkBWySbp5nhrrROOYc0LYZ1EA1Lj8hBYHx4Etl1bnQwnJlCqiJYPa93rxmsmw
JaASgyh7GyNGvjiMXea+7pqRfxwcUa7qYDdWriog9p1G7XgLQ6Pc8eq0ufBHn2FU
4nU7oc8abFOXD5Qy2smPvBgtAoxwLLOc2mXMwKcfDQpE8eaqmhaaKhJznVWZ+N9n
1zFRJS4oYhPabVnzAmy9hIbIO66cbOOF86Z3Bq6XbhA2cjwARVHd1QTG29t1f+7B
K4GEOivJtK3rVurvCmsSElpRs3pBQHCGFwqOMRsSY52MwufwLUs32sKmF9clEYQc
X5beQKdSoNScaVtF/Zj6Yk56ukhNERFXCcrhZHFt0mW0FgfnWS+P4cCuBL8ZS/cD
CNHdmaclkWjF/zamveUfl8wuFgXVXgWP0YWYfITRnU5cngmWjvnUWgherjaVDyD2
ZfiDrWm5CnO0eH0Lr7a2hWhpQqu3kw8Ys2nIoOpHRCr5PMzO340hfKRgpQ+4/4i7
jrDOhDiDX35t80bN/PfJ1JVtvsmqK9BpogbY4Qa5b+OmXtgZtjujI/HWS49HrJPD
7bDojY0PSyEs+JrGb3l1lwLk29x1rm9vMaQWzdKkvXxGRDJxvIahuspATRgTFIdA
JNC9lUDbVzYmCn1FYZiMimHsk6b+Gb55WkImdJnSDrkmp4mnVWhph2/ac5xmNUAy
EM84wG/8nD/D31/33anXWn0DZQhq91IInD5DLNYaAZaM5LUNedjmGQ1dswN1F0fi
DxZ1cZ1WHr1Nb3zet+1VKkUIQLqq3Hp/9i/z9mwj5dyRF+6A4E/0VbfH8jq9lCtn
MIehIwvgOWsfVkmfCtFdgdG9JeFVMoEMm0hyYXgOsePfzi33pzBIEB/XpExTblJG
rkDRBXGMjiiXbh5J7JG7Pz8BREAGA4/c04RbhYFpbu9fddEbcj5iwzHFKLeN5EpH
pdW4GzRuIMSrzDYz5yY7e4yQgYkRu35Tnhk7BLrXv9Tf8fww8E99spOTJG6N397T
24KpSFWfeBo2MyCTGIFt6/2k+WIQhvS4HSG34vhiaee/43Qf2w+J20hXG+9C/IiY
HTMKbJxSeivAfnoi8dbfiec2KNt/RW52NanQQf7KM1vUUm5ot9ZQeWiSNcCVIRy5
tLJaTgP7+ftXwwP4ADGOLjl9QGnX1Vv9jBrX+tdDVwH5cDMGltMdJWl5ScnUr/ue
Y5Ml0z/aoyFPLkEG9sGBpKBZoUkOd9xPy8SSidUW7vAhFEYN+Gpftxze8xbfBxyB
/VF41VoBGkF5EKrvmVtTJsUcRMVhELQD9MLmgt5g9rKjFlu6jaqDYtKDGUXiJgeF
A1ds5O6Y+v8Ivaez4xLGVeIhETTKSMbzJ/rSWJxigb09V3TwPByuuUYloOOeNPrZ
Z0R8GgHTxDN8l3w5xn91GaT9Ut5aOmzsiY54ounUdElkOBlSRWMcafXp1XENoNYj
f6FVt5881XqzHlQcIC/c5gZdjBkipnnzr+nnkwxEHVaTkEcH8Zqk5cKHGsnP1equ
3XXopb//3xmekxB7OTdcLCzvnfgyy452cY3BUWn9d2UmCV+fw7AcuBGu05yJamha
4V6PkxZXWuZc2zzMJ96M0OqjVkXyKl3Q98G4Xl5Y8gkMiuTinnTMbncdhbry4mrU
GaJMoHOjDsP7sPEtkBy5g2LDjud4Dx3dL76CGoYhAtU1Bl5xmuJxUVkxtfSWln7Y
fhs2mouR1egHWQ8FSABG84PdGNCIGd6glS7+HDsV49QqvgMtpdI4zmW4sTCA8/7k
qOMXGkWALQ2ETPMfs8q6NpVznEZomusRfqPconCxQ9hfd1cj/gitNSDH0zl7/09r
xHlhVmxYeI3NFcafiS0tBom8bBfncuIARZaKP5EpmPHTzAXe1uJaBbuOPPDnjcGK
0qgDyEHm8WBgv0fBqasVNfhqmdeF6mx+jPToQ1O/jhcuAMUfW4/k6BmYONcnkJVJ
LEvygtd/iloCdSmb0kmiAjyJObIqJhb1Oa2w3OBjG9e8849bAiTgAv1M0Ltgn7MO
GuzY/gMB5Y3DtOlXPb9vmyAUmOMT1Y3mST+BCeT/CguM8mkpH9cxeTmeMEUiZPFW
8VXRcT3J6TDNATs9v9M9n9ZNFzyV9mRibgyYDYVLWFYMjdD7wrvn2zqI5Rz5ZIwP
b4aQzqqPV2+HJvu+q7OHXJahf78eLgm4JTqs3iM2kO6hvIczzFf3eoYHn9dWur2+
V9nGT1FBsnQPD1W/IKo9ZWIE1bOM+MrfdPHu7+QQgrZIDrBhVZiKRoycBhVCh1PK
GF2LNcz2HKelBANUfIbdwrOVRKISkVUj9m42JXdsjjsDPYzsE5F69VzF5H4QQfzW
TMRyFb6JtJnZ7JBNQG4oGTTj4+bnzNSPfKCzo+DLkygJValqkVhNEJ1PI32Ts94q
eb+1e5+zAJujZTe4fGDcg3f9OQwVoX3UzJ11aKcxihq8F06qcsk8N3QDJmfwBkkS
+HQjVK/y7kPG9HdcItUm0XTCW3UqRJ93Yq92Nh1UQv+jbC61s9PuVHxZByaksn8c
sz7KLZT4gadAnQih26NHIaXl7mnTzn+Ya3r2v7soink1OpAZQ5jI6/I+H/y8qSCs
scrOE8RxkeWirS+c7x6s4M+M4cEiuHHKNIcRl1COOySkO9XJej8KuJtuJxfKd4d3
DbkZT46dd82aWHIY8GhiZu5ouLN0ftzZKaQLd0ekDmhFnzUlsZBOgoi2u9Ns4IB4
QDeMHYe24R2Jd7WtotCGrELtQlQjkvljqh0ur9caWVSo1+MYFYBTxVs5OPvuaoIP
DNj1VeU0leuW0Vm6FVPg65OIUrgzUlMVjkLXcDLnxptukTPdxU92fsME/VQQJUyd
LfUY54/X0yaN3jw0Qi6JdBR0c2S4pM5LX2VGpIMJGgWXWnL9Z2gl2j2IJ1fvl1pd
PkbqHMuMTn47BHCdxhrITEjZ17/aeX5i94MC020gFCebnedox9hxbwQYILkFmf0H
1fvFtcN1mNCOPWnwSyL2XYa0TOUtGTVSJ4U/u9Krm9ZcHH2EKI5fTTa2vM9qpuza
hHBGCThtk89eScpoVPzZFzvnCo30DXIYiMqweVjNGbgBbMyYeYHDlAPy/TmGMbPn
prxT6n2q85QdVNQmCt48uof2v+7dZfrh9NjH8zzW4e0VwXehRhtFhjSDGBnam3gV
3uZbsOL4+RFbXKAXu82q/Q/HDphgMnF7tYcmTHl2wiaxNyskkfJj1UGO6YEm9E9d
oKz3qNeM7yWm1uhhoz7hx+NIafAY3DHGb0DOY5gt9WHSk4JzZbEskMYvD0e+EcLr
hNdX5qE2EoHxPmy+ogfoYY3JTgkPxXvN+BG2e1lXwD0k2YXUzqqM7+Asnp8+mBI2
cmj1FxW+YWCm8cf2Ltzkn/0GMrv2zQiLd7mMo/GqXz39RVRLkrelv/y4pY2dJFSk
A8qasROj3cQWix9rTCpEnTVPLzVi8awD8POmr3/AvVxz71NDQ+/ifGqbEwqqeRv1
/b2JQvnbRLjUNgKcmruTP7O9fyhlK4nZk+py44H4kZRvuUvPF/LM3TjRNFI99vHX
4+KN/fm7fdbl0fDPRL6GYRjWm0fCt/Mtsw5bj6OB4RP7sphuO/AmV2IclMwTnWIK
G3j1JCk13sjYJ17Jriu3Z9ubAW/cHezD9nxa+nSiwWa4Xoi5zYEEbJmf6s3enkyA
bILhUJdxXjQDlGnILG2kBx9Y21ffgw5u2tyPV46Btlwk+4rW3QmxIrgM4jBU6JTE
FM5c2jGfMgcxZmjK43BIybEbYKahySiKt7QxgrJtvS3r7WwwFUzSiJLz9oUTXaOC
j04WUUAMuXJq+XTKd0aRfeXyQPqurL2QKGWWkgi2WERElUXYn4k31kHzBWZbHULE
W1hKNMalnLVNGPaayz2l+T8U6Ql/GfFg8TjIffxeZUQi1CsyinRtSLcAmXJ6oIwN
mUiJ9ULOl8NvEMJrtquBpNIOPZ/U+2cx04XLQ1RNnBYSg+Exyk5JQyvYea1qiqsf
h2HWpakdHAOYH+vQiTe64p+8hcpm6TzhrTsauM2ZOXeV21iMOuK9WZYPDt/2wQdU
5S4OxvPz1Mg75eED8YC4o0TferhJSBvRhFvi9ImN0S69ZUM9eKLH4JXYaAnUMmo3
SzNQYdllBJbw+HoFzhqjqYiIGxSGQoqRhVE6bqBR4lGBHU0QS+ffzv5agvhB63cX
Wes/e6FfFfezHswG96tYAqg/+AHqlnhFEdKsDDy0DvCG+KgwVv9TbGLawEbHv4l9
ReHj8Gkdn/BuJNh+776OYyGe0jzyA0nHyAoCQVolzB9+Z9+toD5keUvP/wcklo8m
af7KLZ0FTNULAiAGOfUJBmhFBzblYlWAGSI1rA3VL1UBAcF2+LoC4UDf8f+2jAyK
lA+XYuFYErbKofWHcvYx79NRKVdgVNhSFnbvK66KKJR2m3DDNnW/QQ0EZOEYcDyu
TCjowhb3wEBjsVV+Aa7lP1PjcDrlAw87SJHSaYJNufoe0y2oxUvnZPLpziZNQ/2B
wAPetCA9zMA3bMTZ5gYziqMoX6CxSfhy/nu+0D0h2fcY2sPLnwV902z4KC/RLsAl
1PejKwzvLByqkAO1j6m73k06DdS5LzxqS4CHEUisGTqYIqnWqHQ9HmK9/TJoGY0T
tTkSBVPGVPCNtLpQuOtODL892hn5GuYI56e6x1755tvF2HM6kxU2c+p5ZsoHJO1R
JDAANu5K433zZzbv+oWM+km99pG0gakmUDDfX41hHPh4YX6neMffQGfqz6xFrOgi
fEmHAVR8WZZ1GAYM8UkKuO67fT+v77KsglDmPIKxHx5OwYRFroIk0RaIebZA/Amg
NmDY90hD8Vmm7GxcqkgZRRCL6SBQP1KZ/5VPhBoysfbqysgB1s5K7hCub6t38En5
RPvbJkrJgEku6p3dRwQWvBc1u6gs4H9+/2HoN46hSwmAuTy76eI9PfxL8ylxyhh3
22YmZTuU1PN3trVn+RXR/w0zdBBggoHYEgQTDY9TAPk7ZHiaVz+i1o+qWvliCMBH
lIQ9DgBiF6A8WzVP0ex5vbx/fvcD/DTUJIxVjbX+4vbBmFMrZZRrHo0Z2PQwVXvT
fxq6SlN2h5h9AOvP/mReyA1+H2LootN7IZZvXORgTOmp3DioOu96HWDy26j/oV2p
PQZTCFaApT6Q0ZUo4PsRaoheB7epzT7XILaCKYsewotNz47SI5zdnPs4yElnzzuR
NAeiSG1hSipV1wfJLFdbGpVMvp6h/vHZQs4XWIJVo1zJnLODDgYxvLq9XfEGXmcQ
tV/JkyUTkySsMwiVHeVbf1fGXbMWZZWdTz2tNVpBUUGC1klv4P6LYmMQrrqDCQW3
6EIQ0XK3GHpL8n6QnvwKmhHZOUyjKNknMCLK35+sycz4McJAib0NtRjrr25Ch3uU
79BPCTd6/3OmXzfApregg7Ux3ZH/qr4iT0ux0qr3uCRvG0Fv2TCMwbUVN1AZjkdH
kjwtQwzEEAKwKLAGJrxvbb0GIo9L4mOPyH1sbxVV0F/HMfGRKkKEmY7x6jyi+loW
uRIvzTbknz7Ugo0SIQ691L6a5JF/nI2cJs8eCDO0fpwh9Y0dTCnjrd9hNPyQW9pP
/iRE2owAO2ZFV9aXtXTaSduJq26MHC3XVndnyXBiqQk2HuPgfIjafLr5ciIiOfgO
0lcp7UAQvWPvXq2KGVOc8Sw+DJHwQOBEL0dtzj19ZKprF0fE/kJs/+CB7oDV2QYt
1diuJ8HOZ3p+6l69SbKY68S4b5WSPENSjhRt7I0DKD5roqoRsLkhVRC7Xvtde+Ai
gCFLXqyhm2vOMQnV9x/uNrmYGl031ZURwiuWusQ1RozURz2phE+VoHKIBjO00exd
RypXX4k2HQqGfkW5MkCGaOciQf3gbf0H1NhBQ65uAvJ8DGIVGPBKYzDsc88EtuOd
LhHPTnEJJqVpQbpdLAhLM85zXFTpof5F7L0U3zssvb72Jf2FqHOovAKmvcA5HDS9
DTQDSOx8CBKCKprQ93yiwylvzhvkaHcgjaeuh0xskI+YrAdcQWqEYoajmj+mAs5P
X5nHB+oIkG0wyTQSg20Y2qBbVH8DllxDZXj6oH/v1iK5KYrLh3S+u7+h13CFJq3y
r1FyVm1CvNeuUAKyv4BxD5A5e346Zascyyl0KMyT2dT2Kahhgc3Ubc59qy82zytl
c5bpw/zxLhFZseKSxcG18+VilxQ1k26K1C+sRENU/Ujm8lqchvyVmWowWr6t2Kp0
XBpFm8VAFnUs5CDx3/p981Vr8ogvLkHs+g9a59ynPSU05Yqx2T3mu03XmxHtwMMH
NY2l/eYMPY1yuuQFjV638fjvMjLO9993RQnXAgcOzKJtLvoPMfNcyNugvvRsJGJB
zXkzGJwNTSZJ0kn1TNf9lDgu+8DEejcu2JfVmQu8Phk0GfWlST+prZkJdTzwBu59
e+ZRMhqqswWh5VGCFcdSCK4DW0Dk3gUoTD3cpngclOxlnJFb4yNtZKbYWBnMPyri
/QeK+O6XUAAvHCQYcYdKhQ9iV0EyhCqLD+TRtZ+k3M8g0xyGeFzUnsLrQ20sL0UK
wmR97RruB45RGqwZUdqVVqP1EeAXOZsrty1CkY6opHkg7aPhC1geHXrVxWiVfCMh
lVceHoLoasYHR/Erx2p7KwsQNASwf24CxtlMEL47CS8BYGoKxpzpG5yOXNe7xfo6
7XYC1VTHtadIqCakb3BuJT+B/S2cJ0gQGjOSD+YWz0/v7LzhwM15nF8Cx104tBlA
bMZjX3hMN6i+6LE7dyHMoJ93WCUMm7OAPE/nvRSvrIuuvw/ez+k0Jexk+oH/DbHV
3oeu3gZUeLVkDcPz3Ws8FcomKitYK882fJeJMLWl+i+oQ8yKWnWYFOR1+2JyNvmm
yHIjgN+GTLSHQNtgrH7OpUHUFdo4taGP6rETLi7p0RSd/V1giWfaA88hZzRfvxqI
7iX6GpVQH/9QOaCgbbKIlUkeB3giz/gfJWq4jgYBtIdmB3dtRbp5s2BZMadKmQfi
WLhq4xGEXFZkuzgM0kuKq0e4YkdB3n7VY+aNcLuch4oAFOfhpVL8ApKSBlDcDaPr
hmy5UqqfduIU/rgSpKCdl9tqKlD1IlkooOulMElsK1Dg1CnVZYrJLxa2//s7iFIt
YaTBPCLMWfrO3RSGAZmBVp7uukYkB2LRf7vnzScKT10JBYTHQdrfx8boREeInRLW
QsRKWrMYFOuMprfE5lP+FgxFlNRW+ouQKFey/LSfeumkRPz8UjCAx6kXvIbZxrUv
8Mw8zcicY6tzue4tblsMIACp8p0k9fIC9zkuNFgldnrZkGF0J8eVhkiloVclE/te
k+UqBA/uXdczzM+xMawli8voiIACQV+H1jt6Mo5Ahj9/wCzqvrXeLfWmAGedUh3h
TUkfL8mFcoRvrXweAgzaPVnatNlpCbrpGr2DWQz922pOW0IJuLRDjKWQgC+IfcfX
HuLUoG+MxMNyjzpp+LUvYhtnYFWZPkck3u47vAQVILvCMzdu5W4nFeFmeNTChZh6
DCe9kHrAy9Jgi/qMqArWrAlzJUoCl2FP46hbwQNZbMHoViFkz0USPp63VeDhS4hs
UJZXUesRTzmszpA2AwS6FOyMApfLFrYeIOmFoDQBy+tFB9dGrL7tyYifDjQheKE5
cD6k9DCS/A2AuJlHCj2xj4spE5ppUl2ErsPtgS4UhnH1pZYSSh8Uy/vI1foswllh
5kzn9ARCyg3EMRvALcucvZkEDQw6CfA2sRUA5g4barSG89CrLn+VsohWY1yCF3dN
uE4i0+esQnNJznx0SKqJteBFaACu734ePGtyFZsNgFaRwHXgU/rhTvicaccnhfGC
ku4p9vITWrH1YSQbRNEqjXKVPz+5Bacsyge/nLTvxqbEIU9tTZrSmMr3El0LI7IY
BqZTwf77izgD6Ir9g+YiP7yPg/GcNtVBBIXGdWtK1RF5n00oqmHNNox5yypYCzgC
dizve6CunFb78FiZdniPu/KBpyMT0a75yDI8wQIH4QJ7FaLMyTIjgYtKcutAjoIB
XABzZGGjKT+piWzB86tTHgUudXSUiOI8aUb+Lur8FOEeYcZaoRLAU+2MucMmEXfr
Tb2IHaMrqi3wpxAcrGm1jlH5HPmM6Den5Di8sERfahYFHqLtikoyMS1G6Tq3G/2E
2L6SjGCXeYbS5+bvHCU9VQi3DMgdZbbx5tKv4rlLQdHq5wc5bokfSsyaYz3rR/V7
j3yFGFHxj0BsmY0w76sWTIFORBpdDGmykl62bCe/P4uTl3EdD3xO7H/lKNWajrTq
AroyTkLVnow24rBfEmm2zqj5K0eW2xv6E4EjrwV+7io73kpOMn5/mcPmOWrAaodD
h9oQrvIGyx+bY+PvdfkPa3GavDeajxOV1WQOea9XzFmUbBBcXmj2kHl15PibTI7H
k354szRZobx7r2L8zn1Exn2+maNqFHoLfm9QFdcRcWKRr54PHkTlKkg0/Z+2F+oW
jcjzMl+XKoLFREzeFTLWNpERkteD8UxqdhWN8W/Bt0dcJuZG79MdejmbCRRwrWHr
8ihQR008GOqtuRwaoGhMkd67gw2X9AwYXsMvRET9dwma3IAmbFCKE0K2gHBtSNWE
1418BSwI37dGYNZytPeHxBt2uXIgkdAI7XLlSIr7Af8dKAojpZyuwr9tD8OfXEdq
az9DGQdrFNglSJrwnWGOgUSl7hWeNzems87f5K+cvCt0MZ2arSDh1euetrKfZ2No
UFu23IfrGLaiZMaDkkHJwux0+hPcgQNvVz3HcCyQtkUOpR6671ROLer7Uw5wgoPl
gtmYguFIpQpWZ88cEqzxBs8uU6+i3Y5e0cWgZkHVzk2F5ebl4zA8Oys9oVumBfd7
rkHTYsERaQUdnqCuIJdTseluCf1RhBS4mT+Gy019rGAo4nKU8y/A+LZuP8DhJjnl
B5vBieCL1jS0w/0PIDBJD96YJUc0TfQRh7FSdo9k7WlTb5fJcQquZpOgYLBXOb/7
UqrYiy4G07ATV6yRDDLuh4TkQo2PvJol/06U3XjQf4AsuFRq/AaDvq2kUf0aHsOu
HHirYzf/ed0/Jtla93Pu4RvCY8JFdK94lY+SBoXKFiMkMztmdhCzArn1nCSQWW4i
PDDrBMfybjhAy/wKw/HyT5MJouVCOYy/zGVJJLjhgNteGReAwcBLmWjpqGSmNgMt
k3OUuc41DVTRJ36CTtrg9Tbi2l5MpuEVQnNIKXb05BwKkduaHIz3YOxwHrPlXaoW
t264jim01zQw8YV1R2wY40ITvSDoWCaTik/yG5InOqTL6zAXNC2nnllSyJDw2EWn
LqNnHCr9zxTv5YTg2m3zqz9/XyPXhO7b9dFzEzO7yxspQkjn+Q5d8hOmaI+2z9uX
eTRTxl/ogq0Ucw17JrFC+S+pEKos/GcbdFIneo4XJeSleqVWK2YLN4MMzdwOvJrc
Vl/yX961CIPCmQFwAa+iThROYfXbHoBgrXj0JFsiiM0oMepUeWTW0AXNbDaUQ2dK
pkC+mOIj1Cd6HYLozuSG2XennJRsp1ORZfKm+gqGiLsObNIt+fCAsLcV/ScDeU3h
rYYYCDyscXLViQWyGMXR9XGzIVirAmB3bHRG9nIrCdeYdXHzAG8KvL7GLHwE9hLV
2OhmnjUIRWGJAjb3R5fMrARYiH2OJ83CudCOS2O7fjCruVW7ZyNqVso4PQbPzjIZ
LpH4ENpYvw+Vn4DwDDNt5Wq1BK8tIAM7um3r58jvswTa9/h+CPAQUJ0quEKdOxmo
4aUI3wbH6v1rOLO55U+INDE3axAEp/idgxD2f+q9VlRviTa4SHsn3egTNJJdua1h
VED0yjwaI5t6H7rol7HSJma0lXN42vba+7wTb98IbSuBHX4j17EVO5v3zifI1WeT
O3jyBgeDffCIGq627jJ+0EuDsT/IexgYg7kLa3bWqpRc3ydwrhfifgaxA2g5l3wL
F85DNFREbHLMPnLvC5N7eLTiu1IxcGXLwEumAbBY+RSNLrlTBQLcg0853wXulSh+
u3dYDv1Z3HmG+WA6z1pkUo/v/MD0HvGbYK82NtwR/vgPQpH8Xj+9vtgHMAA/oGLG
/ISLF4NnBkmtz8CPuCKspZNIcvwtADeENs8SaG2DKwKNlgUsHI6Ic+/l/w9L0Kej
JjHu+L2DoQWiZLN6GnEIuIWOnC+mNtUkIsvHfPDF3fa2KhTSjfiNQLLWz6ONRReS
BeEaM2yKYupPSI+9jV4RgHJjezbFQ12kZ/FIVddZ4rFl5cPCNBcuj2rL+9ltp028
OG6I7+uuIaTeXFXtG+hwY2SFf6tRWVD3XQTkpUGcVEBIEIw3vbvh7CsyQOzp1Upq
Pny0qZt4k2+7Gk6EHLb2gtDH3xLQjiD+RHp5kgRapb/P2AOA7xMJl0GT7grl72/Q
KLyToqEwOKHZGCm8cN+vhv0naOKbmsEokl16p18uYX4PkrtXfR910xZZsqFhSs89
BRFhbExsa1WrSRy0f7zW7Wtyrv/jl53seZusC6dQlvxLwNplzqHxzohkfIDonT1z
BttM1QoIr+3fnFUVqmv8Ud0x/SsCWl/Uy3oSByYgCz9KaWoV3rgyp6VWEbDvv2/j
SESOWSp2QxvhyJOLdNdzQbklY7LZMOhNAzIe/nSu6emkka2bQ6ofhsj2KoqHOIAt
t9qEoyL/4kaOWWSmhEWYG6dRKpH/jsW05Kf6lBwLh35kZm3wV9q8cizdQCZ2ZM1k
bCPGJ+zaLLzYpAMcn8nTkQlqk1jL3H6Tu/buKwmJPRlfgHuVDihOMQeXK197kQ13
VqLt/Uv5CVmTclMgtisVXpFtBGC8R6L4vkyigxKRX7jo66p/0wUbCO0y6ksBMehH
zgvsKtydjSzs4FMjYd3G2GuUPHc7a9DDqn/5GJiNZELYsNKhHZgbI4y3e5VFiCGT
C2Z++3EMt1CDVvoFbuCQcm952DMoxA5AlPzewv1JxelaH0K4+Sb+7t6TXtALUh0D
9sKVG/oMLuoIrVODIYkWXyeaFfN6XaFBJ2H56XIlRfCr07nQiSj/LE2LSZh7eoL5
xpIWLC/sG+PEMdUyIX4siq79jqSZfEYl4aKZLjaVEXWQg8a4CjbFduFyJd2NGmPV
SuUm2R9F7AiprDTF05glugaaoYdBd5TZvxd52pdLeJoXGdHwPla94biHCryil/+J
6ky0UpQKSsj1bbR/SAaRJOj8MjORdOS/c/TTJqMqgAYDxEp+elklvEz/XnMlE63H
M66eguus1G5L09X4FlAhU+l40tKnk2GQZ0rC7WMk/cZ2C4Hj+Ua90z1Z7eXvlexs
I4J2rxvEuYW4DDbMbq1xtX7xbhrR7TOZ8WZ3ICDFEk4lRwLcj21VmXfbiCQ4WPSH
RkErimt9wexbraOSaq6yUVi9DL1M6tNJ5yTq71/07DstuohiSuxekgpmW3dVASxU
b7Rtp8Ec4Rls4nv+jwkEF+NtH2wEw+xdN46lxn4RdmwcB9XcmIG7nvfBRsjkgc0p
CjALmDXJW1VQhstembQ/Y3v4HWCL2zsrBP+Ju3vOLpbKiDLyn6oFVpO/C81UMjOi
8C7NeKGwRXR9ybBcO3MwZoer9JCOJ60D3T+zGKHd4KAx6+1XSWvfu+4lM0TmTikR
cL6+CtYNJc1Cy8ZnWmO+y1ZjXTQmrLCISr1bqp9apA+fcDoDeoXiN2qZ6LxVKEn3
UCCxteP7i6Zb5h32sCOyN6dmfWqqLE9PLEj2owmRohjmvAnqg0Pw+nZniuBGebrZ
sJNITogMTovu5ELnqtdxRx92a3yYkxiYTg7yY/BHUGN/Fra3ZibxQwrS778m70DO
opgWNO7LXOQvyCUVI/m0jjmt7ZxLZU/YIK8zxVCOnltsnQzt3m44OUm9H0Bhf1R/
ScwTgf7sJb5ZR0Yf8N5eyIZcGjlsMJc96Kiph39EgvimJUS8ouphYutqiKmtMgdg
qYoUHomlETg1LXWqITm8t+ninVT2SniA3+QocI5K2gt4pG6zM0LAxPsehqtDZ+Fg
1DWKHIQIeDcxLl549splMJpD+foc+CNDAygUm4umfiSJJhIB8hJ7yzr5xbLGm9RA
BNKCKLJnEfwadQUPvppjoz6Xu8PIdG+JqxMZS2JtwZO6fLAPg0ZlCKlU2QvytU7i
wCZNBDEZZw4uUlMhggGftwkO0ydI4ie8LJsozYervNG8y1QvjYpPoTQJDur3d0C9
I/fdq11JEk29giPKLYpqIff9OuJzU4y0HBlQk9gXhlVJm8WMwe07RPXJ2JNUFJIU
2qPZqQSeyaHWUSA9loweF2VVpWY51UVq1N0ng7PCCoQovR9eP/hR4vie6k3GyrZ5
FTYGBRY92aWNcf95ZOEggkYeWL94FnmuqJamObcrgMTxjT8Wx1cVuokFrG7m3gk4
HNv3r2a30VuDtMvz5X9lrbqKXR7VEpovvcnShmkyD54ets6G/IWu7UhFmSahUSjb
p8D4/wdDtCIAXgPcFOPpIm1ox+Yg5TsQJaDzY+HNcduemPo8bDg1nb/zMReV1ZhG
rrSJQEvBswMY7TkgKUUlXKxFhmFA+2Sv8ok4NZ57i2uN6OCoF/qZQX9UfMrD7+ef
X2bYtfypcdzoOoFRGhrRLaE1N7PZ+Ght5kUhPB++7COPasa562yKyiRZBoLvpbW5
pwoCCoIK+eciFzkMfanWvVkvpzZt2ZvwBUdjlFI+NqusznPKzfslgAqmL8qXipve
AbXILHap1H/uOMqJDD8N9+b66NNsM0x+E7pexoQbYj9crK+z3RtyMRAeKGbL2QzD
XoXSMcFJVLlUDV6Z44mBk4OE8n1MGH7SeQ83/564jc8xHSPQZ9NzMnOL056vXRm6
TLU9sOGGNPnkHbNqrfRwmOgMTLXCyz6e8revrTfM4Y29/SguJD/TSJ/R/afezJ+N
SPoSPNsvkg05BuMbOyUJLmgu5G7FFGFalN17fhQN3/L/FMYT3GOnjIX1+ieiwRkP
y4nCcLRp2aBKxfVIChRpgZZGc5JlXWpec1FxKXwJ2bfmaj/9kS5h91bVAJzbdvax
V8rNGz2ZY95c/uKnBefvwUbDkI5+m59d2NmQwYgra8oC2GVLMwIIiswHDQv9itvP
3oA8y7up3RdGx18QWvOLz9yNzm4UdHrzuVxyl2XeiWVic5yaXyF2ffgFuPOBMzV4
XFktl3g53DxupbfkICX3OUPe+BXb030g7dsK7LSy+63rBEaikz4NQ1PITPX4sxmX
lyAK6qG7Bc4f+w5tIpkfKW5bYiLF4f8SsxUDpfCqKgAIozqew9ecwdtZGiI8b+eT
QRajSfDNNyTKzIMQznYIUpP5E0aC4hrpV/sJEZvGNaeT3YT+40STX5WpQpWHL5z3
reeJq07C/l4o7pITOfiM8QckRer373/HITi94+QieJV/ZbFYBzggkl6NxRaScc9c
oX/kZbCkYM3sKkrT+sMYaV3MTQ27lkakb/mVjDE3HiT8C+C5Ngum8yaKdpF8Nx5B
wAaaw24o0xYAQYzPRe5ENBKyZpi4jjZQad+C+m9soq3mbZ4jfEeTmaJEJcYsEYu7
SaGVjVJ37ACUeTVicngBiAdU6uFXfT/22mJuym3yLyFh1basiasAN+q3u9xQw2LS
/nhMWDan+GVrG3MIpoetqpKQI1ouX8pfKdXnM8NXGeCgvPsC1uTtoaVIQTpSW7L5
pbDnOTqiPC0oqo4jhY2yYw7kuqSbidW30xoKYtbOeTknRqpTgoNAW6YdV1dgWMY5
d5SWNWryQi4deq/lxlz/fZmoLnWkfPyMSXppLAxPp0OkdpFhYXHgkm3ydkHzp18C
Pn9DOMYBr/hpkTfq2iS+QtX4DPaY1QMqKW8QgUd0m25VPALID2Y1u78KFvhi/U/4
8fI/BZqUKLYUgPnZdbpTCPpNZ0j4VMr3jOd2P2CC00JNqPml+/+Er9qAdcWM3Y8t
ZndonioehW9/EcTK9hvc9aBB+J6GL9IjJW57RwZnzcm7Xj5VnjL3Gp6dHZS3inN/
zGHd+z3uWerGZSLmDrkafcKxBuNDSp+WG46tsYGOWMXUptKN3GmiXcZocbYDEvU2
mJ4vT7yGh2e444/P/Q1HTxiUv9Mhwro/L9niT5rPURHTc9bXSksjmbbij1s7BcbB
iYtYhrCgNy3ZGJHvoeNDzmvYcxbJYI2tvncvDCwgpQBnIE2U2BXHVbIGis6ME6RO
AMAH+Ec7Y7ZSDwq5NFMmVqHogpRHB8lnW7MieYT0lMOiojAsyFy7t01FJAAUUTw+
VU4JBqGoXnRiMB1BObU9i3mS3nIkVnDqlui5RJvrI+sNtWtNuQtgfNtrcLA8z3Re
egKAgMALbIF8iJgJ0OXGumxs/2pddd3rH8Gitmpk4oPIIsxmt/Ughwv3a3CCCcHF
CAdaQgQ9//52Kns4wTJN7ccJt+4dvReASr2FThpyFSmSUTpP5cONdqlknVT/0z2U
5Gx5KhQtqWOc/pNiVHQJCUve9Ldli708PkeJmyddgBk5GAKaMH1DHSfPLBpq8dfF
16TGiiYGNHMRABP3MuniktZNNxayNv8TwVGD3AabxirtCH/Fz7WUngVf8lFRLZPJ
XqgsKYR9SuQjpUUPNbgulSLyjTM7trnaWwQfitxIuw7E5lsKCL3QI626Jkt9gmPZ
ywBSHgY39D7IVocnqsvsN+/Xnuoo1JKagXSB/OD9dICtM9uypw0aBZkW0W+MoWG0
8ydysip2eKEcix8nSRReDOa47vfn0SBqRPtZCn5JbRypWwTh40L7qVWCiRri5POQ
O2hTiUfeQddWGJAylzUONMxwoKkItc6/vivh5k7r00GiCF3QHHUDGGqpm6U/zyHh
2i0+Ewu2ZF9c2epNFVRJQaewCNsmooOa8esqlcTkZmDUb0IVjY3+w8OIeAOeouT2
p1Ih+kVMNohfI7y5UuAU7r/ExQQ9lRBJx32hoB9fUgziJ28HwBWQjmUwcQmfwSpm
Ylgef2rQBJSjQoGieywbn4Z8h3/MhCIoaNA65fRg7RzI/oJ+FCwnc5fKJE3sdj8T
fo/XvmnSbRjs1g3r06q6x+dptw87Jj7OSnXbJMuEUMMW17Y3hs6vS+ZL4jSwYy2N
FlrWODvD9hXiY/4q+pwD7MVKKSNv5v5KX+KjvM/3cfixBjLcK6tW/VhmVUxGvPpz
VAswpC2H/MRBezaVRgy8GkgI1WZVQkZtfxeRuYtD2v0aqlLpjNtTuBKPQzoGvfr3
c8nZlSLnsiVj0OSL5Ax9pt4JBuKVO1o0AQodwRdKJRcFNyVymv9jghDT4aCfAWYN
UVaVqFd67IH4PRjj5m44sEWKD7ySWa1UPbj78rtRuEvnhcSoFrQ1iPtJcxcbEKfR
0yA7BwB9vhiiCTltoICkC+w0XMGVrVeWhwoFLnS14oMRt0WYbe4yfd55bX4cEzBS
2CIWhmlM8duUnYrNPS1r4rhJZJX+SFo6QvdHUTVL3t6yIsiQO/mgypi3jivoxBMH
huFMUr1tpu5WiiQsNRO4t7AZRS5yFI3HCgoIiPKZlzh0mJCCmIynWJQo3hdtC9A+
0f7uD4pC1LieFDe8eNONUZjHlhNRGhHAWQRX+6PYz3MoG48jpP6VjLJyB60EqiV4
qU2uf9xeY7Uj7dS4Rn7+PZv8+rM3iQhK//5NQrlPHPvUP0373x1G31vkF0CCfYmq
aRsBUMKswH569hO9ordDdalyue/tj1HWEroQZrYCpaKXk0XNlCVwETV1puzeafxT
Y6h6Vv2nN1aURT8FsHXNNNt6DYXD8ee8MXjkO0NEEW+DHIi/8v9/5Uh0qMu73dyL
9RrwfmGzNwPUMbetGQwcfTOPcNrRRMgiiZafGX1nb7qOWCwTAjTITaEU+kYI/o2c
ByPEvIcsG/z34p9zqIf3hK5GTT4UdFZG/q+fwbqJMJsm4tWkMoxu935YpqZPuE1j
cJEEGjNXly/t540rWUjS3KOlRSiZAQ7z/pa9yO4cYaan8pFbC2X38Y6obWeGM6HT
8bueTigBSFss87d6TdaC27rNmpRaT3YEv8m0AiE8HyanGAO6e5fE0rakSaLYO9pC
OB8UTNfaJzFcMBQ56e/9kYdVAkVUCtIY2rwulWe+aOJ+D/Ye659q98ZmVA8eZxdn
allrnGCm8h6xwtomVoT+xw/5qLGkXyAdbdXapq+fR8Oq3Qj9ReblQiT/L2/htflz
hIlbFalkhPGNZ+xsQ6rCAuCf9v1Eol2F03pHsq/rzjIstsOX64Ro9kb5CEr0dPos
l1aWyz91s4on3yu0GWJfsRvFM9Xe55oadIJ1DuNOlH7PKJqlZwhiFRjehZDykKgf
OnIDoe/S7WZCb0Ki/nsAr8S0x4PpFfRDMkCbItVQ2jtvK9ljXOeDVqhxNymwxa6T
3EDSKD5LmdVdy2tujNnvNC6QgImX2cVz7J923+7TwG8GpTKg7eBh14E0VBd0lBrw
HLL9UfUiNtBOkef9Sdb5W4djv0a5eZtQ0dReIQeDX04uuU2U8GmWwyDnfK2q0mH8
zekZdVhg2LvLAdXx9F7rHw9ybsD6+NSsQdkRI2UQpK03dcjkyanq0eusuesFZMyS
ocm1i55fePphXPPQtrWbpOD3qPEISTFFQPAY1qKdrAPHSXXz2dYBkc1O5LH2l/Fb
WqHBFPE+H1JuMNZoCyzSxA7DpNCEKncPItyozn8zAQvhJc4pYx9YEbIXJJjlFmTG
xb2z9CcKvCZLRTjmJyn1Z376EJB1vFGAtPjQIgXo3+ibmEuvmLmi7luvOC0HQPW8
y+krfwG9v4tr8f5E/Tb7JQ1zCdHmjMvkm7wxq0GPdoiUcpaELjG9bu30O+HkK0cm
e26ro6UR9yFk5Zwdw8fmnJ+nf4gAaxgQqErXf3Jlz8BUAwbet+v6ZR8D8Cr1ddsy
O4pHtqfrfPqvgtN8KVuZmPLi5kCadeuzQrWsLoNyBzeFvGG0q8jDfMibMC12e7Ed
Xpg691vhhusvekLu6/20ddm/PXebtI7PVFLtV5x/BahY5kZTk9F8AnK7bFDKAHXL
79IdscHtuR51uox/EoY0sFC4sC8LX6xJQYDnTNLHbQvwFLCPICj2lcw1DZCsmafI
tTxTzjgUsDAre11UPA7apXS3bceoAuIQHmB7svHbdGFKOHOFvilCw2pUjDTK+jxv
4BvTkM+5oengQXr40ysz6ayG0fIyU9njp8A+B4sVWxReqDCFBQXGqhoqhqknVN1Q
tWfxMd/fd4VJIR8CPvE2ZVZeY/c+dZ+r/dj15smog1QScwfO1pLMgeZ6Nr6HgytG
BxNEfhRaM24nhRTgKknM5ZCXIWPjYAIXtyok8UKaBDnb5PAo0mVzrWvC8DwWtWR9
hU7+00uhrulGRIZP5IEzRCGyKqCGyKBjZmc+CEd3fe4TdD5rQh1PX4onleZv5scK
TczuUa09Qzs2l7iR9DKobbUTYac03DuHVDIzCvDzHSodoCL+zcpTLW/EJ0x7YaZW
8On4aJaUNA2SUyb3KnX/2w+iYjzr9C9YTSK1rs4YqNYS/KwtiqmW9aNKwg5g07vx
88f0RqIY/Y326hN/AcFDkSyRsFI0lqSdfgIQh0n8CnmYzQ3sBRbxbwA+zNieUXVs
8Fc69SsmZTDe74YL/piyPorPqB0HDRd2U1NknYPmrqYQ4nNbwfL5EKt/goQ8aVBN
SLcJh2PlzAnaMlxOp9KaEr8AjGxUbErtjGuSAK7EB+NRsINXM7HA+VEP50nrGGDE
IGMBdaYfs9YNNZI14dY5IAtTHaaR7d7sB0lOGts0cKaEXYiDAxbLaPqOhHCtk3qq
EpdSKuzUcttskVKDdqGWBoEJ6WppIcgIuIM5G84lGHOw1FjAg4jreZIqZey/npnw
ID9hlRa1hoOrJhteqFC7/kV2EjfgwzIl6gX7+P7EMrc6Owr2byWt04nVAsMwcbCT
cdYmBOlS76Z5G/XZSSnnmNW4eMDhO8Gn8YJOKTssf06GHL4gvvr0GWUYkB0DBYKO
Viaqt1f01lzfpV8XXdbwqr0tVS4L4a8Y8JUEowARDC/KeiNmm6I3BZ0pdY9SeyUv
4Gw+5wRSw3uDd/mUCsKQ5kvn66cVlaLH5ZXSG3pSVCaysE2PY4w7+PedU2Akz+zi
tGCtZKh9ItCAl5MuSFVan1DFbzCerqRlVTpJZ9M5/OG+YyFvoOaWKCHFBsNP0yky
I/efPL9NBnvYd4EqmEUXN17yU524GpfgXpKu2e3PUwREn6m1zUACjRvgvC9Rs97G
U99VjIceWb07clHTaV7GgO3fi3A5RO6N/Tu/9J4DG1MnrluHXGaAfXyg7CtoTLvm
+gxUK4nCeCdts+B+qnvfx3DUd9wf+HBuisXtwcN/lrfiwwbpUk+zg6U8TNFWG+/b
bsR9ZryhRLMQJOT8GFGMwCkI4yZl1tAUeI5ijXmGywsrnn+5+CuDYPDav6Trjpfg
pNvZQSv3Fn+2Hhnp+7K8qdI4RIsPW+uIklCnlpLPuAmeZBggYBDhkmuX3tuJBsCi
HZ7x7j+dHzMgR67xpDWqMIWWW8BSEYZyNgnpGixQoCOwFLeO2puFpfLha2O5kOX6
GDg+0xT20nEW+x2ZMZ0j0ipwblPyiz9rATBy5FARUrpBaTw/FzGk+FMcrhnXqCU2
HQWHeY/QOydsfMXk6jYNYeouDdhFkENaZpLc/3sIpVF0LRfAQnF3vv+gjQsWEGEO
kCrcdwEf5vm+QciXYDagDy85FBC/p/b7gTECIM4J05COaD5kuR0Tl0f2uOnZAJ8R
RoZluQ1BHqJIVOakjUMjqTrsXciUF/22dv9tD0qJixNU06PP7hwlRigc10Es38oM
kXxTnA2yRlJO6KPTR8PWXP1Um5qZPkW4dyZCSY8rgfJVUabUBQgFkeNHGz76XqwT
VfAQl3yn5c0w5o7nOfZFR960YNcoX3dXt1QTb3Q4U3kcFLmYHNBctU94rlSn4/OJ
bbRop7G2WZO9EqqlPDli4HphWO0to7B2oGZ60ugoPcrgrqTwp9oIK+qzhckTkjod
Ul78TQF6B3iP/Hx7ab1G5KPGIXpwkRv8esn+l24PHTRcaPXZ19ysB5DSBJmZIfM7
dQCEXQwpajrVDuYnnO/ALPFLDDhbdTZM/i/NzarHhavf3FF6ZQG0YZxjU2WXIPuL
pKUZ3okbuIQcp8+430wayamegqkQrJ5N/QahVIIVVBkynmw0vsgz2+RRDCUvJFh0
zkrnj6k7rCrGwm6MuA8UoEGiYBBwDtNoKbbyJwLmPfdQ3Fyi45DSn0594o/Lqt52
YA49zgojUjHqil3sgPDiOK6EUBgcV8QA5bnE0lAgJ+EgxCPdgWIXFKxXEJBMaNAw
SWO8CmnxCLlLRKJWGaytQuWFS/jdXFvMtXMrOGLpIB5uPHWKNNmhSnic0os6uYMb
onjcLvwZYU3UVK1Lf3BVpIREmLPoojLnv2i0k1JJLTN6+51kosm5rRzou2AFTDUW
WZCzeWg2QkKmpF256sbD/AQ18j7xbQKtaf1SnJL/SJ+tFEvJ2UagWOaTBVzqEo1I
let2DMuOkhQeuWaUBbsY6s1YDppsMwRkC1pYS/jQUqYomOYhoqPTSd4jurZ3+Qez
fJI4L0+fDiRYYhcvx2qkbxm2/2wj+VZ5bBF6/17OlhXTIDQVhONcWI8VkJJ/zWNY
3+D/gJraSb3KABbcaF/BPhnbui9OcacpzwiuhHdVbw/1uMksUKdB9XWJ+6hNvUJa
buTuP33uXHOqy88xab2HpmuUAnf9CBpko5bDn9bTA2VQjPrXDlkf11y4AnsI4rLo
QfGGk3JFwdKDW5SZDpL+VL/Z8c0lpyEDgRjxJK8Ol4FKW8ubwXmPesT33I8qe9UB
PiJqA+NNx34SeMeGJe+px4TryxsNargnuqVL/XaMkvXMEtciqUAWRA5SjRpr6lRi
xV1cNtrhuJshymZBCzxhuJLGHd0rlzJT4qUS1HLFs12M0Eka2JlQJpYRMmJemnNG
Jx2nEr4RNgB1Y2qgwUSKmGM4Fv+8cI392X02n7rwVW+d2JSllEzsdv9UZPotssmt
m+gyDOfjy19IOJQAOmac30YOiokSXeaa+IFc6wHWLnmWeLVUScfOayK3A004Tc9l
5zfYBvoXn9+9xp775UCk/N9f63Gux/H6nHBWk5na5zmPtUfgULxCIHvVoKRHN4wG
cnMNKQxXkGgy+VE00Ods+DsJcxznwVxOTQPGfxfC98Ec4mvTSq9utN76ESr6GW46
Zdr8qHJpHpmo1ngbMjL2OdNokafELPIak8NFkW/a1sFAG8bvlgZpNmZLixFINCiy
qYuXYF53j9H2X2KnbEJqJL1uO5nBL1WVzY35neXVYfaz2VMghawHF3j57NVuySUh
1l8Sh8KzjhpBxd2dhSijxB75BaQ+sP+utb2M1in2u41f/jv2AJqidDcSJzfTX1AY
I/n7IuQj2JVdfaj7fkemO1nc+keI72OdKPTpuP74GVi/kMC9FWLEFuchN1wFUndj
BM9LmM2Pk7icU22silcn2iCBDBVuFrrjllFbU5K4o/si83xA3miANyIKU4uuB1CO
Ru/y49squdxk/+bLsYpp6mb+7LChyb3YzSSug7mIqsiysnUlZZHguV07Rfx6IXJX
dcrHhp5f21M4OhHcwLijx9fipZT2j3BGQGxy/zx8ZsAFkSrR4aHGKkRZvtlcj50A
4omAQeO2+CxgZ+RqWYdJ7bz+RHwT8t+Nxfv2UIrpdX9ltdWoYzucQecLA9+FxpKA
rEirlA0G89EDe8c/cx9rj5Pb2utv8uFRyd5lAWTDDmrlW7Hs4JNW/Y+WNWEJ6xIr
HL2RVDOdqd6LXxD/HL62LTVddnZMuKcBAYw5w/xINh0+DmgYASj/ORnvl5VxZNdZ
OKdNO80Ds/VDokhJs8cIbTuH84GZDrXsRGZD25SRakJTT+JsS3cGvRonNoYHYLcw
/ZE8hIwVsr6gTgydGtaL4URUIX7e9tFjm1N6wE2lzPXkki4anZatqH+TtazvCluC
8cPs3u8RvGKtgH/F67IALGWjZ8yecC81OLAzXK/uFyMwU/q937V5/G71UAom8niy
bEP6gMq9Nl03QqnTa1iGwuvCFhjVkE3HljLSSzpL5na7j/NgOl2TuPRm1daZBvAA
g73mN5uTcR9WpEFr58cju9UB2XtY3bR+scEaRYnVLQFapl4gOiZvX3RGZ6ZQ8Yyw
KS1qMR64eTvlDAyNELsaSifAr8pj4cLqnzCURaY6e6/Gm+a/JIZbaBqHMWd+naRM
WBfGol9VLXi3TSMcbGhPrZCyscRw/QNGfayLf2QeoBPQW0imDTDG6m34w4WKcvjh
5aXDoan1LuNIdC6UrmXBn0xPHFOl4+itIYpcbtWHfhMzdBYdFZrU8HozuZSIZt5k
w5+4rKIPfh+63PUaf4X6n1NgnOVpvSeGZ2c6hWaGcPZW9Oh3iHZgD7BfMAuZQ5Xb
5+bTmvydWEKt1eVnML/21jpxQke6lP3LS7IRXQHr5XnVBD4Cfhd2t4Nwr4wo8tqX
lM0lQpx1aDG+ufkWNg+bpONKFs1vqTQxu0jJJ6GNnDMlgJeViNiSMMThCLHcdJPR
pd1oASemWI8E4fdws6nZhmaeGgJ/zNmJ04vMGDlt4GVwMkelHrpovFJJsnyeSQDC
zZqmBB5aFfzYrhoCVgyr+YJ9KpgA4dQHw/8nn2CaLSLWeD3Vd+RkRZMgeWVxDaXH
gU4OZe2PzqUfx2iAgzjoH9OKiYctMCJ24qoIJ1WrifleL0z0a/byAgr7vbaKim3s
DRMfKkhCVABtTNC3sCKV8pDNrZjOI13/VZTO3cTxmLOH3JvMw4AvvQrXPZjn29um
qOKzvZqIcCbXWll7xdW2DQ3MgE0GGxouAN9N1cazewHwH7x8H2okDMG3VKNNnaFo
sW5B9zJsI0jPKhcys7BZk8w+MKJUGayZjWTkosT2oIJsaFvcq5tqbcI64XPrSMrb
MFUPFznUP1ETd7UY1yg/4vlRm/k010wrBOg4vXBylYzoYAPWahMUUEWIpvVlaE9r
KITiOsheRGprbY7wMUXKNvqHcHYgI9pCSor5CcYkdult22gvlxEuZ9sELMpaFKue
V5blAtJe41GZxESzn1fBmPTuICntilQ7GyiEwkTgfBF+wqSlGlpnnu8012oBpdkH
A3Wkmav15Tim2wymQjz8+sNd/8Q/A4+z8TpL1Sx887kD6x+P9o90tjeHGgmDmEMh
eBDiFHxZOC+9H8hCezQIYrm6YlG+zm3qT9NznhWCFmnoeEcH2GaFWeZ/faZANsA7
TOAuLVYGjtLhWOBJOO6UtEiPqYGVfDRtFy5kNQ8KOlL4RLjPiySMvwt1K9kUo79X
T63gh7KQbsW7HiwH9O+H8X1hroO3zUJ1rkydrieAlObqAkdB/r4JDaIcvutspyJy
4+pKym3CbumzOVAnbeAsECCkaHaoDBbHaQ03f9WtZXCadJ7QD7N90/yq2QNdiVcR
xXKQRcldhQgrQMbXVsmd5HOnjiP/8NXkXKFBZbPYi7yowuRTd2VHtL/t/2fsBGMh
PQBAza6yUw/jdqHzyNMW//Qkq2wgF9rNlVhodw/N+1WMv4ZVdGACgI0yFxQ6W7F9
WHZ2WsybtibLgFBmU5wWChjDgDe2Tv6WS1vfY8KaZ1UVAlHOrMoEY+4/qHm4RMU4
ONSZTuofuowctgEp2iujq1WnJ5jSFznytTNfLaqhKLuZdxY96mIj0I2z6PV8Puxh
Gdk8bP/FDzfcpZ7mMqoyCA1IKvWGupx/L99KtW9rfzv1dgXQyuAwb2zpCPP8KVEX
6gO5nHBtBYl2XEO1pNkhjplUxhXCRHHc61KdUrrLkm825M/an+xtm/08fjwedQPF
qQiVUXeasJxK5wgF6OMSe4qKfj/O4pvPJIAygoV2VqGK1zNRKX9MqXqhn2g9P3Sn
ikQsuZgzZP1iI7e5A/WaCvTtyc5//76FUaTsWzsYOkH+KeREwkKm1DAZOigowz1F
319wY+XvmZOMDEhTmp3++a7MubtfvQjRjcyzlSMZJ9hJN4WRESTX0kGpNE9lDQCU
fr0ejajKETtC7scODu/5BBtVUtOk4q1ztSfmks8/t5eFIOIUDB2Wqf2+cRUwZE1F
8vyyjE9nsGD+cCHlY5LEvGMPUu+0SeHtVPbTwP/M9MmVZ6v410BJ1UiYSPM6Q3R5
jYvZqqKLKB8ppr3VW3wULWk6SPPHLvDS+byk+ARMy/EFqPbnsAebe2ckOWjtEOq/
ecO8Olie9CED7tvqZpAMsAbZzDGybaKa/P6C/tlzhibSIBii+JqhqRNDog6pC/BC
bSbr08ZlZ66BtwIrLoEQcfssZon/TbKomjqA+yX4pdhqDkdFCMVvpL2yibU9we9p
VzWaEoDbs5AriBWHfs9YGT24qwgiFohsMoL1LpHpnCrQqaetHIzoPljhQNRvDqVa
UtVGcV372squUJy2yvPGCda1bpE+6TZCN5HguFwgdRimoFwv5D2gu/2l2HE41OgN
FZABeT92YSCoFfUQY4MoisGREfbFb1hVjqjK+mKnEHTEPn3ppKbC8IJPCcX7GxpL
05DRixbsys2gPV5nOsb/3M0DSDRq/iyZnO9ZFnDL50lk1pt+uSmlVRZf5OZmEM2f
G4Lt0dTz+8c6CP4G5K0NgTuSfxHKWoGJXEInebJ+IxK8Tfu/g6s2MlGUi0QmQdb2
muLdOxSWjV/gZmKbFTnDARSt6xXM7KnfJi3Z0iWCcSBbAeiTRZo9FzL6N+4gGB+S
24KltZHLrGRPyNfcyRtjF25neqBa2WjLm0J2QJY8VdxvQUp3zDTSDBq96skzQdod
NpL3JNZbmBsqOX5jINxWnbDPZ0aFuZJH5DzSQU0haOzIbqlxTH1/I7SeEybhgsQN
zURo2Oh5WlPmjhqsmDdmvUvAN4RpHy38sGQQI2F6ldbm5mM5/qF2jQRg5sUVtC0/
+wPakDtUw49KoKwIsONnm5Ilgh0IWyh0IGufeRJzdQGNL8K1fW0U+jFZV9Qq/bTe
Wb8qHYsoCi66u0U55eGrW0uTcH52oNCHH3FO3ZfALkI3V/qmK2Kbaj1lvkuReBmF
KlDm6lYStRtzSfhm1uFmrp12KcbcX1ScBoLuWK7gQmQIdzXuz4wOOzwEhBYQ+lky
qAjwL2LqDCGSEKHDYBO8fexey3Z2y9YFDABffbiBGQI1O2lN+foyTDfvjxOmBCQ0
8lP+jwHCofPdgOQ4RzrjnXbDn6P4kcnHb0PCWsMOVudiMv7qGS2VqkJy6kEp/JX0
i4wxBytzYCusvN6lT+28YsOzpBImPcJ50wrmkh+8JF/pZS0GAAXjEb45lfrWD6Tq
fu3Q4c7v5v82hpvbBADyl585yG1eI9dkfLCD285dR49UCObpyaMxZ6mhDS1J7JBB
1sTGZY6YaKJOATOU6VaHjX8Udp4RF1zG7oIw70DyDWUIt5IiTeB15bhRXTQUpMVh
WmLfS40cPRT0RHNinOWink8lGhP72TwazzNbN4jpxklbCW7BmYW8mBmsdorNPAr2
auL+EvXdvCdfFQNDyqYPAiV6tOy+lmsG242aDzY9uq3ZZ8abaPpkbILvs4Dt19g3
NYSRbkL4oBQzp1LLHo37p8vZYu/drXF813L8Q0anVqQD0clH+IVBCFenH5+Pjas+
AGTQj0hlcZQ1r0tpspKbuAxEOhq25Jty2TViqQFMvXKuR7ghYI83KCDmPLizGoq1
HCOyk56sBWLnG1cfEZfeo3UI3mhiMgqbHLUI0xrBGXLX2SX0ePROAumH1bdAkTHm
LffEkWgwiVvowGLt7+1blKrK7QDSXSz4uTWsa1Fgf+3l38iXRQmWnIWF+5EkMPiD
vytAO1IHSViPRRk69S2tA6ohRpPp3/r6DSPQJjYGN3R7RrvKHtiwoJde5X/gwSt7
ioVkGzoIIzYPM1kcYMxvR11rL+WRCKeIX5AdMKzh0cwdFbn4hN13S4l4IGWn7JP2
43YPLpmT7Ee5pl5abe6K6K2NF+LrJicdYe9QC89gz3VKKt/QdqgL2AIsH839iLVT
NYGWxf+9YSa0cTnV6GXGq0goa56O72WrpEmXojG7F7TmSonMHAa0CPYqvRWu3d3h
25SE++3ZsfyX1pK1e/5j2cREXbXMOXTE1/lByoKUa5A8X8SH643DIB9/aI+5csiE
Sg2CtJ5i7NHR430qS5NMdpKGwiThmYKMhP4rAeXbJtil+1qL6wqbPRFG3kD5tpUv
1Mto4Hh/8w/ZSs2DpfmE8g3k2nUC7Zgc+8JdpCallfsiQh7ASkDf8irQirlBOUKD
7tcV/tABn1ax23a31N7p2YgcGUseH3NApxMhFy5mm6S/zLw6gOYTTq1Pbx1oau3x
j6NcaUrTi0vcOSezS/RFCWU2zyCjVZWP4Eg5pSSWijU+9azNb4ygb9wRIzAUf0ne
NTVmcXozLVe4Wndss7FCIXuxNaUH++W6fLazuv8CNaJcSQTFzDONF0AcxQadljv9
iX5toX6RmtgOdGr3l24CGCploXfNKLwW5ysDBGxPgM0WIoVHO+X23QwnJze/ZUeA
lEwF0NAaCvTl4X8KqcW0RdT4TEGFjjjbnSFKrm1xVLZqQbXWVIZpS9i/yitUyFu5
PL3f6y6129f5W5r3hhNGLOBnkyvLhDiDuYIu0Yfu2THDiM/ymf2296RmcugE0Bqa
m+O1f/ccwztlYBl8aqyczoScZjXczu07/5TLEd0WAcvn4WePoqzZbvIpx/2hYWGs
iPOpQDaurHgei+gEpf40lye9EhbLWR/vSfxDXCIXIpnfy8LhFk3Y3+s6GWnKy2bX
xra3SbArzLKd4eSW/n6scCGqdG8H+iLPYAi/gwfUxMOgnhPOcNSfFOLe9j+3G002
ODtW0Cph/it1Ls+0x7GWGim3pA02mrbZDbIO1AT6BM4vh3TPp4/PdTbVini0BuAY
JAP6ZSPTqddcUDafsfn3vEDtt3nmd/eBnxjd+nIVRlOFJIT8fZdvob3Q8ngBMOOh
ut7OsY702WYEps7fyrjAcXWjexvO/4gGzm6JSjbWgwUlrc0wPLSg8tyC6BqMr7kp
OAqoQiRoW9U+BwUCKx8yQpyg7rVVehMi3zvaQuM2jG0Hp0bsyd1gv1+wFKyMzoiK
PBEE/UXz5yM3dF6Mt9luGnkL0uh6ZZANGifgz463bgBRQDz0saK/EKmnmwifO3rr
59ujTLRe/0cRJlBM6+vnGMZGyFWpS4M8ALWYl2woMUjVTkQSv0/2c/NA58SU2U+o
WKWsLFUYZFxQK6HYIBq9ScFJOp5nzJfSPy81gPEJxUajva3PcUj/Pq1PcEVVvnYS
S1XXp31ceoO51sdGeAzM9Yvy95Qob7NXAg0Njh/hWiQnA77h1y00UcSRO6rhr0Oe
G2OYwy4bpz9mGb4KM1lfgqSNP+qLTYM+tYPMxQzatcsM9eY5yklJuwIJ8OyXZs0+
RuIlkDuxi1IlkZsfv6Do55IAXpG+mB+k6aGJtsMYSyBYfiK/EPFME9zGQrFXsumh
PBv0vd+8TIW1aNsh4e5h++zFw0PnMMEzO78f41eq7B7sgnR1gRrhnnk14S38uZR9
pTyKW32am1Gtt0t5oDCsx1ghj/AP/u5EV6k3JU0+yitohZdqNuGUdVLLURZPPXDQ
lU18aN4TTn3pdgVake4m3yQKlMOHsHxGWarbFPpmVKLptZ/yUQoUoVy/KZkHmpWQ
nM4p/VQtWNopztZLcx0fs6cLeLyf6e+D0MDXW461jdFI9NO9nlxs1zC764NsNdIb
lSEG8O8Tb3p60/x6AUShz4qWV6TJlvX6UxFGzLcgmLlGMrx2stIOEXoXo6nR3GvD
xD+928rbZ+BJA2tcmSTVSXogJ7DBVhukU2zhT65bAjxmfp14pXgWwYKPxRnJwNgN
2MeAdJ+riYWNtb2d8C00yeaW/+y0J1IyN/VmIL2HmdLWq7LHLHcGAT4+QWsgDVOz
AHEgS2qlSXpKMHXyoIUA3reD/NVDomFZshPhbfD/h3HxfYVOaFJ78JHhbF6tvTde
CTWA2c9A3LvLN74ZddrKAm1s1aVtgKHDKs+dBUI8MCMjVW8zihQUsnNLy7ihg7Ux
W6ZRh0jjAi6g/4QbTSN50Zmf9DXDUNavu1rt03aMpx5HLnFg5b3YMOa0Btt14dEw
fpkN1LXhIYHnJjfBpcmV1mKZ6vBEwOhcprCNGMTM0CyCfgnvoboQS7FN69Jn+NUb
bNHH5WHeDnSB1UpYpjjRrhEb9eC4qsi2qxZDi4aAVtOeJ2dnURGaDNZIgUtqSwOX
7irfndN+8P+VuD+zSz9uuI7WNuIanVjLE3SorIpmnd5jkxDFo+cx5SFv57nuOqKN
s8ny1fW/ThLmn0AkIKJlK27D37Askr+J/I7yDr2EB3a4qdFKOxUEgPzRvZIXXdkR
TxqHC2vOXKMuY1KLuKKlA/LWr85vfJuzAxGVk9ErXX3LBTcSfPBgF8JKhOyVFJuw
go9LWruU0bZd6Hd8tXMW2amRELdKuwhBDu0oO98wJz3YpHJOmj4dlA5cw678sN5O
dnojHWqzvENf7xo+Ix6Qf1uisCy6uekb4DYx8V9XEQvFqg28oUrtP+NFTpNbFvHz
n/qdelPDC0xKNBsTZeObRCwMr1sc2PL/t7HmpFUEjYMOyHHVejlbQy364U58A82B
aMjb1bAUYymhUDBuUYmA8ZPAykyTWI9iUS9mTUhwIA6X/MlJhtDzsR6i+sC9skC0
fCoEPqB3Fp0JsrO6/xdX0ScSL7/GDBlkQaK0mAf/nGbbwV4wu5scg8/2G5Wt5r00
IPh4aDMUKZKMda52Hmf5KRatyuFi5XlAaG0J4ww2BHvcNdQDlg2pk6lCaYtXnWSy
5wreWAUOBFq2oxvrWLXmzmT27mHyfT3NAbrG/nSVCdrSSZVnoAnm79020ojZmV1y
5GSsDBDrwsuMSrp1Zl/u69rQ6mm3B4iIkEwscMw44TZgPKMO8VIiwks+c75V9AUa
5jDJNMVRBTe6P3+n8is4DLknlbnsvqmDtVthmVq0KQ/GNKE8QbNHNk6bNe8+DORO
mIndW/LkUDpSQEwKFjzWvhrTWYSjarkBjxlPD3SKrXM63y/JGhbvSLepYZLslxE/
a20CUqdo7km4OMnmLT1Fkpr3dqL6ac2nDoDBb9KfPst1Hlf1VjXpgsKYEH6J6b9B
eeZH/czbLL9l4BJpFzUxbGjKckyb0mbcFZBY8YLtkTpIQD8iwT5Bie+oXlZzffmf
I5SXT5YOFwI0xzxoPEfek8zRANdPb5071UrFaWu8mwyAch+FLF4iJ/0knfRDidCc
lBqqHBgUFUK5wXJMPJu1EIsFK3fGdruKT3SHq30l2mF2TqBeVZMXqQxt/oinY5JB
bxGbBXBgqA8rE+8Ho8wvWhvBOE9NhqhmbC17fulz7aW0V7nGxfExTUMjLuy/O9Vp
JyN75kX/9sWY3QWEY+2esoLVfG8FY/OgVEGTJMrlxspkkPDfbGSAJ/ky3620rgHX
Q/wcQbjb8ya1W9b2gz4MvdirjF6QNGQYTvOdvBGPrG6BLdWLu0aGUGQRbIIcBXpA
RlfmwpiXNOEAvk/yK32S7u1Nmv3iAOVpYLuWmxiDN9x7rcWAwZ8pHvPlYZiufY+8
Mxp0iskH25OAhoXq+54o5NAsQdvzMq7UJJZM6ZQORE3c+TMK5qSvKxJPbkU3FLmP
XRuGB0C8q6IhFdCbl4XNusl6COpBsIwO3NDVR4GHZ66Bz4AGRhZMmJzVcz4cY9qj
rO4gAAT0iLgQQCegk+sx6sOJt8h43u41+Fo43CsSoUrYRnbjKA7ysPjFlke/5U2P
a/UQtNLTWiWGVsFzhZk3Lj7QmI1YgMEsIEuBqCEwbQ/Vh2awd0/LvenrdVNOf82r
wntQhs8mnGV2A/dw851UgotMihCG9NP62RDhjGNuQbrPOvsyvX/JzNP688m5fRwp
C/CqMM00OLsM4lQRzHQ6TFXrvNb+qc0ZuNVNktEvCGi3K0hFaDmji4V8OZvgb52P
KTkaVMN5N6YcmxCg+0svG9fByCd536ARwrJiPY99Fa9LHct2ASquVxrMaZiQX2nH
ormnV21Axxup85Ui5WBtMOaSiTVuQCCa8pbZaSCuONVKCuFIxDRwzHRVP3qZ38qW
1gDQEd+BEtdG05xVphcH8HrFOxW5BlchxtA5ig2KL1geuxmW2vuJbFCBDB2ItsjU
QN5TGP5T1uZvKnf3U3RFyWAY6NJgf7//TIy5OXo4wzbqXIGX6z0P2/nij8Q0LWp/
cWPV4Sn6WP0PjOZ4Vaz3zaHnY3zBbVxeGwSGTViNuPyw97ygs3firaYj8oBVuNvD
AYGvMcRN/HLzH6m8BskFFw2FO/40FQhqzMx7QNgcqAWqwAop+kVn3+nKmcYmYUtW
w3Vx2QV3VwXvxSmdY1RCZ9o6PAYXGiIS2Iav9ZLH1j8Gi5IpzBBSXrS/gLKZ/2Mk
DmwOOHEBx2F3SNnu9IJ+riIVsV+f9H3HRVC80gOR1zExCNfpUSeirZ8K0luuz8Q2
z+V7/oXd8GZCcUVYFrNH9wWNT6rUS8qMKyHPe4i51jW8IDdJXdL6u3R+NP10uf4C
/eobVFmSh/3NsHnL7Lpok3EFSyoAgcB1+gRb4KC3PuRufWaMP4dxksuv1rG1bfZV
jne9MpuDTcgiIgGGq/3BzFrULsDl/x29i5crlnI+H0REE3ihPaD0sql9Ze/jNpha
/dlpg+lKczPSik+ZyUdlh83GRfoANiUJuZuFZdIwe9X0IqExOeFawPg82K3cwgrs
EBbWptwE0mOEHtnD3nROp0X2u/Xjm7Y0ruAADzXJufTaksLyOhHvG1abx9agPcE0
mNXjYAOwaNwG8/F4yhDVjwUBrYbWhC22Y8HpyJFqNhF4zGagOJqaI9bJFF9WmnfB
N6t/5lpoMbZGXghDlH0Nl7B3yC71LMz5dzCOOFfVfH1vM0kvIZh2J1ncVckomiVs
Yj6zNyPHoVtetzHhGC6OJVhKZm4WqJSAhsJt33CiPspbz/SADSPfrLUTpPOrTs1l
zQJtb1nwWFa0b5Ek3Wr/InuexJCWLBZiExCcYXFvrZbBoIMoKiW1benThpjQ38+U
t7A0KkG30wO+NNooA3x573gb/HsfyC4ja6govHhWvVqLhq9YRvZdIhsJV50vS1oQ
kVaQQ/KKHJW3ZgqjGlNTntCHm4GUd9hhV++gUc18QfylzrF7hNCNM8Ojx+BRr7Cv
cRsKH4RAqrs5BEyZ/kUpRB87LFY2aclzR16UyIsdCHajISfdByeFvjJBCNZJxd1y
YSRq8IVw8LqJD89+ZKEGwBXHmoDdDPS1uTpVbifYdshkcoJbbRfy+hcP4Z2XdwNG
tJ/G/x4sM8FmtngRGO29RaCTZAlMpHr1ZqWbQuQ7d/KOuXMMiEFPtVqniAek+f/4
SOtd1AqjpiEr06CSJZ8xBiCkqGuGEHqeL72LeVRHIsb6EBF3Ff4RX6/A3ai11m1v
X9YBD11mddZGCizNSj9SMI3kqS3XleTSjDZnw+tEvQlfH4AAbdDluZdFkGVAkawG
QMyl2bioAWlylBDf6XiFU+mqEoJQaWNaMUKgK4uFXxlLuWyGhnIedCvcjzoD7Pq4
h4G32kxoddEVls3g7cgHNhC65goeJja4ydxZ0+BuU2p8rfk6irkgi0GfjXdHYmlM
oqNtUAMWr7l6gjHaYWJ+K2EMPPdxtgFS7kbVmi8/51kW7Bn1dv4DUP+jehNRbwl9
ZygK82dCWcG3gROEqCfGY5lAqietgwxJswctDOfGk4KB9J3YvfgnFfsl3A7dlYsw
ZH7PbjvRe7ANjDZzqi6557pSX4+ubFE4bBPKmEx94X7AXQo1ZPOXf+AGWg4xAFwP
7I1Aa4jfoHSM4HdvPZ4eBbzAoJLeffjXQiuYgarLiuPHcupDuvH6uFj24UHtZKXM
Bg0Xhjnn1BR7fnQ1aCfFAeSZqBdebpm0FzvDXSnnoqgV+vROiGmIbijjIHf894GS
MyZxjM1dyo5ATpFIh9VK23rvRe01qwp9i8/BGeVYLJZlWWe8JuNwx2xuxlNjLqU9
9sfcQMRUAmfUQVYAA+Yt38HA2h7pR8kR4trJRjCC1GLm0/1SBrRVbbuO4JxOTYA6
dlBUx+98v1x3f7IPCY51tMYHhKQpAEP2Fbbxlxc7NQBCo4mSpKoKFL3w8FpIr20c
o4AlVEPCwRxZFruWNTo36N3QCEgbtbmHq3tUN79X8EWcnlL0po9dPufqupP9oMws
W9/PhYkKdXV3s9c8uq2BTzC1HpfWECcmG7ap5vMIX8invzEg61qUWy5kmvm2JRbW
8Jyp0UXu+z3gISkaV5TJKFajuvk1kl1d8H1IWRaRHuNRGom2TajnffVwnaQ3Gcg0
z3rGGAxaIYiHOqeqVdneS5V37ynljsTR6cH0U6bRj7mkbSi6CvWZ0Qzre+nEFTC0
F/ww4LP8SmmPZvMaLEA1AOTDTpTXrWJHEFB/4/wU6X7Q/8nyUxJi5YeHaCQ7SJIX
1Wl3CTzm480+6btIfrN5p/mEDqM3YtwhdRDUONw1MmmR5JFn6AACoA4xJ1IMZl+v
wn0credmqfu0VU0a3S47loAh5IFpzKYEGe82LquhgVTBOLA1591v0wjqt81zeJqY
OE72hCARfGCVw9wTvU6D0lF9NQMgnTEvbT43aeGmQj8z8CWYcOtZ05/3nSvLviTE
A2v7YQqhvrnFSM9AE65n1sQOcIEMVVia0acN6DVlY63f5aidOSndsiO+HUem5q/K
hcUFn7xaNhrwYMO3hTfrMuqYPd4Q7lHAa50/cIseH7pMdBoOH0qjFJAMEaCqYjPR
3Gku7mF45GiqbFJyi7aglD8j0L9KdTICspRL7zOQ7SirfWV3wINwsPq1YT7AwDmr
CAd38H9stgJkApBbX7I2my0H9DUxcN1Yb1ga0ti/c3NxF6WZkOlqznr5jiVMQ0n5
CdpcN7FZ4W2Jt9oX+OeojugGQ3e5bBhXPb1Xrp82VxVxfjTZU5t3yvjRrujeGCdw
leqo+ZpFOjpJRodU2dCnSCpxCFoeWweYZ3PnLbr1ZzPzD6E/ObfbiKmfuckpHQZc
EDDrfZo8wog9CY/lefoY+9EgG9Y2sEjThXVt+hg5/dKXhYqvVbauZwXVOQrggDqF
k42RMQ23BEuz/SLyWBZ6N0QYHFPobTluW1XA8SpUVS+jWEn/2JPtnTetYetrk6Af
AfYRNCsDT0S9HlD4DBqudfArBUn9RHkPyyUyDf8wmX1D6bg/uXJFcpEqz/SsXqiT
vecxFMCGAqwS8aA/q76QgSbIV2/fI2oHE+uToTq+d2xvLXQ3n/oVT1kcYYiOSXM+
R4BrS2UW4GDlUTvCaeCbljmuCRARHWXYDc0X85lH5HPIGBTdDsmJGU9lOGV0pVMw
gWSaHwvOTG1lQQ0qmV/9EMEe1zl41zsiAObfQma04JGH4JENN0xCNbjg6d1HI9ie
xWP2rQYm3/v5jkUlqSlJtamvGNjLQBYe3JbYw5yhotLT+naiR5exMQTAOhSGye48
p74za8Y9T+kfGB6hAXO7o/ustZsGR7mLxhoxJTnIytx4mnIgBwuS5+4aaDUudrEi
cLRvlR0wZSbLPO1AtgB2X2UCTTN9BiAEodVEYwetCw2BAmJ1PFoN7hTiabehBTfS
A4vo40cCe99Wh+ZCL+MUImsNeky5jdZCMkGX3V7wr53ImTGfV34cXaRDsPv/pIWg
JGLJQuiPFgO/nWpvNRGsvDoleD38UcUJbY/I5wGo5T9tlzEN5qNF7BleskCSIhGl
dZWcqlLX5hLFqAqvewKbhvwK3MkKHXhhd+7GmTIFp/VSi5KaeLixMHayCJlXKGRJ
x5T2MbhpDkLk37KB5m++ipq6ube35pjIa7jb9yp+O2VbC7vcscuclg4FWWc7aOw2
Wza3jiLSGw9Y0gIOjkBa6/GRx3fxAyd/N/gBsdVWdT3NOkLFbWNpUdIlkitwKF1h
J7DvXqNQfNDXyzENNudHbAFB2NVflBL8W0jRf3950g4Y/WmeEA4BG9dldt9EmZV7
blGjUY7DuB1wJBfFfzy6HB40mjHsc2InAPyPLKupGSIVtsXIleSE9i1IHewEjmHU
b9jAk0jLdWaOxyUFlhuNAlrVCPrnJ34UKKl49jbVgcx9K4YEE/Q41ZA2qUMxn/mU
NyqPkkuFSqASDVJaASmyeiXjskEeCggTSMpwdg/JZFhcvYNL+eZXVwM662MkE3QA
PNine/37AoXEOQWZT8lzOckL8vYxnNwTQBYKwVPcB7P6JeXHgiNEEk1ZDF99KnXJ
MSsPR+UXr715qwmpgYS/xi/WUobLhaIO5XennYVo/gksUJ4WtDN+PdcKndeMlsSR
LAO+Jxfio6xyH7hFrfc6XVWrd/KS3FlecON1i9WMYIxjVQh//HcW/DTQzm+RqLVs
8FZHvP9lScl4jATBN+YUHiANo7/zCDDzC6fPE50z3cq02OxsifTCqFQbesL5g+99
yjjmF4L95sMa9rLyKcU4ARJxQdsTzDOQwkcYe28mYjawDQP7wEYWI75oJnDVuq8c
yEgmfhCBpYIPy0NR/5mdWNSLI/f60pCDELFDWt14znWp8bjmOZqGJ+VKil2xkh8K
Rircx1m3v9G35mSGE8q95hGVNBekNh+p8/FdB8BoikeqR3cpA72/b8+iFwdNfBlb
IlKbYupI+6BKJ9zE7nULYjGcjLAHOcyzmnVbnJlqr/WoitfS3GcatdBrE7CjiUrb
OugkgTunSWvz0dVEdy9gvm/SpTrzx/JBfgLVcO+X9JouSU3rTlALiqde4zxA8WUk
Hu83uHfSqcDqhBdsragWAaxPvgup771RqZcj5nntcfjvnVtpXfGh2pdsbPSSyLab
qfkgO8PTx/g0Ae5OyEuEX8zcGOMTykopmaW9/N/qz4H5zR0/sA/o22FdIkj3xz2Y
h7vYPknm1VcCPEsfZ9jHAGdwAd6BaomGbYADr0oy02Up+NmWP0C2AglDmEbIgIyF
2PBRvyE/pGsAgeKxbHlAFyN5WBb2YGUi7upVVuTLR05pRTC/EGYGvw8Fl7S2matr
Cej6TLL4APCx//hVyA3kOGXgHGUJoZUapTO+07h/4W6ZJGwlWByErj/+NOSLKcL9
JZ9MhTg3JSbV42Z6r0H/BccUkSB8DhvSPfFeG/shEZJ7QteF+BaXagO1GWYd/gCR
WoczuAHIwQmUtSE4CWuht0pKH7X6IHGcc/jrQRiTlfETOkGzSa3qqT+h5NPTNXWI
zIt/fbyc4gnWWIxawgcUHJbwSYXQMkaX/FKZKApOYQ3dr16wj2B5oBdEBE2PYEXp
9oBwn3QCyJsGDp7B92YbKnLz4tciT+oFV+vrpWZOCbiIeBUHEvFHojXWDwFXCvru
PSHL/Bj++PTdVfGP9aSWFP45rlfSZ42T5DVYZyOQio0yduffMXu8sFZLxSCQZM93
liB5hTsyIT9EfcEKUpMX9MXyU2z35wH2rwkGcHzzlAnKUOwV6IwsP93Gi1b8zef1
5BAnl6jJCnKjf+DEcBd1Vdx1MU7PkGnGe2oOG0M+I1lz3tJjWk0yZjMR91298i7u
1PP/0EMrSXMIvcctYQjD1jH0NS6BOnTuueKMXFYLrOd5s54cLj2H4CiPkjlzq5/n
pgmmEGQVsS4Os6yxPdg2Ugw/NrjhKoYfBwyDsr+TGPLeDTl/uD4dYhRFVoBJ69Iv
W1vItODK1eaN7q2xiTMvPtaG/gkvFWcP3b8UZIs9zAozxl9VT5q2K+L7DCzcfAnw
t75xV1RywWIQcG04+HJpv8LjydCSjcWewXTRpyDeJAXdz5v4YjLg3uSVWbEtpIKM
0ZiESjjgZUPj+Ii5fOljB81jKuiHVvAjhkefW+oBSynR76xvpaSjxHC/D01okeT8
IzsOYxWnwi+aRWpL+hgZJsBD1+dExNbZAts6LlWtdsubivPaZb0QRS3aesgYz0S+
hRc6lLsD/Pm7azJ84UVPSBeBNXYLOaF1iBAB2OPlra8sCcftOgejYDoo2BVbPZ0W
qFZqVs4HrkyOt5zSZ1SEWEC+TES6PitIXYNx1r4fIC0oqlPIJiu4A7LoPjtqA+B4
7ia6e0a07UbZWqEoQsgH2vxDiEwM1jtnJ5vCj5lFDA6ewS80NRPVilyi8av+vzB+
cw2mTpeW2l3rTBdh/OQcsRsPDaS40TvmIZsbfTYgqsERO3on1oixRExtoMxIdo/a
1q1YcRyuNWSPUw2+aOHhVSWdF2j4kH2DZdIn9aMuB8bVtsIwH4rq7xTmfu030W0w
Uj36+h0n7+VhReqoiOh0/cf9m80hvluYGGN4DXJXYI9DLJ+kVonThVKhbi5BNJO2
X+if7k01N6yxqB4JZqUrHgmLWQJdZ5g4Qi8tbNvPjDEVuXb7BWdG4tPOkD2u5dXD
kr5ZvQ+Nqkyksc4lwwjSBPqRTD9qmTAnNnMUubx1lPlTthx9B19h/F3dBfa1fw8V
T0K2adAtlG7ICtbqU5YcNs32Kre2VBadEknNNMUNAJ8VVVpBbjtXwimlvoqI7j7j
DmJQ10ykXiyLWZHpTSJNTwSsniDmY3U7d9fiAUSMRxa2OH0WRP/zmQ7SjlijZYQ1
M9C+FOjHzdGBNz852dQCmarANahl1PMenuxo8CQggLCnXvHnnT0CP8LCNBKZPwtf
raeBeDRNegLaVEo568sRIYqLuoq77kJOCbcrlztmRH+ScQaceXJz9HVoAXF1Y7Zt
cgPnkKGSJvVtRqnXefPHGy5lMlp+Vw5m1moy9BbBLJt85jizFVuT/pZKRyPJ1nl5
YHEolNQCxF2zm3IXBUExZk+rD9+E/+m4ZzMvC75IyHGOZdeo7pGy7hYogGmrrx+w
/vQHD33FPmybM6RNvIfn6p5LdPKvf5cIbArNj/hlmjSHZe9SttYOt7G4N2FhcC3c
DwxOcp0/EDMktQZqyv+cNXv9CIi13Zt81GbAIZOwBEagjkpmhO0pxEKld3l9uDq6
33grafL0UxQ4E5xZMLo5/P89YC/JjTCVMuO444cdJDADQ3SeLrc9XNI2OGXr9WYB
pSoA4XglP5NFa3sGh+VhA5ei1zVGCXmkvEcBU4bco8LIouCtInrRqtSxtsoFiN5u
BWPUHx02gTDleoP65nhnFZ5mo3wAaKk0lFgnER/iIiXwMWMI+N0AZWvYCOZtW7TN
4XTj2VPpE77LdG0lKyw6o8LfacmaSbzvV6B95l6YcnWfnvIvnc65swVl3tJNH97x
+rtUbrBGT/5TjBSTr8MkvSpDPmDWNxex1VdLYBG3qINx4C6zjpRsgT+KZS+uVjBG
KI/vbWUbS/Gy0LcV7YUHrg0hsDH0gVZs7oY9NClH2jZjXIyYTX65b3UOywKzN782
2zIAghzQB0kprwZID09eyh9grvmISNABDqSnqJ0lyU1GjlgasNAja5ZqbAp3RGLi
0ldlc8lyn0hbqjRqY+RVQWWSrKbYP+jVcEp1Da21rxzcWB/Xq6TQ1IowQORdYHKv
bhTHf2f/RXRdAmQ4BRkVlU8j22/ORR/11GRPStqb5Plg0y+9AVRp19MilNi+wmQ1
VLXXNofdBfDSCBPIFFzAy5jQ+Ns/bq19g2TZ39QEq+W/83+bCnMwwAMrSc8Ex7QH
uiIuOjtjxkUT//zc0PY+OmcqOlapl97kwkqszoGyGbMBP1lOVJ0MHsha+WmKl/vW
cZfw9//8YLq/G9Tm39Uj/E3dayNvz8tMTQ5hV1a8ljXxVXGm6nVnKIGIWpgRlLdV
eNdDtSRhKPqrntaDoY4yywWPPw0zowsjZEjrvE4C4dsCLt589BOQluBKpg0KZ530
xv9ejWk0JjELywohenLC6qqVLCvbsL26EVpB3ucySOMJElCjCSG1v0jdSLf7TEFW
tUleiKE9/ZDzvGNi2nv5RkkSLPPwDt1xiBmC6+g8rR8LNfBA8xEMDoOb0dNAFX0Q
rsEMxKJf6lvC0LnJTq8tIN3JOfIO/F97yw1ZLuA0mrSxUbpxSbodeWiumAxQE2QF
lZlpPAcyXDbCuWiyOT3p6Mz2wbpIi1S3rR7qbcxa2xugUm7xHMFeW1RJKVFNO8XQ
a2Hf7EdrkQoI1I+IQtbMCCRbON3Pb09i9rLHY+iXstU+mpX9iUtjQbyMkwH7SulL
qCFcRvTj3hK0y/1rdxB2EORfpGPXuOu0E8q4+EWv8D9crNrtNb6oeBoxUQTStSXd
pJr1vsQgkVMoGCyMwY3s86YgdY3E0gL5Tqeg9Z3zEEe1TF0PDL6NEVJqrJQg81E5
87ceq8apPmyKhz4Xv3X6P8sr2vcPevhyRXovZap6hZbiCrlR/vp/KhnxHqFeh5As
HF+KNtZaT4hzIx/X19cosXP5vxDNhCc3czpwGeh8Sc99p4ZiTaVk1wM97o5dZfcW
alWF6J36Q70LMd6Dba/SZ8gl37R6XSUyGSvemoh8p0S/LK4djk2+nR6ulwpI4OQZ
00Cafh0tudrXTknTk/yBFp38e4oTNdtXSeuYQVpZUe4XuOqOWu9eyKGpkJXqUtxW
Enx/Um2wxlClvWFGbonZYN2wg01t/ER0WTrrRjZ1DY/8bckKxcfJHHxsAlF6cHoB
sRUYC/6xg+fSCQgJoc8B7Y3SiZu9hGauQAQFh0eHj6ePXbs+c/1GJc4DFz3qBo+J
86l2DhN6aKsQN0KYpH7SKwjqKkwkXHf2veLlkPSvYZZQvyRp559qB5r835FsVUQ6
kgzeUwj2j/j403OAsrkkRoy7/jG1SwmVXKcsAv0FCUlJ0p4I61Nis7Hn/Zy4gFyF
K12nBK3a5HLtRdHlJG9Rl+NbCOmNfB16RXlbrnDi8ceDYV3HPSkt0Dz9nu0ineOh
5HhVV21hjQZYSZLdtZHaPKPgFZKy0K1JMpadUwx35RBlDcKR1zEgpYWsEkklcnMC
hYKaFAB7ysBoGplvGJpYP8wxNHhqW+FbEFoar0p1YdMXvMDDRyj6cEVDNGyb48vX
Bwm0AiAcN0j7Qg0ky69puLFSm+mNnBpHYLtvyKya2smYfdqFDfo7goAC45ApZoBX
6HdyL0/cuB8AtsJviLq4ULHcDx87PTu0BhzUVSAyKxwrk9eReqHX6sRJZO0BhgSN
bHHQ5MiFxNmEV2lKpEygCXlZm1U+NLhWc2pFFW96rRU9j8IEYbdrOZIaPSFIFQtE
1YjUEtSDnDr+/yBTC6rzuttomvPV6A7Aedh+fZjjysKU5DjUj6EgX2gep7JvgEzF
wy9hdQ6HyxGRCCCJt4LgKFc/XMYe5BE9CgNF937mn/5hXd+brMb9X8fR8+Z86GR3
ITs0HLRZ2FDfGlhPWu5ZBIkCCjOpsCblGlnCq4XnBENhlcF+UGLeMt5XdtzSWmxd
M4jH8ZQ2noUenF5SE3tTa9U/8mh8alHqlb0Pwzh5F+kx1WKgWmyjScfWzMLH6MB0
onMqWpdY1SaEGq94f0fme9JtigYp7tirKydU6+NCX4cnX3thiGnZCkXChIQ/OqH0
iNHQ+lgwUXGgngr+e1nyU//NyK6SrVxPeAhtQHF5/F9PwO1oB9nS3PO1nbmEONAU
qMR5uP3ufZ8ODka+hz9A4Ql+MuiWNVAhC64khphZ4bPp18rEcdwyPiCByms5RpKp
owRaaw+Yk0CgwveOzVen2Y0jL+w5tfVZfUKaKJayYFm6wuqnXj/RIwbXtwZuyY6a
h7JAVCYY4HwTjH6KZAromqGlfS+mHqVoIdEyC0BEyTVY2buLKik4DDLFhc4/4hgW
xDcwGJVTsNwphyBekK9oL8TlUZTfVCXn3vfEtun/wlrbED+1RoFkXUK9OYD7weNC
nCNBJbZRR0PxueCdfzPi6VRc3icjUXh3mgg8PLQQf574OnmTYS7A88VJqjmoxIul
u10aYWt8cuTEFHZ4K0ipf7l7uXAz9VX/QePtXrPZ20vbpLDXd3dXsA5yLrAYwmUY
0DgtCPpzP9oOgM6BMQ3hmT5SppMnTuPv2PoTcAlHa1KdfpGP+ZFZoXKEcB8bXK2k
2zJkD8bWJeqKh9+dXm3noQL6PBk25omeZ7w484lNsfh1hOdLpt0TqPxicSYsUP4v
1PFZCX59se3aOeh00+kvZI4fMOviSY28Tz/EZc6c8StayaqjM0Tqr/AzR4AkCmxk
HYM5h3QUCSovrq/DE5NsSffT4mApoV5NoFfRCgWAX8JDMDh47iLEQo/40pqYEZQr
q2dqu/9jFGEtuWyY8Zgmu+4Z0+TPPHPYE8eanr7QdksUpm1bD7UrZDrq5jD4lQYt
ny4G/f4pn+kVroDhMqoUvjHQ6ASs0QqPzBDHmfpat4CrmnpDDkLyRMCn7lSAUd2U
YVxSPQLrI8x+H1FpyV4FUNAIlFIcLyu3VgYuAq2GuvKghFVoaVzMvf059L22942A
xokROr1z6VHktuzDw6+cnaVYsclsx2zNpYI+FjSBsETU/bQVbYSNNEa9FxXDMBKn
37hxRZKwacB3iwtM7FdAGnZS1Pb1J5LAzoqFDfrOIcgeoFPQOb1YYLEVuYWBCEoI
qzjrsbmhe27manJkcnmH7XGtHdKq6poFKE18g6UTVleCMbTQu8LACthK2BbYbMO0
yEnFQ4XnIdcJl7R1zgSLU7Kxhp5Ao5ncNABEGaybYXftsqUzByqHISIZ+zCNzmjM
+HrMsZwoJOL1b78VvbxtpJN94JqNbsIVqdAvGzgqALUHLKGXNeTT7aYZ4+f7W0AG
M6Se6tHeFUGNhXbXO+B1gxa5RJW64Uok/ytpNnaNGJld7KqbHJc1O4K0rNcU92ST
p0c13fX4kzPddzd2uOWdhDDZdxzbV+snGQs7KNcEJAaFtKSn/m/Xj7eoqPlAWLEF
PnrvR93cxVvb5fHkCtCVF6c9ZaIOLGulSTGUKjwFxU3AlPnhinOPiP752kSu4BQK
HRBaAMChXdqqakWBSxXd8giOkRSV0oRWw7UuHlFBF+CNy8StI6JmU9K8AudUMW0C
KjJES12hLfde1UGFIaA6QUqjOgiR98skFCNA0uoATrWh/UBoR7GllIJpipNPgoLT
QIR0n4l3myDFy001VLQNiCQgrAIMbYmRpIiIaIqyZFhHRO5tCwvmEqFEw9ZdLisj
mgQZbqno7bF6Rcp4zA6vdHotwNDxHxvp6Jfakfqg2EaK/18Xw75DXFlWispYyw85
jAB6HJMrQjj+JSMV95MiCORmxJRGw/UxY9A7JZGp6iW/qOsxMVvEiNnvrbGDLYW+
UgHFAyw4RXmBxmIrr+1oownk8+4uNkl8JwMieT2KTcj2bHg/Frsb3po3ziYG5hyd
JSASpeSOFFYUYeleDO1iAsDNzhD96gUJKgD6GJ3wEcdDrL5QUPydaoJapIiSOWqA
AWw9VWEfkqVyqe+2g2D91x5Xoo/iKeVtuNAdxiAokePOz0mkKMbnpUm7FCN3n/2o
evboo9S/JSUUz1rZ7w3PnDQml2pMhCejrnhxTPqZwd5OIixFSDuoYG40hgsT4g0V
Uh+5g8+5fsHE6b3048/oKCT0ilFo6ySVTAaatarxKHLeOE3DKjyx+dFjWwSQIsum
t0nXF582JxP33YNG6aUCpSz1/GFnbtQaHSCDCqhncoqfltNScm0fanY6ZtpVaSyM
Sm2Qx6WTlaYetpICdI7iYXuJQ77szbvbGQOzsEHS2i33bbO+QwTytP2Y0z33YJOZ
h+sWOarONS+Cq/sSkF8GUzIUdltE+DJ9YAVof9s/rj8F3OPBnGGko1tK9GODjtyM
NgeAt0Uvnu9b1e7HjXrzdIn9AwWlAA54JWKa82TQupPsC+cQeW4XapRDkh6rn+kI
2nPwKZW3uA6DQv1V4cSUNcsTEt9zPrtGKcTezIAN5l4WL8U6/X1jAcuj3The3Vjo
TJ0TXcR+IfTHx60YfHJvxtE0nSHxq6JtvgLuFsgDCEE72vxdA8blJamvrsDDPb5t
pf91uwuQGqbNoc7wVLq+/GAfnocnR5EDfr8+fQNI3FOdaeFjwmkCZs3yUuTM4tlq
fmtsrqvi/QVa8DAW6SSHV46xRJzxu5ohNpMTlpZ3UG+hNjTATBpPuDfsGyZcHTfy
EoG5Jj+t5isbwWbSc+iLKIN/vhR0hchRm//NgBKQGcHxhk9EtdMlZIS8VU/xR/fj
VKJ6VmMhw4fcF5qZLEYLKtbk0rsRoNEzCnI3HJ4XS+TnfVCoaU1ynAFdXqlcD7Uz
M/EHqmaC5ucN9ttjpcaM0YAX9uRbYGjozIWGX6XXKadfS2TwbZ4/MNOzGapVeoWP
NMct1+2wLLeV9y9uDGDNzkArZUgi2hOWLzVgvW6DH2oSJuDL/R2yq/ukCeOHw+fm
MrOj38AotovlLipZHTr1S7ib46NFziGplV5FPw+4oVVNry1j8FbAXFF12MMjLpbq
kfCAJv2zkYOhqS6+rw1RhMzm4WU5LImlJcI4PpqhpKif2QOjGe21h9N12NULuqYH
d2mhDJAFTFRIb3PdkEtBeo636Vemj1bgtwhfFxYGWQhPsXQqJn9HSs7lMnBgxFof
3262ewCcz8zV2by2d0lTN3IDXvOF2WfYgVYH69vLbasABLI0De/YTejCP7vCKccD
TTfcGAPNIQGFvmXNav6ykm3WwGeOU3AAsfTYr7XcmOvuZXDV5wxnwr5wCyQzxZQR
eDsQstcGNrsWTB7Ip18mo1OnSK1U89k68GAOY3H38DdIF0GK8N6Hs9Dis9HHHd2H
VEBE80FwQfN5D1h0Ed3vnfsElNz0LkcYF+neE9ptsLMgyGnZP2113Q98R7+yX5ru
08Ah4m5fZelyczgx4uhMkkC2IAknh6LgPrhgaAKH8ODkLbmfO4zSK/wy4Eh+CpXW
v/SThmGR5qGyVKFP6Ih8oty41RBnPGWaavYf+D74p+/af/rBG4IStFQAwtUbkk8C
vhys5GPkMkxm1FMzsXTBlN/gwCxmVyNtgw2ri6FkP60GuTZf/tgPdN5FflsZC6Vf
S+LGYWnkSAhYq5SUdkLYYEBFVsZ9K8z7MQxwYCGZbm/2sMNoYuZK29hpnepQhFra
yhjptlob5cVIO5R+LhSs/jLM898XMXgMHmWIqp0q+wl0B415iWYKPhs/qfNJC6kB
/U6hpvhfshmuDcWA9u8xPZ0ddgAKxdIM5HW32cWSeZA6Tb2yaqWg+pdFzwacPtUr
kvcgQ5tGZv2PNBnqzYUuZSSMUJc+Iu0FEiAA2Knp3DGy5dlkauy8j6CgnLd05V53
7gfJrV0IG/V7yhiR8dbgPJ09rMBiToWio0kmNVAg2KmqYEwzVe96C13kDzNNQE8R
MHB442r7rxX3o9YFJwpx325AkrlD4KL6gIcDggBWOzL+pyLtfZNwwewU0IgpFohU
UOJ4QF1AsPZwB0DxG2AkJ6POtGEM101n22xfR0c33hSwCD61YElslT6+J1Ub8yE5
g1H6Zw/Y7uRrYOiSZS/oawAM4chyQwXFq2imsT9N4TSrJnOTdRoQg4fp2q2nVcmc
GGhVlkDqL7aprWppylJ00Kv2CTFw6WBy2Gv3yAj4ncjV/2n0CEBbqwxALaFVqTF5
WpBRCzEVeskR8gkRhWq9B6cN0oSq8iA2u7gb0A0zIt4btmj2yYKtgoMsR4AAttdG
ywBhIEXL0ESZTAO9AfTipzdtRI0axad3ylOSJKzTl9Mg3gkBiawGEA/rvcTYgViO
IE/0JnHQZdwR6yz3+8UcHeSDCAOALmZ86ScIwJiOBDQDIn41+/wpHxUhOfT+5fhk
RlorA9mMsveeGTOfaJf4T4UVxWbLicbfOjrvZtBpud+V4bwDlnV0dwsbXgJEW28y
xowJBCtNo9bN4dk3yEVQwdPk+w5aSXuCsqmrHycaH2LzWPeJxuVsFi74Y72RU5Qd
Q2El5LATd5Ix9IvTok5Wi45cfJOgSRiy5u0ag6RDLYj7VKxaHCmm/RR22rm4eEDH
sSSlxMJTklyb8neMecFzL+ECkdFb5rlse0HEHMhSO6mzWOjTacI7r7CdFmv6lm0f
f0ZYY14myJ9xKnjgTvLdUau7mPxK/xaiOP4gir6QNTxGtXeXHzgvat28BOvSF234
vBAW/2HO164EskIP7GK/oAe99JcuOV1jr/JrYbqGR02Kf7AwacbzdVhPOIdr3PcX
H2tp6Ey0lpe63TuEQUNNzaxzRmN7LHUEXmRPb2J0+mL22WUI9c4/V7jSI1kOETM7
pW8gEXQuIlQrHRo5IPUeB7fcaZwum1Lu1kzTCH23NZ/SxSO58PUivU/G1KSSgCPF
csW8x2h4OE1rBIoygN9jScGyajNOwBZDhx+WUHaWS4wP4jbax499hjx7Pl6w8SJC
jDGv4iYYvPZSC45jLGNsZADyQ9B9b+NpsamWmRHtzRQYbaQM0s2GK6ew9dOZ1hts
PnGHWDvhtaUDN602p4QoPbRj8fAVjD6hCYNPd7GiSh77ArRIeSob1I6kL9csAaep
LGXGnaiOqnCHlT06zYfE94IC+AMBWzbo4mozpRFKDljq6vMh3VAGFwgkbqU45kdE
lu40d9a0ntgvhRXXw7rXowbzsB5+n7zNbXChrjZpVDnc+0WaJOW8DN6ybIFqGkct
fTTBq1MWg60sdKN95yzgnwunK/YRRp1naRAxo9SnEUtBxJI4WUye38tqxT+F0zaF
N9p7aaVdAacA2cj7/mbg6cMj+8hugxMNoyN7v/UY2SAeMtD14Kj+eht3BSzjL6W9
igfyNaPvL/19BRh4sm0/SwNXgsewH+IOk1Nw8a4c93waEUBgtBoSOAsxoabOEcLg
JXJPmx/O0xXARzwhJD9o8DFtUlsuGSQc8lBQPq8Q/Bo0go23CPShjmk90ZU2DHDd
gkSpJVQAayUyicjaBexvE1mYdZ2xw1hz7f/+FhOYMue58s1IUgzdu/t3wMbWfYUO
aBN2mmgMeU5lG+4OK2i8ADcXAdQf8O62Hl43fk7oIaJ2MdZVDLTBXNo/C01BEDXh
JGZKNgYpkYPmsTLrr34fVeRzlHamefRWo9jHeJQj1TG60xbe/cAjnCiEDwbH38+4
N6o3ICMdLHhgxLW8J7jzOZl65DDoKypixR5Nc11z1c5+PTaW//ZCiZSn8bQJNugP
yjfVjVR4WZvQ4Cde8czjgtGG/IEhN5GminIFIwDL+4nkzb3ePCsU9s6EhmKwxjv9
3NeNN0SXR8Tp97qDeI/koNRlzP7GnxXwAZrYxm7NEJHDYrIutE0UsNik30o8uRpr
ViWWiITZxq4lhat+Chx3VMQnfIyKKKbfmpfrIu1LM0g98UmgoaP5BtVQUjf4fvKv
RY4AU081mm2Xg+2DryHKCsj/WoKX/wtuxwOBoxNhVil1OENpUB6iFk77Fu6s9A9s
fnPYuS8VeTsTcZtpockLi6xxP3LPuCyz7vSGAFtyfVIrLEAEFnlKOAS7WwUXg5m2
saGp7Hup0HUU7RqMdIhBcGOwf+bzg2R+Oeb0RB1XzUSqFGPm807uwnZ+rN1gLp46
PlZhh/nVihVLhSNKU1V9lVHqBVqyYDsGF2FcfbU8tr3UdLUv7FWFBOw31ZBk1H2e
7I1VckUp7RGogT39Acw5m32szKOzEquZiKqqUUlHeUg7u22zSTgyHx3WqTiOqXKt
hc3O5SCYhb0KkNonMRJpGhfkZb6e43QYtuc0KxwFVY5zM+siZM7N512oMbL/kR/p
HtjM5yyTGywofCw+E4ChM4S63OGbRVBXeOJAsktExfKYBPh/GulrbsrHFlCvLAIs
OmZNiaOvCS3Ky5yVC2IQZNB2dfDi6whzzDarRNWANNopjTuJIHiBa/U/FRDMlgYD
M1oY5bCYQgdM+ceJ65c89/k32fE3l6YxkvIFRqqK3jGR0G/tkMDM6IefrCm19+8K
Fy5INhmQqcqOmUr8NAGUSSLyaQU5wVK7qoEzi3eIOpnMue/bITvBrESCY4qwth9r
12/4gSHS5yBCIKgiGSGuXgBVJ+D2vH4xWV+OrWoSqKdg9OkK8d0o2zu6g1qPOFQe
YOfvlrabxd4DXj1cPJl8nWTHQJl9X+dnGBJCpjCr7dBRrsAJdhR868/CMjntWuyC
+ni6sGvYiC8DX1Rnm59p4FyIiqyXc0WzvLr50mNnAQSU1xHmjCRjQ62RTPA0J2lV
AtA7wjildnEjUZUrAowd9GoE89jzoAcNLW5NWh1b501k6r40aZTnD8wzXKRRHJlE
LLZt3ey51iY3KUYQ74h1TWqiKUvt6CVkhjWlui+frwQ6IxQMpUtt39YzsRK9l9jf
dCPSzt8VWrqJTmFmvD01T7FMpMXDCvIc8Dasfkt+CeCVxNNhtEtV5RXdKWNm92HV
vdZt8ROxL3OB5bZ6Rf5V2/fSzFYfUzL74hc1NYbjivHd26YkDe+SQBFPgAK/EVeC
n5MNBfmNZgojkCjFIjHdQw45r7ni/21pvz+ajBWsG9CJ51gR/s/LYkyTrsVg/nUd
qDWZabZZEv2XeIunf4dPDoqE6wPrGNHoyBGzrbeXKvHh4OookO7y3rl71J3WndTq
zAB2uXQBfMPQpaKWfgXtr81yUlpsufEMvU/0LOo7Y09a1eTJTV25cSJxjs58aEv9
tUaNzMHBLB8tBwJYNjKdQqYF4pvcvZgg0NNlEt6+OmEQF7q3DMNbCgjEKIrmkA++
ngdMYd2Eao0409KdVtygoh8MbnkyqgEcVLBhmd6jutpDVb6I3/d+g+W7AWY9VI2K
GavGgdqAeGjntL0JD0DKzu6MYJuKP/SSssRXlUAl5aaHkKyqczpQQJ/PXf0FRlwZ
JsjKDaWKqfRz4DaoVSI929o7jhy3/pb8pkWWByCiY9whXbac2Wo6mHc7GxrlwS1j
ofhNM++j/XmejM3e4Dt2i0bjcJe5O05XbV4zNEoG9dsW2yq7DiOklprr+JXSotQa
pc63e3dxbONoGQzkjL9IqyOYSainRpPXlXCgg91+u5KEPqs2Z7Qs+x/X942ZesvY
u5Fj/vhAFoG+YvWxg15oPN8BZr3PixeQyuje8X7LDMMGKcGn9Kmh8LE5EiVKPIl7
sPzcRG5Ri3jsYSEBFcIM7AELE5cABoUrbEx7JjVofVZ8LB8CRfnVUrKB4fC77S46
Il0PtYz1rEs7MDzhWzxD0JHBi6B65XRF5PAgO4sniKsN+sDVwvV+4Ywk4bN/WeOa
ylPhYw6paPEwkBrFD9+AnclvAHIiJX0a8AV+SQuAFWJpql4idikf5SEhJaQB1EJ0
N8pVydx7clglMnKGW9U/on+bVQhxBewpcYK5m8Yicu7hfGad6aAklJbZMGQ839dh
HrPJbSPwnG403TIsg6JpG/af7QJGqMdIa+j3ny1vHeK6lVMoLudHnF6dH6QliXc6
vDvKpCauD7KJf59y56rrejZ0kK2UuRdYVg2m6oo+f7mGwBslf0usaM5SzEbDxzTS
fKfGovWf88yv9JkMme54r9T0XcOH4sqD2IaWS4J69kAlYq0liWMgh8VN5aXMkVNv
o/IkJ2TPmH2+TluYQf1/XTfgHP0n7YiKzLI5LwWXwN5dlfvBXjnosVwlruWoJ2ZR
DDmbEKJ4VEkuJYsi9a7o9HYPijrzquWiFKtrLNQWlKUiGWAGUWoRenEs46hj07rA
+DhkjNSIQ1UMtdAjeIRkCrjmzyaSxqTgsD46U7f68AXRDlPn8/6ahP6U0E6PsMFN
xzasPxe856EH4MKm5VoHuPISVAosyYBKtJou+Ypy/y/e3J+CaHsQcO1IbcXxmBZZ
QpwItL/ARwUyqq1FQEx1D7UIhbKC7Ld33CWX1ACPqW1DwgoqIwbHnzBkUGaz1BzI
3wSLYu4AOsZgD6/dPk8AJRn83KHUXtELlgsmCOLR3dhfPizoQ7YKncsvMNXMmfT6
0PNsoYwS/ztq20Chlttd9dnM98ES3gR1JQ+m6YECy3FFvM5HWRkIHGxCy/5pRD7F
16K42CZopljEEJEwMHniHjau5TwmzWE/5+TcIQKCy68RNhr9Ee7ZAqC8Yw2j12Ox
PvtAabgGQU8qLPUy9qTxN2oM6j8ZYvt9D20EWvxLks+gw1fon209TAh6O6WYVgBf
hIFQgdozB2BbnheRcMBN2of915Rk8SXkpSFSBHHBhX5s3DndBlZNPZxjqzm+d9rj
Uyv38j7KAnQrn/gS9vtb9ycnb347kX/RpM1gj/nOKwC6ciZeqkJ7zemNujbvhoII
SLkWB+dKuWArvo+TqoKKCQMNdggmeMNh+Nu/dat96QNg1HGNecQ/AldMqsdNKSGI
yjQlDMhIKhaaEW73UTpCtdxn1laOipHlutH4LxTpWP6xbZPBiB/iX/XyaV+GSfxR
eol6pRkYg9ZK06gw+okYkHN3UugPEXDqee07Ag3LYZUIDLHNKSgeomKW/Z4mAamY
mjepPRiNBOvXRuPCgsFKCnt6md2zj/3iKbSaFElbfOH1mR8zbQlBeqzUTCjjUmXr
Pc2wsOQ1zsVRyYZJFRw5c0Jgig0+V7SzFHBu90Ogu6jlwZwvvM6Zf6kMb4pL1rtQ
ZMLsAb69/x9Rz3pnwGHGYBnETBTzw8q/fljy3rnkiL1TADFQieukqy8K6l/CxBvY
fIZQh/5spRj4/U5eU1KoowLVrRrOmfSNmlneiioImIUOrMMf9xM7YB8+vRdtEExD
QBApGbVw/OaTMBUWS242BAfpppmSm42OPU25Iv13Zwk+53fHSX1PLQ8sNP//KQyr
0tZ/YGdIXfV+0OdytbdNb1l5XOSEGWHatsUCb0ZYNyGzrmPCaWnZVU4oGs1QEi6y
dUfO46vDyIz1tbl+biJynyBgBC19C3Mnykp0edfEJFhWNh8OVtXZwGdfqvfbFSLj
O1+SQjKN1bSIIQPA2m0Xs+DOGhzLmFsbDDOqhqk0CuU9Uu0kvCNQE4sTjqGCsb5s
bub3V7B7HsJ57yDrE2T+uvWGcGbitA+VFDulC068GegdqwogxekAIm/Qedrr+ibc
sDjEAPDzwZizux6yce94570QnvhLm82BoVIeIJ1gpUWsIm0wsZ/SBB1k9MgAwnVM
Vmd2wTXD61b8gsZbnbPdHetUJCkoaT+69ppy363u6NG2igWKRkU7ocLmixFaZ2j+
kzWqSttv8EWGoWYVguN8UCc4+koYhherRq585LMXYdBM5hySxSkXglObiX3VLKbr
max6yAkCxXdfokHd56FDgK+guO5iSqPVaOK8B9e5kepLa7ebFL+RD7n/gnvrbxxM
2d8DcQ8p7yidJffJwHHwsWkxQvD7JLbgNrnzMAyXOIsnCt1ZufeQf2HuldXFAMEm
mWxNu1JovH6L8dcLohCsNIN7k8i1NJV2xe/WoQ5+FSToSqXJwbGhM2ifGKwDMGM/
tGAxBzWbnzdTkMbN0hkLOt02DcAjPbo8UD3UgTSgwov1QjWqXsLExXURknxUa4jx
tdEZ5a4Rd78IM7PK4vNnhLBUMS8Podiv5dQF3nrazBsnyH/lAAwDYkHPINRuSabZ
jqVSkJGTex75UfcHy2aSWHknhv09xIuuHlpJAdf+HgSbafdtvwtWhwC3RGpOkheZ
w/cs7lrXDuMrMTAJYdFapVDgZAjbES/ccaLvY6uddRuBRBpBwO1dhbDpZQaTiMTa
ntNLW/Tz+d1N2mIfqOjmzQewPCLhe9NcrVu/7FESW+CKeNYIqYppK+H9Up8y88pM
3ZeSfA7f0548X0ng3StYth0/9RZlhWWXp3T7sUm4Hk2EMxz0gPb2lA8jg5oK/Dpz
jRmh6WqFJTuJoDsbQ67GVYY+0iv4fh5izDJ+baxwdvsweBWnQm75C0tRLKaQParf
a0uczFJgLcoCG0jKgfjvAdRUAzttFv8//Sjdn9g/1PYgOBdmDXv84jRm18rnrNyU
RXR0gyftcnChkl/rgSo9qi6skvErBjrdi2Bw5fZAIE9hriV2n3Ma8liI3GwmsXX0
u/Bqlz60/t5F5A8s6ab7X7XAa/tgdNp18lr4xmO3azNS+3Rvr8jHtR5nxaGPdwCg
csUJOykGkvcK7RA2jAcV4D8N60Wb3kE8C+RYVeMLJMB7YgSpBGD8JTTIFGwCLalQ
CrDjaUlGac4sUdcyhwmZjZGvEMQWw5dGmTPa1/F9x9NmslERRVWtdRKdItmRaozy
Ta9QGAifKQDkSvDsTHmuY8slJE2kj4eJH+yrvg0MIMoH2z5+epkuf+7YJfR1muBM
iaX1pasHwuGx0OyZjf1t/Gv6JPs3P6QKTHrg7c0K2nTrLMkFw6vOM43FKJT54sYe
BMm5jDG614nGAeQdgu3pxoi7bq4g8xqN96dr25fzV/oYnn+uppQzhBOShYoRWpEf
TjOQMbFEZ+E1lOp96nckP9gxDFaebeyX/uU0YFvQzVGTzALW3/hJxjUIHw+1f81y
Qg0zEnMAbS+U1hxWSH8ZaNZlgz6f3SzJKLT/DHBmuXa8CG4BIgO/RDEqq4OYT5Cd
8QJBriuJF6gk1IcstH4S8zta35BbpGZU7nhG+/T72gFuiwYhM0O5MeN5QrYdxcKR
YZIrV944sb94cVSkIFatVZmX0DNWxUJDFRti5zS0EnZsOJGiGC0d2UInQjQzvRFy
VIJ/OPaDxFqo7mhxAA7XxhvLAfkloeGOhXiIQS/OlDAWDrR0X880mgIpsPdB5m9F
lj7VwIfszl/lGqJuN9KlN7S0rXlvbKotQOk9DIm0zt7Muf5taNe/GcWv82GcmYFr
4OhXEbTn8lqaC6k7RIxIq4JLz3RY+7IZNQkzhgOD4SYJbSulOdgvqfR+gZf1UGuB
8C+UTDGxqf0EhIDDZZvGWvUbn4R3xz4e8p66ZGbRyuX7jiukvHisTKPu0VV7nEy6
8aIvrspsWhs5MdVUTA1c6muufyUiqqovi2sn9ou9U3/9uFVKf5XLCDCwPbBTP21f
9oabz1EtwRFIBc34oiuzt9LJiVdglNxOe02M1twiwRZukTBVnwcRGzSQLmsDQ6SB
ssFHtx+SuOM2j7SlJUKTur3/fF/hWGzGpoIpjVNpe0jbbTKFH2HxNhFDLX2V940M
PptWHTD7Li7N4nFbZKMwslN87G0mhStnrZwM4UFnEzL9Yrvx3fjAah+RhpjGtg2T
iXyMyBhCC7H2kXO1B0u5/4Vuzj7NxLokFe12nTHoZmgRvpvlO9Ik/ZNLmmMBTSGh
KeDFg7TsoiRl8N5Ee7647ptUVO0QfJ7D4tJW2/It78ocSO168ubOiJTHWtgLAIil
2cS1biWOcxZTEgwivYVYGSaupCRjX0IvhN1NpLYAhZLnOHwXxiPbhTckVFXn5bCc
0Q27hjHWHUg+z2h637J0Udc02kwWBdH14Ngz+OMLsK0fozuiqqA1t3aYz267LRZm
bEf90CNCth03zPjOE8sna4ZgHwURiD+blwQ3VGNu+q14A5xuEoMuDsEvGUxkLKcv
O3gIsbFUFF5SHyN5owjc8obiebrLmn96rWLEAuRvIPCuIga7AOuQKrUom91SDNo7
VVBETV+yF1VtW4g4Ugm07oAEHnsx6SG2nv/QvCVIgzU1/JXJIqk/jyUr0GDHzFcX
LJ3ayESTfICgX7nBZ2nRHrTuGKaIvorRt+S7yvFQKl8UVHmOUo++nPj0XNd9ZYUG
pC+/Kf4rAswUFrjWlSEPR4pXR79DiRHqbM2N6ADRAfbWhBBvq4fXAyzUHx3VXteX
ZR8rh5JB/jg/YWvXqy9c4J0rVw4aaonTV0sNl7IkTB7uZTlZ5U7TJjUhW1aMLhYX
G3J64w1/Krnjv9MjFRraUwQUskvhVVDHLepUs6S9zYkK2I+WPnw3TIcqrs+ZpuXH
M8XnPRXZwZGw1oUKHzSOCILShYD+a0oLZb1BPAmLtg4M2jbAo9my20R4YhYmLOol
RWXDZrBixwahUqnHpTayd2uuksLvhsV5cDm6lspaczt4KyfGuIP4fbFcNGHl4MlC
n80kW9wtMVzOPZxxnx/oHUTOnJeLZo9V94lt5jPNQgjWktRfs50SH1YyDtmniFhU
/mmHyk/aGq8VU9GgtEE05zxfBvPEq6yJT71w9NgQsnsONFTbYcRdBetMPfALOgw/
L76PpZMSuhKjqtwGBdA5iXzzCq6NkJc31LcrKceSJxuaMfI84dTmn5UeRYPcJbZx
96G42whf3dD/myrdVZRlWmUBwWW41896NjaxI3IBAAYJ/437O4tK5ttNdvJdsaEj
b2euug/11C3+QbkKGJBwXozohA7RXGhWVwhQpp9r7aqrD+8/hnb+PUgyGA36eHYT
vpi9qsx/zQLVegb/Qz6MyxVWwtBQkkb+SC6ZhS3F1jvnBhn1vsVAmId6ckVSsKTv
RysGItP/4TsRAhnuFW88MFmAAf88hQH8PkCqn3LzBGl0aLPixblOh4erzxJ9X18c
8r8Hrh5S6wfqTfuhNUWG1SrFFS+OV05DGDNWTiFUvEu9g1FNcTBNNtH3dLmgTqm6
l+Pcvftkbrh6XfV1iR3EoYQ+8SD5HzPjO8CYhTd0XK3dWKT5P1pb74kp3x4bjDPt
chgF22UrRU2n+bWW0J+DoteeHfgqFHSSlxyyxBGbVRSxFpaPnh9Qha8+Vml9i9YU
RvudsLPLKSNbUojxSMD8V8CZREsJr1iffaRnfnDNTpCYxjCyNU9WGN3Vh0mTAh8G
VrpWl/r6AR226LpAJS/4TZ8PpfORCOTSHy3wjcRkETaHcEtMEK5Jn1O3VmfrUeb9
Metk/hr5C2OlojFc9GQlSib177mbViMoIT65Eqg/M5e3tcN1rywYG5ntw3SaxDdy
smGXVRC8PhQ/40qg6qxKWkhJlIhZY2zHKzwfIz9VldLrkQmWoYRXKJgK4CFjVzu3
YCojhzAAoE7UJhGhxxZS+z/1saQTMhZ/UbbTQZ10bUM4gsnsiVz+rGTuWW6b4aEe
F2moYGsK2HRo5VlyjqRRULg+CiR31uhpU6Ri5s8q3AwMOl70XHMATXb0H4yRzXHV
GwlHRmYz9fSiIFxuTOJ82vgZ6wc8UUJc4SP0yIxgpZIbNl7dP2WVFh9OWGiqZUuv
/7es3R6cmdJ0teN3uqDzNidrag9nyU18qI/sHNZBHOshQ++4/ttIVRi16z3DmAIY
AafrrjFO6+Q7h25LWXSkdBDV1ujjeXY4p8vm5XsSNixZpMFfx2YwFqeUdO0O6vmd
2Y2jb81S+6034MOhZZH/ggsKSkWbosJmCoScg0CkPFuzh+g2WOz4aIbgLRCJQOiB
D40aQrXCq/cDg8LpGfpqWsO/aG5voKmqpHnv3VRPt640oUJVTCMFRvY/MwqWh2ik
MigFnWBN5Lu1b6dS9euxILVKJnLdnuBiYsS+dy+A3GUKBIL86lhDuw8ZuX5DxSWc
sXcTYlPkfmmimdrrn6KSzjQB8YK87YQGKORjTL5CpCBEboDIHTYBZPQa43m3hUMJ
gzxNv08Ru6J0Ox24QiBHAw5YucYu+JTBocAzP5/otAYWGqYzzMo/A+icRP+9oMRc
aLAbfQ/tpP4+iz5E/GaTnsyj3a7s+8w1GGH6pQM+uZKBQ8rFb+b1juqW9gR1UemU
ygzfml2CZGGMbpYxLjkNxpYUMPpxucCpt2C4oZ3LebsemZBknX2FJ8IEq3Vbjxy5
wWrNs33tMceJKcfWltAo49PP1HQ4fEaZC33rJCwbho5VTQA1wks3Gvwic5g3pW5G
4KxYEkaKk45D/Ks48yOOl7RUNI5TVwzgFnC2FieMlptfXbWSSh09DVbJBlnUYljr
sbHIr0eDEziWBXa+ar6HRfe7UerUH0bt1U+BCED3eZTqmAHEZLAXIadXWJNUq7xP
SEWHvjVJetnKZRh8zjx02H0UYG04D69ZWWRK746Yt1iS+Yq53S2uLmUmlKjWg+DX
kjhsYVGlU6qCZNE3D01WGHztQyCOQ7uydknuGlTixHpLnjamGI9APsPz5yQOhu/5
cHWmmH2+UVsLHN848//n5/8De57J8MggiCEIcqNctaIEpfDWaWrFly9dXkdTwJdp
/s3b3o6CYyAcCnebtL7ULPrg66rI/pNAdwYkCZNtlwallTc+5NkV83srLS20YkjV
JAZ435YJX0YiPXA4YngACbXYKbgNOtm3xLDnPQA2h9HXUWCQbQo3DQFwImSrhAvN
fdv3PI3+etsBcLAN3c0FBPuRSuOQNoSk7YdGRT4kd6KLNV0vvekrf5UmJvHEYtBi
K1FoP8RnB4tYlopE0956zOh46++R7OFfqbACYoOaUMiyobz0kU+ttE4o9V6Gefqh
I8QgD34ddymd9dkXyjlZT+lke3sSm1ahvYcPx72jWdvcBnFg4X0XoGMCvelDB9CU
715mnELYwoF0KZCyLhI6tXNw9pYSMXwuEWTwtoMJjpZ0Vn95oFm6Virh3L38EIkD
Y1dfhqYbl2WTpd4XuqHxC2OYv8IoJMl7yGcG7AJB9ySiJpIysSQK2dNSILGwSkUN
Pi4zKJZufEN3jO7A0IZW7sC6vSJd44/O6gKAWWPN2GnEpoqhwg708yRulHErT8H2
wGhU/zipu0DGhrFqe66kmabF/Fg1f1u+h9m5g5sP2DQ44PzNdVeWY4YBBENh1Ew1
DAYXJZzJry1ICLd9NrzQL2ueE3cp9chg/JnH4shQCG1tiHOTR9ShIXIW8YhaEc39
82oic7b4TnGS6x+fZn1SkHsrWRlvVIJ8Wcbd04x6ZdNuKdclJlCpyWfYOZOsxfFR
fU27dvDTJV0Rm7CzPpPdgiom6oofOQDlCuQJ6GCl//M5ftSjzh282AfNEARrEa5y
rodNI/fPtXNMcWgHucUsfXPyClolFtTzYxaJzS99Z1YnnsaU627r2o9pUb7Z7nmy
6FU/2qyrcZrtC2MuFUK2P6PFbN7oVhVz/DuZW5avXGfxqsTtTu35d4wkCJsyzY6X
pEeLuJs9ytKTehivU3Wz5iJTI5ngcwdylyNcGy1KbDJ9Tnbk+D51l+kWeKRmKy1B
2GaOwSq/lUneWWiVz7qX/f3z5iP718CMQCQOGf1zmn6S14/THYkKT6mv23U50fZv
n40s6mjd/XWpAkUOiKWmn0l/4x9lYxrvrJtTt3fIVqXn9h1ATF+TKfJdADn98/R9
yr3Ojbzl/lhGEzsUQTZT8WxJsPo1tGM040zpd8I2ArYsNBpnRaMD+X0PPofRFwSK
Seb2nOPv9t5tSDjeXLasjnFFIRI1UWGc8QcYqbCNZGYawtV8xshKFQGOFLF8Gse/
eC4P25/1FtbS7oaEsTt1IwNeDi+3dR8p5NBO9Ew0VTP1q2NnG3Ql1bNMn+XyQCOq
sNl/BBnRLTYPFkD4Z0IB6tsU24zxLAgaUxif8cgcS7XWim1RKcQHYbUeCQ0DHgGd
H/9+tfOLenbJYb4pFC+w77n/nqfttAClMfJN0LSA63VVai0ycq3vyPPS2t/FEZwx
UNl67T6MIiJ8AjSsKOiXgoA5AVhTmNitXuiEY5Pe9FZnUQEUt5EtxHEjTRWSFc0H
bVvbmC3hF0LtIhJwJY4BqQB3XTWsM9+zKlslG90Dq1thtw7J6oE1ag5eH96psLGl
QxTf/MRuQFBXj1UpQsxkAzqv+jtaxXTL93nG6tB+gQJ3peSloEF20ppytxo33GH8
7k3AVOwAvptRuUheqZ/wsBixPGexL6RWJpeBQ0AFhiAqfwpxRtICgKTUyadHALyu
6Q8bf6gtH83FuHSrN41bE+PI/vXKD65qvyZctnwbc+H4E1CqRGU4A7ZHFRQpqlHe
VKMijRajixUWyVQrpV5Zny1Jax+nbXf8iItz9cdNUcnKfGRWSg+AEcGRW5JkeXRU
75i/ssaYN0sWDfQJlOqD32Czir89qep3/X6TFNIuT9VuxLE4bM2LY6YAhLG3wn+g
Mv6esYV5xhjosf45Ycg4BWXGpfXhKxZPYu0EQl2tLLx+45OMcZDEJzUbUfSJkibn
n/q+W15Tu1soEEo7Lkeq9j+aeMBCli8QWFCCXkDqz3004WAnjOh+Ej3IcWpwz3o7
Z/5RHKNM2FgMqoe4VRKrl9NneDhEkbPEhqBmEMHFc7ocjJldWtUwtAfUwzqSCne/
NgUvK5uBL9SpIyqpYGVliZBISTXJhGMlTunWwNx7IzbaNny7BLxEWkehV4TlEsWq
9gXhWsixjuMK+o4LLrxIusDH1tGZ+TrlcjPn8i154MqQEQiM3AXpucMUxrOee+y6
nGQ/kiMgtA86CQfWq9VzA8sMpOnVfbVmNs1/fukT5yYZh7AND5esu3SPmon+EhP8
RO/Ab5Qau0jR1L+NdmRJZAg/fy6DMSD5C3HPMU4ha+lfS1HpABmizR5hbC3GuPkj
chnxyqBYchNKaqRF1yik936Teo0xtk4kv+JoerLR2YYDcJasGM6PKA30fsOdTVFv
nLR/NNhRH1yWPt73UOTd58WsMRBt7+5wILXSpabZMxPZWqy2y6KwL96+neAXqMDe
EJxj97d6T3X8b5OD+xgTOWB5R2W9qdgB4Yhi+LljwzkrHr0xpHX4pP7R4A6Xe8ZI
iIMgCZ6aiZdT6wACh7GUZb3v9b3MUrigHhUnk9y+4pz2BKiWLGgrqW/IhcT0HQN5
w/1eCijRuI77otkWO6xhQSkQz2XekNyf3QBq8TXpjlHpu5yYU14cAMoFruLYIvq7
w/4O6WxEgFXpkZxDC9MxUvvIIxM6OmEl1tRR8kdS1o9RRnreHWJBgq0VZS0deU/d
M1MdZeEQSCEhtyxizvCoTgQrvZXDQftsvxqvWJaMiauJ/UewFdW6GVw6zGjaFm38
hnWC+m3NjIu0OQ95Psw144Jisz+thRi+HaowR83nTF9MDGmQxGMarNY5tDbt+HJW
UQNlhhilA/Pymzv32hHalnNWOo8zrXoagJI+1qCGwuwVA2BxJnwdTvFeV5PhRMBG
MUFfrEpHvYRHqogOsg2n16vSldqIzer1T4/mZ7IMzjZCCMlDD+VPMPCifnFLwFNa
bS3vbH0fOfZZ8LnNNqfWVoHyJNsP0XQQ1J88oAbGbEk/tEWFCmARR/tBzHihS9Ls
KJ9aiq4oUbC2tYVwJoQBJRooqKjEAgRckuTSHwJCdlyufIIaLPT90xS5m94+lld9
q0P3aAkqmnEQvjFCkr7AxCx+dRByOf9qaoJcYXWJ13/+yZq09UkxEa/jzB2b6Z3P
V1o1w+MxeRy63oreCBLyCNBBNhS6LCKupz2UKmDH8guVmvyosXdrlpENBXbsMBCN
uBztCX8OM40HpEFDtaLHgJ8qUofnCmTT36k4UvSZg6SgzCzjCGjKxnbms4X4RyKN
uunIG0gUXAsIy0m70SUjO13K/9c/OhSJ7v2/e5GJ38ZuQTJJbhvczSlgyEhyg6gg
YLEJQP1zJDqDmT9ARW7M4xR7W+Hz5J9n3lMX/JKAzQP3KqLCi2JWspGfVQkiVKrC
+6jq1cPo311Uxjolglsq0OB9rJvbgohGcKtynmMsp58Jds5Y4uEaSk5NlOo0e+m8
g/Jcrq/wKr6HlEc2uP6Kf58EAUZQcbEOnny23Z/6BzdFCnNIehYI75+L+f/o6A71
sozyBWMHtib2w88QEZYbnbeTapcaOFfC539CN1IqqCwtxUQETRnlE+wNbJc5tdZX
R6FtW5F0QdcrMZzDkwjeQnOppNB0nmob35ZtwX8DE+VsG5Dk5G0MgRxbzW36h6q3
V9gJ7tyZ5VfMjxK53NlKUmBWCwaekANrwp+R/3r4ZdeBXWCJO8DRr8V0zF1U2f4F
xE43+sJT+j9GLybgtT5AuhTugH1AMd9bVcspbbiYBc74v3HVpfwHl4iWx5NccFK9
qHBLX/aHnQNblpllFbQ2hgfBZK+iwNHVgq4Ol5BQ2Yvs37wOPNkhrrbKkT9kBS8Z
Hy2Po1rJiuHDPZj8CPmMOdSi5bA5s9HtNfbp2TVYPmOT1QQQfOgC9yoyx9TSIHkn
3639+VBfGVyFJmgo8i+yZBRQZuwGlF0fSImffoBagBKtizD7MVA4ggCoiI3b5aZ7
+i+dEGCqC7hBO5kQI77bBRPHY/Mtf7YnbeePie/HT+MyNnGvCmawwNkA+ILJvysO
pvjK26JOBWqlc1mKWQ5lFkRu3h7pKo8GBtacZAglCABXlLuJa5rys3gnoNTZxQfz
BSNUlix3VkZpYCqZRrbsMYy/WaxNWeevWu6DLIEnI57z7L7qRLJFxewIJ8xAwKpS
Ro2u3lPNVtMrprEiHITraunVVlM5gNDGG9Di9Gr88jZlxcPgcjMo7e1FpF8dmt8u
TUjqNO2GxaEHfG4xSTIAW1yBcB2AgRZKpZZT6ayYzUqC8VsEMQzVyiDZqfECSMZ9
vGewzs/ZP+jT2YWCMVjM/uVmHWtyvPVBDhufW8RRxlB1fTuaAzxeMwPtArK4eU6n
KD0zz8fARUeoRIr9VYtiO4ywW56WGcW/hCn5m+lwWaYnZ/VQfqhH29UsQQXrhV+L
/+4B53ZTvUggGPY8uqNSfFj7iGic8KA+9keIOBCIa+Jd2pJpER5tS3f1SOrymCyj
53y4RYTxJO2il+bbwdLU+ACqQGEmAzgXMzEJrWSZpOV66k9xBC/lGB3vpAH8BvcT
hhFtZoXTizSp0vWZ3hAawT8wLZtQj2R4LnE/cbE3CXnNv9p97fLxoeXAJt1XXt0G
or3nfImfrDTBLRsNmjq7HX2ikmnLqwacBHqpIr6/WCWbBzbU0lnB7bMQpiOLnMAj
de8gcwjiR+HKmQYAutuzQ4iktxIwzMO/R+wj3rqWiqNUeYehdMnQWu991nbVWtHr
8a9V7blHL4UxqPRKBN3VtwLjcNehwKj9JTxLubdPGPcRG4uZsSarNkHoiN7w3BFA
jNn+6w68XZ+/Xhbhq/GAWJ2vCItS+93Cvkt8y11OX+wdMAaAb8F03dbpzQgBDq/r
oNfoI8UB3u5pQsN32OhYE30QKErLRapY/AvIEJ2he2DB2V5w5Jbur5qM/Z3CO3JG
crBxMnXHMSbyV7De8qHxt+x/OWyc0RUTnMOjEv9SOLanYTZaUF1OLbF0ayVoit8t
5L7eTLVosclxrSLBnlDBTFAxgnFR3fYkWmeNv401qXySC/vuPDMSbngZ5yQpcENw
QGrEgEaVjh1YFrLvB+ZFOWOmWxosK4+MYIA0whGq63oPfpYGvtqqyDrxvWUpPc6N
MQPmru0rvCZzmuVcnPWlGd/zY4rXT8R+gXJr/RizGL5FCkUPRszb1bTsgxOl6pGT
1k1gRK2mwOuEyU1an/dCMN0O5TJGb3FQzIVETPxuVyFpGjO7d9S8JnLkGRFWXBgo
WDkrQyqD3SzyL5GwxbEOBFwYjesszI7aLz4MacQj3acFQSaJNQO5SLGKESHmT+y6
i56Dz9uGmGPfaTdThUcErFI21NB0BMBLaFyPRGTyVcMSmzpx4iRf004T5kaqdQIT
1gC0ifaxUlpP+IUwmsUhzob/WI6AhBeC90Tcl0PeLLXjQpgtfsJxd5JKIJQE5icA
m1vpp+uTbsSTpf2hXzkFAbNi2s5gxo7tD5ga3TPQ2AQlbpwhzjMctAzirUl22vvr
NflTcIbbNBAiGzBcL8vdwITOtgzOyMeMZmgHyCFXXzqey+ppDbKn97MGj3S4nm8+
8xJXvR1cKA6mF+xU+/s1hlmzrNquhLWHaoCYIundG6LiXdgVTnsfkRXVUQ7XkwMp
LEeAR5HqwhVuFVwfRseGgbNBXl6fYq5FT53k3K6Lyam/f2uoQXwQ9ZvbR6xChSud
j8M5MXwJrvRcghWB57ILislRkTC/rOqH+Ln90MU0koXZAp04v0c3IAOLWWeWlpZj
ByidmDKM8bpNu8gWd3JhPb2ibYWhYu3weTETDdv8x/8oNZGDcwQBM9IffRiKHSOK
tjDjdieXTjHMK/NZgGsLaolpxdBzB26n8/7VKEcnDRppDs9s3/MqH2b1qsfFUS5D
ec4asVTMTu5XV7gbkdlLuW6SHbSgJJLv62Ed4dlXjG1T0j+pqVFo4VTG02SKAmtq
HKh8vd0kf+60+sivcvccfgsWtEcdCfGNGliw9OhZX3hg6VcbjS7dsnkLRWUihwBF
rAOLVE0nOngg7E9NQUBogChHijFHiHFGDBuNUgRsogCECWKlM+m9xKvSzVrpPMpu
0CCe7FTZEtb+GBW+edv7OlHn+/UsOaqAavMzj4L8eXSBzhb23jXQh/gkBRc4CQVI
EHS4HpC9qJIPzc4aGCgbi8aPj826NnvqI7bjmsSA24BdxrWpcP/g133vC3habn9p
pItzWwBDVdoiHNki5v1yYnCKRfgxA+msQpOml4IFpSQTzjtQ/SiiCLPi4hJZ5FW/
LGSVBdGXHV+0Dq0ViLkfqjmC/CAvfppanIoJMQmH+GAbwLzbNtQSTproHrOU+yTJ
b6ZPnP5akS/JbXk7uOPDZu71Mf1t+eHLucOexzhLfm7n0Ge3b2H2QS2B1n4ObqmR
hSLkw/zcFGNQ4y9G2TUPRAvxUYf/A03E35tP6b0L22HJfckKOfEOOUao4x15otTz
V+nAExsgISCHXqFNzyw88i1IjTeUPSfmrXrSwmClxDSKPx5XXAj3z1wSH6kdSf8L
ZgSeY5ls9CH4ZbKRIr+S9vhrJQHjYJHQaQjIGHF/kHrqq6nE0HJi4k+8suSKUIDc
bglJNEbUWIf5GQwmGtO8ZBhVCYspgD8oiCdHZxaajbqEUBfBcGU81JXvR+b3PyPb
qDWiEZIq91y58znXMMMiygFNlsgiN+/emYTfyvQO30Fjoecxibf2YRKWvxJsxfQk
IWwltp4FeHfbMqU7bHIDFqTM94CKLVMJ7jRCqeFlDSQlUp2/kuw+nzjEq1zKKgdP
4/gPr3D+IlzjKsIPMaDbFSMklAZZPD6n09so/emkLebXZ6sEeFrrpkBuaC4reLvx
UmxsV1Q2t7nJ0+QmsZulMTB7IDnYmUCB+PCmewpkVWepOtKwNOM7lZYRTAwAIxx0
f8GBCA+l6qp9yl0SvYr6GLSP48XYo4Msat57r69vQeSm0/XsBUjbVdJikRLqIb90
eLfKJPFPv54KWt0Nf320GAjbF12tIcUPVKAX3FVui6YcPta2c9SVMeHTs/zD/OPE
ps4el2sOiJuPiE3gLHjXOHzXU45sfZh474gEFqLp0NoJj3rA+aXLRbFay1uMCHGU
LtrRKnXSe22Hjk99fPM5IZavvx+47dsKTX27hsKNe3xby9Fzbl78mZ4eQ360uQne
34wSP1YSEa6/52JTj966E2iM+2E5Pq9djjYYAgShTJnIrzlBnWzyFe/f2LUOzLbW
OMLofnInSCEQpJ4JM2KlIJ+uiBnEZzRWVh7bO+5rHDdQXlHA9QO8jpisofEXhof4
m+7VxWsmyOdFz9w3seeG9ArDfTzKrx2bNQdEW5AzKFPKqctGc/r+7WJ+VYuynPi9
r3HknOQhwYQGNBdZSCWEu5pvZ4JU/EDF0OX5YHInNcGaCkSKXZHZBVNuKnekKu9z
nSReRWrHpBiWqasxbZuEyaJpejy6Y0s09U30+zxcVQrYJav1GVvVvLGcUMdVDYtH
hh+g+Y8h91LOBu5W5IwQPcpH5xNFUnoYmwmwv8+GwWSgrSRvJXD4AwxaJ3P7/EPE
ARe4OgvhLccpT5EvJevN/jMEMKSPsVKylqpE52MT2se+voODPQqfjKRwrHKfUXnL
4niHB43pbeD7anYchnTwjfs1mjfQC8YdIF67bAoEYBy8JRAlx4TzGs6FhCv+Akk2
zwRVJJEpcj0No+xNMzx38Z0y0TJdU2oEZA+nvlpuh9mulpXIwvGpWW3oV/ShYxx+
dSYCOWiPQpgU9XY8Jxk4pkya05FJg4KNlgmqqJ3E85wN2lbDfV9AkkrTZ0IbbPzy
N/Q7+I5Lp5/g+SzcArzssgUuTrHBNe0nDLZhjaTXXTOGfbw06BzBtm1HwEzuXzJb
M6c4/KbGvUWj3fuVTf+OVpPtDwrje2KLnHRPu3D+6lfkXDvyJcuBCbwr53+Mn3Sd
mFMrxSTUXHKYO/hMNf1g8BOOIv8HOI1dAf2MIMnWHm2gTRAtzuQA7GjaTVFyklvb
ySYAyD6YKJ4bH7Wn6EVBOb4LlElGGfxe/qehCwDQCNxTDrluBHv4fW4Zd5yIbAq+
M1w0qhoIBr/wAl4rKsbFrezmcqIvTFZ5MV421GqPiqT95/ktcgoQTbDv+x4Xwe3s
CAV4DaCJdMGXcSYtgm0so+LRPcAWuNWmnOlILPwIFE009caFtKOTEsCZPivc9DuS
EYSeNuTJ7KdlrEZ2ybiOTqnq9smRPTuvLpDN0/RbwfHIA1HEVjv7clZlsodxjmE8
XRSym7ssKVHbcHMFBf+qijPdYr7IC95CocmNU5f/BFYhOhZcWESEidID/413PaRl
uNsJuPlJBPtnU5BM3SUIL/1+wtf3vmBybaHBsPtCO7z0pfqQZiiKZWKLb5GmHWtS
4FO4zDIED0LOOlgsSPWQr222p1OBscIX6G4tHCIDNeJxzMh+Xzll5lVxeZ3fqYZp
msKp41ILW2HRwtFXt/zurrT5mKhtKcgUL9OsiZEgYSunLjIktLxoWt14k3qgL1zT
jKzKuVzSOr7MrFY48bPbYv791WHw6uoOiEWM8fnMsSHDYxcMu8WeVZBbaOOwqgs5
s1Osh/G/5LOWckva3jlnVBQslUcDcrhL0Nnhudqr77ROiC0QMU94m93OkkTCHeHw
X6KF8ek+9nZaEVmnxVNkpK9PXdFZe7UkYdEHXxrb36XmQnZhbcArYI/hoG7icX0T
ppsb3lT26yUsCtC6pNLxokngP2XPX9pH9JGyGBdvUAb1MIptym6LlvTx0n7RavzA
+lY+eQFnb5hE4W036fjXHHq6wZD4JTqB2OJmAjwbPq0Z7iFvJ5PhMjobYu2V8qXL
yDrlKYOxadEGsM3zU9k/HkEvNCx5Cm53m4T4BVoj4hV8gtyLJ2sfOXrZ6Ue7FZK9
+AZDiT+zYx7MtX6assMwIgf0BcWb+MPhlvGSt4bcAc6eHvM6jcF3e5toCSB1JLxz
ifuoKy8iNYOfLyDeLHSslkWhWLWNcR1o/obyrf7lxVXk8wOsuOsXrH43yE3QLNbq
+BzDFlDKgFPA/D5NcQkMaRTDqo9mHbzIYQyLeAbQfA35q6/EfLnAklFLqfGQSal9
g44/2MHl+aWi/f58LeJOCBFlLrTYXCvi7MAOvOqGXLNMTwTqx7Amb/OluE6MsWeH
Anwg4I2QBnUYq5BVvmAk9JojWZGdTCNHjtaoToUCQ8qrR9rXmHo7BnETted6jIpb
TU8ja25FjuaPV0lfoXfB55SHBswg0W6h1EiZYCMdfGGFfxulSTQ3ZJ1pbC5BpsOl
gTtBfyb4CjfBSwNvj+39FatzNtKq9i2bv68Pj2S5uKxhX/1L5zUZ8yI/25KaQ4lA
V1glWhFLmhLjwHi2stBM8SpWzDOyliswdQVutEhOPD4rIlA9umC29lB8pos+M49o
sj3MTmhjZ4iBpAKStmTctz7nw0BQFf/1yGcQeIT9yVE9Ngvf8nz4p7TabgEoJTLm
lW38f0bRSz9vV4lJNdr7ARa/dRWAI1itlA5SY+fF6tE/vGPjftRvjollD8xare/1
04F2PwtzBg/z1kiL+5mILkvPBUGtTzDEWW42IZzAzMihscX3jNSLetAEgrGjNR/U
qa2jmnvO0mJ7ldZHUEe+Z4y00Saa9ULMCwiACuHZd80bWg9GdoMdBFGF/shWoMIb
WaMYQEz0MiMSWHP2xIxpYfbUbrgzHuEH03HqLQMQuRqOA3ZQmZmWInKWKimD6zXR
1lGi62S/4NPrUxqT8A6M52wZroxae0syafcBXBVaawpD+3lKj8j/xP8ziiyip4f0
Dk/q34Vn7Azh3ZhgwjrJSY1Fv0M/Ni+4txNiGDSO0BoWwSVNBZQOaptiPt1DhX9V
mL6D/Nf+/Kii61Bp/e+xJZ7naK0gqzdlEQWHlU1iE9nk81JXy+qFQByUthrELIJA
epQaU5zlO0j3/QbeQ++aVJuHZAXbyp7NqnoM1fMreNnUgc7ta3LOMtvj+NmFLztW
9MJKNYSWU13HspcYSrLHrupWxanXa7euHXIoXITRaru2yGSgVqXRbFd1tiizTvxG
9mcbUQ9tw2+/QWv8SY+beiwU2r7zU2oX8D2PbWKZMGrytbfzhQOmTFnu7ZW9Fg7+
vtUT7SqPbG/r+SCxZYUgIl9RiAdpH3rCji0poKRpRHbNkejn++5zUo1Cd7iG8oC6
t/6jP5uM8H14sNOvRncNHW0KSdlDgWmDChbJB+/5ib9sBdajGN5jpnbYkQRDDdo6
CIckoSIHd441XajQ+A0Z0d38cdm4gbCm6aGg8FswiOT8u6k21McCXkRLhNtHEJ9J
qTM7FQwrPxLPtReBPWYaYeyXs9IHbc+vsjwhbexYeaJDUyshHwMqiYctMh2S5woy
E2N9WOrgLGxCPIHP9XZp4OPdGJnXig/mE0N+OrRxaqpZrtKyIjunOSAa1sqax6Xz
VhS+W36kNhDtTUe7G/VPvu+YSXVhhje6WKret6IL4fKI0oZxhWKTsxN7F3Z5jRKr
3eEeeWArS6XzcSknppGwZyh2mh0A0G9AD8mE59jbdwxFXpJ6Qu5aj+mVl9I4a4Ts
p620pLoSUxaaRxP/38cXbepVD3WdLxjcTNhckfrPwKJdnQ78CcO7rVman2tUmmBK
QKLRweiKc0/2PVbboqoX+ejCTwkytonsQhSduXEj4OabMawqYNP2ysnnfPC224gI
CIIASX+jbUV+n3Sz8veYUjrxk+giRepuhhKiIrFnfMEsdmS8ufe282C5JXvnVjvK
p8NeeydbJZFjqPoceM/ZQEluuc9xVOPu4mS/r9dnyrVZETM7Qiat0pWXmA53mph/
rKz1StBdcAU6APRPGxhsUAINQMdX1FO7Do3+dJrSgkhfl9c70UBGt6gzCofGvX63
Ces9W6cDkv8WF/AVoYqknYcSVKogRdlPuN2Oe7zn4oS3mi4gZW56g/WCGHQTRheU
p9BDWXR+6vj2s7osRLYB5zYgh2pEgo1MR1EzrnPlAD7U0XRwnF9BhCzEh6DRmoIe
f52x5h6DyhxOMtNf+EnLmA6AlU4HuO2sETn1NaYRuSxWMnxNIJMIziOczydcXUkR
vjy3DilA/puXAya+OGUQUYgqcNuu3+hEXYqjnM/nzVY3D0+FLpqaxwYmOf/1HAg4
XCCVcCnO6F1T6EeFGVqJosQJbF9CCeeJjXxHHr3jY0ODtIdvQ+dsJIFKxL/6/QZe
olMTUydnVuApHrIdcvoOVu3/Vo7mF42JLRY0bNbDZEih8NfcUvQXbeBOMBAztYAS
wFDsEkVCJM68MjZw7Eja0tLZQTEWD9IllibSm4b/RKp4+ZinNc+kgx+GZjZNPsi0
sLjVIc41tRyR1P5W2vmSRJg+gNZu6BLeT1jwhw+i1vYhDhiq2+t2b+hasbUDBfcc
jgHb3EeBnqNBXDDe1p0ShMN+UtZ0W53cHdGO4Jh+zwJMpi9VAb0a+VkOSNu21fRa
vdBJ5hSdtwVjKu6WnBJ2M+ob4RWc1lL/Nn4MNN+Fu7Gww1OAiQx+bH6OUDD2P4q0
g0EAnhH1qO4IhGm/xyypLEOc5ylEJ6DRfKdHhdyrz1wLnlAMzrxkL4uLPLlW1CRE
r0jp/IhNRKaVP4M5bghdjyJ0LaM02jmSxJxWALTF6b2/pBkhhfZI/dbWh/rGMXw/
5MPjDgey9uO9KN3Yeht1HeXuxhvDHindeBKtrQnzHZuBlpnOSRbgz3zQyZD90av1
MHx4/Uz8UP34YJRBITurSVbVEhcZldR0IhjEAyOs5TExXNC1HHgkC/pEqk0BIqyg
I7nA02wnTxyUrJ1my6SaOVeZHfsYyF9MkEBnFIn6suzMAucF2DE8QQ99rT761N+h
bEhNVghp4i/K80AGkVv9p5j+6EM4cHCcj+yFvMRnKHlhMof4Yt3NjORko2LqVvsv
MJHmEoeCl3YQvYvAIHfuLk7CU6MIotethLyhtX2St5var+qOGoUix03ldoqjeoZX
4d1XYRJLcWjKwm0wOQ0yzQZrTdcV6CGlBZERuUdBrR8G9+0Rg1o6z9zKb/ivz2of
N+CTbkqh1tcITCal9xUGPAhDYynkbVm0UejHnYTbXvOclhhHRl+FUL5egN2LwlrP
YXwg8H3Lcc9tXwIYdcOuTe0Wl83k92SL2+nSChXvqBaVMHl4TyBqHn5AsUZ3xWrP
n5xqeKxshqKXaB+GR0pHi63Uc8fPbwtESe4a+9C9HiyJk2PIsioo+SMQozkA5SJm
z/T9A1LahdxbkLcbg2Cyso/j6q5l6CPwWb13wjw2qIk6jq5Ua25c1tiDsX4kE3Fh
rnm0ogx0A07csAQl49bHeb9YY+DgdLaZqZ1M6Dim1OmHBkrUWDWPVxQwx9uV6wuO
9L9d1eeLMtgbkNHMr4cy2vGHHlTVR29Ue+nGasrE9OW+DgyorQaUVa5IINZ4rFcV
8rUzFeWLtKSmRhAIWzPXJJ40yFcWEnsfnlCRh1nMcVV2BxpjMWAl4++92NjhyrHn
RcH+YbBMMujDs7q0kb9BtOzpY2U5C2bER06AkWVsO5pUtySMkJhqhU15p7JwTojI
IeDcFa7vsNYdeLYxHAeu6GQ+zXp06oU1EzJfPjkHSEWqoQYcZXoihJpvdzZlg1T4
flOHnPxhmj/2fwAAfx3F6OzBccIWT/rtcrdzMXg/rWk3CrmnwlTq47KST8mWJ3zm
O3i29MPQ/kqppicjif9U2NnUCMnQ6uXmmrmsCeNIenQCMVLa3hIhY7c1snWKQXE0
RojdVyVHl1zIkH5IUg7KBc2Vq4+ZujFvY4ijC6aH9+A3TSR5ZPCpqv4WLUF1iSKw
i1OhuYnJ55UdzyQia0sw0MznnpGcnb0eGV0D1qMr6MseMztumr+QhAPadItY1cyc
1h868+/E8iY3IOuMhzHYsLjZffWqB9AYMMmeq3VL0sFNvrEqZ2IoWYkDNG6hp+DX
rEAIW4xTaM0xNHhV4JckAbwMKmlf6447CuKEZaelhUQib0qdUneoSCxwaATA7mEd
45qBYRzAMEeLxIRARQeFXNAehbq56u7hWyPb9+ufSeox+yqaUy42GpO/GSzBAw3J
CElDsuoI43s1dMEIp2/Gsea2Q9LlYY1FS/Yk+x44R4jHkGBF6O5A39pYeIQwd3rj
ZUZ3kNTh6PAzegWxelmw9tpP+Gx9DzKFDPPX8ACIRdr4KWzhvGPA5BeKZFjai4XQ
gWzpM9JWYZa8kAVaGBgHdIfNncjZc2anenCgypnO879PjYCbbDID1q2Y0JdBP5Zl
2+2IY9XKYk11Gatl6TGl4NSTjSccmUpxPLDlbH5RTPIqxEhH1VujJBgXJrqGjwDr
2visD1uLEOnsh6/5JnI44cL9NRroWT9HgauoCjuvhBzvAoxl9GaNfv2v6GODBuN5
uf8uoqSE+meYmWa9jmCY5NNyCsKchxFevXeTowP4XCnV9PXt+xTWIvmDKFDKPoGQ
dEZMIlw/91ZHIwPEVCGSYK7f+jktLLT6JJwR+8PE3xZL4qz+7AH5AkTxz81j5m6J
JtIj0E/GHJUa3bO4BVdEX1B9CddOpWZrEuKxZXi6tAXUjrIttBbqOR+VGNKJBxoa
h/YyOB6MPWAOcSFUFmR4PAyC9o73RbditNU4ARBKgSedIKAkmewjOfQ9cZzSeB1+
VyiWhFLhoQ2HbLKG7DdQJtkgFDyRegTiFK7Mg/hZFZP6ZGTvuIqXJ6pCS+UUY8fm
i3L0tBZ1VaAMzxDpvWtj6i/1BIg20s99gFuNmSLDF+T7Bbr9WTzfI34RElemX0w6
/jOqCcALGqM7AyP/brlITIGqq9IEwPRycogW+yaX6K3hfW3qi9xBaDvQ3GHwhPyC
VguT81lKtQGKE3TFPUvx/G3zEtPTfGwVJtlgmhb0ef3cq5k1AJz//aok+w5m4+XD
3yJtn/uwaGqgN55YKRYkb43hw5ZMVFHaLQZThMM5D7bYoxWFfccHGwB09pPlMeTA
8HtMRHLTX10//0YIAJOop/27Q0INQVuDJ8yJfZHMwG5mZddbvwGfed11yl9dfVzg
KlPbCI+iZ5u0RgbGfpg4QEElkAlBPCdzFJDG1pcnfylaDM4a3lcPJFl+8XS8uimf
MEJjTOmlFqYIRuADgRs2R+V2+28hQRRP/YanS9M2GoQvMWVpFVhhhVPSHfcCIGd/
zzQP5hBz1ty4e43cseqe5AEcb/gFoWuR81Rr7d+LN5KMlWdSpfMYL9ch/vvXwF5J
OqXqTzF30YGaSrX/2etV86AO2IWdXNcQeYqZhXxJOSH83AGM3fBA12Xp9Z5333u2
crSX6MOsIga2gE5Mf3MNP+MfobFEG7GDA3Rs2v2gsu8i09vOlhFfcoMz/iydTeSN
cWg1zSjwdNIaLyYGpUK8l/6SrWcmvdSZ3q1bxAXVgJ4mPf/S5AfDxeNeizj19isN
Cl5AQG6OB8k0EmruJcaALWFK+si03RlcZmCPlK6PXxIEUw10CM97BTpGou8iUKYJ
oyAklpxPv4AFCL65Jk6YwyqLLbSvqY2Y/2Fp5JxDle061NalPsyKO6O3AMSkp7/3
+A9AczcuxIVVTkVfPSgPUw5UYiTCu5dEXyi7zkPrUOWeiugygZTHF9PfMHiGhvlu
9Us+m7yhGp6SHgVw7q9nbaQFddLH7ZTScvP7u7lWhiOygmre/lK8fWaWOazPCVL2
tPhm5HTptSKy5f1tfuV1mgJZfXqDUICoXfto8RTHPOZ2c4+QznCpfwJjDUHkwaRi
G0CeMgE1Du4iKBRWbxjX3EAniy+CZxmdbLZg8ZDKxJz1msOV0f6R7kwL4w5ZRgyP
R+1u7GzzWW60TgmDToMdGSMor333Q6zwXB2jrP0fypbxj5zvkt23GjAuw1ZwVYra
ANJ4hziQD9LKPgNi9jybjzqhE4GNPeT7PPgZyxtfOYhlGQnHoQlBlG8zDVBGbZSA
xk3ajWyhstIOCroMM9g6WgpclbTsdz1B5sH06WdqZ/ezToC6I3mnzWblZMOpUn34
l48G2V6Zs4o60r+CDozRZt//bGD95C+BfZ0oACQlEIHrbi0S7BeHtlo6npdE6sZn
G2Ed37ssV6xh+GjnxOCEG4QFF5SDBIzMsxhW0RtbbU0Vx/YilS80IQQbx4hWSOFn
AYL3eSRraYFyE5zkQwLkKO2Nf8a/9C4HnfziOvgvF2sJ3AMB42D2t7d47UPqzH/G
ustJNPJNm/iTdzE0N2z9PnOrnbp12X0JUyCabiXEx8jAB6rb+I8j3IAQ9QI4Ke1e
LRRmwEQUN5mu1Ez8A8hkDUtq0zPOTzJtYprvy8zoq3TlGVeuFnEhU6PqFeoUehe0
POtWTqj7HyfkQ0Cp1xDAnBvSUjVrwR1OFJM62sUvbO+kuD5WVN+XUf3ShgbTb0F3
6qVjOlwnCh40l+YosYVhM/KpgVTXw2Pk2xiB+dU7eWbkgt2AsoJlCGGSvs9fBEJ0
QiF1Y+MaxdhcsH/m9sqFlKDQtP8ZcEgOwO7nwcKqEg3yRJdT50UxdzqcE0WPIqqG
O2G6k8p6POHlkJH1xp/oNvCwVfgvGi3yJIVhVujfuXUH25LX1HhbnQKF/9EjYUMG
i8+9cP1lFdbNAHYd3+jNh0WhhDd7QtnfKpaTZYI7BiL7LKhYo60S4efT/aZ52DGU
bqacx6UhpguSbfHnCrnXV4sX72spl1F6m7ihJN9Kr4kdpOtLHwYXkftekLl5/MIa
5x50FK3N4XAgzlv3dj7jd15WRs+cSc4bfOruF3rXa7e7PNoaVZ16KpnkMijiomB3
TpSpCy1kdfqTOlsZDcy9zrwyf9MMnamu8fMjodD7AhdM5D+DNR95hy8s6EAm8EJU
tL+De7VE72oRkO4/j1bbA8byWsEsfk1B43vHciE3dJv9cKuwAQDaqdTLFpU46ho6
dq+gH+gp8nZoGyprKJyTlT+nvpUx8rOFRm3SVyGEoqE7oeadYl1vMqzNWcP1VMIU
wFcwdL1t+vunYi4RTcWa+CtFO7S9RP8QPhnj67fURpoilTq/5twEMl/yoZaR5SMG
qoxCwg9BcN29KHl9lWki56woPTB53EY60Pr+Dpv6Oa5DC7l2h/6fzgDbJuxbwtp3
1sCnhdg4DiPGZobsvMOQYT7T01qh68UlzxBvrBCHqJa/pS74X7aXZ0tZz3fFHVWS
sRNKYLcQmFpScHTaKLYITpbSXOO4hK07N2UgHZdRLSIv15Iwf94lcSOujNevDh4J
7sKb0OHg7cQnvC7mRWLYoXuz2IYXq5aQHXGgyPLbOw+edIF9G5/S35Fg7k5PKzof
VhM9N2NG9JMOQSQDAGXNgq1plemABmI+Ea240yGQ0Wq809/Y8+HkDVbZ7rqA7GYJ
np7p9Q1K/vvPIwwvmr37ixAAcpivip4HWQs4AcLVyfq4h4ooYS7v/tRANz54J3k+
wchdRML+SrpRS4DhIhSKBTJKF5KfQjmUrJM+xbgWa0Ry6qSUXEP1jj0s5PGfFdRY
tYp2mXbSHtm+H7RyPa/Zu7AD9miTYutL+m9boCaY3gXIMfYQKVmoi2FGxsED5csG
CawWGMPIxw5mQ5zAaWZ9MSoSrZbOM1halNGKOmoJjvZwqi5UcxdBtW4cYruNwBzR
WTpwnoMOW5X3SaKLlyKdqMpTHwGTwRVJdmK4D6JoEXKPo0Rcog0xstaU/ZqiTVVg
WNQRN4MN3ST+Ka08tlI9JcO3D8s1Dg0bIj8HM7URTZ2+HAXbqi1Behj7iBpgD93f
eTuoKlmClCUH9X5THHpG8VFx4/snw/Kx6XC7LE2CblBt5wau1dEGr8CHRKFMYN34
1mgy2FGkEp/WVkIxPemlVNj9fAwxD/ld1p78DigqSTEN0msdeorw2YzyY+tUO5kz
ny3OdwUZylS/RUER5TBQuxTNfglY3xce1OIPx9aBd8NktcfFmFSfLsvyIuawFu2u
ulwVExyYcUjTz9gegcU/n53C4XfSUF9h45r2nskzsl79vxSwtgNJD3g2Tmf9cbaG
1K/cZLA+6MVZFBf6lS5b4D+48QfizccHQ845XGYSfWjol/DcQppV9KlTil+YKA2Q
5ShJmjL1vOZF40Gr3vOQoXsIQIPgEC9OpygaZXLw80Hll9PE9tl5Ec6TcxYq8T38
pr1IyOiP5qC8QDUK3mm7XjeJqHbbQcdhfiGdrzXTmAHj0KBgmmXhtQ8V0X+dp9eA
NEavVa1NBX3lnyZLwBc7zVoAfmhMig0j6qO50gQz+8PkuKxduaMeIbGLoe9PUpCk
oOJvptqELngHfQFpz1L5oWKBOjRJGIloduDMrI+QMBLDLyARPdeV2s8ECUhHUZ9l
6IG3m0zjri3ND9l3rHPTiwCC5teqpXP/4hSEDjQ20Yx/Cx0iJyWs3McyYekgAo6g
CFDUtm4M7D346yWekP7+KrhUX44B9AzqgZjs4HcvsD7dNPQgbjDLF/L2T1FRP28r
SuB0jK3h423hzufMe5yRuhBuGT65sgDTihBfuGqFgtbWT4G6oA7vRdf5bYUNY16+
GAMyE4v9GVWwxNfbGNY19Ea6wBf9okwNrP1e2mkoQJfOH/EOz6ydgsHS7ndPVu+o
rkx4lOjnbd6rAKUjBInI8UcMzTe4/e2ikbgpVFXZ+0cLaM7EJXrOkJ/rJH6XISrv
w/oJ6/Cp64gm6nA+06NVk3KNvFM9QXN5j0reftKbMnsFS0GA74CRluFEer6/WCdy
dNrQGOmcIvqwfFOeAKG5lZQTfVoIL5QS3EcfRLUSpjXtjfqoNyluJtrovkIglCrL
ERbcH3Kk8axI7Km+dFh/ILFSNl9JhQs+0lilPgtqs9yemikE/e265+5/8aStJhZM
O13FwSvsRZSdjItwjkrVayXnrW6PvUJ6OKMa9VTo2zHqWbeACvHDknvo76Go8BGI
qQfI6oxj1x4j8SSTkebSWSyJZXZ5isg3Te7k0rSlTScERBOuAyw6ej4rWu+q9ZH/
/HnfVrA2ovN0gX1sL4/ItoNQNxUoxmng+D1iNMFQzPA3ij2n2Jl0H8CBni/9YgAN
BwiWRutl3r05VqBD0DSJ8rU4If3JWvGZ+NRKBNEbJ/jBA+i+B/As9IwvL3yB7qir
S3+rUxhPBQ0YWgQ1GR+J+DFT7ao17derc1rNgD9sa9k9di+bJV1U2s+iwluzNdcz
V57PTrVcxQaTltJ9NBSBlTe4HS7cx0SH+WQ/rwJJBO+vhwX4JjSu3POwTcxKHe4K
k/9Cs4BW9Fnu6LaxkkiQSO7ui0X+MxHSbUS4uYQrt5PLD9YG8ZK8OTggXm7/j1Tm
OKRue5j+121DzGYI2GxW7kYV0aLC3BiurZVAJ8CLTFPEds3KmaGQghdLE5uEZare
AMAyHtsw4Jq6F7Qpeq9NK7L9K1KjvTrJYqe6seThMP2IvjTXGOTc2OisOXhNwx9j
26ngClXrccvA+iZsXESGKtgheYAVnXK2BV5mGJZi7TpJmukSPAfpgHFeDxv7vmw7
ABfKNhBRDmYspcg8/mzzxarjRn1SV3GKHTS6Pcp2bo+S0EjVpT4vRRpFqTm+L5Jc
swM4OufFOrBuJ/Rzj+UT2r3LOQkntQAKo4dcRaxRx821lDOUaNKcSR03+JInPhYV
c8U4H0StK+mB7gTu/M0diyya5uK5sacUpLRaq5kMV1yI3iswIe/m7AeHihQeIYWQ
+BpS2C7TEmo217GthFoPIco4wd+N8HgcCU6NHcB8TMyN0qKeUSH3nI7fn0MUcg6o
NIOl8m8m02RG8RGotHBqKv3W11clHuYslhtLHeGwYrn8hh7YHIwqrYQLRx2LSIhp
WPoD5vVHHYheXs5OBUE6f/2q1U2dnvavxTslnkfI8AfyZkY6/9aKAKKVc2y3iRaL
/X6vCrsT7OOcd7pPPWhZW+z1RCztJ4y0ohjZEeftwBe+Sp8J+qSrgsINMxni5z77
p87GFq6cLDYGZxvNDxMk4pDDivV7I7Z62t8rApeRk9OT2s10o74EDJd5QLh2fJ2W
Chp8j3oNKUjzjZaC1NCnHbD+oNa8wD7kTgi4gvqq/2MeOMeSjx06/TKhnj7U+b5h
CGD33X/BX6aUB4UlMCQX0NgB4dhBOq/6HXjrzKmGI3hg+ZxDuPhEh4Nhoa83QhlP
y8YpgYG/SfXUgmHydmY9wENvo3BNQ/JLR5k/0PWDwouXwrXSXNnMRDkxgas5rb40
bFCtr8SA5MdKA8xhrtIuzVnsB1SZsExkkwWskGMTlXpzpPxPUxhLTPgpvTq+eRIp
KGhOhWVKPh/ZEZXIdcozBt2aJ02BXLASeKDW49Gy2HKaFsIuELN0+BX5dHt23YUP
tP/WMGcVlEJEWfqOmKlFCXdFjVhx9iDJUlQnDEBDyqQuEHcND+mC7mUvhmPfbarM
TiMtXIB4XUeNNixEjXmFGuQh3MsRL0MW984yg049TR9okFB4aDgVs4KKP66jV+LX
rR9cxtiC221XOSgDvz8CWYFTJg5hfzOPZdihJ/qkaG5fqoCJ2P1O7gn/JaHkRVgH
daZNgr90v3i6rHR5o0mG9eMsAu7zOehgQhJvJWphM2nQdtOHXXaIm0CjM3IA326f
qXgsmmWfWFqfLQJwzPQ3T3xcG+aupwZPzPAzh6i8WrOXHiULoovapH+fMkWWA9OS
HLfJhiHgtVbLPczUPHFR0KjOf1E4kCPlCTv4YVamUonqffvxumV77Ve9F5uP8eoZ
kw5XZ4fP1dUEZadbgOZC5pc1eYGrfkkD9HTFFce6Xt/bcsb+yrqjcZzAH0O+f8zc
Xt6nHEuUl/zo9+elYwLgRtGfpOxL/NiCJ0/trBi1dAcoWHXmf3+fYB2elzwrXDaw
yEpZMAIPRnEZgB2riRjRpm/4091u/tq5fXZkCvhvcUYsZ8A4lhEZplL9Jwz7h9z+
ZsEw479vYi90zPF7kMHVvXo6vYYD23IhRA01bGCR4Jbe80kJhZol9DFHSlzinBC7
xFIIE62jsWqKNI+eMap0zDcMvWkja/tdgQgBJIbAZ3BV9WwMeLN9q+8z5y2R0NQb
2SCYtDz1aVUEB/fNXLMoxpVCM4c7AGEErLH547MnK3n/+HMSUndx43Y5ed213r33
+AD6VfZtThvhY7EvwmhEwAv9V+S1SMwe1XRo/T18wFJ/RE4JUtz0Qf+IoQvdkded
V11m5lK2H6k0Abr3kjU19PEMtBQcbkbtm0uPrn8zDfqczpQv0Lx+gHZxZ1Qp3Fwb
Xb72XYnINBA0N2HAnfJ+RPa+oreVj/OXJuLMc1mYtbsNtOYABCoFBl4ibZHD8hDh
IWB1UzilWAQSm4R06lOI6hyGmEjXE3d9OsQEH5rCB07dvhQ4ixqE+wSh6WIBsD7F
ik4vcMYvGqcwS3bXfGL4cJRPYEc58AzofMXe+xv6/IVi8LRHs+b1o03B5kFXZWp/
2GVKio/BV4IkoXEaENC/C3CdYWlc4ZllBmfQCMAN0Rvo7TPZzqWaVTe6gJVIhQ0v
bV5143mXQf99zqXT2ORmY/nqhjtgi/ijVi7XH5e0CsC/P8N/DvIaWiagvkWXDVkz
+E6VGpq+Y0dwdLYhSC6RZ4KOEe9PiXzt3dYwDmjeyFg2GaKs9xqn42qtXIquNEmq
nGmJkWk6iL4rCzbZwsPdKcHQw5xTP2nXbZLdayKxjmee8O9VlvMCaZX4K4LaEKrl
cLicKS6JSzcYnqiS5cb6eo35GdG3N7adQl9BejJBrD5UcSFroKBqhQaVtTO/fLB2
ADhUMiIROKZUOZO0QjA3geNY8XNwISSTLPEVtGB5z2uRLtXGcnPYcoZaadRAj5ZI
RIg8DoMMcbGZz3NygUUS8N3eK5NrW3qAIpMMJxJ7cNFr019vV+lZ8Gifl76+3oYP
5T3kDjat6TujRgkkFBYF6pUJ7kEwVhpu/8zaPQYmSQp+RoKuixahFyJSihzgEsk0
nI3ZuyffJUn6hBXneZBha/sT2rtfF9aESwsVpVeD3ud2eAq92auWlttzG5usExbB
Z/XrXJxVWUgGGxr/oO7c6mqg1ljfUKJK6Pk9gz/Ln4TSdIaNcinGyMAQtqSmgpHK
+J8iPYu98EQeLw/MVsrjT5IvTXa6ESk/vm9W5rNe1+w2RZVGTQUVcHrzKqd5IwKx
S3f4W61tbq/GqH/VWdDLrT8qFerwIitfp+rF+O3iQGtTeDpnhm5jDY9a6nslpCkC
ohxR3iLYNm4ccsC5SjBhAVUPHhvD1OU+FuyZm+JLlLPlubCccbfcekP9r63NFyag
JP0qKV6nl0mGcZOkPmZUR/I63HHuaA3NrKs73zEB/Us/6MXngx5c4gM6+wCbWjRz
ejGo817HZ9JkSFJUfkVwZa8ayG+wqrzBNRAnEwxGvQvqEI7W6/R7j0mblM+pvvo1
CFH+xquT6xbAuA59Ro68SWjec48KQaneJrIbMiasacKjvSRPAucJKG+2RkS86q4A
AxT5GwwJXZXGOmzllXiTXxw3JEqi4ZX+K03dp88KNFSxmoyc4ivu7eyA8ClmbaKH
qpDs2YVCs+dAXPWdsO1Jdq8m5Wml0UzonZMlZgV35vZ0anjpNNg/k5z/JqlhAoe6
ZUJa+hdsgIJbdg6SbfAd8eT657oW9ppDaKCmHz5goTGCaeatRdZikQhs3PXtimZO
zq33/vtVtcRGR8oFYlaZ/OLTVNsgPeDY3pq+4aEnSEX2iIzOVxzXRF7ghzzpsRFK
m4PcYDkGa1HP9Dp1DmxxFbmFrMI+6GJ6zTyKc67IL9sML1Z3K/qijw7jSSwxFIF1
shleFEP8ucKJxu3bDrpF7yBYY7LAcDlnO8b0E3BRveaMRy3oyddSmlHHUahadj0S
Iv6IJSDSplA9ZXOXkOxzDG50DtR5gx7zI9GhiQ4ujLkQK+tiXbpZhnIBBbKM6o9N
N2RYoHP33dOZSCSN9F8RL1qy3YROzYGHOvs1PZitJw8D4L0ft+R+vq02KA1KZgL3
ZCsFj2Qe/sgAXNbj9dEGySWhPBmSeAu7XadEdMsLLpH2U7BBF/75oy428g2mbIKM
F5eBTDn4GSoBaaObaoPPTmq6jmLR6sZFqzry9N7D9MxhOtOsb+aMFt/ZdhCj4E51
AhZBckzlOulASBMwqbciNQjCSvZ3G7yhw9kJrOahxcblGmC5dtlRfzoNPTgvRjCl
mi6IRhXWJ0eBI2BEpGLAeeNLmHWut5BqWiKvljj7nidCI42a7N5tcY4UAb2DGLju
1wfvyoQ0/gIuVqf7gg1tQLlRfJ8m5s6MvI585Xdfdt9A0ERFek6FtX0bnTz0vCox
ty5zXV6lyNCVGxMxxrxYnDsjXgUQJCpLqkzqdC0q+pa0wrRaHE2HKFSi3zEncN59
Owd2eF+fjjyYGppATc9coN498JGysvDAfEHzgsONxo5RmhG3fgLBXOgHQC9qO/FD
G1NKXKUyRb/mrcX2fyXxG36R4k1OS5j6ZgrJsgF3DKDYhO99p71/jgLwdNcUrDg9
Y7JsHEGjvuFfTqu7YPUmNJY/6gNYexTRmw8XB3yO/NcjTqQxlM5isHP7u9+VdprH
cWsGIrmB0vY56CxNybGK7L3aSvZHfVuOrJFSZ6FpKl/b8vp7e7LCDt394HX58VTs
jQ8RInzFHqPyFnUgam69d6k6KnlwObeXLwX5gN7AzQOxC0kBG25aZyj7uXIIjKTW
8nb8uDgTrsAEYMGULfZknh5JifaqAuc+194lTVqn6WXRsatNPcoryZ9YnzNM1f2V
9URg234Hrt6LZ4EJUlPNu1Ob8/0kiZq/l9VSEqT1MXjBgvHdKyuCtJXjMmjCf2iA
tUt6aW1pV42Y3hoN5pMOFgtU2QZcG/tpGcF1YMcOl7cJfnx/1QXFNj1DUCaPizL5
XeMKADtlYKNMWZS3FAH663pGVrbWE8BmUSIEyYHjPRN87D1R/3i19z9OuoGwJssD
5DKmPTapjLe71EECiq4BukMkKzw+GKjtVy684gqqq3k7878a4c+6qFRcP86riP6a
MCKh8WJaO77TJiDAJA5fxVmDJAbSlTBfncxwgtXupTA4O0UBQaNhWmAU6rVHLMRe
JwqNqzjppysbfqxrLC6QBe9gwQFmDq/TxXO6BrqLwNYb0A+WuZgyut5IFAJyLYSH
P3N2jqhUtCBj7n3hsd0sZYYGtQkmz0VibHehorFt33mZXwRlC/6FCy+9wKwCQ+vI
lDX9VDDCVttEl6GcckVghC21K8EHZ8tfQKwvo46LRScFaOYPAMu95lC9Xiffd3IL
0I/EKkNRWiO4kJ0H7U+fZ2JmY7P7LVYSxE1dwwOYYXApcXqQ6fnG4IHOoe3W4FmI
8si9wvFM7EZ1ikxzRFdezf9cvTpXpe1x08M2RrQxrXDwnKimaq2LlpaY5vKwmaMj
qlOSAdOOQyj3H/DLAo5nWH48GwClLvaDUFOoabADj5aTL4M5VxWIqABPTAVwU4Mj
jddWEZN8G4fqpgD5vKHOJEqDykYxOyx2Li6rsReMsaqVlKW2xNL/BGzBjzeHHGuV
MkHwVUTg4+X9CTLHym7NC8bJDaqjfePagztKT/bt/155wxD0+ULSJbvSDsDft+cZ
1VI9qbtormX76k0gk/IR8zrT/U2A1g0sY3e6ZexujiGoAKaCBdDbCuoelyfX7LBA
I20+hng3UKIB4mhmLA5UAn9jHF7Q89GxoVcwcRHi40Bw2X1mgC0pxPHBd6FQiycw
OuAcLupC5+OzB+olJnNiq9NYbj+ALwCB5hnCflmIj8hOWwjUEF97fWiV4HZdtaKh
eVoIixkYUYJxAK7HeZe3RbX5b3VojNzgJC0I9IYmjXWyr2J0IS5P1R14Vy/C/Qbu
Ov2Lbl5pmS+kmI66D9pZ1PZGlTvOcHKAPRMhPojLqOgI7bXqhVZTsg6bpacpBxhA
n6Ln7SbB1GTrl/GBQbHJmEEk/IzG2N9kJuOLi1gunJpMwoXQH67/F9dYOvCcD7sq
t6qC6n+rxtT/kCC7r5e+FfeqhNsce7fgjO7MrSoLk5qs78I4sFJl/nSE3GEaji3J
/5YwaDpaoMT7MM1fu1631XwQa4Fqzp0cGCaSQVzdFzgHkqz37SzO/JH0iezU9RFN
ReTvXnte3tTi6Dr7BsdRCxDN4rAlF29DKR7cJgRB2Qq6S8FQemsKfoeZ9wgbgTz7
VUbkhne3DHi73rbRXr4sA/acF00+koncMkibu53Nn+htpyY9c1XTeQyJ/LwxwQgy
fKEcSzIK1gmT8e28VHvU89tkiMWGJUothCZVf+ORnFatsdWfKU6ftPGV6pAEuq0G
eOUbVp1ML6gvFZaI7yHLAS0ABJ7gFzJP0D5kWrM8JDmJJ9hFdWJgGx/TCuyTktjI
ZT20Mz6GwWeuZTZF3Y52dHLmFN8zR14c9Zm7SRJTQuwsWIyKrWhhITV6eC0qj+mY
Kv6unv1f3IfPT6x+5M7CHOEkDp3jjKcKbZ4qDwcKvlI23o2HEX5YEUXQfQhjW0Hn
DtgKUpXEPYeoN3HtS8q68jE2qDxsdbpzgZUvvpU6CGebpXS2Gb6wouqIbMXqfUh8
7jEYfs4NTerK8l1WxRI6Vhst6dSLLsw/EmsPjTbTzr848HCe2H4igKTylXCUWooW
cj02ljHsw5DWzFbn7fUCjBFydsUVFNjmNWv1xWg39Rmckfo6+iUXvGecc+bBCMLU
SCgBqpR1yTBzRug7yhYUG9P8lkPcqnlpcSGwWoLlT6UDoHCuXffUXlIx8szy1nje
9bX3DPkqIsXNL2GIZyxayOBlwUUYlCe3lJ5FBLOlsWZf+CGGu8JBM7mWQKoq3AaB
CJ4X4caHFV8KMC7LFzLMLJOEoANJLrahm2sbJeYZDUr/AKiSAWX2eymBk5cyU4wl
woiAmvWMY0m7HyA11vsbZwQ5HBPXKvU47mdeHUBlmj5EuNU87WAD8uy25M51gly6
gfyHgxPW3vTfep/PzlCY4vUUyNWhp7ICyDJAGnE4VFU/f47CfBAbdam7+85OVxdG
2B2BK8bJyECzDQho3uXWfKc5hTZAgBi/V8Wj9zLsXFouh3+IpTidrcYPvl8yOz/6
Z95U+d3xmmhXXRYwwPUFi1zZlGQZke5EJlri/muGyD4ZAEJGM+215rVd7dzjvlHX
pl//Mow3h+Ujc1HIWvd+gVI2Akc403sWc0/0hrPLgwOIDpzANAG0sYZdP2z6MJVb
Ea1cMrZ+iPD6PCpWx1MRMwpIt8MqGWFXoWLE3ORKcNXrgWXRfP3GMBP34kBzj0KM
PbM/MykkYqPE823P4QX8k93fSCNMW6ZyPAvTSgdU9aAncGPOWaL1CqDUEHnrPI4L
QG6rjP7EVMzur2v1gvCOVX0N8lYPXCMmNGNopwBvGI+qKSk3+FP7b8yXcGXP1OVM
9jeRK+d1nK/KROD9nPwnRuW1nw8/kDzaQWjYJ5i6YgOu4VHZSCTV+ky656xK1TET
vCLepUCiALY5N4Sustare0KWPbgBMjSSJ3X59ARKXy/tS31myNbxY1qA+vVi2HxB
VKSsDpwG53Kl9898toURk2q2ZobEeyeas2/zgrX8vazgiQ15C1Nn6nju3A5h3PrW
nHUCl46vyJy+vkgxQ0MlfoHuQtvt5S/lZn6z+pDTupMp3ckuNfXxKADj8vlB5UZG
WFxhEHY56gc3ge/h6eB2Ou/w9Ds3Y/aq4xyF3fLR/MSCqRT/i1UfKu3wOi/1Ydr7
oUpdj3Lq+aMRDi0GUpcr4xujIj7VcYqPmPEryUq9qxokymFi9Kd96deeCiOGq3uK
RNKAxX27IkelyyVsGj5+Vr/HT51vSmqcMoHhamtR5tQC0Eb9yIyRz+RTNTUZwid6
ZoDvfc+KSKzG916mvyBkOgZsEjcvg/qZlXtgt0Awh4VgYeDvP8aF1MP+3fJ6+juY
STYHi62CX/1sfFAxmt6xcdSXj7Vk8vF5SQT5AsQf4LQ+i8KBwpVCxLP2+mHGicGb
cuWEeI2BlZSV9wpySuOCk2ismVpt2ieERwN8kciJI6EYc5PeIESWFtYRCtVwdFqZ
r8xmBwnrFOknR1L0dQCdgz11og/GGizDd+x2X65UI2dWdGTPRffLuo4qFTjDRbhB
bGReyNv/kCaCx9E1lIG5TjM4EPxFPVGy1NEns6mvkXxxQcrJAsd8sv4RsRzf9x5Y
FqV3ZJmTSxs9r1cLXKEOioBZtImVsHF918OK6lrXo0s/Z9DEQpYGKHQ0YhX6E9ft
n0C9MxfjUUQrzo3yGpGxhNSa2DOKMCP/Q9O9V995mU+GuertBaEEE8kI8fc8Eidd
MjeBqhS7YMIKv39ghURfDaZWU/PcBre3hfHpZ42nLbwzjS3i/t7yXaWfU9l9oU/K
mPqhBE+iFIs4x+5SaiXfUY2R+2SLZFbMeL6+hyx49GJwVaegTYE1ZKcsJnlMR0dQ
F4NHRBnUAv4kD4EZdHBfTH4lsbIdv33nhs2Ac6alZ4dLC2lRZzFXGrnej85m4H4J
2WWu3gsLEb7M8Gm0QTBeqwIAIBrYHvMIXeljINGvraffmdPPnVHwu/2yN2UMeTvs
j8a3XCDzd0DgTKUDhfnh22q/Rswxlw4LMVx2IrKW2gMROS3roW+/pYxE3o+QJato
Wbk/f8hBj7dqvvcg7WYshhyWpJj4ekeZUva15qZE6kWiPLBNMpSwzyOdB8KaA8oX
Q6aDgLLMF5107S1axaDKPGeipjwmEjMFcaqELN6YrrGFOOCGohAoWpnpmkH+ZrLa
I+dzxD3l4iXkvcQsBjnpl1nEWabDWK/dSpcAeVxMDqZUfN8y9YM3+HKKRGzeYj2y
TFE+7lYCkAdNE08bcPht/5jVLdJOBxt/Z132xDmRiMUSoxgwVDl09Gs+XzWfduSv
6Q6zZudf/uzKvsJU2LiWbQNjpUGbgAQszW4Mroa6LsLwv4I6ej2Vo8TNPt75VBq0
cp4HWYYJSe8/gWrkqjSrHpOI+qt331LyOoy312kyeNunjXGk2UVQbiIflc0zo2KE
ICSAnTFRmWbrgWVsjwZTJaR2cKDPFV4A4asfMZ2zhi/j0/po3ARpC7OfAGKK7seX
EY9E2xRsxRAAk33srgib0ft08wi+vdUM5YXmpayz6HZsjFZilJ6o/tRSmmDGpert
sYXiclKKLnqa3HSRmpvEz9wXECvR1arNgMhHebWx7Ssof7WoAziOSOnt3xRpJ8HW
Ec6guI4ky5CVRM5KkYxiNa9vIatE3yY8v/kVsbzjN32RO2eRXXRML4EieF3KvisZ
jd6+7k0JsyIlHENVZKGk22nCupki5bYGUhG2Zx/amhADc/uavt9UE38AuusiPqHT
kC/qxDMRM9+PRwIhB+UZ/SenOU+zl7noJJUwB0GohMGhAr8+ncuwrXEs8S6YNV8A
QvTFM3Zj/jDWyXDe984PIWLqHLaGNMHe3+4qUusWxpdtz0qzsLZ6i/ErnfG0Cn34
qkpMxyIEiDQq1tDSXXjCR+qXYttRcjMVw0I3X83ouKKhVcMDYKhbSfOMZy4KKLqo
TCtPSDa5irlNM0BhcBOYBDSBEaVGoWpmK9sJFkpLFOhi7OLp91EW+U6xz2V8TUQb
sd8aG+rdq+cBuqxCWOKV5nYDq1cdhx48Sz78Z5mlLTy9/j68FkRz+nMJfT55pDpj
I8ron+mb+NqjhLZ69foIL7jP8k+G1z8Dv8MSE3Zy27xdqLdNDaiBDCNtOx+H0ovz
dbR4HNe/bCQQSfbm1edK9u6RBc4437URzA7cxtoh7XrzROC5BnRTvv3irpmvP993
AnLKixQ//RSsHQ4p2RztvfUs2akMkqP0eTzpw/aCRcSam4EaDGR+KSZ4QsIwWAUv
jitXHcI74xeDiRcSF/XKnlzJHYvqjRoWg5Qs4yYBuXRjtRG3m6I3l3HeHLLEK1Pq
SmyyfNgSTj816AgR+JLiNyVA40DWFbqCgtc1RPnSGJF42e4yACLhtIoNY1uRuWvd
hMEsrUdEH1QM1ebdInHA30BJjycB+yLHxBhLq11uyckuD/WwruPYqs3k9Pegg3LG
dg+rmQ7WGenF3X5EMwOQd7x01qW6TmF2ojbt4T/n9F/l6zQRJqtVOR425EEoOIUQ
s8GYTeUsXSISlfkGXPkRGhxdalR2G8uA2M0GtaSsPqaIoVftkViTn8p1Wh2qBlxT
PsX0HT3ADeGE84R8gMWENHCyCb4vMe+R2SstcmF/M8KqtjIUYExuEDJxjpKzJfC9
wFLdxj6hZSojRNrXJNpetmIlkQEfEN8LGzv5nKjf+0KSeGvFNbB2oWQaGk9qgrnY
nV01V9aBmBZUm48yBm0RZDniYKu2LJ3F+YUflYUu3tPXW5+LqA06ojWdos4aQoRv
Fj5RnHepEu+w6Nc45v+pMAY4UH42EV0F5eAMzxC8KcY9S84Sf7TeQ495z1D7m6kK
bscZWMev7PDCRfiDDdDPHguSLwgOugffg04ViG5mlqkpzrPA8s1zZsakYdc2wFaY
lcNDPiRa2ct7HHN11it8v9I2jWuosTlpbv41Mb4KsyDUMD8pUCUBRyMwhqUSN+Fw
B2JlU6dp72Gkd7A5d60aTDCgrjdEuvXMmwcQt6PF489wT+3RPj8MULhQKce3E8JT
7p67AWzo9pNFXoWVf2Dca4XTghuwUg33rPrIY4UtkKBgSzvPehPWdN8uV+iAAepy
NC7OaASVCHGD3C/8PazVfVkySTpNeDiitVdzkgYdXC8A4zaicjaEFH2VfUlY9msv
lHmATqy2HuaZcB4QZaZ+c0eYNK/RVw2RoB3RMzsokFMawr/z5RQPlf2wXfAwEUGJ
blPUuV2UFvzqhMGWCxYyMzxSnO8Hb46Kp28CFGqGPdrTXalu5YOax0X2JfC47YMt
lBBQLu4HZ8np8EaIjw7Au+ZPCbs3J89phVwkZ+4R3bnLEsfKKYswMeLRxnkjr8J3
QxjikW1aR7MrzgyDrzi5Sg+Bha005zXdHuSxpCwwI+IzG5+rfW1+mXIK1qtejLcL
QUnVVsvGFxENGNasWN09e5NJZFB9bSfLFS3B2bpqHnFmI6daAFgKINXkoO8cf0jp
Z/Ne3ci8F8QkBl9FeIUTU82eARkg87cJDrGtvvMGEgO1Es5hVikhpTNDOJcoQudO
C1RMGPtATZX5eHC+jlQwm8ouFu/WQagVLwnqz44oVKSA1s9TD2jxT8yqO/PAgqOs
64kY5YYawmZrzZECe6Bv6UjOXCgb3QAAmYXR/ELkwdtWQjeElWoFGzjLZA7c7Zl4
4XLPxKKLZ7PTpkCmgP14yMFyHorxsOzEckdvul/OD9MgPSSe58C5WfqLHGFK9Y7b
ixdPaJDcL2QAabKP90BpGWUqLxwEUVc5+SzMMSqsdW/k0ppuFhyGo/4NEuf5I7ee
gEvAzJgNW0/UI2B7vQZj7NW0ZCPHKcaFz/WeFdiqE9ZK0JGRnmoh2STM+TF74kAX
uuL1nz5WZNO5bW2Z6Od6d1SRmCqpz4jMKOJD3bDJ8Ruob3DTRdjp6vTgVrVt5Acf
fRL/jGKh0PpkG294blGJQTdau3mZOoqUElG25eOqRmkajA0/sYyFqAc96oIF577x
REIY69qgHLKVqrZoWnWb0Z3um6nQTcARw7jZGGDbhcka5tolim6hemPpr4+21mFj
CATkOLRszNeMwb+A3hX969g/7Lx98iEZ0p3DkORsxbw9ZDQuoUR6QmDor6wOSuT6
Z1U+qww+kRMYvV85sx/2SlktBxq31eQdQplw+jXrLJWu/i/wPfielcUhpbULKe/V
r6Zfv38GqULrhTmqJGI8EtIqhzOOB52N83utZAKHFsekBWBRPF8LUAREd3e6FCnK
uhUDqgfmjUns5dU0mTBQoxj/T17utLDCqbXlZJGP+9g7kOe6djaUl6oK/AjDeSkq
p+ESWwZZO7ChbCn6d+SL9Q7/w5RpVAPpTBNxK9CFq2CSKW1BC3X55yt6SiGHuB9o
MbJZAA1DmshVhLhFntfN3nZiTwlWdpPME1NEVQMJXvU3+XjvUUYt4UDco49fWfBx
vZkJxelBSjueGL1BUCSZ4NeDGf9ILSJgxuLigrx3a7Ojm27uegSBtKCe6l0CtYiG
IdAbL6Dkuf6qoZYI21x9jhMGZQyUjTBqw/ICLDoaN13CvkvQm9Ckf+uKzlbj94XR
EjYjyAtIvfpIGFey3k7s2dqFKybhhLpFQ+8jTrnlvg67x9C6IKufKrFhKlYmUzCH
zsOrXbzDN4JgDtofNjnN9I6ZTgms97VUgz2xOgjLO4M06t52vhmOuPUO2O+IhI+w
LqN+FO0/Sj97uzAIpj0gZ/tZkIHWHDLc/4ZDMGp1lEgwrezD+eu7bItcqMg1bgq2
ijjaHjYWdAwLX62Prc1mE3z3I16qiIu00CXUwb3/afe2uIkrHqmjhvXwF2W6VZf7
0KGSr1lv8CTEEi5f3mISacjJo9KVvtDZ8ox9XHlttkwsNQRYUrGv5Q/ZfUOayE3f
EUpBm+Ft8C0v0KlY8Sd07GJSyOJkPIpiakXDaJRk8FadShh+UwazDZsYyGK2XvKQ
Bol3iyCoAoM6OKxUR6+qZs5NRL8IHlHZ2057fuJPuF4SCCEOVpbm0WPFcyRjINjm
wMb6PijXeE696NBU/zI5qNXd1rQwV+ZnTDuJHzpKd3jzMXJ1jrx//ExSxYFsUPul
D4r1u9dOnXiF3+2lBgLOS7yfBcz6poPh8g0RwlUm5VJmEfTYN0/y7w0/U57Uu50i
sFLNz4pNlWL46bmajIVwhdKGXx/MnsM8pQwTQca75ilzBOn7tln2EuOZcu2vAxk5
sQIrQu3JfxW4M41CQBDEbYIt68a9Pb5PdqhKOeppe6SbvIFHMbMjEJwWBjImMJ5B
mIKaW950ePMK8fD3sG8AlgftpuLDpuhqYosTZysDcs7zVJhgvbblitmP+v03d2kh
BgO8ser3W+87nX9Xv9jmPjE8s8PgyTt5Mwu6HXFkznRsGoMZ/i/Bd9HJwJj7AhVL
OSQiwk42FLiOfLWAa6vSR5l3BE5zX38aBHlXGaVIcgMjgZzVRrq0kHteEQlVXHXu
c+nlTpaLhHPcJFIp4GLzAU8/DJsWFsfntYAsuxGYdx9dHB/JVpQPLM57Tso/Rd4g
bJCidJAT1DHogzcG1b5RGjRTHkwUKTHjpnkO5st6TBXi2adiVsHYMmY8wDhcuVSl
h0Zf/gQ6WwYu3QxbNKp/78D9KKufx5LXw0XdCOP6KCtK5lfn/nglwNMJf19xIV93
ohodLQuD2N6JN34qOdXk2OMts+RxE7jOnv2VOc5JI4I3EgL4kHZmyEOWsfNJUgfb
AttFr0zMx0KVfHefFXqSDfanP/L27hWFpt6LP+cOus8Xnx4VrypTL4ErENirdZO6
cJkUoaqQyxKwN2aKRxqzyXvrqEqGU+SwQPoBJdig41+IVONUDoCerMeVlsSw2FFP
/DWCwJdw78Jn76b8gMJU0bWK096OS3LnghamVi/oJ8miZ3OxlVXpYTJ4jUNSKOzd
Kwziek9KyYSGNjuJ6xvsY7qOg13rg9revQjccgwpIovFfkQ8SLXFi6aIoLP0aqcO
YBlNS3mNdAbz7PhNcwUJct7ORxMZqFwtl1WZDgKrTfqJ+LwY6HRNjFZ1okxqEqz9
p5cwl74k52R0R6EFmfjGYjFWtmz8BLxSv7Xe3yK/wBsl1udE1nHlVCaEPHjq2m7K
agzRV/T+f/6Kx1Ymbp3E0nLp/3Vn37onWOFiaXQ69xX/oc1jywMzjLfU7v1HQ1Ha
9zKo3MGH0D4bftBmUdVrcRQeAV2O70hzXeMoMLmQGgwSwPt109zjah5Mn/bqZM4t
TRgKy5614rKlylp88AHTi2Zl8FNprTku4OCsrM0GmPyqPpdcNF3uQd59SzlA8og1
YBUyivq3wCZYUXGLCIFrGc8kwOTM7e3BRjBcKv8Exy8vFw4RnDzrHK+XR38arbUJ
OsA3Sa0nUJg2UeoABdcfMGa4DBV8TD0fSNGfbYyyrXJwXoIcpRJGEfm2KPpRI4E7
dO+MSsIq51+PlGRbtWwjxqhN7me6MZNYBrbLkfCsf/JvEBcg3ZXWA1TvqhknDvwE
UP9Z273r5Lb15eQE2iArQq+WKicRthmY29RoUkO4xfB+hQKIOcbH3p2h3oyRH/UH
mADqewx6JHiYArpZK4JRwydFI89948WyWcEoVYxGRhjWgxW3kzetn1C2897Fr1fB
u8DnN68MOPelLfzICSNwkhFSKhvJrT1WhzY2iQZfzxZ3fjPGuFkTDPFWm8c0mqkx
IsUIsyClh95FOZ8w8e86pTECpw14r5glFmwVUSfNgwXEayGQM6gxg4t9yURkPWjS
jIDv1/9dMJbKD24UeTfnm+5z7ggD+TGJ5/arwl2aXNCw6hHV7QMgPhtzuozjWb7S
s1koQFAbX5p8itqn3pJByIADyIeh2ygX+LAYVAlX2nt0Re3O+SKM4zPYjEeG/Gax
EvOOdLCLJGYlL+dTB8+5IpYwTqTb1L7Z9DzgdbahcSXlPBp6izyRqeY7hcC02JBw
kwambOrnYfEPWedzZ8sGbeqSvr7iqQ78nr2A1uBJO15m/EiBjO027UP3HSz8mGTD
3Wqr50o6lsfHr7q9PJgZRUbzDPy2ELAeDBmat1Bd2NZuCr6H6040kRsdeM6RIkGr
M9EKS2klnABYZKRKdEL9zmw+OUnOv5qlt/UcTZvworMjfBZsefklleuWB8jTQe23
aAqtOB8Ucvkgo8KN0iZwcG2lENeAE1tYHsZcP/AgobVPkZ3ysJqK6mehft5f262W
ECVfHKS/uOA/PccLw57jjySZIN1mJ5Ids1KoFyl9iojkKLBqo//8XYhY+Ohz69+P
sXHjehjL2WFzh5upptm9BMaTdOHcZYyIzHVHDRIxOQ85WYMIUrK5zYHIS/nfUsFg
foul5lsyYfjBgcxU8fII/T2Uc9bWRB8N5HPZSCrTBm2mcS7QNV5/hLrFPAOHDbGe
06vN0ItZbYhxzrypaPd6AWWoM3/sPCnzreWlmWGZCDgu416JzXsfkCU4nkrqbUhq
7KYhwUYpJ9v/EMzWo7zyZijx4TEgO1UxY/im6jc9q3k2Lb6y1cHuQZHWL7RAZhVI
cIDAidHrLHu0eoxOWDUgOxG7kucOvkrKO2RSUJBTuyx5c/uBCxCsNheP20JvWB25
/JvL3+n0m5oP1MQBhhOV96iRyjRBWnnbY6TSOmva/lGFOd9DXJXWyMnkMLASa4Cf
D87ZFCR8UfnTbWWeDmpA5iBOV6h251mBnvTnPJPxD+GtzaLZc82+CvqTMCOF3PFe
TeMs4g/hHQBhTq+VNQJxypOsiRNdZr7DTilqcRGifOAJbjQvrxTfdyTFyBlXVgwD
gY5KpeeKhqRZgLMkesOiXwk3DUZ3PSTd3lCSnVBoX6tzgMgQyHdxnh5fIDsRvr1Y
o6Ly5831Q3BEJKULTusgmID8Z1mkj1OKga1DLoMRLeqiGheqfmCPlW12ze7AMsdv
vU4t2E3I4Bwl4iWb2UDaJCdJFWRxVT3Ro7sQxhJrbRZxhB331is7AR2K3RXbzPHG
iEI16nDANhruwnZuF5PuvLawHCKupgtfyL0+x+8pMBikr418FG139mgaVtiMJIc0
zgHJ0p7WWDCZeUZcHfQw1rH3BWjEAKcVoSZf+JX7JBtktqWZAjnxIsLVcjJE+eta
l+FYV5VErvTLGg020muBSIkG1pTd7KX1EzQhy0AV7gU0AducQFXrf6+dJomxt6Dr
e70U980uIMXnHwJdgW6QVLzMLfLAeY9YwaNlpNjHdQhd60oOnSJ37H9SwEd1FSfL
rCSKBfvtlyv4WRjUDxuXJdXmNAIlOOPARQ4Dw1ahhB2CUT84DfCa8topugpi9mlG
TwkhTmlotMTZYMcNgYYSPjxBJ3VeC55jEB982871EFcm3Z5+kOdsrx4sUCdSOvD4
6wFJI28FLuz4B70+PU07X55QU/nSMK8wG8VfXxP/PjCC4xBGNPYooaOA2fOcpt+n
1liNj2wALjv9OMoHBMS16S8hPT+V/5NNQd/WK/Kgs3Jv93nit8mAqCCxHIchfLzl
IVoxvGgg+sse/KPlMwI+4ythn5InTwZwjFR9lYEy+LtG1HvFMsSC0+W5Gi/b/uO9
QSSF278Yglg29tsQmgz8+c9G4FIBKz6cvYaaYFwYdmHBbCg2g/ZQUv9u4J7kyx1p
zHVbUeCsAn6gNjIeT2RxfjKm11g9As5VHEyBSxnRQJqx7ALKy6GWeM3EALwTyTl5
MS4Swc2JZvHHiwEY/qARLny07FMeofbUwshdtSgWn2jTcjmuXtGb3r9+6iceTJOx
2eQcLcMLvI3gsgHICCCRG1FwYXnO9ujfey2LNCBrrwCk3kE0ZdDLxD63K7fEfMvp
J8rkzFnWT3V5pZOCfcAuF1fBHtm/eIVjDO/+7NJhpmu+uS3cpCuhqWZCH6GZv2bW
nJ4HnUs69QmZi65dUiWCnCZg3xgA7V54D8Xbj/zkF0bAJ/XEDmLFIIrgDkaKQqVA
7F/qNaN8TfwJ6KeWUPUbyz9hwVnj/QcoRe7/8Y0qmqpYLe0L232l/xrEmVNZd1o1
oHb9eylFUPVoBaLs8BaGqL4FWTfADF0kWMWp+WUaZycRM2IBLri3UjMbGY+KL1bO
t2BMlZvDSbefqOLy+MLuk2RjqeBl9igUa6GHAc5tXpPBH+uBEb04TLiRngw7aPBv
lM8E15aWnHTrKSzDwkdVJSAajjn1QJZMpXApqabLoz/vFqFId3JWbN3imVY6s1IS
zSGfsSFby+Y1RE2cQC4/BahXqydGPvkXDjUIXr7WGLBIfMv+/oigf1lVy5JiqAdO
zeh0eTkpQXm59wDu1uwebLxgQntnTkNjckDSGuTvnL7U6WKqgoSzvPKkEES80623
qtUT/1ohuvvw1IHwM+GYMuG2ofOyXj7LADj3TxZOICSWF68MSDDpRr6T1k16f8Fi
Fl0VyBoWqDe99kIFvMh194Dq2f4neudNP0e3t15QyIrA0hCnGIlDt6i8GK9miowB
LyC75Jg1qPUG8RsBKJnnFLNgJbjPjvPEtq4Tj4b6ck6qlYEZNuIsq3lFoYqzvTcC
jaxxergR0/APj5RHRwhX3uacsA/GQtqZYG+T8Own5SuuRpkeH5gcfNleAORp6XLB
s0dQ2S+KZ2lpU/t+ecxDbTtEIgCYnd60di0uJixURNBsoSaHciIyfcI71EsQAzHj
KNlBeh0jePFPJOEHGewpKhV56fpGLKkiP2k6sLLW35JA+SjO3JQLTkECORoQfEzO
CJw1i7DR2l3DWPeU+SOqsLQ+WayoY4FyjicZ7LqFLc1CqwhVDkQs6PY6u9hjp1Uu
TsYXdRCKKG7gggCOR/He9ApAGJkruttyQPfrpLoC270/5tNVmjW3G3mFQvWdqEul
3i88ZxxsnH2US2kwg/LjIoqRJNiC8MEfZXU5Z5DzU2PMrEQNjOjmUcQ+FWDl0jU5
9xu0GJnGuuF9sn4VjJop6fhi0OcZ44pQdZvcOxC6qzOKJkmfCMo84lSMFxER+exN
3SQy10CzDdKXjG1c/IHksLpZO2VXhMOMdH9TIZ6RxwfE3rnU5QJsgN5d6CFChEPZ
Qb0rGIj79JhS7v0ABM5tGvSy0xWmRq9fB9aW4O9a4fhtYSwoS07vvPd/vXnit70o
DeevxfwjZ/Z6M0WgBjSNl2zrRGaTr84AcNvVg4FVInpMqcgUHXIitlOFXT2pQNzE
ch2f01Rxi50n2hDaEDnK0cSfXY1RJe0yC3AOSfRSbDHlFW++7jmiXsMZg+9JhgPL
D7kH3ooCu8rk/rEUQhKKLONZ8ehsXyWZK7uO4HBvXjfjX+yBpNOxL9wqcccJuTO2
NK+gxCDzJa8kVdcrU/i3WfO85plwzplQzSYAJBdHSqqzWNox38rgtp131EHWkxJ+
jRjMgSULYXyGqlluzJYnbRhXck8DjQZUwDTS+qWrFE2Gkzq8abKUS/WZ1FY3diKH
VDxpd6R5Z3wBEBljIYIBPemXBY9DeGYKh+Pk7U75UhTRUsxifDaF5wwkgXPfSUrY
Ma7VKtUuepaFf5nRjmhTNUKshU+Vz9r1Wr1HItCgu4Q8AcsQZLZZig51lYhqJqdJ
TXGZwLDqIVQpNX9vNallvGqOwS9a144wbr5Habi+baPpKsgCftCbgbhq/PIrzePZ
Q9yiFH686XwPZPYfF70ByyxaiLI5tNsFR7fkcDty8xXzLvoDwsKPvUpTL9MOVdX9
k5xkO9DWRgSXsJRCuApP/wIC90qVTNcnL/6VnOHj0Vn1XJYM2QnsQ2lT48ylOXrf
1gWgV4AqJuHst9DXVKcU/Pj9BL28WveXyf8zKAzsZV8SQpZrw/K90MsIL11V0l0X
cArIdA82bx1FtCG/sDCLnc1IVF/LULHiG7F67owatgrs2p9Z7heOIAx+b3r1X0Sx
SzTpQMm+HDUBoKXFKo83+EsYb6cXjBa0/aQ51ADgjpxExj4MlzeCR3QW+egrRk7q
a5gYtdXs6GnGNdAbnDpFHeeWJnznw86E9I+b8bWWzoILalVsLOJ1giF2rIRL9PjU
JYAZyaEPO4MT4M/QNYIeVFttrDP2pseEgwWnZbaUfi6ey9zH4cd7ysfwQtNkoeQI
N5VqtFjLuOJwjtrUn1VmqI++GseLTc+HGr+6WdubZm8jr7gL9ZGUHB56K2I0Ni22
vg1y3hx6ogQGb98VErvrRZW/Log6GGZYaI49Zuf9Iyx7x12MtH4VjjwfJO2it8gW
DR5vKj3raD7VkZVJPUm2v9MjolKWICm2FYAZ7iIZpOLx1ij46ra6mb12vSfHbMeS
2M2aEowKumVsRcMUirxCe5sInIKK5VHoLqVnz4LCgGpB6eXnuKOAHHA/cn03njdz
Nib0GJG0jXPcHz0xbN3gkKS9BVctcSqpk+QauAmMazHImZ2r4DB6KjqwdfZNf+u+
R5pMqpE1PE7Yc3IgmQ5kABserwfNG1QQCT6Xjvqlnsl41/Rge2/vZm+74sCw93VC
vXwmDfp+zKYZAOnR2PvHm6T/rFUgUf0FO97SgEuVcWbaHXPyJnyRt4dH08TLpyib
kJOaH1FulqZ3ytHR2tznYkmUvqV+LvLx8EjKp8vXBY8n8Wv9Ex+VGYWHiBIF9JuL
9NOwGT5slHK8y0tJyrubpQPFW9azZ9O7q2hgBXaS0paTkb0KpOCOvsHrt0gSlsam
L0/BeNGHTJQRZWa2vLsHIUx5d/paOLg5Qqbi6bJ2pKiOqIhi/e016BmMFb/geryT
gxh8+EabfkDZpiUtPfH9cXyxq+psLbB4ovbtC/g7Y8qDBtl9Mvnba/soiBcKiqO9
/HepHmMPx8t6yd/Ozs/hn4m9eVBJSZLeX2aYNWTnKKKHrzGyxIxQ5QAorNT3+DgL
VFVLBy1YG/dXos0XLZPej/eUZs3SZ8stHsFSYVGt5SjNfzbtrJ5KJLqKxrKk/U6n
Qy5U35rvtfpeRZQrn7rbOYhbMQayGlBBosRveuo72E8wBBTWb089Nllw34x7Ultn
CSAubRIySh/Jd5OcGd88Os4/q8n2veFFevG7QPXVAyM/RcyGNESt0czTy8kHtcF7
Lwrh5wdBnY7c9Fz14krz4Hvaiyl8qL3AAAVogjjA9S5rmPlw/9mhUc9KkS0t0T8u
UpPXW4eT7eMSevgszVOKcBxlco72HS5661YBZ+OQdllsBH+Qyfeb769S2fOM8oQ0
d4Bc/ZJvh6maLZgTuwHOX82bedtVei/G3mDIgK7lGDyEa8aOA5RnDN9JgWaufVZN
uiNbbV4arFcVgDqO99PHKw1yvpDk1mOGTliiQmYd5LMYp6J9DIAU+tUB2i1Qtjru
SfzhZZRCIDMqYvjClLDFhVgCZsSCzfpb83uKmFYex6v3zWo+YLQzK4bgY1NxAND8
YoFtEuOFQo9uFdA3Fca2JjA5O3gY6Kdp2gzZNr5+fWkBApscO6vmf3C+ZbBA7mfs
ubHerXsIladDi1KodTn3jPv4AI/blAj/EM3gBGh9veHD1DjmAYPoWzsLpduKRGWW
5eZ/MPS/ITfEtL0mlQ3JGcee7C4MhcWqEYxkGdYOBVJWSPzeNX2x6/lf21s/n5lS
TuhdTaQ88k8f93uPS7uRdzfHxWrsLMnX1Iu5Q9fSQmuk+FIjFt73gR3ZmF9Okht/
zn+bPwbxMY50GBwa9SkGYqhxFiba/L9PpsnyPrP8C8qBj2vj5rGDnThFscQMwK2d
qXfS8oNUDCJX4VTix0uPS3lK+bXzGoLMr7yhGo8VD0RLUBX5zkGoamSIMk6hmjZ5
2Z4WolkD+Hg3k0KsmR1gLBX/rRnCmDDqCGBajvhpkj4XAEsP313W81RhWDJLTSzw
FcS7QFc1FdCj4vV9zVima9sDAybDQGyknME4tVKAecpgaG2FnPNgL3NtLSvvl5++
rCzQuuE41W61oXWPB6jGz7H3wUNy9vI9nBs3xla/sCfiXcbCQbRMHYWL4ePF4P5z
jfboJfH7im9qEohTmOfI+7dnEI173MZWr5rNaSv9KRBzv9nyT8XULGiG0eM44LyA
YYO5iOWgCPHJrOTFxlckaq/JxdxnnrzbKM2Xh+VF6olm4HRvxNXDb9EZm5bBoJqi
YvO2mvS5sDupwDihJum3fZQpkD+TMwiKSXaBWJ2IcFED7bLiuCz5Lm5vI5wxbgnT
Kpx+CrwpRnC4UhS6mpmpm7FZsySMFUSndc3eHIoDE7bBgYCQbe3s3w1HQB2mbMUw
prd1TU6/TTNBO1xkq+2DqKoSQQ0Hm0+JwvODuHVwMdU2yu0txIHDgMCRRIIU1Fbr
wXinEex5+zR0SCtVqdHbPpePcmlaQeYeLznP8TTJl6wcaJE/SFGlzclUjOTUFqN8
p89GGzc5F4nm5FmT/v/SfP2nsHeIsR6PtL2tcXeFS5PqmGg1LNmpEe6pVUhjqUwZ
tmXbhb5IR1Qge/i7slXFFYgnekw+57Sdb78XAXh5Q97SgGrUkvcMB97SLCRSf80X
DYSK7Lxn5eP06AhC1YZ61gkmNIwpIPNHchh9sF/wlKSoGabe9Wq4EX5PlFssLNvO
d+XafZ+mu/zahrN59XNGpyYmP/w8UCkWv72kxz+8qIMgJiYFBEqHmMxp0oc1ZwRm
LZVaQmq+8mNTP9gXQWRxUvjOnhB/mXu4bV5ORdjPBuLCtj3f6Iw+CWKD8T+75Sa8
l8yN5LlWmLiZV2LHE6H2X9sAl67cAcsUj1OWhHagng9dqkEz+RqA0iNjAjlp/W5S
AUgT2w++a3mMbIVcqro12ilvUyKDwZxuWjroe3ju3m5chdi9AxTolkHWcP1L7Jwn
HGPNV4cEB8HYcVWQAXN6fk5cHeceEPVUaFMbQ5LcrB3JV5lOIYom1ZHiiC3xAJG3
GQOM5JukD3XOpsm829dZjmA/LItUs82u6RKLY0BRlZzkaWRLgUr6LUesEbyudA9D
XRzd/ssu/4FIcjCElhp/SCIUP2rsttnxiIRcGSOv6I0eBqz1JUn7GqOqi3ccFJ9J
n/3rSax8oJfqCN7e6fiit1GmveTuDg6YKuzrEn7eGnZ8ZaPFuyWSeckYZQvCTc3j
7u/aENzwiao/O1XcAs7ltSWMiqP+5cbqLseVztZWEpoWJP3lBmoVmfOYaEDsaXKv
RjcnG77ymM8zAXKgMobrUbOga3+2VgaTNt7hp4izce0Ncx5V3pPYk9JDIzAVnYEr
ZW+8AF68Q91uXJdMdqwQ4vL+V0bu9IOTxLtruRqPa+VUAn8Mi7Ix71iTil+ckSmJ
e+wdQQ+pXYGnPxacjwlIlTB96evib0bFpLF/1CaB1FIzU3mNABwOtwRrmM9Po+zR
Bray3IKGfHwSgBCH6/0cB6PdlyerQ+Ivm+pa5t6tmsPc5/qr3XDB1cguQomccZG6
1DNloBAi/8aZj0gLiWF+yhvhp2/qS2rG9fL0+R4U7ytiAqb5l2XJ2eOhkbsFy3AL
zTXWRbl9tol5mS20vsQ5SY8bpcWD+6k/Gk8c31qBCBRfcIzcueTVwnfk44etddnm
jhu9z0GGsJWrzeCm+r5V5ckCSKMe/etkRzpCIbwBPPPWfEePmP7ASJaYKUX4OqYi
nvubTgYPbGUl3BkB+wC7TlVrSCFhicsobG7TT7lXNQBXAhF9xL04hoJjMcxacZMN
P9mbptauywHes8qDs+cgFEvaRa1YVN8Y3PcB1bMckUzO1YAKiZ9Q+6gaFJvJSawL
8IsgHJFbYVpI6yRLiDxaRHTFWQcTExhh96U61JLTpLUXOjIFELKHFJXO963qMg6N
oNBd6u/vhk6MHzNrhe1axL+GN4rcY0KMPgZHH+t+LWFqR9wLgDC/L/M8YPP5WA7m
M9GlIrWsXdsmRkZZvi2PputVTFgHlUUNNmktJWYFXRcyfQdiNyOWgx7gZb9EGM14
5+YHst8OmJT0AnKBSx1HxUFHfUW6YVBO+EUW+gByCRwvQalMx5hlyq1xs/mnfL5z
KUbIZUblDOaS/v9XRTKU3IRkNihG9ir4yPSiX2iMG/R4qMv5+OtcXRlTlF7MK3s7
QPtvCL6h9PcBrS1iENFAPNjrgNpmEbuasEsdk5vhfNExEyC969grx4uDex8YDuqA
XeAzfUou4ZZ6+MDfYpEvzRMQx8D/2R9sydCSJa2GA1dPhOSY8N2PXdbOP1kCMqme
GlJJOT3qxVpvJA72jfBUk3MpLQ8PL+82KwM1eyG0Fp/6+LJIHo4ps3OGehleTuie
DlJFLWMA7qAzRpndlt8UpAl3xwBCI66fh2eKw10BkaOS8WJKKW4O662C563IULCW
lfPwSNsiqXn2AKZQesqu1d204C08VGzAJJzVt8+21jdChygHxCt738dYNhuhx2GX
SmfFxpSTAMfcIef3vU4mHWiKMIkXhDL6ib/3RTq2Fh6WXtZCBleUmP9iOSW4UGTb
UWEXGhDWf0kCTsQbZXJGni09EI8oQrYQpqkw5yQ1DcGjLR5hxbo3OAm5lTB84W3R
2jabr9CSwl/vvUsM97h56T0yxqew6qH4RLkcRb7VdLoNp5kGVPxqhRsITdXiCYRc
8eSdqGpcEcq3Zfb74xaN2ydlJyvFPnM2DbqkEGaB/hsZF6fyvSblFlFSSIhDGVng
kZWMwiB60BV2KsSzH+imyREMGqrGKM7avWo3iiZhGd4e89sAeL9WL0r9WpkorcGj
Fl/52GLne4QwvJBKnTN1XY8yuNGGX/ecGlKpE4oJLy5u6lga5tdm0ObBGD6Jfdf3
F1ZAO+c72KQ0HiRQMaEOpUeG8RSBhIqljkIyF/i9gSOj9gWbrfa9OLUwtnF2Cfwp
beFu1bwT44C/mMzwkL94Rfdu4GVn1R6mgO2WA7DQzLVY8dt3ox+oIf/eXAOJsK8C
o2hxdKAQAtCAYSayS1tHgVNudKxmn4DgEP9HpD7BGv9l1QiQjQekKOKrsQ19x428
3x8TBcQ872HV9VosEGI6akRbmHBTLxe3JI+wJiSGVJpuPhz9uZMCCHVTl9vvI51P
dEIsZ7wsFPHQXFMNrmYCGwuf4wTSQ8c686151Mq/FYAHhwH/TVYNjMQCLEs5+Lr9
GrrdjEC6tkwRc1eWV8FPPVbCrenxN5TxvssKhESPfuQZPovz/9mNVlPYdZ7jCD+c
WqAzbPQcmr432U3a9V7uGBYAMjo6EEhl4/r1jEnXc3fPdVZz5N7ZUQj4czbpwT3P
HC6w7IGe68bmCeGpEdJLYdZZE1XdVGBfYQr9SRYp4OfuNsyTsumqxaFmMw2PzzIT
w5BW5rN1poAl33nM6fr2iUnvMnOHouGyjR+qCRK2mx97QpKfGLdKIGZaP6+9hT6N
vsnzrm1zKoDJB1pgz8WJGfSr2vaqT6yrhYcR6yN3hSBdEFEybM8P8RC7sdapJ1qn
KlK1PJxofdUH3uCj5N5IY1HOTH78W2PALoYNpAeq/Bj6sGXIQCgmU1w9f5weF8Nc
pCrl+A6EMXL6Y3iRVDknKbpCV4RSrmLBaukzuSr22og73FbeC4nMLwb2dx10PyGw
2MkjmgsBb4E/V2JnvA4HscyFRjKJzgGwnn92pNTGLZbyS/zIOFnC7wJ0Wbn46Elw
d22M/jdFimUTWiB+x0J8TY7AW3kIJB0ht1v97bab/VmUb456MKFkdWzhsv1BYQKo
wtjq1gnNdadcCSXvtq3PHNQsO5KFFv1pyCVEMH/rInB7B7vSjVjPjY2MvchrjRFO
h4Sippa8ds+zNC+Y5YQsa3SwPpP7oztlZVKe+Tzr/wQ4RCsZlzP8POCMp8O2FkHU
SVZqGnfxUM7lVn+OxtJZr/w2up/XBoVu2mHjHS4N+MY60ZMEN682sqBOeKW3L9H8
dpexUSyDjCHAYqLD+5IzQDntcTabCRdHvm8pyG0iVsMQ/vb7e6rcoDCNtxEIia92
SmnZrfpsjsdjr/Ke9xdiTp+4HALC9c2mOqBrQzozr1CWi0/HB3VQKD2VDw+cn9Rv
ubgnToOWm+1z87FRoCNIUeuaWFQMNboegHNLxsl2pzeyre7UMPUXyfd7rX6oZzNQ
kkoLPtLLBuBowXOstRXaoCtH9worNBPeYEWMvJPNVKSLQxdKPLaCmi5+QfgFTjyO
Fn6unZxh1L0+3MEVYbkr6WOyr+NcHUz45bkg8/sO7Akgy7bmTy7ULM1kK1J2USGj
2D2nWOYMewBSW0/9YDKQTQPMUM/PNQp7F2itBT0TMQzKA515aM2zAq9ZJJSa53r1
aTdHnak7PN2ZIrRi6MD06rAmfe3Ud2vEPFiLV9fhu913vFMmOhAalFTsF8uBkhKE
2UB+lvpLYSIrQchQD+y+tNEoKDrFm6kjKMoetGNoFc8MQG5TmSyp5C1CxJzpV/37
Ae/aLbQLQtMyRdqXBG0yu/iyVgLUbjYrG2Df7Ir+KGh/s8bVb+7tJlOrhyChLD18
51m0ydn1INtw+qK0pbI4XENq57XBsL0HhAviGNBUani7GkmcLEPjplZJm+GvD3ix
FXCs2TwKAsLyQk755TIn/UauPiQld3Z+w4ZimsNOEts3wb4gKomwUtyEKtcMJ+9D
BmGu3M6xLhR+OqRr01Ow29IDrzd2NSoCYOUYm3h4DGh5AkVOfvKwEXXGP24gQf0p
tiofP75YPf2KWRKCQkMEsGISyp+oqXqervNvTGsrnpaPaZGZ4O6Lt5a/qC6gnRuz
jzbzybut4k1l39toaA0fTef7x39hXAxUC/8pNcRyiv010NFWzFKfmiYKs2UurYGj
Uk91DC34I49gu+qnj2PngUxMi8EwCLDb6dzKU88GhDPJmqDDk4fUY/1bDP37MVcF
CdRgD+YsOKYxIsz3gjHPAPRwAxV+Lkx66x2yiSfHWNIZ6sMv4cGRuIGHX1bPrnoZ
Isvge290CS4c7402QI6CZjUaw/cZDQz9ptv//VlasT22w/u9uJF2Roe7UuTW5Ta0
AjMuFMMDotyyL+i4+7ewiiDzpagr1ERkCWVT+1MdRtZzz7vNaIe7tkoDFVeeEE/H
w4DIsCS8XOzOIcEprrnPBn1/iKhtOxvsJSbIamk2QBg0CP06xMxaQyGJCXplaanK
YZ0Y/FA/CJb+oW4xzW/AztHSKJAzAfimNstX0XsFiYvdyk2VuzlVUedQuEdeqr5Z
7j8kwJF+0sYwJ6LFS7kKt2FAd7V4lIIBDP5Ye4Eu4pWBMNByujDs2cwN6IMQErpF
n0oj6Hp2adp/9m4oNA3oTsosIPdDHpPUCnf70ZI9F/snMqGeGqK8Dmmpko9SZaLr
VdX8wXqzgxPU+4HR86hNAXlKWMkzTL8IjJzIB1+cHIgs5NfHia04z/VcfNlXHemJ
bKcE9x1fsoDE3dWa+raz2CLAj/RVAevUyGadSyxRVjsiIJdUi+3M6T5H69jaGc3B
FYnyQXzsNVdW2hLuf+cwICDLyrxVRjmWVC94bifCYhfMC4guUlPMYTc3RAf7PHZS
zCpn0vjzoZSNQVpEifoXC0gC0OgNs4mlDbK3U6yE3gy5p7eP/JdkNI7wplip3+iD
7NHhOXB614ApNNnhRygoPtSDUdsy8wjJHeWVyFdrHLafnjRo3bLajwV4DP8qFBpA
X4rMa2rwz7G2bxKd+YTC6BxM5OCCbt1f/iNn3KylE+MysLbU66z/BJx7c0FAIPNb
+ik0NaTGrfAxN9yg9NoaDbrrDsOrOs6KTdif/N0Wc82k4768xfcxz4ESMsVxMLig
JqWRIVZ1vUZfgdoh/qBJ41+8QpVUEs2JK/enc6GJqUd+7XyQwhFPueIWey0fbvIe
rK/qzaVObkMRD9nzlPK9xKPPCO0Kx4PslaJ4Qb+Ba6hscj1eKa2kD7uNTXF7EmoE
x7krVpbvjcqIUDazQ3gYr8V06Zy8g2ZGN8zBJ8PjhyQKHOT3qyW6ssPVvO+BHYCm
lE3bYYcDeUsMDwjjXhKgvl8AXyt4GSmaUKrWkbYMnyJgg2Jdh5VSeG5tx2BBCAuZ
F7Ny9Mbnw1edf2PX0SSoLuwlgF/EHAJqFP7DmV1FSVAqB7mQgATwUPuv4qq21d5b
39uWotMM0H9DuKWFUlc9cS2pqkO9rMTyXrHSzZyxOK4dxAIpVXKe+r7LmAnUvajj
0PZm3uvkrpBWJQc1PDLlZGtE1yfFShTprZIfVQYNtkQbnraT/DLD81ljta8BzwFy
V5dPVagdQjNBB8D9FSoeBKW1bAivYXYhVcbthT9DZqWbUjSQ7APWOq1PxkzeupAd
zDuuNZfTKEm0K0Q7KFMRnSZkrbbJgLCqB0alU4c8uv+ghXMwPpHJToUSvxhPZ9R3
fg86oJBdJ/L1k+kMnFAY/kpPmWu7qHMoIiVDQSaFYV3709Y7R06FU/CzVg5eJDmX
+kqeUXLF4Q7gTYFIIs+Oi3/hHKl81VuMsH+9EFdiCQ9pQlMf4fI+TXLozE/RyPk8
ALhkvlC3xrX1jvs3NQbf82oh4iU5xJ+N2CgVBtf4+Ie5f42jpYcEv1RdxBD7YRy4
oTSSIOXGHszS5lZuXU/wVO3Z6sOQex4HqqY392eotJ1O0GdAP9y7UkMSWyUBUvHl
yG+gx6DyoHmU3f++GoU2BxuEyJSFYuXg2LFBOD6Q0itWUpXNingItsQxfpzQXG58
KBIpc8tbIQSoOR+20sbSsLusbtvN88Rdb10jQULA9eJ0qg22DwYocR6tAlmONOqm
6otJaIzKWAvAZfv8RxcwgojRDdPtedh2npcnPaJSYUo+qnh+C+UA5SN0IvVrCM7+
8qdF30YaFjeEehOpA69G9KV6cLwz14u/WBHnZj8um4pq9w/Bsr3veMKJZM8QuVZY
8GgK+twM3LrmCk4m9smRthz/5hZiC2JeBabM5O0DY4eMIiDzCC6aQ78JzYUPBMkO
Bg72tii726+ap3IzGIiFZ8BXC4Q4txH4JVlZHMm1GNKlcMxp2nEU6ZQKHyKbGe6E
Tg3hiLCZ41k/Ddpg9DYDPBhnm65xf4F3iDuavmoAQhxm4LPOs5mHIqsltXaWnwmu
+pWGhUOhdGrVc4n+bCnfoorDyZrb6aQ1kHeCcvdB7xds6TqUwbC0RAgvgphzbNx4
fY8Wn08z9Zrg2WNuw1e4RaemnM+sI4R0KwFHY9qqVZile1rf0TjtqZu2jJV6srJD
nWw7gYgVCs+hHl2sT7xAY3tx8cYJTvQbXLPcq300FgRsJzypACRyearDj1T1XsIG
CFlvqxv2wpOTEN5tGt//WRZvzJk2Bk6yJl4HQt5LdMZ8bp768IS9acS07Y3eiILY
o332UQEdDIqIVrUUCZH04fwtcD9IjhGJcGypyazlU+fBLHJWv8r1CaqF+8xQjMxD
mxh9ay7QEHo1LJYERhfNDZj2qLM7zKiuuV2t6qsO3mZlCUzerZLIRpxBlldCLAeO
tvNzYL/ELt9YVxeZJq2JCVE8+vfslxQ5raRdL6EVTnuJ33tKrNjieyslnJKsFW/y
OPHPeRrv/odYW+8CIbTNbEdZ6V/d05WkzULanrllVwLf6ZWCDcJcGIoCRMFeBDuZ
Yam9ChjUbBU5BfpHgUNPoUvget99CVEq0zJK4uVvaVnRFaU+GhVILCBgATUfyTDM
LPZ2mLRaGUxaPRw0D7cIThT2ULs+PwILY0uA3cXiDYKYrVY6TB2Ue/rr3of/Qm5W
PNlACUMxlAPC4ii8Rk0m/aLHDi8KoXtLNksfy4jkiTKexQIGPAAtg/ZCZaYMtBQR
vF7BB08Uxaja+0xYXmoUCrRgzwvMRZx9VX45LXn+clu8DXwdEU/+bYMKqXrwtE3a
Qlasm0Slh5tYM2iABIOUtqWDkebP2WYN8a7Z1FCIR877ednObmjzwJWwexXO7IR6
OwhuVk6h0tThJKfxm+45ARAdmU6HG1OXMpqqc8Grwv3WpKLHCzeKLRKK87teg/hC
WPtUw0KTx8Yho2PGrhjql7hxV8pf0Bvu/U+Axmgfj/VAWorVPkiWYfBl2aBDkyLN
hov0Q8LgAg5lVuIJ3mVMtUzN3gxdrx+d2WoLSYmyiI4n3GUoQMX5/De2rBVCDP5a
FnRSfu/vOFS4dBFYol6ZqYacVKaCxYE5eu+f3dAPsQ0bCEVymU6ZYugOUWDHXib1
4R7MZNlstpOCwK2QPN7KhntZAxKfngqGJfmL+RT64JbZEFMesrtcoGSr1aahwHeW
aOSSOSI1F3zEbHdW1OZegiaslbKxymre42VC2XBLNkU+uisJQrkiNl1x0YaS7rJd
oTyJFvGnJKxB+iTJOFvZbysJ1CXD8KRKDDyOK5sPP0oqkr73GDcs9ldJ2LsrsSUh
Ar+S6yeIDjOay4GuChrtcOqdTgZbAP6LqBP7YKJpmeZU1BFilaFW4h9oKSKOOeGu
nHYjUSM1NOKCs7+QWy8jobvh83I263qTEcaAfIEbrqEwJKAP2KkQhN4NqJgKzQxo
Wc38sBmtprBKOyup5kJANA1Qha+3DiU1qmh+TyNOQkGIHbyxQF3mjvRDCk5wOeX0
7aYi7lKyw8qzTDa76o9/0JmvwKyioLoOLfQOqATzmrkECGvYeXxycPJoQscCmIgj
QBXCQ/3X67dYhlbg2HqKYHBuVf+G09y/NH0lXmgr35nQU0GdHqJ68zxCVFqOTEAa
TaGPXRApQZQv7JRwDeQ2KLH9ZrBK7Ax0dgrAfffVmqx7kmepaHH5GGwM8BPkgp80
RRj1epIA8Awg20GzmYAWgPYlCtpfLC8+mNfSCjE60dsGKJREHkX5dbne+by6BgAD
eyonlsLS+pkixoIiPS7b9Vv4vm/Pu5qt5rD1ZBysbSfsMx8T6ahmNIHTr6sSf4hg
yb+ew9/prjpGe0uulcJv5hZP5ex9bV4hV4AvVAHVezopZZmJvSK6NlY1uRkuJU4f
4/qz2eOMHRmg8dDiMUlyB8X+VrrioywP1zMyU6GrcTbGWHkRtFS14LDnsRDfmH3C
Its6CqBA6M3UaWWSR5bB6c+7goRJIsDoFQgo9pxD/1E2iUAy9FNj2/ljShmCgUfF
Ramnkr3GkomoNI9UmmJ5+99hW8hm35hSNygB1WcYagocXBnwKbkjrzKNblIFFjgs
XeTYKc7BjayY/meypNC98V1YsDRaX0IAmShEJnLnANIow4bvmFtH6RIAOck33Aza
y5KwWVLBQckeTvikIPwNp65QUm4VD6SEr1VH5q8R3LhNWnN90hUyu/4CkVjbWykd
O7ZLJH+YFX4xxslH+++OFBET/IjWZudY0WWWjl4econvwpPhPH/2HcXVA6LNZiC4
vI9m+lD4QyhBSgVrI4X40EREo3v2GAopSimcGezoV8zjNR/HesrHqXKEsaFOMzXf
8w19Hr6sEfF3p4usL+Dgmznsky+MfN3VO6eFI1ebdQ9AXqacV5pIHueJhScEL0DB
t5pHl6JPWV9HAnssnmkAPIk4dnD6UbfE2fSQegxQ58bSnk1AZYXnoeQmZQ3N8c9L
A904bej1N1MhV9EvU8JYR/D1GAcvwCSOBP8vgaVxCWpVuib+5smRV0XZi5cXUCPC
MQXoSlu3gFW7HH1cKhCvxLKOlTKuLmod+kJutGMAHxu9iK1DR9hHMse2I414v4f2
HXCFTQ47n+5vWz+2HFiZ+Ru3hYZo6e1RADKjU0S+QhGklDlPrBsNA6Qi1e7Y5+Jl
W21ChqD8/bejlAW0GiCa+WFrbRJC0pUvSoHaVW22TIzmwWarFBt2H8AKGtqAMoE3
cwCi3SfkQXP/+Q3zOr4ylNhpqjZ2GgvkXXIF0X8vTDw76jftR7sTancAaln8OwHc
TzUiBWpi2T466pMSE4JoRjsmccQRlBwOxoa90to5cCVPNwm4ZK5nqcnke6rWA7R/
ikoz/1yQ+zb64MfzSRqGHCfcC+FtHpJiTgZifgIIJyeQqPXH3muEEi3g90w27h4i
ebUscyDUZ75riysRKrgsxqFiH1v5aZKG0X046m6pg2UdYzT2NIjx4JXRvxVuaOec
OWvV3VQmilq4pjGjfdn7YGEIoPa6vjMn6YmhE9emNuOkX7znMnoDWdZSr1Fxgojr
Eu7vUF7GRvVwMBT8ZjtpXw56KEGlUWR9YbLctDdPG0CTEZwqPrcWSI9f2/iIleNJ
MDRA9934rYmrviJS6ONMeILDQC2DQDSM2m4C3aGygf47qrqWiIxlmdPIbp6KY2e8
DcAauKo6BeOU3GhXWQfIDIAXYxfP3HJCQ9IRZrUFJS1UfVPU9LITNntZTAb+YFBy
F7mZVrKkqa0cG/jfOWtkKmPiEvLB8zvAt5VVu461jrhMQrk5EWVO43axd1FKF5vT
JK4Up7lPJ6M9CBJoer2MQwliFGKz9uEJezMM5inQADWq7dCU7hfbGiUcKS9ca24v
bzng5h+vJT4mc+Ii0Nwg9oTQKZbPrSv0y5MxpvGYdlQD5uCsfTsVjTxHioKnzxTR
mbbXO4Pc6GmE4UaF3xQz6jDH4mZljSmBDdmtwXyDczdcT32DpRrPFLQf4C8bwS22
gZvABIhkubdGjKdmcDIbpG7z7Tx+UJ9zZitBiRqHI0tZqbbHvorgMpporUM4vYi/
QlWEovNUcojxade32kuVCR9zb9oCOI7R0YLr+Yx75MtI/xg5HaOk9D3zyatvxjyA
IHEW96Vd9Gca6swTcaKB9oILJ8PWX5OR0yFhvoNqTpwVOKPaYAp/yd3UQ3AF29uS
5NJYb3CneKn4E58h1WlVPq/cTqMA/D1xsFqikOA3mAsWi8vY1ETcrzgPfBLtqyt/
lqajZEa5f/s/11z8Vm0e9RrUGPNiqG3wqnWUS5slhoK/AZ+OKRHDrA3C2/mMcm27
57fvuC4r+cybimtkcDPWWe87qgOVrnKHgyZS/H+756oK78G68/s9pp/zK7fz7fzX
F6amjCSG13V3UVlE4d888dqvGC5EBbf8tGg5F74YPddBliCF0p+riPtSr5Rdyeat
SDQpiqJzQrG4XXhDMVnxtrIarIqX3IYT1RlbbVn/Seghqu+PU937J6uw3E/VAzLF
2l+NONnQRR0nXmqGe8x9slr/vnehL6Llc9IDoDEx23b/Tab3x/DFIZ3zS75+Vd9I
q54PXe+TOWpBafrcntmrj6Qn+h9eK2vyvntPvE3X67ugqbC2W9grSbNJqE7I9OYb
aNuRR1L21LVugRknCDq59EOmilnANV2EB973AsD33xKWIt0taKs0cV5eH8EHkrY+
E7BcYV5sM3tETNYLsdpz5msfdpn45cHLux1oZGSSBJdv2eC9d1hofrH4Y515j+6u
rR1D9wTkTb3C7UuZv2xOOawoU9lUUg3Wu70c8yEJBWkuzUPTGwVLq1qBx2i5gFVb
IE6HTU7ZnfT/9LoS62bpjGMU9SvIlwgjPznRvbaxUPgVBtKJ0SrYFsmXCa5yUOCP
IrXLx8xxrWdt92wTP6JKz8vvqTlcs9EbsxEs6/NEPnsZ1JjNg9AlvWlaNPRosW+p
Ydgb7ndMA1mKaEFS6bsD57h2PnExrh7vBduZ2UgJswM5YmG/SamJm+WUMGZGhHE8
v0FWn1Q/pLGjOUaGfkdd5XKNiz38Z5UCQpOFOuz5CnSMIshz8iYctWyGmf96jYTh
s15aeOpI/nQ5t9Q8p6QMS15x38WdUM6YoJ6/AJlDMtaX1YaGJHntaTQ+E6Jf2vXo
JsP6vPDe9yiW98FF2jdvBSoopp7oQkloX8CE6iJKEctRyzU7CAGnQ4f3x3tMKaG3
MQZInxsruC72zrtAzG5/UMX+3k/S5dDbzQeq15kwhW4o2pykEmJJd4D5DSb1qgPE
oPYggKbVCGZQEjbYr/Dr4b60NfGFZ3PToqGvr0fwKbiPbBTIG6jYTMR/TLmR7Dpz
5x5R8HrntM2KsFkvDg32GBB+eRvu4otM8YJza0wph1jZtsqtUfJwyV/CXEcRXi45
z/Xa5me9sE1/VTj1hqd+q58qgBlT3NK0F1a0S3KY235Xug/I+7QmiQYIU3IcphAA
AqNlurEsh9cAaUxnjPETxgejRo7XHo4pnT7u+zwwKkvLnenqjj3KmAbGTu5TPdmu
IfdhIRY0FjGdMVuftB5QcLqCD4Ufi5aOynLE8ORkjoE9X8LX7VA8iih8ncHY698U
8Ea3rJ75x1B0UhtrNZdQ9U8GfO5WZ9m7VDrVopM99cCCfjYYeYMnBU2zcbjKimcO
Uda9x2YcAIEP+rPnWdj7SAKmB9omr9u9n2n/tqLUABFRlgx/+FV6keYCLkYGhxrq
jnEiyJu4uADrfknkmhD+MoCX8bKd8pt9RPvWUuyLEPxwozV2Yk/tXXFNEgUQnKy0
L9VWzmJoIbrzi57QfJNzP+/N+727oIodys1VTfNNFTXesk7D+pLW4CTJxnUclboR
3ZaAZ3vOviWTdOiNuZB47Xhqce08yjXkbZzi94eWhYREL0uXuxNOUJPRxQYzESlD
ApIcujwY1hHYxTJLVztnJnAcFSxd13pNnPfsu8rZvAaiZeZDScc4pnoSAoCDFp1E
X9NV5nKPKXK6nPUKbXD+6wvUh/m+YNmMn9L7tgm+R1cZII3LcBN9n8LuVK1k/8Fc
Lx99CDEi87kZmyGfe2ceWfH9ZkaN+B2aDop5vmqUv7kPK9d2yeULKn+9NuuU+VaN
/jKhGhkjpFZJRxmP5CvlpgBAB7gBoZKIRrad3Z4PYm0JlinSA/kF0xFVH0F2pvPj
dDTUBA03uDnV6Gvpp7vrNZgbRndp6Wj+LRz+S+hQGMhAxX1eCQuM0mMjshiQiJRs
hHtSPqB0GTrNip8VFNokI+1DjkLxw+8/sIUwXm8tL8+T3EyLSSSa3OnQs4iIYiQO
tAwcPjbWGOQBMJnPTG4hCDgsyPhywj0eG+o1LkcG9t45Vt/5vtMY57QnA3A9f9Hm
dV2FKq3xRt/8UQJ5eik/RdM4JljZ+tkiSJaBvrRBQZCbS1GJbF4D07k+d2RTzlhq
ux1NUic8ozkK4vJk+vyJz474nempS8k7HnrozPPk+qLTOCr560zVeVOywoXGBckS
5sLeDkyLmwA2YdE8eIup+2wPBL8nuVfdaYqsfovcLLEbI56v3dnsGoDoN3XD+B39
ziy4t4Xx/HK4RPJY7MCCHRR1jHxzLXl8UNAW+LV5KLCZU9VjsdkLCyZgf4gedhVr
BP0GLtjzNxXthwkkyy6QRfd9Gc/CWKBZPLKPBRH1OPq8WKQe+JXqXchXCxE4L4DE
wRQWQIHYdGurScM8MaMf3tQr2bpyKmqGcIHeuWE7u8m7I4RmrsCSBtLHbmX8Pl5C
lpKY/cHBcM2qwdB7OJGwEr0rWhKkAADpdBN8WvXl+GRAeZU5n33twh0BEPord4HN
kNuSpRyIKodKr+AE0gW2TZf8d+rh1HgB8L2lL/5Bo9nfhsHII/uRToc0HTCsPQkJ
wjFrS90F0SGLFWheqB3FbDfwokNZga3W2oZMiYrKVgfXG+2HOCZWq3zblbSOctJ2
XLiIAOlyFGTsZ4jar76Z+Djli+s9B/A+FxAQF6AtEbzp3IOaFZumqs729oCVYEXZ
D2IGl2dkfoWvsrbHIdWErwudfYkQ3oNfuT1fGLyUG69TqBcba8u6sAwVNYEoEUUl
nnEtyhhTJ75UhjF5P4xQPbbjOdWXLgQvjYyvxqEKuEw80kWsZRyu5fRLye1RWSPt
kP+Lrxv9p1u3qij/HylKe/2rIEbY24uH7U02ymesjEXVO5Rh2G1B7Gbq3+qfs89L
k/X4IBod0GQkuPbrOBTjqt/wAwmpcdzb4jWyFGXklff40OD5c4l60NumQdNWSfgw
P2QH/CHMMkVWo6BAYd7KtI0QhgrYlPMNFSQnZcnDvQEi0HgzlOC4v+FZhLkAV1wr
4yUYnmfuNbrq8H/D0+dmNFHMoN9QuWP8tQAlMk6cm2ajBgNATwNHUhDGsVekJPN/
TeRIy/z7Oru+RinNZlGH/e8MmAaZJ/F35QhxiTh+alh6rnSKHEEihI7CBXPxRSfL
nhOvkuvkV0QcqnmlH2ahk7zMrLv7RMikROUy2m+vZ3+ptBrPfD6FUmC1ZpxqRA6r
LfvBroxFNwItG1TURHksZN9O4+mZQ3UMgW3cU9N6julov3w0Dqe//4hQBxWGl+7z
Yr2WUVSIXqPbh5JePnfM8L0wMPaGMZ5v3fx1oZzBnHrxj8OeOVncihkoYB0IlrPC
4rydnehIju0boIDOhxqqegAQReQ3kWkEPeHbO1WFsmMXzjOm55brTvopHtJukO2D
Kf5b1toU4fwYonHUS6HREsY4dtxWwluW6HHRtUErNVjTCCUIIzQ3b+WlQGd69Of8
1IXlupo7uXgwpL6FkXI+zydfYbmZXJHctcm2qSSMI+AebOj21iRHWLe77lIe2YHB
d7uhF32oVw4x7KMSLdVl+EQYif4x4JrG0wjQlB/wreQ4sFPAmQHaVq4CNOsODfVg
i0bkS/PfZCvkGowrGtyPPazQ3bFUj+SzOXM0hgfSK1A/Ax8WD5HkUBe0NxKK+piu
fxDk020cDQrobPxbt8O3RfrqnyEweBMZNJUoqUsxEpqkbnphol+SyTPpl6yEOOZL
BNvt1zagNzgCRy5yuNLoCgBWfcCBgS/03zAjSZZq+MGgrLSHy9nu2z7ckAH5iwub
Bmh23W96ydqWrnQwloWC9mCbcY6PcDS5xGnuqFR5jZ5QAKdh7rv6mFoiY8IcaljZ
UAbcnazgJKKva74gDUj0rvauW42ZL36hzj9owJ4nkzeINvXzClPglbXVNqa/drZh
N1GqzxrLfkP8+I7uDELXamTGbVekgVwJY7cApeoORK8UWnVnl8j0jVIfriDpaZ3e
HL5DHVkYGvyiD2CN3tG0GumKdueMFjzTiEcRT0C4PrZvt683G11K9gHtE5mfGTm3
3Gl+JA1gHYiIWDX+4MFym0jJVOYliDEtMqg2vkBXjSdO+lj1aLP9jBoRJkIHCwr7
dGohrDeM4hbKIsO2A+Zwp8PoH/b3L2KsPDVq04pQXcd2sc9SeMJtDBuwmLxqoz6R
GQJcQb387zFfu8PW12GZZSyaON5yVjw+7mdpvNkhziopeySMXysZ47nap5i7dnua
CrPoRawOC6bHrmFJm3+idRLr1CkkY4cURORqbyi0XPtOJ6lKUI1TT8WXRxOSr02Y
CMp7Vvu6h+o4EFT+lngemrbylSQhGIoYk9AL4u/AvHv7iN3MHclp4F/u6kjHXyGD
7qXxQOBO1c9gryPTh0Spxe002TCezKS/P+VQD8oHkZfXzI0jw4ETdQUr97coqi33
lG4QovvhN+zu+R7uqVbn3ltGbrxFhq7J0zsvA67Mia0tJdW1nz/+CW2DtBVZIX+m
aOmjy9AEYGEQUsouoVD+QA0k1MMaj8G7YqEok25hVT7eLY0w3no/uj26AZ6sc0R3
wwxmZEE6pjb3PZVw1P76SfbDJivCbVgpQEiU0Sz64zLSX5x9fbh7qMZ0w05CH0P5
W7uMBB5Z4UsGEE0ScVhso9wCpcpthaTRtOZqN7ZaZFYGXUegfhlWrB2X0lgiNry7
mbjGkG6CcdqOCjQkKIjGO2NIQfFvGc2SDgG3w4QhoSwHBdZT+KGeX3NXMHM3WFB/
K2d/jofLyXbDyepUxpB56ojfTWg5hFscf0Jhkx65zePm9WLe5Gn/55tsl3QsPTnJ
sDLoGrz1eey/wpXMG+lnF3Vt41sm+uTy/44w+Sr9AMo++nvJkuVSHcS/exZHDsnS
bm9e3E99bqBR5FWczQYXMOWjLiG3Wf7tJE6Kuym5mCdnmHjk1/TVuUPe0GfqN2wg
PSvkqwgzKo3lmSuETdFJn9lHScVUx0F+Jn9H28FtyPDsbYlhkRtwuPNmzwA0HDq2
/aGr/mOayLzcUuBaEU9gBXs5Osx7EXS0vhxZaUozV60m7CDi16vd3hMkYeGP9uRx
gMxjULGFm8yP6lTfIeEpiXRb2evwnP9OqwGYhdJOpyar49MHJaiv+JC8lLAe9BRz
cPZT3LhPX0ShaXQzkLyuZACKYhejb/smZPhk9mMkGv31+rVAl+BMycWDEtueFqLH
bOf0sJEcxDFk6TeBLItkujHaDCCfE8QvrQmmEC6hcx3hgkRk4Io+vVXQwDc6T3Xv
HcTbQbwm+4kNEzCGGizKW2RfasKf7bZRUEOnpTbGYbvNXb6cqJ1heEgIkisua8T0
Dr5QBGF1EMgUv3IkZKfiLsdGjYChl5/1H3ifLkYYllpKBimh9qAx4h28/cKOFwnB
P/Bobg+wZ9fa+LkZG/u5HqajKBJrXQOIKDS9wvLaHkU6I6HGv6Iy/DoIWMvtulQF
HkUpcUiWdbDFLyy14w0ZmpAgLxeuQultKCna8rXLsXJm40iT6CThmXi7zR2vTLqG
TeRIesXAoo1QlUz+dveIw456b7sJ8mMscQ6QBIlirmvP08ChfjCpUaPurJwM/F5R
av/LmcKvP255uZV1vWw11FyigvxsWRk78HlzArVdLXw0ujz0pPzgh5GuvA5VBySO
tYVtKKxwj8KtGrjmarqjNywXJvkgVok+WuIzxsDIb1COoa6SQgrw/1BLznwAYRqb
tQRoJ18noNGjRxFAws4k7qpTrqHOqSWv/XEdSZwPU4gT2qk6PzgGLhUtCH2v7BTy
58ma9D5PmkiU2pmAOPN8io5raCctN+JxwJ33zQ4VtQX6IZ6zmOhzMlSjFc3iX+jR
MPdRczFkGCe8mFQoVkzRLFzeNsYtSBVVPmNPWbSSUDI9A2PNEofHJRhZGWxFKq2q
JH7RvQAek4EnU1Vmr/AXwVQAR/VBsFFJEHpNpdhXGoBoN8ZZ99SajeUnbFU8UWU4
pNIPuj3mVFkJ28mUEhq0X2wPEFpFMYuduiazkFbrJV2nh4GtakCkhfFTbtVhet/X
UGzNG3pO3RtL/mPYF8VNqAu0GfpJ3aasEYUs8aivzevUiV8G4GieRpCnJqYyvc8y
iPsVAlGjdKSlJW8ZuisENo96yyitoaLT0WyQfcVLYs8nlO8+Dv/jLv+bjdN6zs3P
DBon/f7jLnPCtDtACWx9EtZMUj2HVOyUNP4Z4J0FDYTLPxcpzCAE2Ljci1TrUjzr
Hj2/Ok7gUpNr1gY2MZNPSZHTMHcPRuqZm3qYUAdT6Kf6WFquZ8W/sXHbOqqkSLdb
XvvgHtEzVthj2wF1iICnPhg96ZiHO1cpmZYzZ4EoEMWtvSBBOD+XTD5vpmTWCTSg
1/HgyBlu7JxJ9Pd7Mp2Ahbyip/G954JGxuoobc0tbLdfNsS/w0sBJ8GIHOkajWNJ
WCJGBCV+ULTaHkjQWYByYP5j3AL8XZAEc3gLMf//R1CHctjPJQxWZwpKXOUj5wOB
sjvIlPyurqyRj28QU04vvd80I9a6BV8xMlrQKFUHuJH/bzgBp5C6dxMAsByN3h6J
PK22NxXUb1zyPNB1C93qayoVeil4zu48+aXkz03dXSkJRpi22SWboBahMaKxM4nb
02gkhq6n/CMjd22of/2gltAF6B0qZFl+97L9gj9Iu6m2IcHOvxWocnH8rjBDNn8R
2KKWrQUH4CWeqANX4khattHVaVx8AcxO9Tn3taYNgNkFEqT+77akBU4OqMOAKCWu
6tbufYSqXcg67sOiyuZ9bL3ivcjGTQ63M/gE2SNM40fA3W3l3gJXeDi87zQXqCCk
iNAzBmLUNERnyHaL8WPlt53zwUf4BS3pYDPyzxS2op8kR3B7Rm9NBMqC+StjMmKQ
wncWyy4Yn0L7bn0mQeFcA6QIj83gcBUml2Yy2yO+ErA3Zmb3UkWthVSdvjsLdSyY
GYT4AN5t19DhjnhW8NMIG9JQQk3Az6cyg0JWisMCVa6nnYinPTrtmV1csF1WsUGJ
27l5Y/66oZiSo9rKBg/HL8+pDZjx3TvOszcLE8p9TSmnKuJlNFq9WcIXhK6sxJbG
iuMDcm0jQ46Cjt1hz5hV4qMliLwrufRb5gpnvs4HMbDpu0kBy27+Aw7/BZVyADIg
wCop+7c19hW/t1wLtx6tpLj3bmjB+Ly3Y0xLPu+MPtBVD/yBj+s+nJJqgK/NpTKi
bKJ8fCcwP6eXflcVKTNPcpDtF15kGANom4uTKVl+K0rTWCr1PTfyA7qajQjneN/b
TZgeZbDY/Rt1ch/QmsrRqwFm9T5Y3oqBuRKYIedH4Wl7UJSmXyiamfYT0ptsuvuB
ZbtZIV2qIdWUgFVpNGHxYaPP1Ihvacip6GaosclipZ9ITohxQnUKCkoVy3pEP2qp
Jv3sdL3frn1erTOR5k2aY6YOSivZ8Ddb2O3bJq+73ZomkDhvTJ4xM8GelEDVW4sI
hm90KQUZ3QffBN2dxLm4dyReI99yKN/j1IGwk9o/mSaO5zRxR+23Bjn4Bih7CPyn
Fci79ehUlEDnWJy36aqf/i7NOG53Oi0+EgxPgy0aY8MvqF3l2k1GemIiN0kLC1c1
hdaazVMI9iKambCkaiqSoVkWVnigUVL0y8Y/LtW2lUSopiNz2yU4qy62PtasK9HI
EtSzGQ/gZasBgJckPT3fWtSibNO8+4jweuYfZjHEdh5U+twuvGETElO1bLjspD5B
2ulJPf451YRN8QL5aw8qFLszTj8splik9T0BRIayZaeHzA19UXwgnZAell7qlwCg
Fy3N4rcmOlX/5iFDEOQtArxabCP8t9L5jvM27bBif9eZzb7uv/gesRgll4qk+ScX
40GfWYx0Ggdn4H3au+SlX9zN1+FB9TYZu7W0ElaRQLoBR/ze5hczTJj0Ykoiq+8Z
/r7kHg+LBaQO1eflNYujhw4B4JriHYas1je/Nldqb+5xF9kLmyeVEEVBhIuFPDYN
rERfALSLGE8cGUYQPJ50tgHjcajLlBPBFDvtxyKxZdqG4yGLcLBunJgVlzWkPyRp
6nDaTmZ50AXMjh83NZBrMIzBwbBzOr9cRdppbhahJlSsqDUgOIs74oV+eT+aNtEd
7+A2RM71asYYtr8tiAslwOjmJnkwavs6T13G1Y/RQA+jcQ6v/rA95nXPRLJa0nT9
WU2mjCwxWCKcWC66+djb86qrT1NdeVgJ4zwUV8M+RaxLgtosAasqmPSKvFiCdwes
5xKnxhBLZ8aZEjJl6WlZCVd8z0Pw9wmidLQuodOPz5DWDgy97DjoFO37HJptDTtT
hRLFgxAcVxFRaC+kTaIXhySzWwyw17Q6jTu7UfqomC4uFKZtfO/39e7U4Hms/KZl
B3842HMvn3OiQ0keLFDYAVeMHNGu3qEgcJeMRHIygaEZRdZ82YCjesxwG+NtltEz
VAhnpHq5WDYijQDfnzdWMdyAWmk/1qR9xOARUzpcZP5jxJA8PzZF6iorxw9UoCWi
Ba37p/l4+XpEEdLLh0pLcizlLeiRKdroP7o8l1m6XgMmPiHldHVHxSFm9qI3JsQS
krbjIdckEZ//Alp0tTd7xBsu+Asob7c9fEPAYVscONBe9vO9G6alCuWIv3t4bv7T
oZwvu2abDkseR0MTwy56FEI7DGbcQCLe8Xrf52zJQZSTuLPDKB0Vq/hDGj1sVbbI
+5V/rEVAzUgdavuysM2fnPs4eVi9aMVI3+l2rDEj7eArw6z/qIOkosBmkEIb9n22
j0uHBXZi8ZK6SFrZBJyRwPLtrUPS9XzSkS8Qp9+cUaISNX8Kqtwpmf4Pu04a7+Ie
+mRi2n68qABzYxMfMCSxFeR4JCRj3MwcdB8wryhB7zNl2Oo41Lm4Xv7XxKZIAceh
2ys+0zF/4u4oi+NGXmd4PD/JkpPhUjRMlqiCWXPqRH16eW5lGrsepCg6jFa+Z1fZ
NEIztNMBEa2RnxoU38VjmrCv6xar2TlxozOxkaY/HkdGVGbZFei0nWuFbZUNBa8K
floP0opRg3DPG4cQLV9PU6wGUIGZpWCsJ/5BE8wWWs6Vw3PPHPohLlhe7ev3YrE3
Zd34CEcYepMUv/vEJQI0P2DLBH/wt8Q3NfHnaMgwG7cbMpZP90WSBTSkskxuLF/8
3wJuDOmorLt0dEpy4kgCI6pbheX7YTwxEcU9N76KF4iX6kAgjcgbHYjI/CgxHZjS
Ce/Q5Afhhm7SlGLpasFNE1oEAxjLXSmgfMswQPod6+wSZ/d/YW/Vo2b/kKJLREqf
Qc59+oa9p3O2BP7Bv2nAMCqDNkPFZ9xEBzsCOaFvYi/DP7eo4dj1I4Y/xnV6h8Aa
U8LlxUOVAKpxoZcT25ZuCgIiQ07ymsCOK4dpJ2k0HB2IuQ8jNn2/3v9dQbsjMjUc
dHzD1taZ63ixo8e5wrKtprcVPMPZDnpl0uAipO3Tp0Y+OE/1sagenWbYP91P3UXw
NHfLPL0hl7VqMpRRJkQivpqZnpzmoqPrUWhuMn0DLAfOve7PLoef5EiLUyMf5BP0
ZwuFogbT3TdpfCOlNGVUZ63NX/H4Ob7DkwaKjIHTzTQn1s1/4961kllYveVad8xv
n8oGo+Du1H1n19v3Jj9WDDJ8jQyGIXrFCDUUONkLpQhhKEIStDPZDEKO5N2gIq6W
zhpnxFhFDkol7PT/pJJPw3Q5LqDkXQJ7zLsry+8QQOFwwtIzsZa5NTXwwi5EoOCV
rqg1vdWO44XDbmwT41VEYejLwrwg7IRuCbGOm5eKMEGMY+mBVyicA3E5Eo4zaFQq
DYnEG3lYppNsgwjPT4ithFXMTVvPI5QJt36EFz+uYdrFGsmyl1WkE+N/7uQMkgbL
Up7oKNuHRXMqzF6DPUyQTNIiPsKuB+mR35qLKcVGZg+mxoFs6Ixkl/srUFYO5UuF
ccs1C4KzsSjUttTZxSlQ/GkeGd0RLG7AsCgxm3pNYyvMRihCNQcOd86yfgu+BS18
kjyl0t3eYmrZKmiKU1CIUmOsIvVNr+g4buDf/vv31RSSxhj2/2Zkz24L6PbPia6V
K3psGFMLKEyZ4FDqV9hHhVWEcTwbKy46aMpDrn5ecztqC0Kzv5dCV2wloGtroRlj
/BRF/lATrPQoZmhyQXMYI2NgavJLeDwgIH1Ez83wIIIhNwJgywD5v4S0DQJQ2jGg
p8u9GpPRV4ihSt5H8XWKt9saJ3E8tMG4sYUtuxXj1GgJKtPawJjNCBLrkufg3eJc
g0CBPwDQ3bH4qbRge3sGZkSMVPCF5y+KCuqKeqt3AiF4jRZ2b+FmgRsbKrLFhPeU
+tT9CQMF8Ommr9iSvQ2QzEpBb8L2bwI5OBqHpHZAql2OCUQ560S2mDg8tZq5piwh
/jIv7mOrBjs584KixPGrbwCzFWJlpaymZDMQaefZ3Ewz0hwzgLAQkD2JMsglHyhj
6BAzD/BoLYcLmzIAXR3xRQ0bXGXhCrWeC9ACuvT+c80yQjTcOJgIn+G1gwBLDXMA
snsOi6a6brhO3IpodOpU+IgymdjuP6gxW2gLLs5Dn49E7KN+t24jLFl4HKO9WODw
YLGgYS/ePrRARGVsr2eqi6rjSjIguJiIJgIg92Qevs7tsb3E794bdcZ9XdUeGOhD
4x1ohxFQY+MTMAl+WLkwL1jIcRTIcNdFkhgnRyhutBS9hJLIoxOMLV+is06VXLBV
03SK6UH4Ek/lApEGOZ6gr/VUbroYZUDf4qnD/J9lYQTvWPOQF8Lxbbsy2DAdL4BY
6ca/9NtDo4lm2fYA8QWCbkILVrOkt90yzcJW6NRPknI5evsHn9acnUEtrX+isyf3
UrmM1Mh/zRLWJhxWWIjz5qPjxzixbzqNjc3GgxsTwqcd0eHxZ/rVVqe3fPdaU0lF
Ejx4WHEsSaFcBWPIxj+ugkjU5DFK3CFjA1bBzKODOEe0/Q00JqXVZCkJhedG7uZj
LQxJyTddV6iTQMv+e2bLncFW5+BMoOjvA/1LiasfCQCwFkh277ONQHVbhp4tPQIV
0mKiqdxdGrEOH/ewO3M4gko7mmoAGdfR+Ze/rXFbGADP0NCv9v/yY20sj0LJ6D8Z
udfkdg3+nIl8Lc9VY/Fz5BC6r/6s+m7wRSoFDpK5CNsM6iqte/NGvP428t33WsYk
8DpO7k45CAS0njt6R/w+JNh/1NXuaT+nM29TGxDK46Dp/UlTlQ4btpZlseJ5z5UM
ceZoc5FvQwtV+7/PjYwYxYYB6JVHQTd+J3gO5r23Bz0KQjUq4sX105hzjqZq6HtU
07/WeGTvkUrcpDOXFa0W5XhL1TnhyGTmk3dlQ0IJNFzWpjq01OThsXWAd7Sv4EEB
48xqJ7F7DwFaCUHE2APGNBn7H81mXjmezDsukGAYVXfQjHneQufsp1OE7eKT8Kib
LtN48vclg4d4/oUnGOxxd3KHbRhEj1AXWnBk6I7Rd9sjPrASyOchszU3BZCix0I+
kUES5vxJE87mB6ClDB2H0rODFOkp5XMxv2/8GNuEY/R+kgHYM4TSlIv5DE9YFdqL
uZsbdtOV7sDU8M/pOhRBgVHf++6SnE8d+yYWOskl0quuFBJxIbTrLDR2iwdJCBId
lV1rHV4zkQLD55qDeqSEyBIyI32KMtKG5ZW3RDDHF95QRUM95FPBFrqaH3N5cef2
zoFBcPTntQkeDEAvo8yPbAZYyXZaGnIv4Q+MARwzJ4PmEWecZrSHpWBYXUmipJ32
MCJxaQJpv29US9GlFzKe6KpygOTzIXRPAR3tSCoKZ4BWuq2UFY/WqRqlW7YyzD/d
fATKF4Qb4Tzof0w1Qh4uxpEL6PRdJ4Az6zeTBYhFBSanZx/xqC5IAMnQjn6qcS9y
53Mrj5xLthuzbyHEWvpJqSDMFi6f26GjkElXbm7VUc/XsxcqUmwTVokgKq5rdyGp
cCeLUff2LP24AS9maRwNJrGoLEuvW08pWNjg+jmbcrfRXfSGKOSHp4H9pYNdyprE
FpqSoKDRVMzfUUQk0Q7iFWx751R9mwp/onFaw2KMgn1PNbvLPUx8I+lQXIW2KG1P
NvABQ3oLMNwGjvRfIOLC+Reae/kFkx4XObgdSaGOf5tQBKraz5WX96GS0ncJRLGj
DF/iflWPaxKlxncjXIChiW6R2QCaH/oZTFgyC/GKoUpNT4UaCqiU4VM2e7f5/O+Y
oWcBj1+HrSBpq64KbitzR0FIbfBTLCmclxWhmV3FjPClgVmHgJxBTbabz/6T7aPk
z9F28TNcyOYOn0ug3QNIanKG5pmj4swhwG/qHSGp/IpRFLqBPMjy/D7V8ub16G/a
A3GVM7ENHlK/NqPmtFM3uDE0pxtyt5wnic1iBdAyHHJsc6XJGvykLelaGwiD6YfX
UkTbusDytMlOR4FN53hfuHJ/Sizm9xU/Hh3he3PTkGRLi1YYKNUjOcr82eDEaJk4
6T5yqX5agMmzmPlg9s6xVTfUkEmZAl5yuU5ZU8zyQL7XLcxDug+FWi3+mRXfEMzS
FSB7GMx+nyQLfQE/s1MA3uD/lIbrUQAgQt6qgh+Zv+LKXjAMSnvLJ/IfbzjV/gmV
teDbAnfX+9LJXE1ISqlJgtjzTKhbd3Sb1otisC2F9ES7q4DAtZfP9oW+5bViyKR+
kOsVGM036ehyjMuaNe9bq4XmpkbpwsfwjbrvNaQsgYrE9UkodJeDdnPTR5YHElAI
P7wr7rTgHYwHume14gWYVlyOl9qQ1kVvZMU+Z98Gd0AiUq6HNozwTwJFGAGCiJjw
zBhA3suGpFR0tCfMlRyScPOdUvzDwLN5wz+c1oL9DEeBPl3IQaKS8imdk/h5DQDg
JyQbNBoT/zJJpXnh1WT74jb2LcaRwuZ5N/2UcSqH6ZNGhlETyio5b7VUvR8ibaoG
q3D4bXBrbs8yak9Q2vNIPx/Jc3UKLs2qNE/B/2nO8pVy6ZOHQzg2e5e/pQPUC5K8
FA8/mp1v1zcNiDGRzlXt7yVWCptI/juiZQEj6gqGj7rJSh/ym2eLz5aqr0Y7er/6
6/l4yIIEfO4x/e1bqlRVknp9VQvDTncIvH06QpMBZ/rkXJI/rvHbRfOml29wC9M0
18mVzzwOONxk7obLv85T9mURWGuQ8UlP4P52CoAgvXFvD0ac2gQDKakVyuwH0MIs
+60mlKwNVF0xjtIggliMp0gFw81dOhj9CWDqq67r9rRMikAFqvNls2Afm1aIrH6u
qwVp940HTAlBblX472IVEs8hQuHMUSpRVKc4GY+4d8zDaD7FhOETrfHfRXIhc9Bf
j3Fz0LHELOH0b/MTxC7AeONt+FP+OypZiLzcVSNE2UZMRihOp5yG4j52AgqKlPHB
mHtyVUS+/HttVHmDuoZ1GPfy4IV9coJlgC/H5iHZVzQTbF3jJK+dDvJFmrwE4miK
pOqwdGTmkc1/hvjCSOeTEAPingG2Gc5zGYLzdO9icl/m33RT5grA3TOEy+iM1hde
hIXC6tDyUowtRBAuOgl8QxjwNDr5fODJV+2yXeKUZm98B8IxJIN2CYF6PakGOqWo
m0rwBWgqhDY/lVRzs6w1LhHP7tl1WZeLIqgNdiug9HsCjug0uueRWSn+s68HOu+w
Wzq3nXNZod2I33uIw3Di6y/4v53MoCKx9XnQDuf2aEKU9ocI4hz07I+hXq900NM9
GKPoFjc23+CaKW3ikWOEWZ8kas7TerJiUjF0bKUVgQ88kd44Pd3tO3Fna85m5z3b
xeRHbzjNq7LRGlr1cCXuqNnQFnzJwmVW5mht1y7vKEVEMoqi0Y9OIhbqj4he4jcA
i76kyYx8Ir6r04SSyowJ/I6mJIh7ZraW0Fkc4une/xwlwUzccsxJz28neVKvsoDy
pyKzqR6Nk1EpbtonR/rJiu0g5XWzCbNG67tVb4kOotlUHUD+V9SgKlrC1Whlu+4i
ZHk9MrFCGBm2+3X975SEQy7B13VS2nWV197uQ/zb9cdw12K8X6+EdrOthEK6Iorp
qbvoq6q+FG+ot8BKji4pCTO/6lxJFMnk4Ii81qisSILyBaxeFJziptmMpAdGCmXL
DcqZwLnRd7wDCV/BgaTnmhYbYkiFd8zDiqqrLBWhtdofthF9mzlmXn4nK5UzuZPU
BT/U2eEEmGd68ukDrxD1+cwHtlGUlsz4mdhe33JeZAvr/pr16/d3vf//WjhA5FJ6
gv3BA7/I6SHfhSOERHyBwwEiOmh9ROKC4SyD3qoYQshZ67Oh1SVVaHYpgqMOULZF
Y5AtJPUyxuoEcjei5rW1HbrVyRT4sXVhKvZQz/2Jlr6v3sd9miD7bsSYAr6fxuSI
FG0xVfs0ogcRzbMSNxU48mD7KYhR27HPMHL6lMfbg9iOygY1aaoDD4g9SDkdeaBc
7MuIF0YoG5gtbtlXjNJocRmZ+7LVTJL7PI3Wk8mVjKtSTw/K9yLDGv1E48cVD6eD
P4guE7DClPQ4g0YZRFxv/XD9SoSD3FjYCiIuA4uHQGDd84kB8P/eegDnJOQRbYfv
dbtMuccKWrOuxO4pwNhxUJb035TD6ek1/LIWu7F0DCWZfBotredHd2alIOGLqHnE
95APR2pOpsw0fy/dJDAp9xq5+QpTKf9b2U5TWdZswEb2CyOClnalPGYu2Vjy+f4L
cWBLE/z8sNi1SOXcOX2JRvohBt/j+XDGFxaRW80xPOhf8YyMXm2eQ14nE5MLRLsi
73VQSbtC70+Z1PNcJGpV3RroZJNTy7JWSbvdIyS4ugZyIPJkjJJsh1YGeFiNRECV
cNpC2Sw7+m4WRmsANjR/x0RBqqs5CaH6bkKrgx9Lx1xlmKIFTIUNs22nJkUoS3ya
Xe79Ev09GUcxTQ1stX9dKnqaMah43fDaNgoXGdUsyneCLgTFsMHhiW6MNgdeBo9G
+Qpa8zFHqC4/i/JZtle4LH1dGE7rhtttnt4CN1u4se1lfiISmJpwYNlA0qNvt2MU
szJCBULYohgUaDrZQRLV6MSO7U0MOcQ4xdvstn8iWaQMY8uHClBdV6wgTqj9NhDG
E+RTy/C8iMyL66Q42nPPbsnWluHYCo60rzDewczSYNrJ0q+J7h49Oc1NRh2CeReM
hJI9pPRcovBB+VVkW9Cssq/RIpoXhMLO1Axj2l1tkhrDdoqfm/iZ3DMuGC/T6lMM
9DZlesVLTzbbgHazI3tcsaA80arAPa1fQHJDPLjkLq5gGsLbIdPLwYfP4ix1YNg7
fOQZazhdiqihA0xzhfyzdcHpEXiWJ0SvXKme8MVmQVl08AVpG8r1+DZQUoQFh9Xy
Zw2voffvI7HjnUyC8KGK8WDm8XBHgz8s9GnxlgRZ6WBiEX7PPik5XRFyDjKz5982
i/u1er9mvBIMxZKw9JKBJrjQ1beFRy09iGEQZ6cVwL6z2mw2X2vMVDdC5cUkSyTM
BTF2JDM4T/aeYTbHfotC2hQniHfKKAk5ovlNgWoA8sSakV+aqkwHjnwyQ7PdeTjA
XScUbxVtyjhP7ouKE9mo/LN9SndNtRXsq+B9LEjcl2gC9luA9xIX/AwuIWo0G7bj
eLNRWUmghf/gZsbDHQofceslvmhBlcEK4hYYVH7mmDpyBkCeOz7pTqxAbXEkXHuk
M7o4Ur/uX3TyVhjxSevYfdykXABXNkLjyi90rd3yBdx+cIU2QSmgZfPqZbm0lcdg
pIwrinmkG5mAKopirHM6oploIoUrhb+EEq7daE2bxGfpI1sF9oQJ8i+QwvRIAoWY
SGft4sO748kcJjmJ317cnhsRdmv3rvMYbnwAa8NMukP97q0h2YWP84NHvFh3WDJL
dEJklH6CKmZirhNc7U1fYVDL/BXu2WCoV8Z8yHQO713w0NkfL9afhJkqr41OWhBP
aQe5ld1WIFcDuATHPFn/NHQMq6tXxruL93rfzyVYVId+1TetAbMmRdqVrbGekEaM
jbT4Ez0v5Q5KTl1i3RN06dHbKDyhdRnSrnaAjRA81zp7PjqpLZ2oOdlgjZeu1Ga5
eRqcJoDz7jAnpATWr6k4wPmVQ/8Od9CxB9gbbnJsFel4g6W2Yvi/NV3sZ6S8cxBs
INRfAROfRC6x9oatbZPyW33yTshyLY85ViOw1jVvVMIptxBRXZB9AVSVYaxoaFMV
5fNsqLVUETB063PJzwQwoSXZ5oxUxYfHFpgC6EBXYT61Yzd824lmc154MFU2c1KN
62i67UDMzdQEA58N/S9SQUddkBXgd9JsZIZ+njGhQNpyXCnGRwMcRpjTE+p7v/zc
avEC5/QQlqBYH1d/OODvE3JEDjHupBSXbRYzy5UdNOG2N3qxQJeykR68yiVPc9oe
DdqaX9myNrM3aDdJzBXwqVVzowOtK9ejJqbmoo/l4LMP82M6LyLUS9uXZ9qd7T+u
p/tfW6cI/ysSv4occFLSx9cIpqqi/OlLdV/tMRlIz4DMsZMFuImw+N7VQfGPxVYI
nSzVkSj3N3DTMUJq1QOyoRHqxUr+6gppY2dZFFwsKPVC1Yc8WRAjCTHr7B21MyRH
zBmwqa6QRzXoKdwRYYUM0PiU2oCJ2MhR+2h0gcRC1ael1eDSPjwewq6714AIJ+Lp
86g/oJgG8F3AxB3otbvG15JuJG8qvx/6M+cJBKhQvl9tK8GK4/AQ6B44KaU2qtDG
0U8tiHl8vhhM0A8oRb+XQdB8JyV6PKHcVVWhXGwPoCqpMHNjZ5WZV7hEXpmPh2Zp
0FFCKXBdVKbTJEuBTgBrTpOieV0HfSZqRuoxOM0TJhUC45yALFp502U9UrtAXMAf
Nlrp9vKyOOC+UVW6S2Ok5qaC69OOMuoprp3A5IyiVo/b+YCOvCqLK9AAraqK5Ww2
sel2KZ8JcUelIPf7g8ToJ0E4npZq+8QzXADXNIuEfgPy6zq6RtNeOc+yMXaOSJRr
dyurTV5KsTQ4QWKqakk62gPRaqmLWY6YhCnEC9OiBwqQd5hBRrOXY6XWrp0LhRyE
IWMHohvFN0RuyPBHLB09DbqZBNtlDdd1lSpJ5dN4EzQJ8lk96GwvbHhS5Rj3V+JK
o6JUC/VvSKjgdk+RPD5Jpl4Yy0rDoyVOYeAfQRP6F+GwDcW/yP7bU9sKIMb/1r65
FRYA117EEoGZD+aVry2Tr/ACHmt9SElMqhdVekC2dNLN6NJgtbuTzJc1Bno5Uw9G
o/fTPpwRT2iEgOrrnGZil1/WYgGRFlpjFAat1T3rrdyQj+CWrS8M2xe/UjS/QfnX
bPZ+vG6gWFRtspNDsxYdkBTqJPGodmEMc/oiPvJ+XD42061sfNxv8+4my5sf5EcH
KRybeGlVy3xiMJEJjISQwInneuD6Wo16Tl09Vc+N4dkQXlelEilCn3UE9xuz+6UN
TRcNhSyMPs985FPmm8xCL56zC/2JjSSQmXs2VbYXXMYPYKDoHU6/tJl1wBgvWFZ2
1+oO107tIyN4B2eTcRuMP6iaKBgwhcVAEbR6xstnykUe/RbhF4uSIO5zCVdCSh3P
dYYsECwP6cykHrWTQsIKZGgC4byBv3wORahOQblQmeXtl38x7DtdhDR8bTjXTytt
ZRCGhlVbNdmJTdXkmWw72R0x4LEzGpw0KwEFg8FgvxLSuHVOlqxYIXrOVSKPw8R/
GY6PkRNQtiL7ufBkZt3h986uAzfjCnn3xMYgV/gsaTEhC+C9UzzphP8v2pLLOefO
iTC6ccw8sMH9mrgLo+NUFRdqi32G0JY7uL3ly26DSbX6itTn9aQLOP/Qs38PE8/8
+ZDcXgsv2+XdmxsOsOJ4/e85hT83HOzO5pAi2nxH3lr6bTX1xIeIZYigoTWjXLqa
VepMDNVTL65vT9lRhwzu8sXrRtaPxtSeQ1EpUGjKoJiXTI9wU/eAVnR/GTgKxALo
o07vnI3Vs3JM29b8jXVXd7OK6gI2oOgqsHAjw33KiCAgEJHsmzelUo5NWSV9vHLj
8ml8CH+IMc8PDpCilncIjpQYq/Y6Mair8zWHFz7mB1FpIgiMU9RacOx8aZIr4oC6
yZ2e86aiMdcBTfDwh88z+Y7Wf1/vWLYlaihgSY2HwH8goYAM0V24dvJQX0v6LAqj
ord6aAK8HHJMhWDiw8e47mdStVUuVRy7ZNVAXhUMGZoC0EsmZ52ut1f6XnG7TGel
e+iCrHBMm9Yqa61SRWTITFRBCqrVOjbMLPJ3JzQE2Rv8mxq18CME/cYX65ojMM+E
5P2z65ZxWlm1knvtGsUBQPZywykycK6AP1PYDYWwLdKkF6gbjimr/cWwhqOTv/md
HYWT6oDL+3QKzLk0Xv2p/ZaxmEbWMbEbLXeKN7tZ93VZvovYf0T4eS/yeDWKE0J6
7C2o2hJxMRynNSK7uf2KDDE+71VSoTYWdiIbUwC5NuvAEBBcaN2//0UlE8WMy95P
2A3gmL6R7dTUnce5RRV4ORjQk08CtunNMudU+z3Vf8nGsDu1WWXLWMVpgyYHcLl+
y5d1aNUXnt2IdIL+5hLwi4jehSkeEjQs8qmBSUxjHg2H9mZaJvslC6mhMKLqO0rN
uKxVsq7tp1BLGG+3fa9DQESXiIPAXUA0QpsGWxvhLZyC4En6ljWQxd4c6gDuALlG
CGGw0YSUJI1DaeAG8CyJHZeHAi8JTtPnhu+3bgxyzwtq0E3WKeqy4Hg2S+jTE+li
kSZRPDZ1Fm8hnOTXSKr8+AeyV74CmF82mhhhEPjB/GwVCP04TkGdi2Rg0/nzPNU8
JxqZDadWUvSuVV8MdpeyDOEW0D7TzKQdb6bXd2xXE4TG2pOMaappxfG6r8beiqrf
za9kwxn2DuayHQk+JRldpuo/uwg9qvOO/BHIlP3PoMdeuwsV7hHpxdlCZzJQc75T
vHjU31YkjgFTMTi56zqu4hLlkGSiMnjtskMLLsp4RbQY1njF8IttLWGYIhTAXYcf
zCytS6D+VbV4j5I5j5TQuVKXyLdgQnhgqp5OsdaotyeNvq4bTZriOvVGwqkkh5V3
LY5VQVpmSByQ31sFWcyE78aW45IV/7zuu1gXPo/plMRJ6jTOM9FB2/sOKJ+6yk4q
ABsSb2ODKC926mrdibg2mFpuNU52T8jnColu3U36KP7mkf/rBpHYGhN5xfD9owLj
oTcVSnKcCbl1bTXrRL+hFNHaSflbUU+x/gN/EXzkuPA96cT3zgJ3g/XOrzizYDHZ
d/TnHuVFazelcN4Dgdf7xen3+t5c6JSRabkfPCpR8UJLZKuspqYBVaLrJoKDCVjE
id7ARkiANuLHRJfgwCs0p4b1vAGWEMCQF/u0A3WWaWa0yt/g61j5OX7BeYXw3ozC
wMiST1T9RN8dAa8EyXzebmyTQAbKxZNkwcgZZSSleAU8PrSheWB+xE5xll75cf3x
6Ux+x6rqYfyNNlgS7Gnd28emonse3HTEkQmHWXSNWQ4Fo3x+f8yga0M3iVK37jsR
x0grXTVXyMdXTbtoCoHdAt4FTxyfuCOm+KBgierHC5bNnMcQUfN5HPGycEMlOEMc
0rYgR4JoJqzeigNpGlEIwJbGJqEnzkt+aq/EgAO0jxN2bpM8AtDTlcnIsdERiL9q
laYoY4aaAWjDMbo/n0AmX5un/k1I5ROteE01fwzR+IvbCgKlh+0K3m0AwH2cM4GI
1jCeDdtZI9ohlnJoqTpGCrjvNPgc3/PdlZ6Dmui5HKJ7X3l8g13sCdF/IlC1UKSL
lLk7nJpfNNs4UcjhBTmPJpelwitCtpT4SvDMBYaZWUfSiaQirOxsonLo1ODFTn7R
TCqrwPT2BKtJ5ZgJZftqRr8twP7TmKWPL7/iRmxgKoJR27XYHx9iyvFO1p2da2qL
DNGuHq7CJ5NrO+a3z8Vx+LLr78aAf+vUMp5Y146DfNunSqSMKp/i5CtVGi0PRhGp
hzqSXQ7qcHerHwLJ8Rzi4lZ7Qbk3l8apglo2WVtNpOhO1V/qnrt5qIJJwJfDsVn1
QC42oXyGPkG0luqAfuGILYD55A2JxJvTLIfOfrlaagOLcx19suD85UbtWlY6aQEH
GLdnM3sSe+taC+UvrhQnKx164Oo+hwPAK6sVuW6pGPGb+WwjCY8NgqDNF8+M4oi8
R/czrCPrwsfLaQEwrQ43e/PwrksKCWsYLKpe00HNBiFRYe5uAZJJsdQz0fD/ZEPY
OaQCpuBuKOwp1TsBjwK5FN2KKvVYBr4YTl5Y3R2Np51Coa16M73WXMv/Aqfa65jZ
SvQPX2Kg1+E0uN4XLOyvJ9/pY2l35iUJP8YfCJN62MuYSzuVZGdL1oNfLFIh4shH
q/CSPckYJvrBUenoUmcAYYcpaAyKiMb+jR6NKKmZtOM/0IWHkwBuCnSZyL57BM+u
7X+ws/RQeQygHOMKTHIaSCxK0aHyGLNjKsD2axY/PcH0FGvMRpMJvKPrs7aeMQXc
SsZYA/vnmgp1tHzPZJ2yxqa00wFqCQEv44r+lenjnZxY21vZrfy7VrOhShkCAdhX
E/p2FDhm5y5Al8xABYl20fOgs2Jk2QcutFoE53tlH24ZuCZ7GGqGehvKO0/UZMrv
JDlrwUMuZJ5Dcq7XM+madcq6RQFqDCEaF95VMHefn3/FpfMAWy0vD08oMDNd6UN5
Ens+DgY0cRjk0eGSIkxAzb0/VAMKjBMAJOAhqUx7mVL4kv7krfcnkpj0s0EcTkI1
Z+Vl+9XTpD6Z8J0VB6JcA+5HKH58yE2iCdS4fgCW4412bQ0VYWFQflAFlM8m4E0t
uoTAfRksp5fDtb3hH7SFBVrRR+5tRUAXOehPZx6begrt4Y/SaO+hAwWoj8dI+gw4
veNLBSEhCIZ6cyK8WckiBy8zvj1eOWnM6cXotEbWyClF6EbiFEfUbvPUaaVkGLXq
PYeQaN0Nj7K0l6NfdheO+cjpziZWPV7I3zsFfHSJrDopRbjhhCvpq4wr+GJdhcsP
9jKvrMCxEJ0TqAMGdGnYaruS7K4K19VrJhi3SBxAC+CyzA026WW5qcPiO6DDNBnI
Gu31LVGFW9ar1AMNXw6m9GGpZSERVnEvX/QrDWKq7qXLEFuloSdHDf7Z1+FEmkvR
dfnzM7UMClcmC/Xp8rAprMZb9SPduag9U9yEBu0FqUeKUbW1MbCNrp3bElhomZSm
fzW889G4XpMcqkcmUjZ4xOQaWo1keo2fu+EKHMH4Z12b2FtLIwghtYoodDrLZ+cq
8A/7POO7TwRbo/IL6pliDKsiZEZujEiIk5GEnXKdTlR2xot1L4r1Vk80j4k20kAv
/Bw8sK2zSuIi4Zufmbkdu+MN2rZMh4NfHn0XwLDa414PyE8q/eI7mRJHGL7kd4qn
yetl0QklWONW11RmM9hh1lkmMCmGpJNructICmfbVE//WgnOuK74TVv/zywBG6Ik
I28qHbO2bVcnoTkYFbpBa8nhhSAKoIb2VopcKkj/yJymtzODwUR4YkorQzDNVQ3e
zNN2j940ja3pfbCzhFcME7SsbyosLuwwdO5G2TU6oZ/Xqh3ZNi183+GR+9OIIAgZ
tAWmS+eMSHcj2L/aGnySTga3sgrCgvVenE6etAbQQw44rb95eTlINpD7NogFEzMP
wNMjxd0aAMpKe25Bem1/CaLHkYw2jNmBnn+eeHQOXSjfAWnlkRLUwE0A27pF5Qrg
alXkbDs9g82VJ+aTBGUFjMsejBFmOmlt3qxjqTQraeOgg6BtWABn/vOnwB73kHgX
Tc3p9Wh30WXaoyZ6LEXhJn+SUTxN3E20J15ejnJ1iDnEKQarcwNociiPyyq8KNh0
9G5DUxsjW85T4d58Q4sQ6Zr8szlaFJn7lwxhpQLoSKCZvTfORrIgOrXUR5YMLFzs
Tof3erJXePKJ3wdaWztTIIf/0D1mqMkX/VvcXZYS8fDY1FlQkmIT93G+LkM2RdXI
X2c8pYCS+QlvCyw0Yz+xwcehbNfcH4C+yohzAb1ueddkGVlcTfXwbAViiZf5fIFw
AKFeDiQItSizicxaZUjWcT78AOgZZJQGZyKuCAsXNDOsthQ8pe+/yQkNmMBG1LEv
1AKzM8ODaErBf1E1CfzT3Zxf8fLt/LoERo5T7ANplZu0H3frASQcvMWQEZDabZLf
lQzwEamPOC+WQW3R9khueZ49XtXo0w0dgJUOQu8ykSsPcWqB8zx+inNS2ZFg8Zhl
afS68we2CvbAQ0JvnCTO/xXcnulpQe5hO9CmuO9zxJlNPKcPuxvZXCbP5k5Cknvc
bmr6w5C3Nl79i4VaK4sysq7Qp/92vFfkQhvWDhinuaf602SJVpSSMJ63jpxj7ksR
hCft9ne5hE6e4Gh2W+Jy8e+5LcHx33dX9rFK47qdMTaoXfp5zxMt6aDclRxcCxXb
FAItSlhCibyAudgnUvuNc4CbWbOR7VxbZmsk0zAAOMJqTA0ZY3ROeXojGZ0krumA
eBlrRR0zHMwb/iu1c5rxCnCoEuiF4sD59H0ho5FwFfimWwAxelQws8pzoYOMcHme
8clkQkA0eemlq8xnPh6ajmRmFRMzRbN1vkjb3V2y3SIw336IZbe9+JJpeA2eX7Q/
OZNVRPhU9h3F7zktwlhUz4cGJDBWciMieiSqUPUIQIIprWoiFP+q7jxHLc0hVgSg
+IrYtXn2kCjgDsyQs1TMM6xm6UP57w0PZOntuM702h5aJwehokCidCZLF3frLbbj
L+CB1eQVUbeHabOilbiLXEzd2W3Zpp/ASffp6HiJtmyND9pJdnCYYrdNAixXiiwZ
CtMwqh3V3Ov1QSwb5dUvThDhN4dyZa5i+q8z4mKE58HYochUbCfC7kR8y3hVgjDF
M/cTrMF9757UpUEOiLSbnxQUDbcIB5i5RoihaVScRs9myBZFGr9e2apOTz3Ci8Eh
VSX8JwAtNW0ogkNDT0PV48bqUPqE83lm0j7Ceo7a3q/sAI0YFVTRFbd/72nnBbqa
KWrN1t/+CFbEBWaHpK7z83hFVVulDkVPlgczt0ZsxP3+Uha7rO9Hs8p7DUm7WB8B
uC+PFcJHwDdWasv2HAPAVhayQRmGY+EZMcOWScAf9a0Ou0h3KGoPQRhalTAAOkVr
EGUkji+39ZW5jJePdOseiOtKaTPYDBrlwyr1K7zoqGGrUmI2Jlguz7uZT70dsMFK
x6Ll0pvr4uOFWossfuqHnBDwYGqvVdvTap9wiux43J4cgOkNRIZwoaQrENS87RrQ
1xcPXwm0fnTM1+5zwCIY8L9C+anrHXSUntJsx6ybYiObOD5fibjZLwNWBtVr7ASa
MTUa7TQqEKL56uPd0uW/fYZE/MWvLXyBgUmbjMsDSPZwXKUPdGtpyTmilNKy9wTF
uv31CPnpRlqwOfCt5vffrX9e+FFGCU3WypJYR6+9/HGjV9mfcBgJgqbwDZG6nj1C
FrldpQPGpSMT1Ku9WczPD4mI+aW1SE1qJc+WXqNm/ox/5UfwtYRFHIp9BxUKEJ6W
j2Ti9xzW01/odqoJyeXMjsbxlTQKtH8dw/NEDM22wLlAsq29eLU1OpBlQaRGd0DK
1CpoB9RxkBzhjtogS9+P1HXy8MSQ/SnigMuMoD2g2sWARTNa/uNb6bLuckFfoSb8
3jL37J3r6bjp9nAgpR4noks+NcfwODWGdEog+DEzaGrZT2d6AC0baIVLyio9IMyB
KXLrzG7ramY2iKfRTDNt/hOTrKdBpKkaUPhcVe/8yysdUGrrlF7ZQ7QrNbzBwL3H
yMNH/oh/lS4nUPcqAPxw+c5WbNVxI9irf9Bn/I4FcZM1jyxZcVAFd9TBpH3+8xlL
AjtoDyPqQEum5/wU7My/uhAZzzsRd9tsYXxJvZAO2a+PZN3kNwXJTbRzn8cH8DZq
Q/IJxubhlaX1G38L8rcn3GRurCRp7CeagCiNXr6PnYTC9WA+srrdJ1r/2RHQZQ8a
DpkaNuXkD3bakHo2f3QlCvroNK9gEbQol5vgl17xZBGevUzloKoKhCxkpGZe3Rr+
db0buUGNSy70zBMsW6CBHKqoTyTvPeQ6ljjtsceMYlnGrDjfjNvxqp2RCxnXGsPY
vqHyNRj6parKG+N8M9RXsdWLCx4jdPLdstLawjnbuj4BW0SPe6zNjHVuMsUF6JUz
CQvbjb2xo3nAKQrY0rVi4w4wdX4F8XvD+wENisWlyM3gjrm/ZbzNU0UF2Uh/7kEd
TwqbQYEu7lv+QbsWmvjmozsUfe3/IuZpAQuEp7bz6ofayMtnr+13skw4Obh7cj1a
T611WV0LBV06G62MW5HHB12fZ/nGtFvrfTg7V9WIdbcE2y0OtdMkMLsaWmPLO0xp
HyRCSS3995pBMN7QGEG8zWaH6pCwfVgtlPQXm/68B5nBt20sntfVzcHDuLw2F1iP
xL2OCb8+QlISkHBsPOU+D7A+q+FYGRyEmiyOkf3yrXVTZfENgZiPAMyO8U5AHrQt
IlWihP8nlj+sZiDeOUusDZHx0gBKIy5v0H4uXi3TZch6KYnsLg49iewhPCeqJYFM
SYD6q3dCXDDygbHsWypy2mM0W6c768OSrEi/yA1ndPfp/JKrr5M7zuEoGTIfZ5C9
xt5Alcd8jipWcCuy0aWoLufRQwrxeoPQN6EzxK/dQQq+l1a0jtc1TnS9Q69Z1DKr
d4uxrwlZnujjYbyC1tFqZ0C9Is6zDIpdtb244gjaHt0wgVplUFtiINOCB81PMoA6
ZwaqzJAw1exw6vzpl5L5NAoR57FPTU37qVWJoT46rEKt42hFpMA7Mu0WKz659xbw
LHxU6LFeEqqYb6kXCZYBC3OK/26nI7AxYghEmarjAlYzkl8ZQTE7GZkDXvveWp2/
0dXb1o/wFazT0viZgKdWEll5xaPzxGnWecYkqoexTxvDmgVPunh8M7pdpZCSmhTg
CyQPVHt6MN3UlFCCopL/RsvFuZQ/ylLf6GhlrrO4fGY3CtokqQ2MyF2e1LdXEFa1
u8FAly3bh5zRI8yqDhVNluxO14x+Fa9Vxe9ZXpJeZaoFY+MdOLhwWHvxrGOU0Uis
MxtBiFdP9xX/7Z6iFfQMnyI75CMU1fHZsJCdGSBpho/VfDMP8DXDtHXTAW1Bm8v8
M24OUMi9ZRwA+3/VcTAMnIkEx8euWGCfAkt2JzjyeAr54LhsDUAPynrYTG3pkPxF
aG6de2fP5/ikcZ/WbKDVhggzSkrstdrq3VIf8rfaFiYg/HGcKLd05Edgqf5A/lnd
/wPlTv6Lg9SPE/EI0re+kP8AMyBrShyUYbjXEEPU2X0GjkFYYOL6IOIXhpHppvYC
XKtm4vNnE7uCX4jqc2mWuQZe0ujxRXmsiorKbZjgy7mqy8PD+uV0gEAR7Y1S1/gA
2ejCRrMtnJ0ap/Pcos8j9fycRkiCrGyfo+3/vp3fUn5eS0xDGlDh4HevkPbRdd9+
Lmr7WMD6ys4MmvNBwi7gNYb/ffwdF4L0cLVG5EiCdzm2APwLpgMvQEZuxCvhQWAs
Y69hRwpUwP31cf60cmv18Py4ux76vHGjVOrPTTrATfx834YxZ1rqv9xfurggIocD
lxu9JJge0tW0AFJRyTV85KTurBSm/PWxr4f8bfJbUlmKLyYgMJ2plWtXztwGUgdo
xOtxJvVwcA8B7QNuj8/e3waEaqfVdw7Fy+mkl/UXUxJ95MlDE28x+G1VCgXOYTgk
znn5RSN3VoXOaGp1VmRHdvgWSX5lRidYntZ0M8IJBkhdxrLXzH+17MUfrqf19uF9
bFUWGn6tcdDBYtAvt0WlzDPKf3n7LJKRFCVqjbJCEx6cCwCtnt4Hotnhrv5wPz8n
4yzZr0PWzhKCc+aB7trTMazEE6a+a+12saZGADjSdvMjHbthAXEPCwuE9YWR99GL
h9rbqDci6FQHR+zrl/pUyqEhBUc1jlGve9yjxP0ZdWtUOj96KwzNyCpHj/9LCwlp
fK+YVdgy7Z6QNn6/4HTS1BA9e6FkQvHau/x/dr2DOX6SXZHtFeMvzk/pDUhcOSPz
yPHvME9dJrYHgIg2N9xPYUwuxeMsNS9rzpHejOO2Sh3xe/pytDmLXZ9bLA7jNJRc
g1jG+DnsT2jlXtNJZlskUtetwDdBYDsaObQtNZxdrvAAwJv7nGWEFGL8KBv96Okj
/WcylI2Ce0WYHJk7FlJoRa2oEcOqRwhQeyasuhnbkpEXNkQgM7Q4to1dIVNqiNCD
Yhyctl+RGSHXVs3tXmZV20AYBxFRZpQsfRo5bRpZztAdlMhkgkME6hNHiDadVV2Y
IrK3KfwQKP6c62UVpu77m+mF3KSwJfOLk2Bbw5mrMX/qcnn3kx4N37ii/Q+LAK4j
OPcABG+bjmrhiUMiZ2Rhr8+gUByAhfkq09Swfbvdw/dYdzUwckxU+o17XnHyd0wh
P1izH+jRdarnEITJZMfi/P+X4a3bCWS+gJrF16BJslz3/SPdi0wTvzcXFIr2rOud
Kbm9jbUuWfUJX2rkqH5gaiex7FDZb2wjcsl/NfH4laL2KDUYgtIN4ro9Z/ikAKvH
kmED98fp3Jj8iykklq6dHe8AwGKpijxIDcseU6Z3UvUokOU3f2ogFSkyKToK1FoI
468LeoNxVP3CTPCllpaxjAAp3Ic1AhOUOI8yabC+NqgPuAJJijAyfxS0/HiWQQ83
xW14cwCxxhk+6IJtLG1LfzuCRTIZPksm8sZWT1/2x5cmVyWbZEx/keR7rdeiqV2v
Sgx6KFU35+cHSt9BEG5jk9aJY/WFcnIrdmtRyJ+aOIhjFEf7bX9zy2aq2SW9yAvK
oRlT7+CLmCCsnvNXFW1WWgXE79IgDyjpQawkwOrDDZpufL8tk9c5Bm4qZDLeLABC
vQx74o5wrcAidUk9OBdsceXFV1LKyC+PlrQinLR0h0jKDMf2D/n0JvLNzJeZQ8wh
whNucZLTfr5Gp7LhaFf3RA+cnNrfEC7+wW29Vn2VFSE3MD8JG0XJ2bT2oEDJEr3I
kWi+bzRRFvwNUyV3Jr1TyPHCVaWDX7mkU+AxMin5z9KH3Yhq8xnANFORyA8kife9
Jy3ohH7czgyEzs/0bw3OkeuNqO2sNgqtRv0Mm2r5WA09GF+GLzRil+JGPm8YDo6V
IPjIT8hpRIUxHGw5FmIA0Fg4Ia5TBySYryMXw92hauHmuvUx1RGywK5TnyEnhJZX
4w1+BcTbqkgy5zOvYzWonLAFsXSQxQT4kMA/YiCLNJ8M+J7tHB7jcYxjVgY9f/xI
4SZIe4bQDr9HZXVXUqjaTsh9myaLRYTI/1/igOVObfyUtIyG4sp4rUusNJN4o7Ie
s9p8LcskTePlpsqYoUBGsmQgycb28wyhhjtxUhEjKm9TAxYgS8qW5KIA/MdNDQCp
02Y7/bb8oY5xcC64ipSF7efMWt7HqHdRwEB2iGezYyMsu4O2eXjwbca/SBH3v9hR
doj4SjnJP+aXlSvEY6lGwVWX6s18HcXlXsHe/r9NEa88JvnSiiu0ZHAev6W4appu
mMsof8MJXgqSXQKFrwJHI0EpVGtFNVcRMOTs2PYQE1Zexf48HOudIIFiLX6g4sTS
iHIfiEr/++Y0BYIXAvPBc3m6FkP5bNVkmG9W6u3fTuPQvAqrpLv1rth7XlCjk9k8
KNXTCHy89ID24bU1ZUQINcaQgp31BwpnPCICTgkVsBjW05k2xwcmju9z1TDXbPll
nJLgJIecIcECSa3vapmG8q/0cmt+MyeNI1jyOLpv+5BCpV3bGa125aHYkjxAGU3z
7ldXuR4Uf6q6W3lIcMIv66B+oVzjiUi4L7kVoxoeMYgLce1Bds6HCggoTfFaB6PW
/i6Iqx1hUt/k3zR4Mgz9c9ae+xh2uuIgtUzfWGRQWccOcyTAQHvTrknJeFEm04+o
pnvgKBIvXpUCM+ktno3KapzrHjJOt/XQRpE2KqppCjlqzhUTMLoEdfA1PZXvNusn
HQ/6OB9TMDmqjarNVJSpBFZmrpDTeHP5bZNTf6kcWa1kO9E5GCv4hnMosczhLEIv
tFhJFdrb73+mz5Eaw4Wt5Se8jzvWan3osfigF+kEL99mFA54NfaQWz0Tsu1rgq+c
/LmM/iF9MBKdxrf4M9f9GtnILCAlmZ5PQY7ofcgjAF8vl8zt6uLqqrq0eFVYtTZI
M0iS0emOugvu5mMd0AUDsHVfQkugZG+bUtVl1JWI/14uuHeb2aZH4e1Ms3LdD2iB
orz7wo7TI1xAbpIf+3wyt1y9aZN/LAALRhzyqlHTcrkOXI1u/VJj8V/RYLU+RKew
g2LKOqQTYzOA8/hj3DFsqBsXus0GO4/EejZwzrr7RLtLEgbbZkZSYPMEI1hN94W3
Q9gAl85SIqkPmQYPrc0HTbJ38wI1kIkcghkDp3O5mZFypt12wvtqiFOujP/KcD7A
TrZVLni+PwwtmWOisXptdCsF7S2dI+a8E1+F7E2yMctauK+iCNosGOm/21igY/Z6
UczbGp02TdG6Wv1S8/rypaj2H20xT/YkgXvuHW45sZNYjDORH1dUhURvNbWNITcY
Ml6k5uSsVgv58U34mDcX60a2kM0+ETGGp15b9fewY+WGGBqXkWyo7N0kJ12EYUrm
fN2qZ8vWP+obeNmW86ytXPLArN5rssac0ykGoe+0CDs4ARMn6yRQx/ASnQveDWrA
635vVCC3ZbvVmi3IhFNgh5q4ih8GJQ6cQp/IH8PjoLE1m/8J6nQQ945LUkmuHhMz
Fhizs5OutVt1iS2lBkdViOaIU/l6Zx7iWLQIjMCTuNuLJkKfatezUs0hD2ojI+KD
QCFYXY/KCIyphaNSVVC30oMOA+MppCHGvNnYHM3bNBmDDwSV590KwUjnNe8dDehe
Wby9uvR16+agYDtKsSzqPnZl+l3UaKbuEzbTzX7iW8sR1rf2GkWduWgfNAIdS2sV
F5vkQDonMrZhJ24+o/s3ZLe5LaDbDQWHk4dKjSg09iwM8Q8rRRaxMNhM0m/ZvCe2
N1hnsPgp1xwbfbSa2PToVGQmlvCe1GOAgn7nAR868urL7t0usEByJ/kUC/8vcxge
UbIfhEFcMhpZA68PI1imIWXg4GxcuaaGX+Y+Ugm9NNVKXD+Jq+eXfJ5mOx06I1rx
cGqs65oH8AkEYZOPH+zJA5Blq+2YrSKhVp9OgeGxTxwOSs4eWaTa49vJlpC4W04e
df6pHhbxGE+BBh2JpHXrNCrYhnX7QOShcb88rAlnwCjvBbuD+aw9x0zt6fkShH9o
itfOEdxOjXH+aI9p2XjXremBZxuncy14XWsf1/aSfEqV3pj9iESt/b//LrZJkRTU
nq+Exn5ayZq56bWrj3bURROi6OcPPpzLJV4+LETOiN4ELibnW82gYauKR5cyRrlX
qLxN6Q7yuFGpYFEegoSVazLmEmATpKtuZ5v1KamFlm1iQ/tTecXWx8kgrBrfhuJh
6aWTIPI9ij2vEISpYBMU8hATRyuNJDnaLktvaHsfrc+IUC+dRKy6ROq7NL47wy1E
v9EAKE/YhjIs8emrOcY/OB8W9xaBrOuWiEu8B9XsP/eBpSXHrYRwjILVtmeilk9y
erWYwfDb2J/P3Z/LmCpGwOxtfXeOa2gdQlQQkhc6btS/WAvjaYF7lzTqxcClnM/A
vlD2wRKt0a50LCOAXOrBAOPgI/CTLp5DB01gwKWLSG5PctNLuO8hgO4fiUvJq8Aw
hVZUr5agzrMLAkzDON/c9+U7C0NCXxSnll1eYQUbnepEfKAMIJt/9miIWgyhYzHB
zDLbD3zsOaeHMXDeDfM2jLJ1j5mpg5bWVgQLLSD/L3m4u/ItoUS70AbjXdqKNp/J
0DGxLZBCD8UsYnrvySU4mTomQuxuFS2I+pk32oo1ZOO7ywxlnu9Stf4J/2al+xLx
Bfn113cedKhci1e5p1jMl15pj486XNLvby/o5iEFa/OvDAJ3+76lYtvAUU7vBZhX
62BBWVR8Hg6IG/MzVJTOMToZnY30YJK5aOX+UuvCIxZjEBA7CJT2g8yWXRC2HI8i
Z/rJzpMFlXsrM7JmoY8KUeQc8F1+HFjZasE+46H9Ax4JysLe4EG51HY7SKn4VeT/
mGmIdGAFqFvN1OHckWw1kxcQcM+WN+Kolx5l6Xt635EGFkFsOgNbYa+eyR78kO4M
J0oOCA0ASczpXkjReccfUc0V3KKoEK6gOnol89tlGgF3KlZxpQyle9aPOEw+6JNW
j1yCNAKR/QYYe2gOgr8fErtU7T3AgH5cYyPNY+62gawfyZI/mzEH8qqvzKHM06NJ
Z3tKIC/Sz/RTvz4XQHwv6dhlLlOQpjOIy/CPlyMeYnQYVn/qcvE3U6rTyURvyLs9
36aL8tsrOiwpd6WfMdI+WUJwTCpWOX3SAQWDsYJbcZVmTVksRS4RT7mz22bZPiZL
09Zxi/iaDnMFFWAiUsOsJJUidJ6rmISGF/ycqLsw8U4IemAXCCVOEmUlKaIULmYG
S7bhqVgZABYY4Qo3Gy8lmzJhTk2ozSY+8G2QvvtnoqN+PhBiqPoE/bMYzF68s3qS
dFxV4JbP35zd/oqeJB4zjfcQ89ZeljPmCt62g9/6Ayzo4m3SVHkvz6QqFMssKJ1W
ZzA79kWqRonMkMfkfpHNWPLPhD68odHzdnW6QZ5rG31GjJEgdSeoOePChHKxt45X
VYCZgzi0xGmExVRh5uKSOPAfiqx83v8ynB8KCFCk93T9Q2RoJRM12zqAJOFdGG95
f2OKSAckowUCioZNlmOhbTp8/oR8jXHiZVgY1muaQisdyDtYZQqtnwj3VzLJioDt
PdcrS1PBT5PEpHmwCSmQgRW1t6iAKBC/25ZzlO+5Pu8IIaPUgXg+bRCBYI2FZ2fK
9s0Np/XZWc5EjMI2/hOT/rpG2x160kOBVW28jWs3UFfWU+rFsqeCx8esOJcMQxL8
p6Z4PTO433jqruAW4DHGFcmqZUVAPTonUwVfzIKNHv5hyg4GsMNc8KyxI5wWGhJJ
KeQvRJglODGFaPJ1jDLah5ONnvGbJBwvt2d84vzXYDBSZ0tWr8PLqbR5gWSf5KyD
D0UIznD25FswxyRErG6aHzFVfcyDQol/SxZ9EDQzDXjg62E6l+b7mLP+WjRLNQkj
9WcFOC27oW99fI0sc9SVRK6UM3mvmDw8qocrNKSzSl9VK3uyRnY43pFcqyIuQguu
M+7AjqacMs7+saATxDh1OhpiLJX8HwiuBoxr0WLV2EmtE6kyjvSUt6Wx+4K8yJEb
zXhHvSMCEuT0/kGoDFdaZOgeynMxYPKPQ8YWHFNqngOZBu7z/qkdNbXVAIj1O3SR
J3bxSXWl8v7DhRqPeZADoGK+c/EjjOX5q5xz27oG1addSb0aK3r8eKiQCLM7xv5R
YJi56WXn4rD1HUBxbhY4lNnfEcaospOzAyoaYhP00m0KGY05IfB/dencVnxZxCUc
OU+1CeOjeJY5AJyaoqzwJZeY+9ANStNqxYemKpMYgOBZPteDFRw9TGseHnFs4SId
R/wP2gMjFA+lR13ZaVKVdNY7uaq9+Cdg+xpO1bmZq/X6FYW+PZqCtko3WqGjheZD
G2eQq6IUcfQyP4J/YTWHmB+Akw1U9FIYDARytGaQT2ilVm3UZfQsnlXcGU479Zkp
mehlS4Lzjp1dDzjiMv+NjTE93JYc07zAoq/Mq8GnEt0qjjzXohO1rIOhL50OlVUi
vylYtyKX6HVYDPH9liHd+GVzCjTkp2ha+Q5oNROsi9AlwC1y2llUMz2m8ZEGiBVF
JtNV6+TOHWjDm1cLjzATKGTNEea9AJiZlYKrcPWOaiTKYp8MWWpMHcJ54p3VQD9K
TMkn4A9oUdBSV6205n73SzZcgu05m5wcT7lfJ0fDsLoolLhs6MkKjmyOskf/0X8l
lrIrwkWALdV8gpoJXvyiyyyJVRFJige3uHfyNbFsSFTaY9yft9cRHSGxhacvdy2X
On6kqcoXNC+mI36v16MfGTXYE2Ia0262QE/vy6rbFobA3t7FrBC+dnCy9IhE/jCf
RNxFrRNlyQVfi4kcY3RG6WbgFJqdR47AssSUM/FAKw6/xyJ1ffQdS8FTW/3mf5k8
4RjzPaKjmz7gl7z9zL3Ogn62Z/iq0N2M2fdPHyblY3IYAGl7gShOIVssHxqP7NXp
82k+27XaUbRHvNfAMzifRtL05c4pWVlIwlrQyzdn0XsNpPFq+ql3KZbaVLVDIy9Y
mQGVxaLE/8uE3upjpMIg9CvsJJrzPKZdcUc1ZpqRzyxzOIDHDVw/Pa0DHne/uJNX
68jjK/DR+p/feV/KIqjVK/xU5FeI984zCrdvqQgT3s59BR+UPMzyNe7BEyzCgvej
vVkdwDjuP2f5r665DvIBTthP+reRkZjR3TYCmJxhHHP1hza+M1MXno+V6n/JaHi/
R6teB3bKQpvvCfRWtRL+ro9GAr2wPbjzDUd7cgNVSu4mGzkNSTGSbWZqYNAh1v2S
XceipWbY6SKgpHc7axw6Z+P0jGQ3hp6BfrNQtt51IVrqCCuk8bgi8YEaZXUttUGo
9Z8tWE+AQSyO3UzL2w+qvuokbPEufEIswuZ5PVcTMy15AFm+gYRqCbTLP/X0PZvr
p4++3iZL5l2lmCiAh0Nl4G3KT4CbUv7KRpwEkzHKUfkSujphV4muJSf/DQayfXuW
Kqu99+WUDWJDKbXD+xtImvkj480IaQSMLrMGWajkIcQF4fK+M46NqE7wMrozlaEj
TiSWxEfgB7RDqUhvC67+e3kWFvczHiW0VEcr1NqKTuu0WQO68s98ZnNC5MfaLADt
zRtCqVStgeQXY9K1CIZpZ8RlqCVLKA1CZGYY8uuvYDVCOoa+7PdHhuxToQHPU54j
kPlYaVdlSqJjVrMgImGm9UX21Pt29iG63u5LDSN2CnNn5aofnYEU3POweg3qLFLl
QB2Bu2XErb3YcgZtDTy8TSkUih9T0dsQYN0++/oC5z+Ufn4Y6SkxN9jVe1HMlW8Q
u5X4domp46qIAbjtxpiIwD3kVQcQEQqD+G4P97z8elBYi+0iaaJJ+v4qtPY8T08h
qCmIiejM1vTx0KYI76EhmOk99iy+wrn/iFkDldcDthKvtcWPW59BixvziRoLG0Xn
3Xjez+uGZTCzw4dkI4UQht/noi8pijdliC+XVeUURaGo2kSpuKj91EtQmk9JSZTT
wm7WVXiYRL6KW9v5FKgTFWdGrMpZXoWyk7eYFHARXlGSo2tOBoHh5+3fsjNBjA9I
JGQ/Pl0E+boN1xK94V9JOmaUFVWQzLXdt4xc/UXhchDYUsBznD9hyWU/8wksxjJq
4+MyT7UKG2ZSL8VnuIjThhb5K1q5EEhgqMWMrB+klO2QjLov0MPfMqAw0dR7zcyo
hW9CA8+58PE1iCYsg6uoDZwMsTCoz+8NhrRkgqz79H9hSIyXzjgjFu8ylG84pB8R
psuOIVVFu+pbeA8CNfxnGIqwpM4G1dhu6wCjDSA1kR5m27l7qbOwN2AK5+/F9M5R
5x1mIoZ/PmA7rPo58GMN1M7r4unfflgIHZF6gvLIWABZqffGlhZzeEDyzt+SccZd
f0SfyDSwa8GZcZC/PXOzQnIkFqjnqyZG7GlV7vQ+SB8En2L5jYGz2GTjEtmGfRPe
QGt73h2vFh+midOZAQdHVh9vIlFXSTbdJOUP3L6gxiM2gLas52Ja+ETf/58HK4lo
x82s5vPX5Xt7+WiMDsCpzhn4LqxRHUfbBj4p1jLlCsWyXmYLZDNBdefS8+Bli0s5
zS801eiaFJp3m/VGPgNfSaXe94EJ1TtBy1Qqc2bXqrytwIFY5Lyo8e6sxImW5cbx
zCy/2eIVtQICG1YH7VtS6pyh8Cn7vL0gFuKd6GQ6pRLpgMmFRpAcbHJrWxyikD2q
TDWfEv2yeuIfDNrOuKVOurw00wYwN4Nj+9kvtKeqgW5Dvwszdl71mlq+5Vu9PpOg
dPWzxLhq2bm5+ICWBAHda9QDoT6wDFF6fsvFGHJ6CXgue+1Ruhfv9FOfmE/+MfLB
cF6i0JAleW74KSvV+SffSrHYA9mFIZfjnK2GA2K+0T2qOTZDBtpmrpN5+mAV0TAw
0YunkYEJMI0s2SuKZ0BkQMCQKTXqgxpt85QIrjXlKQtuCMGStTJSY12Em39JvQCr
tcW0yMEFbvDhTCxT+wm3OAv00OUKk1WOu9HGXazAiHXVMG1bMMN9lyYf0F8ii1nh
iTUSlty3m5Wd3gA0gIL2PmZK8IOp5N4d8mmO7ESIwTBiapAr1BDoDB0YuuDqNtp1
Y23YcLT7V87ULT6ozyIPRJ02ZcOsahjDMSoCUyFKNpYNoANPwBpeJr7/nHFvEQ32
Z+YnXGQITico/PhTOeRsLkY/Ur5d1WmiSrTF2dSNpQ6EeMAP44o4eWQ717t3KWRg
OORnguWIYK4CwU+f/bAI4iRQPrz6cDLhfQIzARkeHw2RqONZsSVuv+8RKlwsVGgE
CyTTwKp/S0zVGc4A44ugguWu+Z/3VO5T/hBFQW6x4vp9f9QU7FpI+X1PsYfpRKtf
85mtHGuREgELu3/nBe0nytz+5Gdw1h4P1WH6LMnUBMxdleXLXfiSVAFLrgmscoz0
CCXCcC5e4AV/c1iOaJxxXoEDhfi4XjpWdvz+zvdFyNs/4DyXc3z2jiQyqUYkv27P
m+bdkpBFVVsumP7crnEU7W37up263o/psnldu3fomIA32MjNmD+/9PlplmCPKZIH
RE8xQVe7LeZy12+cQX9iepKhGaOC40hlRfVAmEenc3TLsOOMt/VUD9yIixg8POyI
OQgr5XM/S4OfnIq/HSZonwhjQV33kKr/RKCgQH8PYSh7tG6gPE6NdrUq3PWPTEq+
NSso4eSSGlM6bMSsrKxyQIJ+oQdWU7Oo0+H7JcsxWcl7CkZsZ8LC5uIVtpu/Gi5U
WSgFSOSbA3/duwgoIbolkoWWrZAwB+WTxjIyDLUAaBRJHSzGfkPpXSAwoypoaXDL
l4Z50vgOEZ6hxJ1aeUgJk1qUUZAxBcputKx/CcXZg5AN2gBGuLFE4/ww7Z6N+lM/
s0iauZMKwSZQFdYzfLCmT8baAMiYPeI0wlT5LeDKBrTINq8xDwIlk2MIClL/CvT4
Es4bviX61RMVm05PNbbSMKFrpqD7r5Dnqx2evxnXy45tFgqJue0aRN54Z5yQT5tG
LIUtr0KznqeX4al8brI+rdZtreTE6b2dXXPcVFZJaFeDIyHnfQOvAKrnbQskBxXG
uUlEQXoANT+xVG2FC9KWi1BRbYb1be7nQq4UZWj9Y8joCHaP0cDlviEZzBCVc9ZA
Fy9cJ+BaLWf/X3JDTNCGzrqGxAfPycEkc0UquMQfOhcSlgyw3bMJoylSc7vIp92X
bs80vC50tILiZTT8f+a9HlarKbrniH1Jyx8YLgGMi95k+MtrwI4jG2mSmf4eijeX
V6wduhiXNPcsGtPkNobYRPZtEPPZ7YGy03y2IWR2ut8Onn7qeqoVTVCVgcjiQC+w
4NIUI6T65/9nr8CRapbw0auMoUCk67yoVnb4JTq9y6/xpkB518IJOOY3dLRJT/6+
haS+EqbE9KDW72C0S/yLvGBhCcpoNjDdlvTDSKukG4C3ePaGew6Edr3mLq++8i7O
5D1zhJqNUivLvITfuRn1ihly7ZcdwJcl6sy3ka7LJJea/Mz207cXlkFFhByN8V2r
SfreGtCPQp4pTJvycCdsF1FQ+NIXkB4IfkcoBSCIW4b5LARHdSq4x2aaRGDkTMuu
KLakmKN0+FPUo5m6JDT1USL71ZITpf5dft1plWxhrke0OQcXHaHLBjPEnjh5eE35
YivZjQMkOmeypO0x/rUcW1QVYa4sro0mOlMFgxejnU/zUsilr9Lq0AgZqG4lkyRu
nvCFAtqgTjjfZihkgPYq5wE3ObHUQJ/uydes1v/VaAO42j7wJmyV2jeI3+KzOrJ7
bm99vnjndBYjIRUBwSV+T6/Z2b09ftdF1bD4mDz4RN/1T0HJy68dndJBQrEu/AGV
z8ub/mSR39kQLkBnGZQzTrLEiMNykwZBVZg/2q7Y/2y77ZJXk2Pe+XhpYMOWRTAG
T5SImgD/cUAVYlJeh0jfufbxWcU/nTN2YbY4ACau64fWhes1Z0Hm0t2XS1T3J9tj
4SLPSsY61z4x7Qy83vh13oyKpqRo/5Jx4IkXer4MliaCoZvXHwuERLW8d05wFCg9
uFHIOg2IU9dRqUK+ozca9tFB4dS7dVFdrpn6Layt2Dv+sIsd3fEBV9VUqnMbQAfr
/djz/qOmLUKkJ4oEQ4Ry20Ge3YZOilvZ7zKHSdibuttOnLCZzHJIl2GT4X1NPOqn
1atc2ZYjKzo3zA1+zTVFH/vCs/G5yYgMzV1+1inRcgFNrGh56ae2q4pI+F1eOsDX
/SWKAvU2q5Lsqq3BJP1qA413g9i59qfvWEoCC+RJZee62cJs7DP/SwRFBu8+Be8J
00pO+StNUN6NHjz8g5Mg10SXs6euG8jy5K58Z7vFlu5+QWor3se9ceHOfb1QZ04u
W+s1L1DrvWZ/IDFf7wK7k+ml6FjrT52SwIss6gQS6kpv2Du9DoERd4Nq+4J2G3Pi
h1b9rJyGoNy26GAegFaUA3xe2pLZSbPqa6SpLGJ2UYduNlJvl7S0VnB6gH8YvV+H
gRGVzvEU5UUEMJ2LyfqXihr3/L74smWnBsl58inRNW3RqPm0xh1/yNRkK7qVno07
0jnQFeVGwzi28f0y52l/Kuj/94qdXPFh44gbpjAklniesFG0KC/HJ/cXC8gJHxy5
Vm+btVLrwhliLIJbXCBg0QQQ+z61XN4mtwlMBtm/HRhSy9K5dH+WMueuRhiKCj62
PhZje01LX8W3+3bNZw0bj8cJoszMuNLbyPZw0ZvE0yTX/8oe07PZJ+D8OxZ+8uBj
76KUlaoruBQD4ttR758lQ9++UQyRj7VBucuNO4SMBO51Ysrx49gbIG06hpVzIMIr
9ZybTq5xeeKNYdoESt/JhqPjiqdoKVJr9Ujm+SNilGqzStHJgmkYYbsHkXwNbZv8
oXs78vXNLAJ0/cfGXXbD44BPt0FchWkckruhi2M85qwZeZVHjxecayX++dUagjz/
01iGvlFkv5UHAnnpl+QNHbYCgZcbqQJFrfJBx913v3Cx3krd20460ZJHcEcfLGpE
zsaVA2uvYt0w1Kqmoq+wnxeOoqpA5iUGx2LyA3XIlNNlwQKqjW/eth6imF26EPd6
a5WolJfe6Tv/3O1n5oDlAwbAH1gGQwsSevMO3z/pjJKJ4d8asNAthF9buhDZ8Uuz
IlpTYHwWJGebJMuOdYDKm0QDeetfroK5hwpjtEKYgcHwXPpDvKiMx6rfNyjv45Gm
Ltv2lqpoKRHD0/mBjZ7VwPOWMjIPdJo8MzyA859mC1vo7Q7hn64Cl1McTDXMrljn
b1SXilxCKCVQ/7d8pUEACzJBUS13tq22tUsoT2h6AQ188mFOX7sZ5Lc0Y2HMp5wV
5sNdkzY1s/6FrdSwgnHaE9d4Z56Ao/PUJvixwNZMFyx2XqGar5LhLSat34Vr/SrC
ldPCq7OEuAqMRosfno78M55BbCLFR18hwGc8+yHvvco0N3Qold4JB01naTw/LuTp
hm1HP/0RVPfTPP54cI+hYIGM9VCgsrhEQZr5gLoMNfMGyMaU0wAvvAmXROD9nKB5
5NMTzzQSPHB99j0CaZLE914/qKqJT2wSZKc7P2kxgOuebFs66KHVCTVT34/LKMyh
8uIPA/0ku070XrZTlSiL0M3k/NV3WI5bH8zfa6J8Hhd4zDs53WGz+9gQr0+8g9V3
Ksycyx4f+o1JDKgDdM2oeF46Fj9qFKBhXf+IVDNRa7XNP77ybdRg8lOC3YQY4rDy
nDkodIaCTB/MCmp/xnbDFN75dq8kxktbklmKAvosUnLY/O2Ad3sCCRIzAM8fD1mx
0KiP01vOpvCgnGfER9iYXeAiwh8eWfPX+2hxwZT4p/9R2RcV7cBZi7o4ToxJ+okM
mslmEFh5Vcsr37EwTpHceJwW5YvG5zrkHcdi9J8PRnZv7uOhCZ9hrXTVlmOQjG2f
6XvaMwW80w3E7DyLtJtgTrzTC42kYWmgYZkOz7RxRgLYwyEk4oTcFyO7C8jg6lBu
89R6Ojh4gMVzquC9g/3XtTBCT6y9Pt738nlJB7lBS9BMwsSIeitVvZbyeG3AZbzz
vQOBxmqzPEBuUbIxd7s+++++spxR60vevMAuarkSd10ReaBH67BFqG/FgrzXc570
VJuYgL1dIGtA1ebHqhCXqhROs78gePbJmpZXR2ey8xq0+Or5BuPGXC/tM93/Mh/e
XDZy5DQrzM/TqDExJrIe/uXdZMYBBK6i5zEnlK1dksIZ4I288MbRqHCLOauyzeJQ
eqCjjYJX2P9MHE6kl2f/XR7x6zQDLfI+DhwZo0tvqzzI8d7RPG0iR1w/JGkvGB8w
6SJFq4+dp11CP+7F2ULW6G3S3CsdGVUXmJmdDS+u4Jrx+MTEM6lFtzSh6jMSWxM/
w34Bjjn2nZoPHNMMUzDNs4hooT1FxamuL6fxUIOPMajc3gHvJB2kPbBjVeszGVaZ
oHkxQfC13MmJtGEc+8s5ES0o9rfhzIOjXTCnV1d2CeRCNY0hKBVx8UHlkkF25zkV
uI3mcZ14aF5TuERVIRRTPhG39Xtxq8ALGjqqPAeweBzeHqnwdhVXFbXxhSiLRlV6
6oQ1bnfeBSBJagtpJwnKplklQlpQ61x1bwF2MXFbezdKbC3QPnzD1fFNS0RrI1s/
4GtCpC2n1VKZE9cIWRghafZ8Z3BTcLa3xKhV7qKSR37JrRR0w0y+iSHaAFmMWfKM
rjJLDx8RmI3MVkDGyoPBlPjbr46eI/11vHTr0q8jYzY+c5GCcLT9p/qowaNGYfco
Tb0tiwRNpIOvJIUUpMK+VkOnDxsx4esw20guuv6ZaDs8r+f2c2Iu8W4MzA+Mtd7f
STfGQryjfccCwvmgpCNR7RHdnM0I5pBDoL9KqGQlGCVtUfvOREKDf9HGyDmnZFrE
mMFbAs3i+C3kQnQEx5ZWk/7cQyv8rEGmyfO+dcM8qQVm6hZMKD/cQNoOoVtmEmo0
PRYJlFm/9upTSsiEHYv+C3Ho7530JDZKJLHah4M0CS3aWZixLrxPaKc18t/ntcog
X834mwb1TwLkdCG3gCOnZfTIcNpPBbe+3VedZSV/A4u9v/oE/7vmAzkZtb03YhJU
Jw8XSF0SE2wjcVQmuIKOFAN+yZM/CNvIb8F7TMTL7V6n/zQt03UMa2PzffBY4TZq
pnP0EkpKz+s7Xfe89erKFU+wrQ/KNWFtPEY8tGktQwuxbiOmZo7FQp5Aixf3s2J6
Hw8bapXWoH32uRfTn4UpQrCEp/+hkgPzj4Kgkb/pV6awmVY+JfvHUEXU1IV7zV9k
ZuwQK0PpvuO0QMCau1YLsKZmVIAtI2LrZAvO937pUKZfySjuky4EsPA3P88h+TMU
WncJAQVpquDwb4NVEeOryNRpdvxN3WYuBTP6CPS7GIobLl/mhcO6mJW45s3+6voW
7mAvrG2Munb6KFN1/fFydC6CCifrJ+qRsvhy5xfdiN3x7nJltEqb1xdNvLqaARUe
3ut7/fdW+QHuqEqLhmwBZZJfGNOWSbDHfB7UZbcZypZEGwhDiea8BbiB0y8nk2aB
vrgUTeQuo4lXp4iL6XAgS2YZUcjuWHHlJ4ENOliKLx6jIxRYS/gtui11eWNxDsI8
IAQegvTl75AV9hRyxavcxadeN46ibwYJNuq+zbOduk9QuNBnTonBnsunxLiLwTqN
OzXbVySyP4Fq8wicTvyIOBqJyhzns5AWC9ZiRb+F/ynf2q27Jo+OFjkgtIH1x/ug
fY8I8tvYniRDiORR4dvZtTn4r126yDVO+TaJTg8ZV2sCMUUvqA64fd88tdyzcve/
m981P2k/nZHLOhXyuGpKzLPu3CKU9+dgL4dHgFOAEkDydCpvTN88YcvkvapcToEj
jjfn1xPbWR1J1eIgzlA1MMlmSsY9kOn5/+JTJx5qNf8wzLC9ubFRI7+K/vFxB9Xn
ISypELXCdda2b9TOLCajtFHt0jDcJ3DLZeYaRGAsUuEtD88wHJ7OfOcTz8/QpMH8
j8Q0Di4VN72A+JkuKOgL5TCFbL0nLkymgXALAD6flo1lVEp/LgwYN/0/PjUVLSvE
f4IojLRWVFKNSIp8KTaW/FYoY7OQR1pGJYpe9/kQ4LWPHBkO2isXzdKWqS9W8bJo
JMv/Zlx7bYwHd/O6fydp5JYOxj4htTUSAJyr5A7+E+WES7kp9SFYKFfcwphduwlX
oIcUD5PWrhyd6gCmvoWi5QnPGKUlsPZUs6Scgl2lLagwzTpeFCDvGg/teU9Nw4Uz
Y5+EDjpoQkAUhLqoSA4neeaTHvrxI2NGWLH8gEP8Z9X3ViQSxHJ4C8IeSam2cetY
vwZC+waVMQi04v7sq9mRQJoXsT/8d2Fg7WdVF4k5RNw6SgBaggsb/87XGcrDFXD0
gqsNNHv+ZY8d1fI7qqX/2dJCRNRaE4FCEmJfkwQnIq6n6aFMjfUpgldFTmyo3YOx
M7XlwzuG+UXTnnNK+/SNTmGrktMTNTgaXQdn0V8qGrrGNpt33Z5dXz3RPwTDz5jK
Vp+EAmMC530HwA0Lgn3/7cWeIabo5xr0AbFJmOPBqyoc/lNhrRitH2NlzVq7Wq26
39JEbeM05HW6WoCDwd97NuBNfIpzPF5RyLBA4YGyxAg1AixLCp+XCZY4QC7IhuKU
+cqv7dh+sgqQwzsSA7e6vreJEMZ9qfzd2aiXcxOVL2T+t33ATCKAY22HSe4Q2fUR
udnb+rRWbLKZCZ3szzPk6Q4Y3E+WL2j0fzq+G5k/N82/+Uho70cCmE6NCW2nBFJe
5m5M5PCWEXRNL6tFqaYxxZ957Bu3epXhnLIv0AXuRbEELl3N2yZ3BEdBYNdrMUoy
d7rg5YsOTEP0c18MHJad6IqadaZ0A+8M40H+a2SeQvxw2hJNPz3i4wJDNb1eWAp6
ifjiY9RGudWIK9vcEWxChQjxLSsyKzD6ehyRlnaeXDVt26+7H//cNnwGlXkZ2dnC
0lA9vyEpuAhvlZ1Cn3GLuCKc0oMmU4CLqdt/4tPj2+qHse2IvGFu+855YDnlrIZL
kc6DLKNq8ctaCFcgRj3U+7AQA3d8NZDpTr0R9zEd+Eb++k/ZUQ0b4v1XjVdcWZdZ
Yppnsbh6HinqW0F7thwErq3muwL8plIYvdeEPnhlkaQ85eQ1H/liZGTMRmmRaFsM
xcwUVQPd6wMbJaqabbuf9fYFnulA8U7ZcT1ao1jjT5obPLt0NoxZ01eBfhvMAHct
ZmrGucsgjGbFMtJAVvhaE/qFUDIlDbf4zsR55VDTyWap+Twazo2YCyBifq92iQh7
+XEAdrC6mmWfPMyWK2SD+yHLKQjgbJITKRlMxSesQFtr4UjQS88d7J6g5UCL8Xyc
Jeh9UXk5XjjBpJVtbDZuyQXZTTpo67bbeC2MeBCO+P+vuVEXzBjx1PBhXCGtYA9s
3Ek/S/mku8ykn9Vt8R5LzSBrKzwpkSzWXqCVWMAERFTN+Awr1nUEPWPpVFZ0xbw5
LRGXKg+udRfb4zjNmXYP/xJTVsWBRhnBHn3SSBD3srlUf31wnHw0mmb/0tcyQFZI
5Sm4c2qXOlSU4jcp/Qukn3dZNq/cZuIRSGUVJv3Cpe7uju0SOiqfSOQ6dZbOUpDH
BSjMdXby6xzSFCZfJ+ZFNFusHWxsq6DnUOI05GM6iJXtCMioMDBLc0WZldmX8Nfo
ZhI6t+wVr0DJJfNH4Elng14KmRV6HiKKEi5YC87brN5GETzAsidAncwsi8l9VDGr
XFhWuphEYSdcC676N0ndjSulC+w7xhlxCjl9PsRVem5JjL4WN2FWme0pmB2yCbFr
9Amuk6AMeNVazKjN1IxBwqSvJbaF85TSywu2LBNG1tVBoIr2/rF0vVTgUp03Vzwg
3WhCw2F+eJyQtuwiHZ/kWtc3tTKmrAE9Nn/zO9PN69n1ppgR2nYVQUVljJo8cp5b
ph8zW8AtLPWLIf4ySiOZJymqJZKP3vFATumWoju72vyzvTUlHVa65Sqkb8/u8HMN
7q83RnlTmbdmkIrVDUd/mdIOL936BE/ln9LOdjanr63wjUpRYR563mAVCpC5IGE7
YDKnhG2d8A3ZHsPDQg7sK7GJPOWjtznu2X308gN+52WNtXBfFwcYT5QAN2Bc0/ow
XP9vdIyKzRbCZ4nwOXaZcw0nY0NBC7nAAzosyjg8AmT59cvyWojVD11qECiyQMV9
2z+GhHvRn5y6Rctx+u/2Ngtjm3fil17Tz7uLdfC7kqcHh7mDzltFI/MO3oim7zRD
KCSvdpb3+qmqBXxS1IjvVjURarNv6xwEBaw3jHNoG3O0gPbYv68eX+bOC4G6Iul0
G/iDS0p3ouYhotr/N/Xrb2HmAWVV4CIaRo5E4Suu3EXlKi+YKP2BlfJgr9jcQIhN
2XR7qSebk2LGIQSXTmGM45xE542+CIUIhnxfVBqTL3+u20fK8dgS6QJ3p5r4p2cA
wkwiWcFxv4Upvk4f3catJtk0kwtYg02aHZBpEf72D6zjegaJv9tycCpsbQP4vPjD
cbChI/XCOGvZVkZwsAdaOUP+P+uocrNCXqKTdrzgo4N4rSaYghrUEmtSGzjRwT1s
flap/KYEpYezbUz06ymvnFatgerGP/iAcwCY6ecUn1E0GPDpibecNrPR4bjE6bEC
pwJWETU2N8OXNYK/UEO785yF0vWQK/wgahM8RMZjQ38prE83O5+d/5VqpK2eKYPv
zQxWCuukTHkb+l2zJnGHDl/esn0fDcujU/4JIXBbRWAkEvlmTV5IAT+VXzJthFw4
D2AsOg75MCl7ElXxGsyxHXLf0aTfwsoJWRzWlEouqfP/yqHMvHCMm0x9WN2gNfXf
fuLdK+GuHBGMAFjAdFmdvMgI4F7rhX43cnrRAWIYKQoY8tRaP4qqSmzEMjWDu+mL
bdbmchBfBEDA5wIgPsNoPV1RzCdgNI7Eqy+yGN0qs3+mgRBvzyCofawKGh+6DMns
gxZyD+cguXvCO1szxlWS0vN0AF8CVfErMnXnRMkWskz7xrUAcx1nfqyxhShmvySU
5rlWLjPx5nAbiexY18llDWoe+BRN1AUPJvmtP1z9lcmM3SkEVDqiT2YTnIM+r9Vb
MN8sm5x5ncD4esfnkDOONnTfTCEmCnZcFlzubScdXvx3lbE4W0RDso1iY2kLEysn
tQMmUR//PY1dfTNM2kqcCbnMz3jx3jEpHyUoElzNAvMokOm7GCFlAItMes91sVYg
Wvk+iyii8/T2dMTyNETVNft0nTs/+A8Mi4N5glFcwQK7M/nfLU1SamKgXoQoFTYa
DkurRlE1zLO4gJdKbd2LfE7Att7eWRZYAFSSlwV3GheSnnK8pUpMa9auUvgZghx6
nTCpEyzV6TmvIczhnCvQz61zI3ohg0y+4rLtkp0vURrWtQ8iWWsoQQ6pc6jDMW1v
0CHZ4L8P4eZ1kz80tKAYV3D+0/aq6gYnvK/uko++nrLa9SOiLj+8NG5+Dj31z9AM
N3E/tieNh1oX0nrakiQhqtO0SNHFPyzG/bZIf6shVyFTJ7eO4rienMPK1E36WMXm
JSPEuHyShRKT6YdLuCn7xI9LnkZPfHV4hHh7IIz5eNWEPQsXbgytUm/q5dKbfpSM
IAeosqyF7JDpa2Ro9nhIwBvo4JAUzOsvoPOb9VTVgQURfsqYSCaadwISHBfnVnyO
UQasKBrrJySNaIGDwsx3wnYsTfPA0lzEO2lBAT2mv9M8/uaQg/CQeaW5ccPQlhbP
FUPfbJOIneH7Mwl6k/gqdjnJrrDe9iNwtKBM+Jnzi8QgqXmvsx9sHpqz0zFabAEq
iKgMzgLjr6TBeDqny0SeflgH88dEAJNv2oLne7U7lhVvnBpoFtRTMKCdUsnNHqJ6
BKfHKTeeKI46EL+MrHL5+DVCO8KS6JPOz2Zm56jZ9ydVkdNHKJqbvMrskmMQYEWR
7pF26eq7FHYhJEMwkRLgnPZ+9mZfHYUc9AhrRtVqhFqxUrq6yRjHgo9eD1uMJ4AP
4pmrT2IWqEdmkVNRKdOB3kKtL/iQx7orE0dpoUSx5R8SvshU/kVnJR2iSnWd3+mf
LbCkvcKFVWp8w8EMwgJlDDNvV8IfEfPc667zxEqfcFmOZ09bvFQ6NEFNRS02wmFq
QYhg7qPf+yg1jBG2P00x1hqhrNnc4NGaWJ0NwOFasPIw6lePkN6v7WOLlzESdhs7
BHB8VmS03SREOG3henRjE5lC8iAU0/J4JjKQ//S49ncb/z8eBtBrveT2lZIIFJnW
2n/V3LRNxQZMPTen2QaE+1oPSKvKn2lfHT9ULxcqtdDMrGbcSWiUJBrP9AU6u6KO
PX9HHyrXfRka61xI+d3iCXbyIJRA8mazP+z8fLaH/kTP0LcR3eWrYAzCIR3Wf8E3
0GI69BUc3xLmc1oDRfYW/Ji2Jvu1J76QiBzcoDFkGb/z7DvEyvbBYuIt+jIrQkV5
bfhN2N2IxVRJy7aUgyUPUxNEUBB+/46w72qbZJYmEmtPtyWTFjKPPXUBruqXC8vv
nNO2v7WK079VotMWm2vVNnNWW4bXOGUHdlccTwbXllClnXahw3j8Wog5ifBTwCyu
RfnFKipjcX08xQGLv3WxqEEtSM3ollT5a/CsyF4JQknkNHyKVoFW0Hq7TfAoz+h9
kLcInCY9lbKHO6T5Fs+Kf5B7LM4dhZfAbYB4KRtN2YxosbvCq5zAEAOOK2bquoZV
uCK5j0t2NH2pqq+6DWwdAyKimHeSQBUYguaWMsaYoT4W6ygwXZDyhl6CeSvbtaWp
PqQ8dRYuiYghlgs7PyHEAZqJDrT7Op3Eo0FTXQVgBWo496VOXbtlPpgdc4inpwnA
Zx8IE6Yff2jYjKPh0qkPfFpOi51GQ6M/jLHyY5HEXxh0OBiy/Y8F9u1+A4KP5+7Z
JNoqVSqZHkLJxn/rviGp571mXYUsb6Le9L/n1ZdeGeIHwcpEgtDsRPVVZG/R/FKr
aB/J/3FepXMNqUcW0yoiJ+psb8FiZdADa4s5wvOyZ9fWMQZavpzjuBgIfRDeYtYR
cjFM+0D5m2Me+qX91c+XcXeQA+EcaSE4jwpF5RdlH8pmjtCr5SlxF9ZX2rTPaf0I
kq+pyQIMFScKdYW9oclQSbHDRG1GRSTfBZWuhaZq63zfnVSjzj72CPMCxB2rLF7i
T0dGQqeub48UD76/e+fIUBVjU9rUzma9PXnWOXylr9EwwbGvqcNPgDFTL5qP+gad
Fhe7cW1kH3s5QVO2sq/4wmcsZKg1FK296xXy9a1I59atISPHCyyO+wRZ5XPFkRkB
suxX9KSbi102ebfLr1vurBklMXmt8G0rH5OnOGUW6mn6ci5RA4DiX6AxBxNSU/IM
W/HmKJYGI3ktTEXD+O0vuUWihcAu10tS200fi2dJr72PUjfA05+TO7PPnX66egI8
D0EhyureecBwSqJQJdGIifkArzU00UabJvgK0YO1J2Xcs9sYTEca8nhR5WUl52SP
FeDXxwxI9BYA8zQNyiWeXJ2SMuLf31XpEH922XOLR/E7IvWDZ5khbpPZ5Zk4U/2k
YUn0pKYWfjmZa6X5O0xR91zHkKpymRpDMIhsjNc7zIDE4AnwWdCIh3DbftIa12lD
yzF1LUxFTbUlSHBZuMSYlUYQFUrnef42E4+J4Qq0/sGtBPnNvIYPrjBG0W4OvUz8
PpWgSrV0MDcEgKNl/9QCL1gQJGHMGy2dEyWaz4IF1FqsLzWRjF/1+xuFK8C6sa4u
rFos+51qkcG++rZINCG4OG6cF+BbMkZymB86CUMb8vXCkjZbJEk+cNzgvcww1KiV
+0QyKM7zm7GXUWEqgUtTbJr+6LWkPRqnsv9sMhBGYTzz8NTWcCaDybk2hny4iWio
ydEZTe096PW4gRXpUT5gPycC/O4iUQnay0/B/lTE6ZlP2E1HXbUbQCHxFc3SmMMZ
30KTVD1BJpkgP+ibPJkEnVjuEnuJKY2ve9Il/OOMg2UOQqWnautTtxIgEcdBzKrl
sirpcr5cbXnPTOmAEU6vVKnBMak/7EJRHjY5UPRwCSUSvtJmbSECVnwWRbtHe0R/
vYVU56IBVSALNYKVM1qN3pxqUom19bpqSr1+DufhOs+/WiTnlH4P7x7XReRj4eTK
EIs6ACbm0nbTMFl1+/mbpBMl++8czTx4EfJQlBrDS7L1DYyzWb1EQ+4ZfvYtpuhl
s9tdAkU70y/NTkBjWKjA9c82bhg0yUIYkBzZGhZ6BVFcv9oyhmT4omxEqyHUq5jm
9fXlPY2ISHIJrnjo6TDhX+NhF990NUtZu+USqUoVwqPyn/TtaCbgXgwvow8LDbtQ
Ca2mtp2v6CglZy7d+EbL0oYAawzVsp5FvZSrT29MP8xhwYntBEVyujx6ZRnCRCab
3ipUNOQppP3vQqfITB9B9P4rmDzvdneSLbiwAypvx8a7e2iRjnlhwe8iVF3+OSgY
5IWf3hm55XWE819QWE194VmSzD7WZRWYmD7LH0bOaKG7rKKo5OLyyM8zKI1+24wo
dJQddxDd/3hVsLY95CjeKVYakte0J5T73shZ6PK6jrAcMDRsqCZC9sBrphoNn4u9
KLZpg4mv3SrbZ63908Jijim2G/ix2lbaC7ds9fk6pjRjTG9qVvge8VyR9SMvBYeZ
xA/QCk1eYoWvlkDuCIIDvSEM2tMK9t7vw4NnusCwX/N6T8Wo5zLsBQvZZloDNfvX
0tyrQJEX8eg4X0MDe8LTi2n3mZsoTI9VI4+DK+S3DOHtBmr3EHAZPEc85taywwmC
2+zKzoW85d9zEGwOjzpLbrfb4RyvJpRf+T+LnxGz+2qJxfTlsVOjG879HsKId1UU
YUssYEDBxcP+Rh8WZ3zqSucaojFHQsLdVtWDjiGRerMjE2rOlpJWvjcJHUhnQ89h
F80HEwfSaLauVozQIyAtd+yvLr2yyfBHmN/8VMhIB+xNm4CBYYhEf/FaqBJBYVqb
+DES2aqstWYwulwi/CFd0vDrNMGSrjCdru8nFmQFwSKSIVRqq6Yu+0ymGIea6/uQ
lv20QSIDQkRp+dkSEGFZqKfK1O4RGcC24h/BSthq4q/hCH79zHOSJ49S0zGrP/hD
NzJ7n7jHzoFmBAVy/9olOW8yP1kc28QGiB9Yn+acJj/aBPp3cje03nCAi9aVaYhG
v543WiUmun5Qary1h1aFHX9nOmoU852h4QM7GJM1FmKCOorXZZxpe2WGa1CWDRjZ
Ja1bcgdXgDglLcQoJnWnta1rNu+CnaFLpLaoWmNq5ILMUqr6V7lAbnuMP5A0qGBr
uxFcduS6BXUJBMy5mATLp0execdvHY322q0ekOgn5NLSraccA2KojKguCwPIWEyY
61mI+12GWf+4vpxsIm4o2A21+ITYODzoXhmgjtoH6zT5kDCTe6fnTLGHBe0uYG3w
Kqd4GIXD8NZJXW+C3s8ZLgrebAB+7PAcMR/zfXcmmM6L19hSF6m9ONu2lYudjncy
K4lP0XywciYmz78OtG+4kicTClnbWcQ4xTxIu/q8EsaSSeLyVNxHpB+cGZ1x6mSm
VAMHYFQ82rQdqMo5rPRBzBj924HxRylY8KL+y8TFWEWVPjoKk08/NBAJRGzfi+BJ
Eeqn2vhyDoez762ECtksvwfzcNN/9t2eakPH2B/HnAU2dowS4kg+RKHI5OCX6o7E
2auLrLnfc3zIgBbfUjUbREDk8IyyctFB484sK1lExy3Cak9zuNbGoMSScNSEY/TG
2rHS1+xa3uw7/6+tfEnqwRPZJ77F9hKFsFQ2iNRkHQpKXpCZj2zqPABpKzCtE+qL
hWM2NxoUs7h8Qmd7jKHKjQOTiShIGiCqXgrpmIDnlde+YRBNYyVN0GKBqQ2ymDyV
E6EokYJ9i7ckhimMb/wxhGSpZIRSLzypmMZ8L53PoX3Z+uj3JeGbL/PwjgJemsiL
usv5HNxC1nTh3EIk7dANXpKo1Xr7iSH3GhO7vFg9cLcab1XybfgZcyieDGe4SsJk
SXlNfs0V3OFk49dY2fG/F7HT4aSln5SYRbhYKRFudI4FEYmTrdNx4zp6xwOs9/dC
9wRBKTRxUU4gBKuIeNYye93zqDKvVbi9/+LYphgImu7GwdJNTOlCuEXX0f/zLokb
QOSteqXTsOssiu57x0BZu4hPqKKVrgvbBAIAv8mPdLPxWz4oUh/DpDIQiYmm79T0
jf8UAZP6rGOiyfIPDmU1qyjK1/2ud28ErLkqTaQS409Xc7deFxKtHJ124XJlwjol
EZaiat6/p+XvrnnHSBmLHFWwOg44kMW1lXIeOntrwhi795ICMbn3YNfhFZJsZzWU
l1r2ygnU2izaGcBsaziPr7Y7/pu8umT3nJx3a9zycyGS1Y1up+9Z6kg8w78oNK2R
9UyPsUiLyIbM/6KSeYU5h/7vjbKikYXLOcDvvuxP4xa/P770hdKmeSQRPLf9Ig7d
MZRELYhBf5oBn/6CGXd4ny/6s3iPZWfOgSMrnc1wExV3jTGctkGrwxIY3ZEs2/Pp
RWnA9imuDRq7vHGT+htMoKTjzil1raFeD4q/EnalMnVXJqjKq3uZ1+SpUx1MzP/5
Ih4W9MvDL1n32C6TzJ8Ix73LPXZqiFWIHLcTC9xnkktec9dj792iLzF2WAi2Mt9l
QUMGGCH9XvCCEjImzrvXJngekfTkAoH3rzE/WS1px93FwxF40KPEaDn9rNPf2V2C
6sid1DXNOgiTB1J1G3c66LlX6EqfGj59nJmS5PSB50AdvdcgrFxinLjKrXUhV6b4
0NjUdQxQJRlLNfRSvF+ldo36ZQ5Q4gceZH5keluFmNkmRdzsGxi2dY1YuniqtOLe
ZW5OdI5QYxANfcO+dMUosT28QY07uSTvXr2k2uWO20TDXYjiKl23/j7rv/jqhPqU
CWTkiXC3IpJn6LFtXBpqrsE8QyL9FlGmNDJYRpIQVCikUA/cNPDTb3uTJy/FQd9N
bduPPCZk+vtaw/5MI8+fOM0+Zdy4cur1nn+BUAKuYA4qnCzUenskYnbMrK7M+/V3
2tcPQdwUH7QsgnJF5vvhveZ7YYhSQfpUJV1DNAw6rNplCk3QnUgPCKx+ZMI1yojL
hwzSwvmygd2we7N/q9jtoyiZ5dB14sFz2enbHpUiBmPya0nxAcHrh6OU6wHQllD6
H1V9jIUQul3QqGJmnFgNNKj4p2V3StWLHjx+ww/wOlxZEQl5DAbtjMmm2znBXQ6p
kGwzv8+7KrY69kmASqJ+JgKJncBvPBnJt8wpThBHLFhTqvANv3MR8+skoqJQGxlw
bT0hfraSHz5+pZAAXVzkX/wH3u4033sJci16pNwKmuYbnzcfAL4IDDU8ZxZwNLgw
saOn2MBIFJzEKEbLoEbDfdLsTnQpmWjmBtcSAwevD9SZJ+hyc50+D2Gpl49MTSwz
aoNq38Q82PHxj8PUJkrioWug7GjAvr3BB7UESRnk8Y4L+izfUq9Q+NRHScuT724B
q0J6bz61kZyCUxn72Pe/kq4MwZc5cdH2VFRxlbTpvlfhZzsOKGgOvizw61NEuu5v
MDW/rIzAkxDmVdYtgtX74wDZWRJnlIgtURnXikxCs18nYUW4yXASPcgh3MTEenut
pTZtwMawOEuTjysC6w/e7YsUDUDTqWL6s9mE1fVF1NgT6eTTnmNd2A5ugsG1iWNc
jE1yVAYMXoZlIK3ANC+mXymfYCUxAI+iN9Nul+hmqY1OpTHjSG4cu+OAALnzAdKv
5nDOJsA9klMnc8iXENYF4Biy3NPojCRuSHsVGt3u1Q6KfglYWoJPd2ceucAceCFm
oUicL5329A0/eGIg3dglz8aANUJpy5IUnj6HQz0Hau9O9H1kj1maolK0uuWxK4Ex
H1fNBZzyAYm5HfSmH5usFTjmc4Z5LMr+mLwNbZVeQIfd51NtNVrtWDG/YY2dHuc4
A0aZsuwY5RH6/Xt/VGRAE6fJEBVG38svU9pjZMHM5H5wut8wuQsu5xR7szMZF9Vl
Gv5NS0RAwwMv1zzUtE5ERNi4WwEFml4GRN4DBJr/kkdi8fs1Pf1nwPbkfeQzFJqF
mPuRmwhAEH6wyA2jXcpzZQVQeLiLLyOKsLwiqhoxAzXrzNkurPicFz1K0lHETMSD
+loUEQ4eovaxxhoHOw1xSiPCLeV9shVfNp5j5z7PXEtDl9bkr8M/hnVmvy0QnrLj
njxBYXWcbKEUeck6vfo7Llysd1liHzWWVF1QJxHyjG++E/gSxARR3WHBDZqafzMl
Vz5/nUabE//c9uI4iACzLFGSdMnPqSzo543XwSY1A55qq4b2AzP3bRkT41x2VC33
WZ86SHVPKzYgSZWTpGCTdjr4TdJNncTCDvUALJiQFZZRmcA1ftondKn3JZ54gxUi
31a65SJn9hwEBxYuYZuTP7MRQyDu8Ot72IWT+WY2OuucRc2zzs8qk3xtybW1FxMV
7W7dyaKB3LUM9fsVqrolSzUHXgALyC/Or7/A8hcVSA6P+UHoR6ZveDoLsKIyOfsY
DcmorlaGXarSkV+Zp81JvdiJekCMucsHcTl9a9na0Fw4Ny5eVv1cVkgi7jJ0dJDU
ikOwIRx2+Fci2HJXchYx1zKMLpUPyJODlNCVVW2+2w8stay4nKskQVhuk312cZjc
yjUbpEZNy/d8VyjsiK5Qk48WziMoswlR1EOgnk99upsgVGioC57as88QZ0spQ2L8
H6uRZwwhp06d21jFoIh/OjZrl9tE8LB2fXV1gcC4jSKlObvfp0C4h92vpG1YCpkD
Re0bKkr1jJHT5DQIbrXv4Slu60Dn3Vyvzms8W6P/JLr03oNRIAHVPhE+MarP2Uwm
DzxKNOpJhzeE4Zm3wUzgX343x75UpYhFzR6Qk4lWluZO3O8XjMeHyiKBO4PmnP8T
opn0rJ46qR09eUrcVqLHJzD9MoP+s4rMBqhAmeqynf91LhO/cdUOcrl8RPsZOmsv
LMlqSiS0nS7xn8L3cChJkZro9I0TJPeNyLFw8k9WT3gpA8FIRuIO1ySBjQDvINsD
HZW2lCMl2R+KGaTYjXxBcg9wY7wIs+6J4mNpjSVlcdbu35T91JPa/RhSvGV9Y30b
8MfbWl3PTxQO51z3ENQZNYYIeoh+YsN1jsIoggOaWbDr38IOUdJsuwEQO8/GWjgN
OUWa2bMNNUWT1qUH/pSmGitg3MbZXDzbUe4pfUt69nC/kTqzFottl4AvR2JyWiu9
/zkJd12/H1yMszg1W4AvsehQICAuhUZRz5ButcE2EFuwZYPIQkW8fw6Vrac1wmID
CyY8+LerzvJYT4v8Wivc5WDdtYKDQTLA19557M1DWt2PyopmP4qsl4oO/clQcWeV
y2nqH6u+p9hsTVKWiwZhmhqWYNpEBFqPWhZVedwvRlF18JgbYy75Jlda9AI1yyGy
GQnqAH4AKKqTqRYIKl1GIcgWRnC/CEO9e5leZHXk1QhGTQ5h9i3ZdvWE66fR1ydb
nNu7fZ4DeWwUm1yK9/tPYBdmG1JZax76vXXSJ45bFa4j5qXhaLl1M3tWyY7xQLnB
2ZEY+cehWQwDpbLP0zlLfxuapFH+ECQlg3dZxOcvpsaN0NDCa2XHC7Vnoe1eNfu/
Bo77qU57tDRZhUGD8Yu5Fp8d8E03HTteE9nrYfC0SwXellIzUW49xVjTdFYlChvW
/q4wnifTXEcxirGTivralKz2pdWZ18wZQqyyeRAtLbqIcEQArqvwUWySMqcG6cMl
ER3P8Y/c+dwe8PwO2q71BN91og72lWUtu7E8SHvjl+tmT+aDn/8L1qXLlxNhD5gj
Q1ye2NxgeEIDPoHtf7dEROCIRkw4UH43/l4i1kmViD/YcnJcsiGOf9HTTIe/tGpC
u9OeooKpUikPWy1/jp+TGvN91ZfjSi74tzcWnSnus9ky+vIJST6nqvERC41rYc+W
yat8ed31BtPBRB53zp2WVtmyZwLTl4zQcMuHpIDa2KbwPu4WAn90MYmaxZZEaTf3
XyvNev0WsjuHbAQGuVmiWtha5GoiAr+f/lVIOVV42OaIYkqQRrynCkrPH9iPRQ6l
kDPAvwgdjniI1XhKjrw7WL00xav4f4rGKrAZLF7XqQRi+O12HG7/wrj7luRcZa5X
8ZzGkA9xMLjNMKNhTCrZthz904c6xDDP0ro7MNm0BPR7eTtW1n2f9091wYmNdF4A
kwZLzyafI1QVj1Gevkk7sjbapj5qKqA6QOV8GXkhspJkWwUHayIHJ2/oJ55uWQTX
ZVtLlRu7IfR+NRtPb7Ueh8j2eq9WMbTcI3SUDHL8CXU/P0lB3GFJ5HYutGbsZoOW
67QdJvGsWC9IOUgIZbwfty1iLJJvZg7X2KOLcIlvLqaNjequdb2o0CEeepAq1DTj
QlnuZkzR2wyOLdGe0EhW3Kv78paolGoYurjyj40AxTw4doDEs7ADeC7c9ZbO+4Aa
ZZ5XFHpmeBAH62Sev8h4wkG4FvdhYAXV+Y9qygyiWrMUXn64tiKAYzqpYTKNXQ5W
jVUg7r2LD1Xw2LkwS7MMADizV4431a3nV641/Mk/ksoV1WkOtcMo1Wfd6wTUAPQt
G7e9n6WLTU6ZnX+zma3FTW94ucTT73F6rTmtY72d+J4ij6xr57SiPb6MMosF219/
nIMa1gbhpqftYEjCHeMCLF+GX7DEcysMjVVLm1FvzQWc02tzNJ/Mq1OkXj3suxGY
Xal/k/2TpdylaeMFj8AxwwGbIxvljvI9oBgtPQIaW9dUTKXHohg/blunGbVnmM1J
ZBTdR+dwpE3urVf5aXExseMjNzlOQSMYVaY5a8MbhqStJ3ttvjwrBJDVBofOSEz7
1ndMOuFDky/6Z31GlRtFmoD38DSr17EpItc4ZThvIxvfylLuyH6EQzbnX1PRGebB
C4P+5C3XoDYFmvMNZT4SfJFOH9j4CSDjiXCmlVyJf28O5NQKAqRK9a0T6dG0ozf4
AG6os6z0JU+EF2woBofoSidqWeuZPKDpjk1Qqid9HqPlIp/ksf+FqoSKK1VJBJC1
yZfUosCOqVGSkwZXLCDjxZcdmDnHuk/Yd2uS3LoKHUAq9+MK/kE79jPAd6MOY0dK
1Tz2yf1bF6DyNhK4xZ9F4u5bEw+G+wmvUte3y0kvP2p7L1wZOzQYuqNltSMXZaDY
PfX8LQihuWQXaDZ06q2h4EFl0Mk2G9vTO0tTqimnakQzOs17I6KF/QZkkJ1lAmEY
sDVW1H6eCoXc3nqQPiXFmcX4AhFPsF4R51KJdR85ppqXJo/vZJK+zIxKgWil8fPP
X+rJbGRSYNx+q4r4m460crSHoVf4P/12hffGIENn4wBttaM90EDoT5k7dXeb5lmc
0yNbJ/u6PB4e3acMQqGhTa3dAP4tJuUDrZCc/H8WWecS0GpWaJYlP+0pGCWXgizf
nPsl9mq5745Ye61+14QBMrZO1+Gt4VL5hL641WHJYVGn3VNTjTJ6sLJb+i15vHCy
odpiMvSCTjWzDoOotwxOHFuQzRGYx8RQARTDxx/teWchfnE5pOUkq5kn4vs74wsh
lhHcwUwzZXALHVkGN6yZqspQiWFxzV08VfaCp6JXFe9yhR6d+7W10QKUkYUTCGZR
oSqdCuzbAzgHNyeUn87G+EP947Y3tE1WnyLl1EppzNBaxHJOdy8S4DnbJ69Wj9Mn
JRNULmqRXZt3hMEjigaHemVQsjTEMyAyJ3ZQBlyRS0WMfEYTt73GOZiIZDOcgi0P
lTUv1ZWf88UMYiIZjNXj+DMcofDnp6OMeidziHPy03GrBQvYnGZvWD6hDEPkGyeZ
5L5Wf6Xb5z/Je2jrP/MHqNPYjETKSvC4vhenvzrUz2yZhvfMz8R8osKrPNRK2pQm
swTwj+5hEaGMWeO3l+mjZTHSuaWtsrx7QsM64BOZWXudqBSH6cat8mwUm+4IfS0a
IUOMAZ+ZYGuKBS+gtYBAVhiu1aJO9nM8OVPYaeB+7hhKTkcO+YKOuO1f8mqjfT34
oo1zVS1hNeMR0v7zIIavMun4y0j0F4NabyY0s0I9CaIjQQRpDILegEiGZu9oJM74
wjS2OYKG6DGSdIlEoHId0+xPxjHYnrHFsFeF5UcAN7mx7EsB1jSGRvAuCH7GAXR7
9MeailUzIXC9JhjTGdRgKtJDOTy9yOGaGkMDrV/U7nBZYRCsgDZd3nk+S5BFhwos
XqZxOOKl/WIuJRSEsDYPFtZr1DLgmUG+qjYcBC37F0MNK/M4K8dIwBNmSG96cbDW
5sJanJdN1mjRHLoyee+jdYLTzX26usf4oPN2LqQvQQ5gKrJuIK1GO5RLveKrqetm
irUuimHREYt7MS7NGu8VJtzDKGgzkmwluUo/fTBV5mEGH2kzK1PhA8u5HxNfWdYZ
2avmungoZnnRH3AwrW0v0EC5ZpC1v3xuNdVWx62ksgjzxyNjACkaIqPj6xYXqTl7
6gkpqNmQdrK2t2wnq0dGRtsIC+aRDwCCcFTiguD8Z8J2V3WmvcHR7qM0MG33IZaW
TGCHNM7WLx9mU918pRwADWYJSHHc8kjRL/u/etWRPTFW75cKvmoC+Mbxjg6tF/rM
+m1sV6iSsRANogLYgf9N30hqth5E7LU1H5mJlNSeT4MHzWkASB8s0SmLMmYi37W6
oZhrXN82Xj0A1Z8NOojZvgdhalGssmRMHUWJJD0mpbtZjSwKkNkIUYvxeqoD6Aue
IdU/ZO/I7VeKs/ZeP7saiDwoygxi1qt6N7xxGYIZwpjq6JMc3ajeJujRUNCE6oph
L10QbFAVQ1GPADMgv8ye3HHsGE2K+77x+GU/2NiSo62N84pOVm+qsNC/vB61pi8n
/xBFIao5R+FkGKcDSAQn79s+MLuZU7fjsNj/gXfdNWWQVLNdaOZq2xh2oMtGb4re
gGABhpbd/Q7CN6rm/KKj+24MiLRuV8lfJQX5GscArk1Qj1K+a7tGyevr5zKkKkKK
cyOgv1OkldTnks32cbW/7U6zyugZC2FUGtvKBG4hPRUuwlWe9fZJacan5A96nKNH
ZJF7x7vzRl8NPc/6wmO9WjPHT+/IVz51JHtNvBoZON5oCXmQj1audQxXEDI5Hq8u
0jeFsh1Om0+kKACoB76GNANTTGcBDXunBW/zWp/AQBQHI71J7OBsZM++eaqgS7Os
fDcPLRNFTOzy/9EkjoWX8954IHkOTVpJx+0g8AUA6eiUCNEGYObivVuHKL/H8YLr
/NA/2h+694wFUysueEgBbn8JIj5xxgqwzsKPqDAsNFGS3N8HrxQrikPTHXqeVVRy
EFzzQLDxQyCgB7dR18MzSX8HbWIb1OY/BZ8J6cpDvyYZpGBElUUneV8dj7PNPYg2
5LmOL9POChsfdk6vUtGa14aIfy4Un6Z9DYD0pmc8eYgeDJPnkx8o8noeC2XCUZQD
VNqGgueM4x9rltruGmEwGlDWVTNmPuPj8l7agO7I1ecVHi4ih6UFAdopUfLKBnLq
zoYQqNa/PTQx1KSJwHhFPoBn0KyZznB+8bS/oY4dKQeLSDbQQ9pjdp28Q4HQcZ4q
xutwegwa2ETFfgpIOhoROujlTMfV6no2yfJ2c8OYDo4x9+/z0WMXH07Vn7+1ZZYB
TGbP/D6EMcwb6aNewatpxGGt/XHkvrIxZZqm7toP3+wPNS7v7W/SWImM/xj10ZbL
xtuxsrsrTTHfHhRSCdD98dhm1XaeOavhbj7YRUwjsYD0FnuEIRZvGrMKAaB4xG+2
ralaaouEh2AckgepvFMmitP4cobaUktnTUjf39nKsoNmIRxYnBfkqO/0Qy7pSc+o
Q0ykznCv6qBZB9r0nkZSUprlaAKY4jvjjNFzY33H9dN5vI1ZFvr3jDROW4Mo5bHa
rmIcS7j1KTNBEvfveJJln7WuBrEPLihuR/XhOGbyvHCblxPIgTBgp5xqUHGCwkou
RC0kobOGFvy70iHRAvtAQLO7njljjtbvznqPFigWCoXkX7zp1yi8KmBQth6mgGvZ
WNoHy3ZchAWMlM205EW/3ip7ycHJk2ui8OSUSmAbio03PGn9XBt0wUKu/JsGIn0O
ndVewJMSOqe/XV9dAWRomWprDbTF4NruTuz0mIgINE2nIbFJCrDxiPClo41a2fQk
n3LhxO8BR8QTPqrkD+oi9Me2NREFy8o6kRp8OVpQwDLmT4d6xFTdtpo5cGA+o6pA
N5UFUwpMnCcfffBzlwjjbBG7deG4pKpqfyAg5gz+1b9xkY/LzNd4+5R6OYdeyLZd
CygJaADfiiNdatD8Y59JDspCJ0OolXW8CvVi7pN6VG++lgAVJzJDHM5DFXHW7wiH
PyzeW6GEK9Q0qrwWlIWiH36q/LiBWA102O71rL4VOPWTZZkqI/Zr78QNFwX6Herp
EbfGpr3hsY62+oy6HXCPifIFvyoxdfq8xdwRI4e/t+FpNeZ2tcrs6X+x5zwNKyF0
HZcTf5nLqWN75pecWF+DR2RZ9+Dp6b/0kGpNvCC1sl3bqSfKmHYdRUQo/4vlnAhT
uAlSvAmh1KhTgOMvG4S5kFbLYDd+mIXrzPB6a0a4XDoWeRBmmV7KvXAvnjbaM2p9
/eZURwp1QVyjRxLQWhNx4cuL1zDgCrNS/6okPXuAx1CG3uQH7oll5aetm3bHD19l
EXu40OHLMLiiR0LCv/fm8TMMYwJe9QpoOuKAevCAM0YmpfEy4aeT4F0jNnT8BUEe
vDSq97fdXNNYdXOAf7kqEZl+mZW09USlxJAw9VFoDNJ5qZy0I1G09b6MIeUS4BAu
YKZld6DLTbTVVYqTc6YwYmwb1lwzGHqt873JODobasQeBTnMe97D1slsjeTzUz72
o/P7dlbTOIyRSzyy5LDvIL073+lQm6AOHf6DQgFYGfe/WbLQ9kB0EXcGt+vvqKnR
V0VlSJxv55W7bUXBWZEJirrdIhVek4UnMExbPCCrr0r9eZ9PGSub0d84muhabdCE
/dlfF4deygymmno22cDWOv5B9b9daDudloGDUJ8/iwG9gJONevqBuLsN/UxHTDNU
9iX1lyH0keA6fEVpWiew9d4FwpJHYYiJrCtRDOXwveTlJWnrMWdyiRi4b//GS2ZN
W3KbmFJUGqL3DWJFvHiXTPfVfBmjk3aeo6aPOqUlPgbiyXYzTNlInJlz0nfwm0Et
DSBA95kyhY5YKzIw0t2DZVT0vmLLeSVfYUF1fKSo16oDD5fk/i22GBnkDRl60im9
XwYnJ0T3hkjAMeU3c6iEDPE4PU/ahW6zq8tCzPV/DbU9lk+wKMjfburhCrax55wa
B/+L3IBVwAOpRLR62nLYCd4QodtKjlvHUdoiqCElgZsI7kcBOCOGpUhz8YrC1IAA
E5ZOq4dv9Z04IL7SLqOSVhRSrWE2wI83YuU2BP6Ec0BBSYW3NcFMutjSkwY9yVdL
wXT5327PsNysjTX8yd9DRRiBFLI2xqmsO1fUn3qcKG6WE9bzb/G/4jZexrmtSBSS
SKnieNCdspPJLt5XG09v//byWaVnzb+o+Oc2eBFk234XPrm7gA6UAWFIGXdfYtcd
PU5suVn67xG6yk6lMsqyAqkAOB2NvRf1wqSAb5ntrcuAxLrGWZzxQvkrnD/iLi0Q
f5aFsOSAI3h3aETbquHXoHFZEK7k0lKkMWE1XNjmRgXrvd1zLojFI5YJ8Djrs4Wg
idiy6peaHMHotxPOhyleJtFx1DmT4tcFU4e9tDk8AlsvV6JKf0OymKojzfNs5xFY
IMXUevggffB7wcw60nuCIXR7dV3LWuGad6c6kU79wO1XSqGmVk4XfWnLS1fSD0fw
gtbNB7J8wDT5qAusMwBsSE59WzLZv5ECUi2KOgKs1HCjSoBP/s7APXTHapQdq8d6
xA0aFZ9nxosC+H9CynEIh6nqQUn2R69nhm2BIcyekk58oZaVPB3kV/3KTiS1W8pF
Fj8nzH/0KbuwmBTifKBjIwX434HR77zruaVZ9CilATBcuINcqoQMO7DO5gokZW0Q
IRZnDpESL1bGFtNa3RG9DFvBKsd2b+gPZ3Oipr8Ykm3CU5eFmF5m9zKILmVe6h4k
lnM/aiNnJtHsxSCiOweTuSKs6DaUSWr8sQmrjCkLnE2DKBvstksNHMA+XD/cFmH3
+3tkfPkw0GK+v6Sza1SyACcu/NOw0/INl7wAekG4sYObmn+CpO1JkfE3seymftFP
dyLs8MzkWJa4uRWxKmLtc+GFPOTpo3zFgQCJE17ti+3tMmU8K9/dv71xi4Sw8BCX
McxkkGhHeKX++MSURqwHjyDkYwBSh0tUMKdDqcDSThCoZKRZlBkBHIEpvDEr0uck
PQ/Rg3Ll4U/PPQ1pFe5IVCm3ypKmDyylOYHTMzFZpnROQTPBv0hqw0ltrzR6SDa6
9tAoE5zQLS0R7ScXKE041mHlcZ4nJzV5wXFSUKhEitZb77HOUCDHDdvtiSDKl333
os4E0CF5+GFkHSbfoP390oo9V2iscVN81+OxlkzvirZKUhaIps5rrusLifpQYvgN
QnZWZ9BbXZW6DkK6O4b6jPbA1ReYIXCDf9nZqHDFAff9pO1o0iki3iAh2Rfj/JlQ
FC/IVE+LMwtlFiZPMzvszscUcLAb2ScDuhEmku6kxGL/lSdAqhm4iRuSa+g9jrGO
WK+Z8YsSWScVUJ1RE4GwRFnl7X8UeRAquhr9o7u6i0/vAbD1B/5m8c6xy8jVOkp8
NsdyWVkJ5I3RiaSACd7qNYb0YwSqJBsADU9vvNLJu1Ax/FDi1shHJ6CaKBtPQ/Fc
JsJZZKKoY31byCBGOJSJp+s4DFezqroMJoF4oY9lRJTOQpQOXYhiqWjL42Rmc4NH
fNgDD77/ZJwvl4Ua0iDqRkEg4jFIPCE7BDCmKj3oJD3tOWW3zFhooU1cycm1237e
pj7Q/fnFL+UvWJPgV0QY9+vYBNrIfJckY8oNojPqu8hra07J6fHb0Ai6HjkD8hiY
TwQEuJ78eLP2rR5cHCVipQqaGO16ac1+rpE8SbbDJrXOAxE4iNtaXO/NWtUpvwDy
REJPJ1YOqG+YsQ51AoQrxLNFp6pRinCPppF7opPOTEAAGaPW+QbY2pclla0IG6Yx
D2i3DTh5GOZ21HQc7keE6oaaGhggeiegFFd1TpGA2pcT3DCmpFexZmLsk3AM+Irz
DAgWaJ9Fhu+AtW8mgwrjbpHSDasOxnula7A0aq/EHk4Mw0YuBUta5qIot1GNZ/+W
EWjqPATlVblINotIoEb3Gm+LS+Lv012FpEbNqhTDjURRCHxJ5k3uBS2Tzds4ewEr
FGoE/rNrfqfzoTJgHcShofwY/OgPAeuJEwW1JWxT8X0e5Ns5eWZembmm2cb9z4S/
y/iPU97rsYqpz39w3J8AMvLr+5HB6u2KFxnm78wzFvCU9yS0h34CICakdFDuzUmr
F9yBelgZNeu4kf7mmnldXuQA3LFXV3U30xY0FcNdFoKseEFLGtClpJDf/2ITIiJ2
SiWf+3MBwzyRjuCMEJWXvzxCe2Ryj1QhEY08Mq7M+lEqFfr+5ynusc+sHiZuM893
cBRdih4q0oP7svRVOhef8WbdtxT1aoiSeHDkRdb9doiND4I4HtWB4rwzoQle2HUr
oCye6m00toypvaQfgBGT7RPs9fUFNQxPKqzdRqWsYH7bLj1kd6Tt6rIqcBNleCw8
G0AEy+JnIjx7StdmeCVT6EjoUT9sIahYBsU8uUMsRGkRTTcI766eGub3Ue5AphjV
vuuDYJsEG3aZWZl0HZD03P+roGORzv6chrgbn/0ZkPjvxc53d8O4JWypxV+l0S3w
8zzQBtM+J7rdBzc7WR/+EsPUc3QUeXiMigWeMMhNm0V0AEem+Wiu8/Wj8FAhYS1f
/Q75wcdbteg9UmmHC+/9tPaMAVOA1GIfDcbSPLxFlKLpog48AZ3Q6FHb3y+JzegT
ZzRSlJwj+GeX95iSESTmuLI7Xp2+4rW0vxpZLX4AyUW7f16s+XzpOpUMPQSJoOdJ
vlAxfDgt3+ccx/MqPSm6JmlkGrpb/p/z29kO01qMIFqWhjRPB1r1GsY31dyArvQN
sT6Kf8So2ORXCrTOljBWYpiIl2ct3ucAUMYjJ69m7Dgyp7wfl4rbO4emSNPhtxE9
R2tzngnWl7SUm/KpJiRYE2SpvoozvGDF1t6VYX8+F5o7g8AuEGTApgjJMGgoMqWX
+Hq2QD4C/c5jnsGkzpgNqX6dBwIZ+l+JiYfbz8vIG9wWyjzs29htfqw5SINd/Qba
1msK9ewBnfB3xWWFB4aDvOMiGdXHp/EI0SOTBuL5/vP9VsxeEhH88W3esNlyQaBr
TdcdFTZlmvJVAd0HRJOEo7BH6EbiYfqUxKvugCvsyfb393omltkaCfoV92d9pERp
7WGq4N0rtguWhhd+xYcXQPMJe+oGc45gqtWkRN4keX8JrsaDwDZxUToRnbDkaVf1
XQSLw9domsExh9+wOL+9cOSKaBmlvSSX5tvFth4AyaIIDYv5lbH0Bm/f6yuXqae0
3LG+L0A2geiy6S/HVO40EwaCf/6qav2OXaDPyckUydZQf+LIB44WzsG/mhW4rRez
j63lP5cM87GXHhOW37M6ApvhxIDtPLdtJx6SeoDs3ln9Mc3SmqFcH35zt91NWOzH
aYj2dhK2SqmLXwC1c7MoUIaXA4UEkPlzBGQ0ioKE6h3MFA8gayyv38iiQ/DQ+Mmp
oSTHr3zOblRP3BD9n46NBpdf/jOj+9GiL/jVIejg++4m65uk+n5wSMnjZd2jxMbu
wE238P6uw8fIEi8nxOC1YRiaNuFOBr0cwgH+uiFq39g+V2VBo+QRvE13gPoOTxS9
BE85/kxWDmTU0k07jZneZt0FvIzbqU3pN7m+6cgByn7MKI2V5tYbcrwLZHRnsxiV
YOM39vS2bBiiiXFdWn2aK1Hmmw3RmMTvJaG95M/X4RUm/rpcWwwwNk/K4Z4mC6LE
h7kEHq5EZThuvhCPxIcgq2AA7tOCDiqbrfSaVPi4Tn13x32P5a8gOQaTAax/0oHm
FGgunyrkHurPpXBViZCRzlWOZ3GJxLO9SIRbEV+jQinWTahtvlJHcVQKuGXeJc/b
FeUtuiAEOT1zfujCF87Kh4JaIYUX8B571LITtpXohPhiqwYncy9S1XL5Zem6TRZU
K9vqoyKx0YN0lM9+Nw6tf2o/27d+dq3fbDGrrSB5UnclhfKepdIGo0y+oMtxQe1b
0aC30GFPGuZzNmT5ST9h7D+f2D/8uchVJynRehTSqM0uwpTwEK0bd+nsCEBn/mNH
BMrl9qrOUbk7+Ewy+0OQ6MirACNUtZThHY+KD1OZPHRYbzR/Cen9yQs76d4HNOX6
SO4avgI9UDPN3sN//Ev5HrSmahDL20Ol8itDVpL4r8aGTD5Q3O/EtfkQvY2tGJj6
JpUfTEdo+QQkdyz2OOzv/1kl6EIOO2vSE9E4Cf7x5naQRQSJF3YcLoRB0Ymz5wbW
fCQE6K6wQwFYySdfulRF6t82G/S/d3NPjoTHNge5KL8DVqWfGkkAbmy/tpKXFEVv
21bpQCksdIfumAffQBo+4BVNNZfX3CmJNWtQCPq+mUZGZbZLnv35fjxkOQsxXv4v
R71j6QUwjHKhmvbGZVWjGH8sqV9atlLYI9RuHnKY77cT614cDWPvuIMb8HL5ISVv
szZOttcw2Y8Xt6O5E/UkEufH+LLWEocYWGQS7gJ2du3W1BMYy9sTkVHLjgVca3jC
i/r319KmP1mW7FMtEFGp4fTdCoUddTwPQkF948Oy3oJ2AXfaSrbCAwQR8/g/yo1s
9jwbPuWBbCmv9eiovuC0EYdf8S/RASvFIEbLYblWqKS7Ug/4123S/iDxEBpgFP4j
gN5CaiefHea75PphhVipukEUd/CPzNKFOifKM10T+aaheaRywIhb4YngsujcvMjy
8pRsiILXPKxkGqPRGh4euaFdHj7d4oaXx9hbDLQrtBjxmhWAaQ2VJC9gg1z3uUNF
kX0jhh4EHm/vJvL2T9r2TRz1rVxBLk7WI7CxcMCSi1dUL/s2Hc37O99kOkn4C8X6
FTy9vFNvriI4y1wTUb2FOi2FQaz2TJbijlVk1psUJAt6VvJjAqovfEIEz38Tn5e3
Ci1ZC3sQB4LioKFa66W3WDFkFcwgUuJLV4YOC5G3/gvNXfw6W2P9jWFS7AJcWa87
5aLugTW3RSJyBpkBW6vs88xBiVWuD7tuMb023vkrqgM3dednFLHbY2K5JNUHXDDC
gchfOrPQzPdiSGQIMtIEZNZ5964+DisgROd1o6yPFiUfjitdUuZfQ1+kyG7Ifzwv
6l8mwwBKA0XN78XAA7YgVZjXvVyPCY9dlXfFS6awSivl8LOOz80tK+i0suaSrxuA
e0sxknwZmiFy4+2cPEwTwddX7m71OGoAPmPWAzHj84L3U5DKa2mRFE5v+WrXRiCw
17XUJa9q7aJ4gvUDiQIBJsB/8MwbuUMhNoQZz8a/iVKsBaZ+DAPfy+3mq9NoYluR
QHJdrc2U/Wjkz1I0SEhfz+ttvN1JCbQhhg8nDvYHMLUE8TTdImV01jF8CvObgWkn
pRK66BTwqtuaMTsPWamxspYAvknWq/Is+8fky/03SlU6XFx8/nOoyO/q+h1Punai
7AttrP2MEOolf97/r/NhClLBLWufpRocznpocsOU/uUkEkTGwFjCuw3pYNytFRbm
UsTPn1Pp93NDuvB6lgcpA6DK4FkAruuFl97rgR2q+BivlucSWesX+iIzoAP6MjT0
yCvej9PzQIjU+kWkJRr8Wo0OxurK4NiFzqzaSY6QblprjV7SEeSYfTjWnjgYbpTT
g9DYdD9aTvwPug3l+mjFZMNUsMxT82tCMGIwIVHYZGKCP0wZ4GF4VY80s52xFW1X
R5ZpfdlnJ8aSXmeKloVTMQOZXIdcdegKZTuikFDqG7XMoLkaIUmrUBqTOlI09M73
kPAUYyWkS5HfDlAH4kO9VZbxbuJvbEqtMEaQ3H9FWMYQIozvZPg1FCCP4g2Pak+f
8PIyIiSsKyM2aq+0Dxt45ywL2wcR6NreTtamiYeoWHKSViinKPQrLXKTR+HAik3m
40KCq4ZmjDFERD8WB6mrZgHTW4EEf4rlH9vHL3d89XYzQZK7CnDs0T+nno+7MKJX
AKoBAQs5veppjeO3JureMr8fVWAwB6cjdbkOGhbun/0qTeBOCWTawwnB8mGI9+1Z
MIpWjh7rKz7/upMaHRIKJy5LdGD3UNR+nr0W/4RSYCgJWnutbJVcu0mCqSpQ+508
sTqAZ7tb6y5Gi6rSBoHZ9eJ9gpbs1GNHvfhOccN5u25dxL+6whsvDayMM6OSyjRw
fup0rGlsL/7YlMCa76a6ju2OPepY6mG6JhUO7fZIYvXRLWw8HX0aFeqW++nrL68A
N+dlRliGiwNLa8U8uFNbe4F+Y8TqkGS9dz7RdcMUrIx2UzK4J5UVOkVzO1rFd5MB
FLbmRHXrSNDLuWThbO6YyjaZnViOzM5FxVS9Ax/6od6cjJteDAg2BjuVAMJdPjsW
lYnFtj4JhpMWS/qZwBOCAlG7PQLUeWkf70yYrfP7Ua9pZK0RL5SuoicHTMrVRXGU
iCLRbvxbLCpESyF5xB74vZyev22pbTLDKmv9x6YAlKwe4TknYbDoAC55EwLpTbYl
1rYuJ04avnmM9/Bn+s0bJP7fYhyyOq5+NonBLf5ZbgstPUG6NfJLqjb0fTJDysJn
aX41US7CvVqAtyW52FaZSlWQhBtMLH45JWeolyJ0kSYkAWCcXlcDnfG3rzEZDaRD
3JdZ163kXOxs1v9fPsIGA0NyCK9fSST08RqYmFABNDUiTrwj4YXXerErl4CKaMjs
gqL/BR6/iVrcqnPOSODo6u6aPrXvcyYD7LORwlO4OBMRe/PWMTbKkZhYonJw9Ty+
fn1owBP9WitSRRlVZCNDtKKyHWrTSjibnt96xJjMyaAo2C8PgpssPwjqFU1ouQ1x
7sa1wXG8s/4a0SAtyyeQ+pR+N/GA5AiXeCAii6jLmnmgCx6HulxfmmagyA7+k6VQ
2CPtkVlYTv8Uhsx9H4gnKPLqLrYEfap/8Aut+5S8PbLlmTmJBxV6ssrusGBr+ZZP
+4qv9wLFOXWB9GNmfCEgwPJzi2RH7SfYi3/db1OSdiTDWY2beNobyPvRkGZGRJtf
ErHTdeJQ7LJ2FcJVjqZyapm9KhGQCIPpmZHw8q4OnKbvhDRbQWm1yZaMeFrOZd5l
lcbaLtKJkwOkdABDt5+u5I+ZkPSIP0MrcaXZs8Rb8nuV4CorjlBZIPLybo+OgYdx
oGH0Q8rFlXi1S6Gyro6gpGTnKHcVMInQCan0tdAUUCz9jkJAhBhl2VnXpoLjFHkS
uBkpeafUdFPCxdTAqsH28hQ1KT00DvKXIpnFBCtUZIEXhs4B0iXK1HwUgP/FwcTD
gqq7+hUPaAB0r2kX++bH8a37ZAAPw/1nXzh+Yls3lub+nllr9DVHkF1YJdPorvR2
m2cUrY0H3oRwaYDBLfBj4JS7UciUAiYwkVg2cuSAtX1fmTjIaPpKNujFQ3Mq0fUi
w7RfJaPh0QjcxPVmiBFVIUXrPuxhu1eqZjvKPZKBArWRoeSBkP61DQmLslFe3jhN
yKPkaj0ICR+ZBR1u29THchsgZa2pNuDggJaoQYjsFEfiQk2UvT4exJFnZrYLmvXR
UD8UhBY42Z79DZe+kQECBEqueSLwAHFsYDrVpmzgqSfjQvdOkxzqSv6Djjh32Cxa
mXiCY+NQkxfT1fTuuFSwFQI6M0EfmNqwoQ71w7yC1OhPnXJEjdg/gEsNhCzbCb/W
XPEDGTIj67xHk1FaIa9/KMsint5TtCXXmLwWhlcWVwNjxXCnBN3dzqu+Wb9vW+yk
M7ODdce5vZCVW/gNkuwWw2cJYebTjWlHyT0Xhg2WzIdo5M9V4m/yGYyFyTu6eulE
yZ/g7utF//35jzt82zz7kDUkMsoCKNJneLhfXkAJz7bPUXPqYCzL0SdJI4R1eoEM
g4S3p8dy/rAbs2S6c2qkXQTMTjRuq/wwJx4kXOKU3PSNBs+f5lgr6Yu+cB9Izfvk
3NeR4RLYzggrEbRNgSr6HBR9YwgS4Tw5pC3SxGU62jVYVYQI6jTcNFJygBpGt9A8
VmpQC2ZtpczfHtDh9fDPZ5H8uQJm+yCLUdhNbs6ioDdmGNcg4sQFuagLoBmdTODf
fxQuRktiv08kECta+nJfyFRjSUOTdeU3pfmw+dfO8vQ3MGzrwzbDeeNdrecCajBj
3hm+XRlwDBYqYgWRc1V0dNwcTwdX2b1QO6NmauzPgUcJQHNkZDWDnJ+G1gVGYxNu
h9WqfqyC83y3GmYVPA5Go+kNuREWK2wTiFi11BKT6cb53D9kZ/QNsr5IeR6FsQbY
iZDfxKMqHI7GUdR4QYfVo7Yn60Jp5sS7wnuDHmAjMn1c5KeqO+/CZ+c/mm6OWMls
7Wra6ds0Wh/wRKPFfv+I1pbeaZ2ldjVGtFP6LWvB3PJTrP4m9ocfJ0Zc9EdzRle0
koXLr/ttSvPzj+sDwgx6xVCKah2zUWxOmYCO3OMwr2hRrv1ApsEzzzviz9U/r7Bd
0NDCc5oa48tU1ST34lwZP9dKcRje15X+KRc2VcvYoIfBXLeKHiIl9b8q0hhIit+A
R1LaKCdkn/0Zsn1Bt0QGEJCpFmNcd908NQOzhXrC522SzA4lH+mcV/S3opuANJTI
mghQZa9zhF3r2YbrIBbJqwj2sXzGTpX9hldjXGbONy2FAOdfp8laGSdnHVu3ho8z
VB2FvCieEDeOebQ8NhSDdoqSfbZfE2xs9gaC8dXgreyu6mPTF2GbyVKhFCR77BVx
00v9ZOjisU4ULb/CujpaHCPj6kQLW1jDsIXMAZmXu6XxVdlhLV8uSq89zx1u7U6W
OYxtvu0P4vV6lB2L0fL2qlvB1oMRX0EhqdhhKNEWXL68uqmIBhRL3edc54EPdh9w
6kD3NirlVL2qRXO9EjwzaZePrbTQWDRWg9snjzN03Ee4trabn0e40uWxl8xJVJ/P
nuHBWCUWxZpchiHxRFYuwOn3E0pMn2U/Nup9J6CPkE4Bigzn0hw4L0N7ymo5AhJz
bIH/oVhW/JWdWI5T2F9wSd/ZooFfoIdJcR3j0Yr8KMfHOokOnN+URYLmJmraZAtF
XwhMn3JHMy4HAfe+sCA80bH76U9pW7P74skJ90vWjI8HH1AqgQ3hPU3dkrYKf0cJ
gLwX4rNdTZcRHUbT8ctOXisrigOTqKnOvkCeMks4rmr0KEBrXCJ63G7VAsdKZFd1
e0jNHCmGr4E2P4heE+f2ljL8bBvVn+FMECMtm0brq30F3E4w2iUts/U2ASka502z
HnLhuZXXAdBvk6CWDmfu6UZr+Ih3wFc9Kefc4bwLEqzP4udu+hyssTqG+C7mH2AA
e8AHuSCzi2vQ5VoGzb1TPvOnobFxRW1uhjBttxWpsEda0WEOen85+ogToPqON088
vllOzxmmBRxJThM2ZQgg2ZfojiLYc2ZDJ5qzqD1AcpSJHIpjkbtFQ9YUsACMOujK
Tg834X829UxLAuZNB7piWxQxvqz95NkwgeA/smHQ17UqZA4P6cfgJ/9UlmCoAnVe
cBB8DzHo/mApVa0/tnbV+bk/QztVtgH3nV8rGBaMwddXOdztDbdjLOoNB9SNrlXc
lIHhxnwZrVMZOrARYtZBPtzNMd11goDGm8xbCZpAw+3i4aKcqJ/7oCoYjJiUCGA7
2DTq4V90fjND8TFZ3R5ORJ2YS9p1/8mrneI5gBkG/2GKDOWAgzuXJx2wA43Nqrwj
hMbzuEliLAxwtr7uaNfd5xr7Twxc88R+2ZA30OAu/3kwAiC3JbT/qI0pMcyQj/Ba
WJRyTuvA2WK9cZCkisbc5sMRaDfYniwsexJDAiQPJXNx1W1PyVm/0GEdyjBcNK84
vHYeVDi3G+u2E5q3a07smgZX/NMr5NC9kKVtaOzlxY+7Ag6x3bnbpRjAZN4/5+RD
dXkSzfTHV4Jehk2fvZgm81RDMrLZQ9FuYUbRrEEFLj2CdmDkrsQAFDsTac07HCwG
eDukUful4nYOqgSsUXYmL8QkHryI8zkxGgw/D4Oz0NqyfL6Y7GEreSWN7QBvhdDj
apbTWg5ofePVljDuhD51MueL9N6lmVt9O298SbW86wXMsFDuwmAaaTMxeQeEbrY0
JvFKQPuGip/tPBxwI3lKXeEESInV9PopeGKC6HpgpBgeA5wAMPGOew0tQCIpbPOm
drKjPinOKP7IDC3ki0ie2NwCaXFeveF7+OUx2hN9xft3P4+3VemLriTwFNSwFSxZ
OzkLHIEVefn1O3bUGQDWAgy94DFH34uXbmdme8yKsXAvrLfecL2OTl97XrFVa6/7
XxjoaW7JPT/3cY5rxk+6CeNghKnPcGBwPGOU8rkFOF0OsZ/n3ekAQ+W3pYu+kWx/
hrMAZkhrMeqmGPoQRr8yUcD9ZovaS4kF1JMoo2y3M8+P45gSIVtX582O0RBZ1xIE
fvstBK/ZhUU56Z0w8wZ8KLYiqTmRWAWVcuXk1Uj1nWvOvfTVNZ9tK7P/TVPLQgGD
9uQ6fwVn15YO0+98ZsNC9P6/2p5YF1j/zLcMh2/mAB+E7U/1WdQyJJbYM1B8lZxF
r/PijaTlT5JpvwK7R2iEMYS0WL4s+Pxx/2dfeLQRcg/aIiv4ND1EGDjr5QKuId3P
04QHw60aDCZYWMyBksguAjErjh8X9d9MvvKqd73/3B7Dd1oFY4/evTmYo6c2FKmG
UGlylZkSgQWNCsw8NiuqnDD53UdjlR5quYd9WCnLljDvSCmy6f33NbWDe1DjQekV
3J8wF38+AUXYM524whyla9fvRZTe8VhqWFdZMhsqWtFnN7GkuYe/elfPoKahFy+C
rTtiFZnbXEV8/TPtvIFANmdtpXyh3/SXTf+euDP/s+DEkrSB7KuGiRbw5c+jPs6K
F6cChs99a8RvkWiEaUywvRNnnfRvHHIxvndlcUc2M96DIScOxHKCv8I82+iO1Yga
XFdrw2NTDBj3bP8GspfiBcbZH6FTU4en+tQ7lKyF0UJJHjGEVPHqURCfTC+EX4J1
KWQYcnaEY2+kJ1rLkZZuESqAmVa8ZYSOjSELmfSmOZqHgt7Le/Kyd6kYT1j/TymX
SRVgdSj7Y2Rx5wQZPFOl5sTvPe4iRobxdR7IOnnBGANbo+K+0wjHeXkhbUHpdIcn
bc7vjKAxjue0DQ1+lebhnMUn79DrLuIEDI4Z7bMIhV7iYzTIn2N0TEEmWDEkP5ES
hgODk0MEmFcOY7FsiHdZssK40/L/LuYxGGzJbtQjQauC/rRPncbnbWT2UjnOKkpF
aOGquE7ubpb9RYEMNdRTT35DTJ76H2IuqtBBeMuJC2BODuuvaVe62fm6Kf1hkg+U
cyujJGYraAoB7pNARa+Xh7fGPyPlZkhgAFI88dRBh/ckN1hri0Ioff7Ry+nOlg01
kuCzXhDRgaHWBI65ErqgNfmk9zcnWUEBpkQRGEUeuN6t39FE6xWHd6+fcp9AxZwC
eJY3LSUfB8E8/FS1I8vo7yUAOWff2hUhcEcpMhK3JtYFU/dctRbVlNfcRFREoAyt
JQsYgB4lmX3L8moktBrnJcOrjIQ7Gk19+4EPc/oXrlW5S1relr/piX9enGM+XLDL
xDcdY1/XdsZVwy6LqphHUi48lCbRRvH26geV276Wi4cxjEv7L9mMyRNh3JsEe7e7
vqmW8WaGUBxqOdO4JL7Fm0nLNB1G9uR9D691G+N4r6SBlhsVAstsyMmZp8oxbVHW
YDhH3OkTgF6CskSQYc1BGl+w1T5HBtTkcKTNPepWriBsTuuhkfq2j9k14abdvBso
J3Gl4XYuTaX4Dbu26/eiJYQ/zDGqsOC3Uc/tjlRqdQ5Ef6lDtbQI1bVx7UGfM7zv
AivnDCd8/dKdxGmklsuGlkrsx94V6kL78T0UU9GBCk+9qqaO0LSXKUFKOZG4sTj7
nGsJWhxCKfjlbcMf0unuY8HyqPwPxWUE1IT8jxlmN+BkIkQwzJ/FO8SyaEV0ipZC
T821nz/GKGRPr+kqrArgwdNzOTvJ9FUWVsaA5+zMuk+7/RfY1C+gS2t6LYSdW88k
vKgnUyKx+RJ7WYukt71wwqgmNrxIMWdg4wKbydOWp0LiRGEWapR8Uky3vNIAAVnp
aKn8+1GtTmg2at61ktrDHMGR/zgkv8nyIy3OEhahmjifcaMpyFy6kIeAU5K8kP7m
6y1Q0ou6N1OGm0nC2G+/Qa3N3cJu4QPKdGNVwbS/J+7oUV+jdoH1qVBkpHEq8gCZ
upGnljazwktEBCAbe0yL9gBh+woGPCOYyhqP5+7fznx0BxcgycD4RtTuwLVLU8aw
aQ4DhULnLXETPFsY909VP4JLAQNetwTUOg0ce/9uRhOdOwb4Ri+agb9U1F5aF1lz
q94yZmyjrAQryt9g+sm9depPN2BNVeW7fhuhVx4i+GxRdw0qvt8PN1G3ZbkBx4uX
tK6henFJYK19dKDKR046cO44LqX3c4njPsGGqSzPAzRWJ0yXNM/K3Y9fD/b+OInM
1NqlXOTeCHpG7teoags2W8NxxPmgMRyCcUNKWJmMYmwKYxEkMiH9yTXuTpiqm68s
Hnv6kkvZUUBzPBspHTlxlq+vFSiIlk6BlUtQyBtTymlWRzXOr9FO9epGTcaLfpWR
0spDmHAoqNr5+GibQ11ZKzi1EHM4afBbYl/fvEnYSZrmaJqZu1QYPjohhaHIgJrR
h0nGJmy/RqAo2WXzha35kuxwpTSgNSF3vCceMZKyYUfq0QI/FvORBfrMPEZZ/LJs
LZ36Hgx0ro4SfdOYmnnwgyWyTqzVI3WsXczLKbhER7lS3kZCcs+v7UAKu0OdZSiS
FiU5SQMGlrzATSc+alygoy/VIf/wzOEKYg4qPTZIrwdJS6Xtq3UcciuwrPIjFK7J
op+ueQEnbCJJgBv9o32p9krjCMtic1sLxG/TgTGwRswZlHo6GF0ZsEioxP50iEoM
BueJ0erpjGXA7D/8TQRpHiisowCc1CDZlMS5fXxueAKm5J3ykBj1s1dMB1UE8ZjD
iLiUPmXqpkqEnIvIdraxmBXIm5h/bZC1EcKgNu0Oy3v5Lrd2NVmSC56luL8HBOfB
X5X6XJzGUn92nZSq2xt5UiQszS5iBF8IpTVk5RfAOKIwzELF0Jl69eXNOABQAsAV
MkNsKm6Pbad9oFZmTpjTkMqhSI5R2Z0/D/9uc2L6iGDGKfws2xk3IprD3dRtqxS8
daHoePwaXbj3FnS7AtL2SRz1rcY14FpysDuaqOXGfFZ6qW9otYI8CBFJM4n6aQkl
v7hcUWcVC3jEyC9UVWnWycx4emNwcdpn4FWjUV3Ik9hGAXQ2c0npSCsSBoRqaxd/
C9miu3dN08WIXZ0nrweeHnvMzpMiAvh25QobkRTq0oZsu9B0bB/M9B+VMRbZVbqQ
zgb9CAdZ/8DElJx+j/7MHKnrso7DakYtEqzXfGsooUhEKfCjZQN4ncGUyAro1JJw
jAouA8YsEBOgKIDDbaBqpRZf/Foan1MY3+/+gK+R0wW7wK2vSgJwwLx3/sVXJhuU
WiTOTmt7kYl+uzERY6jdEY//VOQ8N/vHpob38aH/yxAXooAHA+ibDj95WsbyZPfV
3NXOpiv5KNsx01nJ04ejy7Wg7dW+XOygsEdY6pdZeJGYzf3BbZ2zmBKlCwbKm6NZ
0SpiD8zUl7GtPbqpWwAJzYKDET/QI2n2aEXG2gWyr0K4TNXKaIRv3F8LbH50GGuu
YSaufDtG/90ChKCxJ/Nm/1EX2elEa22+189Pnr75GAYlj9Y90eUGa4RrVwWNQRmr
CXvsu09UxRCIH6bkPT0dDGhYNeW6RMrQ9i73XjceDRVykx4DSTcBFtRpRahGhTUn
VZLLsgOIA0CHnYa3yMWy+MIg0AvzFvieMu2xhbnVr1FG5vV8W3NCZ4JFdYD0/xRn
upiJK+/0wN4qQC0f8lpKM3pMk6TUmO9hq4qVCnR9Sb0RBOOUzItITXGI46Kq7J9J
vNQd5AgmPZ8aQzockXNg33NXFc64hjzg4SeXew40Q03wn1ZQrqOFvk+xCy6KUnjO
ypKx9V1tWdBeaPbcIpq27Ose/jQikEZiKpJcqWHNRjRt+oBnsvjCcV3M3m3cfUOd
+IIk7bD8rv2+F0fRDhJRUXbDgZgMAUhAwe4wUCl2JoJQwb+ehvl8BpSbNuwxX15u
KWScF/tCViP177z+4831KRf6KwDNx6WsWY+hTF26zGN+/jLso5XhPrHlDs4SXz03
qjtPlAzPLaSUUzVmbTrQG8o4JNqW+O09+SdlxheXe1sGziQB5DiDxQEBKc0nOx88
umLIOopaeHm26NzdcsXMMVWFxlp9ltj0T3iWvty0xFDHq0QMQL+sEGyeJCqCGYd9
9TbfcjdVejI0HgGEQI8m93mkDyT56QqgmvCalQpn5cISxIEJ6ckGErE01lRUyEXL
daEu3cX7+4HbryS0D9+E4LdB+tnK1ysrDFejKYHtQ4LgCnv7dUt4segyjXaAGm13
tn+bJXDQ0RV+QMGEjS7mxjefHDEgm0CVJxrAYWoPwbwS0iCx7r7jhitnxXRcLdnD
R5F6N/NDRh6Kb4g5Zj7lkgFGhPvbGICIDAQ0TR1iuCrkUmhZ5XyCMqehNfMNQ/su
dMh9xXiaZn29Dq3EEuf1Qj3QaFzaoa2DAYfPoLKKxvM815uTOvsWrCRRKRauY8Mk
I7pfcCgXJRxaE2lLYS8n3H1hjLSgqtGUcy6rjw6wnq8ah977Mpe+KzX6HeY9MAbN
qQLH5tgT/4HtDb2JEDcFHqTYDXA72gMcyTZYrSuoQ4/ZnPDaG3oUim+k8tk4AVJg
2N0nVFkPSEz1HHotJh2HdnY4nSH2A+OWiNU70uskFVLqlrPzKXvy0oh9T+Lwb1oJ
Nx10pehgQg01z9Xyf0L1ijT5/57oAvYpLj6lvfW3ZPmvT9kOTyeFlv77+EIxKJdZ
BzZ/+LU2sgV+XR5kKYTp9ETAJlEukAkxKJegP96GOGvUZTf9tkGoTWfrtNjAHqP/
Jp6539ahNCqVw3K4/MF0hz6TkO9dBloH/8e7J45sPuulOHrt3wCevAHq9GXiHVvD
dudfXKSk4Bgkipt6RM9AHEEp6U68DbAwP9i89JdT7A+xXmtiFi2Hgk5mju+wxvzz
lRHAPLAvFcT/MJseFCF3PPblDsJ6s3tZiivFiaLHJVUFIsNruLMc/ovVq/vzjZBO
0SK0JSfp8mImRskHPblVg7qyWPY/XCYiHC1WjJot8ncAb/K8fjd6klN7mCxSAVqL
W9kyUEQB4/Vu2BnIPQSNxM3UicXUt3a6VCt9M0uuvzujsukFa/xXyhxCOirH1foo
7FcbVK1sp1DvoU9fSf8MBtjFJ/TCMZr3HBy7LssfrNjunlZvlnGfHeYQJVn/IqUM
G599YH/uLlmxgpsCA6/7Zwf3wJHXXzDe32hEWrygjqSXqmdd9si8bbDdQtTXQHl0
lYO3BrMmA/d+CrGJ992D6KUcXgt4IS5lSGnyPKq7UdW4U0ZLE92vE6AzmB8ey0Mv
EWgxADpF3g87yda6KWbviiNi1pNzbTOKrOCwkD4sAdLieyZMD8REW8vK7l1KMhVm
qt269IUaa7ETrwmqbattcZXUW900Lsoar8cHYCjlmvSZhKqfSJ8fRo1jdL9G84HW
EYugVB5FB7bBzNmvAp4Wh8BwzV3UFYzgX0keq1i6Pt7tYAhGkdOOv1YMO408f28f
WvFgfEkVOAnl+zKAv0LUPJxaOYt0YArSsIHr8vS4z6lYwNhyRvKTeBMdB/Ejkzac
QIz7y+81om5ZAF4ZPhnG+qARmBvKscXWUfadTUt5puePIY3692zNePuSZLwRvSjI
TiKXlwmuWqk5dAD9XVlDmVf64DFj7tA5J7wB5BSWJHrpb4dYllyxRxgbxp941777
70opkF5GGwx0s9aU1D78V8nm2X2HsnK7d/xdHDEA97kMuMTw176chf3D/bO0++YL
umBvOVcFyJU5fitzRQAWlkHGOo9g4Cb28/JJH5enE7+UfxobCVVx6gKp4GdzwsAT
hf93u4dTcKkl1XITJhmxeEwA9M3KkqJxhStTF3JdbrUttXhnb7HaKs75zdNn3drv
lZDUhtAwq1KpQq9Vo8XSMc8uXphEdKdj6S2+UoYXz15x31yjsP/PhS8rBJ3C6Fit
Z8UtIzXVs3JAumZRZNKndfWYibz7wBLNEEJzPAuRDrxDJ21F4CHAzyXnCyl1eCXt
iYAMZR7Nd/DzrHQwljSkxE/SVX3FUoZBIGvut9n4bV4L2Ji+Ar1rSzdH/mMZKH6F
E1dVQ93/7Ny3qqV7yb9pX7bXNLNOmoP19cWR0juKHYS44n5kqYIEYWc//vneinwc
ET/RmRIaSKlGY+VcDrdPVjSwFP98gvZVLDzAbVPSY11jeMmmIfp93zCcl1KacsCn
DN6BD09tlr2Sk5UONieVgUNgBF20EgUGUWWHObBkcipbih4/QuRZRq/qVK/6c/N9
q7k+czvrIdMUx99r1GRKurziKamXN7mFbm7xN7TYU1+SXVzesCSyzraHuMUkUZJK
9lBOuIIjgIfey+ZjDsFliiXqkETnHum/RXKsBevxdIU4jgVe2gpnPKuwjAiw9viZ
ZJVjpuEWfpWG2BvP0jZGXvY9dCuwbtVGdLEt/R0gHhSgK41Dj9W42PExNJ3nYv/0
VWXwT0YVZwrxKPqdsZ1p36E2RDAQaXHfTA6xs1pThUt0Lm70VH5MssclZVRnMKHI
4k/eWvgUOTTDrfPEajASGbqhKkpd2o07Re+pKZmB0CeU6/M7CSfWncLBAbrJ5WTs
LvFX4X326fg22BAyHYrRzKWy5etuu/0iANJ3+ccKWxtEGCv/cKzCltMhI7NQ8IjJ
a4MzVtVcA/6PykZbcV+WoGSqZgf5d90ZGnttmBcDgrqIb3e/VnETbasP7f4WdB8U
y8GzNuNTJRML5aACrrRtyLsGNQTbUNlOjMg/DwiHF92OAd/exMVvCxSZo36LXvh7
B/ZEJeWkk8Z63tRW+Paefz+1AE9RUhIEKVFgWspV2oHgHYbNWuqytynCWlcZvs1h
XovPq/ois4IBCJZ3Smh4TzohcpWzmec3wNnRH10CVbVmQHCXmqqdE9L5L65yjRgz
vn0luNfZhOxVRq+rsb9wnrG15nlUpjQQ1fpz5lbKcYNKxPrB2764eBJt7MQ1Yq9i
UkebmlKmweSIWVDyMyxY2GDiXSCmYxuqKBQIjdZnry6hyCHFGk5ifnm2WHz0Ccdi
udlXBf0ktAnsEwUqyE+TjRXqHIYUQV/QOGAZzL2hGGog+xyf2JcLs3j+z1qdlVLd
J3YFG5VMZEw5J1GhLjcODIThWOG9QTTb/mLXLRvle7nSeE/lAivqcZQM3wpZmS2R
fbL08DJoB/8vYtBPY2qtzf7AdudmHMPnzjW0TpF0Z2dA/YGcFtm7xLn6G7dhLbZs
DiNQTuGGwd97PiqgF/tlU9G0o2jsfajgZCV3kKYCVb6hIGM9aQ4DtkMU0hZivPOY
J4JbdQ3facf/ZK5/syiCMR5JWcIlc4x55uM4YtHfyF1ZohQe0u4ih2z2y8ODEZ5B
xRu/54wh1Sx/GWQ67GMIBE66UIit64n0pSSn+15t79nhNKCXQV7gQBx0nv3b++qr
Q42pYLUpZYM31a/5FXUzzFKYrkOSn7FPrK5ELecCAj8OZjqu668LigPtMI7CSrsk
iIbaByUASINMr7kap+ezF9TAgpzQDson3rjRGlb/6nNMkDDFAnW2bXDcLIw6YWTn
nyZJvxw5oxq2isUgRO9nt++4WUig1hjPhdLJ68pjThjUTHs4PTomIzqPV1nnaZjJ
P+8H6u3YRF64NKM9iFMZAqMeaflpTbm/yINY57h3p1XX/HRAi0DQi8ibgsTZo4JL
vOuqC9R2AfDzEzE6TbAoOJ9PniY2zD1og6Fyogc0B5mbcALhkMBd4xyBIJ0kLdhB
cNW5u7eW4p6EGcaPX19CFNamUQfZkqs+5oeXjnqiC9yozMKwIygHKXjk4v8rXwGb
sS70LMoCfuhruwFApMyCqnCBstHH+J0mtK7Jz/l8LZit84VI8QBkwTW6lUSIwouf
9NPb60hpbiclIumBx3dCas9aqpIEujw2PUhSz1CwuKtnvHmZHqATNfaGwlL4EB+S
SRkXK8OgEV8PQ4em/N0J3PJK1aLbrC3urWipknIMAktq6nVgaHZpgTaX9cT2Vkk1
X39cBNzkQ5a91feFiuDzhp9sEuOBd4Wlt8cc6pMLJ0JuyncGu+FycMBm6nOGk7Fn
cOm/tyZj2fiTMojoy/+Hi7niy0U71vjYMmqGG02XtZyD4eUDQUCekUM/MGRGtiUW
Wa0QjAJj66ZrIJ22z+YDJTsnMtvO9lw+TIIBQWtrUA7P8B4cAN43RJcJYddUQfmy
GQSmsamlbqTwSBxhDqiGBwhDk0Op3XGSPmRGoffwLShf119MI4DDMwd9sJKro+7M
Yi6PMzRNstdtYln7v4EiEtyXbJU3M/k4U2iuyF0Bk1vEw3aiGBMuZvwQWDwtAxBd
QP/cT2OVEzQ/98lILKPoxOdfPMwFUtV8hmByE9VKpvEW+ReDdjHhzu99JhpnthEV
6l33tMCoE2DRYz/kWq0YZme7Uf8LMlZVpqgvIKT/HZ5mJi2/xjNkCkj1hw9r/P3T
KcmdYDC08JpOJnTFOBaT6HqGmJQRdoidr/Mk3r7Gyp1kBT6ubu7RTIkZ7rv0la8n
PeR49831ZY2HMevMSl76oLX8UPF0bw4dECIMJ7z1Ejh+HjWUit+AIUIBPZR7Jhsh
YjZPqI6lompof4sRhAarRE+F4TAJS8D9b0vcGBob/0Y7zNoZDuXw1BVsr6O5/Pee
hApiW2ZILo4RY1h9zVCRAwedLJGy7HmZDyF9n2lGMHOd9lSqmd9oUqmotps5wb/s
F/DvEIHmnS4sb5JoWN1h/zW9EbwAA7yCaaUcOmuQgwuYBx5K5aVTFtoGjgtINctb
FzB3GQYIbS+rVU/QSYxD5/q+7GeMqg4Y1WQRxqxxGPd1yVNK/og1KLASfB5h+qzx
WcaIF8FqeHHeOImDBy7EukRAuOny8pdFbX2Uf2O5bJ9alBvC0x8aPJ8D1PjDcTGT
eja44M7k/SwmORoObynLMVvGzSOoFDrOG2Dat4c5kSHW1Ju7NmZglKlhxliR+GjF
/9swTiu6DbY0gsQ/0mfTdRngPcIzDG3kIN49l0BAoIN/BoJ70YVG3C7KmR7vUGJl
51Zi+F1JF5TbFBPILL5HtGEy0W2e5DnwRD93C9liQsku0Iut3Kovnh5WsHCioNAH
7WMnOoUU5CmboweyXe7z3WRrBi66Zr+70UFqoSS9SzcBvNNs3wLD/vuT6QuL54fI
zGloNMHeUVLzISkxlWbnrthIgLGV0/HilTJ4mN8KDM0zl34Ne/oM2eRp048AGf7z
ohIX9UyqnDbYAMUpaZzx7YahPDqakJUMFndFVbMdHOgjEKTvVJqrwyXmpruSVyDx
xZ5AEktltgIkPRnFemUHqmWegLRc0a3XD4IzNcr8dnUL1IJGs3j8zeNdRHjRgulL
bL8864TxmGevLaqsiWIQl2TsA1zRoWazOCmo//ubMtJ7VayVuyekS/WUuzQRn3am
1NfKynCgbhK1DaKTWfCD+yXNOphRNevTzNWl39USkoQq/05JF3JjQ6/0L7DAM8Aw
ouLXGQ+KSVdOQ2YkNgO4tWdsSszL6A+dz6UAACjNFgQTwXhJQbyJ1jgPRX86i+qi
3Cga6QCLUaQBp5xs2D0h5BvxEgymddoHYREyWm5OcpmU40TrYkJKwICOZ0GEg3Ib
wjVj15/GrCCqaH0rEIqFPmrGMyA0UrMJuiKNzLRwwDg4nZdbNbAOjw3BMASJEmxx
KBJTFYWR8h9GISLv4BId574vz+A37WsPnO37OA701h3hHsz0qkwe5MNOoXoF+CtL
t+C00C7EgqT7P+jod2uVVLXMLKAb18jUci8FS9kPvznBM2+p8VXoKXaRSw/JvEXc
m5QByHKKP3htGf4sjO82QXW88/ned1Qp9sC5ksKUjdcaGa6ZwFMWaVxox1a5ISlP
fmA5Lv9R9YmqHchrj76bhLgKXoz4eFhuufXcmRlV2cFjx1k+uOJa2iWSQLELAEhK
WUHLmtFdheI+2NabK5Uq+Q7oAgKDyv5NMTaprx2cCuclUE8D9+BdEqk5+LJF6B5F
xJXhIAB6zK3EuY3iFn5aKQOLHgYz3Nsmftr7FvXEWAPNMz+n7PKqBj2CqImMb1dg
zMvdW+LYUqcfO5x6oonP3GWvCn6qscyKQS51Z8gGV/ADDP5vCLbJfq+G0PuCWEdw
0UPSuxEFjN+i/JTgCtEJByqosxIP/Zvaz0AauQmloesi8nCmtl4xSskmxWY77/Aw
7UNSigFI4lWDAnxISwme7jy+oY450URAy1jnF7rF30gPM24NddvCl/cvnIJH7cjD
3P4npzMmTsUQPMkZD1g8aRagD7fSKLQZOO6zS0Mfbzrv1SIAdNBtPkGp4vV4Tc3N
PAy5ia0kNTcF5iZ/Nl7J+LH7GfQBnoAn6BzHiya1srF9UEppQU8uNz5U2vMFeEq5
gCf/0x4e7NhedWftB/nZ135H6CRIOMzeJ2aChfeTE8go6lXsevqWaaJd19Ezh04P
UpggLvJ39co9Hp1oCP88SUolVYyYcwCMUB4NFliuDEG0NZCJg9YD8fOqCpu+BSGT
DD0Yd0J4G4v0HB2XcXc+BbRdfR2uQIt+MWk7ysL2CIZu17g9JOtcqnWmZDQmd/Oe
2PlHsropRlKtugm62kZxm72aCKWMzHdYn4by3ytUEPIknq9BSo0J6moTvkvQKaQO
WLCha7qnWy5Yc/9a6IihbwYBFf+xK3urORP/Bnbba72820Z/rWBAABXw7lCsgzy2
mqZRnha7EvaAPKtObKjS9ShyhLD4fZuXqml9F5+qCZUmAL4azex4omHHakUAH790
Iu/HahVtHx6bv1fHegws8VVuXqYvI+mltutIVPgsM//+g3z3al44HchF6OBkZMIK
cCxLfI/5Kt/aMhJpvjI7PqAgzR7yLZhlyhAjgH1g+m7K+vO0J/J/TJJoPfusAMXY
ugzYy6WeIZu4iskMSgvgqmKxxiatLQakolirKcTTVPUlgofw74b16olPnu40gCtO
myxk64dqKAphIKpJsi4UJ9w2gNX0CsNWHPEJD23F8VYiO+nmZYuifDIxE6Z/H8NQ
ktvt7wKqtkdda35/BC6dy2zGtZfNdEFp3zu3ECZW+yfWTQLtmUUCcFe2Yek9q63O
86L3vR+AvuoqdnrCKxiM0qRk3qqHGTNtRA2lbbrOsqnhMhKKkFazw59y+JlS5NqI
SFr4yeklzw05nh7wEhxs/hz7fgN/VC67O20cuuF1vAbo74AUhfPKBz0t7aJnZ9bH
8mW5mEDoFhf9be07Mzx67GPV7kS7FtQaNf5MvBAyrwCuIUAaiautEaI2ukh+H2Xl
1+5icBnOgd3vwQciqvlpW76ZyXo6AoIJoIG1eHqaxjrolBTpQnpc5PSn91E2niZ2
EcjaWI4Zoikpdj2/vp7S3qATu+Uw447cADwwNodR+gxlhfSpWilnwIZMGY4UaRXO
zom6Zsho9ncUaktVMsPYvP1z1QXKiyABkv7yg2twR9cVdRs6GTeYMAdgeyz/Me3Q
Qge8kMXAjRCzvZroGZjPo+J1XTL0/aObuHRW44OB4a77PGL7W9d8CMTaN4OdJ0pu
/M02rHQrWw08h86IMi9CrLYPYtGSldOv756+ua8zzdJUfJpkDA/58HossJk7g6k8
ncrnhUWWEC1A9EROZTSUdk8QE7pKkTjkUQOZFfbIqvRtvdaaZQEV2Ogsgz1Hg1z8
g3sSvk3vWfG46/fgJk5Jh/1fKe9ueR2JRkCTPuIJXcnDvBeSm0XVscSnta6o+FF/
ObvdRLgQE9i0xoLKhcEzShKIuzeRKNA1yLNGgLtmutMMaxlFKUsNUO2pz4BiG1Me
ErEy6/vrPeIvQRXsjNbmKIhXX7IXod7wetGR1BMwIAaNjdkvpj+pUygL2MZKx9Gh
qXQZ1a3qbqEji6KBV2EUhhtB0C5cJ2JbU48R3sC8RvzLB3jyHFyF0jYhMYzDB/8C
6fbixDifVbE+/mHKyZlxL7A9kZhiWn49e8Wh0yav4JMyAhDhtdLiHKMosrcCvIIu
RGBxImf/Rm/JzuDIox7aEVnA0TNLYXiKzpU9Db7q5Psb4RRzmuvn3AQzSR98oYwX
NhKU3Hv4QOwPt6LfsO0+3HEPXvue7PzeKfCt1cHpLX/EvV+dJACE/fMCP+jMWRSd
W28Zh51rCjX1udOcRgKpYdtg2lSjJ0xYQ/EaeG/yN3/usxljBlZb9/485rNsu40y
fPvotYp0DA3WlibM+yoeJ4jt5jtqZ8g2rpcqagw1QdXd72IROeYbS32aa1Igw0YR
spIKzrsN7fiojx1Vx4422ZQLggw19kgTmcZLXw/0tIHXYgL/Il55jbFilMwwsHm5
G1Db0+BTAuOaENqhenG+B+jg2m2P/EH8TGkFflzFqhEFSShtSFtx3VXIhQmT7X2S
D/CaYWLWgI5VehGs0pydBcRWMv5jHLuDFfgYu11jiDDqqd7T2W8pAsbBW/XuOekY
69aVVUrDq2sczXdfUNulHdXO25QtTmtXDFhV6MZpy0yYEg/HVpTooJDlx0AKOqZ3
F2RfdJGRqehOOgCtVhZhsQ8NzYKhLFPdiImey2CDrY0e7UbJHBvaGvRAwGspCseA
laehKQdD+itWWtNo/qTc8HvUhYj61ATod+wtBoKtyC024lZvQBry0a0PKQXBXmzM
HlZXsv0jC+8n0QTZOpbOOMI1ZQXzkAYebrgOE0z9yCCzwxDzDLUseK90czYJ2h2V
JJL+sH8dSqoUqjc+BDIPAS78PbP8cw8JPl0zKKue7+iQqjVMw/9TsoZVKexHfH4J
JJCdryp0vyc0N4w7jfNfcENsJ8E1am73BH0pmx6kHtvLNXk/AgfXVXfM8qWAhYyD
In3DWq+N9fb3OewQ+yjUrT8DWwKFdyAriW91F3AxjLgRzq/DvWhb0ZEbySKNEpK/
SBaQixSumxUX7YaOaQBZSTo16MTTs0ruCgXedtDnDxRIgrpsxIbCdjQKr2GpOkBT
5aNNn5L4Iy03B3HcC2MhK9bVOqkTTweN+ahDax/eZi7XaUv2lz+pZyHflKRqj4nO
aqMJajR49U3wlpszHpGhKhyQbcvACc2zsQhoT5i1SYF7x0dfUA0KRAta3YL+ppd1
DPsi22NuOygn6XCs2t8Uzj7iHPxvcDUlsJC/iOx7m4OLfQbZGn04bqLty/50gRLF
mORpaIgzvIQPICphA5rE8Qi4UetDLDKSCtXdXIjQMvdmIegLMTY9xYIxbQszDkku
5FukZXVje/YnlL3dngQ57O2jwVNCn9jOrK35uRm604oxaF+stYuwmoQzTRAXOaMp
4/KKLi4h4thcU5lvzzxSiMCVuMGfbVZCI3DC7skv617y8NJCryAqA/GV+8KKoU6j
EakR4LbFdEVrEZ3RcbrjgofwIzTrbOD+IvpLp8+37RsfFNBHaOXy2larSc3Yp46c
TE/QyZUodvQVereFI+LAXI2zH6crzVi1pgG+QgDFT0JbJoOl1XjgkuhO8gWQhIFq
uL1YCX7eWg/pUbLPVraMF+TGWVt1W3VnCODSkypcmGR9P3mV5o2ZnldBB07XpZA5
0uc1JQ3tNQLwVDVunAcf9qajqlJvxPCLcjvRb67Sj6V+mnKKl3+VQyVIChjTN7/y
EgK2t17H7EjG6S7YRhMPfLFmeofl5BPOpObKkgZ3vyu/fYopW35lWL8K4agJP5Nf
0GCVljcS05bML0ZvCktXOpiLhSePB3BI0R0NQ02S+R7cN1SgVBzxi8ujT8Bcxv9D
ZP0QvRgDDyLrZSYGhHZuCkAnZEgrRMSN2q9ah2yHXRsylh7KArmq12ZplZElJdUt
OJ2EH3HkzczAfYLkeDDLT75vpvya5mZkEw1BvhflZkka9l45nw2a/1MZRCcu3LZM
FIf6K/ev0g+NwGA/vxDdNnsRz54N3b/nvZWzJ44JRZJH6UE7ht+38tc/gXgLFdYy
nj4lpfyFqTHelvLABCsL7zLgf5h1Rvo1uUJ7hxJCvF1eYKQSMvWwbWRC6KgIHWN+
iuPG/8ohEub9LZX2ok1dAojkh6DBKMMR0GAPIweYVC+lxXd/hLMVsUenunsqCWMO
3BnIbRXoUw/Ldl6iXlQY0/YmlyhJqBMNIu+6GSfBSVP6A1E0KhS7nc6FD5h054P9
XmU39gkCC/IDE9b4yxuF0jmscB28atj7VqOVm9LCP5iTNUJSLJYxjEZlfbdj2yhJ
JGf/djqmialzkqV3kJ3Mh+agZZlEXrPT+bn1qZWKLm13KuY5zEtdAnWeHEyGPeLG
NQnljhT3uQOaF851wqygLIZog7rLo5NEABn/EP4fCZw0NBJoj/xQZ20rVvcFqrcE
91Y6Ie3w60adUAkR+YomoU8CYFvuFxlv9FTAojZWxVPu4H82YuAI1jPDKrBTFi7W
Kx8rARqe72i64YoHuQnZnXohyFqtwHhptxF5xpe9CsOlmdoMBbvq3gIXbjUMmsCr
8utT8zs/ONTKLmMtB+tzRLq9o/RIJoaiQTHX2IFnQQl/RuoSpamoaxIvBtYHOTP3
TKa7CDMmp+K/N8tRel8uKdXYkTuA6iaWZEWsNavMBIAuKkfQt1Nq0I9fJeZIiQZD
Tndd1v67mR4ATGOyi5BQjy1hX25/fMo1+QI4oDpP3VdFcHli98gdz/JKM6T8WlP8
z/VBSmSE3afQzlxpAEx/YXW6nrZ3RKRB6BSX3csAnMi79Btn6Fsc7puPUClgliYd
TOCXNkjE2qVDNecHMSktSpY9WcBHpTUw21ChfXzLB3Y0xa68Vht28d44BJDedlCd
sRHThl3BzX/mo3j/415MrRmpGaRCyyFFbpe+eXRr4zRBiYsFIlY5bze826HElAwk
gK2RjzG8UkHnAZYvyJWfBTMXfQTB43kxJcKOkXymkZuoe+V6W3TrJcvy7oNr43WT
KQnLylfYoNVg9Tjxi6POGfPvzNadULf9vKkwnUYaDEfGOGJtihsQFykvpB7TE7h0
aOZx2UlmlJ3WN5a/DxTiZGQdtIRcAkYx0jU3atESPc0zsLfRjAfV2/EZyqkE0Gqk
bMBBzCrJR55td26yBHdo7e42cqHObrlQyj00AqB5JAqlRLrpyQZRRqvtvtOSt7oA
Sk7JVEPp3ZvNf+j+CuR/FFBtOPCHPrP488LJOORtsjATV+JIlecVEOUASwYVkIw3
RYPeoj49LBjEzRs1U55BZ6qkzwELcYHdK5D0ixe32t5aRvhO+5USUOxq1fTCQuhK
jF0zHrToO90ntH4jpq8lgikVE1Wr6j9hJbPQI6zRPbPt/8IaxmizD//9qFDFrJIW
t9lUzTu6xqyCG4JrEBpk5F06MZTR4rT9AnW3P5lxIO+kZWrw1Mybx7ylDLv4TTMN
u8inF+SgsUOcKqoCyvNarNgxsRmXqBat6HJ8RgmkcwV0aDHdj5k9j8wdkoRrmChK
q6adnsnooc9rLJT/4KbgIHR7LKHRnswYNAWlWg+8VlMXjDUMiVqL4n4tE+NjUbgG
9IUiBZ4zDsbOyYeGU+XPYkeJ2siPi0TSNFjPe8gmQXCdos3rRCErFszSmsBlq+KL
KQt7a/qR1fBt6uzx7DwdX9dMVKNzsOThUPu+Yx8w9K5+ASpj0jrR3b0iw/4eQ3qQ
2Qb4g02jLDQkBFWMvdxM/PddVPDdkm9Usn5YL5Hg5DwvvnE/1BkBA7vHXiuosw7H
y3WHCZhCnSAlp/RJQ+TLupTUOlgwQ8E9JgVT0hqIqMuTWK5rk8QEA3MIWe9gxkGy
H4zsoBW5EOZxPrHUxEJxeOTvSFAm8Dzla0q8mxQudg7QRu7oeh4z9cOdGaudXC2F
GBbJgWDExwH1SN0zNhqWBcm8axe6/J1LXwXXu2oJ06pGEFD2KYlVbQzCn//3xLl5
jQ8bJh8W3ytBaADm7+6d3C586D3ePtPnPQmp4ok0TOAWSEtXhfzke3r+oay3R2dR
xlcIXbuT0X9dUqmmD3lz0YxrSb6uNTMqo4C0ngNJ2R5Juq/7g9WxLqchNhX6hkDE
fQa/WM0juxmYxLjBsMlGekOyryFEi9plOYlzQ9B4IAHVKhUGg917vezf87k5t4aU
1c+cJYbKdDTjlQH9OmQ9uK4GLSubSB98Sq/c3Vik4AbUpFlaYw/VB2TOG9JNWkH9
PQBlBdTXFT1Rvelwt4nKRqpCnbmShfUxVdXMvz9vU6dMxueUUG3ZFHEjAdEOdWzl
wa7dV1iKNGgQdrVd5KeiGD0hE1dshdP9TRbFen1jxLFUj03KYuuZ2xZtQj60f3g5
UyJ/EhAtOXn2WAs1HtXc5P1AnEDsoVoG8URcCdyPZGN/ffMwh48QItN6xeMch4Qg
X1bspIb9kvgthfc2r0XlQoZN6BsNGXMhSbn3ELEgyIFxeBSbDORTixCp/JaC1NUJ
g5ierNq1fhmIF8HdhxK5llaHAxNv6kBhpTH0b/n/mp/9Rxd4f5JIMTHdeqI7Q+kH
SOgdOe3Zt0Mhkc9Nt60AA9g/JzKW1Ibm7BAKXRJmuNo5Sgb2JYeHSU2UFVQS0MDT
BGKWcu19MuNvk6OTxQtN7t5IMjIoORVENueooQKy3IimdkpgUDPpLB57RAkL0BAv
YEVnodkfJFdji7rmaSyeLlM2kLOCQtPyZD3TcqSPU6V5aclosHkC9YUS8DhoLMXd
VNvhD1bjbS3ssnE5roDSG48TIPFXGgyJ/JcSwSeMwhP+X6rcX+NdC67TZamUpYLm
rM6jxS+2eHhzmSnZnrbdSSX3hpDHuLmE227nqGzUlYkvxLNiJ065VaNYf3jiFQdr
hrrn+bNSTHV96WepoFSzb5Cmb07isX75xLVfpgX9AkSfQHkKZxecqrwssvdAtFhq
o8mvfSbAT3rsNFsfOwjdPRe0iaGBnpMOMkBYu/h7iShxNOyjg36WMyplW6o6gOpg
e0khsPbYBNXxh21mGGQJz4NRPLoRD8q6mKaZ7ejcHxcp1SAE1c24Fx1djQnDuO93
4KgFypRBPr8EEEWUWLXGjNl4uOxmqT57GpxQNa+LuPipbo57l8pTULLdMlOlYtYi
UaWZQTveycvgs1wQm6b3kgiF1Nn4iTQuVfbWvUpOORgauBsNnRwYI9JK5KZJuR5j
TMw8/0HBRnXIvV/akVOIkPPo342K7F5mySVcRgjxoyBX/5yyNp29xQu39FpWBnQ7
/dwnikvrgj+1PGnqBCIeNJyCwfnwDfANSTvg8lUgb60Xp3IqQSFLTwSUjo0g+ziv
Gm5dVmws6MWAhe2V3eztG65uSoBXE8h0Ly/I64NrsMOX40VVgyiQni9w5fY3o1JQ
5vb3ZT7LeykK7OlLoLulSOW4Jwx0cCcO7fzI4QJRr2/4IjvZAsWkLFAzw4ZmV9G2
goJHj8R+/7LkprBnt93QNzpGEieCKFE1aS52CoEA7LvrxSrXqerpLN2AvClss4Rd
3n+fYFwyQ6MpywnjOM4g3VaA4fIp9Xsm0j2SnnYmZba1E25YdBnu5bs2Tc9WBdTD
36Tuk451hSWSPgEx9SefYBs2gL1lOoVTrdjxLr3dLratKWnwXtBakjHjBIGigdiw
Uo/KDEMxE3arEoMT0Wn1ejunRwPE3Kt/naTHJOcvQUy9T15BKx0flP2L/3Q/6g51
rr1cbGbqgcZLtxhftKgKYQPyOZBQWL5CQPihrZ4pWZ/vtQNBiVJZP4VFEep9UtFj
S//QuJ1/dI8B1TI0hGXnj7s1is9aSSWSaXmp1ccBlQ4epBdcbmxQtSejFRLX/8Et
E54UbJmDGb9qCX+Qg1U8hh83yx2qsnXsDanHN1T2RD21tupXDJyb9CrS9dGdNx2i
OfOWwrdapLPWrG3x4+ZsSI3JEsT+9aE42k0ycJbEOym0fT/rVV6y7p955b7o+Dln
YAcrI26sEEbJpea+BzJUUm1373JiLaZpD+6LGwCKn7oBJt8zzYvJwQLY49/bxBoX
WVi2ThIl6TMSltUgBBNhjgCZ3+RhArrxn0q906oBxcD0bkbYZhwpL0cxB5cXODSP
HKGy6VOSdrMqaKakP0GdqgcW5u4sU27oqj4WH3ltcVPWI5yopip2ny/KLAm1khIO
umCvbuRJmrIcrlq3f8g3lUJStuYg1SF9HaZIXLNHOFjub9O+gJGK3UzzSD4jrSXp
e5pD0ZIJ4Vn8qawrTdUndFOO0j3nxr8Ip07cOJJI2+zBbNaYPPyR2D13TWHtJvih
0xMBMiGi6mHhbelXEgg+1NIV/O6xMa8XFJ9HopENeDyaC21jVYzC6Fz8hjLjtdzK
t0Zg3lvP/YQ2q/YpXou2+E4ToNo3j5JLHA2Q4XcqxQKyRtq6v7g16eukQzxDHMOJ
K/FkT68mSJ1NucVL66C1E6FY9sjb8f74FbPAkV+WyHnE5aC7gSiVCjBOe7EpJ2Dy
s2gmW9VFBAp6ekC/iwHNnxbNJWAxMnsOXfPE/Qh+Rx/zia819gic00xi+A4LIoSa
ToIq31ne0A7+Llui8dF1nyOmEVv6iaz+ZUJxjKzIOGFS0k4B0Z65ZgSys+39RKrS
Y1DKqjCKbxYWPGixW0WQHNV5GMOB1tyewibR2gmSDxhhmrZaAXpGt4t5KbBZhGTO
+8giACymXB8n4eHGc51p3NGTCVccmCuJJiBo6U+RKTRW/+vFWIEZxXEXUGECDgAW
Asv7emmgwrPbDGQjT0VSLH1fEkQBmjMi/q6y1/jN0ZM5LzQjhpvXR329ZLWuGyeV
l6+3S1tzbDYHKBgx3+usyq8TnSC1CupRQpKTs9Y5cvX3dk/kA2Zf+fmGXv/HLJk+
QI6nHO/t/HdeGMTQO6o7gcPnirXyRwcMQyLln6NQQSPFYr00sFVm07N7NCRJeRhj
f3e/dF669iZgALaARNt8b7Emxxsp3RDKOqyfKDcnsFRqAQ/t+V7WB1OVE1GVUySq
FGpb3uHUMUKt22Fr1Ga07T1OZaDqTjJQuiGMkX69hVU3iEYRJeB7+ZUAuaHVeujI
GUZBXV2lGAI/exPCEcBgo0mk0T/TCl94ffVfO4nVlO6QQZtmuTQuLvS5X3uOOU1i
Af2YHm1WdZLPZ4VQ3F+4ozSfs/ALfniRVe+3oms/+2fRLwbTXsQh5M6vNXkHyOxb
J2ePN/RlPfB2yrBEmgovXeCqbJRMDgDSi+zVzg8McmVk8KpT8+zqVBj39AHr/mcn
zq7aeyRzDawiiJgj3BeB8TQr5X9BkR3Ualqnfnd3jC+az4pFgsOaHkrONG3vJzXt
Swn7S3D7d6GqRDSVZzwRKTZ56Q85vUDs6Y+MZaxnPAQU6yMedRSki8KVDNbWsyRC
EtKcpCKtqatakOHCK6ahY/LqVXwx1TWU+PYW6AMaoubIQ/8ooOgoXMAh81Ff8X4f
P5Pu3dHksr78dY7SrPP0jUcYhiC5aaMOxhZ9YImyi2+4GEzkw9k0SsGxkoUvfy7O
lZPXCCjJv8AVG/2oAvDb//SUHtCxDBbymDbvrjGamAaTLtv01SBJZOaQAX5IP56w
07KkQEu8EYAL10Da6/N+b0TMDwrHg4XEeKrJ4RVimvLxc6ZNVRSGxrCGq93Qjg6N
kmM0oSbAuG4Fhryym9bflMMsDay5nn+ZIy5sLQ0JSXJBIIrykC1I0K0Aoz9SsSPR
G3NhJTQ3bk7H4yo5NsdwPFzfH/V6/aEBQ+FqLLsvaAbBZYDKY2WT06jwHVHGw+00
hgKFwLK4nid5gvZ8rP8eLjVXOC3TYpRVMiKOJmEYTsf0Pe2OxrecQiAbDgcT9Gnv
vAbh6Stp36fTHTR0psyk+8iBC7yOrQKxXSVLg+4TA3qQzocynjwr2kis3z9LJgjJ
/5IBpUVjw+sryfac5rqdzyocRvSXCDvNp2tBMuZA9LxdlVKA6W5PZagG9PrBfboT
nWpIGRJVoL80xRY1vuk+HCUYibOAxLpEO/AD0fpNdOniyR1vtU4NUJGwJHiJWgIh
kwYquJ0net+EppedUEFDEonzt/WHqm0kHD0DHnPMuixpd+xplu/hfUQhRuZBNSWj
8Syjv5Le2fhXbWP3C9JBrPrKlr5objYWyocxvUnd3hz5ky+NqaHThFn9dsjKd0OI
UAn8JWyScYEjuljuzS0pK5IywR6xYpv2ZsDhizaLx95pXKmjGf8PU77ySq9UGHNZ
9LWJ9TL6YJ7rPj7y/uLCOL8+CNHAWM+CaSXjOmZTO7RuW95FPo1B4Gukfac+dsyW
QwjqFdl/36iS7f41jS7t5OelqGMYo4ePdk/A3sI726i6hUMEpjkLeWOvPEtCQ7gR
RFujGcJDD7EXgkaGgtfkrk63/AYIsNPgtIi6tUBICn94OnJTfFQtdkf/3ZXVWyt1
/T0wNrPVI/SJ3h05tyiI3Kf6MSLH8kNBLOo2/coya47GjIGCY0uDR0BkK9nbm7Rt
LNK2jX7sJ+ApcjF20uWjpqFmmdy+k/VpMbIzy6E/sIWD0acMdXKaVVlYC7oLYsaH
PbQo7xyZYg81T3X5xusLdGC4jBiRwnpoOVsFhFW1cllFlmcMblAvmsdI2STYUxJ8
Jor+iJawmM3QnlS2ly+CkNeNaBkcOpxlIzgNzc4tPKbANkiYQzWI4+Lvzy6fc57H
vMGUztWl0y6rt5wPDj212Vxl19aVzIqdW++f8WShs8vo+3ZkvoLfrEgmBKd6ma9m
ARlJcwDKjk/ZGTrF5wp8RGmPB999fXpWHfUZMMaEalNH5u72hDo4EhrZrOKqrjrV
k3b36A9sehoFn1TImaectAc91qCuPizuDL6z5rgYOfxjGlEcKiaK6vy7HRzTlNwk
FS55YW+rWQX1Et/xxvNLg5vfWPwvI+2qJ8rLrwsHWlQimhbTNDiwkWW9gzye8Aab
wQB/kAhhpGmbtjdfo856AgdqNEPp0ubF5cdop/WVa8atf268wyDRlXte+MXB1cHS
K+t86E6ccvMqOeMTeO3BXD0qi2oXv1fUup41hpBSHZsXToxvZm5yGwamXakh/gNd
OqgnyKU+8ebKGVWKxre9fxNGPOPRBcChrh0lWFFtu423OjBV20+ktGTdP2z2NCQk
8XpuE5bKVzHmksM/9CFencYoIPyEpD64I6CSLnC3/o/DJxLAeh6A1KDByYZTRLoS
GoOcwsSigExjlusjwDKq058KrStdokxP5GiSwbfRdNqvf9oPpPWq4kABcVLAfIYu
7bGBrqbXBZlyZ2awNRsjAan/soK1C6PXRr21yQrFxbuGwHAUFx966EV7nuTCL7ps
mNPhRouFmkX0mS3oOJoK/EK+xpAkcl99hAJ0nKIOaBxK3iaZbzEzF2YbOdQTeNRr
7Sir94W5YSv9eKAi6Ztlg0oOJZrbzIGQxmJ5dj1PeYzR9yKGWfGfEHEQqkss85pb
pndQyGRMOH46kJn3UNRriiMynE9r6JxT5TAIklBo1TWBhT4tzsCQnnlaoNTMp+N0
f1zimV3t8YAMYPHuyKTnGxzE15GNRNUj3G+5m2TvZ7OwcVHzJnlKH/FzKflMEtgW
c1U9UoR5lT9hXoKdaliR/C+7rckROkGfxhThyNxSsQcrHxe4nn5JDWTbkRO65MFB
77DpPj/sc/sQP3kf3tdUi37NoNgSi4256FZsztohhk+fVVzG2cwk+WOJe/G4UTX8
kwkXn+GIO+JWX9PVCfAL1VyTEFCoCdoQIuarI9DA1JG60WjcsK8V4EciB387lS5O
y5oQCs7fP2+uPiwk0FTNUy27+lUm8Qf23rU6ZkF2ECtOlxQau6Es/otTHa6YgBRz
FGYHsvkVgzjxIPcANfQx1LVhWIqL2eX8uS/RXzxJv4SgyHVaqVYxSAa14NCwJZR9
IaB2TtKhmOQA4YiTUnKyAWRNXz7WanRU+mL8OogIGUZHaaymho4ugyls5/jKxN6r
7W1JAxeQZYF5yWzSK3AEgR1i03swIIQ91XEygLfGjITllIvBkFrX3iJxoRBNX3t8
E6I1M10K6jHeyyPV9U3XXlKvmn/c2e3eDMGD5LqfEXn53FxYOXYMNnrQQLzRJyHS
YG6GLF+9/uZPTrPFU6jDnAedb9K0fUawWxxnU3/SjsgRh6h1w+YXrCEzHV9NKuBn
ZOUrDORt+7IObggx7K8TlPqDmFq8C1LP+xx0vyn7Zisj92wk5/qKgrroy7jT5PZY
qbSKvVfUeUBQ2sXnd0nAgIf4qjMh9O5jVOasjIIuPvJ03U/RgwHMlvQ6cH53gWm4
pApiglQVwa9Yontzc585oFKKSPUsOwkm4W4ObrqheVflPuaAbrh5fkrLM9efmhrr
Ex0i3EhzfboHeHeljB84hMUyal+jXzaNkPGXQ/dqnx7JCOr47YjWeFFmK76+lngb
oCqIepM5x2XrFp/NY0d4s4ODi86+2Ds31GADZfd1iu3abTm5KIaUcR2WqHc72XOv
/R2J7qvywZH2DdxCUi9BeDlyJRLGoNlVWBI0flooz5MEjFJm/j0q7REEqkXDCHqF
XhxaAm4saItQYu0KJL5LHtjxjUa9gIFRi1c33iycD3zD4Y0c7lmWHsq0pKeI6QP5
Jg3vDGX48HU8mkK4MPhLxM/elg85vNnEGOPAbP6ejlWMOkb2CJLcABbT/QBP7eRj
a4qPxV73c6rGwWahPM3cqOBhxtaceG2mLxEinqPk2WZkk59NSm9kLumuH4yoHIpW
uDzeDE/gK9Ug3sBMXoDGirx+vsmAk0fbGunvbPlm12QQBaBFInNbUERpqk/bE/Ls
+fw45+e17O88YnzF7tCngTt7HthULICYgXEEKFX2sk36Kaplk30DYrkKTFL06Z7Z
v8uhLetHpRchb0ZfnS2CBYg0x27AW2xsk9k4bPOmmFD50xClO+e2+UlXaD8bTBtx
tiqX3PZu0efIh3rDX/AWmTkggPas9o5JtZw1jYsorE4AM6F7iuQAZeaeQHNpIJuV
7nl1u+Sxb2DuLxjdNtNRLsUwVpDFQjKw7+03/RQKkgYnUbHYC1wm4Hb0KKdLQ8/1
WBjLXjyldE71bboDBFxcPInHyT1fKCAarDtkNsLupTJX4HnFhu44jBHeQtMXE5g9
brNlzCWmlnP6EnUaD3n9T80LxoXoxKIhRzrmPWXxXYrH9XNl9JLdUxltt+mIbytL
26R08RrvWSKjJ+wCqpMFdtC6/IWFPQ9S/8VSptX4/K2cJrRuW676JvKFq5tpxH1R
NSqpXB6MqPr3Ec0l7nEq0a9FTLFHalveeHxieqWOvJ0eAb1/Vnz6He6BsZ/sXNgS
9IjA7qWC2oEFlZt7zCzaU8irEehiaOMpNGbd3I0IJJPAr0vm9Vqmhkv/smth2B39
XvPM/+MTJVazJw24WqquzhqO5U+5orD+9W9fb4GXCjeJGHnMNvoo65jAKsMC9/Dg
grvrE4I/b+16YMvc0zthRYrkYP8gAyjnS4M+iILH7rA85hfl5W/yIZXYhJrJi0A7
OsOqLJMbsh+L+SYPcVv9tEoqINPbHUqwq4hNu7Vl1BLD/ka6m7eWKLtC+gL8ejmT
BQ1O8OeGCC19NHbD9vzmXmtEIOywRzjzOuUDpOuSGIGAn20tvIp+J1cVcZRa+pMn
wjPL7gvLHv30Z1UGDD3bRMjh2hJOrAM1ZSapiktq8ePeqbUDE18BTFgjcjZPEzif
A3/j9x2vIBHiFKcKvV0jVe3nD+Z2dNeqv99CEltPFW+KgPOAhwUdvfnVOYRcG5ef
VW1DUnL/Ud20MMW7GbIRjKnSJ3ux5qYW14qOvMgI+bvLwdanleHKuepOptUWFjCd
jRpYagyyYDR+9DxOdSdgV16ukpme9FmDeIQ+nnQyvQreu/21beYECS+n9RYi+NFh
dazJhIFf2R8jIJ2vaRtCpVjtPWOWZcdJ3q6fScs6L2Wb3PtPTOgP4stxrzhO/t8F
oili426DxjkeQrTOPv0AJpbiZtAapT1BXrcXDNE77Z27c7q48ckMAl2kVu4/3Dgp
qNbb1t8xQyxqj4crTshS1id12nDo14M0GonDShH6zECDP5pjF+SzOwqdL+Lu27Kt
cjKZdDKaoscoO6yQILOQLGbSGqfPzJeoaY9g52WeZQVwLaFavXpj21nU0hbLKZCD
CDa6+p/gWeh6lRr+dxHZFgGt3SixXjSw3IcruWqafBhnFDxM0IrJplm229TQy16e
Ks/D52JW7+Q8cDMZI4RUflG901T2MldmavhCAjrsYdEmDpzaX7PHJjRjk6gpy5UF
DnDGPLi9R0c+0kefeT5B7bpZ9Oid4AteEUM/41GUduG8vrooyRWxF9f+y0YGY9tF
/YGVscZutATa7vRrtk3jCK65VFdkpBv5Ssn90TsBo3AGlwTuAWhMbMnbAPvZ3qAj
I6XdK5cfhPoHvN5E2M2dyefHfICyySlUh6+AmLaRCQMl9tSbmyfIMeyS6s8ung+L
wG4ScOF3JAIlpBnNsB3RrlJi9lz4Ac5UPh4m3XW6JfV9Sk4qNH8/9C20X5AeDhew
GsPf4ROAXIOtTm1yJqBRkcqezmjkdjYBK0PDBRzhw6b8aW9z1j/bEk76bld4ZKjf
DyrnyzdXirYGe1zOO6uSl9sP+8rJ9UGxECC7undzka21s5Y7UrpzPSsnzSfw5ebf
+2v7XdLbo7ucFTsUFPjo4DSSAAhoD3FRFpOynJKSKXopn3qvPtLHITnjR+EKqGpY
Yf7KtC6Wneo2Yhq2EZSjef7iep7k/vBKW+yx7t9XokU0HDjtyRQUiI7w4T+hqr44
lGfNwo7vo9uwpyjdEHMmekAU02WQixsRy2/+j3vYPzazXFjZm6re610Ep320uJEx
JR+Jlfo/3/kOo/SZuVGWmgYoMLVC+VxlJyczNoXirw/GTZ4egcCuxCaH6XOBA6UV
vpaWMXsp9ysxs/UgTPL1iX5+qDqVvtA1AcuQwtICpDUn8SbG6fFYXP0MyqGqbWvz
EVHfXYunz9TqtznUqSDCG3r00kmWygjbuTXEdSEWAeEAdjknlGu17wsWF3S5Meze
9FVtYQdTY2LI+Zeaj+++I5g7xuoQt0kaDC5dvbHiKbYTxqLXefkJ5oZUbfbVSkZu
iHFL10LNz+lyk+vaxx/agHEVo5k3Nw2WQSEEzLROs+3H1T/1i+o71giX1q2HPary
IqsT1C4RUrGfVgViKU+AYcnIADo0Rs36dYyR0BGFfEPGJR7KL+W2rqhOLdvXH/j8
nTWYS0nOlEHYhWFBNgDQsnEVp/lKaFTZDWNonJbSlGeG3ghzkfbKBzCHB9qPHiTy
qsr7GPwMu2YUA+M1Sjil9b8x+Txnx1CEA4jlvaPUUgmKPEzUkejcp0yWugXHnUil
ieizS3FlB0n4WRor/BTXVw+eJhdH0k54+sjCd4IEkGp9mwElxu+wFFfb5ohTlx4n
pGZXGupJmAA3pMwt4CSi/AtzzWbSXSy6V3sXKZ24NwdJN6g9F0jdkragUNh2IHvz
pEfdf3sZnmj3QSabGKcNIvaHBCqwpj6q5BOXb+uhjZ50GggL36/ZUGYl/63yp+3X
1SaQ0h+9aIe2FaSh+NgRwLmWOF4o2/MdJz7yhnT07hN55QjIqJJEDc6vUo4CXo7z
Kd0uXVmp+xCua2Kqdd/XozXcnRrSq5OUr0uJnObwGwPJ1FOJeY07C3tdUqc3AjFK
wdyCcSxJj6fOOA9cE63qHIBAlAPTsSjR4HV0zkTPzgnpItazE6Fvkddw0lPnKRio
7WECpLstX4Xt5BGBVheBvNJxTSwRgoDysGoIHgUn8XPHe6B1VdiBm/xnUXDZ2pP7
5L8WgTjii9HagYVUmpntOcvW4BW1CPvjsxWFRs1DsB5gTpVyNuFcqov4h4FyNUfs
x9b0QSwToKOp1jg6lAqTdy1IppZeF+vSOBHZ/8NLXms9oniBm52gnb83qJZoxcjC
vyUYB8vK6/gnrfgfWEbROCYLqh6HMwQLTaSg8KzF3H+A/ssy8WMXb72Pjcr8L+sT
SX/5n2X1f6w6WI7P7go5p1GjHKtRlM397Oga/ydB1xEq+BhnWqPt4iclqNBqrrkV
g7it1JMnGK4Jgr5jj5iF5Qd0cE06LO6XAczeobML4OV8uKBReAXf5t6TkHBN2uqg
yaDwOju9ZB6mjlEvrKYMad+2x3jYplaWX8sy8MwgE+vr8DDsVSfHs/8klkllTwQe
1ZGOX5K4QjjYJAuZGFD2vGbRsyBf4nEE2rbH0DdlnmlGuNibP4KodN9eX18cHB2B
E2TdwjAb7rYZdoM+hcrAUBZSKzOkwD366JAnQATRyzc5sU3gMca4QpAYjv1eFeN8
VE6SI5Q9fsvIFUeTiayohjc7G6WJ1wYCqt7d6iqwR4kjbX2oAlySzpFQHxkHmPz/
iVgVVNx/qSmr7vpEEcGicSHiCp74vBX6fM/OGZ59tFsJbZL5hFqJt9lX5P3bcUUQ
tRQQqYjNsQ9tge7UepHSw3fgIoMkLhZEjzYCLqmFhuM12otc5y8b90uNHZ39km7p
Kt/QLR5L0J1o+4MAu1iomD5ADSP/fpCFBAzVbdT8konwcE09+WujicIgiF6NhvIH
8QSc8BFvnFLnBJ20xjMaOktsbbLygDgs9Kv/+lY4PSzt6s3lYpp4+SiUqnqyyN+6
xwQEVAg76CNXTQJi1vi8SkwG4M35RpDTNnCZyVIQ9GnR0tTi4NSr5Ju9kd9BZl43
H7NqoKACDHKK0PL0MLQJ2nnm4h9PaLGS4ULbyoEXBNN1EFra9iQOw0tcX2fSKNHS
DaGCn1dI27la/rCD3RyxKAWPgGA6uCg8we0M5jkCc/mmrWa9xxRPGPgGzRMjIXKU
ZyK5ezZRXXYrsXX+8xeKdZF6wUOuxdPIpOTLXIOoK5yyepn2S3wk9vz16yRXNSI3
QS+rApBGf1fDB88zhaxCUmFV5rkL/ZM7HrIARpvKcNWXA2y2UcRMIbRIHpU3G640
zqnhR57OSz1xGi1gueg8oW4FJXtqKeSUXv8fY5oug5K4n/r9Jb/AACYiQVJWOmj0
XZANqgLlBSBTBkZYZuCBhk5NXimFlIcfUJoRKpph1SoGEmIjSs3UKsVbHcHUhUh2
DlK6zlCcDLySW3kmXaME2jcloFNj/wPUi9kgEzQI7E6aWkuCl1moDbrwsfHJNQ4C
MaJ5D4NZ36MhSPX/oUw4UgZcPVaXy86jDSxA9truGldS6c7+y1VXh+ouO2S7ziU1
ZUPw+mL5puVVt4eIjAd+jLsiy1J7FLpYgWpQOrJlQ08pooOpYo3h7eJRR6m3ca/O
P6Vj9cDO9QkJuMdtpfXd7iudA5uYHVfg+++MXHm6UD9VATqIG8f/7/9mJRBE/7nP
F/JkZjeB48WMLDHloF9iL2aQJO2Z7S0tAhOsOl+9bdx3ITWwlcZbxlS/BW37/M0b
GjEt/ZICJDB7X7b+DYjx19bZIImoq9sCchioDmSWQIN/ZIiiU6bKuvf7qJb0l5s6
/n/j73lhORdMADusbZmfAwkT5N0C7V1J//8yS6WfXE/1H6tmcZ/yt+0e6Z1e9x9X
6OyEDXGd/zugajyiiuZTjv2UiCo7whtsJyaCqQNLqi9CHe5dnB7AbGbKWl43R1hA
9D1cZzeJZw/QTnapGCUIoWLzFA4N7BFy9YFpn4yiUl8ax+wjeGCqrxFASUfEUUIQ
CffbXquERnQf8LZtuRk0Of7Gnp0c+nIKt3AGy0kwEP/jQdqZygHGEHhNBxE2GEPj
gNZ6KjCU2/bQRLcVIaY7M6NdCy/QblpTyrvz8mrtkzcWpM3mQBJlwzDIlXtFpjTY
SxJtBH4pXU7axxVE1CJ5JTCqgZq7+VWotod5dNIrvln4EXc3TGjEvZhxNxaomdTJ
amxaeGOsVV+q+gHNq0noxn3eXhJYL2cXmX0xX+zbky3m1jER/QYGUAq2lLwN0/mX
cWnDPKmc0BADr1H9oo/Gkhu7ErU/nOt0gwnX6RSf6fYGzySXiQAl+m77d1oBKWHg
TrEVVqzbC9HR9+EuR8PEZCTRVxHqGMoxlqvCp2WDnlAYMOoO+dDrvRAU8bKYq8t4
hj/eH13ffDGA7dmZ/naXewGZYQd5IO9ZULVq6+xbaFgIj2R3oBTj7VGN4L0J+1Cl
DA4bZuR85QUvjfgBveSjLjbz8CY6tB324vDcHg3fusBONMmbrsMWY1QO6sdxn3L4
BThyFBi0hrXLXxh8+VXdJiZ26HaJRmOv5FQ/E1jS0H8EXkdC2RYuHUuMG+fOS1uR
Qh0KHUyerevGyXSONYtxukTPPW2yudjKMxgwbpdNfurHx9hIoi5H790z0mRKilGp
r1hs1wA1sMIsJGx4s+MyktHxAoMEpmfj/w7W+wSYDnWL5lICkBdC/uMLBmJgHvVB
YZxgV9KKC4nuJzGs/xEGZPkj4szkNX8sNBFkZZp2mSLZGbq16BBbkR7dh9onVBVY
X/1/Y/NRiK4hVrqRE1QxFgg5eqbmk9LJSdELgTYI7/Bi4M1CVdf8nsek6/2JnlDH
q3XS38U5MDPvpwITtp6Iv5gr4lNi+8UCyxrrKktr8Ono41LOx2rtDoSYi+0ok3da
5H940z1sCnJJtkocU3TuUQKIfaNzWaXfhvaDyXrQ6I7WwhBGB/JBeYIdBAbSdfX4
o3PV24fPj0TI/u9xcY2i3M58woVRaCk7onO1Or02JNHQwzipBFMJf2pQKCg1qSa0
m8JjV9dNGrRPMYLJAbjqIL822rMu2TEcCLD+f0dsWFbqtrY03KcxTQsmpd8MCwEq
kR9Y7hYDOK9gg9C/+4JSf3ia2hW6gXfyrXnxQV20AfYpVtq4ss/4a5FR4ypA5Zu1
m4Y2QlfQm4EH3pJs4WccAnfpavWfw1LpHZuvn5RPDVTDcCA6835ip3bROoS9M209
bcvSW3jbNBsuXUGJPVf6pkWs8OM70/xuy0UBfUYlXyBUwxACJa1IuP87u8Puqf5M
gpWs7BUc4qOTBAjfg1oW309z8F4/oJTLPgYLqLogdTiasKJsM+Gi4NmoMdo71on9
8PPSe5jZBWgvC48/jC7LbMrZsGGhf4JOSsPf3Kaulp2X9uEhK5yGaWSlHTMoIkI9
cHr5eBI/e8gBGkJBDXee56gQgR+gdGgUR4qVzkSDlS1epMs19w2PgICO9fBQ2AWf
upRioVzya6oi1san/GRNFk4O7d0b4ulvK/XfpItOWLaXCEk0SucR5sq823cOUKsU
CJNGa9JaBTbudXIzBo2tfg1ksfzXByBY40rEMwAjU/Vjq6+kl+8ntJEdyMvySyKk
VNzG9Utxqzcwp78UXJ1fXFkvBKg7fhr8BOxlVx7+u+JQKxZqynCTA8kcgpQFTOkO
Oxtf3MWpIfhTo3e4JbDkcMSgDHilox+yuru8FmTW01jRgxeQh89J2ZBaHwdiP04T
yPpI1OJkM7PTa+5z7zIPP97+/7c5oyXCJ3D+K/RXNTCqGjEJnht90MNyzUXFvmOK
mj+Xm9lnr6nS0sQRTXdI6y9KjEX8UawFlbYR/JJYR3BOy2EomHYwaocWjQ+R8yJ+
2+n9+ZKsskSDV5ruTP+Ot4kbrsMSHoibeJiriXMcKnDxKwxybFS5JzUHEQOzxmaP
r6unryAH0MtadO5f3kaL2duhaEAmGPJMsvPQ6TOEbzMFagC0eGP7ddKs+rbi2cR7
PADxIUTl9j9uoBK75jQ8973fqfCLL+nNPe6ozatzQQeQTcvcn0i1zNTBBD/71+U9
hd81GzsY7z4YOHkqsZZB5Fo18hdLD61nU78rJwacyMQwoRtl06kHSSZ2Jg248SQF
uLOpNBroulEt2oHEEHEdfcPtiuuln3rYXbdgVCDwvf36hfA/NR8BfvjcCX+xP6fO
sf2QiiNKXVUE3zi35RVNlyBGMgAu1b+LBj9H3WGSS/hAd/Lk4+B33IOxI4/A7ZsT
NWNZm6I8kPWJDYAGymzb07W9H9w7t90Uy+rmvmtS9OOsSKLG8s0Uhe8IN4qfdVup
9HbkajoBY3PdUqKVqjWyG/OLCwwMq6sTaqaRueabj1lOqo+El2vb3J7bHlczReqy
ueElO8ymy2ktVb6a0BIQ7o0Ik5fchr6JMhNaEJpufz2BZUgUvDh91Q3lvTYlV2vN
/BZgrHzd1PoyPcBSAx97MUpA+0WTKrbXrfuzkAhEc+01PEjerMWA0/x7Rm7w2rkn
CVH2iLXknjXlBh9mT/xBkDUEmRa4VOQ1TT0Ma0Hu1Cl8af5Sa7qBScSmdH30sQBS
2sX18UTTQtpHUM0rotPVYbghvNIYNXt/fPfOqLI/aImcDUCUK1EEX9i3nvxwrEGz
6FYNQzLpoezVpjD6jViirl2hITYQN4YBkZyRBL4rZTaFkOERVZEdGq9KS3O797mz
nyv8sRv2GMeuT+pmr21XFQYRzkfpxB8Z0mVu3ZTWmKrDE5oaXXx+w05fDQRjCpIf
98v08kOYWTN0w9V+K1gUQIM2eTDy4IS7Jg9Pibm9rQ2558OH0SL+KSABfg4eF3OK
ahWuKgjM/0cvlnqckALuBpi920WsIR48mHUxPeh32T49E9MF105Uc7/Arf2R/GjR
vj71aECB3U7+cTHQLboitqYJdN7Dsc57b9Pm22Ff6bO0gPeNlTN0D6zSx2TZAXuF
5R/1h+Xs3BoStxGEYgA4Qku6+99ogozlnFClqYwT2RAF7yOQ1rPmnVNUVmJcSPPB
WQbLC8hELh2UXIHS1fpacMN/BTeOn9e6s1gp4LiPdSMbpIfAt54PMoGP5lyYV8XA
OUlhCZ5iF2zlCm1gYfG7M8OWFCsjKQGGxAheSSGCB8AC2JrA+oWAc33C0luQeDT2
nQCOwFUtZx3QpYp5e5+FrtHdLDLyWvFjRyciy17nFyYoDMgq67iKooxkm10fz65R
C43h2zq2APSLAluzQaeunNiMdMpwNCPRfgz2iELchEmfYbDy9+ndXBb2TwXy4aNR
NTNdXkag4uJSVDNxBaNCAi/8LGhAftgfNUAjWPV9j70ggfr1uCydfDlYJe7p5WIF
LUFPYYkTUIUFMLhsuMElufwrhejPb4q/O6HQDGdZ9FFe2UZ4hCJo3+3vWY8Mr4PK
h7yb+RtKfJ31aUp6RAulsmoMsiD+c92UaW8K/NxYQg0DsNDyzw8hstbNHmhux/bg
uRGuPscb7VHxmhbenaBaX3il8u3mBwNEM35TdAQ4fxiHnV/mUZCkiyMsDo77OCWF
gBOyEhsuQckgbc4uYi+zxDKE5Hb+SyHaxrGByuToilBv4wOALLDxWfg4DulTD2qR
WEHsPVjQ73EQp8jFhVjbL4oni7Xs+ukEVsvfpmuPZeZ2Ce/eJpD/RNeNZ8l2xU1Y
4Lyoc58oQeINhvWgYKx7rOU5IJSNMCk+wvSnSLBGWoDfsTtizEFainYSEVecmrZq
fTFUXIyWvLlHttSW3azyQNhaZlZbrTtnEDKxLIHJ3m7eJ7KsooI+hRiVeA8jphKX
21tph8UCXsaFsZHA6L0UIq7h7vt/GqsFx1CZp/+eOEFKdWsAxoN64hTTbkPBzlhC
2I4iaaQok8v+VfduBihwRljJST3gzaTcz9X9T6gv06xFNLQFRiTpvnhFkWl42HSj
Tb5wG367bocJT2/P1SSn+0uNSs04kWVnJZOkbXr6UrqY+bsRNb85uJjnuOMKl1PO
wjo2RhfvaNsE0EV3FDIW3C9OnT0J1duPVanoL9B5EIxNDuiMzyfakQnawHYs7ehl
kO/uxfBJlGn5Wx/A7X6gu3lr54a7EZhqrIfmix+xfXm+OS0C1Ho+Me1Oi7x2SM8d
ptDGlxs+Xmz427ys34G7LOk3EBktELz4Qx9xEjfCEOo1DD8aS8btqiJ//ct6I96i
Q/OD1U73aAlA5LjX2X8myoDDC+gRkg82Txgn9TKWy83ZSyY3h1CrIwa+Btshlp27
wk4Y8pODmPzADZ0w1UqHwoaxL12fu+wwBGqj0e/ez700vsxXspZ11rOarAcMD8JQ
jbTHQz5LQc/qd4HIEYk7fzOykB0MeGc2oGxAyzVo14qPucDb3ay3wZfG4ockjcoJ
kHXzEkgu6LkEdxUPFagpodbgeefD70zEtEzjHGaLESVdYV45f0KH2t32/QsAzJfd
ovmQi0U7Be/Q2QF/+EJBiNslDb5adsPlqWKHT2kKG/JS0zMcM0mAsN4vIpxiqgJX
lUn/qrH1WLdFfIrwV4h5VQ1IyXYzpdC0n/saUyjc5RXUnk0P5g2DVQ8WAOT/K7kq
eI3Xf54xpDzJJTwqnbHWtFEyFb9XkDGooaNYckt9kzINf6iqiDZrPQ/ARCEoiyqm
vXhJeceJ2TDdZ95vT7DYmpb1PkJ1sEkvlRiW1g8/Y8dedLpn8MDaeOTmxXlpL41a
BB3ALr6zHwCEmcoErYA0ziAGl3DzEC3s/nvuJqbzkBF4tZKn6dy1Yb0Bm5kDJTid
F2+hKTjvxijkBX/gFvvSL2vfyYjhm6outGcG7cb2iZlPrvkuOFTBiiBSG5UPZWe/
BBZsxHbvzT/OQKjb1xzvFPMkyLeqFe/H8L5e+Rx7TaO4wTgVyvS3caEd2UeLrRuX
z65HCH6ZwMG/so0FCd9Oz2HfceG+o1RDEdbwTZwtNU26vkkZVT/FyLWJBg53ZMFD
3Elin5nmlOnxMBG7hy600PEpPoc/90fijiytXY2FpFtmbRdS+mTrBLZDq2gJUT+k
jVwDuDN2+9WEASpoJ+94BHwVRTPVBSD8nrPFEV4FZP57PS51YM3kpQBr8TJT8fNb
2HHBOLFz/bWdi4dgeAcGsocyjPbcU5MIjDI0naGFCNlv62VpPjP9xiqE7IhVL514
ei1gB9rM9iEALLuZEbai1Gxlzp9BgRZKHYx1RMpgvwvDLPTkxxCI4ygkw2osTkWa
ofegM8FwZ4jcw+VGSKMzkOInePe9cGvgYEy5vRaPvhPloeF6qib9WMtcbRrpoEzh
X1/3MbuzWOAvz5cPMYaDZVtgjwoNgeaB35agDse+Tks1pirXCK5cvDctM5K5e+xi
r0Nm0R1+CpWKw22hA41oWFIjO78I/iSpzdW5dk2vbOOYsy6sHrlgAZ6EzKBKG8Ul
3TGYGCQGB/jZUd9C5BPJZfP3fuDUv6tqnQ7NhUqNhPy70eyrvrLURDM7wKpu+Sjv
I+MRNVpNaXDLqXjiRjAsMTEr40sFtb41z+igTbl64b/NCWxVGqHaeQOv14xbxBBW
xuj5nxMiGA+AHgyT2TC2UxYjIbYrgPX+GP54jNG4Qibxk+65k0FrDhsxC5sxcsN6
aJ8bI2R3EHT9bO2Rt7kZGPO8J3KB0256FW8lqnSq+7VJT+7Je7vWHYmjB5pj5Ym7
h8EFdk/qWUVYiy2Qa55Gtbfi8exeakqiafG/TrOJ7noJXfuhgWMDXJp9tVVUusGJ
rH+WU1YBf+z7jfsF0BNd+tNRUuQrAn2CxMqpiK4OvLLbAoAVFYXhxtjo5eDHWNtF
Is2XfmGRgrKHxlJibX/eG0ZNqMtucJn4nio/8torLohbzeW0LfIDqitJhByTD94S
oTa9KfHot8WrXFCVKQJ+BB+/xNYeE+KZre2wn+MZK3OuEjp6hmexwK78Cjzr3mSt
nh4VXcINRoRISu4vTiL09UQV5x4MVZa7793FmtXltsls0Qz9XF+qZ0gcxoHljhSk
QdTuLJtM1s/jyRewl3trReUb2paNtElQdMBbIO2lHWeynt6K9szhgq+qsIycmRow
VdTbo+zOb0xqF/4K8uTUd+KfNw191hbUcu4TN+3f+LX1A6/KYpm6LAvzY9I71uRm
7rPbxkgqHKRnciRNGvKu82Csy9DGFAGEXqNaw1aBoRzLRQZ2biLVTK62yRgtwguN
Pp4N8QVF+cgH7Lu/LGti8BxnURvE57jNhzytb5J4pYZJdZ8uqOSJe6QPW9kp7tA5
wlwF7ajEQ4a4DMgZXyVxf49JrPbDwcJQ+DbARUo4VAgZ8xLZYbuVrAPTrH+2a6UZ
rwWQu0CW6k6oYLtr0q995CCwDnZgZKud+5OQDtXdxwN10RLYcLRbmPFddFNJsjLH
vl2iOE2h5MHtmeXaoJnBblp+17WKrgJhx/2erWqJlIcKVWm2ct5JsA5xP+JKOkTb
6G74YNlIRbb7upF7MPxfSa0Uph5Rv77piTj+0jPmAR8Ba3tKvec1X2k5UzZW1St2
p7ZpdQ6FhqJOn9EjwMfSt8dgV8AYSYinjqhAuAjs0tYE2/0ejYPPcR6Ip6hdXBti
y1eZUYLtZPe1S+JfZ08T9i1e8duuEyaQkx1PEc5nEYnc7aKnnEDdVjjaOdBkX/rg
bvJDe4kGURa2cUWSZwDAhvWztSeOR9heOHCMh8adMr+bv/azhc5kJ15W5/RtI1Ja
9fbkh/tEsvYnKNux6DUfXdWZqnIwbXSusNZzZp/1JER5PW1x8khh6QMHKdgJZlqC
9mQLcCd9z2LNYa5OdMN2UHFqstN7P2j/mMA1Uf6dxSsY+Is5r+ya1Ng5aiJ4jKrb
+egZR3cuGAPG/IwPBBrvJn6qsoP3xKsMIhbOUhEnXfkp5nu9AX593IoPVANTq1TR
tULs+7uw5tDaZh4ekX2cnDdEyNJnDcI6ZfdH3FiBgJUUEvsm6wca3eLNqgRO1QiN
EPuraW7KhDDMbfqFGUEp4kiLXios3/OWum75ofJbF7gXEaoi1hMnXzXSi7gPuLW+
wcE82n0yAupmlcQJMJdDC9Jq+LUOmCgJCw1HUJG3AD7/ggHwQAJPVrRhBK14Js9k
QCitlG8fkiYqUnXCBgEiXfzc8AKFq0HvOoJiv5hUy6wwSIZatOizZsC4BxBcyBF1
NgUUnMv6FUvcX28KSAAN+GknkjMRSyorxm4ffBN2zjQfLUWiDGwmSXIOOx5YGGxN
DvhC1QBQFlAR5Dte45nUYWuk2otTGp4/UDVFuYWp6fQ1Nnt4a1B6FQFhnunrPwE/
UH2AG5T13dHFr9XSIJXAlThSlljPHz1mRxYqOaXXOV07t4pfiaUq23meEgOpDMU7
rMknTFy5h0iCc3/1wEpmqtLwDmesKmnjaQmS52ngr3K05ewQv/Eb19OgJvCVY8Rn
s189FqGq4b7o4KUDUhY2ugdHppbL3OC6gAVa9tkqnVWzJHkwPRVOfMBUk8MlA4cc
njn+Te5HUsO88xa+uD+wzx28SwVSUmqFBBWPAcwClAq4Sqiqq+Wkfad8PMDpXvoJ
s0DsGrM8qNQc0hGTfvEW3cjYduIAloyhHWoAyphnbmJ/sUvy1Drt8BAueZ7huZZL
it/6GLQQoYgQjkKZi/sXjfcpHvBVzwzbg+Zt/5M5vcXFx9NUPSozMwgSCeDo6DtG
WtkV4kyrW8mMHYDhcacLST8tCw1OwgUE+pMgtMutP49rGOdfJHJ7vLlMxMFmBrlI
IzdoBVPbeCsEwnWmK83AKK7X//HjPBH/UpEI8ZClLlRk7EUowQWxRkEGxEKLL5Oo
V0+ix+AS+VVOzOQ4WaKNg6dkA77Wt+RYc2RmssJkTx/YKICsOHSaGvFmFjBHquMl
IZyuFJbIltfpejD9D7K2q9DEW3SFfa7tm4bOcT/15vgnhcPEjep/J62ILtSXIzmr
qsamrbHkDwz3MiOswLb2EPrEgCaERIHiHlgUfLOLI7AgbHB0UjPi+Yv+1Uxq2QUf
Gvr190O3GzYHIg8R/RSkvQ2TmFV0g+LktUlmwDugrptGqHd94iVdckgKs5L2JBug
TsZ+idugN/vwOog7eb+JbAH0VR6T1GJnjMB2bloY6fWpKhsY2yb2+/4gROYA9Qup
0U9gslIwq9LFC4TQCi8QG+26IxChwWqbUXXSjOp4e/VlhLL3bk4IZtGQQT+qIFMZ
yqHech6TndVZVmxk0VLcAkFQGFnyS9i8XvgD5LZoZu9eIhyUYQwZF03mATXP3dJC
+fukk6sGbvz84f5XrStYkhW7e/b9tjELos9vbysw0HOmRuG+ETwQCPJwZGaTk4R4
BUnjC/TIxWxwAV03xlzhGyvT+TWEIQD0VvrW66+fNv7MlCzwhVgV3rJOdsm3v8Uc
r2XD6EcvEo9yYgbUSXhpSA0/u/1hlqWFDHMloCZVfLj21uZXDAw9q9IAZKsRRTP1
r8IUk049kll7yLpfdeyEgS3ox+39Mt3y5DNOgzk0G11XXKg2rCAtVko5AySfJUrz
B0jtXGX9xGxji2nYdU5jV3ijPliTVkVBzSpEFVmMAbe/JHH2N08z1V2g5/TiZrlg
jaVoKfrRgEEqz0p1O+7aWKZ08KHBtSEWSO50V3Od4GGcSWLvqqw+nZUmN6WcZPrV
0NSWE7nrIlt7UPMmSUzT9pjxTW7YJmc2uHTbWkvkxHTkWks8cGD0+522bKae3mB5
GM+bdmgYpoKzSH8fzcufAzX569KnDGws9VIRf6vx3A05SBq3UwZnbECwYMH4woGB
rDGAamTXDy800/ORSEqFzcg5ZaFtMte9Aw2SA2Gnpq+tDp//KncJnsPzZqZymUFY
k0dJklM+UOysPjjT24+AM+OA3skg4ort/ncKtvcOt2Cmf0AhK0hWjITWvrgPXBKi
sAh4VJ5b5i4rWmbfxNHhf5EkICkHLlJdyDVAQ5df9KVSroF7G/S5ZL2djyVmiAoO
GKvKRs2BX+nhBRob0loQPguZf3TwQ/PpA045BlS0aFEIv1pYd7uz6hh43EgtmRge
ZSFhX7cz2MDAU6oykqUqBuave1CgOFdCGVAe8amsIi0lbB6Oe2dotNuKwrFKxXIO
reza3j5WQHI6kjNY0ng/E3fe/bJGZy93fUXj8B0S0SxZBQePIABk3Emjs/ok20tN
7dD5JiwQMLp8bpbwrzPbMWbFxioKTbWl2Tv3zc1ASyHbf4zSsrxzgg/CS7y7vVQ9
kuzC5Ddp1P34V6PpypKtO3F37bg5/nPKw6XElEHhnzgSSeeARXYelitZHwzqyqmx
NBkQomKzOHoGw4RL2W4WHDAyxxKzEw5wUojeuKCeMafHUlk627PSVAD2Ix80R+Tr
Nh3Eb/12xT7KAHnhh6wTKUGcbZKpRtwKEpn9mS0pGg6jkBj2eIA3opHIhJnMMIJH
kXT54SqhXcO/FNg3+djc9dMyBrZsY40jSWxBjpEFbxiK5C8SPhKsjNtAtbxJeJd/
MHdgwFUN4+BvLQoYPABZFAi94YfRAxQnkbPEjpALSSghdKuIyhcCajQ3iY548/xt
8ciDkoNmyNw5hB6rLsZhvyw67LA8PQ8QpUW8y83L4uDMZzZg3Y028t8l2OlDo6cN
G5R9bSGwvlqxcXq6OnOJ8NXcFZhBirVK7Z+iF5i2PHVxKMtVhwoEm9ergjvTEvgf
tNUHz0S6QrI6J1XpDTWF0i0imaM9nQQtl1DTbwrt/0Gz1QyTHsVpJqC5IlTBDKD6
109V/s9qpdWj0O8K93ihnMsb/YCtxBBGz3vKx6IvG7rrClG+RENuyxloKO0ug47w
e4ev71To9M/aJ8SSYAiksCcgkZxaXc46QBXEWKWsvC/jFpcZ7dR35O4Jtlud8qD4
vt1T/Vdt/nEXTEnrJdVx7kJu3b2TYBrH+TeV+I7IrhcdphfJ4FlY6Y2gIP9jXZUu
mlND2Q+KVBfzNzKPyVm1OLHJy5vf30tv4SqrFdbZJeLvTKAaI/TFx3N49DerZWe0
OA6clYTieE83HBoYSrJs4v/2p5ZYh/8nOpTM8D8nB8Xobhg+MmbU4uBh5nYPY3hG
RB7bmMpZ/Wz9ySiwPRmhPdCwByfgL/0YHo7fpDT45qufZogOvB/HNshLSZGKUMeP
7bojCWOAdkuk9lWSl+m4kHSt5KlVFT1p2JokQc8dbeACecK0w21jtP3pZkaRAddd
gN4S27JlQ9hS/muyMfzO1S7MNDzpEqio7hmT05+XzTvldj8sCfb1ObeFTg+AIHR1
+ktVotw+ZYp0ODYVeXG4CHFuXpz5+m1xAk40msW6qM5IprROdem4ZDABRp+hLpqw
J8dHYB6izLjuttnoNR/0h8ZsxJVEWaxEkd3MDm/zZz4YJ/oCKO/mINbF/oqZwttF
FohuoApqWtzltUPbI0CaOqVSxCWBDo9x7FA4N2oB6CTs9G4LcX89P0q56x/YeBV2
Le+pPyPxJo6lSK/NnM74q8QgwUJpOdaVf1r/XI+lPqyoSaNLM5VmJitUAI75H8vt
VhD0MHf3MnyMDLjaKBDhPbd7a7z3qXmu6Y1Lctm1Oydy0jlg5smpjO55kyrhDKEq
7pAs3InV3gM3x0rvt8iS7+O8EJgui4ZoVTd+WBFF3foPp3rNj7CYHaYMF7eSq0dI
2O/fiszJ9DCBW98ir0eQrtkRq82uOgKKgaDSy9OAgK+gUcgsEChfiHNtBfrB2WQS
WbhszZlmhEgsWBbkDOBqOhUD7KF+SWrtSugDRonn1bmsrSf/S7ziTLzIfy1SdeHC
w2PTOVaE72baLWYx+xud9X4NpohtssNbbjJZm6bRlObN2KhNfNWCzvG7Xt92Zfwi
zE3dSLTNfGYbW5EKe8rpmIOlg8WK5ZqNSwJpAsVd8ejctb9q1b4Lzse/+W2+DU31
1NSriwDd0+Q1f9vvuO0wLsqROl/iANcFifASZes4ceYw8E0myxJ3zeah8Xr3iSGc
Px1jfkZPpYYEZ35fUE+r2+nRkV+0r7vab/ylERsnj2xY6lu58DTr7JvvmSED92cU
TOzuKCCZBx/aeK+m8jUTMJTmrfMNkj1w1u8boDx6xlaptLlu/lB6R0urqZegfklE
IfX7xVTC6lBvuaAv44mYQh3rvuhzqqy0I8glyTSrgxogsO/F/IaP2/43m/diJa2Y
IkHt1F9W5CR1W3hdlPjiu9K3ONAtViUJShCSp1OhbrUGBZzg7IqfMHZT3+5tGuPk
untZFs5OHlrNxHNknDGatEEO3ODkh/8yxaUo/dATDFy8+KYA2HLWtxRLvkHNTRxW
huzs1doulhGbEwSKbOT+UuLTAVGSVPAR0SjxBjVI2GutDc7DQp1uVVegaI7m9MZM
hmhUOmjuv/GxAXj3QauMpmHLUwXdisEMEJ+xlvcywA+Q+mE7Z3rE8PkEpESUAL/U
XlBpTDeRE1IEUOzIOM0XpNZntjDNoPmvBYiEG3ghpXZBg3SkdhGgcBRtxWUZjWdC
XVPob9au0NfAaLysX6hio6m3zZu0HkUNmS0FhTdhbDOGvxEmWSqlUAihyOdx0SQI
bXRG8gyHm7XCbdFZe1+2WOwGJv+iFHqQy4x3H9nR/npKwB/wAyNS07VlidbdKC/t
3m/csdGd21H2pY+WaUse1r4SQgokGU2y/FvUIFolf9C0tdAH9B0gZIe7CNjRNrqk
2oBpe988DgvkJ5VPCQtzXCceJqMJNHBBdolCpyYm5+sI+5vRYHh+ambrAsa6HIwM
jMXiENyyTyF2mTva4KmSQ3XiCDYOZnIgtOVIUGMY7fRctwD33yLLWj/NMrTIQQzd
HaPcaGuiPOXiGWZTv3nmy69U60Mnt2F0UST/y5tnlVSDlBFo4r4cfHRtDCop8cYQ
TdeJKVAjjPWGWVETWP7k5NTDV08tN1hRTdRvkD6/141PUQflhkHfxEBHiYcpQrew
0tYl112IB70O2mOXKVAvxrgUr7fs2JMK+ItiIhv8f0zuqt28xTZIxo0Fs+f3wD1d
Hdk6ymVk9ocjaNR/C6pwqEQbJCST0NIfEVOAVv927tbpwBhIRsucogVZ97ctH2Io
oi4MSbOejzQFRwZ3Ez8ObsIfeEqylN7mSGtr/GLFfRicobgrgCPU+sG9yeUUMibT
vq8KLybg6AEhKpdGx7IYOR8IlPenhbAG1WLTjHaFhVvwpY0uCAGckvHEfRa4SzGc
nBsojFXGv8nMS/4SwZNn9HP66kVRRvW8Mk2WG5AlIQnehRqgKpLi/NW1Jh3QE5Br
W5dRzlh8SAyd0zW/kOQf6w/jgnh9BAUBhop75wiCf1oVizgNX29RYDWApJmVy3J1
Bt8WsWNjy0QfZYa5oj/R+muUDo8rLfx0axva3NFJ3E/YVOkl+Znk+IaSrwaQUPl2
DJECP0SLF/0klqaU+HYgltBfGKk5IkSa4ObZmzZRNo958YmJ6DiiYBlr4ePcBW0a
ZlwcWjmWpxcdJimcShEvKCDC6Zk7WdYulNWMIVYKHFWoBsMQvkpqmRRfErUpBqQi
4d3g8EmQL46aBVRfi8QdFFsJgvLFEMZZaBLcr+qB6whiXboRsXRQbJymPgmynwl/
TcAQaNgDbJgmbeWHH+xUwzvn/bT2Rjx5yoaqFybMftFZ82e2UckQTHR7Ee4cTjOD
evcPnmYNYuA+npBJI6xxIDV85wSh33wqx2GXE60psRtKTDrF/Zu/DFOqqECDdt+U
k2PuCgQ9T51jn/4ha4Q7xmPrZEBbSEk61pu3k8KYWcU1Z3UldpOmfrB2z5fWB6by
qZ0y+pJBk22r+mMLMYxFcVYkSS9or1cTmiIxWDF8kryfn1ru+UbkV4M6R//499fg
O9yKGjgTiGH35Hg2/JynGlEx7+WzwtyZL1Bjp0rLjmhw5d81P6tpV2FdflhXENm8
FBtPuI14J9ycYLmchHTW2VSqt1yGsfhRO3AUTb1lrnz20ePxVqrS2j8UOl1TVVMO
aHs2PfZanlaC7DKAs3mlxnb0de1FGqtlbPRpJRjPgqtBVWpQPJTt/OeqFKNsqvKU
O4/i5ngItcVYOAA/oyiJVGWKxbQFVqoTwFUIVtZJnau3ew30k0GB93XTkL6Snrky
GhFmbJZQJRYep1WR+PPbReBkwjhjDE4D3QRxeFfT8mUBfdgEXm6pKBjXOqAthzHH
QPrEpyOGpx1B080HW3WhBk77zh3d3jBXr/AsyqaBTJd2H/gwJJUaU5TiF5+ZCVpF
tg1CFIuTe3KrSoIRWFtuzGEbwL9lmA6Av2j+vlon8VxiV9vBbPUFPDHd8kqQfbNh
9nH9YKc0noSUxmM7aN05bR8Utp8G/feOtCF/4Nyvgb4jJAkuT+5mn6nEntR/Hrgo
FI3a3oHcXuYtsV9sngi702dbBBqZqC6KAcwVvElB8W9B3eNLIdSE0gELIWun/GWz
b2Cyr7c32lvmEY/K5EKZRSWZvZ92bP/7Vr5d+4TQOyIjnBoAIqMWvhjhKzro15yK
0VHf+dYM4DfFKAm4XophvjxLnHnHeVUkBxQkgGpHoYfvonS1/rEwVOUenlSzd/s4
Idazs238ys4W0GJcwWxSX/i8zvCIak6fYF3Rv9hndFP7dzXbA0o2XkzOAOfeILtN
fGRIKrsp/DJCDT3scj6BdRlRJ6+BxH3zuZKbhCiy9iqIj4fASZVvemMCENld4dS5
D5rUwRgGZEEih/0CzPDf9PwDBq2kJiv4o9PoRyFZa0uIfDsG3rPSFvFeaf8VLNXn
4REZrnPeMtgRa/ZJVoDmGhFFzoSvjJd6OSOMTv+def8uz8aHOAAW0UPdP1p6kFlB
OKRKLBHr105dHbaOEc3ttn8z5ssujPxvKzw/lHkbPeWMzN94EprX+diWfGYXLyiW
ihl1LaOkJiFlMFZL8QV5se9sZT4QrCREApA3jXjIK0/nd0qXPrZX1B3x+FVpF5Dg
IgXcewsBEN5ji/t3gijUiisO0iHY/q/rvTPyDo9Qxc9bncwXEjPYzZ/QG5ozwVSi
52WaxApevirMP7sksbZf3uyw9xK5Jens5PVWGFt2juq+T3Yw/NlpaYL34GX8pqlk
6zu70t393T8nsqBBsvStXDzubcRVM8AIY1WOzC1zW9ajUEl3YecDHtxSxsdn3aia
Ibc0x+53IcDeer7MjlOZz/hrxKTUhOv72BNg0OIYwiW/J9nfo+4VVuZ52gLx1/Jm
RZhCNbm2yRFFperb8MzcXM/5sjpkPb81KF6PbJaLW1NGbyV8oQ73LBm4kryFgFiQ
JFqUoao9E4g+S6vz5do3/yEEhEdpcDpcvNr8PNAlLYaEUoV99TLeFF7ZoQ2+lsJN
qk2C20ECbT2yVqKV6B26cWhCOaK7aDlaOXw0eYCRauh5mYf1fFyIU2NMpktKg0YZ
Z/LB7NDmJ4dogQn4vnqVNMxWTbFO/53d1JtzcCRVUrm0HRtevMtBb6xSKUtd8uH9
4+szSivs0jEYuqRML5b6eOFpmL/y8Hxo9Vhd3PQHp6CjRbxO9jM1n6z022BIhVnu
OUpN9bVt10gQxAdOh+4SJXlk0Jb7IwzJWzjbCVhpGoP2jxfTVBL9n3FTrwTNIUFN
3i/tmlcd6x6KvSyw5BB96kM/PTPPX8VFXvCa4zesyt2q6Nd/MMiLGvl+Eqc9GmNG
uDr5Gn3U5YUuCjtwKfSaz1SfKXrrCwZDGIdWmo4rQ6+KT7mn+xRFmrMPucYVDgJ3
/uRnvYUE0InGhjZkg9EuhrkzRVjG1TrKcHoVjGzUVlEccf6Y9D/b1YhRIId00SW/
1ecHi9VcTZnMClm6aEYh1h0EdQX+UMKY/4wFZp2MemPV0efG+w+Ll80QKnH/u7Ar
Hv68o428cWAsWCf1dUQ4XWGHrLyO+xfIq9rDsKrV2XC7Nho4lVdu9izOlNkDiA8a
lHFiXYJbMXeEGqbnLH56W7OfK19a7msGX2B+F5BxCrKH2xOr6osEmFCD2fidCydk
4NgsZUrro04Rf1Eo03FZS/cknnjtYd1Ml5vP4xWT4aZCt5jObij3LD8U3ghlJ/65
uzaybWfP7Cn8oBG2x7CZ4YJc/vEEu0fQIk1bqaAC31mM1MTxDODk4g9AJDyEqX/8
ij1hsqYNej83Mk0s4h/dqTnXWsDe3igjDBObMPX2GyYVoSFsvwmyvwMZ7yRn4Vqj
/l+zs/Y5+F2RdtICt37muoC5WX+SNSTw6UD/fS3878Q8h5RTbJcdigZsbFG6ZGAU
rlZS7dvWgy/3HlB/xgjKaHQT9RBE5GXHxl+/lvF/f5OaXnarG/4Xcr5va2IeNhgj
fPMUGdKgLACho0dHa+lMQUsjKejYnD/9LBgghhE+bX6HES56rxcOmJmnoEsEvEWo
EyBrVezuV/3WKR7VQN9cjp6s/cVzcoiCTbbtnLPnm0F7uta0RvGDUd9B1GHSXGDO
c586oPQvKyIHEYV8WWkvwQvLEYsgfW/JkgoGFukGfAebkqs6/iu/lqwTKAW9Mzj0
CDukcV56wb8MPbYiYB0GSSBZWw3hgHMQN1p0P95HxPwqdjH5JQu2fOlSZw+6+xPT
fgmyhY1Pf/nwsZ/7q0PrKHhJFOtZ3YsSK1qAg9Xy9JvEQugIu9IBuaX/KW24LNXQ
MHhI9HrBoHgvAAxNI5dpylR3P24F+cOpyn+zY8XmUr/xPbgnRoB1ni8BP/KuTv4L
4jRpG+sBbBTK5iQgLanTDBgtp+pPqqXYozlzcXDL7OmrOJlGPCLvcBCvqiPrGhfq
GoLy56JXgxTDUDJCtuJVQzX/zcIELZxO4T0xCe7TDSNWyH9rIjX4hUXGcv1QgMQQ
5qHugj3kiZR+yyL8NO/1nzXMUSGDmIW2VUvyvBb43jyWUQGZ19KMbUFo3GSt2aFE
4Wgxl/MZzSYyXtFpQsrAXB6IKT8phG9hr6nM68ujsoWXjXmcaUILNPGgHfhkh6rX
CVyg5yT9dBSr0tSHfF7thcIbnfZ3Fq2cIe5D8qs5WT9thYfuXwzadKS3aUIcb335
gNEFIO4XtJJNq9vJ0xLYXUTx/G/GCCMr4LClyNSoPu+h405EmcbnEbPifzxLFJ+t
18c2WBtGHZYSwJ95ehZLge4986AiEn5rxE1MMZRU1jD0Meq2ZK0BK65ZUZOimWxP
xSo/77ZjYaRZtjCdODaB7kzjcLh0Af3ERtDlT8A9ZLBaG+YhsUbYH101VJdbrLZz
M1MEb8OM4KjFyjYV+/p2LtSTkWRhcYzESyQeHy8MvMiF8QgFaoHm5gkN+OXpNnbw
eW99lkfnIVHcqk12I6796Cyhbu53ZTGnYaqPNqkk6T+vrBAvYbVDKOhXgD0X8wYU
1ObqgWKGk7AkLvTLvjrZh+6nscSwFIAFijUOa3bz8cQR4aEf+oJo4NwgNwZsw26Z
Z8D0XB3adQ7q9ivCiOQBfewY1/r8/qFS+0PYOaxHxizDOUvmpXqa7Kj9spQPJY1+
syqZ1h3OBI47pDH73kFdVUSHd36bsycuOnuea6uvKNEpbMY4ABJpuPiF0LzjD3UA
MfUx6J2W87gSGLY5ho9tpaIiNeRR1TrzAPc5Jnk6k7g7KD/CqHtYY274IL5Us6VS
pOF+yUY4hf+LrbzME7u4jl5OYqun5WTbs4BxXQiKFYHjy7s0C08lLNJDRMhwikbe
V86C5kpgs5npVXM/7X63/OeqomCfUNUXkVntckhO/c0zh4BzDwI1eiQUm+rok8fU
aMBhkjT78H2ls4h4vV2BHCyO7gYK0mu4bY9d2b9PykNLXYESaPiYv59oWM/v9sOK
UF2Sue/9NVGMzdPwo+w0iDbInBC/dSHfHzAuJ+ocjrgN2ANqQRHDY7+CQRTfG1l9
9Pl/DNUWkRPTCPBM+q2kB2ZfRV5+zeO/+Yc/hsw87wh8+HHqeKV42erDRIWhMfMs
B2jbBCzS/b6Jyi9OZb5PyphVdgBsR22t4FUQKw0PoRn1tNbP5icVEwVcSqTGBER4
/jaRvs+VFrI+HkMw46xEKI+xSqaqBwgG73QDFvAMrBqXX3G84G6QMn1QpfOG4itc
4xFsVe+2IGm2XOloDI7KuFzMsYG555hPJnxNLBcRYwHreLahKfUZA0ViamNr1fZA
CaFiZuwoE8RiCBXaAamLzo+j2tp6yYUc9rnE8DiecNkgio5U289cbEHbif2CvbrU
TQ0g9bfUILXJ2Muku/f0QT7XuFmBmmnyGlubPF+Sy5eaHuVorlzGEvBsnVaQM63K
9G+Tprn0daH0I+UZTWoCnmCBN5kDDrJbszgbEoJxXYQJXI/XTDxVNn6M4mEIgscV
7XONSK9VA2ZNqRdJZFZkwbeRfSYA3hEoQssgruirEfpkdTMS7Q09K4ves7yNU4NZ
ib83zz6cFQcoZ+kXbZQs6l/pUbUhDt0I7MJjZeWibx1Lweg67A9I6o3CjnYyUwAp
OBJIOikvK3kDVSYfBKRrFopYjAJO7ERm5H0Y9rdlZAKwfMhwr3vLh2yrMke8ZsC2
36mqJUFiboqWdDbUsMSKw4XJuh2MDkSHjhEhlAnRKGbiYj9t3a0tHUXxJrdL6i4/
upM7ZWZD4RY929b06LnkuufV+M6QCY3l7NBL3oSLVt83M/0CqTaKSyOxIUlA3Glw
dnfL0NyLhzfhKblTrb5bHJV51madSZiZTjojmUKKchcmCcxZ+2xERoSJ2XmzqetF
WmHKFmgRSUpyPfL/bD1AADSGFe1hE7G6cinHQJ7J+GJRJwUP5Ijcc5Y2dry229PY
JQsGpNMA1hn3dAN2lyDtYxHPC5jBvBsPQjKcYj/oVaD7x0BVFPTVT8LOsmCiWMZO
uER0Q3gMJ1VqlK8GRhwmrp2JQC4DhGbuBSP6yvYHaR77+kitQ3UB7/JrSY6AE6WX
l+qhR5Lo59SP4QVG/qgxEpKgNSky69TTxdXyRvtbwFOg0GE3G2V26y9g9WFULkDB
8O5zgHwYSN68+4c24yn5tl5O2D5mp9ne7MBG/m+T+g99+kQC9WSOdS6kTBnqbkUo
sTlsErCc7rQInXGY9569jd25U/qXUyE8JfZ5N4/MjNUJd8Rv36bP48/XLXVWKJS8
FzRDmKpOn1xRGeTyEOBoZvwpi4KfA33QIHfr1gPu8cCz/VchhTZyC3l04QsSHou5
UvBqVDn7StzPbGqZ1/7hGMF0RCbfep/ozYMKfkQkIRPzfji+/CcUY9GZn2iKzFC5
k2rX2cChasA107WV9pc7I+TIm/PAMFx4aW7xQZss6qYLXd5gcz0TurM28bAQOlbR
qOHOeXZSbo1X6vSvYSonMi4Wy4kVyBU/xMQKa5hJlHwP85LUADVpDKOW+QcOsivy
7KMmjZMCqj3j2H+c95+rZoLJ2Gj+h9rHtRVI8C0X6jsHfaBU66ziTm3jPppYYOff
WcHAYUauUV/qKqLsE9Dy/6TJz7fRt70+KxsrUGWAQOqgyAak4SgiG9AYm7Voxf2H
nQ5YkeTLwsJBBPv/gFdSetCz7g5JbeE1J3UzZqgpvLjLv21KKkFXMrtdGSsE4rbJ
XpeW4Vd6UirBX7P9xlz3GA41K/AoxvTtjZObNzauFVLwlYWy0H6PY1hcPva/+Okd
s9mpziK2wg9+TijL0TmvYgWkjiGDAO/Y/y225QNj/qstlJqarhxcv7FkzYpTMlnA
9p7uFns/7bd2oCxwkgzQuNCDuEdN3SHfPEZMQtcSPbzQ0qLP+s9pQzXZuXojmqxL
T1EJBi3rTUKTQJrM1gheDrqAy+HzDxbqvx7f95UCuDacf9vXER+mVS1qAG/c4EgV
tqIDzNJGT8oNsGFSunZjz7kaVPfFTgcvY7s5sjmc7tuYJAsqE8MC6scHwVL4MFFt
5j7mdZNB3FFN8c3VzHxbhlztezwBT0DQLW21JANg2mCPpYNEgMisku4Pu2hvVTAJ
BTWT7KMG9ub9cakZ5w2w7Ecuvd/ZixIWQyNHrF+NHpkzJPA+SFyzbj6FojwC1CH5
WBqJE0X9+xtNShkkH0U+VcEyZ9L0bEg9Wyf9u55pbl137ACBA4Qax/X9j7abqA2R
89WsVUkdYYyWj8odNc91rTUVakIn1Mw3YYrjw5xRzyr4QZI0wpDXNh0M8zskS+0V
i6TQXVxJt5x1B7IGJuyhUH8nO5B3TDnaZjUWeL2tDsG1IT407FP0UFuTiT2FGP6I
2YS0qGwEatOoNEVlvQ3+SQgGCeUeRPetAdy73Aqvvd1xUDpKY4z7c+Wj0E0oqmul
aZsYvTGLp5Af+kTqsyHZ2P8t69OFuCvfLFHYW3QP79bcI+ldg1YVF5rQlyheBPVT
mkcOsLWWhMzTQaz5AOlbny5MSPNFrcTM74LSC3TyJQ5T3GdBi/fgPyoxSsehPS+i
Nx6ZDF+7TgMiAhoUKAiUSDUm0O56KwmwoTnaFl7bJKIy/2R0T7sCM2siLmjQ+Fki
cmrgon7vkva/uRBjPUkZ1/0rzMd97FyxGjIlBt/kDt12UFUtcTyClo8pcijXZ/p0
tcnb4e9RH9lhLdNlYV7amuyLrqJ08Vl1tB0DLRgAWWLb7sFiuxRzzMf+sMZEullU
KxynTFfjMJTvhrGz2vA5o4vOIL52XUY7tD4rQ4uKXT7o6Xirb4fCxYLLMIPfYr3k
U/L5tBwLU6LczDUHgohdhQ2hagfVy9t9BhqfOaXsKnB4QeGDhkHJ7cSnijzvlwy/
6NCOeSP8/fx78RA9lhk6V2iA5JYssTaApv3KOI2wGxFb0O5iHnxVEjVvwuZLB/dR
aK/33E9916MTbQYZdLud4Xk20XXWl18523pgZK55TEbPl1I7Lju0k+7gO8k66ifM
Y9r7pxsZ82swbAhyFVIKsyOjAUspVfwI86vn2QmMmQ+rIUp/GFRO22eGHrLMFoli
EEtaz1TrC4+psQyUn+VzfzY3szDoA/A0iyvVNZmE6gkypbByhJotjqVK4dmmmUMQ
156dJBsZYazNPw2qgTh1gbMTbtyDMaKFbG10Gl2oBFvSaAS5RK6rVkxyTWRkaE+F
dg4KQC/dMeMZf4Q32nBWcp2xGcjpmRzfccJpI+mPRVK5QqDCE8PhphwtQ2o92SGN
VTqGNXyOI3V/vga4vDU4Dy2VM+20sqHuHZskXiKxFZvKxmes8mzskDy9S7GX5fFu
xEDZVlUk2gfbhq6bFKzA3Ly0e8mMl3rzFIv0c/cNXCUdOlpj+a5mbipzlBL6wKGk
U5kuyd0xmshvUTObHQQaWil2paFhHhzPyZ1RNLr/nrTv05FABOmoHzV3ELZb2Mn+
Yma1PjoaHfKqOK7P0HOcWmYFY9G1cxWNYkG2iRDtBAY8Lcabx4m8vEAfCOg9UOdy
ZJ5V10bevs8qt6jvjxARJnvMJcFM2PKnXtcdjYWkJVrdwdahhx1IrQtpo6Rh2OBk
w5R+vHFVs2wS0dPuKXT5aSG/kBbZuAyseo93XrRSNmvyUHo6wiMicj6dbAAMYbUR
OluuDnMjM97YvgxMn6CRvXP11Rc1yQzL4xUT23cL8p86dMz/TJ+Qjc/h2yAgsFBP
F8APEe3rY6SCwXXW4+PWU3h7wo8Oul55lau97mj7glppe1AVFxfTAMBiPNz7swNS
IWQWhQIIdmtZ9+sG8aHMMQlYnvrczhjz/edM/2nmUmwNGe9rHr+9UgMz5uGykYO+
tsJui0Gt0KC2h2ytCfY4smUH0ZEQiY+P7kHAJ79QeBw8yQvwlaNYc9yR2N84WhCq
PmbLWvtu+MG3zJg2mbHmGTsSbvJciA0Aaq1e3QLUX4XVCTKn4y5pzGoY/e5eXGRd
MrWwzZY9IwNUbHopSZj+s24yPT4P5LxVFhDZag4oIBeYLErbAUtD/6h8dqLjhgfk
i3wbTIpnLV3v8z9PlzAmFIfQiIlUlC0TxTClWpYtrt6dn0JhR+OCNtkFYeklYGX6
/vdxVnsnMKLI4yiR4NhWpQ08IhaGlmiO2OCIM1nPEV5NiMR0u9FlTKWDfPG0WKdR
5RVKPPHxiDQvNlzOIjMkz3ie/x6iZWp3G4xOHK3RFZjIls7oMopBYmKyqMsMzN6M
mXmSVHJ/w7rQgalY7LFi1/8v3xd0Zg9CATq+e4fRnP3ZToFNCORH6QJodCPGt5EJ
78TN/MXVcrpRaKeEmdlbyoI1ottYvfzHmTYTjVmTD6WFHcJc6FlN8HbQsW3X22o7
C8N2u+z89tdkGQA0/3oKhZ5xpsHAgTPOfgVQc0/kctXdGAmHF0wwaP+Du3AewAAt
BWYPytjjS+I5UmwzowhgWHJ8uMZ7L2DLjwO1xgMw0L1yKWn7jnvP1zRk8+8kQvQG
AsUj6U4cACqwSvEXW431GstwKUJZGeIHVC8Q7tU4MgRQz/HD6dSIibrAb+UHCe1S
bj1hceQEOuNAlAau9tFojcFUag+J7iuqQlDfpQuV6vaDUrF6yjDnZB9zSWj4k64t
Sxe3Ipw/DZTjypOSUwnNktMoifRXQ6jdYXt8j+lhpCR3apCkPleZTg1Ac7kA08HZ
XdqgH6ZsvGwnBpuO4iPxsdSRS6X48+pPAoFxw03cpAmCo0Qt/kYZJ6cGkfxMTY1c
wqTidDz4/4vA14m4+XH0zWl5KIhUZ6I/wvVX46iCC12YyLvDNAwAzLP+eLd4kJLl
S3dlo+gGyThcbpD3Es4biT66KLKN27TlbD84yb0kubF+yAVGoU8JZe4X7EPr9u+G
65Guh/69dHrKa7IukhYTEapw4eR0YDUfZ8XmFlLdAoJXC5jjV5HHjWym/nbGiCSR
T5aLWa75jCUSOJ7rGgDVLiuCodZu2SUpjk3FGOOZiFhmWAqTYPh8W+r4+ubiN70h
CJaZYcACqBzeuBVxbqXhYUHVgIFNXEOhtmnzoOpRhjZNKUurf7XTcYuCPqxmJL0b
v7b+pnUPQRSj93tzlJ9xMmhXMgLAcOiXesOn6vKzvVh8ZnAV+TtKeQA7GCoQGJ8L
hNdyBb1L3+9NC9HlayqoQYYTQUuNRbgrQNRxG5DBGAKQIQPuyhPSUwkR48dl4jwH
fopyll6wT9vlxc4b1Pyw/c0tkHBxKWGNgWPG00f1X+nmVG6hbP0Fh187uUiUxZLU
QQ8yAWRkOfgsdM0HHH3dJ3qoxcF+kHjtDWXjWAVTUvQusBO/eZch0fCOTAEI9zcE
HfcSsK6mfbslZ9/a4YMiJpWELyFRNNTVYtEcAHwYGSVzAKUYkjJ0cXwsEq5yYnwf
Vxt+aD6MXUX7xgdfOn8CN4Jl9bPJ3cVcvPFS5GV4V+jOjQpgM8jmmvSAtPZ7E6hJ
o74KBdOKfV6ZshKWgn6afFuith7u+pMvOO9P5lt1ZEkULKjDTcx9FTFZ/RZqhEJl
2sJbH18Gfzb0kaqJEB7Ep7f1Ln/7ZK/S8A00JDe+N5QEsoCmDtG5O3X7srseJcXt
kaapx+KAwZAKwkFT4fF2U6Je38v1sunnSwJBrPMImVlQoyzoWJ8v1mxKovhwR/J4
9+AXrwMcZVdtTqAfIJPX0V8KL+XuHwztVbPhi+tA+i8THiS//NkGsNJs2gmv04Fp
3/YUZntBWROO/f4EGAsiquoNKBoYBelkP6hUuAJ3HsX5czVw+kOL1y67FdQiDnH3
Tgu8um8yjXlM7cbtRS9WRqEx5/va5ZMaX5aZqc4n3nqcTMI9kL6OYgsZM9qKSkSf
IOgoS2Ssf+IorLmh25OEQpoDIy0iKM/72Gdy3PRboumePAhtLXkmejQf7WstrIVM
CE0sp90rd6x1/EiC7NoE1busiCde47TmFRACq6Znx2VoUszN/iwVUsr14VF6t1JX
d9nxNK7W56keFou+AtT/ArgGKGFV6wDvGrzfc+EcoZkQjQeP+JDXSHd2W22iPxFv
KGWsrR00AJMei6Epfx0DBO78PDsYCYBVA3YuMLAceNG62TPg3lfDD/jZKBwMto+g
zLyzUc3ippGRA6MQ56L63grlgQ6RMHsOthivIWEQ1u3YfVO+oRUbLLZktQhZu/fQ
oYdSGgtvGX139kW2ZM2+7lzF26vRE5k8PDskPb0WahoABtBYP4mhXZlEWrgAQifD
9p7c44SFbVZCrO9eDbY7N9MkDusrTfipTq6/PleJ9tkQZdG+2JdbZWLcEpip4DYz
hsynCCZxJ68tOfDg2XUFvAke8+9YhbpLrx1PAdExx3w+FqYo8+vR3cXwAJ6RgxL5
ImnObwApKXPDv84mnGa2RObpih14v8hrfMsVDuCSK4YoF3324boh6skHXuXGkSzb
hFADDi4PyCoajY2kXqxCXYgB8O/exQRJ1M3meLOhCbUVtf4/PMZenWALZ/6BNQcY
nsn7p8LvJm4gowByF7FOb0jiyw4KHn3FipvC3VA9fixXP4DON4rTxq03W6aEPG4j
m6KJdBkI5PBgdkD4v/pj7OZsazBzVCnVJrMTPpWKrv0ukGdqlCikOglWn927Xh8N
BVmOsUO69t7bSvu/W5KDIcONCL9tRqhxEEQZ1NgkLkudSPfihHKAbhoSYbb/hDGJ
eGq8iKPeAadOFIqwK9cpL7Q4ynB8ZCylSO7uC8yEZCmLHMd/5DZ2fnfVColTI6La
aKf1o3Upd/O80jO+p/4wRRdzsSp6ZhhgupzFTTkEnqfeh3qI6Yrwdw2yN2Em1TWR
MdMZ+KjigzakL1guabzE0a5ZAGc528XDjULRExTC41DM4TWBSF8pvLIEfFBLdeaC
SauB1W3GeqYO/eA3fU0m0yqSe9Ow4B5D9cSmrR6vTL0McsBZLdNqArtCPSjFIOHz
KPprOugJkhwgxayvxRrc9bh6nXaXQdzKDXeEwhb8BuynX7BK6+QOCfEYxWfPMJJJ
hlVVVEZnUdZqneTozOzHvjnDV0PwS+UdMwrNqqveLrpz3TJiHAKGvYxMtPTgHCt5
v1o3qUcVgFvp4BU2YIbM7n+jAnJRKorrrpJCGacQs3X0iC5MMPGAJDcI1ccHWQ6A
UTyzJdn2dsEy8kB3o2d9dNSivHbpmpkbwbyx3KmnxCZ+5GqXLCWyP3pnzeKAztmg
dkedizKgdzoA3uV2uFJD5xO1osZD2JXaQMhAF4S4/3rRn/1rUYwYZzeMAwGeacPX
R6MCDAYzWE9ZQh7ZjWIceuP3L7lE/myb2mCLRDvS9e5IoR+0vU3YY6Fb+O8PG/HM
jvNwvMijRCEwuzs6mrcBezmXWW81qB57Snkx7Kr+T2+nyErFq+2JcQkYB1cDL99E
RYPDxRejGfneV7u5T5F5pg27tVwpkjts6veVC+PugBkZqwKW9XHZBvyxXiqD+Zo5
+QWXRzH70mGb9P79V7gGAFntJt3oVrDyp3BOHju43jpSbEakwxnBY5trW/mlf7l+
xldRE+gwXBES1ViQpP2xisZJsH0K6u8IJhuq63uBpBRa2Jg1nnP3L6EcP2MLjnOQ
x34PZDd28Y2aOfHhHHxOW1HyG3yPEp4STvpXW50LA9+z3QyEX1x06YvW6vlwjt5t
+eBFEjVFKrU8d+n4tRLp66lvQurrgKiZoEVkPOth7pcDzq1rd0CTPNzHD/4D48hh
gG2tDSYDGvtyc1ejkeaV77GNN1iuMs7D2ZMAWzrP2ZL06BwcEFsABMr+uqp+YHfl
FK9Ooy7gTycIivnlzwzMUbz0i6v828m+C3vE1/YR4BhrVl6+CH/tRxqL9hmlScoU
Bgw3hLQxcEfzhu7HVhWoKj0i3Wy3fDN9VxbQbbPw780euadFbRRP71SU7cTU2/cd
G3mRUvptcVOOfo9RHzvUMuEUnA9o4lwFCw+nd8VzhmoCbczloc/U4IuoT9x0UUeU
z7G5yuwj7pd/e4nzmm6l9k/aPds+0N/UOuoSQ8sfoA8T0ouytZJnLrDvpI7TYsj4
rd6wFRqOgua3Ck+aUDA1SyAkZ7IbSfwDSEpBY+YLhCFjaW/ep2DKq/w0MPzdv0zp
AxmgWCWoSAzAxRpn699/+fnq2HzwJZj0UQosRLpBCzh6rETPH7B55/XOuJgVVV18
Jtl4bLR2vy3ih50pZc4WBqJ2FmI0n2H/vFWGsjimWj0lntVmI7tIeW7p9rxJjF1e
LUM8dBtfX800pLo+J7mR8Qn5QMCbW3Amxs1yYLe7XJzqvk7bA3OmZLCTyn3DS8Nf
fq4uG1PlJDV4GTe7NnbR+SPb83uOkDQeYpe+hyeQdWWx7BP79V4CyqJZ2a0dyOJ1
PApT50ajlNBMs1nGWfUZ8CCDA2XJmWdIiUTtYSBbSWJMdXbemQ5bsO2Z05/7M2nR
HogZloJtxJqdFz03mHP+s20OQw2+/GdtrIvSikd8x03d0OmUVQ+UuNskSh5NQ+p5
AfhmNIHlEguBXHzsQX6cghM3ckhisRyh/o3+0aJ1bHtxMH+h+Nnzy6MFQlhF9RiP
pVlfkhP4R/vDeunEcNxSCcqhDPdsvkoBcHu9mfY3HDlNVWFOMEo/EwkT8KfrMicG
BersSgJC6OUb7bQOYqDxfRKVWfmvBR7XvVfvWgoyZKJwaqhD1dntO9MUjjMgWUhu
tjxhNT54/zylDL7+eGPrmw6b7VxmBf2C7c7TV1xaHxMRCMAMB6IBFsigDcoGSdSh
UHLZTNcSOH8jWRYM/JVR0uzf0/X4kwQu2BDe+65a3a+VcMMsz8KbP7N1ZOJmaUK7
YI+M8jOPbVdUTNDk3XtgcBV5yYF6GuHgBS/0fWiM5oOogYGWD7+tqGD8sLgISloy
lctgYuKtLeUZqEFNSrXhO3+ufs3wZpQtiv6IKGuekeeGTA9vMWfhsUGSbAvQWrp0
dK5ibOI5PaADfSSEPm+HEcfElz7zvy44J9MVVg3MZEftwBfBb2YRMuWHHJJeP3xH
S0uVrb0qZlBJkV72xxhv0y94bOR21tHYpOCgueJRXcWrOXzUCdDIMmhGvmfsKP8m
pJawf4AQBkDGHKv5BSYeOAcndYVtRwsBcM02Pg8IxBwbZUrJ8gehIgmAlR/rt/Iv
y5Z9dZMnS1hEmRgoEcoBNRp9H62r3rnVZJSzoR2u2LOWs+1AhPxx/wZOW0wc/3AG
rLGr0/iwPFWFzLVT8/sRU0RGI1LpKFa0OI994eeTJN3D3ZC6fL3m9IFV79YE7e4n
+J6v1mbrph8z+QnOQAKgc5Ykaj8s0FWngKT2fClzvHYx3saMS7rzk3G358sc1+Cs
UYljQbZwndWTc4rwPq0ALqybRcLAsXCHPhO6Lzw7CQl97k2FuMC8uPo/UVLa1C1A
VGKj82QKc8v8lm3XFCgIJYQ4/qGATNqro16gAAGkSh0X+OVouWTbnl4WdOX9/sep
7shRtv+XtDkyY57+9uj2ey8C/d+ffwTmVT3C9JSOiOmmLgR9DBCO2YdXiuFvdc5G
eOHbPZVNn4kqn34D2pu+sYkl9R1yTXn7uqnifKiYyKOIhQvo43zwJZElugiHIi7W
vzEbl6y21Z+fRE5Ng19r1DoXwtqNJ46ZzuORjGaf+SRHdzMxh61HPJwYkUcWeGta
BNf6XBdwSHut32o2YFA3Ab1S9HM8GIL7zdHCgZuSNxRrfWcHvfQpIXpG9bZkyp24
uBstNhLJnMaw+rgDChnSCjCYrE2UQrol98IXqIeBbM+ds9VuJ8q5NsakUrFVLIR1
686nCHKp6X47lDLGm8zJXX9gwKt5kL0/K3Nuse/MYIvc61/7ZpAi87SFZStGJWvV
H03e0D40DENhARmvermLgn3oMs+GpqcLQYHDPxJmXJz1ySQiludq3DT+12K9E0u0
bgVP0ErmvBgjnjJgf8MkpiYPeWQl4TLruXaLIr+SxyCgl7xdgNAyFHXYPlknQt9p
z0xopWFgpU3XtQtoL91SD/Pr4HP47FtZmU2L0qj8+rP7OGU/pMZfN23k69vw3Xj9
RdDBvzqnFuOGIWpE6ViaA8ram8mkQ0t7Mhe7Sa1K0AOJzJCBBFvYg6aSZDwR5JvN
jMQk+kLfXzskCgBu5URrR2nTSKwH9kj/su/KwiE+9evlExX6XxmlrLQX9bH+xr7T
uexpRqY5/52uziD83CeWqvT8fifzI34OGn14/7SnsHSq1Ch6cWQ0Z/W4R9dOiqPJ
s84rMxlr3RoL5VMvUKchK9U46oS6pCVJhJID38eRXVf+Wn6gf00uGn0lISsua0je
oGo5D4TK2p0AvK9/PXNHyDt/jBf8lf989rBVJ+Z6YZO6mwJ1uW45tS/tMDXOH1nF
3BqJH5V34q7HZKaljYtXsVJTdHSFrXExSNbYo7UdODEecF8tLp0B5QCPl5yTygdY
5HisN5SmXzMBhk49KWK+Aw1mobL1tuPPrU45bwQd9rColRxnafB+SS8wgqdPCzJQ
VR+cOCrYArSJayaiLLOsbVqjBhmqYh5a2RssZqyUDMl06UU64fqiXMfy6Nlgb6Ym
EIxMsvv8cce3Jpg2y/S6pQc063kpWgOMEXWbkZzCysuE46/GIXFweFAdYb78qGmT
6yRXWQyU5YTm8pIeVpzTb1joGGudJ8TUGXBSNkZ+89Tw6P1B9EMC8TILk8HgKLKL
dcAi/T0Ipi5gfeAaX4QOsAMvFhcrHhdHWshfZWUhariTn96EkshkSFJS3mdVAznB
8phJIzOBlIY5+PD9bulp3PfFda05YSz0OzYqn9dlQiHXIwxzwoG1mElEOzLI5jOb
UWjtKhzwo4YkXky2TrhvXo9KSnmSdSPGkZY2R607S0AOLw6o4rWm9VWZLsOPnwvK
EF8w92wtIgG9JTAwT+nKQiitE3nnUN3irWmU/hWdLY6l1LMeR55CaxlWbhBv/MvN
SMu7t53mU2I1LP6eDet9KgtMx9QUjVSPsF2FZlk0pxbAK6gUwFdRmXMxM9u3LUKI
VPZrEJrvwDaL8qUgWJG1uwOQv/6EGtv+IHTzKeMIq+rsmbFXp23oiZdaHJ6X1CNW
N2D+I79H3/VdQN6ZiUsJ0M6FylZAIOvp63mrQVY8cR6DpoT8azD3eWSw++92J0dR
ncljpf4rNTAWoOZREb5jQBOUt19adHEkZaDu9sbHBlDH0iUKO7zCYTbRhD2sDLqW
JxBLfLgo9eeQ41TeYKlfWRMj71KcrFn94bLAKd7qUsNZc3GInGrjEvLWodNO4/yT
zL6m2num1U95nkl3wqIsIXJtAD8h6vkHWIehGDz22O9NbuAeMJI/gmXSMS4xrQyl
zh6TK4B0EM6ofH6B4q0l4zvHICF3Dt60ufKAD99eh3JxP51kab+wwYHNPyTDlq1x
uUblFOBvJVNUqIFgmwU4jpBNuYuEMRSHFsrU99P0NlUMiFLOTNzILoTkrEc6d+Oy
O5DhkAXbLxzFHLP8IBswIcEtyt/Ys4LhbenTZmMnh1Tux0IGOxmI/Cplg2aM0287
Sf/+XoAicqAv9uFbJVeqwE8XcQqFPQffiqZJaA2+iw+kOp9GlDKW+tkdBXHraDpL
W07BgM1nLRHmtwSgON1oNXQN/fNdkWZciptPn1eAYQg0rBI6vVihbByYrfTGfglN
wYJN99N9Tf2FW+Oam+qZwxpJx4mFxr4JHyhQe9TReSagZe7K/xlSGoVNw8Ff8uBU
nFirAfYfzzJkJFJUpNmhFsjXBocJm/F823AHchRSnTPZ7wbfeG5/socX9jkPF1i/
NXOWCOPny3y3Y1O8UE4L+imq3qgVymZx0/pASGFzdAn0xETftE9PPylvjYLcf9Fp
PM9MqrXDtwYQdRVMuBb0yH/PD4e8y56ByOLAe1zACsFG9NoTTYXMmqmLeHYEcipJ
bawutBIcLY7UTOGHHpgH58FMHX0bj4bD8MWUYtoLPNq/cQ8N6JcDgWOdm4LKNWPT
nBq6WCO5I1tltGo4x0kjr0dKrH/67SBkYI2AS0BSItjS0BKh65Sjp7D9stdNO82K
H8CxaX74xoOOqnnpSJkbCv4/PLFSYT1DaX6Mb9c1wVOKDgn8gfF9r4iz+GkPDbBM
WtFBiwodvr0MALfMA6mrAQon7oCuruP5joVo1eEfsOS9gYVzhbDHeR1xtp3suLih
W70WnkUaeAtDw9WsX3sa4ncGfgN3RVmeCYRLFR3fS1/mWtKfyaOIvAWAC6uBphsw
XT1AT4UtrULoxyjpQgwDlMyjaFqah800xRMKc2h9nfRq/j+nkpg3gfP/7DPNkzcn
8fK66d1bxTtYYPeR07OTzkyvggrnYqylqGyjElEeB3MzBnANrXL7to9bgjH/ZkCz
nnJGvJjk5KMD+OunNMkt9WwNCFHtkaSFEUyWo+Hxee3+6OowvCXPlzYkAHDm0BIB
pJWKUOQFB7SgxG6P2spfmPTOdJKZPalSDs/UHfQegC+QBpoG102ozAviT5kEyRqC
qm6iiwVHwlPPAHtlGfSh7+N1fiVd18cpgDE9gbwKhvGP1RI2cjj8M/cGhTGITpoy
77L1Ggtt90yI9ne820ODXjrfrc9R0moiEfZ+8InByvLYMtUQbw3ejMyT2xQgOGSj
MbZQbOi0ejnsO1zbSgAXiQgO2GfgFGJl54zfpA5Fj04y+dWrhy86CEJvxJ/84gsn
o096VU1ov3ktz4UwMLCY/x8atQEKaEd4VIWIXolG/EOdtmTpG49Q0/85v6gUhlKc
Nhue/4mbdzMMWEhcG0hdGOXN95ynt4fvvKa8/KN8O3D7Rz2whfIlOBXrf2oxcaGJ
qyd3nI9qZssRyR0XY60Iae9LzZYV7Zk1sQAKckvdgfJa6cFs6UZDYajXZbuZiA9H
sSnAxSTXuOO8W8SZpgV/AFByPvDrK2fx0/4c/SmjgT0OnogVcCXLt/7z36/Y/nSW
T5FZQ/H2sbUqS26a7UfTxwyq2irP2QEFkRbMaLTBcmRvLrAJ68M+O0o7DCNamAkj
9B4ANRXKfA73mp1iIFI4jwzuqmQ4z1+CWyPtOxRMgBLryWSjqxEYi+LbOoOyErhv
9RKsRMfzpazVWeTNBoS/iqRHNjiYESsy/MJFeiGQFEheaR16REfE+R1VArzQCSpl
jR7qcByCLo4mhz3+h/peeLdJIElLU1BqE3Q1mQlpeWISQIABKcvMAEdtWG/vIDVm
L0mrvEirfP6hrwE3f6vRCjD7ia6J1UTiWSsf4h1dn6gIy5F0Qin3vUJVoVSSWOfI
KAxhh9Osmn6V2XUZMg9JtwYu8l/c0y+rnBWjXrDReyUtfx95FSL4mj6h0mGN9PQE
U0A9R8M0o4N8ADRH3fyKm3SYLfwR2KYZ0D765jl34j1ftDs+V4pNcg5Hz1D05riZ
M7wwl+oZ2O8m2a9vvc/GrA4D1ZXxC2G26H26rd3jGTbzityo0KP4cBvnjshd9C6b
xfq5zJguog1SbYzAPsKIrkPW1bXmmyL0e7IM4HzoordUxONceBAjNUNcK0x6eNqN
dzDudJpFRWmaoXOl+AAAVyCRup6IPRIBa7cUO9LmucbutYgtaEAXYvkabKvOBoJk
DwXV6sHMqr7plHlzWuo5fVYDCCtEXybVPlAUOfUKGliZqCJ9KeRKBY/hnXupAenE
OLijMccJdMPamrGvaBxLZxQ3UyNUssIuQ9kd2O+/ZD8NeH1XReqaJlf++xucMUnT
fvSsIX+fIpto8ysMU2hj6a00OW+7hPPeA9jWaPV5dv25gd7kqU4TpNv4RBVCvzUi
CM8cJdW3W+i0hVasblKvAliD80HT41Gzskbpl4Eha8eWh+2tVu6/3HilsFjL8Gaq
0wUhtjtC9pIZMt0B/S6bYVYxEWt1dZG9xiYvze3ST4NgmQZTjahgSLuyD/m9MvIH
xMpp+xsIxN+gRIaxp6q/5wpM5WpTQVL6IiWnFIh1d1GYO7dJj1Ajtg5HYzKa5B4d
ZKERntRgZTtwwQ7wDuGC8fen3AAlhpAAnEQTmll9+ULZG9dBBwx8QcpWi92ZzMqw
ZELUlRVYB6BH2N2V+Urt5kalfaNutYTzU/ZG/LuIZrnRYuObSqO2kUSzpNpRsXyk
DStlYPP3PuhjpxSiAkXvYdXA8bKQ7UHOXjKUQqmIafkSc6mghYxIJZ3UjmGqKFmR
EKsQrNVWE9G4jnnKI0G5FJdg75E8OLZE8oVRCNumMExJ585BZXok06v1YeET/57f
8y/XNb5DyjLmhvEbW9yvSr3cCrrm14skIpo1WZWjaco9Chmmj825uSyIOdWE56yk
EvJuYosmfwvyR4uZbRqSZZz80SrcYEH6xQeAi/xlQKL7YON30C+t5hRp3kCzexYd
UEgWyWR2anDoCH+Gf9kGv/sDqtUpzmgRCJvNnWRUK3oIfBaur/ZfbloS2N0AkcBy
gcxvy3PrMcf9qZmty2+EPWbCTtUNBVQvcE7VKzxfjwIy8JDcXSrXoJYJClzaifOd
zWwbH0H7MimMsS80nyKhIz1ld7TbAq0SA42Z0tAlJ/NL6X+/61fqiSBKmGiJTusV
ffCNfzjKcNKKXtqYU8cJYQBHxXb9D7OgiGVc5Zo6heTUDuIAd3spxz7CvoM+OCJO
3a6LTxPTwzd4zJr0q0fOURkQJuz9MK4ZBEHXgWq52ViZ+T4nP3sDkLSIXGUvrrKx
Iw0WpYtFMtwLKtIUq0dltarc4odtsSkG02jtpRYxCzawXFeGG9KZUsNCpcRJICoH
gAZkC+NSBhIoAorH0mSANCKR1xY5HPeFUIuMGMl6I7uXYxmjI63a41D4L5e7HJ1J
nDaEjUuE4oZU2NXJBWAHo4fUqZGVNbSAwp1Jah3rk4hLH1NnM0cp/gyxJXaEOGzn
fuG6+JEs0OOnffRUoEoBDs7ws2xuvmQfKsxtmMKyl1mgf9PLPgrH4te6aAxyP1Ky
C9rJgdsDhm4xABQhF+oJdk6s1Bu7spQBoNTVSQbfbchR3nl2Xc1fXRS1C9q6pnIJ
5ADW8dUXiz5xYKQzquyJxK61ZsX7hs8Vla38xOAdkhCuNRR/xiJoMjolQ+WdU5c2
t6FRYCetRSo5RyMDTfYxFYsl/5iFQH71c1v0Ch/qjj91h5V+SW6XRR55O1V1hv50
rd+WlV+OU0QF6MiWjO3f6bzEYNe54zq0sqli86rSKmSR3WpYohWuwUPXyV04k885
S219IjW6r181fbIauiRY6xFjsVfonXMlXC/h8xvxszDgd1TaCQTKb2+OE3XMf7H2
nd7oDBZnjD3myCdKuANCQ1S5i5pXE50p3RzwZZZBJ4UJ0IAXdMqh4OGrqPB6NnyK
UvQsjuAkTLLD6yaaC9MJTXhX9SsEdAp4RL4AXjX+fgzlLuGimUoz+ECdOMimNxtH
hoglGvrO4mk7VcZ2IhcCIrBguMx+CDp1gQrlN7dJICZNzVUCLdGjwoFxFqqC4UcC
KnStm343I9I0uh8dAda19feNqznfGqBeWg0VhR4+9USjpFW3NCoag4A8KLEb+DxS
Cr1DRyuEOjYjJ7ReDGYYSLBrGdh+G6eYdJ2qhwxrxiyeKbG2FrkIrsHThNZNT21X
OfPjMyxJcefDodR8nNDByjfMeH95a+689HOjdwFzIUIQJPHtr/6uYTzVWnWq+oP7
82uewe01l6oeLidvE5RRGp2RwJWMa39gi/Vr6M1LC/PzYFOd7UsrC+4IDeqyzIo0
GRxwVBclIux1DpAy9pYezdF2U3yyGHr/cddW1qZJ49l4HmQXjvj8qS+PAv3P9BYC
ymMm389PVJncFOLXtEHpz3ure/a66RLykYxblMRjJql64ftFyM5WN/BIHNABxkhp
0248kXXxf4/PAGFVW8j70NnZQCvS82HxFMO4NYPqTPdnu5iPXp3WifK351+5Ws7X
UClbCOkdIkK0a3PoiwMfm3z0GMkSswPPUdcCkxpTFz8U48RGLDoCcXakHFkigDnZ
x1GxE0xIMBihe71RIzIeeTVKdcjzHUiAbn7QSnFaydRcwiMecaV0eJo1KMRubk6e
xQ+41l3q2O52FX/uTcUnI2JbtcFCt/iBgIfEDmz0sZR2HS3QbdKCyyG41rzrbaFz
jjhG98xzM+ECtrEdtCuiwRw7HKUbeMsgSRqoD986dUKbGrLTfqEtkxyOVSJKw+Qd
+DpO48vL32rc/pvJjtdcLmQttJ+fwHAF+H34oFH/4El9xOF6dKiZLJyWJyAdGdPs
dlu1voYEiUf0LTjnqowant/j57jwcsMryimJQ4XZlEba2BoUkNj86xpXs8odcFDi
ZmOSS6u0VVsajRBpQWlW1UluqrEk2BkKZ5QQYUVtI2b2AJ/wZTzajXO/AgnGADQA
/3YtgEpjwkufBvijkRNqJ4DNyC3wB/XDUB1dygc7WIBaC6sIoJm6n7/AWDGJ62UL
erljTDwRwvJFE4O6PiqqZFA3cGzZdgwoB2NeYZSStXWIQth06KQE8UXx0UhpM56x
0AO4k4Skd/8ryZvCCiiZZ/nT98oUYozefdryjzS04pLI+7zY7iNwiz0UMgYZ8fHK
ytaP0IC47d9SfdFxk4PiVBYIw2g9eBPYZ1lStjoWNnRYkabiRCneYFi1G/EE3mof
oaQnRQG+JM90uwcgGPRwn6VjVIVJDJfpaKrVe90c1cGKBsPxslmcplwl+hynw+1C
cCduLo8OK+Tji3LHFPrxGKagFuapfgRxR7WTa3ljvmU8O+LGlWCcreFvjEkuI4fQ
HWTgIXnUPNvKCj0liHaf8+ri6jkiAutns976LgxmOU0Gx3CUrK9Ie3NT7jJ6jH3L
LeQBJ2lXVkGAxyCZU9OIrREJ8tE2LgELG5mGGzmuYJHh2OKMmXgXp+jGKJOSAPCO
KQI0vOwt/mQ5XHdeaMKiZkn4ihbTTWCvAlBeAjQtDhiKPWY9asxGKlJIYkZ0x7zI
OOJ0ZTNNj2ZEmkmf6WK2WsWNvqTeaYx44lwPS2XELucZFuMUUkAFWoKj60UFBF/i
KjiBi/yCqE/7x2B+S1CKGgepkIJ9jlyq9pkgv1VKY9aK/crz20nB5+eQgJSJJxOA
ex4VJOma2IiWx2R4Kghwl2melznKM3ftPv/zIJ3tMXUiD8Y8GRC5fhR1gQ/5i0sn
heEH9b82VX25rshjIcsGry2wWtEplghmQyCPDikUu7MTlk4IsycNOfbV0lw04K8O
TgZJSh49ldYAaeVGL0rvonEnzuf1/piBWVKiT7iXadI+A/KTrsZXAyAch0j2EFoe
ZX2L+2c1hN2PbnRK9kbFhzjJ2hIX8ovb2PXtMlKEGDjNvJkR5Mk3x9sZLcSvwcaB
H7Lxxz3uwaRORki6cjayuG8C4cfPbcDzeRtGY/kY0nqEnxW8uKeHvNtktVoq1C/D
VMPMuDJTDWbvrip//SK5tfEa5/hPPxE+Xduoxh1uSBYj3TtEPZEBLtFcQ0RdkQ+e
X7KJ9RoJQqECrLAetwiRHeY4WWTgAb9TxwteXASRrfbfbAiWyJue6Hm3GcKUgnPt
E/QRBRK6NDSNZ+j5JOBbaoolSpFb/Dpzmx6lQN8pmbGQSf84yoVUHTXJZ6DvpBxM
Z6WTJUe4w0diYcpvn4wGltfrWcsWjkoQqhRXiLTwq65T43W8CQZbARj6bslL305j
XymLs3+Mag08xjh7IMLFQQWfiTk+IfGjRWZC0MkalgU2N2D1uknMMjo0cPoyU7vD
PmblktZ1dBpCZQqXfQF4h690+0xipdce1xF0NPhl8+XjUM6huklQgeKibK80rDSJ
QskoeqVVRs8rjYEZhwhHmjipgIgD/bBpAHfyrMKs4kpMU1s5LKTQgN/qxmJtMj3W
LtmNDb1gqF8HhqlMgDIICnpIhzk77hO+1hp4/D47ZVRO8nyOhUmekNTZAh3DJR/E
8p9paWjMN86ZcZvyGGf1vZP4G4O3eJI2JNDm1btJ/1+f7vljnSHod4MFz+/IwMHE
v3IsTjXtKHjcenqcnlNYmWcVHkwInkXNBcQQ7Jl6FgwAYA0qGQ5nlG0hSkAHms8W
yzZfy5AhBeyn/cwYM1YOQXZjJtY6YyEcs/bKxnew03EO2fIi5hS1DHdxY+s74H2y
acn5hJnsWIbTyFRXqY+nsuLLBpZHnFBCb8mjU7R9nQem7r3TI9TashVY5z3mNQ6S
UTUdSAvfBXv8KLyDQSdDksEsQUp4e7jNeerNfKBJiJk0NukQ052/AASwnLuKNw7L
BbSJYGFubducbCKuKkPw5bhx2JATZjsPKxScOUqA8r1DgG6JDFccJzrUobbfD1yr
x/mfk5ki4txnnBQP4/LSI49e5QfBxmnPgQBpau9lvuGP1UwvqagEmzA+HBmy09F7
kQjA2KghCTBhH1zGO9zgfdm90vVqqerxSi66rXau5dWJNkyu/qzLNaB/z0z4C09n
LdBWvIV150S9Bub6y76svgomGrNxeAFn3NFkNHYINwY0y26E/M9cfxikQdtnrLL+
+9zQTGT+JXqJQQT49D6j1AG8pIDTBA343NTBBAWOwYV3ETo5nIuU3dNqls1evxTL
zqqzCt3ac0K0rff9nuciYh78EOcLkCrB5SAVFPB4FM+f3j/LRnERVnma/ofqv5VC
LUkvqFHyKUV/Hc7/MJXpODsJfpZbC5Sb1eREZQLfk8zrcMLPnEAh9Kdsq9HS2ukM
mLTcb+bzbyQPa9e4NOPa70mvHbDIztpH6th1Y7P34FY0sjYtcf46dzNkygyXsmeF
ERDgMsC1U2SCcuQtvBW0wQOtNS1/03DG0p7/Yuoz5TG43oc89f2P6RhAU0kWfecg
C2qXEN1gyO/xy3FmF6FP73zcRVC9En4ZifuoD1oYbvw0yyKiIMhIM8PXowZn6MJa
nCJp+Lo1mlov4nEdpqBj9M6qkgL1WZ0ehT28lJHvlKewqxxRglOkUWBa5jhhW1/j
S3a6/VSMXCG4zxgKIyDijEKPtQN5nXrq/AIB+j0VRcnqjek9WfvZOH3CIrjqALyp
//kDxPo6MvPjksDKn6KY+lv/kKvhgBhpEcDLwHKkkT14J3rhqA04fKHuI0Vr8uz4
qbFVYQTn8wmgQ8VKo9bbQBuf+G3Nopg3xyL30TwhSdC1ahHeMjK1FZ/N+kYNaEDa
EeaNlqxeA43WT9hDYDtx0a2zZUA48GvlmnQjIVvzIUKglIGZ+kye9Y1vczWYlris
GMrgat7d4uRtlvftkmYsB8JyV5qq2pXBm++x+Em6jDkNj83VEsex5rSuj54CumSw
uE5XOi2xma+x/wV/CZceHRb8rP36rZkkpAPOPEGx0yv9cuIMYBHnYiCKPThlazpY
ylvPQeuuvnw37+L08oNexG+7nBjNiZdBZSsVFJDmCO7GqytucjS/XYbwOPuJskn/
lvrPXHBFuCmJOJ5dKsguol/0zISOGXhCP+cOp0BH9vsSOkdvwYk50nscCo53bmKY
irnxPGUOc9iUC3B45YUixs7Wl5/SELOdm8o147Bz5C0YmLF+qkMxqjDC6FX4LMEC
KzuLf1RGUy/H13ZSkh3aefvioGpkcDaTAGVffvvM9rcT6WGorXnbn84KnWbgD+7Z
oLLExwIuuPkwgsuEZ38ek7olOJg6nTSqARBxpBAf52PeaHLo8JjtTPvwLoHh540K
e661wQYS82C1Nufm34S7cuwRtRIBZFZsSuKmIaSynZAwJ7pXCxaA63ua2RMwLnxx
II1cCpAr/jVchapTLqY8jy8R+snE0bNu2VAczIW+GtS6PCj5TbjfdRYyaGg49d9P
2/USdkyjyVh2ebXruJlBF/Z9mrOFzsojUd2dqzTaJLr7uAHpbaBKrB69Ss8K05pA
z1UZldnt7hUToDsHC/VaJbNjOPBZjWFuCW1LJhuQ4EiaX3xeMs94I1/wPVWDs55U
oJeoVtGZBnjDobNDoqGiqJnpHRLc+Foy/0yizHTzmsZq0+n+yDh87inzX/llsb7w
B0pDnkSWMtH9PROGaloUhWnyZRXroR7EqzMzoqKRuYsrKASJDgXzKncnWyDwlgLV
uYlAngJuk7SkNoL0+d821cijNGcS4FjOE9UGByJ35LEI4uLsFAi9tmm2rxLX+QIO
FwbOQZO61rCfVUwjkMruiwwsDisu6BTI84yienMnbJba68aK1/F7U1V0hwEk1XiQ
OCwj4+w+xBnkTZ2oT6wp09MJud5iZOJyXlDquFJYwSlty/Fdv0f+UTOvohhgwtCj
uL9ePBug1eviEY/OC+pSeFR2mpwtrH9BtAx7gGh8+ndKvNSuRhAHwdTT/khFKRIf
5KGJIqKsJadEz+30VxwdpNJWIep6L2MbvYS0QdRbTOQP7tzuTRi5gKbmm/YqYeau
GX8ZBFL3whmxQC5Pc7mTkgWFUpDKxazoLPFCznRiXJFT5jpqMe1bflsKPq5IasF5
viMucyq11vcMXldzRQlLYs0tuaFfY07rAzYbHB4vCKoW5Apa1HxGlHXWS4clOodA
UgpWml2LlMF+R416kzCFk5LmX2Lf0EsX2um/RrdTZbXSMim3fIKWVDDO2GUNrC2G
mrIceV60l5LdNb5ASraLGvuUHdMaZXYg0DCyZuQgv9rizc3QDUb7bYlV3IkgydOI
+AetOuP/nIRudN9YTvg/bMGUIwIWLGMS6P1jGNSQsNLxlcEdVOpBIOuvxSJW9ixk
fP4ieulv9llRLsUHj+X/k2FrfCI+phfh3DyOnnIAmyUV2d4ZW8SHfyp176/XJmJ8
REp87ZsqsmUOPJDzZARowzXM7TMTUvB3zlZdC9PHwKtnO3VRiFeEDFnoK2eL1a70
ROb2hOthmhdEP9GgcZHv/kvf+Y/yPwEHuMNviDWe3urhWStwbHzSYRMW6w7g8Tp8
KqxwIXV4WDX71UsdsJEfLuWd2SeCD38eBR9Z44VrUHVWtwhfEz9ENeqIzj5UY1cE
nNA679aBb7X9/JgaD+s7KecaY+lvVJl3/15b/cVOTxBJWK6DxY3ANWDFCSRHzFx4
eO2EyGcdVt0C7zUMKw0QxLJmzD7+3Nvi32zO20U7Z+kyYRN7hDTdnoTb/gXde6dH
nrDb63YO89B8opIleObbptj40wRGFHtrO9ppG3eGadMivZbQ2gAdSFK7wmx/lrfP
16cwEtSfryRUiCaFOh52RyTHgzRFqWz6GFTMxtXTQiURGhb++iWB8J9GJp6LJg+S
R6Gw3FHbUfm+OqcietDVfXvrQaXYausC2GfTQargzfdU0h6MckHl29E/bvriMSj0
FIfFyc9vJIrUTVKw/FFsihglFLIKpDRTokJ8OeT/KvRFrU8jYv4FAjTxbg6u8E33
rbmTyPwkGrPCmRozk6Dgu7mWt3sdMoBmnUOlxh+r3EPwJLSw/eMPCDfyUCNjMgX0
w8DGzIjS7B+f3z2jC0fdVYdGmsT6QoLBcEIZvNmrg5z0Vql4pf0g2dzXmIAHAv8w
knT4Bg6aG9l+RNW1TfYIK5X2HHnOzY8/srZ39bJaNdvMR/QJMF8uZa6baJGV3G/z
wtFQgXYjjhzR8cf4zHgEZGkFXSPZEk5t02CnFIjAhuEbpoLpRDUSL7T6by6ovBod
bu5Ept+kmExxp/8HzMbwAwb7Gkbwuic8UW4NsW9QRbKzcr8IM/7MtB2KxhGg39yD
3++FLZs2oZ5awOFq/w4/aU2/y7hSKAgR0XlzY+At/HJt3DXvv10G+AyJF4WutuxA
UmgUeNfg6tDCgmlH7buqukXW/acmXsX2utjVap7b15aMrwqvd4kBsJ8SMJfthr2X
M/3GC2OfPP67JEKN5KvYWdiMYHVmENdYJyFUeMZ3PncJcBsjHPrxgy2PTZuoCsok
YNawAjBku83AVCTCPDkXG30SkkdI2vvN8lnwu1hat40PQneEriVpITjQnPmUTuaD
FbAcfXqV+xAXkd8DCT57q/qc1+hUr0UyFahUJXq9+cOH7ts1yVXIaKLD5rUEL9t1
vyLZM2NDqAo5zekET7iWv4gTQ8q+L/k6/ytUePX+zWXTnbSXzfaq+rZ6uZ1Zr3jz
0Cf1v8nOhAXar5pDZKO5AdBUltbR/oRO5wP+kPX+3yvcyfh99oU//bzyEIg6bLHY
PQHAvyWNpgVASg6kxXjznaSRk2KZk3JICZX54BA9uDVVo464mL4G/C1s4nKWHUKA
RYcN9uwC8CpA2oaGN8goF8oZQWswPWiLxjQj+2PF3cl5Vmh0428S4GhZcuy7gsxJ
OT5d/FFU3ohot4p7y3jshTLqtkqnhMdy7+8PmG4mfrdg5CBsywf8Po/AHYQBFX1m
EPLjszDI1pM73ftLF1fPrwzdu6Jdr9D29svh4CMqZivjpDFSlODnmRYWqGxW5lVH
sAfOWwtkOkULPZZRkVUSu1vZhiSlMAlK/DPAqep8MJ73eaQCzbKpTgom6Ce5fdf4
HgTwjx+oeuYKd/BsJH76EEuTXUuGsF79BMCvz5cEIKZW9jPP7ydLWXk2zaQ8enan
yzU3uk5uuN3Dpp1KYoBYCojbZ+VsVaUhNhCA1+Y+85bmb7rhoGd5wkOKnPGIx+bD
labWiuVS9MHTTdGQiL2lPSjRaGfgSEzyPmiW4YQBiJiqMhJVWqLtjqzEqGg5E9iK
o/I2Opadsyb8C5se2TUkmjKeRbDa46Gqb1TSUW1fX+bi9WVapXSTc7Lcu3mZJOxK
Oy9wjm5PaupBX5ABuWRQ1J9gG2Tb+QvC9K0v/bTXMqnsfp5cXYwctJoDBad7gWaN
KSLLu0FvKgGYuHaVi+elRgsVGAnjLWhO7vdlDvB6fWONRJyYxEdc/FMh0J5bBZLc
v2sbXQW/MuDjbV1WBEP0oU+paOQP995BSkUGV19RX9vXEsZPFK4npmeknoso4vQH
13LCXePhdBIGJddkbB6n79BVnbMbJ/seTyto7EIYJd38IevW2JCgKnjYSr1kmf6R
FWhQaMrqHFiveXtCAgw6ohkj3i0o2RLAsZtkXl91Wzb7drkQmTBx3GTqaKXGClIs
jfhPdmDE/J4TJ1OxTkFf+JEA8xx1wTbLQmwdrux9DdFv9qw2Y9xrLZI6VeklYHv9
1RXOKPJQx9R3UZbr51uO8pqeVkPQNWfIdNniXk2Z2JU2Hzc/+A3a2Xrtkllepr4L
uq1ul47L9HtYe+KAm6UvhjQMr1n/0FtVdDo8tJ4cKV0c3m0k/0RosFbs6CxnLYcl
MpYJcYVnJnF26ASJXqiZwRk0iImlDXXS4EFeOs4ljVVDulaNZ6v6HUpA98Pgg6lR
MjcjZNBNJgyeb/Ghbk/Z64sftl7J35Yu4lOsgfMjGSgupugKiJXMsT4mqLqrhHUV
TN3N5Tvg5jOhUPyh/Rgtq/44EDnCUBUbyZ4wAuh8LY9Sh4KnY2Fvxs0tQCxezTt/
BYbUnfI9x9APlaFwrxSWnZLk+ZXGWL1mMPTb29+xSbBuhLGHzxFD7k9e3B6dLj7E
NbM+mqI091Ie1SO2oWO8yhrVU7V+p1j/EI+Z24/ksm/SJAJRZ5xW7c//EExRYgPA
uQvEIVU/yHjihMbPNlNyRaFukNa2TwCXQi2gOYpGPX2Mipq/Hy8qOLb9+OUkwfzM
hLczFVsWMil0PSVV/wJUV9zmLyivh2+5wArfMdoHoxaHyx/9pNhn78Kp3bhdxMcW
m16Mstc9hCAa51FH/HzwOcAJ0z87gIlyua85Au67fciX2XqrLuNLeS9uGxgZ09at
7ndAL60Brt4LcTdPbOqu5sSkTYTop9/lwv0uKwwkNHelHNchrLXDMILcCzMXWHN0
SMzZu+e9yz6pkNyaLDjVEPi/VTIYF7iQypF19VhDZ3T/IK1BhS/hGfzU8pJBnCjV
3Pyt4bBqdpD+FaAj/Xv4vsn+9hq0BXd6OUfd1grg+JrAkrEe0I+oHK3J2q9ani1h
jg1Vn7v8LVMtL+6lJ8So1kaGl96u0x2HdpBPCvmSrSaro07PSVHdFrmLFpnnYsRo
zLGQajSDnOK+F/yeedI+RzK+i7D+LBHv1c1Tqbs/DD/LSUF8WyGcTGj7s82Zh5iR
gxOe/A8oG2qrPbQGl8fbSNfvtUNRJ07gidmAIA4tpGSewo1xZcyRSbap3dBiUZll
i1lic1r1QTISUOzJ6zq0wesj2sKAEwBrrlsHI0qvYtrbWj9aQN16+MBXU4cR/0ha
t02g5PVuyVRwGiBenlnEyUFosky4wqj+r0HFN8yRji9W7+JYGmJ+NR+h+jCsGaAj
4VuLETfBWn0MAiecOeJXVV0bVRAf9tTC67f8aepi1GjB7g717EVcrjanwNd2kmEv
GJJixQtmeIslowOTC1WKxF2uCT6I+CI69VlRAcJjPC8sqOjDpArzDkIsFpw3HEuM
tbc1XLZzz876igMMmzhtr1yqyNgzjGWin8/s+LD8NXAnzl8d5AMemt/DU/3rUsfe
RVzGuvv9iWIacc9c2a9o9i6vFWUnYTi3UlibDD19/YkOA9HYod0bTiF5RY3tw/lx
uRrK/Pvct1BZiah5ZcZaGS4hTAvfuBcSnGAeuMbTFQCJ+iaD1RRVTqLNw4oP0qE1
BFWWvdWPkgy1xFlRMqAp52VhdbvcgAMhPEedg7ZGo02wgV7t19ZBblTURGzIu3NM
CnzskfxFyNYtKFg4/8q9rzC5dlqm/oyELiU6Mdz7qwnAL0dlwbM22vHJFQ3CA+YY
tJTpXt6vhzPTl3CGZa3TmGkVkH8dbuyxrviXNcjZwQCOJFi3Gvj+gUEix0QsMXdX
9/i6DlJzlqXYDEEC7ISpxwRRvs3XRt9CdaVCG4aTuwinacUL3EurzhILUVM8zmiF
A8Pov+FIeW0ykCRk3FVTuyq62YE6cK00fHVOcHvC5mKRASpYMkwRrU9kx9SrjRWy
SaYLltMnH0j3SOpd+HyeZpM27bhKYU1X3gseRFDuuQ3biXytfB+m2MrkLkRdQc6o
5sthB42L9Vaqqo/yRenptoMHEknuZs8VqohAQ9PVeR+9M46MptjvDd90JYxFbnyg
HpLpAqljQEQ3BFGhmNdq2he19PY6tZxRbrI1iWmMXZdeMBxL+wNUXmtew1ZeHw61
dcYAILP3wmn8VOpgoF9Pi6xOt5I0CZS8UX3oOIvIeZrowhtgfwSJdTO2q8yagz5i
OB7NGuwgXTgNHMBNi6vPqXM2mK5JbgJWj96bfV0iMRprQ8fOcSPvKTmFQoJoqAk8
pbRGHs9O4lP0EX7bYoB3e1CPN0/60cdA9KraC11ahBIpkPz9bOBH79xR+b4H6C91
atNBXr2lDX0+LDRQ+DkUiePdTjcw+Z4Tv+hWfUPLf7bFLlBYllpIHHQ9s3tnEf1S
1qi0Bi7TV7CQ/qsp5VQ3frt/lFk6hGn6C6ZX7W2ukxXsSGmLljiZsOioGaKFVW81
YqPvK6MFaV2F3vzkuIXKrmeSS5aoMVXvEobrl5IN8aJCnRfGWczYIQTeORPLqi+v
/NiYpXL3Fs/8wxMbMxo/2tj36Vl4ZdlayAafzj/He5TaV7arCKJzQd6qYRxc/ZG/
A1SWKn/I/xNajFOxfCc30rE9HcY1Ad9RjyM/W5IbTGTQZe97LazdeOAb0PctkYVM
zqKB9CFa193foH5YI9lI+8Qwijxbhe6xPbWRHquHRbxhTPhWDrLf1aQ/KVD/ryyD
l8bKfLRAKSAM2J/yMAzJ0tD5Aq0OpnI/O/5vKDTuWlc6ZrCPLyKbuzrJFIdFX7lo
jij18P3ieE3U8Ls6KsAJ+MDFSAke5VogxhAWbSZbHzI7En3xFB2rz95wWIjiavS6
8NcMY2hEvKoTEOq31aWomBle085VfdzkixlwFTYTYtS4NHE5jc+IRSJUv9N/TfB1
pOzP8NOQBPTsFKl5zktpcoo7FSkkpwyFeI2/pkGykkZx1Sl9Q/tQ3iFP//PEc0ai
kPBEIqy5B5RbHwrIP6jfcPOzQJCVOT+8qpl3B0kNkcNr8+HUFVymi6JaCjdQh/Ls
l5q9JF3Sx32EA3QqbVcq/56sD7zmVyl34aRNymzgYlnYOptQxUkelHxXkTtovta3
xzcuKjLAcu/jhywyXBbhFhIxzUhhpufx2XUBdmeQGWFNzvJbu9RFov3NWmMoe+FE
71tL/TIXlCtF5Frgji6artW2DEIyWL4fsLKCz/ygMNXl2C3EWPPccP8xqy12Ek5R
0q7+G/iUVSbRb0cFATCmT3FUCY9RHdaxG4oI0svFp8/s9acUtvjmkQW5mllzadww
teeWQC9F0FkcxOybX2o82Rq8kMSGF0y98UzTsM+4D6n7kKfgp0LGhRivP6dwJ5T4
HijUV/4WWana0IrX+oKX2QN9ljFOBzDoeI5HawLx7f7a6Peg1/D8nPQFsCXG6Suj
kj0hO09chZqLdR2Sikfc7KlFMe5jn0bDOmDNqUnhFS3UwNFut1g8v5QoAwnfp5cl
F9UEdT50UMipo82PJNSCjCbvQbtJPQZ4jX299rXbObR0n3F0UYBDr/Gh/WebvSAt
/WWAJtWvSwl8/K169JqVLJqMystgMrqXoslp5U5jazTJAOw+g5NoORmOeZER6jQW
X8+wtdoTiqjOkVW8T4cUDDu7qc6qOkSt2wX2Rv2cw7Y8ShhgoAOoR4QKpvNRd9n2
eVMiMVaiQjERiwjbC0wvfR8bmtlPJ0Ki67n8BBdlRtLIO9utcE/hXJmggjf0aoir
/Y0FnYrJDK8YOwKK1lbMPCd943hVZqKXCI9rTaowpWgOmk207R5XD4/Xi1svP3K+
3oc1F+yVFN5aqYDo/uFFg34yZOec7U7QimsN/6aHgprAYpNyMlx+RLVNtRYiC4rX
LOaDtlJgCBWS+MiBh9tv+yEGz2ej9znW98aEY9ZwsS+jEtVjlkOwcecNftJLu4rO
BomNJd2jO1A29J6VDtPdNwumFxJg86pKWyYyptJHqgveEwCTg+deTmbG6yfgzJT4
YqzZt6Svx3+QwsnNgZCdyjcmS1ROyY1ZYcxavUmjtTES2LSuDn0kqK2lHVH3oC45
NpOchzDQdZzDHHCGxHmjoU1o8vm7jciXJhcNV/ei/8ufKO7zBrcJHd/huO4uwute
lshc+4W0K5g9CMPI/JbFnjodOI6fuLVT0HKSSXB4z3kb7O9/ZrZSdOUH140jXdEh
E8hEVti2sSWfiw4uv7CBbY7+pCZfS3JZ/YmUwJa2ZO7ceRvb7IRXqCzJ8FuLBFaD
lUm0MlC//KMs6gOQgkGoJZQIqM1V/Z7l89JWYCQ6vpdEfNt9m4bcHfYsW2PEI7IR
GCCb54ub27F9owz4tjOJlaKYrcghrnAIl2ZGpSOlhkdXIuR4bkLfevWvpweShMU2
5mxZ/smJcJvFrj4kiUuWuzyp9wR+oKHlzRDbCPQUkjPUj8zdR2UsaOD/wSQo2W5i
2bDd/I19w6bGLp4cpeF2A1q5RStjE14Qwf1ZK0Ou/49FGvngd2yZGdXlsr3Ijdox
fNCvYo6gnNZIA6Wd2SWQ4r6L3Y+KWrDfhg0HFKzNIm2SFh2QuzC8wc7d0atZ3WCD
xEv6n70si3I3egU0RssO9rdmU2Gaq6pld1cgJEhT1fkV7AAxOr9Mg4FuhM2negc3
nXK6ztZK+G7uqgkHTrhLm8+iMwii5VcWGvCPUY7bgo2vs2hqQPgjBbH/dehWO5ZM
J1ZNAomi0a9N7BMey6mOokdlPFIxYEZSA8EEQ/cjBGqS4Ar5/MLqDIHNCxtc8u/o
/GyV+xjvyOKwG+SPebKfeOsa4Igl/3JNpLs+d/08UHle8iFPVqBRSrmOD+QWkgON
DvLwPHu42gTf5mrp5u9APGiHg4sRnvC+pgq4kmwe65y2mI5uI364WzYvgdp7fISf
/Y03OUaFHcxVBf9Kl6qwyd5x1gMwd/LqZ96UdfTqYTHx0rpUgiKdEeRRQ8+/+w33
vPIY2ckuuambwuZVP7sTzru6p0otWx4coFJpR4f23nfhoNe+s9MQjLittQv2i5FT
Fa/b7qFfn4IB1MFhxQJGh0WQnzIF1hW03VypekwIc+OfeQ1U6rCjFFC98Olu5xFU
ptgibzR3Z67FiqzNbMKEWJTR6dfQ0cftKxsIIKUN5kZlaLXGDneWDnDLkj2DAmeZ
4GNpusZx7FyXTLGKdKtEDAwX8TtGywiQ9V3BZhI8tDqmHVtfHlJ0CDA9GktPn2z9
QyyIWib8ErotF1h8RCrxzsq1psrlA/bt49207xxkJxBzp/2zPvuwhwAjYhRdzNlL
eTxw7xvNactXr45kGME8ug15XndHmNA0nMWpJV8gKnv/WK/GHkhf473RnSSUUaj3
nYTc231spJFOu8Kiqhr2RhTMVPJfOdAC/UuKVQnIkFKUPaGdVq/p88/eoLM4vi3C
kfYYGH3ZrG9Gl1FW90lbT6XBYgmkD3B+59iLMDZJKm+lGs5PpquvJvM65jVG9zBO
GiDvw0gm5Yy+vzH6ofc+jf+sfGtWZG17QAcKf6/gCCAsiR9UiHb/dtxUzfB4jPd3
2p/kuBK+MKUL07NUfWmjbjRerxlPZ99q0081aEBOOPxe5QRwf2eGT+5PmE94508i
Juxd92IVlD+Nza42nPfEbNnuX7mTzL5xXFzKbpLcrOgffg+w6j/JJpMzG00Y7q7b
dIY8I1uewAvi9yI3NUkpeeGunw15gJA5JnMZLDBztH6Tg+vQ49hWUpWkSecPdl9y
kCmGeZ1h4lF5dw0WhhTYasjSUE/f4MK54fF+Hxz10itIs2bscrcQSIF/7Hj1Yv0H
oQTXMD3GzxYuYf7zBIts2i13qvEWCryO/YFuBWVIWHPBhZXvBkIoJMbqrO1xj8nU
+ngDwsqixrx7e61FEZcTCWtnmPZU16N8T8b2N088zDZj5aywS9plpOJ64JCnPYvj
2qe3xq8ly/BysJjdk9J6JNW2qc3JsQ7FPN1kfmRDnZZa24n8KyAndd38TZXmdx1r
OBhn3UXN7hx398pUlmrAXf2GJw1T0WFrhbtLVq6utwwERaYJk2ZMDYi02C5hp6qt
oC9trPOQ1tstqqFHnMAHUQzmvfO/MsENXGh9AngRilgFU6shNGyoUToLF59V5id5
jvlkV/Urvr8p3G4cLGkpF/nYpEwEIkJOjex9MbvFm4HmzyVbZPi3nPRMZEyJ24iz
Fd/sJJ5aS/znjW0peKWWsea4m7dhiiwypPYazXCU03ZNyztoQaNnRN9tVD1tuEAl
eBuC1mZ1W+Hqjh3PsLqFtC5SNRZboCXZFFwW2OlTwc1X0oxl0TRdlmq+e5BRlO+D
wVMJqgU3IJkPoq+rBGgygbFxDOpC33DNMe7dxJxkEXtEko6Xg+iLnNwW130K7F7h
fjONkQVWFJ6fMMLhH5DSNyuIUWiKS5Zudk/Xm9adc+7luetyFgfE6FhCaMSWNLCz
BvRt9kSphLFEDTqFHNfIksehYnkpYbksXCRMYePRb90UW4VBZZbp14S+9vMQCIZD
4feo0VpRTzHvZ+m+IqoBCy6FkJTu8uiWMBEzHdPP1tPMp0UXbfJv0RE7Zhcf0NVn
hcf6tXd/LBM3/9D7bhypLqjXFMugPCChgpYvbSsuprSgyj9hUdiKUnkr7KVQ17VX
wtGTnVS3opX9DrTaMCmwZSj/w4J+3RaYxQJi5oBH3IUFc9s6+LYOq6OFrAep9y1Y
5yeLF88EnHmd1uSAnOigoPaTgzQofyuT42j2/8ZlRlb2ATjOvk39U+mUW4rly5wN
TQXqDb71l9g4IIUYuHbW4VQ+bC9dzxt6XmJ4+/xDf9Di9mVwa/fqWIK6oWfS4c49
d5+r2D+hd13o5pbtGDp90xr+ECh0g4z/DN1sZr4epIGt7+/WwMLXbHCBaGOCSjS6
M72PxwHJCjPpV4i42qems/sqL9n7cieP+hxBA1yjN0rH28YUbu4ESFPwa6Zdifwk
RYVxmBKCEpN2iOwHgbCn3lir8UuFwbTUyuq1Fd6ya2IzWjZVDLIVwTKS1Xrhao9v
pK34NKSUPziyPUoI+VrHmiCC1KfRG95MRWeDfRZ512GakRhr4Hq33lg44FF/m+Z8
/dGAcrEmjHe/d4kANhIojpwVpTJKoRVtvUUCFzX+KTvSswBUsRg9hJaFHPvvOqAr
wpkwVFrcKodRELdpSYrUf8K3/RR0JOpvaA5AcL1jQL6rx+bmMQ7QmqFpqW1j9XLF
R3hLBm4syGhNlwWDvQVPKBalN78/VQiRRgX89vzv4xH6RTWy78L+evcPc5Lcwd5J
b5oewpqNhgw3aRMVxl9KGLKteaPVZ/xAbzhVp5jJ4bF/BvvhUja5qBqWSu9qWQgE
+zPg+jYnXieC8cfaLS2kpZu/JYG5GyRYG1Kc+icnRXzVfrFfxmvWDvzEsXgzcHM3
oXH7LMHKg236rWUG0D+a4ByJ+8gjz49Dtx+XTOjj9EEsVQX7zJ0kO3lVep1W7miY
baLMk7RLhQZ9dm7Mv12ssrPCGyDaHmEPbu3MnzZyuzE5L+phyZlChAmLVeiYOr72
EWFeuJVFwWgpc9a3Qn+yeOzGFdy5HZQtVhEFe0uSl18okJM1ZAguY78i/ig7CXAl
0Ji3KcobXZm9YaG2mQRDRVdPhUtguEqFBsMSyXg7YhafELBNAXyrtR2AsTqOVHJX
ziD6OKUnaMXDvYQ3KQLd/SpTAgR3u/zgtGwdB8Ptsr9uTXi6sW/z1b5QlyHj9ft0
4v9MNbsdbVmlaJQq9xAAUFWLjf+HOFkOVwhuX3Vt+VkedR9dXMXeZNT+1iiPDyC8
GfWxYOigvJkb+zSCIkG1+peapOkPtcoSUV/iQxaQZLl8YAnnleNrMK2vRHhbQcdv
6sWEl1rw2VL3J6X60Azp+YPhAoHTY84U+Q5jwgQc/QmZPdNt4B2niTh9o60Xk6nP
sA2904Vq19ECsQ+NWhWIerXZReU+FYRmKpRpJfc5ml2MDCtrV7cgnSiyswwPDr5t
aDlfPBVqv6m/7c98PWCtQC7qROzVS3SoQx8Khx+YhmtkgCkU9+s/N14qfu0+2lzD
YGieAtWVGfBhA2e4TF2jch0a7FO6ffTlzpUBFMp5Z1T8WnIE4qcmZv9Ux6+Hjp4b
vFcgbEHfQsTvjT6c6hQoIWQ0FGCnuK+AhK5+PeZURacqx9chRfhnwL/22QUbQLcq
sryq0ks7Xpqm946HdV0UgUNxusTCm11v0SVXWFNMCE5iFoW/y32p5gz0U/bs08so
iUwNHZKyC+u160caHWZ+XbvS90AOwWBFmV76Od3Y953DLWlgiU9GiLCi1ZWAqRdP
pU/+H5mk3D0uIybrVLzAntjbx7WAnhn1kbua4X2rwHyV++ksOeGoD3dTZk18eCVu
7JjwzifmP3+x0svkWkQlwyU9HsViguRW9nsiNMEz7wVvaqnXk2yEAD4ugVx9k/it
+yyVIGS2i7mnaU3v6npIlTF+sq74RTcTdXtga0Rix23A46OjyZdeqMtlPwyzzA40
IKcvwpS8VovhUfCW5BB2AaEdfY+J2+aYmOAVm9wz9ztY3Gswasl7LiraL0n8HcEc
T30k6FCaFnwhMEjHZUeuHceLZzzy5mszMQCnPDUdWJXVQ2Gr++/ot9R9IktjJG5N
Wl59R4yUrhLtrvsWr6/IB4c0hfWXxeEuaW1c3zAAqX4AjRxw26w8obtDWT8AvMa1
bm9nkBIfslb/Hrx0CD9AG5XiBPmgU9EPlyFaPXnykYREm74o/SQW2nESNyXsigmo
ovuu1Sx43MAfIzWzMfrtX78b1ILVuZU0CHN3gzkoi6aXP994MwZPVip5+SFUZI5F
1VBCzQjQNEXmBz4NG6FYs0c9wzd42OnRDchlV3cFUS6cgJrCaX9sTxVSzro4AQaD
UJqeDRssmT4Wzpv0eYwoPpuVYN/uo1b21C7S+yggVDl+kgCpI768RNZxPy0SQl74
Zy0hdNHxpGDakeFAUfUWQd5iCaxK68FCQTeZhbYatWVjr8kkdKv+Z7SiSTuHwNFo
ErpJ+ohAyGJ6xeFv77w/kjaKREX08zwuUPobjc0pAZJZGAkc+UuRkvpOCMMJc0Ip
4LCONwdzghg76TMpgo60fOosX9nvrhSVr/7xQE8SWY+2/DFm5jGZIAFokA+7q/QV
arWXXr5IywFoaUwX8pqlHqNSxhajaCpkLV6IJrXo0EE1CepRsZ7pP68YAaIWwlUG
R9cMXKpD5qxhwccOhXjvXlopPfX6WnEiGWytMebBlcnj2ziYWdvd1JMtSdkV+5Q0
xy8EtUxkMZve+FJX3CqUozN++zan1S5CV8F0SAQY8ZbhBwMsLE3bCS4TXjbBG8Cb
A5hn4o2RJspI049pswkG0lrDbYIGgRFueByvp0U3COGBjLta1iNoWbw3BbI3ybfh
wjAnvFS4kGkkRDJPE8fi+tf39GiUDSvdIUPNbcE8vOH1uPzvr4sGzBzG68s6cl6P
RrPwbLBHu0yo3Wo6Chh6NyhKpDGdPH2x5RDFj8fOlY7AzMCNtX5pn5WEEXEZ9L/O
dhzd3xRdS7qOMOI2spwr9POv24pXnNtduA5CTqVfokEMGma9Mg1HmVQjMbLjAmX2
rqT9NACf3LI/100cAelgfDuf7CfZV0jsEHfzaLBjzRYRx4snJguFq10TTv0E1ByJ
Z8vaAN80mB4sbVzrmIbQ46tUQU1u8iycOK3Hwbk6cn+pTc79HjR6oIZ+EIoBZSGD
lh1rA8llritgOo7kCeFS+lKHcvSlOVEM376QLK8qxoC+ttbUVbfvIcAd5/cT6+JO
lh5YBsCopHy5QxUZ9W7M7qSDvh6o5iGMrwLI+UazD2lAo3p+dH9xe/VtDy60+WLi
8ve33lGyb/E4VskhbqTBYoqxKaRu9A3whOqiQe9A1DW0+5VpnePMGHkhsGxulb2q
CxLo7Km0hjx7qD7KqUwT1cjb5irgEDcJ+gaeeLM7OFuJRisvw4Guz9+sIMNQADi3
B8imDRRJhgbfrYxxAQzOvw/uFDblwKXYi7PHOWbpjrPpe9cx4gnTOmbGX4xmrrir
464mo/o0MrLGv67SkJcP062JtHWpLQzEK936d1pBdIzfIBzzZEFIoe5yo434addu
ZBqRKuO2+AF0lj1GRbqWn+YvxTU7HHpwfxjZkQNE1AdIpXIzyUIHHEuYqjiYK4yN
KvFwWrPXgFPqhxWwe5jKOsmRMEcYP5lV9qNQAuUuUqEPXrR4G9ebAf6KKHyBBtRf
mCPG97EC5my9iC1fRef40/kI4cqHJ9uL+h3dZyLnlLFFCHKXA42jPYpqMvKB0r76
gj8EAO2G1uckMtK/FkmeGk3kS5vxKhXFp4DTQCFcgMVhNvZD09OjpYKDWsBAgCK4
Foc1NsRkh4s1Mi2QywC+ds+5kn/6ZRazzI0BCOT2xHILMccr5LHOcOVEcC/Glo8N
WICgA8devWzpvA7/jZAqOyss+Ww+23jMSL8nlvxnqaT0E5NVdUkGIJ2nDEXbKPqe
M1nClFuQkAJJtgGaA/fb6wUMtVKoJ8kqNaAxPa6sqD6gN9jy3XjOlc4tvePoVmfQ
yWBug3SitUymMDlq8YUUnvAuVeieFL8lXKC3+OVt6oFrVdSne3UoeOFp70PFve2E
FXFG0nhDd1FVMAK9uSxjOJVtti9FRamuvJyPi1/UwXTkmCwU4oikG5KyCjJimXFB
SF+K9Af8Ml6wEUvZ58N4knASSWRmMpQn/dRW6ri9RrDPxf2UOfKerU42Qr1WCUKf
A27PkjgD6T2vB3sdPvNcVRrZxa9FAwr0ikrwkD3z8M4PhrV1vogCf+i0vqhGIeRK
ZEdv2O9QAU1drhKDXoL7N+Fos4uXhJp8dtNBHhxBHoClp+2JI9uO1ZO3UunvWBGT
SgumBNLmvGV0hY9N01Igg3nDEbPIzvVZnuDwspR1tGTc1qMVhsbbNH9ZjfT7NX/J
TSxcUNaCP9xiU+pKztptzwohchd7hrjhdc+V+xcsNsh3EcU9fx6hk2DDUgcAVg3V
wu0qZuEjR/8HZEq8JAfZAgnZX4ahJDIYI0ngqp+CtGoz+XnGNpavFH0r67vzeBps
q7Mk8IO6WerkPBXzgaw87e1d9zotky/OyNvuc78h9YlTbr49Ax95f8bLk1bfGSvm
GxCW4DWLxSRCItzNc4+88u/HsNERdBpPGXj+pv4m/y1HaCtU9Gy/78uKB8+8tUk9
8QiQjI5Kp0WNMAkFRzXacfqUS+vVfSgFu4gQXBObiUupfVJ59CN1Y7nht7VKaYTU
R/HvYyq/TQMxGmNlbK0eftOWGoWECu2caxZ6vEPZYxaDuVxwp2UYUVY0TIatYamq
eX8+ng3BKsyvh8hotCwZuBXtnrZya65dw/h7aIpZAsBEZp+/oZ2dmz+eNDYg52Q/
e8NVl31nIXx4VuYNKeaeGCzyviWncKgZii5kR+cR6xrTqzfwtu3A8EpwnL9Ol1Fr
ZpxUXscDg4UgMZNUIZ4KKyK1bCLXFhafMy45t4Nv0iFNPYZxHf9ZSIXiAPfkFxK3
t5oz96V1MuamOHpjbCoDLq2z7UdvwCaHTZySf5RXFIIUA8lb6gFbAq9DX/BLys+3
5roXe3H7FLONQzjiNTKBP0aJm3MWv2azc6RX1H2HjabCdBgDPGHZgiTdVj1SzmMU
Z76jXzHxBlfERxhiqlro9GP+w6Wlk1oq+X7xt/TGOEBkGO6NgJXjCK9zZxUPEr02
hj8vxMz5LQhMz4g2Ctl594e6vhTUn8+taPmxzUFO3Zw3mDIHKAfSvOCGCjErry8I
p6hJl+DA1uRhGes2dnRYQwUsMuN6qERWol0/EPclACYe3hKs/AMTq2pXPDi0PW6U
naXMj4NT38Z9WMsKnn3wZ9NJpHl6FCiTHV9VSFw8Hd8RQaPcfDiFjwxOUsspN4G1
9y4Z7idWElf+29P/pRIVo0nkGY9mJS8VQtP+F5hrWyi1ASKFFRzg2TAKx9GO735p
FKA/k+ErPzZM4ny0wF15hv6mU5SzvtmHNQwuiuASXQyYWkMOKsmNBOu9r21QYq/A
vqh+Lsi+I4XfkPsaRlQJ6dEqP7A/H9Ju/UaR2PcdHmuKUvvCkUw63g3/0mkB1X+b
gPB0dzXFCwTNTSGqJNx2BrSsJ7uDtLPSfovDWCJf3D1IV6N3RptDmj3x8092w6yO
TLLFlWFv3HioLzCxRnP1DqoH7FcEDtVoCbPhksagj6Ck/F9l4+za0Nyg01KIFCMB
bFQGJOfvEi5cwTGMn6shKdeHuywXeGtHG7dqJiR5mJTCVFi5koAAy1yvHyzX2SS5
Gwse6N6obvVX1WQEtc80yxyvBL45I1k7x91y6WbEo/V79P2/awqSLcCHzTf7kuGK
IRtHLypewUuduocXpIJSkxBkRwVR6X4hl7ZeacSNz+N+rivNzdAUQdINEds5WDqJ
vnrEvarg00wVrIgRMfv9zeEXAXQRG7Y/1y2UyI94Ma1hdnPOFrBttD1q+pFeLlFZ
CwR630xyt7JUNre53Hn2q6R5Ra4qKN0svB2Hiz7Xn/SwOEhfA+q05mez0rxZ9oYi
8VrDS/wa8ICYw3CsbE9JnNZrSAz5zWHf8WSFBoR+BXowXG+06R2W/tYCMbQZ5xFY
m0n18I5Nccyb+D9+qO4MivTP3J9dDuDfouyRgmT9SBPhjIPowMAhqBcuCmHfU+SF
nXfuw7aWyfR8bIytDT0rtZvqVbPFQgkbw0Kv0nJrDHCHi4jTyapxVujAbAjYaG2j
LuYRVEGJkLCpS+0o7MuvJrvcg4Jh58SwaxHAoYS86wwpKF4QCVdaGvBYzlT8Ii2U
TEkSfFjPMf18T16kAM5IsQoL/IZ7Mz99N+TV9WU7bvFzq/UbR0nyGeaKXelWOi8g
mkxRmP/7WaPE6WBqzMwmfNiqAmwjYOmkCoDQzSsxBaASlAfdNnneLvTVilfh8oq0
n5BR6+Hd+9WZaHU93KaHLNzdqemrhKplan65goXQdh8a2RpB0HGUNAD76khaDpAL
h43YwiMN04tSottjsLRvNN3XD3MUVVpWpX+n6tEa+VkmKXK2QzS50NcCRae27/RX
ziKJliTlIZprYQjbUWpxjjTJekZUrYuK0sEyXD4eRZLO6Wq0fyxD02rEOF8KbP1s
JjZ4s3PEJSu4QXjnf1T6fJJpFsSPccYB+2PPZHlaOIC0NoKwU8uf8VstpnazbriO
z7Uf6etrlYvZDmwgeoLjtDe2LwzoDO5DmGowhY9XlquCRSwc+6iOX77HrNRbBmCA
AOiLg8DHraFVXAUzvcoJ1hYmG9t7z3uamrdFaRe8lccxzrDIjKTyh8U7GsPgfi+o
stO32YggzF5gMo7Tc0gJyzfvjow4D52HhqFHNIAee4IAwSDc4KWUWQhwhVKR/zTz
sWIdeHtIkV9lGhHZcgk8HapDtPk5dD5s1joJp7t9C/fnhxuzOvM/2DLsC36A3XYK
m4d3L+BRoNKj+PW9pkGFSwh/qYCoo+hjRceZyH8RvvOqNDCVinBnTXa+eKZplJ0N
kBrIiE31Yx1oMSYzhFDwQFV9EY9qoKbV1MZcBIkEknIjthH77h3vhb1jyZ6UcX/z
/7eRkp89GIkayZEQrOLLyX4aGN7e4fQLwwDJZ4Zb3WasVmWuSb8gtf1j8LipRzhb
2lrVEz+0k7MvY+vHJyanDUly2APxeId0x/dRdS/qDvvWEDgbSqaJLqpDVJofWLXv
a/LOTMBohm/5VH5x9py1h3oUr3Vt5R+zpb/clnrjrmUA7gw+IysdozktuDs2uQar
lA+3LgsagY90NSWRxh+AHZMh3OIMJ36Wc9agp16mNu0xD3NgkNpTyJLtJ4eK4tST
m5jTk36RGQ5OPw60+BmdxIWYsrwHFWC3HC2APXJnO66kpz75TZsMNzOukFaMSqAb
1GFaLMWlc9UJI0kLNluzjRsZnka9ZqEjYhuKbuENbZI6Nc+QKf6pYan0qT9qFejj
3IOWWONJtB7sZELD0I/5jvcxl1Km2uuy4UuAtfmmEJ+hDGp0iE2IQY2QxRA0gB5t
fw2smpW2N9BFzVXZL2RLkueW7Pd9/cmN6S7VuA37Mavj7H+Uws9gHq4WRSTjmpHf
Ev2h3g8NfiPWL85ZJ+CG7CSaun2a7KeYrmgqb8iPSkMWcYiw6kTBkJoUJMfFw31R
jf1Xgl2u55e0+W2zOXj16b2ikdyx4OMsvDI3PjeTctoC7Q+H2DkBoFk6mfjfoGO4
QuWt0DmH37YEMKzsCnAFce8a5L3vrzw8JRw9j/fZOPdJCsFMutyoGRROvIdvGCgn
/xKmFYL9SutwAfdzKIDeJ6dqAvwax3KEJ4eJsmhKK/mhpb7jIOO+5+johAIqXNlC
TEp8oMWeoZ1N3qCl0frKp3/tPfAE7at52u6e/WGmQ+zQI2oWd26PmnjlQgR82jLu
Pcc/CFDoLQOZxh8NRHGg88EZGWOXWnSfEnvmmeEiqj67B/7baZuIZ7AhJopoBjAd
M+1fvAmDYeCxHAhKIlMUmbV7qRpoQ4jN2eiMgSGcF6jBT3kc7mJ1QQ/SW8di0SqU
rmPtXe/iS3BqA176M6JYdDtBj8p8jQt0PnL85L8Z7Letx6+mPSxZPorIceTmUJjA
6asq5AA6oVQPhkqOdG1p5znJMLYmtfeUYNdbToDCIWuD+ZaTBalZ21chHeXizGDf
5wQ50BdEzV5789y1emH/9UWFNT9xpz9quHWAijqrdH9UAVu+gFJHyB5bO+O6fE/L
sG0My6m2KPnxaDrRjGgNRf/izDhTsiRUVxYwNJY+NBX99P3CV9boQX6OTgOkQch8
hGTP6sWGegH+TQ1syS0twMDVYTlSuXMffM03VhxcsjyFsOzk1KuzS8QYxNQd3RB6
y+BoTagY6dBhnM0SXWRyMvtolg1yH18hzls36aXexZSt4Sw26CPpB9XOa3uZxrAr
fStry5c9Y57md11HKXXepOe3pq3byWKcaKA72rIlIVMk//ynly1OS9G2yDCmbjHC
Ekt4UFBQAK4j1zfsyhoLFPGoYpqxIik83/nlmRzn/Fvvp6/LS848szxeQoTlw5g1
TVuGVUANynxAy9CnzxOJog7W0CAEsroqzrNt+QngLRFwqfi0fCxgraC9MnXebcgy
Ix5qyRgRpKdIJg8HZQkI29x/B0G/JTgnOwg7YVZv5+fhahzMtmLTIXbq2D4PntJh
JD0RyQOYKyoVsxX/1QkQ7BN3im/CyAK4S7p6xkOYHssxnxjFhdrkzrAvOTVsPYmv
8XVqC5JhoyQf+/IfISn0wctgVtDJp2JD1doQYDrzP5jRXFgBp3+MXS43hM8XMRYP
N97Y/x6H8JOiqgqnXku3+++kfjb8Ia/2UGnmu2simIi3cCmuNA7d3z8rdogOgSe1
Fvzv5hJzqn7YpkfMuXMZyFUSXl2KHIShPlhlHFvo7qREXIvG0EwZAU8eLyxg/wr+
Te9ikPC+Cxszx63vlsLzFy8GBHkMCH8HBqkRFnCPEr8K+KrlOdBBIPlcG5Jr3ef5
Dd9gjrPX2lRlOFf4OqWp9R1pzXQUmDVhvH4XP5PI6cJI31C445+jX5dkFbQlmAx8
r+Zt4dFBE7OjAoflSo6OlhJ1/w4l78ZJCXVZEG/gWKVIaz81fh5l2dyuwS6fLlh3
eP6gavrx0SgRksbYr7F2BKg+c0ULpMpU/gFDUDfOKx3TXq4fTdgkF1bVSJMJ1C/l
hEQK8N4NvhDRi9efjmIfzted2PKRSUABjYOIfNWJy6uHzjWVnjk6NQAumxUGarEI
2e64cId96pcElPYAS3tIQA49FEoWHe1WDPPjUT4sIf1/f4ZL5qgpvqiW6nK/Hy2S
+1+srLTcECPw0wlYauavFsTUAQUU/k41fw8Ome0u5tgZGl9vGkEF80rZFYuD0LhV
AbCVNBcAcZeQdG2JpbSBnZEVDc+KEe3RA192LgF5F2dePgWrONuUrfg61DAjk77H
8/mOfATEMfqdVRk28+5dKi7MYXJUzb8+O9ud5ZWRHzBV172oJeJdmqUUK+ABt+A8
4wpQdiy0kni9JAx3cX1FOleUARnW6ZJOivBdxlnyPQm+uRAlrO7hNBy3Ih+4RzyR
tJEk1FLtzS40caQFhYjcJRj0ux0bfowyGv2YS1KJXeex9Pg0/w8i1vLyZCZZEgEL
BDtWga+tH/ktZD8HQfr+c1ubTS3pRkyx9ARAQvuQGUcyw2NYEQciXTfTWOmUwzIR
QC2LCZhTSQoNe8w6TlfDWAstUH4bITehTOIfxSPIsoglai+0LBIr7lSroRd23i8n
gv7k/dSGPnhpmoWwDb1qQIAQr5Ak6fiBYWuWGcVnf7foU3tfFuYdqg48ENgzPSNO
lTXDo/L8weqFCEMwIW7ZyyObooUnxPp9PshSXbjyLX1Iek+qzZxWeY3e8WBj/Dx8
VADt/s82R3ZsIR90d1ALkGFPRfGAA72ytyVGPebw4fM3iAtKjItLUubJz19SrPq6
YPii4Ekyv7VNkfm7Na+pAEGuNiySPBgFjajbP29Q1StPh2LE49yJFXOrds0sFmAb
KK6E3EZ26POLw74z1ph1B2wjTy9WTJvoNtNZZ4/FcVzhvADih17rXMx2g+4DMtAH
nyIW59ljWDYbotdKoIXp9tN0C5CWH/xfaTMYpLsw+VM6Y/rzEMi86sha7F6hXg0d
4+hLVnylG0+Qa7wSdu2xZ51Q6Sin3XgITTOsSDmQVFPZ+2IakvKqCUyt8Kd108lY
g08Ydt/iLMaH27J1GT0MfApNhePWp6swBb+vV6rk0sJUskSMVlr/dg65lAIm1Y+9
GqNCTur1Vq8wUKBJUewnEE0I9em0OkzPjND39l7nKG6oSnIAyDU8FkKLcgUdngKJ
1qh/lGNrM0M3VM9XjKPQ09aP5Or/t6uaqaR/TK4s+o+YtUtsp0Fi41z2GuxDfNT2
etQL2ehbqVCM5nKHyl0Ew6sf6/bchHf3dJ0sovmn8Y46XEVSFCJQiQsnGpXXJ8lS
87E+2rraj4KO0ovlQlVtrhbyhppxisBu3W+bZN4ssKVS+hNA3a7xEw7L7KFKNXHL
/4/QvKWVPO0my9d+LTzyISVF8FmdE0Xr2E/1rlD/iw+wUm4Quhg1nfjAZlRfYB4/
LT0Knf2htyMr1iR8zgx4Hwzqt8VvqtRe+a2iv/TWZs1cy68HIj8icPefINyad9FA
7l0D0Tf/GgH1oEHemVDufZBLbxEPFZYpkCCA+irPn/j8qd7eCRSUhrT4fOLAwpHm
5mIpk+X9QgvKPLDuAIZGKLYNBgH+ju0qjalcnggFrK0GtIZjfXQ1Qe7qQWhpEJ2w
rOBoOdtRm1Nvx9/oGT/0bP6hLDVWKzx6+oosBP2WmiYb+EmpRuJaDkUWiY33E5/X
JanbwofS2vWdlXZ6I+hWn7kA1T8ThZmTysAqY+bRDk0Jjoogo/igP01Sr2lBv9az
OCpV2bAEXTDmPFXPLtNmz142Ri+auwahu3AOiiAXhWGQ8RbeCClK9ChK9dKnRc4x
o6OnvaetDKMQz5yzL8yJlpb+yjhygGsib2+hjrQmhccXlbUd+LJv/9zeVPza0Sey
R/typiP6OrulnSB7XlIAAeo0XyDHr9fDMgGxhxXPi0q1BcO1JPEwOmdQHz+cjk9c
ruhHIar/cPyNRBOU7CezTcjgGtX5QAWqmp0W9qm5iGG7Yi5Nqu0U8l/A32fIdQCc
a3FUx/BC5wNwhlhQ1jd7nMWb8YLNvruGU/woHgGcDpFA2KwVqSuJ4Tjx4ejblcTb
+mevPAG8/twjgBMoVqZbMqdHdVXfF253+3uY5JqenXuqgfMS9MPfYyANQ5sOhfi/
L/WrVnq+IPI3Z9oKboT8seyA+33N40r61lZ0pHM1jQoo52DRjDEugZGwXUnRfPNB
08tlRua6rRb3AsxfKV+ywa/b9A6rz+cKuaHxUphqfYxHaHldzc+rvuZBpruRH3wm
yh/Qxn1DG+qP1HOe10HnHRUGATBVr5WDBHmRxdGpyRK7bEAqfGsVXR+fI0Zjr8tk
um1lGpY+1ME/Wd/K4WqlZ4YelfYvdgen5qMEbcMGUk5r+Hp1z1Ikfyjv4dq5Wrhi
1etbsenINQYYc08OZEo4NKs6nvpkVkKkM9pkpuY9y7CFcux1+egKsTu1LhFBLu6n
yYzXlhQhhMJ9ctZGQCLipuWmyJueegW9H6JOGsTIg5q5pbGwWN0CbqdALgomlMrB
6Odje7XS6WfUEKoEfQ2tMOf6RnVCCnMlIXnk/qs6VaVoweRaQk9GgFuHrI7xnFmq
Z+eJ3s0/Z70sIjW/JvlDU1dgjOLcr9IPklxBmslFjG9KzI9a2hFOnNDwaH2yali6
yvxAYIKJUJ6BLAd0n7qZajk7WRexl09u0Il+yd6C5D2DsdSwj2WuQQjElyz+UbL0
IXB/16S5DIRO3l8xmW9gg27t+e5+8UHRtUYkI8Bc/C16F2B0/6hptAwzpZs1Z7KO
Jzqp9QSnnjAm0Ib9H5NTinZAa/xlCCoQGaO4wbrflMDjan/cE4BLjd3zpmWxY68Y
fRuiXhsRgl2EVKc8N4qwVHxfBu4bNvoq3RY0fN+mcEQle1XKJbcymxVyGzVEzI/r
IELq16JVIqI74ZgPMW1b69j3c6mQFPx9Hii6ilGGDMxw+dl5CvMbkLHZ9vmB/L2l
3Tf4j3AzEAckc6i1HaMxQRQ5EOGNupHfiTCzilMGPr7Teum21/FDRUMHMyPUZ0v+
O2alNiI/eKyIA0nuFfLE+BxV0lC0JS7TqWVgrI4EqNI/ksVyElaV5Tt92A2dqoAm
NNn9NXrmAm6I4nGQZAN2jxlhkdyhvaSZAihQISoVZ5znwLwfmCF3vMcEDXBvWeuC
bBuYWIjK/vu8drUBjgiGfBsoyrCCvGdopbu1Pth7zc1pDenL1ouPdW6SaqFKlF7a
cpqomdKc8Gu7GsyvXvMBNe3mIBoxq4CP/wuWwkO757XI3u+wBnErYu+Uk1c7XrKZ
vh9QqR5f+oCbRFoEP+KFhWxRoLh5hwXsVdFw9MZEy6xtCAXIN5Gf7px2x8BnHuUY
xK8KL6lQVTJR7K1eAi/cweDK533wvnF7vIt1HFf1ZtowIglFHikmexn6Vp7GCVLe
4jLOE5+FpWQfC83fXs6mLdYh4pqTpWMcY/DTgop+rpsVMAqKAVjaYX30xIClZiS1
36lv9zEdPU/zuMDB3vbWuK6HJlN2slrJmdRwPbf7fvjLEM382/qAjJiejiqG6YtL
eDwe50NO4xdw8upzYICvS5tRrjV5L9AgAPJkGz75Rih/ZG5fTaCrcxsTqhdNAneT
qu7veUwqdO23V/zk+euJNLrmpq5CHylN59bro4vqQOM1chfnzINWp2yTH4H55+CH
/vdQPqYiszVf4yPtnnizuRtVGm5gmnMqy1KjkqmJ18v0ncz4BZuvcamMY1eeEbQ2
CEZf1I1ECphodhbM0Q/cmHY2lH8O6wWXsWm94GaLHbajsPw9g20FGOxce0EEK2Ti
78GZVdoAnhNKP8ULWIW0duBU4cvwgQ1ZI2OEWW9RgKeziwkBkrC9/n98ezpL+3YT
2ZorlulUUgv9CmjdxKMlAPLmv2FNRCMU6Gp4tKmQySci0hnxmcSglsXfes2xb1zb
9nWwbR/aC3CW1w+27zd+KLMaUXRo+tjfYBcTaLEIhKYCdyGe7IF7bzvTrxwYzqCN
PmKQbNSo8YUj1egE+ae7HBtCIsD8H+VpUajx66CYmoWA0ee3B9+W2ot3qsWm+zbL
4LsxybBjIbQXLnwv86gj0pogBFxccZUksRsS/Va/5XnTuNgW32tiMbueH13h+HjA
+0kwlVPmHfNY36D3o7tzdKDicmt1dd2tKewYQHLrsqFNKpN0dlwEKD/dI3Vi/qTd
mgj17CMm6obzRkvb/H1N6ftQEudIIu+z2r1pPTcwKw1R9ThNzE8cyqTpSM8pkGDF
965pO4BmKZGkF6GOLE0vqRIdtfrky8MWInuSYnKBSGtdVEG/9RwXgP7Q9zDyzjbq
WeMggDedO49ULDWfo/iG/qTXzgLX9ZtNBwYrzM9xmPgWMeCVgWtpmdx/nMKSrh/O
PY6z3HmQktn70tpUfQaToYhcNpBo2suVGqlbVT/ovCVNlhPv+n7ayS2j4RL9gJOI
S85uwsO6Jf8Uri8C12QEeljz8oHSZynAGcv23lfGTVQXNl20DPl4gFqIEcV7jhnM
DRCFZOKiX8si/z3TGRkp6JLohTXY3salQnsBfbRf8q4inx4UoFUvJ3XCj/RYOuLO
iSRecpIdxp+0JI3qKNLklAKCVAHG4Y6sK7xa4p15bqv0Cp/rGAh3owG9ZKajO+3C
zGtLwmu+ZjPUaV5QlnWZToO6++6lSfQz+dL+0o7A1T/VnRQImGHET2XvIsTElDHi
7W7jVzRvjONUj92V59pkzJftGYOsMhoB4zVd2hwxiVbjkihC7GsTLwEaswvPknwF
96fZdFeJkcRYleyg6TEMRDc3eie0bYBxAPPwucEIg/ft9RAWLg0VuLLkpv/v3RAw
PisHXPd0LuXEWwoyJYUIXghUiBqQCOg5Sg1EUV+0PKxlpBM3w64q/ULdyyzuTGbT
p59OA9a2DGdcndoXDrqfkoPm9l8F60wRxx0FyWEjEAxYNsWht7SQsY+UhogX4D6q
j6/URmMXKHXdFoUsyK/hYyHPr5j7SKj8N672u1L+QgmmLQBHgZLT/IFPXMPpG1oc
Jw8qh3h0PdPLUFI7AyNT3gTHQW62YutI0eBgFWOicdyi/uTs7GxnRs4iBkpxC+4g
bc/MmE4gKw6kfn1GcpjYzG6GVcNUqSgfBq6yFesqY0rNnkgg5kQesFvepjFCHs9y
wHOYFUMGqMzEcVDadab4Nh+T06rMJvhmfsfOfFUIi1UyhN7wHDtJSQiJl1Yre/5p
Takk1kd4lrfX3Hdyf+yc2yIviOiDECknXGZbVtkY1dJgqVrhWa+Gk7HknaTOpVaz
/5ddc4L0b8hudYWAF4KCXB8sfFz+h4dNN7d+IYDN4suoMVFWpSPQq8DMG3l45hoJ
ET0tGS4pxIToe3RSwYwXxFMxHgvo6xiqzG/SHcPNodUYusl0y8dLtKcF0SNneg+1
ksrTanb6DZ0W+Ndrd/bMM3Ux2v8XbYrc7ru1lGTEVJwMfWncpLDFcE0H4gIC4j3Z
1xT5MK4csruS5K93PTDsEDXgSKbHfOzg5hzpxKbceMaIB0J0q6E1J2MVh4RnvB6I
oL4hYYyrSVobP+ClUpFAspDZyQXujFTBbEAgcuV7FNfvQvfBtzkTzxSvSiL/wHmv
fCMLxAbRJOhhb+F6z89PnrL3a2S5jNAFPkINYoSqbbGwgHEajf2WdbLHkTEAu/sD
XKg/sKZ9OHhEAryc0jjm+8ax1XMPOBO0Pm93DMWASdxVlayF672DPfBYRVZGDVn3
LElTD1f3LqB7J0TxqtXKNjhxDoSeH31kY7+/gxwobxYyNKN+uUiGspTdDTSVbm7/
+qW+aj1PHnCsBAREwRYWvo4mLW8h12uHWeD6enT79k2PWKSaMTmiFZEVf+9vtmEc
2KysUC2pT2ujnt59HN69pZjyp86YW5tZEZQO8ONfU/fKGjzzD+Z9Nj0ruwPIUnue
dObQY+McTHHaWTGeciZlkkEEietGvgbuohdJEiRNAnZH5uwCmsB7VWJWbZRHiMzw
IvaB/A/lGZ0ecT7M1FVz2n8jfJ6dXxFZ52pX2/Fe1KPCZYpEL9N53omXhY7BM9y5
vn9Cxxi/qPuiG8LzycjiZhDpOvzAs5B83bDLCcY3MUdRNOUhX9KT0POIJWnQPp/u
umd5mrMZ42Bx0g8spFpPNMvcTBaVdir40FAFKAiIbK3wtC4eW9aDdKLY8hzL/pFi
zZOPGbRtw71auf1shZtTQb2V8GzPjmMB3dCuDwYKnIcGkWEnVfmbCWZ6KrV/LVjD
MFZMHTf6JZQxiysu4m0MrrNGZrVHAcG8kCr9KVGAbnj/DAnfN+E9M1jB7otW+ikI
qnSdoJ2kPg5k8SRM7li0Z5pE+6XZxKWnCFaR/TpLesTR0TqxOxfVDpjzSOFnh2N3
iX4r1jWZct/qcsOPtqpOd6Id8CIBAiHSo/2sLwPD8oSwpOXw5jadT7SwAX2gy74f
+FkTouHRb0zaPcdizRbrRmS2dbE9oNn2N2+xi7yb6ijOJPdWNbbkuNakmoe8Uxg/
HBg3lnNSH8gQ57MypIV5E8k/GOQE/6iht+cPVt47+6RFVm1OeT39f5PfWPDx8j7S
FMJLHSgbJxef+yvMOpEO1Vl/+ngoWIO7AFcdel/SVnfBHhociQhqT6Q+XtYxYuXH
eT+P1vEwKsbzUr1+HA8FebyIfhn77wKgUhwOIYQOAVz976PgKlGY5jtUo5Sk61jk
gCvOjEre5ufJcUrBdhrnG06rP0LsXpy1X7DWHGHwMur+qxjwQgUtMnfZ4B67vXHa
Hb4I5Mp+vYyB41u54E914T+sjdYCAlMfaP5disvcWSAclBQCKeTSxbPH8A78QcDU
2wwMnL7hWsOClZxUW8cpRGYQYrwPH4HlSnYbJfLLParNfe1D3u2R5pq90PKAUpDF
4Iikkxzf41/bLFAQWSaA1LbWxpVqQDf+2CN8nfyZgBuwvi5gs8qrTKPR/W70s+OU
rrkubwhKMs7lRJyrkHkPMQ92dJSBtE3lg8h44Tfqrz5KsHAx9ZubGlPsjCy/V6UW
pSKV0cECkZpY8oAAI5zehc9Hr17Q/ARAf5ZowFjs7MXcWHWN9hi16c4qisBXfhGS
1GwJKAUvtGJCOUrHQJx4BB9BgrT0wJp2zpaOyvZ4eLmSKpcPx54WzENT4fLN32sb
h3JDjsMCUdqRSzagMa5fLPNeaTZ2UxmpYWbPZMmadGQied0k/A+Gzi6q7HCxRkVM
eG38HXm+IEsp1B8ya9yItry+O8Kyzgyd9Fj7NHI58XfKnN1bEdJ7GDggXbOh5P8V
8rmn1arF8g0a827ECSpoJNiI1pxzJIrdloWK1sgeEWBnwFfmg3lCRWCF1N26auYM
HLWd3PXGPW/rrvUg1CXGj7Cu00ixQEBwHEKzuHn6PmZSnphbv7cuX5LRUtpct0Ow
NWQbevQuBlG5vgypNJWoLz9Us7H+qZbGBk+jY/hsySjK8iNS/91ndB+Mi0s01SVC
Rto9cxtlW4a6BvQxirTB0ErDwrjykKQO4RWUpf3syAL56UxR3uQkDjH9weKL6sKk
NC3Mjx4dyeyLHVz9V2OLzWfgeyOH5Q+gAmA+VKWNW733OWTs3FszJI9idSz4CaHJ
n9OBt2pFrWdJBLwEJbXI/cNjve9lz9c2F2I7ZEdSbJtdtnT3XTXCkTaMtxjWeQAk
zMGcNJ9bzoUy/TsDNmOAbeymdH62zCFHSPxMSNzRTj+kwWzOAwLBcjZxX2Xy0TLe
Dt5AGZqdrALCetDqKjbgo/3QyRlsAMatH5C34xkCA+iSUUhv3mfBtmOXyb24LufB
0mXvbOZke3tvN10srEEfHgOOQEexnLconX0Qx1A0+UKfKstRdWFZR+83Z+vWw8Wg
ztlBZVMl6f5bcVzGA5VuNuTc+MjNOcDq+25WQG572E/2QuuxIic0k6FUG0qgQbpv
W2K3Np7e5uiNmse+uydpJlkjj19HEGrg3uBeThrEckVrXUdEvU9gCBrCPKcZbQ9o
q7+aenadG13l7an0lcxqG9AHSJEVkgkMzI+DrmnhhyMffAIlIzA5ta0T4XHXPgsU
5TtfsmiTNUOUqVyYmgKTeox5YE/KHfS7BPdVkknWo+s1lq32W+43pvfz+9vWtXMR
1AjM2zFzvwJd0s3uOazYRwToZAxeuJKRD5IR09W7g3PdLshFzO+33H+I/MtfSP64
7tC0Fk6TQbxNqxguNrjNgU5b9YHMHIeuj5UMtJ/bdtNZhaYvzkuCWasWzdmp3XSQ
RN3BhXcIUadl3QdytyD7AbVHUwgMkVrK+rny9D4eSWnC4X5LK9xluF+SDMaNf83b
wR/nssd6NWcThr8ttYNRpf2tsOjQVNyHUqsZoqh3PwWN9nZBNp4hktEN6UPyGO2O
AMJg9BHTT66elttbDrbWxojl9LMSWP7Rlyib5uDh1w6xlpX9blsTOESM5AlmkYPT
IXG0/T07ERliOO2BLrTrHrtWaJrdblGmpS8a5ddvhWkBN9Bfm9X4LYPGZcwQIQEH
ZfdQcdeDF7nY4cqqKFjSmuZ+r3hy54/9T66aVU7lB3KQe5dO1Yo17BHvkJUGok0p
4Q+ONqCyTkfuDX4ufoA53Npnqubxgl2NaJqQCUuuQfK2twNkTMVTGA7ay1wXrI4n
gWBufA5zhS4Ku730iVS3Cgy9IoyvEtBsIYZwJ7e1w9FM9jAeSdyQEtMY89JpnpR6
Dih+T7Gt6CbSOLZlv+uD47exE0JDLznMWLExBAwva0XL7dRXNiwuDLD9vFY5PglD
K8EjBaj+LCO5xYCFJ98j5k8w0WmMsVAfkrr3oHwKJhaOFcr9RHPKJd9v1nMFjNzV
czV+so59UjmI4TZIPvtjav5iMZ+Z4ilaWn/CjvqWYoSgs3rw/VRXRdDN11Onlimr
984UFK2v6Sx7P9Ql04TCWXTy8PoRCTbp3oRZT2YU9F0wrFt5XLebmF6Y4cqKKkCZ
z6oD5W8ZcRwnkWHcEYkgDfno1YfTueCWiHdm5Qy9c+qw9AZS8MOHEgqjnhPVa1+h
VTfWDD1MlBlp1dFsxstFP+kJjaPrXKKjs7v4iZhJ6jMBbsn+PtNt/XzcC5adRDhF
Kn4AfJ1cBEwn+egilVbqFm203GRZKMCn6njFvAqXXtO482JQtuxDEX+oN/l1mdBm
OqPyhVK3tQgXxYDBh0KwFqHMi91atN2ODyuBXG7uWhN9Iw/krwDHcpWLM75ukIQa
tf/0cbqQdF1F2hMyyxYeUe4sOA1KQoDGo54FFPv5ttBu8Q2yIrzxASvJ4Qynewdn
iDV8nSeVkGugQXKVTWrtd03C1ra6c7O30XISb84IdRfoPzwnOF6TLdN2U6Mc2i4o
9t/D2hzXafLDp1TnwYHIHEXtVvUQO/rwpZvAwAN+PGvxqeOs5OAbYdP7mMHM7pe6
W3+YvS2lHkUuVYt6Gtr3c5S9G0gsakQjYlYuOKhhjJexS8VIgxcC7SUA8QrLJaUZ
9lcGzRD9gY0QCLlVjn8uLXGGqGCrSj5vsaVXwh7HMQtKoEScAt+xS7QcbHYag1fM
ogGTtmIFgl7lXtU1SehgJEZFxm2wciDKq34jdFbRILW5UJqXC7eGH/bZZx+Bh4ZB
9SCg80K/4WM97HWRAhIkoNCBMRB1B1DulC1a8ooriLhYV89aBYj/HgFrZx1EJvlG
FTlPTwQ+86t80rGrpzAXmCRhu2RTDGYOMDBN0cIAkh69nhpZGVO+RAYWhpSJbHG2
5LX3Qpf07zxvQHMH0u9qh/8hUvVU4uzEfq3d05GbIejC+t9CanANTsWBOSK6wsIM
DBZXWXj3XqLWAEx9yYGPoaPIZqFnXnS2el5cz+dAPF7xRe3kS4eOE/UHwcE4TLoq
gC0gY0ZJnvGyHDemtBGwc6iowx9hOHiCHs0Tf47u5UfBHk3oCnHAffnIn+oK/hba
bKbn08IyD7q8MRRCazDAswkhyK+R4EN+eGm9uooLmtOfYBZFpsuj3tW6ipPcppuQ
pAEoCi2GuIKq4+ToPKvCXyJL+9TsY5sB+vK7P7EV45aIsIrtPHDPkOCammXs5wA2
iC+f3UpWFtsfLmJ+P5Qk0WMwaFjncc0aGwvjqOYYTcRijA5nkDcD13gIdWTfekce
zJrtpB5FqLb0/va5lp1/uBfaPxEnAsHnuF6nQW+WS+84E0bctig2K2TuZBUIvEMe
7zI2nEDK9s1tNjKKQGvpJA5ol6PmNeZBt7kXJsZwjqnLstgG6gqwdNaBXOcxpK2w
0YnLwlQ5WmDcEZLSW39CVoXP3dHxw/0n+FZX4VwXNC3O6Thm7FcjujDn7HRrxZN7
qG2LS3bb2Zc9kCgia9/4MBz6y7vZmRPECp50+UwOOZRp+jVmdZ431PjFjCRDatOB
82Q6VHOdDW76/rvAxzLTpL8iz6G6YGBBwAas0tNc5DQl6jJnESzT6V+aXkV5aHlu
NfxK+0aRbSq8Eu3Ow/zJOs8bE1F8+Le/TmsgMrjsRMk1vo17Gvbz1U07xjuBN1zM
f7/msnidBvYCQBp2afBT5svjPN/X85C/hsrxUn9jGKDrVG1UrZdGVWvHpCDdaNkS
4bxnZmP63UKL8D1uRaorKYj/S9cUIzj1CdaYbxORd3TeOeuN5ChMUD4WWaZXncTQ
VFpBvd89LGachLrHk/ulCxSkz95EdkE6EmQDs2gFHYoju+XDLAw/HEWlcnel2ycm
OhvMeOLDg0nvyLRoiD6Tx6uaKh0FlMYp888FNkZ2ueHLEPaqdaBhg88yzjc98wqM
3xvwcLVQ4rGNZbq7/9EeDb+xz6x/jY9AOFWyd+mf69E4hQzh+H7latvQHbK+18eA
ZN6M0xS9sC4FGMgTOnFoleQ3b/xOU5UKy7kt3dVyKaEULNT9+FfATz+qcG75Nfs7
K8nrSLnhIotzpADSN8Z6Qfw/B1atv6Q6wcASY13P3HRuRMfkL3w1I+OZaStjSh/N
fUNrEtLrPMPrqYqJ8kj9SXGKvV2cVCjiHahuuTc3mLHETpBLiszVoOpQ8FuzfWN9
/TNluQr3UcZXFcUneD8hX5PDDJKCtTQcurZe5VgmT110hWwjQIOjJQQtoydaze1k
4M4DBiXqVFTAPy+VAiBstjY1p4TbiTNCBV3DePJlpexQ51kc/KMr4hnEEFe0M/2n
0keBCSEufs1bqK74A4drPXxqstYb1EDyHNdrs3UsP3ehD/l3jxNkqPv9fwzZxrGm
0nSBvOvzSQPFJ3k+AFuMb9Ww/w/ZXTkrUCwOlCoan/LfpAep4Ua1DHCMWxz8VsIX
P1cVc4uunAK1HGeqlBStlU8/cWjtgnBxY/7UUK9YcWfwptFpOkPld/xyhhFmMCnq
KTLuzL28PcgsdZWH20hFDvaE0mwebLBZIXakfKh3iTi3ofl4G9RVrYj3mxrijqEU
GZlhWtkykIvdSWZ5dRsiFCj04Eela4wiQbuxdXvUThwurxw17FuzcJjIgLoDUIBC
AsQ1MQPNxL/nGRRzBiem1Ez64v0bMkjmL3sqsZiXv9oJD8t0MeDAiHhaviLOG9Y/
hytYhlTEa0aR0M4LMKwSnBKHIfp0dMrhWFNu6UjaK/WsSfUW3mgInuBquy9mcBcE
sKjuei2VK06on+fjQbJ/HZsfeRb5JEQtd46gYclU0R34zDMxt09c7ghs+Z0ZFcza
aGJ55ER2yqmBs4TsfiVnaF5NOQeJqwTyXXViRCAbDdpEuATHHkbtRYsNsnvQqRg1
c15jYB/JrCog7PeS9+ATfEanzB/6qrXOKzTXrJO1NdjHsCdeLKun868HqVqGsXLu
xhymZW/tyexdzti/p5Ks4x7lMEy6yi7n4W8p4x5BNztvumNxVzyfqwjFSrbiJb00
2N1pfCdxJudQIeoeQFmF0il8K5YR20KdnzQkPMKEJqw6aEAoZtIlKS66sIF388L0
tPINtIsvxxeQzPD1rBp25sjwsFS5S7guZi1+9tldoNwYkL3qad88PnLBaHEgqz+f
EDG40rhKQOFWYRVnxYzKmUKFAw0CQo8xWhqw5LLdb1a1aiWVws+EyCtynRAM2qPW
v5AIh91C0rmeFrvF8PFldAn8xmYrizpe+GNPjvT7H1Ets8/YMKPbT4/AHkfYDoUH
adRUXgYbsiNGWQae/rUoy6I2beA4tuW1fRA/Tt7XmUetDOFbBYLxadzATNldgcvh
mvmBtG2Pse2rnX7y43oIPGky0bScrZClJKm8U9rYPYBjOPCHOYC4fD1xp60Q/mkR
CMTjYmGWuuX8/7v8p9qFeXMT3UZmryZCemNaulqe3H8mYDD+OB0TeDvZ6itDcfP6
XvPF6nXxwZLnHfVl+ESGwiobcCHrQRyoWKdcLMr/v/3gobXl9wWp+VgWbswRti9V
0o5QClBSo5U9yfiYYRPm7v1Y6tbzydI9ELCaTngYzd7H4iJdq/1RHHqVfjvdr68J
q4N6xqlNhSHjVwLEIXnrZWh2wsstjSxyvqPGrbkxC+P4rGbu6qkag8tWA3rTmmpm
aOY2KtRHugeMYqg98QRpgX5jrWB3oq0lCSSl/CIaELlMkaF3TyT1lwyiel4YUzxu
LXLiBiq/DMc86bvf0ehHkFNc6CSiibwOtB9xgGVsrLRBlD2C2a+XdD+9FEafE50G
BxvQLs6p+nI+RyOG4riRa5oujboZlpgoQRZDGuPewELFQV7Y5ZBzoO9xYFlFDFCP
o5DeziaOl/RIA9G0tlQJaeCisDkHu/R4J1awtNmtd4ocPEi53iAlJxxVauD2+/qy
5Q7uZdzj0FT2iYVm2FIMjt/o7PndgwPQ6E+f+rXHQYFQk7G6DiMcDyzz2vjIIsWC
oiL2Uo0nlZvj0gXvr06wbTypV16w3x5bXjI8m04ZFMtWjyd/GBXJ+b0n/3LbyQPa
KjqdyYJr0TV4ytiVft8QSJ5WGF7VqIbJ39PGgmPaGclnzUFLh4WCyItsffnS6PwB
qPIipvHEdoQO19Ffnfti92glKiAE7QVq6ZgGaIAI3H37mqHfdjuLGSb2+UOuI6Po
PbLFCt+9x1oxMK616ohvlmI3p49kv90P87dHiKpY45JqQqlYBXFlTVa6eQQsUllk
Kf5stX1N1jGyRt3PcfoUewz7gS2kBIAEf73ucInZmidduXytZ36dJzWci7/qXnkH
nG8uCCWgjZwg2yYh4yrEWkRMTwinWXtjqp6Up1P9O8dne4ZFzqny4BcYlxfo8BxO
qPsC6P7gsUFPafxv+BND1um3LRzPXz7NVWNnacCxKxiWhi448ykSIsJJnmdxes+A
kxAb6OhqVbvD+thfUY5SjUtN4HZ4L2kaoYIZZmzDRd0cpwMgvHTQVbrbcFYuA7/k
gMNaEVcS8FLUcqwKQfAabUc4N4MLnCPBkMwcbDapN3cCu+FNUUCPLGP5fTHsmN63
5Jp7k4ucv5zmoZH0T3pilJ04SBAB9E5RGBuscUdYJThaqs/wBuhddTfWI+8JxlT0
Y5bJouREsrOxLLGKjVag4mvv4hUXOCUDhIToDJegFpEwYkUu3FUPoiKWEXcO1sB5
316j8rsE7ahrEZEuiyJnuUm1RFqovH2jMnVtGAdJKEOkUsAuoG3Eh2uRoHWR3HFy
pf4zUyYSksZ8ptvJWKWTG7nV9IcCTkP6MKuKsMCIe3GQ9sJ1I3sXZwyzRHBnTuGy
zJYcFlJ5JYVVaeMxYULUwj/nZqFOTOnaqgBBROvUqMB9Q85iS92j9Jb6NB/1MHVn
47vM3e8Q9GiJGygUUqf4I9kTz+QvSJYk+Ph29qsLKsblS4eXX49AvHiANgvdHdfN
8ps5CeO13dF9FxcII9XxhD2+oXFxCpcCCqAmOlZ+aT3T/wNnBTMzEo+g1cSlrrwR
IUjUI1aiPxqnWZY/NzD0Vk/cuAUEvaVZoMzKi/MAuEdT1mwFcXt6cnYX+lTnzr6j
RwHKkaQllpIQVtj+SDAnGufU9b5LXOUMf6BRi+Ldzg9ndIsRoqCpCos1O1fCN4vV
otbGlFUcaI82B4Dvd4IaPw9mxUnl6Ajq0M43DLX4b+Vqrkf7KMxqRKKszrl62j1x
N5Zx4e2xZgirKHrzom6lY66d4zSr2WQmDPcLBxHOUaItTKx3T0JWCq0K6TDKCgAM
uMRwGXmNlfrdWtNOhnRw6u3uqR8KPyZV5nzuofHd7Eunc3dwjT10ikAg3n+PEaIY
VA0Bqb67wwABn8KkvEZM8tr+nur+7pWM+TG+OXzJsJeVO9oGDBSWQb/QTwe8SNP8
TLQBlwDQNzE/qO1IqCiCR093cUdff4RufICzME5QQExsQ361m8xk3J3OG7U8dELe
+myMdaK8hfpudwHdmOsrJA3ujzPhkFC28KUQktDABTY2W+epHLZxQLBdFU2YF+rB
DpyaOJid65h0n93ejbsNDTtehE8zlo/Ov9ZaBa1nq6tkVTZsaPGyC/ZEIrGME/AW
1NPH4VHT3IZQeq20g+HnBC5oC2ekkD+xjFq6geiScfEC9SW8LhfojMugzAnRg7uE
ccQSNUjAHIg0QQ7em6RVPIwNAqhYEEp3iroT9zMIzIyeLbRPPtxQtF0yRmmOQffG
fqQAaMlE8BSvv3zg1qwkKOdit2Y22h8A3BUN3NP+VRfyw+xhVTNOpGiQR244/EsK
+TK6sRfs62gacuUF9tvWMnybNRqADuyrRd3wBY2RK3fcZrzmLSjX0gKM+++Wprzh
fUocwoJex58P5zv0LOWLKbA14MpXXGxQ/yNswRalektlUGMiQQmIrp2DasRZrC2A
YQMc5DFg5elpZ8vRJIeWqJCZBNU04rkpcvnQsX4dyZksM6/w/4hy624/yqyzgIUJ
2CDmT3no47NB3+NxD8xFqty3Rs4wxh53THe2dYfsxlTbvGLOF6R8fg9f9kgbEmbg
cKLLif7NHK97mmpcvC3/4YkJtBrqn4JkCmdOtTT5qqikT/MKEMZXOvFi1XA2D9fK
qtfE1x38sUhkRlbzGHAjlMjMkMkEFJIP2AHGWqeeRnlk6CgmLjJhEA8k1pjRyyZJ
/kiB/SwlC+SF+eOJM3yzGYxUhAONBZkdV/jWcoC0N56aEZL/01zQT45bEC4R1UxQ
JKm/aXGE81zNtsvbwRTP6wWU+35YQPOxHWA2QSvDQyQ4tGvKTWyzejuxGSj8SAhV
Fl9odptD/uiuV0fChDYlytfm3WRrSIrwUmBYApOo1bDOA+NYkNgCwcb1lT3rQ533
mzHPonCjNJZt/RgQqIMhnSI5H48YoqufD87gRCNs0YoKqoq3Iil0IpPbOkoaEMUI
17STVPQuoYWFS3skFmzief2B2yhiF7TET7mvmiNhRdyAFm6rNXzrv6MZqRjlhbUQ
EFhlT5+moHa4YCUj6maJ3Rj415zyHvcopPfY1mqqA8eQMr3mkbIc2e65FOQo2nVp
y+a6LOGCh+CfHnZb7sXlxNXGqTzoRXAcWf7z3as7mnwhZo+yl0sIs6cVI0yrojrO
vgFQ5/U37thZMKgxxSXd2/yuyTggQvSl07W3IYrfqZ/OPL9ad7fCvSNAyQdOPwwZ
qMOTuzaHJ10mRevHrJ9gFkAkuP8X1/3pRHLlCebuea5L00O4xyZ3r1Tw0OoTmRn4
hEJ1K7zEmGT8T0/v+6TOiNwDfVNZ3bJocMi8zRevRNOsBYcUaYPoQ4BhiTbB55HZ
XxiozQB4PTpmumopsmiluN1PXOvMxKsS7uJ3LYEaZRO+562l40LgxpZSccMGasnj
KHQeUx8Ss2/DNuGQAxXMH8trPwQOM9K6pJHTXU7LZkPvtBl10EfHvkNEbShCoOcU
SL2ZmIkSFEDeICsOIsRjQXidKgISB6fbSGutCxD2J0jSaPQ+Zzn5nNmtEz5rQEu/
2RDHtcqyBIMxpbEFM+oVMQFz4DJmHMO8NyTx1emMi0cWvNq08T1yqbgPtK8X6Ua2
ntuX0WTV8OtcFC0cJByZUA4VIFXKRT0WZdW4e0EryYbpMGrZeINt6ZxkJniPXFfV
CnJVZ2f9J8z7iQyD1dDMTP2k2o4fh9of3RtPrYVKElcQfcVeqCnhgpZ3N726lAwi
Yf3a4yHf8X8Rpl5g+Ckqlgm9nDoooz3LfWp38qFEVN8zDFOjCldkaT+nILop3u0q
k7EeCmSpHO1faIfF6WB/HHmaP5SMbjplwN0V52NEHA3r8Ge11ydEzC8XdDvmxAD0
jG4Zf6Q/hMo4Yi2TvKRf9I/idOXNdPJbkSj4oPqOqxjl4MXHvmo5XMp5H0ObCStn
/x50lSEao7Cw7uvxdEunwlxAJqhnxH6ILmOlm5e4bPF0cblyEs2uSmrKQAbGfGrv
NXu85M2HvlRLcZyJY3cIUulRbvMRzhxzD6uz3Wn1NVXjyDnqX9nY6282dQ1PdlYd
j6qlldQpnYFhpyf1p1vcWFv8RDJEMWKVjiZ1hPIBb3Y+LEfNiVVI6bBBBHkLwBXi
YhDQCkrIukohzQYcJG/38RVSF1a2XFT5T+OYFGyDRyAwFyQSRk/MM5LhsrgrRJww
YtL3vjkOWuKTDsGdmUmuMU932gazJ8JTkt5YuHwcNmLueAqWmM283HJRZyuiXhH+
pr2rTCKPnUNmIkIUvhrNslPYm7lDzzBWIJyB5vyv0uHanu/PUOEZ1pYC2DLBCcsC
GtcAFhiAHGxYBq7s+QcKA4uAqgToCGy5BZ7KeCZYEH4uDFExCZq7Rz1JqwDNF3c0
krr7eeb96gLi0jQsFDUa7vcXkRLhYDB8AeUlsQrUndFiHFvi4Vf4k2Eg0Yg4P+ux
zjIkNbNNvNdy0G/So2X6N6m78Jgvyyty2+3JS0W5U9anU9ZuJC/k6cHGvj6L5I0r
Ch3IaGb/CsQI6YdounTKje6KxqsUqArs5INB3nLzaW3S9KvNawQSuphfERXUCEI+
qxArFOXLEfcrZiLs+cb0NU+vNuh/JSNNnXuk7nBO9yI8dv4AK8dG1LqfQXqgpJNf
wzp3enIfbk2UE6nxKRe39O19S0h99XuKTTPX1OwFegqpLnyZJm2cXKA67r1x8Ivw
fh6DDP053UPDsWp5D8zlD91FRqrhuyQpZrvSJ2EG6b8Hr0Pkq1fW7GgmTYxOtgGP
NZWeyA/V7Of4Xgs0c9GoqY83eaSLo2DMtmMRVvKXaBWE8snaSTXyFrjR9UKumrd9
uTyhPvriySuU4s6k+aaT4LxtdAf46HobD+XaF3xM088TM6wH2tUy7NKPH7lIj5q8
0q+7s8lKhf/pVGpy7l6n+w9LUZG9EuSotZYTqaV+r3zEe8KLYsTsl6gs6w90wMVb
KGIOzngXmRr/NyQ4gvmM0umOAzl/twnRGKJIqKX5TzxRzRqdydRAlPfn0GPI3oKo
pJnYjn8FVAVY5TpUb9pRfjD9RB/F+tIxHYDCDOKi+fRqMz+OVqMppopTUGUfaR2O
/CMPYaYO5cLU4aBVJosBTI5yND7AlZ5WONMruQMqjGVRUaA9g8FdwZeVVEY+C1YM
cAoPAvDJ5y/oqxBz3IOialqPFCEQsxNx7mcLXtRQ1+8unzI4uYavauctFycUDWT8
a8HkT/0Auo0Kz5P8EKazvDEqEMz6O54oXrXlS40qQNa65uzSDsAvq8QQOreEw/rc
rlxMCZNMEtKYntaQICIBk0ILYJTEp27ydiba608grEn3Te6AYEN/j7yv9J026sK/
wwotlm3SrrGKUrGHIzTIF7Dv4o4Y1ZZ1VLSHtN45UFGYMH0SWgkYfcQSEYD+47AN
Y238CGJB4mnAOtJm6/ObkuFuIm9PZ28F+3oG4qePvUMRrUKoKwBonuznZPrEVT81
y57VHoHqItMQGZVAQzvbI48N1H+OyFtFNwruUTEd8PUw/M4RY4mK80A1pob3WAXX
WPsSMs+Snw3kvYklWTZGLEgnjB7jZRFAbSTuwfwuyRWECpcG6zvkhLQuJn1fH/Cq
6YzJOFHuUVY3gFsXl6kjUm29DcJZ2OTy4XLcoNoef5w2JjZTH+06OoQIap5tPItF
NRjlQ3ImF/KDLcMIuIRkdiFv7Cwa+Jy2CI9GBVgaQqdG6cjyQluGSLHy09MTYANS
tf2ZiQEan6pYF8cTi67X7XOoLEHgn/nyRW4fvuUC69GwqTUH58yfo5rg+ZFl/KUx
lJMiEtuTX5zsMoFnZaVQTmiubSkLyUw5H/oJ/9HyZaXvSVAmsvp3sv4J/YSiehH7
+opA7/Jk1ev2aO/3AwPjQbHAYF8dHgHxYV2ykQZsVk5xH0PHiUMAAvkYkc361AgZ
Ha7YEQQo5tJsCEyFn9g3356qCxWmC0NcE5WiHaEJU/I4xecLAtP2bqpjZCKH4vi2
nvToarJd2Xv/gc3D29zDYBPm2ZIb9eBLxtLLpngvS6sjrG1HsQexX+SM0CtH9Wov
XCaL7/U9h92VuIhcW+YkrnLES61UtLLurnDAoTjyMXcfluVzhAu/WUKTJ+Z3fkMt
qrkvjzaw+pGrRzftvfUgD8y+Hc9DcBrQNt8RHLpI/sxRT6E7iXjfdm1KNOFynVS/
5lQtsku1Ih3xG+dqPF0lI1nkgW8B94RFv7+jduJzZyX+GmD+UIm7GBnlorfl5tyG
J+60dYYTKWKfvYBOL4tp+piCtJARw6jVDPPHtAdStJS1jQ/cVQz+2oXuP5DFYXVt
nXIwVTaDrvjkDYEbWuxe5UH6p8eTn9WrRiZskvcDi1w+AYtfHdaneNGvUAP/F+OQ
+pZjVczYuZVi5j+ff5x9gejtPCtW6G0Y0ejlJIjOSU/8mjj2de5jRSrFpbCE7kEp
dk8Lga2l+irj/kNZuY3Ph57rGvw/rDEbF1PVUi4lrUJV83pIXrdF3FvS7JWvwFAG
OSfF4tB2B4FfbvhF3D7WqRpCt1glw9mGny6tr0LEVlFkXmO/KXmmPBdDRN+pPek2
ziHbhm2QOzeXuq66mT7q5j8miahc0nNtEr/U8NmE2EfOv+uHCLL9m0IDxJpwxx0z
e91k26lzX2NcZNUACe2HkcZW7/9I+Fx7+qrUPAi8e24KHzwLA89lwBS4rKKdWrH+
WHE8wJ9h6txh1LCPd92jFdvKyY4U8C4FQYzQvheZvLS+Do1LS+PufXGC2ZKZPlw3
gt2m18L9WC/JshRapQA+UjANST8SjRUsmAQt2ZL7K4XuBBPfL9WzDiQu0qHjS+Ci
Y8rGGAysXdhK6rD2CAkImgapxzEOm31mG2TfXkLTCOTMNyXfS6kKOQcMOlQxs1UL
c9L1i2dbTLXr1vIL+YwZZh6DLusdojyMd4TC2YuLppzPu/h7m7QEt4hW4njJvogp
VJHYRhPmZfrRwvMa/Ta2Q/dBeAxu0C7tyVRZRGEG0Qa8nYpJQMvgp0MuhnZiyTTX
E6rSP+F253WO7GomLpWrTN94O7tQxREKgvOtbhKfmm4gqclPGROSqG0cGALIVggf
s9yRZDMu/7e+OsVWDvVJ45Bgw4THv3gfbptI10xwtX4v3YhcuM/yMsE2UHscJVgE
sQG0BuhySIyzdBjc8rb+LJD9vye3/VZNV/0odBGRgP8Gm3Fkh3MAKQPYbfuo/Lb/
AxpY2lOzEAwiVIndahPjBbURKmF1Ix56K/s+VmqO1zChx+9K/wYHLziwHYhH2Enh
9euGAqJYRPP7MklzzaP7crEkh+9YXdtT3d0WaHSOmyTsWxK+WKZ2HLk0qN2N9vOM
q5cpXlyOXudJEm2Q/j5mEV5vDMDIr6V8GGb2UvbqVqbfuaNVnDtVLYjTAIWTK/2/
SbnScMWMPEj41MLzvItsNzixYpLNjbcDc4/pElEyCwHg+ZD1lOO8ueSCDr1F5P9a
JzMkGAMWIBrtBhSxZtbTGq4KhhAWpp04tZ0vSL5DeOTaDpCJ/QAbn307zxWt+Z9I
++Dh6RBkJIb/WZcQft9Bfex2t2ivUywkpjJgDXkNnuEdVeJVErtK0HkW3gkzo5c2
FJF3eDx+c6X3WGgIsRs1p6UqKGpGzDHncoH+lfzIwsWimOBSKYvpyvO2YDDusgyp
v7rzUdQCpmZW+MDjIh56sJI56JQP/ZbcDJfWTNU26vs2tq7p84fsolH1x4zVtanp
+TS2ATZgAUuYIAyHCKOn2yHDfwBAzW93/Zrs9/DcsV466wK9WN9H2rD7wPy5Kye4
owf+BIN+dIH7dCaP0NsX9fTqGWfXG7yseq108PfRdJykGZ/VvLXN+w4TqDzz6V2L
dlp+t2k+wKCEaEkI3ZJFKW5zBbpXS/ICqpSvdIIT3fbWjQBw4C0Rb14IOeuUxfaV
9fHjSkpP8OcWUkS7j9e/Uo/f87TOV/PJ3ggk/PdcBHhPD2eNOsg5lGcTZULAqlRZ
f7tW3Qd2hH+ryp8RS5O22OV8hdnEejCdpvxNl72AHtMOpNtu7I8TRythXh/2hnw6
yyuyQE3jOpTgOZqAcxDe+2ymon3fQihMyd1cGjXpIyv+oBh3gegT1xhrc65lB+J6
HQ7MOZiAiOG2gCgHKfOS6zuBokV3KR7wTRBNLCaAHq7H6JM84Qpm2sa/egJjz+Dt
he8AEvl7GOrC8+ldDNz4HBGsxDEA98w8YTZpBq8zPYgkvLmF8MHTgvIfHBdUKM6Y
I5bya8Z/A7HYy6Wcm0FdVRLfSM/NVPDHrCe7nbWShduN8tTdE6JLHMmtWkZjRKhD
BRSibukplz7hzosm8JWRGihaVxeiitdTbZm7/9MICBJGKV/7DFFiOgR3MTDqXFw8
7eXvdUbwDetRc7CLZsosKj7wWhy3hQJ5QSYfE6w6Db92ru2tA8lzDHBqnVfXCHOa
M5MBNhE1k1ryXYf1j8rDXDAA1MmBaOo0W7Sr3dK8gC/r30YxKs76B7eE+iF5hfvy
XdbpnnO26Jz96WPZqTTM16Hsa1HllgnJ4GQbns+6rEk1m/8T2e35gl+cctgmW11l
ReHeqAFeYqGDF0BsgGh1Joy2L1pz/4ZZ4CDNCG2rXkfe+aHHrzcbR6raO8mYgYJO
oh3qpD85tuLxIoJc7+1SI0hiCME9QCrztAAS7RMilWKmzqHqxPLGCOpbo4XfJxMQ
13/NMkk4+h1jJmGPDYOquW7YvdKVYb0ItzJLRaS38mXdxL2GlVPtNiXTnM6a1t7s
pXogtAR5WnSsycrU6lJFEYWBu6dPzudzyBHk7O/9PcL9JV6OlxjAdi5vgrHUVylp
Ds/Memmyt8nur75q8HUFdBBFkIcUAkkPZNcSwDLi/dIhFMRsx5RwbrFLC2dWCjnS
hsAXorLTpnY+DeyfozpMWDJYMz3QDtSD4rZ9OCfCIoPPU8qma1nBh4QxyjY+2wAZ
9jfvhx/ldGNjGITAmTfBhh0VCERvYG3VYBFGpRaA+Pjnh0QheD2e3A0IXZYaKF10
5LkJ3jV0E5vKYqFyN0CthXINOGevnFb5XbaorM4CHPupDu5y+T2HkB9l9+c1Jed5
ffixqWPuvlbacneb9+ywCeGS44K7MvhjOfsWv/w2EtbHzaRYxHy4tWCHZV+wFXZV
FlDZGP0t36eDG2WlUaEqdY80//UxIBvfg2Oylm8REpdVMo5u3bP/0QFLUlc+UsLU
+JRVX1QuU61uR4vrESc+ZGD95pY8PlOdh9y4Bd3n78l5GP9XRGEMsNTCftMzD304
C+tg1pV4tHD4WD9+VPGBnHy8ShoSddiHGCSVx3bC36MW4wT8w0J7hlb7Io6uJwC7
Osh46KVeaBHoDmOglO163w4uszKeUdjyDsCyb7T2SQ/MGgUFrJTa+jkQ0lxHY1ui
k4s1uy62vZnrLpHfJKo9zLM6S08qieeXgGbWkhufAyqaI5OcMu5tO/NitLcVm0C1
LGvziaUDSI4MSb64623moX4IFkS0nDX15SE9Z5YYJWJlHsF+TarbaOIHQYJuVF5f
RfRizJeP5Kw6HC8P5l74xtk/QH7J0OOtc1cRObHqHQjKMwtanRv1/M/hatgRhUXw
HLsPaEicY+146XLAAn/MJxlnk+cf0vgGiJiSBZQIqDXEF5VRPAWt3It7qr1n0vPD
/jEYB898WKPMYWq/uyosApPvynEtNFvolLerbR5Dm6loG4ciyU7f49PEBKhOCWPw
Xe0srfb+kxuIk7EA0zAxWgLvZcmsLXDshBqGer4ctFqTdjW8Byvh5fhIUv/WZPzM
f95uApospveu/J0jxNBhDDqsKgmb/TIOm7xXz2IBdbiOhQRGqkkx+9TmtsLLLtEb
KhhrbYDQqdgOVf5QlxZWKO3wXF1egoRTUiGxnbK+BTjmec28NvdlW2H2SV1NLb+0
nvjopJE5LllVlQhTpcCzAw7ebTUA5mqA4AvrWXGcwE9VsIYEOaAjk0tQUii4DZzc
RFO6xfgAsgcC+tyAd+wFP4IINMXaxdycSk+tDndixfyqKXLSiwlt6cEb321g4FQB
W6ib/yOd+mQZ3rSevNmtnxDCfB+fkWD9jLCyryz18XfQVFl6OKwODO2RVMwt9sf+
TyVaDnxp1nKshy06VEXsmy4O3UuOam3mHls4o/eAT/gqNJEF4/U1Dcf4zs7q6ALS
6gVmompXjawIeUYCJAzk0WwmX0Hpi3ae98gmD1fNKbUMsag2DgdaB58GILLZC+3f
cBMe8oBvghZYzGSMNCEOxv2r9XUVHmLScQ58Gow0O0hAPglFjLOQ69JAz5SjOobj
rTdMv+h2QkglH51dYUsBO0wJMIY1rXtdndJTQxchkTIC/IPw1HN1rTyQfxypLKwd
/heZ83W4MM59yc3BeMIoeO3VtY6LaQEuNEiG8qGnBBQOvoSCDSVfsxCR81cWnlcH
HCJO1kEFmDwaN1xl0naUwN78gEscn5dyFvFOtlHN1CgQuLdkVC+QpOvqr9WzM6Mx
zhM0cZAiajiYkbT0Rx4/ZRur/QhZPQfoCjv8u5EB2rOieiC0d7bQuEE9bYY3EyyM
SAl9ZQOJGw1ptEkv1HquYNLommGaQDgA5khhKi+6NG+GUJKV3t1Nz/3I6laXnjQ8
B/4z0jRh3buIlrxGyULZbBpH/YnXOKQeJY0sm7n5PgSFTtziSGGrhwip+YIa3IsJ
XK6PWmVE2iqntyIG7D4bWgR1Y2bBjnAVSQgbMUQNgnSMi/YG7WkCEUeYihN4xbbt
nusR0KGqrT9lstogTLcpWSXZgAX5emZN+SORPJxWRFfy4rp13PD6fR60Ok1vB1Ih
mCkdO/yAVf2+OxPg6crymWWsyoqt+e/e34EVeYQYVVTBmbN/ZXnTlU807vKQ2k1F
oQxSUmSt5nEA9CE/LZHgHghQumFeRCGGa5C3fNfzfpEACKHkK3KzpORsNbk1NwH9
XX/sTJqJ31lDvRJou50YPjOcoLBDfPCRXfuSdvFWxRnV5lZyxYWE+Pur848+d+H7
g/RuoP1tVpWqvhWOhuKQPw7hheKChZJUTnUa8tmLuSwT9akX/5EiM4RFVds470Wd
e7WPef75U+4DiLsvMBW+zvt3KAqwTU67hus8tlTGP5YlVNs+wucc3bMhWqupGXxI
ZQm/jW5xIR7AXFVR0BdMSw6A+Y3+TH4bbEMxWt1rO5ZRpwhEqvJpP+W+SR1shs5c
jyBeE62aS8UE5jil8kRkOlmxOqJRteSfphASrFnFkk+EqWp318dRyF9nfv5Gx5dd
Gl0TBLp5Ziy1rF3WkdCHo+tNipfvnso8C57hKAeOF1zQuv+dA/5ELc0ZMVZjZWBf
72OxHInNsk7qdWwMqOPp4y2rDmmzyemIn4ZIIW+WSrfSG55E6otUsU3gfpbYMHoh
BGmdSmFGjuylSWegSGIILcmZ2Np/iEl3tZTNyngCRNeg7Yg5hTLWki6oUzgkNVmp
zeHpPze865pMrmwCitDukqwTnYAbNfEXCxobHBN+wliFSgE5TUv8hjlPeLEwDFqS
nDsi95oCwstzxXakDDCtOn47zKo9iLhm96tX3Tmfi13XDliZ7HW9TV4s1zQb6TUT
ADWVfLnVwIhYaEpRS7eMGKNQqNqjF0lRpJngyrLLZhEb+MKNTHTDqoVuKcKQednA
8GgRTxcaeYI198pJrRKUaLokFmxtL1EcfVWE4CLO9KfkV652uPTP+2UFRabzZaZm
nxRvxng3jwyo3oiKEY3TdTzYljYB4h3esja+S/xnihmVYrpMDdkgmsr1h1zERF06
VfW0xVO4q6QNInKfB3W7jwDtL3xIsKrHr2eD9JR0vS9iASfQJ6mT4WXeH6x+zcbW
EwJH8GLQk4wmhm6vmGR1pD9+5XkEZNSpl8NYaPUwXyPb/H8JJ6OqETkewOLQjs5e
9VIiO2EDnpwNEnj8r8jZ0NETQPtSnkoeLrCaZKwlvRRFZVChpXB2aBT2KqWbUDEa
f33CpwzlWKOc8H4wQOvaZGsMWAj6N9vS5VxbJxTNhnzfHG850H+N94t6nLSdXY/R
6zD1FW93Tj92aX+yJLPMHcnnIbSztiC4bwtPq06hWu90MkSFuzyYjME2XS09aFpW
2VTzjxVps4tcEaBTfHxSAwxaBScBKxOVJQzL/VNuw8HGGYSuqG5GmkCQyMHJT3Kw
Knu3wkBrXWQsr/uW3c5KdVZBGOCyibVEQjmSb90RSVrMoAE29K2VuuZ+zeZmIws+
tj0SUSGlCasH3/JfbyxU/23agxMwDoY9PfTVijbcLGkKNDZ2cuZ0jwd7gpNyajeZ
MZEPF9WEFMIck0GJ3mt7vHJFdZ0dO/OFBgUNLB1DNl7p/zxYSt8qVoik/wkMRIGe
8DL9SskYMcVV/Tvk+ajIzyNcPEHTgIE352ny0BSRvVYwoFWEOcmX70ccYCEqvEbQ
YtASvENvtgsSOTxHARBy43uaOTh7luH77d5X3iS90Wmf1KgarEmLUb5EZmbdmJeP
YsitodCMHSz6UyuQZSk9B6Fbsr94LWrdrOOj9wLdvJ1DimxCe8d1O0mzPF7boVJV
z3qA2skddxdTRMV5/DwFhyLcpbKtFMH2G0Etm9vCgmCTer04Ibwn5QQd2GehK5S3
/AzopU4nYMWyBMxkYjQifWfqLQx9xYP/DDbCJV4IXLWM+awFZfp1iXpZZeczpzI/
l0gzZv2aX9VKeGksseqm/A0NWZUD4+5vsRahsQTz3cSbvs45zSwbkwKIjIxn4IVv
JD3KDxBnC3KB0q/Z6z7gNd0KSBv9DP02+n5YXIYtcVIwEuvempqnWQz7kuYXasgo
HZxe+hmn+IbaFU3lXO+05QR8GWLZXXxwhVyC+L4mwa4HBBH7TBwVaTmS6xrxE1+a
ezE9PHlFWDtFrFjBMKQPwMz+ctAsCWYE48FzVjqQkqhPTBq4a4Sz2yq5uoC4t5rJ
SiOLe/egrM2GL4faqe0eaQNMaCGeD86lYkitmwsxQGbLe3HDYebw7YQ8loF9W4gf
DUaziIlXYazpQ7cqMKVz7UatKXCfRQsSc42/+R5H6OlfByVxao8IRNyi4aWaaYx8
5cSzYR6y/l97bHiMnrllvbcekd8wrTznBgzNVaya8uBmhRRSi/z/gHp5YZXosDij
3SFZAVvzAHzvP1P95iiM/uKSemyw65E+rRyOVV+1xQAGb8lyHm2J5L55Pg1NWvVM
+S3kPEAW3Ws6DMPSN9BNe98++QeCU2cl+Q6dFNqx5V2vgGxpDHnNtfBMzRyeUFoU
RHlRPO/9y71ZQzMFhaEVv1f4nFwdxmr85FBKcehVbzpa65AIcW+aoRebxmUw/u1i
zlrUEH5s3rfM7pUAsy5P4CXa4uSIoO06XJ96bOobQKJPdYIp6nNaC4jzVKJAT6nK
wVxTLtOqwX49cdXuH+vzm1Hi0ow1WJ+Ky47wxILxO9EVOiOhp4i3xHMlEQjEkNI9
BHJwYz8DeB4o9pthsZLh49ry63AHgs9xuE5MydMkTxL80Ds6rUZNk4mI+YeBftod
uL3d4NWKV/BBnycwSTe9Y6mSKjzb+QVYnj1sEND8LIQCNq+cVCEjdl/vY+ONJZps
s5xhvlW3Oi+oLK7YVrtD5CwSGsqNZS32lpefaliX3Zy9AZx0WuYxf9hr6ns0lB+y
pmcnsib5uaGOdyu5AliL790T9RSDdh5lDLleYt7rNGmpoNvfu4bWgpU0L8zZGb+M
6ILm6EeV+RkhM44Wsn4w17tTWuIBUowOjQrA3ZPFo1lk9HlOKgZXjH6dfjV66VxX
hwwEa/90VUUCzY1PpIzMbfuUoiZjCV+yVEyR1xkFvQw0/DTBthaX96xqD6mTXX5a
kqVF2wQDzMYG2o+3HushaGAOZFfGuiXNvGvoRamf37N313qMCZJopXFIvc8NreIf
Gl97dmb++tmbz7jAIIY6dkdaxyr8yo/IoUsdFrUoVDPuXIj1Sk+C1N9CUrawVQE+
ETCBwb8JcLSVRqCQc7ZsZLy1s4F2UT7ZTH73UERxZ1nxT4h9+DJ91t+itG7XqCkr
0Ir8+QzyhqV7/U/5HrzA0pYtrxvQaUO9CFb+SMfH1c5f9kUzaUMgLTjdu/7/1zyJ
Ibj8uQzbjtGn7ZPZw4qOODc1U5G3VxHfQoejo+AUI4741eB/3xcvkjb+2te4toVd
v/DEAw7ul9t09SRgI6YZLoonh/bATsqJMWILYkBfk+6U8wDC6Pknah016Zs1hQqP
VxZTJQpk7dOaSTyNdWUf1Be/d3gcLFZzVi1QWJXQDfsdwoxe85Kwf1oIYvofu/28
zjDdlrQFHIkkEXFt01G0PUiZbXBJ0O9YKY3eaJfvhukiZJgXUf1B5Lnz1+jduKNf
z/kFN9h1l7JS3XW6wxGPTxvZDB/7PBXs0bsaH9GGOSmisAZOyYCJY6k+Bj1sbGDH
9JeRF6QnyIW1/Egwq0yiYVmKcLoHcosAsmTmT0FlS/BARMOzoDeH3apoaNZf4KBZ
KWWPhFwuEk1MAEwxeAZ3G3+j7fw7siUmwGMcHNLraVrXv5w6FEVvcYtfa/JdFuwS
LX99yLy0GJidsSMYCxnAHSyO9gQZ/PwqfDW9F12H1j3X6ijzd+gRUY33oZNcYvD4
GuMqcrpY1x5CpC1JkgCGrSUOlBattzZIOSa2XvbCiv20rIud5ic9hg+tTs9+BSZM
3PBRKwNZnUvbaig5xbb50SdTzT3oSEXd7dWs517MVLF4b7H/CQJtpCUWpflRHDgv
nYaHLNAR/wFNHS8ZYJjSElwNGVqVbvLqjVbJV8T00Cffl9rzS3BLxqs7ZF5aL4QU
DAU7tteeohwIjkCMQOY1e/bV3mZEYl5NcPyJa3Zl8/wA0sdv1KsqgFMjPVozH2u7
smHTAzVYg2HW4ugNYGFvMnPbPfGe8xt2QR1rIKxB9a6dmZavZYOktxbbyDMi2K8W
bktq7iNMEOy4wIGcFi53c07N5GRGaHD1fLd7aHuS3uLnRjrIrOtcpfsjJSQfsJMN
ZNIIMROnanyimlmdIWthPL3MYYwY5DIa2skALnGCCsMcQ7ekz3Fyt/Bizz6BkFMh
z4chq9kdYmLcteQ/VKtTE+DYxD4huxNSQ6tgEHdd73FPYTwRp0yfC/DeEtAWROrE
YloI+0R22fBd/NCuQVHEzEjeeW0Y3HBbfgTbbppY4n34ycUozyn5q1qItrr9Mhwf
kyD0SypgadgD/KTNDka4V9Fc6CxAfnPSsf3TyZFx4kyz8pFBTqg16JuRBRSHe5DD
vcvS2yOWWI9WZoq0k8GIMugyRi8gJPZVY4ay2gibrMK/p4JFQeDjsJkTYtVVvtd0
MZdu/2fVM1GkpA40Pa0ceZWcdASQd/a0tQ90kxXDjNCdjwBgvzPiog8CkkUT3ZW4
YYuRn57kkR4koOFaNAqIjnxtclNOM91ObFCByASU8f3BYLikoaG0xcu3bYtwmqmM
cQD0oIfCOPNnmYVI6NNUYBlN5M01jFT9lqBn3I4v7s9r6GQeinMvZd9r267TOKFA
jwGJ05AAmYNTKYiPK+E+OW2j+0bsaXLKEXayFfeMx/flQEfx/ayBQTLvbKOwTTLH
KAq8Mix1sEru8pF0dFCWxDq+QiLaCkn/GC964rrfDLRv7uQnlc3Z6igkpKmJcWCs
jAYWSTpkJ9bwOJDlCBWBIpkIzdXWdrZ7ytGCDh/pddDF54qk0H2Pfrd5/hU2rGky
xR1crgiujQSQGGYjuLbEbLib0iGRARLeAT4hvtiOmb1tkxw1ISlFEEGk5x0kDl2N
Z56PWoGkKjFANFcC29HiDfvToQgDYOvYYsGbId6DU4GthYxsMbEXtKoLzlYowjsX
DU0z2flw5vHozNAgjsooqam8S14G05UYDdfhoipVkx4MHL1odz0oUm4R83k701rl
ynZq9PLTchpjJC82s10T004c0lmbIV1i7c9onUQ3fJR69eU1IexvplNFlc66V64F
0lTCjTnefi8SA0mkvu+qUsczb0sMPRcj4OTGPlQdOmUD0cN8rfvjZaa7IOW7TDYy
DpJueVbTWJyvmn0eDPTCNe/V+4JDeUG/rrhsqNz7wZRjes0tJOFTo+3feS322HU5
LpIGpiUTOpiW0/X96nbHaFZP1Z/k4T2UjRXuq6kw7pGE9cWg/2y5bZ92L0EuIpLp
QLhMhCQWccQiRJmGMSf76tROdV1TjWTlOp6t/xOUXANx2dc2leGF4e5UjXrGWxWn
AWA2/e/4hcfrHBXHvmDHS79MsSWt8tsNbpO7J4Rl/aztSyTYhiGvfkQdvkOVe61n
tuczdhwBa8lWwntPVkrjEAVjCchUr7D2e//q3vXQlCvX9mfWRZS/lL6z3nECGf52
q07YrVp1+24kv1MBNr6WELHOhIR5mKYgc0FMLNTBF4c17/wI6FEm/qdbfyb09u5e
9piRaExVd0MgZ09Ht4yixnQuPdlEpKrm9GnZptm95KbLv9ujkwbAWm/9bzTRRxtx
UTbPoNpmRuwpXFDLOEOqm7WYMfvzgY6SF00+k4Ftujw73q8gdYLJpF8A4M59qMYZ
a/s6gs0YLz2d8edr1gwxZFHAYtluP5M3SkpDZxHrr5ynd2vrE56Ch2y7IeZ9q4Ef
GhDeX8qp48jVzJErVUzBxmjW/YCrINbIH/CLUvowQ0sNn7qFWpORH082hppjymf5
XZuWbgN5B6K57JF1kdhd/uKfwWQmpt+J4AVSEY3JV/EKGX2jXuAaOqOPMMsBcWXB
30lZSxQyqmQVa2KV2kQWjKurQ/OHeZyzrHoDTXyPmzq1IsuqqNWaqmBJRc0fXFHx
4kJFowux3eVqyczMQt99wiGmBjJFwtjRt5HZmqS7faFh3/MZqmPqxZKfJ8mlecOx
IugD6BEQUYjtsSYPA8IDazGru4Eut9DwF9IVvmjcPxMS08YeN5f6j2QNnvCbckSw
jLixgBgJgELS++rE3Z4P6Zj+M8K0+iIfSOx1hXb+9sVUe2BnrqzO7MNpg+w6N3r2
Iz5PZ+lIDP4pWr3XxoAvromgc3YwrTAQU7/WIgf3tUUx9LwcW0gnGe+NEKbWYaPM
eyQ+IeAbm3KiV9Ft5xAuDtbzq1B/vaKonhl9l+eTssxsxyeYmc+kKVtq05yBdjPp
xoTdOSvHu68CpuKlfqTGKt0OfElG94U2/rBsd1/y9sq5bPbPKUpujGKBsdu54e0x
RngPErVCaxaCySaCgje1xpi4TAu3fx5zd8phTChpHRlo40luNggVxoYfJSklf6ZM
GMHf2RW2hEc5gMB8aFkckq6ZSz293Fu350TZ+YvNFX1MfJWQlflTCuKOAmToVDte
VXiMXJ3WC0WUovMfa3V7q+yW71AZAcy8Z5TNRT/HtoYg2XtVCPGIYHKf6xTfGVel
uB6jgjWgXVrFucyOBfq/baSVfG2h0S4DXcj7o/T2q4PROXnaxN4bYdwHoKacHRGL
bUMRen8aHPqXojy0qDR62uBvBIMrcMRmgELzliqpD50JXP+msx4rhbHC65CPPTrk
uVqCS6yzN7Lgyh7T0KuvXeQPicBR44YcG2wtzYoni47ijQrgCBa8JGgSihvGsAIT
W32a5WO7VRa7ASbziPJX8mWC5FnGduU0ejjJKDGitlIYJylJdjGJWZ+1FsTvDuI/
mGE5Z723KDR5C9NiKTBJUwdO8vTVS0mAiQQGHfIYOD0+qe0195gRFhz4QVQUEaAr
ywpJssIhcaRJ4sWRI9WdQifBE01qCOKih1q6NCiKNmjuB8Sbe5gFqy6QhviP/rN1
lfSDFM/4jq7im9VFB1pDUdx8lRhiYrR8kj8de8C3yN9TQnSZ1FO4GtOf3cLNQobe
gznZbukz6KDzNnn/wQz2n9x8WIFny7MuJh81VeKCX40B29vOdn0c8g/4KZuAYMFG
ncAeiDmKOS9KHJuKBRdPnvc+kh3RZC/wVl+XUYakz7Vi/YZbswUWff4LpuvcmMQz
iF9+pKNKH+6uqMdadzhdmie6VYgRsOHewOyRKB71cgxmkgAqBDbDLegZWXB5mlxT
KSURGA/OjVWuRMMqAeIeC7p6NlP8rQpVph05w5nJXMQd5dcOXzFFJjd+T0k0bYI6
PYo+3EcEMudMxQdaL93BQ0GsOgGTLN819umCOAfD6KDm/IokQPKZW2ubiJ1d3dPA
uzyp7/2BTfpMviNn6vUYUj3TSFVOrWkBvwP6QHac5MTR1v4jbiB0Z96L0eLnjLv5
Qcqn+1b/5J+yxu5lU0fDQJWbR6QmHaddOqiRXQsq1ydj9vjii7gpZwNSPpsyjkmp
M/PeDSGEIT3gBCPoS9FziJYDvjtrB5UQRXmXWQGKTJ/YZl3htIXyzhpPfBPF5O1U
LfUWEQ/CONEDYjY0xD2XmCswD0TA14pbQ0d8blCD0QksRdsLrIIXoSFr/1/3ZOTg
yaVK5xL4gBBCM21voiNRGBRTiwD/X7ekf3h1h0lWqUJKR1sGnujPJJ3btra8T4SU
MZZ+1Oo1nQm54PHVXkc8XIUrzNcMIBEKSCfX0QS6LxG+6vTzNG5a39wRJfhsNicr
h7J4w5aM0pXx+RHqr1TGTxwjjiP022stZ+GZ3oIEU6SWvoz2g7e3L7guM2ZmMMOX
C3oHBfwOCysnkIjS/Z8lG1TVbpjmtBOrfCKny0xxT2gxfz4CKZaHzgdhB9cCrh48
H4+F2VL3WGa1yRtttOktFh22GQOtTvK4xzzSkzRAFT52CIxBN16qG37aPs+dQddB
gjBjwZVVccnQ+El44lMHMOF5wEYjvGU1Dtp160eXYUT81S1GFilYabbDA82kbnz/
RgsFpdlZUKc416jgDmo/IN8WYyIQ/sEKThu8jSts6DcoeLQdPiwGLxNj0IGFaGDp
LtMT6WSeb8+ZJF6dBqPeeVa82CJZLoySciDDTBtnw8eEYVRLqXPKqEleEYfvuSty
S40SVhVRoJitdSmeDP4PeewXN/9BIhby5lsgHda0ktSIBbafiJzbKQ+plxS3t5h/
8U2FuzZZFRIR81ZAOEEoaG/OupHwqJDNKFROiserGNDMATeTdjO7JEfXavAaDP86
npVkgyxFunb6T+OVmesoGDR1aAaM7mm3pTrDyZhpsDr+jXRs0i0t2BZZqjYuIvfD
Opf70a5O9zIg7rHlkdq3cL5RLxpHmRfH63qjcox5q4Sj4lvv+NXfV2hjCKdV1uVq
xO4WvKuvox8DelQqkw0h6Fm7n3B4bYjGKek47eBjvVqZ4DPLZF4UDzgoQh3AC4CI
6OXC5p2bVU2tMwom063x1fbMpvyduJLePQfOMWrm9nETamQtGNCENdvyWFws0Hcq
SmCXNx4k+fHdU7Tf/oS2f1FabnkTzoarazQJY0tJoWct1UNlJIY0TKas/WM+qJBw
NULJVQPGcFrnY5fnXq0aIT5N0uxIYwt4fRYrd1hxEJswJfL5GonSfTb4+RlHFosP
1o2B0SS2mYRx2BMmL8pMHcGeZEiwnfWoyyuvF1oE8Ca2ouySfHkMiAcSkjGMnGsy
7D5SnjJk+beSjLk/006UpdFlZM0RPW4EJJC+JfsmgNURLkUcQn6fZeeZONISWRe0
0/e2w3cVNINrO4TXOd90tX1tJrtyFDPnQVmb7dhTWqPNJZNc/mKoLw4KmKtKRAex
xETg3Km+gVaehdnCDeljlaqtWl17d2UqybcidJvjcIznK4QJPKCqKx8SkAnesMAo
i0siQaAM1pGAxTtrMpHScWo9KGdoB4fXH9k3oeIOQL0ek70m7JLm6prG3Uk7tTE9
y7dQ495VZl1AFHZ1klmKxwbH63ZKiQG10tQGTiMayPSZBix2HGuMZBrq28b9sVDx
NROmK/Jje0kqm3XoeRmKKLeMvp6EXsrAPnDEvEFtnVTFDyCa6hrigR+rKHmmPXtt
oew3PHsQN367zJOO95du3y/OowozgltT0+Bf3Uv29hmBEFwLyXcj+7VoVuOc85P4
YCWLf8IgA2VctPjfCKOdPWU0K/YMRrWs91Jz6kIn2z+l585U65wmN4eN+mM6L6v0
MOILOBJfRbNzHKTA4NshcxJ/n3p4rPED65S1OtDONMSy7Q0TjdjonsMsap1ECRrM
DR/3hiuYChC7ZyOHtKVuq0tBM0aI6MKsXh8YjTDeTmoFuJ+OHMHJM7nftqrqA0Oo
Iyd/j3z1rXFF976p2DE0NNfcMTIcw374xTCUb7MYjXPrEZZ3AZ8Kxbnlru3fnS6S
gLZDqigfP52iBlllivRI9CrabT1pzsqSGbSxDakYrIbarNPC+xprDdkTSUrnwu/l
RixInCHZNRmwxhMd5K3RO3tZGssJGKeTVgL0FtPnGvsQndukjUT4vwCAXt/B/sUs
QXbz6Ld3TZMGuYJS69cD14aX7F+K/R03tJDicfwcxdIgTVPOqiaMHV13TikDBaE+
pqbNOpiRluN4eXpVEY0HTZbqwoA+4lUzwS9qmClkuErvKhesGoN1OM8oz35WNODt
3hh5lT2/dnyOQ55kkzeb8WlpI/KK0TTGcjA2R2hemjFkvSqR1XaY2Cwwrf1bCeA3
QHLo5zvRdHIPN+wNKEs9Bgk1kZKATt8W01DxQ7uN8rjYe6zQw5pZfUSY2QTyEEJo
NMeiUfa5xh0Y27cHeNe5qeSCeAcAc3QIGiCm7tvouPE602mMI44w5rl+ygEOfpbU
Eu3myXGYlTEuHdrxdX2kg/FAd4JNHUz/7yttOr/f41cwNm+FqnQTmKFrW9dAkMR2
RrDSgKDAgst2r4sOl7g1y16nvxVV3NcfB/H2X1bC8KoGkiRoOO2mVhbFbS2rURje
WLNUS3YvRqrjATyqlCZXrcqfe8Z6ND4NQ221K38GP8gG4nMlTl6m41KaFDx/nB+P
yWh1Kp4MfmPerqvINITGCqsP6mmYMeg3rscloco+qqQBLrpN4iTA0eTxLJ96xrlA
BEy0rHGqr0IqaCy1J7Oh9jW8V2IqK4vX5F+X16cySEJxQ/i6sPtKKaanLmsTcCXH
PXG2ulBVvqlPP3I8/urNarHiXZWWEqew2ag9g6uAheeqrGok04IH7zyDk424OIJa
s5li6CuNYl85fqaKePy0o8PjJ84Z4bf9O7YwVttYnnqM9NzKBYnkwz0VJ1GCvkT2
YDxzGs3t99Y2cqXtxebVb1ocgbvF9TBtIi/lOOAVOrh55A3PrnIwEIEUYKezrNX5
dLlzTJMst41NeeIPqUwwHbf43DFr8/usybRlra5gwLFELViuYLvbCPLdN7s4pG4i
dNZ4OW4zXKwOU2MRF7DaI1lTITdHyF1etlHNiXYoZqwpd/9b5a1CiTeqihjRacZr
r5Ep/NdfEgTcSrO6/dWVnhICq8oCcxX9ekdF5KMK/9VWRXFxRq17RtCu7ZrEHGu+
dgXY8yQb/I65xm5z0jMOXoLLwaNtVbQsD5L8lp+5StPQEgoG6Aze/JBUazzqAfZ1
4EVMIaxsu8a17TZUv1MIzxqrJlg4D+p+MENIjIQc4DO0ehXHL4CQDBgZv92HKluH
tbsYG4s+c/XBihALnZ713FCGXLzfczzxDv4KaUaCQewDxfGtiHnRLLqlTfjod6Hp
UDIoAOcebstEDzbJZh+OujSy+x+SUs0bUO5lTHAkflDNYX43idZ/GxdoNX+egPbH
kx4lBnI9kvvvY2qd2p19lZmgL0oDa6Qq+GhOI5y+wx0ySqpnYopn8lKvDMdYIQkq
7BPS0LUAYxgFTAvwOxF+bcPwxHFres++M6f7eDC+tcuRlkujzaSkk51MmXyN+4nN
31T75rpBP3blBhFFfNLQuoHB4fsWpTUABLIJTKwhZA/BAthzTkmH/EdeBHiZSRAT
jj/USpHr4cy96t8lCq+jSwMp6R4VUZG4EKsqLvdAWCPa7vJjibRAvnCQkfFGLwCp
EyDEVJU/XwfESfNJMuIU4gj+gnZuRqkBtkI9sVSvaG38LpPZVQF3qD4dU0MG9Y65
pxz7Y0marWO9zf3qe+C0gBbEWtr+b+O/Htp95j9dxqCT0tTyrl5Cw8JHcEoi45KI
TYsisZ3hK4g29bv4/wIh8ssicxgjQIHrNjqYy5VawtorxxbzzMoloHDR6nb9byCK
ntVUlXeae17uN11LGDdUpl2cJVc5SyBLiNvJ6igy32FBWdYngW7rJ5yS8LoyhhaB
PuIZJCdbCMYIqabD1qtmVb2ucNx2UCc4K3A6+9i3LbPU9vdMC6Fhc8Y6WeWHDf/Y
1KR1XVkuJFfzQ1H3rkv5KYM4i6vPNaWgl+p0/d2h/0XcS0LdDem4kVkzV351AsR1
AA1RAb1qNblNRUGAqf4Xn9gmFhZBk9Q6DzxkhfdkMDxE7DiUyae9LEG5dbz5GwTQ
TTgLqVS1EPi+BGvbPwCvImuPjeAxZNzlgmN5ZNJvxB0MK/esTJfyRlT6FEs2PZaW
Oac9oxIl0jwsv8g3/VdTMYu9Ml1Zgyi9wsJu4UiK/zp0sAJf6E2N2ieO/XpaloTD
8knbC+TVlheSRBWR51u8cuHGSWuCHrQFjudU5SS5mnf9a8o3bO1JQFEkxc6WFLSm
b+kxNhMBrA1xVaCh/k5+JLm4MmiD92GvuIbWy4/NbXRvRT/v1Z5b88kS2JKZ+zLs
7Qw26az+CUg1jAw2UnGcZfB0BjChrhqVIKi0nUDbHC4W8BI8PETqZSwGTlYHMVAi
STjKX0Ma7fa+jQvpL1MDBhkCxHAr8trZrUHXn4blkj0nolPqx/K/VxW0uViXncqI
HHqCl/JYmg2FzBP2jfGu5ht7Yl8iuVn1/GZBWkpI38wC68eTSzxK7FeSFu/G6PO6
dBCsB9odZ60Qfgpg0I5YC/1+qXY1kU28nHx8fvXS0hYBiAMfaoN/61dFhZdC9F+a
SqN710ODkY1ye6ihUOrkctUp4AIUVwexIAULs8Z+1EDEHgzvNn0Awi3Je4tQOica
uMNyxLMdW+6gzUMf6dqZykRhDg1I1kw4feUCI9ogumtFhMw106BwP86jQYbcqQga
/40o4osXgO3tEggvTF9QmOP9RDi3fuK7Fq7GUS7blZ2+lOMaQUo0bijUdQtFkHwA
5gPlNz/eF1IEvp8lthqSWBZBWZnHga0goa+UkcoYfzpWxfEfW3eXLRPIwVwjR9LN
aD2qIF+ZaJgHafsNORwe87cR/rUUZWstk0y/KrjckIhgFHq1OQKvPlPLtXiC1TlY
GKs1Uem7vYIZZ0OFMSL0W8324/4hhw0DXFkuA772fgCeH3EUYHjG1A/D5ktLN25j
thkMRfhgz0QzronSOsZvGn0FJ8zbKliA69axwpS1G8r5CFLN+rinY2zNAK/pdm0G
He7YYDXdRjfOhx2v+nWQDpNMdrmxs8wqRoRjhZ8AUk+ShD91QfLlyku1tFO/QueX
iyFWaaMjKVdF2ennXgz8dqJSYHExrFvJ5/o28hJ3OxRdNUKOAjuOXRU46gp5Cwok
H3Jb/vG1E5PMJcgZYQxx6kav+BY7nzSsOjRi8NttgHfUQ9J5QM7xllXgu4di9fk0
y/6WJAtaWDhuOCModlX/eQvRdbFMk4kzl9B8gbWyvXm7s/VGJ5NH8vKRnDie6+I5
AAuyxrPbHvrRlATHsTloXrb+XyzFKZCvWdBdv2J2v3/PnRkEXWJIu183BunHOxdP
+1OOpsnE04ukLreebD59CWircKqPNzqeK3oYouoFPMuvZTCZstGIF0SVqowxQ0VH
PuvpCbA6qafTqc6Qh2PCr9BOvC20B2zedmXqWKuZlMrw5Hug0puv8iJ6NkLIgLmE
VLWkX9fLIJHeemkGiWPz1IIDvpx6kEjc5CQ1856OH/CrqihRVeiw+ZVwfoi2wupC
IWmlJ014hJ1iLO2Pgb/PMSEjGYoJrc/9HRaPUKBvwh11y86VRsCEGJo8sQZq5YL5
i3OTyTyA8HtxY8EDi7MNmX45eJdj6sNvimMM986rA/4SXDtmbqS63BdEnd4wNPNK
7kS6xVHdPsA8PQtxWRA3VJcuEWOxRh8/O75lzuFq1OzXrjEYpJ5pzPbehX1ck2sm
Ve9EDtJK0JsMusJ1YiGMui+kEkBiixNstCU45KWNYsIjlRTLMWcfyyzzz7hrPhhE
D/66qxT8mSmYGKvVPmPZX4a13UQ0rCPizNUPI6Wt07xqtbVdJAr1jcArgOXzpyjU
O+XKLBfWM3wnvXFbquDN/2TPuockSNDGWeUymqrUaFVoC8AfgejO+X0jh0ymsVxL
6DsWmccM0mye+9uljpN14/oSLZP4WyZ30SZ4rmn9Laqg0eGmBEHsDoSzF8MzcFav
EY1SIXfc88msAh1XxBBfz0ZrWtcquuI3mt9CshQ7dG64hTFyTqTltyE3ic1UC1wN
lC0tCfR7WhKF0tyqaOKfbKJq0jSBEDuAaJ0jpXCJOZzLS/Wuu7y/vbSj0op0N7sb
kpPXo6U3yko2J7/5xPZm14qz6b8VXYp9Ktx2Sm5PW6LkBH0pt/O2rwzQUaFi/+x+
xczkx8s6/Xg3dcXxJvv32gEEOswqvmaWa0CqJHJ7hySXrtvO8eG/2n19NvIrVwEB
oYpzTR95jd7zKvkn/hvu8qX7Z4n2o2w0je0ULb+835wNJF7qWrDpzWxpWqQcsfGc
WPQF6mfzZk1onNfdTO5TsEDOZ9m/6SG2fPim+sHckLTPnPkquunAi4NhpuSTeyxy
0l4I7yVy5oqRzR7nZ+RT+pSjP3bx/Atv+gEC35+9tHbDVcbPKVUc8/XyHXMJl3ce
QuTnF8ChaSmB9C9MHL0vcLEuIi9bU6pZC/HYIWNzbH3ap8QJJSq/p/KCxYFl/0xe
99drWr5ri8XLyHFrxbbd2gQ1U+uVAQETSNwy9Pk613tlYMnx7QLQcflEY9V+X4Mi
Kk4sBpRpYu7Avw/N60iDctz8vRC/QTTurM7dF2ZAwU0jWf7sntEDD0NGvDkkmy/w
NeSDd4tNlKbf4iWwI0RdwvMwdhPSrl64zGAO9fEo1HszLs+waJqK2GMwVLgOTTtD
ipuu2NYNu0/65TiqVUkv3rp0UZfluc8J8RCoCYltQhuUWJ8bnBaxRLqkfYbnMjLc
DBCr88sX2Ki599Da8Kt/dTgQ6pd91ccT6kd9ER1D2/4YA0mLqO0M2K7L/4PyeXjB
aDC4dMNQwVs/Qyu2jDge4X8w7jv7eezN3kTwLRlEZfRXkf953KW5I/rLVn6M2mWt
XOJzTHQ2XZeJkEgRTLgIJ8Sgj92LsVMK8v81oEHPe8M7Q6lWkkzOGwFc87jKW6RN
T0Smjlf4BA9yXnKIWN1Dc15x62Y3/tcxAOLkkERjUsMHobC5qFgBhPASEzegzRpR
eX/91dAYJZVxIhyTHf7T+QUUrjZrHP63lumrpzTc+YlZKqageGTWxI/s46sD0ASh
0LpscZj0pcPSLqnMnp/u4Ahq5RRvUFbPsYRcJ06lRzHYZeOMrmNNezINLwzC438d
lW+WA7mEqfn8TaUo8Ru8Ien7R/nkM8CFqJGwpYdIAV46mgqNAVTzOJlVEH2ujCna
XM6E8TFsAWe/3qP2YM3R/HwCvoqjcWX0xSjScsdIJbQjp5tFDXQg6h+RJ1Z+Xuw0
McGrIY8DYn/ICVokT6AGTdNxRCAObe81vJ6zInQHa4AyYPAm0N1jTp6n7PPBdUE1
Fr6XXu1ZpT9fYL9liuI/Msc2O8eOZdR8xa9mi7CT2VvTAmqYawoFcDEONeeYYYvb
HPFrUHbPohDEZGYu9xQz3iiz2yEvNusBCbuduao9Assfxv4mop6QH+/0Nt4rI4dk
25A6ARmazp6Y66zjXpRlpBXXAm2j6Dk97hHxdjTxTZMvdIHGAAT9jW3SmjD9L9Xy
1gv09OfaQGVPeirw95ONdSk70K6wjQLkp0y29PLi5cZWyAMagPiEDMXZzqAH6q3P
BXnF7XmvgywdOwInbi3qKAXR8h0fHC75TwprP5AaFSyI66OMnNjedQn/QD1P0nFH
n002t8g3Mep7vwqDpcBCmedMpBtaN4VC2z7Sqk20xOqTwFC3iAcPQ+MOoIRKTYZM
oc7JSBx7fjKEgxAyGdXyknsw1fQ3TIxGuKO2mtA3mvjvU2Y2L2STpPjNikdq6Xg5
zZDlDBbY3ExWA0n/K/lVu7DSpw+ovp2ZPdfs9IGzN16rbBXH4YuyxxguAvvMSgls
mu5WKqXd0KfKhJANv3Z1nwzhRo1adzG10zcWFJ/XlLQLpyYiINQnm/FxZ815ToEp
XWLo20FiNWusVDXtBBKj4SEar48S/MWHtk7KaB+iHrHRPg7BJ0XfbQZlu3Il03Lb
De1JHnzTz+ILlWnH6NaLUcc4yDduyV4P53KDvvsAMGf8PLOyad5mk+Fo7eYH0wuU
w6kt22D9isdJRc3zwbQ60Bwg+yD/R0q6GIaCguD3nMCe4NhvEEgHDnG8ly8KkdNg
+aUMijv284WvpGbzujAgIY2xwcjlC9X5MBWdtmT5YY54x3t/jAdfyZf2smtPSvDx
1nlsXv5SGYJD65cfDYmoAgjHW36vCnWMr11REMmAuPfvkJWfFaggY5hW1gixOfGe
jSvt7y2sIqigl/pIXsvhq6C7wCWWxABhIk3jOZ91Nd94NaQpHBKAhpgt8hpAt2aC
8ujfa/DqZE0izVVpbPtHqJKunK3d6knvELNfHSMl/QaPAMy+sw64MVGOGZfEl4RE
KvAMJsWtJZyE0VRkAlxyZggpn4epwuVHQ0XtoSvwggks7+z0TqxjMlPCgufUOT4U
fJeo9yU2I/h3xPHHtH/51beHpm5xcF9QckADpJp+m3QQI6BWUKRGq59BUcXl5Au7
jYCoDVr1zpafA7jzglck5gbGAdFIgz3//QHf98bIar9SnAuUyOGIv6XDKsFqEDNA
pia7wY/lD79rYYr5FLWu3f/FvnwWgfQk8VNNBdOimyWDNnJVd/S6v3kUs9w1rcEU
I6mMjNvcz8gjvC2yWsafJ4ASpF3WREvd0T3Aeqen35liOnlRmD36oM+JXOqrPHoy
C7YqYet6gK4EQskUfCu2B4zDJz9KasrG8QbBUuvb9XetOeYclyvsiEmYPSdjLtUw
W0vuyiJMDBp+Hs4rNx/kHfd1kbq6KYoPRoTTHHXMrq/cagKlYWTnvVX85vSPpR+x
9hHeJFT2p+WzB1B0qPeuqUPdt5zwFJQbw/5l2OeiBK7haOTV8BTDHzOND4+IjNqi
AVYLqmqDEkaf9uil+vSOxRDRDqc+JV8CfOpgQSsKOSooA+uRh1loPGARorZFoOwf
p11I6w6QRyxQbJHgqgub2YRfvEUDd0pivPl5A6jArCTTAIhfDC6rwPJg2TgDZbmv
iGfAqvMnIzAyPGIc9gyBg90FGuTllS9nnU/PlCU+hIfguK9tdu1QW+x7urkP6Mrq
VADYpjtaw/bCCgmP5pubbdNl3FOGQomerc6tZ85yYCj0f4IzxMIEIfYbq1OdZFWm
ESBAlhV9H1BoPmxqyk/p4bUBsVEhl9pB04Iqc7MTWOc9kvU+m7DIfWH5fTQCbYqD
1Wv6GgXlsfTGDwODyDXDzFP5C/1ca28zMwgR+q9G6TSvtaBaMCoZZmyCfSSsl2HN
1iR0lVHnrjMZ2x9sc+KsSWQOTXQLTg1ktaowTWYgnjd7xvLRyBVWIv7M754d0idZ
YfyQaSyIhvmBJ8AopRO7T8F8eXO/ZBXgObAhh1kYysvY3Njzr9P3JJKKIGZ8Xri7
jev1+0RBxRVueQGwbTjCHto/Uz4htJd2dvislrI8D/RDGXwt/D4ectpzI5wlhyJS
2eXYYjHgYyv7YF3ms/76B0hKbVYPDZAjIdTy5bVaCOcilP7Swmtn2Vf0Qc5pBUdy
3kvQ6ZrZ9H+lsOaMH1qqo1mmw7FBBbRLnKNx8oShJ4IK4rU5AZUs//Re5yYfk82A
QhyPdyOkq3s0Hw0BUSLGbtFhKGmk6DxLgTwR3wpFTBqEUrhF7NzCdR4dMWWWNHpl
8iMcOlRskA1U4wt3nxK+Lurd9gPnmMK6mBM7mID8EO++uzMzB8rNoNn/aLDdJc2l
bANkPR5jvU7WmfwpELWV8LSczvmivzC1M2yH4wQqAzOoR+bsEs+6KJUqzd2VH2rv
l7l6FgDC7ywYQmiOpUFUcklYEXfo3jEWRXyo1yAvRhj0LC9M8JGYFgcN71Skuovp
Cyu7bcEYphcExPL28lRS4ZZ4JOQopSYtNS4FfKXUv8wINEz0WDlJJbwiO0P+m/Dh
s/4/Efm+5wyyOcjuiXb5Cwfxg01R005pJfkYU7ocwhcTJdTzkuURSz1trQbPk9tu
Z6FsW7Rqrq2JmGDb1uzRLtl2t3NXwEUwGH9Tf00EWOmaSChW3rBazIiolYfRjGgu
ZWa6mTBDI5tIlQMpDFxMuYWLEhwCU8kD53uvdAW9I9A1PKkRQZkHst1YJzgACApd
iifoiCXhipDQWi8cnMXAk/9coClR7k9ysnRRMldd8vF9v63JY4QwBzfI+kVddZqm
ghuXMm/UKcTqpqV8KzEJmuVhMUY/+c9Hs4YSHtBjnSwACyJZ8OGSKgzqgRi5Ebvb
/mo9zlcJ2MZuV5Sa3y97W2R8jN4GDfvVpq1j+8S424z1/JV/0N7kzrXu7W8zChZ5
qKJa/oMyP2KJr0h8n2djq8saCJG/icNUCGvLB2odYAUnM71fSha3Zm5FnFHwVPJT
FkV6cPJL/pe10VaSXO8yXhTSzu7IfymHx9tJIK0BMRKf/M8b0EutCuoRsO4q01vx
1lcmStbtyxI77NLuXFT7Ez6zjeDaKdy436v+1Cn/Ejqx11j9nqxLyAwX/mTQ8oMG
ACOGS5+cNSXc6Wi5et8vDuLDpxF/9Kg1FSGMFD9GtCBM/Tk6oPv/3lNPG/AhLzsX
j6k91f9WmH2DQGmmJYPUsgztgr1t7Op3d4oD9r98v/pT5Hd0+wtScfEZgkJbTAc7
VV68SUFoXpT/3vC9LhkBz32Q7eoUG1h/sjVPkvEb0Z5hNGY+7uoG7KqA77/NOEK5
FnJ9QvUVCUywm3EjvOsyxiK7T9YZ82kY7gRQ5xsg5cjIyHtOda3Hnho31zjOQ5o5
rgbrJfwVQwnSa4fDnXfqvJuV4p0isnOsH9TwMfXXjTjMhxPIlYlNcCJ+6UAuVoaf
ePXj2pNLtzwSmUHo4eAxrKb2IYYc74z8M499W8WMikh9I+uks4BXCZfjruvbS1gg
F+uAhnz/PoWrlygFFXx8/Mj7fYCONmL7goeyY0xQZNybRldJV/cdmpW0UnkICZH3
dy3ztIxy7eN8icy/w8AbnSLEZe+ss8YP6+feNrSpLLb/xXQ2KTs7m1tu1jwItHa4
qthvbWyYSzJnwjRx9Uq8hEWraGKOXQGd5/0jDKrF+mcMrXbh3c7hhnsAZfplzWXM
U6ZgNVr1fx1d1pR15YvSCZVJnb6P7TFNHMqOmTWQj8+7ja7eVx7cH1veT0Vx6Qtl
FvqIX8H0HlUrM9Xpk6U0Ew/nEd9hFrZnIJUu7+Ra6rTX8TkbFxwFNu704KPYqmeW
Rcer+F7GDLYHqyBRXAf9O/ZPpLaeukx6H6L7gf1tuGe0ShLKTp97q0/FgFcfaKqz
oaIZh1bMXlw+wjLOi6wmzuJruocitBc5Zv2ldBuOZv9x5NrXOrnkMxPT7wNmUEz+
/6HDcrEgqM/yDiU6w4tDRJqCpxs/flWML82nSqjaq9ZRIcQotFb6Si+A6D/R4yYq
i8sBkjFtOEPpEglgAmlSZorV99rGE2CWrCqmypfetCcrL8ZEREIgKnR671T4DKOj
KnE3yRp2yYw1JlbHWLM1GpyF9eLU4GgwgvJ9na7f7ezhNaPaIVRYLJ1iIhybz6yZ
xJZwVoxC1lLSvIZdyOEUafeXXjCuumIisA4m25GLVVjV1CxPk63Ewfu42GF6Lxax
oKs3NxFZLkWvCRbbmZsr/6xV1xTcaBafcdW++cHGWdQT7t1UTGs70pc2acHM7EzR
ZZknOynNm0FlzfKnmcgwTTMtCyDR7B2mbqU7oc8s0w/S3zvvc6myNtGs/sV65HoC
HrR+DTPK8y+Oz0oCModOV8SUQuBYtjIxbshSyEzUh8Bh7KlCqLOVz21c2McE/NGY
bpgzj+DmgBIeYh3MJUr7AEUXuCXcHRAs0MGichyOfjonLxQA7EoWaszDnLT8A14j
C5CDGdmvt+DCkVbRCdlnGKsTdY4XEG9tLy+OB//kfX47sulPxG+wW+rZR9X382E5
UPFPdAKclfestqNZ7MDGLsCs7pZOrUplp9NXV9J2TdO/vAxUff6D5zILUAJ7kTk+
57pc2yzE3GWAcTNHpomBvR1kHionXhs9e5GjFIuvDH4f2Uk4uece3nIh6YJ0z4TW
jtUJfm0PEgpbyGrx4Im9ef9jsV7S7qPGiVt3TlluzWZaR6ZO8gPIytbpTvhCUVZG
ikRAYT5+u2e6N4cHG5fS5OgngFVkPVSYoHpKmSFGd+qOnt+0EtPoLyGMGmnv1Ojk
DO8IvIRSKsbZWTHgkHSrzGALgqDNXovHcmv3ZbpIc9IZkWfguaoFOXS4B/JXNsTU
tLXbjxQRqSI2Uala5qrA2OpLskYMnruDO5aQQqeS0cshqgLhExIpvJXEqmIh+wYI
BT1JyjKKGL6Su2F3ug5lyRqMuR4wtjJr89GuliY4YiNwn8IEQp/thiEcMQrwPwZP
HIZVTZKssOLnekRVdAErZ6XWBZjBA4OaJ67JBN1CvK85PYpR60a9ujiirV5WWJif
SNdcNPTnRNIXet2jxJ47ARX3UbOpGDt1ShjQZTK4CuF4MDn7avUFjUsOopB0d3VM
9+oaMJS9KAdf70pyZBdmFHx5OkN5kZcsphzyBgFAVq3b6mN0ivU7tflk9pKDci0P
V7909rOtXqb1zjOlk3uEchYk1tLl/oJcO6wI/ffJLEWObs4uu9IYE3t3v6xGsViF
KwBForKNl8/glTBqWTZFh7UnYYbnWRdgVqiHBBUVXzhWMbEtA86Wm//GlcvhF4AP
5fiX1p/cADSixl7cf0KIBkx3591Vc9SjEDyxzBJjDbkPTmgrFmn/G+MXNKjGDiHV
5q0gr347oZVsJ9iuqeGa9xHWOeG/6e4r7tbnC8OmARLBkYaHlh55uEisc8ewKQI/
inYGsOIq89B6x5Nihs4wieXUWrj03i/8vWX1OId5E6J+Y1erlowdJcyzDMpdZVSl
/Olq8umnsWUGcWjt7aaWQ9JcLFKFwXsZr2bABaKOjkIsuZGdoCaN+JtoN0wVrzjX
P7Y0u7vLl/69OhdwZgWxRQooiBCqLjJGJksiySAh8pwT2yCX/BgCHO0fyxwTl5Mk
yn+70EoCATBs1Mz7nSlmBglKDijLkz7Hn1imRgKxhfkNGJyFfzjIOT1oIly8462T
xmyb8/dmtJYSX1sxdkdVxr7+rmzAJJUSLh6hnCOrdDHGeFG5Nxam4bHfq6PfeeBy
yKRrWLoXxjzm7vmcLH6pdpW0EZhD50zHt6HG9tE2hMYnjbc3lda5ne13vDRmX6kN
6pUJeUiAO3XaF0PJFSdEq9rFP7RQOrcbSK24vPQs0Z8+GifknQHgHOa3Lo1/7vs0
fRGmjIrHrZoWhrenXtDIAS1yAeYerLMJmEhELW/UaNPX1UVPw6gInWDpgx93jNtU
UOJmvLi2naD0Nlye9B7fed/xd+lF7CC50JKPZce4PBAS1MFM6z+QjBYdjUNWsEyD
zzq4kFt50bZh9qyMHQ6wdiTZW0hIWAsySIB52rNMXhvKr7Le2qaKWfXABDeLlVsc
dKnNFnmxdXlbw5mXp5rl1Y9VV8Cdfd6Irrbm/onybIhSfZ0JBRVUSKJqg84p4/SP
JIAMTvL2Vks30rCXglqAQFm5InLH0QwB01ek7c/4ZUpaicbM+kE2IGXXzjp2DGZH
O/j4TuI9B2QQXvZAaoVPgUkefx8aHqzw7TR2nhj6T6ZCFdR6TCVx1na8+7GRHiex
gAZExtn4qkyJsuk/ubvfE2HXJZ8dI554f7MURxCrSC5Zvkzp3UIRq7bBO7ldyP+X
8BHjQG6Zt5x/vMLSENdRsDRfckiBAOwn0cbIsaw+Vm8eIjlQ7+R3SXdZpg0fRLF3
LshLu8tDZf91lcKYakvzHBkece0rE2Mhm/7P7BJex5xaMCCe0rsdGdzFgKfW5+bB
WwkY8F7C/zTzZzHQBMuWoP2UYVVuUxO6MgjGVm0ChAPB8H+iXD3sG+/SHRnLWUcS
jrXn8C4u9k7JUyvnJWxIUF+44aEHaV62nwLl+Qm/tf3WIH8i/iRykoEb7+XYX3az
S16b/aYQHETw1f6/ocb4ws7xEbaWanfFaw9pSmI/E5ErZzdl7xc6YJ6N/au666IJ
jmDnJU4BRr5hHJpLjOcQ47gdggPdXkLqhwpOg+03HYAlBNpk2HVfueQd3xzEvdHt
CCbkGx+OL6RbUoN2RQ1IaoTvfFopQPQKEKnZ7EKoHhnOe5qua92p3Mh21gyvyKCF
LeEtXeyGc05k7LHDb7yJ/Y4NEPGTsTUwV8EM02qVT5mjFUl9QeSMN6goqLlu8Ynq
RdJBECfBrSAneMKOZSBjb6lhewkhPDdiR6wQn96TESzTDohw66NWudLKLueLN+ut
ScpWHBiq8VwjqaDibSEUkQ6eaH9f2VFqyqg9kStmq9HlotRCBWNJRVSZ/q32c0cp
Dq1QlV5FtAxAPF9hhSVT5wkxEXAOiD1bhKxG5Qp2jVe8bGxW5+U8hkcZzojR02aI
0zlVcI/o4Dh3kBFZ6/LhtJFzLWJ+DRXQzWYZPkzr1UM5avrglj7Do+1D8HeDqmMJ
vPa27ljr6O14FDjFaV+iDCksCMljyTaq3Uu4g++MGbREwFS/kbX7Xsvb6FF+WivD
xgh3URvfb25ghDZWWXIy8hTQoDJY1Gcfamosf9xyOGzLONGc4ZFZorxrvh7PdSNG
QI8r+hMFYfI2ptiJUu8k3+6kYrWBowdhmuFZg6MM6fNQ1w7cs8DHt0wSsWUtp59E
cTt4txKoh1y7BUYnz35MxPhJ5s6E5mrjJ7wyun4DorfCdelc8pUh9dAeYLVIbwTK
0aToRGqpEv4u7J7fcT0Zt2pAKxHzLd2fXfGpmjpx2litnG0C7VdlgqM7M2lWoUk3
qRn/i2ZlCCvhZ169AKezUrbnQ2jAcGtJgAuCPedJHQxkzBJoeoKfappYCbxBG2cu
cSdzbA7h2XDCZirJLbSJZoiHuUeTr0AhhxqLVMocgp9uiHrD9yN4P2Pwn30RmDnG
+RosR9Mjdvj76kYm/HRbrJbYFJEQ2LULE38fw+KMXfdBooQnagn/SkayQd7MitQG
WJeWxWN3cFe96YOBNoJIjdrwL6WMawxUIQQv/17rCHmlTqCsxffsV2ujqrqUrHDv
3cJE/G7pQHtdRG25PtOg84BkcjMwzUoSxPkQ+RWK5KTqCqE8kHTaZnrq6oOgt/7p
2QUuMVbI4OuUz6BfMld1zY8RzEzm7lxfHT6BM4ZaZ6xnQbSLOjUWB5ZI2jQ80Jf/
IUyfyg6LIApbHxukp7lKgTFiJsKOXRb5bpTIHh3i5kp5RKCWPVdQtNZ4sSKG9/4v
G7jJhh9uIDdVc/tyzkBiP+HmddVXL+ywfNjaI8bnRqLiUhTmUnN3wRowgfnfnJ74
F0Nzyql/s0U8P4g2/jAD+j936Gz/ur1u+qsgLmvuRFHA1ftRAauYPAuGpK5kYqME
TxNwOWQrnPEQUZVqpeEKuxlNA4XTMoN1Z6Qx0Rare8qnUyWxfUTEXFgaNLHsFI4D
ghLSLys6D92vtly+z90vFlZJ1eM89Qzgu5pSwO7eBhU/nuiALj7eqHwjH15X+Ag7
lVbquS69yYvv6Ln6uxDtHGvlAfagGH41GMPNX7Y8q2ET8dH9STV4uoGxYWi5ZbPS
s+kyBnTZ7FEI+TIrSa2VkZRzz9+4P+ULi2KRNepuQlYO+xFGjvocIja4nFLWhsNq
OyVPprHPyDNSudhpBGFy4iI8EChXIOu6BV3q12iceYLCyLarWYpXyVZGZUj1tM6q
0UPQxgc6XIktI4P3fN0wh5o6vnmK0TKY/z4Prttp/4+XxeN2Z41WtY6zw3yBNTmR
uSFSQJnUjbOGcWCvmgpOZVZvThBegJmzGHaq6OEwRc96wdo1yR3xqjbCXyKCtVlh
LCeLJmWvThjnoCCnAFfr16RjR4M6MBvWn+1OMD+C7Q9ZjStN7rOF7jRkAt+qeHDf
syK/bnFUMLTHxjYzRcPLeQwn+3CQsIp6BBHHv2DeNGxyNghY93J8L0Gi9ubE7vaP
fEaJvCJ/j0yCiXwlNA1UsDohU5VW8x3JUlu2S1nnwBfCdLXkOoU6Le9Y4v/aAFcN
+tVTDi+Q2vUT7U2feTr87goyYY3QDwAjs7dYwqr43Bg3Lmuc8qqfqfwCpQNZvjAu
BNi/7o2cdQnkMC487hcdTTqtBUjJb4qtDToxYo4G5xK4E8Wv+onF7Applv2YPp6N
zjnB09oJZvfAKnP6icKTFSY5OmKye9ARVd2d8VPYzuFLmwYUK8p7DtfI2GTR8XHo
aahsxspmTH/ZGoF7TFhXcCHs+amTuUtpPRc8t1lMoEbSxUrulnQisvNW3u692FfQ
fRKbh87lPU/JTQ7O9d6/GDthBa+d2rEJiXMwHbqeQqgyfZDr2h5mnBenQloe54gW
oejoQRqQwAm6KEaHW4MgGVsUj1+NSyzLQVra9+XGSskBZs1LUBeQhhfm+bVjKicz
Gl8gS6DOoiTU4YlIxkihKk1lvx8g0tjXQLFgWGYZbNL+yk2uLvMki3J/MYsTLDrP
iNzA8gOdASNHe5yMxwX07qTOsbWgWtZa+TPTrDRTF7WBheayo+52I8Z7LJDHUe9V
b9BtzhYWJD70EcwIKAEZeJ6R8yqsmJutV7eUEYUkrjkQILeAH73jLuqeoV4gosXh
BPm027ddg7w4mQ9/4sF8BqKfZ5FWgZH0e3iDc1A2a8wb/NCWObC4n8uF4HinHQH0
T6zW3unX7cZxYTgR1WhjtQSCmJ3/CbfMAhDMTP+NBcZEPNp9XrC9Q87ZRT7ouybd
qluxbR1hPOIOsprOmk+bDuIjil/rWG1U+XY5ekYu8DKVxV3XU38dWuxDtyqaVb1X
DbgoTsTMyxbEb1p5xg9IEO+tDWsZM/yEIrs2Whh+z7UT2VCEP3dWLLWHUeQ1YPuu
o7CMmDtnKHLqy8c4ISBJmpXNDKGkvd1JSeR4S48i1gHkzHbTQas6bGfB8yILsEbI
Gt+caqJWvRDcTeWVfv8u0J4+zbPTBBN6q6fKOfIQMExTfUlTgOGqxc9CNmqsoXYH
1Ss653xZ+MQvc24eupGO4gGFvutbw+0T+ZGFO0Akl5+4lpcgBG1fDxF0yqdCEvig
0CIdHVC8bvVkq1AEgVxd3HReRMJ9IBE/qtXZKhXEuCjaK3v0C6jVyNZYZkQjuRHB
gTxBrbWwEjuoODFNjqeHhLURpDL8cSf9pP5gBUJFwiVaKEO/IJjSJqWNpGJnJcm1
5AqFmjFSLL1DaKb6c5qHwV5f5qLixzrRzhA/MXVhyKlvpZGAYPsiwWqrnd0an3h1
Iqy9R9PRDBuyQaBLX9x8RRRaxMTgd8wQLCSj5sMJwpi4mCIS2GKMMGGjrUtaVJai
A1FFLxIpbw2e0K6U1wBGmXDgkScyCIty5LG1yJMDM90heZYrpsRjHYV+qN4ealt4
nPDQSk8H1X3DITUst+OiuzlxJiAZOeKowBH8t1VQO6YaHM/gz7hNDyFXdWf1oeH9
MXUpr564iYFNFl6CtEK9JCkLJEdQ5XyFYBLFD/BLXKV7X68Mbd0OrDVcy8SO//Jj
UorCeQrudpB6fx1QR49MXrwyprFI3tkJ+9uFpO/tCuBGbiL0vnj3G/T6bcTfGkZV
jknN6JGZMsosQNRzhSpHpTZOzaMfp3q+49EbO+o+9KJ3i2wCu5/hyk+R6ExJJJDV
y4xuPAYBHaqxu9HGZuUOzLCYbnEbewbufK4IjTMq3b7kQ2fRDi++WYUkkwvv90Lb
I9x/0U7SSsafqNgUR+XSn7w8QLQkDGdXbO1rol/PAJbyOZg+wYBkwrg7LRZHo2Nq
V2Kb86vVaQpB7nzsjMyHuWUTvMZCO989IuJugvzEgLRC2OdQv93PRt80kdOMKYeI
jYgFDWxHCy+YnNLfeXhPgXvGN2wZNVktc8Z0VQrQmF6rKGT426iLQVpY5EJg56WA
2+qSP0gEWH7S7oKHDIovUMUo8VE9XaU01VXHfff9XLADukfcMf8RKoMgSRECbbca
edxutGYY+SQ6cXOzsVk11SWMixRQoUKL3WcGA0gUDg1ysNRUTF30sC0rNPPSyV7N
eQPZwoDqKayTpq0zmAzxGmS7JGffu+6X7Myz729r545+C9sCGzn1kRj4HNLtXenc
tZqO++hAv36ncCaIzRo8VMP1NkgnTsX9lgPT8ZuTX0RxpAGFxAHCRm3bWu3VVVa6
JdZFzD4OKsJZq+yiLIzeLG/xlAEKqHIawu6w1VBIuYK3/Rs7X3nd0Zep5Z+52RAv
4J0VnDUEUfPzjrL9fz8CL3JmcoV9SubMDyqd/G21OpLYhvre6NgJ2NmKpJy0b5iW
WQfxn1l6k4TN5fN/m3FAMEbgeL1U7Q0oSAbV71EJWbsdktY+AT0Y6o/Dgnf1z5ik
8QeXjASC9Z46/7sJdRugnFqzbKpSNt/PtWP+Ryz/c/ZTmHwpSz3/01Ey21JcZxRq
FmBxabZB5Z5exp0Fzl3+gV79/L1k7gRPkjU3o4ZswMwTban6lHgz5Sy09I4+LThK
OdpcFhsBqdRaT6teYpwRVslnVx7Y0+Xr6JCpfELpsazSWWFjeqIM4HAxWhHRGuNk
uG79YPe6/sXrAAI7QW++l3SnCO/R5/epYyFLto8crL2W0Mf9SBORYowa3LEHb5mQ
l3u3R4RkNns+sWnp0z+jRvHP8B4BIp4OQBT0jB35ayYUgzoLODokk6LHu/vmGOQl
GMtsN1O7htBVHmFFsdL8v5kh6rYt9si6SzptLty7Uc1TYwAgvQyXdVSvS8P8mqZz
wZXirxrOWB+oRTeRxG7wkEKvVZUyqD3SiKPQmWW9P7RpUjmB2Y83xBX1JDo4dJsg
Agp0eJIzug3pdu0sbAUvLf/miCWFDAEVEgHuzrYOOmWR1iI/GjHVqTHHtQIsVXvv
sFTAPCv6cJRrImQauQlyw+LGkFgES4oRx1j1kq16ZB8rlDHhP4B2JfcXs5QyvhRm
m5p1ZqbEraOCoT6dCDlAt9LaqmPxjTzg72xIiRgCBbNKWcSGnHbDTyAuFSQc73e5
oZYI4D/KCc/3l2rU0ocXG+9xe2gfdqXKtpl/Yp+eLw6AMG51A5MA4tbRd8qkroEl
iqr9A+5UyiFkU8By/U/F6VMdTbADWHZC/52//AF5zTSVKXbyqDuIdrcoJwtsgEzn
bttMAfn6oVFjhuKczx7hcAMkQYfykI55s4RFpEBmn3tKFkS7fExSd2KtlrBr9gOm
GTfPxDaIlj/qOOIa8+Irr4jsUsZjBglMhVGc24aTGoM99RwrpFV1fkoVfcYxamK5
Rg5lqRl2ovblmDgOEDnihpFFzeg9q8qcs45Q8b2NYBYNcdia+xH/s4xqOGxEk7ul
PEJBTXx0asghjoul5NHlZoQNw6mRJuqSSc4mSkqOaJsl9SIRJugliKVtFQ1w7sxU
llK0y0Nj/qH43A0Gj+qSVqwgjZzqycoYmaCzVfHUBhw+o8DCcPdvqBzIMIaQbeQN
VZE5J8Aifhwkuys/d1PYwf1edkAeCEfmLJ7F9lNK/X/Rx08BRvAzRoLsNC36xCow
R5smCaxMZBluBbWC4305/3pKqAQStZULSaH/6aEoP2ePrXtpLOh6tEnTCLMQgzEM
mXp1Mqq8vplBGB0+bpF6OJPoUMPJ4BW6v11olJaU9NUxZnUQt6PROhOX4Lc6D4le
M8zG+RVL0pKpEfj8vXUgAVzIUt/ClUBmvqQpm0Hh1N521R9Pz+o3yXGIA8Cj+U9r
/e2lHkomDDB6t64S7uUQSqmu+eRZkveZDPLAVwRCtY+OATT3iGocQ+CS0pH3+Tpy
8PMeWsD5UQ3LGl9KCbwF/1zk5SRjDSHbk12hd6vdqxSjrfROK712R1I/0R8kYvui
u5zrqKpZ3Nk3NIXf3UpzXyNhZEeyushDnuVnbninLcc5fKjcmlMW/rmJvoYf4tCn
RNADY+0TW5IMk+2qhcvevpgZrlC0raejQAFdhuFEvsAnuhmRTx3Z0br4SaPVf/Y0
JLNzt6RmtgmVDUy/ct14SmAO8U7SLszeHj41pk4JYHFai89eBHdWZMwKoJhlQWbo
6wMTF2VXM8aypVuFsJEKDb0N8KLj7uYtvPWyO52bqw5yXWxZVh9vvSCdZOsQbTzm
exhD0hGHwisrgUhiwr42CGfB07raLhxBqa2HA7UKY2UEy1StczxRHm9hzs+abqYw
rmF1RYV82K4tRRcLxGg4fBfatBeZDDi1j2OclLcNRa1W++FuCuF29gjZ1HBTFX9W
OWTPU/h8bPHF8aJ6yJGjHaGHYNPs0vHlGiHWDizGJ9V6yyxEyAKFrDGXZvJFusF+
UUytNSqJ+bZMSQaIAYVaL4mYVvmX7eXKD2X54goW/+vcoHAKoILzvnOD9RoaCML1
Z17gMq7os3ip0t748fY9V1z5frAsPx1i4h17bY1f8YLQmIoZlP7sC9RRQ+3q3Olr
gaX1UHYUdHeDvXmNOqckHEZxPN9M0FxM2EbZU1dK26RSZETutOJUEJ/TgeiYo5Fm
LkgbCew2/aGO6JaZ8e4J62g/epTVZy4Zy2H86vOzakS/mdQ5r3MjVaE0vuMyj9ML
P54+YK/H5/dzBgfyKZkk5+BZmz1oaSphI4AQpfMAunK9E0leHN+u+9MIiI+LRsrq
PQI8axB3OM1c86y9LTPSOJjMfD1e03B7SHqHoffOeKyKxx6Qm+HmONuyp4c21nFi
jx50qRJlujfGYEg8fcaocN2cyjlA+QdKVP5a80icmk/gCkXyfUvTrExrokIa/hKX
4M3e2sfkjhpvarVJYdxHVatRIp2yRiGDYqfm+qTjodtgbfhlumRPW/G/nKx+dOBT
vuyBS3GylvdLGGhzw7ZepRIs0SbZNhRn0dS2HVYSSnErvpmRZ+31ec/d93bTNJY2
ovBgWmDAY2w6d/4H5BWJO0jQxqudtFKE7cKskUP5PxDlunDpjl2x+s3q0oW82fxf
NQ0jf8LsuOIsMp5LKDuleAOSl4v5RA8Fq8MQA3/LbKB+uxJ43IHm1VxUMsbv7yTR
fUOe3w54relIdXrvaEopkf9gINPtmok6aI2azp7Gl8xAFNoSndCB4ebAp7YtTJGq
EMunmjs0qOFUARPbA4B6emtIpnkneCvyiGtp2WQxR+k1tv953maCo3lyALuVWv3G
ll4QWT3HvbkOVNU4keAx2Eu9kH891iuKVLLoyT7x80n89axUurXAMz6Ls0t6Tw5I
EcojbKvesW84t+Z4Rsu6yH/ujUeb1H3ifBs5Wqg6OIROTcC2FSYqkQy/OPax5lOk
hYjm6AgK4cIaioAWsPP//1FLHMR9wBEVy8RBL6zqrD4vg4sP3E1XMlpbeKQD89Vn
X83kxfCUlvVjCHwffIDXcqCTZyzSOk8NDfsXoNNj3SlAa61+i+ZTqrrVzvf9P56/
aneMwV7LaP30IGvIHi73odzW7dVOedWaWlLhBP6h1GCzgwlFIJGGL1RbQM1BtEMz
Zhr0fDTv9EpgPaotyYbMAej3lsqZ3UmXeV7XOHmUqnELf734qo2Ejhc8IH1XubHZ
XUzL9Y35oL+zsncBCBoPw8XFIzDYrFojb04lAF1o6qilmSP0cEk40fNPUke31Qll
m33LHXYTOlqc9VBdBj/8EgOTKo1Vh1U6YOEkaB8dZizvAPa4ryg3yqiRcNHgF50C
uJgPLdIF5yoj40HEN7d4IV3pM1ztL5hCvt0WAeKyOCzgyXR2v1Yzzca01Hz6l2c5
jCRCvO8jXxm8BMuquQez3WZGgCM5xX5GOrTjjlPbAFTxgztr9+SCBSKMn/O2Xtk4
ocKtxM2d+TWBlgJrM+iNDGoG+DwOSsC99kdR+VzeHi/NPB9O2qvQT5IjNDCND9o3
YDyzRGm02S17vWBGKxN8gXeX9T0BKbqJD8DA+8p7wpwZlU5aQXs6OR2baIEU7Ipx
6eC15TnTu8uD+JMq1rR1VgeHoMcOYPRT4DL5N1jy+QN4Z0GRYxpe179Uv2LPshzb
OI3b8DyQf0nLL9KgvuTE2TXQ76dxkbQU3zI2rOAd0BjUWH+nhmUFjSjWFVeGSUsN
4lPF1isZOGUr9SGP5Ho4h5SUi/cCnnOyCMh60D+bIX/4KGJmhG91NuExON3kWc+O
jk7gOgEslIyt49bDiDF5WqCE6QEHuBDgaf0TYQYoQiydZ0Ojy3y6TbWwxnQfG31u
T9T1cniUA/E58onrr07GkpXbNIWQ2AM+pFFEtEdinJNMNWx2T3/ztbAmua989N4q
fNxrw/jE53FryAldp5T0x3HdD820FpUucry0ATGlJkIJGGbRaoj3zwIH2EsDZE9r
bjSAyysp37hvPum4XvSEhFCjh9Ok6nqgUvxgdK/pEzGfmhoT7hfHNjiNu9JQZdGK
rbbsQcm7grDZ7RTR7ovBZxCYI8rZFArWBjHOaJoovPPYbvk2DjMqmZerY8vO3Vrb
bSFpZ4RtrrHXHIGle48iztZ6AH7rLpewt3AxPjalqxliEIwxG+46/uIDDYo7+U1f
1oFEWVDhBr4JAwHKvygPcDQHN6985bhaL1TDAAXHFLG1TcpJDh8OzTM3Wupcxh/8
7qqR1C8Pxz5tEu3JxK8qt0E8z1S70/HEd3DdJnG4dRzVi/QY34W3KGs7cKp1GEbv
TkP9jnBhljXqV4+ru2HNuCjS//fVHS2hi6xqTIWhGlGKCETV80V+HuH7Xid9qf4p
uIIB9uOT/ZPHOSZZ7pmYfRfLSye+RI2AniUa/fTsqviFdoYjyUdeBX6K/vxOsQ4+
eCZwjq1lqlKuqmBU5ed57keXGqMNqq6OpanT2iV0VyXxqGx7tYjISYySkz3ZdiHK
8cNASDjSnXwozcBGQDbfFEbQ/yep6SChza9TCYGJIeiEvAd2sKpyAJxw96YydfK8
nigR9CAFYIESo8RccrsnbUB7ZQY43x0rY26SVjmOQLmA7r1EavAhNyd5abUmcWM1
7+28+mTz7AxoFq6me8LF5fTwdnxcXnJGOD2/ko7lDea9rmJR6fHVnvFliriDdq4u
e7wePHPpezJAuN2jPz48G6Su7gCzUrnJvLpmlwQ/9ERHumSKw9VMHpik0mRr9MAI
NUX3vdJg1Of8E3oFhaTkAONENCeYCdg4xRkOlY8WZt7c15v+MA1OPaqLDeKOAWej
V1m8TxBBtksbrvWV8JMu4NgPJ7ZwtTMD9qgqWCL/7I6CGntq/i2kODsL/x2DBzdS
atwNdaBkLchDuzZLUDvFVY2ieJqKDro1ddOJONDw0tuOxGpRXXQia/3rTCiiLGKA
b2N/h9qSXINFVxvqfb8XkswppMCBVe+sKO6QlmMQP9llo0iC8jPJ4f0Mr1cjLxdF
HvlVYr+jD9ClkSP9Q7gZ0lrfy1p8bJbFAx+uEMYvojQyNeMPi1DSR5ZCixDcacc+
h74MBuP4R3/1Q6IIyrimEFL2a1ttM2wMt+3OWcNyIU/2GEsDITEhZgXKJB2TynAF
oRPljs2uAfocAfNS4ga5oA/PD+08F1SkK+ziZQoF4KTWmgfTg21m0yxsmE5fQYRk
xs5h5XOK45WI7csAzbzY5ZzuAHswkX6X2/RFV3q3Vos9HjL+Czw2z4BsfM03x5WZ
d5evZ17VY5A8nsjNVfPlghf5kOq6QhYG+JU5ePbP5qn9wUZdqMdszufQsK+F56+l
U6FuH7kKAFf/nUUrck91D9MuFXyWDpx5SnvZ39N4OBmkUt9OYqJc6v0Xt0J4RwFf
mV92ZVKRRUC/6EcvN61CtfUis70hLcN9yRZxtN7Z0sAvnDz4YF7XtBfrGI2IFXap
2QL387eHCdHsbGWbxNLK48migla3HrF86c09m8j/rQGR22QUPB8DF0NucCtsC91J
jA9Z8SL6mwFaOXmieR2uP1i8WmrMBwm4cmecA3ILgJit22dTgGxgvNlHLtUY8kyn
biNOjUnJ/ShZDw3Hz03vAHPe/rPe5Xo/lZhxkTEnqPh4xKwVyr2jUSaJ9zJ7Fq8f
q4E55xWsHW1FOqCwJHI77VJZrg31m+qqK3JSmt2jMP2DBEhOaophGLIWoIcBbw2a
LDBIm9118LwLpWKqLzrSd4AwF6P0od5xS9ZKL9M+kY1uqWJRyGVrouRc2AHfSxg/
G5CSGxwSHjdI20NjVfLZtMoui6IDUGUbAzPh0mQEfaqVtBhrvyUgaOvvD+tbBFtx
IwRo6WucC69F2+LmtkGE+O/NtEclF2QRS5IZqKqP7ZhfG8tqjyB9XW7KcTJtPkgs
bdfVp9uF794feCdXFP/yuzrlDvMH9nieG13rAaLDZY9xx3mlexJ0IsrYmV7+pZNg
Y10StynQgTvzuw11KEraFgcZf5KmgcQjHDhKDESM5XLCraTSMZyvahdpoMb2bgrK
26igZB35adx2RZjVOHHEFSA9KAzQd2Sh1VxVoz6i+X/AvwZDBG6NpMhNTn+CEdrW
6J+XJEHc0TVst/3zhei90+CIg+f7fF4nCNirlisJwz33dcWleAkiJblRe+vfEsRz
BUkgIo+ZouXJTTGgSTGCORSfKeYyl3MGw0fB6jiE03sihMHTeTrqSgYc8UBGarP/
rj9LWKeTcAHV0HQUdK+ypNNpLWBSwQKi43TDNAb2mhimOGLhncoHaYn/p4/rUvby
2SNaXoX74NiABS3omM9B4r/DE+dT5F8z/VGb8jdw+P+fg80PzeIgn7K+hXBgoOGx
9wIN0R0Y6ZGa8Z6Qc131/zTSzjKs9ds6YGbweT3MPJdmF9KM7ouGDrsiRxiBG1Yr
iV9gHQhF/kH8OQjFYD/53EFAsYL0rht1j2x72vJLzDntkmd2GrQpyaU0KxST8+pT
XTzs1UnLrZ29Gr4fpXjcHKeSGFKNPsLb+RR5RdgKpERf0bsvgvDBqL8AgsSnWy9j
p+8FV/IpMHDDiIcC/oZB4XgEFy0jgXHhg5jlUkC8/98snE1ywwVHX7T5ndNSUgfv
T803qBcometttByqoayMGEXf5DkwvBeKRSea8xRTdK548eSCELPmNLwwpaZPedWb
vyFPIYVfiEaoSUrb1xZdRDt1TLiQ8R6mRcoq/lz/VEOcFwPPTm+oi1vmzJfL4D+F
C7pFudU/VMtUwqdDjYuF5+Lr/MHKYrsT0kdrUyfK1sqQj6UIJ+rf2KN8/F3HaL0i
Z4BCzKc+4mH8WU3mdM2+sl7xUYZV6vS9qBRGScvxV/oxkFXgrKs0lokedTzh63MW
bgKq9oUt9MyA/TBYBNn58AuGaZDin6PQ8lezuvDNadq/lz7nLXXbMVHKsIEc6uT5
lb1qGDyFglr9O3wiu0mH8YdpNhqvBiyxchNwnVzOQ/f7LmweynL7DmA/gs3YZFdP
nHDd90FUKLHOwt+wPI5/edP73Uy+2r9nsL8tZ/pdh5QS4on4CSV8eOuGhpCmxcIL
bxZ7101ikfHXoDMoqluV7W9thGN7V/Cvuf3ADX2o60goPU6hmmy/Wtrf+Oy9R+Wd
ixJ9SDzElTNEPcPmNvuUVDbIb6WH/FkWkDyYilN5nRWNWACMG0mn3fGJydNdosZx
YpHCOjOAFW2l7DP5p+cf3VBRrzoy92772Qd0OfYytPKoz6q2/Zl2I4wizZfcy+WJ
Suan6kEsr+2x1fcgf02goEGZDCadQV9HMEAPffPL7FbM3PIyTSwxwTjgxKBSclGx
RvUU5BcGLPzECms+IA9SvQm3FS2uCdm+Hr43ZzVrAAJlgFyNFj3QOIBd+yNtaiaG
c+MpB1L86J3xXSVRGM0Wk2hA361YSAiSGAZKKGotAJPSdYfyKYzlzMScS6gtODrh
pfuA5p+rF5LgvWJ3lQeGVk6oZbgmVu3Uhdz2xGy6yC+u2X1s+/NaNM1yRVIPLCSP
eOmN+tBHSglM/lr1hEylCBw/8zjGzresQGugX6Qy0fLJeehCQJiKHKle2Ne7WoI9
WyhDAOOM/iVwyKZknTniuDDVuC8y3wDbl8uiCGOw4P+3H3R7lv/MqkWF/XxCb59M
+FaoKVnBsK/XtZvcRLrJq3kTlXUB2n8LU1SRJtOjidHg6YS/HsTmyjLnW2pgbr7g
LwCSHojY1c5cSoLQdWw7Ym7QqC11zYlhp9VJa/wO0ebOAZU5rhLEp4L6cmyqQV1s
dy738KxUPtRRpDCAilMZ9ozDzI+R8HtkG0I/kb3kUzcJHs2IAN5qj+Y/Ta0w97kD
v6yoGdNCqUpyseKY2POHJz1XF3VTPUMR3IC6FLODqJW3JoMVwM5UGCPObBw4b4Tc
gpBhkwZaXIAmxpRqp0MkrWKyQOdlu2zl2NX8magK7ebsuF6d7Y6v3mswmLnWRhVF
BEQP5EAGbD1Iv/WXlZlLjs90f14suZkyU6+fqkRFWZwFmL9nAp7kvK1EbA0A0K7w
PGUMqKXH4xlYvuF5MNmzljDDl2Srifa1dxWVLF91ykPOZOg9XBc2nAkvFk8wDH7g
4q8StgAFezDnd55cN+PEh7s21Mc0Cw8hr4kemAS6I5JuJrd8F7ysDjdlyThv2/Jb
ZJaj/qUwMxqw6qSD0RA/WqZitWqhL6US4OtC4d/lg4acK1KZCUtQYFIuQyHiLLGB
fppgzYbL9S1YpqnZf9V6hKlpsvQpZTDpxki5MxP3GURnee97SGye8xcFd0ldjOvC
pOLrP+ohFTFuTUdgubgfGf11QgCG0Mg29Ua7+VKGlXTvjwpg1zA2/BtNAsgSsoFV
R8dYlDUkPRNJUeqfB7Qt8SB6V8Rl5pxjF0gtfa9CNBNAf2Lguj6PyCEPx/KGPk2q
kNXajQlcVOeCM28arxAVx68TBGJ3wEMOZ9vf1/FenF5GJ2COP+ABdzquQS+yT6Z9
sMVBUEK7Xl02MYZaDNsqMJoUAun3tEG/+fsWEeurVs23KhXKGfuNsVZeb+waqNA6
bT1qjPy6uxM3OQ/+BHuIAYF8X3g/RSJ5Wh2jsgkRuQZcmND18U7DLpEdJOwpNH/v
4R/SvZ5UNlNtk8IVi0jxTPcOExnlhNMOzU6eFNXTbQMELhLcLFmy4VhyiUBy6dXi
3Hn7IuNftJhNowiXvKQck4NBNMuzisqbARfIzNIb/xa4ToP1IJ1PDCoDzCCcmCzk
v/og2TrzNioJsWYr8+9SE8WgBlnclHRi41rwX74tyQe9CORXdYeYm6jwAwM2Bs6f
/6e4Ls7y6FCCKFeuipQ4JZAMLRfu2xNc3rn6LkDW3E6Q9heBvNOmFhg4ndumFThr
+M7rKNqca+LQfiFUV8FkOZCDoYS4kaYdNRn31pV6BpU3o5guKJkdc3HQIAZXHDiJ
KXQW3ba9aqlQ0gSqpzUydYQFE77aBQHJuUkmPC6YpjgLwUurzmNpwnQdXLCuyiMf
3xINMfAEfCAYEjsTfMgOiu52s4WiRElcscJc1FKn2XvyCigx50YXcJGhGWxXlAUG
Y4Omeir0NQp4VMHGKcwraMUuTeSKkUdMRMmVwIluuQkYbyoCeZ5q5g1YiPtoE9iT
X7t1ZlJubqX/J8/IzfzYzrKrFdW2tsPfl8iIZLwsWGP/432A5gu9TjdfjVgy84Vl
R5XOzTO/gDDgTpGl5UgFwUY4Agh9Qrzwekr4l+Hrfs1JBegClS0UHqpXo3x2ENFz
uBxaoIhU8WtW00T84yYolIOjP2TRBuucAFeKLBoNTitjFYydStYWcfdxXZTREY6Q
v1sbSxeZfRJJSpyfgH2OgZOdvhqn5EVgF+ky+/kCZVOmGzqxbuVzqhsxklwQJUy/
1CTY4wekP5L1k/LHBlKqRltQHV/Wa3J8gJrU2FoAoEJym7vLEhRPxjyr69IzHTMR
8HMclppByqgZGkseKxbEYImiYup4hADYLrrkITSTAADBylxo+KaUc4OY5OpDQ1vm
NitZaupDsqDUqlQ/6FNPymS/1M3U13N+6z89Ha4dkXkCWqi5vFgQqGgihVV3Ob/g
RfJ4CP5EDCNFdRKjcjegX/78oI33FE/IKBYsYV0ymjzPt3STdes3IiJ0prnpQuKP
BOFicRoJhN/m+tOWJmeVqwbLY5sGtopSV2evQ8zH+3wLQY376zdp+HVUOOnTZ/Bd
PNwfYbyYsb6EoPgl1R2HjXwCA75i9U0i8Vg+PFz0R4roncuGTiHyxFo/jnQBjDTK
0W5s+t2sk7w7kz5W9dlNh2z8JtczGDOvX3ahjOsmhMBBaucB4bXJ91zYsZ4nY8MF
eMmHELf3zNJnYR5hr+ZXPyfQNHgF4bXgPz7TSTlQ/k/rIy2Z7MT+EK9ccsvyHLsY
2i1ozA+ag1g0oi6VE8k6NbdpcZDDbLZEIOUpP8ed1hrNag9myruKSad6mzF/glJS
6edXloijXPzzIHJieb21sR7VRJbK1tiyyCFeLNhUpSaSvgS72kdDjxNPJKQYzTX2
r7sPt7BNh1lq1fSYvT9MaySxP6TW6t7DIl/s1zO5UycFSTVgRhmZTW4mVbQFNKk0
25hgi52BKqJRoKoV5NFSQn9G+zR6o1cTod7hHvvKIyNlB4KrlOqiMOYL9Gn+9JT1
8Jw4SLwIrZC31XRpa6fpVH1NEjtQuVhXIhN2QQ8Dm0BOd5Jbp30SHFQpG0irE33h
wlNxiXpDw0YRM9tT5TBJh5+m8piVf/YsNO866niARGLyNKK5QZ4joLTu6ezmCX8f
RsSUJZiXW13pB1fajXKIoF8xq6WZ0wUJQOgw57YhN2vzrgySW1U5s74ucC3QaAel
7URJeJlHHF4WigIOK92anppOsWkd6OA93qjCeIyGrxanMGqcEENRCthbdSUDEtnL
KBwplLTbllKxXgBBxJmV8ByXXMrnP6U3hwwsvdBeFQdgc9UlFIu/gZZk+sIJ207p
Y/lwB9PBXEHHwIbBgtzuBUNTbgGPP1kvQtVRV8Uz98R+HiJJi7M4af2ph+zmAITe
MtOJS+WFmRAUVDk4ApBcAjDgeZyrG4JlyAfdGhVxbUkHy1MbJXVhc6axYGp6D6sK
c5UyZjwcLFPyihN4l1iGSRCuTEN9zfIBGyZVBFesJKGdDeOKgu4qPJ4g6i28IQnR
/J1RXiM5NcYg8QMZyduwE7sGQX2PelM5PxSvEda5hMRnJ+dn3fgK/iEEz+YY67re
kZzpP+TFtvm4Gqm4DoyMg4f82cPb9XqfiguaThaajZDsfQ2M4ZTw3+Kdz0tzR1qd
7ZOr8cSefeeRdJ5d11NtnpcdWxDZw1eiP7zUn2CVhlMsb/6X2RVk2Oq7USYRaRsg
BT2FDHz2PXwkvegLdFv72tWNqNS58Z0wbjE5ZeBx4n+CwsA9vaeQSoFgYkKOnDls
nchtl+BlHO6/1WZ+LQsD2qO0lk5QhNcNyDNcQAU/MT8tzwEeOvSbffbNj7JCOtov
yaA9fqXdzjYEiTGDeKYKU+cge/99aJwb6/5GvRsO0USgz/Zv2xqZQvOnVN5hupfR
8YSjVAuv+f8YQ73i0IveWErDXweLAzsT2QC7qhVQG5bzymyUDEXK/0myU6Ln1lW3
rRhY7dZ+EF5mTulULupFeDCRXIzdOa6M5k+3h1lS61mT6RcIi5b0dHUO0IYSc6Ut
2QEC7JC192bN9UM3t0m5HyVnm5WeKk7ucfiWRSpkiwUXAZkrOggW5kDA7QpM1C6M
pHbX1E473AS5VgNHz6A8GZ/eEN6c0WTvdSYPHsBeumq6RCmljoq5tJJJQD2pfTMG
Ma3yR4Cr6nXG2DGsLavYJYxaQQQ4FpHbDyMN3kEUT73W46Q32/CkNkJJE7vH0X//
KqkcETNVAmAWy2GrUF07/H5KwiVFrMoPwzSJdvpnnomO03uIUFmmKyMmZD5KTkzC
kmQpM0hTHrEXcnxNnKlKQbAQ/7ARawdN0JHdXGnAcKywO4Fi1+4yeT/2zE09/t21
DxwJVYzPJf8IpPLqQg7hwDTHFHX1Xe+GqA6eDz9HMw7HtjEyj6UsXlxoXNIfwHdY
VwKcAfz0AI9Zk7ExVZJKMB/+9ETb7EC6fZrEolhQ7zL/I2bGN420TwHjlx9t1QxS
dGkK/kSHcNdeYlGQwJ5nuY4dVSsWHS9PycspKSl9MhXDI9LqMQXEwlNJzSo9YIWm
YRRxq8ykhSZFPRzbLi1shW4sg8opaVN6v8gTUDmgKLY02xr/S26D01dOpP0EXvMr
EEWBSDNK97ScCrfPykcH5oCRhSnlOKGZa6x1c2Benn+cHv7iXFwTikhWJy/8Y6W/
VTuZwSv7WHGsZpbW60J7aiqLoxSm8K0KmuIz2kxCdGaQJBJFvum3oMwxszYLNE74
PIqVIDXDyquTR7iXNKUv/NuZfvtWf0y9bgafYX9kSCjj8HhiX8amrbYFqgBcDTKS
feAikb4QYcHTPc5n6FKG+hGP9a6oW86ZjJB1Xqo2BLSXaMlBboh2EqYwHkN+ZM3F
ERGYyS7jWHaBvYfhwe2+Gfoss8fSiHq94oxQk+YZfDZUqxJR02Ho4W5QANBFh+0I
Rvn7l7XLkbxKlteKXI0z4ZmRhtedkhWhJd2krUhF1idtWBYVfvRmZ4310vTB7/Eu
TkMOwdI46u8GBdI5tjimpgaGaVgt0dg4uN+Vt+ZajU/pWOgyPxdRDRWVHJwbR6hh
mTbS1xHrN86mJCTbHf1TFG6LcDQjmGoeCSnmGsXZ9PUyvK5rEcjNWOdJ3ILvRGD0
HdyHhYN8Ysdu4pikLwD7O8WYyXAf8UuRki0+GZV6ON9LKftZuRmSGZc4TF1Sb1/j
w5XmbUdQ0fILQlH5sfJQ6pV9NbOMwpszFH5B0YExbxlLoF1AqrCQ4jlKqGJiAvpL
Q/xI/bCBcShEQ20GKFaaNOVe6eZIJ2SL2MJ3ywtMlROMzhoUb8RLIvbVtpKnyLQ6
Vp/ryw9BC2TPavLewibiuQzNzKg6Xj2A70/hdRgTzo34IUCCenyirCjPN6yfVpS/
luQV2LpXwAwSimJzt18MPMVY3hsKpIViY3ASAbr88OQo/61oZ3domt2bYFyddRPN
bs1EXbOgOkWyTbovsc/S34555AC+UQ8xzPG6z9g3I0Jy7JZtmKPi3FifKhcgqh7U
3VLRFnvmJ8QI1PZXeTso90/PyXgY8N++OwG+KuJ2xQPu9JPi5mWE2yWE37dD7YKJ
fr7NmPXfGtl2K7HUYKPMymgJgLJnmDo9qx3E1wptE37RWNW/WgNeRw3JimSV8/n4
oAMqGyTTAmHGzlEW/G2herR+nuY1W9tCVm1vSJQQ1ggWaxLbg5lwtBO8mJEcKV9e
pG6bwibkWsPn9EwwWnp9gZxCBfO22GFsCaHV5MxH7IlKlx6lvkoJyTWpyoP0/7lN
JkTXSAkqiCsy3TV2PnStsu89ti80ttPSC4Fwi4z75AmRm0eLb9viqFk+QgjGLSbM
5mx8fEnwQRJhNscR9ZgWAnxXS2a2gueTj5o3MFKEhNWNoH2d0aviNy9mpBEGfJgL
ScGSIO3aBoLbq8ZMCSHNFc/oPEImEpee3U41H314FxXJ3ptB72DRKIF3npUIxArN
x97EEqIrkEjbqAf9tLl/3+aNvCeadih6lx0hxH1wqgkp6XYxaaN9dettXoVJbhBD
4uha4Um/dIQpqejCyksE+7lCUkEV427Lsd9p7S0bCzQ7EoWEMifSWTGc8nBMaXM5
ofAs54nSJViBXWKzE7dN33y8hN+4n9IaTE7Vkckf6NVhxDe/FDV9wgej83bVaXm6
MM0qsZjOB29TVvi0/T74wKpGqlyVJIfNFWZhHjlSYrNlHewxl+SplpFmyicRg+3b
uQQBgTMBtCygYz2nHnyma1qhUiCNL8uwlZkxd01t0TNikySWAQGFEzdEXHg57EqD
hfELbI/Jf6nJpJTMjS/oLg5pEGjj76KslG7ieYtxfXdOMsqRA4O+uiY3AyUz7EXv
DJVoK/BUtrQaB1gAEtxfsq1vR6lKraWacp2YDpBWhYVTzjLcCKoT3LYhuAfylc17
btBdthSzyd5TH2QXkKHwHlm1y+AP2VvS2iWvU0z9+iy1/9M+qYiRivfL12o6cqIP
OIMAJCT1E9AxVGVOpxtFJ0Ccpna9ZauTGR2CYhNo5ScdkhftwnmPqQOd63wXD63X
TG/Da42ODmNduHhmPjnblMvqoN4ghdjCgth4+mlx5QVua+J0FtiWO5amYhMgbTFr
cUgC+RryAzaa7s8hlrkYq31Jg/gomdwJj9RdG5cPl6Cb8d75WsPTy2IxBTqf6hhm
DCO9vYraOVkNnt7jK4qmfRMswByb994RW5hU+wEHby+SYPnk88TOEVCsp6nlH0KM
4X6tLanRi5TTMXjbhx1fVMM3+UAxEOoisYCgw7hWiobD5jx5nu4NQpqIzmkcFg49
KhOFJXGMmQhWHQm3VA3KNufrn4TWeGxHhgWZy7Vuqn7ESi16QPFv/DXEzqjMkvnx
cQ0VxWhlsRjXReeVcRJZkGncysXg+jlulnx6XclOPXxSUwHYlOmKo0x8iycyOZ/4
ZpEDLpqFBDRWsR89NQWEuDdGPLYik89Bc7qdp5fnYmx5etNqv1kPtsp03aD89fVc
x09XveCBXyk1u8XHVAJlAdsZGn/FfjqpLKJ0gWhxA7cjJBfNBZJCFyXivtJAW1sz
9GeR9uKn9LqRs8KxZWnNzu+rfWi4L1AtUnSWGixTw/Dp3SCB/uD+x8Vrqf7OsjCv
u7x6mUCGWDBfGSpeiMfZt44fziq97PQA2FskZdhe9pkLEG+k7Gs+bKgotAmSCrXR
t+rGBT1hWd5Ld3fhEghOjiBPSPJt2nkhkm1+G3SMvXWpUvznfz1nlawP9cXDX5C7
WDixf/WBXR+i0keD2myq4DEg5zz3DJZk9IcqdspkwG+JrelxfTFhW7qWeNxgqyxs
lLPtDvldI2hxqu0UiKuXgk7dLIut3EJAXwtGg//HXQx/yMUN9KwXr44w3I6CsEFH
Upc9FM243xe9ghJF1vEfuag9r7sP5IYBI3hjvjiGvBhXWhkldtsoBHZi2qgNj3Nf
Y6n2rBM0rxUKAnKRcjhCNJcVKhJlWgH61iDZ2dIZipt4S5A/Q8tnxtVrxdArIdYz
/VKz/CgTsCCaAPoKKbw7aF8o4ZawxD9Y7E57JHsNwpCL43Bg0TwFhXdwtJYxAITi
hEjpHUXqLbr9vPbKwfsXir1NJxx9hzSReszd5dW7MbLN4f6krvxnZNRG4xpReoHE
ud03KLh+U7v3mgyZ7YzUGOoldq1jzvSQsxauVjv1RpdNM6XTLjsvJapNzW0l9qnu
mOAQD8ylFEVYFUSiG0wNeu3SkZgcszFuKTHJ8IRpg1ZoknnEnB2yP8KAcKGFzAbU
YYcEZ+W2xbi2PVa2E3zKaOemNAWxlRGaizWXwaPcoX1HuzghII2/+Lx4l8O1JBvq
FFdXGD539h/MvrTaXfW66Mn10CgERo/Z2JYx+8SvjGwWBiZrpYY2JN4OGaQAjgp4
Bqy6oeN26fyohH5h1Ps/HOEJBLzBpE5sUiXk8OYKAIsjmQR2/KNxfvd2AEvOw98U
vsXNapdsQaQQ4cTuBbKDcbX/KxwMCDPqmSvdyGCY1IqCK8HGWGm5wB67EamaCEgU
WySdh5yy22v8JTctrDVQdttOpzCRn0ZfIZIO8Lht1dNo55q6LhJ5LlCjZIXxWQPb
aHDH5sDTPt9yc4tH2yHao1TdjoSmicLfRrFHLDU1iMASZxqcYqdWrLcx2KqwTLgf
xAwo+htV8IzckHiQyKCxNgNNmaDlied7eBftAtmj9YJ1WrJKL2gaqe64aTE1wuGe
a7VP3odLm5Efdu1ieBrWZyfKeqHFVBEfrJAnu2ztL6ioAo25HE+1jb+4vxFzOli+
7+WeUvgfpkfdIdRAQZgPvwEvKJJEj/O//F7r2A31AD6BpwJVSbkV3LR9r2llpMcZ
AiLiIbX1cnuGo+YZf3n7wbNE6A8WX4qlNmAuzpj5gbnF3aBOYcttPrGC94QxsTwI
kJUnHdWgfSYxswd4SHZB4tmhcK936/ORqLotsAlQztF0UXQ7O3woL5LtIfUf+Phl
KnqXOd1kzCbeUb648PmmumDnxAwgD3RBTYZ7wyI9mpAoWcJ8fz1ukOjkA1hQdfU3
cQw7WwHXnueNtjmxudy8pd4CAKAFnOM3qgrwV9WIOzeAOctYuhriHaAmy4IaWo1z
spbWto5g2JqvpMWz6r/8LoUKK+5npihW8woEZQzx1tlyScu/Xi49qsvob6RnhiZi
g7iyvNsV7b0QMSAkyPEcoNm6EV/lWa5mcldGmI/jbbKQCkrer+w7GfKxrXFiwfbJ
fEK1zpnLfy795uj1ShSc03mOHQSH5O0gktrIFgzyPj7i02bdjctK9lPX2sHGDtFx
iIWAKoGdQQ1JqUASkG8rKFbjUZo/jIrKivkgdNWzk+ckoCHu3OqZrT9lpn517LKI
MZ5EK3QWoF91FRv20cMh/Qlh0OfxDTl+ND7PXxFvpP0Xc4kYBKPY+mI+ODes62Df
lyupb2Bbg9YR9nD4WV4WZucpD2UYtBiGcDIV3s0aIAHhdjImLmbj7r3zAyW3u7Ve
VWwj2z08+Tia6iQW38CkJswM3z8C4GAfS3V3tSyUfSPS3ZiRYwTsyHkGVeNW+cFZ
LDo2+NRJ7Ab/k7mlTN3J4NRzwetyL6tjlE0cd5kd0c6tqupX+jGsPo6/tHhY43AO
JrQu5YtvAMF4Rsnc66BB0ddPTGfCB3e4LIW4R2DxUz6vAqrmgpZ92Xa8GFG6vC+H
OecP+1Zn2p81L4dR/196v20xiYyyYX4LHwv1sxzaPs2MJlmk58u4Ni0YfDLT+DcW
h+Ro0PdO2iuGsmnjG5qSKo695onkvzbAvYgJxoBPueGia4nBVI5RohAOIZhhuZDJ
E4EboQ5X9ItgeZ8g6vSaR4N9aEiR0bpLUwv9KtsaV8qusnnDbeU8KXHSUWsBqoRN
sWYVZt6T6z0z3uKcEtmoYu43OtGpdykCYWMUrOJ9kvJmusM1CPT4m0IMR6KoAwwu
qC8ajhf7kofg1t6iLDwBb7Lg1gWtO5qn4NN8e+F+ECQ7ZHRzNC1+xmE0RKdqxKh7
9VD3X8UFQGPHoLbNTViu9S0TKkuqebjp94fxE4ohMTFE0brdwOj5+f47LkDf/NNF
tdFpY3QHphQrhGC6uiEvWt4s2ZWP4Y0/rqxCydzT24cJDizhXPW/ZE1NH7ce7onG
xNehZMoKD5SWOC6zDpPg31lJe94C8Bno4mSCFLXlqphHx0gFoCFLqQ/23/pWcaBB
kaToaEPLPUARwVRyZzxuthagG6f6+c5KzM65K+2DGDMEfaGaoIIdNB704yWnQnN3
+jdU+Ap5ouZ0YoEPfUW8LDzOlLx7LGY3V38/QD524yEfSr440370WdnH0UtIlAEa
ZiUxdhg0/GJ9tjd4G2A6L4Sm/syL+qXnYWor/SnU9g5XBL8lE35O0T3BZd10b7t5
vGovGM9m5xIfcBqSnZfJyJx7IrinH2bUoENiXvR+jJ2ImoBqEK32Nc2Rd9UfHIEL
PcYOOZOWjnJWktXYAWwUhFYV/LlLtn64P0gabzA+m4whoOtrih5bFfDTADhzmfQr
8STpHWwsyjqAcdS3xJVnlbgKZC8K0gmRWOVY6g4DSo1Wz/K1DJyMiP3deHNL4PRw
+G6KNYcsjIYpl0BO9pWkLkRGEExb8hcK4KbKwd+SSH8Jjktan3jQLC06CXA9GCgw
S7iW4v0Y/FnerwHT/o1DOtFKP0RgSsC+OYBhIiPkZ+aqqwLZzrvsWBCA9ZL50a2U
UWm3JGqntxc/1M8fHlILM5j2s/vT4y3eod/9TQs+pA7Z1SAjl1s8WiLU1YT8A2Qk
A6kME7nKJPhd2lpEiPuzGDXFut2P7xQvAS70M/0R1oCfPnvSya0G9rGla5KdvPZO
PMl9RSgRG+k7hyizGlwKDRPxrBwkKXkQP7I5/tsX3ORCjtiF0QhFdNXwFyR8bcEP
Z4vLohNgksFf11sYXLfVjPwG276XeGELxV44XsdwF7Tto3r3vpHGlcQdPcm3hIlF
s2N1YkYmaIEgV+zVtVAvkfP0tvNocrMuMV5FiGy07XqtKP88UTaNplpgWpBInpol
MGZWoHxPc9s/ge0zN7wajUad6kCKoDRgVvc2FBnMHImKNxAysEv0kwhXwdTVAkrN
L5v9U3b+p9cVnPM24b1my/kUkF9RjPTWhupQb8a1t62/tSEsoevPV8StTMWPMzOp
bKAE8PRFvPubKTbUJ17Ga9X2EBmi2ocF+HAezi3H/lmHPbxfzb3lAxJXguHKUajN
3VjXoYp6qb9oBvqtniIXi8jbtEv7IbIXKG5OVpBm2Xtnd9oz+ftf9QErcssI/3kR
c2fiV2kyD/t9nKUUIZd6pDm9azNNzydU2CU0znJBRR8ETUILIVGmSzb8h29KIIi+
V6zqj7LCiAM/Ep3L+QNypVCVuINbaAJ9eiOTcYl1/hg90eCGaDzU0VHjVsrWZLnI
J0sR9gPLak2ggIuCulHTgNjjR5ilcjzrUL/pMnZtz2gK/JQZKzyMeJlrnaUseWY2
8Lxt8QXw1mdrRYbuB0HeNrZhATEbO8zs8s1q/I2hBF9q2pR0K2PiEtjtmDeuusqs
+21FMnZAdqZ9x1TDqI6GHLz1EsbTQpvMyoTx9VvAXsTbrhpAepyHPeY/Xz0pV96t
1dCz2q3uK/gBw2puPngLVhKhbbdRUCayJIwDH4xQqPK0B63mJjWexTd/xNy1paR9
EBl9CWIP8kFp6BDUMpzZskUSILvXs1n573DCOUR/plWLBtlP7GXBLw0nbatYlDg6
F/TAU1Ha3UqWIvJzu8DeMpClf0QErxIIpJanD29eZmwOzf3q6PrsTXJsqT7dA/p9
PmaSaTukJgq59/olkKDhQgvcEXIqEQGKswVmfz7Otl17dlyM2NBVj9KaFvzTuFdD
x5mhVe4HZJMD5qgBHNrYEYttsn94wUz/qt/V0aCqEWMWuB+U532slZ/cWAJdIkwU
UJW7Vj03xZmzzBjZqHnf4DhJIyItLk9mQmVpu5GntowbRm9xtTEmZHhcF9FpAmFM
Fu38tldlfhd4ssRgsXaVBSIUfLvbu26sH53H+WIa0RhkL58U4+0AUgYMkWoSiwy+
cVUK0XDVmPvRBVWryZcRGJd8h/AW5SDvy+dJznLolFB0nOZrNf2xm0AjOsOuUM1Z
d6/jFms9e38q7jR4oA2Jp5IQeivPe8/nnBIzd9Iz1XALelFDg5Z53dM1cJ2zbgJe
zozc3fHUv+FT4bEEyS7U7VrchekXmg3y54IBpvtwAFgeuaOHlzIUkNr9w1I0UUO3
xchGoiVP8QdwPWzCxu1u7hgnAxOd4p1KE7QqM9n09NGBVZXOHGD4wlzUT1tSZwOv
wcGjhBmQA+S/igu1/EJMGZqMW9lc+QKmCjklQ9PiMZzeDczAUSXJC7NrixN9i4Sc
sbbJOnIp0yEg9TgHlv6Gu9dyKhgruZcwZXpb2TuAOkUS2MUNdIP+wclR4Qhb3Du/
3gajcXb6pYMnQcMmAGoXDXeqLIL/7VTNmREs+p/v66eeX7x/ptkaYy8z9BjT/GQS
UybsRGy99QtaQMGfyGOr+EuSxOX3Wa6Jzz7cZzhNn87qA8rRyZy3wD4w5jea0d/z
AdjG9ijf1TOpmTkTxKT2TcCZtxcMPiXc4s34mWOQPmFI8FktzJuLp5h/zh6mR08y
dd4Etl5RNaSSKCgNbMQVJ5Jh6GDrDTNUNqql8T/9i7LN++Mg1SQs4ocCFrZCtZtt
r6RlrBWxuMD1BVfhHA2i/QctrXdPNUVvBxbciAQVbLFiEKtJSsMfHHaqFS5QbQmk
GFaXV4dCGSTuQeFXdIe1gcj/EvX2iWRQsehk3a7E+1POiTtNqclhAtQ02sPDLGtY
ptH7MBxQszCnkxn9CIaDaZ1rhqSUUMLZlaDLrzbDFupDA4NmlWpfm5pOeK6YA0xl
1Md4Qkp+ZvLna2vGvtv23e7CABZa3bS+3abRzxPjxKmKfjb0H1HrWW002aYb9g1K
B/EIn/V4IKooWse/99uLMMbkAKoNnaIe3Z64+naxpIXQJp4XO7/Ekfqtv176UOI1
LILgPV+2MeAqVRTViWThZQqGfBtfWbub6/a0bdqdiGavkoaB7m29ziJtsXz5wVE+
GCnkKX+BsAEd5w9M0+7ttCADPkKjRHRDFyCHb3MxE02xoLO+X0JYL5phOiGJWRqh
hfLgv7pdqAaCYvrCjVXCGTSvznQjmRx2CrDvRQC+ZyY1MbpVRhRjyWI8y8/vpY81
br7x1W2fJPY+sXUAxuON/5e3UFNb1wIyDXtZBb700hs4RpGuO8dm+WfZ0i+bEOH/
Kt22agSml646H4RqqlaFMss5WX92cMQmon8LcOLY85glkmErV2+B0UgPTf1qZ/Wj
nTl6Yy/oIHAHg22H8IZjeAFvI85QhC2U40eTy4hCupfoD0wyT3RvSq6o16fHjofP
ZMERtD7acJVNeHoy+ZUuVxyUTuwAXHDJBa1TGA+zYoH6cGmD1xpsv3uszlF573Ek
YoRzqy5NzA24gDnk/KbPv59c8kLUzpWrmHRkFmU7ZD6xviInXdeo0EaN9Gowikxg
cmesUTRAWsmJK6dlkyMFDhkbiJoDx1f+h4QmZfiEXw3NUX8UhNYAG9XfHAIeyLzG
MmU8QjWk9/hOVGWNP46eBKzmbc0fl25Dj7y3ksxasKIHPz80wk8Pe/k6xv1XVcp5
Jw2uTmskEwmWMuyt0WjM6cEYDCN9+egmqPYyv6as6fWu3tIkPi4qH96o3pKghk53
ps0mhI/CicTt59Abwl8y/DhlW0T7p0anEcaDF/JPK9VJptMUrD5QL3XNyaMqxtaK
7TIX6F5CaPqMgswn8ZX3pcqx4PrnAtUFIiHUD2//nt/GbyzPAvr9SDyKMbRdw1en
3qnlPtc4cds08GJOJU+QY7+BnDb9PaxLaMI68o3/BI6JsX+vA8CdZcSsxL8hy8Dm
wPfLA3B9MyKk8pSIASGgi6H03FIZ1bcWuheOknSaeMaC2WBzcf6BtUD3zNDjPiEt
ncdn4Up15NR85UCSS0tXe541tTADoxVZdfx29r7rpjtZ+QEDsj8hJCIGec6x9jEI
et4zDmCRRU4EhQ2NojiA6goxciopiuIEgbiYUGs2J28jyuEXzwWyFv0djZMOFR6V
hb9YWMkZr/hYhDg1PXX9t7Ac2ZAIndYV1rFxIgna4Uolquj6o0LWkKxfSlxO51Y0
bTu30my+fdXDLwBXHUFqQVNCEPY0goryPmb65BBLtwIp/BakalQIcdIrFlr/wn4q
3AER1A4Zpf7o3mwKJwnChk8sfpTKEBsMen92wtvQtRYvZ2HUdjmt30dZy+jnUzXR
Nv3xT+CsVlWMBnqpxmiPfRy+AR5Fp3nHaTIud3rsthiGLWol5nrzaiJvy2YeLxS+
rp8xba5aGKBHa3Q58xS3cIgjGqJu5ybZiIfF8LRW59de3ASijNqzfLR8nOQQtqHx
SgTEkCRllc4ZLmd3MOKTZKozONjly9KbIrRqh2TLcUbMHk2yuDfF7/Avkj+Nb/qH
/OFsj9XeLApw9MH4R2g9CgGv5tzzTWu0TdsGUgN80xN+OTF9HoXm14XxzIFyNzV7
7SbUtdGvJa2lCIsWl+9qWvURHNmB2M+5qikTIQOT9cvnPHpcbCmPSGDk6ive3/uF
9MHZl9nPKwhRtbxw/TeJDv++zAKWusDgGTWgmn/kLLl7gJLY0e6HEY8+q37kQTTK
Fj3/11WmRLWU8CtGCjxm2jlzij29Sh7b4fcPqJBCvBSHXJKyGg15jtElRFwoGP1I
QlPtWkps2euCeTi9IYJH2bvR29rEeQvfALq+zCx46hS/Lpu3j1W9T9VKV6n7OgSx
6hPm1DyEaUzTV+AbVNznB7mzcJTQsQlLVcAly9JBiv/DRDNSYLOpEORrGZrCLDeM
ixml38f2yOsfUhK6v6hRnNe539FtsSCGikV9mtZRkMQJr6U4T7pgiO/oppWleM0e
/tMbhkUJSGbwmpWMGNVgwmqGSTE3am6x/tAZalajzpIgPUxGUE4lEPOQsd2jjLFO
MmZo0a6CKnCP2zPZwnkv1eft0b5dQshb6c1dJl9oWMyK1S8DP/IOBj6i7GQIvRjN
3KmXbscnawPQW1YEsqUrgUUTJdwk0h2nfqUi88l9dVLuzX3Bp3sWPwIu8QWtN4Gw
IL4pAZ8rzX9pCEruBslHkhT+tH8L7ZxnujCq6KhUHIzt6N+Ok1rNdG/P0j73ZFMq
ArVpqM/ZhVwzp6bUacpdJ7IPwY/CtXAvwtGw2c8Lv05vehHlCQ+QtX1lFGBpRrrg
JPvtIOvZhpKzneAXrHXknKYCP+Y96NT6P0jPKE9jDMKcq+msfN84/VaKqRmgabt4
cmazp+cWqUQyk0KcuV5GRSHhzqIxNo1KJCOiVEkhibWSyxdFZxvDK4/p5xbXo1n0
PTV7Y5IupYR8IkFUV8oTJAJRvtZVjFCwz+wzUofp5Zunk3mT8WfUAJ1TL+8dFLO/
/sIDfx+q9djSLVyqMvZLJcrI11egwp8A/VoXoDEwktwULw8pvV+8jgjcsTYL10KB
ETFHhjHj6+5Z1tpvUsMkXQ3yAcAA038NUXVPWsuXcHVzgRpEMSwkY0dqUh5yE18X
ujoB0wUF+0zKzET0ogo6P2xrQhKbed+KKf7a88g2zn7SuX1Us+Jlw70f4PSLVyh2
tQnRDZ4cl19MIbWLMeEFpRjSmY8noEQpTMpDRSNyeLbTg5kiUmm7MngCKzkHoCaV
g21x9yUfv7lLr8NGRGUKnQKzIxyEyF3J6elKBvaPKPLFbEsj+6/73WvLg/ah5DTH
9T/KdP1lSxPSTHAZyqSah9EBvrU3rVyIBYvXqNSTWtHHRENWXeFySM0fO6qdbTuJ
MtL4IibDWxUP/jklyEt6jzdYesUhkyNOiilBHKl1PjyFEGPTGeajAEXAaolRR0k3
Iner4qtZcFxourJ0Vb1G/x7bqwmMB1YFW2JY6kh4zeMMWFAicW4gMRcYcz8AQk3s
Bz+UVmPZRNvhl6VFZ4ZWKO1+/Clxn8cY6ZGxFEKderurbRLxqanjJy1vGYUBHGc3
jgUEwuVuAqWA+4x+uhLnbodvZv59PvOFmkdGiruRJ9nWDiEForHO0haK/RenHeX+
Ye8p82V20bS+jC1ghZFdPFcpOyusf7AGdezHGIZ7qeYAdrmAQKpKJnw/DojG4EED
UCbXE03o2bqHHHXAlxQERcyY3I5wBpVWsxMrsHncVD6TxjsDkrdon2ZBB1LZNB/5
3E9H2mvDjW0rQjO0cteD4OmaxIY/vK/mDFdC2aBKafb1t/G3ISeo8yiBhTjNuzNU
I3lyaLA+FB+LelKX/o8VMqJ4H7IwS8PxXI3FpVbwnhURMlhPstIWQZ+f3Wz7O9pJ
HiTzVK7uNz2jjF0F+iMPPpTfui89ES5iun64B662Yeq7K9XelV2+bPJxjYhmST9E
8jgVYQTwlziheEhZK6ghH4AD6yCzLgW+eaM9ePZGKy6L2Nl+Opjh6mnnweo1bngb
/50tb8HKxm1y0V0/iTwPSG7vmJ5oJ5FMskglRO68v0xrwTAl/Gz2oOn/f18AndIf
Y3KlTZ1rJx+YxO1CNqktgSenBMXbbZvnPXWrRGt74XP+ZAz4N/nq5GWovOnDuqVF
43acnIMXwGHeDv0Uvj/gM0g3d7vUh3C2rwadP+0Mq7ypQ9UBsDbKc/u8pXH6vURc
bjTPltoCgpJC8sLeuZlmvaNxCbd4En/ctsjmKfPmKUX3gyDQc25x+HNssIp6LvSc
WF7kzjlCE9DghHK8el8o7kdsM3upUN9xHf+BM7/OFxNAfzEO/b3LPYi2MVmy0cUq
fD7TUZGzfJo1wo6p8Z7dvCtUcji731U2jt5S0a3Zz4KlsEYGPqRA3RzgSmdWHyOS
XwUs1E+x7iSubcigzLSzoZsJri43y+osSdJ2Gu8qjQboxkHREMHMf2d8OmzBPxI6
LN2kuEsZi3kdNXAn8nxUdbKb94tdp0qjH3kgJs1A9M5i3sOJqhDnAksPCsgIo2pw
3co0p2bFrOyU8y0CS28kQsagcu8W9NOBe0OHNCRATKH68QeES3vHgYZn5rLgNf+Y
hIZ67h8BxuyFfX6Nsn4Wp1U74gmc/Xq9+rtUQPeLVfntK/MgLnJ3ewRidFaRVj9I
4LN2BdHNIRZIYJyqW6UEWg61EywkSzTrPTJk9JDM/DyoWlcFcVPac4huxC/PSaxD
s2eq6sUnz1QR0X+5Kvsx6VDl5Ni7sCn6yrIDzHXLC1vA9hU59E9x5p73zBPXXlBP
iFyYvlLhu0JgsFK9zOghX6V8XLssQwO3Bg2a5PCX5Wxt4ivjq3dmhSdJK0Z2l3z0
MpPbbBtZ0qhTEFOTe0FzNf03wVF2VKU/0Jw0d6hd9JJLaDrxTKfOZoSlhDFfbnf4
67ssi92A+tP8Xa2TQcLFicrQv/9W+OmU+GuIPnbXgoY9+TKI9KUCzUOC5Szr+bCh
t2UFtnDB8mTE8eCt/+C7iWHEGEmIHQjOSqEy1XVu687CSV22yezxCy32IgTlWb3Q
tGh/aOYE4YtomfV7f8jDUURtwfWDNCUzjGNhOV00ZTEm2LBATPN1aR5vnn3RHSRw
6qNJDVKRpSwZmRmWk3X+KP12Pd4EkO5M4VNB7QjnTEcgr2bgxxw/n/QPZlyORc/Y
csPIZMvAe2Htkt9CkGABgtMKux6d1bg3+tTOqgXijldPfCQr7Y5GOTGO9zKB3Hzf
xnS2FTX+QxnkXGPf+p+S3PMMV7Dgdj6IY3WK8IXXpX4yBwhrxLwl8JJiVguyjYrc
9paL8spqT5saeI/q7SuoDLZyShW3+K54FXjD4pJPV0NVAiGulc8rt0Zk6sLjiuh8
/lENdJF+o8Ajj3t+NoYESB9ogsK9wKxaOa/Ne3WLEcKqih9WMBka4vJIZdNv1Fkr
65qC8XJTZJskKw8nlchYTxyWmtruaEKuIlmooRjNIu61ikV07VzagHPacP71IH73
e20SSHr3fwwBmf7OvvGD5jNtr08EQG8AxgA3PXQ3SMJIfeFOm6Castg9XhIA3Ici
cGlJWBbagB69zvNrQGg5+FHnxeBjqp1+mfSq3qca0HqKC7Yv5TdBU775xtqZywt0
QJMVjQ9eHCotL9jEYgsbwZ/rmOBQOWviJIAAOTNtEJG6I/lbnMddxsQD7M+uiFWn
fI7PEJMizuFbnXzJjUU4bFD46f1yUDk6KX+gt4gr6dlIMSGQIgEoTbaGnfoWq7in
eKG3rxABEOZ1N2G5f0BbJmcs1iEXSPU3qb5qmjlOBUaxVHzup0YloySkrp2t+qdb
7h7m2K4XRAOqQ9eFIp3Gn7QZriFM3US1AyRD4JzrtgbrtHj+8/nJ1HcpF5OmdPOb
aWkWKC9p4Wd6fQtg6zdAIfwAWP0i7YwrQJZk3F0MyX/qOtm/gnCSGf/Xn6TU6ND7
kTZ7AgWQwKsgBqQvagr8N+acM9JJeqQ7uJJ5VuQhWf1XYGozsjJH2b8fNZVnpO4F
DsA4EXS5Ngc/SpNph2dRWGjYovBdyN8QGnn9yx6yt0E7HiZqKgoOA4sxDoigi0G5
pEAHcXrs3dtPh7sJxD8TcYHEz2IfFldvB5zvOoh/ugGfhBAb6qLuFdZYP0213CQv
0nP1vh4QW6p1Kn0UOLj9hW5pnJyvK9V09u4Tkt7KFkPVqLQgkip+HxjZg1Q4ypUZ
Z28kpXtNsVzaZ4N+ycqwjSpweJ9zCSBA1YTQ7c0s2i4bK0D03IlFsp7j37BJNqiz
cKRbCpi9+uxMm/7x0ATEVqYgnZZBEGk9z2X36wfK9TRadI5wb5pdoWAv05lRW2GO
PdI5YcD1sb1AXj6fYM+lPwNoFvYiY26gZVp/uIEUTa0srC79cUk3ho4yF50Rqur4
/FpmrcMM5MeOubO3YjrMd6yqhY2hDo5QsmhZmEA9OpwodQLIhIi4v5qNWjBFGIgV
qDKuAWzYXUJDkKInNd+NFn76RCD2+20W7qnlZax+BYttd/sJXsJFIUbARwuCbCJG
A69VlSSaS7YSg2tKJiV4SlPdro57G2zavcsjlOqjsiV9lWIzsba+3zxtgy9HQkW+
GUhDimgV6JFtjBmBt7KCZnKIxVah97nTxb3nB9RGJRYu6qFotZ9Uwn3i01WfuCAU
9Y/BwNM/WFzUqlJraZs46AiNsBV+Cvw6fVJQC8YQgl2CgKNHuayMw+pWWsJoW9yy
W5cHaiFHq7IHpTnN8KIo3cLmlekXMyv8mqIsFesKuWqGqC6zNeIyt+ZT4NZv3+/m
f6SMI8lTs0xW3zKfLCrgUpYDdckbA07B01NWKyyXbHqmp9yfniKsyHnl7Qc+P6Fy
A9+KzUowhDRg1YEz1OyOuAZ4mZnG8IJbyGRiGRMjxVQdQ+eBuNx4OEx4OhLF1pRm
ZGhFYy03OgWFhBZ6MJwxAWM88+wiCPmgRRF4slDJj72xHx6p5Wk8kSXQa3i6sz1Z
KBHaVAYF9n33nty7Lg21bBYnyHvGeRUPPqQmO2yk9fTOEuRGb7Yx0ze5+4stTzF3
NfRuBx6cMB39A2lmTehA/mXwU25qQjZ4N5ZLjgAWffD3SPm/ODnW5cWgXyCY0G4i
y+y+wXsUxClj8jT9Pwg+ioW36YO9X09Kj61rWYc3NZmbLbw+rjCIYv9pJtiVqjAJ
hX8akg24GdeZodsUPafgQjoGlYzAdfM/iNAjBejQ01yjT+YMlD3YX3S2J40sMPBR
y7LZHnIvC7k6e63rCTcCFPXfQ5sDslzUJKm2O6a6bjloTcHq+raMG2RmnOql5PQT
4snYP5p09WkBSXl4IoqBGSg9qaKCqnkJ6bUpQaGjqGRx+gtwxD6U1FbkEsNx/Tgc
lAg+NWl3TSZDpWGZ2PNaAEs+hq/sTld0K8/+WPsErabMmBVBeHABsejvN7rhJZD9
Tcb+r1OC7ROoA0DpaWCg48LHJ21SqSlP6wHlKAfv5sg6U4MU0gsQeytkBgUAvz6b
KE/l0q33kUdUU1KEeDC/y8EyOX14788cYlHiCGT699P76uNKY7MNwD5dyHot9vY6
roTlQI3Da4rjarKd9oWNNmrr7ArsxlobG7s0cPKXx0ytOComyaa+uJpahLlO1h7J
1olYXiVZfIQ7P6rjNUhz9hGmjdKv96CpUSoU2hNdPx/scYpZgyrGZEjIcOVRr259
zjKejkmPFFnMugHNb3uwbT+9Wfh+9KAK0DwmiFojIMHOc1FLfTKVkKMhRt/Z4cWK
mpJjVnn2nNHE6vE0E1QYAoCcuRL0ROcX0tCXAJ45coVj4BROemBBVN9neOTojPIw
mRI1gOki3uGEYIb9v6Xvm0GlT9sp9MMkSYW5fhq3f9c4BmDpeZ63BPV379qt1qsG
GmjcxOlfl+97aKIQRfFs1P9/VOL/ETRa2FwE7gJ8RwTwTwXcOkncEGvWec15tN2C
pCs1qyKk6o/6kMHHHhKnmTPwxgVZDTtNaVMRJFfOExrJHp2CokV1TlXgGYLr4Sjg
cO6pK0uKOJse2qDq5MfMf7maSHQy+f18jT7IAufu8WkEzd/1l2ajEXcqspZlyjCG
NAo1VTE9JXFwIM8cWMpfQNHeHbdhFBtGxG+SbV7wTdTm0x8gRz7kS+I1WxK0Xmb1
Td03qQ10+wP4A70Ml0E4B6ek7Lu/5d/QJm1ASHEK6E+5eUBb1MNsrNWc0BvbGp6L
fVWG+Hdnoi/ZcuWrXPRVmImcRzWy1/Ls5OhTF21mj+mNt++8KiKxEmmchakgClVO
ePbwH5PHrLIBU1VPXxO71YLVREnrcfBnr03q6b8vx0BpJVjzVbqdvWeGqhdZ1gCX
oUszLj7EADjAKI2k0cN7356Oh2MitITEZJ0r4pRUTfkCAcgY+Z85HVr6UTkZ0IRP
3QgBOiKP+RtfhaNumeulKnPD6b0ySLOyV2FCv40pN7WalFpP6mP2TYf7TcGdoaYM
i/ofpR5G9irK1wd9SJEgiH9gruCfLESX+7MMi5RGp6A3xItDZjKi1L/ubLKVNf73
PwNL4DZn7XfkcrwpASKnkLG9eH1zSs5TcT2aSY63qUdG3VGpDhI7kEvIzTcAlwxl
VDMoSb7D9kGRM5nftFq1G/xR4tjUcRFJkfiWYpDY8qh+P9nvhwwZH8ySVsRA3ClD
yQnq1hfgBdSRm5NQxz6HTQ3peO8EtJONuJKPdl45mZPBwdR2Wc2Nm4wepgoUPZhR
5IHzUsBC3AumnPn72XYjB9u10nHwtewGPyMTv3+H1VhN4Z0sMecAl+C0P9VC6iOa
t2UaJ9hUfQrOfLinxjoWcvTjVy78J6m8GoLYRiG0G8HGqH+CMAmkdPtFt4007CL8
IWzoeBRETBaFXb9CQClSdUirBT3Djn8aJXgGsNdagn7KbBnwsgVhGhFwYnB0mxsa
GCRvhyYnXQgo9jRhwABoVewOoyDCbwkZwjE3P+WZPLCNRB/aC9iGmMBDUhnlhaZK
ombLZ7YVW0HE4Hun04ZOLzBBtHtKKGOr/56pa1txiSOm2kFHYLR8n/2pMZRuNSI4
io7nVJh0Nl7GedsUJi4GTtmfTzeERhemugVhNHmlISA1HZpwqYGP/2M7OgUCA8E5
Oz4KYYgEgSbnRG9kLb8TZtH3uZM/qYS9DWawi/jIohAy3LEF+29TJ5j0fH5/GOPi
iPARdpWM7P4fgt3c9LZnFlpBuPeFHzJGTplEzGJEeRou1onnnuAgoaccck8aQaxg
VMVLUFzHI9l+zSH5zK72IAt6Zdx7vx9hIMyTM1reuj6ne6C0v2E+04FB/3e7069v
9bJXnRaLQOLgGC/Z1QrA6jPUwcCyaVaXpPV6gHQyyUn8z8/9VbabptMXX8a0i6Jx
/JAlasE2NuDcVSYrQjSD6FNmW+JVPyCQvuVMHH2vXNQrJm0QXrPeeAIjkdh2NNT9
j8SI9T0SaskAsxrhywsmxPZFz28EMa/cjuaG7kROvD886C/caDAUgu3n1A8+KM+H
L0kXabBVv511RFMoNSjeW001ym71sZ7rtTXxXwFz7F87WbZsh6T0lbDU/Vxw+MSa
O0LoeC1gkKh1r9OA1qWqXvGHUL0l+xSLCJ1Rviy7suaTnvyBX+fKxhWkjb5TMf6w
VLGn1eyXn95Nj517ILWHab9oXtU8XStv0646VDdHUtjrxT+10x5VOygEgVQdQi21
1CIT2V9A0CjiIAgtTFDakXj3tTdCMMnlH5f5FLD2YkZmv/hA5th4FKiiFCziBU4w
zRl0hQI7rEjDyfZVwurgq/cW3G3hgdIKqzRQDZt9nBGoaXvP5OrEcn5zHPOiifg/
4v5xUteXUoqy/AOKBfpkIwYGgrpu6yrGn46EdgUpJ5TKnMlERSfLl7Qmacj2K/qA
v7KTzOPghls9ppN7gPzE06iwJ4LjjNLNEoJDM2CO1kJdzbeUZNBv5hYcIQmBRtTv
D2VOtAgMw+1FaIO8vKOxjXP+/f35s8dfbP3/evsLPPg7ykcBONP8ffltDNTQnqG4
8xMyY7vKcVzDawQbGbaAtVYYu/U5u55mpzfR3TqRPBJu+KXeVYCRtHQ8ieY8g7mb
DQO1aVPvWTYD9Kd7z6qaAsFCXxaf3LypKf4ocsWERsbmfpS1HqJQxaXWUkijduH5
hsx9hzFG3Yxef+lh1JZ8UpXBUCca6JOyaPuzj9vvfKhLUtfMWmWNhUiQgjo3rkpg
XhBIx9ITf9GeWKzckzDIoAgPTaH7Z/dRDpHcGe80oIEOE4+BBc/DOVWf5tzejUNP
5LLHu1Tn/rNQMzqJ/6RAm3NruY/P3nwgx3vFpNUW+N6sPJ/3lPtg6CBuHeEf3AZx
jsyQu4fu4qutXX55rVcmFWQ8NyAEAxsFRY2dgNbemmJlbgSkouAkURvqQvLK3O5X
7an3+8w2Z/FMonm+aXhxM0GQOBZIZBV2cencWi/5mI3qesKRZwISD6QkGKgdDEI8
/DsrCAiXs9csPEreSlW0fiWcUcB+Rj0gS/q53UPgJw3rliXf6vy+bzwHbnvpWQrj
c+1DlkG+RXdLWJX7ABdfzp5wPv694E/TPonaZwIwMYUF3KM7HyDlJ1ATVzvzqFU+
CoTnsV549SogJQ/0CzLmi88rqxELf3B3H5V+KIrC/4p/gHR1ZVksd/gnUSYUpSsj
f+FKudxTon3xV1BzY/vhQQHNgd3PSPtKmF1bGvWggReS5QuZlmttuc2vnQ5H+3EZ
f9uSA8UfoZzDjt9XM1Q+DVyKcG4S94OS+bRrpZyKRnzhD5BczJkjdzNrMT1CIjK2
/RtSyfYcG0MfEfWDdb8drYc0T8JIQFInZUQgSoLMWp9Orqx9EZYy0HwR4uKDFR2d
7RXy+kBtr/03g4DOgYf6t6sSC1mq9GtpaeDuP3g4hyZmI9UTtNTapjT0rN4T5B6G
PNxWIGLD/+7JD6vO2mtT1yREtTz0NOmgF3jHTRYjou031egW6s/9epY7VeT76/AF
qhR6SuBGsFqqhc+FLikhHjev8/lcQHEiIrSnQ5L3Ue7dIqxboAkDEiHIaa1ruDvJ
a8lQoTl+DumxyiTrcB1J1SBYyH+ngeyxdfn3NsX7JSzL14BYh1Q4UqG46G2+XDxi
EklfuDBSe1HM7SxyY4AyiRhoPKG6TeeN3l3WgyC1k6HQ/OLj7LI6HsooOirhHGgN
sYGxwA6JY0f21hXevyx5p3GCkAZz8GNIBOYZdQKa8+hVHcvkA3X7dGwfNB218et5
FA6FVPnTNxgbVeCXXgn5TgYSUg2xo9qY6N6iK1JHDDcKt01ixMl9CVNceN1wbSvb
SYJrXcNCAqbueRh4myn5nMKl+WUUqtx96VNQZyj5tluaZR/70YL5E7tSQ9M0bfh7
f+LsO78fkoR3OXn37dgfxGvM2NCnVaUZmsmTDeWvphS7Ar5Q5ad5si3VMVmRAp5h
90TwWyTYZBxuCxTqhiC5mxMDCVJXRqV+muSlx7f/7Km8OXiS+ueiKfUFb/hmGrue
1ccEziFch3PXOw24TjG4/kdrgZj28ye63HKIIYCXI7U8YJJTKyrO3hUgHXD4jRkl
NZYYHxyBj57N1VVqFdGi/z/+7DKiVDcL4Qd78BxMj99n3EorKdtLwFpWNVWBHfXF
hlwOcsrYWaL623UHWKumC5+ajICduhSoiYzmUqdwi20JDrTvXNXoSaUzsiSo0Emv
c0u3KTfrgfAwdJFRPyf1GSUwhQXxEbwU1yJjQl6cLTiSzKqRS8BCfUgg01hs/Bl8
AYelSTJg3t73vQ6OEsYVkW3v1bz2T9Dpkd9mbm63mUcvpke8HTp/1EmfY9sQd5Vk
nuJQNX7BAyi9Tj7IconigE9AvvjqoJVFRMnpqLkrZpoQpnHg7R5cdqm/bAs9I21A
lR/b8wZ7+qT9liZvuCo2Zx8c7/3KIxSfJKPctt/TfFwNrItJyUgSitFU7zK6MGqg
6wkaHL/DMwJvHYEfVANs6pYV8h2h0TXFRzSfoXc35vKpLWSm12F7wWv2oFyfgT2p
59EN12gLBxrWA/75qpXe4tOHChNU19EfP8fwphyFthETAcuJr3vDD6/OhQbFrNIp
WqmyzMtx1MvctCr0ckUYohyP+14esZgPgsMD1Evy1jaGAEFpfvtlOWmZt1G2AI+s
KSI2ma1hnrlJDmsheeIeQjwc22/4JsiewmMiV/RDG0uKOPr+fY9QIU/xIwWq4hCe
LDyn6clLFMIq11oOIZo+ftDyMfLSrz7Xp2eCxUXmF5yf9nIyGQac+1Nv0UfY0P5t
kNfxMXa080ZvjkfHnZFH7g0nSJ6lpxOIMKsWqayE01x2BKIQioKT1yWxaS4CWhq4
dqnDEPlgH+avEb3XRNrTib8szXVAFezqozL7EvNwjqfvvtnpThrmsshsKouExmIS
7idFvRH/yrEMabT5p1pA7bWVR8X3sKIcUqfIzd5tlcEsSXRxtncH7R8gewbAawXe
QBnZnJ3MJkrcGfmHVZMOJ+96PEfHuYRtSfDZcaLtgPdOdc/XeKeFog6y5qZrmqYN
Hm9Uja50+NHugOFveO39t6mJGJlxIvltdX5ZLdSvuVPEmlMgkmY0UySW0yTUV7gU
tNd2sBTryF3sHYn1KcKGwZsW12HV6UYUw/FseaB//rXXDlu5ondlIII7m1ij2o1V
gUqspqPbSweQw6CTe+Iflov6cE9qo77t0ef4lDHazpuQi6yNaXAD4IYTWwRRtVGW
FrUZmLH+4G18h6EjzYNEiH5LPdMgFNhG/wEdiwAczFTVW558kgiRryq/mYZ7WENY
pIg0qNgKzBiWiFtX/Ub9k6FgsR/10y2aox2FE4Y/wubeYCJwO5rUqWImNwJdwxNN
9NjvMOIBnVqO7lhlN/C0ujWkoLHUdP0GWAixrH72NeQQ4Mag0/aaE/CIMGNIfGlw
GW6KYVWJ/qpMsk2n3lVQUFOk8sjn+a2W+g0TkGWA+dhoPyQ3+rqppWdG3ly8m7L1
7HVqL15ub81O5b4pEUKYWoUa49UB9HpYQZQAQsQScXJozf3c09wwz0dyHWkT2bG9
InvLsB/OOdPShP+4+bRaCHbEUJE+905I/eAtumjQJ0s81RKz6bb9MAgKHq35Lkch
7FN2OHVBFLams3JVL7i6bssJh5Tva4qImUQIkSaoMOyAfsDEALF1EFNcArS2G+6u
xMWO6TSeNoUGVQWpiWJ/KYlj5e+DLapJeliqIL7Z7lWpcmuH9sUWFYjpaSwVP21j
UgVyN8ts8eoks5yah+1nUjr+WRTzevdyFLy7A0YGi/KfyDoQ/JSUoc8S3QgJMpJ0
fb/WwgV/TKZ9/sIX9P2FqXohIpFAsAOSdsrlvmFEofh0zLheyNIszfDGmTo7ZXEV
Q8HZGwCTmRibAehTlgq/rfCpbUw+IffNRiG/z2UtD13LKeFbLPllSNG24dYYwcgT
aYuPwoMv5F+yr9HashcmhgffCiuEjKR+Iu41tXNv8igB6ZEwfzu2JFMvOylCMbAb
HcLmx3ZhToo3fDHTGW9Jm4Q9oI0k0dSsisQ1wc593ZMXMg83cNZrZDdT5mXKiKDU
7gZ5sTQdGfK0XKy3rvHbL+BsMKGL2gq7mZF4XBU+36AdjspUDS9ATy08gPaQIgD1
3p6XC0Qw9PyT9ysmXUSm2U3QSy1GWyJo+ycOeip8pLTSqsH8xxGweySGac/Nj3pK
q6dMcmtF6X4veLC1sAkdRBv+QPWw+F91XJfTmjLK9+yH3xGFoWutFEM0FbKtzLQI
eaCLOZoc7iS7zPs7/o+CAjNpZGH9ZEVzQDHFQA2dvq8d5IGhRXYl642xYgAAw7P4
jUmHgQ50r961GssEPvHfAfdwqcbfNWftK2r7/nGAZ0R2Zs7eKdGl+q0k9jfv4YAU
fxUIqPsmIRfMcelyqM+4i7Ek5/Yc+RYlA6AOl7f/RoTkoOC0ebxVkapkgRo48W7L
cLRKDadWang3ZSwTIg0MEXXVWjzvfsXJ8Cjriqkc7E5Xlj6lcxXFRbYzwQa2DAkY
XzZ918YZ/ArwX0rbAx/sywsjhX4eihOhitluWyl/6qoMNAcWxlZ/r7mRzuEPH1K1
rY/C7s4ag3sLzSWA0Z7Bhhe/TGAty/cm7zEabmbPQqddTdEnAKRjPVcfnFR5Bi7d
V5wCBEU+Jrp5qT6NA9u0omc71Y8wF7FOE1zt0AJTC4pLtVeBZFa/RccQ2ecH9XxA
7BA62OLPcrFE+WJDuE/+Rnf0DE/+EWdE3gfsyea+vte2ZOkzuDzdlZ4pArFb9qX4
HvjK1bZOVO4kNMr2KxGDWE54NDMa8PCjXSpirpnTnKv0vAKoQScsKgX6+pPnFVnk
0j+iUO3S3gBZTqVBJXtnxEAa6yOcIv0LNfMguF+ScPaKGXlheq9hzc/6fIKlG1d+
25RiEvsZStvU/dtRCjkPZ6Pa8/tGRqAhlP1ayiUWgSJFOy3GUy3GEYVe8tF57itV
8ztAYDb7CokuBZJdzfur81X/TpYXkOaPr27zjkxhIgL7/UNO8luZXrx2ADmw2dOy
ii2XA4Agg43M3DbMroZ8q5k8edBBWZ5YwbCKzD/RS+mOzesrS4VsX9pDw6bLcmjr
gnqpY5VSisxGPnfXLHEm8YkgXVbcU5ZHBsYpw0iMBFUFA5NzcAkMFJWFcAtQmGtL
5LL/SYooMtEMjXh6lOz7Ou6llCNdnY1WR2rsP3JCBrMKEvXkrerGcBhzjiFWxBcU
8n6dmuJ5SNbQPFWfXBegAczvFFcRt/uvSfymb8IpSkdrsT3WSp8dQBXsFtgEHJn4
q9w6JwQ7JMGvaGBHRCa9SWqNqU4+oQdKqkjsJeygqqFZxIzW7IAEV4Qzwj95LXac
+CylFVzSBFlTkTqQ7NhzRFID4y7b1nKy951gz5ryGXEmJ3zHNWGTATcKAjYfIFQY
6xWWR8VYrvvHuGCI7dECDXE1rfHrLHhUwHtxSF/xY4lW6qlO20+OdMlJE7qf91oM
UE5KXQr4+p983wT5NFKTm4uoWqbw6ylHBv5Wv+sC4EYQBH2Sj5SijWORyuoMVxTt
+Ht4Ga2IcQQ03gGncDA6mY5NpJ7XaVLC3hQSKqau2Ogc2NfyjMkiKKg9Rn/0HB1w
J2jKc28oJh24DzYXtCmILl9SFXit3p+LrxrT7WngYabXuo5ck+fPY4kzVHQc94+Q
vVrWl/Co4lzFv7KmoSdVQAY8E1jluuW7j20BgS3JImdZySt02svVwgxhGDcQVXKD
N54d8S9sD4v3q6LOevCi+AuOtKfo+ZnETENbxwUja9kmYkgDgNYnCqbFd1mgNPrX
7A+nuD+ceESQ+Dlg8wC5diy+Ce2TSHC3QhWt9LF7jn+mNtTZRQdvdNwRkXXJPIVa
vbMIogNw6SEDpkGeb6mGGqMam9Cs1NPGHI0RYrhogaGCtiUyggSA6zY5JW14Zbdq
8eklciv3D6NxQpZS/oOas1UQooUUm4OsxUdDrXQFL8Ouxbys+8oA9tItXWgmSU8J
qt1mAdOVvvjg47XkjiQCjhKtQBOcBfPmVu3yZlzbTQN/ys18uWwqv86RTj5nUvwT
WZe5FmKGRyOoznf66YQfFXmCbm5jJZavetP1XSSXYIHZhcJGQ92IKyRcOJryScTV
dVdkl0JgC9zFKsD+4UvMS/fAzpLLn0hFNyBP20f8s3YZ1TGkqj9WMgW0QJpkz1+f
dMWyuNrKvA7Y5QGiG3bO0B+0C13zIO/iYsb3zyi7PURISMe89WZkp6V2JF0lzT/H
icirAQOI6lOmYZDwpTV3Mv2v2PKHQ4ZSt9WoJzSEv7Yw2/HIJv48spZf3BWtzfEN
q95haQfQA+DzVUgmCqoWYzRCwWxjk59Y4m+hmEw/Y9rtPUtTMI2S/h70kSVMfuOH
wPZffXHmvFygkkZV9Lqp7MRvpk6hBtlS3YB9QutfZ/dfdiULp63nn80/+b5ILn5V
WHHIwsNCdYghATceAkGVT8LiwdD+/Ibn0ZFxfxsgW4OASSQ/NclDXQDa1W97P5Xo
+Gs6UP04AIBh6s5uyD5ByU+4VLqGOLQrGat7DIUcoA7lGD3pmotTjcphivzG6c5y
bLkGiAxKNtYqyu/KOGXGZx5ZdBCQ07ZJ+m/l5dhz9wt3sjbC2ui89nL3PhINdUyb
Y/O3HkeJ1mGN6b67MaZfoa8EDtGa69q8hTw8lFMz0WFdN+X+aossdgkA8va4i4tT
jXBrmkQZApZUR3Hqf4mzl7rvlFYp48DwIuNJEIq/U30dUksiyaSGXxkx8jmuqdjt
irW1acimOe7Qpmy4Z+YbU/JfMR1xtTRYqs1xgd3OJuU6ur+xyvC0OUxmhUMLKp+B
CYMRPWReiSAdyWRlpv9nsVqgpQXGCYxHrVmUDPs9gwf11zsmNx4GVQ7jXidA3pXe
PnA62JVb5/BTBTQCfY9ph/rcemUnmg+T8us8WkY9wtdbpY8+q1qEMUcTcwTvetqV
jdxRQdeBQ1xALtJ1+pZ1nXh0Sk9NJmbkS3dN1gVmDBZPWbWiK0b8Mt5z6UtqH5c6
YfcAYmOv2I8c4AwuctgT+LJGGwZd4h/4L+2mSVrB1wGRx51cGkNeMc+JmnxXu3+3
CRILqoS58DZgdGAnb06i4VF0BvVj4CsUpolFBWmmQeWnXFJ65fUvTqiaQ1kx5unQ
W+phRodAtokv8TH7kHc8+Z0Ohmam8jUJwc/5+Z69Gu1Qpg/ZNYsCRjLoN0F6rqkJ
ZGEeUjjBI0Wgdx3xxEafPkc2NVQd48TdstBh8OhRL7/EEIaqyV5P8/N1RQkZASRu
2uKKeukm8I8ZUm0qf/WGpd7SefpFRUcXD6tYy1VdwCsCVwGYUufDXwJstdUZmqkD
jNW/n6bS6nYeG8cud5okqtfepNtzXY3+A4xy34MMHeEQt7ktxDtt2AKxUmvUEGVF
sgduQ6r1Zp7XTIp4nKeZTVXrHFUUH2uBy5fwzFn1jEiOchKlSEGEhizg+0zgaAQQ
LT9v//xJCH4a5SITV80mIe0jE5OlPm4Y5N9B6V3TQY5MKz0jQ/hIc8IM4CKH3kOu
9UI9mLWiru06Y1KSXe4x2hBgrRB0/ClpAsfA7igmL1VWdNn8qI//sNQNq91OHKG7
XQQfFnPNV/orWo1QagdQEz0Zizkn2EQxQhYPOoqSvOKefRaNTtLMsf+nqSLlUw9M
crISc+1d0YRoQWfgWX/n3adrr+8YojptnjaKP9iMTY6SRgTioTuxOocomKC4aGiF
kuq3dnNCVe/9T17ujPmox64FgpoDeBZlsF6eNKtHFCNGnjC2d/pLvad+Euzzk/tv
ZBllrj05qfsVogP702QFxyFDRzwe76+uv4RuT53qAh37WZTxQdfsUAkWkxz9cNrb
ewQEEoclkfLLLu9VPvciBB/os44FhXTFKBb/mDt2TVDwyZOyRpI6/vge0NWlzXYI
rMnJ/z5YmQB2a98QEkFmZpB1A4pcomHfAxGjB9YfVDGBls/8AcS1Tiq2BxETDMZ6
sGKunoIGfDYTmP9UFOTxg9l4//dnqKbJOIKLWrRDKo4h8gUdlu1qPfZ5ktdHPLvh
cCOYZq/cetLgaWtmNckugZQUpUj4eRJRKNrKCgvSFRdTppO8k5CYhfO64OW3qLFq
SrOGinAERc0CEHdmJ2sLNZZz61ioLJTtB47u11EXpXWMrteyrQTMPsEiCztNZOG6
Nmu65PwFlaew7B28e04adh1QfGM2zktIMYCKlb1Di5CwTi8kRxPiG9qZ3vdi0OHI
T9RsyjRfpOSB4Uiei6v+Tm/82ogMhkdv4t4jrEDJWaNY3yHzkZC0AoaZwh576QDj
kTcHPlEmfTWOtj/ZcJKxm5Ug1xQbdRLWXufldmAGZJdSXcEaGxrlJ0fy69SSguGP
xsNONdqySEsn6Kw6+IOitqkppFJuA0OtU+WveXspJEo3t/flEyNSpMQU8SsyT5Jl
9hlFP8wLxcGA9hUqtOnHzdSSqHrYd+UIOgb6pNblFp1wlJA46uNBIfUVPJT1w0ar
/44BeMDrJ7PabAeaqnsgv/b8k4Dgat36sQ/w36Zp5UhrMoB+JkSlTNM/hESpTrRl
VEepfBQcoV8NygnNJGjPg8k4q2YgSeNxX3a65I+XR/ofd06B6gPuejlw5u+HTUR4
cr+vMy2HLXcs+21/clrCEJzcde3y4AtGAo59uAEVrrAtM17VOISMv44Afyj3br/D
JQBoNwG5Y9+TUQI8n8fpZ2EbzLUm/3fpgDqFPUeebZLGd36jbh40Bv7FN5FgcVcB
QsSuXt+/rzreG/TkHMzh2UQP+/tXvFc+9Pcz/Anb+v7MYvot3YLMt5Nh7ZaZV98I
WNynP8oZWD6k8fWd5y1SJnQYUpX9KGqzJXQZsRrMI7vlCEAfWHCQpscsR+27Lpor
DJsOxoXAsORh71+G0ri+J8y+GBfWnzrc0FOj8cG6oUDEtnNKOWpxUY8tOGvXAvIZ
OziX+WX+dZU1pj67I08lS59kp4uONJM7G8qbbBMpqDrpnihdJqtDH5iF58gPR8fY
l2YqXFqTdmeFKKkGndcLDDaZ6ib1QmAD5tRvZ7VQbV3C+SnXmtr3/90rrKSPIZE6
VlMzEqVdN3l/jutocex9bqhzQYkI0Yg4vVz368VXgaW77M96CHwtqSSB16Azm88+
v11H60dIlRBuGzTx+HoM9TD/EBvNesVl/uicLLrO6Kvu8hD+Lj9dusE/ZGyyRDex
GbPjZfDy+yB7sVHohuVh2qp2j/2Yoeppip6n4HgAwMihX//KGcMnSvFy2kEPfcIE
+sCSddC0l9gWWh15HQuYcQDj3RnwmA2xLbgibeBJHtOPKCUROKGw9ID8iraBhJNH
RvOOQav27WUcoxl844NCqAI/aFZFr1KFKVci+Jon3G+Y3W7dkCHTKXDyN/sIxsgA
rKaI0Qcw/qj8gS8fwqzXgCER8LAZ3xerlvm8xda0BVc7Hfd6mdK0mQ0cXr45fQfq
nS17ef7pP0CEN/wWj0eJ9J4UrEqpxWMK3NIyTj0du5bA1ZDjR4zRoK7knpOdzTL5
3lwli+yv3U6YsYCoZlsiqGly/5NmBLH4vJ0/vGKpVAEpqevrJ3PiVP9TkN45O12f
kACYNSc0yhfbeAvfBH/favbLcWTk6Tm2lUIa64a9vaOgyaQTaQlLFaCF4OIhkoMs
K4ZN7ngZkZNAc9Fxk1w7FWJiAJJcen3hrVhFaYhGN1fmsWgqm0N/F+IRC4Dqu0n2
G9AF8lkzdp87Zs8zK0F7I6dgGUMjo5noTgpukSPAEmfmLTp8+NyfsrecIEm0s4ee
v3gFZ9ThIcPvmrzga7ywjiscCLh/r2+6qBwztkhQdmO7FXpVFouJvZ0dqz6Ew5nU
m/JBAXSa/M9n0rtTB3HY/+63jatk0RzHbif0gbwqBd5SMhLELsoNRsBA8leVNuZc
wEsWzJEExIcfTNFjiDoMvt9Y4brvQrO/LPEZ0UU2Y/xR87mbsQYfa/NQ42b8sUWD
7s2QxAaa626Lelalb1C7uiMT9GwZcT5/YolXapqMKz0uEmNU17uJ5lWg79J+MglU
Zuv3cpkrbZJQddmU1aa8SrnYbAhLBgIIJRt20MABLUnc42ZSQdTNuwgqUbCjnNWV
IMPMnjwUWWKxdy0BbjPgbYX8jElRaMcjGpotDJF5AtiRrXTmRTxgV2zAmlLyoi2k
BtwScTBUfN41/88jc/hMV+O+XCVD88bOw/sv5LmZAq4fD4bLj2hRVERszJvhLi6s
TFmBaceRNqW18KOiYffl9v6w/irf4GW/l7riUxdqkzuJIpCnugy/3ZhRVtzqJrzf
FGKSBAQHsK3YHAUcPAq7YKB3CGelDvTfudCEyQ/O6u2ZYg9QseJF1prvmQQI9RgP
N/GVh1XjGBp+Clzdeii8gp1RJWnxWlhwKkzJkIOwYdEMtmk3m//XCrBV5CTN1pRQ
3byrfj3F8pBozGB3edh8DetcPa5ZavdLh+gQKNg4y8O5hB+D9BKoTPZdeel7cxl+
z158My3JPJRer0vVapqTg7voSdc7ktzvOb6jb+TV2qE6S2S30AeNTJk1EkTw3Eum
BXj3sFkOouDaPDpxI+VM2DMeCnprzKerxh5s5Sx/lJR0wo3nkwep74K55vXh9Qga
tsTLgswon8DHqkP4F/GLJM0SMm6fOEVjqa5dLiL0naMG4Exl0P7HqE40Mk8ui5pT
+rkfmbpNqLwoOOyWBHXVazGoTqqKEHB5wtRbaClqv04t1xXYQtHpESiCEyNWT523
gkE0Pd9u8neCUSIqc/9qY3HLZG59nFGerO82baGtb2+lUtzrnbd091vnOG1Awv/m
brr+N37Bj8QzPispyzJJ75TMuehwM0YFkc+XAMP/7vfeAZVE1OUpaIboCzaR7ovC
iVeHX1qFRGF8W2BNhmvm1OGJtzWE2TIq8fbY2xCjwS9HWlYNVlL4arzsO/Cx0rHm
mMixg1I5SWB9SC8U639dUur9igmwFdSGfry560BFLjAehkxrHMy9RqoWVlL3o2KZ
WrZZObz9pzZCSf+PsMvOkXqR8BNCUlMqkeCjmHgnw/aCwLEjAVDVs1wv161nXmHs
vK+5FXfPVuQhoO1YfngieIk01PgVO3HaOIvjri/XXRjjNinspGgpEcYY5IcW52fh
swDWPysa/s4q276Lc5ncQJ/RjjwghLotce1hCXP/4Ep06vbffb69ikCmKDMz82nQ
kX/FSrfCx/+83YcFQUI6m6KXh9hzz+k/xrMr80iDx/SM1pNADLOh2wHY/SNEJg0w
3llYV6I0q7v0NqlOltbm6qKlYS416oWiOko5KYfX14uJHSP+XobpBpOiPBlzHe4G
jm/GSpIl3EQwuknHDc057v0FRY8uzipmZKeKK+Rf+lr1U1I1bQ3J6SIoJ8KLqkiS
L8ZiuU37oI0C0bjTpc+CoEffMPYMksaieyxwf51SfxxBGI4Jqez7j5GU7wCfbh50
Lzlrjzmrzw4ycDUsbvoREbHHAijOZVHzEwyZKVfK+j/MWmtKEIOLOJAVGGRjJL7l
ZFLrlc03a5coU7Bl3VYyX78XQEfON/6cNygeRSSxzM3jAKjfowD9cCpv0tihSTNI
/nbcRVmWkCjcB6qoaQgdGMXFgJZgycl+9Wbocn4Evv46GcCTGMFYtdYReNNzdJ0I
uFrykSRFCzEwr6FcuuXJWGVzyrwzTe2AGJ+qgAxuoIC7RkX+sFVuo9yB2VQ/h3qT
21dov366MQ1gAshlK7yuRivGz+0JQYMv/EP1invr0phMtX+Z0M9Iy/5d9ZUWmrfq
1J3HMoZcLGmKJSCNuAxGviv5SfiBISxqEDBAC8Vbl/a64Bq9FmvbH1QVrpUwuw7H
56JOO4brL+jBCVx/5b5E3sZMNVW7RdQhFnEdk6xntzXht3w7J2Txfaom/TiVL65U
Yn/l8/KBNL7ZrN/ZBlOqV6EVA2Obgw890yC5RmRcb3kbmbiVjyY8Kzu33vQMVZd/
Qeq+6/Dfsbkb7G+ANz26oj+gp6qTncByR8m9OxmR910UrD0DlCmsrbaXKOeGIucZ
O1WCDho/qNxZBD1oDtS9kWhGfNC4Aifh1qYY1/s4F0xijRJh3zlGyEKR7KmUtD7f
1xmH9ndX9RQD1QNZyb60KTsinUh4nyCQ151wVBw3rUCXNToHflMXNp0YcGcbluDb
52BVeReyC93v1qcgxULNc0K/D4lMedkvOktev1Dp0ZZNDyFdn7slNdXFnEWcRJYU
3IqQpagP0nbY0agJe9wrcYGHKyOuc1HGJkleCmQk0CFDMNjBdvZrDuvK68vMX4Rt
ouEH+SEil78O91AmXn4En3+GkOyt3jipn+TXWcJt7yDojxbQMia2qnVvEwaJoQEV
CvspGMl1zPsSO8vuZO19mFSnFxeY4l7Uv4oPw4/fALW6zmUNwJgJcl/Wt7iwqpCN
yDFhalJsy4Ghb1hBZQTpGuAqPSu9FzHfIfR+RJiMtQUZOeslyKzQ6TB+1ogXjKDW
F511LZR7c6cERXZjIeTbjtP1QP0o7PO1IybkSIiE1cKg5s9FwZNShV4XOxQrn6ax
p+eTU9+bIlusoeWI0lAU2WTs0b/64SH14ka7j/3feTvgEEVp1E5rkveP78DMj3qd
0lq65v8RxY4B8mkl5SParu/g7pzSdsPhbMz3aa1xdKeBS+RaBrcTZ3FT1VWxoerA
6tAvj7435dJr5pOzynveuxaUPs/v4MiX56OtdV27ekLZ5pr3DlM7c2e9/Vxrn9Te
diaqBw5Cw0vBxERiY/S5uH2wYEHI1/sliMMVLOOgygR9SBjFO86YackXHqGUaX50
xF1SL/UwQni5x70Rc7fa2O49lmXmmZIE4+cR+G2cr4129YIF6iZgbSMmc8KhSUOp
tFWiWZTnQw4CxWBfvHveLv3JqEP+cqFhHUV7MgYllwAcYVjBLXPv7zsE98Mmty6d
R2lDuiPazeya9UNJx+SuiAdyyec5jCCDvbnoLkW7MPwYbnn7zFUTMc2vLsN29J6c
7TZ4/s098JVkn9oXnnk6Vz9qaaqKIYhU+R1s2G+LK2densN4ayvPgH5/GVjtxmxM
0vxn67TBd6nYKi2vDY7vd+wQT3razNKeYLQ+/Y9Y5gf2fZN6w0xPYWEXExeMz223
iQP1Nh85OkiP2Odmly23977c4Iz9Jd9g4aqQSM55Ut1XMOVIB/9dZnNU18RrRxqs
SpARUvoyyI09LLZbAOcigt2Un0mjEe4MQSlX/J15GTF8bL9vXDNqT2B8mlcaZZEa
Ks9VRfofIY5jshYDPudMJKiNYhElnKzTZiAjAmIAHSAgJHgfmSdbdsvmz5i+pb6F
8LBVgIRLXSQCqVVpryPco0CBtZS0taOKKCLECJahJfnxVV6nHAjlWKPaHAphBa/m
/dwSGw6JFOD3qZ0T5stLMvJvJWYNfucZGgsDkmRl7NxBSUxOsgrPED3ac/4GiJp0
AQB5kruiqWiwAcyPvUqzkFaUtyP8jgzJeAzvevZo9cR8dhucN1Qc+ilIE/ABZv6W
9+U4M8eeuLTp+Atptqd4254iS4EIDmzHLzUN4Hbqm0spA/h4MZgKqb8oaXWhP53Z
EErsDVvtkCJ0mHPRDSpdhBsZOLgHHCgNK9/ZPaojIOOzJxsVIuijSxyBu2aMDRDc
vs57LoQsgpUHzsr3N4tBAJsEjqeKGYz7+vc+3mu/azXj4CZ365E7Q3DD/oc39cwd
TGb3VyU6fhIk7lAS8xXpKB0aqzs4z2NFhXnKokJ1otHhAVBgv0stAd4iyDG8fXq/
XTa9k/IFyuFaYe87HEZYiEDWNfr6nQZE6JE5Hy78XGQrvfPbH8yfKJEjMpwYC03q
G2cIRJcpRESXZZHIRmlb5QnxcfxCbDrM6MALLM+xCr6q23iFclmsqb+AFv8DjLRL
T2W/c2DvF2a+Ft+W1t0U8tYnc4wLv7Kbw510YfhgTuLA7T0BzomvUsvWkkanXfxJ
zgCwv6VySswDB9xXm8dAdrh2FPVySqKJX5eHBGrM49UKGXzvd/mEJf52f5L5J+e7
MfTBqScJ0rJ0Z9sCH8et923jW3VkswscFfpqhNvjwJTvQOf52NESyYsK6dd2v8Mc
GgNC9p7t8d9STiKNtSZK2WhaO5fPnlnSJPNeXl1oc9UBrUEh+NjmV993Ib+3UNb9
Vxz4AY5DtyYDGosPvOWmtbMFTzrbZVNcNALrHaSC7UVQH+d9BicFaZ1+RwSrTofj
FSbriDpxkMNiHiGVxPH0m4KjWlfE9/iMAG0reZdBupsK8UQvvC/K/kpi8KVI8iVc
4H7i5BkuHY+LCCgxylAqgcsYldU0EWwM+ui7RhWKTb8V2NyEncL1tBVjIDztYf+G
YPLtQTwzUUC8OU7tJyuY2qPxnPKv8xiqka2U+zirdNTIDWkxO+6GW008theFAuCg
loSy1Sf90huKbbk3bV+NyK8qrDpy55GKavUcO82EkJvDm+zBHBba4Fl3Bq3EnX2C
fvkQK56Ds6xLDM0C6f6jLj0g4pQ6/k4+FyOV88yV+XnVpbLe3BUTtjPWuGYGGIfe
1nSkPCL5Ae0rXjgBngqwTAFUhjV5Fr7hsiWIzmfCJ9llxNNDzGnDcDiAc0cmw8vZ
LACIZyFD7UtsGktAsVMpE1n/62kkphGbTPzcJEJXHMHOoEscG0R03/pCZQnjpHEv
nmjC+scwH8n/wnigpmUvwiY5AcQy7PzFd+w663SnBEvdYxXayXK8Ii9YmWYcg0mH
ZFj0e3YimQH0REa5ZVMNMDEjEe/OIJCWWUcWFzq4jEMwsovTF6ZG341Gdt8tqX8L
aDJmC/3nlNEuT1Ul3onKWNWQmhZa0y/QuMHQgalbqyjWa6o5ObIFtcSAsX5WmUtw
njumeLNLJj+I9fyUUQlRctIeiBq3oVU3pd6WzHxNonMBexuSQCDDaIswlYjfJQAS
X0hzOmjwMSH23FaNJOnPTUPw5ymToJMalUGe4HUlrgIVD0vy8qzkU+6xVa+Wt2ZY
DiA5FPlFtK4XlLss6Ufdt4Sn7lSucmQwzQPtlZi4zIFUQtTqHpyVnMwxDdorFBt0
ypviNjNQ8lSxBNvUt8YTjev/IfCO3LXWK2EOrmWrqMXaIXZynoLj7KwmNZO3p10G
cMyoePPVktix5xNHoQk2y3xMdWzMf4z/N134rLSyz05sT3LBXIWby01xvxosZOAY
xUatXLra1WvmnneWbxzAgnkptkKpqef2IXi8cQeyXKowR5kiQdD0SVLsENexpMsf
goSPhTTZGAQT30NA7TQGcLY4K4xQVh1SQ+/TwdOQPndeWEKY+qtITvdjEvLaN9Bf
X18vYV3mTzpM26UCq+5qSPy0QS5uKzriPbxuFAaMdv+2Jnqz8v69WBBGdMq8st7Q
A1MEvEPRGa02wWWu4Zb/se2p7ewI0fP6Icy9FFHKmdsid/a2UzhmRck1xi3599em
0LEPtBOdb6pQ325NVdvwTUBERxph12V9/aTcF8/BcIb4ewrusTt7qmhH5CdzuiOk
4Vui2j80a3iqtldmYh21txYr7pKeiy+ermRV/w2MJ/qILQGB/cfNwpBghTlAtzAC
xfuq5dvs8250nVmhH55fX8cpKJMXDoQbrPzZvX8s6gA/oATOFlLs1WoHrHTkXBzp
6CKARIVwZMR3BSIVvdc27OwPfjuKTylH6SAci35loaquI2Hx85Z3JMDlmfB8P9pg
+zkVhnDSUR9gLOK2bFEMNyfIkemezhbfwz+SUUdSjMD7Ow4Q/JyuLpb2WzJTJ+oG
s3iGoSHM9i0KJ5bmszNLsqcyRwq/+UKY+c8ck3OZoMTWFi5/V9mR+eh7lSQ/GGUO
iRfTjEzsl9Dmi8cukw1LvajcdZ58aPQvogQxasSMLg4syoWwQUK375LFDdzzlBhv
OhonhkbxBsm2eT58dh9YLE9sgPCthhi6Pl/pYkYQLBZGTHTQsRyvUgUxpwt0Y7Si
A1rXuGZqf7Mv1awsLX2bJhU+r0XOGDd3MS30JaT8wvVFx9Qy6TMc+5ZJrLe85/k/
U80brZqEbHoC/wL9Ifs6ODIEaFLxntA9yFYDWVQmGNvxUuGcDE9eAlP0UuBpffWo
h187AI2QP0Zd35np6kZb+Ts8NFxHdgpd6H+kkoGEdQVl8rbQIcd0GJpEcxn7iP/L
Fxua9tzOBn4ds64EDYzQtnobTX5yB90dZ4tSowwDVhN/tIamCxmsDL5DAWjbPLIh
I62Ea1xNhJEID2WcyWHQkxTj/ITkMupaKvA7nvgsttiD77IG1BeCsSQGmvf/AJue
14y86aCUi0AZlSJAmhgUGUjxUbE2SJBLo3l4QP5/kpJsFLXyHM62KtLwnxUWbwH8
NEVT0SxcKUyb4VxPCLpZTQJr7iFECdyPxJ+Rm5R8KPB1UpHP79pi5oXErWrEaD+5
u8XBVgGYQZdB1Oumaq+Kv5TeKCV3NtF0aDR9x8h8gMMruQlH/4fxf44xB7XyuQLO
7n6tCuvpwcbmJbh9ZIV2Q2v4ed9koQc+NsjSFysCTYz6kqUtM1kJh9jUiEOLK7NH
njIoXr0bxQxGgEQnlp0dOBM7kyA5tSeHe8/ek7AMuaBbm8sVPn9BbH6+77++TgdY
G5+XQMXO2OyMt7u/2UpAvb6spWnRvrJZEbPYAVw4Xyni6UXYWgfiEZPPaR+nJHBz
GuhlePp7tiCrWEAVS83sMG9ZJDuf2MITDow23HDToXP/mvvSvK5sUXKURRccFYrj
vaR2jMraGuXfoLCIu078lsOZgHo8pvoQFTwnD6kWtWmacprnlQi2KOanh1kGtaNH
kmXOZKZ/xmLN5gKOCRFwo01medZoGmFP0rn/WQU/BoWKNxvocF+JEzHGDs5Cfit6
pMLMeKYryZhnMTXPiyHUic+9obpypulDL6yTngMMcnFTU/SfBDqcqj8YaoWwOnfi
PeJHKn6v1Pa3lYh2QcEblC/G/IODUh6sW0DGthAIwrTUiEJ16B55IMGHdupIwrm9
5b2MrSr4fc/TJK06lrueNrftMhwlOkcn0psdWm09k4gGI0rfMvT03Yp283VkgjKO
H1NypFWgRSV1Q8t7WXza9lSeXRjci/lHHLVvan+BqapyKg5lyu0Sdi3utb8oDKeo
C8GcT/Gd0U2fl0h4eWc+MUcmnMIuEJlb1PxB0dCLLufK6qLXOn3aguCt5B6tIOsY
pWhvbik6LoImh/2kc3tzj4CisRFrwHhx+pdQvQM+MIPafQm9D6f6gdJ1jJ+TFvYZ
xG21jBq2llEchDu00csJPxZuU2wYYeQ8m6fjtrw+IbjxMVsvx7GFywoFpsIAKOex
JYxC9SlOoZe5qXPUUfrRTqRnspOoqlqoLZijWI9Z0jMkYp4lRav14HjKeLHI8dXu
/OmJu2adVkHZ7HAH0tjoj9Eno57Z1+y/RbrXDoj/0YIxoRcILj5k1Pfzk8uTL5uS
azJsD8NfD+5npmUTHATIL11L8mbocKPjxIMqLjwaYevdkDNBQ3WQIljYZPy81bv4
nrDM+snhv5C46kTd9q9jzCxSId837iof5/nV9DH3LMq2Gtwy2jISg87LtuGJaS4k
HS3u9pPjAvhflT6XATuSnKvZC3pE3l5tT4+lSBSCvocp0H/oI8s3+kQ/VaFlFoVv
l31T2dEwA60//bIhN8boK0kzkfFZJFhAe7VbuACgUA2Cj1/IW79uMyS1em8pTFV6
gGpEQjBrc8FjgzEI966i7vchEALq/r6x+kqux7GSPp1nScJmNPd5XN3aug6mj81/
G7CgILW38SgtcTs8AzyxQFnJRAeEvCrTs7IwGGaXNmiW6pTBAM5KQPWrhIfqcvLO
ihYC0g0zc/2TyiEqTudmaMalYLzH2XLDg+40odbxfbA4D4STcyPd1mQr9QVrXWHw
evrJKWRPkVOtyiQXefz58hK+l4bXV0mfjtm9wGn5uNIzEr95bvQQF0FYlsda5nfT
ShcRbTSqVt4ZipW5RTi03Y6ddzNAbln168LBb88zLebvYhO1p4He7ejav7kl6mVG
/P6+/FgD//9X/mlueOYP8fzGHGvE4cnvwiyauJ1rPxXoNvpUQnWLwOAEzFfzyup/
xKjd0JmHqaYMl9tPBhQos3hTZFJLM7MAcDKOcE0WdFWOZTTCiBlmR25T4wRoa8sE
gkjXDBbvYEr1wSEKUiuONJRZ0ofBStbBuv6/GWYtwcgQOeXBh3Si6DMR6j7yh5yR
Mjn9GD/XSsV1jDJ6A+6nVCm1ftnZomo20MeMxutSZ4MwM8wKBhgsYnVQxXCLfr13
9WrTJfLnh9bf8hWL6w6PQi8M07lQC2Jlw26Z94qZpKbBMORXluCVPlFmetwGob3W
gIvt2UwO3Vr0aJbs0NqaqDibU/C21LKzuu1N+69QtzVsb0qfdrgsQpi5w5fIz52l
clcvgJvX1YLtSkSblgkqHlaWlAJRvWqANYkdAeBU4rWKv8bJ5SS3HA76+vYEX3mw
SdzvyFh46762/iRuHZygMkCC5LuxUqbE69WID39HFw3qf5EoS/2cr7nOyECHaRt9
kUUZ2LsEZBCoZa/6UGx65+ljtctGkemmzf4eFPY5PcKgJSkc2fR5YrRO9zUvr7Bx
Dcj1J9wQYs32mQqVbtgKy5EOMhAuv0AkhE7e/D/n+BfxHoyf8zukbaH5rjN0H54t
/LRIpfOg8e/EtACwPMys2GaFUhi+H31WlR5B7sheojYOic1HZwlG3tGSG2719u2F
uEWjFE+iZPUg9U/1FMWlFvAfor7NyRZABvZS/wi0BdatQ18/wAwhnz/aRTe6wncn
tA6uK/Jx3dYsgWVFExfLj97aac+bqxoJERWuuDv+eh7r9UAT5sRIVfE/QQbmmU3t
dC+wQtDQvriuisF1NsHeOQYN340q7BULppfmly0KzynyHhMiz2MZXxBLemissw+n
1FBq2plKYcxY3ChLvpcnDEqTedqD92nje4xQOiRdcVk5hfrNfJafJvRF3Y0FGPIr
cwbJVMFby52SmoMscba+z/ScRqArRxo9p1Irg/qJFsw91z1NpNU3ZrLjzQWO39bU
t5cKAw66Ubmh3F+QqGt0R7jLYTgXnDNh9PHB+rOge4hN2mJsRjbt8UHh7p1Z3VVk
ohJvbNliSuwAJKkuyZIhdACvJe0Q+WS/HiM+uUnoYZA3vR1yInm3+TaEW85RwqTl
P91Hv6RUBg80ZE+aXc8T9pZX7tjzcMqI9rFdYUbmwUBwx2wN+hHKflK5kOYslwMI
FDU/Eud2G/Sjx6d5LrE8ZCJe5OJywNTzqCGOPavzweGO+r0IeIE+fipaE+BePC4k
IxHZRWS6wwq2iOD6Il0owvJsHDUl3X8HP/Yg8EwMBNDKOlVqVeIZCMQiRsYOTbEM
WnnBorG5RmxDzZMQpa7NLxrVOGMDjpuE8G5Whvfxd/CG+cD9Lbb6N1WKkSDuyTJG
NLqs9xFU6XjZ0B7JhuE7Xm3JP9/JXk658fj1xNaOc7VVc4qD+modoN76DqaJubD+
GY1Y12VrJhcG8wWszgE3lcEU/2wvTkESSCuJOng82XV99TWtIBgwvZl6epXCU/iC
ZR8hFOpS0WtzyVlD/4IbzFy5S/JHjYXIbl8KOdWBk7molN/lWN1dS+UcZ/TQY+3B
51JaIBg4mPnHUibUKJw2aSSi9Q2FSZrVqSFtIMT1+cQuNTEWYvZBV09AuqyZeyeA
8AWYWWJqqrRezjLJ2ErtC2aCIOZSLa9PIVRZQVAOY4fV6WBS6+k66nw/A+Wz44qP
b9hnjsLzlDWNFI8ivyTQzkkGI2wwN2/S6vEsdeTbiBWDzRvrnCuT0whItidQn4lx
GC9/pTbJE5C8DTF23ncWSSM1jBXP2cJCAJ/qmnPwthYRCceL7DwY1LxqrgCJ/pDZ
qClZIJRXIczVXWcXsH4IKAU9g5zQzImWqt/iLY0CnODRM6Gg2hH6WgtAH++BPO1w
Hg6Urhpq5jFsCTWCsMcBfM1OXLF+5FodMO82GNeq0JoPQaJmNtPZpIvIAXqwFtsA
UqxxvG3w9RCaWGba308Ur3OrxEPS2CPpin3DPOkIA2Ikl20PC1Nll4e7X6j9R7OS
4AQMubuMYAy4JHLg/c7vo6NkX5SqJTWJPpfL2CGDrQagtqwykt07o5HB6L22j8+B
bI/IvOtHjNrSQ1xjjAoAacRLV1UOxZQNrIZM6LaUqXT1Qbw67r9edcV4mrQMHt3I
oerqlOhFVRxDH+VB50fcKCSm48dKssqhqcgcUWGJIXEcz+c1voCMcQ3q6feNEiGm
uLC+lmOaz7S9LVBz1BKkSrjy/HJ08ZimqwxOStr4IHj/dXYguoJURABHppRPeFkh
TlZnRS9AFxQfB5SjUPDJZEnUqlTHnMujRT2jKdPmOjSOvTeEXRi3oEXkaaaw6Nlk
hMOgNkr5Jy+kKpXpeJvW4vCZypJZ7avVyspQqHzHsVDHzIPTY/KIUkySPmjYffAL
7pHGefRU48Qo//xW9nIjJd2mS+ggH0+lmhNu2BLu8zyGROPHIdEKglLk5CnqeLmf
w49LRL+Dy9NQ/EexKOfDLx6ddPRbxK+M45/0Zgm2cBoDh90zXPyLn+H9agLAydjT
H5r6B807Os6XsIFGW/U/TIoYQlXqODHHF5snchfENpf7ggFEMaMFp4p9pZw5BfLz
I9zwvBCkXUzbJuod/hIMKJbyEg2G1Nb2fPPKWosm5OcMxrYeUju00HAKenn3aK5Y
974uW1mXvPu1eD21tjvikY3ytpxFgLfCJYt54c/+Ad9OzIDefdpFP4eLvub6OW+g
QuXKyg0zviylXisSaYUzXXSn0gVjYEX4Rt1MZZ3CteNLszHo3KYp1I6EqiIB2vzz
P7HGKUM4t2d7shpc4BPlvNtHzwmpsYcCjtro9qKvph9cep1V9vHcmUejG4zunrmm
rVUv4Q0+punyBBksxB1FqlypAkH+h9zh9ZT5VPqL8mX8IJyCgVms6sH+G8o06ZlD
kiYkhUpfp/lf/6M1yqmMLyW0WakH1kjyVVVoZicl8AoemY5/vkysTGUMdCbKMN0S
qQhlfrcXbFlKiklYvynfxpZpC6gNJV28JqXtCEiGMgPgX5k2+HrmuWV0KCnZ4O3m
HKo+5Ji9jgTE/6hmxWnS8d8HDHDiEIArDhtEgsn27RPWmIvaYbPeqM3w1vEwCNO2
Om1wrNjxxTzFAQDpcyhU+xM/YZK7ankOmTiASqfeajnv2wuOCXRX534ZB3u64zKi
o3xjkxFauk5jrSWdimhvFhfxuxvSJPhPhkT+PyjHvqxWHabnWVQ4W9jBeYY2V5Bx
1L7/ohvAs76L8sqPsHqECibiQqNDE6B327vNzSo+ULHorukbU/+ETay2aSesjcJ8
SHvIzzSfE7UsgT74vKf1wuQ3n8cCajlKnEM/Aikyzdkx7vNwICC9zcsw6+NIC/MY
JTWRruQeypYTEA25H5kzxf4tuaTwM85r0/xSS53gCEHyTtYB1HOeA5N3bqAhLUiT
sg46Rl8ax/QZS5xBZAiQUgpO0ClJ5K3fokb3whTXOl0azYDpYmxXcTWZ5vuvwZID
c326dI6QQs6yavU5u9iXGeycTAOFTJLU2bmcjCZB9ZalP7jPAus5xEnXCdrACq1P
auXYVZYx547Z5lfi0HXTs4RZWznCm4U6IwJZgerSx0sbcX+Xhszi1LgPHSgNUc+Q
BxOrrc4duEDGnIi8TZLhjlmbUfIOslNfn5h+KwN31KwE0MbvV8f+N+OlEtx+pBbG
GmJA6Ene1dc90Ywe70/t0I080fgOAmatxCd9YFqb1Ynm4AMFkC5qkAtnTlJK5nxF
7+iD/p06LoIj2MIMrUoUFeuDzvwvWdNKiikDA8/2+GzGPc0oYrcBM4/XU1TkoQGu
iz28Gti8Q4vBebhyUbUciETgWd8AkcvwJS70s0hkX1jDm7MRP6nN1QfgsXw8hbz5
U8oqZ9AzST0ZTiRdzG3XBeFNVvtCUmtk4qj2OLYpwepf2aWvjtGqN21b0vEJcn6C
1iMguZLsTw6HK2uO+zVwXSNpXB3Y1dT4fwRgRwEgKzAzQR18oVqmcB2l2YjbJOVd
INYmBRgBuvzZZ8N0/YGPLROvMgSL9iAIxtk3WXmG0RlEt0gWueAYTmHkXF5IsYd2
wZIGh47pAUV+F/GLRLH1pa8mpS8eUuBUykeR+HFme14c1OTGuKbk8YrY1qzMbAYk
FR10MB5/4cQXzBTVkEJ5z3qQr0XFR1FYweKN1BsDQDc88gPxGfPwDr3pNzPGh7n2
e4fZetvqB/3+Z+qmPmjZ7ZkCq0DMXkHQ3mgXTNOf90HkQMRkVm5Ru7sxlwu4z7C8
2GVptKt/EFyp50fnvWS0fvdVHAyIgx2NA/EgJsekpHjbRPr2GiMXiBh7e81K7/yv
aYpn8n2CGl7g/isTB1w08aw1fzMWYvWan+Vv9Ew5UofkyfJwEOsc3puumiZQdTff
Z/2qaDu9lEfmnnqwnRB3hJeOVqNjvSheDlUw9xyoPCTa2fKJldQNdyheuZgjOO+n
C4btTAdosLCN7pABCwNU0OJFh9CnY/Iqme31AHlXKJz6Q0EkrOu4ouk3E7rH8ph7
fWacjXKj5Xg03i01EVufGOWfhNZ/Zc1GaKsR9oBLmCwGX7O3GgmO+S8oOu9IxJ7P
5pEYrsh5D7sEW3NhqtktlVAPb896Pd6pKbmDYaoyrHLGskVI98dks2WwPOhW/CG6
ZjglewnNc46d4hhcZrxJ8Q+SHjLzQYJ2bWAVoyUAZgC7Xp+Go5W3rojw3XH0O3vT
NKd4AjaRPHw6tujOh+veAyWhlPRQdvKBZzSXoSqQ1eRKjEJSX07l9Dwxu6uNT/7g
lecM7wBzZOaVTU7ERqesj/LdmqYvcAqgHWojf7VuSCMwYdM142IF5WnjvkvVOEFq
dbyjfU/z8063UMYbA/U+YicjR/28gcb6tLcRqJoftW2vZisEZw6JZAY100em52oS
HMDhJ/GXoiy8xWddgux5bu28x89hwe9CZQYXeONivRJwPFtK6bXV0ZaTnkJm9xTz
KfgWI0Be8KRxfBM5MfVXmKZ8gXMnTI8nykjnt49J/P7vpHS6qO2MoPHuoDuXJ4Ab
8ro7CiIZSFikTEFZ/WpNhrvhMyD5qwH2Cxv+nFqicS+/R7bhi4YjTuz1aU68qfdw
nUfgmP7qIDL9bdq+BvmTaXaWtUqVhZpXDvC0appHvjyVYE4ZszmkqP86xQD3dq3P
p0MFMC1JZslpEYQ7cJWyGBeNyq5NcF/eLo/KG7T2LAAuN0gnXGMQR8OSepNjENME
7HheVIveF9Ng5MrZE34Z3+mdZizRQjKr2UudGM/nVl+JW8td7OP0XBd0gfvqmbC5
o12jCod7WFWJAcw2IrfjuCUF/Qcf4HkKjFvIxESzqaBvk+GVNqW1qs8p7hw7tbAO
emmS3uNwZYywcon9qkEx3HfhbedTLCW6UxapZ/btmrEchEzX+BXkPUSa7Ivzt0x2
ID5FvV6SPrq11fCKrYO51HrWl4CUD0agh6iiyq4T7u0UnidfilMOLq+o2audmCEF
k8fVMHPAecn0OJU840crDJ0O/RpbahxayCAK1MUqGvU5fm9QtEcrp+VTJV1XPdf/
HXQs+PR/t+EOMSoudJwEGdz1bvN1/BX3+f++wiw9Oys7vTCMqowqKqL4Mjm/JDZK
lnVjPyfFMkKY5q2FjzYGxmj8oaPo+PjDgeDzHWf47PPB0SzHO+bFW57IwoDdu5pt
Il02jCxlO0YStaPiYq3zDhO4a13jZXryksTMtDm60Z0BWb15EDl5Cwk5ufOInv5O
ZOF0MjTsD0I13NsNciJmzQWUypNiIRJQpjgNu7yVVzLyUT3jHlvdU3PkV75sylOx
EdUWNnETtK6KUXdrjdPPmQ+uYNWFzKeVGvoNVlgOdWTJjihSYeJufE5rP1/bmzw5
5FNCtCHiHnbDe+r/Z5cWzKVgRWCn7nVc9pudVj/obX/t92hi8OUZtGD7cKF+DDC6
qP5Ub+zYDLp0BD4OxcttEYqN0/9xOgkecIi5Gc1tzrwte2tZ2d7TwYHRgMvc7XTs
R4SVvDBWreIUZSnCgJWy+zmApYYCRYxI7uk9AkoTKgG6cDL83qYCqq4Df3XaJX3G
q5XKS+g7EHo11x3eLOJMaSEZaDsqejpJNRwkht+80DY4xIUxuGylvMR4YAZD3QIl
6/oh+FkvM0V+cijJBsmtALziWbBq615X2F5G2Taca7QeJazrMh3vSJF6Rz+CxTJM
s3+WY2tZi8BldWT92t3nf7wxaNtjWVg4ZqDqCo1SMUqrxQbQkn3MGzwkEIp9ZSFi
U+YSzDtZy7neVykCiEKSBqXDH/kLD83OLZMri4ngO+bIu/Jh1+fZtDAfF5cbVHmz
T2iVQbBGnUrz/tKIwdGRxrVOMBz0NJgmZuqsbvGM0z+XWiaX/M7m0pDjpIkBOtDp
xjYoPtNfcfYwRmrLkqTzC42k5IPk/INrPWegpuRZqypwbQI5iNLwlltTY/ZSQ3W2
BejPbCLlBrVouZWMKYTcwyREabGZpZWJH3oiqvVBNcuNeN3T0uWo+7HL8f6kfdEz
+rEjihGVQ5OMHurSafeH3z5gYqdHhlq88tFHfUDAJVX44DiG5jPoV2u+RvJKdNZl
xf/vTaz9ZNDo8iT5XjVO18oUZAkuE2tfBVEvReWg3hHVvt73X3Cx8I9CLPJXGSQd
sfqIFZ0hOg+zKwBHVUasmORBLpq7vJRVsoBMt530clY69y7jBmF4gTtZov6NGwSB
iJd6MicANzOujRsXiALMmnWMkVCaTffG2rCBQMhZB/Hu50b9TLQ8hs5K8rru9zC1
bhmo7yvk56Ow9tdOqmVJxfQDmbWJmufqbjVuRTz7a1LFKy0/efof0VE2aI5pPq69
d5e8XCF7MLCXWNUFKecPPHFfRchZp7nCdE71/kGPii5HXNGvMSVc3gf2+A6DUOcW
5AYoSANIJ/HCDfLO8HIb99OGbBbv5te3TYJh6nNvmJcojbgHhVuJgRbosJe0ibAn
lxByc7AYvflTDZnDr/WodC9fVKEg4WPJRgZla7U4EBHay/rBI5/4IvOuJThE2RUc
5BZHOzgF+/2fmOO3f4foVHItGEDH4KMpK4uT4bk00E56tSnJQqQm7zorxCrnoC7h
KW94zIDeja57kWuOhppRL0kthPA4tXMePsd/xb8cRdAD6qraYvGieLckkM2uvpYH
PwGd3a2taZuwgQOQChBPatEaYqHuqwBpxPRoef02NVnu+DZDOy24h0SdH7VVJvrR
dB//abPCF3qVBjXFkyNMU5OuDgoW723ANt1hh/NYBUa1GijzCKFhGsDKWNzPeSWd
udAxkc7i0zzcevWNcUwBCnx42Q6yCAAd4C8GLfbsFAgV9XVMsAt+d5lv+ZOlAxw3
rid7mkne2vY82+234dMNzJAxNf+Vc6oHGb6KkDzqbeyzzGYQRGlrcYQlk5qn1tFH
xKDjZgzrY0IF3f13ynxSdy8TBrMx+rn1eA9H1ezAZM8LXpMwCRBsxEAYdFKt28ET
G9sVFfcQo6m9FSjqQKFRf1v5k+Dschko+jjD5/JUblU531b0K7Yl8d/I7emm0KCP
XYk9kidz02OY94zV2tbAHIFakb+MLyDputofYBEHjnvoGAx57nWst7xfuyrysi1f
6kGxER7jjjpwVUa8e0M3F5AFoFJXkRZEjmh+scgo0e7JNjEXxmD62O7Qus0h1nVj
BkHbxpwRNNZewaQ8Alq8S7NVlcdHsQC4H+xgB1h84kDYieLvAviKQE5WPMFJRUzv
gKq9CtDh72au6vRBmddyc89wtDhjmtTEgMt530BSIkhzIX7aJMd0aDEJkoePlf2G
4wOTAoWFe7uv2Hf7LxXirgyZa3Ve9VWJAeZdoUj2e99oUehF2tLEFHzDdz+WNZCb
cjomWfANpguiXvlugDqGbKKH+PiGagNIstuRWLyvT1auublc4npSselznYKLh+kK
jg/FyO7wKxvrAn7j6BTqTLsX6pmZf5a34WTqwcVxVBz8YcQBkRsQTyx80PeXqfpB
IcVU42Y3cRZNbp0TjTiqYl5T/qt7u4TH3Z7E2mXnEK6EOL1kgaw9LONU5Zh7Dyr3
orBona/PUcy3W0rsOmJzzO2Ft47wL9Y0EyXl+njqWs89TlP4DhfzC8Ex5nTMoDi2
4eSmi5tuKwje4HpwHZHhj+XDZ1FmTX07IcBNwmOkqZ4TBTpA1Vd/Xu+ZPruSUPIv
jfCImffOxh+arn1TIf/I24OYbDbT+cBaH+ukcyWUIkwwVWAjqSYICIYXr8mwWbsJ
2plvggjKorcyayjSVGrLRt5rmjyYyY3Y+niWmZR8kiyGFy8wiVsMBbRYMClPNihh
NjipMeDVht/0OOm60y9e6dNcSKS35oPO+eGOKShtCvxrlOlLFTbH+xRH1wMRyjPF
TVuWv7xZBjif0KzAJAXvVYp4aT/vPmIJjLNggwKmo5ayEBbT4JrgCRGs8GpWlf5o
aJmCwxzqplG5TyPOPwL4dI2wUBtRDxGJNn7JuBcgUU/bDdqEE7XOiRCk0NSOiQ80
HQ4oc51PShYjgBv6OLRutbQBctrwIZSi2O4lhDsM9xe4ypBp3vxk56SlM1Jyyu8g
UrFwEW8dNMSdp6vIF4P4QnRa5tBlriGbIZTGB4rqjTuvoJqbzjl31tsQfQHlstmo
bk6fOSJ19uhZlHBERROuWxp4/EJeC0sgk71o8DXd6ND4gLxSN0IryJSGTuhF5T+u
qC/f1hR6p2BfalIUpV6xrzQkUa9xrO5EmISZ1rFfQWpI3h9RFgkU0ov4bbBGA86g
kgA+Bfok3VF7P93tqOuC5p6JSqz2i5AF1UdTZ1OkZGPCG/eJiO9lOqzZlBsBSYVv
noE00fyP8Vvft+61BITjhz1YpZlsLPPzdOpLY9zfQXeRaKi8enBKusW2YXE4I129
24gWVoQL7IdfY8D/5UTgLb7QQXd5iSnb07gXom8U8DwXuQYqvy3kWLeRz1vM5gop
nWTCmG7CuxySOpuiALOwA0Lgx6TyFtyyJeYFf3wMuje4QWc8PbaSFC1xTRQZnuk+
9cA0W1NpZUTlESoiGybTUa452JqPajWYIlRjkhKAxq1B3fUlOJ9JN0aGTULHAYpv
vo9iTT3obOnip5PX6OGW74JLahmpE2IYPtV2ECDAfP7W7qTPEHTbcv27Ot+d9Z4i
HUNRXsxsj11eCUo44HCbOtPRqcSLo2hbmg8H9XeaakOpdxKBVm9lc9IgedhSyS0l
G/XkVC4XobE/recRvkU8ChrMgzy34ORlJlvkR4YMwNbaSs68BeeG1nl7nFYtu0GN
03ESQkgg8bixZNYFz68006DQJnp1Mpt8bzC+PhS10lkUGSoglf1xQ/hF7auApFSC
bTq/B8nDXvx+TSF7LLi7NV4q82modreUXYpjPyhY58wrYUvKF/RX+VHCgzB8gTOw
Aqhk8u24ksbNdv5uWcr3LyJ1r0T/9h7fC50cwZU/S0Wf3r4D3r9TM2yhXMlUZ5I5
YMuQeqlyz/EOagX+GBdEFaoq4mdda/4ChJS6xeTXY1okUx9hPNEp6otgbqJaqyDB
YnzQfu4IuI9LglVPbTwBm0xZBLevNvhxwYEQSFFMM11j+fSGSaEqB0UZpwhHxXPz
dhBfX3DfhondSf+4qnrsUDr3vmg6aylTF2eWh3cVi07j2uM7CJY/GwpjqsDSJAm+
A7nf622iU0L5jIartRe3RQARcbd15K3PGJ/6+L9w2ukVxpH0NvZecuoMX1BwreFW
tki3ktGQWB349sWCv2Zlh8XOvg3sy60NagQPBPTznRjNnpYN/Hw4iF2ENo/hHg4e
uaL13U3JB3I1tnI5gangMGyc+jx67QsFmopcrTR5jGJWMypbc5jqHGRPGIOJpH4X
UFHI04BCtuGhA0hWSXg45dXfZe5hX2AQ5dAry2oADlEuf3au4DOtpkLIWYRk9baK
6D/Dx0zCavAsjpPlUPRh+XNbn9vPvOHIhThN8Lj4TgP2FUVT9TcnL4weVtZlPC8T
lJsMGpFaFVEKKFxFK5GPCHU1ErJD9v+ea6uxI441zyboZCLjGJae/0uix4RFP0BY
oEkamQQNUBy+eQJn15r9SAE13K2WIvnG40TCBn6xQ+xYefTdvqH/PsFyre9xKZ+M
j22sWiwFM00JJWesBiAw73wLftI3NgfBGpxaIWqc4PaDluQeBTXDKrcqz8IX5OCa
vaqZsXWavsWGqC4j2ud6fnO7EcjB4ViIKFMwfEfdf1PHlA+UZ1ZBrC1na1nWJcn1
Bs0lJ0cesWS2e5o6hFEnjAeLojtZA4xHDdipjjDeb1EAV6rBlJsVuJt4Fg2qwSIA
iVPwvrsiLbMlTiltxUbYNGOrLywJhMPH5WxFV6wKH59P6ut/Fb67wtFmfKv5kUKx
buTU4LP6XT3QB5B2dgHAtF/MP643B1eIysJvTD0AuK/MHTXtCnp/iixUk4RxYKQR
PX2QNu/Dym0uoNvgCEvGZqt9qOYEZbVANQp/Wa1EEaikpoGaJUjJMRZy3RT9Yimd
7UoE2qP079BBL3IBDh10lmxEZQk/Vq2/Dd7arKBhwuXTSBJvNc6Ynpe6g4b3j8bo
bMtBBtVHlSbaunkGaHg68leywp950O5VLfO3zMYDeOK+8Zye/TtKkzxB5nZFguT2
gJF/t3Y+bjLhFK2/71q1svij1iWBTitbrRyj1YPeh3NhBz3iBAD0FlRteNckahWw
Q1hkWwg6ZJ/g359XTmoHNa5DN3R13af+T5jkYFlof5NllSicHa0KTv9kmhwQY2bS
pGAwQ4AzmZvoApVg5Tk8261BpEx0X6r6K1PP/NFu9adJ7Bm65nvCTiV4FwTK6sDQ
uk2z9vwEeI/MvaVsgbunqK0SyYIaCvaxuzmHW/Od1ChVUN7pV7jRJvCILehWWwA7
nk84B5FNteiDZx+dGSXMoWaU2c7HRF3c0V5I5Q3hhSDcbNdqAnwyWs1/rNsY8uI2
b1MPH/2//PUsyl7KgfSJ9Mn9PYA1g0V93cGaLGuS8QrtGQsVHNGeZIcxodSSyqVb
1qrLQMAo/IqO55D79igfhEQurzZmuHtElQ9ea4V0+u41eHxtDSsSMmStFG84Wts6
3XOX3fx5ZjiW0fUFQ6IB1gOF5DTfS9WIY06t6jm8X5GD9gRKpqKKxxEd5aYFMCqS
fHgFnuKcEcBDEAyo3/sXQkrIy9yd0fg44Njm/+RWJBcI0wEcWEf7DLwY4mZAcJp+
B6tSDDk12itaTsqEEwVJ/owR0x8VeWnAxTi+9uTT+A3yQf4mtLQmAflJdRl0Xx+x
jby9HfCY87++2SzVExYzTfqhDFKqQvK2oiZ4Ug++vNNK8INSWwt+WmyEgRRlhD0/
yq5CzPVRgGaBRh7RjPCFfBQlmQPssSQi8xduKNbUPvgokh9DoCoe7f6T7FI8zetG
3BFNB5RaKXTohG217awcam7Vn7Jml7WMizLJbb0yvwQtUkKIb9ngqnQh7WWuu9fA
iSty/55tosy6jAZAlZRQXp/y4JkempDkQgpU65HI6c6ZSE1T+F6Rl+KuWjqsg0Xw
U7xNYOF9vpcfoOFtdSy+m/ccOD9phXRsurZAe/buJ20WrgbIJX3JYb09LMrBVadH
CkMQnNSvm/H3jYXO2oy5Pj2yP98ti3FQAb9RcLbm8EA3SMYqp7E8HwTr2x3+hfm6
vkspYCv+YVvpGsownxlfQE4/fWv0On6KqxrUUzIjXreUZBYlMYHRNZEl4X7Lzf1E
3Kjpy5SnjOZJGNWaXGl8MjbXDDTp2dDbG74F7DxvvQ1SRQsFRSSvMHVv1iXWBya1
ndN71JZ4dD+/4Fdh9+XVNb/0Rt2t4BcEvh70wVJwzSQj/pc2OcaH6amqX8saLHjc
GSQlT6RDVNmxfhl0MzvqnVvoD1ZvRSN9X7QEzAtezJOBNankZtDJVOtyX86B18cV
+rBNi/yz/FtFCdUVwlVxexsFGo+LnjszJWgIuRQB0tXE4yx99Uqo2vKS1KpsGOr7
wgIuSgav2ahY/i8Tg0YcXyZtF95EFc/3gFRfwtvAnNi1v6ByPctL9RuM4UGNSvK1
nIS6nar4ik+EMM6tUyUoVWYlqHTn39RsNsrJoIZd7KmCrwFkEROLSRiSYG3RUHFt
BB7pX7yf6Vem+V3bhwbKIWCovfvTUIKBJklAYBl2T3TMblMm/r6u0RcEYr/XT4vf
Pl7vAQ9ORXooabl0anzAf+S8T8nOw/VgA5RKALjRYz84ExrHceZg57buTEQM4wCi
9RH/s2tAlC2ja9VbzdDrHs9Oxaqs56v4714JhUy/fM3WgXrFeH6EOoGCf7lyQpYc
CyOmqjUAcLVpBYUjamg7x83Kz+WIO7ew9rVeE+XNGyWmV3n+zPHeSuAaMCkjHZ/0
5AK7XHZuLrWZnopXztY6L/1lHeJzUmcPvi6F9zIxcrS2yQqhZXnJ0KO+2HMU8JS/
aFaobZiV/NDrNLXu9aiTo+TE3A7EDabXQc8PtNPSgfPqK68rFyTZVYwfv8WOM1v6
QaNA8IMP0bm5MVRzRlwwkYxYOx0/ZvFQTR+STr26B0I63YmNARxhcWFZVF/ldRnU
7fp0XxROoDdrRhuqKCbear5D8aM+deLpu8PR6EutFlNqUXLwuz+7c6hq4fIVxrN3
bunM1yjjuapZL/O9smqaFbd2r1BGucF6lQSKdpg24zY8zLcSCeZrie8UFXYpQT6S
SITN6owkhFH7aJjVc8HnzKp7lTLC57LJRQCOo3INRPEdq4vFYfgkeS3dctnaUckz
oVsECOctsw7czN6zSXzkopWih+gRRK73x81dKkW0VwpPOqE5Eixohxa35kPR3Sc6
fdgqEfkIyI5cixnhyWpObbiIM6J1slrBgiZQgEElVfb3Vfg7zMtsTPts07cnZw/B
ctBOFxC+4Dxs3G659RjlOIOEB4gAxPVnr7VOMDjyoG+/AbZ31QqV8LcxYob3qAXP
41Rr2FgHqczU5UdvLOcSePPr/w/V/Ub7OgsL2LvQsgMNejTvuCUs8ZNcyj6hv5KF
YlCwincS6Kk8+qYQoVQdoL0IRbbSuj7eDfwjQBCnmjgLf2/ksQ7zd4D/vhrl5HgW
zUEglwUGooGlLGleDyzp6NAIOZJK5JD2Pc1HwG1zHLH7ge0OOkTYHnvyzxKvRVGr
As7WUTCjSJAgJF3NqtJyabHPT5AMf1SN5x+K+oN6QFFVoJNvJCGXVMwp3RnaNuGx
uIYKqTYsYFsDSXoA/kA4bNch4sPMkIiUaUFBMXhl7kRjGbAFKlMkhLGgT49LBZ2c
ZWJ/P/SU3wL6mZLZK11Su8IVG/pNlOn9D25bmGCkmxVPl7NVc5DeWh7Kno18pG+H
71iYiMulnBxjTMJjzWrVeNO31Yl/NctooRgFSpIZXLG6Hc2iW0WpRjylhN2E36mz
bEyombIKBb6AzFmHl6YTsRn9ieMJ5o/6A1F0vGjhBafwm7GuXbNn/VWxoubWEZ36
g2/8iZRuFU2XII0M8E7C6SnlwvVjqeu1zw0IpfU4yMFipC6ExPgehmm05a2RRYJa
HKkhPRyvDpFH3/D68MmJePR8MfEejGQAG1lYzxeejYf4Lmr2glbwJbBwS2VTf1tF
4fAInsBjDPR0JYXNb3gklXU8i3yj+00sZXjqG25urELa9XLEW4A7NuBJwJczCi0w
6DoPqYrt7eV6T5BF7ISFXbfwEEV67PvPCVbAOwHP8c49J2ps6FVzRENf/O4hGJHJ
n6ab7cYPwXCl3VGgbyOWySewUTp3yaWTEa3EiaU7KLUSZDpZ25ZKndyYwDZe3tAD
Z/8R1SOpkKvJ8oc4zXRBATv7ZTo9Kd4rRhjTyrtUL/bEli1zGQ/HUSfotnwtbUZi
KQgOPlQpW+8C2EQPH8DOYKiIE4R7LE6i4CXB7JwOO22bNqfdWkDDqNXyisTeTn+P
mzs96DB/l6nIC+frnUhT0YVf9ago8lMrzO8FNQvuc+wI3hKiRyiQQ2SLt2nxS+Ei
LEN+AohlD0Ex25xEhBj9KYz03MVrAQjTW5FtW9eLJDyd4ib0V/5rLnMmXU9Y6SzE
SbraEbmXXoGY9008Nc/UzgxBagRsnoyZvf1CU/gC5oSwP8BVmQz289x6giQIsWxp
5Jn3vCkdBxaRQNCti/4GM2m8KjhWyDV0U/lPjpIOjKMRWUWdk5hp3ByIpvjLHybx
fXgEPh7MK+acjaW+5aEqBFyopQ5MWQtE0ORnE3R6Xvt0Umfmh10Hcu0xuSVIoQmP
adhhM6/6eMgsOAWqucXpGXl6McIiH7nkCsZDPqAygw+aFs9krsSi1OwYtP0EU0PH
48i2U3lUgLBcd9l4/1eZCJqZHj1JTlsEPHPeFtjgviYksRAGtRCbrYqvE9I85jWE
LmtGKK1GjbxOYW4XQeyFF3A0lmsm7JfgayupkIIpCNsW5KkbIoFzX+fGWEteWaxj
kLonEnah3gBBVzSRJzcvxpQbVL8BX2FgS3x1NckT1PeyqIxQgDeuYeSN73JYlUpA
d+fDGBmLuKUgb2u3TV3bwkmrO18R34UZNNQpbZiCy4J8//3uko5bMevStrFCLXTC
/crA6jt2zJhv4xUMmtZYLqskjqqI0cGa/zkl7mxqxNrqeS51AK2/bjPUrACGyvub
8KVAdRWZRAT3ua1zjO9WwUjaSAh77qKzMV25HDF8BMq8osZ/C432KMCJhLf4dqmd
glxA5vR8W1Asw3E5KZWyx2HJwpeOSwuifKP1bft0DiCMjsXq43JjLur5TE6PjIib
BjUk8uvTpP5Jmf9Ze6R0ldpY2nWE9E78nBNY/2zJAXa7swfmyXFgyJ7Riz2+DUn5
Uf5zI92K0UbHZ95TQqqWk5Squbmh7Vr2s2hQErv2tJpBR1TBjmC6pJ785DsEBS6z
S/BgkBdPH5SNAFT4G44Dtr3K3yS1yfbspxIJTOibwLa73PBv4QFT+tSnkPajZA4f
INUpkWWyZaLyRzF3MkT8vXBLQOkKUFLdjzVPEoKQuXx+J1P0E6zbgP/OEnVWNSsK
Kbo2UOwTu7V0+O61FakBIsTsQzonue8YxmryEdumbzDGqhX5m8W1pdRBeYNn7rNm
tDg0/CR7rzogOiU/jWnhk/owu60QaobaB6Ue3mMHx6KmsTurcJjmvm1tX2VCvJlU
DDqZrBQqCJxTvFmzlhvb4VzqAY+HS4WOhKqzPaeBuOZq1I+1G4nfwsKMb46b4O5j
KmkeLzAOC+mcK6JS7oxUsv7RshF/N0DwH0+r5RuQROChCAR7C7kMeqSs6gl5IWex
j1/wHCVrOIHJJ6n6qqAYn2HZWB8wjIpB0JGPoS2pvc5nP4u5ytQRy1wEGyG7FHaE
HsL3HWI5YMbPQwm+itdGqMMufAXeqh1haju3yJrhmPqRWVET8LAfjCoPjWg7xg+L
Mwz9Kjx7htdTtRoA1XRmuxGtFmlXtfUGx1RXwUP2wF8xPDEE5T8UqeUCrMCYtp0e
/3bdy/yvdUQZOi+TLq3MlkJcc/bWJjwEOON4Ke8VSMKnyfDU4I6trOENldzLcTJl
lw0MquYBuVlsdNuCD/n5WqhuNmcOAVspHh68F28APsF+bkwziY+Tmej6pEUEFOwU
gGpwjKlzBgaMDGnpAJBGP5ZF9m9pYovsFXWVjkSkTvuJjQaWnrSQVwDUpViisqJb
NYThh77iz0rHm/o5a3ONEmmV7liVp3lFuZXRA8EYxEZHRPYbzb6wstI+ZXEK55ro
6Huh5hKd153fdReIhxCCY7gl7tlLnurictcG0TmWRiWz46tB3rGp51EYmIgD7moZ
lToVcw+zEM4Dh0IP6wmhd2rdL41vWsPln60tN6RUaNwo6KmtkFNpLgGYL803vABW
MoaJY1UxmIfn5WQNRrVIAxmdCobIuGCRwNNhpnlI7ZPQVvqUKV9/TxKaCONfMwMs
MfNhdJS183GzPUgomRIKtrHaGlg94KyHiPOTxzVhyEC2a86gIrgeHS9des9h2RHv
LnY3hg1/6WzbOTxFgJTBA+JD4eZMyjFY2w2t69DDjEJTALPPPX7MvTlreGzwFiXi
aw1h2A4cnZ4ubwca4cFECr8YadvEQf0Ftc3sIETresy3rV+TtEaMQegPNuZDJ6Ge
cSJeu2himp94q1u4tG6TqitGtr6etlevLAnRwpruoLYnSgkMVkDkhwocreAU6+l5
btyWXt+xQCyLS1WYUsU+mGYewrAHO4KQutwSMeKPmvRqMHuhhweg5Nb6yJNB3c0v
v2iPHgPYwuTYGNycTAVJUQfTMgqNRnMYoYxGONzvJnOORzSNhPGtyKIeK0Vt1fk+
j+WQBC8FxEuF3vAVk9zNsxlPQIimUBNvN5W4Nt09rbIlNWASrMb6YEcvv7ss1UdP
TQ9kIKST/zMKEpttyjePC428KXLtp3LoGgl/XGj4nFveb/cI+F+BRYK4m4VzbmdM
MjzflPpyLIEC2Yoa+Q7wPFdJoXbnfmi7Vjn5DCHz8do6+RffAltmtCIsXmxc3MhW
Jtv7Euvqgrr0uM62BVaR3GU+ZlOJ6hFZXsGbJTz4NtrS7UruzIBZfoUiCx2NTISD
sXomdjcJeecK0h4it7EMKtD6x9kKejsiLD4aozQeFN1foMXIoEfG+Nm5coOnyAGI
0w669J45fsRIhv3VkYQ5UdqclYn4mUsaaMVEXt1ms0qHreAQdiIkl3lUiMuLSQpI
Nj7TP5uTlAt7XPor6wBvJsUL5jOfCtFy5AWCI8iocEMxCuiWhHvxVGBp73BC5sN0
W+cSd/HSuEOal6OGT+G/cLZ55yb5MPWjfh5qX9IDH0o777olgby2SuwM4O9Rcu/8
J7XAtGLNkTH38vzPmnBJNVrnb7F1rUkRq2LFxYChBfqO/51IeRkVhuP4PiYTSd0/
5K4iUjjf4Ik3LhWXpKFy/MReI5SmUIhZd5CGCxwTtVji6FhtcT8oqCB0duhSTO6a
1XiO4O+qIVwBT9AoH6Zm+6AZDBaF5W6KBB7Kxi3/aeCkXZaqnxeqnys/vnLCqb4t
EIGN+3BAScZfm/S1q2ad7WX0tp91hAGcEkrjTcGCPbtkCyjUcJ+hCt6l/qzqCkVk
pgSP3vOrJgxHWVTULZ209LNcqKvx9W782radYxxwV+gw2pVg7xYu6yetAIQbna3d
OmQvavvCVDVB3wvyly8CgOxiiVW8C0khkdlqeIKUCf0FMQa8lUk3JGnaqc7WDSK8
tD63Ce1CBjPB9JSPbMPGHGfr4zTyCiNuzgzhwJOvmww5/9wjdTWs9z9QUFmdmfoJ
Bfaywm3LTKG5jje8VdXyxNbwtaap8FQpJoABiMa9u/dVWTnJNFc2VwVhn53rfJjg
v40zV+MeI0o8KrrbQIA7F4dj6RdnpJoVxyze2nuerl5RnRkRVTD1j3iBD2Y/cLVB
njST+9dhOj7ObepmnqEXP0ccws9ZgTrn3OiTTPli23nThP/lPVDoeIY87gjope5f
iUYixXIO+kv/hRqO/rrNwflkT6KNXK7pKV2XspDOxryzVVLhYh0rdBd5L8uFIHa2
uSjSSI415G4aIOD7BUJ1iOfI5luv9496VEkwy26nlHPe1eNCVIoNPU3t84Xf/mNt
4PmoxaFI9/bBxIlRxYrVjA1rLgQ+/HqZe+W6FRb6iIO/CXQW6LsA+SO7ANXtG8sP
fcoZKwZe+wgNoSXBkYjS3pB/+A1DY3s2YdeEIaJblWBnhgAAkKSUL6Vqk716ZzE+
ThXAhnxe1ESIOJMzE3gEPsvELWLVd5bcB3mzr10vqukwv+kvjni5B7SzIGLB6miF
KwPmN7V3nBGBFB3COiDCsGoyg/pOW1ZvsWRBJWPXNQO3if5Js/URuLXLkox+tEFw
gi3dZpL5baXpcCvofPSQhAZN57R5uY5sUgQBRuFRk2hrOTmmJmHkM4s0eQ31M9Fd
YmvrAHK5Pi2oEmO7sEda04Xw3eJ04bswX/uL2iIS5PKHA9g/ozuqYxdhsABahju3
SON/j89v+hxER1ln8iwoq1C5DQJLfkjeq5lBGpvCpbXEt9ROggNymKIYoDCV3i9/
xeBCtu1gGPFR0upYysXaACe35kILwF4pYd0F2cG2nGimoUI4Lhax2vXfonvo+fz9
iDrUimmnoBEC1wPkGNvr752VVgwEWxqlW+XAJuq4kxbo3LghcqIDnmyO41EcaMLn
TD4MHfyjs7/DPbt1CoZes6x5IjdqsmEI4z42eL5p1OOETNxIzFRAkIaBoWqnWfHY
jkKxWOzHyw4ZACvtAI+TuClPguldH3LRYPVAeal3pyasheHhpY5X5YN5pEuYf5t8
FVAvqUYBfOjp+HLtHEEGCFJxFTUMiQsBsZ043i9G3UdgVBHTFSrGYvvfK9UWMt5m
nDY/lSTNwYZOiaVT+DNpT3cB6BeJvnZ7ZJdS3GfznT2Ij1mJjrThm7NUAQGzKM8Q
6FjHOOaM5lBEX/3E/ZnIjG+RuzbVuArSZ3WeH2XoIDvsos0zBWhxM2bMSWO3Wy8Y
hwJ5gTIU9SU6E39+HvbsBJyvd5GwZ0rQtL/dbXS1q3MGJLrDZcmQD4q/0xKzhcnm
t6T91JmujdD22SCCl7kInUZf3ROMjIYfjU3v1p+zEgYucoXDrJZGFyr8xRMYMQre
WiKwzuX+IXbXt2UHXcqQ6jUnVU+ejBbCLVQo8DwCQ0R7Ne+JHZWYQmosIQRihs5p
otcmEie7lORK3/bjbrkhKEDUZNm08xi+bESilQ0fT5AthY2LmltEiSURItmHf/7K
SmHw90WUZOY9oBNr3ktz6KFjqaao38lrFlBmCFCs1m19n2YeqN/FnhUAP1oGJxHb
jCedoSL3Oep8dKo6HBSAQfYoxyM9Lz/G0/puYgb11iDapVkl+tMRHcqUcJ5C1ZRs
6Q0HgNapF+LQ1NsPhvfJfngZAqkPfC/m8EjZZyACAA5odRq6tKOY+h8uX9+C2R5j
ZUe09dw60M1N6+LDO1RDBALm6lbIC5aD8T5QMt5o5yEK5UCAQ35nestdNwXHtkIu
NHxj7hGOMmqDTV28gNV/zO41k5c+jUJJoPwI/NeTD8gmsg61M9EAPaKDsL18Z9Gm
97d7ja4OeKIFBYs1WEjm4ARA/p1WdjXMm1GDAgvO2R35s0GkBRXS9l4U29mGD3cQ
E4gQD/y59F8c/+Uu/djdPWxsiVS5lQWC8nPiVNG7FGsJStQGb2E5CAi7LHbnwEpG
h9AHa8CWW6261QERJatI9IXwDM1MSPK4QXIgKBB++/N40FG3vk1C1NT3VG1FXPYS
ya5+7Eiq6ITxNmQb66ymbiBAJK9Jn1Z97fR0c+8Ul3ruZrV6bSxoXJ3muXWvblYW
XGn5qNb8k4EBrs4MX+T/+EmP2fS3UiUcPz3pIsX9hDAewFVgXqT9RBQDBJchUVqD
tRWdFXcIrNFSEaN8+uW5+eZhNL6NtdCMIHDe0mQt9198HmFqX5jS10YHFDf2w/5k
TUr9Mx/OE+hwacrOrxHy4zRGvUh80vD3iMl/UUVrQOAEnKxOyRwZDOp30uW68JN7
ZcOHpHdiP+Z7ej0pRFmbDsi1vZikgP3JfQYz9hIhUkc6x1T9FAljB+O2skviTP3Q
4tmMTYiOy8G4N0bkcxN1GiyoFzQlpfchNoR9fZ63GNB4NAKXrGo2v0JzcIVp0mQ8
LJiqBXbT47FG8zv5cNR48ekUH5dsJ2hO0FHdNM0QQiNJeDpLXJKyKDdfC6pl/rr4
qQz8Og8ZbrnYp4U262gO/x1207MYarfVUlbUWD/ur6QlNknsM9GX/48RloCnA2BS
TsGqWEiAw9FMcdRIQ3K71wq1eN21f403/M7qT2Rdcbfv7FHUWatrxGPqhHhUS5N0
nA1cejkcpCdghR8+7dX3Qev1VN/qxGxzCY3HbwDln7KS2bQiNthSa6LAXu8yNSUj
eSPDGqD18SS7w9h8HlDUg4skoJu9m5fnIuf4y8mWR13yRSqx/Fb1sNPbECrx2TOo
2qtilOWVB5gMIMMqovCeJe1veUWxY8YURX22LkOUKiiLve26Z9VPYZPgVFXbS7HT
Zt3sXBDSor7dPm+E0nxdO4N2Rh9UmMPyR8tWA79sj5ohgbxt/BcMZ75mgn3ddDqT
q22QiUuKGpBDhtxqqD6nL3M6QV1+Rc5LwVR7en+ECO9j4MRtJgnrYuYHOBX5ha4v
oh3sAf1rfcJNJHdCY7yrUDEonN3I8j89XIuwClymyQiWqiH5l8gEaWbru6d8ZWqJ
Sg5sjWQ+WmbQ/1PcnmG79jXslubG+FaVJzfMWbClwXtsEoW/Z/7AZLG5ca23suWq
l+1oIrvEmbU0hdTVCPY17nj7oQ92HFzmBtgNnpGThhUiEC7dX9N91pLOOkIMfZh8
sWaLSnbBEKEFg2mwh8mcuZyVhpDK1O5bKw+3PXplpo4V+FNt42w+jzCgDo3lVZbw
PnAy4a81OVdqH1X2QuOsBUoEaQjatTlJ4eELgfB50X9mjdV6/6bueMjuTv5VyI3F
zpp8GlK31S6bJiW8CoNoBnhNX8PcBoOcNTVnJe7iUgQ5ThO6mmlfF2x1eFOw5EjA
OSWwxBGwv7kgOw7rPuoHUe6VY598AKiPEdrBnEVkHzk1ZGeie6SLS3UjZiw6jhUD
4nruL1OYOq6NZfJ/R5tNvKv2bRDgR5Qr9GTslPJmjamrF3hdw6Bjbt+XNkVfX34O
HavwV/Ksg1Q8sWMsQ+B37//WDEsY8WfwCYPKG6s3uzfS4BfAWCDGNllQM3Kx1C8v
lzwjdheiL9EMY5eKeowj0mYd5fJQ/sZ6d0HUmNgGKe8+4UUAhULsN9uGxWTftss+
wIRZ4eEkZ1gHwq8t4688O9qOEeGr2lLK4ZJDAEy2cPdpkPXw5zfnqe5Ztz/JUeui
CYQ5GUgMru1QXFq5jlr7vh8TRCId0A1LkCz9Kn+irmo7UkEHxysrj2friCNRDmzj
DTVMhvkOmN4JS1lYJBbAeM3IwcbXZDOmulKMaujpteeINj1ZOK11t2YOPqhQlLeo
7M/oJOzUti0NTepZQKfFbOdaRL+yPeQQzaTK+y7PyFT1QpsbG5/EmP08dEi+7p5e
h6odhfJGdQEN0lS/jCuF6+W6xwYDmR0sRpPAL/C1Vtt+zvGZJiTLmh+9nuAK07IG
4KUGeLUnt9v7EYo5SVIDC8P06ygZB0yfh8V06rP4qEtkVnZsOt7kdh8LDT/2E9Ya
juYS/oZPxQ+O0FYOHXcdHOuRfBsZ2ZjW/yBNxKpKOYToaGnxYzOA8YQtJuLsjfNW
uybZcoljmNODwN4jdv692J2ohH1jbKCzpd39HlinqEG1/AYJu6psjC1vsvgXpiB8
cz2Z+0fg5SvXpIJmlbs5ZoNWI/DU+rQQqKrqD2NTupJNincFCGjq9D0V/8hQ6POD
LNpSXeVE2UiK/ruDEDuY2yfSe3SDOR5WWagyrJUifTJDfLbjf9Ivu1zACRiB4LZh
VrK17a/r/tZq3vSJRHi6BX44AFuVElBP5NK/jAOl6UcdUCEwjUqLNfQx/T3LKLd/
APJbi7XYZXkFwZjXp/dk1WVN6taUY8SD9pxgI8FfRYwBuqnd1DUCpJdI4obj2k4K
faAOHceDe9dzdXLmMQtnH1Z0mhrFfLMKcKo3rqO50xJdcMOhsH0Zpbh/1zOcaLwc
5HFaQjOX8MNmuvs+xfJuC9x1E9jbdAwnyc2Ozy6gn/aZiUYJsF1P558FKYBqu5RQ
5ZtwQ52irN0mORFtVXl2Rv7ArQmeczblC0KZZGllx48jkW1ylVCs5X2W+ZylJIrE
K4v1kshCWZhrPWM8Vdym9x0ftRuOlW6zT6Qo4GNyyhmdML/aAQEJ20nfMMDZ+hdK
VdlYMjmKwSLXW0Yd/zq5SQv4kDyEqUsdaR1ZucRy3Ye5mZW+6EBfthG/YicGeWZj
uo8V/KxR+zY2KAPA/pqy8d3u899H041Tq1tYYljiZb9WOswcuxCjJdmC9VGJktF6
7hZdTZk88dMClWjAm0joWPCcWOYKnafcTx3Bu+rNXZIPQRKyMbfYRWbo4cw8pijq
9+Tq6voEZwLr54GPWt/kTs2KlE02ehoIwGAlvAUfvyP58JYTOS9gjq6aiouWyRUQ
+f40/ULkvEKJyhHM7QCkQtTTcC2vwSWRjSox+PXaRJihGEtu6lIqH/LeL1xTQEv4
i2TEbRbkQi9y1195fL5vDdXQy+yLEvMZ2rH7tTQnP9/jZkq0UM7I2KYbBOkVOwSe
hKSkPkt2iv5bdBIxnMmljbPEi+QjXqr5L0DFuZoa/8+qVqFlSsbWCG4NG2qiGIf9
YqabYYkGofmlkpD6ehCyt0UcuOM7phmkHbdZCS5gymXV+4BNXtLIodbSOZtX31gl
kenREZxjQcLksCdTfolnhf6siCbk/v+IX9161FxqUW7ZzoSfzggRWHFXgxWT2SWa
hXPkPFJR+1oP07I991Q9jZ4hghVUZEIrNkw0hg2u03maCqgbPh4to8XlgFiPeuOJ
I5LMftN56WpGs9uMHqSVrAFhsi0DntYAJkq/g4W9/2iR4WEM7t3mpwMcmg9f5KAF
zMBp3ICR9sWjmEHzuQXc35WIqV1r15YH42tf2atrLSBUJlZjGjf/Qrxz3HQBRl2E
f+w72F6yaiKLfyYBko2Q7KoyicrAUJu7x1WuhWCahKkFK5DvoKxnvLE8vZswECYd
Al5ILrOgZhF+NtO1EGP7LGajd2XevB6/Fhfq1TNZ/7o0Etofk0x/thzP1D4CgXJv
aKLCNGerCUeiSnViPAbq7T1XQitMvM4tkzMyYm9c+QrD6C1FT0AddcCQW7BxGRax
PUPo2ZRuPKlHvlJnhJ8LePdom6bsqlh88wyBq7G4JwDtCOYJx34HmqT0ESGOSKoC
6DaG52NcIqQXs4gCILpb2NRIQAgAMf6tffNqH8Wtg/iAaTNVM2pdq5XuKFKP6g6U
V85HSVMk/7gV6mPjJBl3EihiXgldjOgUPewyWIio9ytCTjtIfmvcyi9N1CWdug8V
VNLqMkFYVCsCAL6z/HjJYYfLC7TUu+8X17tT58+Ffw0/DAMY+a9gZoUTtptLJlHz
0iZ90sbI6oBBrPq4Vs9JYpk1d9lfIPpTNcu0Fd8nOX72foIctcgxNOzkwyDxLDOs
QpXAtD9Gpn9uMZNQD9gj/HyvkugXsjF/sDac7mkL/iOYg0hQW56/Q4Vl8UUVZgr+
1ra6tS8nDAAKCztPbc9gAcE2a9ND4hkDTTml/fO9qimoZ1nQmVzCHFV3gNhhE1b0
SDCU+LXn7lGrtTa6NLHlus38aG1CO6RBe5e93M9vUG2vR1R5JGRB0e96KVek0Yqi
iyz0/6Q5J+M4t1kEmsDoZDZdllGcuTAjHw9UpUMWssx9DBRrSzTDE0APL5Ry6m85
JqGMxH6Wnaa0A5PmgwP0Qb7CGhkKGH8DBQBebn9s4nMrOVdj2C5cmwdXnc0bgsOP
6sJznVYTECPB39F5HJbNDeb0K6kvbrazeysynBRkELVxQux4Jml4p+Hc7VMOkKLp
ooeJdr1+i9orp5RU/3v5OY1UoYPkqO8oz/VfiURNO2G+IggDfwfGBXTFbv8HB826
cAMhvk3nqk8gUIRvW9Zb1icBFtr7FWxn6YAJELYE8/vdh662thtSH3yvevIf6ySl
mjO9f93PbiX6opvUu5fWL4RTRPBiDdaYL4wppG2o9pV+3IXQO8wMy1CZHg6VXw3s
iDsFqqbslJamq3k6kgYquqhLIzyICGJTY7rnNrUACTZ4np4y2O4y3Mv7ZpZBth1U
DOuhJOPxIyBg6mD9azaqpnDPR12UpY0f8SJtZ/P4WOpOTqMKwv1J4dbgEzIMqdtJ
p3hlL/5ywYxtx3Zb7RcNHAlglTjmw2Tfx1YKrr1/EzO0R263FVr5cczSkexH7ljg
YoKdnqbuobHd8lBJERkEaOfATKIYmeWWZ444DCkWu0iObjr/nrwwj5yUO0dfrDLY
lQZ5pCjV7XWy5iu6AXJlsFYok/GtzBOd7z4yLUatpzwjd5qda8ArXwQ2vSBl9PDj
bjp71kmbyH4Ktdd/vh9GZkRsIl2e0ZWiX2xufii/qrSMmub6OhcAz/B0jnK7DDNy
VecZ9xKVxwUYCflzYpYP9DysofZXXgnlKfyljWW1pAgsbaP82DKA84LtwwbhE7LQ
zyCYqB5w4PkP9fMRCeHMuf29W87R0eIFibjmWoJFFpnO17Ufc0lua58YfjvxYNfS
4ba8qzHfh1a2xR5n72bfk5ZSAViHz6aWVGKlkssh8p/mLz5v4P3D++VusvDNVAMJ
6ES87AtdI8ZZt+tAdoIBRx3Lz3gB6Hj4wPGPmXcNFAAR36uALam0RCGodmTv/Kge
5552SnZTUyJe7aB4cIzcI0I8CWuRGAJWcVG/9785C1bfCs/M8CwUijtw3jO5/v5Q
3E4y799+KZwcXFt6XdrBvBlGJAo5Txt6rfiO+RHiGHLDt/xmoFdURb13Oxo/+OUc
e/9041A5YlwUXv29bvGjlmQ0zJimFgA8vxwxbReBATSJH0AoJPbjpx6qibtpzHLW
EpRZPRBeX5v5LkqdPbUuLn7FjQFIgRAorZZBEzUjZoo93hN1GP4tS5SQDaXzCMJu
zhGSKaYN+JBFGm7guelFxRNTjktzQKP75oNTiyc4A5v3nYdE+gkS/2xAV1q07kPA
xkQaox3JofwD72esUNIvw5y3PZdn0ImLfwxaBHKn08ns6C+ReSyAqcDZk7E4iR8n
WD8mm5jdI6I6tFfDFN/GLPFK/Cu3BHsJdNyisVcXVt8bHcWtL1C9aoog98JQukjW
LSA0jwmM+TWYb1afteCnyCMi4WpH+CQkoF42JOU6TEblVu4xeRH1brZxAdFXa38P
pqZu9AgkFtgNjhp/gKfMxpjYA4M9pkWx/YjGjd8U+Mbh/gmCQJ0U5p0ccG+H8NkP
QZ4hdASjK3AZBPTfzIkFbgwxLrBd/LDIlyBrrPJb1bH5Y25p+rOtFFN2amfXAGM2
nge+oU6RhMLMZiBP92KIQf2W+IdP4AygLM1PzuM5s0+PaaE32cwZc/Vr5fq804su
eyXHQIcLV1wdpoQPCNZoYS9GuTdvAUfSaXvS0C1ZdcvoKXp3TcNDOCWJfNOg90cr
5bDt5F1lzVOolGfMjiPz+JP71vLCllxGhjpFn3WdEHTvxOVheEi42nA7Leo+XWVC
KngywOxPTGcWNYEm2UgvxaqBjq/JxbQFhqdZxGvqpBcceIQYJseLpYl7eKhFcKkW
inIkRiV9jLJi3DVvpx3HaRRoaRrFxXZb44erw+HZDebsn/hK/fwLtFBs8ctYMCjQ
gGFJ1K9sqS+KDiaVwDos4y8zIgoycDOvZUu8cRo6n0PqeQ0xXVtEcw2MQCnL6GNS
N+Pq3+t+5OLUCkpbjKaVY/M6gMTcARCGy5DksPJ7mfvdjbKC/IQ5/eXeJJF0xBgs
esQpSfEW+fQtHbj5y+aOMmHhyJBY+hu6iIxi/48Ux8A8fO39UzDVt30hq7ssD5V8
3IiTBaVf0rYivJS27gw/bBWONAIREhMH5zwRwjZsBK8mm6dAlZkPYenZcHahFWSn
OmULGqI3dloFm6w7MkCRRlmGFFBcW70fue0xr2BG5m5sxrrUbGW5rT0LOaTF6cch
svq+Lkk/jnF7wUEwzuMYt986wWGGM+Yj1bLVDjI762Upd5WKgMbxbF+4nL0Ga9DV
GkUC2HWITyYalSKUnbwD6LQ6aiQIrbulpid92FUFBOy7F1i2+Iv3wPLs20fyGmPj
/mY+rRNavsVyVQZoLCVzZSpGIDcQPpmdPsw9A2kvC85Ej+xNhtaX4R/wQxlTo/dg
kAusV+yPwQnByqsSjP9vR8E/izslw9CURmf6Vr9robZ/VD4dN84y0lwLUuMntPQT
2BP+2jRl3I2N8gunmxVnwfNsatKZ0s8IJa0nNwjT15VXWosL/OD+OQyHWRujY3yP
9AeI7a6RzjSsUWFDqvIH2eW/H5jr/8DDklfcYQKUIZ1z2AgyTHVFXUGId4jnR1Mp
SWxPo30Zcd/TKledp1YlM6MlhV2+6POkWW4IVDiLJ0D8wUtLwhrwd4mtndWXqZOC
zcMv2W3DnpbFWskWWGDEYCWjFEcogxJ+bhHldqTeMQYYdXuNCqVCilKKjUPaMPjA
0jGI3oMl3UFs2tUz8b/w9/Szec2jGJyy7qS0hiiu7svTygrmtt6toLp/CY2LvR7j
dP72R9lpL+jFjvukIDR8L4xa07+3R2qW0FTZkQZa/ArNFBsr20Pqz8CTrw2nS/p4
LlC8Mq0/Ymv+A/m2F2T95v19VIp5DtM7o1T4KjDLHB+7tiQVO7WYnDOGMRN+qHbP
Ey9qllKAYeLJSDyN7uT79J2+80qEIFOIstfHdHbZUt3/mPw+tUUF1oZ1pKxNdpVU
kkAIZnr7yGnrzzfyETwtMBLQEKYDtZ4obfW4SGhRnZPeit/60FrKAzwjcyUbHlYf
hk8gGH5vTfwbyoVCRpro+Wp8/Ygh/um9EmwpH35YQ0IUZpfoNO/JXfLCj8dt9fTD
hvZSlpCBPlZDdV/zF9aMDhNP4yZfGk8vuhuvgAXGu2MAs58YN6NwPtZXDw0RZS1F
y1rTc2Gkg53x6KcKUPTCgNdITHwKw7KCPMxMfJdz/ZMbKSWDBqTsfPfWJ+BL0yzn
t5xKVkwY9eYIsywvYyUatfIFGfDH60xchpqF7u8CKVErcg/JY38N5G3NUdr0nWDc
MRTF/XS/lt4sx2QdTD+2dlPLUFqtaUqlpWzAD3sm8Fsn3VOGNNl1Aq3Q78oY4iAx
buc2eDJDp/UaXyWDEHZOfq9bgFS2GykoA7vc5sBSXia8y0JbEI9YE94BjYG+PSOn
JBjJOQ48Y6JXv1lQPl1oSGO0gKwfEoLAE6H9bGF358c+IvHR7AT0KTJ7KWZEYDLm
S6lEirsO0AIEyOsnZ5WGrV9hyl/ZKVGZCCju3xlHadKIm/NBINuxaNCNH6jeZ+oQ
37YjB6GbDodiHzrMtBbMy9VdLtpsMw+P7S/VLyZYMHr7Z2yo3UwSabu05HKHElvf
09QZZ9zLd2rBPD1TrrzeWsAVmTqrLm8tfO8bXpBHKbUuO5SjxOy100cMvAb/vukN
3XMYPo2lXaJ+OuCXL4YMKKpOfZfgsjuLRqbhmSm41TduFxMvLHVHvDt9GpNLpAXH
QWpA7KBvnV3VpaaO9ETPg8mr8JhSXslvRyuD5ECWp44vpc8m8+Q+Hl6U0vJrLEX3
+aeQ28/XBsAdM88iWG2zFqJFdNBQAHSzgyoSO9cOQVs6X6HyBEhGwGCstfoQM8KH
XwJcFLI1Qd/pDeHiNjuNOMJ4R9uYo81cb4bkDgkuvgwMfolq7lblGMADL/GkjBm+
hit3eOEMKkQkxaL2DY5tTEGF1xI9OabciX2/MbDkx+fMnQ/UAcOHdMqSjCshC88L
lY5X0J0sltdzYwUJn+NF9WmfA4qrcIkvEuJvNp9A57aQStRLHdIQ9VUEW3g3zswy
6Jl6Y20t4jkm0+fsB48GKu86ZGOnZ2y2F5BzxhAdg+o5sMoziSMcRzde2guE1PBk
7LVeV85aSy5mm73zvr9E+txa3QAtJBJodsQTTEwWdbtUPpbo1NlAkPHK6w0bcgxZ
MtTAsTdnHHhSXdyecHHHhwnBD6OSjPeeGoGn2Ml28IRGK8UAIC7V2z3q5dhsReY5
Asu2OpSo9ZrwirhrHLD55M/sEtPxAwZS2Dln87LBeT1ezrgHHsaEocVadzugLk+5
VvlQZanA2MAXWzv9wx0rjykVIvh1blsXjPthZFuGHp0FQqsDlgqIzROkaVW+OiGk
lG3WkYeYxrBTD1BWMMb9lPYioVaCTGsU6Z9uAfqtOOJb7jfI8BF07Fa7XmAtGGpq
MZxxru95+vBMt8g6hbAZajlro40TD0TIyVC8yx3BLm1DRAptFfgcjI2DY6EvQ5Mt
i8PtNOXQRku9IfQ6gUOjadRM/deUFUx+NC4V77ilGDyXajueDmhKhjP0FGuvmnBZ
8mwnmdwyd5PMvyERZFnn3fJfzwe4M9x6RzKmhCu65PTQdjXXFuTwSHIXySIqAaJm
7fSrJRIC/jUU/xHc93zfFbHVGtVyvDbSRD/h+fUlYPkVCQiw8IsbrUJcffMdzKSE
zB6uKNJBRUuw4HuUz1oZPsJdqRRFWi0Ki3lTnrcHzlZIczlHObE+ReD88dj7XSyl
GWNBDIGVE94FHJVFxwsnaS7RlWAZGRND+sBpnkQFprzUx0l432ZXU1ov0t8/sJv5
tVgcog0ixMJTO1I2zTGQG7M7c8trdkubhkLkpEewkd/wv4DkNVkm1n4QPqbPGoLe
OXjWLCE0WP0+mJDwkaN3t8ZoJIN63KJAKB/pPMzzHGRrugUjbtwqhzXzhAoOofLM
/Ez3Rv8hRY1plJ8xinSXqHpciplS+/A8lkGu2QUN25MlvPWWAiHwqBAx5EBlqRjG
lnwXuTX/KeOZSch0es1kHw0fvEwW48oiCMR+yAWnkU8dr53QSkFqvZ1652wgDcQa
FaZ9aixeOrb/tdjOWP6PSOuQPYHJL7P1hKWe6neBHWav+jHz0/mBcFyFEspFeHYg
3rpi/vmmYC1nO6HhFJZSvg2A3YFKAcew4SymY9qap9eH0Uf+cUph+eadXP15U3iJ
AYjSb8cVYyLU5n1bTmjV/a8wf76g6TbUbtsEeaK8GP8olsC1vVm5MYQlomCXXvHa
nF+bZgOAYfLAyQJhUHycWW069tFOoPkqBnNrjUTn7dDi46qLpODXIsCl348cLgSx
NzqFyzADWv29UXF3DJpn/A0UCaOjvjDyByDRS2Xc0RFh90Ht/7Gtn2sEt20alLju
wsDsliSsdBn7hFdxT4xjOwUXdaADfHW3AV57nAgfm5qmMs8DunpJzIk1sIVXUEb3
xf2GzkKOsBN04OGN+6XO79HV3XQ4PckUv8/WJd2lzk448iYw74FceBO+seO6yjJo
3mPRYiWb0akh2omZuuoOFuB348aEECvL0ziAUJM+GujK+ZdOHaSPM+/6wcMzxhI5
fBlKyaz4m9rDYUK7ziYlBDKtGMNPEfbsVM5lR4fjx4e5zFU9d3oRuo90Q9ITENUu
+l53zLlkqqFoq6K9IqW1fkch4GA862v4YMCTRiQ119BTk7YM1RGwGiH24RLwgf8M
m1SZDukKITnQpHhHBPBwQnBwRNpchSwuPjfnBjQv04WKW3eXeWW0KFshOfpQ3sHk
U5eqGAtgRbgHKwJAfuDRDdZSGf1AD9q/CS85OaongahF0mk/DSXwVo4zuNaBNQfp
sypfRjof224SqIOylfpEvbnzAj2ocDPVGLl7mw3d4/V4yFjg8nzuZOYE/8Xb090U
EUs2/o3dCC5VXB5Awajwu8PsCjGW9ZoHUGwdbhZjYLkyN7BKEl5+gf86gYJi4nMz
52KeBL1knP3uz/+75S6xWPdY1RISLczmQ1pTreD3tfHpfekciJheyPYQKc475+QX
25BULQCZfPxBcjzWgPCoW8w9r12Pr5ssl2yQ6UZYJJxb213XEfM0dg2y1HonSSaq
gcyv8k1SqIH9KwG5RWZOxuuL4XhaosfqVq9ZyJsB1Dw0mGJeOjSF02TIVb1hs9g4
ioLrEmOa5S1IlTIqAy1sB50RTKtKRrlfBGzIXtDGKYKDft0Pe/eONlmacERC7Ep5
BOtzk5a36yAQKYbSO0QCb6qhaqVu5qZEYwHP4FtIrcBrUhPB4OYWZhLuPAhO2eH+
ie14133tl+Vi+YpRfsGR57gUu/qSAQpNQtAxork+trUIqMnQmVgo3xeGiHSDHwki
6KWl7o+BwW74IyEKFKOTRkP8V1BZmg4IYU/FM9tphfwBmFbm0GRpxRhQ3d0F/FQD
OLkdnfs55PXmI7Zjf/BHiGcsPhjXOv+aSMtzxUHOD6LH+J48q6tWVIdn+7yANTY+
1U1HjKmKf3hNMeSjP7mXHccZFjNaA/IR/e1GhovrmnAAH03NSO6VGPydZd6FCxG8
Uk1NSpTjK4TvJsPM3oyRTQVWHaUgwaShd6v+HshSZhN4gUk+R5dLKbjIONzPI4Z/
M8PJbSjtGyz6N34UeD0EvSBf5BAQE+PE0IynBgN83R6eWU6S0oIR6z8kdINgjerY
hHxKfFkV1slTBiGtBROFcf2xHHbznkHYQmy6gA73jcNlYBFttp2PO0gpTa2B/Ijo
i/H61tr994TBenDmRRYBRC+0tN0YDvKNrYXnUJo4L8Xob3mFFzqjI3tevTAub/FR
DoMMoSuElbmmV6Uye6VLgM5eFkwDyz8ZTRWUUTJaE7j9DZzIf6D+WO6J9huPhI+i
hp5Gjljnx5dT4Ou8gcpaUuhCpQdsTL32sVG1wmzLbjLoqZWScfHrdq4BNaOK6Z/K
oiLw2zTwyMJJQzw4GrsN5iQm8GFeiHkVFThpVBAz1itxrzJ3+rqZne8HP7mSR/s2
rUO/5o3HJvUQWsA4Qeg+ULAn8s05dw/QeR67d0wrRk1I+uN19+fhnDhMSZqi7elJ
tmNzDwrDWM2YBn3NxoNy/pXxoP0JAAVuKMBe9yjo2ayZQfcZmekHlsFZ1D0FNcmb
y01WfaiBAFZQ573xyzI+YgZOhI5Rqk2xMUMZoCQ2INr30uww8uF5IWfxT4LcQV05
Xpfk8c3jZkHA0GAQhc6QoPMqQl9ldZuq6h/cPQ8TOf5hU6rfAEOKsKca8iRKgMiE
fiaAYmgwwjGBXmaDchGTRk3t5YehDYL0ws+FRbOyPQisQjVR5aMPS8ERiih6pAJP
9tkv22VtR1KjVKZYe/lajvXd/IkFkRyw6GooEmHlSvUkLmI4QCljUx/qNl4u8iZY
OqhRSdh2qBJjf0DfcL7ReTWA/KGnRmdim17B3pI5GJ0dOlJrFzN/XG1WTWM3fbTt
W2Mp3ZearU28YV2yrlqAt1WZwRix8zg7zG8n4AM/0nyyL96DLPAhE9I6p9VUs/Rx
4Z8XsZx6uY8RwshNp6+g8KSOr47VeT4SY9ay29kHhz3k+WDWfaBhHVJW5YUq81RV
jMyeFPN8X8j+GC20LJ7nyEgYtqwYnfyM1qBQRyM4+du5rrGgNU/b2t24BS8Cg/QO
iMHcP52hzn3IKlgtILp8Q36zyfIP9TPG3GjqDvztg+KOMq97erVnkewKa1T8msZd
HK3dd5YF54fIzCPf8sFV+Ka71VrTJH7du4SkjnvusJ4iBXasQut6PQRq8ARGwdIG
Tdv/+cUvruKpXU8Kask7EblBrCMl1ETsBLKHH7TuHy2yVk/DzSBZNXXKFHmxob6J
ON4HdP5ZWne9OGcafkc+GYtihuIKLaUwEF+9FSSyIIr1d1KYeyjwl1XaSa8YQwDG
GuYcIbR3QI+kduJh6y30NQbCxqzBev8R4/++LnVaKwHJ3dAw7hEMIS/663Z9H0jN
vvRMoaxrDl63NBFwTNllqxxd1oKljtkPwX5LSvHLz7RZid4tw3l858Z+4KiSgdbj
yWZs7tUolaztnrQui8S4LjlAmmTOiXMYB+cF5N9fYWSjOBt2Z8E7FpS+IcYTJ0Ng
/ElouVP8mbDltzHUsPPNq4Tojdf//PZzl9BBtm9OgjFLSxkoNfCDv1WKIOPpwYCb
16OnkWHHfUdcL3tx7tjaEfTlAie6uCR1whtFdKwVHT1bt7vjVylAKVuXHSpPCa27
D1C1KsOnOAnRLJ3siwNWqnDTst/uHeLNdbYYq0a0p/opJGLNL64Hepv/IhL9rDec
dyoDxND4WaIt1TU3QqwIycupv21PsW4eUZeCorXRrUxzO3bejt36oSe4vHYg0YH0
E7GlNK7hYNexdF3bSq0pKzqkxui6/bMsvBMtCoaQc0nT1+ndRISY0ogYzt70qVCY
hGDThLxsdSrdh3Z20jFYKAU+sZVSBAPU+cDUlViCbWj2kQmbPaU7jyZ/Pvol5AQi
vSdq6jq7+V6Yjm299V+fekJidgUol/Pi3zIMxwNQqAXMb3ekE2E+dOeXElc2Dw9P
3UDgiGF8wl6g4atRRTxgJi+HOXk6AXL8EcSuKEOXn4sEzIhaAFD+KNCqTspiGiRW
9Bl9WQAQbjhcQ45VSSrqmJpU98+jKx9qA6IUeRJ4XVGr1lsclCsa87RbEm0Z4AIy
VrQQRDRsIkRGhQT0UrAuC/yt0W+0uK6azo8pb/r7ZSoTWRJOe6BtCJW+ymNAm0Km
lvb1gNgXbOT5Z6U5HBXbefvMAi5gm2ZUJi5EZwF2sICXvJaUkUDgpWmieocjP5+W
A/a7a5vp9u209iZrSSvrtrRfO0GtLDcX4+3bC9TqzklupxKZTyt+dP3y2y/eSQR4
GyZP3ppaFgISp4/ytKqjAnQo6KEeJZ1E8BfMIwC6paESx9e9fHAq2u/RdT29PDHK
5KvcwnbJ3Eedb3J0OCfUgNa1xO9VVjnZenFGEz5C+b3MioA5hjz9RZ7jT2niIXXS
gwNpak1mIWJY4xJr4P7zlxBQ4KaRjaAiioWb7iB/SiEkJpTNCw7OBVRpLX6yKJGa
p2iRh6JmPl/6Fp/jYO+8zS7xny8EPpkb9bODUWplNW398PEwcAPlY0NV/xRCvQpn
ytS8Z/Qz3tcSnkjVxXtM8pCfKXoySXXYuePhq8WqncLdLeLBKPOhbtaXCnFOqz+7
1mGLLPPHN20bjxd9NxAY9uQQIWOp+uiW/ek+gZLUEZw0wAV4j5op0Q0U4E7Vch7r
3tgyocoTHdm1XZ2p239QAF+oVR18EufKnKZicdd9ZZ2LRZfnaZMqmtPOoS552I4C
87Pt/vryUKwzZuAS3LwHLIQ+6+9WQPcXuUEI9DDbsclyg6XM1Tafy6MVDvHQkHyh
NkZoDbsn4A/wI/pm/v0iFrdJ8HdwV7rNO+dxmBsOKSh/Xk4u8+yFja2F7O3t43Br
f6Z4ehL7IEKZXuoPAFCCQU21h+mS+StRl7V1KBEJGk3niP4tlorKBFYkNMqWc6cE
5aPVbSErpiabXdy1+nCL4R9kqAvRl8bT/0vo/sk+84UdOs54iro8HiaiyAU4rXYi
aIa9yYepJ1CliLeqqCqsbIldXcjihqKmN0xfgKtbZGdbQS74SN77SYaJpxY9TN32
VYVGYkbfEfWt73rwyBE8awZVY7PhS4ja53bUCa66zAW+E2u77RcTdGshEhaDF3Ri
V5mW0VgiGvR/uSMvDU3U73UgTGOSwet2PDIDY8ZgJJllu0s0euFo7aggIspjDoyi
MGBOCcLYx3M13XSjPth7rFKGgEfEDLQI2qg/ei03Usk7Kh6mykKF3jWyZASJH4LE
yUiEqM5hoTzZaEcO0ZnMvMOmOXyHVG3x+BrW+idn2BrWhycYYv1rJ9C8ssXLQABe
ADovdM28/UVx36ALr8HXxhwQ0401peFICitLysd+KEoKOpwCUF5sEgfpyX8thIoe
79UwonFRV97Q5pXHGlYtyqnQjfx4GYndUnEmN4mul56q2KCs8nGMTYPJbhlCbAtW
ymGEzQe81Vh8dIiAaFChKGtDHTSyKobXCSarf2UvUHLqr1TEcg1619hFihUnDaQr
V3xfNbHGXACdwus+3bEE/j6OoFAY8U6GQoSKVs1hwBnKezWbd3fRu3L0y6BbdSon
nvFaUUozGoBGWtIOcpdV4ShlpMrHkvIGn0q+dRZCTeiLgnNWDIJMBrH6yDwNMAIU
x8L7/1JYLgfd3WrcUlJXIIdwJmTy19UO3iRG3V+HSSPNNY3/i+J4C7VkQa+YY25r
qGR7n6zYA+uUlbwcPNcYi/gBWDcxP8kBkwcLZ+D04NfcFNt/eY2yyTRfZndNb7PU
IZdc55I3hZg5UiDkZ8ALF8YjEO2xWmwFqCJE5q+NLrKBkYBNv6Aj7WNsvX4t2k9+
7SFWjkHdeyAvtS8nbN/U5P5WueFdPgBoPREdiDdNi3sbAOmXTXPPCMyYi/hHA9Jy
M9A/n6j6ql8pyv+jKlhP1zsLrzD+N34bbNcW/gN3glWlux3YwZxo8r4iAOnCxG3K
grTDLoLVGXJkqqHMeiFraj8nvCwJeuA3/9PC69v1RBzoaITyO8DbPZYT2fyVRFs6
ZSfMmd+BiH8CJe/pNpShXO8UMIuFIlXRxR9k8sjH2syLu1sEuqpxkogW+zI3yIes
RTy3H7pAbNbxpcXRO0j8qbj53DhJ6fpvV4VY/gogoAxuSnNy4OcL/IBI+KNmCVeA
48cj4l0d2sptd4PgktVcql+jH3P39TPlwxRhBPZMXGuR98cC54Ie7ivUmVgz84za
+Re1zqK38K3ZLexefe6rMwAuyaxOiDMvLYD3Pmdipi6bP37LlAdGY0XX4Pb6TIDp
F0p+zHtyeKLWbx5GWidxwFaCJ5qlx2gIrNCf7rCtFDGxVzoqL6eEeCT3wTlooFsS
itXTARayPwthQttA1oEoH/siVFKzJeBo4KV03qxkBa8MXXgD+qetOuk18ZUo82nw
tC3hn6+YQz4cSEkgN8oTeCNop5hu8zxBMARTrWpuP78aGydGc9KfxpIqPzcCT7ke
ly2ETSFlCmZE6gVTC36edHcV8uoSXdJUd4NUcXj+wl29FwTjWSZM5T+7YVQ0tWzb
hdkS584dd9S5x7gZSsXml6Ytf1QX/celpcuV6WVHVHLcr26sohJhgs9DLfJfSSGw
n4JR4EcsKpZEHqYVkL0N0xTPCnBTRRdLoAsDqIYsiWAvptDPvfgKyeA+q/xH77LI
cyRF6vffMIM6SujKt+ixk7TQweI4H0bnPksv6OJBmz3feaV32HK4hkbqtrjdcdOX
sBqoryuLQP9ohKhzAHj7kGjgKdpIwLPJIGNpCnk9Bmw0wFLtUB7f8KPsDFNwKCsL
xY0CQnyB98PbkiAWVF/z2p7IA0odRYxX8il77bSd7zJLdMEKwgZ8I1lVPkxpPCZM
gmsuyz+Yphqx4ifHz0XmzxoewgjfobYIfAxNY6DCwhKBVdkKtkiaRiniL9imoB9k
stjmDvNmok6s+eWJiSEOWi0EUBHsIr+DqrmWvHH3TafVpazSzfkfBgopchbOcCX+
EBnNW3u6YprrC2AWyKlJ9nambH2/rVnr6iiCTsO/93f5zibQA4vcdpf1W+hbIuGR
/i63U3cjwGP7UC7ihMpXr3S9QwuS6hPhU/Qo7t96dqvb/lFmwBsqZd/VzsrLAQ1l
Mtzom4XUGsqwmfn7rDL3AM5CDlxaePXX3EFRnALDx6KVWlza0akZWJS7TshGuBf6
yaKRckqjYqJDKxxuJeBdQwqiNaju1J7PtUwFLUdV1D+dkO2td10woR/QwOEiP5pw
UpUfIG2Jzn8SBtcwTM6gMY6M6nMnvxatkfpnrbOwKXoj7frDXa3xsYVRpV3ta+F/
0adzgitKhH++9NcGXeGTMVzkB3RZwoXO0moVmaqcS+78yggwVNzv49VcHB6nvyS3
wGeZh42CSRQdhE3KsCkuyhmWWet+bFkvG+YjtMTAMXOTgcWtKX49Kjg//9XJOVWv
oFBZj5l9m4evjyZVsjoa9R7C+1riEsQYrfvCXq38lLTw2NdfH3gMfwcd2kHduv6L
WoDKE9/PEm6B6mEOfqPRyjLYSR1rYoRQSEQ1oRmRAgw3JyW9ni2UGp877L2gVXk1
Kr7mlxotNQoKrw1f6Dwd4ddixpGDCkiUwbAVN6SThfG0+bGt1zmzfbssxmcaEFI+
xHCLcriS9JL96IVjAO8sKPW/qqvc35rs4gxrp4/Lq5Fq5GICVMoTFhXtHwxaXuRU
nHVBi2oxK7JdEUMDuhaBPw1uAxnSxlg5Cp1UCrH9Ch6fDk3PfvSyGfUjjxMcWWN3
2PnIr4FLUa7WPatBuCl0dQvHb7jcWwkfo6berqBBQrnQAZXl7/9rnw+XBAQA7nFQ
mIx+XjsLXrLK/qewrKNwRO70+aEsX12jb6N3OAiw8Oa51grMHz9Rh1gC9Sniey65
8xumqbXxDOcrlxYgysCcGxg70mqN1o+xcasn88xMd09QFkMdhCG/4ti19E0uXGat
1HwgqUYsind4Z1uyARrTpo3ytJKMGWIf01Dq5G07+VD16cDrZnil47/412rrcFuT
Ohf93of81Pb8FuIREkgAKt/coge/iROiwrCV+ZEN6nbY2hyJ56f/H1nvDnePIITC
kGn9QXzMUG7RyUeu0ZmTsTe5rJm7gaqnsgzxCDAY4yDvgEXqE9SqVpOUMtNdwssE
XZRNkhB/rqnzqPko5FM7WMHCpoc6fz4hRELJ7ku/mi1kpL8uf37Nh/KPsnVA4w+w
F8Vmgl9QpETR9Ha5vpbCqDSQI3BlD8rEeg9caKANfSvCgUp1Zkp4Iy6x7f+SGgHL
NIXFVT0oQXBmFiv6FjHdJ1xO1jxQuNFnBXUHWvuraiftucz5Ehlmtq8wKLRF1F/G
bCTgZdHfqrQycltU6r/MJEOCo6yyz+mh87e0hnP+UIEMtIeySq+3AUMoKA07OFW8
782gCQZ26IakNUBO1PzMAjSwqizTulq0JV6WJ6LNyEhSKmlXxsbWt5b1+muGnQwT
zqbj5MbRcYFDdKrmGghUeDcZrtHeprOhOIiqIwEi5QOC2jJi2qqTLJYwq25oUmfA
yIXqsc1LuPVL899ftmJiOQbG4u7k5OA0jm5QT1Fnkz7tHukC6snMr2Irc/j6t+FA
GcI/7uS1zPsKcq6d3T/otTiMgTIdIK3gEQCd+Gis6E7mLIxVtWlobyZGfpfTeyIJ
O37NLqg80PtozLqY0Us1+24Fr5PCgs/s4etBkmpqncRAq39f4kA/ccbb6Bubd4q5
EOcObmjbpzqRWc0EnRW9joY62LYWnmuFhiRQGvbXcBmeo4Rn5MH60iWTExYPRyEU
8mYh4PYkCe6smjN+nFnApU0FYdl8yGm1u4bjv9zNQK9KkXidDcF+GWEKkY56vOBH
lAQ89NABFi7WB1LH5JuQuma5Ie3CGBMshfcx7/SRxxDw4MwBMAtvABOvlKWnadva
/we28qGetdtOFHO6cxLKPwCGCc6zIq7ePHRQp/CAdidp0/4jB9z5Om9VfMy4wuIr
cCkDA7kYObmkWlx0/KjXzJ9k3d1FlDRINT5u/meqoQxVXlf5vCHIEuYB+ReKA0ir
/aNEuoOkICJqW0EnPgA1r04pStc40p8qZSn7zJpK0sMPWGuTf5XHi7cnBxvu0aPL
9zElI5NoOAOgvADbSObSA+i1w+rIlZAXQKm7fR5v6iqef8SDkoCUWvAiu/10xnK5
tO9HtRDm/ivMdg77CP/bzDa174dQACC+akyFRGBUTN7gsISZuvPQpKIG2h0NjefI
k+1Nd2a2r9uRifnb2Jsk7X06O62in+wTiHThSAf6j5Xpr2+8zCro0i5kWQ6zay7W
mvI5Na1qYK8iy5b2EG9dyl1Ya94ekovanTfv8C+OkRsh0mHIQGMmjNUzz4s+G0X3
gjD4Sm8v1gLrNRG05K1h0RbdFCV+I+vMfDekS7GZzUSGLau+W37RrijzmTUnHStM
HZL4sueSJKHoHCkdNm7IS4stHn4jBupcQRR7txV8MFT1/wG8ZsnjiWfRj5LJSaIr
SwZRL/7atWHbNLIK3f3wT6uvQ60JsI9qPvRupoNQG8+FjsLrL4IuLKkVxVtTJkae
U4mnt2l0luyOEqOagtVaMcMtql6ZYAC1GHjsXOx34xoCUz32UdS4lVrOzF6HQxqd
ur2FD9j7PyE6UMidR4gHtrIVeNL0TH5Ni+oivnVVtpsy97DjMChi7JlguC3ztY5w
ijk2JuOW/u1D51CRzZedyBrU5urR7mpogEopU7uH8czJAQprmFSDa835iSExF4Wf
8qQNJ4NrJLlzrRvBNx7/fydH6qbkZdBJ42y7jVAfmgTjJO0BLdW72+dxheEDv+vl
7eV+bQX82YuLBxdf8Az6q4/nqm7ZwqY7lxV9gjvf9PBIpPljA3V5LmCd2nSIEc6F
SuizpFKniTf+8pnGUpmm1+DrjGjERJuBx0bN9IunWu1HV8qNHqvTJ16ziKwON1w6
cScOs+IXR97PazUssNdomgskSgC6loQ2WGFDOiKzNqBRnEsVKmLcVsYc14mqEjVE
qk+6PE9+fd+SRcK816Oma/YTgLlGbUCvsR+fd66bockTGN6K7x/wRP9GDt+dsJU6
ylT+PfDa5+KQ+psAly9uFuC17rdb0nyBq4u2cWsz6hMF5H8NsixyueaWMjInimvj
jr1SswkPZ3DoyxFNjuby/tf4XNt+MXTSxiTM2hsQMZJK+WQgsVgPmdsswpUDBtRX
b5EFpkvAzZXNfLxoRfKDDfZ8CUIcjqsCDSJSXMHjXFRc19a4gJBNotL9BsKNQrM5
oOtQCN7BYB6thhIEG5RR+f5wlStXsZuDd2SMSevXDNw4FFYhR6i/7uFStcqdC458
PabL9yWZdp6G4QwMnsu7nvM2XIgNXV87CugPQWSiq34L+3GuDRRkg2Z6/HtMvVmd
lc3O1cXGRSYvA/VLbio0Zg5J3ERKeodhv9du1KtlEIzeoqQDj/CqmeAVd52FmD+H
bVjACrKlN1WRv/zNEzchej/b3PiSyHcVk0k/26RaeK+gfoIn0fj1TRu2NDC/HbmH
gsM2u8kvbOJEkgqoNT7nH4vwiOs++3IYVZBxfHAzAJgAF/tHWc/g3MJ0lpwKEy6O
5LwmN2EU/0jSsox6hyiIXYkRtGu2aqcRbUZmnF2536qwNo69Mt4bsfLOq5aTUsdV
nWM9N+vd47fazKQ6FeSw42sQaRZyGIA9qQdWsjnwX7R7Icwhk73zrMv24zKzLc+c
4ddy7HRIdghWJUUtWM0pHRZLGmq5uhQ3qsiCS/IshFbqQk0m9onqFEos+M+66ahK
ZfZSJnKLaByzUMSpG/l1TUqRKRzyaLa1x27u7TfTQvUVrQc7tPQY4AZqCPDB+iNn
7mKr+L43IDx+CBNeSvKTEKWDXsZlh++5p160JusLpiVb5DB40GXf/+Mnd9gdhcUz
rzCCsZUfzWee1H1PRTdKvupfvXXJumaIbi0aVTXOjuHmRUrt9I8oc3J5ElPqWhaB
+XbKGqeNTfuHYP5FxjC1stNqcgS10BBJfFkJmcG+yIhV53c7hh8NMP7jN6s6j5So
4DZl7XC/5X/dJLNRBDVhbJ9UsRy4BcyiWrDvSqHoKt2wPvhEV680VTGw2giRcvVt
m8Bf5WeYYVTuSw7vWalGcQaDcNthyYAOx1IeLBf6BRIGQV+F3WOAZusd3RlZ3JRq
MeeV+xTk7PDMpUQBotba/oYM5og+W/jNMQIgt++mgqqeaY6on5I7nAqk6sbn4q5J
sfscowA2GjBrgp0av1+S983zJF/GxHxjmujm0bNLhQHs83mSQ2PidrNUTEtAbqsT
4r2bdvO3V1aH1MUMLXFtv+Wc5Mx8BYl4RhsgcJeRDwj/JMiJAJtow5b40hURYNgW
RIFXZ97IgbQFcKwQYP5Cky/LnaftLIotaK7ubgcVUD8ineZhORI9Z5TllHQv6i1P
+Y5S4P4GyoU0LOFYPXfAKfgZJwYiqKJqrxAadHb+0bgzhtBkuRn7QPecdkX2il3t
hqquxd0cIzjmUqmy4IgpxtPqFWNt82IXwF4a03x7vZZQ8bBM/KiGb2vfIYykOdBL
nEtOiwMGPctIEM03dyDIYwJJGZwB9Bk+AGbHqhl79BDcs1IX9Q5aECgJTj7NXwwC
QtDFDfSsZ9e/vkuTj/TlMrOORmmL7HHaNR9O3dXFsawBiMBVszuCldyyL1+Fptdx
/vcQrRswJzC3BD3QwDV9PRTOOO1pSGyymNXCmqPv55QfR0Fr/BxzAQ9jxcf5oeBy
fHAGsYoXIXKp4r6Sk5w5/yMADRr0c/9I1NraxizNXQRjLGREBGPhVo6pr1qb4fVe
kaRXUXUCZJ/qbHiiXUsZj9ghkayUfPhtxyYDYsWV4sQD8flTRjgbEsXwZymszCag
0fwuonuKvus/zmgBuiAMJvCeJITmzdwKTEZ/kSmL8fbGc3Pen1kHhXuvgzbFL0P/
zYVmOZelpqeRw8q4NnyFXla1Z8exYZYHK8DlTcSTGFTs5+lOofnsn1fs26JKchX0
H5r21XckgQtdGh6qpUV3gQGvEO/T3DW65O/rGG7MTVe0Ii+qSYNquKCxYtxYuDsy
0jzCEDSfcHtLzR9cSreVAPMengN70KJ0n1KUSm37OGYiA/7Clzka8sodCJY+NumF
o3w2wECsgMNypLRJzDXVyNKxYCwlgHrE/9ImilXxGR1S+kV9GKVdVVhIx8L2jfHV
8ep59tLxmArgTuaio04o4Kys82bNN/+zUmXlACQXWhf3nUtzUW6c0RsryHdjl92k
JDX9aAanIyLMTPqxuSVtw+uU7/gTELfaNKe959MZL7nLla1Se+wZhnbOePqTytHz
H4GyOgF9WlWS9BNsLJB5MHyAcAnqUuTuHR2Et6mEqK0hbVoseFYlEAZxqYqWpxA3
5LstnroEMVRJQ5C2wnlaar2t/kWgsWQVOjJ8EDr4WwrJORwPGljl3o2f2pue4MIG
2KS1lmN/Gxo41d9dAtAfbfOcJfahKBEJd4pVwwgWTLewOD2DcOjDkNJ5waO1fsnJ
rDnGv7xx7lwDcXCqORmjEms6MxyaAcV43c4o/Zg9KYyxM0466j/ehpbi01Oon+s+
Bx6kw+k9DtTP3SG938oovl24IbEab9vypQHbAKAUmbmB4w4W6XCCvohGdWrQW7Yd
qt1w/wg6gh/r42vfNPYicpgXEUFX0aNAZfqsh+V99m8yb0o4rC78dY84CqyVtmVu
rKIKeGRaOwvdRkuD+jaj66H8zKlAFJWK9bHcZ7X+uF9cjgfQD2fXx8SSFJPYULP3
uM2/Sr+1e2rgW4czz5pM/bsfHHkkq+KsKgrn5zS9aR+et/jaueG5hJ2RVoiEw5Zg
ansubQ9h4HAMuyRgdN7y4C3JTfQbq8yKJlOoCSGNHRhEwtd6/H+OcP6EoPW78Dcz
8pW1bCvB015MKuwm2qNjYifDAaPSUF7fh1qkvdDllryM/DSh3ksz5I7Sd/56dRum
2ri0NVoIX/6fWZKkbz/gCjYarXJL2TBMhDFvqzN93LUgTuvaRdi0OTRKIvko6R+p
wzrb0351ifYmkOMz2Z64lx/zHeIcrYsGkDu3aRuOBwN1wuWjokhcMM/+TjG5+LD+
Qhq/vcUMhNdRiss/4dp/iJotPGGFgSsReH7U7WSMPagmFd5cfBLKOocqrrQUE4Pk
0y7uBz85JD/U23j1G5Jtr9BSS2CZCJV8QQV9VvkxtzgyKn9dB5bEuIKjLwKaxYIn
Ux78gXLh5dvRFr04P8UfWzAwQ08sqQAm8yGifLJ9z87yiinjXnKTSleKT6l7+7RD
fb8zHu7g5tzTi2cPclnqtovsNDP2NOgLQ93urv/oijM5iD+u3gnIeeLoHtVdXuhg
6HffAidJ5pmnQhA9Fi7R3+QXa+Q7SXAuf6XMYzxq5fz60zznAH8LPTCoKuJKMneg
W6GqZanEW8Qo03mG7BVzR2UM6bFhq/Upg7HrVjaVHHgmgV76WoQLC21UprmE6itF
we8Q8gMcQgplyZmK95lH8Xl8uVnS/aGNa2y6HSeGb2VgeXlAMxG9Dj9xRiHtkHSH
Ut4HTCLqpgtOnFf2979qMFi8C+ic4JmE66J6mKmEfW3a6jjSY717RE64wVUJ5S/e
CKKJEBG+xYS02r8X0h9e9NBWDtrrTTwIrm9plLYwB9NIqHVrgk5JAy9T92RlmIDV
1EJ+G8JJn2pyRMXHV0yB83jcp7JGc1srLSkfHh+tbBObnI3zZ4aZQnUqFUrSe0qj
+q2nsoqVLAeoD2xmMuiW2ANIRjQwjJ4zHXr9UokBRvzJKsrb/Ynl/9WGEo7InsGT
PLzBp8Cd68Rv6/g4EmguDt67cY45aCuVhvr8qeht/S4NMeTnnMkuskKUAPNLOIxq
NY+DhUi3ZNq/DZRKc12BM8WJu614BkkfUzPOGHNilpeLMfsErXPDXgkocHkq7cm9
QHwbx+1g+cWp9a0TMqeSxfpvQrhy6ZTXmc1NwEZW9a52ZX9A5j3xNTKiY5APq/ra
6guySLiHbace9If423WoSotZ9w7o8xhJbbgdyP3l0NpAMfvYGD/C9VJhUagQRUiM
nBx4YU+SttIafGeU0nloD/BTVCpEjX4BJTZka5OnJd6ohT943p1EgOge2/84PtQJ
tLEJRdTxb1hZyryUP/I5MPlJYnR7KsZ0UwlumCNHBP4iomBx5iABgGzYJAbwkksJ
tOwXHGtu+zTgzALE1E0n7z+ZtzRNTmYf9qpQ/TmISI0l5p0wfNzLJ/ZWdU1nsjes
DuS9Gf3RO/CY9TMNFWXf4Dzwu3dxH21/NfahMsCLNz2GtEDFTSe9wQRixIVU1DYb
X9fMKL0cJivtUlfxEWhSwKEEUoiNv79ix9ZINt2M4AoStYW1G6OaS4pZD3Wm+ZnX
R1iKa0C8HrENtWnCbhwJW7H3PxLwwJOYngALcaya76TJd3IIaZFSQ2aneleUC3Wp
aI9eV+DKDllKJi56SBq2xP225YOlPYnjMjmKEeYQ7+k9pPLbublsIN/y6pWPUtqe
qR7Rk4PoOjSU8mgYfxBV21WT9zwdd4BqF2fRj7v923Omz9nEQ675ojz/fuSPhWtR
T0isc4zg1DrYKIHo4VL2MOWZpK4fRDj09NzxxqrNOjE+Mrpe23lQbhJD3HRA2pJu
5+jNnaLK7JHyjzZuPCftnCxchMTUO5kuTyyWE/vTWnu3QzQF3VGsjyDSoPxblmh2
oAaqlIs0E7/r7Kte8Cb+BalLl0he5+JO+bJK/IAyH7CEbZQGcykyZZui4+EWV649
BDY1TX9kogIROpzL3GiXYVRATZc2fvvUgGuuDjZaCpoX/nKCVMNACvCcJifDLbzg
vGYgO9ncl5SIVYMAUNAE6+h3Epe0DUbLVvPepUvau/zqHAH0XmpyyDaH9QZpYa0e
k+yD4YWm/F3aHiVJVzRwfbIg96nIKNlgZfObPY7fgfRLwp/nejv0MBCvuUQPWUoh
1aSJlgklfK4fA4Z2LXqXVWd7ohf9s73mAKgHtcsh+rOc4PRDYdwioB7Oy1PqYMc+
A8oKFj9/G2wsEbNZ4uLTY03Q5Plfs07OZUXplWjq9JupkIue37p5mvUrYZl+r32H
i1+ic84vapeIOEralskgQKcTe6a3rUvdl/LEyCD85Ak6kRoSVlYMNHaE4B+5ZkLy
RvgaD2x63J4AbZ410+9c+SbknVods3iXai7fXiybRMsxlI/n4zGwWRhU6I3Gj82V
CAbyWJ5+izjaW0f5CsCWjLWlENpAE95rPBwrid71RgZ/gQ9djEkfQ3kg2FP2V3kr
soSE6t5C68vUq3X05FQ4c2LOES9m/aXsJHk/dfYziwLYIei0+9u6ou3+lWiX6ZL+
Ff6GNY3jY+Ur4Ax4qe4r0XvL1BHngjo4RCMtbSNnqrtt9lBleIkB2gs4ST+JK5Ob
kgogUOdHpBgEiJzFmykOpykGJtP3R7gtOAVtRzw2oMLIVuU7He1v1r6Dr4enlyIz
/0iTWnu0g4dU5SSBOYaMxqb/hJ0atIwfKLFmleGensNGJPZ1mvO7IGBUz1o8CeNH
weQFuSxvXRqK/5A6jjZgVVDzJbEVLOTf4e3zrArFUk41s0nsz/k0JDRnjZOYe/1w
UOIYG/Z/OGkPU3izk/zkdt4W4aVXF7o/uJTsUINayNQ7tvnR3Xd5dcBT6bsy33mq
cEAQ3m+YvKHdvZuc67Ukve8Z6pNXkRqbhOR9iqcBCMWV/Rz4pe10bAUrcQvl+gsY
hETDjSHTLkUr1cCP0awRhhYMZrMtP9ljaYE5j/zcjvsKg1sM4s22GkriVsHFptN5
X2bmhS7si3GnSpP8DsepE7o314M316UV5aBRKGVh4aKbXsD3KrOmjxScWaeklNPK
0b0ZCJ7NG3WULQbrDgVWdnfR6SFyHIpww57Xqt9CRQnZr4U22RcKMN8kASvW653R
7BDVdtTNyEY+vMsyfLrLEqbDea8PLTtM37bq93s/2vsAE1Ab4xlyw9kQP4ghLw80
XHre+KGfxzYrnaU4SXNIrKtfY080I++rLlfYHoQd5/Zx9foYrbQDMx8wGzv1JxAQ
/hGRA3oDOdCpo/MkeTfLB9D52GUG3m6mgnu91V5PvW4uz4w9JCd5OFF0/mejLPIs
FqhRlwrySBGrYc5Cn5lRpSmsadHjdWeiRSErr558KMgY157I4RlqIHwp2H4LMp+v
TuTY6PkM7FK+uV+oGtLbbYzv1OAZfv2Ba72rS4n0a66CUmjTkoVmBl+RTHVhoqH8
7ogoWGnyQfRZhBgqsn20mxyGVTWVeNrHQZtxoMU266OxHgTmY37xqmWucqSwhyn/
8ZEWJ9whJIUB+69l6gsvAMXEi3OUWHIaO14/TAY8TWOn6tcLI1x/ujuQSK6uM4Ar
OzRUCwDMbBdlDLpUVEdjh6lFbNUjqcE+ORsPcNod8n2v6Z8ZKbIR+yJUaydG7rmm
F3pEUEmYxlDoKBZ+eUFS+5kKsz8qE6wF/nwQmca13Er1Ns8K9h/25jAmtlSy0FCF
uEAbSudCEt66spvVrFYCY1sBqR+TFPsrmkFxpaCQavBplj+JfbcZB5KcOdK5Vsh0
YwZDgifhZyo60CBG/TwPZR0joWtZL8IWYSeevt2siPSlLZmJU+bJAbTmjHqPhbG4
4YdC2Km3+UREGfd57ajxBirCu5gPYcW4cnEGt1vbmxfLuZJ0dHXS5a8QKb5dohN7
s3nxvrmXGpGzp8iZJHVA3G5VwfiTsPrFd6IURLR8njEc8lGew8vn6F3p7pJL6L9O
u022opE5nKn7y9f+5dPbz0uIQqEe2ST7UPERaAGQNnnEoG72K1spuW25xcrQDgu8
0mUOHywproatLaqbqzId+no79JhdojtB8Aa1c3TCybpT5FV1t6mfqlJSY62EvoDG
oeAUiwz0ipPhSmawSe6qQTRO6wOTcjk2tjbDTkEnISekxWV7a3RVoOVkvjRecI8X
rnzPsSagvG7qWL7h0Ad3Z5eib4t2hMws51IKDq0y0qPjI22zK7tqTWea5mQSfCVY
INWS27F4EWn3sga+LigliGxtHuT+PVz1lwVdRPz4CX8iY9UfbkdeFnre+373cgPo
X7AeiSzyLyKArTJDVvPWbNgjDNEedvlduYlhZH/Fp9zoyvROlzp1SPRq/6/zJQnI
ujyHU6h5c2GO/74yBsRcge/sAxSUOjCg9PUAt0MRBwFwNEtMUdCiGfXL0SnZnf2A
ey9GK04YwQ1dvTTZoNcN82P/sPFPw68ebaS4GqPd/qn5GGCTajHXMupUCCKKRrn9
tW3V9FL7WU0RwPZaW/2GsuoP61RN1uCh5gLqoVpOBLLmIyGNtV+bfj7tP2ZmYf4B
lR1EYqcrWg8Am3C5MxQjjPSKFypTbh88AKB/2gUiY3fnHpYbw3vw4F2A2W9xfdg2
1DZX2o53XgTfxYjV2enUC50jIO1GIbsLXPJ8NZfce75azILAT8tKHJ4Jjy2hKBLM
iAFfJmGNdT8lbvzknb5wQsZnwSfrlC3UzZMxFynCNbwRXIsqRap1qepNTGLte2z3
3sNHdvhtOqiH+4zItonjvdL2LGwIlpth158WYuvEet5DmimKOiujc7/iXSDwQsxK
nagzYeYg0VNoVoBU5rgQGwwKmhAcP/jrV7Tw5rDkUMAM9PYfwteH0j1yiPGT6ms3
osQuuWil43dRJWRni92dxTD8VYkw6fXXWkf2mqx77kJdYIJrXPeZW2nnQLGxLWea
+H6p6nWhRhDANijC9xgGU0yxzWlJnN986LYEkaZ+jxiifPsXgGyT5HNO09XXiB7R
7Jnd25pD4UXYyzASZQLJ1PWWNdhW2HZ/To/FyqQENICUoLy5if4tMa1zAevBH/3B
A+IV8t3UPglByOorInzXuCAw0d/kQI70bLkTErXs3mcXeWQ4yKpKx1/lMxBYC1oX
nL/OvQJoj+6XdLKwQRU/CHn99gubBB0MFWT0bpRhkQItwK7Mf91M7trqZzJKq2GT
AUFfu8rrO1+lOf5fcsJ+gc5LB7H77A4SA0aKDv5sdwDz1RuxrpDXnL9RwLwVnbfs
PgX7tGDbSWvfXZABiVtmYGX8LNNEgXopGiyKRj+kYRCwzLg2PKFQARHh+1BFdGoG
paZLewSt+q7N/r8s9z5oijdHDtJ9wTObuL2G8RTuKmYtHhFRzCxa3hjnet2B8Lxu
c2WiHpVDH9LcPr9BxkO/9DFFT9oo4ouakbca/0jq6TP0NzNGtZa6htNbhpr8P9aI
mGIiT169lSVZWXB8OENAneeB42XN76+HahUCxEMj2rR0nw1hxeY/FNGh3p+hCxtg
+jL1ANIu9nxaNM9ltNVCJC+VVvqcGeM4AI59uYrMfPpVUtF2U1ZmpI4sD7NWPZx9
7suiDHlNG+hrhnLl9RXkKUUsKVJZ24Qqm7YGMoElQHzwhp47b9wWzPRwahDVIz8K
DTNdQNh2f2blG6sKTgOc96RaNNRMmrA0MntzzGiIM2hQwCdIsO6EN04klMgGXiL1
Y9iaUybzYnsEOaW7khEv8JiCcAYlReByxqos3T8tjLDJIFGc15pl8XQUcMFjyDSa
KMCFVH8o6diMOhcT/dVepS7b1bLE5CAn1+ZvzN3dgjheXoSJB6lidnMVs1oykjaC
+S0ke3L8DsYSlke36Baq6Fi0DNOPdzi1vi/NODnBf+OhdvoGQ+mP0Srrf2FIR+bn
YIlM8Q1wJ6MpVRqikdQ1kA7kyLNSN7CenZ3eCYSHcgFJ1PXG3cravEaxQKqpTWSB
tCAsJbHqM/IhU1oFCYQnmzsa38fAjhsOkFnJv8IYcEmNf66P4STsN0ZsTW3DLDe2
5JQiT5tbLhIiv3Xc13FlqFIYYT3xVFprskO2yYTrB9PNWq+CsDNPuRq2hCBrxWwb
riyA6jeMn+w6fqy/MjZaLoesE9haeBcGXAuA54ZokZdYof7BnxCzMAMzuaA9vDBn
jdXpoU3fRw6r4eQXE4J5uDNGikPSO/0PGAGMjKGbAcDq4keMpkKQFWW/EVSxqACS
vSSauelysRPADrEy4llzP6xq19MK7dqGs3gZedX/bd5TkBFbL580fNzGbMaLujQO
Fq0paNWR1BOariHDKjrEu58eLmwCtc+adcuroMjuA9qIng3SskcvVprwG4SOHipH
zd+MAdjfmQyT0k0ZTvovQvZlQQkGtBrePI0Kg33QNItc9a2UrmYs5oX4FnO3SQDn
UDjNIA1uPd17lB9H3DgOqU8ciDfou08w2Q4uI4O2MoXj2XqKzfwVY2O9VxTZJLU+
r6DlLIftpeEjFVfADwgUOUaRXgFofG7M6k3x5kbc2XnfW8Xo5Nknscil7f4+N5tk
K88Fx4EK/MxvGn8N3poU6bvW5ZvHVnbwQ+X8V/efzLQeVHUJWHDp8lQxipLQFRu0
GrEl0Zxvmkr34QxajmOOthOfZXKGtH8ZE8EtgmAZQDdS/NKaemUi+YpaDyjiG04q
I3P9vVFD2QQEeZeEIwbhu8/TFzm1JBGXprzV4JrQ0HzgA/weSA7GmsPY/ZnZT6/m
ICqBdNgE0mNObx9EVoAxqwle5CWstejH5dWei3Dofsxp1l59AE+EvdvHULxWxM0M
9EePcwdB6G9nsg0wKBv354mHJxvPXoiBh/yHBbRAOf51jJ5E+s0JTp1ZprMAOTKg
hln8kr3et43r1MzkvuQXxfbUBW5fiWFYu2wA/wIVvsSglXaSnNQYTH3ZWsd3vvjE
3k2pvyVudUX6JZCKAeZ3I53Xc1hnHdOgnwtPoL3cnbzxooauD3i1VikUUKAE2O/f
V6HZZzLw0+kmXgYMqX3++RGD9DUAVcV24HiL6/fbk53KdnaQHhImWdXXcHJNEEbW
AGt1Jo4/Kb//D8nAKBeCtcdQF0LxPIIHavoGt50r1+Z9j3hKU0xnQYVYm1wAryKn
is8a99JLHr7hrchOrjWnyjId0tPLp1ufM/B59ppVklpiPa4IXwCJEkJBVTlEMx9M
NVNGNhspWM3LgQUPl2g1ooiaWJehC5ofJSFo7I+YKuaCBEu6+9oZr23oaJAf8Yxp
Y6TXDgQnrhNkX9t6d/7xMA/fVWPwrJchm92JeV/u66NeSxiiBKDnpf8O2dAjfHyF
2jgLpVXtwyVF5nNXsMvBl/XG4AIYGjf25BjBHr2MfhmQSPlEDGALOFspwPc5LCXl
l0URioUrpYh/qLdQB92eyctxCtTlHOdckEUzkVU1+wenf+cAJqEmab+/5yuSKz71
McIy9rNc9Hl4Ye9sVxdCCmEm6c9fGEXyd46Qm7c2GrJE9B+fzOiE99IPbEjFlUV2
p4tcUUI00TMUptre4F9S6NfvYOjoGhGGnDjqXkqwcun+wn0SdSXaAZ9QVKNYfbAV
+9L7QoFQkBCNlUNe8r/agfGHq2dUyzy1adERsG5uLuSL2OMh9EjHsrYEDfWGV+5d
L8B1MulbB/+3veuXiTw+aWBxJYlFEjCWVeU8Ertad5CqMc4ppj+bv/A+/NaGCGwd
GD9Wuy5OoqlLDV/gQQB0Ah35uVzn9zUthPUznyjGxqiMfxpnsWVRZyguepgjBCaR
Y4BwliAyitcHP//ozeQdqFQjGvMX9t3pmenti+XCfaQHHrYWGcFsBOFzJNE2gq58
uSeiqIun0Uj5LHJv4waFEmggEn0zWaZWVQhYtsqiDCZIvYATZ/JUH7odlXNnun46
rm9sVmtbqwGzM0W8abiWit9W49AHboR9QBEJgP0Pxiu80cYcly12F3W4ihfCLSfF
aWdFFmCusDgpddNUVpjGQCAc5X7F+x5nLNLtgMDOxQOesiXN0gkjnY1l1qWhlUYS
Z7EGdY6bihZjtyDK7NFvTI+F4louQp300V9vHWJjFglG8u0nl8HkA6mjpx/cA8cb
vHxpKmd3OnxXXElwrX5LYdI5XPl2lxnFDuQwpL0rPHZwhTTIIEPJylBhc0337iOK
nFoS56yMycwo0RviZSvYHakMbTew3rHbTHtyMQacQNs3saKVf7Bs/PvjkLkztI+g
/1O5ZSchj6ykRLM/BXGOXZyh+V4yYHogQrrava2M7MEXDpzUS8CfNj5cAq1BD8qz
EDPFk8QJoFdK4J3TL+NdCm4tP1Ukq74JzdkG2KSg7pde/bSngJGhAGl5Vf7yClTe
voyTQxz9mwKkTky0xiAjQqIFOO+LvpHDn1cRxnkktVOv+JMCNzA9iCzE1qnTlMbH
J5jJKSpcdueXjMid/GLsMwpJczXdle1HXPHIouT5ARM58l2VDJizZ/MFJfrCoiOv
bFoqBWMcmt9Le1UjOlrWMyoWbXEvoxhsdr0lq7u39NFPkenosV0Fff1RVxhe/0MA
2cnkKRtHwNsFwTL71K5q0imflZ5+BUtVTlEoOsgqijXvMVZDKxgpByt6//t+C8wA
1qO7EZYiRxrgDEjQP3izHgpZ2z4dzLhT48CuoCJGKyFj0AHJvEHrptukBaVYQSUr
qU9NEvo5XX1cfcV4gXWwvSMHzddStExWTyyp6VPdzBivYgtRhe0xq8H2fQU8Y1MD
2vrGC12Z/4sp6uBaexIBBPjmwa0R75wkl5wrJavVywcVxGINzQsYrKpmrAk+gNdY
lwe0R6YjfrbL09fXczoH0RFQ8F7rYlElC/qXbWhWJzE+tHh/y0DRe727X/aTqWDJ
I6SC7UbJd0oDi6gggi7f90LIAsX8b+dDtYSld3LU2+CdNeWQHesUPYBJnm7Xjkc2
AgX1UO087DEkZsm6sskgVd6ZsY9V+ucewV/OYQXLYeFFaAHfs0kxY1yVcX92y2q3
xXrKWJ375Qsmhl0rLi1ws2vh7HcpPukA48x0GWqEvUrNrFS+RZKxQ56pJBjVjufV
JanWsbuu20SSCTk8A/Ru+wY1cy97ir99gtoBdfAgwVfQLEPrCA3w5IC/lHrLiRNo
EdOkNtaGnEZdAa7Wv++i5YX9Zbuh5ERt3gen5Sbq+RTk05WHlVRFckgtEWhZQcTi
JpREO2Sgtg74f+zi99ZsrpqnhRmqKMK9JrxeYJkowEMAlcDSFRDr72Swr2t2JRmV
reAP6G0U7bdJyKT3MsPb0XX0ms9PVNthYu30Xijp5NCHWx+xzCgXEjp+npjRSBGX
8AXATbfz3ImCGVz2T7KbCBmqJK5iKdSa51K8RURz56Sd/I4x2fRKOapyza26/2+W
5ReCkvML2pNdWwhbZkaCjp+DSIpxjj/SAaIyHNRe4MyQ20DQ34Stdh7V56HD71pz
kHJqs00emHUOA1K+NRqVNbEdqQIvmet9SxRknUpN2YPUV+8pe21HBsXYoP5y2VK7
6BZsoXwV36S7Cvggcv2Qs6JAz6WSshlCW5OLUyMpSIp6Dq74K2odi3i8xxCMPVzz
q8gNyvbFeTFm4oskPsyIvUSX+y0uNHjD3Q6tX+g7JOh1IeIzffPEukKDZ4O7UaUt
On1BQTvJrC65NHEEAghKKqEGjPDDDe7/MdxhklmTc9cBXOKe1eT+VNvICl8GDC0M
fzwsHzHkfFnvvoyleWP7Nc2iUOsjbx9l3vDSOh6Zl36sNotpOTl6pkUrSnaYKkH4
o7HRH+65Zt5nl0C+4aL7EaL4Jg0dRK9nMgoePdazf4t3cYgQvPotFRbLQglJOZF1
Da1HleTd8UzlO3cDYyHOucRM7nRfWa9+BOyJlU8lsq716h3JWsgdh3xtMnh0ciUp
lYPZ9YljUs7iUI3Xf+FAXXrPgn7Idxcow0RLNzY/LRW3G8uzlYhjeC9DQtz8AvHe
CctAsfi8mUcvVK12+7uGNZMQRkKo27JZSXPmBGBWBrG58Klx6pQqACFRg0HnNibC
PjbjFLWSEzBk+46wnIfXdhUVIA80W+VwyCFr9m/q3DWyHg9j0ny6JYUlu4Tpn6Lh
e4S/q7fRmode+SupgHx8goYFB1rBVZD/w8ip9RxhbhGUP5f8mjLpoDjzedVdVajr
Nm4bkiitwGJsi2paacGLnTSfSoCIg6hExrkmAu0uPgo0Jdpb7YnSO4HqM8lTUH8L
qioSf+QyJ3dA+PPajLDBpktZeTaTcZvpNefNDRuHYygW5Lr7LEBBsS5zn4n0YQmj
mqoEN7s3UyAWQKerybvTtJf/tegooqe1vF6hiO8Su2gQ8KUfeQMX6BlZ6OoZo+yn
1yLKbw4m6KfvUyadZ+M/wS087/IMqX/HY2e1gy0KwpGZd6Vd894tJ3ZKq6cehWWT
DiMZe1G5xXAX3AJTRFQyZ71yvNoom2t1zbN+TkvnHU+KQ7DH1eR64zjidjSQ9ZH2
Q2Azw7i0olzsrXWti+5r1Cnu49nPd7Lk194rBXtF34yqG5zChnF/bVnR/1qKIWmC
1j0a8MBc2oIlkI93HwwwNZkYSJUeutHUg0bGhClCG1D2lT1PQXDEirMaauKiAXL1
WE/c3fmrhgggD+KqLZv+uTNWzKAm2Bv9ll9CTEH8lrPbCIWtTnDmKuRuU2dY2TBs
q8gXN73bWeIFRb3GDDs0/nW5GOAGpkjgenE54g6+Gbfvu/gCr1TrLaYln0pfJspb
+U/ePl3cdxuhGT5D4cC0R8c2WSpoQa59wHk18AFsrLgoXxTWhBCWjmnsQ7K1Sijl
VmigGKzhJqKysDH01KydVlu1AZ+Lxx43RZM3fRTTuFcYLiSqZFrLhq72YYoAyZjs
re3QPTLU2Q7zB4WJJ2Fg2LwQxUtAPDTymvRMmGs91oS6zvmJUbMar6YzTGRqWO6q
c9t9rGn0pQvxQxA4F4lDMRs3qjV7jgt2tr1wNeky2appMvOEASB42LkTKAN131Gj
Jpz8U1U+12Nq969QFK6sTHmr6ovIvU06Il94FPRK9ncormtlajnQEpw/VPbJw3xO
wHGXJC8lhwYHVg32ND1Rwh1vV/Q7U8Gx4TRzrRWB/55G5aDewKbZ9wxqMWwWAAvx
JmZbuocDKf/zslZSoGzhYJxgON/ydmm3sRfszCoMvrbwEu6zW1URGBGk/FRjdIZE
/E6eexJDD2LJvpOLmPkZW7bfGsplY4XWClXvqP+zFeKAXhOsi2eESye60KNj3n0G
Hnv5xFG0v+5TDY2lYp/9sJU+ynFFRJ4VN2c/RqUYoG3pex8SgVG3DWBFVVIw3MaN
2gMrTBlPZxKuME6g3RB8rEjHhGVrCEGMmGm/5O4C1OZSAo21kJkcOCKTs30M9O4R
o0MkVAX9JyjDD0QcAmtdj4ApWqnqQtozstdOx0NbNIXvIUHdVMeaXbci/qTIfuEs
k6Zm7MKfodP0quEk+6t6jWNiXx7M4mHrdoyhEmSedOPOujgOcV1qovhOijVZi/d6
ZkfkERoEONOkyszQtOmIvsSCNJjcugDO39PbSQy4xGwktTrcwvYJ8l5vzj2Id9zs
ycvpGgxFeli/JK+iYxbM6J61L5hRDZKRnqYltLLm3pdpI0D76mIxcMPnwSggr5xc
/GwhnGdZCmOh4HrL7NTrl2rlCJs3tJMQHmusPt3zojbVO3jvySBMUnTx9XWYqmpP
qLoOzLefI53yViQYnc8JNXJ4VRPZY9gmxsO+/9Xzvm6HsAiJOTR6wBDxQNbcp6cX
lLEU15jEr2yuMxVFAeLKT5ZuCutcknlBZzyRKggNzm/1LwZXAg9qW2ZFMqsEmBwc
mLrP9wOEJoAum0NQrwU05jmWi9W08If7R8n1+Q/VnNzT9Qj2uvkMJx8RZ+h80/mC
zUpGZg2XLWjpSFAJmfGG4dykhb4l20ytczLAGG6UEhahV9IxmojEhU86Hrfx4Oel
7FUqcVdZAJOT4ZSmDWjOU9b2lK2oATzmPF/f/G3QlVynJy8i3cmR0oye2K2PEABk
CVubj4ICqlh13fdLGmhUGlxUWyj82+HdAUFfLhoCwcAwrqSpnDMrCCAok99rJYr7
vgTAytpup0CKG+XkPxEQMFyIJV+frv75TuxLKW3ewjaFWk8uroJTwVGBoaSBGL+a
DiUVtG33dyCP5m/Ftd/ri9RbGhjNqSXg2SLCoj5hR+tVy3UnlRSS7WvqtlsG0Wy+
REiP/LZ/IaL68e8kFqNarsx7Gt3zyGbbli9W+ezlqiIG2+1/q7x86hOPi67RZpkl
xpJROhUXevxDvZSVa1vX7RDfw7ZBFuMNcl7vafgjur5y+0BcZfv8DAqIkHOpT5SA
Ldp/TaD5eQream+NjQZ373rMK2e14nLVXyXjaiM8+v23teTEuBG51vPF5oVDrd8e
tBkm3VmabPHNQXOB0W6Aaqr5DtVRezsxqT5Fg2z6RCeSVI+As+qICibOtrkWxs5u
/OSEsM2LaVQqN4vEjIudQU6by9mLaTfk0G8bZ9vod29dVgqqfbgzbDNHi+k9s+22
89T7/CgAj3WaNWitEzBTUas3LSouFZzPG5T4k3l9uWdxK+90h5jfyJe4vN3ZKhE7
CIlgHLKEaUI3A3HFAKWM78VnDt1y78mI9tjfe1+sSHfGAeqsY3WVa5Ts7npgyGzV
06mTWAzrhLxEqlFv25nrY6xkF6zful0tPLzrITks/nlkgW76bMJckNuHDSKpZGvp
JFNlyl+NcMH3i1BxszY8iKrbD6DiUOtDG58VfnnArTylVyzYwtA6z/9dgsyJnRzY
rL0WEOCUrHvpPNhat6A5PipjcNxKqGP6mBJi/gCoUVbSPJwA6nVaipiqmtPf06Xt
2LSiB+TeNSbJnevUqxet9++Lq1vNwjRxYSDpN5nSoEsg+aKNRkIsr1WEE0Fs0bau
T/GXqeWpSBZzNnWFsGc3C6SfYn7ikv9TQxW1tsz+HwCEvdc9zQVBLYMCsmszO3E0
qTh0FoZhLnUvTluvB84SdOjJ7/dgy/CmrSIeiqO5VlxjX8Scz0jcl17lM/uR72qr
o2u0JCZN1dWpCxaiikkXZYnb4UFS1ezkL++NHAODo4tRlV6G057JkkSXviPOuEyy
mOSk0uhWPU7P3TvG1hARb6Hm6Q67idewHs29I3W/4g2cgF4bSzHpzmWZBDjSVuzz
Pp1Bon+Ix696chJNQo17m2rb8Z/VrBjr0JHvBvb3X7fQAzW8CY5T8cTPeCnt115W
aRRkL2fBRlYf6Mo6oJs8rKCvUMHXRXa7R4qhqPZrMrvHhaqrVh+BY7jCs0u8gwSQ
em2kxyuUKXs9GzhB6jxIj+Je1/j/pHUCGAMpfIkjKATKkt4MfIrYeBPZaYMVd/Cl
hyqLk6a/m6QEfa4s7iO5WX582q6U9qX+BUaeIs7G8LW7qgAX7XPMpXdmWtRgsorD
ekfdqbv8mvtgTG20+mT6sjEK7mVG/N+1iAzO7Jyz+7kh3NLkV6yf4fjshjXlZavt
s7CHTRZkGGlUNSqdPnYZRa7Fvsbd9xy5vafD+M165cGoVzzlGSY+Yd1zFBU1eWKd
MZGV9b2G4LzEVJ0nIlUNkxT4Hl7fZ83nS6kbtvrckkUY5bi0vSl30dDEHQ22MT7N
5xSwSB9PI+B3Y9hPKMr7+RzKEfxYam5vNDOmZUmA+QrB18N7h+rq86QZDW6zrsid
wPzuqtEgWgiuxKwYpwiP26g+UzzXpS6h0iA+/G9fm7NFEG1BdkB86uqmClAdXMA/
wCQtM1Q+uir5b53l6fDqDW30APBTlzAe8c57xRJdySDg1ibr6Lw4WsUt5E8oBwVB
QHqa+NJEALi+qPzxQjcOkp3+sGAMqV9sPzMZt4SLg1c16J6z3BWNbZ6MdbsgvR1U
WLNLCZPHSWyxYtu01+Mn7Y4Fl5lOr/0ceJV94y3kgkIVQBWk7drzOJcCuKST1rc6
xaTOEeNkerRCJiflbygvKizSSCDMZSBnzDNVwAiZin7Hc1H7iSyU+Nbybu/ROJEQ
VdbFFG8Lo7BdnOWf+DqJVz40ME1kWfts5ejSdbtwkda04RuvZSLDsYaEONt2Mq+X
imXKeIvPK+kjilrGeBZzmCmxXnYXVWP330KSQ0AIBWGZ7uaOPAYvDIchwNE9wNY8
4PQajPsvTCV61xWYRa8b0euBC0NaCLxL6LBZuh7BYNTVz/TK/ClnInigB656SgYm
au16Vbth7ZzYCKssIRi7si6Dp6jsaMlyG8oOn670rL6DKUhqV5ESiTmlHTeTb0Aj
JOTC71yW0pJ2txe9lBOet6gAbhYCn+76EZvRMgGc5woPE/NQGs8ORB1xso60Kuyz
HI3Dsp9pw/Q55eGSkVIMp+zChXeHcqrD5BSh7GYJyLZ+u08Od6Pg8/abSdo+wqID
WlB7P+y00TtZ9P6xuWVFaqmea2nDSj7vRnNOSYfgoO1bgVbEeSdI+otBnT9DtUs9
H2GPkElcYjb3yffcwdZ0KW94wCt9X3bozxlf+XgBmdU/A5e3mNJf+VoJcxEyvcro
iL9JiQaRPZ281VrMMxSUVor38rcmokWgyn0pCXvVcGw89dtACX2xE1/vy9vK7XVo
JwtW6Y3Vf3qw3EHpzn5OKIHPet/4I2NBVQP3GsZazSvAz4oAKm0HxDiW96slHLRD
AnkUXUrxL1NdHMtRnwZcuBqbrJB8hgdc7oBhLg1phjbGa6Ijm+ZZQTrjtGI3XZTR
xS9E3onb8jzWKaCTfLphoKsFODOXcJiyolLpveq5Kuoi9IBmdLfPUehdQgAPL1UD
jznFqzP2fMVHh/ly0URLVcZrEQ4fYobVLI7XUu23o2uAl52b1pDli4TMqZ0jblkW
iKDkukyc3RR0QiTcDuloiYRuuxsXqAA0abuwTJrl0HlUwTSvs9Y2uwR3gmAiScaC
2tBUyP89VdqPSMaq8NWz21oXrjaTj3d47pHUxjALRYi9U+LNNEyrwL2E7AffrU+n
r87rImj8LDE7517RyxXYKTiY0EIi9vJ/ixzpw2DWFDWXjFOFcmtXJj5qykv+Q/xQ
1+ZkljET+uAtATlDTz4hWUdp0GFyuC6UjfA7V1lvSenzBwjUnAWPu1jy9ppUVK22
tH8sR0DFEIf95Q5d1iwFdrGFq1qG3qA3DysNtctjAC5zNhmlD+2MKpgSNMGhP3jM
PIT2h5TYjoRLr5/wDxD0dKTOpzzD0pCsZsuIOH5g+6uXMHFFZ6lc8KyT7RtfXHNJ
2uctKcW9b6+jyx7guzlS2s5+Cfb3M4e6XCK+4MtlsJnfaQXAD0NWWkL3DhbjwyB6
Zaj7jSx+nKC1Y09kSy68mvLFzBg0XrxlO8zU+Y6OnmC9Ss9DtLY0BKSFnPZkcU1J
6BmiUEbOfSKUrXlAUX7QSdsYALzHeOvGY1kfVpUesShTmMSgqF4V6rmu3u5m9u3H
Ho4mQQMySJ/ronaKlS2zw9WsGYsL1tEn7CA8WWTSQZqq701eGMMqje2PjdaRyv0/
UJ5PQ3H1KVR0rcALE45QsGye2CgDRFtxMG2cAVuLurE1/22S+hGNXCx9yYgZuTA9
76XmVsCF91t/NXgujycod3G484aVM3couNcKlrtFIJmlZc3UlrmCaLpjHwKJWEuw
yjh82D6F4+1ONEJrusZwmLursr2gsCJeSOkwc2+giepny5xmFONYfGYzBX1lBFlW
2IMVQ4SKCBMFfuntne2C0HaRG+AddbIysyzjthiW7DvNkq1XRktJeFwiPYz4NK5F
/GxvTt0f17NAZOLWcXxR5r0tvHmWX2fK+qIHddSJ6xRdLqsmkdJGTTQPcgDYyj09
yhaK0+YIPBnb6T7JtP7knf9u6zVL5y+tnJXpZZTrpJNoIC6JIyBqVLi/Oy5qt+tu
QhUcew4jlqkYc9E/Nj/OHfc6C1cIETc7ow52vJIM2qxemW0V2RglbRTrZrr1Bp+D
0KUQBY/o+HSP638dWWjPKuksandIb2RjrqHcNgw0FK9L3uTNwgq32iPIDHtJqEqa
L+JGfeUdrlrIdH/aiqXcAeTDHz7JBykdJl08lWal+DCy5UwQL6F9oSnn9zeAEb1p
5DOs9gEYnwtmQLE2K4klZs/xrk+q8ue12CebjMhTbbVgmdBBtZ6SYVZ0icCkDb0l
Ef83AfH0cQnLDmO6BuXoTgZefnJFj1ZNTvMigtg8TeA1bMS3jp+aHZr0CXjbh/gx
h1LiU/yTYe24dqoAYJpJhebE7GEgOdjRV/J4FyLcQf/2QYZdvC8aPC/VeSTVLFpt
EU3850yyc87oScsTUncBBRXmVDbdMsK1nxdV0sIO6fYzx1ojt6HRooP1AuoD/Z/4
J3dCxJJ5uKlyD4/TLRz+UdUaiYLA6eqqhwZ/PFbXMgHWyIUha0tHEdogZi1Vzibu
tuQtn0yDyrVanL5Kkovyd9ex68oqtZb2ttZzgvoKePznD8g4tnQfWsv9hatQhfZV
to4sxmfFmE7xaXz4SJH3sUuAkefb3CjJPyn/xEoAPplQakdmJ9qbRs77PHolxIa8
XGyv78sMcaE64giQbQlpyKqud/XnnvOjDAlBmexyv3hitXfLfwzpnFNmea8mQvAA
TaEXg9/wz17qWxYk+lUM0Mv1dJWnBzMRtSn3gnHKIPSzQigH16CVGwnvf6I6S/Zt
z/E60z0N9fyht1LR3Rm/1oll+KtxDO2BiXpjUb5vTKLFNBMWLb8MFjPQtzxyMVnM
+dzy1/bsT72lbltrg9sGlPji+mNULxEjx3lcyo6FDTs1NHMfNeDblj6cMBmueC+9
/DwOU3H5NGlsEZuf1vQupeLQ8qkchBWyedooc0lNSKBRe3DdVihn9N5P71QhNpaV
3pUTLTPrqq0sirlOAOmCUw7GdXb9cFzfCmSCf8uYovclk1eI5DrWKEAPUTRtTSnv
jW4RhZ2trFizWCfCUnAlkHBwtygVIwQp1JBF4+MfdoTjTx8ZplzjtUVoDmmJQHW5
7VwI1Ak46cfckg5Skc1/FOPfAJfpY5ABYFPZi/q0KBJ+q/FU1CDyGvqAQbJUOCU6
igcTU7Vl46PN2ohy+rF3mfRREiVbNCLtYVvG2uoNal/dNJSkjdmpTp7NhTDvttTR
lmvaJHul2bdzYJEhGs9slwlJwzZFUidpaNUqr1SAk9oYGLdg3axpQpx9s689CcBQ
W4/ytMv/89gVdikTwceHldnOovRjd5+8s2CtRc2AvHZTxJH77+utKD/sixqwgf0/
aD927zwsZ7LUbHqrKhFP8T84VoUk8ZrAaG6O/mqToZvzUGm4HJ1bM5GUHZeFTTP3
QK1A4fzDMPfS4nfkpckS518jsfGOTwNERuC2Nd7+v0ILAhmPsJXFmTlXSG39qyV5
sfqQz7JLD3BBFr4GSdIflRr14m6PG5On7gIQbc5iZEsrTtBSHqDAis4N/39xXbuY
eKIIjOlKmp4rKLy+bfVKvL4TJsumcwBn5V0lnPj3LfFXnDDo+e6HHCu+cME0PIxR
gy709FJN8vTcaQD9TUiHuW/r0WYYw98MCz/NRCZvxeOQqPvAfILvVIlbwxsLa4y4
CSxB5mCSWcv82ewBkoYP3n4odT6Uh9VWDftv2SrlODtNxVIz6XRgnxQIBhvBPjKc
vXQEvXjTsiT5O6K+Z8+aTE8koHKsoP0RKbcd6dZNdKJgVLV1xufyx4pBaR7WqLuM
bwA+1pJm53/z2s2SlhIpur5mvJNQHoyJufBIeK8hDi+O7m1TdI9E4zfKTMzWbXRW
I5OeP8mDZwuiCAQD90ZiqkRhF26uKijCxbUYeOEHl7XCDbS/9CQbIkXWFqgS4GeS
mvfNDZ458XZm2rxE+BxbN+C3Bv+QUXi6pokgiN+83xTQdrJbmWI9DNUIawmZyeZ5
LmLAvplzQglSTX1mM+C6WkonUp1X1n8lG51I1c2HEZs/dcG+1NaWnec66YlTBSU/
JW1xh9N4LQ8LzYosi/elwff2Jozc5S5wFg0s2TwvLsV+sxJIAYrrarYW25yUv0g+
YZ6t/1eZETTvzVCHNu38VRzXvVCJFM50aCH+lXqsSuUKgssSqb6UKz5Cno/qL0Gb
hV90lt68y3wtk3y9BHkwWrELprC7Oy6TF1P45TXX/Sy3wcTUBSo+cjlCSGmlYyrw
abLiIDqAXghY5yTF2mCAix0ukCPLruUekIePxAMuYQnKIYyY4Zqnva5MMHQVz92T
2MjIjfPG7jv2a/Y9/oZMrVtnM6MIEQiuyUWIx2iUyfnePYDp9ukkNbUxsxFqe/yc
yy5uHtinnWCahIOlUdJnCaMtJWQwrG8x+ffw0IT9Ne0ZQK9tVKz6syL0Uw0Z9/Xd
fmulL4yTjf3plWklPuKcFLTNRP+dC2/3w0kKTf+9AmCb5FXcZXKNFoU5OaGDM6DV
MpLBMLyMUExyxgFXxCfWZ4gOKzg3XV+Q1I1tSWMqcoM94P+iyCGWUi5e+DlHna3Q
g033PdPRRmhkqyspMGdVC0t53dLMgyJqb472cIBO3MA3UR195UE1rIt199DuRECU
yP6fVvrh5+tNR6+YF8W1me2i+rxxhROaXUzul/pgzc1/CR99vrPNzBDVLKT2dLyx
4cTWhjAJ+0mqs4/8MUK2zj5COGebVm1lP54MRrKDDB/x1SViN8/UgWBZIMg+vOU9
N2R2+3YKiDYUaIlmR4Xx2DBvPzLC/l5iUcwGgmnL4lpmryYx7sekZZDgHkLz6msE
PT4pxsOl9iIC+TUYXreVVaKsxBUOnKGFecWwZLT85CRkNS0347Seb/tytDuDSW5y
H0UEoIFwQ4uVe6kAhZw0wLgw1wym6ctw4SMA+S2NWz8rryrDoNb7YeTpk+q70w+z
VHV8p5V1mqpG6RRWQRUmuvd/sAw19cfuzC3dT0TafCinKxDplH7cm1RJ+cGhEV2l
WBK3SKUtHJCkYM9LbRrF83P3A72CfnF/1IgVyThXvXJBbzLj2E6mF3ctC4qn60tM
ASb7coCv4QyZRuzFT+//wr1fnOyGo0B9fY3vxD5EzHLinDH9gwr8QgiH/R0SMek0
+Hn9xg/sZJ0+KQrB5Wu6urkCdRkn8IKvprsEAsSEdpWBMXCuq+CCWTBJxGgDFGFN
KMoIe8RBKulSOF8Eb+FPal3EYqVjCLkQTZL3hhC03IWpKyL1IScBo7+jdfuaTDgN
fL0ksiJP6/O0MVeXSunGKQtckIEw+5J4Gu0Vk09+mpdAbkMVZrJEgIlfoDN1yzcz
98uJCkR63Fw0ZqK2izE9otW7fbMgl1bnA8woC43OAuFrGApTXYqpraBxifYx4gfr
tPs/oT2bmyrS9NE4m6sghKr8B1oO01uv5cZj0riezpYvOZsUaGy2F+P7hNgDzSp9
ktrUWa/sEiaq3tUP8L6NGtpu/ZrH3CV1FgzUGd8MlWe2jiPEFutHll8XjpeuxLVF
+8CdTAUrhjXEJ0NztlBxOtfYfToabXv15L321CUBAT82jK24sn0Dt0PcbDCBxhsn
daCUCowosDkA79C+u5Zfl1zUkaS4NfDLqeII6RonbJ/ZarRVQdH0EaGfL+C2/GTg
xktUTIfwa/b0kXw2ofnoOMax9cAewGs126spfY+jzxeLcAynj2ax7Cv371ey82FY
an0STuaCTBpmre+vC/DHtCBI5o9U1HyvxzjABv0Cpsnz1VvL12ahtg+G2tCmNihE
8KR6CdOM7fqWP35y9A9YW0Z8Cg8WQ2w9aKfLyWtuM9/Xp+EXYe0IxX5yqK9F71cr
hkis3FpisUuJTLVhp4YioPwU61PRMyF4tRTZ/WuI96Z1vO6NwUyduUu/2Jgw2ez2
UYGi0Uo8sbfETobrMrNiDw7viqYlXymJC5yS9QhHlCv+C0nqoPe7Ew2vsCa4bV7b
RCaLmo+6x2oWObjGgicaNR0+3EsgwvhYtc7jSj84fN/5s0G6DK6DdHsNcPV8ysUH
JP2x9/U7mCtbabyHaW37oRhqnGvSjXjW1ShorjigjMyup3+wkkUTz9G/ScRhjyGp
KMdwN9KFePsQkgy/gLkxDmTPV43pe653G1EkxQtklEVXHznhu4Ie737aO1ZosARO
zBoym6zzrTWLQxkdYKO3W4GxQmkVQ0grDaOad3vDf1BnoTYfjEHVQI0Jb6AllNaY
8CQ4wVDU8fgVfzj/330XxQtpe7zit158GIgp7iSz107kuDBD389GGiUqRWuz+NvU
0I06M7NFzvIUpWWf5qnMZiLlD7a5MxxGQE94v+HWWzV0wBh5fRFLqdEaEvMenx+3
fVUn5iPkSMSgkMfMAU9LO1saVBDnAYEm67hmyX4K0DVRhd8Id4OKblD7gM4fhAwI
xUWvOF0Q0/B4ICQ42tEL6QJmLfiJ9yvbxkAvheh5forybRzu0OVLfj19GGvqBYNF
fjblCTumsyoamK/QHHpcbc822SBsD+9mMpLmdEwbprnSKA+STCT0WdPhFJw6EAYt
17Y+NOMVM3574zgkvcscb9UKYXFc8Ikq+lW1Eriepgxg/sT+RDzqT+Hx6q46Pui+
yL45Ut0msLrZeIa6j+t5Rvdmypi+kx/+aMiNetcU9bMxarCX8bF54M7A4X4MSfV3
9PpX+xU11yt3wjdDbCVHnnVOkdRVHiE4dVHxbHlr5+PhwfUkvVQwTA/6OMh5czVM
pF3VC8pneQj8pEtv0rapVARXdDzsW/BedyMF7jsGbjzuTK//l88SI+e364zGioQE
bqVkDpRijxgzvxk26unIG5qNS36a9sCgTlmsYm7MOzVDTlwsN71oXgbBIfyZEgpK
Av+1QUfpFzyPz9jfQ+DS8kqAQ6k78GNJfXn8pe5/dkq6Yt9Jjni+z8M56hJgxDAK
syhtM8FiRKb6a2ILh6daKs/hfJlIwTzLy3Qcu872zRTp06IuCx91EnaOgktKHmxa
dahWolsUnGOK/4Q9vNOXVnlS+Nu6au0zYN25Rx0xykuG0dkVVAXJK+nmilA6dDJf
sqgbEbtbh5k6HVqyeXQW6gkJ1snLCTW4KeqyR7byXSJwDXeqgCukA/6Ab4drvL87
oKESwHSMP15fFEC8WTRJ1G9Rc6lbW+3HRhfLjPUIYheZxQGgq8Pcrcc1POujxXpg
rPuzxYWyTe5WEgRvH1veo/u9CGZU7BuanHLMQCUrUEZcDi08LZGrHoH9JE3uoY3W
7q3IC8vQ2gqmOxEwR88eoZe14MwR4zdSpwXZtzLtExwiJO58Cv5ycvt5LNVYXOmM
mlzhIto5hdi1xvVQWaWJmfZRmioA0t3Bx3iNsgtdv4zu+0Zs9qojhELNciuZ5mZX
QRHd4gfyNlv936xhzZWsfPjbNpAtDRFeRoOdDsRDlkKc1Rv0qazXbUTQxcFYxQ01
7Nu7lSz6QWVpV0FZWN8erpY5QI7RkJv/1edWeq75h59uccuL4NkVKmpGB/HG76Ei
yvS7oShOvq1H9t5yBe32acXwcs8OqlzyDWI5CC8slCTxHlYMNM70wSIpgDO35bTb
z6c61pBb8hRLAlPjbgE7qBqlSo1leTU61qlBqlWfP7Tfg5sZVDqkm5bRRJRqgffS
KSIbPUbOO0CZ3WbZRAatQBVuIwTI261foASm9BoU6BF0GH3VldeK1JuPHyA9oMs4
nuVkoBLrzQp43aGBTKCgNoMR/cDAgpY40zSZUHdX2sQMdN+S7cqljt/z6Jrxt7q7
sltifziqHH3/7/w5OGlG6nrq3gbeH+HMgEZgGSbbvQqDz/gk6cWY9/LaEwwFXUoY
424U5IcGMKz+k5MJqgAec2E5kmi3s1gJjQOR/Xn/gq3ckOeqTME5JWrMg4sOQSmt
GWyE8JzpdUZG2I4NWxY+oaxUfNlBpeCL63fwsQiLK42Cm2RgQdXgzh4nq4NzrYsz
EU3QhctKboMLnylOcxtT1ffy2ADzq/hF80AzyNKYhFeK24m8qlrfC+yig/HtYEDE
0/M533jBwQ+v6+XL0Ae6Q1/QcFyEKV30Ux0HTltKMcPoulzesOWvQfn1RfJDZSOP
T/fN6+ONzgUgZpv7mRNJMTFsUiiSbNzHjnQZZb1oxGE7KmJm4gF3ZQTbEcCb3cNz
buz1HVnjN+oeZjlNJin3WRHxTGc0qCSks5fZB2ziSRD4RWxtXsAvOFMkJRcHaMoB
aLLG51cxwLfDd1vL8Pf1qW2CM/kSU002ukfL9eTF+3aop+EoTWSeD0r+HLQL5+vA
UE0Wsz7FS/rNW0boOQwjCIc2q0pHdsD5mCg0yFBDQyq0CdpoE5ktp1qa3Kt705ir
PVUU0bH+0pquUCNHpDIxBHfkMiFWZPNTkze6m34vV+OtKCnEiNZ35QlAvrNw0TTr
bY4B8K2uIFvp8zliTRODzGDta28BImMOA+H02IPwXFagNKwiHvjCcPVmULxjpHM6
fYmD2FT4Am3EMVnSr8IJrOCI8ycdGbb1Dit5CmJhfbeIwv1Y9PFz/txhbwM5l+FL
so2OvmgFR7NzKc/YXKW1z/u5Iy2qGM/18xXXPvpwDW3VIlVNc0HTbkXsFPYsL2Zw
JjvqYoMOIphJLZd84xusNF8gM8hk+lbnuOWd8QEitjbBAgwLlNE7NHcHLLK1JK/W
FSOGWiGCAmqKDwKxdibIPe3gu5tJvcUG79uuXV3Lr9WHJb3XLCG7On+ZjMK8fIjH
yaY1lHQmPqPj3TVmojw/S7VFsVZRWR9tTxP6Ue6yCfzExzqiER9TBRvA1jpYdCsz
Yc36WTQ600rovvdZgVig333SlO4L8nvuL0p2y7xov1/4V+5kfdE3Gia8gBWTSIXd
nT9be20ceg5o6e5HfsmoD2E86vbjM0AV6ADABD6IgPkssW8CoBdwz8FPKhsTP/i/
C0ndEO9NEayhxdhAU77BK5oQvjBH6dKX0Cz6hku0aYUoBwds/tw0WzaZbxq9kuUY
sdWGPjFtHxSTr2xQFJiXtvF8gLFiIt52WdJJemDoAyckvAKd0vOu0ukSS/sI2ZKo
tMxDfPjDepo0L4rMdaR7njvunCKvm5RfS3CK/Ha37N6iSyk1ENhL2siYcgAFWhCe
aUpSyJdeJbXviy9MXDQ1yANXNBRvFkqB3+HPJ0Od1LmmUiHR++BIVbe1nUtn8wrZ
heM6H7bhDaiLvTG1SXF/urPzJJdPGAeDbHJqPbMqNn5s8HgsMsO05AZAwxqXXZGS
GA9pTnI6rnba0GB2lb2BhFDxGP18lSAj6/PqwA+4RcsJ6XF4YvnuRCS1wIBPl33T
YJGi6kRFhYYGxvlmoQDyAx/fbjeXiYQzS470HfAH0j4IfxIg+HZ3MYlaHfSeETMh
SuJnqvPTDcI9XhELdZlkyPEqUV5FFLR66Q7Uzpf7fHYqEXYMtcoSvOQ+tAPVfoNc
QJS+c/PLqyJfdjUYpMCT6QRoa+Xi3OaFW+38NxeZynmPX+AiK+8pak8jZ/C5P2a9
OZ7p7y7R8byzGgwZ0T2YSNgTlZ9j6i7gSitP0UUH/hGyBWhk7FvuTkOB4bWxqLoB
AyTuSAyKvUWFvahNhYs3Wy/gPyKlSOkwUYFajByLaCbYRoIfNJ2ZMFIS89rvJCC7
VkGltYsgI/D8vIgS4dk/du656iy+vN5goGooL0LWvKQnyLOC3SyAI3MzGkhL/rc6
XYaldQXdlgSY2e9pLPt2GdDGg6eXr4Odew3/sc4FQdiE1yNA190/WUpXGk+if2bx
UUEHIjuiSPTer8udF7TKFBEKoxKfvLoRLgnJSL/rfBV7bVphYWmrdDZFNdSXHUQ2
goDh+oitF1FrrrrHmoTXNSbCaXm5a29rpHGDOK7YbACftMK1W3Ksyn9k6F9j+eU/
op344+/osnlZiScU4i0pHsCHI/FtBiEKjaEpBGwBjPxiWzOcU0aHJk33SyaB8ZeR
Ku2fbZUefrmcSwNfsLY1xbL6btcjxNuTblsWyJKuib2EGeMCis0WGfE1qMnyCb9T
INRyBpPyTjBkAg1y9pft/Lp21FuGmNpFnXoJ8bnKR2E/5jFlqjL/EV6GzCZ6G4q4
BFQYF6qnF8ie1BnSRWs+jY6yCi1FbTo0ova7ypVa76CdJLk6G9EHZ6BwupOe9+Vt
o1ghE8hoWxqE9XALzr131h4zXfrDyguTXj0qzJTTpQbuDKJ/iiVtj1ujBLJfdzT8
ZK7DMMilAdehZxra9wQ5BEomPMpwMuisOkti+EG97LgU/XQHnYuhNbHsa4JYwlaB
iJeUbrnMg+REttUZinPwiW2knNOj7QXFEpMwzSkvcyTZp0Cu4OG2qTBJllDxxQiR
knBBM5g33POnorDJGCwK3SxGGxEn4DbmzVDzi7mwnn26S4/+Fdzu1i8hs4Vdq+Yy
K6UNao3TX/lck5vqVtBjY+8cdQhIJ43esHPRDJeY0/Lhms7A5HyYjEgLSEXk6PrT
4j/miJ2ljwfoovzNN2eQeMfFpxnEiuENMmu2KbLZQjoWo8u6iH20En6RubV3rxJK
f/PP+W7pARNPdWOclUbM0AlHwDiK6TCKa9eo3XVNAcNI7ZPhyijK42c/DH+t4vFU
oI02WbSkOAJIp+4Bxfe5sbKmAP1pPf4FmxoSjFqOpg7kCBQflxYC065Iw/Lh64aK
7yXTTYh/1h7F6jYJgaF70LjIXFsxyvOzhwE7SXSWKeXk2WEL/w1K/XPz6I2bD9Kh
jjBZBZtNtq1GanRVk9+jEqPhVOXU1AO6mlHQdPKxMFJwwJ7mkOaRBbWHqc7fZvrb
crrfPO4XX0ffcr/MKqv5mMYHjBia9Pm9o/FzGqFFE22j/iSSFVAmqUkOZmHxCu3d
xloQ8Zj8xM7p7h5n7HdibJujuiEMiaNZvfW69+RlRdWor5nrBqhBwGrmJJwiQU/T
g93M/utCqArGrKixrDb9Vbs7wIQu770FYCjMemKsgpyoAi/4rMtnrmI2VfGCWAUB
r9NBoohVWIE83B4zMqAle4Lmu2JVIAACW07vIaEB45TarMycX16NY0+B0RANRtzS
2GkpE2qEvphd7LZRYnXm52LvXuhlcQn7p6HtZYPZzu8hk7XLOs1gr34cKE1hdyuM
cJXj1d8D9Bmirud+eNccpv23zRCw19V+XU7EGjWJNkrp/T2v+dROqOfHEPMk3P3c
h6N4O+CKGi3AocpFBD3ZpaqnWgE1YSsKuy7ZcfkOIaF4I59k2ccFfTXDy9OLAB46
2jxo9sBaIQV048g8QsEPEm3dqQmki43EugAE3/jCGNWCn3h4LvyIGjAv/h4CSba4
xxJc/JBJOvdy9RcH4ZHCR7ZHlpXrZpixl8+OTL/iYgw1hixFtraE3v30qmtYvzeb
NoYWkoVqjz0FQGO6kdF/1E3MrYf4yJ+WYVSCW4hM5bkFlNuAymb2cbCgWlM0zytk
xVFvC+hOWzoEdb/b5DPNPqnrueO0uRhqEoApYUaMR/ktB8NirTlRIUOo8MVxw/F0
VD8Vy8LnEyC5SkZdkPDFiZ/ZCawiURpwiKX+4QT6kMd2sejCocdKA49gTmm0wuU+
8tolyYa1gIXG8+UC57UPh3/Jgn3dJnqAB6LnizuuWwwNKFsLSvBNWfFbXNyx6TGL
ba1vLtEEaRSKODO+U2qjo1T1JrnG+oXsGbwDiwDURhYNkexQ7V8DLeXfRZJzNIza
Lh5WQ15hiGNjXrWxMjgQ6g7fWu/VlA3qEd36toNMKVAr3VHQdMFbWX30Jimb5nud
qWiiCTM8sjLJiWpdPf6nWrXfDZBbpxxmXMNSx5LBudobTFU2DFD0dS0QLnZkIKFG
HGKRtV/rDJ5fmeNX8ZJqwejKsCI+xWepGQSA2rB8S3hLI6AMW+hEgI9Z3M2zR2Bj
DRG7j1qn8/O7ARd2RWlCaRyn7Q62NiPh9XQYkbMe7nUHbHkM4oySDkoMQEZZ0GAy
8YGtT4vdMJx2LFBaBt1qO8QXgNNbnfHDyQk+oZ9qjq/hwQJzXaqc8wXRO1pFyeyp
NWD61zXrnQ/wDzj69qI/+4jxAImtPeouAdM4vIW/cHfXvYqBPM8JbvtU4hnXhu/9
VvytaYneTzHoIE38JjDu+JSLndlRxHzvg+jc5VBr9LkB7I9ArDzjYXcQe3qy5y9N
b25hAX/H01nHwDyQeyWxmBRT+Jt9+XHKLkylyDVCCprASZBnfjiPYg1gByE2Xlhw
o42bRmU4+YZK6J7knuS3cFfcHXWbvSW0DJmI6dnBZAUV7saAe/Da7UPlRcuzvmrV
VTjEuv9mP+SCiKIc81JIf15k4zeilJgSfgz4V0Af+1K9tQ0MEDlL0F4mJkxyz4rD
NCuIzK0fEh7MlDfylLX3GEH/ZN+YK/hSCoCVR/oIk5ecLGTujkhcENQaS1nfG3Tj
XYGF/t7xT+8gavknqvkokSptLSr+1/Gbb1aeBhW08j4ytAFnODHCV4lf9crH1xtp
ZtTpirzjIpoQAJiX3rqExJiOYgA7y4zawORqsW7Qwb0xMwgy81PC1PSgj0h4eH9D
nEWTlrmzVPrTl1//N8c242QdGYvvBIBChaaIit2RHUrFxvpEqcvDrWg8Ip90AoNW
QeQ5DqCijeXoDpaI8R8XhqEOyIzHN8WljJNiU1OxOezT67CSGi2Vi41q56CFRiKz
YzoY6VqJHWTh4HQbsdBM5ipKtVRtNw5uTDlv5apsOBJTlKoJnl+AgQC+eSsr165d
lHTzSn9y/fdko/TWBh0qXr09SRo4tC6iroQAc5Tk83Ll1h5YbFSsl0eUUOoHsIg8
XDbH+exk7+JPxUQO+QRZkIo2mqDvGX8P+IjnK+FWSBEMLAB+vvthvmeklw/Vcbwq
gFl24BAufjpeWVY4v5dmBxSxzXlwhM3oLy+yWaHbFcpxiu/OTeHVg6MmO//fdHl8
E7j9dJoce2Gr1qkzVP0jfOFGJcKpf62TXSOLOWJtzn2/IFLJ9hVdovaZWbA2jDQy
BuE7NqjHAO5oCJU+u9PxG2PqiVaiD4R3ZCj1UmBzHheYFzj5jpVsG3xSi4lVt9lm
MAi4UyFtA/eclfNe72cb2GHuxOw8vv97P8EoosUyVoDzyp3oxEgZa/21KgWXBMIb
IBiTOTBWtCACi4U0pdAR570v255pfHL65BoAi00COlF26S32IfaJQ3KBriWtxtiD
ATxwVA+x2Ye6viNp6KtV/6bYi6g07TQ22pRAsSYiiAnllIPjPvVEP5ENUfE2pt+s
J/XGhfNYzyHZKv0yvZKzof7mY57820JsSqfY797LU3jZvmeQgq3EcA6X0KRvBcsl
x0OhJfCkkOw1hwSRSkIQ5R0+GSbQp2lGfqkKbVr9HR1mpRGUWPWbMFU8ikYCj4FS
1EIx+g4q0rqdH1Jws8UC19qWIUM5snpQ8/KT+/GcsBHowRbBr+AhWQmSmuHcTFe3
gK17yiK8Neplw3ZADJlUMiP8iXbgErHrRPX6BmA/EqHg9MJf1oCOqWOIIvCiNwVi
o3XYk4Vy7XVH4NvJH2MTv9DeqZoAWyRQl7DrIou/8caTGhBY+pmGsX79q6K9pwuH
/EbdHEK9M7M6Ej4BVKmLW/wrorHkI9jPPc79KbKJk8oU0nZAOaZVCwlvB2GgTVH0
W1DSh+tlXEOwoWy7ZV76xfG7simt6Iuvt9h8J+uiYDY+PhbEBSfXV2LWVkt81Ihb
C9XIJASZgSedIprN4ynk6mCrqsJGKMO+0AyZphwM2jiUkd0VsCZwdP1Drp6Tcel4
A4WlJUZ9ZFb5YGG37V/SxjdUd+0x8iz/tyCd8Z6zZri8w0lLCb3k2k1HmX4ZlI+3
nHC1L/2E105semdoGW1rkg+cxpjZ+YBQFkisEPatESHvrKr9O5dMH6V6r3Ebe0RL
XP6dxgJobjFyIgCSeosPb4R4GunRv4/NIQ5LUOswn9PsnFN+VdHZIJI+kB+t212E
RyzPp8oXHzQWLvC9nwoQVtT6ywo/ypW1jdoEd6i5a6ROV/u8kSIDurEJS2bLoHmg
fOEVU4oWZuKUjMXTZpQgfj9K/ivUmjCNLHzdONXcH0c9uLoQtNrugzMXsztZGiUo
eSdGnUoX/V1b+WIYOXSKppgwjy/hZ6B75s+4HiEE984DI7UY1t8NLJ/5sbLYZgtW
zGxBzRsS5pY+odNdrUzUDbLmfUIW074Oet8tsl8n92er4+RbXI1z/laaqZQ4YWu3
KdppKrYJ8W/fowsY3N+L72EnoSKwDKIYvCqVeolSnwDNp05EjqlDVK/HUpr+Q4Gu
j8BNjlE7WaQkdyEtGgepkx3l0ktefwD29JGW5cwSPOrzCRTQB2uGKxlMHK66zOp0
ElyqdBLBC8oZTKtu2O5SrVSynnbD867UaJrXxj/8v601yc0WQJb7mSTqoobbTX55
4hHGJH/CFiHv0ih39//NgXFsxCLMgc073I5uhxchHfK703DGNi/4yY2WawsNhjlM
vYQsbNNwQHA7kDdrSzROSuUJYKyxbVuzf+wSPIvJOkBuF3SCdhJm90gKpXXXh4vL
8wg2/L/1ZKKH/oRLXIjb1Kpyar/EmMTd1+8bmXzxL/agMIef04DRX1mRajD+WcOh
1b/Tz22+TuZtFs1rfKvSrPZ6/jrolnGhUAvFkBUDzK/x6zjkcvKLX1N7KrEXKT7N
CIj2r/lyFL9OyqhkZoBN2xPlu3L4mLoA+eeWbDC91FOLfTUTS6nN4r4ka62xsDtV
7lz/YfoCWn5F6CQy0fSe4WwiM6SY8GuIqLMRlxcSPbW461xrt0+1OlWLHmA8hSX4
9wSP5RN9a28Nu38Eo5BTZMjpoDQF2gjbdu+FIAmBpS4FhqruRIvqDqooU0H8WNnN
l83vJE0EXAhG49syGv5TiWsNKbE1AedqvaA/t/mbwF9eC2567Kr9ZMS/x9cxbtcl
pLexYdo2HR0xn+h8l9RAhFGRVpaUd0vDoenl3nQYgXs/MoeIM6KcKMAwKvwekpPU
Wm0KcBKi+LANgGAiStAEcno4LI3W0nphNjTycq4aTEqR1pXRH2q/dX443EGNdoTi
0PsQjUwOzYw9+Cdi6mkIFmj3xBAVY1HStiejW4OD2KfZ8xBE0ssPbv2oxPRal0CI
7X9j+wOUqrTA2+MrB3ygI+7YBx3wYuSHDGrovJrlyUhuIM4QkIHrQK43f5Eo71vd
CQ52NTGTQLoMXesVSKlwukkQ+v1MEuYJk/9dy5mMRC1MYQewH4GJbrDARHZXoS5k
mYD9qRDQakYKSgy/D+EDiG8+sFN1rQOy0QmtqhwyK8Ui5LdRR/t3UArjaL9wtb9m
8yclg28CcCRKS1L+NcTSbdAs6NSda9MSZXMaaXk6b+bNDWw5ryXO4xsgckr4/jIs
Qb1BY5d98F8YBGRYqFyHuap91PNxceIilaurjQXMlo4tUUsQeP5LaRMMQTraAFXS
b7VVpRxhPlJ+rzU/kVC84CZMhirqQ779D1b+U9JfqBaIwJxe8+Zx/D4X1YMAHRov
jZaHCTYN1FxBWpUEcNXjUjMJfs3XroMqWH93EAE67RiWIxypGDhO0imgZX6acK+7
MuE5f4319f+Rer4p6SbnFuQsQkYu9EilwFzSNr/4RLQZ6EOzf/zujP4psRYdaaM9
hAoTkgRj2fyFcwJncEsFkTqn6o2ogdQBYxC6fzi1PAUq567CkWWmHhh6XJWcl394
12kGfON6OtRcQV8F9YiNCK+74Sc/UvJOvjET3GYRMOJ2smI81u2EFFMs7wYttL5z
RstPufvvS/RqHtwEwT/xXvK9UMa2BWbXQq1YMfx1V1X/FCCygUc1L4YlsuOSizBJ
g/6dke+tvBwYqanjhe/f6iqKUo0ZpPifpSdhrZkaCB4fdU9xR1i+6omul0CwRyhU
tkrIuHgJH+XnwLsnOdQurvVFzXXzJhEW76tbdlIfTZnCz/09LD3npZRY3kBAQ3h4
aR3sbvDphaSpOP2F8i7agyUFENyHPvx5TLKOXrU7SbBNWpyf+R+p+KQ/Y9vZZNej
tXbf3qdkmsVg/7zCaNRmMfl7jmUz7LVAFOX8LHtKg97CMOEMdHAn5opYS8HGRv8+
DchPuu+61qLrsTRJ2I668n/CpzSyM4otdKJ8zbozEaEIPXCW11/Gys6VZQgI/gQe
yaG/f0WKTycmv8Wib9swvqXWqcPFY4XDclQOOv2H2HEJUuFnCYB3RMS506O+bDkA
Ldr++2LD5QMH3BMAZ5Z3YPmLyOEhHphcKXAeT2ieYiyq9wpAv67ofXjDiZZzCIYT
nrQDYJU/Fh5X6iTTvGkt0VGnCARTzvQC30cx5OuZcFK090BbBE1WZJ4ceNlR2SaD
XqnKuzAnvKCC66u3VbBwsx82XO5MgTOHPe9JbGlckr4UzXhGojTwnpleRVjeTBQi
mv1wp56C+Lua2S5xm47+SnTGodmzUMSh8rPV1EGwSbEtpqhdLsSHroRgJiL/hlyP
vuzF17nOxo9YKaWTOIjHzXe++YeN3UktkuoYWxh5+zoNIocryvIAd4YcqoQs7k/x
WcyPI7fXg2Mte/jF4Aa+tT96NHRx8L0u88T3Z2jvqzabViot4iIVBetvEryjiI9b
fnwKzg1wi0jBSrp/AteKMzftgIniLTE05MmAFn4YKjLQSyHbhUFWPd7JOECDEhpL
n7KQt2FMy3BkuAev2qs72SSnuhDxtds554+M4DMqPFy3GlA1boPUYBdNLb/0syb2
qZWGILCVYtZQF6VQ2hovmbeJQx6OUXtewK5xU908Dovr1qm869he4I2TPbDceWi7
f3wqdAdE5vI4DBnbWRTl+6DzVLmPAWtb815OpiFMg6AdMyVXQhmo/tSaCH0d72Hw
akRNj+tNjN1P4Q/+yHT/cLxrJHxt+SY3NQ5m27vmYkcREhuCpgLkZBdllW0T9mHX
DlUBEYfrhAV5GoSdAAeRoBAvZ+41DUbOG4mg09geMPHWLwQ7DvMuIFJceO5OvhFu
HiwPu84GXhoPwyNzjuVxk5iu/N/Ryqjn9UZ9o3h7pqMlW4VlpAR3G9FNfP9S0CYG
LVIZF6JoVcfknhukh9ku7C3c4/vIxFIbTUFcnSNmTOs/5so79B1TcjOqB5UJ3hIr
cscX0MDv1b+U7CngwJZLO/2s72TXI6t3JzKVgJ2k9Cg6hxQF0F/kuVQ7LXlhqRj6
rP9fkH/6VQOZSVTLTZ3p5JCKdhhuWRrYEQmjI0PAROlsxMJRIHY/HmVxzR665tso
IHJF/CMK3ZBpeSgWsdy15Km4Z/caWj5E7UtcJSaM7pVjKSE2MbmHLR5PmW2HXNfa
G0AQsaMo7Bx0ha0ta8wDpZjGJ9sZ2Q+w+S6ImUfbCkoPvEzLztClV6B+LZCIZhGI
EKCcUEZYVJb9CILheFVtcPsVAWYO0h8IRZSjjld9jhI/ujVrPEzhc3cXcP5+oWBH
CITLGvr9YY///ILrguCaCEsr8e8GftCxp8HF+jZT7rZW/AhM5dseIu3m4IEoEtl4
rZT7dt9sQE/CeNHVWkX1iqMOg4QJfTjzSUP69ZBD2QyJZZTO+zv5km9msGP8JgML
z0Jztjfl/9fFkn6Xjr1oQfds4G3NIfRHfVbkz3CW7+loNLEuehAb9fgPCuDgVpT3
fH7B4jlpFcYE7cyTNyyHO+HJJ+fuuL7hFknZVR62Cj4itVQHAQZvxQuxjN7yS8H+
ik++wNdZ8ickG593IZnfm/HPWffm5DWQJ2yMXlQAqiLgB4Y1aPgSEyXNbXIzyB0h
JQsojkliXMRcCkUOuOBrnXLGb8RDqKYZGT+cTsOylP6LOWxDQyOlIy7r86ImgTBC
SKXUu1LKyItfJTv9O5WUZTAWJoab8Z7BGpVx2z/zWwBeld7RZIn6OeytahzmUU5m
YQvc4iqo98f9gwbnfWckpJz+mgE1HBxxnA9jMdGGyalzVLk/b4vXTZ1Ue6EOg+W9
GvQmTdfDOJE37f7FgGUnplGCuMr3XuxHnSp4q1ufaT4gTetrBx/KBLbwH8RWvmdA
jNq1YXCvWiusT0m304b1jQU23sDgtChdERM3NX02v7UIGBF72RSQOeGJFKikGFh5
UNh1Hw+oMF8+Pvc/VzPY0hG+atQ29E3fW/zZWtp6XHOaMJeXsvPpBvuemBhQ/u3x
hVPDy8VCJ3Wbn6n+yomNWpTjEMU0hk2fGj5Cj87JuXNPbFKrcbLJ47SGpw/hO3Ct
TcmSZoqWcA9RNTTFAFszuEdnRPrS9oIXAQMgKoLvv2cyWKigcDZ2kFqJlT+LoIlb
XRqJoJVyytlswX9WmdIB86NvCmQ/O5eWSU/lMdje+fIXI+KObLL5QTij1iIXu7DV
9U8dEKVFZuxZBOY4KQgAdQzHP+ZQcI2zH485DZSj7vemdde4XNPN9Os9uwTQXfo7
yieHk9W8yJv6ex+sTe9gochEZ2q3+wXuFaYUc0JtU+mueahWhs5NhWIW4uo2xYMt
KRgmxIPsfOnw/YFKjw5Xi0S0HRh9+ClN5Cxb+FhLrJay7idUmBxdo2cJ44QB0Pcr
CCyXMLNNFwXwR+RciYtRL9yFUF9CU1agn0lh6A2pXzolzJWUDBwuO1+qhTdbtTXx
yTjO2S97tFzUZanxOHyGt9co0CEkaHDZYvxH5GoyDW8t0m5f1kPhEerPdjtV3AQ3
vI7rAokrj7WeBju9Lxmuu2aK2wql1mCV84o9lfe1Y0du+VU74pZVc8SPo9iBQS2u
MFTrkcLUTUxcsnkLifT9N49pJERMYnm6Y07WZlFAp1OfffN14o6Cd9z+/GqXBx65
nL4MTGWaSsu0s8el09ZRW90e8wE7QdG6r4mt83oqHrqcEa8C+hj/6RNc7bwEJg9S
b9dbSG5hZVj1ZSDPw5r3O/5TTRjNKcHQbC3qWj/RB2HaVed235usyvrllDZbds2q
aXGRHGw+Ycdapu7iWnDK8PFGyd4TQu+JiwPXx5haDrKm19q2SOh10cU2SkRHXaeA
eI4MJjFTCVLg2aJajQ5keoGue2q0NhJGzHIF2Jb0GLIncjMJHXX0xLeBZ/DqT9K4
pW+ty46LY6GNMUsssEs64/PJnCjVcd9DzU5aEQWmD44iAc1LOJVCddeIq9UsNWyq
DkudN8J+r96YbqC98QN7oQLGVNvvFLk+Q94bA6gjFKladMy8GgvY1yXZnr/n1qXE
f6ZQMmLFm5n68S63NVdkLAuVEgekrJ5uJjtmkhiYbesGvlqhzvsLKCFzi3K7HrlP
VlQhtWLyg1yJc7tufEMWKge0JCCsuykuP+JHaljSYf5dyamiXXA5ap4n3pMhtAqg
2aPijE6dCc7vQ4Jr5qZtWROwnLPG41EmTBH15vhJWti3/hpC4KLWm9TJcRv5EigQ
Wyg7AKzaPeyTmJZUx/IAMSKjL9vWopxuZADcmbMS8TK2XvoecaQTCvQhOLz+P/7H
keaR995fRbFv6WiJV3sI3Ej2d6DQZtK7xhZfXyOVLJIs9ESsgSLhrcMYlGUVr+Lf
mv7kvBVrsy/NMj88rpaska97melWO2XR96ZUxzjG9qsT4+TwzJhe848U9H4P4VRE
ZNMdnG7l87AQX3mQTGBeM113N1LO/+fYOzdoukOlEL91pgbiSmuBjqYOU9wwE37B
WYkWtsFwYWz5THhg8qc0HUq+z8dbHT3Qlaa9JTIEJup5YRI4PS62XWMd2sdzs87C
Obzkh61Vqw64fogZYZb/Oncq/KpwkeImKH7Cd9NKScKwHNsvbI6zojEdDZtDvGvZ
+70gEU5VEX+9XvnLCqxJpRcFCVt5MOmxwvAKVCdbV8tgVs/TQP85qBeSsEv+hTau
ag7QI+07aq2iNfz1PN3rFabUVWLncEyX3vc1eDyf3OkjoPAQdvNxuOEylqHeM/B2
z96D/Yd2VbOJpkAzE5InTzW9HIvD2amasntWn67+dd2ufYeEmQYj0T/6UZLCpNXR
VgTp24w+DMLZD6SCwFoePFcDjMa9Bch/jGZrzblyEGOAIS/7obEV4vurq/xL8VxX
1fsNhCQjLFNHz13BunKvKuF8ePAaKvWcHbqsvutkIimGjbIV+lhQs+cuXR1edIZk
ERaA9JjTH/bJZFeRChWrf9uZuhtxck5X7Rxf7lmUH5yrGQIpMmp41d7SNQtCjacI
iLkMzgTVDcJBzs/EHmNCvc6a7Hk56H5eMziWMex7lzABaSYVGxgVJzag+go+6XOY
h0vHA/LBYoA/sNZVLzmNtLLq5onn9JsCMftBRNYfETnyYmOvA3d/9YxxWRzzgIk5
hdesnW4gxvgfCPRykvIIlvFAI+uxdl3r27p0BiNWKchBWo7hX+i9W7yHajRHQaUO
ySH6bcSzou98RlyKlw3YNedSkqJypPgKHfZKjjz5mRAhwKUQZRdQjtPkjAYvAZLn
BSZK/4Hr5iWiBRYogwCZ8gCBRSxW+aEVxpx8MjyzeNQvf/rwH2Xli3hbZr7SXFZr
jn+7OnySZLhp3V6fq0zN4y52DtaazTJHrb4RdR8qzjnJxoTY502KM8XRR1v96uXP
iywb9qMiRdMf/kj6QOauLZqm3f6+/8JGkh4arYKHt1cfVPKcY6UXDHKOzFlRy6Pi
qPl+vF0NxFvlS8xIrptgCm4QEL+4NfVmcBD1a5QwsLTedVUdjnyfkr39lA+YfniW
1K3Y6LXFqXFeJ5P/6mzcYxQPUBt9JoUFmgkdOtpEHkP+1HE7KDztkupNrSVAMFzz
pwUuq50WyBUQXHeU5vRPJdZzFLyctxJWpv5RTcNh+MRzX/0xuFvwXPVG+bihlLyZ
A1VhLBdQm7YWML5/d+M8y3Ijk1gjrlEhoI0ZSJuAbz4onllut5z9je1E503e9Uim
koXVknDamAVlL41sf2plDVMVj1MJ9gk48yoR+f36Zdje12D/XqHXYiM+beukxcWF
nzlZKLDEyuKRHHvehMsfMX7u4LWf9cvLM9guxkQVGKJBxTU7Qtl7NAfp32KuQbZp
GmQxBkMqE7Q3cvByxaKv8VrgYPzrLQ/ty+g4VwvC6HxDvTNxcFRlktw0oFe0D1TN
MAP6qKNGQfZKuqVUzVWNsMyeMbwQztdQ3d96+FIRfCRLonukpcOPzoSea1zK+ZJy
GyHiOI1jdxxSqbF0W63NTxS8ulxH72MZjWKW/7LnQDp0mZdp+C6SW9OwXGljE4iy
6ioTVs17fKVM/JIUAee7QviPpHnsUmgpkgWFv+q61JL7KUQkf2lKtYPBf1gN5xMW
8hRLCY/XrID3hpejMUGOQdg7lI7gApe4VglN/JS3djJYka0vgZAud1Iq/3LeyO5D
6AlzER37DrnNvyr5WHzlrVEiJjhwKj4PNCEXKsmh+1qfDnkSn1EBHNb6fjoTU+jz
5oBrHfzMAFtQR7gLXDDDaHIY4yxBlQwQccGN6CITjby7ZzB0IN1GYeDrnv+hv4tI
P9kCAU4uf21kOzh0s2VVq4sa/mso+EtcKzCoPy6SD/7DX1V+aJQRGrg1uisjF1/q
qFQxon3yhZ4tFTDfqMmTeLJGejzWnpFDsOgeV+AUbdJv4UqDMnw6heeJ2vsJdFb6
vRiwEGfL5e9/JtboQoxaI49znZPKJ9ioYfiYqSoQwbEwe82OA/HRJuVOqM5EEvbW
Nt7HrInaXExGh7nOLPDr/4UJKezER2ncZ5nV+u0lKRQcxAa39Aor+d4QOdxuuqhY
AMsza8aVutiuK+JWvxTORcVnGwHAdheJdUFONh/GmJEKqUUEXLNYqAUtkDkE9Y9T
GXzW6BdczxD4nt7QuwGUfC1HqpMP2VMZadlapwsQ7ZTsKnZmzoJh7tfSRZdNZ9zy
X+5BJ4DP/VxZRd1oMRQUluHfz20AxhRJovTSn86j978b/kr69Wb0eLrCM7dtREk4
D/DO/+JMPmzgP8QRFQm64HK9hroVfurRCz7SjCLGJr6dXSnXIiz6jAJh7c2uluZQ
Sg5MAdDdvHOX0Q/08Vp0esXXXT+6bPwnjcWdvhskXKpUU5+nDw3Zu+owcj7LrcTo
WkdcJYEHip8ey3MCVNKUVkz+UZQN3nhQDf5pwbU1DZjQy5atN9hk3fCxEbZWChE7
LlnH9nZT3vCZSsh9Z1yrBQvo5BhDQwynAg23rqWCP/8ovG3ShXuDhG8/fXxP/gaq
JuLoLm/8eaMsUts9Oy5qLpBTcoZ09g4z99TYwTTLXXwlt44tC/fwLkOcXbxNEsNc
70kaJigxKOBRw2vcKNnmHEfvs+D3LvW8bdzc5rNnvFdOU2rEiXlj3Y0pEVxHq2er
zGlYrl8Nm/G+bxPZMWjENCmW4tVL8zqAxMXDFtMAyZQXid4t3no1+VD4hcPumsyN
B2ZfLklDux+/LKiVCMFyZXZeu7dSERB+hqgSbHWyfX7ZAFWeY9V5G0tfjApw685n
3zPYyoEWKUp9+BS1yCniHy0aXSDJZqjbGyvv1nXDxoh06zQJr1YnwEkNUbYJqcSY
Ur6E3jf1P8nqnWC4VCliZLhmgIWn/IeVTtlISQvRZxr/UwwfB3wBth0xlMeoy2Of
gVVLdyR77pl8iutmXqRAM7OYMDYJd6EUYkpn7R6iCcP2EAivpUy2+y1lYkAd1U0p
2gY0iVXjDuzS/KwLgyut+lJ5iq2U5iic0ENYpA/+w1pKTRIEhZnseUMQQDdEirES
VVEbiJptNYo0ikF/mgas+VynY6dq7JjR/r85D8OF6XZj2eozkOpqw4L2KPgyWkS3
xH4UXjaJ+3GlNFnVnMDT4mvGwAai02vc+VYKMFoGQQj96S+HLbFLE7WqJQwCf+sH
XWOhvWVPfT9KvMeYrUWnHGsgEwmWoax/PTu1VPqle3ZqgM2PRizGuVYtQmCoAdIm
fk+tO4EoWn8d/X6FOz6onUArOh03suCXe5c3XflSyHGN9IDIXW0bvw0zFEhMQ82+
6splnGEwbf67i/npLYmEPDdl7YOUYkd9yOoM4DZITlT1Nk7x7VKv8lbGokzIv61O
lpKeQMmOyl1gCYh7cztBRQcL8Zolgu7YB8SW/UkTJ6b3cTSVBnNgWaw804CmTWlj
gyczgnaLEFlY3dlD7azYJTQCuroViNrSBhH6R+6NzK+MWUAoCAvH7RXJVBCWJls3
iVeeFFn68reVLrb3UzYZWCgZ1047uqXeVz14e/z8GgP9de1Jg7s2JAKaB+PXhwHR
ZOVhBakl3cBff7sA3oa/rLgi4AfE5JxfVDkf+EOm7s3hyLQpqkvzNC15YMuIA9kA
lXf2WfMeoNfoKC3Bfg0TvdRALFqnLGpHz3nANLQPvpd0/y39gnbL9c9mjmOAnCAx
/z0hdB0rPnVvID3E6+B9xyddxCLuolADAvgdJJ002hZgqDd7U6BrufVcuRANnlYl
tn75N+6+vB8v9Um4kOA1uwdphowrcIvgC9wdaFGh2mLwcRt0Fj7Yq19ozBcxMEw6
b6lAe5BmHZTs0gG8wPGJMT+5pPy8yeH12vS8UQN2OOkW1SAIRpr900xIVmoDQlED
8T6lNPresi4W2D2lasGvYLg9l5bhC3Az74fV3Z0VEtEn/zmAyqEz0dZw4FF+M4jR
zNG1P1WVJgwWWfV6W81y5czNg48aQkh0l3n94gF5VH804o0hGXwn5PhKOLWdl7TD
9LMBdpAoiAcuO2FgfK6nqsTNNatZCUchMBo2ATXNF0S+OJuHuCn78KMjKwzzEtbk
WjiqNQBkfQeVrJJRM7MRieZBNbUutA7X11W/yy6DxPL/AZOT0QP+QI/peZ6eVmX8
YbKbgVmA+PVWnFs21kTrCleabWTge8FyG/SH7ddKfTQDr2x2+6Uob6VsJOAHWM8k
EVv0B+MMTTtTXqg2XiuNbBCuFG/YYAGOczE0wrIelhvpJaMozF3jFRGMdLbZye7v
aCl4zHyXvOP2Hr9IonCvJvPgdelgsADKrA4XufDvx65nwOiRixHnMegilDk83Yk+
H2qlxgf9bojH0KqBnFN0oUTr3UnzEyYBXfcYRKC6UAVKXpzjsU49ntrRxGtIwxpm
FEv4ssM0EiK4LQEcClX85Yrfj19X8j/eZJyTDdwuoxmSzF1myLHYLdJ3Ms5LoAua
uqAx7ELWbP84HouaQ05pvHL1GvFHD1rBWrsciaIbhlsZQRyZZO5iFWFFb9ay/6vI
ITHfqskgWaWB1M1o7FOPhZ4FNoSg14Q66qCDlj7Fq0U7SFZyAXAJqxaf9UWy5nCF
MZT4Zz3xct/a1M/K8vy/rcQMzrGt8PewjV0GoXrDpbEmvYLIGS24CXqgPRRhgyk3
bNCS3HJyri3PHXVakZ75sU8xXmkA/YoHTn3PrYeYSQZQCL/WVOGiSUkx4cniR53N
rC23BL1kmWlKyioeDUhkA/VnuZRXMnXUk8u9+OpToW6aUtA2WVbmDYF9YY/7szry
NkEmWv/gysf+Au3dJrDWsEQ9d7e9PbjnLEnYWj5+ufH1xKIarV4ZscpGaNFAZ9KW
D/t61vyQlMORDEzNN5ISxvBPNovgMEu0Eh1aSbuegfug8pyD7AJr02dqyor2GBVP
w91M//28t27CyzFocmxRiTu8qPa9lyoVnb76zyRV6re+x1FpMjgn0rf+v1M4Y8Sl
ZopSLHOiBP+fHv6AsHtYZhziCwQPkmgTfn2S5ITQIOY2BL/QMaVj5ZtOpbqpxKml
JeUZ/ypNIRwUaqjIkvtUfJ2hJg04FrhD2e6kD5i7YVafUqWVdQY5lsZ0X9R8QB8I
6CFUSF8tEWaL3Ff4JY2uKpxiWkUKQw7IVSh2+fVOhqIfENyWVCYxIobbpsrCZbqx
oIA9V9StfPzExKDAxdpKGtdh69If1jeZF3luhHp0CQPT/2I/ZFx2IWOinv5WUGVm
/virmynJDBBJhhpW29GtM0GGceroidJ+Jz/hboWJwsFhZPFMcdF7387iu0EZofwQ
meXXlzylS/3WC6HK38VbItIwtfpwIrzp3PYkpfNdRKEiWqARLYNqPTJKe4s5Vf0m
uP0lEMXRuD747eABlaGu4ggfPnWbTbRtq7kCIplzEdfEqB4U6uyJDRR0LenxvLi0
R6fvvmC+354dZBIXe8YpHL2aNbZIHQipCL4w5ZW8Tu71SkiAHz6MfKnXvCgmTgnc
mY0wH0KxF7wTF+3LAZ6t3Z7203QfB4QqpXHjUZzLTQS9MyEHOATjBCWb42q5Sd/9
NJ6+Loy7OVApMIxFhWJBpT78HDh2jNjh/x0Sn9+q4UkoTDhFyebYxa3ECl65Iako
JDifHqcbwDPYlzwT/Bgrrzh6bvbGJ4xn/IWPl4GSGBZs7csHE/kXpOmbJDsvwznC
d2KuVM3AoQZjRdOKAxuxGK551mXxOFz+j0AffGhUGYdv74Ve68F3SPgCsB8YApeg
iBdb+rqIsRmcKvsGb/VLVI5nIJ2NRjrAWzJtrSD+2J++aYnMvPpgBcBuJBYO0Xow
zzgTrgA7kYY2FuHQAxvOgkksr/UQ8do6OmFKMp55+JbZCrhgM8mYWIGU6KJVNx9I
uzFpOuGf3p7g2wMH/DDJUqteK9fQCYHCMMmRmCJNJ6uVsjfSNWS8t6+tGUkIO8/G
3esx6BVnTLwcu0RdrFr1cHRvPK5O2nU6D7jbjAXXKnzHxVF6WBCWNSkpR5t7VVTj
S8GflezJRraotGcoEm50y7Js9p7X0W/eteOAbVgordHM3kclorOrtH97gFfeO9rj
A08BvMVa9qSqiZShJVovFjGLb0+wog1wV6ROKLqW/yoBJ4HMo3HCqhyIyCz5RiCR
eRuMl8szQsLRf4UbwcHs4rAY+iTeg8FIF/yLfXtHrejVsyT/pBAaWJn3hbjhbnz5
tcNroUxxKK1b3cSWyv78T9PuQSN4pSDrVMNwkb7mBDHNH7gIHcxuh93+hIp+BcxR
OnMNGhBQCEcg7ZEHSI/A/U6yl2wLa6/QPzIL5fdZVNg/hY4XwPTUYYJenviMXc+k
YrWxWtCC7HWLzBa7JFKLD+1rJ4c8ITnh8zJxUTVnlY4KEje7rIed1JdY5DcKcLZq
kBNxfbOvA9N2Lr5yITKiNDmMWYGrzK8m8nkfC+s1gOqjM+9LvngEB4tallW7yRG0
tlj1jJqgvjy/8NZbNGpny1dDfUT4xvuC/A4JV0ik0ttFlTTtSSeNVR91h5iYAVlp
k7SrXIp4TgsZEwZhShLDAl/pbWOmJBDgJ5fLVOKAiQCY9Hsy0ejVQ5YButnYvMPi
fmDumeX2CcFD9oZvmFoRlFoZ0acWGnrtwnIpwiCol/WperG8OWumWOQpucZyN2Fb
jZgz4KFUHaJMlUuulYD3ExdA77Vf72+/ReE+XWClgvv3wdtwC0OmxhyVmkA+O64U
NKVjFjXPLPan4QjM50IznQBdNC64FVcEXzMWgvbDB9LPqflTHGkdHD6znrubsuso
/J5fT6zVF2hqORVkB7cWkH8j4gTekKOEAUq/wadiVW56SqVHpWrGs6cdWPYkXSxQ
6G4zykpySDziU1e+tICAINU6NDhCE4QRaSBM+Vas/HM3wS4U3EcZGuzT/IkMkTOn
tgitnA7bWlY0XkoIZ15YotPhbwxx71WyF8d/Yav23l+h8wLHqVnqsME1Hytpog9u
Q7Fa9VLI8yrDNGK3GaRE9ulSG5spnqqF8xCBc0IPEBWfSclx1/OWF6JeCcv7cq5m
c/iVLoipcIjmZNJtBOzMcPMXXr706v2PeXCKEg8ZMndipg3ZiIK8tMQNBOfSUQ78
sTBffgpUZ6/eLCEgqhjMsasEIFORlnd5kGlOR4/N7oNxqojFvMkaduadrBSdnbHE
wT7MavKajeg3hLI9fIl7oLjGYrG6gIooeQGb7tkv5cBsdGu/uXqh7jKQjbQKieRu
n6a9AfOIQsCkA8ZA4VAh3kdJdEb/fVGz5hSREt9Z/rSMJe1ED5IghivHz0nn7li5
1nm23UqBxM9sTjzOl1mo7m5mmCB40Y2yxv+kkE+b6DCVRerpmzVVT+nO53z9pt73
cpqeXuDMh5OsoM+zG76R9xnpcV3qEmO6jLmbcHDCIJVLFFiBc2HxBFYtFfDBPOMH
v0xG6r1EBXFBgAzgDoLJKKR12l00of4QuoAsE9hAyVfE7PP+AqOUvN0ZYuI4QjyN
jbuZpcXHFgch+T8BDgfi3yl4XIq8QOAGjfw9CsCaEY8Q6kwRm5IJHBA+JUgFEWYq
0qVxE3rT9U1zwfvcBhXWTdK1Qgej6bvQzIgEG4ILFbm49GQYf9FYp1SThljeCA6M
XpyYQRtqlOddBBiQPXTmv3XGRt+AYz0Up50PhY/B8IGCw6PqMLKeo+jsV6hXTpe8
TDqucrgUPm0xEPoycyw5XESRxyDNH/1Zv/o8GVVVcAHPrucW706cTeZ7QQEi42fe
KOld2DvGsCSfOR83xBdIuSWNOjrhtv7m19Aw9lNMRo7ZKb+k+J5wNET6QnDOm4UA
eD9o5kKsP/Qa4wZhbzrnjMWSOWHhl6ZWxIlxFKqLRq7QeSoUHPwC43R7c/3etlbi
6sLtlF2IpZFoRXXKT2ypjIn6ZHsVCHtRGwBUENkga7QYtx+3Dr/AJb5Rzt81CnZr
9IKkdmCkQU/PqEHUharK0l+TnhccQ0tXrI4Zh98yDqGxinYxpR7LIgJlPc5QBvwK
I6fJdLyAPICdCRaPmJC+rCZqbcR4Cg1bHpKYNrENQOJ6mDPiiuZVp1tMvWlBubbZ
2HKPSrjEOCyCR40ENzClHWn2Mpqa4uZ80S1/OPK6P6oMWifcLJzps12QAPP7eP9w
4yXZL01vq/hG5lUPIt5oNEjFYpJoivIi4V1XAlWFJ3mSU25N4oaqCpqyuDfP1vvI
goep02mI1D/ST0PE3zK3NnHzu1YNwT6WsXFJ6BcNMoujBReR0yUiZWK/iG+sfhaA
yKSlQfHCKxy0StWNM2NvqkOXhTMAPGL1UyJeeN0DDlz9uKOy3U/QNTWRzOUOwiWH
dB0VzGhv+xuVnacCY7KdAOKjtcAEEGiHVjILKEFT7eQSKFxSZjn4Z7LmUcN7RSu7
6op3EPiu2weKGRn5G4ZiniOf5/+tafOyfaXUg2dAxd6BRQjBweinTUdxQhhXC77G
8QRY7l5oahhDxjytANaQs6ZKhOYWzyIu3pyXKBKsFF46lgzZD7xLH6prwUnkPUp2
EbACf88CU28zcFBJ2qX6/70mfUPiuBqFzvyBUWF0nKRrhofVrTZr5apk76vt0qYg
Yw/G9BFbI34qu7K2avLiTxJYst/bVOwmwWkdLPC5ilqbXto6yoW1J/jtxxj9e798
Bk+4isFeaijIgyDpqixhidswi661ELVUEnwEF3nnK9xToclHAxWWos+tLVldu1NS
Wp27DC2N0W8Yj0ObTt5ymHAUbabg3g9pRH/rCD0AtJTasZN7ktN6xMdHcul2qGHQ
J2vtHERt8YTIz0mMe/Gsf5ZcY6H84/ZtPUNbMzHTCAv3j/pMqOSlQr5Tj6Tp2Qwl
Vp6ln4H/2N/UvwQ2v8iv9SA37FLVqaoapKyGP4d65GOlI0bvQ5M2N08QIamy8Kwi
hKNd6HGP2hODCjBM5IE5qUvqzabIBG63LWhW1OgQq6xV8EZyXSDSsUWQzCjxUo1v
kldHWdWI86c+7e6m5g65PUDobZo7k959RsJCfdgfnksaUkAscN7jD5X8bHXMEaJT
/yKJhpo4nPky0PB7TwkVM19nqjA+Fp99+p9HQwcR0oxfTHn750liRasBE7lGtXpM
HKdabpi3tMQutgcvntg5VAEuAadboqZ+VX2BFGyyF5oC0X1Uo3XByAF0MgJPoHty
4fAw1QKNcZVC2EdFPuzBglqnxyyuhG2/6P8cPiRvrHOnrpFWORhbU1jOBIvB/HkO
d7wQ12pl5+MJg3hL8DWxkyrE+lvVw2H6I5F7sGenK2o94ob3aKw+yVPD6D4g9l59
5yjm6eWIsx9mwxxDP9aXca3Ubi6FRYJ/f7hbpQYspAzmMJZTlHgC13peesTLUmpb
4NEai0el05G6shx8l+T4l1fJO1uhtPeh1DxB94v2DdsvRpscyPsdJsrKUPR5bgPk
x2oXnouxm5Zr+jya2RabeOePX1eZvF1Z05z4VwmQq1m9rz5ws4pw2Oq1dZT4h8Ia
2Ro7GJw6/VKsneZzw/Jvk70oLdJJkxszvLIiFfXVkjpFBTqB9+E1qyW++NaiWg9Y
1vQqMc1i8qBA/Ytt+EMP6+BFc4LkZrQVuLpY59+ofKdESjK3zMHeGSUDWlWOLJSh
a9dizueLguNzO8FdzkXE8OKCf0dt0XpatAalMyOVMrZVd8VUAqQJVAvQ6t9Enm90
lyg5rKuU0GZUt4F6d8hYRsqIqlAhGCeVWwNq6EbwFDpivXW0A54UvxKf6Qs48X71
66RIhAwaK7ueFSRewzvIxEUGtrSC2mMdW2pzSQadccailJrK/4N+maHfc5YZmtAW
f1Jlbz0Vgs11TVm8qz9CMuTIvKWQeDHfNeZ6VGdfDU3Mbd6Mkwvv1jTskcNIBs+X
3nyetWTLDWsd/72WkAAqS06vIaBh/qXCyojOMyAvirFi4g/TDc8g9cRv3tMGjeTD
OgBMMY2xih/7vL/McQlLZZv+5vz2uWq+xkX9tvwshxaL+ZmCycBXfqzcDIyssjli
E48rKk03Kx7kd/7FPwUtRr/BD41RNJBfe/IT25VGxKavdBA5MzYSlpMgzxTV0sXL
3VoxtZl3XZiJj7xNp27biptoFbWAovrJgQSTmmlHSuVoxa4GhnuybJMe4P5M/q3Z
Kuey2S2isxQ3jJovWVf5Z7JD2u/IFmBNzvDQQbIkdgjmO7AyDTa0s8Jq7xuq5CSe
fDNqvYlXADKhunBQDglFJ8IhjyGZ0Gwnyhh/kFKYQlTsi2pF48RG+5QIHxAUntdr
RQ33OXg1v5vscVQCTb8SvAGX4imnNSd5LifM5jNelN6xbvLyJoKDjxMo5hNa5ggm
dWG64diuhaCPwAYff3g+3ThFHkM8Utpg5dQrb/JnMT+PhkfJ/JrYiJKvkIsoSf7Z
MY76pVRI/SI+OxM5AOXKPFGjEyz1QNn/Z29uQBWd11Vbtsk84ODMr8+2KppcEDX7
JqvQ1TktPiNT7OM9qiUkDQWk2BSxr0YGh6E4TsbB4PRBCxaHY5mC40tFmM8zhGDK
sdWLAFxMKmk7kyqhg/++hxjLAUzMIgcG+Ks1FyXb9QYUQyxf3SlQNuNeyZVnqgmc
EdqH4zafmfxevCBBvuw70QG8FlstrEMGm3QUdofJGvKlsU3sx/487NLks56piuPd
qDcoTXvhP8RfPRVZ03gCMsPQT1MYfmxepw+rfMLotFUFHyfEdQNog/Ip8htVAdsl
yLLqvX0rtT80qJcyDPv1RojejTKrcxFMQCGA+S/MQlH+vEhnE5aqhOpVS6qQTz9M
lsfbVd9QlhCRpDyRJSY1D+dMOSc069k1mNWlVOMfsAIgP7zSnWdc3oCFwilbVNtz
Rl8xLaXj3CbZkCWPozpTRJLCvKtUkZqgVDFEuielZXgwZruDSbrSTf1VWOyE6gTX
oBerf4u1rjb9b/Grg+z47UTCC5odKx6LiN/33Ks8q09P0TsCEEGDYAbQovF/nOT/
HRsgD/Cn/FTuxRXrQBBJrKukpom0hprQJQ8PyD8taZgeuoqbsHAifANritZhDWHZ
9WgdxWUsf8s+S294NrUq7GdqbZOxe+D+0F5dSHhxzDa9vlH5QMgBoEBJyC88bbRC
QIT/K2G7tZE4MkEO94CRYLTc47s8KrB/ugHb09CJeq9Y7deFNNMFc0EUNnX2FPjH
M8Q1Bh7kVS/TQqTSSdjDlvUj27rcTpodPvmthxkpojAp6we7PolhwglkFi41bEBu
CuvhtQLtHCSMusK6diZUdJHn004m0T9whbJAfills/Cf7F02i+l7kX3yv44FtYaS
HomMcT+MOapgXhdQD9oCS+9Kzrb4pFtd1J7TuKoAYbkmrUtObNdGlqp3Np8paPl8
ph0xndZCJ548lWx5HsCMonYgTc196Pb9wQPejjO/51gRVPjKUijJ6xaR1sxwMFlf
elF92qO33+EMbSF4P9Ypk5tJjAK+SKwDnHZhkFmYSLr0WH7KqFIh4VzOYR4/8Mu6
b4LRHcsbedyoEqU02NSz88ru+7BJ6L9DXeKS2D4eMUy858UJirs0cbjmRAekCJSf
0Q3JaFMZMxxFJVG6GQ01Hw1GKTuZsgrK90u63mA1Mt43zlbzKbN7Q7jttVIQDWWY
BR39O8HhbhKugnxneSVT3pnGmQgXE0aV6S1nkmbvGBpATeXWtAZHfTetNNL1FBj4
EDs/fplbwQyPvYzxjb9JDpsnjLCtw010185RyJW8HAjhuUYyJEtETXSS119us/QA
jcaTCq9c0dyXX84SqZMW5PD1SFDpQur9eGb85QwEXGyzIepMzOtzcsi74dnFBZIh
nKaOvou61XuWUOtb1Q2U+otA5BrtK6zCTEiBupo3prpdV5IfESzb600BhGyE+12a
rWZq2qgCJ/akQerM31k6sE/A65rKSBH61KVMaLT6D6ZqNcNis/rLh3m6yQvoQecx
cDeVlhplCua8AoS8lGaw3lIvQkdNJnZgrv/JgkASyVfjiIaEgL9GpYAvSiTkjc4r
2cXudahh0Elh88NsvfEnKx5SdK4irsrigj7Oh6AQnDdh/gwY6T1PypJM2YzYuGND
LWddgX0wDJUYPZUM0DCZ4boGNpvObXm3nuVv84SIthSy6Q2Qw1ihJoOJgozPQCUs
HLG3pjVRg14de4gJz7U3nijj71gwpcGaOBzkRsp84RfzaCIkgBCBHR6MajSbiwm/
CiUd0NCdd5iOI/hiKNl3P0KxH5Mm2KwT3f0uqZg4xrn81b1jggUJFTDegcSZdWi6
hLhKi4Gcnh1sasFIROSsk/HM23+USKFeLJNcyMdmZphHlSUIquCCAWAL8y4elFVO
caW1qh4DKiCw7NS9Rd9WLKs+jTONOF4NN2jQGoj3DT4c1yR8SSItcFWnoC0cpNrX
cCA360bi0exbWR+6J9qh9lJJNPRAHZSe3/ZyowvcTg7gLgHK2CsT3P6adDJlynva
Tb62N8jxClfTzGi8tU3Pjlc/7U1fRP4ekEFGH4YGu29gMSndH48sG1QT7b9Vgzct
RRqep1NWahzYbrcBVUcRamqSooEDjSwlo8OXi6R34AnG4v8800AeVUFtox7nDvMG
JDJkalNIISDeUDHWwLKGIi1vgFI29kKrm4Qvetp8rhTqoik6KVjPh+R9d5sR9Ip2
nHP0oa9go4bAEIMteWrdskGA/qyGe/cbKWRAsj+fP/DWwnirqB8hT4Jn8F2bkxT3
tI8syeyaSE8PXhxo/JmB4eF21xw09/p7mZVSOcKCAFjXITM3TcTbd14XWgkrppjZ
gRsWehLbiD6f6jYcFtGeRU8pNetFYuedlII6VcexHoS0bujqjQOJyJv/wsk+lKnt
OcSnKXOULXStM0ZNuPLahC+jExXIvRdK33oMq6yBApjU0thVGMZoz1GqOwZeGMOi
2vmXmwyjFz1Zs9G+MzsLFvEq6lBjD3PveUmlnaWtK8AWaSXUjJ4YswPFO5X1rsZq
0sGt9qPnxHhsf4FzLnToPNv8EQH38v9hCS6deYhh367/xYT56EVF50z5Ujx3FHxy
XuvM2QNbbdFdegkzR5h7rasvd79P7W7OkaVspWP0Uxy8Wt2q38vCYe4fl5oyJDJ4
P7v5mJVJk0dWnhYFQLBRD6Eg0nT2PhveVygdz4s9uCOFnfEPhJCyM9D0P4lBGubu
w1lregyN/R9keRGx0BxewLvPWKVkkWWl2N3ei9cCQSSkxFx+4Wz0/t4fL90ClAmj
0RKBmu8i49+mOkYEebUeLm5oyDRTFF7SDGVeoqO+Q50/okEtXJ0mAoTNP0jXMIF3
D6uE42mRtvw8VRzgIvBMvkZdnF/wqDVWTuvbUsO5btTuvNpHGGrEI+GWeMpKqTQW
aIyBZQYxHhb2vtMJjiR63TgxkPKHVXfhUbuNapDJkDPxM3t3OcblBNz+6wrpCJ+2
7BVYGzR5GyA0mPIJ1fgzuXzr7YSzpSoFJA+D+b3iVAH4pmn/jGmqa7KcXH8hWMYA
dfGahYTbuSLIq3J5kjeZWYszMVv+zFzFQPsuBqIAE22pDnfJu6/bYzCPpeM6QmSp
ECxsAA5Uf5f7Noox2+tevQpDUwBQkjKR2Akqvfz0p/wGaaJYNvSBTkv4+MPWFdhE
YAZ/sin8178+Mvc/TQ728Asok991lpt1gGWmTywWAto1PkKFpwhX0WYXec5lpDFI
xicK69PqwVDCI80VJwLaUTl335D1sWuxBTC0mmZeYoL6u/sxFzOKceJ0tkfsAc9i
04BHO3Z3OIBbUE91K88geq9o/lRBHLUFjVGG/IHhkfd1o3XxNK2JMM0TylwXBNhG
tDuXl7ADuON53ecHN7FM+vLALiYsbxDrewKTZrOcp2f4Xv9DjVaqxdxuRWnxJ/gN
C2zxaIesXMyl5ZPu+7+IQC3QIYIeGfszveM3R1R6MMh4wELtsKCzfPNFYTdAHuHz
mQY+6npLKUMHHJmOAHjFQSPFELJkv5HC1EvEmn6ZRwXEZxLaKYbH28oPqsdLb3oO
BLDirj9JHM5edQClWVijV8boY2clAcCzBzbv+OKiX4SkO8tMbzxMTeAjZOkVbE9L
/TYYP3rpdVIRs3Y1t62R0I2u0ad0hkgPjqzPBcJ4QP3dcPx2HmJkRvxPWHfFR/lg
EE/f35G7xXus8XsKOqrunEsA+5kapocgT630BgsZ+HrWeUn1A9xTmgm26Hmwf47f
fEvngHf5LrgAZi/qX+csTHemgfcOlUyQ2VYSUJA9KSMpC03vX79Nge9334E0MAN6
wRoZ21XEzUb0b4SCFUvWQvVVqvjku1Hx6XKgmi4bQuWKKlvpmQxao3YI0TUk3v46
nx6K5ocPvawwDDvMtpRqw7k3VZbRwQOUV43RwcIzeofQkdc7cNhi/PYelbGGO/ec
f2pR4im2CYP1qhMDJ/Mm4z5P7/jCFa6cw8co552vqrPkJ5T90rZdl+QyaKP9Noge
7YmGCysJWTmNxVirDDxpGkyKlSkgBgqSHjaAbOsZHSyXTopFb5N0imChAI3Iflfo
SFcB1dx3WBBavqmdIjZzypzdMOTs6lOod93s47FNqnHpHn2SZgW3emml+y0VZkaZ
qwTDzY4OMDO8Bk/rZ9ljqPQKvJDl8P81X3/7sbOhJdEhBcY4n2vmkbJrybYaR+nO
F28dE0hJtYJymuM2wev7/uYmRfSACKJpWhmX1+2K5bMTuFl1eDiK82utP/aYwyxe
XsesvBJxX4I8KvVuaMrC2xcbQ9aiCdM8g1QMxzv9Zc4nAXbvlZsXyt82q5KyZM58
pTvEiXcbNV+tqOQZGp3sdjMyvXu3E7JntlRFB/NfVV9oULWgEL7F2AxuBcSsr+sE
iY1detUqbLnNZ2BWiKL2u2PZzIGD9nI7HpnXLS8H3+WoUZAb9wiI5onV4C6I1FgH
3vxKjNjFCfbp/cZf65pTudXrAV3SSSn4MV1GwUv9g5gOUuspALLTCr4F4Reqb0Qp
ae1e4HnsuLfzVFR7dtApEmvKpMaC2YxokyEw6qQYbcfnIwiTcUVmVsWbexS9Dm0D
xecEe+O4jdRRMnWa+FARJL/FIC4yp8+jn/EZat5chrWbysd//lWOJQ3qNlQmU7t9
68oL3a4cC8+E2a06pKwIrYidSu5VlOzfWnoeQWwpkAIsxfbZDVooh4HhBxtw0LGo
z3j/wb3aECOOZcNVCzoTP+emHjZVe8dyHUrSnLgTYXnxzPamVQTShyj0hnx+xrMB
0UZNDwvS2Tth7s7zZSvlUFgFILX9/kZ0a2k+ErO5RDRIgMmMshB+hhJkUllH8JXQ
texQ002qu0RiPmypWbiAGq2uC6hQUDk0a6mnOPmOkeRDbBI9Uvm89GIJZINDAALV
T5ppefVjciHElpOkjxHg4uC41zwoaq4LL/TXJaDz8ojhuJKe5xSVN9ijjcJiW6lk
uFlqVrjQsgRLczo70Ho3jYuq6sDdvfT+GQphGwm/1krtuHaYvfYf2JFrsoeULlVQ
j2a2FscIyqZj/hhY4NsbEAzAGF0Sr28cO3O9gM1MbphIiRUJtO298TpSp2xig8OH
3prMJqBdz4jk8RiYBSENOPfC1kjgFBxgz+29ykUX6po4OlhpiXenVV3wOW4RO8ds
dgWj6KKZEnH4Ee+6NrgI3m1rj01H5AiOPOij2mPHhJluvOZ4IuODQYq8TjD0QZxk
Y8JuLgrDrab5frMRTdVtutXkj9i1V6+PCTRwP0SqugDk0Ngi9jOTMX+0b67pGye3
FdfFY029291kOOf8ETtTsD6ZSnWXG8bOGHqsStjTA1uyqgNDvZ5o2DryFyDtJNA2
Rmp7aKFjDUsGPLTlcpyceGtdRZH0Fdn26owhMAS+nM3jJBz5wAgLrYIbTnSolJNL
M5v3DyEztKe6OZp8230Xf7pnzKwDgX6lqdqW9wNDXVD9mBF5nZ7WOR+Nhjr01EV7
wxYKDXT9W37IbCNgB+EnFiyiw9Dmw6rWuCIy2KC+519RMN/4qmWPRTH4Dh27B6Wb
Qrvu2wqL2CkKSbO5pTK04/+PZE59ZF/8ghAOzrv8XLqDXpzjYOWpc2vT+URQNx20
U/1xPc3zmX3s1DUcYrB2JTo5Lz1Ge57biJ1GkdRIDpnX+Ikp3Oxui5qrUkDYnatk
KcpiMXJjo+Rf782YU+tlIEgmVZOtYazWdCT0aI1UWH15fBr2c+2LpwifM8YzCNg0
eRIuQmLoG9ledx5w6kWp+5ae7OESYaN3txveTcDiFfYnzbe3yfIKR+LOXHasY+sC
N6pW03pS4sDE/uSdYrdQsE8ahJvD3u90qaUUdzGwfi3P4Qp8rGWyDf2aEV+qeAt1
zjHBl1pMMDvxXWcYzAyIRwJH29VF9+t85hudO7zAn+ypFh8vSbsNMvu5LMdhnuSw
0QMkTb1yLkaKDNDcfY5R4HnVTmnyebxpWgFtFSbY+J6HZFlDUItn6GOufAEYnlqK
T4u5PfWcq+9CKx8JMbBHvFGNrNr3LgcpXYewctf53z11O2WGm0zgJWJdLr9Cpifx
IJYVLteyZozveshsD79D805/xXcNqglJOag7e0RVKKPRNIYYd9njrO0jsR4T710w
UGRYRKudlwArm9z/auAT2nAPIb4AbIpQaKwlUQgdqIJl1H5srsPjoeL0HyupmbXP
hwfFylxjW6+NV21yvNSMwk27Zb8gaaP+e7m7SYjNSQ5cVsGXMTDVPFdDHfFpGqrp
GEl99YoVS+07nT0K5GZuIDA+YnECzhK/yWuYkKQpeT+mFLqWUpmS6mTBbTbRWbpt
fQPfESFXpBy7HObiYp8Vrj05qBfg4M0w8QYIjGgDdJqGQnjLHaXjj/Ptro91Dbv/
CqWZ8Gh06Jp9osxLLUw9CqkYQPKmGdzhprwZtLpsDk0nFji4ZyWF8jJEVPB1bCNx
tlPhTEGuWX1xByHaa7IRu3/cCuv740Dpy92VAOv5d7O8roa6LbRsL6Hf8q5mkn5+
HaourbbAvmDdE/ld+vEIEwFZ2k3Tlxc3eB6TRUcAa/lJu6nQj2a1lb36mRWnb6Ux
rKtESAeOCcpI3tF/wZ+raPNaBcRE6P+qOthurJNlDf8Dc+EEGUAsLoAfPjJ9pcDe
qVJSWGRgf7gmHfWYp0+ly1Z2fj9snSA1zpRFAI3KNTagVKBveu2DiEOyMc8HMb/s
WcveuNUGVhXP3szk6So00Hq5FIGbkbWMG2y4nqYxcCQ9Z2UFNV6SnmYyPXr0b5pb
sSCLwN4aJhD3Wxzu/JFUjofV1e/VQzEe3fPIxm93IfO9z7+IMsutrzimnY0NK4iZ
g5JQfm5Eowu7pngiskNCaDXZFx+vnDTzG4BRmq+vxM1KfQwxarAPe4Xh7NaiThhZ
uG/0afbYfvWKv6utJ84r1d09zaOh0giLZYPG6gUuev03fv0nM++kW3BnxoMWQpBM
aRa2qk2N8R2FuWw3yYNG1w8JTwtY3enBWLI3hDwxQ4UU315YaCrbOi2yB3xLEmnk
EWLryWeB5qicO/hFojB2vaKWUF2MS3SQErWsW0pPGwY6FZ0MSeJ5pdinD5czDJcT
zYpWcbKlCR6PLoMNaNTgauOdItYlLCEXe0xAK5RuhrSmZbuCG1Pj3LgxfjYtKbwj
FTip9NcfwVhjwecGLa+70vDnWrHJ5RThhwQf9gPsDYJiH0ewUtJmcQGHRCLScEgs
8PBVkgctVGdQ4nnZ6//rm9tUyA84yqOQvBVZu5JGwYuyGYcv6LrvJbAapfoDtxLR
tY2NP0m/pU1rOsv4MKnD+MdVT2VEf/xop7Z43v5mje7X3zwtYSgQ5Vls7ppLhCgs
FTFAFHGt1DyNve1OCNxT+9n9yw2VT37VX0ViZPa42QqDnVSqve/k/S1ol/mBI6d4
lDGtNDOD0Qe6s/3tuM/yo/ImZqORnGk2u+zwNvULoGraa8pgN1cuKDxZMNYw59Df
65j4LNxXqN58C2GAODEs+utIRkCAZuQvOzzJbvrZkyfQc8X74j3aEXqoLNK9cU+S
kBf0Fi0vrZwp2d7x7uy95LPNzfcXbJJoZsYW03IO6xcEE2XdFLPBa9KWFUy0hLhG
M6K+wZWjddVB9ocMD/4RHCq9a7PTrg3hnQKSglrS3vj+xgbi0WLbxVGrOcH+veeZ
5uCYN2GIikRl5GD9Mgjl/lqCtvSpOOyvz+ne/leuRPWAtSYGfv8bZNyCgwx+Tom4
ata2Wk/rikfMmWLvJw0arK/RZ9JzhatLbgVYYuR9SoPvaREHlxHO+zOQMfWUO77z
zXUfONT8Jhw+AAR1f0cqE1LpQ9BxMKQcIXxgtSZYGKAwHvEcRxjgzO+Cns+qsmMX
/+kyn1sPtSrBL/1DYwZ3EF+wbVjTKS6OkVxDY/mW3uiNQYzmQ4+EDBDeLTh8Mod8
g0ULzMUZ80CLPngViRoi/GlXrohKrcogWuaq4w9aXDImY5NnODRlKtfJ1mi4xtXL
eTNII8jmmHiUZrUZca2km9e2ZZ5mYpek8/eeD5EVGmEPdT0i7nBcvecmWPviWXD/
FtJo/QjC0t+5TyhB8cQf5UxFUqzJqCWt6ZEL0eM5ILbWqkO0dzFhHb2hyUXnR0oK
M/naZ1303Koa9cDEYMSUcsBisqSahG11VH03xUoBKM6bn/CnRk2iu5lI9xsVUVKg
0UEL3eXdJxoUzPaTvmv097PcaNAP09Yj2dSQdHNLPDov+p0ibfyN0KfVIEfkurqA
WZvRhe8WEI+vC79BFmYdfv1lBxRLkpeTagvfQ3I84NZBz+lIyGWYoSjQEQOVqZYp
WsvaS5nSlfV/qFTKvX+UjP8C9jj9AUEBTZMxyRfLpGxS2H45AN8gQOetySJVaAZR
PER6Y9WAQWsJmoNAER73teagmEcp7sPE+9BHoCxnjG8q/gg0gatxs/0/mfEndMol
M/03QVOfOr4w4bJMoHE1m0yAZsy1YfgL7ZOSIR0CQcb4MD6kvCROzVnrx5BHsQQ8
Aqg1NJpPO34IFAfNDzlkxECTapbd/XdnMYypIOMpQBdTyMLqmeLs9739jcqkmMRB
/RilivwQ5rt0RvFdC6q/RbDlyF7TX5xrpDHuAVhX1AuTWM4kluewqMGMPDfK0+zd
cwHio+q9x/F2TfU0dvtXXGLykD7ILG9u64tkuJnG7JEoCPO0OKzOi9rLJtdjeaQS
8ZqlpTdGnyECEAn4iJ9pi2Kapbx1x39IsgYn02g0CJTLT20TkIWMJ6dVPap50xeD
09dtawCASYNvYyFqTWKEuZRwx/IyMPZ/4C97Zr/at2u2S30jtNKSyKqcQ2Qj5qU1
S85sNAZP97+d5PhyrUOL4A4exir4ylgw26iR0mGIfe+6CwgCctR68wXN5dxh6MUy
Zb1PQgeVBXAgf/0rGT9hwc2LHsWJD+lyd1Nju10wpHDWdtUHAi7KcVz4LcV88TqR
MaKGN/ZgbY50ioH9+I5E138MYImj6Us7JD8yTrrT0LQyltjUquxpnrsPKecbDhQU
GsB67qfWGbc2rxGvAqYoGIxHXE1jK1Q52MapWqlQ3jwnOqtUv6/pJrmJdkUTzdcV
O9FfqCnOAZB53/obEbwVdYq+tTMNvU+0Aht6lksbe4udLhQCm7CnzT8eLKNodw/l
zT+5HAmhtcnTzaGV6xvu7GNfAKdxQi0zFmp4Ai7Ewd9+pRkA8fEIQwTCT8WyQ/Vp
RGg6OngdN/Vx5EiD8zW35sn3TPa2qHwr9fJSGwHNB1tb1p1rhDOBhpEqpCXdxzAV
HUSWnr8d2zhziLy3HSoNJDqnvXoi/Ssu0U1VTHF806+hySF1Eb+y57kBng1iLqem
ZqgsuZ8yXZrqbwDCQCXPabnUTxkMtMiQogGDFjta5dfaXvsoo+t1NdneftmV7jML
U6AODlzx2KUNl+0yai2MvsdkTkLZRalA7q+8w+Ot5n84up17Bet6OLo6/Y/WWzBj
vdyimz1SOgsBpictbBCQ0cVms3kLCi8J9IcleJ5BTD0uT0pr//1mU8qhvq5U1duU
EXJNMCPiH1ncqEyk7oCc9mcNYdo1Hg0f9h7p+Jj7YJePJrt0WT3MNuyIJL6/rDOU
yAcjgQfUPD2muVxcWwroiczZKGTbGpS5MKLN4cRzKsHkEE0T+62OXq7YZdIR6cNZ
cg2KiAAT6oOcU78czG28f64hRF6tOWW5jA0mC+jFXLHX/G8VwgYJ+yVQ7PMf1Ehh
Rlx5SlmyEobExmaKNDU68WXwCteKVZU/kWjbtQDF+02EmGrf/uQMYSsBIlZgJm3f
EXBZY5JrXcgedaxK2yjBcvvQJ8zp628ASA80m7hioDAcGdXGkHWVyw8vh04kDIFH
qccTFyTYYYSAIZkuXiseXGLO5FD2C55ynE2zGLPXKzzT1yiEI40gVDL7OZXs03Cs
8lTZBzesg87vsv2YPNVORe6IUgAqLADeu/nekFp5P4+fzc2i/BBTQdmCtJX7kgZC
xHGjAXeRIJzZ0SZvKSpt7Tq5ydvLbFOJUEKF/TfzQBWoMHVvBll7Q1AadCGdEWd3
ekgzwV3ywYvDtX7HvjWEeoqtPrjJmyDNnvaNHIBiIrWFL/oaKFPPLmVDK0orNRT3
QmhyiCxanfmuBIdaj23FYC+mdOXSN+YHYkBE43gBcR26Ppzd7wse8XtpJVnGG2nb
Zn4UXD4W0gIpki8iM+Glvmo2DD6QM99XhenjfUPCSQwmokqquCrmo+KwgpD2r708
AiFzp7KYBJUKqo7rhn0aGukLW63cQaqcBOm/IZ29O9N44wKZ488xM4beHnUFnup3
/4pqJp722p7PlSMFz2g2v51g0oqLE+VyeSf5xDEM9/jsi4w7AeGY2N6duTeTKJbv
v6OQMVofFZwQkyh0mZhfOWLrEuY8OP55PFvIJO3XYciu07yCasw3pApHNZAu2fAg
ubXgEDhxPS9Z3J02yzhDAQbVCWKsqYBM25F7oSYBZYOzlogiNPLGqzRF3VAJUCoS
m56JF0ALvg7W3AbEoZYL0oZfwEyMwf9rSsUMtR8CJb7WNXcrrCGhD6L/c4LRsFtN
vCTS1Wjmg9KbyPnVkiFR9w949q+OK9uiNSIFgu18BMQrjDgsdSirt+o/NueSqSeK
6X39kmarHFAT4hMLoC+wtuN0zscKtnKLd+yt9QbI+kWHLkpvwqZ0uUQyC+WLqGEr
nc7ZFJf5NCoKYc+rp5fsRLzywJ8XDDo3gpwyln09wqDPwj4IoiqpRZO2lt+YwwZs
9XoomC7l5UhPCOAM/5zkVpUNZu4JByddoChbpOAZSbLCRHbQAbg/oIUQrWhXDMwg
brT6nEeJbiQiOpuLo8EYWkHMZSu33VvsI4MbRCcBUGmCfIF8uwfOXpOv+hS54Tc6
KiPU7XDABmNZMAvwvMsjKe3ASLdk9dgLdiGZrUhdoT4YOfvCK59s6xmZBzShU19S
xJhI1u+hwJwhnqgDh2GF0yFIDEW0ewkHJ6Hfiu4UoblhFv8Mkg/Xk7mEDe81q2VX
I+KroypojigUarASAJi6GwTWw5J2RaI7m1venQdxnjqtmdUOU4VjByVuatKEyEmb
q40JdifPvJRHmt1xcGTr6LadmN87qDBA+7ktHcYkxdXWamuo1yaZGFSuLeXTvrl9
bt3AfHM80ULgmPvfPXvIr+EUlGiibGh/1qte1sJToykQoEMOAsKHqMpnSV5qLQCa
P6CfLgW/v3VNh3fwWgTMm5Vj0H7cKD9yRNhJn1Lki/Ea56j7zEV4zDPbRCr0Y3R9
8q+8bIUIYCeqWJ47Z4Da2FFCc8nyd6sUBdPYd4zHuli5KZ4qbpq2KXrMbuWp3QSF
4dQnm1zTgy2eCAPYh2TeEZoqccy+oseAO0qcqYrkgUndXF7pFC0RLjOZ4RYhTZbZ
hMwv+jN6vlvy6QgfhE7BC34zA8xWiaumhbXBO2GDhMSgddHUIBY5VCaROn5efJmo
TCAag/lOLzEL6Q+yuD+suVw5pA6Xwvos+32Lb3NV/rGnBu/VkLfi7azC+XtKGkWz
m7PiAnzDpzJ0QIvYiHUAlI2bzb9i9PJuFZoYqK8wsUmyFXue3UkuQS6fwmCI1RPe
FQ5j9sn5yfRdrnWBT5ahKg318TetJmMJsOXNr2/778K4ChVmv3ev3I0fiVvQHQq4
9bY1HVJ4MukyJ2f79wudO1j5n93B5mc1D37tcao7TK4kOTXcnHZxvJ/dUsMV1yej
tCG+p1xetCScRc/YbueeZWHSDVm1SkYvYGxH2aqi7ZLY1Wm5SfDQZhHLCDLhd4H8
u8cVoyb3AHFfcozOJKDU4Dl+azN3xJtKMGd4rdW4Hr7U9sx/oH1TCUzqdqiXWBeN
u4KEm2uXgVMAU10zfdmcbInmJfWplI791kJluBqtsT+ovJzwpLcqMe7DIOb9yngB
uOiO0WX5WG+am7qyNvqddEa0fvXT49fPjgyfQQ8dAry02IX8951+rYirhbEEN9cz
XzDCJUjyuJzhUJk/zfpJk09yO2LrPd2YfUErdHHrr2N8/vta9jXcYzPKYoJ0zbbI
SggIUGdT5+0GnZBeF1aGrPsf3Gb5FT5DZRcQKVqkb9OL+3NTTIiU8NRpaXstB1gt
mlfh4RSGm8PyGkz70lVr2964tm/gNrrCHbvFfukz1KKx5jI/Ptnc6gKRY+mEAuuw
JWlrngKHE+7FRu5vCAyIaZ9HNwt5eKMvT11hDOmFz8BchP05Sxf389vpjIcFDBsb
6Dj/UT9K9QgqzeOMiFeXBnxVDBJId15gm0ZUUcUtXs3Rq3MCjk+gMzIEP/1eiLCG
4cGNCWv4Fe4SVzzKmGuG2uISyT9JmRgngc/Eh9noQhCRaC9a5YhE9mQBeRfybgNW
vUkme4Jy+C4atxGYY58Hta60aCHTVLysiATO9GSjOJ7bU/dEUymBAHi0XFU5L33u
Hn/Fr+qdZYx8lBQsGBGb2hesOpk58gAlT6y0W8jeFOfUICBvgxj0S2kVjNRn1EBZ
1+5ppnqRagIkVS6Ty3At8ErxlUD2g954oA31Y6NBrysIQfuJmlw+3LPzgx0QRrH1
yRiYkfOU//DghnD79bXIdqCHoQTzhwGtX3eJSeIYCX+Lly1u/FCmT/9bbyhx561/
bWZKjqHSk/FJe6yLuaoTdCnbhrm6o500/JeZIbkNPGI/UyAjjLLiw2oa74fsFte+
njWNphe4ynr+Pw01sEfZNWD0WiqPWpL8K3hlZj/4XoZCpc/Bwy4Zqkd740e9jAOc
hMFZfQQWH9+AZ/7t802l8iWBtE3Jto8xx3yhoIOvo4m2gbp1gCSG6URHWM5BISzh
q9sbVSfMVnYhIXSd4HLQuxr4Thbw/doGlcEjcoQRQDim5sJ7pb76rCALZb0oRuFm
9ZcWZv3M/BRWBE1hD5qkUWIuHbmlF+w8jmjwTSgmzFw0p7Xq0lyVmQEtc1gpQ8Tl
8xAAamU/55W6NqkFYtm0wrrEQeQqimJocmYSpNOvKO50v9C1RBO+QlD++vgs6msa
0otfU2VFaGK21hFN8Ixqx/LXAq6zMwIMlW/S1WthFOnTEbJDSI30pdKpFXuyWV7y
X6P6p2VoHyIEtDAsE9xwRuRFL3HDs3YfkQDJEoCTSs9d6rpokRMxHIjQoB2k2ulX
7y+u1PIfuWIOYCOuiXiIgLVMPvH4Btk4W5F8MtZobvjK79ysW2fZ1jcz98YER+Bm
FyDvSz3Bnn7RXlzHbC+O5H4JVTDb6cDhYY5liQzZAN55Ywg16bHYHR2g132c/OiV
e8L/R5v6eeiV/xMwadzgqDKVdQLPS1dnavuJchIg9r/KEzYez3ANHv6zKBi5Fqe+
B6ungurK3McioIvpWvgz+3IXg9oeopk9lj3DghJb1Y3HxdzNqSlo5KKGgW9W1BKj
tgOxOtWdqoFVtJtW7rXnKfJjHvk4T6TQVfTKvlHsiH+siWxV4q6EicJzU9mzZd/o
G06YNQoM21flPDH3aTUlk9KlFirGNknjdVMcLbeq588LAtH9GwtVYSXDiaVSk4iP
pZgHeeNHIVWlX3TwiuLLq0O5UHmcNgRiWP68f1LQn0TpTuesfYQHKgedPNsm+lmL
KHa5w5/04HOJGRvzO4W+iqEBLAbG2twWsm+GUQPMuHYK+QPVH5qn+KW15ngtAmE9
81JcNLnt9BI3UlEPfyj1VSlM1Oz0mjvXrREbigSuQRx3oIDrjsvhV56QX/Ssc5sy
/IfYcf6qeaF7wVF5e3nyy5wk0HYNjA/6vCOPC7v7oSHTnHO8inujFTP1if21X61L
dyLvL09vYisvJYqFomkkdfIa/+bcMjLyVQtI7rFwd8M1A7XQ9DXuKa2NEz8w9mOL
tFk9dXjNQojkoB5G2itSFYdQMaSPt9FaVNAPQuUR/NX8l9iaKtJxxaqMk83oaknK
THES9S2ZLsiVJiogH1Rcy6dhNMZOI9p1OtHjxB7pl+HN4qsIWQGXadW2CfRefhH0
tBLFz7U+iNN3fUzzgONscmOr+adG80Xy1z2JBDxwhXuc8wzjZEhy05VNKGullyj6
Dh7ImG3YCzpUXUrmNqdvMqlV16FrmAqWbVb5uKGTmG2u6hcX9PkCcr/Duooz7QfP
k6x4iF8o0oLhIjKF8PMOYgpon1PY5c3G2h7VnO98AGso1+wProJotvU2h3q+aC6h
WP2iHfJkkpV2e26zYnS7bPGit+Hb2HGPgUbRRRjzADErbnwZ+f3lCLOSTdgUWt7d
lG3eOZLvpBXBtIZ8/2akJ+fkJH5eTTrFZS0xW1QTaFN1LzizGOV8YIrEAYboF/PE
WP0FR3XV5gQZftaowHiV63I5toaJGNWQSOMeLL+RHYXPrdQGcSFdrnap4KM3BxxS
PEo2fyqUf7Df77dTdHGW7pCskgfOyHrI0a2ysl52ZLnyvUEjaQxBeawXd0z4Ajj2
nXKhsIoVSHBFkH1J3ud5rdBVbMGBxCVRoCV0H8ZV30Z1nUT0bkDPU4EQ4+4wTzlP
DbFPaJNn8dqBanLEGCDZZ8wbY7VjXHkxnJip58cSMT7dGDPUAQOcmRoCVaHQh4VT
VkyLoK5wmrFgc4cUM4WncAiJskY+c4u560ngFwbY8lwKgu09jb+wUDiyTTbEWeXi
FOZZbRtScA1a9ThjJzsV5sPh1MmawlDqQ1As1RiAwOmntTsIRY80XeNSpt6X6eEJ
5+K8AwEx4kbSBS7+tTV2WZPgiILfmcOZ+Vb1S2+kcJLvKwJQ/rUdUVeEg1zV5S0Q
AAchDEFpT10JdemVRF7xuIFEfbmDnWBQGUNbxbhv1ND64jAGphujqfG+z/eFgw+n
THqyuqgbns2qcTeUIj0E8QPeXGbeiYwq8YvP35P56FqJXRHXErdOqJp6mBRo6XsX
UtbB49+yBV9ola3wA9EHwJae+GYdnq9A72iAeyFXZ5/3CasbROVklfLjUT2YxVZP
3s3NXZj5Qcc2LkIcjDZ8uHHiLg/eshMqCmD86I55wnYmb3pkzjogcAq/+xC2Xr94
GQZFFj9Ux+tpA6DhTcd3W+X8Hr13XOexY5YvbNzsPxNgT91mktK1z824QID4HHx8
Mc38M4pCxpeysPAhMiVd5E9aF4gL4lp18ks6eJBPV2D+oCmHTN9hHRXjeVyUhgKo
20io19VKx7noemrKoOJZMF4iYqaui/E/YZIK61qohnMKrD4d+FcjtPO5XNJRcmcE
C/mmqQdajGBQ1ShWHLXmgKde++82vHhj4W0WLi5CowTqIXeXYpfBb0dDRn0oElZX
JxCo0vJfGE8xPJFQG0bIiJK8Q15NRkzK2ZKUwS4B2zb6mVwpkhzYlD2YXbI0e+zy
lXHqjWqbh9OpmEt1rO6W+Gzu5YRAkfe1akTtB2D8m85sBgaKAh+qe6fZqBdSJZFn
W9OSa3QkxPwDnxohMIwsWew/pQJm/Fk14vjCi6okiX3Plks4ac6fKpHtu7ogk2Tk
eqSrslQRp0yQF/1ipOt2xwLlUdzC7yilqRYMM/fW7gXQEggWF18H+ygTbC7VSkYS
Ru1748ZifY8fKTWOjdkcc8AEKaIdDS+dOe6YIIe+dUCnxOvWqQersXldMWSU5JR1
xQh8jlYqoIykemeIvS1NxzXOUrQHjBUMxNc+mCINnGMkW0H6Ks/d0qAqwz/ZjX9q
fNYaBiNcgNXvYDgNP4ShxJHAsr8F1fubJHrIFycRqQzA4rLCCF+W8IZF6KdWzrHc
b3mQn4AI0oDOYXQV4GQOgUOS+uOUYGiHHqmZQfqOP8ekCCSPGs9TMjm7G0SLpX8W
fQTmQeNb/Tq3QnaWPAh7Y9XW5/hAKJGgpnInSXBHD+6cCekUjV8+3j9Vthm6cEq4
o/wVaGix6X2Z4jibxpb8xzUgtdxzLDLCKU/gfJDxAEQ6Wv7PjVdrQZ96046yvLaV
YpAzi7LSVZWyE9GjZMKZdP9JY/tILMRHOFW3SEbnPvsk5/4x12VNmHMB10/pmxZ+
hMkK55H04wWLs3hRg139G6tV3KKvHkYW9R644r2GDqdaFsqVGm+ZsPZsqXLALeOv
/PJiqREEFeE3BQG5auqqJ1FJ92KMVMXr2OIXiqhXVZScRKPGN8INg3FEjN9D+Yg6
Rc57GegMSR7KBRclxo8UJQqn3E3PALDKML+NtuCUFJfcYGSLgqaz6LfvIhDxgUvv
3FWBjYjcT2DqVZt54Fmvc1YWPgOSrSHaI9CuHKutbnuTECMb9cWoTFIQLHClFii0
qPFE8iVng8O2OUnJP1yNdZFmU7nDVEngG6BbIu00n9N/3ZFQPz2y79+E2JbvzVSn
qm0JrDGZyKVd0shEHVzelQM/3K0PQI3WLg5O03Iz8r7QUkRahUIftFPZbxq0oaiT
5oKD//WjdIGoStJQY6DzLEZ5MwdNHI1arfi+bH+c0Vejfp2Ib2RYQJw/n1A86XNL
R0fdDFL02dnd0GzqWOKhZQhDig5yNlSpn3EWgE/EX2acFzxkfnMndZUyqKdsh3OE
243nAhHPNF8F6w2SbZwIYYkIN8lYmRZPDn4kY19/ijaB4LcBtznM0U20jkIuebQL
HVTxjuPP6JlPn1h+xB4Th0GiDU9e7KNpwVm9niCfI3yLX24Ok2rdHLcYHX5WNsRy
MMcIlUmtIx9GW3fMf68OukT32ywgSjczyTePbaxwF/pYNTivOotzyorY48/T+fvV
f3ThR744Webd0OSytC5NjOG0IIIQKuBDCKHu0zgjjiJ5GeegZEAD/BrbkDLzDuNE
BodAQOiAWdqLPTaJSTjMRsYO+Xsecq8oFmgZxDmWL1PiVyVpa8BDDYqUY54XKzGn
gdqhSlTCVjdwsnCiJ8pFY7BV4kWhzfXvVgXdToKTWqmN2bZW/4Jc5bNs/x55LIzg
oH3W9oX94Irx/9nU4gRgRM7sybAuuIvjLnZA4ebg+n+Nk7IVQ86nL7dAMNzNOIgi
Dvf3sP4MUmA6VaPlUVDtlME2WL3r0vs1KxZgW2wDnl6kOZV6aFu+6kAfp13NDRPe
mJ/mJRXaMdfb8W8knuodgroMVBa4HCv9DCgbHmg4cXjPgOS1CRgHcgqf1GtAKS9q
7o1InzYdqZtrGwgHNcA8CXFbIJR3ouhXqs650f+/OXku05CF/DkhCLvyaQcChWqq
IOLdNJ7k4dVmCj3Gz8YVsgkBB4orBM6dtk4fjhFQDPaeW3M6rtbeck8ECLTlHWEr
EFljnKsfLUhcpdHpPD0VdWrPiK0u/Wl5i0vvN3iknBu+qxfeEQw045X+YsAxzSVf
RaEh0wM+wC6SxEHOUIDD8ylvwkSahtj3kiWTrOPjNwP7LAyQSMXZxuRITfN+z1M+
orH6O2mrx+vdWjsKzfSNyktIpXZICVSe1LwxZtp9bfxNDRVqk/YppzyOl5mu7alm
PJgpPO7xSFt9U39sZfUz0txPr6DMf0hjVJqEifqN0kI7a3xTuuz5cK5iqWxuw875
oT4pheweucRVPF5NZIPrTlyZsQL8s9aohg3blVSVgzbyFY4ebC1li9NAkoZnfakE
nwxFa1sJQ9D3uAxnaz8GJUOY8e94fmTgpOqsR0cBZu0eRg3Mo4dgm32RnciJmpkr
ZWm8UQDX7cQOZ6s7X2fdvjhZjikSfc8c1cz+ahTpSCqDtEeQrseLE0H1hdRmQ9V2
IPTMk6HOmNjzfwtKgWZQ3HUIhbBWFdtTGCJYhh1n1X3NhzxpTQQmlT4V4QsBk5PN
tauDdU35/DWo9bHi1ZzhVioc3ZFS2F+nUw35ZEsdhZO/eP/7JFdfuP+E5wW7hkGi
Ou62o5ZvQMRiOJoAM5IWC/Et7Ll1xgs2JQNPBpzNvH65b0a3I3mXgb3uZuYf622I
GlAymoRbql7WRhHmkzPrt4g/2l2sFiASD4KV/i3qLyJJ2aSqnOr3SvJMU/Xu+R/8
h3ubFCKi4r8SYRD6GLHsw7i1xyCHn6g9R+qS2PBD3zABNXX7VnkD+xO9kfefd5el
6DUaP9dOVjXd173/tEIatcMB/BsymPXO6tIEgPOewSI6wLWn2oAp6KgHwTNdhr6k
nGH4W4SY1l/EjJw3i/6DCp4m/5W2pJmmqYdaHUiI2nuFY+5PxiQKSd8kELFtFGw6
daMlVkuGaxo2RvwdYT2kloA0Wt9Ho4WD77WCeFnDIO0262xnXgDe1zzy0XkBctrh
7kBb3EyARJpCfoqDcxi8uN5jGNJrLASVNM3ODUZzS1CI6qx5lYKrrAlPwdVH0YqP

`pragma protect end_protected
