// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
okKP+R09AI1TnVOvTFpekv7vY5dH8IakejIdktTLeXm5H3c7n2+nWUBsKYxNSaYE
51zPP7kaqZGOCiryqu7XCkkAO8aCH527KiMNJWjKTuYkh7qrIiVR4fLE50541uPz
ozm4XZoKWzrLzPGCSLKBt3AmWLCl3XJHGeYf8MNQbiYxpSY6IKGRUQ==
//pragma protect end_key_block
//pragma protect digest_block
r+V8XsBza0qO0w33766pn9vlFLs=
//pragma protect end_digest_block
//pragma protect data_block
8YLrHq6jpSoCoybEOuTZCTXtOllS1tSn7K0B7a2HvvsAc95PGqBhffDMhwg9BTr+
bvo9Q/+UprfYMrjZBQrs6fwzrnGE5VAeyEpsU/+WtkTxR5uiH5f++MMsrvYOp1N+
YiILsMk0z7iTMjrV1TrkaufSr/y2POIYTJvJl0TchQnZKr3neAbIvLZwiILiAcw5
SRcfbvAxeZMfVZOxQqUzwloj5U7Q/58t3/DFmX/YJQo8d9N4mlzB0Y5n9IqykNXh
GZLWsqu1vardfUFLY0tpxFuqhLT+RgUzVfFVoiKylPGJ8JiCYCX3qHQ9dCQX1S1m
Jg58IIlWbRgdE1EG5Xl3xE1yTSvt77UtTTFwFqSpxerVWTvF1AvjV/NalOlndWOr
9xkB6xumBqwZh2t6lHQZEN38M/qWD9gVFr8Q3ZoT8WnEdU60rMFB8n+3n0sseRTT
lPduxTbuskBerIlNOl8yNv5Js2KRTYfkQHThUxn0dLn9chT5ePNsIzCkRIDUJETV
GfB5WwwEEwuxBgCblXmsFZ+xsJoGWFxYXNYrTv6g8ESFkKV9V82fcJrN1CIeM9JG
5UBzfhPidF8fPqX04VTk7uezlFNyd1bM8JOQnR0PFoItW6JtdvlFnk8IOJXZZjAo
12ryszsJlfPHChnN9mxHPVa77j7G82nq6FZ9drXKC4XcFshdJKkaP04kTfXtx1Vv
7CUdS6KVL0Dkx4W9oq44drYvZdcUPuVA4I/XzSbma+RgJ8K/pTXBBLia/r68q+hE
PB9lxoQGpbHFM0cdbSrbJpv7exMTbZE1BwHZiRQwHqCP7vhH1jpKOPsWwNjtaJSB
tBHetFLFz6QfDO4JPCsrZ2v+jKlqM+hZFPr71LCEUUncJQbE534w2eEwxfuDnP32
9aFRHBUncgUm1LsC5zJAJgukbkBh9MZCUG/gyign+DGOFcNIUCad4lT5IRUI2hh0
I2+Jqz0lhJwiUV02b2bTjWTenrkBn7Z95T8zwDxez97I2oHDEz9LS5ZyHm75tGPy
kzh5Lm15iTEv30jZH3V7yRpn5p5Hs/3N0oquAoJzCLbkpX46dioSSjDZJBN11GVr
iFkJwplj4meqAM1dwLbicFcKWCQ498Q6wXZHwsbTwMUmeW8nw1rDJZ8KZhZ8cjQ9
kHEsxD1gnNT1vw2gVO7mpZAivGGUvQ1VzwmTBR3QEa2ihvxciYGJPJ9wwHE3A78T
y523C49HE+hXmZVtRjnM4P5VIWhJ3gzxIXz2jrai83Xuo95hvvUnyBMVREQq5s2b
+qnRm5bW7wHJtL2BD5UyqWedfiY8MIX8j42PAbxFWvC3txpBE16UgmqnrG1VUoDx
D6RUFasaK0nTBKooiWE+Veca0dDZYkLTbmtFQYkOMOSJGHQGPCkMV/2JT0Y6A2b8
iEEp9kG76O1XKUxsg9CnJk0LPMlLfEdq5BIT19nXB4XMsfriacPz2rv2EloaUcPy
m6U6hS+h1GvoyDAwEqPvKLpbQrV7AbXKInq/ClRj0T5GrPOz74q5VOAP2UZ3Im5E
wQbY3uGd/l8rEnY7/32fwGvyBXaqXEtn9N/r84TSjeK2yNbGE+2eOoDS3bNYODNH
qbHXV0FV+X1nJyBYLTMWx5Yyv1ch94NNN9ccdO1lJPI6D6Bxk3dVqG0SH3Nzy4ky
1EsofD2l025xO33mnhu0aFL9drY5kniOu3bhxXvQv3wteqJBxqPN+hQ6kjovIe3E
lmWlD3Nf/0IJAAPFGkLHCXf72uI6BZ2Q509eLQayWHH/3BJ3jq4yG2tG0Erg+IVr
jq0XhBLGIYGEJw8OAirgqOxImyXw/Q3ypgvepDYjNXzEvv6dIzmWKGjLltLgfH50
kQMQamyBmHGFKPK+r32XTrJumBNv9DfMxdxzY5nbsR9a+yzeUhcAJbiEedSan9AV
guuKvdHeAnHmHxKNoKIowKHNCoMTO5xoBQDnyMuN5szmu/Gk37DyLsqR/LFvHdyl
RQkCZUdh6pzMS/yuf3uXSoDY/wQPyPd4MjKXWxLf8+ojaWB66bhC39i1xG2O4L/i
nWvKHKznhaF/28HZxFmeU7+PbqGE1QOKzgLO8/QkFH4aR6Xv/CiorqSgbthOoDz+
YQ90rQJW3G/IOXw4cXGt079SyCNFttLhwftoz1fk8IVmaU+BK8j3+CWArFFRKC4y
mb5GXIOsx3t9VQeYVHo06zgD+Ss//sAFwzx11+O1A0WkJZVTV2Uw7Hr1zbKM21YO
1ganB1SqkP750Afbeumj+Nfigoy5QXW7PX8wqoHRHHCS9z05r/Ifdl4jHzddx1d7
rakLIfwFYikGIlceWUZeyZ38d/+Cvb+UhWuLNRR7JszBq4AuBilxrrPrgSxqekI3
Leg9psJhvJ6gw2V2fzL6hRgaVgULfzOJ3sdDqPO3+Ga0bpRkZDwy7HL7NoKeQm4V
OfOnU3e3RaGC9X/VK6KgMvuhlA4v19qLs0vbRFh6gNme/ixjt0wvGfJYNwr4hYeq
6AjXQbfjCpB1C9XHcTyjL29DW74MKzDuBYFR3SqDygaWFsrjIwspehlnFQbx7kD4
QqiXXuBYsyeZHwbCBzjjzkvzEHn8Mfe9YDJEIST/9Rc/AiRHPbZJwSpq1uQ8XVJl
rrxQ965EOCHqhoMJd6benzxbuTMV7zDIhQoeOTlxZZ80a6P3eNvH21bJKRcfjlmb
pIe5oXicEfF9+4mgWQ2tieX5+8u6OhqCQiZoK3tcVDOUqosontIo2fLv1o/WZAnw
tpL1/3vItgwmBO1q8+6zs4wQu9sy3l5SCLsv4wXV9hYvw7GfbRxYoenLEEl7AwR9
YsZaEbO1KcNch6pFGvo91kZCJuax5NWemX+u5hK7eQWtGUHmusIBEL7XuJmxbA+h
KlyL5marCTcW7cKjy+cirJZPpOFlrZsROcTVzfMlJc87tKmEOpInv8jyOQaSEPME
HV0EUCDRqd/M50uaLKIkxWwA1rRJTJBK4whktKaJ8yBc3Z9jU5N3zDzoHw545bFu
7w1JX3IyWQS05kMZeD66vINCxL3xbbt0kgrKG18ikUOLl45+R5U+4dF0tousiDT+
A0/oKtFOlmU/WP//TirQInhZk4spqSYdN+nnzs0g6FhLgnRp4SGBHFQoOKn6LGPN
DwlVp/j3bzhN/8huRcGEY1aVO4MgHGqZ3IkLaHpxKAyRGw3OtjpyPNQ+X4Lk7o0P
NaCO+W+uKu4t9IBNO1ZFJbjvlzMg6NvU/n4BR71ugYapPoUwukY1ugEnqD09nY/e
aq4s0uuEcKEo19t08X2WF+hxKeM95uaV/Lpw3UjhN6HnTkTXfpKixbynJz5P5OSi
YOrJhUsMyI+SrT8BdSic0VScNdBRt0hRu4kMjusD7/CF5OB61zZdkZEGJHDsIEU4
9xfRB8VgCZAd75TQcyDW4+rKL3HVOp48yOwu/j8UeZ3lBjDdGpoJZ6pgVPeVRfdD
yoLHZq4jHqyBqze5B2/SLWjMAUaX6I5uIY2P5S3Uxq54NkjAtA8Kz5MTD+QVWi7P
Wh/1drTrMV+5k+XUlBqldpvV4+lf0zy5tKMWy7cfbBYofAQnq2BSjPfA2Zv2LFBZ
cnYEFMz2c+RSvcgCp2EkPvpPmUQVQS/V4PCfzkb8aqj5Fk+ApkZ1Le2oJl8+ShZ1
Yg5vLpZBHeNTY/NI+qlLEafSUp/zC/rT+tyMBWuSEEoyqTpjafAe4SQnvmesmbQD
1A3rrDzBExhYWTfmxQbNgfiYU2OyE+RPdQRGtPu0YUZFXOsF5Wysr3/IZmJ6yMkY
Vm6fe71vAWpd5WlG+elHF3mzfi1FzQ5GMU7ee+GOJFdcSsFltahk1Zrd7GRvxO6e
yHrLWARRIzsS/y/hbR037P/q2vPf0gzV1+Ig+bd52GWIgOeBEK68FrWxmJrkPI2B
ycJxoVS9pFALXkBC6u7fcGqw1v+X1RaatvQIH1KJmMDvBEcJny25G3HvNbmV8rfA
4m4JjcRW3A6qpC8FMStxJ01PU/Mi25PSYWrAK44G3hPlNbTjHRu0teviG5GZD7bg
3EVPQO0PjbhzpbGcCn/mGnU/sPDL7zcyzEvFjk9k49VCjVlReCmBxEB0HLR1Nsdg
ilHgIx980ddHV4AYDBxp7oan/G3KvZORMHQ1ms3mpb8C/pUAx52Sq2KaISwlSxMC
gtjqF4uXt45ZuMiMiqggsLhiT8GDW8F2DU5gP4RP7ssGeWoS27UjEDqWgjcdUXQs
Cr6jZ/4hNvjp34+aAb19bazFkqxRbA8Nstra4MNjtmDoQLu2Sw7CEcC7nu6PvL3x
t+CFeG+BQJGTDS9BPeWNi1iFl/MAMOPS1ftJuDIHiCrrv6WgO0fYZ6PtGYgf11L2
5wQUCYwXH566cNLx9lqmzyt/Us1WWvdbb1oeDvJlv31ZKSZvdPayY1t1CE0RxhLM
ixZ2V7YOn1vt081Da+rk55mv0vyZqUFedpmI87wNcu7qZ5+YUwB7jSVntDUCM0K3
NNKioQXYEpmeftnvOh5h24Z5PcoeoWGtBmRS48SQUqkvA9X3u7+NprWzDSmyZxbW
xyFcmS0ddSn0qPhPK3jpqb3z93iOmrZ+7HnF8iCSZUVX1ouwh9Px6RHL+NrXpitQ
EwRLCpBVZfDB7BTjUA153XgDCr+Ys3oLPiGUsMDGx7L9xBT8YskYHAHKuIE1Ropq
lQLBVekB+48MM+3CAjxBl6dTIetol6MAmcc4h5/m7ZAhDL336XuqIhuwNnatc3zj
BqsYcz00y0xn59CgJoilcnrWIf5MqCVCPrUNip6uXKoxXDLiT8DMXtIrBAn8dcoN
e8HRrWgUe0MwAq5+nKRwyZmzE+YwAwlBRvGYTehT12YSMD1pqIynk4Av++xFz4U0
3yBkEiqQ2cX01ARIuqLU+Mht+t7eXOsR0gw611i3t9FkdZW/G71ZOKpNsQc+GYp5
coASk9NLl9FK5oLNcm+H/cY5zkPMQ1hsuhYb0sRQoAWxOgFCTOR4Odfdp0lj3TbC
xZ2Cj60N8+AoBREi45YniRVSuyFinvy1WmSdX2Y3FDclHUENateBjSLE8hA9OQVa
IAR+I1VQCb3yn+9A7H94zyFI7EmKTG4cKmCO9cq50Nfh0cdcW7UHzw8QxO6AUYhR
IeAKLT8j0kLG+pyX5huNbyFTqeXGgh7RrOkzQzesDR48bRVO2Dis6yPBszcpIAIe
gjVj9e2Mh4Zgjr3mQWX+v4Pscji544EhqNbRWXLTv1AIGUL8XU3T5I/u6mE2Wcio
wr5yKcYbuO77PhM0pzp4Q3TUq1vrhgROsnRdg1s0/lSQ35ysB4nVda8ly8+cW5Vb
aw3CNgAVDk+JJETRVqXQP16puWQSqg5oMLPl/blnpegWvRhC8XHL2UbMeYIypDt1
dNBXnRvc7mJDl0Ddat4CMlgmyub6M5vYVYfA/Q9IwHQMkyeIhJR8dJcXAfj9XM4q
YanNllom0YsOao3vtgR562UTZQj2uv1t6yiujgO4f4MnmrFSnuQPdIKUxCvwJQZY
KDK98e2htXeIM/PYWpiZydfzyibraEqaeyO376wIFHMydhOaT4vZfOR19PpWLd4W
hg3EjwcGJ0P28liwQQJTe2glCy89HoRZoUdmnT7zxeMT40iklyL0Zs5HhfO1c6Hg
mSfzM2D06skU95LxjajXi3dU4wjtEH7USS9LdxRxNYSMLMzzcQxQFDLRcHZn1/RT
OTpzWaUVzI5RC83EjLlT27mIhrLvvPEz1dDJf7eQ8RinCfI8w3EWuUBySqGC0U7y
crVFRWEyAHHWNBF6e2kEBaM5g/qq8OPASwDmDdzY6BDoPPrzc3dLm8Ar1KcSZke7
pec4kLTB7e4oi6qYkOaHPWSOt+hBXT92vszelPxwwkX10/+U3bSbgO60l0xNlDPq
581LVoqBEfp7LCyqzUSFNNxhEWfqBeELWpPxdqf+bSfD3K9qOqXRzPUSitSaRozQ
yu1gcR+AWdMM5b+4WS7xBBgNQuMBDQhQ7wvIrstcEE08+czy3Iu792FP8rG7lNjh
dOTzuQ3YbK3DvTZsf7JQDQ/z4UaPbG7fZJ5mGtJp8fSnIgC4PbkBkBzY+JE6FNqN
mMGZ3r1f6CUnWBXhWaqLnFXdlHDoTFh5gntM/ApUgJPgcRTkDW1qI18kZomaLR1O
P6TTnqs+qjS2WHTl/cWIdgW121ECj6Xcyimo2b4bn8RLeWuRiE+TvLOlnH5o4kx1
zVTydjn+XeZXg7gEvei9VeU1Hj+yQOKmaKzOKxEE4IBVMtV5i8uOFdLpceG5JhRU
lw8fLmpy6DSmi+NG7jIj+tul0o4eWIAC6pwOCdxmMcZmr2dnkFIz/Km5d4JnDUEI
Rf/sEOV42GKxWylFD7aecm84/7ln9ms9TW7o10ptxHGddZkbHJIvJRFz73pe70S7
nVIrGJ36cjuFGJtRZ7hoKtGADra7JEVTwJH+JKiWhQnZNrZZn+h5EvGuJEaasn92
+GB4V3KmtnJcJBwwIkx5My6G6pQ7V2DF7ha2gW/tyNLAkqff3jt2qT9fuR3bi4cW
0kkneu9X+0FHv3gVyhKuyCG7tmLRLbHv3DQFRflvz+z9Yw5PLiZhK5P7s95KF5KE
E7gyEXAozVPRAQOei3Q6TZh9KQaQFRKqSogJtROynM3keoxc0v6i0WedvhEtkrAP
rCpJgwldFdk2eearTVw14aZyADYZrV257D4lANb281sD9OwsHGUOQC5bAkGipxoZ
IWAFVJ+ZXPXb1Le5+1T5acNBtiwCWmO0Wa5s0pfGR4/haMG1BrIO8FklTd+Cl1mO
ICwpZxPtVtqdyVH0w57P+kgzh2RQWOuPAT0tgT4A55j8EB+/Dgg8qSdI6B6p74jg
xLymZU3BxtHqOoHf1gR+oABzFkx3uz+15qk3OB3Ll/knVNkUAhFV8IXwXKJ0WJYa
Pdnn1GIHKft/0hjp+C65kiKDtRz6YSghkHDOjCBINKHAEJqNuhHhQV+jYxzlf76r
jxJGx+jAW+G27mCg5dLd407s25xTzpHJ1GhsZIKgB/U8PGIQ9ZN8Ym8pXSOFGLmF
p5dJhDQEjKPiZsbJ4IrWvttL9mYGmETZg3ZRw492MFhgp1nADV6NWY0ocBbYrHnc
cZGkhMLFh8CQpqcoSvkpSUKE3TsrpopFgM45/+1xN0J+adtntjXpPMSGu/nz4nlj
bJY1PJRdM22eb/4DjLuzrnuTMRw4J58m0i3ra2hwziQOmb4u2vZVmcK9MsWGOK2a
dWitjCtmKqgG6kAR5yxUrASeAruSO2HlolK3gS2ccIgylOypzG3Fw53+FfQ8cnjm
kHoDsUvf6d0J1npIBHFawGyIVQ5KuC/qwkwEBrAJKj/xPmYBvMwAH2iEFMpM+NEa
c3RlaEWty58WzcNZQStOsFAFRiD+pKS3ZFFIscx7RHLCiks5U2L9w38bC+uS4w0M
a8+fl+qBQAnNW1COf0ilvLaYsAjmJGKoAF781+ipMGLfKtDYEEwtwIhNXCN4SPV6
uFEXRMOcpt+LX64AliV86WZ14pIv1563L/O9KbJjTSkZvzkr4WaWbHgn8SYCZtkL
XsKjAUMLSxvVJiiD/LjYNBUIl2f13eER3TLn6X33p1TmuVZ7OsVW4Z0aDFffExuC
n4M7dLYX1JsoJHECxvXaNHOPKFw0EiZIzmd0GbvY2+NqALWlKQcn7sQABXYllYDv
zoBElCtq1osnQ1pSSsGk1B4RxsTHyoMRun8sI0NmTCst0Zz3esiE1xg1fA03LMis
A8QoW1RvQR/2dLGZXNOmTj8yQYvzqb0ly1mSaUv1lRH2a7q6Dh/0TTG/WBB5XxJT
cxZ6I1soGNPICmRV3re2C7oVg7jD6uAhvTbcDKiB8CLFsu9mTPjj+mSXc2+8EXlX
GDde1vmt+APmr/dYNhA18hKt0gFpbe5kVAwIDZbpTH3O91G75i1Ik3gKSga5WpwO
wr/gMNAeIwFV4k/PMpQfQDhgv10syiTKFUuCo14/4ANk2aylA9uLg3iCZdFU70Ps
982pddqzEwto1brdyJfQFlASpkmaXWtMtcoua8hrTgXDID8VQIlRgVXkvCm8MLUC
YAI4n9rvMn3JLjFHT5ZWv63e6UYy6cV7ZRzCqH3Dxtd9u09npZ/AT3TZmZIdXfka
xwlLA2PJwrE6SnqWN8+sOumxtUe1HAAuBdRzOX9DioPJ/G+FWArkeIUisZCfrM3Q
9RZynJIhPglt8MyPajFmx0GO8m29QkYf1y7BA3lQXCNWQsoPuhiScZo0Pdn29ca4
7Krrvkn15qFTUDSov4hN3xerB4anmKyO3JQj1TQrrFVpEJKXvWsuFCo79tl5D/xU
9VijXCNbgu5HwNPeFOkVnnMd36Hro8ymYAr+bcri4NnvNiG57Eiy3/gSUbeFfK2o
Qjn3v6OypwoH3cZ1YBgdLSCzP4f5tsLJeck6FkGrbNgdjzLg1TwjnVR4u25cYoPi
05u21i8L9KUh9XjSfVSlAtgh596YFTOPKPrg7FYjBTTxg09QEniVQWGhBcd2hPMn
vuKQ/PeWiJ67L/iSbi72YJj8gnaU2p7n4aerEAPUkev72PKYusqGQJT0QyLwKnzH
XQ60Q5mnGVoGMoEWmns3FHjzO3mcCsxr7l5xUiUP0fYvx0MGiLXGIf5xvhVE/8BX
SckJ019Cr0000q4El4ZQUWJ8Y/caY1iC8yYxlqB4hNRQMf7ktM9/P2mcTIdRbHF8
dnQcV1rYyW6U4N1EviEF5s6LZmeFnyoHKkzhjsAZDO9ZUlU5Fd/2sI/GyI4py8iQ
ihFqJxCRVwihManqiMHB2yR+TfMVlOmMM5ryB0sluyHFrcVk7CTutt4nOLbztMdn
HezmJjVX9/A3igJRD+3A/hCdBUqyPnwiCK7qz/0IBIKUH1VrI5Ql8kSKJr8L9wGx
R/hV/773VS8U3tK3HiCX6pnjarRHdH9g4GYaTepuYDvYsvg8fqsd3gMsNvAZ1BYa
bxkEWugmQ17IZakIgNlN5WNnCzdgAT1f+naKe9a5XiyT2Q4LANlOnwGBWm3QFLJN
qj7XWnsvURM3wvHUw1Xivb7YKBjRvxt/AAJXr1l7W+Yn1TXilhFmLn5nrCMZbdww
uGzCp2SvBbOdMgELwAng35yno0ZNsTbLrxR6k964U27sPWTHhNkKh0c9/X4LH30T
A8fDWWL4mDhkFpfIVdwU9FF2G7FK4rH+WiXs1bNCcd3GyI32kGZz1Q6DKKenTEf8
lBO6PnNJleInAzjQt20qJHTYkR+ljc/u4NxKqqaIaxhqKrnggOw9Q4bKq3xpTqgt
Cm/ijVUq0XMKt2AvtxE12FE/xBNJW9od1XfS7zGjf2BY0zNYRZNK8LGf98wdIP6u
/shJrV2t4qMma9CHJHAF89ZmVD3SbkwM8xMrTcaDP8E7s1iGyDwqfsWKlCQTDEhV
WPKtlMTRQ2ju8E3zU5DscyypLq/31RkwDNaXglrijxsZij8X82ASQfvNQSXVe3po
83GS+lWNKK9u//gw9LxWBbniTI9FU88+XDQvRL/QG0kcsNMS+Qod3R8Ab0u5A3NB
7cn34WuJfhZcVvXCkhb6W1ItXwmwKMoaRVy7Xk7rj4AUdacG6lGx/QKmC3sEjGXq
ZjqqGAuja4N2kaND2rH2YaPkCwJRRrK6uxtNC6tXtfeqCnObqFQoYsJMLUjq1KED
qysNaM2K1bbdq2q+BqcLwNcgn2iyduwAm4Pu/VwKzFvi8wFENMPfMiQvxXFf+c5m
BsFQ4fRvDObTaiMwGnaCSe+j+m55n+ApVDlfiIGcbx02pYT8XjLHDwJ4ZBeEEpjp
lldBt4XEPJrUW3dMeHkKbFmz5owkr4FC5eO0sFRH6DQ825ekArIWrx82Q5Bn04p/
VnY9OALwUqdn+z163e8ZPYWiS6nwmMDTl8lWJK3reFV8MDrlryk5BV9Ll0alY+34
54xQOOVBbyR11q3tUIN2A8XIBhfJH0W51xnTCUhtRXDk5K2qCyQEZC6T3vmYNBz6
/uDbLeDo4IdsI74jNI6QeAD3729wbNUS8JAoCUK6D1VFyCzvEW6R6VQZbsSSoLYr
Mh1LKW/zvUQf6k0HNjyasCY24oYTfqikZjJkIXxqrb8d7pWmW+RYAMofub68i7aa
kRxiYzLu1J9xdzhMEFd9zaXnv5ZCEiuhHY5LheZpa88ZMgwL6Z/lg4rdTiD+I58y
WuY6SHHyQDMV6X5OU7OvzvFo9nx1adPlzb1VPtEXDHqHIUfayKWueju0xMM8nkWh
Z/TSE3PEWJDbccXSv6fjxo4i7qWcaj/kX+yBVd/iQ6ZlMf3CEhu3xh8adRJr4T4A
HGuPfAMzgjp1cfUdFOXRnXVPjS5r/HnA14b+uriEfiDgNQbl7NFUWtSStkwFtv+3
+PDUJVLa/aV+P3ruQwgm8EjdTMka/b7G/8+DxBXI5WlTgGg2sGbjORXwYpJX4ITP
HwQlVFxI7gDOoqhJ2bIw2bfIlJA+NxRb5R4Mpsp66dNMmpau424C3dO9cmZOUlnB
utysUXMN2RKfs/34fEj1uDfyy1h5Yl+CIMA701rZKToY9qp9/UTnGfMkg2NXk5Mx
+jPzg9TWQtt+F2vc7Mvfsnz9UCRz7/DThn0i6hCt0u3oH042mtaPE/qDEJCROalS
tAYRK1u1pfRHpFNV/blNM4n7llUrDq+bQMacQjrq9c369V+jAeWj1aAMXxQvsWSu
ef44jKryyUmrijwfUPNukZ2NK+SsDZQpEPmPw0vVXlm8ODkAL3/PL0WRERN6CsUr
xPI6Mh2G7S3xKUMhOZSXWeeXPyg8YZZN0l+1+ixkk1SCKxyL0255YpvyEtUzFs8N
Tm//eeh2+FVTYgIeN79y3UOI8dpgn8hMALCHr/VlLRFnSBBNrPHWb2OJ26INiWPZ
QBswoTXUkC0VixJ/UlEumabPBwmBAGOqTRsDv/m8JhG7ZfA9GMhrQrMvmNbOnZUo
ERQr8UPXeJX20LxWu603rO3AK/xXjqEHc02mhp3c4a8lwF9g1aoJEcp0LQOJi62O
QtIMF+MOTff8NoSWwmmRJ5cEcl9eZGXyJ2jqNM7h4iPhPOAe6pxntrRmv6zhDeMZ
jFYbl/hbUPpPl7CcTSRg4MWjZ6ejDsInfC7/ivZCWkra8zzP0kQGVzPVDUwAG5hS
qD/BkHXH+Q7FPENUb4Rj96yueS0FcKx6+xD0v0GfK/6a/7Lw9dITS4PgWXAbsqgx
vK4PQE8i7aHkqwEvFoz9O+ZaE8TmEetDT3TnxAQSdI45MUCYy9nMeK2jWNraGm+U
IonZ+AiXwUt5gkV61/xdWrrBhtbE4rj3wZGZnGg1ohsH9w7u15qWmzNgRiF+1cKS
g47VKjzMUcGsorvv/evRH5TNKwFfGj79thx3Ey/2ZndV6uhJcQs/AFzdaT10FmE9
s2NAfiQ2/cGyzdd80lwSZ3E/gt/SmZ2165+WeSeEBuYjycmrIgzQBDTIxPuSeHWr
AxrcIVU8Ewwmynu1NR1Yz6ifQafK6RbJzzAUHfwZwyurzpEt3fFT94MPqIVYPQpe
Rqe09pmlr27PnMEptAfNIO4rLVA0j32ixjKVdOz7Azv1Uxr188yi2oHdHk/lme7F
OPLFke9IM/Ubox5+MYWJOg2C8V63TnghaD7gydGg66gTmVAsV5t6WZD7LaYx3krE
4iZFdjDuUCYSgSXBay2e4QYhqPpbpx0QSOOJE3eE6UuctvCfkb784uw1RUDWeUsv
9dzdtzU1BEOOWheIPaLze7xVREV7N8n5+U4/8sD/BXwLMi4H3nonhCrFXhjyNie6
OVHQwQvz2yZF0KTeKUpLnJxogboK2vC+p64QZYDbM8lhl2Ktm9ZpbEfNvrmPDcN8
dwe/lot/F8+BU26dAzR4XrjiLZ5NAA+QWimgCO8E1hUp5+V1QATCCw+UPXssXL/p
0YVSiMcfcb1NVUzQPFCRleH6ebBSPd4gWoxiaFpOgCRtiBQ+RGJMhKfzRRhOrpW+
qkyuKi8DIWwRW1YU7VrbUwoUZP8IdW8/iundrCBdGXwdZh+qhViHgdwyVWbOravq
h5CUsn5zf+mWt0xStxJqODiy8/HsBzOSWwsZW15MB2Gzo3KUxfLcWRsVllOMcFsg
BXfeSu96yfqe1bs5vY114y+LaSCmbBFKjWTDEYUxH+rWV4iuy0JSbo8ZwdichS/X
ue7lqLzuXK9agU9Wdnr1ALe6oLEsHMMXb6HwHmkyumAPLkTWVtXy4tXbL3uy3ag2
QnQIpgXo5DYsbUqhcAMUAVXKTUMPOFHBubP02f/oNyDMbd0ENMiY16NV/uzg1iBn
8TEWuU1qgJ2OxOQd9BqfTa40hkt9N4x4Dl+aEpqT8yE+6ZThswzP14CaWuxRfBWm
i3TUBtuHAEUjxZMJ1z9P5hJf8a37T99t957Z+HYKK/9o1l2LbJmbuvBvFF1cOvQK
RnMGCGJ2MPfoXLjOGnUmkxDYp2xU+NVQ8KpiapFZYd3oJmkQFR3B19WflYeiA9BH
Uaerz5eeRbfSdsH4M7AzU0TJpZx0ZwOjgVACbZ/bU0j6Qp8mlc+v6xbOtGhvkiWI
KlNTxDm5PaR78kAT0SsOos7kiWOm80KJBNMc8fXTJhrfKnlM2jMgoPwLlEcea8I9
4hZTtNkUNgqYpaN7BmnSx8J4B0/J13ZUUPwEl4hv/M0mkDuzleJSv4v0aGwAP4ca
i80R5S/rRv41+Vh/xaHRqiAG6ZeDqwYEQfnqjV5we9o/k04PtxvcfM5VckJwPmNI
tvVatbUdae/4sGFdiC3W9EZMUtlCxWxdjGlht+guCJ9Nc7G8NSi/KToQv4YwTAzj
oFWaKyMpegCGKlS3MBdyu71FWu4HFjEMF9WNGv19v7nUMF00FM03BzBK20/gUOm8
wCJ3b2arcpIFMwv3qoKiSu7cxYrc+gy8eR6HMNuEMA2BShOWjHgvjBuEzSzobZWO
QqT7rwPsPpZ/zliWz4r3WB/+8yXepCBsDF36DXrlnaRzIbk2z7pwvevpJDLvKbh5
skQOkDPSzXMO6xC19vDeqpLjCvJA2wNxOS94vsBWFuDJA5YW3CA2vJGJB/AU4QbW
ClhbssCWUQ79a4AF3LbCfaqiLS0OGpN0KlPBIwA7E1t+Seu/ppz8UPOTo79sKSmr
QvtuaCVXR/sPfrNfyXR97Lu/iulh8Sm/EAurvpBqqzLNpac2nclF58JmnlF0+fjR
44SKyX9IoOBmcSZopajbQPcytBPBQJ7w4vYksbVBEUW4zG3XlGUN0xfIt9yeT3Mg
tm32kbA3NOsuKsSr8Jb0KzdQZgzYJXwtYRTWx5grYZkp+wq1VcoKl6gzbukf2UCg
ARTCMxBUj0RoPg0xnG9x4T0fGp2AOE0U1McBG2/ec0DvKtWRSk5LTNW7kfYeMSDo
a2EbijnbnqK4bzHcTCex7+VUd7kFqx5VGr56gjPsOVYH+Z12xiPXzuAYh/48aLDz
ckcgIRZrF8ZO+L92bhVYQblaMYQZhrqSaHsWhKI+vCt8Il7L6QfI/TJd5EIA9hdG
SNCH82NREmz7P5r2LCU1We/wo6I6YYPUPjKluCeHMaA6juJybBXigwvRTo9iXMy5
xQuBH4UNMPvOcv87fJNHXlmC/BrhIR7HRTUd5aPdhR9dAh8ZXn6r67uJo/xVrhsl
g7t0dIridh99yvou1Ftg4fGNdZLiaUH1TFIdIUueqkVfour34+iDrZ6BMVeh4yzl
lDueBgu3VjaH7jd/+2Bjs8ttEs8885tyEDK9dsj9a6by0rvlreJZ+xSnnR7WbZOY
EYhLOgDvwc1VGFrI9PFw8EGRN0GWVbjhJyhBeAmh1ryRN0kSAudsq66GiAZzMxxQ
DWjCcEHK1c/k5Je02x8ehz+5ftRZ7bFlRcEgng+gqS6ILEzCO4E7ZpDRdqeUyG/2
bkIarm7rJ/bdgZQiuTX3V/RK3r1Iy16EA5MlHg9CPXSbM2JEKIanz8xqwyBAv5GC
rLJ1mYN1Wq5Uu9/M9uhgYUeny3B2dvwhIacjfnGpjEwB2p3abBLl2Cx5DnmP8X6/
h5gvij/l/qSPT9+z8P/z8NXcwFS13nVd4oEAGKnWoCZaXgmxh5tNrnZxKjSNrL4v
/m7KG0HpENJguGe2cXsAfxhlK6A+Qy9FmOKBqFpUPEoFnMBvmChuGIHOyOD+7eYQ
bIWHR08HDQTD+VVDJmg2uvd9AEP3YPpx4/zWP38IGRU+DMs2ewFShY5X50dYBvzo
hpQC3t0p2pp946fvPkXnSS2FAfPkz0Y8NlObVHP6Kv80oZtd9tu/E8xDrFuJZJdM
7iOx1LF1mMDeq+MfmJe7pfepzJ5YA5VBCnjui91vOlwFeOQyUOLa6gOuodRGlP9U
ilmFnJDGtp49bxwkUJgZICV5ZVTjnDnmX8JVVaG1Z2+mz3qAh7W0wM6JEdXDZIUY
uD7D42rFtZ/hqakIyKXWhjn8x0qNp5sR7XRbGZhHW9D8XUhTuX1jDvKTaNtGjUMe
Z6B2n7B1XZhSjPPM1dR2nCGnNCrr8gNSv6qWA6dfbYyboDcFmr64keXzPeCpO2h9
HY1U3PRCdzTGnCUOVe98OrIM8PFhPz4ZHy/s3iAwvchvQrI2pFuGAuiLGQNyxeNl
MnKHXr4BYCQ+/qhqrCoCsTVY7dbgaurSkxRppYSDVC+H5OABzOP7yGVZAUW/D7ef
KDuabba41MWBSjmC3ue5Gc4blV6+/Ry/5qZDQjyIHyJMajLkn2gt7adQzyCmeeb/
8H4eaNMwulTcP2U+MLTu6T1wq98qye2LcgGorA9fO2OiHE2ymvRa4+56yCy2JyKU
tzrt34ZDeZwKwQxLSrQDhPWz5hMJSJACM2PW29HSZVeeL/3KMKgWO3/HsF9pfhIZ
WjMM5gb0YCobcMC0pcXqGVJ9saqIK2RTsn+63HuQigBb6P0bmGKOcCCWEpNqHVK/
Hg3aJm5ivns4Ev3gyfcIgoaQGq0Ft2KGOndIoFREzkGsm4BJ20HiCUUMIraXtQDB
pYY7LD1TNzKmiuZ99Q6oWbu/Xn4CvH/7IKEDKqkzgu5mRvdZXS0kFTW+xbPXnqt9
gY9JR903+TKcTN+NfsWAh1ajReT7+LXSbCHljt30yB04k9vJ7vkIsx5zKDyk5xVP
Z2PPra7puxR0f2S/AzZuq/770aLWs8Dds4Rc3RMm5gZcHZvGn6OWtY0HmSYNu9VI
TWsCaykkBdIeRXjTIeWREf4ROljP2BojFbCuePLuie5/iqefer97lujOUUmgGfMp
uM+x4MmPRqJV1TttOC6GyL1JJliHGgftJ5KabKy0wWNZPaMwCayPae+qjRL5nYGA
gxysgyMpaB+NeyCz1ItBwrOTr8FSUoE/Kj4xM7FLDbtwhRUvRO6XXuTlV+qe7ufk
wJuMl82pr9N/e8K3V/yi1a5t1ofNpVk4SrFN0TgfnxmD1MnTo8AzNRyZn1OEhbdk
PMCaPG2K/WdN8+c+hLhVG5RuHFrs7Zob7u57a8J2DsIyMC2KLhpQjIu2u8TDUUSY
LTV24eBjtfnYTHP1jbJ+8uSAIrPS+nd57EwZ/0AjDgD0aRiD3eAXLeU/2qhuoc3e
IID95oUKiLjkzu8HhAAN+aMcK2OCv8aI0yTojQXIz3ylkkymIKm/8sJdhS6LGJ/c
YQBjQPchkNpczgGchjPlbC+o5UxzmZ3MUdf43i1suGndoMKAbdmkSvCMcX7G7OpW
tkt8cIAm2HppD/efaI47drAFsMfBuT0rTJZQeAV06R4e10otXXLatDZS5Cc8RPiE
OnFExs8C2ZU/4aOdLE3Hxgr4kwxSMzu1cX2CRnJcvdBB68/DCIi98jVYoKSXPu/y
B+W+NKLc7kpzmHiX9fW8C5aFnwEq+o/XA4+oBVIrCuESE6hSjZQ+1kab8aw+kSlF
SPfeWaRLVX/0CbztJ1qBm01xmJilbnFDfYvKEYgcs9tdvr3vw1FW9LCncWDckb/1
qGNOhguSvnKN0VYU4Y3awvkSma1x6/mdIn9psbFOHvQFn3UpRuU9MqSU5JC+vHnH
IiSebkYVqaQXupk5jgl3ZhzhVvTolO3PgFmAkrdfA6o6z1kbvpWgdSNPE8lZNskG
JNK1gdt+mbzgeMDSd5981mM6Vutvs0CVfrITRWl34XBFlCOt66Uv1SZtYn1vnreh
rt4BttWRhRkkIXyGaAr5ZNtwEMClHvl8sml7Wlo9garDYW6OMEUnO6qWcBd6HRLb
5qcV0L23XQIs3sJvyEC0uN1Z5+eHMU/XEpxxen1wdtn8YDzq+RcFVcsGyd5XS3/G
H5TmWee/zOuN5qz7yvwEEBa3uFmGt5IlwOWU7V7k/LfLfwFqHBvXn2BUGlhnFSmo
Ay8vVRxwVH57atJZ7zmFwcNN7iVv1NieR6HD9XOGxpy3K530+s0EnX3gx46h5Mt7
D0OhwBAVG/mCLphPp7pq8Rl89MtuQJeKiHUydKIfIRd4m05z2SB2BJmED9tM7sgH
ARCFFPf2v8ER+QG2uxbb+q8fNYtjbNldg3nzLyM4oMzYCLf0L1URp7nfSv8/VJBp
BiIY7tCqNz2JSK5dX5xhhgH9RaRpD/wlDmm90EaGgpzDmv0ADoLt6rl3+JqUkvO5
7nuaCP/LLByoQXYD5wDu0AavKkGVG0Bb3B/cMgQofa59TVVwEEvAkwUy3bsnxrNj
/XsN0rvnwPvnGaOIHH6xwuxwra7jty2zNVXKKDpytSnN3lrubtRTzDYkzxLJRsUb
JDSwpJkauFl63FkTD+P1x4kcUXcGbVSodztMsqIIonnhymKmsnLzQZygS4Raxgay
qIrTFE/uAbAFfXZgAWUJoeqKmNGVtYSX87KOqP2CIt6XY38k4m6cBxp+kMjHTMCC
mLZdSjwi9qX/XT4gaaZn+09I0M04qk69ivxVAnMl+CXp2UWcAGohTxGi1rOHLkzI
U1jb1fiW+AUGqJdaRlZD12ADdM5G4p6Qo4uhJbcwn/CCTlu/uymGtNlKV5OPaGPG
kn0lyqyh1htuurkqlpljW8PbbwAypdi+PHLcvi0aX4GHghLGAYlPm9oDAbxH+yU+
mh/OxehoJ2j6uUWq3gY46Zfi/5TI9HrzGjITgLfLnl65uCXlyIcEk4kUcYdWky1n
CNAdX408NTJZNx9Wtb8q8q/PB4TUieo/HGG8ei+thbHBD9RTKAXoqjlelb7UptOg
8ysmem9XYKRLGEqQaQxs+0SAGEYPVcT9f62whc6wdM3tlGt11xFAmV/Tz4Z79kFt
D8sSLOL8odckaiI4blVfyY2kQDEjKLTVyy/fNXtezi0/cVC5YBTsumMpMA36TksO
d/gPFUf58bj07RIQ+L61PGmwouilxvy9hykbLVTp3SfKxdt+i9moocdAiPJ/q2Dh
oHaHisAbAgPHgSbxxrdP3LQ0+EJiqZi/6C2hzLyMvaNvxiSzwUO7nVBvddvWRWwq
jqEG/ILhpQOkorZFaFmReyUx7jRxxc7v+GM4JWpHhEVEPlWFjf8SU/7OZzQkbwJ4
kbkccnAY/GYf6W1z0Mv+jYrGvEzP4zMQhGuJGBKl7PJN8XaDDun1Xd99yU6/sFi3
k+YODq+ZLJ5bucdHBG4ZrIUQ6T0hqU/pAcRDrodfAz73m79gLTwmakFSNS81dZXB
8Tx4NJIG2j7bm/jLJkSqVxZ2wD3o1k/X/Q+vmWjy/CLRLyNRDanx98ayxMv04wdU
4pZMTqaaMrG9TpG+JJ+EYlPHMtkkVuE1sX6kgcp3gUjB9S8yKA5gk42VhrbSle/F
gH1XcR+sssxnCmfIeeRGfkjGdtW3b2+P8k+5i2erIL4cKvoffqRebvpfiTEGjuLn
8mMITrNWwRZzTzvUkAPToX8CgJgO1+Luul4N/Tpk4Uh/kCXugpk634JYpL8Dpfvr
VngbLtoYwFSFYW1SgU6yvcjcicH28GA3KnkH1ioJATlpQQOKLzbJOLBgON100TkK
FJ2wJCPH42qTCTInWoSs2lfPEmO0IDn9uaPna9S7PxkiNTf8m9KpGLcbHWewANQJ
L+det9rtLbDo5P5PMnrAXL0SM1oIHlJcuSr7JitZe1Fyl/u7YqaALH+Z27V0l+j+
2UucaYG5QUIK+r2X2MYaovN2g5wA5zn36xJ8iJDgFQyCLnNE4l+RRNza7kk1mWlB
KEex0AhOZc1Z+ktXYRjpvwP/MVpVjpsGaLZPwIOAtQamgwOGLUSbKCH2uqSkNnyD
vbpXW5pZWNx0xrAMjrR42Z6h2jG/UD9hOk6oqKQG9JFVImAvSSH3DUKGFI6/AK2Q
HoqH1A+Nd/kp7jOC1puVCrg11X5NGGeHQdDdiFsNKG38HJLa7JAMfeWhinhzzJh4
ACe0a0oEq8FuAy3o7+3yISUep9gk42h78mq0Ka6FDotlKTUELUosHyP4BjMSXfry
ObSgmpsuHLKxYO3euG/VzGfFr0EHi+klshhBh4jleE+hhhiAWHP1DOQrgnZPN0LA
4yN1u3eBXZiRB0viYVw23qCf0f2AXEaDE36kkLv9UdAZQAaLdfmUqobgau+YjNDM
TDvOdRjci5zMbIu9Be6G4XU0gcg85oUxAGkzvAcpv1ZwDaXQ1weq7XDtg3hJ/XIs
YeEoefo1yQsxX3UUvIO0Chg7JI7SWs0zHJqHvs0XxZt/obg6fvMhO54QvZ1FLR5w
E1YlnjFVFzUfDsyLelViMwY77dQxa0dauldP4r0skVv++adlYz12MDVq0khqAHY9
J2tMRbzX2z/cFwZm7J/PXTkV73asI0jxsS+R3uYhOel5tE9VeKKOkYGzXXXifax+
CewkGr3Mzslve+uwEkj58HWGs/wIdkGNcmwgUC5FiFrcK0o1/VlVrC0FIJZFUkO5
ItLBdnseUNe5c0SfswFibN+mHYElEAYu5mDp2zaf0R9C8jhgNCNPodaW2uhL51fm
vdiwYMNM/p9FaHJCO29rmM9O4aPcbt2gJJaHKa43IQyrrcwSmituFi/wBtDhBwbq
8bXRdvIRZkMlnbA5l11oXkawFf6ocPy1dt01Aa+fE/LZe1vGB44tyVBAxl5rTOoT
qbg1SfafEOf+oIPP3UdK1NyfLgOJjlCWHn9/tHrBQeDmiRD3M63qMhwz5URITfNo
eyPI9N6swPgfJAJpE+fjmuXmWyVa/Mv0jXhn+4XRDey7iBRgZ9GtEe2ThXIGIF8F
2vfqP3gYo6xxaFlus2mP7D10hSVNugQ1IBOkFt5VNdJXxj9lIPN/GrTfFiqZjOjS
gKZalrh0Ck2s2Bbmm+XBg9yfuQb3JZIGf9YSowoB6UoLE0rVROhyWHkR1TfTttd4
xofGMf9ugvVN9/09W8MBb01Eb1NR8m1bTMt5KqG0xEDeNiktN6kLVvkHcVdcBYrc
WSj7Fqoc0Av/Ro42Qy+s4pKho+HYLRhalAJ0jtOLLbuzNzJFhZxTzsz5P/YdcUCD
9mZuqPLSXJ3q7xnAeDtF8pd1UsPnYb6tbIi3jJXGWlxjWvvJ5RUEZhOuUFyemc5Z
8ZAX8U3cFhDTiWHAHMoWBSofcAlcci82Yk6a4TgjaaJ567jpioR77CVhyUD7nRJF
K3wP2p7HpWLcv70mQl4pkwXdzi4lqvricRncnuccTEEHM7rcG9MX+bOYw1p1Oeac
NOgxv3o6ublU5K2tBPCGLxjVG2ljpANSpWc8BbPdqIe3ravoZbHh6XWAgAkjb4Gd
Ys1HoRsd3ktO9PO6U/xyP6coFMCY9lkVwKws+hA2cTA11e8V+CX+c2NLGLUgvHRL
pk0aNafw5B+sp1fbDLRni8M2Vq29On/mpenTs1TqbGPZy+N4ni2ZSGgPiymM7bTw
Jh0nb8G4C652VkL+rC5WUw4QoUaLJvLVUgTh+wUj9aJWE7+fbI8DpFYfQdbbec5k
XPYezV9Uh94b6SC1X9Stl1D8KUG16uI7nviQGoM+XpH/KDPkFw3vCyCDRlt51pqk
P9gF2BPbYIz5RZ02ZM9wwIbH1vnMNQ1MOwVxqYjYeF5WHzXG+hCl7vN3Pi/FQaxe
04qcUbEDL67wqsap9Vjb+rVvg4Dy+S+0++mp8OEulu4U22qskXNovHP8zbHrfFP8
Ay++MPyBOzUxQcHJxHRDXxJi6+uKxZBwRm0EGnHrbayyKN+fx9eJH7vajvD+cFPT
7n7+sRNm2AMGKirT2DIG4ehWBC+R6unafekxH4iRMGwBMOGeRNWX8nEHDkud6CV9
aM55mOnefUbrdlbUJ1GvKQRJ+zzF9GkNeijpKm2atNpT2wIg6MKL4RNVbf6SXZ6s
/NMLIyPug8LEtvE/xKmWlpo3400qzJ+/RSD0m9reoegLTaaXP5z+g62MRJrDXZlw
rZLDKAlw+NeJyr+IiHCdHpLMA6GSqGiqf4BBsuE751XO7nhVWRZPw59JMA0T4+SC
dJlAiUEJdCI8kDiV/My4m2rK9kOyBFRSKGDH4kCDbEMFs81Z7Q1UUmnLS7IxDbVV
SHeA5+P9ZJzIaFTGRA9JwgWhE9QnR5QlkB9xeyUQ2nb0mHeGj2ELMSrKItkArsFO
oSMPfhxH8L39zsw9pg9M9WI1zrCEtytU/u7W0DjQRkqc8K3YdkZWQtR8/mbvVI+3
NX5zSAxP2tTspsGl+dTZtfVGNW9tIb9BmCHZrfhvLalxBZYG491tFXKXqLcnaJj+
TF6mtTYiU0wN8BuRShdtQqW8BI1T4Y9CVrPOj33P95z6Rh2XJT/4lF3l0qZuWOWa
Zh38nEVsmOlkdiJ/T/cS4FrtAQpcIyHRSaaCBd+drh3JpZmEyMZM/GaUraPiibLq
TNiwq4dL3BO262vZzKtGZsZ9qfGRCHm/OQKAl7GOUAbcapBFKkveOGW+61m/q8cn
N+szeYpXe84IYak7tTZNDm06Pi7SdL3HegZLgyJhx2qf5XW/AO0+kj5NK+vErv7h
CuwFw71DRViT+HAyOlUpmeaANYUNg4Kdt28JhkdV9YgUTll7xKW47bu/9A/FbjJd
o7ZDIKSNP+poEaf6eg3l4b8hHo4v9d/PTfwvoDsuimOGMsXHEkRW3Kd3gwFVQPIr
Nn8myBY2e1jtlaaDiKqPSXHd8DWwt5k3nzQB9bwKLlJ/mBoh2DjqLP8B5GdTb6fG
Kr9aUd7RPzvVAhdTG8+fZtIH4xCsNZqr9f0rH6AsS/L+6+NQCQGTsJgqQcfJhh0m
due/qVJ2yFbY67KWeYLJg0c/8xxDzYQPVGam4BL6fFrufG5fJ1eiIHAZyHevFts0
UegB4Npbe+b8sbODFmMLHAHcy567OUq2jt448n1zIxFo8w4oLzpnCCgDpcgQeMrH
pGtnctM5UioVSEBr/bxopxFdebCtfYpXvYGMA4pnL04vNpa/i7g1wm57Rd7+aCsd
PpIDzR5I/r8qfcrhhvwhEGzxDBCDKOyINDh6/mPfgdmLjKZkSdjUUXA8FGyewYev
NCRW0AITKAB+SFHcvquL1PcFxsGUNsBvtbxvv8urWVvLHsF/JwtDoO2/Kwxx4WL5
6xz9GfL9H68l+DqMnBu1B54oLYXj030XUUNcodD+rXPTacjQc/+hS+aurm3j0c/F
Mv+l95iwHv2BOH48wdLaXJCsLfs63yUDM7QR8KKVqmGVKxcp4LGtDIzHjTqI6oe0
425boGe3+4wYI3JTVxcqeXEAgLKedpgLeRlTitsue4s5JKqISG2Bc7OASVfke4tR
vRS7zm8vgIEpxdY+tapN7iy6BYIijN3GSM7jH70SHdR4wpSCnX7OpC5voXt6H+ho
4WJzzCR15LyNS88/3XM1/SSScTE3NFnQddoBbMebqzbatUFOah9EdKLtCdy3acTH
UElIW9hnwhU4UsFWP/Q4U1TCnce1vVNIGRIkTG3rBY0Qn8Y0WgqbLjKVpGfrSl9R
YOw3m2Sjd2fGdzSbZlb/F+jkVJJ/XUjYKyPE5TqJrllp2lqQRtm3E7+Q1ohV4IBT
4kj79eCj1vH6OOyApdc+qRq2o+xN9bLWn1m+jzzSz/m7YsXTS4Fitsr+0q+cXHDr
n0HPT9+b9JuLqeufcxjfz8yGshPisQA8UIZVGj/zbYJeclLJL29FHz9PEvzU6hBn
K6UchUz7/cWWZFs8H8945v0wATmsOjrdQbPrq6KMoUW0yFUwLxw1CRA0spK88Dil
IphgYM7W9YgkBfEbOzJEnc47dSDQriD0sDhaNvejyV7Xaf1lPPXZsgz9YcDkB4Md
X1feaejLx5uFmZkOtTMl7lvLdyyonWq+r4OcueaCiXzmbzLWiKl52dAl78KSfJfX
me368cZ1JYEMsxb9NB93cvIp9Slti6ZZAWus7Ggf+aVYqIWglARY909cBiUKgE7M
apyt2ymJOwVryWPctH31imoQp6m74CEfyrL5mhmCyIcgt3/Gn+/sjy3ESp0Cd++a
UjuIk4dC/zQK7RX+i+rixzKtaOa1q98bLQdmqA2Ot8Ow8tlq7banU8Bo3Uijx6VN
BYJD6QkVpTDRlF+VIM0QvnkJM87fvf44tssISptycbV1GOAtYsYOHKHk11i6lm3A
+h8/D+LB4afzZzS/LB8lL9a2duitV6S1DYw7f2kCO++DNuCsit4lf+cOCqzsYK1C
3QlacIJNmFSoy5V4eCjmS6hcLlgwW7VTmRt+tvVEUcIFZpdPyx083m4OAQhcJ2xq
sMUg9JmFmofdLk0bnimnybYSE1oaSJGXaLPk68utu93o0hTBTzteVzNoQu1NARsv
b27E2nMqVWzi7dLR5ceT0IoTX4UsSXu71byo5VX7ZFFX5Su19Q58cSEI3qneD6xI
RIVsfSDpZj/SYJLwzuGE1dDlPEFc5SstZCaZ812hP+Qt58z07/A/5O3JU6+PGLcJ
gg/C1/w5PKxmEkqxlq63U0GFjyKNTSNaIR4Ls4qfo55igDc0p/CqLgVr8KESa1at
lGicXkcZl6dt8o7NxOXziVu7RZf5+H1Z3vFu2648vX5gQus1wPhsKgN/D1Ry2LfL
6+OkHlopb1V6ehPawFrH+3vtTqfzWywx6zGt/lP+tP+8QsWSdanNA+Qy/O9mDKfi
qoSrKFteLAtXO0/no1+HII5uypOboCk9/5binCU+gZ8tHX1lekcZKo9yQjkcyHYv
xoUKZxRS3DN5wso7V4Iu/WWkyM8tBGAcDwSqlwrDQ2kmuhfqXUF6+SbDzlspicgf
8tKLKwIsth+m8It/ywGUwUu2pY6U3Kzx2QZbCIXI4JtxsjkHmqHrsK2D/agej5yh
X28+8cpkiMw/gyJxeuGu5LM+Sa5lGi0Q+1HYw0PB9+uAD7oVcnXA3uDi++KeDbmi
7tIU6h0fGvwA7/vAO1xu21NzRiBUbFdK8AemElDBWt77VcKFL8c1d4O74Q6a1kED
k0WD0h9chsxuHTk4R5+rTsR0zCnRkwg9FZUjAOPpCUXfFtW149H8uHOCHVOi3V33
Cw6dgFt3Ntd30ao2yZb2oPB3mJBIqU8fzUknaiYPLSQSznajUjWKZ2jUh8gzkVpa
p9OSOlbIQDPYh1r1vfqcXDv9KPfm2kQ9KEyXj2e+JQdmYqDolTwD0MnW3Niz5Aum
O/V2NVQR6i1ClGpfql/+8knkOsOx8CnF5uhf3pGhHQOVAIuZ17WJamp8jsrmB6f8
rayceMn/YB/gNHYvSBryJ8TNJBfQ6mFxGjRBb/Y2LBWxiqNhbnocIpzS818b/Nx+
92KPzfqmTOgP/GfMlFGthCE7t9qoPIj/2BNXFi9XPZCYpo7BUmwdX5V4mZmMtU7U
MezqHg4DJdVfcdIPlEgs8hfxM2SQfx9r15CPsROgOONDjBh1sTVgG4kJHegyELVF
BWFoZz+HZuBDlM77DMA1B6JRS9SIeyPFdIkVNjEsJahmZrEVS+tQGI1+3h9pgIjn
coKaKrxU5Q6YvvvYCqDxbSoQFTh/+jSpdqLxX8Ff82iFZbrpAz5OAqPerAEOTUoS
X6nQxwMc9mAnorojNR3o37NTDy5nFuN3c130BkLUHXN4c1hyRE5J7HSZDUv0EXe1
8gYvvRQOKuqRm37Knhvk6LG1CZML9WH4q1kIocAw26PQWtty4nH15sCOotzhCALd
0k81LMwQLliqLvgD38iXeAGZojL+vL1PLG1pTPwFBbM7EXVm8lEGBYINmwuY5q19
naevFdxKgnz4YuLw3yibdmNwYKPRhLk5QQCBit0/T5tf1BCMIS7jvV0Kt0X0qgBZ
6+/Uk6eztzBVutKQ+OqJtTx8cMUSsNJ4GwCwGJMJ8vN4kjnpWL60dpK1dXdJkYvG
6b5Uh3ipsY8+8QQ7M5xsatJkpRd2Cu8Het4Jk1bn4z3CsJGWGsUCL8lc6CJLzF5J
6yDaDoLOFy14CgK8f2JsMXhOycWu3TmBeXAmlupULp65G+D7aUbiV2m79xFEV/Mm
OQBBL+lxsO/3RyBNJZm3YpRuGfPgIrDbizOI23agN3pPhPh+pjEOdDRoI0Rz6QAG
sxUOLK9obL28mm2dmVcryUWfBU8d78MMOL7VOvC8slHdQlvEH8Hiu2eiMDJkSVrw
wZJ2D/Lv8V9W+4vFqpv0bOP+Q14V6wwuGPOGepqVZI3JC/EuwsCCu4dhmg5x34Ox
Zz9As9di513cNiG7ZE4UF4SM79I9Zn7baGXSyqBWiFARsJ30HeYdZLxoGvr7TNxz
I2GdyvqSmiC4Zsdo8HwMkHmi9g4WH9iBuKoEw59DdK0fvi2vrSR3eQxouha+niLS
Jks39zQd+bNYoG4owUoOIsHlR2JU6DauTYwpoBN0ZWx+brB+gRSCfvA96vVRtyLo
G5Yw+d6J4UbF95IH7rbtYTtUX2gB7BnFmRk1TLgtlv2bg9S6egCdXHO1l+SlHtWC
eeqVUYPFZPP/6mQTzsKL/cGH1a36PcGd0YyHdkh6F1lrXnlrgO2nPbR5xU34oiYU
lROwyBLaUCb+1ehNdio80bN4/BwblLLL5wGWoydGz4KilpseNA1R+Wq/iYkNUUSp
zLYBCqydtSihA/Ja7WYmmRmi+3l7YWvPigCU51dfeS4471SlAF5Tnjb8mfkQvD3s
okyDWVditOSCfbFhTe3prDs/qO4LceitpTkkML8b+v8BjJJyFZii0VmNYzJSWvlX
uwBUrPLdbBtZu1PGMmHcPJOc6EDuivfNGeUEtnsI0epjZS8xemc99DJS5PGsupbf
iC0u5y0lT4KGPOnmF1AzLpqlp2C5Uxx1ET/iL++un68kAwQnVN1LMXqri74XhCbG
5xjajLWHiMPMT9M6XGl1d2FDRn+KsJFHzOYsFb83hEhQcAOYVlmVmPnS6XPyi7+6
MD27QchqZyCnXHvhaI1lESRHB+9m6gOu3MaqTqR4GwhwBkCFMJneyWOWuYc2q1AI
9zEAGTfzntq9cQepIabOrQh/Iz9frp/ZHTRtRkvGN2b1uYTNdSqeDugZsgTBcN90
T1PE3sZzddmmUOQeFyCTrW/rAfX3M/z67TlH/hysXUTT6AEa4tGPUPQ5XJfkv2tl
Xexh3MYc3qs4eJ5SyODFqbIlm6EQB1JhLyxk2f9VWzjdIaUMjzynUbWq9ElSeBy3
2LcFGi8CyypmDBjbzm3vxv38KANsiJJMZ+xBCfewg5X19COSkT4O8pK2NOjGzMjk
RBIh4ky+2JncPoxuxMG3drMb6tAoZT78cAhtyZnaU02cAIvH1Emzlasf8jDH21By
0UWHEHDQo9IszPJCPdQFgMnAHwL1SDQ2CpJeoQIt9IcdtA3xx+GGUzP36UquVnXo
YE1RIep9/DYKrj+Kj4CtD0cP1GMvQkcazeZXjLqnPG/DjyOmPIMSA274rFeJzFdC
5KCDI4arStsuNBg68DoZ+QS2UqkNvIn5HdHyRB7VwUhJedXZzAS0Uf9Z/ib+HmF4
f65B22qa/VGgO7W7dIMTotTOyxqfMbrsHC9G4j46NRPZOISmaTMwINbtIlez8VA1
3DmNxi6tRwzks79lR1BpILHb5UueiQncuc68ZjiF0UwDTkwPKBxZwYtqmaaIH8z0
cS4QKFGmqyFEOzAgB609YVzqUNhbuOHFqT8Ui9Gwu/iGpyoqxulc6DvEQ6jJWCGE
/qvcgszQfZuCXIAPb+3YlimSisVV0h9kGBdOCBFzvRsOE6JLJlGj7OhS23ruTQJi
3c9jxBrgu/amDh9M/xGzTEnB2/j4BRcOrnJaz0gnIdhN8dz27aCfURu1cRgZ4A2G
o7ECaJlcAKLLW4aJxndKdfKOtu5sNW0m5z3RLmKkobbWRRU6jeZkR4wg+D/ATDj8
V5/KhP0sF7VyuZuW1D5E+5JJ1j4zn8jLsSFGuWPq/91FoudkkDsCtXBP+dxfQw8n
bz2rT7UnmsOK1lsBDGV3oIeOqw1fJU/b5ZBwNFrE0E2/mxfu8RcMdymi+BReac2N
I+GKabV45SXtkXUqk7r9bjmWiDLY8hULpSIAK2ovH/0Hn6trsoZ2/D8RqTI5baYc
/MvQrmA8mo3YJeMTdeE1AXfAyWM+TypuTfXUVI5jBIbElxcXc99wzSzWM2NEsbjn
QStwqD2E5yfRm/SFSACtnFZ0o5q+1sIeiIIiURE9NQznP+q8V7GVcABD0xCJOk+j
YEaaLfqB++V0CkQeUVrId3NangfAQWbExz6arK8wI+KoD/bD9IBMpdGGW7CE9RWk
Of7NOf0EK34D+Lw8xH4xIIUiSRew/hv/sohhjmlhYNEjhxsSZfGev/9X4wSaQ0w7
t76JsI924eWAsvG2mpfK7YIA9+wQiBDVEJ9t5FF1PynAxd0D2K2d2iKIYl7utevD
v7tHECj0ayKDkT+G3G1qxcEtcn4sCfb1pTUfjyJ0V7K0kSljJLaO8VaEIEn6n9zT
PbAehWquh+YBprgJtgc1CdZawNz/NT/y4o7Iy6atF1lN49xGTf6bpls48QMxJhll
plcy5PNSskT/o8lhOvPYUn1nmovgICg4xjLHwrvcm7231mlbEg7cXkSS4Op2z6ym
tzeaX37CFjwZ2DUVH1+1zvvTnMjTZUhhxtRzjkk4vOk3IAV25SpX/blwvDA9mL16
iYkeWR+VdPq1NQvTbMs/AGptFyW6Skd56Ka68FTX5TARQulTFKUqFX9rXy1sg18D
vMijz8OT37YGI9pJ7bzLxDq+nDajte8Yak9Xf79fn7gZFMr0DuCD/4+PzB/sMtun
NzzoBEHeBigDVmUh7QBUiOO+bfx2xZFL/TU6QplipUueCxh1STps+XwTcxBe7DmK
CzQl+H7aQu8AorBbfNqneQH0vfIS+M14GRtpPptGWJ9/Sz3u7CvFhO+0MKTORjaC
bdxX0N9e42c01d9LzH5HFBB9Igi+WTkUfwb+BMuR+QEPfE/fhapOiPEStZNUaLGt
0n589ozwqIMftc9NWplwNByp2yvYZoVIGunBbO4dAkRACBGQaYHSxgYuSUOvvcFP
lrM4tFTvWQfXTCt38UaPMy89Oc+Js/NXykT7Fh0VlZ0YM3XrB7VF5YLl5CpckILy
mG7JX5t1rZRRdQxK1ubAOHDApsZ0Yj7foWw+m5pJ+Sbtn6Car6iVvY8o8BNtBGIm
vFjTkQgj2afnL6iG/H65Jt6wWr+HKNNK9a87bdPd4yEPmvje0pEMNmIEbOO8OwTo
XJOwERFvpRr/Z8h5PmXxKEGPSrQB7uCrc0eQ+F7NRUzxwu4VrJ737xpYnrP0KKww
uom/sRDEzTqAKBNEXn18J/4R+LxG8Qd0vABiR/msp3j/khsAwoex4P82A5EYGmyr
0WO1ciXHN6F9dwiTjYBvuY9nKiQa5gvThNPOlkT3luCbQ5FDG5xDqPD7eSi1AMPA
ErdJdpbBsSlR4kzNb+bnAX0UA2U2r7GA+bFQwHziXwlemZbe7CwSHVjz6y2lkFdL
dqO85lZ8outDt5Fd315+urATZ9o2yaRMgofbcv3kl1cTGCuzX6Y3bB/5xyUzPbY/
tA0MxQatY+GabuAnfMUg4PWA5Kb1jMZ4buzVNPkfW9huI6r4wSX7ydZ5DAoqaWJW
pMeX+KUKfmCK4NkzJxMsX5uUafwsClZAYfx1HnRwOeRwUIxUVTT9tR+fVs4aCL9+
wzKpTPW9ZrGeurjkNIjMG9D5T9QD1JzM2eNG5xOBTJ/w7kyA1/c5n8UDrx1LwJfa
i0mnK6lYCfGX3ZX3YSA2olbLgYSyTAh7E1Re+JQ2eX2u90WUqvc1F01L1nf3P3kO
/5xwi5mRx8O1XO4xLjyfP+l7XlszDz3y6+thdP+eW7i78pclbCa4ShKDKJ7gpZp0
DaZ+BqP+6pbnczvM1QKyIi7Wxa8dnjcIgWiGJpz5StJ2G1iaC5HvJPU5lX4qXaz6
ZjMvuDvAPiC69VoxIOFoCbn6dhln2V2EOPhQnD0bXj4kXyhe9f8gjKNviNOT4R/A
8fWGdr0OJPvFWM0K+BHyO83w459U/vX1+28gI8uYKGCZI3PtfCz32R/YQ+eN5X+P
fTLd210/IennY6Yj0zy6eWqDEBV2SH6CrJnrdVU1FOdUA/EDDyD6czpLowlaphbr
GB4tegCD+eLupmQBL7eXwsEVvfS7HyYVCNmE6nKSIKHvsGd+aGGK1omgpV6NVaGy
C8L/akjVxe+fUyyjcX5bQuvnxYaJOnm7WJpWwgaWCNYKNz+BNkanf6ATAjn7X/59
moZAiBkRTQuSHRzcPsvAxrXY+38p+MU+uLPdSyoXCXKRnHD9r5mwxGkF7sdZjOx4
EDdWdzWEeE4qTKVAwN/lbfPKCKPxG47HYtWgGTgZKRtaEbFZST4EYZhArWrjqOHZ
Un9GZveUsTOCisu1xXyAyTAv95pGcmFn1DChtdWPC5O6mCbmTRbMIC7RC2ezu65z
kGWTiFeFX5uNrfvzB6q9doWxYYSLvCPXZrGQp2OHH1rD8ViBF+470gXWfivoUlyY
f1Cq0sdmgWnG35UifiU14MIij7l6m6x1QpgYuO4whk+hudez3rQSm0J8tNakxGNX
21db1fdnIzEqvrobLCou7M8iUfm2T2x4xcB2flkrFSzYSShZHnB4OvzYnXVdrYG8
lX5CZ93pAWD1sW6dvHASu/HmzPhCviz9PXVR7gQj4+tlp9zZ5ex4a+sWWBa534lK
jglL3Y5R7ud+UUvbVRrFefYn5rX0HSy8YYBxwbQfnFW6vrYIWi9iZfWREgnZjt2F
PZloOPjDs+HVEAAhGTGf99KNbdmvhzUcxTCbaRld6Nb7pUu2Mpm7kMrPr15H92Gd
NeGLB5oNR4jmz7IyvPDY4OH4kYbSj/1tRkGebNIQ504EccCynIRa3MNWvy7HHeb2
DWL4KGnNoBmc7XL08CGftdYJls62eUlbbPxrivmCtlHQjBvm3h4P8chXWwdqm6XA
rMzBei2MYtynV1DBPe88A8XUSeNj9o/pTBFPEDaUqciBOSsJSrR4wKkNzZUk+Q2j
u5OkJXpGE8t8GKR8kHGdSGOlVR9/Qx2Z5EO/xDqJ0LSIx2LMH45d7fhYQCBJUP1B
OjXP2wnNiiRGeRlW+blHQ477ne4DnMlb/f5DPSZWzrSJD2vW864Flmw6DPXH02tY
8qO9r5JYGOLVCBOis/4EBeKw6bF39knP9D46dn0HVXLp0ACK4hxJhXaCxoDryk/S
d+S9vTtJb3H1HYCacWz1QjzgJqLxnzlTqDsEhdfm95j6satA/HAHLCCOcVnJcm7X
c7DHKY6YzJD1pcQALjHb797KC1d+fTj4dH9B/kRzpFQdRTcwRx/IPzLxSNWCkDvT
Yo8z+/D/yykhnuUhyn5GvmCyErTJ+svYc0F8/pteVJmh5MbRzd7A5QVjwQd4qG16
3KGatuleGhAiBquC7CAjotd/jCSSgIuv+icvHt4GcGSPeEqP2W1OtRVnJ0A8Wd4c
Ll+k5TbL9Bg1rKdP3IQ9OAooyUbh0GEVKc/HEF1GF4Y7aBpRcIw1oWtrmIfxWPzJ
YxJtu61R6L6xnedoLLnsIBVi63/s280YGsEwAaBLmHLGyHuu0hdk4TayMuZDBjOI
8VXsICkCIYJjCWGTsEsxuLnUfVgu4o1QqwdTOG1LCG3qRu9MVJtBMVsMB0aj1Ydg
IZhh7q6SyeU6RsAFwbSLepsi41to46nfBUssM8XqmKelLc0r9R8Y4itMBbQ/Vtql
xw6wmXV8cwC6d6Pi7le0uT6IciwgLMrUtnGc5/Z8j7W4LkM2BVEq37F9sehMU0ik
af3xaEk9A7WlJZzUYG4FIwOteFY05L6xAW4N5fPdES+Gqq/DVJStSylf40wL3PJj
OwooMKO8N9Y0fyd+Bstqa90BQaNy0KNE9IYHWTsEx6uIVgt2AnlvQZytA2cKnMk2
UsVucloq6kHyzObo/+jg3F+L6jTxclsXK60bMICCMZo+55b/+hJX3/2mMx28zvSC
KLwklwwnNz11SSoDXS5B0Q26/oL0dGbJYKOtp7hyAZ80Gwe3Q5sp3CT9xHNGvULw
hiupec3t8owPbXndrB2z99Jt2gtpzVNJ58ksGF5gXJMfv05yVWv7FjtkMt93C7Tl
jv0KDDbp1D7LbK8dyvrxOYK62fuusEq8Y316n4NIamfwTnbHS0fPfkdJFark8ae4
4yJz4WPE10UABaS6iCPqUv0OaQMiAueVZjzhXaoJJ2Cu5sDRxVSyW7IzcyshMPjq
qOKteWtpQQHNV/ry7KnUVmUtbMjSZO3qKZuarU1wZCqTRh1BGqgKTroKj3QFu4tG
4O5p6CH65EpRybJZ6fTt1AXqleDsOToCnSe1XPLpMIGafVy1nCxFH1Fd/kqelVaB
Pwwaiqc6c0EF0xa9+HRqXJyOR8dpeVwxZgcAQk3stFzMKahsRudC/x2RHX1ZFlkx
VDk8TUQbYrFNHa6kerQzMqaGMx1c9A2hqf27DQ+7xCJ/FUwAiKHwRB2afBFPR+01
gPvHo+At+TzQ/vgHM4q6PWVG0U1yG9qj6e2f8PKKUwJmlEvAFoBj5FB8KXbzOIGw
8Rj1fCkNI5Bn7YXOcIYCNG+usah2I/wwoddOhO5uarMgh6Kgci7lTmqZ8Bt0umYg
hg51NZBp36BeuN7I1z44s165EPCVqThxiDOiErudxgrlvnRMEKT+hQUweiV2lBMI
DEiwbDCP1ogTQXTEqeTPJdOdfSdkMNlX0dxL6kQJPYOYEbLPGEZ/nBxm0ydzBra+
KqrKDmmVnOB9Xiq0XfxYE+c2OjzWxKdH79h1CrakNB6PI/DynxEei3ezbpryHwC6
fOPYbvubllpwGiXgBlJh/xHHf5WczP8wQxhVONKTg5kbIKjHBAiSE6icP9Z+sCne
59OJs+HSyZH5CQbUpIJRT/tbzwtvR/F+aah/o4vuK5/X73OC+d7PAuNxXGpZYSAN
JIF1DUoJogguBYqtHsdJ4KMmNnlm70JHARUqqGTgrqi31UB2Np8LbJFTMvAY5NpR
UDMo3VsGn4Z3DPLqB5D2jCDUA240+JO5uBbEuDhTzpAcGqhe12LrXkPHaRJS/KzJ
vvgpGucFCsIaxOa/a0+OIu2g56FezKzKrIn+5QgGAXmFOKiQWKg0HkXH4L6aIj6C
sKVl8eYmeRdEu6IEUHO31c1WLgAA/C+7DjyZ8v2iMU2+Ks0AraT2uvBe3rN7A5eA
5RRlYjn4MtH/tRXV10YnxOOlo7x2F53Wew/bVyfvLxDfeRslPRHWaybLy77/LBBU
Y2mR9i4QvJRs6E7wRlkbQp9NjUJkhtyCP0u9XHhKUYALZytFCr5dalI/OZFHzrX3
Q86eMb28+hxwlD2F0lBK0GaaF5pk7++Jf2x9u2pABzq0wbgggbFHl8SI5M5sf98G
yeAvCEypEsBNrhtFg790SuElslWoiq/Mb2kHjKEzOMImQXaJvff9KnJgL0T7NiJ1
xIJc84ITGcp2UdeFTizyd9x7Bn83xrlZG5B59UQayQLLd0L5ZPe09aZml0G0P9jL
3H1ObqayOv0kTBnswvmk9nM/wAApdl9n5TC8YBZNMORp4lIr2R0PIgrgNP85J9kz
vae+UbfrkoGktPp5GUETQSfB+ajslODsTI8KLa8iX4TMwQOnkEbIj6OGKyQ7s5q5
uGyrW7yjPPSkTcGunOkCeuaGVpEN6Mn1HkW+QZgUiuI6gwSHvuWxHLYaFcWI0IEw
9H+KCe0AAIGE+kbFnBo7F3nGslw9GPvh/Rxv9w7/2fJyrxnu6EZ5d4zyyGc2fFM7
T1lXFlSirckBQS01Tx5eaJOJpSpS6u3dSnWHcOFllYdMFC80duqLZFZQ2NLB/Zr8
OuAKA9G1HgreIwBkEhE2FHs0a1xtm1uqg2rKTuibJ2sEklCZXdPrdAldH4Lzie6A
qpGiScBWJ9mnj8afD4VsImFI/H+Uizfp8bBZNz0y63e8b1qR0Ggky1QH9DOUk96w
BddN3wkQrx54cnRSING0aRSarcTPmdaelB0DVtWzBvr1BavyKVJea3Uxfb99VUaM
ny8Jdr8qZUUwzoX1/vQ5A3UjDqEZ11+sz5R4ZIMHu2By+2w333DV9PEJ4wodhlMY
CkriAJp5Xtxijpvh/CCrg18tkKHvtLPyzHpx76BcugduEsP9AqsTLMA2eWQqnbH5
YtaRVzpNCBUiOaYoWDvNWIbvYH2aV6VIzyAPw0Sb7jSKufrIuv7W87yQ0TvgwPZn
GHWHTjBk6pCv5rNRRofpY+V4tntpCyQw09+HUH4QY3Uvml2wAaZWQR/Jr/YdwsGa
Zig00z5RwymfzoLvqpWnDlM61fH9udXUwuycuK524y/FRjVoQgFAIGajtJNKCJwV
6iqRLmuOsSpmkM5kHwIr47BM1sJ9fQbSMvzHYY4vM8hauZxT9rpq/83oSZnouqlc
HImGy+nspYPX4Ud97cZOFrOkjPptNCT9zxS0Uh/n9RySpliKFDrkm0aSZMZkHUMn
Kb4vgLDRKyRXC2ENJ0vmd9B5Fv5Vk+sLnUIAObc6gO6CEQajV2qC08ypJdxCwo72
CNc0BO3p88rMDdSX57MldDXoCk5Q0mK7IWDiUKv/N75mw8GIy4rdDUsWQIgp0iFJ
3ICef4QDXxaaHoNYwMbcsYfpMI6uaLep9kQY/OVJNz2/CEGeq5Jc/fq9JnoQEyGv
HYXnPv33bsf0Zz7e7gptb8ZY6BWFj1BYCFAWH/dyM/BywisN3htrQR2hB8enfyBy
HEWUu1gnIyHzCtAmIE1Fvo2tdJI2bN22BoB9GcpsWG51Vh0PMuv7Iz2W3NNCWL3N
51V3Z79J+XY1OCKlOuPv6qhtTXgAQMnvopjDVfQCpQfEuf3WJeDmzT1EOrHvf++J
AsUsVim0Sav+7tKNm62NtQ5Lix4wOlD+HAJg0SAF4Fedbn9Gmjt9QHC1jO1Zo2G4
wm4SGxf7ygtAZWSX0tKWBPU9N4QRJ8XI36F0ciAMNalzH0gvyEBINURcg5E8biV+
zfLqpbrAgb+fvzTS2mfAij0bRe7vfsdGl8uR/OBbCcAKXCfG3HfPYqGBLZZutxTk
tJqxTN1yTWAqY859vavhCawZn3bfecy3WoOCCQDPD8MW/yL3WOZzl1czmgzzRpQY
hFhkzGsWutD2kcf8JdkFC7MEyKY2r0CtZRtIgWpkqNRjnrTj0mjgB/jR9gYj/gI7
J6z2fyCUHBCsygIVkHij3JvSRs/cr9xf22KmNRJ0IsGWJE1fox2R2SElV/NYDzQY
G0+l+lq8bmTmyTNBgbMGK6ceYJ5pbco7nipDEvRr1xGaPOTUFDm0izUYDNJLUN7E
uMj82jnIHMpncZ03DmuZSRrDas+JobEWRBfG2dWeEb54XymkKJX9fxjF/XiiZwZq
lZiRmxM3QKE+NNENkVux9o3CFBcAVG4ZSxO+LZiCtaIzGNcCxQ2/MbYn61528CRw
VSMeOf7TcY2VDRlmSOLZHKJZha8eOtIXAPTD7NosZHR5dsnPmuUwqkAmjxDy4R8U
IqHfb527mpvv+zjJU/OpWMqsK8vDTGF+tINQL/qHJSmfrXbrLL6h83vp6KcFVnsd
rzFjYse4a7kxjyHtGMZ75JJlB9Tl9OFUyW+EGr5JBd5j0Ld6nKZBDnNX+weqa6mT
AMUE8R4CzP3xkpoI0hL+YMODntU9IlUPXpWgt6pvo0KjnXkm8yvwZEFm2Dz15GOp
HIuUZsgfa/wO/c7WJFuafXVHDKeyfhsAe3AP/LCs2HWeryQjgHS4sQm23q77iRf+
U3XO8xNmtXTWOLu1vsIIXrS8R3xiqErboHOMAtW+BDZSFzFS6x5RGu60/CwqQZr1
lPxEydkPP+XyaCvVWPeBYwy0HKxtHcznhXK6HjhqFh5x5NMeHofAMNoZjDUoHVvt
Ct2YG/++CjSMXUvTOFhlvCL7rBSmij7LdDVrXR6Bl5QcncyHQkeXJtXKbQD4XdL+
vGeM0LRx1SYuzIFJA4jvkRNg6px9dYrqwGG+c350XVJqy1Vrk2zb99WQuPvL84B4
4P0nxumOztodGeKIoCQyI96u6xbt6l+ArzVpKjPN8ndmvqMxOi51hs1ciE22w2HV
EhRGftoYYtYR83lyvxq4IuXuKZsu+hcmYalgpcgGlZEdkCMmSmRO6l1hHXHGvwao
k4e1XNM+0Y0zbbx9XvdxYLx7q130wprD7tGbuWlYdGWprAkD1o+DYSdSZT62DAah
gELjmwjvuSXIT+7ryuA2s52L7sdss2WHwIEQtSrMdNzw8kM7big+7w6Wxttzgckm
89YqgsTeH8XWbPfxYKAG3laJyv6biyXkco+6TqnSnHd3lD6UBedpQYSXG0fFQ+qJ
So9UFS9RAB4bawPZUQJGy/Tb83U1FT3MFVy0qqC+qpOXeiaVC+HLrSo2MRe/0/ll
jhg6unF2xBfHv7z3n8JvKBY21AJzUSXctxIyDEoYaIOIU+0BF5mEi1WTrk/ESWbf
nBVa8zjg4xLvezhN6OFZ6T907/d2qrIEAhNIs6OHMwzcH08TFTobffPUMiS4xggb
n9zLkm+O/5LnnvDAzRyTlt+0fbV7mUd2UDIpRK15QSPCDwygDVDLFbhQ1E2EgUze
uPAHbyU3pTCANDjQPFhtznq5XWZ1EA9dhP65BLY5Y7YQJP3i4fWs2nOn3GrNCy5E
ygNudgXKdgDtx1F3fPBs0ytKF82NcYT67swkkvIWheW6x4/W4P0ciqxon+HJXerP
5QbER0ST8pS3cBj3yHsjsTbtAaLSWTTkw/6EfwhVbLF0GpF9hjVIi2F6O6JuuF0r
Oq4H5hXG0mX8RE6GPRTQk4Iko21iZPS16PkeisutX29lrj0m+zb/OQ9Pwyf6EgHR
kImL6XuZ+Rpf15Sm4zHno96P7pXtEGgu0VqplbbGGPbjqR5cxceCspxS77fiRhBW
6aWo1L0S+qZiDZyQhc8fse55v60ftYKEvcpcbXG6dBDBpfLQhcatZ0jCpGkRTzFA
LMH542yg20zeg//eeBDJVInbXOVcgWiBKqsKjsJNABy/UjUnc/WXTrKRyXzf254U
H/NTl14REO9G9F3Nk13im0vv56TKEfpsjomQvakVSbRofw0FD+3CYOtx2q1Yv/Gi
ZrCEnVjxVxQ42Xzo91jAsVf9MuA2ZycI4dcS24ghtJ+n4MY738HRHxHv8LH2Bl6v
uI1fNxFviB/wc+lTIrpL9g/Px0r4Yi02iJWa9aNSQ04WDeUKn5Fz66lUs79+pDPl
92Ks2GJLut4avKqjd9/6fJID9CA01/EGR4XCj5Dvyk9m/GzhkdnVV0kHiMHcxk3T
mN+ybu09owwSwmKLjXEdh6/Ys0DcMhWnGlQQOEq97UU41UV6ibwQmCzvEbDvZNFZ
25kGIjPNV6K/3mqf88mBCwUCSA+KtxcXoe0NMs24+D0ezF3DqWhZYguyoqnT8maI
2HFkUWbdWwQQombBYDbktSPzcDdNkCWJFFzPbDDV/Qo+um10V5chT8QJecwepNsQ
9MB4xLDkKGXmos4HuhPRiRgLegJ2Z8v+og3cWGCFBed0gXR/Efivueja6Sf4jCeJ
bfnn7uLI4ONxY+QqnEoOnIGPyPpYzl8Jp3ugnYDAMDHK/hE3PHO9/CdjJjCBOJUu
3nWqsoqnPtuCTiysSZYyGkJdfXEgRyxkDDM73n+LAm3Jm7m5FNsFESQVnRqhatqX
i0Q7tVt8NNZSgaaorJXDquEN1f7hZ/NHZI8erNaiW2VMZ5O3ZUwv7RKNCX6EXjXy
0NT4uVT2a5WHnzQzPAaCAritU+YpVSA/2ipM/4h3HsE8bd4mxBqBfyz+hoE3LMpC
HPKv4OYrgzvIcQ2BQ689mC69y0HCjWzWotnQqU4qbEw64Sk5O2meGR3mGHptz6F6
81I6xIpuQvFzBTkQ/SwRJ8h6T8UWmXD2DoajAT/jJ5lCnDikuIz8P6fWLcWzpvCW
SpxZvWVPHtyOjXV9wVuP+l7/HNZB8X9a2iQ/8asn+QiT4zN35SfmdmZFIaxx8wFs
nMXdDeeP4yJbmj3eCDJAkUM5AZaSFFpUf26AO38F2jVStAiAvrpzqrCT9HuyRDfa
x676j323yXVAs4q7SeFQo/60oRydp74tx8DJkBSSd4d0IsSSVwJp6sXCJSi09wvi
I1J5fxis1prS1HRHz2MmGiCUaUBeDMrNPUFa6QMWBi969DI9s9v+qXaeMOhMspJO
jEz5nt+eVgGaUXm7rbNKAiSD0RaSvDjFUJGR0LDMFbxSJ5bSQ6m66LIPpHRFZF3N
q29Ws44KAL6qoKCPtLt1cwTnbdaF441db0Mz37Jn8eBrVTKqnvdMqvUTm3R5kfHO
6xxut7hYbp1DATDHhaM+uGOkhUxsOKwJsqv1SjG7CCEjXvsTbEhktRGKvwARlnkU
VkZ3i5PXNEUqyVbvpzjgaBeYQmuP+C0PT1fAQAyy94G8IdTd90ZBFE14no1RKw+M
V30d6J+NQamD2cx40wXSesmW7HblGm/lSH7JJy9vFzqY+qhNAf9unBB6zeMmvOky
Y7FR2dBafh0txyQJB7GZEeUWslY22PdhRDaTN+GyZ+LyJ6EUqFOQ8p2JcXp5ksuR
1r2QonmUdvnDHexkCHLGrHZ5cjLFYRBPEN+0GjgBaahKoN8diZQm6QaGAjC3RR8t
S627o4N9+zFSL/qFBN2wSpp0kudYQcvkbuO23eMmllh0CS8iwpvwxuPxoL3MpV+T
4LxMPdkzZ15Stf/Hxzo8KJII5h/3NE8xvKEhZFA5F9+GQCwnukEaCltuTKmiPh4x
fa2zO+4iEev/fmCI4LPBkdHPwp7UK2uL2DCzuEVl3L+MCO5JjYX6LMiDjhFLlO5i
vy+AZdDk/7y7NOGfblsFAOGTv32lPJZo84ANsz/uSgTtA+GSzMyy8hto4xNHpDWS
ccwQ7Z+PwML7/W+GMEv+XIRBC+J8Ny9B871ZDw8Lx8UJ6iRgOsaQxR9g1OOA1/6E
Fam3gS8WgZk5zbiAskUwD8Noxetl2wOws0HkqYHJ5xZ/892iy1bIEDRVMqs1Dljw
D/4qKSHDyutNVjS9cChPpIf7VO4dsPCU5awDpixvfUxs1+h6u2q8aLJHvdXKFfsy
zYIvhXTbXSIe8PnJzW1R865niHpabnRr3MAQ1LHTNXddurGH9/Z9FMUrFZsOFdC3
0W4pT/yh26OB2j1+si/rjFiJlTWadz6Oz33lBCrtHR8j5b7GBi3iof4zjV5IzUSB
L67tnQh8XrQ1J9XJaqodKJx5VJ/4i7tCaCtwymtT3hkSVjLRMmGcLoEQ/B18YuN3
x9+5ElKPzC5cOxeS4XvFMD3vP+tBGH0wdS8phOPsDwaIHKIDlcXO3cTh+nr1NHsJ
rBGUXxU4+Q/YpxbwsehuvgxRXhIm7u/Xk6THlO0hilbn5jYRybk8XkNvBhGpBfMj
7yXkKlo0RWL7o78v+KDggdDIQx4Dqpmmk8VclXlIiXqBOZdeL9ePYEUhZzUcdCIK
z//d2yPNqQwwXrxXAmHXQRh1IRjP3KY3KNRaCQ6hb8lLXenNoJKVD4q4HMv6ENtu
gBKljL281JM313iPFVmZCbh8SjSzrU6hdGh4oTPQy2Z9HZyXA/Eh1q7tD6VzLgNt
mYE98MyqO22tq+m2bcNLme27S7C9YHPPHr6DysAJJjKPwfNEX4Vbi2Q1/7TIKm6I
+0g1iA41IclVB05KlsGMfbgiO3x8TLDdl4yWBX6ebjYx4AVCzq9VfTMBHL5f+PGj
0pbUPGDuzIxHOjLSOnIAdMjTM0ygSyAf5J22+H/cfHLDKRLOdMPKpzNCxPoL+/a4
BP/t3wxqJ67ob5oi5vCx9lGFpB+P7llbryCu2DRud4whJQYO5cf3bqpVDllEg8qZ
VkiPPsBsmDroJPWAnoHvMTmSqz8c1SXaC/hSNVOdeEmKOIfbOJe4J8s012Na1/BG
RttV2eOCuQdScxT9oO0XC3SSdRnOkdvw9GzrXbYuCEPtBP4DjUIh3PIRfLnsqC7d
SbP8K2oxgwLriA/MiK1OlvIBFbsI/oaRp/dCV7nE9fwLG2gy9cz3HSRNVspeHA77
oQ5qqKJhCwzGH8NOIp9dRgpAtazVt2aj7IVPxybR8eipbawMkef7Vvn7c7Rve7Aw
+Aw8j8gtckEf07NPBSA/Eh2Wmdf0X+QyOQ4Dgp5uQfxiEVmLebLE7rNe/T9FKX5D
DfiqgJQY7uwpPyh0mLNocUD5wlBf8+lINOS2FWESLEYFqI+ICSOKUlAha0zpXCfy
Et3XNWN3lnOOqK0UNym8uaeaquxT94DORWufzSMWRBGfKjqvwTTA9YQ0TablaInY
S7rxPRMHjOGcXJS581qvJ3VFd06229h838qw8AsW8ALtIoPF/wUtuZSw681+rZTS
VPVnAFmXnAYdpBbZBiw38wC0bSl3qGKhaVcXqSW+tV1duqOf5DIL3WKPJoF/WUqb
1CPwuAlYPjJQzOdzOjKVg3TgBiXltjMbP2wMt50bKHOZnw77JdercXm9UclgUu9q
RaqvwxDfkjVkA5eUEroelIZ+gMRy+ttTSJ2VWpJBVrsmZH4s1DoXCaJqHKm8sf4S
IqVWbdJYRc8oV30Eu/8UtZL3lltl57aN6P0SfFH5WusQBuoJA8z+sFLVmCpWLMZh
hpXlmLCY6jUii9fEMV2QuWfuqQi47PlcllQzYIThwN8ApkfTQwiRJBQ2uRXW3zTR
q2i0byxP35JZFaVlVY/ySBZt2AMfn6UdoM0K1g1H4Pi88YKrl2WMUVuaqjhpS5+/
LNctaQMq3W3S3jwrAJJu7ux1VQn1Y+g1WA66gZ8blHFZa94eJUzgrerUN6HjbTrO
VX13Up3lmXuXCYQV33fwvtqKZMrmIYEzSgOSjZu9TJuDeqJHZa/MF7yJ3bDD0hfb
61JTyAZZle8SuGqyPthz8KaOdeBx75FdW5bhjL0bLDVj2z4t0XjMf1CwKP4yPz7z
Eod9YdHwnmFpBVeIdz3Jmi2PP/gE+tmxx9lHWAwSt5TRQpBtUkYa0uFbF0tl67eI
CAJQa5cr5eNo+39QVUwvhkX2dbwSbc1+Ea9MNYL2jELMVN07s2pRDAoV+mY4rEO7
k++z0hcnP0/H3eodW3zI7xsxDTUuHvseRqkyk9ae+KZn4zbnmfd7o6yHhcIiNTe4
Svc2mDR17cyfbyiB8HRQJ4qejaYLprZwUUhjEnrYXxkalDxUMY4UpWPuLtY9U64d
XAGm7IC4YDA+jvIZAH5q5gsdJRlv27jnIwuVREbso/CF6p+uc/SVABg/lQSLYJJA
pxMiWZ9KFanKsUL/vPIV+8WvzALkMwdqEL+2hF9BHd3pzWNO3NIFEafAJzz8mArV
laTh5vNqlm7iRnwoASdtT5O4ioiuqsTVdANEbT/Alu0ithb53BNYJAr2jc4ftZSv
84Dn2Wy4jW+BdK4UfMCHPPI48/AtfHvW4XIWI+T/BT6UcdZNZCBO8zHv6PnxobUM
hy/KkpTU7K8L3kfGL794U3hnAkHfayE/vZENmvF7SUckkirxcLE7fx05CQeDJlsd
xRD115x5Z+ypLUzUOYo/eZr74YATzbD1XS6w+hel37YdCS7MSajzn8ckCQRub5HS
oqumcq8vhlL+ZhLplqgRm3kFjqRM8JI3TD3aw3uXYW7JjMA5/kXFClO1PtgDwfEi
e5cMqT1DXNWEKYpKNujR2r7SVO6Db6FSMCRDKTkDW4u92LnuilQZoTs7ZjIMaSxq
joSsl1uVp99lmG1Z3d/x6ePlYMOQaA+OHzf1LpDeSP9ciG29Enf8MG3uKD0sE4RJ
+6Zn8KQM6B2rCVtNyK5mLdMNoaiokAg88XHOatVeyjhvKc0LQnTAPs/CJv4sqpSe
yn/sWR/c/NGm0J8irBC4YDX37fYcVaoyyp/24/LtyllcDwJzKK9D3AnuXx9NdQP5
ZAuRQXU//Jbl24q978gPh+f7s8O8RCufHhMglk/+lkxiCrDdNnghBqozL78ZNdRc
Go62XIT68UUv4MeZYBKdO2ogU3lSb543ZESjB49U5fNRAAM8gtDMABT071fRgkr7
IBiz1BId6d3mhsu8k9+AvlDdQYzJE1oYFpu34YsA+Dctt2N1kqX+bruNE/408oA+
SoCAoskGKbVPb79g7h/pTnUcsfLpXQaWU6lh+XuKmX96VY3wh79ABBj3bX9dmXaa
1YRgPugzXxiHRcADSH43Z8MdadwSyx59UcfWd7jMzBRZIxXLiScwarxBxl5L6f3Z
YkPRX8+yEvLUO9+Zo5m017Mk7EqBCawOHXG7WjlvJijCyj1XJhIfZ8WRbtlw1M/s
yqMYLojpfO6TnEuSqNtxtFoiAhPBj5JpPhTqZgpPdupd1QSwBskgb0yjkfYlvNta
BhCueNJLT++xEbaalC3LSNXawgBkRjJw9+Uq+TXDgkYHy6XIMcBGoqOALt5K4GcZ
/mTml9DE0Jjmygdl69eONpDXfeG//pX/ALeNWbG8D0NuzjFWRgie3ZBejuIGav1n
CORAuXX5YXacmedT5odQ9iWqCSKImpH6S++O/RCwyNDkMxNLHYMPJQx2xK2fuvgU
t5KSeKt+FCb7UP/so/0qw7sCvMAQbIEugmhY3DXJZUH/o4EE1QnkvMutRTSz32+G
aX9NiLl45cdWpvqO232KyPg1+2oJSEBWOOJb04LfdQzOph6fWwJ0ewFhf6jvhI+2
qto9wY7btc6wf8LciAzzgnYaiWcLjGxMQjgpivLX67uleUXy81AXkvk/pl2QpZJA
ifehiwrUnS/YvKDEkgRq8RFfEoOIMgJbEvK18sRcixIWIthp8+A3HtMgc1pYP/+9
WzYo4rulssgfprqICoFW2n6fU8jGqC0Cej5rC78KPbEcKXGAYecU26fOX+T4UMX6
GQRzSB8NLH4TnHXAI64tSIrv9ectSxEdZyzfRB832eOhXHHViG8qHr/rTuwVkQC0
F/Rts4H8O4MmGkatdQJLv0K6034BIp1uo6xPQqVpEAx5OaI2T+2lPFzTau+xD1OU
hxwCUpjwHmBowg28hZVVL4+MwJdOu9hCe4dXe7KRWicEXNMZxE1hCSsQEf6t5miF
tL26LyWNhA4mf+fD9iSQ/ouyTs43WVJ+kVOpQhy3DSjHf66wQBdbzDs7DhIFSG9T
rdy2gOHiCmiDxcy8igeT/O33PGGQOmHD+qzTIu1IwBNpvY1B2h2vkIpOUmJA/mXs
Bhj8oZipwl0+HFOhEdCdfsNdEHnIlfEu0CnaSZfAzpAqD+/fQvwv+KN/Q5a0ZhgY
peQzGJUHDO+oNt6Nw4HUxWiMlLkZVYs4TJz1Wev3Sskj45jShy0mDoy9fue8ZdZb
/9/GZFtbz+zc8gUBExuJ/ydFXr4SPCYlk6w7mxpwF59xh+xsD/lhpvWaY5Pr6/Aw
qszHUpz3tbyU4v1kI9NtCemmH22WTDr0Wz4nBVq66ecG0PXDSeWjdV2I67Rz1vgw
6s9y6PgatfBp+xak7pFp8O8pavTA3XyC+P+JsyMfdIneXr3D6UOtr1mrKGrWhjpU
KzlCan6TWCK0YbpRDyiYO414eMuwfLKw2sln+Zc3f/dqwvwGudsMyrcvFTvazqRF
guENjBKjtNT5YSPTc7uEO2y4DNq+yNthTpsV/ATGapzA1PeTE9jp3BAS5F+OI4Fm
/I5tVJQwHfs2bQ7M4lLm4stfZvSlQTJsdQFP0RWyto4BxzmwJHpAWohJDv+ZqwJx
gPWZqghu+UNzED3OCqqHNyIl9k5GZlhqZrbVQePYzAtN1zuBiDMmdpxx0WEDcimp
oKG6H8Uve28R7QKhrDn1FA6k0rioYw/rpJKuDSCToGIhCavaDPsI6YX1ddWHMpS5
IZp3mdk/fYDk5TgDYXsGg9BEt5XG1feIGFVVI78d/UwuUc9ZSJ6surAlMfJAkdhC
KlGcGPjGa4A+5qQ5y3FnbWQC1jDZYoK6JiZVswsNOrXpwbgYoY7iPwMbAnQ2Bxxu
D4k0JwX21fHeQcvxS+i6m7mUlX/QasSYCHI6rkQKWwyqqYpJUtaeA9ZPeZti/X63
NuiYsrm7xLK1Y9Z+CeGKR6D3nB6ZRxawyIcO/a/0Rrn3aozmxNXARci4af38Psma
Zjdf0pE0hSUmVbxjL+25g8MFkwm7K9C8x6O0csJpMvtinmJHh+HVOkrtWTeIxel6
ra7TbUjOV0/jHmYClu4qzxNsLUvawsUbl/mBr/GaRdJ8lC2DAC+2uVuOVHXm5CH8
jZHW/xtmJfVY1BV+d63a+K95RL4L/eLgL/WVoPPZtqA9fe0IuHgwQvjwr7D1pAYu
VsM4krt+QzH52SC0BWzwLxIJWMST6ufi91tmxCcFUQsDgjKbbdHuzOY5QMYKQwuE
BeNeXrIHjLVpAUIgOuOO8lVnxouU/WmSBNaHobRlgKNGuzOF4CfZKW7LYM3Qj+LC
JXsySnETMH2JhsTv4vsGyUgnlpx1uLuOitJpCtDOvzEk6UUj3aNSsq5+MpaZCXiP
Qi+4Wj7pQo+culjpbrqCp4irTkzuRt3vMMa380QJUha/7DXXn/vNKGRTObmVb8sJ
bacTiQ3jLRBaXcxAEVVcXQ5ORABVQ3Tju5Ynd6VEpxaYU/oEb1DMxwSGFnMo/OS/
cHqC80Az+88AwDFgxHm+mq8HNnQkI0aVAfFHOFEBjlIrSk5mGwMJx9wmmghWRsIC
m/uuKa2bAosOKTKvRwKoQRzlONDt3I8vuvpJMfeIr4eaa7WmjAMTihoGHdFP0LlU
3jkVwKS1HuJsYITNIAfblV8lFmvaF+P0c1bSpiMx6isA2OCAYyZ+G2oblSE61EUJ
o72sZCEzN8Hdq44S+xPtVOOTooKDooNY7xm97rX68qE95QpUKxAryx5pGCu6YKgN
W3cASdvzqjoNX7Z66uIwWWVz8R5cv6jju9tOemh3RHdisIfPYo8AmsOFNjgI2UxS
hSKz6qcOECLexkavKULNYXqdu3NmcKZsFOLPL9AGlVdKfFIvJXPY2J4IduddNGhC
tkQQv0OXpSu+Y592HQTWduJEmOYFq3YWFBtFYXnLbYFXIHBVLUAV0NVzTOogshXA
OwrEM7fKkk87OJNQ1aX5cfc58kEV4gxbD3OkzNLaI6zFHpE7a8MWO3vVU2O2kGJK
rH3LF/mG4W3Pm01AGQ7I6qjhx29m01T+3I/RLuVumRPeSTxqSzwc8WjEidcJBSV8
kags9RK7odDy63+zLPgBhyzGmqFtZo2jcgrDAnIgFbb9h5qZ/T0+S+QWC36bfNiw
Tcdhmc8HFdxiusSgPHR/tqb0B5CnykKEQetZbSBtW/FGqSIMA5z/SHTOETlj+ybj
psuPDoVKvZAYPFjf+M9LR/DPP4/i4oJ7hv3PEb4mhwNSt0GzqQtp1MFy3Z251nI7
W4aRFdw6CoFplJ/XiTIwKWqgWIl0AyX0LncXRKlROwuSRrG0gh/6ik7TZN+ztXfG
epwyvUv8X7CR2moe3xOotH4AUjeEDQk9uvXiyl4f5Z0zga/sYbiOhix10e4SPq7O
g9JbmrB4j2MZ5tGud+59NcG+TKWuMwI4R7O20zokDO4VkMigl1d/0xo/IEZlbblg
/nDAOmcZfwkQRsr9yGnamledd6YoYy475+UpidE5DoWYW3mON38i1KJ1UttReHFL
/XTzgaB22qwNe1pgOaUjdCXUZsm2x92AJ8pzAy4/FztQ2oHp2dfCDU+qiTo1andz
N3RcO0tqM6PTb4tQ7sW+H4ASKgTP9nOoU/diPSzuH98NwBxm5v0c4wjbif9L/74C
hJwCWN04Iddmt9pQBuQvtO9p5QCFOTHDskHqdTIZgGsGIP72/p2OtXNpgJ9ZxGsx
a4N2ZGsSXM01rolAs+Yhc+k4I0hQwEnM3PVkWFiTtYGnHyrhspyl7kofU+2Ca/E3
bvKNS4TwQJhTU21FUcbz/MM8Nk1ZrmL+B5C0Q+BB4ZgHe/JWtZE48RYeP8M3fiZc
9C+RFRrLnchsX2zJQklkGhclrNBuhb3aN2tEBUbOkAme6xLwyxaOCjM0SAEDmW/7
H3jaS0SlDU5qiPg8WAyv/hs1/uiuaEF4sdP91/8HNDyFM/n71TPLUWF6SCaWuCoR
Ag4p9op2D+c86fU8PVTAzp1ZrFKZXsYwmcRAxpnyVQMu1Zd4kjNjgzHup5fSjjp/
KLoYlg/GoDKy/8nHRSMKsc9DyIeOx6BU54hkLKx86xG46swc4A08/Fqtvk63fpUZ
w/r2r3LAju9cyx5wENJZA/D3NmmnLsCWerSPC9KGTKK5t0OnvZOcCm0yd9AI5DMJ
+O3U4UQu4GW7vNxHLzqMVVlr0zpGtPSul3MRxdzMpO6eU7zO7xBtR/oBLC8jJw90
wuDg/OZUSjdaQotIn6Pwb+Yfn9q/X8JMjgR+rLgeR3jYsl5ww5xmhNeSEOaZmEM4
lLf90QQ312I14FehR63r6I2bv+Z/1ZjCJSmHNB7ZsW1G3KIWFxJa2wj8ndiMm5Qg
WRiwm2LeL30aFKSP+wYZ11SAK4I1YzCK56Ez5mNwChtX13O+1wzRg9dhgQBtJ6dL
KIigdYf41s8GA/j0/nNRVU/v9hTMqrKgHc1R8ipPGxHM9yUBbiH0MS817gWfh07A
dYqZJXJEuHkuskJYvKeFDIGWw3pmWLomLQCQxi4UImq2DA6cj9fpPkPukbS4dILJ
+j2BWArAmAIzT8BtOExF3zm5+E3LBtDhgfyLXh1/AiHKKD4j3PsqbC6DX0+vXduK
GchwpZK91hIs+WBn0ExYhhfozrjdD/LrdHj5hOuCzPPxsLyNuuYL1lXrYbUb7ewC
fxt5YjKVZBGkirlIlY3QdyiJoDQB/VhD1oN70C6WQ+cWLTQgh0+bplxRkRgz8S0B
Nu/r+D8QUMiztxPBGJWCTgWH9VCwR01zA7bmhsyowCBcQu2jwrrtXCiLkSmj3REY
22aA1ma84PNjUOXyaFxEA2WBOO+AlR6RJuxTGjgsWw5YGtaLCEgMg8Kq3CWXCDmn
cYK5mE0nbHUXHD+YR5Hl9DCLmOmgfmksyq51Z5pFn7zbom8Co3ZLmHiQXbOhbHb7
N7aShYHxL8BduFVyqn6ZJ0rDTrtagn/gOdj/7UlxpqhSGROWrpuqZDQLxKuW1oVV
8myy0NCId5NXgROHHvqjqoj4xQd/rumo8lt7pYYSOJLJohYNdFDDVPL+MU2DaEx7
WUIbn8V4fHMfSUgpqI1nvyB4mXHEngB+qcLG7wq22MHLGE3nP5WG2b2ShExp2SuZ
6F2bNBYEz3jryAfDAn6tcI7zkF4BuNLj71Wo6rXUVcrknhatK4qQjUzibwmIaqim
t/z5lNwEYYJ+joeMX/0gf6bD5sJp5fF7g5aqmq0srUia5OD/CtR0grXRVpzsqKNp
75XJu44QvO+JTyekXJFY1FcUuGAnyPJbdYni2CQQlAvT978wa5+NCCiceennbVu+
JP1gvOOccFBsZFr2XjBj9SMAheuK3lGBCh5vpHTk7glFIi5jReZJp9zey4+P4+Cd
KIdUgKXZ0qLaPAGgfO3pwvJ4sryi3sZtExL7wovf+SOsVcbH+Kh0ykayk55y/qmb
IbphNAIMBMWV4Mi1T9xidTCAV7J7opHCCfGD7nPXSm52ciKaOFJ07J5fKypd+25f
ka29kptVAbRb/9OBe92iy1QZnHJUUrABYQHkbsm95yooggaOKEwkYoxG3tDMs6js
4L87Pi1flVpC05BbL/I6EatzG8ayS/OMldbDNXFN3pWHurzHrsJ6tSkJ/55aDM58
F3rlvzmnzMDoAa8QCRL0EmF6IW6cce8rHxut3b3ah3Yd2dsoxumA+iSLWxxkl63y
6y9eUeyOv2QwghvTqoPUkcgi/NPejxQX1FMWQjafEIOUmGGar5VHM17Oh8eN5p5I
LGqW/K4CaxoGizx0zJBJWDoVm8+of2W+RO2uG3iTKEZE2lFP0Aq1MJrb3pk1HfED
ER6S0n4DiI81nhnUwQY13uZ5EDciGsLE+aTWt2Ve4Du3XNnDM+fGxGfJqoVbUR9U
yGBEDTc5Zak6LWFtK71rFMwcCSF1fT1iimgjbgKWJv4/rm2WS/XOVls2FxugstnW
kEcOmZRDjiCkNs6PEo0SHq6tfik/DHd4stKP2blur9o6g+Cw3LB8matvFr8iF1T+
ytZ8WDniOEFAI2JLqkHloSFYvllrFWuZ8yWm76YETCn8DNnSFb+Lbl9u1Nf0qSw1
fav+y63AiUvCWtBbDXlna/UDjZ2SE+sFCNXeV+HNmSHcXhfZ0av9qWVZpLo0D36J
B+T/YPySsWxMMzHh8YSmX+88r6QXxpEsy+Xx0Ms7avsJ5Fs0tvA6LSyMy5qHAQGY
ZhlvYUmdQD2J4wdXEHelcYxrrZKgJCUiN7YX6ofUpbstJOIqfBWycAnXBxd45uUz
NkAAj/NGgH1tj3zqo40ESybuOnnETeqEObZNIwTQFRC2t9cCrNrf0AFlRT81ZwSD
SzTP+XMswkzJfso96hnm9SMjSG/l9ZgQo8FunS/7ki0R8p83aGM0vF9KsVEeoxig
UcX9emyacqTYa101SAc/YrViG4PhlF8lJSHnR7nJoUCGQRxFIq6W/D4ybQSbOWoK
auSuwZTp702Z+UknWAIpNvzWCWXmJ7U1qs1ndy9SUlOiL+vhlpiStuz4gzjVArL6
7RPJg+IK+6w4Hp1Pd6EU6CSOFTRdfpGQl9uq/JIGOqFAAx9rGQYez0q1ah1yyAD0
jqA17pql+WpN/iiO3M778Rs+JdjMdMrBAzM+sFauh0P3537OnZmKuFFzY13doYCQ
eGHZMkBtsMtzN5O8boCGDOFoeeBvX/YO5JvtxAPAQhObrRSblgWSBDYhIush76mV
BKBmvZI7IwOoOO9VgGtBZNKyAIduNIKA7ISyDac3uF59kp2FaHQf6mNvet8YeOP3
RCPE0w/Tbzj0Sp5onbgiVEjgSRpGUIi4CpToPDZ0tDMMyigsA0kRGd0+11We8qSZ
426Ggemh4W00LjwsCIoQj67iZbsIxpPLTNe11CwNQq8fKFiJyTNpsonCcu2AO2mr
YJ87U4CKcWBdqrou9Ghoq6ts63es9abKe8B5yVGmN6fhe0ugmyMMXF6r1V/doktZ
sMwWa5ENyjj+L0wAGppi9aKqLyW3sjfjn5JmRAHp/ye9KZS15/ekzk6zU0YquYFx
4Irmarju/BMYYHi3l9hCEbRBotrHxVOq7/csNSfK8PhIwSZYiw3ZxhMvczYMw/Rw
XNphu1JOsBhYWjhm3s111iv5UU0bo0Hto9k8xgPmNZk+OeXvWVDLJW2YIoQTi8rE
nWMlr/3A6kiT2atFTj00h3TwOhgUGg+6WcZHY/+khTfJcpORfek7BPl0XqWCV89F
ZydDQYmKcR8Hee8Fq6/95I/6YQCicIRMwOUCGmk4fpKVNj82NIP2pmfiRgAQNL72
MSSyGOETLqTTHIbD2bnlylvZWU+9yFcggN6O3vmrElduTM4rpF1IzTu1O8XFzv1c
LqlgNJci6B6ERoKhI8M/KIQRwA+An+6Wi1ILkH1mv5QEaGiiyRXxE1Md0o0+00+Z
ziDsATR9l37KlFYOASVNwd4lZfvB5DtBqyg3LMx37EGkeCXRL4X7s0L5+TVXS9fu
cGrmsKN87HujOfCQTGIyrc3azShhy2MxwUypL8qTUi8h3imGJrO/xZkYUQn+iC0y
z659MGwgWwxoYAszImHZj6wmHBHn1vo4OZ1gXzDFlrzSIkjG8JxKmqUA5PGo1nbc
5GFtKffkNZbHTJW3XYZ6kB5dLvc6Kb8Fn5g9WIE/sDXWaymrRBefrsbnn69jxUMe
bIJ92RsB3BsIabPv3HifX1xOImo+wYAX/ruJ1AwVC3Nm9lpY5oxDWn5tiiDPAeMx
WLPpBSgXLBEeBVrPYbmLx6CA+fQBF6qgJcxz9DS42/pc4R1MVKaJBTcBr0/QXOAg
mwMVdxqvsmhPRX1SW5KRkjhpywyspSxITOsDc1xKnsu71tSJo/Y9/PAnd97SJcL6
i/+ccO3F6ocOVqOwNpOeLRuHVqDq7sVVLSHXKwxDsspXhOqaGbADg5/ex+EPvcWN
4i5/qLsrXrVfAjfr0yTcSlMICMPpm5ESwuWMpOYEU8veaAlxIXq8jDBjSV6kB/9h
7VLL88ghZ307wwnsqluB20ojS+5yAtQ+QKh4CA6v+e2db/MnhJrKAZmCpDeqgq+e
0giJa99L6qwUZlr3wRILQGyM1Z3EI4NRCGLi4oVzsgdPi6WfNsLZMEFy4505vMK7
AjTBx0/WQgYssidU6y9hc0becorl5LV2Thbbx3IH4zkNbdZAjbGvN+3rHeaNB8Wf
ydw7R+B509eb7Hg5gjPRbB1654hOWyaQfIamqx9VBcPNNny9QrBE+swWFtbPtr0z
5ehUMT4bASEhp5e/9OenKssArQDLLGTXqcrPZYdErFNiaxQUfUKMQsheVZdc+sJO
C+qyh5lxMyZnk3pldHfo4iLTlnioxKtKylUvQYrIuBVfO+NppmLlXNZRZw/ZAWSg
X03isWoyy4WQpMFJ2SX7J0b2UbCHkH3wIgz4ApNBM0QtgaqWLPGgj6fTxjeCxu6Q
XBkD4HIFqCF5WQv+KlsbNcO+lq8VUiwjmAO/ALAJ3hlaPH9U0PQqHGfFQeGnyIBZ
9TuiHSh+0Gq4uOQ6rf077zvWKs3/7B0DokXJG5C2QT6tyFqV43e9FKg4tP9feWoA
QfeWkMJMN8i45vK7bOuO+kKUD8UYaiAVHdP9BqqSuBO1qXvkkrRR8DNHu6G89TX+
OH4B81JSkzg62vGrmo2OSpXb5noxN54l8eXjCV5ZwxThY+oynXo5Sq2DnP23G8bm
yY1ZpOPVH+UMwquVZ9HrXpPQnhYzoS4T85vR8vYmejz+S7R7s6RsVcGC0DGlyuzu
EsPql8UVFENsIKAJoceS5coG0RcbF63nTvnzSZkEIHCn0DyYU76AS3k81+HGXclo
Q6du/jqPZcXDrBnK4+7HZrn0IJAYcpw0Bda0kXeCG1ZOIYQlUOUHv4733b3fnBK2
vySlLlFpYGACUmFlnmxW4AtE9vESe8DXF1vVU5j5605R6+l1CifbpVjc63ZmnXIG
6bt34Qj5uk937M1TyCM4nq64eNQgHrb2okb/Rgzjodws+kAGjgyew0VI2a+NZLDF
xIvRPXcJDL2ODhWmWri44rhuuTZD09/Yf7u3E8xmrHJTZDZxKVitjl9UU8oy/XpT
V764XvQ9xkIFI/WtW0LLlSJsL8p2dRmUyWZcPiLkLJYsdUSTSr8J47lL6Dujmg6p
TlB7QZ5446eN7XboEvDKZ3AXEtB8RhPGWM5BAXpmNbBisOAAsuLaOvNUzzE2pjWl
nLlp0dtuChSShV7HUCeIFC2U3SjcXt7q6db72ddZZF4wlL7ya/huawPgegtGO3Ow
LNN3mFokgJskKjPGoImkcB8mQxpz9QiI8Pp2av0EBoDxByq08vHHi78wsHpxMT4v
W+o29f/dV7f/ihoEefYUKD/BAd4rNAM/bUKgQdzWASdNH63bM87nqUNpZUgtmppv
KtqOWUCIcIMMZo1ACH8oq0sHewxUYNAnlm2e/McG87w9zeQWbjirb+4eaegEitNF
t10ppKk5/YjcDrWmk8PZx4jdg8FAW7rmCIN/wotmDJ44vT7qQna0H3GQ/CM4Ks/N
tv5g5uG6RroYj/JAiyfyyn6PxAX0T3SKckqGrXI90qafQ2aUhv6TOKoYclHDrrf6
X2R7+y3I1JpPM9zFu3xR4ll/x3jyx1FDohMhpVTFe4V3TJfrApZqtPqvBCHVh24c
lcfKsm6VW+NhrWbUcIhUkbiGKF8siTZAHYJ5bFOWkbcaF1FhC5ePuGJdFiKRTa1I
agO55gchepKOzvpfYroAVWQJGmjJJS7vOASBE1xigT6W24I+TJDR+fquV8TF/vXR
vAkNwLVyZrwKPB9ke86U9xVt6PagdB1/ke7G2zx7IS81+pLknI6MsnsMkzbGJlpi
qp3lnPLbggRvpMLtT7/KouGy307K8GL9xUoXIkQibedE5BhoR6eESussX4DrkE1O
d+b4+6ErH2owOEcJGxpmt93oj0+GbQi8QfViNk4vq/li4lk6kt4TZ67lpN9ad4qb
3KoP6vllXDUJDkQGnx/frjQI4SbrtiEXMSLwR1N6jvKWjreF67t7kNPHUipxCC/d
Np8Rptjl9dDl+w3hdfFjOepADI2X4Gpdk0SuelMJQHiabFe9W+iZ9PO8WVpRyoil
4IxPfYeM3ZPv8pbjpqOuZHaU1cWb4i8zsqzLGxlVt2oOG5ZJNgFxBGyJ/n5hGLP9
j6OJF3IzOwZmAdSitDbBKxmMNvC9PHghvbXDIVQpUQZyk88stAaBAy9mxYk578DL
t9eC48jkY0b0DT2QBpyb2JNai6U9O/MZGhX9Dil6ofJSwSz+SuQI20dv2fVSb6bJ
Jd6LUXu4HodH2M9NB5/WacGWSBT5G2OSWkPbvDyds0cgZYUQ1mbbhI803aKzWxZ/
bCBQWxwD1w/IKQBGfqlq6P5mO/iSbpUjE0XSYdqCREKqrwEwb4dsziEFbvHN9DRz
bX2QVIbAGGlFy6gqTC9ZRO/kDrC9JXhBwd6DiQoElvUV1iiu+q72w9Mr205klQOw
3/y6hCbS18VWGPWzAe+zCInJvg6xJEBL5c9p8wMFCqWnbWpEWGQa98itgYQ+ujVZ
m7iDtQyxPrlZz63EswDEvBwH9yze6e/Z4dsupAMJEgcwkoYLCROhjuHf8PE/m3mY
aZDqrMeiO4rioj7w4GnDhN09egUQndt2yFF8lmnij+uiBSkrUHzXxu5uwh3EZTqg
lqUvBLl9hGXf379lWggV04y2sLW1yovC+g429kp0G24wWh6tD9HXbtHfgw95Scqw
AU8ypQfWjYRNxlEfacaOXC6/x4VCzMtPaFFaapQ4MKdPqNZZ9otOOUb+zGSwWBEC
RwwXDxVfJopRwEMDXVVrFfoH/exH5BTWP/fX5xjkgHCeXMfr1FarqwhD5ya0ncVu
oJhpEeAA11/Ip3oa8IUoAs/f5QWH0fDCmtPK4xnFe6P5ePEaolotFYLukyGnPm14
7GXYM4+kVIVkUv1pxO+ZtXGzNvPaKEehZhGTgY+Uh0p4nX1QnKowcRSKMrU5FcKE
Ifn+k3Hptsz5uTt3w57t0UcYKq8s2P3C+ucjtn3cyEISgUn5NMxuKMCqBvL+n5wa
+JR6Q8eGlbUnxKX1hKmHCSwxW4itcV7shlTTRGpM5rrbh6+Qa/fR9cBU52phcELZ
OT2D9jyWTACNfoh5au3LLWKSmc1/imdP7WVuZbzKPxQiKfNMp+HIwLksdJpXll5A
AOehE+UXYe0aG5kZ1q8G6FB0UCsLStY9QK7RbnOngF18p05jAYHhEOP+eIrxLVLI
eIERw48jsckigSxc0pStyJkbcnsceDBYwaOYhwEk/olbpzNBGSUmI3H2M28tpmIH
oVFWLaEj7Op0vW0k4AP3UISINpLvcKJOXaHmRVEtF2xK8M+xsS0ONcCgNY81JSSu
h7TdVNs9YmkCq4FJp4QM9i6/qMBWLEH4QDKc7kuiSigcZ2YD7CoF+uYXWdvkvG9Q
oK9B5OGc3SyRBp1vOTB1+pvSGiTXOiReK8M7qjXLeP83NOovXrBljRUF4Tlv6zLp
XvlNA/YTSWzjes7Rpu4bCjubQf2t8sqGweZKjpBrpBKguHeOQD7V0KSfK3vFmzft
gBNTzbvPSZq6hRe33bqn+om/Y2/YsBW7cJwFSd/wMRiX34p0Alc9F0HHL8H8nUOy
5Bc4rr253XXDS+tqxqtjZb+ciZiTbY8ATksoFyypjOtdMX4TotFFhQPKtKHBjVLB
XwFU2Tue8NhGCcfUen3wERnyuatPFm7vxueYcucmX0QGWdTpCBy6XFkGQ1PFFTxt
gaMem2IYBZXoZRPtu08yTtS3RXuIg707CJkgeK7HAX4HRlvAIEY4l0t72VaVCgRn
VGgyhvND1H+Tw//e9YsoEr4rPf84Z1MQPQIkTZmU1hJo75rHNit7nAhnjTj3LzFW
OjStmTTFRrlvsmgKGcbaqRqGtRVBYFu9AeBEojERo35fLtJsTiaIHafLsk7wS2zX
WMRLi+sxjJL1LMB7lf/g9Ncq71GkK4VmLkP8usr0Bjc8bhhG76hWpbZU79qyGCJO
BFvV/uysksTEtk1HvcoFmQWhRVKyRi5th/RC37n2ju0OsgZ/ClFvmLDnI1Sb3CqH
B8Xf8SblQO6ClWlBQtmEFBkw/ME4eQ8xGPbTrdNJWzIUmp9GeyusO+tKaJcY6tGL
Ag/VOVWYRDT759VIFPjozW1g1SfiZYrbUhLQ3SCpOns9Fh1JcoMtrxwqisLD+vlF
hKxG4j3PRc1mHNs5ClKn/vLVkgUohjkWfMKu1F7gVBgyO2ilt1w1zQzG8vBFY8K2
jCo4oU5nrhPJGhtFuq1Nglc+8XPSmIPzBUll9vFGwLRp9dz1dHgyJx8QdNmRkyLb
j9MpAadndZdTEcvkdsRecvUTeQxmeoX8AB7qwFbJFDwuKZH6+Aq1PMeZoiIPmk96
YXvRdTJD9w5qoWXJmpjRiHYvl4Ua3zvR+8ViJkU4nc+DAkYP/SJUPdrJFgF8fHP1
oQv2g5lvcdiUm/izLSXzRwpaQtm9k7nDyQRAy2MdbdWuuBtgEW92wz/hu4/Qh6Hz
HJFL0FaRZH6LdDco7w3I/Wd9/c2T33aZ6T7aa8DQ0sTV27721jZFuToD6fRMRPod
BGBrYVyWt2F2nj2sOeyBQY8Tt64EN+qH7wTIDZxiGOmgE8iFx/KBRYpToUx3zi7v
ui3OspbgBN7ayvx+hk8vxg8wMn6pnxkOoxokMRnPZcIwAp2GLIBNdR5I5Y/XjNh2
nua3hqWI0a6K1TUjQsZZ9mi8Xn0Zef5xvVVC7+cS8O3rek4r4c2O+PCrbNyBJxpq
nc7qL2K4U0UluEU5SHvk7CVqgE434/FtQR8FjPwGuPHwQAgHkOCk+ohCm89bTbY6
5pLn8xVH0elE14j1dEZ/5j5gixf6eIDP/AF9UFaUKs/1Z4gigxw3lkv2XJa/gdK5
9LZBnRhp2+og0sVtfL8fs86aDEfzdj0B/s0ORvcyCBkDw6qw8IlKEoS3Aukbv0aU
q0PepHjNCHEwefIPxww10jMhzygANH9yJ2zof24QSPFnGSslK03WgZGktVS2Et5G
l+UsocDdNNZVE+2jUNi/D9PV0ow/mZN4jUkmhFHP44TTQ5lE3yS+jGVC+Mivy2jh
fI2VkzfV4Ksj2+2tH4zyzsfDtPW5MgEkt7TKxBOtyI+BQnNH0bNksu7XYM7npfkk
one0mUNLOHoRvWKwph5skRAt9mWd4v02ChBAeN7wB3TW12kjtw1lVB8w0aUxALvW
RnaiiQDCvm2gDqU8ImeRLtXzPL382LAd34k3lqzAo7Mg6PaSLd7pGC4x0PJK6/xd
jlX6Y2Nm8BFeX/dYIdB0HTIQVoa13FTahDIKeB/Rv755pnXlJ3xj05N28oGkwbOB
R0/4dNywzhoiQgLDNJ38on/YFWT9Qp008htnvMHGP3XsMNnSAhBxiFQFbJSU5YC8
MLoY0NOSOyj8rzDJLSHcQBqBbbbjdX5Lu1LHyzKrIs7zEjZO3QehIp2O2DQIXGtZ
Juf+FMqAZxFG2w24NZHLZ9SeDkj02yulPkLxRpYgy6Q0NAdFsJ3NS/M3vpu9E7vz
hUJFIsfBdIxZ46uMncoBvlmGoyeIWAhdr4qPt39z5rt1lzQQLCSxAwIAAZDlGW0H
irO6ZLTvbJXPkL3FtwhHPQw03132hJgNrD2Knh+UnmWjab+FJ474nNjRcbPwtFvj
i8+wbSMXv8HRFFE+hln8E/83frbpTi8+QU1W6eYXiSO4baNRhOl9yg/9rCIkr6jg
iKyAJ/swmefZHjdspgULfHVMZjF78h3iG6jRNt3C3IzFUA0SZkTBZoWQyOUbjCdt
+wZDGdef5dk32WpMumQrqbaIx9OZIfgUiEePG/O7iya7zL+JQTbmWI0hqg54JOtR
Y626sBTYWDPT+WoJOtAIWkT4vSID+91chCContKmOqhQQ1IkQP0oNZR2yZd56/5i
+p89/9GIbyNvkkqSX47pFbHtjwWZiCfDIcv7mVhCSRMFgqwDyYcXDlTD70/L434q
jsTO2ngsyLMizhp/LldnU8FPOwbMI3r5Grh+Qq2FJvgbTTKVqRV6nSeHn/zL15to
L9Pi0IZuZv6bmRBwx50itd6F3aaNMuBV/ZVOP2EqJQJQCriOL1mnx02gxQv5ibHP
XoIyprmDFD0p+9Dz42P0pk9sLq9BbkCf7bjqCgQTVxlXGe7uOE7WBp3NELpCqijN
xK5MlmLGbGS1tIojpzk2BprsGd9CWb3gsJEI46WDxTsTaCnhZ6HgBhva4aH/yyh1
VWxezu8cyidPQJadKd/KQTgqHsEgXHTgOubsmBl5+M3mjiXHTxW7/CKKEpEHdV0O
26v7YxGbUNFyzJnipo98PbWzxdrabxHFXqeTZZFlX9EypIi8cl6Xdecn/B0Zk/L4
bHdBcu8wvsOb81xnaYG7dXGU+VCofHrgtGWC///KyYtDnrrF1gj8LADFBpfgBl3p
hdda/JiePjusIOEnHZZfI8/BFfB6e2bxMJQWefQZbbhOapGdrPYqrwSeDXlZWHM0
f6Td6zp6R+Oug13uVnpLQQ9HI2633QNnH2yO413EHWyeDv2nNXfGUGtZ6IxyD28r
KXyDscYBHjMt4fwgSExuJ2u9EXz9Xn8K4+OTtORSsD3EAnfs0KIcCNOAb8pNmiBd
yXWT62tSsQDYmPWD91JowR6x9MqXDz5oR/fqBybKhAzvoHiGA1e7v/rJ7PnuV7/t
ttfp19mklfYN72y8CGRyW+rpk5Ub54WJgp0O+JsPjOT83ICTar+uNErvyQVClw+s
H0ejrJ4xA18oPQpcvuN2In+Fc9BF9IeVib43RXQlCyGWdu7QLIAtvg4ek35ccMn/
h5+zrRnT0dUfKKHH/6D9/SUWNiLePsgK1lbEEWqWv+Q/gPkPIIWGMQgDEMlxt7it
a0c9FIhpnmSg0ZD6+5lcYtC3ENZKflCkfdiRv7YqE7gmjdN+ZbgghSkO5xMF7vwX
JQycrS3y2iU8GO4JHrRm4gB/vjt5tIxjCapq+6yTnyFMXIyCfVnXank9rKZARrvn
jkbMC/tMXYsZHjW4Wy9rck3hUV4MY7GTe5g0KuQQ1Nus+VrHoyqspwrVrYzVmxac
pdaa7w5UPRA3tlDeVVYoRtGSKZeVfT/oOybkZE7bGsBpp/h4C8wPXsSPJNXzEygr
RZmENpWYFnyiUYij0SXtbrXL6x5MiiKWh12hlmKlZrPsUKZy/J3p2T8qv/or0XBF
WA+F+usZKGfOK+LMGbRXJoL77boqIIz//7h2OsE3p+B3JN33wxdTx04pXvSr3y4e
Pw7q0hFKkntOe508jQia8QD6VEEtpxCPzsRwZFm1is1ccc7AhTeTnwaBzIvFkUHR
qIPDaOTHv5IYyEJB3K03ds1tKuVk7bhQ9KxR80lc0k7SOi4lbRDt5LU7swXV6aFW
3tkR1JL0pSOItbPWQny4oaGlYwEfE4Ah60gWlcLyZQRCPkeI3SyZsvdDn2DFu3OI
d98SHU6/ujRa7gGeBF4GoNVyqvyBVKlw/FVuHcTF+poxGKDEk/s09e6k5Tq3hlre
dN9x58f3YYVp8QnGz4uTevXSEVnZVXnM1t/RJvxUbu9nCJQyx+tfqDYsgj+fn2/L
BH1YSK4eaoaQhDoJU4u4Qc434PLQGHeRMEKXGFh7x6N1T2qH/9UkORxJJuObCiV1
oPGPheMCLXdNFVdlNC86RR3RsCF9auphKDvS2NKTTXUg3JjjW+MuzvRJQyoGmhRt
W+aPwDDUmR7fS4QKgc89+hy2gVlu8by+zGAS5A4yP0tgGs3wiAMiCpV+k5ipnI+b
c8Doyv5XkXrTKx+oqePmxTYQgGb/XFNmNW2MG08bZ0jexbouH6ZeVRXGz+H3I563
AO+UsDPUe3wryovaurfPeizpcI1BwuH3xjxYnhO0B8ST7eIONAO35QywDJ7Baz9X
zX3z7ihLwK0SxBwujkRMRHuPZ3TBvRYu+EpRuzUiNr4AHvmZBhGtbk5kTzh7PnHU
pfugY0hyoP0B9fuqzgulW8NKHbaquKhI/xCaFXPzoL8bjmUxz0yr2mjRwA+q6b8C
DqIKoMjaG8GVFEgfU1A/+xgcepiPNnC4AY5w8fMbv56Za3KGUBZlBr/2MGtfS627
UtTiUkMtaLcA5/bcEMDfBvSW3raeZh7HI+BfS0S4aGtWqxtOAFptgpjhgsqySr3J
C2CgO3SzcKzTw85gM7BN+85weUlWfGUeNgHFHvEyNzDIkUqMVNFg3blTtCEPnyK5
4qgvf7Re/bGUAtfG9L3yMbY4QvO7PGai7fdCzYw3e4QPqDNFlkJAPtI2s/jQUKXK
s+VRpc1vjLu1C+vSgJKWCVlsddC5Y+oH8j9MlHGr2jVMZXPR96lzeeL5LEaxmSx0
omjhUZzfvAmAHwZ6fhfBXjYNJVwtLEoL062WQOvzjs6iwG4lg0vRjOmoNNpgAxnC
pGVvH7u7foNxQlmtkXN43J9vn+fotfj9ENvwTOsi0bjnH3QN6w9GxMRsmBXqHc1z
uH5jmEHBWE6VbntGFDLytoVsyroeoqzX+FTRN2tRq0jAGEucuHf/GgbQC2zIpyjP
xBGcG/vBhGylYUIx7oH/Qbr2viqBz7Fl3PzCHrUy0/VyleXaTKe4A9zWAd/ZZxqN
v/wH/1YV/ORICOBwaoVdD2lIZWEp1H5OKAz8tpQglUAmsbB9rWZuYmY0KLO9Mq+J
VLAmd3Yt7ZppTTLshuUjuqqdWqk7aH+ozykALczRh/FiyOi2qtJvlhHQYKogwaSY
li5JvdxTVLjprFSAABnvRYcS+SEKNaBW5BSiojnvWKHg3IJxwgTWmp2sjujB1CCW
gkvFmrOTCPxTXIkU9ov6vwx1xlrk7X3MN5STwA8dBgsCysmeFDtlEYehOpatCzBy
5JGBgXfnanx6OwQ0D8tQS72LYygyWXqgv5ut8mP+w5zTsfQPGaOPhieyBojNDbag
MFMWyUHSXEMJBtOJsAV8IGiUaFE5QMZNXns/HLjwTgqYbplNAqaSzO9S+m9/Vik3
ri6fVZ4d7QbWdZ22V8zxlip9FiLRIDtlekXnn7Sq9riDOvtJzDPe+x8iu4D+hSLA
iim8syITSR4tPGOOeR5keYZNonW4VDiGACGFD9lD+vuDd3MXLAUd+6RmAiESLBDi
rMJN9BtgHw+7aLN6kDEAj4Gzb5Sz7MsrcpnojaNyx8VtmsKFMArzX4YJJ2CyA56L
xJgPU+HUpw2brWfkzndwG1G7J+JMQWmqfyuTmDwAjUOXrw58TdVbiV/KIiiIL7Yb
LH7y1vA6v85pa1wF4w330STtjJJ4Vg+zpt5OS9KWttus76qMylGZQOKa4jvkS4FE
Nz0GlczeCQJlUgZO7xG7HqEevMaxyqa1DO9R+asQa+EI0RdqWxb9dlSi2nVrqtuO
TNYcRB8slpP95R+WeffX3K2reFFCLs2/CKpE3ABncZbTMaHdzYv3MWq8B/pUdqaE
E87ZzwazGKmIYDinfbH+zN0UyocNV2EmSYfYP4BP7XQrJYUTEWx/4hX2sTAy1T2z
iPGAoENCAhSouQE9Vpg/rgax71WWQ5g23u3lYhKhTgtxM8fmGHxBBgF/IxdKT7vc
S7tfWNV04uzZxkyx3zmtOVXwprSfrCiQOyMPgwwG016d7f2GX0/ZZUPVgFQEM8oV
ag5rwtcbeQMM4V8xnilCmyxiy3sGRAY0xLY5kNofH7Bj4OwBOenbvksAEZA4H/CU
SjoRaSqVvqmHwb3FBr6/tQlsZAQ159DwlB5x+gEt9ax1scUkY7vB/uP2uPdQoZip
qyzXuYPWSv9qr8aImVc7xZvF7WwLxNDx6QsjW9Hdzq5m67BH/gv8ssZGYhvU/W26
H0B1HXanrt9kcMq+xG7lnF3I/XsTzvQzRgJUYtVwJDy6PfjHFgfnTW+nQL1gOa8Z
aJcYnBwS6bYzDkMwBBSHpJviEftiixE2TWlIfT2eJuryAS8ze6dOAqKk9HrR/GYZ
qeyF/hmtkic73UPDg+aiVaa1ckQeh3AmqUkvjKbN03iiNXEXaAbUA/7KVc0n/XoI
tNi5QIzq1thkYiA5R0ePAptUzpF+E8ApTt/eutuaA6SB/QFObNxqNb7KR+K/VYkO
0P5ApGeIbL0mxC8F+qy6h8+RMsvpVxfuE1V7oK+fGDvU7LpXqtFZJBLLpCUZ37qk
yUVcJtvNmsrd5QuE2pqzPh+xg/UI9KRt7uTs867LsXkn+qT90cLBMJLqlMmFOvOE
QrkHALX2Trede1dnzVUxQv+QZthejJ68D4CssQzDPgYXpZfEeWsc8szrMjTOxy4C
kQYmq6abJ9Nz2LHB6CFs5kJy3xZkuI8A3ApSY11ToH84JbX+I7luqob4oS+x3mN7
LCeUlEAFCUesQIfpQavSW3bppuCUJwxGYD+49A80LS+0xp5LREkvmBuxcWMJwMMQ
AOVncpo1PUhz21uBsWcyDhulAPeqs7Rid2j32V9kHf2IrURyXufQZyJWKS4uz0Ki
P8VpovxusgEdQMqAJDHpVTr6ybQ2hTyOSURj8N/V5MQjvKEYa7xnWM66+vzV99D/
abFg03hBtbuhXI7OiowGNKH/32sz0g9/zdUxmS2pKO+vPPH+MUnRZof7KC0hlVUl
BSC54CU15T0gPGhz7I/9Ay1rM0s8NKRqDNezbpryaSW9SNhvVuyvVmiRHCpDhQrr
twFcbkDR/rrSCoSob8dRlCVED8BKeUj+UQ4aD46hSWFIu4XdEWTx8P6gtF7RwrOl
m+bKdXx2nIb4QZhWuwJweLWjmW89lmv5RYfRKPYXbWnpEhaZyajyMUr1IvQiVu1I
dwmRBTBIEe2q5r33l8s4G2IfnCGCmJeisG3UGOwT9GRn3jHJu7rOMYr5kGEcqRam
r3YhOLamaaEp/gwknsXpdOlotPFkLiKpReFZgEqQoV89Fi0oazJ2WBaaagwc8e2X
0BWM0Su1ZsupNVUV23TBImq4En/MBR0Bvj5jB2W34i/6+ZIHHDFfRVf32o+BJoBg
2JZ8/YzTOPyyMTxQINSJhnmC6wpIlTH0EHmWcvk/dNt2wrTNF07lDUXynO4KM61m
QxEMZyNjbXRk975Z/scWmv9sRL7yis/GLJbbFH4rngz4EzdCB0ra8f+8goZIiMmL
/JzVw2LYyGpVfMabz3L9WkfSxU9eXIrCbJQwxSGgtdpmrQdZcVhYCuim7e3b16EM
CI/fNihhrO5Bg5dXExy/XVN3ZHohmAaOqzcB5vYsEIw5Dm/LQd33Kf/M3JICOILs
8zgpJ1tMwzYC/3FlgiIq44hWDcgqBhfDgmyGa0OHg0Im8ccGza4hhfyJB07wcjir
UquyAgdi0/i2fRpQ+8niZGpwbT7AsE0LxUP/sWo0oBk07whu4k34ewf9PmXMdb4+
jcK3YB2k6SJKNHQLw+lmlDXfxFsTySCSohdBp3P+iJa4OWdPAy1fMu4P/9p0yUo/
l4UoDT17Pyl7HyTo34/cHzezDNv5hfL36myaPzjyoczr9xCMCWbP5zcEWB3BvwsI
2wcYPtfuEAHaxzC1otqkzWx3J6f+0kbDuh5hj6mjycsu7cWtYgjQbbWpzY1Prx/E
Rj0uxnHKQcJwRdMo9+vsV8TU3RiDIgaQa1rp9RjcDxt3LmfVdGLj3pucIBXfusBc
Upnoqvu+6OYT+UOLDl3MB+XLd2Win8zV3jA1XnxecCtVkxGIn+YTGCRqWYfAbsrV
A/kCcoj4zHQgfFGBOFWTMX0asizwauefq5lSsuXLRfFV95I8qgjQe+QKjzcJlhhU
A9gwb0gayOCnOWgZbAbRxzFL42kcbHItPuvuiXeU556oYpxTZfEui3lKelGhwsaN
cfdEzc1uolEtuwLFKMR15TdQTFir+UjtgKL/a2fW9h12LeAU83f3QD7zHNhACHgW
8cbrGD9q/hfKvJ/966AoC5drBuk+DcIJ/Gat0bBRtDYNP9hww4XqkH6oxKRmO/9I
D19qC3TXh77mYClFEHF93MOmvOkwgu7LB5GAuRNNBsPFknE0WoYaobzjOdvXYv0X
AHQBf4MgANlBOWkwWQq08K3O+WPQatwaWXWoaVBAvyaUu1SIElMww8u4nlVxHpZr
MMyIXqn1/vbrZIlTllZnDMegT8NRVig/RSGIAOK5jfO4tOnBTghmmGNGZ48ckMfS
qYn7QuAFNi55IYCd7T+PDCXkuZ87s8r5orux1UFFiYnaP77r5M7puEIBi4zdKNh/
omD/6GDLpY0sup/u+zDoWvJD0eYZthguZWbAh5CFQKND/gOAGhBPWoO03CTHCmdi
sqLUiCI05L9Ng7ne1PmRBr+EIsuddINCHkbbgpcr/yTLvxO5xT8cKZij72dovGnH
PeFk+i4PiM0CI/2uM/d/afPn20gBVl19a9gAKp7kLMRggv1ZF/jbfLnWfvoHCoZ4
vCnJCwzRijY0c7qD+GKZjscnmBRcUqRtwaLirWqTEbgyM9Xr52Qr5ArELdil4PBY
KhMGNny8uwqzf/+DxUDJ82xckldvN/M1oxlOYSghluHS3LZTfMqRBorZSo7cVy/D
NuL5+JkLy2nQcpSDHOGLOczUopRV9TqB0Y8uh0OSFx+/Hwy1u1D4xQxcIxScUNC1
AnWHiUetSXUqKNJ/zAzAzVcOgOrluMRgfeRfnCdpOaQantqUU93JGrl/e6iedrpa
xOakd0lvPilnYNMx7dvR0RxkHoPgNYqblidtx5JAodMTsQhFvl0/WbqSVUkFjbHi
1ruvj/htUGyy8vlZ75XXH7pmzmtDO7jID1thvaCUuczBYs/YEuAajS3WiabcfeGH
j2YNTAL1GF2om6tKSJFXOTASgXIh/2XQwVglt8+Rty5xOdOttRq5W7+MQc0AUS33
7hwKuUsrNB7N1k0b4UQQ2inf6LZAKdgs6UjLvPqtm074gGpgpREM5KCEHy03Eho+
643Tuun1kjE0fIhxx5MAmQQDcm2IjOQfvbtqk09bcIbfqKQuGjLzhDCJyQ3A+bW/
8gUkhCYYaZUfSuboicPjRw/2zTJyUuXGob+9xVaonEcPGlsMoNBwExPBrDheOE+r
hVI0LDtHjfwur0l86Auh5bl454+2xS7sUHOSGzpIj7dqvws7GF0BAfQR76L7ETMP
NW6pUpLKfQhDzmTSFvk7CM4rXWNgoRP3aqT4aFWL4CRQg5tx8gzUF6BMWFlYobGe
aSYRn62PhYVO+fysilCr1QejXeM3+qDD7vNiIURYLPYDOUwzUo/ee+NQEUdcvqPE
801eZuy0BglzQIkhW6OwExuK759VURL2ujDeKyaupbd6Uquu4BYDun/ASiSIYUJZ
fl9cOeL1s57WeMevwuPw53bTL1qa+yOakKbIqlISwj64vlm/+1nf933sx2k2Bgmu
6Sd+erl/Aqe7v7yzLZO/beLreu8R2A65plK4J2t73A0Uc9FpkH29Db+ktFw0HGKt
HpMcQ1Df+QFWJlxmSKaOyqJDKtj54Zrxbi9FPeDxH2qSRSnqg7ultVSCiHBn5uJG
m11KT5VWZhiYLmmk9Sr3fit5c2mFDM5sDSpAq2Yt37bhuhSeSkoYVhII34QvmqLV
gerohV3NUciuJMieJ17z6IWEIYA6aUxpLpMT/IbOnTqfWtGgE4ZGt0/QOlTo9IOn
LI+MxOTDA7YDBH0KYNbHc8GlJXH/jvtuKiLxbRizOvdOQSM2gN+tqDN2L5M3O/8w
ycyKqDmydJQckRaHIj+XAA==
//pragma protect end_data_block
//pragma protect digest_block
8wOIKehG6YRZATAjphgOH8t3jvQ=
//pragma protect end_digest_block
//pragma protect end_protected
