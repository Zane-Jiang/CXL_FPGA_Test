`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
E8H4E/4kZIORC5qMlWU5uzSUIR1y3Ib9S1/CVqnXVXsuHv7l2GmkXw7npqC1x9V5
svaF1JqvMAN0Fw1PXxGKlv+tjQKPz7q2WalPQ9uIjFwQuqNCbDCWETW6AZ3D9j/o
agopMAxtkT+KLA4HbfmzH3m2m9cXZNqcyJNbo/3rvmE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 9616), data_block
6EFvpwLMnp+gVcMCYn19ajce9wYa/x+qsxfLKdS13QxTqmncw3VZ0GGFnjvoge0/
rQEgjOaZULc8L/Ty7D/UDYQruF3Fw7ljpYSlNn0rrDp0cWdh8hU9sILakhaNrGUm
/w0S96GHJK534VkGA+a8dGn96TKKDyVhL62PLshCngoh/MwZPuGFjdrmXcIufe4B
msCWV508hSFyQE+sD4uyrt4efcAEryJ6FUXgN19baz0xS0Mf1aO/8zqhgYpRxuXF
B03avIddXLQ+tw/dNPJ3hvhb/A42f0PKJjq0FPJOQpa/cMPf2XZte0oD80ZJMBOy
bY767FT4teIsqW/2hS00uaqUApsEyVgoyB4vVP2pjUqLtFPpk4ei6foiRkouwSWT
Vg9SNM5jewR3BRD2nnCHTcwXtA1dU1HC1VBG9ZrZvIaewP9cYptIGiFuYJ4isHwS
EpikVc2voIdkdw9CMj/TomnDBfewHjWTH4mdTHP7zswwGJS5NcK6Q66RNC9vO5ln
UmJQb2bcBgtk2Ekd111TyIh4tGfn804vBPufoYcBa53bsyKP58JKXPTvRVmkNec3
l7uTWuhoYBWaySY3ZW53wUtY+0n6PliiCeNk3hJIgoHnVDZmeshmTXi0VOEL+lnh
6sHvwtmc7foJERCT55I6cI0xi2iQhrfc/RgnwjS03ouW1yrTMKtSdlYu+t7dmKIa
cBVvI63cqk08R4tMX3MwRRuZ76/gCU3HYx+bmJjhvDISl9ph2WiPTqdOG3R0i/bJ
mYkiz3lvMPpDmD9e99iGLslaCRyITl1nmYjZqholG9ed0PLcTDDRKvCE/J86N0U2
PZc4Xt0znkECUKQy8ZnownLbtxgVKp/6edDU71MRVWFW9kZTrJqQOzjwFfGi/u8Y
hj8QQiCstErlzoC8Aph/T3AjvGiCUNkS0Vdao1DeK6ZausLfNLD/lVyRSqOZABUz
esM5eOs/NOl62Qsvt5q4Nv2zZXiribFBBCGrOyHhu9tHYwDJva7tUDLVr6onFwfl
QshWiGWAXkpL6yZxpLOesw2pHOZihoIUUu/2delvYyAGPYG52JkF0ubQmxvFzNje
CZI5gMGlACtJ7aKfbgiUbTjjP9UMa+nB7654YY7p8iDSd+xS4nGeMvj2jUVQ6VwS
31a0s/xbqsalXHsPWvko3pzV8Xl8uFjxqS00XqHcVfajkl5bT1aZgIyFhX6p+Np2
zeYiKYo5+Qto7F5gKz+4tEsvSHfJaNhrCeDJFahRjF7hB7IyiEUL7LK2eS1ZK0IS
e/Xq3mB0xFEqXXjOkJ7n0MV1pVXfwkX0RRNZVxrk3+AdOpvy2fmZY9hyPRv2hspz
aXFafI4cMFHdcftc1/TYBrSxmadf3j/RCchJE/8aMLKsMzPF0a61UMJP33kwexSf
UENaws7va0tOLSjVEwx4b43zhiDk4cx3CWnjvy3B2AJThfot8y1I4A64VbjiQZkR
xDGadf73LbMnxWU9QeDfN3UCnWD3n0cULaqP1aNwompLSyj/J+nErKCHq4Sin0IE
QnTkyMY6o2CaYZXTkFwi4vyvRFyTmqSJWHGHZtRYVy3JJ1zuP5Z26FzRhzgl8Wfg
Xi2OJPTSxMmYzLpP1sSrlcl5UPtStQP3P+PVB1IaiD7HV6gIXTDH/O+5WwQqHhdN
3uieUjOiEVEzN9W4YSAfWIXMBWTd31NgseaT0M7WspXHv1dA4evxJTKjulyYx/jf
keNnlVUb9eCr5xMPIw2ma9X4PqgQKwu+VPEAOpRim3fIpA57iZE6J22k2ROP+QeZ
D46dzQR3EctSkSZTJ3n7ZLWHOvLFXB75Eyd3ZA/5zZM29d+jWlmIzfkUo8eKCECf
HBNuB0uLr9P8DQyqn3TKPGG40RZTAEHfQdeVZYE3kpM6D5YCfehQ366xf8kfVLZm
RJNwbY89NeHJ3qe1c649k35QZbwmZsJqi0BqYQTz+Cj7gXxRd1aeGYptXopgMA1P
fGps5FN58q6DplPLA0b93dm/F6BTJ8y9BWOPDdpz0f71fbCWnO9z3zDJsSzCn2IH
9OYN4R0EzLRySWt91XWY+Qg8hOdUg/TzGPlW9HOyWbnbQQbgDeilq53DTRWAOnCB
p5M4c2qymyMoMg00sGBj4f9B7duyEJl09O7e5tSXqkB7j7zXSa+ojunyRhD6PUgl
rvJS/UiXsP5Y3lnvv5UkSNNLL3Q3OF4lPIYjhp+4hjAVwvAAdXeG15QqYWPKGW2V
sVwqBYj+nE1MEKQV8wtXctvLLyy88IReWMzng5wKLZ+r2lQxK63JvO/0yoVle+AG
p3asUEVmmJOMvZ8Gx6dfjxtCZBl99R/VUylEF6riGwUTuDqmDQiRDBdbkxB1mIEj
zIMAucQoHiCtPoaOiKZf+N26gwgoIJ4ZS7GetG/pyD4/alt3Uewt2OPtJj4V8xSd
P2Di2lxrTCPgcsDQjocWOxUWixMUlBmn6/wqYBuaRSUA87rxqQtr16feehyc5+sa
4k72++GpelzVDsX25w4gZwJ5vCe4T9+qU3YA3ye1KE7uM7vDeyiQF7EBaugE9rIz
xE6cCxMFXBHAQGSEBpZgCgP31f44Hf9TDIdBbx6rIxzdAyLXgFN00PmmjoAR4Q1+
yc6tl1DA736ZOIqOVK4keuEkpUcOQNJZ/HRpkbcdI+7hen5QcTf1bSnDIX6DiXtg
sRcanZPcaiQlLIA0wqUX9b4GaJEfoexSZtLXJ3uMyiswDnvvcLc9yJOMZ0UHiiew
3fViLJM707IaSzzNnlErECP/OUbpmTU0MDc4FrLbDRXNzZ39r1leYrFi1IX3J1m/
Wt8+BWNhRfW7wE6ltEY4qtv+lJTklIKo7aEEKEF7jnxgvf6s147DAvuHCLZ05aNV
WKR2EsFe2wNf6iGCOz97jozlpy1PL+70WxTpFcEkEBGYOE47U0pAlvYJyz6LhxD7
6Twaans5Ga8o8V6ifhxvf429KgdSUJuzTtGIKLhLQqbFuyP18RSIFTo/iz9+qKxP
hPK+7EgU7r9li9CAV08nSI/5LEwfYXsbsQnaLtVMSIPNRHMaQPpST9KqVcfAkwp4
WNVeRIUPXECyMF6qp7At54CGZpHH9RFsZ1q+a8RBfZkofIHeLPOkQirDVbGpcD7S
rBtHni0k80lsMsUTvxHZ5CTsotRGqIvX9nWZBIpHXQJmoYWh/Jq27WMfbAy/6A6P
65czZBMHLjeXQb3zyrHiLSJd6H8KHZ/NcaF5LCIf+72cB4ehdPhXiK3yGgxNZ7m1
AIIUfwS3jLrXxl2txCwocIbK9brW8iDj00DhPZrDVnrDXVZGuf77mRbL3XJas7dB
/jBHgWc6uBAys4QA1KM2YL1HiJ85+SwHhnBvQCINSOoRpjEP0kXrinGWVzwNS5de
el2n1xe3YZbuOeMHQKdPBSTCLiPsNdLOj7s5yPSuWjNk5JFaLEj2FQya2dulQnaW
yDvmg/DFDE43bEw7WxI7L3gmx/IsJPoTFxB6/xgQShtgEkbgEEHNJfn1l7wyErfp
x7KtmpSoD1Nimb6C3sND3g43YPbJ58jzkWdqN9ci18AicqBYmZZDr2MMpLFIeNE4
R1ka9yxOWKYiT+cQBkM3FMUryWyjzxx0OvM9iAu16eenXX7b1xVnxat8KKxy3rJR
ZynUKhBkvXkK0J+k4sPkdMrI2yAvdva1mcdY8W0SLAy5RToG8PxCS7JjWaM5oXOt
k8nnX1PBc/z/YduESGA5hI4onOQWp9WfxdMSV3AjF0tt8b/Dxl3+l/yPgdWN0RZ4
5R8MxBRIep88dvINz/WD0dr5loNDVw+IXpnAZcINmpwTpC0Bdbc5ti+cnNStna2q
vehSmC4kVahtzsIzaxLzvnnZWkCtKUcm7oE7o+JV8ep6uhr9nxgF+or96uNN8OLi
X5I6VQUiNFSwckPs0GmR7wA1ndyn0sqDWERfTtJKOOCrpQA4W0gKW62Z/rb6XRq/
JqkJBpWiEhminxeBLUZHM9YzkGt8jgKXlX4LPyp3kntFBEu9MMceELEosFQrr1w+
SmyznnWtBZcRSUbySC3cylgxhqxZEC3fGeNH8FjyNQmN1a2RthNLsszEbzOjHDtM
BlaEp3Sp3eDULeS5aKArXu24OWn+iqrg6xQ61rVGN2Jk+ycwtRycHhvT/Pf1Vwgh
brShhQ9xmvOyT4z6MkShDXVJrAIAihz9daFBwlHHgpn5EYsIGyKqXnjAnF/J2u5u
YrnFWn2mfgI4rK38faNQco2eMHPEDkSHURbecFN4OqhSSbCOqkT+/la2kO1dB0Gk
vC6jU2A81kZHB8VREiN+VPpuF1/eIzPuuWhTopEHVvqlufIf5hv+svOGv4QiWuGj
OKx4igYlfZZORcRRX2ocztIeTY5gWBtFfjzzPGwrcA6AamQKykBEIZGpslBkSi4Q
uKEmgMX41TIcSwrzDV5sHAQ2YjhthTv/c0sNa+SZVEtummRf98rJtJbrMvumdgjf
UgnMfI/T+pg9vIn7CVk9iINVw6e5W3qo+vs9e2q7+iBy5y1DGFapXOYaQzomeJnT
ILcHlw9v4Ac2ODdLFZUmuUvbfGs1ti5n31o4CMmREhu7M5g023BFUlSFRd7sJTrb
ju1zB+cgZJS3UsYCafNHgLAFPyYBRuz7KV3G5fe2NiBwWKh08EeGzhnn6Nc6U4gD
oqjO+SS1Mo4teTJ6MXjnSbs1tRbv/nMwr6sXrPpZg4/aHfBysrv8McqFqkR5E+K/
nWgfxMJEUn8ZsxS5NKQQNGrtbQm8kf09pFtZ/Wp9/SZVoxaBL67SJmIMokQxjkEH
V7+ChYRc1YGRj3J4oyFjFP6Gmi78h54P4uZy8xMnFduVmce58e5SEmp3E19bmzFB
fjjV3LZXU2P+TEi6ZlUMaHMctd12dtmXTMxNbBjf2+SXWaErhZJs1G0y9s0E1lWu
s83IJBJQk4mfnNqOjPJyJF/0XFICRW+XYpolCVsCKni073/5JFJm0LoNmS0Shsr5
xQFVb1ZKSMK70kLJk1OI0nsncMUdGWaK9xcgVs2QTHyzPs+81aXirlyg0elwChCA
/sn9vu+8HRJnChmVmjZ5CfmCsxaLK1ScyaIq8Q+86e/zKOYsRVGSpVw9PMEDhpOu
j3hibxgdQddHZCXgMBNs+2iFXfe5Pdn1P95vsD3VvruWXG5DMIbMveuBGMoPq3Zx
N05Mu0SCRd+AyAWCFLjfYM3whcvDrRn0eMXKapzLRfO3YPvtsoqSpAGoLUMuX8gG
gQ5SnP/TTBeDFo7qsnWLx1tjZKLEFAHvjAUhZ8Z23/4bMi6QkoKQwZarXezgupEM
NHWaj0E1zIErG/h3wk+E1Mwoyg9p9u+fGjSJnYR7cyPqfD6n/IbfW2WeXWczk4Po
MhJyqRdgFOCrStBNx4xs4LCsUxFUADIoeBYpJNxpjg4kGEqb8jthzbPc/T1BtEBh
CQ8Y8676LmNuGRvNQr6XSWDMcfiVGaDJ1RwcJGjqDP4+uxSI6l3swsFw/6Te2yyx
WqEyF4sFDBD1iolUqiNiWYSVz7PsFIJun/3i2Gst5jMOPBC1iAfmM2Yo/G04MBXz
6w6WWKXw9JtnNzK+T79WZRx/EyiaLjlhswIfKlgFLzKG/L7B2YAg2iOEYjh3ZfpP
K2nN1GCDeAly/fNMf8Nn1JjZZnAq0eWYU1A32HeJ7tQVTc+FbyLpMyw1Je0MuGDX
hzH1EdrTP26UDXtpXEt56DTMg6uXzZzGq9fB9VHTGMpCbkP/jmSzX8bJj/nb/HWR
C2GV8494CUhGmrcRASfaAqpmHCEUP3dasMRIld8nxhUCwkmNqgF8+0IhsbmcvrXT
Vn7MRZk5AWTsXQC6ZHZyrriOx7Sgq0gWsNpmwzZhSTMgjtJliIK8M8gZttlL7BHs
RmcdLtnSO2oMTR/CqZwrgNbZPm9wAQBasL897TkP7aa1PdTUGzcRF2qbfizkNeXR
dTD6eg0rszyCEt6i8/Yk8MQRxDiKRSDpIQqIp9xZoFLbZANxCdADr3IWnfA2Mjy9
PtC3/PG5Mtt9Hn0tVO/lVKvlMrCWoxzJrYg7cAMxeDvaYq29F05T05qaeelz35FU
T+ra38ouppymZN0PiMnH2ScLMe5ynn8EWDTrMdecGgNEt+HKbu8QCkZMD5+YurHQ
Sh9MgAiRcp46fm0CaQFaIExINB6nIgJKq52qiSbbzzJV9jblNCSbvqIxg2U6wVBD
gPUnANdd/+BSukg5Tpy357202lxGWrgdjrI+JPfrhmrezyLSC8gn9CFMGnBSpyrb
obQptkJX27F+mX3PKGFJu6XQLWUdxK5TYyE/Rdr3/KD5t6kMCaX+xeWDzdnSR/vX
ugVoEffL9c6GY6Zsc0YIKV4N/I4ae8TpbpflstVBZLS6uu5tTgvPv5qy36w4BGI+
EPc582w9CZp3I9iaADG1P9G/7Gay8TniE60gtiluNFWYNF/2TvGAIMExf+6GU3Ms
QzITMvIUYGatgmyajm2+IktGNrHrcIsSUQF0ROGD0oQCsq6GtPB4B5xCAoX8J6Hs
usHki7shFSVd1TfHeovTmlMPFt6CCFEFoxQ6bbVZDa6+kpeBJs9lyxDPtlCXxznE
8JumUfa0DMvDXUSKhSnCAgv9+MlctZ2+RIs1FAVs+Z4x46L1qJd8Bl9LGnvFuNu6
Xn+kYySWMQYoxHE+a7vUmISTlQefjU4d0ogI3U5ba83dqNV5D5UzKbZtMlEOFmof
XTZ4wO70gTLpjVBZ8X1Xe9qEdZDDSeXuu1uVm/dMPVf8yVO249F0ViY7O5YwoUNC
zsvl55CWdStWWbsYQyILluB2Q1V8d/fhzl3e0e5mfllpEyzuFF2HgFJd3iF8eCaD
pHuE0A8Id5z0AL+YwZMQoehkm6IIGP+nmcU7KzxXOopoIDYc2c4KUilmQ7Nu4hAn
hg7GRJ/BBmBHJy5PyaPjrYte1mJnj2b3akYruwkZwh/166Zje9K5nKARxyEpbjuE
O61YI0/6LcUfJpXcBDhjF2HNfQX+8Cmjdud91xnaFOFNWJ1KEjdSocNCZiM1bq9k
41GBnPrGtowiL8VEwzr32M8jt2HRlX9Xm1QS8kzok0j0iDfqwzmDCFplowSWkHZx
hXToCqbiLnAWtV301oe9bC77bT060oAJeRcyFz82LAnKdDyzqcoecsEhEODUonh+
y+UrE+/f/GlCp8SOhlzUbYyNu6zTGJsaOt+j+4Fe1VpbK4kXnKe3mFW1cPlWc50W
0JNA8iZKCqvQLKdcl+fngIsQKWojlB2vyr6b0HaWy1fhGIwZR87j7HSQ3gLjL5ib
tJFQl/TnZCxjfc/ijcg4oBCgjXjIuVqWyByz+HjfNvrpxtKEDiqVNsPJ7U0viGCg
nH7e5TJ8tUuICF9ldWeT4hp/ZhiYUinv5kyUM7kTYcm36ouSYqAKKXShqHF4kagP
wol42jgAjshakg9afhtsGhLJE3awMKRYMiU2VP14qihUtek6CLgX51IXUOaVwJ6m
v+SuZztu4aUnwv38BnwOuJuZKRZRE3cTndVAP1eyqAMBv2lwm/K+zuVHLBJQJDfE
35ct3WwIzOZNhZZajE9oO6SGr+C+MXCv6ElaYGzNjBwaVEUHea6fJHxYXg+HHy+K
p4cF4+rITIOkOt+XiZQuGK6GRcX37z+/0PVEdXaZE1b/C9wGR1WjDgCvWgetDMwL
L9nU5JCIT9j3zK8qRIn2W0UOoV9mJNlMhOm+v3LWeGdt2jTOKyahg2GFjV38K3E3
FrjY6oD+lrxfv1vJN5QJYyF6s4sa6iA6eBw5UoZBA+D8GXCSqMcGXj2lrK2d3DHn
3myaGVxMaDiy02s6nwvkJ/v66ZttTYcvGVexCNvndVxvLmQVhM9nafT1i/zHyCXn
IfTkFCx+fchBWTN38x+OQC25oa5HqLh6PUZex5IANTEUZxwKCy5R8bgAuq4B0JoN
lXkP7r/GS3bouieGOZomZtqpl4SZWXwXsqjqqfjsx3WMxDB+IlifOPPEu8Kcxkdx
JS4/0De0UAzkC+zwl7L5PCfy4FBkQH6oioNkOgAGkdrCwfVAvKMgHChymmU8cXDE
xM0zWZU4Hdlu8OICkLZw8bteW+XrXwmJnj1nxlQyyzYpDuSnUX8lZY8xlGlmljNm
YDEvm5idvZJwSP5LRDESJxSL6WLaq0ZVX5h+4Enl2vsGR28EY17u0KshyPIw3aHR
tJIZ/StiSRmb2sJRAp6tTxioxaWiBvVHaX1msBg19DaKotf5wbPigf2heEb8yUUh
5P8WganfjyMZadEqVGNReqaNtdjE9WTeCrn1HPCZeg6niY+UNd86Z5lFe+W8lIY/
/PmO37EKrbpx6HTdAN9Zcqwzet8Ch+heaCF4BaIcR1qsNUtQ3dabIFVpqfKImpql
wTqWC8wuJnLvgbO24lYZtFxtGE4zI0vEFLs/TI81+sbyB3xypH9QgOD9zQDol5jd
MHlyH9n+3/2sKNJ3BYbws0qzIkgKpUZMzs1TPEgYcMZE1S2mDPoKazuAz+EroUcP
P6in89Ik/fKGGtHZAM3ww3DbTuof1+7oPtaAnAGHglScxTE0+pOqiImGM6+nDPVi
PgGRGpuyftQBsyib6TJpDQToK2RkvvqaoaAfXYP4tjFDon4Pwyr0aEk3eHHbQq10
fSAzflRdRBw4Jl+rviXj87/X4ZkLkosEHzdWm9TzdaGNMj0PpzdtGS8EQDi/9bD1
2LwchZ7Jd8pa0GZLweCB2QRfq7DC1yBg7kpjuGHu0HhBFfku/PSCuEsh0GUQ2cd5
XU7YqUbgYUGZFllZxNB3QqQs/7aKPmq9fZP+IGbNJ0ADcLoouxblpYGAMuYyMQe7
K/G4qOV1FkcwvZWeWBQJ/2Ld17r+AjMqKiRJyCeLmPNCXx5ejU/0OgfMXyW80Oxf
qSZL7fzFspz1WQJetiXdBxZMzvRo8PA5qt6cEf+A2wBwUbTYtgot0p1WT9NqE0C9
QTqaiGbU9m867h3MP4oITbU1z9HOszYPeyW0lF84U79vAc1/aHwvm3deJ2Ct46zB
8NXJDDL+KwA77/gTTae0Vg0pfLKhWLWJkf/xSF2tukgVL/NM1pbDUD7J8G7/BIT2
XCwoDwwgsdTBT2ReNHsitPfKxrt6m9l7J5ysWmOX2B2nT7UUHhThrTyrVTeoHr8j
nBVXECIUOik9P9SP/oR37/n579h2GXIuRmJc4eVLHkfdzrXxUoIobbwzP8Bzn50L
ev7yj5S9KdqQzlA82Atc0Ucd4jpqFArhVbeBuOnNmXL6BNG0Ki+XWlv0efycXFwN
EiqF6/JmIArcjGwFJ/67yDYDrQVlKRvJ2MkzoYG/ZkJrSBDHslW4gDS4k4o/YLOa
VAu8DvXw3GrbUKUm0jk/2Td0aBm/KN2bd+dEoTISp462jPJh9a6Z8FOpOgaJCeXP
4e4gtnHxM97yi0uwhtei0eFHuvqVfwYXfHwkNHSFMuoYe/IAqn5XvfM/CfjzYEPc
gKuieX7fh+Z06Vs8796BvdOrCTMpVw8GclRBxn7twfSdjODYI3EhLa6+3oJ0FpUS
FT8VKl1Gnu5SebT4J/q8i8GObtFskmcOFae5WPSz9UEoARqXnzX8v0+lLT7mLd0E
a/aaNEXehrfsQrEbtts5BVIbxPaTmSBbnCDaGmISG7n2IKFckXCmBC5g3Z9OeRh8
CDrltCLu9FdpJKxwMkSIQUADgf2rYVbVSW/LUB62gwtFvWmfFV9bcCm0R/VZMbmn
vepLZRjbFS6alVMjZFpHQ0yr6aCAz3tlBNq+YggbyvDTGwBFj0v0KsQVpTxtRopo
Zph1R+rx5gRRZrDiaCiWqoYpINKEUuQvMUhluhM9zPIlg5g6WfzC8YphHoyFQCu1
h3kip/IsukpjcGRdkQoSWqjFrmgGTC5lroqvtZasY7KZjyYAjp+qolk8ORuc28TV
l5YGmWg2BGLy0Hjp3w0pUbU9aZOs2kB97GOsT2LADI8oLzyBm+fh+UnmpCoi0kT9
uazaNI5iqr7BDh58d/YtqP8hxD3rZKQemUdsLLnLxZhdDTpJzQnbO6D9G2+C1MH4
fm3ntH12mBxMOf8vELRry1Y7J4Ura9QSXGZBypuEZKq7gpmpfQrk2ds7L+Hy+I7l
LFUF6D8nRYaJn6oEVBNkwJNUdbqN8DtOFWEiv5OeSUd6pkBL/6Xw7jGLlujh/HgX
l3VGhUEJ7Xx4XDRo1aSJRkAcS/4eg7yp2qs9lPl2FZZNUzXwiYdDLlBibtWnXROQ
7nuJz2lO2W0Ua2rvFCzUub+oTTj3Vp+qyT9xEyTeU3nV04eSpDxqKktRcjuosL9P
Xua40aJkIQdYyg/HpvAZkoWHcj1JacRBOtrrchkWySl0YLpZ008sp0nkkbv+pyfM
D//ORb1MIhp07zTx2zp7hXQUvj7w4iTgexEcR0Y0iZ4k+9Zw5PIkaGh/Eolxms+j
jxKMW/qN9SrDST1VTpNOFr5DBh4sXHu3JDkwDZIqiw80WFCY3w9Tw1uHVu9i0AAk
m8Hv+oK6Ea0AWYgSd9hWcW2CJoa/yksPBNi0H4OHr8a3THfGu4G+GSMKBxgn9Wxj
n9rlmGD/IpkQIV+WJTKUX60Y80m4yRCCmebpzQNsyIHD1TetmaIbmPNZ21XLEYvE
3x5BGBlU4oogwgGvlv2kmj+0X9diycl7TmNUbmO4DqNBF0Dwlnia32Z3C3vhXCZ9
5Yf9Kg1YdQTk5XpwQG6UQU8tP9bNBek/FVBhgaiWVyKjmUbuGTTswt/5iZOu0X2F
HFNYweGhnb4FU4uGltANTDhcfDJ4Hn2wfebQ6Cauaj85xRcWWBjQKmzzEWr5/iib
ZM7wTh4e8CrBKtuGcJ3xNiO6lu6yyZ3yyz/ToifFTnmPdBQcNXHnDM62+LosKUb8
bRNUqJmGovikOmEZmi1nJTyb+x/8PZkpyD0dl/JzF6CXXv6kvuB5o9JDIGnAmGGz
VWzrXbxlFzy4MlQTaM/6ZxDNSe1ni8gMhQvtt1g35w0OluJjhpiWGeDuRejdQuf3
ctcDSWACTFNkVZsN92p28TUuo/gO3scou/moD0fPRgXsudh1uJhKzd8Q3GEs6aHa
w2Le52Tq+J5fJiT/sRrO1CFCeearl8U3VAOgSszfm+4x9KhUEf4dqzJfnhx3CUf6
dpkQl7wTEkeU2ARqlzpenHMkQ3Y/AmQayfQNKTcQWwEWeu3sSTmPh9ZtxAzrjOZ+
QFdPDrw87Eh3tsJMWn9QPVYacPfBojZyZ8Wslw4JS5vik7299RhBV/g18lLab1Bl
v2vJeCplFa89oz+pnpD380zjHeF3p4IsPYr3kDXBBdYcPb9QFx/lSrjrt5w3m+op
NXALfVr/lfYMxXR9BuxngLLVRbEkbq2uGa90MkfVbve8Kl8d3SKjKBCl4aX6NJWT
Zxs2QyNJ2t2RTVHGmjf7pli1I3TBZnM7ogOdUiXG/FjRJgc1dghXN7Tn/9HIe7xS
74DRp4yTtTlwaUIZ9cDonhuRBacfMuPI9FskcK7WGoWtQvpaK1bMdb/qtqU3a0Wi
B+pVaggx+loFNk6dkzqHL1nQI676khPcyZE0Yd8ltlF/mh75Rq/WZJFKjCp1MIJj
dxgXkj4ybtF6z133/EO17DLiZNS5KiRojPhhv4mGKdWuD6D4CC/QAn/05f13te8J
E2f2tr2OFs6PjidK6ZGeLk3gqrbBT1FmcmLYgfur0c5X6qnEVRkFqYBc0GjJAtLC
O3bm6yGjbTa+J6EbCm04PPEql6SwN1v/SScYSJT6lybHvbrWBkcbcLfSsZ6trkOQ
u0fNpMqkeJEOrNf87tawikfhuIa2NCcouKWzYCrfb+lIdyE2/1WBCqpGUwxYDs8Q
44w+qRVu9pJ9pf1Dj0LxMcTl8zKeHV/Japzsv9naDGn1ppEWM5tQRQSnV7ZL9FII
77e8fVt2FVtLRRfV12H4/+D5n8FG2uzRbH1a0lkakbvt6zO1lXjhnS7GzfgIbyum
W6F98YjFPk25zVhDCky0VEpOhOYkESqpsXZgZZ54ddG/+jyk2Otx6EJlEec42XkM
v1ES63gHeYSzuyqbjsoNSTz+5EhTlsCDrplpmWq0V78Q+lQLgcoMMTuj2i24rIZb
n6xXZl6CmLRtg8wj0Uqed/8eWPb7MNXnWDxmYVthZWobilvL7NcCTO+kz2j/og0+
VZhtdy8SKWQKN5ubFKGnAcJdK7j+kWCNuqWBiofKZJKP4O7Y8o3ay6abZ3jUOJIx
ff1LdryH7QXbACHVq8/9T8woNo0qqdkAK2S9e7K/e7whWS/Rfc6EDUt69/w16VG2
zRD2eXiGNfSFNdK9Ggr5lR4sq8a29yLaDSVVGnayCZW4tupd+U9eDHxnukDMHSAB
Op+RXzKwVD8CxJrc2n+A4BECLW3ckmdpwa65ad3VlqwOfjNQOJk98+WTtgkahD0P
OHANFxYM3U24h9hKQUaUs1zMGR8WvX64lZgiftKxg2cz6CriUmUwD55RsSFlzYEl
msuUJFRyzt4Y+AUlpsTDLYcupDdgXerLi3d9eqkl1RKej6E8N75MvbnD3YDmiPgb
T+64gpM+hbbk6OPNl1M4reForHN2BSt4AVfpbRpQqAxVDFaFRE7AUuOYPUx+/MJk
Hc5vLbEtEwnEf7F+v3WnOG43nd3y/Zdw9ECJMgpV8iMvnglonBAh1M0eEg1mnQsG
N5la0p/SDQft3Lzjx3Ok7YY+osjW98XKTtVNoPodRSl1sLxE/xKQ4wtzkOlJUc0a
upe1jJ1hE+lHepw8rlzFSuUuG36jgAGMf/KjdpymUZgVjRP81fTeoM4GkTTBIvUk
pqdEAh+pW4kN5xrFGLceOQ==
`pragma protect end_protected
