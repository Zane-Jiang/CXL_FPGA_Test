// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
ZVlk2h6tXverihGWpVHzUp8tHjT6Qt6w75CGUkCKfo6nIlp00vgJNmkOOX2wHhPR
PEspPqStJPt4nm6GDKjv8Pg7XITXBUWodjZ/TDZcilvpb3loPxINSnX7oxrWk0RT
nPK8TRjJD1QG1iqbPeH3K+u6NXueuHY69kp3BOASpz8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 20000 )
`pragma protect data_block
pKrLrEUF8qrCN+69lK3IbvymL15EKPhpKqW+QwYPgTJfzUD9AfxGIe8Wo4200TuQ
BJ4Y42tRKY6p0NSENcrjbdf+NvUhB3FTnF+bSWHMgxOEUnasmr8IcGxY9HAkOBb0
veGGFnWo/6U6PdadscaESznXARVmvqwWAkYhIqjVl4KDlpY7NESjKgVAJStm/Y1p
qAcltZZ7FK3tqI809HB5kmGNJC/IkwBpWgV7LrIzFW9boFZaCg1GgwTszi2DktqK
mCIfi6R3/JKn+KNjmI/zqnAsMBRlSrKeYYLupWd8YG0K508uHYU9/HekuLmvRKWH
Te2CIpSPR6tyLwwzfidPcwnuwgTIjbbyXKcSP23nEL5CSJwee2usVRkfOADxv6gz
oI0VdFkbU8JZWMaQSOriwuiyynbwKEzEhB2y+uvnlVpzOqSn659MU+l+anwc07Rl
FiWebK+BKevxccyJsL8i9ljFcCZnbwu8mGtIM00tSBmkHOuAdoyKjMdUiWpex9AW
Lw7i/xfx1WDNxKfzVP2N8fzn//1g5IT+hO1XA+c4QgSO4/Fh1gDzdktUwv3XO6dk
tiiWR8RcfdXnCL/jxi5rYhpTYtVc4SX0j+nObeciLlH6++WC6Naek7Vc2EZb0vhH
tPNYyU2HQIcIQP0kDhGo41DrRm/yFBLE05ip8JdvmyEFgNV8A9CV1+bHoPiR9Wn6
Qj2oMj677lHfcdLf7QpaVbEVIxoWsnXPfe9OshrCozVHrWVL7iOMf2oARBr4yOs7
20kMCTqgQiZwUKibpSaVOE2QHtcIbqdmUxh5x+hcCzoONoUNH+UGNOiCu5lWexYa
ZxL1JOeI3ngqCPMYICyoan3fiNS6Sj/n3CpzgCDnxjy+WGGpq9Bksk1LmGD+NHbG
r17OlB400ThLiFPDvtjJe80b+Gd0Dw2HlPHsWa8XZBb0h5be0aRljDUUeMdQeUEm
2WI+VEq5QH0qTpgm8CQeSfwpYisSK4ypBTckhdu9DdGgO2u9UUzHJPpRE2l6AqVm
VjdR/ppewojsmeVBeIzgAiUYM+KZgr+2Fq/+vbW26R9AbYRwOikpynTJWvD85fz9
AlvCXl9AG0hgPJDWH8k3gI6GK9phGrfxnC7hJ6VmF0CP9lLylSwtgNZ2VOTDo+Gs
PWqGW92NExgpLsATzKS1+/2hmxVBqtbhlgcO22/5W13Ru80thLol6g7WYmHa42qf
49kDAu4Q/TCR62/eLI0lJ5ZmN2c3RajP7Y2y8W6uqop+Y2Qr1tcK+bnVmNkpds3j
NCrVu8OJ6PZwewpu0OQkCFcZ5tCqlYXYS/A8q/kyvuvk+t4pb/iXfUM3zZjqV2Jv
FNL29k803JzcC8kMr+n+63whC5eIGUAtTHHrVHDQDNnRdi4+I1Jzq/Q4Cin+pHTz
dmcSklnhtFU34NlUwITZ4eCr3gP+hvO/JrKdtH2pSIOUgPgKAj2xpOhVAME48EKJ
r1hvTshu3+OhdqnurOwM8fnpSasgsIiS30skmqWim2WnK3hG5/P6yG3kG8bFqFtK
c7B8kV+3MiPXMa0JEFfBaRpbgpBrUCRkfpiKbohZSERvS16HrUr743+qmHfZpc03
85mlKeydp/SLSsPNkZc/WCUpngYuMl26Mvxk0c0M8hZw5YjP1D0Zz1cpcNC0DTsD
XJ6XspR1aPeWPVP2EdJ7Or2/a0OjKh6oI+TiRB94lgMUFD94T4M4TETtYGXjukDT
a94TXWjCF4wfy44n0raQfTFbrD7HMoK+hW0pYQ2H7xdgW/lYVSZtRVCflffyZkea
JDeYqdvOzbwWx98UXazRpI8lTdDDrfcYYTkuVpMIPcc9e5n/e6UI/Ri4p8qsOrjQ
215vPOTR1HIPF97XIlpHcw3U7Rc197NTBhj4qmFrQDe7Eur1mMXpK9l5nesEvtMF
PVrElsBS47WmJm/qwoQ0b3M93/YAvrf7jS4oX0ZEofvECzuKKnjk0vQ/z/gggqlv
8q0sW8giicxc978XR7PWpY6L1V8aaZ3Myrj51406vqf3MvR1EYY6ICbrLGkIsuXg
DxmrhryCaTz4YMJf/Ly4UNw9YHoKTfA8jb+tb6/MwOYJhd408pSveeiQIPTQA/pQ
ZOf7MnS4vi5WB60egbbRKo65kIamEqfSH44j33l906fFgApq7J4ksTrGF77TQigh
bRgHTxrLOOluk5fRrWLZYHKPmd4kSZxbrHhZ2R9YmmIsVXX2S9uCcNehxGugAHnX
sRja7FfeX0IKTVaYH0RYu5ZEFbvICGzcYsi99joiO7ubTCY3Qtu0scgYABhkuTzR
O00I9Ul6929k8UrYhSrhzwfSc6QeopMKDApHEQFQnGSTlOjRCNpQ0V1DCYwiDF+a
bkGNyhw0yCNZgw+9xfZ0pSeXjoOjkgnmnGXMH324JruF/+F7OYKmiEbpyr33i1hj
m+ExHFIzNLZGKJhPoybC+wo1Bo/kg70CezeT7Kq9mC8oQTF+bucVs7uKsuW9fv6I
VCvdOjRMF5j5KpfKHVG3TgC/HplwaUh/5FLlDnk37iofv2vVfiT6S+xUeQ1ZH/J/
xeMnIwUQvmL5BGY01XujHiw7ggdTi4BnpRw51imtWd7oC2UcGmHRsBi26ILtpEoL
TM98GF9CeslTk992WtYzyih/l6Hf4wHSrhaC+zv4HBMy2eorleDW7rJGFUUR3hOh
ktjczI9UGpliRPKMb+G24RXaX2Nx2jxg4TP5DPbCMpHks8WtBXrLemjTbM9s+1pY
f03djpHVWoM6oyfESjchS6FrzDFeQSYjHIQKdU6ATVuryZdegfxRFo363V9E3rZK
4NMAJ/B2z92hsWA66KEN4jCh+TsRfEvrm/HpJTlZb9tvAO5NwTieEwVM14tbCtlu
BH/ojhAVrmVgPzd75/Q2wTFaqzpdATFHtrf/muw9KsvMIgAWacM5nrhftHvokDEs
cALn4TEpiA80UgAxwQJeO+agGSzmcvERX2/xhf3A4FC+q1+++J1zI6gYAyza7SP0
kKFMYKPuMBukgnd2JqwrqO4ov/KderWiTDZPG7qkcG5WDFAe3aY4S1kqqSWgNRHi
PD/8zaFvirTOTd5Fjls4RscIW0LzYQGkyXXtM8OAnu5XDzj9nG6vBH86CKzdSBET
LDsZxb6+cIA853lkpd8lVsQtdWeLdviiQTri1pgG85CR7gzdOVJrgT373NMDknd3
jFzQgNRWz+o36zFgykf8unzWE3wktb1uLA9UBjMxlVnh2bHwna/pxgNYxS516R2R
s28D+rMutAZDxNDHPJA21r2c9TOxLiwxPubkrMK7870wMG0d1qE2j1ViAHpPjm1s
A9ooaogFipN7BzY/WT5K/5P0jplL7UWE+I521gqJarPDclvV8Irtu07m8K1FF6/1
zVUiol5PXHmN1m2n2f8V3YOoRtaMYDTqD5jHhAW8RedHieXMUmM2RxNBtZRQXS0F
tpIKpV8I1cGA67gB7KqXMWlLXse5CUg3ZNF7Y6pqrdVYfvfRjLItUsyGlON8oUNx
3o0GuQjYNc4BheOGWcaQoQCXd3pMQgBSRr3hOeXR8m0DIthcwpaX9DG0hpgn0C89
CHIVZAlSIq6vza47EBoP3O+vfysLkgSl6vkrtrN9cqH3iD6bAskCXyg8sCZ/dr9a
5mPqndpcpS8FBXt2nNcQ5pXeIAQrm6fxG2tWx1O78Qs5//HigC7kSEgmczUtp9tv
OX5MKwtSaXpysjCAFxcvaMYRu22bxpcBBDGfqM+rFMiPkglh94ln9KFgRJGMdKuI
CLFIa7/I03dzuUU3DIk1mtJV2Zn1bl5ypTEO+sw7YMF1epdmXpKyYsoQn6SC7+Ky
V4vcP45m+oUTJ+SKRqTf54/VFjYAR4cnJz96IkjlG33iIE9PLHBf/FGjWn78Hvky
pz1/XzZOTGStGUojGNWk9XPCHlDpfzZwtyq45gxcHLj/sSoqhVOn1nsKWju8h+H3
mVu6slAcDQSpx+w4uRIEPW90EyHfzQHn2aiKhAeR9q80cNDz8k/t+gBGB1LNE4ys
wJyAfyJSsqKu1KzCWrDTGtHKClEu+mZtcYfoBglmdWBELrqhTbpIPxUWZ3HQFlav
hbYk2Tx1m3ID6O0HN9/nymnwaEAPNNdULFc+Qw6uWC6TBC5/LKy0AaIZlh+eU7kG
jlrpQiA2OAWaMk5OmKzk8MlvzJ3sTcYPTrAz6yom1+6tdxuWHtmaYaeJM1BBFHIG
+oyOPy90u+2ghqim4LNbxJFBAameNdV1hNo6WJW+vndQ6sXmM4HfIScaZiQ5q7g8
gCcCRzOIYW1QtLtF9lIM+4V6sPEllyfbLqkrcktNFRJNiCjbYfaH+PYmMKhomLv7
K5AKCZbD3jLGFvKS5FzaNox9VSjr2pWWL0miWrFWc3c8mnOICrvVvuCPoVdHr4oq
ekulQgBRD4HTzcJarSyWtJFIQ9VlhtqoRPSF4HsqHmVM0B9sSIoqaC0lvVNPCXop
VK/xvtzQC5UIqK3CSjAZ0+oyr/CJ9O7FbNCg8pkp52usiuem1p80GjT+pvq9/L1R
fHGGZhQXX6F7cN/mOlcUuuBJcEb7fbQcvPp3kf0lHnGpRLQKc5GqCwc19O6f9PFN
QKZHNXUxzBTG54D8hEskX54ov41sfh71idLX9ZZOtUfpO4ElkgFHukvDXN6XlDac
mINB9c/V0EgA/yeYjAwUezMy0EtrX+hLTBsLSDxmDpiNtNAzXzkpDLBDxCJ7VwVi
heqQEqGy1MWENjaBTda6fUfk1o8I0cQyP+eQqU7X24T6MztS94RBmAV6R6VfASOG
MATGFMVjEUELHpLJlD1/GwwV0/crUUijn6YEI3SvNScdwVdLhUWSQ/W8kti7bB2g
U7co731xefSnXXy8Ere81zh3hGQiqwZy6tvEJp1qzzADzEzJKpwjHDlc6YLim5bF
MlBboGk8u5AwAtsfGgck1X76mY18TpDP9suxT3xFBaRx8rPDvTZ5I9e/MrVfr8PE
/KULiz4zRsfzSLYb6NSdEgxGjHGfX6CqPIxZ9LvADHSjQiaGuyCLxEsO0RoBA1aL
fh2VIIc/HsA4qdjMAPAE1nll/leJK6L6jGrkVmP1grhG11YbBIjKa68sL+zX2Ru2
gtjRHScymn7iXGQ/C93HFs8YN5IsFPgXE+Yg3JMyy2ZMhLrlwlz4hGGQ67UMjcdQ
lV7nK/JNuI2PWizZ+kk2QX4kB7Y5JMM0O6cvBCpa2QxtrVmFcwVFy0yf1BcDx4dT
9KcTVmJEZ4qXLWfDrcevhuh33rRqK1f9InISS8QRgAoExzwlx/4I/dsBCRSH3t6w
d/aIK08pUTJuDPRNreB/ZZ+msHJRTVboDCAPIiiJgCveR4HZlJX5CR8Rn+pEuCdZ
0V5fQMzir5dUAFOhT+ef6pk3Nq2u8qfeujtra/4j1Qyl2ZnYWsezHCh2CncY6bya
Zi8oQ84dyqFyuBfNTbPYbhmZPjPflvjhzBoHFmSvH72a7Mc5sNspa6O1niIm3rjr
NcTsOrkqzGVvo8M72hhpaCTqNbp+1w12CoIOrB+lVw3fm6v/X0mdltMub2CMzeZc
xV++EHTHkmcHS/eRvVO0TADUeL9BF9xkMxUfxnadrDcrFY4l7dZvwSCY3w9+i5/4
ZtFuO54PLLxZvm4qXdGIo+2hEEkTA7BoSLR3FNW4+zWKAJIKKuis8cYx00CZ9QjP
lxtlFmpcijbM2sLFpQMmP3dHD5HfsKMVW/ilohIHiAQDTsMsdWaoDybfnJQCEcc5
JWJhONJ9GanFkiHVjeZ1qFUBfU9tJ44OD0FhU++RhMQLrIWr7zkvfB3WHLgnR4SM
xPeTLoEnCEkh7KH7c5nOX1bJrHIBSVQSpi5nCo7m7YDtg0A35XfhGSV+p3ISSD3S
89swfOxw8SQf09kO2hSiMU0/njNlTDPsu39rimmpDfZja4KNwL1aO4I6JT2XrjH+
vL2WYw+GTSQTdrOGigte5YQvZErnTeoLwGXKUCbi4d271/ASejioNPGnJRcYPYAr
r8mrHICy2B5WyEtXxmgZ1PzpgQqSDX5oZ1gKaOEMPKxGIvhCAzmvn4bXtCg/K9Hf
zASO+nRVYyp3sJVpg38Tj0gO079Ig0YLLjz4/miRi7S26FNTrPwDzfb9Ddo6ezej
b3RwDwzdA1TufNKqejM1AZAb3VwsBEqbb2uhDrdcgyXjHHC2UqTObZHnIugwxOjA
PfEgHSeH3o2vHU2vik3tKP6fSZgtLwDjkBl7KoCLKDn0OTmesufoE05o0g9L5sef
BrDTIi596r5rjFTV8DF6ljZnS1X+ooSUaMSDyfVzCRdCH7pPhgtq3fCO666klKgX
7WqTcmUY7lu2p6J4Wnk/bzLGHDJtbM5aK6HEvmceF8nkd9F4aHhEhVVPbAiSOao6
tMCk8rTD9U9uMy0kHBdJZDQSlMj/dQ7yjI6olZOHkWS8rNLQYzLiETkNo1E1xqKe
RImpTeKvaxl5t3oeoGZ0d7Qarp0UJjyUInXPpYX6L2F32s37U7TSX3TtzZfwGqRn
sSrE5lah9pokhuiqBhz7HQFoZfmdDsMTwVsZHllddqGNw/LmCzSMbjKD9dqCnfan
spsy9K/FkIXyAgeNtr5kfWgQwhKLNNYIuWl1wr2PMuhD/SZgrM7qnGO4ynZ0SAEX
WsyEWjdhfGJ1uKfMpo5ww/9wyQq/5RENKsgZcz9zuyG7Oo4QdUBpVJMjaQQMVIc+
70syhQQYbz8HDgqZu6nUqi2lwpP+orY5YNLCXAQdTkdcjkeJIbIkzIeyRWdLBbE0
jUjbyp/x4VGHXcdhH3TvXvc/AKWWE5RSfb0PtuaPCVRIRgYNpi9MKCdd4Y6rUDHQ
ai5tNnUdfhr+gRb3AkfXuUT3Llao8ncWSPQTiZrNdjZcATgxWcIsRI48n1EGUnjV
QSfno1JkgOTFPqTaywNLhTetHQepUsdPzMvnGWFzM+9otvvA28mdPh3Q+ClfVoP7
YKPwa6z6/22FR1AWPUTi45HAvuxuEGPayfdGCGz7drIfvc6S45M3/mHCqXh1Ovat
5Hz7ZYlEDyO3jHwCHgtjyFmwroLfy1F9us75m83j34jqn7T2E8TwNSbRCIwZBMzG
nMGCSAz/j4BQyibC8lqhCCUQSHsEx3w9WS5rBMwbPsz+obfVNG/x5RkU430Qa1e2
xh8t+EifmavRyBTmqnWGlpBNmv0AxGIFDdKESFjctZB/+pjjvM113cjGgGyWtab2
Q3IhaTOhtmWz0RtIage/185OuLhxdm0UCxxkzXbK5FtEUa2Owr/NAZiQEJ6lEVLU
pUK+8jNbcuiA0b/on8AC3TDP7X3lQwgZmQk7O6LMpPbIAQVh1ke4/cP4aEUilkbE
Ib0iTHeKqS6BjMtJ1c9pOvptP4Nu7LDMfCmuNDBLykn/B+5an/e6j98fCAHyW53w
wkxIYTSWUNnJUHa2/eskTtlv0P0oqjdnUw5nSzicfg/crRlAMF2XywfAb7CPit+F
ilvX6A5x8hHJfmFv0ONPPKX6Y7CBupHEa54g1LXZShGWnA/2DmfwUQU+KEhmtujG
7SEyKDvhJDYAQJYslXHQCY5Fot3YNjwGojIKDx1rXvexK+txOhK0E08BLeHWxCjL
1ce4YqH8vXFhvD/bYGOrN0L+XgolIH41mxpsnnAPDoxpqbr05XejmyKgsk8yaTK8
1QtWkkHAbTJdItNlqh54gjGtEYpVDtGAj+/G/K+mH2B82HvpYN7R/+7X1tcFOd0B
gNIEq+oYRoWUjDhRS4lc5BWE/fx6YKjgbIVDx6ns4Joy562PiG9E2aCm+4oQJDYV
SuJkNBN8RoXRDN8baM6JIpFsa2vBeYzkAGYva+mrs4ez6WSKCwi/3Glla4I7DOsp
Xqh8vohO1QzyiN/s34QUd8gUUpGVM7dSCYEx7sl5njuF3NblrsaSkoDNpx47w6W2
O8JnO45P4uvU6AKxqtZcfmh3i/jH3xD1be7Z4vc3GTXorEmmn+/qUMzJLM2bJIIq
MDH992GHAZEr9DI7ASV61Ymry63GP6FLs2ykd5e2Jop2p0nw6S4ePjQbt1GJO29p
LqbleXbTqy6/trj/XAIkktVtKfGbubl0lXqOi1GoYRxdSUwS+wGkrxFl7/5bw9nF
yp7GKGVE4hGWXUZWYXiRwfFvecNFf8BYPTJSyjEJ0IXTF8+sKmmIlYi/vBJwYneP
SFY+z3ABaJoPPTfBXo2o6ZvRhjVFuazVTBwXgOEiEQVCmk1WP/gggAe0eMBBhEnT
bgUgcy6Lta3Im7cqHpVYMgLanYuM7d3XU6MY+SNG60HQU4XPdeIyTyn4xk+mgNK0
f43dbbluHkb1R+UReDeRBmJxpahydVwAqnHd62RchZU5xRDwwR+vFJ5kjd/yCqtR
8YJ+uZwmDqbvZJDvFOZLUu6sspTKIzSXvlP2Spm2oQiqwH8rNWR7ntYSnNmCNT6W
pzMI5yy4D47SwNaLTqyjAMhntffezgvaiWeRym1PS2z9GiotYxKN1PrUja1jy7s1
vKMVw5H5i9OBleZDPLnEP9ogkv1SMJLpzeoJqTrhVKeptVGPjXIQTcYa42LaHLbY
i/7ZBdkC6YVWlVJPc2sJ+Esl1tinbC+mu3xV1RzEZ6WaCiUwP5tn7/v8ernndRgc
aQ4n69pk9O/33T4b0d1sTqNseGmM95Vd14YDyTExaIzZyMg7DpyKnA8+Nq0V2wq1
DRtRurS4AhCGLWZdRZn4rFwD1d5d09jMHXY5GbAHiSWTAkpIEJa5qDheIti9V2Ch
clC7FQ70A9f8AuXQw9U9YIoDD8jshss4hjGrvbh4fMPfSthaqnUOF6ysbZUSVH1f
Bas02Urbk7kz+AQfjL/fHrNGfu3JX+tEctKPuSSvLVdHaZiWqKvBZfYHG5OPvCdg
L+4K2Rcgvq38BoM1Vo5071FbkUWGUrkoTzEcGDc4t5QKWe5Duv09cHtY+Ur0j8u/
wMiNCm1B26HkEYecF+BWUSN+vqesFzhV5evidnNCB3BFrerGowcEb1hpqUM7WAlO
J+AaL3p5LZuyKfeuWpekjhaN0WsRDtbm6wmLsJAylgCy8bAOS0gIjns/Hdv31XeC
SZoBbtRqvMpy7x3j5NrMrMWipj8W3sK8hpWkoS1F0o7KW17xDyiowvvJGsIsOWGI
MFkZVpx7TBl/HZUY9+IvpqXjK/cMyQS9XtaiwBm9ZggQmiCeAWpvIgq9K3d9Ha9g
tAXM8KmftK/GmUASfRR6XmO50NkFf4os3cbuJABkyNxBQl9MoihtIizpB774Y7RB
pYekMnOPNPJ3x4q1m+Fgw5gveqNKF+l9XT/969zztCKtRxXpTz9NUoiYsd00qPl3
VangNZE0Um5zbSn+pY6/WsUnLdDApxSS/guTdSEfjRC9oPwRxx/965agAiSwEwSD
4jiJurrlYFLGRn41wGV8kFMjTKRPzEl6US/xILYVm2x/QKvzS/KHazgc7Mdmwtph
+HBVvSI8Vhgk4XvOwx4rnjIHKl8+w63TDfB4n9SCvZtBqtuLw9eh028/XEKRIYyE
JCTsIyOvGcaz6nkfD2hG+awnLxmF78r3I/qqTOEdlSs450Vk/n1Uu+15y1ScTRpE
t+B5wBUs747HK9I8fiRaT1c/io9HVkWicUDsz2mayEQp1QOjAWCH3b/8khDmtASi
BiS+COMF97HBFUstni7pvrBOmNHpP7liCN/XsL3TIR/ROhxQQhBJV6Z0sjw+MCKR
Ng2wEIUfJgYZ+iFfM9HOnillbDWV1lSnMXh8S6I1NlGySJknMBG48n5hbWWdKMYt
Sw2SkyhQ3r5Od+VOv+IfOHe9r1HOR9I3t2J67C/BFHhbqFAuv30Jxtm7Gq6GaYgW
ZCnq54oFdT/tJ9FKUCLT7GnSey31xcK9PtWqOWafNHeOLNG7+9vCqqkGCtb65yjL
+1OuB4Ws3sdH1JuYAN6vaCIn58J88XqN61yHtXX0/624DJ4B6U2+oho8BWvBaj21
pecB2ffvkRhEYNudkM2mUmEj0Mt7LbRHi/aFQHdOzBW/c+ySGXb4rrGIhcfFV+Fs
/ek+b3NNyFBHoKTfVjt7kmWXXZUA3o79n3WsvrME3QOCKZTPmEsfsp875UN49eKp
gR92B/2z+k/mzrcEMAeSrtIetRsl7qHxMDlmSyB35Omf7R7z3cF/Ubmrk/vdy6HX
bA4hThPqJwkmTGlgDnQy6YJgQta4TM+B+lGOQiH2M+li+eoPZnkG9sBRW3bAGRGK
7f8LBpNvU+W5a1YUiSxgVnKle7NpUZuTMT2ouxB3UPqMbit7aMQ1n4nvjh3oiJv4
XYd7BGB4lMJ6Pc+7W653iWB9MKRhSnFHl5J9wNGTAxitDAnNNyYnaEhCpzfDF/VK
hPeNIF911CbnXCG19VdXmBe8qGW1CSPTUCS7RYUR+fVYJk9rhw7Gb3ghLT3pFTc7
KMgFIFKE2GYgD5aN4D4gMPpH/+I/gxJaiz8HgDg77alH0TX3Gc//luVIlRVet7o5
R6zz/tWZOUu1zJJSgY791dBbdugD6gAnuwUJH70OOFw4mRQiy3QIzsb26r2X7bmb
OqDGei7uCLBvGO9/hb1vOFV6tjlkQwH9IzkkwqcJer6YmLdwAMiP6HNXt/O/MHuP
IcbpLfEn5HywKjLaYg8XdpDnPflUmBR00A7YTPJCc/NmUBcAMvhysujlCg09mkee
rHmgpu4A2XnOAhIg/O8SWQ4eOp0M9wgv4gkw2W4LFvUVneq/nVU9sl/1RhgmseJq
43neOC4NdAItrvbaHeHlo640PyYUdP2phNEQZe4B2vuzKsG3K+fgjI1ph2na34Wk
WTVaIqUifrCEPLGeNTb9+i12BKv5dok6sw+9+SKfjlmPx3EhyYBVMM4LAU7cUf0B
Dyh2rTtEP7k7RxXvd9vYier24EiqybHJuuc5gEwz2KcuGpjBpgH9AsVW+3e8SpZM
9/VO9aSwq1vp/RsOYI3FQjSBrfor8iG/k8g2wVOAD2DY69YMNmgs5R5MjuiC8QMF
Hv52/wTDAxTUwkZYTNz7/AFySmQt4q7c4Hgz2G60OIFGoNkhj6C3D+4iRDxVq0ce
EqCAVU7q8DPhpH6oF1gVwTSK5Jh9AnGToJydprALFmikeaHjix18Nuim1jhRt678
XeAVdR5NV8LUlW2pZEmmbReoOx/83gVJKjKz0c/HhM6y8VSdgL/8IgyacOlUt0cw
dntPnpUG6QElw1RSrB5yzr5BS2OtQ4MwvA+D+KJOALDTs9w6vDsuKdUEj64gr/o7
W/ZX5ynCOFoj4nBy8Ig0GcP6sQS5BrQBaBVkJQl2CnlqMPf90ZbfGXuGgBp6oQmi
uaX/Gn3f+PREMuDX/96xSq2ThILFLgwRoF8iLY/tYpY+kkCHOWcc02hxPkjfPEv0
hHwfGtN0qY2/Si1C1XbvpIflDAdSFe6jBqsM1EburV8MZoAX0bF8Vkl7pswbXpVf
AlquDO4wI/KtmYD/WJLT2QklFGoi/T0vGs2/6Nrc1w6o2yuyj/fcQDx72+RyRxoZ
zdLqQch2TYBkIN/EvrDRGFj106Q3Ho0VX67vEopyCh6lVZ2S5hAQDjzCSA5aMTvH
sKuxsa8M91PL8a9U2cs2cyKEd+I18RfyIOQmRfCL8Z5yEoouKc3tTezbM0iocCyU
iUU5+mxoK/579vAXHP32v/vAk0kVb51CiM18SAdd2l6153c7m5m6QwyIx7UDPFjy
rRTtP2UzkXvX5o2tX4qI1f4aVFjKprTWOjyY75ZrE9K4YqdqeOWbaBaoyzWmwMNA
P6binxbEZ+Qrm0lWRJ1dSQ0frtTqLkRi56ROIXkamtDHeJCEPzyOrTSwen43x5bf
uNFs523tlKIZRoC4t5v+5qjn1vTrLN6aXCA2TKJRCyyp94/7Ka+VjhOgjC+RlJVJ
E+ANv1DBfyUUPjMba1TG1kDUx+mrQ2j5Pa8Nm4/BFq/fKPUo2ek1JokjZ8R++uAM
v19SFlV2AkMq/YITOS9xXN2doaHCL0DbbonPfOzT/fp4u4U8f3KsD1T1oSA9vvMS
4QtE5RAG4mBxBInzpV3GsoRHOBHK8csLL8dFnCCaqiKSHE123kb3Y6fIanoAzdiY
sKVGb19ZJSc38t23rLDI6wVPZXPG4vAglWotCGWwJxDVEB8ITqIB/endK5HqUyU5
oP8/KIlt4Ipfe5jaI/8/J53BFAkmruUjAsZAF7+tq6/Gm1U/MT8bbOCX9bAHzDiC
J76uNIpE7iZEseZtwr6DlTR9IxtxrcjhFyndciTYs7YynguxdTk2hvz1VudzV0vg
E+TLd00YbiXLc2cQi7cdWeDC7fD+xGe3kfXf+OAZDArf2DrVugMFvmBFwzhK7aWQ
qrS1vCU5ENfHSmd7X/OMSLkfvpilCx9wwZZxzePfEN0EZGWAOuJCbbwYffr9MY8z
N/MYeLSbQIAhFgeJt+ZWNPuO+GzI1ky6EvPrCcZWPzhE3ZCyhGwSg1lKBXtCxmaG
SzwZYl8s6561q9jVZ9OHlfrhNSquIFy/Wtc7NZuljtl4T4qHGn8Kv/HhNzg99hsm
6dHyZNqD7IRZaA8HAucC8yvpZseYt1XywfoF7BxAReAFSb75FDOK0Pro4TKYYVd3
fKHr0peMLwyc0FDoXvhrV33ySy4WKVrNR4LCoJ4IQPWQVJQqM7bwhPTWZKFTj7Tp
Sr+jbEL4/9XmPHYZkO03/eeOfW2evyTjonM51OxlGMkB8BfVMyMXcxCFs9saH0tQ
AxBbdf1z2+mWTv52MfVyKbJHNQd/e44t7sMFDNNskhSoa2tOPSy6ai0wYoIQnv5O
8XTJOKhZU6nsuZ2gOEWwzJd6GP+a/krq5IvvvxSAJGWDGNf835wsI8CmGdDoJ7DG
5rgl9DS8o9qP0kLdJn/PbM8+cDg4NolRCe5UDHobd48O05nB0Y+cYyLLg9+wEYnx
thfAT3H+OL3ZSMQX+ct9fg3x51VVWbEOyEtwVZonGhLhcvd90ufZD6HBqM5C1GgQ
aGAvt+eNijheoog55pCCxZlyiVKrnpjf7Y5+j4+BUvKlpynibN8aozquHuk4r14t
Oi1nfFnOqMKYr4MBcAZF9VeaM599PKgdMIY2IwX8bbVhdUZSfggCdmSQqtG7vEKV
jMnT0gnFuSS2K/v7EZSIMtOhDYKaLk/9NWEDPwtWLdZFWoq4+mY4gyiBT3paIwl0
dRXwoDtOUDEl4QMoT+lXAwG0O0/eUB14EmlqNnFChNzkXuviH6WHkxk8G/GTzd9w
pJWoyXQAS3PedcpZTh43ZhtJ3dGzGLQu/iCpU4Gr+1RkPVjygcrAbha94r1U2ulb
bu4WkFv87wQcP9BjqvBnO8E9TNKZvQvoUNv6a0XZ3MVbRCSzlYGkeFaYqCUWRpmg
dlwI651xGae/5J13LLU31bdF8h1WKJSQ02Yf12AyWHL7wUNQH5lQ2stWIYr8Dnap
WrqF9H8JLSSraQUfTZKJHJ51P2FY13UWuD/NI9VvO153wBgvolGnNN60o4LXJrJK
XHETYViDGP9rrTG/6GnGlOtULcS09oajBy3mj+stvJbjyFbz9hdCq2TtFcfL9uAG
mVHup/Tk7tUuhA+7PHirL2I3mt7L4iuQQD6q/6IqJ3ZAc1HaD0fGoz6ZPlHqZ+F1
LpbWXvGRqPsdX2n0ibFsPNAsxcHFdO+5lKtFOG9xohgpfHe5sinv8qullXL5T1EX
hwP2nG83mc9Go4FRcE8tf0gyK++ACdzYm14a00JLlmWYXaCHQBigT0d8Pm8u+u1k
1Nm+a4W0oUuyLBq5/yigPBJCc2NH3HtKuw+UJc0GyHodg9HUhNVdijc/ISN2cG8k
VdG+wDQuuPyoUHCvIRFTwWNXnWLuAZc12Wvhp/g4SsR3fv5ZPvyewj9ltoI93FlK
GO6mip52MsyFQ3wNl4L0FAAah0LwTsx15U3oWObnfikV57h0g5RIbeCZ1izDh7LJ
BkDVZOK0iSP+/SY6lff3+b1/ER5lLJq12YE7Ww/VFgW59W7YTEoTwdm0AnGzai2h
EOxgsfIxXpRrajr6SBvI6heoUO6caRL16gIQ4nXAF57dEHG5TW6aWg7eaXcuhzTY
HUVEC3ldwZoqFktsFRvdcyF3et0reFMENEZtl7zAbCwumAvnje8ka2kQFy+T3x27
vuRBP0oyFj0SF39Rbnw3zEbwVEvde8Nek/SK4FQMTMd2osDMyKm85zXmSUDuybKb
ildHimgLvmkN9liE5V0VEKXVrFsU6a965s6hJCQ8o654rEwCHzTSAieiTDYnX1fg
DBj6J3qEXF2o545JJIvOZQSiCneKAtxZMRb7nmsO7rFKAkc+bi4dI4qxqaldR/gv
19tlnhqoY4vC+hTeQphkSggsb0V2XbuNvfeJSId2ejMHsiKLl8D00mlL8/a+HQOc
23Kzd9kc54mG64tn99FVV25d7VS5Bwb+dm61G8KFf4clNXHVIAAJtxlnb7Uf6uYM
gRM6ZTu8KK5OLe93d6g81DbqYbx59u59lG83ZBKzqoQmKyfJHmsOyVCPaP9oNi3M
ercJduQzyl/vP7vUcN55+I4Okexdz8DeRe0m2a1XW3sT2RkoL9d8ZJWxDubMLEI5
15OvOOCu9VRO+2NPQ3wHV/ICpC4TovNx/tsKxGZCXfcPCAtafyn/mE3Jn9MSOTrm
i6XZV5IOC0iPo/Bw/LfVy1/zYnfVTR5oxjGpwQS5Hq6Tgm6ETEmBPFX2ZK4iq7dG
AjfRbal6kyR34MUqZl3sOYwTRVFiF1vmY+GPxUVfWrKyZ2KfsbYGBiM2VNfyUqC/
IjnZmlw63DIlHAyNcyRc52WhKCB0d1tU+m3PHVjNH3vs93l8dWkunFjbHmugIJa1
1//Wpewz5uqnYmYucEC15LOwFgFHRuSRhip4lN0DnP5W0rP5ROL/wU7PmRNITi5I
43NeVl0mC0bxusAaWWQROC1RtTPWZz2dF8FtGfIKwGelakQke/Az4+rVxUl9YFCm
r5WqliprTcOp8FYsqTIaj+//UDh7hHHGx1vusHGoeSg3VKjg7aRvCb2rdX0OmWRZ
SICkIYRmzAgO8pb/kx5dxAn9TL3BBNVCdLwtiR5jTrEi8AcPOh+8mlEm4OzLkqI/
pvsRjonjJgUbOCsL+dFH80Rpxvzho7I+/3prWzvvte2Gd5YJmO1h0b22FFyusiW8
3fFG69fkz98T0xcx59U5s1fJjYQQbDcta0PskwqrDcWjl99GH1t5aLmPGYlPe1yj
tIEgE3z3+/EyGu+9C7AdlSbMg4KvodwG4nBsAI36LO8cu0OSs/aCTphCuwDckMsC
liaI57NZ+rRHN1PFuOep4t+3IMiWYz9qHVVFROnjPM/WwARqRX5I2S+JDlXaKDbA
7fLhDMiQAECzxLsOT9/jh3gSdjzjzYQOQAsni/4I3yem6wEy832JYcu9ANWVDlyR
g7YibSgUykJWIZOAtS5DZfYmt6KatSScog1fVkDpatJaqFQdOYDagp2ZAblb47zV
IHtBNTzZRz46aReQzjxQuTkBAf/PKeTjFVc1Q1pp9/78jJiFg8r+M+WTtGTfDF7f
wQ6QpR47fLj2CUxIx1Yz3wd9RXlHlo/hxHEFYiqzpUT0yvsfLAkvdE3u7fZYQbud
+yvgAD+KHLIBH0HJwt3GBZxjTYOWiruTIw6CIbrO7VeZQJZgAHqsmGopBiAjTq/B
TutWECAqBwLM/wPAxLrdiqQfhh66wECtwnbI9QOOoMaXgWaR1MWE7TyeWhSQLKx6
uMnfOfLXaRPLRx0/KxwUGyu5/334AjnV8LDJquIRE4hPsV/bH+xrL/+mLh5mcSYO
edTQ22usmVANZblfxLYcoFbT7zrg7kmPXsaMn6J8pNPzss6mAItb4Or6/W/BPgm/
3MHmLIR7TahfMVRz1gKrPhHHnkLIDxwBPcmhMHLnTSuvtuEfeW7/cUDt2VnChtu5
60US6Q1JWzgv8R/47aO/snjJZTfYwdURnGNV+FEedDzEtRkLTfzr5fh6A9bh26cR
g56Z56pbgL2k+x4XP3hyJh5pqbgYI5cByXPr6tvBZAhw2CivpIxS3xzjq71fqWIK
UcF29+0s8xn6JkThMKb23CioXglYcBm7fVuuWbgzbfQTP/RvII6+TiU0yg87oezd
M7r2eRWd0UxsJsgmhQy+El+Az7yeCHMPkhiAYCu2N7pKyt76SsKsVvGLAkXs+kem
4zqzPsBIj6XGAkTSTlI2gBz+Hh42tLqOZr2rJ2bfCyNmU+1R8TmwvJt+i+lAGUtU
6uj/ceS2gAlP7WjnIOfSlSsb/lMg8IrnPJj+TZ286p4+RHTuO1CK3wxvTkNF9+t/
E/pFgBR9vMO06vx6RZwQ3HcKqdNcXbLqpz27QzmqkU/dJifQZgpJSlYu8HdPEV77
e/iOMx7fOZTQCKrG6VMIMmf34nZK/vdKOXpdUB6pA5P99xmCBKEeZU1HoAI4ijSs
e0Xxq1VsPnm4rVX2Kl7Q4zT8M7L58/uPNxioigUNfnVppkyAVyJxG+6L0zPJQ1ov
q+pwREJDG5W+eF3sxXtCscYlmulTXpEdGkeIssjqj6yqHcR5Qd0utnxWuhqxsyDx
0cmidqu6Z+q9ZW0SuEgVIzxo5AxbgiuDOADeELGoeAVnsY0UJiB5yRigqcd5WYwx
xXPWHBoMwRan1vC25IHAy2q7sNGHpj9U64Wp8/9TvO9rtL79Dm/p/lwok6RwHWtc
8KPP0qlOIyqMAcwrxFjXc7u/CJSlMDjlz2s+Hlz89pT2mcYWG2ModV3IyHu9Xg2f
uGjfEa0oriNy+rFkr91r8pXDSGgckosGlhAxx4vncciuQkI+3P+wniyI6Oft/hiq
+Dgv0a5CEU7Rt9bw/bOrMi1YNstkuVCpNU65ANMDs2+Z7FfhKGOCR9RkWJjEQKJg
HUP/MGX1cEqpQe0BWRVKKugTPcrcuBSKUnH47Q5ERvQSIrtV/LEZDVYNqFCEc/BR
pYUVxKf6SYdbsU9QbzkNiA1J4i6088mX3xcV+3ty1gU3E7PvLFrji1L5BSBbD/Ki
pD8NMamVW1rbMfUHuy721UA4VSBchrNdzBEPzE6NqwggJkLL/2dHcj1t+NjorUb3
SzGEy26oZceGwN+LTzoaAFtj4nnnmBAVvXzOl3RN1X/uxaVYsHMvPnKfSJrMUNaH
3dYZhrZ4x4CWEh+GCPJYGiTee+zpxvbjZ7fxUrJcr1r7HvojWr03/qA08CihyIr9
JuLaPVL14A/3ze/iTQIhaj5eCNJ2otWqdAuM+HSjDqW30KG5ijQMcr31F6GWKjHP
3OB3fBFymf2a2CIAJ4acfujwQv4ykwVYGSdKkxeAhPlh12efv28m1XMphBC0tCIx
nUkFu8MciJA7RFytrX8FrfM5BHyCwSzcW8KowqFoq3pTZzbsZsg+ni1yNmw+xREm
OByDmXSycyy21NXnmILGzFKZ+F7DzD1GMWNqGOPlMX4Bn/Pu3xPRjnBLO7H0Gu91
NI8W1p/Lmrxvsr1VB7qOyr9qosQ0EIim8OEL24nN2TgzTyjLIrHEnMmTudyK33NE
UCd8/u+gqoufm67hcnSUaiZzmdv8hC2ddgtQfU5NxWN5T5Hta+ZmQx8PZVDt1Hbk
Dl/DmC2mKe5OBXzkjI1T0SaIGTmO8ysDvBxSsUD+gIkOa2kNRa7PWTNYL08HdjTm
hXQbSDFOyV7N8XjG0YtABSoiiYXBfxAkPhdAqa0FNTTm+P0rn+nUBTMwWO44AflL
Z1/+ZJdiYZbYokyDkdu6K+oi/pRRSLeh4Lp9/qPdUJzHibA3LD3zo9OpqWzK38SN
kI6AKR+1DM0s8AlFUHMenfqobWAK6XxXBHpNf+1Xx4pRB8Szcla16Z4z/pmz7DFa
b6VSBoNcHjoP7ZKz2Spc781fMrd2wx0G4835Fds8MVbBsR1+ILJd3YIl4b5sjRk2
mbQlm23I9bcHQpE2zzwYZIbrNV6QiLWwdPSpjkJk8up+2ukiPeFMAlhvq+tylAOS
iHqKRVeU/WCVXw3uU5YxQ1xBFLK9UwKF+jFqoolNSp84/tAo1+iyidpO/wQru0HK
HxGweijW3wTw7+mtKP4444FU3SzqPUDCTCgtwN6RYBqVQ+heuW2Kef9MAvXWkmIA
1a0Kc4bQdlL1uWjwBL9oFYOZlKmFsHwS+boM09K/Wyfr8upily97JkdT+EJ82foV
EwIYtr/Y7OA3Sk6/3ANEv/WjxHeyTghYKcUDPqgrbETTJzI/I9OVb8Hz4c+1z9lW
c7bWZy4+zFmnjy/I/kbei8Mt2J6u4gDU6vfhD1djwJAh+3qtx1MzmASdSmiujZ/e
AFJAzWKEWKhnVx5L2D971oc5xBauzKzF1KAURerhbImR7w2yOUqXYrOZGn56xusa
fPkn2aNeQkVvqU3PE68+ECsFLRLDQbhw4A37Xj9SbFUw6XxWvzgG9UTQnphW9Gmb
2rZlfW8n9fauWNlZpCTOnVZ2c4O6z8KvRV8svDLfuOp9z4SH+W2XRxp6bF14llAG
6tzufMJHpL167rdMAr1+MuLXSEYN/02xXySO7wLqD49gsZno6TNhGNfAgg6ITiOK
7+qM5ZWsrIVkdFgri8z/Hf4G1XnQVON7SRgp0CNTMIsNCA8QJbpdCcGR4DHs3vDp
TS5pz2Lrcw06QkjKwsmVUs0msPMwYp0gs9SJxC2HAVvQbfPYkIgpff7FjJc2IBtn
kt97HMSRJd0ChvMYzYWVMxfWZvfU610eoVj95vue1GdSo3XqKkMgG7hgE5I7Uw5C
94kx6Xp85SXJXmh4ui1KbY6hHj21gD1YosGreDjmACzChDikp3tC2W04W/OJCx1P
lifFU0QMEVUc6vM39bzQIvoWGabO9gcdkS2+S127UoRMVtsZb+EPWRcdn3OsGcjZ
ROlpK41VVvTy/QpNNpZ3c0u0WxqqFc3hTY5QHo3qh1cefuRuthvHpvwLPSN2S14T
RRnHcmoNCpCkg9pvyJmCdp/ZKRvXyq5uk9rtFZwB2C6pT5kilzGYlEZqfNgdrG7R
dzDkLZYaXlJww9S+5M/Pbk2zDmr80SySeX1rqgNA4h6TFUfECRtlxlUAdZ41Pibn
bOOfdk8I8jLJTAzG28dC8TFdWjecjrB1AMbRXzgT1hPnrV0NXiVv2m0NbeEG/UvD
GZiu+sHlItjarSI4o1V3/jbPWvxjR5lIVBdvj2qe0zDRo844xgXM1W8yDYCgunO5
nbcpTlJo8WdwDiukjBxa44s6MwSL1lKACEd6Me32HyMTOzyYw01FonLgokh6aobM
T2U9v6moqT21x0Gu5IZ7KHi5Io67ygat1HupK+T5zCgG1QwVG+mE4LM/mvkpaOFA
Iz+68XxE8fcdbRTavZPCTUSKehucBTPIEv7gjzVXIorvkl8DDkWOJ3I5VkMSjwYR
YR3XjU9Hs8tXmI2oJqhjFcFLCSo2NFunAAP9qQAp/d5lUFsozcsnUa2wFI2qVIw5
ouVkJecDw7VpIqzp8BwQEClgCflX9JHRg/ftmEhKfsJ4K949MqYo7QiEw7kP0Pu8
iXrLa/4yGnOavE5CZ96Q7YNZFFEqx2geLpBR2naiwBB2TT89Ozli4IUy4kDRSoTT
jS1+exGyHNyXZiyVF4sayCPPP3rL1peXyts6yaB1t8rqEgAJF4pnwGIdcFv0ekGJ
TM1HufYrLHNUFzye95FALfHMXYqg6qVGyJP2FmaJiam85706R0h7n47kLUiUU+1/
uigwyNND5qSvraS+o8XzPPXSw0GXwW9h6aAi2g2wNawMk+Spe1Pl4huos9opxcd3
vw7G8mvkr39oLVi+srjiO4KwxEWU5NbD+VSE9LlG2ex+270M/rOwq2FSNBrM3fr2
RggIhUw7a6uudktsEde/jCI8Fce3CzquEnRfbXN8vbFUPoWn0efQDMG3ca2VAdRs
BFxM/YEOU9Ka7WQxWSA6TG3J8v5qzvjEhjp8QvNWezMPQ+zqyuNaa1Jca5oeXNWb
M6v4TQ0jDV87hf9GqDwGP+VbCDj/jcE6XA9KTUQl490evc0mtBzvZpiCuQO7gf6+
F0b3lXVx98vKsAja29jXrDM0EfAHWgKVIuUJWY4KXIlGoR15KwhVjiCZ+Ucwdedi
qhJD3dbfn27gR7DEGvR1vebZA68ovAVpm8p3PjnIbghX6Hdjp+CmhOPmzz9aJg01
7VBOEPIWPRRKirWU6SzzsOfHfq+mSRToNZpHfvZ4nLY6UBXQnAgUcWioI+fwlq/4
F9dXoQcnUd2YvPtiiBgmN0swWhcGMOMG0u/oiSbf2pWcz02KUBYlJ+xL/7BHFqnz
NpNWtHjY0yBWK4xJtPXqFRnPOdB5uxRbUCRRIpW8MCmunZt0eh+XbEoDOdjzaXqP
iZ7vE/92b/Gqp/WejFCTSJmdQSujBrLdANou3C432eOhqNsCLS6dXios/jCzOOUd
C7Dy9KF8Y3ms/SOuHTRL5U0BLyZUPZSJgtg+exwd2cujNEwiv+XQvNolSpXm5vxc
mkPB/aFA4GPpry4L5/wbpbi9Scj5rJmkRE3uZE/bQbmWlyvxAJnP/jZ9i1eWaRNo
uVxY7vRc6QCM2QYYJX/sVKj46FvvwMFjwozb7lSmkVIu2+inDoIkk4PSYmSUwqsb
oPNRlyakaXz63nXBUg40QFlBpyT5gkndprhudxXUyv6AXklV9sG/BDd349+Xf4Ma
OhsguaqLP/qcGih5K/lq5QgDhFvHopk/hMDeHTkgG0GiCqmwrS/Tqldo94C0POS8
JQ+LSqBzFZck4JFPPrNWn20cjWYTHg+v36TR/zwk4MEOkBGddViRLtCJ+n/2Kk8c
MREOZN1XqAOTf2KwxPOptG7Vk7rHsII+VCCp4uSJ18bQdB/GsQyosaZvzW4a0K65
zCRODOeTZPfU0/50B6ZxZ5F+ewvnJ7O16PAD3i8Tbrv2pGY8el2d+K3/VsqrqYt1
1urB4QASfpT+JTR8xTn2Lp1PhZOW0NhLq03HBfplH+HjwnFJ5zAR+wc/4oP6dybD
3X40CmPTBQ3J2yOOStFJMMZ4pScNLnbaezvAsftPHeYZLxvSQYqPNO7mhb8hiUy2
Rnl4X2qno2DpASPoXwLQyz4oqvZ68JWoWcHSLlCP+tnVHTP4qB4GUN9Pr+TLPKdv
PrpZSHFLzS3ekvpsVdY7hLUUBWSvhJ99nS8p/VQGeXQycbtjUkT4uYTWmo5tA0v5
bdT2T0JrU3tQ4L7zRS0n306kIbBW1SWeFoNanRwWnoiobWtF4NzuTPJDZVkMtBXb
+6CyYE9npla5ue9sVqt2cmo2TgXL4OALaUl1Huh8vhViKXZQgnvVmP0/2XUiATcC
HSg+qVh1Ko5GEj/bCotJYSe1+KmoMm7CLYnTtwh9RN4xVvg2lLgFW6wOxH08gPR8
0BEb3Qp3v1wHQzlR9JSshpReFHRWekRR4Kas7+CWBwyc8hxmPjm/M1k0KHmUqTb5
gm2bD1GcUe+pPwwSiXwRX4KBHxyy5RPQl0Pmpm4UyCs6Er+XDfEW3N0KqItHf03Y
0DPZLmHOGbvnwhPW6BPdVdXbN2CzT4JvoADLBl/9iYTW/E+ZBFDTBkB4Q2OPuKiD
8wF5NENZaJNr5Cch7Lc9aTLzVV7qHa8PAkQ94XEJLRNlqVqdVnTKl/J8/5xKZhgB
C4jKgC9VmRmp9H59FjDfe1TtP5a0jsZvLCZ7BTqz8tECi0gqQ3CZG8Yqabc+fvDM
+HNqKP7uoVHH+Sbpch6dhoQJE9A+UrlT0D8qbC7w2NgLIYKkjeJT84tLterE9HyL
fGIz/R1n8wtOD7aoz1mi0IpQ7ZARLhReAC96Vr2+VZddqNPzYTLj243PAIHiJfH7
l9sYPCcn1C2lvGwLRL0+NpMbYx0CCxbA9EdMm+kBTeVa+bhwpSPGoR4AGa4XmSNP
uPdMBV8YEO9AUqD5ZfJ2B7tSKoz+9g8TB6iDhar0t7RXAz339GgpZCdgFdV9L0hJ
BzESswoSZ1EsQtA3mZ6pa6Sth4lQs00QidONfaMeGzFhd5bP0mfCiCFrBV6GnNFC
BrWujmkzzKgK0fdjTkAXe8wSP56jPgaa/KmeW0QLijoNYjTKY7OS8TYyQ7aILdcW
rp0ehC0W6YL8WEGFB6eDmxq89hGpGzFYu0cjVrrU5kua0z4h+/nxq9mty4pGkIrt
IU74xOnwNJzxkolHAbzwYjsSaUtYFvp4Fet2NJ7Q96/3ATHlhiaa1cHDn67uGNZ3
VjQDF4aPJR6j4BXHTGh1aeNJr03Imr+6gEL0iON/dY8++vKyNwqzoPINemsNPj/z
lRm+956pBgoIcUBxehrIss9nX0Fjm56h7/2YoqM7b9j5fSg4rMkRXMi6pe9/x1zJ
g9BpUqjhcdU0iCy/x2ulV0ZS1alhuyxWpVdFFjErwqcoDPKR2DeKsfgY/oomERKa
/YotsfnK/MYWDbrGYtn8dYjdHL9UHrWukiuT3kiXPC9hYwweepP81y1pxrGkO9HY
9iHtn4XQW9DM12K8eluu+F3NN+kKdfau/tYiUBNEQQCXFnBS2hErSnSsuSAD+AZB
ybJ11EpPEtNEBa4VEIDT6iyAgb2+MKcHx/+tS1njt25vE6IZV/6YsCK+v8t0xwcW
xtRVKtMKpW/zx+Xd96S78PjhT8uSJSl5qPNhgbwDNw04z6l5DyBlXFszdIpr6pix
XnOrzWqLX8ZPspXRIaQZ3zYT5OtEf1OEdP/WBTTHG/SrybEJOH9awu8OF29od/pu
heiO1MRCfAhcRLZA75g8rREM40yj4RT4GPFDRjFbi543/yUHJgR51/90DQEKPlcU
FbT40vKPtq/dO+aJq3j0bdlIfXhd/gDrCOq2HETsjH24tIt85DS3Gc63aIJAEt/h
PakZ3ozkTGfeJrvu/OTyceqpvBynVRFqbrNgsgN+xXpmdLtODrSQCbD3K5x3KemB
KnJaL8YHZZ/OyPt5dcoecsLxiiJ/kPXnYmEpV8lmPY08sWRRITqk2Z+WizcpvHr/
Jv4MOitYomuphd6+qaAmkNxBcFeA1q8ufPZfgFgvxhsNEkbVX9dJ9BABPDBeXKev
AGuinFthGmMFFl+9Bw0Fi2q3FBIYbYN+mdWn4MzBhN1HI4CRvRLOaZIAfrUvlqcu
+OYA/jXw0pHd4M2oXZqBLgaQu2tx2Vqchh+AAHLDT/j5KaRq2y6OwNtqdiJgxrMY
61fOMB08GZX91xkZt4GQk029bDBz8y1lF5An21LRxqsv4pBb89sA1/vhHPvVlc9d
6Ig2ny52a/f0zyf+Zfyvo2dQPOzFpHNIAtvGJ2QSIf5n4BzMJm6dhO1OlBXErCdA
NlOfR33bRvgxtsRS4cuxQvIyWpxmnWK05rd/+VGce2d0tek/Jm3matvwkH221wSb
TuvNXemGZ40vjXDqlXKEhs5kHNG40PpnQFQL7pcFHZdrd97MGOTo2VTUbA+d7OEu
9uft/rT8gS15dKIag2x3o3FmZkjGCzq+NPumUSljXTVdNMS92GYeKv/u2keu29p/
uwW86QKs0MLG46EbV9Ikud1GoCEaHQ08HN0eddn9pBXNan0yZNWmB3bVrP5dRVuh
ze8yDgZCGuvfCtOpLWr0XNlLnhwPY1wWt7p7LBietHLyaAe8KJikIsjCRBBra1G3
sAZaEDAdyaQiLxFLDEFt7vA/RcHILb2apgQ5G3jCwfND1ZBM2NDNK87JFjvLxe4f
2Oh/VtMDbj6p17u4+9SmnZTZo7ACyf43lUdSXbMuK9piN6pLPE8pldjhra6bQlT2
WAbzPdZ/KLvOzgFvMMQszXlGoesdkig91+WjdB/hQ9juScPr+QCztfdUCa1jluEq
sH92y/hhoVkVAR+8xXOm8e7PozDa0whjHAHViq9mTbVhjn+1n3yQkrjY5Rzk5rpq
COhlIIpgzJsf+c8WS5+JCKX0ll2hFdszam898x+HHGTIZj8Vqu3roCq6aAYT7QdI
xfv3ko3bC29kPBtXTlPz6ukJBrJp0q9PY5eoaO0fc4P5MJ8EPOZdFsVPPeT4K8Dl
zcE2Sqh/MxLsT7xOR/1QHnRFW3Ce2EJg6yTfABIKCLjZd/+Rrbv905VZ+NTmKxlt
qSM24hwKoYFEJJdeQGxPyABtMj2aApNPqlkbJzy3rodMRbvKeDEDZNX99K3pHjzU
9MVdFIrFFXuMyw+cStU0izp8iK9gQvN+mR3prVXi97cdOJf96YSf/hYXS/Jie+RS
MWdLXqzD91qBpHWxtO24v1SB8tIQ68u274pdIWLLfEjIt/CKfLnQD9EYpxj67dsH
TFjThiFZefzWD3FZCAe5+tsxlx+YuT6i5K7/0SMvXS0e9JVJZ8vepbHOA62Q72cY
JTEl9y5iLu2uAFshB4JjvlReYl5i7spmAsuZvF8F9uQrQ7U/dssn3dNbeynpEvf3
xafZl1a+OHT0gT5m4DiPbkKAMaiNkVsW3AFgaIl0zC9lgabsp42M/yPuStzIXFqO
P0bpB8ai7hXBFw+BGU26VW1GYlwJl5rxcQddBwlhbiukrLtqXrEgGaJePXN8SrT2
aP2Osa9T6lSRaEs8i9LbroMj5O8KJ3f8G9XAwWldaHM280dn6J4UQPkdOVE/vio/
DmP8ApOPvJcgQn9lduBUnI5rI0XkP7gY4izXxZK3aNPowa6aJyyW9Q8MQxRsI9cl
617vKlB/6VV2MGBQQwPdR/sT+1UX7U0dSoWEHpVBwKUQXWWF5PotsbTFFwPCR5zg
9TaWyFUh9fTFSCeqaM63PAjyg+wr6ijTpcvYIXDRvNf48wGxCyJ9eYDOB1NSXxq4
UPVPXirNjrTQeoC7KeLNA9BA7FVIx2Yjc7Ckh3nyP/PhOudjjjYrgE7RjIh8/P67
bHyfdd6pslyx3b3Dgc/ivce8rnEm70F6dl5rCGtGUJ17SgxqWmmFM2FZxUYSm02E
u0jInr3xk2T8O1wPPHrrfI9Td2lG5jmoSy5mTDJ4U02QkZ8RW5UYZHVsPlwEdUhZ
Xem47wpD9QmUPq6bHOZ4nuj/9qGMnL6T9frEfzlW/yHAgd1YGd5G7qOUisul9sJ0
tiBSDKbBY58TlS/PRT8qTMWlPpLACKD6lCIoueRjVcNV+tYtu4bX6s5mvl8KTYwr
aMMGUnHvHvGk3fUKXW/InbAIbzEJ49In9CJuTYqWxSKOXPUcDCtC57tYLGcAyiiI
asfdlcqtjmvIg8UNA7s2uxoqMMA4Akzbh62o1BD8csecSvR/0VDqxemMrStRr0oC
YJ2qi/ajX/cXfVIuaSzf/IyKkNxo5FBG0gHr9I0NLxBK0eniGKmlmAt1n1nAd0Em
KbiIucnF/8aOZFPCr3pFq+2brtnyNrzkJWeerJSCoqJUbc+TKeCSfy2HOyaFZyVV
GN2xg6cWafYBvsgKN4o58EzJc4PWD3DMt9TNuSA02GO7ANIwCarOO6S/EHX56FEf
VMcE4+w5NHQBTgumjkiG8JqF99HxIv+MKxTKS4GJC+vrVXVdSb9dVptJs5pJbIbY
GNlup4+0S3eYBSn3T27XlHnGIws7VjESZU6ojejKeqmNSlSMU87+NPWKNZxGKAmE
cYlzj9V5vunomvpGmIGgPSwZqV0JBpdlE6YIaZnBfR4NZ+5zmOHNmtB5XIVVYqlk
Vz3C5KFnqFsEp3znXeoDXRo0Ya8ajnoA59ljruBKtnjAPhbY3dEWd7mWuaT1T+wy
eaVgNrnFwv+smzvHElz6P/OZ/Wl7xIZXnfE9f0Wz0tkwvzlmDh8feOnSh80qOhlz
YvPx6Rn3wcslnihcbKQY888645tFcMWD7sS8XhwIiHB51yZnH6uDHUeOQNMxdSqk
ZPeC7VNTu4zWQKhX3yL+aaRwYj70Cnyh6gYP9NZ8psV1isvfTgdgxeOem9bKW2DY
aWJiBFRdqQ5N7o7XOSUGgrEG2j+1wpd4MS47i34PfKBakj1pz+eeDmRSQotpT8Mr
UtmCl0+TRI6yUU7g0bFU3ctUlOcjVVL6SdgbW7p0Gszf8WZiMmzikTqFlG/jS+uK
2W5fxsYNq8NOtq+ep8DUaZYYMWkaeeb2eFte8Bm+adsrB3SC8D+tTKhNZA0WaLnV
MGTWVw5Pro6lLHquxK/USotWVDHqUV29WN3vnt633EpygA3U1LPdcmorqEpIIp8p
7JJcqksKKR+G0H2CgSqqd3B9/yMl2U9euflGGms9pEoQgp7mY3XrVSWAK3c7qHlm
gaWiRBS33aEKuPjFKFyEALJ1x+wAj3Rk93xMuvi5sSTcrRe8uZU40F7zr77fAQVH
X/sfBPg/iUnHVlLZdjSpCTDTFBE8N1N69Dk9zrP1L/V3bVQ32/DuoLB46rFKrdp4
3Cj2hnrLTyN/0PikzamFgXVgHDPnYUsAPriTtWYS+NbWrWx4CqxYbpy0JuArb2vs
mGUi2zWTUqNLyClz7IZlofMtztJHsvs7jVGHR3ApfmYJLZP6Jq6PmkAOosMg+III
XjFQOzaSH0UaWKaCXCyz/FGxmg1LyX/s+AmS1nop8ZfAwF078F8ckp+XOuM4iXpM
VKlZAGmB27p6IsO4o9B4EkiQqdqE0sMwF4C+z2Tkttk//LtFc5yDK8uc3R1I5T+0
hXP8UvCSONODO1UzRpXrVPvULyiY1WbGR7A3JLcPSbGYNHmyZMiYWA3oI7XO7yPO
6MrExjQ6j/fQw74gRabsGVffkueZJRvKKi7/oBjunoI=

`pragma protect end_protected
