`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
e81sw7RTawiX6xRRoWp2M0XvMzstBryaorTDDOLwkwvQA06xulHCSAC+EuUR8NZ0
Ymv2wr2Fu9rp+1GyhHU4SbQZ/FqRamcvuoiwDNRl67LxVRC+4SMBY5RMtv0/EJe9
w8OjfCm/QYBqhqFE87Ubjr22gJxHIbIRJsaaesUu4Vo=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4144), data_block
taslohXWPo36vDP3jjCZeq6ulIh1eO5R5xp/ipq3uoomoKZIAcZfXln+HoJNuQM/
Zoh/rpx6Ul8zNYXW1dqmTHLION8E+Bt5RdhvvRccqQRpRjyBN1T9ZbXXlgWo/WGi
Gfs7FdSBsujlPuJLVmFQhaLPWTVcTJz/qSE702STHvtmdSQ+piWvW8oYaJWZXawF
J680bRsZD5XB2KohIL6Snvoe+efe4l3Gy6IPYyUgsTRhY131pDxn7cS9mmoWKTnY
6z/iVV4hBrJex4Mp0rN8s5F0gmoLVDbOOol7wOKZ8ey/cg2mu1oII7P1CcDO+yMD
ffp+jx6rfg/kZ1rkb9gl9rv4pydTIV5XJhJ7qW9SfUGjUa3U8DsH08MmNnYQ/Wlc
tGax9mTgwaAqso3Mfs7A1wfl1lM81I7IWVQ5WC5WpKryoJm7wQtYOKPfGDgzMBJP
AoxF/zmtoDzEn7y+eP/T4zdWSc0MlIDGeJX0rQRTIMuflRwO5z/5kmb/g/imCcEe
kmzdwKraAjHRoDbgWrjAdZ3HayFKGq6A6gNUBrEgyRUTcY3UhhgUKE3PI7Tf1i/L
7yFvNHucxW/Uw8ztJpBaldvaEfV92jbnWQ1/MHu1GHrdnotmL87/65OD+o+4wPZH
UP0o8tC5cE/t1LoKbqcH5ZEvKe3QhoDVK0Wj33ccYe9hgooEq8aWmf6KyCdo4QNt
NkdnGLSjGrIkKcUKvK79WcdA16TvYTQnZd5143Jo417H0yAwO5kIqpcaMNinEPyE
CVapI7AwRO+AhAA2893xEHti2OzOud66cAbUChtArEfB22MijWThp5+g4RCsFbMn
bbLK+PxtXremM5DQsiq5Us6bXToVVGb9xUOLBPoCTnXqqiqECeShsBXEpw73hOfS
d8LxhYwhK9vqbKGuj72/3KFyBJh7CcEWW5/x8WFHBsRg+hYk95F4cxtn3qw+Ari2
jzIqx38XHQntj5pLjAy2HzM8X0Opo6bwj9zHTfdiHmCQ2IHyuCadhk8LM1b+VS9Y
5twHT9yh/y3E2SJw3cn6cbI2HxIcMq2lco4yuUhxjrimtV8oG+oE4v3pgwaHdLJe
KVZt5Fy+IDII54ezJ9aHPn8X0CPZm8qGSmAEc+HKKYCYfFQeKHSkJa4a361UFzE3
HcoJlM/uwy8jBjZkglv2RyZ4e1GyqetAdk/AEmtNHRAxMgPgmNhnxDE7e9UlhFTI
BTnewDJc5tP63rRgw+e/5jy0PFX+RAolaMfTzqdg8WYKnclbnELF6ufz8ack580l
Rkgzq2aVwB1hK+/5soUDOp7av+oDwexJf6iJ4eOo2QxxHK56QYrDtM5VKb57xIhT
swwKbfmepoSGHlgQ08Wt0IKaOODqn4peCuUpv8rjtzn+8sP8QvPxtHsBCj+hD+qB
kozX5yRsDqS7FHUkDtYTY+K8K1HZ5jJirF90lemR2hRtiSY+hCCxQirsVoq/gX4a
V5jZKYvZ7RrYv5cSPvrCYjgN/3cGZeC5cPB8gm501YHoLQd6M2f6bnbUD4Gep8Tz
XoX4Q+j7mn+uJS+i4iglJ87/Gd4RhXXrulqXreV8it2U0DMENCHS5K8fRvoz6zUy
crWgqcZbvvh8DAD6miCuhCEbWQaXKSZjxsIkvHI1DtamykrCyWe20Obisx76t3VQ
0OgByEWJwwoOpPE8R8DmjHW4I8jZqUF2OmgwsJYfGHHwn7VgmmJjgJXmbg+rFshg
DWOHyIPiGrSaHVxKyWzVg3C78xdCh6mw0DfvBpdWkrfcwlt9SvuvP4EingXArIHD
momVUzs369+Wd8Popd86CN1806Jw9S2yAg7lzTkUpZ5lJ77aHo11DuyPmLCn6G3n
Q5swnr9T/ZQt4Vjn/RzkNrJEfHPTwJd1Q1AuTEA/xvaUPq/2Hi6I1fCx8DF9o7JV
/9bQ2lfi7+cO6pI28Ix+YAS/NPi2WjdwNatcsDqi9sr2NDG8pCYU9lo+SziM2wVi
ddwD1XjttfJR3Nx3MX+Atw87tqIpNmyEPxhNxQmBm6sIDMiVfLSwpmJ545AgDQ8T
gY4n5EBm2tcrXyycnLxYEWsM2M4jUoNwWY5z8HSZu0+Jwgalc2ZFBzav/YtIwUoh
kigchv2c4kyWWurx+jiUDrJqC1a7+pdjlwbxoN5mk+j0leSZLm2btJmD6V3euztq
TZSrwVexYu/82/pTc83pUMAy2PgLkMKqS76TGnbfSY8M83IVJiMyZTGbuKyFJxG8
25fzcXBu+mP1WiUuosNS5ABkR3bowKKzzdrd8B+T/idWTEZp+8p++j7fgux9TNv4
61T8WzoC4wLi7pSoabJTE+wG6E070pUd+Trn/tvOkgCKJ6LG8z3Za0t+yqAWYhaz
KZetK3Y8i++TvA4ReQsU9p4T7vhlL8ETRnBxh/06zM/bsjhZDWw3olfheR/mmdsO
8SAi78vP1OTzH2aD7pHSxsnJdT5Kaj4E5OvFOHKa0Fapb+U6s5VcjRNjsr0y1s/Q
y5bU6A9v72MlORss5HuZAxpgiMJwjJcjMgFyttP4K2JSAmCJ/mEALIcg8RUa76pq
66sreu56IMRzesHbivyNdo6Rg342Rm9krfxO9vihhPDNPvrO9S3aVcSbSAgjEPSd
/6+evJmnq+3biJYCdsWGXurpczaYfGI6BSbLJRojVcdCcDpMKBPRJojrb1ULuY8d
4EpITKEdbbEogoiFUwm7eti9Jdclp8UkRVuKM7WQIYOEI5cIsoMESxpNDybq+ldq
mqhwKw3eA721mwHwZ0FgMdKj7XdKdy6YeTOJ2bNFqDy6LMJxhSf2kwqLV2DDwvtD
pO1qguKzQzez3kN0yJBcmBz0YkSWShMtXvs88nmP+sCDzXve47hDY4GewLi+woQe
NEID0B0jc0fM1a9JVqsRIPvtRVd8wX52QkAH8p0bez3YoT7F66ax46XELjyytqwZ
DUgVLOyNM5SM00ehisCzpOnZWZHQwOwXWSwNdzGowzyQTuLF28ZHIEs1Q4x4XmTq
NuxmiGL17F2sKqQvXvDNB8Rs0Hu2FDSmuEo1OgqM74hyJWJYvMqa5Ven1gGpkYDi
qNrPeQ6zMGNgRnShRkTZSVmmKTQ1qIyoeIL2BtfREnJgnZuGHrJIXy9liKThhXll
Htj0693B35mj5HWr8NI8va8QStL89ASOxbGflfkah4+/qh/YGd2udpD+1ktJErmM
GVPWDXvQ3MsTKixW1FAOulJnuEfeNX6IoyZ6rfJkXZbvMKiumTAR3dPR3Mk2AgTW
hau2eUz3tFMLE7WZHsJizFKNVHmMmNLG2UH131hDpuc7qL1eG2qCWcuI2fCihiky
nV8e9EhpgBjOZVzNIVPTC3VUyGWo7mul6DTHVoUVC1PdzwsL1JT3Dy6Rk7bry1+d
ErIA0IvGgXkt7AKNKXbBpBhOY0A4amNAVGemaqFxX1LRXUPOCL3Ke8iNAP+9WuK4
FLuTOI2wfvruDZHu9rYuqHWSnNtGbptU2sT5zFcuZi+xx/tzJ6nAPulnMFWIc3dp
s3VHTHXnq9/K/PSTtZJlYDtGxjfidl2s4Kd/UE0n59OFLgDmILl8HoYdlnaUqh+9
Kx6GzpDOxjZxumBot8xEwzq75SGIQppkpl4DZoePR1fCcpnBM32fWsUfiCr19xnE
SubCnWH060dH5ey0zRgZx6TnpwmhsLN/bncxuOZw2PLFHhuE/2Bixv39RTjso9+B
yIq1JJ+30JJ6zNEXYS1s/3N19zEtfoHqC4EnJuSwcNNqfElsjzXfk3wpM0SDZMOQ
N2tJSy+S8m6pOfWfr6my2lhF9926F5CXLKY8V6jyugC9fFVKFG6gNt9yez8ZgRsf
dA/S1mNRPhrY9lOb40PdIYYGEsJbM435bb0jEaaCKe7DbBEqDUFpS0yLWZ9dQaWH
hefC8lOmw6d5QOwwVDNEoQyJXSFYrA7bBW3X4HRuHynsbMFhe3XfPVZCFABs3XgL
JqnZLpb9Kw4zfEqv+Igxttla7Z3KszrL1enejKxXfVHix3bEZx/BWC6t2suOahLG
XU4uFI5C3MpVbuRE5Um03ZTma4BBrEmFjR2QaKJ5EE8Zce2maEgGwEDSddhX//iH
ALs0odOD0yKqQViijQUtIOLyfj8L/x2KH7TEyyfatwP3bS7EnLHJy7sbH8OhfVrA
nxz7r5IqUq7MYPYRoNXmHZEPPOAzC11JUiPwc/EvcfhfZtUceM1Ye58YjmiJvQVz
uXgKPk7GDTnOU4h+fG/4tTcSJwk5vPihxvUwS4YZMmGvkcoHT0EkhrAzwjyxpRqB
eD8xSvM6eDz3ABM8cl9/pJrMxDTR59KbDpWjcla8Gd4g38JaC5XRRQV+YN7JwbMQ
vSMsmr1necD2i6e5EamOTbhi/1oprHfYfWm98faTb/FnSwC2wAdingjE97BIJgSl
WcaZna8lsqApVzCyZ8UnluvVaqadiehu9O5eukaFoVk55us9eo+ZzB1OEGZnFap5
iv4sFSRWRGLk44R/cpPRbAMugTQxq4GqJqi4VhEOaziU+/ijoE3I3WkbHK6vq3HL
M/GsjBmssFznqUhwDMIlqs6xJQkdibaXxSwyiKvUiZutWoEJ4dtsj4BOW7PfeTmY
a+3s2LDaLZ4a/2RDw1dz5rhsNGJnglE9NYE6X9CLPRwMg3YO5xs9iyKTy7i9eDGh
c/X0xOEn+amMSFvjxDto7Gqy4FL+vSV1TWi1JpmLTekKWywpIVBIqmBpo8z3KOBU
l61Qo9INH7JUpVsa15iq1Olxulc86v0PLnZVgLh9CXLcDm2/uRZpyIs7ZO3D3Yow
Q/Z287YXSY2aZ/M/jUTgdfccA76QxKBJOWcppOIgrwiaXkI8t8hunlu4rL5xV7Il
M2VZN4My3mJMlBUSQdbzU211HQE6Q2UBXlj4uXiJ5ZZPrE8yFrfj5NrnCXM12WVc
cd4JIZog+xj4HNqMOQKrzagOjYhM3i5yp0VUD56C0lNrjorglSgEBG8wdNksEzWj
Ew+KjK80879SrAhbh3+ucEPyDHO52GCSZsi0cK46liZd5ypcccJyKDqGksCBUWjs
Tq+u6ATeUEULC8nQOZBppkiTAvgM4HeiwjTqcK8mxCYJKASztCsCl2iCHYPvS+WT
pTez9MHkrzqw1gHNO2W6bovTfLDO0HB+4VNpk2OcCwgVlfxbVn9pSNRgaFXbe82j
Ws/aUg20gc9GJd2d6uum892QVcg1/ynzZLoMh2LVJFCwLuvqPNkjpI5LafPgzI0N
AfUm5SkGqfvQ9X1jWZRCJf9hRQgboa5xZIHb0IDy6KhCPS75Q/9w4R0A44KFwjNX
p20aToU8Iw2HxmQTSb5tdyfK9v88JwwUhfyipjEy3tTdKQH/KxwzMC4dR1E7IZuG
W/LoL3Wp6srH08l1Bhpyf5cWKf0eSInCzwUITRpusLaXfyn769hzBz11cGSu0TzI
qjUR9k3J4GF7oGioNauflcChtTrJXDF9r0ZZamafymHny5MnwXDHUhZqX8UyjoS2
9aEK5gl5z3ZOxPNamMPnoQ==
`pragma protect end_protected
