// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Sr8qE7ALroQdR4OE5TVOCTKfgSUzLwLYAtAEKG4vKHtDdzNeOA0AyBLRpePTRIGX
tlDDUh5U5P326djtaXGOU0EnhaLKQ/F+jVy9ynPOjNRdgTRZ2XifmtPvtaOJtaVF
Q+GHhHeMGK1evqcsW/DocGzM/YRmSiF+QWopo7K3NUM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8544 )
`pragma protect data_block
uJ/NAPr6W+nn3FZNgthXObGCHTtvGi+fZkOTw6Mizl3pbS+2F6AMq8bwLvvCzrQj
U9/Up40+L2vl0qMszXViVtkUrKk3W33tpU7GFnv0SCUz859inLq8elm6d49Tm5ls
ozRpPK+WqpV75bAYzvDwsTu3FMsJ4/x/8se94ZuOpOD3R//DKau1elPYFbgNrNH8
59F+N+S+Wxfah5Ib80fqij0tH0+2+awqf99hZ1iIeSHJk4fTN4D4jFuZ5OXtGmWX
Q1AU35UxEidtYxmldQn4/hAcpO60a9NK6RVx5QC87HMzRf+EYWb0ycti7eGf8wSW
RJXJQUdVNUTw4x9EaL6Q4mIQEGtBYSSIkGQwdVBEaAcJedvfXWYLcjjCy/2uOnas
6eF8Nevq51Rc07gJGOc4BucQh4EL+yTw/+J1mxAHDLZchLVGHkRQ2D2PCDOUZNDA
i4zRkcaRkqYCJzjaxEV+TXSenLmN2xJH/TAbjehNmfwhJGXyRZWCb0ON5sJxpzH3
oWAmhkTaWrhJEg153yn07tvSI4AJzpuN0G9zZc6o9Fm+gKZGFkqe/vjkFN01Udie
PCYlimB2hpLSHP1FkQVsncbEzi19fwvBF13Rm7GasCEMOudum3ilOX5eHh0ATd+s
Zj1m6TuUDegnaugNeaYFE9mAvxaq3/WHugHffWxOoPOWwvE7osL40udJV5s5jhQh
arTGCiaSazbWUQJIiNv1E0gXa1k3mvge9hPXBlsNOdhIKmRHMa1xVnaq6s+TB0FS
jzT1VOTL8n0J+6fGs5ffEuVOt1Cbi4oCyvZUKTsP9i2VOP9vGw1akwR+JL2JcOdH
1rscJKVUKv4/4jySoN7CmDCYPPpwnqfXU4EzwHA+idnZ+nL3OBjVYkK1cYvNrr6J
v1ZEf0lFtFww2NgXq/rDrRl2SggDC079f2sqrlpdiqP2nMOgqXxjjAkp+aUXDdBt
1l9G189CjknOS/mXcBHGHsv0OsQ2nrRKAOFVXGUJS2uSWJRSy2QIDrr/KWGpO3WW
vspB5gzAPkYqFsRFgMK/q087v0cEodAm4984KB6+QNCsi7ASUcVv9ONUEwYCXqYA
fN9dgG4tsn+240kJ48LQgEpco03LATcA7LOx65e0BfiBm8HJpZ6ehhdXxN86MvuM
J7mGqwG8eoqKuNAkZbSiQFxB0yr10iSUQGsgBw1K6RB6wYcuFFzLNnZe1dQoBW5K
Zq4FIuN4gdvYn952e69Ta3wc9e4DI6Zm8fugPEcjoDZVcaie8Vsa6KLltf5zGVPJ
5i1ca+85rLQgN2gk5BrPjf3Y7b3MeL3si2zK4oUBg5by/G7yp4NDDgw6BJjCdhQ4
Tc62Us1P+oEu0HmqNZa5hXJGU699YldLEZqbn13gUrUNKzRWUHAf8R0Yh+lYqEP1
rzzZdTyJTcztRZoPH2IPcHx1uHHpjYeKWu1ZJQcoSrUHMlFZgbsbLXlHWXkkq5lX
CzDGwszVbXlv4JiFw3xc3WdYyAA5hDdS4cPE0l8ccRXWtms8KG4ocyIqyKdXpqAu
NqYDuTAjON0fNAfMds2yn/BdxWXTa7DayRtp9hClnR3WOteBivUef4yPPAu7NTpT
EXO+WmxeXXMgBwEwBA+3cuHNG7SAGoKq6R3cnFVhZdO5fXxDvquCRXdfG2K7sJvP
TsDzYv6ymqaxRuqxmXPJCVdHpJRyryZRJovB81DABXbmHtB1jrSVY5k0Skb0AbpW
8zJioNApZuIlnzx/bYVRM9UodGUBD/gic2CrQut6rPPReE9lBX1fpFtDDgQkZ4Pd
tnW44u0qH3l7qIhJT8NTgV/VmqmEsiQE7avCKuUETXJ1CMbGuQQTIxuYXQ36xc4y
Dklq8jXqmr1R1dLFM5VfuWXqFLhdYCKgSj+AbjMxeWgvTgS9ECBGzBdmiU/0P9kb
nG/uD2htLd1bJV/3AZGgJbjA09ptU99HBtTJRaaew/iW8CsegM7V8FP98iB36HAN
aotOAFZND4CngXTydJ5pDS76mwjrATICMfUGk1OZBsVnxKW3VfWeuzC9Wl3+GzXz
JtQJ8kxRwIaOWRRQGcXY0pexXo90g/usBf9sZmO98H0gLTBJEkg7Es6QcrmzdbCl
IxGt2NeICzRIjdQcwwaMVWLI4NtbjceOPTedHxMZgp1x5/f9+0k0GhjWPgyJqQh1
qXNcsTXQm739eyMvgqfkHszcpkPrfkp/fRl5Hsff3pnIiwYN5TcY13MlNjPXwwu2
pQ0q+6Ff0PhMh5UAA6PQ4dEcCtxGojYGbowyHYGiYZNfkmwHKbgMZRdfHVmxCoa9
s1fkjnS66eRHMpPGRpKJSJuWHcZgbFZ4rzssYro9yFJ9XhV3BZh2leHRd+31/Vj9
JNwttA9jSXprBG0LylBm6WHDODBMK9VaxX6NkAbmsd8CnScvI4bz0gQaXLUjV4Bw
mx3B60HMXkbHP91bAtSQ6MARY8ow1dXufwChdTHdxRxOBcPR/E9W7HDJS7S+IGuq
3dGvVanK52zj7z7JH8uUb1sxMGNOUyxzcgGrGn2b0JAYEc4BiJuOI2eNIHR0zXMc
+9ARN+XfjYA3+hBECdHrqbdx0YK6ND5UalASfnJ16rPaf6y5u1BYKzWACCElHWZ6
W+LQtMTHsHrhCR1oTKcU+8Wjl7bqMMr5GHHCCA0t6CqfqDPxhkol/TOGcWF2GHsj
pxEruaahZZW78QXfa3dBEF/PZyrN2/RFedOzpUYSf5uBXmAm4Yx7mMD+4sJAdmY7
zT8GxfAZvxVo1zshDy6oYMdnNJoPiiPaQ5DYY+auG6+v8wJAE6kKExJD32dHMpQj
b7TsBHbWIyySt/EqSBZoeTVUeXLEVivk21x3oPJM3jM10/JKiMGQp8h+RJpMh75o
6iO5EqDozRCJgupDx4cjCAWdRrFJuK9Yi+CAVpuq1rdIan0vOpgAuQ+PfKdVuooZ
+uBETCBi+GFMn4eYV/8/3Sgl3CsCbFoReHg6wEZyKk63K1Rdn0lpprHisNEAoy8k
53HmEykCiJPgrUW0u77QyE5aSrDhYjkm8y1dqkuLRnsM9D8wNV09dAh0iAEOJz24
yedjokHe+o2IfE8Q/zWmlrNH1BgoOGhf/0zDNvlYRselVP/xaaW6QHoySUNCTwgn
2OJaQz67YKiGrBzUZ5A6fu7kuNFegD1PEwLeQaJnmRR5XkintTshWP8hc5G2hVVW
VUbayyPI45okSNdBzLe+6r+tJUQU1prVlQKWB7KkBCKkoK1PS8rT70t7ArM+DGFQ
565hOYlXWvmwZFD4l/tQ+H0Im0vv34uf2+YCVYB+uFMJpgGSS91H4aOrNDbo9v6z
CyYhG8A5nIKg54gsmcgJ6xCwUu8I/PEcMvgCV4gq9sCz9+1cN9oAaeO8ie6t5hRL
ZoP+Kd0a+tAuwNvTqerMpZ+j4k2pTyDCVhm9XheS0zNwDCDOhVSDr0BjcI1VmoQw
L3GorKVJ6NPjZvzqwZwf64kEXmLUxBJEyjI0HElbC97YQ/A1bm1Fn0zKQAKNmJ6L
VNH+yfzEA4PqE9KbjO69x0N7Qwq1gJV2tZNDPnjAtUY4x9sfssnKUhc61AzVz8M2
uXUry1tIAbtVod0Pwiq0XOMeXXLyDB23G43yXJkyr+7D7SMpagkQRUwlTwiAPLAB
Wbyloo2dhNqWCFUY0CVcAl/4ULqZMXGtzeMLrXzynQFdc+V8McdDBNt3ZsE655GL
23JrzjLDmz5jjDG78JFIvIsAVsK0m9RcO4XyFjV4lbgEed4MsmTgz9tcR+NG6OSA
2IUYlO7aJiGkP2KwdxCBDbWaEN64P6MxgxJYoa1Nfd86mEp7p/K7x/QcimOU2PNr
EBbkSF9VOpGXpyqKjWFp0drHbGm3h0cOg5kxxs/REiZXP9ifC3ItSX4k9RekiJ6t
wYC2Gs1oi6iUtdIyvwWEQkRq8ISywSShtTJBZir60qxQ4axPbhkF4Or72SdqLpsG
xzkp6Kl+47nSwUmv5gJqFCHDuJf4XIaRwyuxkEwWpqBlxR7Ncl9ezMX4NnEw1WCb
L2HD3ZEmaQYMc7IscMZtHNhjMIGrhBQFQh5R5Q0ROLez0jN3oFANBBAOlQ9AiOj0
BdOfIAeT2y60a/vG9v61bII30P8r/nX54UY5UuCAFMExJWQpy9ojSR71J8w6w7Qz
+O8nEFQYAtyvJx2jUmhLGIQTyH26Aurx6bxr6PyEBPP5lECqrzbWkKuANPQ9iAFy
OmvlX5pSmwkQo9IAwj+YX5GTiZPk9BOYlnVsR0wwqLcGp+iJn1M1hQy9pdVS/UuA
PlCHomLlDsZ0wDqZcjcd//bSKTONlYDSQzELzuQhk+qOgvmlGfwNwR5zQqWI8w/j
cfb8ghuvzzb2dbmQYp7iUUjSTg+UxBTy9JhZEaqqVoNk7bafV3v7X6dZ+i+SYaSp
DowqQlTl9sxlEdmaAXjkW6rh6PNaf6g/z9zjSSlOrWMber4MdATFqxp2qp73opWf
+L72ZjqRN/xI3ZpO1iGcCnrO6k6ahm7vJf2aqLjH0Qd03kM76eiF6cI+rvBRRCso
ShIUvZ9Np3qT5IASXokc8SPZkFJpHIOWgHecTQRSjiS56G+jbSdlKuy1a4miqo2U
Ap0BWck3sSOsT5qxRjgPzIAHf0dHQAUJBntHTa/XDrYZ711dEF0dVobQPmLgJkSx
VH3B0DLlJUPBLxopy8EhEdHY2DV8msvw7WtT0Y2F5A8f9c0PzNsEtUcLX8KeYDdz
D9sH1nSZgU3rzMZbme+CDcajvhNdbG5kb+u9jmnFh0bsKpOP1t4oB1KDcD7KZcgJ
iThwL+K477n3bCtbiFtOvfeGgbOUbTgGbIfUwySVWl8ZBEw8Zxn2ecH5ls3TDUrG
19opgaT/bgdBI7qKTRxVoSmvDwgmScq+iY9l7/kA8PAEtzcfRawEUqC8OMlQ379t
5VGnnJcVC2NYBybnkqs6Wfc2n1KEDw33t/+txVzc54XH/zAn+3syVhNiRAqWS43H
YZIP1avHI0104ElL3wv+l5Zcym7A0VT9R0lmEiNXoXjeUISCTxnd6iiEhuJBOVJL
l9BJMYEmQT2sLeuQDIZtwTJGVaM8MBHroKhhLR/E3czvFpw7k52u1f9mcgGX6tCR
uBgJ0p88w8B7SN5IOSjwdMBP6eumT4WHjF7Y1jtuge3FMwcF99anoISkKIzN0UDO
EcE5Ax/gmSVPlbkdnzMa3tSqOI2pDDa51qdbwo+Ex7rRI85kO+0KwtyPMomXyUNN
59f+3FFVgKKUpwOBIgilqZNSWz/1x0YQlE1ISll1joyTUATRMB90453cMQz4VyrW
Ul9ltXzDY65lqZHf8z55SqoRZnFfbkvnIseLz4dKkNborK7S2yqQ7i4jtFbDpr/6
6feKt3d8BHoIzeQ0WHfifsUJhtHvNWo1i/sfh9LdIoCncB2p0z4ooqkpyERC3J4e
uz1z2Ugetoofvdqd75pgcOnfbwZswhBNgzhN40Xo4N5cg0QMva52eagPNvRcJ96L
1U8PSJ12TxAuPiJKyLPZMPr57gNpwXjuO9UUAMDnPlnG/aeAka+gWSg4nZ8oku7p
sFrGjpa0i+NpFSzM4CPSAlfPflyCHxswCEWYFqTfHjKueXcben6Cncrf3jZANCA7
qHU8eHVdppwn5HGrJ78fb9n4LruJR79LEb01ARDguzf9aqWuIxL7thIfwHpem3Tn
M5pT3MZtZ+EhBt2CE/06rSw4lOY6lpTu4Cd/jY/IXGPR84F8S7Z019CPdjQJ58hb
+immSBu+yZMnalrzaTF2GSq9d3L0FxLcQNgRPfb/gQQFA6KpJSUWkFgkQi4b6988
lLCULQikQQg2MOIL1PzVKXYVwYf3iOTsvQCXM5wji8+8t3YI/ojT+8DjY9JLXxDD
kuc0SZ3TFlBysTLhKS5L2M7GAaE2DDE5FeQ4OXdp2I1lxl6fNHyIP42lMojTHRbm
ygaC2l/Swn0D7yVYiwXVOEbBzffLz4Wzds7DQTBgwzZNu3jYOZcB4qcqqp23Estp
5q7dCUh3XvU3QDrEZBbcuzRvZjbITaoM+dKLOqnT9d3xivCf4NxhEom3WNdq2CtY
EA7qvOq1jWqDidcE6UCwNTSMYapO6TzshMqPhMG0GAEelwe90oCudhukXwO1QBX9
z43RJkfQKoaitZ7Ifhj+zoujSGf16rt0HTmkG6FAm9dc52EO51oyCHq7teFxepVI
B6nRGQ8cJRdkR4oJ7E/IxZaQx+hfIQLOviuCKqgHe7yXzcfwpAJ00UKmcIaAv+SN
tuk8iEc7ZxF/dh7lWyaOeVESBS4B7YSVDAr0qoPIgL+U7OwlOi/T7s8sR8lfcrwk
+eD/XR57xNjV665/GweG3wq/b8tF8Bz27lA0o4rvmA6OimGLniuZQlMkhzlEU3sx
oGBBo3JN0jIKuW8tKDfO20smYscOiCa0oXTUtuUcNpgrxL6QT3zw228JZK/n1nj3
HpA47PWiQr/QnSGcaS8HH+s67SUtm0CTAW+V3ZhSxJN6tyH9ymW0+O1o4dGt4H27
Do/TFmo/oq2LCkSDTHmmzhA8XPfxci/siqIk1fU9RYtE4Y2ghICsxhWjc2XE2gku
UvaX/brhLusIlXnubLgFWtADCgfh6JBlHfMzzH3KKmAn6VrIm0NC2AAlvnIDqhez
VOYfBa1R4qhBBw5imT9lNt/FKWCFsoNA45MrU7IjeqjQGKKlNBEqQ8/0mzqmnIXs
3WEkMUXdYTh08GtjuWniCqnNyC9s+6FayZHB3WbFOjuqu/EKOcmJzBr3wIW5JrdC
+5lmE82RzmTYD4R6rWGuHZgAo7AGppL+YGz7mhhODTliUJoaByY+4x0Ad7Ya0CUZ
x/0BDQzte6P7HmZTEu4dxWZtPWWwJN1kyDbuJnJmKjpVrcdr9l4VQ7j87dXeXnze
d7GNYS73yoFaXVGDPxtxIyplFY9bw7RaCKds3XGbhoW4ya86sDm3zF3SV4KffMB6
ooPr+Um5urTNndJJiJAYjwTqobsDgI3TkEMO/JveNxPu8G5xUJZbHt4OgDThV0wP
xfFastDziP+F5Sl407CQlKiAPZ/R1YY4z+OGMTaQ8+Bd1bku16PyY87JSBB1dZ2l
GaL/QhH/vDpgtuxfICd9QIAjP6tRcXMiP4U1TcvRDO+LySmtPwGNyeJ+HsRgsagd
oZG8sd02zyl6bvLLdX5o0LJHxQj4WsaJQMGn6z9JowgwOve0Ubb0VsETxOEd5KYw
KHNtAczGRFqtLB3YO4zwabNxg8wJFs6lCC5VpELAy7s7E1hiqj+N9giMpZnKx9o+
fQMNUH9C0QUeFlQimXpNa39XOmcOnOVMVuuR50rzgaSCBZ7YyGuYVnd6g45JEZm/
4ZExsWEAliB323GMA4h+BqCoikgkrvwLzGKB5Q2Fo37HhJfeodzRRiHn7/DIBRnD
wRhHiLS7TOpGvf6lsI7Bg7nLZkCXU+F8l29Xh8TdSTuUAX2qNG1PaW+qYnF6bqqy
fCQy7Dsb7jHw0F2zuu7wSguAK7YGt4u9ry43TF5EufNxRY8Adr0yC6h8fQe6yhz3
hcB6xq1o0CxbggQJe/zN+WBCpQHhOLOpBmGe9eDG6lULHA+Tk8dgGYkVK7X/HqjR
aBc2Mc9GIeWNq9ptuQWJ+9e3pDBDGC1TXiiVB4na1LhSkzV+HPMJzJ4uUBBzaDnc
c6ophmFWyUr3zvYSUBEXYViycaoQV7OJ8j3aq8kw8Kh5V/YUJtT3izUfKxJOepcH
5Bk/XQR7aJ+BlYSjPpo4pGsMxJGHPbyYcHX3UNDHHihiRC/cblMgzTFJgNIDh9nt
G6FsJa2fdTLOavGvN5O1fwY0HT76s97RE1zvJqvzNiaSsxyG/6Fmwcb4MPLKyr8D
EJ7O3pwfaYVCZb3p+kAsOVNxRGphOrT7Nh/mbPbeRkV6D/a6YrXIl9jvUyIZMgGm
i7JlGtS6eY83hoaLUNyg7tAa+2cE+q91TVqsDnh3Mg9MuOTOvy9AsHtJXxpw9T6T
Me7Z9fTkm+AOfD5dhtMpJoWr5LMXz3MwNKjGHg7zmoQNh+bTUzop2hhZmB1o5pTI
l4Hm64w6Q/Xjo8JEQgV/td7JaVBAd6NMHk91n0bPn+PKRsXYNksjQZXHZPCf05IG
AbadDIBy4EmEseYcsfJH7peYrMOAKGvAjrjavScpnrPp/fGiL9HOya1Wh0thX40O
hJgAt5enE8ZJFBv49HZ/wXMC3js/A1Q4QSudRmev5FS4hhqUzWVP3AGpJjFgvKXN
/wG4FQGqIllrjgmhHnE+qcax1V9HbtuBfdNp6aGhyMmCF6eXQUUnZXuLge5jKRwg
KEv78lSAQcPSZoO6/3cOYSaGLAbX96Mo+pzlSvJRcPkwxlQetvuZZnxXG89YDYVq
u7qpz1BeKsE5kJpNza7cJGPb/lvggX9Tbc10uRAzXJqALgqTnv467a/r2hEV2Ckm
Wf2UaNohlB0AK8J7ODnPhJb5SV2wM7y0FkqS9I/Ourgw3u4+TsqLSBAYZ94Pmq6Q
LfRPsqpJwR1NwrCv6egrTQ4gCWOQgdDQR/OPdcSEYvQJ6X3gMo2vJn/1TOBBoUm5
jv4uS4Idkalueq8NZcKEQP6g0niCPB8RA5gZ00AoxTAnm2mtU4MRlcqbRTuFZdV0
N3QkSK0awgwGaprjswJaGU+7eH7EbRAwgJKGxyZkiDfadMR7WiLXHax0vVWku3VU
UJ7/kU9UagZEV2uOdwdmM/J9DnSBSBVbLBa3U7zffMYXO4oNB7PAbtukBbRTKOjM
b9oeLutlErKbi3kv85RH9qynEzPSgsJ0LDmwZZ/bdYel8pmZJ9Uj9jfFn7Y63rb9
gKSq/a7t0GM4K5/f4Eagtfa1mQw2s18EFrdw939NiO1IPEzZLwWP4BpWw58ZnM2n
qhz/SEyzob3K59GGTYe4SfWG9YEW9T99yNn/QPd78yodqSTIPHDb+IAxQhEfRgti
AL76TBDdB0+dA8biIndjDGEv3FHAS8Tjf/+JNWEwtoL/N+uR4SGkEjDvwEv9iKXa
u2ja9ZWrqczVMZpJYEKo4HXZ+oWHO0GzEHyddQoGnDaZDbUwRxkDDFcFLgWodlCv
ZIi1VP4tWyoNq2oArHoePuRMdbfQcssmMT1S0ZYgo4aiAmt1U5qpPMz8ZXun/pQt
Fmy2nDnKEdFqQw6a4kxk4RuiG/Pw/tqO/fGT2od2gX2JByVoflwDhLIeMCZwLBG8
Mr6+i8uo0u6XWLQkimvjiUcE9yaJDvgbWGbizzJHgAZkonVw1DPGmoi2SlEOJIJE
IsLOwWPgWd97NUOk//2+lB4PPv89y78WcflHLvLon/Kdma10Y2OBALty6/ntYThw
/k0w+HgYuQtTkqJM9ytdS9lo2sgXxKoT+5fZDLHo4RXtJ4cpkzv6nWk8MJ4fvJxj
52pffLgEvXqhhbPTkPRDagLgVS9+U+Zt4yt04xsG0tLIeWiHcZKTkxgXzELOpMfq
JRsGh4vPUtKn7ygvDhEtTkxPTqvAOtq4iRFjml/0E4n9Bxxw5MTMbapAY5zY76W+
1X0XVQYg3USi+PRC739EQQSOCJn6I8oi6nV+8wq2S0h8hHjYezyUvKMke36GpSbr
m8f3G/iDQsv9VG8KXHJMQctcD4so5Ajz2BC2LfjFPD4StfDioiW1kmVttdr76bfl
F3MZG5zgR9Fe1WjDiCyE07KD4mHiKYnqIcj2qKhCmO/er32d/ZDQ4lHdoSN2mbWp
6IFOMyqjlb/vbQmgwyxu4rptt4NRZxIxCOaLG0sAvWaS91PnoGrcFpBypfFQONqZ
P2xu93joGK/5lLJOiDaBnQrI5QE6yDmMAxax5rBNzP42u21olt+xeBBENHTZu0u0
IfHrk1w7ASOhGs4EOm9XMnUKuKP9YnXo2+VaeMCiot9Wg4yW+o9UqMrjR5GERsc7
Ht3W50FVVHqi2jc1ppgMSKq09gbZ9/iRt7pE9EErYwKDXEwr3DE4XdXavGvr7esO
yoeLRIVKtJQ257nefK48c0PZB0c7O06rSMq/ZQwAx7ThGhuD7maLSAwTA/adR6VY
bUMG/xdi6ZNCf19xwbGT1nPjwkpmxjhwOffLfhZgERldgX6x08yM1g1pXcIoGCkA
31GTeR6sR2v2LXl/EgCVegxC4mMcFGpQR2yUy1BYi5xeaRFlklXxH9R8B2d/V142
cbs91Omc1eogDnY9bsIPhkDiFXu4DhFfTHcE9846QW5gcKZwK8iS2bgnnmPEOdKy
JiS39VOpZXwbrrtRxnrwbwijF7o5Xou1ktxwM0JAZhuqFA6QkGIy8ulGZCxR3wkk
zOiwqfDq2rojA3EXFUpegmNcLZZZmhRz8MqLmcT26uMHL4HTsxzEZyW20z00MrfT
yA6/ctcRBKLPtOwLx4uTMighqDFs0vjjygOXjLbpsj9wWPxmSsLstVpZJJPXSOKl
Ld1MoTp5d+6tZN7+n7tpuZUEnqxGwD9FeveCDU4ChkXD992sQ7FWU5AqS06HksYL
PQgbFIFhaFlYVbvwfGHt+C97IY3jM59hSXk39sxCN7Nkc7LgtpM5wZE9r3eL+KPo
DLcujBur9LdJFNiBSmrR+Hvt7vG/gvJ/R0MSCz5qNrYV4iX+hWC/nLRmEiR99LrC
YAtG4x9NpobbIgO7imjy+ySRvrgwxHd3zfTL56xJjqEaWwgvFSfQwe6lj+HmBcFr
RnA2HwauXoYDn1xMrWfq1ZyYIVjNlTWqJfiO04JAIUFpTXPVttpVQ0nSyasnKm1N
KZGfN/71UgW7aHi+I5VYRhVy+/5VpXNGQp0+Kzm6w5iWWID2stJU2pJXdgRPOXWw
TZWzR6g4HNmw2GQX+vUCsb5X/jtZXdmkiVDXjKRtX2JeZz5ytDtUd0VdvHjrz9E0
GXNDkRhl+sMzjlv6E37s4oyLr66iyQHV19kqzxy4a3Pwt4waD2m2ylYBDCbNzO12
iA6c2qGHC7WOOn5b8VMyVjGQBWtFHRqApRB+tcAxMgPSl88cMKYa1ymbhlf3F2en
dFZ4B1L4HLGo7cdGrq+k9ZUOUFwWVZhocY9SvZNhhVKadaC5TCfqk628zPB/9OT/
gkk4mAMaDmqdXTnraA6bsa7yPF+aFPQW7/QECpJTXm8/yWcLonA6XBef5emVxI7t
PCmnccCcwHW3W/RKIeSwA9Fni6qUuFFl8sN8eS4/CKofStGplauut0fhv3H9mfXh
bNiaBk90GT3amaA8UDmGEqoNmkk5iBCfSyQc52T6g4nXq0c/jt1nSmBxTwEBV6v5
+ni1VmGiJC0Ty/C24d2E871ngXJJYVYSVA4vvHQMgWfqxoFX+gbQmhs8ri4/PQYC
WMy4xIB9z9AAz7YQj5Cy8vPPvqQip5RYbbyyZj+4u052hssOkhhSZXfzOta40EEG

`pragma protect end_protected
