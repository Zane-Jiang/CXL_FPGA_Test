// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S1yHgCyfg8U8Zqlfs+87MhAAlc/U0wNbl18BWnfNL4bVcyQc6YTyjtDgDcOk
9P+T1llz8TZ7aTJFui65COg+ZK3zri8FFI2H7QZ7cAo0KEYynjv+2gAUMUT7
AIDo2zaN2uFlrtzeGBCTjdFs4jnrEUDos7nMZT0LDD7RYUfAhUCTl/ZEpZVo
gsj3m3isHfKXM2I8HsW3o6sMzJsSnJzf66u+OMh34NUbT+x6F/mAObR/wPKB
1pLt/8NQ7QqQRMM9P54OFjeuq63vPK27LVucSwEXzAq34ujHxIkV6EA9HCfl
dF6MuQ5Kx3JfbS9CmUg52WtAOTfm5zyjIw1mGzIddg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MBkiOuoHa01oMqKMXdGT8YwA286IPPVZr+xKkAqAVMvytFhYd0nKo5PR8/h1
Y0O7fxr7mq19KcU0DuugRMm+SmhQP2vDjuFoTjf8TRqHVT8PzrBLdZ2T+gnk
zMdshsXt/FLR0RLwz8UapglxboeCBuz461nrrt4WmsDpgaW3/gnp7l9eov2E
bPy1C9psPpkydVgAySWDI3orYYhRxyOYTmOVNjee6v8aaupno/AKE6wZNGBU
o/aPS/NRVFGAAd5E0X1OxMSPelk98rY3IntyF3u81U0/78NSTY8NG1bpvznW
sHIW+L5gSTLFMt0Oleajvi9zXD/CukEd0hJ7Dr3EQQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XKIM0ndK+Be1ZvuIs/hXKtqtHNhUO/4wavdilm+k17RtnYLeVHHyK0aIhu1u
XJ2iQ8fuNPStGi+UgH0RLGpj0fW1RwKzQF8eW/wq4V22YQCauR8nccm+Q1XO
ZNwKOny1jVgfQFRMsFT4zjtWo5++WTx8JeF9Rp4ZgTPpLfwcxkUq+HSCxuf6
4VLXl+2WbFlU8FI51lO1vszQ9ZePy22RZ/hdGrH0zDl76dykzDY6j4GXSiln
GxwEPkbXKepMBdXbG3eKwZVqXHQ+xLD4bnuM/IcPtMJXbL1KzlDjReRdTfum
x/03tAgYklGdtjKY3i76W11F8/1jXgFN0HKEhRbEuQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GZ7sHVvATcz0K9zkf97IPInuZhWIRQ9Bbhj7C+izKNiPCzYBT23EpSq+5jx4
6WythOS9zp58yCLoEq7gJdy0pbqgcsoByzP29wdwlrXvDvHz+GZxxCzAfZJc
xsm5jycfx1hMgFehsjj3knMzarYL4k6LVTz7MQsnuo06JL1Z19o=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wd47OjpfjcapFvFY0aqN8TZ6Edbv1YHiyP/bQY23jpc3EVHDvnR6W2aKkIIr
OhRX5cQt2lOwxfda8I8jagBKFIcqcbcuXtZHyOvyv7Rgx4gSb1y9qAiBXYWg
P44wjixAyTfKvYmVnsCthO5uZEI5JSilaU6E/1wvBhY01aeW0rakNdUtV5qt
+lUY6R8M/bubBCx3kOLAfbQzqoTclKmy/vDLnBwm0NObxyaWCpERFF8tkEMQ
kJxnelpKYsp+2TtvE89tIwYSbUD254Fu1Dp4yrOEWsoKIvjge88LxFXROsEy
HkkzOpBij/kPHVoenjflp6nDBu1B32tU8SY16ysjKNnEpwZoK2Nmd8otlLav
olFvWTah7790NwWFIIdMu4aBdq1oXxIv2s/ilRWzur2H92rhyfPWqLYudwi4
3jaVeZvognmG3xuQ6EzEcJpdBPiYThrkjOt7FJ3rgoYBFWF+XEZm45BuC2fb
CCucZgH+jFyKphEOHrkAMVYYzVFOjGgf


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TfhbARCG/MJt7xFIXKdY9gsNvsFiGOs2F9y1mM+rlijwLIFBYefhPIxjOuTG
R1hPkgLLARWid+9GHlcFhM/gAiSssn8qpe5O+Jp5DJkd6SXXMII+fVKT+UDU
joy/8dlsuTjhHbNTat6h7wtCxi8oAQRVHDbpirI8E7NRuT+OTUY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rdSebQF1Xic++h3WQsHH5d6Z0zqguw4v1o0gkLFARaPxIBIYZY45rphGx7Zt
EZ7kWfWNvyQ0BSjs+kAbbZhYvfSujK515Vzy7bJWxmXniXVR9SIjiTX7deo4
HibhIiZdWBWIDFHc7EMyp/nZFMMHKt/gF8AFoV++BmApqZnX9Vw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 5968)
`pragma protect data_block
H/JDHcE5crX/mCl8oEsWDDb0t18uW4VWVGXdWtQqrcbQUn73LbtECh39KfMH
/R7CLlGxKoQVTBVbJVzqodSUWn7DQ/mdVI9aUMS92XE44fBdL5MgKoaXYijb
ynv/Ni4usGFNqfhWM/LyfWdxKOdhUfNk4sWMTFOVvb6gD8OocmTsWovS4dfg
x/5ckqyV49467JFCEHdDX4tfPzSrryumARwZWjZ0KVAanLjL2655BZER9NrQ
Lqp2WZR21RMnmnlQH9gNc/MK5B9hAddejFgBuMf3vRPRfxMaqxCf8rIPbgN4
nK4vwoMDTFMiuKiUiKvXZ4w3eRz64M425yCgUoGnGKPYOVLyXV/1nqbYX0O8
MgAc2E0PwzFwGc09DNNjYhuK/NUqx1wsCoSzGW1JrONGApXJ3Mbhg0nGbDDZ
eWHfaeApX0HhrG/2Szhv+ZbA8/v1JUN2/zoOF5nVr8a6es9pDh4G+SuEtQ93
1Iqg9pWFQS5hQVXeavr0pUGohdrMMTjHWdmTwn5IqdfRxpLRG72Xt+L2kHsl
Ezm4ctnyMBLFom7GqX4rXy5oMx/U/mCBpxxnIEBQ+Ru/VXm9kqoPsagrB3za
5PfQcY7nJHtKJunhHGF4xc4vv9dMWH7sgas0e0IPJJWnJwlTDSEtCdutNn5m
pThgcnMneBF+ckf7UvEsQs8hv9XJLewfMnqh25kFDMa2/i8ly2dfTYFQbCth
kQFxAQ1sChC/IgdwV3eNR8hSSe2zHHr1gks8y4avvwy2YdAMuLFf4PXt7NTP
LXpg1XW9v3FTPxLdU646YNxGZ12mmcVXeFx7dhZoc8WEue6hCUmiNmXl06KL
tYlo3rf1XcNTlmyMvcCs8CurWccjAspDU0biqfVsZDVhUKQFg5isEpyaKLS+
Ew15sdAvkQ8KqrDW0VBItbLkQYGw1BzztxVNJFkyy2m/jYu5jxce3u/DXjKG
j1gtUOJRfmx88rZNVe2jhFU+I0CcINjWP5Tt6rYZqowbA81fgJPII1dX+Zy/
C3VoAmTnjNFgDr9Q1uBIw/e9374izPGDWGa22dmjX4+KizCoN6K1Yc2/1epZ
ddVg1W0hMchMc+fx3xeXB+iV9yMLgFHrwHPKCF5oGpazTtZnNAvQ21OHqkDq
8HU2zdk+g3sdT7rwejbm4TJ3T2pyvcS4WApYJ951CLxVh5NXOav9d9Wwlj0L
+9b6HnW6IGGLri1MX9zFn/Z/7xEXVZzlybfQQyafcLANebz5AG9jKNCQqRJh
VZtGcQ82dHz7S2tgRY8kiVcsHUG/NwLcZfqyM4uzfDQrF8n5fW0pAho1wPzI
nNgv0VoNQAGC7roXbiqv7kjNe3bw551jRhg9QkhtFaq7y2nMjrLp4OjYnXxI
nYJEuHYtgZQKf951w5lwyM0WgGGB0EbMcugE0LdR8p4SgEuYBzNr7YC4AdU7
qj6tZx2bq0s4tLmZhdthGnJ9BYVxtmmv2EGycMkjKuUuPuJC16+OZIMSj+yy
RVli8IB3GbyNKy671qGNU70ptqXyDsUGBtldK1fai1uO71a6yrTjb8lfIUpH
6ytTE/cgn3xg4Q9kzJDClvKyG8DkmknaRE2Cx2tDa/+0eBVpbdpuk1EBgSf6
bjLZK8fUqfH5coPMBoLMLcjvHbba/w8HodzYegDKrUKuPHdEGeUB6qcywdNd
d4aoFYOt7gCkJWbI7/uxqjHzvd5krWS8/vUPEESJ5SnmmO0b7ekNH96ZICrR
x6d8DP/YuIi0c3/b1SWJedfiVw2duvyUkWquJBn/e1WRFQ1sn6LddW8g2oUN
gYOZyqW/SUbH7f7IHn936mu4zxrug0ak4NvNLSJDDb7nsb4nNshPeZW6iKVV
lUBuYzLaoHp8en4ONR6SFyixqjB6KAt7CcPjaMCMgRCxZri7V9S+GAafHERX
sTyjxUt/cSdAYvCCW8d42vegTlBbHN3FPcTwbRcRUr7euFwbC8GHKxPf2xdZ
54Z45T8EXTIR0nvyrYtWrqWABYg8S47YEfG3xyDgMWspnwqozWYaTKxdfacM
hIXNbdFGrv2J92KBA1UN72vsC2NGrLOIiUPw7SORJO00OgZ4PDeX+Su7LAH3
KnXNaQ2x7qJp9NjNHWK9mgDYqM1Go1m3vYQ2UR0Y/wPFmKhRpKkz+QD4Kpx/
EenIskmsEJFM8vshE64gEVzIYszzJV971E7huAdnS5/lO7mqrUsy55OsVN8+
Ub26ayzj+GeLP9mPyuNieBG2dL1/ZKrAJnd4BAaU4prY4oSCcX78S1j6KURe
daemjKwSPBHabxs8vSpl1h7WQsi2GwRr4TombGiPcNArnYem1kc7d+ZxpXwp
dDdEIR3PGO7J75wXHUptXVyz1noZ0tZYejLDf0CGbHKnFc6bY+Elg8GT9jdg
AQAkx1gnxVlheX565/CRloDfwM71K8jDiHwb2ScUM/zz/MGRrxLplc5LjBMZ
SLiQ9G89dR5w7PO+gw0MuaLu5iX2vXdF/Utl2ye4hGm74EY0/OwoqlgnOCY2
/5r/8P7mhhIo3pszpCxyFAEYQX1e3SlOwu+2RAaS4Y/Ihx4uS5kosFJ4HSi6
x5LFlTQUmNn4dF2ou0EP8FQwDYoWweuxQbCFL4b778Zqs1TtZZ4mVt0H3qNx
FM/ofPPe5QPNCitfdAofRA3XbzfCIsgQ/rGp7IVZDx6qGnahU67Qfo5UPElv
VAqjudxYMg6aR8QtKU75wzeputTqYB/rRBj/5cSCfMRHszhr8oXidUGaDFtZ
uNBT/rOJkZSahuXqgAZQFR8b4SIBNOlCT0A0X8XuwU3Vbag9htCZ9LTvRHZf
EfFCgxHl4SbVqLBKLmyVLE/EKvhIXOepHRSXu4uiJWZoMpU2ENoSmw3CYy02
MBCQkUPM8Bny4Chjrz3wWIBLnp/+EwW0bV08OwvVi/UgNPdlWiMTDSKnqrsA
N4KQZuNdVrkA7xkIfv5W4OOr4F3vo5SomOduRv92JELNlMozDhtYJoS24PfB
NTPV+eJF1BcPoZ5fxTebalrXUTGAusJBrisYNu7WPYgGDRW3PpaiQjud1O4n
YzxyTGbek3jUj0JzRgmXVLqSLOtMbiSllAT3IbTSag/pkIPAM+j5aSV9Jj2c
uuoldG1KPcOfy5o52A5Bb362p+UVQOPA5gzqsp9iIHeC8WTPEwakKF+WuUEq
Y9MJ5TuUwbpM8nfkurNGHoaCbxOIPjbO5tD5PYI6gC+WzgTSGfFbYpsWezaT
fRg3joCO6Q+Km+uph2IAahcIThyTEJkltnfF23BQxLqFHF9gP+oYHGuxZ+S6
uPTixWO6AgsoA5njsCQQl0oFYDDaMEVVCKrl7TTrLUV9q0eOEQ/idBB0R40D
z6kV4cX4aw7J6EDYom1g9Z8fbD3SUr5q5CitPNxC+GDoB1YLGNy0icyDk5QK
x3/ziGSY41RBl08IN/PpgMxavEHDzuII79ibDIh7cXtb4ubQTDFFD6c3nkDQ
vrGSQOC49Hga02n6Vl6dqeb3BmZrQpPcszN+t3LflUQznKEdeBRGK3CqTq/4
76X7EYRF3bRTxja+DAMMAzSikoi7kTid89TS2Q0cPU6O+JOQ0Ff4ZOhl7mEz
RcF99e0MfUS0RzkSbOkFr8I3C/TThOL/pFHlK4PQcUsdx/KQcudAXHRZhv+3
/q4Ig0r5UO5zgucrEC/F0b0X0WzE3Ci3YqkFaNphYL3vEz1S5XFhBBjKL45o
xRcjeYZxrBmmrVelSpPrPVVKBOHZbMWgmnvlqy/MvaS+6kbcUStw3WDC6V0t
3nagnr0eVWMfqgQ4Tmyc6cvXeCI238HzgfF/HWQnZBrx20elRzK3tOwu2qUa
M8aOHBa1HAJCh0S881HPobsy5azWHvLonMTHh26KPa+CHJwBtZtBljq/QI3H
5ez2evLz4RM7lA1wwYI/WpzjGiP6NXj2lCaGX81NKzQH68rI3SisEx9tPGt2
o0LYlowSFfcvipNtfswsblOeRP3V0t5RpiAnrAjpbaKGlyvVGvt5rDreaOE+
XQlG+YxW4wFIBmOHPwrvZLCS3JT6o6at6cIS7JoGQBVLcW72aFNUgZV+hPbM
YeugmGsMtyzjf9C9HROAwzmROkDmnMm3g7VA5TDMXsmme9+n1cPu3uK8KDnp
smcemtWlwoILVKxUFx0DDQrhdu0VxpbPVFEZrFw45Qdwx43Y1hc0iAQVvY6H
yYVI4JpfbU2fuwRXsQqSUmmX5UXOr+yIyELuqcxCCfd4h8lIUT1vYMz39WwR
TY/5q0o2Jkt1Chw5l40ClSwJR6bsyazu3SmjMqqFQdDaOd0I/KsLUKbgBfR0
K1LEYyljve3FJt+3h/9gnhafNEfVDuf7SufXa14RgA+nkCEHkx9gCVgitt6u
8zk6deNUe/Na24GiQBCnOrOHB/UwdapDI8+9KeiwD0eDYME1PQpaN6E0j14Q
4FUFHCx2ePTWu6pm2hNHUcfpaxwwwCRzQuOjY0AVF2IYsEnWggHmTJqA+4b3
4mY7hKljUSfQG85UJfs6JSxHfqFaKHTW7x2+DXIRgmY5zwrCgCUyXE2Rx8Pw
Ww7ku/lxX7iapdAv9+mKOubR/D2rJHPH+Es8zT6nSBTkfIyN5zpV+ahFvq1d
sp0C8WHN8QpfEQ5Shh2kqKSWO8bTCfbymWvCL4Vuq3v2C77dWp6uspM3hIEJ
zggOLEmSAXbVjKtEMeCsGaToAtOPxWqBwuP8sLzjW52jKiTNZblq9rYJE6vl
BP2s5tyZexAKy9jIo5UIcwVkiTlEi5sf16fOF2caJWi7SGB3d8vqWVT+wRQ5
Qst5VW8WbQSm9MiVmBX4d5mxo2qR5T5RjD+lq6Tr2OpHCy4oefhnM0HADYp6
wIcUCJg48FD2dJ0QkMgSUyL5h2YE1oHpfovYEw0Q2UhYG6RGwBVKfRsyueG9
cTABqo/Pzb1q0cbqy9uM2HpKLv4lDRq8fvdTMZX8HYzHsRyFKL4AOE0nVP0T
NuXdD3Qjpq+9Zl14QgtPMJ9UVAUJbhdek7BueVhtY1YNjBvpkWQ3D2j0gFXU
RmwgdICacvh9KHugNz4AqsDCbGtlbcoEkhsOfOTnC+4a9u3puIAMg6BIO3Fc
DmXVLXju4dz+vX+sTBo6NegnE+HMJu5WMSzBVhK+SXfz+7BVEZzYpDnzgm6x
NXcDiPwMet2M5dOoXCXh42xzcD37WAi92riiBvFO89icZtoIqhhja/hRvotP
FI0cTkHQh3AQapALgX4MQ4PC0eWhWID2V9cqUSrCoRhFw5L76Lzxgwo96Nlc
+6unG/cu/KioVC5xNX0dWYF27PXKdTfGDKRmJLEbz9NvYyTWTccHZZ5YGzrp
S3fBzu+hnJGoYWKScxjeLn/FZSiG+hA7nBAbwy1At2q3dDsGl2oPXou5v9os
5nKTuI5nzcAjAnhHuGPfd8gGIpcYZkULNjHt0pl8rYqjRfMKaknpT4q/Oy+z
fFvSIIzEVHSOu6wry7I+CyFDLG0O21b4dC3A/0bR6k0tKo8PE8lGuFuxRAOx
PlupoAcD8VDSgbou88kb9TKBfRzwFp06nX4vjLXP4bjvKEBS+cW7Dl9AvCQi
WBa376kbeyDrmYO0AFdtC8aT9Vx+ZFo2ke9ecUXQ6uE8zz+TlPmQhAYwMDUo
bSFUI7BIMNtm1svK2yvryhQ+ClyXb8tIc8vZKk2bjBqqMC2Jv9ieaE2c/kt9
O9PYMInjyOtT1DVR2Q2HKgzrtsFQanXQuVUSQ/KktQ8as7sO6hKRSAnIhWn+
W2/3bLsCWGDetHyw5n07cawu4ryIhtjx0nwpq7+LVqxwm1j+D8gs0pQonw6j
tqaJdmDKBjOyqnGtSlY/Ce104atLcsenz4CSOAFNyeuubDYuJ+tLsrlAMwR3
DYrTCDwIqElS2asDicyQe+cchfaymAHyJMf/rSpHR2bL2jeW+6b7EZlW5b1D
1unV0kQrKardMz3ghWNHjS4rqxmGotvShgvDV5hjUpwq5VE+Xsb36RBEoqqy
ZOwyMYbPfJgudyyGpqhsotqhiHks2jiZDlBu4LWMqV2mC6kXAviNuXXcMtAv
l9VZzKJ898GGEKnZXFeX84WjGgDO8J2lj87TemSWjkBaLPa6rR2pGN3/3qG3
S3OISjA4zbK1jjztjr0O80hff/XrtunOnU337Q6jFcEAed5SE7fVMc52BBaL
cVXRtyo0sBCJblvMAvvcb48TDsfMletQiNroNCU062Amux9xXh5q2HwlWQRL
NPsD+vcc0/4lo/j1Z6TPH4MAiUIEkQ7n1nPrHNPKSMkr1XQEHXAiHpp9+qAO
+09/weDNqqD/nfa4lfYCr5g9Vydmioxe/w4qnrgKmsZmVcuIuxC9reZN1UEZ
Fs7t5r5SjZ/Ax94nkc+WJv96LPV/uBSLE2TVoGS+nvDPW1I7KqIo5zcsb62X
iVPizLPVc6XIDh/RO+L4825mBpspXS2oD0bxxdPJWRMmzaEdHPhqBSzQanih
5+U58Rkwbk924FrYcJqK2RdZLFFwrioDncY8kLoOfrnfzs2CFQ79MfTyoXl8
kQvQfUIDoLcLAw+KMY6ZJcsYttCx7iwrQW/IE4OitdIe3suWccE71JJFKQ1p
TcnD6F1e+hN4wHe0BBaErQ7rasS67+/b3I/gbM/lUCOiTBJA3OJwTGe8tUYV
B8wFKXTmqgvMD1j2yTGfHcn4TjVh9TJqY6ehi8cABE5PPz4z9UfL6uJ78Hc2
KjdAh1shEFrs2ajfweQ4kW8IFktBEKz6WiU9nRTzUlOdnQQa+1K1XtHg4yjF
hy8uPi/YaBPTnVn6dndT8yWPN3yGZBUFtrpRX/7pprXSp67H8WN+qHCfprW6
pM0UmgAI0DVqLmWghRZhWdbAtNbGOXkKp02Cd4g91RU6GvV0dS9GTPDKPyAi
M6T9VC824qJsBrM9Ce49SvbSa/jq4EiaS91qrWmSmiNpFF7uaUPOphAtPBrS
+jtY6YawLEeTfCOGjIO5NU9FA8htgTZMNY8twdRw53HhHz7NViYA/oC0sbQj
yxiYI/vb19BMlLCMmVc2weZbyxSyFAdGsfwnK+FZTaq4gI3bRR4X1NLk6tpx
hDqYZjg80VCJ931TSHISQzmWLmQvTe8vLa8N7OrQYrJrjTMm992LpoXA+9gv
Rd5ptEnZ4WoWL62gwtT4jLmVOs4Rv/j4MKQU33RVSyJtWJdtwv4f4bIu8l0x
QG1fHCDmNV7/xoBnzQL8VkNlLEMjcRh5VS+TPDBtuHRTAJnlU5RPH1g8Tu79
3pu8UutTiJvonWU/DPN0n/4GZEmY7RXq/vMucNBtmoIfmw6IEqYnVXHg5TzP
XSDW8NwhGoDNzxhfixBTSfIN2Xecv7tOUiUEFXLyIt9HMgWDtLlqnHZOQ7PQ
kDh4d0m5xHAGNIFCyBQ9zTG7w/qkcT50qMcG+C8AuViknN1+/iqShkRnLmIH
JrVXF7C33L/Nb5TSN/Cj0rnM2dOpTMcZQURVIb/dP8Q3wANQYLnxFZWGm1JJ
AjrXTwkKS3urbxZAmnngRJXo7JYG3hYQihdCya4ybDdg9OYD5eNPq1aDoa6s
c9KSPIQx5B6Xvgq1RRJVYvTAfj9+S/K9wdEwu69jAk6udWAv5d5T88WVSNmZ
YD7n5QRZWhti8SYw0iYbQ3P48/TUtn1uu0cOHGhOaJwSu36iJnAjfPlYCgml
SF1jimyHKu5nL7v8VR120AGkmYY/Dv1lHMzw+zeFen2aowcpR2zDT+S2hFMb
5JoiP5n4x2mR8dlfTSQkZQs2Vaw6qb7tZXcZ5YCNIGx/y7t4UzZIk+LjrQdu
wtw6Wn88ZjU2YLc77t2yMKIc/oG8M7umeySYr7FKnUR5nv+gOLC1wzcWT2LQ
MInV8VXjwABXzGv7ZTg0F+GFxSLDHA6k8+3GYUOj1hpgxzfQ4k/1yw9n1n9S
+mYuDXJChifHABZXtaRYYdycsMwa8lek+ywIbQ==

`pragma protect end_protected
