// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IRwwYp+CNCKSbWu+4CkusLc3qfX/Ygz4w0IewfqXNgBEOtiaS5e0kgqrs4Sv
tC2lJA3+b1aE+HHLEJX+d1/4P20YZ3uBjRZuaDygOtYC41NZF9+KL5yXu6nW
6UqEZCepkKSYoaSRS7jgqMMbSrStKNwiBFUHYkEdno/Icq+W7HrWDQm7QoDO
oXnZK7hjk6n1Ye2ZjyfTRxceaT6bBKBqobAIV7S+oRYkFwChfC+WQz4Mmqg/
NStqWX0WscGnkSc+vqRUQ0aRrhwKoK4Vu1feO5c4DkFmvIVbsA4EFhVBUvFp
eQjMjELzjMZQPoghtzqB1keqVb9Pj7y1OBBk5PaXPw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZUECj9J5y90OtzkMtB6ZcTec7hp9pSR36jgoW8mz1wU0iDnqfYaWajNvHP2V
umITc0FKkWVmsXgonoMfMtZgrcvKFSzFAeumPqIexqewAQGT7EIlEDeFwSVb
2i/6nLLI2io4mB5g82GL4xx0bJke1ZGN92VI6HBfN4A8/G/LSo4NsBEFctxe
lHBtUYDIUo+LbK2/lr5YmDzM1DNcPTIiz6gJv/BLsZmW1/SLjEo3Pqlj54rA
3aoW4xOIrKijFOiGMpHI+kfBUWGJCg+rRu7/BSgEpxNrTPQX34yQF7Q54Vg6
1n3pMy0fpVHqLsPZSP4Fq5arU50C6Llx25d3hpCxLg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ODJu8XXvjWM47ph1nWSLMeNUn8kCnzD7Ptd8vSsmn7VQS7ER25csn26WgyUY
CFkdGTprfOjyBsLYQpqfODDw5Ussbr0RdCdkrmdhITTc/RlYh5vclbljhdzf
MgZkOrxXMQoL78att2M1rczMRvObJhnt7C/XK7F+3LjUB3GTXE+1ppv9nlg7
hy6Nk4uSmLcqYaQhYQM7IMYjqjGIUwS0IiNpzVh/jnh4Aw3Dc2C9g00y2qI1
cmnV68qB0g7mPr8/Uqotl8vPvbuGn+seAtFd4A52o5I6OVc/++kFqHJx+lfq
5PEI+uQHU7sn/qbyoGSax+Tb1M2C5Pc6KgpGsTXb4A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
s+xMkn4iLp5y+AGv144y3JJ682b/sgDDXXrU1ajdFc2xogRzZ+k+8lGQTtvN
s/rX6VEMwdvmWdTaGeSLs4kfWzpN+9B2bLVuOULW+eq4pvY1DtPJxZMCF/TS
x+GQGvjuipQEls4dWfg5VvR7sUQ8Cb7C0nzCa7ZfMzjhZxeSeIY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LPOxwUIA4L70tNAEZ66az9x5hmJtLJB3txex+IqTW2kWWNc/WCtE74KY4HeI
IhGRSa4iakrf+Ng6qwE4pQwZx0Zsfauo83vnk44o/KQcPPA1IzntMMms71Eh
XbuJLp4TEb07bLkrE403F4Pb5VE8WcqrPNipx9UAdojhi8zewmtkkwGzwlfl
o2poKin9AeaHPqwEBsGBYejW9CDKOYuhZsWZyCEG9g4R8Mmq1/SmUTH6oGET
BjF1C84x5yrlls48j9QHhBdSZxumamWx3W9KCLwTb/BqSREQw+LH1uO+SbHI
1PMFd1VG8mBPnawpOyZYAwm9JvEZA3lBpnQDJ9wCQ+L6+gz1zqeZQAufbWxD
rfw2nS0XxzWWnz+ZyHIyjcJBefzCMJEdlOLRw+9xiJOlWHtkPcdp87lQipEG
tpP3duqrSVf2RVwYB8+HZahy7pZOsGsJQ8xypKSqtRXhIGsQBcHjyC7g74u0
umCpIfzvEv+Bc56UntyVqhM+O0x5NBCi


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BwXPMgGZX+iT9CfQpxJ7hAR7p1j+lFng6Hh/sTSpN7DKM8OJGWECNvDiRBVU
E+hUrL6UicL/8iK6ImmYZYYR6/voZ3q+wzzWsMJZJWKSIoqPI7ZS4HNM2F/c
tSnwbi5Dfz0UttISZy7cRMNOQsjby3zF4W9uOMxeBljOw6gIJwk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BiIBoEaEYUUInhToadmjhBIo3NqfeOhGNrNWugxp62eQIYzn2XgaOT0reAN5
tOG4mprIcpjnf0Pbng8ZbREN/yhcztzTCKxuzYyDtGNO8cmU8SFxtwTdAHRc
xNtLwP/u+07SwtMdzjO4pDKI0V51eTfi4aXxKapCojn5KgF65c8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3904)
`pragma protect data_block
k1HQnMRVhiosYH02fy6VW6OVzC3BhX/v2a/8wxHPu3XqQGwZZpaIHdYn9nat
mX+dWoEYUAKv++oEcKOOZgVIloFfQ3qmF9NSKkO/kB7dRZgDKubhvcbKLA+1
9FKW6uWjrHOq38ln7rKTyZZccHTgk1zPqU5jNczGSDfY6cvXioViObEWAnCA
91vj4erR2nSg33GFl0+uWN8NIvBumAhALnnkjnrj8eZoCXFpUMo1I+1+X2af
OwqqonApAXMydzJ0da4jkUVcfTMR2aGUB7i3i7YJDlIw0Hyb0rMrXaqStNSD
hIMIT1WY05ZdaU5A4+/9QmrLhY5JwBsRCn1mTbpLPBLn32GF0bfPYTpyziLr
XTe5eDJojee0eszJgJ7yYttOi5oOUxLsohBbxDbAVahzbj1yKtTijqnV/OxM
euXIFGTFTikbeRVRcDaNUL0P4yuMH6EqnfDz3h+8I4REYiwRNHmlxUDqfUp/
6mUZdKKxso0wOyRDQfP3A9Bj/qTcUsHUWRWSivmnHiKEti//PoyC1s4CrT9r
bI/qRkuqekVeH/fx6rX8JX7pkh8y7g43Kq63WSatxUzuCef5RyhAOyv28o6g
Z7k3HBjNkLmsr//IyOJihO2kDYJZaQv2xe5MYGfCwQC1msGLOg1yy/2C6ALf
H8X8FFSU8EpuR2ITz7oNaToUTR/2i+jAjFYSJa2TsullpMo/U25moMwIfEpi
+oeJWLIyuEJQA77+Y7QimtU6TipzZqh7geSQH0ZLqi5f5cBkXce8NRi07D15
ybaMhIrBCvP6VznSQ2JTveif3HwBq5zxex/+SSx5oaFJdUs5fDKdckQEM0Fc
EkqROwUiRbcHo3BKC9UzwZ4d/ifA2z6pPJSA6yfWaPDJrx3Uwo6W3DFulEdW
oSdlri7FxiiMNtj9+N46WZhwoyCGNTJIYNp5h5Q0BvzzKNXCX6czveVgtXBv
RvZY4PRx+H8GrLgnhweHmekvQkD8p5WD5qvCTcpeFfFeneZlISBcfsh8NVk+
sgeuY4AJJpuxvwZ2QkCGxwCbugWu5+f311FXqyWaDjaiOaOs7k5Tuqth0xW/
qwLQWvy5Bo43WDPSMwdF5PxHEdrNgi2ixYJhZnSN8k9kP7e+kWrwhFvL+NVN
9F4Le+bwLXgOQlm4p0PYaou3sOYC+8bHaUo6bZwI0vlixcAfXRJgi4Yj1fZZ
axTmKjmAYGmtg/xORQ1jVv6zzHMTZzRu7WiA+ht/iUgcIa8mKtTT2ruv6swI
ew9W53n+6kzMLk1izwYLQ+BlAuoTGg5nozP2bl+gogT8A80jbpHh3qlqZRBp
ZXDYT/kWrZYlEk4xC5xB2N1lLf+zOaF75ZsucFh6ndg1zN2/m0Glfsyqnl3v
vSEyScNV7LgRS/vekJ5jCTSkj43B7gjql6lYSmyMXPzccbcb/LNXpV1/27+4
JPC7WB42wE3GQDPeE6uaXzarWJsV/t/BizE6acoxXVX82CGq6vvMPnWKHWRP
sxbShBxdluM3fE+a+kCa4kUjK2ZBo0VmDtrcvbxn/xKn9QsOmSRJDYLFQ2wW
LRDF3b11x/Bzmo9sp+Mfwb4+gz787YVFywaPWLyGVLNb8keyiDcCG3k8cVpO
9C0RChOsfu7d1zd0Y1WfCdZ/S/6pLxDypkHGAgIhuObdtUndr5zzF8O6FsGz
gVSFyy3ohEtVr34bKClkzBw6yq9ZZdaa3cGGQSqW0MhDvbcT3ttSWD/VMnlb
Z2uDDlBeo6/m8MQ2SizjUQRxo755fNMLmXSkJ1FQek7qYxbvcN1PbsNNUDqN
YuxKkxXtYjT8r7eDGaeTno7mltRT/8OrDhx7BMmYW1ckFPRZ+jWPgDrlLugG
d/FPMHHgsrr+SMZ6zcB1t9/KE2I4i9ohV8JneHpyLk4Ny9ILQl+gN+RPP/6R
h1ZSlIy1e2b5CPruFami4TleFiHVzJKA7XTCwLP2jb4nRtl8LUWvlwyQ6jWN
Xi57Jt0p59gJo2bVHzt1S6ZSTr4Ql4nNqDwW+D/G3iRQQN201sh8RsW5rNDB
7AtW3+HTGVVmO8aSVRXPOQgXXKq9aUjlhwqasAZqapVlG3smKaAkkX2RuydS
JiZftjL4sYxSvNHdlwPo8uSHd57F/E/WjrCwLOukBe7D+Xfc+LtUo5/UaLEZ
GwYYWOO5lhxk/WRCmsf1S0bWKlLnhYug1P02TzeXodGXgwJMthBMdesbux6A
07fIIdV4YhgoszhrBSrbA3da15VxGUr9I1KLZbtKP+OmtYb6gQniZ++mjC7n
MsLzp0cUBfitw1Lw5tZZQHKNcDUkwuku/sgaX7anCjKc8yGIhLzdfkD4pvUP
5CK++Q0+Ecb9zdtfJ73GRM9zaECWjOL1ZJOc8meSeyTZ513VNgFhcmo/ff+c
NnnGp4ZZe3kzlUEpm6hAZUPVH6mDJaN4lSf1cd6cqyaMaZbr8o++JH+20Y1g
1Z82c5X2fz5NWiXH0HC3ndngSZlHxrym2RYacyiCDBhNm95eCl0AA5DVtI7R
IBZbsNFqTXGtV165XH5jxQUTop2UchrqmvhPPvuMz9DTD8wkQH4vyMJqfRwm
atUTpJnHX2DJvDuXzPgqNZJiXZB1h2x6OKwwr6s2DQ4RcU1n07Vc7DOTUDUJ
9zWcdTZbdpdVeugkgvn7QndcrekpMCJ7jnEubCFr6uwOENTal4QYP63FwYbY
1liVHshMk5JLkmfUa24GJpPAfMFIzv8ghi0BAkXqB6+O+8coRbykGo7VjqeC
smT5f9amw5kFAOsaQJoJDYTXJxKef9MweYeqe9m5jApC5ucnW2uzAsbLAIcF
Czd6jBPxFUM/vCikHoiJg3tiISXK1lKLEsAqMv2fhRe2+LYvbDjpIbbRN0T2
miomDHdYDNrxrDUp16T26o9TpCucsjYVtp0DQcHGTviPl+Xwu6PBaqGftwzF
CMzKCva13lcFXUxRQ5myDId5mNgO75wf3k/U7bCC2sQiQFgWVdTf40UiXVHI
E82/lsKL+sjNvQc1ui7KONLdVZe0m/x75WGQJpoiFUmUyNRbxqr/0mKySSnJ
S11SD2W4VdLByUZ7M5FzbNnxzJZYRgrB/A2TCzVfo87PbxyOHUFY4OmI2Jcq
tKA6ojhlTJYI0edux+yY6nbW08/FNpVsltP+478vHTKE/6vH+lENsIQddpgD
zoFJgVN2N9NbuRTYM98/1D2Y0cy7fRIRj8E3t5eUx9+sfYxudGwlvjtxuuAm
mfnpPfOW5T1zlYyftJpnK/iEUtbb7zmz3nAoltetVOj7fd6XkYEP0lN5xX2y
lx+2eeTF/UPgfwfz2dte4tQdg4sPgBvcxObCG08oveAAYYqpHkkXJpckqdrn
sofCenTGWa4iGeWP1MkSO8Jkf71jGtdrbeMwtib0Ds2nWw4bdAHcy2n4eFIU
OMMq2Qvd22Dgi7d0Rdoib7cJ8Ig6of+SYdas3smZfTtf7dh2g3dFICHJ+d5P
ImiwzW+x9Gylstd4nDqtumg2790zrk2pAbiZTn0iU8fmWPSTEXCiUyYQKG3f
DCpz9+94wWLptA6B5YSMb49MMzZ/ov0kGFqAQM64B2vLZ5x0UEe2RA8itW8l
0UmWNy3HIKeIJhUfX5dPFQeaT0mctTaEkap3VihMA5GbheZGPYB6E+qG2EoD
Q0nYu+3FiKKitOs64zpmI0pw6VvuPLsrp+ysilqQPbA3LWHSDiY/5Vpf7DE3
x5PZVbS/GbXPno1WD+TxxWRw2PGo56qF1vprtBsAqcqutEwrqRaugI2Dkz40
n7nJH/YX+NeGhaXsgvdKy9pdsaOp1sOeqXhwl+U75lGhPiLHH1En/I4NuRM4
MSp1hw4EFmlQmtu8rPU7s8hE7l4JpCIQ8EnKXQM3IOhpHRE/HoL9DAPXOwjf
H7RVdS+TCOeRoEJsDwkYgRSmanbGknvD3k8nKsyr4txIE1mx0CabH7vVImR2
kKOcUylFMShe6WuNOzZ5rVPd56/DHAX3F2hfByYXMFRM+L1YaWw13b99zWgv
qecGKPt9TW0ZbpnKUXP4ViZS1QLuBeWtnpcBJSGy4mK0pXkKsCkIlXlwBCuE
lSbyptFPGVLI1kR5/DaTe+L58BpDRibg57bFULq8SbSJ7NYd9QZpZ739yUTi
MnUGgi1Ufq04F5TlFfQo4sRW2EiAPRQbXhk4y5iOJY74+i3FD2WqnL9a42Sr
HD7lPeFE8EzcFnpZ4mo7H4+KcLd2Ir+6jzJJVNbwUPssK5CatmSnvwPiiOr9
dMW7p/0FTXbptkSF35URoNHTNcmyWRZ0wzjR1/oZrlVqVky8/ROEDJi69sUs
gfQ1lsi3NPiz3TlMA2WWukSE5a4aU1w/D9JzFN8i//Y/VOHDYTGp0ElrWCyR
OVib1RMi19eApphZqvACepZzxcPX3viszmm5+LI6JX6dP3upJfQAIHTav8zL
1qCeOeDafmarC2UhKRRR2zMNozqsfIdNtTjmSYyZ2uSE5X7MPIij8JNSo78P
eXqZt/7RXdyHCL04Yz6ZRHSGhULfhSjItlApa+XHoPiHCwJVCojJqObT4nBZ
To0FNQ4nA6cpnlau2HPIjyWOA3iRc1gMt3fJrawmS3MKrUTkoSnmoYz1NeF2
wkC0hDmOULKaioiYsMShNBpe99ReBuuDRQut9Z+Rea9duesH/4kQyokyHZKA
klpg9Bx+L6pIvrkyXeRh0bcPSeDB65zB5mVcM4DbTknA+a6LR5HKloFiaUTk
BfNl9VAWFwTzrJVFiUk5QBYPe8JFybmEXCTjr7hjas6h7fDQV/6qTYDmyzWG
NnXnEJX1cHUy3OyUhExfNBmJMOaOEFIGVHjgc6Ek8DZsKjbRyLRLBRXBjMmO
XHDECW0qjxAuw6oqSFw8H3leM+5h/HTpT+aeh7U0qDIncqUr/t7FMVobXdJi
Xv4Mgxih1KXHEx1inCmwtR2Tsxq9vGgHPvgYon3G+P0HR55dnrjJyrWE7HR0
T4misv6a6QgxSRhit86LkH2ZiweTRM7V+mcvYuRxVNJtGxT4nzr/xIFyQFJ+
qHeRxxFlvCHsorSjER4NjxoU8Ng0F7YR8YiPNXU25B4HZS/LIFOUsMjenWUl
LoG53/w73te3dAq58jWxXIwgrAWU5OiQW5c8TGDauNdzkUbYCnULnwgMG/EV
Tdchp0WhA8T4OAY9q1HT6QPDJlR5xjOAv/6W8lylas/lzg==

`pragma protect end_protected
