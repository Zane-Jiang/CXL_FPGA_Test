// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
nhM5H+ksDqNGKQcEaL41YTwuP0adOZKdZuOxTcxUaLAOAXfCCfXvtKQB0OOHCMtO
jpFX0tcgFw6Ius4LsXbTaPI6w/7iMHJt3XaZFHeXNI1w03AE2E1xrP9uAVyXDHdi
X7nBQlNleSiCPw4YA5KS5oJznmHXUFxjxs7+q4V10xCvfkakz1YI3w==
//pragma protect end_key_block
//pragma protect digest_block
nC2B6A63Lze/7VavhQ99hJto7AU=
//pragma protect end_digest_block
//pragma protect data_block
nzROx1jMYRLlCytAxvhvSFiEVrkjgfBcnQTuTWpjUjfN3y7f4OxM/PrpPcyhQd0Q
nszLkAr1ZlZV1J5Grb0ibUGD0US8gLiiRmgSVWG8hf+Xj6Nk6xuUWaJJEFV0zLON
BYWHW1/4vN/h4LBxqnDSqqIj2uttpI2rz+hI6dOr7DAQlAe2W3nNNXzF94wEXgNx
Xg+lRz6agH+WWrzdyUf0in5WeYEXLjQSOdVTn2KdqEe1ib/bHdVWki1k+Rnm0cEW
tHGpQgAQ5jEepVpzCrAvyeJXzxL+OFGagwlxs7N75TlZdQWUBFpPx8O8HB4fve2a
W3oVgTOKcbHjHHMYZTnCmYwv8dQzcWmF7XBmlWg928ZMxz6o1lleFoEPjh5/oFz5
xqX+UEToXkkBFHroLipNUiz7RN+VBFCtqswQMwOqWDjRqgDgI+376j0yvwK86x/q
kk36zJGPtkiApjf5S3EfFZnWkipKpORQa7bib28Xk0RUKyZ1JC/BWGVXKN1mdud7
inBR/+T8Gx2elmwyjUWx5wWfinh4QZ4CTb16ox8grKpXFUiheVbPuVEerU5Z8niU
Zi4MmRKNRyyC4weRpLEwNWIk9pWI+i16yy92eU2pWSFyMbE97vLZdvv3EXFHFk5d
rqEdth+Ffvpjz4KG9yaSSCf+GLCrfzIF9EScWVpug5eNJPziQDI30qSrPdNFS3fn
an2a9uU24mJ0psAdgK9bgc66H8ZbR5jXUSqV5LolDt+cxl+7GOdvbLTVkVRDnLM+
nsoia2+wHixI2wDqbFIYnzL/Qfe5xtt7OPJymHQ2y/o20jzD4K+N4sk6WiK3BIC1
lUI3nvlGTkbkYKy6K10v8TlzS7BznktdIhgFcuiM+SvrDvwyDyl2tfLIzbSmtCd3
NKf73KuYPRBxT6+7ZUM2tws8wESQgsOeBqijzYt8vkJQ/eZ+MP9Xwe/maO6Vq8BG
CDyD1EgLg9G6e4MNNmaU3Nv1+9GF7BLJGAju24r0CgmgzzmMik82Qh3dHVNEqzD2
v/43TFalJF9ECtrIKZJ7CCB2uwBHcumgm6m/Cbf0cMpI/mwaXvtaA9t/5adwhoaR
S0PhOpxhr0ioYmx2PurKhS63OZ+EoCpNC3E65vuyTylBl6rt072DPZIsYiEu2b+6
9y98mQ2OaXLProu1tISOgjLR/mnLKvKYxl6o3LjIbwpY49aqk1TpQjZIcoNim80V
LBp1pCD0RbhLWOp1w5up5KfAmsTq03OumbMJbMCgRHA8k6G6toX9X3ffFaFr2IH6
6a2buLS4EZF8nfowQMwgQpR9H+ZQGh6M325dm0ItTz738/1MIxulamAfG8sMRRpG
KSC5juILrFdgp8K6/VSUZ/TLCTIbOpUT63tZFoS045636FiOrAPOJorCBGTwJh4Q
MjtxRbvrI8MF9M3XiS1ERU/K+RqkxlsRyF8kwhIhaihZgPN5bQduidliMucsTPuS
nzjIpfIB/b0mGV4BVWFlscKmD3gRQBVU56uMHWTJ+Np/kOzTJPZ8VV2XWv/2eMe3
blSIP96hkqYXnjfqAtcclAcB+6VDwgLGcQmnLPLn2yG/xa7dFTS9ixtX9WCD77Ij
kaXPNEqJh0QjbBSVX1XWGrVdb1UmqS1bjLXzQUwpGvRXyHqzKEfHCy7QSl854tCk
yUoed3KCDfYSv7w9kbD/bDXQZQy88HcEaIOS8Dyl4QV+RI4j61DB0RMom+h1NXcU
5yG0CcV0vX5nvxLcFTzBoZthdI/jhGIqC2t9BL639acQQjssCUWBMsGVxQyW0m7D
AY97Bc1Q4DBe7GFAvO0RrKAi8TQFYyzGDlM3fv+g3+POiMP7doiqBB2DM+DJjbRS
B7g8jF8V2htNZC+wdth2GEq7kgEoVedH9MC78U8nKJ8KTsgp+bzuuuaEfBX25Qca
ki+e1h3L7TgGO7qHOBT6OdJSR05Bdvw8zZwtSFyetwL86JTyx7+dlkspYyKVg/AV
qHBFIBjVupqtjK84VRiYwptTOYlL6KBDxcKM0LUHdCU8ylQXiMTiyytm0I4xxb0P
ttLxd+p0hJ/vNchiOzUQNMwOSoPg9lbQI6qL4BZE2O3j4+ZWoF2N7+IHbUHPvKBa
cerlyeUG0hUKtUx8MtiGj8aXG5Dk7giGNnXbChJuQBww48VtIZc4N+G7aHI/YS7z
b2aaVpAI19GmSbsi7PmtGkM+I1643ESIDRGVvZGljUbw/Zrc00n9WTIOJfGuhXJc
ksrW8fGDSEND5H1UNhCsuhgvAXpX+t3nBhGxHW32NJ8vSIQBEFHOV43fPR4nAxQ9
PS+06BosWrv/Z9C/lz09kPo1yokvyZj7BhQEkhsdf+wueLWMWhiCd8r2HIIJ60Lu
VISktDSbwHoQfecQ191JJbY+SXtFKM4pXnUFiOiiaWXnZIUsUqEiw50M7IiyrC3o
Xlx8b2X7hnGnKwviDyOAYrrI/uGyGlzYxPjK8PT4TYk2wQYb/UUKhxG28VYcyIUP
XixqgXWOb+UywgdzkgzbrsKBQjZ9etg9MN5S0xnt3Gd/LQou8Fz9YUKOyGyuH1BH
QaDGPpRtMZ0TqFoQrvxxFVVrK6QP+FTPyMDrwEh6/YBIM0ulSSdd5AUxid6gvsPe
eDLs2coJXQGpMfpHoZI6rFgWcR9FmuHtsTLVNXnvuSmf4csDBjPhxm4pZ3+YBhx4
rT4aAcQAM+PO7gcMbIOEh1gJXaW4HpxR2MVS1aoUnq6n723RRXXSjWlazU6Lm5nt
2Rm1Ehmib580AjNxg73cR50ottAfbkfbXXTmbBfOlDfmoD8O3jDn/3TNuvzr0/vj
i9x/Ky+LzFPhNSJWZ8avhQua5kamjDAnebVl2nOZ/Q7+4iCZPLKu6mz1DjkzdYKT
vz5LIgQLns2ORYcmsgzIX+9FapwCEhheqy590CtF5MBflBnjsWk2n3sx6ciDcmP9
uCZIJGdKmZjSxmpDISPElvlRdUXRE/5BHY3xEjwAF4+J19SQ7lD4axeRI4NQiuOQ
2Ln4k3A+g15Vb1VR3SHFB8yUt02XTBy2xsizUZhEj6d4xO3kE4dPkEgZ72OI3qtl
P1yhevNBnj1q18tM+wyINj3h26D8PSc6pfnHvTealecEix3NEHyhVX/HM4C/qYMY
B6R/dfbpGuq+oPQbv/2YavK0lxNvrB6qcNfrq1EKSvxYTRPDwoF2Y9WUO0ug0bVk
j7KAxG55hpcVYcJCgcXcqXDkEhx4piQAjW4nENxzRNkGMh9VtA6ERuPiXRbyrYED
SfBrV0iRVMkzQ4lYdd/zq9Q++UUGBsk9yOSyCN+431rG9Jak2ZbuAkhXQ/QSvPYT
wz5mtVf8KW6IIOdmTJvUtDu0Um4MIDjeS4UjTQZKwg2QE9Yr379zM3m2CMKeA0L1
H1uvt9GjUw4hYAEi1P6PJLg5Ihrl+45YAY4dYZKRKlR2sgV83ZMrPbxK2ec9DySX
KcZQY6JJRZelr7Dr6O8s0dDNAeFHvA5jRWs+9Q4iTCjJPM+QlIB587TrpdP7skJT
CZHyc4FVt6m0ktcQIJXzleEK9yNzEqAlguKswwvLWQUbjvn6Tq2bWPdc2bNdRuzf
+GYOSXxDQEwJTJt0D5jf7AbQEkPOp9CnDfREMmFaxEUpg95sLJRVkZfJonBtj7AH
+pUXloLuTMXIauG37hg5ESFYJlthy51mB34Xo2eisTDW5yDCnUZqwIHodgXsMQ+d
HYM9tD/0JPf6LdZp11AGDJ6CNBKKKCAPbZNHrlW/YVdPfggT7Zi6sraSpxE/gnxb
3BiYxm7/ukZ13f7G4hh7XKbzVsor+raMkZm/wWO/nJWpU2HOE+yOenJ5sKOy9B/9
rBKZh4fqtGyTSAvhAHQJNkChP8v1hx+5vsna3LXsLEQ+IwnjMBEfcrd7xsvygzdS
i7n0l0rCexXDmSNJhDqkrGPVCnVBLos5PfikbsoFPIcdQbZn8ztooJlCPoS+q6WA
4zcGmvmcY7dHbxFStnhznW/1sQSS93jI7SXIzusHnGWqO94gDFuNwMJLNiQhkrZt
XlSpRqo9kNgKoX6LFSJPAIOpxxtujviDZk+yfV2iaIn+kcE0jXzAWP2pAwpsbhXz
bz2TfL/j2VP1r3oKgBQN1hJpXIqAUUZwNXsoIfkC2Aq85day3//S2QJS9PCcAYAT
FwiPqIxAQmuFS6cH6pkKQTtLn8FFNoGq6pN66iT8EgJcP0p+iLbd7/IoOzhWv0Ua
VPGM+2r9Mw2kvT9h0pS/wZpMzQN18sGobMVK0Wj0PpFawT+Ad8fU75AS4gauD4kK
q2aKMdLdHlRHl0ITLR0oMxLUggiJAYFDC1ukUQzuHahrWoRG8WwVttGbX3W4e744
YPs30lUalDXcq+lWh1+c6RRcV2PRsURmtt8G1Mqh5DXeyQZqhr7ZtVgJA1zekql+
5SH+S0tZ9gHKUJtQb0xm+yzC+g5B1JRqVcBTJ0CiTcqKU2W7mrbxjmnvIWr47PbD
hiN9ir5SfE+BRzosU2t5t8lwLXhUfN2llxdZECDOsJvLlFarOERkwR5X05aBoyS7
M30mMU8YUvZmBUax/yHGqi1IWwXK2pgPIztEq/nf673S/88crpCzwxWqj7XqIcTc
yNc4BHsuIeebFGUw5wAPlnZDjL+cice1gVSRknmuzOiabsyfmvlBdKOwT6vzezcU
yOdfxCaRDOKDIbNYJwVI+5lQGYEMr2t6nHHaOdyEIe9fNhafrZ4cMrUHAoTXvBDA
74m/jPxiUmx6I1kEX7OELjH9HCfCd0Y5W8z0G+hEHDFxtRS0eziY6cjmV5cXJ4Og
I4m8RG7kbN+Zj4ArGYx7mq40vXXPvUm80Cpl+guQk7ID/Kn1+JVCOqAojkC2unow
u5UmtDDhHhBggUiuqcWWlDGQp94KAE6/iv8Ie6Pi4JPfQPt6KJbYM0k5ELK9Euu/
hA5I7790wZnhFAvSzCP5LTwmx3Y+mLIf7mFZq5n22nPvPXiIFclOExOGojRj9hOz
CAeIJVPWdixRN7vrMUCwPnldFNEndsTtRI/ZK0xHI9y2+ocS+tAVLYlbztOUDVKz
y/JGM5PZ3bw4H6pO9HzwBGNs5vgKeoo0eZahxNzEITFmhsdS6wzqvfYjfXJFKbWq
0uVXgJIw4xdm8akx0rK2SYuYU8a5yB39BzclfBrFlzUoPCmjP8FUXKyIk0hGnrFi
KhRzWp6+D4JuP42fXnxpqWxLGbmQyu3OqBhslY7lzsFviGJykyZ/Mrbbahjd0Hgj
/ad1kYarcMc6jT1Cp1YT1nS0lrOxndeuWRA8vl/0pgp2f69Lin8RQ3Z9bPwJdyM4
njIX7UcCXFhyL4WGPs7PBj935xbeaSpNi4ScmeILDHUltHfv5O2nyDCPR1HMqO8B
f/FisrUBq1py1w+nAmp1fBfjT/rgrNlzDfdQdzY/U6QA6V9VLXidMwMhtLd3segJ
axR5hjXOB+ZEvpieOn1qL6bNbAEKT6iEtPfkPIcCASUcwkWo4rPeo0k2dxbNQlW2
XNe70F6McmrwmnMy9G6se8yOqfUgW+SKu8VF0G0bESgEdRHIaIt23es7sdoVq9ee
yptsIjYMY7r9FjtCMb3MlGvY2mp47GxzijG68KkcewZvBrRJ57hYSqhOqjnFeQOX
ET8gclkMxbcsI0XFVn34wEmTOO2daE7BUwxGHJaSzYTbI7JjQIg6pNJJvpB3maPZ
l0p/v2cIWrYrqXNU9COsFNsgMPJUzCL7htazN7kmAYNXbkat7YX2wA8fKfMPT5Ul
Zw++HGUqSLlWlTFdDEZxLYEeF2V05i/NqyQhLPOkOLopuS3Zf6xMSs6KHzpMgOS8
82sqTr5VJfZQJ6K0AMVLVxyiU5TpX3UfPOAeeYCIg0n5oaZ0oAqJ3x5UZQndVl1F
5VLomvCEp+7zON2n8SmNc4kgeKjFI1EIrRFOfvoUN90YKK7IMeq6Wqy0Le+MtqA4
JfSc25FsI0HZ3oGbqqkWbbK4t3T4LrxFPbQkV61SY5TRepURQNnRLDVcj925vU45
cC04Z9aWi01lLdozpwYcgi6wUMTARpG2/junJPk7bRHoZGYEFUrErjxreLLdrBpm
e3y99l56ECrbwuiEwV53tK0qjzaRtW4tfLQ8694gJahNkqrYldZAmBnGhq/E2Mx1
L9rp9mzPFchMherpf0zlak36JRy0uZu2s54eJaqxvMFncNFyxxGhkDVb2ffC3fNW
TBOKqsJyrKm7Wtpq6OxM1iEoBVCFZUjFHFgQoIcuPPQkj+1MyYoz3upe/Ifl4dF5
mbe477nr64GJU/QZseCd/kjV+k23mj3lHHzHkH2YGdT2pa5X5NNvNZYjuqHfLz1y
6HAUIHQntNZuYsvnkS+SLG23fcyQRJyKpNI/vpZNMFmneTJGJDmhte4JiKpg4UxK
lhouMHtylkf3BKFHyMDfdLd6PHEPxYazNLkstQSYptk=
//pragma protect end_data_block
//pragma protect digest_block
ysdMY61LuVJVuZSNGjspzM61vZI=
//pragma protect end_digest_block
//pragma protect end_protected
