// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
bxxgENql13PT4eGTMmfTqx5ATA4ZW0M8+EQYuxyPcRbCzrTrsr4DJ9I5LpYCYX4DGH/XpTUUJwYo
/FYKBFJbwpIuXpb8odXhowLShuYg9GbLIpK9G2cIPa+eqp2gc22AMcWEyqMAsJIDcCBuz0wDiAei
273KTo5yGi9Ud3CHduEd9Ya3OkG+pnpX7cpzT6Q6gpFjDDvlRlQQLdqdTwkrvgiwCkwKtSWqMv5z
508dqiuXLYvEe/3HQ+cq1Jqo4TgEChnJeUIm0NOZ2/2abvUVHN0FFOsNb0WNXlA7/0iiV1VQmpYO
ZH/zWc2v1MvBDfUJOVJE5xOeW2NVjYQf+d4Mqw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2272)
6nEMRG0+Lh8gQaf4JuURBXAOwcPl13xOmAN0QN4w7x0MUSVHaxGB2K/gSztYLVfMdjMJYCWVda8F
GfgjBSRQxzKnKNgiIQNe9VLiCNG49cGg5IkA29z2YYnJdJWbs8GX3VfEoiWq6HROjIKVOJwOXD6s
Bb0kVJzWpSelna4Vb21V4IpdFxj0tZLo5BewXPRKzKKmObNxG4L9fhh410Jh4OGMvJzCXhADNw25
vJ4Ct8nt/ctGV2fX7liw4GaF62USQJdl+pKI/zFlfU4qA4VT70V/b4G+MVFVHvZTGpxQM6fXOD/L
TUlPMOlCkU3p3bv1qUwBiugfOE5XTLK5eqClU5gt9uzPItghX6Hw2tAzZ55g6pQ9VCmXFdOEW7mm
EEZvJmRDvsld8pggKqUMiPIIWR8Gaohf8YMBlxibaPk4znQ4R42rH4q9BljGqfioH3btIfUg4z16
Y/BzzTo6q70CqiSacE8uhGuP9goI4JiGRZ3WXze6cTWSnAjq9hLPAa09IctN+ImlTiLnx6LIFBus
+7P1NqFI4NFSQpR0r1+tiUkbfa3YcuUaYjHqHD3xHysrwiEuw486ADbE1+dcaZZBk3RKlcwgottz
q3iN/E/O+nQD3jNiJ6F6H+Gbe/eCtRoI54YyolGFR9lN9P9ut/R8B54ovKcEgTD077THnQJEbQfW
gGbMDcH/Na4alOFPeeOlO97VYmgC4fkOBL1mztp5XnR58BMktuM36kkwn6hMS0VKZsm9av2rmM5h
PwziM37x2ZP4mFJl0jjpaX8o/r1dEXNyA3ZWVsqRvoLS8oxnfHTuiA4qWQM2VgaOp9IqplrYECKo
volS8NLOZx5FIM1ki4D6rkCdqhme1tRFnPAMUxBYsQaB23Tx4arRqYWKvf4yx2HKFNLA/s9zHwVz
IGbFP/lUpnYojCwGDZUhLO/miGV+ddYkEBylmcX7C016xUNmKjCa4l4hUaxCJkPlxDC79OtIFvjr
iE8QuazSilY6UkYye34rOLUtipdE0iSQ68jctpWQwLyzDlUVYEbiC7XQwInPTMbdzWgtkG/xC8H6
1HbT3BvPOE63NeMA5A/rrXQolKeiQxIuDOAu3wp/yiRKUHTYdiW53r9ehsMVWQNonJDUPgfU6k4g
X+Ifg/FMxqWI8NuTlebfsdgZbs3BanYBqDIENerP7wkvLeRc3bkqAf1G8UUP9xv8yWOKBLODdZBv
sENzKWZpIS2xOr48fYBijWwiEmK3IFzRQ1PvLAvyUa1aDSivmUJDwQlpy6B7P1rA5NxXXsVubIRd
h43oklUnRm7J/bNRdLdCcLICBx6pL9WqcZ0Jj8/T5r4hiY3slnKUGADqFYfcdJYHi9p12naoYkqN
YKyH73GZ8zOVnSV/qQOqj2EaiOYjJrcfdoB5DILMEPw/jS/uGKrARiAGdem1Nus0T9+ORIx4YQT7
3ScEg2vcFA5r/+DFBz9LRVIumWlQeiNCPOqHb8IMpQ6SsOPjD7yLeoDoH0QK0dmJHWq9tuQQeUWD
5oyHhSz/MFgXvnRJIzVpti6qpMH2hQMdaWb+3QvGprgGQmAPFli7nr0ImdcFlLZqVRYS+2zHxVi1
K0mGwwVlQE+FqLAR/eky4jR/BujUzVavhhHdOelp/G5yeahdeyvc5V/pt6sFs58qQFBkyywesNHg
DqGDM2ji+W5EgcAgOK2QKbYe7KeFWfQj6J1vosp4gTE7xouR813vu41XtNbomxtPpTRDSGT4V2BR
b+hskImaphqGiP4laMCy6lUHFAbnH4BcplHwZB8DK6mMUy0cf+7ACRm8XSq0JOeZq3MqN8DWz+Wu
i/fmiolINZRtysZXmOSTcW41XnAmeM+kxGCPTUSNRtEPH4A7m4zSqUaf0IzK5PjZqS4RjT5yRRwj
2AenRMPRqfKs0b1Bu2hGFqNM8E4VLJ/B5yBCcAmrz2XitoXHRxVUs4/Nx1Hcb6u3C6zbhEQNJJBU
4qLna3Z2MV9MjDdTAyDFKgVUMMZPa6WDCjkie/zpgeF8GuGiK/lF/0N2fWpGv1foDYbDUt4ZVh7z
V0NEB58dakLAYnaZm2mOhV/v7uNfhrcNyT+lCTLhk7EN799pHYA3sO9AqTm9nmRVSAft4pnbE5Jd
dBvto423P5avF9e+3lEWUYZvkRN2qHMr7AXFUtyqyVEzAESFX71BEQFcSQlsCWinb6hDaxQdpbi+
BsOf99gYEKECu8JEdz7lsgr2p5IwghNg5p38B3fEoMjzHoV5HuU+Iw/rK42eJqDesj7nF7Zc64U1
cBUfpdoF9yfnfgGKBL/KZG63JoH0t/Jouo/7N1Nf+wKhZyHxsS2raNdBh9f+Rs45/Lk4tcVPE1gS
54dcLSdwXGt8z+1sDyqMoUyh/tlR49+HBjixFmJTxbUKNxovmSaNcQ8FWb0wYzSScqdhqxOH586r
+cnb7WFDzG+x1+Wc2Q4VB5AmQR1tY53nlWU627tuRpPHYYze9NutVymp47q9DwVycoazmnHE+jb6
anXi/p0PU0Kk5ut2jcijmJmVVeVTZwmGlUtMFozrrpXInsEdlcyIoVv/nO/k1oaDBJwmWoy7KD9E
a5pxQmVnSVxgme8XnQEsu3VaDGhk6QxOq5K2odIXt5o8jPndcc86LRPCuzi+vRKQ8HZWcq0XB/Af
V0LWj1UFpJ0jLDioCaCCRfffPMgU3m2ZOUBylXmFNaghIvlu0VaHgsa9uEnkIojw0eQ3lxDWFjtF
FjS1Z0GS4s5F1qoN3LmL4LKvpdtfcQProq7vn5drMqXYA75Ob/bB4PWYoaPqTSN/0w5zo3VZEdDS
pkLIDciclRYYPyhQshvUnOaKa5u9W/UZGOx+6L+0Fy2W+mcMOwo9iMl6JoOrFNGz0rh/XkYUVJD/
NsyolI5cFtK7L+HbTJ0gRDdg7tRkkxFI21TOhleX3KHGdiDQ8FPFInxBDcE7dXgUnZfKsVBROr0/
Iumkm1cWAuK/smKCrUfc/3TAXlp2ABaXA0czDgKVkghU8O5fA8qIpzDroeFev7I/9A==
`pragma protect end_protected
