// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
VxnHs2ppsjSwltshvvRPFNlDD2o3E7bw4wVtqa9hMEDZTc7dup+P1Q2JiCeWHB8BXaT3T/asgbnJ
zFrXRG1qwTYmjIsaQAm40brB2/qhbHEbUwwjvj+l/ZPrBPLPhWxnbyHvbBAk/G8Z55nNghFGw4Wt
eL8FRziTkgSz5Xh25sfcvz3hEoz859Es45Ks+U/m1xjW/LJnW4bx8FPCHzsi1gWtqig0opxwB61/
QpciQwPEPfZSmKWKZS5fVKcmPX5H8q6ptKMQ8kTeteQ8aR7gqD5NsA7crBePBUxrX40gM/ghslGD
JRBPswgVTUdokHekfF4BK+vqNvPM/KK+kh8GyA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10336)
6FVdkj0sqxoznp/XpcmeS7OgRQvAEMTkVN5VNVn5xeimi6ad8GoI+PuFQR6Z2tl63IG1laq8t6oh
Er+wgXpdCBaJ20yAHR+cJOPj9XNFOCIBjgi1fK1SPvqAvnpYTOLKu+7gjxtteXFlECPVjYdAblyF
WxRagax6XQ/kxofok492ACWrjLCVcKkhLldn03nw4G7uLtl9spms+k85jm+jB74ntkVHjLpP/B3g
AICdRIrsd+Zqdo1caCwUJDovsXD16cxoGyYY1oXYcCQGE41kb8lTFmdr4w+NmqwnHO3N/SiuGkUC
4gmV145/wmTau0r4ik4poBkCTV5lVJ+8QeaofDqn4LcaSBQN0BVWz9h7s35nThL2bH4Qln0X/aJZ
TUOAW5ZM/HsQoTF3Rtq8zn8zPf1WT41iQ1DcGOB75XiXZSlz3p3NWxo1Rsb6BB7yYeTU4fVKmXm2
o6Rjwf8B75rM4F8nXOXPziPN5TSvourKwUzMU6VX9Jy1IeOV/fIrwBuw3PSRY42byCUp/PM+TpXu
Z9vRwa8+V8v4H55xCRRQCGI70z64ZtbX4uLftwpRgdFkB343A/tZdcAlR7vqYyvL0D7CFLwXNwRd
KxSRx+ZjdgkpZf94xx83nXe+fOFWkQVK9IR4eMx4y/3KQ2y6KYjo8brG9m0Wse7ysyzR7pRheeqd
uyJZ4movqIadRKAXi9hEpH2jATvx0dnG7NsbNrHNP7QNMDDUfhP/P8c0cCDCcTOMgwqaYewlQtVw
xl+X+bRTWQR5DR/QsyspoNphwoyD94GFg2jf4qdTiLYFheQ3yO7SqjfFi5WR4hbFxaYJBYySQhqb
XzNiesP8uqn4hnBM3AcUxIcXf3yCVAdl4632oKANR8i4DSyPX4Gsl3NEVrWSoGtQshnaTEParAsq
2RmIgyRhrIUpzObrAGiPlvlVG8JoPRzB/jsikaqskZrT2DUmqkuhfFxkXhYJ213OlgutsrCdRO2k
Jx902mT49xbc2jhZCFAF5qxGRfnlhG+030GPdewnEbs8nhwTa083VjdO9T7CQ+5M1vXB7HjT6wTw
hwcJM7rLujTAhpetSG3kTYDEJveowCkBB0r+kEnOo9G7O/39iXZxSNrbERBlSDfeiZuVD/A3ylfz
nuIl2Ba7sIIpQP2aTwgRK/MzIb7DQRYAAfrM4KzPbi8u/aTbWOMKZArh6pEroLAP6Cn5GkE7RjhL
ucNSpHGGsxl31p0tQ+Gi8muLhvICfm+vvnvmx77zXx46lmls5mP0+B9eQIxjyvEeO0D3K5196dDT
lM9ou4932e9j6mxAJexxdYC9rEBS7tzc+3VvMMhgkHNfnRTuWhWXon89GN0yZ3hNnOdOObRBxpU7
DQzBoJMRBmk7aWM8DEMbpLG78RbNaq7bGVJmitdn61KHwgfY50eYBE9MSFaY/foDcT9oMJsbjMhs
hfVLFESLJqumNh835dDBEVR1yCPyJ/LQdmggyZ50Y3E1QevVYmEYKjmY6slTgJJntqRV3VlBSrJL
FxQTnXx27k0BUmMVRKkYwsUJmuR/Lqhvyq0v5KpsxV+5GsAXjxMeD6tE/lqHp6TTEYs481wxTD+k
wmFwpzUOBAMDXe2pov7hvisgwNjf05MOfUvuVaQu/U7e5dwx2UVaUFiZ0jPaPlmE61kdKlihVP9l
GtIsTJB9LkN7uHagNuMp0gq5XNvh0VnrsmndVrMDQ3Kcru53M7KlxwP3rJWKlktGC73qL0zCwh+g
Cz7w9hwG1m2OKbclR6puF6Ydcg70GmEtPobnWQYm7cG+E4ZXHkJv11pp48bm9RO6OtJ5mvJpmw7Q
YCRQSrvXLODDKWQjE7GNHkNMn7S0CAPX3SkhbNBUc7RZQffsYXRxpmAMu2EFhV7wKnvvVA5DxwHQ
itMfIzSJewo6Nq5R3yNxNpNfpA3+wZpgR7yrHXlBunox8lcYtQpL+2SWGFOSifJODZEr7chf9eea
SaEGFn8Mb3UpgTbgNGtONKVI9UK2NNqUvAbSDIvnXpaKGhMVxgl3Mge4KK03cqwk8dT9lsIkEPzW
XwWwFmsY0fwwgf9qyfPdJAlQPUtr6qznGN1qD6U5Yh+kRlkoOPBjtQEuy4Yy/ZzDLgXMg5cMDFrf
YRkpm5nkbJeh7E3biCZQ4Gt3HZ2pnSOfy4TVb29h57+oGWNe0vjtEkprl3s3IZzfYvGk6EOet4CM
8hvMy9ApaQFnGYCQeA19w0Czbgamm3iXaMeHUHponOz/B9sdUmIgbJw7PyLuowUVkTyUt1fRFIqZ
DC3H3VqBfotLs2D/p/yXnPEuEV9WezsXGcGK7Sx3rGZcQkGGW6JWoec41lZa0tYqY9Wy9CXs/QsJ
2Z5FaNVIWdeiML6Sf+x8BMJXZAu8AOKcEYEEvzz5C9XaOjbSzahDWLCqeys8sDd/8glwQonWpiq2
44XqD6o4Ed4C9Jl8/EyQpNJVdiE4YD33C40u/DwXzSm+x7qAT6xqcYUY5KPaxNolkK/Ax8Vyt9O6
+I1yyi1CkV2rNS+zCSsKWQKiJP2PddC5F4G88KExhHsL8NAXswYvyBM41z6JJhK8MAbf8WyWb75H
TIOKj1r1hmwGWhxTIwla5bwr1E5VuEKpNjqRhbPQlpB6WbppT6IC4t/oMBGr39vQVEz++0sW1l1W
n8kJNDgL03C5m+qHR/MGYIbL9clgrE3gtYlr1AIaVEVlNo9sWLykS+0tcyUTp4EMJufzZHOJbciN
IahGcBsufIMvSBoAflAyIWYtsqyMvaYvpLg5IdVoeeqkIK3BbsGwbO1/CNWMaCNDnYQegQmPpERI
OpSVNtCsCwpJzcSDZqToe2WUPetfdaq4BTFaxp/lE8H86RL5Avh2zTNh9th5iD4XE0VR35kYFBZi
Z6SEAXnmfKdF1Bw6ZH+vz+9+rSchnknuh0Ro0ZfJ4Ox0qkUbdxagbgPizbPPKXy63G+OVCi12bFu
W0YvEG5MMYQbUsTOKf3jtdnKtcPJHbpX7Lev5nRS3wRL4tkalUvFCc5rv6SV2bWdgZZvidibLN77
8JAZ9Zrxkl/Gdut1NGw84tOCYaQuex9IxVroAZnqrS1XuSoUQ40cVx3MVFZc659WkWRuNjW91Usv
BgV/OKOA2ixOgxszT33iZHjmA59rCl4mOjdWG9DEoSibvEX0dQyH9GrpYsEOl4D7ZyNTRBa796Tn
4hO/2O50nLxZDW/t+Z2qZq2gml9KIsH7usQERu4GPh0ybz99nzpXTcAQ/eZ3Nqo7B9dJpnz9e8mp
j58ApA6LfOuSssSpey5w0GfR8xkQ1+e8KBA3ZJmsb9FZcAkH3zwz7+j3mXN5VhtrV44gb5bleZKj
pFuENvpFb30R7vbHCgB25QLBDnhzLKC1t63FLuLN1foekcQf0vxGrh5EYX7KL2imxkrqoPGpurq+
YPVZDRpVpXRmLN5VpJI1gcED3D17wItzLgeDbrpVH+BeF3M9k02Li+MPg8AzmRttI/+stLDSrREn
hojc1VTliqsGES3pMFPv3+30hLP2GhoyfcVgVa2orKP2gYLJ68uAGBiekQzEh5u4WPeLeKxYmcjw
Ig/QMskuclKSleJW5cCLrKdsXi3mX2vboD7aoxP2zxW41pV8mYNvcDqOR73i3+31OWe1FomQnHDD
xODM3oDg0a13C3QbtpSWqRSEAB9LCYUetag15f2TixrtFQFSPhN4CGocb97jwghbRd6D6hojqG3U
BGBtaiNoUDmvCgiVaKr6NnJAFS5cc2Jg/u+f2pjPz+QJY3Ba7B6TXda57sZrHzaTQQe8T2RiyAEQ
3TOaj7wp0eELmMIXytE0AzpSigyBsqu4Urh6l63vNVo6ckGgAsdF13JyqKV8rl+t6CjwPsTRHUq3
VLolDWPrxq4Bwcc7q6QVTi6+3urMC4t8UIfe+WkVg6WbsZrq5ycer/0Zs7GF2Cfht2/Kth7G+nvx
j7enND+Wi7qjRj8J9U7QS3H7MWZDgspPFvtFMBXgzNEmlj3K7HcxcXt2lb1t/dJEV+9HWHXT4poA
TcgKI51Eo4zHxDffr2r06MDu13TtvuAW+hSZhxxSlxuLyDYKcJmvHrnnPrWKl/EIb5A4EV3dX0eg
QB2bVbc6/Vc37DH+kkYIJOeDK+7oX2K0XTvJh0zRS6ktrJjmGGXETkwFiACMAcqw7Q6aCLRp+yNo
MkBurDKeY4R3/KyA7zbsFupVA9s5ldI/JAQS+vGYRnb+o47vr2nGIj6OnjRCrALTO1HFlG/oPAhc
QLOiOBeH6sVWUtIg8XCV6mXIqfDexZY0elPkKofTj3M0bytHwixlKj6CZTtIsqQ/D6GyKchAp8sT
p1+8S/lMQbFUxIPOfb/rSIlr4nHSkW9A8+VjFwu3W5gY1CC7h777+tS32lrbyKczb964kmCocvPO
Jc60CtXFY08ds+EweuaMwNVFB0IdrhB+SwbxJD71S9+8qXJh8+sIT6dXNav769Ng/UjqkDArdSnc
DLQ0lLhzLLXXCHCk48aIPcfvOy+mT9ByYF6S6SIedsi3PnwpbpJ49GtB61PGyP1JW+5TnzznaMyg
OpzOmAlAs/EH7ZSnE1hi68h9B4hVQHrmj1Nu7tmzhiYox94UWUg1nfvA/29bqkevbqk/heDbHj2V
RSW2zOf60A/B9BTu+f1CJio54Uw5JS8RVM2wSts92GWjCLUTO5EB67ai4OIlzPgpZ6vLF3Friqa8
NfvVnrqMLzD+OHnsUjrTIgAA94QOCjiyKTbhHdrUcoJC4GflK+ACo0uGd4eT9Z70crs1qhKe7oNs
slahi5Tn/Xj8JkJ85wvYjBw5nvWtX/G0jDMx47BKDqKlhxI2q6AZNHDL6vRDSu9HLGcHeu6f73Zl
ms3EDBrIqt7VWP8yJNoDavHma4t7Xp1j2u04HWbz8EXoClPBNeWuwYvQD2tFkV8QuyV9ACf1MKmd
P4duhAjnwrHUlMnBGRTHARYlr+jmcq4S0f05+i7yXe17Q8prxRX3EoHqsDFxy9OCQGXUONrXq6av
iEuqur8bi4tCDRf+QcV/zTOZQR18anmvaZETaefDxLV2frVc3Fgkd8T9DBIjCD/zNcTfNLTWKZ3C
sAMx2ufKW2rMUa21oFQXi1He5YaJ6tabzj4Twi3nhiM6MU7FN12vsKc17Bwh+iJGDzgT6jF9Nbpy
lwPvND1BQqtWJcDjTeULxCiuZbPo/51r/rfmPa2MTwBW4JA+bqvF/U50pWtJ5T3Bpm2dZO7EcYmn
lkTkH38GNghpio7vGQKHdw9WPppcWeR+6OSPP2Sksseye5bx7996mu50rTvgNcvKECf68DuVCPJA
c5fUyLfQKNrYEV+Ze+zNSG58hcb44pHS2CUREqj4TsEaVJE2Afba9PpbnJEXCj0EznR5mNUwiUey
C2Qkw8r9YKavDwlFQH8IvYq2IUoOmzRD85i43zaPzZ+N3ZoKPMsuEM+0dyu4ATf/r06+GKni/Kif
BdenFhfyyhZTjqpfhDlrv/h/PbNVjnSzFauXA8awt19fdnbQh1EFmfwFVHnTeedj3ipmLXtRp68t
l61MznB5W/V8IioipBcjdm9BC+b7qTMnG46Js44vsNWUcyOPstFW0SwfjdlYSgpAG9htng714bu8
uONPqYrcMxtn1mJIuUZFjNk5nsnHtPmummG3LLyuLX7UUBFuh6WaqsBALrpQotxNQ0Cx5z+fHpiG
xYmgBinGmoeRn7jhoPxDJ11aNabqo8lowx1dot3glUC/mMQ77hGav7HPcSyEOSRe6di8YuWg/iNf
QmzbjcDMBQvtCIWRSRnCjXEiS+BkOqDpDpfjN2MjeDQSHldM7Tpdee2StdbpwyySS1l2gqKSvmYL
z3JS61qJqNDB7GnJKeHxEh8JsL4DHLdmNTHsXswG5keRgkz6Stvn9w1e2gDvxetOQ7Ip4tsorhge
bF6cUV2TPdNRmWlB34CFWzam2nQK/4tNMO/1/NSL0jER2Y5nXBUhH7PM+aT0ROktJhOTRnCkPIhU
iaeR/aHVkI2zI4KFmHBi8+hz0tXgjPfMTRXAQ3rHkHnKc/jd2kZevE9FzmH13iSaXf5DytO5I5MN
KbvPJD/n3vnJowU1fuybYP9AGvfSq7q6PA/rsNlSR6yJCNfq6kh/Y+t29669gTrMb7sMiz+sySIM
H1sIlurYtLr0qBpMfrHD/5xUU5lEpaYQobdLK2IZEh1unKK37H/nbhf8JCO8sYN63w9AOAOide30
nwLDlZQwCli5ZcrvoaabuCX7+aYwC1wPC7/jlmzq5/6ZUlWgFQlfASbtUyl5YqQHZyFpAHpix3Sg
RasPFGHM3qSb6jBkvsDCNJfCjouTZABAYyjHL6rZ0uzbOHqYrpDQFr9gtWoftvyEpwAg6lDh6YLi
1bpZt8Di4pEQxQqA3RTBFHowKMA8jVQCRVe93OfNywR+pVdX2SMZF12T0+vvSRePzw3Zrv1M2/RR
tP4n0Uc+VD+vjeMYPNgTZOqsBV0IDI6eWLVG4QAEgBukxhRrgEswjDMzvzTFLSYCE+NF7rX0f5sy
gOhUpm8ULGfaluBorJU0WuV53KeE61iuLQsH8wtYAkDB9KDfuCL6e34WHaQGZJ6cWYLPQmFedXgu
btr+lrWddrguFP1R+xKf/OP69kmVqQUsUgGRnd0npexBzcmQcjVtb31PyTlyZwDzv2+ruUrzr+Ml
LGd0/eHjTwoowcEBIjOarOjpNmllANO8QTesSOuTOkOJa3VZpXkfRWl+rBVD3oPP2hL3T2gCJ4Xb
k+Wcr2evEyw0EuA98tKZkd5Sngz5Zqw5V3Gpd3YRS9X4GRmLkHRYslKvYG5OQKsxQer2uVDGCqa/
ohGgxFcHLx9Tlvlgb9zvo/W+RcdNyAuEFumaliX2RBr55f8Okh5/TBuER9RWLiKTmdj6O9fW1dR+
mcGLqH/RoGhrXiiAaxQyeU43eCYe8/uL3ZM7q0WfsLLTJsRz+pzvhDpWTplopZeuksV2KpU34EiJ
SDGr65yD8rsdqnW4ckKNq2dOVxP/E69vXKpWzt4gFVitm9DeDYaAA/d6DsNBAk7VYV8Nz4ObKGul
RYL/emsjZo9JrXSiRJNEKMdz3T8/YvpHPdVCmP7O40RdS3EE3U1qnjPveFDJl7HyW1CAY5E3I7GG
NkZ7+9ZYqw0Qe/Ui5S2AjGR4jsIIkAmYSdqcsgX1zfu/CG+LV9g4D1tlPhsP2I07+x59UWe490Oc
j5zMfDFSKITVsPdPNnB7avaGuWQ0S9TE7hdr7OJa8+dhaCb9eWxCjmwojz+xcUo4NOKy4wIcQAg9
sc5hnJcLMX/t1DNb6IR4fSp/fntT/sqdak8LLND+NhR27c58oNyYHvRA2bTLyvYtTYLpCb4RoX+3
pgpG6pTX7/4Dj9cLgvAlpqBxSCcYXKG9ha0GjiI3vK+F3/5lcv2Gu4ZbTM1Si1p/W4QmYleXOYSy
FJ0Vxd03YvTn94utaWSUpqncVfZEMzd10FAt+yXwYyKjRHvIeZXBq4d+4B0jdc/oVyIB3Pbw7Pjh
TDmLyndy9zITIxLoNNY0hvZopLVS5m5rDNDDbNz6IRYVviXgwoUl8NOTA5v8qBpfZwC91rl8kH5L
djQ73BkX9G1Wf/ZrM7ABvTy7lXPygD8C9R9E4vZvDnCLaSSp6WOHO1lTahGFwVAnEZJ9jzpBErS0
KM+cKYyLK8g6PHP3LpHsqcLA5vCBswjK9tL6ipsn/SOf7SR3SrSSy+TSyubFDkINPlPrm7oAGzO1
Pc6mCnUXQyBdNV97GOKEBpxTdszXReOrxwUH1jdINazQeuy8w0MVmSOcqQC8syBYrIDWT0xXeEyh
w7K/Qb6YXmUn75Y2UvNlSDGcG84/8LOu3umo7lw1StoBG4sqGLU+J42wTdtb33zj1awjlew9ocuD
1l6fCGxKLHh0afJhFKxX0KX8PBLmaroZ/MhFlP2vHEaEx3ryMSkCD41KDtnIWnUsoT/ylRoleGFu
6SDQ135Dqt0lwTNVgRG/meifPNm6C82N+xyk1aAnqoGNi0DZEiGfejHz+yrR8uBQ3CH3eoxZovrI
NTjhKY/4jYWe3bJ/UFYONJeUVfnuC0Zp/QbtknRIjQew7aWd/zpmvlSyQidYcn90+kgiw6HzPrlV
iqeHVRjHCrdH2fgXBYWPWMlJXXy+C0erx79G88Bmzm8B5Wc4w6cfteEnq49AxXly60i3gUK+uk5C
WNFYvFSB6/0ZlKA8ncq7q4fEF4Uh2nUoXmuMfCF7m/K9Tf5WJcoM9LU+8bYxpGxe8xBbYRvH6eFu
OqZ6HS4lpOFflyz98gH58JATqIwWqLq/9IJ0iCIc0cGad/EkvKTQTEKqTkDFUJfJ6VJR5x/bJsVI
r068YDuiKH7r5bBMtVFaFBC+DL/EEKK7QGxg/cfKKMbrXv70Zly3dAcZM3d8R2UL53teB2iGPEP8
MnLilqNf4cLstsoBo95yI0QHIeww6ezDnv9yIEAKl8sg0GfrEKhJOzsscQLFCFfxVZ4SdsTIx/8m
QtmpCL77OQT4/7GDaaAafBBiPr1udOnH8tjIet9U36mts/gkK4y48JofRqYwPPNc4PBYvWEUDaUy
G6AUQdBznV0hwx3WvoukQJ8pg1vH9g24TgsbsYFiua3RKf9mdQNLB0G1d0tpd8W6FzwKejwLg2JN
0MLvy9Atg9TLzYA2wcaT0Y5SSjEqu/N7TNh1xXJS3+6I/kflnlmfBbMXwSYfkqePNXHIXzMKEwq4
4SgS2ol7qLxvaUPzCOmDV1cbw45jxhOCTnQ3thnkSml/bK2nfySEtIBC+FrOf74W/4h4d9mysS7T
rcIUiBj8StmIX087Rv0OIodus/LgdQK4blGHbEYdw5JXJTOWeeZyGnboszPWZJZ1YbhaqLHQF6YA
+oBY0MyAtvr/GDCe6IY2N/eubEeW231lj2urX2upiGfIPX5Ei2Xw4Ianc17BsgVSTZEGWuYQq2Z9
JzEuxvc240va/CcrCK6rZrxSz7081VV+HuJ6VgVBdaS7xjvAVc0K27WOdYIVbUBesf3buahiUnWR
gXecrcnLbiQcwRMU3PMF8oDXgkM0TB54Y4lK/q91qjQOb68kmTG3xM6dWF+0ccPcOCsa3TpUS2ZV
d3F0i0bG+Mw1aOTT9yAUBOqTtWtNZwcVP+UAT3Z+dKaeMOTw4BSIlofftwk0ExKK9jyHOK9As7Ro
rjfqA0AB2KY0MCN+8B/i0WiBL7h6u/iS+mkLwdFhEjRx/U9AEVimZw28DpOf4pkhwL/uOx7Q3K7O
j8h7Fd80DQRiHtMJ8oTUdSf1kdDdph1GTHpua91un22q9f1iJh/FMTrJsN8sxXtnFDBLo2Kxcj49
Wy86qEWfzODvsn6577CUbpfRY4FeYaWuQjrkvOEXmhqpvFPdlTV7knFe+TTfxyEdwEZncw/RsV6b
pkuzZc9WYXUb77CW/Afoi/RxIMUVXL6t4OBoCZlPdv8hQKaX86Mybe3lvKCasMeyitCDWcT3Gh7J
d9dHzyL1lpT7T6RUOx/BSGQZgOTxs3X8l9wbZ9oHyB/o/KJ/F40Ty9wTdk54dt1Pn//QuYlzkYGn
Igh20+YD6zfpPIP8rPBZkBZbwNZeJnPZk4mdVuHdlZlukpeI7QUFqWOUlWyw1j0BX9kpyiL2yXSl
BBmxXcdsRD0PtwT1Hb4SDxcfLl35noV264xTiuoXsvFilOnArCcRW7FPsBRFndzHogZLAYeIfplv
4WkcZf6Phz6mEFAm4pLo/n+a06Lm5iHmb9yVGyfSX46XRbjyv2m/tMa2mUIUnbHLi5cJkjRDAx+9
6NDwEehXJyval2kurQQW0koEcO5ykzLeNg3aNMStmBGnEkYquDeqIS3qc550FKqSORSVvP9DrN7O
1O2fKz1cIxpWJSl7ROkdxIs80hinaImjCAZFv6esLKyRL1efnL7XA/Lxln172LNL9CAHMXxyt0yU
tvSVT0s6YoZOeHhXNeWT7T/SZ81S8NwyB+M6wXE8kxrWEFke+SJuRo+IgKm6Na826HHCg4azcHfW
8J470c2E+/m6Ms9Q+2PfN3LCspP9cNg+SSny/nHZi6eZu3BQMnIKy7izh3BOHsk2pguNm8OPlZtq
pimt0ktQGjFeEBxt0Hv3iOTEm579xZqyv4lAM2Jq8YhHc1d/y/3/L/FZbtoF3F4bVS3tp6lApozv
WVVdbgKDyouAL2zb/22K7ztyLEYh97jvMEWhDIjPZFY7kn10Opi7pFUHZ9jpqDO0OSzJXwH2qK3g
B7N/drZlUDu/qWdZW0AiSvpICE6LKxDP6NIXeh7CSjdtttR5Aeh44d/JOftdxXpPATIsmjHkaZd+
i93RL/KCtgPmqU2Y5gk9pGf0orSkgv4H8MKFLCUj0jyfXX/pwIzHHMyERNu6BvjqAeHur4lt5yho
BGcinbU5bYLCCusfoIEIhHopQPjGas9ZFdIfqBQtXz+DtmKFyM23IXHMg89+5p5qO5DL9edh1qWs
+xASDQYVmCCLx6+rqtlA7D1FlrDBOO0qPGLT5r4+RnnV0FXZlKGOMNfUBIi5L1CnM7XidgdBlrk+
rxODSLUgcrRjvlIq2gTdIalhLV7OlpU79uQEHXGcC+DyP0YoLBdCYzg5bUH87LkNJiGxhV68vOKM
uwgvs+kTkMyunpbPcdtwXNn51izuKxaG3Jy0JuIuh3eeaOPtREcoAwc0MxW0HDaZ09Qufw9MZsZW
ZDoTyxCvgeMN5sC8XrlA2xpks78h/FCaC4eIoJNCiwZbODnqUMvySWlD9VCVMIL91xmUhVdYqDf+
fJZHEHwUXgZV1jxXUZoDaRs3812x3uJjvL67GwxzXERSfjus5tUbvZzD9HT8D42+2x8QVuTVupPi
Uy09je8V9e29OVBPE9eaVsNQwzQAGOK2vFwtiYMZcSghdGoL9i5FbjRbv3VXlQofkH/2ga5DfP9P
iM7poIfERc0fVO0XZTj3782rJ7F7Xo2FXjXr09FrZnnlyyzQTutlkpZjrz42keqpo3oq4ogiaZZn
WbDJ+LVwomkVx+Avm+jzXRVItNKi+OXI3OgCyfPMlzIdghJ+lwCW0qFfmzCY4EpUwpEs6ytAe6ny
GdwNpQGbbgpldutyHlsLjtsv05cfZsj+RSOJw7mfe9+rmkW/u1YB78HLBcG438tCtK8jWxK4g/6i
AXwssFHAjhHv55bf5+9+OrDuRMFoLplU4Kq7uVKU0ZlG48ZfaW/A88gTttX58KsX1EeT7hnkA84U
jMhWlh1TB4Hwfv2Ovop9eJvUxk+1B9GPbozYt9MbgbyTz2frkK9HjLCnbxc6pU8nxSOC065xPlub
l9tkp8pFvH+OKuOlqpn05jdsuQOjy3O81OXb/cWP41hUsaIsqfSfhN/Zn/SsANRfW1sBWqAjXZ/x
yBHFcVJ5DdI0a5haBLjUIp5dKO1/dU+kPay44XUfw7Ea0iumY9Hni4K4Y2mMllG1idJ6rahxyhRk
3XqnD28sgPKyboWIwjn10+ElM4FoI6QCSlhvlwqwxFMX/8YMCsLkcycAzV8Wa5TejvSZLYVCb9VA
b5mRI8j2ybbYVj6DauiBpRvyUOD6M1Gb7l3/Yw7DWDdmyixSArfIWhi2rflO5BKxIh4OUjcnRHk5
NAcRBRrwXVZa0olUU0Qxs39v5jzzRaNGC/FvnTa3WhHOzoKvf6xCLnb36wTa+IZVELSTZ1iIuRHZ
VwJ9RUsce1lxVZM2eOBJsvvvi1f+cKazb3vX6UFiYiKRMAtvmNrk9h5b+Q9Pi0MfpWKDOZHWtPRv
k47lJoX57Agv8fFPqyRk7wXePw42NAggBfPIH9jk2GI3r6Rf3aTN4DCbX8hVo1JQI/FBAssQYmuE
LTvDYtVCb04uGOEUNExErNH3/pa/j5YtGfK+HF3RuZ4hslF9LZT4/bbJy8tmRquytbGlIl/wLzD/
eENc4VA1T7Wumb9b6iOCHG6S2B+nqyLF2CCYzbJrbSf9bkeRYlROrLq+0LaN7gmlVgDIhbgAQuGJ
Wf6Pwpe/+vEDzbQuJpD0wY1NPq+zij38BhvymheantAixBAMljrmgg9SJC7SVjNFaVl2uO+AMkja
881Jwqde0x/j7Gob7Nw40Dd+6h5EPfrvUza500Smsj060iYtWaKxSaaqIEAbNgsfn9ynKqBRP8dI
QfNakoFsfJO7vGPlqlxrQqBbNo7Tw0Cy6DDrRzlVvWRlSvczXpI9r4JQYlrv/p6OXM/nX0jMhC2U
v6Y4co/nS+4f2cljD3f9xBl6dohvROiVLDGOWrZ0UkaaPuCdhtGUtIEW021usc88xvuOp8WX6k67
XFW6/gId2hZtvGtOdRAqOO23M979ybpj3esCZwxVOs8n0NHVCJvgI0jsERNrcTz9gw3oyclYgGpF
Xs6OwxkWVcniX2sSJ9ZKJcL6A5gB+0u67dWRXWxXX0/z+1979PPdOaVb35LEW8cRCqBEgP3cPe/6
fjye2Vdj8nOU145SKCIbmUo2CjHt597PPw0gvA7mlegfg9XuFH6fwYrazW3DU183QCcFG0K74cgI
zXOMWBy1zAA4bS6n5qfLzhdF1FrfmBDwkbBOnRy1lWzxUEGHBKa+Hb8qV4EwmT9y3rNi7Von0Jss
MD4DIIgY1vx5OW6NUrc+4w7U9XuUYxDwQEhblkbkx/gsVmVEgRktBehP+M1lbvD31Ad5PdFhmSFY
CduAG4kU4Wh0CDRHLQzIX0v+8lvkPEBmznxVvWiRKVStGY40I+5o9rv6DfSBKPU/FfGhaTt2pJIF
GyMxN9d03MM3PkbWPCY+dmwojW0KZfL1N8V2rql0emwjJ7CzPUTnGDBnv0Ez3CaHAkc+wPrbHsYW
b0CCyTiNEN+PbGWntzrIwZQXroxUcXwBANV6ynxLmCTFyhR0URCxh+V3bRMjXo+BXaVw+7EAFWTY
TK9FMpCqf+jaCAXN+fRMVvg3AUK+PJbzCKm9hiFZ02LjjDx+mfJVGtzNG89r8dQTv5Jez7q8taLR
Juz3HedxNijFW6ptPaZ6TtqMCFF0Dyk1uw9jx2wvgnGass8gFjDxYIlP7atEs5PbfwvyNro27GuJ
nEZXQ5pYeNANyUdgz/RihtHV3VI0vWCXDrDge63ddBRSxtTdTW+DQgoJfbEAUyFNIAm3uY78IbsN
nKkp4WhmAVdHgIGjhctBawVWmA8c+gTjLCEU7ZGUuqcq0YRc5wgEO+GuiVDIvEU38NFd9GlfVyzH
nWROl8DU5lRyBLNj9uFwC0DbkNQZfAeIXTqLet+s9kOSx+Im73jUIZvNLFU6ybQP83Qe4vrPuQ2c
QdccbgUlLjQiIw/7A00lFtlq6VgZ6P51cPHkfs8V/F3QgallsE24sX60SDPkrpiapJQTqoAoFMt/
DibLIJV/O98pnFU34x6JnQ1nTIzf4WGlgU+koXAXurKWwLFdwP+RV0kFaakZV5mX7Vse9FZ62zhO
0S2hS+88HJpkq3N5ymX5zxH67yO9TLC/UCvNVWVNTAnjFg17i4ZuxVF3ap4Xr9KA6zmHmiHK0n3z
7cYYYh9CB/c27wSPxLtsyTf+k1YdZlxwkmNN5i/996CTpsfx43EOkbbJ+unoMcINmmduYg2f1s3a
aZvdireOQooKR2Q79pgjaDsBIj45RY2XydxYa8aFimmhrdE5gO8Rwqd1gQVDyTtKX2t/WIccnlL0
bfkfKgvn4Zfc4GlHTgjmuRSyLL6ehsi33JWicpiMPUhkJxKdvWh3zObTGv15RjxPWKsk4ioc34il
s1n4Kx5YXhpEAyJN3hRNRHPEZg==
`pragma protect end_protected
