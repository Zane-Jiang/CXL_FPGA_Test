// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
F17KXvL2y0FbLddTqrxjAy7gawV0QL1A3aCnnrs4T3xhBVSO6wd+XZL2qVat
k6eGnBK2+BST/gRFvJ2Ne8fqMV0ETL2ouHxl99u2e6JGzcI8OCwhstVVXiaE
WKpPWsCp56ucDmzhsNm0hAhmdey1whMQ7CKsTuxp0h44rTu/YCOQwQYbYmca
d87FAkXGSh6vEfKiMrlCWXwpgJAlrLILx6nxVI2Vr/z0S5OGI1UThtqnANhl
ZleMJ1G62E7C7S/raoFjjqjeo02JVxqm2mqypEdOVhNiIDqMSIe8aArFriWK
pznF5YsrIK1TSYYMsSmjN6RxxBm3iE1DTAUPYiDVNw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o0QmMvyMZvzRftBtj7Mh/l4/UfrbDPWJfTo5MW+zOSxNyOlqsOZmJaF0yVrz
rwxS/m1zXaJjsjExNRN2WcJiUJln22odrPGv9f3JfB0zObyqWv0yQms0K8a8
/h87n7qQ6zNfv8w7N8+iF13yTnTnQl8YY2uRZuVWYIkW9A+FXwBCnMwb5Aih
+tnqFIBxxhSUjoSYQNWnHJOjy7Of0VC1QYVF+qU0Ubkcbcg3oYTdxrvomGlt
ez2yNcqGrAPvlWW1jVGUq0IB3H8UVH4bxvijRi/fDIzMkCw31LdwPv4zyqSr
1rtNhhUDTevFqFdiFKnE1Hon/7FH1JtSDRRqfya8OQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZTjMqzJ4Z57mW6Go+cxigoHh1WFEYNT+MrhkWiuuANnPQzG3Bis435WQs+tr
I0dCxYb8pMF3321NQjI8fGz69QodF8M/4eWMqa0jwwkgvVoNF8RqGBovF7/w
wQ1iohp2yv+60u6xD2avRkbWLeB80AOt96LKhdkNRc5ZhFg6dspjZyWqQOGb
DWcXOM/1E5My7kWaUw5/1fnLj9twlnSdNVyXhz2ZRoC/x6cATZN2KCayE0dQ
xCFTOxilC5i/5o3CKt4V2KDAFjiVYX0n8GbMVcTk3c4VE4qVGkYSAjMdBB9a
qqPr2ihiA6ixY/cabeh2rs4FNeOvo+bL4fzuxUCBKg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eSUjwxCv1L01ZpSrWjIRSa6uSZrP+RR7+bWIZAI1u8Ke+YdyIhrlnk50oLmZ
XodOudmEexuZpljlPqzuBkYL6tkaui8tJM4DIAuNvkDihVgctf9XYjoXoYm9
gs3Rt01GGXQz6TDqESwgLnl/ZnsmbcQBReyjgY8VDONZF+ieJuo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PnmbTfon+6oOa1vFgoEOXxMekiDD1gqGw82AMTDoczbpaXJV8QMFPvNMjKrl
I8/zDG3X7hgfiZ83esj2+0CCWhj8e46cRyP5Vs7JGcDyd/4evhgoPixEEphy
O/p86S2zSttdx7yTh4JxRAroX+L2LBb/fQcY1Xk9y9zX4MoZlTs+5yesQGZY
xuWJTG6pvt2hwxyXRu8YK+qE/3hbQZ6+i74jmlApQJWTPW9p/cp5s4vjB3dI
eggo2NIcu4R6JkwHSPjIteml1T2Mu3u6FG9NJcFV4cBGSIMJSnmsuCKh97OY
D7PRkR7YbRDWcvQ+txpZZFg9tEgLWYHpJXI086afw0cPtyxOtmLsbNP7LjIH
n2HGVRbQav22o/RNAR5MYo9DhzFtephdxlyyU70UbASUAvSnTbTJ2EuYqDT4
acntHkEYuQYeLeYxumY9zt6C+pAWllwi7wLIdIyCOxG1xHQ7M2orDG5nOcW4
GzriT67vRLXnqm2KXl7ndUk/zW8Q349R


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j5ElzSjLKmGXMlI+DHp/BIkxKmaSLLeBjGqoDz5KEiQR57I2l+2i3n2VSg5d
tAfiDDOnOpaQhs5CLxzJL0ySEZaitv3aEr+fx/y5L9IF5I0dwyz4qOOMb9un
FuVpR1FP/wAm/88iaY4lT2Util5q/c4CxFqGN6i8vYflrW45Vjs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AFWlTPPYJMfQcPOC6v9LEXCB+AwKTSya8qSX8g1NCb0s37nCPAGetS63t+Ve
YK6VQXMzPMPizT9571spk2/DKg6e7pOxnvK2iaiUwKpEkmIYvy3qSxhbI63y
3VXjP066iP/Aov3g6LrleSo1PDfGYQbVHxgkT+OhXK7cfyw7PbE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 76368)
`pragma protect data_block
mWk1Z4KtJ5vQIKutHYpEqvNmT8FSahNT214V0wuwV00TbYwW35x55YMLywYZ
UeHi5qFEGk5A5ScYQhIFRgAVfOYU+Y725gD0OUSWXcjKFyva+DL5T4541ytg
Y6EsI9K9U5lH5lJu3M87NN9ManBLpPgxKPNhOFX2sOlnLdf6+kuf5m4oMC14
KgcSkPAUZjhfE7sRmiis6GqJ8zW5nZHjgDLWsSbrNSv16kiCos9Wjfofnctn
cQyJYMDS+IVpbgsraLz7M+/2MrTxZ57wt85nfITvlVGyu5oOcSZJYFRsOuTl
JctLWEeniuGGc0Im4FZpqRacrflmU09HtAh0d8EoSVcFQrkTbNkEbFIPiaqH
nbuIuWUblVpyACTu1sHZBXkBQKWuEwvte9v5QC8/SxaZYR5Yi3ONEmyAJd3W
NYN4M9dfl4RHU6ZQBT24M3xw0PKz7LNHAgTgSVAcSOYA94noqkafTwiPfqe3
vSjaRJcxSxZmJFrER4bsxhXKLDMf2+06QSWXQqgFGYaanlqyd/IYTmDKpxwi
59DI1BLp2AEGd3bamU8YWF7YZk7YXVq8ayzJad3GkjgkTyb3AkU/JJTIy5YT
PX3xPX1SKHntIZVdzAdSY76EsrSju4HrtBGMzeMEBg0WMgpIvxR4Bk20EL2o
p3CcRHP8ZF5yXyypPXcqyxk67jmuBNKKbcB4nm2MflLrJ3VRAURXZWpLizJa
OjNCzyVetQPiibnw8whUbWrdBYYWCIvfJ21m4LDWb2hyybK3dhp7564DcMa9
GenoI2mZfzPzbI0FwOSO9O7qPD9IJLuBU7S4Pplr+z1FebVKT4EC/5Zc1S8R
ctbUkQMhu0D5nkSwINwJL0ii3QyPeXjxJtT5hnplgOTZobJBjL9KRJHsvM2w
DV7bGFHlVvj2iu6CMtUaXtcf25A67WKNsL6sHwC2qY8xlg7E2rKS3aCnsvOc
NJpscmi/nq2zZVSGUbNzyYphF4Xzycm6MPQPHFGR/nLlFKanYS8ilsTIcOTx
m02lb5y2xb5V+UHg9t6B1YNg2UawMyt8miYrtLnjv29GtHCaRRm9AV8dnGaa
P2WG2SwqwClBNq8XWfpk2s3ABnTIBRmOGnsvYu8OcQO08mi/73TAituVj1Tt
ye41T7FKeskr3IrXnCi4Vdys5VqIMxJvL8IKo7zFXfuxwLcxGkFHJYW+OsFy
l2UDtME67Xq53OoPx+SD9eQWRud70PXNpdoM1Xn2jzubkeFqaEEEGSv8bI6I
uSgCZsPeXeFJ7Aa7kXH+4x9COPjMUNCYlvscJLw2uW4Muy97Dm9ZhD4wXqVG
qmUK4u6TWVrWLET+T8L1zvsvH8qs3fBcuQ54035Q2Yl0B+lx1ZPRuQddSw4c
bUyfm109kMrJF49burT7+IvcqPtPi2MFl34cPa+bBnadf+525q/sQuX40XWJ
Qg5wH6b7htWyWx0r2cIQcHDJwSMTA2/TfuyJ3BPSWx4r7fXStedWX4X/5AT2
xOCdwh90+Rwi8d5/0B0M/doiNemZGpvOC8CCVB5WGYNQSNOEA3SBPWZsxIGh
htBseiCc+yzicyoVgpwbopb8pMvMcvdmWtlIfi7mlb3HUUpTvQtq3J+O/XgI
R1NlhvwSUedoerfqG7/Z9IfbTIyEaDSRnykLrDmx8PM+EGAHqFOI4TWBANCi
A8MloZOlC5rJTLg1rCk/7K+INoO0WYeBlwJxk1AxKqIWEdJ5ZbSoX+7JENiH
TewQedmKGk5v1ZiI7SPM2QY+OUbWe923LpnBLrswrbZg/VsgBX3KtgmPt/c4
BG9S+wKUbwLTCYxr1WsjlO9q6R2GGm25LHfBBQk/2tGTuyrqZJ9lzmNDGTcx
9gexc7tmM/uZ1cAYcW0qW/ERXtUhcOQ7Ic9MMUsz6aDluny0SpzSHvHrkpO7
yDVMJIAybhP3CabsjHsBhayRKhZqNz30O149xVwWvHL/yGRb0KpIps9VeAXA
nZ6B+g9N/4x10Ymn0J2W1NmDoiwc7YzppPxR+6re3HfZBQhU1+eseZBEK45G
diQUZYrFK+ANrFI1bei5pOUEjtE4zZezxpxbfWvtF6Ch4H6YEYx0i7kmKt8Q
s5svJ+8Idc3D0JjmhKWvMjuXb0WdKnFvvuPXYJ1T7HJgpKrxDxsNske29D8V
9HkqmDnhg7lRU8wK/VYz4TttFVcrytZOVUpVP6voyPSKr4FOhuoObwVLsxvd
3baxim3BG15elKj3T7APpiDpk+1SZkOgpt2WIEbQlQdvlJqkOIhsewpzFIqX
m/Pe5rKXDX+TGLmk7ZeVTUQEEbcWav0bE5npAURwFStC/r8qtA8GQUAnQleG
OO+VR/kSbmPwn7P16QAv7sonaHVCAzyN2T/CrHhATQSIPf7eM9oBZTDIgMal
eaiDWh/YT8kxcqwB3U9EF+ZrAJadmWYJsRnKTvF9wstRjxStm7+mlthUVjYu
9T8qtX7Kn9rI59z9JPX1rydCHTy9OzzTQGpJ01ouv95jhddWAex4GLeBO7Cw
NgUxpmQ7yDBnldtvmAsODB1z84JptCfzh4aTAU9Mp+iFBrw3exFVUnlCCdTs
pVbrWYz/P9GpF1eXwi+4ds6Pog8M01LJTJsE4xZGtCewuzFm0QDWRLX4VEYn
PDSESn1r+ecP/iVG60yfwsqHhd21T53UhzYhHC5FhZA8gu99zUOMmc4WyJrs
+WqCbV1L+tBT2qe2srV6p5YA9vGzPv+yRYUpq+cHq6z8uC9KWuDQvQora0C+
CZ95+Ia7tmMOlj92NsDV21Ji32BB9uf5bCJssiQuv77MK6CJaFZSL3bCqT0X
0iaiSvw/79+D3AmdZVd09Q2iO28dgWtzdenkFn6oiPPWrKotBDOn1SFtLYOR
1hZQ7UBPhN/VPlTMuG8/YkInLXvOTLovBdFCpPS1CAXiyUYCk0ZTOo3zPYqA
BP8ldGyfoITrrJ/B/pscjN0DRgda0nvyf/hDrzMGknd6IxtXuL9MWlUMdWCC
YLK6fSqS73NaLrk1VDoHtb7qKGbjiI2XQcQ+8pK/VOArn8NEL7fEeXJZ7qRk
QYXdIAA2qexTXfX+IEBb0VnZUat/7M6oPeVvkwPi05D24UwpSfBlqr9XNmJW
uuSMHDh9fKT3TrsbahxfQYVSYoIg+wJsbIfArf4qKSYj5x2nWWai21WVzhTT
qWaE7GUdd/WKd3Bf/CrHgfnjsGZhoUT4DneJxFhIyGWY5aNxN5J7fY6Ds+Yh
osVyzG24XcnZUb9hsUlxwjRSKlDlKpI21MO6GiXnB7LIEEUoAj7wpzysVhaQ
tC6Xr72BvqCsTDw/pD+jYU6wvgY11ryxR+O+E0mHubOQXRcT4HTIM5lZbBGe
XOEN8dZWiHlHUR7S+QdHOeMSEcuYaFTNNNsJ3dQDxqI5TNicN9u7FC+rxooy
KoMryLK5MQWMwAuQ4rPQYV5q3GsCKnw6Fh2ypaSDrn10d+I1ZsOwf0S1tCIv
mhRK/Eb3SoDfisPRjVRkeTALW4eRSVt8e81mxrcvrKOqJyUow3GG4uiWAFgb
OKKNjHE5ERQbOn3CGV054+vckOLeEAf8/5I2Q5NnxNua3whsD3ReOD72YMST
LE5SzF/0/vQX+l6l6Q9g/scZ3Ue1xmv0425cATWluB+As7eM/oJ03keVvQLk
AlFFDFTWOcQT1VSolh+T+hW0gg04DAmX5xN4wdZZIpEjBFN7KJAaGqq9hRZI
RS6fXeMxMAXoA7hkr6GtOwSoo1Ddr8dPxdQgcb6rfkePKWCPe9yi1U3a5IvQ
HlvsiTFbB0pg4hiAgB18HVgni0xpm9+5TEn5tWcUKl1DNPAKvHCQDlpzX+Lq
hJJycjTeG7PjIKFlu81wdwEWKpRUV38yTs3m+bNLDtGK6TrzOv4+KxdDsBr6
Czl2kPAGMBGfoaqA8k+VGY4Gqrt3iW+rOx9lbB90/Hwc6tGT+c86gaWQlOVX
vpNBp8SG4/5L/naZ02QCWUISi3OXLJ7/r2xqmfYXEfQQwQKdvTL5bXIegA0i
fR2WzgCSI2QmWRvd4TJBtSJumufvSLFc9E4xoGRCAt3VvtC8SLvwn9wOly8h
YIwIsHV4I0W503wkYJefGeAdQXWzSLkAukIqZo1LU5H1JR10kOi8gyBryAX8
zrXgwKO+bz1KaxSZI1RyAk9ImzKaRiEAJcBFcLdJqe8hhS1aU4MfXzhexIDe
+l5kmhtNwedqICfkN2F4te7I6rie3vBnoTX/dvKuKOq3koO7/DW/zEJt4ltM
ePlJ84Clnry0SPqsH8maXiYor7P1sGeX94z3nrvP5o0BQygJyOLUi8pAuNXa
RnIDEoa8M37VEf6k3GOEV98Bp3SiuEJBGLgHdYATXq7VTUUc1fX4XwMPx4xg
jpem3JJCx8ztHFoVI+nEhtYpkEHiaVwXlJCArmydu7t9q4/Ixq2Z978qiM5D
modJTGE4J9fdzvGOADaHlryJyGGJcILp98TFZcdHmcJCpApjb8ZIDcvptHZs
ksGvvIixR7N1Vz3ZUCn0JaL5dwrvyBDyTAL3VSXfOK/vRA0HzOJrEMwgFEuv
LUCOD8leYG2fpOpr6edYhSHHmGufPtn2TFZ9w8FhnIvY7LDssW32agkqrUwJ
n9NXk0xzEcfEMN3iDX+7uju+k6W0OKM8EpLS5ezBt6+zVsIUUr45boPN/+Ek
XWTXlHp3aiBkQ9qmpbHDycJyYwYbcuccTXSELWEkBFJ1hSApxR/jsguQXYLR
zbjxKRzKsUIeOPXZcnMBsbMlwQLQtdpCtWY8UxJVBFzeNFG0npxaQNxI4J7j
cz+ktsixFm11oP0jAJ3R1iS67hdcwfZNx7pinlrXNTIT7mZShTpS948e9D3T
0K0hu9F3G3zgrhbBeYoUjsyefixKQJY5TE1e0bYqyXAtAwtdkT6oMOCg8BIp
1irahgQrtu6GgZQugsmyYBtOdlU2HCL3ONDO93C7dG7WrTzUg8WIytVig4HY
/lN2OZxPIocV+7O9NZIgegSJm8mI8TX1ma7ATLlQ72mcTheE9R1W005siVU1
fV2cDG89jEYhrR8aOvkPWgYoJ/oz7mFP2ZS7D9aMibgi0tu4Wy3DtKW9L4zz
kUEDwxJe9lHWpDPOlBxmCoxAPjSDjpD0wKQP/SFuKHRij46PIVb6NQ2zArnP
oiR9FTHftlHLs9U9/uGlQMHlifPBd7GzumcaQ2XLDyxjUPtpHZdgslDKWu7R
YLbw3K/UBpqBAaZal0R9IlWVWc/e4RVkvKbETuAdd8HvynSSYf6KJqt5/0sL
Tn0/PA+6GyMpGdwY+lgZm72GtWGMg7L3sVloKieVKR6MUaTSiuEyNZulJ63u
T/tLLQYrQIwIYs7LQtlFV5P32UYLWiKesuNt3J3uvmV/DwzBj4i+yE9OBAp9
MDWYye9ocCjbeha/CWZwtVTCeWNJrmx6KTNX1BTGiN3qSW2IL8sSUoLRSX5v
iEmOTyTuqRWr9M4SJS5eLezL/EJLWVYfhtu/a6u76UluRgBlKRHQLxv0oC0n
mNb1snOpuHXqIX8KvOpQtBIe+KnGmUIqYWcUFlVCUOapTiJCBu9kHwY6wkz7
h2UCz9LFENwjKEldA1I0U8i8yf7Mt5qNAJDHwKV5rERFSyXJCP1hUJP9vZYX
JFqeKceEACavDFGSHvjVqUY4E5yLEUU7pf76nJCuYzJCtksACP3B98R/PE+1
9YgJNZDXHXTBEvIWpOGkmog34Jcfzj/zL61QyhCrud0XL6LOPSdbcglB1mtX
PvVTDawFPknRiYm3L1Bf7jBdYYiF9LvWQqGdkkkIVp4Uo9JQZGaV+oxU9LAX
nOQ4+2pkvjetQWDl4+G8uINzI4+gvfb8frYs6dZ9W59N8pcK0Hoe3rbpPdGo
nKE4F3YrRVW/BHnPqR0LG7v6S04hoypguhC5cXvWGzerhZFtUeya5PZJv2k3
AXApR4F9lwsgKRHLIn6FB6GNg+4/EDANqroC6gAWmZgYnEgGsQOOS/YrrQdP
Hm9pOZ8BgB08tKsDSWkK2hULrV7YqdlwATEL1DmrfxCF9uxvHz5L+S6zJ08/
u/aQQYZtM3bI/7BWnyA4W+vC+1/7fW2WYk6PISpUlXSuu7WoDfJVcrtB9022
GyTcxrxnN1iMhCjpQz4mF6t3JRrl/wgKrluxtrGjZgSI5u67EiWCLdoMWOxN
etERI67ItW6K97ENaErBuHSreHckiV3dpzc1DsvkpryK9lOWG+c/bLXHMY0D
TTGnzBbtNB8hj9zNoLYXzs77xbNTCdrxDP6ukmyA8SWPFnROTJmwLjXOUK3n
DfrXcKJrk2QVLQCycTIaBMYtSoZr73MKo6qYyo4ysmAcKpSTSMUWzTc+INZg
OaH/tZQC70GCKR6qWFMIFfDR4WBL+wTOtQXyP4QFsZxdkk185T/ehBdPzy6J
vxR4F0tKtFlBog6RKn0Z5vHAJxYKpaaE8qi7UOY2I+aC91FifL3gA1OpU/fR
ZjDWLFDf9Pzj9mgytRLB9u2QFTqKsg9CF5Q4XcQ8pd3wNpR+bBnfvFDtLeQv
FXzZHNYltmJZm22pF6Z6PFelT0WUv5BsslXPmdIP1GoDA7k6UgNIM9/pe6d+
tu/SwwD5AndQl2O8Qmrd9egmiDULCsaM9wezl0gmjpQOF1aG0G8FC5KXsLU6
GutCXQ5geB2vWSLzxPN3VcH57uPPnfYxgAuKudP4y60/+auYv1UxvNllKA5h
yxYjz6tLV6mbUba5vX2uHOPM0iJWODoM50nftbSj6yvHOnoVz0f0IJ6N66S/
PbCzhV2RTxWZpIeuxvQ1fcSTqXenCZUTN3U5xtQ6/5VdIiAyquHaMeukYGWX
j/PQeM5jsLX5IT//MilWnaob3S4kLEwPKbmd9csxpriueU1jEtMNEOZ5YEd3
qPXgrWlO5vJKNGdbGKAWkEsWXSatKq9bTD2gN2tXhEmuPa1STGdmH1BgW82n
vjitBSGKFKCZdVvck0mN5PR79yCWLchoKVtz9pNM3k+0XpEa01DOF8XuZoFj
sH0BmXmNXQaMZazEUaHuNNgeoFjZAsRYL/vw/2aGPcGa1nT4TkQQ8NWeM816
ZZpyuHyi4uNiGXoU3Ov1Arpx+2sLNZ7Omy1Vhk+M61YDZUP139QJ5l+RWC2w
aGeItHRqRgFI3Y2pPp+4H7DVBftB0+eGMWnCdFU0Br5nj6FwBxg6SHVvpPFY
x6nsJTP7wMTht17uEKubKZsv3rwSNnYZ/IWtW/Dd8/INe5EMsvWrzK5rI1/3
D4H97tJPSNaZt6T9BgFiXTQiYjixithBrIcmaMtgOnD9D5c7nlvP9VNW3oD7
v/sFsZfbeTmWcsm8zkh36wtXiUc4Dg8hw7lfQ9IZUve3/7HlqHc1FxrepJ+A
kGjF7drK+HgCO4Fb1Oer/5YMqvRyexlg8A7J2v0Mk2Xw2YVyKE5SCHEt2CsE
Rjrh5+AJ9z+PgNb6Adjeg+ikqe3xVcIzUYXKXBQGyIOdSs7zo4Bb68pyw5KC
09OJTWVpf8t67IrLsHtTiT0AZLflmibXPXC53VbWXobEUv5qq1KrLQFPDj3G
kQgBP4QkKsYlFkjKGX6xaZoeFM1hXSth60EoF2tyYjBuPBwj38QpqfWZBC4z
DiREhcfep4GTYJwFXNY6srQCmhHh/5B+B6iQTPbIjJ/AyaFc5pOk+uN+jjja
NziRT4MBW0HY448T5ApIkemeCaSXV/ig7zOyYme9bnByevjocXeb1Lzax43L
wm+lEV2C5mOICBeQRpCJXs9tj3lxjhcrZz7cokNZMtrdqtvmgey8M9+Vmv1H
+ARSH5j/YCO+tuExkv3oaRPnrEYgLyuir5dwIU3coUOW9lQ9CT9TQPXLvx8F
GIbIJP9zl3DarYutVrNtVvXZ1Ganqbn0xVCYOjQa8itcIYKQZudX9FE2RWYv
352e7qddll8hBP7rAJF8iCylExM/6I8woOG8yIuQZAaEkfbnNr7sbJUU2VG2
gco2UGokRB9yo0aIi4aj9jerb6yxtSuzlmdsu1NWly8A9FkRARyAvMXU0qPk
RA0yr3m5JanPxSzdcnRrNFYOs4NltSZ5qY4jxk4k99xrmx8R7PVMIeQ+NURG
PkrYur2XTrPqy+aVf6fsq/J7TKU0E+UGu9MdFwsL2aW5eGfGoox5eC6RKNSn
AAKPiQwwk42i45YtVslMElVUhGnWpwnmsO8Rv64hoeJq74oxOYErsffU7M54
E9OPk2I4T0+OAB8BjIew8krc9uZoQdMgK7jdvggGgaQKNYNZd2LoFLy/GZCJ
yv1LPbI5cSAi2gubY818XT6Sb/S3vPMIqixa7dPo1w4LVRnV6AT4kDKIk1Pd
zB85RhzZ9ibI0i016I/xky0A4NDKLmpTmLta8br9MFmUJtRCaXpEtzP2E892
87ToRLVSLus1wsJ5PnE454h7jHiZzsF8A05lxKTnwIWoj9Rcft2oVQ8S58tK
tmwLk35p8J+bOOBC2AulU8fJ2YT6DcpVXqJtlmyeEZweWbRroXXio34hUfP6
W+0BGIMwkmNHQD2VQ2n0o3Q4VnJCVxYyD1kMgCE0AZTqy3mDUKXYWlu6s7BG
LqlTe9o/Hmu/OzaH3oYC3yC3NAoSybPd17/SkGwiq7yUOC3/A5Abit2tKsE6
5YC+CKWW5iXsJnjUx57GxcjubFhUNFLiWy9WWtJm3nWfvWH5aEgrFzDZxTNR
2a2qdyIJLgcejqTHRG900MlxAFQcAbBdqq4ezXFo6rDspOUuWJT4H5hEoiyf
eNFR9aOQHBT+oKDRKTEIYSKPovaS5qx8Ht0SMONL6nHlfshN8BDJOexL3brZ
BngWUrOT9pp7EtPFkSWrI96TiEbsDk7IdIqvvd/RTd4I0K0ZCZmhPZgUpfxJ
btg5r7bk8nx6C/BvK7b6vT1h0WrCRZG0WqceoIw07soF4jYPgS+4B+gQg0oE
joggiGOlDYaueOVM8nCT9yht1EvnQUkwZKz2dH98HNuMlCR6I6hp73K5GZSf
WuUWk451Sag9zgH+dLZ1IbXgcBeOaehAA8HZ4HMF3+IysfAz7m+oggVHhHvc
Tm5mP+JQRmtTpPhkYpyk45pgeneZXkatpX+kjRYOGMK1e1lnREAqomcIfmfh
k13/KIjBrFEkN/ErYXfyPWAe+Hrojspz5qI5OXGPN6gbAdmuyDP6zE9zhG/M
rvZbV2CHhzfGHPBD31rOm+oEfRa4Iv8Cz1FOzjYQsXXwX+2giG7PV/uamfue
Ynw4oSICjRkunAKYpB8cvICvQ0Uhubbw4oqpjShLyKqzJz8Fxa99eNdLpttu
YeVMjtlqOpPy/aeQl9q4TX/ykMGM4XLR079lZjsA7xv/PRa+IHNHld51NqQp
1+yOt4P2RTua9kWdS1fKjFOqV8i5LmZkXPblHlBFKLBOI00R+r7veOq9eVcS
oxGboeI9a/wZlrdEfWR+3RKBzv55QIO9xtC54zJJ7J6UxDKN6ZnNeiPZ8w1O
CHFDwO7gcbEG/Uok4nmcgYO7yBJMf/0ypxAUHq+gz9c3Bj4SuNGCUsLgosG2
EG4cSQ8ayGxHZiW0DvhBDxpB2092mCAiGXnY/fjeNSvaODWr588ciqaZqyKY
JfUvhiqta0cSgrW2a29k55tvE19JezCu1YKiH6VdCSOlKwf4P7EaiDNFVCvj
mLjNq3m9dgSEwKZ0N0W9gDo9/js6hqGqqLlG6Y0RerubYGXy/yXUShzDja6U
tOusrGDbGV2UHxfzpQ+F6gCauwg0nmWS6bbT0r+0U95KkbsAZUXw+/pXLefM
Fkb7BC6PVj3XqEyXLQohWvbzJim7i5A4jb80UFmSPzeFzYDfuw0k6hg+Jw9C
2FrorXvchY3XZW1BxohAvEMZrX+m+sB2DOJe8VO0vPGLaRBJNt1PQ4aI3i2y
AQ44HeJwzes3L+Q4sTSe0Wlp9jDAwQFGg4uF8O7QXcevpDeLxxxg4C/9Lu7b
sRYIbOYUTUJRP0Ww6Q9+uKg9HZbaQiwyoFyvbxz2mUZiXVufL3tFuh5fZNJJ
Wpoc4FkKy6KiTSnxjeuPO3/BpNBaelqrlv2ejw4ljt2DIA9Il3b9IGdmZMaj
uhThZTEYhioxXbznpDjGbV4cfHp4S6bFIgY+RevU8kqrtK9/uZJR8cOCy5+9
r+9ygWqfgh2V84xiJD6Zy/GPGaVKQO8c3+eYf/sAf+XwBoqh6yTIqW9Ag9TQ
bHcTwhxga8lDQr2wB2onWiw6CWgKzBUqgimECa5R8wO2dRgg0PPNwNPLVp+o
OeivTNblMpilRShzwPnDWkrlCECTYRK3wc6ZgM09N8mEO+G7a6I9A/sbVaHw
mXAaEW37SIk2ZbsWqfcVGbNFEQaLmEPVY6EET+IV4ZvAcCtudagMqjBopJDv
n7ARyNF44Mi2K07KAdyaDRysegvW3byw7PfFHbk325+kNtA0oFutR8VG4rLP
NDXaxtQTF9Z1QGBM3g3IfNDY5kRnN5mSXlOYVvlwMHsJVZ4t+YKkcuKFuYJb
b4KuK9VkO8Npl+G/jYpA7s12p6LNE7p/FfCt87/a/4it4NRrvo9mEDD2raPh
PBrK+NHF1Z4OOCVnNlaZRiY3i9f4kgteKPFbY+RSJWPGAr3wJ/6qBZ6c4nC4
fc3CL0zfCLhh9oT6WtC8INnb9yLkKeCu4dqbWfOB7J2dl28OLDIZvL4cqF7J
aht/aDtLWrC9E0zsOTU4qcVVWnKz/2sbBVgZ5/fDAc5pNf8LUsw0uPD8plPB
jL44jJHU5hLfzIgchM2jvnR0yeYngrVaTcoB0itjTweayP+1pEhkRNz28KAb
Et7b96Wc/0Rb5VGImFLqH4P7eajbWwWGghl+rGqP+XLWGVG+qLvUlbXBCQnq
tkEUMXGv84x7kFRDVik/iS1RbNNveYLTVNxeoSKxGW29zneQBVeSU/eooPV8
7hdf+rloRwJFtvVZlVyqIpAEdNGiAGsF9Gq+Cpk6ekogTYD/CSyMakcsCZon
XfOZN98eFR84YhIBqYUMCFNRJyqrFW2KpRbgsmwfzk+r3Oo2w4zZeiCWZaZu
go3CfsZ9P7iLKA3wDDvukQVxiXvYS9g9cNMvZ2dh9x8x+TOVNYHLKpb8nTuX
y3ziUfkr7a1BlpW6iuBnH8NCB5J0AL29OueKsWfVyjD9KEyhpjwGRIqW1tKx
EHvx/jYXrW3PRX+BwEd9F5jojT9cgRrvzZmcQFaYZQnoqYZwnnncMlrCIq6p
nYoepgQ638GGMEadUcdu4ph0Y6pYiap/GPchi9TjAus79QQflLviDW3ADIIN
2cEfkCsHvhoWzMMhuG++EQf6X2CasgKEqlu3nFdU3waInY8LKTBRmNSFMQRW
y6+NK3U+t9ZY66Dr5OmYs+m+9l1kMilXmMszOv4xHdlPmEKQz03Prcjri8YD
g9PtsDE6C1NfiMrpuM7IitllfCwMXgpyLSFB9lQWpnfCiAjrejMIdZuW7jfe
dyquck1c8CDUoN1yZIf8Zm+5C9Uw4yORnoSR5N0dYYj9tJITByIp1VOsHhjJ
eIL22gH0/JoZuOCYPy18gguWwrR9Q8ZEip3kJUHsIf4Z9ufQX7BeGZsqmlYm
WZ2lwGemtIdbSn7kPh+GkmP1AfB9pIpOmShSWlAFMetWcWxNe7Wy3Dz/RpWv
lct+YyJwloKja76Fihcn0/8wvcQMWmcqtEIzAj7JlNg5/MQAct/1TKaBF3xI
/x+6z+m5l4jh4C1bEO9AW8evUw/51GMLLjxO7jPtyC9mFxpT72hci+thnybe
oJjXg6uKgw7yl3PL0BBUJvPhacpbSc88+WLaYzDVbRHozLjQrLIZDvwM9Q5s
BtMZyvbvk5n84UjcLkGvtKnocR4+yFr21wNr+WrGem3dt7gt3k6+JEKqG+NC
FCY3TYR5w6IRVr/DxSoPvbArfF+rGWRooADFQhx+Gi3JsR16aTg7LwEUIo5k
OZhRXnNPgT8CS1B7ZvMiEC46fg6RNYmDyE6lKJrvkrqmDq4QJQEJ5PRclfVb
jhL6o434G4M8elwt+g7DWu+Aq3tg6ubLsYeoV/1o6vM2KCyZc72Un3+Vv3Ud
4SX91S6pSOl7zNRdf9QB2DLQNrEqMEPhVbe9nEMPn5gbLv5cE0axJgyquRVD
QoAA+FjWvXbuMOyhzkKBSpG6avBHw0pFMkjs3G/O/jOJf1WVLgSj89BYN30o
lGOM4v9cbdD0pqssgHOGb9K4fWVPfula0pq/svZ+2CZM8xK9uUM117sMuLsK
chFVSTNHmG524qK1OBqNPYi8aWD/j7TUQq0WNECR4pgusgzj8y0rSMFmaB6M
q84dFa/sOsFfhcUSot2VwDQxxGNROI2o9Va2pDrc474GEAAPXHmFKX9A0WhP
BWt3FZFVVYd9vq6gfw3xcVtA+i1RHZ8QIb8+M4Nv5dpqsJE6CeXokHK2LDXy
Z4/ZaGQUwljCrRgvSVEWaVDQNAEpzR4u4SUUNL/QALeHyjjowvjpYuFz1Td0
0MW2gQqho/wOcxiQ/EKvZz5Zx3XiW7H/DWlyz5e4zVua9WNZwNPeW5ulUugB
PU+14lHlM2ISZp6FhnYGhU3KG0/FQHnm0paXKDS9PgrTXCqsgdnnYWhH4H9S
Pm5cmmEB++9GeGHDDrkPu2iHNHMuDElQYCOTzg/S0INBVzI7K/2WJUJ0Jf4D
uuX/BQfPgvS8N5M9J8O4BqHYeLLjG12qIo5oUWRm17ZGNZhn3tx4R6exfd1q
CZKji0UCM6eKKDwxyOBZco+32LGzAbPEjbDRXr+itG7v4ZE8QtQ5HHBQGNjV
UiWdgQfPEz4mFw1cH3tBnwn/EuF9LGz0Z6cQ9Y/zZshhtZ2rYl+nl4bBdXRu
TFp97GXcXuSke/GUcWfTPIahVO/bskudCdBi+3S8Zn5oqoJWxrZvetU9l4YJ
Vn6DHM4TZjepajYETRrzUhs08GrQzii4GC2sg9kYY/L+TQUpwzGHnl9Hrxo7
7AVQJUBXI2AnEdHzgmIwFyEQMSbf8xd+XLo5wU8e9E1WsOGdq4+UfbF561bA
zYp2GeziIuXDw7cbHqgVxasXOB8Aevzk8g8IxBSLQy8VUQtKHfcsS6G2q+Nf
tLdHxiZI5jA9adbLC7+g0FAR5fAq7Wzx4zp5pUavfLVqHYTEg6VtllpAcJl6
aRgG2GQALqvDDRRKEBY09/idjm+Z6F97OOz0jo4If/0frjwl8RXaNZo2Xe6B
sEmIsNa3kztDIQcz72egb90g7hFToZvQcqGhz7lJGHzVH8WTpLumI93uqVUz
cxp18RgKP7Gmc7R+l5JTOeyLhumv4gY/gjut+Qp9xfLij+hQ5kvOalZzHc9/
GlTXpgEZiV7SgVoJrQnc6DjrtU/6kZrVhGe5tZLT2aobICOaq2Byrgv3BvO8
OE/9vnBX5zz54HWbqkIqSj/ppk4HJflNmFF80fLmaHIXTo2pIw7Vzh5c3w/U
yywUyaUgaTVO39B2PkRMOWUfkgEqm3A6oJOMQcIqdxiPY6ouOCn7z9pCcnWM
ahtuVL6tx+t8xSQnjEyaYBYqenQtCH+OQGK9KmAbejm62Q2cHRXxJ4iB+E06
pMjQaVdnweRfykjNNB5jzN0w2IsiNe8/qNYURQgm19VA/L1Fh9ToSIdKtZpT
qbtazkLVXGnnTFBuK/Be/cD/Yx7g/++BTYyzNFyysLX1x/n6pyWxjI/E99pe
XMzjrHXji/mk4CC/1TINY0iK6t+7HxgtgAlA3cDpCx8O+G9APMuaAbjjKHj2
LExc1qL+XYmz/mjMU4lOPyFnrjnwAp4dDA8CglJE59yUAYOqNem1ESRO9DIH
rNtX+b8WjKKI5+W0AJiGQBohqcOhU79DO6zRqbSJxZZz/BNtmmcCTgIzyScU
4zoSXVUFJRQfK9zTiK/SrCY6/KSXNEgDpyPgN/RVzBHEuoKASN2aSlfZm7Sm
rkXllspxpZRWD06wPsCrRoGvbzwzntmNNHd4rXpiM7oZWEse45WbDmcjEjoB
SQzsWO6Wlh3u4f/ZtxTveX5sUwCvsVvkHps6+VgDqo7HVURFsWfrLdg0GJid
/ATr7dfIoxzruUE2hrAVuFJbYPvoM+uQP3MIpZpGx5X5mv6hql31DI9jbzv5
/nCMjay4bWvbgdrLgjgimYqgIAz1xl5dAVsV4oFo/z2OVnTptPd64n+yeioP
7nyGmvPbnpoRgpw5vULcXpeDzHjIdHCX3nAYDeucOOW911s1gTSVXNaYt6vL
pdvBwbs5Dtsi/u9khsf2B/CK68ghddmmtRW8pQ+Evz+espRm750JC5cyN/RL
GsgpuAR30493nrpuAiJFt6RX9rwdt4uMn6KIoslBGinrNiz1bNo1/89U3sXe
CtO593+2cZvq2W9ENqkQ3dCVvrypndN6u+W7ZFZrgR+vY/SxOOKXa4YsotHP
w8qNc9d2/j4/McWtjvkt2I/hOcWmlbudXM5huGOzyuvszp2vkgitKZW4C/Qi
w4r2Uy5Ibys+nXfQHLKpqbrGT4XilQs+jMy3npJSzlPx2okmqCD6ls2JqliD
BD2K6oqbh3Hf2lE1FbfldM99GaY0CQgdusesO1AJzR72d4rXJEx9njsdfjKh
vWjaoufaUj67OLHBZ/S1NfCKL+cbom8vbGFvakRQjZp5CyVtGo36boh8tvaQ
OlJkam/Eel5MAa/8XuRY/TxCs8iJxkoKMid1cKQO/mVJ3MYIQKXHZHulZiS7
COhPYF90OC/f33uKYaaFG6TJKks9coNK4k2DWKHaIv7LR6GxtusUZxyXqXpx
TzyHj/sZfH+2Zsndsr89efcV7mDLdbuHmEF5I3oMyy4XvbGioCAsgDBmCa0s
7uKBtGdrGJ+J1BNOvUR70uV8/KlcPlDJTKrx3kJnV2LlHT7JVbtRgQuDL4Kq
PppjjpemM632eMG0Ck+C0XtGzwi7jwr3qS08da7dBHFAIHnZ+CmIi0YxP422
lIwcF9ZVDMtEQcVX0hmlwQUqxlfm27nZ6tU8UWbVbAK/YDt3FauXoNAdf7kq
aSp6+9HvAXP30kGymeUlACZLnJHsh6q0AvY1dzqemwbmgRg3FRGBtkPVsI05
XbOsPIDe2f1Ofn5ARK/CTPvMszZj2aB+3FiNdnpMnwDthpaTMulznmCbWDpx
sBuJxTr+gLedA6iN4Yx2bJOzamiN1LOPFavhf45byVxBtTSin5PCvmMQ2Xvy
0WF7s8wD5xzBO8QHxUuVHcahl2KVdQmRcRyz1mqTpopAA85AK9R2/e14KThf
DoR0h7eiiWOgh7fptb8Lv2Neia5EeoqHZDUjRxeAUixZ2C2n00WmHHGkFZqa
blXF5oTCUFXxp4pJaW0U9Ls5WMPzUPRfYnUY4docCydr2uHoZUf6+zEXGxIg
5BX21zODKHXyViW2CYvYh12M+aGLDETtF4ykkjH50MSkxwWklT9NyVZlQztX
NiqYYqwMBDdSVUG7E6PHu4tUWtkaEcz80yRGmrh8ee6QuaR7AEk25bg5f/Y6
hbw/HQZdEpWL1orE+QOTg5615s+oR7LbRprCLfAj/Q4IX3N/kzl2FmlwR7D7
ZUoZLZw3P+kJFCRdxRd8zM2Q1gnPwgfp0H4boEKmGePJlcd3iWNzKFbih/BF
LKcJfWGj1jZJ5WgjqPfUkVyrpoCm+zH+ROsg/pld1c0aYPEVdCjJJgENtxHG
ECWwmNYo+WjgES14nwc4tPKwYCGV9fGABc5Ekl6+kL0/Eb4eoQqu7iY1DDKV
2IcWstDfQ7LUew5STrUO9aZPw4n5tZGqI/PkJUisf/fICVcDI1AqDwiX6pgn
4ENJcb9NthA8XkajG8DnDbea3oyxkXeH3CPbT6q5NUnJYQhYPn4nLQFlQMCC
9GQ0tz+o2rKNSWiJwHWAXO1+sogEQtVusFpXcHAm7BFGZ0oqvNKeSIsQjq9O
ECU3aYQE+iC+6tWlEJFuOx9HWTeePLKETrRQkOrccMQMXMJi0yDN/JE4ZMot
rVEGHmrctueRRTkw3xcXLI9XNur1nH3i/O+skb2tJBPslVqrqJfm+R2FoaAH
c6DRwvyJoomEUFOdEIxs60NP9I2+SDbJlywmFdaL20/B+X2+NYXe8PKgycdm
3CILt/6MOYGNEibhWTdR/b1yh2mhWx62+63x/T1GuwF5xpXMiw97miu5UODS
IKkBdoi3sRGGNH+pOwikUcAJyy55zfMKegXweXV96xs6rntyEXyDbiHkSfOT
H5NlcPBzsJKOLeK3sTeZAeAobhQ0rovQVMha5oV5+8JRlKI+qdhdOA4wVnZw
9e8K0vfYtNV1R5Z2Nfx4FaUNpmO3diAtyuGeeWvviqpLLjWxJoHgyY6pi3KC
VA+R1PoJqUl1AxZu92vs9zzknlnm9w0su68eOgAWaRGocBc7b3WrOrhFZ2C0
ZKhZu+tAEMz8LMNouuFZ8N/PlJgbjAFabVApR3F1MInXFn9sU+WTp2U0wYQI
rHj2JEUlaQxp7pLJyfR+l8S0XCCtLrLRrC1yZM7bEKK3h+BOaqlNrBVYOuqO
P87AhLL4b7WX0M5MVc+hRK89E8U++IGWHBR44oKVX3D9aR4IUKlsGik9MbAL
1Da77OtSqOKJEb9JVTfJlBEoApuVATa4ru4pCQeudU0T7NLjkjfCuvvIbPh7
yABy7QDcawqQRKBicORg7gXoPmoPaFH+73tWDpMcAXyLqHAT6TcxM16p8mCE
is4g5aqHPHA3auxVp79J8vT2Re0rulCvAENIE0W8HrYLcE6LHnG9MnsEdW8z
He2kBE0EAvNyo8d/piHdwnuq6g/77EBsFezZOBxYGdstm8N922E7SBW+gzZF
364NY8WT/OxOkZeuu8NGs/jvzsJYTfy2TmBzQZxDs6TbY5+jaDUN5vFUd8Bc
2Ng2ll9u3qYuKRVZCuwD4lDRRolUYF39mp56Ut17NUv9lCOcevlZo1thUzpE
2FihzCeOYS7Vmm/vcRjcUk551Yo+hIt+ZKW3OcYW5cVOx1E/OV6MM6bFEcie
5nWsvu/TEH4R12BWJTuckhPxwQIFO1BbNk6HrOss9EAlsct1aHhVo42BNg0T
t8eOqiw0hjZWBbv5c9Ry6a/0TR+HMvjZyI0k/TFlKe5NnpGlVWfWDpWI0OZZ
kB8Zn9bchQYqEJElknpnOX/vyVG3gNyzQZGjlT6tdoJMOtU3jNlMZDBUE86k
5V5xztJqdZfErJ8Xqf3GOAVMUfoNtljjVSd44l66VOsWUJ1ON9iofKzgxoL5
q3iR7aRy2NBN4J1mR7EzNdPbHcoaOSpLdUpx2+pj9Nu+nA296FR3WJsVXfoV
Bb+ZZQoBS3J4bY4dIij1hB4rerbHlZKgbjEGX0nlenCw+pCr5s1DF093UGvD
I8up2+J0Agfcyp7WTN4WnOQZPVmnP2WozvGv7DnNvlpX2O+tjN7u94tKXVBg
Dv88uUPjgv5lFdr4ClRsUuMnoUG7uujLVQ9f/8aE19+XG3ECMLN44mB4k5kY
hDzaKcx0wb3JlGpINX6dKedWAq6Bdqxl44psDu4UG7RWhatBxY7vMs8OZGWp
hkkWemkry9U3AifgC7ZF1ZgbfB+P//wfmLJHaiKDd8jGuhnH1W2fAObzhw0Y
/q9lEzbytUTw92JWwc/tQOAvXuGFgy9JVbUT90Yd1RqZII7GSAUflIavk/Vu
qkqffqUnHjrjoHbvNIZfSkvQbseejkiol50tJReEi8Kf9S2RkZpJWNvSEw0a
rz5M/E1FELTpEBdo+3prtzT107i5DmSkEOH6bPrx1jlE9yiWysuRLB26Tuhz
uWpC62LHFc+VDU+S5RRHYZ9V08PPTIfWeb8WgeeDBddKMFFjOwjdYrya372k
fXt/MEftnhXg13N2zZBssDtyYM2Pp8S5sewtHTpm57QNP7TqdaBLrJ4DfEVb
6zPi7Zs4wDLQi7i6gyc+EP9JtFBBLztuTkrZslJneamr6pelAo+j2EaLzVxb
3S8oZuSoEm9Y4eA4iwrGi1lFhSlCll/F8lg4d7FpslyDc7EX3VBulB1VOPPI
8He+EuAwLJwdbPb7vCK7aJ0cv7Y3MinmYSY31Vj4KbTaWBGpUp1HOA6j21zk
Iz2Uaueo0rx9Td+5KCW2KDK1Z8pLACN+ImGSzxhFB1YbDklxRrm9zuq5GVmU
nlRaJrs8a2SUZRIJ1IFVS2zRI2CHzmKFdt4Sxrw819hinxXGKxq8Yulm21Gp
0arOCkCxtwRiPkeYIMqMxhD1BE620wQf9In7JJbuIVTZqK9pB48dDwENlrXn
cF/J81+ixtkI5HEZa4FwDmLEYrXYcrgT7I21jyr8U8qkNvBMXB0kZrzcPEp7
JLFrot0OTb4s8DoiRJnrNyeW1imsP6DHTqxya0pC4vyIgYTbwK4b89paH+4Q
lY9OGjZWYIudnHtJFdtC5Vpm3OR3OI184rAYG2gZwCTZtxZboSB/GdsNB5uc
wC/FEPIgHIuJMBu+kasYaDtPqrP5KDxtFoA70UbdmocSdKejl08+ZliNMxkG
UArWPzQCmBtK2K+PqjxLY3deOrCBjlv99Xd2JFArdRsyOPl4PtNkAuMrHkQY
TE4uy+zwoEMvtDCiyNr6zrA1+0rF47uUhZgfI02upvJ+cHrs58GxgSLrGKEa
5rPjd6zOY1eOfW6GnAqzclZBryVKwwb/2AL1745/FrEHX2NjdKRxrf7NQeVT
VyR7jUsDgAk8HmyYZqq2k9g5vf5+Vuns41jEkkOfOMdueCbfamueqegm/Yjb
CV7gcTaSOsKvNmrZdt8Pk3/qyMcdhLZLCwrQPHtXKjta79RlggxDC3jJfWtL
epz8Cr8PXGGjYJiiY9VV9o+RN73fRYnUtb7nI9NQA5MeCdAxTxnEbgqAUvEL
WOMNV6RL/9iyH6uQSw++ybj6/zO1vQaOhM5IT2g8uno/jqKqcHxPSja6xFib
xJtYrnPJ3vxesPX6QO4Yo3a7sItM1UONA4BY/UQauqcFvGc8RFuQN5fWhXy4
J+GaU6NLl6KRyvUNrWMONLQimFq7nzKuRDV1cvSehsyZpRwT2H3Ziu0F1RHj
5B5vDuJLblDPUlwbBciy4KJmJRagXum0WsaZeu6+Ch30ks04aaGLmP/uo3+1
8gAzFSfl1HR1Hb5Nx64KLdY705Kqkw09UZHm6S/jVn3vqxzvS04mNkssrFx6
LYhUPbr+IqrYUMAx/A/YlXXIRwkRhMHyuVpAFrEtnp9edoVaNBz/+FNbCpTA
VEgxbWdsFrq+PEioQezaoXPUUhDQTnYT41Jt8YQ5VJb2W0NcIhgtvyB/RpAi
EDOOdDlFLXiSfs2fN7TbP/WMlg6zkHRChSuHB7AI3cbrw5fqYBN1vXp4BYlZ
jAnZgHyZthNROfYV6mHylFlPI4KrRd6yX47NIPitctaBhQ3+1EzPYuhvl1iG
rIAk/StyGdMvUnoh/QY+XXGZUiNEIwB+L9vG5ivsxHzO6rNyHwvo2wf23TXf
JTu+62WxAMDwyi4qdXqpIvNAOMsdkRYBv3ce7X9gqnn7dI6AMYJitZt5vDzY
gGH9ZOGETpQbEbrh9zbq6K45VU28TYcjaAiYFTS7f5L7/JIanyy+Xy0arq63
mjqDk933DW2oE7RHpNdb54CKhgdk/ZFXu6U4NatYltUwyu9KIJtv8v8V45VW
OK1Tr+LJ5/SOuFSzUgxoTMiJdMKP38rUI8JsRT58d2xjaC2RENo9hPZsRFec
qTcM5jvno3VNkkRjlehbOOgiEr6TL5uJTk9ub6oaRDhcFU97bIqC+W+FFyRh
/gavyAYkTJ7phXmIU1+TowuUII+HL35BxVVZi8K9OubPv5TzZ8KdGfmDV6dc
OUJVDDo6v/DMJ0Dwldr9xf2PtzT5taMxilDLGPb1PvARQ2OP9GHHy4muudJ1
5oxCcpVYgYmcKC5t7YoqG4zTIbmpxgObGuZQUxbPqBF9mDq0ZLqXDfgGTD5Y
ZDYioAMKZSCnYdqiJXn9HH7G6EgpxJZH3nSbUz4KocqGZQ8rUvPvMtceZZri
HyhZ4P0uQJQ3yWsn3X+obELg8aiD/kYOawW/tzCfH8ns2STR7rE1MbNq/FY9
SHXR50kPW156qGPr2ZPXiGCagYOc9Urd7nz73epzw+6bbUF2vVaxZjJJst62
47omRRxtoWDoCORivxyC39p5zhObWRWvLmQGzLxpicoZg86qAOMD9zOv1Zxh
HY38iyhOP8d7f5eNG1Pb4vcDSJSdPfOkuJwe/yXsqgXHfEv24qY4Z/ffY2kT
RpbpPjjORjqOjf8NQWXExWXB6JnygkNE1rzTqdpr1b62UPwLo09E38lnrDqs
vHVZhh9tdQ10kU43LA02zdNseL9FAkUQo2tTW+4Kokeq/JH8JMLMVuGakKnR
8kDiJa9L3ThtiI1qekl2rsCYDO4enUS5e1KENDbcoRsdbek+d8BUgdqqEuHg
hOnQqFzHvEKaIGA08Sxkn3CfZf2X0lIx/mCc067cxPQHowsnTfiURFEAjafq
rpjE4240JhTMD6KMyb+Uccn3yNtxBbikbNMCcW1QuS2Aj4GzPodE1Yh7+Ybk
vHZclfwEgN/KQA8j9e7/ugBwSrG4dxLqRW95h6GHGJDOMlFvThHV/mwMS+oe
q9N0wIP3QFKkO6rw9tZafUGcLy886Gqmy9BNl041vJ9JxNvmKwzyIcxeqdhC
gEWzi/xDoMUHE/YoQhvmBRpyyjKfQgOgen6uA6Izj4CalIVqkjY9z3y0mi8E
ktlqg8kku0WCSGE1NBtkocyHUxJTbXj3PmUdQDKbw6Ik9HV6W13GaUOg1JxV
WbmDpkTECleY76P7SZoC8jJcP5f9rVZVz8RwskCDT6qVzmqf9oGMX1dv8IZA
Fqk2Ds8Q3EXinSuB1hYp/3OXlF7ouTX0/z3RDT9DmbdLJjiZ7v9a4RbHrB7U
uepKbTyGtz0W8cWmvasUJWvm/K5gyMNsuc7gQHt4GnkPaV6g3AG75AjEkg6f
q+Evz84tgr4MXvJhxpmJRoof37iCYHs2PKRensp4Du2fYktWKVnApbHU2IDo
ZuGDiWxgJE5Gf8Qw9HRrLltt13thaxnRTNyfLqPiuKUoBON3yAscTnweLXoS
+/PUDYPA8tSaaDfQcccxjNvsCu5iv7SgLNyPQfwx1pouqTeaFDRsv6cfQDyv
HRgX+/DTpUlSiovgyu0pcn8C6IibleVpqNgg79o0oLPxrmvCzJAnj0wzeI9v
T9z0C/HjOEzR4HDTQ2+BDYF2vSGJyFRpfkO7hwfjx+IOcgCA4E4QkWwvE2YN
gmchPcImLqfKqn+bN6/0KODXckOLQVIumsmei7bD+FoEoTYYDEthLAmM/LbU
x+qWHxDWUHghtYSBg+fNpZlkZE29xx0G/Dhv+O/+CwBmLB/iXJXqFC8pvOiB
nXLXBjxysue5uJqClP6ieORzPJQlyinLfZ+PkMp5s+0INvfKsUSGKCs8BOf9
SqhEgIJ1HT3AqXymJNg0APJ1n/dMGglkM/NgBzCz+cLzwfcNZmLaP4ovjqSa
QS7ijsZrJNDBd5gjhxua+N6w3V9FgkVYWNrmyObQQj6YZnL1eT4eoCA8cRYM
BbovpVCBnwriFFGvJHThArUP/WqOgslQN4cv56R99LkCTxW1PQtKbVKPY6pO
wMlcIR1xcdT8vHMkPsUrdDGwtbeZn5rrt0mYbZ/bHqsPhVmYdRH/bo0Us0YD
w6UNL3M+XUrQsGeV17Fg3NcNzkcSNhgJaDKyknAmFCJ3/rCQCClEjrYxqRoD
pPaLGb+AOmwdAZvkvpjOsOBvuNtwqtKORXXakeMKKrU61CsdcAnuBpc1vwpn
ALt++DoxZ+ftb+PliOwbG1EuN7o4L0sz9V7sqKul9+hY7mYY0vkyFCsPLrgY
JlmyC/FDI/FGYV19h8Bg4x063WzPq/6Jb5L/vmKGA3hYHT1feSIY4bn+QtPr
taj2bxWRFyGfjQ+JjPrh9BkTLZh6aLSuDvV5q5AapXV5jBXf8em9VjQZ1YQB
P5m259/zmwzpaH08O1pOnD/gCQXT3i599CT0Xnx5ZZznOhwATqSGioLJ0WCb
1esgqGxnAOF0XfP37L3AWhaevOeuBxJQPAtndT8BGACIlNBxy39QihTDUfTa
poK/EgMDIHU4c8HTr40We2qbu7CMuYJwlxHIfzOjGnvsKDbsufmg7V5hHb6F
p80xSBUCw7Wp8D3KH77nO0mbaJhjGFX6IMPy4fNmYoDecHcSi8HsoJpl4kD1
VAAokP/YQCa76058B30JutoWpbZ3DT2hlD8ltiyDoLPNksip/M7EmabaNglQ
F8lm5/iB75Vkh+P3bCOvCEd1U5Z6U25rhCVWXNhr9+OGhLkNgEhdzo2JZu5S
JA1Of0mfIhYtrBFefDSMGXEIO4F1K4igs4wxJadEjA4GmQ6kul/uVtL1zKOe
/dxQaEVTujt0sEt1a46u8wigh06bBxqEE6D7qTp38i4yZSUpAHgjJOoAZjdf
QR5ss7RWFbcfO4WTdH6deHKUEZLvSFc3gOKunBr+aZ9G7wnJpGq+1w54d0kx
QmKDDLDTOmANdpDp2R7f6UnxxghjpwMzAaxIpcmsxe8NSCV7Q6UfpgCyRBoy
0f3axXGgMPgYjU1xkwKJtdt+iE97oXBa42lwnrVYwzDAnjNB5pvGv7/hOb25
0yt4DFXpe8rK51kUF+C3sGJmNzjILTYV08iUznZfXwZady1jYLxdGV4JnrP6
N00abRQPrLatZqYN3u8VYUPrwztEHsGSTekK7SJFTu7ArpPSUAqH33yB6eih
iMHz2d2bNW71YK9Mk7HyyTfmWI6+/cDD1dl/Eq2OT4TFaG8hFHdHN42XN0ge
MRtYkvcECUPw/Oc/JDIFQ00sLUaXuhI2DRsPiTAKQhM2cXo17C90xQtVXO9v
V2Q0P8IW8yVFHyTZS9nTfhhnBd9sygsnf3/pLYLKIqEMqdQLNUMd4NdSRwpF
f5/S+M7t3JUYV/GKW5CYuihl1c1RUFwBEKe461hA/FMEMFnQz2WcFwmiGgMC
y3qUDSEhRJoZnTZt3yFwYO6CCRqQkxEMvG7hokpcvbARisaPyTppJjMhBgi0
pOkiO800H/KFo/dG0tCAjcgYnHmHaW5/2rmZbjjZ1Kf7cmFCdpe0hVm2Mi4Y
oHftz0yEHRRvLx2riisBSSXRZnxOr4CeNr+EUuqB7DbJIrK156uYu9qmLc0k
rrT2tOrEpfmMkKDtUcOH51egDZN6Kyvn+rCk4e0Ux6UF/HEJp21y6JkCXOwV
q+y3QFL9LQbRP3unG7ahMJm+aNq0ULDKoCAoIudvwtl8yStbvyCC4afZF++k
mHc905evxoZZxJMy1KHrL9QXRd7TAh8jnN4n7KV1iaCj0prspSGZw41nAC9j
sh4BMiCpuUeyuegu/pXbEan+cbie0S0QXkYzNOvNRvmYvicAyVZiOax7zUtt
S+TQgRxGSSOVQ+WTkh0FBm81bIAHX3Hlz30qIk76xapDbn27JdXfdXAUPAjD
yeoM/13a4RFSAwXqy+DT4M3z/2AqzxW4DX+wLqP1RhWh8BeQgcwzcdSdLkoO
E5rn1SiDScw+6H6UxbWSq03+WZvdF5ZFkXv+TpMPJD+eBtifwS0IfcJPSRve
jTzMoIPs14s9mSCuhQV8ORgz9pal2SCvyL+y3HxK7tZ3zCFP8YwSmhd0SBjD
Z5/DTO9L+mxGS2SkXDfL2Dew8OzOoAy5b+dsRsdROxc5u4yzyIKY38DQt0Tv
NQOD2LwKTmqp/abN7Vp/b8n8/wxVUTFx0U1Gx8yvLgCLfcpkuqdKolQzHKqc
N6a5urhzjYBjqz/ani/boZEKgnHb+dGg++S8QXw4w8zZme6ifJ7i2IGamt/Q
czfouAbbg5sUbAJ0aoBNs1EjYotCu0qBSreFYBE0v7Q2wrh3Xwg10Nww69vr
0EW79N+DTlRxuBekNqQDH52WOw4ikD6qv6OnZlsgf+Ab+YE9Y5LzxFmIcTdx
2F1sZ6Y3J6ytMGFvaW8iM51NMVrvpZHf2xpRuCUgIYe7IWt82wz/fk/A/X9F
zYFcx7u3tABCtDBZchoB/X7qW83iWNqc78EuT1nnOZv/zziseEP+O5vxMEUI
uf5vHrKLY0AB6MfJG3ryR3dD0ixujon8oA8D/JOkkVnCCs5UxRsMVVW0LwHO
x7FggY/2fMXNjkEyQJ7SN8HHTFE7G/4lkpb0tPEWQc9TAcy1wj21Qd5J+/T1
dNjdx7vcbps8Y6aEnWrdDQXB6iSoZrj2nkWMqGwd9vrWjWGiH7QazmDqzNWU
MSkLL8O9znIBGKv96yDTOXjaAIZIC3ncYRISYkLLU71t9q+52x9JUeHMH8Rm
8+z7R7H5ztXP+eHS3eGMUZtBo/VjjXs5xKB/+E4wcjssbwLB4SQMWl/VYYaR
zHTkKp/hh8LRkH59XUrUkIwLE/+3tFChhDN1V753VzCVsZXWN7t/I4zIgyYB
u7SFdtyT+kmBz7FCl9UGaQ+/yFOPh67pQQKcB/kdtjHBYln3EpTn6nH9wWdl
jXy5A5aZF/kS0mauitr9E/hWN2a3OOt91SvUbXvOlViaOiwcVWLwWHPb73l2
Iwc8WDjBqW/b+sXRnvioNowZVxMCmPkflRW3iqFjiorPmjJtr+jNGv4w4v01
VO2Z42KmrVTW10/jfO3X09KOr1pFDuGS+dwZUG0Q48+mnF34G28pdy88XFYn
42u/bykOo9hindHYq5QC0vXgOAGdZVaVwsJGIEAfcPBKWAm/xtrVTWZx17IJ
r641SVNM2RGr9vaay08YGRUj44KWEjVIMneylAKwdThUsCwz3rMokH0TuGMj
tLnPWpg07FeqhSpvc0BX9TuCV7macPMwIZvwWM6lEbe0qQOKIIJZtuvX9SOT
tB/CxtHlBQnXeE9/dXhREdlGGLEWdbJREtVdBh2tAleEs7ZVutqaq8MfLBcx
kMBMsFStG2oSgORwO/rDlwVRalKDRcYSw8DByB10/0hxZwHzD+I+8p+bJuXw
olRjKL5VyNUcJb62xota+IcqTfva+2emmCYQZOM+RxX90lYoRxOyM3idKXk6
qESt/0HTDHfLORShNVvB6xuNhHsNDWvjQTQ0+sB/7mHl1mHiHAk20822N5N+
+069i+IOhKv5Qc1EgAG01kpbW4Ef1Bzez66TYmeBLa47NB7bSnyJmaMtwjDu
H6k3EULvUlwCOA5tehpTD742eukEGfMavOBoTUNL/acbna3q4gp4hfKMmn7m
9DJo79WvLK80Q0P88aI9non6OM0G4R114bb/Hc/QQabhNoz2aXSF2ihGu3Q2
D3zYM4FTjOqBXbdh1NAD2YO/6g0Xld04NswPBND5u1zQpxgHKMQxBl0Y6MfI
uxj7+SmOItv18AHouc7tq7+S5NvmDTNIqyZDyqzF/Sbh9FTZ57EMTZLSrDZG
Pso9gdcclLSxLg7s8ifmeKixI1EqxFdZFC83ZG4e57D88X92w/Scn2dxw3Gx
52Oh4SAgQK30Mod2A0OWw4z12a/Ox/vMEfV0X4H/i2do8SXcno47D3mmcOo7
7St8mZCil+76IiGGfHq+R669Gml99XT2uswgt6Zc/zurixhuaQew4yvQWRY3
2Qs57iU7sroS7N+p3TPGwRBOSQRAhfltxACJNLoBnH7Ke3Df+gpcN8K1u8rV
qd5qstNhf7J5xIUHDFlukiIX36LMnfPisLn0fmk7WUJOQN+2e3vOC0x/NmLz
+WUniOuFrsdIJg1RLzcAfVbioT/q9tvsG3bMhwzpkHV98AATjShJhOvMN/Ab
kCB6MZU8J8SoQTd2kNV88epwf/bpowFbOhSuim4g2gtWFjUq5W1zAiSi7E0v
zDaDFFqEivNVVme7u/tEsbcxb8tKOXDYONMzXTILzDu0xv4O3DIhuGZYaAYF
G/VC7RSEhQLTEeabEFztK/koUD2igzRPt+Xto7EGDm7UNYChlIWf+ytFN1BH
ubgLuB4jDxDKcdy3JC7ENYfdpFO8Bo1iNm8mnHxauxG6JYldeTPu/glapvMh
OUzW6/D+KBYcyAWcPzRzAUG/wewB5FQJW/Y0zNvT3G0m2EAJJVu6UiuFAeTo
Dm4JGm49JJzqPQOi+0e0kL5y3JAc9JrCnPi823ayQJvTmSyCwG+/Xgy2nyob
D54iQMD5E3iYPVKynYD2SPeJgk6ItWnUs996b2gU5JjcbGSUc1IrrgcEFxvz
NwcPNLqI1VdbNDkXdZv9iWkhs5V8rt+FBJgHmhHjUJLw2dzV7wXDSBLugN8R
u5yXrk/LZWryKd33zweNVgoat/1/kV8ml4EOvWV1+KFeFbVRNR4FYvSj5Z4x
Snao6iBKoQqrJA1lhS2JbOrp07nGaLWAkHlEAzFReN9zQ6bah5Cj5K2y9Kdu
DP8helmt83XNNyO14f5k9B77s57tbmL3FkKc/zUs/h6ornUxPwsTX6153Ux7
k/zWr9nhQa1aUWmlcdiB0TIm/xg2OBaWc8/zpNp+ZqUiZqOO4MWSrDn7AMtz
xsgVxjD4dpu3KAoqM5RTiBd1MqL92ElFEDxQsFCj0ttG6rggN310tOLshovt
9M81MUYAntRgifQ7hE0wyUZlsxRGLlv1cvof+wM/AXGFAL/Ut88b6sn8BV0K
VONA1IgRsxOSdU1VvFFmwc+Qb6tVYOaFVaMN78KY3jLqCLQiXdhnowdddowd
qIBHWnzn6XisgrEM5rcCP4T10cgfqx+lXiAt+jaefJSw5prkMxeBJ9NWPl/0
h6g3GWmEUeWUxTH0lLV8dPsPh0fW/OwIzP3YmIw4FS6iBLrZHIPz1MCyraCT
KqZNw8TVaDiTa0567pDSmz/YXy2LvphtCUsJwm6LwKO7kjOH96HShGgCEnQ7
kfl+LlwdCo70IDc2FQHiYfOLH8Mx7O1Es59QMlPWYshxqUNU6YTfDyWbBd4Y
QdLLgyeuCGXTUaDxo9EWtgK1oqDEScVN2fEpGNb6NRlj/bdduIRNN8KBqBsW
RZNyQsJFF0jhMHALNqCGrhlxDImMp6doJjpVaZJ+zO9wR6PTnVmEeIpIBsAd
KiUZx8FnAVhErs0g+N5izbiTlwLKHvVp90OFB8vbg+ZKriiGeup8KW3rbXc2
3Lk3KIwyr+8H6sh7HDMyU5A8go8ARTvElU+xSAqbYh/VhLHI8LeDyftI9KE2
n2+Cff8iYzsspipDsaG1tJV60fdWRFo2aFFk2AsaHAYZMsAzJJ1fGNN+2nIU
1RdeF5yHIq/4Kc3Xy9aNTXYIv0nPZyAJOHGIYpQf252M9wxYcfsm31wYlHRy
oxwA9EnR1Czw4al+Tvrd81NGqW3GdRn+Vpdb1yP+Zwdm2Avd5gSCVJNAqMye
eP8NhKv1Ur60Gh6YsVCh04wz/sSjXjon6lRhTONwb5wpdef6Z+grGZ5LmR6e
ad9bwGtzWdYZj6Pcm/I4Mb3XLVOSXfPN+/YUcCiZi3JbPKTlbSPpEvleWf9A
CoTm53EjWpDy1VJu3Cn2mCBkA5jThQnfONZOWTyqgNN2ON1DPja5t3wGdDjK
m2zgOt9cgXwEjGOU9G7+G17z3tDBlsoTrcFSmY4D5Bc9KPCcsWFP8SuKHT6+
Q+ANKFONcQCEAH1NFtWEiEoO4Djfasx45+p1LL03O/hQO8FgRzzz/GRqmmhB
Axc7c9TipU6KVPxjEJaLn39niAEz4S1mqwPbHKkU5P/6q9bcmrrNcf60JK0S
9RC056lTOts2tMWZKDxNrqDSNy0WyowXo67zSvCYu6NC+fBc2/+ODG8UVP7I
iOSXGFWipgYtsVPgVs7DXYwpWRhwrkuOsFfDh+kbZEST1kughuyRgHkiZBeJ
vBBOvgJeBr/SpfsfRniV84KRwGW5iMHYJDX9v6Oyz6J7VR6zVdPD7GiBs89/
XrCrnaym1l3Be4ZGqoAX22UHK3K7eEIAofkIwOzwvOD7U4PwDbR+djafTkWI
0iTSEItX+TVqp23ApXikLhAyk8UAWL+lPNgUlDD6/SDlNF9TtAruyalCUlUo
dU1XZc2/uXvojMAaanojjh66hstWO3AlKRjdZcVeBzA5mX8IeSwWS7Oez0eM
eYRVrxaNRPm4X5zYaaTfZl2MCI+6aexfCqyA+978gmgE8T9BK2eIHnkDml1J
V7zF+4I912qhYXgxyWTJHnuzTO88do0x3AhZYdtXEVmzyeamvuUQBsg3CHr7
dj7iUKXqzvprVeK3egmmvwqmaipQp0oSUHNQIgFb09bEyBDIWxKUYjX0XQT9
TJ0W8oNnM76UryXMEiUbORQ8QR4xjDeEZtVImqLuQLBP9dguBaL5q9xigBO3
94YPcdY36axUF42NDT1cPGsOqbQcWVbV1A9TQ6azngp2sTJ9alPaXVjhH7U+
4+JGTq6WM9TRTG+Mw0e97tXV6rGs69ePipedVfpajz3id9vfGH3FxJwNq3sJ
NF6P2kb8JatIxLmaycy2/BVc7PG+4O5QFADlFPer7/33E6qb+Rfsdp8meH2m
uS6BVaXsql8CgMHff5MA6P7m65uytYoS6+W0/SF5ZUOeKQHIdjRGY4ENkkWC
OkEKpeTvQcR9qSYloi6kbWnlXcI7kBMUYa/xxB8bkzp+gTGWTVRtNFECD92v
fnvnL85uLpPHCJl7r2AGNgds5v341PbhvNZRQs6lbVRQEP+BsTBQUqe+wp0X
fdJZgK6cA85vpKQzrCFO7tTt4kd4sABxWzwnoVljZ6ufPb77lFXoFQFudiuT
a/L+88bBxvYOHEc369BaBjXPw//Us5g/LM9Qxdm9nXzjA2GnLhSrtCNAiYOu
ugfb22U5dXS9CW8jSjCddVLiKPt8BupOkQVFsNEDOOfBNYYDO5PrR29BR5Rd
zuFC9/zZsEjNI3IRoErV6h5bnFB/KwcgKpj9lvwslgv35mjzTj/GKNHj21IF
lpsO3oLggnU2w8nT/m7s94W3lfSvzeVQSKYyp08BPIyt5NzLq+Lz1GOlwncs
2Quj0wvx435h/UAoVB9RXGQiFjpb142K47D528RjCXVqdmKu5Fbnx7spCrAl
dRzrAWMRW4BF8t6BEZCwIOxiDul1hUvbV6/t4eQQ4ykqJxDEiQIgQADS0P7B
MBG9eyDi0q7DHnBoQnErIxMP6X7LrLuFVw8cq9MKawLqIi85wUDqBcXSk/hv
PmU3hLuPIgVwWmf+DMNwXBrPr4WzKZLBDPvjmlm5OiUrvBZ0LHUaeCuyxPN2
fua7uTjVmM2AZuwCgkSH9nE91XSfNzLJ5E3WSLMjkXBB9EYulP49IOV71JY+
MLs9uqNijfeFphiW5sa63ax0fBfzTlXLj18K+jG4GQjUSaDpj3yfSP986Duh
lAZmY0jro+ulwOu+hvp7RvMAL/gzth3KFQPwC/hmKEBzgxkr8Vw70FUJ5CBW
w+PrTmUgBZUjVmmwwolfcj1SVBhXxqwDF7KuHZ9Wsu4VGWcXa/EtfJQ4nqJS
H1/O+TC0H5CTGC4BsuQgJXXDQx/t+NxprX4B1X1wvoqBu0CxT31GR1sE/7DL
rgfqIF8y1GTmrmSV7Ril+HSfKpCVVRVINfEfratPwBVDUiJ4oIt4fABng2jq
gi7OtsIETIPj1x8CbH012azsDhTXaRHIKf4zyZyxFz2USvxpXwJPtCcvoG7U
MLsqKYhmGrKrVGLV8hFPdfsJAVsp22bZ11W98opfdfVlC3Avx3rAg8oMkETe
4qJLShHrSYJgf4n6w3SI7GpRTuh7/irpNhUWSKVNn2gowMt+4JC7BMGuaSoC
92TS0pP5ocdBAaWX/yfSmoHbRYZEZ6L2AhQWA5GW9zLLBPrapLStQsxsJ19C
SCmsp2JlfqEI/cNAbdiRJBiaXMywQL47UFVIa1g/TPk4mZP2mCGZeFP47SNR
sIpOQMSq3QmkC4/SinvaoSXDTvlywn3sb0R0tmeoC4tGGAhCrPsgXsQZs2Ej
87/IvYn6v/vR3kXfMq/sUpDoYkQ6yjQ0iTYLSIEtb8otM/w5qmrze+FvGEAt
aa/2WRhOftv6gZ9pFxQqyW3mD+WbGD9Ya5MONvqmu0MzYWvo2ltZx6AW3Tfr
2St2ONxLqaszRhDMA14l06wA18+Zzl3xAhAavDj5tins4SttJNdJ8QhXRxW3
71a7VdbMQk/MA0PdJtTpdfsKoZgXA4nBCjWvO2gP03nl9qRuOB2H5YjE7DNb
uzv+hiHVELHKbf6oMQgKp6cX11+L+Eab7tKk+TglLXd3Fg40+917Dp1VuoLw
7a3xpr/Hu1gy78lc+ACJLT81k+9jxACeBl/uxmfALqpLgptRjLESRtv5/UI9
s6gLPyHgmOQaG9w6h3/5DUcG2/fcfZscTQNO98op8qtr2E+8REBX7eW1kP47
Y7Y9kFwEhEykq0/HeDNC22uz7TFekxFq3B6hFKpkoNcJy+skbhhd8qGTsf1n
YxWVlcTNqCJPRDcH5l6AeF8RRZLAOUu9/cHjt6cbkqt9LtV9I11I1R4jhY5m
6odgVUBMVTtaSjnh/QQWwgR1Eto9qx0/Ib50yNQApSW6YypSRffFsbEK296i
zYcdv0VKhcJL7hZbN5WPzOvHBpj3g81cyX5PRAK0xXWsm2mtLUW6eiVdZVLd
IL+RhcRUeSHtMjryyksFMX9Y9bmojb+AePxEDaokk22CbmBQ0r1ui5ZLWzw8
Z+/s3ODPgamHWJQzArsrGQ2cJXrw5XUkWEDMH3O9nZ4uP4Unxn1TDz/L6X+S
4jlqYFp+EKDhX/s6YsIhgxsYKS8Du8fXNXLiMmRQqUAxuHCJwhoSxNTGAE3M
VAorFRu8ycjuojqwnoNjDBSxa+y0/YW5bEOMW7iv56o9I87Cnm8qFu2uBX+i
51tTpQRoJlKydtzkSbzgO8yLpb0bBosZBVsTtmOLuFQjKhijop3zO+KrOWMU
ztKflEkq4ObtqMUM5pCnC2uhMqd3n1Qb1hVzaw9yPTv5fNAyOaVSqvQc2wSc
qpDjLDAyifc1y0x6P0csd98Y6IJXvqHXhtetugclzlI9LSUDCA5+r8f8O2O2
eHY9+UwTpJhXbbd1lSMw32wpbPDhX1cCZQL/2teum6Eq/5Tr1ZXIzMjRt4nY
+9pAuMsR2eBXsT/XOAPgD5pOZA7DXYa7IqRbihMhB/ApO663CbKaA8RDhaeR
ZqofxpP9FhsMJ8Fih3x7hLybpDZBnSvXY4ZB+zW1l/pzSoYMV2QH8TyVEHK5
tGBg7X5hpSq+4hYIptd3gXkU7TVZJoSItLT/0lX71wtQoJFQg3RHv47oPelR
uF22zeld6sYklN5l8bjidWep/ihv09JftkDlu38CTpv5duRYs9ZnNbYUxmSW
UjJYwV1nKL8eZTjvJddZNelXhVUCQ0h2R+kObGsETjBt8A6MMmJtmLDNt0qw
wE8V9uJc3PpyllQsGdD8MCRgaW+2XSpNVJWu00xgxu43p0yjwJVi9kj9Ht9S
+hEr20itX/I1e1UebO61+B0Wb2s+TdF0IIW/uEyRIa2S2LiZpiOOYxFvAspR
uG6AhPMDBtu0L18IItRBd+NYhnp78GBMyrXxMKKsTjA08ZoIQ+Rn7+kMNPX6
VWoksJula7lP/dzpe4YKq25v6wIdwwsaNBjXxg9mzNP4x7N1BaX0vzFLpG8o
bbuZpYsYFbIIQTXu3GHqxtLD2NClOytuTofIhONLQTPbL9Zh+4UMjTGA8XUK
vQqEWza013jNpfyqTZtuqEgXpqIY6CjvugO1aQOQiuL9c+qKAh9Avrz97zWn
jd3cwh59pCQNeHC699IOoQLw0qd8Rc/Am2ny5BudDIVosGVHTym7zag/xZCg
7o1lntSmQEk/3yJMgaOCgqu35U+K8r69CyGDG8bzjPAB1iCWGdLu271+43Yp
WHRcMyDoiGokGN7n39MLMH3f7zx9bQ80xKrE0apMboyhVq440+JJzAd1ajEB
h5ACzF8McEcQP5kA3S8yw37SBxToAXeL3D0kgv0f0nx24XTWus3WIyHdWfaz
LufWgPX8WBS3BH8xLmZN8LZlDlhCxm3WEpwegFQWo6dG/742J+o+hY9z5IKp
yDWdh2ESeC/QRx4le2KCCbtGsCMt3gVb6Y5Y/mubggWXSfDrh0O4JS8Dwwl8
JqB4ZfWAYpSP9LOqC1s2MGrvb69ETCeHzob6kp6jIMDCMcdAEGgAYR9ssrGJ
9+az5bCg5Bl9cIEumXJC55vmgjEq/3drd9Wrzg67jJ0eswp6+hGjO9/82sD/
fdZPWfX4PZyU8/GEe3SVpnIMbD2rrZ8oet42sHEhcybaBC0tOB0DXzGUdRpa
yWsqtpP8kh/D+RrLdUuMAcUnrmaspDvrFSQpsKJqeRMEtZXkN2G94lKUBLyO
WA+q91BcvRAGMDWlHYogyKXpsYrSEyHTXHs6OvgVBlIOOa1kLxv3ViN1mg+y
Fdv6ndhiQov27EKukZVlhcmO/gCJowXm+XOMEJh28+hlI2Fwbf5P7jc7D66p
sAX1A4O2FRHWUHkExoySE64xHbzmlGCcCZMo8avXHfUVZwFQID1nlh8SoBI5
VhQltMg0iGKRqU3aJxYWF6f4dBD1YEB/DoTjgh6pyRgFBSvdiYsPH/gDvG1e
YJnN30qISElBwzuUwBdC2iATeZ4bUr/n/6tSCF5b7Jd+mQGBu0OBs0ZoD0UF
dt8qiFcOyGJWDpd+itZqY8IFrTA9UsDV22OFtNKPAaapGLbwGWp5IY7BYtmm
3AghrdeoyyC9gzuxW14Tzaz2rharyyP1ONsS+SUEY/33CzNvFgHf5F+rHHLZ
EDM714Qnb2uBzccScS53mMfqMk/N2Qp6ZxZ0GW6OgTXt8xo2UzaRaXoUiaxS
KK2NuNlP03l39WyrvS31Lw/bPR3bB4OsbFHwKZdgPqyETGR+HfGeVnR3BGEt
hl83GA9Ck4YHa1ZXKovffG2SWV1GIWsG19T1cpH/g6PevMAmBztKjXMqH3Po
PPOexznjar5D4dn4e0jkPUxuS21YVzRrq/CKsUBXexrKuHiA7gZlaccs/xNT
LOxaUa5sx7veOW6RgQBZAVD6EqzlRmlxeW3a6mSKHyt9DNSM99eHLW5qfsGG
BP0Eh138TAqKGu57gLwM0xpYAOWuy/umFMF5ybV6uH0S0gwCKeZOJlRitbHI
AVQ2134i3KrFo1h7CL+ajICiHOPOEMFXKI6+TQwTPjImjOdeqt+ieg8ts22r
hpW7sci7Cc00thq6xU4RFVTFC66AxZURYA67Jr+76fT/S4+qoJ+c+mPCZUfB
dpfSDejEzCfSwaRok4o5MyalCo4N9NVKZ+3aub5PzgElc1yVHBvRCUD/0BIp
LY/RQu/zbcIubh7LSU19ZwKi3mRQ7cOPcGS+MBqHHf7Jo5Mz249Uvjws0KcN
F5wz1pP82sC8cv5JbnWySS1X6eTHKxS+PgLcR8eKmJNCtEOjSap9Dz/nyUzD
Ld8QmdDhkVxjHnPDTrFuttKGiI48CEZQJnVfmWrH1wtlzQVq6/HcZCSBtPQG
iyCcxD34qcHZbmgBbUeqFa3mnJoyMoCPbyt4jeJMetZHOY5sU9fxIwO/7eom
lHq0gDP3y3xWbvgO9dvI8v1sFWHvbmJkkW/t7jJqD8ysOLtteN6EXnY9UOge
22nj4De+3ytZDfH7KlFOlw89j4iQXqmvOmDvEeMuhsqIdqNEZ/oDD+4ld2qa
ttRTvizb5SUFO9zVe+lVZEM6zVcH6yrcaPkpzEngDt525wg9GfWXIq58EY42
S57ijvlIiQEdGh907MaDLEWThxkMzoDUmNSjuIXUyO3VCL7OmlZvrgCXYdms
TfjbfJeabX8UxmKLkZPnnjpZ2m7+ZFEkQpcSiZwT02JhfXrLncqPPSmO2KtQ
EZ3WhVOKqbHg5eeHm9aMn6eahrq0aswJ001IT66V/dUnnnHfz+4oNwjJELcd
AmIuvX+HMB8fr0QwvpPg5em5qjfWbpikmEFc0jEdXW6AnfS6NXVvdB60Fv7b
wIusoc9jwoFdzGZIKD++1gykGOBpPS9vVT9ikfD5dND4JZzWgvyg5Cq5x538
/6UxGEoI8EHiyltPkq9OTaU5LHwmmQVhbRHcTVJzGHF/bTptkAfpqqsExr8/
ihfFUJoexWHjEy9LO+1KhFOYPJaIRDI3QSP+oCr95qANCEVjXIZa8mVhRWyk
RaLJnRQ3r3gzvCZqfDz6ZkQsU+YlL0bMSMxyb0fmqUtmQR23674pIU/id55M
rT/yEdJ/UmKgtjcvmu0Q3XUEZF6fjuUezmd6wGt73Jm7GLtELJYtkKNmhG/h
duA6QRTuiTDNAoBxasfx61/NbTt894x+HVUWNN3lBtsPHKC7VQ6v/zxOakMR
vxJ/IlA3lEWiIYI0Jr6iMsmLu+WICHMnH265KZGNrvUeZvPJQ25ViAnIXTAt
AWPBS8V543lPSMVcfdyB1XcRo1k6/DNH/tLaG+doFF4uo3B9DyqodlqClNEy
KiVlFUQZi3iQ+w2oCHBVWW0hgLnfIywlc9yY7YeflqtDNL0O+Lc9G8qvsr3P
qajmz4OlFPnN6eGcHI8H48kn9VxEaB3g+g8L3JWJiawgai2a6r9dYL7zvbDx
pt7UPAqdbIzcvjIb0VjmF7bFn6DkbEnnJ5C+iSoIXnRN+wYAMooisqnTuUMh
v4dpa6CRiDvwIbJxj82cdzXcEaMgV/TaWw+/ley+dVW8zmhVwboax44AQnm4
T1mV7ZXOpF9MCG3Kz3Buoehm+6gjbU+ka9MiE/p9AQYWO0HHfl51CY+iy1G1
LJ4V1xndy3Xv8vDLSRZuzIbT5ejM3hOwEY7kaAsN9j4S2KXiqVi8PEcB/eY8
sMAEnGlNl4E9JwdGwJt/XZRVp7K+yK2HsrZsoSfPslIRCNk6cNAm+OAa3EbF
eVVxkj6QOO0K+Pc/s/V4wTJuAODbFqcVE0vyC77hmcjCr0JVmfpLa8c5dOUe
7zMO6QaSEeWAbSEWwrO2HKs6Mh6WuwjTSwxASrehq3m2q/27vp7nucmp9mgG
LLj8JWWo0VkVFAZ8RzGt1NJvNhB/nQ96VGozqsXieKvERdfQTPSta71vb6Oz
v4HNkRYfta9hlcrUGyxok4BZojO4Wb63MjTzEWh12VvtFZXcjC6ZYhyizJ7r
sPkHgj+vJvRqATB/oLPygL/va+UQiqrgXB53h0tLTPfNURQNuOIgPQg3byHs
QPB/PI782Ej+cW05ospo3ZcE8rlw7FnstITa27YC4yHV75DNc8a0S5RU09+3
LoxczWbintyjq45f6jFj8LeuuMl9C6Mv3aJVhsus2tXrddHHI0Hrs0Fz5WUg
cKii2QqWt1DFxh9LUDe+c7MqdRLdS7yZUWvvfZu2RHgBjcyRIsduMewqtap5
83BSWaW7iL+c2ehl3uFqyMgMDARvV53xOfcWRPKWsaF7oGchwDCMlzKbghyV
k9HUsUl0f66Ro6xyfUPBcCfNfpQ7dlJCLpWgqa1NoT4zTsEwtcrVNCyY01+I
MVBjVmhHWF/WO7AZSh0gOvQaKTLWohQf8uUwSTFFtbthWE9RzBQbvMGiXiUU
qeME/EFZjTlHv8V7vb9e3i3aU9u2wu8HoWk3bc3LV9XV9Hhcy10tnoD6hZ7Z
gym3BxUWoi17I/dFlOk+MtYDUYhU3if/OjeW7LWdnsv+ncEoJ4Art7VA5m/g
IP3msSyTZs6Wow/IolH9TJLBJp5el0CAw4IQhRLlaBO2MkGSKA36Ypp4VfKc
YLj0Ou2YtYoSsWYD3cLnuHJt7TL+usPOIiptYYGSVQtHDl88VaWsYSz7ELeL
rmAZVU7aTV8kBlTEkEDTXb74RDqyDVgPsSnTMtY/ASOfn7m88ewwF99UIK+o
pcp4pTzdYXWj/sc9oeuechBkhpPr/CRz7KLFgAR00wC77wLCJi709R1XN6Gs
iQJYpFmwKAWrKLNzLz31XPsv6j0EOuXRnp354xS72Z1m8EQwNk09aQRGdRtc
HBxgDHPCp8o5h5J2t4TvKfLVqou1sCUH0pwYM7wscDWv/+4zZjfNlyiYNZxb
EtqpU4nJu7XLb7TbhkSN26kwfXskWNX2PL+M0c4zixFWJvYdoIfuiCXeFvYU
uqB9ltBYPUHoutDs1dc5N2iGyU4AqmBexrzslh8Nrjb0EOF49Z+dxmhxd67k
1FsnU2pkDO/1gcYs2IyYUzarr3eSVMdUbh2Msk2KkCymm5pJ8sjHDQs/LWcH
Tz9+kT9giOCf5372N1wDJc1rU+JMj04I+jDMFyiC/s+gWjYRMIp+irtF96fT
gwSlwsVpW32pgEah8oNNNUfREiejcpqke8i+Yb9DG6V36Vljze+SLxlOk1w5
JAp8PLjDbTlTfgXPCw304Gv02Y+79PHLlbTMFgckYssrK1nMUnZiuH05vEXx
XbA4AT+IC0eE2D+uSXFLMVAOcGmOrqmsptS07oj2ix50+wESRUaIW3vGCtlx
bDp67c8/2oN/AbPUmrtoi6pkKRrMQ5gIHyaVElnWiDYpYUn0r3VsbINUbX+V
07U/UA7u9+jxt1+0wAo7c8SN61SBxrPNo+2tJIurJXvojdz1wvXlDJVmsYby
TSCDzLR+DOttSsVyBWK1ezDGZvro04gR8tXqHWxyJVjvBGYlYU8Gr+esDzyF
dTXa2v49bdNghwGHBrq/W0uKoq9xVz8AfsB2/zAFaHcLFuSU9ywOG5v32Dqm
Kz4AvNI9MEuee5v7qrv9CSbQRUKWkASOJJCkjG8QimTWw6ol2oB5Ls6BYl6y
9/ypngphvJop75vEA59iL2APWIu8BGkYDZJ7gBi/+dqir/A4ADCE2o5Zhh68
LhRPbr0d+h8Kik0XfV8AcGxu/Ona7nhnLfdwZvwMnmTX69CxGtna/sOytEXD
SvKhO4XuPfhEfqC2t0lJSbgi7oqEGc9wy3Xw9Ui//OqcwO8gVPppLMm+Dz90
4ZHQ+Pl9SJ2FPv4gxbp7bk05zS7Ml8RCw1i0ptaZ38SdyIYKrlob9+RpP1LE
8D+XmPmgv6J0469CePLMcbJOLhi5pusfgPzFDWr0/5rwQfZ7AUmC8JlXVLyP
ylyIqrnj6IQnTA9nfHYCSkgU25d/GYnfa41ZLtDfvkRQLZVtQ/PEoGs3VRuu
DvJjE7wF8ZISVMH6nrFQuDmwMInkhyG429jcFPYOkWTlaJXr9KxLhel2B71D
deuWKIITKPSNeG+PghcqtLZYzmuw9XaWCCePLSJin987gQKXTWAAB6QZ/8Pg
PLb5hwp+XQZmbC1vK8o+1Cuwm1ZG4j1e+5zAQb7+7aldKCI0CyBwupUI3dge
P/J9utBscixGu58HLADwe3+bkEFrHbFGuJI/5eGSDAt4iVpmVmGp+EgxzM1k
wUToaS4fI28HLqKSt+qq6HLJuZEtoPokaGiLm6UOSQTNhNfGFBUoTuN1T+nP
QQdJ/EZjJOn1jvCo/P5PWX7hPfZcfMfd3051pvQoyd31EP056sZJgpTbp5Pz
W1/citUnMNPsjgw94UR948MmraxQh9n50TVDVJreDSo7/JIjJNdcCUHjoVeV
NUCa0UicSVYmRfrb/zOMw2WS4SaF5ZsBDTz6OORPq7p+9vvj8luKbC1k5bE3
VMQGy3ZvH0Tx5wM1Is3YaRZhQ+RK8LkAeJjoaqf7ZWkKrpke8F6oOm/2Z+xP
5jG6Z/7p4yvKNpkXQRrG3R6I2Re5Lvb83rngJuG8O6MIPNA+ZDgYZwF8uLX8
vz4VQurvhvg7rZ3dJeDzUvzz3+vpVh+r4gRx73y3p68uwjMvQjQzZCr10fmb
8ioaec3Z0bWPySfpg0+/FjkQWe0LMnqJLzSZpOmS+rVCKtiJ89BL7N7GigLu
ivrQHGkCQLS+dDyv+NEZ/YBBhOqGFBhc8L/tsza1vv0RyqF+azh6T1I28Hwl
yGYMJerUV8xRehN3eKpDJNg55HxJSgtmIkebi2MrQGc9fimq4ViiHYCKZGX7
awlgrZJIBs6MgQUKVYROJWNZai43iAW3vUqoPOwms1hxszA3nNuofxNC5/t6
KR4Y8ftCuoYjeL8NPL8+wNMkeU3ikrlEvmfpYBxjvf6TFxIEnzpNOFEBE2xG
AypqWqGvDE7CeIICdlI5HtEgO9arul+IwlvsvcS1mlj6aTbtX5RUL8vpbYVv
7pkybvcegJglGpss4Ddk2nmmIzF/gQriReALz0Qh2vwLMwC7DiEIJWzosml3
uuUViOrwNDGFaYz5c+cbVuIgixEAwdeN7OYzctggM8SmRaUCSXCjNJWW848F
1mdC/qbScKJJDjeBxRek0u6re7CCPvP6ThepCx3Pptfd2gze/PeVWt0ha26y
yBWnedRqG2OePeP0azcFkhq9mlTw+WsvQPvcn2fQjA1lr6HEsVTtY6pP8xZD
AIm9uCNcIJrm6lHXt7B7UYe+Mmn4hRJZPRSbKOO5zCoRHRiIWuWv1p3SVauI
xrnXxvGyErjOeeZ/LQo6qW5oM8TpQ4cGyyVzbQjj4dcy+HeLEHsA3vhL0qQa
ifgmBciwFrj3eqfvx39ubyDFbUzVLv+VA+fCZZEU8H+La+IMrPevU3jJWttJ
MOuEjtBFcxpDsFG/6esfMxHKzz6wqr9480oufmIOpcxPh445vGmX3dpMmt3A
KPaTVUuEFj5gQrDfVovmrX1Ir0Bw4w5er6Z3Z6b91qJbxNZfwbqNCySq+IZv
GQSPXF8QhwXSru+bIwMhoALvXUCZIg9qX5vCY4YHTronBaH+aFe1ZhSTxIHP
tRrUk6/dKwpGLegDHTiuccUAwNFSfORXiH5Hjesl+dels5EBwPkH8jsRoWFk
tXTHOvItwMMTq9K1fb9xzCxqBvjHizpuE7pKlbNACEH7TfrBdzG0DK9TLqSY
DPfAUVK0q2T1uu9Ttbr8j3CJOxdVKU4cJnPiZJ8cN+p8pMbfjasP3D3dqKQ2
xVuoYb0dSNNCRsFEE0idpNgaw1aPWfWO3FPh5ljb1RH+pFmkhOI1kQOlC8Ag
+gqseFdbLz4aHZKXv1NadgUF5frvLnxrnHUnzvD0iBLfACnoSTGsXb/vLHqL
EtPEAxUEML9tVaKKxRvDaQcIvqwsZsi0Wk5+CpURb3a5KnC9LVznYDI1sBcs
ZWW4xutjxSHMm0wWsb1XLH1CF2GmscJghNjDw1mJpyBllKeFIlIQXHPTUD2K
nP60k4tarR5nNfL3TQa1gXRHOrllLF4l7rwsi+hXZJxyTcAP3NvMHM/tmsNx
/Zki6gX5q5guiJc2T+6HdRwA0BM6INSnVk5px6Fp1l/Qtqatfuc2Xjg6kCtk
KfxiqiuXMyJZCkAjyCd9yY/hqhMyXW++B73SazBFoq1yrXX1sKDX4o1bfhr2
vka+8LPVSgy37oqc13vOQ/TxJKbxB1I4jcwlpmlRkCuO+pdsIlWoxC019qZj
2Zf84bwsZeC+0Ufxd7v12LBiOn+ILOPZmazlyOSKzSKwXMA8zcqdiYSAorFT
Z/ViDjT+V8XHnBv5rJEkY7N8e6Sjf/ouSUqkdKJ+2PL9U6bO89PSvZkL4+PE
epQX4NXWYos970+OnW6z9HC1SEXTibZbXML6i0EwhYKjUDO8shmn0VBv/rIH
rNJxFykT8vpVas4EuIt3oQNb6nHU1ip/luqQXSUU7yGuI3icHu6n1GI5/98e
gB9Eo8cjDdBo1QIbz1ViAzxMDTGgBffdOZw23l1MLf5nHM53LHFX/DjZxAe4
8ufGfnLaD8Xw+Cxu4tPHMZtTPPRst7Hfs3WLZZ5/UcTF2Y3woeasSFuiQ99l
I7Ev6rkpVhPHcKkReTOZcI9+WgtD1rG1i2MjbJy66NJ4RxI0OQGAH0SBeHo6
prnJkeGgp/pvDMu9msrCATpTcI2fnrZ/fxPlBfCjmVNw+MAUM+JRkXFdXzKa
/1ccX8ckRlt7/op7lykqKk7YRrV3z9EttOLe1m4tznwgZAJjhK4U+C2UtKbM
ZAMnGOnvOaYHgjDQrHG5mjF4aNLgDcepESSBS8OVoXH3+1zj0AHTqNeeQYMu
O459ciOV4MXLleVgyv2ul/43aXmCPB7m5saTJohmE7pZufUWMy45kwQTRY8Q
huoA1wH83B1k0hDsb8o7m01Q9H+ra9fXAx9ya7knXsDLcRvnvSWoRPudsbrq
EW4aTQAOXqRoPLZiOfazFIBvD+BJqzyH6jLokn7MxmVqN+cIkR/xH0NIIgK/
z1SWgSSQ65jur1t+X3U66jkJ07IgN9l9KjCrwUuBYqZUYD4fmf18Xz3v72Gf
ciRo+1ZhV48z764GGM751eM7TRwQ09cXq6ibCYQ+PQCZzsiLHZPMsFJp6dnZ
SVlfgFfbAnJKx8XU4spQwjIfK86GNaliE2T8shvt2q6hK8b1OWRFdK8SfNMg
BczxwJa8GdB9YtKv2mzmL97rnf3HOhmmly+tIL7d2zNKDsfgcd1sVwE7q8UN
bEvk9DlLiL1AndR/rroZNtgLSVbZFGqQ+2X7h10jVsE2c033i+xZoWbaFEAp
iXdJkmvRK9D9thRCynS/jOluurtgxXSDYUTX3Af6uQzono9/WMmZWfPiTM8+
VLY9tifTq6SLnXSZ9jZWdv0h1Fif7hDAeNQjJ8CQLTfc/YuhTwDqIGquR5KB
rw8EWnQ+py3AQJg5b5npoYjmJcwVoVBErHk65YyfBHwrQK0Ngxj69fLn86h3
8QoKHaavW58DMsS9GM6ZuUZG1RhuU6yD+hwCpybhB5TwOVL360+U519I/QzV
2brtB8NT3W+vvravtz3SKh0jqzUZZtxIlZzq/2tvpK4LXnZbg3DJVv2AGH5T
0+nzP1RjzW5Uxm96N9C4jdIkV+Md9Y+0JQF+J6LPgwaxiuxTBGED0v5u01Qg
oikEn5qPoMLzAa2ShgaAqeOLjnGmfApbEUsL3OBKwUc0zDnhVhL4rLgELrVN
9a21WfSGgx3ZsYT77+jsczNOWpeDzbXJ54ZlNCb/uUjkiXVpVCLHwIynENnW
VuikDQ/Sg/65faDXFDYSt43KAflM7crvCIlHimhntNToLa7EqlNX2BdOb3DF
wQUC0IWF9oIVqVfNPMunY8DhI58Aefem7thtflKtcA7cuALADoiW8D70aJbT
j9rGAIGY7WBwpwrcERLYatP2Cfos6Kja+v7DPGojf13LY+Tj75N3htMh87VN
ogC/fts09Ryv2b2O2sjzg64csQMujooF/wWf6HJeAuhw/24xgTs9DrXYJgYu
Z+/GXx48wrlaQdEXVN+iBp+mTRKR0ScN9g/vPgHr5Rd+HW8RK2NwtxM30BrB
n8v54f2uUhHgfdh9YBcydwvz6azPBlLueU2Yy6c3AY5UQb0IJIsYYZZq2Uz+
NmQ1x/HHLwcmwUIwfjnw9YiaIWMXY9abG5OWbNVXp08/Crvsm+4K9Sr1v2EQ
dWsmv1pS8a8jxkrbeoPrQS9fTNjZq4s8EiqIX1DdsH6Os9vQyd4e2yODy6C7
omBDDvIZ6x7uxmkTqi2xID1M8V0Vu9DT7FTNnfeKdx1GbqdhlyWyxAZn+3Ty
lAdmpgtY8+LL7m2ItJBclhQW7/bH7x/U0SVdsdyMTL/61gWGEX2rc4n7Es2X
gkNLeT3gG9poY3KMJKs60aumApzyh0jZZ1SrLBuPupWmCS2k62irdx4Cz0DV
Xc0B3cNYJ8ri9WcV2toou+3pTrBbRwJHH3lV7nyTA8mNd3fRRBqdoouzEez+
l6V3WqHzUJtrFsBFXlnZGQS5/pC7wuE+NbieBbic/XhRS7hVPy3KQQQdE3Uz
s7t3KB5Sgd3Es6qYzXmufMy6v5JJQ2LLgFtTMnq2O24gr3yHUCqJ67ajZJqr
r9GNZJ242lgdu2rhycn2pJY97iT3JIzqr9EaaW8Vxt8qOKaYdY4kSO2Dl6Sh
DV+vwJ8njQcgAXUHmhxcWNq9IBCO2XDCEL4Dt+35J/qtzkW2tGWrRlZKpjHf
muXrBjmuyhsJbsy1SrJrLMXmjD78dhv3Olbp+858ZWfT1nbj3iHZdy8gnUoT
iYL7+P49Sy84mkwLTXQrdzxOdd9ItBfOWcHCvMnJn4eB0oCLPex1/1P2XK/p
MQNxdjjfb9UsdEHEgbHYFyFdpE6TfYE3xaxdTGl+HEtSzDaKLURRL2hb0I4g
uN9pqWCz2iAIqpNVAJyJlzl83huCqFI4U9CxQowyteQaKEUrM355gQ6Hkzrx
UPCo6whfUDhV7070SQ+Oru/BOyBCfz6kBhRbETgvGaPEMm5s982KcTCai55X
FlnV99anAlbBXSgFZ5Z853HbpzRXHWMft3/QUTRCk07c8kZ6W3n23JwSaGEd
1O59qra8DMDd1iNEGPBIel4vTAHXDpa3qX/eoShJ+Q0/4RD8yvxDicjL73WW
+Q+ALRlK+Q7aAiBxyv5zEEGm9ouiEQpaKMImsmH4yl50k1eZ8VzlO5vYEBs6
FCeEOzvidl/+1XCsKQDW9Wa71fuaPw7g2pG1pBqHe3YG1hg2vpm9LtqWOg0x
a97EskrgL9piPrxrq6NoXzA5awxqSpWDYnCOUmFRXxZthHPbaOVBs0Zl9wKU
dVHzf4V9hObUDoEhzTroXzYrk0oyIj5iq5InoLb99nlz1iGGwDojaWfKpMc4
QwvtAhezBsYW3gYazylnCMHivvnYsBcdSRSre827HuTKfcHBhga5S8XQLhIr
zpd9C4k2tTJ4X9+yej7RrRcYmSoYwXUEwt5ckUL0ibrBl0IG5vrbO2qP4jsP
awi7SySh7fmXcyc4uGwcQfFh4dYJb/SC97BbMjUCjP5aQ/+cPqvbL7u1/oHp
wZj5xbkeM+kTtVZmC5DWwt2/hnw3UmVO8miosSH9pzDYKsICPQNE2jgkHR/s
oFjOlxU4wq1qV8c/oGfURLrjDRzVDpnunDAhDlKtFceu7IyWxCu1kYu31AhE
tCWQRKfhemejp86l4LFjlO44r5tk7IHMNQdMFmF7V0qjNSTLn2GMWLrBCSzE
3thL7EzwKj4kIeBJl4JYhiPwNW/wrW1CQk8VPSvnLMMvN0HXcwhuGbYysDhu
x4o6H258pHb+G33fDcEDrTaj3uNhxvH3q3E4pZd5NOI0//rqzmhqk2wSLSu7
olzF8kWYfVTj4qo8CJuDzUbABlOTQfP4JkwxUKNFwN+DsAIaWmvS4lbLeeIG
p2Emtz8iTGxssF0RRwQT8SYE031Gp6r1QgSKzepnBGkGIHiFF5nbmf8br+ir
NRSTLBSs9Tk2rEvxBaqiwiL/V0yzyx7pwoepqX+emantmd9kufzAjtEdZxT5
DdBnZgNkygEIbh6/O5EVhOh8fgbpjYe5VkTv9Mrku+eZKie6HSLSmUgx8Ycx
zUyOzUIAPgiJU7ZB64PZfz2l8ZQU8wcE+lP6T8T5dK3JG8vW6NY8VVXi7UTY
mtuhE3Lub8zP7EPIpYz9r+ICnuF7iOSQ0s7K+apTFAQC+VA7xodv3YqBs6Oc
vm0N1hND5XIpQQ5RRxLnOHUFrWOv7HFIi6YCfGeVtYj4T665EZe1E0upKA8N
2uH9gMEwuPlhLdUaBI9sHNCz+cDH0xcow1S2msH6zpiZsEhpiBFETMemsHMS
KOdVEP3c1mgL1WyDlOAv2mMBh7BH6MsR1q5K6ZRHEIQqi59Hr4NgOQUQ/n9C
zYWEp0pLDcL56toG/tmGL1Pt/SwUqdLD9MxS8Rccd4OpNUDS5N7SNRngTtnj
Dd85SaNIbvXlH3wLE1Z9ywWRqzxu/C/XdZgHsAYPMZ9oxEwzP0LvvwyjurNL
5oYcRqkmJZ6NIhUXXzvBxtW3T4+3d2JxT9051K0piklTewH+7Y7Zke+IpCgE
eBZcelthuIl5Bemyae6q8uFlP5rncUuSq/3LmbmlcIyPxbxUAoPvh4oaelBg
ti7jNzacKVYeu9SC/phtm6GqS1v/2592LOZovOpQ5TFkGDsFuriJGQHE6qNi
veCb/q5AVs+d84QokPlXu+dZv0KiNNonTtpIZVqEDvw+JRLmE722SwGOfinN
xKEHBD6BoI4aOEIp+luRgk5nf00QclOFrac8s3e+TFPzQ4SfOQH4m7nFHdqC
9SyfD3njU3m9krpiFPPnS/lkkKniWmB6JapbgnmnwQcjO/n+P7x+0DR4Xblw
RJhhKSjD+U1ICJJCxYE4T8lP23k2sdsJFc+plW/2GP45gt+znra5iDnjwInu
8hoPPivGRj7BIB4nyhUSyW5Tyn33OWJNtULKdAFK8vmJgWNypjASGh2cCQo2
rjJ9rM0aTQ8A7FQb+Boz95zGc9yALRcq0DUYgZB2k9Q6WImy2ZMSJrvakycV
UbyWPMY4Aw2Wff1fWmOulRiGSUL1fN02GgZbS9aybfq8X1KzcSUVgCqzpeIN
ic9gQrfUH/AeI+TdGAQl19kgjI7EERLk5Q8x4Qp1MKkonjsmayfqbSHJzKlK
5Y/oL+duWsqA5HkypGMxZf/5xELRcjMgrbSBWWODX+GTGItgWuvGRbTdJsgr
W/QBSkL3MgGyPCdg6/HnRN4TmP02/ILB5/Dn47CUKnEAOFjc9gOk03bPNOMM
5FGIzjBCRMBhjUky3eOhRfQ9tZDeaUC0oV/Rt/x1NFSiwyb3ZfWBhCZ1qiki
TytLRi29QWGp0NC0MnJI9KK6zW4sMhAfMWM0ui4jPfTiDpdwqYhqqbs8Rugc
60NoezrGCnsZzP+iWXhOaY6yxXY764rNPUFeakwrW+SPEodZjryHjVip7T2e
T3Xi33QJHhnsBv51RNU5oxHQPg39HAHF3w38dL15pHYaVF8YbwXa70hqZZ/3
hCPATWFyXuQb7zWZtic98eVEaVwLk+uw3guXNHQIItp7Eqieiqrd79FP6UHQ
Zvfmx5b18sJeuwRMUIV9OwskCIm2ZE4dl0oQWVX7jC92L9dRSxTQTifvBYTJ
WPRPqJGn4dZ1uImb5vEZ20ik4i/7xPsorfvcg4M9DnOMzcHP8fYnvQmsnC2r
rC5iTX8O/9yz8s3QDBEMxfl1gc5S9eiBWnuNSFyr2LCVMqnXBdzVSWt8URZ7
b6Bm/rjiduoy8/J+ML+As/L2DzCv17PoJ/fsLkojJO0ZN0OrkBe6QH6UzcSk
ZvvQkUKCGOR7hV+bGBnFTXFG2PFBgtvB4Rz30rFRgHYbxqj8Z6FSgpcq5EG+
mSukosaL75iSKLxtmKSK+cFyn5OsysYT8JEPfA7le9BFIwPNrrO7Nq0L/MVF
f0CwLYTucS1geMimDQn2XedMU/bwm14QSK/86j5spZ0J+g2j+jdLaHlMkoBC
aB748M1QaY3un56xX0Ex2C0PYIqK4W9JGp5BUnivvS3lF0K03rek9JwmCDCR
jnVUU/bU7ew8tuyN7RkeLzAjT+LOfqFupUYdWUqJHBCRyguIxx+C01BuTjoG
mFj0SxBPuY6TRrmXQl3ElC1xT5pjQ5t6JRAjaU1UOeZK8TbGAZ8fzOjmCssY
rMf/2Pu3/U9Smc4MQRyGBWR3jQDLhCKoUJMz5W2WGpWJAHJH7hvJ5xaOOc/t
svtehQyxYzcqX38svD9vxnDdjSOKYs4hsmWebBEbjJDmJxaU3lC/iqyaamWp
PztVSnoZ4e3suyxiw0LfElH7czqfclHX8rV4N/xGeYaqJFUD2i/fl6UEYIEQ
rU6kfONdM2Qjfvs2nACIB12dffZ2jonDNPFWFB7G1tDzFlyOQ/3wKEtwBwwp
Z6Xsq4jDRUIYFSIXRgbMBSVBMDsBe/WaqWkr2pZmJO00P7v6b+CC3MshcleV
AdUZaVA1HN9nZXUq5WcnPZxPoTwll9q9KJCfONa+ooWbHooutHSBGj5fVHDb
eZwUdB/Nhz8uCwLNona8RLMfUkRIgGt9ta50E9ma3qirmV6Ruf0FqJ8RR88K
Egx7Fo29gTtJ7ap06wyJ2xLXiue6RDh64fJg9jhdiTqIQX+DefLZtS+RZWa0
OD7p4nTzBSJ+rT7dvp1KbPFo8ZusRasKGwBAdRrAJ5+WDQsnBbBMLVcPtz6c
IsP+gSUVmfNkMsKCpbJy1r6Bt42qPMjF5vZjvtYuK1TqkRK7dRdYn6XGJ195
dgsb4qC5bVQsRrDQZi7cPo0tXbHAOrAA5wb1/Kcalv4DHfL4fHJKPYFrqR3H
nGJl/YWvwJuHANUSRjj0vdP0oA3zlLZjaaGdGatuXthQdMNawIf0XeEQ843C
Iy8F1bgqrqStcDAYZ26dkOmjMeR1i6HxUySpNpYh9ry2J1fncadGcZA1XLa+
r0RPYQl9UNTh4IQmSA9u+Ooj5kDRZi1eM7BZW9MNETD35v22VS3OpQI/VmZi
sENET3uDCbSoAu1BT8bXezIIIDWpt0YY/2ZjSKx+9i5e0N6SHmdQx/q63u5h
47eHM+O763b5PpCqmKbnPQFZNIJanMhw1/s7ejVS7WmiwWA+Ipd9ogi8AJMj
XPhXue5UCeYp6NbIx1fW9VRjv72YCa6CuxpCBifR4qQYpl9p01BxRs+UuNcL
SsVjNb49jlc2gDkZ0is+zTM7vFCisy0eMfhzLvdJ+2Rw3vMSMra7XbVXg/nz
K9oCPqTcElDp4Q3y1YfdE+46fjHs1YC2ga+Z+0VMv0JnzFjGnBTpvJnB9acE
qxWrvKrXwV1pm+hEe7/AVT0oQaaRFJCKG95ubNRcJx46/K4e0HmPvEgkmXu6
CowBThDzILxPTfC0S33ZvcCthIrofUoSOgLKKyCe+eOSl4FxnG8jsEPA59gJ
MApASXEfX2TBBC8mKFMuijwGnJF0E2BxFVoIZ73Vb4A8AIcx8xreK+tuEWNT
m8Y0twDU/eNrqbNJ3kLxDMXvidKrrsvcq6QOCZibIVDiHeA3K4Rxr1MUGhaD
J87eXQuN7xzPxyWphkzlDFvBJ3uhWCvTZmnoT5P/Xz1zntK9srXkssZL8ztB
SVWvhPEdmluraWB7UnR5TnmVdz97MTh/EbWdWw4ocV2OptVU/ufjfljKPCid
J4H8I9Al937N3svDxA+HuUbZJjraUxkT2MseB9uN/jrTjiyqsIzD0HP1NZI1
yWvFl3GPO8vwZEL52Mpe0R1qjNbCDxxFuqjDgtDvV2vTswosvv7sZEGPlWHl
DXfEC+t6UtABKMKozTFJvTjqNMEmNg9Yid9LU/vQ0LKwP0EWJXNMaG7+uC6t
XDLItx+wnHF7jlW5JY7cIlQJSm1TtB1zU/Nizg7MkAaBr3XaGeANTEt2m+ER
gtgv1QdGSyR8l6Xx7wrZtSITssij+icJnqymc4iM/4yzrcZS+qlWhDsDnWHO
LOm9OswpbN5oxJ3VeTZDMugnI06s73m0A8ya60qh7mtpS6y58rAHNikabutB
8dlqVqBie8+e5+vo6fimy60YSKoQobmhbnfPUCuOzjZjcgNLFy1Op59Yhixg
b3vPV9ZaWQ0jIGSPeZwsbb8clyL9pvXng7+WtfaNB3fc3xBDYY4BXLwyzybD
g2A6NtbFmGqwicdCJayRGc3LRblQOa3nen0fZRlCddw2L3UNt9CAXvmO7O9X
lq26wQ5afL8+EHbj42Js2bkp+zIlzY0se7bBv+to9aFbvI9aWWa/KwyIJlqm
K3w9cQBOT8OtYw3QZd2Resjbns1NAVuY0bDC48jo+iwy9jiQxyr3ZDbw578b
DYnCjfUpby8zqRGGSfQSIFxo1/3CLY7WFF7wJ6KoNwG4TVo+bM9cZ0JAdyqR
7NBjQ09s2LKsr+06xIrh2ROzrVDbQgrui+inkWKt1mK+KiOAaS1Z6pqFMTF/
SmWzS4DI9ukC0W6AlNyml1PuSiHvCvByKNP7GuN9QHMTecYreKTlpgNmf6VP
rVNWc5gHdc91Cv9bk/RwiBC3JII10CuYZM8KvDRV5A3gAkCQnHGQ1N+MJTnv
atQDbdCmM0ZjH7UOBbzqStKQv2SPLpTY5nPg/srPUcvMQmc9CWtR9CdLVsRN
BuCyd+a3ly8WSOWShVjfxMnHlwLs5gNZwNvM7KJ9ZIycB96+yD39rFVATlNc
tCJ3VlowHYWjr6fH6VBPYPkSWDpOibgTuprF9AaiMnGhMdRHZqrbpB4KyeKu
D8+Y1GcqOspEdzhm8hVX+FMeSTVOqnecIjCrnOEs02MCfxcaXclvzmtxBd+E
Cx2437m/uD9oB9AD+/26DJ0DBwcJ5WNKZ8afLbkJRxvEiZMbQ1XPW/2Wp7/K
Bmi/nX474CnzH9+2a/zN6RHnptzClmtYpzla9HlpfjCbfyHFobKvZ4vbMa31
Yt8DFuHUVTa6CWPiw3UcnPooE3bWJLVXvmv39o5yFbWwBvtlv7GeLca7E3u8
jsYsdJ4DpxvRFydl4EyrNZ560E1GIv/I8azuK6/wsZPWxyZKbCWBLNXcNnv5
h7Kf8ZhCV5IE4JA0ZPjk2RxRDW8c64IwbLqiLHiF25AqtASR1/O6cRqGntqi
H5gPN+cK0YQc7kwyXOrO3dVI53u06Z8Q+rqw9wteySGjfcKgss1842MjeCab
PSrEFOuw2+YQ6Anblm0yHMa/Nx+KMuGJWFBEzkpDjWQ3BpySQpl8ONC3C/zv
rKBw7rNjLVc7L38pcS1ZPF8WY8DgKocQeF/TBx9poXNnT3Hl0CWKYKFDkT2Q
0FQb8UXIhxl10DBpCd+qS5XIdutUFFutgeXgyKvS4/ZEimdcPJ50ZK/U9Gxh
8i6abu1/mA7i2t9sh5Ky3a+aNv1jD4b9M2NLmOa4crSKpWosfWTUY060Pudu
Dav7CF8fYK49CCwImMiSSoiVE2GRAT731uhq0UBcRJ3jonfp3cRGxvMYd+Tc
Ctw4v+Q4Za0dZGcjK6rmglUbs2fQwh4Rr9yqVxFZaT4CyTdUSybAA3dvLP/h
y8DS31XT9iUBmDRG4f5LtpbqyscaDeCZYU/eHUs4zKmq5oz7bWxC1TsMYAij
AyNv/Bm9d4aFz3PtHYB4LhFcbCsgZ/K7kAywn3Z2LV28dduDmR89B64OAWPe
05bZmRuNkJWsNabV73ZxTrhbhdHT2a4ojiYRWiw1EMzv1qwPO7a1RbudIZQb
TTo9bAJcGFfiGnBDU9hlm55Rl5duFuFH4t26BIGZ243jYi2LElfixk4ETcez
p51OcBXWIl8G6Vj+i9vyR37LLcBqEaEtU6BvAtkd/pO69uxNlLfhApykdPT0
xNryULX97dH//SRdLNqWeXAdTjpy/jT0xlrI26ML2Bn6Ol77jnCI/xt5RVBX
oX//qu8xUhjJmGcYWqj7pP52put8sQ0NrDG6nmC3BW7G9PXQ+sJNi5jElJ9I
kUfgMQJ1hlO8B1mREFxrqH+yBbcjp4n8dyrKM/DMAB16Cu/Ai/zu2OrjCsYH
iGnXWprTni+4r2/EkBAFyp6bkN2tk9/Laf2LyDwXmkFUz/8yW+0zY4UXXobt
ZxBJ/DBakyWcW9VKSPqmeUaXiI8b3jEBwc7U/suPBU8PMPzWDephtceqKblf
v736wwD+UdmBuM5YAyVMeSZBtVyL6yyrbPPGtvKc5/yyMleBn9uK0vO/ftbK
zzpofG+wonzeE8qLzxuhzQXwfSDX98wmlF53IFkH+8c2tkV43+1dSA4Tktix
J7+IDPF4VW5NeSP47KNLVJPlcNOIC8zwbKfyjQ5Ubyt15oU4dkQFajG8ayf0
6RJRwl9A448t6h8NKD0fjL9w2ZGosCT6dru47eXhFKwL5kf05O0BJc6MrbKW
/m6YiID99cFySOZjfMByVdFd9Pwd3g0cBSZdr98p2OkVBZaFFnZgxYDD4XwC
untENP0K4upkh9rk947++bKHKG9fWh9n7tNs5QHoVMxdLm4aXPswVNcsOYIB
WXwvG9vVZnTdLP9Khtu1h3qvwVSfQlfy9gkMkUPjbtewgVofFHBfN9zHkHhL
VCbCLjjOXjccGaC8JixaJ5I41GqDr5IlIw2hrVzCCPKJVe02GxDeyn/LWIpt
zYhwjxA7wzv6QSpB5BkePTW6Ri6Uj7Drmri0sBeysJ+OlG9AdePkwoBb15PU
08DhMq7MuOzpuVIo+ArhxRRktMoLJfjmSFRgWkBczW3Ou6Sw8YUviTdiQuZU
wiNYjy4doJdgbOjbWhQkmpfzGs8Z6oKJbfjmSupB9P4qbZkjs9l1JJ+hGmfL
MRzP+dyBb5kEfKk+ubddywFHdDMd13FjQVJPMYX5RUWkT2D59rVFwXVEpsBl
7ngGIjoTm5Z4H6GndJzVzBkYZj+2g7XLDDJRUU6Zj8VC87K1FqGN253rmFGR
qGf3Nv7/59Uh/RB9vPIi2hqHSqRBw46l8i5B+tEakHpmLmA3WlhNMGXjk4gR
yrlhPwADWWij170yVJOBJGVQI8yI0yKQpnJgq7ncNrYJz1qE/jecg39Q6kdr
szmNWLVTyWzFYVeDXWxkGY//Tgl4GGVvUg3OvFg5024WyF/FsPl+zC2wRSZ1
2I92kAgG5h6icvU9O9E6OCqw9t6VshpFJTRv+vhkNKPZA5cNvG+pyCP6Evmv
aLZ6cG2aQ3r14UVJMvz1L578jlcqUFknrfzPCffBuHIrx5BnNQnULypkrKUK
ziJ4RWgy3ueHQYErti+tvub+SVC7HhmhF989l986vATpwZCFB+77uj2+Db6g
h4iXIpqLikeurPvJgvFd71acm0V8iwdX12mY1QxTgd7pSiPrzA9gPum5/dcQ
hQEK5BQLa6LfB+8VQDBXFSPNv0EeHqeEe5oRwi660n9+3sozL3TFjwUeAa45
g9g5uIfwYVZtz6pFCSl4+nbx6fhEl/GW2OoJGrbx8PRSUX7FzBVWwrc7SIBd
oF5PkuGI6MOJH528U6rBmL/bmAkPuQf8+wsM8Joqu8FmW9I5bhN6XMDyNg/V
LQam1BLMkS98StRtteoq3Xi4zF9XyLuteR9qmJak50kYNzrDWjAGNdHMHyXd
kw/tl3mZM1tLTCu1lgtKdM2IWTO27ud/T+QlixUMWe1valMP3NAO7wmCH/in
Fevl/oJ+UBvlxzlBQnJ/7JasdjevC/Le1l7Z6pxbUlCMhhTobLquZ1LA8sOi
lT/r398yIYxfPmnFw6AnHvKZYDVY1FIXy1GMe4KYBgoEm5/nc1q3+KoYXNYf
SVDSTB5EbHvn8jAsVryEWRufWTA1weDO3c2svxsRba5nbXCOH0j8T0T3TGQE
IVL0BvCHzNgqTcyfDyB3R0DdzT6yG2FsGzvJ2fRxMvVxg4lXdGi/2r21RsYP
vOvShotUdlA7WGKTg7WI9goBlsy28NKLJLSnUTsSohlBs3mJpvxwG2L1HM7L
127DhKOv9t3bEFn9eGw7EUn9zkyuNHLIQH0KHbDbc44KatyrKF7jFUN/ctJc
SEOYmPw1BnKjbEeIrTnDNZpKjDQhuyVgFyEBh0zv77zajc3RThKp1o2O/gPU
ncoQaAZhi3TNmrlbaOOhfv1l97hyVXyu3PxiL5A50KzMepoB8nAxirq9Xixr
U6bk51GMGVzqui7ggRmRrVjlGAgcdDZkGXmGvZenHfmKx+Ej1no4RhTAxOTs
KiuS1X0f0qlRCFJsOYOT4aXM+g6tp7mXvUgzsXt4qRbDZctT5MueqPg6GO/M
RdpGW7jieU+pvq1CzTWqBcWoK0rrWZ7PrR6Zqtxq7J1rtidlfryZxedY3EWR
tzBpJwECCDkUMbGaAiSdIpspIj7lqN+P5DQjqwxTawOe3J/DvaOD+1EIfRwx
JBwLxWoPIjkFwDVTU0Cp3MhdIDrqMJ5UggCBzmN7DhHuM2CI8ulknuK/Lu4S
F+/7DVoWI27F0oQ79AdRETla/+7DTFl5G7PnwK2XEZEFwoyJFl65XLnPxRlF
0rHtzOhCuE6SON6qF2mcj+KckWQkFnh9oF562l4y5200x5X2cM4P73SgWtX/
UKzXaEwHjEtKHWqnOMAgTrWjnqT6M+DbrCuIKxWixXI3cNqFIgl9Yso+az0t
uLHi50UXB+PGO0FAKWBmXMJ8GZeK6xA7WF6984QzEKkjUag0kdx+V4W2KoNk
RY25f2HL2vHZlgeGELvQxXZKVLsPU7ycRBGGxjR+xHPs+LI9gdv82N4N4Ge6
GXtBB25LOF35G9z+w7Z2jgtRvYwJXs4LGfEkBowR2CR5lE+EDQyIAwvRknci
o33TReMLq4tWEL6+QMhQnFG7wKMJNY2cH+1XLBZYfbL0xvR3oVuOG+hCcrH5
PaGXsSIdhGeAS1ZKe0yQHVZyQkcpKLpy/NdD/QlIVquP77Tt7+D4y8uy8JQ9
2T0S14hR7CXRkhWnqVJDFPRy9pIHxluDvq/o7jmZD7jjZOu+4sm1a+pMXMwg
KutE2NHg4BMVK7tQxL8ZsiYRb1ywMxhH5p/VdJ9YwsTjlCXps6spWJynDXa4
w8tttIu+ZlK2upmfzxW/SzuMUtiCW7KuC3Yc62CcdmkmiZQC3sNVdKBg32UO
oQEX+BD/XylBzc8Dsnj/6JIKr3MHhtndROMwqaYI1uAUoJ5cLC5Ke51tg8ad
NzGKDEZsa9Pw4KJqg1G8IOCXK2iu2BGhEAZoMH2ZeBidu0C7ILEjJCEwq8Db
WBzJq3NPDj3m7KQ1N4GTR+aHRYaahy1YURUIh3jnF4c2iaoWxFOLTEFvN+Ky
teOngcPQL2TUVtTCvXtXvQpKVFhQRgSATFsH24DK3CgHU/q3mL0vipNq2Foh
0EmLX7xX34DPxr28rSso5Uquqt5RYBs7V223n0S47EK0mMv3LYDMbh1121iR
WtL2YNwu9WVKGLOsCqkhmc8iKKvG55e0/Q4HINFQKEx9Iy8HyDkiJw+yd/r2
k9gTOR3DCrQGuArmBXH5H39Ov1Is17/Cg4VzdmzqoxzzHnmD1eUHu4JnpOGi
hCgim2WbYqgA10rsEy/7coAl1ifX26cSYYtx2NcWk0OkWsum81EWVzEaJPjR
TrU1audm4cBnU9aJA3CqZZ+YS5a6ws9XOmUqnJY/K0WC+v86yFIWrfgkGFJl
3v4dvlWUZy5NRSHzp+T/RRJNYkx2fJ1slLDf32C5UCNxiYT/QzGwJhqZgTnR
y8qZW1um0temWYJrX5zZjTkNo4oIQojDGaUVwO2UnykruzmeXOwOOeXG0CjS
r2Ne1xyGjouLyENJVrHPUuOM1Y5OXCLCcVyC2FP448+8gzgYzV5gcSRc+6q9
s+iPL7zd0Nu1JhTn/bLzpoem2wE1KAVuI3Cd3cSflr8IAeHOYIP8XrZUrUkh
wdMBIfFHtsWILq0GFzCWMEZpHnbP9tHiggeOTzMnpqvVTAfF9b8m7DHYhdl8
yos8R6OwQXklXzNNz+jEAmXfFvxRX28gH+UIjoJpgp6H/SXrMbgZc8z/+/I3
BNwHLqCHtwT1GIQ3JrgF3g9pz/K1Hyo3W8aHi0hB6VOEUj5g3YCGnYPGK6W/
ndRclnS2yeQX35/doH6eB3PkapOG6Q2WjQGDk4x3gSVPoih36ksD7MmSWDUJ
TPUmt4MkyHZBFBEcinBROSM0Bk+DrWtH6OnWOfPyHxeR4dnbRtI1/diANFbz
xTv5X65wCoaFX9vpzQu9ng1xdvcTAC1OgYRKhLpQJuEDK1vlB8gng9DjYtZ0
zM2mTYsf828A5NkCOqM46qwvUlLO/tPhm54y4ZU6vbMhldxt06iWUryOyq3/
jLsWsLdkJLoImnBYla759xPXC+Un9uyvc5TH8dL39jiJXLWuQtc/Te2RrDxy
hCdznKiCcRd0QS8eJ75vQgiBNQAlEEOaTOTSVWz1kOR8gkM6bMGjHOfACqXH
CEj4oavkxrOclkEB7izCwW/vMZzjJC8i3hG/3ZI+/0EnWFLaMaKRW1EhS0iI
T5oGK+ttg7JyCEUdu6f2mnr7V5syBMkvo3TSLavk8IUb6b2ilhfOVhgdWpa+
HAjN/uXS4s3ECU6fhbvkwecZGLMeK1qn7Ky9bL4bbL0cQEmkF2exPK8VaQds
hieya/VaHKkFYG8QtOwiigx4vz+2t6f5vVdBpo7hDwJlXgUakesBsV+qTqfb
95qabC7PfCWOaraaXvBKrSPqm3GxWtJi66k1CNgCPu1Ke8AEwDShJtMQinHj
ZWkxF7Uy1lBmtsLICE19wzZbLKllg37QHVTCZTpTmpltnTZTTws358BD4LSb
ptf5drHiDE+HpPakFYoTltKmIG1mzP0DF30jV/yBVBlnz2sinYszxieyz/7N
NYUPqq8Fu+E5fgFl23QJkEz3VkmAkCdORX5B4PXYbRZjPDxP7XPTPm4ZFMnt
4LiIDeqlRTTNg+RzxWOf0ZpuWWKTGgxA5cCM9v4i8Kb0lBLHUkTqk1dHBcFn
qPRZAUARNVES337UCzwWnfeDd7qVEY9Rnp8FK4ILO+MgI3ld7K9DJR0/qLVA
Zh/OiWPPV1WqBDea0fC6XBpPBcG3GLB6CTi0OxPNGVlZ3YlYBJaRKgCCOjp8
0swsjbMbYUIXhr2qUbOCYbilp+UCxl0mTtaiFmyJADcjn31Cqf8Fyzf7x64R
3WL2tq/RGylHJK1a8qF8MypUc1jbfdIl6wmUkygy8vHW8R45bkYeIOOftE9+
0Y0On+YbIyH7IvbBJNUQFfm8yWcD7K5CibwNqVdVjKKZKr+s4Zeiz6RCxRJu
gxKNgdF7ZqxuSexj1FB5Lt3yLZH7LfAwEVurkDaErYLLv1WKnXykcdnA72X2
Obv9j3He04aYQyBI6tTQJ3xB54lFfwiSe+ZN2UX4w2KVtcgbEA/G/oRKWu1J
TdS8Z6xKXT5F8pU+h6FKVnqxmBmMXq+2rhYiN4n6JM9inAcnulzOgNVW7Rr/
2R0X7hdykTkfqcdzJ5FnchyP9Ax9YzX7rqOpfrMRV9ayI162wVnsMTj+aSFQ
yzoxv7Cs5lPjvuF+Uk/VK8bdmQ82vAi4A/MN7X7FslbRPwG8PYoiGyUkaEgu
d987JZr3RFQpvCvDGDH7QUnZB6MXiGtAEDA694kHZK5o5vqAaJXokGCF22na
LO3DGUt5qX563s/8NF+DTfQTyDXHqJ4/+uNA5EYB3R3lmv6Ftnd8+6jYVa7u
ep2rmJ+xrkv8j85AgfaKkD1RuLKQotMEU2x4ws8BYaKYLeVmUUXViPYX4pi1
CtX/OXDG3GAXWhmUJL/We838rxI54mHj/EHQVV4e8lqMQ/9gGtDds6qNRN1k
NoLtpot66FycV0/I3wwFVkIHpLb6ZNPUWjSWR8k2denXS7SXeZNbstCwpvgs
Pc0AJ3h6U1mOCPYPHtJwRdmKXAwX5Gqk2imYOKMM1Gbd9QVXsy2C6/NnUwiU
GgBy/bB7v0sMIQnis6pfF5R1jpB/RqbURfuxH/t6qVysDxNPvSMlfQsbrOod
2V9YXNbsuE0/HeK8UVXKV1CMH1TUw6jxW8bwJjZELact0m3ZEM9YZ2bpfSGP
3m5dMNSLoDsX397LVziZcfCzxFjeWlbCz3jS3X5vIQwrT+bF1+zkYikFfKXy
yOe925emzAAzA86m43799+ozzaT7eDoqR9p7XF2z/0G721i9Qo1OjKzKiUyE
ItRvBzOgz6SvqFEHEXHn5NBJWSEhXyjmay7CgI+Z5CdpQDK/ym5a0WugDBt6
pYu2EFTD/n77utL6ffndRa+h1SmAKbkc3QLzL5QYMvg2pJJl3qCU/4cUwT57
Nv1J3vCl6FmoleVw0gCkvhlC6HlBgxz/UBLaNit3eijMCS97Eyv43FYyI352
aVtCnATipdlp2Ah9xHOgty78FQQO6LplcGQEl4i10OMEpNSiiyK/6Gi7ngD3
dDYw9SQaDNSMy4Dwpzn1RIX7SykOLC14FRVw6OSUQkSiIBHmpfJQW4mKWmhP
wlSjQhSlSg0D4IYYmq7DXpWKXrZusKJiDGwp4lmZn+DTJqjq+Nzz2JbE+Fqy
+p0LwjxL7LXFd16V1iztf9D5nPqhsHR7IMu4MdsVqpT6M61p1SeA7iToPOKA
/py3e5qbpQDY2c9i7cR9rnF90i4Pro6MYDR9IVi0shKWpujIvYwgxIo3lGR/
Ht0pa90e0z2FbQpvVsuMBHD++LBR9FWH7UQs8xhSoe4GFWVPOO69Fwy/XDC1
BtLYPMB/vpto4cI5R8+HviVSsgdFpaxcxwbLJ4ds09Df8ABxe7+plScNimqL
ZtIAspZSdtX8KH/yOgsdxMIrFzT4aJQOTsSnnBN7Fv3C0uht8JIXVz66RmtF
GxZDTvEj0hNovDpOSvy4PatJAIZAIJYyy7C2RJHLME4F/AAlUY6bwQeVtA/V
xFaLqjFyGPbHJaldVnK4qBlFSgmlPAIbnR7W4PkvssCi0HIad2FogMFQZ/Sm
YY7L/OgzBfsUbkkv1WVPJJ/eBWvOGMZ1TuRt5UDyDD3HZDtcWYg81izKZ0tE
cbHIjr5BSm5vPQS3jqnqYAgq5wttU0qyn36oY7ZKqkJ2IDceBs/imdOjpyI4
lBquOZNqCNBn9SEqbOs2WLAbrsfD6sPxmBwpFLZTH9l+cCSn5uRDNJrAxLqZ
J3GsxrpVFy+goKJ0IYx8SQQdqma/Ydbdmr5iiOZp+gZuKizJnRb55ZGWLxgr
i8pIU0F4/qRooKfIXe+h59e2pI8qoRL70A0GfyVC3LBRV3ohqYaQ8v9NQqtp
V17qNKQVFqMAiPOQ2NlBQGb+fqRMxaM0IXvgb8Bb3wQgT3ErAyVnZ4enEWCN
PCnnRH6BdUBvaxVIbXRAmbQ0RhGdmwmcWOxM8DW0/bQeXEKHyRp0NdlLoRjb
cCfaeb5Y1Van0pfSa2ewcMcAOQmvAZ3taa/oilZJCMdsLepEMba/0EEVetoj
w3CEwHptvxg5D/9neLdlO+Ld189FvBedQYHwnxgjoFHo3byoRpjYkTb8FB8p
gGy3ubu7HQQ0Q26s8UtNPLPg+4+RvVg1sXfzcLOuATRHWv6b/OU5x+FC2+ZG
+yWgZLnsTgUAhkaoTVOWBessBWitQI87XxrD9CxEzqs61qczGuKUuv7U6EdO
Auxi6/rZrjYpu7H6Hc4iBoF8E0eP53Rgnm+h6wEHo0o9QMphePk8HOJWwNam
MDZSKPJYoJIwiVXrbJMMKQRTuIWuapwuIslKmpJsVHJCGZ36lS97IL21/qkF
DdLNA2uO60htSXZMALIu42BIZb1bfhdB4pNIeG/XNKotnLsqq6ykRhBie41U
TccinY1J8FKyWeAmaVgQUaaCPJMCVrhh2GFYXD227OFmB/+tLWzjIJh+55La
Ylb8BvUCamN3qU0ds+oHbeFY3FbMQINVatpgQW8AYJnuPtkKWwNytu8lTFLq
EGoirkNb5kOhaqF1jJwAZHwNd903f9Zu4YS0KbkaRrTclf22b1HGgBjAjERS
p3zLgErStWPMwYwtk0/vofS3BS9rAIevEQhIVcUj9HqprALzSJ96PRm8bFex
qya5ZVfU7WHmz1fN54fWd0+CfyQc2UOTFGra4iTLfkNyNjsH7DrPKoaclvDC
UzRym16RmYtoVEYxYfpRumqdt7JGk1aCC+6ydH7R3NdwgLehdYozVbfj9QPd
WqLUZzggKj3qmZtjtMdV/Bazcdyv3C3dJCLiMt2IMogeWwMxfnFVLSTGQ1A0
DKqMiMWaV0ypBOw3cILYPRLrmeMzA+HiPjkEInFalSeAZkcVX2sJYjvYJRMM
bQV2ju5ZU9G37RHBTV2ETN8VNh2d5g8ST7h8dVHV4+VdZS6dIC1MaOkfITjC
Z/z/FeYz7Ry1wPNTuoE+p/R0jn/D0g2/ODxjFUczrrXsiNrba7PkOPtpo5Y9
NWRk223GsLSg5726TJitTMeC2iwOCsuO0mmn0/bNE3dr7fUArFex5TEEVneT
CrcPm5EKEZ+mOo5s+oXynl2WgSxnVXoCy3vcz438MUeo6IPP0AF1OQ31FxpJ
kNLoaKNA+7t3lFPHGtIQMd5+hHdJWENT8Nnd/cbWQdZlMezkYPCjNY5vQUjo
P2Ztu8912OnPTNinExuUiFgSDWr9roYlqdPsW1TZTVJgvWFhfMChQVdz9l3g
85dvEmdVtXc6cQ4fV+1Qir/AGwASdibkURHNy9bNhRchli2wcILKSEkxM2v2
bx4wUlRmhWn0xG47FuqMditkv/YjZi8bhpFQWaI4QJJ7jtBWmypHPCQA3UUJ
s4x2mT243CstKltNjHHU35wKPdr2FMHax6nqFr2LJpZB29saKIqNm/nlNii2
k5YOPOZ21vId9Atqxvinq4IRNAAUILqSEqgeOyTcQnjpvChPLbeuMd7Ap5G0
9WZKg5DMkR2cY4SyWJAeZ4EroIRj9eTH3l08wiCRb/+4lg9UCoZdCEkDjr4P
ycxL6WdYR0viUgRiXXqkaXwpuKFqfVq5msiDk2JLLB0C5h5tfH7GXCODNJe6
hxhankw88nlNUIdjogoeBodYD6j/2G8oN/zGCnW9WfN6fGgIh+xiH+e3cMf7
Pda3nzLDQG7rUEePJ+cPnExtg0uHXcC9Gto/fchbHvTuj63o4IfNwR4ZeCv4
B4Vi/69G5yiHdXm7Ff6kRnAggqKCXeNZIEad5I68so5/oN0yKsypP2JBtIlN
ESCxd3Qu/FDw9hjOIyiKZoTZBN7RNX7CpK9t8D7G6Bq/fI/ugcUu/VAUh/gX
pptXauK7UKFhq8/efOH9Zxh2rEzAzHGzvL1DPYE8q4M4ogdAHLOLZu9/P8Bh
rsS4Ja59tzWDv0WVP6esUVeKaJORMERGhCIa7JPoKlfyzeIRbZ/Lq0yO4vG2
ny3iSY43YGrx14R3ljlqWe30wYdbIgEegNiS9pc8prFsCR4YhUqRX6TXdrT0
ct+ATbTSsIX99TQZM//uBgWWPBMX6Gn7+2nHhtvW983zCY+Bx0IM7g2ZRpsU
tYLW5Dt9vH4rY1mxrxKZwOZ4khG93mE3w1u2sNarzwfhGRFJD3LhvY+WBCUQ
sPw0FJBZcFvX3p9icUie1+zrEIPo6bT+2mWXWylHyo3ZDOzSaXGHK3fPTSdj
4DBF0Z+MsAaNcm73/jEseuNhhmdTJnaJ1VYbAMPK0XQUwZ3fztktI88JadKN
+E0egMGNKvohbM2zWZuclz8uiuISney8VYtpYRleRzmMHw8f04SvArQOT4bq
6QjuGOCkJzfFeyEz6axJQ8y87ayq2Idnj8+faAFPYyYu68A2q5Dt4zff0rOk
FrqELAzVF9RdqQyDoi7DpA/XRFueKbfghJcZtgkXqhH/0AaTpvPT1Gw5AwpV
mOKd+IbSZyrXpHdQTJlhE+sv1KJ9ppIOI6Mmo0DBWeKCx2NJgBlppt4OdPdW
P67Hml73NMa3kLx3W2LPev+LImmcfQw7SnVElPQnOFWZhGCIiChq1Rm3ZjPV
MEryzSK5x60uYLG2U2nz/+XdusRqXibu3GXJv/cofblPhKBA82POG4cgoy6q
wZrJgtGhuJKxOvqJDNmB1MsGfwz+97FeVGHYB+CFfRa1LN5275HT4yZaA6ZI
thZjb4UDbU8+jbMZb9YX0vdk+oGHau/z6tW7SOJ5L82hrbH1wLV0n8WkV3nB
FM/8VTOoEeSfWNphwbrgSAXf43JjMskS7qdYT/72M75jmh1EtV/HaTYWwsN9
ons9mwTSizrDr4OK465ys1S+mEtVf803oJc+wU7d5SE0w4UZ+kZ8Ul+z73L2
9NksSgG7nmokJ9mK0xFD3BqJ1U13WEQ9IY8NH97opbXcEte8uSQSvJfaswNl
B2j7CSqPYRFM3W+kdo/y1o3mp7wTox9gsvWUURJbzaeIQFG0erl6F+eXRZ9k
FCmenS/aimJ/pR5I8V7gL08muN+vVCGfSMhSKB4waQs+osVWPrIZmpS+w54P
RQXnwYRFbyL34rxogx2xj5kHDgzQkKJU6PSaHQ8i4+E5FDNquHuWytJOpyp5
iERsElPqhOqG+u1M93TNzlT63wXbE6lkKEoWI67rO8Xegily4hMrb6JtTxCo
3VggU083JvJlQmH+lYUKgKZ3dR9rL1W203RKM8DsPvcvCgoI8fAw46pJtiEn
esGNFcUOeE8pj7Rg6vTYXX64gIL2OqmjzR8KPpmgNycOdn/Hvi0PrymxWaC9
1UDx8sWIAN8Cr9GtBCpRaz0RvyIRV38HovtVOQhseH19y7v9U6wveIsRajfX
X6U+UXkc6al3CMAg9+6mv2YhI+Gx7s4B1gSYlTLCg4s25glkZd34MQubiDPQ
mwFvq3/6cJA/CPO6nZmvgNaJ3GtxlaPu9QVNsgMHVbFXaKdWUcPYbNoIeFQ/
m97g1I/aEbxukWI6EZrUpz4TfN9539xqOMRmC3mfTmdLvyEiCjmWXbTeJSGF
eAas01vwE6D3iWoX3DKDB1CmtovyyaGYmFsYiqTAm467cP9VrYAP9kebqPrn
hkCC1BoyLO/3SeHMeHL8qzG0u0Fa9A17VdIL1At9DYXVGD18D6JITkFFf2hz
Ujf5nvQ/UXHi8EbGWYIlrON8w2JuruXS7w/UDBrIYQjOwrV1wCKmPPS5XEwq
GKYNADm1bSnDaeAXmSc4zs4yQAx3XfBR3b84MISsDTLd7cFGWfy4HZ3nfPvY
UT8Qo+SSUh+LSrDeFphjgClQ+fKmNVN/MxEZ5e8SfCgvPt6Xsy2M8sVxZQUK
20R3kYUgE1qrM2U0Hy00w+HF/iTbuOD/7D+IamCznjma1jnVwQ4XVyFuSCHt
JWMdsANALpiPQqNBtskLHBzVrHzBwVo+qgBivToMzfhfXroLX4jz/WuURsEZ
iHcFijRR3Kiw33MmJ0+N2KdJ8i90VIV5mE/mYzEa8+7MSJ0oBGp1ElnzSA2p
u/2PGYka2CTufFpGU2REf+1IA6bk/KWt+mELprMLCwbDItUf7i05dDqC2JQl
u841D86Eb+Ic1tTszrC3WZ5FPGIXbSllfScvJXxVtInsSUNQeOHC7tRruoYa
Z7+UgfF9RjeDpyV9mTZns184KgQwj3GS4XGJw1Dj0JbqwjJTD+jG0lUaeA4o
2InbFDLrZmRiFfrnCNA0qDjdrMujP1V8PapqFExIvudN60WO/5BbIikWysO+
xMkomODN6R2aHKrzbX66NOOGI61p4/R+NJw8AjedyD+culmHA94nB4hagjPF
zHeIppkQhajbIP2tt1cKV00Eo+q67nZrbEmuSNszrPZ2S7/JnIs+QCgyETjx
bHqqF+LwlTqiMjlzA2Bg2FkLSFJYCPHhgfz6WuCpjVwO+lEW9zLX8QiDZUWR
+4vMWcLe7d8hbJt0hfqs5trSf46N+Indtq3JQ+xGvLMgjyInnvKdLCF/kgte
KVmEMNq0wshqn3TkUVLobli+mOW/ww2E45rpT3dFT/7j1Jk9TGNjBDaaSOhM
WasxyG4UGvhs0pEkN0DWsDAnyEDQLnhbjk+fE95/4Apgb0Gug0a02AfAFrZc
7BMYBk+qQy7HsMAYKZfSUEMKmY3Xr7SSBa6D5YHo+JPMoarh7/JbhPkxx1ry
Yaa5hnwmzKbT/GxXozgdGINxfcUzNokTU2LhqfUJXrw+H6fCgNU/y2jkShW/
J+i+4Fn1lV/BND9TfTUUE3bDbPqDcjG91Xu3gbjlSFfYiAEUOZ+KwXTmaJoC
Ce4t3ik5zQ1queCEXhem/fPTFWg740ADm43FS6Fy0a1BSZOrOahiS1T6gCV/
X0QenBKx/tpHaM+An+ouahnoIvlh1rIyrncgIRksB9DQh74tncZnExSt56pg
Comw5HTAyGF6JBuVM+iiBSXssMSQ8cPIZSH6uxkF45BPP/5G7RkokslJgLQ9
rFo3OQHrSndbR5N+uXj8hM2/d3NrJ3h5b1u7tLM0/9J+ezvcvx2odxH1bmAa
fAZolM7ctX09TiamCq0aDf8fyjvZd2fRiki2gGDo7/O7BwuVuQaNfM6KnHbo
ryXv7LWJwEruUhbg19rI1/QY26+Ca/PmZS2satNUlTbJmNa1q7/HhBN0txXV
QMVLCxkr+lPLMzMw+lv4DhGsUALba1K0pGrBjRBtWEYBjJTDm5FEUSg8hr4U
Xy5INRTP4nVTBL8rtSBuYf97RLaLUcK4VvEeDw9aOJ/4exlrPCL2jq4EBGRL
P+zRAjq0nlueJuc/YncjA+4Jk9Za8CKw//lT1DyWci/LDVKgZ/JajZBdvsuW
OXpGHK34Z2ZKtanari7BTZXg5TCZ5wMkxRN9dxFQ7rWCvy+wNpJt3o+pVYiR
xSyNiyMWFxHvhZEVtFLiUs5kMo8/ONvHppqeV68KqvMgZZucoIcmQxyzZMvc
jiT0YcTKFT2AxxJRKVNHK3DJ3CPtxkLdl1DYlzVgVbTyP3NEllKi38Tankw4
7+iBAWlv9ULjRUTTyDGNi+5wCVq3Vrp5nXU6xM8KVAEgNRT3ZR9dnZMwfIVp
m/Q7ivXrCsm5OoNwQyHebjSQG24oZkigos1hZdJKB+jVt3elP8pU/UN5QGqQ
Z8flghObl/qZX36MGF2XPT8aZt3kAMiIKto5QKsBVtGTfiqadhbtOBj++I4E
LWvbi7TYT95j5ZxbyRkK20+2rYYtIWKkLHr1JIBlFOCkXPgo9w4uTTpvryRB
27a0QGGY7peXfg2ZdFZutsyX0Kpsix9jfHQE7JfawkFk9HHWJDfhBFwVl8BP
Pzgot+4tmCaFrefCfI4BvTxSFdZ6771H2D2A9MK4/cne7IPFCc4Wz8DbSvtr
9423JRanGYP7BR5M0Nt8DBDwVHVDqCjRkzXLwn9LcnJG/0ft8u2Vjqt3f7V7
ZSpUaofO0HV2pYUXrgQIjdE7XoCTxpCLN76EvbQCWwPbFUsMBnVYIFhhCcvg
mXiD7MNdvl3Qbc4ONmqBO5tkAW660W9DSc6wVTmsMcCMpUI51xWWw6wDFIAJ
k9RIVpMyGmPGWTf7wVHIzpBwd7wu8tSwk2KNEGyTUi3nNAeduTYv9SN0GWbr
PCad8aFDArMCeXawsfxiopEpCoOM8yfHSm4auSqdNEAHXE7iDcb9AQDIEl+i
RWgR1eIM2DlbFwB6sVVtMRcuVc5HSE3cIu7fpD5SnhNn1wFWdJrtWTY042fC
LyycIQdlne6hjcCC573jsCYVGA/aXLdnJ9LZptZJd//QaGqbFLJSyc2i88yP
KnQjasIvguxDjsV5wRx/QNhxLJhk43flTthBwK26fIhJyVmt3Mnltda4LtK/
lRfWcShNM+yXTgUxn+M1qTHRGCxrvxTwulaOS6FNv77SMTPDUILVB/XWBDh/
0Os82tDUbD9HxJhQ/wIk626YeCN6xZApA4P15vw/Ct1zy2Gteq1YSF96nByE
zJ4X5mu+yxIWUbuxVHP64aMgQevC4mCq+M+A3ZNneeqqLXlK8GfHZyeNr+VQ
G4OlwWYEtfcBjFm1u0IdyTvdmfyL05itCQH9kcStXdhm4YPTSfPPz1hqbxz9
xsrxi+eetQ4NIwNvPyjAXaf4n1g6SJg7F4AtBWTmJbKs0/lPoW1Ye35bBL3y
Gz8KsCNyyN6f7sqWThHh/7PhzkCIjl8TY7etwIfWFZIuoF/XQxFfrPeqIzPq
77xFL5XIK6s9x+xYUdwXNtQzuH122Sc4XyLuG2sRZuXMhFgzXdylz9XvvXLR
8epW/DPzYydcz4F3IAWjI9F2RG7bs8Q4cXedD2O5UQZGOud3+li6zsnlpmzp
55nd5O/XxLr7ZT/mKo0ysG62LL6AS3ZnsEnvRCMWyIEpndmh9sxqhzgzq07v
t3Eyk2It/MUoWYoSES3duaPC2YlfWYgD6+wN/gb1/xL4RIdk9kv3VLKmMI/z
C6hkQTzriU8wIq7aoIxHS5UYcSOcSKguPj1THNT0GCqYqXNVBvMRlPZNaboV
YuteVVgMOkrNhe7TOZfm62z2OokD2d6iqjpFmJoDTKs7zhx7/RWY69lFLCe6
pg8t/O5tqFupo6OtyA2MArPUAbSSONpViN/r/pm9iGcE6R+ONQE3LB6dELKv
eFElV7fLbmceapK08qalf/9jNESXXWoA6ZY9H3bXp4+o1QHKgRc3GXUEEusm
n4q3BkHZlFxEySPgrkB+caItp5oeLRSl9ssVR9CRe8WueBrUVXS5q2ef8kWy
sI0wgTKMQMKAF7hT/pnvRvvIns09xArS/eV+McetX+NS+ObRT6BM+1cFGiMD
CGBszYG2bUFMGy2cl6uhXMzSHefv3+IKvy4LvhJtWK2s+eTdiUSX2drRRwLz
N4m/5xTZC5oWkTezhkjs2odzeQPTHXODbIaUWUT/FUDz86vv6ODfkdFsMpZX
/dG6KtRY4Uqe4+yQVN8dRCYVOTBNq4aH5VJMekHReXu8dwwpbO58o3OejH6Q
4g6TSoSbC62eKCjy4pQPWlQqYT+GUkynPvaKkFCRocpylflN4CLGbfYF31ve
LbAuTzN5xYFsZElvjPme41TrGKJg4cVX2MfPc4ibssfbhyzkSufLRavXRVJf
qPDrpwxPxfzd/t7pZ5dV4RC+OkhL1h/2LXlf0j3iP0D6D44h+LMIBpNmMtxM
zukI8knBRujQpfiHOLCOeJDvd+i0BPxBGdU845SXB+eFcZTEGM5PpLHxddS5
VehYjcuqYUnbOzV3cXu964m6+xxZwtSIkYaLNnUBiIN6eudseYv+7rIorqmB
ClEggC82br6mOoC7b0QkfRtnJjwtaqSCMfkG5y77gsB0/MVeXNvBI4ItGb3L
DpjNUpTI2SqlFbDcRjjK4nWlHDg0nziWWzgjo06XfHfpXxW47GZTB/frUROp
AIRJrZVS1eFWP6AifErH+PyTkN9hZVmT9UeRbZS+BBfuShbjjHq1dVK34vgs
7F2vBvB1+zSAw/SbO86XlB7BZwtQ954+GGAPHqHINEhMsxRZCHswIzglMxMF
vIZOzzhIn3Q2F1wFk6Nt0GYEWAfvhuOQCeM7u0NmuWdI2OBeE0rooJW0Qnoi
2A+FByd+Tbxnkq6P7ut+1bmyvUDIIgDKs/idBepF1Xlw9wnK+7oyJ5BP9p4R
R+SAAboX4QS+v3PC/e/lijTPilC5lhwHIgzpLs+5x0G2aazKuosAux5e9Nh9
ARASL/XIk8PUTvxzFSiMcPaJYGUnVO0sUpTUf/Rvf5CO886oez0bZPDkjca3
kM3gBIJCiTzRGiyJwtMGQM7aTLyR0keE9zTB2Ki0ajzwMSW8E11b7T1RYSKt
K6lRyN7dYUmddSoA4WJVGMyodQi3lmbykM3zznWAa3Vp0/qpwjMk2CpuP6YV
3UoD/u69eChlBJ75E40B4tDyR7KaFtQTVd9+uR1JbeR8v6iGihuyZ6NzwXt9
Ru3/NfzTPTOvDJKYaEBOtI4yCrsbFskOIskOThhM+7Xg+hKPucFepk3d+rzr
iGs6USeVH1GFCn4B57Cde7ZTMKmNioZhicYiZrYA/daCurEqc0tFBnmHSVjl
caYXa+aZjzaxJhod7Hy7bdy2azSOiYfQzwcH8mogehn2Qb+jwhhhSJVr8fjX
6qI4VZox7WYwhL+LXLw943+QD2p0tV0bSo91pcwLb7WLKxpG5km4p6gxj3eM
pUp631J/cnMEUh9AjcfQh3YuOpSZtvPxOc7p9Cn1r08BLN/NXwGoKvCxQyfP
Wl2i+XNkPLkk4Muyn3se84iX8cCl+zAW7xeaa5fGmiAh/uLnheC2dmDHEq6V
H60I2/TRr+K+6FAhPZGhgXT+jeaV3I7cFc8cAmipxPcItobDVDIRpPBUOL4Z
8vGSlAM5gSY8h5bUbjxZKt+IpcT7I3isRfZZd2d/RRSSTGXbolZQndkO6EWW
9Rr6BzgwdcJ/wSDuk/bJaCSP/Fcdg9KeNDpg+6IDe3CMoQXzYn6pUNrkDSir
oOb91n87upemZ4kJevX2HMFYxmIIxr3MzC1WDcz3e+Jnrka/INkyVBQ3ZVbg
J4oTIDO46FkrkYdAi56UQ7p10wy9m10OspTFLbXz1nV2mbpc59dNeeDjMgye
UGdg88zg4X2HzwUlQVqVT3XntJ7JafNEHXOt1rf3BOVq2YTUO9eWcQ5uP2eh
1IXbL06+goQ/tzJH9khyq9/a/GLSini9ut8y70OCQ6Tp1KQT2YyYFoxuZMf5
YBEvLjCuVHKzZny7Qkf9neKrGxifRTPLFOt2jWv37VexFVi3paChylgO96GP
aBTelsoDd5uWzi0H3ZvBExSLH2XTidh603ooM52Cx6fuy016WbqwrpNSXJZk
0SXbgIVF9lKLdrWhNcgJb1yUnqf+7GSdNv++qWq5pCTxqH3dWilj2AWUcuH0
B4YV8EDURsOMY+k4b0bGiuk/D0+4fD2f6IplMsS+rRyXcM1ZLAC27qsN//8V
pAMyrly0Nxte+wlefWOA+uYbT/HYxoTPGXcrd69MJhhAaM+O2EyTRldKAknm
Pj69B27he8Q335qHyMTCVumd3l4kkwvO7C4gAo4mAzl1ySpAjYFt/GLf6GK9
sijSrgg2EStAYajfocKHnf0yQC+8Wftt+cpd77OUv2oI+LnehPHuY1EC750U
ZFd4vuTc+pa3gc1QFkd1qePJxx8QCb3Zc4JmZwm+w1XSIMXsRQxKgXuZdmi0
a2xqk6dc+lO/RdegVO7Rh6gM37LlCAljWiqS4jJEOF7Y4qIthl3AKJmzywrT
7aATeOVl875ZuJo15OmqVv32Q3+NjSS/TAm2hVHOV2aLsKVh1CN4HJH1QZ5y
oT6cA4ysb7s2NVZCNe9N7a08C95nfnqsldtVimhCg81GvBLLjGxpFxt1f/6T
+3GS71MVlrZ97j6uKodDa/q5NjIu+oMiYdGcnPGVGWpej0v9Rz8KY5QzafWV
GPx3mfsBUuDxCHdWp8J52qRYyZlqUQCqsxIzJuZ81fuFtvSLteRDvwobJ5Y7
ISKKC9zv3d05EK7fEFEaepJL8MZ1H20GuHRKwn3wNc8he1JqtN2vCT8AOEzf
ievBB+bbOu9I+MtEnb6tSvojvcMhx5QlXRPnD1jAJQp79s3TtE9NLt7ijOeq
JOa93Y2qRRkXjoEAbNIzWBSQzvmCstiE1t5mW3NZe5Ihf4+Z22eE4rXTyA8J
c/LgeK3DfB4qfSE80+SWQ/8epyVVOL+wDmYavdRvcyoCQhuLVhxVGlC7xzwm
/oOnUKM/8lKpH5ZN1zfiwDfNdkj7/S6QGllzRTKqn4bAI4jTIjspf/82Y7IE
ChS32FmharYrWhzxgY6neGYl9Wvgqht3S/dp4SIbRX7WQ8AT4mUz9qKJ7prq
h83lyHGyGETU0c/aDQ2TNsm3Y/2o8mAtS1DCDM0FucKb2nvaiKUpDfVH6iIZ
ynh66kXpSIMVjc1wqYdRomObCrS5POmKdWDuZqgmmRbIQ7aTlXxtrge3TcW2
/AbTCd5Bd0coD/PkGi75zGifAFkySf5pkLWef5IwyFEzNgeDOohFdM30DpGw
1fXrLxB43/XO1BjPQdy51pFGWixy+gq+TOKJCFRqBVObS19+L9bRrZP4IumW
pTl1YXdjFuJ1wKGZbC9cMGXsV03GLoHqDGdz5mdUsxuWXcc1B1AJhuDeMt88
lY+3/1Pz9DXDKDLSZAR42l98Mit8L66Q3mlNItiUTXkCLF0XiBEcdScZ16A+
6/1wjuCVovKFzro2aFZaAFW2LlGgrn1r/JIfhqvfFNRdr86x9OUVDv8ubHBj
fGiUpP8NewRZFohZEv52X2U0ULN4fhopYnhHAkwhYP0ydX4+OM19Cu62SsP+
BT3pg0h0WryX3/yseAruIeGm7aDRITQPtM9jnv1tCfEQUF9I2LXsZUUD2FwC
6qUNd6eEfcPQaDxSU3weFcMBXGc0HtinJM0KoILOel0fpv+PRYHLtmpmQUjf
kTaEsW/KdZstocriHQXLaY7iFsEnGrybalskqLgOZhZtnIJTy56HVQUsZQyX
vKY1aYq+4H+HvLwBxiGO8GdSS0bfTlkLWaJcZR8pwpf0CesEjqvyv9SfkRfn
2vKL9np2gEJ7fU5EFt8MowuCmGBJvCyAV3tr73K+yjUvLvhrI2xRnQdzdxYi
Shkj82PCxKX3n5HwcJK1lIco/pF541D6qzPVwUaJvxmrtppidmt1gBR1TUSz
l8l+xjwF1jNDY82LLiaqwQiHl5TbP16QLX2Obj0PXqWl5y1OoGeuHuHY9oNv
4IOUhWIeXElvbZdAJc+w777gAdoaNHGAPnNkq/s7oIBAAkQimCnp1uVHPHx6
HoJ6xTZ8LMZzKZAF0HSmiOemzlvC/An2d+t0dibSKTCmkesYX8g/6KOSjWf8
nyOeyajw8SQhOlxSoY3xwqjklRKQU5GnePNBcJiRNxmGFtlMp2lcZsNrWgXv
fnOU893EFWOxkw5q+f4kWJ+6PfEWkxZw9oScGYnZZ1BOihhtKO7D95KMeu5X
rK6kAvRFElKPYftOorB/YyfjMXnhRWCjBHIY6XGIGHSm+KmlAKp+a6BEXhl6
3ueyElm8UuUdHPK0Qym2vunyyffsgrS6xmJ+21BZI5fLAKnaToOg2QJXjMBX
mBwM1InF1YY9y0CAMe5BRMijF+eEkaIY7K4aIcYd56/pPYWk8/+qyhd6o+L7
UHm7ud/pD8/M7NxTgOCR8CJAmElCSbh1m+CYsyt760JxBsEK99Hh4KPCL4jk
4yrORPMUa24l1tO9A1MzJk1G3TRTY3YFZn+PJ31mNrP+VsQ4ABKxjwE+F+oS
yCELbVdDMh2eyML5HIcDKn8xjXvuphbrM5vKwpt6PAWnPxG2XMc2CKHBmNGP
8ln3kO9EUr4AQk4uyS40MTB/BiDK1NWIiWTnaO+iiGeTm9GvwBSCkRGEhmcJ
3Blc9gEbb/5OsW4+MX5NXRyuU5hvp++mr3Nrz+t33lCOZO7ehBVMBzWGOSZD
1SZjhTI5CseePMWbwoBDYTB5L9Z4O9zn7l/Khp8w+KMr8PMxfGUjYv0qNuMy
3prQ6Se88WQtH+I/p2ZXjSMmvK8bi2oG7Kqq5/BnEEMiDNnlpuZ/I+d9h+P3
BE1+4pokOOGJxnYmdw5xw7k3Whw4ogWdLsHB7CUrvBhlMODPCsugZM9vl4lH
pKgwsdZ3AUcynwnAVY/HjaY7GXKdqQQbIpZzNW85RvI+r6gHqQC+FaM1FU1+
NFxwJsor063HNCdq9gdgegr6akO0W0p+Xrbrv2SiKhTwqXSjg1ofYnpU7cs1
dvKe81xvRcIQaACzN+rl1QN8l07u7/kvmiWBuqaNrjSm3uuuLs3lY6XLH/N9
GOR1GVqdjN1g6KiPqSmtaAIhi93c+luwkYFn9Dy2zpy5uJb7R2xY8xIzxTzP
XHBKub9ALukgJ+9PB7/KthXupBn5bDwQ4kTAWkMP9aoglDhKCrRLEa96JTMk
O39T479STnygI1t2ZclmoYH5EOsMz4KiuoQrq7z2uuJixc5rY3wNHX0HFeZu
KtZ6HZ0KU0R1C14Vu8EgoNLehehdCHDugk+WwTyEXHD1WbwIVojY5sWmYgZ8
evbvOn1V/MXT02mslCnQzKoxAU5zv3CqBisS3Xt8mO6h3PEEAteV2gl+oBya
OOsLCmPloTxvLKbvO4rCm//BUyojp9xUDMskStKWKlnEfjuCmeYA1VyDMSOF
E35CCzITB142XjM0RjMWSHI+NTRku/uTvAWc613Sh+ovxUhbLRVvu9q1rd+n
QhVP9I4KFylGfleYcstkcIG/IO7GcPMF/nahuDLbgDgbMj/pOXRJljAmvB1h
MPY/MzEDrSDk3xrf4cfRZigdmy2dsjwl7jdS48brneVLjHITEnH65b/diEug
7TDMJ+kUQ75Iqu7kwyINVhWlQfpsOPr6EwEFDAHsOwWPPhQAm3jtUGzsnuxO
B7KhBhBoTFEwDfXnwTiLVaR0U/qruqLfAbyRK4vpbv2TPhSV41Vg0FkSFN8Q
KedCqyI+R536ZIR31n3NfnnCK/ABeo6T6ImSTGxB3IdQ27+KVQRe4qh85goq
MvBGcbV0/z3Wm7fvID5iNJtSk+VUDCB755CtEDvgjdKSTp/K4Xwe0blo63z3
/tU8mSZg8DD8boaHJweQDV9LEh+pNcXA/lM8j4e+L5R8rNT1TXRBD0ROxR12
GUHn8dZI/NEkxZJYgZdz794YQxKJApmJbo8KAH6HwI1YLsTZY8nRu4dHbpVQ
dks9Q/LxFQwp5iqF0+G2fScyQ0ofnNL/4NPDPE83BwTibFy5VxoISlc8QVnN
5dLDBbE/nSwTy1Q+RoNV8rlM8juEHf0ynuLUDMWvo9EdqjQPdOKk/F5MRth1
Cb/0Pr9TtchIZymbJ/bYwE55LQA8vviRO6+04DkpqUqJRMl72xHyM6KFgc7X
IChFmEmHVJK+/wdc6n6bsMSob4YWLGPYH3nxGBsvPNRDdgqx2WyMB54EOFwq
5qHvjAGcwm+k7iW3PsiJtarbrHJkyrqDZ98bcAvY3VjBFBtHbkleCsyWCm1e
qN/4g4AHBhVOhJk4imMrcszd0KzjJmMuHjFZ+EorQnwvWmONgbhcYyi+ePo5
CGpqZugdBw47/R+rhLL9xGuto4voZDdCDdoXqFepDFKqqVZeRnJ5FFeII9yw
gzu+Q04NG0BkDMyOgHITok8IFCQ076ZqLsF61bTx5Kb7Bx7TsY5thTaQrEcW
pxYJihpxJoLlMv+itSVOKijdP8ByzXHhiabCvVCLmLIB5GvIjyGfM7kx34Dc
+c7+EQkwcJ1Y9ZGSmF4/fHm0Mb/kr3jcxIVgD8oYBEl6XBRDWmftjRBHtSop
7nRzCPgRGO9uSdg9R/vpvVi8Gh/RWlxpGJJ07xi5gbLxSHVEy9HbEwx9YNAq
EAoovJjvZQYt1ItlUudVQp8ZK3oY1qjxtnaJPo0pVWajKUx92sJBNn1MgNad
NL/haaT3Xf4/CyjeRZnhaMEUgCEyxl1UWLgG8W1ScUwT81jZGRVxNFmwZ6mH
z5M9uq56uUQKDDfllP6h4rPPLcpX9pQmoUgv99dcUwSqzvVqxnHt7R56+WvL
/TLjlPFe6fG8W6O8VBzhdYqvwsLqycH+FW9TdFjcKhktFlFmuZRgn2+x9Yeu
pKbAKSHmCYNjsNajm3HlT6LDFSwN0V82Qk8Ioxv9RezyO8KN4GYedJ/TJ6JC
JQmhEWQIHcl30RUhAwJHbK0R4GUzetPEz8ky0HfB/dTt+avAkj1lUvbCgsQp
3dXEr486yDR7Yfv+FKaM0NhvhdVmbMYdxETajrcFQHwdWVt783ZBwZhLH3vY
TPO0tesS+PK+mFy6F4u2W6nemoDRriDdx7CT+4w0FgY0/mlHw7GDCRyoiLf2
J3dZfYyfuLKESaX9Z2JnzWRY/Wyocz1xB7NHNKf3vvayILJEaSjXouJ9UKgp
GcfwMHF4ZNwKF1CQdoc68Xm/hA/7kyJ51rc+9N01qa75yu7kG/U9MAfv/ddg
1jVhR07JhIAq6rIPK2h1GMh1lHrvnIzBxc2U/R7Ns2Del+ieyoWvKXHm6J4Z
QA7k9r5EpTs3uQRkz8Ak0RgiuCYO6F3OESWGOg7gdHCpUhOiCZtifEKGOKlx
NFwUZnPo/Y/kxPJJk9+SYwXS8PtsVmTuNht0wi8HjmXsf5kQCNMo5I6wm0Ty
S6/0bu2ygt7u+isldYmerTuGM+bbHDr2poAaaZcx5qBLICyrB5zXmIfPKt+o
HPmOxOkP6O0oDWBVAo30O5Lr/Lz6rbhVJmV6uApdG73kkSZ/g0E6IJ6nOTlX
xjSFnIAfQrlJ9PIwnNPUKsu5dKwu7PaTtb81rxIOR2PaqV3wJeKL7t+RX/Xs
KvkG688hr6hNDJcH14y5GXB9G0LS8rCVXFO32t4KrN6cSN0L9zsTvIfGm6M6
/7WAGBxGmsBhtk4uRBgeUlrPx4tNa1LnD+OeousbcFtT8T2V8/mhc+OsYsik
vvO2MrgTr+31emK9/aiIIL7/HAXGZ3z8CGOwr1V8Tuc8B9S5SCUaMtCGQ51C
RahEkTRaNxNxWB0gOiONzZIVnczLR1TfEFwJQ0lmSAp7RyI1McAF+o5mQ68U
0j18EYVbtzAJmHiVvNaXgiJ1LL755yKg9oG4Dpt2HzZe2vxZ87HG2wDoPi7M
rvx+t0Zv83BimNzXrgwj3z9EzCnLmblHxo8VnUp9TyvdPRM7JCCoRdTGz442
ywSbO9E2l8tG0coP75knhjIdB505LWi5M5QOOOBJWlMg3Hi2DX7pAAucCLRe
Z8p553/RPkcZwF/RXyYHFu7KS6QkvYnR7hp7S2tF3VBHewTOA7KzG5+YpJNL
tDF1IYrbu6KF/H567C7VAFhVmvUGqW4firpioFPXtWTjhfW/fyLok6wspZy5
Ev14GHqnH3pASKIAaj1mkSwURYc9fupIF/iVyXwvM9T2lhnvbzSZTnP6IJ2s
hMNqRDiF3Ak2WlWnDkEZu03NkBX3wdKsAh3okyNyC3OFDj7cLFsIFnXWSj9M
uuiDfg4qDiqaOVMGbNKRGKVMi4O1aNmxEpiXoZQJzvvde9xFRcz0Ple74tK/
wxGeLHDyNj8ufk3M6xbnwkaYEZo83Zihx0IfXGzwz8hlydq4QoY8lUF8KxTj
A+c9SXaP/SD8v4NKLV7Kve9aXU9AiYaN3eh+BlDaad6XGdr+dwsyo9QrQJD3
rkGfhQpokv0mbzktQZFOKHFTzPAtpjcL0SqkKWMTd3t+EvYuYs26HT1PCE47
dYH293y5YAlwqPaAA6+TnkbUfXk8L7PKhXBLfMqeaIENTMdZO7CZJYupqot+
hYMzT3F+omcyWfb02NfKad92mqd7rgNXpPkY6GIc9upIGiweLoDDCak7+bAi
i0izftKXb68g+zvO+z9lMHplv8cITbXy+jM9UT1cFCdQsIWsrfPRZCMiQKTS
WlNwiBUD36HzXcwLbwHeR15ZkjCjpUyBQvyeP4sdBX/PHnVr+rwuYMbkltu3
h810vyh8Zv6UCjrljHp2tvZNxLCBUUrv6BE/A4liFsO5UOMmuqxeAc5AShno
M7woyije0rCYDDWyEzJ1kcnu8k3r4hdb9gvcHl5y1z/xsPXCdpJZ1JpvBSgY
f60TB73qzlNQfBzhcCQAhgnLW+ayn2CRaHD5XimehK2O0lxNK+dH9qog4o7q
/+2m/nDUjZipfGjNkSZMAb1yERXvw7wqrXEHW0NMuc2TylhwULS8wudUPtG6
nY/Eq/LyLuEEQAm2RCXEFdnOMnTSrShhf8vu6jtqoLoVIxi0xrMXKxatzMyA
1UIpylNC82aSK+IDbHExRVKGQoL7s17KbgeZSuVB5adWsXD81g+nRWARbpj2
M4DLBbMpNhrTOqU7lXksQcXOdb1Sh6RoQeUVplRwGRsYKwqRxLfVZXIbmc/2
pZT3VHzpIAW3aRSzzgoa86ToJh4tZrfqjk8sJTVkTpopO+CLYn6W08uSCIhx
lMFc9PrYuHmt3KG9Y5E3ZsTM4iOe745ofeoMhzR9GQk2TJQOtIyEkvHbWT4p
PHPE+Dcun9L8UMPj7TWc7Z77kuQYG2ZMJecaMSBWWFXXsU3GRDFl6APJRm5V
evZaOSshS/LIdL26judo436d3bgqAy4YGpDcSlB1SN1e9ykMyz0ESgKAMBPe
ogBV4O8i8xsPcEKEZqMlxGoIsB2vv1ufoDIMpZBaAl0oYHm3LNc0jpYRf7Xy
wIWNDcyu7NJGodvhlhy1hjkiTXdaosEx8IfAMHwUvXM06/2UQcwV50ru5/R+
LirmZeuhcdi8VZOPs4hyGA72PKJ4GG2k9M3F81S7/P+1qhbtNukVeEhopEgk
xn/zPQ5/I1rHXMQhTQRVu+MS0mlsvsGQRxGI7+8+t1DE2ySC3TN6kD7MAIoU
PjdkroN143B0opq/54ep47ALCOmTASH+ajPXvb4PmlVjm1neSD3DZ0bpaKZq
OECmYgDaJSPLO4F5C/r0m6x6IzfE65sx8boE1QRNu3e/2GIB6YqJngjE5119
MMbLUXjFZ8cLpKG1FnyXKAVVsmB/AO4612lo6cLygU5Uw+eQrGhjSwimvcrX
ezeuhaYXFubvOC1NdABgcy5IAhGDcE7vHwpYzrtXRpzF0/bY4izvzI+8KOwy
LqNOPT/JsHsEkMYnB+ev1ovxW+hgAe4rBR7KqFRiZHYXCwpprZzXMC1nGb/p
R4PQbgnttnEbNBqfTE70keIdxPg/KMBGReMXL6BE7kiDxmraP2+EVS/jDljP
z5cReoNyy9KohgBo4jiZrmmSMKTZBdUi6GNWqZcDI2WaCnUERUVxBpdJJ4yY
garJWw+5QUSwphG+fRMYPLhHuNwv8Mqux5WXHCxnCknlCJZNNHR9y4S5jgoo
QOIruwVakSv3b8gdAHAb8IP9Dt3Jtda6G2gwAHgaw1jIQIVG1VQf3k8se2T2
I1R2xB2XVSt9mkj7N4CmUbLjwNrAvGMZwOLLoWi0ufKn9Opt4BbBGgjBeVTg
Ay7Lot8kTGjftp4HX3RdA9WLBO1Xev9dL3ICErYO0YPD1LWvi87GTW/PJD0I
r+FORbnrus3J2lNB3vA4t/1/E1224Kjj+xQcFsQcrcju6CiZ1w5BxNNX51lr
HuGfZS+sWfzKDfkWc6HDzliaQNHm4gZ7mbEUSIHlHZJZh5gusORpja6IcKpQ
CXAicbvgYCYU+xm9N5pgNl1oJnkn1OPDb1R9ufKih4KHTo/R+Ly+osy8d0C6
U18F6iFjfgo4M8vsrvI+tUgg9WJXd9uDWuWZwkiMjDT1j3E1ShPVvr2a2X2F
JrMBTelmktd9F/969XP7aZzEvsPnwTGBVfRo/+2Xidrqe6rGXp3ZJE9/Nx64
pGjsceDTspi6cF6agqN0EZmDliqwcLvIPG4UZIbyIkw6FNC3813KXnV3j2sb
PcwjSUDMPDxZjk5Lxdw1wzbLUpDxxcbFVY/odH/VRKAhn9xBSRRcM3Nmu0nE
IYnZF2ts08GfJTuffGqsMzAFsSKn7ajutBlkVnPv+FW4QrtXCwzVUb0I9rBP
J+bVIwXn+RWVQZZY+EDV8Pn/MlgmKTGWF/CY+KzTwXAiKrZGKmIw/7yFUKKh
xoLkzhT6eK/kaDth3IbMdQs7K8Dneu9WPFNiRGbdzq8IWM8gJAFnAaouzN/g
GCu8jc7lgAEcWS4CHT+qMl02JL2JLWbk+95wqXWQSZ3bg5zYuRSqthyap0rA
iI2yDbVGILAozODC/Awunf0iAQMA247Kbphet/jEekrSK1cptTOZKGnM5Xws
P+Dd/oHsZ8kjDhsRBzmV7LEPq5fZCx7VJnO/BFn+pzjoga77jR+80RmMpHP1
8jyVwwo3ocP+oConLnD79bal6F+OXvueKltIHvy7qEdEyEcA0n/u/xKEVc+/
7sL8aNazI2HnbIKPz6t3fE7WRm+F07nR7nC5s6wT89BWJn+3vQPd5pdhAhph
Jd3UBGuvhEfMQ4V9vwfJUqfStyUPovCIBJZT6MD5xTbbqsOVTGWESdIv1s5T
aIauCk9gkOsDz58UuxMpzdvk2d99tOStRjKksqGFz9lxsx/U/nKhu41aPlbF
AfirYlqDDOXVqY9DqWftcVPcLRSmQBCkVVhfV9syQqTnS8VJfc6OSD/SCX9C
NXOK/1Goy5qi1XG0jCGN+I5M/4PqwJc8jQ44Ut6kRcXgwxN5loNFi3mXuA9M
t8Mu1gG4B3/fq06BGJiS06WAmPNoeTDp/zGcZK+6vx5ThUBRYhaiT5yegCiq
FKuVrlWs1+IjMCAjb9SZsxwB1SGT1vwoHpOvSDPSEEFYEGX/rMcjYYXJ/J2V
uy2/tvx2QNxS91ldh9/xzRW6WTuk5pVoX75dSt6OJ4pHBzOA3ahqUFVyeHni
aTXAznzMhQDjB7IdFiBoeF5m6pTL+hp8OHT0Ax/RwE4gXSjKTNarmotIpTwc
nVxoEYeq9ZxC9JbxQPnNalBG0CCoPp0c4zKUUDBaAd/VIhRYuH3haG0LBg26
TpRLSGQYuyxxdgHgXipLC12MVxzqTovNOysGpEFa/G7uq6ulDkejBBNlTQia
uwzmTN8NTj2LE6KRbzUPHPZdzoOaqb71NhBEuGwWLY+2QOin4Iegum+zLi3N
Fwz9tiWvaDa0SmVcQq7aIUJw1hvH3TmD/5WoSQCDptL8KN1FJFP0gEvRgVYp
h5dc7neLWa87EWpL9gqwzAHSHtgUjDSobU2ddGaQPUHPdA+wylxLWDNIrKy0
SgpgsuZKwu3JK2C/9k9EXE8kjBqEanJVU++bkXwZqSGHN6wn7ufU71C9w5Dr
V25gpymtrKMpJl2icyw2grX6TzQ+eosWYALC6YE9gyFo3WzTXlFek90DDEQD
0XcRixA/rCVSQIAKGZAp2oETf3ipOOxBWhNWChwlhSBvw+uYV6m387qdxYbm
Gtohw5Im7lJayEn9iTymbiDMlrnk4EYkdeErr9DH6csgwkYPC5QBuqzkrJup
6i7M4u8u1LZbEW7E0nDDNq/8EJYcyi93FO0YbKuuUl+pT6sVh6pe2eq2iiuw
sailHdtMTI1c7XyBYQbVCFv7EeEjiiBpAeSu2wbPerHb0h4KE3L3b8HQGFe8
lEhW0rcx5xp3oPUIbV01b+Rf3E1ChITDQl8mB2vysncVH0tZBnOhkmYHDVfz
NWASre1VcyHGsdfYFoMroic7vnq9sa8yecQ+KgX+jdVPccapIJTg6OBJF7XZ
R0rdX7bTAYu9nl+Xs+cRm3VlZTJnhd0NqANJYFn1q436HyngHk6EY1anS7tS
mui1wftGyxZtXJE44xYgqUdHQtx4qJtehysPc4OvcIQDlz6MeiBt9qx08ob3
F+R3q2zso60A+RvmkAUPjhM4Id6ztBQoC//iaZUrT5gBryxJkiUwhzfybaQG
gqHCrceWKovXDxPkGm39GIfaam2HHQ2ziXw+d+3YWuD2b1BEVaw3MmKFQBrf
LdGDRZIjmEp4CA1q39Zb2niscSXkl/TLyiK+004tj5dQcE4vLx5tpU8oY0xz
Wix4Z07IgHBhHOn/n+c51s4+quhkELskVdw74wwDZmfR7azyNJxig8ow9D8V
in452iaactB5i6enGRZu7ZpePa1VJGi3elxb6JBBC+b9XuMbZo7wqYePxziQ
TOh6I96z/5pb9Et+EQnuHLujPb8j/XPcYDdnmDTPK4tL19JuTyN91wgO3z3r
zxvJSflocENJeoZ0ZvU1ccrIKp3I8YjttyMm47KG6Eb2hmuKo+fEHU1DcVAS
SraqirNeI3vXDc3wsG3BbZyIU1vJk2nb8loBHIeIt+cCCbIV5YLU4Oibz3Dp
BT1JCoTGVFsgcjF8h0+ZpO2i6mwF3LWr+o1uYkf+AOWg0fQsyhSCcoKkNbdL
WPrF1PudjH+okcM2ivIvHg2Mwm/wcNr2WNmPnUhJuGxwbN8ylZf5C4nHsMyn
lgYNA68ChTrAkf/c7ya1774BY8uf2ghbW/iKYgginbk4bj4OI7vAil3PCsy+
8rfU++ZPAyN8J4RSbbvxZc7rmIvVFJYcX4Gw7EXwVt0cv5G7jechAA3xgahL
XpkAmGThH/1NazXhOFZ8oh8VFB/FyQjowaNC2n2nkgOhlmh0QWRhAoH70Dmz
Kn4+ziS/jbE7YZqVNicLCAK1/x2zC3RKhw0D5wQIyYQE1wT3/GyoIFPyuhn9
hmmiXi3ZmfXkfKn1kbXWSVKDKGaESc14tSqTLccfzVbBm+WlFWzE2G0hi38C
2u4Dcl1NI9TZRjYVH8+52ozaeZhJH4hQ4e8t+Ke5eQyaU94i8Q3FF35qI773
69FoXvSRaPw76KHGp2yKrxLJyiaL/wJMT58V4b/8NJUSbwW88Czw3Soq6zoH
vaSLuiAxOLCggXs+srej7wMlXbxRYmX1F29QbzmmGbD9e/cGXSW5oSbw1teH
vlXC/sykvWuTW5T97KxVl6mxdwTd62RpB01RhXSi7syvq6rRbIEAxdj/EEwe
19D6bFLRv2R1tETC5z/0TMMDl8RRt3MuDBRKLvlSHwZFs3aRzJU9h1N6VX39
7kNMDm2km5un2rWyXGTabzjDUbaF0k54+GhfBD4INEfrYmvZyGkQPa1fg1fc
RhH3N6s1VMBzgNqvxTcZ7+3UY3iypVlx5JjFeeRpYYmCybToMfIoCVUtozZk
A3TjO/p2NKep1zN3iesnOksznlOaGQak+zmMrFmfiNHFGfjYwaEuYJJGPDBD
8sdyfrDbn2eDp37r6nsJWxQGeEf7Y4C3zQYGq94YWx48UrUjP0DWlsMmaV4/
5MEA+vYMdP8vF5m/dUveNq+/vPd2qgpnGRYAJpnWHb4mdo7UHs5yTiMdBXQD
rPI1fT417AmosekhGFh0og6EgbfGs7LQsxrxA01j5qZapiB6fAAEuOZEy76H
6PY3jkMEHXU8f1egppT4Vj6BnIP1pnrnIolvn0bzo/PLd54buXnU4zRf51yB
xi8VZ6xMDzZoR6+v7m0PmH9XV47KLQZTaGanmwEzmwOHBaPWIVfmkD4arULT
jV6rfV6EyXgQKeAJm5OBVrcER9TelqaZ+eWUfCqluAXE6TgU0ZhnKS73OFCk
ZpdRoKTQcj6d90EJMCkt6Re5Alp5/gVY//fqOlavuhiYNDMA6Jp/naEzc4dO
7rWc9TXFUEXuMuCWbMnNU2fTYqBj4otGGLF7/p74F2T6Mhs9jRwWO1JmygRO
VAzoqs+8Xe54yE7XAEltW/0aB/rMITtSkkvuBX3JbY9VCS72k/mdEXoLP++E
nGBqteHq6sDsEttCKWrUgV5JVsx0IhMkeaX1e9J/AGmE1Y52S9uZJdN/Yvth
BRkK5zMJTZBb9JxxhMe/QceVVekyHPujvvhFFY2No9vuu5OiO2h2dPTUZ9uq
ok/o+5gGoNNabK+hr/A2XKNGVcTrHt9Ct0UDX/FYySNwbtE7wCeioqB5pUoh
2pYlSfWY5LxIx690eXvMXDGFu0q7hK7Jc66YZsO8oFW20qbkhaL2TiI9DAkG
Ng2CGCK4R9vn94CSbN5VEAEVIXiKLEsSVKjBHVw7sFT02GGfP6iUJ9HyK8Sm
O+Uz0LifRrQj+rR48a0b9G6JsrcOWBYlMbd0HNimNoR9n82SKPha9MSwNgFj
fxxb72bti0u+iwVl0tCCjVWx48kH4r9rBLtbOrXme7gKrQW79R6WJMlFUsM1
xEYG3I/csmhuyB0mAsyMz+5O2cE9E6Yn/tWfuUAJPVJPww+cVf2QXRuxrpIe
sZgbdSmLNm7t3Ysh5lHll/MveBcX5HTWrrCf104CErS0/Z6jlYBFVX+Ok/Hx
RZbWVUvazB0QrGb/VsDLn/RyCa/ms/i3lJsXIrYvZ86fI+98Grnea+nHSyTD
T3jBLNzyUoacVlACqQ++HzvC+tUh9zj/gxUdqcQfqXXhr8zaCek6FpNc1nr+
UkXdjYmu/OLVOqEWYArZTBj8ypZC59ely+SVUniGQ8aI8nkE9PWOpjCt6B0X
ql6wIChxk36lKPMJR2ZWKPASx5OaH5EUNYkFWXeyTb51tpKL5AaHB5vzjMLV
aG29fNBPNDSp5DE9vjTVZJGnJhzW8T0oUYmy19wNe/1aFnEv/Uuhz9Uz6oLP
9MRMdbefOlUKBQBLG7xC3brkAWlV0u9FMJZFCFq3e+mpQvWjtPAtXtytFEJA
hcIfiV4MQXTRBuQ8WEg7Zr2Bht+aTquFUNQqlbbVLLfhNZWFGS4RPwoUAKhQ
3ZqGLtPqFLOC2tVpCCjXzDMJyQOFq8nBuUDbxtQn14OVKOsPVujFqDkHfLHc
BausnR/odd1NtRw2NgIQAiRanRuxWiW/lOPe92k7Q4RIv5xDDCAPGmCM/xig
kM0Sm7FBA1onEBikbE/Wp5u61WBaZj+1Lk43H2/Si4qrsWdcVEDE7KPWAw2k
6EfT862RMsDpG9VpMZ65/Y7g/VihFbcNMN1oGXkTY4+rsjENQ/0ap+vxNRCI
4+3ecoMuBL+IRNEjxicHzCVp7r86ZAjPvQZs1E5qBvgeukliF5ey/RES97Nm
PnPPtAoupBJjF/W8TX9LJvIjRIup6BYKToFQhxvC7OGIyPZz3VttUXtoun+P
MYEvf5vPArrY0hXCWq85Hp7iUl338ZgSc+9rxn85G7LElwr2SmzTFFKrcS0B
weAhEbhUkShBkjL1luhh17eT2Rgbk8YxfRLjy9zsEyxIEHtKzCkH1xErxqIi
pMfUWfVjGQb6Qx6ta6VEArpnPGr2s3Ti3j5WMdnNJXbix6hhK/fDCZCOhAUc
yRstH1x3athil9pwuUvEn4LDNSRqm6kLGo+VdumD309Kw5kMoSYmqjny0xf3
LEWk7r+V9c94i8x+W91TREPkA5KI24X6aGdFipKnBLPf1BKr/mpYOUivbq88
p2lUIddQIFd55iMUWwV0ri0Xfm9T21tIWowmf3ztqgVNaIrWXJUs14zF8GsH
vXeZGAGJ3WkV0/gLapMN6m1kP6PQVWuXNR7aXVYTWxH6wfJ6nBfgSVs+rsu3
T4zX/aB2PQwIT1ibIh9sRVEthywPC8pXXtLwZS3JmRwOMOX0LXvM9CYW7nLh
E+oUMlR17klGez97iiR7o0SSQCztvLJispd86UloX53Dv9/RD/m7xtJRa5Bs
tUw60ZJyLXukG2qqjZtvbey8yxsPSUDR64RtZQi1H6n6Njqrxf0NZyqPwHrx
UOo7D/4qFX8kQw0EZ2J3rRBWsXWaj3TgrYoK3FW17sQ2OW8R+s+K5NVQ8n4x
ZEoTdb3wFmw++pSeL+7kLBO5z8qzDMNaG0Zg1Ztu7SpG11utEdm3NyeJ3RL4
lvN5IWWRIuYaX06KfyB5W0J0Q6AY7g4kaXM2Z66+o7CJ8XFTtG5EhLHWaS8f
KOxonQ7TZzpIjVr/8uDrZnA2aV3MSer9+4xAl2we2skxAdGh4vGShUjvJ4mt
gv9PRHXsM8t+JUgiaa4di9Fs5ggqlGnjz6y9HKYSZPrVRrXSeLpWDDVrAQil
I4hgLtJdalQFl/kAywMwGPlIdlJrRLruphDppmiY8Ksv2yD7NlBPQPNEVy3u
xxL9REAdjdeXoYfHJEcFdhxj2C7h+lAcwq1LxXuZO9hO31oxNwMI+hlMZ7sN
3BdPnB2iIVFEp2noWg29hEXCAdB78TL2VpId4eiizUGaB0Or/bSz/BOn/GYP
f/ul8RiElA/SpKBv9y8slsbQoiHpq4FzMV5bbgMCJ+azkay/smiTgzqDWaQf
qZbyIrfah6HbKzyultS2q0UytB9QeBcm7GA53Gn7QEhth+HF1eOfEXaXPAC9
+8vZmVLd1j0LUBWqx0vzfHbv9YJu5b/sVjcl9wUD+sLSp6+JutEs8uTw0XRz
d15d7/SPxf6gZL01cNs789HWLxwoHRUKyzo9LbWuzZIxaDhiXLY+6mWQSYqf
GdONBvSvpYLgX+BCWlMaB25OLnG3k/Czyt6x+nYLbXl4xnHzGKceLBKueAip
eY8ni6o7wqvg4tGmqbh1MK8J6ihXH5mWx9rwNnywD8Mjg67SlEsk6s2CXRQx
cEPx7ql7R+HKn3axtahPCKxfBFHnPnDpmBpnR5IE7JwpYNTT5xS0rcHJkOCr
NJAOjfiXZYM7hW2JsEOIkk24nZ1SEXyamNIhfTtyt/pYlfEh0RIMCVlI/AH7
oSlLHfpN5roSX3Y8TyzDwbMpauMHYN8x/9xEVcXSH24wndPibbVBWqEfv9Rr
Tui2VBOFDQmqtm72pAVfDnIqcnRBPf8vGv16DFIxd/hKLMimvVSRMtPYizNY
urNc5Yxbh+7Wc9rnusCyDG09tAXv4BwleSaMGS7QR+svCN4VTyV370plRq6x
akSo2+e8TnpUZ3yYhkgdUPI59rufnkQemVn9jMoyUD3YpAnDvIEh+9t/c4fd
rwwhO4c3fAwfCWUX87MhwluMbLqRHPXbmsMXxYndVRb/sLJdyg/fye4eT6sj
uXhZ+D28IKDURGDyCFJfQ/HaO1u7pUR4GNdlgvY+9MolICNclONBS4/gfNxm
IKCsPfVdsTfHtKEtUv7AahyEton+KpJrJYDewz+om5fb5Q+V2XALVcARaQuQ
Lz2jAf970CA3AKX/a5FzZWO87liIf5jmW66aX0Qjf47/moEi90f2PLvQzFZl
LnIx6QR8FfAEC5w6Hl82LMiDDzH7VYlxTMyZHzUFN8O1y5HpM7aPiuMTmyqY
7mljuelevPiIVP9k74bAvEjwAKL0ruRzIszH4kewFISE+csXbf6z7RyxJEiG
etYyeDQT2l5ux5/tHg0spb39bLtJ5akG3irx0V0yUkLSTmV96caR2Vs8apes
0nC5LtoqlPqjspJCYq8WhdjLqrncM92UT2dXTEkENz1utBJOkYL70AdFOgFO
iW4bVKYZM00h7gqx9IoWSI2/F19mkkxbuJAJVkC3aNrVTFf8M0RJQIOKBX0D
QkMptndtlanNlER9j8t87YVukGSiI7mN5emYjkLkR3ZZg5ui1DOAPmh+BWkI
qaUjCSA1lrQS2YJe4TZQQiHmX21XysM4fgDvgRfDRbCwYAHUa83GKzaUzr5p
CtuLJLYt7/W8KySCCgiN8QlQ5NSapIO9jRbII4lj3vqAsTMKsev5DSDqzpM0
ppFUcYmIfyvSfyHJYdL0/Jg+U7w0o09g++2VvMemUUV9KLbZ5RgWGpDMpGaK
d5SdpYeM5tnbRdWCm5KKOiNUMpyd1TYtwyR+lVQKdzxodE5hSDX29dNexKz0
7zY8ho8Xq9fgFT2zJvoFaU0NC/fGyOAjh15IJKioIBoYFMa3apjnqhEe/0jT
xDVVRY/uJQ26ekhVX8QIqsXIkEw7gctFbNIvUXJQZEcWZsY3nVCy6ZmWT9pR
2c6I+FWh1xw/geCwBcF8Whq3+3rwCNZ2f9sjVCEO+K2NTv9A7wLJJlRZCukl
dMjqVaxS+XUiVKSBe1BOl3sTMicyXbbUkMmgPL7bL4WRLWzO8yOTru5DVcRl
si7mV5/OBleTqsn4hJoxwd6fAdVt8QyGzw8IkaK6Wyx1x6zfO2x9QT54oQHW
70qjqO+OzZk8OpZ++f6DmmwrLu5oNFt2qRokpzLeLyUOOMeQXs9PMoWGadCj
UoMTFdUkoe7JQRLTAGmlNfAFkrxeV5XU+rOOStzh1eoYuHWtKJTsl8wCFhEG
3tkXppxpd1HWqCyXgpzakEZMt/Ilao3sN0Vu7TPtrQYf+DT0gmISTFILXqDS
qtx/cm5Xm/OW8C8eHeMjgX7yx7qX7/MGulrG9f2d7kc4EParhRIXXxspQ/87
vMFBa1vT/jrB/3TZ6Hd2GsluAxhQBd5EeFR5L11J6eNDwkRdtJer7g0Yz4mp
bPS3G7qoxn4OY9vdhgh0QGuXrBzlz1Oqe5g7hGsgGC5FV1rgyvx4ku6dI68f
JLj/v/RhDwcn1Ug/eE5Av7VZQQd3NMwgCrMILR61OfrdJUb8HPf7+ZsaT5ff
FJK+FwTjdN1StL1CLz35Zzs+QuqXdbP8qdIh4ESGe52cHjqxVYaJ6zo1eXMV
1mwijrAPBrQ8sZzsDEmu+xmMtkZK9QFhL6yo4508daoknE+wN6hsiBbw5z7h
l8PsZLsiY4WlCJUnq8WRVGO4vXRSHkSr4EE01p+AYqzWqhoIrugLiz8yarZ7
LVVyqE//fo0COWclV9oDi29uHAmm2so3lCTJVDlFGtzDWGf4T7BtVEppp8Se
td/yV6e1URSqhzj79rlDTAoZuA83bJz00pADmLWFt8JV0FBKAZcSW84iq4Sb
e/y8HDDspIvDitk4KM6GSeXZNZBHiEas6t0i5EBBfnMuDymrkaUBYdiQ4X4C
RWVCk6SBVa73CQjsPWpnLxo36uyS7iJ419sqwxUBwLRFWwNIATEuJPJhH1Ol
vNV3XCdoHKpkhElotkn1UotBMbeoTafQopfubl72mMofS+UuAITdpRVIG/n/
reONvjwwJKz6J8uGq8OtozDRKQ2loxikfdflmsbygEAYPOQRuzHxmuaM8Y/w
10sn9RWSDC9QMu2fc4JRXD9i8w6LflYp+3bII9JbmbZgDkbSmYI8ehd+U4fa
8FrCCkXqY6ajNaODzr2Tz2eRcDM8fP4M0DEi72vC5dFfJ28B8f74GQ3i4Vkv
m7t/OVH/yaxQBIclXRZkN/ZcB8CacbwC8jm+JplHsU9r6JEbBc487pRFgcU4
/4+n4QZyZ+Lqku1hzTNvMW+eqREAQTiGZtcw0DmXfrXbsUY85Uvh/icNptjp
r1pqwkSCkPj+DxnooSLfji1UMsr1G9bSd7MSfpmmLl+zpF1oL57IEQRJXqcE
3X4nE02W813nuhZbUPQZX8CgfuJAX1/vpSIYLlpc7o9+f2pilVLxoa3OENP6
8p6HJmpQr2Tx/OhSAIz+JwyvICLUtcIBsjT/+j8kLym5dZ+fDMl1v2jfjypE
m8Avv9BVrUS5G8x3Ns9uuYnv8ySPYW8gX65GddyAKgQ0Rbm73+OdaGISny5Y
a1KV+PFrtvIYe0oZs2XD5+0K7splY6HcA54/0YCQ5ou8SERR3/QCgryVEn0f
E/qlNdnCGhDgo5ndG8K3DQcwD3G3G+8qjeTfrZygG4g6PN4K04vKqHCEUZmW
AtmP/Ea3bC3CiHCqz4yTW7obLPrUQ1vEcAvUbBvmykG+J1rHZ++B0cLp8xf0
YowS9trEgvXFW1Wh7FxgPXoda6EN7aVC6obnOV9QzJICDkGwgBPL6MlTb3Ft
oKsoICAyENq+WcvZW7s6IgNJovefdu7cifyuIOKZs6f79ODTAeSHspD1kGpP
vaH90/eAEV/JOayRsbgW0SHBS04Y3E53qm7K3o/TVEfOK8nIQ2RtDJwlPzDm
I2+PDWxgW+qUS+LkyHi6iicFnk0ARw9YKpH2+H8qn36dZsqmmkwehgUXl82P
szyaJp0xGYMbTAGca9BitLAa9A+eFhpwDHBsmdP9A444cxn0DVC1PO0V9QSj
WrS8E+yizbOeyNLPF0j87Gdml7/vpV+Uz2XNZdjK1DwSFE/VJ6KzqnJS6OAi
vWU9Utwni0j1lEQdoNjguhBxAYo3Rgiv8R4ndpqKCEuDdofsSg8oOrM9qcMf
qHZyKZUB2L6gm2eDlwjYd9RGtLYPHFlav5fIH/6KPtj04X5dmtsR1xhkpZ87
ykOc4w1sXuljmXGJgcyK3h3DrgfzBSwho0dpq/Fjz+HuNAWyYqNdTx2guF/1
fLCWj4c0xcwFqyh+POh6OKM54ZbOzUHA7g08N6R9iMtfmYYLk/KQZiyGaRLL
jlPAmK7UVbmDE4gzyn5SbwQ314c6mPLc4HQEvJ+OP0g5PQEAw+0IqIIjEoHH
lblhyM+xCN+tu+29wd0Da9w7WQjVyDownjDx+WUOWSV5r8iqPJP411HlbaO3
Ul7phyRoj0mx5xXujDZ9ZYcPOQLoIn6B63A0p7IjCiUFvRx+rC2k1surWpn3
KanuUvaAJEUGasihQH7cTI2JoYkyGYNQMb9qrNbxc+0aOfOxvtKA9eTNPjov
BfoV+BLwuUcMnOnTqt31QW2XlQq3w/1tAtzCXkKfaFSssUC+rtFE8vOPstiC
aGG8I/pxs2XUKuIMDgmRozmp+C4OATlQEfXlhiJRavkQ3QkSCiZsmhughu6r
VX2R40LiQKaOOi7fEUR/2BN4R7Av4z3TZRjcmbQeWpMyb17K/I9MGb0PXfEc
37xhAQ9ds7A+F+5o1iNxO2C64EkrsIOAESuNZvRM5wiMOiJ5GgV6jpSu7dag
bEVTCbr+bI9C7PJXT9UqUpdJVKJALuT24O4NGhjieNc70B1vrvX5v/1f969w
X72Wx7wBxJccazyJbvZTRhH0UArEe2vHElcUlQCubgBmFwDJ+eFMSohUi6Wq
95iiT57YPgrRqabbYwsoPnVrTPwzDbLpYff8fclaqaERA7xVVuP5qxfMiMXD
9xV0l1kh/IYZ8K5s0hZ3CfJ25P+2FgLczoiW9+J5sDAPgMnDcFDp6RbASTbp
vXlpLvM4qaMWaswRiyh5Hgy7L1Ra/mFqULqptTlncrcwXJDSvhDaa1B3d06i
VE4OVgITYvXFrZlAsRB03VbJ+ViPmCDey/GsX/bTDZKd25LXAmIBmD4+XqKX
H4C4EvqrypN6G+HnXiB0wdVbN/MMfvdjz/x6jXHCcpbjbijD05bPDnO6lb/8
qQkzF0Ksro0EtoqxAk/nT3oj9sR9Xb/wc1TICc6Plnb137fGAe+RlwSrgyUZ
2DZI5jsN3LJBjSEUTUouXk40l+l3QCOw8aajnFtl0uhDASoM3E3/UrnzvHch
Tb90KnY+LZeU79fSGsQuwAUACb3QU4/oKxtca4RDlEM/ALJn0NXn/PjtQaOi
IiO5vOMWeOVEyQo6ScZSILLY+F7tW5SyTQp9LtFPykYAfZ3B6w8XVHq3maKS
icyIA8LyGY+snOTs0IVtozA5RwLPUSUxsxNiyEl9I5f46gjONFLN0SZ9oq3L
fCjbU0PLpM+eyOy05tcg0j4sxPZJ5sSCsnL/4cvDko7ca0bO99eBwQeTtQqO
OTjJywQOzEsGPU9g1A9xtdjo+W1f+BrsS3zHV/XK1hK92GHv9N4clj6jT3lX
5/ljUBjcmShb1OJ1cjDozPFJKw+dQdX6A76dL/iQzxxEbWcUCgH2m28d1zuS
IxLT1kVo0qBZDmxWCPhjRdkPbJaBpRrpgUyO/QKO1DdASa/4BxVn5SSJnyrK
EFUPAyuY+d6gYgYoRQ0IT0s7+Vjifbo5eU3CGHGVULAReFuh0sqmkB+vipCE
qcPvaVmfOjONlJ5oYqXkoNzCc+i2fVHQEoB2i5LwkWa8Lw+bVcWZ6P+iAVhx
6HPb+FLDqx9GaLXW+W6ZJH9GYSyY7OHBZ34Tt2MgjAvEWz5WAOI9/sJrgAoT
UXNfti48vcOaPGdshznm60PyGndQeEnhKtAuHlUO7AI1o/csdzt9WGKcaRyJ
tUjIfionYGccxIPhULlU0V86EWSBkKmW/L+2Bj2p0YEUiVuhL5aDhX3YBCQj
S1/LsUtqM3LYHHfwLIHcct7IUUe2GDiMvBDYpE4Ev3GRDjhy6apAxHXUYgce
6UoypJNUuaW+ucGiuBy5qu5edSnzO9LO/2bJDbqG5EUFfrJh3ekXJzzBqEN3
MSE8rtjhQyOEZGQTw4P/YeHjTtFb3gedwupU/+GlCPHXqQmdHIjYTdloSMxZ
mMbOPf9sUbqFNZxToRlP7MjkNA0nyXFmXpkB+COkeYlu9BQ/nejbYeiw51+/
lH2lRSTgwwE7UmjJrCutVGS89dYee9ex6VpiWakVmpV9tP5SYWfbFUhgS8+6
nwwHnxhgqKgCEtU+xIavI9Ve95QlgVbjIVuFsweIBB/OGEJ8n3BblYvBtYsa
129VbY8uUewCMuUa4LL5uInwwXJTLDo5R7THT1/cyGrrGtO1TSji7AtBqV/z
C0+NfnOVrPygOCn050gu+P6SQyIlPCnXo2HuR3OxONnFPFBENNfCRhlLvf+S
5fFANYUJ0BzEGs7bKuirKozG2mUWQeolwJOJD9jyu+Y4v7hK4IZ0EhOIolXh
eYUg8U2WCQK/NmTWlHAwqy504LT+BDaGGzM1pkCDJ2Fl24b0iV9eciRxedk1
Iu09un9F46Qa9txPozA5bCAsyFzZrYrZ0tax5NY914vL29Z76cLkTdykFdbt
JwYPPmXPTPy9EMqqSj/bNlBuRH7z3lG1OzulbjpiT5lrPUCU9Ekr6HsALNZC
zRJso/18lBpxUTeFhgnKezW0c+b0DkowGxf7yw9iGXVMon+7BpHLpksADIv6
8u9DD44K+vRBMdZhOGoM4aM3zN14mZuhb7myI3nohpmmfQvveBaEp8Mk0gRy
nGNOFZdq32/iSv5m3SMuJ1Y3xRwzCxpLY7wZpkthqe2v5vUokzV6AqNJg6hg
+ww008e+UsphFmvJek3B8lfO+i2ZTSmAuN27fHQC1zxI9c41APNap3VKxy1Z
QAjvJmEZxguhJoVayGdtu8KvEIi5SXdHHcFM/5jm88BWyYUp80XxqNOaSQKI
27lcPos3pWVkR/ff5E60fCTn11U5rwNVyZRXyeu1eM34vRVAf3uUV9W0h9xm
e0Q67e+qhkG++vGH+Q8xEVMSLiIkUAORMddbpaR7PBPt/0BHA9yPOHXW6G1D
3ILZAN2CTbEGqmlcZw1XhQ/TvGbQCO8muwqwu2kxKc0y8wBcNw6a3dibnYyI
h9sKItaZ6uJ1UIrSk2yOdX3Ulwt0f5anA/sm/R//+mXB0JLIuq67AWlxVTof
JwHNvk5KEEbd0konON0ISDudLIeoryNiRDI95nfM1DOtTHhzb4OGcVJdGanY
FJE277tZ3yPGKs+yKNro8+Y7dXnfKBcr1MHX4n/KovN9ZovA6DcSwtd8BsHk
FWVGdXN+QleYk6fTxvgjbTNR9rMbkK4VRi10PoyrczXVi3WA+HG9Mk14izm+
DRrB3SBOFjb09B4SjLJHPNWAzPbn6FMtY35XM3ryB3D5d5RrM404uFtofBJK
fqHTQzq7VC/WgDPU08y4gTlKGy8yMX56gbgcx4AqObp4864Ef72BcC/uKedH
Pe8tWfSwty1qSI43nZ66rjPTwJkBJwdbaKMb2j/ysRYHijtFu8vnQDkDGw8v
WgRoB9NpTUZqBiXShGMVyLWpfXkelnP71UJWa+olv7B2UH0noFHlNbDrSCIY
O8cr9fjSEy3IwIf9xVXxTV1bLaJXmsbsBVL/3hKBWvnz4Memk3R4UQYItfQU
56gP98DJzEcAE8KLJUFVllbkHzeC5xJ/2TLq03hx0ROCUcDpmaQaYCFZGZpu
AfwUAo1AzbsBIMSqLvOacwEDFEz68eQashKqP82T0xBblooS7oafsFf9Yn6J
/AGpT2jzg1i47gWk+TEwmS9wCyYXV6T/7xQXbg26YfXPiykFujqzGXyJY+xt
WGu2TUebNBcqqZ+p4qefguqwVksBDbhMA/bXj8XbO0uNBjhU0IbwG03/eMLK
PJZWzAMnHX7nyvZPfRZVKbLoMyYtXMW5rE7c2awNFRN26CwEEmTLK3f1qHBE
24Ybrs2Qb+RUqlhcqBWLpVFzKORH/tyaQ2DmvxWaoifjettd8DQKlk+9CVPS
c5KQirmj+IN4VN0zNgDK6QNy7oa3gEVJaK0lqrYuIt7gNVbqCgaY5Dpj6NcX
Ths/VXG0wWF9KMsreRUAZXfpd4QREGtiCd1L0jGLn85gwoIuBlVzyxrZRXym
s/tIadLAdh11CB9B5YNKd4YG8U7ruR4EAc5GkFTP9PJYTsVTRVCdauCj0IHL
hcrtaj2HhoGhOliiU7g19ZeG/wfoeoCWoyAymEXPT7vocL8Gp+wermxXqnHx
1JLdcijQdge9v9N1LajPZic0PzfgsrWQ8Gyz8Xw5YBAb5Mj3XbRlJZa0PQEl
GknlwAR8Di+yDfzcI4B7Pv7GEpwWgdOhRk2cd1OQmAkFW7rVOzbAsz/EuDkK
V9zKJfuC/0ttlVh2nuwbIfeLeyH6xARH2mIu645k/jKSZIh214vwKIvzQ18w
DgHBy8ox0pJzQXCx9STt+Y3bBlUXKIhYZ1KveCoe1ic60jVcUzTs/Ag33XjT
+1J5cny0YxZF+/cq1LWDMJHUduJZt/zJqmlcAXrfOu+ZZUd1roAEg3CLMXdw
yFLIXIHFxIoatuSrXKOLmKQTjU5u2hY6Ppw5bwqq1HnwTmzLq1ocrsEj9evg
O1tM9n1QaDr9J1d4lwbqN+Dj+0mXVoCuVB0OuDw4ry3DU4hHINbaZiVr/DHh
u3OUdmSSaKEukPVYERs9cfPCswEd+Z8DVy9XJLW7aO74K1Mv4k3cxrYFbKZU
I6C+SFMbM8aWDBn2NnUJ/iyYLbGP5t7P8y+lEcWoidNp92V1RznpSGtn93gg
Tm8WvyCx9zPe3XW0Tc18IRNNTRbIr0/2+/Rp57oW7G990M286uww5kHPYLIP
oKlQyaocQNpaNH5IKL5EdFNjXBAV2U8B3vcMdTm7m7cvzxcbfQ58tY+XK4+K
78PYZSRK36UGtZJqvZGSVYGjaMoWpt+hbXAvG+eoyHgqlARw4CCptdLLVmvW
cS+vfUoN1VaeBAegxhXK89X7G1ad14pSC4zBXxRXxlQI/s9SRlyyCLLA5MbQ
P6hB3FkkJLRW/lONcI+L/XLMbAPBB0+b3+MiqSbkDSjpe8vQBO0OrUy7Yj1t
LfYBo5CzkjWAxyzbGCz2CD9suZjwiHabdKhbfFT7t3v6Ut/R1BTzLMS8j51x
roOCSuuu2HLO2Gs74Kqn2krXn+VOaWPiZrQrGylvwULliKWlYoE+gNRnEbY/
6K2ssiDwyD4maB3UBxMiv0l9vcm8UVPmB7FS1SGu7NAZ659C3shw32od1Ysg
5c+HzS6bFOxCp5atOq/sjEO4ylmBYdwRJk2S1R5SG21E/NawtUTqG6wWKih7
0sJNVl3tOssuxLpwVpEalgx0lHzwlHeCgkVb1SWc7MSpm/moh6ukG4IEMz/H
fns+rozqoIS1JAwWfb0J7dctzET3CtdyPkgWt79Vh7ukSk9i3i9c/y8LkSc2
EP3xAoTZqloxcuy0t8TJZC+2c8QarGkAKeDuHd4sB945UMRuu03PA8CzIUaE
dcr9fdYK/ZdJ+nuYhep+Z7V1U2rIfJEsdkbL7vRACSJ9KBmQ0yrZnr61kU1r
uCRLy86+Yl2X37cD6AK94kGCxtGzLbbf2aQyYSuqRzsGVu+LeSLH5h1oALCK
jy+poufy03RuD0Xi2YYnkvryTjuZYAMVk3rnMrGxU52yOM6ABzTaitBcanzu
FokWqu6SEcPKdyR8qydu4Yy3kYtDkLpW0dIxSj3+AacE4nkXnV2u1yM+yVCu
Wvb6bsIUoLUU0lg9SwT6Ms24q2SPzrxD7J47BTsKjB80aOdsZhpOE9F23gZp
fMWr82CpozlAsPhvhyKihjayIcNY0wBvQEZ9I8CYlXojjqlRFampLpdCCapx
m5BKRYZQTtclq/a/9s4+svIEybToj+grohuENoPgZ+6k+MD4k9m8KnL8gR1P
W1wCDMXMFMaK7yj5gl392iFxggOTmCEci8/4+RxNnRy4KrG6sE3VWEJ7YCSR
+HWCujYaXSFZ0kY5tGweqDtc3LSNzXwMRhQK9pNj3YFM6keMFMXA9TLCoIMl
pKopSRXCrKlOfdpGtQLZbWkH1c7FPdmE8TJk1vjssjkZTosiOQOmjxtPWpBs
BUi0S6Gjc0l6g159HU7DxFB/6vZ82v6UvhhPSW7I4KKOY79kpHMTP1WzJ6H4
8byLhq0kKYoTg1eTMY7W3k1A5KEhSmhY8oD+8CM353e7vwgBC3+NDtkMB5Kt
Ee1kpgMuqg2zwi8K4+KGUN/4lNXKECJNzwXjAS3aQMihaBF3AvmdL5WwiVAp
REljEO6nQ98t9EmXkyWfy/w6g3x8SBTHtCTr7EzHFmfR8PhvIr6F7OmR6Olb
9wqSJn1zbcvD5F7buKbgaFeOF89meGmSCVjVbFHka+Xce26oyXt1MekAvONH
qGusArT7nRJgNmK8EM945Qr/pofOtmZiRbiF5IPaiUUYJm6iuVnYNqm4oFh7
s079b0siE4LIKs0TeJJCuJrZT2wjnaKrtwuaK37VsDUd2pEbe5gz4LnFraKd
q3B7fp7u4PGUW4v148TMmjRQxVQHA7wGgAhGy6IRLIYfoOBm0Y4wmmU8Rv5j
QaycqJDyek+WAs/eRfgWp9ye2cWE4vfQASLhH1aGCclyDn6YB8h8rHv8iA9t
uokHcAN0WBIvbmK6QeJ5ZN21lseAwar/QpQXoI+OX+pp1eiuBoZjOQypsznu
SHDW1uvik+hA9XWScTsAw3JkD0T2WYOuvH4PmOIZrpiRr+/Amd3ibVLY12b+
UJuCTve3eqGxGFcLwY5O7YPL0XRcK5DxiRFdoI7xmd926rmTpKJ6p4GQREg4
tjA6N3/x3+ysL3jifwexrqV6UAMPr+mH52vXEIUXkpxptgPHeuolIASfiMdH
o22oaviMOAb8ZM8lz4zLW21AS7+y/PNKuwEqNlsRJCHw4fwMKVMwWfY6xCX7
Vhu8wM78NuiWLjktKhjE9Kc/OoMCMTkJnQeAA1R8x/Pn17sHw9WIFiQOzBMD
OrOw/fXNwWq6uEGwW+I1hbvQKzLqG9A4q8sVUrR/DRGv/Nv6SQhv//crioJO
ehucYUM6jRMGkom3u58abtduWU5mw0wYPj4qMo739aKNPRKwyweHzNSyzDJT
vlY+iDyLA8M3Ikk5sFdo79ZaI3Ii026n7c6GJWVj5AJzCYp+5JNWuJPZczxt
cBDkE6Pif5x9zisVAYxvf+Dvb2YatxGnA1VNsDhxjE/jEOHDPHihR33qeSij
iUurdnaShh/WA9f/ugzxNftitshMuFcVwmR63fC4PdalXfzoF8Tx4HdN647+
9QoITKsxAIQ+sXBjMQB728cu4jWt3W+NF6TC1Cq+4Mfd28usoLshP58YfwQ9
SRcaI/Y+3rycZijeU7KCEq8pXkZczKmVtTzBUvZJoIxRtWeq8U/EPXQW9MA9
lHgbUZf8tj5GrzUecEs5coLc0eD3GxVZMJNrGCggxxxG3d8/7HjEkFzqUxah
OGvIMQO8oP9GFLbnh8hiQnpwRpmIgWQ14TYbBVKz4peRfZWiaMWmfyvoIipz
nXRfHv9Ey/fAiFXW2l9BP+BHiy6lDuLXEA3fFpG2JaHxMijn8e+HKxPaHmFT
qyv0DdYbzGjnu7zrTzH1GEkqRQfll0KB+TCT4xx8MLhiR0UhUJx+JT1KWOOB
8xNU7AJJMMXSF2askhEuiKJm/0GHd81t/C4uRlRdRqH0xmE3Lra0t4+goAUL
SSJdHS7RBACaBy7mEmXv6kioAPxrQxq/tWW9Hj5Dbqv3IxY4cHQExwvheBNh
EXb4aDYBudKnJ7dsHdN7OLkQHRkNFwUbgEU4GlhTA0FDKI9OJa/scCi7EbIc
Dnjk91Wu1HFF+U30TuE2EY+/ZtTG5tg57TckH1TMSZ+OxgPMTIC5NyzmLUu8
AS8zojsG1fT36dMzQQk+xGb0uvPDEPnPHq8fDDflZ0W2nyIGn8RHhCqhVxLy
j3WntHkTPZYtzUbN6t6j/+TgQVA7UrSV3cJnQSTl2FRbeSMlXI32pVyFYIqH
4fjuitKKwjEnzOxAMX0o051W7XzMbeM9wYBOltseb3anm+nnunaafIg1dWbQ
3Hfcz1VUL4/Bn1tgK0GlcIoj/Ele3rJ1qETisvjq7NG97K2A3909Ax5iWWQZ
lfH/G4x6WBLLkfup8hZGgrQ5oR1iVIQvT4NFCI+abhV2h+xKwTKfebT1yKVd
wtYP2CBWvllmQBR5o82J+enzMjkzTZM1MdN7nogZLoIC03wFJzXLAwdG0EkE
n9MCdzb1xyO0SuxeJs/9h/EG9Qy5VPqXuhhwg08udo6XoBT0iM4QsTX0mQOR
VC29og1T8c+hnPmyZQ22VevYLxlw0Q6b6WhFk61wCePXdhkf3HlOzpvXMNKx
YOoP79B4Y1WQY1dQr28YAA9St5TEyEgeee6P2C15taEHi73B7ljwQTsZcXgH
Y3+/4TJAur6jttGQPeytbR8rnPeAeO9XkoP+RekpJB/0j5fFDnSERP35d/tB
CU4Af6+13V8LZH5QBpdQCHthIIIbK5iPmFoezKK+qFykVfvfICaJvOdBXyuG
WUC5HewQbDDIpZtxpGSfWSQBLpAe9ORP6Gqsb2pJCPCbl5tY/Ag7O/HCZjCw
JLjKM4L8/nXhokI5jOHYFWkyMQW/ZjeYT+mYlvzC/00/9f+CloyPMg9wPmbc
CHYcsJAUqv9mQUAQcgcEu/WEjEulfNfK6vK0S/2C5DkgAI0IF1yZF2RASNDJ
jcVuUfLih7rWnjDbHW0/m697G5mZZagK12BvzNfJOkAWZhP+FxtlmdJcLAWT
bEC5O9VjWzDNMX61moVyNnrWdh7yOIeuxxdWDade+ZiN7kyG6ziPDYFZlZvo
Dzz+mTKe9Gg9t1eYn4OiMiWYhsgCRmW1pgaTzDM8RrZNbnaguAVFpFoECK1J
4Ub+6LLMCMdilz5daxhPIzVm3ThDItq3rrq+k5EJsl/XHhSJszWGbg7J2qJ9
wtYVXSzupJJGOXEfmms6CqDDjrmbJhr9Y1mM4wY3pjZ/gTP7iQSkfm2MNvjL
QaxifgMO+Dovru9bIuzQ90hD4YvxBEMKDCSVxkEN0yBI4Oax29on6HJmOX+g
1wEim+A0rC6c4REOdhx5qTIkIetNG36nHOn2hGMcpjFptlObsWt9m1c2Xi/d
moC4o31ufdx8E3VQsvAKbcpnNy7ZM+8N/70bTu2ATCIRWwMTM0h+znXHcgwD
FW/xt2wjLtgeqQHS0ISsVxYoYTd6y1lApiIAs4P6PiulnMsd3X5KTqImJedY
oFACSFC9xHA+YgS6i045lt6wYPcYGtdlIE+0V2ZBy5DU4KaP2kiZSxfRaACy
e5Oal1/Vxfl/7kh6bFNhW0/GF4It7WX4v89Hrm005Yvwz7f9dXb2JrHfM38I
f3g0FMPvLgDyc3WsdZoTOOLSzbYc6KCpCgvClyozwSHqt343HOITUxbo41Vg
OqqgaO1bV0MD0o9AYDOMw20JyoZpzfNPHOCjIqjuuW2IbrKcnT2rOEE/Sr/b
3cCRLHz3ERCvv1pwCFFle34yjmS9h2nfrTxWXYSTi6qzGTdWQcTqKhMIGc/Y
ylUpeii/61gJ/eiBlm94TlOP6NORIGYGo62tbtbcA0yS7VNDPJo5hZbOdl8j
mM1Pj5U9yuslvLq2jFPmso+EYXJy9CpkEbGVd3v2NSs+0+MPhvzWrky0gFFI
rXKN3IRdS30GdQ2CCXQJS6N3U6ohoWL339T83l6MWPBkeks5LQmQVDfcasI+
/iK8ig02Td6DdJxVDJKLhLQ4iaZH+iVMU4bpGnqwe+zirr0tEUQ9P0O1BD64
+oN6m8U3n1rurJtcn4NUITOhNWPGeCwOySka6eySr7q8XMjAkQQb7z5VAnLO
7Mjl+ukhDTRb6FIjWIVTNMKeptqzDML/UzrZtNsaQCE79plMCFohV+8JToRF
ZkEkyPullB4gZrt4wJVrvmGpQ/Akp5zDM/uTOA3EUK/iaxfRxr6mD/JjYFl8
gYPLi3ikSGJX9P3dM5fsWkqQ7yyXbY+0QOeXjM+ZAbzRorWvcmbI5aysoWos
eoQ5RKALhzfIlwf9uAVblVmJWclMzeIoEAjcBkyirWIEv39S6VqN6wS2VCJn
KlN6LsAGv1oxVR0ev4C7MS3uzhoJ+vjltql7snlcHWRMVP2EXkQid1ilnUr0
IBYR41kelW4b7EkymqVM7J5pPIXLH49pkN2cHZp2f95nxTGEyEKlLcsbNFzs
40/txxUis82EUObz7IEnw6AwhNSkwGL3pKr7UmEKi4KNYCu8m5Zd5h7Hbls5
WReQyUD6yv/qCY0Kb/pLbSe1r57wcfFoee2Gje32gS4f05M4QBW2kOPdZSDE
JsUZhqmsgheNJSPvNyJd/nWeaQZme2ImCJPnkfDwEgSPfqe6YQ9yV3Pi4x4J
bWSpEl88yLSnqz778mdaCJzJkYg+0E/J4nvjSOkDRTL9mc0KvGO+bxUCypTW
G2Pbhr55fiIxt9925nvICZ9r1htIdTfzjD/i/2drntuF0NLtimSmH6lhJqmw
DJp0j04pn3HUXiheU775A0hkFjjuD+4GtZBbzql6Fq2WUqs19zEUPlKYWmPC
NMD/8r06yYRqc3I5/1VH+ETtsbt8BfyiAW9a5XaUD9A6ZM3/xz5TIwtZkn69
nm4f+yDbYcAPCdIrqafnnzYg5Q8AeT1jc6G2wVn5cupKJIbJTrMgK9oE9iD6
NNSS7IjhnYmY9waYrjJyXDHQZVygZcAQh98cQT2dI7qoudm01ZzLOEkCPbYK
tTfyF2o7sgv/gkUUrPB3TI++/vonWxPv4KTHbpQjEqNZ0HcqBsaMP7hJGwga
Cf9W41EjY2wrwvYxlwnzP4xdG3ciCJpIBbKtOYwXJMZue8sfEIe7Dn7++6mT
NCn8t5rOPRTXmbqLPFezGGROcZejBr8KIUV9U/QE9oJC6wDevsZhy0r1JT3Q
0MnyzxMnwBH8VTOiNgNK1IEfcDPq/vcU9Rbg+Jxv8AI+2TegE8wDVFiPxRB1
utbYLI6ODKnUjkt6PW8KFzF04M0r+3+YKAFZKdTtw1XcFAmX4NJBZ3tyeAQ7
YusN2+VXW3di+hjyq8de04JOfsDnFOYD2bm8h8+T1/aRWTFfZ4JejgAXQ1ZM
WNtknM8ye0m0/teFm2M7olTpT81pEmuDtM5WJWSBoDgkwy4YmGJWLrjEqjKt
uezYttXAzAY57BGNr0ik7gqfwoli43TD+WMhNRakcgaiO4WQTitU0AU2VJfC
pbhyaOGxZywxezFKgeLcJcEnS4kg1XE4XQv0xeslELuFDjRYomHxsVIoX44F
2+9FnuzrfZTNyUEpLafh7PD/yEChzRNVWlwH1glhmnrdu+/d5dRhSA4QtnKz
cPuW5C0RwSD8JnIb43q7/zwZ5mR1p2kStG1Raewnvl61xVw4csGm4Z9fCcwf
zr+vdtSnQG5ttTZbzFkk2p1FtmFFPMk4Nf49Q56B8kMo5S6AvL0RWqAS2BbT
JqVhQnc4jqdfd3ICy3NnMOQ66vP/4aYBwNQl6RrSBFd97qZYxX9f/fJGJLLz
mKuG5X4LMmDahSR4ikI8Z02QkQ2GUkI0lKl8rIxCG6uMAq4DW7iIznFLU/ZQ
bdenvgAVpmjW/we3I1XFCOgGLoKj4oZVpUthkWyDskeQYYROxVhNpMuvgAgz
WBmYgN1w+TmuxLzCcxXz0fcid70Ev28pNM6fjN49d/yULZragU0pfkp45psK
wBaxjgRMJ8XyF9698R1SuTDe4VoLBHavjXpmZWuL5R0ZM7zzRW0TJB64offJ
aN0gTYF0xX/9+CN59CQI2tPN8JHXshrvSAiQsFa7mkzvyXaTHlC61nkJpgcV
AcLyJeXhES8okhtOyCVkQRItt6tENoWkR1U5XHVbBHVeJd4nbl4qbGGGhtjk
5hmP9Wz6bSWE6AOI+H69E4CiaNa5XP6R+N+MPcD8Hu7FrRvO1XgF0bU36lG2
/xbBiZfBtNo12VcLxTZ61odPpTDtOndBjYtheXK+BqRLRMc3r/F28SSbh7sD
lQnnzrqDvsrhzrxnQ3+5+pOtV49zgHn5/l9VbLxsyhQhhhSRjINSoe6tznqk
S0pvL/v6daq0U/NIedqRzoGwMRTRQXTYAD6aGvS18y76wcxiea1EPeBoOmzX
NnW/aE6zLZio9d8JsWKYd2yIueCOF2Up6OsC8i1jS7Iu5EzuWSrR+Bdw6oTX
N2qcQX/iImtx1BFINz30E3a0Ocv4TgBuDDaAtUCGHAK6lQ/EKerK8DW3NLum
89EXBr5Z3LNjsWLcGZaHcOBzBmhkCB2Xd3LOHOc1ZG8AaWCt4YwopPXZSz4v
ur2CMhFit1FKX8TVX+yX6kgZwS9OVl/dTO+53XxlcwQu0ouNm42uYf8wpsJt
B4rR+tgheVyQ5GmXPl/qNqVigEflZMLUpkYp0x/uLUnuEqQuu1WvCCzV61xi
DoCcbQ93Cn39djJmgoBBgcYSfzTicdGBheRA/LgfAe0BSu+w4opE4iNMe4j7
UcW0cEfl4h8b4Golmy+D7O9ifakNG0m5Zs/iIMp2fFD/FreCobQnmhq6OPcr
4kw+Uug6cuA5dtAcjz+fcTfB9/5npfSNpWiuOpY3p3GxWhDLWky4EzhUCZfK
8jlJ4E9N4atRJaUGxdjCOiioFbnzYvSUcomdcjoRkK73+IKUBlix7Xnd9cP6
LGq7xJdJ0jxOTX6H2vOYbHOwLsUODDBCwYxtntNRBuVg+mKYuH3BJm53/dd/
aaORGVAkJ3oS6KqzX9FalssQzYk43jIPhFcT3QHFU7UYusEj8C1OhHvFijdJ
nwCPOEsxeY8Q6ZKEH+D94pObTAIgfd9CRuHEUXB8Q+5CWmgTSud/lDZnxg1m
2Vt6FOAkVVO7UAPvRgrNij09V0mk5satuTwW8AEZ9xNr3RrrgUgkIeRXBXJs
Rm+B9bmbai2wYS8iME4EarNeZhMLqpSZFM9+9MQq41643RfwnjeKxG7YOwXC
Ub4lFcHambRNDbVOr0JOOj+54wmaxG30nPxwgtEpWMWobjxCsbZ4RncvwmSW
0QkkgZ9IvxtL4LzFLGaIIiBDHYLUX4qU6C7BFOSZV254sqT7sTqXhgt1sDNQ
krSVZKs5AqTVzeS9fgfCBW4NnuUaC/UxKkjOFpvPp7Hz+JjKd0vkTcwNBPkX
pHnzpu9DYcKUG02BJX4IpsnQ9r5IWkZPkl1HGPZsWwh5daJEkwJ1osF1hHUY
yVDFfXpdt6mO8HH09+uuxywwwZKIYiHjDpLIjRIqUjXammMFbsRV/rIfcpQN
R4wF+MTno4a7Og+vkysJWygcxAcRHNctrBS6cnqF2GE7D45v1Fhf5mBri0da
7qfKSScmYMEiYoLb+TxrUqVe9kOAobZio/ntnrW+EG2lB6+BRICyDm+U+0pd
FvgahnTNR1l80PAX4hr2gVakPI8cfEjLnukzBz5aCS1il0AipVvQCS6xG6aa
vumvN+a2vxKr4/pTgrUAX7R5GrkT1+8pJkCIAzymCAHzlnCaCjtWk6xMFyw0
C/yU/3eB7R9G97Mcmm0f6i5KYAJzW2mAxi0wPRoAX8iPYQ1LWbm9bPDmJWRy
o+X2h0q6fNSG7jLLzsOe+fAI3hF/N2csz8T/KOL/KqQWtwM1l0V1wvaTPNYg
W0pL0xW8VS/F3mZL/PDfjr89Zlg4PfBSlua8qs1uX3oh2OIS8rAzF0G45kuv
pz5IhhWcG9sD7KPRq8EGCbChjmC+u5nXEhGYpTPLhrIwjq/pdNqtX4fJDPBa
gGBCsfnwd8t2+WfcgXjtNH5ReRmUx8Q06KJZYiC2bKKID69z2K4jswpal+hV
XsYSVEErkyohTm44JZtTrPKy7OZzZj3zpfa+WoQbx6NXY3Xfp+rRIGAGrydk
WbiBkE6mW7/sGUxQN90CSwdDZBd0lZH7QDtq6P93JtnI15IvZZ2Uiq1EIXG1
3/kXtozRD1RwA4fo5v2OHjMOiDOugRMBCHcJamupiZX2LiiFmG+9oKYafZqV
CEy/mEpcv1Ajwm0fVJjO/REOiMRyo45C7y+OGieCJqJYKOSUgJsV5VKaSiEp
lzYSPwIdz9ECX2JzTi8pK7rPSDAbb+qczHwmVTZxxnbYgJtnD97CM0Bhc/BX
WL/xDrBx1A036QCI04uE97ojYhzZAC8xCqzsJ3C4ee4b8zVg+1+wWNVHmO+7
+bWhuoOC9DOKxPKoNKFVCOSs2DGUCIUImHOPxCJyfhNMxN2YCumWiVBAZ9kQ
nbd9n4a0B4U8TChY1/XVLSwj54S7Ho+2xEgK5Cq/WK95AtmOKxC1VsNSPZWW
lSae1IZ7k96gCVFOTd472PNB2XbZB1EAQyv0jBdDNLnC6tisAuNTK85iHWLq
RvV+fdeepxywA3mgnJEUnb5bs1SEQdHkzYWJgz6xmz566933duPBKooAhhXJ
QP+TWBWxFVfkHXNQCOzd2fSsqdfXYMi9brSIhL0PQzwsTxAkHa150WF4Hnen
IMKkIsjf9qkiQFKDiuykqD5pecgXBhbF89kHhtXHd9vHLZcNTybKxCqQwMqr
5/VVPaLjtlc35KWak3vf4OXgA5cZyRflQ+fWuW4ws4ur8zQLpCsTUZE4eYpZ
MqqvboA/qeLUzYiQH98vQuHVsCh/iG2NyiT84Ll5VoRn6UmflVMLeuBOSVtL
787JeWqqZ1oDpWk7D42FieYKoCsODbeTemFVFzqJH5FeUYS383mw1a2923yE
wPs+M/vm3OvUfoG2XCwvqIDJutglgVm/rnp8fjqrNLd7fuRsnnQrF4hC1Czs
UCqiqawPYSqCQD+3muywc0CJDOzoQjqrM1wqWU6SKcHm9HYfUY9DUt2wvryK
mJFp26mwILQK5LeD4I9rA4zejVSe1+O6kfIaTGm0K1codesZP98++T/gIq9X
2ceJ/BgoNoB7tAZhCFLjfF0GGic6eBg3xUPa8SFtz72EqXIQLnfi6zRgBBdB
e+BWcDnPQ+fz6hVQmFwb541+pdTK+dYpDzyEIUqkEeKteX5RXgbyQy6o7LGc
/vSaoqOWqqjvVRtfiGVtYvwP/HXs98g/17xQvG9AB/jZ7dvOlghcnVpHVKCJ
TxSQ9SjXxyCGOIsbsfbqbvsscZDu7I6ixOk49mR6Jp+w49MNNhlbuwgbkACm
u2Bdb4IEy/b42GoahgvtrOKMuHY393ATt2QsAIQ3m4ocpvI2ig2K6ry+68eY
lFG0QjuilwjlFhM0Y0Haomne3GVaxoIhMAnwOjk71qlxmqZOmPEb3ZDSdQ5Y
K/DM0uBu3hj2NUqRCVZ1d/+UJ+MakKjWWMdFWibMZjMoP+qe9xNnbGQp3ryd
uRJajw7Pyr0eoYwtxUv2ufmyOfGwEzmYbO9wV13Vo/dG9GSzuqCfAIHS2XQZ
GC9TadfuyFakU5bzy5hyqUdsYQekgPSmSbtC4jRBmTPgwJAsoT9IMLYGk0Td
kITjXuYdTPrwcoF64l9Iorv8vkYHECgCGIslwhVQz6tHwvSYi3J4JzJTvWRX
OGr7NmQPrr54LiFeieJZjiwVhy6QoYNyBOzbeu0rG2ZwQX8xmC55Nw8PVAXy
LDA6p09eEOJzRyJi/DQL78Ck4teq6JunPMe4PUjpUk0lq0Q3LVNmX2axFBoe
7eumFaIK8fSprhx83jLEJe1zaEsog7ATKFxH4jvay/fbHahB7V5KPz2wHqNi
g4qv/EaJQ0ooyEANe7hcjqVDaPFZveMZUYFF6/jQ0XIK+ZSw51G305iXaWkg
+J+h8pq14oTe6bqjojYBs0ZBf1DXLPXH+4aWkgl4Nit4k4zXjF4JZla+DSIT
zOhw85RU9dulH3qXeC77OGvW/zOrR5Top0V1No/eH7MUqtTPPIs+OaE87wIY
ACGt2kUg2ehRRRkG0BtBhyp0X7lRNtkQt/uHXMDrV89EJCh7Gl5mccR6ynpk
a+6Z2qlM876IRXHcg5WtmaCbUdGPEk1fKKry9/vQmIqtxGlZ5XdWkpi/0jaJ
3Ja0+0phZ/bUy0Y071fCeFssbfBZuvrcwLWCBLLdsc9nPRxnUtdQ7+JdrqJZ
2J0P8oPxz4Iy+f+g6sZUK15telfIK4xmICSs4p0MoRTyYGAgHtb/05IpnGOz
+wRztjeEzBJ3C2gWQNyMYXQ5MYLVh1Z49f2qTdr0Es6aJMWSR9rnPLC11PRq
6CB197udbG9OUP2qoMUM45Emg1JZp/Aiob7yDejyR9R3yXusB7cpc79/nU8V
BhOeA7oZWPVEJcAL+y1EvxaLvAn5ToVX9zcXBpvitrED4TNa0BeWWGFUHwT5
QcslDIrF5qLl1MwH2A9tqfL2tnQ6dE2OtylykTs1UekhBlMbG8BMOkppujRw
NUl89zCI/aCxeujfIB75TMNT6/6nXSmsjvn0BcoErvmb2R/iea+qGtpHzGnv
Rj3LQ9MM4LXMdgWCy7xhgv/WBIyrvJczW17sn6f9PXGizyUDgN3Bk/a/cNr3
kMXbbMlrsER1JmYu/P0Cdxq/T6J/62+p3azYIxdpsBgLD+BJYRJluuAOaQED
khnVWOhRcgFmCsq3obUG/O6eRo9NeYMqqNBIu51VUmCF7SyvQaCNYIAbW0S/
PURQVYq7JCymN6mmvPXxM+80u66+T6lY+X9Ry10TX2r4fAP6kk2rnUMifsm0
UvREoXTXBsphwrURwcgJYdE9N8D9i5aJp506KPi5Nfh4ZUJawP6hskvuRRj7
MrI6++rqbq1mJuLOoFEp9hsPW0Z7C7EiYaTCkIzyBRQdeMxrrfNZfZth1G4z
ZnE1aJtWFbNWgdJtD9R89qkopgdTEn3/Vwkk6ieGbgkEg56/c1Nj7wbLUySC
l8Aw1EjEG3Q+K5gnmmVcRGcr4jT3JOMT5zREUQENOjD6MXpslwMWV2SmKCBe
zgwM0PTPX1hOBK9XPNsjjvY7W6EiiURXr5vXiktMnbPi8UlTW5rAtuveQ/85
Sd0lhy8Jg1J1sj00pIySTr/HJfY0WQSOEjcoInHK36xvUbRtSCqwHRqPOLjQ
TILXIoDjMpYW8h+q549T5/3mZehIW9MK9gR+/DwEbc6ws6H0Nj3eFgP7B18B
717NPH+MpIcTRCbaTmgf4smDu1wc5zl8h6SsvUkKQVOJscwn5f0KyAW9D/It
l76qC5da24HOCMDqihUF2vtUHFZTx/WewQB+E2IIkqFcE2aZcNigUITeIRES
bZA7k+mHA+EKJTMxmDrRBZ4TTZuB1nwfyOKIjHyJ3Xq6AGXpISU46MgupXwy
TCIt

`pragma protect end_protected
