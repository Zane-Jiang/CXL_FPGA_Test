// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vWU7DTkMHggBTd86cZBuvBMA9X6g9BOk8WvZk6p+T5ufhL4p8mR+uDmLb9sx7O4tO0OqF2S3tm2Y
EnRoCxdGsG25gQeJF3g9/lHex9dwQqWYvUVEaP2I5wAmhFNZoYG73TYeWBuE3q8i8BBavuoAu9qy
VVdZd+MY9j/yXqVhHZ88Z/KF901pGIvzbDFSpNEQXgb626IzporpMbYAojTwD6UdgXJWuSnSa1ln
ZtTzkfLD1KKPzaQmXehDKtaUdmgUsoR72zVidN5QcmdAscx8ORuoaOZ8pqF8QJuM37Wu1+ZtqjQ4
yB02OJ0iasIonEliTwMkBF+etohEZsOOAfG/4A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10000)
HWNRZnRNvNzNBq8/AMQcEgYAMA6pCBFMboLBFyOBwOCVjzRATCOq9V5cLpbVWpJiF35vUldgGigB
Y1QUN51vCmzgCYdFFCR/CB2JCe7b2G7G0dSmxjMUpbvQMJQvaa5BXAelbXBbErtbyi4fI/4ws7Wd
40Rpk9odqjKdyJHZWY1ldk0KMUlaUkZVyJNCAWHL4O5SjyWdMmS4TltQJjroKQ61rW7bnqpb67/I
sZUoHB0KHfVl3gFVu4rOhHlxnFxn0rikODwwtsI9uTPO5pVLw3UdF/MLhwogOf5l+Ay4AMgj9A5G
XHdiQJlaQyN4Gzz56Eg6kr4gJTITELwW11thO8aE0tQsTgqRzw4rwufxHhex8EnpTUivUu8w8uQn
jRGY4sHdjWMT9e/NgpkTfnwYsXrJFD/EfDcVp1uErlz5MC2zmn3fEXGoz7qrIgvqlS3ArnQK08Ox
3b5QgAblq87bZMGLWLVmVF2oPwWOwLxOhnSR0cwfB5BcSrqYpwkIKYetOzRzGnQvyse1PvVBhMO0
ZVVdr4DjRG2wVq0e/5F45ybK74kPS8SfAqpEwmR27leBHb/Tw7AwJsiwseYvMMQE82Iqbj+hYVMU
OQIl9e/dMoBjNlaEV3M0RD8sxwCUEBNfUPGCRjzUCnMi9DhhURCAGXeg1vAMaC6s9npEZTc/Ie90
vrq0vlLet0C8ckbSSyJ9/v3yn0Ypk5fqI+X5q2EIWciBHiL7oOTgQ6LzErz+ePv3ys8eoiv9UzaG
nvKH+4cVozmtQZVUAIikIQmWPu9mrmE+oRDnnjXsJkkH9O6ycThlfMFFMKmjTwwckAxlgNSIgBms
XK0YP+aW19SHK37lpgigCcYEKAGQf0VueijJsgX8rq+p9cORIFHbkDTcEVmsTDpAVcbo6cwOhKUV
Z6Kd3tD8doLnsYbY70oFSxqWx86KeMWHLLa1jeFJHPuQzLMOVJsiKj8gbBT3XDMFq1nETvvWMLRH
SOjZmmrZ3upDbdrJrgv5mkpMuPmcJetz11sF2f9kWKaOok0U1AUO2iQuiUt9wFIkoDOz27eiZmhU
nfH7IcG2wB5TOoAFVRblojgypzVv1IuKB3OnmRM6FfXxd8e10UXpycSagqQblnSupM3waUTjPdt8
SHgXGRSl5ZoR10IiwnPppvowIQGOQLHuBBli+Asl6nTGEV0wPntHHrIo2IdQckKAImCin1Mju4ZH
r1jl2VOJ/3pgjxF87K+BmqSDatNCggWx7kkT7UVhKz19OFDZjWMFSIBROVwYTfQAobueuly0TXXW
a2Vmk7qVO2/B6gmre/xJ5/wDbedi6ihUfgj0nq+k3K+dRTDQuPI3/vUel4kNvAvutuc65Ec5uiF3
t+i0/e/ddBM5YLweKjb/2pVlo962SPNlioqjGOuk/NgOhM6p7bnB7gwsEqDJNjwoqPXz+FwpwHMa
LKXrgRbMQMFsfOgeg4pIhskSFfJtAYBeqVmU/yzIzHBtbccmet5SVU09Csz6BW3rCiDnYr7XKRXy
3LT0XtB+3O0Y41UekMk/fOtkD39cvx3Xj//TXQhnJRf+YLqaLsG8/W2Fc4X84jpkpLKOzwtBxCUW
+2fRiCXt/BaAZAyjTUIuC3YgyyDD1O85cwP3AvjMTZxISSdwXIoPFunh8YQxRuNrbqgWmfnsikKM
B8wMOIrG2BQUteRiB+YF16APy23ox54ZcTOOObIgl4hVyGGKIUCr+Rbcuiu6B7XnFCYUcGHJ0xb9
Q6O/4sEy8u4GmqCkMOcesQSK7HuzfGamofpOCuCkt7FVeCIj/00EZrOSzUfmSD5NNSS2zzqBWZO6
B7vXv8Xnk6IC59XiHIX2/8lLCqM01SVA9cWH/t71zVvTJR4k+KLZJZpjdEZ8tC626jZR/3Q44jks
jL55vfGhANFXCnWg1y1mz45Xm/63dEv68PnMvX6a+2lXkfYoAIXLXsGoBM1eXfv5XbuO6E18gwI2
jo7vAveXiOeuCKlPeq7jMZl40ZBZjyOdSkyUcvvRklDog6MvbtBNCb5PHi2UVr2iqo5Y3eqEOrZV
K6FGqbzLk//enfGpAn+Cu7vqFKIkUTu9xxk1jzzOFCBV3uWClKRP/Z8YsmVSZ2Jl5K07iEzbUe91
HDTlBm2qVvyx1PcT4WB8uz2e036vv1AcyyKMU/eP/ME45V54M3bZhdRWB4lMr0VF6vxVE73L/YzN
Yb9sUkkW4XgBbtQE35Vnv+SUHpFIqaQ3Xg0Q/SrvtyAbITK1E/agfw4dQBV0gN/IDvzW+zxoF/Nz
VLVVDQwleWJ7VHfkWHHFPoUcuL0MNzuqOPe8Zj6H+RkPPNUzDDNxMvgUAcL2YCNxHyqOHyVqPoWJ
irFPzx+XCYNuwUGlO/EY6t7Jyn9CMXoTvYvYUa1VlIFr88bMjBOQffLeUAS7zwPoA7evUGj/kTla
/qbz+rNslk+Q5HnwF9eAI9y2vpzmfmSlV/ebjnHcS/FGySdpQrhTCgpe9+FlWRAzLevXSZ/pXAnS
/mfkoNl5aebMm63GGUC99MFwjqfZ7GTgZH7SfcjsxhsAn5OwzIAdIAB4d77oYQ0lkOY6ZtRT7dHb
DJo+h4G03T4RVU5i5Kip+ArkoJwXnFhgyFa/U4hFj0TC7EyjsRB1eQ+VHvxL6n/BLEixzV77iGoL
TmSmZN46qOZgFCli5Ww3eCnUqGRjtbqFhRT7vO0vcxPWIv5ikSnuChDd9xcMCOPYuv9wZnjQO13p
VWHVxlOuzi6xlnWrr7SKTCP0l+f+Xv0z506JYDcIfUPtiBnYVxd1XMLTvILXgvuCZMuxodK+Oq0W
clWw1dJ4dA/DWe9cOI9zFzI/AhWyKlT9TiiG6/XPB5rgCQr3G6JELZQWD7XEVXRiKygwvStFYOeN
ftB+Pfz18wWRctxp7wY4PBE+h050dpG916ijfumuoyV6F64pIjdAV+riEG0QxMyhtZawIP/MhKbr
gr2bWiP8FLMu4pqQfKTkO3bUBWwUMEcRhd3R3XpsLj5faV0EXxhvu/p8a6OHL3jqE2iFFnY0HVPz
mY3+RnQc727BhNOhR38y0lJQhBN3uWKm4Ac424MHy2SKLMdRVi0drTBCh5lRRMjywDfYsimLJmy0
cS+N7edkYTi67VMsX7CS3nACkDzs6UckWm/IMiHnXMNE3boeygV/GZckkq7ULOFxv16gUhnnZU+n
7sHQvpQ9PYpq1xQo0ox7VLZmE8a2Mp1AKn7LAfCGhjatJhFLNQDTZABxyE1wMCtVx+n5iOEpJWO6
OrEbwcZgVGzIWPJ7n5dXFZHUH/+j2Euwz4mBEIhJL6BsbxgljE27U243DQ3uFRb1PQTaHJe0CvI4
yQzu7TVl9yi5pQ24fW11RBzwF01qAkujin2pbsLWAze9Isj06OoWPjIt5t2LuErNIeaU3eRGxP8Z
u2ay8qVmnEEEz//fIkNdDjUxnNnbyMupjSDvTMrQlJOvlSvtCQQHPVA8Ghv+nPBD2k8+OMji7Y23
lKGqXvjAv72+7TNGDRmh3odS8xyVmE9QDLI2NqdSQRWMbtUaSSQ2J2N0z/cu1iOtlVd7GBzrv8+7
uDIGstTe1vjKAzo6OtEH66cwEtm7qOZjJX94G+lV9hnzO6yoNF7NSvOJfCdkvpfFrf72Cw5hSsNj
KScfbL4DwmcFdNLUNMinT+/JFJIH7VnzmVEancU+Xjl98v+aiCDBTGwcfOziTKE7w9ui5CcX83tO
7SqCCCvF+ls8b5vzgflpDePf71+FxjDzg03a9NlKyamoFyRwuaMqGDYJGiiF1UcyF9pu85tI51Vl
sLQqtse+PTdT3j979ETiOSHdJbAEvol1PowfJIUJYtTE8W2k1q6aJyJQ81ipqmWGY6/WQ9Ni+gb1
ET2iBNUyWL7m8+WOOrkxyqdsjRMtSXixjxsr6IASrqBTt6qlSx6yNNwDqn8t21EkXrrCjXJgjv+J
Ffn9EB7Xmcm7RpZwi/DIz4RiXTTfUCARrcpQXtkOI/sQFQn5KRLgZ9EGk2lrn6EJ83E45fx5vYEn
1HhJmToLjSGScQLGrtFYDDDWx84yGImnd10WXsoboBTNYdIRLtmyS8TH8+PPRBcW9y0SqXjyva/g
1+rSuJyDSXm1Dp8fgb0P1h9nz44B8wMkZqHM9raNklI1E3BX0VyzLo7zy/OhNBIi+rzuxMs6iP3O
MRHWAESH7FyFhu3qrK0KVgTwZK1+cy1YRjc4yPmSDsGuoDjjSKAdYkSjQVHEhLl6A2mrcmyU/U7U
xfzwH68TE8x1o8u6XATKFnJQ4sbo9pdT08tIXl41jJeNP+ChKZc3WN6oYdnCaBj9di4cskMO4H0W
aMfZh6QkJveFOeMY8fOW55Y26iGPXJbSIBrGPd0ct0FM6NihaANHk3zbZD9zc5MH2uQJHw1Xy7sy
SYUlgKSeoUZeDQKMPymF1LMLd/hSqJaiXt86SfGHhHZnzgTzDBLBMcb6lT7NxqznBue9ymktH2cq
qU5EOgzrKK3bsGMJj6ViLcYgrUIp89a/3srGA53N/aN+9LS2qn61pO4aHCh9Yqm3AJvEY2UJVJ3y
5bZ+qEPKxBNE5lWaZ3M08mV6FnMZysIP5HKN6U6IBIBw8QvM8Yr59wjGReD8SdKA3+YFXcdjhQZ1
ctBHe1wQqRRivuq5JI3EKJyj0E8NnHPDqt98FSVPKqWCS/V+qLsYydEv1Peo9UJ4ewk6/Oku+FXh
WD+tVnFLqY1WMt1aPTQ2VSVodBAH0oT67qxJM6zDaeHLH6zpQsOWayVrE0ZMhTHuOI8iqdBXTW/E
TncckmmNHOAlZ2AHYHc2+LnMVHhW16HwMVWe5Gpp+kje0D898foBGw0UDcjTA30FetfU4bCyctzO
rj5cOMJqbEzCGsY3OQwFRJEUlOF+2/beDdaqfDHTUvxdJBdl7K12rTYdZpa8yhZtVh/TG+Fy0728
LNq3LPG0rZXyaP87qQdcXZ6To1U5z9bHceKR6zFgE3ii5ZcfPUEdJ+T75q9btfqlAkjZsKHlE6QH
Bnb5LrRXtFMJE9+ytZRyvcZnfmcDzWUHMENd6xceSO7f+080ok2nd+1r/UFYfO1VjZEyZtqxzfFs
ykelO9sgr1BOCedN4IXPreZ62tlrSdY0dp0SLflbDgysvQnPGCJBaY9ZoBokTzL7l1vaaMxzj1rg
8inTEGhnUY95gC4/VSOBqmQKmCx/LU6BGMfAXp7sFr31YfWECCC1hRUatZOpaCsPdiigUm8Hh6II
5Bm+dK4CdHfCsqsO6UmHg1pRSmyQgjJQo63pbOroDbX/bamG6K0FOssX5HUESHwV9M1+99ZMrbuh
uj16b58+vAc3vJIO2tra827Oa+/y8jzSp2nCne4/4Qk7l44oHZ0KSBUNx83q5LV1+j0SUQV3CjLi
Q+yALFOKk/wFvLdnV6sghnqRFD5BPWNGiAlVtTNmM6Dg7L+v8jZHOeeuhP5KmJPPhHVQrZwqnHKX
BC4XOYpbFXkj9cpvanprg3SBgUSA1J2m4m/3lYjDXgnkhJgSMAeRNb4Ckiim0mS28RfFtFZNKjKd
V83wRg9/yiVo0K4Zgt2qXOK6aZYKfUmvZoDmiV+rIcLrAVXM6o3zeKGMqq2oHZix0SB+e/xCDm5j
5psgT89ZQbo4l0omvMK6qVVAAlQoVdEjkcvK8XxJqLwVVFcKpq/s+tuVE9Z932zMrs5Eaa4cWVCz
9fJb3LwA2wMdxPF35Jjx4JhS9b6c59XvPh2gXUpz4m/HkxvC/NWf/TjVJdk81eCOUwkbhTRx0S8B
jNEvQgpq/jE1hkjb0aoOAQwdBblMbTH/83FUP2/SCHSjElGC9aa+9XlCoqGXxU+1I4cf+wLBDoj7
xlonfNplq+V1+Q31zM0zKE7BXBysenCfKm09otGNqHI0TFwFg2pPY4mP/RIka9vudSxyruT2Vka8
0A6xgfa+kaHy8l1ybt4MrS9J89sZ+3BGT933WPNdr/UuxchP8bFFOAozDIR5SsF1BPfD0gHHEHhC
EQvSnsjywscYQM3/WnjNs1tsVIxSOBw0V4uH797Od98n0b3WRZ7Xj8KUJizeBuMgiWB2Pq7aLAAT
oNv/EutxmNYhV2K2tcfuemKwddC6hd56gaJDp3n//IDlLsV3w+zf1RC1jhZJkRjoQ9zmDtVCqW6T
FCSJky3PvPiPzlFGG5u35q498IzZFy8hZH+XWD3zKIlyIJWRUUggmAzLtd9DZxxG39HF3mhut4jr
mKdCjoIFdJvJwK/L3yJWUZmtHEMrW/N+wLjFYYMKpx5QNuFsPpmD9V8A75f1KxmHelmPoBBwXINz
ewUClDPFQhyp77b0PhnKPeDW4x0QH7zu7ZTyJ0gGDtBzQCrPHnTnE3Tb7+D1VBsrUuaSjBbq/dUO
o7rRIGnfRYk/6xIgyT0orNxdgnE/LtbqAz7m7bEWynSG9FiarXN8zIlhqJ08YDR0kdzYBIK1YEd9
KLkyrfK3mNZm2yTMh3Lsv8JWXt/eUbji6maqDYIgQfKtscAvOcndT8+e4MpQp0TjKbSnae9h6ug8
o93QZ/5yAIpnP/eNHIbPHK/ZRC7Cz+gSr6/tVvO0tAk6IlYf3cTAgq1q92pdSjYr4vMer5puf5tX
wdnSSP6G1b3ToeuUPZPHREnbvUQ1bGQUSSI4R9l5IXqyd85S/HcHhcVT/MchDUAIxKVE4c6GBFPW
44pgzLbJ29ztRGeCJzHrRmPzV33FACOylSz31JxRO9jDBC9aSsiVHdSZWsJeV/uz7rhRsSvkL8CY
HICHyY00xjeswdJjzsUyo3U8BBLVWOpmNZVwtF6r4e0RdSmGYq3t1n5Wp+UOJaHfZat7a1bQISFr
IfAZVGeyTIDvk2xYdO1OUa9WaSvlW+Fzya5I8lCehff0G8He4uO+HKHlF8o408ZaqIDSMRxrF2RR
Iy80nYDl8SVrebu8yXVxpReSI2zuhkZ7Aq7MtP8KcEI5sbynL57tqiE+Vyfvc6bTK8EkGYne1ajn
vYDs5t/dGr2g0GTt/2qsywkNkUL4pVg4zkNzVPg5PSYZMNdB98vSbj4kl3XUaHfXcpmOoudDoyPv
JmIpwTKGuJg/QkthnggM6jNsCfsvH7v3vdu/oum6bKMYDjuWCUkEi5LvVPfOPoGeHIADS6Tac1zr
l9Sw2RLzogOQcsuFOp0PsGZnvXnRPTSPBJUmxlRkeYvU0w6L+YGo3Cf5p+3R1VbGLrvaZbwvK+o5
7lnRAS3+Y2b6TbFC4InVbr80XVg5iLr8vtT/VRFCheCk1Cssw9aH9Ga6IRu4aBNFJ3sm+GY/X6Bz
hNfVZh4GEIN2/p8w1O4hqvsG36Pg0Vmla4CylC8FmLHpONLpgXMSvZbSO7RnKvG17UmPuYwcqMCz
1z8IP3XP0gydNTO81+4N1wK0EpiVkT+xKl+SbNjlUQuz8EhFk8TFJNR8tlhc+4XBa2LPRO4fV2wG
VFd/5GPCR5Dt0oWxN2XAkSJzuVihTXCoUm5pCLEc6SOMT0s3yb8gz9Q+5lsfoTCGcYdnx67vMkBn
T3PEx4/Ha/A+ie9UQS0NKzIYlZd2jkZSWVOMnODn+0v23DDeQn+bTDqi7G9a7Mp341IRI+cX+Fog
TSkcMcxAD+GwSAFV1/9NAfVRrODRw0hZlwuLA8Q/cxnkXfYp7ZvRCWeBYLc2RyOE+/bUzJxrlvpX
GGNURb4zvk7Vgc1mYHwbyajm9ztg+wJIZz7x4ivu9vR1GQizwrABM1hCobLJdeaDCNn6cRJTR9dw
uBhPNZjeEioBsevbqjGZ1po/UyPk+5xsEBTOEHNI620X7YFWWaEgmqOt73FSffBde8j5Q95GfGpr
bYRQdd+eH/H6NsYUsgwPyPxZ6Dxr9JvVoS3C+ReJRWvkLjWItPRT1fxc7mdV0ZooATvnqNM72ffH
kUR8pg2rkwgOQkdgEV31mpSlhaPc1c1oityGHxf9xa6lr/T3TAALhVL8s8wnKNj/+qx1WYYH4Be9
qrWdyFIMn1VFSTFdREkb3HXEF1kWSslILCji57Q/WFXp9KH0WBsazVkODzkYflSeox9xUtk1gyPE
CIifs/HEBZS+OlitDThhLDvmP3qh8/+Aq6cClJYUhHSZ1hPYH5oL45t75TWFG/Z697jrp6FT47cc
Nt3ONWHAiYYW7YTq/QFjE3b8uke4Wxv23rieN1uPgxnGWe52JRL9xRcGEVYbFFmibZg4J/iqJRpl
+Il/Sj0iTVFQP5NOAwu8Oy3Ohkh3IC0u+cdVRbO2Dm+dhn5MG+80KUb2xgy72upDr4OfDHe1oLA6
BqYC6/MM4Bb5Y0Ju3gX8TkcLRoKtEYMXV745N64d1sYLB3rIKB84FgQAJwb5yKouRNRjm9dzaVZw
Akahhy6p6LtYjAEkJV4RO/mC8kSqqEL/scn3plaZxSNVtXW1Lt83l+nXSzOvppYgG2siOCW2B1Pv
vBagIuWtMgwO1SMN2mHieJD5YV39WducgcChI83T9W3M7Qv3nHYMcBZtwVlYi/UTJs6cgWneNq4X
NzKldKb28nX7GW9u9TCGczNfm60sqco+EDxcRqCXlgGrwz13KBDmKLWvTKfEAK78lvQlJWAPJ+af
f8+jcCME/vTkCXCsW5/JSLglMPjHDILMT7R/STE3fTy+oaEvrXziLVLuFNPtFTs8jwMo6cmFpJUL
+vaqLixZ/W1VLVMLgFURiICrjMxOLvWvDp1f5Sk7ACw7Ep0cyDNRtOVVyvcCj3PKOKfqCKlxeGWW
4hXuGArnaDDXdaJckKu1QzJcyKQF97CjiLKBUPWj5pYpkHfQ2JbBYzVtBpB/3kDi75S9BG059zpw
D/tItz/ENNgfCcVNI2ODOq+cfGAWWhh/5kniRUHLHHBPj6wcjZsibztYY373DMKDAjcsckoEUb/M
kiOo/m/m3AO5XYyfdzP8I6ZRYert8OTwmqKzKohnMivXdisfgpYCsEUFDSDTGxFrFwyJuuDjTvCG
vakEIp5c342gXtcJXOdeRY457H5qtrkfZFXDb4NEmQzF9IDZurmSQS7dtZsPdfnhprTBRw/RN2Ux
jKbJhTVyAAh9Rdvhu+mwnnRxXQi1HEoud3SVISOQTWIJOwEYtNEmvLZFC6pI8mNHSW4OwwYpxbDC
+uGlaoaN8ray3CtOJyqKsS02IZpk34VwHUC7xYa661eQVNkvJPTvxchOfFSLrQ2YhnpPB0j9+47i
TzYjpT4UEVgCcCmLIXJL1jtQofRkfmUcxG08CUlN8FYbOkwlnd+dwPtNqK5o2WgkrZl8F4Gc+Rv7
rTSu0EZihQc18Q1R+W3M2vbbhYs3Kiz1JIzCBZpU8nS+9lxKKnB3gxdJ8MEHAoDpFC4UyTerad9q
BbWxhp1BAO346QJwN9TXtpe4mKr06yb+0BN6bW7oOsMCxIZoj+Mu3WNjkOqDBCt8My3oidplXd5K
3dVWfPbOH8s1y5HVCwY2JTAeh1hK5Zvc3QDuqwSHfUGuIkJBef8f08MwaENa+mf4kQuX3RgHhFmV
nqJsgDR+jY0lqGVcd4RqNzlmijy5hDilMZd+DP8rpmo39cRJ32rXKxS/IAhsyBQxyNzJOB4sdCSm
HAPWAhVWMhZR8kZLnUHma6DQdV2sAJZjheFgEmNi1TTFF2jZYp5JKyqd1+ddAo9jcquKjZ6eFVY9
GlTihQQqV+BHyjOB3RTffJchILLkDti2eKUsDcLRBy9lkU/m3MQ9DUSqOUPupE0FNQivS/OwTR4s
z0SUBHyc+BMcZcud00ZGEqX6JyoyeRyznj9jXOrIt/MConB3u4xVJxyNaA8IsCSP0RXQ0GYZmrIJ
Jz4eGJK1g57YUI8WRG9936Gk1pfSN57ywh9pvIaEwBVRujLRfXofKoy9XvSaV5BaTPNvYGFlNZai
U2XnlaRjb5ULWpZcVkiNWzDRo/+o/AMVzp8ruUtw116yO5bKe94QQnFOvrS0hNCeu489o95vwcqX
itpKdlu0kGxMyDjAEsdKhkkBEwJqh3AoCYHCCocNa5e9/PwhnJ+HTYCT7R3Omxi4jc7Ck6eQTsXm
oQZobvEuPD50t+xwnU/OyXc+esSPSHZHZW9ouQJJ3Q5gMqfGSUrQejn8qdJVwzb93K4BykVQbcCz
88EnvklaVQoUqqw51eb0IxYT5GYgzrnWqQXRKAXciIbaAKcrwqJo2Oi3QF4qp9BmdCeg2EAjOFH1
fuy3W/D+4Y3nxXJS280eVv0cPChK5A8NQ/Lbx5w09NqsodKh46Xux4zbxYRgT223VJWVOkmMaqgd
TJAvaCSFxT5h3H8ySmj5JBPF58j/yNOMdvgirEnogOQHdq9+KmjIVkVSXR6qj+ekoNzQ9/TaXlyJ
M6uUXudfxualpzGAEqCViv6GBS0CkvqG8ZU7g1wB1yG7v2RBoxJSlZj66trna30s1Vqxcm9qRGal
vy6ycJ9j7VWT2uTf4l8EoadrQz3zJaUs2MWc2TWIAKJK7IoOZycqVduCh1x0rDH/UdV9MxnbaAmY
4OY8u0z4QBmWybAiGGFV09806gZ2+7CwBZlcgAJTfBgs/u6mKf6ZpO3IXzwVfI8ZeIfwA4Hc8sBy
GgzpdzY4QJ4Lrfq0bckb1YC9M4+90RaPuzacXWF36T7ODNP2bKwAp8Z/GBxTGJvjhcNhJqgrQUwR
kyS0u6ecG8+HSJ55tU7QE1+RAb4Zxil7gHwbRUbvHZmabryp2FaPheiQ4oTpb16lrSqcsTavqE3v
4AWRS6AnytPvarN4EwXlX0GKn1I0CIAk8LNSH27mIP8hPhlomEfvIzV5VUROV1x4jkohRXU0a7dp
9CF7scdacTq1xm+kFrLE87x1o4J3xHoio9JuBHXCFs+Ye/eiMCSVjltq+w2BmC9U8bKjOQgc4iTp
xo7X9wwJeNRWBlIF6NjBy/mb9jzurdW97Lrmf5uRZbGMjvsIl6kw+GnZlIUKPqeW7A5ADrTYKCd2
ZCoAElMiMEX96XXC8qZQWwn80RZL0CrAoF1J9F1XNhMBmgkwpviJ2+1y3U2Vmm/Z3Z9LJKxPLWWK
p/fDrq/Yohb6GrfzP3CZ6kdCvn9NuAWr+Bm3ioECb52GZaE5Zrop73xj/OBTgUhAq/HabC0z1d/z
p2H1dpx8eqsDA6Vaca2JYK17QZULRsc/0lBRJhvIGA1Fi/XcRvF5trFm30gajeoc4/xCIT2pIqBB
XRbYVcJAFZxrBBQMeCGWW0p1auaJqB1D1gDd5k6ImIO37gH6e9ASxg+mhtY7XpZxeXfhp4VpV4oC
gIbxO+OAeoOyeSWm4afmI9iKVXLWUynZexvKJXiZ+sv7YG6AYqCxc82HEWijqWX2JsPQ+wqvsVUT
NXCNkwy0/PRGN5oUJ1iryKsgLyFHBr2V0NC6vWNbULLUhjgpepwB4hJGJdYuZ5OrNJvio91e4A6t
uU/c4W4LYVbWAZapQyP1Ewnx7hjUhJBcOQ/TXWET98qaOCl/37VIOLtoM0BO+4vmoPbkO/qI/8qA
HIba+WIpcdrYOFMVJ6XHukfcPxDukilbmpoxe7MpFyMXZ5BqxLyzeDw6p3AxT16Oo0l7G9GEg16l
5P8cnkG0NgTLNBc18alHvMT6bOavAkTo5Pi7SLMvCVlUUgFkKaBQME6EMy0ZROG6YD8gAvP2fIxk
B4w9E6R9SSxjwX2pOMeq1/UDM5dW6uH001O0p3PG2EcBNmNRnA+UBU+k+PEOfOxsiUc0xUP1q6ZB
z0j19uIxyfdaZDtfSnOZY/TwLNZsaz8kRueOt0MHcPNhiv5jBcfKwFhYW26tUjgKTAsjGwwIE2EP
A8aftSbP0J/OzRxqMkP+Z+cXvqmxrEfCWP5RD6AGizpLkMxOsjs/gIzg2r9Lu6gqYWPu1C2EXnza
R6WVOE0PG+EuX6EqkYQIOD98zWlCgZBrpO+Bwd4D28hJNAvCX2PnBQlVWsrCFgMhZXxA3xWVBDiC
5+fGqx/k91QnY6B0guroXcUIpXZtUY2svhNzDyuHDSWFvrX3sc75sEaC2QI5BOP8xYTajQy+r1DD
/kuTiL46qqUXfZb2NryQG09R0GayYQshbtPc9+un5btsg8T6HVp1JNpZtSGTz9up2MPUqvES2aq/
+fdkBFE0MvoUprfiVQ2V5G/TDztk1y80FZ9pD7i5lovx3WnI7HjJ/PIkYvnBcIksbCNZa04qdrQj
7+m7rc2lAGxWnsXUm5VqRWi9+ek5HqfsY6+LTGQTlRE06RhjjWPSOv2oN5EQXKLH9Coh477heVDe
9YBiq7/gBz5m4/XNi2Y2VCvI0HsGHyCw7QnCsHK6Xwkrwd2AHSb9LkIcIKPGT4caE5zuVr39ItUx
5/JWwFrSrawVGY40iOPEmIG+its+pRG9ZC/OGgOeK+wndF278f41te4E0ghBoI93JBfSnLzPew1x
O9bnMNoZVy9EPHceo4CaIRr2kR8updIW5g7JdK5aPL7of1IP9krPqDBVjSxz3RyhHwXIKf0Xwkun
jJUtwUoAmYZg98g8qN0wp79dYeKiaPVWHGO+kv7jkds6SPFCqsQQFVoPI4xiJ6Ba7llbckDsaeeu
O6sE+xMcsPYE7pjtD+QSef2M4HkDcIB+miYSKAxlPirKNbV+ZKp86JxnfsD0OicFC7tmL8dkmAKA
hsSpXGjTHfBIj/o69V40XCJUKNAW2Ko8UxAiSx/NbRyQUONPtQf5AbWUO5Lg80kVzb4em1gMQFyy
b6AgmJ3KZuGMYSr1gmXFhYabyXjPQl8Gt1oESPz+z9Mv83HWIGSZ7JtyCZNirXory1I1HqO5VbZc
wHae1h+2PSpH2dzRAlI6gYtWMPkH5RHIBP1Ov2mMYIDWMP6itE6c6lidraLsuallgSgE2jEceDYq
F8pPZZxhlIzr6WlGm6688tw+FbSYE2NTj0ur3QzuQUlV8El+xOm58U1UmSBr9jp0Vn9CjR/vCyPd
X0g3UmU0fIORIQEjVokdbX1pY6ll0ngeSi935XX0XVQC7L/qUiqYBW5nZPkxfvFceN6lNTA12Rsn
Rk1ufJtSXAPnYhQhf0Jh2p1tyEI7HdncPBTU+FsZWX3EYTu4eAqG4Q0aCz0L3m3DTgMyAIYdPC3b
ev9yZADDjDyoe+rDJV4q7YNid8hY9w/+M7u7nUUpc4/cneOrA006cyYe5LQXaLXJiGknXw0NXKar
fYr36gN20NvAsbehKXPNh6l4dn7gc/PIvuBNgEz7IMg7HqYJus636d2iHtfJjbW9ZbhD9Kk0o4W6
UfvCgxl6bQE3Y80NU+f2YeL5PWzlH6aqCSsuM65CP6rGg5hI3S/uOEi/Z+YCCVOXmFbivWoaGGeY
Po65pYQoIeWov3uf13TAqjtkolo4uq56LQ==
`pragma protect end_protected
