// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
srbdG8R7jOgFodYT62pe22+B09nMiZjebkU+PmyOZCG+pdoPTUVIOCkxXG1WPp1/xTdBW2jfvHn+
Q6zITZhbMwfpOE6e92TyoQLZdEAiELyBQERRcepUi5uHQXGPUGXoJFt4hOuP9hTwN84iDy4EdYvW
IR+Mga7UljCh2YdWS3XdjKfJhSODfTNwAhXJpBz5eUPBno3oUHIMd51X+NbITyJil1OenP1vDCiq
ECAaVyvLoQB2PlFAn7BzfAu7TyvizlZ6z55eqlS+ILu7X/NawxobgLwaA3XOPpvUEQeaL9FxXmg4
jb9SXObgwjqT2L1VYEiZX/qS9+q9a2qzxmWDlA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 44848)
0iaZ4B07XbMx3I3oyk51sMOfz881OCE0giSas1WAiAwjr9vEIXUnLZoh3B7aCAcFlc8l150GxHvZ
Y6yKYODlUYg6auBdZ+X1joI31TjnAz/Lfo5FnEMlujC9oGPEO3extBfe/BEq1JF34w67KkpXH9XM
0GE9m7IJywtGWMXym3aAZnPP0nZ0T6gXgNYdVomflreQex7MuD3/4qXUN08WKZlkD5MRp9ed4J0c
pNsHB2289RqpUcurvQQ4NHyQ+Es7FvxfaHkG72qmWlFVWySYqems5phI04I+ivZSMZW7d+o5LuE8
1l5areJ83aMFgwF8VLdou82q3v4SHPha9g+WLjgi68LISjqryUSCwoO52qWvjZ/U+27HzARLdI8I
HqqaTviX/raqYULndf44/YYbA3pYqP57a223X76kgxRfh45XT4IiZPNG+N9MkZfqdNBZC2+1JUyz
UTAr9nRgpMtMNxDpRv8XrsNf3HBeUL9zT3gVgoK/sOnjKZkCt+j7p4Rp8oYa98QTLASe89mU2lf7
Y68yAe+b1SZRv9b+2IckpmLZUOCLIUavVCEGrF/5FnSX/FkWa58qc4DGOX2vnmvSBNs5EtzA091+
u8hXiU0zFqUBndjFEesjJSx6Ru5q6ja5Qgfv+UValO5eF3pot2pT5U2mL/Z/e9BMO3WaaEbBM+OU
wFkyg9oDF5HGIpYodwo1s/6g8ApnQlH05jGW+Oz30mXPFN0cEfyDIrOcQ++Y6IWedvYFldyW8rIw
ksQNpcn8OuuLaQ3ycdgvRNblU8+aQViNvgYyzHLJmAsGZqEw4t6xQQWzue1/8dhgvbRXh2lbNQw6
7DPIA5I1YqQluqSGBnWJxuRfV1g1XNmm332nzMKTmMUbA+2p2COE4YcpC0NqAK2ci+Caq+oFE4OK
OCjFIpltPuMvSzmsi9jqV23Ej8KE8cwT0K7IqLkTkHqxi1hMulI4KoNy8VaiiFjPdfSITsbtWu10
HVSBb2G/uQ3j0ONt+PQobOyyBuyDfs0rBzPkS+eqoFEkcNb8W/yhWM4Dmq09xT7Oe5AOPl1lntn2
z8iFmHRMbG2OLGLCbIrmK8hw8uOdeXsdCb8XSGcRJyMA5EjTnYj6lyyyQ9eIw9az1nxevD0K27Ob
v7PdLPLejbDaSA/3ldhu6avsfI7n/VNHENhXDVPiBG7MTrbG3rmKtBpR7M9IxquHIqh49ArASYXC
ZkcdS4PVbBMNby2ynJELt5pbZF8ZObs01MsnC/vNTJCY4+zeDHBSTmakLYsOm9g/tQjok+1Ljjjr
VxzxyFEKu8hfuEBHJnpyy4oG3VhbwQ01zgdVdVvX7VqkBOrZC4l+6ZPS8WLKoW6R8MaRav38hIsa
O50VEEfhWbMhVruH7UF+rSTp+8DGFlyyC2oAWgSAzEPQjLVGbDRQNiQe1xobAqVzcBdOUndXiIVc
0WW53dbO4f+rgRPmmt3Rc8XhWN3+izjYKTDwrWRwONDBV5dJguIz90XNqsEUkUv9W7KJ3cbvkZT+
5INoRVsglv2evZdlHuDSfYyG1n7MSlxM4NU4yZS2TAgATAdA8FvOcxX0c+FKm8ODfZKi3pl/CP+d
RiW+4zX8SpCWXFSzVaV3hArmoPDKYBJSXStFgm0Yz9r4dzUZro7HbTdmCsDy1hVHWrye9MD413Im
/3QDZcqzUld/uqOGPblW2mEB1TihUADlM4oZeSoftDOf9lDm7HsNuUJD+elUHIoVfLevIV7o89Va
FqgmUV2QXqIuZNVyZsUE7kIieOaudPf583NLQv47LLGcbBEK14ToKJrKN5BfuH+tbArsDQiH6qAZ
DtwgnL4Zz8jD6nR7w5GofZikL6vz7j9OH4K9fj1pSTxJA7Kp566Cxx5PwaI8JFGiRujm/7ktjDVU
dFN5m5yOU9oZ9JG/pu1gSZWG3ViixRa8MG4KF3SLhQdZ+UEW1eDbJriJBY05BEkVZQudx+VFn6bi
7RJiirbp+Wy9W6we/gQuMf2eSpiSmn+lBpL/GhYzxhmw6Jv6Xiin5wJYkXY4QucwvRexbUBO83gd
QV1MpFzSzvp3XHPfQ3G72RtACgSGT2qhhHAb2y2eiRafSYHrnLecoQzoqY6gfJRGoinWdZcKI4aP
k3n+8R+AJTokVVKGLObAq9MDkddQ0UN6b8PFD7fz0L3jePcCCJ4lgP1H7CDN61LvhGLZVQC5GWZn
6E0h3jgvcHJ/h3JiQNQXXZnO45U/yu9hDux/W0tZxSrTmps/Zyp/x+20f+qXad2gRwIVQFagI/IO
uMOhePYsgAF1RATS2iWNlZ2xhPLG0PP+QS3IiF0ofkCIn4xUAhhQsJ1yXh3qNxXx9U0QJRJG0Q7l
oAI2dG8HhpakO0kFuBkcdHBJ08hSVqfIJaxRLwtP3XXlXUK48O2Tx+FkY4EcVk70k4E0Nqk0WKse
HrxYDYsA71syPXJyl3X9vsxpGkAVda1jvGTCcsPjFyFiEDpCPtuAoTv29phtrgKKqZszv0ZprGKQ
Py3Juljb3242of1MzJFaPYF8snJyiaJC2S0FqRwZEN/e9w/mITMwB8IK640JB73PRsIj5b0QwPAA
QR4ryY46PBunCYWU2uCkDmE140xg5olllH2jri85hvvp8VYV+O69ebayZPDDVQdTPr+GEchddv1k
9VDFKftSWpTKFhbT/tj0UhUsQoMPrjxE5Je4w7Awdcs6/UMyhmfOL9Qj/HHNT0IATOCokI2eu32w
kl3T68AsgrRY4fLQjfgK0evMFT+oK8otUYsfS2MUv3SCDGPvSTl+t7u/WK8QIbVHWskECv6AV0iU
RvO6ii7ils+M0sugnu3O9y0vunm3qd5WdGKxz31rrQXFdt0RlSIRurqhplTL5e5N0jfLyLon/svL
wZx4ZXyvk/16adgeqwdoTKnXwzErv62MHUZ2ubPB+1VOfTa8jZVNY+Udte5laMkOwa3wHkf23hWS
tPgG4yEXj6JL82bhtuiBGWSVa/DjE2SniAlKvu8qa/eg+CvQ6HC3+4E2eHEsZRVGLMjXZccn9V0V
jZKm/tUqxdV8hNz66UAHwtGDvcRucxQAcj4gGuCNJWARWh7aMo2qK33xXzw38m1CpEF8O6A69zEk
dZ0TWtX++d5W2xZUMDvYsrZRUB2CIMFweX3EJgvGtVDVji8hAHSw2zSx5XNwm/w6VfLoJnIcRm2R
ohiHfQVjWRaz5qjIV2MWfT5JTNQwsTV87SxX8rFpvLzSkLTnlIlMSNbZQzoCIrKJC1X7huC0DFMu
S5nVV2GmAp4qjgKLTb+4O6raPmmHME7qmI7cryyps96G6+WanGJuOz61M0Y6ZC8JAf9n811vZeLu
M/qe4iAKTrlFPNgTq49JYUiZCuAUgIdhSkkqc2O7ZPiXS1rvReG+OxZoXAPlU+zWkAET3UCXzewO
mJfIeO00DjsgiDNGO1cnHsXVj1zTB5HY9Fba6aDBytZWVPUfDrdlY7XECw8hWTQz7sjcP9baiIIk
F1Oa4w7WOKVnpOPyC/Sqm78D2ZctvVQPzqaxzs+YujJRoP4qiqy8eBRah4iCCNlsfjVfawaB3EkT
/vZLIpPuMyc3S/7gpAfgLlE+JJsZUQfKxUlExp8zQFDwKZKo+IpVl2ufwZ1cIt6e9028O31fO1uU
QLzpuxBtfDT63Qrx/yPpt7GyNZ4ttpWqcRobC8GTkxoIW77rpBfzPBume440S9ms2xmTwd96kSgc
l72o/6qgoyGhOEnYuklDSO0ndw/NbKN8QoAh+OuRDAMAVghPXHexgFmZaNn7+5XObLoAD/BiDLfe
O56/K/qeXhDJOt7OWQi5sdKnyAD/iXUtlZm8aPV5IItlshcipG9gvt56F/sppGoeMdSEybJjv5Es
FVfPykvnx1ZwozaZEW+cTCzp7B3eWsX0uzTaOHMlbPJb62IZpJQeTDKXTbN57SiVFpiZvjTO+SFr
K3uECUl4vHSHHQHYOtF4hNN4Vsm61ehxq2+KxN7DjR1Ao/a1MczOrDdtzfK1gUgSkNLZllNVfqb5
guyTgbgkAMaN61S3o2FZ6ViLFdw4x5A+6pXpZwoAPvE8ZnXf9qGAy4Xw8DSXbpZ9XNYgrI/fLI2P
nDUT5/fSpi+Yd1TwsI11d4GJBOFwVqSS0kxr5bnU41J0vzwNpdtIbq6Zr/ykhaNJY2a/02PPz7jd
gSM76O8cO/5DQXfi3VCYGaz1IKsr04zi3oA2bB0lKuVjnX12KMaNPBm+d3KGZYmq8Y/sWQHk0Jsi
XvcQ6Ocuh74dkc7LbL20VtTSXoGXZum1kRuvjdwFOS62X7ZrzYP9xbBdxq2jADSFsV2Tgs6NyRVN
4tCvtPN16LcMZjGFIJZ24wxtbWPXvB8epEC8h4xVO1FJvysLc84leWgs8tmDaMwwAw215Q54Tqom
cCcy1hW5621E02B6yvxsIUzts9dyA1g1xhLIhSJnfr4zMiO+oPEpA13N/prMwiHdqhg8uXj288DP
AGcpXQ7eH/GmoqxCgRuhxtRdEeCvEO1YEB82Yw+H07paErpyzCIWxHFqhiku5x4K9ZiIrGVSAm+Y
0UuHoXmTh7rTwAqoXcUUuF6w5G64l8ZMSyOVmH6t0iO1NQmH7+8GQ2NH+EZYLDf/Jf792q7Y6Tvd
PiWZAGBxyDiwPVVEdl5UZBUB/nUEO5fvEAd/NkrHjgODDk3LTuEaBKuX5kw+SCsv1rSQtmq7LIqK
nB35atG39JrSKFDkT48sjpid/8vE4fgw48OAnTMLpWpptiMcio6+B11NjbXcfHFQkCLpV46mdmaR
iPkfO+kh7SmE8K/JC9yHF5ZzL5GUx7c2HdgE3Zeso6iIHxc2i+TNJN3SKldhYYhvJ94MYwSIgShj
WRThCNE5z1V0P7MvocMy2Ij3l/AJJ40mfMfQGyv0QmMUvnIpvaFpn/gjXuF3sxDQOehqg68Mlmib
Jj9PBN1R5seTwzFqkzcpTqrxAIMVXA4k3BN3gy70KqmwRyPI/rC0lr1YDwOQDqo2AE+WNnEdPYdI
GF9bHAR/16sNYG2vPvF2ZlgC1L83vqbd2OioYdsmUOUyaFcrALK8XFzzcBKwN7g+20SZ7guYS1jd
AIiAnJEQS3clT49T8hMeLkdl6sseligD0Pv0eA96vWvyTRDUqy+j5KzUKY17YQz4r0JYthlRN2VV
WCqnmM1akRwR9r0g4O12/x+gozKVcfMncI4D0QEmMFZCVUIH/0KhNmqYO5mtQaXY8Ar4kp/sNwFu
+ITesIMWBKZF8XDytKVSeTa0OhVppGkUZT3gURlzeP337VQVp/06coTUs5avWBKjsCJSo22CU9Pa
hXDldtTacmMfzF1pUXTIOnXtFBfpONRanflDcEzW3QRQ3RXdYAnZ8kNoB6Ppz3bNAFf3qSyRddgj
MaNamApgkoXKPWvQir6ry72EjpN3So9jpB+LbZP2NXQYUL0+zi2WPW0vhYBMy4qEEJc0IvqelQ2G
ZITtKxNXFm46jYmJOto3veXihgSLk5PmoXdz7n9cMOxlyZUIYjB7PcXtDPtjNyHXGp9uRIW2MYeE
VcL0WazDoaze1AtuCIspX3FLarbtYl+4aWz/0IYNgRYytao050EQeMBUvG55xVYwosB9dls2LxSQ
nfCqu1o60MHlZXmjZNQYJjwCRwghgB+aXK/vrtsxqXKUBSFo/kqKw1d5502N1uniwJZhs9ITy809
A7lCW+gVcYqAiTBXP6dig7tjGcJGOnZPUtn7LcjxQbZ8lAoyUXL/YdazoiB/fF1xpHZXuOfwoQ0i
nm0LWXHdLpmAf4+S1qf61/T0putJlMub1e27RVZuoJr4O8Xuy9yHtJP27N1sADYObWIKIGcmxbm3
DBoQc4NHbtNdrBsbAPP36+6g8jhZVEVzN3N1d63SVrJ3SCcaHdMYm1v6+qekZJmUaCxFdcSOdCZY
AAJPLExdK/3Ra/+KHYwvIW91YHqbgSjMJgATbxcKvaPJGAaYAFM35d5qFizAzbZ89vJekPs/A6n6
i9LecJ4bgGzrecFQ1f6H9WYAR01AdJ/onMvdct4/+31Rp2XrdIZvcmBaQRwdD0MUwl5n1WFQhqrH
bQlsdxuncOhc4SIilksSaAIO1CYTRKCI9ynTxE3qUSfU+D7Qq5mUGLTMUx5grlJ6o1mSUZJTSFW1
Qm7k2zetydmFMXS2H6jbRE0mDHEMjvWDI+azSj13nzoAKHaw41XcjgKwZy1UhGS6nJH+O0mMrg2X
yJn6DOoTE71JlSy4hklhJHa/1kWpLmE7/l2NzKQ0F1fobnsJx6OA0J3/3cHY0mRohFFCfsoceIvR
2AaHqXZEztzvPYWK6EjgXUQ9kg6JtohCVcbajKwyMGnUq8++zasYzhK1Pt6sLfUYkP/54Bqke6cI
tHKIRm89czgddINkUNEFuxIvTbs7loccGr+Im98LuZKMGn4ilKXeQouaumbTRFQsM53ZQQJVRRTs
pBUm29TeaTMDTr7YbmYDDKuleaaHEl9ujbNtmZdFNxq5AW1AG6yUJlALC2Fjc8cawle8JZydvKMz
7bNZdSo3CI0deFunhBQi8MBwNEs8wmymxnuH3DoYz0i5nvCmB//ufqDajeQEsn7YH0Z1X2YAaDh6
1ehc8TYmA4gznx4E8s4TMzUzSHCEnhcd5b/5RWup1fsAoHY5pwp9MfPXthaCQbG+1bm8kHDWQiaH
U8TwjJwHUO/UJlIwfWOzS+w67HfBpolh74WvCMPUTKsptllcQThUa3wsePveBz2KOrBoc4WtJp1r
jxeoXc/bUhKfofy6Nwq7DXMzbTW766NqaILraqW4cDXm44FlcKYHMP0/hoOeqNOgC/+wtl0JFssy
DSK/Bq9XviBMDXzOu6kfHMungQHdRSxDY5+gTRW4Os4HTaxwjOXGeIcyRquIuGOQ3/iOlNXbgjlJ
iYuPt4si17mw/JOV4Lslmiem/+OsiRDNJmxXNUZ6R30sZMRhOMyLvouAj4hFQEQDx5Keg912UT7+
SjglpSmMBbvEgxfmLHT5Vql2Y96BDH3G9RrjAZIIZw7C8OMbOAwD6kpZd425/eUjrmCaOVxMeGdB
NnuH2aW1ZywrknccMQFsybvx/6/WvrT/r14nTfWSaPP83EJFVSAzG7iQax+2q0IuAMxos3Nn65kP
iFpwrEQJjSirVyp37tlua7hlvT3X9r8uaDWPVyilG/FMx1JrdxvOINq7YVK5jWzOveJv7FCBNesi
Ri67104gr6O/sHq3mTb8v+popHTbMclizml4HHPu+Ol5mtDW3LLsYlzlMuHw6/7bSEGXCHqpp8Oo
3iFJPtL8Z0S+mOexlXDQcsc1D5WO2prTTsGt5VEZ+uMT58NBCcdKmdqHvsQa4X0ZvHlEDGT9AlR7
Lxp40MJgb1yPcN8iZ5+0aSdtGmmAXCkMYzJxGzXufKuUpskeBASBjwdab6A5jNzjD3PXJBkrx3e0
cekZinT0VKDoYx7pc7fjVmar3gAOsSyYSV668ntpgNqff8McgI5vwXyAV8+NfIZqTx2jyIKyDyh9
K8ZXvEiKXdgDwMu3r1S0eKlPURx12PhAhVGnJcxkBSiQMnR2cPwy82iHdckMvQMyeMagVevdM8D7
frxOORKgGRx4WvKnch/uwYSBp8n38AX6mjNE7dzEY81PKhpsguk3aXSxMA1RL21d/FEGeya0WknA
XLfvkDEMQOpWsdsm4mdabg84miks4mV9aH/c21K8Uko7M/PwIyPL08R2VjKQVGFVo3VQMun1EjM3
mD5u4AqhOmWFU/wAr4v+Yae+7A2xpN3v5ncMsTDk31f4Hdy3e7b4+Go375UP1Pejh4uZ+SwuO92A
bSi4raEOO/mban/ucS7CsNz5/hXrY4XYhq4u88MuVcn0vger6kjkjfBaqbaMbEp+WCmHTaDSdjhZ
ShbZn7bf6Muac5OtvPuc2IzvYCoIGFajMdJZHY7LkvkpoQypf1pUbiIA/f3Fs0/M6XduSzuZzyNa
4FJqWixkJjaN2rSx05nGNq/Hk/fOVwrwpY1YWI8YlumZy1U6dkFmjyq0It1H08O7BrrRGEAgoEa7
OgfgTChjjuJ4C4g13CGprvvaVDaCwJko2B0TNaOQ7UCfxrp+7kTjY6bujOrGB8gvpDgSnvlWFPJr
Q7drAlV7b/L5LhXwelRchKixFl7bJtejlXbr61TZwb4ajIwEOGT+a7pTgYxYP4Em3KKfqWT1/xEa
f2ynqTTBx9s2jpBf4z6NKUeuIZUCMGoJdQkeJLPN7q/LefqbK3w66YzNoyV7iUQZu20uTLcW4/KU
fuFz6ZKCNetUaCAlsm4VGfWtsjLvVPVDWqeI6T3yefQMTlze4bQEqyA1oq4SF6Dmvj78cybGVcEL
Rn9EYJe+kTOYEuE/itiv9QU238BMTbaH2Rx671hVt2zSd9RUROVzpCG9T4RXYJeMInUKUHU+s7++
CUel8E8oDp0MNloWeYroOoX1xzt3QcLgcfMcwvRHP+mT1dx2qIslIYSVA9hkKM1qd5YqbpI2W8lt
7SYC3PZRRjNZGNdRtE9yrpGmTz8LoS5MAcJVdcL9EmPkiwydolDRLxIAVFC6bMP1s9lcls3nwsaM
hzzUn2W2sl7BkSmpHfwxEcea8iclYtSCjD3WLBmhOvUb2UdZho1BgvDJSofZR0xN3z53LyFj32IR
y7rIggNWI8WSJ1wN18Z10uaKUvoeNZrUj34FZ+dYQPHDCeJs+NdJpkH5j/P5kVnBRUXhqVn4DcdT
ANkCDny2yHi/LgE1U8VPf5gSrh664WcDdvO+oTmtnl5P1yRDDHktGYs26OqZ0efJYJNz8totTJgv
j7Y4B9xmApv2en8M60PiPIsH78D/FJ7diWyQaKiG0B2dEi0TSx1+nRJTdkQsOAAyh+tM9sJHEHUo
553t7ncwa1ix2u70t2qxHImKReSEtQ6I4EUUESBH9AR7hm3beJQ72IDczakLgZ3PD8VL4RY9Xjtm
HlGNwj8y7EFxJVm7TY8lYSz11aOOBuZfYRbypltGmFJrlaur71TZLaZtY6Na6z2ClvNS7BJ3oYT+
WzzJ/JvKJAnoY9hJPI1Lst86dV0Zaq+IZonq9e7Suk8A1dklaYX5GWpZ2rhqmkN0U4OVTCzRlZ+H
Xh3V9gxOiHhdigzNCD4kO5FX7cFPddIb1fFlf/E5RdbUlPDpfSjuFr+XPCK9T7OtsYmYx2tIMl2c
YRNXC4AtGoy4YMYmnDAsGHM9yy2o1/4R0TLlbc7cYKDR0An8HL2PNWjzjBB9ZQfzTR78tDeUrRjC
g2VmoDAVg9HD7qTRQyaJrFYgc16ipzOED4FlkO8ruYub0Rg9mNRoHeiVNL9DmQ8oaDgu7UZbfg9g
CS1ivH3GiFvQ16HxT9P4Zz0CGrf+roMCjO/H98+e+mWOx/EUe0KbllP56zLLGUhQH0DfFMktQzRA
LLs6MnwWcHd/IR8gWTy6RL3aHlTWQAXc0Gn11VuIjsLaTj8kOK+JrWZW2fAB0+LPeNqwz0z5Q93P
N/8XqBL6H9nQRlQsZZWGq9yAnTdQb/cSs436yYCQY6NIKOfqXDOUqOuqczuFkRBeFFLbQlQYIZj/
GIRm5BRxFkAoI52S+0qhbfS/e3t5rq495B9jgj0h7FHJynmDZkONIU1wcd60Ck+kHewq+VGzzZHE
UvN+KQr+P/mb6lgW+wj3ZjI8E0E8xlaUi5Z/yFTHZ9QYC1bOq3leoIdpFAMHqTh09UrMp7l/XvAZ
c8D1kfjXQTf/3Y808O3z21gGCcO+hTAWix7IFFBIj5W4raRqcNAzvsq2zM8ZwiPc2Ho78SF4UbZZ
BuIl9ar/NPSwf6/mxviu44llNOoolYc63gb1HdHxVPkesSX2qDrR9mccTdir2FIMMWGUs3y8Ki4Y
d/66iM3ngxRtjj539mA9VQgU/TNVjbr1AmYu9V++ttEMVfuB+Hd4CrNWpqUfXfRtm8KZHq09P2RG
qtpYBq7nfRho3WVjTYGaEywUJxdaTZ5U7sHXD5eVAOq+paEy8P3xv8RhqSb5T4vL1ApR2eoGR3J2
z6R28QQZXZpKBL+Bq1KJtvDktaLzxThbyosT7/74ZUyn0cBAMoErZ986JOQRdzB9I7O7XCrxztPp
hN7zu/fpLTdDnKVg8WcqE5WhPakJ17G4pcxPnJ7EtkI9UGwmoLwwYi/NEbtTy91OigzvI1r6luhq
niMUXfBMJm9wF/jjJwGCw7eYbCt0lPJxT4/BpBP+mQlamn/QrkySlA9pIvflcOQdN8wrCquGyIVX
57yqYH4+DAJ+8xDahWMkf2l/zWAqiT6vr3emKIcgPALvZQ090X3bIvhzNJWay13SUEfveT8dNIev
vD2JA7KIqahEKNYx9acgn6zdBGstHWLCJmTkQcnc3l8i9shNWXYK+QlPPxOAvpgSPvtBz7eIn+Mw
KYAnjLipjPLRjxA6DSbworOq/BJZNnh/VbbAIcLMsFBsRSADWGuC1c+Nmf79edxjDHV2NhtZs4sm
AiDdxVjt+DBR7R5YV2PshmhFSYooZfc2EqmYrHXP0PKujOKfld7HFDISc/W+XGtd/M7MOa0BPoBE
MpZXf0k+/OquDPeZe1BJ7SyxUbeosWRQ0lpT+QSFQvlOjtGDTx18sDzrG7CadF5NFxZCEnGu//UE
wuKy5hYBOvu4Xg0wSp9StTEc4zWAdEyaHq6bvcuYFLxiFQi//rPymiT/t3G0WoHBwb4FbKeRFJXd
rc06Vo44IhKAQmWK3cconhEBzwcQdNAOJAJhWJvRsRTOxiQAiwiJn8h2KWocEHJ6vpbN8KQMlB/4
ZKGPk0aSbRraxz9Zx1Y7re8f3Qr3PiYfUN9u3XYBwAwMfNizRg2464ZOIqbQSvTsnurXozY/qCcT
THkzROTKgR2xMfgSdE+9Y2hnK8Z1I4/GbunOTudJHC3r9Vc9FnWsxzU/rwJM2zn/PFjDjPMYbDGF
zpySuATt2mVWQcky+cYeDpaTDqqii/cd9keU3xzRPVx0syiaVnxxOSc7xaH1SNm4UKQuFVZ7f/dG
091/JjwZl+N6k9ZlzjXT8poZx9nsUqQlnEpakwtkowgaAIeqZQGc3I8bZ0xDfh5Y5fkRomZg+miB
d8iu0ZiAj+nN1jbTnTJVWi8n36vjNTkU49RDuCccBM10TdS+gO51IjwwXzl5+XBtJdckmm5tHBsc
itLmLwb2bkMrP2p8syiudXZndeRFU9eXXiLh25spxL3dJcJPsj3vp/S8taB66nW3duw8mny0kik+
XGYmChPQaPPxGNOn29uEUXvbyFFMr384ZVAStaiCZAN9wcHxst18S5Xt/BGzNzrW+9OVlptw3YCG
3Am1yUHM2o/pWbl7oCmpxm3fTpus3SgJk0MqjxYcHBbAQWcCa3/saSnGPFyhCDWdxju439n7pHdV
oAcpjXmNl6wb6pIvXrtW94P16tLsNbmpP5yjdfVHlg1KeNkrC/gg2MYFCD5Zv91GH045USamWyRc
YzK2frd8KjpdXPV8XY8K6giOMHu8kIN2moMsGnkNcMRRCTj38F3s23s8BQGlaFZc3AGVsboYY9Pb
gwFUUUGjXs7SreQzSZioZRl4E3oHbI+V9ZS6JmfkjW/BbcaS+hrw19mrBLyE/A0L2cy6rCe51WJj
F83FJ/VEntu/IJIiCi4ARbe5hLOJFh2dECIkVvdVUt4cbKzKJhJo90ULEKNc7ml1lxxmUNMPG28i
azA6j17VvcnAsLTexf0XQFzxZnjMh4a2Q9RYacFskZW1M6FMhbNUox1RNHC5GgNRuCAJX4At3uln
bFqwKUluYntKuR73rhxnKpPCgXnQANzvExgy+eqz7vSjoPEcQckL8+0bXkcb9bCl7J6g8RB1fO3N
paPAfxGFifqhqEhSJJ/dR+xchZ+NwwWMcGOfZYQtHNW5bvrPHasfFh4NSSds/Ql73NjZOi8QEByI
g6B5gU1Z95mp7NpzbGWgu94g+pzjRVPr53yVL4BBOvaAQy1ZFI1wYVgTTGD1j6+8fWC6mSYdKcuD
WhqSZFRpz92Ayl7/xXE5a0ZB4f5LggP9npi2++d5/F6K/1AG0tY9uw29+6ODOYZqfVKUmhp/gFJY
DMDLaEY2n1mo1MEMd2Hb+IVlq5/i+djyIogzkUtc+VcXvAkea8jF4TdR97TmYdRL6BJrsg1CS7mY
0DdSvHHWPBLcgOjRC/888ECQZiIFmMS+hcBOEAulg88sHvixp1aubICLQEUedAfJHaJ5JQkkZWR2
Y5JWJfaklpTxrzQHm7Ayh0gnoeZResj5L45PSMs5/ijh3Uge2Lb+Z+/Wlp63+RPwKK+WbOAEnXtT
lKNlVOoogEzgD6fbGDGOAYL7I/wKRATKbks1IS3lslSs08tvHL9QnuNwABioCpkjKAUOzxT3fnax
z1S0x1DoT5Cy3Tzz217e9bzkGGR40Vsh5mN5Aa27VplBNYeLbZ9cECJZR0bJU2te+OD2fTdriGvv
oDdmfeHdwAdTRS4nMhr+KvtVzVt3RnAdcQzPSQUG+xdWbOGjlkjduoJHj6JzBhkfmNwHP7M5Lt7F
hTxLkSrVzyAuycGM25F6+UJiw1VYM+SO3obecd2SaZVgaHI9HDG+PmeiQhirkJz1MO8xflPX5N5x
QeE5CTA6gz5rJty2lWWgXYHlTv37UQCNrRJ8D0+TD1QRnoaOexeh4ohHp8xJYX762ze9EcTudIO0
8VNukRRsER/obAcUPnUXDZNu/gdqzDNFkl56s+bb4oTL4lVdq+tKniNFqZYvCrqdsGdlW+c4o8XK
YkduJsT4+jjO/dAiM8IFyQhGDSgZXA+BGqsjcgN7DG09PEiLwApzR5l+H3idu2HtbowYZKmZ90Go
3jLEbOxFU7sDpgPyMMEc5OO9AjAN39fPxd+R2CCQoLgQixkp6n2qPIAIu3D/S8WUXjGqfd1pxDYS
BA7WCFT0IgOAKVQ4Hrt82OKTaAbwPuGU6tCURHi3/TSUwlF1M+N+moHVUaPGBmwXuk8cajFUvApY
V0Bmf7L2p7bc1Xg3wl/SEdiTzUE/KaIIkp2jH+KrMmROZofytIJVk2bTeGMsxcJkJXGUxEAJXYS8
8Jgg/qMJmHLdLLNrAwxepUP2qbcXb0io/ociq1yHbVbi1DcVWEMaceQxTOpng22z7YOK+g1vRAD4
7+wT3G77uOQQmWwLlfA7zdusZauGX3CNYtOkB1VEi9aWeKdPclyXI9P9AHMcC3bFz6519nBPtdSB
GfmkyTafVPzIpHYY5bWtosn76HKC2pI4tSjwUeb9WracOePNsg9BSTSYHvK3EU2Za153uIatPXoz
DHvard3rYIiyH5DKJp1i0CbrGyGAsAevJmx9nr1JHXxpoOULuBYb6D5Pg7lPtNLYrWxDtMIorYzc
uDqxqR8BXWJ5KJ35vhVWA4fPWXBh0wbHIgbIQlvtdG01McHgARGCXSbQ79mIWTVID4BeSGxs9nB1
KZOw4zW8T+ifDMonXl3eULb0mjcxg4oJX3+hmGbrtYtD1QX7ovkM66OdwSj520sjBPDFOW8g0Ikp
l1SGf+Uv60PApkZpI1aI/bF1a2JRB+wM0FZlPFNxl+ZeqtCYWmso3/KnBTJwzwAe9W+99G00g0lp
54bOgdD3VvcZ/jpah5cPWB9wWLh7OEkflsgFqCrlEG3CyzqOOupd51TSqL2ZNPKUYIwPXPxb5qwI
fFpIif2p72GcaHvALMuLzOeo97npFsai008t4ZdlnIY/a+HrztVFD52pnEpY/RRvmqdv2Xz3U/sJ
r1IW4sTScHf8wLr0DzLOWugumQoCtcSPcVLDLhzm4kpqG1DMjchkQ7fxWoEp6Skvpypefmq97/pA
ZmMSONXqMXyqpWbFw4X9gL57Ig28CK7S6Zn1Ff93dOme8M9YJwqm+helh4ZpmrwdbiLPaTdNjR7Q
w/9dC/9pC6rpuoE4/5zrWm4zIvVw4uAHhDnce5DE5stYDWLgSd1I5QFtzER3G/makl34k2K9HCkS
87PcAI0QTzgig8mtci8PE1VohI1B3vCguiEn0UmAeT1lK9lm+2pv615RmebWA4ltGtQdjTdXMrox
eo+KGptjrOjJz7y2r/nHTDJPV8w9j3Pw7MLIX2yAO5RAAO5ByCGyG69Q6ywN9O/yI9fwUaDp9Obc
POqnaz60VFS3GrGm2gWzO2A9p27P2jWyTmax1bDYZG/paZecBBa98EYdZVpUulLudRvXYESvQI2M
OLyHKfeGlzgck2X1F7qHWpRF4MK5AfePHCYcZPEQvFpogurx813gk/jZ9rod4sKjTHs8qJ5ft07m
I+961UxgM5c9JSbdxtn2vVyZi2sp+Mqk/JeMc3VMIDgHxEIks/0RG9a3jLgwV3h3yUaj2rPcxjJw
5VZ8toywvPxHUmeL/TgBj5cGy5y2jHG9pCeEjFVoZJ4a3ZWYTrgggImg6iIJ4Ej2XTIMuAR9LxUL
b7FKSxIi5pCl99g2GMiDU2Tygp2HMqVaMvUgP+ovqUuDV0tix5GbKRdc8V4qqQBlvxvYjaPW+/Ja
P1xGPOJ4DFDAcGYB6jPMcr5o8mpBFMKI5oUTSzjPeSfgcYjjEFeXAi4uiHhVxidil7odLSJ3qSL/
HkR1UIeOcyy6UwByvXNAqcQM7LH6b3BbQoFDS/5g5YY+XJCEhPuZQWHlYEY31/yibdwGPjaJZ5eY
jbfSKLSwwPkyPA300jLCObXZuQdK+nVFt5fPtBc+i+Q01yeRMZtB+5o2t4hdRkVgoBggljo6hcjT
vRH2Ns5jAVsQ/uRl/ElThAhn1YdJG8F/M0Rn2B4nr5HO76EKIKKj2Kn4OdHRDNj2ErLb0nxAt/6c
jvNnoLS4rIAY06UaMUkdl8po6BIcPP50wsP2domLXGTsfiYKPcN6+0QvOrIhMAZFV8ICYnykIemi
ebJhzBLwsquiS4u9F62C4xtY3G7zqMF9geRQMBO3X2w1jnyLjbidvZ1il6TNtTGHVLAJ0Z/PFKzh
pKFTdUcKB0Ic52ojXYvwL0C9NEEKjbJIapO6LIsqENzDkvpXoQzFjOyLZ+d98+UJZjJAmcJE3tV1
xGISwzHhi2qdmvJhPXsbgiQpl2qDe2i7sd3FtDWVClZS+2e7QMMytHIduNEjRkuCj2ZJC61ZKpnD
8/+bGWugrwO8Thga0ghWoBxHXsZd9hW+nYRJe1Gu6HbD+nPdM1yN6wo9PYbRK9ALVVvimgH2+ll6
Pw6jFgS/uTQgOZSHn5SylbrM+946ywg2cxp7wzZew+VkjwJyhaYnPSAgwuAR/t43ZGxydKI1L9bQ
5VEVede3SX2s+NjnDFfM/7Z/A+0Tav7avU4UZMdFWWP4e/qKjycZ/Wy5Y83ACL+NYGdtB7qKaiDT
vJw1Q2fIk3AFLdysazbufm5Ek4ucqAaH2Ou1sYX3i1O8MJdbUO8S/wwjtQGsq3I7ZhkUJZIh42lO
wI3jYHdvLv6huW6WRPtVIuCvT+7JwLSYaDFXhU9R1l+2GFFXvo5b/AX9uDHhf2lLnvrVRdPNiFVW
+WAuTWjbdIutvlCKCG7cSTwP7H+n0wPjSiVczhbbPfwchk0wxSe4NKJAj5nxv2qiru8gn4lZwk/K
EdNwToFFMogSDEz6SnYRfyaNMdhDcU2Ja2mmlygJDg9JJtBh/yHe52Vr2OBa3d1aOHjU6iMArMSH
1B14gHLAbO08wI8Xpy+a/qvrnGFcN8k42A5iAUDs7rDQjz01axaxefpF8YiB2iIzngt7d7W6AGDw
4qKm+oRxY+5Y39vwkKF12HvXEquQe7et+wJMEJUtcUoC4AN7Bg/HDVY0d0y7DGlKn4brr/vqcXnb
NWYVlziBDYN8LgCcxjegGORfVhJxC8vIGA3ZS3JgxD0nfzgFGRic7GxS228Y06EckbVYFAg1umVn
ZsHXFw5yJlWHB+nxz11GW7Z619JLsRIqXBnreKy+3oJdPkPyO3OYPTok0j3BzaeWOmyp+62r8nZi
QXncWFvrZvA73HuC2rBNzGsIJLkiWcUhjeJFvUeiPrw/qjjhukKJBIvmWaaDiY4cFp/fS4SeZuih
4YhfQ+EC0ORFS1GeOx7N9JqeDTavRhJM7AjKag0cKhak+5ULB3oW+KNPsurbduitAQFUwGEOgYN6
6BgCRWq1XEXVRBWf02omtwRruC/aE6TUWK+s/CS0/f/90MsligL3JHZHV9yyRvvOad2J6zrJFd+N
Fgf3FhSsbBDnatMI4TnzJyPWKcBFJr1A8jXOHeOFX8miXBy2Hd4e5HxSaychMVDKLP4gTACUubSk
Jw1lLoKfGtLFhW1qwmDWdth5YDpklKJ9kafApIkV9RVMKpilA00nXKUm9TB9CjfA9FT8k0n8DwF5
izHnqP5p3KKq/1G942pt7t0L7jCHtJmmNj2ekwY9fNGBRNpqdJyKnadWjj2EzkTsj5iZxIOGFvwZ
zImdsb46/rwXrmmlJ8JTDOKMNbEcMKAG85ovjPdrqoeet0GTLouhx6fNipRFfTR8w+tFp9KOcyr6
xj11BIQWVd95AtNPFYqQeh/gj+5ySJ1Xrp+pWm97q3guvztIy4d+XLMHRyJhwEJPtgGOX1HDygdE
/pXmo4GNcm215iFzPyY03y5vFCv5B7iIG5YhZ1ozSY2HtNKDEs5RCIoSdwP+4BCN87yeLwRJ8g2d
eQEfThifeYPh8BUOLnYYnenADoNkKPrnPvqWxl8FjrdmsSV1XK3aod5unPRoPRswAE1D+sUgrLKI
hNBRHdx9Xqnlvr5IL7VFOlCn5jEa/rlku+7wQxxKAYAZE3sY6mt+ifip6xyOShPtRHRwIotCQ7pM
95gmWsfh/IElV/PLvBFJ6Qhrnwl4iX+zhoVWKJtLYN5NYC1/KIg5kMs5zi+JLKUI8mkUFXMr3c41
ToVBI68kw8JcdsDT3wT6p3GNwaU0/m2Ekha8nVfFfoqezRCt+9tGjtigWfmy9sNMA1k2dCr9uA+N
a0Xl7U4KlvEEUJ+Q1myN9bKAIk8L3IM3A2pM7ItzWdEfuLelIdmhHRKHUIR7gGKdS4obrfrDgRoF
nQAPHwtwNeeM2TBAhJQZGUco9fW2itcAo0IYa7Nax2fHWTLWv5Ho+maB+JbyXE2vyHxGiAurEHPp
VDTdpSgIj7C8/g+Ja/zZ8AEAKNvEZBOO+7LuS/EaXmAddLb/0V3nipwcL9Bl6+R+WUYPFZJSh27f
g4jdUHnJEbIIk1jjcopoFunc2KaAa6VFIQ3qtpXHJscoiLgjzOWn9AuFEyDQJgFXMgwfe0uExiWs
Th+MjKN5YmBE7HXqVqS0uJJCzre3YG5rTEg/AnkonepXi1PQcnOBLxpBI6PdnGlNZZjeLdH3Q/Ec
opgYkd/6Xc7T9gRl9rnr2E5IzhmLMxhQQM4Egg1F2wUzTV7k2DXAadnBExH9Zv2cafr851oyh98k
Q2Tp0ipxFBp20A4v8N/CYVbXsUCAFSFwnhVVDOR0BsvLWT2UBWKe7hs+4PlZkVg0txf3XprNVEZd
z3W00leR+uk1Wtfzhwt/kO1qVtqGxZp8/lAexfrdm2FwkyGroMXISk6ftc4mHaeo8BInhLETdQQq
eUSdIcZElDoJ1eJQ6L03t2coOvmdjqVbIJVGllWROCTyGdNDwG801/lNscJHLUiGw4AwpqgFDMLN
jV6o4SFUOwsmJVayL7Htel7UdpHHGpfC8KaCJHf5RIgVa2ZUDpLrf6ZC3SolqeatTIS18rj743iI
0Za7KSdtjvbLBno4ARFcG0qFSqyCpRGAJjdMQKnHygZ8/meSS+9sixNvHqZ8UvCkPdSu2mTCqVDm
CZ1wwwwOtSaQyHVenjRgXWYIUj1Y4ojuJ5ImUmX4lYbQVtXDfIqLIBqVvLpz2TaTGBG3lc1Mhj//
F0JDtdSOaJltNFZVjDmSwtM9ibZB5I4wqASxYx48WvonNwKX4R4kzLxakaCd5XQ1fiuKzkPMLZHp
a7BPhrL7unGELORnCujpg9rPfXksUmTI9NQzIrZZQkW42kOXEyovVM+0QpXMNJ0dEqLYSfR9g/hl
55uTDEFwRTKnPlx7zlFQE7cEcXRjn/YB+Hz0JawH6yY/zmUjwjnDl/C0LV/11QtDnH4jjQSUJtEI
p4jEaKPjWdihOmWg2tJTkWJcyAaeg95auiHX8zdGy/aHag2gGughXYbBBdhd1TXMdJupD+DgS+CS
sLGTQGT59BJ1S5qzFXoUZPp6BF79SaigAt3eqz2W6iFlHSgwR0UIrHxP/EqXK3jRZ1m0aKiQ5+3g
lp8PXZLZ02ltTbqGWbK3PBpOB56JCGd3KhAsUkhuzkEeDSrN0QgYCUtRV5zCLLJHqyuM1gzDowjB
zAcYCvn2q+Jbc2u1e1t8UbSyjbvhiRdyb6/vzZQIMUdi7kw7KQ4Wo75WgdRtsXAw2lGWQaT5O3/M
HR1bhk5aUzmX/mN1kNzX/RN/HJM+Hkf0pEXuN7z9ihHyWLetPZ0xkkmJ4gI/Ac0O6gKQiqPChP2A
LeDN9Ll5oW0bdIe02LW427jatpVYtfH5Ije4LHqdTVbLSWzIq7apScmqOGK4TffuiIlyFuLi/nuY
gTsWzffCNOEsFRInfJsRi1y+XRN9PhbUrhg43g/clNXAGoQBvOSTc48Ga9y2kXrofUg1pBPFjdna
4K/3gaarmJWStyXWE/6lnoc1O6dRx+z4Ig/Scj+9nPJ0Fv8apTnXGVM8yNWU2zOxmKA3VNiK/3eg
9YSp0VoYoY7cJy7EK91PWNi9wddJyItJx42ucxVmI9GEjim8b7XmBCmkE9ePl6ReQsnVgwAOcvrC
VsH9JkRMxnICM5r+F/Q6IEA/GgraDor3HWo5Dcmmqm69eSGxFmNHXnjGTD1YPaKgrGPMqV+0dZSp
9l1s+ITBtZWjyZ8lYmwAqZZtmdpcknHfcYrNmf4QE7dVh3XRk/z59GLNVzT6Upkf91Fz3ERNi26/
qbTqQ2LtKwWl99o/j+VunCeWr7qzSNUW4jNBnFRiXqCjs+K4SEGW0mS5iEeYH/zY3u2B6PJJB7rw
3WEfaXWoGw/jZdDO0Bma7q5GsFB8IbA6sz5N3ATwB+eceiCMNxlT3oAtUHPqyHOPVpf+cC/oyRPu
siyU4L73eOLDB1V0JTGW4amj/mUrJbgtNgRvulGbvYQ+gIABDpmu5SLPKU5NBylSIot+7t990xx+
N6lndz1JNKcJGkl+PhOFO4m2QVMzXb5L5YaO9vqtmDJMf7F4sENhWLFNtRYj/IIklr1vIoikC1jC
fmBCWZMiuQ7+ATJLCGuZyiVP5oL/D5rPHowV1er+wFG15Rz/qRK7Eseg15G9MvWTIqSU5hb996Mc
UBQ/uRkF+I5J+eGqoqNbUi3KHuEVhvywxeDnnDJib+duOiK9mRQUKLStuk4WrKVWKkFFli9nWuom
k/3u2x4Ubvvb8MDOfkAO8l0KowcJOSytJSTF05ModTcORnaxf0Qf0TDVEU4mtFUIzEgq13Sta+mp
60IZaahmuF/7bt8lZRzSOc9GlMIPg2QKHChZPSpKML44g88DgOAAz2glWLzQNG2VfsJyUKApovuA
MgTqFu1WIn5/sAzSHhaULvt7A4AbLWIxV9YfxkS4fk8cE84eogYClEocENBvGGvyzFIke1ulJTop
llgUvi9Yv3Tw5luX+vg+JH/Y96VCX9ZoT4f/O+X4hpTuNI5CBknSowOA+sWNk/5Xp8U7Lu9HLYgX
egzujTaoNdcFNmtym3pdZpYl6nxro8GGZxKeW6ZlSwc8gd6qTf8ucyvjijOs/0cGo/dBuFHIsjZH
mT1fuNum4rmA2oA+GcrJMPjz0ERWcIhE+HwMhDHQn0OuOLTSuSCfVg79a+0m+ETrNvd+Y3S4CYeN
Pwc6oLjtMd/1n3BTwjkqpJMQ5ULX82UpWdnxTYRmeePX+kFupjdy/THLlkUwWHk82EAqalAFfmKN
mTrJYxUu8PCGdTboOL6FmTrMeeXao1NAoXSJfTZrldVGRKZv7cQ98CKj0jjP8H/1JRu7V+xv9fY4
24SmPxd38a/pgv77ITreqGTFdyXUG02J8iyy1RadreMmr9XFR4fygX7rar1l9B0m604CawUMHClK
9NcqQ8f4r9VSJDwfGg9ZxuLn3lhQPSzZXUgE/sYOvLTDAEZhO2/SAjWJOOkeZvpWbJvWZ66DqR6w
ThUc+9X+bgERGuLTJHZmtrRJmKtmAXEXji8/rroNwSVzi7SP3srlhK1gIKNMe96gDDegJ28IRk/1
pa/9Q0Yqz4MbNquLmtkyz4aEAeDUuem8bXYNlBqoHBsryYLwh0MwmVasgN5dG9oMqxisWo4HT7VM
4uhm7bPVCQy9iaFJHtBRlch+WwT2yc55p7rqZtAdTL7niGb0bX2HJWBK8DUy04p+IpzLc4l+tK6Y
nvyJTVccu71Elz4CzoQHxm2DiTJeXQFf4CDQOrT15TITjg6Nm+X+Ywa34IY/GDQjkFfNMfO+wwot
gN9mywR5/Zjjg9xIVvZst2X7fsh/4jI5lsbgEhQ1XtdXswqMnTFpGq6akh6hm4QTI6oNMdnONTeI
ZjRYod0AgIWTZITY3Jl/OHPx8Xk9ICyzfZfm0o2saimszuG0igm2c4OPWpD12Bxp1g/lr0WEqwRG
B8XwtnbXYUv4erINGRbhIPqpeEgRM33f5iAn0JvMqzaa+Cz698kYNgA7nz+YIi1HAKHIsXyF0t2S
RXUbOG+JMlPsWMGP+B9++dqYsR0O5I1FlWS7Rm//ruHOF9QYVEbuD2L3HqrFxl/1BvBA8stmayLp
TS6yQlBHWN1stFwBQvtpqhWSksu3jXlPH51PWaLGlqz1OzEcZ48cMY10KukOn5ggpVtXCIOaeJAK
DlaiTUPTXKpZVXyHHN+kmEeeA1t+UQdUKRRJsvYC32ybJuwBlEJKpXdiTNyggolpDy/Gc7eWo/0D
g4xMctQdwAlonjU6QuRqRvMqtj3c1tPxvz8n3Y3la97peZTWYpW9CmCnGuFzbA2n5LrY76XpvGTJ
VIRTK6E5ttaNbMA0JPbGSCPrc2Xz7m15aBCHYdoWsDHdRnOQGow+1ebn/Rt1Nyztn579mINCHBoR
biUF3L8gDD6ZCq2vPBE+Iy9I89jlTEQccXEWC5vWBgucPmysRxs1sXytcHgsc1AHta1GF5FFJ+Gj
xJm2cENCQsd4FrWspFBnOS6jtmcXz63hJ6rZSuMDLyoG/It35dmwK4Lor8xFMbRadc3LRcvDr2Sa
IM8wZYM6IEAdI34DbOdbrXGxLDnncpNIM4QhWP/ifn0W/nnQnj/UWukoeX8PhmhSQnGBTc01Klkl
kYxpEbQP7dwa0rNBzTiEU8GqtpEOwFuwpPyCRg428zmfFzDHoxkfoFi9BneAJRqZ1eydKAjJTrtx
D2gpi9sgjrrzdI6h+W+DTQ+PPi4gO9FB/V5cYvWdJUnRK0rP5s2affWg8jl+C1d5lN6UmD8LFjFq
hih7lEulCEpbncgiFJvIFcW3PafmpjCmz0FUPlhvU9FUJncAcfJFKX+E2c5m04qleryQrvuLuKwd
MZCgmndZjvYQGkPR+uzkHjXYko3wPDTWNJebW4SUSrfjaKW6DGLQP4sRLN29uZ0MUeTFrHHxCSFR
wdD6jp2lhe7ytjpSVOheHgnfN6syDpZ8kzlQhg1yZcpn0J1m1/yX6hWmheoJVfXXdQqqaU5xU003
9Fook1+ywZB1UN+NXCEiJNH+jB2GmOdKQk2iWFMDy33butllGU8dN3GgG6LC92NuW/BJ78tKtOd4
LLaKFHCfrzfZjcGKtPBBSQ9r4WwxpWZxYncWbyiqwCW2ZKX2ayV/dWogZk8UdKVmttnPLlQI3ASP
RYHoDggD7uOnD7WlTft9SB8Sti1hBKII3nJ3a2nw53vlv5d3oSghP6HUe2dcQEYFyaQADw8FhW1U
BNo/MpWStmDnKnGL4NBt8XNC+W1kWjNbtmfdmaRAZRWJCSZPwi2OxaljYmURgUCWHcQodl5VVihP
9XaoRwvEe0KoNv7URrk7Sa+zJ8xCCoFOSuAqv+qibvPr3PcjyCzeC3kgeqeSjeIwAcpBvZYMzAdH
Vup7H8oDgKYn5KfkHGlF+twqT43hz1FImX75dtsXDTHP8GkFpBylkGSBkkmVEfMUV+9PRZhdD4zs
1AtTvRp/qSYvjWoMA9h7kWr/Kk8BfZhT7yaOS5CkjG3PaQMWP+/IG8gTocErqLGP8PW5AZvqPalg
01s/lBtPWrCyHeQ6AWcpALNdBVbqNIEEraSy/fKxOaL6mcEO2wkYCpkHoEdBQK3fLQCnheI4DQSl
yPUwOWBqq8XsndyltcxDonDP/qlrsie1TRdRvxfYxW9rvMHYGgezWFhe8n8AyyXX3bJ6CEHsfvFC
yoEMI9EJoA6SBDItb10rQLPF5Cla41TVH9gqjglWRbpC6NWk+UVAp4K9HoU8Xyo25UDGFohV75G/
4v1O5GMawD6zzovFq7f+wvjOT54SDIyhczHj2iymAaUiJHz0jxbbPpeJK+WBIEj/QHDsjx+QawFl
SLthHkGaTuLnooz8dZMWgvuaRDOEVJ6FoGNvQea3hmkF6Nqo0N0pyCJ75ISdK7PnGkP/ur0rdygG
fEV8Lk7EI/FAsoJXfrKPpuVw6ejFzZ9fl+NsCLUmDz3YpW1cS09QhHYFUl9bPwgsOiXLJruBKqM6
etZGHXLc88Q87dekLG2+wOQm9azRnDs7m7XorPFN9QBsAZQsUgoBCgIlviipskERd57FD5ZtpkcK
8xs7H8Dv87N17jWGk3C3JOU+nSiNi94fDF6pZ9B50N4Q3AGbEWc/62W3PmAm/U/MgJARnxqF7Wsh
aLffIju2+bkAoMOjWW+Blp85K3VJXhAoqM/EZBim79hUZPCXHfWV5HZONpOPwdSkSd3LBvsculwx
R/T/Ji2vw8RifhmYXvgrFACPIWdj8MkxYGkZ2wlujG3D4z8YfX6GH+8MLCpsOgNmVGwRPmwX1s+X
vUBzwpPtZqNbAwHoqserCOBPVt1Ta6OC4Yx1LIQG8q7vLvM8sPBpFA3p9SkOUfifPbd5JI4mK4WL
UdS4Rg2amrFhDw9K5QWV/f/Zcp6YAWLk+Mm+AwyKD6VJdaodC3zZkaktxleO8uES023/JpUKKGZI
b3FDKkkzhtaLi7VmiR349hVqmTe9YUUrzfW5zExKteLOkbBZMo7uQMeEt8OfJHQah9uz6dAVXMWO
8cdNtvaLtTkmb4UqMQCwxlhSZ6S4JV6atTszt+OxosavKdXkmXS92BTPmbjhi9OmqcS7J/j9zEJs
uSfeE6QF3YNxxjLINfMo/Q10NFD7mH7dHBvlh5Hn+QIJ0tOPu7lH9oZU99kU1Y5bpmZiBkj7Vcbr
/MoF4WA1D8ZbpuoPM5X7H4chtHSYeuqPfiP9gw1UdwaegTm9yWwooiZCOxR0hkNsqaUMu2h17Qup
Y1BFJLCWY0D9O6iY9v4ZzVAMoeOiNGp7LHGFoqRbxzBeVrt4OgUIokOfPTA20fKmqJ/tqH5fJphA
VJIA51t+cxfu6hnL1GMBdvhkV+MndUv2NmGR0uGhgM7lnPAJ7oKhXm9cM1gbYfl5ipImdae3BXYd
N10UFhNihiIfd4FJ6RbQcT7KNOykKWPj6hSgUX9wM9d4uo3ZWfo0RZ78WOzQ3vBGH5Gso5j+Fwnv
TdBWBNXrMbcnQVhEl86nnpLsbNe9Fhea0bvRJ2bkHVm4KA0RhEus7YWtIfc5GlCCwtnLHH8D+CMR
TJ+2jIIx8lkokO3mOCzmsiIWGAg4vfWKPpws3/Zb+HDVtA6yP+7ks5VVLotglvsbkUcVdKuS7Kbl
CPmSr4NT8y4eUGkSe+1dEngRTHmXDEYwXpBLZuxm3eXbkDT226iQQ6UFVdsK6Ep2BT2v61CxwIkW
0hVdVczQkxur8MaDCAGr/QcN5r9uJCMGQV2zt4AoDwF0uHwxNaf8AwInGKjiP1t58+tV2AjC6dUT
0z4RowT8Ej6QJzAiRQzIAXAFK6t0UDKM8RkgYEEAm8ZUNC22IkuQiqObf3Afa6r6cjy+nMvc6yXh
j+rqZbNM3qpRQ7axyHW0zCr7Jt9PFJTro4Lhoo4WIgL5wlIa70VNkyX2qnPjhtE6oskWCPwny6GZ
UTB7vLiy5EynNGI+E0KC3kvrhQz6QcFiUW/WqfyZQjeRE+ugnqVkY9DbF6fNX9xKAvjB9pkI+QHx
iSwWXmv/WZ5pofwmJ6AqnRrKTfVjQmsNFatFtVZ98oOWqsqAo570TfYR7nLLYP3xxwjIlB5m2A6F
frn4/OqkXb/d/GRqwoh606egNn8kD51abn7UAvm1Fo4M/+Q8Gr8QgDyK7pIOnYyc9M2Kzq8exAdX
/7J0UFReOtRZo1IRE59S3D84fdFmAvwpCz56Yv0ACn6P5v4DweKBiWir2rIO2TTfj7Wn0euPURNy
GJw/d1h7DuFR5cE2Ib7qJak8wxgb1W6PSTQ/uUFeutQcXyKPu4m9bXQzzYR7Sz0hAtnqpUul66MH
Ui3OHri8Zrka6k5kBuT7XOMf1wbJLNjmpJUr1wLVrnWt2osKQC18VzUdIYZYKItftxUQwK2PFzQJ
8Ysei5Zwsa5yGV1MlzJHKDVkv3K8vFNASE3c+6KQVy9mrIYO3I9RD7VkhJP7ABhXwD2OL8uCbvPg
EV8X+HfGwxT1wVghKm/jSfDNOpl1Ku+LZiVd4iTCVpaAMJ7IfwWWKoMUDNelWetu+sqOADOHr6wo
xY3JsLavYPmj3bOS+i5mh0tqle2pqco4CvjpaXxamNik9bMTsvl0hne0/1Me4rDnAs0LrTvjz9df
7UhKW5bAB0PXv6QSe3jQFp8VHP4FUk4vJbwVNpStZIBrgbyhcc4WzsZ5Xr7oOkLFdLaTX+5zgK2C
J2mBNerAYganHC/xhl5hxAdEuYLyseSh16aTwGvH6sbNZV84zjS8fqXrw9z2FatpxQSU2N9g0cp+
yZXR3LWJyMOQAG7WQA/Mbd08j7cjZvTuPNJppMMSHrANCim3yFdRQJTrs4m9Zj85cpagVcgb0w52
EN/MvFEmFyqNM4Oo8nem7uucno+ADqHkGxqCOHQOIETnWrMqc1AuT7x7DiaBkploY8+hxsSQbgPf
B6djNbtksxQ+CpX4ISW6sCeH8B7pWmhfvhXWoKFfxMN3P5niuW0w9F5nBsDqKILZ8W10PvsmGVW8
Gamo7pbpA60/0h2t5IUO5yP8dHbhxeRUzbV9/8oWFJHehBEJP2nCcrt4Tk5NsmwQnuW5OZ+w38m5
6dCrnjvxBplzg5T/iOpeVrdZq2pMtjy5OI9NLVA9jfpMObee0gOioIx+f3hzV9BmupQpme6dtA6Z
hrIhEL7ZgtRspZsXASP0ZEQc4gdHT2gniocKggvfEjDm02GxLtEin/eixVV326xGc5KkwlEcuZcj
yHN3ahmoBbnPhtnHje6WUwNgP2PBdJ+6qTZGVAHZk6vi908g8FthDCY8F7O/eGZu0uoCZqeH40Ib
3AjWS5YBcjzfaAW6TDDyHrMX7ohARiQ+3D3EeZIekUVthAneEFZGOFq2B4fB/XskxENbJiTVadbi
2KJG9pdlxJ9gtLNUgsR8DDRB0VHJFDTVB4STpfI2lLlthEe7vmdJEhvMw+Zxrbk5raE1aprmTgJv
gCm6z2/zbC49UDXtArZb8h1j1Ok+g1r0t+5OALoPSlmVx9twd/S4AhQyhVgIaq2d3+j9sY7ZCtFn
3XQcX3NlmVJI0IQ4JfVh5Z+tYYt38hoxNI0WatY+DAK14wEewzVRs/RlnrV+MAVSxcIOzQyQ+5MQ
7vpoP5VdvLtTvOdbetqIxuW74hrXxVbJLStWA81u5UrQVqh92E3p9QJbyE6wX1DEvGWQJZHOaAm8
GIYGzONSRD/oEgeWUes09lhyJi+u/UpPJZSQ41BHLe14ASQTlmOD0/GWQ66ye0TzZSFWF2xZEvo4
mOu+tjXru0TQgua8kJzIqMhfUXhs0LqsSYQjdcAVmW/tfJw2JO7sbFY7m0+G0MD1yHG5XyboXXte
hCZJXHEPCyFIkKYW8Oxo81+CVjZgDxQRIhoVoqzMnKHSGNj0SA/hWYuSjIPtm79Zv8BbaVUdT83f
MG61rjZPltr9s+1KOzMz8RpTZqqUSsWaTGIj0xpSCUdu6S/2WVEJlOcgUSiLQlYYZL6+Ce9AK9aT
Fk86xLgQbw95PdX2+XozBbUNIurZmVhwXflQwyohaxVBcsFDV4f+Sk0gngmD1KFVTlHTlt2MNWFw
UIwIq6nSW7TS6WuMaTFx11LrDp52gafYhkABh6T89a6hCr0gI4WmGkxMj/BcLGtq0JpPaKtbl1j9
BHpNIOQKUokrK8IXghIyXAhh4P/R1MrqcJzjCLit/xGoDWdxMeEEiV9BhknTTkGGJvrVWbPqP/Kn
m7Isstfh/kUhssLZQ8DTklRfE24qOOFNjUk8ZgEfVh5TsgK3ebs+/it0aLgDG3IoIw8byVRw30OC
q8TEOUPxlPGAP69XXHcaqlmr8DlLm9tJIEAsOfXkfnb6L6+Bhyaoj14MRB2+HRMfZm5TTHHtqj0x
SXpkt6f7yCvIIG2S5Uk79CVwMSF4WDODBWFN2FNvdgW4waguRu9+VfW09oB/Z/AgRVfgy+iJClIQ
VP+3BMowSULIILuoBxOYouk8fqpSFHY9aDdKFkKkbZrRU54I5DsVIF79JAbFvryeQKdc40UWN91M
d6FRFc8DhcmXCzIa24HzreGzIn36qhROcPp8IUNDTVs3VYeKj6FWWJdpHlqZ567+f0llPkRL/xBl
dCbg+IyU/ZZ0Uak+ZQ45+AsNLR3u/j1b5rM5GAGfWpa+1+p8uQcSC+uDH8vGEi4qohzU7pWem71+
6ZcwwI+nrsy7vNxI7x2iTzKz5VJFqslhl+8RD6EZM7wMhFIcEVrJc8cmCh9NaZzWdZmAkG6DcDQP
ZhAU3zvh0rYzEYv1SjAZyCrXwNyMjovNmPs4dhfDUN26kKThjyO7kq0h8TLUzwqU9TlOztJdIDbq
jC9tCCUd/n+3FWtUTqXJfp7ZwqpZ3i/SC9dluNwZXA/KmYbfEKT43SoYNNS5uV31ujKWLnx/laup
ZZCbNmnENmOUN1ZnyXx3wpgOpWB3vGie+ny4Aqu8N4FuxuMe2O3IgweDDQ/kbq03O891fMODwUqk
Z0S2z8rO5UJZVR8GuwELTOIrA753350zJZc2VP3+h5JXiFAf7zPf9gtMTIaCnZYPem+FRQkhji5R
0UyVG8S6jteIPMHtP7rcuzJCen4FhMSJtv8EZT35iuLGs3O19kMaiPU1QPfFX+WZ9v67ku9radw3
akCJGlMZsIwiEw3skJGu9zsLpm8TomITXhHJQZNXcQBTNvXxRs3wQdl3YIfvXE+5mP5yANDR3Ugp
YqGTmU1vayko1Bx2SqQtxHlyd8z2BuU4WaHlsVxQLO2bGeEKAuCUS7NcR3q2jUsNcdHURO06mYvs
A3gdvpsLa1PNQHjbFS2G9DSCa0oKycymXiNYHt/3cqLTHrLuXYkC316BqrKaOw5ViJDKS/XDmcOQ
WWKLrBgcJDZSGub6jnw5IYZSPnjQ3hs5ksP27s+qBY57JSl4OXV4TPq8wcu/xWvnpX+8mQXiN6CG
4EBLyorqLLR7+umLuRLaBODwTWc3M9qHYV4fiKZdDaYUw2rYXhN5V5VJcRSQgAIif8V4xpLSByn2
X7FQeIBY1E73PrMYED1PjcfGw1UQXCo3BfK76Ag+bWZ6Dgq0EaL6/LBaFwfbkeVxM5I3y75uGBgA
tIOzcm1oic86EN/n3XAPyEhI5fXr1Cw6G3MPLQrUk/ZbJcj48R4qSS6KX19qxoU3Dm33SVFWZMhO
XZFVvmXBIZPRK/0Hv7lJ1syZzYqcZY20/7kfaNMHzJT1F3OiRSjFeNCEzC9ZsydfW249MfIAiD13
SrrKG8dgNjLwKxgQrcB1Ry56O8PyxARIWN81WDSrSLfYEhfY8vqBY55RnkOqcU0brMyrrhxd/6N+
Wlbc1RIfVq0fBpAdl2/gVhLOGNIVcx1XRA8ALUK78L2CcivfC0jf+1WyBC9Bwex4LjIaDeoawswh
tIbAJV8NjAftB2AsXo4tcPErtPzbZ6xfUEhqA/zc5zBRlfZQ6T2qubd+MCD6U8woXnByhFsLMUe/
eM6TmtlQtc9m0nuKiMb7Iw6RMh6/dcG+sO2Y/52hh0tY/yEnO4tknoSAXfE+bxifnmkFyGmVimE/
cEQuILVPR9EoAX9Im0V7TpXg0Ko9ifzA0Lfw7FcwqVRtovWBG9NBQ+Yf0boZqDy11MWdDq0SHUJ5
+84HSP7qwI34R65tMVJEm54agVhK8KEZggiXgQJ1MSvCEuaTqWTVciHsPrLLPNXXqHuwco8VEkL9
5m+J0KqbKfWPnUFaS0ER1iPQmKHVzT+YS3bWb1A9fzMJliF1GDfH8XsV7A+bA6ztTKFntOQdYvFS
XeZkCsDYUtHTyp87UA2ASsVrWpECXQFkkCH8p3w2Qdv7js+EsvMHJgaMRIBNMvYQW+IEsBZAk+Cw
01MSsWxQQEt+TQHW6yjaS6mvqssZaU1tgQxqMsw3zgxn7vF5nOaLGkDVKNGI/0k9IcrG/m20Gyhz
hH1f0DsEHVBIM5WAHAIgKtd8TfLPHwQ74hp3xlthV4ElB7krZlMxWNjiyPVB3B2L/qAnntVX5owx
2FaHYNw6ze4xg6W/TG7mgI2VPIeFXBpll2pEGulvZu8pvANob4WV4SWjOYxS9pdolmgLmClKyXvk
0bTOpyVqlmFFryKo2CpbKhkjjd2bOHsMt5c0ALGOvvntN6EjDFbmVXx9r7PQUD/cJb2cfETch4qp
1Zq83RudFQecuRbDwK3MeBmnaz3+MuhNLdy6rOVHyaXRSy75HwE0a/DAd03HBQZWrtQ67axL5DRJ
hlbKYDX2d6tsYhfOmFQfGIzrhhEJtWXJrWI9R2J1w5Fv4NS9KWR7c9ScVw0/UD6Tfpm0FTIWgU2b
w6sLaUk/2yrN0VXHJw+0YCW8kQdVAiPFywYJp8Pa9pN0EzTlbS/HbOu7AFQiI4vWmqwwMdrzQuAR
VG4oaFpnUz9/CLGRGswOCZeALba0TIJXYUa+eBJR+Z0Xgzn5iiKAm5/8CyIrLliYtVsFV2QHKMxq
Ftu46z/5KYFtmjJug6DCWbiuwxj6NHlyopCSku3+BRFfQJTECCVnnEdmWHAly8eRB2e4Es6JiwBQ
nIJz4CLQ5pwEma/4etNVcp10bB3LMmxY2mV4BV4Boii+uicwA4Buq+EQ227HxYtXFk6xnA01+I/S
8g+lIIQN1mtfrg4bAA3aM5rAu7GHeeNoGl2Chyt0WlyExbcFCPtQPg10jeMNuH7gc6H2rfPUorZy
GRo46FXcPWvZzpFneTJvRznhV+fTRBeetCY1MYYX81u6TIOyh1FFamfoA5xFUrHbBoXUby5ayhb0
q4wUKESNdV6nzt3J7do27z/X5MilGdqHos+UBbyKjfOhLuu7nAwxl9W4piOuYjDtEbLpTMRlIZHc
Y/DvW0uUfkPEnJput1K63PLyUWTsrbXwk6wKiZKBTgigK2ifSTmf9AAJaR7CLYpQknRImJPEMIuc
n73+jr/n+7yFARWA8NyaQKbU5P8HPR54ooOinIRiOFhngIMHE+jo3NkUDuh/BHSmtUTJfJEkkdS2
Sw8o8DjBrzgUki0oWHpAvYpfm7LpH3Rm1eZVLvwfzUTr8M0XVutSSL4eDI5dactDICs8uVbxxs8+
raOm+/K+NiJgUXMwHj5zy5Fj1aZ3XCwXCsdoVccvvRANwt645NMoMM9Y0VCoxPfrg3kaipjfwxmu
mqI5X/ETiitRcDMHpSpRxIPPZRQPCpb6wQ3GRPJtK3guw+5F5WTCkeWC4sRVTQUwe75kknspg6NZ
HeLd3M7a+7Eb7amKwWvRDxktt8aRvJSqjdCJ64TyoMK+zbpiBiYpr52L2Y9Hbh+fgGIgoLCyfiZf
F89fMEYWMn6boQn39R2eIK6PSDXHo3kVEkp13J+Z1CNTUknCCGQNx9fPHIkq0wYa4ufeAIqPvfoc
aHDfeBK75OhOneFSwUIshoGADgXOiwlg5E8lQquI6VdlniTTP7VHWko7Lw+0Rk/Lq9LeVfP9NhUC
EZvhi2IMnw5tfxF4+uEpEtiEP9h37jhIC+vKhZjmYXAWf7NAszZzwsWB2Iiz/OI+jio9qc6R6c/D
YwhpmsSC7FhMdezCW22UEjKpzfn5D8PkAx84yrhJX4KOS8P4oZ/9lecIXyAvzwJn1k95FPqKoM4r
xteByFy8YX6VUPLvEclCUjioYGh5fkfsENU7uQiiVLcVwW8ETaiLvzPftnmqia2aQfeKUEKaFbAI
c5R+O4UGP3C56rkrr2kh8KO6J0GWcNK2Z7EXK2kOegBeualGga7z97dOVndgin5yYmmhLQeYQKAQ
1lws15BaV5CeJ0Xx7755zh7azYCTAY+/9f9XJPUDaXKByRJFjdsolOiBLnBFHRGVJ1URzRiyS2pb
4Sxuno4tEqDlgVeK5q6X9jPAAA9KeRCZD9PvMHOW+bQo/l9g49mwojrxKw2cTligjzhSKuZD0VMr
b8NVowXg4pEaaD5gMjPLfv8Tzr2XM9rLM2IKaSq2SSlivlsSGQCwy8ArhYnp8qGHBy3D7S1+xc4s
lZVPaNf8iDFkArghyQiun4/ZKpcctzsGvRmVfwDM36Dx8cDrd0k3P/ce/25eHWs2sqvEUGpkc2Ev
NcyequbgbtPcYGUAon64nPiTsqvBLz+5fTrcurTI2eLxGMhAHC0dBY7EsQkXyR+C9N21iJmOJ4p5
mZR/gxn0HQgMjRFbgNZXqr/B8kehhBvVUgbUZnza4Wr/5VGjdg14xjMvSU4Su52TFnLvhC8H0cKu
8/7uRJ7v9qwTxRHVc2Y5K8A/b7VT/trX4GbUvZE0VW4REvwJ9sZTD3ocouK7YfVvZsm1WDtlP7ZF
tYIVncA+1lRDr8FhHNE7KLy+NDhZNlUSPcBJcLOTzWFukimlDfXJYxKWwg8qErw33o+eRILv90JS
PRrnfPaebs42qNxKK0dGKmfIxn2khaY5r0gvenzn8Yr43Yyj5pz5Ed8S+Bhm4yIVWqLf2XcXlBqr
kLpRJjMkcQx0GobcpT/w7UA6DukoQr93eEWWE+gU9vc7z0xwHdxluDCcnbOBMNqRjNtH5oPnVI6o
caGbtUlZbzjTiCcRnb5CPB8XO9Xurn6aHhNgo3SJX1PpuqtMSA9J2Dm5fYCfNaG+PBTHktVCLqOp
OK1XQPWpWncvFfIUebgLwwybcXVvidQeiNjc/9y9vRAAWR6+uujdilUSy5ZeFnsDcg6+/hpCADz5
D+zDZeQE8pai6t6JnCF9bVFs+5kBXmKLwrIoN7+qekcKdVObiCZfoMfGxMLPH2cZXmT7euYCH90o
HxgUUUKZWEBxWwRzRANav7+HxjGgjf0UTjmTmPK85iIaFQlS8Cvaus3bWE5HVK8qwg5utfRQMbhP
rTZukL48IZwlRST+zpKVxeVwmg17XVHFWZbIC84i3lHEHF8B0scyvhInCUn7+0FRTJcExLUpqwDY
fv0khQ0BW35UKGJEIlsEmvPaRcPuAFOmr9ov16Ohmao8w/+oUU9CTNG0tF4fa5CflQER8NSW0H/6
uRyhQTthYZcMmjluhxrzgv9CJxYwhy2qqIoaHsQIkNw/rSHepA0GFt+x8rmaZy+TufzKK323EaeM
0iySwdgXbyEBx2vw28Ka0AmEUSFF4CU5VOJAQGTb60gVVjRSb1rGOb1kFnvm1p8X2tkwJeWSKRFk
vvI0d3dHeCn2XP8/IBMfvOToO9OOf7QnCWRWIgv39805hfcDIt1VVnAslns02YxBA8J2cEtkko90
Ylf+nNeMbfAu2dH0V2n7T/TQSRIgfWW4s3Ofc2lnr45g0T4zkQ7tfKosnY15E1yd3zijkYDkfpEj
LXtX8qLS16wYqOd0t/KF4YQ1/w/OIFWXYoqUxEHFJcUI5BtnX00WXuk4HhRmLV7BnF/sAUh3d+Hi
dKZ5xm7oiXNnn7yIhwLkKLpRODdX3hsZpHEHZSeIphoxETLnqKHkkciWmswiLKUXjAZQ3l457ZUL
I0wxn7uoamtYHICXyGhAqNjSapgoOx7muxKBXBs5QGRnfe1YRdgST+NJHx8gJyvPK1JOxSVr/pj8
7PAdLY1PQriFzXHsY/UD6RYmJMi5u2wyQEn5zVduG/RkbH4DdNIs/a5das8LVT+1YJrBLMy8U6gZ
KS4HEd8uEG2lfGZdyeZs9hgeTTLjFcj01aU3Hj+5UfKc9AkXgI5SQYAMdPlKDHzCJqk9szuyg+fq
+M3EehMAMZICn6XRNWAFM7NTXZcgM6ZDJuzi9kccHKC7h7DuEYCRVQ88P2s6Vz1w1G/zXJ3hthWB
zYdwmIWO3cmu7bkyoC6pIq1gLQJZsyl/sefy8GorMUxigD0g2HJR8n3LZMmiRUPJOt++X1A11Frb
E8D1mxDkYm09nbKw3114VawGN2faNQoxPWt/VPQyItFCcrJ+N8Ulc6ZgmfLsa21J4phwconv4UMm
rU42V8PRBHYsD/220D/mCBfo7gOLNbblBn7jAaj4ewp9yBxvzfs+0YJAB2v6F1hBxlhK4v99MP6N
WbCMAp1wm5UPEHcFA3a+kH08zX5PIuKgmRLUWFAfX3tV8g+XI9pXQ6GzeP0PBZrtnC3+vGqs6EJ7
0AjPGlfh7qRgnrzgUa4aVPeQ/43/XzQb3KOPCVo8pmtT6rzebweIrgx8MX/C+JS5mmC+dIn/A4TA
Fsr+4Aas9JIwmdg3UqkWhTjk+MCI59f91hYJR/CDWqDYxZnh2BIFGhEk3Luyh8cb1SIk7aYmtFy4
H+jFrXEmQBRNrkI28YT2H0EjcNqmBP+9CwgADgi9f5BtlXm+f5PV2p1yDKYetXkezmv0KXuSNBeT
ccwQtgxRKOCFGGLL3dMWXEo7IVnNbjQgRiZq+YucIDX5aq1tym9th4z3iI3sL8NhobpD1lVKagtB
Q+0j/2rfEwS48Q9FAFxTh3wa4VM9Ke9oRKBCwLOuL00714SjwzHUxB2hdPacm7NsShyoNKR41ZuN
mNfk3vzlX3MRJYXF2rpknKf7aMLqBntnx57c3cS+ZjgFTKdYK5XKreJUruntM5QR5Ao9ULsPAO6g
spduBrjM+ix7AnMnALxdR0aEluM/t37HDDy4OPtH58ujn7vDnhlzetn7rIHhMil7XaL0HM0ip2Im
KrGD58oZM31xcZaVDp0AGscDo69tZEgS0ekL44ZLWgLteE75dLuQ8CR4rTmuyKizFOeOHMoWxBUB
yIvIuLeO7agWmyjpal0RdU5uepfbBV8+xCONRqus5uJju4M/fmWb5r54RthW2iUJEQ++H8+KCAUG
dGlvxNvSNR90sU2PMcB4WCnkH5ptURC1FsFxLU1ITIaeG3hZYXRwOsR9J/lBySkxcRphd6ruWxyd
il8JcG/LX/fIt9WFKiURCcPtQI0XE2e+h0+/fCTrwR+Xl3fjmP3liF0KnHQDzYxxxu/cw9KMGFeG
JYinfAaCakSEcR7o3/9m6vjwpfSyMV9t2r50Ili3Pr4UVKlDMf8CH5bRfpcizzj1W+PyU0hBonHx
hwa33AY8Db7XhcvVE5mWakQWxaxXmGkRp/bXJaXPkBvT8aufI82oT1+m23ECk62BG2BfaCxJwl8Z
ZUJN+xS9p0sCPJzMHn1xvR/onlEXE+/wtjbu8byjjQMPsouzhEFsgcxthAkihL+MaALysT/8e8ja
71OabzIEEerOBuUKnSw5wsTd1FoNbVI5n+TN0wn+AIhCCBgoQtGRixEvD1NigS0MUQGk/Hifaw+I
e1U8H1nCh+KGiDG9GXwMtnuPyOvwC/eOonHGXsfA25QfatFtEg36TusnDWZA1W12/AzbYIHVQeqp
gJXd+RYYIrIC7S4WW0AIpieagd0KeYMSuhL1mmXq1EPNsjzLapr8zhHhzEVhqIN64utLYdVmEKLr
Av53AwibTH/kTE2GeQS6C54NltldaHdlMnBECLnxmOjE0gP/5UewGXLZfniegOm+bdfXS385Oj8G
8fAGF04RJp761OwGbcQWNDBoqpcrTFqYlWs9/W2LOURUPrz+cmoQucX17K5BGr0Wj//dB0WGv1zp
3Ca41yxgQrB7bJa1xZVeOOprXjC/FS8XPYRFqffJHvL1OC841Tmu0gLAf/oGnhcAShbqAN/1vC8K
38J6tS60dfYsdxDJvr/97bmSBiEUskYLvHzZHj1lVzXEM0Xc/dcvN5O4tmdF+bbjNudcImBz1gXt
jnVYGZcrVIBUNWThSG4ZcfNKHfCvBze5JrZ8pBmPp/nydB0dr7oGuWibJ+d5mb6CncpZLsSiqurj
/PMS6pnZJ+KJasiTOe7mUS3+9gUQFqIy4NtvbdQJZBzYKUL09V4ZAIyrEibTdzYE0WMWtfoLGshW
60v1R1iKQv0UOx4g3oCn5FECu5bCp+7Kur3SjzktYqAtnykZXO345x215GoD7HQvDRSQ8zRlOBYC
buOfXMj+0asIoejizZMtIpVnXAEwt4hvud/yK43BI8ok9u59St0uvP6ehQni6c6U1ss7ZqticCef
R1Vz6clvAD1Ygscr+EkHaOVS9dilb/Aj2icrRIqPaUKsbTe4bLmuhymXpil4suDUoZgFGVc4Vsun
cI+vP76ANW0meWxs64yaQMQjGGXvzkORNffX/p9KI8RlahH5vmovTsMjcVYk63BucuuIdwbm2O+X
fvw/F8trBxR2n6qOtvrUhOmdtSrkwu4T2hgsaE8Qq7FqIEEnrNc9LgpRuPGp1HE/x6KhoS7J75iw
zrdV+oWA3SCvQFqfoBU7LgwuzyemPE+djvPc+/wZCP8ig5jTiqK9lI+IoS2Y2tp9MjNDU452Cpis
kHKVsTkWDGmxU5NjNH7e6J9q4FqMUpq4WNo7hX2PSk8FgJAsO/8tIh2f6iZZRHq3Yp0IkvmGelwV
t/3ZkaSVRoxJaNnL+p4W41xL1OvK/6xSJq6l35OAdmEmo50evLOvMN+scy40AmHIx4knBb9ILmhR
Ak7+VBeHdeNff0EE3SHCx6kqGljHtnyHV3/IHRi4V1IP7OzdIPVenZ9MvJt8SIMQ9kfZNd1F6Nv3
xIq/WLLUUTmsqasFusXmrY2cBx6SkskF6lQdj9mUk6MwAWdO+lrpcpnWObmYJRYXG+AyijP3pNET
gZHOSHTWuhUSCD3V31uHaPwous7rc0cgS904VlAFOrrQWrYaxCF5MNuQgMFDJkfInS5B3fKPhTLf
WmkYOmpZzogmZfl3W4A6zKW94cYIpAcFZgMVVnNK44FcYOWm+q+sJalciJjHsudb9fbDTdfP/25m
Piuay6GFeuP7fJeBCCL/x04qyU+6DbyF+99KtTYOQdqYge/4EyzvtEmYfjriJCsN8jdXT5r43O7Q
3St2ZrtyqdNb3PkxVhYfVPAi+dCD+0kURXm+icng4KetETZ9Zf3c0pGhChmAa9qb4anlZIKlUcpn
Uecdrj2LLhq3FfZNj3siwzxjnw+j1WiWu7U3dZCy7msJ1Vr42HHiRqy0QN5Q1R5jniaaOtGez6cI
qVcl/ZJUGJtDShqTdO5oG7ZuH8mpWKK6985DZf+C3fQdedLckstV+Dil4TRdCi+ZiUok1UVNp6Z9
Te3G7vg9VmhEFgZ4OACLw23lj78uUiqluFdVpYwXVEIU4SlZ2EuKuvD17xTfRBgdNKRSZjEwzSBn
7gFaeCsVdyl0be2JLN+Jgl8b4J5i0EHg82JsX+EVHMul3zZ60f078rq6H3wYyI8M/SlDUXbcMGKe
shYtjY8d6S+AtUs2oqsYg3P4pPQ2dfEe9xWMaVh6oG53Hp95HJckflhlJuujJqXIGSnCJhh4oN0Z
BzRQxYhuicBea5LChQTlOUDfklqqid4zHhAbgfUJRFjfod2gfyy3/MQgsYM9HDX4DiDNuWHAHfGo
AsDcXmxnaDZ+C0o3jv8hQOeY+YXikZWpjvbu7wO+S/iUwLKD3iCd+Pd+Rs2Uxiwtl4F4yYsX1t+D
GGTqm+432kTkJQLeLjnodj0Jl4CuEFnIRbwUBMKlZQJ5rQ4KoBKDEROl1G4AyVY44PSF5BnWxMdq
LiLWY6Xp5BV5Kh4wHKYIptn3FEpOWGAZAMjBjKFB3oOOiAYOHhBNbHZ05Q5aw9wyC8iiBb/rLQsh
480yuTpOA1uZHPB9xJUR0ZR1EikpSlfKoGs9ZkGaedjCqCjDWfyH9XKdmkAoWOk7sqcAyFDUbz4K
xGW3EHQp4hKqUCaST0Rr8OHlyre50V+Zw6Iz6D3nN1wwlmwB6BeouI9r+lh2oQDu4eAg7LG0gjbx
XzwwA/7HCSGHfPs1OI26zuogR4aa+4a8rz5z/lQ6ZmyVzzBZ2sQi7ZP1Yc8MjioWoCEGdl3Smhrb
OmhpMFYUqE9X41Zz7JS0HI+w0LbcxInwmsj4yDQE2GM3+Kd1txlsEmAiLGAaaz2CHM4bMT5dqUvo
cWzMF1mdULVGPDolsI6DDlFfoZ0OiJ7ygqNgrnNbOyuInwaPnAT+ef1cx5/QjS2LNQUFYd4SjXr+
rTyehiDnIyQbxmvFyR2rhS23v09FJBgjXPQZilrpRpuEH81+/Pc0l8u/pszG4bAibQn2eswQD9Lm
tAehTOJBUMxmP8RAULoY9cvBCdwfOE8WMzWnLkmX3kdvR5eNFeZf55ephuK91uKSbQGjy7n4Yub8
gwtwPMRdwekUpCVmZlrNzThyXcDh+cL7hqMFlh2lD+huFgv2l86M09leCjzgajOwMIf+SNWcpaIz
fPURel6jCPV01eGbAptS7MteRCmB+ddlnLiHM6cEVf70Oem/1qg0soRaAWqr4y5R4wfDih3H7wTg
6EucVaaFkcRGzWcg6dHlmtm5y7EQE6jk8xSb6GOCKTU2F5qZpRLtASqmSEW9cSSL7ybErQhhZx+x
8AJc0ZTcJVAmFO8Aj0mdIZI9n6GxCwvYtR0aj5wOKm1HC0Zgnrtbx3bOhx/uunkE+gacHhh1SABb
+HxM9QOhnWXWjgz/jwALIODqtswf/nEjA9eEBVvb/YqsrRZCZKcIR2HQNo8/LyF++OhLoE68uf0H
KZWz2k4klJnh1YhMPIXwtYeBnWvfPnFplBR+/dTYzYEPDcEp0nuA3rIua2lK5Sy7FvL2kY5eSrMq
cdG4nRh8Ar7RZc2Z6pmqZ8c8fvt4wUi77p3YRWECRmLhDyodo/ZnYERjwaFE9Z9THFvjeCQ7DR0/
LPx9Xg0kDBebLNsbF2BPxcVEMlrDaUNm2HYSTS7ultvwPE7pj1GInED2XiLq0ZDSMdr2R1pAVStj
LTMo/SkNzaL0opiu9xmaJw4WyhEYH1C+eCHPkjp5LZ/sw9awNRXBuVGM91rbrVuAR4EPGz0QzOTG
wHsJUDg6v/7MdHRpcVt5gJtCmiXey3VCWLmMpBASz+4ItZSNnNMR9OAq8RbOvahBiAqTbHOwJDvl
ivy/NQ3neDoWIC9ZZKfob0yc2x9DqWlOzlMIHBvwfnOPBfbI+AKO1h0aOWZKPw7lH5zKgHQKSngi
s7STFF5BvNMif4k6RxFGVdqdTxoGWsAu91c7YYvHfZSmDQhNSS70sGhuIdJbDp/038bdsS7/jVj2
9sEQJcxQJXsXn5+G8/Z/ydgQATFPDmonRXZFETahmkaAx8weR9eHKlAfsBMPFK6WPorFlCRcqVYf
Oda38nBMHVglHz/A2QZwGaJLUJlVA9iNLjAf3GPMRQIxaErAsW+zVVsIDVFr7v2/I9Qxn45wkoyf
ll2KGaDT1pPtoJvpCr35r4GgZ9qntXmCX6Q+qQovwGyvcJdxRweeiPgjSVPqz3qABKDB3Bv1pMlK
a1kpekDMOPrUxKbBRY4qgwZLWUhd24sbrycCjikFz++UBbkZLh/EoJuoih9Q6yLZPl3ATKozRyZK
pVoGj4+B3NmI4y83Pk63GH+m7PP8xX8gDOuszEJoe7XeetUDkuYgTbJBu8lm1MqWDvqZA3RG30YH
jevDJ9gm8Z35rITN+ck0GgFdUPzP+OvrVxi4rmXhj1Fuji6xegSd6fkek7Yf5aPVN3qYFSYp839l
RVkIZ1sF6zefAiMVFOk1fG6M6f9SpmvLLJ/TRSKHQEuS6JioZcJgVKVrHupfRlHbxo2nzHAx9ElI
njpDmWf/SsTrHoasb1RVh0jsexdWdCjUtAtKa2LBw0cDSnkCZ6HR9NNsW5LtSVN6F35abwMT1SDR
rbTON39JgkfMiIrK0J30wsWjSUlRG88NEY4Con4T+jmpkAV5lgBuFmwFAfhyL/qWHtVFL/q3qKDu
MxXMOWjEdmhB8o8rg7JrSuANSecKOCAkUO06tYphg1hZzuTGY0ew3ep7C0YES/vGEI8if+8G+nAN
+ReZTnznBvnooZa9LU6lDzVNQFAjWafxdTgnaXwlLQcBqH7jlkts2MPDVq7P9W/sf8f8+t9BtNv4
rwlWKOXtmvBkvrs8AbPrA8JKDi5BPKx5v1QAs14wR6fmnQ/vxdJIXHKcarErHgA4ym0pB8gNwlVW
PXWS9TWT/0Hcy3a1xmQywgzahGXRxTLEwttZui/s7PncCzXL4hrouwddL53NjOW6tAYVG9MKJumu
vqYiwmbZHexI9U+JecPcA9ug+gsdOlLXH3j5ZTtRYSB0aQ5IcotJozcRVN/2yb2UzqQS/lY7ZVZR
xby6gddK1/QBcxZ+xX8jEsx571XBzNz9wFDFv0JICFVdCTO46PP/lwSo+/VsPmuBWNvwNAw6JtAO
VoQPF9rKoPlwi+oSG/UVBnRLzcFhNnJreaG0Y4V0hO7KfFxLL2ZeoE0htZj+i4DThSqUmG5v4mlB
1mnsWSz3uF12k5QX6JjrcNiUzLkgpqDjbHmQMaoIN3jK8jdM1H8UuhoxRJdXtFgM5LUBxkVY+9Q7
jRSmSM2mCKe3lnB4zC95vD4zWgdOSzWbUUoTOEXYn5Ses0q57H8sIlg4zNvuzyJkrNrRdggvhAOF
y9ptqw7fsaw+ZB3oAu8UXW3TEq63bOYwmN9a9ChDTXxdVnubXJzXl2JXNXN8P8FMZNbn+9xm097k
RNj2gbSLBkmmiWLId0Fc3WPtwDdFC5nrMwLCGKLCDvwVKGuGyklAOjmu5bD5mctaz5RxXFbGS1a8
5V16NISdQHnLYDTFeh66Lm/VNXjwDPGpbxnXAOqMvisn1B72LRCdVxV+K/HVmWXci0Ol9ogBRtMf
HL4kB642incz9FrMgiCDNNCEdq4Vq0RGcpUpu8fxi9XkT9+4BFwp1xHHAQEZeJZMQWfQfDehZECb
yqwhbzql66N/KDD27QDlw04Hv9WabwxSYSOxqDGpCRBPcdE+4i3kV7svipkevr/g50Rj+GJlzjd2
DU8iyoLsk6sZG+Ze56uXr5QYC/hY9f1QxNDniB83V883iK9k8CcYibvHoSMUhYS6u9G/OcDdIpBl
Netx2dWIKXUCf20YZRMj4onZ38HP0Ob00l9iHgEmOxyXD6+8jk122uuS6BCo6ouPDQ+89il/SjtS
bD4tbD3iyjSh+SrrP7yhHMOuwURUrRrW1A/wdeeiOr2PHJhMbs3bFRvGs3Y6pxHSaLzwIRYY+Zx1
KCwlzuzVEUsQiKowNtSFvpMm/UEJHv8hSL6aJ9TMWXWqhZ7H0TMYL2VUkpe0LhxQ0D2EROKXYj37
3Yb+Stp2OKcmmmMk+ZovvdgmPdDmPi/lzATebzOLtcTMjr2FuV54Lx6lByAO4P4xXTZrFR/qgUdU
GwW13FFBWKF0i7SmHLq9QH+9XUWpLP1Evfn6Jt6qcIkvwItSFOVxNKukwiWkKbaGRb6DjAUgkFgP
bfCGs3p28Pv8KVnbykX1O7sjp5z9dG9bc9abaaezSw2UxN46gf5NEbWb6OGZmzkKILCBhQ2gOzOg
kqKLu8HP2rVmihIevXODKmoK83qfuje6MXZKX7PEnXaFz0lg1uycgH9r6lsrpA6J8Fe4uwa77I1k
uRFbW9ku7Q4jnywFbDetI60d7cF6DVaWd9HSW/ncU/hElVWq2j1lCYs1VFAfRvHK7piMBqcwJA3U
ZLfD7cf+eGuoq+mxYJqFZVpCiPhQN51ItdLLPt27zM7806f+/zoyIvAzEIlqS4jakbolMX3S1aqm
z1F/rz08Ui7yWhve1eZoMRe5kOOdVOLqlMAeT1DTLlDsJr1T5mNOh97gR6H8qVmiwqrfiBNZDWYo
3mhCSSG0vL3hdx4eRE7QvY9n7L58T9FZoKmfg56yrcIP5iN3Rm1JzpkCqtlPVHVGw/Efr1Gv4LzM
yAxQvoovbvFYLHkPlGic86ACiBKr4uHM2J1lmL86dlnox817swMwjVtRWQLhwZQis6Y4hwio+Z3K
41qaRBPvy9NcH7CRJSjHuIkQ/S928YyaZnfddBjDT6HxjRyG53hXdPoan/WZ14RDjXtSJWPFE33M
Za0jN1qxWV9XZaMamVwvrsPL3dARe7qpQXHgu0uurYiC2t0IyZSjsMZxLjCYswkGsSN6CxfKaRCl
qm9v2GCbqahZcJ+3mAjMrk5wbylIap1mnVX9ERKQpiZpxsOVqd7GNdt7iPNdAaPkQg5v2vjLZ72B
WIqYtjZ2ryL6hJsXt50mzpcK1cvC8TRAQbWZW+AscMBeVIzJSayyIRo32Jbu7+Ym4GpyVMra0SQr
y63fE7bsJw00XnaHSoj5FdVcKngGVhORQEGkaQgieKIVGrzM4xgHPO2H8FjqMUFbdyYMydDom67R
whBTS9mTigVpPzy3Jq3nlU6sdTfeQTG1ZSBugT94BX/505kVd2TGqg1IhhhWsJn6fASBDCne2jmd
rJkwH6CdL7b8GjQCpqT7+4kzRKTSMS1bwRUGBFjlKv62LH2/lV+QBxnJllJeuOt9SfDh8P1Iw0wc
qJH2Ji88xdI1jaiUCxMzCoZXZzJ2cDfWcDqHlqhixldtaPzQPK6X8s0T7bK12DDS1wifT9mcVdEz
kfxU8Jx33it9HY6hk96zIjFl+U+SLGYn6QuTb8QB734BtKLfjl1ryAfpV5nrAzwcWQE5tRJbmkDf
z18WWK8sGHDKrishK1F3TZhI4hxJthJJnsgNV3wl6C7AcFfB/rCUw5oDy0feDzx8sYGDcxxr3ZD7
57KUcKFUNO7Xe5HS1IuIfDavX9kwBm5zdmLSv9f65FQHkVgIAY37I8XuUZUcaHYs2M0dvtvkMxQ5
LKoTh3bUnzXdwkEBxxiPwxWRbZHaEpkdXUyRUJ70YIhdQWNKE6zyUNCCgQEVKZSoMs4DpGnpGcJY
XHYp8xfOdthrW1p9She+dDXJ5RSTJi8kI+m+9cns7pA4gG4bcLQ7ZvQkd2vVpsMsOWVVZjw515+5
LfXpb0gTuLq8Q9JrnabfdE8WMAVqz5q/GnqrD7h8or7xUSL1GnTJq3KK9b+rcl09aqvMyp9s0/8L
dHUJkq+vh9gK6FiO7YriKV2C7rKLfuf4puWNdX6sEhDuNoRobJbFm5BEqy5lFrY/ZjYo0pQdRq3a
1MRaWOF4IKhWGSaZxuPVGJ1YRj2chmyi/WYXAcOpK6SsiKV8cueN6IH+OwvThXqfx/en4hEjtdfN
nB827c2yQeqdQQNiRv2Uo7owhP2WQcEE32lG4B8mMpgYBxWwoz6qwK+24xtDavp/7QWMFSQQa2KE
4gU0aiBPwzJEclbArBw1M5X5vOsBKehn0xzVhiy7c6OU2rBYgZ7EkEZcZYHNduR4yfrcNqC++Gzz
iMr9ty8J8Z0O3+Ao5bxzc5EwtaHTx2Pa0y+hoExherx+rk88l94rr9vAevN5aZLT5aKUHEJ7D32s
FUEmpvx3Vc25vYsShmYOrccxiuZ+3WJzWnNkw4AYvr2y6kuyZKbL7XeRdFw0xtXM8jbsBO46FCbb
rKNws9R6OB4x1C6We4i9q6BwC68Bb0BLRaeGpF5RJxl4vSJTtVjO/OdsJbd5LsSNmHrIPSxKp0Dq
hLLzIwpcGCjuJvLlgt796COgGRJZrq67vyjJIV95UidCDpg8S07wpl0SpYBTKKU4FZxqJ4bd/nfX
y+mEcreJAqheLidWno5qGfYV0rV4kwlIRK0NbQUX0N+qBvOw/juLf46t/0kv99sqJl7v0FFRR1k4
WZSuF79QREhBtMPSFPThtQw5GQnybbpdd/zrZqCKgLnfTCAyf/w3lfITSQYiyr+EzjX51qtVtnVU
PodzC/mWDm1f2iVbnBSr0h6CdmUQZYjOfc6NAJbS3axkZ0Z/hYOAPXiWTqAHSF+r8Q+OtCdU2qTm
n8xUKnUPvUJbu7zELY5RcvU7jUWgjRMFnzmSc79k5dNVCSFSj/znqDgjV5jt1jNJW6amFkO8OiGJ
QyLTp4f7pkMV8lDAU+s6PII886IMOqK2SyjwfsdR59IaZNV7KOjNhVZsnv+jtAcmnyFVhmoSafbV
l2f52lZx0RFij/F6KDLqf4jalWzqdExufvY6PGln8yoeCQSxCrX2H7qR4CI5LENLWWxMvbUJH1lP
QEjjHkvQYJXOSem08/ko3oZ8poA0M0p4gngqWYm3u3Un9eoR/jKG8DH48PM2BpdXIqbhxsxumaw3
Xi6ONGuLldZ7GKylMK0X0sSz/1vXakDRi4EcjUN1/8VofIxEdfM+69fPhAfhTRf3pzCqns3OuBfi
9YtcSaSly3KQ1VyQFi/q0iEBVX3/0iM8is0lF1inj0PMsjekilFjmIOFnxuUc62aitrdeTHvnuGX
RyiDZCjQNgeg8Oe6yQk7kkjwAFgmznkoDrZJ5TQA1kH9RPPTxs4VL6o2J5nSqySii/fkO1jpY/Ld
fkEZMWC51zb/w9IJeI7SWtbGTT1Btxjhic3Jbl7G7DUwwtlJYZxGvZKBEBzdDTnpktMnfhZFybTx
BdUWGehMxusivZhAhZgqtYemazvjtZicqzrMiY8+T9dZcF8CE2+UTqR2ZvVhH45c/qcmj6yoxp2J
JVkp4anri0ZL52cHfC62KyVmzG1q4wThiW5Ms39mB/6wpJMSbvPCi7lFnFEZO1PdToYJOa/1wlNH
2zx70/WrHDroLpYBtk0HhF7YP3HDxMlnvczjvdU9orm/Y5gJFiPiTClYYDVB7OKOJopzI/F1AVHa
Ah0jgbBOPHfuqviSMuaj48eC+JCyPmJVW7wHD6AVi8hDcM6V4zsM6+nebv21TQ82YELcTxwJlwl+
Am6teCHSbk49lWKpVmwXa88zcjUoIjkgSwnUEpsa/IvE0c2o1kObvHTEy4N+sv50cLLlb3ZZZOn+
fC2q0ir8x9C8b/vU+ily6NkTSc6G6ghEmbaSVsp7dyhmOFvsg2x232yJVX3Z1uiztWMjbYkokNxs
0UERuEmsGM30e7+GUlncQ95J2Mw1OqL78fEkGJKO/NEhzoHw1UmlwgdohDh1uSXik0FB1GF2b7In
3358STYe5OjAs0JJDfEXwSd+FankpvL7l2e0n1gMOUutI4/Te2h9ugWpJACF9TxqCGPBpwJoE9pS
xlt5tUl9qPWhr5vSpRC3fOKWOFR0G+Y6gag4TbKHktVta+U9ZYxga/JuUafxpxjVT5xyCFHiUey9
JkmfG8a+DSy2xK+QKHJMGUaCUALnP0ZlqVtU0d+LQ0ah4EDN+wNOqnwxtrmdMPSf4/+mXaVzaHrh
cFSn93X+KIwU2IOes/0RXyhGKpP87HGAYd4uAMQVbgp6B6LxirOKoCGF3N3dlFKNVZZsvnF1rIT/
jfHKLPFx3tSArRfa7gPMg08z7VjD+FRmGgGyPqon5O27M1xzXV1CJ86fDiczhFZ4rrytZa+bzpwq
STGxApnsCzi3lv0YGPRQuWTck9DzIrZZnXPCqUBSp0E/C71vDfhwgaSZKV0XfB+N9DEU/HDu/HUc
IDCPeoGDO8jNptxd9GI9Fe4YqwQPbhdB/4SobeVwJBePPed9DNbSs/yqGlHFjBWvqwtiG8IATpP2
5DDp2l47z9kk0kryOz4DigmZNTpRvbF70wVQqWwuOgfcMxR1sOXplIgq6r4IlE+edbxfnrbg6Lpd
p4rHXvo75/8jDy1mUvYHetiH1F86fAj6TGQzgyC9VV8uDmgyHMWRu9Sb0Yw8CPN8TweyehDjH38e
a9MaQsAWGtuFxsh85w/HbGZf88IVEWDPbSXryrCWmuGQZfrJ5i/fC2XC5KjMDrEsSBRrmZKBnuyR
yG2JO1IodkZibJ9B1RKfcO8nFiINNKkhGy6o0DnJGxOFr67B/VMxIh5EjVfrUpjof2S3NqPMQexw
p4COeQOlWD+4LP5lFPkbLiqaHaGPXyg3khlibqQDvgLJ3tzEZrsVd7dCefTTe3gq/+oYs8J8FFTe
amIOLctb2MWnyB+tVohVShV3ceqN10cKc2rHxlhAwV6jyuIm6O9TJJmTHTw4uEiqrrF6GfM1GMSh
l5kZ3I1kBB6WfQTam+i2hWB/P/J6Q/C2TVVV+Uw4kfUiNWU5ZI1lu3Svbld30coKah01lRPu/wS2
W7srKnASmtGsexmTaJp0q6BmYsd8yxxxusWJiktPsVVz7Hb+71VvhJu7j6p+VLfM5gragd0Ot3nb
n0CvTCSlxDv4AC8UC/kOBiaSmWtRtLQxdSIE+UqNJBuW/xODEtnBd9g2csLuAyQ9YvgEkRReaWAv
po47aYn/PqJKXVclkqn0l/Z3NbB39LKyTbvZUfWK2jUclH3nrmKL8tFSD/lIsynaHMkz40tJRm7B
/3p4khn+BbAsEW8P/SP0TXPcR16pqgyOALIZcNuVQMad4Em04Uq11ZdnKWaXSiHmbyrTikAopYr6
qtddErQb7jjJNoJCkxyMV60NGCjZj8+oY2HGWvPpMWLlSrFC1I88Tf7nLybEufK7NtswFU0b+UR3
YiJH2VAvDCj70a7BOkXbtvcDbR4EFsk1zw6GqT6AGAvYcJyRefBHsBisoyIqexPqm2FTJ44aRfDJ
xvXKLiY0iReRYHxVHG5n/NuL9QdA8DaRIDmSA1/DkyjX7x+QbcgwmGgJ8u0F7XwTV/SkQ1LNd6e6
OhEGJVNGxeIQmv8WaicxMK44lMFxyWnybCGrHfC9cYI5dLD/YHg2A0FgJofrqFCIqt/YV3yHEIhU
YsMjulws5QS7uQuVzxaA7Ry5C+DAbmf9rquB5M+Iljuzbnrorb0eDIo9OGMYEWhm8a7wPDA8QzVb
CNTAoP/fNXFEyOh+zreueLSjjjd2NV61Vd/dQWQYkq3dPWCutEhFYxKJ2ZXSkZzJYnu3ONxe8EQJ
OeKr1EjvOsXTFcOeQNjs09G62p/rbU+ALGtmcVqPszXZpl05m9nzJDRl3r+VAQ2YfbhQCbWWkXJ6
antCohYK13RmbKub0Nek1Ozx9uKrpu4D9ZSVErSLlCcakIXl95CSkL6Th4g9qGzUkTDFI+4ubf+d
+sIkOqJkJbYc1+eE1nfY3DMjY9srI1jFYLEp3MmYzUJhqgR9XMXRb2EYHZbbC7M2MS+v7c2kmU0C
R8SPSqYtC6WLK4oS0ypX9Vin7dbpU9Kh+hjqMB1UUuilQQbXa8nWGLuWimz3NoyFP1sI4DVjQTxu
OOX+Y+6CRjG+D+AzqlfGEdFzR507pzgPBiBGKCeRoee2v7KvB5/VHGyuSbuRRUxRYZUqLF1hJylA
CLe4y9lJdYOS4NOBYPFRcHNln+0pfOaYXs0VKnWpCHhlV8w3mUicGFFy9d8gz83pQuAXu8Dn4gXv
b+MOjOUqT4YGOnN+Oah7ewDvJUVFkdsekyp1gcrjPRbdfLrMxprkutSwWDZC4u1y29oo/FVmFO3+
+5FIeip/P+O2KPfzWGbr3KNrsukZYG7/lZ6RNfO0kcO8XtjatN5lqXWo6bf4Rp9cAKsUkMmT3oqH
M6dk+lYqAC03/fC2Y3BWb9vmsmQz3s0ocm9ZrIG3GMx5yscEIO/d5G2CxcLGz7imF3ykGVbdpyte
aQuaBX9c8z+WEGwLgOxwPGjJvAenYSZAl9z9W6FRJ19/5Fx0VxfKGI60HgaXuFyM3qAkImO/BRkj
BzeDQob65uWGuAAC76Oh9uXB8LqpUbkE7NFWzGaVZd64A4Ee65tqrFqZeWE73aNsORSpSGupb1xS
MKtMLJnziEkeu03rd4OgJMLHtUvpymdAA25mtN9aIFvrVfP+EBPPpdRwfwJ/glhRYSvW/82IFHt1
qX30Nn6SvTOuhZAkMsc7QCjKQiIZRluv/3b9oSlmTg68eJAL4jnHobwrnv7b+sufF2O/LT+jFJ+J
A+bNMcHt4zX/KIUNafGY7Vy5U56QCbW8tKzitr+eAfjVXUkVGn/0ugmmSKxwKizOzOA3zipCAjTi
NmhV57cKhEE1QXUCrGbuS7qXaCpVy5RxjrcXEqvLq0Vuq3wGzwsVH06ivnyPGQzx7f1zxbpeg2Xp
fnYAGCjpjDyzbW+7Qk1Y1hKrfIzGntd6YoyreRCtcYJUPLn0pOLX50n6Ox7Mxsqay+KfjMV+hMes
VRipZQaNKMz/2eUnQwnNDRGQGsMitO7881kMmnLkZQvQcrHg0V/bdsv64b3TBwwzXwQRgiTqUeaq
cnsURzlLslHobgmqxBR/DzqcZ8jX3kjUIrPt4yre5eBnU1JTn9M2NnXTUFRORSo/Ts/FIJay05TJ
Fgct+11rljqNhfPugASOAkTx0B+BhDNN3V+QD1jNNArGJaLhi2ir8WJHlozHf9BBha7/NXgybq+I
Pa1GTeTfmHzLRgi25OO3Xo97YL86H4WIkN8UOWsJ2OfrTHtFuvtZmy0mLOMhJBV1/cjudaC7kved
X9HNuSb7YbUJCSZuIzG38TT9X3TT3CrJOVY2M3DLESsV6yQfdjUl3wCRMqbBYl6UwF5Ic4VEdaWr
Oe4VpyYoZGcPnoOw/7v3HNpyyznAuySR2EkjPJZ/nUFl4Ol8WaMnOKy5TYyzXPF01T+uy0aEL2Vg
HJwiRJfzYcOefCkhLO6XAvnXZdzRWXHN5ZgPKq9JtW6/onDng/QOey/CN4uL3jl96zCVgpst9Wgg
btmAZrX5Hyhk5BcuML6wEsuMRgWnfQNVxJZ6f9RVAYinz4j7B3yRPMPO3hefSBQO3pdI5K1+mF8P
j7JXIEDnYBwKvzqikqzsQz3NeZXN34bmjECYfLEkYhIH2CzuPMKSLmozVZl7R+M3DTmp5t9LhuGT
uP6SZiiOafeGkMw9gDzWuOC1QzrEIaqURGIZ6/nRwuvv0Ef34J00I+/K2tiCejWfpaudPk1odIiI
viv6nkU+twEdIlG5P2kvUcMXSwKjOwnC2M/QeZkt9HTtJZhZU1aghNwYdG2b3SkR0QraMyLeJuyb
sl3GknTpvw9nZujm5MdHVa/bcBwNzBQrOuDIRg4D8P1ZFNtorJPGeD2rH0io2dGlp9NDOUpocY08
DtoZlr5HoN3iAAfO/x/JckDpyHezLIXUvxcvio7WdG4+Jnq7ShaliGxWZjcNFfeerBk8HE/uIgoE
MMUXCOfbt4um3FLCwq8Hegs878ZbXHidJq4zpYmqesMbo2nZICdadI87omYqf14pNT5/8Elm6CFX
ryoXUVSKROQScnZPwqUC4oQhfxIJVSFqiJp1Mk0zOEklr8dNhD/1TH3nE1rwDfw3Hl7VwggT9UDC
iUeZ1X00nMYToqDl8J08Z4jSmnA4vNUrhizkeKeRQPgtBn4WeGsNEYGSu5VO7XkZa3cE+KZ1ss5E
6RGSkbIrHM4DsUDAPcdxJMZULQnfg1zaKFf5KdwzusrwBf8eNIiYJ6aChQHe2z881kqy5Dh3bJ9B
sz9Eg4xGaBuXCjPhdVhzQbxMZ9YG84bVr4gTxR4a1ihp50zrO7BNKic4KZo0VAoFb1kHbIwnRpOG
uG/o+ikSww1nF5Q/EGicFE0l89psyeQ6Y2H9rh8Z7+PnMdFPGWBkVoTR2Kg1vDvUWI5HN1Vo5BLD
cRO3tWX5MIZimhoipLWP2xOSDKaWo4aAtvr6Dr3ayM0Sz04Nc7kE3SKYt0ZM8SLzkg+Q07rDwN4N
AOjpDGMTFeQYYD+smmPkJNJmpTCKFU8hunVoH3pH1kkWoGqujjeZSrdm5sOjEf2SehmKMGCht9Wg
3MsOEokmoARLCHhD8AkLduo0Tu9wrrBZZSeYAnlL3FNZH13opXpJYKdxaNm+lfrbaDaDp6TGYSnd
FBNvcB42lRQHuSrH+d4C9zGhPxQQiUts91y+PP1/QrmsdVSYQOPpKdVhJK0LWNOAHIi1xXtAMAVc
ES/CJrHTMjCiTlS++K2VkrkHOH/PTh+N+iNkWAq/XWfDcG/uOpx9W4P/b4NMPN6yOurCnFZEP5WF
7Wl3vjy4WrrfhuNRT72sOfCCrkF1lapTcabFpFFRDk6zSu1kP1ULG/DoDajyUc+ie88Y8Z5p4rVK
oReQ3UM/qgQ8qosfMK5M+BH6rIURYWeIlPAv4u4hPPqmQv6HlaghkKPXlpkIVUKVrrSEEl/3Unxb
DB53M5ibdWFs9i03fM9cTgE880B+hpY5cvE9WagWioA7+STWfPr8hnpt/naH2sUjDikJ3jbE+KKk
FAzjAxsLZmMPWXACyluqorCyRSt7B/Zw6mKvdtzMCWA2edxoYngwv9MxjB4fTI7TGMXmltHbxJcY
dUDyV0AL+z5GrWaqmWR3NsZ3FwRQvllxyOJxP3lGXMtbBagpslBFSgoO2n/xmqoQ4jIjEDr5MMZZ
ekso0ezQNGGsMUkCMEogZoTjc7DIqptUfhEA0FFtarAICzusKalpNq5rNwr6e3Q1NP+pjDKc9HvB
0A5Sx/9QRcmXL6fBriLMUou3bpqBljdMSfo3h0etQxyFODLVPhIFoaT/qc03gUmxjCBMJ96NzzWG
oTQoWGQV1EoX3fUJI0v4PA5F13dzHcHKDzzuscjJgysq5sUhLH/059Y7cYi6wd6RFo9Pds4ljTWh
5jH71aSZIt9h3F9XShpSU3U1aHx7ZHEm7bbLBU0ecUDYqyymUR7pGWOpM7DWoVtmyT3BPyanpzHT
XriN0uZezyaTxkSXtBt1qu/KhAgqshiwqIOiO4uQ+I8c3Lk3duL1oRvbaNxAFuu3cfhfmh4LioaA
jVscbhpPAh5hkot0UaUGZFHijUMh/4iEIlyCzMnfx4QiGeW+c/yPw0vylFGizLydbM9K0QfMWsAL
tvRA2Z/tDwYzdjZd8Bk14zx+TS23xnZ7OsfrYmYBjW/DCIJ7mkPtkSFaRI4rCTCzsED1sS/6ZzCQ
v6BVVQJn87V/C3Bg1Sg1iksEbf6ZrRbAxSGXARVt1oJO016E0ewoUoIY5RS0/zAL5Y1OYnCB8JX6
j3UXpXQWn1Lo6VZh/4Uui4Aup7F9uUGfjeoe9YH3UEkgcqh0D0FTACsBCcSPd7kQGGmKCJsTiwfI
pmZeffGRd656KXOl92r7kOH9f3/u66afQBcjXExkhKXIvxDzUa6Mvp5hgGkq9/XG/gP2EysZhiZa
frkP12qPjk0Uz3Mz5J04Z1BZFqsFAt0AFYa5jBHCtFBgS+YDdtqH5GihtoMKS36MRwP8tcxorer/
mkvvGECjBCxSWpzt4V4hxEl2NkO3N+yPttYengbdGTkjkjxMyZ4snCtNDMbX6ZHGzLvbH5I/6QAS
uvuM7f07YVtwn1KUpxBD/a7QzMQSOHj6neWUOnvcg6PGatVHaHvDj/D45MeOjUE429a8Eg9UugHm
BAqMeq7Cg41qSPkdNT5GQdSXvo4DPmOFfS3XpsUIp0zHMCLvLbj5G24PORF8j+uXwfvDA4iPC7jg
ADWiHC9r7BqimxiNMcRy988G6YYUT6OA81Di+1lIrGYNZ/BPIu31zH1B39zQp7w0HST38R4p7nKW
5GIsyZzfMeKrumKUUaG/RpO2TbIfitVe1seEs4td8B+nVlor2CHXMAIHLoqtUMOkpx5c7uqhhA7c
s5l+C7AE9Txct1jnfZHKl8/+mbt0sswWUmgAadpi8Oc6rL1gX3/LM/kLvqVkbdJ7hLS4hvFU+Oyq
w9YQuoU8XRWZUrJQAMADGxcXxcD4ZkwvYPFvTX2vFWuIIJxwv6zeYmyZOCChQFBeN1wqXqvVKchA
DQ2Hw8/1uhUvR4HpEK72W4ufD1F7N12kIaZvgpc42VsohU3/r6op571SzUreLLsZSc2mTxC3DA8Z
YOtP35sN4lrOJtG0SBjvTEG9oYkAnCG6RdtCEQKxNMKiIEPZWkSsQ1czKj1eNwgR3QfFy5DCDOQH
C6JxSwdNeHFBmisPc51+dRAH69lqdKC4D8EKDs3yfg9QI7V2+0IZA9jLdyeC92w0WTKK9Z8xv9xu
TsvpkHvICx2F1PHTQ5dU5ee0816FHa+bWjTDJURzlZe0wb8rMcNgAhqldFzauWBGB/26MtxyOuDD
461Cuvg+nTGp534kIqLzr8j0spZKx6o/iRrezkd3lSN437fL/C4nrMfJUggM3SKrQ4/BNGcDkyDu
tLq8E2eXNvNSfCvlwAcXxb3xHsnJ8ioIbT8hlAqmW1dkxT+Pm9G29DW2+9TtXzcUo1zlUo3lo3Gd
vTiMtt/LLVno8a3dmYoM6u3TJ8d0arZxcvEoksUwVhvGFvYnmbLZfjmuJJ3th1J3xa4Ln3/lisTg
tKCyUP1v8+PeslAjxRBsTzG7RnF9m4f8EnNtgrnGqsF5Vsu+zvOuO4hRpTR/5graW6Iey6M9bvXu
2DfieSJwkbRSzhYXSRbUAsoI01N5Udn+MCprPwZGNyZ5nXHoA30Co1DgRGjFalhUxEsM3HcSsiDN
JwMbtmMdpRT7IQTutHTSnVqxztxk79ouz0D/yHF5uNn6HsVz6ufco6QtTP3zjVWchbksr/T3PFOd
X7CvGqnio07wDZ9MXonCAiEFiQYSZsHhf0utczkzXoH9DwjWdvIpsha7NlthflCo05rgRR1a0uzq
HkAXeW1tBNwlMJTeS6mLMSrvvmjCOeFVP0d+ekqPvArnS8RRT+1wjJuJIziEyQ/65S5Nj8z8xaLH
zl4VKWkX2P7uefpCvENJufFHKeibkuAvwb5yiVyN/+Uer8fQNBa4q7iqgoQxDoE6KiZXE3jrNzQK
ONDS8WeWNHC6vDRlXWRa1KarJO1LnqwaxSIUqVMkBi86DaK25aVmMZZAvLiRkukjAFktLqNlk6rG
jI4i7gt+TnF/XUBXddpcAGecYmCXWD8YwgEoKGq/6pRqIXCi/jaLj/JBXU72YYaGgAf5rjcZx6r9
gXgZgSp92InlEcUT+iQJTlCTDY6lFW7oW/tNOj0RIMKYmH+V1qnsS3qVSe2mRC7eEsdeetNMLEr0
3Y1yU3/qO1iYtfIRtcSfOgPeB99bLoxl8oVWBFkM3GPMH7M6a3f2p3/cjHkOVxbn//yKGpSQhQ/Q
mzYU6YIC9aYpekh8NGrv/OWyw/pUXes6PTQv/KmDWCPv2NoClLCGOGo6ccigY9z6SijsPw/677Ke
SigT8rN5JjkWfVv7r6sEMR6bbyTXT6nJxlsLt/8xTaLJJv+vV7yNR7zzzmrrqQgtxD+uVPS8mpBo
WOLXjAFMCq2CIx1SWXz53dRiJ/dUj+TbmygjV4bZ4sYvzhFiJb4DWajznAqAhu0tTXNnwT2mesBk
rxZohiUKB2ZnjCxfkr0VWeY+qUpiVhfbozy2SLmmOLKXMPTZUBSZBdBEma4IY8c5ZVUvMFWaCRVl
S++pRHRXbxZn4pck/uyI/E39uNJB6Fe4IbllNFATxmg9WXJx4lY/t1sKyDds8kqwuTkUezKrIE/L
X8Pny3+zO/Un2n4TrysMeFVAK1RDub/puySYt+9le/6GrqwubrKGpC2cIkrB/mp0sNFwc9svD57b
/qAQzkhAt/M7HrxrS71c8UGXwa/Aj5Rcil4kKAhvH2p/3FG0n0k8bAVGjynJrKid0iLrvaix2ztG
40eipwfmm/9HrFuGrnXVnnJNRm4l0YX5VQOCkUCzauKzBISjWpfKoOwAa0i4Ga5NzGmyeShqkyMm
rtJWlOnc0q4mhaNAN6CpH0OoSoqQ2Y8FGyGcXwTI/EE4fWx5NX856Wpc+A7j0mftpqleTUMP54PT
05/E5BiyeStHg0lEDknLaveNbFNWNHzYqS9SiyeTRBIdqQS+yRwMKOPJZDG7heUY4jq1smS3p+hA
ttTCEQ9cRJVe6JuZbiq7V1nss9V0nl/d6vkwvT6uqCBZJq6VARxvGaFvxA+seRy2/8lnYslVCB0X
r7SkkJydNa8UTYqVO8YY/10UOWLWae02ZMx2oc9VstE9+8jcnACf9iMz1JMh3w92cgB1fvqZZmzg
98KwlY3JownxkBOFanR5TGG5slYyh2MNVAp6IUsx7LOOI7Yi5bP2BBgFFQtvcLaiZzUog+qzGhCe
nNBoGyvqXMC/o5f4UMt+eYvegu35bynKUH2ivYDcjh4fOlL+v65UfTeccW1rixDEV3OZYwuzdQgK
rbtEdLt/SBGlkRHH0P8KBlnmz6ScIiZnpOt2HZj1tobAwnm0ac88dCGqdmJnC2+74zYtW/5K9zzO
bp+rBmORUscNnKppFtvDnOhkXtHgUghIGDpMwvAg/y8Q1ghxdv3ucpQB2mh59YRo7NBchx93N8Eb
rNHZU4CbKoJSGCidxs1Z70iKWqXgtkbc/GAceLjIp9hkET4ykSLNe+oDAMJsho8mKPg8MG1YuDSB
8CMurFnzDzQlX/+hobp5qGRT3s2vgIPAzoHwTjfX5doJIvVZ5QdeZVZJ/RIOXg1eCgvXcnkCW7S3
SQS3VlFh9hEaUpRuIykKqOiiokrSEjwTcme8rPtk1jK0oLsLpvTmvy00/f2EuI7qxjTO1tL1SgIt
6WWujLe0n3+NU6ucsflq1GUjVdVYo1MIDDD5bqmdCUwPTi2xFJjXCW2am2qn/fj/pAuI5HSmWURf
R3LjMJ6iHoL70T3q3UtyBoI3telFsPmhaLIuz93IB4eR1VJQXueTnNLRDYMs5tLD6HvtiJosFXNO
ao7vMmVtBAN54S+IxN4NXTzuwxJLze/ZhkAk79rjoCx0H+m/C0kmuF26StX33whrE9AKYLv2CACz
Y3AeF8xjZxJJDylLbguOeFpjjH061H2cuTAO6SikmGoXl86oWd7qHHCMFkryBDJ7Qj2md1qHp3OJ
/mvtfjk2RJJphp/9tSZbvx98Y1a5VpiBJo3lIG3ESBmE2Szl/sUPw9ZAvMrbmd2C3S2QdBHUwdft
Y+vo7+W4DIO24RV5BcZbWi0sdfxy/7S/dywGmDygTFG2pUhDkctoI7vMpJXoUocAg/hlnMxyJRQX
6PbKLSLa5nmJOlHpBrTikv/jTs0v7KkGTFnWOOAaB3YP7w7UFRlkaFeBqbN5UJEi4yDXBqB6b3B5
biZ05LUY4JaJUeSHmIRJq/NDIOIJfxX5znl3YdtwcLGbFrzr92EgL0aBJ/nNvPr3FvX00WblH7gH
MJdvjLGrQym6KyJjyji9xD6uaFd2RMeo8c7ulaHeWt8jPXjgMTGlk/BxPpW22OFpS354jqCHDBfR
fwcdwxpP/uuzXneHZVCPA1ElTT1U4UHWWpm/mVsPmOyHGicI8XdkgbZ2c7zavSFZU5cpwbc09zyW
WEZQc26Ggb2GFDQHx3We65QL2g2TxiiIUomtm0cFRxjcOy4F7YAIR40eHDXV26BPukcykkbz9StK
Gy466n3rek5BV6Wke1jnyHzi8NBvMDeGLSXl+I64J3owzzstlHp+aoMCDxcpjvAWJES9eSOUD1Ox
tjzNa/QZEaIx4K3SCvsZIWvFSW6Vu0RGWkZWEirNi8wCQMFFE+zUUqSmulIK43kEw9Z5DFRV7GxM
ydKE1OjQiMT4IluSHF79OvfWEGPz+5a9yxiNX/fwAz2OlFZ41lhR8vUAxvevazxjNP9SmqNBPNG2
yH4VfRpoGYLtmUZVYxpMYnsSbU3pF8BS7uVp91kxkrYOB/1M8B4vbetJWcjDr6KOWu7NoAvEuTjD
LgnY5+NWHdZW32JuHsXSqNcHn4Zmf1NTL6MSFotJsN9mFJTJm9N6FaLWfSEKblPgKeg44hB/czDn
BJHFGh+YBvrJJL21Dv5/AAfbQ8a2kbQH+eEDJ/zww6lZ+4kjHDf/7aqFnc0TrRXee8QL9qNItJ6Z
6O0696/KOJJPPdKhGc+H9NQxeSRL5mh+9mtiKvHwugG7eIwU9jpXdsv2ABnFyxdgwH6VRtBemgHf
F/B/LHnmblasx0PGCefp5ZPF62PLenOfK0BeoNbdSWqpIStrYtDsNOg6nFnNXdmBKgiK3HJeyPwB
Ga7458UoAnCdCeufjIGXR51MIwQ9ZAxGAqhvxpQh0UQa6XUbOXNImqjAvEd5aB+9yzQJFgywQmdQ
Zr1gTkazYeddIpHqlv9SIy9NkaMrKXUZCcuOtfve8XaSjd7cv/IY6GBq+GRha4ylrN39mBZwMoc7
Pj4wtRDpOOSJj8XCClBd5imDoyTw4oxmi5nCYdilA+r4qnA3goCvg6EeuQ4S44SO7U/F5bL5J7+7
ZaKnnL7n2Azib0ud3GYYwCqGa4YBFr98VnUTrtWbDD0Vf5xmJS0cLGJbD7bDcVFNcoCa1TNtGGTE
3WIMr7mf07dFZptRU4SPNTVXsa7euqYjrNOTtPQ0R6z/KtWXqT3/hJeAo2s2J5XZ2jfJv3Q3+o2i
W01I6HrNWyDFekUrgDCrRw4aQnQL76GgNax4q9T3dDCzR+AJ0pQzq9EB+rWM7E5KL0QcdbQKX7bx
fuMkKZmmc+HDn865kjtkz3rku0W7qT6OJ/Lj+kMBwqYm78EatjoMsL8UKrvE8v9TXDdelvSZP1pp
a2AOwU7oE89Zbl6ynJ2Zpe2Sk5m0Hge9tjbyPp8C/7XNxJigPfHLot/3zeSLa1MqLVmMIAV9xIF3
wmK0cxk8EbMUMaZt5swh5HixY6ltfMtEvJyjs+KmUFVB/sP60Ju2qYXRKbMuii6eAEgKTAiT+4sv
CnaZk3Y5gUh3ZW+VbDMRI8NAbmrkV6Y0FYl+nc6kHjngnm3gJjHCLPDWyNRt+vy6HJVyJVc3kcti
swuo46zRybtNp/E/7E5MnoeN5rVUD+kvLwt3lDztX+tb7VR8DD08bWEr46/kct+VN4PDAVEDlmUr
Q8oWqYDx22rdhscvA/TmSEvhE3fD49figJLhXcxHxF5Lgx7Z+vjxGM0hyoeC8UxJJqKErIR04Jpy
AHm6NtLbSA2F8iNeV90hNi46ruOc9zIax7LfAIpIMqHr2nb9opOqX9JKnG6hC5IhSfGe/uvsudqE
exW2IDNBYbpvSxKE38uF1SkTWuZunfeNySxGt1q9TdTys8NbZghsJEWy+y/j7n9mKhJ/5uJPtOhT
d72AUTjTRa5LjHE+RgQF8DgGI5fZ+qIKMYVmiGPCe7OjGIn3wTIb4D8nL4rhgWk72/Tt7E0nttZJ
O3+FyvfRAIeWTsvnchLHzb1SCreo0ZkpdB2AW8S67XO96G3S1n5G9M7ImmkkTTDXtTGkWXruYj36
U8aQh7AEvokbnhvCHodaFoN8gh5jscsrRLvcS9VS4mctXWOr5PLYzS/OQn9CSiDKOmswDs4Ji5oQ
OIO9fbCzU1uUTgV9n3ldlJM17akKrEWeDm2zinQVruaVPawnBPV7wh+jfLavFPQuVr7YojNxHMn0
JSyVzZrZB1A5rf3axM1y7f2bQVv7Bb1SzrTNJJ11YpK94sFoi+/nQ9wc9Y2nsHQi+9oaGl5CNDR0
KP7sKx8Gxc05WQ07TSOfgq6imVv4WzLqnxpltmd/ddzrFe4dzG3YPIdt2ZnWaBDgBCe9GS1KOWOE
DTpRjGJqPjzDNhSRMAy7t1hJm7nYXoY2irDDbjj6j4kNGWeXCxxHDTy6etLuSSSV/46H/wKH/6KW
n6Hd9rYk/+9mlZCx8mlQir9jjVSVIJP4GEzwyAZSXz3wHIS2wng/+XcoiSxAtgUF809rpol5P0ya
JPZ4fKOOZa8x//7+xE7igwybieXOK448s0+iSw9AsVrZB3rrLmMb0MjgWGsp8NevD+r6FevHiCFw
4G0j4z7KoWFukv55g4T+hHBIsJhBiMJXSzHq3hhUU4EP8RTfy8Idc27fgD+qTIJtJHNyjCp6iusn
9QdytHzi3fAjdyEeXwRiAOvP2Oo/7itAghOQBusFtKqN5/k8BMFHiE/vfxuU8OP6YfpwTT0oU/Wx
7LYqOPYEW6IVrejcbojriO+DN0wAqf23YG7EHzksRsjM+A8fIhqWzMahiJvH/mWlEcA6ReMNEhB8
ooTmwa1SInsMpSO/3KYiKETk8U+snHzJnt0gikFE+VLn9SXSkMrZY/GkzAN6/JCEPigGtGY5dfS9
LM/BIVHAJgNuXld3uoV67BC50QSSpUO5BlNLN/yziVoLNkBOhfzsml7BuHYcawbWBdBmZg2GgfA1
LyPCFKCxU5dwVvg8tlkYScdFFTrIwk693zOMWYU+gA8sRSTsoX1LlN62s9cZxVZZQ25kh8KYySP1
a9NfrTEJiLbxI5N8i/JuNNbXv2YdhacwaQqka4YBIIJabu+uwsUhleBewlF9QtrEJQOwZiWyi7k8
YsH16ZMFNYg4bHF3IT3ovquD5Qnj4iZuz1RypR9oZeHXIPOAg410vN2Y1cwWxORwKbzMFNxSpOfZ
81zTbelluI6qjemIuym+/YV7z8XPURIk09kvim6vcOGnIJpO9+ysH9Dynp5/t++nsi46SHWxUdu9
osqKil2b5LMfLF12tLzAmJbBHIZlfUYildd1QZnEbwBgoOLal03luqp02hCK351N/dA22lks9qIt
OhcvgbcMKI92zmALD7aCczYBdSb3gz0khcy6gJZDTJSBN03KpCZMx9FPmGMaOAQvS7VMcN6Anvsz
4ARXfzDlD0CpMm/alkH/pk3CqHRphnSsGfCzvc9633umZrVHXcJ8pnFDSc3uwpqjr1FdqqfdKYpt
tGVa2+xo3qXgS05xQIItFcxn+7xoMhaw0qjIBNnVGxTamT9X5ctU8dqrNvIIkUAvsy/2GIgwL1os
EpZl91q/in5EABKPiViuHY+1y7pRXtdbvBaDNzYe7b4EN7mN1lM7uw5uLV4PPaL3je/s+8Po/IlS
h+vSpoEWjPTmHFG7XVLa4AZx9bbmRJ+9FD2zHWkyrgaHSCRaTEp8aowsLR5EpztvtsV+smsZ2z5l
dlQzwzQTiRerEO4lgqo0JB0Ha9hgqEbnrGIH8YkfsdwAK/A6nfjZRh/D93YiCy182DDj6LuWXdu3
x1EFZ2yvq1pqURLjUH335T+5Plt0zBhix1hGem2miO7e2KUIqdP2xRL15qNCCzW3PEfNy8CyWqfm
wQqKGdP0x60QnlkkGnuAhl7Bd0KjK79HriDVNJbokk/H9acPHb+Wh+Znt4yupPUFJ+B95B7MBHmG
itRGF51BsPuGwhP2CPMxEUORGORttZdFGjxvztDtRAFYxQSSfmkMhQI/AnsJgF8YDrm5bwbLaiz0
QGNhwyRCCYF9lHB5MWjp8jov6MvyJSJOocJqvRW7ifvMNzSrJH0hPnUetJTn2qR2eSoAnhyeva8L
XDalv6KuzJKdqVda+bOgfcblq62+7F6+4/9U4dzkeFA8Durn8qRf/ypSYNxVjb6BHu/aJ9FS6oNn
jLE2JjHW76/tCgnXlChaSgcnHj+tikZSEmcDn4tpaIgbqkwM9gad/nOYBGVpAQ+a4FxcDN+tn92k
TSanbU3bjbrer8ubnsyL6wkYGVvWJJEKbDli7dhyAUR3A9O4nKHx9igd94rl+Om7wePF4ogeTX1T
Pu36GLmkqAd9zvq4MiijOJ7V/nWYnjasgZbL+yokWusexP7phTVjwQYPNfLUAvOHOlifJX0it9+B
KgQn+8E1KcnKNKPaKTkl19d9dDSaaoUU6f0zcOyoPIPqkC2lDGmDBn7YfAFAJJpm7vEvMrZnjtP3
o/c63nNSNsws+VdgEs4wm9j5t8lP/hOtH0+/5O4CNrFBO7cEJYFVo1l9vS4hqgsWSb7Bciuej+RG
S75ApFxHK9S6LtTuUItyChLaMazpUzQyzg1gogE5hH0f64yW8qHEGEYJWUBsuKr+E9gg4evof4yS
+24krv4rhpL47VIMIlNR6iYw1GSstsFhhoVPo6gcbFDmDqYynUrJs1VMQBp37WPc+eFtPawhIWwJ
fkJ8QZuvjaRiA0wgYCWC24SVzzlEplc+eRwjg8uAHx4G5hdxpJbMsUj92bl6Uq02yh22bLxAELfa
YjXWsEs+oE10r5+uNAW5ii8E0voDPevmqt/idKliEupXbD3OcZIr1K082rKN0EUH2x7ElHBSWuxD
Ks/qqxcHRsgGTvvsXPyE44ZbqUZMXtAOAKSaHfYGOiV6mqOLtgQGXtpI22Hkj1w+fOe97jYl5j/F
rnW2/TO/A1A9/CkRgSNBAy/QSxCiBepc+t0UIryWA2NlMDtUExjZHqPj5ALSY3qVWALiyx5tYQAk
FCZV6Jw+2AWBUQHGRVcXfWmaph5a+A/DR8TSxSfO0u4Kac9jRU2Ye80YP7u2/c+c4z7qEuYCjoFR
WbCMQh/UgPJxEW+EejIvt95XAWU8+FmX2e/RjlAurfu5WS5w+1oOYfT271iJEn8QSVjN7usqXhvU
M2JKsTXXVw4MLdjZGtK3w6BDkXcmrsDS+BwvsWJeXJehfMi9Z2i6JC/+jqqhaq4ixPQxcBdLbqn5
ZcOhn4bzOmmXBD+heOFqN+C3ZWwmOo6YUlWpigdx76WzDp0dXss+q4awTF2dFLgw1msLfjaYaZLF
/hQlcKTC9fhn96o3m7YLvKlhRbctbFNX2a6wNMOTcwucbyLLGTTP+CGFQ+1u1J5OHKVeEHTjBzQf
vBkBvfv2Gju+FhOL6vopn7nTL07O8nfEpLGmA3hyycE0IGqhTgPHXwMFIhmP7WsMTc8i3Sio9qbH
g22KaCQQjZBkm1LfPnwI9W3J8Fx92u96pg5m3wDflaMn1BvALKMIE0ScMo9gwhWZLX3BaQzyB2ce
r28CXPlPzjiGzQvjRzzTyjMG/1dCkKUrNACFPRgneD1/WaDCaAi4zHhzxVWKVnjeBjVoGSyUk7r9
gMHYoSO2QFeSH//03Y1cBcXiiS2Bz68U6L8aQzNxI1PJEcpJligfqY0Iy0GpH3VNNfGZUZ1b2cTJ
RO9zCERw9woc4XvzIb0HYhVuSL7dQunzlw3xq5BhmR2P1tEd+/kjrBo3CazfcJQmBIsftBz/ChfD
/ESVbc6MzZtYmbWdUSHu/aF8TAIwgMOrbFQm6YVh3EAHWQi28cSf27YvDDw5MGHjvxZUj9DkNoyp
+FFL0FL5p+JUR1CNJfwgDzc06lLv+6Jt/gG2oPCAf5tpkMV76JZ5+ye7ow8wITHzuClDZIUECgQL
VzhbJgaj0JxY4wLpRV8ZhIJsQJyOsccflDz0kXsnBDbmPC2ZI273qy5eLC1qDfXcPG+4FgMy7YCD
2NjHmK8JKAaoYEG+aWVob1KvP5TmV2ZNn7JNYbo4br553iZkP3pESh+8e+Sx4yZgmwnVk/lkhL99
cZTzrwjhgfzls8gDir3N2mEOMMOnS+BUPfkT1R+Uj6PNqPwF8hiSfnK8LhiSDbAEa5FxFclIWBJE
fNVQHzHzR3/A08GTqj6bUHyoB/jlNzGWw/nGd4+aAmA16ozh9A1AAUAToke1ERr4ios5dvjH37LP
I4D6hQW+qBVBwBn2dCzuyN512evVGIcr4WHpw7+S5zPjxJK1GDcnUxpk6Vanratzi9wOBNbBnvaf
zD8Yo5IN1ur2b1ajjx7TLmEHNBykpS5GCZn876cClZGL/AO7zdwxlWdBIldDKzs6Pta3VIs464R/
91zhPezpcq6jK20SbNAdhMSMB9lVzoqKaEOFJJw8p0+DFPEci+1+d6QblioGkA==
`pragma protect end_protected
