// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
zCCr6W73Gtz0mVW0sBsDauD5Pelkf4H7LmBPTB3kKGybn+Zy4v8HWlSRyo/IElEDha7Eq37M89wJ
18CAgxI9+/3wpfgQ2R8iMykW7sSxvtlhpDavsNQ1lidgVxxRHhXH9BB3tnspH/HvhZ7n+erO58XF
JOMCez9ypikksi8M7G2q1gpqSZpHULINK1d7CYNUNOXv08eMoQbG+Jd2IyxW7Th7SuMEYA/ULAK/
SlRtMeGvTu82mIRdLFMOwJabeDOx6Jujy7ieX53I3nkF0p3YxFlaK7e9UR3EB86r09zwR2J2YT2I
4giZYB4GzAu7m6Gby1e7siomSEyB3dcWRmKnSA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10848)
zI+ht48NQ8zaRatkM3jvsWl5/toxJjsFco2iPE7VrFNkEXq6Sk3HKcWzeGfONkQ4C/zPpvlzsFCw
KkQyuOhYOof/RenOS8sNz/ODJUisIl9tba9w0wTZjhu9VxRBnpWYsbFLpcjxA7FUCtNXYxY2amTc
/cClx0LItYUUWJFCNG0WxPiFvQK5ew5AA4H7MqHMXi7GXnWqd1+u0l6QaU6VJI6s4J1cngATlRua
Qy0yB1NgCFfRDwHfJPmfLHLHUfJihpbZj30KmCL/AQLJlXVrcpqat8ccwMpiW/gvPW8g1qsMOyaX
SlGzeBOb/U5UfMKMjfeqlbTYDR4i8Mhn4ASrDJWvhCHjKUoh8uSbxwBngYoRL07ZIU540dbXpYMN
5IlIxeM388d++9uqtxySQeT6ald4yQAfNocBWfvrRR7i0WoZruYChksn7Qg4oPBpyvhmIG8k0CTw
FdzDhezWwram9kOmXCjc8lXo8PNEx9gz3S5s3zfnHcW/9nlN0hsL5lXADn+XlKXbTEWyz5xRQFeT
hHWEtBByce0pZabqRaTPP6PzE8qnkFxP+pPhYvv3qDZt/JvASSx6uw3xFRykNjkloZYNFmpOfUAQ
nS64CTbubU5ldKfYX/mM10SZ3IeLj+NciF/lR97EGjuARFrR9z6J24lgo5s4vbAjPjgeg7uSoJLX
vmLjb9PQxqOIi5f6scNHxStykCEjWDZya+BD1lwsq744MQ9vmtMSK+Gr+AUe5SxKp5jB1mj9ZkDs
hIWpCT8W0Rzq9AY08wB0aB6DtryYVmmGjbqBwyb3qfshs9aS19bf/3ChqtVtlTLQHMUlFfhuIMzV
nnDn4cX8HKYecPNcW+u1kbDiwreOfOCKjDX4dnIHoLYiGydUyPFnYL8iKeucCDdC0Vitb2UxJzTP
fqy1vlCTMWr6bVJhDYL3NG7BirxjYKRkL1PPcVGimdetdPNpYWP4pdz94QvdISio2hoNiBp55OXT
Hfod3uYSYgpPJ+PovfkAh3y2xRPjcw736T//Tk0RUZjhhykJQ2DZ0IArx9H7cDUz+exBuy6QPZhH
VleqJBfF42yewPa/Z49kZ9lwS+OMjPtoEhKNIIVHXBGLt5vAdH/4Hm7Dne+57D/CpXnrAw8zfrdB
3+IGTERNqxg50FZz1aEKLfvFG907ljL2ATsWR27LBCFt6nP0pnXlWfAMB4OuW0vFfEUBN0ywz9B0
+8NNewDltNfts6WyGREtHFv7HGMbMhU0NtySorNVQq2G1582ADI6mwA4SBNn9wTPlwgO/mTcz9se
iFGVUaitCvCW97g2Furz0wvhCPpVuKxtVyRG02s8dQkkZz1Wc8ZB9Tle/FMIxJ5Hbol7E0VAfENS
GcsxOl2wK0in95vmzSaBDXgIrNyYEgjman+tdRv9vc0kj7QP8ZjwYS8NN/dIyG5X8DBsAxuvTRHC
D4fJR4ztgxoxrqp6RhX308gE6wEgrmwgu1qKh4DYXajPo0Ib+O3EF1eymmihQJeJv2jfnGtLtBjR
IQmL4c82fcT2mpVFRNhWIuJNOB0xbTgQ4gl+FMmspXQgBKOUhujMWv2dg8CMiTVGSpibeM7J2UO0
EH7PhmD9T8jVLY4RXLlgfqAfJp0dbeWIRW/qo+R6mMtIfg2BjP2/YDqMB+NIKG37IoeNvrpDxjXj
9niRLA4GrpRHwJC+OII8kAkXDzDoPt0ykdprSw426l761lefy7Y7IPnTJIXAxD7YExFtTN437ED3
OGyun5a3u2/xMlnQIcgS+ydnSxOQvo6JQn6Pzdsx1EoDDnrqZ7Jyh7KHv27XCYnnSM/BbkhrTS1S
VFxm52vlvwMsjBVkugAgcjdDf2wnJnpbyA4Vjg7kl2QNEh7MCDdOK2IGYN5jmIhbokhI4BAUxRq4
G9eklqbrX+6Gmm7R4qdX66MEUvzcJukRznxprCmgkdfo5g0/1ZDK6ZKQGsp8HbCPVpK3z9X++Sp6
HZLfYDxiDPdGk3uQIOxerwem57J7+K4vow1MXkX6gZx6gAMat7X+wppaWxhHJ5fojkb1uO+VnDJu
5ikpxcGL1bNQGQBnfqCFTIMJHAnB9yTEi69li/fkg92gylEuWLDExeW9RGrUKx9Zvq5DhKonQ6dr
Y09NRRfrHFehlsM7wN96D0DWM3vSKVmk/jdVij2Daer7Ds/so6NOP954BqEXGdewEbTsLVEv0371
i1f0j8pEEMJOCoZG2n9TiJsj2vhWD14m7XE4j26MtsjrUE7/aYWhOjGvwiDLaIvpWDOKgvhCNVZA
8sxSJDmoOhRlkBPCgAM/vu3aHDIiFS7EKzfe64w13VK9R8ogR86yb5EPHLFBoI6enCRbQGZ2DVBV
TZ49Ui8H5Yhxq4cdWX0XrklDluh7wqkQFC1hQUXef3gpZqhpfI/HGOiEa7zdRVy4JH6m2E0qh8+n
SyvmUW9WvshCsLZZ+wkSIgHyTqwFN0cHd9QykTYcfazmWtimZnMzq7PrKQL7ypChbMHhhRaBvB+h
Q7uXF8CeIcrEJiQSJ9c5lZetY3lEuWQycXxAooPHgOfUHLIgOe78l844xjaG7/+UxLh0plrMfW4K
yrUSSREaA1A0k4+Hgu3v/lpzip0bfGOITPjLtH3dOLnNSdZyqd0rAqzEKssgnVYKzmJRwivFnQJ4
6u8gZqcrvtsVXAxB290JpJt8eUIvfRKLK2qnedu0iPYmJXC6kmE5HVACxpiJ43oUGogOJ9TAeSP6
PxAtjY+sIclHx1Cy38bHHeQXtWimY6Ez/SJaA3el4j2pN5SagV5Nr/VuyHU8gwA5K5ti48LfBMz8
28uEz+J9XkdHxPdJTGSYawPTPTTw9ecSP7hAIGL1dTfZaFcybSy4U7gX3udUb3sjhcHf2TqdE7R6
dRThFQJ3SpojCxfRDPjfMxY5covBoCoQrf86U6E0a8Oik2YVDZIjx07zbrw5x5VxcK0alCdbnK5U
LbkScB0Nh/JIR7ri/RlcnQIM5HcBl7Awnj/oPUcD1yACPtSCP7IYcdcO2IlULnZaJw68PI88BHea
E+aS3JESQ7g83A2xY8qOwIIIr3gDddRarZQTPds6Lak1BjpIIDEQqTLS7leIsNo4WXFifiS8yXu7
TSTNJ9Teoyxe30ril4GsCDf9MUYyFXZAHuGgp7o4z0WqgOLbQLCz9eDbpyBSUnPxW5PNofo2P2aY
TZG1ZXaErCTyAOanM68k+HUG0x+Q+41KEBF3jg/aqev5IdSUrw7I7Gf8FQy1NBPQyxN6rbQPIoZ9
6vfoMRvLlNPckaqU9ksqR04185zsRJymzx1UdLg9ycK570VyqUouZzYAfkoj5/HzIDXLU2DThi9F
+Pllbb8C9MJ9Tmb0/XccZCGyygViruugFPi9iQa1DtI4AzVP4BJe+HqCDSZmZicckRO/nyhKEH6D
3Hch8cIcZ/sAfei0KA5u9N6W2IC+YU1TceqEkVAq0YMsQRhD40zzfblklicTqUT3METoIO1CDU5v
+AdDf50CafSD/Xfa7LoR+NVHPM5JzWMjf7h6uHQPEmsj5ypVKu9mC0VWgQsDd9dQORXYsbLKh+Yy
n4ITIPlGEQPPNhDqdnxYehczpbtgEppVB/hM0FlbQU34dsUL1JZzpYz8mmWCSyre4W57OxXh/JhL
tW/Kmtiw3WOTW/VVY7WR5Dj6Rr6nCS8BC8GqvFSvndiTJeM8QQkOGBdPAavBnFUnKrgJHV5E3sMC
LVr33DmVzwinPSJY4POduMxrNYlcO2OjhuBlmqLpZ0zF9hKJyHcVgOMPxBFkSodTPIGyAOl4zYEI
6Pkl/lq+zoQ98e3K50FE9bnVZSDQ2aQu5S0A/5+JpUAVaxJssNI3YU0TTD7VkyvQcgXGYw8YBPNv
WlIib9mSOzxV2Zsvnos80w2jlliVzuGpsYZPQ285UbbzDITWtAJQ0quNlgkelffbTFcLM7L1A8iz
tJ8m+D7PCzuLqT6ejP+9yYE+CI+VtJRFgnaq4HmQiK3NJByw6+X9SmDb+cagshWjjXA54sPdDWKh
Ig7hsNgZxQp1lKFrDoXsXVFQ1V5KyhdZPW9nIV9iQE+zp2SwNa8mFwgfRU5xic1IYZvf4y3lDKdE
69mEVZJmh9LWsodDoXKH8GMXYL84rlGR88ZCOXjY+jYh6w03buCZjE3PBtOFI0YWnIbUApnDsRqR
uK/TuHGslWcMyeTCY2LiAzQ7dKhpeKgRVzISrCklSWJ+X8C9OxLVvBN0MgO3hVDivwhxbtJZoCdm
VIku3GLMBNkvWUpnWoWE0A++6fpHfLFx4Oh0VkKxqy2ZmI6VLKjD/cxMl146Po9NvI4ZXUMAIVFj
zlJBGwZDa6KFyCYRCc32e1FnHS82RXvN1o7YZ/pnN7vQniSfQ1lJX0JVhNZmDBQIZOvPsGWJW++0
O+6SpLSzs/o6X7vgM4KJ5oGCZgSyirwPQrzkbINMzX6mWP5iV3ycIGl38nZ9Bo77ZEq4jY88GZLD
p8amWOd+nMGgVaVNRc2ywvzv2p6yX4qY0CHC/90zRzq9gXaNc4A3LLA4xQcPEkKDqMx9Y4G2GVLD
a3IrRfgm6X6i8TO/fgLXT3a5hqCzaLiDuwSrurAZunNqWvJZq7LvrrDg7S5nqezra331VaYRYO8c
AnVPF1fxVDZwScHRNl/8zl+7TSc4UrywF/fhPN1yesU6XswKAHGIeuNYGY/0oBOKG2RtS2zv+T1Y
DIL1ut1dc0YjByBzQVPJFtdKPVHDXG3DDZI7MYAJn6nYS6I7kslpTdeqQ8RJtJXatFcD4m935Az5
N2bxjQPvQ6k2hw4sUU6nEtt/TVBJR4IGpfmUdHcQeQnu5KAkjgEbQvWvuGG1ok6e/iY0xrZlOeFn
aC+1SYlAvT84kW0iXNbDJbnF3A07coEgD8X2gZyw+MCT9IyzgBgTxPdYZ4OdN90iUEV5aFQJgDo1
+/zJ78k77+eg0w7Yz+vUox+uFxiiz2JNzmYPjL7TzIOh4fDOFc0jlPv/oKSikzFSHGamyjZsOm1+
5mGM3Z46JSl1X44I2MGqdw30OalEOFDld6jcymA6c/F0JiYdfpAVUyKJ1BXQZk9F08v1BnlATMRU
lhgRvnu/4eaqByjS5jNcX2ddZrZYSgPngycPaSpsF/A8DXW37oCTdP75tnu5hXXfz80IPERrja4Q
4EBBxJp4CVeep/hjf/HHTpvIQ1akdmh4S5zDOkHv7cMcsACdHfi3QCn+upK3z+HJVRp+XBtaDScd
7SR9/qdvmMbJDDjgxpQLqoiWor4DQd05gv9dtkJHFdHvKnIQq+psLJWwEtJGa9LsX+aUVHcMoVGP
w5kERWTPh5bp+14qAklfF5fgsgnrOzSEIqDbsTWS5nS7cA8NSbv3Ro1joRlerke883p0v4JMvjCg
5xZtNBzug4Zu9/WDiOHg7xeZsMVaX+Y7mJuZckDWYZ7SrBVbquRDIxfnzam8a7ek+lCP8eONdalK
vnILO0S0EJrwa4GfV1YtLxBVcJxHrW4bcgm1UKHu3cyYAmeKkUBeVQSOmLSytFL74ZwcTKmdOuEb
S8278XHIZ1h3ncXa9sm0qUmXgGoqKNV+V3wvWoE4t+1H3aKr1S/nUbydiJTb1AfoUMukucRoc47S
OTbeTuTAbwZDgj6cd4B8D7tnL0c2bL6O9KUsRXuYf/kMlC5rB6ezgxom5gpuGs/PaFeP2mN3Uir4
ZE4UNU5q5J7KLKIfZQMfWT5mLZYZgFTiAJoC2m3P9xNVmC9HhHiJFQHvOw5nWhUATxWfi9CgFI37
JbnlWzKlcBoTADJ8dGqYWSFOKBJ0aeH3rm/uLKXXlBFCE83lfNfCgHnZX+dPErC1XzM9D6F9MtqU
87UTcVi7x5ryJdzevKFxkBbB77QzaMJLF0SAM142hxzJ0C0Zna/1UxXinBdUPOLYzujCZpWAiKPY
CAFp0K2OPy7/e12K+YliKRvFTD8CRcmmTwv6NJ3Qs3nlQwv7AtiPveWRx91v9XBzFXq8h7XI87Ef
mDUx/IqOWQZeNrpdTvi/12XR55YLoJOCdhM5NIMj3FvXU1MaygEsAGP/zLdx3TE3l5B+1B/Pq6SC
NguXB3sWgTCWoDPIp/FO6bDky73Z21C3tu1Yv7BW8Xz7IiFwJLrQ0Bx1bC4hh7Mp5Y1jW9Oz5I1Q
F6H95NH0zGhaaFZ4HDbplGvCR0gp2bYPN17fJzdn3ShO5cfx7XujYC/1Rx5vFR3wimz2GR/EdKhK
BbmKTXAfKbK4Rq8UoRvi6grNJIHqORR+JVMRwOMTSE5lE/YdP2kqeIQ8wHtOJK+ep+dIHgttHfcP
7XEu9BbzEb2IoUBOg3ZoVQ2t1CBRvmY1FqGoFzEQ9eVVo6OYnD68jb1A0DQgJhGhddGW+zcgipjH
pMdq1CvFiGiRgl1NT8Qx7KxT5oGQIDZEdLZ6GGYmEpQE/rh1waMyhFGvltRtgb0gi+wGIWHdFvaP
DTVyuFMkLPORvZC0w51a6kqWbP05PqQz2VTKML7BR9/38glWUPZ0bpecDB4QMIx5gbW4+etvpNvl
WzEDCPqlzs+PIJ5QX7PbFd6OfwrGS0fC90eCu5rOb2bbA6bE9XO1Nk8DrgkBH6CWVP11mZlvDZv9
lCL6OjZOasImCqQp6G4qa024wEGhJo2Wk6yQQgPW4+vb166Z6BxOh2vflGDkyCy8toi9khjPpoC5
PpFnlN2QX3OwYgjRwva0ahwwWuJBUeH0GOTgjqSA7nWqT3Gd5qd5nKc1d+IRr8Y0LIZih3KzYone
vGcSEN2+4aU+CfeXApXU/kd3bqCCz0opLpo+MkKIsiV0mpmOF9IcHoJlVdDJ2AoGynDO8AX42Fdh
WDIH41Huk0uXRpA3DJGX4ZaU+V2FYw1dXNi3cmculQLfmdzkr4BCVq4ns80DL7BuUXLpEiaCIycZ
jK3pygRVvhFsIq5A8HTV47JH567OeZg/3Jc7Dh21jTUaI3eKxLo7jiPTRUUndWn1SVrCTP+WnsQ+
cP5nDQnsYPADBDNRjp3kkMAzePjYUJmV2ExwtN475BILLPEe5mPAEQe4rM/SLu9E2IefH8ssyUFO
aA7FLKOvmP7yhAgi8hXj5ErA10JkzD0Ryml/K0mBeBhw5cIu0P5v+2SmurxwU5BkEIFpldEqglXY
Zc7sNRGu5sV9uM9bMHGtPYUKVdjrL0oZX9Np3xgvlQdMWA+bvImbEwdpEFghZonZ/iVIwy2I8EuG
8FqV9N6SIQliT8/HGxNcDv75+9YZx29B7mZ2pT0RgsJ4Ck3ykf8owg770VZwYnj8PcVexV/wp6o+
j+HoSO2U8JT9y/jbwHczw6padWcc00gZfQkXZJt+dbph1ZmdBBcODZlLHoSP/MKTAKGZpEfOfwwg
Q9pAV5D1GK/T+teTjocbDcOGkqkl2BIDk3VV1SaZAAYYm9SKYxSNOZQDrSI7wyjSZOxVMQNkeOkI
fGR0Ed96okeBuSRZPP0zqziCgbBpr+xITO6xyj8eM0+yHTZsNMhUkDXe5i4i5mTTC3gHKlTDzi9d
W065HNua5dL1KlZSS+hya9A9PwQRme5B5PHG6i7gT03/s3kzhMCnXt1xg7vYXTqUcnRshaz7czDx
+aewtJFtn6FVBoFC5ODe67gh1zmjEhOoTwVJQMHVULmr1bUuYkNIH86bpIHEq+VwV26nVCOnT0rG
fNrnX5m91v07sBeTgyXlRTJV+RTh/ikxBADR62qANu9dYWkUnSUkKa1+ROA1GTLreaVF78+NvvKj
ElwCMVb0NQGufWN8Z3+QBk3AKCjf5HfRPd2YEapC2R230qoxmR8mc36qi8LBJFpV+kout3f1AjIE
DvTOGUirDUs01atGbaZdJxCFt6KIJCuBEMvoBO6/5hxC5Deu+lf6AKp0qyI9tG0Yo9w7U/ZUD9gT
VU5zNMhwGCHXcf6gVsPVcY1imbGczDrjH0n7IYUrSmwFtgeH6FeqfYBy2yeDPvLJS4eNqBsAMPxd
+Vg4AhfckVwi6X4BgmZqISeezT6822qQhQryAb3+XcX1cKL46Fq/w0cwaD699P73hch7A1UMdZkq
WsyI9yAm/iLRayTVdXVFGDrFkPUtuXKe5HTxW8NtM/0RiU2EFLHVtLAEZeJB8SIpTpS1a9UhDedU
b65Pv16myk5/gFn8VPIG3XdSob/eH514rWNT0lZ48Mg6O1vWcVBLPyWaxkrYPp/R7AhVq78ddrUK
6RrO/gRmf5gfYdOKn7OA8vg0+Up5iwpyovJV3HxMIKaxjRzil71VYCsljb0891G3McNXfILbZE+J
IVdFMt6PQff9VQFMQfRqLcyLAZcT+NUo31TXmlkqpsmSz/EJt7zxFGjCRGD2rf9TifWag/frp569
w3WBejcoB0AHgdmdp5mepft51k2hOmENHdANylx05+51GuYqSVk6/519srknqXx0afHiecgHQSzo
DEMjflvU2pvUdjpsx7YVn7JlJ3lol5+nMpXJjh9eep30GXWP2it4282Mcy5s5T3llDGbyIDBtuEL
CUIRR83xYQ1hNcIoCA5EJY1diAXyORCLqN4rrvmcH1h23rktiGRIlDVRN4BejKMugwhocpBxMeJg
XPJW1RF2AGPj2C/99apJ6cgsHhsN8CXMHV/xzPFG9FoKCIFX7nv66MM1HhzE/IX35zN34g4e3BMw
V22pMa+xknJ40v9Z2QfvFz2oSsAsb1k5RtdMVHxz6vsxL/67JbmvjP/R8ix7abJ+ZHsjBOwb+i/7
+oippvadJjOdl+D4Qsm2TPF7eFSr702E2P1r8eBC1CbiscO0DEdWrS/owd6om+PFaMzdgSSCOPyM
kZtNJIm1Z27BEnl+bioQ9haz9ipvJ2vFIAON8Z6WaUgTFF4phpUdXPypVBLWI6xI7Be29lFdp4vR
zW2aEOx41Li3DIe6T5qzt6CYlA5aG5nlN+sE1ckpcCSFnW6jDEqU/62mRxnsQiwcld5IiIfhWPqm
NSTW7iu0UK0ugnCkWZOxVfzPju2igGYmVWUZbRmwf9E+zKaUTr9kSMyeUFkd81k/rLB3VOiw7IFQ
MLvKGghiDIo0/v6MTDrwta5SQpAAHJWtFLv86Wn0PS3CP6TpckP/m/ZpnQl7JStjALPvTfYM6CGJ
dP8c6Z+C9cjBs1w0XpqxCzEgRnAyekss66wVN3/dwedjRRb7//q1ZE67C7axAtVKXuO4IyytWQJG
hbaUChRb5/rdx2rogaXIywRReXwlXJKhU1NRbvYprGiRcBjS/NusOYa8AM0gy5F2gqXErkFCV20K
pcZzdguKfET8GhpFaac6hUi5uMqaw8KCDu4HheDI8aj2GA8YkEr3KAEsiS25o/3bU8lKRgI4lcQz
CTeyI+7c0aCJqBUaGBOD3W+6Afa0oRGERfXSf1uzYOgMwswOlLoBn4TL9NlXgxZ5EmG0cEhVp3Cz
hDjmRCeiR3B5ZPUHxAiEF3HY+EHEbHHGk/c++q862BcQVaEOr2lHEOZ4O+5colJW1BXIqjUZuHC+
m76EYzR5AgiROXBtQbKvGXmY5qRfth6sjRPlGEScNb0DR+qUoel10jicIPdyutXYv/VSry9c5wvF
OtEN4tHlPsdrMQXywUqhlWxp9yzujiKzd0z5485A7MUauGM5fRo5FX9MoDXzowdHdlIunLp9zlWQ
1YNRpz2McW1H+fSaEqLhcwxRtEZygBs6MWQnF/5KrUjjkdkNFoni17zjKrT3a0BmD1La9zagG9r/
ARWDFZpKMMp+0/SLE82qK7NahuwHC8eR35zhs9Ml4d3QVJEJe/Mj3+znL1Ia5cWJdMKWiZrfG1s/
zuN+gUkyd/neNL9AiSxW7Dfs4tILqRwJ/cMmM0pdH37KysEhh/4WMITLs67PRRyulvB95UHgXVCU
5oTrWX/V6pIOfVSLP+JsOBOgZS2sdJh4ZRrxRu5buBzGj06qLNQ4EwfuENLBIUh0VoTLMUJjVAAB
zO/jtn/C915Tg/iCi0+tXGmNpjVBv91zju/a6PfyJ5doxOOPRp71xKDjbIqz4Nw1zYtTZ4e8zRJj
PlxxDpaBjkpeQpvUiozXUbzHdXdDATIansGz55U/W7TYyiN2RGg55UMLihFEOwLXuGKWz1atfpRX
bh/hGABzB6SOt8DeFlsoHqap8/y8K/lkdvpgup5VLrio0HhK00sP4A7XRLMk7eRrYXn14HwKQTGe
0L6WMr280REaJeZb446K5BAwEsDIUwljyX3YEFbNt2bfSt/EGo17Fo8obF+ICqI/V3dQrvXIILry
YtXcgDlh9f63V+Lius9CvgSarSu0S+LMkDFaJ6LfmsqMenCaMF9yPBxh9HLChGzt/0HwkfNNT3+5
qBw4dUcr3gNS828kviWtUFU1MYhKdjMr3BvVXN9bI3BI8YdJMvpLh/blzJk/Rf82ZgRQ73Rc/NLi
zfH4BIFpoqB0V7SVLPY2HbttE6K+qN/b99RrA7oZtkPKN9HlOyRNJsj+RWD2qmbQpthoNvPsyGCC
drpoJgs40j/5Sfjyi39M4hfhrr8dfKUZwxETGCYW5zoG+5nP5zcX4fVzHTV36Am+lvTxsg8gDH/k
17mZqcvNEE5ITiMJEmDfHq667sT0OMzywPNPSdBIG8cxfFDzBzhC1fIFGQOv1fp/J2dGOoltc+3g
5v1sFW43O9y4ta/XV/k3nQm/DT9OA5+7g3fxgghl1EAgzdN02f7Dv6OCSu/olaN6a7+BGpejBWwZ
L+dwrzzKs2k7GPvvw2W+tqfyDRhGAqRvtEJ/j7lG0fiRHVU97VtoYNN+pRiXcwpJgoE5elGNFPjb
SjSitLSO347XtXlpJWAfuPA4sEzVzkX7k7idaUMHJTLszPSTg0ziq1mfcnuM3Zks/jqIQmG+WRGh
V2g6cLLgRx9pZGwnkpOz3n8YpPIA6dMgIf3CjhCqxduXMb2pL3Tk41qumREc15ewxLtPXlwDFHjN
VHjphV9wJ4Pnpez3vsIwCbUMWafV6VgQ4fo+h1Sm0bdRWZ0MBG6Lvx+XgF6uyzGc9WGGMB4I32xW
Dsagf/4h9dqyrh/sOrtbO48KnrpWns8to87up3+lhlJWnGmaRatrOUaSIoDr64+XVrFhVYoTY6aS
bs9TRa1vTS0/Z6I4FslktwiQALR7RSZQSJdIkRjmERAaJ/sRZs/srX0+2CT0AXxrUOgMb0mkzgNt
OBw4A0/Y+B6OzdFwf+I0iDPhwU4uGrhrK6gGb1qRWo2DlRirXidpJILcMfLMEXn4d1wOrV/pnpGT
RbTdVwpfxMuMxvKH8sX7AGlGHpVjDAnuP3Hhmqo4BKOXNxy4Bpwck5GNY2A9q8U+rJzo3n8CAmID
i6QaVL6nVgmtcWPh5GD6DxwN9MSW7/q3lZpM6SRNSvbMSX18F1MfmVmF65RVBHtVmyO9O8TztYhk
x5NGZbRBQFFs0G9/sC0G7Vxw9kGtJFfW6dq49/tiOaSPjsXbp9eGIyeupbEacbrRX2i+lfwKGfGW
d8cdr2xTzADjSluIksYVn5NUDkHNNsuSPX7PDylzHB1RB1fn0hjHK6VZDJ5N4NsHIE6Mgjas1jKv
dAF9QxURYUGa8ED+QruQVFw24yFLvIqSLobIRpJoGGugHGVltko/DwTl5XX9ZXNzZdEB8MKh+oiy
PpQrpHZHO34uw0UDBQpAte5Obuzi+fHI30t0lFCMRlu9ABFqx1NrysrknxuuQgZc+5V9QCQ3C91b
0M7BvRoTcEuuk8dZJhrZ004x82uBiEdp9+0NGioYIws/5kQmB8bww69IAK9cHKEPLeBBESZF1pva
KD38EzxdLhPjjaxnEE3VS0P2KNexmsnXEpAMj1O8/S1yOJSHHSLjT3S0j1vn/lBrs0CJ06nTjN1C
DdqdxT/R0V7/Tos5SPVH+pFN9VGZvzYO9mLJwGw4Bad1K0vCTjlFS/hBS+mP/FfPDHnA51WMYaE5
bhxu1NAHrq8Or6vM6Z17P05t/WV9agfzGAk8ltrCCr+icPJe0Pc8rPVe1S03JNzUKv3e6cu80V7n
x8sMCO/tsoPlr5UCKXyon2ywS7XeJIXzS2VRV3vHWt1flV7ZlgbfkN4kpS07izkeaVfWqlRwkXOY
zM6BAvaL95G8fY966n7+eHksgPtqB85t/ndExa8tDhaeGcm8NLU1fzxPYVVvcXAZyT9pGQ7REgbm
YLSZc0PEUSLGx9tWVD7p+k9Ts5lg6o2ay9nxVqHnqsL8DxLNceu9XS/mNBuyLKQwwtulakvZ29Zs
eacsiD3AM8kbpMu0uoOn/rDPrwbfHUIW8wCp+MFg2rMa8CeIAWfZOEtbmzTFCBq8wGfzz2T7tlwc
wdkcOrunzK4nEb3QGhF2pX+enM/kFiT01Yw7FePEo34dmKOGhwQQqTkawxSL9tifYbwTI8xOlg04
2XAhBeBNN9R7i0RT6dtAl+R+OV37VOGWxLI4Ah4/9L/e34iy5wFAPx0QDGKaIKIzjLqtEGXSLxI+
9oj1jigM41OHtgw8951uMaksJpntlsEGK6ugF1PrZPYyn2/qL311ITq6yYcclpm0HDfe+QWz3Y2C
hjvLB1W5odOoPVb2Z0P/LsfzWYJ8Oi/dy1xwrSoeIUpRz5DaV3f7/9G/YJlmuiKYXXYYw/m0Oc9W
FvT5Fq/56x/LYWsDtRBfCgfnZWdZFQzgHbekEBzf+b58Tdj6iWqpo9aKWaqT7p6QEvJsv603aJIz
ZVSQ6Jw8DDU0B2zMQi8Fpfgoc9q6T8g45O+d7mGlAjR4CJV6odKjmnqDIBHdxqqtHV4m3xjauURd
BuwmX66iOa4v231zrveMsnB1hYOjNsZldp9hkMTOzrroR8eCWFKTf3V0fkb2XO4B25zf3cMCk0pV
Zhbxx6tt648ZADXJrTLLPeBKQcwCP+73Fl6BZDG5SpuZTWibe/urYB37N9vO+9YP/IqLXUJ8OQLp
IK2y7MMZhQZXBvJKXAeWV2/bcJ0pAjzG0XQL/onrnkaEh61PmDi/UOjJzfqBxN0m/wIoN7pqaQt3
BPNlYnbF+HkOGjOVDTIij1jROvejrdovNIKJOHTy7tJJW1q9rCJSzGVic7nAoKtye1tRgmIfpiHY
K7agw0/+3+vm3PqEITkO4FEaRMarunZ3/as9B7nm2YVC4XE474Ks1rZDd54BXvu3RD8uBCSFTUUT
szp8A+9qISvI4+xRfuLZeKGP/VKmaha0j8h1q8a+rEj3U2JGXUGFHU1Cqi3Zx/jiSzhLLxeqW2wN
UzjUOV3KPeaJFtn+DSaLkIn8iXp63U8OBcsmcBtccVpmQosMllreItZxwx1qy+UjCYXBBVYJhJYS
7/Th+TS7JcA05Z+xkYyzDTjFGBZ+fNlglzlfE6e4yX9+9YLVJZ6SdKn5nJJsMgD98UzvsuRXMZCP
JUVk0oUp28UtqoxudBO3tqug52Z41+qafWMM4OVrd8E3KOZqyCJAPWbIGdSywEcaWlhyYYetSWxn
Wru0uQnHnFJnv2IPW6RQE8cbzVv3CiJxE2qVW4rBr+0UgzpalBS6yz9+SiQ2gsMlIuGCqacawylN
mfw1+fFXKzdz3MWQPWVNjZtXDWj3YERNtiEqj/6nu0sQtoqZCq8hmb/O1g/lL4xAt79gGpZMCo2Y
k4JfOtFprY1w7kGtD6EvLqb5WPe93lhPaF19E4uENT2W6NE37GZwqSOklR9zUQNhqHFHoO062IAq
x+9pQLHRyLAntsWMkc7mtx6eac1eNS68K/NXGx/kK7UH8rzGNczHObgw+Bg6Mb81yamaPn017M55
RUG5uOoB0U0HCKftQ6urx4oohfXECxkTYifDMIyuIJXEzrQcaDdsfmRNAGTFjjhnd/koXvFdYW6G
AWkPzpUtNoUjQxzvP4Jxvk6QmuZaxu6h1QStFuWpXqMjk7VJ3IFhhint4xNCJdIpP8uKf09SMTT9
P4zsHiU0i/dG9JUH79fA+S1RFGPP64ozaxNL5+sbSNbOR4UsROHRbjEP5Wmah3pextYzJqpiB181
9tLy3aLWqYHUTTzhT4oqrGouoO868rcZsC1SZube2EVI6VT0xQ6/kNjW4hNOmXSRzj4bjOfM+u2F
nXMzey3/Y9c40mRVm5Q1h1SeKeEIbU2qJqpaQPbXOHjPufTWMHln+x8bzbX1EMgQo13932ZJjoAc
AwG5u8smzxZDPpThwQZFioSQ2l7zbE0E5BfbANuMqJTBBUvt3vTyw/dRwNlfI/RhQT94PPRV8oHS
ijyRkG7B0jn4Wb7wWF2bpbLAQar1qhv4nVYWBicylrFEYKYrOGKttqVJLIfgXz8ME+GycIy4Rei1
Cm5DxFEGKph8CA1QoeRRAOv0rVuPljVcVlq/5oci/Zu84cTsm10zOxgpd/9qqsIb4ROBfsUfbeH0
EK4tEWETcke67KXvwZ86ORadtKuNZ7bjmlCauGYqEICBJeRp3mIye/MY7M1EqCDFu2ytMnvSy4h4
1vmu7XJtmn3VuJRdFRnj4WLy
`pragma protect end_protected
