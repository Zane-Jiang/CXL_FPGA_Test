// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jleUUAfzwuRLluhL7HbhPnx+iki8kArkMtEun2zzSNmdn35O5tVv83FWnF5W
SOEPjxPU/7v776L14rV90hklaQoo+4v0PxzcHd65UAGkcHJY6LPBydQBmi75
8l4XGkjR9oHUcEN1+7sJRa5RglXV0AVHJ+ib3T25P9qN60Luot7/Yjlcy0fY
sFYFkfnDcn/yX0IuNK5cmQ+OABEP3Z/gUv0WFw+cdLVdWoumLP504jPt9Y9r
etnhc2LFTUw1l+weYUnhQ3OTjYMY0HTUPn034HQYbBZ2RXLMVgC3leaifjJE
7YdOk2chV/vDIwmNzh20osQLT7JDOwDantR5LeSwvQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IxhecUvOLwKaOrsy2+wsshRYUwp0VbayOK//hqpCss6oDj+xTCkopn7f9zJ9
akZ/NNGSti6/CDqzLfSshTzTfOOMMm1FHDOne4i4FWZ8hCXw9OpOaVKZnRPu
9iFpDv6URz3oMlsXu2iyFiIS2MirzmeyLvjXJl7ddzpqtQlN4dgTGVZqnzNS
oYuDjLmuLVbWvwEheq40pSD6rd2JGzxQ8d9WZBq4I7GV4f9s1qRbC1veCnzW
y1Q02vtFAwLmtXWu/S5txZYW8wLOCHR3I94NQW90ngZ0zkTe/Wt+kfkiSohX
ruq4P58p3n/2wqLtBjuKDttaYAEhDLGsbg//cdJang==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ByUDNB4AobJLHoBMzXt33cId5w3gtzAHQc/JxFSrIIk+U0dbFurf6EipnqbV
ImKE4pfkp1E35rt2GJPEPE4Qyn9cq4aBKmmsM+QErb+PZGXgDHG0mhUA2qeS
2hByR9XS8m/0CUefUa4UF3+TfC10rbp5MNDBrzWDrMiEJl2qdFePGAkaAHaG
GPfX+Co+rUHVjMrsIPOsHeI+stlPS/iFGcFLGR5Ilw4VSzqsvEQ0Pky6BuUs
rvI0CR5lOv0o1m6DEjm5nQurW4GCgXCHJt/7BfkqxOgyB7broj0PgLu60kBi
ykvvfOnk049r49SRyZ8+cV4gzdZvlF2JpIK7lC4pDw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rvwddKfb3SiJwBK/Il+1nkBuDs8FVI4CivJbUVvWxRox5X0unyRilvhO3l6Y
wVAsYC/mhPEc5JUGeC7CegqXeYIxaqAyaPxqhD8tl84cabEmjgUarPmlqDq2
75EOgnAdaUuJMksaVNfCbfWxxhvEz2oLYPnpUokv8kSzCAZCQO8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
s1KzStwIrXj5DXG4zKd/FdLqRx1COKA2FAXU6gEINJQE28f0BSrSGPc4yYT8
Sk9GpV5kFdlfhoeyc2NbpKbs4O5zfg5y9PgehvXaog3wz/23BsK44oEtY7yX
wGJA4fdlu5qNxz5W8HbJWWYZZt0XC+Mi9bavQqmVo3WC3lP8t0mru2Ar2E8w
OfleDwkqvWAc8p/vSsSEzTUEnsInbiQpWQE7gCqTfU1Eab+36m+di6y3eXuc
FyTZTxcAZgn5oiQBbvDho3dyJSf0GFjRYlBjcbVGkKAfi8xqwbgOtECzLGvU
6TKirlKEOFjS34207mZCT+24nx58RJuJefr6Vdalwngocw8XBESpYOKKzp0g
oKG8nHmnWcexOazY/YdUES5jQBlogR6vG/VfWNfqdTE5Yn0nOG+meS+WXJ0f
FIfZyjXI9Yf4Abj0kOgMWpWg3qyRPVeLcI+5DKHqeiSsm/aUtKHbXkrGSidd
pZ6i4khzWNEKD3mpCxzWKaIYfZ+smNcD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QrIg05aChQkRudY5W5hsBqPiso78RUy7MhaWBIFylkbjzEfsg6dEk7H348Wo
zCdztxUyzHTuH39Kv4uCH4hZz9B8JQaMPXx3Xvwdh6UmXbf+zFy/isivFlx3
bRgX10fN0cVOdRCaPAiHMNJRSrmLtSQ78V8o64tzBdTELFobcUM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hD2qlRhKnZ61/txCGUPI0XFNB7NfngWzwgzPD3SJrE6rDXEGaHbqEG4ji7qS
2VE5fI5saEzWKROWSb2pa1ffOVPQcPrTDsx4BEhYbrKSmK4clBWpSM2IBL/o
RAvZrtKD3iALc4N7aXIF5TUwszGqxXUZKZ36/T7rhH1HVS0F2a8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10816)
`pragma protect data_block
9EIaxoyMqTAL0ES4sjIVuLEKAqLUZ4ztFXX1Msw4poA9KEzw+PWr4Kos0BXd
EV9OhoDek9KAf9gKEHhkFpG3WNPU8wF9WneSngtSW0fRZZ2VJsvmXNz/KIyS
939QKKjHQyMDo+DCV4yGwM8SJ/6UcNGrZXnZ3yYvabNsXHUl36Z0z/IbUWrF
owcZ+RwuKaaP27drHQFzDllZk+/wKcqwZqosCB3ZRPtXwv94i+2zhlJtnSc9
oW4nSLsQzMjIiOGD5wGqg47qqibEITYsSSIR8e/BIhES/WxSIwe+MsUfsfj8
52tlxIPfJ6y5nc+p7GbftjhoX68agP76abw3BA8Z2Nvwg1XmIAWlvE4K/fgu
aU3o0rhopOOJARhLVWGhhUnGnEun8StJlttRW3rMcWAlT2mUPKVJhm2G0qAI
K9VwbauEXx7Vy2fZ/zAWnNwI6z+bZvhO1HgsWeqarhqhVLaEY9N3sEZi8GzL
YcGieHKnS4wARDaGteMSO6MLCqdTxQp0M1LOAnt9cWW5+snbHpgb8gEiw/uY
ukuVXDl+FFWD174WQL2s6ZJbzMatMtcqk90jLKcKKY3bpmVL5cvw7UIewVq9
eUuFa5KiD2wK5Xvj0/R4iTDeFexNKBGMAL19fm7C1H3aOyZ4AVGjWTDHtc/X
YfMDfbqOUXDXhmfOqr0KTF1gIn7yxiKUpcu27so7de+FN4/Yrn6wGxA3ItJL
OzAlb/9D0tgur/HFwAW+jRELRXfrs/VDaKJWw1mUvMM12sPS4HVsqmoZf7uN
giKxZigFBFEjm2DXXwQ4yNPBK5x+ZrIWm+XoMkRDouKU05a57PKH9ANsRT4b
k1vdfxuZN+Imk1ZnzxRy0xlDmmNA7vbNd5cAHuBMQ6vMrhUhT322X4x0TMgo
paoLU11TzZQyoq9yn1RjQTgJaUPhMT/m6q2jWyZvQD5Y0ONstTZJARxCQIkY
f3MhOy0I91w3jDoFMk/7nr+ZuW0L7FnEaLTNqjAH0G02tHGQ2Zk+of0xR+ta
RHE4Ci7RHMzY9CzRp/CsMoe9OHrj7phn+uJZfgnNlC3yX+qzvK2cxvqVkku/
Hv0BaZLU6uAacVgTst2QGG/mtfLgOxsxjNeurrVhHZvZtP3LtVTJn+oA2JKs
GOYcWWa9OU9SbT1oI+o88XyyrkxvaEh90QsSE/nIS6SESHqpuLD8mRgxk8ki
BTApEhc+IUVgwQiRKBDT148ZXEOtLVDCgOAaRnu/28C+66Ak1R2uqtb2hZr0
+AZ2LrCPHx1Y7LRUgGvUOtGooy/y+xK3C1nPhPe6DsP92gIVp4nCo2Ha9oU/
y0xgevMvcQUTmC4snMVKEx17tlhTdzr/2q8DvSZxzMYIHmVGKkxCGfGnaSxJ
FySi2otmkm/dNMP6aAt6PtlhdeYhBXI4TogYrivzbuGnjBhKmiGokmOie6ic
S2nD2InDva1VWtYmTx7cpgv5An+iIc2qmzbjZdkELDaRBomOFIGsCiCTkrJy
JwBhH2J/uIF3R8U1uNMijSi2uapwVvCGVuJbE+PEy1+AF8kfD4BjIJciKyvW
UuxTkP3sZEzDUiSs0ImXXD4i/MI2z77GkkOpmBDkpSyNAGO3kvjeV3QdrQ4w
CAjfHxjVETvNW+INjs5MMTRjbQZ2stMAuAlp6kp7JXqIpAWqMxZbIg+AwgTM
SRpRqxaP2YY5HUqT40jjeYIHYr2Dd3sTcwV1BhpvfcoLVfs89UwoaPAG8e5P
PKJw2dSNKonISN58TPD9NRvxvDUuFjbDXeGChnFJmSYXzbpDwlM6iQk/yPLB
o9n/QJlvIzwxEZGk5Zg00nNxurwmHt+sAD4os7pdopGQCeAyxVD3f8GV7xWl
l4Mf1+7jGuqwXNWdLEu0tz9C7f2yLz6lI1DzLMlHlIpR0a8drUXHz7DxZ2sl
41aJZMoJOp5PsEQO0+03GQHIu7ZhBC2pNxp656dR9UQ+OudO03i1FxmX+FMa
V2Z8fJ0tuFm9L8kJo+VzvXPNIMUc8HSY5E/bWBrIyiTthffd6aD2P6mzw1qp
5agvXuGo1ejp28cvtGnZQjMSaLiVoKXn9UaWmO74lhQbAPLRjK6eGPm98GDY
AvEpHc8hKVbTc6YMqelRKTzNczoDO1u+EDvzRuPQRNsp6PleU3piUCvavIg3
LnQ1XEQ1m9C9d0kb+nmZXyQG2O3uVVTDVSaOnHY3QoucCEgO/pPRlNqgHL4j
EQBe71WGeW1hJP3dEzeNjPUV+ispC17sHDM0fJHJT1WdG9MJ3iomCznYkmhk
oGQvFUAqdQsusgENRB19c6PgIqAlXvtg/7RpWYocGbUkH+m7Y3qZUc0lp0Ic
Wyn77tCFZZwaCxkwG6Reff15C5bP9RbQd80LqnJMblz43kYw11OCgeDjfYFD
zDh66Qz9KGZ575EpUv5zQAeeczsFxywZb7TKdhljqgYv1CWAPAjgpaRrT5zf
wr5gLJhClLNt59DoEtIzQGGfkYHbRshGx/AQ4pf3ucJl0W1lI38R5tM3NRrv
U7G1FYPXzBtbfqui44hV8gB/GDvYkUasUWebH1uG7/PUUbBmJUZCgjnQ7TGP
Bvi/Gk6TCo/ory3Yp0pea97oiG56MLZXbT3fc8YEfG4HJIRMnhu0iAOJ9i8E
Yk/gi/QicpNKcgv+XN9zZ7wHEDMYQl8U2JNfLqF5kkwAmezPAdAe0MZxxJ9M
93zMsRovwJi2LK7v0beu7SiofdK1sjwWgHfqdK3QVJwyx3cgNrBgiaSB93C5
Op5J/IPBaBC4zHbYKge1lRqL15sMA/zjbdCOZQt7e7UFIFy9atfFAlSEENnx
QGb11KJ9VKCOfeQO3VqYGWmwXqvdR+6KkN85fzJbU7KHfhmBzp2UCSyGfZoi
pudJUG3I68sb8HFgh4UTwysml5KWWjExL11tO5DDuyeBrR3xQxUm+44KIsTa
VkJyJ2P71De6TcyUGNO0IC4scNM8Gi27uMyK5UbIGzu1XigX3D1Te5Groy+n
0LHgxnJub9TQLQet4K3f4r/g5B4VvfZGE9BzDrGaqLO9qim9ioURS0J5ghoi
D3b/SN+fUp8j4bqF6xuWc+NnAzacoAGKDuyxyMmxTJExqh+jH6/tQYer/p8D
CyJaxwc+SOhMhmCCHht/0EMtlf6cW0Squ9MR6S7/mLp6VC+TTgDc8J2yYV41
srE3Y3rGp3fao02lL8hEkXCbp4iDtzTiwninZDOBM9vjmTsRX7D4+k0y2Q8J
GEG0cruqZWvtlG9AEVg4VhZellryKIbsx6IIk/KHiFNxWk977mm5IrOmTu7e
kTVpy6y4SeDIaE+ESlw4tJbdqFlfKIXy5HAefwk9LRp6R/Q3YQAZvpODxovU
7VGwSQeK+odM5VBrEu4GJYHFHwHNR1lL+TSYfMq3H+SaU+i+Edx4ShgXcetl
DRs9RdOhdJuqI5Nl1OCctyBXhtoPkhQVikA7GWNTGAWRRmt7o1MMKjJvTEpa
sxmIWxtW7LegSlYt28xmtXUh9kWJdUZc8IICCbofkLdZKBmTeTSA+9Ow3EP5
ZERq+G2hZ+pD9RWyxtDdVG066W8iFXRgvGcD2K7Qyai1qYtcolTT/lWZThLS
OJHPhbAms0LiGvyn7rrpRrDl8YYRArkzvrOXhcWwYZFfH6yhcfPI5NK+wTwm
EOJvV2+/dkair8ZXc05BEvmbpLr1Ju+F+lYPXFIhNylg2tSdfeXN35jyb44y
egygKhJc4wSJH2uDHUGxONgai89xHet4nSaH1Wxe3ahNIAV5Ms0eXcK2HeuP
gkEOdRwR55VtOsxWBJPmkeVFkhP5XWjqTtUj91uFbAXjg+F5P/ldRN+nxh2R
EbJ8qiTynUL6z8OqMBKtLnNYzUhF6xx8TW0hfv3fsrrkXsWU9dzOJGQMBbL+
sNWTgYUfG7278pnXuZi2+ShEiEflxDdsE/0TJLp25bZjRUhi2YBe8sho/3FC
Cr4G2L/FVDRmFQMZJ5varW0FeK6cKkeOKEWP47JH+rf3M9+te+iXd6zU78Mj
lsBQyjMVXpKKWZEIXAd9t8MkSiHrqsh9J/BVTxNhOee9lA1TtST5pZlVFfSS
fxUTpUopldYv48fVeT88S6vh3phvGwndpSWVr3xwuWiqmG3g1DZdUSqv8FYW
lBPqEqU8Qq9Fo3ZAb78IFRzorum4aA5WJe6pnAGY5/mDqv3Q7rhBtKPJpjUJ
2+sygPaAhqo2swTrA0QThFWquuU5DKnQ9RHs0PZumEhenUoQph6f3Fvx/UEw
jWe+BRmNdReZ6Em1zWrzFpW/J7P8k21Ehl2UxCrYBl2b7Vq8J2oITmTis/4v
vR++4amhyOyKEDhBjEHvOapMebWABQjm+g9YJEGcf7xJ9fdq4c2xalCcH2Ck
sDpzI1BxQB+Vi/qbt86F6vgkPW8v7lHhZct1buZFFaoDPMRirHZn527wFVoI
iyy7TCLf+S+xEoSosCxX/QfAcXXcuxFfQM4WwZvaC1/lrlnPuNpwRmhglfM7
Iv64Zyr7VpriDtq81ao9WYSttsaKW4Zmjqua9vgqGA7YBYFiz8ewLOUpz6g9
7A+9VTcPQtwGtUyQqwtS+AxPYOXYnGzGyTgo1Zc4LZvCmxVZT1OuK2zVha6c
dXtH9g9ehIe4VfCaH8pPDe3FWypY9TbBprq18HFjA10GAipRY98bpqggONQK
RxKM//ITFwDAAT7lx9SjWG/0eqpLgdXrq/XRSkhgJIENFwzeSYlW9bJzGnGU
c9FpD5On5efR76uCvPiCkqvtauBDFoWC70QFyWHfvF/dbnJYK+GDxghT5eOg
45Qxh8jg5/WOs63qMogN23a1knhgBeOMBp23WagolPFgAmubn9Vp3F5Ybhec
4eiE6ORDxc/35G9Q4ZthBvyuYHHV8drUU7tZKlspGG2i/CDPUvIG8MdYZ+3r
pL+BRDWO+6obOfdWA3ZBFCb5hQcMD5ZshJ5eyiYBfcepUhnrbUClCVTjX8Zn
tb39Eym0raMeypYxzzImU4pZnnooBHrJD8THO3Bq4b3QjyjV7zD4ZxZmKHdx
WKnDHt2QJpeVhfhVgolNSJ1vPS1IH9U+D1XKn3cwwBKAlKjseHOZyFZCTl0F
TJzZJZAwwicL83I8ArqcHGJHwpvyMNJEuYwhvSav5yrMjuCrGTXmv6RGpkvt
if1+p99seiBq67Iywo/cymWx6TgPCaAqfGZ4lYImSInlpCWVh6pz4MrkiWlI
PJSRAER1F7YsTk1tm5X7Phr3XNiF7dB+Ts+ic/JDDML0nO0N/NNhAWhdxPJ9
kB9Mo5g0+6ZQhPYux+sZhrmbNAKGseGFqydPD/5jWh1ux0nKw0nkijesdVj4
2rSDU9KKT+tcIqEgPzVGcmcocyeXvZn7u9RS37LVp0jtmJ1qnc+5241kbwOH
UTP+j6p4A+9+4C48fIkpQxg333QfR+UuuhIg2bbiAz5GI1Aa/PBVpdljHcm4
mbZTfRG7ZlvurF/eKnwpiEEscgrNF0wYTVfQGmMBA3WA84wG6oscoC0knnmB
yaMi64dDbtSB1VaX7tPLurowKqs4ys3YnYpbqEMYct6gSmEkOTNNffp56h4T
Mb5IZlHwxYVq5qf+C7eClw9vL1sFu8ecr42J30A8I3JUmV3MmTDVeAM1hCxX
Pmcg+CDBbvCwpQOErve270oHUlTvddglOrtiXiWOkDWcw1UeslvYStwxLpYX
bv/8sYZrmUxwf9xGgzMkfXT4PT5e/PGxWa3whTR2Hybo8Y2mg6m60FvOu7hy
LTz1hPc9ESXWoWJSLXCLNoUuJrlEIZfcXSSw4+e5F9MweskdHqYnOdV5KY1I
0kSzIoNi1JfPIQRW7Gf88G/MJyyhxdpXVFTvPqUrGF5biKQ0bw4krI5LLxew
pmUjmvo/iPyAdzydj0JIyOoV0UOR2cC+a9Pr/QOL6+LINRY5cf3K13dww2cn
XqWaLuJqrdZMA3OvwPXb+HI9oQrKrryth5IhWdXgkvYYokaQicr1Y6EjPVkl
rNvWF2w1rkdT8QC8/TGBvWJHKsL1IZXZSkigA/9H0TnQoXms0oxzBzhjiTiS
bs/Q55aSyLaWNZEeXrSQhdVqHODgCQc1kpQtS08Vakw0WMjKskp3DcgWr7h7
yPR9dsJUBDm7xE3hcXyB4nHYVoT0oYvj2yXjvDmYogM1xwijGwxLW0ifKyI8
9EfMTYJvN6fQpnfEZx/MkIkxrtYhjPHGGZLXzQvi+3jvapGiXZ4Yn5IqUTMv
MaqYwlgmdU9tAWLFfO9tgFuezkIO5Yjlq5R7e4BD8FxQuJMM/updSiZ2T6fs
k6rexWOvo/sH1goh0enzP0a8TQOY/ky1hjP74Y/31j3YWeaewGT+e0PejzdW
TTVrXvF3SQTR2Rf98Wgh6/HS6QMY+/GnrErMPIUd9aTuFuWkzurFVQhIc577
zlV1M/e89vXq+spbPgBg9GHrvrnFGfLZOgqTE51PET7m/pU2k7W/ZiBDMNBt
Ve0d18/IA3VEk/QrN3Oob4cKhFxgoCD4QUo3h6CtIWgVCh9Ws5V74C59CUwF
Pi21pXidnPYQbPbB/or/aoy/I7Jt1VtGqheHC+bsDCU0HfUM7H0R18nsiyes
EeNE3g2SwfvW9Z9y8ZQYvqg2xaqeuYi9M7uG0E/RWZkCrGQgsYDnmsHPKR/t
knQCrtQsGl+Ekc1zDnbP6ftUxNqh0o1s09OMnkS6CUGKjdLYNXvtAOg4GaRn
CdgAR4ervJvKs9e1Rgip/zlKL8gGswK8klPc5Ff/FrePpf2gZsOUeTRPswX3
G00q8BgkX3pbAl3QB7QEC48Vid7IXnrfp22NwvmARf7IzXjUIZZetf/9YgLF
/sF12D0H2vjsv/RH4ZxMwpfw8alDM5oBMnDJ7Eg7hSSQebOOsmrlZtfzN6Z9
S1LtSkOq73qd4qCtQNAhWqg2Wvhl0GE1HmDzNQexCEKcaudRpeFm5BiBaNIW
CqUnI59yP4F8ZxNqVRE+KKETnEdyQOtEaoMUNhyIun3VfSFV48Jhd0Am7gZl
MFVP17uA8tZQyo7iNCr14ETCcITZvcksaJnR3GLb2eg4NicpJTl7T+69ydkq
LrlcB99NKNm3K8q1lPhEq8LVYqmAEvkg4hwYFWkfj7xwrwOL5btvk2CDya0E
YPAL6IhlDOVxMed4GeNOUQuuuW2TbOLaq8YJyKryQVU8V9MYBrr2sfgQu99m
LsYq75Rl83gbeEkzdDy6G7XhWLAFXuJ1OBlmj0nSIcHKY2BYkpwxOW70UmpG
M6RGPb6fZOijdhs03KulcIFZQ4OGLjkffVfkCw/+TgjyTbXk0grP9yDVZ7Y2
dmijXH3ukqkpoPsPIsTEUc/iFLVSSBZG79ruw2IDAUQyG/kcec1oN2vT99yf
dXKG7jJfuraip0QYwmKEc6MUP13+9rSauKbUj254AdAVe6ypf3IwnuvJuH/r
s2hJZGTy28AMdVyChlQ7L+Wkw8XCMnC8dWOjWTpTqTjrdeAid6InB1rNlfAu
39szOvrNplY0G7qmQ8PzgbSZPxJXmIDnV0kJuMCUxK4ESBzVdN95Gxqsb8HW
61zgcG+o8VCFAOL/fmUzUkaVWyMcbNodLoUwapj9+0GR3fgCcDFnXKvUq8tZ
luWnk6PkmJfIYtpTaw9Q48nagG2p8N8ctZprmEwcPsQQRPVYTH+pBJJDfYDV
rv9muwRPCZIE9/RShTB+eXAZNxUtwI2YTGOMYrMCLTIUQvq4f99RuUTmKqMq
Rf9Ewvh00H1im+ph+6DIcdzTWp5SYtLNbT2lGyW3ibFPQu2B+T/23ZCtYNX3
P6bhBI7Qc6E6eUXfcZi6o/s4NN3xusCCszmHkLrTwiAvHhD9WZpvnAb9diu4
oTvZBG2VpJ2OgxMYg1DtxzV9r9y0cUe2QvPjPnlGc3GKhQdf4zpSjELXhAvw
wXVhBVkUAwxCviV+PmeYL/yML3E6THvn4lw3cIoaUgsDsgD4FsHTuwmGp0kT
7BFak34aZsASvGbkRiS5LBqrhfAZv+jTrF8Q7X/bYcm01ljDhiHTgbeV4vBe
EbHI2i5gnN/bjpDG89Y9oQ8RdzrNEgvn0iRrCj+bUkh69Eg2faVIG8hijPjm
fl8RzXaT7mSVUnZRJuUARSWAeLWd6wITudQpDYl/CCd4lS3+BQEkWWJN4lS+
uzej9DB3A8D4SBwlTPVE2R5WMEpzvN/s9R5qhdrH4rSI4+vJsC+JDqaKYMAT
tRRHoPqwNkr0igwcxppvpJRG1NHxphImJsHpR8lEhB1BY9fQMsCrKxF4d0U/
DrlWUYeXMhCqYkwUaHJ/bn51M7McoEc1kcF2uU7Du73U20sTxKfRs1AGyZCb
Ur9NDH4dgz+F5Ca17IX/nf5xsOOfN2UdRZ5zmvaU0b5hf2eQl3dRpsSzclIe
v1sGxJBs/Dq4lswZtJAnyChXbW8I85uF0GcjGZKNjI6Og0Resz5DnRB6WYbt
XxU5/cmiCqtkrhoSCB+JLuUjJf2aXLxV89ftX5FAp5M7mDhunQ5Cvv2RlHkn
BqYjKJTpN9Zkc0+llHl5aiwP82vBph7P+Nh2R/RBNwgn4lqn2ZDpB8yupKgj
6PuatyUw9q2NPTDIANvbVt8bswRMlUPs8KmijWI8Fdtd9bZzVe/ycmyEM57X
aJnjrG+RJCIuQcCIHc/XnZxbktGKHlxlnVXHw8jZKsWeEQ3IxaqUmRtEPUqy
+fVRqh41AGENe6Ob1jusxbaK+/lgIPelb6A8FYzTgyR0BZNWLV0waGK3JMmH
YN9mRMwDfz3s4k6cw5igayRDj0W/EusuFYlDdrtKzf+ns89AFtZN/f3PAdhM
/wOp5Ax0fInJxCenaicEmtcPz9psVoyzZtaMfM/No6dpjiNcn1lG1NLA75Pf
x8MlYcA8yd7wx7PLs1xUhpbYPBo/S13hm4PLqEkiLHFnCd8+oQIuHOzDDrWi
7xa1jHV6z06yZX5hwEx1UKJu5XqIz4RChRN/bz7kZSVs2Tqzj7APbO+fDdkw
MDi9qVSB1TxizDhtpKN1JoX+JICer4MHiOxcX4BMeY8xzZJ2SzoVqJ1C9Scn
zQ2oe4r/ZY2OEl4cWqClPhEg/BgSCUVHd5oO/tDQyPpDjFlcfA4mp7JRuJTG
UyRd9xF+P1sDxylgDKXpB+4wG4J0bfKhQAJGwpTxdwTHZywlfpAQ6bugztpU
9B7Kq2HbRGYjXU5tosLmpmipugeFFSEH4oi2ODhXn8kL4+dmI0M9xQfIkDZj
k2DuYmC25KUuotyq9ZQ35+e5MZXXIyRil+V3wqbXnJATeZvMvKwnsOEIoF1W
NKIbPNrmjx2ldMEM1XGExu3upYUWO+6VzEBH9WvwqPbfBnMjrfez6GIZySwj
DV2PEpMZBxHL7yIynXojTH0qN5swNQJMOtIT6XMwTAqULU67mdI4Pj/OPxVc
euRaMZm1bFIgvJQyBB+wViorWu4zWOfaMDvvhvlxFmNAPGNcb8uGx4JlDp3Z
iCHMFsCFIyj40yOo7ZE02q3BHZcBqXqrQ2W0sNh6Dwf377hDoWxZHFgJAWRE
d+tg7wmHgrW9SqQDsWhD7iknwAHhYNxJV6ZIuLxt9M3iNpjsCbv2ZSHo0ijq
M9s45TMEWe1tfbxF+5DGeXV+rA+6AZ20Ycu6+zyAyMF7lFp2WB2NqxzILP6/
ZSpvCGspULiRJkVIY+qSkgGuKDFWw2S+dbmFtnQI4m6QQUCj2mSVXj96d6md
/tBgsTcWBNiLYaUzrx48MKXzI2KYpAwdfLkNdxYVUPeyG+P8vJIcBXi2nSir
gn8XC7xLK0PKLY+DtCCbLeAMyRArO7yNV1XlV9UFB0q4lkq4OfDzhj6GM41S
6CdOMtgb/XRYO4cIYkxwG6cg5NqM7nVim37omvvnvobE3hnaB4uRHWfpkDDa
iuoECj92WsIoiHfoFZjYWtDJzm6zjfjWnmrntvnW5GDmqu2v7d7ibJm6H7QE
n4hkzytzBYfi4S25Xv8X7kskKjYjAo4+A2xYCfyr3OzKqPfPpTKRr4DkLEeK
knFHwzYYOvBefBVkvvNM8JpIQCSJ44j67Bx/yZCe75t5HAPilZL7BERc8QvV
j02Q6CWF7R4nZvQ0OYUVp9DizrZLhyeKipe2e4I09cbgT48+umyxvUXupCNU
ABphqdrenZe3N4CZS0d2btyopPK9ZEwX9hRVd6MucV7n+ngO5su5dTsnaN+3
srsU+IZYAGfQ2BqPq/F9G4qLhdPKYprKxDpO5MdlWhnXOVp0RgoHcoL9+w/W
wxyFslFuP4m7DsyDcsFkw9Fe6bnh7pH/hko1qwZdBsBvngm3ZT48+kwffC1p
e87SUPQNl+3nrjR2u4TtiT0Vf4Qy22zHCMrLYFh6G8HerjpDDJ/c24w+BD6p
TN4KdPw7UjarlT6YyuWzJNGSlindPFLNkzMqPFJOkally0XHYZC4KMVpO3x9
E2ySjwJ07r2WhvpY1Y0ZaY/nDDibjIG+Ox0n9KZz+pnDt9tglVDTL4TM38W/
dRL9ozGL2A8IyLGbMmR/gKllJgVTu1pzyI8C0n58tMVy73/lOaVd/OGhAfhe
N1oBilZMmHmY1+U7I3UYUKk0EwBnnjaXq4GPNKHAM6JYmAO32hdg5IbAuF3X
EhQXI625BGdknpZwKiXvmXzBLM8f3yardOJgxib4cjXSqcyBV0uctSy1i5F1
4/FBWeZ6C3NbjVVaoDaKqsQqpeORbmpNh5wQfuMkp7BTZFa+I3wT4HU9mUC7
16uzoYG4VBY/ePeTQw2LFzEVuKKVHv54jGhjywDy0KOq/132xWqcVkiiRfBb
s2s4g+46kQkFQo1U2yBZrcsup5K48R1mH36ynIe2LJMTmh56Qiu5KzoXfhDS
p633cIvHpl5v2NndhYCr+2ZqGj3jEU/1tcjBY41gPciQ7nRxZtmo7kaQ//wE
Mm9FiIz+kmkl3DBajT3K8Yo+Ft7tbq4LGIJuGXmGVNgsDKKklUFTdC+fgPz8
Emq+DmtNIe6CvRCI6Gw+CpMVqTYW+EBSKh7ibCN0JZ6QUkfJ7NGazYpWRj44
QZT3DuL7HVPUgHUIzOU0tVFO4uLgWIFWIjtcoWcVLycyNifDisnZma0P9hVc
rOW+P/FUYpLS/LOryArQsef/dEvio1fX9W9FFX4CbPU0OAG6N18pNPC2kpmL
XQ9ykTT9BJcxtgW7dQPGJP8jUyzT2jpA7yfRLlERrvUncghY1zudA9/4PrSZ
rTBXYfO+4m1P3j0xTTAXtwkOFAz/KesGxJSte04+urAKKV6DJ8hGVYNs8sMR
B8eScwVR0SIjT3S4wrKtW09LXzkegzXJFaqWWQOUiwFEzSVaDkQWypfDdsO4
EJr0tQpjGKWJbzPKlxvGD3XJRWIWFZTdT8HggU+Rdw/2EhOSiK+lwj6/bOQ6
WkRm3asNjAu4PYWhV4FaNSmuMurjxvx2Sjqzlo46lmf+ilF5UoZ+iDplmKoq
xDP/pzOJJMOAOe5dP1RxRXZBggk7yZCSX9IiSUK0xenIy0UxEb6dYBgnljwa
RF875dpcPJExWQ/qisG5zde8pODbUDjPDzShkg+wMaFYAt/AZqLVJpBx+7kg
tGT4pYAFYinM49zyyHcJ2ava1KDfItJfetzweoV7fZfLMZAxvj8JDq4Sb20H
Qss7twJ1i+DfVfvOrRzpYsvxxwCi7lvmg6y8PtVbcJv+0+zpUAH/F9Jw23dF
9eabP23l8+82uLxfYL6lCgZVRAuucHurtsNFB8GLIfnRyI5BYnIVgF3MpIqb
u0GF8siW0W2pwPsqU9q4cGOcgfi9t2yYHF0Eh1sjtISo0VdPSuBkGKH1/h12
nIILcUJUgjVUZe5Z4/rR3R22xhDI7I0k57I2fn9dtCYxFd8V+OpvUrStSEUw
r+kFefHoicz8tm0mduztrgNgoD0bdvMzTQQdvlgc74NHLnJMKWwyZ312DZxV
XP/feLPnFKGC/q+IHSwR12TcTmmIs7Lo9pFReSYtoP5Qr02RMUBO8vxZlYlT
JTn2ZWZyAAyWkOvOepqBFHXfskCOESMeHnSMVbl1xQLWSljnfC52JjxgmBux
FABta1nkuoxHGMp6lIoV/7/vuKvIIqPDHaSbyEzi8afaCi3x14Z7ECiZ0fo9
1LyBAVgJazPVwfQZpbxmnQn/ne5Xbzn+2dtg92z1esOWruTxWx7hWIlISmn5
5TIH4pxrgYBSh3yVBH+CZJLQO8Aqw5zd2xQyuFojL+sowDuYRgJCc0LNkOJb
MmO8QLw77VR+Dwg2i5yLxvZBHmZ4iYZ+WvcOX7ruRg0Z4RVj2PXXM6ezOiWI
qHLE6FO1YZRjow1tFlKJov4zDDxz60nTD9PNT+W7CXqFn6neGOj5bRGWiv67
9PmbueJV5JEPalKXcC60KFJ+HHCbg7EXaZO9B3WLdGRIGmXpADW8CtXRQEeZ
F+XxtXQqZmjeLG1mDkZcvvD5uFTfRE/C3tXgYyN4e0+0q6jukxQp/yao1u7a
q8LtubnzWNhghNq/wDy9Nq8JIZWJNuC0iEJQvKaCT5/W/V/Bk0U91EaK0gv2
EZ7qQUtnAMkKdyHBImT+EPp1H8l3AXr+Au7ZTago34f4lcksGJWooTtKlDEt
uNrkz3wyMwI9CJ6NMwWZBqvMkjd0mO0HZznXjLP4ENy3m9E9bIq1txG0jHag
ryguvhFE2rVuiKKRWnmnEransVM8ij0z0Gk09afs21hvFUTMLomH+PxWX6NZ
ERNUPWlliB4xHfv7IeC0u5jpbXPBhhkO+BvvZOAYnxGcasa5FiyAnpcFj7d1
RLovlI2zuFrJfUaq+M30udDT/n0jFxy+nNA5du8I68RiedlXtfCu2bEteqYN
f4qoeE03vDS9LaU/bC4SZwWmq7dItlDJymR9Zq+O134ew5KxMgnL3u7Nildg
Wla1n6gbAXaRnJT2fMEY6dmFQoEABS6SRLSgIp31Tih3jr7I7ZLPpheU1bMC
cg9F2JqBYWTmw3lwemJVW6QTpFhArq4+xd+1MfL2ISyLB3qaSkTs8PNnnMUW
jO5Xd81FfkXzWr8tA398QXBSWHlnCg4kGo321cp+e2afLraUwM2EfmGOU1IB
/tS8r2mnIP6tJCvTY2wExPMe4xaM8CVGoctAzzmeuavxC9oX5szhfoxSxQxC
XnAMYLiNl7G1GXmVz3lZJRmwqmv6ex33EOIXSY8NHXqApXC1iv9mGCFlNohX
qwYiUdazfLH/h+POUUu4CjZVOwRm4AqgU/2AK1y1iRkt0A1gjH0X66ZrmmOM
kIJK7i3OEsRLQ0OlR1Q1eMVpnKxn8bd+5avkYhSKrhbTo2rHdSLXr7DHNKUc
daMDPdWpKYmn9sga+VSWRplR/gajFj92fCBdlzDNxoAM0GI99weNBF0oXlJa
cZD2pj8bJ1LimAsUSmIuc+s5lDZB7EJZPj/ycsaRLYOCit3CGrnMaXo0kvok
cJOOnPM4tAkzRCmHzQ/ScbeLlxtw64F+nPFZ6a9QizpRBNZ6pKnzm+xQfuuE
Z1YUpAKjlVC/OJxBeVlkMqG5nzVTgbfVFryKPmFza1vJifVj6uAdaVxIr9Pg
j6kwLS9ts8WirH7StuP4dv/HHUROTz+BOtKadrW6kJSZf7UlhEx2k3AjlkWi
jo3xHq5lQQd+TclcJ+Tc8+mirULZX+kOczhQJDwqirztSy6Xi5rsNrNGKjAM
pLnx9AFK2l65oq1depUkhDQ8kixJF4ovMBYEIQUWwwWkaQRj030T6UuzMt5m
7YjlKoyWxtit9nyIC63sYMkBzXO7zN6uHrdEubo47qJKC2yinXlWOQ2hf0Gg
KrF/uZ9prN06lK2eG5nmu9oRpOJ/jEYXsTsQM32G+a2RMLpHchyU8m31I5oJ
2OhMEqjGe74BY29NbjndBRMmoRGhAn41Og7PYXjaKTs6Z7VnxpyZ2yIfOMoR
mVL+tf4hMHF4rzQ1wG9DtcN02Fwqu+h0DqGqbJDZFrqvLP7VppHAbAUTVKKg
QjBHRxeQWJNLPyk3MIV7uyWEd8gNWPgu1/q6SQ8ZuU/BpI93VYGMY5/gR8rh
FBOxYLWC/j4E6H7Lyhqj2t2ley69x75u5CSAV0sVKM2kreR4eHz1k0HxKxwF
H5wVEF7LM/tS35cmtZgFtu017K7MCgOubl9MaV49EOPLfXXmvVELIlkLa16B
cOsxAyNtn4w85Gl9TNPRqx3VK5Q1A10GAz4Ez2GxpnNWkapJCOXRrtO/Z5oa
cek7esfUabkkGqX3zC7OYgTJUksgKRu+FNqfnsW2lbxg/Q+IzDRlr1yAcaPx
ECGwnQu6orgI5CPVCPgL2ufr6gEEJnKijB8Q7tbU3kq/yTJd6YRiMjSMnucK
h0mPqSaS6LgvXEvvfSXguB/uQ+h0ENbU63Xb2+D2vSHHbryGMiWZS1cuoURd
HA7sBshbvSAhxp8zAqbRKg==

`pragma protect end_protected
