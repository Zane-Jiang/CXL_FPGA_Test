// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YLI4nqH537drqz2+rsCrDK42NPwF6brHEAffwabviDHAaecOzbcOQ/zGjDaD
eURQZ7tijGJRjohe/GoUzSaKWEh7XuzvZ0Bw3RYn94B66FvXz6Ye8o/AmggY
dvUV5h2CXHuuDdmBDP5VPqKcEBd3oCzchLywn+uRHeaqxzxtVxe080QqlkgW
ZyL6hvLjJKGuaBuX014990UV604S3VL8LOBVrusu8iDUfCzT1au6aqa+7bY9
8l261191h1wBwuUNr1VHMyeThxhlFfN/ieEmDsbXqsetDU9Tflxaj49kE0S/
u7niJEU5+teXExVdYhYlrFonuRq2pBh1ZDonAidj3Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xswo85ibG40UphYoyKAfuvgMgiUmbS0MTLCQG+hsNc6h6/EFpdjGkSqo0DR9
vn2cZCScEIGDWdWycX2WcMnox2nxSiY2x7/Nbd52QY9cNjDty5rr1H3M2qTK
Cpo+6wA76wlJzn3yxi+HwgIynLYqsH2GYC48afusnqZNwlazAOxYxsfRc7p2
+RK8LyiC6ZASryroUxikcKW719g7V1vfzDC7CQnu185V2F3DWeb5cpGe2oqd
2QGToSC3oMMNkvC2GZPqmLQdW005SGo2h1xtt3BwseTx2ZNMfS4kdtMYd9hD
J9wmtjEp8EkjTCN3qIZea2Guun9LrZBF/IUSA7uiYw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WBF5cj7ZMOoVw5WeWYsWXQeWdccZTug7EmGMiGUebdQIGoDNM21vrbObv1Hp
6BvK6HFpuWnc68xlaSxQkuvaKnL+UQdsQrjr+5e7CzhO4LdWV8JOVf44iHC+
NWpz/55Rd5ASs8UpDVNQS7umIFGOU3xibTbn1irIirNpIJx/aVGT7bE8fwEP
TmUvFUHoYpTxnD0GodIOycKkpN6KQN/Sh+DiYLnezhKp+tpq0Grchk1mfgi+
aArnyWbGMk0JTwDxeiaD/Gis8Njm9qIVgvYRgwdsb7ApYuQ+C+Ydede3TDT4
4Lpqbsc+kjfQTHN5opTsIz0bwDYRALMZ82IEQXVXaA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sJjTqc5PwYrOiKSMJ2OvEF6g5EkKJjnddGUM5h9Pex6gh0T6ChgvClvwzZnl
bNJwR2foTwnVkCLmSWm1qog/HLfjNimjzXHha1bS+lTLa/fUrkx+vNkBS+x6
YfRwzmG14qojkL9TpIdz6YYk+CBxw+gzZEDuXiFypiU7I1Vbq6Q=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pjfoxbEh5BV4OdDIZcgR4m7FmUUASlUJdVYXgBTnguNCKl3OFw/VIpZLH0D4
2XjnZn0P5FxL+aqXNFyD+aWYI2sG2xuz9NP1sImgZlUj6wjdIvlEl7qRWN99
J6Zdxi1zsVw7ng4X5cpLisslMwf7e5Cb6qFZiW0nvNZU2qLyAI7E0a81wyEb
GtBeGJoGaPrCKIccZtkpU7N4T1+12KNll35M85h/n+FhH9FJTCxxJpN4AeZ3
kR3zWB4GrDB8FFIqTcFzu1DlzJ5WYKZjrX/5EzO4kZEE6nApCtZAGEyZESoC
HQliM5fNbyboXDvQvXYN88Dci2EL4piic9tnWCOftje7w0g2sOBfwJskcxhK
IB3KGs+jAvgvys9sjW89gQn5mdxMwbmwZylo4blUrVHF/FhgFoLPdS/qa2Ec
ggMm4KB8kcv777BsUWC4H3oIWd5UXWI2oC1q9T2Qgf48KK13tnBbECjqIpn9
IQ2xLrc9L65JGFlQei5c65jkQFBANjup


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PXESxs/aedqkTQl6txzMykVxHH9EQ6N88z6vrJ/WPBmbjmNZ8jqfdPg5G52R
z+n+IJOy/FxR0xSAHtkitztjYOX4T7q+p09TwimARCjsrQDHWQY1izCG4LmK
/TzHWATfe2hsBbcptYrXpBYY+o2sOE6bM7AWu/sW8CaYqG+2VXo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lmHpLRTjacgdHkIxQHYcgnuKMhjRUQW7GJoj0QUlgBYq5dCYyZnKj4lgV451
Bpg68jjICvVkMpmixv6Qlq5R2BgSON/4AvVmx22ePUGSXKyQgAmotLQZcIb9
wgeK7iE8SvMouPJZpJxvI8RspusMPr4etlJaheHWpbshtNDImp8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
e/r9yoUVXDmzoXYfBqisEnUv5RSF2QWyd6VW5DFyZHTrod4Dr+dwbNTmtxcL
I2FPkvyVxrJ6rPP7ZSHwR0+oQ37KKdvGr4Ga4ffrsgkQIIS50BQmbWvrkUhS
pS77rWYSqk43qWWLTxcu3AzdEuY3HUsdyb+qXOXZeFkcE8SWm1zfpHD0P6Ip
zhef5csFVghqzSuJlL/pRZqstqOy1Y10a1GYYVoxPoMFhUkx816ogjm0mgKo
U2sT02kEkUnUnwmXqJViNu3YnNg72rw6zVA+jDstufQ+al5GjLcNJoXV77D0
tNonH78vkIklz7Wm2SvwKL3BySqcB1OAH5omJ6yDEIw6fhzRFytPdVJaMGZe
U9m7n6lREalhphIwJrZnZ0dnrg7czl+GKquBFo6ZFBVfVEGzYaia/U2BTzdT
ElAcuCov22fR+UGOcw5hRqzxYGG5hspLaDd577RgfVrFOySVSyGqbAA2dzh3
Bi5FVkvobRHpaxAFSh++OQJJ49hjK9Bj+kT7xyxXm0e0UizeKdsuhWVTQAE7
7oebV/5RNqPgY6x6qZGSvJvOt/t2WudTKepZ27SgG2lZJLFB5ZY+hNGOj6cg
afuNU4uCl8IMTZlDEG8EmKMVch2s243ynQJZFHyqfG/V/8lzGot1vsOy5n3Q
ob7hYC5dsFePdEIuDvZe9DzEC05WnmkSIiyo1v/hrf72tincxYmSiZ5JrIDc
wVMwnngYcDyvRtKqKWL1+XzrHDL0dT/m1t18wdPk2Uji5+Hto2SdsTJjRWVa
AKzaUURoVIG4QVU6rDMFbuEoc3TTVGeBZMmOHZyMvQPtIkdOv0jYRfHWkUsJ
pVnf/JMTBh3B4Ig3nU1AMuYkLsCe+89jsDDY9apRnqFJe/Tz0SzJhWK7S7sb
0VQz6naPSnYROz1jyXavhlAk1EjbKwBCpOqv0fSQcHtY/s1EDw5OH0CawlIQ
fP8hskR+YJhz6/G748T0oB6EBDYCHc01KkgSzlkqwgvr8Na0+T4IORjCK0L7
gdqhBFtyni1ISSj1ZvnubEOVyQiPfGDZcypfiAKFZ87c3nYPhXAWz2qmSOeF
/9+P4bjubFKUmpjskXJBj2pc4viKuUunRyYtpmd3jGFrJckRvaxAjgUkEZ8s
5+Vilrse6W8HozrgILYPDSQXuCG+wMWaZ1QZac0lRc+OwvmxR0qpjVsSDVOn
9TyIlul7DrZW/5tu2x7en8Y3YXBpPRo2sXINmRiD1zuS/4cDC0UEjXL+JgMf
6SXmm8jIiBAzE46sTqDV7Vsk4PoZRO0usg/Gokm0NyqvfCMFEcgl7ziTT7Cm
oooeaYgRVCkAr5m66dv2pNckArhmUtRP9t2ySqu/eFSt+USnbNFOnQDh/sTn
djhhplmTzdiT0agFtxh/VXLfGDFdQgl4r6xrBZh+oxQFGcW03Fnd6jRff4mk
TBaFMpVwy8MvEw3RJmqtxK3k6fD2D/h6myj05TVv5Q6+dJ+jM/oICU9wHuzQ
RlvqFxPj4YWU2rUxUoGNSYgalx4VEIiUWHAOVKjVlbsaEcE/bQNTDjNsAm0C
UpjtpIYTWehCGSXsSHkr8qJnTPZ9IJE6unvgV4y0D44SCuvRHxck3tviqAgF
HV0GLWDWlVt9eRQCUMKXVzWJLY6viwn4DIDZakvfDIwcMV0IqywzckOzaH86
NDqa8IwOZLjs0KOOcE9JQyn+06CVwwXMroxnTuHDdrWxyd9IHDc5S0IQuUOq
0hx5pJt7+09HOYbKjG7kfROniD6Iypzf89fSeJ2jPwkpNCJG4T9AdfWLI1N1
xdzlXUs3eIKofPcTxuJDiEj+DZ4JFawUkZ4=

`pragma protect end_protected
