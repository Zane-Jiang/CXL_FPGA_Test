`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
bxW/NTGFVLrdMRpyrImeTldqg+heFmR8K+Ywf1hnkoWjK//QBPm9dtuysQGOBkne
u8G2wYm9/icRPv7HjvlZ9FeLIWseaxuJMvCVeE/ii2gBIeGfcalqQzAoMHcIoHYm
hepQPQXNLS8Vuk1bGnK2COXo/kijsPGbcUD7CskzftA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 15568), data_block
+f2riXpampE/AhhqYm2FOp4yDbjhwG3HmU6/Ck/CO3k72HwQXUA62MFgiSZSYRW6
K56snOiJ6XtHDnJHLkQZYdBkKLNC4r348vco2C57BIC6ek+Zf0tXUDKrAZ640wse
gmZuyeq/7XOCjqqgxVQkr0gXIA7hqCjolgm0j9kNp84CHkr4z3DCHGhYKK97er0Y
C5Hx8qf7LrnP3KZiKWed9haZYKkJjEHiJheR9+q9u/vAFNNxDsVhSJLNDMXYcnWV
a8XcLZgDVozb8Ax96txtTs3WUj1Fnp7LfMmASPgLdxOvkN/yLst7tlF6OvNvOM28
V9dyDd/37n3lj4OcYXS+CcjVJAfsVt2VLcMXOWhwJ5TYjpPeqelt74crOw8DAS/w
SqwYaWhvDXLTzknowT2t5VG5/dPLjUG2RpmggZhFEzlsHegnRT0BVkvnYdaWAuya
1rNeuVd++fX+vNxNyUFkBB0q9BEI4VvbVbLqqWfuMTCq0fBD7AxC4fIP85+/92qh
Q4oCfpMgtowtC4OnC9GmMJ1oyQmijmI4UOzQd2nxTDlA0QuBX+pSDbkQ63Upeu6n
/qrXTr3TYqk1fmPTZFZT/IU73gNXELqGCojdamMCkbNPzlBJbuAEGiaMpfW+dHQx
YbpAGTPjWVPOgrFjRlR8kXddy/3r6RrZ5LVCbmL9ens+YUoMnRYqBdUUy2qO6A4M
DYvzDCMgiSpsAUgMC2jIZZ2iwmDSWADgtppzgDxBhPEMBdHwQrvUtpHx5N2AQcCc
NRFshjhjpmTWTL44fSBDC2696+CxI4qgxuy2AazyjL4S87dv84gAMDQLBLNdkUnE
MsWZqfd9+rlXh3dt3jtm+osXDsSAuGhJED0y7je1tRIhVfGd9/gR1zbQds/JZIbD
ERr45+4seangMj5uuuSvhlS4AMp5AnCOM7zD+T2II/C5s4yoevGLFuxBuWc3PmFe
bx0OCyxBSLLyWeLyMIS/UfWdZUZMBM7RaCYVpFcnXHg9eq0EZuOl04SKOMQw36KX
NyZyj6L4z5mLcKG79oFLsWzpsAOQMDX8PtbDKZ4LqGMQHJyujCyhEbrEVsqAB3I8
VVxWwwv5DnjWDjOulOQSgYPs4JPcipumrS76kycQigNMCcLPpnZxD5+0Y8Meh32+
3PRDAK7BVrKqGaoXBrxvbl0vtmjXJJDBvxNB8GAypCb7gJVBCf21HeCjLYiMDlPy
WvnwY71n+2pNz+DWta3R9mqh0Q3Dos5t0eihNLZNmCFbkA5RBJjtPyF66ed/zdug
bJ/Nyg/sItOoYG1Fx6YfD+UcpaKQAHubhtQfFoXPSY/l5L3XgnF3xjurAabKJLEM
mg2wi7edLT4kIJTtTmY3+UL0vsW8z4StTxRoiuolqLEzBapagfuk6zuXMrJIaY9z
1tGD7ylyACWXuit2V1ykLHy48jdIiw+LTGEhhMQILiwhCkWMMAOKutyLGuuSSq80
8p8NNyD3+aqrbZn19c7jgW0+GRN4QIrrCnFGA5KVuCy6YV8wrlc1Z05IhEP+b/W/
fLx0FI5VG2RRzPBaiqF8SEBv3NapJHr+IGP6jn3SGeyGUE0XuDDuIO0XGm9M/pNV
xfJF2jnrvslnIov7f9MdZW2iM8xsKyqHTM0q0IbZ9GbicKLHl70R08E04258Gujz
IDUk/sIAyLv6ke6u4PZZbXF9382Q2lvyOIwEWV7xnMJHZVZMpdM8qNszYCQ9Zyf+
0ifHTjTvcE1EI1w+wK3YhXONvDu1flIGZoRk1X/7/zoSSC2ct++hz9ltTXuE5ker
ChxqbORUEKSynBX7OS91fbxsRMRjScBkN6ZRaZj3YtrV2230kvgHjhxiEWzWvToL
sA4PF7TfOwV4RyhpIWQjRQWZjLsJms+xFUeljNKsvy1jTTwn/WetHEN0rXF66sWD
Xz7Fmd0JON8yFFx8ptbR24/KJELajiJnfxrGeoftLg2+z4CCfZjOALjED36sQpt5
UGamypd7vqDIiby8gpMAgpwet3zgRphtm9MAhK3OtLHN4YyQFuF+nxGjTDGcss0S
HuAc8uLKwY2AWOa8Bgco9UuvHfIKAi6q55ElogKvgOoUEqNg0zmpWXKsMhcx0i/8
Lq2+Mk3lVKcGilGSuagLwv/8eurxkLvhOP5f+8XMj50gjaiG84x/8NwQeMtIZr9n
JVgyK16QKmsvag+/UdhIoKjHN4oEgWgEQ8jBJuwTL8iw04t+xynnPiSzQ1DACtN1
ROvljUi6zUHGoMI5luD7ZfUCUCFvIOcqo9aFVoG/ZQGCG8GnFhHGN7kawBiosddc
EOVzJi91jlXlyD2QZn9swKR6faEIIMot691vqn61APz17ZLjJm0nrGKPn8Bw2OKH
x4ma62OwI4U8EP6ZbTn2VO03vEAWjvkSMGae9DNnEn7jr/DbHwflWuKKl7BQlrqV
P6THsOMEfrJMFS2EgIz0WtBytOGTJDGEk+o5DsF1mNIeqgz4C4MktsvNHkjkKaA5
gFbF7Abb4pqKpQ8bIeGAJSLs+m9VPDBwmfEbHhIhSs0EVk/YWu7y654geP44qnQ2
Vi+DuEmPxQrKsBDZIosKbnSh6QJlyMbUoFslzsxRYyz3gIS15j18ujwrw5kVCs8t
O2QVnGZyAe/uJWx9DfjwRWekoUMQcbwqolvLZ/32CxUFopB7FLrPUyenIkK9LMj1
CvumQHXhdW5h9rW+1Bzs12yP3tO5YWp7NVN79w22vylTsjTReq5fSU1rt+4IGVGf
18jZ6mWpdg9ZhdotDUMq4SruxcW/nY/t+xwqGFyB7gLGS25I1moeouBr23cCL/SF
Jvkj0/8hRRr2h3Rj7WQvPtkn1v4DDVZkUySWmeHWBghZC96fyRg7+WGuq+jRdj73
LRe6KxibVBQxbChoomxcm0PwLfKax/b+dfFsXOcnqIsiK049aZd/r+55qVvWJ2Gb
f2jNRWLjYaqbAA4sVAnWmCWx+xKF1uELpQCyYvRK01sbggHTfYKRDtyV6DiFq0/K
XeUfluB5RVByEDsCuFVONzPZxC86OydbLQh2iYUkH8B8rB8AJj4yGoSaeAv+Bjep
9g0/FSe4zf4YSyHA7o6Zxsd6ZS8fzQaL163yDUUr5SVuf+gAKhISCeNmppPq93Tl
lrR9Lcob+skf6bFAGPYhVw/UcoxOit6v2+XhElPW+kHAtxvJrr8vh19d3QD8o+iJ
5ZS7xAqPOjPoPc6iyvwF/kkxlW2Glgy3E4cAMIqsS+fijebGYzzens7edDY+Rivp
jm/gKccHEuccnEnG1mhaYO15mXzxqkpYSh0gznNOIGGhExBe3iLGbD6Hb51++nFA
3r9riQrnIukMPA6PAnlPF6QHmCxYeeyBextTe+NAe1Blbp0TWTNdTKCj/YrlZ+EK
PrRJF6G/1a8F2RkwB719j0YTfznI5VgJ51Z3iC5eFkCtUo0Y7Mct5NxqKPbGRLgz
H5GxhdyiOYfyIuMm/uz71l1lrNAEXChko+STwmj3BQgv7Xpwto2sOABUttJgBiXZ
Gh8TE9D03qmLjs2GzhKKCqvUsYkstQeunyD5+ArUwZJ+8V26YVAfKi9XsCqgCU4D
QlWqUU4WH/hgom7uJ7lBNOLbKeUQ1ZFyBzROYiBrUv6aaYyQXw9Ka4e+LXOw1tNX
8iJdo2sBaLYa71r1qERWGzP2X8/MOlvzx5ihZZ2Z3Z72+Cdz1l+HBRxHrvIcSgWe
Y4clW3UNSmSYwBENHyhO23Z6/Xp2bFTkWnEeRelc1uk3OS3w0BMsIh/ElTBziPVC
aYOlR2BNsTNguDl5sow3VMO/p4GemYkKmvhFTUl8Tg91C/nwEXZP/vjdgjbAzJ4o
17dbriTEap222YuFR+pOsqZ3F4fLkrWtRq7fNpYU9UaDg9DH8SoZ2SvZfNZknyNG
70s6VLEL63EbmtUR7uWFElncczS6ngBcTvL13tUNNy36jXS8z9NQjBJ7MoCYg8tq
gFKycQ05w0WqJ26G0Y6qSgltL4Pil/VTm4VlqSz5wXaRypDCRMKKGtLxqwhgeYLs
qMbilns6dNudPUB9QQ5nI9TqVJeqbrLpcQkLFfccdUI3kbEkJ6LzKDKrtqcSamYW
hsYN6LLaPWZPLQEcNMPVnTSMZKxiwOcOS9AeP9bSbSFl5MoK4alsZfZM1oWnJH3f
YRmD0tQO+bpnkwPyWZnOUWCjt+7dsGkhXx8F0Jb9eDRdiKjHbUaQ7GD5fML5ji6j
TE8wJthZ4PZD278iYe3qOKNHitDSGCf6ShvlqM0VpXjbTJf0git+2kXCJUvv3Tpy
sWIjbrto968TcxwA711a9dm9c6hH60VUkCN2auiotIR1QzBHPTPX4qX83HgSkUXV
KMlyMUNlTY4xwFJxrKYB2JpmQkGLI7+Ou2nRorwSkdORN9IBLWUWA305cdspuZW0
iOF6+dim5iguoouPAp0cNTfG/dnTFmH+LK6r3cQMM7qOL3NqEDU/+/0S9FZAha83
8sqI57XT7OtpzCqdE/Opr0iXfR+CVuSTlCKh9HLUSMGBocxpxGsidLRWtUFTvMJ4
4MHBGvxLQxms4krIScruteYFidDBTANkQFTrqJgIlJ4JhRzweIBaLCHt5nfkaS+C
HAyBlCjUs/loxm5FnjCbaZ5xNCfHsQU4sF1EgF0vjoZxUK8UEypS8jQBtM57DfFZ
/PZEgv+BbGRALg2RtXPA1wUB9cLpafUnXqc69cpoa2CPkNSErHW4NEnxSmv4+3dT
hJ8xOI+7XPPKm7IopH5DAhGyKBc42rIQQLPe2/pzqurvNx5lTeXgjTTKxH7O0N7P
95b5imgJE/6gb3mS3O+nPfyeE+BlV7EeEWZfxgG4fXTPFj585d14NHhnLyaeQ+TC
uxUPO6ytCxBOEpGUjI9KVN999Hhea6Mm2uWhuwjXSLcXaJW46Q2fm6W8dVqdhS1r
EWgfYGGate2ExoCDS2Q/PPfJnO8dmG3rZ8Fw4m59eVYY1W1XIVWx4/BcrJsyRjBJ
gFpS8jGv/fUqcdowvv34EjbyTOcOjQRTEXBqYKueslQOV27MfRIUg/qlXSIb/Mvu
N3aE48uTpbbf3I+FVnnC+sGacAdkiTgw0Z35rQJRMZYSvGazycYb2SF8VKh18z2a
u0LCULST+RLlrEphCmtRGG15l3N4zy9ANHNN/prU5kiTvaqAhX2Is8weoqNBXDPw
+nx+QA3xOR4QB3fZszy0D/2ZlnMN2cFTknCvGskV1jcuTVR6DEhGcYn92ANpHhLP
Y8GdmPk60b6BdIEcrJUpwS8ldGOtUxmYIdGSLsVYJr12DayeqwLKbdxe4cuZi2wE
X8IQhFAOw7fGzMerYaOrZPN45EDcCLFnXLnpQBHTuWCIdSwGVgS7X97aoCn+ybKW
xCESr53pU/wdmkSvjIGNN5MXKwA6OTv88YbT20DJhiiEHmykGUAYtSfFgGdOE/BN
qlfcyBYrhQjVDClwL2pLQSJReCsypCYr89x3QWvQax6cuag4pn6Agd8g4QwCuzMT
fbOyftTodfi0Crbz8YmLToqdSfQVcFcQqrYW3R9lW9Hp0G5+CmswrHaVS8Housf7
bsV1XMugD2eMEskDUg9yFeGXVKXucEBkpiQf3ICNJt/eEaBLJdh+h+zBtol7PF0X
HUth9uEsV3MbgSA5eX4T8HvzWZRlNRpiLJnoxQP28L3UJGsP/x8v2XT7df1yyBOr
ro5oBfY3UCn6uL3zYq3WP+UXVcTGzwnTBtWAebbVlN6h3ioFTcr44UylgBH9xBx4
E8EVcnX+6ATZHerLMRmbM6yBcrGOHC9HJnoreIepcfHIhtYBs5FqQq61ctEszOxg
szwtNJ7hU+nFI4h6KVflK/pqEZVS0rsG3lMSYN0VAIdo/uJy5lOfgAmowj2ayJZr
kdZutjOxrq8dTsrAhRilV9qrITYMWkQ1gK+0kXzgu9Kn49H/jCKo7T7+CVwoPrBQ
EQXcCCpWUFoQJT/WiWsJaPEqtejoEnnySWhxB+GNlG0hJ5fXaRu8PY71c5SYefYd
FLq8ly7D8Gaui1A8juDv7gtUWpBraxM+X4RcyHgM3+zWJJbK27PE8njqQwlgljRi
PpVqbKrPQ33JU4vGkLZSe2L4dppR67QT4kPidZzkuCu/3NcHNwyO+DnWlIPcpAYE
9f95B/zcAPmH9gEg6KuyIqgvPIq2EsQmXzLXd1G5mdm3nQ8C9L4JKtSOECbbSfdC
WPylbQlr2CROn06/awABVXxApRo000SNyxsbsNjVnSoLa/ccYgqIEBKBTCwXs+8W
X0fUbpYvU7hdRkKtfGAICXTdqVJVVh5bHi8Q+Su3X4bs1LbM15WxLtWLznMTM1JY
+3E7Y4yw82wl8E6I7tHB0UCbggYAAPkf7DqjNMXNzXPwmx/4NXvnJuLBGHASgVQn
Zg8lB6q3RD46W+VrOo7ah43XJEz37b/9hA/8b7pTcNQrNBWrEJbt7WecsAILo60X
ch3J5s5t1hrcXbPHcIzW3Twrb0j9UIwyNyyqG5gNEARwuHbq/30y1CdHg1qv/zWU
NUPKOHNi0jIuaCeA5kH3YB54hY1/uadu3J2Xa6w0F+WtAnc4WZVdGKMiN1oH8jH4
5KX7MIaGtmnM0p6t7XUryUxCkjcHCICDC7+nU8SDxbAmKbT3Fwytz2YVpBenyi9x
C5lCcS8u4xEaDYdnDuynRCx3rJIDuO7yy0nSfRiJc3NsTy5xqtXqLWam9E1FgC3P
UN6KmLfTU7REqW8Hraas8oV7yo9QOq3JPuL+eaq1Eojz3UU98Uqi2ERADjq+gowu
IkBf9E668CDKz0EciY5rlqmXogA0LnmjD169RuGO3sCV3gYIYZ8HHjwthRhm14t7
ud5q67x5t0ASb8hHaxmHEjXupvdHxNWeqSvd9o5Ztbw+OfxP9bHN4bJa4C53pmaB
YUUalaaqqtk5/LzI8osLWL2HTpCTyRXmJjaSKJGbzqJn1lBBHygWNmx6YJNaanVa
3F/r2xbTiaRJRUSc39GOb/TfT6ZmhTOB/IK4zgA94dVTclxtV39nzdEnKmX5D02W
mv4VECvYFC11fC4hUpGstubgIMzNIshXZ6KX2m8CBUrHYVwgHxhlezLVbK1Xha3g
bQLabPsrW6ajol05W8hjDVf5CXKJP+dQhaNTuoRAhfZubZsYdlK8Jin6xU7Ps+dO
KRRg2/YdDeXsOceroz4w0LMy1oKzzZ5aPYIahuqcxR7g3XG/ocgcQeZlC2murlKF
gL0NPPTr53IQuXZZaVJsm4Xs7ZiWdy1p9yzaSK/sTlNixm7vhYq6Ht2Z5wpGff2z
SswATPUEYfQFVqspBzTVu5gONzrmgrMDgzLyJ91NVs0FET8HjBtHQT+sgDGIdanx
jrvpeMy1eoIVJfU4EzXHH1/SDMJmGS5wxgiy87uC1yJxyqXwmwrJzj/igt1SF7vy
PFo7DicJCk7m1WXq60UE4SMzyR4pVU6E1Z7awm9jc3WQAz3yfLaegXGM8slx+L0D
w3uRk8zXxBt+dV6nAi34rVDSMkkC9F8lWiaDZUiHGyF8h5353VTZkjQmmzaYzCMe
7mwLUNtcpN6n/6bi+77UYJt+eCvHvauIAISVV8JbDqgb5BjCI3EAAxV2sgya5XjK
w3QHVQcadzrVnD4p279VNxU7v3xd/3r2V9hCXjI2fz3efMrgkZUXEHfabNuweXl4
S29le/+i92kbfER9KTe4+iODs/Gb5J77E0+5L/o4+xFOV5UYr916InNQuofya96O
2vhZ+UNjOvQQaH7/zM+ls+/E7dZe7TAhv6iMVCw2IMrebGoSdGvB0MZBJ9vTcFi/
4Ww06JCpJSrz3eBFzRC6AHMMjjC+PNHQjHPDHByIH72obbEnCGVS5tnxepDHvhbh
O5h0TTZ81eWVULnR6u3J1752suldjb9TAKPT3gJAWEaAGz9VT0jPWwQLlP4aglIt
2Z5OmQEUlxVCOY2bjEOlR5pkLlLyT6XHEgi7klyH61/yosOwF6u4jV2S5Gpv+G+e
5ZdrSJrvllCrUWA3t/z9KdJFD4fxp9Ksqvx+bGmV3jK4fKJK7yve7/dpoPEHO/Vp
Tf4zhmjiA+llwat2PrnIvWNi81kbJPQ6QWJf+v+VIqRVTwt7caaM7yTre+5hLc1P
owOZ8CFc9shdXzK4JkgG14aS00LEriU+ndx7ZDyOCuu+czjh3YMCL/IvEiJhOMn5
BobCSrIDI++sasI+bBHYCuI9itlOPRe9nfQ7Ts8E9xlsWbrGzTjMkiL8U55BorJ2
7MxfRj0sjbAt3gYUHACfRdbkpnWRPHCxugsP6EMFlCvx+k/dv4mTD8aCh2h0HEeW
/feHq69ZdU3lueUujaoDtxquQDUKn/SmreIrLOgSNNCvyq2upuDnMVC9zrk5bED9
54GB//+2o7uglNk6jXGnmMG8jL3bcWnGT7gKOHfr3jhLhx8fyQq7D4+0sTcpE66l
VqlFfHAd1Sq0+cz8waftcIJttrKULbI1G1IAxfGYXBV68z1Mz9MErgQcV0QwWznm
6AKn1WtsbwVzbwDFoTuT+eiiDuF3dB0aukYd02btd/3cvxSC0P7Wy5AQN2q0hfVR
9fGLjU9lHb9S9SVjjT/tCS75S7m4y//bTDPHKqN7KJqaHheHnvSaR6j4lW3EW2zI
kZJfstgnCF2AnwKjpkYlkWj39F+BLcJmu2Hh37x4nDFa3SaETtPBVmACQHfllGQ+
wmL1mvonO9MyCCAY29zk6+tI8r5IoBsMa072TsDvTKsrPykD9wVHinEn1syHgPHU
jHQicVoXYCCa1D7q18Z+9mE6R5qn322oJQDMFTet85Va4D9QKpU0J5/eekSiYFZ0
zDWc4q3MybXNLoSjFtdRuYV4Dfj491+cxLwazlyhADhCAIMngnfa6gQ2JTCQEXxl
is599K7XQ1m2FpqOkm03aqdPXLeFIR8uxiyNBrA3u6qqqQlWfaSRGsmah//6khrY
qXnhCFTRxurDFnCZMRH7FEGZ8FnxU/xcxH6qB/GMPuo1kYZXvJXsvskJba5PM01O
+gDYjUypNKjorYcP43rvjC1mMspAcbPNRyl2YkJDwIPoLGyz6kQrBh4d3odGXuW7
S+P/PDEZ6qSwSCxObaNm0kZAIynfwu2Z6v1dDMCQ46a0rMfiBKr64nhN3ETTAhv0
8UaUTHmqU9G3lK1/p5oNw1Bj3AYZRH8o48v0AJRpqi7OIYmgI94KD8wgm8u9aIaV
BtuiPQAX+Nye2zlPyAroDEpyG9v7ERwEuEkg3ulFwm32SfW0/RK4CwV24J2oAW7w
+OLD8m2kprTpNu6AlJgAU/uPcfhNsJ+ELi1fPlQDCNwhcISMU8zW4TdrNMb3kN4S
vPDWGUwaE391hcbimtzZYpsLqpdzVD3L4kvrs/Qq0rmY4PuvmlTVOGOyhyilr4cF
Rb8T/oj5v0wGuZXoJZb2HGwbAMU1MblBwjsbYwzToAH4ptmDJ8ZIAjD6mL69DkAM
/WYPrUc51PTeHqEjwmknqrPpaUELhlM1OTKIksraDhKrRQwnBqhfMgZK7u2iZKDa
QMJMLSUEK6MhDQEqisdMXnRctq5FZRQzpw+l2xHsFyE1NFnhkEuasiC08b4XCxZt
uVZB+H+ruKNnf9PF5IIcSmyH1hKcd0TMYj1eK4bWAE3ozawWPLJAuKJh2jf+2Sti
doL7QPyCrBTCUxFugdVnh4K3lcaBUh/eubjYmM0XgBCO12a+jK3GYWGnbOvfa3he
V3QcIRW/KJmuHc6ifkLWiQCGlSayzVwj7y9J7e0C+UooR0+S186h69hxRkIEz270
2KUlno/r/FkY01/p2F86Migpfik3l1k3E+Fr6ej6+HbIb1PWzM6gQlLqHU69mvw2
scVPxJSd2iU/A7u1TWFN/BLPMidmw85upj4fwR0FgxusLWk2Kn9ws2KrsOoFn2RL
gwy5YKkHFR38Q2dzTMrepGcCWZzuDEaO0dwDE010N6nuja8CK04HMUhgnV4Z6aVv
45gxLx8Wm0/D4xT0K6bqKDBex+eTE2Xad6Ep5CxAQ9ImYMNYgmOVpf3B+5A39b/V
ePGSLJYYRD5Ipma+sgMOJN7wAtRaWkhrue6tQJqp+sU2bveckHs7ku4g4EETqCvh
hH39GhboPjp4ujX8vo2xWjSm0pZTnwaSnyDzz196BW44q11qgHf5HMaUM4M02zB7
mnNpTH4k1U076u6UOWXPsC6tXpzcTW4KH4ZOQmK5iCp7IurUWsUB7SaZlv/d2zJL
9s7JTneyY/EVf3HRdsZxsKVT/bpY/7t3Cfs3F2Mua0rg6XX8llnMQMoc+h0FJTly
ou1Io2jxFK6Uus/nMEGOX9ZTq1LefK3xBDN2tQ0wGS1WybUjfQSCWS6hVi4/yhT1
V5zcTdhr62ffKRLVdtdwpqz6lQYWxxgYjK3qzLUfF5vMS4h/DvTxGgDtD8FuzCj1
CLSF1y29fuLCtLc4Oty9+6vBWKeELaoZNePjbZ1u8RJw4eazxJFq2m2Kx33JSLVX
mwCy6ed7KBJKusMkI27vIuD7jn7r13HDUyCRFMD8hxSlZVa7UFEt5z8B0q9twhLB
exqigggAXW7Ho/0fhLArPuGmW/yQQmREui60HCGYZQq6KLiQHij9y8/l8jYKpZIy
j0RmZmIow2sNDd0MW2I+WFyLooYDor8nrf97ySp2BR9strmH7+quHaMi1Jv44Fan
/Ck40trskKK4FVX8zwbmwmtgAosIDgX87rI3GQqsF+c/rbkmw69tZujGBh0o2lsY
SUqonCdxVmyfWHK4ndXYZUVt7z1MDj6fM9c8x540Hd+6kvYgvUAchKAyWuARpyNU
9qxD/uqn/LR4YdON2LlRr3rSGhOhAum3dsu8cY3+xSACpyNHNZw4C4xjXf8cXyfY
JIFz+de1s/4VI7YXHCfP95iiEGEPgC1Hvijf27D1EMibo2zoyJbT/PEG8CokvNaM
VnGDsj10h8yXFcCgtV6C3+zcz9qkylAwON9vbFg0H8G8tUs/W93sN9ih6C/uXwX0
ibPiV8OaZqCePOYlMpz0H+TqHzYJwt8VDjy5vsN9yz0hO0W3Br3TRi7T9nBHmlzx
bJeiMTsZeBYpymli3C+sMPODS8txgaQtDHUj45E2amYPhFR/t0ZzcyNELl+gVZSV
jjtrlp9H7+IUJZ+UzLAw0tMkHB6kcOaJfZ6M2LYJuQXtKmCUHWc5LUzdKkBasBvR
I3Vy4n6vg3SqQZ7V66dwINlzC9uqhcbLPKSCsBP+t5ExelTvaBHyRPSUJPKeizZN
XIrhu2ga88dGxQkrv0HaILPnKG9ALXujY+ees+nTl/eiT4EaCvMsksagDVPx5D5V
f6Y1fMGI/0Wsp68PNw6mk7eQaZFgmHS1ZWoA9JuvopITBit/KSnNutyDmUh+XQTw
Ry9RJXdhev1IbFuLdzrpR203pgl8le6m5dSmCxTygPem5RUhWf2P0wBbKbts34qL
sN5Ez5zkr59UPT0JZxIMCthkqg+PJR/4WhEe9sP7eqdExJH7fHAouzloPvtTguwh
LIr6s9ibW9Gyw+yNJyN1LLpSScokZ81Tc3i1P6bi0u2iPZKfMAF3XWc9OIUueoFk
fZGDTDyvZLANilElyTXAiLWRe1otkg+BcXJs9FD6qjQVV72+Ge6KLKJtewUEL9fD
dgesrYgfHcGawkWL4rGux6PcC7GUQ8rGMynkAblTEVqoQLh0PtizhwKk7tZiNM6m
JsKsehqZ3OVTnDagoxFfwpuOnHJRFfV3VAH7i471dgfbemzWMG5A2/hU/03SDXoC
8TtiY3OQObBsimCSt6VePdmFHaHs6hrgy7b9jdQ5HCdNemLbAMYVIpmf7gVK2fZg
S5O3zwztKqCNj+WFW6FDw80HO0IXq+PH/whAFBbuO7B+19K9wqtKVwTsym61pGl2
lh1vFbRy9HGKlkGqRAKSHQAdXFRYEJ4zWHunGLxCTWW7PpEf8XC4oAlfNKKsF35y
/CtiKUW4i5wdnegbtUprj4j+bEcUe0LW3pjmAA4dyd6rRB7SUaQfRk0tBNOIqGKm
uvQ+G3Yb1rHU+Ycs0Oa17UvlGRQ9PdBh1Z+8fpDgh0z531dlkV6DRi5Ou49RHtob
crR3+eyTfvIK/n/n1PX8UlH2kNALRqTw6qI0/8NqPaBjBWe41PAa+FQB8FWXNfTI
8eMIb2LSLtPSG1Dii3Ots5QI3kQxIEsvfI/um7dsyR+EB8QneXvivZHsJ9d68LME
+PKa2TXR3yyBPTNZ2evNbNuAN306MK8+HNHAWHG1CU8FwZpxW4XPMMpfa4cOA37i
r41vkTpblKv1TZO9rgGNisL5sGaSbLkj48nVhIf+kIjkZDieFFhqEMH4dq3WkPPE
VvSjoHR33ckp8toa+z04SGdxhq4uNgFvcsvuU8zp0SXn5AyB/uloqlVCkYIwztg/
m6hSqJcOsvBTOFLI/RC1weAwLkMnT8lXVb9CWc/62GdlsNSYzU4gjFWWkNgz2G5j
onjaT+E7D/l/xAXhXOMaCYbk1SsGq7jDoCeI/55pGDB6/q069eGixun2UrLjB1uP
tMSV0I0gnH7Zu3GYtr+DWjlROaQ6mc9Bjtva+PQ6BfyNSu64dB67iczkcsS7FzRr
zdkd7Bl6wHvlaEQIebzEr+ATecD1AY2q2bD7ieVgGjS3KaaYkN3tbjsbnzjz8MMF
dvZCVYpFJlZrONVgsle6LTGXjTgy13fFzCofLmhsQEQRF/uwbyy2XoWt7zzJM7RE
2+pdbIv4yI3JyE5zPWOMKdWenTLlB0HfKHmFbZ2TRKIPvckKiTN+koYqG8wfa1Cf
U3WejSDrMJtCsM68QirRPMorGkE/3JBoePl4hmGwhWM99QzmWXZL0H819YQqKwVF
NHi73MWKlmBZZybWgD3DZC+KqTeyPK6aJMNV3ChLbvaBuUTje+S8+UqfpkoBC6g8
qPr1LKFlKxwkyqCJtfJ/yu17zTgQy/NbCJDWmHTuPc6xGMcI6URPKMQ9a/1Njbwz
XfsGsxzT+bZi3Wg+w+hTVWJ2Ifs23QCMf0aT4z5sVWiEUIIui05iHpWWdX/3qA3S
xIsdceTAIVUcuZV6htbfeVS4bYTdxUluHA+2u11RIFqwXWMOFUVzZpVglyekShaa
L0N/0v0dkkrMpAiPfCRQIyxGoFn1IgA6K0WRv8eHD5Sl+SHysOOU+qFp55sAw3du
2ILlcI0TnHEtIj5KWgDa+yRrfqoJjyiHe3HkAZXvDz7Eyu5Vht5I6aW5Kbtb+b3e
4VrHaj0rOkEBuozgBV3Gurp3Ruxcp5Lc8Jz49yeXocyBRdj1itZcrivWRZOsRQJN
BWldUN3iUj1GZ+oEbiXqZInux12JWd8W3o6luRyO3WumR7LyGQX9/SB+k/xpFbes
86dTmhJ9JhjIjsN9vkeOdrk0uql6R/IDpnq3iwFCZEHFtAJrhYtdsecot9r3iKlA
vpJbfU6NwORkMkOowm9Sw+9iy1GFk3VA55bKWpiw1/OOnfKL5TPcvE2/y7uL8Scu
nrpxUUU/Y0Nk+jOt9OY9kWU7SBcZQj288NMV1VfV07ZvUvwTOjZFJvUOEWUjlP73
NJOqAVfbhoJVphdBFu6KQVGJ3Lf7+EE4M0WFV8rbfPfiqGbcNlOlV8wl0G0A7zdp
P8JeKqNZlZNGIXDczzMbNNRy8P87qiHetdUnnc9enCxxtwLeUBXHbLWtGiK03sW/
D4rw2gjWDAP+Ml01CPHCKoV0PsP4w4N6p/kSvDKKmiDMI9Hj3OVWJgsQOCCSZSZF
/Eto7WLJZ9mlzaAGyyp6DHsaLtLPrbUHqfpb+euZQwLYS8J+mcyIvedAwrpA3CSh
vyhxxoZEwauRROxL+5sKuPIftlVo1X/DuwcLH04Abu/nLp4eC7FbLM5rk9KBeGrn
s4v4WnuJp4v3/nW0B8BqgkQnsxj9xXdTQnfEQXJMpgBnMK1B7N7OUOmEDtza13Bx
y0fXWwjbSSC3S53ZlFsz+g5pbZelhT4up4p7c/lHJ7AEf97bqBk9Z6NZyYp2qfzO
dGvu0Rb/rsgCNJYF0S5ylPLX7EKL9yZ1XTNIgjcIpTlTEDuBq4X9+4mgq+j0KZMO
C3OIveZC3gqDkIgxtHHs2qWvX+7H+k08T1V+7nuvW+FolRyBvircPZ/ko+1uWEGd
2Bva/DfAFbfsHv/n5El7hoA1xz1+cMhzF524JfwJ1A0NfGnuW2DAlMQP5DHetUja
4xGLEBbm+wk5bIjHGH2g48h6ioMykcgWNVJLiY4+pWRMXiJLdMQ3kBwyxj4flumz
N9uNVESKGbB106oCEdhkbtcWpygRwz2zZ/oeL9g54cvK8Jv6+9bz09m9YaFrcy0p
9PmRO+XKyAujgTaC29t6PPZzDbhEMZsl1e9+mQ/VjCG6ssQmBl4HYfnukjok6N+g
V9XX/pRk7eDRR8C1pOcsWZ4e0cMS95pi5WcBWl9I8Ktg89IQa8ds01/9b1PYTxma
wvLbKXdJcElcYVTFKqcyddur2Jc1RWwg3D8gTNjrX2NYzyBdUvxsi+V/Tawq4zav
3tCdlHZJJgR5hYnbsRrxb3e0kQ5WNBTBqaT+AFjYefQE0MkGiZmxYHXfoyUfo+3v
BERk6TlywPqi6XKHK3svWySHTBqJ/LftRFI8H6TfgG/xhU8s2IiRIyE2iJucIGr8
zPODcJWjc5X7huYqKZsmgDgq63N/sVtYskIZIVghGzn0Wt077AfUVvaw8iDCcvbt
QOS39dbL+Tl8wTFe+snbTevGqt44FT+yF1v0ZSN1Sq0caZxZtc31JW6acm+O5jcO
s0hdKFo6LzLJ/dMpCzPcEu55KukF7/IHiA+QQBMXVmX7hdv3bwpooH4gaYxZPuj4
uhssKVU5F2j3u+lZxiHhE8j5/kDWo9wa0FF7gIUA6CqMZx1QSE7yMObllTrBCKIQ
nd1FYKsZEDgLEk9exEG6hWM3xfUxlpXg1k5MOOpFsASRabFe0KAq2TEnlJWxH1er
beJ6h+FMZMfkSYwqRTvCBzdlpqtTi3REO7ilvmu3QGu7AEDL228mPufqbhm69SfP
1XXfNk6wAILCN78AbXm2S1nGkicfP2BCdh2dhcUlnfxH/aXbBlU/s6YW5u0md2UX
T9fAfYz9WBvrqF4uzcqvUDSAFg/hCf1uQHibaFqPqnHPDKmBVC6ySxRjiANuiEjj
hYfnNLO6zyUntNLOo4XTxdb/SOXnEYMK/EsnR/Zzgh+TS9dOPGzw+zQgUm/zKpQx
ghxCiT1aHDu1kp2m24R0xveL78ZwUwc3bBGGD5X1xIKfC5zw5RPSPSdmzwo8begR
5vtdATU1oUPccS2WbUlOo7aUC+k2Wc+jYgzmH3mOxFPwUyJ7VMIsxWUmRGGnzMqD
8BcwDaGhdVvrDIR8YXQH3mpu2dzblM+ATEu0hSfUx8ZZ/mrOxGSMS/lMhpiJsU4r
w6Ptc0EEnrEt20oDBUZSdMdQd0Z5R8VsotP61YKzpRgY2OEcAznjN27JOqImjgRT
7fgHFUs2XCLtwB32ADZgTyxuAieIh5heXXxC1wXrTnwQTqLoE3BT6VypZ0ClRTnu
X144GoriR0t3DpiU1+YUvTORUqQeQXXnuAh3Zgt6Kt7Ux09RkC6PKKiruc+q/wRv
HmFXD9SWznM+QNKh9I4NJ+9ymM4zxhMsxmM5FXFy/wN/tutBd1OadIwTifEQfiyA
eDZ9OU/NxYWwbg8UWrnJ44Yn03qi8SmQ7+6aJQSCErguJOBXvEyN6ZAE96jFFX62
9MT2gCHqJmNt9qfgwERM7kWwiEl74qZWzpXtUosqj69e1C6v2fmNGJJKNmAkZP/k
BrWbDs5TGS2xvM3d0fL678EGCVjjESb2DY1GkE14JlpYWdDCb6rLek0JNn2EPLSe
PSfWVZg7fTpOzH5d+vIGRhBlWZQVu0HDBz/V/ENVVVCYxldMW4GEwFldkYz6yw/r
aKE5wHFufUbH4eg9eoRZtsJWaanjYzD38ey6dYmCd5kZq1csilBOer3M3sjOQ1d5
bOvBZ/8I4aIh4A8XSS+YnvK235G0DgWbElqX0TSUsZpR3ye4iWGLHaebAnGUvIS6
ExIDOFtra4ihe4kOV+QlRyRu68U6t+dVgfHOfYZ5jB/fzcCidOpW1gLI0Fly5dKU
8wRvL+iuh0lKvb0v5yQZ2XOMj2HmxN3ftMwvvgDtK55dP+fVbg1P0edXIxLvl1tO
71fEa3aVQrWc9TVayZHQDrmGMOLtj5rY3ayeUPq5a5yiNyeQFQG+Pa75ami8aHUT
9QPfFXxF9Kr78Wi0clvOCEGJ57XBJOszpmHnP8UmyyuOjcCUcrn3uG4L3hB6ZAy7
3xLM2jPttnuDlXygK4ur6oq+hW2QIFSAv0hizno6Y7hSIpRY4Omt2ZEcrwfcRT8I
HAUTb+DcehJGsvo8o3PGrGjFkpswMyVyW1wL2/hoXBEb9t1ycJ1vNohgGSb3agiy
MY/JmpQIutqIsFZeSFrArbYg5E6ILn0alO7mLNsIHSP8tKc1oWcWduc46M+RxGXc
mf+RgOainbws07h4uPrNVX/2OAJWWdbulKBtQZ5baaBQg73k8gD+XQftWrtXv76r
iGfwC0ooAu9Dz8CKBbyHqW0anu9FQS8TiKDX2zNXl8fF+O1yAhv7BwrJa8QIMVLN
l54rO86U9GtCa3y9UYnC/BzS8q3fbBcZIlYwT179AAXqxQfb/0Cr1mtFzXSx6gLN
YfrSbfukVWXf0XB0M9TohILKhsULylRDS6vht9A7LJbuOTs6QjK9Wb9ac/2CTrK+
Zkva7sdVJHH7Xj7fNZ8uRI7PV8jtFKwCLJGRFr2SBBgg93+9uuQEQzD0RX05QnUn
WdkgKV7LT2V6hv4uVPIg6BXG3dCKzdg62H9zIyCovpNPUCxZpVirkcaQe001YmSc
IoWpku+vfVVcxtpWWdkJGjhh00/gbuhhXwgFXHpFOAqQr8s7+zTyKzGZL7odfvf6
yS90hQljLrXqlq5z+VTsCLR/JQVoDPpuL48C4NsLbAJRgpq+22gsOPQYZuXB0bNI
4wjK7AT7qvnxtZiks4nJ+VHNF/hgcbC8hbQ0KjqOjzSoegoeP6Hf3m+OQdJ7Uje0
7iCywpthETJwWOtb/F0n5jszemO3BalJGApBxGXVnjn+6TSDXVzGN4POSg2BoH1Q
LXgmCkIjgKTc2ctsrUyJ+KvubjqGBTS7NRCCjhB0zOYpZzFUhiX6AFECuFoCaYUm
FMdFUJqNrg9Chj/P9z5mb2IhKeuUFSmic+x1/iCIUUrC4hwVODd2YqGPTmNJcB1F
TqRV2BflxFlcnvIEid1dKoLBUsZKsHhrCYAkih1M0LrB7D1E6eVhHbF7aW+DwL4z
P/u6h9zfMyJmhSTnSIKwQXMSjeYPLYdyGbh5vSKT4GfdQZTTGQwUolvWIg/IF2ZP
HCzZggNb7dttqofmOnLF03/slRRGnMlZIZXxlXIovMSULDMIEAsFDpSY7HY2fsCu
72dUhv5WrwJjLYO89QFeWKYoHusO9dB9vQwMEFtsP4jhLfIV63g+qOFRKmw0UmN1
e0+RANWd1Y4voji+GYSbmjH3AS8LyfCEYkzaanYuU6ozffrhTitK1eZCDNyzq9xD
Ss7lBJRXmqUdpjD+xpzgZf2l9Upjs/azOxm+zUXP5v75MRwL+9uzG+/Wy7JVShIU
iRJYNileAF7wdxAAQ98Kw6n13/rcwwviMHlp9XnFVx4q9z/dHPLuApmVD7k2ig6Y
6zr5q4uwTsUAiOaOAovR0tpJ1n0ZfV7Z4bHMw3zAqG3typ+Fx3YbrIcKbqM5V9Ny
TOyK+J1SL2cSKS/rzAu/F6o8d70X7a74JoefYY/OcExZwW9Y09FyE/NgkGWVNRLD
dLp9jGKMIourJZF9LzD+LtnzYD58q7ERh6EeFsQKCx7rV/veE0LIyN5vvirMTyeu
5RREQAiC0+ElM5PxfhkdiGVMM5acjTTfrI4xFlHaKum4yC374cEmIejJZYc41uUf
ed8YOP7rAvKY255i+s0mmE3TpywL/h/niVKExKKtlLE3r0DL++MJ2viA3wt1RpG+
48a6UclRKqQ5K6E7YlneO7arijCv42hP7MBOkFfYq3Kv8MGXXIlSTK1ruDzO6d6F
igOLpQ2Vw1DSS6mKp8SO5xN1xc5G04/m5eHowg7uWKkQuOKEjjtq3iXHhTr2+Kp3
dYBHr5OIrkOAJzvl5DUhVStfAv0go59VBTtfQtLtMvT34t8YcYTSp0DxZ4J2UK7C
Bf79MyjEe4LkSvKfQPSg0BjMQIede0Z1dTzFICI2jocSi2TpAmMxjbcJn4flD/2N
scS8h6pL0yK4ggd5zF3uZWJyaCRngZHuxFuJNS6tySObdx9o7EuYQkDz81Rte/Dy
+gJe68Vz+GniyjqJTEFtC1Jbz/vz17NSnvcaa07ouMUMMTRU5Nkw1YE/AnAo3RLt
8K2Gio57R+I78LWRMuvWaIOpKPx5JIi06ZgzX8YW2me2JQTsHk2iFboEPLqqQ5ih
LOO+Ky+pLB2DCqS8zVe8RoVBk4pozErVuIysNIv40l/aPCuRMMVcAV8uzJCZNrEB
4RM2Dv1nxVRg2bxb6yp+8PAW1GGdPaPACWlLyoxPmhIqxNzm6oLZfJaKl4g8G6qE
EPaXcwhnybxxsRSwXfRLKYAaQvFjwZ/MQLMVKtyd43P+koRZ1iNFd0ELrz/KNj5P
PHcGgphnYn1u98XfXhgQJPtN35nPqJFBQR3khOlO4JadffFt3Wq8w3qD7wzsiNPl
TvhQnUfOr+ZxWmAE2AsawRflzxLMPT/M2WFuaa3Whi95m6J3d0rrkOr45DNP+tPP
YZSw/W2D9V9ByoOFRQhe9561ssTEid1Kt/sti4FFhGtLlls+UCPWpt30mLXXpz+p
eQKkXbI3ZsumyRLWWGylOEtHEFGZo7a0s/4AP/EJdvl4jn/cvliaYs/rorLp+8ep
e8jaJaGo2ZpRjwPL95Gky5pMokokRWxMkjQhe9Yfyrvk/RLk00ljPadK0Pioeltt
52jqMgwhOzQmkaPPs8d64tgbriiRX8O7kf0B8NccdC504tpLc9KRDGmS3iSsz8xi
Ntg5bsLwoXXvHV2jmythZGGKxwI74/+CfvzSpZxj3PdWhzuUFQ1p0iKh3xk4uLbd
Vd00DKbuadoURPbyokgNhW8JMgYtiNfnW1Slhf5BPMUB2fA7zk9d1L6VwJE58Z8m
mn6GidJA7fiw9oPt6auqni6QvnQ78ejT5DKFcAFcTZMacSlV+GAx5vuzHQM00Zp+
piZPrxgPnfVB0+HZ59hMdOpz34LX40OVwIiiBm+e3SD2lnt+voHQxM4RJsLYQnhL
L2uE+YwCoAPJ0Ouextt1zRs/XW6yOTS2nHDGSkaxh9Xj/wOrkHAVZ1ZXOqpUz3kE
9ApStv52tdwoVBd0Im2w49z3+RERno/7751H2GwX3iYeoHpJxkumM+SllPSSmADV
1NgAwhOB+u9eRQVEU6LfTCVSV/MEGk2pDwirxdMDbF9ChcJboi/6yEIIH5qpLRcw
LyDpk9Bv9Y4I6xqIA4E+pEvhwkghUSFlA9tcqG2PCUPkVeoC3dLY5eOg2ytoBscO
x812RI7mHqdhWvNVeUQD6z3MvDE6CyflLbUXqtOrj4tUp2o8Wj1k8xQr6hduOCz+
0rnaNeydzjJWPaLTZt0KuspRabIqzLmFQDC4Xg7aJUOa29K45jS7+BXo2F/ld4T4
JnLGP4yYSGGa9cY+LM9uN0VgOhossH91gUogETOQxeJ+YFQ97/DnDazK6S1DI+Qd
oIJJn+73BASx2nZ3XVPgXJr5N/+caGcEVM5eMi2oEoAlw8z0N/72AxKgSuir8Em2
G9tYVx6P0yx0QpP6gWg8nXe33zyH5StR3jIlch7qqW93hl0BQN+Gh1xWfcXWPmQ5
c4XR/3v44X+CdOR4vTaKKCWkO14sdFaXKC3x5QrBylP+ejgY9Uc9EOmg1lDPe4nT
gwz+9nwXD451XQ9H1xjXlgnN3n77nzcxv/XvaZu7UcGLQin097+oNfD6nmAqFFwn
FiA5Ue80P8zsLLDNrBgcaZ23ta2Tn0ssI7DTCDuDIrplE6p+beP1fdezKez+e43M
vJjvESWYmupZ5LZ1ER0M1Twy3B7DA6hGfiMtCfqt3eJXOK74Ne+qlTEUkxla+hdz
g/42LdZ1yUKBZfzINI2fhSIo9gFv8BQKewZagTSWALqRhKsXTOX85+N8c5Te4IRe
g1gZ57rHXzPgUh0ROFqWA8NyaS0RvYdtLhL/ebRwZtk8+BoDXGn7vOJd/FDxT/zb
bsOq9ZZDJoCfGCKorh6BY1Z+DP6NETpMFikeQszw6JqU55HTBCrjbKVqQTXPt+T0
n/lgxACC5Cj2x94Vt9GLJCmc09NanRDXmDBtlyk0Y93Q/CHSNB0T+AT/1nhzFNiH
g7B3gKeKwyDNSFMSrw6zlZRm0jR4aMbc10mKgXSfwc5Q9Jb708KKd6DYsHYNZCJf
DM3VcRk4eHczgdmcDuKd25rpZAfjcYP26wWCdhdIfzPaMsHKr0p8uKUqgZtmS121
xmhHuDsO1cr9iTR2hTV9ODCVoLwuFDgs1MQUE+G47cyemxUEZw15lyL2XDHV1a1S
Eeqp27RZ1q5eJ5lrMKwaM32kLxIXTigDNkzUkO3j8g+EpHpZA6tr2cPLoeH7XB+0
4vK24CMob9lNZwu+VfhnlvPg/DGzEj7NVwc52Aoy/48QieieY0kv4VySKCJUGesJ
+iBCH9BihgQn4Cl6SH61ew==
`pragma protect end_protected
