// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
gdfMwvVyJBX7Dc0g2aJRTtSj1M7r0tiwCyVvAe2u5m3GLCSVo1HhNPWuZ8JmDOSZ
QTKrzhYAtQ0hBYvHHsOqyTpysOId/vWtH33FQA02XInLq9cIz7RwRq3g/hLsOLJ8
khV4FKJ6xrbyJu1+4bdYhnieR7n79miButpK3oAMMUXlHtpNZDK8qQ==
//pragma protect end_key_block
//pragma protect digest_block
7Em8vDLOwvcggvgdElxCbcFffzg=
//pragma protect end_digest_block
//pragma protect data_block
lkBT4FgLW6wqguxdSXltc6MN5WqyUV4ph2QqGga263sR1AVtRIj2CltiSCuBOzZ/
W0QZd+StJavAZ7MvsxNwnJZdm1guDibkrnE8IrU6dz844gj/pC3cVwA1DWiwq/xW
5PyXDfNY8RLTux5puh39XXywmzTWmpYoXONjX+BKj7Mdvv+qO1BBBnCddina8N9t
Zne0VbVIrH8FibESRmyQT2tz8slFEdz36ENvTdDJlwHI1KScoY25LsHmDX+wf0Er
RwO+YssXFuiTKcWsIdCGgsCYONRvD8ZCNOSzkZMCKBN8hO22VHxfHhSCYNMb3p+g
CcenyENOVq4mDi1zmt8QrX982x3vVpq0SD8W18JIPRtYLymlVgNHhWW4+bX4X6wK
p7J9Z1k+KaykflF7EVKtjFJE21z7Cv81JAbIdhaB4CBZsWsFaWXsX209vPUZuZfR
yaFcuaEGls7L7h7Ukd4fcCZypXPTm9dJUE/nJr9HU4jfbdpuRAjqS4K5w+VJIK7r
n1LSkLDCUglqZsE0ov9uT/QmBH6AZ9djaBBZdnOE8PZuVLCSaguGq867k1LfnnWK
ukJsHkHzIC6GJmJ90WqccqtzpYl9q8FJdM9v8omz5x+zUOYmRq7jrJcmO50ZsgcB
oJOL8zvzadMKasysSH4rxyVeX+prEcTGVhfitiJMWV2vAvV1+x0ntTioPU/cSnYS
452mAhi/c3pTWrPw1kO+cTErVogdsZVLoJcSn8s/14BGPNBKtRtJWmFvB7Y/2B7Q
kFBmSgNur2UGVZw6++J/9+WDUQivN7BSun4RIh6leXokoA47nVXvRLTvwm+A0UJf
iH+A56Flo9SK0MSs+IBNU5l1flqoLpUqIh1Y4J+qSFk5Itn6z8dKItuwZgP2smbQ
cNicfTXFpKIhFhmiaMheBWIgyq7cCTkeaXthJIl2F55yJRwzsJEafSCtM3yhevBQ
DDes3/QZM3VrK7MaTwwvQM3DXV9bbNEiM5nH3ln/JYDyM+wqMv/B9EpbOymVgJe8
ORsJbvguSo04yX2EFzy6B9dbM6ODpa9mMAPKf0AOtLqTH2rHqn4tLLy91Dw1BSr+
O9Z11vwF8VyylQtwh4mmSzpRTjeeAmpXlEBVsWuUtyUl6kGBmczv7tIoqjpvKs/Q
echGhAh3Wuv0BXukfIFtNdIPryuOkIL0kqLVDfq0WtWDI6ifSjWTFPrbd3oq1XDA
yybi+iVnpfPOHCuAaiTyy0vNO5/RKp4+iHu9EmYLf8iP/dRbJVHHjcCiF+kEbzls
m4OXrVdOM0DG5m/57p+Df9zDtQjEuQkPKl2bEI10Jhwi3O5c81s7XmKSwqbiPdCf
sxzt0oTLW+q7UD9VCliE018Svm/2glIcMs4jUkTclxInz2zeQOfSOmbLoHjop3Z4
coxhiSj6u7NN3ZNhTcLgjxZMYjpJCGe/A5W1bS6Ylp0LirHmif563Jr1cpHFknGT
8je6M2hwO0EBWhP5ImBlm/e1LY4v/GHDAL/fd8PDybhkDtTFDH4E61w5NUODVj74
u6HvzYn4XAL5Nrdh7f7CObWORnvik5kvfnCVn8D8magKPzR8MBrXuTgEoF/j2y8Q
qLRCpZnKv8XUISm2dPz5srQSShsAe/sl2vIB4vmBrg4QJMwWguRLGdXQ9DA+giLK
jY8SSU13ZLeuTnb9caGg9LxSkCo4mjG/LC9f+rxzRBnSMVq3CcEIMPiz4We5atJx
4IaPp6tC+bzWl8KtRvwhYy1QcfrcENOukoZcKKU7N7VDtLyxTtzcNeN2Z3KxTQ8n
vgqCoW9H8whBPv1YtR5nCSu02VdXnoL7YmERbWf2bqTqmvqB/0Bzk53DkHZWOcaD
aiO6/Lum+9NZ+D22Qtoy5YQauzwZuRYGI+htuBpdJGYWZPo0zS79YWzCaqlxAvML
/vGNuYjSabJsPxuuDv7921fJM8LOk/8xhC3oUow9abkex9bXepkMZL1MCPa6YSxp
4Yeh4gAqnHJlQl04b9BW60IL4hxOh+QMKU31L7R+w0+7D6KHZxN9scyMQTxkoepF
lPziD3XWrXhF4Spn7Of9VxF2HN5Ld34hBWiccTWldxswqY2jYuanOE3O4vEl1sFJ
77yFAjJijhIFHBzTh1xf4ZpVV84YEbVo93cRFdSjv9BwhG8oJVH0TfCdrVtgs1ts
jH2N2vXEWyKHJU/l4Mezd3f6mi1Aj5ePfaGGjr4HCO3dLzNS2RZ7xgFy8K4g0seW
5K7S9mihKjYjgu1vzr1OTzKUpb6uQ7oty5rQkWTwSz98UYB1ArP377lQ7MR2WQ7h
Kt33J4X84IAkof4Rn9FUZy0g0dn5W5d/MoHIcjk8c8seESWb9HsICjM5VeRrM4Ou
ewFhPcJJ5N7xu4bS5bxAtDblFbVcdt+fUq/oJ5AwDK7oRC9FBDUWmbY6UWgDvGVh
8y28nYAov8SvhKZN3PWgGCjiVFUxHTrntN3KXnkkKv5u4T44rQ3NIo/uyLShwzbt
tvPIGpM1/9pXzhUbAD3O4wqRPGKnSDYMRDHVdmNGdDdvVHz6oU0EWYo+GFmC759N
GjByROkV+nYWki4pdZYBjj6+XjQtjMTS7ESNm5MHBTG7Ovk+PBKBSdfZ0WaKs0b3
ndoU7nkmysK1QbXBf7usppx5bTWor2h+5FE9v8os/wNllVomyv1wJiZ4uh1zMzoX
m2Ihi6qLu2lO57lIKoS6ijJ5M+2jBl3FDhUbU4mFKErukfXihYN7YmGdoakafr+8
1ftc7u2y7H5kgT9kNcI8od0YqT5otuBsUlhtmECN8QhdaFmY1WHaSXWl9XxP95HS
VnlyPdwkW0YdwrNYSQDZYfvpsJlmymGHB60xnh5PphQg60SFjQebKwPNDnS0ejNn
cS32G3r7buChzuFlG/8Y0iN14Kj5YXXr/evRBFkOmJWVSVlDoKSrjjskhcZ4IY5T
4v+qaugl/p/5R9Rr7ynV2OkDylcNFakLQUJwOmFSF6IrHNnD/T/62SvgtfBEWhx6
Ujprn5w0o71BBCq7u1LsTlOwWIqUwr5CRGBw1oeiYaU3Sn76PHZL+FsO2FuHxiAB
9ScQE8tBQHA1h9/UPt+DxqSsTabumDT82SbyA8gZqXqcUa92XPM8nmMGNVNaXOTy
OxZ6EilMfwT2OSkahoYBsRcJ+DZRwKjXbvr1qk0Y8acxRRAI6GZ0djQsCKTGQAv+
l2xjaIneMzdgqeC0ZXSx6VaoiaURMToekbSKOsBEZD+WgYD7W3SBxirT6G0VPC+E
m8X6DCfTssLqLMvxKFRrkBLZGz6OJfIIK+Oh1Q643RtGZNjTSoD6NL/SJuHK0+Tl
4zU/Oe2dOegCRPnmtnANRIryiqZcbizgTSdGAcMhQuW0cqkSIzqtOjwGoAWjjazC
wEEa3P4ELcL8j0woRw9SIAIOFErDOLF+DpU1mTN4aswaLOrDJVZTDM9oaZem/9DW
t9wcewQrBrqLjvwCsnlrytmtszK9WpvN1yKRBp24FsEF567ezDRCT9md2IUDplph
dKJcumRdoeuqoJ3IUP6sQKM5DTeKaBnheIdIa7IO+DuBZ9iHEb2oiBob7jGNjYWX
tZKIC3q4wbnVAA8us8SHG+jkbSMRwAMXW69uUq6dnJUFytjGBpOxCnVVjWR0jVQE
KkxDIbwgTjFOBkDT1TP+dyPpAUnUIH95nU8YxKg0WY3lSCig+GgXMwyYF5FyRJIZ
86rg4CMSqvFKwg+eJQIYPdC03r1b2+XMG5svd5gfYEcCHvc3j7jHEw39rLDpj3vR
oXspgBlzMwsH/y8dT21kSfeaIsOy0lLTHCy2ShrJxh0aQhS/pB85M0osdfQtSblP
rayCBxZQRarVLGyUMiaxfjqqHKD/rcBF4+kMh+TgvwsOTSTG7Bi0G4n1OtrFQ3iy
0ghBOsx7y/hWeCTqbxcpHMfPPjwC9FwLioUbANcoDkdx3VCREI4lS3JTUbJUewmQ
CUGfBhCQInvCVsORiZNGeMolFojvnuaftAIcOXo3pH55NTReL97OY25Y5bKVnGGN
i8QXLejExv+lqnXqMUjYKHH8wQHN+q9dUsRCqQanU1IddbvBwaEWIsRsL+0vU4e2
uWR21MiLdfblitwCa0cv6ISIG0S5jBA9sq36LKLLdjfGC0goSsVDFluYYR/CUu+I
meG8QnB+gnC+LctEpCs/q0CmkiJTqGd0X1hXmd+GP9g45Cy+NKa9vjSvszD01pYZ
+Gyq6cZwJjEwEGHTkmBnbn+Ap6G2u+Spw6cJJDkvPZtluOqVtWQIx/+jtCNDYRgQ
E85obKIEshxS6uLOY8V+lZ2CNhNeUSAuSVzWwOM+/EDuPdbf6I12XUH3fdCazgek
/LXF2UBXBcIhB//ln75pO3T3rN5lG3+KXzIRKrbJ5ksG3USQ2M9kAONSww8NMJT+
c3yWyBzgajUmGyRK3O/EYcHGcZ0L9hQA5heZzQtBB8uaLVS8DDRbbKCrud6fXY6V
Ut9NETLKdgOIP4zkYmpTtV95lol8UJvr062YYcLdG0Ht1yBqcrSdP8CoADFB2r5x
xYP9WvlbTxjW2ZOm0rUsjSpIoboz34rit1wKpr4ZL2oWmRLZGYyyDG2EbkSXEmfy
zQ6D8T5VuFpvv3kfM4vO2LZsdsThozGf2rH+9PeKffuAKdttlhnFE5LlwdJAFaeN
zrueqWuZV1QD5fGkFODhmk4pVSK9CpQntYXszNIycWg1UMkAHGXQJZmHmT7p4S33
LZD8mZrt3UODPMd6cSk1s01aeaOXIsuQ+vxBshw7DOIr+OdzeGZnGLm7wgzgT1av
1yG2hg8PFp4kbVyHl95P9YPPcTXpXaf+M/mBFpkivRmaGMoFlBHpPzc48v4rEGPh
rBMqTfM2aLzMz7aJKUk/6LyhwYhffd8VMezfCY/u7yeh0xA7PKnhYp+yM0yz2MTi
ucoPz9LjdJi2/K9YgqBCfv+TQyxe4tL2xRpfrNrk6hadRA2sjwTTLy4g5JNfhfv8
++eRtpRUGiOW5peDiNyo9cKQH/cS1fvVdBbRK1+1tDA5lk66IUtFUOMv77jfMCJB
77N7uyxzzJ2gM/dAE24uE1t148LlP+gLcujBE4RCnKAUjYRIX3rfS+4v8GTSA9DI
jjem63Xf81s5PJa8rBunaWX55DLA6T2iaufq9WZnTtJ+yVTr1sWDE1HOJbVZkCzS
oCT/pHw2a6AU9AeOTYd2Kq4q4PqF0OLgwP1Toghr2s18jm6jMYyojYiGWC/uRkQV
F5tb9gX4ivazmCq4M3hoTMzHY9/P+hsZXjOLKtaG5Gpy8zgWUSvHa8bfM0y3OqOV
WcFYEmPCvAzZaTLvooNuEvTUwFjzBMEE3QkXGQ14qMV74xNzJbwZ4QpLjKl0sIHE
FGgKY+JcNv7NcsrvwT9Y7yJG59hoMTJWA8iRdmRum7Pjjm23Js0ZNECfjt470hHM
pktdrxqVbmNAYwIrVLPz7MDL/e4s+qDm/nRo1B3mtvLxuUokJWuHAKCtlvpqROl1
NlszdmnMSY5OVHVFuRX5IqZqvvuvBRSBpJsipOVdglhKvUSPZ2Mwr2dw7cpYuNRV
+AqT8nmQ6MR+t7ArygYOWUERGr9kEd4Li4Bnepwhogv6mQ78xFggDSnqD4DFDYAo
6g34DObPCO7TW7sUtYVffPyPZI8g6RIsMgac5bl3sIZC0/8nzBziBjgT6kZXIT//
/2FMabrDPSPhkENO5rgi2u6TTQyYK0qZibQqyNX/yCDvlJBqwGAQPZ8YGSdhiZkS
rwuLHyTo5OY881c8c78d268/6s+8hTxvqvije3QuYWycX4IYh6rRRSM4bQIjrkCY
ZuHZSf8tBcm21k8EMvuvGJNgLaDsxN2MKsZAtS8I7FVe7WIdNTlsS9pl4yLWszqz
Nn//ReddHCsdVK+S+IS42boerVSaHJUPvP5BDrBGz/v15kufvWoYjiIdcmWdyiLR
m8ommtipTqRoM6U0ZyWztUC5V3B4yBDLnafb9oymduC12pfh/dAgNr2RUKxO/Vy9
tA6jGnqV997nvvPsb59X8zIZwR93iR/J/w2X/rKNpmMGY/aVgKxy/5pTLhN5eozs
PfoAb6qtllXClHG2J1xBCrl3ZQdtDqvxXoCw46z2wY4t6zbJhtxfzHNRcrKOj2Be
O9LQZDoRgSC4mZbb0eXaSkJ7AB6j6rZA9g7OChTCCJfFZdF+4ZPUVP5oBGfO+xls
zyC1jgEsJrCZnCPGbftGr93mxTY5jUF55uomIq9y2ZzYPfw12J7WqKDTfDJLS158
LNIKngQ197Uhtj1sAfau+cDhWgR3yxR5vY36vLco/fI6OzPBaP8aGrrgCyS2A3FA
UBAIWjvTqVTxlIhL/LfRKJnBfs6FYl8xTP5JewauAQ/IQUE3CXrYbC6lfjpTOk8z
QL/qqWYd79xdV17reJT6bMewoW8xhjyk5mnQcZ3J4fI7HoBDI4QAM82jRUiVANFr
gedWLX8Fe9Ms+WF8dCUdWMA795oLL00vL4tS54jti1dqmeL6JVCi6BBOKF8d+39f
C8qEia+m7K5fI9LldeA8/Lfz78HCYtiSX+ACqkmLTuLZpf1s04UOC9ZcqvVk0Urb
lZ8Mn7apw6hsJMeFmDwlM7+URYQnvjodoWOMWq6fORmZq3tKDgOYxE8/dRG1IwDl
PI7O3Tj12NzlYyOQ0xGeefibRzPhwLJCJTnO/Xdk2CzJfKytSFcnvSxt5Kg22ijL
vCQ5h4VBjhyANSCy7GICpc4thBcz835qVodRRNN4r+tSi7LPmz2OaDDTAx/Zi6L5
6si2oBqDm+gPBQ9NhyKMIsf87UOKB0ltO+tqb0cU/D5HmpoGrwQ2xUcsE/Rmc/au
UI2DWOYx2t8aEBCEmDOJz1qjW0LkAvWfrW3dhZZjudRCh+oaUFHhq5DG743T5ric
9yUHL7p3pljOgpOtCaekWiJhlrvSaHHXy35hygRgxfeTOcYbgaHAAqYVrjonchg8
oVTO9QzxGBUDEp/Abu8EOoHFkQP+169ukdNE3P+lP0vjEL9Emr7RhXB7PfB06WXt
KGSS1n07KoGRfd0V3VbIxvJQqOosAbIvEzrJF/Mj+aldmTqNtcZ+lVNwpG9xfo0n
HCeP/3M0SclfyRzQtz1HD24qhq1aI9d6k4JgPHf6qP7ZJ9sFmYY+uk1Q+UN+UA1U
6xC+eCW6bIvdGESUHBEkhqy7yUiiFoUnC9a2j4G2hFrloCZny/xYZpU9pTG73k0y
VlgUrTA7Rip98QVaTtm56OOtlI1PzkD1z8V0rtHLkX4jaPiQ6G0LswimR8/1i6W3
EzDzbbXknymOIx5LL7k1L3Ka34cr+afn1wS48HLGwMPwb77ZQJNaBrtm643ijdWK
okmEwpdsUEEvDxhbFIbGYDaZ3+UHa4+5RWaxABQJ0A4gkrvMxNPTTLEIHO2wZ5qK
Ob635JddmuyAbsyk9BknEd55urvoa+7UDLGutR35MRFLwFjmOaoYjeaHXASma2KA
kFvnNTRXsnYm4tvxmXkcZrIdXg1+chfE2oEqoHL0c1Ga+zh/Xv+V4P4c42DqpL9H
bJ9ddwEJE3cDWkfBWcMNl0qKqJxGXbkx/ZU6iMEXlu58ymw0BrqSeacc0f9iFnn6
CT+NGxH9JLfaMbGd2g/GM1UUqIeL9yn9EV2RL+mSJ1m60XV3GgCkD7mq1n+NcEc2
Oygn4qgskNqSv35KzlVYWVBH1H07H//77H7ZyLMV9+P2+HjdEZyWPQpkOPHBS4bA
L358UnauUcxrMnpRvFxaXhfN2rJAfSwbZe1Mal5+z9a/tFN55eQBV2WzI8NJHkVZ
MuTXJtx9DOeW2ezh5J3nAbIKHRtTDQKEMtnlSjYMVkeVCWPriYX3CJQpPN3Z20ud
zommHeT2KSF8vlHHGXicyfKGFFGuF0AKNw1tmz1E8Ai2xnem9NUnhuMbtD2TY5m3
xSn1ll9JZzakogjQRqQ7YbYoopX8V9qgNujYCzEVDvgTGT92suiPwGkttlsBQCKn
7BOr6o7bI2XMN/eqpCroSW3/dccjchsiOkv2zaBForlRCQ6UfPGRMJntczyq8xHu
/En3TfOD6u7VwhjdSxKNSV9IqEpVfS0CbQKXzOjEmR6H83ia6FX2uV49p0Dsa2pE
qJMbQBjUg82WvEGOge8fgnRghOrNBaV1Rmq4TXHmbqJpj2lUPq1RWUyPOh2vXlvJ
Ls4Hdgsve5IPYIFNBhvFbjws5afADLyU3UUPPN+Pi7fDqjnrITZJMVQ78YfOSR+G
SifTMAejK5c7NmNMery2fY8RqjXNOBNLE81379ddHcdUCPm518WxrbF/HkPHFsA2
lp3o4OLPRwD8EC5PvoGbCqPgA4QQRRu+eeERz5m8qS+hgnG7X4uVe2qcVIcZ2LS2
4rq8y4rvgavtceyqooUQk1pOMWbj8KbaUB1yvzZzuVvwupMwmgFJJsaBjZDyrHAM
WdGx42gyvEhENjwjC0ekmB0WtWkGDrrnhIZbZzVKX+Noji8dFH5/KM7ypT4+87Xb
7yX7pKDBYz59Yq+XG3ffdrYM2FmrAV4hnvts3I2wlc3l2m8AAQjEVX5iIiNkBNCJ
QO7dWJRlnBPt/calnmiNUToMDIuliE8xNRL3ZhdY3W2Gjo5A9k+2k1R3pkGT3/lZ
BCfJi+LDYtKGW9TetqWfDOrzx2cVP/Kfz5/80O4Cv0ah2oqe/N5N2rpzEDzpUU7u
AraBS9HlNA2DC4uTNt2wV4pxxXNeHh53hjqLbPnt+XIKQ/p683cYXKIixnXBbebd
Hxxpw4dXCXn1c7Giba3Le6cg3x3tPBf5pVMO+CjSTmGYZloBvP5OK5aZqI5upK2h
8qrQqg6vpCqiEHaR7WdPTIY4V3CAgh0xG5DmxtcF7dAApMkV41cL85oRl4c4o/TT
Xeh4RfIGRDlsRZ/VVx6OmTRz+a2aXe4i8tOrcF/qHmqhMfYP+TAV/jmH4TbuU7cx
dYwsIARiCjFdrxJ6IXWZ/iX5zMv4dbgeVuK6+4wXH/uIlETt2auHkMt5rpkIWYIH
CK6ps9bgNL8nY+dfIGScsaWgFjfThHKdGeLbv81NLudUbMroRbyIaA+KgZACz/LR
LDEC/xxKplwADNGSbUj/sT1UrRc9WqXKz8CZL46N0ZaUVKnb7n8QXYYo5schB+9g
uLfTWQZFWfMbNyR4hyIoBLIAGXFk8dmO00pX29a+avwxOEzrhIxfO0wbO6aU5EBm
CQsIGTvfJb8bFApFh1RAYWhD6gl5ITq3kROJgXz0ap4gBMtubz4c9P2BKEF96VSH
i4bSkS2FYpZMBDIiq22Bhe7xdlUjo0QFw0gnQhhUzZuCXD+OYbA2IaUi6tBPLdIf
QfYSqMER5j0qy6MUyNEL6k4pYU+9C87WR/m+iXoIc9TeBvCbZ8/pQrD7DKcEhe1N
DVSqIKc6FIVUd/zi6tfAkTYMr5m2UvNSJXxPvD5+eTKtA6fvwDeXtmOpiT0+TbPR
Ntm1kFirP9qnYL5LDMvlUoSV/ExxY/Evnf++zbTSUIb/O4MnldoGl/jguCsjvAQQ
4mptKHpi/5OKS7HjHZDCYA7dKl3A0jTGz/yWkh9mKmmcz6THHqsZTBOA9CqmlcUt
18UWlmpS2gaCJJG153jDJVzQUD0Db3NdRbgkxZlzeHPB8+5V1rhAw5GhoYB6hOtQ
+H7+TkIFLCse41m91MS331O7xo7EX5SawHMT/YIrem41O5gPZtBSJRa2jJxnotcz
V+raE4RmdBzAXNDetYqhhOmScuBjfOFOKv05v1hkQ0fTwIn7PXvzdgN720EJV7PW
Vj5uC7PWIU2LxmiXzYYcfGHxCUalWZDLtoZjJ5ptX0GnqtaEKUQ2BJnLR6UWe3Kf
7awccswaK1M8I/s0e7DE2YUrO3y4jIdZyjqXX4zyQOjIowgPNYeg9aXGkI/JmfOU
cdp42udpjKZYulyQ+hrQeN8IzIYXgpt7Z88zTs32tZdeXQwl3q5KfCMQIS2HB6aN
YnVpujTOKhK3mGccEaxIqPhU1+KWg+TwSDIx4iTNPbmaEdilEGY9s75DvjP1V4Eq
y9r+7sd4iSou7PqOuUtSR5revAewN8kfi+yJ7H8L5VIL5sN7wYXZqsbWi7vDBTXg
h2aea9yHtkmc5+wPl41c34cqPZLECLxQGK2DiJaRbxxRAkc2+I+gg+JPSosUISU5
gqBX5n9QBeDmrQkTiaXS+QmsfY2VmHL4TYQ/k0KZVk42V+83b8fnqUVypdfMwH60
f4Qk1uaobggM64QPRUAx81UMx4zZIuuGD6UCsyn1cSwUYnpNf+UlI1OIXdAePzB0
gRH9/dzfARuokQ0vzrJw2iSuTjhI61xT/Oc0EHLSEHrb67Nct/8/VWNs7cIxse2u
uN8b8udn+4WCZAqb2RXrp6ADHGa09moCwQ0P7IJe5GfTN3qZu8hBjbevVOx3+d7D
IEnBVGhoeyaTwrXZAp82qENXTnnh8jTXxlOpgPf/yG9f3U38xLelfX4LNwj4b57p
pobf7Khu5V0fPJgBE4gaOVhupGmj6C+UUFg0aHt5E0Z3g+/cXEVAQupdUr3KE2ze
9ODh81ybtcWOP8y2Q/fi0pb70Gm7RzP5mVJL8h1P1sU/cbQoOSS3Q0Z6zXLYeDqD
azNRk/uLl2+cqEsC67vzcTdQXss1Zs1WP/aPJXuZdH/D66KYdVQAbQUuby7ZhF2q
gP/sJFms1PmOxzFtCyIVv9TrdhDTK9vr6XfCzyeoekqF90Z8+bmseTL3qdOXjj20
WpO6Twg85TTtg3T6jlV6fiEWLl2UrIzdG9UV0qTHKZT1reVjgM7ZiRi1b2sZ87Wl
TBY13Gzu4A+l0heRpor9CB7KI4b8ojcQQ5aIqheFlgUfaoRkCYeVGdjBsfTxYu4L
sWh1KqmNH0Ev3ZoZeVVtBUKoEHzJu1ubbvAdWx8BA3OkiDaHzdQGl9Y2zOUuScfL
8TSgYmZ/57NhvhcDagFmV8qL9KFaUnCV8u4yofaOnUBgwNXlVIU6Kcrc0iko/Snu
GZwl8Vb0ThXckGNkTEdKXNKikqIUALSxu8AUkSaMvXRWK1vu6v5z/piGnL/YWozC
kyqdVNjvZV88t5DEBICMRtiGoV/s0QgPYkAj3QmmHRjdjV0FaO3JJlu9U/0E0mWW
yOJcoXSbP7eDaedej7txf5lkyabxpSyMwak/HkCe8tYIS+vGKSILKmarvkC+rkKf
36yGBCQ6DvbhP9Xryiu/yt8VW3dFQTCwYjOVXeTly2nU3gdQiTliJUfem1kI+tQU
Vqfk0aN0pMWkh5iMV1lpsJoNkxxl9G7Iz2cTwjf1DJOI9aml/3CzOH3NfcwKBQOz
EPTc21RNvczKN8DRtSRN8cXvCy27Yb00G7yJWxdkPIMNsODeqeQe3UWWZAHrEjwY
/bz6AuNmFxrshWzz7esTMtLdcQvCx0z9SGcxSleEToMHhRf0/Jm1lGGBzw4+JgYM
aZTqpJTG3Yfw7cj5Hk/iRBdDQ3Wf05XxLlPnNvhLiDm44+N5/iQIZ+9P70V1CIGI
3W+YJOsm0FBFr41hVydBMsSDrdRN0eCJb4t7ZQ9DDmrjjbdGnaoM+CXjDHuyMCjo
4S0Z7adLS9hbQBKBYU39AzEh6rLwxo0qgaxS5RAGdW1Mx50zQT4J6rNnjPMxciJn
H3Kc4MnLr389pFE/GMpa0dlAajc0RaB8dal3LOZaCfoTwiW/yI1HUrOFP91Gwp+r
ozOmWlqDyNJjfICKY9vLsbwIDx9Eu+yNRKfvnNOxXuub9l0TkInc84zO4JJ+l0Gj
5Od7u9rARQyOp5IpXJj0GXxqNIlWxVjcQzmps/7+eQPAMseapL6GHof4t87+maOh
BPQCmwdTVDTnRq/6VwoWrY7L/tMfBHyx+eMKuru4uRfiCXW85NjM0Gk+hULSpsO1
YYhfbP97mFc/Uc1HQvRxeO1Fl0xlV6Sznx2hvoQ3lz0bX1LtkMqu72yoIvrm53yN
/N/W9J37jJ431PRIuYicQ9U0/uFv5td/FJDGJtpEt7gpeWh8PZ/M1E8FgG6ZCzov
5xcKzgK07sTRBfB4e+l4Uxn4lGn6u9/KbP1LJB4tTBpV6UJ8DRdd3/7ATj1MvM+2
oAKlwgFEhMLAgMoPdYC2kdvMdjEWRIWLnmJE8i367vzBgfK/jTh3IBwvuab2Om3k
6vDC4DveJSu4JO7U+rIOJ7FDavZCL49yL1NOl+q7ZfYVmjk53ycJq30iNmVXCuDM
mkQEVbkOHZ+iXIBVgKbp25/FoYU4+o1QJA40H3y327D56rAQb2RXRoMHuDIT+rFD
fXMP68CKK4XOgOn8Gin3uXI1GGa3J58ZCFNNgHYSW9CRFo8MqIy65+2ueJhR6vTF
eGWn2eOfZAlRz9Fw6Da582qkCK8SWKyQ2XkClXcfkaIgLSIWaJA6tIM1yBJmncCo
feG8nKhl3bSq6ChqinfKwriPxFnFTvwpvG0v7hdiYgtKz0nIU982wVgtEJzW9QV+
ChuRsuMOfDHTHy7N2NpzyQYty32yJLjD01pUAYYCQSiY1xbicWVA3mvRuyYcWT+G
tisdeWXScQia0GSGlkJPxeL5Q3fsrJmmiTNXUqp96xf6zDFO1ns3GrGMKqD9lPs2
9HuWsL6EJOwlIUehbu5ctpM/Th8ZW7zn9DiS/TscFUP49v6M9GPEqq8kp7RKBrJA
mKQOxfkWbDCR5UqL4uWQWpCUDvbIBVn0oNgsG0unCz4p/qmMpN7pLZQoLVeLenEq
bn6mIlxfsrwSKCdrNcqxUlHLBJfhOZ7SF946RtS6+OJ+fITivL6DFCoHB/NVnkN/
MR1WVQnZpawNeejmlIEVZU16ZwDvCWhWsVSv0AXtjngcT81MwK/zIdAuibwc61vR
Z96OSf65+lVgW2AquwHEW0nlUOFogfMPAi/gwXABEeOlYptLyPx426tkkw8q4wP8
YKUUPIkkSzM6BZRbfbPipWCX/ykZfivC0TTqI67ub3WmM6yRTI8HLw+iAu0C06mg
hlZEUF5p2OTqjH1dSDeWgi33Wm22fxqYvXeW3omicYeVHZpxqU54e+upTNMc8xoj
omkRUJgcKiowcbQoSzm41LG5cumsk0xkKspTTFoifcf47k10Ngb6Odor4tEfvGWB
yXJQ70sY+KAXPk12RG0g/HQ0gMVWYiBM8Jn6DmU9LIlTGyiJ3cSFRkHS9XPwNaKx
xKyi6gSuZE2NR3G8Cj86un4Nb+lhqk9qRzmwsUE7BVz9j9iw2xKWYdEIleTNmKHr
dwpb7tYjrTQnsWPp9pHQkwnOHFtPhCDju5br+H//nU9Z/09bV5/2yEdC3HK1d/NE
Q+Y/1hH6ty6jTYodbbGv5akQ0H/hi2CWgeirroLmWDrDXDA8gciT+EpAFxnD4bfx
afCk3Bp5eECF9XKB03+UZ3yXEwE9Ts8e9L9+4mkJQAtds8JTgf5jlHZyDANc4PS+
jOcOOCX4YYIGMJ6ydo1yqagjFC+NuUGar71EoKi2rMbZYCG2pcDv/zsSFkKCSKNI
i/j7cAB+qL7zsZ+k2RBO+hcKADznTOAaRaTUZP83YRGlStHztJrhsCYYM2c/UzKu
3/CBxHX8089zczhaPPX03p3CZbzPxJpF3QLdYV8G7rVbPW2U1JY2BSxy1AT8bnrt
UPGIBtfe84ct6PevLGguT5a0o+T9iYrn8QMo8319McXK5FgSXqJYKfUq/UHW9mVP
qoXdyIuOO25nU/raFhNfVyDpLAn94P53uu+QW382I+mOh3CLRL127fDpLIcG3UVC
5prAtkIATDSnQDjBQTkrj8CSX4EzfJsOQ4cfnxu9odYf7Y9PKGsPc5bYoixC5can
H7AbS0G7hH+lgYc0CAJLfCn/PdjYGgKXrCBjUyTNXPUcz2OhuHQMLOpk/H9rJ4Bk
fB0hqGpAJLBr97/7So+VtWeuTdgGoJtIAEb1DG3sLy+tngBcaBeDYBDem2RSD97i
yft7yisDN9dn6XLg/nA+xiNs/Bj1FJioOV8ake89S5Bb1WzTwMh2w6G99xyso3hn
yCpErYe73u8Oraf5+yZsdkzf6SLbCWVQxZnchimjC+UC7w9i6SJ+VLXMmWrK8fMP
dl6W66bU8JBd9idkvg/rj2lCCR9+yK3PcL0Sr+ZJ/Gx24nld+q0lqxR1EW8an/ev
aKmhLc1p8oBlu5J2gZYZlDulVjC5gl1cgQ9nalgJUd0FYiJtzNJ4L4ibcw5Upy91
h8Qtx67k8RzVDXzpZENpOYBsoBJ84v1uVuc9G/PuXflTlQoHufRUSJqKoYFKxc5b
HNcMbeMuti5gKr83ogRiMh+DZaGShixPuSiC88lLCySmkNe0MtbyWGYkwtCHlYlX
BSGacuan7+Xtkw9yBvmGr3kiTQdNslEwPoZvEQUj3sXDzLxoL8zdEt5dKZ4x0Nl3
OrOpwgOgQVc8J/3qfqtWWUM1wpCK0sQa0j7WpFCY8DMvruDQbKZtrXXYW1s/3bys
PH47G+/Mq9UP5PC8zgta9euXHvdPRn7SOorbxSnAypXTHTcM7EcHw4eekJdIqJqc
nj+YohOKD8CkTz3aj31iVuRBRv0yY8rvMSMklqC5ciR/0uVieF1GC8FHUnN5QwCC
fHuGeAiKiMkPsubLC3Z/oSiWK7HNuaa9Rt59uLw/OpXo2yMvJ134U5VB5zt5fNyX
lJLTzrYZoniEn9WoV/0bzg4MNiUvXJnVCZ9X1dwP9cnHK+pBmmxhwKfhEGzEcxLW
RHCh7G8e99h3M4w16ZVMfuL08gQxmzW55HPPDGFzcgZVrekniGK4Md0ygMomP4u4
DzAvUKYw29+TYWcXtXKZN3DluctzkOkYV8FgKBKN/as5bjLuQOMU4dpFHr8J5dFG
JcB2gcsctkA9z6q5Izgyygk6KqDZG1HNShyVOH3wa0AyMUfcPr/h3IDZHCDjwTe8
+CIHMpRJFJViOfaNbGhWjKegbQL+tWwZiXohjIsJkapDBCaItEb4U3HD6L7zafSr
NGV+6kHHn34EXJEywTV5cHsgB+Y9KW/T4a7qkl2H9Qu98KRzFBmXWtJfXJCoqMyA
s0UrJBx7H5DjHPIOwbXG+iTU/30MnXWSH+Ja8B/vyPcpJkq/++qOrKPK7VAbXfpA
jovyu0aovIJsvudlGf+Le1Fc4KtEQ0ArSisDrDqyVUo4eu4N/D0ip4cYXiaV1WGL
wuqokssS2sIEQ0y6RMzVSyzm84rJ/+z5pNnzeQcsAUqqz8X2hy0qIXDnylP0CU+Z
0a2CB0fG7KWp664tqNxY3APznfddS2socc0OGlIjD60Cxl4JLkU4jYAbnRJCK4ko
BnP0wJJ+bIMFdppydeNUUkEMsUXLw2yzLOnhifRiC5s=
//pragma protect end_data_block
//pragma protect digest_block
JpydpozlwUOJhWX/YHYCzwzkXWY=
//pragma protect end_digest_block
//pragma protect end_protected
