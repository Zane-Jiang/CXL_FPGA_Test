`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
SCwkcIQ8csnP+TTR7Sd+ugQe1oXFOY6bVvqAfME1hy5Fpn9vlmbUdCUwYhAX9R8Y
NN0q6QQUIUFroeTTmBWlOUe/2b+6I16ZMEHs2XbRniIY0Mr/IqZlCadP2vobpTUw
YNea+BYpSqyXWmeeoQc4oNXGc8q2O3QLlNM+t32lemQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
z5j2N60XW4p0misE/UhC1y1VajHsrQ3K4YHYgmqhDA6athiVpjIZD2ruD2NOpvke
Bswu4/y6U6j8w+YgxA1/MAzlRkHu79kvEAUksaab5gRyFVbGI3Q453wu8Bn794YL
M/QVJgh0bDZKeB0GWGZ1kqW30IatPr5pYxw+BKxqWJtBTbIgLKQIrG4DPb9SqwyH
mwwdfIsKFj9bdxTfEG41GZADELlyk/MgespcN2Jc+Sz+VU016KK01h96PZ4HOEwx
nw9+it6+4YFTwNb0YpZnr6B3fIHlMW0VMfN/TBPgROaY1uRe8G43NuoK2DBtny0j
gNahoKADpqRkyyWjqRq1pcL+zwUSqdtHBroreU6/PNlyxL0/wnuNnMn/txoceP5q
LNM83lZXs83CSGvQV4jK4FaOiUQRKEHI3FGUeBXW+AUzEB2aeJasEe1ks2aerncB
2hIIceukBV/0ROg3iCn5Vjo+BAeq2l/B+b22JX/yseHg0kkGRZd8q+QM/KObIged
2RP8HQlDF0LBWJ2JlniHTXlmitydIaDJGOP88sBSM2qpzQPidroHg0kAlbAe5e3T
KLjpg3+fMm9Rz81aDJ7J2e3RjI440i/CcBcHqJc/e54YGRdbNpLis7Z6SOw7j4sI
d9EvF1rc4G7lvuiuQMOrkVEBZdsqN+ujfhO4Gi/RB3dHQ5QCa227/pdK3VYoiYP5
yKMfzAyWNpKobz/ct3518jSoNk/omHS+xBW5KsULestgJoRAxHlBg7RrOgayHr3z
9GZCq9v/J619bs+eFQeDyQg+i0grjYvVxxKeTTZUjiSbQLPGb+LBcf8bYUmfI4r8
KrCWQFHBU8qqDERVip5mGXvsQ9w5Zc4TWNZeK6k1oJpRXt9d5UXw28Pqud16I0er
4U99FxWV3od9ysiGZNaOnVvHBwpymCsVmbUcyiaBsYlESikzeyD4ZLyp9RvFbd6G
UvJ1wsG+jHG7zYObHsl4TPDL0qNMESDxYX97+1uz/M75OI2Ic0E0IMcla4zHjXRL
gMaAzUK+xzhiylTWu2Y0Vh9Ff5mNJklC1lX7WYi/ovt1HdDtuRz3wF1bXNUgrz4o
BFYey9M4nRoZTzDEcQc1XROG0415/c3jdhlfONq/bPeyjV00XjCAykqSrX7j0jbd
eeg92Hl5Nb19hoFTsjUPT7mt97GCu4v+t2DnRgbh5m1fsQLtWe0y5onOfzES7MN9
iYNQTsWYZW0j4KMZhvjXRIiWabpw9Cy9zkg4WAQ3q6XcraJ08sClk3bnO1+PfWsV
oAGuGZBIZ7dPRwFWVdjjerJQm0KEAAh1+sDuuKdtj/uOufJAkmPTDCghDYCpKM8h
ezYn3lvS6OwL8L83/g8cbje0dQ4e629PISMsZq+bH2TG8sHqTpvKOn8SkYF8A+ec
nUjFvUNalIsjWPjTFMU54RWn+bof06UeSJQNS1iZvQ24ghe9ZodZaZHe9u6geC5m
FN+WMtQKxTphmx7B6GPawNyLVkUufPqPuz0KVl0X4azw0Zeyc2WrnqOHNfvKNaPX
MrhR2wCB1U69QCF3DSB8C5LTceftPS+dbtCxNk0QWG4u3YOiSvzEhegEg+JL34us
tL8YbtXddAlEsVaNww1v9ZFYf/U2rnoxt/o0/qumhzh9LfD3c5kvE9BYSJCIttFI
XSDu8QwUhOm7zLdJi08xG9ok46u5wjfgabmrAAhwleks5MWD0IOtiHWOZmkpHSHg
oblRAqR0wV12gIpspOlZ1yt5Uy48Axz5MfgDgvW3tFSxEXseYSaa+1fGkzfLMui5
i+OrPaMq10YyZxiubGGQUgvjvFIA+M5QUHD7ysEc3b394KNtE+3QKA/qW17gtSOw
H7XkxrrkZ4ga0ZGzV0Xlua8XRPT+DoNhwh9nfmEz2nC6njKQQtfn/QntEZGw944/
L/ikfITRvaw5B5R1berd3vA2MJ0VLZgXVRCxXQyvEEbwMp5cIze2+ePIKJcGbQ8A
7S5MejRbZPQvJGWuOLENiTgPMjNWAsi6jhPNRbjHCiqqJUBAz/q2JdDuWaGF9bBc
ltHYviUvNmxqJzz670y7jCgEWTeVBS2+RXAa4tQxPFAVntaGGmfeQwVfTXVxrto8
u0IlLmJVYXIl8mvio9yfXu3r7ZLio0FcTOzMl/HgHyUB4VmHRUU1scIpAu6gKo2+
MkB6ReefUIn5jY5yu2G4AKdARvoTonfkRNIZx4NRVYF0E4PfFw4AxsAgSi+ygHL6
6+ezwfQB8OPezwPQU7EGX+78pyViv6u4JAixBzSxsuCld4XseDbXAy0ysP/kWJ3W
449Mhzc/vDEAQat+dcOM7bKWtfeQUiS+jvWh83+iNpLeRj17vS4CHoBTnnPWVbCK
K1am6JOO8N4RgfsLcIEQQZ0hsyWMJfCo1v6GAXYh5webCtxL3aHJTR2qg5UGhuBb
u9pfXOmg8c9fxlKSwwljoOlZuGJEdRQkRgq7zuqU0nmiAVB4oKozfjki09qVKHtV
O0dAyMC5RG4Y8R0m1QzB2xb0ECw8cboOD5gosdQWYdzSZ7YA2+DDqwf63jqAvRFw
xbulqHQaige1MSloeNnEMb60KVrGvwBtLCCu177WERlQ13+LVVujemQHnnIMoSrg
qHoZ/yyjcEdpT7Wm4GcMAPwx3MPFjSHPKxx7N/t+ij+04Egq2i8hXwu9puIAyZPG
Vv83cJFZUmJu8GU9Ekbd7bbHP5FusDtzSPxKddSsDfIVo1Fy02nATvN0k7XX9aeo
WFMWlAx4zapI5XYN8N75NoETEcbvb73J/kLmDWCbQL39Hn8YuK8SI/K9YaAjRx9t
thZyTzD1zhoVL0l6oeAE3Kcloy0yQFqqt+XPm0IuZ7fUm2Fp97KNE9ex5ONCH91r
BuKqjKDtNHnYILi9pUS6AT7pFqxnMRVCX8GNUAINOuNu2v7uzheMAy9O1Qx4xi3O
O7JF9bcu6HgyhrcJuEaWqtoojXd/Vw7MPTM7Lyqhjv1ABMMee1W8Newxs78pl1jq
PdiiJjz0fgpadsELHJy101vr7gGUFu0Hvl/M7g7PcGZuINjC1Ty/EhvCfhkJirO9
laaLz3mHtlAUJQV7U2ZAiEdNSJp7rxJ3F5+knLsP0mJKAgl1daLneIGXIHKtYhLJ
ngA7ltYMcyd7T2Xbr4PzTvyQBBaXeW899IRqWS2wrn+7h0rYxRGSygEC5vIHTWp4
3L+6G/FboWJ4rJrqgU1PDQs9bbd9eWedVg7GNOORMYYQNKorb1HnPaghS3Gt65KI
pejlV2ISYInC/Qqa7WZDxAaX2oAtJhRNBBqI2t1tOSG0hwYjKBDiUjcENTic7ZKV
AbClVI5H05pcz843PqJjAeFpZrBfkeeOJP/aCG/aSrAeYaoeKGsk2m76Nfg7udBn
4RvZpSG9wfLtY7MdozfZ5DgRXWWObl04/B7j3jY3f3jvsZ84rnXaGjqAz9cRQDaY
MtQ+zR8oRea8k+owCQlQFwW4CLAZ7G5Rufopb9pAXSZ3o+MeDFpND6Es1n4ycayL
JfzXEJj3glG1F3vCHr5qiOaXplcnn6TggAgH2ZeY62Yvnkg+eg/DzqF3mgEQYHOQ
tyoy6WA6sBbmBGujSFLhT/8Wj+MQ+QlJF6JZB278M41mAHRT2atSI33/6GT0sI8U
BPV6Ms9IpoyiUo2858YsZzEN+GK0+mA7+JrBgb3/TKiUQxaeSxyv7SKAbGzjS/ZL
PxWlx+cCnBPdAktPEtNY7ZwPxD4IgBhkk488/rWxhw2bXciGmLiI9jLC+J1c4cvo
0uQuXdnZl1fI0CfUrIRIN5jcBLPAAZ+EBsIxtzdozlsSRtu8r1mFkGTYVbrvrfS6
jBnfcm3nJB3Q9MaztAWziydqF53atGN1yOMvqCAMsASL++Ams1HdSp68adBG2KwP
T7XBDpwG/fAQBCtR9XFUhHlE4tUoQg7FMv/U8EzbmRjQEFxZAxbdNLaihLSz5TOS
Jt6gwM0orla2fcM8CNOfwItLNcXPUA7NJ27wE9LFLq5O6dQVvtEfcD7o/dexrhxr
DbeyeM1GHE8+IziJz7GNEcm7F2KTjTOs/Iq4yLtfUjoU8ol5ZKFOLXcfbdjKaioY
RudpY2srj27oBZEbWNAf3xV01wb/1FwLpLN90rpYBxMAtCFGxHP+BtYoPZ7b0itn
9j1vlzWXZX3UD95i+w3WaJ4qSc1UdXY8aa8tVfeLz1Ha2Sy1NhHU4xIH7HJ5dOj0
BJZhpzo0rKSuuxo80ubwSpS0lR8EXZ1MW/7tZupUgr0uQq7iwjwsb+Bq1bSY2mYO
0f5HuVsfsOAVJtowXxr3i+VXYwn/OtVOxs0l8YZ1E4MSNX0gCyKOkHTB9ACaJ9iH
qHtX1Ngo+lR/nBnHKDP8Iu5+1Pqj72VrsSCIfNXdE8/9W0QRy0q4y9TgYxQG6Juz
ldSEIcvW7gbDPFNciauxXhTEO3144nRrsqpb82KAD2RHK/fAAckaaIQ8XOY9azwN
Y4+ux44xVfIITURkuCdy77UXhju+wZvTuR6+l7jtKUyFmD7Mgtdw3h24b9e9LbyM
n5mM7Z//EXngMUo+9PZ5UfioIwehprD57JN8rFUNVQcSDmSHQ44jUBBn74qsiYx3
qWmlxiCG3CNcrdax+lJqV3EZ0Ic7wCQJYE0tNchyl1IFfzHOSiXzsYZgYSkb7Syp
gX5b31nt5BwcdEjoceo06XVq0IL8dPzougk4k1z/etPR4Doy6A1Cjb0QL0jL3WWG
0qvZRw7uG9y6F/x5l7nPupRbgQLIKTR/DqbL7r2eP2b1ZFriXhK2V14+xknaLiaY
xmEg2ywTXzChDXnGv56VLq3p0WdlGEKQBy/RHkugOCSN5u5PPxPGjVdxWzS4tFYB
vh4cANOe9JpNHSReqSeywa87u6O21krqBMpczm0rB6CM/2wxfzyA6CexFTaSCEGX
HXgS5xG4pMUM39YtEprunKDttxWSYjXPB3KeoddBZYHAOgYVCVD7zqQdjIQUu/JE
oYvJQu3V9iYmXWILxodutcuZ9vJBNxqC61pF+Mv6OL58g7b89/mkXgGGoCnmjxdA
SuWb+vkYruZCoVjC7ym5kXgsAw6tDScj0hdNRZ3Sofjwbubjn4bUoffPpmM/rNK8
RV8jt5lrzMiX696GV8oueeFgL2iVosHhg3vQWdlZj7B58f67ffZ/RoIHmcSnOSJ3
RxHMjQ021qavhaYTqLIu5g57lXnASlJn/kgjoaSf1/S1jBdAM/TKn0g+TZ59SKU2
3m8MDLTGDlQ+b5rQlnyLMTsYEvfLS9GfhqlWQjr8pFAOfLKPJUSRWUxDNX+ZKDf+
oEvPIAJzKJxc2y5WG7HJiZ18J0ceQxPTCEOrnirKyoVLkZkXUT/lyh1gF4pR3qNx
MuAdBZX7d6U81Bgl024H2vSpGOyWosNV4fVnsP+Y7X2uAE0iF0wYzw3g8KAQQ03h
b9IGZPV46aicn55OoIdKHNrtzT4jtz57iswRCqD1rsMJd59SNkdB59xKWOsyduil
6vjjbQyPl/uZY9xwyuw2wtBhJWjKyPW0ur3KMrIhbFM3m6Bxyf37H4aJ3ldTZA+x
+7I2OQauJwxENNslItZCwQ5M39wyRqE/NOXVRHTachu5VI7BwRkwZniYm7Z59pG3
wWgO7k+4k1oCsipjqiPFUr0q+Pr9Hgi0w2Q2n1UTIwnDIVCU1i7Nbj7OcAAPSJf1
Aots/ah/X2wpg7haHrhgKReUqIr71Gis5Uakn3tvKNvclEDr6UzkX33Byc4cC3og
HU4MP/g3dT/nsvYN+zbHTwhhPCkX/9g1zZVS+lf7aqQNr0/As6SSFEwKZAcB/hFF
6S/FIVPPsyNE98H2zlIk592iRVfn5FJycQ3Wy+BBKV+u7infiEmkA/ygFCSrIN0c
Tkb9i+LqReLDVaVto5S/lO8AZCqGj/MpWvDZdZNv7O7ulDJdYUNXTWPxdt7aCpn/
FHLKNmEwP8osKOKSpdD44i0CxhM4+Pa0UvyiTdZcW37MBGYrYaUEr8Tk+Y++mGRW
TK6o4I9NcQ489I+3RWXoF6dbtxzjuI6jz3dFgBiBaD9HK1mJdynPpJtQjxnTK8I0
2GlAwRaiMnYlKlU1ZRnRq3FJfX+GBHTp4KZiFUukp40aJgzzcgdITLsulAJVWhAE
5mTkKVx8lbxn8q5ECiLswOV7EQiI3CU5/4Xbg9d3cXvxWjC8JNAUal+JL62tGi6v
wcNDi/R1NaqF8z7i5WjGseroefue9Eq7uDjvAz13R2oBJYXWKctpCdqigIeUJAta
uzaWvUP6aghOaMG5PAmCSSsSqCe9iFAbG+RFFgrB4Xo9kEzqpo5XfbgcDVG5U/jM
QFc4Y6q3pj1UAnHApgdgYP79+AkRuWaCUq6oJwFxXmgzzjK2eK9QWx2Em0LvNLTT
b+C6q5QFlOrD1rMR0F2R2AUd10xs5p+CPxD0S8rk3KuA1oMaiXe9vA3AWZ5JUkYf
f3bx9EzG+wcycUEAFwPmY/drkyhI/Oph5RFYyJ47ftRvsqe2LfQ2Q2qIgPdMGMGE
jfDdRgXHDdLUEEhFJ9ABx8FTAk+Wm7Ncz+0bDDaj3ktWnjhEx9GcpLiDP2XZRFjb
pIg2u0RVM5/krCDcuKZ//eFzoiVkZ8edGXs/TA/5vYSMOk+KyDROsMYh/YZk6+of
ZYouSpnNfm1mN/enWwGW3kxOw+0YJBMcV5NCKnPEdphFHgO2taDRjKNS67H6lpna
LkUpGCRxnnu+3NSzL4kI6J1G8jpTKMZgcSnOslUipvqq7r51CK8zjj1bjA66Rgao
pniULb6ISJss37WPteO0qBz2G0uWSsxKhEF7WtKCRXb04uE6Fr4Qh8apDrDL+bKR
YlKVGd9WfkEfg3O8jPh2ORxY6eS7zSx9+e6zJ/1uxne1nOI73DX7ckRadJAp/KVH
RDvsxLCcAXY0y0WS9AEBE+4eP2Z8ciBQNV8TXsYOakf/byjx7qaZnpkBURaP2My1
VYMnQZh5qKItoEN9iw2D17iaNlIHR+nIoSHvsBuVwiUM5YAVkbuCMvuoPFezTWyK
zxCj+JYyMeNE38m5ferXi/7y6sZgr63xHBe0M4jQdkEkD3Tl4iw6Qhi94mJqFBZV
rXRKhn8IZkQ2r23L7P+8tPkUlsk7TzM2Lct1S9tdi7O8rctUPMLdcwMl84xsSXU1
V2FpspoHs0fzDnGRKm4EoZAWg5H0S2cPd4N31J5iM8HAO4X+r3+aDj30qz4XEhpA
TbUC7dUth9s1ynQO1jaQwP6vI89bakJ62M4jOsE3565bwxZSa4WwLy7RXI1KRkFi
VpT5rOBenvPAr6s5nSMu9f7jsR5kq4wPxkFQn8wzDrlv7u5otSz+LVdfkB2Kchli
CBbdMRl5JnAxq7YXoIv/zCnG97LmjFhONC2/aEjBQTTTmubBXQCUElpbjw5GOUwT
Mhysk2oja/oojhOTWGCSC10mZvoKIxsSA1jUN1yIxc2ym+uqfnUDr5njMv0IGdjN
xNi1RDjYWrFzoaYbTroP7egLBHPjHzK65GOho4kBGCEHASaTA5ZBajNl4EgMUwel
CG/HS6FT+Rl7vE0dVU0Nxgmfgpgwd+gx13ZAkoC6dDOap3WlawNtk8ymJbDVQ7ET
Nt4tU8U8tfsURROCFpT8AwhgzwSi6EFf4q+XkyKCp7RRB2YAUz4VO44YXacV05HJ
l42y09LqdMLUafB2bbIbfzpq89HGdlAcKbYdcY6Ro1v78bIHWhfuVOhAiyY/RzrI
t8e+Pq6pWMt4XYdj4gnHteOscK0SZOlgQ4QRMC9mTa1GOfDZPv75i21CfaT8K09D
btwKEUd6UphsOc1Kp7al39ni7B5i96FtjShNuGSN3NEqyEcA33vBPubGreqY1j8u
LK1V3N7Tr59RRfqu7NxwSp9f6IOG5UehbJOuZVb+5RGZcLWN81s9elFljIuW+1Io
wrs79MLseoEQ69hDohKaAkhfza6wvYOOcr3EoZRpwcFQC9lUnmiDChZI4U6eFl2b
Fgooc6tXyzA/agl1KZjsPHqLxGaS0hqXpT6kQpl4hFsYGKKIx1W1qdiTMujvBspS
6DJ76fwVOWnLf0A/9YPHomptjyDkp4ZDGBC4JRAGoSmdjM52EkOP07Tnj+9ym4Mk
XcPNYsjWT8L6I3akCCmOJstpELhFfE4L5VQ57MngaOiHnwMASFRKTiOajoIka33j
VH7THQe+4SAGu7ZNSD5igaDkk5yFLn3LuhyubBAdZYHbXkkpyr4n8X3iJ1LDauaV
UWUqgRHsakbPEEuj2mu+fovkPbaSLYnWjqQ1ArTRrB1O53trpjL/UcxUgsEcjKKd
LtIddvYNtIZczh2TZFsnihONN60pz9IkWhhly2c82nTfIZGB3r9W1jKT0aBSAAX3
6NIrpFM4KNdoftQGheKhPKMuqxqj4c+dxpn4rNVZ6b/VL2V9tcepN8DcDgOBAqk8
aGvkYAR245EoRqcqy2K4mJ+MykzOjFQIHPPn9ZTlIkapHrrQSOW18WD0QBVlUHzq
rU2ag/Kzr1SRowoc3fSae+db16ZE+p1bWJWis/UTsqHpaLs1anG06GJSPLe3FKLZ
PZucV8pT6VAS6dEouUdKPj6wu1sR2EpAqaAlSOz9F2tzYBl9nSwUAk4EOnIiPWiX
TXhYCAlaIF64YWK7trARZxhY7JO50eQPF8YFtT6z8aOyvmOZ8gfDWHssHvf7fpd4
CATN3lWQYl5NWbj6PS60PC/cG8hTyufvZtxDM5t2MSuQHiWaN5ytt5grDETr+98L
rnOuxEIzqRdj7B0w3zvGhzUHT6Tg6f9TLguArhxF3p2e2QAVqNpvAI880kSwVAsb
kpujGfONoSX6ZSAEz9Pf1A0TBRSnsv/zvB9ULasyn5r72aMqy7yYEz7voy2QvZRM
93ZSNES2a9c/CS2UCUsvDS3CJFaF/IhdXTXGfeTPFvty8VRuZCOFwF4aYpBNLoXG
msP4ghbxj4MfXLoIdywcDIMbsIejyOjEJtuOTxffb01PkJ+GuOA/nysIbQ1hvNEP
Gf+JzqGL3L/8yhU2HK4EjFgTwU4qPlebfg31zNiRRRV4JawPI32XCiG478HRcaux
/C/kVFhlLOp2q6uIu8S0xL/Db5C/pfcB0QB7RhXWoZkww0L30Gntd21otD0ThniR
0JwGi0Ksa1/9RDsR0EaGRhanu2qiBQ27RGN9Z25C1wAdy7u868PU2BUrBsO2ntcw
OohbYS9wcxA6h4vTKxHD5vnhpv+O+mVFOv6T4a9KBYGSE8fN39HOTGLTjxuS7DC0
T/G3C3wbBNRAhU1g1GftodCu3W9z3qDiUqP+GWOHkEz02wNDIuSDKnnUFE1O4X2V
LSscGGL1FK0k5t0lb8sl5VEwUVFvfPB2f/i0aIaEWcdyhiP+d5Rk3wUbNbTTvjBU
77RPljukae1stisHjPYilg3JMlOFMekTO1rv/Xi9brEbrQh4VQLWH8raNxsZgyp4
G+r0rDOxcgQjGdZC+juqfZnGN01nu2Xm61louRqj4QzvvBlvniWxsc0dWnBkF13m
LY8B8VBCcYP9UARPpaFP7MVJgwyqrXQgq2kfOstmh+YyDSQBWognLvwahsENwVfH
r7k4/q6dxC7wlE9EWHj9pQ+4qD5n3bEy6714E/ezX+4CNX5Nl19sER04M58KhqGN
AfD0n6kqCDkbYLYWm1HLtbIfFxdTyf3+GE4410gYfQHbOE72hFvgMPdn1GY8XXin
UhiMH9TnvMY16lFjBI0DAusLL/R+P8G8hpitGg+2YJyFZTyjSpUQloFCAAiihvCm
mPnJa3s4Jbx64HdJHJJbvYB6hfvS193Hm40icYI/TtMohQW4QBzXRJvSG16Zr6ps
GLn4K/4UhJyL/KAg60gPQYl8GaDeSYfHs13RDqB0TLOR4uH+fzOj16dcg9yjL2Ne
yy3EYbs9aDwyA61GCnvrwP83HupJ5uFKfumGBdvaAmRn6iQtLSEMwJVB71O7+sXY
U1NOm84DqEqdyRFfOsWxoP3GBYS40UVoEcxeXBl7hxteBFT/kGLKLjDxhY19Xn57
c8msnv0KaeFxupW3ZZsp3y/BahRbJm2qL9odbKS5QqZ9ui1a9brLWuWLmq36U4Z+
9tCFqYyYQqn8hPOC9ujB6f2fvTCc7CsrCafA49jr/HDBFKlbRHppo56q4iANF0MR
1JLFsncDcTiSM6sEKfga6mMItrhKOajuWHmLxYJCjMkpe6OokYCCX5dBpob3EvJX
TVEYpGldSNUmTqs8o0fBo31/QioyIAm3jzlTOvzO1CRCpCGp8FNrwhjnJfvelaEx
+55B8eh8pVAGVN3IXOAm6oArU81+p9/78BsdPin00oXGM13K+Hnl026qq+OolToA
oWYkrPH2puaqsGoz0hESbdkGAJztsrgwUC4FsFCZtTCQG3P26Zz60KY/UF/Y+RK/
qITQ0cNAdNdrLbQMHE69Iv9/mFZivGu0JjVDKw0HQI5coEs4XjZ+zID0VlrEF1MO
2uPuv32r/aqqzv5vtAIGIw1V5dB4uPJF8bchINawKnSkR7KsNIOF1W9ExoRTNKfH
uJ6huO6t/HsVLa0pHdgEhEKB0wR7qPaGBkH2DyogrVrtWfiwIdCIVKB3XoFkDZDq
JuFn1K4R/M27/kntGLIJ1g0nYnNzLfZn7S+lcQBdHLlZ4z91KvswB4N7jNQ5x9ZZ
3iBHj3LNea7b0TonXQ2BxYDHornwiJthdmVptCgzX+dCMud0ExrmfO8kUBRYFUyc
dVmJl3FVEylGlaLY5YWTo/nCKVbZgBcjvdyO7/HHcEyfzbpvdPQbroFQaY/CewSO
yOANI/LpBlIWmQGi6rZ5j4cXBQBVNg+bvUBcCqFA9rq/wA/Zj8tsq04tdC2SZxyI
n50+CFg6ZYcSPkvZ6lTidGcSRmZUft/kOmwrT2ucPSkEzqkqcpFzgqNY+fA7snCd
jJztLl7TNenBda4WcbuRC14GOX7ka1eMSRhIsBo7KpCBt2k0xjAb3ODp4hgi4QdZ
dnsyToaLx2w+gxxi9H6LwCnGSu+WqISvvuNs+Q7ETgADXTXrlcJGJLkqxoNjg4kR
kNWQkAhsNqhZslT5qYli6kmrB7jtGytGzMXUL+AQq4S2dwOEqaM9e5ybIlc6MUho
s3+ZRGgPlXfBXuCajsZwYFT/g/O+A9YM3Z1Lf4eNEjNiiDyMXKcRSHuu15Jp+QZX
FKribsA2fEQxEkaD+2W+bmmsSVPmIA77m4hlYS+2nf/xFcsYtj3kxRgISNLRsj2k
V5jA4CBjBggyjY9w5xAkG9yurp1VTy0KIurdJU/U45XlTsQ/AZzl01XmljEa+G1y
Q4Fn+egaO6fGODukr1rA0Ijz5IbQFKqu6mBe2+2tN3NxAasft9WJgW6ebOJorCjE
g+6hjSetHUJaO/15R31sgL/kdnCsq0sHBvAxHOgs+3Y=
`pragma protect end_protected
