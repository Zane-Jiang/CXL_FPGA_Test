`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
drsbAG+/0YL/bKNwQ0NtyiNQNuryuDSpJbRou+k6WAGXH0cGdh07SZsWJelEvCAZ
jNpY1HsUOQ/tfh1gfUEjI7HQh36s3SIGdeGYILTY4jL2rFB+5khePwjnllv98E5c
hkkIS89ZLXGsUZsYh5MYSPFdWPcOaOz9dtcpuTzhHHA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 31024), data_block
+2Jw5YZ9A3dSlHIhDDuZmGdGVK4aM2ZopYjBtL9RyAjsYQkBJw1VPFE5K+ODzlY3
O44lCArVriX1pEl4Pa36IpR4sYQ4zqo5Zygz+4vlBuXQXjJeppuyf03gQZF0tSrY
ofmS93aAL7lDliria7VSkW4S/AxCgV5XBoIMjmMOMhYyjPmX3B8j7+LNBZefj612
b0Z2+C4mQx1b/h6AkFk7aGkqaxWqk1IBaS5xLKbN0pINtkhqg4izusysfcIncxKH
V6mo6CZrcY6nIU9p72nYofV7veFu6T+nKZDHDhxzRl/obVxLefcw0FDoGG1Hlzfi
t5DBpLFp8jpY0Vxa0wUgRCCBodnMORDK7lzo7ANzQuX4xwBtxoOgu0T64gHi6QcU
MbU55gS6ZcWAcLc+n7XJhKjjdaBbmdz2kMqQcV0dt9THBkWT+iqH3/vUdKSiCxES
0GgXtVcUiPWW8wSd5HiefRB32XbLppm+T1Bn5/pwH0EkBVBsDhOGnstAZn9oVSZs
t/0J9Hs0rwtlcuIFZtSRo4/hGiV9fLTu4V+e53HQVPBDWlP+6VE1FNcH+MNNDxU1
uQrNs+oJEAdTmbwMPyEXeQ6hgLbkfGGuBBYN5LN5ufYexTD0dqVtiG8VCvzPI6yG
5gHTp6TfRe/b71d+XNCUtmcEw9B8F7O3FqmLjFxw+ER118D0z0ifV81GmSIjfpwz
Hp15e7oVtLAZ1HnwxHU9UwFXHzKlsuRGSsbFdXKlAqp2IPE5O9sDGR/1k5Bn0LXK
6JEAkslartyAimUcxFxONUw7yTajJ2A4lEU5jxnMXGPvG/CmjDIz+FysANXwL7yp
XBQlE24juTU0XpKqAIu5mY7R8hP3C7POF5bJ3MwOaXh4gZmE9jWTFrsO6tC+nEE5
seZZPQlEswUs7AZhYATKJtHgJJeiL4uIgHJZxjL5MgJx+SpE2y6WYSYU5RkCzGLz
ok9nYWmvxTdT/wcWn9YW6mFu3fvgywslQvgXFJoXIex0f7dADjrdRklDPlCGUxjy
4jBnCSByqIn3T5zkhDzOeGPCA6KLjlLCw12NHZolNuxVbzJiR6feeZsrNEUbGmVY
QaJaUNvr2QMcT3eOzQnBoS+52JsLx/YHg4LXcjkNDCJZZyzajwaMt9vqVYWqFiYO
tSn427EVAULLpCWkRUdfUq6c2l4JjYvIHiX1Yj6E8WNp8ooYqvZmzZ8OKx7hfOai
I6mkMCRDqGlJqvsuP+2fDrHpZGjBs4nQmSPmrt+hbKIlkMtlfma/6ceegF12u7am
ss6rlty/yWWoB6EDbfnpYuAd5aF1lBOz+sbuqW+v4L9qPxXw+wLKKo59UD9nvM4M
MvIV3+ath4jXffMwghzsknRAXSWR+4acixtXGwsTvP3cOtdHlyCM+JDktWwPbg0c
fkUPjQ8/n4+cHPzIlsOyyq2JEEeewwQ15B7HDvcCDAOYyXcu+WqtlHCPZDFN0CMX
qjhCVQshpH2LsU6zOCywPWbbImxrgASustyRcr+gQrh1WMbRjIc6gY1ky6xOrh5m
WUo/hlEkfo4nV6yDAx92jdDWqhX10HcocknPzQ09ZrA3cWeyZv0sTF2ucwOomj/G
yb7n0c05Q3XjmSEbiXGklk5jheMsFmQELYoprLKbmxNseSdqPa56E4qGQgDfSP2i
zit7A6/4HGYNQfjX9OpxrSpXKfjgHiSDn6sO5bhfhtIlXeSz3R9EoSl+38oo82nI
ELtMbfIzlTprbdATOPhh/pkUlDJm3xZMCFVnWNw0Cd3lMJvxpKHeLgWe+EZu3r9E
KMfv/u8PHaAZj7SQXDotoYJNEcFByM5EaUfP/f+UGzTyd+eSVBgS3pVHFVSPTipg
GE1dK4+cD57YdUlwFSLXuJCqn3FYDajhYnW8yYJQP8nckHkNm3IRkg/ATdL19ypH
9RXpav11j3xT710bqQM7e/ypb0UgT7S8edM9YAhhFr/9P/vpAHa3fbUplfqMYr5G
IvZKk8gwM6wKQH/NRp0KuE3YDJAypO/rormc9z7qqIS7SGFpVaXmT5pUXa6/hsL4
V6BY3eVtfsn1BEU6KO45gg43so1+IxRWlqd7SPclqYkDkhWAN5OxczGN0zmjILSj
kVe3cqGQHJtAHuoUZKurs+ta0ZmkzZS1tBuWIwgoCECAhqw4MgcbHYA5/dDmC2yT
9OpTrz641JWo2zu26tdcXRS3OhsiCGjcxXhMDPTi9cIcejyhZZT5DoTXOK8CWeLU
NQs57XfAiXyDB5ioTlzFGrKHc/jhad2dKeVp2X6UNH3FxaX8oUR0uTiLY16Rp15L
EI+ReNDD39voLB0VQEtvcu5ZMx6x4cWjm179mq0Tll88TaLdrGmIaYATllbuSnGm
trJL9MaUjjl83nMv0oSJDlRW8kZsWBI1sJkuRrxXg1rTvYOt0uETohHUanpJS2mz
Ssj/KJTH44aPlur6mkjC/oK6VvQB53O9mZaCXz6hsNNeDuCEabnWqtrctvArVDgl
Sc9uDLCd4l+LgHv7OC3MIRi+wlMsc01twDSpyKE3ineCRQTBFAuOq5bhD69YTAJK
U4FARQ/ENKOFqMiIR5YL9vZx9sR8B0H7Co6Kzbl+alnmjCwlhuommwdwHaatUnCy
rgxCyuqEGoW4fQPDVawj/6NrZcvDMJclh8e1mq8BFwhd/Lp1zWtp6wTbdIzSbIlu
MReE2+Dsw8MJ2gGiETBzvMXxJymKWTayzReF/V3iv5eC4Llloe3pPn3iC3Yy3Hyd
MkJKFypXU7/ds2kQZxmbOvT0uhq5+BkAdFFnIZXj1x1DpGsMKjHHCy5ZlnzM6tzw
w8I67nM/dxd8q46ExGUpxbLdiZOLoAg8vxBUB0M6A8YN9+qDBxQFrUg1GqcOVmpf
3sKzpcErkTs9d632X8nSqiISAgnPd+fOzvrTqyNzyPS4Q+VHRY6uk4bGHGD+02FO
gg65M8HRBbM17W9CuAVfMfjEcwAzU5MYvLwWfEUvEe6gCQkH4+oMUcHwV9tEvtaJ
RmokP9lWpMOWq4SYXr0NhDJpG1NRbNN7sqQslNFyyCmkQdbT0dF4FklsVfA3xG8h
FlGr4HBjn8CINcYrPkNzpOFEMQkob2VJXRdLMfPhBV6zM2xXhOqObfFKD0HRFjSn
nSh8vo3EyNTziXvKNLUhLscYRzZn608yGUcWmqvpSMAH8mYifM1MprIHHt8PJAkn
8I3m1L4Dmqx8kZzeK40r1AELf5ItZHdchRUwIUqI2SoPB4eaNOmuX06QL3O6X/gJ
EIvLm/LWPuTp4xKqW3ppVjh8bKfN5H5Y+hcDKL+KgjM7XQsUz9T5Sf+eX7fe29OK
XvKuYdqRrPAWaMVWlE9hXaTPSqVVUcNht64f5UmzQRpYRh8S2xY6E/Hcdq4ni+m4
kGc6UHxRprlLa1JSq0fBBzKxl4HZfErqFiClQ03+p6fDy7z709Bi3vsodxNBHmDZ
XzhOgxiipSDNWQ5p8N/wSSPxqf0YRluASLpMfPjarjgbmEAJAsZ8wYH5mFLk+h1D
aug9YBJza2aRkBiH3ccXAa/BQiWYV45rNFMFr4nnivgm/5YzMNQcqagbBuQiTRaK
drkaxq6Zykf0dWWWZrhlMo6WHZaPNmDkdZkVeRLqNTrDIv300gnlokY84WETxirY
Gq6y+ucOnqpatayW38q3fN3fa7jGPn4Zjp13qQggKTwTpTjK5gDiDJoW5qGv4Ws+
GPZCOctFKDanZIYvOJMvnsmSZeF3Oog3PBlSopKUSRoiKblssEm8B/hs3etgiQbj
uqVSe6FX0/R++gMzFPZEBum9tlQGImMzFJltG05F5/u2xOjd4MNJW3QNhM0i3Nv3
iJfsb1VhAG7P+amM+G4Y2Rxg/I48c2i9E/HzaatiF7HbcOWsun93FkZXYLCv1+XE
26yY94aPQKvfgzVafh43n4k8dF8yvHsUMdqgV6/S81WSPcX4qYgGObfUXd83tcKA
/q3qp4B7GB6/ZwsQn17hsGtSgWnL5eHa01U8vbk7gyCSSJqg4fZtMTedpNL8lZCU
FFvl2JYJJsNvDBx8F30lyLvQTiAz1LJjJiNiwnSyj2ifWypt2dMTANgK4NbePEWx
ErP5W3dBs5RGI/AzHKGO8v+dzlfHddO5sKc8Qm06Yp04bEb0MVr3mVSIlqnYiDWc
eNGeE0PM6AycAF2/zm9gqUGOTUz/2ZyDAMUBZiCvINHJujpiTnsp61n9OmG9tr68
FoKDtabJeMuDX8YRp3SW8ivAgv8W19WsM1W5CuiUCyn7KplKx8jxJYf+xOjAto1I
pBf6/quQRE2QWH8Z76Dhx+EbU3FIviQRPq8P6+FzJPKid45oybGEykvA/6ZrQDi/
sJJlcmCCiyvX46RTC8P7JsM7Hx5rSOod1987IZXdrjnmwwXghVOcCsbWtglYRh+K
wVL3GMV93HAH3BkRsdU/1chX5E5FxtztZkyXHZheIVNW76DPnt2e1bNSpJFYBLz0
3knFzw7CrI5XpwSQIiYoNe38+2eVat0uY7I5Zu9ubM26NJqMjJM2pWvYQuruV9tF
KO1FPAgthHoigxFnHf2gJKUmBbD3K8NyYXfU5Fc9W+XfLJjL18js2+p8XE2Sxp+m
5KbZ9V0fq0Pj4AaDHJAl2xfZhlyLqsvxNiSdBNoAsxRnkHlu6U74JaMivY+qfH/e
6HU1yyrrHj2UuN+dAJijz2caHmtJk8eeW2kFvkDTshtA2ptd3Y9MNoosgbtRgTqx
a5OIGid8ElmxlN5G7PQvIIOSyLE1J0iXVtbMgprFrGExgSriPRxVs9NefAh7bwSc
vDFJfcVmDJ+UctGZ0xlUMCFLKuw5CyKO7axhEHxDGX+LC3ZivLelY5SOga7+kdek
AawLHAnk3b5KuU83JMh8oahQ81FXQTNjs5f8doLtdIb+h5wGzFMZx1J9QibyTm53
IPRHiK/Ac5saffFReIBZGqQoJ+LReVQLGukHiDhlQj2qo714gf2vFUJ9DcFFLyQ0
BqRcbG9wHz3X7TBfGZpX7DT9W7m4x4NgUD/zvCvTvip98fvRzNzeiSIhw/gURRfk
k63K75I/15zqX4oF2s9MSLAbgeU1Yf/DOp+0FiwgL/81utjAi1/J9lcyX+5mr2ho
yrHlQpDXBmt9tLHOhF0cnu8Yoo4QcSM/HhewMXdz7k8Af+5iwtH54jAwa50/yADV
s1bXHfTcbU3eV733BUwgCP/hHzcH9XVKHPAY20xwLHEl7pBfoTksg+WXa92Oe5VN
YUpH/br7oKYmJXbA6nVbb+P1zaC7ef756IjULPYCLf4d6uggYQwC0SnNuQjdgjjJ
qIpwyA0uliTfMZ/+8PSQxmv4HR1A124qGba0DcA3HToAT4EBlG1BRcVvT0UgMLQX
qfwkb6WvItkiSD0nvHT6ZKG41syosm66DA+238pIQl94YhC5w6zx+05Blo7H+AVM
o7FfP266NuueRo/gsqhkenp3fkd+oDAC6zEB7KYoJHU0E5RsFy0r/BnUSUm5qNLq
1PdTruKxLnrB4Hw/oxWvwm2YrxYp+G3zQzFAdrM8sXQk9EaVnMyBmOXKLqvQg4q2
y3Ls5egbVSlMyo3n9OLNdBJokoH6qnb+r5JWgE+gSh/wmrRmt/9mlFz7BB2fne4N
ct69x9lSDCPZuGgUMCifFEhqKNnGDNVaGk6d4JyDLmM5MtAm0odowU5Lt5gnunbG
5zz+taBkWvDY2pW2fh/3Jccc0qjQbpdbNl+tMckLGvarKW1uuR9S4JV3foU4rjZb
gkMuggXz0IjIF+jzopVtffkBPUSG03hu2H2CDXfV9cxpNKS0QfJKHln0GOL6EH/K
8S+V20mynmkmSZUfmUJ7DJDrlswwsUd28s3vQ02sKMeOpknMw2nd6hsb1k6E30HA
2NYc9F8cCNpZ2CSYehaCdpXqAmR4Gg0HNXz/bi+i9cT9r3WaVKRk1tH8K/UpI8B2
N68BELkWA43ffOTWhqTAPvVhxLSuBw7mE521HDYQ3Z1LT6rPM9pbX7Jck594n9SW
fmKWoxxtPJzDu0l97bLwkmpemghghBPloiPNwYDQB6GjN9M5o/JIQTRWSvMm31pd
lxguVUE6pzWjPv4ICvn/m9WWHWII9/5duCHjP0OZGBNQiSaiQRdmn3VFJ9sX6dWv
hx9vvLCd5ondY5GzQNplrNdd6rzEdEOHmTZHkwLSjtpneWsuXUPCfrBj9Jt5s2+U
AyFcKT6n5+Zc5HBjMrIQ5+1cER4wVRnmWZnhvnuyDCULtBvZY9gybijgY4vz0h4p
dzjWRqdyE5ekLmcNeTAvsms+yr8BCqD+yQ6kpOkqAyrJu9ntkP+gz1XEjUSxBlKb
Vmn9lFVZ24pZMIQxLdf8YzooVBvMnO/y8um2QiEM7rbSZec7hB6XbVI6bWcl2o9V
bRvOg1pdmAv4YT7wDIT/yoaLYrwN9la3rLvGNXaZ2552qpMpqvqWA+VtrRQpIWKB
u0dj7kKfsk2Vk0788V4oVqdir/mWi5/DOUdHeZST4DC8small/+AUODKlHFKkyIF
zf+afqPDUEUjSJuMHjbN0gSF9AczH/KcAAkSEr4oK40uVpFUa0SMNTPaoiB8Ukrq
ELsHhaj70Ouz1ALaztnmQHnYvSH3mqVbDtILO0V1EwDGW5iibDTCCoiaXXhGjep+
zncfy+FMH7iIOq8I7g52L/RM4agenHZUdsJasXZs30y3GMl55snN1en9ODNas4RM
BYvDIxtnilStRRFHTXklOuGwe7xqA43jsvJNjQ/YzQxXPEyDfOozNIItAGHB+TCq
jUOyuj+shr862f7ekJ1wmTLh7DHSO51CuyaozJJbmdL3eG2GANduAjDUBySns7Uc
WWMOxPsO1+Ml3sfjvV5HJJ+SrIFvip4vbbBgNqz3aHw4rNxZbrtXOp3FGexoFxni
KLtV676EjrK+DeHVTR0AtzL4kB6HAJYdS64mgFmJ4eapO1F4+D8TBem74ta93KVs
TZMJ+sjE4BvijlUzW8t86ODCP7eCqKHJ/RaT3g3RTN4n32OOe9AUfwgmcv15lnNA
cbZUJeWUYNx67uoucT9FVW9YegDw8ZjDXLeSN0Yw79GTp2ZMTLpI2sc7vy16J4Rl
W2z2VPOdTyE6xT60MiuSY/fSU834YdIIscdEQjnfUwVA9nT3AC4YMj9VGjlQFS86
9gC8Efj2IIoEHD4A2OzBSOSD7ZvzsT5yGzEixscn4iDYnzAqN6X01oDbxPACm6wE
sf9fhM1g8VYXhKHcKX5bg+0lGZRiWgH5faHzfNxH69+nBHT69gkuerDgXY9HanTH
bSD5PMnwHZWd28XXuH2MtLVzrSn/58YkOqE6sv2IPPjbhGkRO2NVu+llKYz9H4OT
lb91eePokZEntmtW61G9ZC19euEiwkvUE7QzvO7zitBFu/U4VDjk4PtE9AXF6g5M
Z6qs5CCVJ6/6ZS1MB7z6MHjrStdoS69hcS4T5oTBWOda/pm+coXtPA0sySuItEtZ
1pMvL+Hwd+phAi2JoKC6VJ6RyR5k9jhmughEzr/4n739W1VSTmXVwVCNUih+GzGi
mbclcIiad7/IU6+4LYiF/qG/wJtHwnT31kPIKgRh7n03Vn5fIbe1nkToWqVAZBvT
pIJauApDTCYcPZrDzyEiLbLjqpgmKhlJ5P7smjjLf5BVb9TzBu5mQKJ7lsVuQVwt
EzfSS0MRn4kkav4U8ZqCxgVWIdk6v3fjD5x4rQt4ID3SqxqGI7vsAJGWFH3NyfdK
Tsw1F2yodTE+QMP63q3TR9xM3fVBlU/NF7AAmmW8EArSm/zZw2hd7mk7dmWnHXWo
sXDtdrP+HE4UXZ49f3tnObPMdu8sfFuD1nrm4dD4x/ivlo18BsX5c4502/73YWk3
7pGT5yvNWkZ6To618Lj/4TJPKl/BE8/P7aeE3q3wUCPIYZsYGwnTDqgFcSRJxefM
bYLvxxA3iajkzC/rjLt12QC3EASUvSTsrzxc8z09V6rIzCYA5cWsH7/5C7nze9PF
MIES/AEobF3TNdsvwPhHzAlZQlsJfZtmQkOdgGVli0WWHVIvRh0L0bI4UMA2Sxka
nhVAIgYW0+4GV2EBrPoOTIW+ZyBcB05a5kPyHNNKx08cpt/uCe72qtAUAwmWQOpY
7sM1Yo7nWH0SD70MiSATjP4gK635xwHIMPgE2l2IwtM3+OaaAegzefBVCrjQMWvk
YiYbeBJmd0CgJc9pAzxmI85D1SlRa3in/abnwvQkZR2q4KhFTp9TjphlQwoiQzZ0
bCPHE3T9HByeC7zjAXz7Cnnhb9DQ9y21wq7WZcIqnXG613Cd9sS1rbuNknCizKGt
zl8f77lyxFoYMOupcXbuZgcsPiW06uegJZ5dvxKNWnl5AVertfLkRPr8lOusO+yJ
sysdWWfHEfzT5xxdog4HfRG0O1leumHtX/vl4L1Fufm7uLWk51tnwPEX0q/MAXX7
U9EwKYhF2fkWCgpQoEshaV3PPag5nVS1GWJt2PLoSRQOqa+9raUGsZYGT7kIG8bE
peR+DpyRMTLOqYK3Nmd7TgEB5r0QmxD0eHG7a4MOW+Trq4tTulyeBW1EW8ubWned
O6gHeSi4t71lBxy57TDEkgadiqle9UyM8M8ncU1SZyvDbBnIPj0AK5aE+Adbc325
U5euq4YW30i2EQkf1xNQaL9zrOOp59Vu1lwBRE+t1iJ6oOBNHhGl7oCZyArxhXOZ
fEpzytguqxzb3WVxEdZ7YwnnOlzvaABHda3SS51UCHDC3SzFkLLDR6ooGWPXCAHR
NX8GOQCMO1wTzZ2y+G1DaMXFu8y+rsBo6njUoBw/cXOTmxpGcos7n6qjUjL7T74D
H2k3nEvz16pYU6sqkcZEhHfAF1C3JBRtzEVvLxXp2QebkLpQVT++kuV6ND0LP1Sk
lkEy8lipMpkBzHGalHs7mqloIGQr/asp4Fd2gv/Dq+srqYagkkvX16Q0KbG9Sirz
mJd4tfOtQurApWJE9duTptfshiiPLK7W4UTHjQIzMwspWJqK9YzE+bI0rrBMwsZg
r70kAUXtgriQwDlIGSuPxWmjnGuA2fD+nBrzXYkIaAlm+c6nIBNHgRWPC4YzKgOd
OcUj1gJqy8BbackBnLxmZLv+JwX59OgQ1PgsW/6b1tZrtGVbgacT7cqJioumK+me
pzhyrWmx6hSAgkoMtgbLUDuWDTknQIAnmBaNpDUxIzXika7RfA6AyP2/j61RIG0p
IsBNKEvKnr/CLmVJfU4pb3nMpSZPbCwnLiElmW8YJLJIZ+YnKxJD8jalvAtv184y
exqO6tywlzM7We1cdeoVeTyRWutESId8U531gEQcmOVawuncH46ez+JYswT7lEyi
AxwH24mvaRmSs0vuiE6NU4tfJ3sxZaWaFaP/NQ9/baw8CY8Q50sm73GGapz3QTkW
oJqVPHTopmcIT0wAc3tcXxbzzeY0wdUha/keARGVcKxWJS8E/HJ31KuFoBSwe/7P
CuxiarcxxZRC6vG9FRBqV1uwNd/Xv/Sgu34XnJQY5tK8sEpDePDwD31VMQCD8x8m
+7Vla1Ktii8egLxQt9AzFw6qYw5lmQFmYo25SGKd1NCBm9wzE4i6A7hnsb2s2UJ0
SirqJpAtSFgfDBnLh2mSAgNhe08iGJR9AIso7OP5ELzSfd3A2/w9jTUlVUYPYOfC
amw3g7bsec+MBhSu0eU7Uj3rXM+1gxHQAZmNPxOLv7cd4MoDNZZhSHfqoYUM9Bup
6VvqefQXkT0Ej6rhJV6bSeldIgP/j1R/i94VlQRPctHYySIC75BS8Pw6n2m4g61X
dXizDKTx2HKoLOoHdEcGTmfZNkyYaTLeOJSu4NVrSYsUGfq2Fl7yqeSv3jhW/836
WZPcFB+ZxKvMfmJNC9W1pa7KSoXhygFCxBsXFlPyqWBE4LZYywj3BRm6Qr8ybAln
jeVd9tShURDHOf0dTptqBBuwDPmlRZ05IsatlA28/E50hPajjkxZveU0DBCvU8QO
jyC+aIlpSlwfWmdNDJJlXBK59EQHSdAasl4Oom2Hemkxn7jO2XalCqsat80MgouV
D1xwQ7lg3H3vXnsAwzxfqFxCnvX6YWPWX7mDvUlwQE9pE1WAq+ZMcWYbPb9CTKip
CV9UZFS6r5lgIVcT1+gBgrLjV2zBIw0YKcaSPXi0RIdayMSFGknxVHyj0Z7MEWAq
WApbhxx+7eDaLl7iN7tNMcTFoPuUcqlbYH616T9NcVSgWm3PH0O3iGi/APjHHbk6
TrkRUmHgu9en48u0CtHZc1EV6L+1fpvdVrvMSOTCU6HRaPvfRv3TsskMl3E22ufm
genWf5LbrpG9qVUhz7G3iDyHjC6L/LKuIoYlJjn5YTkR73ZLETxMQ9q2Err7+3ee
3X5zIesxEC06X8dA4GfgWZhr3PNsN8PYDrrCEqeMzQQLfNq4WhI5XT/tVTJCOq4W
xUx1ALtIjfYNDqA9erDBLyaETDN/SuIn12TuFFAmVaIeYK6Wcqqaub8x/kaTSiL8
YLARS3Wh+pJFPpWTrXk16hPZaEnQ/11tc6Gq6Bl7QmluBgvroJGIhFp8/yKf8iXg
E/3ZkLanjO0IfbAJcnf5yuDLPJ4+udWGL3lIOG4J23I+F9kkISRM55N2vhBVNcCj
QvBWiWoRDigoez9izODpxUR7spJ9mrzflT1ERhb/CYM5b1dR0kBvDTXACvFVAfze
miB7FYwpdVyDatT8blNrWya1tfS/0yRavsXbkx7zfLty+VWSWuuPwLP6KpcK36m9
cx77kMw/A7OmjsarNIwfdFCKqtwf+73neGtBxWO9C68FIx+qvns6yW4twjL+oo4M
rTK0Elv1B1v5F8KfimZ7F/CsQeXsQt8nzsFO+yz5CMwssamoEIYbIpWPeDmtzwrL
XMMz+gbePSxqOAICCZu6EvyLEhoCXu1xAjfsinyQS+iv7ZvLSPcZqdA1wb4Go0t0
ua08bVDqlvRW1134Dqtviu77IUw9ctg2vbHJPgqJEiF72GztZI935tLtE6Nov44Y
9N71Kei7XhzpN9RESLFFMheFD2guZ+Jq77wIgmvGVME9Uezpwg39I5F8AakFzAuB
G4yOjUuvU09l3P0AHOesGoqCa+w6fDGBPTsfpLMV3H3QEGG1rjYXV5Ove8S3/q8w
tVKEgVGAsrS0gV0aLi81kUj6+ihXYaAksCS0BUsj0Fqh11QanTKRy2wZKxmr6TUY
qVWiz7qyupEJ/vQb82F07SppF8N/6l6LKbuftLhB70h8V0Xw/6DU5eGBb5YKbaBo
h/Yiuxl5pdJ67jpJYg1PWzY1pRIbWOyRzD893VvHnYeHWRtJsAmBXCeKdkdzjQfH
rvCiJC44ZWJ/gzykSJdIouw+gsOH+8E0JMZBXdIlf3JQVyNZ/NSi4p0PEttx5kR0
bN9v33dCvQt3EJ4aEgyTdWZPbnHgyvI5ibun+3v0Vrb/AAsdW3prcMvBVk8jfWVi
DBPI3tww7SMAAIYid16OKKDRmsbPpr4aPar06/Hlvb7SAWdCeu/0XsiLqP4oKsmO
SSQn42MWs08N+M616g/s3w/lR0odtjox/RH6knzgA7+hCibO5M0A/VM+cNJNz8He
x3Q9x5YtDFlJ5X2KmEqB0e5PgpWR2S7NveMYtSg3ZG3hqBN+xQP6bj+2lvVvtQXU
1TgZMbiGPdz4Y8dljOEOpmB/vp5Cf+bKhuEq0SlNVXvu6mCm4UVqWvaD4wtASxz0
Y4dAATZCqx8IXayphd55CMaxPIQOOzN4IwNLkshjiFHzOSzBz0Hm9TnlfwxK8fyu
JqHq6dAo3FFGZvAab5tYlaQBJchEmwMqFBmWmEIbwVhILXqr6jFH6/RP8mjuSTJz
6FNwfHchqQuw73xq8k7e3W/rSNlLKxH7anwgpstEWul0RbMPABLggfjjekqyH47O
zEwz3g+CN8cioLOY37BT1CYAlQF+xYnIldn09nBWCfv2lEmQrx6W5GaV8Z40MpwA
u0oGwGQctvSxvl0vU4Adj9LnTVw8jnv1FT33UyIKvAztqn+ore6yFuIeS2l8j8+J
G/dIPf2hA9vFi9GO6ttNYtksAV6EiCNfIVfmDdE2DeZeIBnLtf3gaoReWXZtTKc5
NcElOGBpDCg6ouXtLqvpd4rzpmObqMsezML1RtDvAvUxcTYGZ+DqD7tFYWwxpIAT
9bvvkLcQ9nLbHsNFm2RJ/ovC+DrfM62I5OxRfNOT6MnEgZRaddBYnpaEv+cXu2vJ
fHq8HsyLidsgZxFIXOMmhUHxeSTEfyaNb00FoxJa0VF/I8H0ty1OQORletHrEWTM
qojwp/9yYXVzm12hSNnZKa79gvjA8+0wpgxc2Pj8DIkdKXTFWiVedgBdMIaPL7dr
QeV3vQFGGrKeBFgnkJe8SVIb137NjL2WfxCeKCd/xAHsQCh7mEKI/5k7zhrKt60b
/rLEO4qdqwIEg5JR6+PHpacbTJKNySLrdzAiXnWb30O6w948/2hsgkpJYIStyxRV
+/iQPlhvjJdYm79YWkPTIDCaztlGPC3+JwfVubdmTlpq2qKfH3bdn5S0aTzbkcC6
8QXesNUwdZiTzN+YCoavSKjB6UuULafLoImRnt1WWJ+BrHtDuI1GscUBzBokgi2R
P5tZYQdgHaBcdmQkmebfkoFiPuKYGtaCDvGs8RPLxb7jC0iJxx0JRvMsLxgMbf6T
b3gX1HMelK7IowLiqOI4WxjhYF0TapF91BLB/0gtKgsZMuwnQVvJhkKsIO1QhOHS
lzUlJuBLOqPhEEgPPYop64y5YM+FLQuPltMlvR/NtJASrHhP/mfCsYc+MFMRrNeW
bjgOiZKLRGgArGssV253bRBN7L4yLzUdg+UvmUpfKoug7pt2bSPaRSUqDUlobQx5
YpLUMHR+TJ2pnBdkB5UyVhg74122UBKZERa0vIpcAL7VR924wWvLHsBsHB4lKcvX
s4tubRyQp2Axa/5GacJQes5mvl3ZkIJ09b8dqjTTwRQUGh5ObseqQzCTDgSIdLeB
hZihvbgp+oyyGX5idtSBbIDxwwW4a+9Ss3LQr60/r6R4qQzECt4S4wFLP7jTmeRz
iQz4p82GP7oWs3AXyo2fplEB0T1iVCNRccMunYYknEz61NNdldf6zZZR3r5fPK9M
/HFKKP7l9NOck2QjsWcYIJMS+eXXWo6XdHLnTdfFOelU41nlC1FTKgdUw+pMFvEN
GsqSnuMYaKQOwXI1J+aXyeym8BJgwyupFySCut54Zp/guy9KnXnNXI2ysjdul53U
9MUVKySgZZ0KgLImwhZZ/x3T8LkghK59ByJSzQ3imWoFTJny6P9UTvVb1YRrOx8G
ARVg3C3LH2zemvQrVNKzfRxpE/s0pYLENLeiN99/HgRimvKkZuDBzxYOobb/x8V5
dvaJM1Lr9iEPd3tBjUMVBKvrYu6ab4Gihz5IwOmDcyxaB44bmGVHx3NoEofS6p2R
FNDAHyK+xbK88FVFKqLVtbvToNRkCWadw5BlQxq40hUBxL9m3yxwNYYTedkAc/gX
8dpFoelhi1EQjLPRU4/ZFc94R1oGh2N4ozzpZDFi19Vk/qfSTYMUQdCUmPoqiG3P
STs9lWQ0L9Cm+H+/BQ3Oz+Q1j3RBn2L3MhPVt+KWa1KS8osROsKhFfGxs7VAljpm
oZNnCtNBVlPugB1pfGMMYiIVXRleciI7Sf5CmrOP5MRocWP3TVNs2zB0nTog6nvi
w9xJMrluouTmzdvQu7JPeZS2+WdLVLo5aDdwSXKMb81hRj00MUWXVuxq3zJm/5QL
GW9MLZI2CmoMkf18weoJRf+LQbScgL+OC7vP1uPxaKOYc2VtqCjhlVPtC3qKTxts
xKm5EkRCd7kKT9ytQtdTG0X5Fc9SxEvpcHn1CNHIEbvU1gcmi0Q2hXnTemQG66AC
81xxjtaReuOWLaAh7Q+oYrJA6mdXUJ4mnz+7AMv/gPF1ogYTvbarZfJyz0IwrfiH
QBevzPODlVAO9gIhot2igfNncPe236NyIKhqSM7HE5hO1qgMWZ0lV+OhCnggcA+/
6J8thLlsPhflZZvobk0kYH07gOuZLqYbnjTTljdtGtiS/6csMYyK+SjS35SyqQnr
ZmXMJSZefloa4e85bcbS4fM+YMM2x+aEsrdJ7TtO1ucaIyMuO952q1rBjx8W3Iqu
JIi7qDD7o+fFKnzFCbpxNjFeMcSE6mvaW0kQSWIyDjyyqAaPAxgQHzv5TKibhXRU
fCJ0Ma8MHeIUYnEMEp5Nu8JUXUM13SGs/UbzGlASgK76Si6BY4lXrpLYp4mDBZZN
EuQtj0/EAoKWP/mlEN7ITaICHOMtF/WjXrcC3cPENM0ynqSZOULinQhIUilVrrpS
NTGBFtI35pBQ4HYzZo0uOiCAR7AEkXTbAcCbssVFsRQzDVyMHyXSm2nMqJI0yxPt
dcoq28gWjc7Dd7P63qZFooeapB21bigmtj4YzmoGVpEjwT+5oXQ2U+C76nZluiAJ
G/GQrSp57fySWuO7KrT1Zi9ZS3IdpnUtLT0k41hSv+mHuCtg4NAfTHkuUaPdZ3s6
2673TJoAdTt26ONRblWlB6w6PBKSP/ie9+XKdEuuge2R15F4EJGP73v9qFrHzcLH
kzawstvmqk72lLYda87JuENCCMWSOG8VV5VDerhhrNAt7t/mpo3jGqo9aLyD9wGF
tSUXRXqllvmQ3cZO/z1uNiJci1MDNGjobDd3u5xp/e7ZLRO3V/ddp5ZW7c7ogfVz
yvkGq3cBlFD8IoPdo7oyLKDUMwEPZA/lvc4T0vFNVrKBiucukv6x6s1Bq4iUJQ4Y
lf53mNtVVIdLT0tP9fW1dUNj/rmlfH6fsVUAkJpHVzreTLMJouSf9/vAH1IBFN4c
TqgXV1g6X7yYlcpt/Ub28dk+B+PuiLZEeVA5L/R7wWeJDhP2mUQSQaclXDL9KBaL
A3ZY+YXCq7YAuQUgeCoh2MJi3BxGQ8sa47AAdyX/3a/0WDlwY3XPLEaBtrIzMtrN
yOeQcByUeWEunz4rBgBsdtFGxO/36THfAJqonqG9JxIqqNv9JpMfqKYoi4ZPLCNJ
jNnkfgoFY143zz8KmGozr0uZdrMzmG/6GmpLFTwnCm+/+xNM+JHrBEvT8bNXfvcq
f0fKkZP05T5jy++DmA/yJ08/wjPD6DHIroCcKYpNM6VFr30Alw0LLFDRXR7k6K65
TDclCnsfm/9z7T26etbyF9ekLWbG0RfBhqhu4YNmzT/NUq4QEZFu1EixD/jDGpq1
3x6rtsBGVqaqAYKALovK2QE2nLfKX4twuV6pQQBP33yZvT/oNCTb2T9pGqN248QN
564VVfEJM6sb2xvoe3MR/FEqVgqLlHyvB5HK2xyLb8tjCnyC6iGt+/CQh9DrEYw2
Krv2ZwVFPS9rAjzA/NdKNNaME+O/g9CzIf3tR1r6o4dQi9FCBQ1lJQfBIWeYPQT2
i4jWt17uevBZtVOMJVZq/EuNC2CTHyziLg2qP+DK+g009HESJrdQaVxIlaj8gAPJ
8FbUqu7qJm6qnj8tGVrz+3qf6D2Wc/9nLknPGRqL7G/oMay7CK7Un7AtxJdyvLlE
VDUim31wYtKownCl5cmf/EP3/xeEh1jAROroWQ5zfe3KoeBsBST+d3IockbwmkJ7
9yO7YQurQFdBohWCzULua+0VtKbhMzNiOgu5QzDMJsgpTUCVcdu9tZ6Meb4cUCxY
3BIAJNGB8Go8DpZSlvMotaEux563Yz7ytiYkXRss2Mi7xzowc84kP5QiaARo6j/O
PmED/wZUnfaFuZeWyMdi9PvnDmmjR9iW1h27zEzjUy3EISCDyUHZK1DsJKxIDBUL
JZSGcWekuqcb8GjGhVnVx9hTjrTinZsrSrWO16bU5yoTXmfQi5WW8N6VK6Aqv9Um
yvUkvslrjJtrNxJr9Lb6nBP5Gcti9O7lZrLT27Bdm1LFLAsdQZY08XzGafx286/v
mGcKsoLffRK0OZxEPufUyqITTWk5zwlQasmupc5HAPL9VzpvRyuNTnz/WKpYc7l0
7LzO4JgAWacl27yF27PiWc6VTN1LxvRJLhgWCzSVRdWK6Ji6BwBkE2mpNK8HauY9
NLf4WO01jbj/ZUir7S6QCQPuQ2R5z55miFLrFg1mdGma3O+xp+YxYDsrauXIo69+
IFh7bKjmdeuBVZIYNAt6kFCJ8xgpKmNDdJlHIOUcEJehGl+kkvZC0iXrAeBjBJ6f
A0w6/5hIEpGeZOLIcsafQu1e8aaLEVelQorNlYUZQKCcll5EiFqBjlO2tG0csjiA
nHwpAwTw3KhXf/8CYwkde8EBnILTclSpKoodH7JrbMa21EANJyVjxvAsnL4FsZIq
uTP35kYc8vs3pKGjmH8LEy+6kIKaQhG1ZzVFnEW5BVxlKrBlXQopcDHi9MwAKRd6
d5SHteJBO3SqNM34aCcEf4vSUJhMKBid3N2Z8MMPA9/3+ru8hd3PPFlkH+Oc45D3
31tFZAwHQasfROSTwXYUk2G72G+pTI8wXPNE/XgMrd30UZ+KpVEQYxqpMhDp89Nr
nHf3JGTe0ZoqmHTf4h+DvkOpUeAKG3mhkHw8ncXQUAHDACh8fzYt+nUE6+PIU4p/
66kxLWv1d9ntnGPdgHyJ69Rk2f7ZsF/0T4MVnI5gSNSFMFzUScgtzVVO8gDEdop7
ULtnBVG/OBopoyV+pdoJTXWPWrbWuY6GW6ErnTDjKt0sBdSiMOqQl+CwmwY3IKUg
jkAGEmiBXdRTa/fuDxidOa55Q2zeZRgqL4L+CLUWr4lTJtJXnUvLo0jJ7hcEWleJ
8gm93yrPVIcCwMR0YR+qR0T4rbZo3p/nR8VNe7cdUhzi1j8Ch5T7R4uQxtG1kSgz
E0KREto8CMjFNZZggB0R8Q4+kx2JthnO4dW2r4WR/G2Yc8fuK6uasPc2+nBbiUxt
h6Y7XAou2KhToGlJcNmQbq4lK8KO1q6Do8DKKGl2V5/wAsr6ZMTnd4CVPZizDctJ
BPUQKLpXVQ1cHMX3r8vtZnXV3n0xUeOeiNxVvaZn532P2Aam4eNJqN/gS54q9HKe
KfLhGLyF4mfN0t1pPySBgGRUVcNVUvUk5tRCBd+MEKITzmbMaS99vbNy1QXIuHE6
hYzUKpcnb0sTo87bXo4xtuAKmDw/1AfNswokXGX06X3c32scRb6Y0lnZVfTZq8/K
UaQItVUXnplT9cHbnwHjmGDhbb0MqmZ3u8mZr8OwF67H5ZcKNdE/udDAT/srMydb
sE5z0p6dQfOj0/PY3rlSMoQn8b8rEAXzUm2tCKBqDUjQW+YkdC3QhcnXX7wqUgDP
3y+rfbLrsgZcObO8k0QjmUi6FVkHo1QLHZPtd5wqXIEPLzz7rgCoMgxsbaVy5J51
WX7pIotdBAp8RBoX0eSE5JZluFmKTQGfu4cUGPJ949askgACppJdsS9WS2cFGczb
oclydt4VMdiOm4o6tnzDTz/nDw0/lSyf8s6ulhTlOht666Ei5b4f1ROsYgHdKKj4
VFMd1L6Q0ApUu99YFiRHqHzqWzH4RKiWBDUctz7tT2lDQ+TKVhv2N2HZVRRY+/mj
N0UDTSdpYhkUwlNwzYoVzRc4Oknp8cCZwaFFPkpvHcwG4Qom1njVI1beRwE4T/Xy
lAfi3Fyqqer+v+/ttvrcAZtqBkgplPcxt2yW7qalGlikP7enpTXBdcgDKUmp/plb
Rh2sMkN2MMWfGowrZ8P61SxtUjtoEybXaSoqwr05aiX6NeyKu1H38SuqTUfNnVo2
0DMU+5tRUk5esDHYDd/60Ju7QdWKGqHnmPS3oRBIlMC4I1DMNw69pddne766RAFp
+z7MGCfptYtypEKAKjZq17Nuruy9hZd9rDemB4ffq0NqFM1XAw3LzzMIlHIEvFHr
/+RmGPFOF90vagO/mQK7ZgtSTBJ9DmHhdKgXtTorIXA31SofljDZiTBvglFuQK8L
qy4GzVhwNcEelKoD95jL61gM+tAn84WHL9ydvs0vlWoGDeuyJwjogOHi8Lm+OcBq
eUXAkFkkFNcrHJH8BOKFI5vcPYxYbfdX+hT69BFfJiiHVv4knV2PrmUi1em03iku
UE6zAdaq5UXXp6DZnUyO2S2IFSAQP5JNajVr6hA9icNjGxLi7VdwePmzfMMmPbAZ
EBYpG3ypeHaEZkX68jkBpGuwlMC7xPOPdDlYZ3On4age4EPDSGqnodtPyuD2KCrp
sAC0BlbwsQo/JELg0+AAMgxJVCnPAtjJJ5A2/Kk7sgUTTuSZ9N7h5JF8v3xYynS4
2Vg3agqtjMt7RIzqoL3Nyltrc3BcUIHWtG5OnCUmBMva1V0yRoLHo5d2M27AkrH2
i2OmRitGH+EONopyMT5g6FGuvFHPZj4ArbnrGymvNYNHBul9vnmmZf+FUUEFrXOQ
kn6g9hlOZH0eJJliFSwcf5Qj+23Bu5AsxyU7FY6Z54GID/v/I41jAVCmU4vlKjk7
UPmv9NcQJoZrZL/ceLDm6IgFl0eq/H4BmQ73kwf3UBn6+Q+htt6B1yhkDyFGr+yd
kWPEx6raKUY521e5+S6t+Q3rdtwmG7sBfv04/ZS8Kz3T7jeqkhvyaOGJS9Pd6Um3
LYM+YDWKPJ8Ugy9t6W2y9ZQhEi7e/XTgUe7YKQFN6omTcFDz0/v/ZIxiN/2brHba
tlgl199J3bf1ud/S97mIdZGvvbpAm9E9xYcckweAfVwrUSOIjcpotzelTyTqFzWE
9UqDwkRpZ4LMp8N+mZhiahN1J1TcWXZM/09aEQeUVbGuhD/XmxvbSSFQcyN3KQkN
wPR6sv3EFnN6xm80whufm0TaOStGmzhE+zY3cNNLGQN1Bl7k91Xv6Kz11meRgq6/
OBuY5DVWPiJh+Mwc9tUzASb6i3V7E16e7Dy1NvLFPDJ4d7JjJiZcaRDrM85lKcAx
woEhqpXMGcO3viizI0FLoXzqQ7SShCMUUyC1TAhn34h2dF1ME+0kFXEck9jY8Mls
Azr6HkD/r2XYpTnZE1vOOYvyvxruSd3Q78kS4W01aEbs9bNINJusQxz2z3vsrI31
lHafzWfOJKjufwR7BakDX8SocZZrC13zJw5ty0y6NGr3ef/wXIwRYM3IHpnptKbq
hw1bkyABBcTQCnMMJJG2OIYriiTW1Jq3xJlQHBI3ffM0iHcNF3FCh6+A0w0SoxYm
zX2hSMRPlAbWDvNRnLwAQLaQFK8xFGW3wla+kAB0Mf0W9RqtZpeOLQxBbA1RJz7o
IQgkTvYyJ8olxGnPkfroRFd26fvTcSm+1D/46ZuO4tb9+cJQhoM2CWIYyVqeKmUt
93AYDYwHtUADzQ4QjQ6Gempy45rsUudDluqq30hXYvr8NqPtKrXni5lV3LuBZR52
Ke3axTEUyNXZucC9wz6gFesxIq/9X2WzhqVOKkS8l2zqqs74izPuUoghlcRngNCX
yVUQV18VE8iTuxmhLu21f9ESA3pTMHHT/hbCeiy+lrCtw41/c/Y/IGfUUuqKmb7s
USfOv3vW/7Ktxnhy0lNXzakUnSHIGJ2PqFlZ+byxiBOcwyuKA3QTMtSNfabASopA
My96/LuqkPi81hkQ/nmn0sZkqkzZaY0R030WtddQFclGC2EOnaAGhbZhgF7lIhAd
g6VdBEB6DM66I2U7g445b+x5qkZpeX9HI9eCCiAhD4mz8mL7eNQyNK3BwarZPwdn
vzbPF7SamSC4V8PYgukJ28cdSHzt9TpVuMh86BGMoGG4pCLx01p9hVf+ew6i3J3i
740odNkKD9HZozb6xitOoPYIF9bxu/h936jg5mshSUIV3LX6M+FQpz66XoRropnR
iT3sDvJkcQtar6tLiL1OPvVr1RK6USA+Ku7L6A4vIXVIJdlhBEs4fTftHbZJ3Ipj
Qzzg4Gk6xcP8f8JiNPx07FdXyx6ggyvI57nnY/UjrIpg6UKVqOsQ2HzWMQmmW/W8
X+SqfldF9SxZ1hfj9WFpZwn3wNlL05EO9NrBlcYvDqLvkprB7t9EGhzeMaJdSiej
3t149Y4iFA3RL/13WPB992NJ1rx7vtIgIcmnVRRXVGJp0RF7uuZEqZVaQp9kFLho
pxAtK3NGAa9KqYPGxfHPRhlW/q5z2is5o8YZQus69xXZArijNBR8vVNqTGGreyv7
e/lsPDTkr4SNmOvaaOI5PPmQ4FnDu7behUzbpvohJ4RhUL40cLHQ3jzAZRAb+dgu
/kXWxeDO8xoWgorC/ixKSGJC+8IzRoaGQCn6r+0cDafhaTa7XpIvwAyl1NPkJV1T
XhUFD+8sK4eRkR+ZiHbJWhcdpIA0DVeVpl6M8SLEUUE2Mm3eLeDUnY3nYIS7pDgl
0Wnk9ilX1j8GYRGee7H9zyITUvaoSp2xzDqOfLFhSMHmDLkqCAawmEGHHWZW+xSy
IDReTQ9cHQUk1VSA/PjFE24FPs1xrg7u/vXUG5afghcx54I0WoZe9Mv9822q32Zz
W11CkQvjYRt9cAAdiII55oxtWewGZI/P0CEZzwtdY+KZ5qwkTNh0TLYZYDha7l7E
wGmKzqZDvyonCJ3Q6SN2MATDs/KcoOl5/qZXjIKzwVKaxwag82ZyDXAMfOrFy7Gk
mWdzjtF8M/GVGQvTbsfNYa/u+15PS/Q/QPKfHTBruHbq7RrS2zsNxU2TIeBBmZ+O
aD4dgDZTAdGdDGXBuS0VoxfaE2JfJM++K3yinbTC++4M/2Gi2Rd3YCWVORQYF0FO
sM6azXD3jr9oNcm5RlXtn9OI8RrxCe9uUPgUtLmxR5oeZO3zvxrBazX5n9hr+oPB
aFZAr+fIAnwxm0wXJIy+CCLhAesoWRFpQdF5L38GJgKiNeAMbWmQbs9StuS9QHfG
9we2Qoi/UM48vxSTgSrQQs/Kc7bIVqQFo2GkX7uMiVbrS4uELrP843/j3elj97bY
2Ypb+7zaJ/YReFw1FxRRvwDYrQpqIv5DLf2yHkLEQ9R1EFC7rvt459nw5BQfKZcI
TfQTw4jRBd8lHH6SHEzpJ7m7QFtBi+D3wt+I76qp0Cedt/QhIZ3TsJcHQdq2cGsJ
tBeqNTHisGqDWdjs/5y0cjHN5J9WsKp6FLF+X94QcEHqNJooaZmsVx7pysulMjvj
C65YNwZcmkxV3zx3tc2ffu10jgf+XtPSTSn7szrVZVdfecB8WAMPe1wElp7j25i8
EjzaPGCz1ZHTxfSXzE+e/zCd2nvuKS13nVFK1/+aV8NpcgYPThXGpLDLkQzdLxzv
jy7a9kaV6OpFjBZ0jmpaYpRMaVk3hr9Lgz7oGTlKi/ZUGKVkQpv3O+ehjmLfeF2l
QsEul1hNwnP8ZSwG7DSIK9GNPJcIsyWSLQMje7QjtwCWvAFEwQLPEj1lK/mm1C8d
aYyi1Ib9AbqBUxPw0kbP8iy1DGNM1UkgK41mPso1zru5DRC+7HBgETVoHNOxbaxz
wT/MbVTVYVyD8OKnJlEVy94iddkiNpomrcVWn5ZifRlFPbYpX1Tz39DP7g5mnF8e
z0PdAc9XTT1ZZneFcwbBtvxC+5Bybns5QVsQ9pDmnrsnKHwV6GMwGWL1nDlNh7vB
ZFA3hzLQVb0iVaySV++PUPGofdL+BM9oO+ycHHO8Le+uONsdjXm671QuBLVkFMHc
ieXAGb7VMoTiv9CKtNnpZGvq+LZx+PJ0PrAWh1NrOftr27ktSZdXIuFdRwNjSw9w
AqjnYH/FifJxPD5IWE+Wapt+Ti9pVAYLCK0Da1vUXgj91SagG4n22fLCmofA/IMW
QjAsJSrIgTj3sMnpFFY8w3j4iLA0/vPbEdTNByjfwzvkxA2n59s6rY8a83h9uNe6
Uxhy7qHZm/vsD/Yd49BXOHhzAD0aMVpAlfAb5fIBQVDwTkro0+CKoh6Ta6uDJB9N
0R+kFhybxiATtxNyFofhpkC3T7S86daXxN3hs15192bMiNN5MZWCHmFWUe2VaFQj
fQYlYJUrpGQn/1gVSuJ6aVFgUX3Z+Z9QP/ZZGDXqIeDanoPpSZTtsU5AKh497sFG
r9jzrrDS58KV09TYU01YjNUr4WF7+kuNPP/0kzYDZQYsLRjZLouqxedjBN0yg7fG
0KNHph8YwUYkaYnrP7/fdvJUSRSuqJMSp1ll6IhI/qpIuHEkSaD4n8OgRrUldq5/
qJA5rYQCmUIRcXOI6gh9fZUQpkc1xtC5wyMQzcr78qBjtqFHiL92NBfBp9h2lxMn
FdIVNHGUx2OdkO27YX4PkqplqTdWOK0d27YtK1oK5NM1A4e+bawagTtP4hthKHmZ
TiZysrGupaZe3L8GpwJvcZCTPPB2FCp6H+oyOjngXolACf+AkB2OPUbApNWNASXW
eLBMYxufdIAuRumBpxyfuEAPy3tG7Z1Ivwj3izQaTkqvOgQnFPrkfMdeXNllKKcg
ahH4Mz+H7WTlmwgtqbw0V8+4TIQB+Sk4cDFi3LH3PwpQbLYhtSeVZLRJ7rH4FiPN
XxLRLer1IYfYQyI3hzBajpgkftK9piEAm8dN4noPbOb4VXYpwfbFhnKsrlFLHeg/
PxQx4wMn2Fm7Mx/XWfn355p80INWVvmm0kT2ZAP3dgIxT5f6He+jKuEXBdRZ3SLI
QvxxUdNv9t24/5sPZx0Gc4ZBlKFZS0Yf0BLxO7i/Im99hRwWfIwAnhuz1GI2pj8k
5uF2u7oJgpAgJCBo7PUWId7SysFzAcXzstDdHfWspgX+VyefBQGnwEvMtdQFlE5Q
fqPEBk2UVaP/v3tynUn0RUuEwYwijBfIzEu8rMZhaB+SNQjq/QT5hZPc2iTygHVm
057bWKb6a2PjyXrFK7iCTVQvdsqZmYbiBYtfIobeGbOpB74ULL77YeNuF1N8ifiP
1NCs0WKJL+S1IppEmNxc3c95mGg3FekwCpLBqFvVwssR+TnXZSzyYOwDEgOYwJeR
VuOaQosWAKYBcBH4SMjvyOkuZIZt/Q6vprsNF61kot53x9bxUvaXIbzg+ySIcLnD
v7MYFolPooDxlMgm2X+MJeE6WfahAZ/m7DUFCKzzT72aBGw0W6ICOGFcpVHtPoMA
8y+eZZqnQjqkT69zn8FbFhlhcttV2Oe5r/AHitYO0E9jncqhtmioKxUWZBqlAJxw
gIXxPyCUJNXxPEP7QvB8fsJ8nfjVmKOQSJOzofhH/YlQk9GXS/zyhaf6MMI1y12e
FkqF/jq1iZELdzK+w1/T54rf3OGMJeuJqVRn3zcC6OdO40E32Ii6ifR2QSia12Em
/B044MFJO0mPah4JDGLAGKGsowMPDTcfvzkUGiSoGRj2eIUX+Pp3Xu7/ocPPbvsQ
Nrgt4XlL7+JMW9Ifd4LNd0RiIvT0e2W1jhY5Jcy6M/A3t55U7Zzl/s9ZiFRihqz/
19JdfXkcFg+JmiZNlqBEPbYEkAvtpZQgL1Vg1HH6JTTWM41PgzHmIlpWf43RsS7e
ER019AJzfgDw4xPR5j3s4X5lLrk5yF8KpCh4gN3xlr+ab7UmJHMa4HSuSSjLXWLj
3BGSyw6/DwsGkhQUw+cznZp6cYZ3uGDWArmAVzGaCkQIwCg7QmcoGiWkKDqiJCka
uYl8d0zcuhy4TDvRnrbnWHZxN007Q9ZddlRUCe05R3Z0917ZDx9tsbz3V5JrqbVC
RfinMUVRoT9Xktn32l4iCYBGu1C5Z3hspHL6vGFtKU+hHRTCrRhZdnAFrHDCS1cn
dbYbLYyOJkeDs5zXIqAJGynr9eJRxp1W0VPGYgbjk2+zTyfDP9VeHIIxR4ngoqCB
PTWn6wAHWxcMrxC2x315cXeXKmGKTXDmLYL5cofoeTpBaJH8ftonwgiODXrMMnuG
+1g6rCc0VIfGiGj3N1aNXzE1z3nb/I8MpIB/Ocb624cpytHFqR/4DSjilGobsTQH
PMtuabhYNJ3kaihTftKcqWfJZkvJxT99JvWuIIpazkxLk0rtDrwGSJTKdfn8s6sP
gjVJKRpt9tT0DCLuJ184rjlnFrounUzEnCfHYsRxcr7tIULr7zIWoX7Pm/RrCqOi
Ahc2sC06tPjIz0RyWjaDcrfdAuBOViQfR769CQrDB2Q4sUnfiJT0Lq0Yr7MWhwjN
quZdCIA42VsptLCDqtmYdTs/776TUgMjIjoD/ybVugYipMtOAVEf12dDvdjMM94H
eu+UUWJencq3PSD6SN/EIe/bR4nnlMEW6VqMD0mJxxBLw1raGbumk7sazLQzSkCr
WEZRJQkH5y/pIYKmPSaPelV9U6n3k6Sw7p1Y4gDjDAZb87+b8uz4N8utgTK3K0xf
U0Pf5xbShzQC8qN/5jmpvDh3myApY0qwSecaXlQ+uTS6u6P/ix+34+WA5oX0YfMQ
ncWgWswVYhjCYLijIbucfLsHvg68X425OBYyGhGSY9KkcaIwV7Yo6U8BF6hJpaIi
dhe8jAQlryUREV/eAnCLksuhyxr0MdMqS1NQ+Qa8V8tvfBfz+3IhRFH71SX/okQ/
42BQvVjKjm2ospmC8KOmLkwBKJotaxshguIiDAb1BpSWOn6PaI83L8PjAIBSpgtK
8hcErQiGY67YtqVUbwAXV37pdSQAzrZR/9sQr0saFbXqrL57utDB144gdEfIn7TD
vD5gnUl7Mp6p65PVfiQsVgWF6MUlpGgMrBCPczY9J3BJzPyHVy4KtPpAzCyavxMa
el++xM6UJBG69Kg7JFFZV2Q9PQMHNR+XqyfSzsEalTq0tkm0LMpFb8XN3gw+h/QR
G0N+ephXsBx95oEZD90sYPr7pC0zlCNc8F/AvIzuI/lsDa7TG/h43wCJkpQ3N4iK
xm7VmocaU4Fz/YyhwY1oZCV57F+VVr3T15L3pUGjUWCAZS/yuBmOkGxDj5zaXPzA
cB9c0SZycKtSBRRaq0CQyTe7rnCLHUgimJC+Ekv5sOsambvMEd4URdBOz/T40gZN
OkZSQ/N3WXQKuKB18Mtzq3hM9rth6tUyrNn4uJtyV15eSAST7SV9eu5xl/Qr5XPm
+8fFSuSpLbNBcu3DtSxJkSmmiRhRzEOWb3NYwCpAYHU7o01r70RS9Y8NBVpHvAhq
5N/NDhKNBvb6Mrujqvnlbl7QcXVgAPxPhG42NoTYlEA79heLtqgj3dLivLVz4pNx
P2eJJfKg9y5R01f9S3E/knKDFr3jAUsUwsckkkDA7UVXYw26QIcsXvzMZmfG9SS8
pmT+6VxosNfv85krBM4FbnJ3rt7wVhJa63ChQZM4UErUNnfNBP2U1KD9ZK86UpH7
xeCXR3r9ba49ZJxkMiKiQBp1IY7cp9B5gVhZH/uBElcuVg47pebRMeqEgEyz7GPe
K3pGF34VrWWw6tdTknDa72uR915noAgM7D21NasdzxcIAnQ1p4yLxB+01y9b3DVy
UUTRVohJuLfiae47qYZGOgfLpdbXxeT3Ok1TPXIiR58zm4aYtNOeOSLjZPgzJ9KR
WEipNAbiWtOKOOGEMEJunItkBFOiXmRXQW6JIWObVH+Ti8ExCKMgVkrXVq4wz11k
+4cBGVM51Oo2Y98vzCjkX7VGHPD81x1FRxLjJOmUn4O35x3TdMUMwaNFyJrQOPxz
uk6ijnFcNAVEp2xd/fwYgIE/tOy6uYBbBBkqbNXIzISOnrERgfWWyT8VkfWLfzVW
Jx7b/xJWPmkWs4F2mTXhqP3yWkq0uz6lEMoSzlKJZy4Whiyo6pkJLw+fYsRM7wS6
GgvclNBD9cJ+fXPXuzr8uSRv8wP8ONR5naGt0IOhjk7Bp/zVTpW6U0rO8S3u7bpL
vgEuiQuiykBwtqY8rt4uu+4DlcCd+FhTxPB1h3Sjp1SZVgNOJwTz4FCKPVt2MoqP
yHuTGX8VCtOg5CVfzoZfYiPUFFKKhC+bYnZBA/p8d3tLk70jgh2kTIJoSo7rFT0E
SUoIovCFT8kZpFwVW2vJGZiydx56PqSvodXV5aqR71rrmD18jPiNmMG7B9dp4YJc
U/jivkKPM+K9DqB2xHZ0zFW5v1oKelH7GJRFNgrplTc87yxT1rRZ1Am6gDVYnG6j
bMZJZcomYLw/Dnsa/qOVFH9gj/UT4xI+leOW/GwACuryGvR0A9gLvw2zIt9p4Xm3
VJHEuGLH2hsaCxvU32vKnJxpzaBsGxX+QotX9RsYb8cXCbduv6whkNNU2fTAeDFj
IvQFenYCGxqJ+faWI4EVj+rpIFaFJ99LQdu3ZRkwU4aioepYj9CzxkukvkoaVHlX
3b3gMxOzC7W9F6uZ8zUVWS6JA5KAJi3iXKg5h4xbLxhjLzDP5UZ58F6ManDNKUb9
F7w2iTWTNxFmtOUVBZMdqQlU+FB/u0XabzIgmZO3iqBAA+bmEPw+jv57uRR/onks
fY6ZO6yYFMeJ99hgLi8gF1gE+TEb6dFmfmax4z8qe0hctcytzVggzwPGazXKJgoi
eB/eDS+wkIkoRIQcZDXWD72UGbcjtfhUtiPqNLD2yLrAJNtNio7iy4ZWpgjaS8nW
cvskGYYcbzjxK8IW9N13TTt4l4mhUYyDFcLwjdABs1VUVRVx3sWjQRnV+fPOjG55
eTDIdfzWz+ca9Y2StqoureFJOcPljw2IqMKh5Z0sB0tWYoJdg42Dt7jYjUZvIFPQ
YJWZpNmHFb37vKnkfVTeDOEmdlrgAjAnEdCNpgeb49F+bsiifodY9mn9buKLyD04
cli12NvIb92G1oHz4FKYKlUh8Gdl0Ix/n63/UCafuZPPXR1NKnVKRgu6DJzdcFqX
b119Invdihmh5RAV3hkxzcIvEdNusOshUgY5cXk6Vbrqq32XSeaRdiEJICpSyNaO
w35N5XLWqBQ1aXdvh80RXvHMZgqiKm/QqU6u8Pg1MfGojn8zkNmfSeQVwhqskeDm
ymfKIwKqfHDWTEskvvpzzyte99b8NDcDCmG4kcPE93HQwo+UdJ37OqVN5EDn9aZ8
rrtMtY8XRr2qXnHuUtIUtkVpvlbZvD0rFQsGcJ1vHN2VQw3Dwp8utfPI6i2FBFv4
udWFuPStt1TYKHB+tCMn/E3eTHXx4dnZ9LPv74RMavnhZ23Y6riqTje4glXbtnrT
HUjXAgdPSLc1yi/TsmXPWI7zIDP+oj5hXW7VrTudCGomjrLUBI/GsgfTN57xSzF0
O+i0aW0XyPB4l6BCxFauG2fe1oXH10/8bHib749TxMPkZoaA4UEAQtELTN3nTfMO
9Psr7i/nnx0J7qFuDMG6QMPeBQryUwdur937omt8tAvBBWmJAIxwGxQFQkpE2eYC
rsgsWFQaSTqOvQZF4K8NlSba7OCTh+LFACui4gr2sRmaTGZACQx9qpOmI3U4Wdy5
hpGwjRua9FLSyk++kAXjV+BIXalKwOXSg7Z6JdMNKPyP/60Kr2U4MDSSR+LtmkSi
HCc8H2H4mOsnGeRXV9gaqbaIeyU1MsNxN20daNczUyO9WuG90Ok71djQwhcq+E5N
rGB9ylCRZT+FaRmda6ZiXZBMxNvSWQFvufzA9/8SXqYqeY6YfAPnh5RAiBlk5uu1
FMGpcJyymlB+k0dNcZvXjEVRZp72eJfV79udCx81xYxjvIeb8Nz1n+w1yf/W7Gl8
kz6eV0pF8AKdhplR0yGUAbx+1WdUkowFDrFbCECtTZ5WN4vbrOWO+aMptbRNFrgf
X/4FarxnJHPUqZnknx+GSc6ys83WnKqo6qYiK2D6rDDQS7ZZIeiGxsYZBRIPU4po
t2CUf5foDrWaVPQLNfYOb+RLBO33pPWHby1YOPCLu4xvN2Y2T5rvl7cPwfOJ53xV
cCdfHQv1dcz/7orTRDS1N03EXZBe1KLDpjloOOodRCA3/x8mi7B5tRz7V0H8Ci46
NAwkNWQ0aVbqIFRSVhzZNxcLK0DPFwEkeupyeSKHo8VEbeDKyVDRD4DVkgkRuOTV
zhp4dXJCVhT2gNJz2J83VeraafzeylkmTyeuMjEVP9K8tQOXUE/cPQa/1ShLOhHP
Fu662uSGnADGXcyz2W2rYG76Wr1ze2Lgx9QzgpyAoK1MLHUdzMf2mH91cxtPdJiW
aqcPYxmHynyKmtCEIqkup4mn5gQAbhpbaqVJF+WuVBmIP2uz9T0THblN5+GUpQ5w
mnk3YcxUL+dr8kfFam2mVSa+PJVnb3ak2/J9/O8A6hFipC+OeE8UrenFGNvn5pPh
pja6R8X8SF6GQNYco1nhEgTOnjIMAjkCnwfxjkAZtK3a3mm7ElsngHGm5Q65w8u0
d5Tb6DCkKYil29CMiqvjOEhE7+ixY49v+I281HGO1cjv6v1Nbbec0uLcrsdzmyMQ
WZXWz/RFoG8IJi/z649GMZ++Pd6/wqjfCyVfUIJtAVRfRIDitigiAxe9nubql7nb
FEt9o6j5UVVMNFBBz9HIlP4lMFjFpmc/dKwLViL26Um8Rkq/d4SiFGA1Y0KIyBLD
8uuGBf/1FbKDooCE/YuX5gq7D4zNm8fbeBhUTa23SFNIMZw5GU2KdR+FnHZCgF/Q
Y3ciwDsHbzVfpt728frLGWsmOTcoN/tcCZF0OQZyTUUs2SvDbITIwg4s5Mhitdm9
DgpcWp0D38wxn8bFfTsP+NvsqkdAu6waJdkK/nKBAdbY8XBy1GiVCOM8rESRVk9Y
tf5hoGj+8LRWGWZCtU6GegkN0C/YibzEq3p8jnk+7kKDEx4Wkx6rO5UQaptMZGLx
12qnPRFTK+oASjaTGmU02BJbeAGj59dnMvhvcaKvespX0BfLCO9mWitFQQ3hOq61
QdC0cibGvpvdGyNft7Ip8rxqflVrb4/zhGDfif/U7TdTv9mUpm+ABKJEmirsct2K
vuyROvUJd207PTzIwI2pHMKjxpxrcnp2SMrGv6U8ZK1MAaUmf3vQVpPcrTHvoy2l
De0k19a+46Ty98D85XFPtAmFNuA5GlDRMu9o5XP9qt/hZP8Tls9MMFrBL2XTFi7H
Q1SFbz6BULbsGqZOqehywTa6F7brG3TjpHi1bKa8ZUR/p3eT5N5X8PCa30uh6Sx2
uJthhkNf36+a3XjrQHbAPLKBb/jKe6D/CniEkwwSwwQpxp/ln9sD1Rca71SgBnjg
dcgkFT+j34PLcSib23czT0tB9GxanMIRbHct8yVrNVlU5jNk8kXoF36DZeHQiQRX
lJjzqjwPjCSBmMG/9inpQ3mBnTAkrdYjE3vnJHjrv/tYC+D0Q9bDh/BCK9jqMF3Y
Tric/1TKmFdKgYpwudSjqi9uOp4PUxGX2hv9oEfhVInpi7M7Mn539c+VXTUyo3H6
dikyoHDgvbp0EIE+hOMa1CYVh02+vIsxTEFEaRvhcjXe1Ry1coviS5OW2kVGWa4D
qWDxnmSPOkPERExckpoqOu8HU4TlODA2qdz3lfg6HsJ9qBx58R8jSPIjTiHbze5b
vgy56ulxGa+BYsX/kdXv9HxQvu0hRiXgR7pSan9n2b/FLwLWVcZdrKbKShnOwv8O
1/68w9qyW5tkUKr/B3fnhkDfsTzPZdYY8YX1iPB//2z6XHys5bKzUz4a1v0Q76EY
aEEHFMFJ+U+UdmvgraX/B8d2NmOJkCGChTJ9BX1W8aJqz+XwlZJspVQCU/bcWgWF
mu3u2TA8LlUZeZV7jhPvPCnKzT0XnYmqExVXhxTgJ188FgwxD2br07pMgAy2doAO
/co1ZCNUxtwm3K12geyOgiiUpAU1V9BNSQ9vn7gSRrFZZt/7m/QPUDnNfYAvExxw
VInxvgqQbt1rM9vs7kLRJvqltSxtFQVdypKZ5Ii31ftOpxVvyzY1+OeMofWfS87f
IZVq3PM3Rw571/29d/E+t5b28s+pD8nWrNb1xu1yGev2LtjMuA5SvOQl3m2ZfMBT
aHZg9PDHvn5PbUicpekk/1h1lLsvoPYc1elhBST2gvaWDjlclRQSK7XO44xzOOYT
CFPVkF9LPGatFpBRBdiaUdg80+bJyV0VEnigSxNORijT7XBNjfksnDr9p3B+iSo/
on6aCkGew+o3Q8e9mghtZhmYy6lW88pmja2XtgOVRF9VBGBM8YaF4NFyKSUSLkWo
6LUZWfun1G+KAQSmzWNrv/HH0TXEqGIfDMBPBXP54LxNSwh+OnJZm2ArdF6rdMmM
JCKwwVGuG4IyTdFymN/ChoB7EgEQ7YknmiefSNVvUJPtNA0CRerN6o7w2mP9teil
fAE5MeE4W9/NZuHR8LQdVGXbH0Z3vlb2NCS5dAWt4MFfBuCsL7mEjxt8ZdRZzRO+
rcnMhBlsYkxQpVqULx3rO96B3eINEKeD2xHF5IqQDrHhQxD+LYnVZ7rADP0RXpwc
WCnYj0ocTYkGkPoEy8xoB2FaW7PbGV8qk3I8YfgyenMir7rGTgqraHGCr+rV1miD
xNVLNj4z+MsZSIk1BYmi0OsxtPNRk1HuIgkHIgQOuU10F/pzuSdBnipD8Qoc3WTx
rhP42j/AzEDGjRnCx6PuCd0VhN1CRmlQYboNy28ugYi4PiOTDLhaR/xzU+thtWBM
bCKwJzCz3+bCwMigjaqWSGS8mgNoe+3BnZM8l8QBx6pWe7d715y3rX3EZVwIG3/7
J3pCVFNUfZMyzMgfdE0Mzf2o5icVTb9bvn51XnfKKirQk2Ew+M/C5kOwPPjXICeo
rYComlvIHaksuaBE42hGObeXlyDK5uimFQe1coqkB/3LyHUpWjWpzuhKrF2NpRlU
98oCxmFpDuW2FN1JY+PK55S0FRPXsQGjZi/jSQySy5UVLPkdHGlRz1v5ff1iA6vG
+TZc3uIlebEgnWRodYiFezzGilI+99ZvjUyIMhSapGhxiZ31DP83GWUGgbHfxjU7
uSrGRtEBX7HF8AQt9+l0Feyd7GHV9NGRdJ9K2HvwcfmBw2K4MhqdjSwoIjK0mOxv
cqJ9Z2pWV6/m2vhr5wf0ddG/gt2ZipJnjqxnKgOoi5s2wlQ/b5G5CFb4udYP/Dvr
yqbOdGN5DgfzKWjxXaIYQLcfckg09A1ltPwpYSonWjQh5+Sz3MHfak2YwxnXo2K8
S1Q34btdRLLddEqvghqa9HQGS8jhXHX+jsMkSC3Z1KWMl2M9e/64RoVre+2gR9Ib
kD3xWDbrosdT9AKYo3jxfpeDUoMhqMsSzhGJgMcvcQ6sMapGh1m1XC2sUmluUT5u
iiLIsUtoVhVR9ZL4ArUDAoWZUCckT6xo91HgN/ZXtGQTsJ1Ln2PImuqbPPO8Jqza
c1CZ6pNtiQfCSRM7skFPE94uG7zw3inpUcrs12MRPzTZfNUqpBdjXGXSsqcisdE0
k4wkriaekeMRUdwQy4D2d3kc2LjmyM8RfiyBzol0qVOsvYgRqIMwwBLcI6m1JLxz
/Mt3vIlWiBt0W4coVo0MHz299vM7fgoSTS+3f4HAPetGrFbmv4nbRn11l0LgYD6f
HNfBU3E8de2Px9NHKi75JQLOD9QDuYF3RJxnO2IqDFYoWT5qQvWkcgl+WZEwlKMG
OFryNa+sk0Gt0G6NEJ3vi0M2nGJ4o0nKSUZ30kyD8SMgen9ELBEGrCPEHiva9WCr
1zGJ0YX5IeDsKxS2RjGU3TopovGS23u+a6SH26rxclxwSDzi0Z88D66Lq1x5ryOH
g4Z6muEAyEV2qQNJx/spySfmoeCsO2RYzXTe+x8Aoferin9A87MfUuOegfxqW2pM
lS3vUB0acMD4hHPjP1cetC2wY3Ouu9oEC+/MeUthnkoRU4rYeeDe0gfchC5omkrf
nB1V29QMZV2tS7kzCiK40+uXvZNTQlIuU1YAqRanUNFTEb8HlOSYaedbyMUjz1J6
DkJhUN3sgWD1UTT5ONBxE0OV2QN1Jmdj/mvUos7d5R1PSymtBZLpcSIZkZ7Z20kP
/BqkFh0c44cGpm/nqsZvUo+XyEshjhUrOJbi9jRBpj7BO89dGyShofKVR68L4EV4
eeqoPKa7qHVZVulWie1Tz8SNxfVfAi0LzeevXeIsvk9H9Ct/D/sqEESflmjBgGSD
akQOOYHwWe/+piBnsJcfx4A1C9Immyo7GdGSxiGcsORZ45DPZBwws6Zg2P37MV5h
3jlEtlQER6gJoch/6MYVLb6XwfU0GSRmbjhzYOARRQk2W3wURjPhe6SIXOH3ayfa
kaT5LMGUHREs6SpnEDP5zzfGsHCBw/0kiVTNcj+hGKec4k3RAsuijH4cKu0RSXkS
W5UQ9wV/irhJYwgkRY83TIZIXihVglOrOgLncMTaj2cCUKFfg0ui+n4nA7N3pgS7
+Kd8Kk1fby4YSoyMN5G8tPsVPbWxk/ZO5fd5NIeJVY5Rw970DaHyA7n7l9GyeYvz
BUhmogC079Ls3iCaOcIxm4eO727fw9879DkKQoEGufOpRcSVYzh2I2pi172PaA0v
Ynjo/PkBPD3hlpYasexJVRsv4r0T9IeiYn4BghMOWkZA8hQozk5IJ+xTzROeKtjv
Zj2AuS34HGET0jMRgVTS7M8G45MAiaHnoB4x92x1c3kmMimgHGjljo/1hxStM2zf
HQU0C7Alpstm2TkA2i/su0GapqoVYXSh2p/g1IcgS6a7GO9TFhcYRm8KuSFDYY+g
f2cyJ4N1Cz0+b22E5ZJLRzyyxIjaCiK1dvyDw1+AEGof++LAbDRE1NLtsyLJesEu
vWBA2T8Bigl8p5K3QZ3AEDF/S6mEwqsaagJAFkYKitXCtznw5dwCBWwV206yZTkr
2/kkNOIdBnF2Y/cWSxJtmLO2HNRUrdHrGgC6DgBaiTcRNszaytox5u7kkaj1xQeP
SJSHvHy4PttNqIL0N71M5SYL/WEJ6lcOQi+Sf5YZ3BYUH48hbs0WTMIWWWCQeviP
g1sM70zd+89wO6Ua+H9UEj6oWs7kOmbQ9ldZMtlrblIhGFX6nUuRxzJTvYG8jNoi
0b0NMTy6hcbF99YebxA7S/8WLFWTRNJi6O4nlHvMbkjA8ZstqOd03j2L0OxEuUqi
eAhIwlAGYEQDQRCUq2dYpSZtRcFeYQR42bvVHjwzjFXo4e5sPS9eCjew25GoS/lx
FJ6XFc3aEnCWSEs3ks3UpjTXSt/rHswOBBVU6xFwQAcckDqDZ5UJUj0J7v/toTKi
nw8zGMcfOuzcQ5YNVsDXE3f4JpqKngveRK/BmsTbJU489p58NY9vPCeCK2GWgMJD
C9+gFQ5WnsHYUCFB8QB8x11QSnHnvihEJ+QINH4vSC5brf7UTU8TcjNxlF+KiPRi
ttzzEw0S0B5Z3wkOWHGjarlCmA5bTFaZq49uYyet54CQBC2PrgFvbfMv28z9S9hn
FBcO8r7MTPqL5+b6L3hwepTnawOjJalkXATfYUYev9W9+bO4nWmiTWwCHwg9sCUr
T0RC3AzGYWIixgIidKNSK+mJcA2kJqtdo61ppzQfpUr7VCHkrAgh/UjKCCcrLZ5I
rWg4ZfhS4CNiv8kYbktqQrm5YC7zx2qKbbSvN8nNM/EqaGEFDYcNmDcxkMLYrNbw
1U7Mz7qYFXaqGhOrtQ2k8SP+KfH07tZuTxgAGtF4FyI+4/8b5VWd1dg9feDSSnlC
5omNNVBag2sHuXncqtXkR620ZH3LZd3xedCOo4LgzmD5Q1c5nCGHRDcWwMrwypR0
4lMLmyHxvC/Xd82Hp21qPKZmOzdktYGBKoIIrHPyVOzVc773FBoD8cna71Jk984V
FQBXJ4KBBJsP4wfsR9w79GgZryKOG00kubcS4iR42wQagr1/PEWVRk52HTkISlDW
ZPcgwWA6UVNBGFR8Y9pF9JR2p9mgTILboYst0SMM2MpX/5ElrMNaGv8uGzunp6TM
CxPVSXKNiak8f/quIazgenvJrdBBF6iwMuHTDqZq2ELf0f2KadxULiyTLTV6NGkr
Hshc4jt63dK+3RH1VbWiCy7GiHXY5pPVwLkTbzIuqWoRi+4ORWtOZMljuMKEgZGA
/RiiDTZWpPEefNchGLOrrcagzMKlz2AdjZRhqHutGMapuJgNNt8OyRjMUc9CpdOc
xzrRsz6RX2U+v0782eioykq0fB7C4FxXawWFKmCajLC1Zau4oRaWRNFkDmrD/i+n
SDBIdWWNAuJYiXn75IYdjIpuSDfpyJQKdx72fcDTC/mb/wGynIoXMKINVbiK/ovN
OUWgc3SLSuelTyg/UKJJVKkTNUCV0KnLE4AJ4SsFZTctghdjUl3dj7ND5i8nVmRu
pE1QCfoEpUarCMg6lOrPL7bOsxbsLEN168sz6gT7xXwcQObjiow1zwYtCit1B8zu
RWTpNBc3M7fKCmczn+REpVtZYqwD1alTNS99hedWWhqLsrPpBh/0uQX0oT4HvwsI
o+H9tgzWhNhzTIORhozMIejbnZrHI3hKIMEtdMuFP6Fm+9wfRvVtEvylXfSRKAZP
MIBh+sQYUL5df1JCKI0TbCvsoP+7feY+oxEZZkaXWnkz7Cr7W3dluYDonEq5UyU0
u3tZ56zkqJKb75FAISkyM9ZpzalxVToXhYF5dRGnbaPwSZUMoYIqkaaHE6Ilnazv
DgHn851AypdlStX9SNdFckNaM23p7asQm9eccczK9OY3KHbj5WMXZDIZ4SvrudAZ
albIL9JNFzRn6KdRtq2ZHuq+pArSTXO2BuC3Sq3cExQENre9TuV41/6FUWVJGHb2
y7el7kJCJp09KPkQym17uQJYb3IBwWTurb/NZ6bytnLmCbTCaT+YxgmG5BOqu482
NRwjRdD3O6Ma4c0F3DMGEeUSbSuC3m7dwtDovinPAMvgYLFco18hzdmvWccLmHrg
eJqJEluqMnq/mTAJvZDaOPISKTra7/cYkZircybaArcEWkNITbgX/WZOY4VL3UPv
OYKXL3mwWXJOR2vcMzKgrfoW1MGFpJp6WFx6ge8dUFBb/W87t480xpQUw9tBQVe9
NFW0DWfcJHDHyMi7lRIl6pC6nMMts4SUmicTgDrfMnUd7WoNBBgy4klRKYLlKOXl
kVE1OUWawPcNX+JL+HtXDZHetVauGXpWqgAlW31H2DrUOw4bQenm9NhDDCcLPK8T
OKPKVQSPpQ4UJ8GwktFqCpnxAHIwMqwxQtcUwL6hNBpPRxgCm+Kuqth04X4dzIXG
zukjSQ+FY34q5RQ59BMLJCToO+ze8Z5M2VIc2UVm1qzwoOF042P+5zNfXTBM0B6l
W0R8D8Jdgntg2ifA1b8VhZ2m5saxy09LUT59zy2BPcwPeBXM3EA5mb8c2AGECewa
V+bKMB3sFiojN1iJaz/i7zyoXXNBm6cC3FdnrpWwIiABvOvngr6ICgVoDPfQO0ki
P9X2oaCkg3jEjRd9tK8ZyVDx+WLC0A0lg8XQuCFsEf43wlf8LcEOPAXkg8DNKpZE
+ycG/ggvyMTw122uFcpwJNXlwf8i6Ukx8lqwNCZpzKQw4slkwyyK0rkjEAwUX3oN
t59c4a6qvWcO080NZPdj+EBxLv5zwu1uPugzYq7fwsaGWe0xiAB3/FpwmsXj2LWz
7KmE2O5t3PsJ1+wv3tyn3WC1dDO7FXxH6nQjJWhEQguDzR0TAjKNd6GHItaxZqQ5
YjgGqMMhqv0Ex5ztuR4aYYpo7WOb8v40N/Mp5IsgvNAOPeHgg6DIJzszERHVeb8n
jbHorx29JB22YQ9FypA2DPOljr7gRhvYw+S8kq/iVHtEiHmTlMuGS8qRnCWk93sv
B654WLVTHtHhyhc2UlRDl7lbAmfttUJjz0wvgYC6p4gh3Nk6AfGWjWeOwpfhHrJz
Z1jsr+oHXDEXEV3rMZHLPtrL2vE283krKSa3wp43wShLq8A+lQhDEi+qouq/aBdO
CJYjsTwKKb3N4oWPD/pnMNAX0XLq4efTNl5YNWhsDN6Dh1ME8DLASJ4DpXUhwrGe
1ofd2C5GFnjoUkIKT22TS06mb4lTFmsLKH2C4tvfGviez2VAkKO6n8pKGeQ8YQuh
XyA1keGtF1XBwqLIyK01FX3EJ46kEgIjluVrqv57+TK6nGMkt4sKlDo7vhV58+wp
XAvvjBdawybxjpZXsdcC3/M698kli0ugUw3Z+IpIuTC2q/9SolT4cl3GMzp4OFFJ
39R/eLeF5dP+dsZElaxABZclZJgc3RwZ/JUCmlIqi8mvlNlhKuG8KrWMdY9o17lc
MiqJqHDhlgZCBfxxSks3N6NXVARTiQAeKG5V8mk/av0ciXvm209qukK9H0+mfMo1
oqBpHV2wq/S9mfQ5wOpXTqNtbDVcOKyE+wsk6MU0mWXBMM6vH7DkXJkWNaBMpzZf
SX4sWYsnO2J8vOH/Of+3rFXNGxXkyTcBySzmEOHyF2smjskAen0/klCJuPdfrFj0
ENxUPncuCtlMEAeURQdRa9jZYxd9RhD29xEazVzlO/lKHYb0Fs+YHOLEWcD1EbtH
ml+wX3YiEH3ckDvWUNrK7CzmpOndkzwApc5yi/945Waxt//fXkGrmNHofiWojksd
oHnfJ+eXX7qVdQNtWd4KfNVMo0BStEdTKQ2UJHKOhEA050bQNkgWdYjKckpWJ4Vy
OlX0SWfzLp08KNzpCWSXc82Y8yRCZnrvud5FdRBXmfGhC8SxKpxP+/FMpE1qd8nL
PzATGGM3reyQjb+Vg+1FxWxuTvPhhcNlMvy6sxo0srAFc22vuTM/uz1QqcPry5vX
4QU7dF0JQo/aS4FZzdgaGGlCq7G9kKRmz1lGVXE0ZTTskpkEt6dFB/QWfk+Y7PHr
zxPd9kKC6VMRn35tRW0BeDQKobKSYidAzJcDWav/fziPwFYMEHdEP10PvExyyjOp
AJh4P4BoTniMeAKu7BYWsfZgcINj4N8niuznignKjiWmobASDB/7Sdpgg/d+Syar
3G/28kc6eIU37ARJfcz7xIe71Z5evC10WD87OzlGazIN13a1SYPgRd4CmImvTvyc
wjhSbVqFnf0odmtTMFf8OT18klrc6z3dYNPnU5ERwyBQiBb8romW7sWHB9EHhz4g
rjHtACNktONa4xIfg6SQLnfzVWN0KeW9QejiShpraewlHk8wL2eobJAw28DSGhRU
OzXq4osso81SGcVsBN8Tw8Jm30zmashMJEVgQAS0h+opFAtQ031+NdoOL8OfvC2F
erVq+X9CfuaSFy/71/e3ANJTPl0aq5bt3QF0TCbQQjaxRcLmDPn2DGHzWi4E9/Ds
hv6u8NfrSaoEoJjN+SRbZGoaCx7pA6DgC7D/9A2cizcWYjy26mogan3Lv0+M0RIQ
KZT2s6WITSQTi5a9m+KHxxUzuKKfEzWLnxBnKWAm+Up+yLu569lkaZWn6eASQfR7
kS4HmrF6L3X1qKAPyhjIy5poiIbRrtLQHkIyYQSJ2uG1PcVakJRU2GYlxdWDF/v7
RxVYOAnkEjmDx1h3YJrwxChgOfpwC85jggjq0ULtMU49G2OD0mw6BfQ8uoE5pC0X
KqFhj7guKelUiGVVEWqS9uMUcCafOht4apfEzSpNz/h4zufqefzpsKpl7Hu+7W4o
kz5Iofr3nuOeRwIQm9N4b1vynayFW/kUTwpxIMorSumvIDMGKm0x62B22FdB6mMz
MY0x+HzJTZAVL7eRiVAk+TGoScFj69rioS83UDv+xqLk6I6oFnPwC9lW9D2+pThV
9cp7blpCyewsT1hxSPTfa3fqUU8jJDAJhO/dgiehYQlHNuUCnmEoLmFPvqZTeKOl
yE1V6dcD/K+CUFKnyLNJFgyWLkpMvaMyEFTAQQkWz5AnyTPGVXcx6loPyHeCpvgt
L8B3o+FVVHhJkJPOQugLq+DUBpeXdsYM4nQ+4HWJGrpfGDcpjY/J07WZGdWAwAhg
vxT4/sLbuc/GiCm6Di1IfzSAHKomfScv/Fl0ih8zKNZcj/DeTRwcTAknBdUi4uar
eUMziCcCNi37fb5IRwJaeiEfnZaZQs7IxRw1ifDrfEYyqMEUocGzvd6gdUF3mDy+
FmlnJ529+eB6M1TLvDqujn8cAdZVTPana9HHuY1wEVwu3qGfQwdxV/O1azANIhLe
2Ky0PlLX4XB3MI36yQrtHDaqkIiJYesHKRVpuGOu5P+rfBSvvYRLRHki8K93296a
m8Q3BRRbSl0kKXQ2kNcaHpZPc1OvgugJSilqysu8PZVuGUJhp9y571nEmPeLa+gZ
Vp9xjGc0ANcByTCTX3DoCU4LtalJKt0Q5Sm3P0zUNf1TLFcYIot5BEIoxqbWuUdF
17d1nslS4at0S7dq0xPxbb83WFCegSuGC7IZ22Lz1viC0iBJB8+clcT12FjNp//s
jOH71AoIaqlNgCrrxoo0JNYqlnleXGUfio42LYTbIBBE6eBv8vTiVP8QvTdqH2wo
EUdcAx3CSJg5dVesometQc69h6Yb7Ldu2mjHxgmDqWM4Ry4yGH224jwg+5htbe1a
UKy2EwIfn+zYp1bp4XhA8biR1GFZyE3fq8KAGPEZIJMWoOi/TPtqR+1QUNhIY4DP
1qqDyk8NXNuQMCROShllQjq7QEt29h4SiZYjnQ0SWPLWFtKTnXjdvvCnF5IfcL4P
GOPCDS81pzwchmnN5N7EtVyIN4Vmj5nB31lAxYLmHsL0M3oDp8/OFkujLoTahjL3
U5ZgbEoMQvJwBt5XZbO4DiHZhMz7fO+l9ElLO7lUByoiWiusMivPwGLmRmMMztN7
rV3aZ94N1A72Ud+g/hLfrVlTBdPE4vgjol8SkzqCD2EpJJiIUQ9V7UynYIYcdh51
QjFcPOXglkSCXGk5zAbuu7CSczXvXZA3LH2URs+E6ekrTYOf82Squ0jWqvgfoENJ
MnQ1aq4F/1rv9j+FO3E96gsEqba/Gh6qoe8/ckMe126naowbrY1sPyU2Za0EEh+P
WVj8gGyQdu9NWaF0vOEl7cRSR2tCF4sdQAgLQKDof4IrBAgCKanoyF8JhkmRH//j
aKySTw8k1mVM4vJemBMli7guSyBIti4BW5yEyErefj3eTb6P24ynqzAZvmXbLjCW
TbHee6/zSRt+egOneRH0BdzwfDvSD2vS/PQMIhVdNcAFmfWNkysFUk3D+fCNsB3t
UJYd7sFq6CCw0JRT7L7L9nJRbk/mPyoOjG2ZoMHrzCha7hZHg5o/MV6aexSMQDk2
as1yOaXCPp2Fh9BdxVY/6Kizn7FxysQdsPIOnInX8zHNKuHUr+Gb7MeUpNg280iD
x7rS0qvlKWUfz6FTyIii0+OY/99oT0d0eom/f+YIXEpokU6ua1zXmxc+VyFRjf+d
ZtwaDpiv+X/uplJy1ZdwU4TEr0TCcP2s4Y5aBvUobz9ONSwVratr7+SldYbGCWOp
44bfhpCvA6DoGVlj10Zotbd2DqEb/CMZkXNr1HhIAnzZsSn1H+25USGP9PNw46/+
LaFh/Lf+cXwx/5+uNiMYZwrMECIoiguF0OFI822GgLYiHyDPk2XShPujXcfyA5RJ
lXekHkmPv/UJX92RurYWtVuX2Y2ovzpQG2vD+q1pmn+zmxnaHNnDLcIhTndjJO2l
vYIdgN3dHB2IRv/9pTrAGt8xNrWVITxeVvm0CCUmC4Ysblod9CiLLEYI9lodGAhP
F8rtOlGrFFYfc7U2lytkA37/hhDwto62rZ+VDVzxYpEfMrNUKPsOR+s9ZwNDUDaY
6OkEL2LIhdrZrRwWAydi317zB37zuwKutRRxCKXTi3sjTP40sScmMYLl32Nu1YmX
4ZTti/M5di3xO8D2A/cOQSoOqm0ytqp98gHXnH9/Ccr68XuRgiBcyiK7lGHgzgc0
CBtyEjXtUqzLdLtlptzE6Py51ieUzb++LFG6th7LZIdGIvV8j5JvDPhvmE1CqiTi
F0GB5LYS470rUvCPrGNs3N8U8XlDAnjLkMQha2zvCNM1Hih5o2i8XCT0ay62i8i8
G6ITg9NvSqpapqls0TG8JhbudhiR+DTK6jImNNe3Z/6noDc/M5nY48jVP7/3Mb6t
W9VI4yfWeJD2XDGigyo5VgBkLfmStyvmUFo3O9/47yUmUpXpir3oyFUU/p/EB+k/
u9vxbWQpNSI9RMDIlsH2Wreo0KZGpsRKUU43XiXgamcXTIifu+pHGJNWG+WKs9Kq
qwRAll7fFXV3spqRnZ/1NHz4SzBWphd/9S7welownn17yvRCWXtK3tg2vhKOFNQI
SA4Cg3ZmM9LYM53u69HuVaGZNoREyeSirmYcAKmZymULmjCz1S094r1piQtpHDrJ
ylH9cIDuTfjEmW1XRHKhOtshudm3fQG26o9eobkSIJ4z1oJevs0LUKESkVllY1/E
GuDXuTBvS0uY9Yx44UejjrjddBwELNe7W12CeVaurZoyA9kC89chJzTPxbrhIbJp
pHguJNW2ftsbNW5GuQNMkvqOIX0AlJkv6Gejzs2u5It3SZ4LlNx01chaQowOBcZ7
Uqk5Qv42CTi7Wx+qBpTzCJiINdPQw/NwT6JSKhPpYDPXPxvjylTOVvdZCcnbMHcW
MvIErlDEk/e04Cpio2lXmS1w29foIYz+37isVz3fm224BP0U4G4Y3+kqikitB+I/
lC1bF5r7tIqIDqpXVUX1IrgkeVRSAhv2BS2/0Erw/7m+Cc7bMNM3t4l+InfbLTDv
ycrii+V2oDFg+IDQodS9i7gLnjx70NxYPjUqRbyeu/VxE/OmQvidBu/6B+taZbKK
QtZvmalluJWUC5nuqgEul+HOs6behQ8TifgqxjMb9L1cFmJ5f5L95hXX2DcZ8JOe
8R9vFwt5CyeOJAl0FEGdc9raG3v46hY3wjogNBesI/GZMnOlh28Kx3aJUjhP9Q2p
NC+gnKOLrmKwyHCk5lE54upH/x4W5VXLt3XEbQy4gJKf70XvER/BMuOjbw87RDYK
5dX4Yi89W031E5HiCfLS2PJKauibpAfq3WzX04RYY0nWn9YhEg4/ButGbevDl0+8
/AYNR/QjlWcULpPKIIkIBtFTbzMGqs7K9t05qt0YeAqcyo0r1YUvSdEqSzqIm7sE
fJ304QRd3e28FVi5aqm31bI0h+i3wA7YaVv/ewB791w0vb+R/y0+dT8Pt7AxPx4Y
CJ7+2654k7TsMmhDU5+NARGf24bHdOH+PrXz7RvvfefRUysiYcmEIXUg9/RTId3T
dQpwJVPqd0vCHrShkcyr7Juecvz5RF2wrRMbvad/PXbYH/Xett1dUmRUgIjveYZ7
80FiH+HzwR/mKpUY/U/WmnNeab/ut8YYNx5jwaNzN7M2OVTQ//p9k7/38Wi4A/dD
m+xLf7n9ehcH/vnpUMN5Xk0KSMOwPfclz2IAGEXPLJ0l2jvf7Zrdtn8yGdTXt775
8mtt0c3ncOgAy8Ynhdh1eJ85PjGhezBmfLj1cK2LXYnWUOfJ/mk6kxR9OI31jOH/
plIhJCJfxdaSzWM7yQnDzxCDUCR8+fKSnXB5VpCHtOnvJ7P32EkLL3iu4nTzQLAK
VYnLJ6YkX6fNlcmgC+F+9C17uO5dPjRBD/n4pWEdR28BA52nZUyFsc+XaFdnovVO
LmktCnc/DfgUOlhfW1R2LySOTjvEZQ0AIRwqQAl14NyH4LuuH+Jvet/EJVoZgcwr
1OsrMpBZyPscrWQ8T3Ndq+eFM3ZxlEhoo7FAU0H0u+/lIPVOZm1JNZ6sXRVr0YaM
CUnbUJ29WS+TLpsd2gE69Q==
`pragma protect end_protected
