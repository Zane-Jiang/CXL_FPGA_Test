// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
AYiYaN4oPQKzHg42fkfweLNkBenzR1oRB7FGhUmtANgXD2oahAwDtbDS85ibfX0L
073OaaubwT0dCyb/4CTJrywPipJyQhfPQhvC8lsvrLdosqiJlDO0HITP1+iyI6nC
p3EOPHekyUgmLkDfRilG8UHJyR/642eSXTIdaGKZu/A=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10288 )
`pragma protect data_block
/aaGqseUijyPODdd7jzY8EqfPgGrzSTFvqZZUlIY7DnbDVxWgAjN+BY7sW1VZH8Z
MlEieawGGXuFuv+pBD6gNicm8QBalpCSPCEG/jY30S5Fa1oj+f7kLjKR9BubbgX4
rOmlZJCC0jkT9CNmeM2iF7DhpE3AmO4AQL4Znthtw/3/dSAtbH9FiwQnBfvDZVlz
VJNiupocDSVLeBoEpaZefcsdCu3/P9BDE+mUsuDQtOl7s1bRsSX3wmvr9slW69M2
Qp3JOLnGfyZqHGaiXGtOa/3RHCeJAvxz+EY83cRi56ekYot2eY5Bf33rtWp4hXx8
W9/zPZJNHAqT/kh5IZd9C4R4klXnDJHc30RrWFgqlwYLZY8YMEVusIobzYbhfGG5
vDPTl9lGRPYTEuoaFwdLTf7LfcSNsgLd609s9X4ITNxh/4oPoCxc9rpxhyQm09jP
ewZJOqri0WqNE2lXjJpbX58s8tMyJxaxOSEIllVv8IW9Bx7ZGa88WeXUBjxnWRfF
Eb0S4oe/4alvtgCCmY8oS0A4YRdlk52J4cO8QuB43AwImmAG9bw1r87IHRGECoU9
XG9wCa2kLYCbJinyP3lCG9EXo7kOlbWCzsVL5rhZlQbNMELDS0onH5Co1gmilzrz
5MBToNCvoUuPFSeR7lIN1c7G4r8CLARh6c2/5f+PpqM5a5b1cmKAuhWfZGKXmZ3X
qPaYqFAFUJQ7/o1m7au2uiYTpzGicx6mIrT9lh+1y9LsXEektW+6hxDtnE84wgzC
XxYnmY4GmonpPbCu687E+C2plozX8rqbpiuSQqwy54VlpUnzq+eDOoqLzUf3p22L
HLaHyrCkQaYRVDFZQLp4oXWSUvZAc2B+B13TzhqX8CRIT7DuxKuKrYroeKBhfoNH
fJB+Bo6Mlv5xEhz4fIYoRyfTtakaqvqtlwV4pt8GmJ60UGkOpN5XWCyQFdWOuZId
pvOEkKlmu0UoKfQqr+b+N+1piaxKNv52HdA289ETmW9KNl0rWLC3Y0tPTLVXLkd5
LBpydBrkgvNgTDSntFogbuTcl+1FpzL52s9F/CtYrtunD1jAaMudNJQ3DU33Ai/9
Kvp40YNK+xv9A5QMon6OmyZSGaxsvJcgJeZwRwIyFlOYlyxxipVLYCtiNi7J4sIK
S5OuEO+vRwYEru5kWvhaL+W/J9pPpJnkweEDLtQiQFcl9O1hkYYQiZyRWyLRw6BT
JW0PF8fgjJlagkDQMHpdNQmfrFL7AAz8oJLzwcRUW66f8/6qUyuy1wNUr728Hs0Y
M+NA+ipw68Azz65N9HigkcVmAVNrKv1F5jjoLCQd+NzE+a/tNEt3TQzpSskJ+D0A
PARS4Ju6XHhXMH1XFyc4fPijI+rLUbcf9hkDBc2p3dnBJ5391bu4RMlSgfruzroR
Ef/vx7jsJG0Ww1/kWQCwfoi2H8IBXAGS8uRLdxqc3FwZ/UjW2hROGJh21pHRGpNs
WkOYRmr3Sbf3oXxxbUxjDfdpSd2TRnwyJ0v8s63N6YQJYo1DWDQ+JnYGvwZT5OpH
3wKvOpoqYyeqN0Kb75vKB6S80dR4jz6cWpnrfcGf9KcqRqSrCo1AA/qjEP5q1Bsi
NJQBFnGPdbe0rZpDGyoajymSTUxwcsKr64Yq33CvGqn7ZXGgPwM9NIxOR0Ax56Up
SPbJQuhWYJ6aU7qjEgMZaSZXoQvlUzwEkowVGSHNBdz5V8NTgT+RiRaBIA1Xrt9Z
+tz7F2QtBEbu5K9kYe+5NF5n9erP18GTNaKLXYbXdvGnbg/rrBGP5UrORyeU/lJ7
8IRolSAuUVtr/Zt3jq4DJNoGb6QB3hC6cM0pZni3K9QS8uND8Cw1j1oCBABxXeZv
RJlv/4j2SsI9Imu6DCJ4uDecGzv2z3aC39CMOGGdfwk0K58OAzZow1weOGG6LV9e
o4BC1xF8+TKsG3fvLnu/50tdGUouIXN6cdjImoe952SymxaS5WdUO8cR8run/ja0
Zd/Q0qZc0lz7qHFeCL3IQioRpaMvXuUwHaomeGuZhIFnZoPzSbHEttPuBmJ5vYvD
YzyP/rxwpHfJajF876rL0aXIuH1GiVvL7gM9cafwYIE5W3t1x2b6ZST/S2SErk4i
IACQ4ijUZ5HNbydnPrVKHm72k0vqrchKCK6QYBRyYj7tAymT621b117tsvLHWq/4
zQPU7XR1wZ4Pk8E4JRoG+KnhBu8VrpW8nYKfjSUyIm/fGa7pOMBO1tyH/Ccl/PLV
2FP5kAj3WVZVDh4B9ajnQ4jJ4yqGpq1UW9X1QwKYS59dS3Qw5SE9aIB6EweoP80s
6G2LFmPonGkWE3+aZ1xkNvUZe5KHU6a+DLVegES++rMpWbXmRe4NX9Vscz6nFXT/
1mTYM4fOfJsDfc+AR8sNijgzEbd4Rg95gi3n0mgxEGjL9aKoAjrGY+Z1TJ5lV83M
ouXshW0ywAQpvaEf8nxRHhfsfGMHxbKUjHEEk3bUWIfX+MehKPlsaj/ryKg+1yf1
L7im2c7AFoee59fOvtwrEmsZlxKhkMPB12ST2vvu9D5rXsgDCFTzAker9aSyfPkp
5G88BxXCDmH4kjWipyeqVSWoZHQoU05ECYUFBPp0oBnmSpINP8ZY+3ClCZhc+HPD
XU9Tk0IFuNi8NnKfE1F6XeGoo/Lzf4vjrhY4uuh1yTrAz9/oPAQk7G+uz75hw1SO
RoOqZJFpjRLsA+5BVcDmpBwgc1EQ1xVj/2oCy8ahjLAN6J1XU6yxkR5/Q0sHwv/J
6Uq8JLRcT3IsaSKYyA3GWs4nEaX+L56G9AUoSxDAbnBn8KeBZIUTEfNQs9al8wSY
OtnvaFm4ds36Q2Vz0XDjB8J09yAg+hOn4FEuCpn9sj1bbuQ9FpYmGPAu72zVawcb
mWTOuYbDCHs8UvR9nReK8/za2Z+eyeFuAoM/4ySq0HO0Ur2qZeTftS74lWa+gaIS
GOlEPcbI6/yZYI8/dcw/3WhU4Nt7tRMq8gDy4MkG6LQP+ECLtn+wkIGzwgUOouic
7sS57LJZx/f9WjAWVK9NQKa83I9DDSxaAyYnhVDKTPti8s929WLEO0E+6JM4rMFC
dVqcXLbyLL2ut1kWkVCEKWa6gW6aE7kkscsZdSq+9/ojUpTTPSqGOmDwmrtYq0o0
+dygXg95i3Vleu/cc5gSnDuFVMHnZWREnv7ZMQEpv/m/ZecA8B6ZXFA50MraVYvE
4sm+RSv8q90SFVP+lxDAWCsrS2qHIHj8k7qk8Niix7WSmsX3TOdf57mF9BQ3v29b
C6o+jcS6qSAGfkXzh908EKEfswiViANJCNvEkkvfqcCLkPahH3FarnFWClSzawYK
R5abxthUJTZtYR6CKKuhcPgZXzcPoQo6S7uUJ0M4CkjMKIrf7SdVIJJrLdM+UbNS
ayAN/I8l45hhf9XVDvg1/NrXpXafbc7iyDapDn+P/cD3PHr3VaeFGu4YcHqJfGOT
5A9t1m0W3pg7iJK5tMFjFKvpNXLQJHnvLmCbBpcJ80DywkXKZbkI9BDnAoTiLktG
gzOsSiCg+Q82CBhO+MYtDJVytMEKYDs6AtJ2f32XIkEyakgidTZPSkShPWfgId9E
8vw3/GdbAmyeSjA2G1ukdrPXn6VP5SkxqcBt33V0SAGvd5d+zfq5rNKQBG4mcYRP
wa2SX374QUo/YSURcM/SVRlDEu7eNWH02HshFTX/ucYyUUcGl8dK40+Lrs+la5O6
Dh48F6BbSBnNMavyfUZyeTWW9X3VdTYCsv/YQnMCKq0fup6RlKP3/oPXZMD1Spzo
Hmi93N63ycVGoVW/NTA8fyIVW6OIGayRCz5r7LZ0pLI4WIZr9p/6QNBpiXzC6Lt/
zpEVM8IQyWAx6Hb3JD3ruXgSC/b67qgTAJG42U3nqTS6a0V91PnWe2MLVZCPmNZ9
ikv7H+GZFhbW1jxj9cXO5adWS3JzGnlUxjxNTUtDwdbkyA2ctkrrje8bvAfiUtn/
1Qch6565hVdVB0IIDAQ9o4GIO/j9H12QV4AT36r5egxB7yR7UGhhCFSKeawTGBhx
VKYm8n6c7jxC21E9acdM/keiVdgUr23sm9rh/orTyRctqEeGi3+UnYJvGRdWpWTy
Kq0qF8j4FZFda5DGyPMKaqyJJTQRYZqikSxy69fJ/SeCehTvW/eT0bOWsuZRt0Eh
YQLs1jenFZVPmskSTi+RM3Yn+MUQ2w8FYYkEz9AYhlMOCcgoE4y3oUMCWR4ibxDj
tWYkiWSWpbNXX/MMu1fUZFzfxnvL0NSN6kt6EIXTBnTCoG3MfyKRyREgEtL8BUBY
ic5Jchn0Tdh/FjeOz9Wo27qePAphtipgVbC8cs1cI40Rj8y3zsNAxa7Bg3DA31o5
wxmw4f1lcQlQl5e85XlFEM8dM8jiIhJ7u9PlcMr9B1hE4UIYz9xexPfzPqWM3TNL
UWv3obBNVuWjWLwVpdEbhaAeSwj4LEVnY/lgvYOlPRuC9X8joyLf2/bWlS/oLaj/
d3fcrr/+8NAuZtLXO74vbEgoik5TdH0QK9hDQoSumTlPc7fm5PiVlNwLmLG/FUyY
mw3KbvjQBHgI0CMTZ9yaKPP38XMEX2OZcsigoUxuVeFCll+qycITjfl+NV+11/xl
EWRLGUmAOJogyF8f7AYr4pQQMtJ9VSnuisLMeG4GohLrFmS+ZrKkrsS5slo7y7v6
xEwNsDOdS340O4gqpyLUYQrMiZPaWNCib3QpJVHq9ehU5ATssyelJizOyNwvUoFz
jM2Ncw1O9e+Oiy4YSId2eTOwsqGkkhkqitUbbah/fTR3Igqfg2JG9juQcuT+uEWI
Md+G91Emjf2dTXluTF3UyBjhqMY+bj5hyUv24CYPqF8aqePTeFhIwg6RwPiA3SmO
eP3rQ1tGEpnfnlFRlLZcEzoyLa1XFMSaOpxuO2FCj8pNdwJlF9rg0OV/1YswQP/C
/XiwCeJhXfLh+5RrYXxCWxp5csCTwIBf02HDz3M1xO/fEGAtIY8lYH78SIuOuucW
dZGneQlVu03wXb6HRL/r0zX4gV+t3n1n2OJ2tfWXV6LdosaPE55a+nps8qaVFT37
SXVbAYOcCvhWVUBLwp8hEscT78Vo0u/ri6ilC3WwxQFlYzF2KDWZx+Aq2JoBqkjz
/Zxi31MHu1TGFKrmTimccUy0s5V+z6w5h5kHJHLA7nLxg95Z2TkEQk8FV04wKnFk
vzclOTxNw27b3rf2PSJx1TTcmxP3WSveOmTffM1YVV1qq4eWXZfd8aDR98Qcc3/q
zJb4HrwUSmWERfTsoBNWZlnz0mxb18sn4wVml/K1OfCTh6wJJb1WaqzIXfwec38C
5JOaqoY8vDyXybQ1vBawEDZpokSUrxVmyTK1+5tQM1mZD6gVxhogEGH6ZV8b2YXP
ReHdzR25bq7vJwx4g2ZwslfiNdw+dzjLLR9WFTZ0bPqBNnFJXJnwykVkrZ4izcNO
wRdlzcEqFmwYVr1N/bZb4uQNMsja99W+FhFSyezGz6roYhBohApZTh7MjLlQ1aMJ
K0sVQ/waskQoj9GqYgHmL3UuU/nD0UJcZokoDyldKWQThlY+tCyYZXKSSlXrtHMp
QeVmXF9pgpEzfzXrufE8FBsK/N3rqE4VDoTHNpidWRq0mZ2301JQXoK/UhBrpsa5
OTffyr/F77ny5R/8nI1AFyI2YhbdRQEpl+l57uEQptbjr7QUUi2H0NgWtKrlwEcW
OTbBFu8C8qeKmTj7JGZuNkd4+eSBidWW7h/JejGtrkNzYi6w9uqfn2U/A+Olvl0q
BcAoeWJK5h4DtvZHpNXqSf5on8N+DbtL/p7jM9oTiz45wVtqKSEj+35QyfAuY3NR
+Vg+3/YQrDVz8shzoiOnuaF3hUdGUWHt/xiBJt3Y//3NTL/9Q/XMzp/F8yAkvHcT
F2G+rtXoO60bW1PDJ3QIX914vUNl+iYtRkdGRENrKl5iNxstYVfWJb9sypIPS3IO
6eaUGeJVyS2fAxVa8/RC1zNpqxFdNjkv+SMvydBwoa8v4B4zgpqaP6BnYRnIMSSZ
Ge4T5xIEWFDoXA9gStJ/Q+Nhk7iZRflzOFKToZ5TzTwAnHwmfRPGcovrR198WWcs
8hPn+o53Fa1B/PAtyvBpAyYD/X5XmenMQLC5W2LjO4i9SyXio6ZltCbua2MmouLf
L4kOS2or/dJg8Vewcz/iDQDva+oLFdeTQfXJx05nlmc7lzhJDokKqvMvEYAvZuDB
ipwrXr3wprfAPqq7VHlz8xQYOGb7vgRO57QQ4WMchLxGUiwdU9A7uE/8JHUoYRh2
IgAnHw2SXUARUaMLHiglPU0EGLGtupX1/wjXviZ8s8Wi2a+SKyeA4T45uy4KOpGb
2cMSSgorwOJdW/BNas4lFDbDvmY6di0dlWAoc6IA+52Tp21c/9CDIYuZvtQNrj/J
vYQ4ph8G2T19ESFdR3ccIud/ETwO0ZiloA0bwKFHbCJIx+J8JDPhYoOdSXGMust3
BKBi701USRAOT6BxANypGdK2O0sHvbdWV3GXlc5m6cwBjTPtYE+0gA1FzWE4Pqe/
q/x/wn3iczhs3FzijEVIAU/icSSVmKLYhWN39TbbHovH+idnEdSef/mRsZpiCJwI
1Q1yl51PiLziDGAQmsi1XrUabX08RcaESau10Al9vpIzEqOXlrrhrII6wjpYvNh5
PRLzypb50EIdieh3j4wL2Xipz3aQYUQyngJe2SjuDI8iD/1JTzNt3hNwlTuW5zU0
lYVoUBnGmXFr2gZRMrXo87I4GvqjywM90If7lTpox4d8mlLqHV/cOsi+WoocvmvM
8djgB+GjKjmoT+z4jFnB5iIO0zXZ4fZB6MtVsBIpUItSZkoOMop8fTQJ3dnB6k67
zGxuNxbUNrjvbukZfIz/zMoXgf46Ia6wgHpuq2W+NNiweupP2h1Q2RThXWAlrxEw
+gmb4mzwJNl0f8bvUVniOCSF/bWSR/M3nTxuO05AMGorbWubVegFFBXooZOYOD3k
tlg1za+Vh4OaEqy3GHrOn9f3uthw4dDidi9+3qVzkhKuuyrSy43ftOX1P0JVgCDd
X2g34Kfe9WkEbWrULDTyCRqML0/tWO9KaTx1y+hHf/Ai4lHDkbRfWKQP02mj9HZ5
PTDUignTAN/oeNDIsTKjijZBkWOvyRCS41PWltvTalL2BuO+NWlce4r/379gw8qf
5m8DFbPlEIUfbDFSgA22sdvu1K7sKc/oMer8DjZIzktAZYCfakNoo3IyWDjR8dZw
GF+mATVXRBTsB2SnrXxIoZHlz1a3+kMpcodezYk1wSC5cZg4z8FlrjGbF+tazu5e
9XHqcs3evAs1oTl8ewliZqHtNyki71gZ1LN2yLnD4OCob/7hOiJRrc3O53aGo+LZ
mUvb2zl+4+rhhR7EQUvLKHLrm6hvB5snP65+mMef7q1mjrx8a21WPvAlzNv4rJCu
7onAjGwdXISvFDe6DlUTmzzBIh74de54BYHyqThO6TvTDZXRWcltxeHfqZgxJZD3
XLPExhs32p/9P7kgoubzKjLULiVue3TTjAVPEsiPTUfZGvSMKreq9O4OOkd9z0Ui
+B3LvWTxBzCYtjm/sICIPd0wls2x5QKDRvsCqm9DlGL7n+ExpwS9fDkQOocYoWtz
15thqdvYmyjP0H9z3NEGfTsyydjSqHw9+OppBOOa7/D2KHj+oMH8ZJsnIL1uFV44
BCWsmHwFUAtksEsKRZEBOfNTPGMJyursWmBqdkcdKWtCaRBF2sxnPnpdNKn+hlL5
H2dukxr6Ae0t+SGETZNVEu0hL0yhXKjmKOPRAZNm7uP6chpkSfcYSq50mkRvhKwL
ZmJTo9avYola9dWrOAKhMo2/HXLlZnhMkNXzK6kxVMW6ZBMiw91asRfpM0WM8GI/
61dvz7PAPO7NhT0ZcjlB04fmQkmR+6deJELymAv4upaeLaFb1DY8qvlx2FxGhjR5
x65+OhDJyZnl9HNWWQYXXBBQWgCDtU9EAhUgT2lyggkIjGExcDXtp45tyZXdFLGk
hV+uXIUizfQtyYQyrM7ar5fCG2SO5fhXn5yz6MerqhP14LXpb59FyZ6ffUXTUCr2
sazbKmthGebde14R17uTmrjszkWaSKfr3tiWdrzjmrWuINAxnUpWUpKGzLTVSWTd
sbNkFEBBco+L26osw78SFFGTd4Q5k/R3qKIcEplP7zRhmKRDuWAsnRTGtcIPi71o
KUy4ie7ruCGUuRMk0Lpj01ZPnRmFDnEI/mGqalS49oPzoknCIioROn1b3F5G7Mgl
xuJJ1Y6y49T88WZP44K2wJPMpV8aALgRvX/Hj8GmTnHME6++A5e/WcNrNDfHsDce
nq5yNdJ5Dj+k9dzTzzViVnggHwAXjqDxx8BJ3zv8SsxuNuPWqOgWoaJS9s2+EL/+
o1LIVRnEzzfc9prCHBDcmoLEZ6Tdk23c9jmN7DRGyxWRwfnD6Li8Ex9XFtZg/QPp
blGehD8UgmYOxPnUVV4Kx+lA5HgHczkigh9HAMVViVNKmO7hDCXUMGS2weDsk6BE
xE6eR59gSJrJVwgp5EcvxT8Rz2wn48Moy2RHl0GD718u2KEIjc4S1lHWRy7KeThm
TUxoKxr/ygc+LkU5+WyJOkdsqA2lFqdHecR8NEzhlpdwvS2pynvURhKZDlDw5lLx
/JRWd06z1lzXsmmHDGYpueNzwG9P+D40sXnFMiCElKarhRQJ5xE9dgb7JaI3uyXi
/e8L+f4KnCuL/HzNuZXiXHOCl4krssHT5vJPSf5KCcsU37jO0d9Kf2AwdObJbCkU
sweqodymYRbXwTx8AbADAicHXDvMKBlaL+ftIkI2o5zXEoyLgk/VfSRVfFarvSBz
L4DV8o9PnJPdXAGhS7HAK/pGcaly1aak0mwoBUu2bnCiXMrNHeOSov/AHpEksF8w
Dm1Pumbmpt14AXqHRdG7b0JYRqwAlE0FDvOyLTz+msLkTvOszB0FLQX+OhbJCT2D
oOQROdsScMe+QKDTUP8trKb2YYhLmultEYHUKFprLA5RNVqvT2kciqhnL+U13oTC
8vWRck9+aHIxnXYkkOjRPd4aLfkZUoTDgiwQ3H14d3P3fowDCMSH1xZgIuhAl3Ue
fBcRgU3OEQyPQu3v/ix1So/a+FrNA+5YW7g8PPXf2o35NtvHCjdtEnJ4A2SvnJia
O2G7DtyMovpmrItJAk8NPYJeMy13R4ubr0G2p7286o+YtMz07T5JQFGLPc9vRP6K
xSMEczfF9UHpoufI2c8RuPxHJ7IuVTJtyo5hXhXOD6Vn4sf8L/Xe3mtGAKfNkvWy
bIPSZEHyzr09l7M3/Z6cgT683a0BhAIW4hjNgjoY/q56kIrOS55XJX5SB7XzLt+0
D+vJt+qYydz/iINRtobvEHbdN3okPOHh6gK0islNJr92WnofB4qxNmFaeb1/vICJ
D6oKoYt+2SqC1eo5Yfg8UbO/jpaPX7MRYgY01VU0qCoOhoRFYasrRcERP38yV2+k
wJRL2k3SsDdtt3EgxwojcDsjQrRb6gJti9FYUL7IlelbkZWM2SIFBoHV2xv7htUl
4gHu1XonCrIaIxqfAJdbSku59KO/ytlz1fqfg0PzU6kHCbvNp4pIcqZWAMGizVsc
/0VwNL/GVDUP3BS28oKhnxGJCP3DtBf8wMsUe7hjwhkYZ8FEu17c1lHIIxUivv+n
G1AiNBQ4x0EEcc+RxLxraUEZRLnSAkX+6lzEWbnO2zSdTSzdnnYThdObVisycgZC
WSPPmdB4xc6JDywQBYCKVBPF6/zEor/gHFvKzTiUJhIoQgTCUsBPwgVhxc4Z5D/X
9C705NZI1tEqZa+UCao5RyNESKLmfDe5MxHwqzJS+9hBaV+o8G2lYKnVfEcR9UNG
TNkAxdwEamCQthAK6lffoossjPCigJu54aeuGoQp3BzTIDe/kz2v8awVOm0SMDAs
BNKN6oCzDQVbvnKjd118hQi/GtfkpJ1JvZTpBQ9Gd4dVtMuqJijx7csCzFb0lyip
te2HOQIPtnc+eKNZjpmIRX6SNqBG/nOXHUVY1piMLzh2pNa1W3/6/IsM0rCdeMe0
cqq9PIoIUW3yyEos9SRqmCFPuRr4RbZSTtO+vFNic2q17TKDiOjNEGusdCoQoVi7
boXTz/9jfWFpoRC+Toc2nmoWNZWa5M0Jt4c+SNc15YqDVyhWAQ03A/jMx7xL8c8u
GhChQh3r9ZZF4vfYKkjA2XK3LfHbZJABp0LEEJb+rgMUTRQmvRARCrMwTabpyJ/Y
BZ8xoU9ie1AbGJWUC9qRB9T5Kg2pab5R1102h5P4UpSpvjTPo+DVihzy1+0ntz0l
d+tNtC0ukq08Dz+sqg0BZfUCjFnPY3su5V03OWAc0WsGRpwqWbFIqqIlCmempf7O
VyIu6kLfjYJOq/iIz+GgJ9mUzYq6ZCmNusMgsZUjMIEZCdI9UslRgpGOGvEWIOT7
gCts9LCr2xaGE7eqRto9WHKC7yjuqh3nSAwbYRJQ671+a8bP0jwpBBLoMx8G0xXv
DUyfTYPELuPrZ3BycUbWz+KP8MzUN8gqfx19YKY0DKAGTMwkAHtTU0C0k0NKL6C3
MGgHcAq1evpk7ekZBQ9LiiLdg9I4g/jwZggGNLYJHQOg0ANC2zCNFUePlccHjn9L
1+auGi5SZTDep53h3AZ7yy1G6UlwT/Y/kH2gZ29FybGG3mYI3OGO+YuAmTnqJdHi
8Qmz6usDIeJcMQf/wAS5Apq7iT57LOAkIsSZZaaJGWF5Fn/a3J2xXpdgXAJkI6Mh
exfmPb3fSoQQIobkVhnb8/6svbHKd1m07D1E9+UjKyfzr9G10MBzWnVOEg4GiJQx
OnSQJ0pkuT41Ba/gCY34H61AmJ7hA08wc6lWuLlGAoNAGfjItjOTzWRzaXL37W56
SrbRv/aZxEi15Ne+8XHy/IJUoTl9Sb/uvG6mLq3umCrVXnDfEkz0/wi3h7OuXXt9
uwsksD9MnS5Hfrj8B7v7P2PsAD/fQsnHNup6gNGliGY2Lsw1qdPCuNPrgYoUfKfq
24mhBY2U8BBAWf4XuKktkVbSY9TLkVjvHi82YSRe61oKWGTQ5Z8Z1qsrImDlo2dn
QhLhPLX/5oiNTWQcua9qYSp08GL725FXCtN7yzJiL++O5Oc/LSWacgtZ3kIzGMeP
1DIYy5rlxk3oK3qRMUEqqS7cggdoGvz2SYk3WWKUIIXbJqMpKGm1GQHrYqjEZtqC
IWCmbyEdCAGdKgbqktaZ2x/ay6abQVBBcizJJ8z7JRK5YEAi84YxGmmlLKlGnJ8I
xcxTZQxxNNZ7OQ4H1w16qgUd8EZUr7fDzHmVb75AqgkC8hZf5EIUHc6g60I1TWkC
5y05ZSvaM01qqM2Z6iuy4XgBzGS6yF3aZIVd09IZq8A2KL5oGA/tcLqPPY2VOUP/
rpMboe3QHQ6L98kjuvVUz0WlUhZ5TTHZJ9jT+2c8+InX9VQ0uXz1Cpx+QvuRukFy
4XmAld+8xQWrRvP0A8uHopawZ9mRZy1uUBvWKBpwaFJzaqh41OARkcY++0FBsZ+Z
WP9LtZ1/PXwyVnQWxtZhORgeCZ7gCbHiUvF/nUw9e1VHySG9LE6rW4fAxkAlEIi8
THpdUXRrewN5wrRa6XnB8do/oOUM7x1/N9zZFHd9p/spNG5PmpxvzF9QjkrKJb5C
2JOjJupUArPsV2cUMiDXSsMbjT1eGBVhYxXznpDmIoYchmSbbmla1NGKfiJZgcVa
G3CmmErz0SrXoG4hOVXJIlarHuUBHKh4yUcpOSRo07/8ZjCb3TZEASbpzPAuSZ+I
pdlbhBw8k5hJGbieVi5eJ/CbxDDWfnvnINxAP04mpiaf8SFntmr9uaBMja660ZNB
hdiGVOQlJOwEkMtm6jPxO6XkdvfsxKryygnRY64O8QG7D6RSHC7hEsBMwuTjqc71
M3NhDc97+mbroCTeG8mIFKNnlGF0AFhawnIWJuqP5Be+VQXsjpkeVUGYZnc4gOmO
2tVqaAjx63Shlr51gxztvXqvZhlNd9OaNaeujOerFM+hFUB4/fOkuZa4DmrUhZQk
M44ybIzR6KEackDlyoxvaE6fpDSMGcQQbfT+8ESVZWzxboA5kiMvyi3P6uFGjhB0
/p3J4QTs11XG5U4crkf0+kNijGjWOjAaorhj4X6oQkoirV3g0VC1uEhfyuUF7seF
ZJ3PQvfQylcIohWgZK64XkBDfKRcsc3pQc1KARNFj/fHau+7dWrfXN3M67qGtj1c
4uYQFnj8frOVdxnGFXRWE5VM9x7EgUNDT4soRivJZqatNTwVU6J5+rAK1dRDWeXh
3Lh1AN9D6rdrENWahPftFZnq0zYarNpOrsXm3oyzhFUKM0eTyoYhR8d33qCBS7iN
9Ld/3UL/RvrqxECMhLvVGdj49w1LbuPGoQ6vV0oOiyhjSveTEZcR/YstOBgPES8K
8UJB68Azpze5UCL0XWtnfMZ65SjQRlb35KPus+7fKqSNI2POCXxdc0my2uI0DdPb
VBpmVBc0y2JHZ05IPdMlkpIvK9RirQZfC0x5kHEj80eMlcKiEE6JEHTIDhBIDhDC
zHmkTlQsq0CD3mBPAFy5fGBrPyoZIw310yH5D4j0MbK9MeAGmHluaPdmjnOw63Iz
n8mMVlUUX2eHFdp1rTJD37mFfGKpzHuzIgZLQB12SHlbkekmaSci7XM+r1BrqlPt
94sb8dT/J5AW9usHChXPeOfgqbgnBW1GmiQ2NzRrwn+yWRfv8a0+ZtOuVEnm2IzI
sNiWm9p/XLST83SjwUbKEMzXUzuKikrdsbHoc2RFoOqxoCTikJBBLYzhJohAMldP
68ALlbq/PthX0FQKpiAF7K4KBerVP/T8wXf6ickgI7j42GmTbGcc9DrQQJ2oAvD3
Y/il/OZonl09vvQKcfIezfsJIIXothnexPa1agbS/foFO0klkQwOMSe7mAZyExB8
SDGNdP1FkZi8A7q6LUaptaMSCxEyv6h1tOFTTozRoMeoTOqrBjOk/wcetyFup7JR
o28dML6+fRj1dqMhjvsEIf8mW5MdxuYWvA6tQRyfKRnben3GqjJWTDs1MknzIiQ6
60Hd6HiPxaI6h5C+ucgersVuhhifh2Kvm2PJwz1PoYqEnEuJVze9uorthQSmUD10
hb9CnNJgYzszfjxPOOeRhuDDbtVKzk8+aUWn8U+10E4YWU77soLXmDxSDcVNRpLB
M+6vFaBH9n9/xBYm510LF8TN91b8Sh7Y8yD3zdU9tLA01NTQx2kPxYLfP1jNze8a
c83qw9j9fnWg37PREn2omLEnxcWpi1alaSNaGYAg+Ij/55vBL09ulQEV9lSmNcue
ejCep4wuykcLiJzFugelpC/0dUIO4zg4CAqKjI6MeQ3QeeNwAUhDpL/xskD0h+FP
lCRLq9mSvD2WpUWc1K2YsEPGGkuURLXtXf8LnxN3GMt3s5FbF9ILSZNDtVpWbSyT
nbN0bhaO3ieZvmbd3eYdTXST1e+5MR0KE3kfL4YHzKB5VwT81omVEofjp1fETYHA
2hPdml8F2xG3e1nkzO8i9Vi5xGlJvAqxE7W8VB8f9aE3EkS3VwT/QZB2CaX2D27t
PFYJXNAS1vvY69A9tjWXn5Wd4WEcDB3Iq1kU3wsaXp9sFaLppZ/tMYqPBJnvzeWo
4UfUzKUG81NMCGvba8RaGQdiZuDCGlDDqiuw7mR9rPIj/wOldKyH+V8CZaeTB2FG
gSdZqr4oKTPRQ3+JZcsa5w==

`pragma protect end_protected
