// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
PduKI6l2t/8qmRDZfWOLTVhZBJ9hahwMQyHYAdMzx/iisjt8hKhgcZf0xFmHkPHk
SE3jEhL5VU2VPtX1V8IJRuCASOa01snibeqS7jaLE9EOju8y5Np2OU4h1X57Y4gC
vJqoaHma0ear2aIGR3P+t5raxTU6epf9IZx7nI0JrQc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
gFqLB6wajJqiWfp3851un38z68vLyUpvrYNBG8Dem7AfWdlC+2m+b0yE+1KiSY/a
5j4OGT8vlC6O2580dEn5hMxCNlXZu/HpRsAIQKXJHJFOI6ooTrtGs39/oqE2uV9E
PcEHtT/EkBPXZy1QLAB8RY87fpOybP5xUaNXiVIRI9rTOC4rMpRVixL7hY4j2W+W
GfGXAJmxpJuAujLd3MUgKYSnwRtlT80jhNYtl3w9SGs5rWQi1jp5jh/0mNQdafMR
X1Gan+ApASI8RqomyyDRZ1uVmejhRrlhm3fWfUoQoSNvLY7JlAhhBtzCYjOhEOQr
L8EaRb/x5LQIlzJ3KHD40POP11qz8r0Rk0Gnog9t1FYhVcHgXHRCOfNMYJ/Ru5XE
/4LE1TVg1sKqWKABJ7gEkXHYkVEbVcelM2SgJyNwuXfD6Iu7NwioyPasEL9Jx03j
E6eT3mbqusQ5W7/7SHDlpE6THtWbH1VQ56XWc+Q++AkxBZ8nIh/2dYD2vel1Ww8d
NF1VDtPOFtc2baFM1QbUlLU1peZPRM2oCh60T6VWnQuD/nkSkgQtajLD9Xa5UmHU
Grp57q8b0L1eR7ZqdLIfqZzYugMsDh7Ft5ioC7hSF2aU+GcPvJ0maSxykbnEhtJ+
O4QAGn4NNaDIJMDtVUKnpDM569Az2ovC4p6cWuZpYLKfyiUwBgj+seXSJkE7fQQY
80JV0EmfbTM9XBHX9ZMcyPRbjvZE2icYYgwClHyPYnwEUo1IlkBqQ5Q5l6nAJ315
k/jwEYWoFSrQ7VA998aJ4Sd8T4Hg2zroE6hPhlbGNf6sQ5VmxboFZJR2pAUWEHX3
Y7pf8NQABlH5adJZdVO4RTyFKVEuj4/M96myzlI9sO9dVBx35kl0gVsLcNFB+qxR
DMsuzTw4mw+6yQPzP2YyerAUXtTTsMlYaxjnb/FAarNzP2zG5o0czbG9nI5XndQ5
Q9WhZwzP7isHL9ZUM0QYOMuhsXD64VQq5LTdtdNyFccvOPEwI27EHjzrlBA5cS4t
k8yFbDKjzU41b9TMXKWOPJhBwcMgEs2lWgNM0EuroTHA3cFbgCKm0IyDL57E4L4U
dZMJrvb3w47wgDeb1wBl1Y0F/LceI+lvhaVZRRbedrobitZP9wouRlX6Q/5SAQBZ
kAEQXrPlM/craWe3CbneHguSRALOXVFT+nl096cKHgvvrKvDDzG4pLd7HRmF/4yp
nBchuO0cdkfr9n/fPoraazuMFs3CaakIqHflgo9M+j06kn/83sjZ4Zj7rSWGUfVy
27S1I7W8WFPS4KmFeJc+UewdbABj3ggrML71/Nl1BP0Di8JH/Bat3744vZDzEOeT
baCENt9ZdGakstNvOkTTqwIMPyGorZ4c44TwoxvM/SstqyvObfkNJOTaZyYpf1pC
bxEvE16vgs7E/R4aarsvm6oRClMwhr712Ke4X1trkeAjMmnGcKge69IOqyHAYera
AgBtrwA2DnKyEoSsJ8BR5UkjfiA7jbs3Jf2zkxyC+BVRRSsmxB/kK5pioIw00quI
TmFzam5Bfzs1eJmRzZpW/yoHuWnp6r/5CXE85OKzGjoaRmUtx5km725a/3L68nnY
EsxNWYlaodgv39UUASoBdqjIiHWMRDRzLwXr7WWaaKCuMyPwGDP58WHDdxnxG2op
YmWW8oTBEdFBIu//rYJIvUfGcScMkk7c0kmfEacbx+NUrSe3uL77YQq15Vd67aYG
dh20T4BIXTRXAO0FXuyY5e/Fo4BTHylBrdH/KFHnknXKsSqprOdgXqu1NBFwr9NA
xn3lKeyxC7WZsP/qU2/4Ob2UmplDp4H3NhJ1KRjjm+gyFEPZWGOcYABt9dNsVrTK
Sji8pKQZFF5FlOWZpoLDyTurHc51EmeXQCjaLhSLbTDDKOhWRQtUw9R1zae7leOb
g6myvyIMSSzdVXMTOUQi19phMrXFZ/TEoEg7kOee7ITeGYay3yHeXqzyuQDOcZlD
xFjWUS7/iUhgVu69lLAxhBGTC6k3IXdhpACAKzKrg/HAR9K4le35GGsDu69NPll1
CAmNWOuetKawIUAuk0xVKzxHovMIJUg75iKy0t2Lov9OKJJH5lv98H9rMOZAQrh6
glU+V3Tp03Ct98eT6dh76YovIlHcTR/myHPhbANqORNhYCG8VBW/lcSiZ5+if+1X
z2F2ijkb/1OLnmOf7nqibuASbH260ZV5U0vuApvwvtSnsHIA3R3w8ANn4/rNUl2b
OJv52LpMIDblfx5Oa1ypFyADJxS0QfMoqqVGLVdztcP23M+bNn3T6zzO6HC5AVKF
J5jAPveGlbj66qvaPcq0Pn0Ic6s7fS1JGDB36rhpfUJormefDkl0OW2j/qShh4u4
fDBYuV/+oj08wPEwlLfB8a+1d+z0VIedZniO1n6d0Ifp5WUQv5Beq/NI/5VhWFLm
SjuOQ5cFwWXq37H0YShqe7GYy3u+iMGOoVEDx/eYCnbha+AsDCrAXNi8Ha3fj/g8
KKHMfSZnx6A0UC2fm6L3vE3/6ysKrERM7Oc5z3d6bWoBTvO7MDPDZdhmIgdcHhLp
GYbd9Wd2m5AYKpR50LzHGJuC+TijDBa60bMnMdi64dLiiSCCIhkAZ8K8q29Q69E7
YuZ+oh6CoKADWH35BSx2GIUNMTk28eD9I8/mxyg4o26hQrU0PJio6elAYUIcyo38
ZRo9IS/DdlWiLwKTNgGcKnN6hf2yFy+jTyU9wXMdpI/YhyaeO5vITdCRHaqWhu+Z
Ysdl1I79mM7/xdjFZNaXsfV+1PD8/H81CAX+FmYdHflNVErz55NYlD6yB4QhYxAi
c/U54dm9CQ8oqVm55BG3ZnbaJVLaxazzb/qCaOQUDkgvh91hj79FG5Y4NcnTz/AO
9UdHc2Is9h9PSezTL/pCQykvjWVWaq9Ddj1ivgU3UX6514Pn2uFdEx0OPRiDy6R8
4g3gfryE3sHDKiSxboVP8sx/LwdXJLHSobj3OBUDRUaioSFD7Vv4jR9CUj537HEN
lfX1f0lVSIXTHu8mpyDdgl9gLvzBKWil0N2KNiK9Eq5TS8odmUZ8NEl8a3MDsm26
D+jo0a7QnD6WqF6trYQP3MAtQTtGTQVi5nDTFl6+x+FX2fFbNUPDNFqhIVgwgelh
xfoBnzJJ6VUTFI8Y/6qERfwGNZklVVSqBGF0PKVtaCR7Gr9KJ6YKf2W76rk6d9Jw
pCUtpzCyzsVBzhTtJyD1YR1LvOg0TujQN1OhRRi5rD30FKe20T3uMz+5Mw7KF85V
h2EiDG6f4bz0gke6CZiBjqckWIxgcjwa7eL6rQx586l9Q+GuSXHKa0LDgeW4keEW
3W5nY1v7+G2ErW0+OcoslW4k4K9S/WGq7hGurQ9F9WOFXCqZQvqk0T47pyGfxrV9
IvsgGOZdW5G5y0KHgqIn+JO5g6+kNRj5b252girdyh3GyRIlL5HAHC4OBx5wf4av
WO83lct1Cqtc3Xmd2xvpYrkM26/mxOrVVbedSGIh6T6pCzejFY3vaipyZ1uGQgF3
lX9+PwEuccd+it0H79bv/UhZTkTZmrJa7ewTFml0hRrMH/a31woet5o2HvP8h80+
IUv8LZWpfw3l2SPTfaDdSw7s7DFAF+4xVHwp79wpfGeI/vv2BuOJR5SdTPqg/cxj
772UlyWorvGiKK6bbEdOkZZEgkUZfI0/omrDvpVCjEhbFk4XtpdyAl2/9SN/kHBG
jaUQ73bWx+5jaDhrPW9M+rY1iKcHYuupPQvBEWgv6Bwo5MOJUXWlA6Yeky+RNHEB
I7xgF2g8QfBrrwtukd57BqNmBAXJPAsjT/ExkkPnotYwXOnUBNI3tzmdhj/b1yxX
7oFaIM43+gPe783YDnyLEk8xDOqroPSKB/oUHdUIYYDIJF9M7Gvd/uoxf+Offdzh
Uhl+j63zZx7c3XTDdKBpQDQlDqKZ+NCYqn+gaL9KQGeu5GT8N++F3RhxHtieJdlZ
wrKNluyLfD+tV6G09PtEsmLSuELG9l6OEyG8kyormcgf9mJ7UQrXuzy9qW0OyhWZ
hbYHlc5byqZEWo2TeXHxLHIOot13zZcf2JYRLo1g96IzHd99I3y65FNDPwqIE1bs
nIgmzcld/ewfLK0H1jH4lMnVvK/7bWPBRJ+A76UfG+TFcP8qDrDJQ/S9+7ks8cYz
hXsRKuKOlfntMEq131LW0qxpDQTQEKqAy7xHgn2ILkIYR/QQCIAQeJF6uGOj30gy
8gV7AS5w2N9S9NnGLda+f7yfVQpibn0j9c2VTEO9hkRmdd9i05eeUkkvxaXoTSwG
zoi65IqQRFkr4Y6+IJ9fIRBSVgZPKtfGtzAzYeDK6asKaYH3+Vtt0Coxe2KR8geE
sxPbd5oZ1R9nU2xkIvXxkeqMq4op19IhCKXjYISe9HiSFAf9dkDIJQHJYbdrmhe5
wUalJKW9KUpkzNTpjZP6LQXp/DiXyuO6p+PJdUabyVWtvD04PZOZGRArR7pv02O2
c7cUep8VX7NME/r1IteTSFIssvpFgatq7XtAOuBF8I4xXsUc7HgF2GQPc0mXWbzc
Txk/IAZOFyGb9uyd0en9FpeUb/CJBPfZjvxJu1pTY8PTixqfmkkHR0hjd303jSL+
cY7b9LzV/lphswRvW8UGSjkBPznKnnD9EnWebVSumAGeY4S0wyhEhUROc59HxpfI
W+sqKN/JyV8iS8P3lftUlcmKhnG0n3tT0lnNNc83qsNiYc5xiI7zvBAGlQe37Wsr
hy8AzLtRO+jyYxMyHTahOgeNaXLfQiR1FuReMqemhA9Jg0TCSLhhZf243HSjZwTu
7wKoRSkj66y72k/QsuBMNIotukaGnczGlJc6KKEeGaw9YzfRL7zdWkgDwEf+qHg0
2HimF8hx8xJQsx8sSP/mgNXN1x2w1yf7ue2QAB8FemHYghRkLLZusOlqd0LqS8AS
N9hWqVt8PIWLNJMY5+SmvTZluSoKHmFOsJ6SZwa0aXiABK1xVgmtQNcEmu8MxHG+
lW/kIzT3h8GMcCmSrH0yV0nL/nnQ2V1LKvBCW+0lmM/+hafOUad26qoS3pqo/gp/
Jncmm4sSpixxZhjWeM6tB6AG5NCc9svJMqQON9tG2bAtDT953xCJbhGrjhjbHxik
vX2HTkPmUFF3ICz52sHFqo9dVtlaXZQzPbN+7tP38kQTNsZylD3I7WAEpAVdFU8K
GNH/tHWgQovGNhfP0s/fG1vCKJFwyScGO3g7hQT5mrW8oeOc7pkNkLjEIqC553eI
zKHEUFT7B20ZjlhlZRWFfe2FJyrixCsWF0qWZZa45ATFip+s0x5vbcGa9uVzJX+7
gbnpxlAzAeYd76CSVM5HRUTdOt5EDv/ARx6L0nrMPsQ/LHv+xV2GBKtBVHQhJsjW
RBLiyFHcKo+y+oMXQT2sl4iutZ8qbGuLBlu814g12tPSfpHRIww9jLeTcSljRzO2
A7IpQqrCQMprNJROrQv50rkwaWin4Nqlk7pWcdmTNjvdTZuAUYj1C9TshN0SQ9F+
7xyAm6tCeM6L6toPr0FrSY1krhFAGuzXjoMfwlJGMOwcxURkUmnzORYdq8nbu5Hz
VpPvnnDVupuH1CiI3cSVp7unoxtzuxrqsEJwjyZN44u7+MMuuaNGZ3IC0mC8VwOS
EkoRMcBNZcOgSx291T3YTrvvgWT5t7e8vdzlg+/tS5wambfhe/NqMFCYoUN60pxg
CtgQ79R0FF4ySzPA1ItVIxkaM1rwKpNpKDYI+liDtfSP7kNUDz7nurrZIpZYdbob
pe5Fc9eYzC2mCurSDqXzLCd93NOn6FcjIelb4OPE9tnbXNZx7ft7Pxtz+/BkU2Wr
g5tvdWDgeSnnBaE3WPqgAqLWC7kEd5Ssw8gDaJGBPWaDI/w1hmI30KIW22UBR4bB
BO/Oz9hz4CNNFPt0wIMNoouc/YLHAA/NMXG2QNFYg1HGbg+jcDkgJfqeZa4YaABC
zd2PjX9JeOTZ+f0n3XaWv2gGQ42UypoRF8FAStRbIgAZYLDske5mwFHFPT7Z2OJj
BPAz1iiv9VveM6oeRnFT4M2d/Bnxq02xezyv9mqOoa93x9oj2OdqYVY7KHaTbkTP
z3bGyrH4jZjfxLbKt3tFEKEDDkqhtq+un5/UVOecMhFx1aSnLaCaSC4L9wFAPlru
zDp3YM3R+IB3JIfW6pl6jwz8LIpKEXm1EthIjsps5VGEo+Nj8k6VIPGuxQINrpWC
vazQAhdsb9keccafL//rGhU+p+biFfHMf4pfRYrqL20iFg/8mO/jM2QNj2VSIMrQ
L4POYgwvYQRKYdrFekjvuyZEi6paFJl6E/NosVp0djnchJtOIxlx3o4vdVro6uDL
kVcfW7nFomNDU1UnptJP8P1cS4y+/tXWQPNpqOBzZMNCQLjopPP4AY3L2ssKwWyl
BW2ciX2QMpNc+GdaJO2pMFiagEO3cBlQieZX6pG4oTTPmie4mXygwqLu3zQNFlyp
ygGcvzxZ3LFDhGcBaeqRaioElXALA4EF9KduLk5WF+bDw19QpoePlBglj1aqOBRG
9FnqEONbaKp/PPD16xNDaR/Df51KQ+D3Dey/spxprc+knAZXR+RJedA/4krBPRLM
a2rGT4L51ml8sElon+BQi8DLB3j/BHPR85Y4XEYHKif21ONRzO6dGp+UWTIOnA1P
b1AzqI4yfGHjiwGQHM/FtaGvgC5h+jH9shcPDTuWqdLqe5h+2PviWxkZL80AzypM
qq1eA3dunLFjO2WD93rBBTEKH39UeZcBsYxy8b44xW67VoOtlaQTu3/gGKgjvJuh
HKH+Wg3cdx04bYjcfOuCRv85TuATkKvhlwbYU4mQRItxOl/qjQ109LLQ46kWh3Ze
tmIUWui9eC3eUrVPfnr6rQKZLl813ragUt/32PhPuyc1oU9V965UE5w78r6mO+VL
Ey+CyAdFeSEKSvoH4uk9yiY96bdnd89RqgwPM2bHoB2CGJ1NpcXFTU8rAk9XXJbm
BSFr9UcetlFFnfgHlED9Ai/qK0+65OKvRugfKBLdR9TR1UhhpdwSmcrlq2Khz9hx
CdqZZVNi/UuIeHFQN10zJGxagY8WwtIKfOSanM6mg9fTGaUu5OCiVGT7JvcjUSIP
57c7+HgFsM2Qi7HvPCc8GoyPbUIWg4C4pyxgHVeqsfnU+xp9XE+XSoyH+OXxQgC0
VaKGW/NN/Q89XMC7H1QQQ+ivbQxEA+ng7UlMkUPs/EsVLdqhBVamJPzu5wi52kKC
iJk5J9rx9ZHa+2ZtlM8JoQAaENiH15pgooSSk4ZA328WwcghIxPXVFAWdbI/RbYR
KaixIDmPCy2/f3ohEXY5wAQTdSLv6oG8/Lm0BO6xn+UFv341B7dV8LFmjZiCjQ9h
aKJHWY0LiwoNhkCanZ5jf1sgOigi3WQnK+sIilp8O80jvx9bxlvcvzVEiYgx3YGy
2MTbzAsYK6co54vhmnvvWSjgSCOZ/vAR9nGKqS64HLrTlfUaM8Pi+g3Cuzah+A6T
W+YywisSPxVNlW1NPU4m8lHWdGxWu6il1EQux7r/XISbTBs9zGxn5RaWxOCbP5wB
rUVkoy/WOPAXGPfyaATZkH03krO2Tj7X/lP/zDpl5jDWdILnsn+nEx6U5BKb0xsu
6zWOm0X5e32n6531OzogCUTgc1hsU64Mj2Aqdt5QJ6QzvlNWBfiCmvull2g4PdmP
WYrpELuAGOMXK+892tdm0dxNm0nbYXVt5Hov2T875tjE69TnIpU9vKKUvoIRbh11
hVEP9ooPL/Ni7uG9m/OkvNISZLN7CNfCEhKnQt0zBUvsT3Iop1E1zkU10B/bCYoK
m3FslvigNXx/x13vmFHaRuiIWeiwC0HDPTKaOWeqUldfVmhuw+nl5jfeVN0l9IFK
TMPVrRz2ZAVwI3vg9sEH+SZrN18B8EX/Q4PQbMBO5pXiw73xVf0URrweMYH1uixA
H2pFVOqKcDWyr2l4T7+C6zV1cCl+BwxkQt1tf4UAUhbtKTrNZ61YP1ICG2vxTQsE
Z1i+Pi8hRqRgYOhgQqpxpoT0/XJjivNZ3UZ4sYS7v4TBZcA4tJczdLV9PvIa/xjH
ERafkMIRU05isNUIyZldrmdxI0/CnPJSCXIzT9bRfQ9QbhSimtKD0domy9IZ73WV
8GeuhaJc/HviLP77udDijqBZ+L4W3VDYcXfIyItWPCzHP+Fo0Aytn/+7ShQfP/Tf
FO5h3VQfz+RzwSyBIPjQu2zuuT2h2bk30uaJhtp3mEL/xCWCMLyE3acsj1ML/lTm
ZvsRf8vPQE1kbWXfni5UF7TptbxirEHlnpJAJF/Ym/HjsWo5JUyvROf+t9P7F6+K
htqHg6kzD0xT+I6FO2Er2SnsoIBZviQWP60ccnnEBGeyZlk7QDdiDpWXYPYDROay
RMYj1tDP1wuwbgEHlEKETdl8yHZ24Ix11CBaRx2BqzFQSti3elg0Lo8rpNmrSvAv
qyM3DMX7afTqTwM9v433gRr0xXK+7Sh6rg7O14tBqjadTdQr0/NW4BnDJBFRUfFo
xkJy9uhh1zmyC26kTzKfkn6QAOkvrgXueMM0Jl1PmlwdH58wEwvoHLAkFja7qZ+w
4sXo3qoe87rg7bgGSE5gVmntg3B/F7hv5WuRcP/5iAS3v+Vxui7aGEwZ3lOdbzsr
wZi10v6FxEV7w/GoShjOXUwSDB6Q3P0RT/7FFpaxuqI0SKmB5zzU8JqXW5qtBTuV
swXe2o2KwwcgAHp68aqb8VM04fVguOTqqse/rqSnZFpadmfK+xXtlzyf38c5iKH7
lgtKtpgJ6EaZ9lGO1Xx+6Sk5ok1A6OtatBm4BX1bp1202o+jwxjzvK0bFnA3nVtE
yCeOBMYueZ4p5uQqhyDSkwyqrUDjIiLFfFSiOWW1NCtNLFfYlqxFD1vQyj6JktQ1
GXNtx2UQbXV+GKghctloqevK7bWKGJvbFXxH9JygOL9fbTYAtgc0Q+68657Nz2Ak
WUSWD+8pHDPdNjI5EBQrI2vD2Uyn7h5a/pgCi2cDwud7vNcNtW4+1h9JrC9S7ab2
Sddo0jvs3cwmxnSOe+WO9rqI+V37xCiAh4t/aXV5WDQHWkeRrjD5KlI2MmZyrmDD
i4uO13+wkIKJ79RXIuI7rSpBdxcbB6iOMetpNvPzATUetBWgl5R9al/ty7+IUmuY
mfLp03bsXsNJ2KpLh/oBooMeBVm7GYxTBSaeAHh/Lt6aeG7BiT+KLdSjTTE37VCC
yo4tGKpaBZFqdMrezKCmlZUGPG+oBUYqzyk/EnVwvTBa+ElrBwSrKJZWghqZmWgN
diavA/u6YZJyBn8Jf/YF9+j3XoHaSj3R9ojJEZqvdA7aaZQH94sUZV3HOqA3EoAc
aqGTE6ZLpcbV3ZoaivEfShrXZyqwhXkk0hGr97taoiQDgNhm53Zvy/eJQjGClSPP
0PpHxyQ4jONZR4Cg5UrK5/Mq/QfZw00XMvvMJBTr7o+l5NF6ebd3nYUgZj+gBE/V
1xkyYeNURhV7YYvhMP6uZ7KivcFlQBziUpp7PZgLuQKqDdJhJIUdxolhHvyXY4iW
pFrwEwZ3s0XBdIlTAc4sF1YTtt5AVHtMqa1SYsHWng0mvKhAekcVWPHhIMrr9se+
glIXk/wNLufpSpeYPEX8gen6wxXOlIEf0nYg8Y50bvP7lJlQ+0JhhyjyurDFp+k2
wL6rRL8xKxJyATqr/jj2aBN7lhy9Dg+w2eEu/zvA/vAMvQx/nA0/9xziNvFUkxFX
OFQJ/ck+TjWrVJUeyb1BCpJOhZxz5TrgHlIKcCoraS7SH8I8NCoIJPwDMAN73jWr
W8O06iO0yUfH5EKQlNfNKObTpixLnivUtM8VJKK11L0pJs/nGIRiX/N/5GUZYy44
7pp9qx+iUMxspqst9wAAczJvDybL7USDMSoqlt3vpacuvY6LKEgFfYrF0Ksi22fR
n7Wn8IV+EIUO1v4auvFLY0S7cI3eHPEbSF6E/KKPpq58NlsoIptauE/GpYbkS1aE
IaQJ1j0mlMTkzoMpIRtzJ+DpGUOpqlFdxTc7mN6w+weNI+6du+j7fQnI2bqmQY2f
N32801ZmE+nyekGJG/C57yUo+i7bXG1O2YDKWirnydEOjNHsVvBQN7FjHcmrQh1D
vmfyuftpSvTq6Iv+fV0uIRaUkMds0/A2uNVoz1IzoCRviCUjoMIs3p3bNRUaiLhu
I81C000IimaljwtbtbFPbzkzK/szw+i4LGhlOHkBYXxOAnwe/7RHz4MDBuI2AH1r
QoyGElRFxSelqOeAcQG6mpKDA5yFOee8BK3cGNtBPGKqwnv2PIwG+NaaM1AGQK/C
PVUDzLseB2Wq1lIKzBJcGdQT9WLba2sykONZp5EuUVBVnBkoWWC5aC1cNKwhnSUK
JNauLqb2kA0jH8E/bLdROW0kS3db4GiDb++iaqj688x01Pvyj1tX86boKhHBr9IR
P4JdpBSch5GVFQ78khTJJHGKOgsiJ/lqerE0Brc7OOfQEU43CpGLubFl9DOEJU0S
TbB5FG5TWMHFX4PbkzFRZhnpLw5AMXW9i34wt15CGG5hD+KYYTHZHcBQuV9Xm4Kd
RQKGOX2dPySUsaCDEVCdeKhcg/nkMoRzytLdpiZCvV+X2FFt4iJU8o3ad672mzYM
EUzs0E04ZRkJFvvshplEkKE3hQjHrWaCD8OQvpJVS1A/kba2NH7v04rSS/Y2TmpN
7tTkwpNPr+vf0fN2k9dls2FPqT4ZkzB8fz32aMv+bqv7tBK/4AyzePx4vgP1l0c9
tYHa2wjSZq42Q9fWGkNAu+3dQoAOUglc2WnQrrMZ2gTLZFhL/tAqYa1wQG2zV1NG
NucHyISsiqI9Gx0cL1KgHLnu8orLykdxZvjZhBySn+oNizkjDzFp2fl1d6bhYh+A
LcfQ85kLB+kljO8JkS6iZN7X0OnyVmRufSNujAffAi3/0weFLD3yqyCL9qTaFhqC
rs29BzckG/EZHihoW5RnegLG2YzCUzOepwEXQfZ1zVi3pwYdFOkS25oBuj40dp9k
hifqJbzbs4zdwB3yUb21AQXjEWU8EELr5uJvJ3TYCrp6RRPVJRsaVRZ9UKqI6ykp
x7UJJOmJtseprVU9iV1fbIsf623kCQlZ13lpC0ylGWFtW69auwQtqYfWiA9J8h4G
aNFS1lEsnGpTZMYPOxeVequqEGYGsq7OoJVf4XVFAu8daU7ApWq5Sl4Os1AtrPCX
x1zczzW/hat1RgjXSUIOoh5pGdzBUhde6Kk3CO93itTsc6gH7Phj/1yXb6W2BwOr
+OvKFKe1gtwq2RoKZOKUu7BWAstqzvx0dcY3TK9JAfyezkGKGrJYjkArMqnmLNUO

`pragma protect end_protected
