// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OWltXuEw26vmvykWbBfHWm8u+W5dzH+aAC3KlmmudsTMKqD3YzJI1nfxfogf
ILh7o5iPpkWTD6UaKSeq0ePk1/oIFa+XWmMcLp6QfGxEM9r5+VsNQDSmRkFt
bXrWhSVjeklTMfb52Dts+gjX5/3t6z9jpCRYZ81S3WGN9hHvFlYzDHB5icjO
+RKW3KxAuMlDxRYafoxqt/V2wloYoaZO9Rx0RmEcuKXAxBwYUB8SopR2Umc/
ePps0vTLoDgg/5gGr7UTy2NgEKy71O2K1xHZNojD3fIVi3UON+oiSpZQzQ0V
gA/KyhJjD83tpryXRhOxasutLE2pIRH+/JZGnbF00A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XQiAdu8D9nlz6p3C/ac0CneZ0T2UbNnQes71yO8jfv16zGru5wmQTUjeDA4K
iv/dJrQMD/gNHKRT4c2w4DEIhTHAVR3sh0kRB+jkNq00oVba2AG5eRSdnEr2
IAuOyu3vzOWtG1UZUwljslNTTTlH/Xfa4GJLbPtZVx6RX14ydGVnXwhqXxa+
OjT+MlGP2u1sAXDmFFHwklFTFPyuY4yTV5F44/Zs/H4+ekfUr4/WIyjSgeIV
3aBVOAtN2Bq22KIz5rYX3zBhmc3bbxH3AZ40N48Ir1JDnKJwSR5Yc5rydpdQ
YTYqvV/QdsnOruGgQX0GDQ8lBj3Yee/Nm343Tu/VVg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pqDi0ECAe6ZJBdl53YeJQvZFKaGsYuRULPULcMd9DcnNzMD9KGg7Ok6ZAJwP
p/fH/5ckhhhQMrMrj9VhC63n3WwDT9HLEB17zzuqUuW46T9moWOGHu70RpYO
JTVkGhCjNb5SBH918XVqe4V47gcH1Ew/nrDrDo+I1kxBBaL90wW7e5nCPeyM
jo6X9fK1MVwUG1RNgwosRPHkN6zdHg+9XbUxnDEuB+uUYOmgF6LtMlq8t6ic
ww9rXLuXacCKpI0UA1cNGj7qxRrKvROBknvhqMGt1LxqqGysEfCjtKDKi5WV
pFlhtSDgJWObacmeo/EBSXemawdDFX2mD8q3tN2VzA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EXeqbEwPKchDwg+TUcB5e2HcaHUplR5ed1Obh3d6VNtuPaP6S2KC0eTRgBMq
M+3NFIqIcfeodNs9pnrsYlTkc2Wcm2Dqg1kHcr2wTZzNNaePd6j3AH+nz3pF
KWkDXTj7u/8FriADac2eoFHVbloV/rVXLK/fEbzKbaYYNd3aiXc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yDcO9GTnBn2s8prs4w2R9q3JL+vn+ly/Dmuqx9TF0VuN/TASqJGWO9oE2PUN
gYwtGCYDyjk4B64U6p3eaCjg6gq+Kp8UBRoNzxCoUCQBSZWHp3gvXndKKKdR
1rEzsdVNZTBSGSzd6PLUMJ4rTYFEAFJJ7pILtwvnNPr2e02EBcQI5hcXk+Kp
9N66BeEfl5fSJO/A4E/pCrSZ48Nabk81U5/7dOnh2KN0rZlhycFJgxKEZwJW
obpkXB3exlKJAC3OCBLhaCB9cyzzIOESyvCB+mYGH3EWW1FH9XLrx9h2w6CS
iMXXuFmzAjRGftNTXR0Cmb6H4uKk8HTODh8KwkHVtQIG/neYKl89zWGvM9uz
PXBukNkV5020qTyO2qPJxOrdXH5T0prZOFDUXwcJu11FAZoSJjYZKb3MzRqK
HHWg8RHSeC6MZfTHJo7ZRUmeYhZQOss1AWOjVrZ5uhDDcQM9Ev1x+Bud3QKR
TndqUPMjV0TkBxbk7pF9ZoA3jHmo79LA


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W04V7shHg9hiybWedMMiZX8AHIDcYtKy5uWvWkOMpUIcB9ST+EaJKKUi0wDJ
X7CXbH9FA1arRMgBsW8NOujHoWfc4MXErqZ+rAGnmvE9AUgYGB7IOUCQcI97
X7nIFOxwCr7fvz1LJlVLn4/uXLdghY/qrjDp0Ti32XMCeLMbtxM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IFqCtBaZw4su2zcXN4m66TfzQ8OMxS8W47igNJFGH+on0bv4XclECV0i4vD1
ofU1u7G8e0tfgig0XwlahKArt4hExyXvw00LA7rosXjUD6Jw/8iE/NdbJotH
NF+/889WAwvjyjHy72MVt/u9PxyNGOMvzNIOnYwwBJtI8C1z5CQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1472)
`pragma protect data_block
CNvfjs/AAfyqSR3cogw7DDzMppmvyj7KXMfHKXZEFDcDvly61jxhg9H/cLtw
/2t6h8oiyUS8XRlWZwvTp3Sjo5O/Ay+zrBeERqw7cYo9MUW6Na0TizaWGcYx
GIjUrGcvSBGVbpVpXH7UctAtIu5ng2/qKx5GGVAY15jSmaA0Xe6AExst/Gpq
qFv62pBPPrbtenaFryP1zvozG4GK65HUpB4SRPgiVgaqZqQx87CcajUOWKuB
alUTZ9f5QiqOcgy0XU1BSizXh2sr6Y/G6KmBRI0A5l88MpWIluKWpvKjgKx8
t+1Uo0h/ZiPAh6MKQ6vZv5rjg7UBHKHRYYHTgkpZZxoWCR9HEYBaN+V8jGSv
DozYtaneEh1/OHWZ1sBizTi2DHvjWhTsfPgurSwbDEC0rGm0JC6UID97Stbq
t4rv03KUmtRUwMkBgvvJhqRIqzKKfD4pQMZAsIE8pgmvk2gSgb6tJbMMinD2
8WhecLicEoLL3V3uDkafFZ+E9Byb41mHcWC5/K8sgCKs22ATEdV6GqIqXszk
jIz55ldK2hAL77fTPFM/CfHzK9qBMR3Odl4ZCU4F8JV0YZvn/FuL2OQGLM3q
sxWi6ULWssFJ4Hm4CmNx6zfu+GuDpGYBTLxQ+KoS5eytbKu6+SmzLS2t7cGu
+lKT1UR0bbP28+NeUhf+6GtPzaqiR6dOdHAWmOcD6B5sgJRJ2MpokkAQpxhK
BikIrSJdhDAhWW2t675nc7yohc4pDtSnKIne2nmfP6vV6y30Hgc8mCEpu0+5
xYECNUh66I7gWsG6VK/3eLilIkFwfUrZfG2OyCnPpBis8m3hgA/SpiFVcN62
54mmrYZtVArGhzMsGMvja2js2El1YpIOmTVoUCBh/TmTP6XtfmA4FyAuV+6K
Rg2lm7lsj1GI05b8TLBkA2O0BdpIwTGH6tsfZx/UJ9gYeRUG/AgO5pvLLQcP
8NJipqXdo28DNuOw3B9rkSRh4bb1D3A8zybbkZyoEtCfBFSt3xG+vkYhIgEZ
T9H5vFEPJtnDdP2Nfn+L+RykU6pEIYpjjPK69J0VctTubZ3FTtsvYTIfOKAv
jOiT7Z7mCbvnFA3fhc+Y+tNlI3l/mskjlaO+lBISKMIxBscsgkJccZGI9LUv
13y6ZaiR2C8sdQyJ4PeOcKJHJYHaUH4gLtKl4j/esvm8voI2pDFB047/i8Oc
2DWReF1LjeINv7B402BBcBVPXIZIQiM2H1qWg4kvVAUo56pdAZuMgMEAC9mb
drZw6QGNnZ6zyo1/ccfGUCxjh+oi9EoSfhqXW/W6LPeFrod09iEVtr9f8yf7
dv+gVwtk5fdOre0jKv9mY6ENJCDGdfvTw4cwSsiZSNlS07t5boI91kn3JXcM
MLQo8iU2KxYoDiVRjFaovr4LByJgDTxaMm6CItOHDqFgBCx7hWTJRcF+iZCe
HvvuORY3BJNxB58HLy46z8D3lTN5TxUnQ/UW/jqPnQF5uSvBfJwsCNbH6yYU
xSFopZVFUqucbKvuMAaTauNLxM5KVFApgPi5MWDSE6pbUkSkIHzM6xdeGTwX
Vb5Zu/nU539wXxkiVUoxydPh6XewjokFROHiHrB+PCzJMqkmydNQzxyNvvdJ
1/jDcWh9VrEFPIyhkAGBjxQmJRwIQU/qLZzdQZp+9GtHI0mVhHJ6PXD1n4Lf
7OMzwyQ3ZJoxl19ipYbzef/3wzJtucqDACxYvrAabYOA7DniOUOrEkRQRgWa
9N8t3i71dD5o2RUyuDOT0n/VoSYg/GSOqD0I1O4JvrJYW+XZfFoCasmjCu4p
75FDhNdXcjWpCoAHS3/tVsg3MAaUwSWfxDw093dnLce34Tiw0F86I2D7x2EG
AkOSV7wJ17IuqOcOI/t3yElBy1UqxoO3cIynXhrubL6IptLm5seX8JmF6Elu
JSrNNWuwKqM6ppaadxlRyRNatv9gKQgEJXqZpg7ovAQ=

`pragma protect end_protected
