`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
XFoK4u28/0beilFgvhbtheXYeBqZUvKGjKElESqzqo9M7tpb2brlNMHXTn3UO0lx
K/v6rd2ZZxvTUvqjYVyC9PZwyP1qZlq8v3mLLgDlnEBgmyli0G17dDnhgm+2TO9X
MOaV3h1au3Vp2+VOBNjxdRpyif68PhSAUyhrGaoTzak=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 25808), data_block
J3Qpws+TIpXsdejzcQiphwUouHoQC4kA4R3zDMzWBWOPuS87FdmG1tDdlzaxw0tB
IpNK9L4Ih83NA1/hy3QipxWbv6rBe5BKt6aNnrAioXf0iAckoMMw7Vu2K51ZuZpV
lT8x6of39tDUVeMw3Zhlos/jCtcZ0qTMPtFU5BX2sdpBd/y6sfIse3ChVcpaMA0z
vxisVzdQp7qrVA8mjZyI24wScGwkM2a6SOVZJMJbp0CItq4bGsoo/7EeyXwraDOq
h0qnBDilpRB32GDlAlmrpNAjSmbCtT6CdUJ91MGE8Cl/eqMGRlJ7pMVPANAho5BU
QE8avjGrdryx2hey918MXW+GaNH19x7maMtINJJXOyYS1fPQiHGQ+5AtzBxkZGXh
Jh4vw7mVjvDpB36xvhDAo72VZ3GLQ2zpWIPiAfL85KYpZeUoUNNfNGsZ/LVcwGk7
4yydo9rnuRGxPXjJtfTOF68ZfMePORs5dsP+9iD+B+O6xdEXvob7lb5WWUO5ST1R
gGeYcbODlvSBDK0KbpdUMKesK/Fo/zFanp4kX1oGjPeE5i8diKzldA5mivuDS6+X
tR9jY+4hcJvgMmhNrtzUzkNDkUqW/X1wgawdGLR5lL/Eg7LYJhTQ0FvqBHP8l3uv
C3QPFrpwK4mAa2WZ+lo3o94wGf0LFMXqICgGW2aDI4qksluo78yqvAHDpVx6Bicj
hzkQugyKgYvbhyPsTgSl79PKPb/uCjsxxrBndUwQjrJGxKeH9Ox3XUGwu6CuPV5y
UR7gxrmeDv0JNGLD7CpWzc1naiLcO1IbvR9znTIIA2wOc7nKCHHFFjnyMSFAGJEK
GCiEAS6VzkVTR/AHTHha5aOOttvurfI6jB7xE8olpXygWGcxiQ6O4ltwAAYNHDXJ
KHV8xha9ig7hKG5xzlfGp3Ua8NaJsLSp/7UUhIS+2iWw8gqM1GP/LizGlGEnqClY
7rxk56Y53vCFSkelCxgOUoKbaLTQttnFd8oJJYxwvSiL1m26qQR8yDJvSFahuWoy
T43j5nWfM68emypofurdNnnMazalSsd36GJEum5ZxgwMWRzjCxDUU5fKPVSlv6P8
kiGFWQ1SBDeFkQE0TuGKEqqB2/l+e3RzPlLxmMGyqS8PC1rTW5TfojWJMyxwFGZ3
JSypuDWkgyhQX1NguyVCMmd3zR7ouxa+mGOb2PmyIUhTw0hVEDCmJIQX2xaFHBqz
jNTa1U9lMwYsOB+FoghOQm93qn7cCRqwRwv6GXlX1SEjlRo8+4Tx7Jl04rG91FeY
vm6ubMPIuGGqqlfc5jUxxSYQ5LkV3oVcuXekq+P9DrF3czduKFP6nyeU0C4PvYzH
jMxLNL4KqBRcolEfcNhBgilS4sUSjERdQ1fhZ6vNmMfH3BAEwiGmmxAj0y583zzE
uLogyxR1Ld1sPSpgsCpqYbrHXk6M/ByxUgjS21hO6DVDxVXD2MlTpU0xHMpm16h1
5EHJqLPW4nWo0DbWeCpt5tLocqT87h25DbnoXCmGDOgTn5u4ti1D3xX0BgtrHt9T
cpJhm/wBxO1p7YXK5W6t00QgnhlPdieaH7Y9Pxwx5/u6FpUVK8tnBOyffVwwY+GD
7DCdX4wDmuBDw7powAAXC/aCrcCwMTF69TcPCHnbWgV2bh4IaiDdmQ/r6/tFwhDH
DuTRadJ/pHe40b7NzRNYRHskS2grXiV5MJqxZP11uzA1JUKo/PK64D5XzYa54Q1h
oubTc0KO1XH2hsYaFloMmoHHCnHFY+k2fbDMaVJKZgLwJSyPn6MNTfVcRFNATaJe
SaXLBmdry51z/TyTfeDpP0QC75LSXJNDBEtZ85VKgaIflR+PyR+GuDkq+FLR1Lqf
JBLSVab0yqlyco0LEt09ikT1bJDTy36Ym8/YMt7GR9GXt459/Mlsqki2KBssa6HX
+oLvPNhrQlnmWbf37jYyKd6JdzDDxFvUMWwLq8FSuM2tYpVTR4fpyJ90lIRGuzcH
ZYGwrwENekWsvz+e2Bj2NUJ97gMmbui6dFSUhgGYqr+Lxdz60qLUjZGQaBC3ezSG
cFn4+BKJA8jGEvAk3SS3snN9d1zJ0i7A7W4I90sX9MVVU/6RwNVgJCEvHc1Psj4c
FUe2yQv+zJX4NX4QKBP6CQVfu8FAQmSYdXOsyIRfWsmAW/X3AiRnh9YSOm8PniJr
Ciq5Eo/c7oANO8JWxUBy7Hu4gyqAgTN+lopRB1Bzisvtyxei5nBb0MghFAnG75Ph
e+TbvuFUccJaX135jjMg6ZPchLSzfMVC+OzUJ8hZyeU3uspPHhDi74ckNRhly0ug
3rgjR6xpCnNNbbTiIW7MdxauV+cuJWwfKZWAg5DFLbiNoh8qCqkbLzJVtSdHGpM2
6VofNWjfYgPCvazKIsqo0+2LaM66kJ9pb5WIUeGvhIe7rzCXj4Br+wT5yDauePBG
nswiLDZ8Ur5H5J1X/QWrJmi4ry/OB1GOBy5tnkvZkuTyxWQggrCr/WUdKXr78KkM
l8BAk0HbjpPFViiD3TaQI/bQjEvvGDT/3MKywxHzI6ehKI7GGFNSSLy1dIFbuxZV
Oz1l0iYJHnHyNvhLtvS1SHs0jO5TB5yyE2fmJERp9OkTa8diXKXcoObu83BNMbrh
X3cSuV02eFYFBZHQU8yY4Iu2t2Xvl06dwcDYTmDuiDVrUkkRb3klJEX6Zuqmatik
hCw8XTPurYp9aCFHMlQbWJ4ACO4uSBK6S6Dl3kyedFkmkvNtPXJ7mz1vCE7CXamR
fjaLAAcs7rUsXYZWfWSOnYEB/RlDDxMsAHeZmWAMFc0y4JXNyZBCM0Wsa9cDVWZ0
WwSniUxktMBHDFtx5F0yal4Rz97WmGBfuGkBnFZ7Uu0wSSgw7S2exSayl3GWl5qJ
QgBVsNPYOZAtFbxIMQhM7MVjnfWxUs+DMKbuXj0p1HEsSpTY+v4PCyDKJDSFk2wn
liDGBW9dFVVkTWJi/daky+HEdhYD8GFQTZvcuR8SD2qKMtsmUI0Ns1m5I2KM4272
KafQGuHbOBJu3L3blxvbHfwH4q2U/frTI5+Nzf2FLTB1jyC7yqsQk+dk8y/pZq94
Ndtu4+z4LKmBeJMVFPiNc4/y2dLWRlUYsVafllnn/X+Ph0hPiQcEhYqS3R40HlV0
w+OUax8nbyrOtDYMDMI2jK6Q+n+d8xlb0FuctQcv3RVMoJ8VdL0BrZ9pxRMGoJDc
PybhzVxTZSdks1DzxvpmqScA+5rme+4F/6fL7raQ77Ie55bsYLY9TMiphdfilBoN
0dP5vbJfvmWfkBY1/66fRK4DC0WiKwcIAocwfqFRjsv1u4gvsFy/ZJwHBcs0H+0U
LOVza5mz/M7TbFy0iez2Nvyya7gCAShdKGr+PSYZfsUtkNy5Y3yYYTzdK0de7x3q
bBCaBfNvYzoZsDf8sF9OSSc5ThZDTOA0o+rBXbU2xzHzSQO+3Jhs9xLYluWmF/fc
gRHtpFFUVfOWm2fp/ev+YsRcWCtolej+qwOwneJaqo6UeZM2HOgGDTpms+rf6TuC
Hj6Uj7mTmV5C84/AHT/LvoKNv/4U123uScOOaJUDLJ+FM90ucNQP1a5qZqQFs0U/
E75WkCq1rDKp4eMOqUde5coqHrc3mOxQddYx8neJu0ZhOcnQ6i2S1r+xpyxq17nq
qGMJxK5W8VkwWzcqUCN0YblwLy4IEaRI6jrDAJNKlBRr/yxA24hsqQAGYXrhv9CR
3xQFgSavQLFUUpeDTjgl3kLX5Ub/pMMJpMABHaJYM7vLdr4L/jtsurvcDMAeIZfA
MLUYqwqKpDbui1z+B2WVXG7D3izfochEq1zItQF91kuu+BAB+2X1KCUB9sq5BdF5
YLUChGxo9IJeVObS4TpmjS9pT5Ol0C4vShrWtTJaRFXUMsQRXSDJ+gX93T+YgNiK
b5zGz0i5UT9k2lAwZJl/iQrh4k0dpAp0unMO1AP01Z+F4P2iMHa726se7OtiWwml
XCyLkrCOImOdhLxFc7UVvqgjmu0Lu2wZC45E1LIZ1lKn9CoJi8BzmdJthmR/8TGf
oIO1pGOf2f3oeqad0BrifmlFSU4gqkhKVWfMWXPkbrLZMRoLdVd2Y7grg9TzyKlh
7U8KNe2evQufsoEiZRNlQmmd7K1Uq/U/MBOJVGYC/Haoa35QmyQ7UtrWkP6JVoGP
cCDjoM00nKR9qwHOffA6JuXs4o2Z2ZjWGlwhDCYQtKfZY5EC5XkeQyBq2BfpFyGU
NpeVQWFH7lCX40GrpABNfkmvCZBOvTr6rohhIGNrBIF7g+pUVcCDfMhs55EVyjm8
Lzw6l95ykw1tJjvFachl/eg4v0/hBGmRyHyaOgWOts53CuTq59sEe8kXRU8iLd5F
gEZJm3XCXY4ukhfNvYTMhOzW27429zxmvb4jpG2JGBo6/GcySFTVJs+KtxZd++NE
w8KU+h6KBqgtX7Zi4P+UDJwnwxjaWRo205TabK32tHF2OGnTn4i6Xjth0TiVKs2Z
mwIP5gcUV4LQOR3qvUE87C4aEEEKcdgoHjtUmKk9U8wK8aG2qj3XyH1Q5ERtaaP5
MZbJpCqv3gkMSBqnnDoEphj49pDQUpvpfd4LqQSKeS2bBGuNrwDQVDXX/cS9ewAd
SAMiVrB15UElC6NNA3EekV0fKbnl7UUq47y/NxVwaDb+XkPkeEYCzPMIQ2d35s1Y
LJ1rzY8K8eEopPooqS880MFU2LcSuDHYBW0rBilZ+v6RSS738msmVVBC1OzkLgw9
0duhVYp9c02XHyXoKmj2BHPs5dqUeRWALIg0UMAFUims//iAKm73RN8VaU/jNDlO
7X03nm7CNrVSH6wtm6nuzMo5mAZHbTaZ/YCaLLSZ48C9xudXWMLZJXrDGi8RvUd5
kHi1AQqZNr7VslO0RlLs+Ufyi7ORH525TprLCL5e5w/uijvRufnVwbxK8vUcTKFd
kJaWhSkCRnbWhbimRLHhfgIu82xZ70azuFQk84pC1b5JkDBjIvaOQDco37IXP/w/
pIG+I5EZilEU+SFwd2PWPZxhLqA6oHUhmhsaJQvldx+I+pTHvfPjNYbm88QsL1GP
eSR4/gq5fC/E3EAmQJAlhUJZEnGghdxgQXJ4d+LHkkzEvNEVtje0dxYEYDsdVYW/
0Oq21FJ+ZkiGj/89ktQuUy/4psL7+tm4rr3vvNM69LKn7kmdp5fHydh0ImDvG1pN
Oh/q4r5OIMy3tWHh2hEodTTjk5cGBMXzIkYvcgVhiESVP/Wnd6V1kX5p4fQ9gt1q
yR0mJnn/6LRENNrXLM4/V/O6xC3jJBbitrVRvlDex2E/9/+69TwyarzQYEjIFzHg
raa7KjPJHUMFTetQNch+jz858bzikWD6fbW5k+OeKwvYPc86W6FIivKXW3Eokbbh
w0hYBrPrNso6jRW2QV/qnYmJwJPUHzRbouI3XpXsDlNHCkJ9yzBIITu7cAxCLn21
SJ6fyc4cpCucXhbCIVj4/wUrWjjB+fajDWWE4va1SgikxfAm92Ykl8/yUg+8K3DA
cgsty2iy8ELSSZt3PDjF8r55DW+prYkDzLyorZZA7PwJCQU19VCiFPcKRJaPrzQ+
UFoq+RbhBCWQixKxSwNsA8CwjQd6EZa8WQPQAUOoVXs+2rB1r0DXTOWPhB1MlUVE
lynXgmr62IoaVKVlQFGlOs0WaMOM+JacGqVj5RsKeGvFuLeUftk0nm6TtloJs73P
issJG1/oi/Lsyj3lWPSg/kNETK2t8Kibun3AnxViHTB3l1bHyZZ8NUBX+fqWEywJ
36os71OnScLX1yci8stV5RBfIPOv9/NnvL5i/5sfPv1iX4S+nsE0nl6kOYt0gM4W
00ZB2sRakA24XFjvaNq6FdGuRQn3J0/trAAlmvaKgKtMqNX1v8JVPYKA8GF7Sz5U
9YOd6A0UphVmx88+nVRYjoLQiVbBZLlW5+XC8p0GzQ7e8oy68qWL9mW4pALQc42j
+w23HiLnQJNcsFLZJ6NI8H/gHZLQ6mTXw5MVc2GBxFI78UItbJrLGgYU23qD8Gdd
N5nc4OtoHprG4u+drF+VU6SO5audQ7Ny//oUncUigMIcHAxJJHnKxAZZx4M9kYl/
MbDGekjWSKSdVJGrexgBRyJscdmufVlF7YsvNs+jFyhFW/52Yt74c0lbEP4VJgoN
FZlTriva3KMI38qgLJQ3g3BcSFM6e/MDmBwUcO3hIKLUw7oSV7xu6aMeGpBzk/e2
j+A07yrkvNjGTSJb53V2OvoCp4sAHZ+i+9zAgao1oOU/N2kuRo5wOtLqSMhdr8/3
B0P7thzDIOoSKK8YPn4OM6fwIXI7RU8hdr7Ba5brk0r8XnPCc3uqHMAbEITt6YmC
smxCRG8Wpof04YcVFUp7RoHa4aMJ9sUTAHw9w7VQJ9SdNksRiT868m3xoQ4FSaR5
shkNm1FxEEj7++BNAZihW92SA2PgGU92z5yKFb5QLb4M6ilq412YoFe1WAukMS83
+zr/d5OUD0A3OFCnWNEJEhWoAbO4mBTcS2sVd8rUNDDjtulQzFJF0yUmvD1Le4Cw
SX4se7BwBGVei+zCapNNFvXLMLcIqIvNJgDPak+u85MRPXvbpnTZ0cbjq/sUzpiz
/yB//buTSWbAL9WKAvuLPjacHLIGrGE081brKRRXq70XwHrK+hpsISzNjHMdMoes
E4yz43dkMJwjHgaOFqVbTN26cEqtBtvrvojqDSJBZ3+g/xZbwEHzuohaYnbylFO1
M8Qtkhm3gpVCh//RTm/8M1y2j527naI7Dy0/IYei6pCAX1PPiR/CjcaNqAYC/oYZ
MQ0WP8e8CVWqR5tRIsCqwebrAYxOKAMS78J5YS/4MkC272QHq55pBvgARnEcwSP1
82nQuk9MKvzi7KPQBmskxi1L0Gj1BEu1xdSVDNVlyqhw4X3rUpeha5+DGhQ1gPyr
c9LtArWVxIAQnwLtg1qfbV5XmyUpM5NgptqJgwo4hnV4ECbhxgFhhCfsAteuQqO5
n4uJM+WtOjgSBA6/sIjeUBtoiBBypCIYpDPBw5F11WvtCQmMAcsJ8UlXiO1qdy9p
7wYpl8TrJPCsqFNDQmBqrLvBN5s1cCWFnguv3AtYrCJKXB3RWD4pYPwfWKYIpB2M
V2MbihCDGfA+rGq5HSta4okxGKdGfsUpYcsoYTZnA8TaJ2L18x1D5hh5S/S4X59p
UO84KWZdxmfoRju2/Jp5MPMxLUWb9qF8QTd9wYCAvJARETfHju3od+hgci7To4nT
vPlKQT48sVhjRcm4GSYHyaqhPWbou5JCseXFf9F4+MfOrhT9Bud9RZewheTY+NW7
b/Iogursd8YZcVnpnu2i6ePY5/OdD3P47BadfyBknXuKFrPhe/q1m5d8G2ajGIQB
/4e6NkL9gGjFOHivZyFtKmRBwns2fXwCToyBHZ1vA4tvZnGV87YJQm0+uGGqBVnS
k5fsutLg1xQt7Y6waKpe7ZsUQtwbrjZRgBFbs5S7DXKb4uSXqhxH1d2R4usaM1r6
4pXKaCPlI82efXFPD8FL8NJTvDrJDGF9glefxeSPyX12fRTIaCiaLU+cqutk3l6D
mh4nKEK6TGg86hFxm3wRNNFWnafao/LIPW9Sd36yAczDGGWaO0d8Fw30vkP707ko
7+U+hlxQL54GoiwPZIUNmWGMJZ5a7OLvDUVm5ibE5FymzgrMG/edf9bwwn+rTEiI
r+NlP2RGYKza7J3u2SB9nH9WFKv7swK2RFj8ZgjsXhXxnnQAOIbjpo62nxjgzl1Z
sWbImNCOCPR0zeAlqp/uNz+oKOHpiYSp0dRK9KlGMuN4rhmA/yS8ucMkMtepnZSo
6jzUWErzUKrGEplSIyZxQKiHC9r/neKbC33HQpoqHBQX190X8By9cJ/tSnlK4MVv
DDmM9b8ZzUd2OJvoQDo9ZgB52nBkmy1pQMq89ljnuod1MhxR90kZs65xCoe72qbx
yWbOAolq9YHC2N9vJQVFpCn+ukPJIXDfF5Ob0t1ERG20W74APKQZcwDwEflqqC/W
syY3RU9nb6NJuxTb3AGX1eHVPd39+Zhbd6czv09lZq/zI3KdKoUeRBky2o2kliG8
fpBxegVQVssUn5Y5dkH2AOg7ssuT/wN4ulIFdu6EQbWchYhOVgQNakGFWGlq2nqk
0vA6Zd6jubcUdxxKzpQP4KwbNYJuVCbolCAkjb6cIoZ+qf0tnSyVS8f9U3GpT8LY
S2hd/fRhDWJrcYSihAJq6azSNfRuUIIx5JJCTnu7J8w/vhL5xwI9QAMMusF9DhxZ
f53y9E8oXRiugmdUNfgfzkmrLL/PY3bd3wr7UKABsZFOCHRNNjhRBhtjuZilfXEG
8JSmuO7NQ3oZS95tCRDNSKTZc6uZ0kxOIkoU35RsyK1CctYxB0DTMO3WCH10cAdZ
z8Z+IuHYh+qZ5j1aD1QTYPpUY2JrkYrwnX09icJuMaQLhn5uqrIWEWiHUrmaJI+b
Qoaj/TwKdtZDyQ6UQ3AquDyD5kY4sZadpxaI52Iu5yUzWco25y9MgiJewpOPZNYY
SrEyCwj9iEG4DwK6/9OBUlhVUc4hNEDodDYm77O1SMYvu4TolW2p0H1z9U6H69/M
O5EKHAURq2LjBTEVSIdr9WK1Qjdhu+PiUF8cK6/b7rTFMzRFU3k/NCG58YDqZfAA
8QBA64MuRlDVhPYYV/1oWdMtLu+gXqhePimiq36W+9PuZ293ubNCNhxKGONxnkYb
G6B7LMOK+17HSLcsfyV/PV064Ntsbl/maRmcsNCgxc0mEKeNx+OKwPGdRrq5CE1S
c2BCa8OV7IQa7gYCn5pTMX8HL780nGHa4PYNTfEPnPDGK9ro/lIG++bX5EDtglZs
FQQJ46KqY8UD3UbgXUUV5HX/r/PqNNt/B3jDldLijG/prxnAQwgv7oIjFq4r0iTK
w56vaZvZS3Zox18HzZvwS9G5cIQt6ssPNLzg4daEPrJNIP3Oa3i1HfVYq72jbEWK
HIZ0YS8BXbNO4HZEB1lzeDMHZqxegjKk3PlFiy+G2cPm0LyA1VuNvMImPDIIzh9G
dp3KYbpEaerGTQf/l553urlRY5nnZ4OFgPBeUOa6QirVlaRxdl8k0yYQtRgTJh/3
kuTS7/TKMJVWfbNszN0hJbQqrFXQAKyY3PJW85cRxHKOiiGn8V32V4pnWKSnossO
22zZsX6LD7RTuoIbRRmVDW1qyJy8BmxW1Wohd3PKkd3asOH4XA3+zwNxidvMrgdQ
k/6xquQFyxXqPrxgHjoK2FSKh4ZAyFhlEaNDXLM6qr0m9S6G0+s4woouifhiKZKX
dQnWFW1e5Z/p/36pT0Ry4JjsENfAuA2tuILG6572CRn4dSsDa+RbmE588L7fgedX
eqvsk+Gfjgp9/gTv3go9JHoc4rcrAw3i4c/CsYx7dFqDJanAgfKm1I/j8Pao2iMS
xezDqKsSc/8NUb0gFOLZVO82C4co29tQvWM7BfazBfhpmdRP10/iaGAXREVX2gVH
rd15DmYVUZ6EdXf1vaPv1Bs3QFjBo1JFVnOfbQ7dmphJTKW9avfTv3YdIAZ1K+Dl
uBqdFkdpEFwLuRupyuoDtNcpGDmKIroFs3avTivDi/xmRsa8L2NewTtBez+YMjuM
B7cB4UJpPN35xZsPOZ6WLUtLZJ2Y1pNJx9shzmauud5pQ7kUJC3YLNmi54GHfvHY
hdNVTAQstgvja23t/Fa84XBYTmuBZ61/w6gYzFtMe0vR6Y/+20M9fPm2oVcwdvGj
tzFCnhduZEklOUhCyZ58+TCvIrv5TnM89WkpO5J6l98kaT3+TDzvfXZ1JF0uyonA
bixMaI6Y0CnAMEhBZQLwR6LewqYgWWccxIKaZrln440/W+jqWuC16YyJPJNMN1yg
CgXVCckdE+7jX7/ApZ/hnaIcd9sHsH7ofyxfvui4g8azuxjbo8tWcsmRoCRVGdXb
/DhUeG5aRAMAd/FJinH1/xF3AICxUJV5AMjbdmmSV8TEygRxpaydpX4GsrXfqLec
c7sT8eUhc5tE4G2TYgtXJaxwZP624URwBlzSGKX+0YT6R8b3GUdUphtSqYlRTmeC
/EZhRcogLoUJ1HFxQPHiFpHnKseNU4aFaDkXVGTyH6f4OtMO8MkeCQarL7o6EA94
SoVRMASgGcP05uKjA1pnKQGgxLAmttWlIpowa6lizbqvYSRbQtCNc81kKeyqve2Y
yKkaz0mffcsUILCyCCkG/fIgeU05H8sVL5PJjTbqjfXppnkU72cHJkJS5g0H1R0I
S11pfNcfTTVqopSwG4DefTc1CjE6jkksJRLDzClE8pC53NwSTLtq6kswZKMxK6vT
WFuxU0qQcE211qcCnrCupGxohvw1K+XAm1ACYAIlURGkOPfHvnAn+AzqKI90qfxl
mIPlwspgNvLczm2jCQilW6OdgXkCwmleuogf1QjhK+bjgR8hfEAMJmQy6qexXmAw
QR/6Q3HJVKIJGFGo+oWk6S/T0PXCjdlJAcWke/RmOb5zyHJqEgwhj7TJuuq9ClhC
dnKTEWc+eTW1qAfODGPlWXSNnymG69u76451G7zXnVfFyDkVcdDDqaONvNtIAJUH
ncs95puI5ZpsRKFut84dNrwRaDhf6omVtir6i+HO4seG0F+CMMgmJdxdEE7o12vF
DlI3gPOZXs1b7z/r5PQhMtzQHjPc4IQ/WHs3US7kr/1sZy5/z+lfErV4Ap4nltNg
8s+y2l8yi30E1ckWONZ09/CsD7jwiOvf4DSuHRuzwHnakfrCvFiQJkW1WVBhFnyR
de3vw1HmorFdZUVPK7R03jI1XD+Nsv4OO9QD836U93L9IzJPJVmDXmHBmFp0wgQ8
UU9clbh1NCUfYvWT78yn/5o4G5Slj+Slsw6vCUYbdU5UGUVIG0uc5ZaCXD1efD5V
mnHftYkwmhnHFgtDhuI11V3lcagaC0qs6nbs7sqm9553kr3fPFdb9mvFzjTzu676
BlhcUAkfz583ZfVrLvKLgJcbA/VJ6W5GbLS1G4wNAA9MNoh+lTaQJ2UwZus9Pv4q
/QKAGvPgSvk0QQHn1sSA+yC+IBUpV2Q2I4mG6RJua/UD9QY95eLzPWAoYkuC62ml
F6/lonOuwAoXoh3hNg5WRqlZIFPjCaut2RXAl7xR7kAbdUZ5/WIRIJU3cz95kfY5
3njjxx80CCE8AhzpibGJnW6/nxuJN2ymaNWDfCHMNj6gPj9rbGRmnnc8bLG/f/W6
H5o2B7Xx69wnqjY4CazEioIGMF0le5sIEM7F+v7N7mh2MLNGRN9Fzvh5Q9woUbYa
0KNSDeyxDHkXb6Pk/qkNT2UyCTZExxYCggotQ8rJ+eegL62y35OgGS6C0Tp4uAI5
k+RKhdSq8Ggx9G3Y0USYwi+pZCRKI+UdqS/2H3U4NJZ3yZBC77fQDgCnSPP4yttD
GvD6p4celgN8cL8ldZbxLTVm2LDfTYEwAb1HeDeGIYBoeKQp7DU5ZZ5etXdK0IXR
c7PZoBqBDd0p77XfWE7r6tftdUXV63YdNCfs/T5/qAPsElhlqBbQAhNks3nR8EWm
A1Gco9/wtRRVQQMyIA7klg05Edx/9NsnGyck9/qDvivuUaN40wy43gOlmkbqzPI0
I105X7tLQPgo+coIZhUYY4NhxkFSxFSuOxIhjoYxPH71AIjkqcdD1jhiuRN/2POO
EKWjMKweZyo1FyOyavFgjozBzhsJ0ML+N7sF31ijGzKeDl/v8fJJ9Hpk3EhViF2m
dnZ2BOi8rjR38Db2MtSXVWvFWkXvETelcBOgVV/F/j5RaKJTPjkcbyFVFqPK3yQC
e+A3pkm305Jf2p4nJ/cHjqHEDSF3/AlRACygowusZ3o15UhkuZCxayOSPD941PEp
a0ORkx4wcuLi5qu5opjGKcRMJuo5ONsMG24wYorsVOOnxUEAEHayYZCXa4JJxTtw
tCk8qvSB4CjmQ1hEl6N1zXqdEM32Hds9H4VPHSX8WgGctRcV6PVc/ddusDmEJvjM
0ff/6gq+EMr/gSpawHRfGPtHdmf2+b1Ci/FqRR30yHDwBvFpZq6FWJrOLeeMjLLA
2QK93g56obSX0uPi0tpDPgVkIcETbxD1iS/WoD/DceWGmRqkIGAsvkZZgGpLrqSP
v18xJrU9DUGPEo9WFyHfTpkCGHR+0h5mvwxlggJu/uGaxSlQ2mOY8e3ZvMCqgoO0
MhJClnzpf1DvtjQ3clWNmnKuwekG+Gws2P/hyO7Bf+LwI62xpRNtrjTRU5inSdee
/LvpitNQU1T+hgi0d4p7njXX8GicLN4UkUCbFwMRREaahL99HNdLEvgENdGNuI2f
JgIM7+4nmQ1GunETEyIijlLTYWlN9vBXqlIpJkJ7XveREvd/nV2davipbYacH0B+
WX/gI14RBWFum3TtZVYD/TyCTmw+XqAH7j6ldCBytcEfdLJhCcimszx3/llxQg7N
SOoEkbYQxmFbRf38YYYdO/8jYDDrShDbNQEhkWFYTJi+uHWWHmz/g+HvaMMTmrX0
q80UxdBK2vIJiXE0LOJbM9XdJX74TbJXxDz1CkR9oi1GqwnRZj3A30plCnbN8+x3
Yh/1B+y3VWofRMS3ypCmUK6wbwkKgVYJ0vuSa8S9v3qt6Z57JU6FEDr5PgaZLdmE
jDfvTrJSpz9qWGe6MTToQDzCYsVrunElVLuDBkjwJ224D6WgEhGn/pWyJo0CzE6w
KNxhoBAbGM/jqJT8QRI4lz8Wcvz44H6PsxHJu8tpM1f8zeYgYCu+eJZY4LW3zWFf
bLe84qggzspJ4prHmouB4keUu/HSRtb/xlBdKS3lXhJ3yh8fJAWBwMZRUWFbClqz
+hzHdaJP+0ChLkK3FX9XAyqggd65mVJFjziduMKCkUVgUNJrgjWaX5N2rdzPP4Sc
kLOaGta5uBcBIoYbc8Ft/VoUb73As0lmDbWbqJMVR6CVXRoGsHSU/84bAh6qNisA
cVsFNo30FS17Pj5xQN8yJ91N3htdxWKTpHA+FIaon7kf8+Vl7WKD1r3mAcZZX4TO
yDqO/ung49nZ9YF7mP4PnUHpviUMJW41nWSy5Da5ANysPIY3SVwVHlCJG4cebJdX
azCPXMznMeU5ESHg7S4gXUwksfxdVeaXSQfcXVTHCbRIvpBerIuyuzEnXS2nC8u1
hym2PDRvQgr6IQSyJYewlo2aOooUubtiHleSZpS3+7HxZhgR5BDQk2JTxCzPHINV
8vFNBry18pORzHHxxK6VywdNybNLsixK7Kln702YpikE2B4tMkTZzKhNLUgW7MoN
ZdscFYXgruAt+BS5VpBcLNXCQHRkQa20x8c+T+zGVxOXqZnPz4JoRvu7BVGP/JfK
O4+OUq6H7/gqinh6pcoy0y+ESMfTW3tWr/rXo0+bU6jabv1hF+V9pTssktc/7AQw
fYSTn6ZXXT0/T6Pwc3QA6Nsumm3pxpyhu33HIuD3RMIxJ7cv5jq5NCHl7+4m0sns
y4kcrFtZKrLiS62KhWHCc3IW2ufivCy+mrXkLJydIB031Hy5lJo9jE3NELKlNEun
YhnGsYlceqk94hIJ0rUk4jjKO7/wmTq3JvnY//n8BJ6LlulkiEpZ5DKvPAI6KHax
usqE15vqQ45/JKdiHlPLe/UOaW/bRsab98XUoXU8yWpjq5sPWtH431L990xTiFdn
GHc6yHq5H8/XM/KgzjPpEHiruR10Jph3CTEbnEnMCi5ThWkrI/d9TKNJfV6SU4pk
BYzqYPTGSvuZcmAlLWkTMDU2WueV+JvxG/wVYl14xvZlGXjhb8laoPAxfq0f4N8H
oZiBolgX+yBwqFT/DIt9aUPWn/8zkiAIV/ivMptD6EqTvrtSNRyWEj1CekOtMiUy
oUJsSIV/OpZz60dTn+MZxnylpdqLDxYNQJLnUxp0qnjFZ+4Bgz2szkHPQlRDybpH
AlALH/V6TwFVpsrh6Wi/pfQ4BgKBndyZezCliGpls+xDSJBofQrc/pmy330TpelY
few6XGWbc0Z1DUA3uSaBi83cznTRGZ0SMydxu1N5k57In0y87Myj4+O7vBZkU31h
OG6rdXvJeWk353PFZItJ3tGg54haxDwfOoJyypNFCwqMVjKrud/xVhDdZgw4kWmQ
YR9OTS1n6ZBMeqKqk2bMVQYtMpE4QiwsfQUXwXYkS9GA+GCFeuWPe83Mk2srxxup
CiZNmkZCn1n82LkSfgHjt8e3pKmelC6EiEe2zeAd1OLS3542yXy/XmMztcBh9WSP
8GlPYYyYhVkMl/RyyQmmRLvTYMd0cMRdrmnMPM6dcalaq+ndVmoIz6OtPNaPY+Ms
R2T5Le3D4udSkt0Izub18SVsW4xeuRdbnTgunGEmoQ9yCX3YT44jC+Qcvwhts708
xxe1LVTfx+i1OFntkk0LoF+pbsrrqYgfSF1anSh8syi9mGXuR2DIdJUCvUbijpCi
LbQ8dvIAK8OPbeiKOr/3vmJ/N6O3Wlci1hZs7oszQH/y4GSTe05m/44YOgwX4xGF
b3tARjTgv2ebXXLEAqtTDPxDIxxPu4en+yYFaSwsbOjpaSILC5F3UQ1H/oyb4NzP
8KkW//ynbin95GF8OHVoCiCD1rDfBXtkhbNYrD7CiYXQDAUAb09KS5Gyt3B2PvQP
BkFcpbeQcWxRh+wTXhLBwHV0k7PCjVQ1y2uqQUsTpSrtCtEDabexOl+fXm4fGehS
WUEmH+i857CrLB85NsAhhCqpT+ZPn6LDIP+q5l5tLkJWzZZF42hZMKIfHSbCY9eB
bEo0PxJo9H9gOT3fTJ1kuEC18ez2Od9COjwZcq6UvhAiOO0vTtByq8HlX/SXQkBQ
ZeU230tTiPVz7yfyF5zsLznprGt1EM2ESnIJ7XrCDrKdrrGZT5lbYED8/KB6JZkf
0ZwvHit5T6HYE+o/8tsAFDtFD8wulscRF7UMhNAPEQK9KQS3BS3gRpWmryYbA8eQ
PH3s/jNbPw5COwqkAZjZctmIvdhSJxZeTmxJlkQyarKpeEboJHEgSrt+hvtvuZab
msh68iWP+grMkr0SuXv+VKesZ3/ly0p4NUHhI6/3YeC+TfuielSfcE4ochEXFfJh
yAdBbA65bEMxfVL2NcLO30P66PJbZFftY+ckOzJJYEEYLWxTJaVYaJCcuKtYKaKy
cJ3p2PqHZOyYTy6ae12YX1xfH3yw7B8kA+VXJkOi0uk+FSzmbF1qqOtAupmc2TyC
89kl0L6V9WPfrLMdZUXPEZ7Siu+p1diGgVdkSBR1Sarx+7SgDMeI+Ko4764JvyXk
OU1F6B2XfewgL2zTB1cVv0CPnOIqPVcMvMylL0lyR9urf7SGXcfwysIaJLqH13sp
k3wdLnUXLh15RYwFIg8r4ECHQKzkwt1C8Kex5JPa1KwIIkeFJrxY4LOrITNmeqoS
FpnCiiFGXVXUZf6btBT3qv8PpkeQhFxmDH4qIij3o2xk5H14t+fVeYOcFqTEMBLE
uAMfwi0XmgGzhDeuA0vX1NztgR/jL4phIEWwFlSQd3GjRREV9xvjL9u/nZUe3nuQ
KI0vRfwO9+xatFrXvGX/AeEUMA+yZh8pEVbtmMi0wW6EH44ReOkYbo4cJbd1Ri4x
wCcJ43Vc7mmgBmZ+LzdV27UhG70P+Va1A1gFRvaJUvCtUwOrBNFuDTEz/l0HTLXv
jHrhphemSBt6qZq0q8beuAoMWVXoNwodM5BMw3JmyxxPvhcXPsI2qN/4J5vo4e77
Fih1Ry2JP1AfF3J7ZfZ8pTzKV4qyoqSfymGdf4H6XRYynVZ4ROOmXPujg+4XnlIZ
KCiPZ3ilLPOELHROdzIlmyyKvI6xreCmKXd3664w1GGuEGkHB3OJ0sx94gC8ch1q
OHlKCRJz+VSZtXa204hQLxugSnwOPJkQslEEsFrkneN4GcSbfC2tlnlvNjxDc4p6
XbZ0e7FU2MrpMQ56paaKFNL2tTIYOAZh2Wsv63/mAC6fwHZ1EqnK4Hq+/H9xxSFi
6Tyayy/74B5syQPCH6XnnaOVHvS8dsSKkEJgeB4C0cNXN2uH7d+h54TVbG7m7rey
9c8hMKKaNXDFDP8GEHTTajj55JNyrKEYI6ovXkyKIO4COVTu05nw/st9uSQPfu7M
WRWn4rHUxjoNChbMEtdLzXMQ3T0v7RVtPyDMuCrNT9aXV7t9KpZFx1up9FEuEDdS
AAFM4g8Wn3Vsgpiq6WTnNkVH3jkqmnX27m27EXM5xwMRPowMeOqdF8gwGBwFzkxa
LAlFaunv8WTSsNLgPWX91x+s9gySJLu+Iv64hEQdv7FK8H3zi3Eix1Pa+lAThHGu
xUq2DoErXNrHueW51D33qBg0Nf9p5row829qVSPXf4heQ4sdpn2pXvxFQwxgwe3+
glHb0nXFpk4rgeM4w0yZKtQ0gWQqGWMCosObIWbV6j73LvSnuYKbg20ZYYEON11K
ga8/nHKqBMdo6Rpiy8+lacmr/M4mGChi+W1h0w+AQeY1VPl39BYG78fhzjbv3MEn
sY4rm8nYBaboU9g+PCURBnmLna22QHkI9FduEMJ/JK0KyLXHEEU1HyaLWhL956Z2
RiBHS8LkWngc9eOKtuAFMfht20lvXacUXYgXtRcSzrwFSZToO71tq7lCLH383hGv
RUQe8MfZpU6ebQ1LlqKj5AgSyhRARFhO9PNBX5YyYwhHHJkbYLkT8tUKrCauhmyD
dnEfFmLikzVH34sQyOB3DsYeKLaR0pegrm9hUXsfA8593XhpZEXDTskXtgByWea2
Ro7/effRyiWGGPWoynP/rDmJPN8lNjRB0PK5Hlj4FOyqBxglqZ1dSeDvXjJKqHKi
+a0t0AXMrISM7Vf79oOELLXlY42XcO9ufF5A8iS3B/iYVCe+bE5Vt16+wp5or4wm
KrIFsjNbV5wzCjOrUUJCHPQnntnQiQiR/2rFxymLw4sa2ZySvGbTwrctYasvJ3BV
kBqSFrf70DizoGLBECMuWkItAeECtviLEQxrtwEweytPEPAlYHZG25QGULhkBL25
s7F0MK8k3ZZgeHIpl5Kb/M+TOUpPSC+9/UJ59q8sWsszzhOoe75S89cmfjm1RIG3
2zQM0Vt2DeC7JurMqi01VKDRTSMwjUijrX4KeSqyWtnBKEIRz94DkIMev4Sg6URV
wPucl51mx2cMiFTyKHYqQuwxh1VSZBMjnkWnNNr/haQesTzhoLEynYUjkUYcBR55
OBMdEGgSozNcyyCN1W3nI0dVCHzRz8fCCzAU8F9TWjR4N7ejxLmVsmJEv6/bB397
e9OgxM/6P8I9gFWjIVc/TE0Q+cD9fuCVjBeRR31rvQhHriG5KVau3skfxfwtFXGv
TmtxO/SQR1OSOIvqq7No8PPEPw6GDISHPPK+jfZ91IYVbkJtCugyeZOwO6SkdnSz
Iuj+x+I1lOaSqgvT83gR/A/kI2TWkQtpJvAA4Y50VarFIpJnqgbHDQmxBKcJ7u5/
w1qerFYNCohHfRdXgS5Kmmx3zNUFA1mcdONlsPxc5pTkPQHdm2MC8Bpvf1BpGMrq
Wd1LcncwsN6/nzDEVc8YwZe95MBHWnd3ZRMHWum5DdiXfwitKhH4m7GJCfsPD7mw
/DoefR/QhQys9ks5ot7jaAUXLl/gShnZVOP9AaE7Nl+cJ3kCuaE7Rxs9Z1l0a5cd
vvW70yBTZQMbTCeczR7tmvry9yzhHNyExgQelNZhYRhAADp+KeLGTgVg+te40RmN
GQWfQOAh7h+aLMubTL2+6+IHb8cpvE+NraBQAQxKfQx8acly8K6ECV2qDUv6aqTo
M69WXwyTJIQiv6x0ZRBJdSnCmC4ZBn8+/dPwCPntuDCY43TzvdvtLYuSSsBiBlgE
aX//BL6Hi8q1HKtksMCc3FOGBAeATZfIiTJHakYCTVecnjPPJjLMgSBBZkQ4SRTL
3pWOTEZZQUriqu/qq3B5S0iCUIh2OSbqtGXABooijR8bZT0upb4ZLDNjBBArOLWa
fp1AqcMbT4xQCd30S2bcmr0AV63ZpjTrNjBbo7KjeWdXME06BWDkV4XizNIsDakb
3Kf1obii351m3P2Hc5CgA8U348YArxMoDV/qe94roCLPKbDK58kyiSAzbHk4DT/I
u9taQlfFzCYB5jWhN/dsRPqFdK6gH8ej77SV7v8B2pqo3k/1W/NwFTySKo0PnBkz
o2+txABw85UBzFzKZntMWNjF0vi69kFSDkFmqtPtJO4uQAQQNFMZvJLhCWxsA+Ht
1jYCZb9Iz92JqXUMnuDlKYf64T1Q0ZGrW8XCOhP2CyLGxsNvTJS5Ae/cIw9l9HT2
Pu5ZMTfTGdMVKAsa62p9XU89sED01ks3FbOdbokXHliLMuB5wqu50olzw/uEzu83
IWznl+0NiwQAmZSCxY6Q0fub89zZOL6vqbQycjgg/gfBGXHub01/TSZgZ4PEPCGE
RfKwDIeq9mWqM9oAj7Z1dUNLv+7lk5pH8+FJKlLmbTY93BOeYiKMGA0dm1X+mPnY
a+bT8RTdCROuzBMHDwPEzAMnYXJ16d3jEdho3b2lj1BNSD1Y86bbO31PRK5TvxtP
XGIVxXLJFuTVb6okEMUDgxZBAd70TNquVklCzfIBltquplylPLNmd0PW/rOSI0jD
4BOA33cJ4+i2a10bsYVNdpAu5J5DhFx8RIsHI8+EpQioaLHHf1vNWt4avcsOvplA
Koo/GTIifEm5583se2K1PGqPiElaJIqMtg06mnr1bTi3JhRuojWmLPWWOofj+H6S
m1LN9E9i3Qt5DC4cCxsv2agygNQEy7uFUWw5j/cOKV8RdcBilrKyFwusISmWo2y/
IMEqWp9LCKrsf6sD+BMVeaD/z3b7KZGO/ge178ihdodq5ts9n3ipKdGJXhzeO1gp
R8a0nBRtcbVs2aDEoN6Hebyc8To0qTgkRjcj9QBw5i9E52nJuL/QoHhB/05hZj0H
Ae9CvuYohNZYPlr2a+68y3Oj4CRWaOO85ROyRNXClk4wG8YLrWnOTpeQh5z3GzMZ
8flCkeS6SS/FfANmxCjqxmCCNWTong6exth4hKeNzHUcFhA0LlvRSrM3BVieBMpC
TJSmxy0Z6455k6gBlumLLBtMZixmgh2c1WgaW3ONaG4V0MNBcH4RrZxpv/h0UxFq
6vfnENg9Xe8o4coeR+1IO+5Aac40FqmcqYmgJ0k/gkOmeGBEoTGKEdBXYdnaZ/5A
qGx7iU5P07HvUsD21VxGSz3E5dfowtcGrw7GzsPE4txnbP09KXZlCZ3c3bYhdtpY
WuxYXMztbMfeHMqMCmQykdiksp2/I8gAkKKBzgeFAIfRYcuBXmIExto6BnKHzDOJ
7ewjQ6jhiw6VDVhWyZNQygxjHDgHw/mNAlgfCy/wmbqKYK3rcCXmgQ7ZoHh0Q/o+
R9dwPYPQvgSFwlUWGYNzrsV0yXnMqinTk71a2d0aC6doUt9cSg0vb020TsaNeOpu
ZT8qmPMLnnTRJ8MkFFDMaMxRWwJ0gKj0hfjs5QVykM4rPXdc1K/5USW8basVb/oN
WZRh4Ec5oQtXrUdz6ex6puIXUgmV7lgKD+1q0SqNEg35Z5z/Q7KkmmDhUW4GVUXY
79SrV9lvq0jszurVu8YKqjGAVZ6rDON7WN6LruG38AVgiEOfl18bBG3MTVtdoOcj
xfDUrTdBYNXe32puZT8mVhTbSJlfbeAg36dadikoPaedFJOU5Pwgg25CrNRWj/ng
slnowlcZoh4SuVfJ+a80A1+ewPQ5Cy70meLbP0Uz5W9VzTLUK8NG/i8HOgodc3TD
7JBWcS8t9r3pzCxe86Rjqqx7vqBSGJKN6u/mkYGdN1tWlKFZst1r6/wZx32XFu1p
WKLBgPGQTJt4eeMZ8uoArL6zLxo+OEFhqjwMexGDbKhJXkYXcbjEDIcSiewMtGOC
HJ00Wp7VrwqJ1x8ylmlMIM3Pjjrs1WPZIuuz60KN1t7MPOdweqZdOOMfphoIpYqb
taXHl+X3CjZq/hjpOPFrmO4CTFTLJoz0cIUW2TB/3NeCoEfU/gdGwAAhf1/dMKBz
yY/JeQboJjxuiToxq26L120qCE8G/pXJbuQq7DKLOIfYtlJwiMXPa1uCRu1MsOwH
TQJXKKMKk27o1jQBNOkWZncUw5R5j2yiKtXku5lgEjtUO14WHEYb7Y9F/CArgazs
vmTF7S4HGrm4KLa5xjel8C2FLZMCbMFY+Ef5kPr6J92aAH4lxbcPoT9QwrOYqlQr
TGeNy7LezaDU0K9goSWr2hdj1WzYCDtFgb1pqc4BQnjmgWNERWE9Y32iq/P939LF
YnqKU2a+5cdeQWqgGAg9kVzK6kUaOSUYM+Y+gZvajAHa/EDLLktP0iuyZBMox/Ne
cAoJvVDBVO55YtjxlZfQOJ0XLb4LCSxJzlSDvyzJyEb2brA5BIe+6WmM5nkz2rWe
EGsoVeKro01gbYNNwC2KxfdJladBBVLejQeC0Qt1s9UU/A20Svl/RhiXeCLI4GKO
ZUzq3CkWOy8WeA9uJ/O2Nckdz8RFj4XB3p9J5uA51WKYZ6WBeHPTRT6llgkS7rm7
lHvXjKWB/jrLLQ2E5gpnztiXGSfIPrOmp0CuEbzyv34W55YQlE6Vbv94TYUW+pmn
HVi3qz3aoB+hqI3nfa8hjzXm7kheZusnEvOjr1g2Kp6ZHZb5zqfF6u19b6S41kXZ
usXbBAI5M1q04uCjVKoDNE0MQSyn0HjkGUvZ4hPce4yGWnvKM478d2gIqph1X+eb
Oc+ayDibGeE6x0WuZBWefvKfiLTYWCME4HIRf1nM17Ufd08CKoFsUp2F8U38yLmV
C6nmW1miGlWwXDo0u9ouEz+mWDD/RcLtIpUgb1HMNot8qRUF3NfszsBZ8dzJxgtj
uWSUUmVp89VcnblwTj72MY7m21ZbFMvuFXJYvGVxLXLUpB3MRpetb3iZb/FnTFa6
+NPNb5gb/SVp0W1+vChUHFSj+J2e1UaOnDTwrjrcEXSW1HBxpx8OWBoAYE+/9uim
rVnaTcd5ech0DuLjqwc2pkVFpv2tPaAFc7rj+8f463btBjJFpw2xtmSoFP6ZSAaX
+Y+1GrXmMErt3DFD0p71aqu8fTQO5VeQJ0h4cN3iNRDHGgs/we21YptlIGcHP1/F
R20t0k6UdjQ0HyzDLyZpThE2eEvsTlM5ekhiCGAGYYP+W9CeYKaUdBXBeFxLEcmj
O7shpQacZ0c6fBH5Z/YKoN1d7TcapnNftWbI+2ZtSDhSJr/R8WUqBeKBlr167Jfc
p8gS1Odgtt+pXZMvf1yFqcWgJjHw2YR2xEzxSv7pqfRsEPDjKiS1K5KmaeG0PW8u
zzo1mIFWeWUocUHstMAt/1r4gC/cH6Q1n63KpUMwdrLeRySd2RfMbr3ERmWgBMSE
5PpRCslIy3d1dxz2AIwmOBizqwGD0kEVfxNRtc5cp/aK/UysQM0KpVTZKAYb+xPT
SMkgXuqwCLAEZ/YjkCpR/WX5R8u/pr1mL8mgM5nsE0QyZOMh1NwpLDit7gWL4xam
xek3+S4qnAuuZ1MIiM2py+mZgyzhBodY3Dfb3O9OfsZqPfAEm/75byMXCTP4QzYw
atIlapwYlVrIUCGqgau3+DetgtiCimwvovrgY0J22tEOXmxTvmu3T/gphJ5BGDoU
ahOYfQp7gQZc1VibrkL4UBJ8vBNKrxhUYiG3TPO2HXtxbSaxmiJPG5gunG+qwqk0
G7JCKYCfj7mw0iHHrgsK6oIeKvHMqEZIyGEn+Pi/Llg6VbthNIAZWQijh1kuqTac
ymGg6pjhj1wACGuF7ZYIDMb5TeoouXrYB9nqrzqs/3fwEsDtvGPtnRayQpkTqinU
czUbYoAppswKlRbwyGZGiVQeN2G9v84xthHnkVTyJFsgWWQ+TjkbHX7Zf1DTOq+N
mUskUXAbCNwhe+0nBpO8D9SREZNpHeNvIEwAvj8RHJLwCqczOTw1jNGjIuwARiJj
nRgQeODiRYzSpPYdVA4O/5+Dyy71FdV4gZ3fZ6mP9UO76AZVfqpdtZ5zPFlyQpV1
47CrywaxLFvyCYNPp+Ap93sTN24EpzO8R23JHC6LYWrc1mMimBY1Y+NnayTqCNdY
1tldaHYM3gA9+SEcE6oX7wXlV1HBd8SJqZZEISjCTSqPScwT5417g2U9upze55Ye
QFfApbxyzJ98Qlhvrkt+TezWMqMUm83dtV6C5GjIWb1GVUU47/tUKrmCsVhvMNbb
mNGoLGgtbqBoQdncVGbsh3hFb6OyhyV7P02+ehjk7zOdRWuXx+IfzDfYEF5ypEux
tKpjnjZn/At+Uq09HsQacYioinpACoLjqDRNYAMCA3crOaZCLgTGtZFeJxwl4sVW
oTbGJ8KKHakj4vWQDnxK9j8EmEpxIESQrh1PkAx8Bkk4B84T2ZOXd9AsPyfBOeBw
7f8V6kal26ypWHRTwoMb3IHZkRl1IBuJ8VbLpe7TzUeyLSDIxH7iaaY2wBjuylNC
q6xNd7QoHbA8ceVTRN1TaJk5MdH7EsS+sQjA0D1fIDV+9kLCbKCXawipG6wiISkN
br+PAjRvM4ap6WG3B4nKmGQadXUI1vv4HIE2e6JelW6GHKRcysZVIhSe4P5wRFtA
iLuuCVF4O73G4fxRtLaQ/v3JHiflQDBPpjaS9iBcIAPZSVnumA4VXrTTZKtKNGXa
s8uSSYC8MO2Cg2xo/Kle3wOwOh0Iwhy7zH8GWUFZVxxkmpElkbau1/Ub69VJyuma
AExet11HisWJH4AoHrCBK5vS3A+HTbKO9dhY4p6EvxBTsaOKC6Wc8iVuoOdvXNzF
2Esr+IgftdJilaBv51JPgP0J+xjGj/7Ie6Xhx3/BJ973DXmEGcYt8kiQrS5ZYN9V
Tu7mTSlXGH/Y4ShL03VjlyiECIhY8oDGGfQOINLjT7/sQ3cZfYpZTffRo0ZrBdtZ
CTCIzC+H+O0Zkm6JOQftRC7SfgNNyz1MnMl0hrxEVsLH3DEatGgWuWFimff6YPsn
tK7C5IfHFKUYYror7QCA+Z/P5ROoW6ebUVbtBEjReWTyQSao0ofnQrpQnnHeAzPF
LiP6/zbyFE9lAF3i8HPcMgHJ09YpSA4mGK9NnPLaxOrQprMfpOubtSJYvdubVpN3
np+rxFnrA8fGnxAtV9Ro2ky6j8YZG5zILZYY7whL5N519y9Td7ERc8tsu04AM5Uz
opxJt45X40x+KyOCwj5EzeU9d3XPfGUJ5iJ67TzAtdZIPONgbbTTb7FRxAfzw+6V
92xB/XKoWXZzuVBJJTIIp88C8HOKfdBQgJE+hke9jXCVGNtzTOzF+2cwilg1NY/B
KXpkOr7SDuuEefekDni38ja1cuWtE7nrme01Xzh4GxzBk7OaO8hQqmDTPz7y19B5
W7xPepAGl0lN0oLEaHlTEbwiHN9a9mRFFD/lsfahHVn+Sq3NM08OV0h/l1g5g5AM
LAOgmjuX7eEcryLqZgHS6nRQAzXwgsmPWvEBiTO0bf67cQckr1MZyN5QYGOJSLIK
o3jNR4ZNP2t1eYFz9McAB3hxlrQHkijLBfqoW4H9TGy4pAcIfyFlD833hwrNpzl0
95CWx5/3HDezeUYOR4QyjtfTiMTgRYXap7EORzJhKHHIL1Wd0D29OyPWoavyn8Tv
rNY2s+Mr5KGtBdy7notSJkUIvWRrW3zh06ACjhnu5T2wdbONVv9r7KktVpbPEndP
1CR30rk+YQOjPJwKeQMzBCERTgIOdkH7uRvGaQ6R5hKmArlnh0kzORWyOpcJ4cKm
CmGttOvn5jLV8UP5RZmnndXk6MCgAN3/HFZNNvg7epLPZxLlKiuc/sulLp3l0eNI
jTRASgu4bmCtFbrH82qQfYOHNPowTmohCUk1SpT1KPVFjp+CJZOA7EwuPSUxVljI
FMLTjixixvClkmHuvSyKSFkNpotDBMx+3id2/EgoVKSV+5GfUVhG+EIuWfTfI1LW
ZNXbU2d1yifXDJgBUo4gqAkqoBi6A8+q63/WwkkR1IEUlj9lqlA63aeduh3H42U5
cSPh7gdzNnEz3JOLQ1FbfxBWu8ENpEAbXdWWzJyo+S9/GX2Wp+AJZJ85IvA6Hxcz
K96BFWtt/TgOffKnEi8Hj+7W3v3i588ecGYM8aCsUPz4BXQIH+xAtc6KP8fQqeHo
llKltpFEEStJbSeW617zcgxQhZ9AgYsWZ9WKoAhy47P4FB1cn1xZBTr4PW+SWtOf
fnGi/3lopWRtTvu5VX5ByCdTJBfQQOwWGegf+HpSoO+zbPKktaG1C9Uzbky8GODP
sXzlAWM/TNjbRGcmb2IFQQaDtmzhNuNYjxCq6+Mvj30TPVqTF6JOutSD6Yf3Jsse
qeMmUqZUNOpxQ++x8m3cPeFDSpI5PJwZkIXrpyIztfxpisHDLqTtbSpPEwxUdwuy
Y9Lrl4ytT9B2ojVf160gAbqoxOx/6C2ucDHu8gBJSSCzlZAAZr53rbuQ4mXGGzp0
g34m2OETsQqw8JWec8mzEnEjnpTz4f9zuGmi9cHxaa/Jyc9WpShCTROuzwCCmLFf
yVPZ2dtmQ+zoZagOvBhE42H6XwC70GmV2F3WxjocMty/7wsOlm2obPHZieu1FfQq
BEuBsQTbMF0tYiNaPG+FJaZsSCXcW2YArzJHXTXeIf/a5q76fetthxUUSqfq7XdJ
Bb8n4OKxI/E8Bg1Fk0WB6M/sGmhcJpVcUWbwbn12cY4o1hF3bpaMjGFtoD3X+eNq
FNivTRxUpXn0Pg06QfLrF95+qfw//0zy6dJzOR/1YVTkGjpeOCTGoDU90yhFzrNV
kvaHFm+wfrR/GI2SXcdF9T/LR2v3/j+x68EVx/XY67YBbHji0RMiQaSkNzBBXzDd
m9oL/g0MYvGJB5wU9EMqVFeVUuY4HKe0UeNJCaJ516EfvrQ6XWY4kSg4AGxsSnwy
3iqiOzH8YsutPiNmucAVOXaOyJAlesjagilbHZ+AEduKMXAbcjgXS4gkDZZe9ubM
QDCiF0cZS+JFMS42V00ULViXy1GVXdbObgODWL5cFN9PEwjKO1K/3zeEm/mmIIe/
ujqp7CBEYg3bed6vKYc0mWkRPY562hsIsnaCWh6lgDNphaUA7u3hXhmj0LtamZaQ
uS1yQXyb7sGVdhbRkO17QfSEewNfpqxG4Omc2cI1qzgHKA4i7r4BTbhRyGB+f27J
bP+CbzuKUKAJLXT4qxrVfarF4kRLlgR8gblgrUgyh88pAFHDJJgAERAJDxfYFe9M
/i1GHbdlkMxhMJxaP3CKG08BoAIQgPVTJbzxZtnNjhjjZk8f+7Dw2d/JS0sDMHqO
VRRuGIAazWj72KIcafkNrSadYJRYwKdqhsKzO7xkLnNx75z4umtTfXAt9D5Y6Fl+
v3yx0PBIR8vImOaYXebzN3SvyZi/d4TmV6xercSWbQxxENh1BuQhgnU/N2jazFvP
qo9LXWFxi3/ahgZ9vmkQP6yNcStUE9sRAzKwwblhepmju+XRLrSVdBk0rJtA7yvD
/jt0VBS4lL7cq8v9XL1XT+VIZTdAOzUOYPF8gmK944oOgRZGC0P+DC/z8R8G3vja
ucjNuMFNJPFnzw4x+T655ePu6Au/LxQErN93FhbPfKtW01RoLlXJRo7dRI8MIO6A
ak7jExRyptGIlzmUcSLOLEvx2zygw1qUqrJWP4ZYthi8Jv4rBiSxki5o3sTxENn1
0RhEuYpexiy8/G+YuRv1+JKIkvh1Fw0d37eYkLCCfE9Cum5kF3s6o6CIcBdTGfxP
jW/lbzVpJ+UC4dIsGEZXkNFTgWCAl4N+m+IkCrZdMiKDDTVhk1FcOCX8DaLXqVyB
XQ17dOilEhh1tUnYMFP21W3lUHF3/lMj1faDCYBgtFKhDidqPYEWqRU39FMu/0jL
wWTb6/22hQ1gJ9QCCkP7EZ/pG2odbhLE1l3CNTuoOZUeRV1ZfVf4oKfUnBQ4AGMT
Y7WKr89habQi0alY9uxiAo+f96ksAuPJHWvLvjUNoIePcaRLg7/HMFDHz6VGmoAA
LauMCUIbT0g3UVC5h2ohuNfTGmMpXWfrGU2TddQ2OAErR945r4TlOhjBMRZFlYGJ
/S/9a8HKmLe7Yp7JCpUlvKNeN2hnbZ0bKCGRSeX9lIGl6Ujr2b4obwhRwwpCtXal
oEva1IOIW9eT1+Nrejcr5xH+CcYOzrGOmHTecqRbRuf6qmAytsJTee+f9FQWrpoO
Y6Bb1W6yPrKqlk6xEfZr9btESSdhzAKZ7iXG+F0RDRyA6aYUTVOHjMmQ6T9AYdTI
Mepv7LA94ePGeOmuUWQ3mMliU2EMSZvgGm96x6lKR0O595BHEFOn5AitEtesKmm6
kJ05VxfYI9aOZe1gZEUW0KS+k6e4S/YylF6szZeqqY+4U0iK8jlkOsUZ9SgrTE2T
EsX73q/52vrqcigJtLIxOdhWAdaiyUabx9t4uLm4mvr8CwI/x6UtSVphMcn6XNiQ
uicqH5cEn5YkRmWNbmi58z3lApG8n6igHPD5Ef2NI+jH2PjExsYuI4oVUMJlw29M
vAli3zqL2sDArP4d4PVoHKbrod+87hXoqNW7xv0NII6QXRTdK0TtX3cS4n4nrYzb
e04kEOBjUU5r5OMpJEvvTeMKKzHO8G6bh7zq5vzulyyoK29iaRmUgS6jXJP06rOo
ZfgAtzh14gJ3z/yyEsRk9hWhffrvCXsnfkMUKZz+GD1wfIaImpML2ID3XtSOcbPl
kHknKE1+7gzleHEGY3nijh7QKW8WjLT7Lemv9Fu6n5RaceSH7SW2z4CImxoJ0DwQ
UtTDFnc1q2shfWhNyGXLOlB5idGdcwCjYKxKOM1CIS9Xrq4JnF+Z6MOTZJDaRvra
52RMogUcx2onugc7mvpMEiIrIX9teEpr1s/9bxM+IVhkUA7t0lefDKMR1eyOeXFG
JPvblKixDepN/J4K3syyyZn0SIAp771a8C+cpY5MtyJ7hZkTgO1yaP1iq7hwF0Jk
7YBtgwUgkGsCdKiyHQtJ6m/uTavO2Oidz36MgMCM7rxTIlljUR4UE31QoSSXu4QP
+cghRVb/uZOx+LBn5dl5hRZ7hhPP68NEVbKzNMZH4y+ms1XWiY70rvKqLFhVn49M
DVBlrfDp86HNds466SUcH/hS2DebWqaRdm8CJb/6XfCoLDIQG11TmqZdI9qEyocJ
U1B0BcHMHYFAGSNyWJa7p0X0rgxPmoqlyYFkI4OM72xQ53YuEeJ3m2DeOXyqNCtr
XpBLVN2FRPUa+yjV+vVcfJY7PG/ybj4CdL7UKuHFXLskFTcx872eKmRNUG2VFAit
ZfvnHmnuIHK1RNk10zODbwqGolBnO6CTnUw9rp6oOvBwdhq4RKvttkvH8UTPehfc
EGW8RBNC5HdbFrEXPbhumV7MDnbaMLYVDc4CyV9eWZ/OlVzZTh+R3yO9soNUHYz/
yDV2LCTR3JBR59ccYltxjFUHgSkHhlGNYC5j5Y4Kz/daXfcLw1AUSIaUDSHqTCY1
SNg22daxkeWM6mfNUhmMovsjOTqXAAVrId1ZNBcZkJAOivHU7oZOpNNQ+V7H2hUB
+lyG1V1sFxipBqZ+TTIzd1cCrxD2J0/ADnp9HS97w2zfp+h7NrUExAcIvRfQe6wt
8S0y+wYjXhxLxqruElnPxk+NMwDXtHiafE9mQzOh/UfCURZA7gLG1kbF2bBRheq0
v4/uZINXHuQJJAvUFonXZBw4MRepk295JvHyW8CU2XwS10tNVC9QS6f7zQqpfovZ
oh/3Zw9Iz1C29DyWUogTmfNP+ZpHGkqFohMtmVZjCDAN0ZmqTMr0EfNlnTOYH4BB
QBIuSl9Yfv8k5J5xva6JTllu3H+j4QsFxBwxW+i7Wzgix6wg/ME5Lqa/CSxRMvo2
lspL/yc+3zgVTTKKxFqXKoqbNf2Uc9iE4+YZIxFw8MhVzZ8eDRcKMv5Sx7rkNzVS
kS6mHFJ2fJ15dL4ngxisqx6luf3SARhqEmFlyVa/1S+G/Arufecihlm80OBXGBew
mwskND3tbXuDabGogGHKuOtJd5qw2jG2JKX7Y9Y8DkB/lKj6+sC0fem2hTowQZu2
qZKElYqUlsqltXlMIVyreTw7JEsfq8EAJcYc7UEMydkfMhxT4vUS97IntTHhYUDG
b4pBpQl1ZRUxMHVJVOD2CSCClSXbVhJrn4f/0C2ocgcSFPqqgS3LVuJCz+WLb6mK
aSn5AZyne+5S+sHT+hbdvQec7cxzQTGCfccM04pdKBdc5p0TUNyDS48iy0fTtXyQ
LnY+x+/yYqWp8ELn1VMPCrw48689t7eb1fyPzSiE5W8IcCoAoC+/6s5Ch70ZU/7L
sPXfe7J8kmyZAZ3U1lrDUxFHVTbkqcOd69sr/Z8k2FG6oCVwROU4KylcoOoh5QVP
Aju29ImU3Yn8u+9kLXZwoK89zaZGmMaIOsfsDtSE6YX6+btjMnytm1u1p8+qqdga
66mZVPYrIfIK516xw/H8MWECzdApa49+70E+GXy/fe6K155IiuEgfTtbGZVjX6FI
0SktvqxQL0GM1mrXpOk4pC7BwDdXmlhpi0WyNaYwg7kJxpJdjpi7Frk0I4KFLa8t
hPntE0JFHI9XI9H5/pt1wCN1AADXV72cpHwUKf/QOQQgTZdkGSZCx1+8gIZooh9A
UcVeKJmxGECHiJDyBRd+0/938S+TY+EZwB8j8Be27kYH659L1CPtHjE77RD0atMj
tyOpm7gynaCTaIX84ehwl7hOWVNuyx0vQPhiiMucoAsr7zRGzN12yEpS7mDhikga
y6lunFh2YHKo4gly73Tjhm8TPdWjbk3P9LfiVlLsPA9oI7gLvw6dsuhsLFRm2h24
3iiAl+A8o86qu5YlC1Jvs2j/ghsIQVXGhQbsZ5HuEGDg3Oi9fm907mQ+ODlBp5Je
mW38BiUazzWixcV7FaXiEan7Lwnaf55TDrk5smPZIWHo+Xxk38XFC67Oc4f7DaoD
YsnKrawYuFh+oBHxg9bKYoAbkuFqgE3e73eHExLUBfJ3A1moKAlw/o+EajBa4FVb
LTWrtckojOlinlh6orKSDF0ARVNtl0gxjL+JauuH0ViEeWS2ruxeL47psqmdW0GN
w8Pe2cP79kctNgO8zsCrKs6S/EfcX3jq2slr6oDZeuAkMjvzizLvmdamF3Yq/bpA
Hx8Fxi0fnmVUPEsL0mdFLmxZs0IlfXpXGj5PPxOumJSDM/7HMTYfw9fRBnuj/3ec
qPcI3DUirdzQBdCOo7rN8U963Fknwy+Yx1xB8bWVWUulql5ld4wA4I7Ni6DeADyr
d+afp+RowyuvlvDDfCkRAfzD5LF7Xz8lw5m99xkiyzwvkAXcApd3NztFR4wW1Hne
O3doHY/aXjUmPxiQzPYfm4DYjaLmytgVOxetvPN/nyvSuzlAmeSGBzMa1vUQBTGj
Jcm+Ly/FHXg797XK0XmCOrklJfSjs6QmCAd2lEfuDbKbwiVxOJ9Ov2aQDfpqF+gl
HbcrSZDT/NT5oEwYOU/6cm8+Y1uEr1khxliKw7dpOgJoEhLWj9aD4Fadq8HSKEig
Eo9SCb4cglqpw8laVhGfWUfPBOQW0hx0e3aQN1x7WYOgYghfhUuXwsmNtTVolui6
p8AOHBKoFNh4l/SFh/pxLL4+t8DQO+vKab1QZFy5ib9wYIrrEkiudVj4/XunMulm
+OGV2bW5IRmBlDRKM5L+RFm4Q+TPQtIWMmX37TPqt2BiNw9KIJHLxBO5HLkDoATM
N2VtbMGlfPpH1SUtGuncix1xjYAaDrd93oszhr5dPXlEYzFuX+a1RiGEnPvDQbvp
aD5/Vn1qfbIgj4iBDkSZABoM29Je0yEsHjyvFiVZkHtMnb+9BTexMBE4UIZ1b57G
n2sspCJ8DnOlylkIqOoEmHTqPG4PTOhv3OWcDsV4XgLtXJxLJb6+Uy6l8En4hD+S
Me0I5w3ua+Qw8HFGnCzTFmwv5mZZOc5ayU4J00qeaF9j2GssRlPOddrZ53MbNzts
j/lHnkRn49sWBTEJ0GWevdJm5aSRk7nvMkdfCPCe9uOHXJNRI+9jBASln/D3sKDR
jAdBGkw0NcWxxpmZSwQJqb6HnB/Ma+5GwJBRwIRJ1LUmPDaxpE39uFMFlFJFUpUc
Rr8/Xmw2Xzd2ZuZXw9XRHEIsxaoY6OD3HlXEHgPUdQJIO4qToLATHa7VvoVbLs/l
n7h8XjF8mAHmE9cpDt2OcpvbjorojVdahRccE75CynQciX1OnNnZ3Bvf+hKFIdnC
LoDrEzwpyqLi2bKqXSWALspToA+ZqbzWb1Tq803URI1+T6DLz9JyIUsR54Q93JVs
7OQiNA7Qda5fhHWPeIoa0r4xAi6LrispCizjsfpYH75grF4OK9UI7x27AcOncW1B
YZnCaOskZfPpJiXKGtrY8S2PhvjjVtU4UPkF6Rs3lKaSyPnTnpmxOXZ2l5qsLl8x
BEmv705aJEPeasZgyYlLtJ/oe1ZDaY7m9gppFQjQ9M/0344n4EKBlcf5hk26p8me
/55+vWbGilGXRWzm3w+qrHRw56RsUK+y8dWwtCkY6z+b/kbrqBnWja78dCeU+pZq
UxvYu+vaO8ntXYC+/YJg+3knyZ+ujP3eDzI/VRtI25ZB3K9Fi6SY25wk8W2E3uqr
OR6rCO5SVBIb5HA8eReZgvX8zneZotPtwYB8jS7tPcgRxw4+7BvE5HhJfYtEM1fO
bJSStW7Gns3mltkEaQ3nF+Jazt2qAlrO309dBoTJZDItnunUulVMZDZEtdyvwPf8
tubGBY1Stk/WPtArMHwBcqkWgOkQohtsYqo/NHiQd1zOCdsDvgQromBVOCGgo+DB
1uj4zAjI2wB7G2DuCiuH4mWX8p5dwPr7WAMYQ4OvCdgcMGhiJLLfHpKPzdKMAawR
ZNDM+7jl9JoM6LcHoxVSnSGmqbu4It/JEK91gjC4O0Uyysgp3nmcM5FjX93IU6Za
vyI/7V1PZv3CYtr+cZPW5TkE2CqwpcfIQRl+7rvM2VCgug8sY3c/qMLxiJx/E35/
jfo9ymXSGRKNpddNP2ef+OXdZ5bdqTwBI+QOjlyehLvWKxE6Xc53QFN1i8fUhQnt
fQtgdeO8yqCnQV2ZMA19hdGsiCtgytpiMZQ1kNWE1TbKDLFy6vEAb87AdFBZAZUR
KTSbNkys97WDV+JK4Ew+mOPSx5n9DYKp4RPEwSG4MNr91OXwCGIFgpZHLcfGIQ0W
uHGxt02KWhrc32UBVoHuvsuvtemOqnQUV0MQDTFHMuFRIeMPC5EFpVTgpUOq4zv7
uHcRSM28WhCphsb6WBh4JGF5nmaardeADn1kf31MdYmpe4hBtFsHv+Q+IM1rZC2A
Vga4OtvtWyFUEVNkMFpdzK9Tbi734w280vuLCmDD+Ih+SDqgcT5URYZ/+HkdSKci
v4THnXqrSkNMuK34x0J57mSbvHZOQy0poo96RrDXyJsUieE6bz/FQL3irwWW6XLO
vlYgpPMST1yI8s1ChdZ5S4gfI0zTHeDlCQrUKUcLZfC+kkDobeZsHA5Kw5EZyK/a
RsNPamO1XI5bQtZgV1sw5nTRsMzbGfaJeiHXln3lCCUyvRYCmC/zgc4zt0B2I19z
t3mkljum7sf7graHkCfW1CSbFoJG2JR8QGQUtOfTsO5iG0rLZltfchbHYD+zB/vQ
faqJhnNOomlF17DXTLMk9yy2utY7+VCnN5hAXcHogRz15DPfh2eImJDhQJhkCg/O
xtyKRTL+HO44pkLV2L2RinUz/jvUALjeJmFS1OI5idFksNqfKic/8+MVst18duEK
CeQSG9HY9y5oWKytrVajjVgzpCdTjLbq5tOsoNnVN52mRq9Qynp/XbTMohjddUjN
OduDzrRMb0afDHze9CLzilEBiu40aWFbvlIltxfPQm4nHOToD7TIToLkFvvoPH2I
zrRsH5W8Kc8c69sF3njWMaYruTaZPB6dpDsxpc2wzc1jfMEToR3s5rM3HVioexeQ
2r+U4DBTZUCBj2jMg4ketLXF7W0xd/AZFOvt7M7JLRP14//lUWgK/pzyf3KmW74d
Tr3e/rLw0dUN+tHs+KHuajOyLjDrblw5wjIRBQrnWPU4uxr98uMtJE/eGt36DYU2
oSAzwKvJL8j2kWaxJKA4M0d1U1Ga07cGpHQeAiBndZW6LK/rMBST008wFisKActr
qiwIrbImg7GpqlZTH6Ah9c1ObzW56n6m0YnRME7dG06HwnOEVOHcZrIehcKSbJJW
XTlA8RYigY/yK1G/DkiQac3Bv5lhldlGSeV2rg1Y/bZVwIy89gvs1kF/qOCJj48+
Vb4ZAbcDY9bQkgHL2opqAJbNOI8/AFV0ZPD534NDGNaetO6ClYcvQxg9E1L1GYdE
a8A1DvcoAVnxpzKna0n3fDeM/16gSHC40gq04GROJ44t8ZVIQxu7dZwkVR8G7HCk
UoVeLDc4VfMPb6anF2Ww3Hs507LlYr+FoEWSEKxVqiP5KwKNihmBLvOMOXkY9YH0
o0gSm/Rufz/rhWFxhNlxS5nSJ9/qOikMs8ttImYxByUP/9t4kana/t64zXVzcNjO
reU8VYw7di7NF6FXp6Vj1EeEfKELb+o3UXyHtSaylwx0JKm9QTge1RWkjLnlwG9G
N1UIKD0JQ35nvIiY48vI6Z3nIuKEqG/DdQuWQDzLHMqjYi6fFt2WNH+fazUs4/B0
BKxyjJJvj3/Yvd1tJnpUa6cK3QCjOoURMeHtA3QLDmnaNGz7saXvbvZT5Jx0Yzuk
Tk8UD1kPmnwhDAHRfR3guQgVnJZFhym9fdhtKA2thFpumhwwVVjhOZvXC4gmNlaF
en2uKOZ2kG6RH+AKLRyAEw5FtE934ZQRNM9yc/YtXiaPkyZmB+pyEf5jp+eXAdJ7
Uzj5EwCjSEsaMSkQqoOUhF8En97auC06HE34kV+Ss84+DGs98bFExeWWpDmsQWlv
ja8jgdbexl/zIKdRB+jOXmzQXK8D6ZYlN8Rt5ZF9eD7EirUUGobU5Qae2Kup0zJH
clKrhI2KpuBGEPxLNN97A/ymxfJVmk6c8FucuJI0kGThl3WshkYsIpmrVZZIQGBU
XGsyYOGe7yZVdWNl+v/U4jf3iWJu2g5gckTkoLBwzuDv4BCegf/X05gWx/W8oxDm
nRGt77FfKNu6PTrM7Fbq2nBa2hTckex+P9DcsjNCA70tYpEdBATcIwjUx6OK/gfl
iJTl400/hPJkSq5aNtRvwLCoNpeln1ZRyriTWXMfxweTjxn6kMS5hExDlfMwphYf
n99Oc7lLQN/+Uw0450yZF9k9Rq7h0CaGkNoX5jCEQGhKZIvXwZao6BcpT7R1JkHg
xIihMxnanHf6dXsnTVMNyj/Ibrf2xeZX8pTyig+qxVQWbRuclaMIHMKq3mlZItpE
36N5y7lKwYfnGCoEdZOryiSjykaYTgiIxlGF+CXfa1uXMk4yEnxsPTOqH5FjKcf0
Ox5Z2HVHQmIB34FUvNqJjcv/ToSnBD+F+xGKrul+h6uviC/vCg5ETHSIEpsBb2Ls
EAmPYj/EOtdVhjoljG8pB+bO33kXLuM4vOqsPiwv8WoMGib4QV/nMYdgTL5ZweUR
vj+xHpmEhQHYv705zPBRhlcSymNjCPsWHyt1WohGA+u9SDPy/+nu22CHjU1W3DmE
EdwRSkpGRrpCM6dF8/yZa4ENz33fFnmOwobjWQMDmfp83JWG9xccrkV1R+CZfjHx
ZNyGlISgU5RXHWE9Xz5XN6oHQIehM3KyvQRkrlwl/hvHhxYzzEb+zAOW6VGENzSK
LNask7vIBY01O70X2JGdrWHJb01x5WDZq6iFhwctKK33eHLlDk0tm5VrmfW2gOZ0
BtbS7HT/aWXrXDaUBATQr0EVla+3cu4sUUJydnFGW2W+ktWRLhDSPN3ZgQNddGx2
GEI1Hu1AjAbJ3f/iIRM8BUoIoGW7nq3ICLJU6PzBnisSkq6O0EgL99EfsO5+1Wpe
O7syLA9MYobXBbbR5Imz9si0aIk0ykVZilvgcZk6eT5Myx4gsHGoAsvC1ZnNjdry
WElavSZvJ+cg3aihkEapNqQrFFZdN4Nw2gLX88bA0iueOr+bWm59fXWV5rRA6RVD
7U57U2ewug28rYgKR/q/vFRkldBZkHLoFW+tpeYi264M60ouQjB0TL6AIn4Drkj8
TXHioUkpYCQR6Bjn6CZA53DeiswsKU6d4VZ07k4Fo1k5R4hUC2esRHNwGRqqNCnP
nnCLE6waO8iN3PUQ5iFxHXm9LWv4qmvcLgpZcjCOCx0bA9IH7hXofh1NzG37if6+
YL5/Hf7o/jSMU/nNQC9SgbXaILoIUrC5jJ1dbRpJEmmmyUGYbyjX2NJ5XNg3FrPJ
0M2M3xhwe8BFQocuw3OtMi3YbHqGLVBjl+/3NfZFfLFavuDJ7guD2vZFWQW0WAPN
LM5iInOfrsChtUXVk2zoZP/nPD3u3xjdOtiMlETJNDGZ+XV8c65nr8QXB9i2J8LM
A7nFmVEBlhu979GkNLMehdcTieWoqcHyr3mE9mNDTU0=
`pragma protect end_protected
